// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
4SZwofKfGpwkgmY1lWkFphFootp5Xpa9QaPEpI3znBR0aubSuRQvThqfJTw3SN1T
PzETeIyPVb2pd84b/hp6QVhdGvVIkWhsGNc814/GHqvACFU6HZarsL3XgREm6q99
wH9DnomRPPunNcREUaVR89EJNlcaMAAB4ODWtyTO2Hk=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 1080496 )
`pragma protect data_block
NnPXmzGjwMfTFuxx9dcLkvXF9htITgCu1VRuRISRv6Db4FB6wclaL/9qc4KhSdal
CX2QBI1bv4suGqZvo0yCmYnV5tdG+p4U7bXU9mnX4jojsAysOaWIVLA9TflLS4Yc
irxEYFyqvJ+z9Oln415GJlf5fTlgUWpW4G7OGa3A9fl3a7rnbhBBdI3vZf+HJtMU
rmfxkdYj7ufenB+d6gqo/nZ3r9I06X+cy8w+uk6wgEkdoXlR1yJ4EUMUjGjXjwIW
lrpTZvb5LmlVEJgcx/yW31n51gAoVwK/q2EyxhrbpyGv1VKIfM9OHMzJobo7rsR5
eGbpPbEBOmb7tuQOYoR5SIrhZ6GlFiPXLmOxJBMbzZjOUQ81qECmHd794J7B3qnW
0mwsiHLioo0eV0UAKh6Zwxi0esq3I2PUaOGv5TRbp3xX2erqyfcOp/nBbhILO77V
D0bCNjG4UsWrHhSNJKccUon2Jd0AvR1490uTMesPm5jq6H+2cPf3XNkNL6ZvqMRg
Edt+Hj95HL7YicF4UU1fR5P+HBeA6g/T2Q4LhzfQI3NCTb3AYDQv11d1Od4L7mOf
g0f3t9GgwiF4LSOAesA8HpH0+w70LmeeqZ8vf9gm8JCgtu9UmtNKNVyXQTLXZXGR
4ph/jAEOemS7EnGX8ZqgKgq+7ZidKu1onzbh0QjHnMJv5al6ncXQFPFeonKxy6c6
1LY8U7oovzilWxpKJy8c1P9Gf/2PO8fkSiVDm1QAN/sdpeNTkGJMG9yjhrwLLcHd
EYS1SjZ1Fgq+lYLfmDDbc6Qt4tTmU/0WtWX3hZ2Snm16t4CCO3FPl/lhhxT76QB3
Ryrs/vGZnI3iav0+bV1fNKAT7RbJ+9ZbcifAC7dTRB9sgoVtKd3ElXGIqIbJ21pH
g6EaYZXbQuKCCTGhKQAXzwYpuJnihomavU7KXaRIISL82x8M+ai+TiEW28F5ZRfp
EGED2Xgx9xsDpZH6y8Ikrf2HQZkvfUfd+uqEG9E5D0QFoKOoAESsIqzaKm1bKQ7k
ulDwwdGZ5aJn9y+Fp73qYSwgIHrDO+KaXMt8HyVYvxkTjvTGIQyJvDgrnra57QUQ
VSD4BuQhG4o2o6aoen5GwuoPQ6t413bcE7HdCpEBkwJMlYEJoIJHvSIvcpDCSRfB
4Or257vp8f5WlNFU2vaAH5bnIvx92Sw6AyWMNPbg/I6i/7AGyBCmpsL/ZCSp1+0P
D1OaRrq3nfvgcG6E4JB7Qp2o6mS3EW9NMUBpzVLedpCWnwVbd7Gh3aPYd5ieRr78
mOzPv7UCajVnovN1bgFTc5fCL5+HGirshi0NutxTp7AU3F1eHmXSWg9nzR2q6pYB
FwgWqBJP4A6mP3QuSZHFu1l+/mVXP4DwATFDgIw94o4Og40kQIebfm6MLkcCc3Oh
qoE85HhDBR3gUmrvdJAR9YNMyljlsaWjF7s5oOfdovmXftORdCQBC9ra5FmOnmiG
H31Uc0NwOJbZGP/UXP3kg0Z4Zw22wK0z3oT/7XAjhcf6qZho+fV5hLKgN8AUBjPc
+dhswo1ImOHCFwZTkWK4u2BqVX3BaGB8PsVihnLngmgjFSlrCm/6UPu4tWAGz33A
jC859j5zpqPx2hj0I/Dnq7Gb28sXU9pkynVRLY2lw02awWgBTGVPw+1nSkzkNsyP
+r9PU54f3AUOOGQADC4joxWpOlstboz9qvG2eOniWL6USrGEiJoQZRSB00RjsAvC
d7p8ZDNjE6JsNY461W3O9ZqEWYOj6AssMq4HIQHVua2TzQFQmVSZH3y8a1678SFw
AiA+uKU5jmXsFL4C1jtGPIHZYq/9KTMjKeNc8MvyIlozfELqQsCFt35dbEiMg1di
gD+JLJ95UfzQG7p2PjCuP6r2RLvm0FviuvC6LvFIvNPNPxWw9QATpL4+2MzLNIZm
hYQRVd1lNjWvIdiRWR/GhTpFRQY290d4N40sMXO5V+fP/SVMSVrKP+tf4GDfmzGz
NhgQjH1kYt5nLyv2rXwPcwSzibBZp5RYVsCm66Md3fTdLqwauExCm5KD+d9YihTr
hYTrqRosoRw7JwboRI2NMy4j+AfdniOvGCAxQ9DdNUrNxn6uzwMtz6WfDijB4lii
cLRn/3I86gB2jpi/SkMq/Fv9rM+7bsmsJmF9Tln0NESgDXqCGmZ/eUfzXduPlKer
JinTRqHQm7/+a/vTN/Fu6M52d4YK4CecOYz6ArBHsmRuv4+CH4ML1Jjw7G5hEH9x
iOdzYNABA7rh8/H4MoTuTb5ofMapofMeGAmx4cxoWUEzjCpdvnEmAB0LuaDNRUGM
15k4yoezTx/lU2Ea+OqF6W/nSXN5meqh/77DmiYCvUjyb/DUkYxtTL/sOEEzFbug
yq3IS+Ow1qyYRwIxpddUHNuRlwuVc8qa0a0ir48ohbRoi2Ve5cQRLksp8s2BVY/j
DZkGVfF/EvqA7crQm7Ko5rJjNmRLEK9o64DZcLJe3ULNHMaHIXDRXHgfP2oqgnMb
vRabHg6KkM0RNZvtFAAgIXyHbjvOGNbB2WVcsrfAD1hKCjRJjSbsGhTlEEmWcIfh
zUOxru0iI+s3MeYg9Cc3QXgtFNezZ3mKOeo9rvEPlQ0I8gHYhcrFmtVvjNPcYlgq
p2q/a+xdxJBQTkaMpRzxV04wnoAMxdU7mvn8r6QZ/y9M90Zq+J6jSVBV0zPYxBHA
5hVtn48YRbYtSzHU01Rzq0nGEOt5xS8diSUjoyaAmW0VNzTg1wxpNBo8jdrQRPiw
/yc/oKi7FPirsf0BBG5JMxTB9j9FUcaprCd6Gsm99xkVDoLzOcA8carPq8NeBt2Z
kLsO12HQemRc5Ne/Un990RswGf0rN8UZ8c0VXOwRJtkEDb46w3L7tn7FQZQ0GJUW
Ek7pYlipH6QCotWcktsPFy3Gig6UxrKKz0xtYPrcWmfx4z6F08Ds2hkAFs43CID1
Pl/ryrvtu9edojtJ/ulmn3oJ9FRq3I3s3TmcIR9xynii11EjvE3Q3z0mITCCXO1Q
EyPMqcbTsgWgrdYvzcCjR9QcsIpTfrKhv3/73FwvQI0qBJuOk4yUcOwKCttfrCcT
UFTY/v0rhvehPddxDlA196zkKaf2brAFyuYY/aOEaZfu9hEn6+6Zie62viyXduI4
cQIotnCli2gjvOk2FJViEBG5blWYjmcCS4Qt3JcbPmC8CBBOU9XcVWPYQ4FW5E5F
0rNyEuBCodO4IMjJXzfrZS3602ISxKvGYJT+Fv+2ffjMgxFbtGEWUKHoJIAEgw4e
ur4jI/4hpSdGnThyFCn7s2ggHu92Say/NG+bhIuwq0kzV5A+H2CV6WVVv+KQNGSH
NVyAe8gf6+K+ncqfakYRrF5zrIbAx4rLGOwGpkogmlodorAQF7whj2KYmEn9qQED
h3bOl6in8438Z47N+8ANWnhuq4bfdOFCeSTtRCnS2L710WAAllegeQ2FRg90sFS3
j0CMeJHuHxkrJRPrc6x7o890FerUIVSyCczYfORSmMi1PJ459t/BOlmHaKWaYwff
NUUESxHiyZj2R4c3/paal2dpFu1+6jn6WpkRmBnq6SQtcPhAzo6yCEQF51M+tnb8
UJEkNBol2D3U8oPKWuCz3tqq9MywyJ8d8P6cj/U69mx357CuNUCErPbaogKgPxnG
rYryWWxc3Y1gHpCwankKKv7IoQ2Knnf/JtcLho24pflq9Q+z8VMXGLVV/2095M3N
0W8pTOXpH/NFYbGMtLyIeR/iCQwUyI7jAyntGsvUddGoDMtsJYFn1J4wBptpa7l7
ngU7XR0BODF5xm/SOzwepVE8fpVvnDzxdJ4W1c8t2hxwWUuPuBr1w1UR3vYC7x8m
a1i7UvCDWzjOekmBZOmDkxirQI8xRwi56isVSpoEez/gcuoA9gdA4W/OEEKV4v1D
VOgjK20IMWUxcK38J/bCDzV9b9s4wN1FJHrYA8/wq39vAK2iaV9H7o5Q/pFsATcK
um4CU1tj+9QxK4xbfjc5GguXuXh6Gz3IsER1JJgk0W15tIxr7ahFw1MlShb0+5hT
qw/1iesNbcvT1uZaBqETbckQd0MScZ034ui6iRoMquW0LFMIV7eGXtpg3KPujEU/
5h3K4n1l0X3vzNijS8VPuKQmyviKbA20S0Zm+0yO40/AIl8JkrJJ8H1klLvkuWHG
RT+8NBX+AT5SO79EQXEMjFIkHVJiKvoUvUZg+DgWirusVsRTIGnkcoOZhDOxqmNS
4QI0jvdW3EDyWFw3FI/pnIlY/DyuoAZm30Hhh0v+VZ3x6RuhiHNR/y4fV8KVzFlC
x0k4tMd9k7RbGP1asA5ABc1pq2JXuh0JUxLHphBTLMdDEc8ke3GuFqg33CD2ueNm
9SaBM5Tr5pq/SMq87DCDmaGIOnfQHEziYjHNa9xnscxndGCzg2U9Y78kq1MIZdrn
/nJxeDtyorAB16591vYqP7zsFQ/SuSoSuQdV7HPZPQEve+3iJ0m26PB2JMEi1dul
5XU754yUftE6c96F3HnT0EKY/WonebLW4Cl8u0+UvovvUHFG1AxFRdUNMFwfgQFB
26QK41/reJSNe4I9P1esbxV31TjKmL/D3PPfeKTeYDDz+FQrX3ewNdmT8z8cGwsT
AmnjlUzS1XS6J3f65sICF+yg9v5Ko9KcRb3e2GC/GSwYUOrZiSDGbf8nVNRKmCVf
T8UuZ6jNzWjLgBEp9rZBukeKwomyAvLgswnM0SRZiZuwzq077lsOqB6E46uaSeOB
+OHv3zEz+xdx2nsgM7iZzttl7H2l7LELHjNCzxoBCSwyBZN5uHJ29slBqUzbXkgY
UiAogvcIDU+bCXUvTG2BJ7zgLuLFDFqkWcCqhbcWNIShrJ1mhwlt6te8Xmy/tw0M
NxuhHJdhp737w9UU+bHj8HV0McejibGew2ZYnG3JTqmP6lkr2Vb04Pgi40ejFjzf
gc1KxhCpPEFKiboUVXTkaXYmQYwq4gj488pcp6xvGay2z6N189ijID4fOtve5oT7
HM10p/jgm87HNH3nh3lZ7oQVUtzEs+EwdhoQrUiUp6eunR3+XzebgCPL48ofHgaO
telYeiL3VT6drbPKMuVnOachM7rksxenJsFmEEOz8Seqv01YyAiuD41e6iWdcpXT
Fwv6pCVPZaz8akW02SuDn+MZUf6VrzZukwe0v+9ShmlDG3XaUHPMGfFAYgxz6yAg
8ykT9oVx38XcbswdJvO+jPIO9OwA86v/fmqVQjMyGlfVED3VlkBiq0J5cZ2Fhnnw
sGDWxezTJ5FihhAHpbXjhyI9kzlRmEpFKatuEv6yEWd5XKwd7x2q6KrrtKHs/wyC
9tpg3L53DvMCiRLRCKQBFWnDrj9rjy96uvaOBSah3sAGKvQEzFxgWEM9b8VsveIj
whZbF76wNTWgdouwDTwIwJMF9BcNXbxnKa9n4eq6TVdV4RhCN1GwPTJ8JPMuQA/5
9pddd/anRzxSJ8gidUdKgfFNsTIyDPAgfBwqoWJErYnLz1wxYbI+YBHKnhhwWAw3
hbzjqXizmtjKqoTyB3iPQDQUiVSIG02jR91QxS9f5M86dMLrcjmakuko91eQ0Xoh
JrRI5HpCHAC930ZQeV7mMBp7HjYkMAPCdTy97i0P83yH/y9g2J2RlRv/Boo7BWO5
QbvwbQlPetnRbxRTxuAyb5EXBgaw8vkump6Cppk4Rl302GJoaj0UmNZQHEDsTVTz
gahFcF7HJ0W0ogTpn9AKnykpxPDoaYla48LEmFJTfSLn9ics4hACr5x46ZiYTP4j
ZHq0JqwLFfiNVigw1WFa6go/QtS0J+Ly8pkRRs4RHOriiyoJ4ForCaNVBnvU1lIa
qiR5lAMPXftlZooY+3Prjwa+LdkK2s/KKlmDVfI7fc+u/CKcdu0Otf5sqGkwTuAF
00E7SPHluIeEGTpBMu+IYIYoVp5F/QHVPlUhwvhq8VwCuMgSbAHyYvN5eT533jHG
e8boqruzApMVuLY82hrevQlfalEuDtsTHc2hlQ/Izf7dp1nQRljxS0RcNDoXQEEG
0KtBcBX9Smv1lC2hAay3LSS1YFRj/+N8tOo9S39FLmQkMWJImvF/Y6XDkmwZtb3H
WGJ2KimgAgqY5vm0x1Orhdwh4l/E/eRMENatc8YFOhf0u3eaQkOw9L3mmHqIRoG9
VrcG8CT2qSwLib5I6iM6X7VLVVg969lAW7OJeX6g/VY+WZDUJPBOCUV+oiKek0o8
23iRYx1nlp/J+BjdoG4RGnwKweh2UHL4rmv6oEOFfGjABOpAB7gmt0bhzQFmoRKB
+EB6oXCbNcmsHTWgYCYoJbAfJarcfph1x3ipavirvxUG5NSr52cCQM9nauZdEi2n
QyFewVsEwRP6VRpqVNDba/iLhv4H/1U66qXmS9mfDu3wYajD7HEUG4eHQlOEHwLR
/FFsYP0I76CJM/A/v7wHzHJiEWuZORJ4dNd47JcA6063S1QIBVh/+NQF5o4pBJF0
Jnh0rPlzEontDg1Rt9QBit3GWJvBrsoNV5S8VH0WPEeIirsyQTVboufzrHZKx12N
3r6KWvm5qNuVQ8fO8pBSRRVqF6pUF2dQadjEkiBDJs5o91YNG3r8Dl4wZLatx+lw
QG3kK/8aIvD4kaEh8vCXhoCfC4FWHEqB9WaSgHL0+d8dLq3Ox9rnKIgMmqcdmXZI
wLW3AvCucvst3PRcFDaOPApefuLpeyPUBafRIaxcI698UOAbekVtlAKPsNCnxaZP
cZgUze2FAMpeh6wUdSJhw32+0P6nTrOSbuaymlRzbbV7mLNP5KY/tcl3TVwRaH5w
BAnr0KGYyVnXiXvbMWcML2adIzrAupntFT1lC1qANC4PGO8680FD5Ab8bD7msBYG
+ZguRsueRqsyGUDU7vrtJzBLF1PFq4R4Y/dc73+NojNJ3UMXAYluhnhOGCwmHZwx
b8mFpaCGMqKLbgqHTBVS6brGmzDyKaprhDwNNegXP9vf5m7Dj9zi02I30n1Sz8XS
SXOKUR4X/kFgBR3sECoAGgBA8l2xmXMcPDoDSEoagk/wfObSa1+U7UAF7g9Tsv3i
3qHoyHIan63Y/MCZlTO9ayqu80miYYyCkvhQgre89OCvXlabrgqCM4yLLaWZLsvP
Pwu/fnXZIfTcx+f8IoZR6qMj+462jd+zQc7xZezqyMb9LQXGTbbXOgZ3UpCbG0cW
hiOIrXihDICyTMByd9mn2qB1Oa0VHJHm9eZX0ffh5CTbAKOE3vNOrSfBm+rzJnJ/
KZ/BHyqyX+64Ed0nXbDvRqBgpffkyclTdvuQ6km9r7QnV+cNGXhuo1HVRjoAqq8B
+ZxSfmrL2MsnddOxwK5KTv+KXLv8NjeZ3CPvBbb7mQjq/n5i/0czw/UzgCgyFvF5
e8omdwUdm+Oaw0vqt/GPXzWN3Bw1evmRk/aaIhrHL+nap81sEkhvpUJ6YDhn0/Ww
9El6srOjc/iY7TXfwSRVPp6OfH1vr2ob57raoyhAGgcO3ISRBbv1VJkhaSFaYNE6
KrVzEqQD4UlS9NouDhUktu2TekRjzkXBtZJbGmsk8U/5m4YTQnX5JroIllaV/Csn
HT08jHg8LPN/1ilzsk3teZeEluHSo/TmgM+uNI8CkdmTOFyNAyx00qwCPjZ7z1hx
79eoB1dYTmTeXSOrl7shcEpty/3h3hf2QGpBhdLWcNnF6sk02AadYeVl/irnkKNs
hzxqZFH5d6K7mIqsWh+95RwGLd0EwKOWig369aUkn7lpvspoKLj1rSn9jhlgaTB9
seoPbIBSTTQy5gQWDJzWCdsLsWSFaMzJmh5wABx30ckeJwJpJGusKBU6qipTfFAs
wBRKXH5kyp9XY9cVIVuwoJ2/feRxqUvvsHf3Y6PdA5h7xiVgXYMKHoQdmFd4fiL7
Q/E7PSDRTGcbNr38j9SW7WdtoG6YLC9gTMUJBCpFwjyo8apO/kVc2BnCckyw+56d
NTODa0M8Bhx9tQgVUr5aX1YwnOHHYBEK3hZ0tJJdITMqVFs7C8uz2hbi092x2WcT
1XB3qwKwB+pVx/iuz1ESWpomRh7cY+L9Uouvj0jNgbuGQkXRGsxjJg0dDPR/Jgja
YUZ8gLKlBQVM92FtQybOfnmfw4QFRGETksNdOk3rb/+Zaowho5QYQ2GFYcvrp7sb
AwIncVUzJ5leni+jfgNEPw5zsy6QpbzUn2SBfc4O3XlAu8znzIClG51UAbYN8FV5
4t71gCmpRt8d5yHdnKat87xYuGsBbISEYllyo0vuySPAzqiiZ+Ll3FtD2gOE+nsF
RAK/RviqwgD6kqseCSxZPYZ+4gIDRCLBpx3SpzIR17HJZopSTLjU4tFbY0q3EhZ7
9Lz5CbjEG4GKGHE0T95pOAQaD3wiKVlDxmWnxbAPoEJMdACTo2v4cd3uUPIjWKd2
5FpW75eWRl1U1N24ti8WcwbEH1yw6EHTlkg/sp/6KD0N0ouYFkq21ML22ssvKRPZ
AiIJ3cR9JPPHT8N+S8rBWhH+eCEMIEQAuKpp5mI3ykJ6E9oN00EESl6lkZYXavzr
56Do1ci6ngTJntrJLkwhTym6qqyNyxh0F+OJ26/Pz7gOpy+pzf+6qczjMHGgRmRg
PpVOEREAkzPZDdx49pt3zycOLaKAsj0UW1ZcySKLXW2D4AkAlnhGcktJyP6Ulflc
0M6X7xc26NgF4bpXOU9lG3KzojmnqDWbCtgHNltJBFIcGmZE7kkb9dmmA09HbTzD
QAbrVYIT8TtCXES0nlMnckIpdTRqHAL+sO+qeYqVLS1ndX9nmh41nICWXdBPFdZN
dmrozBIFf6VUXn14xoJPuvYPrESJpXeChP6Gq0Ol0fIlyEMMAlu4bs/7vamUkqQC
QWX0s657D2bRnEOKpdC4aDpdTpUfWpKv4gI9FxZzcjPaMeqVflGCyHfetmV4EHwW
Vz+qTT330iJnCDuKjPTkYKlqnqBvpilkbo/+z0XMAkEhmp1XwXBDhmpi0hvS/huK
/x+SAX5Vq8xsHzxVAYVNfcJ1mBXv06T+lpMzRcv6S7b84yiNue+hrHglu6d46mRD
9+OrvVXOHi8A7EY8DFpCeLNA3dRgU83P9wEq9IY6FpkqgRnwKXyQnwa71CBarBS9
amzxM0zB27jTaMhtkUzVXL5xZ+VUWdR3K8Ve3oJoKVFd9cIpB2OIBhDSR7pcN7Uq
BS6p9QJEfpZvdxE7iLHGndYusetKrNUIVwVXlfHnbemVXF2fg1MP1ksdKPbmQA3s
ESSwGiBnph4FiliefhYIfrHONEk3uxoTCbGi2xMU4hTcgdc9Xlcv1s8XPRrfhQjR
1gghaKYk48jEgthi7hiW1gvEZailEjynrDe4HyOg6Nujh6oZ0rszm80kyqflOgzy
qWFsjLhJc085ualbhRW7J+RyXF2YY96LFRp0XSBoKEYjZRmxTZLZTS+1wthH33Eh
OeAuhSLsUMtgNHP2JvJ2ys4gnbqF00SsoZFf26Tt539IsyZq2Rgks9CmS92Aa7Df
bA+2EgT/JmKzVuP1N5oSA7lsqb6AS+IyhS56NbhpE9+vXIdQ07QJJ0Od6zD2ZeCQ
HDGC0Nz7BZ/xew1B5I4Qi1J6qla1e+5FSOFaIfrL6PfQljkXTr1UmlkwLeloHHiz
cXpGR21avJdf6AYTd0uAGFM+w3UTcQk3Oq8j3gh64NpXs57Qn79SdKZNE7e4jxyN
Rcfl4jltFaIFWzbRprCcv251WOkWt+LsLOBxlJecsioxVqqZE2StO3NtHimm462y
hObe91mGzTxcVayASr1Dnx3ILkuq6lF057vuo2rT97ruy6hwozl8jfvm4WMdJMNC
rv2O33lFmhiwcRSoFi1rSTb57jo+YIbHMYvn4oDIG615f2erzdjX4X6ORClgH46i
UAqqkwcmcttgOO1WFXyyQ2BCFDI1gyYFXB8prXCRLjStwLlv4EXeQTtEmUnYJ3N+
8YmfkMGiN6Ed+t9T7b2wVbMOzNf2p8hpFuezkXnyvoa7fYJs5TbX0mWNoVShid/X
BE1GYmyBkhp+j5zc6X/QfeVHuqouN/Uk7NgzE/HR08cNPCTlaKN/1d3r30pJNqfr
cpPUoqdL5ViNFH4FMmGL9egs5+n0bOy0e++TBT0F7DyK7Qg/g4JFV+viVYvRauk4
DpwozyoBbVp+j7D72u6FyfCLXBl2qiXC/mILajU7PvQDdyvKWJ9r388v17TvtVeJ
/vsXWPKdlq0PydrLRjQ6g4deO7LOcGmUZ6I/Kn4895E8GHPK+dUpvigevlHrQXOM
Oz2TxjK4XvdJCyyLzZTxIwT72kRYZ7xIDYDEpw0EuYUOW94AsCo9TJ0+jXd4rI1A
uSJn9GqWASqOyKvfCxiPQqYDTA85aYZlGLUUM1CwtbZ7cMkXcJdCQWmy7XVBg1Oj
pXRREzSiaANrZeqS6UOkgo4b1qeR21C457hLuApvFMGCH8IPjVQBFS7VwdbRwFie
wYoXd5nA3MgYkD3wzVNMOLJyeIID89Tl5YSkix3b5oNYk5qFseyzufS97kzh6N3t
EvtzLg25/02JIrbd74hd15GosV6WIAVyoKLhTpqdK0jdEova2bEzLvKAEOK6D95P
+9ZnQBIn3B5S5r1icrjOy+f/mf5qM6czq5zfKFKjhrNE2vwSkwXmAhbfP9NAY+NT
ZPi1LGskRPgRjIjUH25R7KVXpxszn9vgfDrCixr9NSOLoOZj2WAyboQTKL8GYils
2M6dIiS3IDyVbUbCook8zM4NUDR+y0TgS1YHCFvjzwdGVOlT+uw3hzle+jU62/Ty
a1GPWFxWYdjOtPrp5g0c7MTHzwDrwbCllDkDibXFJToetFZkOlXfk6Z7c6dQnclY
W69g9OC+osHf6MVYQw2TPlCddZy9lvYX9yqHLjNTf6pEbyX5GX8mIysL/PeQHk96
fhUnH/NcpOj9GKoUMyYwSBCjpy4DA6iZEZSqA/H7d+NHb+YbWDdg7mz/ggweBs09
rezMvo7Lm6OejLbKqi8b/zEt9LhkDw+KeYAoJQv4LNuugQaDBml+UMMEJP2ZWLDZ
PDAf5Ow0qSaoFXah6EDVlPQT26LC/wmsVK4SQ6KA8FMcH26KP9Y1ooyrQ1ZrKKUd
miHIiG7kE0dN/olq9e2IHtq9u3Eq0BO6Cc7/hGw6zIryyINpRkSK9NKIs4ocjgq6
0l5eKpAfRVDhmoIrFVQghwIiLF1e6xuxq7Gacwh+NsE7PWV9XC/SP/8B/NT3VkFG
X3bxVP3Hu6Vpi29JT1gs7B4yi+Ljno1DK5Lw65bozs32QRAmq21suM4vcmv9TenJ
jPHaT323NWuJZL4YpGjaKw5QqXw5X9j2qnBFERh1E7QvptzW0LX7QmsSQQDKfEQB
hiNg9U4lwZrVf+2cFlzWY1ByyOZ9cj6/bqNQFAg2Zwc5CYQc1/3B+yLz5DNjjLfb
9ZhxtI7XbKMxh1xkxfuzBGg35l6LTKchsaH1oVEWXnFqvT1BivGG9i2LuZ6TJF88
fqIVHUYyFqjzRLQV9U1K50wVyKrgN0jjAy/j4nDtw8FwfT6CoNfPaJMcx/H7rsPW
Vzy++pmf8SM8g3PPzMkOTDcjlzdKOhaaxmDOp3jsb8Ix5iAZOJ7LgCSAdyhevPMk
ukb2sKDMZAGQKnmXT4PFc+1Zb1TG1npBV4/RedKuE/oR5kaJmo2rVGcL16Ivofsk
faWKj01d6i2rTW8KvqIYOgQ8Izr0AHoeRKrSQ0Gy/wvhsqgCgiXErQHII3Jghi/Q
4N5AZyU+CQvlIZOEQztTIZqphIqjHuD4PIqXrldTB9Qd8QU7CfddilTQBxCa+DwT
/swNcNYX52WYeixYOKYtjV4jJp5IRwqjzPD54+QMjBlrgaDf797rcnQZDDOdeVMy
G3VwNa0N6LP4AhAX96ARSg/cuyAH5f3rW+xs48QySo33ZQZRROLTNnPF8Z78Vf3g
xr+Pq+DJZpVlrdrpGekMkhjH9adyJ1eQ9dfbAG0iDxhaE2Q890EA0gW/mL5488lg
2c/eKQp9moOlZLpu3BeYOKQ1RxYtIfF8FZZF1Twolo+sWPjS8LEJeI5aiGBVHYBr
sQwiSlpDOx0xZSeB3VygiwB1B8p4KlgDz1EgZaHVjO/5myLhitFKPXlvMz9+BoHO
JO5401Sj4wYeypZBQhaTTSpEFuwLW5bgQ32rWP83DD3osINo2v5VplpNNO20MUYm
tsValWGqea/wepmrv/eEYfYYwkY+8b2oQHzihDHvxzM/oXRDJsFym5e/mGCvZ582
6RPIKFt6bd++JVxMA0r0zFt7p0OQfIm7Z/s7Tmo94y2FroC5/alpqHmG/g4tNXj+
xtncbqixKASIVV2LPmPS7Nn0RBq+qvqkwZ/STHo+dpGzdkMBsdVWTnYRvAw8mkLU
e1En4/SgYxjTGifWZECHmFtlMLck3E/XcYlpofpoh9XwALbjFSGu+dMfnF25/zPY
gcqbj8RJYt/YKdg3FKnIIsT9u57jq0mVKc5hUNZ1bz9g427BR5/XqRHlJRWHf566
P99yff9WDuuel/a6Rr8Tv/XixqfJISUmlK4KX3y+cMy9sc4uYyRDOtkdZ3iCuVZe
R4Adl2WVZr0dHV3kEiCYj69Lk7WS0SRvC52K9lSyCbZmRMBuXzhiA5Ivbo++WblM
Mx4dgsOFh6YtGrQyJPzTRnxLxAWnB4oCh6NHJQsKA34vcWzjtBm1hsQ47cp9ZVW+
UjUMcucbESQz7n/MGxefdUig23j7b6vNDELwU//YHt7PFBXHLjXHW8xJMS594LWl
ZFTibZ+l34hyPwX7L5PLyOP7FQciyot80HRChHQ9oQ+9KKv/hX6Em8PIkQl1wqy4
7bXbN/xyiV1B8to5CsstIy2s7VXB3o7E2EOfmcznUowS/+2m/A1Cfs+k5LCMjBNV
i8yDRIpSq9HOq4U8mohw+QkYd6ZX+OWD/GerAH4Tccn+o3zWw6LHOu/6kGjKHae8
0GhKI6IQPbhL9YZ/eYFHVq3eaOa2qZ19Cc/z4KdSYRvv4GrmiMc2LYdn6DoDzNwo
Q1nGE3qnd3I+yW7eUpVgVVl7Q8igd2s8mJtPzSpol0wJf7E1GtiXodcM82Kpxxdc
m/La+x/msG9KX6a1VZzdNejYt7/8KZ8l/Sg0lIMh92slFnbf2yG2DNs1A52icHkz
+TpjisUCHlvBxL8gGN9aMJZhPyFywNRgIu1b6a0Wzye0SueZN+loGE/x7dcD6ECa
j8ts1p46dMh5HVbofJeakWqprJZrJ3IynsM8SbP3W3wk00P3dZxFatdF9v5WfYUY
rl64CNWWZ7jh/T2t3nnxplwwFDkE9c89AcysOcwIWEWhOMn5gbf6jTGVLUUxcVaE
z/F1P8qslr5jNmksQxvUGm1f8WXNIPgrcDg40lqYvRazRGUaTGDgihuadHzflgK6
aclNN9dDnKvgmHSJhorH+Q+PF6VuJ3JL4CF2m1Q5MG1Z3hBn3RxBg++3XFt11DcB
CJVYAO3lVjkX5fJ6kT/ryUktsKl8aguIg2m30lJVqCxbIiVNyXUnJpZILOdufsWT
M311KxOrJxtdOUgtH8C7XH4fq3opO1XDeJRfA4ele09NVg1CwoSxs/qDsBGD74MQ
sSgdXNsxMSQRQvD09d1BT9KPpjbKwnrFOc6g4u10P6Ycg9MFIhbP4MDZ+ukGJZ4c
6hHa61/gD6MJoHFM8+ZNw/kqjhVIIaJiv2VpwzPUkUUEXijxlmf0/8raFYdzCNaq
ogqo47UJd+iDUmH9IKKlzSZexiqpFClY+GVtj3nL7zpoMU10S0o2qkeZUjiSLm2D
9DzMjAYANWeyRxl2zRuzDnDwo3eSyXl5OTemXp74EvSa8rF4ucrORrVz/P6Ag9wR
GJXddxZNc3YfySq6ikhmnWfzIqzMYwsBWgauPeeXkjEwVWwTUiwLbwzgHmyJWyQ1
zi5Q1IOCFvXMVESxk8ezKRf8phyGomNobtnsV1nqoSEFEG+zS9bSa1+2ZUFqnhej
uQmo5wtxsNREIaeavlmK04bb1vrpxPB2yolCUbgmYPq+J5EfH1CvztIGC7OMivJ5
2xVHh1zSkzcHVPVi56DrEvXEXO8y8nGayfdl/BeDzlTMqbdcoEnGvGAuT+0eg84o
ZTWVTVsY9OOEtfkhUPmK7Dyzq3qCWq37tpZRufCvh+09LbIAxqFdtDNjz1LZNwYU
em5rLoUuLdQTnsnTYZ8H+yozm3JC5xns2VsrNtZbgqpUMKKtTZFqK4jDGzmrYlgV
TtJnTVc9Jt9PKf+PchzSGvjHhMv6QBVRgIFgTx9i1JxxKznMakYSfQVKxbErkc5F
HB2+hxeI9hiDdfxHCcFEcy5x6KkLvFY3wh/MdNJb4vn0N5cNy2EWPxUWEZeLQMju
pap9CX9PGymb80+mdCCTQq/PJIJ5ex5DsBCJTo3WNK8kxwz6nZWNlSjLxJkuTZ5M
2paVBRgYlFSf38qBRIc3xcw7UAtW5sp5KBkwsXKqfAhO9p8lTsIrzYyH49zQrp3O
T/yL7tFP65Bc0jQueAUFwSv0DbyLerUOpdSk7uX95LnbxaYIwZhfF+9dWFdNBqe4
uY+Rq+62VI0++n+6t9e2ZdoqbJqbBPJYyY0PLyD0Nz/LqDZ5jA4KAstyaxowTMbu
eEzoBXrV3nlL6QNKBvrvtaa87gBYAPg771EOQj9hg+rhe9gq3lSpX+NJcW0Nd06s
VRBxmtEUCiQlzktxkO77dFQEmwepECuDs69nuk5NFOrivJTvTvgdAutse87mrjZn
QGclLsxE/9rBNw7djs+Xk0PqgOymB5/7+E+uxPH7/0yDcEBaWd4iDgyuXuRda5PE
1lOqTou/SlnvCqeFjJS/gaT+SMS0cdmtvu3l52gMESDG3ybaQCB2drHDo4yJ4zWX
N5ofD0C8p1R2dgIetRIOGyn45KHff0A7HY217uRHbvHIaoalL9YgkosH/6XaisIg
qatn9DgOFa3Ov4purhlCUEgp23Yuo69UPMhDbGI90ZHzXhpkil+H7rP6yjXTIlhj
2BzxjVd1FpDuh3VSPX8RZ4ZQW4seh3Iwag3SN2qJwBpQsxPfnEd6mv2GThmNXNTr
5L5jlC8e72Exd4YfUTmpHcmeuBbLM8IiElI3JAt228eVWHYpl+QJuyya0dPaYZ5c
NOeHV86/AGwpwdebXee5s4QlyfyYqc4yqxuEqA52fMeVA9EwIE1xb71OgU7kbCqy
rME1Fe4toBfH1SdwauGeIWUHOocGx4PGxESE2ZXNBLJv+514UC4Pg/DLzP4Nz9TG
SX/gA9ylbeQyCypuJhIdhcQxgcqm9LodFR7/xJImJplIAMQ1WeccgjPHIQooTAd0
xXkIlc2YIDpyQUJzA1b0ImthnBlv8mlrURcvtU2I8y6Te55uWBWmXoVYg+FJ5Y6r
/O3B5faRM4XqAHh79iVV71kHHbDqLPW52GNTBpe7QTq3684jLlSN2JTPdU91PHUP
Eamx+Oa/375RAj42A0Ec/hlbgH/oa1IwADYiZvt4ZqC8imY/NuPC7fLo+qQtCJuL
JVAORkgVmff5i3auKYegJG5YELX5OuCUgZLV+A/Rex5E+Br8FlLWTuhrxiPpwjFD
tRZAzaAxuQT5fK3OBSAbZaN/yVo1W5XOO5QtdZE6UPK3DjI5jDvHDwB6UEgZyYW9
GHcMd1hnkPgf2pmzWeMSG2VRr10MYbsLs1Cio8hZuMtz/0ddVVqMiOnuEdXeVG3H
7XT9+kzK/F2lXm1D2V7Erh2UM4DGcI9/VEJTCwDVzCoxeyW+TqcDUMdcQ5s/Mzns
8bkMVd7EvuqO9DeN5QgQRJin9+hKHva4PQ8zr+fyI1gybkj8dPzgO/DgFJSvvELi
gFeD25ZOcEIhxcn8H+TR7vUo0E3WYMSXYZU5Q1tl9XNzP2tIJueH94BVrL8nG066
6vZPCDwCm1h35riBqw+z04x229H8YYkKbK11/n0x1AbEO6pnAUgx9ubR9USvMCZ9
3VVtzan/tuo8l5/GAw2svfbMS4kgsY2FJ5ZfABumKhQ1ET385APpIrMU/OF6o67W
RnBlsCV5QaCy2KrcLtn/4jgw1LsKXD4aHyCD7xsRTXjlzJ4kzfJSQ0OCYif4+D0q
L5aD6ScFrZ2e4niA1ffL5Zquot/ysJzVNQHNwLhEZC39uvZ82s2GP4GyJvLeB73o
JWqQuiv6j1QGELBoY7p0/oMD0GIbR4MMkhBKHku3p9eUMYlicmcegbBAkZpLTwRg
OE7WZD66H1ZzWVLrJzYG6p3s4y4Q+xSZS1I9Xe5/QMTuyy12uJnKriLnBvLxrFPS
UXGz5Aek70nG3UkI13DUmXbFjOfrSRkajIyPJjxslIRqgJK6Rcu347V+Un0O4Qv4
tiRW7QhGKINyrStRlq4HkY3N2+YjzvAqU7WltfcyZq7VxBsdXeUnMiZyUaZgYvNL
/SgiYLucuXK+Lt2OiCyo8wXc3wEaWDG4Zw0nXbxVAJKda+Ob1g3rczBv3a5lyo0F
8iXaOXH+l2MpW1qZIgF6BO25ej54Nq9fFSwlJcDYh2l4SxuX6cTto9CkqcoxUNzN
wFh2aMl3cx2rbDdGuD+l4aPFBdMT5NeET8TNz10G6RFYj44LUDaEd49E718NONoT
wbif4HimY6QorzNPZN8y+c+UJBM66wrDbb9mZN6Im6tGDiY/KCpvVNVVrl+AfPPT
gohNt7BRQjWZ433fKAWckDKAKuok9xDhw8YQlz73fsjlejvReCLbOpG5ty93gtB+
vg1z+6SDE/refATnullIBGFhYZi2jlhER8Sdx5mJYmmrfyvWZoI537tB8NTP058v
5A0gKPp5ETMqKMdtrEl/6AAP02chiLG07smwdJISPkO7+3jqF3e9ENXfdiMlEu6e
9qpRUjk1kPOB64YK+HhjcP5PT4NRfpL2ER1zb9SVAwobKEljWM75JSNkKQ/WkoPw
YEodhqGL7s4xQg/iHe+TZYvIeEtiBvmnw83M8AGsbze0Vy35yu3ium0+wb3vvO7r
+27uEx1BWOQXweUy9ppTws1EWmE0c2fGqtRbc8cB8rZDnp6ccTbsgNb47eVwgtIl
th/Aln1QloozQrQrIj4n7ZdO4PLd0mhApSsgGTrWSwqt93zLmQ4GrPaw+QRybCmz
MRUMydQCwGPrvr3o/nxet6zM+ART2fFUAz6dRkXvg6qoWklS/NSSBOMeeWNzC0bt
4lsnS2NHDaEh47hi3qOmA/FC3b4MkPTiK8MmPvbr+ynEgErhPkX27vdb4wChN9aw
LWc++vzRLSubFhHXyu2MEL9KO7VCz8CBWXdLVYjSXx+3PXWNl37cK2JONOMxvkGF
lHvhxnvuLuUB6ui58IU1YMNUH3Z0ItVBwFk/9V+yTY5U+Kx1Zt7wYpMTuE9WeNzf
z3jx+gma5DMZKzzcsq3C2bn+bHGWqNcwvPE76YNEkSgxse3Nark0JRa9+JurngsV
6RblkBUMvw9InDHvMK9cLI1QSMSFLKNmxQzrCg59murE/dU+Ap1hrIfPqjzNJg9g
xgI4FP1dM9GgdAD83B7wbbbl6DQu1649V6Hp/uD8PNZDnwOhtR3vHppyTVROD+Gd
K5RrNtKAcwVBJdo8tlOhajxGFqNhI4sD5UZWT+Fh/H17sxpV7NXjRqnOZhb3wLKH
hwI/dVwLYVeHXIcQbEci1RRdEEmW5GY9/+u4j3lm5RUoqCyOLuursgaBiKAu2b0r
Q3UA7J49ZN82UIJpqqn3rf3OmxKa8MAclTk+EEhF0Q3eQhXvljDRVrqGng3Wj6p4
TdIJM4LmyofJvMUGI5OEpYwTL9gwR85bc6hGCcTfrNfqngCtCuNFGUp0DdcEH3pp
9JLerLYexrxXAO70WIdhMCxPRoBwFkfzwg25u7FThbDTNAzcrm4+5+Gb4w4t9/m2
6L22o5vqvlomvCqoIkczH4Omh+COvqMp2NB40Yu0BfHNvOd+AS1zQWIWd3cdlYeD
O/3njudOELmv1E+hQsZu2boBqcDaBe6BDJzONLWt+CzFSUxjSY2RO/SvqduuVHnm
V0XcYmgTrtJysxwWgfz+9fEzap7+AWOErHsMcE5wTUk4Zsh0NVAU5C3SU+llxRw7
m4+GRz3KOyMwi263GgqbIVtpn7Iw6sXrzSrHldo6KO0zjkY480bNDVTyHZDPMPzn
Ieoo2qZ7uRRynp4m8juvkrbHn+V6XSS5XTe2+3FOCTj+FEokuh89FXrpG6ujRUeX
IMHKYx31G9SrEaAxBeV+4ioCoP+HGIaKT8bAPIk+spHWdKsdNSxPMNSKMaxoO8I/
fdCK4iZEniNhSWILZEsGkx0WWvHFQHPTi9O+/wgP7qoda/Yc/ZBVaA6sN7juI7Sg
SSrY1CGVF3LFLXq7Lp8EToofoHDda835BHQdm8k5pS8NuDTXzTGTUkIlVBJtF172
+EA23Mxhpa+OdqVlLeyGI9gonxYJSgUia6cqRKcKOQKMWUeAxMVLH+oz38dODLkM
9z3pIZ/91Lzhhv3b7X20d/7sdFh5yNP5cPtHGAJ22y9GILcgw0kIvDjrGsGMZg1/
BXpN7EbxLMci1v5ZuTVIo+Q/N78zIsnVaFtQJKQ1ie7/rZIKvNjmNHFeObO+3VA8
rMe5HkxcFHo2bO9Xv9BrV2STtZxZqfgjlewl7qk/pVwh8h8wagYt7W2SNuljSU0O
cfNo5l88rpnrDMrukwC3P5H13crEcemVEzxCzWuHeEVJ7j3+si7QKYHvoAh/wYb8
lVL7He+SAK6jH/mpNwOer8ZafvfYxlwgqNdXvcdWRKRW/so/z44lsEEIGwvsfh2q
b5XdG+E/lCvyP05UphvS+sU7qPNNrnnwzdhSbk1IgCr5fc3XwE1iLES+eHWEOJ5c
rM+bmAEBUh7dHeqaeySh4uOvNgCyUhZKpd7Mffuz4nfGY/ne0XmPc0lnGNu3rUgZ
o8aTlIJ5H453N03gOQCVo6BrypdayWwcya8xmXFiFVoaF6fwxxsW46hnlOebp1Hq
m144I5I7Ke8FGAV+73P/Gd3r5rAdgStcrxVCbmEnfxkCgx8MX75RyDL2v4kKIr1m
oFcZjevhdGn+IwxI31Ul0W/q5jeChFKIZ6fOg9z6eJFPx0gjtiPhwwzKUHhAxvxn
8bXxE4fMotyOS8EqxMkbED/K4iHtekW1mwieFhk4WQ9G+JcczDsLRS4YVR8VBS82
VbrSEeBYooaNorQFIwRNGUc96LKP2/hZNlw76DbQbTWRzZdHCErNUZf2znM0HzYM
OnKJwqqEoS0WSSPQ0k3AzZG/3QdQXPmnhoglta9P6EWLOfFOv7ifdZRmQ1yG4k9E
9UhHwVKtqJ6EOkNBaE5zgFVuYFP5hFmqF5KbiGBaBsHPQL/zZHbd9MTf+qxWlcAY
MtRSaLyT3oc2SgGm87RxlGjf0CPXJMPdtRFWqXD4zcCHY+hTnbn1dhveaSrlIbxr
vzvJTfuBEtiB5/dt4hILAHc02ZA/0XcUwFaS92N2CXlgCLUH5W+/XrZhHSAyMi8M
2I0feAR/JcoAj4B6s4erhjbDDfBFed+/HyAObGIKANIvhanoibV394z9NARjjkVG
FqJW09KwggR4FraIiSewCGoydL/AlWaZnRcdAgFU1/CF2GR33/wz2c6VZO7xhpWZ
0IbTU6EeEHnINTEXOxXIV5Q8yrdD/+B1m2PIq6w3Kkn9nq8tB7+J+mLGxMmcPnvk
KrGzchagX2VQy9TY8m1uGeGBc8n87cMIrYCi3sEIaAqXzSLlg5Y+3LlsVL+u1DxE
suAPu5351jSR1DI1XAVPNzABIBuFbbIJn26N3AY/lCS/BivhqGD3irUHzxaUeH6z
svNCPtbi9jXeLiu9IJGLhhp9u5f6jkzDJqGjJWO1wLGHzJeFjukQX129MkESXVno
dz79cQ2qRnyRlvEUmAlrP9mws4lh024rrhLwbRmc5lC6UmZp+riAg1x4KReznU+G
yBpnlbDocMNjbO0zj7PnV6wbAD0b3Hmk8MRqREYZnFSXx6332tBspQLjWOx8VNmz
TPxZmneVpVzQV9udxvss7n2THFV6iKel37TK15yLIM+VptoLvKQta2seefInNIJg
w5n+U1XBdAVb0D9And+b6hSlxqAseCHOk8jlgQ6P4N5dVAw3d6rKwOOY+V5hlgiw
TWG524YG3LQqvVCqo/S+7ZQRNjQhTdnOSTy8TfT9WHUk3OJqK9wWyhoD3pi3GXI5
nPqLSjjH5kyQglOwd98mIflpfOEvnBTfGm9SNs/bphZw3+cy8n7ahB6oRouvTR2v
hs0PjRolFoiQujoBpaoaOFrIcmnKGBVUnf/E8vsfIOcPqVBOUfJJ1Y+D3XkqKkDl
SnSnJ+fOwsG6h+s6zBRbX2OTuQGKrQEiXERgrxwVBGfIhAx+DSeQM9X9c1IEqird
5ml8C/vjuWbdrZuLxDMhdYmz4q+RZ2altHeZ4xZzARyAZZ4Z6VJ2Nx0EQJcj6PTQ
fnpYnvGVcMJ1GFxbG1DFzFbaxQ2eiSjsHpJYWcKYu7C273Ayw7pHYF3B40RFNGEZ
hTNJSyioRHUUysdDiUZS4CzYu2EaEl7XofKwUpeNCPxVSsNyLdyY1WlhmfsEjNqi
saW0yfvo6fq3GDCItIIGxXgJ+LJzH+nByp4rmbZvnTgkOHqUEG/gIjMitRDkRrEM
N1WsDUBDs4V0fcNzJdz0dA/GitjU0WM0NdLEP7dUMdJVUCl40RWuZEm9YQBGmzip
BoVURi2nLJgu3DJR0RjvefVWS7Fc5urDMWYXo/vDCiUxg3ZflOelLdHrfECRXNBN
IqIqwESoMLucAlnJ4Jk+stAQK5b2VrXje4JElkhgkgyvJIabdQ75Ncs/TlSlZmEc
MHzvxQMMWC1/CLiDvWmhEax2fRNcxTYMGefGyGXQ8khxKfaLFMObjovH9zwqMn6o
klnMCRD3+CVAfjuELcR0Bznw2cqQtw4JvTzX30ArBL6wphZRTnAgwtwGIX0d5E6u
q7s8sbw7Y1AO/ubml1jbiYQarBN1iTYJDtNZUQLxwZDlnmvhHTtpi6lvrKEyh93Z
Tr8YTIbbwowP0Lxvi0Xo4bZHS0GNUxQtJd0KvSL6wobSIewrSMqUxXx4Em1uoE4l
kFVcDoWuanC51U4H1w9QpChHyxID/pBIwiIZ9O2Usb0bU7zbum2doz81Wtk5uI5V
650UTs3hkal1IOe3DPfYMcbErh2zo8gs+bEHUVpcwhhhyZsb+OqTmMc7sZ792dr1
DmlUB6C5ObTkC0CH7Bfvs3cR8lR2KkaOt+ZmWprlgoRrjyC2fjWzqnJj8bjb6JBF
YveEVC7BQshWzOREnKF/HQhXcYV0PFjR4UXJgg804vnQyp/IujACuutU270IipCW
kCcNmoktiEUjGbifOiRI5AcE6yNlQeyQPs8chKlSlJvHxEZlLsY3X/7mW3IsmD7n
VfjTWG7fvn5NQZmdVgCtVRk5eckkYeC3VJE3oelqOW2yfvZc+8aK+p8YaSP6qhbw
T++Utl19NF1g8R5K4pfYDkXnyC6jSeNS6DqCabP+1i5wy28V8dCF+hYgOcvwcQlP
xznE2P2LKvWSaKBVS/ddJUgfyddbUJhKlQ9Qkxd6eIKhWjPTKD6she+AYOhsA3y2
dz7vgcIEMAX8VGTdQ6zzQSrastVKtdyPniJS6GCyrHMkjM+wOvYj5d2Mzg+6kjTw
yscfrMgf14czY674e0EhPEF+18jZxxpCJ6vutPwI1MQYhxfpzNQpfAK7fsuI5awi
g5/1MckxcjVkLR6fqsZUjV8nv8z0+7EcvFPRJsPjoRC7DuAhiMkvjWnm8rC9ybK+
98ZcPJXws2a6WLM7UOyDj0Y1DmOod9GQbtAaA3fIhRBusrBAvRa2AXvzEHfaJhdm
FxlWMI4puN13xnFZpC+SRXbOoCRN3bEnmFPqBAYbB7Xkp8Tf9hRcPHWU3y0o+koQ
PfMV42vYYRRCTUTehfECflbHTs48SqcoJ/qMlESYflFN4woFlKBO/hheBBZzNMHI
MDVqZYyBrPlMyozxUimqYF6p+b7URkcjCnqgcv7Q5oLiJf7RkWlQcO8WVntcqWS5
VyA4AfT9ucGACRIhGAEA66QsMblUexwMe62PWGK5Hwtp0V9hKLKklFeQl/icyzG2
8yxhNXaeC9y8Uhen4O+3daV3l2FYMpV3Wa6qfHICCCxupzmdOH8qXSaCoyhYkVJp
/IdCnVO8bRHhRNGXnSU7MuARsZwID+I6N6iXt3GDW1qHuuyvA0E3JOeM9CQ9s/sz
qAJhY2H/QAVkYsRC2unXzcbXjN/gdztZ4W9Nw6IpZgDIpIEr9lbRJCzEyQfv41s+
jVlxlPP0dRH6eYPm+XMjDT/dRULoiWRLwMWC/qnFaCyKatqUvjlkEe+fjORebf4T
xvVWqcISo1pwB1HSTcMWmUddQYVDbSiCpAphcoyfrFX5d1cZrmguz4Yp9nArFM/H
xu9nAM0cs1bKMpajvlkjh7AggMzGf+ISyQHvuWGRJlIkIsXnmr1zenHyLVcfwvGA
0+5UAtY6g71brAAdmwEqNxIfNkIb0oC1tehVlKClwqxe5C4MY1NZGOTFnZ1wnRuB
FsE5AjcYeTrbFnnCNfB7g8Z+0bNYBnqb5oi6f2aYn+X0X0me/C2KCBj2Y+qjYgx2
na2Mq4tAIr7vUU1BMTdJsW4mqYY0avb8X5Zb84Fv29FOxDdynld19jT5RxdgKjdL
QnRcGl7Y9N1mTBcET/IIMOTBGsJ2EX/ZJ915vdQWk3jZqkGc3Ad5yxd5mtBF/gVx
5oqUQADXs00QL5hCHyfuenH5PyuzYmO+LT2CB+IDWuA1ZvfLs6GFrWNaAvVcRcpd
zQSXA13P/oZ8oAbDGhn+h9pMYSm20uFord8AvTeDW82yhbXP2rg1F7Ophb9gxv1U
Y2WYVBYDMIV4dbpA9981GGKlv/H52uFRH6qb51Ba4tKJLIvhJnmE4zHeuLAkM4MF
vp4TpDWno/2hIN8EXnkbX5DLpOD+2HfAFBQ4Vz6qKClX45n1CawE1p3J72cVXkwO
7ouG6KrN9mtbaE/pamKRdadI6MiznG0xGHnhUatzqeJYO0cPHMt21T4J5/LqCfm1
6m7EBaiOglan3XYI6vTbxSPMpHdaRMO3HG/ORdRU4AOo0DdxdRgfX/QL28LETdB9
vR9SQhasMzyxjKbOu5DQwQprnyfB1ulNLeNfjAnNBMur+etUw64+HC2xjB1zK09p
1CPKiVUc0gjNk6JgbT2jsNVNzJg5gIG9MLmIPzvgYuA+Og6RYKHL3+cAPGVXw7dT
ad5wyO2zPi06gKbr9R+SZrA+sIQAsUkaj/VavskfYZMsqn4oQGdpgIp1TJuOOqyy
L1lSvl7pOMhCwCnFEas0zjYtjMRcNZKUhXWo1oWiq01B9jidWeKKNY63jo8Xfcgu
qTgE6qQwHBlW646E4UTLQKdL7+DHemaRi8BIPq6VtgJea+DVAzhEDk0XwPTFYME2
ZtLcTJbYYT7P2vO6BczkJmIc8dIDZD+iwY2Pkj2vQ/TZUNbDmxX/o+m6HyoK+ofr
qhW/YIqvVluBWLbs+f8w3oct5kGVuds0eAPhAknk2eikYc+TI4kqg2qhaIWVZMS+
CuGxWX2IYtPQOCUJBGEjPBiYuc6Gy1y+44pjnFdgAYXJ0okx8n1y0NYbTRjiPSRK
6QfFQbQiN5GsMU7xz0bQQGR6zlkGMCt0nfdLn5h3I7H+oh6zdluR3Jmg0uSSyR6P
HWUxcDDocKm+1pBH5Hx4QHo8mYnxMmttdth1M9WcIiTuCxnGOgZeghQlXIKjruPO
ZCKTUuUisKWG0WJemqZIuJdBkNwI4WnV4WKqJMYNz4Z+APQBuxphCm4hxRjy3hY8
iq3doM2jR6eZQkEc9J/HrmYkqCUGTpxwSk77FKNzgSSpdf5hQO1ki+Zepghsh5st
ebPWclGwVI+T+EKDRq8lDpVhC+gqnLvKhTqO8sjzEqeL9xyRCXEozvBIRkkLPHUK
kifg/63h/GCL3OEQRUfBwJuyyZOwqJ1VuUC6PjwMPHSmpgPwvngjtVc8wzGGNzhc
hEQWn2XBJ/66MiS+M/ddqez65Wt0XpwFCAYYZslUAjWOWSABcmvVEtiiVvy4Te1q
FQJT20Zl7dEF/IsBFS4rVXu1GWYMqoiw0uU425kJ9Yan4Zd24Bc+8guuutUGdBqO
vV5qq9CbnK0AgEtt6XIzdDglHjgYXgObVDl+8fVUW6CMx8jRvgaj7NdNxu4uZN20
FnTl+xhhVNsn4BuVHD0j8kwAwSuBuEmDQOrv4ZDKAt2Z5aCRKHYrO7URBkr++ttc
BndSK0+drG3kW1HTUw9+b2PaAkLd5fzyt1g1KPJgW5PBHIOK8W71qLWGJGFkFPrL
7mpqcJF1AhbpdvAXAGMJveY+mbnHWycWPlCA9pFgm0K99xbIEpimiB24iWHSJRjf
bAfTqRmu5uaZ9fOgw3nmxk7+1PPwiw9bM3xAaYTHkUQ0MXcViXVpn7VDJfBVcvth
CDJ3XD3W+sJpchb6A3H9hohheLsT796nj/tCwXqrSFGeQnpVQtpT9Y6B6K4kPoPr
H6MADkAxmhWTm+ziYQgbeMdfxy0Br2gACCnjZeidB67cjXP3ZlyS0NctTbJWJBz4
JJBZ/eqLwB4Q52GJanvbhw/g2jDvvPi45PuuYFD7bDcgenBsTnykobHgde2ciIRf
8AHxBOaSZAMpdHBrNrv+qG2tJeq5YAoMTcRlHmUUh5zLDSH/Cs7vNbAH7W0SzHZS
X8g75nOllpj7xNA+jNrwEiETyX0NtaQ/7IbirYvKukkqe8zztRJAJt9app1cqRrj
Hkyp58Q6+0eYirlYvFsIPzGKDOeM9satSCqXvORtCpW7X4QJGyaSODuJNW/1pr0j
PKLSFfCj7jnCbGuVkiv5goAzoMxc6i2MFsXwkCZ9cOsVHFNKoqf0ku5ijyCs8lld
T/d0G6vBpfv/KZmcnxPbPfpKB45IJDfQSAWDUn7qo3d/VNZdDVDiDqYdZxZgYJCw
IickhG9mnPfkt2zrbxedzf6xuJmLGAD4SPiuB+ZBjQD+SdMPf0r7ByvBFkq+1m8+
XxEGfxTvPXI3+vaBSikVNRxw11PndmqZl5aVZFdurUmvViLzj7zez0HKeqfjxuWV
eJ/Y1UWOijvJnclz32DSSDWUcwZILUOe+62EuKlSH0sUaFNY4bINs/u0LzS6RmvM
PBhFdBeWNI9ZAKEMcLQf2tyLwbCPFAu2UmaMggplEQcbV0LqgWcEEdSycE/HFYMA
wzoG1TZ9YtH8neNxOlxtJ6RZ+zHCHysg/rhu/dtsXS23scWTBNrxlp4zw7H7diY7
dr4frrmAM//Mktu6qeVOg7CdcOU9KHep0hbpqKiK8oG70lBH5j/vEmBg7Cc5lHd+
tdWFdWEUjq90CmOpURAAZkW9Nhzl7S6vKUs7FTEdpSqb0XJItGD3qwWSf0ddMWpO
DAaZDAgENTPs3S4oKvS3toWoGBHicLCczaLr4R0k4/SOUWiTEKef9QuSm9oXhHCg
mQst3PlO2p8ZEQFVM9upwBxVSblParRJFKm6GkYbaSfYHGV9nz7WQUI09Og16JjZ
VMGnwFpqn3yYclIJUA8ltCvEJ8Y0v+F9SiaBE3vMtl33OX6eUjikRDsVlWJeeh08
+r0QJ3+j6g8QXGcLxAYUIQ7VlaWyzizh7FP52BdJvjSg+ixjqBpIl9PMQiHy3ZmP
j33hWIUSwTdz90N/DAUB0ePg2uPhMaxkfvvp2/bY6kBVuIuQW0sa34C4v+Ht3C44
Aii/VpZ4DrocBCW9lwTbvJI79aSGY4pOE2/XowCgh2pDU06FLTLj8B4vasSDwjzS
m0oEskNEz5jrd74+Ke1ezl2iFnFhhROCnpKJEtGZlE14dxT+vnEhHgPKCRGZWD+s
AWC0gcPadf1Z2V9jEmzfu6NU7geRLX5EOYumlyuCcyEvxYOtdMMqaDOOnlExvFLT
p+YUipLx4wr7YyKRWxtEoDDzo+QzMAeCqpAkY3LtBhaOp64SWdePMv8ui2TaEvvw
mJAU3iSliDndGMpPjJOyp1rNT0oA1Psry3uPDnck0FmHwUA287fhXEg9JV6U9srB
2MKUEjB+Q5Q/juTNotGN7GBAfD3rcci1oA2nn2gbEZTDTQFIT8kToCuVeqFtdFqm
QwWzJ/21ieaiIJ48Nj/+5dgII+6EqMmeIJs8PFa4hS4f70RsiEBbUhPEjtI+0nTl
7Yrr2oTOoHQDHzUT4msXB1qO93b0RGZnsmmN9GJ6U89g4DVPQIfCWexwmv1OXrfG
MMGlfszXQ4BKd8WOyHiPWjfHhIDR0VUVhIHXwNpxEtxvBKEzoiHhkG/SSzNeajb/
SFQpGvsEZUMiqj/9oVa50gM48/eHfUEZ4G3wYegvlt4HnY6X9AgXYTr7kBH/mOx4
wFo2uR8bJRcRZtidiOHtksBFtLs1S9Qe98QDQfVojR7ebk9j2gfAx0SoHoMA2ThI
HQenT12lJ+LpoF3pw2Mp+lQZWzsNCQScqU97d7dOHkHMbyxF6phpYWXHR2i/owPi
eHlP1kBzYQ9V/jPV7Pd1WlEGmO6CDs5Wm17Ssd7nhtKfOJg0XpuyshG1ZxLuRP7t
TmtytnnrbapPxLf2s3vBXSePFaFONkUBX/Je9y5me0HPEMwiwEaDdTyPxm0gzGBr
X1EpB9UDE6CZv9In3SgMnrnvV81DMbrNjl3+x15z2xlimihmrLCvjxe21wE9zjUc
Ab3dwpwraZlFW1rvUBTEpDcmAJi15ttmvQxqRAJUFm6FRNzzetoxn7BoOTlvABKj
+4Pqd/3u5/KZ9EK7TnGfZwpBr1cq8XGYr/ORgOS9aC65y77kxXMndvW2gLpp6VH4
TiSQte/wQpuu32Te7nTrBa/1ca0KKkkP/cc/DlPrQBj3n/cwPiR7ok6EdzOHE363
rRHwaZaYDZlnO7Z08JQNy4o4dgrHpSA96lfYN2ot/jEG+uPP1pUK7MrKFBzY8Zwu
AQdolPCXoDVcuqsmrmZh2JySqC8ssD7haZqL6NMA4GgAA0N5KI2/kKCGAs7Ojqpy
wQ5mPELUOazqdYG3Tt5a2iHZJmsDW+9gNajdmqnAMLBo0ihQqM8YIr1brDefZE97
lCuxfSp0bxGrt6X2gaToD1PwJGo5hfs3Z34yYHJWRfG80nfLWUhrZ4ITZ1jVEd1H
MU/1GbkwJqPrCLIFq8/DJLkuZ8s7Y2xtOfgnZPujzeV2Ii+cuRh2JLqz+c9c9LwR
Dk27KGJW2QMpIisVfcYHtaQBaBKVXiz/fcPbt2YlbR2rzuPWYdAiNW3E1Z8oAcTj
J2PllsSkZiKHChQuPUTVmWdTHEQ6KSmH9JfiWiBms/BaG1iIc7zAmtRC7AVsb3Kz
HR7Gn1KXNC9H57k+8q9JRihcYzwKFVxLM/zfDrqKFGn0h9rXKHy/xPPOCnVRhgWW
WRNPT7OvdXGp+62k4u19geO7DBQzONcAyPbg7VIfXUG65d9YMD/qaGrQlqiLshHl
0QTq6CDQAnHQopoPGfKpThknxTzkg6JEovYrQlrtNamh8ox1skiChX3wIIdRgbgl
oSs1PGiAhBFCLI+ygpjK1capKA027hl3xZ2d7NFxa23oVJOeIpZmtb0scexCfL2S
KNDCdRj29AWRVcprncYktQGbqUiRexDiiyOc3SFOtdwVIErAuU9kHzmrAwvbNPZ+
Alhp9qUL5j0W/vFjH4ZX5aE7HQrCePtxHqUUIYRgEdH5WzTxb8RG6WvkLeO63daw
fN/EaZ0kg7Ezhcrm3AEUov6CnB9GtCAl4bwZQB51R2uyP+iizrrVLnByic+RLi4S
Dk2en7eWThF9Um5WZK4CPK6Sfi9KzX1g2UHw+DPnqcGSUizmJoIm20L5wXbxNod2
VgYElAhUb4CaB6yBAnGjCoNgdq/KRbDXCYhuH+m/sgFV/GKWSTmDG2Jfi4uFcQtm
iNp1408qPavLO/R52Yv26r6+qUUUcQpBoyxEuor6DQf7dtCf6EvJ0R2cSJYa8KFO
8m3ezrOPVkubWBwQ+V1BIl4mObULgtHJpcPHBnsA6GxXRJFFsb/sfLKYQdKyGcZT
i480EAIUcElGWqOJ/0lfuQa/JTfhHxwNFvvcrdhhF6pzN+2YFW0wl91eYMUkh/0z
yMnVHCahpC0KOFfUZQGbne/m28Oe+hnsKyugGlF83SQz0O3poJNRcldr1X5tsEBy
oTf3ghW4iT7WTWRT9JBGLTXmxZeTZk66Zu3efyi7PtVHnS2dU14HZWyHwI9pxcpP
1DpGPF23Qqec2cvEDvhrl8iC+k5Q/5+o9sqFF76yKkAzwpZogGbz//gmHBOqlSom
7bpP2WYdYwkTfmj3XNnmNxSowo0y0zChd2iROubQoZ7MZ0xhDj9CIAa5weZ/748K
94x8t5C5SD+ovSKyuyx7i9uhnb5oAn+zOlX08GDI7MWUVJeEk0wc9c3N8lTTUgkV
aHcMoNm7/A6h2zB4216FF9/VevZEVDk91Ml0cFPZzxsHTJMnvq943oasXs0QyxLR
kMrCRrGOEmvfmtVks4ur6c2xCXH1v7ckTKv2BsLluUCs5W1+5VuCEZnbKPes2an4
VTeZx5Yp0MARfF2MM6q672QmtnJKRL31kkPtwkJ3MQeBSn4eyGVQO7aumGNDne7b
NUOX/Cc284HIxWsbqimYB+oHfRw4bZdal7/AIFqC8bHzqXCW1db8lTEjP2cod98j
6gKdw2kmVUzwvfCsz3qVCzg2eAF5hvTlWgEgeum7pMwEPyf6ZJKdpQewaqnbFhPh
sfiZvpx2VZWbzvlAFS+3pA2pr6ol6zvKmLFV8Ny2eZv6mEchXYIZx/4jfjtyv3l8
UhQb5YLwvc0tjZ0PBy3A2Y1hQX83C+XWENSD82bvv7y35Up8Kr7uL7RpJEc1JqmG
yfOmza0mjEhKPcPrOQ1iPXUTs6G+okgwP8k+KiEQi2faw0Z6iqoJ627opx/yUJs+
7Bm37RSAoGG/X/q/2nRCjBHq4eTQSwB4dYn832Wlmswe0JrOai/9Mxz6JJ0DssgP
iygwTwoQYfUL8zjyGsj6kOL/n4zR9dnXhlz07GJihOPpIx6JqxnnMddIALtOJNJ7
/hqeAaftjlRV0UYmCo3eDhrei9XQN7d4xYDyvSDGfjtwn3BVqjBXHd7zFTUDHcPq
ZjVbrxtbifQ1NOYXTIfBqzybau+KmYTq6NC2fSmeIw4QwJQnTTeelUx/zBFTmK62
Qw2pKAaIUJvtm6nNbiIPSudWbIVnjgpLaYaZEry3pkeeJuQ9V0TiJrViCFc7vmPd
9q9swWM1IniEjSuyGRPntKEwET0DhcRmjC3ZAbRCd2AnTQaBqPEQChPs0iI6x8rQ
Bxg0xG8nsM/FW8vdEM0ir4I70KssVrXDWDmNUnazm6fFrfs4hLLozDnXqXw84syG
Rp7Br0qG6MbAb15o+qUAEgnT5cWJH9EKGTewSuWUOMBFMU5rrk8AJuI/BEjJzKwj
0ayfXQRN7GlT8jICseiG+OHPFcJ93BLBiPRhCsY9fQzPxw+pAd2ahT/KlsCgWfRl
wluIxfkaA2CLQkuQWY/5J/dALqSxJNlrihTe81XvySJUKutw/dOdRvp2DoGfiCAz
VIBWB6MpTZlBgw3ys3wooxwUQzbQepdyatY18UcBHtxlA02xI0Y5K2iGszvctFaN
SUN7/QgPpHqxCY/lZa/Qh+thQAq8ylb9bJ0sbjg9tECGjEzz3LAbzbM7Od/Y+qG/
1AGGUrIGPuXRjCxjclemuAlIUXhOqHReDS1d7v7fm2zFbJFSl9GHiK1tA8NYGuqO
kXfCYFTxqloJ4Ykm02KKHvbbxpbGS9H0o4EZh0w4SoeMIwlIxLiUUQnh/sqqVUsn
HiatodPMYyakodGIWx2jXoCT0bX3GP0c2UZUsiRf9HyH/qp1Cx09U1Ui4g6it5AS
ZKsjY0kkSRMz35Dt9TAi1uMy7vh1hkkktFJAP6DEaMvt5DIMW19dqpuWfk/3jTUP
RXC9tREG5hyhz1WxChEV5ZQdLEToktPz8w8uU0LRwkWdnqe6R8pRZckRQcmPlu5T
dad8u/JQeS7d+M8wt3SMNnRC5nrfblsBSW16Yy3yC6iWdU8er5GareIAtvlYtoaF
iRCaIuUOzlTb5vxVb5kIcRr4onQYKHCAg2WsBVldj2aTpgSEpBAwOfWEDfWqONUn
PAIB2wqvvIVXyzfVDgBHXnn2x+DaDipZMZ4o3WL4FyQ/l40brJF1kulU+GxYYJt7
MQ5LxQBOedD8VpqEdl/zcDV0qriGZ41RV0k0RzUeKUz5GrHOgYQrYK85ym/F0PMu
SYl1t4ftoZzT2sU9l3brVQI2TdsY/OVi3BDRFL+//lgoQzZNI18CW4tqYNxYqqU7
9p8w2VAYdC7t02MJKvKQ6jPPQ2zvObF1KXovNSOamAyy+3jQYWoP5fpSeMZbSuxx
rqCnw1eu4PzTVsKVgfKAHwn4ZuTxm6F7C7y2DpW2H/204GQoHt4cAMxc6xjYuvM6
fAYhaqaIBmR+D0yL7m2AtCIqSZkBQSpEr+wuNjWXk770ylwL9gfvbS7Li4UJ8oJP
ydnsYe/Csrq1KuCgH4Rl6EUFdzsg7pILg5Tr5aLQE4q4H+BdgE9dJya2Ckj1m7fb
4UMCfVtqABvRoW6q2At/ohi5lhbHieQ/mTqZS58N5FrYtQwlIDjn2/JKXMReoicw
3wkss0UJCtBkmZZ1MWRR91KgW3ruO5wOVenkkAQSwjT28aNtH6OH76pSS9fEEuHI
PV5Y7T6px8j/QPpXufU3XS8xnWNsm6oZpnezuvF/WdkOL23BFogPvq40eexyiEVF
6c3NFyWuk84TN+TAtHYrThY0sT+ix6VtqDXJoHrRMoZcjHSG/e/LGu4F/ernJ1wx
m1AYqN2Pdb2TG+b4rc09KtCv10Zs8QzNXFWC5FX0rNfG5ytgu/xyo+kjybnGWDFs
PhEXNiwCetH8GZtmXBdVtO6kmiNOrc3SEDY9ulwppBRNF3DsRmbPhZhkf9+CnFvd
zGPF48+umiteMMDzyqxwyYF7sZD1i+v6Ti4RxjgxdXx+LSZMgJ15utiYwQ8lAHVQ
eCMjYrTndWaLlvA0xZPpZXCO9fPoUlCThagEcbCwDJETEY77HCIFE+srOehWqDHX
JjYpLhfhIol3rV/4R/U4rJHZ0CqjU7aM/wBUZjD/TPxUAd6pKI/ZCiLoRoXwqs+M
QAB73F6xjLhU67tA4iH8vAmHNEDfPtjeXjmiuES1R7hPV2oTYZc/+2+h/t7F+CJV
D/C0CnP1KPnsdU7VybYn3eCy58kJ/wuOdSfN01oPl/K/H74tyovColaZ2JBgvrLK
ZDbuGz395BGARRDlf2gBA4szGrVNdH+MNh0ZmPjTQDeRmA2m4Kqw8aQ22ioqOr9e
mffZ5VdGHnPF40ZBP8Dm0vIPu121iqCLrpEap/UbsYLXh+fKciAtMR5HuyjAWqWF
OacnyoJ5OvrmygiDSNN+gDA9qbc57zkgyofH+1fD7D+uAYE2GsRFACMQbVMA2J5B
gn7SA707V8CzQU/y/sl9p1NEDWV57eIsDUCmK9mm0FkJFad8b+lkjKWlLSCQFFPL
RnCYni/oODpWY0iZSEx2BqWvVX0BJnXVM5sRoN1L+loeCL186ob505RdC+jkOOmj
a3JeEio9LhDFS6ZZWQ9yUPCGAobPGV4QR0RbC+b4unRe/6itx2VaAuwC27Kt4nxg
2yRhPVd8TTzRT3VjEGRyfiq65jpn+IW/bakunPuwyTqnKXOz2sovdpMPovMNd853
HjPpNL2pSTDLRsq8GOTSOsXd0wDnPgETymWGnr5wyIpFB9xJdn9fFLJV0beZ9oqA
ryx8t19nFSdNWtzcdxON006bCJKbycLHQuCClWWsfZiN4YDxlQOGX2wJ3VjBfuqw
iRFdtPhe61Zq+cE/VMl3kcMsvRawaVpJuyWph8Qy2gTQJRBPiJu+5xztZT+Ul96o
TmIrAcYhCWc9NcHIR3jKTSp9hTf1IaFnzR+zpa6RPCGCSen0RPTuP0fyGa+quGtF
gsA5hK9mcq7Wk0syGwpWNQxHeLt1g20oLkSndrDs5lzXn7vtYquCJuJNPJchFEl1
3SjCIQRHTAJC/oyzhe7Zy8HvsWHC5NVLTVW9tvKDD8vF/uJEbznaCiWRQOIVTkkg
u6dTKFIww47k21eyFAT1HfVt+52M2LVahU++IfRhIXRv1PYwk/oEG+WBSnp2Wxn/
caXAtVDcuZ7/gE1IOckWLkoJEZM2Vg7iHQFWBjuPnNie6aoRpjbHdjqlpcvp+bCW
aztTstfkTyvBoaJqmVJNUfkqPxMvRV7TfZqJNtVGuNailBtlP4OjGp4b64Lav0hK
yOT0Me5h3/dW4K+AqSNELbvEkklbo3Duc8DUvxLIU1oMh97HRAGokyfNxItjjk88
5DKcMceBj5FZOr5nPL6EvYfjptSaV03xZ2Wk7vm6dE+POx9GokDF7m/HCk76Rh7G
y2OiH75Z2b07Fdj6gYPCa7VuWbOUjKaHvoY+4eaTU0S7PRlG+VzXpVcyvhNC5gf2
0OQdKqbhpqhEqglXagwnycJ9I6Iidsb6PPk6ed1gqT6+HBFsCHIIMDIpmKMA7Py2
3SMxZ+SXYtxhWDa8ABCcoQ39uFg4RbU+YcBavVDeUT7RGZP1d1VhIeb+SeP+6ph7
/eAaq0VO8pLEnaqcXtTWb09cvfQMP13A9uiRmDW6VDH5Hz5LYMRgNrd2ZqrVbF1I
4eCle+n+dhWNo/Jhk3jvQq2pHF7gzUyII39VxB3m520tA9up/gbTVpl1poNVE1dv
j+6ZPX6peeHsdTutZBVFcZKdHUOSm4PdzLE7FKaKPukAwChnrA6yWdM6jQ50poAz
TAep7mIg2HcYAaHzNiNjS8884NALmsrPtNFGSCAHP8+Q9N16cIKzL5JHd8FiLRQn
PKl/Kd3/R3CpJEea8ZSbCgciXH0LsvnrkpLBgnmNqkFf3LMbXk24WrVzWLEsmIA1
uccZDos2mVaxkFQvVFC9GzzxT/MEQUJo+LpCCbQp48vEvp7IuwEizFk+Z+xsy2HL
hyDxl9goY1wpZ3JxJUpZIIdQe+Xh9RGQTQXsnj/uHfrECK27c1tloG0ADDy52987
LNjYV/nymPrOTsRV4OzKadolRfo7ev8vXJb7eArjeCFsjAt6Rx3kQThRYg/4nsBX
yseSCBHBYLGtV35ubK8ehUuP+d+oeI53fRG/ClkiwsQ+PTULSUor+F1cRDISdo5m
YDr4R22NwrY11oTDAs8P1WyecE1YDTbDg3VAMVZItDEwFcbCzdRtY/u2iNRATCe1
KiahQcX+fcexJuXlCGAfv24cCOeEvZFNRJAdAyZQJJihaczX7vWq/Mmp+6iOGRQb
eaR8TK1dk/KimA7XHegT37nw6XPe5Eyb4j1RmQjn6VMFGmD4nIXNKLOKNptyYd/T
XQ122RuCTRbIDtWR6Nj3llcBZWKJUucbBe7xPnnlagDzLQPh7ZZRjvBiqMo6Y8CW
5ZzSxm2zQdf9GNhpN1di2996fvKhtREOuoWkcMNTM95XnI54efn6eBrsC6L/W1y+
ft0b9QOF4JCZq+YqIVUQPo0mxYL7nAMokc06ZwZT71RBjmILFFxgWLQ+MA9O8XGH
ChAo30edvtcj+V6FSs3/Ftiv+OFnKJsbF4Ysd4KwOrI8RUU94ltYOweYqwwmUwCP
X54jvicXgCVSLey1Zxz/FHzNihE1IhfHb1YaII0yow3EcF+o+KXviJoTG2TB+t6/
fAAGOnyG2WXvzPIWKor9vFLHAsBaBj5chakHkAqqjRICnSh2QA+iT9B6aQwUPl5p
HvFk4FKYPlPKux1Y7I8wTAvjzN2oi+qjjkNHPt41YSUEDgTzDIh6pE2ppuA59fh7
lhYofcyOmqcFBCV7opdruT13G53P/RdKO4AOiVT8UQGfEi7n1/lcxatEZPf2IdEY
8d6+d9+86PE2x7dCmYK/pF814wWDiYv4QmxpYdt853uWzUPi3IrozfqdctNT2YEL
47WxZ1POQfALqUicJ8/AaggsysZbBylQXvh5hFlQigMwUhTAdcDEjPy7C2gVN+Wl
4pPlqYNr+xrX82sKRjaaAeT9cCL6Ch31Z6zXzCV4XpjOy5HggfI63XVO7A3/Z6s0
TOzXVOCiy9rk1Cm6u5NwQGvzU85Zi8LD4cMZsD8ZPUVt9FiqaqfVeh45Mld4Qzhh
iT4lytOvOjGuNh4FNVIdAfo94JyfKTUoik//3MbztDskAXXaJnXYLDC1bRjUjf2U
NW+tDMkejMmmUP8JNHp3sUpNI7z9HKfPLFWDbcwQ2i6ATQu8Fw6aDp62I3piQXVJ
Rg5/FxLcCwDxcEo860xhMdTI/EY5MIRa5AT5x8uR52pGL3nSTy90tLb81tVgcKh9
cGHbui8TEoeBHLQOeGVqZk9IZC1UjZwTsvH94RTiyzd/uyK32Xya8ihVMP0jOvrl
k2OmXsFE2h+eDQEbsYTpQV4ssUyJc4KBFOban2fdOtOL9KC76xDbRS+asWsmTt+v
SALCw9EvvtULL0a4JCm8gdSAad54Xd1WvIXIB4h3ePaW1+8G7L6cnhkGvi8CWCWW
xqtsiZ8b5+inYPQx3t/eljdBcaWmOg9bfZnIlB92xsB8nxOqV4QsqPFgIYyGX3Jk
a0TDa2/eaDTAH6ntNW+X5LKO79HmBxc4BPiXWPMc11V1xrpCIOYg6po1SUmJzr0x
uyNxl8LPK5YqPOzzfXEwPN71NHIWPd2I30LWBv09jUDidzV3V9yOeYyuEDHeTY2O
Qsf6ln++GBvOLlAKAXomHMgPwoSV62CFqlnVBlLFCIdbqfIFieu3IbCYsmrwZkiV
bRQ/ng+Oz4IJvGxpRLd/yBX12pRWlXv57XCMqgYLk3Zf0WBt/upsjO6E0+QWKvgP
6lNQJQqAmsYbNQjL+6S7pRfaW8HG1ifGZ4bz51ppxSsOCNsQv1XCscIYGpY9+Y0k
zzU/Sj/JPEgQFVX0gpgfK1zM0/X6CRmgKg+Do3hKlGTpjmKcpS95LZCWJJgsaDoV
GpquLQ/Mbs1cILZQrixz81zQiY9X0+bQj5cW9nnU3AnoUpVqJbRr0xEW/NRZBOOe
CCcX/H5uOGwArqdXR7umEezl9uM4Tik1VnNF/TuwXb/+MGZmyz7bxVEO267AyIVN
mga3S3eQF9ZqzoBU+IUYspeH/9RQAZg/hH5PKGgB7PcURybsAIVfSHedtXI38Moe
pvB5WKKxZuMvw8JgJ/RII2SDuR9Ulv7jO0uds0gTc5jnpLYcs3nej4yKUkrXXzN7
yqD8ANvy6j5V5UUjusHP+wmvh+xZBeTw8IwNMr9LgYA7ICOX8raLdSvrPZ8JGqOq
jXWfBsjMPqTwFGv6cUoFOgdYE8dfX0tm85GDgxxCenOwCMSEk8pkfk12q7DbtLaF
Ee951JBREH70DFJu4fGxCPtFwXOakHAHwCEG9q2l8CgsX20wv/UiTw8+BV393LFE
D/P0J2TLT1SgBHcnVz739MsFGxO628rYUGXDTP+LEtN9B74wPFyxQMw0V29UnJWd
hJZmU0mj/G4+F+fUZNp4XRGgOfONjvNJy7mlca+W3xOHhr/FMJlJ9XHIXS0PpV4B
PiHL8WFuUlADZCAWV/lHbrbK7c1dW9/GbknYOw/adh//9edXOEGNO5rHAuiKimrX
OkGQqUJ6lhXnHt3NkF+9ueZxh5XNI5sduMX7ak3rokH51pElPH7P8q417PiTBENK
ZAjGMdXHhsrApnyKMi06e0PZ8z3znEo/L31B+RsBa2MrknHBMnpzPdZrisEdJfjb
djeYyMpsf1xnBMIVV0OFCWb038iAtE/JHgvIS/x5gLXY3L5KSSybrjRGDd0YsPWw
NvCTk9u8R4HGOGlarlPYcXHJj0gnOofxWkJEDAUA2g57MgIY6jBFxbalwVScaotr
kc+oOaMVDg7sy5QVx08OJnytfHsFWXtWgZYZQK8JgmeJQcO054fL7nMjEc/7fv+B
87jiYYsJEOT25tep97mW2/lFE1tXSEFGFyOhe2m8RAcR7qFux6OQmInKAVJvK5CT
mcI3WfQZCvaSX/ZyVtK7s/SCKB9asdRc9xVXngOFF0CEXFFKqr/d+9U8jmhBLXSL
AYbIeg9nPcGzEI2F4gV6CX9xCvQIUfmC+9kqpar0bAySo4gzJ9cBggb2TDB6l1jf
NLV5dDAuv4lBTwpjx+jGw7agW/FBf29EZrV1jCihbhvm28Yi3SdFgIEPYDjRcoJL
l8nnyXXZJmwuF8VBwGcpsiwn7tc7jg/wOFZ97eT3jJmJr+SbK1GsNMbtf3Z1p9w/
7KyyIvd2fbd8MztdvyrqR/reWYuUuS7MPMI0CIeppwFpdk1HnAubVQ0fN+ZuL/tz
d6nQ/hi4HqT+LmDFzxUOhITh4IMf75ruDvzcLIAWh15Qh9hqou7e4q7xg1kc5FH+
eeOe1eWK+9oKXBA41wt9UuE7Ni7Sf5xNrCTQ5po8wUP+J2z4Omhwm+ZMxlKBAFeh
tQBU3RidLqJUlsgKE5IeGMcp0pTDHTlo4CNMkcyGp/G58hSTfjJEeBQObgi0KgIX
sgRz8MiQAeHWfINEAdrP9mzRbYdoM77Q8GfkkDwlvzVxDCfGWSf9LDgqpyAHf+k/
WNX2p2GG7Y7bFbx7nHE9haDTTO+i2yCQAsdja+DtL7nlzYHUlaPh1A0vhPl6rZIB
5uD5U/xdHrgAxAHEMHLlHdX4lPKvLlwZAIaD2mowuXIC03S52nU3oYL4US131jCl
HRxDW9nKAlggqmYeavN5Gmoczdrq3zov0R8Ts/tT/gJkxFuEZLwpt9ChqgQ+x8zD
X4XaXdijZuJm/10Kd4R8e8uHKiTYr5IthJ4KpC9Lqip+d6ZnHkBrXfYTbXkptDZr
LPQMFxZhArgQq09qSOldRyYb2AoCgfBhdU2HIGoXQp+R3qH/f55ARpcDWC0037AN
yVv52ZxvttENLMFc7fwj1ePOwlE2qtZPQHXH/PO3SHz8FKBaZawPdt+C9GdHEown
xR2WlzjBW1yiTkZu9OE5uiyUbvq+de1il3bi7KLCQsAUsSGGPvn7I9d0+2yJG6wy
KNqhAzo6dRqZ1H8vXr1mSDlbzSh5mMHs0qjQ75aID+KFCK2C/pjRZSTIg2yeF5x4
3fjOSAI8mpRm599ShlBeM26el3HprdUWKkjXwVKEU020ox9HkkTaIkooHljObtFy
bIiBdqb3/C2jgJo8J8BKDA9ditqm2gio84/4nF9EMauLWZ0Xi1e0GJOAZiYQaAL/
lhp+2lHecSyJ5hJQ2ZyHQ5lM124E2WtaYTkV4STWQ+65w5JuW7qBLJJdyQdIFZai
GBa3J92MCFPPmljHCFvvvct4cxekPIEVWWynF9e8FlNF2GlULB8vxs2+3lIu8+u2
HKvlWO6f1/09/iQl5DLH146TymA9tTYKhnP1uiC9Zt0Xq/tcKPPudKwEir8r0CrO
u28wq/qMSPUnmigIN8460wCyFuNT1vdgXoQWHdB0LvV/1hUv8esUz7kGPJyBUGVf
Q07KpDVxysWvV4XE69uq/e2BQeKhP6Cc2nVU+fKDcWhaw26/e1xgsYDywnbrPlyw
kdV5gUHI9D9yH9rVqPBWV62vDTYE0+EcrEjxt1VWB3cmjHMYKYjyQDoH8W1o3tZv
ZqIltjaPJB20ptV4TYcyv0f71Q1BcuTA6/4dSmehXcbew+p1S2w7HbXltTKFWNwX
prux20Tx5mVD9TmR8via+sppEp22vin8d5zgSGUEDm/jaXbit/o4AN6zUyy+gyE0
jGeopGwrnI+OhtvWHp5/WJJa/0K3qrD6UvXm+F9ngvU5CNvOQASK+FZSXXYh22Dc
culEZc3AobhhZuDgXVaM+j/MWHsCNi+AmRAEN3ObQPEKZeI33Av658C6yBhwHEsx
ESYjQSEtI0sdXOjrYCUC38Gfh0GseDRVHkbXQwrDryGBwnl0Vl0Rc8yrBkmABCwE
L/PZFw5CMyFoM/wRhvcV8SZdB2cetJe7ncxlOqVKHwXqxsvb3mQZ8Q1Crq5LiC19
iMrCcS7tcdPAMbfKRZZQ/s8l0a5PBjzN2JQxmXaP69BmwkZVkNpcwarBj2aH7SUg
aZNmSQ4tR6vOT5zme6eAbIrx2jireFcpqutHsSI1ZGsuj03j5/bSGLJADla9ujs6
CzmMUEt95DWGSSfE0D/NNvfIrPmpgXiQWhOAePbVpRJPuYHHGbVXLvC4x3cBXoHu
tUoJn+UPEt1XZjiYf+6+7vI0wj80R7YBnY5gHhChdMTtb+MzcqtFH06K97QSdxgi
HUkIV7y5vTJUDrhNVslYFlmGtiPE6tnyjnHH2bah5HvUAMegpqJ7B8AaagXFbYN6
8JU/ScossCvSH5HP2BIQFHlV26hqCBhsiozS1TeuXi7lF+GrM7odw7GfJSPqzrH1
UV7J9024n1g2KswYanqkf0x05usbkRsgZmoqWdkFubZQFUJcD5//ottOVLTw+nW/
4VXiuyZ2E63jV0PJrL1/2dua9b8tgBEF4h+GzqrODuSWVbGK2JzCyAOaCnbRcfQ3
gFkiZS5QaFxdqOKoJUEZnRPQvBTlgRsUyEl4UFv8bWi2n3Wzd8rnA2FIu0geKxo1
QMy4ONO48+9PCKglPeEY48QaEq2NI2qMeZlLu0h/VhoaZxe/KovyjBzRz5QZ5uPH
xXz2Pb3NFqhiD83EK79byxR+qPRIIZkZqbw2ZsSdkUjB/SuKsJHD9yfkwb1NjeuW
y9jRpGc0rDnKvPAFD+J5Uwoa2PxNQqN9M4WrNGFoop6e/9FNN+LgBbXJpz2PnZM7
GYa0T6ioX+2XzBPKEzvn6T4iXGWzqepJmEeEeXMc+sA3Ocsz8bjYDOET3gcedxtz
76+GTdwMwm31AEvzInCsEWA610xpHCr498YumoCiA4IwSUVBtP3Ek3idTbjDh7a/
lXdlr6KfHBBday0sYUPTAFQA/oNGfNqGx3HCIXLjldLlXwULO1RMv8cLglAKMsnj
mSKMqcgGoaga5abzfzyl7FfbSrtd+Bbagz7lQs4M9aJtEVCHJUz12vex9/S3ofSG
wXA9hV9rYSVKt/dkiU5mX0D8lRiuye5Eqesr4IaZJ2HA/wPoyiJUNuVyzUha57XG
ppX9VzmSMx+XnA1F5/x6kreSI8FUp8hNBzU+fgEg9uNI8/TPSjLv8/mez+3B19rT
46hV6VNMutnsEbgkbgT3KC+WIiyrLuZw6DtB2CoPV2XwE4sPbmvWHD/vvFk0Y+wa
i7jSIrz9MboSn6CPtKr0hpwNnJqjSAViifWwHia2b013pnXFJ3tIeLrwcFoZo1Nf
huAdZ9y8sDUPBH+XsnZcchUE0nY0FsBHLuAAFRqtU/Ko3CV7DucXPCHhuJ62npOg
eEMnrYcE4wdpLtyeu1wCUMftkhWWbCwhOIOzSeiuDzMAefuIauzEtxy/CE58SB2s
sxUjyPg91eU4IaNVZGylI/9jvu4e2Y99+itL3EptuE02SqWDh2rJrQkG7LoSmPrT
kuKqlzBT3UUS9zx6qSv2r2cZmwGiyAOdZ7rBvtUJYrH1q2KTvUtCwen3wZcht0ZR
qoPSvUcQyCGjuFPqcuvBcGRabHcExkNzs1yQmJo32eRuhmqEX9yd++BIuBDJkspp
Suij3Ma+oi93bdLWJj8EPx//H1i9uAU9zOZwFZXfpPOvs+EMpMwwu+Y9LIthJstu
TVG31wEXEjjgAUmNIt+P+9DgWQd/flcfW89JqzSPyRasVN7jtL3nS+rzLu/7JR8O
rqMMnzfL/2dqrMcioIaytz8IIge7THghgUnP5GZpx+IjfKo6p3dWYghkzoXKwl/r
yUvn5gyQpIxc/qXZ7Td3OESD/Y/Q5ex06T/Smd0P1zrzW8WbIKq/oBbk9X1pExBq
NCSk64WrNrxddw4OSniO7f2X2tvUpwwUSaNoV+L2jVXCDYc0kjMhHYp3XTp8yJQz
Pcau9iDryNHRnK5iVGBmfSn3Z1MzdFDvokQaspYIfGFsrpMDCCm8zwLoQdJdTBnk
vkd/0reuxK6tPgqhdCcrKkIHQ0GLJlEQefjuYT2TpI5HqB5S8KeFuq7mvprH8REY
JJ+6tbVLJMMZBAQ+sKQ9ADw0/V4L0rYmDO1K54r9NnebohgulntMvzEXIvYVszDC
fIF4TNvifeA2QZ7l9gS3IaFzqZUfDz4Sqf/IFpsCa30kVMmdzbzHwT2J9Z0MuTKh
GDHSAJRd5/13sxBIt5JcIvswX81sBGzqEanjU48KdjkuD4PiH9QPMoTF87g0T1+h
bPUMW/1xmvgFe6pOgyeDnKFlTYw+FZmWlawStq1fXXWj2HcTb1Ux8TsGUd3Mb/mt
SFlqtdsGA/L/7gLXqSCbirIG8QBIwRXJEnSaPil93zkI15W7+DNdoalwzvkYVC01
epIfUmD+jyqLVSvOwRttnzrGmn7qKz1KL9PkumKZWGN9gLz68o1d9bwoLbkgooVO
TWByFZdHfzPAMxWZh7UKRCquOJt/a6cGT4btFzr8rEhl0zPSgvqUMSq8XRz++iJk
/qXLILyMQw5QRf4zv8rAhaFYi7nElKur8s4+AzUct08owW2adjFapOjqbAPZJs60
GVymt1+39Zr7UuTZ5TO3G/QeF3d83Acdhkg94wjjGu8WRp1Y9Uy79NsPvsZkIkgU
BMKllbE9lC+Il0EiDcUpsGBN9AKLIIGP+R33TJpEN3lkyPbuSc6ahfjEvmqsWiLs
J3CVZAgQ6df0Z7TI9oHLrle6/Yj8CGX3liLqz6fv8jQEVGCbC5/32iJFZIPlYcH+
vU+7qPtu5zB1ObNT9cLRl5/FEySk8LJXW2Ujt3ThyUvMII/icySJgSlTVvrdkKlt
VTYebTCjpwWiMDEqPt0F/8Qh7Dg53LksEjuRrUaG3HdCjgDNqerJQ9V1xp2C+lGQ
jN9Y/oqExKBFQNk0pHMXdzG0slCy1VvfaiIDApknZ8KLX7y9+IAjs2noGIhElhn5
RTPhUCnRedXRY0Umw2+Ivv1fJreaQFEpfisqU88SrBD94Bc2QCD/gOuLoyFxvadf
mbRoc3tIrwet004o1cZMQvJZJ15V8NZjBN3Xc1uY7zDCHBrWI9wfwHhbG9uuS4uA
Jx1S3Nje1XfMbcJGpqdjOgD005PrN2AwP4I8sRYa/xvMd1BYRC6wDBwOb4thUFKQ
8WGbM2caYt/mkkdYui/Tss7M26Zn0WY1LPcJw9xWA91nlVJkfZuQOcvVXp5Lmc/V
siCPNFqKVfEZMccoELClf+I+X0LKEKnb01SwvQI2Hq/DBhWmq99lT0j5mJmcSbYp
BIbFoN32wkP1lHkYik191mylWRndXXyXygkjBuuNwLGt9P4IVkuep7D71yCm7S7E
bqzz5XkbDF4PAWqS8ikSFgNHgxQKb214V3/RSUHXHPCcE0Md94Qfrw9UqKXH++VE
zr99vXY4bRWlhEAPCwz/iCi6kX7wEgEiV/oJvbdM1xVIYqN3UtXXu1/JO5J5x2X5
QubNGypP4bn7VwtdICeZwNnWKFFVWyj3CLH29hbU4vtuc9NQCuayLw5a02PobIhF
pW918cDd85V+4vPqFlMgvkrgdABq+b9gwtT0SrR/IFyz6zSJNz26KkqEj2/7mHt2
W30pPaLt1W8Mbro794lcd37CXgSyBf1d0Z8SCMo+C8ezAFdSQ6Eg5sDvJEZRLntt
5djKS1Iasaqa/1fVo2VM1Pijr2EJ/TKQ1+bhx2PVAqpke3j6osAi9pC9B8VSIbYv
7jduwmZjjlfeSypR9Cq4KB3ExPcKRkIVoyIorevsmaFly8/zXOMqS2d25Xa77dke
/k03n7esR5CEjQ/Ly+NagUSSqG71pMSdjgiyScwHN4jv/1UmRxrdZtoiKmZsYPtl
KT8SDbJVk6faAqYfBU8AlMlf00dpBRKHzJ+viw66UT9km+IfAwOZ7i+CdB3qiNin
Kx7QvnE7EyTk6wOh/tZCHdJy/VkU1KNgrPkWdePxFZSmJ6cgAgO4n0jgZlCMjOhF
XZvSSK6WtFFi/Uwg+1lHnUST/uftccyikXNfVMVce80xfniIbCy+bpl0gS3QQcTs
YuFo3ADDrqJuWAfxIiLyMGehIRzAbLuVGvM+8TMyIx5Tv7cPiw1XVg+Y+9tby5+b
WMTxvs1GVzOmwOFCvdfVNLXwnP0mPsdFiEjOdIFiN8vngyfUiPWVk83m5e/XTTxu
qxHzcv61kFF3xH6Q3cp/YEyiNYgWBdW0+SuXX95TsA05JJ2x+KYl/VCFKFqNMwTN
7C7sxhY3h6Kgtx6dktyzPk7psOIJZuSoox2lBbeDPO7M0qA56PgtFWRPtPBGvrIp
fIq2xH6DRGvjRVIs7EhXz3Ci47XFsRKLFhCE9R7kf320WYq6LYKMg38zRTCeE2/X
uR+EEyEGGT5U30Z1wew+q4tuQG7F7+nVqn7mzMxpNMloNOxCEBtvrvU2nHg2PHfS
c3hHCaAqhFeDB19JOQeYsqoo7xb51eFGeyFQKEziYFFWkVy8nZZMDf+1q6VUSkQa
tbRTamcrE36Su+G0ajngmOa3UFW1r2sTsmKK4gw0jUOlBG80UgYd7nUa4EFf3j7J
SHPa7NiGpYj7phiW6yxMcKLJnrFzme2ox472xQiyzyr9njaO3FgOPXWUVoCSELZ6
q/xqB9x5Tk0j+4rjlvy+syhUJNkXQLWLXDAfA1r8no/LMztLSyk/Jg0OSCPWsLV9
Kln7k0+1vHXxikaZxgPjWQwoEQPGxi7WRprsJMRMnMRByKKNW8kNnG6DQvX8BZPT
vw8INI6lN9nzvZO+qZER9FMrly7JFqM8TEuc1b+/Uv7ugJA6SQeoxKI3QccB6aiK
/2XkvCsI0/bZp7CxpZrZccWr5fmgKGObcEyngA/8kweFNAYwewxROfwHTzyS3iOc
mMiO6AjF6/4ETDIql6kFAUggF8lOiAWMWwdK/aGB4mixgKSKoBWfg8sU2Z6UL+rA
8oRMBLV/ttRPRctS7+2+Z9yD//31r8rSfCTmHL7/4TtTcKbPrwagkUL2GJtKTK/v
KFGrQn8tHtmgsSCgQc+5XSGRT6SXz7wFlFTb3pnR3TEbq+gdcJH8RtZJOYWCUetM
16LJ9Of+uL6jkNeBDayKFM/CPf+VkFHDYWLd2AQgCIPC4UTEmoc1YlqIodoM6yWZ
PQ68QQb5bUuy4DCCIYKIwo8FNYvT7TEHjl4Pa5eDmRy4FENHYemrRO7X8RkcMxjz
ENJUpM4UoPrF76PWt3dOHrxjt1agKNZDEYKmmufDLYo7rfs/zCEpQ/jcvzd95PyL
GkyzMkfOY/1k/dJiu3DxP7z/aXBt/kMyoxZFrwr2OtWwhMM0fiITJcYID3EguGmp
DhnYZS4vi7L5NypDeeazGP/EavVXzbiy18JVbcmFpqwSFZdu906IWvAVJe9SGxxn
1SGrvyekB0m9mVg+JkhnzpmpGtXWSaI7mKBSBvk698Gx67RUrJKwx0/lfMtkP5vu
LsudpP3aMUS+azF8l0rNZZoj74coSvU2y8sCp9IH88e3Vgkw0/fNg0oDy1x2nEZ6
dEiO22nRSXZ3oayDfR77PvQdLQ+nJvBubFRI6Ur3zBn+Te9TuhLJ4Mn7r6JLxaFq
z7lI92AkWvpDfSrloelW46xsi73Um9eTAyuaJSKgg+KE7pzTEiqxxTBHlDFn6jZX
Tym4Th2sJkO1HVqLMIsqZFTls9GJWNNp0lolWulD5Tcfb7YJA+s1ABTC0Wo2+9G7
Ucwe2PQ1JKiKuC08eLfs2Gr+SU5BXoa9OZwdTm1c52Sf60tQBrKVCBQX3bfrqt+S
2ZGzWzhJ2eFd0isbl0fkx4nZRSfobZFM34DzCPjSRmKoTBV1VYKZX71att2mfn8M
nWiHTFO4qAHWQPZqdTY/qcMn8sjcwrwHRbiPY7XVwAm/29nr84J8ug5z5BGTrvsC
0eSq7F7QORJr0LHF2+YMMvCxiOguDpWBMkSGbmBXfdts8wJZKpmUVUBXU+5vh/LZ
2H2Nuvzax8ig0ev9Bp/Og38w+YDXa9b52awk9QpCspjb3jrsK4YaY1URd4rDjlaJ
0OKYruOfudZafnE57DUDt3WyMcNJuh987nzCMPalsdvOA85gPvNxa4c7wDHCipBC
lMFJQ3flDvF2PGa5kF9dVwsiIhUoAy/9HQSU8Af9lHru3TBdXyzQTqPbm1GUOD7l
xFTk0i4hTiokTwU6ik827EXjGWO4hoz5H5AigSg+VouuNYsD8SguW3XPvVGPgxei
faFKTzJAcIRCei5MNyeqJnhD2rBfyTlvwAp3eNYOymi0WiWWAPd3s0o2b/Rr2uzx
qFUSQXaD+ajkJc+ha9OdXzWqAqKxNZ/Q1nO/x74MIHQR3E9VrQ078wijEF9ZqzVF
X1RbIBH0UrF9g4y6gwZ5VAGifzKIXmud89EMz91+J2EJKi9MQszvmwaW4hY9W3PE
mpznR4nq4+/XEIpfxRvGWT4axdGs+QyW7if5884rVy7KWodeUUXqdghnOX9V7CXx
FVYqUN3TStNYkx4DrAioTsDiggsLoyGQdUD9dz+iU/KUklkeqCWJzrA4fTBHXznw
yCXh1OeLKfgX+r45HH3gT0PomNKc4JB0aVE7xab06BhY6+610cX0vJ6/81KWWdk0
3k1lcZR032NkfjKrR48mGfXkSUuZZC0ltONRpw/2q7WjrW2i2XUppcs2kd+VZWtM
uBue2ZxNJ0xPVIKlgbECl+l1vZTbgpLG67K2yNNtfSAVymf/BZspvdFq9NVVR/tj
YQrH4sVxh0h2TnEk126ehN/Nbbv09KZOFKTldRichBZLDj0EbvdcKKBhpi65y/Mw
zvLbwdk1BFc6sV+27VUBEYeeZZMfDz8dmOfL9dezEQpooOlPAZRdaY07rBeha3Fd
27m0crTx795/PvemQuHYu5ZoYVEDXJccfNcRHjD26MbwnJ0InRAFpgUgcj7P4Hhe
Mb27F+e5XqgW/ukoMpRk45vTtbfK0Sdo/oHq7ESIw46KXP+R5KQAwwJjxvmm5e2f
qhH9wMoUBpki9/DxuwP3c5XwCtOKO+txXH/tMLH5wAy8ZdmuQiWgdvlTrwwhMl+B
KYzcv6j372/Fk2Vnirl5OawZ53AGXF0hrwXZa4LlN0yvBT8NDfarq8NGZVQ0BmYe
IfStnx5V3KIF+X2EVCXVTN9JUcRJtGzNWy7Ei+1JfsvikmSf/l5e/Z7A6KRW2MFN
tkzVAXGRR5Aub3GBALFlcE6gquT0KmDDq0cvW+n4CLOE+vYZxQtPFzdel1jL6Ayt
3P0EZboashX7z1PUqVHmq2/2D8Lp+B+a37sszyHmxyN1wbhvhvM5to2VYdkhw9PO
mb1iACHCshJwbnQjDdx73Kebowh5nVDCSS3LS3X8M0gp+h9zBY7CSfbT6XWgV7wn
R8XwiZlJgpzb0gIz0S7ETUJI+RbpARLRVyj822Y0kKGLv2Clr4gYGT4lwlL7IRsF
4Xc1ANnxOqlbine6WRFeLZqHoZz06RT0WUygvv0gOL1Xmot2qE8NFWRFMYzepgJZ
XRgDGraXwfLwd8okzUPS35gyRc+qSyze1ULbMRFhIsZzCWKJgmBxaJzYFOzp3fBv
pNxztZTSoeQGnzeXiLg3WeZQzswrrkC3USLsH6QN7f6drRVoqVru7l8oqjxyE10q
AyYyVqUpaQIaIKz5d0nuAlGFhw8vx/y+60V/fCqZ4Th/VP7HiIJ+mMDVCHBHKlgV
l9QrSiw2sDf2QmaTCexp7v08CXM/thTy1356pQEJmv2YBsYrbQhTJqG+sc/pK1Zs
xFqaDCFugpPi2LPVHdf4fXJV+6TmeHg2ridtMHwzOh92Qghkl3tzZKZgf9vj9rlM
e/2CXdhkgcc1fmSQ4kv9iBqq7mzflZ8kH3aweoUPS3r9RPlwjFu/1h1i3O3W/QR5
wdYb8BBwltPBMSNw5BgUoCZUytKpyAb8OaYzU5EmYCqRzz19GtLIqI7ivS7ARB6w
Qa+TyN32FiGoCwNK9dfh30e2Fo0VpkGnjrxmIvOZjpYXpyBfb4v3GICqHQHwb/Fu
FgYXxz/zRZZgjTiwj2qC1XEiCYMVLTx8Av0017BOjhUqPNiQyAQ2MxncXsm2msP9
brSMTQIG61DuhZP//IRzeha8a0QDM81Ga7NHRh4bbkjRvp6/daM0waRbP2sF+rLo
MqJyl885UJsgM33fJTGH3v6PWEBkqmgB/kGEBkfE32KplmwuNisObyINQadPmUKr
sumWNaf+cXy/T9qW9gvE0OSmAYrxUOs6PS43pna5YFU3bB6F1ncjzMtZmjBUJEmo
6K73cwKugSbTzSNr6jBBgePPgKRRmsSUjk9+8TFMccoodhO4Vli1ge/ediUMchnL
upL8r0DPlZpj6Ia0yu1j7OwirQ1GExFqpa5zQKRydMHP2KybWhyHcvf3e5PikSyZ
h3e6jwnUhR/JbdzLSRsl8RaPYxfFs055fSQotMhQv7OZL9CJLbLMAhDDd0OQKyN4
sMNtI/N5gzXe/8gJQHBYy5UfKW7fUsobNzpQv3JwPQUiUv5iq7lpElgi/QWMezeJ
ofCkud/XteKZRWqonvcrNTP7lGncfpVtbbZ/19XfL6Bk9+eoIfriQL7x0JByv//x
HXf6eVEmnv4mehtJSCAqPrBVSzyWIleuoWM5JQqXQ1YBioKLJziiYaNKzPXitsKI
tFHnM4D9J3U767t70DNdBTpnA7ACKCej45tQaEtjZwuqrsGTDLERSPUngRjzIxqB
9bPGmc7j7ZEfMCdxdfxVLtjyOIhohGiSymQxALgDaVc/mCFbmgs2VgCaGHz1Qduj
rW8nCivQDO9GTQp2BEYg8sLCp+n0igyGpXIentpHIOglqRg/cX+2n0cmlUD4RtUH
jl+h0ce/zo2wO5lG20KahegVfhQZDba/sH2CKuFN1Jo6Z1v33+avFyF7W+EUimqo
jbSEp0hE4wgg7XMByiXWGsj9m6buAr27euGDAtrUonj9pfvnpjNk2ueatkrtVQi0
gFcxvG6rA4vY+l7b8C8dZUOYmHtTUijBChYLzYhHpDC2ry4SLCbkFgoUVNxNNXKB
7CWR28m8nrFZrgVe0f+qPEhkhhe8OxHCPsM+R0lGOIrMw6i/Bzejd4Z5tkeKxVxL
veWcCrpKpvmzyPUpPn2XTj6Vm+P7q3jEJh6wNKL/jdDd3b8NxnLYs8RYR6IgByWg
Ksmjf1dGG8r+AvqIK+SQB7GDHLSwGFfW8UccolwbV7dBX38EaP2NorRpOouYhMnL
jhoUhydb7PYTS68MpZhyxAUQRV7+eQEIuntiIrQOsZRWeYVXe/+NqUUFImuhvJtF
17/1eQPxx/+koEH9aktPd96z89ApKka2vg0Ovo3IvyzbYJbf2ACHgX6mUtFUs9LF
D220LH7GR8fM9S0Df84xfBzpOowX3GHBNt1wSx6xuzKCy4uQRbq2pv9gZfxVxBcX
afohiE/4vP23xai6Urpmgo2vK5MBTkN+8F+wxUKz5c2UisrzAWD71YJ8h4Rkn8/b
0LgFemEekVAdX+kGlty7ApgCdtuh5bVogfwwZZprTIbo0/8T3P+vvurUvkUxrqxX
VPayhN0HWZl4tm0a3XwcMbq8VfXnoFeqBl/Gcy/XNHcV5djEXWKlLDpWf6FSTkIT
Vfkd847lJ5MB963/pm9AXSh+Mo1KoKyVuTRPHWZCNgE6MXjj9h3wqMNldm+T/bsi
boHqizNzm6JTS2XOHe5FA2LHjTJx7+LH5v5RkLgdllKPIO0b+ECaW+cVSFk1/Z2Z
cJ4WpOpKnBLcO5fZPXXf8Dq6B2WTERk9QJlla1TT8zEpqB2fTwvQfLzv+ba6VOvO
P4pQ3Fd4cvU1hWWYPPTwJsx3tIuQZI4W7iR36+5UouBi2jGZuYERHzXYw16B5yzy
pMbcEbduct3612/jb4CfcLlVd6yp53YzfoBtheJtnGj42mh6Pog6pRtR+d1zH3zq
r+vItVXUSfAz4D7HJd7j25YRyd7oj0Yhggq4VEwecsLqq/AHiUVDcRtKJQTPVCfe
XhfWALhvRfdmhckKai9C0V0QcOeGqUFSmX5YVUmD2jTwCAWwEdpayF8lnfafB2m4
0Br1bVZC3i+gfxcLZInmbvPKM5480fLcvKm8l6cPFReJ9Kg29pgg4Sv2cT0N56Nc
nuE86wYoJxitVXDHiaCOM/hLeTyQjULPPsm8ZCJnFTkeVt60agozZrhFwl0Of7oI
0pUAnUcoVmllnIsLnJ7yMahe/6uXQaN9zZT+U8GPCOn8vKfRt1rtk6Ltlq6iYTaf
nEURb9z4TTJw+5ujTdZAbQdRbec5mdQZ/NhTU1nf3HWTHdmIwyzTs7aYU+lbtTMk
kfcvj6XlvYmTkJ2XLZHLNqrDLh3sEEwi8WcKxjqvQYc0f1AoFmTe6Bu0vDi4c5nE
v9JAIqjzZ0pbYHNin35GnLCG5bW8xe9h9hwiMRKUlWgGw4XETGNPyETKM6AAUNfh
ONdGPzpjhcHHtxC1Sb5arONbMTYGgPy9J+I5bvHsUnGNu7d2NV2KgqXXZyVl+7xi
FNI8TegMbGyQSTlHd/DI7ItvFq6Z5NVQcJdxNJqkjRRtQdgdu7bV8dhoHp7p2Hb9
CwI06elmt5hsge8Im+U5sYt0wvU+oWdp5gO24I8FVk3uQTwu3u7MiEIl9ljzs06x
HMhz3bpzy3dwiwHEsZYT3+o6pnkAAPrNCm0kXn1Hl94w3/mzOvdfVji1uNKdxrLU
0rzMZPjkD7uSosDufDwwItfAAm2sRLmEOkTfc3ccTvlRRNR3C7r3O1GAijm5wM5p
5Fuxv8p+9i92Fcif1gOHkexd8Y/LVGD8w7qBPOBndE3Qkao4DHXWmJFMDFnTAS6K
/J9ixa+Q0lSP95MNtXJy3W3f7pVzhf8A20c1x7U6jZ26Jq4igjj6d4OIDpLJC5Lo
ymNMOO0ASx1L0eUeYFScMXJWaw0EazWnEgmUYpBbIRgV4N3RVgxIyCBrN9ubKzYq
cYWL78eGWW52fD1f9pCQdrTS5dqZGVJhWGILazVTcQ4+q69FUShHjug/cKdrrmEC
GzazAH0IcNMjaE05Ycx7nnQjSfGvFnhXWPQJIxUrUj3YvneToNhQwocmwnNlOWH8
R8Tes/KOyV6VffoqHgMMcFQFB6nw2rmCccEarq3pJMaXgnEnlOz/2RoKYblDRQ66
GeGTlNKLOKNL4oiF+HlA0a1ZUBM4/up9TV42Zy6ccmDwZpyEyo8zwylrElAZhYUq
cL18VAmyJpeYQmlB7vvZTVlo3Vg2omELMrLUMWaUsf4ETwwhK8so5TAD3hHrFokH
QbPwU8gw/bCryScNonqg3ElMPzaEGOxoLi1og1mLmMHl+E7Lih+Pg6aF/+cDqNse
iXkSy3PgNi8fhj4xQ12+fqrP4rJdBXCvLxU4VKPb3Hd6jOgK0k09utwaJ2hILxxt
ihwvju9WsZsMonxXc76sHyfsgX2umRID1r0UqEye6XeKlDeNT8zJMw0VxAb+HAUN
v5Ot3Q4/rvsYe/VYC4ZR9B90ESbZRM4lq4AsQl4m4Nj97tdrnZwGwLU9qckPbKW7
b5jatT2NG+HM4uZ9/n56k+EJEegtVZbKxLDpSpQvZyZQQAL4WwdwfNirwfNj1EYn
PSnp37BFJ8jlY1xlomxbjTVHlpoLdyAtqLjN8O2ZxKU5keBWSxDs8GTgAp35D0yq
FnwkMPnthcWcuPL3cAXtSRFQi9TJabJWxpxq5kLA+eYTwAEy676O12tDLFP4o1vs
JS7PYU6VilfUcmGK838cJ3vARUbOkaSDRQnTbd1/xn0I4LnhTibj6CRRh+w/HM93
oeovddrA32Eaz0uM6sGCRkW2mXWjJUxj0R1Htd4etYSGV2ACB1VBfXO3GaBmmyMa
dcUUm1hzkoPcMqPsucMjI9YL6e1qIQ52iWXPfLK7POORG0gz3nXGXfznWLRj83p8
kGdh/q4LYC91hwSucD3VGgIrQ/XmzRbWJc21i37dJdjEPfL6Gp3GIzaipMRdUP6W
hJoAFuYiMLeHSMS05sf3GO1HFQneAyM4WTTRHajJFxZ0/RiNQ5ZyP4uPgt07r7tt
dB185voFPemz2evDDjlnzbaUgUa3oOviMrPPBjKVNewxMuTbGsKs6zoqoP8tPyI3
KOuDe6KDbtgXuAZuqcAvoXd79smAxkMvvauHTufkaJJrfHcbnDFXfrsKTV/HzJns
8UXOW2BX88/V+FP6/QOfq2VSgV5qqkvQO5wnEnHXPJud/ishsMH6bC55GhUALZkX
gAjKTymYUg4A+xYry9ZqJgZ0IjGym1Kyb5Sd8igmYLKnH2qMR0+MJ27qkSZui2xm
s7gGU6F+24H2hUnCsykcMrskXgitT3/gfu1RLaEYkYCbtspJv7MziRiGsfDyihlz
F7DYAf9MerrYbMNJm17rM6zulLB7SICx1wV4iuHWDey1aoPac4HWSyxbOwgFoXvE
5DjlUJMfrNzSvd8i3M38iiMVURrXI1Ok+NLTYpaOdzuSOhR/cRVRSKTgW8bPe5tv
+A1t5yfNJLh6wSIR1UjheeRTQ8f1thNVyvDtOf9jseZkXhR0SwaroATqGxT9O0dH
Pj6jobLtOog+GdG+8DMiWtIp4lhB68YLGAWqRxb/8nwaX4nSRDxZcEd0Qt+b8Spp
iEsNFHXbF0zXB8AxNv1LAQHgN3BlGaXWe+GjV849rrj0Wt6012EyU5HUiAN5He/c
uWGHrNtS9XpD+LPTehogJ4ZEBCN/dqytUyOT0SDIdC+MZGOwVwN38FxRlyhNVnFM
POrZ7QkE0nPI6JumhRYahItTAbF7QEECE1xeLK1hcjxbarQJ9hCmoQ6mWPGN5YZZ
L8VHDepkC+dfVb+qnZIIk7ed5JkLONxn1mgQnIjAx7ScONn/fh4C7/OUbFnMHT3C
LFWQU4Bm1w9KAiPDgFBaPtgnLDIgp4dkOa4sBe4J37ovOz26j8zou9Zw+NOlzq6g
xrgvfKiirXeuV7diCuf9ITSjyQs+NG7FS3IiXofZhSLOvkXvS3Cy9wOwqgl08jWY
eG5Lgh+CoqDwhaGA1ha+JiFYks6XY7bhbNxTzhQBnjIQDbH4mx9WiiaNu0SaE5f0
jyvLNibS6LChHPSqSzp1RmeFFZaPw0+7SzgCqalPFpTqdWryPBHje04CKoYDNSTl
8Dtr8/hA+jOTkUVd+cMq9nf+zmD9phgW2DW3GGvogV6pB1xs2usrpS9+KOZmfmuy
BYpB9HAEvr5hkoZPOhygS0f9nmQKOjtK3XvZaW9SKfvpCfOsgvHYetOyXtyn4Q0R
H1xDZ2kxU4OXntfxowTTBF9MkcXvVCkfSz1dJ8UhIHg0B1k76XlJbKPSz3Ve6uMQ
9WLYfb+LtWdHB0YoBnMwoFMojQf2CPKXqcvn0j4+yudeuinPJF7rRF8S50gz9g6D
tgJ01s8hWtuEU3k6XLU/PbH9XiCRambvaQBOMAL+BTIS4CqwHWzuTBrFYsN0iOi5
qWyPEP9BnpV9x0NbQVVPS3aMfQ7s9x4kyZdWdIzxDHPC1hymGBAS+u7oFvucryzh
lqKoTMG1zXQ/14On9AXJouo1pnMfFP8KMaZG+8cH/v2xLiTbmAI8qmvIg3Qtbwoi
v6U2A0py8b6zcyWG26mq2xHeE4VxSB51SJh1bSSGWCt+n7ytKSoa2he01dSI+MqR
/7HHwVNIc/P0ENVE4R8BV36ckknprxRzZwVM+pvKg3Fe8mztroNta75FQC0jV8Uk
gjtHX3VTuSALKl3dh5XhM/CDAdINyN8AVBUEwPLJkCAIX2j4cQtIT3RzkS7ALirx
rwgI2s7kqfqYHzCwoR7bIlL9x7cx4jaaiDi2TfXXFMPYhvX0UhWIxnxYpdX/Itsr
n3j1Gq91yxW8kJbrKuJS9QbrvCFe/CTAMZVb89FpxJUsfDYzAZPupZK2ndLkQ0Un
P01Pm254qm6RjHnlupBp36dWjmbpIkts78y49nQgk92Hlat4WrC2BcpPoVNsCQA9
n1HEQwsRF6064FeFAaElBc3BV6cjdweCOeFZ2x4Hz6tVVaXaHVmVpGx91HLBlRd9
6N7C+bf0Tz7vl+585zHZ6WH1jCkeoYk9RfiP5KvZPlmGFzR6dlSt5EdSr+AP5/9W
0d5d0tzJ9WewasHmOnTnRTticKDiZj5wptb5ZEI1a3OuFFrK/vk2Uvw40EbRt7oz
ONDzK0sKSe9gtGCYAGjfWV8qdv5hSurNAh4xyGRgSjPe9EZb+4PRtOA15oxLKRse
q4VXD/yoZBGEOqs1F0qTlpd9K8w+W//mZONvgToIRrKEaKH6v6PfaePAa0vB6dXV
7iKAwodXZNtIZd9qLJUjxD9yTwBDUhXhtVBxTW0yAvT19b/sCaRctr05hn+IBfty
e94zQfPLePX2P3r/10Y9B71ifbVtphlE6QvhNqID/YzqsoOcjQxjYaX1jV6kPF6U
z0LK6E01jBRXEnfb+HkpCpdfmJysJC7FGiBds0tUY06hQvbsjnf4mo/+Vn7ncuhC
q7iats4Hsb+wvTXcHICKaOCUzEY4Nz021BJmYJvg5B9ZPX1xWdfrnvT83l2Cel7D
Jsy4K0G08+YL2fefxTNtj24Uaz7GKRDyX9NXBeirkbqOAS3yvZiT4/tjOUidjguw
3grWgPsnp7jyY7R7M7VwJnx+uGRPWhzEPgCrFt8BXQZiZjLEx8E7b1/Z+jPHwUZ7
E013SYFtpSr9WVmB48MrKFaze9pEaQo5w39CxaFXjuUuteNCR7WwUYlYJRzUeoAM
9oQ/ONd2bQiHPsIB6CgcHW7GJ+2GhUbtB+/P3vCW6fwtrKb7KEOHzvO2MTVGXzcd
NI/zzG91qTif3EaUVYMWLSjqS9/BoKE3WEhAyzUkh2GxKlHCGeh0t8wfk7SZeQ13
Oogj05KmFuI0IstJDRnQwsZIRmPkSVbAYIRL3BZrSDq87b4nL4vYV4GN1bgWBK+W
nNhMd3Pp8gdTPyHLuyKvy+UYtTLACTd+4NDpeyxGTn0yzXuSA5eTKVBtaUaFXLJZ
/XkIr/ONcaLsnsR5m9jEaYxzc7j2zNvsNFIPMtiuFNvPSPm6fwscyY7UWzwuUJTf
hkkfytm8xQlmXoeaeP3D4xDwo71gpviZEvIUqVh5FAo8ER+ZHjwC82NxTvIeTDza
vBbtuNtX0S6ZQIxruLkTFW7oaxY/LbIYRNkTQdfjY0oVQM59sdW59PUouxolT7w9
0PrDGVeqd9/5yWC7Q3EQI11gNQY8MtwTnrBpZZTOU+4GMuKUMg2JI/Jog5U4j62e
SI0zbr44TM9/vms25yAO6qHA6g4z7XQ4vtRW2FwnZSyeBIcnaqW0ywwnFOMfS9sD
JOwN08nvspt8iAh/0pny+r+MvxDD6JToI3IoZM3l5hwAQT3M1+rmCntNlKh+RHlo
yUxaZYLrAkrGA9zD/66Xmmod00t2hO16xutpPRV5St2OGSA7HnShrM7bB05cA5hE
tYyf5U/+AWetEYrhP2fyuoyyvreK+RFoHUqRjqPrwdlDnhzIO9tvz4w64CudaVWl
MYg5Z+BGD0rxjY2S7G3+dt2QQeX+v/Nu+YaaRiCpTioAXXddnmCYTYVRzNiPpX6q
/xmoHPQsgFp4CyWIjX1BbHmDO60vpdxVcfpEsnhCWDxcqNY/A8taM14kzX+lO526
cEE05ukUwBh9XQJiuACg0WoJ+xaldnGs50kV/piv7Ek8ook+K0+X6joks0WVgprb
256YMLSUhF/+CCfqgN6b2qQGVmes0Zw6Oh2lXy20J2Ly/7CCF5IneBx0z12y1C3a
qF386noowoajh6YGSMZmkP/Kyno4HKGn/cnJi3eaga42dorgsWeGdgsLWd9aVD5Y
9CunTMrlCCMp14cTTlfvLDQOWhTF0wqEIZQLPqJAZKLvgObeIv9DFxRzqf0y5VbI
/ia4Y/yC+PFxulsfygK9v3lM8FPaoo6vRGcVo9WcgHT7PffBJXrIU0FN1CweE50G
t8TM+1VBv/MdeTdk2WFpGrR849Xq3Wh00YHPazqIvZVeObOy3V5ndFxMJGeCaNec
+wTEnYeioRI2Cw+dtclZJ6oWzZeoOHmA4ZTF0zYb5y1YqVLoQ35kZlqmjcUzvVAV
pJhJL7eQXneg7TqvNl4DQGOjeAqIwmUVQBRoHkYKlSOiwB5dzC7GgNqG8KMDSgCl
FzOvo/UTCkbaIlIV+W5mD/R7E+fyqrGitxcg6k/+EJZeK3YPB9S9SlGC7Cr2n3u2
btg86Phv3OszG48DwX9N9cPo1e9gJCI/alvls81Dl69dXYdobwABzbSdizZCFUNS
nLvvZhnOHiue1FweFdNekXGUObs/bQjWqrmaixn2xDPF8oCIsmeLHKJr9jWE1BRa
Xb1VO8s7J4+CUPGW5/Lzk3BL/RKqRGuWQu8drE5xQVp4f381IVrrNmQV3vY3NB96
ozFJ7vM+Itkgb4EtufDKuJmYEPtpR3jqwMuBQqrZpyQ15JPGutBVHDltfcuU2kPf
nP9M4NC4LZeR9lPjY3An1Mnt3b/4Voqa1kfoaCSk5W6D3NbkVaKogW15IN1+F+Hz
we1MMzQUXq9vgohPhlenMY320+yArGtKT8+herAYdwvIZSr0gcQhkfEp0Z6gfL7p
gxGQV+O4zoFewCxS/JvfE6i3L5PP/hqVAW7OR65ulHKwSJb+fY5p+faOcDexUnD9
KrN1A/uyLS7/5gRI4nZdeMeTRHGO5AKlmJQRYttoBZ9997d0w3r4aqgAYxEopVUd
L081NFomhUF1UQZOUiqxizAnSnjKXuazmb/p9ClD3/odLekKcrI3xbeY1VCyW802
fFxHsiRi4pDiVTtLw3nrA3CFMNlW2KJ45TIimX6OaV7f1Lg4bhQ4n5qhSgjjo6KE
2JxyqRV5ZLsysfI+mPqZbFHU6WxRJaHSqowwT3F34ihwkt/gcUqVsxTNIoccyAJl
naRdK05TIfp0BKxvfYOoIy+lFbukAjXB1rjwgP0et7VNbPmQDUR5cBzv6V/iAqo1
SyHIY6EOJXOhI74NktwvLt0Kx6I2uHt+Tj9Ma3Ij4NPyK+77fW6WsJ/V5J1yLPqT
vUpQ3nt6Rzmxx08zN0lMA2r1mTfUuDruqqOkPKFnDwdzM1AFw0Pwx0vSAfR50G7/
TTIuzI/9qnnFlKe8rKdmwje8qZB8cDaT7vKeE7VuZgITlFGcIMGp+Ko4LIXng0X8
iGChCeBvn4jd2nEsISSRKee5J/LP74c/Krw2tCH1IyZjAehMzd1/AwfrvSKhjZGJ
n0nqMcHVfrMgfcxlMs1lVnj/W86rvDiw9u6k2d5X3YZbAahHbU4XryM8wJZ29tbC
phYqkRQWxJ+5VPnbPrWeps4mRrKKCcfLUwS84YuWYAudTDuxIqEM7kC7WUqyD9vH
/O5B8TB/VAshfV1uKnNzmy9QxSp8lXBAhRNjPW+WIaDMsYB0kYW+xFGBlc2qKHVh
LX8dDvTx52VYBjoPbi+gq7vi0OBIUvx9NSnzz8WbNdiqTGax8BYRpTtIR4AHWFtK
CGVxKJPkFSkWhS3hPdb9rDRMc2q8l6qsyuInx3SQRgg2ONG4aPE3a2Exk104SSTo
twN4pU+drm+8WHKwzZqZpgVQvNhrCtjFCB2r5xAPNa+tV7JWi095Nk6Xuesuf2rZ
Dlt2Au88ghf6ZZT7qBvXbXT2gyVKurhECVbEVE9OJwgFQTQ3cHJwwsA3qW0mC0i4
dZ3ASP53fh9wL46wElrI66clCIfg2QfDRkna3KCScAgbuhIOUbeVKeT0igQQUobX
tQHPYy1WubByBu9on/hrLySDcc+/H93rsg+BJHR0U4u+reR08wJ5A5Fq62rXsaFH
6WRwEVmiK/owPPd32YvjaXFWvghMqjHfbEoxEr0pZJDPxDmJjBzBjReo1bxIc6cC
rI9t4d/1iNpo2OxQQ4FIuMAVZ0cn3hEGCOddmkJDZXFcE5V7GAQRf7vZu8zzeL4J
uQ1lmS/LaFfVju4f8mQJMzTa9DXiWxMZT6p6rpmvITQEn5vqEupbs9+mrztlbVjM
9TgVbd/YY7L1czySehJ90EsnLiYAnjherebXv7TaEofbLLUK9RQJVan+A6TdAzff
LzyEe3H9SVYUgZf984RAOiwXPi0/yuen1yKB0sAyDaNhjG14HiNY88qH0CGPdCH5
RZNQQo5GfMMDkQsiGV1g6TtgmL0xSLTHQmvIoMREG3BbQ65AmoJUImsUVuySds92
Ep4WmAVyR+Fx/XzNP7sG/oMRI3ZZgopjvEESZWzzgSl4bfTbCHSDz4m09z2b6Di5
0DfzksX2sNtgY52xPS6KgcOcuDSjCXlGFFtXdRhH2U6n/jWnubmY9CkUcCoA68E6
+N50NBVMzW3Rm66lBQTt3LSIKhrPbYlnvHtngBaEApwNrcdmd6/KQLuuWnYtSeAo
nZds1+301pp0tXu+6eHwzkvJ8+m8xJIurcKKGAQS00KsbFR0oZrFdD+ElUVZpOVT
JINeMSqunqpAmgJUoWyHXgO6VwwnQq7i0ajxCUsDYChpBT4xk0a2S7usFIMKJ6oJ
KbEEycHJs7EBhT/1i7BVy0GiWNHhB+qkfv59uInOpppjqa81PtjM/2J+RMRV3TRP
+jiU3rqQ9yn13vxdEW7RuCUtx3xrQbm0Uigks3+fPoAWL9jYQDxWkx5/5ZmI2hB7
+W4nUxePXmajXlR7ossDCQ3n6gB/OnAh/VHS2TDSWi+/riuYPFH/aqxLw/KGEGV4
ub4o7mgxFyIRg3rEU51PsDMh8V3BKxjeP2W3WS4fWGN7bGZuf6n3aKZRUtgtR0SI
36JCLGWWWjGupKToE7p31rIcGiEpWOODkhyazqXL67W8S6V55NaNuaqceux+5+E8
e0qwrSqkww2BflZYSawa3VxhBa/4KmiZnygVol5YCYlAtvlM2B+v2WoJZtL7JHAM
7/NAq2gModL20whOtvFWuSyRrU43/gn/mwTv4nWAGHbQEmX0NVOtxH29xt1WPaEY
LVdTm2P8nx4ugDFws8mxfP/uFeyr75A20VEoUN3Cu+PhcQlfsqzBey1t/2FAbBn5
cC7MiwVYsS2TfVgyfAMAEwS74SZBfvJLve1q42ZhlAqsAFzntncouMIEojDnnI50
3MODf4j4Hw36PfHdJj90uCG+8hmoQVSGfW7Rh8M7gPCKLxoCJv2WrRUx7JoXcKSl
A5p6ScLgGo+r5gvJgmyFRJdcVfrZvgfkrqxvxbye899Fl3kCM+Dix7/AbyuiI/TB
p6+otwx5gGjmnQ8mTH4v1BDxoeuppXL6hcpUn563k9efezymt4Lw+BNg7H4RGQV7
/Dsr5onaqjwKcmX7gj1d3ckCuDzrbda3MQ/G9WOy9p41N2nVl5nQylylh8mC4h+B
0wVzAvIPQhcsGziKAUneVYMcr53GYaRA1gtNYo8E/EBPrXYF+c8nifUajzYqgNh9
//idypCHIfcLE8GAX8Pc7utG0tQ4+3EU4hCtuTZ47AF9KIvgXO8qX4+K7xXqklUM
mSEbm5qyBmiKYcsyP35vZMn3Q09UTLVKXo/S3+6pY+KRBiS8NcWZA72djwjVCVUB
MsCJyY6XxXR45YP+91/jzAz5KwGw9wePi3pAiwSbe2ACxG4ZGKzgfScwF+ttLCXo
UHjW+z00pZBD5Z6J2TowsdUSXtbDFk3wbvCefcda5/ZXrWmaawGY0Ya3SkmVDxKo
yAfv+IvywCMWmTcyV0+e2gs7Ypg/7wXdDze0x/exG4YEAPzfoI1ub+XMjNQZQbQ5
ZS2L/EIDxzUj0b/bbtZH4JlWqAOAxDj4EnhVRZTEFy12Vo857kFfvBqDrPpgSEVb
QtsSWeUk/Whdacjv6aunewHGvukYhp0u12juPQqssBwWm+TOSQ0cq8SdUnkJrOE/
MRetopLPEBz38tMEpiVQjnv/FBNWDyf74oC9P/Q1qc16nXC/VmOo++i4N65fcwob
xzOWS42Q2clmBXl8qfZ+E/M+TJ5XhMSeYbmfPPLrRv2S8lPBkXhv73B+PWAh9DJY
mQnoQ9bsQjI/Nj+NVEztrCRubVZ51LYB1oAqQYzhkaaWuzP5llGwam+w7uuAGeDk
fcGqhhLN8qVOha1fzHAtp3WGOrVCUkq3U2oe8Fjlw6xIQYW6OVJNyOXK3pH4LbC/
xBMKhpwxIQI1ScWE1GGzzTECf7J0S8vEh6QqC3m1PkOM8gro1TlRn51zeJMkou/v
N7p8/zb/ftWtdSYmgY1px/91ens56g1EVBTJ2aUnwVFfRYlYf0fF9HpDW2MfOUo+
sQL8gdobYIfRs7Wlzw/Qp2qqKwTcPPBp5ddLA300CULu6QyCGCDGmTV866CrLHUI
cQpLlLhhJyNJsE+g6N6O8nLPa0GrYTiiDUHEsaGMKs9ZKPtCTVbc1EApCMZbBgm8
Ru1debQcyUT3O2NmYkmTLWCOcIBrjnBQGoQnm8qrkxIeIVwSsGJTqOIOIEqBIzjR
nxDUalPyeerR0CyjcJ01KyM0HbTnnafFt+5aXzMEQbBd+xNyS81WLLDWIYzQMkcJ
ZfKuwGlUwn9yw034GrsiMtLgscjugkeETwIYsw0sKP3BKbLEC8gJQqv19/bR6V7G
+we+neL+ZlVjlaXAcLFcQW4vblEWB+9YQwi4Jchq/D+JB594JiaXWGLix5LW+HL/
DghSAb669ktxOp3IO83JwzhzkhODcVYVtUM13L4C2mCDS13flVfOazSYPmrGSyNC
8kHJH4xoxHWN6kbQKkSTPFVl194ztvYHty5Bkx6BSdgjW5c1NIkmsMlElHrb4BPT
s3FKI3dhFFmwcU/G4K+1P7mlRzCnSls8KlX2TY8wL58llAzyCZ5MMUJc8/IDLQhD
KYge+QdDP3CvgZBN9tirC7Q1woTUH+CeKgSku1I08k1fWWjmY+NLKCAMfL+II9Qc
Og1zf5IJfoSjLdyFX7n5As8qfFBSKhgeyCFJa9c3TpCN5+Iq3reG+VO4LRZnTYjL
UFx8ej62xCJow1almcVf4ZMcet1t6I4dXenbm1X0q74zvuJzxQNVpi8eVq5cD34t
LxYJ57iC58tzv5UUUfGdqocZgB5XKs+sIYGhcYhcBNMaOaRfIL81ftHv/Nr1DXGp
296FuEVztG8MTET4/MvFA+GxUsOconQ3ePnRTzKoE75CCtiX3BKqUBBIEySgYdo/
b4jScDNb8Ku5/IiGGVyoRQT/w/bdJEn1N/xiyH8gLdSHInfacyu76grKaJ/3HSyB
sJ/v1Vaflr/5YrtJUjvWcPL+kx9pvZg49E7D1w9G85hDX7lMDm3SRqXAsUflqFE/
qQjdStX3uP6Bg321KUDDis7btUJ3JK3dgKqWbL/NsfYN7AatUIeVBDcI+/0hPcSf
4lCgU5L1ZofVG74xw+QMLfnH2Jhx7pti9+1lIMCN9RZV4RCYX94MW/oUXgMLETDl
6NjRT/kvy9K4V1HCyaj2qYqyZmzOB9AvenpvPxzfOHwAtwJBey+fXNSQEA4QTabn
deVMILeecJNkvK7OY7Fc3rWRpqDhRkw1B/D1SkLKfwIMGMc/d+bBsh2J8TPPP7cq
djHFaTSuD/6eSFp53j8PYizybVootxXk4t4MO21ZxZWgIpUOjJkYcf2HkmVo0FPy
Ivxz8cf4IUjskLXN+O7UZSEgRQnv8oUQDZ/FBavTL98WgaM7TKJxUQCNER7PA+QG
bbP7PyGstUFUbAEIOYSm7WCZspgF3SOHNQF+58c7ZJqjbkiNtKG3qsbpjb8MV7rC
ef0I84zwtPnFUDBpc0+WlYtXbf7p8mKRt+LnAewEHuP6ut4njgC+Fo91/FHU2bMW
touuxT1tUgjlGIN88MSUl9GL0BJ3hGtepGEuysrVpgbUO8zsyWbloASXnrdO/h6e
uLKfw2jFxh2hv+jCfA29HT4EOT3V5GUC5P6PFCr4o7YQjxvUV8VpJJrutSloVY7y
PiMcToxLm1Pz3Bxdy185fPpwvhcEl8uMm0HqrQf7IuoVksRSAWiH2lbb0AQ8KwTg
EnJF2MMEU/PM2nO/qOhfRAZo14Qxw4HBt5OfNvZEBO86oqhQcOrO7UaYp8PYb4Xs
63ydlQSZe3nN/+Po4zsDWRitmalXLr0uEEPC1E8SrtrAvAGVXQlZjYB7Zz0AqNDg
A0qtkF1db+1mk25xN6ipOkdWTxK82Nc990FQMNevc88jLjaEgQy9J0jKHNPdWmFP
RUa3eaJkO2YJtNca9JznynAVh56nzLkzwIT+6NKtsfPTtDNZvVYijDeTfkz9M6vR
Q1wkE3Vrk2JT2gNOPy4G1Ub3cMEGUrP6CtbW5pRxwOSSlkKwUMVzsDrEmd1qsH1r
Fd9+OY+Va9rJ3cs80yMGNuTEq4mod97XX5ZRNmWS+Z0L3qMWB1Q6A4fq1RsfzaIU
CNzEqKobUZSmJ0LneNvps+eW51Z7CH3nmovQfi3s3ZNJz9EVFBKF7Iq2LLYqs7N8
eLgWv1TAdurYXsxFaA+g6CgLltobUnEH02aooc8T8dSnHu10TImloZFpYcCX8tbc
JuuKiSVFrt4n3VV3OBCceyxdAvN4p+bJYN3Z9WZlvlgfHX4rG9vXHjRrwuvLLdZy
8rDENFYLvS2Ih+eK0dCP7++0hmL8nUPVUNfydFRRWiQKoWvnkr0WCQTkGgGya098
1WWFwSU4b0P1xi3sOH2e+HDRUpahIbY2W6aK2yLs1i+YXVhW+0PWXdAq8QiDUUvB
6ojAqRcRQwqGWgAGw2QugzgKeV6oxUIhF9RMEzs0Xjr9wMKZw5Mp2GonTq1CHwS9
bdz7UqQBk+ZgOVkcIkmH1lLxZzehr/eFokpicopueKZoBij/DYKCfyRCt/XRE4J/
FLjfDGLLh0Lq5Xw26fkCLmHIGS1IJp6PHlRMO/TCY+R9l/ayYq0ytMqA9A9voNRt
m9+bBklM4jkTtATna8fZqnZxRMj+EdjZ/QbsCy+xIsZocwK+K5xgZY+A5EKMT1dS
2bu1doLCF7UNPOw5dt4BhYUMCTH3Okq5ImXOo4H4pr5Qe3DVG6QdXmYaghWuE0Q7
qJgerEOfeEXAnTn8gLAUDsPxec3pxL9BpHiu+3kTN1CDxPVKN2WMdGrPDIhj+Js+
+jvcHtGEIlYhn7/iPvnYE6ZX9icgAY8KAcuEBE3dV9NJCUO8wWQ7s+DnrE2+j1cF
Rq8wTuJ3bLmMrIevcgjpLC6qYHcZDc3Ns5qlV7PxvTqdHXwNeJEbw1sLMWRSIjw9
Tca6VI564mHDro7a06lXQPfkc81/HuBaHK8IOZBWYm864zJOQ/9ribIz3RtXzv2S
J9KbsRlODU/a6BXWPc3ezi516oqqrUSM3cOT3+to/RgYogAPfb/bloyHaCvEpvSf
3iblq62lCM+MlupIetjUgfL59962IzfJriJfVmAigTgZzCY+mxhC9vRZ98+bQhiy
Qgyaw3WPdW0MqJKaOwHS68nUpfv0CVEPYRFP0cDry3/gIYGNuMJte3Tgjng/hL5i
1EDoPn8Guc7PcQ6w2yh2DeTjFq/y6qD1suJvGLgiPN6H2TYtasiWhnXYDSYRsgd6
lkq3sLx2yA3lUCSWEwaoOghxDa1g/PjnfKJqSJBcjTHc55UMzcYAGngZRTWhIGa+
iplm9/gg++Yd7r5CXUSOu5RHzS10dYVBHcXeLZmoISFCHfIAmPNgP9tkgeu8KOD0
4Yz1VkZF+J5iUk6OH1nHClv3D37R+YUTXzfl91Mfbst/Bw4TzYgyXDlOVUlcczDw
8jMvYiWoaeEpTFvjlkvT269QptmUFe0zlmuisN7SxksOBMfWO47kr4GORLKrrNSu
yz3aY0ftSmxYZIdS3W09GzwVxAYVEOOiu+kDhRTtgQeuEPVRqTFsBDKBA1JCgMYj
Pb5r6tT7nwdOgp20u7juRyVt9O85yqdE1pEilHOt8h4RsQlreul9vZDxQ8lTFhho
KLnpGTdxhHCOmNje+KW7AvVOwhCxHqv8JKzjARFFTOPTEGUFzNeip0YpUvQQJEZt
sZBkMyurwVBIqI6FQTjFD6jhI8LozFVnOzAmFpb9pAK//R9uJaqKOsojg3W6jXNj
QTQYY2cr/l+nyBikGdxVlntksSRYKQ/oJtj4yZNbu6qWKLNajrYxZLphVrFKvAQG
DqTEUTRHvfHCHn4LSHqWoJs21B5g2Zmj/Gx3MlhxW7F6NcpqFHbiSiAn7jl4Qhyk
+Df+J/eX5IeItCZv/RHMhOMOxzcbYUjRhNkEajrQT2u93l+f1dujlmnxepgcrx1d
4O1RNPVG9g0/NM4ITdtt0r1fnpDV26HOEfxWn2vUNqPcOz0kDNNqf4wDw60Eux46
cy7ksr4YyAaVTHmx3mPbs6hKR/BIB4q5rDgL5FcrvbXkYOpjjewYmRgJCVHcahym
vGI18hRxd4WoUxujx+JGnBJAE/srbyMNp4ITkUPDwVOFJOIK/+X0PIFtKik0VPtc
30D1BqkG3YfffMwxXkA4w+ZhFvUamJb70p6TuoQccQI1pmBQ8IZZ/uHexm8xFgv8
giTAFDodMt/iXKUlz+Z0zAaia5SIiV3zUalZxdqQGuXKY3fWdNhSQEhYWyRAUSCJ
BsLQw/WDzchuljrmtVViXyaHRwO9r6aCCQ2Y3i5YcBETOu9oztmsDiouCulteM3f
rEkF5RRwFwwlTJggbFq71fuQE1U0cMDY4sX5RO77/6hDVB1vnY/3ggj9iJECemgH
Au23Nk5YSEIKKHowwcuDFQrq3Gl10vSTlGMTCzFY8Iz6B4DIchV+8L+Iq1/FlPX/
gKZtuu1jFeUMjwcHEgkQ+vHaKXqJeQueDcBLeGWzGd4rmJZJWWOn/GxdzIPDvqk7
FYxfq8LPn4d0FhdvBn6XXgqUKoitEbku2m0h7m0qohWGCm1c08fN9ZPTIijDMxHp
tUcH+c85ErIB3UCKW6ElviUDZ5ga7eGGQA1q1SU0KeG82N8HoZdIcNXGz3hqJCIB
sSksiTCOzJo6maHu6fl2bSfjZVUPAWxgHUoo/CgQ8mOrZLdatp5gyz0WG2vLmOA6
RKWS/BM3A9w7EvRfCoQbliGs7c59tORebjjtlXBpZG5e7FI+9i8ZCnu30kwyiQB4
tiLHaAy4AapzYCD2o/BcS8Rw6wBbNi6Z8OZ0UWIfMMfILE9nUZ3NZLaffWiY9KWc
CS5PklIxtqHbmVP4ouWJoD0bfXuGGJyEJzXn89B1W330k+vhSOOae8FXOab6ahvi
UKXd5YYGFq1NjiOhCG2t8ngpgR1hZPvAHs9xyIlF/wnBpHketCkuO8kPU42RetLt
TxA47kjdIDd4Ocm3FmAiW45FD+JNf7fdPwayUXspvC7a+njqw/GkStXNdIaxt5LX
ChIjBRNaihR8EuXQSuiJYRLF2xqgEf6y821z7VhJtwb9SrYahCLmuBlD9mMOo9El
WncNJuGysgG2ZvrlT8czy3y7+MDcx8i7K6GgeBoBGhlCz2tUNUttDRMxJcyFe4km
2A8JkMyx7pp90wA1TPGgbIy/AQxpohHt1jhZcpZ8QTOeH4TliQc+sMDT7TfkidV7
+uB2Sj+kAL5Hl+pGlaGD3QCWGXud7nuqSx2Ew/m34ZDWPwQCK72+NL7hQ5ag97Ck
HvigjfBCSdKSdyeNV+wXjcnPXEjlza+FCSKgcbXbR3tqV7YAhr8s6nrhqRWKt4wI
ZDUeJd8RyGcjZZicSOuAFiuhX0+q3ASMYNwXoFjuJUzIQWZb/MPeuIr0ttQ4RT+O
I2neKUeIPVqMvPB5oW/vMCZhHe4pIYZ4tBnjfIj9ZN1SGzDTU3T54ww9r5k54pMI
3b6DynPFvBRf5qyI/BcsqLpRwcAXpXvnYcl2iC5fkgB0xImxNCLoT4seDMfD+25z
MpislbxbqztyY7YSd0THsrngCa1rKkN+5h1HQcCqo/HE7bot0xoQuO6Dvwzy5QUt
xVPqXhz1SDQqwbmYRdrPJKie9P7tcxXfowOIn4skn3z6KUvI67NOYUTu+rDzXtQW
yrR8CjRz9Vf270SaJCzdh4YGb+raAyTRXYf49f57+qvfYVJDWoD8b1s2+8+tEFa/
ngBENyoEhVH9yWff//Qp739iMpRJDyda/26Y4bYvz24lQfVBAO+6DKGxspM2hr/o
9rQ5kNCJqdYnbfTynAuWgIDjydmDuTu54RYbKLcfXrlXqnrMxWyEK73gXe2OzD0v
McjViaUv08exEFzpkfEWnEqmp4YzmY2tu0TDFMDgiPUYMhdC8hMXXJEKuLSajUTN
BO0NUu2G+zJxdqzEX/Z+WgSKP2OJ6abPXa8hJLuwHJpPPobiXYNrDnW4nGpTtmzI
iQeGZ+X07xvlJXCRkqwfrPpdFOTJKZsEdQsFX2AYiHb2ZpR+xOcKo167QO9xfaZs
D+CiaNMH5B0H3ygO5JFPctsYCe4sZGRNAkRksaNxPhTBaaBItun543/16JPxo6fA
DM2YN40uv81BZrrPgKqy6/YhCVpRAWc3ijS+SqjxclX2SNWSORHAA5yuO+V2n3R1
DW6idfQi0EoaZj5RS/Yw0ISX+VJMOdj4ZjkBuc0EtWEBLqt7jnW5EmLAn0HmudD/
DdYylu6Rp7PoMZlaI17pA46WIlmL3qSrlTz4cXRna7hHrI0l1cysc9CPm/NyP5zW
nu8mpskOSmZHx6o30vG2D/FcIs/QtXWmAjmUg8rjMyddV9USZctGhuMdaOYLbFZo
XJZ1SLY+2oAziX6/YMpFTXmBx2Y8t1+Y5g4fFi5faPZILH7WLvEOi9jxTLSdxxEH
2Cou2IRkKgO3IFgu/+4hBZ80JoeH6YFo6gS7ckhB3RxShWQ55xmD+CErEf3Egggr
NyMZwkhpuTGOUJunftapG21mOwb2kzaUmaz4aUp5Hk4gbuZpxjBiKWZuDhfZJeCc
LzZtRNvCwemYZ7aWA+cy02aa0YFMYBACl84LN+ldY466WpUpC3WLL+Mi4AE1AMnq
p1q76iELpT7t/ksa64VgbJHgxied21Yjd8ibJjIZ1x+xPZbYSLx0cZFnvdyzP94c
ZnlkmlzzSdhw4MOe3z4V6j/OjNPLovFO7/SxEubxTSzA+3fo6uLfqX1na+bgzsHq
9N97OIpCeLjW0ZKp76mY/Wm8q/V2MEoL+vMJc+oKUeDv5b/rR8XfAfELpr2NsU2j
2Sry17qD9A9aOw4pKjkJiEfC1HZlxRq3Yn8Bn5p1WM/+d0C++OvAnv25a5BGy2y8
tPEACHbf/GMd5/kNcNweRy01ZM2Y8SUZL93GfDPNJofGmzVYw9GnMADdHIpLHzrT
2xpWOkEEQUKryaX8dXbcf+w73mDxoq6ZIj/7Y+pv/6TTI8FngXyX/F4sVQi35tZF
c0c9CdSap+RZlu1zIcgJQr1Z9AXMBnxPZruNfB91xbLAJN2Bdaesqix13G1K86dd
SngGrXAxDisuxKW+YarlLwBNjQVyn1VHTidL5DPnrYCXRUGXVuZbpkQ/2+EwlUOV
5Tp27s4sVXvOdajsn9indj31bc/O50pM0QlfNja/3jB+SepUdAmJRe4O8HUdbxLe
OZHyCFoQ5ocfpHjQN2P1QjKEzfZB36FM9/ueccdE9z9y69D+37vMqHglZhaViLIp
NYphixlCN8bbjz8M2TBfhuIuwSyiQSLRneYDoinDI4RNixDFrlra0vvqGTsVn65H
yZjgs4I0NAkN6c4pCj24TR5kDtB0DcgXezR6C/+datrmgtYUDQ5c6WeGdc8uRMle
DYExbZmUZ9F00b+CBAPpXoj90FAbyF7D+3Cp2oWMKPh7wXWgFbBABIpjOcBsNXNL
9R2kQcLG/FFzf4i8A0DUPYad5GZqyUIo4ptiXXH/NgpsZhOHG6oHTiAD3HLpn/mA
ime47O2fK00GOvkuJmigYh/jcfeWmC9bQC0/mpt/Gt8uw/TD3c+8pZ4vVwOGLTnK
tTLD8mQTUrC8eCA1nKOjW3BCbBiG7UqVcJXo09u+CJI1hLIqLvX/ygW8OAxOXg0q
7x9agKG5U14HCLDri0gZF26mQgn/P8hQmEguEkw5n+b6jJ4560EUObxfsFCT30mH
j/vlSoUubpozw0xTJTu1c6NNDeD9X73VcOLTza1SE/7YYzsrgZfGiTwEXiUaqIWA
IbYrjh5kSI8kIow2hVVI5wabKChPssyzRr/eAzVmHDN6wuUvS3dwnKbxHq+9nrZM
qj8zlbJN9BzjH0NfEb5pQqM6UThvPTSJl1eN5VS1agTFQLm9Lfag1GaCxEnLNLg2
k9gxU34v0h5fVy1AFQdKCSLmjCRSdlcvYhxfJ20KxWl1IwmHKbnUFzmdONX1Qsss
unTYWKmG7/4N9hrDQM+Mvom9LLUSzlsb0MsydNJvbP7z+wVOFD7CVxBVTunLn0Lf
MVHZWh+0oAqNoj+IVO18tSLVzPmUhy70sheEU7jQRRMBGb1XYbf+Nwn2xMi7WgI/
cXLz7LtX4WLMfGO9QOmwzhgP1qQNvIW8NdciJIU/oAN/hCOj8ruMP3epOSYVHC38
tiVgivVpUG2xptbk5p2A2wyS/D+idOR2R0KwBNbB2Y20i+m+AHKmXtg7zkOAIN44
+y7vqfrgQej9oa9DWdE0IX2lU6ztDEOouT5QlG4Re3jKp86P64Ef/4WG/x3VkiOT
Vsx3O0PcudQvsSX7YQYhuCu3aZM3iNwHBvpKstzL7gKiHTa5p5y0Ov9lsj0zFjBb
gFPsv5Xvklptt34fJBJE4JG/2+Nyw8dqb3EZxPahFYW3lTIGV4DZjazJG7LCVIaf
yCrMqYOfoWMMnRG1osykzar6a/Oz6u6c5kMOvAXic2Z1UE+H7La6DAVCbE04ZB8I
j+A4BBB4jj7ZZtPOoNe+um+Vz1xAfwpqYjwPIsifqxP74Hi7Af+HchSdrOHFxGrP
qWirc8OjiCkwog+5RTiBwPGEN5CVUqe6wUc2dhq2ijQ8KS2LVJD9oJuuwY492VBX
cCW575YuSlqY6ekbQal33993WLNusIOqWNOk9bszUF29nWbztZY2CY8f3XTK7eeW
Jc7VcG/e7e9BfIiRaBfvSuoCdDkIQGtC9GBG+QVEYsAzE9XJuUzK4+lDm5n1ZjXa
HsXxH+yy+Q1I3qAcvyRox41iX0Rq/lbK/jBFcaQaNc0IFqpJZPKrVwq9yJrAVq1Z
jjb0vxLH0s1q0Oa0Ps3UiIuqaJRYzPUZk/Mypq0hnuveiCLjXAktmUNUW6a2a9+p
h9GGV9ljepuSSbbjUC6n/67bK23glt36rAm6IadTBRKr/9wW2jNV1E2ZtSdWhAik
q3ixKH0HANH0OyVaEsQRggb3zWx+A2J0Ajvkpcdp5AdsjS2SjHB9vKJJCMxLiE2s
QlQ0eqzN/CwU+h60jtP4PWxUaacKaHqfGOEYc+CljDm9NhQGNvmo4Clymqlf+Yn1
uR/ehF3AvPpDO6WAvpVHP1KaAIgwbKSkiekBWePR81Crgh0UEuYj+dHLIcpENQH1
RWL7NJYPQFra3Om4uEjBcujkFnvChkzs2m7Br1KhvX5IkwyY1m3PQpk3plLn5uY8
a0vXhwKw0G5CJfSVq/NBZ1zf3O7V1B1QBaG516UZxtEeYncmX0mLcoNRj+bc2Nvu
oJgxVw16h5Bk+j6G8qqfGH1hIwLak4Of43TslTGreXzXDpIMsc7qtrlodWK08BZ4
LXXnssasewqRFB/J33ZZeROtpggmTJ4IXE8K8o+uMG1OYYbblZw4t6GGndlJ94/6
6x3FO/DAGPkbvP61OzdjyFX/M1m5tXWncyrUBk+/56ix/f/oVRIE21ZxxkyxoA0q
Tiy8eqYf0rdTqNjRDNih8PdGy/J90+TxvPGfubLPKSBMP5JYr2DzRxnNNzuzOmfE
nMQ3qyeNNDOtSSostxNFHN9PQe+A3kUzvr+zwCIKncyeN1DmHtpmYZQohLaOXFrB
6w+cGdkAPvGHt1rII55WqaWD2H8iEU9eyPCRcnQN/Fq4R6wZhB8ekhhcHmfklyRf
XVG0tvt7FUumnjgnFnCAL689CZaVqUG4ApcVVN7AhiV86yUxRB3GzJsj8Srh0/P0
wQI8JDA8ECLvfOhg9y0hzpNzQVVN0F12x3t6OO9vnZsVo2XZwYj+JvC6cjCdZsyQ
DkcGYKE0aDrH/OyYf2gC2obDbvUsWTqXJVP1vAA9PtvjKWYHnEIc/TUSq6XYkGmb
8HiGoSRkDLxYkIhikX2C3lHsWZskpBKO7OryBGN8OdME4m2SKfwWghxE60t9cV6M
cl7LPKbp4rq9GTj4Y9O/vod/eNkzWBDphGyGUUOWVVhJ9jpQ6EL5YcW2QTiKGFPH
j99Iy3mWtCB0qSQc5ynk4kfxzrxYG6LEeQ1P2OnJ80FsxJVcdixhDSybi9Nw7Sfc
1K50Jc/1RHURWpBHbkspHQHJjw8V6eVwtAa0emNU54h75CqNou0fHh7yurATlSyl
J+iFiv3983fqeulzX3sn6Eqtc39JOu56VRKUFU0U5rswD3XvW3UeDzZeD35krItz
lsMrU4SJVoxIh7KA8mru8jHuupbOj9XHZ6Yvy1Rn2Wdu5vI7D0oMaM2pLCPG30gH
60+FhP2Xw3q++3ZQk7PJreeMednwVM8RHtymdH4QUmguikANDDPZ1J6WoN1VVGND
SpnacrCvPvZAT9mqyDnvrlWEZv2G6CUs6k2FnRoPPek4E6exDRsd0DVRyTrZpoMq
DDfBS+tbyN3I7Yh0Nnh8jPUDtCABOS/+M9scKyIMWfXAXvT3cslt1bAqts1Y9437
82rHXiXrRH75t1jpJOyHwmFyc1gwAmabGLji0zrHZZtpCpU1CJS6O0wiAcQ1oFKa
7QDwApt/zSh4IzZXnQqR0fmkpaBjViHrvmkMAxmPud4FzKA9LB03KpY8obDOy8DK
NFCf2IadmAm8qLQLDxztFrMlxpyV4Cyci+jAxwwZ5qazhaQlHGtdQBmEQ64nO/tR
IjqogjGrCScIOVDNxc3JT0oUFrs7DHumNmXbKE0xprLoXH+4SjSZQvGYEk1QP0ZE
Ej3hreHXIsHxeWZ0k6WEGjA5Hh8Wwvbdiz0XOuueoUn8rGjyM5AnfCdRASXcP/BL
5ldurDAzghIRdinLCrQoEgS5osrahrwBuZ1NiJiEpZ9MT3wEjNfnI0NXdLWsc88T
ioThn4wXE8X5uxouADEL3Z9GePjqrgGY2qUwo66UgJFM106Kqh5kGyahSwUm6L7j
rovnLlWDJuN9bvOPf+o5YRDIbT+Zvyjxy1aYNyZnf//+mpkiFtiYU5FDBEKPcoms
tge1LbEvRmNO8Aca+kdJLChfWWQG50VQjAQrGn7N5IsDs7GlJ1x/kFyo1rmOSDCI
fevpouNJ+B4TE1bbsuVy87sZyQMg39xvqzxdcc3KZVxVrdHMaD48rapy9wy9elVt
Kk7Oq6WlXAs4Vy8rlw0+mF/f5PnYOAz6CBMtTRjKcwm66ecRjlgUZWtHzMNFxJ/U
sEi8aa6tHSoxLiWl22+WeviKMeMEUgvfcv8qtQO/990HrH0TOGZ1FSOYGyZwkYkg
mPwHmKavWmNTiNVJN6eVT4F3BGri75VET1Eq8u70tHozacoTfZ8KVLYiDEaeQ7+D
B5OlIo3onCD2fCvpQmSDQt31Jsr/WeuZ7kYKawPqtu8M8oIy9pfHPSYkg16n1Qzj
rBNdJ4GPRZ29I79ppGKtQz1DOMYz4fkRNrmsstUqIqbnb+nwY9FFH1t8mFAoQih1
NCEiOeI0KWPuQNjTq3X84J0zZz5M5zvm9vORYhtMyZ0vq9bef8E1lu61SW1D2erI
ofxPXHC37uTAgjGTvnnkzVk0lY9TpUK98LHp+yoq/udZyjrU2orvbrq02k8zgu3u
WCNNB2UFzk6xrJg7SaTIa6SjLm8pSI5V2/EqluXJfokwIKL97J3b7NPSCVbTFzQx
Nfvs0lYB9s2g/p9pe2jHBBypQYUgUQUWq20d4CiIhdRwgZWW6SB2jzzCZagT4hUV
kmiNvfGqK6HLp2vYcQ4H8Z9Rhz5CbYVfdCep4WvktCXJsloQw8xOvQ8OhePi4YVV
5A60Ph4vR+CRfRC40rFg1GR+2FeMpkElHYd9YlBVpwly4NGDbhbiMcwHIaJWUfG6
3B8uuANMe+F/5PpMXOiXfN8vOmwVUJW7xRQaHOl89BhT3N4/lrkuxHmNBbZzwBzE
2Yer8bXPp1hskOwZHtxIMoYQSnxqctapwMgiw8jyvTjIytQCd98l19IzjKonVO22
MWR+qs6AbrKHqVoYlGuFGy0MSBUXRDF1pZrwUjfEUGrX3x4JIOTZkSfHgvGpqJ3x
d8atee2cDvBiX4dSrE6P2cRdtNFg+memOkIAyMBRnczKMopJaxF5wn/Yxn68uwZu
jxE/vsXdqYe7wldY1S4Cp4E8bO6adK4CmFiZZcKQPprk10OEuwa3wyPrkObNI4UD
9OVaPCuH5wWwkup8Ymhj0RdTd5epC/NzJQ2UqxplfBR2HN3iVxso9QvHVpqu2n3T
Co/zA1WxwL63vyLrTZPOOGlZH7Bla4uz/nGGDvLp/OycBI0bYNyYWWvcn6aGNuOK
GGuu/WD5NclcSGZAEf1HL4pkjJpSob4NE+oFDi7qU7T8gcDB3WPTrTCKXG4RNo2x
sqkVXiUC7KQu5W+iN2mFAZRnZcQ08Rpf+blwKWR9u9HljlTxi/b00SZeubXjBQH2
mYQ/kkwa/HCKQYr7UZbIH8B0ZzeNZw1uQuwyBmUzbn2esMc+TKeyxw/upb/NydqL
iKUZ5cTBJUv1GohsdMN3RQd4g+bEcOwniJYYlHNbQTdqVt7Mgz4t1S2XvmmMLIBq
bGB9NIRRIUqa1bB7kyqER6jdAhuVHzDgJ682YXn6Fqok4HyziEDp3yufjmPV+xPm
qbcb+D/2fgO695dHd23a8E3ygPwY/ZoUgfKv+UN8GENdA9hYhTlu4UJk44pmV66m
xfrKsgo5DnDBCg+J8kAaUOZQRxIpNQzp+wMrUth9psEP8IYaLXhKQYaxmDdVv3Xs
VbfmL3WrIOysA7Xarbbzrn0xLk0TMqv6UxVOItmcIIsCeT9ysYGIkqCK/xGMY5B8
Hqzk4IiBZkMvRn9qpjAIL+lPKrA1fPw13sP7Jj5bhPTuKDVlE4PCZSD9Sc2VS+Oe
Plrd7M7u882vS1un3YnyHRoWODgHo2Ajf7vrN5p68NQd3c2+WdqYPWfN9SrjJRzV
QHbZdsCGJY1qTDpyX60JSGtUHLpBrV6/FqWAwmGmJ6pZuqfzL2u/jp7Qj9lD4RXi
XxfnQ7PAeyXVzOsRd5/xmYUhLBhuTuheKECzdiF2na9cEnJf/hTpZgbCHyK08wBN
yijORDQ8C88DPBK7Bnz5sXtu8EZKONjM286hhgxEo56shlMXWhCIgpk3mvavlrqL
sB//JSg9th1frZj8XbLTm9gcU90o62ZbebEpyXDvt32n3v+J/0pwXxASyrgQY9Ak
iylwrqwlTAXRslPRzE2WjsJ9VDwmWpKP1bR8GfnwJpTQHdO2EUtfzvgpP3hJyWKv
+hRxHiLq2MU4SO0xsOI30PAx/hCDRs0qwHMH0BoFRD+OLBfWj/zM3WM/ksmfI+fU
nqvBLjTJIUt880OEz8QOBx+HOiOnPexKuyaPcE/xZJh8ULMJFFXwL+8rTeqvol2L
JM/88hrffpndaRjNn3ES8q81bWrogs8hHGGLCwlSPKmOwlbRpelDckHdlULUUP70
mYwYKTVJ0iMX5zWqasWnfbdj7QbiU5I0j1xzY/iwLfanv6XX4hCLbU4M33mVnV5W
U/FBfItVBi0PkIAg51qjKNjjWUDnhiT/qxRrxXsVP6ljImcV0GOBdq3ucWBYK1LK
Ot1hc00Co+nkeY3OnFmDuVyMhZOxJJY4sCfadixAc8GuZMfYzzsSy+hSCqFHPDIS
+WFuH5h5uDZ8zzzmrEPUVh9EWLwycVY51EQ4IUUxnmfZMuJNjpnXv5h26BbQ6euz
63G+plNVXjQxg1ZFxYZJQb85B3PHnMCKZo/aKQJxs+ICgSzWH+950rcbZQ8ocD1j
19eEyrjtCunMxT179j6QUmMtypDrNnLX8XFA/OHVl8w+cai/GdK89gnvQIE4Vc+m
ytY4w1SDOUdhy7wxrH/Fbb4Fyjuhh0gYcVfsAOAGnayym+lSc1bePxdnSZXdk8cH
aZp1kUeDCommB5Q9fIXbx9KGbcSy7uY71+Bb1VOaEaJyzcMrbVU4jYjHRTiNf8bv
7cjMnX2He/JNF851vDmwn+n65hdk5obkT+2bGhXrk3fG6VMYwfqYXnZNi2/eKIf0
7yHFE4vSPLdsxY/CxABmeK1vKTrFERa9OFvr7qWMMa+nx28o/S68TJGvgQ4iQf2J
XuvT88IP85roVPOYHoxhnGs3fnT+2+BwSjhYIzSFTVvRxIwg/+H49faKUqW5Da6L
Ip5+CqOQGC67TwFjJIBPZ0Z87TVBzV37ly2AE023C9lApBa0vWaW5h6GX7wJtxp9
oWT0QMFnoSqaRi7qBHp/JYu0YzA5KADPOtXrPUQmmNa3ix6DCnFU4Fq2y63E8t1Q
pbqrKvRiCk51MAktXDMVoh837zSbyZS7B9MjdDHSs/hHtbdjSavPn/VL6ssY0ZFh
opvI0K9Sa7ZK4KatQw24xW3nyNH459PqlYkiNeje4EzZ2IqK6GqEweoJp7yHibsd
hWW/yqTAHGqDtOZnCA4ITYpa1F6jkoTjj1QSLsOKUtu/bbQCtCmjb7w0ByS6HgWS
0VTzYlg8FhT7Ix5Eih7+omTeIGmA+8GyaFBqmk3lsAqK2vxs2Oe+G/mBJZ/m25EU
GoAZAZ7be/1Zr0X4o/xaoT6h/OvDR5BEmMvVyoDGQhAKpXNib3nyMNzi6r0M65el
sYNvryHfU5qeIOFjBfG5eSoruNgr161vVO+UWL5h4+yhBfeN8Bqu/i7SLDY4X523
4YhUgihHzcodzJ4bzUgKjT8k0wwYFhcWsADFhOLqGnNuB8Tk6KRC+Dk1OYPekjHA
LeRAIetVe0CF/tO/GjmPYY89UL4hHHJe9PoN5nxoohfH8zQQkkkS3XUMZ85TLYh6
/FXApnO/FKt2iy941/4YBVG7MhCyHcJRWCejui1DEmq3ws+ukoGo9qip97Fg362C
58Lpm8S0zbAAB5YeZOLfPThNgWaSykw9f7ISrAcVa4oPZXPDt05OKFMi3huhNkIZ
26O6jScc1GlQLAGJYHI5wSP1O+TzqONE/gJfXtLXDBVzpDN5jAHOMsD2L/dKLLDq
m9M0TnWmnGP8An2DJNLvPe3fNCFukLM8HVJuGJ1OpMXj2ZmAgfWvX1Nvl07ABeyn
OI1YxzvpyqrZZqTnhu7qaikxNpiDV5cXx+deULCc4WE4fUu88bWDdq8RsLYlM+tc
iGBvKaO53jmdQw3ARCozKHBzs4CX9BZP4ldbk+PZEShKPZL9tDm2YStpSbBqiOT1
5y2Eh6zUr9+DcOu/EESN9rdq/uTUZlS5dYQ6Do/voouI9ZfQjznLiyFqX8XdymIo
pyWFuPHjmrAbD6yF4HWHjblhGf38x+1YLod6h+3GIKh8nD9Ui6mWNlPVD2+AZJuV
o0kMaKCsqxLdpnOLjHBGQPLE3qObumP/G0wEWtCPfrj9ANYNB/Bj3a2ASPOhXwBS
8ehIJNKZfYu5711CbAYMyZi/sre8VSo2yQHZjgom8lxICXe0VCzhNWnYQk8PNo6f
Z6wbd+WNcXj9Ujzlfn4cj+Tz9vW4yf6G2r4JFV/wU8GQWhcApBNG7/Rf1aLrLKuE
8pzVSTljti4VyJ0teipBOayOiIyZ7ZcVXjMlPNsdCDnT/71Hp0FwcuZFqngybrDM
jGJGP3pdxzGPdG70a3dPG0ZUtF7DAQ4hse/kgjQedfeqFipArb22u8n42FPp+WNp
sVevya1VG42zgZ4aAwkY1RLfIDSpA1mEivY7jECE5pEjp6WuvYclCym8Vev6jCnr
3itYTwzVll7q6D3+APT91CXgQrsdq8AmLacMHMDQxMrJWkoowAvGQ81F0k84Z+Ht
ualK5Ot91/ggxRjXxlWGIWzFBs8e3fSG2L2C2tFt19rBR7gQ/nXNqDN5zZIkiDQo
5iwQ8Uhery55wq75uIhhTSPIvnGyCdzWMmyiHotGO4gyG8fBB9LpIZGUz+j95Vur
vl2Oatp8KAhobs1BethoW2v60NmMY0VkRYl+5EvpNyQ8MemTkasgHgSdGH3w1hnT
Y5YdVFLrWevno93Wd/9S5UwMn/LuPZ2n6PtTpE9tOaTCOQBDN/TZ3AFCbNmJiyBK
gInw2357EBkpdQirFYgDDpaca3VdE+G70CQrHq5F85ACtCSeCpYMKHwdoESzxWgz
M3RqsHMQBMwUOft9OzYmxjDVpKXOJB4YQWE87LhtMlh5tLH6+VAlLoQKfmwwq7Ny
IUJT9ZoKXVayz1Y4tABrnSQH/l7njoAfWFeX1sy/B44jyl5Vd9M2IexZ3P4nK9U0
MFj0jC/Wln7zTAK9Prr6yYoefqKLs3Y2z94sW60i/R/+z3JZ3flw52t84P4so0B9
QbihoPabCBtBPgHhakBfoi8hUJ7UPPVwb2v1QkY1GaEDAAN7xVT0AAnefXHVjbry
ixxomQdAlsKOOb3Adzf4tcuY2MwE3KUDVjVUSUCdjOAwqt0PVP53yt4WzdbASeuD
9vTl0qFacbACCUc3Mf5+RKZErK9lPV1pZe/cc3Bnb5qkNGlM1QaoDDzBtv31Lsa5
h/wSvWi7M4UNFE8ExvRq34XpIXH4ZyXB1wpYKu8QF7VuUTz+KFWliMVu79Lh9CDc
PlBgEYv2GXqhkEtDzJBt7DvtAjULKpPLuiW4o8oHjtUo0nsTHvABaGaKVBpWOGCA
sdnH/B99EZS7+y3plbAQsqSM4S59jjT1yOwZ6yj03Q7lhqRZxblNeT/DPqZ0D26t
a7/m1bmIMmxDIpEq37H2GzuInLZElR/huloxMmHktA6kIuYWRRXKLB+k2mThyZm3
n8hP/p4cMTgDNFoevtbpDbePIhD9K/QXCH03DC3KmBso6OvGfGsZk5Q6GNnLGHeI
ovzXk2pRgLzWzj1LOsKZIlJG6Q+HiGZsONyZDGwQgBkllRc0hh86JpQPe9J1l2nq
QO0pQU2ffmBIr4Wl1MJysRX6E0wMSSrN2EPJB5m9ek6G6HiRGskKnnFFzJtLNO7A
koX67dqDxNE5tyGiNkUFOWskUohxlAFgOdwBGqmC9Kwob9i7IrZwgrFoRbg3cahg
io4m2W5Vw6YAdjjyNXO/7ijMgfTDS2j57ROrw9xsHNiDvizLLZGmcJ05juIOHkuh
aFHtoed5lXD2nMIq4vg1q9YzqXMONlwXZWE20Netd1YIXkrxNg9kIK2LfvI2CQlD
Pz+q8EJZZ6iBrystV/p4XK2dW1Rnazg17LCcsJEPpUHvVB9pRFn9uH9x9BxRNq+g
7K2NFKP4FVBlPJuLQT6aKn6m2vzn/lX0c2pS/5JVzsR/s5HW8WrHbe65BTSdf5gv
aSpmbtt0pu47nQ0Oe6heDOv3S6Is1Xu8eTja7qboBMl/RcxDPRvZYxyii1fKZH9M
rqoa/+ojK4gH9k1lkVceWZZdg8W7/ICrj8ouC1xpw3vkITZ/vZY2PVjJeqNvJ+jT
YqBC+SgLYxPTh/w9ZHya3usXTJRje96iED4gN+QMQLlub4iWj7XBU3iXWv32KE8v
HvenlWQYfScEeO0TVwI3UW+S9Z7Kg2f3GrITMluri/OZ6LFeKYAhBY8HHAUZtQlw
tWaNNCmsunQ3sUh+XocIhZQKTWl94iXahU/fp6c/SfrmX54nNCLAkGBVdVHT0WP9
/cyLZuxDEJpqcesteUpFD3G9En8LXB0Vkq9p83s2e2p/See0aDH+OK2SnUerJfZ4
pALvJqAlrRNTGdzPG4R7dz0aso6ODm5M2Sgda/fr37HLlfyXSCOodc+Y56/m4RRf
QRRLB1WeRVpL3FGjMTQmQXa+PkEq/c+t4IQWH9GRL5qqTf8WlPF5H/QADDB2rc2z
+XsWwvm+TlxmIYAyOIACjCO5UaZMn1aoLH7TsUSTS+819xaQ9xsLrJ5ckuhNZomT
7V3Fvt/0AX7zLgCUaj279Pwnn2OMiRKhurcuOVt5FG+7DFBvCKr+CztPv3NR3Llx
+xUaZZBISOIP0A7pkDW5q+yeeeRvoleE0XDLHVh6+ne3UpU7j2aJAG6Z2niey3If
uXg498cOz5YygaHOQwIbgjqxy6GNaxEgSP/bHJsafQcU9+I/esJ7Fgb/qNeUPMLn
cS/0e/flAOeSqyvAxTyWljhBbDfO0I1kDNNX2pCs9oGgH3n5nluIcuKGhf1SVfXQ
sFtCFYKdcZhHkOY0mJx3z/VjGXSz/BByQulB/NgttNxXobaSWnC9nlKjyiOPBYIM
nz+7zD23slqAnXp+HoxgLoPEZ2pgZOWbIjxs8eIpAgVjJkgfUjOjS+tSjAgE2F+G
3z1rzjWO2UBc2QYVdF7HOhHZQBpG4lUOknOVU4qJV9akHKV/NRsJVrwmRXo6GULA
wQcQYATH9krZUKafixvgTnUPI3tZfkgW6B1oBJKjBu53XAmJn2R7Vbn3leF7jz9f
rtxU7zjuLNEQwOr89FQH3NOwj+NUj0hxPFoolbysAM6rg9Vz9NLzu13W+aAGSNh2
CgScciVyo7rwqQ3bpBrODTKkKvz6ZjRPNhAc9rj/bcy/vDTAl9DB+hRAV6sDf8SM
xos5YruZNcIt3zlmVwhyTc7XUhULNeDRMid3z9clEHEdC0Pe2IeOuIT6G0Fq5yeq
6L/3c1oIgRjb225H+3ffoJv1oq39oxhgvsGJry893u50N0s9dI5E74u0XJHKciR3
zCoDFYYdLoP3qt/JVvWmSdR6ajrtHWf3ZH7vtqdRtsS5Ak6/O9QijGP0An78yyGi
4tcj73jile4hLi4/bL/nwIY6gpGPwC6J7bi/p+tuoRfM9E3jA+eT/0HbThXsrB2N
3dpBKF6tPudDM5GGPVSDEifZvRrUVPeQVOMoY0ufeolzXx8+n2+Ne+81kNXy/LZB
6qNgmYqk0ubHVZVJhNHdfH5juAdJ+Xe/XaqF1xfX7QZP/SPFn4BtFKpPhlv9y/NR
W+ZtgTSDItby1bk1SfgHR++TGOqCzYmmj7mgSpHdi4FIOCSTFtqGa7vysX8hBaFH
vtI3FeC9FEQgsRgyK7GMpqL8kcuIlPFt+kwrkh5QxyDPq83dGuft0IZWWUUT8mbY
aIZ9tm3BsLrxsQWqZg1m7mR+UQtSjLYziqRsMOERYhVzWAr+pJ+RAIcSe6t9vnDB
VlgdhHxxI9vxXFhuqUH3J9Ra6EbS/FBRRAkdUoY24XX0uKREHES14iUCStMXaGOR
ark6vc4LMi9CKLFCb5Zs8JXckl92X2AEQOs5W7eYtwPd19hdL3vynSHnS3ISv3z6
ixaxNjNujqIKf2KdC0+O2hIRGPkagx7QecRey6QOdMEgJIhA9B0rki/ZSdvYyUmg
y97gLda/V3QZbcgVJke1dNSL2Dwc0YEbngcsTDTvi4qjUrgXycdYsKXPBa8Bzeae
YDgKiJbEZdJ83uVIXh/vKuDvrUa4eKTprBpq1W12tdNZpOmD3xtKWp6ypFYy4a/v
BePFaX7MmiLeGSDLjTQXejqjTKS4M7tvkQwggIZehJ0wdsF/omB6lNxi2YdpjMED
OXADAwO5iP3JkaNQ1rH/dPmwDfMoJHfGt96NCa9QZwBQQRk1wzBosJwUTb3dasvX
dxuUAz3/I/xL4SaEOP37ZVN9VB3fOJu0G+PasbTvhP7wpTvU/WKbEQ1vcGEQ+5Dg
4TfwdQa/KgSD0tnm4CIWrys86f10ziuBxT7qYle2lwq+MgLsTUhawJJ6tM4eQm8C
z3H6hTrNPMtGPXNxri49IL3VZ03bNleyR3cx/8X2ivV2SVSNElmki5GIUFnixms/
YsCkfH5jYeY4pb8/v4FdalElXkbtkuV9HokO3EQjdoCG+8db9rn00JYHV8BlCB6g
ZJF9wgpl+YNFK0zsrxfsHG2RwTGdDVu6PDXDylFL8Y2jyaVDK9T3+WPRtsRap4/f
lr6PiY56JGcLU8ZwnW7GsbTEiGlxImTg6S+oqrOHYWTvwgDwkUmDSzJkLrpJDUcJ
W7byVEFvdwsZGma2J6qs4rkhxAqss21pDy5fRHLQXQE1tdPYhpZbglZ0YvGpzPTw
WFcAMOa6cQhNCl2UlSF5jFbZehDaCAzeTvfNLN00eKUEEGIpw7vXrykp6SMjCTjI
3zuBmtujfVsfyt7PiCB8rygt6WSpxIjyBs0R3I+ti44De8kQ3YYPhUFuVg36E6Hz
1iWl4aAQAy3rtO6EPMvSKCfUond6zPzXRXNydVxXp/CUc7DacoWd1SUNJjG7xoVu
/9T6rKu0sS7AgB9sWod/3aD8+NxcjAy80OptYfH3pGZDyUJHIov6Cj+dym+Qza5f
jFdlUQerIv6yw4PwsDkGg9mb9gxP4ihx6gX7ifDk23i+MB6WTDNq4w9I82+g2CRm
9ZOpj66U7f/+BusZvRaxRrhV/mXH/XuT6cDDyQF649MnigtiW7+8XQo/6v3M5Db6
c5UgteiwbX/shkP0VdM4MNX8HmK1CEa58yKYtVfSoiLsNaGGv9K5MbJSuRgaP14q
pno+hcj4jU2OxjxkU66KTwujKXdticy7Pk3svzSdZFYJ9I2e2lTm0WH0SBG/07gr
jTAX3RmE2tVNVzLzqs2N16JlsyYo/vK7/Ftgruo7WMbJU0boq0nKz9mMZj92ebN7
QzIHHqeTezTK2f0IZqRkWCB/Qxu5EPpOre8x7i0M5vuJwo17nVU3B+Iiaq+DiITY
xV1jDG8i7C2ppWH7Is4COn4KhwkRr7mTRYy88Ds3PjRIm2SpC55m5QIucX9DgtVX
MIVUHSDQ3ABuaP9Cu5GQ3Bv8iGJ9J89pxJ2NcvwrclpG0RcA0I9pO2fN9vckqB+R
OscvlrTEWN8L3JTc9mjhob5pfDSQrfQm6tylNpMU8DjjKtzpQc/ysYfkSHbJoqN2
R/UJz34O3vscRwaZ/XdvtX1QZt/gUsUU9TL0YVaN9vv3uBRoWT2N8ecKJaW+DoP/
z9+YIcnPUky7Hr4+1sBSqLbC/1PooKqgDryplcACv0gwkA+yyRi1zuaSTGWqEXiE
wZEiRKL6JqLsGmlDQImKdXIDus1g9DBEWYnR3LUDxwjQVoqpRhSsvHhD/blS6gnJ
m2hSFEEZI/QtEtPHEikAoVoDB/jdMTH9tgmCfg6M1Mb/sp61FzBEeTIXQ5o9/qu7
n1wWjB/xFRlwiH0Gf1Ek4D+NzTHaWNJ5bahvqmQojb6bBuMAVkW9kDOD4EVjx2Dn
vJSZ2jKlWRuCZ8yauOnf4RhOE3ZpRthZZpekhz3IzDmFzqH/zrHE9rQXyc8trhdV
cS1r6k8ulElRJogN/DKBeoATBgHyIQiISj9y/a1jcI5Fm8pfYmCyY/1KTH0jF3JX
5GbblTSNKb7E3GRZXwjeohamoLWYq4O90YlOvFCLoJPsgndpcWq57df/gDHan+3E
WakxGQA6MBFcvETa4qvHAyymNX+CicoEOyVb+yd3QY0SmKlWGIQbxyLhLKMIRQgr
GgDoamSJ3LTKpW8r6aSHdmmfTbXAFBRddNHqFzX0GQyF+leBbRI3OcQiwOkr3jvb
0rUu1b5sBVNANKv4TwfwSmrfI2NEh8HTm6dyBvS8GAa+Vo9uFpmczh74zGFM0XzA
0D4LwvtvRpts3Cv2T9j4OJEe0Q+8asoJ2lNKdXDD76NA6uKSHXa6CItNI0DJ5hWN
PZh+XQPrpI0cYOyr8whjcf22qBdUxBn5MMs2Mt9r8rG3EI4OLj1w5njoxm+ZK//h
K+RPQgZAJjcm1/aOf6ywhCRRk83+eIYsM/7JlxkuKDLFpLpln0Rs61k2PYivGiRV
2+MyzS4jyFgAB68MiQEa4mljC9ODtplsuh7Z02Ri+SBrZIWf6RMhQ2BT5slUfCHG
JsVSixbImvjahXmsjWUh3Yd/sBmmYLW0YU8quZ2VBL9a9ybU/OkQIkClcVbW0okH
sviKs83jUUzv+bP3wo8q7qEmF1SXjSjKfYk8cNza9xEaFTTyynfxewZV4bf42r65
p/OL9A0br53oRLkhbTIqL22bVjaCEcKVE82FG8/MDhLJ8OPUJ6MEDTNztzNqBBs6
nEfrDIQepEU1znA4UoFcgoylRVDPtElxJkdNxN4syRMfhmlw5Pb5a66/S91QOdA2
dCEs1UKhwBO9V5xpWkAFrYpT9xAd7NjpNqdCUqIiOyXdEoMuZhTJnjir2/re8Ml1
wyFkAnhR4tZbiznCxbbPFsqps1oxQGZbPLU5jlQT61C+j9XjtM3Zz3ooeGUuQ0cj
9weiNAxefEiu/JhFp0fYCSvzLPSXKTKAas5KieSDjRU1ajt7peSl93AhqmgPF+B+
QMbMOhCNDnkrrDSG4hj1EWUJOTES7eiDkcSnCC3kUSoAGxiqtwiwGnTCuVBmclLo
+C9yKM7vcdPrHHOLgO/wQdq5+s9Rn04JFVgiyeZ3mGa1siXlURr3x7ZSuRKnrZmv
IFIf6/AE20k4XoFcUIPNIDTXa6HrxKYkKDvhzPwUOQ6qP3eEIDHLm6H5+cFECCZ+
Z0IVzbCulPsP52jWWCo63/Y5Gf927AFDWoF8o2a9U4aUVKHiQXNIWVp8+/MTC8bB
pW0o6izPdFA77oJP68ivWCvce9x97Cj71M2Fcg/MQOOwoyBprb59ADHKyXJsVyjE
210eFfGfJFJtaVZhbX1kPDNZgFA/tkrgXTK5tP0zrlsX8/tO7pCA6DG9CX3oN760
Yy11R1teOTJRLJ5a11t7dmSJNcWrxA6xckmmcZSca1TY8HAhwfF+j8fAJwh5YFXE
6Slg9JAamw0r7XkXaLU9TwysGXYXyhLsBmEUFQpPSY4+a55HivM5w5VvxsJQCjko
mWVfd/PZpxreBGxqWrOiLgnUBkwtZgkZTE5cmAEbTJvCLNWnkIXgz5sLg49XkDBS
rmxaYJUxBhvinQV2KCPu1TGez7QGLys8ghNIJ42hdoeKFrG9bJrVTvgK5vqlqqsc
bOnNNcV3xT3Y0+vKvmSkUP1fBi+YKaXflAm6UGvolBlZDm2JduzReO++pb1gMLCA
ndQ5q6VLchupWPfcoCuAtqaHnfn5bPHLaHQFzyKlIuzwLaNUVl4MYDdiSVq8gVx6
VX0Fxw8CaPMNOb8BfLm+OOjeTS9NpWlssi+W3tkjTcyjx4+IXBmK82Mm48Fxt2Ps
pjWyb/Jc0fnVW/UiBaHKasbjysy0COpZJ0geSVEcG1Lm+8ToYPOdOs8vDk8wT58K
+ZusZcEiVsPCZCpSr8wEm9p/uqJoMQK/Tx4IPVKWSnRPC2xoYg6S6j6i+aA/JNpT
BKLyh9zMirHiSYZdpLqcxUwe2jnfnkO43RIocyR05qGr+gUTCQD3x5fncu7Y2UPc
A7Zer/EAyyq1D5PJdM+SItUwt66+BGkrA44saFyUSSwkcAFYGSfnGtZeEaYpRaAg
eOpAB0mA4Czg/QMhSmiTErkSP4osrxgtbMxGSRUvkC8rGNX3zF1nRoIlgg+wP6DM
psp4mpLlvrmTqp/bBILnPgSd9sKGhclJXt7BgI1kKHXCFbiob5wZAN1AP1FsF6ro
nvB7lNYSROaqUFUy6KhFJ+2tS4Jt5ZFRJ0sXDLf7XHSjNcMjSnA+Ld+/7qxiOWHg
sYqZGhCjm86izXXQUzyrAV29IM1i3CLo4zq3CoWjmQ41CJbA4OCgIYgxKCSwEHF4
OhM9RchFSzY8bhz5yzDPd9rMZNS2qCW0tqiwKo+uPR9/HYa/QB5RBXp+aWLNRsQe
JP5spHAhn+VcaBqUSy/kgw2p4eeCu3N5d6cTNAT22AWSfEoAXeaUGrSDAi8gc0Bi
KLXqjn/OoZ9EsbIDPG11Cfy8AF/6NHRDKMQyoe0OD1MdCycZ+Tzw/YvyehmnzDFO
oMrOIBAGcVqZoMfHYU6P8OSQhLj81B2Wace2GSn0PmE4V7cvQGlxfvjDotqeqw68
eAc1e0/aizE9xQ539bMPRcDOtvTHvu6WiJ/q9uaOuxXWbDe+cw0zI+Fc9VDr8krB
2sNIokiP4dtFyxe2Mty1Xgem/VkQ/qrOMVWEYZObqOhA+cSBCVQNVoJyNf/irDDW
eaB/wTpswZ/+8eREFFOe6llwYR47xcR04IXUO71P1M3Ojk0a3rS///ZDc5QiyIMm
5J03Q+1E/6qfecaSc0dqDJaOHaEOvD5+CS+1JPlitB7ihI6IerlqjnT41T+psyPR
IaiQUJRvDK5cYVNBsqQ+RjJIvlbhhO9FwzpBB7J7L+oPbxMxXW9WScNg0BgUAUuS
43AJY8GdMUFC+eSK2r0HCBsDUT+e6CWmHUgu9BlHtLiVSc0iYXVGYER1Llg/8ws2
NUH2qmrk85CFun5OZUdFgnymbtgKS+kICp13zaIW0fNPe4vcr2hEMWdYoGXoHG1T
tSFZmJStUicwxj3KPpz1c1phkgiwfll50gPyq93cQCocfRH0RL+O/FP2kU/WLTb9
lzBm9uAbt773eIQvLTK1GFFGPlwylCTE3nZ4H5BuNmHVLI7I01Go5KMIkErc4xP6
vAUXuE2hBo+ZxOGk7za7CiQXfCaBTQpyZh+hqtIPagV75FSssyg5mx1Rm4Vc6+2B
wywuVOYEg6MnglHbRNJ0r/gyHfvle4yGSey4KLehRcj76mLS2q7iDTWLV16NfDcT
GD8jg32LqeffEBF1QGCCfsZYDGCgePTzvU4/HXznt/hU7iQDNwOVI6Trasef23ht
6EIaoLmWMUqkqRW+M7uP06G3usaaFRqyOZCEeKwomfMAueeNvBNNLq9E5SnX22tv
fxKNB1o8AvtK5wlq5Q2Osl33A+GheUU/TWwsn2mwRHXVxylxwZpsramtkWgUO/Fv
3y8WjYUetTlcdrTBm4bEY1h96JjLdmPpFcbbFM1DwntVd1Ka7OwRiFVn+EcDIIsk
9sQL/mtBp44RZL2giBPrhfnKW+2OYxcnd3Ch0q8q4BBZTTMM/uk6S5SroD2WoG04
kNWrgHc5567FONuyNls6Xy4akyoM/md4ojXulQb7O8qmWx4PvjABRM8211vrAGYo
TnCSfyajES+Jwroy+k6vU9TQfSdI8FKvBajvy7269AtW6jbp2AupQY88QwE0xKcm
2casHMKpSBbyg54CFEtrAkbaxO5otyZ06gSpcn53p7HZFtG80dymIzUfONWeVXY+
V+WmZj5Jw1cCXBsOLqWw2enzq1tYrCvFoNCTJfi+I5VirZl7c03gHNv92dH1hpFp
yI90jnDl/QTIwNw+kgpRy3MTsdlltAOiyUJ3VdP0MG/VmTR1p1EE66cPluxcHlJA
hPF+r8DXBCGZKpEeBo2OQSGkFapoiLgHQ688/+ttIea1Uf4+nQa87ymA5pE6fHoe
nAJmJ3BISQLIIJ3tAkizVYMJYobcQJeql6Gaw9u+2vVr0JRsqgYaCprrIKuckz1V
Bg1jc5v6S1k+lrVKohcSOFDAGU3Td8pXZmgA9zNgfo2fSB9nydP87RdDq8qjcxZq
fOidZRxat2BQylxpaXy2VWR8EGGWgQ4YClh5qrNkQBihHvpnJRAPmMEHDlZy72kz
ob9R20cTwZihSl9FULd4s7tMwroHa2Tsbic6tfgBCpiIyUwdG2qOJuH1qk5APvjP
c7E/TXnvxANxFICvtY92na/E6TURt4FpyjDBCYz8E/dLNAkUHPBhZAWpJL/4I/A7
otIHH5ANq1UqKy6KH/R0mvQxf0g7XgW1u79Wxj+DHkPwelWdwNU4e+hR6xHN8rqJ
IREDdwwiVcV+9F6LfZd1J6u05zMeyVRaVkY8n4MAcdUqwOcmEkK2n93/LfIKNSXU
/1mstzPgswz3ogAv0qiRFbn/fK8h32PbjtZAZKVnrO+SkbTXqL4VTbisfM56A9H+
fpByBTVFUpS+qP9bseR6ZdSAwDP8rEMM017Lynio3boridFbcLh3AllKGa3nD9e4
f1qN12/911EynjTA2c4bZqfTbg7onCznjqL1chdWIbkf1Lx3up3/n7v2gYU2IHw5
AC2pX9poOKp8IICYBaVP9xx68UX/e/gRjNEYWBuLnWkv0eAvY+kYxosx2kIzfrp3
nmJVoRE3PXJRUV3/tXSMcwDvJTwnci6K6Cyfc7gHSJaZnWW7cJOMPCt6Eatb9Bbe
qm2ffsw01oZKztzM5L3DV0XmcphYYWOrGMWzeQzNeBzlE3bTPQPjiQ5RlIzNrgpx
EMb6sM/0H56xM2JGvuPps7COxGOef1XriLYeRlo/VWhWLWXNDkRAKWcnp223nMV3
DVcACj4VWRcija1haBi42tp5JypDrmfFJ6iG6JZ0fUmOV2MeiYqfxVaHwp/kvj9p
TRb3ENG81pp5SiPkp+bBjeQ67JHhTAlpoMNGN3IKwMwmUaIdLoIQjPqzybAeORt6
YxX1ipck/Bi50GyYc7SgAIg6Q/j9ujBtbFbTa9jh1h1QGZGzjr9d/le2gqrBc2gC
8YM+i36P83BIaSqgO7Qz6sGM9ooVXRCJxgMeUR6wh/fvg88JSg9FMBsWbW/M9+rz
ddP1koGq17Qf3vzqnaI0bRnZ0+J8gNKrLibQlMs6Uemlb/qHLYPwrPG33SbBKX4s
+BuyVCmkqrntJgVwGNUvCIiK8n7xycRDJzX8AO6L31YUzs29dGrk2AR6gQQIFbXB
BcSNOgPjWlki95t858dNdRAXv2c1t+tcWwrRY4KcVgLVQG7XKrC16VjG9qVpyYHH
ibUD/kj7ulkqU0I+c0bMLF9u1bMhOxDIVYt/wyvFi9WZdWPHmeQNu+ifid5KkI37
xYWcR2909/74qK28PiCYKDUcMBugwd+PTTynuSAIPo7sXxsqYM4ygRUu/E+UTjTb
DVzQOG6OS9PGmoeDqyLyYTgOVqHjaibX94TTjG4Md5zIg1+Oe+S2AEiNpmjEq3rx
C2f0+tDSBGdWGgNsxtr1pjuk8orh6g36GLVjRNIISgSNkcOi/lY4x8EcCEtlsxne
u6wJFxQ21qYgQCGAhDB0Opb+lsikLp0eZHj0iJ/P1CFCoN3C0tfSUccSL8JPhjnH
bkw+xz/SYgc/APDHyiFXA+0bMqUTIoWOZ4q5on6w0/VRZ5h3b8NABVaMXTrR/dgc
IG38FR1flw97RHdcBLsUg00ihRW1CdpPVdu35K1L8wFnGla/aNu6hGMjmVR1JxT6
j0+OveCY+cUd7aYZHA8rprPBwYue8NR9uIszeIWue+o9m0l/vKfWKGdteY4sVWie
bTnyTo5GleHKko2a2qIwyGQuVxae4wQUMkNBD+mjEpZtskzszIzUraLK78Z3owpD
1yTgabbs5MWM/ToX9hhzM9D1HinzFXIRu76FLmqYY6KQg8eCr8n8hR58EdEEYfau
T0lPcQiRzlMLYlrF86QWkbQxfAk4qS1/JMWDeccaZE8ef34TycQOdkw3ZGc7y8Jo
nQUW6pi4yba7ahxh2w1ujE23wTOaTZLSC8Ejrf817OHwnii1Ztl/WqchFCyAjQ2j
yf0i1Vzw0zSTdlTVPFvjJGEHN7kXvQ3Bap591c4XT2I+N4TTENsmBzz19xC7vJPb
p7vlc9+sy5VK4SGMtQND+1x568Lp22gFUP8KOExAQnH1QC8OIYZtdUJmpVkeP8l/
AUdYZD5ZhP8TP/rLMzYnlCEJcaSNOzJzBKSn0ViMxhk6aFuVKNP3vx31BBRFX9pJ
vekSYvABj3W5l3ZCCZJgv8zqfhK6hw7unOi8pU6BZAi+/CC4PiSMYURTG+cXnubh
ZqyL2/WeU1ghdcusCFXPDeLBTa66/sbJN+I4mgNLk2IAL7QHGybBtHCzLCPBC8rB
kus2ibKI5c0oEBsQPMVe31LJehgLf/GD2t0BE/+p8pPtXwlJ/e6owptTtBIj4R+A
8oEmoXnV8pDH/A0eVTn0hVb+e6AQ+4hMwXHfqpqj0xZQU3nWz2+h3SHoDb9jemGi
AiJEfcPwc4BCalY+QSiPDNE4AIGqWuLjSJxfUZhWjcyhSzaL6OhqCJGiqOnXAsHf
ieoSnhAyWBc3kN/Pja0mzInyx/GJ1o8RAMqTGy7qWGC7npn3yUHGWLNIRROoeGIL
m2eSiT3r1yvILGyKFgck7OC//CDALX5tJPpcB+oyqrwgY6hZETGpfkffgn1RbhIn
vuhPQv9vtqy0LDHX62coOG8r9B47VHp6v3W9LbBmR6tY+8V19mbGfyPcyRNvu04f
Wqk2nP3eHGsmWpKlkHq1iYan1e2ZBgSwHQOnVgsh4SJRXOuUrz5xdJ/pA+9ulSbn
5K8pzY3blwgr9k8WFXssjga/FiRVXWXYSp974W3I5uh9AWn8qIfp+AAcbfDUNSkr
KpLTZPULHWQtudC79mooFLXIAaWhUzng67E34flCpxJskx/ivSOdtNM6McB0rB04
ByPrYaPE/YBFmz0p9x06jpn+OfrTuuEjSpUbOhg4WSM+zr00FWD6FfX8XQD3TUZj
8uuw0lUZzaaecQvDqmPy1QPu/JTECkpjlXnkZ+CTjEouGamoxwImw9Im4t6wPVf6
PjoayQjAAIzBCLxjIl5NCxZ+/Fvsz29ssMryIapXNsOLQYuEKtjIrO+zNWeKs1Ux
X8A27AcZNMtuvilJ+KWUeKNt1TSbnKGHUP6wHt0YnH2DnC7EXYZm/RqN844PEZVu
i70lZX+y2t/tdOvq6NDaOhSexhgLcg1cCMvjhrBavXfaK3KxYTPOCPtXT20pXB9r
ezb8ea7VCQH+8yLxRnfVlFgkkkWtpgbN1H0/xGpB8HdRcel3TL1dz+5Ybz8NpNQm
Q4wLJHpuG2tq1hhDAZUuBgc2YYnNIRgF0ptx8SEvsXrGiBtVzflUM2XOgBPaXgUk
Uf3aAhztCTCaj5SDRk6B9XhxPyNLnTszJLv/NTRKBeG5kVZ/Vp7kDcfKtAvuQlWY
R0mwVYsRDUV6td7gdzfPUl+DCkehXdxGk92y9x75xcFCdI9SpYBCUHQZAUdpTOK7
xwmIfaEQORLpw3yjvdhFzUxzoTD32mEIszd9P460Ei1sry0uHdaU+8Xry2hO9xzA
B9OGqACmiymI9i+xEUF6MpXenY+dsQhqLm5I/L0mgMYShkGVTnrUNHczUcokVpQy
vHc+OEnLRanG9ce/ZhT6LBdOnBfV1p8Olj6GidntjW2Rf3cZmrcZQ1kDQDSM1SIE
WB4Ke1EmTFDnP6My39nBArPnV6gKex6aCbALtZcI8Y6+SwudsYViZn+6Bo3yxmXU
TU43fL30IlXPF3Bq8jh1Y42Eo0XPcCoBj1sinV+Sm6oMRcJO2FM8mtER5HfhQ5bI
6cwTxolZB1e2BLVS40Z+pr2/DuWvglc5Bgr28PTOHdhLG+BxwY0Mt+/roe3ZcSmv
zvsnOXLuTX0nSjpCclRqbPpvoYC+9gzloqpFduwKtEOHhwP72SqLeoqgwTmEcQ8D
OmrFxkAcLgcblJ6Fz5QaHh85LO/Gb72fsrS2a4IBvyXJiwybS0yV0n5iDlIb60VY
CnhFKf2O3t0A/xu/Ln/nSX4WuibbmXtro2JuZ6YKbBSXxlcHWs4nyIctmJ+lpPm0
7W35iLK0M462kDxOu1GIk+uh5HTwdES1POSrgHNQI/4/8WPSBBYtt7+9hdZaS/q5
RkRNieKSz+4uQfl28F9M4rzhHQmyecSSSjoug6R9ZraWyZ8Ancb5L+GSqvTAEkCc
ZRs7or6SUhDI+puAF36B/uvfOtQTMjC0jDN2mA79BBa4XxFDTjTxUPZ4Yce/LfmS
MMyDiUFPTPq4CQ0lQKgKUcYxCNgBc4G/s3kN1Kk9UoDLmDpGBA/ECqF64Vo1VXdG
zQenjWRp6b0DUyqo0JiBkvDQzBXwjYMRpDffShCKAU6r9i7GO9biIbbBVNGaSiG/
g+MCdftwRwHitr1u9x/ozKF0IijZKsnr1BYoaUT7TE8gkCJmpCoj3ADs4C12dkFJ
VavnjMD8k62a5c7cD5nspx8T4fCCfvZd8Yp6vWMy3BU1aX5LrlZ9d+a+MFwCujnf
XeMpV5oaM++I+2Bx0ezMQ0KMmNJG+LciXVzNnLzU3VF0r2NhLzQR4M1BZx9WDDV0
HQO1HLkQXkyhb74AS4a30emQBgVmxFcK7WtrmuZ8pL1GMzz6hkC0MRB7kid4YABu
DBjhkwB64rbqwDYJBjiS2GdP2qC8NE6XnYP6jGK3oKaLd4UA8tdJ7j59ho1SznYC
Pk92xVOw/IEg3o7dpOfZF27Y7Va8poxCTEWL2Chc6Dod9Z8lxjpaHjlAuZh6+SqQ
r6cwBY8Rqyd2BR063W2TJuzPkoHORJaP3IKdtBTDu4towve2Bv0iPOoWpb1yZxRa
cdusnMLDeRKfnUN0BfSEx+3t83jqSEzIrVSHJafm2kEev4FpcziHjW2ktX+eOqt1
2iRh8i5WP+0mr2XDqyCgFaOLPoJ55H+iZztyuFtZhYVXrkEWUhFxWIQ8cDyz/fa4
zG1poF+GXkMq/lisK+/uQ4RpIHuAnT/TJdIS4AItpE0HzvBBoULigv8r9ouaK6zv
RBXs0yIAZBLA7fsLewtFhhFkMkfkgSn6O9Y9/pr4kZaZ56fhaDTTn0JxCJ3xTsec
B/VFtDV+BPBV+69II1X6Doafgd9DlAmQ+003JdT7JPp1+7+P6/tvQ26+8MD2iZAK
wa03I1GqDJEsTUATe1hSkV7VNIOGt5PFs5lKjuP86xYhBiQ9kUVBnrxgaEVZk2Ml
JiNImBuVCgUdK9cxC1AgRzEmz4ATLFPy6ctocPRexMTReJtjR3WAu1qT6oryvUIt
du5XvAD491NJ3CZ4NayMLbt3IwPRqyNELf//XbXNrfedMJd9SrzZoFsy/84B066X
V5JV2E63HJXLV9OH/Tmiv3WawUqynPDWG58qy8H2vpaErUhaVt5J0ex3Y3l2ca88
zWprWna1u6OL18zHmcJJXXKkUVCrpUmzCA5W3O8i3egJJrQAj7WjAr+O++aisFSU
xyUAFruSk7NVC6J1aQ9I3IijrX2zhv6zd0vqwn9j/ADT01jMjRsNSc9L71u8kvnM
7rPGlhEARrUhlVSf+bEZC20GAou5HYXD4uGJfDExKHuUNRvE36dMxh5vtjnN1BoT
AtHQp90znOwG0e8WwFWFoI4PjSu8HwbulmTu5xwSnBT0G142EbdlXT01kI33Gpo0
6nLgBaxJfLRF3ktFWIvzIaOHUn0WQW6glRL902vfjIo9S186ELn/UNsOAfaZkVOA
e9Nu5mMRbDJsH8TVzLIk7ufmgCcOOzAqBVx61WUUNbFdi+/dcArIuOQpQbATbwvQ
EJbZwgUXFb7hf50Z8UPnErJYlrNwoLRW6MdzFO/AjbkRy7uGYiSYEr1lhudm6Y6s
+oRccO9QgeETSBa6GRHSS8GROFfWpk/JnDw1JSpa7dUXIIeFlYbMyWAk3FKI7nXR
8N2aF1m2DOnRQj2HwUkm3h5lOctcykDmpnJq6gvWGvHWSiL+zE5dNQ1AVMkEoltX
UgfA1Kfirg9LCzZP+8D7dFD6WbDvQA6N0U72j6lJ7d0w6J4QZNKGxTrGScQz9PjG
isdpoHn+RKMp01s0xFIsCjDyBKL7x27+Guy/HVmofCpdZZUMbu5QKpnUE4YnYxum
nOkpBKhvc6UBf5Yja7aHZJLsJ/K1PcreK+OmEn92vtEed4YeUSF9aKs6mIZwHixJ
q6VBRERzdGc/OCCmk7HU3c+5JilPE0Km1XHwQ1aseOfPyGumdnsTWzyLZPjSo96c
y/R0ece2gcDbdjRH61plj+3tT53JZ/jtJ4yG2uggK9BHV/Ulqvz0d26i8PFGSUFk
jW5QuEa/34myoIRxnylshbRNBlMbhJIuAwcxbO4kBzZYpQ9vKB66/xbBk+B6e5gC
iokBp5Kw+XLArTyDagbmouuidIV5nB/matSYp/z3CaLoZMbN02SGxfjLri43bJuE
cpsTO3YmduTb7tncaG3fT2xrcIHNmm2f4TDWn27vZkFFZMIk6dqbNo8xLuBnHagh
Tp8EgoP9Y+SMeYfnwrI7O8+8IaUqtwenMa8b3/qOD5hVPry9xYhmuDhodxt7mhXa
6n70rzfMu4FsdlYVE4ujzY7A9qoZlr3Wnl9yL1Y8dpy0Jb548FjucRmQLV+mIbIi
4HuLXVVh6j4L1yamKC4DF2uIXa49GNQi/cItMuM0LV3sZccFFuHiA0V0LnJ0n+8U
1KKtugRw6UBPP4y4JYqJsW0c6WuSnkXM5Z0wG5OxHf0y6v2PShSv0aVIsBXhqade
XwA6H9qH9Lz4GjR+OeA2L39EK1OcYiCWAzpoqJi1VA9006OscM2zoobEUSjArN4B
Wzc9fkVrck+/GN+q5mJ3VPZosh4p299adxgCj/jZn0fClrjHtrpFasACzLsTB7Ip
sBOYGQ3xssbZCsQkopENrYVk+ssdsvFokN9IBq/FusESKjFbvvLCrVaEmN7iYyxK
WuLdcVSu302NRwcsV4D015fAQyKhZo3+gCfnmFaI4tNakuRVfwC9ylyXq1j6SXbX
cKO5l7PKSwE+SVf/ZV3KaqeflZkAvWx5ojA/0LL9PHlCxQEhpxFXmwr5POeiXBZv
j72KDh5KhDNHTbFkSHqcvf9G/dcNtcA6bLZp+6MBfQ364QHu0erqcE+pbV6b+4v6
TJBtlbD+zkdI1g29XKCIA/kaQtqTUzKjIb7ryaZpo8bPwrNP/kuLyI2451KtZjNf
3ItxeKjkZUSEuVNNNAPYtlDpI7GLu+F/GlgWIZZnHvjSHzEDniZ5xKKf7jMMgVnt
vJgMFdKUTEJs84aggMYJV6MgRwdsZXvwP0TsfKFJPcc4b+fHUy7O05YFB5n3zlqH
53Qtwvtvi85eI6jPWwsvacmwKZE6OnZxP7w/ZZ0j3wSI4A0C7FTiSP1E8UVkaX7c
DOTST64RZmXBYlbGhj2KMzDY//RYzyN1JXqsUW2x5m8F9LAxQcevxBxG42usrLg/
vwI691MLFevXcOR/W9+yOfQoSy5rhC6kkOPrHRZMkJx6H+SoeLhhc8o0yuvp2MPK
VA5B+1IkNAJv74KWW2aU6vaj5/4nt6HatfJHXPiJvCYveMw1VounGTxdIYsaRnpw
XSNQZ5zIwQu/KIZyYMZRllDjF3arNo/QtFhjYEnQy26Msce646TlKzTzAhFZADZS
Tx/0t7gmKcmPrJ6H03Jp0j4mYEkJAktpntePldSEpjf/ho2g/gmZdOqSWZ6c+HhR
anTLqMM8bfLu0UFrAVku93UcUxE0lB6QIHtFsZamCu9ys2qFNGtN/UPSc3UeAWi8
Ckc/313gDKsMzA3VjV231MiiTU3K6Gr6zfHkcOUD6fBkCjeoNVk6rg0+MYP3dS+q
F3wOn75Z+S1fuJB8owv8UaFnEH8irFp1ZomnBLZ6lI+QQmLuyvz10LiS2nwZo3rn
nVMOaBg7dxdmvbId1VOtZJulyM5CjbCemFy6XnuCbBAlil5N7CIpTPr4WntEmHzU
aG6pIyjm0lFHir+eNfQKwndHrRrWsOdoq4+aeslj+dH3u0xgZXqFLv/Fg4UJTb4+
0LSgOHejDDuDYx4gR3ET2tUJnLG+8FhgIR7J3KOWNxIUABig8gcz3cCw1Gc/kIAL
kl4W2keVe6KHCkEjk6TnzanBE5Ku2tDjBR3bcJU4Hw1htsnbAhsdVwgly0J6tExJ
s/I8Loi3ZivM7146eeM834xUWRPfkzmjOKNeQfPbyUxyKD19uByMDkYW6j/brYsE
0xKxNEool8IS4SWeWFHLKjXnxqn5/2HhMReVidoxLXM1QhvvS7KrLE9NxfrgexcZ
g5XDCS9AJnY1hQ5yO5Ch9ueinR9JmdpBqQGa6YyDW1JxKtXFlXMnGEVEQypkElSy
U2JSVkFYBpn86Lu9cPTi6CnyJoRLySeqaXAeyzvGsWSmjAlM8Q3L3xuDlOONx+QH
xNJ5S3YeWanLk0f1sxHz/UnOtJnxLFg9kjetRODqiLuPXQHK7yjC4Zf2uMeZBqSZ
PM/ReieXE6U0OPk6li31CHoTuQL1q3oxdlmflHucuKiQ6HuCd6ztZwOTOTyBqbqb
aK+/hlLRxFu4BLnjdYUL9Ha2ikkDLwV1uBKtjrE1lsdobDeqsBGxuzwzGpblx7f+
S4ZCdE+CjZu43KgFHOShi1HNGZrUMzFZ5srGuA6BscamuvojpZ7KV5wy89QvLFZ4
2O38NbNA0ShN/7M/rlKbao6aQRfQXsQKsz6SC99LVD6bDIe7k5qOYvW6q2zO6Z90
cMxGlh2t5qOvmHm4+7ui9hUauYMXXiAAs2+JUgDTBJ6CNQC1jqKY0nbsbNcQo1MY
LlJaaGwWt7Ffed4404+45JCuVwpJp5RT53jx0YOFlLOwMm9wZbDuE8ZL1hINoHn8
GvAtk+ch3kDP6Xe2sqF8ZVcbLeEOnb1nn+PiOYRfFK4sL29EmcjOqSb9FzarVFn8
6JfweNJt1I4MXBz49vQfqakleMhCPJYHAFLC/xpbmZa6yUFz4Ccwh6ExoJ5tVHi0
12M2YN5INyNLpZk9/yXHyL9z/EM6Urnnil16diaCeQCcUcnG05ZqJ4rPj6JT1UUt
Y442NK4f7+w5pz1BfkstMFheckLjuDVGegzFQxDLGM+t+iHIl7xEfb/PVpJWxE0G
0gZYjc9Akn2bDv8OtUSbHz7/tGbmAswhp5nKNgrdjyn6y3GXcyzJY4LLniCr47H6
vD9nPlolW5Ixz4Lg2V/NXoaVUJc7m+aHVCbj/FKc7gwClcVca2lB76Hva+1Lmltj
u6YlGunvTgiBuZBdUsj78s5BVkxtz3dvx10yxtp6xDcmEcJbOe/knOcoYLo7wy7H
2t6Y91fehx8i6w+IrxK0WEzVAYuvWoVnbRz+pavhh7mlHwflaqDEb8sk9TwIsupD
w4DwySH9oTSycq3eNCfx1KTGI+P/HG6ONVNDu+PKDcn9XI1xIzQW63kmGHzeGbBr
AGgYiZrtrHF0dE547KvEmJwA0gr+Q3rwgoxHXkLYw8lBZDb19HADVw01iGHZPRYV
vUUe0iDXbN7UBBEflfQg83ATwdENNz+g273KnqaU9NTvjh0Hn6hAocNtin9hdj88
h9NJOLSVz2v54M4c9WVc3KWLM+7uM/mJOdg5t6LdJrjbhQtAVne4emztzLsv+GuE
PH3xU5yx7A6ipPbuUG+SzN1zpZPdjJoecWGAvBdCkPR3mxQdc105aWvwC/7xHjNk
tvputMOE3Q+OIB1JCkuw/LZqopoPJaH/AMFhszDBtJZS6jksXNabIFHYdJbg1Ytd
EgVOT4kzLfhSilpmFM6uM4rlUBljoilYuVyEJEeZxWxTBcNaFmILIsfWFfiHAEBJ
C8MEuU3nfO/3HOe3t7RltvNhH4sKgYKhe03xfeteDIvRV5G+GSs8Um7umZQT54Qf
4mmE1kLIqndqB4vY4LN8h3U4qj0DoXXkI8E97I6IqU4tVDD1rtAMJ3hOV7a4IZce
xVtCr0B5bKGQcpMAj86J+RDCZj5LCOJ+zrnm+59ilTEROq/9JcGI2qh17Q+jwV01
7BRN5uZkPwj1Adz9L0goc4tiPh9ELrE5XOGQwQdNbosy34DG/KjmejT7j67KEO6S
b6N6Xg9eWlwnMltoCsmvxGW6E9YaiasDj6ins2nkQ1vJ/1bRd7JUt+ekNuScOfDv
ymO5fXeKTu9fchSUzmCKMlICyBWAEGD91qkmUCWoDUMZmZRtZPS1EL6HMXile9ff
JdqqYVIM5abnyedWgpenfuu5aoJtEVQy8JHi6ZVaiV7gx3ITKqm1R9hkWeIxx/CA
Tj0gNHU86AB6GWhx64f1inlOwznzvbCHBhLjlRXxmKVH1S7R6XZEmQIwy3b4m0Cm
rw7feFypga0KuHXxsT5yvRUyPkyLEe3NmfJoes6u8FswCDiMyMd1le47TtDfTJx+
KfbcWb3cKidqYTDTMPZttrbyLffQXz/jIh20YFDEFQL5e4vcox0fMbikEhwehRoh
bMnvgGCtfXEbO+8WrKmduKLlxo4PSWQZbngzHlkmfJPCFYv694eQc9yf46pT5EmL
cMasOtnx3RuBV0JvRRWo8GItWtfGLhCvu8wWEOt5xK/07gyAtsx3B39AfhOgUlIz
5R0MzQ5z1cL0IGfC0UhGeXkLOIHLq02M7KTDiY7nGkowY1XZOYCAxN5ldlVa+R9v
ecqdHnDVNGB+t8GuxTjd6erXx4sEWIPYrRoo2CAbHEj76/MrB2BAeqgiCmof1tZa
tQ6inYPs/Iq78OvfPjU12Vl4JK2nJ/EbDZlWC6yQ2MYD0sZ61Wx1HWHMfjKagwcC
ieuymZyM0VzOZFwUDMnSwRP4Cu8v/jta5jbygIaXhO7ghIr731hZag9svJny94vK
69nGA/rTjkhTPXgDbwUUmYLTkOLeFK41DRcRwV+0A8FNmYW7JJg61JeFZ0tQusZD
NCb6QJAHXZ2V5mpWaZy4Jl91BcDgRbkDMrTXME1Q+WG8eITSC9FvcrJKm481m2uN
CLp5GjLAHOg1I5AoxzvQCBu94tyb7p3QHXHwHfw0v1YuO15wH0f5RtbXhm3eK6tj
7z5dIz5Uq+f9U4tHmAqeaelk8fwpDbh8EeMglOFOzivm6dKIuMZTgatFzMKbDC2w
rpJZFbVgRom+/p8h4LZn9hCNSMLADaQsZrpxcZgV8UNewdbvMLxwt7z5KEWBNOaM
Z+eNsQXVWOAA/5pULdRx9YQSmw9PyyKvT1cVEATZQ4twxOLtNpgYJFzQU7IsrZbp
gvCL4JY7v9tq2LlpbSFqNN026g41xSSfBbS5CQZGherKkL1qjR0INAeiEjmVBRqw
7FoJ525jas2AI4cNY/Mx5cH+D6mEJR/cuxzWCmHgTpRfNOB80XX46CyFbjVctt9k
9LhEzwfypJHGAjoHhPC7wpcbHiGVlAhIUP0B1AE6jKT2XS9fjEp/SdHjRrtO2wqb
Z/SFlZzFKnriBStJqTtBV2Gr0xxgbuYJXio6q54ZNOlZiXb7SpqO8mi7Yc9cWV88
Zy60H0AienfY5OCj7hqlGdpIfyp4SUL6KLTy5LifusjE08+bYttM6nszSOfKFWNQ
lGp5VcfLZ60uXmTstUc4JPUhxoRGZ1/YsmDuADApubDT5YFglNcy3dRIqzIpw9S+
uNoNgeNmexvDYiwOR8rdObcYcSLkn8k3Hb3Xwb5wRI0UZChy99V/qouNxeCrd0kG
73/b7pzmuRVgtP5T+pCzLz13kK90D/DcEPk/R+mDASuWBJPZlbQefEv0VqnPgnJV
0650WNr9/Bkbl0cYrezRdBD8BsbARlZ0Ei6JJTqeFpeCfgJk3nKGXaCLwJ23HGgX
yT8PZsal+84apVkX9JxsKYUnm2IG5wUfi3FbgGx7fxpeE0n4O/nPJVxopja8ZjUk
ST45h0BKXp8bMBNEenEA1RXc6whR84oD+HWPeZ7uPuxCuz0JXzWk25WKl/XSCewF
L3ChD/sES+KL489qNioIS52ywDfDeZBIAqHp/qYrIrwOE9kk4V+wGtG266igUyMs
Fk97rkuCuBPZrJ8vnzLGKKX1xlk3zLxvAfIXDgw3xvjyJ8dKA5Jb20JgUJJ9YN3R
CWM4O2IOMBPXkd8oVnH5c/iaXyb2B3l8ja6iuk9g9GyacJcZFs8+rTt/hXKk9oyl
ZMgsGpjto4kjyvg9I9IsBO+5WqmExVLYGMn7MKy5uSMAGqPzvnx5r0RW2MF2w2Qv
pOyipVUmANKjuvfIW1zqUk6lq1VoZlSpBoHIDibE0n//gy6wLlNFjN79QZzhmJpW
QiJRwtYykj/kMo3fINOVbgRAmx715mCqmVxVd1UGMgnzjMr9+eGIRlL596VQnhq0
hZuhFgCQiuVk2NNE0jZ0ZmtBp3UKLT1ozJHhHGLOZuO76L/q2KZssYbazx9QDMeu
2NJisBwFpgtqml+OaqD2MRqXnkHBClCXrysJOANimQanquRwk5SfKGPtUWu4nBeU
WVljxjohqcpnq/q/wnoTTUVNIqfMbxMwYmUvlccdsHTAU1yNBFjWMA6ncy8E9lOh
cVKVvZw+YyqvkypVDpW+EF02Yuks4k9CTXkmH0wqlLStOCKdlynTp9zLdisawpcH
YUArm5Ijzv+T4PJrQKpVAsidW3pmaj6MgTQjy1r+6XJxZVo5DBkEWBLMmrz5MNUN
NQtTUARi2zsxzfvSq0q4D0iUHQiIAT6yn88F26JnUmU+9yIr8DaPUZ4vvn3jfYF3
KKdfpELQf3CYV6LQRZoXIjBCUpOgTex0ExVFnqc0+e47OUNMyMGFO5G08srh+10h
pHiUSGfP8w4yXGUMHPpMWusocZ1EjGUtiReZaJ2lJFBGr5Eo7j6YbkYNqS9/sV3d
yTvDVt3T6afpnWtYUkzsUhzNMzVyutymKLg/OipHMm1FZFTJ6HnfOmvdgHQUKU7g
4/b0/RiGtxedXAh/bbMctbgE7uoIBv5jjzqwUW90e1lpF4Rrpdhvw6LPLMHyALJ/
uiFgZj3oM1Pcvv+Tf14O0WnA/FoWl53WyQBzBc52W7Mf7QVFaXyvdKv+TZ23QnF6
UJvnVITAwVronArZHazxpb0rd8t4NXxm99OTZiipKM4WsGMDATij68IYBrKOI9v9
acw9wtaZ/qnfIBIkJyL/THOrbpN7qzdEZNMdaregEK7k3Xt1IfHW/bp3Sv/IZ+oX
A/AD5Xzfa87pJr7XwjNPl0oJSO7SP6Rvjq30jWboH1JJDjPSgpv9SN4mN3n7mm+8
0WbEn6CpzxgXoivVgl0ZxCOpuVAQAeTwG2hkZBnEmZbexGc4BGFwyBBS7TxJ+84T
8HKBFB053qnkb1hywm8Eb68ghSsHWVjQgjHL8zOUxNq2SjH8/FZqR25B3YOtm6Dr
KfB+9hdnyLZJf2YA26ED65H3+RxNEhHGdMPjb7oSjBGDKuowqn94Zc5d4ueZsfhE
B/FazLMUSt9DKsYw2vLFXz6GqvoXRUPAUGiHeVdbT0ZLyHZcdsM+ns+kEITGyZSr
SFune/e3S0jVPmzUGFreGLgRUQVeAB5oM8yOrDzIu2Vy5zwguD5CcQ8PlP1WSpLU
PNrpXU7frsfIv9T1lZoZh+n/ZWPtICc7q76fowJkbW6EPc+y0LjjvjE05B2Z11Yo
ZPmD5BfgxDTAnQLo+HXC8S5N1W8JTTDF0HRa3F1j97mq8ODMP7/VuW6TT6fAg6yi
2+1UJrIFAlG0+oEacpehZtSbrm4oO+ShHOl5LlFPMZKsT/BQTQtQdO/5G+30+YfL
P6t2b7SiuVIoTbsieq/vwzL5QJ3FfnC4eeggAy4RhlvwtcwdmjYlOcTyWpJHRgod
udhlFZrachsFGi9Ek1+80BewfjvbiJtZtnx52OUoPxCmjui9KG8veF9prFCx/0uJ
Rj/J+jRjxLTCnJVX7GKRPpqLFNwsyaAPEMozsB4S5S+cXZz0HPp4sdQBUtQsRvxT
hR0fM+E3+qmCHY2C478xPQeN6morcEuGnBWdiX88xgQFzX6Z12xz74bIvSNptmax
4ZxxoBqTsEDECgiKkRH+hxemlvNqZGKfbYYBdk+kyaSoiYvLT//q+fyvobU7p2gJ
A2KkOd4rwMNOKipx1ZOiBlXmPOXKRPXxF0cyqtOwwQRJ3OvSRoyhpyzclOsHT3Y5
d04cFBkxGB5ywOvQjVQnoqKtVb3lhmVvpK6o2lMA/bfW49mrbVFkn0OtTJE2TWZt
tN/qS+Xg/HOOICqP61Bl2VHLGbnqY5SeETOqDcyGZoZ9dOmYBp/Qgvy7NFxewEB+
hMmnUZPeKyaxIN3P1NTmb5s2XfQ6zBPzNRbwtsyBr1MP03ioMR97wc8AW6vifzWx
EbCrXhut3Le+l5ouZtZc/55Joc6otlBJvh9/QUVvhbwJpO2mF7YcKRTZat5Ol9lE
Vf2gx7za0EXL4eR0icCpWSjIra95s4RGPEBF/F+jRrQYck/kp6santBZijMNVRhH
5r8Wmapql8n0V25YxurTOAf/lublYtrE62e0Voqbnkqkau6st36dTQI2IaZU80oa
Tp6lTJoqD153/g+yOmVgJ5Ku/9MROQEBHJ7086D6sVtwJQArz7E34QwF5MKo/KV8
v8qdgMdxzyeS5F3gBU4xjmWmRau0SHlsIW8vsUjmhzQiYryUM0ZWDuBnl5sUE+JQ
tduV/sR3OTQCAWbbV6x4duGMPgmVKu8iNEwn6iNbGb9eMCDam/BM/I1kXeRkvXQU
+OmdiJ+TmZX/pWoqZHX36u0EyREjbf+I+paoxIw4/R56ErmqVGb/88vUenFNeZ+z
hlEb19ox06P7bL51AoVS0c4B/qJSG7FhFG7DE7DbVkAyvsAMcfSPhDyay6qejrPL
L7yPwEw6Z/J71543sd5D+T2cd4UzS4Jznk5FJE5oRPn/7R/ijJZSMjv+Bc58HVyp
NihS2/IQkfsI5kNapZjmz2IIKgMWf/y08JRYJXiC7NXtz/ZxtK3uWhQzzr1ircb6
TqiwPNFXoX94Qk9He8tABUKIarykIgtOxV+KtItlzkDxZZCA2NW+0RUAWmUVGpbi
2cO6IFry/p/Dkgw+TaD+3yDfePeebrnQd5F0bGzmrB6uWjGDgbesKXcrhViQj2HR
ze4fzkoBu4GwdEd/sHKED5SUw7Q2hFDgWGh8qtMPWo7LLQqwgXcSsZVlABtZCyFR
HtS5eUyeYJA+LseQAoxtV79M8i5r1Vd0fmc/wwcMu6rP7OrRvTxNj1AiPhir6wGN
znmnlFA7JKWOQ6H4Gw+qvrrUW8W+y9kxFp33Nq326icfOhy6ijbS2/EqBFNxuycR
idwEJHs0Adsbj6zmAEPoTEWNnylkzMQ+ifWuIsJzO6Mra8+hV+kDwZ7oQRAAmZQR
1zlNzrmLmhd6t2TiM5WzG8yyEujIEC+oWatfQ7YjduYGY3UvFmEXcuIv8XKydKqU
XwUeSAJzlrZK7H2blErYxEbd0KwH+GYCgMlm7N8mrB20E+p8GFvqzGytN/063WgJ
fQYt7J2WgT/xWtZLP+wBbV3+ix7SBr/6ofWW6Q5f03cJNcOqVCwEQFnJED3AfK3B
cm24LaWjPa0qiWaTW0q6Ffyd6o481hax/2oFjGGDANtKl+NuvLjHeDCQcpPusOGS
HL+MFcEscIoCaUBUP0b278Qce2GidKe4gAvMptp9+vT9+FFRjO0vAWiYMoazAOdv
UeN9NMRIGANF1l7r7HtLT6porAgFG6N8K0m/PD1ZU6iUlxTRVnaFOjs6p35W3VIq
0g1lZL1mOLg1W0Y6VQoT9WydmJisvuyMnImLIkcwp7X74vsml+DltSmASXHND34X
HArr6rhSD+LtT7ip4YSicbl8XIZ/5BDC28Yoi9pPzZYHLa33I7JN/yOmDmqAg/gT
ChTpGSn7cH7TtQCF/V+VdekcOa3WcaMuuedE02p8l5C5wKMDzyjMwYst5IcRZnGe
PO7WSH/XAD7ae1O8LTgA4ZizxwiKQLf9uF6QHHV1p9KISi3nKKY2lyXLfsg1u0Sa
GMgurPJYAuPELgGZP1oZT/s0BXpLv2RpMvAda2+KzRoE73iqgdjWOXTOC/9CIXYt
6f4st7wDJI1HVyOe8o9Mk0tgl9FQSRCrj7kQah8GxFAA0qm+uql13k6n20FDnKjH
pMypT8WKNoN0d4+uKGctFcVjoHL8zrW0+miPvI4E8bn1KX61BUSs6dfDMYxgIiu0
ZP4S4cW3CvSdwC+8gDwH3bj3lBYws1hvoCwavIAuBhBqzux9R/aUmb2td4Cql339
5YlLHc0+z/fAZLMIXlV6IBpNgKXs6oJWNf6dpVEDaV1skJFi2ptwEoUxRzsX5gjU
O6yAbhomIKDBGXd8VeVKCFFAytNTHpoLeCRjwoqkuRLFvBNU3qbfCz4fvMH7Tjtm
xLFN+3vbtEk8WBvB1129KyAFTdh6qQ8TVNguWXe9fOxRjp1spqlNPKc7sYnXkFJC
mBcZhgbJiTY1hCutOzkIirOUxOCFU+Aqn+hr6V7UU3ZJR6BDaeW99BxFncceeTWM
agzQFSqy5uqFCNPBs8J/JbLt4Msixj4YjUFlGrW3AR+gWcMYdBMn148kE27zl0UK
L05aW1tLpeA4sFSRsQs5q86UKsvX2tatxj39Z0tiSrTocdaZJXGx4m48qkUP0hdI
MtIrPKGOx6CBzWKLmvPUr3qKuRrCGtr9ftjjuHaquwISWYW8leKR3wFTuOscTmsK
U/4QD0va0dKNQMizT5byI7sKvUAEV15Iqy+psSBdwc/j2O502RC5WbOIpKCiSUER
77OqYO0Lu9zjD+RbdvKmQgLIdYc1XAjdM8tILDQqHVS8kSMKR9/YHIsDE2QldPKs
X9g2MGIuNab/G+XVnfQ8sN7nM9jt8oln7StDtb0XdcaHxplzpK8SkNjLBsz9WKmE
zG6KtF6F5Fp1MERgq2/1JkAzGLQPRiv8mhvLV5heyJ/8uLYV3k9o28QCTvGHaMin
jVnz41PC8q2mtPuxlj/i+LZCxa6bySWbd1+7VHNQ3cVLQKtnclCemDSrldCOVyVb
5Bs1mjpfJAylDqdp2in9V/wbqF6F5vGdM81IEqF5tTT2dlPMzRl6pHWrBEcvw2ru
ccNIRLbYatkriM0+z5Ur6GLcsPXr5GN3be3tNU5TGtZrQmaYdgQg+bvrgXYNudBr
Q7WN4MAwsN45kK3fxNXsoiC5zyT7mr2BwT24+bdkkPGuwgoHuVW/H1SA4Ywe2SuR
kCbtiNV2Pfq4oGGqUI811LhGiL+aVpU9b/X15f+ihKS2rL3W73KIS78QimtRJhg2
Zvra13mJIC0Pxv9r+lgeRqNt9zBOSYVskalqfwel7VC/wenY7kUOuGGwhV/JhO5F
zUPw+v58xD0SmO+wjQTfENaCos3lTF4jOw+Av7VGXAoe2KTvz20H2Rt2v8koWZxP
/ZuhgSRVpxGvPdgTqYVzps7kuF5OdGaa4qLr1H3SgIE5wMDACSdYLRlOLWwvTyQm
eJtJgwJzk2qaz8Rzv9pQqjarYcW9oWVraPYxF+TwCR/TKz6grM4rL7Vjl5HDvp3h
6kPLn6noNyKq/K6HUVbmz2gwY/E29AbdOgO7pYDC3jplRlJ6+He0lCgEzIYNReWG
slEusnluReLWL8KwSyzvbDXj6pPrm8QRjYWSEpGZa/9gqHOIfh1XjP2YdcBPG7ba
98HkVY+2xU9aGPaePh6/XSro+afDE44FXKaGN1A5/Erh3SORPve3GZKUwpRtewy8
eZvjG6GPrt9y1+u1EyweL64XjI8F1LEMR0taNXprzQOel2m7bh7TvF0w4XIZBVwL
1LQBZxThkhIphbr7U0MNopFLa5Q/H9SFs4CJh0mPhwxjfoimfH56V1JXfNgo0LxY
/Av3acbQEXC0ocU/5ZcxDkryhljPCxEjUdsbcwQzDfdr7Km+IAidMSiWwf6yAfx2
CvDeZeYJgNxJLw3B4TnQ3QzntYg3ugyISVqzLVHbDk9tBJY8kaW0hdyAcLuKfHBx
B7HnFSTia6zmvpQ4QZpt4npd37xW1bcCPi9y/usHIfXF0Mmguuv5w2cAxEuCtz2t
INElaMUr6q0y9Fc4kqWIzAIG54A8jTPrp7PWQhBYjlQioSHPY3EAKtSTIksuevAT
58iAz2ipeVkqte4apmqUbdDL9/fo4w2+PCdijq4VgFyfZsZzrvl2SJp0GXr5/fVY
AGeS6Nit+tryXm0LdE3qeJcNA1iB/II6VvbcoiWTrpDq3jSxuABf69VTkdgTgInQ
Jt5MxLDHbJmn4FfRJgpdorGugZgmXkY7TRpvIO7+A2s4A+TFfUQfbtzfLHZA2sfQ
OA4582U20Feynlinj/tpUcajZIbZ0NNNwQ5kFyCOmXGf+qCBhgMqJl5T3XG568+q
hHmm0B/VxFxp0AgosCqfChYs9/YbXDHf/H+3EZHUA08OzMtDLE7lIXQERoensvIb
mPemfZVwtqQxhxdP1dtySNJmTjAXBox7zcJicmExHxQiOI3kHvy3ch+NZJZL761K
e8UdnbG5fmJj0se6hfZKUQUNuTqbLSnLqY1A+ENBviugLJVM01LXLzn3GMFiFW4y
HD/fkYbvdxTPErLv3m03YxTqbgnFQUcFUM8ftbGZaOkv8DwmyJFm/JbErX4UmMw1
T4Xp5ayPQQpWzmWrb6jhe01N1ecHgtb+6nU+weIsoVudGZSe1BMF+gxZVOEJf8SA
8ES4VfTpqALpW8EzTLWPsYukjRFqx7JjaSbb3ZMm4/YO9aU3f2a0E6qYr2obDJcc
fVs09pLWofzw1zEi6T7Y4HoUIfGp4oTbHRD3LQTOhAEDz5MmtOq8uXNxgPew5byu
9ItWi1xZ4+1aeAeoQGSZjKp6mnchJx5RXa+J09DWObO1v+RYpsfw1QP3azrJ+QUZ
IMzWRJvkjr9o+sSL/Nu6lelc2SexVvboes+0ZhujgGD6/2IcR9tDSFogVBRr9vGS
QWoLAO46k7sFRuVU8YbZO4QYqBk2x62V3wFDDprH/WF4lGN/e3FmkLdk1q3rs/zb
SLqbK1CJGWEFNjaGT1p0PDh34sEtwnR+sLUVpXp9qe1YCEIzCVU7wOPK49X9zt8B
OxGdRHF9pKEPt8W9qN8utDi+BB26QnD8pZEnuNiIk3N4qaxyVzLeuN8ZnmUq1k7V
fgnuBcIsKXV48u9sNFZgh3c7+acKPrihzdPFlsmygcJl42h8JsMRz7dTpFrOiv2K
PcVB62ie0EI54pNBVIIBBifXCtb3koyf5rmtcYp+hjTRig/TENnVkK8t8KMCKOjt
fD3pyS7LKP82MHEEMFARahPp9ApD0yEgA3ZQ2B0WbEfSZjkoGioxvVI4QOn2ShbI
IoU0y7fLQa+bRt0Tm36m1ISdA5fSRjla1xyNsvgdMYfv7Gdebfi7ye7+mNZUrAw0
B9s/U3CuvxVOrU6uv2Th5dVFZ5rk2C+Q9fFUGAVq5EtAgMWY1sM+kneueUFihIaw
bucl4nZra17owCOHyeXCgV3okGILuIxnc7YGX776UoViRrzkvyGGtztjI+T7/deP
kS6n5xRMlOWAWZjqo8EwgWP798HNAggMBPjKe6cMKQ23vfg/aofVRQEtBzp0rkaF
tSMEs/3tMXkCLLjjNkWtWhIuLV/diuErJqAMtLGB9r0CWE3B+jieuNKbaCDOoM2m
rstLUB6qaMbMC+QlIHWLVhxzxLdlnlCUFIzzJOf10C93F7yeXFWlE910isT5uE+h
ZVhq5KhALtRXK6oHn7i6UTB3W7F/hiSpTDKILTEKFBveTGF+7keGok10BnWRFlVV
TEQ/CL2ulWt3xbhXnFtI0mUfL8o/wyg9O5frbI7adHzD9Sl+JNdXYkhgKgRp+O98
yks7XaJht5Htd1dByT1cY0tlkVaFhxL/yMx75YTAy5RgYnLJQjgi0HTrEcaO8daS
y3ae3VHFIVcTKpQ3ggw6qldk4FrwbCG+brTl8tPcoCJFwsGTvaPTb/BBr/YJARWz
sETNLn4qEACArfrqL2Kawh1BZ3nOzLU97SHcP7WmuKCa6ODJdj4TCZPnPH4JYS1O
BEDpaiHAFTSkEkS28n+bwBjEi0Qbhaj4iIEhZVAoqd8CqpYSnNBFU3DN4m3xS+b1
NjeKH7my2U8dBepX7WA+LodMvKBMUiowZSJU0oK/+2awTj3FLRDabOlAI3LgzI2c
dC0h7fj9d5HU0ymdoTXYMxkyzUrxW8s+gC6NvYZnJ3gRxWGRFg7qv6VUKmOwkrCr
FrFPcNZYeAe239uT9dcxIK34grySo8SR7E49611QpidDXmB1OeV89DYGebtBny2W
oeUL6z1BUDvASM5FCMq6vbEPfVz+9bvxGWxvfOwm+O9ngsuDz4PnyRxaYIZDh7Fu
dlbYpo1t1XrXPflIV9WRat5fpXLxPDxEOnPGlZn5j9NE7opLzxwXfIoFMu471WBA
pYYG7ZfhTFSxbZCmUk1vbRHamjT86zUBH4FzLMLvnhwLIXScFuXhUcWExDjsSEpx
gOtRU/NUZj22ggwVaq/qpNWNrmrZ4T4smtmEz+VdQFXmeHBDF1yiuHUV9k6E29qj
8OGtzb/7ERQ/57zrU/60BzlGy3CRxijyGAz+h1ZTBYx7rcarI+LYv6l6S0HrtDV7
qef7QM2eoLFo4fOoHOZsWuC8gQo7jsW4Q9G/gfdaZSQVRSloufhwFFteWjaevVu/
SV6/O8KNn3ba30tRYgB+9EzOqlZeag6aH9264pxvl3+TPa74vbTNUpkTx433376o
lLZUb6bkHvmXr4ZPilyCzYQEoqN4DTmZBM4rgvB7rzCYTnimQjWIppEl+daIuERn
Pq5JCKYwl6ZoaQzrm2hOotud9ERT6KT3W6hoM7fzh8lZ8/tSG8t6opSgpODbIcrm
mgB3sWdFxRBkBxwYASFl8wRYBDdPIgpfBSIq4HtNSkx/inZHY/6JJ4x61FTuv7rG
SGDYpPTPVhq79xS313S5sOE+arC6seIKg/BuvIpRN95U62g5IkeouNNJ3NTbrw4W
oGTuPbu7osfrIxufbZiEY3D9bqioJjKKx3URTUFO9IKO7YB/vegRGvKxIqzeeA2e
pWqL7NnFRdc/K4ju7XyxKVBD6luvr86UizIiPK6GfK9UmuTRfkED8U99CHfCbzvw
umHDcm8Cmfn66MSqR5NqwNBYlw6tTeDw9OewpYRA7k/mv4ix9PkzVWRs+TwbezDG
rTrmbbAtDIHeE8PWjEP3b/DIfcvKYirbyOxtVtmLOsBOEAea93QD1cMLzz+WKRMj
yf/b/Vpwo+NYHZdlrcsbwpmlw9/ZuYn7wd/cBgZFMds57yY9fQSEYiq2KdkDHQm3
XyJPkkg7rzsoVoS7qyeGtpxqM1g05RFC819y4VP0xD/9e+JvB3PWZjtRjqKK55+Y
3pSmho0JwSAEG2KKCYj6TbQfq8lLgSt58a5dHFYxpbs5D0eXUW9U87b2e5Cxr9yt
vThzandTgWg9F84Jmpt1QI/3xpl7LvHuKSsDnu65COa+24qbbNffvtKcMfA2hxMR
PHcXT5xofgtMNy6YGhZSiTqP4jHQvJ6O0Cr9XsAHzIi8gBK9HxKpVr/LzNBr++t1
H1oLEMRUVGTlF944fiWbmgN2R0GB5oHiiWh2t9g1O8GbqC1ntD4luKwIvQ1MbaEx
F9Yd1BosiepPIFpevdzTa7EIrkf6g3W5p8FK6OiZXf2fpW/M1SYtq3rAzDJ/Z35v
KvEWDCZsZf5YkCnRPFprCHqg0kgU2xY1k7gNk3zXXxqL3Q8neDkcxqP9jEy+wu89
fK+WogiU58RU/4lg8jyEGWKmA7OKxfp6/EuiG0ZdSgbptZYW/xUTp4IvYYB+MFy5
3s6CEmnVG8RBssLO3W0pVwSEMYDgF/hfdrVmYFQ69j+kOsqtlGZwNlaUZ4tf748Z
0tlzBQIL6fnvHl6re09QIaSr0JsxzwB8fG1koYKI9CzeM6YNihKnOzRCabw++cnS
oZKfdpW0gVJ2PVbnjn5iTNbeDACqh/L447lapGqEIAxGeso4yyu4gaH4VK4uuKD/
S2KmaFEejOPsnwqG0Gj+1UMBd0L5/ZXfGeZVIeSShH7en4xz2ahhY9j6iK8arPvm
bFuv/lEjEBZBA5QFGKYNwJJFPjAFuFtKfMdGc82/7pBYCDq09dIGFWC3uMo5tDjw
9D+ExdWzyMEJ+/mSqsAqZMRzYG/nEsZammWyvFsaQKeUeCKxr42m1RM6A5mLQdtS
HeHg6FJ64CKECzQ39H+rib7zdVfemOyW9pS65mx+bY+pQG8RPByurJ0Kyp+sWzY0
NJrX22ecKcqRfi+EO9Fhz9Et2gBXecClvVBD9ZBsrYGDdRGIffrgj2DQRCv+gVkd
SYBb9wzIHQ+PSMivNQgQyPCk9LMlJNIFgCOW9NGpMwnHEAak3b1T4U0r2lpqnXn8
VUKK1cGDo6/FDvcJfOKEXWWhMya8/9mm2QgZyOZNw/ZjwHLed4XI8eegC4Iq4h8S
ryIX8cLQJnvAjbd47rtOBznx9KPpgRrWVx4SEunv/ZDNx9cappdQNt1C+X8YAcjf
CXvCyvPl8QRW3qu4hLGReWVyWitrxtEBFGfeR1zfG/V7N8jFvMm1NtWL1P9TVvSE
WLgo7lS6/DHSgegihn4BBWoDD961/DKt1ywECT79SbWRzLF+axh9PbC4cyu02S6V
bjHw0yOgOvN9x31wqMOPWEYd6PXywNA21G7vH1fd71wx8AOUajd2FOhhMjRbygP4
m0Jx8Sdz1b09i5SiKD6abLN5AbFbq3n+Lyb08VDAbtgkz2PMFa718rrQZhU4fgRT
IE9BqoQ0uUOqfr8vKKk8IVIHWhaT04pOUo8lTukuJlfJGiZWd+b8+JnldXrcQs3F
IlnaOee0iqIqNkARTE5Iwa5zAFfjk00CNpveBHi47Wd2BDk9olMdwVvLNBaaHUbX
tcv0db0NA1hKiY41X3NolNArS606uENoO7praH+fZyX1HibwaZsJbUCb2NNvyWbA
jtufG+VtZFo8Ny/rFO5wq5l41SkNgVf0hBo+KA0e5F0fuXnYAttB49qGS9CLrEIS
1Q0THuubVDl+vNPxFaDc3h6ga3S0wO74N8V5yQ2QvYdsc/sgFsipWY6rW1eRPCDi
1y+x17euvcapvXZW15p3BymlGoBMu8Lz0w96FQlMZ/xZdFerT3abBP/iOnfA3iBD
/iTwxXUg260mSuo2HdQqg/WhdK7ObgibHAidNfLhST7uYFUjPlWa8kCoBcmy0efn
+EkA35mved1VZzqLumPwHnbhKg/4yQHUGfnCq0xf7FQs9sfxGV7iegwMo6UOSg0D
oxMoqET8ahEM14LfKSk909SsBZAWBEjBdu4m9da5s/U1lZPxnOkC0pjOPN31NYQX
5K2rb5c2wgXOLJAaGAq/F8Do2kb58YdB7th8OUBNhS+ioi1x3JZ2WjEt71lbJ6dy
qwH+j6ANcITERwlUJferIBMK4CSwdN4RO5Mw1aYMBNZQ9es/2sgDfIitxZ0vMghR
0+9rq2DXZMC3Np7URvhBnFQlXyTVOPraacdsy7W08A6zBF5yxBL99kA8xP5C6a6O
WFRHfhujK5957nZC3+ceZ7AX6nifEVVtILDpMEKLXZlSZAm/ullxC2XmltDyGnUP
NseuQgODNaFa4PUe6dosea8EjOxr+9oIXR50Ob7xqKY2S15QOuTg0KJVsW7ad2tn
FkyLfMLvIlMnXaZQj4d9EF3NSaMP3Qc3RJ5jY6ju0Td0bUJszdTzTPsY2O5DTs3z
Kc1ufrZe16cdqR2ZDcNPmy4Ww0lg01Ky7PJBJngzTDWmnWyMipvohnr5rLngSolS
OakqplxgSky4ei27GNgyY62FY9MF+bsaKNHAxdkUlT4dylWWzLfAwoRAGehtjKj3
ejrq7u1roFjwQltl1alaw30RnzTcJTC39wuQMs5KgfnjFwq6lEL0Do9RLWyxKSj9
17o88xM1kAdQa8UjWiTQhthb5CI4RVT5IYNXdEgyrKuz7juq52UBHgBm3w6Bj0fq
mwSL5Uv8qagwUSb8AyH+Az7N77/PvYB43eVzmK7z15guVGdaHiSdRUCxnceafpUX
s7os4fNJRw4SlOVYzWZs6u/z3FZO9bE+e7w/8Xf8n/vY1lOd2YplXHC5hldxm9Ro
i5LXQcPKaUe4Sg3z0LVfLTcW87HqT01WUh7RnOlSU00a37942sF8PCbH8QtJPDK2
Bzr2RbZ2dXrJwNelzEtwLhmip/G0/4G4EhTYiWk21kvXpTtcpCaJnCGBZQ2Oto2X
utSRadi8i87ufeoo7d16aqkCsdIpdyPXUvF9CXK0UZkQHcsvGl/v7K7q67P8iPAc
q/7s/cIQhUFsoyiOBkSoTTSafQGgXpB2XJq0ewkK4BGKm980VfJdB87SQE4UXtxC
iUvKKKKtT2S5ZcXD57YWV1R9poVeTQ8yyX4oggO64nrurydiV9zZZE1V1CX47ELz
9zEhY+ZaD3Yu1oBAfm+d5cPmuJmZ54U9FZ3WP794HWQV8FhZQ+cSXN3XH4sqaWHp
MhfOBn73xfoBkXESnIfcWggJ8TCj9qLPsIcIX4SImoeH2pUnGxNpz0EDdnJ4rkZi
bfWCO74rHPdeTrpLKjovHh3d1VHAMuPU37hjTk+qw/4nBXLVqvKyUSkSRMmksHr8
MFywr4w6ZTFmzYUdPk/LIdHPtU4toEOFuPF49glcltyoG8MRgnSv8kw7oJmx4+2t
KzHHPj8lirtq0Sfua+UnmrQJQzZcyyLGlje9sw7Mr2rAsyT8J4eUZWAfCc5yFOPX
iNb3TblbtDHUdAvPYC/wmbxiYlg5KbRSMBPMX8NYs8d1aSkg2tJF9h1li/E2Srh+
AjzySNIu4gHYaqw9dLWzqMrf3aZM+5/+pj2HICIBljDEKMYUdpFEdoHuRc4MoA5O
BMaK3VedLIBE/MSlFzT+e9pBI/ZJl1u3/Ig8FJ6Czsm8ESY4PTYgc0HuK7ToLkk/
BsJ8lLh1TmT+3pn+Es3sZ+1A4acEnH7Mw3SL9tBXOpq/ylF3C0Em55PieXQ2Z5/m
4A9W+Unf5NwcCsAKPMiDOEnYp2osvtEMGn7gun7WO10HJDWnz37gFitRrVl/Qi2n
1FfWlC7fBf/yPadifVmmHYcNWx4M990E1iz9X8n2LErEHrnS5XIjjaRPwpOU40Kj
AVyHrRU84c2W/h2kD0kSuP4oP0SOJf+xxYYMK6mpnmY9w83viAtXJLvRuX3NBEG2
1WD/FF9wBuHc6Wq2n/AR26lfJLFGMPKNEd6GrvpWasz870vj37nMAz+RV3Tfiilm
+vNMJIYZwCjIlo5cxPLAFnPCqWf0+LdGXj2KXMK5sqWc3Duurla3+9BPdeYcl6fx
u7QPMGT3QAk/2h+DqrIziawpsnjOhdWbxIxk/E4NO3uLa6lmNjlsZpBotecobl8B
FUmfN9Hzgnnvd+IFQEaAkHL8WhfQSs+2tEqQTnxF2R76+6hG/u+VksYY7iOsMXmA
n9jFCa7724pMFpnCrFQTufb0Gl5z3rWy2fH8PEV4rjzMiofanLDTdxfQzIf2Ktte
9r5NMLKmOzoWTUnfHDYbGGY1gUIv+noh8Ard354Et2PaKnmbfiFdpFCo4CKDc/+d
pS/Z/nCYlQDXvGGThjjbehy5yzQssRFzw7YDz6GKPxc9HH27gxaZ6hFXFi6F5MzP
erUG4JHuskUo6ow+VPa/ezHSkGFe4Jkq3gspCFFxjZ5p9xJgN5MW5IzLAvB2luN7
w1w0OOoS5rr8lX53xigV1AS9/6lnzHzlXRNCjAeu/SgzQpLfmTk4usc7saxUfc5t
V1yNj79hdeyBtBRD5vTDUoIvP0ylGLzKnEixi/CvvoQI21/8TRFCdH9shjJetbxX
MqVkdNSuyWKqJ/3SHbDwS97ekIvbWWJEzYBzjOpia9iGvBcDEM1RXMwOS+JrSNgH
S5EZLVbRHwKV62QFU1E7UQR8innGlw4+SAr+yq0KWxupdmIXHYtJThiWj1UXulDf
8UWSbZOAuHJ6OPZELoKyScGjEakWvS0BMp/T2tLBmfOs1AM/UNp26Jm2pq6FFZdj
fVq/G+Vt4ZphK0y96JfO1+po4QhDVYSsEFRSbE1W0MZJ2Ed4lcj+WTVcl7NMBFAs
/Z+ZtsHy50yhaKxbs7+dB5KLUVC8oriER5jJrm5xOrBpEG2wCHy8fTvlkf/QTk28
UUOVGjhTOuo0MwElqvz3nJKSAWPFwqQoDWFAOk1tRvFq5mpebEhlREYrWQY8/Q9o
yVqP9yeD0kWr9MOsJ2RQ16fiAWmZCE1xqvgLJ1VgIMH5jsjEcFP3qCN78zRNMdgp
khyrr7zhpvBMsvpZFHBpA00n81EpyvcHV1rd23I4bpf96sCzYiaiw5XvoZr6GSHi
tja4uzqb8BZ5DU2T0QBFOEpIthwV5rH0bgJWi0th4ShZGPNcIRs/EbkOlGqJW0xz
zTHMLtZXkwgEfbrx7lPA6awyzqRgs+TZRPitPNQWNJzkImIDIWL0v0Ck+3+JATbw
mNPfKMzyAUwssaCMn/Po1Bz0+b1aCvm/Ro5ah0Bp88LadUJVrw8xkMwyS4K0Csh8
K7f2YWDvt8MR7DwitO2lPfIAnR2FlLj86JzXeA5EZo2OE1Kw8/SClKUCDew1eIQl
lawDh4J+62yRIZhJ0LEll6ujmuKh5pI87dkJwEtWT4uMX8d+sMc2QrNjsmwEWZHx
uWgmTuLxVuf9ZGPok+XN+RBpOfBwRPeieAAFmuEoywOP0i6pBs0aIcsG5tMExtw6
RwHLcAq1+0kePDV9FIZpWopu0g6TY8F0DOB49F9OSBkim++1IAmrDS+8RPgC2NBH
w+PhEyXf0znG2r9WHqvwyupwzTeOJansld5QqVLoLfkTDh4JWB0StpITmbDnLXzl
MgIeURyvIoylyWJ92PyYCWo6BVty3C3k3InQWc/BF/WAKimN72VlaWdquw9+Y3+j
lZ9qYO3YW9XxODKREoB4UqBX1dwm4pC/h4Hwg7u/np5LPDdZ4HLk/9UzfsIhRLvc
CwYJudkESzQclOQvFEBLr2gsBm+KPXaWsJbVoy/r9ctheiXqIXF4vIZbPK0vvVYo
JfiQW2f75juwZ9bl1DwEMQlrRkalNauUyvDzm5sUPMWcfUYlN0I6b6+aALS0ltCc
Oi+lqiqMsnN4xaYPiHdmMzTSxKKYoctwNLb9I7h3rGHMNNsS7WkOW6LB1J8ZNRWv
dg4uFKnfqzGnrKjhrcED3o3IJCUoF8ELfdD2We3xrQendJw9zIyKwm85sGzPV/0F
Re2A7/Vfy094/pAklYmE0L/Ynx2OtFICLI97deAEVw+Dm8GZxwsbROGQ0vLeYIjm
i9df8Wa8AZpl6SonaHE/qE5r52gmxkxC7HNvv55zmynxGYXMRYsfadKePiAmHdpp
HxQVesco1X9LfpQgdVhUV0nxzFaYKGPnqXnQN1FFR0I4UsLM0mLkjHdmLFIr2MlO
s9Jjs0H29wrFPpqE4IrgLB8RorDJgz4HG6MdnvblWsKl2/epr2DzIrQ1YZ85P3M+
KIRlQenS9uZSL7xZ0a3S7ANIHFY4FS33CxogbWsEgF6PK97NJrK1gSUtLnRHHmTK
PknsqW8IimNSfXvPRZDbYHOSFpUaFi1iH1q+DAwe5KU1BQa1KlQE97qaW2vATxRu
vmbUXOsbuWvUewHubSyFWv9Ic81Vb9lztj4LJKFDanyPpQEnN289TnMm5xgfe2HB
3NrPvrxWhEmTK1q7aPqdRruBKJ20dUcEKkH6f3usBa6G1xVZwa2VONiXcc2aOM92
5C/vfcYrV8PhVmXGJVACY/wdk2RdEvkX65Fn5QvPEHR61LHzUrQUjvLudWEcvhKN
nBFnCyskMhS0LLhUD7uq3c9XfVEWjI2NwRSZcOQD5W2Jx2OH/466JN716Du68iWH
o0Y6Uo2pRGr2kxcXFFv65bSztc1k00Ae7XDNxluz1aszQaV7A79OxjjXKKD37aCF
q7A1AlRnaEWOF9JdX5CEqDTP5f6PFJMkX5iruJFaypkT99wgmKDvGyPkJhQX/NR/
FVP2yUN9M4RBunjzG8t6EtV+/NUwtNGwhRqdVKuSr7ofXiJc5zDyIdWv2o4YVrzW
4RYzXf/OEl9vWt8BFPMYT5qf52H961HEVreljoUotKoaDu3G54VQKV2Dg52QSpjV
I/2kr1kmJ9jjpq9rTECVLe/PnqyxaYkJLwHSBoLTbQ36SKMtrYd6e9OM+N0GhdVK
EsDo8EKd28mPvE3IksMevvliv+g2uHFGXVEDXBgkwMgHroxS3Q08ixymVeXHyljp
NyGsy/hM6H6gdo2m1N1O/sr5Z9A5M5snACptZOk6CdjiPyE9CentMdKqtDbD5w4i
jfpHSM4l0UrOGQeyp2oUxQpbtG590yN4UnNxohB8cglutILgySDKDQhI4AhWpUEz
ZTTK7FjlxkMB6veaqcJA5mQMXH1QYIfIuWohzUPjsKgu53KfpU0gYEGqCyMZDB0J
3OP45nVCSEKfDB4dSLMFXwGX9xikLABDbDJ9Zo66B6k4dDLofbpInAmXEHvgQ3m6
ZpUuLSwP9LseSlKMwQQb3ibK1vH54L2NBbk6l83wiGCUZTVXO6mdBRylpuo9p8JK
cM7ZRagk+QPWhU8vRN+8+/sPZnGx/aWr/y8cV5sgdyh0qleaqFyvNL1a1DyrILiB
mBlu+WfXhfpArKqO2s801fYe1Ppj3OMS4D7py/lzFHnAq/R+k1Ym41HKA7ow96A5
L0h23Uls7N0zsVARxSIwRGIULAnzvN0EeCJ2tmeRTHzBO0i6ppCV2BNieJcDQKku
+U/n7ZLsfjf7WllT8mx96MUPzIz2IQWQElEQ8U/hAKqN5jh7nU2tJNeGIYJeTx7E
3fWDkWHpLHN3EDBVvfbR/tlQ650biQB7K9kdxPxbX77JSQ8pMusqFy3iS2x5nWva
xY9aGomruDMJbyLs6mz7LrPMjjj3fqcKHb3MB1YKj95u2TNXOQWO4DGA37LkfAaM
5LINiX1oMTZvAzzwQ2OvNjOTPQeYmSp8mSx0NDZcM16AtjvmPIJed7Ouk8SFBoF+
qicGEOaY2HtxMJda/eUgtcv9WPsjmarkySUQyGztOLOCbhSz49ZD25pGo/Xl4zt1
sE+DePc4XbG4zGu5gDpyf/lDDrkNMjebFb3J5EQDStDDgAdNRldqnOPvtphXoLLM
8GRlZaXZxB+olvrbNlXI8P2QEeHP70w3FfaQdWlZoIUl5kmjRxcwcr+culZIxeKe
drbZPG3eTT1C89J5pKuVC3KHTE3ai2/T+bDs1ShQQlDkMocUO/3lst2K+DVwcoT7
UMS/6+YCXgmfChh0e93E763w6GEtMoyIVhrKq1mp8bcxL/pzyiWVXzGt2MrloLvD
oioY9u891nAtQpxDWRsgV2NSsVVm5C/7N72dIt+IR9abXcPmZVnLkDQbD2rEI3kD
ray4t3eLq9mmVuSMAOouTWo/HyzftKoiHi7WZ7mrYdJBc0VC84A5KhXoFbOQGp2F
1CdpudqUdGnLILF19qy1FC60Tb29lm3cABqHSN+DgntGwaib2U0mLZ2+qJ2q0Nmd
+tQgqIqJWXbajgylqqjbwcohHgbkUJ6MNL0JNIyIu5Tb5ixMxEVKglwT6EEdY5xp
M19VnrM5mLAec8vI39soP7H5Hjiktn+MphNbDnVbcw5wiTzOZyXpSny4A3ldrMlA
IUEL9IsQ8DphsQ1Hjxj971z96P6+XVMe5HADe8LNl4adXuqz0Rve4c2Uky5qtuwm
QPrNFOAM1l6yIfrZzs/SpSwdW6oGdhfXfxfP6A+xyzZjnb9U1SmmTe02fxDLd3m1
HW8HxCpZk2eLbVKYpjQGE+PwTmmoaYJiJkNT9SLpSnj5wv7iprFrabB7kVUWDRPz
qibz7lDsErOmacMv72B5aQ8Ae5MQlespjTgmkh1wYAG4LVPCS3e9s5VHE68cFYdq
W0K7cSn8t1aa/CSAn9lASJL6ponjnK78bHAwswaoKfxnLMJUjV+F+AnqHCHppJ/P
2H3IzWwE/bLDgD+F6+8zZDqTx3Gom+SkC41EQXKU/VSKPPsG08H1MoKjttKpn9uN
+/P59GaA1vB0YEjm7vwQcf+2F5r/z9xWsweuXedkJbX0IW6tfW0kghKKetA40JRF
zvKr42/SR1zSdXx/XZ8CR0LWlD+68w9EjefgaNAE5zjmdlONs30EGPYROE2yvXdq
STVJsIl/MR8BEIA9VF71a+piVDLgrlQ3xQVlXcdVoP1IaD4m5UgCK0EdSIIjWwwi
9iec15vqrT6rINZLOQtX9t79drTUm/t1MpYNk6VsV0BCmacQSR7j298zwunrUKZ6
y1pQCRAKxpZGFeDr0AkhsWPdpOj+bfV6JrWUJ9QVIEwjnHMT1JxLLN0gcQqJ86O3
QjDZ4fyO/K6sF4uLb9E87uIsvhE5LOhtj88efZRuKTynQHUXn/VRzOb7jtp6qrx8
uXNMOCGnZeVolW9YvTXjWYde3SH/SnmAjfiIRgWzsT77gSSCsyXYbcJ1DxZu9ZRq
H2x0N0mtfcfpFX4ILQCu9BMJCtAAUkm3HOpreiae0RKoHglz9eQoaQZ7YGEMwPIE
gczCrPMbpscEsm1IC/9esVnyvdLWt5hO4Yp4t5Py5sF2RL7yPvSPu7FppnKzdtn7
zY9qSRW9LdFnKFJzfz4lfVCiuB0YYlTPwo0XHgNG914q+BGR99LdqC4mueI8ktwU
tn/B79zcXgqQn1bKkLSl/mweCxEwfm6izFnbc/k8/Ib21m5gPWwURBHZHfvXA3d3
FmEbrxJexxEEoua2Nj1y9QyhvA9zJXFy0GFT1WjB4e8fDOUvHwnRHPAR1g6jBnMQ
R71GFo80ImjyW4qzJsIdsKdQjft8X90OPgZULT/EIv47EsoQLnUYC1pvxo9/RDdL
BBqA0xYXQqEBRZALXOHQLIY779RunGFV3NiE2ot4GKQp5RrIBPBTlzy2CziQKI4W
4iUTQEzl2g+w3uDnsAc86kCitKwktm5XetTdtRo5hNCjVzveSSSWeVAoKFdRn6Rl
CtMXKnicYX9sfN7dkKCapgwpAsns+V1lk6ShSAiITATvXHsOB+0hSfIt5xwvfQI8
2KPLey/yb6VPGEWfKnB1Kp/0/vgvdlUGk7/nswGmo0z4CyFD3l5snlhHvRpMeNdu
PHRVUC2s3mqdi+tyawiL3kRWVA0KAoqU8XGttmBCR44tIgYH7rGW4CRvmKA1tKo5
rQuhbW4IToYmbnbPWBDKFqC6Iol/29/EipbJtIItQJY958dIMY/XYuTXfgZkJwWE
rZR4qEyeHJ4h4HgS50Ia3NH5tmdmwYuYHPUslHbA5pkVmYSNWGDZdy553sgB2UdO
CY5TwpuJKa+hNc7vQ7bfSmOhb3m1ETA93hc5AOSrARDr7XPZCRS6f/RsqY7y+2f8
4LoTxU1BIS1uQJHSqkUTNH7Qlp3fnqV/zhBRriKPHW+F34Lmh4J9wX/5xIc/8nWr
20iEPn/9b1aXAXeYJWw6l14GrdsECjvcx4p85UqpB9EjEmQHpW7xQcJz6fOJkbxj
J/aKdT2XPWDiwBKcKvMlhb0CEKqIkIp6gh6CuV6OzUudr7mvp2Ji/IWjNjt1/Mio
etmL3YiOvRW4qFzG9cDqENWCd3aQ1TIyTc/iy8BiLoKswlRGxox2liLr9HTpF8qz
OreckJHWQlHPSk8s44p76bt5A3F7IKaAP7elI1FyjwFU0yVNIo9DCebwq4dndpSE
+VyoOdwe9/jHVV8+tUOI6EitDpASOuJtDgoHvIRr1fgLdfB44G0wWbtqqhR3Q9hY
yrSSp9aLQO++XTz3PmNmcK1a6cSSv0DihG4222+am+GHFxAu2YER2fAXtkdt5HWb
2FO7Jcvxm8g7rzDKM9ftRQ3rtDKkymlnpk4soxlZLdkLV01tuUItget2QHBUazXS
jzuYqqX9wnK2eV1XgyBWKWQ2b6j11LCdtzARHsE4yZ7GGjKRBUHMBGXq2BfjP+MJ
2qx0/fNWCsKKiaUCZZtGUVbx84M3piV4zpC+R5jyO15n+4toP8N+cICgNwdWKZDn
gFvrp3rucq+WlTsAwmysfMVK7YYKty9GgfA8/b6R+A3U+0KsYst0FdBmxYpITwPP
rptV7a73it/cxv/pYrIZNXqLoQ2YqRJkcI24pvuAi8ZYfKs6ChLZBsEkT59p58oH
hmp4s0Onfh51i+ZikV9BAP+3eVM1/oEg1tfYaickQpHJWusnikSsx0LuPJEz1Xg9
a7KL/AtWLBWdq6fc2vWjwEgK7dkkroetgHUzAOMa/v0uCLAoYtd7aWyGAL2mIerH
yCkn+OoaVFjfvmK4fiUxMHZUVTVPBO2P+VxEmjYxTbm2PL3VAuGwxYVh2JGf07ZT
mj6rMa5Om8BE1Ty8N/tUSmHCHsmXVk9qYIZQ9SgQ71y+Nzr+m+sj/eU2QUDArqpY
MJs1BLWp5KlfCuZaexNGTVbhP7tLdLQfC+grAHg3iLlcDz2PiiLxzoqSD6rGu+z/
vkR9A6LciWfMQ+MiHmwP33cWViujjrzT1xf3dt4gFuYkyfQkjUCOUICh9ivMpUJV
zMs1e543DlVkNPFCgLPWqaKS8N44Apb4prqAUgyblIFJqGr/0ELZW8bKGCqXbv93
SsJPjEk8Egzk3r43UQ/835HoEhRYqiEl9F/H0N1q8/v5oPLzCYXDEfYCIGQFsoHm
gYUsDFBYaHzkuT00n/SZlAQfJLwVw28xn9mlgDEKH8551vff5uGZu4b0Ob1yu7OC
hVtCngSyolx7bwdlymq0eUf5u8zX8zFgIVt10FYPNwM96RHxOEmHo50rS8BrGF1s
FjI2ScK0MhMsaEipskB8F2gaYS2Z0H/+XwubYd/KqJ4MUETStGR8a7MP1wEw55aG
33WPd0uRboGnyIMJDPONwW1lxpfhlBbCusaT2ek2tjt+TyTELVpTqDuFSw1j3jjw
MsT1/kQyOHAwaRBjk2EwWbZC89P+2Igpc2DA9lroCZLMoOFDtvt/Z9T2rhQRbTL1
obCZqHAaJsptOlejOqn1gTN1WoZ+HbnR2wRuG+nn8OezLetu66fZfepaW7oP6nFf
7JCt2LE9T9cdITf0xofAM47pLYrtEn7RRLUGFMkDnpxtUEj0ovufUZCrRkRlAb4x
wTcLt74izL3S3mOh3t3Xjcm5cJe2ekIY8VbbGxX64xyijjkkRKkyx6OWx03vA8Xg
+W6e74MLd4U2yy8GrE2iMmsvPB0qCICaMy06RnUJAoPp9g3TuL20e4wCGYFW9OLb
oaCuFqaWLxWQSy4Z2eVqZpBcxDhqkk2/ppKrJGA94UdP8/vN8pXlQW1RmGdzr30s
RuzZYyNTLdcqZFbZf2uZ/Ub0vOyHa0XeXmLPvH7UXBUZCG98gfPQF+ELhusPaOOp
HEXKhIiIgrGmLOXPnOuaaHI3mnw9UQJQaZuU23WkBmk5bimrOMVpHtyeQiXEkR5n
X1maYx0YFQwBotnI59u7cd8VCEHH0wxWcqD7lzuSa6HK3K6fPmpZZ/ONqs8ewOWp
1hAtohYvD+S1UG6fRiVqHBjou3RwhC2Z9ZHmX7s5SpciK7kMfB3xEcHJcAlNH3vp
MxlK8lwwpaxF3I6oGi6jCpzDhQn1UMqgMsVdJU4Ej+YqX6yBSnwC/DDcB0aUHgWV
fVIl5k5dFNSmzv3B03n5oLxT7jo2UjAM5VlH6BPUP2pZfIMI6rAxMlbsyb9IVL8L
KpmUfk5Y2p4DnCwp/2bM5fdbmnC4Lo96WQy38FWkj+vSPY0guz/ELVdGleOqc9F2
a1ygFLprlHe+wQ1jj9+YC/M6niLgz3Dgh5BOyKAZQPixUp13eeah+V5upb5d7Fn6
t4PSkZ3MG+Tb2emTSGi+ruANpNMHzs6Zg/i89gNvr94S67chgmtLSWrvonyyhCeI
cxZJ+LPdcB4hX39cotZSDVveb6+pbrHBreNQSTFR0K51lM3qIlCd+Y2LyTYAb5GI
n4xVIUT/RZWh2VHjYJLV71eqmj9gnaDqBzm+CiHuH+r3LeemTQHkjOam4KTE+U3i
ARJqHjC9BaZC3Qi9kkQyM3vVrvOz9yzoIj4DyIQyhXPLzcQ0z348cLal+GIFR+67
2c5AEQaKiBURKnicWhVaIw5kwsSzZ7dodomdaRSyi0OIamRB8ppM3pzf70qKNjGv
bK26btM+7//M9ju+w1D7KywbJNtH0Ly9wpZhZfeKVzz5hZ9BqnFZVEgvxDBqqn5k
2e2JLZ4YjYecHwzoykW06vSvdvmwGTi1Qf93mS0ocEjQzUPWZAesRy5N2uR7qFY+
/UG54tXesT/KWJWrsX4aNKg2hGGMqV+Zy0ovkSx6Afk3QhzMm3TGp2fzq9iZX+gC
owOv2x1FasJX5WMUCOpQYRsP4O3Tvk8kt82pmRe985IeP5n8CExH51Rg0uVwZw04
xDSqNpUChtifmclAVxvtzhSgZdo+bDWlXGornOP0C2g7H7Kvmz8n1Nd3VUdV97+b
L3Qos5eeEDF1wgLOrKxwetYzLh8kk4s0cMjZnwoMTMZ/5muhR0kw71RBNyPBbs86
oJsDmO973Jl7Qtp6Jn6nTtTK5ukc1RCjxvfAQy/xsEj9/CWFq0ey5mXafJkxTbD4
qXQDRfWeMASfTpq79rlbLuSjkdHj6GZhwrx9mVHLDZZ2MO+CbTEs+DrMfvlsGup2
MdESaY+xu338AoJwTSjD8O10looKsNqpA3o7ZJJaa2co0/MQOPIoUEj9JJjNEs4y
QPQd4lVewu+ALQ/lcmOpqjm0zxyDOjDp7NiVh+D771lUSpaYw/UOGyYzCR1/DaQH
JNJl0jzmW7uJF+WGvvd74ObxQ5uvTZp6H4WNPx09mp6EEUKuGEv1NGlekTS5dvLy
QBvFUBE66G3yIaf1xbY5UreQ096GltyDoq3RarZ4br/4fzJFvUo2ezkGbdQCdzZG
zTLHLmWgw3Z4pymrhIdWPoDzUWD0akO/GzkVEI3NZyamjZqKXr/rYOQXoGouSv2D
4+ODyhDaXE25ilwtEItDFXLyG3jxX8lYpZuiBNrYoxBHFjGpoq+y73B77RyDAjg9
3xwBnK1tkzLbEzkW+J1JNVC8zhIDlB/B+8fZJNupwZEzJBdMehf3zlC3ztO/xVvo
nhZb7hQFE5LygDQKnvj+l5gPVHAkCqVlEt0JQAXxxAYM+jSO/PWqPTEsIn3dG8jj
XKqZk3uR99LYMa+NE0QRsNgglSaTS8lo/btTeT8jd1qU70lAn1cQUxC/WLyewtZm
j0ah4J5bDNTyM4lObYzOvMvIJX9QkXbPcxLb83W7u/lLRQMnxmi8GqCuHGmkbJ9f
5QxISPG5rz44duRv7MtKUE0L5+TqSMMjlp43sdcYRBqTwad7pU+bPoMgpWFemXiV
PClRAOVFF5butNTERq2vomxxIHIOu3Gb37NW05s/7+zOh2nTjDhRXdJ1FhlUrzrK
SqfE3Z2mAUi0VFHiRiK/pS+vEDJOZbWOkcbrHRDzlTGCtkCao0xJEgbthayHh5PR
WcwnAk1OqwRxzEtNF99CmgX4V4SUEjczhpMhPS31fBeoXRNNxTehm7f0c/sueN0c
APMTBU7Dz8YOEEToDedJeABDQoIxrG8GpOJmLGj+jUbAbRZMFty098MCfQCZsftl
85QZnPvItaKx9AVd8+hXZsLniDKoiRaGRUCnhVIGwZU1gGNaxD+pj+dFnPzp9/ow
pJIxJ37mC9sX89Vy3OA1lRH4xq4YjXgwo32UW4EZldLBGd1qjr7BpKrZ3uVojWda
TxnP9p3VvYACoDxVLoKBsdCk+VrbWuhgFtMuNYXv/KlOLUnpgUDgAxvH3Skej22M
RAqrpm9kjr23WkBBKl5oDjf69SoBJiidAFSp8lVpBmFZSNXD9Y9aEyVvAIhdseIN
asrCvJwSdoe0ED/G1BRnt0foHX/L6zNHKUhcn5BX+ppMK1bSaHjG2y8wrCnG5KNn
B++orUg+G20sYsTtjjFUQwN/cwuSR8sRXMGpBqP5A2pZq/+Eg7B/gYB1Yu8hvL7D
QPZZzXXljcT77DN8iEed5JXnCuVQZJ/F2D/HzgVsFRvAy4CvSD2xLyEWDLsUKfkD
rtXuu+fD1MAhhYdMBwgyfX7S3reTXFO4OjdITcOkcfcB7TlYCOCd5/KAHwiMZoGp
D9Mqn72vdkS0JFnJr5ACGGF32pAUyfkPj/tZWWCHp4Qx43rk5hy4ed4kbjXRQdR9
1YgMpadZ94oLAUXUvxuVi8x5BToi4Yiz+5+vMlb58NeVZIHaNfNb0gPfQqNv0h8K
/9qF3ii9scExjvoq8hXyK7glfR5EUJI9Kuy8Uq8LDidTou4tpUqivvhtyhww/YDm
mgdx9yyekzUZobyp6q/g8Q8Oc7vHO1XQnlTGcfu64S2r3oUkijzU/1xA1UPKsAVl
f3xcUrAcSChzaFz8yOMKI1iY9Bonatpy+9oYiKaAIqSKfgrbjJwrgcONWOVpyLbH
qqGxxqDRn3tHuEW0YoWm3rfc2tZ1ll8B9uDeMP/Q7hy5w4nKtGEEvuesvS6lyFZw
CEOP2I/b0NtwtTKoGoEkqN5NW4K9T9Z2A+skTWjFXtr+Oi2yLjqe56UwBw2mRzyW
TXd7QEEZDm5le5NZnb8LH8sPqiae//FtwUPNepz78TLRM45ises+O/iQhjUE/XkX
5amJQfHLmhqf33UAkd1KctRUIz8wl6tI3SCE7vHnz1ktYq72DdOcEC+O3Z4l+PRF
QXrXH+KQ8xMMxRSFqDyas/bN6vVN7pl3sFSSjBAQ3WWiYedYx++r5GKjK37Zn5+/
3HyRLzNffAoiUjNWTgMAM5BodNETtYJIQYxSD00czLerYm4wOspM60cm3+2kJZwW
dxhJYjgURMu7S6KgHkjd0Pi4O72mZhfYFW9PxIqbx4vkDbEhUPlsU+S7FK5dGt15
SpC6qe2a3vv7UXNsF7wG7JEN+Ffd7koTsZ+t69KS/rmp26zR4pxdl7z8Jedw4gSp
EcwswHHh3Uvlo5NYzQ0pi/qY9e/qkLgdiR8XZjQW90H4pbwgURMYD3xLxoPtfowj
ASbwZtl32ZQUcXe5bIwd4QirDIMqdIXxkVcwxXk5mQPn9o1HeBTMcCqNrVkXZmm1
2mszuXiD5CQzMn8h0N3pkL7ZVLbJfSGSZvzFqBGF+aTZlnPmiULhAG/OkBr10acW
kihUepzkKfSW6pK50WznV/M5NhGbYkIXzv5mDn5gxbxGggsKlIZjWoNN1VK4IxRM
MmzrJUS2BiRvLSqA4KQlrm8aMa6k8Nxm7UBhvmrKoOr5lW+gIJG9aDEb0QQkTRkr
KwTZbqTHtyo4cqFY6VA4uIwu2Ft33p23BK3QlM67T+uhGRz4AU3wWta6AkCA/T3J
VN8UXSFWAyMqB77hkNHJOybbUcypWcZPu8BozTc2eajTwDQQDh5mfJzg/mIeiPV7
DF1+emr4W28b6oghCzdFHTrMMPLGDZ/gqrzFP2cCFJzkuToDJAqU7Jub6C6nJSAp
eZHxTO3neVDqhGb6x6GpZni5Fw/zHMMbCIe53Q3rYgefNKk7kQPtfVhupEJJ4jdj
oaW0hsnNdNd/VNfD3FrftgYJCWXUOuf2TjR/zh/D+ijTTOi1WzKAzS9VO9fG4ohU
t+nud0lF7RJXz2LirSJ+lGTij9+uauHOCkziyXEYHqsJ81ab3ETziz2a8+BmA5Zx
v9QJEQt5RJLAkK8odbZ+O+L3DoLBL6jkUo8oSMo5ueu/8RXcgGoNQsrccBlgz3eS
VFWoWPHOYvGqYg0ZE93XuUtcY4pOgc+p2rRUSV6SPBMqkd9aa+Uf1stBh2QAYx6G
6U+WTJ/FguoHzCxF7iGqpFljhjKy9TA3Fd/6BG0l/eZGGBdZDHvKLZCjVSdHvjqG
Tzo4Rv4USWP+hWFVkdPXLqor/OMdtWP3ySlfngusPeLHSVBHpdftf6QQ+H9EwE4m
ipXz9BmGVWvNUDpkTsaWJ5xAt8D5O4H0AFCDTDwJM+MtusD+Bv70/bLhjaIcL8pe
bmvQxhyjAW5bBvaLZo4MenXLvjmlJWv7XfqVanyWpawtGK3uMZyxZsnhWD/NiOGY
jqhrHe2slAdP2pcl7D9nZQNzdeNdiQfe7NWjwORt2l+UQwzyOmIrwgIKnU3qhC5K
itqiqzZzGzBBui5lU/BA5hVxxenyFz5ah0Y15NWl/3mJCQfUs6oRQaMwbVuryAjq
ClkvDtDe0TDNOUBXsmj4m+G8PhwJjXthUqbpadGta3StvL+Ojctrhka5XIWZP2by
MJC+UCEVsIq7stDthD5A4MzJEWaCBNp3jLH5oKv21y/qvHDOpQS6y98xQxc2/A3e
2XRe0IidFWY/3nvvjmXkVCGqDp3zDpjSPEzot4zFLEUpXRVTc23nb4tkonD3yilQ
gl4mjCszfBgJLmlPZjvYmiMfuKP0MMul14WGbC8w2AvBNtc72n2JdXwraCct8vuK
/lxN54q2oApNrYxsR5DNyxxMOA0DOFBcadnq4RFI2lyePZuPEvtbFtosFWx+DqZq
1qyctvNJzLnzgk9ZWVxorvVoS2EKdR4R2/Out6D7LBDGH/B2dKdoOogOhthDft99
5tV7Y/C2r5XH+szVsvlKGu/KRyYJD3qL+ISw2LEWWrXydTsx96tK1cLedsXE4/X/
ZJqvwiKj1gUIU6kf6aoQGSxYnrU/zrRzpOAEB/ZHshe0ataPVHOkFYiZaZGPQfQI
xn7AsD0EeYKmiKY3eegRMKV4JoanqybaUOADslJDNrULQgf4nikD1TjM3ySDHbUe
BuM/6gBC2TeByghFT5UnOQdhZWkmAQWXAPJGBAA7kp98uC7dPAzOLpxVbDmjm7Nn
isngfQCq6yyHcs5+gt9SqYl4agnx7CMcxcySwC+vz+ndAFk60c0iEqgPvg7F0BdY
EHYeZU9hBh2le3BIn/+qypC0yw5ZMNiRRM4MGoqL0IXXb6SuJbAuA48z3+Kpxu1s
gGQo8Cn05R8GeO4gjJpSb0eyKp5mh1szyDrls0bUDBQcmpTrm/ap8k5rmbiFhedO
boIUURPJrGF8ydR6+W+sH6UvNmTRGw5ahkXx6Z4be9BXBf8jBj7HscMW+Jb90Sfa
W0IO2qM4DiI/zSQGERKga4aEyJ/BJ/t9tWZRO/8WjiUwas/4u62JhFmSSSyNL8eg
LYmap3oP0jNUcjU85cL6VChC0PSGWa+PYYcGeA4CqoS/u7/K87SPyDJcOQjf+aJW
nEyVx0/hmPL9LfmT3p+E2VfY8Drkmwz2p3N6ka36DEuzmb+Ps/OsbeZPp1200M1l
tY5Wlcj5XmzGGoEeRujpbLuc6nkuGwLgNF32ZuPiry5wR57IS+1sikW89iF6oetL
0e4ceR75fpqJanVTF+k98WlHYlu9JQzULt4d65yuCQA35noKma+Tzo1U3VlOliYD
t4HwVx82U91H3v4ilBIUapUaifx5EERlAAVX6GkP8nLMcHpLE4YlJkM58lHh7TDs
bD7zPFz5XiG95z+ETJJI5BUmxPY6MiHCuqj6avBD79w+2rg+R+jVuuLlHPkg33b5
XZWTRWmKBle8bRG0qzMc1H5Lj0GAbspKqVy6w6va+zXRa+52HeL+aXUcwQUTJLjW
WG3XcxbyK8aH95va5b2l0/zazBqBOLxczBoga+en5k4uPtjJPTllmGfDhc3CH70m
Rf9G+RSDFgetut9dFkETJxHfmfBUvxSHA07ezk0qJqVGsRaxEyFfEMjuIzQKbzHR
RaN554FJPUg96ZwYSk66wAHXA/6V4dXDlsA2v8xtPwErpgOsuB0p3dlQquNRdr/m
nWJ8AGbnhIm6zaycJr8YIRJ61qy7ej1tVCLCMmQ0aq+Jcm2gtWGHth97P3CVTDkt
cmVWAkp1re+CtDtp5PJP8prFV+IOx746fLHpRk4USIkvPln5Jll4lgGyQWwS0x1/
k+kgsuaigsNgdaCdSTcA88ZWp5W7cDioW2PWzW1yhgpBUGovynXaCuoQkiTiy/8G
5wxB2Z6BBJ98uXCetttB0LJrA7rcKuzwv7B3b1spuxdhbtl8rrM8b8raVNv8RIlE
Q0hRFlPoV8axVChmovkDqHWtEaJ+iKbFJ4i3QbOe6812NG7/CWtO8SmnAmtyJEQM
af5RO+0WcIStdkC0LH4fmn1v/2JgWRWznZ+iR0fDrAzsTt9hflNUYsQ0DndZL8Zz
C0WO1IkdAgwnvn5doHCbxyeJfTExVCpyh+BW96eOoS+yNVT8Bjb6AgimD9mD7i2x
5tavIf1HfkDsExkQGy5vRbQUae1iResAibLNQd2A+fTHk2aUhneQhB+bRi4X99mg
VaExOo3tRFfd28A2kZEnxKWnGFlqtc4JyroT41i18HD03sVqhVYUdij35U2/QOhI
NawQxGzi+H9CZiehjrnZaEi2uiKPuIiBA64lkfseEhXPv7KcwljVcfdpMAwMoOkq
0e01V/12g1TImp8Kd+ifW89KKLVbgieXg6G4aSu8ti7EzL9O8xdkvJ+Bc6iuk1tR
HDLf6eknAITaKmDSSEVDjmuT4hNqKkvJrZEVRdouO9zJz0zIJLMKCuLnFz11HM79
IEnti920LN4ViC0J+UmkM0YV58IxQm/ivadXYPmuWYVYi40MTAWLlJiFUe1TXZDs
FdptIj8jnE5Eh9fF+XQjiwwKrEe3CXCAOMjA+vrF9euxnMKQCNx+6v43hQHuLniI
PRFj5LOpELSRWsZRjzn1w8KD5kUnv804E5JY+oX7BGWrmBFg5D9IZ03euREPSgyt
hQLXn98YmIQiJE2RLKVA9QMeU366Vxd+45RaPxg87MjgOUPwMt8G8fzB3tvX3qy4
zj59UCd1xhiqiTF4JFGd+uSjqk/ihU/lw1pK1x82cHQ3K8NTeJEYhQV9iHZ0qIhz
fLV37sJzmcRbBGEAcQU6sOvOwrTCc3i/v+jyL1VMaHFeIubeSciqXRbESlxHFV2U
cAoDyQddwDOHJ1U7zXh20Gn2EnDL03VlUdMlNLZDee+hI7DQb92BtLC3JI7yrdhh
Zb8rt+WL+4c8h8Gn5rAz3cQTjgmPZOjaMdOaoWcRCKXviA/TXIxkGdq97N/mKwJc
Opj9771Uq/dDcm9qcbHHqZFzvp1fm5jb2KapLsq7Tbi0oWX4nMUoW9UlAlNGeoC/
yU5KHYS/pF9Lt2VnfMWBmr8j1KAbcY50Br6V62KWgZsadiyru+10KdRXrkgHNTMk
sz8yV1Rd+KbiVdjO8VXlW0swIiEq/VvHdr6JNZd85tRpQvp7G2QKbAV08nSn86ZU
cf3chxOhNnNZauc8d3HtO5odanmK87B5DI/CDfNjc6OfEwfjY1dAxP2tk8dXxZsv
pt6K4Evhv1Lz9YAiyGfYmA+IjFKecnei/4NJtLc3k0IgEYqyxAr33/a/qXjLK+Wj
VuFtpUX1hjZJ2aPeRlq9lHOMUs0w7FHNOlNViLO3FqKwZJrRhguzcscC5V+uiqd+
ijxfqkmGcAkdUuizQTnGwtPvwnj4AP4iGKtUyX/qOsQf7vqtUPafcOhvOseXVDWe
6QmlG0EmguXhqPVgfVYjskXeeqmx26s/e+syJ18YRRNq+EPtwUfBWcAoc6NrpTIH
/CyDUuiTevuDzVWvsKIUCZCa2bR1yicjZ3R/F0L95ERt10xBYvS2lWOrfwthysqM
3r8kh46WEc6K/RALA3G3GP1Vrpm+Bg5uQh/AacuUn+X+ViFlgYlePdnYh5kQTL82
NjhtrpDcwag0KXy3MFNDoh+5sDO7hYRkNaWeZmQLp5S7998eLzHRUG4Ced2k1DLY
JSjd/4ZXHiqypKGl5QSaSDkuUq2yynu2Fl2bfAoB+KlrsDDT4OTx346Uu/Aisf4K
TJaQ6aJfBnpZhg/yoDB2b9SRuUr9UA0XkJmMy+1N1+UCUjoL+yLwF7imkHSC5KeP
Vm+ocVorKsoIX5u+qDTecW8g87mjNhpyeBwn3esYwEVw2BcNYTZYHTjvi+Y1zsct
iWa4D3/XTQU2NnqtPo2vu0SnXXV7Fjs7eWFBGAzo/CThHZYPEgDsEBH6KYA6FMjX
BqFTneZ5TnQ9ImWmwCE6/DMkEkEyv07hoI4eh1qjbFDtKGWZIEI6ArhFodVSXUS9
IBtBb3xVTfx0Di1+Kuw/D0/T93a+ZaYwCQb+Fp+1qk3KriKajeiM7dDrYOC2mpOx
VhfLg1ktysAq6cnp84L3aMZuTG1qYj1uARV6X0rZr3K8xN4u9C8DEY10XBCstChE
3Adl+f07QzkWtHAgHQebdIW0iN7izX0M/pLgM+BGGVuGbN/hm3rAiBHZC3qTV9uT
wkKyNvXaELHwhRnABmfWlvGqhlfEeJk4BmmB+VK5x5ETVW5OzqYouuzSYW/NCySv
ETQ0h55YqebECvyXOPxflYB+AMa6fQ7zyKDv0AVrhWMmZTQ2NAF5OoIj91SRUdeC
kGzUId0M8UlxrSEN9JLtPgfnbt6ePJNVh+deAZNo+KP7A5hgD4iwAF8kYtttILHc
YAIrKCutlORHdNAd+azx91E0HOqfBadEBKZnF3o1ePC1Mjstj6Qsj5pU5uDfZzBd
rp7jqW1y/z2zeyb2rJgusjoKvxLXQ2pwlyJj4LBiTmB8cYtklxkhnlVApztTqWJC
LI+Z3EVqNQ2/fHU+4g56do6mG5vj9oFuNXJSKfJsTejRxiQt7keJzfXl3Y0jKAOy
1a8iOxxjCMs9oRcxlCvnWptWiqEoFotW7k+/CC/3txvF6n4+TX/xnZ3bPGaTwb+u
RZv5mNO+VevoHzFreKaeiKr6PAg6wLg/avO68T1GVVDz1uK5nBj4/rhvvwHp7SQ/
2EHVDCbgggFdIkkzZbyUP4vmcmJGDU28ItaH23Nl/Ii2ZFE3GWJata3nnAw6h6Rn
X9MlH8QEha1D9l7E7QN9ZEHyxtSuW3zPd92wmtnvbeWIaNoKN0HTG7w3ulVvxyTq
oyP/xjhP7dL4p7lbLx6BFv4oywNMs4+6gA+bq+oPA24vbeX1gjz13rdKfYsjShYp
YZH5Hc6xJm8ZGt9NlPc9wqrnLr///9lmqJMMzqmc/BKr9oz+LiBkyS3/4uHocbwf
0Ee1sFuqIXeuq7EHrjGPo356+qzKfvfuq2kyO+TuDdh2Hw2Svoz76dxZx1nt1fOP
pw9TnCSsEPcGLPqOZry6/iW3TfrDIQYKvB1n8QecxfYrBo5NMW1kB8aTbLGzbVin
vL0c7yYWhNBc266dbSW6d0/FMbtpngw4IsWVdz4X1OfCsjUv2ODQ7pYhTwX9k7w1
UCtWvbf4om+8XmbK4CQLW1mcaOZYQN0LpHNmPGaYp/i/UF46S5NPaPfFAZuTkSDM
xsOHWnzcwsz7jI4gQ147vTQuHlNBI1ehAvg+SzKknhkPsrZ+vZPtsk7v+csERgB/
fl9BIQonoqCFLug/HGmUx9RTEn4tcI4RsUef8i5jFpl9LuMbC6bD6cGqw9jglvXs
XmLp229KPMjZPNF/orQRTKp8hv6q6151Suk+vqKZsrcPMWX5qBB0Dmxo+gNrXakw
nqK1GhvwZcFw9IMjw4ogSZ1k6BQ+0RcjPPe25HICC086JxM2Fy4DYhoX9ezgOry1
ASTcia5oGkIScKyvo/3h1EeFSyEjSNo66D4pMZhcqwd0fKbOCepyspkps0V4r6WX
QCQ3fo52d1615MZn0SxJRAU6P1oxNEoUdFNhmY5F39WQJGhvkSMMSiVa8iSzOT0n
tOu0G+qA7fxCs3LnRZLWqBojt0T5fuSMOStyJgAkRITsJwz9trM8dJJMjqyTt7GH
7w9FUyveYDJmzQiGUjvoimkl3UeOrJ6YF6xm10GeFUJgIKCARFuGkANgof6iC64v
tbosZxqTeo0F1e49U4WU5Bxm5Rfg3fg58RQruLVC0DHF+nX7nlqlDkQKQt1fsovu
nxhl27qp0VktImd/CAEEPH09fb38/vu0VqpTPajQwSA1YBWJAzTCcEdR75O3KRy4
OiLzZMo1JkcwNW3pwOi7SdTi/saVe5n6bbkaSjowgnqTExr9FXQA9RdB9YzDOcIK
sX15ziF93T0yf8j3pdvNL0vbbfyWJKnQuLuJotNSsJXDK4PwWV+Fx2lTdpkg1PJd
SqQW76GGbnXtHNhpd+THz85mg9cZPsL6Q3/MUVtGRr7O//ddAc6cXOGngmzxZWSs
I5J7/lQ/9AzgRojgwSRvQ5mgWvWgwEbf2LVZE2zsSVNy27UFVd6dppIpgnHvAVKu
A8+cBmrWqhMM87xd47MXqiENGTMxHpHOq56vgLRygVE0GDY7vgNs/2gT4cmvb/yO
/ISlvUycn2XKrrNNrTU0VZQ88EBPz0OTpGSYKprYMFJV1d+LX2ertlD++sKFSu3o
YKNatDruRW1c1SZErjyqEevNdpPJ38nacDtEN5wBKS8CALFqusUAcAPiNKvCzvFI
oK4h3XBzCWskh2Teu0Ycjc9sMtLBpr4zW5vFbuK+VQSOlbO7+Si8CCy5r6nNh0Mt
aDge2QzuuZG1MMAJHuFcBy7xTUvRYVHIOBFki7H1ZA7bQpUmbc3rU0afT0t824cM
c65Om2Y4SZVcBLHFK4hjaJQyQbp80sh4Z0sUhg9jZHHQOvh8/OCkdo9x3z3U5wuN
1DIwTlVxIrvizUz6FRRYo7PGO1b1LdQAmiHEim/BayLwZE1bsqMOXev4GceFCcEp
ZRlRP3HQRTrBBItQbki6MSJ1l8wi4AkP0T4qPZ5bqYwrfhHpsjoAYgamlrT8ZXDx
+4vnPoezs3KFrIwFOUbGdakYZrBn56ARdqQ6bhtxs23PMwqe4uHPwzVlk0S60KdS
p+saUS2kBB6DWsj4Ycdkvik9qW0bwcJNdk3alNsZ/Gf69sygcVWSzOcMJT1fBBCz
LdpiWmDPRwoRAAbFkpJbVu2wxSgNCXXjJyHeheygkYRH/9CwL82x4ofV3jcV1l+M
5kfN7yXoGZ0vG+ywIBbHWsNYes+eVchhVSo9MfXKXM4/VM/Xd6O+2L519zon6OBe
j6XRb7E90XkzLL+JANg8+Kf+hoSrq4qk0xv/QYzN6bQKyIU+um4h1ZY/aRYD/PIn
H3hIRcTaH7cMEaO4FV64v4vm7mh71Uqh7tnCLSZECkvOFLJAHmSuHdGwS+BwbzRN
aqcEqSoMxzBT2cVgyVdK+cFOS3lHfkBfdrB+B8RfGxi2MlwD+aSrRNsqKgjoLTam
q9AR4qRncPXQ893iXrZS6YbxivpvVUFme4LlM02MxWMDAm3l+GrdXMWpF2AZf6F0
AGtTseDLHfT77OUh0Ij3zGfbO538FE08NHrA1kpgS+VOM/RgIEff3ly/HyLgvilv
it6bNL1b4M3N7moHcZxDz6vFnEV4uIOCjvlomI0sP5DNOouq21fu6DzbuovMZIj6
PNDfhtpUV7n+7tZRx+X2ZvNQjJhYX1vT550Mjhx3PDZSVHYaHJirZrBrORq6yOzJ
ssV6A63LlN3mRYHLWIRk1tFbQ2AqhuR9FDptuz0EKKtBjB9zkjD6LPgMiS0Ry6wV
BDr2DMeBn6Q/hdVmdEAHUbRAyaxSLCGSMAceZAKHj55RQqOZ9HSTJwgoylp3jN5t
LFgqhlY2+MC5MCpBBW9Fz37WN2bSuo/UdENNYe2T44tbL4wFvcNwIzq0Hj9KmPo8
BHHXJxNqISDK7XdOh5lBtEG4mkzxRfigfWBMdTxPgYq6DY846Wly7s3TDsosBStS
8z2mP5f4QnwBQz4klSqCIXruqd0WBgDditszW+JK60U8GRmllncoO8B5LtsPnMW/
4R7xosYJwqgK/Opt5Ho1g05TvcYM84PlV1TNp64nxcIoNyZBomExpofs5JP5qb81
OUXbZmQtETfOCPu5oGp3FlnIsQnvVoKxaoKVxC+LmRIu59MZj1EdlbnqDV7+Ke6s
3te4kTTN+GpCx6ar0OgBFQh3Ye6/fJV+bt4/gW3/zMwvo+5JK58QInK2Q4Vcne5Z
kbvWkrePzgEvI+spGdpR+vduP53YlWgeA+0gAHQ/yS+r3J+qiTn4satZDRab77qt
X+OquKZzhQm9Iref9Hr9HPEjM3a4TnoXg0I9FfeHE9NNs4mqSMhNUHa7sKuViNeA
86O0DE/eoVXCI4yprWG6GnEKlhlREStRE5HHinlLjurunmv3c3yiqRO69u2WlXgk
LpCIp9rTZMsIfjlSFRDxSvnPTwnMDhY+Jh0P5mXNbniRro5DBX08QzFltW7bLLAX
fzxSNENDCGHKOdkeQxDAIgGIlo0LT459DuGCnCxE+OjOCKmVdEh2AVNU3FhELWre
khPayj0IbQOD8cWXziqXZPvOJULMZj8SRYM5Z/dVmUYN6wa5ZRwMofzT0P/pF0k2
Q0CLPK8+zEju59ccUvv0ZsgJpukahrXosf/dNR5mSMBk3qJRtqdogzx5jsmKDgwi
auOpzcL7HTkYR1qIakOlB4bCymwA1VGwwkKISfDLfJVZxQu/L1DwyWh98QIfvj7Y
0VBtxPv9x9sIzgRdWPEb9HzBF3qUzY+yIvRIBahNyEXsTlkxcRuBDWooSZOLPspS
m5Es92ZSZSuUnwNzpBQZXMPEmvXTmWyTunQW7vIJSlgeEz1piZ+zTPhHQc8t2oJT
0RPUPNNIXNrN1j+ZFlvi3kJtLuRKN2EOCGFssQjQ+q0gTjz8C07IHxIdRrWxFf1h
cnuCSfVJaZfZEBv+LFfHfcHkEzlMmmIjtdRXDIzZLKHtswAfiq0NnYxQ11MjgPcr
eoS4VvOo6TkenBNUzCCXCaPqVOirBPhSyn4R93S218nMdGBwAVBYhVNundC+0nBO
xBoHXSOtQUrIzKBo6X0ubL62l47HKjT9DflBstE5o9CtixuV8XYPVr8tPMbtf1dY
muAx/bDWSNoL4Nn3p7QmkSX2rO63rKcYPyJhhCmW6AOXITLTBHeRdC+Uny8llly6
o4qi1wDwidH88E2HiWtwmbLjUnIekOJu+zw7TqZ+RHTM2H7dqPXX71VWT1X/xlB4
iGxUumAlVB2UqDxtYJDjtr/Yed/4C9jMIF8kP3FQ8U2B6zPCmphf/9ARECOuEZD5
F6AxdHDznbi671oRy+gcozAqCtdpfdtc37+BTlkKS5DfsEEdhr8IOuKSb5OD1P41
i5YNUUACHlIs67I4N3IIcxi50ZYFja+zB0wERJ03+q4CXY6LK72wR1hYJoippElr
zfgZDtkzZhnETfXW7GQscSBlAUSTeCF2DGLtvvlNZnxQmg8dkFsJCz8c47unmZOV
xChNn89JU+d/oQXTmiLfL2IsbmoR5n/Aa6bvMu+eeWKw46Z2Dax5H9OuRBIuHeU5
aSKHn8KQYSzb7S7+xzfEjh6WKgJLEIzfTOHmUU5KlnBCjQhDdBoxnnwS65NMEInt
b2QrRcpZ56raXyxpBQKCETwo8ORnPHcNDP/ac/FC1srJfsV4mE2bH7GpHYaODPZV
cAzUhBs54+xjJPlFvRTsO9130cbC9usMfV1c32pDskDJoA93CxERqYDtJbCFaLzG
DU958VYxdbUSp+qtjLYf0pB+fKjXd04PeE6x+OCLjQEfUJDaSoh2Gc86TdmF2IVe
KvA6vGEKSCR1/yDwgwO7cp9t+sMlArpxbrzUvVOcVobYt3XF3ATciM5p76uyfHqJ
5Jppza9EP7tAKOQrDQg1HeXGkyTzciaspxk0KY5kq4Wji5tap3Z5+dA1ZR4Alp11
rcH0csI/JL5fIHm+++9tlRKEY+Qx7R6VrtZT77JYWaF7AwHZxz+0nAke/fODoqJ+
9h0Ab3BYLXog+5clK6zuIroAbDlTPIg/9YdKhQmDA0Xab2dn0QnyT97IevfeAH+0
j0T44G+XFdB+vMpJYrCsHurTZDfsOiKoneexozJqR7qKCz4aqCopExxQlpzBALnF
3ORy5H6+ep+6sVxofVUZy7y2gLxhVX8VL/jMAZULRbo+iTxOmYASNypovXQkSEg5
gArwtAYPfyNLEWQjHfUM93zjP92z3mP6cbd6F8fsSyVfkXVZQn1+UxpFGkYS0Z6s
i6AUx00dQgCEK+jBdk+TF7mmjFdrxJPP4cojaHvvMEnCI7c/TT3KXzTbjUGFj4pX
ulhO/A+lJ75kcPV4OyJbtg91TLaiML1zAOZAS1OBj4p7LcvgwCMt70x7kq2oJoUn
d2feluPKt0cx9zS+1gRXDgl+0hwVu+qBrhmjMMQ38/WWJX7EK9RtIV9d/EO0UxPV
cmVq6lZd7zxmMmwGQMRJ/v4b7yiPOBzfueOrbc4XMBeQAFH9gb26qoTQgeMqwXgg
IB5xFfJ4iIWo8oRtSQsgu0Txig3blE66C4qpRjP8RQrgiQPmkybLahJx1dcLGKd6
ieglDzcevhJiDq5d8S7Cm2vwrafPV64/SytE6blYjZ8ZAIAf0INZi+n4L/qdRqqW
pWHG5rTJ4B2roOEZBcuxL9+RiNl1fJ3tO2k0Zi9feAjs5dMAxPepXr9Np+fMlNy8
UXYVFqRf/rP0Ofm/NN/W1o6bmmcsxb4j1wtEoIBzdwbpQNjafsC5LLTASiuWqgCB
WZ7L3/t+ptZHF2HqMKwAYuJUnjlVQZb4EZd4DX1pqQMvyL/LicbuazAL3Y0ooLpD
0QbwTW4klT/NwyrSiTkVtTwiup+6ASwM6BCez5ml1CY/6Pbv4oCOT0E2Sm/XrKjG
c1jaVt+TOUxvtMNElI20yjo0aNSnkVUNpUIfeMaR9KKUSIB9R4PBw1AgYHyqPtPC
eAPrpUtyghVZKPD9ZB/RTHKFOSEc9BW5hZaJtolxxOYEw2dNt0AK6wfho1q+tPg5
P1EvHbCEAgJdQTFz/ryHG16gEZazwEyKkcFsJ2FjRxx/0vKJPD6OkHF72AA/tU83
1WFxNnwqb003+VdOKLAb9uVJa2D3BgtxbEKbF1veNo4VLCPTIHg6IDsquR+0kmEL
pbXvedNByMZ6LcYuxLLBCKHTr3Hwmr7iNzVPx3QH3SWS9yM1a8tBt728WGTa8fGQ
lvTchEPUnmBkCevxyiSIsI586clFgWZUEbJn3frOC8zNJgG1H1jT8HmAHNzBQQmm
gcojzIcg72HrMGvU+OdzlGCPLKIVtc7Dg6saetBTP8ARt1B9hHrj6yX3xoleLFUO
2UhRQkCa1/cxbpJuZGlDTghxeQquEO13ohAmDEk/UMbBcpQ/cG08LaAqwvO2Xmd0
K+L6u4K1HX0sITx1ryulX9bWiA7GKhGWiz2y0+pQsKDWyrg3Cz7UPanEb3Cnpyw/
4KiZvQZiRXOwa9mQhRwZ0QWrH0nA5M3+CJnfRJl7g+Cwftx0Y4CINHoDplVuqFdd
5gWtOB98z+RmVS341BvOSujxm89ljf2LO5ZZWOoZDqPyT5qCfyjE5k9uv2/Bno6D
RRsGdAybONKmOxVI7jxhq7pi0xBtu9hHSa+kg9lvL5spPGr4SlSOxVpUnO67y640
j5y1plMzmSVX2g5ure/qJpvZcMjfVb5ae6E3ghfQCdNAyskMjg8Tp+MdkQQGJ0ue
hlAkyg5cVuEgRQhVbgAzJp2kv2ozGX4cyQUqVI0MGV6UzgxHqgYdEvBJj+Pq8cMQ
rFjF3s4XPjL5lXNbg+H4N2VbOfsz8rLwipqA3tjeL3i8Yjxx5UFNwtZJR+E6WYQ1
qPH60r6SEDJn7ci0yxFvqFeDmWAuwPwBN+VR5HBd6cErR37/Txp0cpJ4kFbYdlwq
leDNFExh9Wh8wb/8x9uyz/tcLGC29/CT0bChHZ58GvDAIYgtAqOLTIZe6f89AFnN
TpuRox417xNcJhJJS/kb+R0E8L2lJbKaBQn8ap9Ucyy87KyPOfdx65MWZaugQCAi
RfwPZcyXkT3s2l57dUUVo9eOr2uYu+Q1uuKzRix1RlxnVB1RYsMxAhzJRQZ0tRsE
uxj5Z9nFpQRG/oOGuvzmvEa+vzT8sltCfAHavtGy9poNZ1KOsu/Be7HauhOFJKn6
0csHk+skPxekIJ64eZPD/IRvEEEb00Qv0nCcG52B9949tJtCw/SuVbi+P7ql4vgt
WvEJcihhOoDxbF5wkACiUEjfvgtb4QRW6LnQMZur0gGD7FW5sxFR2So7Sp5zItKw
n98Ou8n00lig6EYDhqGGiBey1ru7UoJt38bd+Cc7Zvg+wZaLwuy+VP+N+BxNq+73
MjM7k+8NEjWzIV4ydXI4ebtXiAs033Rp0lLARqwfR+PxEYs6hTeL44H7dEMpNrwW
qhKBfrJKgjhIXbvHBHm46De/wwpNYsU7u9+ZEDmSaqh3FGf12Y7Myu/QVq+7P2wo
XAtchMi37V9fUp5DFWZwghJTOajEMM/ZqNUUux4u2yigePTRrvoAn+ghbiaMw3Y2
Hc+IpgW7b1/1S/NmKj5ot55ZjLGY1gXAk39aIWB58B6O0qBGk/556KjdNdszM+qG
Y1faldNngwLBCIMRFPDWy976vIGLZ0oYKtqxKlal7YOej0uxi9zJSnK859sCjXPZ
5E5FB1XUFN2vBTvfygHG3JG9xdThlTlN+ubaSspkyO8F1sCqj6WYFkSkf06jn4oi
gL2eYwMrC2GnIp6t6ZLCkr/MDtMmIwg8R+wN4VsZrke6bPDOEGzlK+YJJOvYpt3K
ym+pFQEp1cUs7Emv/BVDV6944v618wOO6j25QzsugxA/t02ZWQoRZprzhFXHpa+n
ek5D1VI/1lEa9xXkUDtApB+cx7QsjQUZY+cYwUTOo5RquZ5Vgcbq6hnlwl/ux+GP
N7hUMSKwI0BHqcjucSOLWy4FIVlUOY4kcMaGp5txIAPBpOMqwPU9CWZNbQ0mQ7CX
uDFmFLnAZJ48Sve3oD5ur++JZ1q69HMFAK0ORJ9gyHkNFjurAgmRbpVkFtdKMP6X
KZlsxQ2+VZwKsXpwQsLIs3DdZIwys/Fha4utb3C/ejOCu5l6EGnoPol4hr0RQ1eg
84DErT1mcKH5MFcZpzqqiNohrRj/QbYPeX5htwNkTaHMQM2/xCJT/8SQRDFVn/qL
a/utZ1OJYGbtM8U4Zc5prIg8dINza9z9WHrA0Mjziyua/SxxmVvurF3DUiQdW34h
ob9cApHpvv0kDq/OfMvuSt1h5avCXNBiTIOh7oO5ICfYYR9CpZMvKv1sYJ6YLgnk
gcAhIe4eabpSP9l0nLRpXk7LlQSQTv37OgGspUrGXrPFoAtkE14FVlLowrQMu0AE
6Pw1TGRR5BBNNBPDRfiEJBuLWdcdtoSYAvi4FLLD1Y3h/2WPyjSsK2J2h2orRIo8
qYAJ/8k4vetGHZasdF7+a9fg0lIX0HnuceB+AmcivA6S/p5SOwII+XlMVGlAz8pR
HUFnZNK1A9jgrP0RpKzNmkQ0VXaNm52ORIYckXZrlm5qpYG4mpbeiDbu4BnZlij3
3sN1DFuPHdDpTa1Y2zkoTIcRodD5PYoci9Fje1zd/d1oE5aS7s0Qwh4Odm0HAesc
EkggFXaX7X57gHhXL5iuahjTjbtDHnkldA1vFmj/zl51Z7+zoRTChkGphhRMLHcb
/XYoBRY8q5gdRxUvr8lEXWEetoSk7s9MA6XuvgHDFRe5Yq4mpzA4vVJaKOY3xgHb
qIvFyNefTucnAvxlHrDOIx72KmO8OnaMV473szW7380FH4fYJxGZPTh1wvurwXLX
ViVSDGCdfgdMK1PCuMnFbcijFBY64KG2zuoxF0O0GhQXUT0cU4nOJE9ubgjUbuYZ
jl2sgqllnZKOmVjBPqr0awjg+iVtFEDA0qBI5mODDqZfsr2Z4T6YjDl5/zHA6+ig
0Bgli7bWnfz/THhoN3bGVXzzHc06qVJ2xIFz4quM/7RpmGabtVFF69R9ZlMUPwi+
sy1CmLSUbl9QO8LJAbNmkcPsZgUekEFS5DQU7bdKr9CFKbNzPvi3pNwi+wxdxWw5
0JDCZVGj2XLwRuvQdxA3EgdBxSa/eHrwbJ2D8BNjWm84/U0mKwkhNURshoyYg699
b068B2EthapxKTvfwOQUhjZTr65PaWAr6CgNxwcTQV051ftS5y722KrTOEeSb1LZ
xD8az0w1348sLzcXXBA3FD9SgObCP1zY19Ts29EDS16HUZFgZ1DOyeOnumAV+95O
6eEqqI2TvBlIVAPyI/zpwg1xKnK4nhaDc/yFbhdVGLO+nyBhz2B/sjKIprEU9mc+
bXTEdrM5zP18PpGv7LgVuHvT31naJ56EIvTsJhRy/ULTq79ceSntnIx2M+BdPAWt
eCfJxtFGDdEPl6DOVRD7L06qDiU+KOO0Mw5kzsbeJcJY3b7FmfKvLe4xKbgEnHUV
q2onaVpYY84NtyZXRjkcA891yAisBYpKBDFc7e/5uugz/TD6Mfp4aWGx/u+845DH
msVeljdare62sSG8JdBJDXbZaDqVZs4fmn2LYiWNUy2/5j0TptxkUikHBtB4GkTM
POTOvgL04T3hJSEDuCNG0M2h6TjgfM/Do7lhiziubwN96PPnKBsZFwM7bbWBU/ni
atZTIVMXJk2s9os2ond8TDjLEfSujgOHZpf+dceiWsZOs4Xd1YoKsLqsQCnr3WQ2
G1wwJCsgBq8lXb3LtGjOxhhzJmtWHkwYrBbc8kOnMoC/kj7dpagxE+71bBSw2fwc
poUCHkZHwRHqxPwOzYhfznUNTZ3YkXTMPWz+/RjRa35Cvq+O+64+OHO7z2XH4nyI
1sGFmBIg7JTfTdAr7PoXm+gbOsna375fePc4VOJNFh80bQ0VSXOzwrY4gH1eN4HY
BFN1wtgE4hd2Eaiwm0XBscGnj9pXWzDAAPEZaDRfWHwsZRRs2tVaUKDK/Dklt3Cw
NVBeI9g0Q4Ye2cGA/XmoWQv4AX2NqqagZ8Hcb8+9MBuKmPNlbxdfp8Qv8CpCwHrZ
NNJIgDnrsXheLk57UlaM3WEH7ajSJlSZma+N3mR5Py/M7GY5Ilq2xKfKF8VAEJsx
6XPy0TZ2/CSBRID5uDmgm0NdD4uXHBqNbblyozquNZjqelY/plJcWVpXgY1snx7l
DStfh7dHRputwmzq5W5qs5O7f/UrjvbcKLfN0/cdgGQxUcZvDPQfR9EZQ1z3gnRI
DnrQfJIFnqkV2MYahsAxzTXkQdnn1W5uaHUk2ngEY/nHW7WakDlJdBSx1bupnos7
X7384ljDQ+1bRb8LNAvQw2MThPvvasRAgh0+10/KsDd7UUCow/55TntKAThmlzrF
IJjPmZvhKNL/HLkwY2YaH8k2lBuV0uZcWzTftYS5l73gnyYv9vA4/caTy4XKpe82
FDdya+8KYLag5T7RuycJTX7OPqeJxKAv7eqp0KEgrARB02gi5lIv8CacioyVYFqq
6AHmfecFPqMmSHgHO6lnC7A9Q9ywEEqKOvXminnIo3bRiL2tsRSilVJ2w3YtxLmF
CNdEwJAuyJJFyPyd2JBnR5U/TgWFvDucr4ns9pHEOD0gFsqif8+fMqBBh7Tg7ffm
8NLTWlOzf4Z5iv8VTDd2ckSK+9sQyAlER1b0Jpncg9KjxTvsbIgGj2rYOT6Orb2g
Hj2IvY1aTS6sbXLsB6ubCX9HUP9AZGiDxXjM4OOkcqL9XKuZrT4vV9Cv8gCYIsXa
LxOQ9CfglEIbu5dLeSATgSPJtFfkwRkP9Z+/HDnfp3EHFrCdqqLpGA1ATZtoVIK9
bBuCxs1n/nymapkx4w8ScabjTKbq7mxrPLEkQCDbkuqc5q81gFu+G6evxbobR1b8
zPpix28RqIDJFjZrE+OXRIKgOFVzU58g454Ooxw+CHPlAQYV4ZsHQf5Mx/Asngja
x+EpH4pyCvzV//E7qVhxIWCsX/FOjFDe5C/GoLq/uiJq5ikxe5ShZXsws/6FWjgx
YE6f+2rimgwn57NvGKX8hmwj18GNPhJ+ji5afEMtt7HfbEgyLibJS8fIuRhuQckw
Gzhq40pWhhrQoJWgMQa5/ZZU9YONLzqvvG3PB2GuDDZSgZ6H1Gv9eq+/A081GlLl
kq50gsocO8KkaibIxzJHssXxcnWTCBnOHlfVVNbaYHORoKbJYU7x/pcf7O+jwtsf
gTQnn1klw2YVGZQFsQTGlCTLvnISmDiT5jl3uVLKx3766e53LLsVfzT9cfoxpUZA
AEXcafXkGVF1EA3qppEqNCCeqveeHsac3RUnYsj7k/DrTMNQQTl3z1+rNFQG7f3V
pPNhh+QprfDYJ85QFfoUAU0YcwI/VobqWchzcPZl7uHZROv3oHimhSxuWafSwagj
+eb3Wsz7JurwiIw5RI6HoGZWrpeoS53cBaT0PYEDRX427YKmyHBz3A98EkUEnFR/
E1PCFrevAhvfLnJhEcFvRMogmcdKd2ixY8RZo5UAdRznpm4C3ZT0GZGqcvwtgXdf
vziHjdepwRjdpuR0jpkVhhMeQ0HUAYSPVrHTLiOG/yNQqJdrsgcBPsKVuI2R0pfA
0ZOJy90Ghdx/HElGwidfBg0sHiD2CPty2T0iG0LUPCm2Ix/q/M97tEhv/jTUkW4t
MkcpuTn8kDTRhBO6xuU3XtLb1aP5w8qZNQfS6ELOLiXxAvEvxI/2IC96cSzQL+Fn
ZnCx1b5rNcCiV4D0B8/y8unHpMzixc32wboDtX02fjCldSUNlM2L5RxGbOTG04X7
r5C9xTPxCQYPymlSwLvCWF5fba7+53Xd6ThSo1RT26sHpN7fLLe7O+ROMZD0dVJN
ZrKb14Ea3NiR+7ghVhB3a+St+8CAooBsGnjtdIa17icTLWnW7ZgwfPQqkyXGaS0N
UqvYjWNERfRCEGgS1/4GZvvFb8L1rafUCRcECirgvG6rG99bq4GYAv9NGbRfIkD0
jI4ysIXsfYt1w5DwZD/EsgRbdNM0H0MUgn+Y5JM26uA3WXIpXKHHU5RPbpHlmlt6
aAB9noDndp3X5xcQLtgHKaTi/L8grJttC7gpn9vU6Z2Y9N125dlio3RtDBKfmbyl
G840951CvFOpwdlP5rh0OG38gMJYuYKt1QRfoUmXDh4PIKIrt/mwoELs/+Y1gZV4
sp6DQB+sCMZpNfqJPMINlDALzTbsaQPfFtCEnI0I7UXznygMnT40MYtFJ04WRZ1d
aIYeNge/U3lj+2OuYaft99hF3+PMv6apNHBUZkxq5SW4itr2kqLIpPZ9Hkr7jb8a
ho1x7u2Q97fpOk50/lYxCXNMpqubLXgk1eshaq4SUBSz6Vg6PaRhXGpPiKvCI+Gb
6Z40rED5+2gyH6f80rOT7GnTQr/WCOSLR6HF1+DmcFSW3HAStzLixIbACklTmVwx
6OTx6eBJleyvJmRxbVBxpPxz0GyTVWjWNZ4rKPbfIROxFpDfA088Q+I9pRxVqxAh
mUS19v+3yzampGLpIQSYa82hDnEw/rDBHTeYsncpf8svrlWkgUd0UT4qfJf4Nvzv
CfHKyTJRooELX+yEdr7WUMMuP/6B+brYgN04uhQEMmhALac8bs4JiQzRU/dccirt
TIa2dUyVK0GzAkAcVrrCf3CnP7ndi7mA1l90K4AeFbUtoaX6NY6+m7uYQfLLvadc
OGLWlK0k+o1cEHAW7fjKOsROJO6cQ2YoeDitR7zlMOOEqysbEwI0KpclN1YcGWKz
T7mdJtHF81sYu9EuD0uW69cqIMXgb0As0xn2QklQq8jH+w0iA+9U2zuUUceA8El2
ZvrHnhktNoj2BjSlV1eSPxmLNFZaLo8C9mJmX7fDaV5Ay2loGZsC9D+Cap4/fWx2
g3bdpw6N2qBHOA/6+dwgpvkFje2m9Z2q1y+19p8mzmCXzvQOLJRF37BnBh14JQaR
RO2aCPdKpegl4xu+Zo+6rPCzrXLnjpeOr0Evd4UyPxZy1I+924YZWwWoiPypfcxW
yhAMpPVW7Hov/+ywzIMB4CpHKIwPObM4xvuUw8uwBZDswwaAJs+O5yxcb/ykkJOZ
MSTQTKIT/DI4zlMT773HPM6+xivMYe+LB3NNruTENtTTPE5tk9FEKFcPL5RaxDJZ
qRfdX6eafW1kjSH9WGiaL3sVN//qbcMUwX985R+e6yLs4lVfH+2pQjfMZndAtYeo
KJyS7U6gfbQHm5oKjQi/B8SEs0/q6E4zmOSzZZVZfyoF6iMFKj/4OfbrX7zFdYrO
rVvhOsNoXJlk0ddx6ZCQOfDCufFzJCp9RTrI2URlMgJgjhzFZqzgjl9AKEkHtKZv
e1OdpboBGD0oR4Tqs7BP1ccO8OF1o9PNi9rPkCxFCaRiX/+tTVGXmT+DIOCMl4JF
oqgKewBEhp8nfcI19pF6JKMkDi5Ky1ihyulgi29JpIW1keZ1ZpdsOiTgzOmzsWNo
Oyi2QPvrWO0JRIIAuQF2XnBeYriE2IFvtNUTy7LCcPnCYFZ+rBKx+OmoCkOkaHbE
y9TdVZx3BHCkV178TRz8dHm8qLjbUl8QilLGeOM5huN/vI0pripGTi3lrHZP7kJF
+VHKV7BmSzVkWK8P5MumihOd3MkNh26ZG/+sKhfDlWA9v1ovoj8uLY011T33aAhw
Wm75mn842GiA/KXYpcvg4k5BhiRWTuRMhZgDsLUKAPko3G7mmHlte9GK26VGjJ1c
Z7sVWKuBY4pcfkXh6OuKKHEHuKJ8cnd4yrQWInc6TQhK+fIeuCvulxqgY5+hD42P
O1OM4LI8561L2eOqQe5O9jG9HibKrh6vHmbJQyjcncu+8pLaW4oSMmacfioiuK/M
lhYS/bfT/SJu3MACU+tU++ofvkYXbQYmUGaXp9zgxye1tU4aR83+Cc215Phf957N
kS2PMb6i1WlXYFNnHGiFGzA2fEJbFPHgKMqteyqqFu/vgoIR061U3x7uWs8eekse
13dpy0oVRhIqjg+hM+vB/ksk78S7+vMRqiEkh/+qtT8mP7FKZzQY71vdVq2ViVGJ
7TaVhgY2Z0ZA3pbcFs5hepLW2020eQ/mIHFwsw6eaKynOo50VpRKhWE1HHCVF+Lg
7/K/LnuShT9YWdqLf0mU7V1/mHcbkzIoZmTpvVSwZ/XLqGZORE4v9XpBUYCddJZn
R5kOvDkI71ap/7V4xkiR5mEun0SIeb6adFja+VEXdxS720QO/twugyHp6hguqZVq
+ZZCq72gW5t4A2AlrpbmSuktBz3QVpnhLTViTzuD/OVJPc9CQ2OB/Sy+ayzmoHv+
yUmbFqkUWKRVrxT6iA2A3af/ch2y8vYlARKs+ghJJuPCNNs54CXFOtA+Tz0+dhGC
ssv4jEhrlQCkUTZfEoESeKHayuyQBUwcThCK13gKgfZxjif3b34ZtkVJ5F2R4zEb
v3+4I9mQpojQ1wUK4SrVGwcyNtqLonO/Z1XcZ/UmQWKMVQbhVvJ9ksw2PK+N3SbE
hNeSLAaiffzxfI8NVHX9baQxSQ0ZeH4wZHQvO1UJHuGXrqY0iekQiBx9qdpI5zJz
lYdStV4rQ3dD8kQqIRwnd4ys7lvJ/WjNjr2fFqmtDPTA9ztQV1No4Qdz/AQiENa0
hZAuIR8aL8iEPz6PERBQMfLV9oX7IP+EyCexAg++Lu+RXLIyYTUJ8H02eouk4FDE
pe5R/tc24EAUTeKxNE7D154WKN1Buj/ZCk40/Ju5VphZ5M/IuigNaH96UDy5cBBD
Xuq1ZNcxmLT+FR8y/EnQKLFiMCd/V1m1ZRgRC95Ah7kv9gI/U1jv3ex5qFWvQF6x
gOp7sgKAJ3/LNCx+qpyhJLIHH7Wn6X2Uuu6UtIPxmRkoZoWvC069auJacGQkX1+K
gbsMgZWIyFx263P17f3yVywZwJq+ZEEmTSDe/jnWqjQhNy8hBiEaq4p1MWvW3YfM
/NToeJgu3W1CrxgkXocywx1ix96KpIeybWPd/rpPKCoQpP+STm8N4NTS0eesgfID
joTwti23jsV6kvmHp3q8enkRA3myBK9gXsP8b3q6KzY16/hxHfpQf4nFgS8lZfOy
nCPI8Gw43sl85/FPYR/yBA5pSS0yvAJpY9/tb9QCC/YiXF2NWbZHX3mQYzw6EecR
OJvKoHkFB/y3CAI5FI29ylFVFRenQz8+pXFQ5zovfX3VEB8ah3Sim8FTYWycik9h
UEPqnheIRNbB0ixOUFDls+79lGhFzhGS0NAGnErM42ZUi4cb6FLSC/OOs40if7dW
3ohhjMAQ1hl8uxd9peEWADk8g6B3ndEtk1InX4l8Wk48Tfp/tMusOFwUntteUUjy
zjTom1QRpxc+T30y3a8HZ7UD+wAPEKvupUB6KX/DoPEA2zujfpK8M1IOygyScHGI
m+8+8WiwqiEZ3Kv+d24KVKXeO4rEDl5RHTd5z3DQ72rob247RaQLZkA3N8sFFTmW
tb1aa1i/e5ytXjG+QvuK3WfqhG4OmhCZ1j40uYV0TQXG2Dsf64GEHe0Qvhuvte8W
Hy1S/kNqzpGRj67Cio0YxePk11lqvpO9VMPqxA7NeFTKPs1oF9Ds2H2qcrqV+vZh
y9Vqb54pQ1OEwvtLhBi2TST26ZtlevqELpya2mVQsiNK20D7+WAbGZbfJip98AT8
sXFOLEwALFgo2tpxY1MaLmidmnSarXqIonlAiYJYf55KT14tthAvqkN90sBDljdx
CSzC3zUFMBJsGRvc9DOJDY2f9z/ojhM9CX0sa2GcbydCsBJRAYLsFoXCdgXN+ctp
+Vxwt2BX/hZsR9EH56T3od+ZKpcRem+euJh73P1ZlVDct6YG0BzQSiAUtt+LyY6W
4p8IcggUuKzPB/vBLeaZIFf70XbHl7Hqs5Nb9U8UyzHIR0ZGks+a3f4apWikDIV1
2rf/CpiRpk7Ku3zm+6cJa+G5zsfP/YdJ+/H+4ueszWaKfRZ1l1JpktQuwt/iSlkr
pR8Youg6gY5Z4nDdaIRdBw1kAJ+zf5durX5Dy8bt3TFovo6Z9PjAtDqAM6rI7Lct
BdCNH3ovNbLdDYnI7u+FWr9ktz4320JtTxbjwh/fDEQLVFzMoYiebcnov7uVLO1n
PjyIRO+jLXzYZom6ImtIOnrhdF28FIQi4B+uO702asJoppRCxkN6mhftxguevpDB
aJnw/S5ceoaAeUminjlYVDIX6ldwCu+0F2UgDuGhf7CYgsbzcgNj0CeV9hiho9AG
wGelTGaJivLySiX+vXReNkTsH+3qYDriCiadx2ot+s5+IipwcpK0hndHcoxeqhBP
zytTTZhorUuGAniD8Z7WxXyjRXUKtOJMaiVLihT+vx6iDlYbrwVaZ5dtV2tI39Uz
tWfaEMfYwrPWO+QOLKJg5f2usTCl/Gd4+ys024VJxmKAglSW1AmkOjK0UVsm1COK
3IcTIEPpHT+b5ZG8z5ukEPpHh1TjPNhnXY4k11DIm5qN2xUl7C+iBQIUJbEZOY8c
s9Uzsp9RDYYmCuL90atbmvbv20SZ5cmKrYpl1bKWFDmYdQXNbAYHzOhj/A3I5EP6
4BC8uVxqgEeo+JOMY+9D7eFP+lzIISkH0ZjPmu8z6wpchIUAGvn9XsR7aOfgT5Wi
qv9lPZzaIh9jWfe4pgZCAC2DqP/JLJ824hb58Rk6sRY7swMVgSU1S0FvwHFR2wOO
9wJDxtId7ebRN60japydr8sIn6Qv+0IpBSSAYV90xi6oS9QvzD2bgIZXYyFdofhS
yh54pDgEIYRGGqM/tQLbWt5291YZhhq2sSLyN7MyozjVhzLhCYb16Hq9rY1aJCi9
c+AWywQeouV8Ir4wCigjbdsVnVtL/FYfojfY8a9Tv+W+sqEdo2K2VBX9ROn4Wo5U
kOpVquRKEUsiMFeNtsEekjAuLoHbwgKlW2U4E7934Tgirk+h6ncJ5X9LdzkH5lvj
aFrSHrzi6dTsexfK5/BOc9HLRKBXwefFi2SzViC64MO2qiZTn4zdEEpzQ2wAe3bR
83S+1jIUHpEabrZnW2Ifd0h2Q6luQSmOxBwRJjCW4tSrutpGe2Tnp39bj1V1198Z
SNNXE0o+H9kmOcTlxCxaVdASidPP2Gsy3s99I8lYtpNSFobHvUBOX1DAmvd+HXiX
ruwCZH1qgLyCw+9irZ40xncq/02HgcNIQpy+N25NFCBdIhS6IdDEqPPH7cP3/Cco
HUJw78Ghyq5WFoiMHrb9kCChawJ0bAk5235dgx4TyYumplq2l3xe/qpRIMGlFMfi
FWDiLgDALd3FnpewmI1+ew9ejjLzaCK0VS4xgVgOVChjayzPmvM30EgjJCzbN4/D
k+xeaL7AhGXlHlgnbKn4oAjNQ8k++9rIXhhTCII1u3vFrgfPFwyzdkqX2+DwKDPo
HO/fiDNX+v2rnUhlRmEAJYXqUDTJO1UMC6QMmIVNauDlApfuvL9B6WvtdvmwCW3+
t3lc9tQHeKMUOziLZSINjxbwgcV04/A9RB9rAZmNEK1bFvTo2CRteyecSMu7FA1T
dCKPbZ4NGlhvct82aSVc/+j1/lWEp9zb1iNiU9RbfiL8D7EU3SgpF/2aFWArraW9
WKEVieWtvzybWSGpfIfRGVGryPc7yVUFN4YtU1741BHVJhLGdzQ0ufe2/gBiT20E
ffhmER0jOYQzmqNYWzefv60xBn10/6uwIeRtuM2GYNwF8sShg1ddBG0lHFAnkIq9
+udeg3mCGKvmTb6+G5PSGrid53l/42GMQa+fizqLEhOqN2osMRsxfoA4IaAPJwZQ
7Ycr4watV1Ds3tExfr7Hbf1317g9ObMXFE+cbC9WVw5KqO+z5PYKUBrS8wrn57wl
JcQm38YOLzgI7qd3bSv0MAjaZ4/px0HrwXYNzCQoL7eAK5clvEZF4QP8jYJdf2R7
mkR0uGlUuDHA1JV3ehh4XIT63yP/4bv6nrkNCCmvjjIpKnuIBolRuuG2jUIvUSV3
kD+Cb3XPwekex1gwlMQqNW51Wlrn92GLvFOJBiR+Gj3A6Tia/BT/DzjR7/BZ/BwB
3nhCteoYOtXHxY/ZO9L8nCFTY84ANTKkuX2lcXPCQzgVhbn/gutLGAflvZfLmmxj
o7ZDZnc6/9S8Oott8mooL6EKVHew0JhLbUgUcBupS1N1g6PPDVt4mevu2K+AI8kQ
+rcGZNoCn2fv8bH93DHKYPu+Z+1pBjxDlFiINHY88nmWBQ1aInKGNNxVPRpRgrU/
yhO/une4FV4+rAPAw6gbHETMua21r8BDUrmzQ2P/MkYjiOeWbL+ZMXCByD99AMgR
wtfKdpxbwkEpCp3RWQfVL+lLOCt8+cr2ZLzMjauVWYObpxZoa3vTT51RWKuMk6ya
viIw4HdtQAw++Ry4E1WZxSKj98i3DR8DbtNgJ9QwWUJGOvURNqJzyqWp1CrNL0YT
PY3Fntn3sm0aLEEFdNW7IzbrMcWKVxThSarhADOjxAnjdgCAi7lBUI2GZs/twlpw
APaidwawwpl2OuH1pXNT463aGrCPOKEvD9kKJ5Vxg0J6nFIGCJjzfnM2mYZnjfYc
yNhwCjkLM7y7HYJ2gYKatouMZYUPh3PT80Kb8ul76wPN4m4xNCNpgYkite19aQDD
BN+kustuDg1oGZ96/y5zRu0xTYUOD1Lo6v3Eyjxg85JfuDcXCWdBkt2VPvn8tvUQ
A6NVlgUaK7zxo/iGUZAPrnirQY9xeUcRfa5NpDg6ITL+nJlV17r2wrcYYQpsIXHw
396wRHAZMrHQD4xlof7yykqFzqe0343k7AoOXtriJJ9CRD5Ifq8ME1nPSdGdJL7t
JcaPZvMvWEUR360970O1BUmVFdayfQJqW+0NnDdlJ13IYOfsAcE9Uoj1qHurWUSi
yd41riYRRyA11hENm2i6VNuT6uGLKUnjRgQN47EYqtv9DYbHo6q0l3Bb4kgMTRHN
e49griCtB/fQ0yZtKWBRm9cpaC6xsGrApWfjMGL6BHiRYXaqPLc/NwS5WuRwDpNp
4Z/w4jnTnjBQbLyFrAib4E6Na6F9azwTZxhuGYoPGjkqbusJK5HHXmF0D6MqBhHu
atQhU6/rzzxn2vwK0Wy6fOOmm/OZLvc2DN23TnQ4rSh1zkOlWLG5020YCWVUpzb2
G7qeiUCqzVBtZoB1zAzsTGsIPvtEevlOlLrLett/oxF5JhCcRIL/2ZoJ9swQkq3c
coEKNj9l+Dtzz2i0idgXd1GmJuQru92cfJ73IwUKxHu4I2vWN5eb1/xX9FUzx96M
St4FsHHVPqy3c4wEmhf9gKk3b+dSPl8oM6u0lKx0lBqAa/46SWnH836LrUk62qHA
hMdbKRSacSzvwIgFmjBygHnRFmmzxYELv84XSVy9OQLFxrN7XnwAsXuu1FXd/Sjy
suoIGJRnoizugp9lz2QRLBvWK0rxgKOz8iQvwP1tLcjhvnghEMHfgsjL+D+TCJcO
+WjyISVRkUo9Ud0EGPJL6Dk813i0E8Z2+ZQOQWa3kBspPoF2xdJ2DY+QfurIi06y
TMHUlYN+Gzfs+TxF/dQHQ5mDP5W4xO93EQm+codXst+++fp/Hga2tFRITei/2Kus
Jij3sb5084WaGE9ouQ8ZsqFQKBxTnB38/voiWrU/fWEP44Q+CsG+ohA8fR0sGKjZ
UGkLcHHvXmswWmwMzmtTzgh1tnMr4TAz68Ae9ZuChg8L08tpNNe5S0SNIBTPSky0
YD8Oj5Yj2uBeoopXQpxp4UgkdAKMNNeD0QsKFZaGX0tXylh4MesOGTk0XD8azUP/
PrPKNtVO3r3Fyauz7dDFbjkC72uxfagPxxjBoa6qa3aJ8KXsPvnDPqgOcNP2mjky
oOhpDufbCOOqS0DppCoQdk5q6q4NuWEzy7TKRX6CDNZEtWWFIT6aEqbZhUWQTRfY
p1sT0qozoioPz7P+SzkePxqNc4lkEXEjtZuqwqhUemMLXbdrcl3t6orU7Vw+8eLF
Bxb3bCj9Ohb8DO93KafZKI8PNGe+Se6XMX+Kk2fgtKCscnV8mt8KQSGTskyIdX4L
3BiVjUK6cV444jiO/IXv51AXfZvW3XThkDO7bL4ROhS9Ko3nsQnoosflBezoKlks
SFelA7ffokZxfViIdGcgouic0cnq53XM5qcE+bTG/nblvIg6KAS3shetAuzU/lQb
gANOMEsw/QzyxV1fSqAcKkmSWB3udLs2LEtKA9WcbFK1CgCoZ5UZKxGHDheBasTY
jQgjY1PSISCKGk0Y7rI7jhjHNLsBO6bMF42CLa0+fLVktvKnFBp+Ro3JxZ31VSFG
syEkREaS+xOucO5LG5fGmAZHCdzdy//oDP6xYlDayb4G8TwZI4otJqRN5/reqVSG
t0ZHt+rwFFpihlzXdLRiquzHHwrDASFF3b+PNMqdQ32KzPp26eQA5e0+a4q+QXUE
GWqLizQly4O5VaYBIlXMtvRXL9Kadm0fhx9mmalc1QSgmPGFu6X1gji591XRcr+j
l/PkD3lq2W26Wjx7vMja2fLKKOMUNA9jcB1LBzGY5Qaz+WsGCrWFvVJfWu2+yTZT
KwqmanilOMNviShzVAWED0EQ+w5NGsKhsg/iKeRe0Q9bl3ETiAiimp0srDJLff9n
+CgYJGpbpdZk0eYib5Kk7IzWLlYxCSRSIiizGmfwLLiczTXRsBSnePgGGS9wshGU
rlzGNsuEggFQZ9dfNd+5eXdWxK5fsk6K2LWhAH2jXuiW9Uh2IER9nLlJU/TozTEf
LmPxQTX6J6zS/n626mC8XloJxf/Te040iDc7C7GhbSl0f1cGsGD1yc8e9scB8e28
SN2V7Opp6oa0lKuwwVNO0Tr5Wh4L/HxmPp5pMKfRNB+xGhyfDCl17FtEQ3TQQ9pQ
GZYePaVJP5I69N1ajBP/0PaOsC2ouSkYV4wIt4evStqWGFYDYNYlBmvmiExl8uBT
GvGxdqiVqSuf9DwGSOC1+MzVs132ZcdMdRDIFcN23m4tlbaHbsbgdFDAlXYVXkcZ
jBEw2eXcVHdcJ3ND1Nidn8O36pCAvrC6e7ZOQbRH4feeXg3DlykM9tQzLW9mbrb3
xWn1c0SwRGwehejTRTQCt2t2pEsTVTMfd1Gw+hd+cbuSquLRdqpx+b8Pk4S4rbup
BEvqyixWhe01o1nihDo9YtKO/uUWNcCddcI5YV8SDn0eSXnZsvqExtdRmX+HXqHp
tUBMV5gwXIJgdLyDmfmd3KxUtwgCicjNFJG0P9iyzsv27yI25+zqzmgQZWCVcfnt
HXjZ9IVNXPVeWJl6G1mIdLyYQM8k3yxwIvIoA+owsPPi09EYecXthZD/0Cx59+bZ
3dsS3xl/kL5F1Nlx+ABfyd3mrf5btM97yUgrDO6KoNOGyL3I9C2nKvlpr2/mKgzp
hGSmiMVufcCZTL1kZWSky3VFgSjNMWi22vq8xkRBPLdcdtoN8DX9WZZbA8Iyo3QK
zKX2GXFSUfEH2WwKZ6U7bQcQO6fsXkowNP7rlThR+6D1oFmaMqXnBG3+ei26gqSe
HIoCK2X5wbPBrHYYUPw1gjieYDw9ML++wAngivgIwLJu+0p2uWkDxzoQmJQIgqmk
hZ8Pt57VNKj1KGDXd8MjEwMJ0uEcmdBVYl8xMXEYH0frVzHwrkXYK+KiDtQaR+Da
LL7B8Wg9Y0v1HW0wA/wwG0Zh1m2hD4s8blnh0uLn0EYpJarhmjBnBMzTwvApQvRp
Ji2L+2OygPdJEKUhaHmdx79HOyZ906GEeW9IVMz0UjEzw7H6tT8x2tCxqWrDethM
HzJRNf1dMMkt3ieTCB8zdZTast/6k/9/Mle7aIhRYbnqxkyE3CiJX6h8/2eKbIiK
I6d41jE3jitR3YhM0+X2z3DqsfugVU7p4kXJh7q+cDgNfRX8AYR9+HRX5zZIUbHG
jBMUtGYaQ3+aHWn9SxyHCuyXy8yNP19dCvTafnNM1DegSmerr2mSNbarP46jck6T
uiaXazHjJbVc1oA2uMx5j2WCA4G52wYX4xM2QjBRkyYKdECNzkhDbzjtMIC4stmK
B/RcS2SoG7Q8doftD0gwdy+laRiEkMTisPLbbwxP/AwjDqT9AvGdDUKvi66sygIC
4x51knAuyHAnf9Vq1yOLXDB2g5G7Fr7VRMxWu4z2gTfcf8NDoTcTDEmIqf104LPq
sUZikAyOSVMy7bDkL/rwzjsp8nZjGj7FkCFJTrgu4sOgxMe/0+AUkyENSb7xfOeo
m0WIt6hUXHCxX27jn55qjrLfuUkCr+SDJeyz042CcsR+wVJSds0PBnp1hfPZdbqd
M4a84sFAYBNjpO6w5c9AE0n1DrpxJkbl1Prn8yQiNm3GM9PBgydnG735OEDC/nqM
le58Yj8xajoWazTXRl9Ojn3u5X1RJKPkr09UMLSkNZMLOqZ68On0d6Y+LGtLJEFA
ttyhNg19ydn7GwSTrLSBKKo0EoTG+ITBTox9S1e5R/0awPo+724DaHfKPLxEbHBt
yCueBe8QTBDubR1CgtG486VP7M+r4IIF9VabepUrxN6TJmNmnxLDjM5YVtCvJy5c
y5jV/JPibJxyZs4qmXLEp0N8zywwJMmFpzDelqPJqp3eZAmiGgwyWTEE/utFHiNi
mMZIlBbBVIiZffrnwSFTm1SPazg9scEA5rrlsKSsnv8MeQbmE6zbymujVK1r/rnt
MzzA7tMzAVJAjm1azpdwemfiy4vATX1Oi6kIdWxWkWS+r/qkDpElyjWor9glPHHX
g5Gwr1sdc0DfcDyd1uYF7szC1xP1jSMPGl+B1FdGVKMKxYqVKnDcsN6m56o31grW
rlEv9ln/vwaNvzsAywM9uSv4wAwO7mK/dzc2Tk2cAUVcv/luazuQEXvT5vXBodRn
CWEAgwMT/dr1sCGFGzkOghvqHLN00sYsHBYIuCjhpcrpk4eNh9D6fcQFywTpgQFl
1+RvrU1e5ScHJlvQ7GgYLDziX1XFU9qLlC35dGGsKUbLVs8mvkb1NZxqFOhxgPH2
223DNiayZcJFWxW4GhMTCTewy7LlTc7gIGp6fuRpcHDLltZhP3chl5s6leAuZEhs
DW8pJIzj9WifTHj62PnI6mdnHL60Lp10O8xGg1p6ufOu/zkxXN7G3qHQrhHxxqSb
jrvzpuq2zcLdSaBpCzNrydFwqenp+xVi7v5lMS1QXuLjdAYqQh2/6eCVXa8TxltR
LF2MqlP//GFWpbKMZO/Zz3yRqhlOTyL/2Xsd3TWWPujPKsVPGHsYahTK49fTeowU
ajEhAsNuvCsI7MslQffCTIqiRZw4dEuobumKjmjLEkrsNWsEpnoKaO8kfaAYbJbK
OfSjV6LLVLAjdtZR/N7brFuWD2njJFCtuAGaF08frInaBu7Op3O+DObWanu2ApGp
/xLQpjryBgHhZp/RWS6yKvRaQrK3M1QXZKCRXmu/RGSlZkyejJE8LF/hdSXESS/U
vo9CbYo8fen0bLARKWrIhHkg3WgLwU/EEpHdqxWIb83UmJq2rtnwmTCsYRAkKb1/
FBNX9CnMKPEKxByMPwXuShy2C74z9nd7LdB3gwlAg1SQFPjn3SW6AZ7h+ZaYlU9I
ojF0UrUgMkTD5Fp4wLDo01P9wbhg98ijq0nmJCrbuPIF86JbDS04r1YkmIzkqE18
9He5DKTXYz/DivTWDZamBUEKFw4V4UiUVovZtJHbUerFv8RewMPmHDr4MtzSmKkd
S9WGtdI01odWYFsDEp5HEbYly96rTHN426NY8zKn0GtaLR4Upb6eykU+RT4sJfJH
mHYBzFE0jRBiLQfUsbvzWJScyACyVqPp389H9wkRlnt87Aglx3X5swRaGEnJ3MiU
f6sD/X+UvDnSuHwwccDcg4YWuQBobUrkKRnP98YpTy1vC/majaLhiF3UEQRXxnmv
qFjPCv9b7XTQy78e8JJ4WkYhZ/KzaFXGBjdxDRnbkdIYGGWHMlNdSSDlGXLoedJh
do/VX/UotttUshY6DKXjQUTzd332HRwDZF8ZrvVU9/YaK6kJ/Riu465bmzGS05Y9
qz71sv1BujbjIpReNw6tymnXZBxuGTxmeho4Can6sh/N++hRvFx1HtHbHF/zkXvJ
hMiDj7zBLTv//9/9EtZmNFbZDUSiiB4LmtTFPFC5AjypzgAxtfd6P5dRnKLmAnth
e0D4m0oDtPTsa70tkObEOs+MplmTatqoIHcKaqIEvmnQrmRvd1L8XVZkjWaoAJOE
0k2tuU6stdtfhVbJf7NUri2BC6FXqmOLqCAhR+6J+ROpztczmarN7QHvh93eYZy9
h+DiFN5vbP14Mg/HeOp0Rg5fvltavsz7n1zqf632pOrtLd/MzfYfim+P2aZXFER1
C0wo5o+FsUXKW373/4uDYncj61JHGBxZlalLTCx1Z09JLKU9ewo3sl8dEUYG0MTS
ZEs9kXxA6grjmIUDnJlWdvpx88ldWENxrv9cgCBv7aMlggwueLCriZkMlClNhdJ/
mfu9V/kD+Nr9NfoRMBQaK+zjYta/GbucUonYRW9BpAwbpLHP2N0Zj5LGtV9GMAkA
PrBNF05RUzHG+nODe7FbsDd5H5bLrsO9MOfuDeM8xwaYk7W905Hv8mg2p/j6QVcG
TlPFmzH9yKMQTzGtklRcdVO8//ipFRyVvHagItVTjFa68hPsJHWpWTPYo3h+KnwS
2kUF9Pk/hVLI/hUGqE9yhveaPWNKtVE8gr1V/1fUoRSBMOd4fnb6rZ9zBOHO/vh3
Qyuv00jFn/mOSCKEkby6AwAOdHj1c4YyURoWUpDFD3zcYhV6lUV2U15gWLhyZLEr
/Mo+9L0m2qtx9gkQVLtWOgw23G6xwEgIVN6HPzhLV1aif5o8WfYaXGUQHVXpZngw
W3Nro5ILOMj/S4REuatsuhTiwIffhkPhQfAL0FrE5Fx98on+UVbb39gSXiHVwz/F
XgLX38dmEw5x9TMWhCbq2bJ+VUghIQdo9dNWWwe7TRsGJWRFRF7sM1+MPBxUsTny
k8alPCIZ0/+nRbeGg20p8jWtbpYIZGGTKGARSDsG1NBGCaaQMzLC/W8/FIh347NF
vEPHYydQTDz3RRBuO9gQ3/u5hQIL+R7eLGjDDgQiN57LOqmOO2VFibpcVfs2Bcho
Ks8pAyYtbLGS41I2NN7fC/ZBasJq0pPJ93rXIcSIe2C2HlcOTNNFLQWFNEBVazl+
KsmbKG5XjRbkDyzN7WQAZgBCW6qarkdYSDHWv9c+QK3moZSqaqF+84ff23sdvuds
bHJJtub/6mQFX8S/aMwmmU/bmrk598iI04eeifNTOOjfCOaE7ssHSJZBzXQCsNmV
hDOhCOtruYZzfTiGNllz/DFFeDwmpo3925kGjpqL/mdPE+HSvCwryItmmFcgGVg2
HgUflDYpFIJpNXoo6QzMxn3DGj02GkWLzk0aBkdiTmiHak30gZ1qdmhJ2c9DsUAf
y9fkVpyOp8fvCpa8X1O/He9wd4UKTNjRHcVUTReKoLFLDjhEeSBY+Hj6dQuAsqg3
na0Jb3kY7hCQaGzfTntdj07DxUinjRBEYVFueV0lhyhqu57i76Z5QnMMqc39H0Bb
1DYOHwkWflHWi0iFr5do8a9Y5j9GWF6/0tcF3JPLz3sbqoC8x1a4F88bYodL13wC
PZ6tyDYADlGuERPWZA06OrMSJDE7vCcvSYAO6OGJg24M4izAsMtxy2KcEHZLpD6A
msa1vz8KMdBgs+3EHLt39ZAYzOFStQf1kWrb0jDSb2pt+46BniU2DtEBHqE28PIg
mjKpFD1N6WadyhNXfyHJBu+GTv5N8MA+sXLGvlec5lH65u+dnalvp5M3wRK7nwFu
tG7Tb/jyjh0zxYtUckdph97NCo3ho9IXtcIvS+NTJor/qnNC8CKag63guyzgWjJM
7yAWMCJ7NsFEyA9lCzcXXyeBlYKiXRQMyKhpDCdWmokET1BRrrrBqufmYuJ2Ledn
WHS4q98RpCcrimMwQ347ju99Els177ZTeNgXKu8/u/6MI8S6+NEbSntYG5OlBOi8
lWF/t7eIXL85kGMWm8CgsqYZZK9CqYPkx8D3kpaurn3BwNNo/cE6Q+CzW66rx2/v
ZzjI4Lwhk6SrMkgJo1QgVezUqKQP4Inx9NRD4BQN7lX1dXajEeWIf5i5gOoLRZ4W
A3RMj8q04Ih8FiadvEv7TJkrxKQyMQwF8sWTcg7GD1m7BwhVZGkj7eKOddjzCpFd
gIe//vf3bqmn0o/KS0vvw5ZT/Ag+FaWMAfGqa4RFaMTPSOHyA7imYUvf94ONFYN+
Xv8DAOveQ9vOfBsWld+CLN5LvGMycKWP+hnwKfgw1ErI9+B0/IInN37KJ+ymu4Bj
9EzemHBflfChCKKuuZZPWkPj2KZkHGmkfo6fqKtzE62ZJkztr95qgzhA8FVtTRuU
8/aveL0+1uFEii606BQWkVzJPqzqvM2xixoiRPpDp/PloS8YT6vaTSNQ0JTaGOmA
k5JLxEnDAn9ZwSdKfsq3rFu2iUCX1+gvHiVKS6zkSceoD3heIpzWHR/sm4QL9IQW
rtJl/uaHkzBiX2KUf43t8RO4GiQxIDdON6zh5/HGkim9ub+cA92SUMKGqb6Q4I7A
+0AHq4776h8RkZd+L7Yp2O7BkCvNspVFNaNtp8rrFm+4volMdtRtNlCt+83t8a9p
TpDKoSjfT1zZoTibtS9TvsCqVTh2NIoP7RaQipMVo/Rsb6+Mj3iohzhlmQiQK67b
ohCLacoGzgE3YH+3iiWgk5NQhAenfWaVITIazg3V2bSYDlXmmxbAtXhY+yEFVaZl
4jNq+BE/+uO9V1L2ZxdMFw9OMq5LDsgT7Kr3okh2kG6/atUtTTkgAh0mAYvzPPyH
TPqVGIOXk01NkguVz0BNtJXUPls5bpnXnAV19t0YRyHcF66YX/DawYkS/W/41IP5
6l78TjQZz99pEKuv07c5bOnPmrvbOgrkJOCPYt1MZUDWt+NJpafZ5oQWe0ZMon/x
B4wDliD1/a0ogGZKUFdrRyr8H1mr8iZ3GvHDmyzkgvLmTucK6ju2CNc1+hCwyRIu
nVrOqfuKQf5jXceFopW2rHhgSJJalz4CzPVXWRBH3lx9oSP7iQyzDzF6eXk7MSqH
CgFFlAvVaVNZruh1aSFb1WkdgrCPuK1YVS5QulPsxLD8VbzQnPVndE9StLH2E4pn
b2y+y3wMlf6ca9BHqjdPt1B8js8V5x1P9gOO9Kd8CjS755p/H6F0Ft/ufIY/VoeZ
6WkwTczE3oEU+PIkJHEI8Ox01ARR5dXliS0qMLQAR0lbtNgfCrvzMpBmyn1Ijh59
drN1gnjL2l1Nv5w9WI76/Bzh4gH7xsdVM0Jv2BaQ0Lc8Ii1nD9weGfz/oYF0ECEB
fbi5VoqY7McQoe9hgYAhZ3pkBqHHVHCOsGVjcREut+JrHZMf8qek4Y5PpT2bej6u
+2o9OWDh75xPFEpSVAATE/X9KHE5FBhmApBeVPLcYsKdaslRcY5+EqZ7TUHJRwTb
PwaYabguIrWURscruggkGxlTTJ0FjS7UEiPPO49iubS6UxN4N4inW8a7OaPmeZ8f
CZiA+3ofpZfWDMQOlDsouohNPhJJxcB97jz3t+2IpqYR1DJswbnPL5To0WyQh0cG
Z1cF+UB/VVCU+JVP4QcJERcjANtmoFppVEVg8h0GGGsB8UPzhT036VMO4oLwghvP
VPmNMgY519NeCFCPRmqP4hfg9E2kx2EydEHBz2vtl14sXBcQnWrAPIH+xSCQi3xw
EaZEwpKixMicKO1uthCQugEBQ5iJeX97eoTqIX/mqs1fg5S6RJ9blphDpEIsuKvQ
sdssxySk90l4Tm5a4L/o0WXoQqpFRRXoY7TN/UFOYA0aTUqNoaWbkMSdLGrFvrzR
06QdOEn4XjLqCznZ0lk3bxT1ng21WDG+PdTp04bhN95shqMhFHACCujiCeBQh/gG
GYd5TSQUr0nxmM+ZrzFt6XBJRD7I3ZsqGuvcacLevLL6HSRqTfsr86i/jzH1coMK
VjufMjbikRJ1p0JnFUg6EIw+T4A484diT39+JNmnfpJaVRZqVKs2V39I8Xc+TZ8T
1Prk5AGwj1NFExKsd1QS+Ee+rLDDu8Hw4zCDksdZOt2rHjjrtBv6LuE1+QhvsRz9
M9fnowYSCYQbI226i3jBaq+V24X83HFa+LBZZF7hMt3WxqMf5qOulokHhWYr0WEE
RvYxnFb/YdBWZXQqTB3Ft88ls2xCW76brsqwt5z0mVqx1DugyzedLqu2tPz/TPge
5AJyjphi9evGl5IQC+GzEw6gauQAgAqoMlJOC20a9OIkzRO9KDP+VOjhlqGkvW0I
dJjhD4pI+4bLRBHQLPqBysUDeFKUA7zBmirX2hnb2S/fPp3/GcqOAQv8vbvESfnr
1g7QHuEwnI9hUa4Bx8Y4BF3Yj10lP+Ay+uhny8ls6lXlm7VYQ4z/EYh2Kj4/5sxo
LeKBNcdcE0IBAkgFHOdc1bJLr8Kb6S5HXz3cyF5sB9gXcdQVXzXcrlrBvaWEAn2m
HlwFYwIWPAcLDLm/nturt4hfwjybJWp7+rFeHJH9YW/tg4ijUAiltgaajepy55fd
sV4EXKBEjqneuoIYsvpT9k29H08K+Wg3PLZzHWCWNefnbEr7p/jn2uv53V8XR9k8
4pp3/Bmse07jHiIXD2/KDu6frbL5F+aV52z0ZyUETV6H5fm+fHSGXa70p2wJscJF
aKTZLPlinF+7Bx2j251ePI9ybku/J8z08FslaMnXZU0pCsWgOUG/P1iPo3OHFZRq
VdmqAS1aseF6bQ4ybi2GenRrlmac1v/oB7qWc2PvQQ/joeUCT1g8orp1CwJHNqgL
JdJPEb9kQJhQkFzNrRAapdqwd6nUhYYr8p09CcB13uKiuieQsoooP7yi3376HRDJ
2hgNYSG8jSGXDlVEpIMj2HXaVN16YjoiZJcSUF48JhRk4FyLr1BkyX210dTKj6s7
CRqv46wje9NHsX1wFwIq1XzOnRAw5lnn0OQvi1Sv0OHVBAjxRFHIIX02AvY/G1iV
tkTNfQu23XT3JRAjKMkh3TAP8TSWOQIHR/4OtwrMvJpO1q9prU1S10IMUCdP/335
RKkL0jEXUYV684MdePbg9L862Ue0+4IiZ+FC2EKpLfv48iQf1/oIoxgYgI3NKsZ7
RyABG+gEXXO2AEee/MKK6JrEtmae8AtQzGw4hW8dmcwoVvCxCLKPt8x5WjmnOiUl
VxxcRX7Inmk5lW1rhpYCqtSp5mfe6xsHJzpEAEADhw4AQljPnMh+MsZruXLkwcbr
eXoWLM34oDX1riSqJGUTs7St0USRgAqLOmSrxRt8ZTjV9+gT2VAVTar3lclWmNVh
zplZCi9sjOnfbJC9RuTfmwK35g8/c0ZO5p33qK2TVpXjyGpSZEgjsr/Vx939j6nZ
C4jqsqPAH5VKUBUHBh3zHPPef1LWxd1YztuqULCtI47L8Uc1fat/hKyj9tJgmSHG
HBDEDDD7cS8rhtr5d74X8/IPFfRhBizjy962jyD3BaU/hhm291btNUPbgHmMx/Xy
Ui1Jhf/6PhFBYlwkuWsQPfkKb1szscdNjQeuaLnK8a/QkD7pVFg9ElWN3xBoCK1h
M3JBosA5tOtiCl51Fvvp3BY4koJqksuV6qiwK/CoM4Zuy8hHi3jbn6/zKD6t1e5E
bpX0Ih3VZM664y9XlAwVU+WYVf2nCouXvBC2cdhjHGmQzqJll5pW28qDJjA0W6vF
wiVKlMkeybTk2DgoPxHBP+LyMxEJurDAUFW63dgBxHAXfchTcB8sWYOzc1+2SWM4
AYZObnvfHV0husZIjL946476+2wwua/5Y7Db0SB0kj42mbdpfTZU9Y2WrFAKstYy
raaE2DwDSd1TbWiItkha3XxyLppc8iWGUQ8SbOqMFn1rkD1/aQQIBw4D8eCnjN6j
ocqtqC9C3cYw+omx7U83LVozDYvnFDyT1z+FAphRN/7qGgLf/nLx6h8NkvbsKvDa
Rd5o4lBUEO9lZFICpOPb07046jUzsrGWIKpOBkWnK055+QSfhsIAsDnVWeSk0zST
D7gzIfiFTwbo2PMgPeCWRYNRBVJxsZX8UHIIKS5hPzZPwR18jciYu63sHw8To7f1
dMOTBRVOJUc+821OeE8JFtQula688+pyKrPY/6jSEz9LsLgdxJ1KWWuQRy89CTgN
wIi8Hpr47ZjR5CrWA0OxrEgCE6Agd6xmLVXbgfAXaWZ2dZTVtZGOhx/ylyZrteyL
dRkIFafTCvfPiggvNy6VpTLetqossJicsLhygCNnrg90sUI/ntrIezQ4vjHYLjlq
c2O0ZVjADX1pYxVIdeH1dOcEQ7UlFER6mRQE4piqHrZZV9d++kRn2dsaPk+glpzr
JDPc8qtXVuZARH9PfZlvwqktagrewqNCmi6nI0FKDuHa4r12GtqGaWVlJL/5ftW9
NDtiw+fSf8p7dR8dyd8qcFB3QhFkNMetUoW0Ukk9HEh3IgYTua0ZJVazF88/3VHW
ebmxYVOaXhN5zAQjMdtEz1ganqKba3YegZqu18ciovwWI73n+fKbjY6l62zuCt1f
ecg0Nudzu+UR+K2aQk7wFQMp+NVtKzm+0Ucy7n9ApGkv1rq5Quq/wYSOuYjmr56O
x6kcA3CCMVatFts+G4VPrEq24kyZQPu+GJoiaK9Hx3hrTH8hJueYdVAReDVGpU5w
YlCpdITfcRrauNrb8iuVsm4jOvHhAOaKcrktEYSPrFzPcB9qFGwQ/O21HW82rFXb
TtVKNUEkFJbpTGHpOsTmozW7ncSYq8HTHmbPBDhzEAjv4rRf8T9ECc5c0MuieGuA
Gd4p5nV0OFi9oxwQnZihW57GdBnEHuPEd1KBj5JrkfRjdKavsrp8beHoFEzhk8pk
hwjHpEDxIqD9KElFAYVU/5lbYewM3Tugg1UvZRVaRHZGEibLl1jkPv0u2aSA1Jke
GZDl+c6ZSuBcpKQHoPY7PFRDSILsQwd4vSdg4Yg4h+M7bmcgc9x2moorfnqhvuOU
31pbzs8+aJpn10Ni8EixZdMdF8wych//DeZjk6i0MRqNH/8xytTjKTpgUwBpgAg6
y0y/HRxPhnYV6XJV2eYLmtrJ8zqvJUVl9Lx/486Ml89AufTHXJSrTkeneqoLGrG5
nizrNpKUuOMaHO9hz3uZuemhAupeEKvchyLwpd5cEJDJAR6ijU/qpajfEj9sSP4S
Y8JexP1SYbb1tktTw0/kQCwUY0jO3IiKcA7KEQolWynxWqmBpXANKm119QXMkVRQ
3IQMrnwDBlDJgKGH8lsm3RnBv15337LVMUrdgHfJse8q5wYtgNVRwwU6rwAclkfs
E8decCGWFs32CL3PfYDbrg6nJwepJ28fZMWj+668LjffK2leTJSpvyyFPDY4UpFh
/ASfEaFa+9loOcuWOP34lu61+Ac8KZ0r3wMBvRkjFCHjaJsPou7ZuflLLnf+BtRh
psMJtRn4oqWaZ1Y4/68zSKmWAbnGE47IKGF1hpXuyMYvY6UbPpb6z778ipJLrYL+
02F9CqbwIGee7OaLczvt01pFL6UWszCXfq8wzc/QqAdhdLEGpJw4LSc13qtZAQBA
shej0sLMRHL62SryMzYAippOoTXb/vkDg5o8HDwcVuo+E7rPrdASEN4XfWl0sorP
tGLBFqOBPmboHdAIepRHChU2zJtcsfGnYpc+6nLdOHrbkxLuZ/UsFUEI6vSHcMh7
QIiokFGNQKUKei9dUEycrdZQQh4RdXAbB/CG7iYUPwdd253+wk8QOQDYQtnOH7lv
YRVeOpHTqzPJp6BmnqVAXazYQn2g0O6yV2xX0PhGDLO+ALD5ZkfrNv2W3scBFuIM
lkXNAtJ/qT4uF36UMAjgIZXxrWbQkJY94pHkiwq5VT/a/eLTN/DBvhw2E54qQcKQ
+VaSCLTQxCOzbmPNX1gSdek+gd4KDYW/lo+3DtgJHxp2jL6UgIX/bjEHBwa3eI/p
7IF9H+fyoxA5IbKkyAhaepwSR+xR7kQDX5siQwXs+HkI73i3pOWrNNjOPqi80fFv
2B8WcX/oYQ5CEPwlkzuFu++8SJPc9Y1XqdKpOs0G37z50qyV+1PC91Utt4rVupAu
ifHIRjI/MjUa4OsLAvUuqFqTLYWADwt5yQwnJVRShPaWu9kLAY5zUvslNzlaBd9M
59OIwEr/PQPHJuCV+aG/eDpsBDVHTH4KVpvtfu3XRZNhCzaq3oANKzROKV453XlS
xEQYk3A0cDdm6YFF+d4F2fi1o6H8b2AW3CAbiN/DzmbhV88lU0RexkHGDLe4o3Bw
Wuykht+WFkr2caAJcbXmJHLqUQ+smmFzZO6uJvKVqoL1suGAUYBjk0Ad3BWRpjy+
dqG9dGb+DUzW/5xc038ba0JHA9kxfTJ2PCoOWlvYb8a0UOYZdE58Ys9FlOXABCjA
Fb58pJVc6oV2x+XyvjlJsI84LUl+l4Yt3LWQVugCT6ZVwLRk6EPDzKPAz6TXTjQj
4bV74S3yFQfkI5lc5PcDEVU9A44YjbgifDdcNMh9r1KHHPXtZHv1AeaqsUITCtvN
fWKV2+AvMjqEscWY9IVqFqZqYn1wqAwy+iw0OwlekvXpmxWfo2w3dwUCzYSXG8tR
lgWNoJ66oezSR9UQ+y6y3t7QlWmvSOYCZPSrGV4HKuHgjs5wFYESX1J/lz5NvBZ8
XgYPjPLCiygxmk9Rbx9q+tdoPVoJv7owo/Y0DpRbVVhhGkmvTzcml79d0FVMQX5j
/ASi6dUXidpOF+429OQxI74CwCanjXOGH31NYZG64XbvH0LKaabK4PvR3u+H2ElY
wDgOh35sISQ597W95tVUeRzwme7bb5u/8jiDBUjB/eJlPV/Irw5S8JCDmiviYxgZ
Ff2051UlI299DYiLKL8cMBjP8fOUfN8iBgv8O5ZkM4e1Xkuhn8LBohyPQFTn2zQm
1ayUKgLKDDQjDNOGcxv+pwvUdMQvJPrIGUlpE9T5Ur/E9qtU9qRe6chwW0zbTil9
riCRQbzlH0aMj1sIZk+JDLaBTO2zN6XCEQVViFc2l/sw0iMu+9dhlU6jyffXw2y9
hu+QLOwfNoraEFMf2Szpwf30pT3y7G/Rc/EQe+mpP34Scoi6dkBIU6SwD8rfEXf0
mXX00mih2fkGFT5Kh1iXSU7TOX+j+rUpIVBsLmiDv9/iltftWA2UxNYVw8hazuvD
Mos1DHKVXDTy64VzoCQn6VUhSDpPv3XNEoTNNVlFEn4gc1F258TOOYrbWz92CSoJ
OpggV0H8kM28heJ7Be9k5/80Pa1d5nr8OcbT2A2pNa7/ltgzQiP32vbOKq1ROqmX
hTRz3t/uVPb3o61VuMznq3QCH+gWfyuoTJNtDL6aUVE7PFGKPINtlk3KG4Kdv0RR
LhS6k/plZ38XE2LReUcblrLjFSIo/Gzij3EK5ZDaLkMpI6zpyt5CZXAbiJy+9FrL
UljIXwUC7MHfgYvo2canwTPTZbPyYCbuQlrX/xMJIecqOtsVpwxQemdNknnbv6bE
7tR/VpSHW9TVpmdoEC8UEpOEmKkThjFxc75/Ky4PJRO6ytLFRbxmWPqvBym6rKli
aUnvgTv9EDira3PLohYOBPlhSMkRybkFHGQdkLbVIs7jS7E6Zif8JJeEU3CWUudS
JPJtVhwWAHIbUNdh9on+AakYk/Qb0Vb27B9AEOHsh3nFSH/aBJ2PVkxOIOAtv+s5
Hsf0Jr81xrxf/lB4k48sK3bs3bKYcz7VsA0ZNBbWGrUgVTfXIQENRKt03zSr6/gF
8J0hYAHlVOaDXpTKzUE6ET5l5713HXkosa+XTYKMRQMYUCxCkgTv2VX+p1/ttQDv
SQDaGxzVu2q6o2XIbRf4ti+QvD+jhznE6LbhJAF+hyYG4Qqe7Y8ya+d/CuJOzwTN
w0iYskqtUclkKRARzrDZ3EtBsGwritWbNPFSCYoAyphrQ2Wntim59oi8j6FxbWER
CJmtMPudQ4qcJVOVVo7IHtrBxl2ejcH/FaiU+OgqMzrD55D1J3c+u4OLFJBpU1vF
vj5NYceuAw5Hb4ZuixZaGIL20xrM/CKoaN8yDdPgaAwblEveshvClR1yqVPSMq0V
7D7XErNn2Gu8QuxNkfaroSHeAfc9OUs1BfLnI/hnPWIqvQA8bGi0CYD8ix1f747f
wD4mxK9rpYU9CF54eJBrDf994bV+wIEZ6iYINL4IKbKiehwrQCFKrNcLWxvGPMpm
hHAcEkn1NHJxm1gwz/wLdwXriFJsBx0AxHAUk1Z+JP5b4OVwOap8AlYQQPjk4fO1
Vq9yHi817lefeslDOMi38IGQIYQC1U3Bk+RK3DH0/Rb7/Lp+WAv9d4trx5/a9z+k
Up/XVCnUBfgzre+assUkXPDe62WigVxH1cFP9jc+rKhLT/sraRWcMXoSA/FK5rSI
OSnb2BaQuSdh6EL6z7Ij2emmyq0Wa4tZItYfH9rEVTWd3JlA8+w6Cg4dzyHxa4hD
AZq79/iCNNiJC01sRM4O/pJwGxbo4s7tquHg84Rj8J/toVNf/NVIPs/DCcCRqosn
F2r1FF6zG3okIchSmekNDgTsYmEvfdExtUzs9eoSwzW3o5F0XBXqwDfDnVc0zWJE
KhDCejji66jUFLAgDKu/Cg8RTAn5alg93bTxkF9Nr6ZwQTLPGUVIH4g+KCUIIXR4
9hYzzfoR68m42XTjriDtb+OBAIlBBWqJ6Kz9RIFraJV7ofAUXoqo/kLRmxafkrvv
wSzatKGfBmd5wW99yrwNIx5YErw5AE9k9pN9J1Sydc7IDJeSevLGGicNHDaSoi9w
xtwBqNxNd1wDv7vNc4oOy0KG6WneBQLjFOA3nnJRcp/41nJ1SSEKzWZwgPbpiUcc
S1Poz5PB/mWMkWD4SXa6GsQsm79yZ+gDWHFyEuWG8T1bwWPZD4xVQsR6ZG8N46zb
N0I7ZzDXD2lyt1DdYV5ijf5Pd+IiVjVQ3l6h3jaQIj+uRWgbexcrbiS2s3Xz0qXk
95NN9rHkr6tuNn98zoscnqaK2XVz/QixSzjxR7DoCGX6pp7ez2mxdGJYsI03Ls1O
DH38HEMFbNIL/0v+KKlzW3K5C/yNMAs3Ou0NBEodGkdtG2gPBWEddnjAZhCNVZs8
lSB0xq849YRrRu6Tio6mVNfaKzsweqDeaNWG3fpJ386pc+nuqRGr4+US++TJ0ZXK
uA5mz4NI94Tgm9VpsaKgLE9IOPKkef0D70vE8fB8EmCUMqrEI/yHpxQPNuvhfuTq
JFOYam0bkmp+DEyDjJGmecCO+vbQXbBn/4/eO6hMjaUiMlyZu0/b5rI6MFtRyxnm
cOGReGA6wkMattaPfJjuu7+tzBOmdbukN4IjfWty9tQomDWVuKv5QWC23xU6tVwA
8ppsdFwonCeDY1O8zx3g3EDInw5ypd8Uu+J9ACOpok6Kq1Ux6iOmav9RM2pft8AM
jZrG3nnd47mmE0yMjAbEwPi/E1s8S6A63W1FmQZHYO9GqLDY4Kkjeu1lZefoPUak
JaJOXia7rtB3UXOUyU2K6xf9Mn/6QTn/2NZdnUCEiVCyIFoSVqsYyCeHZrKho1oV
Ts+c75tKtP7gSF/hH1kGHPJmhErpxSPtQXYC8nY6qIwq69dX8D+ThVShGD3wY+BY
pimJsXrJm9q0Ze6okI0krMt8fUjq2zFD4gBA6YF8QqvHhVLdRzetUlX0YfRrx0Fo
phVuOaLGD9HkfG97gB1UyFi0UzriG1LBUnJqRFQJM2lgpkX6ByprBne0hJBdVDkn
JPCbyBVcO9jFoTBbiPdBiR2lQwaYCKsx8LzZyqElXI+T4CxHgcfaXaQ2H7B5ICxH
ajZXXEKt9yfHN7cTw3lIah7aAfbLL8Bg18e5uCH7+ZK3s6h3VuLpSVqOqOJJ7yWx
eUEdKAsAA//VtZSDsKnc9o4RLZmYYUAEBN1hT+ib8TXqMmlzQrScTOu2fJ7g2Ws2
PGG+ozykOvjnVnca8T7JoSXjA4PM9izqhHE9pOKSlrilcmQqGrRXAlh6JgFSwi2D
wieEk0F1ip59M1XGElPRRBhaOK/pW7ZrepyQNGf3EAfo7wtmVGb6qQ3wLGtfCbk8
l0DUiWoKfbgzKsxdXX6dCF6CCJ4FNup2PPnXMLeaNlGK/tU7y1jlBYmfmRL1NzpT
+83mFN0IjtG0LmYQRHOskJQZ8HlqyJJxWALmxkc21blqAuKl7qekoyHcNE7wE7oC
HrVCirhtNTAuitZOlI91F9ieI+euseQQouDtPwWPeeI4gYPTBAK9DQMa0ISB4Jtj
HWrGztyaZH0a7n+h9JJg66WhUkRqeh34KPdEQ3OAhJiEjfyntt5IGYOVgI7IUzaY
cixPjg/oFO6z4N+hnRqEK/GLq8TsSsu5JnXqUtReGaI+fLAU4ZmZdBzujL1hVJoT
5O7QIFY+AUXBKUR6oCh85zLvNpZ7NsrjYMvgYyNLfj6JSWHV0jGYug+u3Ki0MctM
QHHKaKFmJZ9owUtq9gtNScIJqhbm8C6pY1o/6W6LLxSqrTSFcVcKEXAuyPXftETj
QUKDIXtJcL4dcK1TAftes8AjQ2S1hly2/wP/Hm4G8+uTzJQkeAwkSVreabANR2Jz
0EHwvo9VIEKb6fMPy88d54Hhc9Tvj36cuf8U0HIPl9Jl2eNmrIBGlwjLW49r5Bkj
nIzMD35oOHRIqX84/NlaTVd0x2imzPQsRCW3gv/6NjwTbG3+GwHja8dTMqD8+JgY
vgNSGc4yRTozErVqWZYidp9LnXbJKm4WsA53qTIzpUTTj8Zf3+dDXICR1snUEi7m
ebbXwrGVxpRg88dDc8GL+qLXs3cSLM3/031DH55zMCVj7r04wJIXTzJSLERj9evS
4aegWOvRjk6X1R5y1SGG4tpsMSh/PV/1j6PA0YdJnSYSlBVZGGDHu+/YL/b2vt7C
MoK7mOD2eh4AJweiQQXgyBsBdo+xMKU381Ya+5HjvOF5siwYr0AlWRupkiirgz7M
X0S/bYvUHYocAbg8sHcevOL+f6OwB37TczhaFyR2ui1QwsbgI2D5RYdiciVW3qOu
c3OJePqSdSV0X8z5HPBt2Lc1Q3X42Z/n/XpCldFcUipN9PfINDuOeRYwjktb3lqG
oM+kmBSPwWXivVt3ox4vGMH0JIwC0K1mv7eNEzMa8epS1aSu/LsaOOXYmhmGsr22
2vlZDNrgo7l8bCPqTYkAMo30ZrAKqGa8njOchjEuDB5aoTpqPtMqjwCJ+9HKqfqV
TEHiIDBJyMP8OSIkYZVnM33ZPoqTYdV5cEgOZWcoMxBZrujd/Nlv4IvBWw2sMPOU
R004imSmb8eIDD1KuG+uYwJpM/DwHp6PnT/llPx3be+RxPRM4lriJyJLaPiaBKT4
9oltIBG1MyWCAdmai9eCiTanwAyC0xfyp1cQBIMGTye1hgrNp0RIq5N0VKmdKkd5
hRe78tHavs2Baz6C3dVes7uEUajalKna7S5rnL6WtH24dUPhsIoLLXn84NGNrTmF
/2WPumbOjOKpmP6XCeZ3jUEIbOq2UmRrK8CrlNstv6N/iMU1DcQrchmgJcZgg3gU
EemJPexvd5s88qGaJe/Xk7vUqjXCVK3BoFQZYoHjiMc433a9fgctMyIelgJ3fZ3E
0/7vHA9ix4arzUFg/j6wS/c7lJweJtCf0onoiTJ9xw0/rzd5JETcoNRqs0KW5CBD
ypQy3gQwbY2oU8UPCP368vJ0rKvR4s8XeYl7TLxhsanBmheXSSG5f3aSNbokabtg
gvPcn/Umc7ZXiEkaiErh+I3uZnxYXcb7P7qEiLnLm0qZgHjblnv5aZYTb2ssjfCu
meBE3ZSrZ9WaJ0kDh9ho7OZEfGlP1pI9WTk0ZmEynL3DOjOmN9bUX3GPsqUryFTm
uOXimqrUoTgplAuCYqFAr8Sqd4c28Qjl76eFLv+Do6sWJ6sRVqnPtJsxArXsgRw4
pUnt4gHOhghSglZK1Qmg9ixmsLzN9ldlUyciCBh4YDFr9FxwqM2h2WriZrS8mekt
fdRVsJrQpBwqV8DTlfk8s6BwrtpXtV1eJqXr3rPBuvo25hS5tNh1yyXQ5d9UWYWm
fAl6bxmzNi8RoROokfheEEpuf8qgGLyEMMDknriQR41rwjbu1JyPywKF00S2dpaa
nb8w1argCmHikcqCd/101kxdQQK0KAbvsU1Q4fcKlsWByR5DY8nt3U18LZ7rGoEm
rXv7Oft+pBHsyEvXKK8GnI5sRUQCBZr/+eYaPZIC2lLIBGN+HmBOxwdfypH+toqW
qbuFEz1loJXomfqm4CSBOMLRmkmiBn5xvHXRh6PHWSC8UbV2EeYF5nZzlRRfnaY6
e9oorJAEVxyCpWFpbRxI0W89+kGHpmAkBhaPu2VpyxX/L/N/o/2Nh8wkymciBglT
2LZHJ/xVykMY4BVdLg6rI5BpEYI/G+oXSgY0b9Ih/5aknl4OPoDOPb2I7q6sHrya
yAK86KMIushW/eKZ4xsyLAZ3fgI/tNqqiWDfHEp6PX9wiADXQj+QyQ7wz2QXdV/D
6l3uLHBsC2AL0cE6oCHXgxpksWHjQAAYCch7HTqMm62in+qiDeggnh/HEMZpdCLL
Zzifu2xotVaiqKgPcwXO1W7CR3ZhvSnZeLpzy1Rtm2yjiG7R0Mu7yAje4OShcq6Y
A31KcUPX4idnbf5fApwvrJ8Ycnt/2OEM4vTkSniGg0OplStVCJRsfaNsX/gCpvJV
xm/MbfF601QJxLj74NGSdmxOW/Jm9ts5CC1ccUxF33SkJHid3MNzniYgD1FigM9N
TEwJSyayDMaOg+mYSxz8lyfu6Pedh6ymIupDt2M67i2wOa4XKVSCrc9VRgmsadnY
1TPoqDE1/JUYta8YeiiyxOLICD90rTwASVCBXCUlryvut2OGVqdS5bjIvhCskJT3
HI+Tng2RBI/1SGy7nM2l6mW/bFC7557lBETJhb+IIAkkSI/LWmaQ56LOicKm9kG9
/u+AiimZqvz8uoiRxXix2fE7DBLQvfaiPLwVsHaH1RI2pLt/3mUxeP8G1ETtETNU
URDyDRWPewNf09cz7cjcSX4EXH5Eo1zSPbQGWiy0vr8E1PiMwGVrvFJ8cYEvM2TP
MbkDsSgDOByeMIMGp+8OoFoHSBkEEq+jX8/TAdz3q1S2EXWfWQEwVYe2Vp2RF726
aT3QcmmvuK3kVI42aqBQoE3AXbPD4p6yaWPSKvmtQxBi97rXyYuE1OFu8LMoKpVv
RVI9L43vcVY6nxcxRezGHuYC7aZcTCQGuAzbdJ8DX18h+jBf/GYItXyTrS1lJnBp
DU7SL77rPEvXBArEcBuxlOwAh8cfTs12Eq7APFCNdaqTy/mSFRXmlGl5tdaWwH6X
P6/eu+N+Og4XS5y0RYhvLex2tnRosbkOe5W7wX3GaYdormE/j42gbn5Bn5XLmHPa
U1MijwC/wTDShbH5eEe+P4bvfUEDRmhZePtCO1oj6PT9+4OPDh/fE7nqnhw/sKOv
VxwMOGg+YHvaNFiIbyFLB7tKrZ+AI27Qnkng2/HCF084c1I4Mj5DEgyzgxOfSzjb
yAuKm1nyp9q8aCq8eub/A7pRdV1z+oE1gU2UZYomPYW/yQ7GamAu0hhzAoiKA3uJ
LwirV8nM8q7YBICJ6YcYiQtDP4KmORXSSveHoVWvJ+tP2BtiT2fzz/dlzLasFqHG
HDDODMhO0GzKopseFGdZC2LgSs7ieDU5J7S9/Yx0GbYXiCPwlo/wxeMXhdiX2uu8
uI5XKzuYLCIEynvIXtDcnBYr2sFyvZA4iPEL3orq77PbV024da1FxnMiQYfbjoJ6
LU38s/rqBDXV8BLV0MWZlRgIA2e4pTk5bcByE0xoXLnjhLfox7uzCmTN0y36x+oF
JvNOHOrny02raJTqIiLkkpElLUsg4iB5kopiZ4mNNV4SeXVy7JWD4vQpy1YXBiNf
RkAg6fzTelPVEFc6hnp8ouAZkGWt3BIvWPAuwNygi7FUxo8BOrM1wOh7nXBluQY4
iygv1JDtkEw/EIcEKJBQG0GClMQdhId5hqWIavRsHoAWgKdWqhTCBsfvlBES+ONw
e0m6MdnEvoe0lw//5C4+2Wy5FTonct0eOtWnlHrRBYa3nDwgXq3Lls9MSqLGOSE1
r0XRRendwBa+WjUiWFTOc9Inmd+LmoDjE11Pap245yICRxL1jpv5QfkK+EP8JqCl
8ZqIa0U4gk33bb2luTcu/GFgfsl7hAR4MeSn09O7ibUfuMM6MsHRIwQBMr8Sn3o0
bIbrs/S7iwNyINA0XrhjOBFvTJKlmDzTHAKxncugLURrKNZ59/nmvfPToilfbgpq
ya+jFwQNrsXlTz78WXGtTSGuI8W00pknlIxYdEL0+MzM8z9qO8Sn8KA6QHeUSR8v
kcakYXHPhfbu7Stmlpds/5+waVpbE0gjPWqN1KFovZ/OdHq8bGlaSLLFaTRajKpc
VeLR1cLCw+MpbuzLeryUt/Ysxefe678iJpc5a58fLalQSeZhvb5u+Xm6VqnU5L5V
6fBcjgmYdaajw4FFLSIlTwSdx4O/IyQVRWb9P8bIsdsrGyR6DN41osIE2PnGG1ph
wNqOW8yjRKE3YphwZvyoE6kSVpZh0jUWm4dL3ViiKUKI9kRC3MOFqd8TDmtlhu0B
3X6E+XaXrzA++PkzWotHLH4Vk6M/SCXM+Sv3caI2cP7glEzOWggt/zkuJusyAHsF
YzJO/Tl3S0fSrP+ZSF3cfn5mk43/aRLJuZyS4Pfja4IGYGJcbiysamhUC0IQGEKM
bxqCn2XbFpSyJdYfyULxUMlp79KagDV/Tjdngs/CSGaf4dO5F7vjkQHXBdoCtjaW
ug5WPlJsbKRTK+Bhmp2taiBehLxbDUx3hLZE2QIsG6vIRm1L04kClWGNW/uk0tn4
eioSBkFTxnNCnVjKGUQokT27eZw/jGFeH7qrXkZJ2BmfTsB9AkgBiYqOFFmPnsNm
bfN+LtUhyYEq6wvEJOrsAaZwtLkujknk7Ibts0Evmcs8W5kN48O51Y9uE3C97Fdj
x8ZqevMOBnxxBiusIfdVXYhWhwHH+rFe4L9iQkSkTZbRsdRNrst28A0Klqp/qRzL
NXNNC/FqqtSRSYZxujoKZEb9OlqsB/lZBK7crSCb3zEfz04a85tyEwLnTWpxHW+a
VFZ+0HYFeUeOH0CfnOiPb4XexB9n8cPwpsi0xgMdrk1GsnfTpZyZcrCCheHDSxQJ
FeJbphIpeKensJEnzVx8cXDSqY22ENjejFTqIS6cF7ZkppkefKXrfukOruZyvOSy
TBvpOApFULuJpT4KgJWyc9gjA2XKCNb2lv7Ac92EDdGSBWPx2+QYgtAwIIHVaYdi
A2tuynVNUf63ZzQs/IDRy7m/gVQn/tHUNeBM4lC3+S5Hhl5p5EuW7xGr9+U6B4pc
CZJFQ6qTC2uztfsrf6fQMKOsBvBCnXmJhTJD3fd/u3lGcQNDoYrdsPGPR7iwv13W
u4FzuVlUrQ3UgQKH7Q6X8JMbZd9pGFex2h4vU3PSrozWS86JBhdnx9Pp3I7vTbJU
uBXEas+P9f+PXQjowBfw6pNRCzOtV7wi3H/Mzbwmp9Rjk/5UaP0ZtFpM368yrL+V
3JrT9SxwHi2AhJxUnJ8pRIpIq5aHkcPB0qcEfR7+M1mi9gCNmxfmUDfw8rJsrDBs
bkDPRAm8jQotb9NeV2VciCQWm1NnEBHKbMfNrre5F5BANQ9l8usPeIVnHi178DP2
4iQoSGhGRwvNIQEfisfn2JGuqAnpXbdiwlCSJcpIAXsGHPLbUtxFDLiGvcifLUy8
eF224PbSOJNwiqulidhwDdekYC/6NlBCOpKW2b5+wYwX/YOPkK+hBxKuWVBoyU6y
UvdGk/D6tEpEymkgBT76U/oVBNhlZkiGYdHB3GfAQQu+RNi6Eq+Eyx/p0G+ynSCF
z0kBPGGbTVYHNr71QvnYBYeG4UQmMZQlGnvR3yHbXmfqIciBdvC173r/vnhRqehw
oY9shGyJ9VVrmE9W1rh0nW7C4Awz011rGCrITGhJIP0qk7QpWagaG+11rRCNE2qM
mo81sv1Y8flPShuMYwto1mZdOh7h3pjsHOfVVfM2KzdaRTWIO44iTj4JaVym8L6f
fql2qOgvg+b66HWZuXszBwOHQyqPZNxPGEKQl3G/bf/WM36wukgd0YOc6MX69/JW
t1IUgqGeFobz+au0iFrgC+P5b5AEhSArc+I/KPbk1LersdyJb854pnxhLcCFiR8h
ijEBZ8dqlFw075BmEBVc1Aotp0mrVE//4ARxfo37E+Oz3FeZU5JRkI8wzqsJxTwk
r/qfALzx/bhAyTmUp5OmTxZZ+h/kuNgZYxMq/CRQM+oZ0JN+TqvDvs/sT1y8mp3W
Gh82raOMkK1EWm6C9pg9K8RKZrZ7VBAAKsiPN0qadhhvBi2RGmXduqtQQO1e62RQ
NW5DC3sjjkoix5RgxdUhOOJE4gqQMiC5UJzGLcXVd7kGUwXcL0cpk+GF50x6Evft
yos6aLl+kA1l1W6HnLkbxsKL27QA7sO5Duszpl2q2FbSaTByrGPzJdxtByOaX9jm
p/WLZy3/6jHG5qtH0K+ni2EPtZC542t4jSZ1ek16pUK0IzdWyHXC2klh4uWbTvmS
yocsY5Xdx1RtlDJPuNsKNXuUXm7mgwtGChmfTdIbnZpk51IMbyvSrmwdxAaF86Ei
8SFTXsN1/tg9BKqVOMgO6RNk5TygGiMB6e4qOEa7NuG/BW6INObtuLkvLNlqUETX
mScEG6SprQpayVDm5zjBn2dwbwo/vO533JrUgQAHFC/m5LGhrULgMiCZQEPmCyT8
2036ePF8RAx1a64CHI6ntk+5uwDz2A2HQVaMIx4TslnNpmMZ+WW7sP7WLGv6QbcQ
QZ855RjBpVbbONm+CMpbCirzYPHgZw60AL2uxjGUDm7yP67EtwwzK1f2B86MZX4F
PRU6b0bZOvUT6k8h+zJm/ElfyBqNi5S+dhPZPCQ9pTK/p2SGbgnbWN6odh2uESHT
d4CsX8o8tnCq84Tigh7g6dZXym4dDMXbryNGDfdwGJNUfdFzvE4xqKHtujXBuB6S
1dqH+lwQGdVeajBUi5RmrK6bhoX3XM9Hr5F+czZ/IFGwPTslbpHg4XlBaIAh8GHH
DJxgpKCtXDAcSUOpIyygfZK+wkjEjw+DyKh4p98OyXOSahFx6jqYpnNS7hNAp05+
kBUrikIgAYFQCJznqvFEs12VYZCnzjm0bFCEnI+bATijTHl/y579sqIS+0lZ2qgZ
XKZpvJhNekfr/kCaOZa+s1VtbQ6vi6rEgaBsKH1XB2VoMPbgCXdrNJt4IeQe1AzX
gHDpsp94RTOF0blqw1HGVszprDlTzNyRtSJy9JJ0S8VAc6ARLCu49hSLawGHpscc
lUm25lc2mg4tLDG93277XwN2pvpEUxBDjpvsoB8FC4LY3S1cpQ8oCmpGyz35PkC9
tlq4oCHLNBpSPwDHS1FFfLSOGlaamYihmc+pVwGqK9pzntj2VBywdtGNq7IPapNA
uG4pjLuUKcah0QN+78Qy2PoRnxHx4TbLcVRsRwm3t/xZnB0+lmfcmkQsfj2IQ4ps
WnvTJw/yY2FFpay8FPbnjLJgR3HA3Zb6V8KT7fZZxR+RGNqfgGhfc+TvjNK/r09s
aTs1INNOhrx57Iz3PwDQ6OQ8xxyNk+YpXyOKlIAy/+BBcaruGePrYANSm8vU8Gvq
y+EySBGU1/xfnEXmvk1lk0XWACdVR2vu17fLIK99nIvyZIZ8CPQPV8D0ryEb3O6E
csohPfJqQhPaeMt+2jiBOy6qu9XmzyegAAy2an9xNr2JD8mkkjddWZBXWdGvZ3/A
aoocnIs81CLun2Qp8MGmwLFo8+hkcz9m/rFi+KRBLiDUZDZQray2AzAELpmWCEXv
oG2pf7X8WnMAC5cALeJQoDpf6LEc4ai9XAASPgOeV510kTsawh+tD6GcfhBDwDvM
9/3tWq3eWqu6BusgriThkx3WUZI9BTTc33IqLNLVRf4eUMX25M0/LeFMSZ10vO8u
Mj1vg6E0iltZbmkR8G1Ova/qyhLxxg7+H70NWaOAalj+wrqACfvI4W8R/FOIMKku
ZvmVBk/FiYlCivwmfSB07qIdd+zT4jp0KUIcrP/NWWullhhxTdkZx9h2dXp1lb5f
5PI1bwYSCmw9fWzwJBGgaE5SyKDMckpNLfmy/VXO/ocn+9V5Qa5dhWuOz715lM7N
cemAA5cQaUGSufsvRBI87XbFDVSZl6cjKUXLjw1HBr/9UQjuRfcb9l8lN2HJYLqD
ez1U7dnNla8qagTcWniGrfFVhuOaU24v4ViswEotNZb5pRvahvj7010xZtE+PvKX
t3KfDVLiQFnXP92TDIM+rimvAK54ztXdmSix1vWMsz8w61irVli89msmfnTLqkmJ
ARCdNyEi4sfFCvzmAcItq9lxz4XQdtuqhbFvOetRl8XaDmVzC0IT/H1HMmQNvR6J
tuJS6jG+nIha207ucEiMqTPREeFFfl1xwW+Qs+TUiDCPg3DaQjRi5G045qIubdcr
/EOdnTz69QZv0CpklG5b2f2990+bzaOpKKpQw/5vPfv2hapzMUx236gvzHHsxUfu
rQTqRn2fVdjDVaHKqVlzss8HoL9GOttDh9dxFswvKlC9CaKhEy0uKN291KqmVziX
dgxhel3lG3sIr3HzOeTjyt7vYIez9haXzbgUG0xU3LwtrftCZHBv2xIW6Sd0sR7i
ebBAaxM2uFP4y34XFkEoM9YW4DIqOellUdxSbN7rvz/zPdrR9yq20tkFY9nwZkS6
GoOuXgW+jxuyvw6nVk0P2FSxEylZooLfXHwVCMlKoOA3yk68p8ccT+zGT4denUf4
XAoMvLH/2erPDTqp7TkQTzYNDp79XLyqflUKlzGam6Ms+Qd8fTAUeQKrRRHgM3n4
NXTxxpA6mLFYcr6w4oZxtQRST7UezKnNhPYNjCf8Q41ERuEb4noh8iJmbgJr4ON9
kMhvvipOGUFiyS6qXBpjPE4MkorBw8WIXJCeni5Kgvk/lZXe64JlrmOmt1d4xYJJ
tKNaQCLe3ZIGt1SoU3D1Uaju0lWak5B3yI5CQxCxuP43Qm6XfB7RzQwg+y44m3TO
ihUmyO2/SsRx908udMiHq5qqIOO8Z26yvUh4AFeQQ7Df7EHxUP82imuOkAk6L6/g
2mSRjrXcoeXR8YeyUNg6lwgwTACjVXeVWnh9Yp7X1lDh0GUSDZ6B5jDEFxF1PRVK
8rKNfoq17Sa7TnV5eJ+vSWvV9LwuHYWkwFiodhzwJ21Y3T3ZM5zVGd3HRr0okhWZ
yzFqfBZnEibnRoPK9r/BB8adrae4s/ryyFZO9oHCSWOhu1Z+2SSDpq9jbtXMly06
N0Jg23m031+CFKyBQDErd9IUCay7LH4cF2E6HFR9ZF5B7BAglSog1ymRE86z2d9G
r0xuAmD/YjhGhr37cBdU61zyZlH42uYwFcRUctbN1m9tlJwMxtpIzmKuykozwXab
rpi9rEvFq+0x2haLv62dnz3Yxp1CplCtv6CncZsTCPFqmn7eEuGerK0B3xuVvLWn
ARe5H3hPXwkiWRCzq52kOe6xwUK/atXKkwuZfvd8JNr2qURAaxyU9DczLgWlxEaP
ugZ04X8bwC5mWIPnJFgd/Tl1zJDMUgeMYgiIquD1O1S7zmKUHUh2Bcts+RKO5oC/
tmskjm9RhVzhT+v3X9/WasnOxy71zDBPNUYcgmn+98BussSYWIQF1wyB8/Sm3sAE
o5TFdhjdOw4LKPK85dUXITS+39TCDhiOM9I57lAdxRw6qngJOSZuo2NtMcKIvL9K
/tku58u0X0M2b/BbHvbiImtj9fHl2FClhTU0GUekG5kP+JRvgkTn/xhjWUSkGvJE
pU1RyGp49JbryeA3Qk2whbgKVbwclrV/JPGpagenMhytbUAQegcfKpPyr0BrCBBV
SLS/iOs/yS5IaZ5y2bOsHSGUeQDez+RrQaUwUHMDjSwr5ZIA5yQnaL8P3ehKZqBf
ZGFr8YAhnQAJJqXMDni0W0O9WrXW7K+YcQx8U0iellYmpsXQ2QfwN/PXk7LjwZj1
EG7uwvUJyysVJ8r8HPWgrd8k5eYqOBm2EP46izti1P9EAKYChcn8TcHBqlURpOFW
6YTn+k7lCOZaTxvrV3iztl1QK3S5BxP3ypC07b0vwf7ir/7lG9YCQg1au/CIL6oj
JSzsT2QN3T4s5Jw80/gl8ex3v5y8Ytv7pBWj3jGSTo+stkNmb5pOU30s561Luv5u
db/9MJofxUdEkLvxyPtJbSF6WQW0knDFj/r5qBupBbRQ5DWu1haoluUGCkxMTOUP
JEleFl9fM677+hDIRYR3KjFezeKQw4xA+Q4M1yjHQSbcVzKioMpj/G2QWP7OrUpu
bCDIPG7p0j4Gmp6Q6pMcXQTJKbpcItvswOGYmP99nnFA4jtITushoqraUqbZEhCM
PONzWJAKuHOfq14NPBQQN6m6A8t4w/lnQNTpCVU35KSRZG8cqzAzx+lYIQtun27g
Q4mApPY/egQJH3xVZKVZd01SXjVO25UZ+STaxiJQtFSz2hv/XMmIlhdO6a8Qr75O
YC9eveJ2D6BsIRU/ts+OYDo/7Rfrwkdu3QVxFu/UYm5yHkCVkR27rcC4TQJ5bC1G
nCbM3m/B4B93mWuZUd660KWJklQcJQbVMKfBR8gKYYGlwVrYXrwdtTCCjcGFmkrk
rj12XbJexvj5z4GU3jzskkXJP4TzFyheDNyhEF87UlcmSeaQPOnVYqzesquQqTx9
nvt5EaDNbHlH+F76y+GXmUV+dcF7QO3X0REdys1DS7dotwNxLqABQhROy0ysfi97
XKQzmAp2Dd+8tEtbZtVIKhHCgM3QrQduPBp9rASvkGguVucIZK+oiue027MLB36T
+RD80oGbfqIujnSjnCUf+3gXxstHwVV/gPtgFhTO7vPMnh2Nb3RZyvfVnhtmgAxR
bqKtgCBTtowKZTNgDFTcPXvqk/0EpshHLjGJOsIRZyJRUB63doZjX2wMlB+Rcffq
JYgImh263TXH4dd3oVWNbImmcnpMlCgS+lBSy+g9NkYiD1fvNCSbX/FoxgPjCwBX
QofvNackyMYls4WGYfw5Sqg2my+jHya/GZC2mFFBRk1VW32WzWKWkDNxKxrzBSP+
I4dT3u1nvfLRadhr92FXdYO4Eo3B7koTYHq5hfq5UL9hrmpTDgK6a13N09S+EUrk
xu6HhYTmsv02hcQ0l/gvijY18GcAG9J1UH2VCZcTSeeXXdwQ4IGEkDeGB/74KjG7
onaRiye3f3SKqbTwbpds8WvoVJI78k99KJtEdUi9+SvjJhG/jf/zHjZxl0HxWCWg
0uUQhtzeKZnYKYT29BJ3EJmE4627d1qlP1TrCiYStAiiaau3S17Li8sPEUImSx7n
TP043cYa7Pa7qweRjOaGJEB0f+eK3pU26sfhR192aiE9PCWqe+HAhs0U+CGd5NAI
qHNysRo9jf1a4fz2fltlEYO2ls2d4MwzsNu28gf/bCuXSHEG4t5IdGVXBfOTW1I1
vkSaZSE3Psybjj6mNp0ejBJB8nbVJBtCKQu/9ZIZ2ryozotXXRYb8RLPafjMAPI2
ZYN2V//bZe5f3N5cAxcSZGhmun7gu0M3McG36Zki8FiamH5iGxV+z7WLrsaOWJR4
7vbuR2ICOQ3W8CcWOtnMBtlGTuf8D4BFeHlPfoJH6/wZBpFpT0+N0g0od6zB7SrX
K9JojJXvY3tMw3/HDZ+XEiKnAHOUuxV85kgtd9AdR5laOtpzKP0zT75E7bAiYzQq
DDLFWw80j1ayZAqspqmKvhxdGisFr8b9P9cp5LDQa+Au95IHsQM8TSFnVUugKtxY
/Ap6ujZULaiDenmemF4NOKoJ2fz4nlmqa2wNXqJWBikYoFwGNfY7+jUrJ6zZG/XY
ZS/SEsenTnWFqngXmNlz5q0LPEF65YkOefqqgisnR22k7GocLQCh7bWqwIkUhmmv
fd5pgk3qxgLLOYWteYB830XAAZohOsUJuW0vBKxkIeaGiEKU/bdVbGqIYinnH42t
RM7IuJHineU3TYoMD+cxCnCvfhmZN2bsWsG6cZZP8MQ137pmKyd72FVtq+OaoWaa
pPOVPjAdEJ+2rJQnu9QmrN+KyhUm/CoS0cK236s7LTdmMSmkfmTTFyWNIRCanJ5B
qMLJ4f+MB04tVuN0jXgpjNAvStBaFxTuGcpkuEuU3BHdxGerbVj7ZddUf3kXjEyl
QMu1mVbonUAl1jSmy2mOszaR5nnblrVwN9olLXIrdDJ/GrOZq/6fSMDZLYaSLUod
eeDvXgdSGHNq43CJYaHONQJyF3QyHEDSuyFOaKpWlSd+sb7YPrVz726T7223Ov4a
nc9hiX6kn0SxbN2B1xHIKcx0aPSWHbf9N2ja7dKsU48vNPaOS8OHViOK4dZ4/kLR
ZcszG9jyjwx3+ZTQvV7YGN6cRQvwV+YyWIPoTxylk37zxLMrtr4sBqd1ePhvg57p
gEtSlVQSrDQRfL23GvwmQUCgF/3xvwB15q/K0WhHweAghiN7ZK1+7mO+kcA7lnx3
8m5TT70vEUUoEh+6v01SM24SdMKBuH5SsGPamBe+vp5o+9xuKvxIhhsQIhLyORY/
jpgSQH4qT39XqOO/QakNVojs60ZPABldI2oiMIABHb9HC0N097FJDKYy8hYKCGMv
4TY8Yj63Q3U4v3DHIkTFUt4svx6LlHMKm/kGh5nqS/Lk01JKUjBlAmQYpj1ibPxo
cFFmve3puamD+o90c+K/XLWTSRNNl3mCWw9HmxU9zGo2qNfn7s9N22pqPCY1BvZC
UQOvLlQkrql/YYOgO7LbfxyeN4AVPdxDfT6kj8wPBPWvXd4xBWxa+w1Pambj0Blw
XUW85CUOJs5eov23K74h83NTWd+/U+Odl6H3LF+XkDx3eJQ31BNJPNau9HDr9uHH
E67cudJVaRnuLPTuCTJwdu97m16TDzrXWproq+a/IdtxX3doRUwT1s3kEtV7BzBb
C7A5k78KNrWwA7QpQtnyMBXLhlTTtXGrFZxC8s4cAPo9j+qH1y/WwLBkyul+PC1n
KODbLm6rLYQgt2N54hY4H13eGN3sLm0ZV4tUBbwW5f2GSD8iAADRaD6G8mdUCYHM
uUY9fdbi3zneTrk8jL3Nbciw2GsykqPPWqOZ0+BCaL5TN/YQmW9YE/WBdCBz9AIL
QPwE7JUEs4aikHUFNAbEYqJFSjjcIC0zVRZqlSlquPcxeu1goVhRmciu0n03NqFD
V4WvAIvNqjuQLAuP8LxI66mMAxj3Ina5P4ONhRkiZGQbDVF96/vYk41OxgDog/T8
1UqWGnbSErX+qHgWwPe9Sqb10cGurJ8tsT2WUD7a5dplPBUy45774un0st7qz6UK
IHZfgogHdnLWwj21DuI12RKN059MWtz1Fbj2bP23bY7QTC36UsPmVaeO+AymZ1PM
xZQ4scBKqr2ZbZdOOUX0l4tPFUv0BcWJvpyPgieWfaeK7brA9MV5xv+AF1meanPF
FGFnlY12V95BRZF1GoGMIw8+65kUd60nTgRZMeksqR9o1/xW6YqPED1CKh04VWzF
NHqxRQFGu2NEEQosPXgO04Kow929nC5qrJiAN97HbB6xyb4iAjH2vj0Bqz6pelH/
ObXdPquMxBl+1dL+UxmC6mPhOTqhnIXc9io6xFc8v9sqg6rw3RoEq3b3I/1Ai9Ga
U72qYGbbKs3UhsGDSCKPS/SwgJYRJBUGd/wESNaAUkJfqr1VHGDflYkEiJ+aQ5OP
EZv9rFWLmeF1MFpghwhFnE/MKpfAxGyjwjEM2RtVR232g6XL8FO4TwDstN+L+ihG
Bm2BNKgEnuYrSG+emvoJm+YCYNR/1yaMKsj283kDj/HgJ6JRA26P68+exjYMnzTN
mOrwHVFiztXZnGhsrcCctNO6IIsKTyodSZIKsng6ttA94yyQn0dSd/6l++kcj/Kk
joJu9I4qA+Y02wH4MjVUlnuXV+1m0dprOmh6L8APU0FMMbuJwVE3ZvHlAF0yNQ2Z
FXaZug8vToHwb5cZf8fHsMZNys4GOGiBnvkHMOYgu0U9zmlhQDGKb+L6pJYz99yZ
H7+GKhxYjp0Wif3HKmQSApLimE7D5aaNabcIokfXQSHqFhV2szDAfbUcfqo0At+/
jIi4SSAlp6t9Cn1LElkbR7k+DToqDMvPjZfrpiVqzqYrquh5DvmtNnFXDfbvkJYJ
DlScQVHE3TKlnMZNG7WSw+StVO6fSEDFdjx2aVwIGi7fOQj5cgU1WsofL2iKBCea
1TVtVFWYrv0CRzZ1Hye7KQpbAmPB7iUjTvsmdwITXaPn54gstjrsR8xX8o/YsQr7
j1DN3Q/EpyQcmibieRcXjgWLLECFJ8mnvt//XZJyusBwFI0Vwo2P7hq0fY0EzrMZ
OPV8dWJ6lGDh4fhwInEskVnDnaABIzmTgB4OvlgxjZi1QN9iEKFKleSM78OPSQ8v
123/QljH4GvO4rzZ70dL8Y8yfOC9oviCtrcrVNRDdE2hxv0iP9suQ5vqF47lpG62
xjCiWLczUEE/Zf9xgh+gl4nAriIWyKumR7eOylly9IzgPZzHgd0bJlyVF/7/7EAo
eXnEveWGsDX8Ko/Br/3ILAp2AdVWO7dvnAZNRberbjXnXs0Eah9LPlOarmSEGcQO
OYqgvuolUF3DBYpDa6EWGDNyiMMYcMfD+5nVymBcUpiKPxRlp81BblKPHIKgqIo5
VRWi+iURGAc2VtKNNNpj3/8MX468E2lG6ISegfR62J2E6DQ3s/XVZuHV8ZXxmebo
qVkrYnwGiX48PyhIVF7E6hifnQyusW8nuaeJdAm4azkTko0ShiWcDwDoMrJlf75v
fwncQSc0KK76O6fcxuP9gU+ehhItSYgEsuCS7G5by6bkkyU1qMlg/ON68Qr+pZAz
JOsfofRMIa5ZhQDcAz/o/aGLPQ/6VmoMSgH3HCLrF18+30U1IfOOQn1xa6Domu2D
deEBw5WQ5dQMi3g5jLoFd1VUzsqA+mTnLYCJXAfG4l/vTJyFGAAV1i09PHzMWQEQ
OQzuspoM+a7AdvoEssawH9qcMJLgUriTtHMOf94cExkrcj9ai559R3FX9IgM0E0s
ZxLc/ltaO9CPsJJ9mnoes4JMLicHIHFLoEBQZM1ZmxqXMkjnhxbGjAaT/uZpKzxi
vb020clFVqlRSrYYz1yWxHF2fqJIam5HWUkEIeL4n3MVswMY/Sz4Fbbl3reKfCwW
UemYNYwqcv66Hn4OXE5HlgGTG61/b8bQ3H8LG9GDOMx5x8JAK8lAMx3duiALWVQV
pwHb32H29HLpzaWY+unjSmEBg5CwiOHL7zbm2jRXW6nk+q2gugAqFAazcj34KjmK
Bj0oHCybRdlpPdEAPVR9DcwT1dfwBfPu5/ow7WHnuQvk5tchI4qOEip+uLmxYdRa
7PWpl9z7E7dTAHyPSlr/EM39OG4bIJmQ7qtk1cLY/7lNU4gn7nmMFy2Tzj7d0W9j
SMJpGiD3O2XCjcMPTkrggVm50OY5LjU2DSeuztHa/lXDuQ3B/ZG6d+4JIyjgwnoF
Cl7zJpUxe+0sbEnkq1fVt+oW7N+UZGlP88BVPjUQt1E8xMGpeGVJIVKG1rFa8aYe
mvNxf739aUdHQtkJ2X7WNLGr8hvlOg+M5fccbYDyHyRTRm7JWYrKuAByyK+zCBU8
GYjFwmA0UyHB+fgBpEjQ/7k/PKQ9QdBvT2QWs7/LNlugxc2TCl32KluOW23DdMpv
RqxeP7a9zs1T2rZlTm5716r5n3d8mcCAqq4IZ+ySsIu+GtwWDUzDn/WbCWpSjitf
p8/E5YI4B27wBN9fGhb6XeCErfPZglfie0IriE/XvUm8Fr24/SloBFuJhDOvggAI
QTUu4mB5Uzpx6JuXUHTEgVxiCUZYFNwTWlLoQgPv3hrl3dRDhS/xuHLfVC2ax9PB
6P46j7ppQ9g/k++lfZazKSyfiqgIvyMkk2A0xy8/4++Nc8LAGEXBbmaCf/LKeg+3
OCw912XijGLFymL24pmy/NR7M+3av/tk5GQbJzw16i7R7K8z1aCt+e+lBllYRBrH
P5nh3d6SXFsZfNA/uq3LZ0Ch9LBKM3f4Rq2OsuddnBjlb9AJvWa7Av1Up//q83P5
FsOImbpfMBsSvdbLQ7puke9jsWXrzqOUznSumnjFTEBpv4WZBgyIhNkavX62sz+Y
opfVjS+U5/LeAILQwFwukk8wio01of2E8aRSoJRAv9M4uBDU60oXtAkHmVPPeiuK
DBo4yhKxT94Cd2sI7hUwhgOIVYkzSZUQZLjKzA19ZAWfhJQ42HncSIfg6HavFOIB
aPdG03Ca9FL9TEYP9HIqBH1adCU2f9S9O5+nvzt/wjTuyr/k65RrF8kXMdArFDTz
nmM99aPQ6uTf8MHrUeWucaQ3fbMLqTWcc+HXzRBJTXve2A0PF570GzAMcjn57Z/u
q1on9IwKkEij0tpUBYZn3zuyvGRsQxyJDRp65FCqbtiFJLxl2N9LX1Uur8hRYplE
XBg1Wq8CLK1Ed8Hd35aZOXjMUvi3gzvG5HyAteSILDDtZWcKblu6omeZHa/Ox94m
vL8LSYVzFxT2smhdEthnHpVt1YBIhGx/YX38yKWbNDWD6aZHbSBGuBYxDXhBA+mk
ZqdRPzeLMTNZQvKT+yqKyDzcajTxuetOkhzBX0terVNSAwmvriFZIjs4s+2Fk+Tm
DEH+g27O3lz0NhcWIoaF2d4ZIBw58LpLmuhsLsz9NrPl5tSgAEMNPBkb1X9XmCkb
C6T11UDC2y670MZnXPfssOk9u7uIqMHTcQLfb6NShZcUkE7t81ttPVHFxRgKGEn1
9CGog1v3duoPTw/2DyRK9rAlJKGizdG5brQLQqUszE5i4VrdYmPIps52JSEM57+g
osKvaEXXHsjlutkj/WZaJ6d4PAmw1mwQAWZ4SnZG6IsXeQr39TPZncYDgylnVTYo
m192Rb9SpQPKXmbvCDs9dlthWPHc3A+jKjWwIaoqADCLp30j1CUL78lQqs7ASeW3
qd5Gr0UT1xdXeOYQMQnzHrtFRKvxa6WSAuaTcQjgCfcTBusDVBfaOBiHiWfRg7Lj
cyQM0TUeNegL6cbi8HNgdd+9/2iqkjRLSFKCZ1UJ3qnzDCKQTftbTbg+oKvGGU7I
OEkF1B9cVH/Yr/1vJZBWkUrjn2oxQSy7Nf09RzttNwpI/nsVlgMa/R8dVG1OBaB4
6tuLZaxQpwy5LNt4ERqrOW92KBVQ5wBgO6Hqa9vKUm2+4tAMKuMGzzKAjgkmx1/I
XWJMg9eLrLrv1uOWJls+OQX66IoaruAwEcmVqtcBX9xSBvpmd9CVciD41w6LK79S
hlm+uoatvvikOSNdABklbpr/hZ0WL93emrVGYurS/ZLPOUzjYbutoUDDlo4V7HQb
2LgXea7xZ277jf87wqpahR4ql95or0V/W3Kp0/Fs77HepTA7f8wkxxa1GurMy0tT
0c/OqoDBJelq7gt4um3J8Cp3Vo6m0r9oF5mUNx90iMfJp4Qd2ANKi4J50+ztGuJC
Cuv+uje6wgfbzLuB51S3nJH0gpMUanH7rFO9wjpVR8cRkkvrrJ+5ABHm1lY3liPD
tDOuhVjVtDIyV9aYJUD94vV+zKe9Wtd/9e4Mc809VqCA0CWJle6W85q2Y22a5hNQ
0upyhKrkKRqBEofShuU0aeyKHALSeNfaJwjzFTH7AkCBxLn9aKy9ywwSithfkPGs
SnWsUvZbr+JEpJdZY98hYhTDcCX4Io1qAzkxuYlvRjklWRP67SDpwPbiIJ02Zqte
/QmH7tbGs6MK70xBK2mMuNPB0vpgn2PITEhcCDMohIxcC6BrFjoGwRd2SY8lEUF0
HGgVqs5ei9INcTR7am7J+awt690Fh1lnMqAk34Cs8oIRNGzBzZxCLjzE/XBWDR+I
MCs/+IJNONzp8PKUAAVOOhH1+akl59ieiomvLPbUbL3NXlX/LUa/h0qk56+w8S1J
xHVwCkvjk9usY7L97giMOvYqAfKN/OHIQL3bMoXvsF6swIGvKfEHNhdnDGq6hOCv
mhfC4OhBAK1iXXXXvH6U5MC+c1ygBJfsDhpUe6w26gIvHtP1iWiqkW/hyChMsaVc
W/lf4uET1FEmBkKo/3nAfeWAV+ERzichG4Y8QMa/3BmWk0bDvM52pruNmtd/V7Jb
1Aq7nC0jmDJ04xghHvKlBNvmg4prR4IAxVM8ZKHrCPwyg4oWIqHrWDRDJJ9nCU9U
1FdiVHQCgRDTvCO0xEq73TjnStt9ZIwewX8par5AVrIL2qM8cTXqduWWuEDXQCjc
c/jRYpz3XZSgrQ62UnUSNwdkWA6cM+fFBSMelQYXUzi7faBwOzGuqxGz0KBBfKhw
h8dlkxyj6PUkRF3igd4XqYsX6kAQbqSZEk5lHFmfXQcw5K74Az1dmyYy7vEjgww0
Cu1xeFys9iJt1wXDNw+LwhcYgediY/JcFVvH2W9p+mg0R5kn/tJd5aaVp87pp99h
OgeZXhh8XhI1KIjmjTlMOIygOh74fOFqpnhCgqGE83an8jorImkEQSdxzTRhOqf9
SArhfT37deRnY9XqYOMVgDoTEvmWsEqBkvrlF3BL8jO3rPRZziP7pcgirA6uXLKL
pzfiIMhik4bJuScVpsu4Pvmtj+e2lyWjzz9PEho4z06AbTAMgbifOlEjNT9aCuvF
1+zEss8kbCzpv9AiT/Fz2X8bG8WBZEWn/hNN/RAGWg/b1uF4s0JjwxCGmus5hArv
+3HR8H9wAvBPaLbMco4BtaoEwqsPBY3lMWrux0jhytvhp19woN/KiDX9NRXf+rJP
5arxKQaWUewmLXOTK5CuXt4NHt96YQgwg6MJzZMHXdDNkt/hKU5E+OOLRvdoA/eh
HYe60B0PtZouXAIwnNACBFeJupJzDZKxE37H4VqnbcBErjt07gmZw+oB0pGLYYfH
sMDL8faE/XjuFKJh49LOtOUx0dnTwHABYTDqvdapv8fnq5ET9NwoOZa3Cam84hY3
XDd7yvVzCL2G1HPzVMC6OJa5odw0ddihMs7oxwMgbpMPNWealWncSc1YTNbEplcU
302WPXgT+8+lLg91pBw3CEZy7ui/SWs1TnLaI2oUWIvRCkA1m6hKxp9RQ0tytZDI
Gc0Pt3Ke1pRJe9Mh3ztVygL16NfKf5ClgsbTb5hy+Bwtwy4LNH/q5rP4UA7hiO0n
irbjF2o0V8r5KqQf9pZBBABgeG499c9Y2DuTPdEN48cMmJTWtWgcbo9c2FMqQ7jB
kkzGuzEq9ZmeGlc+JHEoS2JVo0bddWTlQuCp69ocai50wB7s0QlUm7byEqm4pAUi
Y8tm6HMYdelZgVpRffZNne0D/IW6TNxdwaZeu/l3NvJCBPJ3bfBVhXs+4X/AF/uB
TGNERkedDLwcuOroSH6idPXH4OP7l1ct93MWhHJz/P2czRoj9b04hHv+jnbeb+9p
z9BYZfj85ZNX6OHg1h09fK3aFdasxefvi6zMsrVCaimR8VwRFSmcFqSkSvi/xmoD
2YChWg20Hcm+zrZapwU4v0SUF1Ebms/dVamwqTNhlmDmb+JyegjaQOJHhZlsYboE
tkHQkA9eB0swMTLW29jt3X64VJQ7LIbwuZjLSQE/8atrwY6aEhwbhYoBnAN0Pd06
o2hSsY7105CPxnvGNW4GJF+vSzRJ+rbqwEelKEJn6CWAsF9pUY12zkfeu4TW7AZ2
ycOEabNGAyB5yysuwDV81Aso7+zwVH7OE+YLtnVDHEaldhr+8n2H7wzgIpye7AWT
YI+ovnDokeTN79hjjxrjNKuJ35tjNTQzmsI/xemclYGIU/6X4zBB6br0O0bXaQcy
nYZnTG5fMqrhEwPlB6oO4k0X93S0oNd4MgJsaKoWSE5yO120PIVRuXuHNv3X3hZS
aZg8pqleURnD2bSXi5jTmDM+7viO8tPdCNm4OZfCXuRQPliQWOfoGEP14e54R5mn
UAA+rkWr3/HYgkvolGqLrAdcMtId8bzUa9zjjM0xifcMu8qrYI+lFs+XF/PcZ0C7
aDfV1dQ7ahgBsaTckrDgzrPjmxyTBP4KOFH3gh2bCyHN5LQdtcfrz8+IPJOAzQuN
bEOp2KBaFLMaZdwqQU94lZusLFsvhMmg5tsxK15EaFv2HIlwyxwPBtqBjniBVhGn
ralaa/MtoLbnC8dar720dZ0fgraS0ExwrNaee1g2b/1MWxJnCS+8rUwGYBlfuodH
umnnabLrTzE/90Tbq3PYiyaQAlLOEJOwsDAozSYtaMQxwYi286iQzr7ZPuXonhDH
fwR6uR0Fty4AmEIlBQMMxdknzlNZY/zAh/EilhxtFmzQCcaCks3rOPYHvgMDC6T2
1nNLCqzuUEDZOAAequ3GIGPHK7054nKJL6UJUhECtkaHKr4APmBHpOJr+DMUt+8m
U9RZSwWO2PuV6FAaIuLfr13GIjrmSOzzI1SGWhjpXWbfzeBOEqgdNMS1Krr548Ly
AjW3SKuBlYcE62SXg2tUwcONUldmeDfIW9gQ9rrmGzowz/YoJRZoyqGP1VwDzHEF
hY6Or92V/wCawYklRxPZQkAPYrclX+K4JO9O5Jp3OQ3PX7ad8chYibwFu58cNYRd
aDgzddz3Uv/lPT4TJD9qEZbaABO6ylD/cvH1ccV7k9lA3mlmbz+wHB5gQQ3oiZRW
bipCkvT8OAUWDdho5IwoNF3ZZ++lPAK4BrUi0eNd46EjfWt+3iqCfxvBL3PtQhzU
SZUV4Bw9Dde+fRREcDSB6F0SPkp6Q1g/q79rX2vU6EbrWV1l6+j0KmonmjJnxVCT
osg7Hcz0RKJwXzDgJpGazAxyPEJh0t4zPD2/G/SsDETMyMJmrceC04TITO2MCsbb
+aw77+CLeJkSPECF/LjXNd5l+0DyRQX+PPyVn/LpOEa12QY12wl4JKxgxMLEDJvS
YKUi0F3c/qYhxje5tb1YMqO2souiDxRgX4boLqLkHUfhx9z9cWMSl6XTWwGC33mC
BaAK7ht2eY82PrzxnXSZfpIAmXgMo9zgNEojMHujAKMl+5uUO3Q+6Cbzt79q9Eyp
fOrah6j2I0JCoUF8fUSxji/ZtETM1RwRA+Nj71NfKH06VVNkeXwiAyaArNsusoQb
XioK/hvGwlQjT4CP69BNfZIxO5UOVmiBeM5+bj5INtX0lX6rg7ih14s+Qd/vv31A
WgS8gtxWUgXg+eC2ZtVRWxCjgxJcfU8rfV6TM4wjQgnNhGotFh4MegnMoaj8bUWF
kBVO4zqjdJhXBjkzO3rpdysAB0iVfxby+48dSOEIVAIepbYeC6Wfx3kgWjIgTLF8
LemjV+LdROZicyrMfzEjMdWfmPYjzITALKjmKP4upfYmKJk4VfggWp5dcWhAOYHd
0bdPFAebvzBWidzRWUtCNSr2AqMiaLIUDKjmJS49zc+OTUI5OWPnp9l5Llaw7OcT
sk1Y1SrBDK4KSuPIp6nLOx0ANKpDQhMhWROq4xgXt509uksU4bDkmzK0XznSve7z
lLSEOVFYRVZ6wOgoi/XvgGV2Ip0Rnym7ab5mxvL5yItZ658zN3EVYUYP13LYITRq
Kib6GxCvY7NGM7nZ+Vidh2yb3cq1C6+MjIpQ2w0NuJLzKv+V3HJAc+SFyLJ4MH9K
tagcPj5KmwyX9gzMcTOCOGamMsWu3wGr+07uTj8HpgVJ/pkt1mkiwOPeCxpvGG8n
nR9tJJu9TsqWhoTVfLKb310oMCvknC4ywUPWw26FeiZ92tYbxiEnhyxljxymRwhV
5Zzk0STUhCfmgOXEfChAn2/sX3mK1GEhM4I9VIFycf2AUhjJA6EGQvhbPwdpXxjt
fbocZi5ZhqJHdaVXj0ESZ56s1sS1BBlMASVCcAzUCOF9hFkVlfPIvaWMLShYVyQ6
n5uo2WbeK8HoLDivWN+XOtKrgDizLwJY9YrGA19WFyRfjBxSEwW/pLy5xqv2wVRI
SzC4ZISZurd/wREoxy7B9zDA46YidHwiT7PFN4fz3N8K6j6iP0/yjpKvWLd715N5
pbYKrGiQ0Bp7AYzT64fUhw685NlORsCOv1I6qnbE0lrALwBOwiWYpmeWsLaIpRNu
zAbsqzUA/RxY9j+rqWsdQdafCH0rryDSZpnlnYHlb84Uy7crNgYYnP9ZTpETXjR6
zqZ8fhPwb7ME1KzVrumY/BjqmqpfmoGBiKjalOBLrQWfqQ+UnzUWIBqvVTTQMmF8
VBH0Y2g8Phtk0HTVfQvgbNYKUDzfoG3az3cZaOT1xKXc3LR9BzSNQSjG6pnYLSIB
cMTGe9ei4NIc19urY44BD4gSzbEB12h7Q4GpJsU2zBCeWof9TuOz1rE5dwYcb8zP
OEjoPK11res37eA7W3ee3WQU5kAE1Ku6VemFYK0CdxLFpMCt+8aFQwKoIZxmXW90
tGlK5we2AyDPapB1DIDXFdo+gEAN0YMH+aFfl8LaHbsoR5BWYReF6yOyP8xC7E/S
PLERWAskia/3dpwdKPMowJzVG4Ur6YJvHN0FO0VsPU95eyRvZ8lYM6KBft3CqT7g
YWlE8vvmDpUNEDNAYoojRXaF7eCLa9oGvoaoFa6JGaCx+Ym3ICQaGyc4+wiNBs9Z
gPyJgXHA37O8I4I+ggI+n9TQJxk7wsxRM2SZYe5oDh7YKwTl6eJ57HMWsyp/jlWc
YKmbAtRC8ig2ZdiWgfZDQNFdXJs5pPrzHrmbSH/j9KJKLUgVy1uWSvErdY6rdsIS
Y6b9tuYEnxtdUAL8FDuM2Q/RKIHiIrwn42bZ54iOpWgZbPNrRMgA41ll61SFP2Zh
B3YOp4UKZlR04oMmwHYgUcaxAokjTNgdirtnOfpz15TB5z4Ceywf4QdqOH9phbub
XV83yP5liRJNx3yJdsUFzakNcAY+S6RusxKbB5+oJh9Bi/S/tI02H/B094EV6/DQ
3KutsvfMuRkQWtTTwKJtqcgczQ1zm3kF+ZHqWlRuCssa87ttHMmAnAvxFbMpYgX5
fJC02jfbSwxeswZKiaiQu1VEwrWbtfs3vJ9cgpQWtsT1eyoGRueryUS8gD58fv/r
OC9Zim0ICScBoQ5lWbVmwvg2rwN7bS3jT0Efeu52j+g3sxm08a9uyaEq9UioPXyn
4C/w6WKIM36JgPAV0fKmYXAxrBZMFV+4ifeDes/kAmcbRBXbkgmLU/iXYSQLhZgO
9DeeC12mHDu7GGggXCIB0aRn+7fG5qStsf60Hcjh6H5Lr2P2iX0b3t6vUg7fVtV6
s19keLusD+uo0Eci7s92JlWJL59DXbXXbgLzjZZaOygAEdOf/VfZfm1On4DSX3Pe
wP0dGQ8aLz6m/v2bitoqacQIJlitgMFZuk0SQhqQIwl35Dto90HxVGDfGigUMuoR
9S/HvzCeOceT3LmYkpAZAytyx0is2RgnzRrFT1G9316MDNaR/uZCdHqo+rs0Dcpj
uaUAelq+mhPjCU7CU/pWavGmbPZ7zRahUyUI3BuyaGwQeLfsVtlV/+edeKARy7fp
PlhSQlT6jdgm2jMlTNq2XOYNl846qfgwsZBrfSYKW2BBdyYN+6xffTAzYcPmM8iq
mh0Yb67sK8ogf9OP52fmRvYwPL3gBqh43+9x140OkaUD1GFiLEI37i95A8MsCs1a
vWtQr/Qq+ZfKmix1W7ve6jnwxi9RoxTrMt5SRl0cjAQpKsN0As8byS+NrdDqUgSH
iElZf8ByKzLW4a238yH+daVUTVKJZT40nAJDwxc9FKTxPx3B63eOO+MLvo1T9d3o
HVsNLqcMy3Q3t+KP+j9UDEid6plFkN7tNJ8ozfxUIhjW14Pu9vG3+hQyVKqEfT/D
cB0P34kJO1sfp0kHb5+bngaTNc7T2U3zCWM4BQkKnmYONguC6fyd4TttcvUEW6FE
L1PBgmWjUoNYaNbOCxjO/cOKGlbwuwjZ9eNunuLfxTuEZ4fmIZxusaisAly4df4c
ZjEhf72IfeTXece4MnU8YSACkHrOrGYuyXoo8PCSG8N/zWp69tIPcRxHVfxHpoTy
Av/rg7cQAn2DmrNmCSF7vNy23gifo7YE2yZo0ERmCmLnLH30Rhh0WW4/2r05GyfJ
EseNwCWZLlGsYaPIdClfZo74IO0ju6lkXX54qgq5uOnvU+TBJQYiXW24iy9VjtDm
r1ynikzC5xkXdHKv62RprOuhUMpB8UeG53EVM4ho4mK/hTp/iFMNZYEmfSUT9gP6
JipMugJRdwcQsYXlAUPOZBKIQQBr4bUQ+h/6Y4cUqTW72MNXhtxzflzgm7EZ3WUm
IjhDRGFE0Zo3Td7iDDP+FwVw+85ecgdh3NXnm8JUvn8L/xV/miDW+J9nlco0Cc/j
YuYWXrSCihpVrxPe1/jLWVY8c6alXlyjDcY62+39ltFVu6c2j4Hp8CaRxRMaB0Tp
PPQ8tdSwi/Z+8iSItsqsX54uWzcmEcXworD2IRCVso8Srzf7UcEzcMzDo4tiPc48
/E4rOkeihFHK0A6vaxEmpOVsdXPy2O4+fcGeq+fBwf/hkx4biOL40Wvn55x1uE4X
RNYBqs/Sp2+MosMWyX1gskkz9f0lLn3Ylt+ODEzlpjt5p7HUiKaA09i9IinU1Qg9
Mteh2G2BkfBooRCViA74sI9VOXnKIAb1fSUppwl8rojekW/xaEtAzZL/AKewBlO9
G/9yFFzZUk+sUNT/hAoaZ5vHB5uXbRjpyzNC7T5qSg/L0vjfwvqI78IGA8mACKiF
jf1Xl9H1US+MKCBMXpG3QhmDyufjzseOpt39C7c2WfPwIJaazKEWDtl997hADUAH
pzOIxUWkH0r/10ES1YSmBxWTxkG4g2rH082hcnTPD4rVX617NV35Ega/Ikg5gtE0
GqTh66bM5j44pFwMqYj6X7Dr0nXqOjBfKfEUJDQtH3T7NlRvRhP6KiVKr7u0VL7o
wthYERCocN2F6CH3DAPfQcyOHl1ykYng2XbfjI3MyqNqDi31U2hCE3pHiuW9Iplz
ycUoQ4pvisQX5a+dQKam42j8aYqPu81G9Q55G0iWdnKmWU5tnBKwp70F3K9YH0KU
z5IG0Qbwua+uKArppS3lPTcDjiI1EjaOvRuUEzQoVGbjRf31oljLGYMyj1HTdP5z
kmCi22wJxOxr1wSiI3EKqKIAPxbYHwu558G5G7qARvNJtLEikIj0LwNDHADk2+sP
6y4tIqg9rg1ZKf/ZkRjyDRyXMgP82TZHDrO28lE+dLiFAlQD5KPqVfZaNf7biHWF
fHyZvX4bDvZoeqoQCEAzY7ljFnGQgMCn1CEG4S6DV+coZLlD8CIkryiOznpauC6P
Bb7mqwYws2msEA00FPK9L9ybjdwRugrwDpahsL1zvhXCseOk2CDiR3ErNbqs3XD+
w1EsJL/KfjoNWvA9X6CD45wfcINXrUG4veRIHj53msekowV/JqoJ1kax+xmJruui
4g5th9tlKRYePDBI5iumg6N3T67In/rrf4qYPs92DmUx26EVPJlrPRp2+AWKQ0lZ
v5yKxzkvkCbxZ1bf8BAHOwOOQtHRA2ut/w6li4hj7j0ex51yEWmM19P5GGUlti72
SOwrXIzOFo7FFw3mgMGJm2SVi6GsGoRFgP1RxCGcs1pk0/IfOqO7WMOYtROWAT7f
aSfqHM+M4K7ctsqMsD5TZp5GBXf62pNn7Gs8P0CjBdED0hetv357KJiVQpI5Jicr
SYkOJWF8D94tTzzz3SZzPoLSJHRWZLGGL5L5J4GAbs3cQx5w4gMkBmzT9fADT89u
3acRfB5zVW7msd1B7H7JAAofCao3+fTPOeLHCOT5QHSQmC8hyFnKNgHPSNXdxchU
loGhFtDgx2H+dpUt5QPu+eLeRR1sy1yGUr0QWMvwsSvppXqIvIBQoSXh0rQFFaqe
g2FK9+D6TXfl6RpfBFK0VoL1u4y/Wj+HZh3ORXxTndZeGac5EVlBMsi5o7gN21u/
X/NnJCsyzn3oo8IN+Z9RznHfbn++ey3B3qN9KCxD3p9brOjJmGqn/yJU/HvJRrke
7fLUJjrvgpCNs8gHtLhNqb85MEq0jmZ4JmoHgbaP0UzeN/rdBf0qM3354BKMFdA5
1/q7Ypbij3B/vQFViUkRwcv4mTkeKaEsz0q2AWsAZfDIt/EvLkL+HbiB9HDOQjz6
3hN+1qfffKJrMuLV4om/82pMH8R7v5JjpJDkwG7ugJyZ5809tc+akGIQlEa5Dn7X
gNaka8IUuEVbLNgvc+GtZbf3aAgQ23AmjO2lG5vfRQPHHkMDJh2jpHw7HwkjnjGg
tD2zuBiHGHiEdbUi2YuWRznPMfVYLvIvo5F+84tZ84zALwuWI0umx0i+5VmvTJC2
1+9iuzduzZsHk/38U0K6KeQghPHihIMPDJ4Tx/3r28ixtXk90Dqc8qr87dLvd7qk
0knKcO5fu2WZoEhIkpnNj8FY3gMT/0vtWr2uZc9YZFPaMwB11Tl3gSomk8UBWhwS
OyjaDlMy11v5m5PJ3/yiGqhwk2ST14G0jrFC/FSOHo7vRwFyeae/MbT/rhDyAd7H
fDKHWkbeXWcXIK/H673DyTWneP15mg1eHrnm4pxrriV7NCm3+1jsn95TSD1tVgEY
9b1AUvA+9hqlQGWg4YN7e89qIFjwqYamZfzR8bYdyH9xhw/kql13zdHwKN2Y90Jf
AZSVsRapdjX4DveeLs5rPNCzJfxj5LSYgmUKu+cbRQWEHkgqs/1Lr8LvseuW5Cfu
22wWyxrdH5fdlylhHM+/r/KfiamyTv7NbxrJ71GlniGMotTFDqbrE8RNrupmRWjS
wSt1HnDktSCsbwUhW8BLMDNRvTBGk6eQaDEppFaCn6EdjRtIMXaG4W4qmw3hCt53
A06/ZLakWObocyked7crtLslmsZgFAM4DcE+80edk/rptRXS7DP2igqaVuDo0SOd
UZ1VFKGtZeZR0w6TBxWruNlLb9z0kzqc+/yxmd4iIylRjom115UZXdChQ3bkdk8U
oml2rNMN0O0DI7DAAUBBZ4rYlHjCqZfUIYAT+yMTKMDyoBNTECYfKl7TmQiQ+1ee
ngM527TduJ6qFqufACrPEcDRfIpMP1Hf3dlNUw0u67N+BhQ7BRCa2Q5CYR0HodZS
c0/TqACjgtGLe4OBN44ZvT3cfbL4E2v7VhYfMEzgWWrFsHuDFdjp618lzWRx1HT9
0nRw6njyYk5kEW3kz7mWllqVGTFdUjod7uGIE0A32H6fIJNfQJW43uEBFaeIUOJh
QhKSZHz4VI+Px4xEhuVBvhrqMbw05Q5imm0LykL8a9HgDuVlC573VFnq5PnmrR87
znMoNDIj0Sr4w97TBU769DhzpPD/8hP1acrKZEJvE/G3N38IBYn9w44I/+LZ3Gfo
yexlOKukb/4WxLzUW/H3FgVS+/6fvzoFqqshxyo/zLVNMbnGHjKbjiwCR9JGfw0s
pSy9ZeqYAcm4L3ObsR/O8EbH4kgaEa7Ip31uRObIyWQ1nWFXzZkEc9wi2XuWSc4o
vMIaHo2dlbxSF1nmY9Z9MbLTXYOyUatwcpQ+pD4Y66YKtUHqwY/WDfXx4jBgcz61
E/nsATXl1F5WvzLMFy72XJH2V5+Z/KJ6O2ges29oobA/+6cxhhxG1Z4UDpqNkVEA
uMvEcZcVjqkYq3fgYaTSbazANL+Pz7voWtKmRXGk9csyOhoAi4+rcxA6tB5SUgPA
v26EeeEe0pgL0kgaIindCEBOoJ20JVcUbaG1xORD7NVJIDGeoLu2+lgWGqn6Ws3/
hRsKuZsiBkjrT9hIiuDyB3ztFU+PPneG8mCsODsQ+UXIGLwYzbY7gbvSgkzjUodP
HYt0ksamAXDXba4JVGTBCYDvTICpMsxwgnKOPd+09GDXWIEO2kQ71AeT40pitGk6
AN5NDVCQUgHDp8M/Nj0iIkLaw0bI83ne1RTk0Cb+vn8PhOweeZC0uhFslz7CU+/F
c0/5UGJDkKMVHcUH+9kkE2B+2QSJeU26bF1vIDbtyEexwUBxojdvKTmVfYK5fGQo
R3EO9oX3WusXs4h8iIbMwwcjYga2NjOlspeH/RsNGxlBDdfAMd9IuMyaM4ZXNT4H
rDoKmffIshCxBK6I66jl/cPr+jxNJRQlHaFT3t7omANVFEHTRF5ZoC5jpgNMpZgr
pz1y1/miB2bo/6+gSiDSaFj7kcsLbxQ7Lptoj1wYOTp8UXoFq14sh7ThOha9dyaF
tMyGyWLHrGfqpBx2PBMRXizisdmZKxI5K1Iy4nClcJcCylLpDOyZ/A79KNo4KUxV
U/q/sqX/y/UL+eVBC76d3aU4fMflo0MDC4tnvCQ//DAME+P5PJKwgi88FdQH4Lic
NQvHCFRdsNUXzxKkP0dN74YDy3ImPwAfYDEisX9+BMh62KZOWIxuBR8bFTLb6EtH
mYWpUyBo0loSk2Wf5+ZqSinxV003c3bbTckPAaFnlHuhS2EkQZB5nYiyylhVYHkw
37/kmSnPEjq3syOAocQhkb1HA0vUGJyinrskpwMYe1WlyZYd8fwW74qjZWRJqlou
LKdTdyqHksUNxGpfSZcahqWcOKXrYbgIDnHEyehbVXaaqyOBfnPJ307hgJYgqkYc
MxT+QuVu5sQ0aDuWSXvqPRtWgrCXF/xFk8nJyupIWcvRosxohs6zcOWK7Ja0qzMY
/bOT+eeqTFORDKmbix0DmyIywSmQG55sE9TquT65UDzfQ9yA+BH2q8gevZXjfBj4
q5QiebeoRyVngr/Xru4rjRLBJyonVU8pe0Pmz7ThWejF6PmMXZ3aH2qzCrSotRfx
ly0fNgtkWnImqGLpL/d6SJFHHG4Rk9IrVC4LADARheg5juv2K3D6hCrtkmHYK8+4
irLDFmbRbwq6ZqB2RXFiJ648lLpOaq3OynJ9UfGCWNYSjz6xXaJifrUyW7bVKeje
aouZj9yJzrHwV5RepGZJBN6uL5qifWROHwGYp7ipAaWY1lAcPPtBmgX0IEjEr09I
lrtEIKwLtVjnbExVVfKiiMEXTW3sC4FlqNb08MPiRVC4YhSMMs12Y+gyeOvnOl2r
CZhkIp39XOrf8zLarnAg4ts8xaBxjq7pBVFWEd/AP/mOuhEBWvJQShejPH5idDf0
/Dd27cZ28Rr4G/sfIV2KKcbJR/rYYiDztn3mWu0gg7npff99mHLgafT8sKmmn3oV
wvnJco0glZzScKEU6gfzTNFieEeotSPnih/8Y67+bMJczl8jnPBBNtJlZC8XTT6A
1UZ/JFNQHUTi7972ZqLicJowautLxtv31vwRzb/WQ1RJQQHUx3TAuQ/qIWt7sJUs
99ml9t0XNoaXR0tKAA3fxL3r81CUYG0xXEWJBJgFR6k4PlcAclwS9i+8brGSY4CX
Q5enWq+MMDhaY7NRD5yH28HBtU2I81JtJPsFcRpx8BJUbhNgCVEIkYezKN/wnrcR
cKSxvzdgmJvDEQRNMnAR/mHZALMNnA8S3ed2vpZ9+5PpKc5N3u2+6X6XDYeojSUK
c1GIGXxW1mvUfCXjqsqHxDvDy+Fr//HTbZEfLeuN/TGeFpI2qqFhAIAPcIWBbWk7
jDdEDEUh/uMQAjs5hlNGuRANdJGOx1rxC1av40lQ8hC0/k7CpsuNWf+wzMaCNLiX
D1UZB05Q/h+L1YdfAZpVT7vSpwOu+Ry4rqBMtUjrP0Oh6mJfwQB6R3OxhXO/Qkem
S+5lqJG1LkPIHvvoojWVCtM8OHF8fSpWeB9HVw/eNKtY9G9cU8J5xlKoztRA/MnV
yuQOV6EwPkFaMz4D3Ym61uYfy43fFF2Em54IoaDAW2czpiGdPYWNgHk/CR5Rrw2K
3RRpG9XeFKN+0E/Eqtxlt/0UJA8OI5FTcBc8vUPoX6D+U9SP8hkOTMAMejh5TdiS
C9bH05raUHG5QqhqSV9xgZJgQeVH1hB8FWGYsjCsoU/EWqIDuHW6DW843SI/XvuV
RYO9BIaMog5+jgqZUqEvf1vxNUpndcLu77vZAqj42xCu0KNsVM9AZg3jSD3SWDZw
CLNQE+V20TsBDMl1AXX8/rrnflX+vTXx9FJ7R9kM6r7LmC17TQDz9l/D2xJnzoV4
y0Q7nFcJsWTubYNpcwumQy4ewcsJIMeQq4zQquAxTfoxa/mGQrz2+GFWx4fIga2D
JOfyFB2dzkZI+B+ecv4HkfW8UTjkCjqQ5A6zjePxpZAmzj/ODMaF8V1xddZ3OVRh
HDh9KpHkwodLp3z+TRVBWopc7l4WFuhhxjGWqSGhI9WgdpurgCmZ65IyejsBvDor
rN6vBQm0NLehZ8PCA9Nf3nfpAeZ7PdQUISKnLrqmo7KvCBb9dY0pqDBmVHCe4bq9
h2JNTH7r++4BS8im47UM3eW0NSJVEZXhD7qMkp2mHNNwwChAjKS1jvHLRM2p4yLD
rcbKwN71ySUUlSLY0i91O6FJkMvpNKe95eeZRpt81db59/TdlmPRUbuJab64iCZ+
yaX84q6AAISlzM4LezUcc7813uK1gkYwSba18rg1fb2IW4DssGxb9RXFPa3ZUvZF
PQolJwNddcrpn3mPGKjRLJZ0aJRIVaRInm3DJYvk+9Ycsi01S4s+gxd88L/guXFC
RVfno5HQedTFyuXojaoXNws3Ud5OtC0Ga79XMM8Bg8WHBJvCFZ+4ifmYTPRnaziw
c1pQ5r3pGq1fzuZqj8SkD5JtW3x92WSmmRSYD8wjf6mdR4xWeY8p28UgZbZ3v4tF
DX3/4W8/WsZ5+8XFGnN9AClWgB+Qgo8lPU9uS8J1BhkAeqZKzRrLSXn8vKBRWDhh
F6eJhaXJwj2QQlu+5uRm+PYBsanY8uaQdL375vMK4pl/6MAtysHDMFNVlbENiFaZ
H7wVqUwrHqDfMMQgDFL/aHOnph4p1H7Jt3AOiDMDfRjackyH/b6ru6kfF0ReTGtu
/AxQFHysiqkks5cr6ttX0Zeq/ivLIVuePWYc+25axHx2gvQeHQzAscAQ2sKa56tL
frbbHeP0wcveG/TxV7sfOpNo73jJgkSPdOF47xmCL99k6LYk/lsfMgJuWw5qP0UX
BfhZiSikdsCwsSeWZN4i63jd+JiBe+DtR+1vXHI4GlL66pINYG5F7O+BMjmTX2D/
K0fVKdM1BUD6ynHr46Yha0FFA0EXYCqFlzlbtgMGTUwSODD5S3MANTK0vivsIFdr
VjinUNqCt/TjOCI/FIRetFssoBsEXMhHZMsssZlwcvLsBqQTlvPXI8GeIMfjdjdZ
+y5l6B/5bK/nOxdWH/wGz/joIf4LlkI65AhIwA7H5LgPbBdp/lFc2RUGddp9YnO2
CqDS2YEJlnEiEBlyk5ikrNaW3JaCV8mdZOZmyDjyaFd/TF4qwwg01S30QX4MrTEu
AYJl3SLvMzTqFt/bKAD0ngrLJCZ1SwODd+V18a7TJvavnRex3HBMHZYMX81ntNZ+
BlGWPaqbALpHxbNxTi3Nbd+tooaDy3a4UFYF+voEdUsIqWIRri1ouFCcwUkZzxEJ
V4PQWjasuX+v/PGz9Hary/LPE48gZZl1GfkF+fNcFrgcXChP+V2zhTd++UvP9nZa
eNuhmioUwTS8On2jxkMBwhIXwtMYwTsQOk2AtQVK1wH15KlPN5ieh1LautwQ6OSx
DztWPE623SPNNILI1VWFSLQfek87SlPeNa4LWZS4tZfUmnVRAmqzCjdPef9ABK+/
p1/9SGh/DKxEZ1uYQSILlH3qVxQFozYrrEdY8mEKq7nxaGKMbKZavMDQ29txyG1v
QsNcO+m24Zof6F5lTh3vx4/g8DEu68M1t10cF6aWNuqD+gIlSoIUsQ+2ynBuDQit
4xhL3UkT9zCwGXL/ZEhoJKdfpmNHJsiYDsP+oKqE5uOpyKQjPAgjv7Gx8AgWGjsu
x4iYMjClp93XyUMeiRgMgZpQikH1ldUNNdrFXJ/jQO6TpR47Str6LON/SwvGKfqn
Euex8KM9sQDvBwrJgU6X4RCxPsJ9rK3St+4vMMwQBro096BrgVFP4j8FecHVvpfZ
8oN+21MXH34TehK/HEbdGlyxipqD9DZI4xMKQ0e1gHxPmkRHe/EBOcaD3PwmiynI
egJs0dnMVWizpJT90Wt6eci38Cr/RTeSQwp0eYv2l4NAsxkYrNmHpiAaOaGRLU1f
Q0M14CC57OTbVHcM34C5SbyGRrieNQFkTEzH4SG0PNIx15wxgNyksP2Hpwm+tVyd
/k14ECe3AJ6SqLzrwBUTCoC7IoWtHa1T4kthBN2cMSGxrMwhW1ay0baE5s7QY3PU
uplBcph5fZkTAPPa2dWjF0JtDQhQ6wD0XZJyBJBY4AMElAW0rVlw51FjNrK/69eH
iaYHYbFK00adaN5Ik5E61NXfPBTzQMWP8IfYTIa3oTie1D7HS2lraKJJfevv4gNz
FKGXko859V3WO3LS5R22uVzqkL4gT2dZIvZj9bm2wGvm6hgHctkwH6nI0M9QriNa
6n55QV7y76QoJQADsnXmWMWka1ZdvBaiDAIR27yOlAzrdfBkrJ8wEgEi5ttUSWRs
rCSo9XboLget0ie8ll10Qp/WuiSptpIit5BTEBj19kqLQwQBN1KXwq9rHiK3Uknn
Dy7b2VqkACyup+QbJ0vvbBKIgkYTSKectdfitleDSduwQeucwkG5kvt+wrOEp39+
mGoc0t9ELMLoiQNgJ+x71eJV1PPh+ZbntVbsEv0ppzH8uSUOpdQ9CmsaqmGor/8y
TIRqUK6rh7m61pQoFvgovjtHU2O0ya9OiRTwFasfX1mDRqG9h8DVebyAyh7FwZMW
RgKJQZ2Tz/g+I54rjlKQmuy/+WnaxjOPQktmh3XeqQG9C9XR7CbPHPXOt9KwLJM9
EpxpeRwe9yU1LD2ztgPpiT8OjNPESDOuRnV382u56jYphk5SPSItrX1ZFc4Fnh6c
nzonwNUr0pTbnLW4SN5tPuQNs0ba5tiYh3bcOxT5xZitOcHLrvd74aZfLcvdOLwh
623DQUKt++LvuinTJHrLNntu6Of7T0xFrt2KKvbDIWCUghgQ7AFkTzRcdaEj9qk9
t7uB0j5XPpFAJ+zaFJa97Ih61X3vG1Pz/qYfnWOgvza9mGWVPssFhdcZZWB6c/QP
ETqm+VeRx1EWzXqNW4pydjugbN9cz6u2v2TZBY1sW/8avJXlisBg/oN8UWkHev8F
at/+Oi7qX/PDBMbbFyd1bXZrlh/SrOVZeoQH+e5DaoCVii9tOIavnupOhvcu38HK
2jXFFKj20XTdoPJL/aCNABnkP+bTq2USu3Ubulyj8ANluPrifUeYcv5bn/Z/SAYS
kEUK5FzA0dIkI4R3zlAtdYxKJq/9TxJ/Yx+cREGU8sDcDvhXYe14gdUrPQoL3KzI
6bVztnsKs0FvxhxdnYRDLpXYDqAyWp282SYlGlDsxlkinbWTf+XnWtc9xVJPHd9G
1FKv6qy8xMGS39erHavCmWkLr0F2q5zMySO6Ay/JQgU5bk7YcO1AYR89PFkd/ok2
XebtTrX9Qazf//uBsqc331qc3PxwSWUBFp8nXx8bV25QHIKvFNmuDwaWJUAL1YK5
cJC1zVUtmr1+Z3lZPpYlcxOaVY+w3m+oWcXwvqcCyuItUx2jzneB4fyuXPCDhFkK
oGad17w7wIerMjF81taAZ8ppacKkx/IV8Ccyh7nyTfKHj619QvnAowR+yDILwhPE
Me78xtetV/EvTYbTjWl3Tp+lt5cWJc/nrPrD9R1RZXsSfd0lNN3QNN0We7EJ9nNc
EoDSHrnUFemHV0d59hHi//pkxt+mrPJ2zLjmsvhsPoK8dBe4dP1avRMDUdp+D02f
3cH34RAevC9YpASHRlICJqnJdWUFwffnLtKE5dCIRh2xLqaawBDxBWUfafOt17Ep
ith8BGsm6RFJfb/ZFDuDKwiYsl9iKofV/3cP55qAyqwcdhPMB39O4o1cxoDymETd
NLKyvMAqVfQ8NexBIGIEsyHWv+AEe2R4XT6SpSnORhU0jghZ/nrRw5jGdKlGOtJc
odV5IWq1PtegztcoreNMMnQluT2WCJgzyqqxwEfUcy8XDexxs6SBgWxX0myjejHI
YW5dQTEDriOmh97m3bWmRqkyzq+YGKQssiOgBe0RosCp6ylh1pQC7yU3mesGMamE
l4G5GgOBG8B8GADf2hwdHStRkrrbVrOO2MvXepqz1PoNT3aQ5WP4dNGLtsDRkrF5
rc9iFBIOAAYbIFFN7WGE/7IRoxsyeNGxLdaq/Zem3wFgjJn2mjihkYEjcLHPAF93
NrqHqqyN/rgiYbuu063/g0MTu4wGcILOBCo78PJMVEWDuHbP3dDKW23V7+ale6Ya
4cZxk3xcPftB4duvf3F6W+VChQWTrkkQJMnOx+y/U7Unu4iPJvC2DLtkaiWNtbdk
CH0Cjb5zhH/V178hF5jH9N0xM4ShReoDLT1elPX6k9ZPDUWv/OqyM8qoOw+kY0bE
TkMK1vyTL2CF0bnSh/sslnxnwrqzm5ENvIy9JBfzBxexU56c91ptTVK5+/Eav5VU
5fXNqky39CiI5tpEc9Or5P1nDllxmlUBFMcHMW1wbvfABErlWh9SmIGVpAWzOtSk
XIVwqjfJSYtcU60A/Tjz8zbtrR2rnWeVpHtepVfSfzhWNR1Rlcw+JD2WgM8Ka3a/
aBC8zFTk1A59kgMBi6JLbUp50Z2k6piKflPPi92DATAHfJyfF7or1HcfREHJO0UJ
Kv/Mgq3JAGwR+hVPWb3EMCPOocSuCiIFauQVAJcBcOZDURONYU6fI47bsi/wFmmw
c30BPOB7xo4p90+JISPpTTTDbvkyYuYffoq0fxk+NPEX+bbmUwawZkonFh0BAtTE
rs5lV0rdwBGWWXYHYnqX58qzzP1QHACG6z4NQ1rAFU/qr/9V9/MspsMGc3XUeJvd
Mzh2iKxy1xrpKxERb/ag8qIsii0hxgLGKGukeJFdW8ZKz57kQZ14yIls22coCRqv
egjDPPHDlx6QBeiVy0oTB5wZQ6e4dDjR8RJn8sm05qwodq005xb9npWtAYRfldry
ViIDi0dTE4l6jUo22f5ZceEhXQmPFdZaLIQkE5eGlis3K4AOQ4cXiLhg4m3PMd+B
NqQfpR5B49GhkB/4rtUbwmxk44SgN9RvQLCRLB5N6jM+Nyhcal4TBy21QE855Pkr
Pj3wmGkTATQPmUkE3pFbB+igUvlydAIJq/IhVApIrnifWRE95HwAPVtF1yp2Ckpd
Y1ZuR7c8yUo0djBnjvrj+7Nm3857JXUIc3iL/Bo+SOKcTKIxTbH960S4B8gx/99+
A3zwHCVb8Ta4UJfVMS/YD/DjKNtckdkflyI7VvKNBNm23cU2BCpzgjTMnTZB9hEZ
pLmOW/x7jHOeYJ2TwXdyidnwMbz0ihrWZvAv+OQfG1XHMM4NE9YQuYYvTaVweLBi
jKCE0VZvFBBTQL+p+RKob9joPIU+YQg3BXF/v9XIM9h82S2l2VYp9nzqg7jsgQhq
Fs9X9ZGG7Up8MxqBQ9uTqVfWahU0ly4h/hJW7ATqbYpEVHP0KSHd0bmGOCo5Qaxc
56cKInqcKgXapWWlj6Sy18k5DC1p0BPjHVr6WyG+mVlPWEHMQ236SFmNwN0UGzTC
5eKbf7Cm2eD37hn7IKBZoy0RN1JnXH3SZ5Pw4CyhhFwFikmInu26gx3gOYgWS26L
yni54leoH/i5iXs+N9dNnfLrGFmSRO4JSK1G8CU+la+1W7+7iksjGamLhhQQSKv6
lndIPzuAM/neP/pLjTibLAIExcoFcv4ZjHJSemLoKM+Fp9Qy6t7CDov1SiVW1l2U
zZ3UO2N5n9ntueeKtq8yFyziYRQKB/5EnZWHacFGC3CrFXaXGfzlpjaSge5hU/J4
5veWEgYBLF7ZHCFEKcgdzWKfz7GMr/Df+tsYOHPCyPCtk6I3LyFKd1vxl3IQyT8F
za7PGNWQAo1d9YGS3at7jTG9caZKbiw86U3GwkPMfX/QrjjIAWYkzaOxBm12fOyP
7cW9txrS8KTQsBvHoqs7iHXT2FWM1BjnpkokLAwHsjCbqb1mIc/2v9iFTo5CGMYI
x/3AzDSemD6w7HPecpDvqH/dlxbJTicTAgruCb/VEgxy65OgV9vSkkfvABaQp5KP
QlicK+aTTgpOYKC0VE468tmoO9rODtI33ufkvFUrbNebMG4kAiEj8lKwX0ptUg46
Ayo9LM/Tv09SztsYJsqXeLc0tiE6rdLt0oRI1xfmolYXe6aWVyiR5tCQlWK1E8/t
SF8wylMi37oi+4Ofa+BVH32wvUIhwvcBuLubsR+eK2j/8zfVXUd/idsqjZvxpjp/
HpXI4mdkUeeJJVQa7GNAIvay/LhG2w08QtAJKmVRPnigITodRZ37Z0tM44oG5ptF
16CNUUcWp//vSz2ExxDPPhz2cCeEpB8+k2II49PBK3ctjylZdVcxVoLtYiVt9sN1
nHLwO6NoY5YT5MzPG7DJYUqBBhykMQwlq++VTZ+phT2us8R4HHT/tKJGP7y5Vljh
xSU5RJi5/6R66kJ7T49bhM/KU3XS3Df+JSr8potzKfyElDVLxVSwpGsd6AfNtajR
J1VEX2v/EFNoBInx9eWB6eWRA9Wklv66arZJXJ9clqcr5q61U/WU5LTjA/IFsp1F
gag89Vy/nFHISbkcw5ZRQ+TT1mLsCuYSD1SXLHwmDWBH0RYMlI0/QC4osF+YO2Rh
N1cfJUOCbNB9sKD782brJ1ei1qhNQ7WiNHt2nBXxY/6G0szBFMLKkvTUnAWJfOIw
7rB8s9E7ORStwXYwQNCI8eKYT1jfgTCKKh3mikKwFkkTuts3ucCixm0y3+yAP37u
LJ4LdJW2wU81K+EwQG6a1F78TqgQ3VZv6K5ErwNP72wDyQu/HTrUJ/DtPksh3JYr
0/Zvo2o+/pWVNJI+L3m+VcXbyrFdZKICM/jj8fDK+dkEVyB+shuwG+337uNAxBbj
vtPRTBcg1i3S7YCVqgUgjh3lojgMzRgXtP6tfK0gkgfIspr39V7FHbvkWm2vzgKj
kf7KjEjC1e/gAlTCl45VKa8/n29WJFxnuuD8VqnYkRtxkXTM54nSZapPVcoj1yi6
Nmem2tfCY3PYUDZybAbWzlp/bzOEIPTTWvwSM8AXewGs5l293xLZDYSF/G4m2BFM
+akHDP6PyYY9XkVfz1OGbPXDgOsrLkkLym7stGx62Sezooo2/afbC5k25Mkp8kAi
k0dpMmjzTUIfgAXwDTmoS7g5YSHTgzYBy+TZnyRTu8VG4ZUMbXWpG9z1WiQjJJOt
qeQgYKZ+ckTEPBJZZnsHuQjZuAeEcxWHfefM4B4Sio2pR/xmbqT6eAgWxxZmhSJy
kbOw3Mi7iHKbyIui6VGwBpX2dG7AfL3gfepFD8GDrcSxI2w7/ThpJFBNVuNevDMl
AUheClliG8gQpT8qIRI35Hxlnw6Ib8bwta6kxjJnbNz3YDmCYFTy+wJseTN5gFnK
epE9W7Pz+3Y2X2HA3NzoDpGljNqfp8EXHWnmdj5UyBjIf3t4P1uaPwfXq1JnxTJG
U4Tl+09zdjXg4hLxJgwBC6cT18HPSM7Ajrg58WHRn026TQI87o6WWQ6bEE+kH6AX
9EVYKFjNVINmuvvts0ItWi/NErv+UZW57htMU8E9ZVgjpymEl8QBqfFEIWTNPWnR
07JSjZ1rWY/tbz/X3xtNxwCu+TO2vfzTJt2XuJi1AxCvR70iPFQQlLcjH9XskU33
/dc3/jc8PA4klrq6Ais2bOdBf/yMLHpMetBB10CEdixwHAFzRWi05GkD5KoPGheE
AVRVkJaPmKMbbbpECU8Vaax+oVWBWaTJegybZUGFtQtApsWafsySboDozZosvieH
ymp6F3FNjU+F39CYgLAhVpyZQFL7nvENdcreWHjTx2DF/sHXdR5iVr99bnkaiDdp
K7g83MmWGlcMcVUi5e3rm31A/lBKsxXu/VejxRYk2ym2ck95nv4SwkFYXeQim+QH
wY2/CR3JJzUE0rYykCaKxAi2Vo+Ug+5OqbFQS8AokZMDZ5wei0Q12lIT9cfGmcG0
428I7wct9AP/EX4WW1fpjYcw+s1upivtZSsIh+tU06zCD8EkZ3KUnxzeuc5mBxg4
tLvVMOablDVXH9c75qxAkqosCJWodptL6i7CxfOi05ZYsDzkWRSP/u1WLszBcT4H
reNoxdLqHVlcRBHUECshUG2xvMKXU/HxbM4Iz69TAKEQmXk5TPbYr0OCj6jXSY7k
qwW74xYb71Y2OpY1EgieJxJuNotB08nq+ET1wjUTmOXbARWT8TDWienRvgf1hXhs
Q/fU3QXcfvXRjaznt06cypjV31ojBKcXNFmdd2DHjq87tfwHiVvN4NynHz2M8AF8
fyOxGTFFtWaOf5yNGh+Rg0M1hPFyo1oINd8rltwCM+79LmD7CxUiqzuIiXew9coj
U8gs9mrIP221mPtSFhsWAIJNf/nAeqBgnGE7wvEy4eGXVTNphC8f2o/+Lqb3OxpO
Nl50NCnE/5kbTNfZDnOvrfOsTP4Juzxjk0Bgfa5UWqszBufvGqAryePYweJhnpPX
XAx4nzfZJHhBHxG28UXb3o8DViGPYormoDzvPsmzhfRgiXDpZ/b4IL9uGCRmu6l3
MSLQsLdrV1M1Q4JinYj5rncta1uocoJI1rHfOVWEKLU+wyU1fxB/6+vxe6pzfhnr
k0CmnMu50qerwc6nKtOVdjIwMAYyZ9KlxvskQ3Ylz++xoJ17qF5gYf3oLNe+z00j
TdNxmNt6PeBCWNR9chxutEYomCoZjuFPc4mfLjDeivGXqIqCxJJzXMs10j1vcgW/
/nXiM85RTae/yt0xLOU9/uPaW0aEGoXp3fej5ig5otq06X0fbI8UG1G8sMrrXa5e
ahqagiyQyXdWJMDadUZFFaHkLDvO+p24hoESfMvrSbMBhHm0qCWlTMFjC3MUsgDK
cen7PHS4RsZDwGpPZbp52yBKivazpff0hD8MeuQQ+g8EdYg9qgddOYjIRUbm9ntq
hFh9i26pbSQmOazv4N+eQ/Y+5MSniLs5CIU92RY25CXp2kZ7fbfjhJuoeuh2H8Up
V5prMGPXTOETzQeJ3l4i3zaL/og79yf0NSeGMvM7mcmpIG7CAJyvSZv9K6LccPG5
YJ7LxkRGItRFBeOTgLu9879OWaLQZ3ZOt/6zyd8Wu3uo5mLkSkcdbCJ0CdRq4ByK
5W74pXUN40mZxVWki3QYlZ3wJTKCXYJWENFV0j3sspRLdGlRSlWYFEK19omi5PDf
zwFd39rbAOnf3Zz/N61sHHmDFu4NCahJHQQIog8ka+3Gph5UmtAM9G3nqXaRlI+h
zeo1gS8iNjYHRgJdMt86WnIzfhYWDqtesOGQQIpSXLqH/6u8CrJHIlhmIOS/kUI2
cBXsvCPHeaNk7EWdk3hd+bpAub54/CFeM+rsNTNkOTOt4JyFnbVAT8je3UKaO7TG
chj1v5+bycetY5NqE8N8AT+Rfpm/65j0RlG7jg4EInOtnxs0H3kl2EXpC6DH50uM
yCVCJDLD2FrAwmbaOW1ionZRxmOgmzjiehetgwQGk+Y+sYDlIhcgYrJIf8F69Nzn
5XuF4exfHZuws0qu4NiaeAw/IscRRJ6/lqk2Xhm64UcVwAFMwHND6L/1bludb+Pq
PxWZHmCm1FGIUrJuOPHTZMunojczINBOivcWkXRvkUyIcUQUr+3Vta9yfB7V6FyA
gLQHBTOMjDb6VHEouv5Bnb5jq4yV1X/5BEFOgpXNuJHiGpD4qkZko4S6J5DO4fdm
pbUvQDdhSiDsh6wticWthHqPjgf8s/LNl5IPWPwGDKvKzdThbQS/CM597EMNV0y6
gBIOG5G9ssn+18vwSn/5X/8PB1yfJaJHVf21B57ptSy6Ls22hOE4/pZkGW1EX9+x
1+CfHs8kpAxkgob8gJbLqFX5XDHSM4KrVdf4KwOUYWOnlOlB5lsRJtf/arx9Ahjo
CAl0bTL0lKLZobvsvzEHx0qTB407rh/RXpDQn+/OVssOA7rGaxUJ6aSJJItb5RhK
E1Vp07WhY8ShSoiCbauTzTtz51s+g4nSh8y9VdxbD4RPPwOc4NkUCTFUaobSt7Zq
u0qQAvM7Kiv4NSm35YMzx+tKnSMFvipKq0qsIJNnbyImc8yzI1rgvGF9g7+7efye
PSk9wN3L5oUIezF8H4ZH8CE9Wq9MqleYvMxb8dDhNcfCLJAKFtoyr+IDFC5MPiKR
qGiYZI1Grb1BAx0L4BqMFGJuELOkNj30J80d8nDygVrT16wkmCaGCzrp2iVWxKDC
ZRfoyYlnirvxbHmHbD92yU3lMlk8ERLsZCmf+v9ZI7s+00x4sOM20hDJIUP9jL+0
g/RPlKMj5GLrIdgsf7gBX354/BU8xhC8bkJSDNMP0Ic89dhZGW2KXQWNSblqnNqH
SLAgw8UgqVFD+1tNPmk0/5J0qG2XAyf5OvJE4MCnEWTzuH3ba71BuM3gEqrRi2OL
FAAU8QHlErQk0nQ5jnIWIb0M27M0iZb5ORliKfIXwmDHd5PxkxRlMrD9WuqJk9L5
QthpmyrAhYWE1bdhCsq2oalEtXyZJxn95OLcO/MRCAm27TCY+YW0s1YQgvebzi+Y
/ERAO3VZfNwh3sS4YzxbuMuuGtCiqvxgIrWMiLnfS4tKwY6nWqEQfwtmgYiVsC2H
lhLOSZj3Yg9m4zAfmOIj0PlZnM1NKyclx74O/Q1pBDyWOwkqM8iXsmvUI2aD1ax6
kr+wn2DAzZNgCRhlF3oXoYphiAYytrY28jTee06KbohA84M4yetrE9svrBhoUOsT
gMfQVioBqo9nvuDao9aBj4CDe6O/ZS9pIWt0kXmnDiR2UC9CYcVf+ADPU6Kgszr9
WWaR8C01JlGk2TOZRAzzvKM/T5fjFQsx2ObqUnDpUpytRZXBFgPuWP1plNF9x5Ds
FqGJbwKM9pLmrpbt/AyQNB0u1kfi/ZbMaBuIk5451BWioflkqH0klVy5uH44arS8
GndACO5tx+VV1EY9T/jYGP5Ovd5gy5jUi3c+NoC7ZJNunnKfWwVMl4OhdR7eKJMB
XviDA07/oekCkQoSULOefxPgZ3ZYzTycS1X0+84EJt2o4bXD+Na0EwSed+RKkfU4
a5byFSi3O5XPGsCnZhbHtfva0iYh8fUzzPJTfMTSjm/YIPtwcsp6YID4b1AtgQc7
fGEe1PiQpxejosPlhg3DCueOGHo5Wbbg8zn9jtng/Gpzjk4EjMgANZBrVW8w65KB
io34QGJtp5/aur9yAB3mAxfVKt1RV9XQMF8xRY7df4eeYZL9GJomJYa6Hu4a9iFq
XgWuj5AbyBN18n72+/6RMXuCg9qxcfyM4qaazvhy2iIrXtbxkrOcXsnpqZVnhAIc
g3cD+9N8c/EaOtGXdRe+EshLZH3g6S0Ho4FPHx+QFf34e+B6p9Vk5R81enOVppEV
nmyOoGQ5RnwLvJwos5KBtEk/ynBgHGxuQ8Sl4frjnSlHcqiPsM0znxyYBErwE2CB
DScfytk3YKJC1DFYwGglE9/11Mpbl9ZK9+G6iQISyaB8fkBlKE55e3ZONVWOa5s2
u5+mqiu6prj9LwM2rmqIS2GTidZ6pfF84eCwAyQlMQ3ptew38cM3aUVpSMHo78eP
ulHft7qo/HWfq2TQZfNCB1v6wcjXqy9r7eL2ryBp5WiFvKAPVu84sMTJV46FwsMn
SRxiaCljFmci1lQGuGrrQ2bteMSguOD0NxT4bhBwDL67PoIdmegYMdoPHTRi0c/f
A3WoH67CaQCXBWgwIZMksU7wMy0ln8oII6nnIi0DbETZKVeb12rR36jNgX3AS9TQ
hBCLGanOqLOPYWLwmtanq63LSHLhfl+6nBLlOIPrY6smh5CLvloyZlsBHyBwTgeB
RmRBLhp7dqwl/Zd6S8SFWvm3kaUw+TVxXJ3jwIErpkN3xbDNlvCTAAx2hr+NXjLv
JPjFmxOVNwXjVjTsi244wWPS91O4HfPtcOY7Ez4QjB7JZI8vULkkaqAksnftq8m8
kdmnKkTab7k74ZLqxxeSMsi8Z5DYqav/DNYcLIPKuhlTYn144Mq76fERLiE2zI3Z
QxnhV5Ivc8uZR4ps7GiV8HJHStEH71NnnWRcAY0zfPFqVkb2Y+ge/+ExGN9k4Occ
AomIHNpYGtjhrV5RnlVFWxnIEPtXOgDzEgixkqFwC+6bX6AojjjhYk/k/QjUGaLy
eNhnlpWYnE3R0HOffQUouctzZiH7/FO91j82Y7a6k7r0PXoa/+QN3YCtSfjhT/1v
NVIllEcVPzdEGfmBDUFHTAM8L4v956+SVhkLPM+oBWhyZB6RvIxjltnBfdIQuon4
Ob8swOlQQFd9gw8+7ql5bvaQHuU3yBUgVB75duZ9nbdk1IDUtRoOis3MEe8egxTW
3/EoxjmqwoQ193cOpJfWz0MiorM26TTCizHmNHgRdoAxWPt3BX0X4opWQCvuxiwM
E9FRMFw2dphBIgCxGvPB9Ux6LTG7NMgPHF7Ti6RfTzo5AeGyiHK2RUoPptg660+t
7FC+4dSkUSkUEYZLrrM4sCJCon6SdJHS+iYAfWosKxbhhTEjCZM8C/NJa0JPt3Ik
BICzf8GvxgTpVd45jrxIsRC9rMsPoZB1POh8UGtxOvk+7nRyc0DkJg1Lcu02vpB7
+F8Hm1HRvXJoOKXjTFZH62rxNH47s3JhHMafw/QB4u0X/j8tXiGwQpyfJB2KjtOe
H/yqJDBM1oMkE3Fd0MqAxuDumzKDLREQ2OhvA44WjbqZs0mxS0ZUDWqYtxdXu4kr
CJ+h8ugrDjWO89hxikwrlK4Gv9Vthx9Uhjqbs/PQ/vKjX7602Ajn3Dya4hATzzoW
NLYKduYCqCoVVjNSu7wpi41OdPWfGqHWoKk/l6XOq0WeiOk8HMdfsQyKiIhB91ks
0Ap4PSbtuDXOgBWBZbhwemAzr5RUgXtS50BRqxZChssmbah2uHfIetNehCCmwIj/
jkRouT7bMU0VmhcS3hkj6ooEFcc39qhq66mQkyKI3JoLvbsa9zt2Rq05B37xtkvl
spLlmFSAZj//H+qKfTlq8oty7K3ghRLX6u6xy72EUxqPgRUk2a9zXwn8ksFYUMVC
z6gYCbCZjcaCQ8Hr5E3H8Q1r0cyg2XYa5Fi8VJDkxLkQ8xqiK7Vfn/Iw0K/ceGOV
RZsYYnZNgIIPGSovgE2DrbfcyTAfkgDHgVzwXqd1028XZkJrRNvSNIZXsEmMZIvM
6s4AjdUSRiHKqCG6UIKt/LOIO5lDjVn1gkrkqRNyS5aw0qnm80vMk8sf46bz/ds/
8gFrpY8QJ+o2+VhhyXy2sFKcVsHwzG0zhW5oUm4iq1LkfSA+vN9TAOIHS+aLbxlk
thuJkLySGu8OQTe2nyKjDjmiGBKHqcitrDulglCq2uSo/s15Zys/Ql4vboEDNDl7
o0ZZ7SV/qVZlFTH1CcHDMCWsmNuSzpuqpjDLo+z7JVacLfsy0JRb0d3Zuvdzrkk/
m/WmbssZevIzN9cjVK74xsxvQhznp+uGqueE+Dv28HBgC1DpaUTiwJnHLVcPPy5d
u0Z1dNQWVyDAJ0xORTCcEVsOACsLkG8m0gjtR2HGFDficVqFe8gece1w5NT4JDxZ
/w1UcEjCTOCsvCw2CYeMKhn0f+6r9EpAyl04d5qB/w72tWiWyfNWGIfFsHsnoSoe
ejWTIJS2AJiXERHs4q9jzR+KJFBfMNj7BVNW4t2uQAr/0/mJZ1yXUaN2DjPr6TLc
LJ1bo6jaDMLnfhK4Bbb9PSfPJiFvGDJH28kJe1ZBNjIBBEzPcuhRd6sHuwgQvE5h
sBOzVj4EhaaupsFmZ2XMMvQoAUb6vKbsP+gUWeJ2rWahrXlcSUsjC63Xg2HOX/Uo
JVV4sC5M/ujxr6ajsJTrq5C4HiwfmPKGesDofm+yIEKRgDvc4fjAv04HAGof7IqH
PWPke4GGADO/e55RMbseFvgh7sVyhWwAMeyJ2dbYV/eQIu84yQqzLVgC3vjkObwA
9EiFPm1c5Vc51kxlsE4sblQqB/3KKKs59ehRLJ3u98v9EQYkYYxBDI5EBGGL5WLA
ZiOwS5U9MJ+ZFZHoRh9IKllRLhRTvmOQvj/XY21cG6ikT3ilWi5rPP9qfbotSJl/
kmsmw8/qT0zBJcs/c1bak5GaaYTkGJff1jTahwc8UGl6fyDjYIfxhitqdwmLxAh8
jXA7cUvRjfshlSmi3M1c+GexCcEgVu56p5N3Qqep8ZMCRXjOwkoguJ8Lem0ycnu+
ilXPzqR7oEwofrvFb80yL+7giJarmOskomg02uf8EeiITdoAXciYZp3IBPzvFdc8
xsSogI6M+FTgx2P0DjPLDmYC3GPSZOEpHb7pcVP4XqDX/9b+H2f5VShaeLibpekA
Ck8i3MV/kP8/N+nomJMsq6D6DYDJTmTn+LBN766nazA/z3xZhJBgw91daPJD03/x
o099JUYQIWj1uJmQ+0BKl1jwk1EOy6SZgvGNrHhzlFQPwKwcTBoiym+mKQwO6Qw5
67Z0QtFgg3/8yAiPlshtM4DlyIQliDY1Uzo8KQ3ZEpYF95WPzeBOc7CN2+GWpwhj
ZzSmoQPyoLtUENcXKD7GR4AP66ZcxGs2TIyIKDKB/2XRm6/Oa5+jqMeNclWklj0Q
GkaNDiw0jfcBHMPqSrctpeOTZgTxSwspqHBbi62d0ZHpiyFxFIMbsorzs55OGGW2
OXKeM5O9sAq3kvXExyDodi2aPVVo0vGWD+QpvneT3uJgsyCYvUh/PWt6I9AdpvFg
4QokrnYwa7XuESTEP3qvXCfc8V6fiAigN6i4L7RMrP+dV+ypUmoRUaddnD6RJUW1
ZL0jYhYLwLQILWadVxAK98lgQMgL4hvymbxJQglBSgwH6iy1ibijxYYHo+Cn+8wU
G5/GAdQ2/qoQRaZlxpKQMEFLuEaff26KF06wapQCsO3g76nfJ96wbQjVHMLcwxg+
p5DHvWp9T2P9570T/kDzkAujJ5yURqlaCBiLiO61wafpHKRoBwgG4k+VJcvFu73X
jJs8727WH8xHylm0RrkoyPQtl4f4Evxcw3eyL48+jMMbFogGX++5ioIo1xVFUzye
O23NwKngyGHFYYLtNF2Mo4xGtoRcncQSexIqeXhtPx+gaepgNrN/o3nyYk87uGUM
OYvtjTiIj+eoOk2bJyDCLplBTWvpx8C2CxJ8w1j6UoNZVCzbb+9fUbB/dkaX2GQs
bSn/mH/8px4E6AqQ2LdN2+9fMboYUhmR6byro+SycMGTv1PqIplj8K1KusQ1X3qS
NkxrE9nTH1yaCBoyVyyaBmHSypVrij+LXHKUY5HYXm5joDtEJMluOmQs7y0TG+Yt
0oKRquuTHQSrNbgNYTRXTpEnkCzn14hJ/lepCU4Om+/oQgCHUlWcuOj4109qRVRv
PNshn8c2NReXDFvWTYpmUb/KF+RSz6OUfr6fbQRfEUEt6V2rPf8cim8ntjDfuKYG
WuY0xsWX52eWOEU8GALtbj8CuA2kyWPE/CpomXCHweAm6KI/gDRrK9TXOwn2xim2
qz++KFGWFx92M0UJ4t9GXjxHrt1TheKAcaRrdu5jvo9aVJsvIuHwZdZZDN0WM5Ul
LTHTChC8Shkt1V+KBePzVXEEDMxSIlR4mfyl1lz+CqUO46cN3zmd1x3xLiitQnSi
CkfxiV93viwQyGc07AIjCk2iY3YRNdzOqmo7eMrNaKCP05b1ufcWBHrDeWApSDB4
MxOiE0Ee03naFNc/NJX3sZWYaIcH9LJOYDD4BAGQgZmUn0CWW3ibEZ8NvI1STWgR
d/neptksb5VWx0F/cDvLWsEkih4eaHneeSCKgQroWQFn1UTCW9jbyokYjSiSQp2C
H87Wqyd+yKituiRfjRdc+aTI6yZn2/FiG0LSq5fCCCC/LPrtJNcrCvIvleNufya2
LRfLUgi4DTbzXowIOuOfOmQEpMXoAPIq8r4ZuaIsbmq+xJR6H1h5Rg8MNPF2IWgS
50/qRoGGH8nEQJ9/nVrAp6J37DQtEvmpH2MnseRhSXT3D0vZBRiJUud14egMTJKK
X9o65W5bYBTkGEOlE0c+g9Dm3LWuqXZE6m1yBnS4mJXO1+NydtAPppyEadT04M1e
8KHVxUPe00hBCCfI7QCJNvPIp0RMHG78fcXvsiY06WZjGaHk6eLTmV48GPSnKvPT
vtuz5kZ9G3U0GRDCWHpwHUfHWPgeTUIQTMkPCN/a2Ite9P8OUD0/Msfq23mC28jq
KCYOxLQvqbXUZnwkkbWwpV6599lxMd/u1aHRMq0xu49gUineMsob3KKu/9QtD5Bi
cOUrZEVBa3a7X9G4wfbnGmgdU0I9YCFawiZ4R7oyzf0dr+U1wT9WZ5QbXJZGK8+Y
e9lNVqeJiD7EKWmXxImaEpYe2Miuos8J8W1w+0eC3x8i41FcfYnKJ9z0HVoIb4aB
Czg3GRZ42+ObBL8z2d3JGIFcIYQWGM6w5egkT7O0zNuU5ekZACGk76OxQgt65vKN
5GBbM9fHdN6mAYASq58l7L5lcxbYJo+N2jQPKieXKN8lbfwSVr/7Uo/u9/f4ewMo
y0ZC24Er/zQ6shzyi1zSXSGJ0snyjd6WmJyjQwXH+8wftKEeqzeWgIaw6GaqL9oD
pDrI5K/6maTfSsgpL69VfhmoztycM+owcM/+NUd4HY3NxwJ0amP+oVjRZgi50Sl6
lKXdRWx+kOe7n05A4/DoPAlWX2jGyR71/OJJd7VV4b9nyg8kvGEB+XxmSolSFNWZ
ZFFyAGiCnGZRhC0epZnK74LSdroPYPeJv+4JHVsMeKmHm6J3TfHlUNmzBHr1QUpH
2kLtqvrSMkydCHR0wjmaybZAqTld3zT0cIDfw6ytRqPEU+evZGfalSwkOu4bBFhc
4AGqoDaT17pAqdfMIh3lmItnmjbVbFJlVfUmX04uA0+j9x1asI3pIk4hnxEPeXPM
jeZNUC6q/sbqysW+yb4MNbc98O51FjBbt5JTDRFUXKC0loq0i1DN/HITCdfs107J
pD5k9P1+XvNqaWYAYHQM3ln+zzV9LqXeVT4u06tHzUW92g37xT2m9pChkrj0ggmX
tXa/acsRxVxTOpRYyL7dtFrownNWoIi3lgZ0pjQ4ZrjKq66IYpbPD6EhTON2akp2
WVHF4TlOcRYsLqW3YrDk350+uo70Vx63dDBS/SVrpWRxoFzJKKpqGpkkmtRvUJf8
BP5oL0gjXLJYvani5GCa5nas/8SO74EphdMlhzYZDzpzt3FI65sBdFRTKgz0e7Pe
4XLnONX1AIpSYNMiD7FTQD9mtbrVwwlRpqkT9VR5dv02pVtCvwprliiysMixRf8k
YwZ76lu11xGBfyRwRs7R1Zka+ziMxhmpUG1WK1hU1+FU9vbWT7RNWMNhfEw3SnBk
ak7TJA7sXkoV+iuVJSaDOjxd1reexz6/fmkYmke8MLGlf5rnKWgZmzboDpOZ3CnX
SZaeQ/HWrhP2KduTX0f4T/5lnRZ7nFLFx+jpFsyQuI2PIyVp0qcE0uckpc7cbt0W
BZO38r8/ua3dON7pp4PAKxnV3xAvlfiL6mQxSNTZ/fhWD/jKcDmPWgmDtqPPIFbv
De1KhvNwa/8N7ds2Lc+1SCiToX87yPZ277YJcYtAh3qJLqETX1SQLbp8ZzVEOquc
LGRxQXUydmO2oZZ2jipHS554AmoETadKOkd+Ces+7VEWYHQ8wXDQupjkWCC1zh8E
dcnvcQtLi7byZPE89060G8P//HCCMulhP4WQYFcEzjAGsqwH1EmKX9ZjoZuA5G3q
1ep4hqn8HB8xujcRa5wzAVF9hYUZOJiqNraioo/OYzFpj1+vtZ02NS8Bad18ZN72
heXmwmZTNj9P+3IR5aXVYQ1hDPEA1DX8Zpz01dVObdZsi6jInVq9bGiDgeHBra1h
1SwuEMRGFMAQbn+aw1L6gBtKHYbIBHRl+wG8nNhdL4JKJ/42AD42ilgxQkxp+dg8
80Uoqnx0C8Uv0zaZKNOJ3wHesKBTLtVvLqZ0mPGavZpD76mvlUBFHjwdJcctBLyG
/3BNRPtVmtnD24XJ2oMIxuNwuJf7nlumS0IHRc3Zphsxmfoh5Gx/V9f4YEvy1QXK
C7i6l8IzLzSwCeUJ/kpBFNgRghNIdz5nDpk9QBGsnkgZ8m3bKP2+90O0+8S+Q7i1
XRvkfzl0mYMjUn2n5maVtk7O2oFZTs7LE2IOJqVOt5iYB7BLmgfxdR04ypJvW4ZX
B7fhMyIf6899rGm1E3gi66hKWqgYEIo31DSy4zwAvQe1MqNCmPn0XnBnyFYGhGl4
4FtrrgRDHY5sXsSdYkujllGAoI2+2zTK+o4Y8Xe9g/TYYSTcV+WIy8Lsnq+nAFGf
weJ4rlJPhAz2hhhntdjKM2q3zo7Fo0Czsrcek8FcmsF9IkBa8L5e7p9gdCFWguVC
8VNWSsUF56dpfZbHiDOpL1Zq71xtoMJk2iw6xsA9DghK6T++Abc1OpU94p8gsFog
C0lAo1Bs73wHkVFX6qBIlzRTK4S4fokc/4L3sKCGB18co8KNiKqXrImkTv174+gS
23qeopro/116DJ4Sjl0sVh8QtJhfHQ/jcwovcCfD2AZVLlFGWnZ9mLPqm8QuSD0u
QS1EnnILeYFH0QknmrshDuefn7REuHpjE5dhDX1gTJ11QA8N2Vy3+YvDVd5aFxC+
0blBKAaz1CyLspBizy5MDfVDyYdi5TzssGANCSkJ/+U+AjwfgaMQg22bSQ57cUtG
8bbjj3iNE1zqI9fKRhwtKajskfRMXZ6ZAC6h7JiT8Zx0XX/LfrDyEpUr8vv41Esd
KP8meZSmMb/uJ6Lq6/6qyqaMEMBidCiB8O8Mbs3LLQJu6d/0f/mHIZa9awkCZJOy
4a7Swt5fGnGkf9eB3Px7lQFOh0DtF1lGNO1q0slrSdvtJtP0Dv32UTzaqDqUfjbv
cG7bPpNpdRVCtVdZXbv8KSb6npCOP69vAt+el1mnMBESaFGScwHr58D59TG9t3fI
WSwKNIB7+xKW0bL5i6K8/3uRz5s7PgvvUVtViVuhYyVZAfY0brYEdSD4EsYWrU1t
k546oCmsNlchgHx6Y2tVABMSthGoLEwDGlGVd5XhqtHNPqw2aoOGCDmNp8VtXpVU
6klBGNvbm47H6C8fughouz7pkuvJ1C8shh/m+l8FYGVqoQTxG+3Ou31uPi74oB4K
LzRUVRDVH6T5z5dq+xfJ/uJfXaxCydXFXa5s1lpJkoyBxZ5Z71M/d/MrAuGMJT27
hgCZjfwdYCp1sEmqorJePs1NHzSGWyKrQAfUkbMIa8yVSm26sgBEioYU2Q2laTy+
knzmXrjNJookQhx7RMGVXWwT9Dx5dwZVS/eQ0m94gUcVMLDj7KPi3MJ3GNvhvrhr
J8E1WpueT3XkXPUda+waaEVJOPGd3Gvq1f25r00ycqBynjOX6oNJ+Xj9eLdiAf2h
gjNrCDiUuHtVU7PL4cIKFiwIdrIRgYO7Sr+/nAZaLgAcFztga93TwxBP7URLrwdZ
FHLqBh2B/97Xbdjh87j+7eWoKH+1HznebU3BUyRBF7Kg/SYILQ+BMYgZtMXmyz80
RcRHnQl9uHF6OBVswgd06/3WDstsysO2UV3W+nSa8Uvvd1WEbRicRWW7+j1LbkQO
nWco1pI3MnH0ZzEyO30/rRY8tcw3aXpjnXGJN8kBZ4fqIcLbs0eLYLsPnESweD2a
epthwRlS/GPVLw8+wFuL2roeocCbv9KfieSeYkMNlgI0sgQ34ZzSMHyKGOQpsbaf
a2U9ZaAQzbK9pXEMZRftg2cYx9ObsrUZ2l5w47Kqm7FlJj6rSzX2edP+GaRYLlI+
uSsm6NVhXc6EjiznLXx5fdQMymaVKVVgDTUEby7TzI4uEsX3CjcCaWXmRiQhxdhm
IDS0Ole2kUA5aqiW9z5xUhRDHrNWFAtKCHce7plQsdHlTks6SHrhN6Jr9ld/6ohV
ThapOBk1Q07lbBu79/dhgs7EDrMTmaDde7G/bJOLeLtYOn7LdFrOU1HPomcjzXqX
r2AqiDP64X26s8As06hhCST/nBzxjS/jqgoMLzgWH4uM0C0i3zaMyN5EQxO4culE
m+USDjFyXgNx6CNIPC3atdswaYPv+0/7z7Zn6lH1tbx3zQct0SWtCxz3UrPeh3fW
CwrCMUbpCN2DRcufADhrvYPGby//NiANhaMITGUxUtxgwUnyxLOmM3zfriJxOJ9r
brqWclQ1gPWxN00PEdBauxSz5qf3vuMjABXZgHmtyw5P4wuCBJOq0ds86L5yvU7J
WFQuJ2Y7tpUNCN5e5sXwdxAaHVOu8b/n8STG8t4Xxp/43b+maz1SQdy2w5IWHmrU
SpaNtIm/Ay5TFcYenmyLgFM276JB3a00E7uEeK/oKDPeVolzHhJuy9TwTkjqA1BI
g8ON/2nggJFv/6DmkNNY8SJRtt1HYsyzeq7LEICIQOzkjRn8/WpXOIQzXjcwIyb5
bIpqPyoeY8djVGnD+B5F0Q0ZWvExbTpYCydT4fY+FaIILYbWNq8YCodkj/wzFJiH
OUsP6wtJtVhhUWrIkD4y52I2zgqCxPRsQWdY4tZBwcsAlF94PO9yEbcS8Mgu63RC
cB7ID+M1iOYZ8fULm3DjqT3/yscMfHxrgK51Lv9v/8L/KpTRT/OTSXv91zkfRSCQ
rtELY0hK52CANceU8ftB9LIKZ+E21NLQ0bRd/WVdiTqHm7FCBeODbf6TxVPvbewH
B6bj/LeexsN2uzQSGDLBkJ+184/evyqYkw5WY4IwvBhdBb/+vALNR8YYrZBrN6ek
0B1vuLFs9UAxfuTPyQGdvO8rHZtLr/GwmCXqLLZTqPp5Y3KuoC4Wrge8z83DXoT+
Xtx3hEB4nHPjXktwiS2B0myw3VhYTvZXlQDLomq64uESkvV4RfQ6MxMbDSoi2pP7
l8/FcCCMFLEPrZjTkbrMQ6RPkdkpTel/LDvK2A01zR3HQjpl9UFbkdrIofJUJitL
rc59Ugvhj67ija/Kys6aapYUiRFBi8WjqKWioca6iifODTJz3TgOLZuyLQD6Oyxj
4uCHp8j8VoCmwLPxDi8LSWyoOMTzr8fumFhFWRUWI8XEfAoaMlNa2NkxRxdHwrzG
nhga5pgohZhYvOE5PkmZc2OcwPrrWTqeEGe4yaB4sKO7IuNrp5e3BAgp5TZNPBq0
xybQ8/eZ32WIjivMpzVDtmV5qtaPqd7Wsa2oCwZ8MGquTJqABvCiuvrU17ke99SU
ft4v3acOJg3QZgkiUyUzRXbRIGzSnFyPWryh1d1+KvoTdmjuiZVGjql/Fe+DA6NG
W332+OyFTsK88GOktUZsJi/WZlBV1JUxMtTP3DlCIEgE99xaBmD2nmbcMVUndgoz
M+xHV9a/Vnyh31rLPUSGFcnzFfZh4j8xYcl/6iEAh7ycBckOfYFCJZRSn0ROBhab
1scoGU+11W6+fnKKEhPi8eOPQH8B8w1+ZUTKAM+j2Y3Eo+jiCdGh+SZWfCcP/l0L
/F7UiGhnBxaFntLLVXCgG4mIQVzrL5bCLHH1jzqSv1cXX7BJdQZi6v4OPbIg/bEe
p11K3/YUm9Js7A7UT7wUUUr0gHpnfPYrmksdhm3AiqfljosPlQMkLhO+D3+dVoFK
QMYTCNykPVNFlojdT7NmyTSzwguAzFXzxTpXHvq9/dRrhe6ElUZodZEF4x79o5kE
dTNqrArWaXN5/J32YS9gUZaM5RZ5TeBm6LvcG0Bdv2dV2FqzLMq2oKT7SW/Xvea0
cXf5M6+TVK1mvTekIU3eTDbGAw9KcjR0yojX31vGDr/1S1vL/zh5tBlDk8uMBO5Z
YtKatdCxm6MPIhWgUMUb5Kjc6/fkAGQ9qGfyPNyskmJehblPCw4DOwXuu24u2/al
8CJuMi1LaU6g0NgnXJxl5ZyTgK7hIcmdfrSOGDCzm3v+vCn3N8mFwsd1upOuRVmC
kV67wMIn4x1DeXcLiTXJt/NYYbCmciMR8S708BVgPswy0MBkfrvUQoKkNlQvGNd0
lS73FMqvCewmYpV6s8msXCX5UbE+93HGIsqxNeyckwsQjQNF5nO4eLyFvAD0LbaD
yGWzCEnD0UsYWFpA0A2s7DSQFTDo++KqN7EmWSJX8tg9IP9DQlYWaPsXTUHbYXqB
7b46MI8ptnxLCSCclD05e+9oM2rtl/p664L2ipEKUxqgBEELJuLa1yKMBwnwrFCZ
sQEUo8r3KJ5nMo/MXKHIx4a57+6LFulsaKadv4HuqQivC/ntrCdV7lKZTt+PtTrK
P+w5EzOETE8kE+6czFjI7CLO1PAjIyQAo6Q7Zzqm5Pz/NGvctjvc/AGBpwK1VZGn
lRxHbji0RNHQhyeGA0pHwU9KLZ7BrCsBRPziMNJw4XPUAGRrX4Fdvc9jdefU2alP
JCjCvuGogk9yKQ3L4FUIOq7GVMMtq6qjFdw9RAR4uh85nlV+gqOJAtfawUUcFwED
iwBWG+Eb1ZHLB9xBJ3rBZmXZ1xp654gaVcszY/fqWiPCNCUFAyJ/KYThdWUaAtdh
zXSWNf001bmZ411Kqr2fqDG2L+i4hsU1q+IS5jgT7XhBEqqVR5R/R+S9f4rNE7GB
eB4ZADbu9FN8QcMcWeZY8JOdHoeVu7SXAZTggpWJVgEGvIoL5dQUTJeV+YWWmXUU
q+ysphSthlF2urOr/7/YqxmZIo8dwYfSITTE/KKuD/Y+j3FJfXCqeW3beWyiU+rZ
rPiMB3s1KngUMhqBsQrlDdPynN/LshEqHU4o8Dox01OCAVlfis3cMV9H4e4J6TMC
W9qSbjruxnWSKIx8jqa8z4LotOpXoXeG+WtV78AYD3XtBIirn6RE1xUlx9P3Hb58
9R6TnZUeB9mQE7Zvlkfleq+V3PltZ935kx84sc7BYDn74NSUYZ2m9La8QfaK1A4F
y4lCShNjFGmNEm/4Km1ql+6pdm/OlvbVdoNnNLy2eHRNkX3ZtV4Rrhulsz8Nq9Ti
DIgofdBHI7tB8ceFP/G0Ln1Lw8piGabahAaG+3S4z2hhPdGjY6jy1Z4RedR4L37K
18Ng70HRRFw02zbLtGOAU4Q9tcvzCZX/R2I8dvEouENYhoFKaWnXsJlzhcaI3LWr
XEMJbBw5NKHKyhqRH0Japc80Sp5UTn9NYVsqLbY2YX/lzPIhQRT6zJw9gtJWK4Z3
XqLhjsumtd2V/ky+Q82bsxCT4MpWQggtAwwx8UwINRf+sN9ZSQ3W4rJ3SLBSc450
BCllM5RlZQLhu14P6CoPODX1Ji7hZZH+1hG+KdB34YNyhXHUa+Lg1gX85LOc3IeC
/0eHxtoHXDXiN9S69SYACJeoKIOLkZ8nrJjQ4rJxiorIKdYeoQukDLl0cPAHMswB
r5JwAoUJUNt4GALrDJn2nwEJhi1PQbE07Q9p8NprdUvlcH/xhVmTDKmi+Fo53yp6
sta+8VL1dcb806AqSnn281pG7ZADo0G4kTrWYgoetRAsB1Rttp/yPU78rhOs9yX5
UjhnM3pGxV/IDQWHFHeL/mp/iFNTxyYliUl8dwyVru0gzuYKcShG/o51XeofDUPT
Av+qrsruAR0sfaI69ffZ4rurree4Jtb1AsJNAuS8dexcSDn+uuREiTsdYI9vu5kS
Rs0zlzeVCqKNIEFEilr6q+xjVy85U4G1lU4QAkU3GqZWVBEHeKilWF5ofnZoth5A
Tq29ONl4ZYGyZLk0Ht5B0phcNgDezvJnzXxf/j+ZABRW7nA+SwZyrdlUZAki3BfX
95YFo0WeLBteu5M92qmfEYNqTQ4XYwNLaLDofvz8owTiGNyqSoRs08afFY74rWCY
ccLAAeRjyAguoof5mjYUvl60u7CbPcBvlYISQk6tfOhH9yuGFrsJg1SSqreFN1pB
XxRTQHGfGjI6kYr/e0Y7t0U49s14h/z//rRRcVg8TLFscWae1JyPUE3FJHCDoC1b
gwcFDrhp+1d0JMe/pBHJTX+HrWVKgG/wvY28QJ2yWhAe53Dl7x80qTLB7r5Uwob5
ZH8X3osrwHQqNPBlpMmKdJ4nCPOnvzViW/oZqzVbqyPsN/omoQ/zJOV4sjq2fauY
9sB/F1od6uTWd0gxxl4ivdpyuolEuoEN1pS6yfh+39tYJ1TRh6P1fk5i1rUFHS9A
XskJKNiiZ87n6oP5OzBRHzQy0pIH6vh/sc2+Tei8a5GxpcRes7+vmUJ0sexmMDSW
mdr+6YCndBSD8wKOn0lJW/b9fZdNzalP5ud3K/lrw8v4WeLPwnqrMmh9vv0qZvVp
vaykatIAorq5RQIscW1dmTRosxjsyIbebWEcI23tILTVNuXdLoTE3GJ35x4umXq/
ZgH4eGFW79SwBI/f7+Pm+F3Zj6iI+zdIphoeUaHgCeYmSZMSvaQkr9lMI0IdHHZD
t9KYmckgqMlQsM34Ipq/q2RkKqovdQhCFhNcPeJajq+8Kd46FXHus0tYTCjqdpm/
o650OoE8J81pBbDINKp8IbABuDd8F9M0e59dozqv2+Ld6t0JtkbBKuZzdIKRA7Ke
xxM3aAFzZA0Yt7yHUvzZ//ve0qy9K1hNBcgaX8iyPjkoMToPlJwG3ZoMmibbR//D
4I0bh2DoG2xLLiaxIya6s6gbXCezkLVZuPnZgIR1EjljpvcKwIGV+cUtDLGRyjGt
t7PG+piDGvFDAYKb5XC1gX/ZUEGRrdbVLFbrW7a7aldUaQXMjhwTvTK54vCrQ7eQ
XWw9xaxOYCzHruLZS68FPpw3TC41CRjzTfLNsoDdEvWLzZ/e6G8bPDsutBb6O84y
2vLVId0AIuu1qMAWDbkqPvw/W2ksTf3Cc0xS1didJH2PzHEQYi8efYtxbB1KhoFL
kIcHWAaiSkdPta9dB5pr9kglQvbOs+OSpQ+n+6DfX0Eyih9pE3JIbSUZpDZmEd+u
/OlLWZ7+RK0jTgzi1sa4xzsCKRNg8IJzaoyC9sSAwLOnxKr6Y377AmRq8MSsiCmK
GkZ9fCyZ3erPvTBn25XJ0SeU6HlhArItqkokZ8uZCEwTiTqLiR2o9KTEYw7zY/eI
1MEw6gWi7fKnVsSF8Ra46bNKpLxpptUJDwJvXEkAaIsRclc4MhwrDWS4AU3IeJRF
ARDwUZGp77ajYwM8uVS6QTJ3gpc35WeFLNWNpy/siEAsUqAjIWULmF5xSqie3pC9
UPotMWiojTUb8+GFT/JzUdY0nx0pvb1gYykPA1WuH3got/wDGKnB7kxLmjk8IfLP
IclBYs+Umo5B6UwE97R5figQZ+hq/cmJPwxCDox39Fl+VqxUhb+Mf4v1Nmv3JFO0
7PFrgnPNpD2LCI3LPQvqw1NYCFq0P9xS8age19q4u5hYBclHJIPgRz/W7O24r2DF
ifsbKJPVPGKIcArn1w66/JKeOvOPdL9IAvWHz1nUW718mVon7Z3EHy6BwXmcaBmR
bBbhrRsSyf5WxVBPmT1CxFgfX5BLhUhN8gCmNktxvqbkuXqVs4V2CWFCzNUcY+ER
WW+QH7G9pJqAyLNy+aVgrkp5PuG285zXJ/bEjrIe+8FInxWzc5e0vZplqXcyymNL
UT5xM8TKu/gJLA1DI7wWKB5GAThBrd6RVeltFQkGpTBLL/qAI9xF8mH0fqkzf8eH
WlfLLD/htOer6iUeZxgdZ5EOJaEctiLgLFbRMCbPQ5C2cxBjvaRAE/mupvk9LpqG
/SVfCQiv2rIsnencavF5IQBcTSu3Ib/hXNtc1IhZFz/lpeNBOnExiwuHxCIKiSyE
pGuviurAfzLRiSzpJ4rD0eKe3vyXFtAkMDd+EuaXsUgCYjSLDyi5BQpB5My/zSFB
RR25VImHQc1oJA3a+E8E9S6DKFGvSKWxNs6adp5Okdho8EpFhmZQaIK4FAPuCUya
prUC9GAIJtOUlzRtYYojIGRDU6HUvhIZEPJi5J8r5CTRQmFwsq78t905n9Yu4T9t
fS2oskHsu5cEgvrTXE5+eX1OQCAHLOg8PPu90TAw3uVldvQbilwiOBvUKydoSJJs
SmndvtIXf/8IZxQqDWNR+EpikoZv1hNOMfOwXIPQ5kNfTlBhR6yXnEW0X0B06xtt
JMv/g+yEfdsaZ1ElLzk72U5AJ6MfyeV0Y6HkqpxgpZOfive6VIjygyVMjmkEQcc3
GjxM2wrpQ4UhVg1s3Bho0UL78nCDZhcRXfnaWmzwxJ0S5JVzTPirF30ydAoOIGPs
SWAU6EuGEDyWYqTkLE3XEwy/XhTQLULUSMKxLCe0CmSJQfjY+XMADYyYgfB3uGlf
bkSc6UKMJTSLWMkFAByd1dZThRH2/AO2yW0FLgftVUfVxb1eI0z9pKm85VM6rIRt
eBktp4hJIXnxs9PkzpOco3x+uw/KrdqDs4cB7yc2ykoEYDc1EobvT65B3Q1V1hxU
WCe0VKjwwNJjKhwEXuZd5WmWhRzWRQfktWRRo+pGBp0vYhS1PGbIgCMT21LcPMj4
H6I4YR8rMC7DRS00xGHovpK8TZOEB80hXPz5CT2hjsiPQSZxDKEwKGGo74WZ3fzQ
TNCzLX+fwzKFKTFKNEgY2UkQnG8ToHbBJq82RAi7h/ZgmNymG8hZ9ze1PCw63KD/
e28GsOgOBZfDWGjTBq72pTNhPJ8elRqt4tI60jTcG0gEfR5lUWTimLCB1AtyyTAA
m+m5pxpkr68L5HNacstTKwkkiyqMjAZomUndJt7cgc125emQ70oXBC6U25zbv7Pg
Lrd9q9VuDM2qJPc4w7lmlbjCU0B+1iBqtbowRa1nIZQEbtLaH/5PzYdPaJZP61m0
LVmqGGkVqCaVR1s+vGb2YMvGZWim3VnelCvxESYWkT7tPcH1IZl8n/+FUzXXE/Cy
ji9RbFBgnkd/jwJkYCTe3yY9Nf27dYkKqDKuTMX/0y4+8YvGvx6o14UGPH8MJTNs
/me/KsTqsGmKpd7Sz7BSFvl+G/51iMuvDFObs2WgoNcAylDSrAioOaKCdhr8TCws
RoAfur2O9UdhKAMmue4ZU/RLF6ImbGezOtbYqtO8Hgg3bo8VmPj4H2XSmiyD23kn
pIiP/gFO8yQRp4k6dYmeQTWwEJI2kYjQHPzqZrN2PMYHKF01GfA9KWP917y62C5G
tEzrdWXufZ5F+SFl4N0b9FUeSc2GCC4VVmkDZ0wUsO10+KDFcwLG6lq6xH7vqFOS
4Mv8hASzftVrtkBkElRgr0d4tBmOujc+trl32+MIDpqJsfrMKSoY8MFgQzVuPw/N
swspi1Hr6d8caqgJwSRzAOYosdpYMmWy4w4br+1RWWzpae7mGE/h57hG3P4p4qDm
jFRtF669Uzv8ilvPXxJa98IBq43dCAtgtsqothYTuFZiYarttmd4o/T7s6lbolAz
cc+X8GkbyBZiMruPZtc48zkGVsgr2zjTZMn+ms5VvIhYH5affoJCSHzD9uEriXKK
gXral8wjBWvCB8IUCuhuTiAwd7Nrv/9lNv0YvF5yyCY/BhuS6pu7MJQpXpXMnJG2
zYMzRqDjdI72N4KthwyqMsdNAwg5Gz2UNTfyKkIYZKmAx49WwzL7RxKjq8Vr7yoe
S65kv06yTrfV4XeFYVmxNdmO29MVByfG2eC/5DJvAGPEwN0ebAa3UMlBk76r4VE2
bV2Didl9ipd/CiFstjbI4R1uN+3nBPePtISGidkSzFC22jOXt+DlkgU7x+EXZtDC
hcpLPN6xYg1lLcLEcNdHvbpCOmcMc+Mt3XtaBJEaQTbQjeFihDW0QizEo+Se1nZU
V3RpcGa3p+x+6AiXcKAeczeZ0Jm1+Xq0YFZhBcdFA5BioQn1DDbCRPl1x9e4lgMw
FE3xiU+9CC80S7ySfFYXrrHUdolOXqTqZn5rexZ6q78TPJQ42zkXhUiXTlLpVXJI
vWAGDvkRrpTcIs8/R3uEijjnCuqjNMiCt4HQgbdLOsWz4RA9x5Qr6r5ZFObgXW2r
bQcsD/deG64YElwZitK0Qjk8z68y5pblPtaR8Mg0HpHYkBq0BX3lI5GS9OTs3s5d
gSphkwmOMFwgTuT5tLIXyqJubANlyh0SVz0HsZB/pwWwCmUhF6YBQdqrIxEC7sBt
azH4Lk4cvfx7dcx9bQ9/t4QwgLq0eAPjl7e7JecB+lnKFfX62VwY83jIB83qwOJx
lpGg2nZ5eiBJPcv1sdjhB+GQbaDmAgew1afqkcd7W3ka/IDK7VBdQmJXJsThb3An
9cxaeJzZ97w3gPUrhYKmKxV5b0tmX1o6kAw9ORpIFNl/cmdXnDcooP/q2mDF6SHB
5060Ru7yq5KX+6mmiBKQDm+u4b0d/RUcyX2FJwYYBm9nYWn+Ygj2pTWioZPG5Qfm
6TzvYgFceFw2GuMffcxuNseMA9FdNgUYsP5Bhs4kDiDzqB2T3tFQVZ7DqZNn/OE4
4gfwijzKpphM99btIJpxT5kXPC/S3XZvumCuL3AWIwlQD6QhFtrj+4AQRh8qE0UW
/a2sUXpRP0UMqWP5GnzTA7Iw3kxsn0+O3PqhcN5CNqn8K6/CpZuCDiOWRiLswSEs
R6F0s5nMtNdnUv0aLAyNS8XO+g/U2TDhUgis01Q19QV3qCQyQBqL8AKVci5T/MGD
Bd7LmYzGoX7r9Qr0T8cc+t06DmYXGgon4PsVvHWNrWAQhj8PTa/PAvKaxZL84Tso
3MpYffML+pv+iqo0Zs6nMAPQwo27yUzTNxueXTDVJjVujbvgjWYOjK3Bn7dFHz1d
xEryzO9mzMneqjgoReU8tCY4+8JtRdzXBis0U9xh8zW8J2ybrC4sT4n/sDzz5aEC
LZxWFfJL0WvjDVaM8afEOl+fsuoOJvpSGjykI7XPkOLlQuWd2JICREzAVdjGNogy
sKOmDI+dqoevOjHH64SnXpqwNKVFsNQ3hQVudNzwRRKCOQrH2LFuz271iNnEBz0G
pBqLU8sWztX/sABg3bDidhnV+sFDf51OspdDwXVl87KcKiTmNH+SCo9465uS6JYA
tUpNeIE06qGNBJmRlCJucozBIxI//ztuMdVzBNu1kxXOdiOkPBzfoPtWl0sSc9gi
Kfnn/DmzpPvGt6cpTl0Mfctkj68ir6bR2ANwIwWzbnLtRTAc59+mPcOElNETCCVt
1Ok74gx/toygDrxtvCs7gWMzxYBzBfb2ANY6ZbOR8DnYMHU7GnUC56s1NozG68Py
G4qwwtkj8YS8LInPBB14CUMpOcZDtdGkFf1dCIc3sqSokiapEtYY9s0ELEtoabSP
Ec3nPmwAmYcdxEELjrr5aVezfwnlUyK5wmtBLMF263pw2nG3PSnChoPjeKwhAH5b
fPNloJ/9Rr2pOxF5p85ZypiODVYOFKBHTVKclvBtZGx8RP5GR7jAScQI3w/fjlOx
VyXZfbzolVXNTRQtLjid6Jy1TyJiXCSVxJ0NdPVgAgEvajh4AU8fHuXMol83A3gm
9mQJ3pCfnaBoIjv6eu08ubRcBZVJQlAV/Mcj1DGLuYePJkxeVUL8Vxviqati/03x
HRUmiah0pv3hSj+ITsvW3GQO4V/pJX9BQPpN4CYqlpABc7rlThUF2//C2GgpDDIq
zPBUi7qGMyxejIbyksOVe5WmUheJa8YflsWN1Ti1hotYT7DenWtVk2f6IWvhAhGE
YmAo7NleMNElHKOECy1/vH7ZVqtVWvrAh2/9QdyZAQvRJ8QQogMeuJ+qp1j5ufSj
Xd4MLAYxSdKp5XWYpj+ENC0vSFWz13blFhd4WodJrYkRpd2igDgeZianOSG4IbXK
UsCbpH8v8enibep1beG+iW+IuXImGKYxTIryqBhLyhx7EPGO/e4rMMbaah/s3V1A
vEz4Flf1pwWkLRg21aPyPRLLmfGtR7pXJs8YdE7FB5nYqQd8+fAksmDHUCW0wMPO
WMN2PEc4ApGUf5fs4u24ApBnp1qMjtfb5OM3/UEGZt81FgrMFUmUcflW01T4nX66
TQBVDYzFkcRBW6ZcQ5bG1guF8fxjVL0eoyD5LP/N5VhrycqNKHqy9y80Q1myHOvw
CN97ycPUv4ADsxOzNQ6RXtUCvgHEh8px65cj9hFTEzyBGZj+rAGmzC0z+GrdY9yB
1RBCN7EKwHkdA1w4EVWyB/3JSzazT7tVLXlK3U0+VfSMGOA8JhHsyCxwSs6kNZ/D
5eWyFQle7CrWD7hrbn42I5CdrmA40QN8CVbovUz2cSFE2/XZrhb+R3Io3AM2ux7i
J+STxmIghdFQG5SF5sWYt0wWvi0J7Lmq4D+46jMUfCxUIfV34TgO0C6aIqZJNlHO
OCuy6eK0PstS2mDE8L0BiPEZQLKIPsVy8T1aLG4dIMHGPaVtScDVVQ3WUhANhJH8
Axwi7uM0SL1NrMWAmYP1MkMKsp5+vksLjZnIzchrOnp8QRcC2POY0lDJ0DdU26S1
e3P9yZvgOjdwA1tMDI7+Qm9M722SH11shDjrd10ZNLgeP2bSy3AOJuypN5nW25yC
97FExYXXiPepIuw6fnmzmVfUlY8HiLSQaEYJ/VKTiUxjkgnIEYTyZVrXeTx6ss/c
LxYi1m26OsgbIVF0b+W8TM0Oj/BMc5jVYtKxm43qeY4HSAf5gLgwiTeVVs0p1UJs
kFFdZ4nZvxuy3BQTRPk+cGl6FB0hW60X/JdXG1+lbWO4IWv9ADmkplwDcugf/7Af
TMJmDnJKJI4KX/rZH2EHM4ssd8ntbDlZ27b7QLCruHO7qUv0PG0ANGMCY20X0EKQ
xb8mvqfEMy676iaF++X+x7KDSIb3H9aise6atnHGNw9Y8EXKCfXhul2SNcRYiTAr
P2eMbABl0aw4y/LVypYM1AvUKCdq2zlxOmYheNyi7b6dpZNhV+r1ywo3F3SWNLec
7invlcakkqflTVP1Px/RiuwfI5BswadidHhC9IZpwUWtCxwN61K9ZZT1WnlES1To
7G+H5eN6gWamcll4coycZy/Gv1aqdwY9N5Q23nNIJTCg/M2k0EvuMXsH1z3uIRSQ
qsaak268SItRJtth6fRfj+/Mi6M062p7XMc6VyApXUawnmkOch9ot5hH0IJfctvb
+Sjuj8whyedFdl2TTigPsQwSxFAr1w+nvjSO9Pxevu6T/NaK/j5P6pfuKAC0J8//
VxZs9J4bFua/ag4DD635xoWqAtwFFqVRRt5KV6c2HQxio2COwvvBWhEoXd93XbAY
gqL26OWGFWcfMxGBwSs+YfQf7Y64mDABs/fNH9gpidd3s0LO1QHwgRUNGpPCJb/q
VlZZ49EbAJMTTcSTA1V+MiZROfx/e7p0WcHCFx7XWjfSMHjJFKScMvOnZdRarBit
gnXqBqRoMqlxrWEt4Xv8aGgtf/ZHf4Vxs0EqrYHp9XK5zSIVqzUUQ3+JyylH9Odx
EaLeKttB/iWx46GY779DCLy5zLvKL7PNBNRSTM/dixWGbZ3eAqRSwYjI4Y9QCSFK
TJqXqgf9wcA8L00Ag3v4QINpyQ/rgB2kxCI+mmzel/BqqKcwiae9Av3U006hyxSy
7djD2mgM8qWLlh6oilzFKStTPGvmqMcUTK+yGYyNu+DSuDkl6RHl5ufTLm45/RN5
AxNmrVYH6528z8QiU5UGU+JIGyBNBlN0u58bCN5Soi4rW09tRtpi+OumsofqLfUc
mNqwj2G9LMcMt+SUMRUWPujukG6ksVnqFeLd2jrDyR8geyVTSIlHFal+HVAIzF7P
Ol1jjVecKCbgMQV643XnQ1uBUlT9elfDf2gbxDnkFkWHwOZ8N95IdN+gTtnPnR+r
WYKMbErLfIIa39PiKOkjwt7kLwWJO5fFCi8vzH6rcNK38IjOWzHXHgsgT7J5FtjS
seYfSjG5wcDwAEh+Bp4/ryuYcMiWO/Zgmx8Ngbpcfk6VgGBsme5hwyCYMNoWaQuE
iAJJ22kgMiNKvVRennUpwR/QVewzgZ9lGclIFRXVQJ6p60DZiS+W7o3CVmFkkp8u
ANJXk3nZuCJsIvzUZg5XwX/h+d/KOHyPEsIG4JE8LyV6OjnJ3vaFu0MhydmS/Uq7
ysl85w+dWYzKqv+d08QZy7lKBGS1dILGaHDn6UmpXkt3EYgRBf5iESRLqn7ELT5z
b6LDln1Hw4b4OfDT3eXXlOE53++NLZC+VFAubZ9pGfKqSJ+EYEErD6difGrz3Ct1
q2AHplOkDPBQ0m0f78UO8NTivFUWc0zYPssKVIkvbixlKHTc8bl+x0zoBcqPZDO7
J8PXFitW9PaH2sXuDiuHBgpsKsBgaZJyqDH9wW7LLyFDLRKH9nu67001fmV1hdwb
dnRQTHjY82PVFD1IkBZAKsfQEvpuhmmUKE3qjXK4fyd73Ogja3S4KzmwrNuWEmoO
Ix6QRn6Sc1dziCacSZvngy5KdYOd8nab0VhwoxuTMQiOBWHtDxD20YGI34zI0oT5
lo9evpSs+J0OCYY5Rvjeey8+cfPk/o+c8OVSXHGp/jXkin2A8jsde6fy97+bkRq+
EvLN7lmCoudHqFkvCy8uj0bj35oxroUKjFl/yEla5BIRkD1zIWiHbGIagkitVjYE
sL/YOEBAox6loESsFnAcPSGArsRlfky2j7Yf0qptu3jwDVftAtbGPj92P2lY6veB
PHjQfv9rL5TDizRzvKrEmKnzHrM8JTKF9j7Ybtv3Rfjk3/L5HUYGhJPEdaLi1YCc
3g48svy97IPXVTlG0wM05YIxmI359o40jnocle0DRm77ZU5KocMoEOlIrG0E4bTj
J+zR3j5wLSjxgwbZXkeFIj2oI3RMCWKtKI8fRNS1j0RbDyz6mYA8JxGxnyRRUZzR
uNpJ0PKPylE82DfHPXM/+UyqI2z98vZ52Vvb13rl7/7XtDmNs1M85Cx0+aJtbckM
PtkgvPJ9bXU9Q2hqFs+9e6BN5adxZ4XIxaN9kT9sx67HOOQIzkUx4A3FqYFkg6yM
y+laB3rDNSJ194SCi6yolPGDyCR8U3UeBhOowRD81uMvRgDvgdRvdbbPFAXrn8kK
4v3QsC/sV/CgDY3HmEO3Qk0SQrfiWR9KCuPktRd1Df++FnmJrDwz7U6iqm8Ab/cb
E2dcstjBoJ3/SLYrc+Itc5HmoEI2+PlFN7kipkBtjrgNMapDIKybgCMQhgAWTG3c
kb6eyl3Me9BJON79x9HU3bKlb4BbUAQVq/zjxSKiPlm64buqs9chZ5BzX+vzl3OR
AO0icueJUzflmQsxGCSkTgpDwOzZde6/1eL7sWLkeojpV38zAeooBRLSKozhlGrs
i3U4Q3jP/LSX2CI8zaUWeWQb1QPX4QzSOvXftuIYwEWmmf0kBM9yxTIBxrum/aBb
XZCtJU6AJ9Fqq277mzOQp8MM1TqiPCbCoSYCXXSPRdPwc+GsvRRuLlDzJpdw2yoB
NubAJH4MbO6IYT08dYhPIdyOLO1KywL/7pEWLw1+EHdBBHEFm9vKsKp7UfJTcPmz
DjLfFb2z4TE1dQt2lpydvCJRVgz/JM0xS/RmhH4sABqF1dwKAsbV+EI994AUp2t4
Q7C300ZPmLeFJinJT4rpbCKZ0tpDmbOEpbvrcWh3QFbw4br6nlXJhIcNQJqj++3R
/TBTa8Qk1eqsiSOH0RoF+a2vvVZv+IARIrWx9NNXNLbhtKC8Kft9O5uh5+gUNSNE
/n0Yfaa//ib2K7Za9aJx02Okcqr4a6c6r6A2VKwspzo72jgnNWgstECz43Cjtjff
XNWMxlkJrbVfuX+d64rXrqS/PplLyVXrHbp7FyclI1CcSEXspsyKD8dpO32ho2/+
HKHAcYZsObXMJDDiovfnZsyhC3H1QJrLlR+2FEqRZy9Bd25Wu9muaxvrjc+1G1Ww
kQaO4iOYXg/ILuUPpPXilfBqBnmr/ouo2wAHRZ8/OiO+t/smbQu3Ri91tk6SxAwu
9vKgztI+1Ew+y0UiMqTEROp5kPtoSP6y2RB2jpp1FNJmHcUkk7E6xFrBjffgTWk+
b8/+80niE/T5lxiI2CeIo9Vvvq5DNF3kDc/VbEHkEIafrhLUuWxK/Ry70hFH4sKd
qA/ksmTiIw1FIJ4xjvE6+Vf+hR95AlJKYFpbZn91BTcIfjd/mFuhygIj82BqUgOW
z8rlTHKuUHHFElPw+eLFYZtbhnKCmKPHm413ht8bkQSLulYasAIFP2xCMaaE/PCL
jSnMev5/k4TADUdVJ/8m6csDOqf8ZoJvbTw3ycc9BZc5J7suaMNyBIbgEZcHrJQd
R8sWgyTGgzQClLTcVtuCyMuHazzd4N+xbbjjJLAqvPdOYnHU5vSE6bJ+unnx6EnX
fOPbHkkTNNxRFkYtDaVoe+p6y7Py99lwB8Yt/C3kq3MPyECNRQZfAnGH4eYlcUrC
bUlBRNeEz+vwQSmy/U7UmMUXpu0W6uGWw70biqnSfhk6lyH4hoYsUpYCLvWlfVB4
/b1GzbK76i6dQllNLB5eo3jrak3e/qvcSX8/YRJIpRELae8Frk6jlFvdJ524BSSl
ILm8zJgR/1SYud2GoA6VDWWs5WoE7/asJVuioPw3StKtwczdVJM8FCeqNKosKQlg
5DhDVoGwZ/ZC9ekdwh9z0+VZ9cBdbbRVW0R6XBCnsgzfrWfuqUsHz57SplPUAeZW
7y1TyZwsRa1qrMFBNKnsKN0amcfzPG5SPsb/MlsjeeJqtrmLMvvE4OIJVe0bJRKd
6tcpaJbtRxriQ59bUOCTT6wkCX4UKPUz0fGuPGCxxiI3hE8pxlEj2RaR4g2UVOXU
cq0M/ALUbBuNyIal3QILxRULsm+ItAzPcv5v1V3DJfIj9Es01ZKGNLk/FL9mdi6g
2JX3EE3VfZ/KoholMuuOMcvnhlIuwQkVcTda9rpP017uu2G4OwPlhnLEiUUR5GGk
MiD+UQ17h2BLd+jCmQRyxlBBEa/MYxVH9BNYy1jJavHP7e6axTgBE5XPpI2jszTb
VBkBG806M+R1LQSCKojIVrrdSKVWj3v+1VwNWZ0KWe4ELxzCC2yiKCteTLztwjgO
YItCCOqT2vttYYu/aOf/3yyHOK/CNjYciQdYLXo5V0w2NgbPnWsZWnwgKcAKD40z
djFw7ax8WRGurmE7CVjGNOEmESZClX8IDslHC22p1QHKOMwfPiT//74ACUIcQIs0
Mdajocxf+RWAXfx3iHGVAHSnxcRtYHVFoEf4Delmc5/7pcd2HCBd/TG4M20H2ClY
FIz2ZzO+5OiBoDxch+4xFD5G/ThBzVHxwUEFlXPeAaPEIbRNAvTlOyHqVopwUyUl
k+s7dreae03Jt2iKENK7zV1rz4JZ9vu6HWCpqiKXAAdkly839xLB56B9YW95FjrU
vuvUNhXq6TdqCrsuQXgUfqAIjcd221GG8WyAYBDii5cCPlzvWCzEaITjjpfhm8Ls
r4h/LWQnlIXuV56JGewVFJxBNzVMTOeeGltJXToaZIejZKcTQGOhTdy+0qCIitO8
JHswEuwj6LIvi0lZtSm7ZU0ySb59hOx0t73H2x1gXAzQLG5aMt2o7F2oS5sUYCH4
nYC5FmGuJ84ZZg+0DsyU7qqRsdAJx/c5yuo45k392q1Mufc2G5min1eGpfqxqcKP
QTolMrEw2yUln+T+LBznjZV55LhdMfMttQNwjkb5FZ7/1NJ8+4/+4LISTv3PJXEi
USjEaA+4CJLTIxeR2jkps7+tUIdhXZkf9r+nTEKTYvVS1JcqCRgW3r0SxJdYJctT
SbNcPShUEg+V5mvWic50cu+RRdT7QIjEjg+lM/cOBDWn9spMG+2B4gffdEIFLh80
Sa/Cy3OHfYrYaZ3QTqY/5tGsZEhBtKOUKkSuRiPFuzPlOKNhlYTfb8m7E+0+GV9P
5W9bM2QYKVjDtQXWBns/Th2YEqa/MPRGkQhipsO9FkcCiIee4V0To4H8lUmFRqM+
nk8UgcuWpmn87SSo8QGJmYxaeVl0TBwXNnZZORuMT/sKeXPSzqaI5kd1trgNlaa+
BC4SZI8Q4OfeymHyLWNds9D2TE5E2320jH392tEPIwY/6DM0QlmsiYYAG6Vdjb3t
tfS1axn7qNdXMaRmZovd5i3t8KYgrOcRuGTcgscoFKBYxuloCJh6P2mrdP/JGnfe
TBPqc/ZVgoxAHolyu9KMKhg3EUYItNr2087sLSddeFhdvNg5aawE3HzykS/rbtys
Vg+lMfmFWJwGVhp5Yzw0ydWWta8SqpQSfc23jb10eNOYLR1wrdAWXcMEHAq43S1c
TS7U6vLA7JR/1CgUsdkLPMUSGVSMDsZzeCC9+u4opgQARnO8KH3/jVg48mBCdqUc
AHZnftHCku2pG2XDHc21B8e30ACYpINh+qOhOfzT5kZalOheicElvOEt/8L+8pjf
q7Wmmpjx131vBgiiCPiLfB4wKTyOco+VP3J/rrAN/nCEWDMmrQz2IICHhUzzGVk9
uei6og2pySL+UVQnxA7lyOJ+Re9dPwkpFW0jvl972l2gENI1wdwx236zct7gfBOw
ojVLgmlL0W+nFg5qUacWpxRAJbXNjnPosLJcHG01HveQUxid5FcXcaRBmO5wxEjy
kAKhHESzs9TdxFJsdHkg90+RVlgKbmuQns9DsXfzK9sdUlINEOOOucZEcb1jYA7+
FES0An8k6pcduzV6YwhnryTTxNocueDOPJfki/K/bWyyTSe0B3s+IZGFn4KJ3J9N
Tf+0HWxTDQHcRMqwOFe9Tvh7jIEI+fhmvxEbaEBp42rp7kD5gwwuf+UMrd2OEZKe
YJw7Ar+04QP/h1kEDmSVGHMj9NddDJlBUsDZ/M6J8manEjSt8cz3HsY4QVWyn7Ze
0+TNDEgHSP+yRt2wRnxs8NUZFlCJ8hqHRX4Ass1j6Pi7QEGmr4k6lxIfORFFRqMO
OM5mBgefBJPFmWtBFD8u1SAnLDp4qFvo1ejuLsLF0oCr2npDWdZ83L7eyDA4fhQo
P1+GQk9QAFyKrhfZ+3WsZwbPlvWXizVvWIOL6ZciNHUmcydcFtjzpe7x2jO8W6Jg
46ebFuhOuES4Bo9Fb9V75fYgy8Sd1tNJwWcKa2VR/qbXTmjaCBsxRsT1KiQqhWHZ
72ShsE6ZZmn6WrIT810HfT6/EzoqlBMxiemDtd+1fLhDCm37TQTQyl/57vDjoOiL
NfHNS1wC13unh6FFioR8UM2F/tdQskcEMFYISntBon8G1eyzLTy/O1QSpFVjCrCw
i17OU5pLEEiSTxV3lCzPbbK0KDchEt7dP3KN300W3e8di6/BUPcGunmni622yqDG
cUv4WQ8myjt5OFvMZ76OJJ9Dnp5rhz9sxTaNDnPTycM+EW5aQvIh3fK2WvZOgsOH
OgOa/lSjYB5ih8Gl2e7wEIWV9TrGhF3MQLhoAhOaDh6nVfeoC9VhelyHzYvJHXsq
6XkZFataY/DIqeoVx6W1pa7+YCaKNOM8r+sba/DtsVuTwhE/pQ7yz/Ax0hEMi9GZ
15l7qqbDq9cHDfP65gFKZrPZIl8VO1XnHNMaRhDBf8xYi6HI7yfWhQBXNyA5o7u6
GyNg0kxaKMxgnb8LtH54H8Bg+bJRYZvdG+bn8xa8AeeAOEuHw2V0t/BgaDFlqB/k
W01dAGPKOXnZlvNPTyToXdP0KHNZDqcnTPoZfHA+Jx9TIa8DdnLAupGjM1+uBH1z
A0vgSCMrEhjOnilQuN7w84qvZH+nfPB+/Ybt4D+a9NawCc9PN+dJI9d4Kzd9EGAG
7ZQmTKEsSJq4qek/0wpnqMxpie81wziWxQGn2G0CE6SAj1JVOseZi8fIvcbZDalZ
RMl0Y9irCqrpEif35Fx83ugB1fP4TFQxyRkPxNR9LE578bbgS5vPJbYFdh9Y93PE
MLB7TM111TAm0376L+kNqRc0Osz7659AD2fHW0OCKIS+ZfnkfOjVuhwfwPYF5tLZ
qAfyVqa2MOPf8fzUXs6ha10PzCI7MLFYRouaqNQxV1rafjcCKQ1gIzQk5wGs6HMB
wkCHOvnhrL6rNvT0BIjBf68Tvwqfg8yJPI/ii9q7hNwXqRCA5qdPLUuj94Rp3ZiN
eX4t8zJNsoW9AFc3Oi0CNv5j7skigpG/+zGGGZvlM2DUid8MYgf8o3KD3wEZCmV3
5lb+CSKElL8k1zMyEhpeakItFBzXxGcB2llKonGS6aJqc+QAHqvg8WUXRGGHFNGh
XBSUuT3GeOzaHrsOTeQY3uCSioet85je8XaDr6Xb8KOxRjrtVm4VqR23ARcZ7xwz
Qqt2lrEXPHxaO9k7Ios+O250vDCRPfnhpqR24EuZqjtCo+8yCA8NG7LX1G7w/i81
gbec4BtYXBfGpiEjC/M2J5ET1lDXuGTs6c1uVHetbaq2VQj8GpRCNAi6Ggj4ApYB
VGyV3dBWhxfqU/2r1vQJsf8zCuUuicCIsc5chbYyDtslzxHYBWSolqzTKRIabFwX
PIa78czuU3h/JPMRSLk4yUm3Gb7TcFsSQ7NMkXOaX7X7529Kfih0veRNxNLC6B5F
EJiD1BN6UW3u2EKqv90jCihvZ+goZrWq5LRlosOUrQv5oaxefXB8aA/smon35fpO
q7stNEQn7CMUWrUT9/m+bESHyDqt3+mCnTEi1MAUmxOUqYXNwyM6zD7EieIFFDaN
RdJIwnjRKYB6Qtyq4a8d67mZm5XG/1LmahdS3LfQhfDuZdLrTd17bZM8lqj6MH4W
OqMeOzykDJvOO9jnjhImnOoEgM1xVN8cPMri6YFxgKZI6AjKuZqJMssV23HGuuZX
iHcifvozzkVgdedvzRK1BnhAW8jJbN5d3bvLMekg9iyffwCduN5e4YKzyAmYaOOb
u2hUKEIdzZOAk0lgr7sqU9dM/8yRW6pTQ07cgmSHKp99Gg06TD25sc373M92EOkv
J2d/Rt1Byws8nXcUq9tMTdw2eP6e1GlYfIjZzOUEcI5FDpKmbv2ZvsCLgdiaFrWo
av0+AjdKmdHTdeuYxt/2cBC52OWMQbslrZBDJ8Om3nO9PSw+sFGFRnU4dF/O8St4
D90haWU2la5peZgaL4WaVT/r/m3eRj029EpMH3VJtJmaHSy9FkIO88kBw+PkdI+R
oOvEy68HdhM4bNrvtOhzhhStitD/2Rl8clCFMt1CPhdAG8h8FMhP8QkBuVzZnLQz
BBz19TcWESP6hRiQ9Tvepw2kXtej3GvCMU1JMT8SZePO6MEf2NF+dA7ZwfUeCNoh
6MCCnNn8v6vJcRZiXa/bbrPZKjHiqbbI9qP0ABrQriwCJRLMdNdrXxfMYfG1zSEz
Gicj3bmeV0BKZ4hNW7ak9iOv3vr7xmlkJM7RYldYOLStt2esUvsZLIRX5/CsPQ36
8EZjRJuLUNbU4G8lqunPlpT/NuVESqbdy7SeUyvzkpnxtJajNYnbZ/bK4scAZWYo
lVbJbEBvZMxl0kpkp3IO44JkSLB1wQkUOZ5jH/D7XkHiaKhjJnIrFfflFxhF1lid
rJ4GouV9TaOaWySv881E4xW/O4pbgR2QAm1y7HLGMAhb4IhEB3r1u9TMvVgdckwX
S+E4GdbC/QIABRGONdiOw3OJxcUHYPHY1gfa+spgLTpLDfhspNkNQo1GZM3QGOQt
RPXkA4IJA6ok5E9bVhOwZ65cIVnT00cvSlxDS/+JKWnTZWzrgfRiO9hN+tGsBYLe
gAS/Pxp5pSMyC1wLD+y0A+VCSMbM1wO5XmEPfmFj1g/ulOv6Xyl3VgR9k2ReDtp5
DxOFwFxRmA5LnOhUje9yRoudU0gRPwZM6KIkfWdLrza7zUeCdv8koFHxvs9uRGvX
pizg7kdtKZRTs8jHyn9MIp0TZiksq8APfEod0Oi9ySuCD/tLGR1nsZJ2Da/UBWOx
nRr7MbfGWcX8obtHt1fww2SOrHUmIqu1gqMk/IevkuD1fCghF84k5HfM+vH73Xkn
yYaAgBNEDPc0lc5E5PW92clOiHcK9aL3QNUzR7BCFBveIuXLx9dJOqdi1jZTPgVe
WOokwbnZgpYc66foES3aOI50+Hq7wBDaryMJghj4EU3vd1SkUjwFKreedXbWcAm2
h5mwt3WX/VRSVJw1QaiqHSsgyAKLPQG1gMnxV2zodc5iGUqm0M3/IL7z5sxMkeoE
eifpTKR9kab9IpktzE9ve1yhkriw5944J40gE44tsb3OTYuf5jSOa2yY3mAfwE1X
VMEj5Cff9hjD2ftluALK9/NY268GKnRp1/snwFtCqgILzizMK3+M/7mDn6QHVRZK
YGicdtsIwZ3nxo5ACzzu0/oYcqa9ZPf3ip6VnW1vn0xwY2ThHkhEJ5QFxeBvgiT2
NYI6JXe+rxnm25lVs5Wf0lgTiphIWbsRtX3Fm1t92sqtDHTzUyZFiVLdvqFf/kbo
eeLGWswvEwpBJTx/aZZ6UsW2zjHSv2xUNiqE6uyNelL6ADGJa47lCexU+vnGg0zk
LUWsx9JbHdcKGdq7gHsTChoHftF0P4y1rchZ3G1uttpVjuw0eP8aUQhbnrOUV/YN
1yjtfk/WeUF2Cfj7xjd4WYocnJ3CQ9muTSz0g9VfKEhy+I7rG73q2oUFmyD7ms+I
4BvBDgACSQkECY4X1MyAzONyas7FFnJKKEF7db1m8eYV1624+Iid5MQc2cJpRaQx
41NMf52p8UnGRREFxUJpRRarCFpPNHNr7IZDTian1vr7WbGsP+BuDCwNtznR225A
6xMmYpdcHekQ/aUo+oEZ37O7MKsusTF3UkQjhkk6Q2cU+ScGWTHJQpW2o3gdLAki
gpsH39lYY7x6+JrcPWpG1llRjq4DZX+uuKpgdMeyO8bu83RHkcvICdITCCbAzeNN
lRiyQ893sn/xeUJazlJG82bi8o6RTHIuuqrvZhNYZVkznRl4YMKVCJUx1zNjXasT
L3o9EtNFQXVx3MUlLUrXhc00A+cohntAd0dSg3JXKZU0Cy8zToBvjB7mHo54Gj/T
eFWHIhLJhKSqNo1wwSPnzorNgDH7AmzYDy8COrd2FwaH6LfmLbmDEwYuqg8tEKRW
mF9lcRYP6Zp5GGQ2BE9sBrHlTfmr16CMDDO+hij2d7BZM4kKvL7HRmwOY9LwGuns
z/35/B/OtKCeaBfAcwNCV3m2cdaJhULkZCvCIsPPPQIbC2kd58Q/hayWBRmYmHLG
GTu+pvjER+3B0Q+m/of9LAe+ZS+/DL0tExHoY4+aWe2CnAeA9NsVEYa+cd+RTvl3
mOMUDd6K977lb8TjCIfx+1IoQxrdWVpgPaLl7c8oucurqOt03KfLQXqLkpLpZfzr
hY32JgUwVqBlh2aVpK0nO6ljF/AAoH8Cpg8oafQpZcDUiuy1rZ8gfiUgAmYArjOs
d4/acT3pDentoOXu97ueE2BDuoVUAFUBktO0LcFqnwbtBEXYNYr+VmZnyU9YGXPt
RIlqOqHUBQa95g7BeE1bBQjeFuCWb8YNCpzIlWh349quXL8XAR91LDczRBAAkoJS
zJ7Azm5Ucx57ucj2b5HikNUiwFmI++x+ifUyAeUXdPhQ2lcgfxrZXphAV2ogKL0s
8Ir+k1qXmsVzPqPZznn3IIKptAebXCfXlw/kv7MnL2Wycb9ZnYmEP2Wn7gUgV4aL
2hxzCec7pRu+2NpERK1/e9Q2WMcXQnTNn3S4KEzgo5WL5cJJucNECfhNXXIZVf5N
bG9sWN5KYzuDQkeyDaap7E8aRiYx/tkd30KGHEPvOEAmjzq1//kOlb38LO+lahrZ
69Ka8EtcOO3rD9p2CBEN6dgk1kEjfKxI0HFyx/mWnmhGMzedUUAzggiIRmdLoDNO
Jc+fnPjcmtWcuaMU/F4svWlZ3b7HqmtXzrO30qXR5d8/0h1RXis7vUzTUZQHhBiX
H9KiSsp8JtUud9RjkMcdxvpkrhV/U3PCP6fO7xn7Zli2ywmMNQhkrtK6MTfa9Eqi
Xz6N+e9jP6hVXsumJ/ebxg3UWKUENM0f5+NtTscrrTpDlFrBIRqcrBQW7TmRybTX
JSYyIoR46FfpQBiASHeX4XOEiuYUoJzQ1/eEzg/gyzkF9gjpCaoLszivAPgi6uub
Xol4NuABVr/ZKIg+hlkDQtUgG4oaW0m+QurnZsMDt8PIP+Nb7yi2RHqrOBocZfUy
5qC2+p3J/r1LzyqlYlNAu2GtJKXHCnWiBXzz2O+ey/UljMcUzZseoAfu1a+1r0NI
mnqDVhl3xhiANnBNUSgs7U7HsGkEayWDgiI1ZPQMS1FSu6LaoIPCNWIJLjCnaHdV
ZARuZHgRuFyVl7ydstV5lo/rvwo9IWkriDe7cBgWzl1kXV3zo4oTD+tHbnkxrR9Y
eRme1iukzxPaMjDt86eb26xln8kMBD+DcgzE9vcb5gNET4yO4SORvCCJ97HJEqbu
04Gpiab19/t9R1u0+OjddtLJQhYWE1hgMIiOQSY5herkUyXYWD0+3JQHC1K0tGZM
rJHBr0GTiDF/dFefUNUd8L6gWpn6q3DYYM5RHdSzK/qydetmXCMevtoVgL0XRQv8
zlgQiMAAmeGvQfkHrLc/EFdFLlyS5p04RHlF6WemUMHW4YnuyI66+Q0KrzN0yMpc
gn2UUuschoq+kgLbcqDBvqE9ulgonRbbTpLQweZfDTY+jsOWUBvMM9ylpbNmYV8y
gDPBUAOszWB3nlUL2jPmMW2BOzghWs4HFM8bb57/ny68N3uFRX7Lf4z5xivBn25Y
o8xSQSlo26KpwjAYLQNWvNf4vFWKQh4cdRlo5ZIsS0b+qMOy3vdg06ZWEGGy+Mke
2PqlByWkSxUjXpaFqE+Qv31teWRoAbXcLPcS/B/SadLjtJuF7QgEp3xYgPdKwCbq
t8KyqlnFM5YiuqLIRtw0oGFVEi99jP+hsly960bg2mOnsanVIv76NuWlmeLkeGMj
iwNlUj1o+RpWl0C2thJBaBQQvxqf6TR/cGqea6xzxjiD/JHqk2nd0UgGafVTL6f8
ny96yxCTRLCreOKTYn6A9UBNcHeT0avNw1bRvjT5Hs+kUsnriDFlNzdZjpaVP8id
j3UGbDA8+RR2+ylFpN/x61UQeCTc9/Y+fiiqyEVUShpiZiWNJoyLOuFGHhvs8GIL
c5HN6ffFPwmIi+h//Seoh74wZ4sjXCIfifQcZFDv4BlwDi5/1a/EZkzOA/WYAd1U
9mfRsefT4BsWwmAwXcYxd6rhMM49GlVInxx8XuJOOtG/paFxzj89Jt8/0EnY8PgI
0pWTHdbaz5t3rIBN0TdY+CSnEqjYRXQdD/7tVN8b43FyGM8wbAExYJ+V/y9y+Nnq
IIg3XVtQGSYvG2cUFp7yDyozLDl5Bl8YLpu20B1CV4CxgDaU/H9HoBhE+vuz+zM3
X9nEsSnLdpwkZBfVCJpReorWc2QqlCpcuBIuXoGpNztd8m+SJGPtriYCjXMkAnPt
QwJmniGyZgz4spfCfsGRqCovfIp1KwiEVqbSupJpe/Xq/bhu/qBLSQ4nsVh2Q3iC
1I3xZEkxk3iWQv2G5YO9zgLlHdjm3K5jeZuYWdxfx0TON/nk5QVDTsX5KUM3Yc+T
1cvMXSkxTLPv1LFfz9t5frszkCd38T5LPWQsRODX7nvHrcBCJMB6pRi3fCfQ75Ky
ja2fqfyuj6eH62/r5IRW2K+xiGRqwawbMQ+QSeGdtT8HlKgmOxiPHH/PhQMH582h
SKz+Tt1YV5EFGjwUsBVz9nU3A6u9GM+vce/w5QP8xF1Fb8EHUcLRZg7Yzx7UMVVK
/nAo0Hn0+JdD476kJ2dT2V1suqkuQTxyaBLLWAV9ykc5Vt2tCmlQVa8B1aeLw/gd
fxSyaotxZkTK05x3Ehz/z7z2mYInqSTUZt8617o3KecFBim/lDJn4ZFHFUCLjMvB
iBhjN2R93g37uTKOCWBKBHGbmGGehV13rcnpdI8+OrdXjHUKBBV9f4LV+nZPHx+Q
QpQ3+A0nOcZZarVgkxnVDV1knQ1r7HoaB6vbHAWMgjsJPjb3XsDNaL/T2C/8zvvk
qJ6kYh9QL5V1zVFyzWZSk4funa9/ZZuj5woCtK3BMcHvbhRKPb6mWOPyH4m+merY
9wCmgHgDfnN6sSPk6XMZl1vjBxGWGonPv8OR2Eh+EoAeRrhVVA3OY3HxbbdHnlBR
rovsOT1/+axgbBKB2eNYJRViuqfDLubxOEie6hfme9YtFE5TRdUMZZzFHOTzU/k9
9dvut4yB9rNAOS9Vxg8riLD3zOaTECFIj1DOmGFQLDZZ9BuiNmvi7gtztwjwcow6
nESDGuSNQdwdweamCDjbBf7IK3B9AEIwXKaxqRwT6H20nRbaaSTxbLP5WCyaFnfP
JlEjJAodBfbNMgqNPK1FZVXYtTgyMjgA+P204rQtvphnDQUOLR/0+mbctACpFfn9
xQyWDj0+63S91gfUO6t8VAjzOd3OyX5MrtEbI6Yyv0L5l9WHQN/YAYS7qJ9grN2G
p7I9+AGFvclkI2Pr/WEEWkAivCvbpvYb5UjCP88CNZ+A7NBM+aLhyD+3FFElizeT
oKKE8Lz4/9aExLYlgKd1cMRIWreJrxwBzGLuJZCV3uD2GlPgqOA3M+tfemOFSOj3
xTWMXjaEPq7yx60a0s84b1XKUFbjHvMJF9v9c9nlT5z4LtOIENKBtgK6LBKBWS73
dQJAHvCUUktPvqRc4d4GdlsMkO9k36+rJ5fBF3pK3frYKUicO1agQFA6JxWUllb7
FX1dhgp57NzU0zmD0lsmUFxQKtah44N2z1ETmWFKr1eiSL0RLljgmAdaDIPXEleS
ovrw2uGHhThj5Ton11/xtcvu5qhjhhKz5zfL5TGusOzLKrBqcYIlx5uD7SRV++i9
sH7ZlralVMjFgUUHArJ7ZVXMAesu8xcSJV/PZabNZD3WjnEuHdurDUeFAdmDSgb/
DL9Qp9XNqwNmIkTh35rE0pJkwDIRjAHVuqF0+CWZhzyacGAUfjF4+wAZbrmB22QZ
8L1bxjtuP9eSJZGJ7XNLl1bg/dm5C0fBkM0Ws2VOOMx/vuw79K0pAQayyVOK1Waj
h66I/+e91ftRUByZ7rw1fIu3581loIdP1j/tb3zhw+SWN4nGRtaxcmuVJT6RVzNl
GMJ3xT0HfGC3BpiDi6zIRpPj4w8aPifoSybQqTtGjKozTnOsjq6bXEMsq3kjONF4
y7Z6TAz9kVNtXTkLGdbpAGubGuaaHy2drsAglf+lou1+i9VPabdyJefVWlAhsoQK
LNggzjYJgNIjOB+l+fLUiLXsK2THITUP3GuyaDV3WTwbVUldkHrCHyaZQS41cQmQ
/csGZVkGh67aGIHjime5kSgxZIETQIiQSNPo0vW2Xa/GCMTqNXCDs3QR+f9P3iIc
ea1g9cWPkYj2fnit0Ak0wAwOkLW4iGMaFj47NNvEnzHdXmfAcesIWCVqwbT2l4kv
jXb+q4bsfsm3IrdvKGRCFKQiyjYJQUIxtfGd91AX6GRi/9lG5u+rzPfNWlpKo5AW
DYd1rqLEoIHXixtOaM//aB5mjk7+kD6bSDXgjGApc+bi8q5cdXmNbhy0Z/ILlYtJ
KSINIf/ugY8TL6SkBRfhBPGW/C1RawCBdxaoW4ltwkjoJl+h2z6MXCSj/KiTIswc
cUYnpZzyVzd//ACA7m2vm3wF+60EzZQSqV+vL5xcaEDby31g1I3ebcBMXNdr37eQ
9XOnqGtUFtPHBgqRIib/lglIpLsYiKPXNXOHXM8YpsjtxG2wr7vegRztSskjwKLj
1rvD5ip476UzcnO8+gG9R3Bzhecz+BbX5+Ly+RgZGnmAmmFUYgFcjvSkCY33ksyX
zFIxTTNvUYDD6i1H9ys9Vzh90uGCjRX+SHStF9IfMZYqOVEDgUST9M91lzIqdSvR
jaafp/q9Pa1gMOqy3yHDwYtz33IcwCaheD6JlhQpfc+d64Nl/yL3OdAJS5+s6PSa
MkqtBVQKZYEAYM6Y2dSSIsxvjHNA2ttnY/32XJjeL3qbURtH2nyYUXMAo68eIDU3
+qURdBwoZHAre6uMVQZfOrenb3xQhSN5GSZVhBpWvImxRg0lgx1B0EBfWJzedzca
hlEiuuxJIz1AKZxqaGA2oVCW8mQHOXdzDY7vAtGDVsKFEaClqEX7sDVpgzAo/BY3
pDCO2kUqSM2Fe8iEUPcWoGgoizS2lpmX2QlC5dkwI3jumTwPuc8zfrQD/29z9tcj
AZnfsCjHkxRSUiqAzRCA03M5sonjRtBFggcIghDX2pn4+lFqomIAiRzSsOQNiKGx
dBuF/VVuuYRd7EtaAvr6c3c3RPEU3JJrhZlx9zTOmpBLvE6Yy0gJkav0iHC1Q2TX
Tx///1tFve/AfO95UVLMYxSkJFX1i1t8DwHk60+7Sp9IT7DIw8CPbMFla1RN3Iz/
163Tzwt7bHUcPf+mKD+VgXgsR5YVvbgLZ7WAT6chtSNRvOVBJ/JExzt09IlNsQ+d
sJrC+fu332QVCyRFhYvKuGjppH0AGxnjnTPjpmr5fdsQ7COtsW8dc2qtdGvXS1MF
dhhsddna4KCbDwfbgAMOs+nr9cbukdh9hOADyrWcITmyvkkfpuaHEdN6iEw1JzcP
UZN9Gtqjlh3TM6XnJwFfn865dv9xSP6OLpy55akIi66Mv8wWA6K91nSa6A42L6VE
8aaLFD5XinquiREpvB1opiFGliELgQDLl9qXgOUE7DGW5bbjxPYFbcgfsJrnfgQP
15cFTnM9Y95eV4fMwKSpPcd3upMVmxgFSaXKWXyfBirGPVSpg7JbFLOyCISYC687
MpTZ+E0Gr+7WZ0mkID1vj0WIkDfnrpVUCG6iyG7B0YByuz0sT3b5ZfNzhe+0oYUm
9FDU4sT538LF4xZopu+o/rZQMflAQRilE318D0LCrt/gZGyN4jq3ktq3nTQGdUVL
14mDF9ZGxcyLH//HusgyJPddgPWP1TNdg0e79lSjXVFAKUOFsx/r2Me9aQB+RoE8
uupZUOWaA4aMd8IhVI1yk0+5vWcMpquvKXs9dSgybo7K9jSMggvU1B0iBReTHYPw
/qlS1O6WQ62H9q+6AcKWdCFSJpa1Wm5sCgGJi8dY5PKItxt2BQMQohoVG+zI/Isk
59HASMiLkIWIo3MtBn1V1heQM4dM45iM/nKKDISYUKBKTwjc+MBY2+GYebT/s/Sb
VsBhHN6aJRMLmzzsw2pWwRJ4aRoI0GFCymEdcNPC9GqUA5jHJnsd68hjjMKtcnYm
KniNwGK0JYGRYFuFP+3Ty9k7WBtxEr7bGTsoLunQ/0HjQ4wuCWpXNQPUpKhBPkx+
QDMqanEpK2kcaGQI6e68cVUdivQxBgVCp49CFy9SX1/mIbB6+I5Le4duHwu7IduY
E7xqMRKksTzGAioqa2bqAfrGqQORxBpL8SkTxGX6TyXWgzKs2ttIfEEsWLNTZF/L
FzQfKKt8vKl7kMPQbwcjYEbwdIZFvqXL0x739CC+sY5q7gFtrAbaxsOKvbmuA5RV
AlKvRz4Hm3f3IKmwoDbNnTH6jddMIooX3UPuwZY1l/HIz6k05jPkyh8GuRge2URN
D5lb7uEq+wV+9H+rs3ExQU9Kjp2WxYwpWH3kbC/Q6lB30jcTZfnkQhmdfy10o0fT
+zMePCrlce3vOBtWhYyExt0Qyjs2Kk/QUXSKXMEoQ+IpeH+e4qb8QxDGds/w66P5
iby9b3YmuNkQhBZX9hEC9srU2CWRunJNKeIc/A5eZEOb/nWVM/doErT2kLt23b68
uRqWP6oga3ulaCi9ymwHLTxVtxTK1t3QAMyOxAIfLyk5PypGEBj9K/+sJHlZCIrp
TES1FX0dd0t8pufq7itMPjubfKfSTACVid4cBGDdRROMBEWYYYdfzMcfvYPsNxYP
lpYvYafQOwJOAflelLSgOwRHICw7JxLcqA7ovsPGaeRML0XeDcNyRXFEuYse+Su0
kLQRM5Mdul1VcQ9I/EiUJyn+MTthiY2pgdLHRxm7/FPwQkVkhpWg59ViJ2f0pR9S
TxTDNEPIELVZI6DyDL6wE5NPwClTQ4T4cmM2gactKO5gVeBzLzXf93U694IGGRaZ
A4sJKXGoyBfUwWrUfHHmbhv+wk0Qnflvo7jNE2ALB3LAmOpt0qIQD3hVye2g8Ydw
VP9mD+8J3SWPO3r1/FX2wztmpYPtMlIm8jvJff4bGG8l03xb8d/wTD+9+c9HNX70
xRPu8pzO4os8al4YAt+TZawhylRH0AgryAZ2CfcdMDkf0+8TXY/TCBjgwUq5zhs2
yX+0eOS2DViqv1npkTNlbKZmRxAkeSoYSuI+V9CqQcVGipS3OOrsVE8O2cyGYnK5
l+FlTifcwOpGg9eGmTU0zg7Q6GovEHWcWsWB5UygrbFujIRR2pnTuyw7Bechjw/I
sHjK0IJOH6umpE57iZZgd4ZLmdbQvSWq/KLJlcQEzxQ4MnaySRT68y7hmor9OuDp
vEjm9w2Grg1kSaZ2DcOCa1XtrnB7oTbgWNFJTO8nM8mTiV3MTbGHK+q3RSPEoPgh
JOfEMcrLT8IrvEdAJFTehn6P5Vflvhb3PKja/AsVBCOIU5XI/BARyCf/5EDe4dCG
9FalX3gk1H9fXUYGJTl7LMDt3+0Sp2PxjEkYPWLn71FxzJv/YjBXli/x4U5QF+Tc
dlG2WKORhhnJZABu0fTHkA+ePYv/X8zmCFoEZsoEUgYMTL0LkDsRH8mV8RBGC1TS
NNj26uYay0d0U4/DFCQP+XB3I7apKo9U6bbAWMvEnZervdnMZhadofIYHiqU/2Tr
SXJbj+vaM2skk27VexGLQ5WqztAEMDz/0FhqACLW7YEByeW67ZoLJo73uRYf1iid
GK75UrmV+7nQGj6TiNvJtBuDbBGE3H6y7BAF/jNlTP8uEr9XPthcsPiS3JVlK82z
dwz4TsMqdbXwnU0oyhfF8Ej2QJcHIJoeHHLFnI0dT8DDyaI/iUwe+4DSRCdkDQ+Z
oftFdUS6VoLxrHlxlYmlVGeqRPqOX3CKuX05AME4wIXCHiJW7u5mAeYQSstIzLjU
meamxBqi2zdQRGKEeZ2/hIapYJODaweJXukNyR1zFM1ZXF0v5UyY+6z32z/h9Y9U
0TD4UHLT4ZOKuVZ6zQ+iWBlHeYu8wuXXAo6fZUMA3H/4vugtmwX5tQniwG08DE6+
liu62DICJdz4SpkAXbJjO8gd0mxfB26yfj0QtjPSBgIEtvjGdoXBnccniSx2Wo7Q
xmMAJFXGox5r9YZVAqiFyr7AbYBUg75fGuSRYePiE10n6NzqnQuqOF5AjS9OAO/K
Uf13+lioiIllo1I+N9iQCIwC/6UTcnWnDX+r4kebXRoSZTRezCYn1ynVpfdi+dkS
a1qRkMnYFPd3yuWUQIjK6HnkZf6FQguolSQu0tP8Kqmf6tKZxQCygFBYUkXGWfEj
JxDoIoOmJWL8rtNFcrkonjPzLQJBioCgmEHDESjWOSAkqusMCK8dKaWY9ZcbCW1M
3Lx6AglZOk/PJDWvcF0CeFc1+FIROdt49OivQ4JuP4jef6bRNoQiHQ0LfsAfNKEu
uPf2/E/FlgpuMHF3e8OKcG0haH43X2QShx5uKDRYH7IZfEvi/K6QXT7SaYA3HYEW
7btHnWMxi4myQDpQJi6wheThBVxFPrzeoZXqn8EaKeci/WDKvUdCXCyfLhF4mZHH
AkXATrep9sjRGUBlwIQikHCUuvaEikIe5KYvCdy2kjZJ9Lsw6J2Lc5k6TP1Nhm1b
3UoRyhbMFqjBZa13mZ3EZmM4g/QWywQPUtQljdTLExd0OCftgNFJ18w4uZx7v9Bu
/nmiXOMLjCN3XjhC/LX9rIFnFZA1abyGTh2tm5d6fdqSNeGLioqH63R9fjYMoEkf
G9DByqo+werzWSarhRc2/cJQvua3Li7/OWBVdjmi1DkfRHlzqHGmfi565gLQTaUH
Xxd4QJqExPtZH8hCoExhGsGpZKQXthr/4cnDihO8m/6vvC24uRIXAeKBU66uqAFQ
V2VfnmOR2Po7kFoTUf+3UvoP+J9yhRN/PYyY6dsw9aSyqlEvbgZ1JsL6ZHKB9GWu
+28Q4GlAAU9r0i6p9IvcIB/ehl7uMYLXLAfFB608G9SQvaeThM0JMn5C8QuZUF+h
kVQSdiGzKiXE6O3x4at+UsOQhBO06NnFtHp3ocdNYuu+7LSPkTzE2KYBZCLDXILs
oF3JUqRtS++Xj22WrXMLunce8V6oQRNn7Jrjrd+Tcx38rxuYPy4TOvv31Rxs3OvU
iT8BPGUn6IuosvAtfqhaaThG8iTZmLjRzBkI0pJBdf022W8kQoCY/E1yhZuhhBmF
k30ncC5UT9ibv8Tqk546XWSrKPJ7wVqxuDbj/kPHt4RgRZJ26XrcQmm38ClPL0d1
lALTgSDxM62wEggA5JHLjFGg7CkaQBVTtxvbbasGsxxaKmDjLuJVw2n0eJE1UQmZ
KXEl18sirhLR9L/tMX9jmeRZfCKJBmV2cPz+rLrW+/cbbRGvQcJKsI8RESkp4mMJ
/ENdgyzVB7bKkrCjoh5nvnfUCih5GEDYdULYvza198RdN6mFprs7ZFBzXmIOhixC
0MKrhliFWw/x5Gp7N+2x9KeAbpsy+FD5bm68GVJ3J02muB0ox5ivDb3LR9hOpCFE
UYvH7On3BSaR+J5xmsq0t0Kg5gAdLGbha4l33K+jsPhTgTl9bkfh8urmLeolDAQ5
QhEkgglOGNqZLdpvSUFxE01aCE66j1Glpre4ziq3MkVfea1vfyj9qeCo4fVkRddx
8mApD6ZEfdf0ktzyPvkKxpCjX9tG3a7SzvjbAtU9B/UVeniy/f/Th2uyvfFdkXHQ
+E3W3F+xFF6CtFI4t/mRfgplMuOE9LEg6KG+MFBgaBuDc24sS4mfKOMG1XarW+bj
o18mE1MgD2BtrG7I3ky/ZuhjJ8c4DCdJlmxxOC/QgFiDbLwpbUCcpq5gRy1NU6Bo
hZnTdwpI5jkDbx0C19QrecKSv/peKwSjvfdMyMw3oYlxjqHzDuIP+q7ebE9MurFz
XQKIULQL9aBZ2JMoo/MSaRblm1Ib2PRjkfX3ez0M4m7ZG+dJa2kE91ShTfH7RNa5
e0oJ3epM9L5KfC4p0zj4aPnVqZXaYz+COd8VTNizvWxBlJGP/EnF2bJYuRe7Jj+r
rfun3BA4YqcYR/p45z+ddwifJM2aGbOd/6JCUHy3UFZbKVpmPQluUN/ZCCuI3JAm
7AcktZ8zJaj4iZQsbVWFkRdQzTZvpX1dILzMQtsWT+vi50RlPeU/0E1TuMJTmE7w
nNFS/Gv0OaGeHBIYt/dJX8b547HfxNuOod1PcRz0dx26NA3kxM5hD6e7VN8M7Nda
znWjq9x8h1UI2xucwhqa5T8JBweT+v0Pcp00WG/jiNcVxehp+8iGiEP3agndEeqG
/h26WpFZo5O+hfXCQHFMmRiX/TJ9zS8hYq2gkQ4llZHJc1lxc4TSQr964x0MO2qP
aG0avAZy9YVEdFjAkwz+YL0fssY2pi+a/DXdXYmdUbyQZzCuQWV2T2g1hbrJlIri
RlATXJPF7VuyDBo8p8TPOauzr8rtwedWJ5UmEBrpIEH1M0rGHqy+FJExyGdhDzAc
hgSiOBYbQZnuIFQTIPXLMviILqXEr9rAAWM+U/DM48T8+OQPPOsb/WH0pRfc3Jwp
odU3Zg31f1eBGoqJ3Sinl7e4I88OOS1FYGFqtqy5ZaFD4jx7l3nPNPMQT0cbusrf
TGDQauhcw6thLmrH3rnwP1uglipdKvKjHtzMXx5bOQNFASGYuI54Ds1reQGhQRCs
tihX55XadWiNJPwx7gOaOFHkcFafBZlTpZ/+biwqNycV97wwWidDNaDXILvGYnWk
GueXN41MuN6DGTlpuZWrb55rIDCPgwCCbYt8vKlBt24oqOMVDLpujm0D5UIvXKUm
cMuupflvUVviW1IBlwkOolqXFnFXFS7PrIWPJDwRjsOt9EJ5SRNH87w8IGakoG3M
8fN4y8Sma8fjfm55OCap6RiVHPZ1SmCsajeKiQzJAS3P/RYug/EB1dfHnJ25Edon
YSyvGieagPxGmeo4CfmG19R9LLUOO/HTNwuFQF98mOZPiGhE7ZI6NejUrNPD64pk
FIIZP7YQyZqCuN+S6xys8XZXjA37kCwvk3Ud82qjSH45vdfJt8y8/W8HDGb08j4M
R5AwZdUTlU/3uekoGlzrMFeJhwBYxvQihli0mEG/Hn0vJHWG15cHguyYU9b8L2DC
dz/vXqynrW8ubnAiqYEZe27nMrmWoXtxycLgq/Nk8k8Plz/J4uVf0b+gJZx++bDR
+NkMGZz4eMdIBIB1w4Puk+MXm4WoMuG0Y8HyKf38Zt9mLBsZjnzTfaV+wwN+6ucE
AfhAqJvzr30iyS6FTY0vhBJ2ke6Gs7oIjTYXMac3dIhufd/PecDrdKY/cNCMLzhF
wisZ3O7O/RjXGu5gmpI6RH7OGF11uMQ34HBH/5g7pU+mqfe5RuISAkalJoX5tFQw
i+W3qp63w/RUbHCyrtOevh9V9sLJO6+8m4Gq4liATfyDFFVXHA/ROJ75JCCb5ahz
rHg3LV3FOsMEbkhGv5c2r9HEE78dVRAesRsaOdteyqn0gwVbe/cE+WCtfbf1oLt2
Mt1mFAC5LSFFzGmq15JVZakmpSOoTdh4oC2UPn7N9Sbs4mgN2jula7LTiR5ROPF+
/mz43mprLCDFKCTfxpTCuVG8f+eVSLgA0BPKRl54auoS5fWy7q2nOdmro/M3bwR7
1W+PE2d2dzKAw07Cv1nKIRDXBrrbU+/Lf9icwKxMZ846P7/fMFLk+l4aFH5TmUFE
b7jq3k6xDe3yVXxLEmuSZdRn5q8oZdb0lD/M9kxKMJFnCtF9RXU/eIAJxh2KvC+t
veBoNAxOWt9adQQJO0ucK260DXINzNmBWAUeoDDl+EGSTlyxIpriaipgwty1jKf8
QQ69BzH2o4keeu1wDpkwsuUqR3xwealG23CPuC05Ut91FZnjRYXEhgYIodQkDera
bIPpJLUNUJcGC98TikMYiNXUs0qgVPZHg770tKTcYUEafaENL7MBptA9WYppvyQ6
WE3WrnXLGPGfvJrIGxVfbdK062tKRtQ1KORiLBTPrDAzdxIzwClRNLd1dJ60I/F6
+VL+fMaJlq3Daia8eLVbKY299wJUt6DJf8Wvs68yy4j2MzRSjOQR4gTWdZPZ55XM
NqD9LYf3IKhtZxjiQe1eiGX32ex0kpvt4NkNOj+BiAL4sSQGDvWo4L0DwJ9FaT9Y
/AyZpN/DFEyLlHypyMsWin21SPqSVpVmlmH5af0d+gEKM9ua2+cEapp+UYbRUhnl
vhUwYm2PS3LXss6FcX8sHglgy4HjYVfja1UNJ0jPP5nwYKv8bu2uoyNxff2NU72B
dHGxkFGrV8P3Nk8J5E/yu+UdXrIzP89oFbzS2oRou40QFPX1gOSWaZ9A2JZ4uY+R
bkQMFgUs8dkILl5zuhR7KC95B1lGHgaSF4EfcrADR0cIgpG2xnkFBRJQNEJtMcRR
uruTAxZa1IlEQq2MRHOIzsIyrl3Gx3pvC6ylyoIPs1Fh4QcNBESljgBf9c06DdpX
3qpgbh10WAY6L8X0rQRBbsA05zTXNSfYj0nxtu1z1MQLUwdyRZFzHjonxh4CLrtp
L1R/83QFa/kJ2aMuHvTIcNgE4dFR55r9mH6/pbbPqEkLCcRADsmAZBBu8RUsgEUF
0Eqhfp3lPzVB/ByO/xrRMyzS2NFKDw+qf2iKuxweGiWhmZK5Ro/oysjUUyMSmoSl
pw1B+0c4PBrXlCWtj8u/Z8bZzDbtbptw3CXa/jU6XcWEGVtjATU3KTT7OpWaerZg
tiwB9rzcCtsaUD6dnEOBeZE+SqAghH4HRNVRW5P5ToNQaMZ4mbS635LZxqxQeppn
/SW/dFEtgPBT1Ha/SBqnL42vsNN4ddxLinIlz0kzeaVkYPxcsrCOVJcRoz52gPZD
IIBX7OiLSWPphmFx/nrJOe8pvrWJK0cWd1TjLEAmyaHyoiKHiWt/RIetSyKIQs8E
kFwcby2+8l6RYpXVoymOdCShmNbNomziIOSkPPAV4R4gAzbooY/aHMgXLdRnS9+j
oYiQSS8YFBIvSDw6wzhHBDqbnXTYdz1zOX1nEQKbhR0H51TsCDLJPqCKxehoSo8c
4NepNEKdX2HGgyJIl6pEAXhH2KvS0SxsS2x9lNw9iNuM7HcCPrGZ5GHP7EvjLES6
5adJdeRg9nZBdKteAPATnzCuhhchAmgfmRHWFUgIrlIf2Quqfa48sE33pb4EueNS
sOahS6HlzS42aY5PPzHsW3BATeLnKMb/LP+Mm5+RgUpczzA+ZVngU9oMIBKd5Kka
Iy33dKi7opNZ7b2xW2RjYeJI+EC7/B3acR8uueUlhyvA7A1d5HIY4cRZFAcya08q
aWsT4Vx0q/lwqYTH3u/XjrPnpe6TwXsMSi9ihpdme1ELCLsBqHAj5ftFHHeSHqUR
kx7KAvpzI+wtDXIKm8F7uASe/Bm5pD3NPb+V2TcXzyf/8p8EUErobsc0+KVq5Nct
zx/lkRmILVV/9mXiGsCok7IJMGbWVrcXVfAogk6DmQPfprYMTHcpe8OoVoclwwFP
8hV5hEOO/xv1P8/fzhrlDTMdFIBTBIEcy/HGZf8NdBYkWcOrEpgKN+2kK/A+gHNE
lm93rja7wpB3mo3CnmXNCrfYDmRjSfa817ps2ZeDlHlZvnRA+kPvpfU1zDfa71t+
1/Hu9PjAyo4Cm3iOJkhLFhFAXyN6Oee3xcJ29PDD205TE4yNypXKVtIDBc7+sGCT
glJAWZof+zZtUFRwO+FQtUTuhZoV6/Q72FWKUT9nYyzqXB9Kb1orb7Koc3Wj9tpH
0mGxpvsPJZaFEYrUqidNBdH9/Nclo7I38i6cmV12eI7Vf3CL6ZDa3hn7B17OjrXn
L3en528yQkjEnUcVIzLiVojmEMw0YqfSW3xcMcB/JsotM51oT3ZU3HP8QuWebr7m
NAyVYJA8ilWcbsBWcfaeIuyrhti2tBvHskhuNFiG/itbBUXru388xMStz/JpA4ce
1/gynLJkjJM29pUrP8FaQG6ZduWakporGq6s1yQxrfLjAz0tzsmbYGSGXRzbMDJm
huxXUjgloP2zwJE6/nvI51baXKriCcQYULvYq+AhmnTX1vga2CrODS+jm/Hazq18
/IQM2XdKhh9rApoB76S7cmGCtuJhd98enwUwZdmmULR8Lf4RciPUEeS1MmtcxBov
1/Fc9WyQnJJJQUUXyNuI9wZcht9CvCXHYoW9vb98Cb8m5dMAo1e5NbdbAVrNE46A
cghxehpQPVttkgCcVy3uJioPSA15rn6DAWhOwoy4/10QakNKbIL/H1XYp7jNjkQ/
kReVF4Nv93keUsfcpaATehmK/iZUo8LUzsnFFbt3vIOd7nxVFJmwVaEk01qKptDn
fvpNOnFyuNArYUPeWgwE6mQU2VdFts1OyxcQi2idtA26JSJNxZU3ztIV1/YMQQCx
1PM7QrrN0ZmnGsD3YNNjGUVC0n7SXqn6WSzj9gWfr87P8vepkajLX9LM8WI3WNQi
5j1dq93iOP/FBAKpIonW/Vyhxolhf0y2Ue6cr1+wnHDfZAu9zzCZuOCqgbb0ZVbs
FK22996Ljl0WdO3A/06jfZ0zBDNhYH2LhOWIPfHvo35663wN3WWWpQDvH0xAw7ON
SXClCq3buT1MqqhZI1FHYokz4LEzxH0ARjXUbzLAnTwp/E93FHBXIZNJbpJ0nk+Y
XG5QZrrJhtY1dFk66ROkK5K0a9e7OeC9qGm4fadYTXHTOJAz0A3R01OA36OOBlzZ
7jHY8AWcqem4nioxE6Ct9I9qO/Gamm5os4uRYfR5idE49Ci8S2fI99UzfmDbNOk1
l1bL69txObvloLsorHqGU44WgjNjaNDrZX3Usfo+u7xqLgwWyyRwmN3o3uBRZREg
rY2vOT7M2Ns5P1jiXxvcQ0/KyxTStbCvueBTGwl4TkSnQlIE7OXgSBYfb68DTJm9
Oo43RMHAnJhb9cDFDr8ngFkjivtBMXeYRZ8dVhh85bGFHzInqqN4a3YwvzA4TK4j
/oX/wI6F3TEVshhbe2uv1xbYIOshBNKbnIp0vnqhfDUNOdvRBbHWQzclDCmJL/tY
HsAooozjo5JD9fznzPRMqx9Sa/GYcmgLoFTtica6LIbUPsfBtMcLHYci8by2BdX3
KSXIqNmpsm3/te8IJcuJtOV5WGNMSgGf9bhlwwx2Rj1ittweCVfUdA88q9iU+EOt
t0gRzhRuRwlc+qb4MVt2Dm8nJ8wIgIAMwAYTw60OPF2cmDLCPjFnY/KfO8I1g9Ag
kIuP8QBgmRW6NSALc0WN3JR1FwLwLLkTTSYBvnyqzNxeVDDjSUzBn3KXutcTDIUo
3HVLerigDBDkhe0YlW6GNZE5HMP3VMxF4g8z0HV3iqHSbhh5FZ1E+ooa5c7L2cf9
bPpMBnIU72QqH2y065xeg7/R3AlxZ3M98qfudLrOUI7KE/FoDrYv7bL5ibDsQMe+
YFzl21N592rQzY7XrX3fB/XmUB8FvnZbrYpxB+dOc2Cn9JzOPUdx0QtFN17fm82U
rFQLjolLtTFPQ4dEep7IE5/RDnupTF32tKnCSE/NeE1bKz48+3wluuDS+b8emgUb
FGD2wFEGxj9JhQd1ZBXEGB8sbllgUOimMoQeNelyy7oCcukFAzEErzgkcH67JbtG
Q8AwP4twslg4EOpMYiG2AKlaCF9J4Sm9hXBxkooKgBn4Lm4VQg56c0QVZNCjONYq
yX4qxJis7CVxkzSIRRgBCVMW5abX3cNm2ksSN84VMM7kErfe5qqDQK5W0a9jfwwd
5/HFTLKrBa+wHql9IwyOQPWHIxOsoZM+R6OrGfS7UkhWQeICEMoI6JhQyujwGJmy
wtGGNeakRa9ATywnhxpHxcE0ZmP9tJFc7/xITZ2A71DmZY+pz6doDaP05J5psaDi
uQh6MTriDdPm4DxzJz8pgN15WadVcFooTDFr77AJXCBD/1zHIEkOECn77jDxCJ/P
+gVZQhKFDJ6ahjY5EMoVNK8+NheDpwOM0ewzF+Df/JmEw22q4wlyWVbeBFc+70P+
cJFkn1ZSbGkJygWkOJdw2ZNaCNj8yUbr0VwstPsdRZFvpyBOW7L2rYU6E+NnPOUV
nb2TfYQ8zsQ6IJd25/twyBhsJX0plgtbWuMQGapgOFq9W/P8y9zNaRQtj+CuLCGb
gh8Y867WgqU0d8xRaLe65ZJjdXJzX89tfmsgbgw5csHoY6fhvPTVPNwTE7LbA6SH
fBKQ/Ecyh7u1QsT2cEwxoIxr6kXGmz1wl4zuoItLklJW0deg3o+L1PZKUI+Ziw5Z
fAq7f8EB5fVIx9d9fuK8eZvWsNnXKUCRNUyYNLdDgP+IxhZkNqLSOrDgEv3Zow5P
5uKy5mRSIP6B4f9dGH/B7KREocqR8ZXqQWagy1XtRlGRvn7lXq+5+YvZMMmJJnw0
U5rDFBwALwoKke4+yM1RBTewktlhj//U2UgIHXCfusvCmNVxTg/I8ps7jBrB22rK
DTkPsQFub9/VKYZDzAielrTxPzQ+IAgu+WqqHtGSAdIRPpybH0QXZ44pDOKBJ9jM
5sGnoc8rGHIgww8GY8fSDZecJItitIKPKFgQJ6R55aElrLaqxtg2g0+bWfQQ7/Z6
IEJwl4ioIVfSbkgXj7z8QGRLvoA4mOTzdR57AhP51P3jM3ydS+WFPs7ACt96UiAp
fcxPomp1GnZWKgMtQHsm/z8gdOFd6JTCAk5Od9XOkytogayjpXnkYc67SE4fGOGj
v3hx2NO2ZpayQQsaHddx4o99oaOcDlmfALe2jjyGZnmFugJYviYGohYcif7K8J0m
Sjd/JrSLv4HtbRbTxoVhzKldrUi1ynbSw58eeMrd4J/Doppd2fy7AnXYQdxr7tzJ
+BOn1tBcFv0gFIgioA0yMbs2ey0D0+3gnRAkkloO9hjX733wKBgNkJkCDtytTPYp
Qv9mnhLJugbt5kMH+i3Ey3U37xwbI1zhIO2czGzh2e8s3o+9/pQ1/0QP+gJ7JCM6
Jsbl++pVBJG+bq7gxb2kyD4l07BRPLVJYN5z1S40uhbD+dOpWsDXAy2FazXYNNcM
WyQtx/JnCA4zKiTploNZLLu8l6mMNS5suvpRci1uNvzZ8vExSvLybJpNjf2NJ3nS
JMGjcqRtG6zDbfIEXaplAT8bZFdjv6NrTveWuB3vrIODOmnslDg3YUg7kflZKYHC
xSRUEk9hyziw+o8NGMJdaB4zQ8tImHZUakEqiZjH6MunIGpleXQ704Gz/t29In12
Wkm0gNHTKnUPzFAqmXc8fosOMx0UZk5agEWi1GSulsB8x34CEH7Wb/S/DNXoEj1M
HF7CdhsHMeUsgXNmHe1bTMdNGM7q/oPWPwY2G2jWxE5WXC1m+zvNZn2CUEC9Sk71
svmUcG43JcpaPbbME9xa9U7smuRQtrnz3G4owqFRY5wX0m7ICZPe0Q715E+kG9LY
LWbiLT+c9w5Ga4rRTR+/GHG5Jnz5zg4DIIj2llo+2OqNpzIPspM0kQjrJe/b4Q2r
scKgaE2Vf+1uzDCYy19GIpgfEHuLS5/gxAPur8g2MUTgEeYfpcD4L1WO5xlI7ASK
ZKrlhNYziQsoP0+/1qs2Kdj0wtSkWog36sCTrqqwtOZLDNtc9rTBVFHDhtKBl/uI
e0M+GJfmahTs2UZsbcFK+a0isNTYPS5OoqmLUiCB7QY3foMq/BgsmSAVq/PbR/LO
y9mUxcNEyF4ezrfcoggRrQu8GH4wqCPM6HaC/Uhejy38rHt59HWvjXIzR388whe2
DJ5yq53d/uNfOnPQ9jRyZKYM7n/AQMLzla0LT8IXhOoB+7VrDB3jML9lhqv3lOms
V8U353DGwPHk3vx6UHYaS9gJsjhCzR+fu5aTKEWdoagKG4I5HmiMfRl/dDicDWCu
1lLjYbrhcP30UJU+8suPG9ln/mQRmv3cWn44XIZzO+z9Jxnuox04HaI1n5FZZ6KF
Abn3RLp6idNjlYVhuNF9FAd9zCiseOBnA3XgMmhACYkCKwOfp4nXWtokFYoZYPvA
tGg+QWRz2a53AIK6/t4mvYjkGuiH7uKbefnm3wDcQu8wM2cEkJpP/QWvQrFzJ7wJ
LNGoyuYyq9s8FghRLTuMFvzWxy5e2OvQ9SltzsYThkdOFIRPh2Wc7K6g55Vy1R9V
crFeM3N1vGWtTfSzRYgZ1sLKU9NWUe/8aOyqS1+t2388mvMtEk0WJx8B/cRtyHoS
4lPVxESvawGNo18VHbJi/3SzCl51k6aUx1AgJWXOWw69qxrfYGTS2PDOjtnZ8sON
Y5PotWOwDVNsaXvFlaUpG041MLXNt/lKg/jG5mL1+uaGTWCVAnYV53FF6bRhENX8
MSPBB6GSS1fy60q3lzrwZHw+ObxgqXJv8xLXkE3QO42ju+u5k6WU5VWDgeysMpnC
DhSL861ERtufzvGdfTCBwgg7XOG0pOdBmD7mKY1xg/Wwg6j6g2boorTEIzGBY2Do
OUHYBte4O0G4or4OR3/E3YZdwkWgMjYp6Wx5uKowT7w9M2bN2uPf5ILrZJVPFSAb
BYGzVlC1ZEyPazuJJcrh/JRJDfvvy+fWAgIfBAR9uobpFpi1Zi60Ivnwjzy+Wac1
YaJdkXriErn0UCrIJlM6wyAoThelR8hv6udnMmEnqzRoO0xAGUGwhW3VKRT6L3y/
+TZpDXE9YvQdDsj5fHAeaLfWK0qPQdX2XqB5/bKLZ+kJ2V/5YM+NyWFsxzCAs4iH
y6XCbwiYrLI0cTYseAoKv0e4bmdo+DqJftDkAGKo1FYFRAMgexLgfvKO0LCpBukN
zETKY+yVM/yHH7BFo6NBbAn9xQfr/TiI8yCiViomHGtUK9eKmYhHvuc8Ip9Qx4OG
6KTuCFnqZzg0Sk+/6frsa6curWl5dJqEB67ow6b5YLG5cXFAag0ucWqsQUyyQHAD
NeJbOMWCwVVDDsBzFCaZfQU60+EY0MGxcdSkmoHT4qaUC/1rjiIF1fv5CVyIjR9h
2HQoA9sUsyLlNQQ/YpS03nEDRPpFp6zFPDSt0EJTjdayKuiRh0hEsqrD6Ql5e8yr
rHb/nrB1tjHe4NG8SmDIvO2rviWcPCS4AoPnYj8ujIfUbqRzF2KWePbjNUf0F327
CbQU8Gb2mgzPteX6REMYNI8nYK0Knxg6fkiFJbnL07Sx9JqGvHp9XxN2IBLj7rid
diYNixE69Y5zsR15q6kgowhS445Pdzmo6iozQxMvD0MfGRvxeJvy/4gMOZtK9p5o
gv1oL+zy3y8h2zcIXOE8I0QVWWCAAFJCXJk5+ZVO6laED2H9hDKvRj9NZKvs2VNo
BAor4W6iuKs/W/AaYJfiyynDilnDOp7er+n90bePXkFhvf3FvwRfGh1uDmanZGz+
QwcAdd0RjRDGx3QUlupxP/+u+Yx0wLfEi1TaRbscy7HpyyHI2B+wv1W54iEQvi4z
/xiaHyPU9E1PuV3pBBTRZpTxh7+/3eHyNpdxqfIUQycB8u+Hk7Wyvir9+dZC7jVE
BqIE3o/ceRgn+3jE6d+j4R6Hyt8cUDkN+/0m13DynVIp4VW5Su5bzRNZCtfK+1TY
2Z7TWu6Na+8+QIjhLxl9B5+aQOl1WCjZEIh6QZQmc+shwoOtFwom+rfC3HVhivaH
UPuJCybve/GeSua81cnvaewy6QHTEhPBvjEsud9+HKNbLJUemDXRdZFn6dEboIvn
izZCe0tWTkPGOOQQ386GfGpahj29atTXGsUcGnpR7b35mwJlceUGSa39zX++cc6h
09n+CgBeuZyq6pWFvkrJZIqoY6L/+ZcsfDsmnUKFFu/gP5mF6uaJoMQHPN/Ygljd
YN6udB2UxGg22GUsdYowam02aIHT01S1WLAnRQ/CzUmJOEkYwfidBuNl3nx7K2FS
eVu1qxxf4Gn6A/Bf3qLfeGUDnfpdfuE6SNECNXMdkGkrT03HzMEDW+By6hSu3vvg
Fp/PQi9CJjGNho4QnlHKuKUYB90roYu4FGgHlIor7rQjoh9lNNgwBiv47PVcj7O3
mpKLD/EbRXOP1MfAbkuM/OgIzINw6AvZWYM0uTN010OhJb0imgd0Sx6FgU7HoLUI
t4iulClWJEN29YHMCCXvBnKJjl/Wat7m2FeJZJ0JKw5V2f6jDsIffvqRrGUa+bBE
uM66K4Azk1FXwNtJkNVJyLB4LLRqchw9SKnEMGZjhZ4s1GiGAaW5VyUBmEoiLnBW
wEB8iPZ1xHEDvgZDvnROP0EhHef5FH41gnWGj2xYpov3jmcfd+f9FU2Kkia2w6O7
9mKTTKy6BMHBIMra0sIH5AZUZ2TOYuf6hnaChFC4YF12EafF0yOkeGS9uSdNbKxH
ZlxtGC2KfKPmH3IxAdlNFOQJyU3dOCdlCFYBDuESI9I2R5N2oXSFBbmDcbyGrJw5
MBqRfstKj0kAbaP6lThlHlu1sPujkImoJxHTwBmdVG/Qrh2+SzGGcO0LqXqzZR+A
enYoWxPfAh7Jph9tfEWnEIuFGIY4OFLGg80o9uwfxvxjY3cbF9egITeVSeBDIw7y
XY+z/vAuv6//6MrJUEMWKHW9jqbkyu9Y8iUKukPTYVEFu3tYmndhT57ao+yxa1YR
82zNoyv9m/vso4snyGGf/avxk/cioI/MIKeZg8m45sHVjzzwbUlBHu5tNL7qdE5S
dg09rXG+0DTIlg1omIzqb9KUZcQkaCgh0Kt80BoHNwI0zNJGJhFH7alH3SZ3WdIJ
xrRLUD2MW32rpqM+PY+y8LgnOQHlJt1eRwSU+mWGln/erWHuKXDvWuIYChyhYFpA
APr39w8rpXtNK9OInxKN1WYc4tTKmBilRJcsnHp58tw5XS7+SddX7QYGY5pHnxxX
HIkjlgdQpYj150N0ws94pZKq+C9yBuuWq8ryeZVP4W1wMwWm7rBUHhUNxQxwKsgk
8gAZ1anxFaeTR5udi45933PkBq1DV0qu/y07DVUC+GlGGwSogx8uV6wED6bBC/2h
6w9iAvPMo4TUB7kxhmd6mu/WFWlTbtiDsdDwaTU57Q+Bsy3AWVer303ktc8qhfVA
6+bJW7AwV2l42MrBYFDH5wDEaTb57l7J7eQW5Hiw4ERd0WfgDYJBa4BbveJ5PIth
sjINm882MQcTn4m09i/NwgZ9PmAy7fovWx0IABX1I+Bb5CL7LzTPHmW28lik+qMD
KIERdYbChw62yNYTJzo+FDov+7NSzgXTofxCOIAMIanPNkDiXi86w2HsgrK2gltt
MmfK+1dRArNSb0CYIKVO8tIBFYfS0PekJYZnveUMjRII/3OjtEVZABPWu/7PZ8i8
6GnUabY9KRz158aJntCuBDwOy+lzyY6zskaI/cyqr80REVpo9SZfN9y/lN56RJMN
8notOcCMlRUqrsbU9xUw7rmteYaFeeTICrA8hYg/D7YDlDgZ0dUHgyZUUqeraSKr
fAm0y4kymnq3Q2vdrtx/y1eas35yzavGjFGh2UJbsGg4CRTiOB0Ol7ShTH2GTJeY
0pmM8ss2/obxkTL//THEZHQE/+MKGaj3tNg6pOH+ecut/rSs+XLlBkCyVnAj1zZs
P4+fhBoPsOkUprEHEzGjPvvjEWuk4WqXoiJuW6aG/Xm/c+kfkmePlcqi0/C4tjzv
CO1N0vvAIzuktwm7281ve4gK39PftZPlEvyXDnOwiszuroEuoXBJdmARybCtYcqt
Q82Jf9Fa9vIVU3KzLNrcsbJOWC+m5EMtWrtPdoTVDghB/i9UQIKY+D81Yp/qkau3
cbdH/n0xybWx2vUc8mML4KuN3UO5LafPfhWb7jW+ccWzoCv+SeYedl9i/sac3CyW
UodzPoNnZjJVNTGmpM/BVYSgXY/5krDtdRryOTr/KgxjpEMzYzNKQFYvit4a+UQ5
nYU1lHKuDl64Pvz0tIgQgnR53iYUq2/9urIgMab2elD2cqnCYPwrn4rOVEBOl4QU
lx4Udxlw26SgeWrJOvBB2273d2Fj2VbaJY/CeiapA9LYHd65vqW/6oIc1yRAN2Y+
Xk2wwWrRW+zpdnSUQS0uvoV15smE1wJi6if99OVfI4AuyDqW9Uv0VZNvVHVBz7z8
nrErB+JJwtLQSMWhctbn6RDBODANzOQVLWnkm7KYG4dtrHOMxUebwdlHNZBU00x9
t+ML5z54u+IZzUml9iranfQFAWJoFWudyPo95mrvzSys+w+QTDklHxRtcH5HrWAl
4w/vM9BltXXRk1bzx9hp6AKY1kHtw7D8dhmYgajPv7jfwGmIUELVP2cFb9De5Hm8
D8j5099ydrBa9LxBu9/Tr4nd2DKq9UWy/EQ2t0Ib2r/oe+YMCBkM5cDYiNU0yUse
g+kav8vXEXzpc+5h2PRzPAFCW9ci5y0u+YDUGUtY2GuRI6J6yR3D4+UFP3Oh6VUA
2/W6DbZmGvvTjMwMFyq9gLSO5x+hRYsqyc7XTRnm3pzqfJb7Sd7IokCt7XHXmFYt
V6Jf4GBUoiJPVvNLyGzD2ihsONzzxkZaorx5De0ZTTC5IuxjQtRCwe0jMPtuIkKb
p9N0BmkERnOb3TWwuOq9tsQv/2J9gsHG47iJBlhw/WQLKwFXTyPWLGNPCB2em3HH
kETkLGkUbTE3XKgu9IbtWkIxw9CT60WZozAfvYyV2jFhAV3gKDRH2g9R7vg/htqW
J2X95RngGpo7/xNoMkUnigtT58Ck0Wmp2OtXebHQ4QzG3sCycZ/N91Mo9pt/8a8R
T97JEE8uHuXPqmtU/QtX4Gm2fr3ntT9dGijY9amzERXnNkYuW3ElVyDKc3dqE5aS
/uLpra/EpD3Kq5nd2VQQjt24N+IjHzMdXzHN57zXYZvatlkVGRAM814OA7ORgqc1
iUV+zgbMC4fWZ5/o4fJuuwXPijFF88P7/yrDRUpaYYDedaGmMR1NjKRep/kkkko4
Had2EQqlqJwpAQI6eucOkGYyoOOhT4RmSe1kQOA/31eRhCz3NcyyPIGc9Bi65Nc9
EvT85JbsRCQvWIEllv3gIYIaEcOMXvKtapFgtzFZGrHUsQ9pKzpuxm1u4vW/gOTG
BmbUIb/52nB16BOYIyvUqrQRrPqYxIfLrJd98c/Sgr7xlPxXTu47ltGso7U8DnnF
Y+XoscTPOvsA09G0mlhpkfKjT/sAj2qC2I4bJtUjPW+cEwHHdkR9NiQQT/BqDwiP
xG4TpalB9piX9kuF2F1REkMhq9WhXptTsTGK4xoNvbNSqXOcx4BLswv70N8uo73h
L8W2YgrZKDWAvHslCuFBx1u1Vv7Q1vzzrUjzBoUeZaSXAIhF/Qr/womVX/6UiYoI
dj7ouxKKhxyVnZnB+Rlstgjyzm5p094EJNN7AQsbpxvOTeJU+Fg5ZS6sebe0Xwja
sTbjOxgI4U+XDXLHU6IBZmn11cTazXtc4GFr2zvFk71vVQk2aIXS+F77a8kIxoQJ
aSxFaOLXmub/tSv5tRObVcGCUlRPGfExYhgLAGBhrkcYELXnf1anJ0RV9WiPm8lZ
//ugDvTDmoPYOkUEmtorh7TgJHaThlvAF4Pz98uyyyvWX1OAyrMrq/PaDOu5l8lm
muim3Ud+v7mOZMilHfEbBasphRPMWG8ZQ6UFZ3/vfEk2nGQgbXcCUr0TGMUidzpm
5gyeciQZMOlf3LwQ2/5zuuUfFR19oIsScdMDtOur8dKsDaauDc2TWngEN/tbAxEo
x1M975wMn4CC/ANaX9qp4/tD6tiApQKw0DayorHBDQ9nlW091uDSRqV7GHOJmej1
S+7qcL11v7C7o27IoXXJVH/X/aeEdgXaAD/NKg0Zsz5ML/IIeeLpb+bLD8guPKBj
Npd1oZjGV+9PdhOCUWjqJoGv5mLWjZT1ArC/H28Ac79pinfdeT3WgcaSEJSikrIU
AGO4VbzCagwXSJg0xEGWn1+975I/9JJUGSwRZr8bRU1ZGBAKbkgdMCq4OvMlTywE
NRYRxFhatwZegO7RgC5N0LrbVbQWqJQ7OVYtJj6TGN/EKjPZxOpYdBCdu8M03mOu
6wLKMr90Jkegpc9ZIr0wICp9i7TRE6wlTyrSxyAqLmW4oSvI98+vXTioERR1Zoyc
4YqG0akWIEWurXTYZkDQq+UpWCAeH+2tHrZ2rRhsn5IVqA8+CWGjrvCeBrGkKhUg
XOcz4zeWBiWrtA3LzWQolxBkkcgiOpFKvjAN+NJYXxvdrzaO0r8tphnYv1GMMhlY
Ev3BvgNfahuXyCOvSk+Ag/mr1etwmFQEYMz9b+7IifGJ2y4zhnqzrUxs96jEyCfE
ow/iPprbhv/pyuo4bCHReTK+nBcgqVb0kSwMbvLHhUO5u5MYk1uVo3jZS6TWRV2P
SXGgQLsHIv17K2lFFf2U8ry9LcAwxMzsi5UoPohCxObiPMXqawOlKFpkFmHPm6gY
UO4AthDwcYFuPIQsMo9LTXgk5PIQk+EnHYyP+tLexbFYhhA2THqomSPpQmER93NR
b/Q7ww/pLuS62RCMdCa/AwIJmgvJvXIesStV4vbEURl0pUbUuuHKwJv+QreQP5wS
VI6/fvFYDiqga/fYUeh+NW2SGjKMlxA4pGVBGFy7NXgeMO0BYf7KbQIpk7ME7UV7
PhK2PB/jyL0n8AxE47mpXcUId+Fy35JyJPOKRTsnKAXTVHPmyYGokYAlz1R9zRib
p89LiRvzESaOCwPXGx9Ftlh6l4WhJPt4DxNEoRbNhwsufs4DsoEFz4ZZmrBlmaiG
Vu46r/9PdAelZgT8DnwNr3poSuxhEm6Agv2Uqcj3N3jxPwPRSWnGyt7sLh14lrnX
WQJmRdoxwQGGFUbZNVsXohDDZBLDdb0VdBA6EvWheE0czh6MIT14rDI0QAIO7SbL
ILqGIZcChnga+GSXdXt8KeChXK/l5N8oXEe/myQfJFEvpfajnrDe/sY3hWp3yP1u
31bVbbIJ+V1P2BpHDax+MDGwVxdECCfJeau4R0NVXZ42QJ5x3aSbw/qaARMAe/cV
LCaVYvgLtTrm42SA46rmeUblNNmi+dHDcklp/eWqS77pnm1igsRy65uRxmb+ANyZ
b0jduQ2bb5r41XCDGL0wUqcTlvq/6UNGBtReVfQkhxL9h+gzWhzzCrukK437zp/7
kk726Ajbt8iAltP8cSkOYlzCSkwL7yqExjTfYEQpL8iSH7lsprmSf2QYCL2OsNi0
/646Ek25pKFUm/RCWF1qhwoxxuRmXq/Xy1mmVe+AdA3hVEBiiVkqkC+VjLax7L72
madIZoY2lEI1hLvqGCKJ30criVRrAgkwbHehk0Of4hCWR7/v8lBt0rdSFdNgQGLO
BZP8cvemCNCFi9mm1cMVNv+/1FdmgAXnfipY+OcaWk4gc4l4n05Qry2zFLiXIBDP
bvSDmHBLbM/ft3qSXFBhIV+1Sg+Xkhsjm5c0ggFQsVrbsXJLcsSuCvnlG2uRSjh4
1QxWTIKcx6vmDyrXbg7Y16w+5eTgJQux6BscrO0tKpeqWEygXXwYkEp9MXsg3dL+
oUbnUgWbl2tDVDV6HQb7pAxzzwDAoAGASTN1ewzlphzivUcHVFrHjFSkrNUJFKeN
5l9IKJIPhzu3VtA2TIce5YelLR0BITWkYnebPxmaUdErNJwiqLhZ3dlyvhwmPEGt
FFe3HJYwMVC3YkRoMqlcbIiwMvkXhy4DGsFeeo21RXln9GSDDv1JtJ7lfrZsZtUy
JbZ0+Kji4YHH34XdVxvjv8Y/GZHLYj3rPE3TKcOiRK6DzapCMcNdjqkK42conW0x
0WJJBN/ZNoOBZYrOM2GCr3GwJm+aFQ2X6sAJ1RLu9xJoeeiba2MdlS1Ei8D2mTa/
owYyHVF14wkH9XSiAWD7MNyBQUf1hye/jNN1XsgTyvEWu9+5al6v1CC9ZR3HhWaE
NlEptZorKAHnuqlAdefETAXF0YpnYMHdur/TFK/lA8XKqNT7kU8xEE8298ueSJdD
fEGqyzYBvOkMi645j7DtSBibZx6SS6toPgNtslSfOII1yV3WKtkm2WStE+RgjVzz
pmfpaUKDn0HRooTrk23PosnKoe/1acJSAweEAgB15jtb3V9ARmaoCx0hBZ14MgOh
7LFP+89ebh/l8NK7YxfIxKcgdvyqJ/V/7ifF9O29FRd3R55UVXvbjRysm/uZqeWb
2scUonqT/Tpwh8gEpf8Xq8gwVUulc3o2RPOA/7EhWZ6aLiJnsyAdBybxKWRbQEvQ
87R2ClF7HQqkZxsGMsxOdSE5/x8yHh/pyGfCBbn9nAHHqXXI45umCSgq0Bxueh0O
zDKaCqcmz9c1AroeFBfYy4va1zK2Pbx+JirZsp36WdB9pz+mln1P0+nZ8PjBTXz4
nwsRYmFUGdB4m4DKkfX7VmvHa8uN2eEe6zlDgYnI6uZjvbZemF6tiMuECCZtE0pX
7ER2+ci0AUqpbBZ03lXzDasS0efqR7gif8fA41J15foqS1/RmdH3tLe2HR/4IQE1
RkTaNuVKn8vLD32cR6NQhNimjTyEkfv18yEFci3igbpiEMpjurQ5C1HACNy75mDZ
p4HnoXIK3Vvoyq5q67Ehr45wx74fepFaHuE77dkFxFhEiYRhRF6+hRHF/geEo1Xy
MftMFGz2DCtJE5lJEAr0Ok4263GgkfuZd+4PeLNFpaXEBVo3AQlFTibY4/nFW5TL
auReWKsS+tQAI+k/9sw++bL1LCnXmPh3V3PE5tYBhbIM9LBOdhE2U4JngYiOuV6e
y6jnVAsGQZbwYdJZGWH0yg5GtNwQnCjr5ljiQPE30EdR4JQguIpbgzjtIl159Ohs
LFhR14O5Z91DzIK1p0z4TvzgKJtTIUIDhe3WUdeTSMSIvoPKfe4chZwIbrPkBvU4
DSginsgoe/hv69Fjs6kcKZerGFZNVNU5z1bFl8Js1GHJ39GSPW9H1FRV9ctDWv2G
Fn2n1DJxroNZnssZCD3hvg8r8f/pj0TdqpN6xyRY8+kPUxUWA5exfiZlYoV2MLpl
ARlppKRDat7P1rwTwmkEjA3Sc0jKT3qr2IDOfG+rwqMBy/GU+fjxnusDZ+sBveb5
dED3Yi0x6s5/e9K7yVOLbypLaqYt1hnjLcYNf9GQh2ZVTSlA/pHuEFLlGD4tzBlj
FDSsKiBMvDcCeukcWomgvczBP7X8BTTqRSUHsayKN8+9JWYGaqwdbT/YYsLMYN4b
NBrodvs1STHzb90nsAq3a/M/P5xFwylfvb+l3EHZWF4qlv44zTiS2LrAG9NTm5BH
5OrmHc682GG4D83+1Jkr6N7ZMh0IO6apI9C+Clwksg2Nph6cHWGhy3Ff9tpnj4Ay
t0so/QZKUCyN0mHb7mpB7Qh6yro8O3h7c+oc2ni4qwUwcFS18Kn0bQeqLO60/oCY
/0eCGmaBQ37sR50fjeU8/BUgaIdnECeSkX5m1zC5FTy/DI35/9F+tOmzTG0BR4jR
KN1W+UOHccSIY5HgJTRVnrWDQl+QtPcJJkPBo9wt5Qv9plNNVfGauYkcA0viUPN4
Ifl6A92hOEnooDje95WiC5xJoUqAHIrF7EYBqOa7rI581JUQY+Nc2G1DxCTquzM5
qmtYKJYFMnFUmsGMLhkVI4yQ5UEASRPzJPMmTQ3ofxhIU/dvOlhEbUI3Jd/upl9i
GPk1TOBDux9zfuEbs2FK0ROytM7It7yWv7PrI1yO0hiu+uh4ob/k1D6DYUMNDK8/
EgYYwCEOR/VnwZkeChA3cTiDTX09SoNUOvpYxj1UUqSg/1nGgP7Bpckjt1Q4pCAr
YAVm2O500jtlUnB2JwHfKEO0/kO++JFI4AvD5ArIucAuilGLX5yTMkA4p5tV0mvN
im7rEb+OShI7riZzBuL/zVtMyrjHE9kqzHQ4V3xu0I2NgbkY/Nhhaxe7tHUdiKwp
4Ft3wVg4m6Orswgf/RSX3E7Eu/iN3JVO23Dr9cK5TgBYX1Vg+DHfBNObcD0TTqWs
lcC8bFY8daWGUePLBULSC1UMFY2azkDE0wVfOUJBaYwUcWz3gGNu3E6H7AbRDfvV
elGo+HLbNZsEkN3wsbh04Naw0X6LtLDJosQZ3Zg7DILW/gXJL/tkMmgM20rLxYBd
AFz9AYhKYgzeDLI3QXZ9u3BbK4UrrHt/vMdOn88L5y4K/59OufeH02UK+lEstKSW
/DX3xnRk8D4b6FJDOFe5c46CeEW9HOPOeq53aNRkEzzfhU19ArfqAfm+DnXLlBND
UTDaxH2m0cDbByJsZ8SGyNfI2L3UACHzWy+xUuZ+yBlQqTqQeG/NG04MxTjyrTOE
iHDVYyaLlAIxUOzGFx1IgHkOEZfHwf3NkEoKcsxYqJEByUDTOzG2O0xizVBqkRkT
dePSA+hNo+fWr1ym334UQSzWKpdofQWKeEfZSe00nsWZRq7+a052GgFRKqGBvDcK
pzrK9oKFpwM5qcUqfGKEBWU1TcOoFQYbp0AM/DKxQT3jk+nTodlRp2NpObAXPGdn
YahDjH4j0jMeTPH+Va+UPapLLY/BBFFVfHRHxGgoewJzYyHwI4HX9bcKY5572vMw
Y8DUTVWy75PncRxg7/E5GTHPt7Cp0m3vdFxhdHxMl18iM2xcOqjXmG+8A9UjsDAo
MjiB/6stugBlSOHnggUjjTHqIkZMSbol8Zdqo3QugXwmzq2qWqVENnfgnzVF7bgq
HyWkhX0yMPhId+RVIjbrHB+QfL37CROQ7E2LAWwE+RrZbgV8yJZ8CFTJRSfK+f1d
tOPnuWt0qHlHEmr92TaNqQtPouKPSq9Iz5NV2XtOBTZH13PIpZRz4SVu9E1tI/1q
AQ3EkhWFWUjndi8HKhdhJR6QdgZ1xcVgzJJfPPm7v4tAQh4MCZeYuGjwOFv4gdh2
6L/E58XVCqfk8Zpb50QAbbIdIbvLnwjZd+PgBfi2U2s8jKnDQrHYLVPCZCatKtFa
Z/UhULWssw8W9AG0abO9aMyah3v+78Eq2vqGVZ21x8p92z1rGdWxrmKYuvUC1Yk0
OaJOkQw+Az1ebA0vNEmokSLt+rki/mQoj2cW9N/4Qm/gFVLrgOl1T9vLhQaz4G5B
+uRxHcRiociaIcYcqDViOSfikjHeJ4mYQT/eExEWk7CddkaB/aKGmlE4pi/HAXxq
cBSkkkHETDDi1apSLond0cWd8DELLgAW1tRQ4bMuzkbzf05V5SrSRANDmEycScHm
c/aFEZJWMHwu+AmsAh6IBARXFHtRLI0d8R/A5OKKWffA8khunSFbZ+B51mZDFelM
TGsvB06DV2SbK8HMjNPApdiYSrV/wuYV1Ulfro6F2SdLXY7UL6ZCXTfKfVkqCh39
1yUz7x6GDaF6TxUwMdPcXBeuQt0XtdQoLNdGMiImoYP374Sf00HpxgdSc4p3wSBz
oTZBBc2KmQyDldcDSiKKR5GrytDpS8Q6dkAXJtdpKdTldWdoA+Cl4zlRHggHEhZ5
imuwgQgExWKs8QxwYah+yJd0koi53pQ60cVKLW3KX/4z82W1waARHlgvQyDCHhOX
aTNxPc3jkk/S648NullINmUF9su7hnE3TBAf0VX7zFTBJfAyOOKTaBFI9L5D7s9c
tA+O6FIgD9DYwocgwgtjrUqA0v5/F6VMXHCO3cGhtPN0dRgbGDrVSBib9i08vyd7
AV5ppXRQIOS64mR47N15uEAvtGcFzxrrGB9fCFSlK+VOP2E2tX0pXfCS16byCIZQ
qgHkMaC5bnLxhPKPXIGMyLrbodWUCP5bifDc2sIwP/Mag4rdC0KWoHypMRP90mPv
vGURz5dSXq2Vts5aJfWHT1CJPQ8GiMPvdVqzH7ltOvy7REdbmyo8M7JPrtwLqBgt
0eEXFWz0+q/DIn75eTWIFfYl7zURT2LlBBOaWnOVLa6qKiupuoUK5ro6XpMofODW
ZhyP93UVKY5TffyMN0lalFT10/sQ0T/QqrZ2x+wgHKHZcfwrcVOH0/2B7j6hWdSZ
I5DJrridR1TmvVg4RAL7jeNM7TyMcKoX8TJmXBsZb2Yj9NYB8OcHxPdeQUl8C7lO
/rMlyoh5EM6JjqAY0l69H5rUg70JgacGlJllh9LdK7ECgJIIil51jgxMiyta5tNr
DxuUanP2sxWwrTRhkHHNgKRn2s/mWUkoTpQx0tA8zaaQMVmptOlEXGUsJjSncBan
R/hftRjrz3wATIl5UVPL1jEj+7s3aI6V2ZVTnp3EDXPj3jisydYPNL8gYLNkRlzH
TT5yGT2yprUo/0vawHriSmqgTjSsATCOAl6UQO2LX1uH1aPNjhjvL3tf+mKGuiaz
cE+F3EKeljxYLzzlALpWb4zfSaU4bm6Y4pv/+lvAYwPuied3XY+FC+gnjJo7Jj1M
qm0/VaDTXUjY3LACDm6pZLhN4Fyp5UANCQjSANKSrzykQH+pbZWKCXZVjX5kWY26
xT6P2/tuS5C+TMxZserydcbDjXrRgeHYHL/TyHOt/RVKVGo8RVUqs2vZ+4hpigFQ
3FVo7nTcTL6Ui6RCSOQ5R9Y/H5XadUDDzkYex5L5l0DUDLN0I7KOfok0lLJdJVkY
Fs/Hlig1mOMFNooQf9+AyCmNxZHfiHsQIAxWd6b5qwqRI0GpY64NNwpxv+iCwqqE
rBjLN+nP88YQA1fowAdgJ2qdxSULDwmi5rCBC+LdFjzPz1J6DJMTCmH6rDkTsIqY
ksf+C2dcuUA0eY17AVUVJOASs6QhvDzwvMuZhmBC/VaEekjxtllvgnrHWzQU8hRs
tg9QR1oLE8L4ngmNJEXq5dVQabxIZVaqvpuG9RZnkeljyiGnBZXYgI1DgW/aIZ4O
qvQ4PABL77rKq4RrNZYQ6n6MsQ4gvJK1TNLqNYn/GXf++AbvySpm2BeRqRXOHxFm
iVNnC6GEhF8Fpz4rZHG17kyR7I+1NV4aluQZ75tR/XHURKph9976IQNdLm2Chw7W
pWcvNxAKO1QkmWA5FeZQWrMLEqf+aSDOF6TIB2Htz9upQMBX3siW9FrwPY5ULgy9
fCmV8H6BSG9DuelHciaVWKlNiGA1l9GSgYH47oVUOKebQBy1MQlB23de53zr6eE5
MDvETOQ8RjcIXycwr2cR/cHpS3k+drnR0EWOcPyxzt3+EVUi4Y954J17FCLcgcyZ
ZIHxmF+49tH/9LbL2mEvkR2GQwW+fxjEMtLadEVmb8OSIM0zu4/x2Bv5vRPkm46k
SrLQiCZtMfaDN4E2arDLFe6sLJPPNlQ1Xb8+E4goU+b4JYxZZDPMSt00WbMGqSDA
A4YizCJb956Y/LifPZIukJNEzeeN8ytI+UvHB4fIcrars8mqkxUFQZARQNhqBWvV
FPiPYWvlpzjjqrxBo9WIZG34QN3ADV6XHf1MYxVOHBpTsRts/RYDovy7qTP4PE1z
SxCjfK3NLdwSvo9jRqzD2eVp6stgW9T1/dZ+CiEcMT/Uc0Pi6+l+oJk58TFA1bWU
zNgjSdbkTd2CKU4ZaFmNlDyDSRuBMQ+CTdHU2NQeUsMFt6ggrD68UlPwlRmNkWNI
A56V+ICGegX2jLlaO7/CNu4qMbECb6iPA2gxuz0kRLAxX8D+2ksa3DrsmmLILhhJ
Ud/W8Y98ToWtu3xjOwv/Y6Cmx8XtomzczFeZ4wgtHGHKw2TQXZyarIF/DTWu5wXY
a5m0zphaAqHMQcmWIz6xHHRB3cCdpWqganb6O1LOJxYZr7SIQJjVfAazcXwqFxjC
hPgszsDO3FmdakphtDhvPiDiBy8691gH8qRRUA4+7Si/4Gx5nrLGhIbboC1Xej5p
b5d/ucENMVxn4XzIq7SbspZ6LVFLgy0kfIi3DSQ1R0Qj22d9BrDoa7apPQ72j0eb
A6C6eoIsvCKitwt9kHIZxGpDZ1I7NBh7W5rcKonTSA5ShS/BNp7sBLHV+l1xDoDo
/+COTZIw4rzL5i2+4WfJI75Rz95466GymU6cOaIWAyVffXVOwkpOoNb4J+RnL5Bt
ayqI6CMuq3njHjbyQXkc9xkRPQHPCVRM04Msrk6MYNMNoMfFhe3pAINtvbDD6J1N
a4JIWF4HU6ZQZt93Bt3rZrt+Cyc0CEVcsO2sF/XY8HDrETgzk/C9Xnjns8A1PkZx
zsfX87m1QS7yv3YKzLLn9QAETvovfVAxGelHTB7tVsy2J14LP69zORsKQV5qjSaf
0OyJWOF7v8FQ/fT+kHqmu2OfRFMQafwTLajVzkdt0cV/KKXcOdTyjIFobC837gd4
JtCqSorH7S94P/SOaOi9XNjofV2g89WDv5m0cw1Q5yj09ACLZ8dK2U+dcNvTaC4o
is621ZkuSBAErUSdinxBoM0qdho+Mn8I5ixVddMbAvTuSGGi95IjhbLxALNRbpGd
SAgvLDyvOnzbEf5sd6gcTuTa8dVZwTcdvxnJQw4bMC3NJICmvSTedf2PF2bkZk7I
TpwMgl5UCABQc7VgUw6KpZbWEhe2dAj91RlOmnuYLP02mkGAED26sJoVT4DocH51
oL8gZ/j7CJCxhOqQFCkFtUDXeCGlYIX6xjPwV9f4u9//ccIVaM3S/K1/sRmURi2U
AceGdN1iNvleK3bfmvKuAKZOySUsxed/BkzsPCbVun76mpuPerFl90vy1S2kHLNW
NxBKVcT1ZXIi9D36i44vDWhKCO4XLalLIE7BDIiJrCQlClMaBX1f5C7Tmm3OPyo+
g/mIYQ1KASH9kisvR8WGrIqMiNxlxFEE0SBFJ265h/Hn+H8+XFMeJbSws4A2Pmdk
GEdw5SjiokJ6m5g55rVs0zzU8MiSNBiWwaZHU/rR71gJaeZaDG5JQMn0ZWmwIMr6
3/UZluclAH7sLzsbqJkskF+aGTu9PgyW109wVRe9lFHkeYbBtEoGYikbHNtUqDJ1
m1SK22kwyCzIOjgo8H+ud25Y+8ZLXY9ti0NMPaidmJc5x06HPcVWyqTMDeTmvDEA
lR25r7cf0/dIEvZcS4M+FM01H3jrSi5e6Gw/Dmvlc5rEhEoDSBRGBnhqFAw0/HZH
RsHioyeW7AWxSgKMUjKfvFKyEzmwrQtjrkDMVGS+4WkY33PPGKbPIghTVdHVobeB
sBcTO5/f3D9+ly11udbBLFSgrO8Yq033zZl4Zmdz6PSWHCN5KDH+/oJgIZhKI/+S
aMFf+9P0F1fyx4U/GJ0dJTQJJaWuxlaA0txPr9IoWSsFSDPq4d0bEQLSKjwUcm1U
vmeBZ4ygcu5wkmf7DnYKmGP8yTGsudrebL+oNjUFz8Z+maeOJpoWSf0e8Rv024Oj
nGpawlKM49UtOd2FUUeyUH9byNgk/nttoAUYGfHtS7wYEbOkVJgCoP0VjKY6NyCF
1fBCd9afabzX2mWPIu+bnKyZMWl507+TAekdDsUVFOahB6LyIoLNEOCHcilq04w4
f6UOSRRMVkEiv6oFOobHNwI4AOBheVjlijbrZ39k2IDZ6tRQpq+eSVtM2Ro6CLqy
ZD2yHCqoBt/k6OHgIJJtcnAL27iYtOy9krp9Gq5owz3/48ic3DZkONm4NSW/gjwD
4UUmLsO3l8A7LAmNX9RFHfk42BPzwTFWZkiFAw4hPEQHWWSXoiEgtKv0k3ZZTN9K
YUaycW5KwAPO58DY3QkFzAQuE4fvth08QTSCvPxHBRdMWIhmL6AKno47Bnxi0EO5
ZFBRoKqgv+gmJaluhvuih4PgkBaVWY+Gec+KO6Bt6wAYJ/AhmvhuD2EIK7yAhqah
uBW/2Pq74WCD2qQSp4v+o1rrIxPjk7Ftg3XPglozQaqh7llM1pw5rsruOjWkfFnK
mkQm3WdNmIkZuBtbhjiPGf7amLSG8dA1//yPlNjAtGHtJddP15DJqH2e37ec9VaI
Nl3gFETKU1vv0BP+dRenTtZ8T1fFhh+Imssh90JdY6FTdPVUNxf4+yKtWYwQ+jkj
dzXRJTzvhty6+VqOpXKCd8gWEGybTfo/OKEEjMcG+lKhdwzg5elahLXrjz3VgSLk
kT4KV2cFoeciDz59icxtkl2NFiYYdB/4+9ROg0vDR3mwoImCsNEv53YbQmJrDp57
b3qJ+1HV5k7YC7J49QtmUMnAvEmZVNLkptKVFDn/Qv3CmiNcCjkW+gvsTIa/su5A
Gs6wG4a/DLMVNOmrXNCgXc/p+p0YLlNeo1ui0Zc3i1h/ypJ5FXGlRtKX5MOmrVwa
mY5+z2I9NN8FffvlrQ9PH6MhkfKOyPj5mfI9QVLVHwEXqti2B4EADQu/o+umgK5n
xtbD18tUGkAwWFw/3KCT4tPcVQ5JUVIdk/+ITMwDS29NzQW6YqU5uu5aTBbaDY55
GeBIRkEuc1Z9/+zLcMJwAbIfsLPU/HTLovhQPcLpInA0D6dQvDuR8EMAwgLp7VRM
9Rps6AM9oEPfnyWQ7QAGKO8BCCXBr4/LgW9lamB3wCqUXpQgmYtMLiEF8eVGJFTB
nhcl7xLYZOqhObPchOA7/7XWfk0jJY+rujms8Lq2ox21DgXsa0tvy7+nnBJqK+yy
yyxGDu/qI1QkHqI00k0NGnDPn6dtRdxxUJyEWdcix6UN8TWFjwaKGX+9KwJcr1GK
Xn3ecc6xpKNhfGrj+PywSGkYa/vhFfYUbIvmKzyn++jv/rAETeE8r4UTnZZr/hSV
EDN+hirOxyFT2zC1tPuQNmqjmMC4rHWpoZigluwTf34VsLlnK5eDJQIUY/dPRvLj
CduFNcCHz/Vd+CuGEJ7OepTrOyf1hImiHbqxf8rkn5WFOvHHD8eTeYtr96KO7DLW
EUTzgGu6ePrB5k/sHcz1EFMWTwMk1QDJIcIDg3qmB99tsxExGrqWhxXW0GHQhgSl
65tVgxZsnCz3iJL3EqiSB1HpQPYDudlrA1UdYm2i4jznXHsZv51O8Suq7+Lplq/a
JucIQDj3loqz/10jvHqx0ltnGnMTROikcEaVdkApPi5p2HDLUc6OlzAZD0Zku05Y
i1iBtEl6dCi8R6uV5Pyb2UeWbDQR7PAspYBLfPZ9NsgmJbgXoKS/xQvRDmbt0A/2
lGGR7+fH/p16YmOohVyj2eGeDySzeudYT/rARmRxXzjk2uIYef0yoWBsBWgeq22G
c/Eg9WvXyem2R6HxFAW6NEZ8qvcPPNl/0CYHJUYvUN5gVKfCxTWLZS8oAR3Xh9Zn
2dntTrFQz0hFuMMaelRxuoax04wOCstJ6jlzc7vnSc/Tf3/5z8uLRO8PTq3Niaat
mh7J6xusQdNLTqwOfuq8c7sXoVtFvQSD5I2pvc33E8c1VExWviY1AAjPTyfXTOPA
a+wL2/sYVAScvb9JJ8OAnUOsjbo9XygxWiC0Athis3Oh8djvmJFQAlnzIfdsbnYV
I0rwdOfNKofcMBuw1mUYvnj+L5ADYOHMAP62VVTNgK5B6xSRjmc6xqKX21qf8eQb
lwgScE4uU23ZGpYy0HlrzHlk7HrG6ZrXJQIwU0ZKB1Kp/J4z+FmXeLyUMW8hOGTR
quSHbpSLPCjSQEYCsO112JqOWz/3OKASn25aPnoFufYZEbJ/soxyinUivJZXnPKt
TERi+0YcCy358SSUGhJUL6T5VNreA2kbViQGOIbD2pBC1dDVB5KNdoE5doD590f7
f5vSjbcdfvDzxzSUQDsrPAKGSnLiZkDbXh/WIgXoxb8F32zrQFM8acGRk32IfIyg
7HpQCHth1vPbDCJBAWBQiEnTcu0reQAh9lv3+DHfk3jxm7inh+AvRqJQAD9lsMKo
FOFAvw4kJLzeayVj/STlpXnd1O8ZQQ9K49THdDDPi37eLMWlvF4mt9flnmoTpDc7
knPfPJJXHJfQTEySLT+UTk4oF6L3R0ge1DzN/WF8nXFS7SkGlaDWxofvjgZUFSir
2SM9TJme1jydLFdHRyadobrMPL/Q2079rJL7Bag0ioxF0Bn6AsoqZq8Eh+pHP4gk
YHi9ZLm2xmKjS3F7ilWQdOsK2SUS8NvOJcBLkyJ3+OzIpSvkZjXYQxDtR00NXOkt
2Z56rFfraQ2gYXt8XuNF4/rEknlukMpz99LtcaGQylvu1qvq9Nj5+P4iCHk457fl
To3cvcDlh9ysW+1CGywj24Pz8F01945TuYj/GSxyAaUJF6mdRqYUxNgEhCPk8RPg
TTkngff00ydss6aUsNQM818iHLx5pxxbmSzgr+JMXbTqmlvG9m8B6GDl9FV2YgUp
4ulcMpT25ujfvH2U2+B96c4cUVBSUSPbmLweieldckj5KGjv+Q5ZniggfJFqDeWl
AoxdKElrXN67ticx12PfpHmAUyUHGHIu6yJeDJdwt4hQvxfZP8hlIuTZ1df67PeA
sfIqxuZecqZMFJtHWhDKmq2gEMvVEhd8/46cRgGFhhQdkA1jO60fuBd1oe3VpYl7
t7rbKD9EE8s/E47pG9Zku3EgSSacr2Fu7WDfcb1tTx7bkaKpEcZ3QGXQLGONhiqw
cOn1xtmGa6FEga3In8kxrvlumWrmYSlBJmY/a4pRaFpYl3kRKrkvIpFSLwESR97b
sUSD/r7mR0Uss5s3gsoeuiSNp/O3q8Aakw6fELzflR1k42d5XcmmJQLTik9zyRM6
GzxqeHaXpu1eGyiPErmYcZ9ESjvgpHfBrTPczKumb+LFC4ISncXiudSQk6RRroR5
13KGcFek0yOg2zjC4d7muQgtx7Aqd35pRcohuYruvDwpnXpzuYCH4W8xECb7+FX5
M/DtCnJbrzQTnBn3Sklo5meQ+aXGErYvoVoLGgA+B6hMeemNOcTYoVpxJuOlwEqB
WWCnvAgcKj/xpKtmRpeNNovWXwNN2EVq+QTU2XtOLkC+oDFQDRYqZ6dcYxyx+s5i
+3NnoQHtwjcMmxsUgqF0VLRnh3gIT85+bJ/AvSVguND8F7Wz0Te6BUTCAlJCC64a
MdvzBRHwU4RMQv1Z8d8karL/etTJ92IVB5KQTlgnDEPiitgYh0a00L/52Noz98n0
86LlfvTwWBeW8A4PrrKPZ/gG8HSdbok9M27lDsyozjYqdNgXPGS9iwSUkuRx4LWX
/rUSbEFKpyPC+0+LHDMIlCkA+BtTMPe2KJLx30hjj6fln2IaOSZtatiLrmr51KYa
DPKYx7HohTRW+do3/+Soqo4pCU0Q5Z1Xhontn01TKoBUrpV6yb4lKAVWEbDMzLOg
FcY4UvRrO7dWutSBPGpMBWykhIQQHkwP84ukj13TwJ+RGXNa7gP29EEeZZvfM3F3
wco26Y/KRnMQknn3JMdBr9MevLIJQtIH/txtvzN8MY9RosCYtwL9YbwSpVzI9zmL
9chlojVyvIPmtw0QW0e2kdx/X3Ju1BtkLvZAE+dshTqQY54d9LU05C9vQ2/xqeVC
NvrGjncC0NvwsiTF+vaoezSlSC3HpfZJTNL4vrzs/ck65plQDuGx30+sMcKtwjqu
TGQozRZK40vYq7MwS8U1VzYEg7aGaPX+Y/VBBrK9M9tQblv0qpjnqYbV9szZpmYm
4UI2efu+yR2iaRe0omF/gOcSHOn6CEbxUw2IXv9Vf2HBG1s2QyEaw5hSIPx++Jeb
wjN5zYZKtzTCOgTDa7laodtezyvbBv8eTio2A7khJUGD/x0Z5kD3rX9gFVhcgYBr
HrhLfwu0mJT5Rd3/of870689F3CIgfyGTX4XO/ej9CQIIh2hyD/xZ/M0ED27zWUz
At5iucR3iP0KpBjYfBpRQylGUInBzhLfVaEiZ5qGW7ywbgO6M+srzkiE4nP6fx1T
Qqdh7QCEet0S822FzflUeR9cffBmvhrVlf/GiVrlbdnkzdjD5CpVgML7o9KlHqf4
HI+wDOquchFuAzb1um1O1UHQDufo44lMH6mAFEEZu9LSwr/k7m7IvZkS0+Lf1PaM
0BVMcroJ++ipOlXKen7oo7aTB9vCm/DVp/oggDht0LRSimpZ+3NsrFhjgw9XXldk
FIWWFJeTzZK2FvGuI1CL+PsaiFXtKb4OOv+ZMa+LWS3zJo4cJJ0Mdg7A+eDyHxV3
SYYgvZ/+Z5XZKwSv4oC8iWG2GMdIIzwAoeL4p8GGxXnFh4CZGHtzF9bjv6w0WTuN
YGZ262pyW8YnRZtzC0I1GnPaIjzXn5Ym62bBP+5vGknGNhMG15pSzhpmOLTiPBWJ
l/TDe1ARZnjRQAslyRd55i38oJVQr9kVy4tSMl4WpdAtSS5oVm+oDNxviuuXaVx4
ILYIwrgOGF//CJuYJWv1KkMvwdvvroP5+qOjCAK+qgBAY7ANB4dHcCGZueDgJuqY
CP2JwdrM3JL0G0uNlZg9x65eZt7tFX35ZRpgZFpMCZfZIRHxzs5sXJ9Sf0F8bCw3
TkxqxzMVtRC4+RW+SAc+ecl7NsF6zjrsPIPNuyka7CvJIcw4eCKG9QH0SL8Yaw/N
su+LZ31FmLtyoeJ5tKVZuSqanIFvwAVTzGJbptGF1pPRewfrNzksm0iDYaNCxkQG
U+sndEQUYND4kWNley5Y8cGKqMDX3kVQCm3ZXqXQu3JZKE0Lqv5Uakv8iejMR9GZ
HNDEBYXxNjYnyenSOR0e9MtTni0ZtjHGD7HdhzAnHzmmvMhTybFdqWU7jpS5vySW
cZFprJbqPhZNnFIzjFdXNyAu6T9FymALtemFhdGsuCc+rabvzl5TYUJzTwHrtzVU
bKoWQgTh5ZkUzIVtPtpSenEHcA+asI3wKrZPkys7NVtwya4tpUO2kL/T4b5slbrr
o5UFnKrqEMZuCMMedYSA2ZnJ7fP8nrDY+3zuqR7d7IJ5U4GOZghLrO9c/U4oG+0j
wjz510HUedsiDEKB/OSV0suNMnW+C9Hl1FWJDsDMqG8eeLbqhItB0Hz+vgvj1qYR
q8YvXT/eDJMS5HZStASnV6jp2YTIzUPRypMCP/zuLpfN3mTPYvHTfB7xvyroxhLR
yj2fRfaPt8t5WuAMkUrCRxrZsQodegOaGzdfjHiw3r8jDaSd7sY7dumPXrrCYndh
49HJnr9lJhk5k+nL7ZvCxtyXwG29tCtt4txANMuYmcl+96U4S0bhN1ks/SgB5s2H
ZWTwgaS+9RNoEhtKfvkgtnMpfW0XubZkQKZ6Hcr4e13ibr9k4cphgtZjMNpqhIFl
ytMQ2rO5nys0imQ2SIf6LRkNn0AsDjz81QTeHmclTCybnfKFQKXoualJo925uZ4t
EWQaYnjLZMLuiF6b1h7FW0VXDwiBp+VRvCjAhRKpI2xa7Z1jQc4v36TOu9pWSuG8
DRapa9baG+Nj2EKWZe4g+hYan9BatR6AzYnmvvafEp4E0/9Lulapx03wXlvwo/p5
tt2nNolePYXdNNjhn6NXpgCy/7KYcvfUaIf4OW1XrLwbQStYoDWi/AP1AEBjfy8E
/SIyF0OHGKffq0F5pVr5goEA+GzCpmXlOI54WqmCq++waJJDJJ6nqigWY13cKL2y
ZtsBfGBI0FhX/jTJEySgcAlMpEXBRwoD4A1JLvDhKTC7Wj2s9YblwKjbU/JsEeaR
ieDZjwcyDKGZ5+Pf2tWErO3mrCFDq5sveWJQsr53yC/O3hUKqfj9/7ZeQ5UmS3dg
eiCHQFMVhGfxXIPJLkhR0VyR2m3U+yZcqyG8PzldJzO6OmA0X0+4lSEGGhcouZYC
zeRu8P2oTfPC5ZLIBVYuUVsKjHOZAxwCGf2g3hOAITCn4GFr+cyTds2iBf1fxmu3
l1FA5Fg6g2nXbKdn7WNiUTMSANCQ6UKG37VlYaS+/mrbxaRZhoOwvt0gUE6h/kMw
OnUAy8tHmEZnkRovpBcV4YMDK2D8gfpH6V1nMZsFsw8rNSsCWuQHWTCYlHTmJnWt
NyVlpW1BaSL31tDHgFScDoD+7NzQBqPnJMxbUo5PELzW8s0Hlx6E0nkosGorOO38
UrKopCoBO75b/b1tP3PhflEVQleMFTsfL7QG8reTJcj/PrKFe8nyWSLX4552HAFL
N6mOuX+EpXgQMwhhXJ69Uq6XOw8kImy7wrRGhEgUTtnOcbqNNFHalpB809is1TBr
MwVEvpwa0PjyqK7H7wCQoDINkM/m9aHrT4wOFNXrIk+9olrJfWFvb5KhWqTFOY9k
ybb6k1rHFS7k5r0koH6ravQMzVZQjGEMgi192j2S3T/fTEsZZvSlQYvqDFP2XXaF
1Jz7BYFWKRjQxWVNnYsDqj3TujOxgTnHI/Mh4l7z4Pd9H1daiGgPEp1L3E4CwkSN
1v9DyeTSGzEhQunov2vO4lBZwKKD48rGyZUWQVW2+544GiZeP2nBylPOUkL7a9Ia
FwmNXA+TJOGnMVEAd6zHkcu/EQmrwYLUBzMVDMdyegfntH8n8NiuzqngoTbMKlyj
R5CpDxHMKJ9KD/eS+GICEhmzWLf5roF8pYCa58WiQzVE8jCxqJ1SWo9k+5+4gBvN
sI/73YORfl+B86yre168VDokxG9P7+BkRDbpoqSvwBSDmL3m5BLwCGIRwmqfEOjA
icQKaHpkEnbDQI5R0vtrmhl+fBmn/mVmIccpwl/FWF0ZuBl50H24jN52pUeEgoIt
XTKbgDsG3r97ctTa4WFHLcAn+uggXO2V+xkiM8TGd0L7L9NCspaPB6Yo9etLnq3y
CQrsR/vyxyRZFRiEhwo7GB/quz0KH+acoEnF/+cPa04jYY1WZQKDdIcUkwXWVbY2
c79mW/+Vf4uVCPSZKMC0o45BhufXA1K0KDPovdiH80cvy6hgGYVJuwqhwaGakRDm
l2gfhBKHEKc2hG+m2LklF0HW3yb2p5mpeJx7G8moncmURTMhxrrhzGfOVsY+/Q6E
97XW447m1fhZzbBeQCz18Ha4LeXkavl0m9y9dPpRUpAHpE5R0psBSiWV5hlxL9YP
mfIsiHy05l/4qjW0YGVYWJG30bqfxbwEjHMi3Ax5RxhK3AyrA5JASbF1XLrruHKL
9tvl5/UeGVrkUNU0T0J3rxReDJzszfPAaMptgBMplzpmUx7g03nWNOxppm45/ULg
jj+RiuHxO19twJHRZ3Qp+9hXYaboyH0+aIVhSOvhSI+DRKWWNMW1fVNs0yxLqmfL
tnmvux4Zk8GxfmoVLn+NrI/JTzay4igqCJXraBg2MYidDLB69TryHg+pA+g5HN80
v7xFCxpHEYLApJiD+BHTfzPiECI2gfAdiEm9thnzMyGjn+DQ8xuQ+ik23YMFK31k
KyqMsQn+3hxJGhbNQTQdLSm1DfsHXhhD1fPq55O2mIvlfueoJEKrDTQa9ZEyCsBh
E/woWKSsWfZi9RSBvScpKLvOTmZ7ZzXjdyFmgccFSsmxALd+YgNlpVkvy/MuUqzC
DpNdoP+WodUlRL0R/MnoqCzjUJqfcDBPFiBipQfc4PSesa+JgewhjhyyGEtDAEzb
6NloyWNEotIeCH4jVwIKw5ZyMUxiII41r1RTTfJl52DL0WxHjhaahnHKut4jeTZk
CwGlaDKHEzrVmGjR5x3I8Cpo/2efcMKmHQPG/TWnCifdd5GcYQhQ+2MhJmZlVm5i
zuQ6pKF96HfM7l/Tjp3OctSKdazXvvcgSVAh0xQaqXfQbmhHIDz3LCP9LYPtjqU3
5D/zUclSwllD/qq0dqAZoDhYPhPZWOucoby/+L7Hwin8bm6mH30dfL6tysbz6ULi
q10QwcPCjgSRKxqMsBuKeSEvkQmDdkuFicVi3jA2bHJ33xjnJ2wJ5EZIc2jIAr7U
WRK3YVax7mn97mf9E8Xr2IMAKtHOpO0K4IDDyH2U961iBaGBC1MrYSjOq/60jxLN
8nwN4YSwk0+kKlOqMPv9iCnrxLFsxIXLiczQ4TCvyBQNFvws8AGQCoDhksWB7k5V
ceCArFQj61DZO9bSyv0kHNZzCL3bXswLWbVNGB5fqjZIPHlTv1sFey8glq4+j/JK
Rzbd2Mky6MB04cVOU7nMunmazbWdPQ/O6BVVM4ltAGPr2IGPPzm3AzMBz69uaobt
7vc3RF6TEyFMHZXIWwhvP5QwBGDo8wMnGikaBsbsYtdYdG1Ym7Yf2HU199mr8wEW
L629IOODNqLPg8KDCPto6zDVx9Tp+/S/3YTK41aHos5mj76SDJixFRrTBhgpNeM4
HPsBBPzP9q/uHku9BIQaNY2ENvzZ9SC/PHVO7nbfwxWczpXwTwu47lAkwxFvCfmC
mSelw0Jv0TLMEr6X9/6YZntbsUa1eCOw9kfjzSM+R1ipiwOCqBrlpPtGTdCj9XUx
1vIPqSGnnCDkpp5szISOO3UnW8oS4k3JyGIaPM/LonHorNq6CdOYqCVanfChDBl4
zsUDchAZGzIEeD004kDZde0o9zypH8Z6PsBDy87kxYePLfG455VSGTc6pn+xR6Q1
GTPiI1aVJRy0ECSs24RQ1CzRK7/3vypZdZFQTci+jvlOa6/1lybnqvsl1RNuiIa+
vLkJqF5mkdqsPKIBWKpHfwvYfTwqrs20grhlLguvEKAwTuhAABCTYtwJOExo6Nc+
F96dy4Laq9w32AT9EJmppdZmUvRt7LXjeaS5RhDlul8d7VO26gsJcyvKShIP/98e
OOv+ZfhJiNPwy7YGPkQQyHj9XFCX2u3m5KtpEoK2Rog/DkNxoC51ezLMWKh05Yg3
iQXyxsJ1OMFLanGf6ORqzCVi1eSxBMkJr4ROf6sc5GmbM4cOxSh/wtgL1BAEyYjI
UhGUK45wk8J4wCpgm+RqYoJ9dQh9LsnYzGvRFmIYZ2OhXBCFPIlOPa1H3VWeBObG
ZnICoTxQuhCuu8h7KIWFW5E3GEGHe4wr3XVA/OIUsqNgry9+XiPxCf2KkUkaW/B8
a1+VedhkwKl8Bfh9JZwDO/qbxIaA4hOQunlfplKoYqBybmrHkhDIFo8NHc5EEnE+
J/kRcge3Ld7+YYff5QmEiq1keM8TJr62N5EtYeSVgANeFohQI/VmjNlQ+q7HpVit
N+GHnokoxcFF9XjfAa3N4DD2BwHOHWgfjzqcHlhIBoW/aVL1kZ6c4RWzHvo0huyI
GSIyvbMFBiHzgDwdHAX95Fgxj15o9GngYwC1E++cRk3+784egsV+gqk+etq2+8CB
ltf4QQ0TnOylPwa8TIzJCuHNJ8th+wT+dd2J2NZrKuuTCwHyuC/VRYCk0YGL82Sj
jxtkdoEu4AhDZjv0mPOvJxXAjYOJTonmAU+IwGGPEWzHgbSLGBso2FnO7OqxGmLv
Hk79UEVZazgja50rj8O58ZBJ5ym0fSjhgICzOQGOUwZfvRD0Esyr5w39D9MFlGMj
IsDCK+E6GyP1HzqkGj8KGqmhKvkAb67Mh8N6Y5l26iUPuFpWBuEgosnPw8eVQQnr
8FX9/fCrBSdVrzdkzB9ADkVwPwd3uRxIRix4TFH5WEGaQ2+j5aS8heHbW+N9riq5
eIaRZR+UNuO4PRV2PQnbBKHUfYlV8G4lwzIQwmtZJHA7WXbDeH6aD+l9kFvB4GV1
RVl3wwy12p+5MFcNBQjYhTXDoN29OfUnHYk7H+wIv+V8leZVKOtCNYhqCzxRZtcH
ireaUIGyAkG0/gRbh/CGtnlsA44kF9akGrUBokAegNOB1R2n3+h+9WDbwItO7wIQ
pUxek5wIPc3g2mlFu6eKOZBgJiL69I3TaY85BIJEHNPOoBRx/j3ZfP4ov5TB/pCz
nyzLBQsqLstKg3qHuRoS3/a7mO86tQKukQoG3dlAnXe/kakrwZy1Uy8XIzYaVmTY
ACTdEvCILdizE96D5AuaUL0Ofz9k6eDkzDTw89msaif1aQIWnrn+uRw6hugz1dXX
W7doVQkjW/WrcTuBBBZQWvo9mfPG3i/xdd7Lrw6pbepRYbZF7bSe4gUYR2U/8HYY
dIPjWMeMP9noaquKhNONK/WT0zHsUjbFQ4ugvCKCekScl4EbVrGmV3jHxVZHfmbe
HsAkocmwxmfD4F44vb6Bk9hS6sUPhwP1Fyt7Vddhhw6XYevM3JQuue8QMFz6lnYN
II5GUbaY6sbL8WIubFv/YVluS0oBjBAKPRd2Z7DmyWilpuS4st8IvOdcTlpjBskM
id+WlTDnRUlsz7rHl5fdTTAcf4YXp8scEIn9Tch34esecgP2EsRLNJ4M5XppQSqi
SYv2QnYNo3EIVaAATtDjwsl6MujHInl9B33lLdYbBYXO49udLBO4GMYnMh8fCmwD
qh1MPzwtcgkAAeC/STHcsSvMHTEM6xO3benSUAMp1+EWxqgHajmDuhgXOh+zMID3
0CJulrnlNCBvU8OEcwOxPowyLsGAUmKev/wbrwrhCH9I9LQxivh0cvSGGb9hrYx7
3qb38dQDHj7PMvjGEOY7njjTR/QUXS0yJWEs2xwBHcgGuFyjWuGVCnzycN3wOhwv
Ax3n1R4dBzW23/PkxX5oYhYU5P3x6ZvQxtbaWVLiZDKiyRb4QXe3mkHqYidHf8O/
57IArVCAQjisgzoownSeqjzRjx5GcSUXtrmXCgUsRwc3EofxQgXi0TP3rnOCgFTu
Ktae+RL39IotBXv6jgi+pAEgeg2XVbf91KsxshQllA87WBR5aF9SrRo6bX2gRGNP
V4rjNYA+VJfsHwCYnb8WhHjuEvnXNJgS1SnnCtzFtSpl4sYkvqPLwObLa02Fvho4
4xRwjcMZP6ENbA91OQuac4qczQYFDwyhnm+pNrmPRdPSdpZ+SJw66ak2Dg0OoC3+
zZauaZ7pBtzKP7ETDl5Mz4HecjCcq16lIamKSOPJLXfzbXpZrysVpSUg0IbtQJYr
wKI3tnz66h+Hgf3EQX0jKWmXQ8s2TF8Rxe/0TxZmYkXCfLaM8na6yhTvyqLM9l7M
2ELPR736HErggRyMDmKEv1Wy6Qi/P2fPAu9wbckQHo3do5ap6DEF9SAir98dgWbe
w/ODUpjp64d6SDQ1PAkvClVxAkr4AyEQGOPx1rYw1tjYFfiWReVkyK579wA+6b0T
vNMunCpswFJxe5eTnJJCG+sFPOvOESA3ak55QuKlA62BLdmKDczYtNKT6EZzHytE
WWbaIGYRPJm5ZoFWOt8D1pybLRqP2ZUdlYcvbohePIaRPckBYJdicpH28/yypCk6
Bux+/CLef057Q4gS21/aijTiDg2fruvWSLsGKTnKwA6D9Qix7vHJp9kVsIhrdMV6
HXwfr5+VxFIXiGLMsiZVj7LWky/tJ6HwweTrCFRvOeuXPpidPutj+T+vl06RWPN/
aPJu4oYZqylYQl06JReyyJF0WMtHNZc+PyQ5kOLyYfBpaXkGQFZugtHobQ0RIw6K
HVC4IqqwE1SLwjFx0KLAR80ALn1ZVWnEo8YCVb2E2Uy/Tls1INdhIedo3gT7Z/s+
v+pIZhe+xyCQ2J2lswp/Rvnm+2doU2jp4MYcQ3opQkax9xUtqdi13HCqHO8vvYh9
M3yogarIBHjieEZh/8S8CTbEnrLF5UvlrOht9rGeiD5m/a8J088S3uyNESE8Bf3U
qSdbwcooTJduk8EYSDTskQ3xlavD+/e9TuMek5XEq7QosuW2QjlCH79ZyCScfTae
Vtqry2amDY/vyNCvvqG/yIAMzdA27kBNKjP3XmhhWsia94oOiKKXSdOljuD3FFkN
nbydWLbVyviNtPaRYRmzcskj46O2Xb2L3N/5AMVOpJUtrO7PnwFltvffHsFzn3JR
ura+/ovPa+4UFVZWzOv+c648nId500zywlaUc6zigM6mYpzOfkMwp95dOfQI7sOW
XPyAPY0E4eZkyenxicTVlLcDuvvyg6Wosz8MGcjcnyETKLSXI1l67yUDbUdNsfMQ
W/Lf6UyJ8Vcrx0W73PMGkwePsz7zpkRs2iwO3qT14BIjk7GP49NvCidywKfceqEe
ynLP0rYdkCVJwRAATtQuJxMJMJ/M/yBqdK173jvUu72PCcYqnwDNZLbIoS4bi+mR
yXFiPyrARcFZTgd4J6HmqAxQF52Wm4WNXYLYk9KXJKG9OXxGNcb1/wJ+lMVhU3NJ
VsljL0hsIt2Lpj1EMiSnzW3Im9ZHh26Fg6HBecXkPWvyLXfD7AiLnh9RigkpBNpw
N9FnoXmZiA0fA5lMqx3X/C7XFUXSkpMPosSKf5DQ8TLJ170ktxWgpQytYYrXAVYV
hMzJBw+fZbTGe1UsxczxFKYcZcJ0s3Mby7wZlxx15gWNgNGRma5UvsH9bgYlhdGO
4cwwn3JdzjbFMSQduhUr1ApBmCJiGS2QxZx2OVNno6q6P5j1HYSUAdi/WzTcCbXC
OxoSGljvyfjd5HAcnsGZ4iwqLL6cu5N8y6GL24XvOXsT7y6JhRRQzfd4Cy1lr1bd
h0GU6tusMYRBWccau0wUR1qoChxw1HV7FeKEYdFFzt3VfXL4e3OEZ+L8D8XzYBGn
57jFH0m1aTwEzY3oiXXClduUWHSjxD7eCeckTjE3MxmebAN699gGpMTo9SCWulJq
71GdfA0cy3t2TJylNCf7LKeUGL6RI5stERAhnW41zUMraK9ZzHZfT+0vhbeXWPFW
BRf3WzjIBz7d+RvfujZZCXI1DHGSxNgmpev7Rkjg43stznW7dERc7CtwMBTNplv/
IqThUa/VwPTv/0+xx5bsGU1HKprMqEmUraElVVssQ3B9/qW3gggrCuvqszfeK2tQ
vpfwSXC+6pKN1GT6o9sWlc29tdP25+Vu1NeGXXR7UOQ82cs7JJdcRDZm3LMntbEG
Kq/qtd1JFVjH9dUvm/u8ct5VamtwzwPwVAZf2No2TNTvS+mi61IRJi1Bn8pppoY7
KdOLjz4N5JYCDN767OSnTL4yGh8NPvJvvMq+HW9LcU7H3GOF1NItm1yGxxJTIxBJ
M/5UwLjE6gfK4fs+VmYJEtC/iJOB0D1AYuym8kO4/zzJQoo9xoCNbqb/W0uQcz/a
FOAODSPoNgZIX0xjbDS0HKr+5rFxTmAR5iM6KdniXFMJD+rgIkP8dPykeyz3CBxk
dFtqCs3tKP0RI2RAuXEz9YFxzupCurQxD5ijSoOptv9MtkwVccPCA/5bb/YLjeUJ
dA5s65ZnkUlOtbZ/rIjtlleljrSxqSKnBqxNFX4CJnv4SKcT1vksG7RjKBOA9DAD
CO0S6KyzK2l3fXvdg3Gz8QEoWaD+Yko4WansaxIw8mBW9Y4OIT1ZjfQLdTRg6GVL
tIFLAhiKWsEJ0HGerT+CSz0PlKF2O2kHvfMRrkBfirwp1PAXZqlBeZjdr6VEIDH9
qtEOTOtFRn1WL44Dg0JAdgn1W2qjZH6QqTQ+2yKdVTRKShL3GlFviEh/ClHq13/w
miLxjUG4xaWyTbRKoI/gPkB9vT43c1vRIgYcurNQrhFc72/VXPfEX7zfmSRz1YBw
aOlEYqh1HWGB48cLQ/Z7vTrSG54b1ulA2rKkvpUElpyaL4lAY9ZaGKbiBLpnq4ng
rXHUTaCQpoGUrhzBmLNV83vWRbR1hwkfbHaObdZbC8+UO75sthDMUA1T5sOQJrx4
Epu4F5P6IwXKWYFDP/xu5z7IcJEahkNn5rhFIUSL9HVcjl012yooDN6BQdoCNbuK
ckGSeYgcYbCG0AruuJcU0pNo+6EhjwC/+cnn1foIV6qqFR6kvfyKrF3iZXcQkS7o
/fa9dR0kaBpF1KNK94pZXtoHlwIZH9qrxJDSDE/r2DTsD+LmyburwwAy1IN7txYc
xl8beXkD/Ho4ZbP7df0SjuWsmnl8wefrnsn/pLIS7pzzZBLNvoJ+gMdm/TEKBluW
LfMrYdMzCTfygMlxObaqcAO7fd8JmmYBImQfqrl9UfYGAiMv8DB4ec9xmqI3wCSF
BiWEX+0iBbo2anuvIvS5cyiIduNbz5XBgMm+uKlPbgrRN9XrMuOYzmNqn0I2ZVW9
6YGbJn+gtnSf9750OO5vMX/PxhFC4JdvKBv4j7oNrAgd0LoAypfVVYP1WSZfaq0p
Zb0MGck7NsSGjDFjahbks3UbeuY8eSvQWbvjrZD60TU0Ee4eXXOBbDwWZxtIOcs5
BKOcqvjVGWMQgf3AxcLyw4LNCnovtHO4Kd0cW0yWL/XHLWtx0TKngXTLqywnFmsm
mx5+xhYrALRYTErE0zFNT8PEZ4fbaXvw3YgfMYVg2yuK4p/tdieBPH3HBoa4uILU
X19nvfA08O0xDfrVO20DeKkm2fZm22vLOPimehsWHnEPf2gkcoY53FLwDcvtUJL2
N7TeOAgoFgMsWNr7Dt+U1Iwx0b0GD5Wt0atCDrD2Q+Ck4WESBfcNfSWmc+NRP4En
vXbc+FcDq0n1px/WnEi3mZ6wcPJ6/5ImS7Pgfe8Qu3Q6b4ZyH5Nj/Y+N+cuXy3xS
b3ks2lE318Hb/P02aO9+jra6YJjUU06o3nVUYyzqgThEorcHgAu9O7cXd3V3Lxw2
c/dEb7z4qaA1wWGWIkoH7CcGIIpOQMrp3csH91HVtUG5OQYNUzhcKsACXh/VWceR
SpPugdlks1YRV4oYwQugOkyJrz/4uhRdXnKPD6NPl+WZ5UoO16SYP8WNRKH07TrJ
OpTJxAatyBwVOibzp51mXJIk0wm1WWZkKlBBdq9+4XnMGLclQyUVuF2khRB+wqIG
5CpzbGm304Feo1zGlBrr1IYrI3JUWBuHT/9TnW/GND5N4f8TnbKDvKGo7jAsOW1j
DSxZSwRiVLdMGHevOVR184WV7PbIBJt33FxPCCmqniBpP//0FLJorQIeGOlOmmdy
nAnSt4XsrRDa7LgGUYWJTfGdgtoI//6fsyUYaLZH5W4vvV5ktoLxim1ILxaASI//
dFHeV3m8Rd/66HJBKK5ctGqJsefZcfn6YV7TR1UrPJS1yCi9ycm659dQtq/E3uP9
9H2N51BDNXc/5McnE9tXd8zBnpMNqWAg3RB/F9nJP/rIyTwvnIFxlLU4WHmJACFu
LT8T3vxu7Cs67bmti43ZinIkR6KjZrAHAHqcEzS6vc1+1ouDthr/Umg1kh13R8qX
EoTEWI/4MJL6qbsmPgjbjkoIg+n2CeibMXeG079Gqykv2yBOT10R2iNjXBRBrshM
Yryw5DuAKT00J8WkrZa4+4zzbiwf1oVp5iJ5ErZeNUv24RX+/Ys7ZHQv5fTzkGhg
vemgrI8VoqI8XNYp5u4WG7qavFBHlcXKH+jzqlEYLW/zpiwhcHw3p2nT0aG4vfkZ
zAsC2i/tCCNpMlwr5+v7io92ODaEUCD+WgszVFvVEfSMMVOojoWRz0L2K4cyMi0V
aQN+HKF1n+cRumMkDJJTMY8KniYuZj7KNxuRBtYwLiSs0fjbCaNBB4Vzqno84Rws
A3rdZFJ0L61WXYBa1c3wXxB8SwiXOXA+kwKQ1DTPkjgfs2M7iX62wcsZJDAAoU5C
3RY7OkLd7pmHy7ax/CDjfIBctCK6SqcTAhdCv7+zZKuonOMkww6fuljgXqL28jfw
barDpfUdL1wz0EnpSVVMxHbVQ7iA2FWc+8PvkiwMETxA1K/ciQTXONvCdTmLtjY5
TeVcpvJeNP/5RWnztv3Y4E07hjQVJuq7uQ2DGohzvAw2AJmp73ke4kEHDh9XczcC
I9q8DewilREwllpqzbKGD8VAP7TeFqG3V/E2tpzVl+iYSjfH3i/X8GJafT6kBhJm
JLgTp+1Qx/Wthtyyne1qP+m+d0fOGdgd8DTcTfZIr6K7wdxoRQIU9mkO9DjUJeUY
bt6Sb4+TRbNnbRQY+EJmOVKvMJsviRA3nvwFgU8Y5Tm3k0Qx2VVImCi1bPSZUSup
KnWSP2oWrMuqkNFFWQo0sDbi2yxFF3kHoSsOPBz/k5EnD+HpjDgpgOmeM1DT1uHI
DGvGtbjFElDGPLdrfe4GO5yufmXxeUqK1n4LocAbjK84ufipS9kbOFRwjVKF+2Qq
XVd9c2j+DjrQ1KMNpgnLNUv6VByWAWAk1oPVvBvWVtgda72bEOps6rrjOudruM/t
SsAzOz6nMGnzns2dJ5AC+I4pso7i6bLBC7Dxecl2k0dBM7MvAXoBEmZ0KNunfYyl
m+ez9FqGo4E8aFaXpoST00JRmTxAQChPpFqdVn+IlPtOF/dvVRoPUrzQuzPWEG98
0Shrr8e90pZPn7nZvJOVWRuYAR7e6SuX88miyioxxYR6f9IDDGIWzmgWld9pdQVI
lsZZB7xMNCLHIUThOQf90eNrki2382Whubqws0D/i8ijgD3EzpiWscOUDsu2I7W1
btUYmTAGWm4xogiqpSyq0n8w3fxfnKDa8hywQeGSy2aDqMZGqzL42WrBsvitm/ix
SDrNJXgWqL6+8fEfyQ+3xwuB+sTqscOia79rRvYicF0U/BFIWO6XDr680BLBvYcK
6Kd0v48lvHjh/mlDMQuNWUQhFLR2rEqwywUX/2qCzr6vzEiqCMZmvqpEEexaYyPM
j39A/1gTR8B++05dAuu2yYTvWTlnOaOhqWQX5op2ljzmeHcncLn6kSEg0hldsf/1
aF6cIk2MhhZCvkIKQfmwhZTy/16E9t4+cLCDoYYlSeqWBQW3d1ocQfuWcy4tJdJ0
FuvRN+qU68OFmir8dJPQX0AB2bHi8bNEunIFEadY6Xq1y6mcMNsOabd+aRAQip+m
lSAPxhC3r+d3NBGz7Mr6mxBomy3C+ADontfO5oaTp1wOlxTnSqNwZTtBrHe6xpSg
rcQOs/dVqnqNA2MYicocctiW7lECH0oDLTIiyi85N2IXChpq0VpreFhtiOkuvp3U
PmWo9p5DNoNOFsCCq3CeKCkMDrKqcG/TDGceii+I7QCIOKBKIiROXFGpSnHj2phR
XqH7Wyc8OvKtJW5fVxE5X0QyZKPhKDBA49Kmy5/YpsvoxClGqm1EKFppgX69QxOz
jG33jl5el7ZEDjqGyobXP85KrKJ/IRa32l9oq8vE9+S40cVbrW/K5pUme1oBstM4
NdnnteafY+/BxEnqLAWyl6PEjD9UHVsADbaZ1uo1TXzefeLTdyr8VM7txr16/c0I
7QJp6b19Ac1t+mf8wBGu6czETuSe9/PW6R9pVzQ8e6gbYH18JeQ78OiI58UpE1ZL
VedZLKFOM3XbsVW0I5O6G4fqwHmDwV5OMwJlZftRqbi3r7r0h8UsS1x5vmfUm12a
Zwv5QEZ7cwPhAMRXShK1fGTsalZqoWbEnQ/zJdYSd0pz6GMixxMJCuIz7N8MuE+R
kZaqAc0bO4/nhdwhvViUHOLxBFu8p+SiR+YhBr0U7AP0qQvrP7dmMoTVR20af4Kx
MFZgdKRjW7R6VhLxPSqVALBytZbt9MxSmyIHbXtT0lvfmKrt123+YNWYW/RAbFZ+
v0kJMaCb9AfDKt50V5KRUWCYN2zRFLPJJcypxjADFsQGTxKWSxBNHrEBhuqGmkzN
JApAwV0IuiPnoLr2brlDjRsZYOsK68QEWybNHJgZIjNnkqzXZX3bb3iV3Ls5uV3X
rZf3qG3xitGAcoZ7IOzyG/hwEFnbIA9dQfVwx5hAdv9j3w5ux78hICsXt+HHXMqf
oLzojIfL9Ys187o5+X3KowrOUl89z5FRgO/pwOspfoBEAR8hgDaikmtTS3M9slu2
VhnR4vpYFJXFvPh5e3b7CfedqndkBZFa9ZlrNlukO3tkIEEdL+Lt43YtGZwjVWwT
n+/TNwERvGL6MQUtqRLrq/tnOfSRHAJanaDsIWGz3qaSald8sFgdeav0NkVOZEUY
iSpuB+oiGLPjEMJDuNlTL6KLOQ2oi0f4kIR0V9j5H2fUZX/y0/qFW6rnqbhyAhv8
6LKFNOPMr1k409n9JDG56LYt9kCxOFqVjadxQqTvjW/yqInl3ez1uZxLagDmffEU
BN0NiVYsmvd5MUWctZR3HphBpp2kbRd9x2Fer4P2KO2OraANsBnv2x5r751HS43c
+Yk1PEcNh4MZn7+qWKZFKvDnxYFdRnMiP/Z3THM66C/tr1srgBNm/lT4zJhOwOod
dxXe7Hc0Hjmqg5fjJVRBA6FLCoFbnKn8eKOJ3L1Gz6WbNXxA79fATD4N8A9+UglQ
P0ELCLFEci4vnTBaAidZBm0qEVFhntPaenzkk2jEU5HpxIK4NeVQHtlxoDEX/tY7
OReGKb7UoqCIn/ACSnRRYyPhZBhwiUlyVS8RmIXLEQQ/+6vIVi/Jy5Ii8bv3RSAv
pj4ue64xwKR8LZ8JsFBLAPAku3TIXdXF6PCCavj1lHY2i4wAPjArlDZwVlsRNvTD
MuCu7MGQEKolQDGW1gN/T9Ao+HFE1ryaQSgjEP/VtSK9IhFhvyLbe/2jq9PU/PwD
kOo+sRtn295xW10R1rfG/Njleyi16koT05ogH1tXk2vAZzbGb5CzwxvMafSUMctL
HfSfeHAQWWUL8ASYlPlBakR9Iwi35Fkx44gCkIkSB+rnFzRZJl4V3QgfJXADnP54
ftB3ukWmUxtUiaWLjqI6laudfSlb5YX4+57qqWOUbun2QJq+VU5vmaCIlzaAEdbo
k0/wN5ZHU2r1bI63v0LkR//zuxlptcA74IeEfie/yjq+Y+AdsbPDPgoZpEvfa4Hs
sN2/mo6EiNqB4DL5v1UQwgTjEipAHTReTPngnXfHZRT8hxyjF1ZFwTltLagbfek9
ld1/RaeI9v+G/pziHO4/vb2ONBm/0320KWNqsX2uxNS6QrsjKzjg+L10eiGllHhv
zVFT+/k3e/syyLuUwNXKvt77Yq/zssGhEIXkWPKUTvxJIm2egpkc5S0DrzAXx0hp
qOKzYC9ECeg4p3Y4m5zNtte6AbZ24rOOtTBESch8mZd6qpGUV/RbS7pGXeFhDF1q
IuZbpDsL+fqOHyKanmR5P925abxzI3HG7PBhwfmYSKX7zPRmSMwkzSPqmqne657j
KV8qEkl7Q5IM5hXPEG4AobURNNusO2Dd1Hyy/nlLXpG9Kn7z6A7n+K5LYw6ZAKne
dck0ZyNGOVShiIo0KrCNWAs/Cxc2mAEebKHxGg7JhvSMW3N+2j6MCwvbUZZjjBVa
bQrfoiJAxo1Ph148cx+utsEwGjQk+C2DpeolQu1evdp1xa3v5jMOmFTCR+DEF6sk
gHgDGszdQSLWm/AJEp/QW9EcP8Rbock7RDnC76ab3W1GGeS7Wy2KvSeZIQ+731Ku
8lo9uNVZ/nEX7mgQIlFCDQZQWkAfpEhUOuDyqtkjHWJNujz71N+l5qVigXUXioYf
0OhM8n3OztK0Wj81eoEgvjEcVWmF0LREAjBZbaNOJ6E0Z5w/7/dB/uqTqjEzGRuz
UenL5P6dzejpNUhQ9v3MFWh8ZwqwxmPgbPYcZ5dCAE15SrN4X8zMNAWV1uM5EnOR
tCkVNa8xrmyxWTXxzzkvFO+bZb5svhOieP1tZVvtcfnKzakyTY3i2FUhcG1+KOk0
ujWkJc3Ar7bWBU8uhMku1kamPOFqmCohyFWbQYiJDtgzOwaQ0dRoQV4P8o7QH9ea
QKoBR0fxJBPcW0TR4JhaK+psTW+hg2dkaZX6/ZgLRnYVSZFL+eBnXR7LlUIutGzW
6UxLb4QWvjV/cIyVWzDMsaxBuKwDY5RbdFvMsDMnZnk5gjt78LSXm9Drz9Q5qf9b
R1xH+rRQscfg/JcKtPfbrVvLE+7ZziRhiuQe6G+QYDhUK410fM/Gf9+fKOoCWAax
UWajDQE5goAWzuUFVYDctEm0iKuZEeqK0Fk+xBGjeuhPf3BbP4aaeqFJkqL4uj5w
OaWI7GpnJ4IoJvZePSXuFMMKA34ZBniY0uuhTvmOyDtuBsoNOliorx6iRdqTCKRO
A2qMIUbsvdBOESeVBq8yVBu4yqjf5cCBnAiU6+EoHmDbWBeV71dfF3mcZwV/HZLP
4nOAndfd2ssISBlrExuxtN6xpbQeCw0pZEeWfGHrfI+DI8LDrs2FsVSmKrgabY3Y
MgVQK71hv4oDWAawkGrRy0QcCY1RvYTfMagSwRxdIb5oRLWZYIbBwalWI8U1v3iD
hYYR0lZJDl/1NtXJgPwpbK59GDPASJOwrARZ+LRLTfRln6/BnH0MNEdCpgBPxHrC
Mij3uqOq32oHFqzBdUzstsbHAdpwlYPZvbQ1eKpYGHyo+YpxqqMTTUyR78ABFxR1
572oS2rdQ0+CdCx0AcNKdIf15WVJIrNZsrTM3qcYQq7eJq6Ep0i8ZUYl/3JOhonY
MAaMpYYUjJY0VQaCzgiXWmnUyMbZQgBY5Sls1y7dpROatg8DvQ44j4CAa1Tl2kdJ
S9qmHvGPrx+BlNGqj4NRNHWFUsb73/WJBj7R6ps2u6m+mW1pCaPvSai4jAfdZKyb
DiUnQq1+EJRq4tULngGM8msskyZGkHRrl6w17k7INYZcXd+LT/ATpDbjL1EjOteR
BCaNUyz0pbK+5ugv4Tcxl/om1fiAAc2h+YLW1m5oNRzB+l9tK32QkGG/5XDDACg0
OoCzJNKAkrFNtDVM9j/XmeoxJnw1E6hutkVB9u6Qo3Ef9XByytLeNCzk06FQCMeV
EeDx44EEuj4jym6OMSk4h7m56fgTetyGS61unr+OkC8EX7fttxA4xrJPjskRDi8I
5vQb5A38g+gALELjW6uYdK2gUmTurQLFcjMAnRblshHFo5DoIXw0qhHwIah/t6JI
yMe9GzBft4TaJkhs33cK+oYEK+7Nqbl5WlTqzB478sgBPwkGZMCsGPSPwNJYqgnW
kLoRiQD/WGviMoG8DUzfMkqfH13xMaJgac4H5AMGdt0w2BfBMLzuVXfwWAy+ERmP
61aY9m9ATEhhqkfQb09I4rvDOR5DfBVlMJ+MzlRSpnNjIdzExCrNRgQI+pvVtFxT
H+mv0mxXF3seXAdadanunJTjv4KYhlbZlKgzeDKBpw1zoirpomZ1YXEWz13DV811
aJnbkI28EGXpZrdcIX7Jb/JJVYUX9lEGD+u3TyDX+0+IJDpW99yTYREbm4rHevVy
wtnvsvCgbIDFtqS3jTwfnNycK4EdnefXVDFVKwSnUnB57dsd78ump50N3RZSkpIN
tXQ83PU6jIZH9mft9KnNv/OyaQ6LKFeDTcCvRAFl6rqUNUu7jCkAZOZwsI917SYM
bN5CpfeItNDBbGlnnfiqd3Nq4WUeCQDRY9Tm9glP4krWHdDm5qQW5fyX+V+wny9K
Pl4hFheY1r0zNsvi+RIr7vNTvlOiZLE8r8DOxh0PyfdzE4wEoQrcshEDcKJt7//5
lC+B3/zEjFK9FlUbDIuMhbAy8+jxVwZts72H1eoSO5moJ8A5q4ZQRoP1lUibDNw5
k1glltdYdYhHaEBtehny5eP10IDygumKJOQcQzTz1sSu5+yFANzYkY5AhIxiVU7n
dDc78obi234uyHFL/6g4xWWA4A6zn8QwoA6E4JxGd3uS8utvTtdmMKL4nAZhlSsE
NTR7Ep1uA8WQQZKN5Z7LOA5Md3FYjWz7fhUj5bgWmvurzWkha/EEqADj1pggToS0
okm8VPNVI6/LYyUuG+Wuvx1GrSfq+4dT3Ca3gLHY9imKkJGC8HTwec1CNuS5DDie
vehdJOWTLajLzRcGDUw3e8AQtR9aJmINQ8hG3DN/UyoDnOTtSpogjDLMuMAhL6Xx
s6CP5MYC9BlrmcWPvG4pEi3O40yZwW2n0v0hyGuIh7u593zxJzPUK/NsbSoOh9wN
72nICVKe3l5Pgm8maDXQwDwIPHXOeQN6RJVfNayUmJ97R9BcI5pvMyJosn/Tbsxd
DnrUfo2GE1+KzBwleq6hexskkGKLzCPoLFyZKQfngUX1qd5bS4A+2bChWJFVQCbB
xGKn7qv8y6C22y5O/vCagUEhRBJQvHQ6bLgY+VuqUe7nVNHI/OE8Lk4cIBOtJ872
uJTauG1BLgp2rHBBy/EWJ7f3G0+IeYEflcreE2bYnO2gdIGgviQTHDY/55HtGGSS
Xl0wyL3s7wEPUX0c3YRIdTx4gdwV6AzAAjJVhHpBQql/h/Aefwq8ngues4Uz4bcl
lKwvAQPQutwg9Lb76HHn/Hf5pBNIOBBIEY+bFh/uj4Bdli/Z2mfUA7LZs1QDsg4E
S9Pf2/I2jvN2As5yny+TSUzz6WTulv3HOh8np/377c7w0a9AyGKkFPYWN31fa7oO
HOpFlLMRpphpsczRa+ti5mO7oANBfOfOQ8wZoD35uLFKrtvDhluNDRuRR178Ws/w
fWJ2pL5ztyQXq6wb3zf33N4P9AffM5hlP1wlWy6je/bgQtuMMOBZ+RSpSOZ6ns4n
wSqsL/KJuHRPRKM7I7KMj1rrrY0FhR7twJbOF4fuxt57wnvtD050od1S/AAMSZM6
tSegMf/gNpQ+fsH0Ft2WXf7kPMjupe+Q/KlCb/sJIeUFQAUKR2ZHzjtTPH9cEvT1
nFYoRnRU1M29UXaz4R5JgqoV9ExW2Cp6fnibh53yXFIqHLhHf9TSTqoUMEJuqW/4
+yTB4YTgnHIKia/V6z8+wwfeYs2mTUla5vwvZES1mfwoof582phPIGNq4nCrmVvK
Ry7UfLVr9BS2hwdlXfdKHKCW9VZRNByu39oc1nlGW1UCO8hSHk07jPRAzPmzgFPn
LJUf1yvBCI94aAxZ0LdMYltIg3Yk3j7+1WwoYlNfUAZpOfbo4xzBE0wDit6GnbN3
xq9lTRlta+8nDlDWpitEOtXUJQLRzUN4LUSC/nLh/KjxhRvgGhbgkjnOO0+3g8r0
XOrNsJBEtvtMC7nP7vCIvAw3/ecddDDt74x6KwPx1XCEPg82xIMlJEbqCMktrKk7
uQ6HEsPpdTRFSty0XSSTO3YksLKyaBJc8YjmvO5rYgwfyHgrIzN/7ewuMrJ5xviP
lhUI+q0mDWsagPNRxRnwpAQNlWvYks8MQ2boFfjELncz7Ez9Yjpur051hRJQOVzP
a/VSh9hLtsLKLsLZyw0MlMgaqoMMtFho+17GiEaMsKUSyUFzWTVQrqKN23IshRas
szlvDvt5TNyY3hEcnr8aJPJ6m4m87kLIgsfF1NvP1ltmCiDlw8d1wEkQrDEMWsNs
sClCa2lCzyFE7slvFtINK7cHZM/eYuvYrbxpBj0RZIZm6VDB15aVGSjf7gTCzpOJ
euCkToU0vSQ4EqXOFGIi54Rh09obE5SV9Bx7Ro0tfXW8nJPZ9Msc4vHkYHJOMQY/
lTWdl585yEhO0sL7Gf55x7+KjNAstRl+1xgGKcGSN4b6vef5tOItVPgq2ryCJJTB
xqohmtVVS7C4Nez50vg5snG8fbWe+AdNnQOB3R7ijRGbnIrRPJiJ3/ifpM0ZY43s
g4ZGHsCX6ZOAcNPviiJl3U+1YG/+MUINIj8LskZm9SMwD5tLAHkoqC03ev0Tf9ZQ
4zES5cgOCRla+edZASf4ygq/cAbyfuqXRJtfq9tjyfpGw5/cjkKeGbzT5ZNG5PlN
H4wfZTRhfUE5BlyQ+HCLOo8NCRVxHtnP6KLEqdUpQ59Ji6KJKdYeS9/t1wN8SlZ2
aLq982XiFVuc8HMV4pjgf6eZzVcicSuiVC2zT+9jyVTj7Td682I63EvGVklL1SWN
EefaBXJS0/+knW4ogrVy1GDyaVPG/kRap6aVF8jEPiTVCjKHnREatGzuhC6ZY7dr
jdJdVQ98fBDS/s2yv43K8QeQl5MB5M0SF7ODEvJxeNcq/Z6dfbdHmGJ7p7/lsL5U
nHZnioTAB7i7msU0L8ZfY5minKWYEdfUfQTFHxW4tH+pCgTu7ZPVnLxHQIN09yBP
vWTAlQXcO7tCGecxxBQMrRUGZ56GPkjru/Rthf5FChKXZzVixNmVlY78xzZXRycO
FTn/iyaU5+Cu/GSwkZ0rRq2LwtGW3jSpFs4OiKtsHlv6DZUQ+y4qB4P6Up0n4lIp
BJGU0cMrl2sJNPof0FCxz5I1TOFTxff0fazbML6lCakPSnweRCjP/dZ7Bl3MFu8Z
+i0d90KKPr/LjGePWZW93H04DnIVSwtjLeQCszW30EmUppOo4F2rgaLWoVsmrjTJ
OrB+6uPhQY2SG2FGZX8OC3Ac2JxpEdAr/GJAB5bMRlRRX5Rnr8DerIa0ga9ltw70
mXeVVtFWzECV0YVTxFmA2rN7lZpA7CZB5f4Ck0aC2j7XcDreGo1IEtOlbdFQc6uf
VZI7n3aVmluWM+omXPsnJFZZsZMI2McpXf7q1buQqqiWIIcV5FR0CRvm/0Ba/PXn
d3X1quaNd/9C7HMfK/5bqDBiM/KNE0f7zmpFR1kaE13rWWebjS8M1L4WWY/IrfR7
4l5mYux0PWc41kxW49J7Roei/L8x57wdm5dyOA/ctu69zGGCmHXiJ6Ycqv5F/3dG
qIRT/lFi8M8nV/dU27BacfaO07YMwwK2SgLc+W1ENxFQ8xlGL6MqjvXT6KnIovwu
IPcZdjdRSrOA/JxWuk6d5NB8288uDHvCor+F10PEvAN1VHzykehCfTLACufU2pn5
aGGXEbt8+Bh/Ztv8ZDUW/xJIfhbRdSYB5x7PgQ/oDC1Z377kHJnxum+Of8z2ZRyZ
rn5/3FuoAwYuKFJZ98KTRIhp8DKhrYlKmorCrMsz15kM0BiamVrSet4Wju5QzWxK
a36nOqV38jNPyWfIza6iaqQ+2m5NE1dz19Lm7I1zY+471fVhikeubzNpzI14hCOd
/qkiIjcPh8hIZ3piCo53ES0/DbRJmkiSgxpj8M1b1P1xfIQldwGQSNM4MW0tWWo7
MlSNaVtzprLLa5bg2NN14AdHY9QWcQ7TGzRbaIYLMPb5iTGom8A5c5MROX80wTkt
wJwoouqNlyXedyZZvwuxC87jpohZIGH+gZxq2TJ91foJvsZDWH74uHrtEuz0ZbLu
OvDNi6FoJD9lmgpkfU57fmlOOe/+LbZv1CuCqLLjTgcmBVwLSDlqeHfZaMjKu2cy
Z6WpYHBrvUCFi2xV4eiW0cV69TeGX7uLYVFq7/B+7NgybkHzQKWVpwmqPAwQWRLw
6Sh+DnMCe5e3iGcYsQIFn+s7eeHCz1s+pULDzl1GX5a+J2PhuL5kusBl6UQIHG60
5otwQatPF2t9aiTuijD6a/MLxudsmYvPkM8sjwF5KDh3lXt9b6udr9NtxcLjuLFQ
7TEEjaT/B4dzVv4iYIdX9+sP7BXt3Jh43GBzo6HoXMaXoGETUhsRLeF4EQNR1aPE
8Fk8VNYLpGwH4x0NnQw7vmThJ+HnE1r/lVbhMcy5pU3Yem+95oe05qa+CONtZDV6
JXzUDigO/6VreDZnqJXIzuzXUcl3q7uCz2swmXDSEe2H5pCq2WQPmOfvEvIQxncx
zNt6nIHJ6tfz4/4Yk/t1wwMc06mWCq6NPdm0hCr9qlGBPKtzFTMQ+MJ+OGC4RXuF
Ry/GUyOD1gGsJMmxehLuvv1xpRpAS/JUJ6Fj/WVqw83bZ22AV7B6MZ8ZmqICFnuo
dgLyrEeWfQt7Q8gUb9HNHCKfWA6FT0OL+9wj+FO20sfZiIbn64REcxI2kyeyGn10
nf2N07feG7js0kabX580Vef8qrLh20twzR2wBh0WJ34TtwO4+9kRGjdGaHnyPxZx
Y7yXoDgYoVfgx2rbsI+zZBWj88E6B2cczpL7F5qyViZsuNGqL1bbY5ouIutyc4DI
9E6Qn0IgpQUYll/+Bxu3zsgw8zC4ryczwCfYBvIox/qFTYs2YTWjAkVCWd/ChIho
VeVc/8TA4X6vIhlBHgAGDy9i2Ka9OCu5YrbWk0Sc62MZFTOez5H7hywq2d/HlcfO
hMgs6rI3e4ZtXtmIQYJV018rEcGCBkgBm53sZdnkwAknab+iTf/ZdOTvjtp9FB6H
S9xLY8k059qbzdP5wfxWZRAUrP01LPTqDqJUyq2U1/fHjXkA/YSPXr9ES7D9YOit
6eHeJyNJ1Mn5Lj4T6T1FBub9PlB8NLBFon0DEVAHEmCALaNjXXh4ulsdZ5EcSMXK
a6+nl4HLYAoCb4Z5do9LVdFb5U1XKNlJMIhFpK+vVPpgG6e2pLTqfcxlqG2TU825
UT1gu0qXP8YCegj6u3Oz2AcDwh+5qDfkKoLK3AwNPuLwqNRcSP1JgrQwrHGYE3z3
ygxuh/IIs4FH5VNmxHYrHJ60G3VCn8gKXXG2Sm2t57dq4ePeAjZD0fGfGE6W0ny9
v83hYYlQ5ZYgG9Wbcy48YmL15BdCak/VuxammWRlSIdhFwsEE6MHgyuLweB93gAm
Po6ahiZvgqKn6G4phDMwS56cMkJhKGIczwnEhb363MWrBgy8HQ+9ioiuU7w3G7PC
74A6uJfSJoUsuy1wpvRJxdqyfF8yR1A6AjhNZKvY2Aqt90aBsxV7hZdOp0meG3Mk
N2Mr2nIfGepn5zH4/yAM5OmvgwtG2g4jO+Uz/XfFU1Fjc2PgWoIYxz8CvyZ/vhKA
eqiJ8386GDdIqGifjvXYBX+eLRY7rRLCOEQeK2uS0i+WskbbuqbYa3T2duhp9z6x
E3mQrySIIlBi9WkltesxGtUjomkSTzpcWVF+gtRPtW/WaH4rrf7hchUERbDv9QxW
iUZlOUBER3e3k+sm4l0ztBvaWeTDd6k+aEu/VfMiJgM2dvrfKaS821PAGX0haCHn
Hxx62Q4KsRrbCrNRi3tDgI5KbNqNvLjHGsLgFIFnjrzFQoip2X91u46yMR67ECYN
FBKT0XzeJKsmz0wKc3q6ffTWNw9O836t5fUxOBdX1ApoiIjwQrctVxVmHf4Kd49L
Jf+UbzhOXr85i4m1bSY2gzweKiksQkHPZklQiph8pKue5Uc/13gTHSZUfmz5F5SA
kKMxjqX9R6NiIPykNULWO4ywNn5hzGCpd3rUpwV1irbDJSLpK6R5nqMZnMhSze5A
wUoGK3zRxEbEsRLSHMLb5o/Wa24ugXeH46e42xQgOIPgqzR5xr9ccjxlk8MkDUAZ
lh4f00mOhTdrWCgh1UpOlLzKo+80tFec9jUVlOe/Bb0nq543wcrwL+0T942/S0Ot
e0oFqZe7yyvtqcv70UtQ6pOPZsTsYqypwcd9N14k678yWeM5V3gP8jYtcFCB301j
pMBqw0FkfoUkT3Yr+cuZu83Floed0LXq+zrHAQ3K0J8Onl0F9v8peSxZEAzjkcGC
QGSfKly5jZ3MlLNu72um0Gg1YHV+xhhMbsIZ+9LwMyrs/34iaXX9QNoweKWaio9H
mSt4OJC5v27F6edHa+XKt5TYmwpnz17thM4/54uW6ZfmvPBRKzqJahY6hCw/eZ5f
R6ldR+yrS1svf3BQyi3I8LLugi/4YYsZJeLNUFRTi3nBISrE/TAgCpuov5kB/LgL
T+mYdiKmI7h2oexOfc1+4I46WyvZ6ivqry7Gnm82cpFE7d7bLG6jaE75Py3rWla6
3ct62f2b6oK7Vxf+r+pKDIZw+hs2KyCAuVetUYOui7uWH9iiAp1SJRZPB0YdkWUa
Whf+AMpUykNtwEIH+5ID1qZuF+RQb60D0UnRPeFoWnfZvJERLjnxkGmC/kCtrwpg
SDdCCJ8fNwYhhMxXR8q0Bp+JU6G2U0jE/YMVKILyRzXZe3hof00GSz9EwTHNXvlW
Y0AcAadescWMMB3orcPhxxEA8UhmBqizA+anrIvjUA5K0TfcInB+NXXpzvyG3woD
wNzah3Regif5AFwRnWUeqhVwJurPjJtd2OSnjAlf0Kb+N4s+yinv4ZF7TswOJPrR
IbxDiWkKKKHXqhNJjgBV8IJqrG3p/azVxlBaYMXTID0eq/CuiCdIbFuTB1RrjPeh
C/hnXYnRDR2RDxdKebxgt9MGRJyIm/GHIzvibGHs1zh6uXOY4xIthlJYpe/g+nq5
vzKhNtamrxo3g1OgkgA8CNb1loWCHJtcurz5xvdU1U1pODWrAYiFPnMRpYeyvfc6
noYhwZk/0gzHMniJf3zRJMrP6sVHikB5D6ruMHSqPOB92DOXG6RmajH6Ly7jdfsm
OAA5KRRRToJVFYBkb9rMhT049nQsvLSmrZZi1ABFHVGN9p15ulQeWMBU3EK7DIZ5
ZEdQydECqzQ+oK91KpIhnOZrd/PnLxODqKyi5xUQfj8vDKGXfn+FR4ZiezYx4JJJ
WFSJdZomK1LEK/58ucRTuHczgHgXHS5krvMgwMV7xvgW5wDpJwxsFoZ004Og5mcq
GonswstkxbI0cHa6ewFH0/gMMFXmoUHRxmzY9Wy+2vUrs9mmQUcuFvtzGJruTv4b
aJIU7obUcUnunGN8RHWsMNUSyj7rr09Eq/lasWWa3JV3myLFJtRbkNixYhJ5WFqv
yIIuxtsspFTD80wJK6t6lhlfXNPTCNXfXTblgU6LIs+w9RHibcEhqWryjXCwkIce
O+dh2QlhnLXFonpWVZD/hoN51Wv49tQveGrIruW5FFQUeg5nGPn88+UPiKIm6G/R
3Ia5pgBRGPxjveG6arotVi+P21EajhXdguhmAOsJyOX/3OgWXN6vTY/5oumCh+qo
3LbTu7DH3yZkw/HLvGnANXA5bmmToSKAzCRhuKUhrRkGQPWUACtL8oVxQwN8vIdq
XfyP0qZ8UnUb/qAAKC1fK/df1LcgTfYIvwOW4FNcnxT+7O2c2lBZkeX6tO7y+zdC
MdwxAMxfpL2wIVXWqI/5HpVgeqKK9TJC2WsRsVM0zpBZj7iLCzXyckUrGJEFYmCy
pmVJixiD2g4y+GMAdu83cG5Pb+jKIHkoa41zgc8Jo/uTivxvMqpBjDcwettc/rJW
njiS5Q6IoP/o1YnP7QY7B7OX3yVwNOJ5n3mCvLmT3vrXjJFCe24vhBNctq1cZD0S
LVfMbvJHtKJ56pQojdbqko49WhYskCbaDLlzANJeMAp00PyfIgFmBZ1UYGQ8TFo1
E1BIsayRMpEvNc4XhR71KRySPcxmrofsxTTx3mwHxiA5nufBmttUH87p3K5S44i1
/gjJrC5L9V8gt18mlNhiXFALqvqFF2zHOFgdCp/qkLvL/gJJKN5zwfxPllHC1yBe
kCLFTHjKnKvskGZtkgwTmOtH0px/ZXgWR9O7aooQgb/S+sq7JppRiuDJn1fHhoIQ
4XPZAdEInLenNPGw6YlmWRTihJ0XcCGHOZ5jJ7SXh6ZjBBvt3/hlT//ZPSfZvdyr
BEe/90YZSAV+kcd7FLczaDHUCf/knX2/9kvUeXr+KBTJHfWQpiPwfMFq7gEqjyHg
yu/wVSxFSRDQ4FeFhXag+q9VUn41TkSEkhtm/v9vUybJwZmIE+SwMKMGSYwrIStf
4U4QaCMFagNCOvRHU/yDHfi4dTADtAADE9RS8SM5mOt0HYmPvrqDQsANyD9ln6i1
UkTYtcsFti77aBHB7eQCCTXYtE+FeODBXvGxOX7v4Q7Ug1iJc5nvB4Ci5mTPJMlC
VCG/zDPE/b5Ve2rp6GbuCFz2IVJ434DXyNqsd/ijzJUeWMM361YOAv4uwOsFrEcs
QNXKolO1gNU64xJfTIK9uspqNkjcgFBO/u2lCPde84KF+eaYvnd551LuGzg78n47
dfIZzrorm2Pm+CoVADba0HtIwpWPNno3GHYG6rGACcEvNRXBcTgNoM8oEjB0bZr+
lx/K5sxN5J4eEzNYi0dFKP6981G+KIkrfvAuOJmR1GF4N6E5II1ZYqNFge1o5G7U
+vPbgy8Xn4egDujnLeeduCw90+mLa+LqDnkO/j0JArexPrOuU2NMiG4TsqBlQzov
d0QQ8fQGdYcZZQFtKl4Qn8MpeRSWAb8Du365mFUsPMhErPCl7ZuACsnFb/PseiQN
qEfhXNKkzgPJxlbmupSkBWQfolApe8WooGKZ+0bF3fRsRJ/F+Ov3v9UFMNq7KnTZ
hMuaXhe6//J+rb7cObXorfz/LDxh5Epf33YpJE7L6VUZl5qFqj21wifFnipJbS+p
WvEl0bvvFWMmE/OFVTVW/aYyzsakrlYmhxtZajml6NBM2re9t7OCh3B/3bTB7hXA
ooMRe1WnDZFJarLo6diYYWah4LCtfk8x7ZlU+8vtyLLxUlZf5KB7EiQTspJdB11F
43RuxPOU+VS4/FsjUs4e3GPK/cjsHj6MVdniF/I93ZpioZ7CBzUnVpQOY1Etf+Bp
HfCke/bqKXfd9XBv+rfGCr/WW+A+OXlNkHiBc0Q0SpuNidi2fEYGOHyaPA+7FRvD
qqWNxh5FQwOgYt6OQ6IP68W0bY5FNN7VJ29eqVaEvG2iOHqHE3Y5bJPsveZB8APW
djbNmGbkMjZsY/Kvt4X7BLlS4BeZ83onRDm+pcjwckVc4L1t8FFrG5MXp/V0qaG6
q6C98O9BjaS5OA0VPKUjvVve08PZphdMExy2Qu3oKXWrvkfePZeuqMicAsvIAkW6
RRhJRYbhChG/Bcant8zZYRDsCEdBTEebWfZP1CSjMiMSexTerBII73H3XHc3k5jD
Goa2EyKqKLWXzbmPXG/bdsj7ADKW2bDXBwhDMBNLrvroxZMJKDorwkmQM2g+NHHP
Y2yeSLr0xJeDDdsivP7m4EadbDRMwKNpVmDHpEe5sjiPcY692xbJTGAv8lcwjQZr
hC9p156jjmLuUNbJZdsSfdZHXHlda3OQyaGeMFX3wXopuKHAX/lEcT4e9BUCyahw
SrROBL4bxyXeCPXO0MMgeT0l9X+cY358R8qCASMM3mhEQH1ZZsisOvDONpU+U6jM
gYg7kfSV7uSAO5oydkTvi89E1XFlOZqnPZDqKhs/KTrHKl6LinciuLNxuXYqiCxA
FLHmwovCAuu1k9YSXNIAjAvI8iOFUzmMpltstoM1GtMeCkq/0hx/LuDU49oDZpO1
MeXDxIVk5PK4YbBc/SM0JuLllHMMG2zKKT7PuIadkOagFStxsg/FU+JCjDPJEbIo
aMDwvi+nmNAycaInoXFYpHayyKUOxMYXFnGDTEZAeRBMMvyEm2lwVurU2ufY7su6
yjFTVeZk+zazIGEzEMfBPyMGgLdZiATaboriOeYegGUSnv8zVjSx+mVlZKrt1e2F
UysZMushisOu0C9qV3UlGiCOpnwnM0hXfqWxj/UsbBEqyjSwVjUektYUDg4GDuoy
iWAS0pIpyuzAx2JN9SIqyNXtmPX/wsu7/MO5R4BOSed7nhYuIcqMQf15nAwAc4gf
Q3rQHVLWYQDHIxhr2hQsuB+sx+UZqjUaT/VHzpl9lea8AY+kYrkqs3G2gurcSh6y
SxrYrXujWMnqUn5KGEHrscDb0J3R410Y7SMQVz4GscHPKaRO9pGMFGRizNGf4g8W
w8qvzQHHnwEWd3cteAnhM4G0sdq5Ih5fbpr7zGbMUhHU4gs9D3qoRROFxwC80rB3
L2hH9513F6WQ3n1Xsm4Hl6ek7+Pm+hmG5Uj53jophM11dt8zZ0h0nqzC2N3lf3HJ
9gxKisuzMAJD0uCULvpD8Npi1y0fQGAOkwn7Iu5DzY+Earb9p63KXkzXf1WbAtfp
YPNr03P4mFdK/mvrwgxEDhEzJ+ktuTZNsFM855j9zTS3QGOLcMZKpZLE8yhqkEBl
+4CaXX1eV0Ut0Dk6HW4aFYjHST5do653yRt1vaJ0HPPXQ/TbpeboQbvbqSt3E7jQ
tGN518XapnRclG6iohYGucCUz1QVt9iloPpE5jHibPqsovRHJRwyXc8gPoGpGqNQ
Ina9j9m9i6LOmxiFob3yHYB+A5cj1m6gRJlwVPCrTaGwpeNLIKoogEqB9Df1YlLd
X/c6207W8rA6om9L/FFeINoLbzJuoCM0RZNg0jIN7mMvSfNBGgJghCGLsocvSjJJ
Um8rM6UkoqRK+cNx4gbp/Mjcz3Ck5DxraSJaupmFU3vP3qo93kTT5azimxZvSJ13
Vs4U3SMpHWmC7CpuhVXqOafspMssXnyxMJxx7M+IhCIISTh5DJThcQ9C6vSUHMSL
9m+imCU+ghxvq/VlXsf7KG4NXIwJ33g9dW5B3Jw9mfUK2w1yKbc3p8ESrp04vg/n
1LFzgneQgNw4srUge7ZEN2+vEM7VxRLU9Kmy6dW+XoeP6Vnz5cJxS3Q2rmIqweoU
pPFCKQvHnNfEneTCrv8DYQ3xi5gXVylpQGQfgMblwCkBHWGW4yUjwPfgtmiMIzC6
7rV/YaoFVdk2c/LFJVPqOFf/36pn8Ggr+01t51TNjswa5ewFf7JeGuj4jcsfX1vJ
Q2u8u0aM9DuASudnV8JgJR2L4B6N6JKArNvDCCMeSrKNME51yu7obk2fKtG1UngG
mzK2tmqFwPI/YwtRZeZnrTAXmC73AwYS+CJ1hcfoniz7FQ1dWTPYnIFsX7VLW5es
Q05Gap1zEHOT+/eR/Z7B2fZsRSBmctgVpg07x4KQ9vDvyJZTgrIDWc7VcUYIwdag
uU+Kw59sfNOp8ohcRDHZHEHad4l8ih4dy/AtiYUZzDYJGOEfh9qgdI/ExpuyBMT+
r76ri7Erf+iqMWf/zFw1J1xV9aMbULTU5iMYpKMYiaZQsz2UcUz2+B/PCXerz/zA
MmJTDtDHb0eTj/9b9f/1RB09E5WT/gV60ZMBqsa6qGjrv2b53C5CeqnytfzhNMr0
PKhg6AlpoNWTozFZAc/HVwO/AC+HHQ7YF1MGH4geoU3NcUCyok8/Pp4d/1WrIhgw
QtiQNljfrre+lBAKaxURjZ8n5WrELyRPvT/nLJquaInjDL80AP6oOAjmG/P4jQ0q
YzywELBliB7ThvDgI+zpGbQhY+9uP72zjZI/nVKDq8T2AdrOiAzR7o4CU+1eDNAj
wURWNbO2bAAnzeie2REf+5LLZ4WsHdJzONi+rfTxPYYKHDGXtkEP6VPxS/IE6xE/
5iw7ViR7y0Kgi0YhvdDWc61B4v0yWR6ELc0TAQ4oTYanGX3BeN8MGyZkWwBBkaDP
8D/wP1wTEz8WNXp/gsPOx8KVVr5KzwcbLUFVypZNbwqp1k79Zc0gXbghXh4rNNLP
jz9XKkGWwKuLc5QK4qKxyTpsJobuC/wR46pGUpeAss8MWkBTOxAzwYKVBtc8XQLj
CVv3ywUFnikmbbziV9RJcHVFuH3Kuq688gH4wUqHByd0K2KMxcBIOQoO2AuredNC
qAGCXdfaqgxKvKbxRGE/IfnvEx8RnXnI6vf/lOT2A3RllQ6Upsyw6rfUZSTh5ypM
B5rux8loFAyhyZ6uWWjcZy/0JFF0zurkbW551D2OfXLxrInf3s6d2Okzh3kbujIV
Hv28AJNBGsxHBsBMEp3QfWqsmQiYhi1dioToBjPynglSoAICn7tTMtHeYT4DRY5I
0qv4qJXtac6TMKw0W+9CJDlwHkKsENZ5EB4J/VXVg9BCaRV/aj90beq/1pg3IWvA
hPsch4uJNmxjp6YtasuuVpKHmm5B9rpVfAjr9ISGj04ETlL2YwOiH+znHqpTW3z7
tlkOOWyl274GkmF9okLRAHNljScieOZk+flEJ3N6TjRkvJEBHK1nfA6VlK7RHVeJ
mgwQqtTfgkb0sNhXhygX9Ih/ISJGsMRYF8XwWtFt88bxbsVQ8WfgB6OfvxAwGwRs
LkHTOYQYgfxoVUx0jq6mYxCyBj1Bap9xpbmj2ALzI/GG+XVIl/hpccDPdzwA6rEa
YZtdM81oU6FEwpG8JhocKIzBCGiIWE2kqd0w15f+8YFu3JFRWCiCnsel08XX07DM
t/suclhxn2Iz3+8GkuWLATVBFQ/kyrCmjtsHXSt5gTFmcIXAOxcjcoPPwYMWDseN
yJAjbg0I5aR86f9US0eJD+jeDxLOADPcQQCZjjj6El4m7/EWV/U/eInLGenEkb6Q
xqv5L+fIzkohUay8hz3HraE+qxNzqUY60R/dLyXei9vqhKceRS+Er6IZd7nwANWQ
dKpBsyNeqiFeHohhzpuEzOKtsZsouYzMSp/R2De6SZnu8laDBU2H4xHCc8oLxpN0
50xT/pgLuFfYAduuHxY3HjWyR/szkBYWpCxiQ4VINmSp4iS2GAQ6dhygCtAOPbWs
oCugeqTNCVOIlndn9mnsJdfpw5Sb0cNvx/QtB0zMFMARQNyOjIcjTm7D8sdwxeA/
gCozcYSDiiPZzpJIjxQc7uQVMO9SXmtxURSAvm4BESx61eAalzj7SVWnlC12o20J
l2/3XmMnqsp1X6TvFzKGKAzaCpCgkOD42LNQKXpzFDbRGO1ZgGsc4prkbP+ONAoK
RRgRl+2jNWBkSmMma9ctn/wEyTULpk4ckeOEeO5qzedZ5i2ouhZZz1RnhIMXZeZ7
WqMHe//k2uJfTAP0LEgixMExpuZX3pZOQqSqm/8jB/iNfurBh0rFTR1CjCxuEuJK
OL5JRf6YC0N94k71hW3rJPT2pMutGyuR4yOUCKnX7p7QfA4I6W81Sw1uyWYZeLSH
vICDDLSo9vOnCGZ7mJFQexWzrd7roUMVj/0rFDcIKgk9NKsOoekTuZKQmCevKudx
vED/tgvm+KakerbpM1KSRATSONjg74a3V6fuh9HJWJ0zLYViSNVxoBCrRIv4qvUp
aQmLTJymOVxgkTS6RNIyRL/Q7byMyHOJVNUQF1zh6hlpB86FQett2ZwDL/ZZmx5L
jl+dCWiQrnAwrBpdXVZluqaAdLlWGRn21YusIJKEWK4rpB6nB5x9kioqynqCyrhl
5Sqh5wm+txTlXSGjgRx1C1ybSIkueYeCrCWMnmcF819IijpxVhfhBb2XNV2CXp2d
aeGBGuoCYlIxyLG1/ePgXv8IoLHL3Tj9lPhZy3KOpxcRxgTGzfqVd6xwqdrPcVqE
cct/U7TlXWkgBKhEJfoTTD6IJ6h4gwnxI9Ri2T0AOAnKSLvwUJBCkv5CrIG4jN3S
sPNYvfqifGjD7zpZILsTuX2gm/Nz4BWMUsVBVSJ0GK0vAeJaYoN2Y0oieeRuXzBl
lDCpmy2T7Wg0IGYwqz5a/0xoOJlTj0OoEfL3KDWSRuqCGMxS0yPBvtRdhWQf29u9
3erB5S2H8al+iFl4cwKITSirwq/p20i1c2za+it0+ekvwdNlPJFqBO/tC4z8J5cI
ugNuZbv8mlKIXiCcOXpQeuV0rIkGqbwSRz8n92LikiU+dvmnDoXPvHzhUtAyLKLE
vrEMqGnRQQ0yyAs7XOP+RxFYQoUalBzvVhvL4n7i8wBknpv/ywlfLmGNh331mZOF
x2J6Se7ZFI5ADHNZjogUPzkxo1ERHbcmiilqa5FK8eiUhCY1dtaaZG75DS11xZSf
rAxbebo/7iictZpTfGwhCZPb3H5CRzBB/M6vI7rd1HOHy4AYLqhNcSV7MF1F5ad7
9wVe/Xfk1smumwNwvmNjbd36t9wdrVkt42TNr75dqpt4sCxXYaxT/pj8/fpSf6u5
mVgNKJPvfHxoadzr2xZPS7gddethyr3wnyCgQmUvOJugYEZCANgFwU2fJXTu99Ho
Cf9nyjjnrmHAuu5N4gPWMxp82aeQfeAjNBvUym8j+HMzWkRoPICDZY+vsyU5jBjv
aaBT9RcuJ5ME9X8nOrGU2TrSbFiQX8aRpCSMjCCpr+qO9rEviC373RQNztQ/ll7u
KeBkS343uRvO/gZWpKDdKxNPuU1AbW+qHcYEBEon70iAr3CK6mb9sdsbcpyH0uqU
sDijmvLlXRxEN60VG8Ezb4FZd6nnRLRJHHegKfaqBedf4/LP/KpKvGo8f1oRrhit
Oo2akLvW+kXO/qWMLJitZVE6uY/L85Fm26KiWBmU+qlkHrVah2yrnD+5lMBm7Jx5
+IGAz8oHigiJ0+lsgRgZT2M3S7oj5ZARBCMT+AcTioI4V7aON9G2VdVpRfGtH9WM
hJZIRtCWlFFothWAfepSXyoVei7tzDlUxNlbFmOInryoEotm2J3Ai9IQXzus52Fs
j8wPoe9y1qu2mUZwMoEtSAYC6ZHNITsbs6ah20hhyyG0AYrUhK2jP1+eZF9Ei6jK
2KdrD2Ie37NbrT5EroWqHlNtiipSdZ9fpG0Fm/XfnpRZUam2YFGzST9B21eWPP+A
YFl88z3oUy/b6ClFXQoEhCokuZfsXM2PrUJOyFPRRnCowP3rrYJ/eQJXQo++qIXz
3ZnVJpBKSqoUfTR9JMUJ23ZCAt81FWlt3UzZ6gnfFbk/c1jyoJ0rALw+bvJi05XO
YqdVEtmd8pPrzDNHvo/dCxoNItswypR9im7yJlnLA6kQdOtTGhS1GhrCHh9oklxp
qk/X4OHXBJEORpR4H5xU3ENEx47hy0c3X+NJhBzV/PYgpJ1Kfv4GI3+7e7ULo22w
aByDLxxO1hJ28m0GOq4QdwwBbeEPHttD9PdS6pLOu6uM8UcVPyKE3WrupqNsJ5ge
saWsjzCR6cI+EyEW3AdxwuaaCjQZnM7sOXZG9QVEuo7KSIBC8pdW/fKeoY5z7HOG
cceERt9wX5Hehl/vbzP1kQ8EKkvfRA/amT5Pj788gZuHyEzrOUNjMJ53w+d9wUVH
j/Ozl66FQFPzbZ+1gmVE84xhYrXsR9WCKCPoT4Hsrcv9aD5M15TTrK1myjupFhIR
fZhmq9J76fip7bP6wagrr/7klGSJVXO1UTvoy2q/UNPEeu/bwKoZTki6sOAWPH1R
WA3h1pC+Y4w10xZNqC9KtSvh5CeIWjVTbHamjDFBM2/dnzOo8HSJsqG4+yTNFC81
9pe3DVtFuMcjcnM3mn7bvhzQM0RYnbOfaVgXEptughH7vYcFiOm7TemmqbSW9oIs
CUfZz+ft7pK+TJykTrPktjzOAR3dSO7vJ+ZqdEsK74VkGUJ/WxYFMDxD38qB13vf
Q1IVvaoHCRcR+KPDzxDy8B+s+AsAglJUUzbpiEgkXFPMNTSq05FtotrOlzc01upr
DFs7qkbc/Vn419htLzpS+c/x1X2rEtJc665E0T0Tuoqz/ErTNlSJGagD7Ek1y35x
2zooePEgzJyrLgPkalLiryHtaelKwLb9uHdWfUYngElEa2PLlCT+Ea3RM5xGEM+l
qERyl0hp+A2R1orhm4m/cdLislmrjkK6+C0tcG9zQxr7F0Tkh7Bt3SKRpnUJkX48
JChM1XcZuJz5LNCs6lut7yOKOxAn6LLFhEm7MAj2WIk9TZUKylk/Pm35AuJzPAXK
2lfpjxezx3qIMbP6yALD9uD1EBnBu12bddlDMJFJHluwaFKPSQXV83MH/yBwLdW+
Y0yFhQ67ELfmS/n2LKHsHGzOWbSZjWbz0hlMfi08ADmt6RNuYXobaGpWbMbpDmMw
wGd8AaFXw0FLj4+6+Rjh1nCnt5WZxruiwNWrYMGc42zXzjxUofpnj8GmfXWt2rnp
MxQMjW6mLJnpPPiY96ARq37JunGc1TRBJOXsQ/kqKwfDimnuF1kubrs1/9dG+2HZ
kMVU1OzG4gLzx+C2kVOhtQoQ/vruQehuvZ74G8LxeMoM0UIJ81v8LjOEpdRpxISP
webiNLHw9Osr0Z+iAFl/Jzk2axlqf+pr9eK00+OcAvizjeGJLaL0qypo36JOAwbN
Z+QokCQ+fxXtLS8RWsCZopLuNbf/LJ1DDRDwOokFPhFojv4vauGw9qxaHYP7vF0Y
2vlulh6UPuHWDOPzOoiYAZMDApPjhFrYcAbNaZ5cblpp5anXX6n9SD55mGADBTdY
N127kKGeM0PAYyWjBymjstRuWo8bcP8rqwk+5bgVSUS0JsBStLmqLU3KVJr/E8NK
qbX3c88HnROhRIMeQ4yM5iqvzaQnmDh5DVt4PM8q7ZeB/hm3hiEctcO1eti0Ghnm
Z0hubd2pa7IsPTI+o619oTfgrfxk4ZonFmjmQFauxcNRCNxvk+Vdbq3QrhpAG52k
+5qntf6JtVjd5ErG8TYYQkhHdA3OT6Eb1VCLupoKXbTDMpXKiSa/g6dpYMbX/ntX
MipPaOnEcNffPRAn4xAGZmyDuK8jcg8nmHhJ7q4bXvJm/AtVbU9E9R0CNORLUf2C
omYkrxRTp7WCE+7oGEQovsh8inwHx/xzY8g3lmscJRIpwUaaNDOQ0eWVrLwOEhgR
fZN3kxck4WvvAt1tnf7LiC0QVHH75SAwz7h8+P4zLHLf220OejD0uXmr8DxcrwaT
4ClM+8acl7x5c+oyCXg6hoQRhftrwVa5JKrTgoj3zDQXA2OFFvtOn9WwYllgUzO5
+Q922CUzb5FCJsvliU4HG5tgKAU34Nqi+Kk6JIorBfWTYHzMICGTy+1yz/v2HPyU
Ki6xF18lgKOQLJlniAzpg6p2p8zZywFdJSXeNBCoCAToefiOTjiOclK4OJt+mepr
N7ACOdKHAOK3vmUGxv6Zrv1LN70kH8btWV12O0+DWzsiJHpcN0k8yBIRWJ1mJIln
pupZUlznnvdtXmvhdjUWhRursS6KrQ3rfkZ2FIFaGEnfAfuej7S0rlQBHn5j7VJs
zYYwiGkrl7TCGGNZnP/UAD22mlgoFT5hXcup7AVacVLAs0/10pmgT+KmXNPxdCPy
HA8iDTNu+vKSQ9/uipz4X0mlch/lLfkI0lWZivkF1gPKTlVz7ZstFl+UV4Wm0BMW
dHDqmCcRmZaLEyecEWio+PJTownz3Q3ofSlEY6zaL9v2+CKsOd8pZVzFXDgu2POo
8eAhJicOwwJ4o4X+2sLMvUOp6sGQBEM09eeXGfOds8q6Rmr51QLRmIXeHyME22vC
Fwu+3sB8zr8r8fdjwuQaz4O8+tfwf1tC+fUcg7H9C+OU2Aazg0ibLSdHk6gDNNOf
HS3GM0LS9L8OHJQX9qUMjZKJuznu+cBT2pNiJx0dem3GPFhjHueWFBVBDJdrJeaY
FhzLzgk8Vhx3baq/yqArQ2UnPWOMUPvGuD7/kWB72r+M3qvjEuHZQzNzxNGPQNFN
QXsfBIYl1Grk2u5oSPbr7uYxJVh5ZvjoDMaUw9WReLVNvniIukttE1MpEOhA+MLB
G9668vDp+q1Ftr84rzZZV5xuw8YcHl0Sc6gqsjoZVjKXn059Vsgis20ACGP0rpP8
hSXMuAgIvONVcPzA1tD+ggFG9EgCsuiVVilJn7Ni5wHFH9HXN04oE/LIuEBA8gQq
7SP6XmaO881FEk5qmTzdPRTLvVPielsuz/m7iJs6P+Ij5JWC4T6wbB3eVx6DCGwV
SJLLHMgS/2diRytYBHy+J+CUi5yOV3Mat6DXf3yMruCy4/2lV0NQVTZUA/h7VYgz
d+Tan+rIuqhgRDlFX+ManoxTmysyCF4mL7QjAEfse0ukeb1HtfIeVeY3r22saX4s
XXXYWVU7qHTz/SqVmXu5SPWrawAH0pR2lLGwkW87CtVkvRRT2dnCe/zcz7EiOOzL
2s/N451Chw9UB7CR//H6aHL90EzIxRedeIdlkKI0AgVmi7zat/Hh8Z1G2xr8nH44
Bf1u6uSYHNF7rpZhiV33FWlNpKw5hxDzOm8JGeRPJVj0tC4esrWXzfbUdBcpub4B
6N/XhCLAjt2DAhP0oylqYd5EoH20Zz9Kvb4qCHwaOdcSLUW8xD8UUXSRbmd31eaw
N0OTu+GMuacplmlFMRKgfWmuq6ciuVGsvt80jfxWWaiSJc7qWFxbqsIxLYaLCTQF
lHnR03FJPeDWyouOJ60ZHln4aSNfjJVJ1Jzma25w/o03ETjLS7/WM+03cYEzLJ0H
sLRo/8fHHUfPs9v86Tx/m/LToMH8vpWGbzwIoxGPw6n1pTPWUnjmW/FTx6UIkQlg
1DVpBIU8pO1JiXVedd4S2n/kJs0G35wY8BmJNry8ZR9jNxFxN0h6UA53GnQ9iz6S
652/pJ+nM8AefeWHvjSpFATEUW21U4Iq/knXkUQMx+SQDENLJr6rar1p8ukz+fSj
qpeXbVIdayTnNc55lGi5iWdLBhQ4lpLHwwAVxFd0rM6VtXarriXSHXvoqZZFOAY2
WeFkKoPoowlFkouwt1rIecbq7vbOKJZW+lpHPsUSM8liv6gT+VcrzXxVJRLQxJYc
F/G8lnfE/a2mr3sReM41d/NyEJTelxxu45P5XyeNO+YmpSpuaaUeqE3IeLl2Qm0/
w8j1ZNiKku4cIQ1vx+H7ExWhELjtPhUn1zVEuM2maaDAEurSokFwKibyJqxMx5Jc
8s4Dwyqg0guyJGfUBypANbnUOTR9Buzm6Y/oau45pPtKkuPvshrQ4KuQzmV27c8B
OeradBOV/GwZ37zqzW1pPfFltwaSKLXI28ngSGhGpLpjepoQjFbB6JteMGB+kZVQ
ILV0NOKXchNImJse7F+LSCX97aMJx+nUlpFZL9sqDmGktKDPrkf9cHzAXXoKvMA7
t8Beu+fnCAJ90Mw3/30Cn7S2Nz1goFiQGI62h62S/rLHYKnu/P6amfa3RBmR5ibf
i41DXWIV8jpHzTJbyexlZavU4kLjxZ2debi/NIp94Vb93Y7HZAxzYAryV4Kdm1k8
gWUJAKPRwGqg1NAPEqYKf2lcCCYQNcZ4zrctNFbWjnhSB9C87EqcJErfrhrdjIh4
/2KSqJNXDlj+/Caz2qp6Wy9ONCJ12lNTX2gVMmqlrZ+lhnqwTg72AOO1SBqEPM/9
TkJc4/opMViW9JzZx76OpviygciX9rwKjl1B3IX5YiTGILZ9ruG9BSTb/o83kKGU
xPyRaJ2HKKGnl6UikSK/PW/y71OedSHKvyFMadJwIGpZIH2aRdrpacnknaVtXl6x
Jhb62Y8XwkKMeqPJBLhaZus1iz5unL+QArRl3tZA6xMBBMzQUJsL2qkE6U5ljdmj
GeXHvwFxev8IhOiNHyWNqLgYBfobYwfc7/TyWt5RTg1pEzSuFeQZkyr/h1q34oXS
4K94Cn2kSvfiS8xasqmqKwzodaLyG+l3Nw5IFlu2Sy8GoKJ7Lq2zDBRrPUjD+cFb
Leti/uTBoc8dqzfcdINMRVkHLOBtXmevr5RfHSKDe+gXYCxHCJyBMILZFGg692nq
YEnfC78Y0ZXhTh5CcWQNYfDV2xQNh+edTNwUUDNbn1zmCPuTdQKQXfB1l7bXxTZn
nIbedFMRcEM2dqKyjXSAskqqRoZS5/quKuKKSc1LgsRv3R6T5P7Di30kBoO8IqwI
8tFSv0+ALvmRUFeB1KYb19aetJ6XGp7uX99sPdC62EyzPb82K1Aw8OY/cmXKo7fU
riRNqn/zMpA+l6hVcQ4QJ6ICpKCt5xBD3K9nEYauSfmM0I14q6Dzh0CUhY0Ng9aS
G2sMGeoa4Vnp+dSVZmd3dUaX2tBg/XSFUyiwYu6YFZYLFPJtnXUKCDgLVFRwHnbg
ZNLgYeADANTlPcqbB1b227TmzF86SisnlEQ8QbhA7JJq+EMbbGrTWUMmmoiuW1Qm
7VjTsGYfCDvmQiUX7Vd4iE2VNVg0E2hGxN0twBolFb1EDQGa0cU+XJ7uEbTlbbcP
3haEGBwJOT4Ke6Sk4sqm3nfYjImHnMZNAP5pdhyja1n61qB6crMq+WluolMfskZT
TNtq57KUpDdb/DKcgCMdOQ8W90rskAv0okd0LU+YodvKJzfToJ1HhO7PWdA5A7h8
CY54zXUIFLIyFIukScNMjkEYTviH0MwGk/eWa+wIF2RXDuo0e+nWlUNNjkmTK/70
fwPTEXGmFuQJCfBHjQeL2GycrH0M6lvEOYkVC7ucChcO3MNNSkF52h0dJihZb6Ab
RCf2TGz95iFdFliT47PnL0o6HPwbM+asUD/HXpq2SMIJA2PDq2Z4PXfsUQAGxdzh
q1oW0Mr4ZCKXCpb1kwlgnlfF3/NHrRHJ/IjjPqOQqR+qwm1myIssr86PaXJShHxo
tgT3OKqXcJbcpTsSYKsvhnlN2+Ao7qRRCyLsj86Ningc/kMu6l0XXwoNpP6hXKvw
i3CZ4qhQ8+3SOvBCz7OGzxJQqECWfDrTlTYjDIsfu6/qw9qVzuMUaYXS+2Ypv5vd
TfJnerg+aYb7OGmete3a/ONrXa1IGnvGTkoO/aLKEOQY6KyWKw5/Qv+LgsKGwpDo
w7HqoRVFtSpLkFkJaPWg/QRRsTZ8gp23ELAG4QgGKR+6Qd8u0RQrmk6KxIcyrgCS
alUNlJafnqZ9aSaXW0twGCCS1A6i/zo9mZQCSt0UvJhfxd3iSllzlkg9MDG4kKlt
2j3RKT9NIf/nozZvInYx0UrHNzp6APOLqOJN/MsWFd7ZvA6ukeKvQZEDCOuTf07p
ob0wHGb42MgyxlZ857o92yw2IXN/dnLob+cUJAo9wOLLFE0DUOaIYB9nQkvcakDb
HHSzo40nHCu/3/O6+d7xi7dy/O1763/D7ERk1kolRZylHsPs8zZ6ghzC0OQM60xQ
/IhunotaASFkcMGyg5FiYmlrUutzY+UyO2sRMKqOUfKPrddoiWw+BGx10SUEdxFU
ZEwV1OydJatidID974hU2+KsZip2S7gDt2uqawc15PUjEa98OJ7cdawa4RHyYfd7
+0JpcFXUiETfwq/B44gnQJDzFCmUlp+wGJe7IePJzDceEDJS+WqJDHZRkvnyfUBd
r5GV02TqD7lJwOi5wZTCHHLrSHZibgeqeyQjmzMw/OfgfEg9rVBtEOM/YRjbApEC
DZHTY1jww95E9e5gnKQy0Zy2pZEhbSH5dFB9fzvbwT6AApuKC7lZy1AQ7xfIK7o3
k1m4/7mgq2zVxmDY9AZfoJ1HU0NL6E7SI18S4gWdEVHKBq5Yyr1VmgMAemUp3WKm
V+p0tIIAysLl9Sv6+RvGJWyIT6iNHTj+myMvNZbCCWqTmmCvzk8UOktHK06mufEq
xhf2SZLIM0gxvK2IyUbcu0HJeprFNlCzl2MYKrQHFaZQtCMhuJaqyNFLnGqqpAfA
6LuJAC0qbUu1fEOxpU/NCc7zCFfbe4781s7JmxlKBrt8usAlSAKtmErGmNMcEWXl
dylmbAodNCSpk9giUjpYb6B0B+znlPhEHm3enbiIqjfsXK7RhkF9QXwHEZ22QbPX
fyF0T63Mk61TqWFhFQhZJKOpSd6Cc9yrCUlEIVaH9HBQkAmaltu7s9UneDzbawoR
hWmuUE4pwxB1MjC7Se5nCzJLqqKPep7ZcrQnM4vpBxHsxcZHW4kbgY0WDWdDZ8MX
XmQm+BJIc5TNWJ2QbrFPsAxHOYppnb7AKEqQX2cSu6ZnklEJpJrQnkl7QZK5rPsy
GEvOlFbt5SqI9Lfo+zchYm98Kpnk7VJgiwhRR2N7Yi5hdi1i8z+AbQAIrdHslTq7
S3x1JtKaGP9YI4BF9a6b3O60J/rehZEDXM9g8oGk8mN1HtMmphrM/c3feFB4E3Ya
JtjYOvNg9aKDeqSvQ9tqnpaRFa/j+oS4+UUnG3j0Oejvw1iFFV4+W9GaTmtQsH4y
bj6qso+ehAmP+n4NCHYj8RnTmiE9f1vQa4yCJJBxRw/Q1/ODQnf6wrIri5QDrZ5A
LMCkkTiRW3ZyV9rBYfmA2EQFk+ir0LLgu+m85ovCm7mEss6SVc8RyXkvJUo31cMj
IECImoR4lLVEvxLQ9Fy3L9awi5zFesYDXR/BrdEtFpslD0D5tp6ZudpuSItzeM2b
tbhsPD6+Qyp08Ff3uefUnHyZ87cUbwfOdeg4aEZLRCfGusmyomz/9V7QLkjfQqY9
KDocsGlNewCmoUS5ewHxSfNSmXz17KXVqPy2uvxXBo4rcULoiCtBJqxaA8B3cQXK
fv6IriTO7/m3Qwr+2T8iewwY3Dvek9WAIT6oQ4YMex3NZgPnYLr6xuguPq6U2uIa
sjz7EE77Yia4h0EfNPacnyqkzb5i2S90jwvcQPeR06dKpvMYTvXeGthMA2ghZr5L
t4U4O60FU1nB7COZRtWfkq+1g5I2796u9eVVgXv/a70LQv283gAbQaZUF+oilCYj
G2+iUUWN83o6rwk3/qSgbudrW0hNpwmvacUpFP5+f8H2CcdoFgv3kzrXdke6LthV
QNPmF5QvaHkYJN8euItG95TXWhytTjiIZntxKlYScyfkp+vR2gI9fbrfTt/9/eGS
Z5f11kdYCkdtamza5SUCVIg4UVWGlb/I5IuPOOGRcvVObN1D1r/K64Tfofy4+mJS
rMmACvYx45iJeE47mtWubcadKFiOIgtfKESyiMAv5XE3fAl6ZAz2hWLCf7WN3Otk
127XSMvHLw/zpif6Tttxq2JOIp/AMkjrhidgoYImGHGiHU4aJBHzxTRtgSU9CAOc
IYC358EXYYazfYp2BNHY4CLDHRI618hxQVHNvqdHcDEv+KSMFW/ZEQsjWsTXww1J
z3pM+M0P+4cv2C4tufTYgfHXadeZnZlZh1R4+Yc8b1xUfj1027c7llJycXp7nOLe
b4Xa+7yl/ghWpaq3PluGp73KRb4GJB3RHPyEKz2J3Lm4VdAq5Nqfkbkjs2i02J2y
V/ZXpLw1eEA/4In21OTVFD5mFn6qU/+GBbMfbkF2trj1jrRbRBCTRC+jslOZx5Bh
edZaFskDUi7MdVUhDeHMZbDFaR9Xc7LmZm+DuambeKPM0taLZebtRzPqD4fh66vP
cP64LN3QJQEeXv7LtelfJq74U+vPKjc1CaS/9StGDC7GdC3yHaEkmzsOscxUZoBl
QBlXShN8oWrYyvprUGoGCGM3Gey6rtDTOsgdIlY+D+U05mwbpKbqrb4QcTNRm5UV
v7iEVOQDVdHAeck1+J9WfhejogD1nDaSVLH4Dp1HxWtjws/+uXrC7e3dKFuWZ38w
AgNqQXkfb3KJ0Gkn2C20z8bkULgsKS0i9imjXF2lP1d77S0XuraGlWaoCQN1htQq
qxi2bt1mWtMx15bFcsd+cruSF0ypx9DR7j0wkXfm4rgI16vayrl0U7bU1EdRqvFp
3/Mnt+I5drRz3miJvs9OAnomrfCs9mjQ3oX2weCMjhso/0AcZNHSG/0oXZanMc+2
pm+OKxLFPWsG6xtKItE0BsiHfYglVJQDSOx+OrtkoftA2FBnbQccOguPWgw9YNtc
caHTyT/zFLCKYcYSmyflWUbMmlGtWmUTEDPuRkJnixktHrHZ5L3Paa6iCVlJFVpF
38WctY6ak3BqK2eqlHR8i/gvF+Ia7V56tDqQS/dbxLeNGS2CT0FBMdGSPfQuqd8o
BpUtWOi4+ZfAV2TrHjVonrl/Iz7LN+etHAd1eSdy0JqsCDRBIA04l5Th5yDN72vL
DGCWjY9IJmvGFuOmLTi0yoMDTxz6JAeH9AbyNVTaeHuRhXKeWGNq+CB3EJjlqCEj
v2jbObR2xzQw+QgHLgV7afg4MLQSDK7M8Cpq/kD0iUCs4nywQGH+WjLFIrawrzFo
W83dN6iofKzEjE5R2UUKyfkCBfBVLLgZQ5qd68Gilf2VsNKMbi488Ozf65nG+zDl
JcMnKr97dbMPXWd6Fv0P4n5wk4dorsalCb9i4YYA7W/mch3q63AEtSyAXvkP8f7A
hK9O3nVNuMMNwGM/q24VekcpnaB6Z1TKKLmcLiyC1qO+wLH6IW9C7Udxky7ZyGdj
aiC3rQfhI91FnJwN6Om+4v6hSf1F31I0KUgPfJckB9ud+2+XJfEgbFt0yrwWcDeZ
czEEMILbxKpC65X7JMejbtLpmI3uYqHgutne6JvSaQ4+A/MH577pjbS6ascORILm
i5K6qVOoVZW5lw7A2VQnrsLfbMYhM/yz5PlIUiUAK9en1ARL+hZ2+cUMVS52biFQ
sUFqaHDytlSNngO0W9miN54t7s+GUWkYxQTReyBJnxeoPlnso4Sjqv/ZzP3cBNPI
w1Il8qKF7Nh9yBVKGFqgK2yfA539e6cTaM0ul8jN5yMnxYnVASBgUa7OY0ES+kuo
my92qXaYviy/I/0FoB63+jN56E1tmP4DHzXymTEVyiT6QH1ziHtV9Mf2r+ep6v+N
hhaj8SrOkGoPHcUZ/UGv980qkZK54nBmEEqf2L/vku73eAIcWDzvYxd48x2WWk4/
eoeZ8Hy2f1is9SaKGQ2aaFMFf9EQe/jymBgPwzP1KHfdKMqd5iBPvJwYQyW8TLky
dNwaFeLpQyeLjCMuOEiwUVq+AokC5MJljh3gJBu5EuNHs173Tl7/ybTJFV/hQrOw
3Dr+GYxyzM3l8ZnemAUmgHdXfw4vl1FVPndzXhvOkwpbn+3Lbgb8YdUPz9PQrZ0r
KVbi3zSdPm/kDEDrIdHERlTmpkhNpf9xshIiFkX22JQYgFaCm6jAzpz/bRxeTQ2j
vwbirxnUQTAcA+K2uq+rIifpZP/5zuex9pv2W6W0Ig5FM8tU8HsqllKvYXU9RLzh
f7zy64Ts39Hx4rnxzKGVUgzv3XCF2yCf9VqkBcWb5kYN4GTVijHoW9qvIiA7Ld4c
4hXlQh2uvtdKWahpQKJC1P53b90B+5aw2yX7Gr8bdoXLHlRiviZwbG2EN0ndnsf0
DW37+mMCsS9tpU41dtRk5552q4iopWO6r7Ml6P60UdQ4fa8OsytOfhjcNpgV9VhB
OMfCyfVZudWuczOogJbstrNoduLY29TYVBIzguD2+GvMoeZd9oYxnk4QtQt5CTTW
44KqJ+TyRqZtuCZ3Pc330Hhl4FFOFK4OyoH/1/0ZfMxl+0wSzB1Z0yPYK+F6W/R6
2c0Q2SMoa+Td7BJwO64WZ2e/H6WbM4UMW9SfJ7Ya1x9D7geGleU9tAMi6TvHZnWz
CqzoCdFYFLd7NX3YTEEpPKLSoYd9z1t4qr0jp/cTH47GVUa6JhJpdCMz4keNc67f
rA/4L9uwaEfuUtXx+9YsZtxCw/FMsHdFRr393SKxglvJ3ihSbkI/e+VXaU+iReDV
S5UYL7N/lG9xXrAdnycr7uiIuPbcCnpfdeSNJ+TcApLZwcWUErMNqvTL/TPTL9kQ
89XlAwEAjf2rAPyEYBhonkSgHDQRFd1cQWH0zNcdiFdBrd6QwCdkDHYXzY8DCRRq
O0jKWxGtjZ8iy5H9XNQKo+OEpWkbUaqt64QbFGkxaWtVfbD2PYix7MyXOqPy/LrP
4eQyrWqu6qfP9cNB57xWZHHjtoKolyeReGw3CMB4dKaxwAl/xmhC+jOZIZtYxSUZ
1WrsOkEcGWeOuPsPA1jHnj1z6OgTNl0lA49tsNxtWEoLRXOpHwVcaUEKz11MiNF9
TTPmrvIQuglIqjbioaScxp3Iy9JbBTwaLRvonAWv3WsQqWIcVNHt8+mJRV89tKWJ
eC8QlvaFiDAdb3o7Lm0M5zGhdo3CxBuG7ym1Ng+WQHqmvuJ7UahlDeufqPDVE4TS
NsJYTXPd8Osh2oh47g0ty92wW/3JqUAH0NVN5YMG7g6wT+iZmM+87jdWOSvRZgAe
05Ca6MBJ03paIhhp9vyaLh1R6aBGicZY2eHtEQ4oR7bqfAUYLRF3LvSD5/mfnN/7
x7YKYhdMZJsEtm5fDLHn5bqFYM1s6FtUQ2ScbbmjSd5MdZrVKA6vVl+bJjT8mdNi
y1Rnd5dfhxJwl8mctzRiyg0p1YBPeCZgSHSTRmdk8prUMi/oCjSsBFEk59l1jUnu
FnFO+SnxZPsZni61Ew9JSUS3dImhsN/gFlVBxoIdygMxqEurWgECD0prJrO5n7/2
AwEkmy4kkoxOrznbgqUjSxe25i4Icr3gR1nDRuZ4XtP7Rfx3psxQKHcBEbPA3XAu
Jty3wHEh9sDWyDBAbJevTmqHU0s2/rctgS/NU6CtOITi3YzvAnqH9pWjrWTZoTKt
QIi9/8pwOuQNrSgfAAKq+rQ4Bbfz48CBve1un4jBgTYaEM2CDQHPVUCGCRFM7nhC
eMtWnDrZl3QX9GI0x77B2WjyYHWzPwRu+phUv2pDWeOOuJpumOfbGT94+RJmwrz1
FrA2K1bOL/N86KSmHg81pi90hBsElfpw+boutRN9xxswfm3y5FTKQmhmeoNBrfVx
Qi7p8lVnxMlvGxQYOl3iN0lRf5RHCJIvEA7sTME8ECVWXchFVCO315KnCKB8TkPo
N+mYlPK0t/gSKwYmv/AGc31josMPCpX/E+hSuJv9mQJBVL5aYOt28fS72IbdGM8K
9W9vnDXHsD2B6hbqu4Rz2CbW41FB9aqQ1PpLAM9oX6eqeOdjhbPK/QLYrdNJN3AU
ibuZ4E9ql2Z5mCRC4CRhcm2bxf703EVSER01ifZvmHtaUP+Yw5bLP96rjYpnEKrT
5oXoHinILMFRGK+VFIFYMxHHbh+FT8X6y5xt94COX2luyyoh9c4QZd/Z7+uQ8kFz
9iXO/OTUvtjp9+vxkIrTrMkaMM7VnWZE6V47PU+JHz8P+Y1W/XxLet7565xpSdBp
pCNk9r3NsukZf1qV1MkHnNGVwAmWSSFpoanT8k1Djgi5C+a45fAQ7+H6T0eh1osd
uAxpIlXyjZlcXmUDQgrIRZRZjeOXuJwwmo5Fgrp9vh96+GUahbEXBRL7Ti/r+HyZ
LdIHuO2Clo8OvhG5D7zPp2LShhs7Znkwcp0z/cfWYjL7ee/j9hxc+2zRR4EwUcFH
Pzp38X0bSCSVqSIsPkLCsqraufsmrmww6r8c1Ey4RVaZG3JlTXE24c7iHfSgR3MG
yq/B5sWSzBzS+9CTtKqmelqHJ1Y3KA+zWxyF+qSf/7/dUWenREXrHdKNR4BLBn0C
Xsa5I0EHf2GeNIA3Pg7QxESkdXXbZRT8fMTeJrhXPBNwfnzx+2WbONFiDp+c0xvR
boWJDIVtwxQk+8DDIMz1bDlFVo6rVhNN+J9oelT+04ccwh95ENkicnXdItw7+EhN
mvl6SFt5YLHrPFLTncX2iiS1QPl6G3fV5d2k6OPU0ptwGL/NiWu8k3oNAVHsY4Ic
PMNE7+8v2XbCY1pqcADdxIj+RKe7rJbVvEeyC5/rnllkpk2TR+N7ibo/v/Mg22mv
bkA0C+309KnHq20wNiFl8Kf2ByNNmSXcxHoPS8Ke0LKYC80h1I1ikqt51ePZ+GrZ
cGW8BiniGneE1rUH9mrlfiBYxUEs2eT0cx0IHCiyAueGFoZkCv39Gj8I62dQiHB3
K9E20AC1Jj1Pj03iAGpz8F7XJeB6yKSTDi8kGvj8oUZYy8hT/9GDWFdG3biE882A
497gw0aQ/lHUS98CYiVvMW40zg7nthujv0bpYkxe3ogYWuy+RMvAYu4yxD+LeC0P
KLfDcC9LLL817Npqcb3fckfMzeXkL/zLLZv/Si5DpraxV6E4gKxDogFBDoiyYPOs
hRJxqJH51leMrIUEvnWUaMxSktnyjz1bDLinut4YRHXyEeikx546qjIz3O6XLypr
tSFLZ4FczNU7bk+OvFjhxdjOU/AWsRzjXX4OqD3v3f86fOBLfF4JxH3+mSZGkjGt
NyDht36G56PoAO1lEscQDPwYr8ghziOGJ1z3bjcI9YTKCXllnMBxK70ipRHg2L1u
AUNjF3ziF8FActQ6blcOxJZ8bufKcKRbmwQUHL3WEnL4pFQPgcciEXMq3UYx50VA
Zmj4edpHIf6Ha55aVzPWvUfxTyriCBfL7ycbmSLo134Jf74BpELUIDgk6XXi12qY
y0mhVR1JPcqEcyKJZnrh2bZmuxkq0gF/y68DSqajaBvE1PQVWt//sE53Q0d8Yb5W
8N29+Cw2m1939tLox8s7CBg/2n46wRL1XO6/ImgMFdlevVcZMcd8BvgA3VMKmPF9
ub5O8XISJOKutk2Qphkq2LHwjoGZ00IVtDe1SPuK1B3S2wAnXnlOpTc+vqriJXb5
EgzQ54WjrFzh8uxaTCDiV8A9GKBV+UQ0OH3+pghp/FJpDl+RnHLBeDwzSRvfR8W0
ybCGI+5zZnXU1oyy/Ez6myaove5WFeCEUgiYlLEGTaxN3ULytK+Mal55ppsEQyeE
mcU6/zJzmZnR811dqXFh66yJHR+TB5OWJ6u6f9t7k3xM7x731l31KaFKcX/nOcVf
bU448IHTjAU0kpudl2qRyAmNvsDv2ud8ualJNM7BoDZA5Wtdr1Bc4noNuHPL9S8X
5ddROvRDxo0nAqNVJ8QXJdlAuyKEmyJTk549D+9aUoKGhyafpDXJSoEuaMGT7vcq
MHjPrp3WP0PM4676TvrfBiHOaLKwEobBk6H2oS+T56dxNsVyLgJulJajknruA8IH
Og6SCLuPAk/qsYkwVVML5QqbAqk8MqTjaO550os/5xoslRKYe3LWji1cPqmJ2QLb
QNcbTZY82hITRKsaWwoSUYDadlULe/vISaDujyEaQDnMbJDwSE7hgaerRMv2yg8D
QbsjKC+tckg7wNL/P0aOYDoT4psUx/9tb7zlG3j9yMCohR6cds3uwBFM4n9whTqp
aD4HvSwM6dyEr8OLC805/CAsQ8Fit5blCEUac5RhWPTwyWgJKS4Afhi+eMIU3Bdy
75rulcEs9GkLUWeQ6dnINAuxlY9ZbiVJ1P/wiuNsN/qz4NoCojhGkWSB7Ftk0cUP
6lCmcLGDUtN4ByOem3NKZjVkD1R3fB9xADXhdSBAfkoqxHuhS7Rn8VCJ3ymaxEMQ
MSBsUoqzPjAgKWpw8UO1gkncfwPLYdHkaruB8effwN/6PU4zIGBM7pn/D/dOsEy5
bqSWypk8xJDnRRtnC0an1VpjEnUtosAfszDh05i39fNQ9pmkV1wRyMj1lacc5rM6
FNCK/B4tf/citNR0EN7oualpFnfVV+Z4SIYxA0OUCpaNrP1/OiygLlfJ7mbRGBQ2
oNWvYhHklq9T56DPuiv+VwdhK5PZNgusG6a38vPWCFAoqmWp2z8XtjzYSRjEVUqJ
pXDK0eO7C1aq++ogY36xU4OPWMDk5E7TBiwngUjC60eFbyshcOVdTCPGIjeFIiO3
E0CEanH7RLAZmnWUwcp5z6oKINXaWcflADMy4jzFswwG9EY2/kdY1Nw+s33vzjYE
i5yLPyxqGki52QjKmAMxML6FvgGCP86qrM+qusoG8tsgOpW+hykWcTs9wIbbGDMv
Uj6G48Wcr0qdRua6WmCZPBbBnzHR+ail3HVtumw6UbBkCA+dXUQwaevvSWCX+nNr
ixks8fxBAl3om9DQ7pFiUlxRY2e9wPt+Hu2UXa/tNGYVCkOasp5Bbtt+eWJQUZKA
/rhoT6uf0miXrxlLEpEhTtr0qCMVaPKcS843MTnvFy6/UXU3QRNVGs/hPbZTQxOG
uUbeAeE0uhJ38J0nEX/dNLn6dwyiEDNguxfnP4WLu9e5q0vLl3mV83XVQYOlvOXz
D7NYCEdLL16CHLt6+KYbfw3kvKPHLXeFg9bovpM1adThuxJIXQAEJ+s8fOz4iV4a
x6ETDwQB/C3yQFKY+IxuwjtGUw6epqCfZysADq9h/Y6y90fK/JlbtaKml6wWEjbY
uuYeS2I8kb+xyJmFj1yg128VLdmZAKeUAcIF8Znh/yZFaEBhViZ780BDR3Z9zIv9
fxPWroRFT/uBQPQZMCv1Nh1h5ygvKnJdSrifDfY43EwZvhPDxQs4Z7RSXY/4lesL
XT3t0dxC+Zn53lhjOUtw5gAg1CLObWvjTxVjSq2g+H/K3h2gYAYA9EtYPKfmp+A7
nZMzEBPMZfn4CQPDKJLcgsCRRv9yM3NusObSN+xH4ugy3b3XqZpLS4UOaM3tr6ci
bK4kzFlePXxY7p/WKw4l9lziuqPz+zo9KvXSul1DwMe086osUgzJG7o4wAPipxFZ
VQL7x+MMvNNr1+Sbeia76yu6RHD2fn2TRfA+YDUT9iVJup5SQvXhMKhlTrxbINE5
ufyxVM9WM4e7OsEjDtyfpBfKDWcj6hqLsTKFTccADMnRbxlpp8EhLnRyHPVcmR79
+MTCOMZsnoHYNY7bUK7dMqtGfQFuhKRDsPTJwn0h1F9d2oHnniKtwrFmXrLvGqyI
x4zNlS8RFtjRPu6rv/6p4swcId+pPNWN1YOTC/gtc0nBCvprwacNvkrF/mtZ3wmf
ks3U357QA/A9DcjxbKFoQJCkbj2fLLd/BHzuVTL5USG8jHmc+546Cyp3gDeMjhrA
0wHGA6f0FaqGPTbr897Hf058KdnRO+5v2C8tom1u0Ecmp9uGXgdB9Cz08b4aCUvL
5vTrvx0Ot/s3Gkl0wHkXAggimR47M0S9ZciCbyxBM9lMNbdsemE6LRM+D7pa0cMr
ybpvy06ELo9P9hB8Vm+LjbfANyBVpqnSR1x/ZfFEfuA6YsU+l1pYq64kgs5CMLDE
w1oOMTF35CGCqFettsJB3wXMyh/ziBQkxLH8GKXbSlkV7f9bBK04eRuMOSNnv9p3
wS66HU4IrFs3u/je9n3igVoVjHBl0iQ7M7PsENgk7xEIEScCxekyZdfkwRNyLf8D
6eb21muzuyfMqo5EXYN7sWgrKSPG5Vj1shFt69KbI7+NBkof8dDPKxYJJ4oqjBIJ
qwd6JthbcxJ//JbXvaRkzRxO4xVPtpjQgJK5VT9WgYWpWaKoYDNd0+X7JQxhDK7N
BEW46cPLqUuuVBwIxBbef78KIU99JfUMSaWt+BfNr67Y1wwxkbMMZOoV/+uXIeXA
/wmh4Oa5GpGPhnURNg9J0FXtBG0XcgW5hbU0AZyva8hNCkdFU/rfxDmmPRa6q2n1
dzrlXxnvF48KLscsMvRQJOSfFTf9xkb7T5tXqqOXx3T+aoXuYFY1NfjsAKU1LyDn
DGDRjaheW/TtAwXuo5tvZuSwb8J+fVTn0k8MUj1aIUkw7Y5oXf8VMgQPWWcYkIKG
9lhAnBSLv12AFJ1y0CqVbDUWzjFEzScKSqYc/ze2g8T5ne3qDTUeF2e7+hRNFUbA
bo8UTYcZgf1jJWQZb4Zq3fBQTXLdTqhCoNd3Fygz10/hnhRnSPIZfVr0jAugTzo5
I80YTuXoqUmU5HFXkdzX+XW1phBreRSlXFntdjFlf+Qxwtx/3RpnW+4PhJo+Vq2J
kTnHQWsCFDcb4AlgP/9rECaYE2y2CgZ4YmJrntuqvhWiz/MNld6958AB4z5aWJJs
3fxIPfO0UHeaaavg087CsqiwJgG/LXGuwKYqMe+F88y/4m/aqowY13PQMVxPb0v+
f50v8Jh/KDNCRvFKFmppdQkcvTbhwhxlAlR9T4WOjx1KfXaPm4j1k2NWZOOkxJns
INGHSuSDQoLifyBcqkXBB620Qi/NmRcuJ1Os+LmIWgYRXjHWy7DChmsXC+/Ug9pd
xN7fcYv2JP58T884uwLsCUO20rVkKv1/N1D7x+KlbhScvAaclprfall6bjlujzpF
of0GHdvnULPbUVX5JMYv3/9ttWF9H3AKuuxHlaRXjjyY4rpkmtjddyoV6kCH3DW/
9Bqs6AdWV3Kr6MWmYNl6yrbi1fh+63XBZVJGvV+A0uuU7jprO5u5AOVii8NUAsDS
MYv7FzuO+0KPtS5SqeSerFcpyJJ6yv8sf+Wykr4XA6HB6iDG66SW3K06fPCE6ugj
dTZAG2GMyg6gkSfFGfyws/CAdi9Be5mcHAiIFEo7yTYbHwm+w+47mUQL+HJ0T8Q2
N0RXe1Vwby48ytrM4Y2mljmXTiplLONb8OFaK3csoOUnYtvgDwsTignNH0KY7rV5
CZFdgR805AYAGFBpDX/bcxXiedPVjZveU7cDkbRWVETw3UwDBbFrhZdX1QopTzrv
g2zJPxkLH2Inzi0kMLgdJaK6gp4NXpfy2cS4f+hE71dTWQWxWie3KsSWc/9a0Zez
vRUit9l+8ZNF1lVdmX16hE3WsQGqxpk8yBdos+1H/PuNSqBe/62mq58sjQVI/enk
pz/whq1ya+dwR48xRuT9p9iGUDcuOsS+Y1/CeqK08jWeiBfn2ocfw4Wz7k9Ay+RJ
gGc+a+Ml2hOUwz22uhlJ8Belf9us/WedS1a0j/NIszBLvOj47gzwIuTlmjD1L0VA
szA9xciDXkLAHdGOvpwbumFy9zboorZk7r5+JQOW2skZSE0kCH8+O5w4B+IORC4E
d0YjHdVkgo3cPXtG3UfJiomVpEvT4DXiu2QVEvgGZGlLvi68IVEmAzRqszfqH0vM
U6DHVml0ovw6WWc+4winxCjJJKKpkFIpwAwb1jbhbRcO2jsSvCEctNA/e2kAbDf/
/Cc9sL0ozxEGrysfRyHnYrFA0nIbNaoQueIgTbwPd6MXOlwVeGZXAPQAknc2lK1Y
F8yNIDXrm+Vz/qHViGaDp0iV/m/CYXOYWslnX1YsYl+DgeAW1TRqG0PKk/6eJale
97otnmbtrLLoMoOopiA3UGbKCLHIP0ImGdKX0Mx0qgKyqQNSydXjwcrSW3cN97bx
3KVPAynxwz4Ah4uiuPwyDCNYjghvtpBTZQEmazCY3UaN/ixYP8Yaljh1dzfHXaWr
8sboTh3gDvy8PRvT9Ex87trQRQUtlNXpc3iBq/DMIb+tW7IoBpF30GFD4lNh2YX3
C2XzGlue944LlZYT3ZNG+tNbzGdIOkPRSZKcTjXVZ2bi3x2mP0rmgqj7kbrYrCT6
NRqKpnAQ1XRyYgq+JhzgoGV31eDmPoMfxZiRFcQLUBfRb4EBRV5QQopbdCsz2cuJ
c43CGIJVsX95zVXn7Kx9szpgyPGayK4sWqM9G5jK5j3nCxaxZcB8Qrw/vCRktby2
AsF53pTyXiCbz28xxD6F2DyFDSQZd0xNN68qhi1Rw/7F2QFgBiWmWbiqCg4+gKO3
97QMRkyaXgwBMt2DoPHIKocjVYBSgXWSXxjR+xDrVbNt39/cwMULOrwV5u4XEg/W
gJWew7vUucuFltb/aERqELbwNO/6N5//I1ChwP4EWCUwbhGC2YLCGb+Rtqdh8az6
9jzXmSSZ8CQY9IbYKL28MLNI2YcD0g5FezCOMGlPSrH7jt9YobE/EYbn/NZQ+ozL
ClGGoFNQWuYKqeQRSHnMqsj7hgSOB4pwikdwOso5gJY+dZaVm2OG/ABLp+e4iSAL
GkkWEouWA3rCgTuotN9lUIk71VNFFTqHCttcmEy7983yzZlrMp0a592vSIeki6TL
hCp5P/C4NZAW9ElneIpPL7RdacZ8N9YSJl4Cy7UTJsntObEnE3Y5lnwY5WxqBwpD
4ktyKrRQWcGxYgRwcGhG7h/DHv7FfTN+8SmoHh/xwiGacrxsU/lQNxSoN+r6HgBA
KijFyf8qFLxKPKwjVD5Z6+jcYTvGnp15mYwu67GbV+pwV01HayK4JBVuyJbMHZ96
rSOKI/ImlE32xsqqOzTursQMzSdCI6F0tfkwVMcCbFE29C2nl3BfL4V4IECVRC6o
S7LI9DEAh2UWTBUgNWK6vwsuSmICdBd5kxxsOrx8nCDPKRxvY8fyTLtSe7xDVGdv
RWtYulPmO71gGhzQr3A8FN8XuCPTkwTnvnoRTKnqrXK/t4cn8EnyI8rl7Mdjjj7q
aGJverJGelr6LrLb8DjCD848YpU8LcHmY/Wuka5/L5bEscAvJo9LXM9JrzWUuRs4
HYZZHDLV7CXIC5XBq+cGHoUa4Z4tNbxTvyk9HvJIwaD/hyjSgFMqfNSt/vK6t4wO
7pGIjA5HNZBfLC5iXlhqp2CcAINTczuBjR9QUrU6kFVncGRJFABAnkHmiomHZg5W
xB+2Mnz1S2q1fG9CgARzYWGyX0kIOWpJdQRLM0HgsqC2UWuGtxvffXXdlKx4xNqe
by0WQSW8KDd+TEVzTqYQeNpIM/EBoXdvmTBZ9tfYgfcLjeatqXy5X2LXJfyBxC3w
pj/ttk1Dq1RtHSgHJ2FYsYsZN45ITLjXPu5DAQ1mdSG43iP+8SN/gyMUFITc31rA
24dW87tSkgscnX1KiEhXr+MGDFzd94oXHgXhjp6M+o6WItX/KbxEpQxtv46KUgpG
tPBPl3ANYeK+7e2twTZjVvL6KSy7J1QPS58RP9PSAuhDeDFQsfu+jT8gzUzIMvSM
GUS0i/c6FXNUP9Y9OP5fmqAbRRpnCYF0DCappzLK5AdXXcZXLOLtsYKVgdWgIbi+
oHM4zL5tDYMSaCkMWwWBSFHbMDXDu185Ea2EmF6hiMVmLTxKURxjRagvzIcUnUe7
7GFydbhPMglJpzEtdpKgDhLetiWtC6oc/7wERo838VetVDtBxYf9rlcSvIgp5W3l
cT8QCFI8BIGGDu3T85p3z4qoN/nT/RXBVXeQYkUZpVWCy5I+55CuggrMH6MdmnzH
i0coJidQUZ9lZzFMpGWYaQBycP7MBbAQp2YAmuKruYxBLupbVNvB9yzBosjBsgIW
6suEvwVHr9bG4wxHhXPben3qjZVbH3o0iXs12ejXf8tq7SSFrVtNXwm+JzyrqYEK
Sfa+XBKpuM45UF8KHeEr7gM13iP1dQMGzGApajI/yA/8H+zB6fOSHMTb2Sxv2UB2
I+u997iaWDmEdKKopjRQwzKC+juk2wP9TMtIJlziNnS1aY2DNXDp7rFTQwPlw9tl
VjAmjNDYavV6V7gtXaet2yMxgwtEfjqx6nhTuDjh83VRaIR6rfyjO48UrvqJDDWj
BkBGWEB5dMLl/letFeW6xEt6QWeRUXIA6UvtHppzOGQlVNUxubIltfCv8/83D5Q2
zBmP/HVIHOCaMSmayHfAbkbxiWyT3acku+Ahvgow+LHeiQN//ku+OBCYVaWtZaZI
+pq6WuMZs6WQKCH6mWQUIyPfmpR1ontSxs7ELdy2WXupBZ4FDTi7GdeJZRoOWaii
i3Vg47KKKUYgLG2iIyf7yQpU+Ghwuz/VLmQCplf9cRmniMTeoznB9l8ACJhaFueo
igM64UKW7GTGeskNJtzi5SRkEe+CUo+QwEEaChlWPsvzDF68jcYOsOGNueeDMP+5
FIuHnnh3BB4zW58rmqu8Si3LVAjuS74072QcyiahikfUbRZDxF7ASl/gY+NnGLz9
hJ8cfAXsFFYzHWUcZrc6NxID6JqWJenQ5ylGnd2XIb9gEnFU8NDt6920XJzCDxby
etMEZ196JVy8RVMne94bhNl1qgSZRqtZ2wTfdO280HB29WLeBZdzl9cf4PaFsCJ5
8BINz3Oit26+41sOgOZSTT9LwGUieW+ZVjWISrNuSycnlOcyPwl/AWdKTy+Iif0D
V74JjIUiBz71dse6adMq+RiKxOEYUTEvgCS/sIio6GillzUwMEFd4HHZEvg0ZV0k
ir7O6zLoP+ujQM8UVynyxviws/qtZktsOvWV2pqgGs6s8OgQITvygUfkVSSMi//P
rPYAlxZ9IHIM3G3w0bUXDtfQaShyfLJGxaz2nzSP0hbfL4UXFQxmzEpAqgtvOmli
SG5ZeNtpy1mT0UjZ+c1eQu00irg3aXR97tm2FCz0nVm0hwXCIS/dXHPEQSXA4zJN
pIbokEjpYZhLXXbVgSBD/eLpIcsP3TDD1v9iJ7Vs0N3hsDsSNkheYquws89SdyrY
B4SSUowkC9ZWzGxOpfCxeex/2uUWhsdgrJb/IpqTnEgbmRBtKB7iyDAxMNcRKsnF
2lLdQXtVgorm6uUgR7fEnu5/mH38zg+KHy3zZYB8sJMWO0Gl5C1q8W42ss3LhZSS
J4rQ600AeCA53qQkEE6RqpYNXZkhWTBNaYMR72SUH2XEIPu1fP2wy9DTNamJHCSv
xz0W1xJfdNsm2Ryd3k/p44RDk8lt6yBEdc6SRYX5YzxZPPy89di00CpY1EKjUCLt
mNobYvjGnKTaFE/FdOb3ZSRI4rHVDNRQVSgzvKD3ONaLfSnOj+8x+X2PuseDEBWD
pHtrwVtHxM707YEBMu6oLKwcVE4apDESl6bmTql/ZsCOpUBS5jO6jluTSxprv7/9
vImtZamjJxRWXgRsp4XHtlx+glv94KOXdFF9F+U9pBqE+wWSSsp1jMR+2PeRu347
WPu6O8KJpK3inB1tbnfradmed9lDZgHRKPVRT9F7srWWZ3vLvEya7c36sJHBXNQ3
hWEkZR7eOVs+46sg0W9LTHLnb7BJ3EoSd4WWIut0yM+CHOtzMBvH3+D5gqHME8Jt
QANKMsDGKMxEHs2nP7HmkHZlT6XyK3W9+XxsGBkbVQ/WJHgTLsvUTalKZcqFOTWm
YWx8jygK6vIW2TvZYOvLDj2B94KCM1mEN9gAssa+vNU5KQZxVptCspLWyoaOQWmp
O4g60seLZBRIKePM1v3eW00EEDd1wYWyHpzfmEyKla2AqzNEbrDMif0OSCDr64CE
4OxsGU8q5olLm7H81S4+DQEmpZ3+C5MG2qJlfbx1gEezrS9h+COpBDxAcLt29diC
1I7u1XmIhCGQ2VmBz/I0TinFS+I55O7OYs3BF+WpH6cR7j11PIJEAL83bAAJUi0m
Y0TbFjXzzu8nlm31ZtNSQDHa1MgiugEeTELyB5RB0uNE2l2X66e4TuvF82hI7Rzp
aEeSdOD9EtOqvo8WQvQes5WOfk0Fe4kkdP/A6sERtwY7yyw/9f4YOAlBI+d7IwR8
gO2Ohkjwtw1xUXYJauFwX3sAUyVOQr3XGyX/TF2N5DCFswYiVh0tksk9t5FkbYKc
aiv1C1y2j5DLYKChAU+dqZmi4Bj+qSsctoGQy+jq6u2Ula62rKqjch9Wv1aW8gIy
Fn08XlvggghxHwqzaj0BR7fuGgXqIc6QV2lT4Fd9hJVqwHNK/Qm79D2/dYV2VqRq
fcwfmAJrNnIm0ELZBUV/8q+NCLDCfL9clv5fsmoiauEa3NXt7jl8vKEogATM9+fF
Gt9ecX60o83oRUJ4bOP/0hJHK2cXGxQ5Aadg0vfxX8IlyZiSl21xxTsEXFa5MqaM
Do9siN0mAZSPj7aDDGvbFSsEANf4FqXFa27V1mzdRItPHGAvq+oXZaGPGW8/Dsdj
5GjPWdfiDiiefabqXgSSGuOdgqsBILlbe3bDJFz0ljjPiZ3NGKGSsj7DgzfsdSkL
frHsPsa1bDHbhsh6EsY6yDZyyjnD835mLn+yTs48I2D8Xb8p7IrrUUtNijoJEg03
hD/K/mIEY9PreZP9KPGa1qkPZyTrePu+x1NYpoXa5r24DxqF25sn27gglKfs/7vf
7gqTMLHwR6HAs2D9pdkUjB2zidOXxYlwnGipspriktcgNaUAQtaG+2UeHdG7jW8b
d4JRuqZU1xMUmbYpwfx2TMsLKzNhwMzdDIhfgvZfQ59P/EK0TZ9p4t+TIwck9TED
Jp+VbRITBRe4lKtN8mSPSV/bKBFzYaVuuSSqM+pkOibnu2lGOIH6P688ZHkoYVMW
tNcxc9hWEGeZcA5ahz96nDRFTEMp23n/5PIJ53ekYhZbEeGEmO30QtVcgZlYf/dm
ODvha18+grOF4h1665aMANuieprAwYVOniXRQ+N9xHhsuBdy0pzDDyFgAVNAnxK/
N8mKfGh/NhgiLpNYkIxFlCHKcyZDKsnTEX8Ce7QzDPglOWQ8Sn3tuiN4bsI9jfp8
DbIRJ77qX4iah13ye48gqJMXrU0/vF/zpoRrxboSSnjbOpI2TmYC6vaN/FIMHn13
x1idtfh4v+YclnJt1TrKq1gOtljRnZoyrbN9Y0RO1M0Dpks0MqNE9uRpbJsv5Pvg
jG2CLZPonODYX+MEg/lJu3tRUYhSkQur+J9iw0JylXIbRJ0hiwAJtqwsT4HIEb60
HjjBdO48tNAsdt5zJ9P+H90o6xB2u7lVsHgnsCavRM9eM0Kwo72yenTm8AY2L+3E
f4rtjrDi7RYKI7hZPmhfP2MoHbBex8jFjLwApWAEjhPrjbZ7Kb4Nt9GGSYyI6s0k
T9dXaiYnydrKODFqGvyVw10JaRUT6zNbzaN/Vfg0N/HE02V1ZPcwHipqVqMMk75W
QxyIyuY/UbjVSIMUvx3VAmYVa/8zkcpuj6/fuXowdckgI83cgLMggRG+XIuhEONk
HPZiZrFYbI3CafCue4HjyeoBrUTDnFCoGBXtc4jj61WbU9md2wPoR/afbmFiFfV4
WPCS1fwCeozZI39KVuSSLRq47v/FSsb3bzO/lw+oXeCZBkLJdxQaaXeWcyH0lML2
erYN+EhErMS7zF0lRfefZqV1HmKZ1WN2xuJGoePxnbe+tQKaHMRja3vqaSgcUU0p
g7k5ebfxwBjF9H4iJBPiokUVlFI60hD/+0G+00LmgpWLQGZK5xmNC6kT56IpEiim
WN05KewL4rZcss1YnBbRWY/OgLYBUn8C7+RQCGY1jtesVDHWu3eTKkngutso9d9E
zJU7KEZ1x6XvdI/sq6FjxOK1sI65hHwJSKyPTxFbKrrPp/q4mXVD9CFK59JFt42F
3kIWvgqx2L3Pq4Y6zWiZXzOrVZL9ky1qkVmEVGU6SEroZSMN78oYG0bGT1aYyBH8
5XEC8zNcN5pQml/uE5f7s+xK5VW1OvXI1opbz4IIWuRwQO70mSbzpedp3shsmiw9
KR7OsP/82lM+vMUyvdWT8GBG2iW4NFt5ek9cSNgi1XPjYPfaZ2fXpJiFoksziTIf
YW9ujwSWM26xwnkt9ve9GBnDpRbQX2vYpMFQWbViAU11ik49BXM+W0XOoMPdOPYZ
0xAzqznUkp6O7pOtJB8XltQBtjgJyLK7z4xPLJOZTtc6hg2rA46LG/BL3VlxtcwX
JNznJ9SzolXiV+e0/gsurUPQioURGfejwctO2YwGRkY+OCVQugtQo2iNmAUCR0SK
6PDQyHHYJLg0mA56yiiC8heI9WDof4omDSw2V45bKb2ITK1F2DHstzb0lElZJY1v
YLu54ksZbiOQq0cGaqchqm61zZqnaawatJL7ZYlWjA0WPTn35BT5W7Ih83mKWODc
KbPwtw1guwEqM8RovUtZT2e5XnCAY4L8fnWwZ/uBD/Il03x7+tkqvBovgkxzqKfy
2J4ZKpSkKj6QAvIRDjsN87c39ID/6HdJ+P1+u4blbgJrkB0K5lhajHPmeapxDaa/
XAtrkpknZOjWwX+ag+fXd2ZFHMie1TlLHSJrd9XZiFvAG1Wv2AD/hCZYZIxxyql+
8Z10J5IXfYnYQuLOeP05eV4hO/V+q81CXiPUrt4v2ccKmjCDQDQL+IH37RpJ9IoH
wppVpdIi+tcrylpjeA+dXtijFPwygcqMXvu0a5KGaqi2pL17AUuiU/vg1hdkUe5T
5ysvYygNroh0bGKLKnka83MuAmVyntTb+rIaQrFPU1zyZrmCQpwzS+RcOnr897Fz
XlmQJTsZalkEcBYOzMr1zW3OyOCTv6TRjo/bKe6T8RupHIcnnx1+hBMgbHKxFMgu
5s6cNCEtyy2UiPHxXlxBJrsoGGscMWUuOVgkt9jNZMOaHTY3eydJpZOXrhR0G3O2
TUv+UU2WxPGsuib0IqcgpH8bRa1g3Id3dLyfUuFimh/Yqhso3f8/j9Fydds7VMUC
wMistXsxI9dN7iF748dcNv4BYLwovcjyZ/xW8EEImPrIBFIbWIeRweGHGZeKrhEe
NkPEQvNH8nXQtU9RFDbT22hzL/EvDS0ugjxixTvM5OODPRDYS4LiwGdw1jYdNw/c
WRrusqr7i4G793S9FdXhBYQavF7slte6G8gsKLpqAXpkC8ezU9DL20YqgKumaEj9
UmK82ib1oS9SC4hH29qx0MT5iDP5g8p3xfaTNxwY35IyYj0pYnwP4J7ZKRvCBVqa
N1vs0I0CvC2JGAPkABpHpsi7cmGed634ne7UgZBu/yIF45Nxo7gEQkK2XThzqq0Y
razFRGy68CeRoJXc4JjKjSb7bKwtxuskog41yAaCTSQVki8D2dsI7TsoNSZsGFms
irvMowhMKIqSPEBUd3DSL/0BldVylL4QDejxOL3HI/TzYuBDT93IWN96Wub7ja+C
tyBwIoDqHSoQ9XFHJtw5lrIaKOePPtpPUukNfyi6qDlBfncFu6ZlwnISmp1Q2+7G
mulWqMf9L0QzS+GGVD3HkY1jqBGQ+wTGX0oEIGKb/cXWVs52NUgbVDfubro+B/1f
vNpLiG24XpbdOQcMYO1QEF1+5SbVGpWRI1K7LJKbe1ob/z4wDgubN6kxMDiTnCf3
DBgQnTRxasAMmQyJTMPxZvZL146I4R353JSDN+5gWfS1tcKs9BmNTg1wHLQI+JyY
BsrGgn10jCVmeM5OQWZ2TLfiHiNjOziQHZiDqhS3B9dTW56VqbNoQJ/UuLX99m6a
IYmky8KNRIt5s29srLQu56do+HRJ+dFAJZqeEpxqUuhkx+R69LVfzf5AX7qP4oXm
ZxVUiWim0ED1CQorktwhYaVy3rCR2gUZZiUyej9qXPkz0e2+XvYv/DUyugHhrYKj
xaQaQbv2LS84h/9ETK1mHi43lcDMwCDMbyiVLtpq7kOFc6ZNy0JNu2+3Gfm6RAlw
+rm9NleWid3ZuO7wBg1TPIqTqa5Z5xF5jSU5uXpSAUtNN0L3TWP3lZWy4P1qC/UB
JAfvcs2RNguubORO90fdvBj+ZOEKQiZ5E48UWOO+ZtQS4TSjZ6E7A5KPqdrb0OV7
0Zyr1+zJJ8gu9BV/0B8hRzboqHhtf5laBO5JhlIGA/mzaEGf583SCD+tS1HK2la5
afGnxlpr+jkfS7GRRyNcjrjD9fDJ3fs6tunriHctKVFG0O0r+Nctq+yH9o+7Jdh/
UdTWAr/AgcLDoBjzX04vdphn8m3Ck1PZdD+TcTQQGqhO1eZF89IwKA7tl+bZhHDT
k/jrtt2VBCSUwvhIEqWl6U1NJMcCryJUa/KTBjktNqUOdhxK/3KJTDX+ePkT1tTg
0fqCBXQlXlB2+2HCfxbT3wbHqMBu7YVFRSZWT3p8WlyKVLCZODqZybCTKd6Q1Sh8
KD5qdqKnh9J7VYMJb9H8frwEwBXCnDoSTAbND1crmHPGLuWMZOs029Igpe+PmFIF
nCf4IYydBrYZtSjn6USGtexkv0sbJQ+q86POees+c4DmJ4rPNiU7cw1zyh7eMw5G
FI3tch3Sr0+CyEMD5e9G+kwkbF+WDluIP6CGsAEVkZnq8/9hmyoetSW7zwWpNHtY
4pZY49PCRtw0s2gasumd0wVjlfHcN5g5DbQJvZuRPsRz9K/YIEZkIlOOl4t7YG5/
ppVOatySeEjaMFDYLXPFe+7s6F+xtv4gl8Ia8GCIHIHCLMphyGWrM12FEoitWMRt
3arjGGP4+Al/m7Z67FcZDP0c2DgPz1vd57jVX/OHMyr4E1ZA0DhDUWV82NgCTNPt
V/1g2DcCXEaAMcPwnOjqB1M5REdjb3K7PtMhQ/CznOvGJ01tCoiEzBCnAmVjAiMT
KvCgZCWmkAalyOrbtRgfQK1TesfOPD/sy9d0CbQPOfYRnONq2Bs0lfSHeqbF/KM+
01fhLMPkSwA4jIJ7FsX/SNNfVgUQNTxwTyVekfKNqyxD1DC7xIRwScODKVewqaz5
O88FRdp6kXXJ7wvj2HRAdZUuLncXtim20M7B7pe55vkmJGuR780yASwj/rIyZEgZ
uxoKn9lFns09jltXdo4tknM5c5uc0wISz8F2GH2UerF5mtRwh/ybpZErSJCiPzya
E52aQ7sfbxslznX57vBk3W1Logpzu3Cbj8CK+mA8SCUuSg4hZhgfpus7qP/3sy84
pSRKHKRsf7hFD8iCYIjp4T94X5nF49Mza5up8C02yTHrQgSrtnthmgX+Gg6FtZVs
Z564K3m3qxqydBMt0fABF6Ba6sj+z2N6alV8QmG7sL4AoUQosLw352bYF9N56T7V
vBK+YBIAPF6tNBXb/X7Z0pnGzS1ozzg1NHeZbfO/BrlosJd3GpM47nxeACmbof1h
xkOzfs0KTIUbPjS9mcrNrwXmzOcsVSyjI+Le6tozV8Rk8kICi0lxMW6som47+jPg
e4XY/aL2W68UQw6jldN+mqEQ1QyzH3n6Zt5oGXvSl2stHyONGe/LnxmG6itHDnli
DDb8CLiWvwKcAOTGgEDmwfPUvh+GOSk0prrG7PPLXtRPSDKv9wwJFwOHhxKCe57N
NHsN1bLCyhuzFZEra+edJ/OkHI+QS8Sgvqyh9xOkoSjIeWCi21OOpyrbASSdmq5e
KL6GvUCI4FDHcTi1EemiP7Gd9NYvrkb0t0buN06VpmvqX7HB0JqKmAgsfay/1lCl
gG5OMq91viVpqsvRKmG7zmv4QoulIheMAkdgA+d9S7VB5BqQ9VAa2JkCleUlW2EP
D3M4thmhZQD6AfXNbTh0pj8OxyhSmUZVrzB1q7fjCPCnfh3kLBSbRM2DIYlMpMHR
lyqJ1goTJbJXv0zI+DGeVtFlcvtEH+hBhSp0aPa0gkiOYSyK2XXvuJlZHR77ByOo
qUAsDulS2H4JUZ3R6iyDYgsTXTwgWXGMQGD+gkRT3FYQY1drt35Kcn3FgfdOgVaZ
8b0205Lj7UWn5xjLx12YQU/PsaT/JGrFxQ8bh+SE22wM//jDQwP4pPyqlpHp7Gt9
BDueO6qWPlzhAat+ajadxORBc1QX7yVD7Vlq17BGCBn2aZ/DotuaUJk754Wo+Tx3
j0yXFg+pVVKR9tOYzibqqxavmwD45rLvu+eUWtQlThG7xlBINjkR1H+8nSpCGMG3
m6ErqViBj+xYW6dbTOIOqmBNGhlgL+SVDHGJol5YWxW1uap3shNs+NvfqhUKPIr7
5GsDGF9AjEAGp8lFm/2CIViavzp8YIAsFCbqh9LzGpfcKMCfkIM/ZJjZc+b1sJmE
foRN13pymDnSpfZjFBv5V5FUTA0VTqclPHGvL/wwh4pDTbaK+83g8ovPHPoC52dG
uFMgUs1dqgoc30Xi1F7+3p5IPQsBsRndfh5/j/2tLq6p1v90luKypLyfcoyJUZsm
x303FIbBSGlWkXabx0YIDyK2utGtD3Xa30o+BhVJ2wKaRkSDTlsnukx3HDuA4x/A
uHAuOeRH2/vpEUYVI/f1c7vDLnPLVehimxYXGRM+2cAyt3Mp9WbdmZb4M3uvUnZK
iZVNWUPifSnUFCI9syAlv9J8kNlIvmOdl5LFUX1xDL3DT/qhsxTiMkFRanSWWcXq
diNsPcBuvs2OqkZnHngeeeTTPLaLLh1z3XPmno1qr6Rkj7nVVJ3PQJkw5qAiSeSO
a0WYF9rP34okhRyZtGCNiTW3zykRkLosiwh9hqP9nN5kEUdDiSZ3wHfApa9A/X72
XIQYZfYYSmchyzujp/DtkyLUrsH2DTEf+UZ3jUd7zM7zHneccj/ZQy+cNCr1T99F
CcibAYG5yWebU0m2TVynXKg0aQGsWa3z78GUBEBX4IArcP9/tyUaLcZNfyS4v5Go
r/alOW3QZVufqD4HD1lC8QqzOQEYG03Vv2kQD3mqVXHzAP9tJNFmJLfExiZ5E53L
OBzjKARiDvtdd3c/IIpGBnmMiGy7SWp7A9gnc0f+3s2CPAChuLpRRpXf2BSbX/WU
cAb5PQq3BTO1ROlRMKQjsGxGbDO1+PuWnOvnN3b+G8w8vK/Z7YPe6qPOaW6DRPfJ
oTo/T9WHluITorUxzqVHlsD6j7VHJzwMlZcOjYrJ9+FyBaq9/5Jnww5rKFPM8q1D
hXxNWlMINXFjCGqBScXaSj96JFFbj9bo4gythRLQi0p/B+vn4urih9TZlj6guvbP
6YLgLeP7Eii3o9QuOSZYgmGBgxD86qogsfAfCF4+5NwQt24vzqsQ/0DLPq5j6qAJ
2NW++7MQazH/SUyUK4MN94Z3ZThG1eGo/nvml0XUljJdCwslJzsjYk3W9x7E/orG
JElGj0hrtWr0CRUXsuEgxeZHdDvVS5sl/QTRI1uYAW+LxtpjMh1K1yGfYhgLrq26
XURV8mA9axfSUZlEOQ8oFtNRHU5GScTlOxsLHY5VjDC8vJnnuM4hX3bQxkp4f+DJ
bpx07RDXVqAlpyS2zGIwwoc+hkDPqLtDFJQEpzrOrMwYAU09Whj47N1v72hoJ+GQ
FzqDZ6/OKpH4zbWi2hifCUM701SzaXCIJFCev8rGi8fXu9RrDW1MPUxQQoYHtskr
K5rpa2RZOHqTzkkuFFlpyfpzMu6XuHp9TDdjTxccw1fa+P0k5Y58dRj2I96ppn+m
NZRAXDDBmhpGrIlG5LMubWWdkL541oq4mCLQuDNTiruDMr47K7HjRrC2Ii/M0aQp
R6Z6HGIYxPq3e+MP961t0rn+TdKqMgC3kH7P0vBrg1CUve9MudYIlNDxlq5LMGlr
jJGQLI8HP8zBmP6/sRQTGA5BX8WuGFWZWFzR/b8fP2m9wuPcWTo9KUPMgJhlhQPC
/dLVgX6OOjUH0uGw3t1pCDaUQ112HgtdCiEvcvJ/0Ux2vNI6b98VAuBR480zg8W4
h6/I6z7c3K+42jbAFXDpR+tTmvqJoBUDXZcxSnEG3n4P2vBVAj8731W96G1Y8OiH
nbykExSwUjqNyHFsWedKkIGQXXgNERyKQTic3yeuCYMqJ5Q8dm04pzjVtNoxuWEK
lQp4Xz5YWKg+LVAWRM+E4GaBdnzPuzX1VrI9OOC7ehAIpRdB/q6mjirbzWD43+P8
3fcjHYXsMJUHqDNVert4NSYw4Tx2TCnPx8zH/ErrPE3s7VuZAKTs98aFpCpMaR18
QrLG1GlBRM5D6LjLJi8h43IaLCipL0U4qKBkOHjosuN/Zdv/BFRCMgMhhR8YbTdk
+purb/2SNF7ZDCSK0cE8O9yhr01Js7byCsanYWl0rrP/6cvtnfqt12H/zn7wKkYt
pe/7YSvEVWytnrmP1Upn/9BnXCDKNhlf5Z8Wfdm2txnwyciO9dwRiBcVDQa+cccC
tOG3MKuzB5sJAxLNsFHja+9BIDo6CeorwarRlObxukmGsSoLREF5IdQWTJd7nRs8
qlbPqX9Lg8iXGoyAqpNF52JEm1c+kFILxgIKh1qeW8GLJ9uYXNXkckcQV9I+wgN2
vJ9e4kjCgqrzO785sC1yFRIj5FebB8R+RjcrBohhxOpWrU9j3eIkSZDmr/EzOFmd
6/pjQB1mBEdq3SseRrri9p1MFRHEXWgT1uZ9bdIvAzDqGRsRWZoEjrDSi3ufeRyA
ET7e4S/2fcp/DjtAy0Bq7C/qCAR7MRwnSmYtjKvenLyuENyVSFaJ9SxkThglDuPk
H3/scsOWA5qTwpekav/prCbfQxKdSVUp2UmFwNDnDPqNdgDraaCXT6NiJ1965HyX
aMxzdhU/Z6tWNCmZOFjmRk7s6eeLdh5NSG+Hha5nYSKpgrIKBHtbD+Z2zsoTDl51
6+f1OzktH/YuTHUXhY0ycbQ/KuKeWheP78lump3QOt1QDlQ7iTfS4asYkkw1C4Tr
H8imUcpCoPT57rksuoTpqR+ZqBTWXeZAeGqbaKojfzEPoo6U7icH4m9vimhu8Xon
3ZQQasfYzjh8yKKDj0T1lh+vKZ18Qfr4HR91rGh34l2H1km5UHExqX/P7T3ecIrb
796jykMxZupoXzUOwsrIkgcgq7FZ9HRIZurLgTbDzSafxi3sFZkYWTtp8qGsf4o7
DvZ6tiov9kASXzQ2DataOLvQbs9YaiOYaKtNV5sn5YrtkJOpm86+6RsVEeDkblVC
0lOkwn/VBh0LwQTamvrEBSNVesfMez2f6pC40CMBFedv8YM+NhFwtfto+6Y1nT8T
MIi7ciTAip1u0xEpTedGSXo/695k9baZ9xLI6OSRMdgZyCRzgDC768dI/9TziE4K
d+RML2CXXbuPKbwKmQhvBaD7vDtywF1t4TUOh9LYzMtFQfeV9GcCKMGzHkxS4ejq
RsZx7TJdO9vvtePguYR1GxYynJH56K5LRTh6DGBLbGXbGLPWfXs1dLlRTsOeDLPV
Q5bfYYy+tNFaNiwmDE8ev75ocrGDBovhBavaxj9t9q08NCpRWKrDGOxQeJECs9hC
ELMlu5Da4JQFNDtI3SzhyjSEPz6O1oHEJxWPKNYbhiy42qlMXUljjP7+zDgrQ97v
saDYPeF2IvOvFI7BqG6H3c2uAVYRVSEwdGyRM1fBcLPjFe4BcjBc1d/+T/EH0Gh4
mxynQ/ckVYrqgrZcPNN3ej4D5yFuQQuXOadj+KzZgG9vpyzKEi+eiLXPeM/7AcD1
/c/i+NnfCWLKDlPSWmiOObJXnIzinhVpJqIBFuy0LVpr5sg+n93r7t8neXULn+zd
dKRak+FM7yKj/8R07vrqLrog2joMUJZkfnc84MNULgingz1KOBw7I7PX3Fu00CzQ
1EiWuaBMcKCf7U9ZZ51hmZhfWTPK5YNLqSLkXjTtAgbYKlMKxIXWi/1Bm0keizum
aIcFFa4GrYlUBk08jVXX463yOXNvNyjdzgoTEZ25C7a36x2eawerm2Lr13dPaMkn
UEX5cNr93k752G3Pl46v7r2E7HBgBmiEaVIYjnc8DmimcH17MwarKUmEd8yDzMLf
xUb023peeQe8oXplp7ccSaHKNfmjpv0QxT910enR3PhXHY7C3uh0KUE56JwjAX+N
ee2XfUNkCQdNQ3x66poWvcuxX5IqC7mE1ZJS56JqQbaOdu65l9n9diPk1S+svWFA
KP0p/Wx4diUlAdYj0gNfLUAXmVy/sbHh6WQLVj0jxte7ypExksBeNWKKPQMAKDjK
OPxmntkbtMXLdQvjW9JRLpY+KoVIVwddjsXyrVwAmZGube+Xhg/7y05r6A9X6iF1
n+HHFW4tG9wMxCXd2TR/YUF6bwGi+kKiXPu0zMrUxeQM9A2hy1wrNhBYo5c8SRcv
5uOIcHqk12uPcnjVBeirdfeJJjtK0F8N+2WF/9wcO1l9AoXGoK05MYBGRosh96Jj
GVW+NGVvjOPMo/sJqvWNwf1VkpUsduWlxJxDpuy2eLreR5cQZeuFrqEVw5V9Rg78
fjq2R75detXjaHj538t1isfDqStz8yAYW16EoyKOy7k+66y6uJweuiYfzIb8igVR
aShTN2qRvVv34iB1cbRx18Zh7UNx7sgEp6NeECXdBfOlHZytms8A76okYihNP5qA
JFP0XDnoGFLthcG3E2JXTphw7vUj4vxoH44tSd65Flc5k+LnIKLzDgpSebQq9d14
GV3Pl1kAZjSYIC9ZWQT20eIJFzzTjW660thgs8G7mhCO8EinMyEFerptp4Dcup0J
tFjJMiBBXIQWxfWwwk1AYwRsvSFd+Thn2B/z0Rin+2xJU4nQuLBfsMR09P1YbXdA
Ide48HD+wKdjH37i3vD4H9uJKmm4SErCh5LpXYu099nh+330/iFiPwXw7ZCw0WaH
AUovFIz2uqteyvU01EUQuuobUko2iBs0QR7MapQ4/UnqNP7RUlhyjUuI5I8KDwf5
pZuVC1qr17aQYhLMitoZqF9GYLPEksJ8Zmk5z2LdwK7Y0kVfniv2LQCsFT121nXj
m78lbeMSrYded/IpnRRQcS4AQ3ADJnjIG+xzj2QTY5kX3JmS4pUAwxEPfFqueicd
tMOG62cnh198KMYsoePqol2OX28EF94ycwjxEiIRGeoCinRhPlz2rLJnJi5StYe0
7Peyl1VUxeUid7Bbh28K+4GHhltjCos7lM2tVeaNzWRbx/9X9vM6QxrWlKPJPp60
JyodNCujMrJxbGSdxuqig3PsZhK0jlni+jrKISw4jw43mcQyr/m8Q6+1ilRd8s6F
MHl5IhOkUdPotwPAxLZrJVWFUtQBYVpOu9bMyoXOeJgIYYc/paEImsSqeSeYAJyx
/HuuVJW+jJb6yU8KaX2gFVXSE+jplIgaYsWaxwrdXj7FtssnJjd0vTbG0iqV/Erp
VC++rdNFOQYCBdhptJX/HG4COHUZriHZW3Nb4b+15qPQ7LtcYK6UfdfyM9mk9b77
3bCKwFQ7jFYPHvJiLLkGIM2BTdJAWLVIXgaDZMep9yzZdJrvYJteQgnHk+3awZ9j
guSpMs1WcmJT6zBhXWWcxFVdwCtCqbC+fkqByzDAfte0yUPpvemsJanTKm5YKgL6
EoWsPI4rnsjbhU+4wrqd0kTgSUhbngkLvyga8e90h2EOtD+KvUoHfa5Va86bO8g9
QtsNOeN2gSWgmd2wGpVF3tnFeEhQ2qWN4X1Ib2z/bdregqr9tvk6pDnQp70QFuko
V6Cw/LS6Uj+VmRTpuUudJ+HIWge/Q9VX2cJg1mpqbQ5tUZB7IUSDEjkAnnwlgSEf
buJu+lor6Abo+D+A+8ClFUf4t2KB5azpaLyGNeXoptjZPz23OiqXLoHi4EUADizU
0cwMc3t3A7fGe4+w3B28Ic+ZtPb3UPTYM3pNgXAJuiUDpnFYUgm9lZgtZ593N7j1
ZGXc7Fio6gqzBgTScL2NsMpYiDa3ofw4L3GtdpSDt3XdD8jcrzcYlx4HWdK0mxjS
EKSAg93t2uIa1DY4Fs6zar0thEKk5Trz/SSfqLPwGMR76VU2J/CKI43bdxy/jP91
YGiY22c4CLnixrgZ1UbeGnn8ZXV3v0rJ1f+iSux2K3BvG3uG/xVnKSCb1+b+8o2c
W8IWj1bCpHB/KJWTEtbGFhGNCKxUXjkj+3tsvTz66ApoVkUKgmKhW/5OE6U5TW83
OBQwAK+Xf1KPlWb2u9qvvaqUPosez3kxiAWEs9hK63AQY6Gqp9Z2bJCKi1lqAhEm
Dp8ot3O1G3y8s8daPkozpn0+lW1Uhi9SqFB074XDjTyIqnhbTGQTZR5dk5JlqxGu
GynCS+KbW7bpNgQXi8qksglpU9ntAq9uUCs9/squ3u3VG8YUuPFYjvyaBEDXz6Fg
l1+9pS2r+UD2AUvPkUCpdu6lxfGsokv8jGpSi/5zeDR3R4GnDdtf7gYiwBmpnPJd
Feg9//8i+DdQimB2kpqxeXrDN9TdpzL6WE+ztMWRaTIyVuAXiW4Aef5l16j8715P
5Sli7GKaxm+wRNfGQyBZuKuzxVCqkkaErY9AALK3rm5vBvyNPPutZVgfvH2nbgCD
Obcgk7JrcD5CeidgHdEGZnYOXthOYj0Jb/8e9vpkLcANKGeIntTau4Btz9JdqwPP
YSe5hHn5JdLZ0bMtSPtorsdPEYcP8HetOBrcPPkPfUrr1m1uJcsQjZWax4GHZjHY
0VuHEU6CVTZlYFclJmZn5KiuBW7eJPORdY/omn/IhTOlB/5q5en7ub9m4wPQjWj6
pZHpZklWZFXXgjfJif4dYqx68oVzGCzf0mBWDSy6aJKmXLho0PitPUvuVZZISJFA
ALkWOkhRlKg4XzpsUKHR2neeFsTS9VKLi6v3USfEgUZT3/CLn5+l9gtixPCS12ZR
TTw5L/MiVKUXtwE12FsJ7LIicbDOiHy8l/1eShF/eNLsBliNlyOtbws05PXVTV4+
Fjp9A03Q8soJ+W7zccUnShJslEu1frb/zLM1u7scLlIUUHl5FSPCjH/5gOIGmwbY
2f+xWO3+PG+5HWqWf02UGmcDrHRSvPtByTBQ+HktGh3uDMaSBWDjnyTcmG3YVO5Y
7Mq5X2yiNeyB1On8ge/VjyVKKJSGf933/xhZgu68hk2o9oNnDvfWEhmlpXGr8X4i
STnXguQ7d63FIQ176jPB5tqvo+c6xSxEOjehP6qJxLeNCdSRM5UNlO/KPTVwllhj
uR4ooJSQFdtW2cweskGxg1oRBLGhi9CVYj/6OUgy48+cGG8h7PK8IOF4ZbWKAdeu
awqxVC2hsJxqAIZu55nMgK9m6rrysPWxcuwa9Lv2yf/xYaivSgjRmcdfsNK2Yqs+
4gf0OBnkbv4UDNbY1XINzxufrz87PwSV1hkL0xpS2SQ7Lt/CMGAKxu7/r6linGGa
QKQDpxa30LKIVbMSPBiPmJFgrOrFkQclb9K8IR/lyH2WviU/V4TqLJ0rVFNAQ3xM
Xx3maRcFyU9ldb3kd7xHbRDQjI9ISYLf/gTnXMWrnCCM/ofeWB9UnygztbA6vZ1W
Ik+OPogstrpbIc2LuEzicgr7k8Awz1EuqMsqVhy+AZOrzWaoY1cXITvBHFgcRjQa
pavgwfM/wh574lCzu4Bg51UjL0wLv8sDqWMtelMV4bWYLgpzSSOre9dPZEo13GuR
0cl+rarPvFr3rMmwRsLBcReO+9BGoMqNJASIsV9bWGuegf8GrUAkc4MlbKRsgjub
Vo3Gyo/1NtG0PFDBsTOTLYgyMQtYTyATC3reCAn23VemQ8H/5nV0/9M2DlMbxDWk
ltMHkCik5hUU5ln/TKzbmF5n6NCOhqshT/IztR4yAUxZL/7BJXFr7o03yeZOANag
jOaYfXWkYSGGvLIz3ZwF2i4FNbhz7LpCf8nZgxK+CJmi/xchZTkZnPnt211gJxd8
YjN22QthlSZKA9qDAzke56Na3EjED0L8PDzx9keSMbVEaUdLIGJCBr/V3eJ6l5PY
oamnOybkbwFW92+KBh1uAZ9+J/l/gubxgHoMkcV1ja4hc9fZWOH9mKEqT4QorokZ
37zc5Rxz0Nb6PudHakg41tA1V1dw9XMEhdBjS1Qr/pwwpX45UJt3bCmcY2/PJ8it
fIoAssytdw31tZnvBdmvmFX8k1pGqC0cX0a1VPKdn5nxlzQRmOA7JMo2JnAJsOaX
buTEU06O+OrZx8dsbHv+97D2aCpRMsqfG17NEml8Vo7RcBCjiWLSmC0+0P8wXh8k
P5vZw0AZPb0QtTf83Z6abOn/yx7hSP7qMk0Eb1u0bp6w7IOF2XwMU9E9nofCFHb5
1KFG+I0/OZ1qWKSx+YFkPlXQe/8jowWOZ3v4I9jLoEaXNhbJb/kdnTStAYcR7WTg
yF89x/rNsw/bNDPWJuOSCqhB/mAWbkBDKpA7ycorvmtisdLFPIwIUt7VVkPa/dnV
MIR0eRwuPg40k0DuQVCIFI3CZAKM6/CHsIoXHAtJmH6zr4zL0pTmYr9Xi2Zp9ySk
AiLRUQSRqarvgNcaAOH83nRACMqTvub+hnjccgxhPa7e7t5BwVEs8dvvunnJJUcs
K9SXkmL9DwV0zgsEHf2jEyZrs70MZc0MszDZJ8F15ShQL3TkB9TtEIoeCGlyEA7R
hC0irD+DfzBCkU4Pd0yOfo3tokdIX2HdO4Ihwbgpipw/kZ5n+McCRsIGNk3vm7pw
XtYgbK4/xFny5f4YGRDx7w3vBebBDhMunuLrCd41qTngo9GkdeXnSbpPJ2GPGTI8
uNa1klcJdYagZUByNz5Y8DDQuWnSxJUPRkolQBBVjk15KwhYic7p5Cj3teA6pF7E
6DjnN7patgMjHm5ycrLtu6f4BCQAEQ9dzB0jld16oe8qZ1OCNRuaPRMvrCZDMW5V
2OqK24ljsniDbkO5QdMAof00BzBp0z8gtpgxjeIZepmHqy9U2K3AQY7gcyGEApe/
Rqobmib9WQY867yDvEmV9jUxc4IeHPoB9YcUy4ACvRg7hDMbPiiIUA7weXRswhrb
TQFkVZZRJ/vEHfNQICkm5y3x9ra3ZPHzGQ8yDLh6sfeoopxSm6Wo4zwXPxblomE+
MiNu6pMIvwXEW+QXeznwKZhiki5Rh3SZNEHOjRovrhoOzIcYM6oVwMF1/YxFiRQI
YSEvn8LnZ7RbcjpH/h5PQBq/v9zWpl1Fr72DgfpV2tjHpwQFQ/LwVF6l4FDBFajb
zihfRRQJtW0GmVAGcv0EG2wVXwgKRD6O3c+JiBlqJWZPeIHmyLTGK6QM6GC9Han5
IJN4PavPZceQUAuLDdxuXJsaF7n2lWIQ5GwZgiHXjHalUywkQZkihfYgr8a2RaBf
O+tXu4ljlM6yMHRojp83h9hbTuZ5Y/fJ2Mu6iT2putXj5SI8PIfFoTaN/YlWpbPZ
LJ4QcFP3OPDVWLOeoJS+qBjkmiZZlUjAMd1hJS3jiNfcluQjIqK6UHqxIC1ZzCjO
eU1yBqANknhyr5Bt06uNs+lXlWQ3detmxhvbk8jo2Ne5FjrX0K26sc2F+1+etEJy
9FQzhBhTCVm9jqB+c4mv7DTpieq/Weg3XtVtZF7hGiG+KTGUeS0KQseQsnYbwcw/
JmHi/5WmGfMNAa0OhqY+shKrKYd+xfAKnm18MY1hcXdreUguGt1jO4P/+xRXQs2b
xw3TOdNPOHsL6pPlAWjAt8zHrmtLqH+KFxFrRkWKPFytoFDGCDXKgUe33hM38hTW
gKzrb0Toez+sYZxfPGAQyUQ3xOxetLREwnWg1tYj/DzPo+w4L43wWcAdiZW8Pkex
rV6VVL+y6plaLH0SLAM3wex9r3zp+Vqkj5gQv4lb14SfYnR2fqaP/wS85KaIG1CJ
z5xErhG5WKKxwwG3igCUTRNp8ep3hm6TTWMTaexc/vj8NtGGQSyC+nolT3+4Wt8q
B24kZ1JKkkyO6LXdPQIsqeakLBQfLggRyxmGy5pbm+Tlc8/x3GZ6ORLMty0vBHT9
HaJR9BWz6vGcU2UvDGsJrnQogMkxRnftBQe3r6nzOLcOhTQoADbUyv94NyB6C/ib
J4oqN48lXLp/NnWDU5KptPmyuchNXdV5zIoNsU3CmILVkZhGn7iwjvZ1XA3hkwaR
1QXD0RoeedJxUXbjaFF3lKW7WJj98vZDdIjO9C9vB0asCe44ej4lAxYjs3LqQnkn
Ydg2hTGGnJdAhsfKeKkJXknulWjGRGt+WFNldlJTd8jqO6kthzm7KajLCPcp2sQR
Vbau88knWrdopzj+bzpSBZr7uj1yCZ58GbO/feu1JJ3RmKCUgyT1Y0ecwDhpOzrg
c3nITEZ/oGVTthGDtwkPo5YGhIRc8rXQh10sknWZi+9NqVQsuHBCrMxBqZmmBaqJ
R6QNiiC3QN3CCIkWn/solqw3W0J5wkTSQMqYMzaM55bvb5Tp7dYO9U2MmjtkEtIE
IP9VB1d1jG+Yatg3Tr3gzqzsTNqdBB0IzHMczIYoEDUS0/+c5/6cwtC8OSHkCBh+
eIqiy3sYFKDZhBhnwsStXRbUX5+wodF7mhnP2/KiRpM4RlIB8GJZcVW9j8JldYuU
VltfRqk88uo1IAwcYmiSqWE/B5rVozgCD6K05uR6E/DGXETg+F2IeH1gn8xmDp4N
omW6JQJwLCYkxTfy5m7go1CD5vyQqGMwMW28KUr9bvOvFSwcesWpDdiKjrLjpQkJ
vg+yvYaOddVQNit4WoeTSxZ0qZQWOugAp14+Ou5s+WK3NfnkrCDnHE0/5L6wBS6J
B6a5Gk8xjJKY0NgKw/z8Mt4x3GdRLvJq/eaSm2o79rGhg5yvQG67/xFHHCC/LYga
1QDp3ZXnNGtbsWjtShZZYHe8SSlhr8HykFQ7Kz2aXKW5aN2CeC3HgH9XocNMfnl4
KvrEDfF1S1L0qJIjizAguPqKrEGPx/3FnoL9IKHHUh3lz2lDAmXwzSMS3n2jLvtZ
70L6EM9+vgtlEUK2BijbCxaTaC+9Vlz15/Z7PYx+fiGQePzpFUH2IT5AFYUsYMTY
LX9oAxo8kQFFyJx3i+QTLihRCsBNEgt2s029YM72GLCWPgZ+CGTEPeeeaM7mwdhS
k/nZlW6HTq3YB0GIWbS6x0SSGQjmtXL/IdwMKLnq2KeqnHy+Wt/opXBxrPpIk+mG
B1+xUhAYZlGVBmtSnu+tvqqEZNAv1A11rgnAqT71NGtgYwhbNLit7XyrnpqrDUXh
RebIXpngGZQEA1WM2xIjvvTaM/j42ATLxDBMMmw7ziaMBU+JvqoGRSbay/RkYBuM
OStixAFLCM6QpMwknxu4BZEM/zOgt6aGgjOhIrP6roF9pPLB931nAPE2LnKZYsYl
EUQZuc6w3Ki25bg5ym/hqSMtCnP7COCXMhIKOXABZ+vrjTq++uoxtlyAxk/Gs0Re
/vM3+VB56Pi6Yu/vCYKU7Gdk1bFebI6oMsa8kJXVZduC4uSzQbsAtzoLxTvRPowM
N4mU7gCXC6ZDvMM3YfeNuFZpdpC6sXL0RDaQH/aQR+TN1mmokLOWY1j7+NWz+m+O
PtAGa+Sxquymg2yAJmFc2MGA7JMIEDUfgoZVEaIsReyxvn7P1YrCiBGjt2sCRvhE
zRJGiB3FQERKv+DkHPLCKzkGuXj5aCyS8drPluj1zkSLbmC7UutyE7W5YLsjmMlj
H0coCp/COzU/qGK/hNZd2ckmg1sp13vqmi1/ODWz8OHTg+MImJrCje/IgLcRuevl
nK6apdvJZRFBzCya4FoPSEzQITgGhmv32P0YJtxrZkwcqGq129LoiG33MKCmBWQR
lS0FieVfc05GR9CPaTo08NTbsYk9mSRhMSJeBkXSbnaST82GPEUt17sO/4UO1g1s
y57Lg5rbw3JAn3ApWwDOa8eoRYllW00N7zP2yilPHeg3gTNjTWmng+4ZfMXASyoL
edscbAAfYEacvppkhHONwbI1NBhCsyzQN9saEGsHCcWuZs2lM7QqYOegOdPl+mkq
tAF8E6FCZHWhvSSd7atw41h/9gBMK9EmJFJdjoYetbnROlnCgJ+vCOEPmEDrKHbF
opBYiGZFTdHvp35CycJTWW3+IDWdV7dVvzIXU9/AkKhHtPqmx4HFDR7UclzaZr2F
TsnE7DUnFfImg3iGYE7UoUryUkQlOjvxw4cozYY5+uaYIXr91HRiqOxhOwLOFL9N
5U4cMLAbYpnhXVdo81c6wElrwDneb3igeubgkwiNBL7StK6z2syTuLCG6Vj4t5cS
qmy4NKle5qNaSM8MOd66yK4PJm7pzt1Nv2a0nD0igdsiHfxW6rgPn4fDK3Rsimxx
94DiIMukLwDPTkpZa7RAg3UZxc00ALqQnHKXkJakypDQ+gftlSssgY/4ABt1PoeX
3MrghgppgiosW1EJvf/gC3vpw+2MUCBgh6MBM9XNpuYoFyy+fksv1OJkp4Rp4Zsa
EJARfzIGY/L15T1+FQO1WgjzdRHL+a/E0uwxLNuugqg+THfgPJ0TmrtACpAZTYoe
hUtpOEACZdx3+3QIH0+1WUj7boy71Y9wmPrC4S+yNthYem/KdEelS/uhM02bW/8c
QT5YjKqtNt70LSX3nKP8iVoMAP7z6UDkimaFakxQx/nouxYTN/8jAXcP4F58IMzc
+37XVPI9GEsOiXcYPIieIeDMydmL74OpDUgQlnmlrMKjIe/8+4cPQGGAWcu+uewV
UEyoAKT1PeS6Uvuv45x8jqVrKRHhVpf1syobbHAof0UkBll3Ck8s+zcUFsVL5xIn
O5nGfH/+mGCBdyArqwsrRaUO+UrHl3vivZjRTr+n5LFEPO+J0OK9LpMtGLf8MJss
j+sP5xVTKnrXKzQYbZWMrnLfbc9rzegb1bGMKGgCVwiu8UmFU5/uVgOm8zY1A0IY
ENFHTYRVH3Vc0v72TLGjPORzJLuqNjOupD7jNn/3gm2eV02nEPX7mQ4cnuWjwUD1
558PbVsdqWSSl9NqjXZZTPyS493mL3/yhPbdrUEgM5jzuTproiD6baos/w6GmOlk
cn1T+igv9bF0isKFPL2RkQrb6dLawnX7z45DO39m+XG4LXR0Xg7bn3l4HNnwxnys
vZDLm4tSwRO9ziTpnzMn+YBZImOuOGiNq71bZpKrxSRbjrMaPbGrU3bnA64LvpuH
urK1IYKpE9VPANZej+Gi61ymwwv4wa6EslXvHOS4H5fRBd5DoT+GNlm9ha/c3QP8
DIXskUizod2y0jhzp9toRMsRUaN8E00IYdx/HujEuUmYJ9K9KWykZuMle4ph1DVw
f5YqCLAXn9Yjlw1BFhZAREiYu18Qd90gDE1VW7b6jZishTVylrq6Oe1qYe/ZtGsJ
/m/4Ikb2o+2KMV9SJBhIunk0TpBGPP4b7Ydg52xdpmN6iIK3mzL0MQZD0liTVAj5
uEmQmqPAtrJF+o4ViImh5VWH9frr7IkZJYDb8bVZsa+IfXe+3wDZxvDiBnAaX5Mu
yimZgeGMwJb5SSkHqGFt4K5S0jygpd+4SUl+rquTrV/QQApwly6sAKnwEn8whap4
1kcz8/7h8Kb+WorPpXWcgSRqGJWBetjSuZaVSnTeDei3brN5IRjKdt0qhdaCGc3S
DMwv8C4dklooqaNiXfLjU5hOvT6NonQ6RHj0HYwWGUA6Ti0RHr5p43fAbyPsSBr8
y3PvhEcJ9gHyGWvzsppVG1+4yWWl3q3BbGbnmlw2wHoi6gg4udhDeCEepveQ/UBj
sxwuoeQPRRtB21RrxW5i4lO1MnFCn0g3psYhBYnCl7/g617FMjm2QpP/iIILctUL
mlRLfXRG4aJdhYTBRoJoZWYdVEJZRETFcstdm0WYx29lfEqGG8KpPS0E/tZti5br
FMFZbhzYI5IS8GeO9rkqDQU8urfuM6pD1Dn66vP2dqWnCshxY3LDd9N2a1b4v9DE
yeBt2Tz6TjQIzIoDZ2ZC0kdnrM2fKjdmYH+vlp5SupmVKzjv769IzmcTjsOM+/UZ
rFqdDRiCzVLIg6jkjm3g9yh4sbUxQ0Md+k9jSYzq3vgjm8RsC++whkKpCbuUggVK
4P4yw64LduJpNXsP80ac99cVErQvE4zDfnN1siFHLip01f5DXZw8ztnCjWabFDwn
5QtLaVWH0YjsnvMyHmXKNSZcpmVw44NMhQRj0zUyBZaaEsI22aKJOQDzMc+Mfr2Y
OS+irJ18kkxi97+cYPXEA77KGfwrDMRuckGiCJ6v1qbzR9B0A6VV9mj80jviqWFd
VcAgiW5n8ugXRq/eu3Jgz9YUevq6W7gqZmGtwcbHI0mMLLumoAnXmNUHSPm+PcmL
fwTKSHWsKZtaDneztMPe33WwKuZ0cng8eULVXrS07xReO+dEHsqo341Z/BQbvV1F
TE1Zb5gX/9dAEYeuZvbqaZdI7Gj2/rvR7sGNmmcYkudZR9jjORw+TMuWgtM4D/yn
z+I1xGRgw119NQxjUDOjulaAhrsoMjyI+dsXza/sIzlHYCwXxMcaj2wvPFg9Q9Vy
YaFGwBCZDFqNipmt8PPAd/fpTT2lW+W5xcBW6I8RzzJesmRttX2lXmVS0WmU0zzl
B55MgrGwELA3P5LsFGKbYZZMUEymRgwARjjNkvBPo/9hlt+WG1Nv+IVripYdrzXj
Fe3ZmY2OMa/GBueoQSYPUivmsi84nRztIh+00UwLvA9xE+0MqWVd/cho7sfuEMYB
99CSShOx46M+5JK7ozPA0GC6B3idwNlBwfVT0xEvzlLWTGWB/3Pa4WjZjiJWUw2L
l4nDtFfoRlny9MrhBS6N1XHBnE4oQ1PYWzSHTw7PCXkzw6vqO7NM9u/oRfLPA8JC
v3OXdxYGTgRpQwgw2LK59sUM7Gqg41nQdR9N5d8bKothu3lxNxJHkE0050tZbY0q
uSoAbDDw2Bk3qQMxnYmawYFK5kGPOrTbgChN9i/fkX9Dt/pFYsd2bsJCXhjeTgsr
1KpToBd4siWv4/0PZhGJC1MCLTzcUIzdQ91PN5JvPam+nZ/kuV/UHmX8u1xhin5v
W1a/XzXaqqp6ErysFGMrPl4BmGTh1BQwEFG/wV1FVhkhY9am/dstvQsw5n4w6raN
pTzvaHYBeeoSBXXYCat2X4KZDOXt1a3RJFMZK+/iysNM6j0vTbN8qJE6uFf58gbD
qy/QxSXktZO4ALHx6E38MDutPKAhX+ikxBuXSVkxURJ4Y2seu2rhwKXljITGj0e6
WHe458zH13SAHXkvymuacLz0j4IObzYhCAYMZDmqmarANZkDqg+ATwpA6zwQe3xf
ZJlfXLGtwMKd15GhwRPqAPS+CW4lozilGD3STPgg1aElhpJxsoK51gOUeCJ9A7in
hSJCoynNQ10Tn4eyRP+3Z8GQzmGacf5KYRngCTRZHw10FKQ+CVu+KpsCi4DXnf9g
3NJcASMdirIWDtew+KM/DTmRXDvxBmTho7aupK6U16zzUpvgjHkV2t3dVCh7wDOP
jg6P46j9ghqvRIju2jaVb/MNPMJr+WGql80sYVEuH5FR6daLKeRukRb7ubQmfKbD
fjedwXbKp64M5XZKjbfXLRVHyRbvKzaTkHjVNOrlFH7GrCqQFuuUAfMyhTe6O2o5
FCtA3prKoNUxaJ4QX8h66Deqy309trd7vDfzZy0OYOY3zwB9hpd4iPnMWO9sbLvQ
sqB+d6UsARl0VkWjd749jgIBljVP3CeimjeZvVm2yqH2HcH+NFNwjGpgnHk/q7no
dW1IXJnRjhE0LmROMtPFpFMO3CfXkLhXly/wInvxH7JgBPviujIM6SZ44TFu3po4
4MHcLltf9K2Hcz9aSqoXYY1tRvAkuk4PwotKHgeoMY6yKj/smjxBwXiDAyYAqIrp
wXPnQ7OoXNrobt23zDGc5FnN6Fht+hGVt8jqdXIjEV9l1QB8HrPb35NqL4Mm1ZVx
nivkiMcq5291Ln2c9von4lHVR2iHojy9l+FrzbNNk+zEToFbBOGWpLS6vBa1rYL1
3PlYz7WF/EuU45ZrC9XglVzeJbD5HohbccILD/DivCR2/3uF1Y94QxRBvFpVwrkA
CljCAHy7mh5VaY0AbCDcdYseO7hrri0QEgctN/f2TBCxKx9uf+DWI6/cLevbVNNF
Wmvg8vT8V4i/zMtqUsxyPHWVAj+JeKvXeqUEcVThc7P5a9ZdWWlAzvARxx5vdWGk
tL2aQwFMexf9nV4fO+5rvSzgokO9Y4NbbjL1+iHlmTrVIelAe1Lc3wgPKA7kHCES
bObeLRUtHoaSeSmxwlE5ebVx3aECQ2mwWVteLB1P7NSk4tZcGWjKQtS2qii3934t
8icWBYY/2Ai9RN270NvnQE82mYtZDyQ82rDb6zITo4VrDoASPeuZ+D1iHsQDLUoH
IM/EnOiOIqdyD5t707WhVGjJkkcChzGpPipnKE+yPe3+j/scuG36wx3FFsy4I+R7
qNs4A3f16MNYkw+FeuqiySm9DD9kzaN8TGmsT5gZidjM30wxEbEmjyGFVJ1xLR+G
xRzGN8W6NzsJmvayIl0TcrD8X2Xg8WmnQfdgm1ACFh57yNwZGB52+MKdry5s3oyH
C25c+irucesgNGwSjbOoD5RgD62l0Q2nmRKiGqpgGQK26LLbB1BdBZbVaZKoW3T3
ggf8Gr58IUKpZsknqW1EzE94Nx17x3xa/e8GN6gDDEAB+Dx9rf7wu5WKWECYQDR+
LGSUJQhGwvdW2eDy+p2Lu20CCsThaOzFKhhe0O8ZJAAB9WIKx+aPJZfQ9EeLuMud
pxbfnmSTH0+QvRfCnI3ukmWGm67Ivo5uBA/b3ASfFON2tru4OYjFkAxjQXZzLvJT
bNKUndMXld+CWDc6hMtqm1Ldjh1K3AwnRmit/PqAQp+CjrOgv6ZXAKz/X8MjpW/l
DGhBAhxk9jh54zAe7Fga+N7xyKfAhn5b/1D8ApbCmPzCiPRmKkEbdEaMEMvcTvaQ
p1zKvhIT+AlZUKqG81ydASHh95AUTrIZcV60J7dYx+UHK+zjZEHj823wd+ZuM0WM
DfrpdNGMC75sxs4fRJSyQXanzNhytkddQkPkWKZbHDuGIgTnZ0uYYJkH9Wh84WuB
tMF8hin8ebPJjd/I4VQT+ud5OIdZjfKTYeQ+3do1RmcyR67Z8Aj7s8DcrfTIwCaB
jOrLoJFRD8KmtNwxlMls/CoYhu8t/BVjRw4ailneV/Tm+SQUbRmNkWJEZFelfcM3
p+Sz1HgPMzaO5Xx7sUdJx8mI5izgYfeU5zLZLwv3CSuqIEVvyI8IFZNEqhe8HNNf
pFGam0mfbQirLsxMpw6E8Mg7tOML203FJsMsmgus81ZwFBOxzo87FMpZncW0Lskn
hT1O+SvE+CIX1j/JcGKi8wNUS1ZoAlDSAQsUuHPJYVAZZEmdonCSWYzwDCPNLNOW
71eLUgO52qjW0kTEyY61TvPTLfII4ZJ78rKaV5lkEDRCkiJoWdnOSaIjp+LvrnoE
yqLFfBb9zxKaHA1pBls8nJYXxist8vu5W7kxIWNt/2ZvAQr8Q35UzK24+WEIwgq6
ytYifepa9xThZLq1Isy75UKLQmyfxzO0fee7gzyGHxxwkcpULiMuFMg0Kka3j7Kx
/zfxiOUaf+E+Vn3c7k+ZAKhlaPHjYfeQXFZg4mxYITqOThWTj1bhs+a75jWGjZ6C
o+43DmsxudVr95p5IyyXOlHy+babkcvoJ2K7YRKjhLz/xtArccCC9S8JuoRH1my9
GhUaPdKA7INFCYQsvvm+j14udDoS8WWPEnDtUAWKUv0xbRh7r3P3xpDfzYulVgOR
vtqmb7t1pu3GHW3QbcR4NUDl0uHOlFAPslV9pwIPVz1sYpkk+I3EsH3ppS/swFQY
G48YUIVZqiNyi5Zkzmi64LKpT1rPrYCDJbmD4GzBZc4P5SXRzsl7ZcrWf0hG49yd
sYagYx8Z5+YXHdiYNBY+kqMhyQsJaOuZIRBOsVCx/MMMO7m8jyKcdqA92yOjirh3
L5wFSBoLDk8qMxezHshHjuWIz+cHN3yATSNjHyVt8yFNDxc1aRrqQX8Euq2IrRyJ
UPHUbL6GEDvfrgtkPAvPkNarWTmhkRqZASfV6JfeOipwaBjAFHMhkYYHc7EAQup/
kq9Bw6GU+6NRwtZldh61d/maA+7iscHcdvM+HrOK6vTCuTvPtuqzc3sW0cXgbPtf
vwuiKF9DvwW3Eff+mN5VDoBiitUbYaapQuPKkXVEcrm9TvF+zD9Je7B7QpjKLbMj
k6h88HEg20k0GlQ3FJPR1gTvgX1/UohewFJw2ruaovHUIi8OxIjaZums+U/hjZKD
gKYcLLVhJ2Oj0q0I7UkMNzNnjhDAYi+J+tvaErzACSh2R9dzCl6WQrGmUtz+4b5m
wqip8CYBrOIDmu0ado7OpkEKobpbF+i3wyv7tO0IOHBt9cBH6TOHg2delh2nPIal
gikBSy8xxFZxZpFa4EpPyIrWWZ7US5BqvBocvCTBb+5dQTnYxjXTi06ESkccgoqx
JL5T/vmbaZhPwjxAU8z/Sid84/Yzxm8SwccbNfwR4epeR+zcNpR+ozOK4RAgn7rv
zuQzowlHPN8sZyDOQdm3BFJD4jWvdENCKjEP+lS9koEd0vZIg3HekuH9BpGbro5D
LsudGQNArMT58yMMoZvYUtinxRctjxz3oVm6mgOWXRkJ9kSi/Ye+peSip3pjmgOM
E69/fU8TpVJErt9O3ot3bRj+XqTTlPX2CniwVxwOuMQu91b7FZM7rqiI99UhMs3d
eckTXHcvm2IFOJDj0yeVjRzaDJijL/TIOyPObvizRaE5iApmAW650x7DtLyWPG+r
LKYHZg6dQl8ZyUz3zCL6ChnhqMYl84vdjoncBNrhf3bWGaAIUtmLcWMwVVgtLvg+
PomYNUQj/g6SOgBL1h5O3w/EdedaxZGvNeGatn8OIrh07J6jALaif17aWWqNcPca
LyN2ijOhw16M/WfLrCIKSAzRR82tBs6TD0FCZcMjmSzoZYzERKwjsLyrHl1H/Vux
My6kppsiyNZsrmPY2keWGF0E2ilfHRuyUw6SENl9s2SDPkiKzKV03RwX4re2Obub
AHXRgNCkVOPfh0Wg9S1y/fLEqLRk403h3aSYIsaaR6cDQ25/gv724m8LyEEq/eRH
aOxzjgx0g5EubWbEUu+cHgeiTrJmhA+WXkWh4ZKqCPgvi2E7YlWHeRowUXhvfzEC
FpoQZfpEMectbScxg5gHcKvxtGct86IaphlAq4ZnHproTVTWzXzDkUbHqppnPP9D
IJh8XBvZ8TbbQ6aa2S3Rmmj3LZGNV4Sg7HsJPmTpRiKc1XxM2Xx26Ci9hyFNgXug
3CsuGksM1G/GMQ8gJyOqXxnOUR9a8H8WhGa2LEFrSvZGf8zzNRkAKn6x+ZDMci4S
s4cVfuTRBTPxys4p+yur442D5kb+fVVrHeMXvzDg6BF7cg9trNmlR/asP/V2mNjD
lnpUBmdgpxlyPvMJdeslsXNnUR8ZKOa2T/wWVfnHWH+MvbD/MR/pzRTFnk+4Mif8
2DRAtbA+Dyf4NbeUXhJQTqmpY44LbuewSJkBiKrQBtIZ5UOb0xU3fN31/SQzMk5V
YOcRGfRPPm6D2SPUl7p6R5SnCyOYZq9xgZ8lIUWslAgJVuUvTeBQJHEx0hVQHYTT
eZBLc+8CmDo7/4mHaU38kdkuP288vXxZMVwe4CdCMe4bLwHLnf4dZIsvhZGFrE6o
CFSng9pHI/MNb2xKcKNEq1wfVehPOuYuZ+gfVRO0FGIjgshCX97pkf+d3UwKAtTQ
Uf3RB6zXimB7zWsJwJcZLEf/CJz72n/QaaT32NDpUbFoz/vj9pn98uCEhFBSL4XE
twc8fjL/uBGn8dRk0kwMpop3TRNA5ES5fdFaXDya22ujio8sKuy6vB/PgdaYmheC
JDkrNd5PLiwKMl1lB+pqaPG8N+3iRpEzyVA8eVECsgKSWRcGVibuqg3Z1f27Jrf7
tzWnb0ySIobTssr7jvgSr1kyWawUoYzUdbBoobwgseaFN8MHicdQksID2pG8EnQ4
qC9EMgVZh+GVy1KcrIWnXSrt5NRLsAFxKSi211Zi5J1Wv0HttQG2P3xB8/eilXy0
iHEQ/q7U+x5rzNm817KxTGUhz98N3WRwltmbpn9kZGbq3DYTnH4EtBbVvqvzxdAS
SQ5IrM1PNiYIFJYXCy44ZtZRPpNj1LMaFPJZmkcFAbMfzRmX1Nyr332HZoDBl5C/
/2kBdBDVrD7bLgqGej2AD4L3YBF2FHFfsSBMAZRq10CTQjs5+dgPR5i+PDNwGY2N
/NwBgCZHICyfd6CIbY2OxRUh7GrvN5qChahbIAhPF+z/j+zALpw0+6+YxGXZfCKr
yvGYW+6pfd75TMx8ezikF7F+uxGqn6PC2GlLTa/kYnr3rXEctht1AOhy/0IjgRtG
Lgyuv8MayOA4FZbL2tp7uDzmXPF1xqZZvSMFmnRBiBZNVouv3rWm8h+a/1aTiEOe
8ESCK/1QcEMK4uab3rxddyBvqJqpgdTHs3Jlp3jG952I4Hf+Yo3rOzz2l62KmbJB
jO8CdMLSWJWkWmoq506DApuh9dBVHDCkgHPwYEHV+Ug5wYoK0fUBT0eACKsOHAXr
0t/ublVNr8pbTxEYkv8Q/v/x3npJyN0W6DZqJ/ZHRi2NRhfZdNZaQnpXAm8loLte
gIZPT6rr1Jx6qri3X474F9rz1//obXT/sCAq3S2Cf8vbr+CmVvWTE8I3Bl59Lpdz
Tfda3gLN3qc2o5oKqd+XVj5899DISUQIXYgXzvbleLXeUySiHplvFTX5opKTKrcs
1REryC4GizBAx8m0/tNogVCONFPN4brxNSBQ2PE3RsSojaBJoMdmlp4KjDTCzclr
kPPWicVuso055pa4HTtxTPpBZyXVlra9AWeEBcljWMn7mdgOxai2rFsQ7Tecj4hX
Gm285Hpe2J8D10sqKVrStU6PytwhTgp8Caq4rjrDSMv464aQ5+m+YRIPFVckU8mG
wH9i3lhP+OfSx6UVuEMSBC32N+9kKnvG+cDdP6PfGP6RlHDM1wg7TJr3qPSssTE5
/kQqmRHanZbc1IAf6MccgUn7kry8M7flk5YfGW/RubKy0PPwInVaNBe6spNtXBPX
DF6ZuOjrSk0hBzZv9D/w4NgBjpCnT946VKYzEuMJ70My7y9+8Fe28sc8vO4rJjF3
m4UiGi729+FgddGQLHcGaJ2dEFNsv9l8navNkVoK7pcAUX4TxBtdqnaLdBX7avkO
7s9CSIA3xgYCJF2GsHkp9CZ2dYzhyW7hpwRNV9oS+XL7dSuc+Tyvz5BMDG2xCcpR
jaFWdzb7HixQEb2jIJNOT+y+t/sCrf/jU127z+G1Me/TfzJnyZa7jXqzVQuZ6gB2
GGg5LiJVXqaRxhMaKNJ2gSNvL4aDqPfHZcElk+iSXT3Arv38kKQB/NPiViey6FQO
Rs82ILL54Lfc2wTaapFdGphTXHaVW6qp7JSRu+aVJ9FNF3OhqNh2IMR4gxnZw7XB
bK/fFwQHv+hS7WVb176jtmxmJ6gEQatv7HnMBDwmLrnba6mbh37iQYpZmWhyvirp
KsEA7MzQ91lXhlPW897M07V/ky3Ml7DgJm/bQGRi4thSin25LcsdkVF6yTBuo73/
hOFnQ5zXU/W8a5hsTgv/2xLnrDExzXwHcbIJsuTMF17oFeOfDO6o7aPQLiwoJCKR
OJDbnoqFI1HYfjNFigCEyL+GLPyd3TmPw8lL3o3J9fsLIZevcB2/DgIvLsKyHbwK
ryzbUe0w5Gg94NfGjQwZ8PHqiXTnf5c2n7mzL8mPdLrsI7rpybA8gZgD8y+N+mue
Lrqnr0RqckRtckl+7f6G3HsKjqv+XgKTPLsDzGAK+PRGIwEsk9WxaipMYoe0Py6E
5pqNgCxuw20DjgXyy4WoKdsejJ3S2KxpLVksCiVqJmLCBN277hHXN7YbGJ/rlTtX
PhcsSuoQ3myLUt7+wiFlD9HntFQ+5JHZ95KCjteE2QI1H1LXdODg4v5Ho/h1MGNY
45P3mcy+Khs0aOtAryTxG1lQJDHUdhpu/0CoH6Ggkj8obowWIR81MSr/duighSHb
+K050XYCUuqp9asSb2cXe7BZMukngTH50oTXYjk0Nk9CTvjq3dkaLensSWU9Ugd5
+lAuWIVHIHsXBp4Xvc5Jeq7lNraBb9v4V97H2fS1Z4qP7UuDezjrNxBoX0y9Jo6J
jGeu69ra3+X4XpDFbAr5A1cp+RPe4kpc33ZQdbjYRVOIV4BCIxMpipeKJBCfXCvS
ZZY9/ewKnGSU4kr65nxIAdwLDtWXBhaAppuABYkQjhzG1+MC+HgMHk3Fp8SUqWFn
2D+aFpR1cDN/OXrySmRNDi4fvHQ74Ja2T8QJ4YkIf82jPymHPb6nV/dG/Q9fljZq
glINSe23ZdMvQ/Ytj2FwT50WAfwCA707TgphZVQsIW4CwnsnrNaMqSAXzG+gUaYr
tl0G+wKoValxYWVuGmGck0+ffa3K42lbTnZPBnLBI/kWVs2ggE95+obbhkT9BUkY
V+s9Q+CLM6HGfritgxMR5nF4RWAiQEFzaXarL1riY/Fiqx290tq+A2GKv8wA3AO+
XmqTZJekgwdwtrbESCqaCYCsupOr0vvbDpKA0fb+9ppOKsXNXLOENg3aJSNvtaCR
Sgu9wq2wC7RnuJZemqmdwNoRczK5qg1AeU/kHXkYhi9xMwFQ2qZeHD4brj98nwHm
DqueKIC7AYMJLE+F4TIc37hidrbHiWJSKYBUcX1nAdlHxNDB9wa6dMj7DPy02JGg
rrp92BtaknWXkUsxzmXYzFVldkWnE9lS8Iw/vv3OT82YRHfJeBTtyu0xzLaz6c1l
EEVaYtbjSoU9x7U0x9fJKB5PLv2Lgg+N+vMzFngvjbJjrurt8Wd6xkAhwqJnWfL0
B4Hi733pkHoJk9kPPpKW8iLgWAiXSISHQ7RZjuE+X+0w3e5ZmTzEk5dVkdbThzUm
AMAeN0iQySghCYsh2uvEWjsm/cpc7lujX2qOuvBOaHMws/PwCFrnygDj35ta1+mX
XgDLZCSbvklMglbiN6DXOdpV2c3txJSVwOQ8W6UroI+0UX124CzWG11Eco84NGEv
uZes4Zv2HEe4I3ulozpvD8xrkyr8V4q2L0q+hYzfGB7zSPY/vRtngq/MsZwiUaVO
I28J3/QRfniieyPusShank1WSEuOA/wTaVN/01nmvubSn83m+h0jDSlnGOHRzNR2
b8865HAnI08hGyqQkqPC+/q++5hSL2juVuWQNTnVKsKJ9yY/6XExXjpSMPBt2owE
Vt9bo85Qu20OinjNVVjmQGMiOpLPdvGr0C8tDHpchoiszjbiscoXEFYrr9wflgYk
tZDJJz+qMLSM0JzoIfmMsfEA/YSuiqs0UF+sG2bltg0K9bQyCZMW3v+93fPjyiSY
iP/+94wg+bJQt4VaW5bLmEkeN2gWycWboJ0T8R08RrlqxIxxT7r336HYxBYnYE+L
ve9bKbKGzlaOr4aqNDrE8HMoQV98tMAA1hBhzIWfx0DK5vZSz0k/NLGhw9Adngzq
ro0VTV2a1ar1EOtMubOYyawSCN/FkwKmO+J1OXPa30/lcTAF9oHZ7NJvTH/ce3tN
dMud8IR5aKP84azWJk/aQ07K+Z6ZTPGzN6rLWkPitxIaXHsV+oN8mt6m52no5b1b
EV0vrh7uD1pmlLonUEqjLHVXLzThKhgKa0FLAAxjMVx9iXTcwl4inGLzCWghGH6Y
b+IFPm+FZxsF/h7pVdQXpvwO4OgBKWY+ZDyzl6R0L2BuHjznMkgpgMPnjLUQIneM
8WpOHO2rRM6MNDPseDy9gaQsi0c9wPYwSos/PSOEN22ZKgqX1ALGZkVJ0iX0ru5/
wUxqfpGPbG77+eQbdgaO5V/ddvsEGd4i21vKxEGEG5N6sLp012TpGrS+uebuH+t4
2v2wKZq+Lm7TM/EPMVcAftVi42tB3raleEo192n1goTiDoGORGdXbHXYL1KEFo1Y
42wRzA1VBkvCtN5yvLxaAqerJ9Ww+xZnDonmleGRBKbJJh6NJ7vS6zXMT4mcktBg
L2SYkAoiDKXTkmz0N+X/K5jIpuZAcSF8jtwxoUC6xW3C/opCs6csLWwkGDBZGvoq
OaDZgFhVItMZyp+vxhcHq5x4+jSV+YnXVEQRW7fcfbyx1rpFA9xrAEXjEE6AfyJV
PzTcHZk+Lfqr0QNeLZdl7H9EDvbaWjobMvW6xgWuGiN6EEYGfFD3JoqIiwQ1oYwy
Mi+X/6wfEQ3gKPa6m8EDrEtUfrQOqnqZ1f30FVqdtQxe+6x5woZHNo3EeuUXq7TP
ndyruzpbjblOweMfn5RrwwVV9AjNsnfZbicjkCqW3YG5fHIpFeqWQRRzBtlW05sY
MXz1ii5Ux4h/mzqYX8Y2IscoC8UqwYDq7vo/BXUoKLZf/0oLBKcQz5FR0uKQiHEc
mfiCv+D6E3kcvvQBTlU4FM7iBZbVNDgcL2v0IndaABmCIRfeYuNZddG9kym4WCqN
ZVkaap6RtTBrus83wfUSehICQ5yIH8vBsfvsR0Y+2Y4gXq2xVHIm/ysVon7wg71C
+ZKSegbEWMbYJ+AjTSc0Ivkkv7HgdIgKqiu4rbA6dk6lDzKQd1Po3i3fkhdLy1YF
MPU2FEDiY3AVNgFoOTPyBzZL+BGdHaTUB/KCqu8M6+qde0po8YSxOUbdXXmNSYKL
EghL+sXJPZBBW4PuAC2Drhf3EsCptwKD8F0t0rrTR3wyk3x6xTuQn9trrxLc0xvZ
1OccH9uIyEOg8C8cGcsXAi9IW2u9Oztqjw/C/AvPZ3pngLIogv7uTu/nKFXcVbhV
GpdFc5J9YsKUzmxrurhtYeA81leTAiMd8PT6zW9tpe0yGxmtLz7DpTL083dkm8dj
NawzbL9uAqEjc3zlZxyuYZX+kWKVszTCqnEaBrh4AafSSQf3LoszuuH4uCpfXzvW
89RxWFFyMwfewq51YC2+MYgEHq/kHp9MZWQ6NWfscszJbwR4YiL0Pm911IA6F/6B
xeiOPJ0n1pLViaW+NFi2uk8i4hdCGRuyzByyXTlMDw+wKiagLV+uBQXgvUYNtdgF
tz/Ld5qENUpkPoP9EJZC6GE+qKe1YRbjkLzEnc4UMSCtoCo+2IX7HqJynPRwczDJ
DxdzEXAD+LuZG+2iDapKatLPq23WZvqlohVMuF1BGkAiKp6hlnpFr/wOVOsHJ2zF
d8qfj088pocxFmimquSqIS6zzi006h5eCLbDm5PgMyvHfh1PgSrpokl/qGh/u4DA
CHdvqjvQJ31+8avhTquMDqmi1bRjZAn7ub0cdMGaX+3I/lQziKlUXJn1Kq61uCL6
LzKu1ZS6mWksNPNVeurP2IcJnoYbHvv2jcH+VgHHKqZ+bHccNT5eswmqZBBDmu/C
Rpd39Qcv3gutSlGTT5sjEYKNqAOIQ9Yp0dLUbHs9XXUbKUEjJZRnOvUTEVn7LCRt
EHlGh7fVLsOSt+hfDqSxY8EQdMz0xNPOZkWaTMVdVwQcJdVhihpmoAIgHLhileGS
8HvHddgGRPVdOok9jndHCcc+qB4n9EmfRzTF5DZR0X7f6k1rnV8y0zGQBovWLFXc
JDREyJuZ1Jom3rxA6BcRerrX0E8ay3nUW3+W4E5luqLTW3gkaXFL7VJMnBEFk8zf
eHgF3LLIL1AF4iy+kbgMPYarygo4zVG6yqOxOOHE0rM/JSfTqoqaY/xLnNLnJ8rf
M3/v67tF39HBrGajnHRZkDcBdjUTa6yleyrhsMidAwpD65ZFG3eb6QZdwHgtNIMl
ShkBIyz8u4db1N92pA1y0yrg/wcolYiA/SxCVv/REHx1dX1gneYQGs/jAdujIgPD
5JRILoXLcXjLYRnHtPC2bG+zXFflev80Hf7WW2hxrxTWpXjrt877tgtfOmrtLxvO
Av7eEDJSy2f41xOg2c09dsl4dv7KD3zpV7bstcTquDzabzyj+EVmAmoq12kvAM9Z
z6MXQGVwuw78uo06WvPEZTX+diZIYiVmdtAOU1WlnIKkNT5kt5d029Ho+nqp1eig
i1qvbondFaEed4lDmBuUhNvXvZHE260DaJs7ViWoUHz5emuPi55q442fO19jZTug
KrDhKlFzcpC4ohPei1utLPubangOevEhTdNigj53CMYZyfe1EZEvcKqCi7XFca8t
O4b2c7U9JwbCCvJJVrzqfF+txT9LG4H2hd01/zqDfZQ6WotscFQh1RGTH3E6VKEQ
s+alAlvfl+x88Yt+1uu4TF6zDUJOxqBgZGBlUhL4zplA2xgoKkl6F4CTBKFIDCvz
nwi3HnhmdjVVAYIyqsBCcwEOpoDX3mK6nIWpsnWLiHEUzGo1ihFTomhNSERDopo9
Zf3O7UmvxOUx3EMK5KiHyw7WaIdCDFOB2yB0wD6TskEwvpgULLRif4+rntULnOpY
cNCBaY7FI+BMUvZNs5CCegtlG40l1wzxCBJMFzYd3dudVawDEWAg+J2AAEhv7vS8
4Fk0Q5YRpbqwpP9g6lCdUlsdFA92r6u8B+jE8S2p6osCUdRd322TbtSR8sYIjP8J
wibIzeW2DcUea0vJIIh363QvDwc8R3o8keia5IepdmivQPnWJpNjYYI8CNSORwbM
+GrUdl0pC54wF5gMVuipgFN5ho8XVAn6PO4fM9cUMA+8lQfdvVa5CKWLz2VqvGHN
WqdsZd8XCFDGeX5ezFgF47n0vfdkVFQ4PiPtHnfJDTrBta9dCLdCO6aQhwkla7qG
1N9ZRn3pZY5CA8k/A+OHLo5EwIOz3jixd1YDE5lyBTLsehxLHCk+/OZ7shcixzQ5
rIXcxLkOgb4byKnFhloi+zF1QyUEEo18zwItSocqHnIW5FyTuKFOrU5k+pNM/1pk
SjA+O6PJDD9paJ93eBtRYgFLsRc4DneBdk/as6mdtmC5Fodw6Gm92spiJMT1K8rP
xFRyzun2+VbmD+ry1Sahe4BnOY82TLRZDAMCh7eDbtBqRVD+0+i2Q70coz9V6dN4
9gIU8ec8rp8Hs5L9KRwwcMua/8Wy9fC4q+/pQ/ckRbFgct2yiG2BPvoVs4xRwBn8
tZcBAXbLk3MH/Dh4V+Y6OGq9wp9bHD696WGL6CQnj6t2sMirBoBT8uJEjapgN4c5
aCnFnY1Gw7AzmqrtvOCSRgCDlSasb8hkHR94l85acS1iJwWfLq6NsDMJzn8AerG6
DBNKGCTBSTwTBzVyNigqLfHXEZM1AXb0TKNkWMrBkLri/SmQEeW7nV0vBqwjwrD5
pJg9LBal7hzeeMfhf95QE5b3s+HT1X6kteJCcDthMcB2oDI7f6iZTYkcdL5FtejN
n2nKvREHle2TWIqXZ7erk/QEY6kdPuVcEaOHXP/wm37Xvx4yg74WGCIYLFyrsPzZ
71ovKHevOhhXFt+ubw1TGFSTLAD6oL3Xjt8xTm2zOJOrnLUNPW96kncY8SiGP8Hp
1inmEPf8GRuvlSDJnIaacLjtKUO9yNgQhK0HoeHddO+sWrMl217xKeDjoEgobyg0
INIYUPCyGpxZsz/g/wcQS+dwZg//EBx8r2r/9KElXdyMgfBrrbcRo4/GZneijnWa
eyjtx04880VdlgpAZxigLpm1URvUotlWEzFJzd7jyq6jQXDJhFZgl9EUySD/Rfx0
8GTdZMNYEdVgDQKq01s2hFzLKviO9jWnH2wcNw6oHx/xeaOY8CcEdx272Lf/cFQ+
4CU0qQWiDOgKpDhTnkJ2FwYP+TMsZQNPAyYM2yfKFZlAqlT+ALbNccQ7Kvux9L5g
0kzN4D6QASNjUwe7H4FlO354mqNh9TWkFj65IWrGk3c2FlgJuNTJ+6BoVv+xxjaX
mtJvYnWKuKLJcTiA6nsKuR9ktc9tQMM9ENCizc3QuW+vsyP8wzZiRobBAtaY9vR3
r9v6QWb1QJ6sFSQvNeCWfA2bPi7sl95INdnYgMwzT+iuU60g5i+Y3/fiEbB0plH5
SCbDmh+6Gj2I8RODF/IVXYgNobf0m4ba7fBHwzSfx4Sbf2Q84bC+qA86K10PniZf
pM9lompkO/CHHjAjA9wDjJXxGfF6jLdzoyv6Eu8dpIL3KsR/n5x/SFmo/frcljRI
sY0jff6g+EZPedTdEeHCHcJoN8a5k0B1hiqwNYunwixuJ6Au8rO3PGDeI70cVrCF
vZtILlfeyZ1nMF+Xrie1Bdt1iD03VowObY4eO3QpEVqIdBypCtr6cS0oP63RNH+H
lucRO+Nz2+GNOhhbBDfowA84i8NTNpZ/5uux9F3rGIngzlOBhIOeQhey7tsyPOdG
szmjkVlCsAtzczt3laKnlc42vqQ3K29MthENS1wvcbS7/YKCLCnTVAPiI/Zyxh+m
PaJ9xZ7ph5SLLAoFNy4woC/B3FxLV1kvq5Y3jGPZ4F118U9+TdNeV1k5i100nAb5
hCuQpUXB24Ss2mS4x/rug/X9VraCx4KNOZCay/KukHwvVZpoLxtXkDVdDSLMiPLN
oW+OnJVLdZIvFJqY558GLBFesPG1E7s9TqknwXIwAIgo1z2vYTiTK9i/l7iUo9fh
YoENCK7k+MFerlOvEEmde8TVFEGnJ0Vv4oEULGhrUH1nErvpcxX90SCQ71wwSKaA
Y4gHsnn4eHFzZ5erFFQ/5i6/RkOA8fAYxaCRSzQBXCHaujL+5jx8TGPYutZq4Px+
LVxeVnGToMihqQtrTwpw/NX///VyeWML7rtTsv70L6AactAzfRsy5bMReUDNQKcL
WRg3+4irPUiQMD88ycU1XQABWIsTzfFsppBWm/6TgRPq5BSF3jMMbkKyzQZKiv7N
4m+wtR7Oc8Jk6j5gkG1F8infCc17/+Wwl27z9L0k2n1za/e1jqWsJ/VsWpmYfv58
VI0EXV9V/0DRslPCTEaPzqgRQgTna2iEoJ/4RhtA7zCf2Ofql2tDpI6a3B309MBd
CCf+soUe25XT1I/1ZjIf8acAhH/twHBj1TsmsblBH9pH2ih9UNzeYy+EhQTn+M53
O/9ZS1hZcAw9sKONDmiYCKCsSxY+WYiuY5zW9cgq9o6edPYi3+rK64xgUjPTG9kV
nJ3q5bk8eMNaiC/6Auk444C3djNYcuhOoZC4HfndrOeb5jFwQk8k+I2ZZsIdhq27
2SnrJhqVj5vHv0VSaweoyNq4BtiJvXIL5NVY6QwpbYK5sW+8B6GOSWVtrv5LclHn
zHBI+5fiZKnx94f43M1RH2a0j48CpSJNwcrgdtSe7kgyYarexIfxa3UbTEJ4t0Le
vG7VftCrzdPRRY+tzWvKuYnLnzJ5LT9z9B2YumhvdOIki306g+OQnqSll3WBAf6o
7HUVJQ/1dwMSjb3C0CMaA8qtLCVevPxRRGcyx7S2lYgnwoIvVzA2XOcgTTFzIHjT
1QgkTJfXa+tcsZFkrCGDZDpCw7Vo1jmJpO2UTkvJlsbQExO0pnZWlqoD7WSR38sS
p6n2bWiVP21aAe8jblfCDqMxfFCSNErvbvQ1oJtHHDisrBb9d2DNw0Y86KV8jmzw
tw2mlhBrL4pBuQG2QkS2N+eWk5bdK4hhlCqlIGd+QRw1rwh8UTkyUgNLtdNd6pRO
QqZKu+HJLFjUO22oPErt222NTz0rguVLVigvhv8kTTSzhppCklk+zsGEwnuzuGYS
NPP2JJfYalWgWKoGGz9+xceBgPEj0lUM//8oOf2oA8j8efs5iffzU2bJbNTpGpG7
tya9aEtVNmVu+pUCIS8eybg3nitJXNf+vJoM19zKILNgeVR0IwT3vHR9IeQk7t/G
HEFE3OTSC559TVoZWzSpgsf379KE3qjmHvKyqe0FGfr7dAuCNVCodCFLHRw0beXb
HfQsjxkIokZhJlo3Xj+kQVj70tLpgZJgUSSPzOw3CDpP/p4mM+2SjJEB0WT6CzaX
GP0GYy7280/o3P1ijAiwetzZp833GKaxq7qUehs5ZDsP+IcOdXwku130VKDKttVE
3QY4nNVwYpxCpCiK6/wlPQ5PIljpk+aiNSvF/6kwmYI4bGIgl3rRM6PbS+gKToVN
7G5df+tqJhRnXxskCWRYQxyPkyAQtVloeVxobWW5V0EDL5fNXwemzYLd7iCVgiAB
t9L+eEAVnicbw9ewRo1UU7ptHJkM0LG87Tj3LEL3gfPFyHqF+/9ghaZrb3f2mMD1
3eozltH0mcIX97yE4dDOO+F6rYCo5s+/8SVh/7im9oU9crnwfpz2ShNb8jLKCvfQ
RcHrB81OOik5MsrlIOcf3PMPQZ7w8CERJcQnko39V3rIsX0CXRZK1C+Gbo1JI1Qa
BYwdKkRjXl5stcG/iYV9E5VT106rb9ch5D2YPFWKoCShiBcuaTmcTKDMTsjZwC5d
+x6YOCFg64i//9QuWleLU8oDVRWx+cjefYyHZv+bYvQlRIUFoz5GpYh3ngtkzTmP
NB6Qw6AwLoLXx6pu2nZ9aL/lHH2Ccz1TVUl5sxObwiRG7vK25wBIwrFQaenWM5O3
jrWoFu1m8jFH6VoDTkZuB7CqvyyKYSxvEw94NO13OnX4BBO5vfYvjkEOQk01vWra
hE1XOQb/mIk0DJ2691TpJ2O1/XPe2VFUV7GgL9jO9AQ7PGjpZpujiAJW9hscOWKx
Nc2hNbauUFXs7HK92G7xk4WxuLHjOt1KEcl8NCELZpX9twvuTgAr0HYJPM9k0mgQ
ydCm272SxXVrUrS9thJjOjF8hVaH6w7nrMiiCDkfifu2ebsLL2M9hjdTMJ94oRDp
PQg/NKKiZSGePp74WBf4U/QtPMG7FW7FhpRLwMX3j4401DUFu8TTlAyfOkPBYRjo
iMTqd5dJ/IsiD3LJ4DI/vqlTCFuzjz4e0DmwGVNcdYCUoNVQqzprTuwIiwmWjakq
nIrBsw7oEOsmx5XZuiuZrjrcnPOMnf7r4xsto++qYRECd2RyP4G94VrNXl/dt0sS
Fujv0FZHYlGUNG/8PGHzbJtjeZ330mNuU4cQzN5yGtp0tQ64jPg5bvWYYH4Y8GyS
Lag5jTfKge0eiNkSpns4Ef05kahLQ78boilAirHqmhMEyELSZ/8U2XHDAfubIUTi
gMT0oiDY8SVpzsFJdWUXNQ3G0gvR9VK/54r60oUO2VVlUcRUQPBonuD3ZTD1Z9xi
LOVICxgbtEGyi3Fd6rlDdMd/pk3H+CsoxmcFD+YE3J+V5HVysC6/S36EiIq4pyFd
3BpS0mmLj+i25/8+WnsE6OKzQ1HKvqRArA1w1/A182N1gdqie9HdHSvMYKE32Z5A
tFwolDMIV05dIc+O0U8yMeRz9G5+eF5jWHNKZTVOHcNgnra6ZUOoEgMA4L+Igjh9
gXSJ5UVJxg4aS6aVY/dsJ6XBfbAwl96/+cAK4j4Y0LPgUKaw/ZSVnBOcssyhY1nB
PJG2HtIxmdxWgLBEn9wO8B7ahpZR8qfsqVHNLG7ChebUPWF23dQ3OfbbmSm78q07
vOpeOj0oomMceSXl7rKHerm32m/0rjeO3EpTUehYSTzsrOpX+80xbdVSZ3R2TSJP
7IP1rr9S3EIQ6JRrlpGc9XBwU0D1EVfgzb5mFtw4MudX3eYrGyrQA4wgGLBk0FKN
7UCIbXwpR49iix40WLsd9iBEYhZyuyz3LJP5e5ciUjtQjk9cMq8kFUs+pfo/7fZf
UGQxFNNCreccNLiW0LK9LyBjbNWZ+sWyQu5P/jAXQfCrdPbICfg2iFm0Nc1jZpRG
gWjYuDdkvpWSvjcg4+NKA9S/S5D+Bj1w+Pr0IG5UjfRDVS9NZ5Osmg+cR2eHVtl9
D4AV7c6wk7gwXyVQKJJ8FwaBuRthjQcTDCp8pzhMMPqhMxEwxfGhNCftvDr3DmUV
u/xuJm/yDkwlBswpfTHjRv40TGFrAiOIa3ndd9Quh+F6WNUMBkue6kXrIe08sCpW
gT7/bkCmluEV66Up7X2hdA55dCbTPuzW43RBJqt7885WD8J2tzNYY6YSmas+BfCV
SMCmvafjvtqw96J2MdP0Mi3/KdRNMJdygrhOnoalRW5Ct3WUtya3MDMmLkAXddFa
evXoV4ns1OW6l0lrICh6DspqN3CKCTXY9To6EYiP1DjNcMMQjB7cyd4sHoR2e6TH
jFen1ZvJrBMYBLMVy3j1XT/P9vrGtXrODDiyBell2GFxtm4MgKm7RWHHcev6CKpz
2AGPPZJg0/P7NaISu3xgzwDCmBTWUQQVwEXPaYvnXM139boenXWXrLAuz6d0x7a8
zKAJLNlPxeM59uRFb3pEPYujw+pe4YJ8Pz9kMveLflmrz1qHFDsBLSzHX+8Lypwm
tbeqjMJhAyF9yIdJmX9rmxN4KH/1YQ5EQBLKlXXupOeVkPU1cdngSrjDY13+sXsi
J6v5O5l91OsAO+0d3FRUgqyYdArWuu5XWYwjZeFKu91Ql+j6CXhZsfT/uze42BY9
4eLibyTZP9eMgLufF+xVCq7v9tILUdZ6w4JjL1C+yUHI74kfZhF9WiR+KuIv2WyS
EKDaDvRkeJtIi2Y15ALoBCCQY7r8h0jIZoLCHsFme8okfDdUpD0xUbhn2jwvTEPB
wfv6q1Pa6ut86J2NZ+rsqwFV1oryDfOoFi2MdTpjF7bBVzPvn7cf+6OFLV4diR0H
wD0+Y2kM+AonDemzbZor2f7FMjT9FD6tuV+E7EwEkDhaZvxFaEQ6TZxOVzHJQEl2
pqn4jnQTwNW/ikg/u3WBohdbGE8EirJOQoonrOKPB4BR0JKBh5gT7yIcXmpsY76X
fQ5ZfuN4jf0V2OzBwhgCOqNuZllbWkZwmPl/COQ0OhE7/dbYPFvUn3bXu3br2ttB
zi0omGIiq0LyUuiAlNvMUYGLjPIEsSnoHW7OKdPqIzGOi4arFx/Z/2+4MDTqLU85
ldvkT+2966v8VF6q1FL7nRHePYCyfZsty24DD5C2AdWL6/ELNypBeMl6w7sbs0v/
23UfTrHqkc/e7v/zxVRZGYN0jWXSdEuPycuhoa9tLAG+dJ3rIOkxez+QMFmnZC4f
Xa6KZO16rCFRd/Kp1HZZy3HrJcqc4RCHDm+fysSv52T8qI6kRcdsn4i+X/+NqZgv
odpfrSdyaHkddOMFUSym4HuK3qs4cj4IuZZhcxgFpGUfPqHng7uNrFrz2v3dxIZd
wZLXJrmZPWQImwqYx9QBvnokylqFZvfM4zrPAE5gPXZhF/4PPdSkQwbUXJ1m+QxM
axTk47bHRJ9hInMINlln8YHPmX3GAtuBsvqVNcuUwkEfRVlkTQDNusQ+cH/lrpeY
ID0mKKoE8KhMInTZruQyYv8f6a0YMhWkoHkupvma4VsKCkdMJGn8eZ20nxhbeP5+
hzExphbSKPFOgsOO8WoftpiB23LghAr6Hx9GbyKCinZsZSkyTJyOUUn+QYaxaGoy
ssLwqZKV6rLJ7NULmjIx8Pu9NL8HnwLjULl+TK6qcbXbcagA4fdboQm3sqq9EWpC
Zj8cHwiJf3x7nUzsvcDG4CD3t+J/iov67w9o/8hRYXBgsxPNEp4BRxMoCYMjaWjG
14m5vJUke/XaBkCGvn7SoNZ9CDe3jgaYX7TZxrPiraCQT0rkuAgJw8AR2Sft38BO
OuwFoiPWcq9dlajZHcpY+ddyK4DnGG5KqzsRLo8CdQ/9yqQ7IvIYzbu9a/A9T03g
CaBJeAAvcX43JJozXtYn3oOXjYpVZ4CZYpMxhUGx4IUM2nglL0We7yvDLWEhOnRw
cqBw9dkAKwRwmKICU7lV1uSzln3w7oKt2L7uwqOfevEjGpH0z2eN7fjmQu0b+zKp
qZSvRFHynjP1HatGs6m4RYo4OWKKjnTml4JHuB6FjYMBT0nIZgyT8DXMB0YLPB9N
es2ffJWv3SwIsbRMmog0Vv4GtaPH/uwhOY/HfcScXBo5+h749yeMFmD1E+sHx6Y4
tHDFMnE9TPF6ObTn6sWPKiPjR9ULMW0UN+C3WMRmxKF9pYmjPpb2Mkt5Gcv1/zgo
OadNkXD40qVDv895mKDVFh97o1llVVuQtgUr7JTI5L7tFVSjIvlvdLm/qulU1gMI
EbbewkweVO8gBzh49kUEDETif72zVUCl0XXt/qESzkGxVpUqfCEMfJsJL76nh15V
YvJ7Jntyxd13cxHap0u+D4jMnarrZikTITUM9cWuUMk5HCc1RIyEXgBnYCVom7Bm
oBkWmPUi44Gy7DwrxRhgOJKqZl4bgaxWiOUCUfgnoPQUXoVEI1xgPL6KOy+a9KNS
/O1qiHtdgBaS97jDf5+eCA1ekW2WA2QjYU20l1Kl1KehbNGH76GcfsHcmKNBclz3
S+ScjM11FdqGSFoKfFvYbgxojyrQKoZ8WwgbHNvayiE7pbsW7+vNxbBDPnC506hj
IjS0XsHZW6YwF0I/Mt0ar1pKW+61H24AX+3+MSDbROPpxNCIiSOUm7CGIZbgfzaw
g51lwTS6njFYZgl8t8pHN9z4Meg9FU5GxeZWiFrIgIjwVqTpGrnZFe8XnJNN1WZq
v2DI6rYPc2pr3RwAnCa1BNzI3h5jW5Cp4tqUC4BWcKCmozJGo/zK7DXhe7pIgwdn
7KHzVVDRh4lQk/sNt6F1mWrJz4e/Ha//wBWYMZMiHxOOkCElI52+v3W1BEK+67vK
kJW7+8Eh+eBr7GPzQvUkGKP18cxBxnVlvSlpKIl3DoGL6EKYbZxvg1bWIaivpTZ3
LE4rMF9QzL8+i1uVIQ406CyMDFW+XXOIm2foXlTbXWuzosUJDuhbDyA2qQxIEHMr
sqMN+TNCvWY0UQd9Krkd9pZN7su/jpJOP7ZAB9NGnnYZccBzdpKYsH/PrszHHHRc
Q2v/SsglE/EXe2TOHPaqF6CMTJgASk9dk5Wju0KQQYjxj2TnmlTvidFEqqYZCqoh
3KXNnOcM4i+rjHKOtA20x3FeYDKtNGjZGR+b3FrSADq7uCCbQpIS7ZCw/o0pUljK
I1/4amiQrBXJniv+nt8t94klzWSyvoO/N+jBBtUccozLn15R12DZaJ+Z30RsGd1d
qULGc2mDC8psNPiVAur/GeBQGr5iBDTVPXQvxrZzi1OEDDj0coEXpBOEgOQuRi0W
zhozH5JevhSxSd0fG0BLQroAd5y3HGZYR28GBUY6Eqbch4TQ0vXj3qVFiJQePk0K
CwjSJEAv/0hLh/IuXUqGv1YECT7ab3CVCfLGn2gYNz5kdxeSW9ccDIwukrtYG6gr
ScJs4ubgcmtGG0BZbXgYtor92Z5t+OfSDaeNWYLuZesXHWAkiLcfWL7gpaFeu8Ud
bCqwGCB2TyjXSFYf1d3/E3L8WPsWIBDe0K3Lm6XSQQL6xLJcDIzar9Wip9TUfhtW
MskyGJJ6iUksmOfWnWFYu2pG8h0f3/AwLEVBCt73RnAyyuASj8+SWRs/dAffdjbl
TY7/NdspS2X2EAUcSsj/bSr2JFcTfP/5vLtH71f90aiWzWA+qs/iWcUctT9s3+IW
qkldrTxW1t4v1ldU04ZFUEflSGtLbY/zgg2gEEqhWgkyO5pRKLpAQDwLII1E3kPi
cHgJs2l2IdFEMRqXU9JuSSkO+VFBBuSMHG7hUDrmbd5G+6r0PLaqOdPAi+LQ38i4
tx4FGg2hpkIdAnoD/G3QEVo3k/saxTB479JTyBmgog6dhNORLpQHRJkhs6RzT5Ew
6Jgk/1ab3D5syEOBfERknFNFsee78dFVqKxKCxix1RX5CixgCXJ/l0TacYTEUZyz
n7VamcKW75r7koBKeL4pp2oGUshD9sIHMGfxgaftPoR2Gl/5cBeOXEZPOL7LXbDE
mYDPq15/M72VNb7BRZIS4pYlEtpZCYyKyTLGmhpXaR4XdUOMMO6PoHExI54+ceA1
gqx8ThVO7T8tA8xfosTfxzGl9bR0U19EtKIx6ND4LArxHO93b6PITTvi3S4CGuVC
effkdKLLS3TqutKEjkCUi6sU+ZWQj7DgiCEiKnSHbmboJ3W0+pKYxm4ukggsvYHS
T2cJhoCRiQeu48lQI6OuMEz8InXEedAHrX+TA/LGeKBDWlDGMZegaL7YEXkBIB3m
2hPP+Ke/O+II8U6xBTnZOTfuL6Yxf6I0iKevowYlk9WnTo311dGzVNO9dqR/vnuq
Fh/5kDf7MOemUQbUm9WaAqMRXg9orEBWyupeDaJB9CMaDu1tzW4yrCNaLRCwkmaD
SdaGyLmlgXQCHciNb0BVEHBcjDn08WHxrWcAfD6c6nDaGOo/3l0WoG0SaHZRaVSj
2sBbmMCTuBtrKg+b/1gO9N5rcqMGKE//xdxCZ7mSbrIN9gyfulBUmnr8Dmagkz54
X7WYV9ibTgz0ZNBuLCX7ESBUvfTlUyqb2mJwc9/tWJPE7TB65SGoXb+jsm2twvCa
KS+JC1hlNYpw811cwN4TnsqGMMElIePcfyknFsGNFoQsYdghZX/YqhgGkuVIa1o2
WZrIomvSntXT4jvl0+kMjsEh0zHnk4Vwe4q0FL/KFNBKNIGS8SQW+AL47NbshuZL
BhDbwufTNyBgvclvZs1RXkNsdh0vtdnzing/L1t9BDy0xILU8OZtNJqnrYAEdNAu
s0/DN/qea79xOT3QbGiMpTTcjlGD96WCn7NCH/2lM5LRWc1PTQeBicc2je/JpIZF
5DyosV0eDRTl4B0t1VfOdUk7OR8VvTV7318ZGlvAilceJTDLvr0WvxRRGh0e83L8
0OkiCzFhKty/J11hOzQ5l8rnocCt94K/Z+y9xKVRjf+R1l0NVorO9Bz3U/SvJ4Pt
12tSeAOztNVia6mqO3lIIyi7cbOeIQ4xo4n2oG7t/zO4xtwf8k0tG9iZTghXoxnZ
K3UoHbS9cn3Z9UuNiC9qsg0IbXEUhehn1ov3ld/r52y24hBgP0j0FZqBI1wrMeTB
hZyKW6FQdyHIqSNNWxa3ZU2kay1sjGrO85TjdxnxD/Yg14AA3d8l5L8/bGwp5SRT
7zTWLwcAmXa0CqrWTOgIwY0DNl8mSRr4b1XPyUxBr6Tvg6imzRVgvGefrQuLeLsh
Pcv9+ZkwaChX3l6kMRpI73x9Q1yBjO35jJVpiIDS3ljTBniAml2Z208JKwSSUi22
XKesw6s2JKiIYy9JVKYDmosGufO4dnp43SJcH6zH2FyrFFlfnp6tNax+lNXyc4ne
TMkKwUacxjs0qVrlRYrL1omgyOrYZX4Q08mpcyMUszCyigs+x34AFA7kZfS7+2Q7
3NnZynf+Nhg0+cZyDU1eH+5SXO3zOz7MaOPUbg/LTJSW5gi4uXSdi6b6EYR2D0Dm
OwV/Ag3CChEVbyKvP+qCdLRmwBn+eqYO4OJYtnWgWYwK9Vl43so1D/qomCUc3xTr
4a/vAJndrHcXz5e6pGCmFcTVsBfEbrRA0vNdo1Icu4srhXBrvrAFfTIdnMymR4jX
6czDIcESKiWn2wgVOrjTtwExQLYXvELw/ITsKrpSLXt3stBz31+DpAFNiaGUF2wb
ACFtgO+cJofRWIc3xm1blj0sbgLMovV31Zew9Bpll/z3ItZFXinK+eXwr2ma+JMA
IYbgpHxcA02XN1vSpfzknQANLYKFjojkeWPAWxZwCJUxCJSq+n/ewEAA3tC9Noyg
DwvrIxG8aExW0GxZknaiDKWq4uixHgWQWhmNA0ooUBND4Vi1/uUCpu53H4G7k2c6
2NXpaOxYGUXsUGdft+bltHgr9kQNvr1zSPksaRtTBsHp3Z/JcPiD/PkDGeJuKmBz
9OPu1Vj4f2rWrnbQkKsBOuACxzB0E+nYW2XkYfiwCb7lawouoOBkEJyKROgcn80M
FeG4/qyHkzuEWRAsVWVkPUbwoaCcXpizePVWXJW+xY31AOXbcLQZDRMXslQYyjbf
ppvW5ckUvA9xGJhqA8FxVzm3hLI9XlmNoOT+gdGLxb02plcbG+pgTozI6jVLyFHo
sNQTLZLj3xQVKbzcs9KMggpszhNkfNqIMLSFWBZ1pdvO/oAD9XP1P6c1LthoTqYc
L+REahk0tzkWry3sXBbLBesPStkBh3xblAkO57LlO/fTSx5LSVUbeij4Lt25TRMM
LJrLuDAt4Q9mpe/0JD9F/4DADBNu2UXWg1EiUfqnjNfkyO3cfeZClnbcAjGlpwS/
rq5Rs0+UTP9FB4W8YICXpbaTRwBNmeWaAPwnt+8PB9LrmjCo7bx5blH4Rdpmfg1b
zSOW4t8zBLjGcb9fJRZhcAVANY5LXgdpkI0TWN1PCql9NhlwwA+EzC7QdV3eog4A
sAuoTRnTSSmHod63+n+qRrm5MasQUeNws9RA6BcuBI4kLdKGGwOEKS6CydEwNnmt
Nqevy8Tx/XJ4niqLNveJAeifnHtCAN0eZ2V2JRTAk1clVFNZlKIv9D7uZHKrsxGo
I2GoQh+0BkFxq100KkicUhh8zwkmH4KjcsKAofvGDjTLcVROplXBG3suvM3yYHWS
BXADSfFkw7VD/mwPeO/YUgYZMoUpBG4Z+cC8CJRuZgP7MuENUT3ZlKQxypu3VxY1
mssZV2IT3P/8QuZBEa2Hf4c02mGRdvGRaRZYccrRlbQk9ikvrGYJ98CHMBRmunHS
vg3ER/lhm26Er5yPnAxF+mB2JhKY6N5aO0OE0KPZag26dld0XxwiVtLA3mSxeBvC
eAzaYdEOdIDlJ2G7cFQ6rC21ii9kGJJ7Qr7m9C2dCFCfmr0FL32G23wfyUIbUX7l
0bpsJy7GJtxb128hpeds70/KP2xq0ePYoQ90ePhqrpY3e3ne461gYFXAGJOpfjdH
6OT6OOXjBjAPa19hBchwY4ex/KUvQpuhqF0ewTDe4zv4WZaqhJGXIUPuKC7ovz2R
ZWdLV59Cr03mt/UKFE2RE2TjQGId2qVaUaes3KwwmbJLiHlRLk5sE2+v7DvwqyAj
0p+Tf7liCyVF29JxNb3VjyzupPoB4BoJFtze6Locu51MejH6iaTocdqmoWDdwkLL
zvBBspnzFXFdec+gOJCz60/anty38iTC3e0fd3fygGwRcBRfrdE7OIRS5pNnosBk
Zczm5+9cGV4w4f46U4TvE1JhBVLMXJWpHVTu6r2hlFHkzzb4XNW0oM8c0yM4bIE0
Tn/cLLxrV0AA7EkMQ866LUt++9xngCjfJDS3HGzq2kvcUby1iHmwdll1TGIC6OJs
Jdc0PcdPz6xGY4g0UQNRU1PBzLCatFjZ24SHJwZxyHcfGAUkiAMmOtbwimPcDreI
OOJ7PDZanr8WHpMZKDSHYE9kPq6LHEYAqzlyTfQvZS/Pa60Z+Nl2xiffKE49KE7X
87Tx4mbRkg4PP6e7tozbcHKj88Sz7bOW839U/ksBCYtbWw5OmT3ifYqRlwFAgxWY
w7UIXPcKgABHMCM2W5Py+UEHU0Qv/l1VREt6aMv2BrYeGg69FskZoPU0RHDXlBMI
Q9UWvvMe7KOf4s2pzr8D8jysjyWkcfHwbk67InO0+M7dBLxwy65s+VYny6+9rako
IaiKOyhm+icfY6Yn5D7O9KGt89NcXleq+j8CPa+AkGMjKAc0+CExVXcXseeusWcb
st71mtFFh/KncYjk5R1LCv+sFUQ7CjuPWKkN1hWTOcVCcGJViMKQjFMGsTwqBCh7
wVNKDptcP5Pdms9AyI7VoI4UB54jwMIfZ8pB2vjU/Wi3kCHkYmzK/8Kz8w6hIJ4V
TGdMOSBthfx8p0HeC+zwQL0x6Kh1ngAOmiNCgFY4JakznHDyhgG5cvoqB0ofRtrY
jyV4eVH6Wmi0dYM7+awPVjPa7JKht6TMb1eoX0HL3CsEd42z3xmJxApldZl+1Fd9
2GoHf1EtxSylyg6pOaDQIe7PAFrrDcWg1gCoWVVM/bYF81M0PJS1O3bzAfx/VJJ4
6ZG405DW2OkhoB5z0ea3tMKS967yNOlTwfd2vhxJR2W9LmWXr4z1E7n3YkKnYqAI
6Ix4BeWSWMxRnBnyVTHJ3+qyUW2qNTOVUL59allROR4rHsbiMenuS16Yqjc0UY/M
FR2hB3s/uw72/FOv9XzcV20tIBBU22dkpl0+hWHmaiDE7XXpIebKnNEFZmWN/jgd
pkEfeL3xUMCSFoC/G1GmemEx6ul6eBAe3vrBGIqgJ3rFykzew17hYq3wuOUiDpc1
8Gt0dWM5nA3QJUlQngrdDaICKhc3Er9QjhJBNYp8Kpapr8USCRWXeUg/7n6E+xji
FusJEr9phOutSmXeVwd7aZQFaKPfqUyNZsNwCPUT2++c3LAofeapauDM8kVxCCO0
7o0/sA76u/ICbJrvB/0vpANGFusQJ9ZPwC3+520ckvnEm3gQM/u46zdUrrEXWxi+
m+0TO8e/O2HLX4MflZ+VCo883SxxneQCy4F7JGxMQytK4PhW0J5Hicj0JbRL4h8M
QXktdfQ4gH5SuiPH6YxODSQ3FOuWkdjn4Tvqy3RSMz44JQtavtLtZ046eie+XeG8
7dvSrMGR9H/3bLPtyU6V8TvcZCTI6n57Wjd4fvUZcsdmGCAg5YiGFMC4rzIs7g6Z
z1JQEAja2WSnAZa+fRY4Dn8ve+HyNvLfWQjpkFoOWXKtZB31y65YcfHZX8JgfanV
rXQObOiAn/eZsF7ZqkV8otJZ6bQLERU97IVnAh1rK1+bTP9HGzUZOofQFkfTsMz0
IAU259VZBsXzDV98Wr4wB2X6iXN/nrZYu8xlmjm8puFlebdRSGQmhYU1YY0T25jB
G2BIT3prGDMW+fe4kkV9V7WLd3f79UE9AF8bOTVEWShVFRLb67N8P+mSd015LcW8
zL1xYenFrUfpf4TWk0ZTdSdaognDWju3x2Zz0xk1iewCI+XcVmw+PuDztE0p/U6d
/YXtbrd1UyI7oiFQhlvFCuynDfyBwJBBeGAvj3YekE+7C+4k7URtc//hSK4ThF1C
5VmOXZo1VEESF6hBVUgDyi8DW8gqHjXa9d6Meb4VgVL4Zdbn+SsHhUzeKLU9JT2K
WnxrbSzARjlbYP69HrwBL7yOqJ2Fbx0ibToUtaDF9kEuL4LaBDiuiIy9cvwL990+
I0XfhHbfNlqvbyIQnYgUzymS0YmHCecBOw0aGRmfV42pi/VoY1J81NylxTPfDk4P
xSpmmUzWzoaDXE3y+b1zgloo0G0ujxmXrBFzeGSp8KtX/vUBx0CwbxynHa4wLJXG
Y4epQtA6yECYltf9Tv1Bl/GyySoH14j0UtgFtxk485ltudMD+MPc7lF+NcISs6V3
D44SBtAPRTG8B+s/MUaC9jkrBVQyT9H5c8pqXDfWdyc5gKl0ZiYr+nS8Lt8Htsct
XRKA17RRS4NVEU2p11FT+2BjaBOpcl9CDuxCUda/xXIxrFB2Kf97eemgbVVET1vz
SIiw1irOUiKh6n6b5qOg8yNDEFZfokM+kzpYwOwyAXRNoJa0jQD7UYKO+nvtgfEH
4/gFcffBMVDSTyaxT23lUXGEY6YxefZ/SmPERcUNpfO9SJV0ayxdv9c6IDGHrr5e
AZdAH1n+lixyhd9ZAowm9rQ6xD49gSmfAMucpgP3d0S8cU2QN02s0xbWJW9XoQ+Z
jPGqFskRGsHSh2WlyKPVyyECNp0gtTgS+dQ1EwakfkaD6Fj9JnXQGevD8WsXptLe
RQ9ePBbtGkVvvd9J+WXcgmngJIw75HBNou/otx5vvU++1yT5zwhgMfx1TgUzenmL
FBSX9SkbMTa59iUwiQ44GEk50qrVEh64ZswBUS0uVhOrmSpHxRNQLwVxKtSasDVA
z6dJf35p4m869PVUKxuWTBc5MGiC+X6uOrIpK+gbD1yObAQo3ozWOgEoSxQjZuwR
3tXq9/iDIskbPXKOs3rMS7aZ3Gvfu2+a2wYgX1/a6h5toqPEEOvjHZO9cMJr+lR8
7BtnlFqQoBwnpOCarMguAuwqoLfKMw/Fqo1bnePhHr9lukXqcHka/tnGB7NZ4OnA
PWep3AsndoLeVZEMox74PN9JM2yenza/dmThdaDkIxKaKlSLzfjVMQy3rzYR4rBd
nc4TenXgywYOrCJoU2laTFGT/ac5Ja39VChuK8LFEEnbm/cmW7f3jevdzsV8hCDQ
G7M9Jhh4OUsUmWo74gSq+OlMcwtoyJ4JaVBsHZLe12fSB1vQOgZyibO4WJhmdW3J
Z/u7RusiCVQoJSfPilG+CrV2+x9iM7IM+VpyDRkgOtIPy8rH+JXMU/l0FKsS3tj8
af0qoWykRHEyZnZJdYsG9GXSGGqdaZq/WyKq+qoqkaxkb4gZkMmwPcnI0go7OXJW
hJ5bSqCHcl7Ug0Hy//olU09FeuBSwRW6YGsefyQ6gJShstlslKc2oh3MxRbZUzhb
FSAydFgXdWNBaiTPBZUKZTrAmrbArZLOTdW9zRhumISZMr8g9qJq4AjCQ6IS6osB
EsyuGsuS5+/UvKpzwJNEW6K+W6nIzc3nZ8SfWqiQKGJv81YUx8Ffk+PekvK/RwHD
TEczdYehCu+jbpf3795nAAzLKOQNyTjDuFYnawV4P5OpKGWgpEzV1z1/1apJQUhq
1LouL7xX5J833kgK1bvk10aiFHH0Q4qUVlQCYKx4PpFJfUpIXHjN3CVQqTT3wVhK
rTa3xuV4s50A5W3oooyqRujEiblqWp5uBy0lgoA1iA0ZWWdd5TyUxB0+Rz0jv0pS
MZL/8VEZPsLt8iYni/45EZuafWY3NEGm+7a6P490BpgFBerrCvhangIASn54vaHF
KWOFC9Ihrwy/JlUxhf1guW5QoFED7jc7Z00ptGZGUDYPlDbR057I/Pm4ZrJfrMJ1
Jpw7qV1H/kdlbsi2nYPPxGiP+BXLWhksA6gxxjIEJIUqeGk/OyprKZ9DzFlXtD3o
lmdruprGSwe5lstYn3Q0sroQjPF9UwxdHN/QdsP3WNCq1XCW8j2vW9LmGxAaNOOD
E6g75ey7tyYkCGv/fYUxEJMrnYoyvAH64sCPq/554LSqHCQfJgV0zDGh1ESN6KUX
lGEoL24PGBb40h4w//7KfZNwlH4tstaLkG/SJwk4WrmSfTSSBrrk4DPSZL48FKmM
+k0lUnwPWs2+306rBp67hYZPFOj5w3vC4o83Q9V00szEcr+gqJCq+G0ty3IPWUfN
Os5qYovRJCsR+oZe9tfIgCMLKM272DtdNCgCcXqUbfsyL+KmvCgaaKEwe6r/hFJn
Bd1Ek+4aUe5HodqMMSOVFvRjxybozTW5Ftkf8jPayiY0dALdIInMtwMQNcFSkP8/
vkNXEIjeksF6e9lXzwqLO62LkikEcbm4FX8u0wlKeNI7K5tRB6OiMcuOonwMmFM2
BEiVt1yv99bPCMazNAYSO+nfTj/VH48d44yIPyTTVwUXf8gnyY4rORoUAmMonRpi
VqPm5w01DsRjvux8uY8LhpJ7CtEBZZZRWRXEun4qb6cEbtLyCXDnV1t3v3MP53K7
f4I82jTpDANMBITncOFoIaj3YB8NvNiQAi6hJOQOq4DdPGYXmJxQEF1oD3aP8FRS
pGtInaxgm7pq1uKhSZSJyPDFo5U4FK7fIPceRhy4JpHOOtOg1ouk7RVCn80MK4f+
1C/YswSHuEFL7yzuMJblDP+dpuHqNqXpZ2u43f8gXkCXDBNIZLBiwi+Nc1WAhAvI
7yc5NkOIUxsHn69gWdasICJKf2FKbYjz3A0JZIyPfVUB0lmYP/1bS4ZJzoOmfP0t
ytkky3njde3SiT8mxEfG4689Zy0ZQ2ZkXtQzwP/FPkWvn6EmPhsWPEEmITUoxK4U
uBk7L45KENvddsDMotyLLITRIOkAHkNn97A+rET5sv+PzTuOfWwvH5aM+FhMF5sJ
CWc4uOLZbYX7s8XJouVCDrb1PCQ06WPn2R5Tgil9iBvufk2CKBML8Db/MoKrp+FC
gTgGTjgUTDyX2yPAzf436ghDqWvPJhLMzcbSGYtQDqxwFLB5y5B47JphNwXW/pFH
eWMJwsRMuICIOB11LIrN1vuA7tJQYUUCxQIu6EJBTUjxzDm3pzq1hA1yc1FEW0TP
jnFQ1eqlCxhG7ZdfbOYMu4frcqKLE8barhWsoOIb/SVfkJF0EC9JmU4YYpZq+1nN
PjyTd/uUKUvHRYR6PhKwKGhKAIgD+xlCsmiN8Wq2zdmHb0OBKclJJXAIznmG4m6v
unZJyGz794KBfqTbfncgb1cQqGsOu/PRHsIOFbYJPt/aC4+ewt+6fJtYI/GehlCM
Njj3UwS4DI3Fgm9zQF3M/9U3AhwlpDhyXxu4AvKYZFd0cCM9QSvr6rMFsI1cKcq6
oMIq5HQBbghQ/TbbgoSrF7bQaS6CNKzl/6AiGan9uRmyLuqwIkqXfF6uxDpZOElk
cJ5LcPiU5oPsByaEzYU0hnbsiLZoqm3wl6fiB1kYnUd/WsNvWdDBFlJh5ZCQntd3
aCLjfcu2lLgnTVLd+63LI3Jjhp2CCYxQrJn0rNsW0OEzVX+CmDu1/X8/2ABBh8VY
mKVLx6SyvWwwmGL4gbgdRFOcmIm5XEwunvxttX1w98O5uzC3IPlrtsjJb+JW0I7H
GXnUKZTvosvOMR7ynOj8mnSWDVbCsFujI0beIfDQYKLwoSeTsw7SIahYpZC5aol0
91T42RO6KcffvAtut693g5iAIrXg9+rLpmHzshOiDB2nGian4EY5bBzi+UBSyE5n
U48NbgLEXUB++XcGmMA4cRPXc083xka5l1cp4rqwx/5eQDujF0kM01IrljkWSBmC
fW2a7IcItM+cx+DlDucRmitCTGGF3Syo494mj33QOVFga3xUeiiqBMBRDnFr3GFp
68acOLFEPoYAZPMYMFKz2IFfpPaqKIExgX3CcKIZPfO/FGhYzg2w7Df2eIL7Nv4r
QqbIeITun9S4Zd+A1gdLmEV9MfFmkfj7gCJkJCqSPW2QD/RbjUUMADI/z0Ug6vya
PXedpZQ/JIpE+bMcmg62cnV5JO54Mi/Mkjfed8a+ePFvK8sNQcA1/p7F84x6ETRC
+z4S2gQ17ePffnsk/wLj5TYWRCVLeGsi+6q2rkW57lO3cunMcTy+HmxguKaYcAwm
Mw3xbL34qi+WjoTd5rY2OOAIcPPUIghsmPKyOffJYhsQ99YX2IhgU7QKk2uYTJU/
L0V8Z3gcQPZRkoXhfAhl7rVPMlQp8L0Uw2QKlK2hFtp/yFZUn/vPt6fZ96+PcCav
RF+BbRm78o40LMrICCpPHGKgJWba+YnroAhKpCsAT+UNdbz9aH3fa743UmY8fBsP
IPmzvNXP0AARq76To+clMduxlgmNgmQrFk/ma5BFATChvVAOJiSDtGAXF+QXrG1f
dMM07TIc6YZXVIkdhCdApG9uT4mQbHYDk9/lwfQbxfUqaw7V8FC9xx8Pv1Bd1HRW
VLcVynWsY1afj0K7CjIJpsAgHxkeG/o/Olqb3qsaXu+GT15DHO9MTofLyNbYTLil
2gYNa+0SdjfSTMfHLbhHlr5OmecxQZcq/FeEcPS896ZoeoAc0vMmCNcOD8gguPVH
17ZK4nqzgbyLEUV0RcZebu9wdQBLXa1t+d5tg0KTdRZ/6xwbmTULKYoEE0g+JgSE
PhyB8VbNeU6XaHh9o7w26sHMLNJRLDAUV8FMR+CqSU0cBu3NCnN0/UrtBQVdAEkZ
BYjXIh+Wr9r9WmKVhXOmX0taOHCZJe49rcGRUDh4eyXo91k/v4lxUNZJBLrM6oQL
TglOscRgHabFWhPyWMDbfTtEkA959JjQeD87WuKFGcVc5P2ys6FGkrNWENIqK3Pe
dsma0LvAFe60eTxXInF06oPAXOAi47+GJbP1FjtkaWndMQ4gRh9HV1IPcYPaD0S1
VKePBUAony+mfRHHh9xbZh5QpLVzlWaGo/5kP1bU2uEN0jmI75+c9XmxuCxK36p8
mr5XEmXmPsoAJCQWfPXCauvJOi8l9kHXVNT1LkkRBYU240ULm3m4GX4sbNb3MP1c
MFwWVPpiaeAfBjGo0dZ2DnwNWWZ3fuoS7QJUi6wGgL/HHXgLkGRxJRqxZEizMKtG
R+4tLxq4JT7zKitnBdkBL4PAkUh1NoZYz5zSJj7SIKwC2wUOmh4iytkqAemB/5Nc
YwDm18qqA7V3fKJwJ2bvaayVx4MFJPHN1VDFB0Y4/4Ps2G8BsDz8Se+Vw3nWRlPb
/sFrab9pAMEuEyIWQA2toyXJ7ugGkdR1BKgZnviHKkKN7YlX3MHWVBfePP/f45U7
kzPZBTNSB+MiwtpMPR06H/wsj2K2Nq15l+xOe4QhtZs6qqlfe0haOta7Gtm2n0+F
CRXwrfHrHadp/+835kbkN45ekE8EaBRcg3buDjl71uaGq4cEGmffSWBeBZm/wplY
fkT/utWVliZQcIxltFwiAc4gP/PKV6pil8QlPiPvFOae0dBoJqfxYNmq5HBoP5Rw
Dv3aymjh/X0k3YpkNlTpL7SKz4eA1vSWBfV8oCC6StuO/BlJvW348JzLVYaeCCEl
oo8wmg1Jwxa0UlFhZ8MKavqwcBtz6Dxtwgu3XibHjL43KFQ0qB+4/cM+/3qT3D4W
e2NJHTEFmCOhdzDDG8vYq7UIcvpR807y42tDAU4kDnaYwOFpmzyWzBBK/dqOozFA
bTI+7JprbFEfK+pDqc1TWZlG1ZzSZ4AydiCZIkYP2oowUOHJGFIcORhfeIirF5ls
BJU9KNWKkufvoYTDgEeAgmdwlKicrIamW/y9A9TyMN7q9g5hJxdEi3gqirqMTOqf
Rwsy/T+pOaN8yWuruIf91pIiGrr2fnOAqFFwmIEgbozr/dGb5Y8+J0CfDDVZegRy
J9C9+0q5rYNaZvBsSX0rAPNSS102ZIGb1vMxAd0vRyV/PZouM3th1s33uwqTGwZw
0sPuPRoes+JzYC2GAJWTFnrwuCMDzKB7Tg4iN+uv2If0eLSW2JsfeOzQd+cav7+8
ph0Fl4iWXTXpj3Jsgbt+Yqu8CRXGhO4CqSdP+qfx+i7OKj1r1jMUUJSaK7Db120t
w8C4WW8twAxp/rpdWP+WIwTLRLlwfINMoq0ZDnKpeafPr45/2zo15Dd/550FzMJb
jDsPXastrj/RkxcqOw1MVtZaYpyfFsAOPpKWteTF2MmCXzcKKWJ1uGbrjwb4kzhz
HtYlh2UVSqAu5wywP4imXz1feara9Lv5CwNZ4H/9VmRkdBhnp0Xq4fTzTbWrkHt1
ZVm6AkFEigTSwmhc8HuSS/vUZ6btKqIvc53nWrXN7w5JUGasLqHOWshxkdJg84rb
1lhGSiIytFJh46h62qVWD3xN/XKG35C39J7+x0I1IJEMd2xKJdJgM2WDlM/X3UDb
JLeqPqeEgkLIAMC+uShSx1L5nBGOUe4jW/AE15OWurLJOjZ4D6d0LUOvutuhiE2X
Eq0pAVrEuXclE4nITmWe+AMEpgVDwOm/tiGMgQ9EMm0frkfoYOKpo6itQTlUmNsg
9cuw++gBiVp6vjmjHjz15zFHXeP57A1yZNDMUDShNR3zwpa3H8ULiHKchG5dr8td
VX4WZS7ZXxhMCLB5CVnzN4kvGXFZWyCs4Ke6oDV+CD7GtzbyYHKfXZVtu0vgl85O
VGglHGgGSC0KiMEEYuuDeeYj1iwcVGlWy5rSFU49OXnZPSPyI1FcJJXhJDV+6e7d
uhZHVD0ldTkXH/h2Ork9UC+ft5KXYzQnXYNgnF5yfwh6B4T7s/Xn8NrliSJfJRqm
ymgKMB/EPtn9TjOEwL+hJRbOX1cs+2zGwX3qqAVvADuAtz6UrVtAe03xgtZE9QOU
52VFoSq22H7FKl/7lZP5XGBnP7IYtPchWqoSfsfZmiTHYTWoADpEGwMUXDzNwnRo
AzmmhC7eZWXa2CRJaE+7GaX+A+lSpaNqk88Kr/ey8jafkXWs6oMASFuMyvXyy9wb
k7e7R1Abb8VFatwQ9PL8LKfaK7/hZYszPOnR0jn8mLGC9V2o4Nq6sc+f25JfuteC
Mjeo7bSY1ZAVEBjRziuTqC4NMwvp8zTaUq7pVfcBbYKa7iV8zc8/CpWC90wOcG5s
/xhSKBo8OHtgTSv60h2mFvuDSLKDBLAp7X8dy4bHoada1PXFlKDXshAXnSwHsI8e
lfizd684gzhbBlx/OOaZYshc+9r/QQRD+pIt/mrD55bIZ1twyPJRF0TCq2MqiTgV
CDP4KoLgN7sG/aX6Jrt2E6fbZAP1kHSaYTVHmPZu3wO/+ympL9g+AJYmgFCPVycz
TzxjAVbVwGEqTlO2atAVJ/+X3v8MC+jGvtp9U45kblACMXZ4dU67mggvf2KaJE7K
m+ePXZZ7rRA8fmO4TlfDjbJgVfwe6L9Gq3AjBl480HLSFRQ9YXeaU7biRRMaSase
nIyzdqLWh+DbD3QU2VY24Po679J0Rw5wfzcjrtTohJASHN2E9p+8HPb2DGT0CWwH
iYjcGaeYkfGhwj5BaiXZNp51+tSStG6ukxLPUIociDconVBKIB6J6MuojHTf6yCG
f5mVl/3bWfw1Yq9VU7+OU4eIPXt09JbvkLhDFjumuiuLJJjSeEJxkEeUpJRo7JIW
euDCmKWXwtVaJBcRdFl4w63p0bNxKhasKD++15f1XSsX3PMeTsIxKS0T12TC1cAw
wXbHum7mr6hfplKTkGEWoaqgRO1kplhxd9KjkbMSjAPfaSXkUOxxktPj16YZC9TT
1Nz9wojZuDV+3K4C7m4XqmgH/zpqEg+0hrCoJrU3kJrzcuOuCAb2SXo81JXMEN7Z
qUkRBH6a0DEMRM80XPUL8eIaiMY6MRy+8jKbfmeUfn7feVBcPMjV4hHrmz6uAU9J
w81CqkFpc+kQBNc9TCxzBtoQq5pSpxf3R+ZwX3Hd8WnFSzDF/mxOqZ8nbBr6D0F5
z+ZSL7/0Wcc2hL/Wpxw92dxj7Q0XtzBYH8wy11+/cgSJCJX9xZmWIZ8wDfS00Vmr
rITLMPYZGJ0ZHautauzEsV23M2ShqQpzjpuMYOzl7Y4NOujkCgO9l7TpQIcS2SZJ
2t1YrtnkgNIiLKDJWrUpnnoBBbf0kWPl08FIlZHkhsf7XNrStlaQnFofn5ksoe27
YWA9dlxTDDwdDY2QDPiR29XZ58kw2tAYXSmhtD+m8yFxfMlf4g2EDDmlK1ccmZCo
InaPBAdQbo7zp3hMW4qmFQcDDWSRenwWDujfkjKafTW5Vtxb7/q3jJ9hd1sr4Gr5
l+zBk1Sq6QygkSEX9l4I6Zjyml9L0LIw8QiW+Yraouz4ZYuSodC3h6pBh2lplwyX
ODIGEkLiMFjZ52twJ5MeNf2dL69mpEiz89YBDXAjQmt4kgDXwLRcF97XMipR8gJU
Astwft912eR1alcDAoP4Nch7wyjxaKi/MeX/V9HylpQ4E7wZvWXl9toXBuiOFbtr
KactaoS4ZZK6vd8OeqR5cPgOE4W03bU8WVTo0lnbJPh1tKsO/lgrV9PyJLsuD8aa
uv154ODv6ZNMoZhnmYpB/U8vUGeyBcMfPT6tK7Q9Sb/IZJqNwSMDQ6v/ZxckwKsT
mwluWRm3qHcowQsPupt/4lOeKOOecnkVt4XEIN+3odDDBc+pwVkPKVFkbCNAQVYt
WdLknsllMZ1JTWvM/a6OGVU/c+RsMaoi3dtitON5xJLjMf6fnHtnrTs0BuiWGIJh
BRNNcJZP6M/ixdTByguRL0gG2RsSY74d86D/3jMEd0RIQT5AoAYVfQ91VjFk8Ji0
7/njj196gVkpW4EnN9i6JslMceBEYyA/0LK1r6U9d3dn053A3zanvIK7ZMCeSrye
98bGj05Gzn4aQFxJIJLybcCQpU4M0R1KDb0uUDWUh8iY5zyJLF3+CFpjwfPIRxBV
DbTlK0CSwuUN6R4J6j/Cb/cjFwwXha+03H6ovo8DBcD+4gJbWbXIDxNbjh80Y61B
+TzYkiBwYu3u+YCDFtBYYknng0xqIRz5UQIX1ZT1PZ+86NUo+OxMOE1DnE29DTKs
hTkO6c5g+Ec+HRrARS3UurM1RSlMvFQQb1z8MGK+QTkyoEhvaCYab9WCoedYBbve
ljnnsfZQD6SMcTtmwykne0GEmtmN62+S0lfJKrkSbH7BbkwJOxwuGv5P//jB6ye0
rENzdK9dTyvzqij1VBbc6MjpQObAlmMhKJ7cM84q5GLhEAV512WsG787Golljp5S
M6FqEyzzqMRxkiiA6Dx/ln777PqK/4VwNRf7IFnA3qCkUy9T95+11xPSnEtuFI1n
IIYpM+aiDEfQHeztNPzH18ztX6evwRW5B1zgMTis26ce6nkYKdXjaubE8WcZrtZG
4D5Nbvhr41U8CAOf3ofpZOI2v24yPkzyBp/wjPEwGveG+BRTKnJul75BxckCjb2p
tZxat/u51e255HvR7sM0rllg4sRkR/b18NWZ1LMwKT7gsAIMWE2wZuWr0XslWKE/
50xtXRV9K0XuRi3KW88CzB/Z5IwdB5pK1TSKntei3LLo4JAfuNZNwtyZfY5g5+yz
mr5iP3enO53oiZ/tfJC8OwH1oQUcGIcMHPTRkoJguqwSdxs9nY4eRbI2KYeIcuLc
CVmQU1UwvR/J+6eKTqlBZ0yxcmFOmQjlKbaoogcyp36b+gaAo5JlkpDqRlUd9Vkt
2tnSGdE+HLJ0kJL5KtU1fPnlEb4UuVCrkJo6EsHrmvXeyA/e/3nmlux1MXyoZ66O
pRRhrXfa92FrPuj+iFRtr6qBTvY6NuG4fov7CyTrmjGvHu3uHuLOXRN0kMvVtl30
5fN6vbtwQrXVo60gLSj+0LglV2ilh2QqWRQIfTIngGzvKgEiYCf5gunwYeMsG+xn
IxughJhgWuzfKrr+4s4ENfTEm1EEZOChV83DoAsW72/8/FFJ85A3Ro1iKE6oYLSP
6/rej1B3qKUQWOuilW35BJZ3U5m0Zbifh8yPMYc+OelaLNaB/Y/Gyph54bXK2DLG
3UPhgVqLC4ALisKUEWbVVJJ+acqy4TH8cXMiRcc9EQA6IyqzorqcC2CDVp3zDusR
yf9KVNw/tw7Zi91INHl4k54tpT4JvTYKcCLDYw9GyGmSwV6jxa7QvixIT3Aw1BW1
0qkPFFruOuylkirbB29easVJKB9ujlYy8dYgTk1uNJqs/3Ubk3GXQTcHimCpvoEN
hhfLboQ86wD9WSUbxfMf2JwhYRfQTZ2I1JiNpu0kSU97QAIKAXm9A+tt9OcSVqzm
8pmVbg9jq/MLm2Mg2JGXwk0gXOxZ+MvIE9Kv7FJnqCg6+FRXZXnbOjznNNogGrd2
X9Oldm3oq9sMzARJ68Eff5FqQovI5WV1/mrpVPyhNVrC3RdS+pwkO4lWXiNDXcVY
R79DHL8TSiBl1OuCv/sJ5FylJb8Zk0rK2i9tJIHUxnEbv0hRJEeK8th6CbZoLUQt
lh8pCLvt/wEc2uf6MAHPE2b4n0gbEOMRdVcl2I8vwLqPsm/G6eUsA5r3J8GgsJLb
nkge/QBjCtYasy5JIDoar0I6ldWeH6GEtTk5ccuXcY5gf28Bc8MNBZyBx56Y8P7z
Lwt3rW8h7vctJJFU1yKU7t0+oHELBJLxVESTFM/xxxMVOwXGPAd77xjrHSNdF8S5
ErXafSDVr8frpLVIsPKz/oj2OiTQNK+n9WKp4RRpIULPP+x9rTpsM4LMTtY7DcsM
1Z5JEsB3ZzbtBf1B4MM7cTDsvuLHA0cICGKKYVfGLYnKqODOsi/mJARuBZBqGgKB
RWK0JVUp2l2EUIle7qyCYT54Ipe3TwsF6iy/37wZ0s4j9oSnQmFh0ioIwivPto8w
Sq3eH895c0qY1qaEPBkNTL0prPs+AH2q3Fx09q46YtZg1iOIVywS4GqHfu4PY76Q
3fdXBRgKNWqKVUX71HxpdssncdqjWVEZZ0NYHu4UDVN8apzjcXot9svBu0pakB9m
nMHAjUeI6zw1xKhiwzol1K/IUbvIOM1Fgc6+aeAdBnpTDVPLob1u0ETlJUiCUC9i
mMRFOz3uSLIORgHJOk7bejZE+4wfUmAFW+tTZFkxegwHW0wMmUtKIsPS0Izrdcwy
RfnOH7bzuR1xTMyp3TIBVIgt1N7DR6ytgE9o5zD7abaS37FMfRX5uYJqTGS3fnTs
C+EWbUnsxne296x8VHlEJaC0dwTlRIK63zXejs9pJaSR6R2FnwRt3pjKZQ0CF9K2
f0Xwb5KCY4pSbSMSnY3NzOTGkY706Ne+PdCqzHG6HaLJmR/2rh0aNVxoQOdntllt
ZbBx1Wxk9ZLEaI6KZy2nSS6DXkRYt6ny2vy3p/EhpSETzLIa6Zwp4POIj+raQJh1
/72JcT3W9dD+iI9BAUz2yNc1+6WS2IKUPSTYkc22xDKvkbDg3MRp6PJQwFZtHAOH
b6yz7YSv8ZB3AFiWziabqMq51+5JXcHxhLVGhiaW8wuSKsDk5xIjOaQlCgcVJcTq
92KdL+Gza7qZwOveXUx3nt4fwefdfbObhBda+2bkGBRElV2QUYwI0jucmonbjWPG
woa/K7Nd5pjRv44HfjC+2z7JRJIZPxbKrsuCb/D/bcAYFe9qh6vYUm8Q7KMPKVnj
DyqUYKnfQdODBctHV/p3TJyUaR8VdVaUurOCNqTTOfMzc2Cp1nqKcIwnj8G6Cttj
VulvtZRiXuFITvutreLb2YYzf4mG+z7ocziwzIuNOyOapSFQcPtzJLVlhrLTXejb
SkUeBpaQ3yyHd1GSSNjbE94SBEj+KEUuVDp1IYpGWDXTwsFeyeFWz1VqWG2T3oXJ
jlbHK2a5oUmscd+CQSjDucr3fFhHi//kau6+SgZVSJncsX+KQZLlbhKjYeXd+sPw
lAbIc4c5b9xaMGzzgTYWrbr44KltJlznVGhVSfEV9nqYCeickG4OC9roZibw17we
4G5L5sqX/ugHihHJJ8KoA5bV6fwUk6eiz5b/AMdAMAxA1WpDbqjrJCY62NFZKRna
/QMKbBP05Nb/yZONfocx4avEssIJjEzRL7MrT47BoOjo1eivZeM9dDG0iOLkKYbG
BHI6FpOWnBD9S/MV1UJQVcRDEkDIJNhP1m3W7FiMZ1smeiKVveCD8kAGEzyDXPNP
K8qz+0BZm9rs1VpqZ3ySwvNIO9EX2zA+qnZaUo8c1tNp7meIn2pdP/j7JaHmtJE4
1OkVZJElTzfebjt/tUA+eqaxV1nmFjuGIwUVM/+A70SM+U+A+CL49tgYsdDBzU15
M8TWcsB9WHyTxYDt5Y1Kes9DgJirDUvpvdCEHRBEJnbAHjz/9Yo4S+vX+ZheTFHj
G1yH3Y9SwWb+X1W1VdXoO35IfmhuiLl6DQA8KuFAgX/edYvOeScBHVtEG82sw5fY
k2V/kCQTVMB8qqMxTnh7J0Z731FMtCdAZyzlrNzH1AKmSgRnXAREGQCjNggXWB7t
Dipr+a59Ppj9GF4qaa1+cNE7S4x6H/RJcUn6GJKKX0RtZMskwpwcVCqoZD2Ny9Os
Nnapgy9gngoR0oBMO3AGAAUCC3B2mX9tAjIYkMLxSMXSqWtJfgOGUoueahMrqolv
Y/4gTPn+WO4+XoTtgJgYTjpGXafFqrECm9UC/wMEve8OSd+3HeRtBJHQcFwusUww
6JxuozSQzlCAieuMv0jX2CBMGNqhwIsDlVKj0WOnbTUJr3YqZmVOeervUJE7kkwW
iQOWP8SwE3DRhEGsN5efJbD/X+nN5dDixnjsiYZD9txHoJHbvfaLwHS/6n2tsQyb
6EKW27w3a6E/5c6UDmXxZhAFQ8TFooA5lvyYY6Z3phjtDQ9jamMqbKYNRMg+aR7y
fSUeBCo59JqQw6SZbpGlMC1Xt4aOThbtGs5hkqXUhQ/1Zsl998c0WDs8l728MezI
X8jAB4CKGd1DfmuKH/OwzF3gwMphNS8/I4naHJMJMCEmJw9W0DIQSlsXPMGhi/si
OpbtARtdg2grLcSwXYUm/IqYMXNCmXyhFXSVpQXf1JfeUQj81SmgOXby2yLUNnkp
9WpoZOOmkzeXCWOowEMSqvE3ipotFVG7Jq+o39O8az0IT7bsKlJrE6SnjnQ+Sm4Y
w7iFgUlUp0d1e+q82nuATlEFTA5ZBrEUZ7pORIRl4QPte/J4XVAS3KitaSnuYwDQ
KRxZk1h8OCLxcvpC1TxILHUVzg/CoXiihowkpEXSj5vvoHYioZpfYPSuVBclMLkg
wreIfP5dK3G1tNCWitrq4bkCCLbI1owVsspoqd9yhpfDEuKv3oZ26MaIqydHtRgR
7hwjbXpgltEoLmW6rkYUxwWquVIXFnQGSv7wZDyb30e8mLMAO3JNVPrbVkuPl4Pg
1gvyD+qSpaziXBX1x9mdMKszXcjWxSNfrxBR9jHBh5Z8a0znX3RuchDVtgDnjXi+
cBOG88fFGEFndkT9+8pMS9bjSi7SUtiCUnXYCi9iIViwogGTM4lZCxDKtDpQ4ZBw
eY0b1+Q00+kYmQ50c2BPvkL29rv3iac2tartZfn8rp/nt2DCeXiyJRGGidOGjlzi
y687k/wzRrrIHMTKipTzN3ZJGIrdTrg6k+4LFWV7+HUG0x9h+3DjdG5LX9D04Nnf
OtTBlwEzlPBBaFfIvatLvixYES8uZos0rlBX0oMto0QnFjy3fRDSLwStKdjyeIxC
abZVpDBETT0DsztRTN7F0qOB20O7TkKA4gAf/i7l2z89q1kOrgxRta7PSFzLzb5c
8i/PAJZFkKmBaTZHC3aI5COUEpDJDAwL+RfBRfgiROAEjGOYdlzJ/iADX+k1D8yC
O61/clxsBkdgAsheXUN/JHiOjzGvm1oiM/5BOTe9HyVmmymouIsIsZuIjydu89xd
OuTKPv7evOgY5dJExWuwBnbZ7L5VUkMRw84ZZ3R/FDv7LpGdPysaFlIyhY0slbjq
wD4c98sZsIVn6xCXp6eJJ5CDi1kCCkjy/taaZ6B6vYCZ1E5r6IrYlmTcPfgFYGpN
C/AFReoVfvZqvrb4tUp7NU/YZh29si/XssVUPBIJwp37K1gHiTOtQdEdH9kfNiA/
ooWZnqbUPCK43Z0jBL+78eDWozdTuLi306dnM3uTIi5oTtBnXa8YzVYalUKGoNUA
54W3VnGnIi3vK41k8ialcArDF86vQxv5GfGut/ZpiEMiPY4Uav9evUbllQYz+mQ7
k0HWP6d3/WZT5yskaGoyBT/6y0LomGV1C6eabWgDm649uYFWjPZZBDUPt6FOUKLN
9JZrT6Wr3YGag+4y5uItCQwKJG1mHETidtBSAT43WlRkaKSuGSTxHdGv22qIs122
gwra4zpOio1IqpP30lPva33JeVPkjl8bK9hLy8UA7t1L1EdtPnz2O28UOEowtEIc
9ERVBJlbjp79PrB1iVLKRUPZdXBvpLC4FS/fryEDftfFBritCYbb2SHzRBTO2quN
xul3bJyM4QWKE1RE9cNzZgZasBldsmLErLQ5ndyoYdnXhIqKZwbJP/dg1aPoHfFg
drMbmGA7kUouGECSddEkI6c5Dy2/UQ/kPDArcnC6Yy54BmObqlWdMAOTYGWK/Tul
8je9lvR1wCT/T29DpTAb+1t6u4u5qvhsRD+WN66SfmpC4T+P3NX8snRHVg2KxKbf
4jqSUSMP23hTYT5ibtCmEcw+sOu1vOs5E3tEXlTvnBh88bXFTCT0tJfus245/KX3
wHr7ufDfcrI/DmYz9ZHtz4Gya33WLCwBPbb5NpO3WfrmwfDpZ+8KT7I784VIXrhk
cWH2OfVoU7R185foNtF9yGOjWKCkGNCjprpr5eq7i0Uh7nFO/aa76S+AU+Nyryr6
7sNMxI77sw40AAtomHl/G5Dnx83kTmqdmdeR7TZMZPdYTAt3o3F9b+7WIJck5qPE
tOC8DbfN3/TPfJWWYRJYhJVbnDQwxMitGBZsAlu72x7ipE+rAF9xqRu2KBzNbHEg
3z6in8B2juTiUGCRSoi1ecr+vnpoMH15fxY/0tYmHxFXCNbcDssLBq83hYux32A0
i5mVHlvDOcJbeS2AjvlygayYpsAqZ1jgDa5QsSj/zVWjA23XximJyPZpyIjTk9Rb
XIf7CaY7soqN0U9w9CnThi3OLQxFH+HBs708siCI+D4+o2ayo9hBEqmhKrijj2Cp
hvusgekSEj0twflO8SKGg17Z0Cqm3dROMHao3Dh6px4Jfg3oDwu+ByB59creeliJ
LwIf8pwBgVG/RP6yIzkUSsHnYEWrwwad/A3AOZe+vGrv4e+syBoYqy0LbH1L6ica
QBBhnVTn4iXxHfujjo8oz5H4uyPyuOIJMwunA64tFI+ComGsCwboGb/EAqQnoBYY
x22yIw1/06yUkXVetzUezjnIP0tvNIpXZw/3rdrivW0rK2bj5N8QMvgmI9ScTTtb
cZ8sepUWnsz+KNRDpveJv+WK8epucxcUa+TD9w7GGrUogyJ/zRBEhYch+h16Onxo
ZBKf9GEh+ukSLweUIsY9Ji0fqOUhEp4Q39Yjx1z0eAVUenFEzaPzlySS6gZ+4akN
otE5jJCXEzQ72X0wqgQ+uBYrgww2HAXLLHiqeUBuamI3Ij3fI6SIf3diulzRtxgS
sg1up4/VqxwDoQ8pQO0XfVd0DbL0ST9d2dLgbW23tB3Xg/Ln6V1gAFOINeUPBe1d
LKoSlks+CU3ptlrMSQZfBl/aFJ8CLDOaohwVqAha/5FmCht/BSnY7zebVH1jEFk6
wLB5dJhmnkePAkLb8bXdWvXdULeXTg+Xa++Y/p8f89Qpz5h2V74Vyc0ykKQIXDpM
MWat/zmB7o7lVOCn3LJ08XTau66EK/2c/LdxeE7Che/6iK1DCdA9Y36CRb4qRhq6
Ivhe1uVI3BrsxxW2vks3qTgKUVRVoWp8Y9Zv4g2c1eaJecsgqqvdUfQLaVwMO2oo
cyLtRd5Cag+nplAEde+BaJXJfr8OsuWBfNSFuYjiBhZmkr3eaUg1/d2IY4OyeHnd
S0DpeFFGNeVuo/pOU+KxX7D5XBDG8fLIOaNJoKa9FluxkTGTK0CqkaIsdpe4DQX4
O1PT1IXXr4bq55PzMQiUe7Sq8FbMJSPBSIjEMJ5mbDaNjl6EASqE2pT9ZgNgtLyQ
XxMIy4FStY046odZYenkXbd6sJ+welRLHpI+gslkkg8YDsSzU4DTvslY/nsx2WVw
vByoFOTvMMFVZd8xIIX//LFxxfJIs7j/GcLRIMetdD6hwRphqdHSlcMNqev2U6NI
u4sv6GZhTjJMT+q4JfszgLc/rrmsrAu+o+51kxXBm52476Cv40Ql6m0hK11hHMn/
ElPycpNPY9zbfCHfUyJaipvHDb+m9g2awFVs4Vo7xlf2yhPoAD5VdRNeSH2b62b8
mbYR4YUBqML2ARajJcKK8LEElPlopVznJHmAtrkFXYbywjDBMs/zOla5WBRTm35A
wD4Fr6P1ZMYsJamLP8WUI6qk+t2K7hiM7l9mUtPpIixAecxAtYkZZAVhBlQ7ay2i
6PtbHeCdy4cCKirVWskMVx+quSWvlACnHVgPYwf71oYNx0iInt2nOytNkozXgB9/
LZF35IWUtSYWYPJADj5U7292Wxy+drvzVsbE3HNHI3t747uLuSQX4gobXuJ3vrxZ
sPAJCZ1+Tr4Am3Y7pSSu9VXfAMYXm/V4u0AzP8uJZxW5mTmLLEJkVh2PH5hTqrMc
qZETGuu1kAzzgHG9va7cVmfiHbGft1OCqUSMvXTjHxOMn88CDVPvH8SlpBhbOYnO
T1qkcS8kml+GKbZ6u/fNx/L6Yylmr1chQay4l0i63KDtbjgb7kepQW65plsg9jJn
4rpxPb2TNTmEWD1e3Uqb7PQvL74NE0Hx7+IPl6zMHzhaf5Q1YU6pXN0ild3SkV0O
E4wcELS2n2AxWORLRNTF2d39ZEhsywQtph9m0G6F7WOUl1F4WPahcd8bQ/EVLG63
1o2whX1mCZdybQOFUH8adewn1Q03Qy7/8bYU4Dgs/Uu8OBQz+MVGCV7Hfm6ezCw+
SOVXyXXyNFtOvgBMJ0hmhWOV3txphxKu6v6zasrQpALAnLDRQI2fD+LKcE+Gai/7
QEnlyeegZ0f2EzUwxtBBm05iEImtQinO63ghkb+ecH0KuEtefZfTbNy24wbzx4OI
Zh4bWC3QMgc6dVkWSK9ZqcVLEW9H6cnRCONsVQhJf3iCIeqzueiOJemYnLq2M2jh
SSoedb8+JyhD2Xj5gvtpjObJDaxshtIDftrMpm5nZFGSUvvKDc/RrGHEubWmB5eF
Swd3XwqJ9luLDVqkw6laljEEwLPZK21hzpuFFf3+SF8o0djLkskiGbvQAxgUIOrI
QJG5ziPzVlaipqXIJt4yxdiJZDcll4BUrUQIHFcpQxzWAerkRfsvoeCW/JRJ24JU
yG94AeTmfQtp72BHHp5AfBMLmCOCaJ4rBK8drWEvuRWK8mkuAEx7gO6eHciObB0m
No2fDLgr7FXXlkBqeEo+EJEAQyhkdiMW/w2hgryffUM21rRDUPJRku6IX7Nxybg/
TXA9Aa9ocxUQuwf2PnRXj1oLGRO0Nze8iQ9nVFkOxmZla6Rh3m/z9MCEgSTlHRvO
4LkhBV3+zSUNG7M5NNgCQCthk6BO256ajA9bReMql7hsCyfwFtPRYwEZIUn2fQx+
cKYhA+6LgXxgmuGGk3G+vfNBKpkm3mTyur3VdgNMNUypXAzKhDFl08PZAewOWZgd
UqBfzewgfXcS5ya/IkA5+UjTc7R9P/W5sbByPKGd3wK6NLE1cYTmDKYQapSm9b2r
tX7dqOnpkqPwv3O3kQRugleUsrT/9iq8fEjd4MotIqR8923Ttj2bdBqKlQRqPYP0
i6+m1JOZHZmQHalTN1xrEjRCcZEkGoT5tLKMfZSqAhP9M9sxzbAVWX2GcMeZ22bS
v/jvoI04dk489ZSa4/C3h/YnEYfnTp+GAv1qiJbIYnGcGzs2+Q544VACQ025Gmkb
BNokJx9eP9005RhgGAW3xUcz/8SJcEhpy6/wTi2Rl3f/6CHT8wQbxUSHOWMYUzRe
yReJ9FW9xMCg4pFG9VPWYbrsDFKxjF425ZS35824j8wZgVFjNyK4ckA6vCVo76Gp
e4D2F/gNMwY2edE08JY9ajIxLaQrMH9wlEaa8TOdKRmThcOYIu6SkoZfOQ1pMAY5
QaVknpTIB9VMsWOVYOKmICzSF26W7WjzYc2OSDXkgOaSZTC6i+kDfRWZ6H57KZD+
emGlCTtvuhxGsFJ23xpjL6L8Cx28eLmJzKzoxKqiiGWJOy4YanpTFRBQqH/Fzx0R
m+sASbVuKpt6L1RDhb731Hw2mjXZAO04bVVQ6SlhHq8+Fkl+Vul1ZCh5WbWcZskS
JIrzgzQp+aNC2lxCOFjklkQMQmLIKk7gOHgfQ+TkpbwHdoxT3wTvBJEb9JGgKLSn
0ENgZCqrC2T4naLicXSTwWsaMkB6QlAJy6esiyULR6oFcyp6X/xDQpWAlFzwLcFD
iEZJYqOeYxilLadgBDK4VJJksdhFG1mhjx7oJ9PeCAfDraDGz4Wvyk0uhs5TlNGJ
Igz+KqktAwOrnpw3ht31RiTHvb4jAT8Hr12bXc5RxqTNHtgS8v5FaI53zu5kbuYy
AZVDJpPifzaxrjLsIQ4pIOZbcKkb19sDIC8fk31Hho+FKNrmPcsTnYLlSI2fVKCS
R/CpllAP4m9wGWsSJHpQFPVZ0xKi6O18jZpkmk5jj68+A8bG/54wMJfYMh5fMIPf
mUp32QZ3UHdbPo1tfqg8WyY2BR2rBor9uD69Yd6zygUcws1sq/KIJaMMX+wbTzEt
VXuzYlOZFnFnaGo5eSFcnMWMicn84TBDJumToZlATmfxu94YycbhZfEyJ99VULDc
NYriI1nCjwKl4DNFdE35EBRjnTd6WjK76U+iJmXmmwTwObaFNtBjb7Mlq796i2ou
Zxrr7bVVcyHXyTyw/b12VyEq6fQAC1ZThhXb8wZzVjWvaONnYacM7L4aVSm0hAM7
MBh6dSJ4fz8eNfn4ReoGhXDNOK6N7pEuD4lhHiuNhFW/jOOnwSV00AHi2kZd4yVj
VDCpGOZpNLX+OTkLt9YXzdNHXDj0NDvlugGeBCBg8BvaXz2WYlFOv3+an9fsbADj
PHXSCsXTEjNVo5wF5rdg00JUsEAaYN2nqz8+Fe+YJPShvwnJFENR52y52dPq8Sc6
UrAwwPhkenWT2mVP1RY14UzHIzBoJ5VG8zZwz88vjiPtrCT2ssQQYVu/mhjeK7s0
B3Yd6tLIUGPyM/ZHYUhu3mZQde3hQDp9GbM6/pU6srb8XtI3JQj4ab3DZflEUL04
uFGDooxgx2ZQjSui6D0nWGsUeJq6L2UUHEkPiEuUfjG6B1vQg9pHe5CK4pgwQoGB
1gaxT5dTAoGOmQX/5jw6ZqZfH9kFO+2dMdJ334SXwqQwETOT5HDOvqNOwiB9x5Rx
Rz0BX88BrqfEBatVREkHJtUdXICFVTLc6AwONFiONpsD9oXz0WflVthe6JUn/83F
6XZ3cmIRkO1PGF65X1GCeovJRe563Ni66+UDp22nKERgbO9I9IMQNdA3tdPWoY/Z
WCDL4mt8GKFNlMEiR931y8LntubEk6jIOFsUyaC7j3TcaQ4yUmNb5ZZEWiRpEtjv
aCtwjNo+NxffkGXRYei7SLoiK1W8z/fMUBs+3WE8W8G/lPnzGp4O53wz616Z90GA
RGlsVrPFoDFOjl9HCCXevDVW+Bca1lZUYPeBeTsY95EhZx8sGd7GhqBpmqjTduD0
yogrufmVZkvEFvnZmmjqYXslJ497wX1Fq/e1qiwGaPTLevIcviz+7ILclM5tVTbG
nvDBN6ll76WD/r1cl/v4pKBqwYq+zs0HqQFMnsXygpv+JvF84ddlNR8qjeIgOjDh
MM4ucqwicJ8FMdj3GRPSn04A9Ill2zymIRtrE2yY4gTAtYqiaMpbU4BUY/EijNaP
02Z6zdRHcoI8VjbqIIsxmyEyPmcjBR9yExpzP+cNJLBsvLbKbMZdPpscoG7HNSC5
6Phb3z06gItcQl0LOMpa3KMttKcwFPXWTiRqguHN6oadQdMFAqN7J0+nDcBL7A8I
035uphy7JbBUJQ1UBeXXBDxbBuFneWsG+qujGT/3JfY3p3hUISyNY5y6bxDYi8t6
Y0WeVCBDfe8NfbxWeGt5YUoUDNd0URwZVWu7G1wUpENYHck0WNhUNqSjc5oHyoAq
I2GscBb1SoRvo0PVXlW9s61aCb+3opwbFibs4F34O4zCy8pkUUsihEvTdX5Bk7k5
18uWlApP2qfYTIQbF2TJfylOD7SyhzAYuZgmFJIjXVnDE7MpPkofM8r/OeLNzWB2
KRo1m2jH7aG0XsLHawVgD1SrfzKtkRXZ67bnUi1e0S9AUfjs/h3zPtrcC9maUbpD
GB+UqV+d8nFxLnE4zog7HHDwzfHDaYqrsW/fkqtRaiQvZDR2DJ3SR8ouiRfg1cWN
b2cZKtlx+c6YZEbdCTh1jvVzXrvTZIqYEuLGh1dnMRsRg2v8D9xeMA2PlXziXB1Y
QqEuSwielTYv6MA/xur7Vlk/b1/KRVYv9sOddy/Pwuj+QjV7GyWoXWExp7g05mOI
50VBFPztcn6IUnFfyFN9Q/NxxqH3/Wv7b1UQ1FF0MLUEyXC27CjKLnuk3ypjvN8r
BNXmLct0VJUB9lOp6WfwNEhv+bkXtrFgfUIkSqtBmaFPRLAjvsAk49PcsIvGpbrf
uDBdOuZjuG+WSrq6pujMoxMm1oeyQaU+TK4vh7xRoBS+eNTYFVNxo31NNT1RKfEn
MEAUBcBMCnhFpE7S/OhyDoOsePdALmKsEFIqNIo7LmnVCISSkmzVYeUA7p9BJyRQ
RbiHZXSu0j9RO5Dks/riNMV1Q5kiZeV5Xxn8Mw5M1NS8+5nuXVvbzsv3lfP8TqD5
sYP5rDEKTdge6RillOWw0l0mtUE+HYZzjek+fjQVGSayWK3QreB92BaCVp4gQQH7
HatT8Iavsmzj3HFGhVBwxO6TcBOe8OnifVC4830yWpgpLDK50gouxpfQMTb48sNV
cB2jt4+o5RCP0ffpYUJn66JOrHdWSqhRdHA+BQFVN7jo5oSOhROL4dUn4p+790BL
zNj8y1iHgOVUKFP0hRgIU4bsl4JMZ4l+jzPHuARxi6vXLInYOc/XssBKnA4gX9HE
X/9ZFgNxdQHLFBtfKEaTMZHkwpnuMs6JsllZGwHYrNw6BTbhbczqtgL0fLPtZ5FX
zgAPtZTiRixwDsJCwwPSlRou6Q3D0iHMOBfvVrZ/XEvdpgqkGDnL6brdFZlvfreg
MYtd98gz9gaTzYvNIDokuBqmmgtaYOL2jSWvvENQZD1+lXHhXG5zbx3+HIWu61jq
twVQtR00MvKejFbYuszi2hMMRLmzui1IziyBLLM6L56wF6m4Ide/u/DY4GNRsrou
XCIOKSJMMeShsZcuQlTs4LNBw67TI6iUx/2+9UMKNjj9zKJrAcxjA/q8yjElBW7P
OFfhP8GKGd9XFGx9qLyU3RWjO9S92X7yt9EWsfLYhIGXGo7PuRdItAeSc0fFSQ7F
6Cl2UkA0pYQ+h4WS/1PhDDL9K+QeunVxg3FC5hICh6/nEjJFcyZScE+gz1f/B/tQ
IKeCELakYDYktCBTxJHCVvu5gCbfmurb/hjPFfVkdpo1ico3aoOPMWIVC+yfrTTF
QE8LRORFMbhWibAR+DIsptgmbOuIMsWVy0kq6SKoClh6YcBdtK49eEiNn3cLuVDJ
gAhC/+Ym0qf9KOMeIKfyIn1VW5Mk6Zh84SxmpCFMLglsX0VUIKCv12z3cC8qzzhE
r93jC2bfYgoiDOMn07wUdI5jSy91g7jhM7QaGCTclhjUQvhxp8SKVgmThwXpmSFo
P/5ldXFE+/5ZjbniMGZwtRQteISkjq6+3VedGh6WYFy4ETNSQwS15G9WpRz9FK6L
kgS4qH/1rIgMC7s+yLFCn0GlGtctwWrrlTuZ9WffBTnDSNauZVxJpeBQNxoQPAED
xgwMBZD4X2ZNSI7U6s4VC6jXPYXbrPJex4yPy+u9eqNack54PpwefCFjsVpO0dMl
pc2NfO3DnbILpL3LrwcjqWcuXhh0elZAOVIjZ/mhebZYT9mZTXFWgtT0spQ4h7fM
ldYQbfdl+AHQnQTVGcsq9dCiZmxupDtCXuqREfbo6Vx3tCBe+fGgnTJecXLzmVod
If3OMWKT5Nu/B1obpCFeX/G9YYvr3bS8pzkN6V/Wcui00a3NH78dXP45bTnkUsRp
bhDhRq9OQaP/yVNf/tw8NC+71mCLeL02IUJG0Rc85RjrTmbuYchXoHFNOYH1u8FN
8psuV7NejsYvSciyMgEmLEAK09cHfgIH/t1895I6jGItyA7tiyBhXriZSJB6Zggn
orwxCCLFSIxEbWLpaMCMPomEAnU9MEjoseZSgXj+2C2i15j1sjldY7w/OyKjf6ST
4SLHPj53He95UcAhnxOUTIPDxZhJLcph+j0b0oTcGWYcvkLHqapxygA+j7hq5kFw
2LhUYi/yx4/qL+z05YFpGOixZP8tceKZqZfAby8EhxWNFu5Y/y6gRbJMF2yATeay
nLl0fEmXUEiX7nSDhiNKgJnJQ0A+IQXYw6UrhICQlkHAR45bV+yPokSNqotJcIcQ
umkw0PxdTVIX8+v8fk6vqBGW3zdqKC2GFBN1CdWCOqUWYHKoW4Z12PnqdCeOxMMY
wo3mCPba1LXWhIbMo+MTQUBawRfjykFK4uCPJ/RvFZBWCwPtRcWbKT7E2GJrvzqe
Xuxycq0WW3XxKCEpvQiypdyIXbZRJCzKlkfIOhKD6dQ7HhVMMdmHesarSXb7eyNz
gsNAaSvV28MRvFxmDFQ/0Xqa/FumngAOiwWiAvCihEAeJhi6OIVDJ1RqxvB55hfT
LTr0+BqhQmW1Nxl2Qb1m2QAqT4AdeCIFLxmSlOdnsUWo745s7Dp1nDTpN2O2v5yc
1svlAJWyho9yXvUa/8TPe0kEZLv5h9x7wbUAH4obIXmNWpjKxtfwW+tYDhXKI8hg
i/5Vpcscr6ZyNKPhMzKhKUmMDqzAPA4dLuqRXELlWuNehECpn4KWAP/fdFBeT3Pu
IA1YVs76e8PerO+fxSY0sVwgU+EYVdPiBUvQ1++A7A732LdcArgnzYS94hRJvyoc
ns+CHXlrsVt/q7O+bzkxHHsaKTnVdJqJAUwBd5dOv0JW5HAWwRPJz9u/IK32In5t
z9pP+knijjFrRdQHf/aNZyElT/PjvyUJx/UWLnbrsKZJRvZERI6Oyox5xzSb6YYE
4Tjz2BZLfDaUINt2wdvGruG9ZnkkeVlFsZ/9+bHvrBHylDvMeZMyYXGTbYVbfZnu
71aqhuYF+R9W0ZXYUm4Ka04w86KIaf/VS+x3k/ayjyhb5seG0q7IefhQerineUB2
b57/G8f+CDAlLq0e/rDa//e58BKsRsJQ0WdYSJCZodkUNfhXb/AOKMC7k3SI4D8s
AkOWB0LbC+668CHa1x7YgPDgYI35mW0CsaXjPintvJmoM0HrKqmRoZvrxt/LSCmS
zhGOB3WUWAkvV2RKzjY1CX2TP6bRBwvU1UAwbpUeF0AmcYoVWFtTY/D4EUlbZG4u
0MBg+s7zUbAJT6nE+KrVMlZme56q/vM2/lI2vJAGFxPZvE6TmL9Ct3gS923tLGGM
aZni7BsXItTN93QyArRErQuupJgUlX6dWWa5YhQa6M5vpL+3Tw8sqJE6E01bVpO+
TvcFcEI8V1na8qYz9kgOsTDz3ygRIm0GczzWHnah/fGS+SgUwhRc99J2gfv/ReGZ
M91THGAQ4a7YuFoB0IBFg3t81zkF7GPTNg0NPb8jY/rf/adAOVnxo7Pr4r80OVfa
E7FrkNZICUQ//bP5MhrVZjtYyNieTWQgx6Ct45314TqPSfLwkpI3vH5c1g7jX5xZ
BhDBg/nnkRnkbVYEv4Kwnn2YqpEeMxKGSk6EWoixnKCXWOrr2FExqPkq7EblxVDA
MzutWPVLwKk2lRCEx039sTwbzQC6I7dn+fMJQsY7m6g/Qlhi9LE4bG1q+0kxsxCj
VWV82rkKWlb4i5b7UmCSIuFV78Iphg0Zv+Et6t8sDv+RmeEMVoGloj9h7U0I6LJX
7oY3rhG0+DkpGbaXbeTTFXasZkmYsn1a3RrUZt3DEjL+OpGmtNvR3hqULsNasZRL
61+P3cccvlGPQy9BIhQrd+fjj7EsQ5qGC4O8ZNeYQ5/S9zBAMvlxn2lzjdmwSYpQ
BWmPEuwNFqqyrs1LgjWp056/YEWuYSVah+ZrhLHSu1flMdcXqVJ6P2NNZcmpT57U
2Bdr8AhLpz0pnKDTz5gV7MW43Yg+56jKtA3RIvrtvBVj1lEuW1X3aCm3QGwt7B8B
CQ4iOIlU3aGaloWDUnposnRni3XxFWOfMccrJrbwv0CrPv+Njm/oQ3abI/kOmNF/
auhGlUse9onA1Bfx5LunZ0T1j97nFdj58QXPt46qzFyCB0GHg0r7K9g8nlq4AVhh
504GQG3VdJ7OEVehaeqCWSIMd22+Q0F0jg2ffJQ0YQ2cKEU55SGbLpbfVpCcMUxd
obkqhPDKNLnY4m/uJVTcQKobSBE6438bW0Zk/nbacQmVhfVrhyuSvAujL9Vp4m+q
1v26EiLs3FTvuWWdkbJLUHaM+I05vWMen0BlgiYYEgJl8wF2EONw3Fe0Y5yTzEF5
wk56ti35pgISveeBzm9XczJSO8v7ZGvJjngPyxVz6kQGFU15gCFtriXIKZyTXshh
OQ6pmuFYP1B5q+HwEpDPwvJHliud9hkUIFTAqgHMIpHvOSLOKjeBe/tPQWh0864e
2h6UiNXzQGJll1+FoO5rGGu7NSiVRSM8Hg5aWZpztnBIXcZUOPSahGrAh8tBexti
nZ/FiXTy8HZ507GJKZ75h976m4SIEBSijd2eAGZHQ9Qr7Os7Hx9JS3ZQ8wwJr7UQ
XUr2IlM0A4wbYbjz+iHuHQq3m9aPg3tVc3bFYEqWroLL/GZ690XWe0ScX0sC6xdC
IvSBHnSk53lERQoV+Ix4l7iY6RaesS0tCUJq1b/5xm/8gKMnhxv0qFgMiyhmpaxH
/6/9fqqgdVTXynfT0ia8zDRuBDMoZ9gOwXG3YWqTg+4wwDFG/r9UIi6Fq/I4SxFY
DiFm2Sn5H5J+pWzmUIm5SOee9Gf/wd0VE+RuUlEXGSUA5NrZ1vFYkdoxsJjrr6N7
zboTXnZ1qfNwTRfe1hXHHS6POahsEDWwBsgR3a+z8I17LBLOZI2Bg9ZDtVnkbo/7
neDoG59NLlbWDJhXinjyVSaZoIJ/HrKCktqrXnZYLEYVfva4tKHLXfZT18vUm6MJ
9GU0/aicehjgAdvHm1ztKMUx62zDmr0hS9z6RJ58QM+dC785fhwzCZUgA0NtI/EK
iRNfH/0MAP+mFBWmbqKu7+FGPfAJ/Pt4tohi/4zsZdgSHpQ3cY0/pfRjshhFkUlb
gRV1pYy5OxIeDkrPzw3wFy7gmzNSWnGbPMizJcVkpYDgxp2rOEeRO/uaZiZbz26w
RNJLHVKu9YdJ+3S1vISlykNovLqkG3ofhzxr/reeECBrChWkSrGSL7Q5kSm55JJL
UbD3oUzA9yJsrvyU9lWnThQebcj0LjqYOA53U3nc0tBbdV+qPu1aV5ccpAa6vGxI
cj1ETZq8nluYD1mAmswbssG4kQ1MgCnfpVxrDFWtQFfB6dEX2vqV+kki6oXIiMnL
Yg6oEzFm60JYhXU5IwSuTePoQwRoB3dOzjSjE/wDDFg3XSEI6hi3Gp3O3dfuD7dP
BopnaiMZkb6UxMrsUQwZHTpJi5/pNm/ryOjHvNK762sjAruwR4c84sAXSNnt/bSZ
zUcnNK2i+iaRMAHEBpnN7szs8eJ7CPNW8rI6jpC94rPccRSObN51g7/zbqPg801i
s7z+dwyTGAVuZpXABPwQ5GllxRS6TBE1pxNU2YMZ4PnJH9Vf48QKrmnodrfwTH9S
6rd3Z2MDI0PnuA3I0g/K284QzjHCyfH6zubNHzNhX962409OuwXLnxTJWYMSQvUG
ngdVl8j74aeMhpjAklubIJ70gsFrPWkuS7RJc3dcQzFDTnhRaVk9h8XA897PB+Ny
9ak79n73uuSuOjK5hdYYg4z6YgtHxSxL3SR/UdqgDKlwdQ17+jChTyvCL+2PSJLs
lAkL0CNAqdP+NokA7GXwziKR6JZcUpU1ytYVpQ7jpiu0hX4Cr7YMaUjYmJWkvW5j
ssrdrEBcQpeoB165gxca5T7G2CMhzdWwt1jKU/vZZbgyGiyZNlJl8BBgmwOYUfeL
l+2lyjQaWwgnBgu6NpRVq4Qwdu8xgt1GnauORFi9rxUng16/C+xGxohl9lq5nMXq
5lQhoPVao8HfwtNXE9QtwqrioubcD0u00bb+k6eqGeif3iVQQfWDuFpfTrlj3AXa
oAD2eqpLP5Jh5ajC9IisHxpOkzxAeURK/eFCSCkV4AX/pkLTJ0U3b3j5jZImFV2q
KhGFSVftpZrKAYse8uIb7YBje6mKRbVFgNhKOR6cLhcNt3e4XpUfz2zd3a3wsS7h
97EF2SDk16iOUp7K1XnY5SNQixJhZAetcaQw0xSAVBrMHaw4nR0H8aXvJMw7m3L7
i1LgKoXoQ+uBnyjZ/ojFJFhsHfnzPSuOPsGo1jP6MWOPYM/h0uAN6MItjk9K44GW
vuHYCYacQRYRjKZlgmwB9t4Ux1MTEQfd3/zHmV94Y7p8ZSv5pezLPh8GGkaOdWBr
/zLvyI2yIPePMphUglvwJCAjM06wc+fncl3W6ttG30IwpAQ/V/17Jn39xekR1fTG
YZq+crShW3p0R/7DlqSOtkU/CEDBRVfBMtk7VCsPistjR7mU9ufevyTrxns6BIYV
47K7jUMRiO6gDOtDM+bHkUuiOlZPQmYlBKh2nKJ3EoI/nCua2nddLVEj3ANz6VlP
F6Dx0scHeG3einpcAUqNuJ6v0G6x4V8Pllvde5FqIl838VaWX0iuvND9UXo9XOvg
pG/eYU+zzWZI7ghN3ymqm1Z0MJQSF2NkEHoWrKnGv/t1O1ubDgHrjPdXHGI/AjOe
WmWZO7o9kIP9bbnP/J5uaAfhUXBZEqMBCY8k6/tzUs9okJW1GXhvGmwvy6+Q/bJV
VDpX7hducg2OzwinaVJk7qlXda5ZNQxmvCQ7KHHUDfNvTm0w5KBaaBbQ6Ory+Ejk
pq9EdlcYZUOwAS0eP/OIuuqZJ7bQPJKwucKxDFWPupTGjBrT+Rx1SF/Zs5RUWiO9
E8BPuNDBc+JmBoUVMv8an9u7HyWQ03t2Elr996e8ixvNh84wCtQ8vFbqOM1/2WF+
FItIP+D0aklBuQgXvYKz916v62bN0Y1dyQLuBwKT6s2D2xqgjX2HoCx2vVYIKzXa
BydEAd5HkIzLc7yPt0fhhLMcNsWAY2bRLrsQSjv3ca12WHj82o253e1D50HVgY/V
BR/bLdijKFZ9tAUoGPCIh3/cjWF6kC9WkBtIdy9ryBTGzeAMN13GOBg8Z52dhlXQ
vyahBLAL8iEVdopqX0h7i1X1P0YZVqpNupc0c6TYg5oc1mFfAKCVJJbJk6nE7sbF
p/MKbP5miKFgSHzytkjVNtYoLT+dwFOWyKc/7bIyh6iwyIm5NNTYSMbyI+Uq+GLi
SPG1irTZM3LchtCJMslXGgomPezgM82nD6ZJw53wc1AA6DASQSQZDScN2aJHvWgO
j6gJn4PNfpbUHvT0SoVwMcq6PVwzqkKhCe64yvG1e6c4mvlipHk5+To2OHVfSlMf
ehapd7vv/0ftOfnDkJqPRWdV3P6EAj64IUpy5kTAeqENv95hzFn4PyI5SgmCTIsD
rY+y6/KnT7XZdbxpsP9FU4fPLdlaackyrhxJvrKGbqkoUf35k2vzCEWbsdUWBmmu
+oAHb9BFTJ3XmAbLd49JEhWlxXul6oZGd2dGUIiM2hei+UmupDRbjviXjMW3S+Nf
MgxOemwVCC5pTlKgtldVygvIZ/xMIk6wRqD7AzUHBDzH7dbX20RSlUaWkUeMgLUF
Z5e+t5+sR2zzDVR4eJjozONFrkE2B7IRAXxyigMgZc4dGP8NuGjLoiD7FrROXCHc
B6hnVVP7bWlqNzbAz/WqmF1Hr68j+//p0FblgWDgfvLDcWXfHgpexTALvuXUhhd7
nFIevEouRJNHwcQ9o8sEA0X8lEbMaIsYVMoptTWXq2taVMBxowB6QS2eKrvErMS/
c1Fg2ts9/3LfaZqECV4NH4IOpYckyffkk1SgLEsf+iJcdLE4HldSmeTOW+UpGGeC
geQObO+kboazHnQMyFpOE3LqcW4rFzXHh6E2tHkzHy7XlXwtTVi7pSElBb/QLhyH
BLxm+NSJ9kP7DTOT9lbyH30AGrRWWo183fbhBvBUkq6Bb4nSBJisTo8ZL4QfjHe3
N3fHDQzWNTy/gjBJzWquYkPqR99uICxxQwhOQgMFyKjpMdI6Jy01S+ACNojmn5p3
cm4PGmeMsqy2aMmo+VE3XqL5qZgPJcw9v8RaVdFHs1NwKBBfy4rnG/qCHEPV09uR
q/4EmaffRRXlLFf7kSJwqOoyjsYYcqBhrYJFGOJ6LxNByvtyXARwKxKD2JgkjeGd
SiEWpm1JG1oMdaK0xA+yAGq9ZedTt7zf9v40V2x7xhKHfnwET2mJq9kFdaQz66sv
IiXoAvCAYXmK79lRNb0xKyt3+l5lZ8JbCdLNX68wuo0yVPRrAcDioQmKceEVzyYN
BBZZINhMTHeuQoJZULY2zG88jsei00D6O7KOdZmYZDIe7Q034Pbb3fd1Jk+CBIpq
h+gkzUaHaHR2GlUnKUWKw79QCCOYTXEAt/9jBbEVV51M86SBNNo9ALe4yTkWyB4x
dvBd7MybXz6xufaMj086KrTA19RbIvp7WmkDB/8ubQ2kSEjZucUFYmkJ/OJoHLmE
v7ei+fms520ExGdHvI5TYXASzFEBMvZn12pgS97IzsRduS2twj2yr8SKQ2G02gu/
/mqwFQ0q+GUnqKxH7OITLT/P5GzlvhFxJ/ttALzb93bLjPWjq+3OJNVxXj14QSwI
XaulxxF99hCd2IqW0BshwPQMCNrtBFZFJY+Yb9QYGfw4a2uxohYUSmSEKa5PwKrj
J5sbIldQbV2UMGiVMMjDTgW4zu3Sj4x8n/rUmIo+AjRryQY1a6BBEc5MGmTRq8j6
Ye3mwebrxDr4taTqZwNXvF7VnD0eAaH8CtPFoTU1dy6PWU1Xowbomd3tUvEWiASB
N7KfQA/ekiRSVopE7sSIGi6tSgbNx0XY1Ly+24BNEVIEEwgJJbU8oayL5dl9VYH8
wVZU0DcHvBIkG0J6q0U6l7xZ5Cmoq41DNUUiY3rFjeeiUQObVN7AoNWF9t3MsrUH
tNeoTVnHPts+qbGFVME6gtvrQjeVjk3qXjFDzAuebs1za7128T0hQMY9739eLQwl
VSy96maSQEZC1+ZsI2eGoRlUxsTGk8jAWB2IcDAmCaAGaCF9O1poH9jvLLuFJ5vT
E40dOlZBZIvQSRNYJ8Vvu1CrrcLo5DEJC2ZdG3FjFXFQiTe+uf5uRKpbNNv63A7E
e8xXmt8/NGJS3NN2xC+y5iHpnO5lUJ5N2qEwMFX7wPx265dR0OvCjndcvi2pFiQm
jNgkarF+FYX3fevIXaStPmZOfRd9hYZ6hEqeddvXd6UFU+MmSshaUWGLVLPzr15a
2CtEh9D32YYXSIr3Sokna0X6R763hJmm/c1RxNdqWwYlCx+aOPT+PMAcJ40Fm96W
DSFyupWnDiCCQ3BcXVJbViqbkJGsE3SZk+K1IexOK5FOYiNTmeY0Xg9TfhozqfOs
Cyng8FZgNOgDee6dOyG8jrg9BJC5cvAx81Oc3qXcNlkVc9QxvaRJ9SoQ5rre01kB
SXaIdSXCFGsusktbAj1eJG22iJ9iWUAZED8trf0RtV5a4S4vS3ktIYuNADL8pLl+
HXqVCJ6zvLKJ7UCg9K2Z4n1Fh2Bqqf8z9qU1lVpcAFzh9n57SN+5QMnMEG0aQYmc
PkWYFwstC4cP4fz4XK10nf6VvqpXQ4ktBg581ERv5jgF8NCRiA0j7vFDHwWCLrwm
j/QfGCLD/WXTW0Lw0fNoa+uqi0JbVwq4v8PXk4yoTtJL4IONimbqBLb/24M0K6WE
Epp3mQHfwAZT6wOrb4+GIEL+b4/a4Z9g7uGviv+IzvV4RcGUiCbkmVIDkwqTswkl
sAtaSqF1O6CL53jimIeWwcovlRbaH2RnodR/6igBqjTDY4Cq9Sg5ubY33xR4R/Su
+xVDSWphHrNMTHDrsY7qBAB+fs9bhRpJYFSpITpH8twqTaOEBRjj5ga6N4as0iMj
9HWYvY9Vegiwkw52TTmifECbYGWITCpC2LEaIP+mXR8LrfMCE7Iop+vax8r8v01l
Thij6liY5aqsbxxCLcR5NwTFqwc17y7qwoTXp7lxkErTEG60acl4l3ydFL46KdJB
wtudCjjRyWb+Qn6SqVKv6cWi40W4BsRubs0pNAK3U1vSjnTe7+iZZQc5Qfkw5RTQ
C4Xq2TDoEwElJhnFw3ktVb76Ma6HdCvEOIBXYA7PklnGZxLvGnJvrimvznkg00qB
6iuQokrkTfh7pPAfZKiRM6iH7QCA01Scfloz7l3vOOSzeOgyrLOE5kFL8tVqM0ZR
3FhTpPWAsHE5JLnqtZ9FzbF+Ielv2/7suHCylVWDdqTq5/Geg9hpD+JV9ndtLZ1O
sDFJt7GYnJ3Ec+AbTdWgELVNlDAqXMVsH7+XHcWAIMMTv1jptYBig1ogYlyMi9mU
gSlNg1Cq19smSOSiGwTcxORaZ5QKZNbX14E9aVv0vVHoK6PaOoqN2UYA4InMVLKt
pdzDoMqeMGgVA6UVRaR3kbbDPMJrZ/IBeGqz3SrayMqXvCtk7ONrC2a0rfHqEIZ0
BZwJVFA+2ORlBhpXT/FHLjoKJCyGBfbXwKaTxSriRqJRkj7yLcqlzC6+iAc3PvbS
61smqCthRwmOBknnFcvFryQSNlMAzoIdHI/So7evtlps9INMrXir7QxAWrSzdt1j
iSY1+mejJglGSKtC1r203sF49oghMHv5lDwz/3YxL/o+hZFORKeJSQUKCBBnL7VT
QnJopYbSHvhQwpdOoF79XusmGHBL87B4DoMHPQYePoBnaTare7W9S1cTCYwmXWV+
gM08aWY4TW+ioCeoOWzPmUu2XULdis20yKJxCAXxxbSFumVn4EBasL4BhLonfsn0
s0RTObVUKNWuTMnZfE1quzbWHtMSl8OfOsENG5Ocdbzr47tP+jeIhNtYpbHazpo3
ptQx0pBqd5ZN/6zGPRXp6ovN2zt6Lm1I/0YLLqjL7O6VCPFePV1n111qoUV6Uy2G
sioDs5dJuovgSKFou6OcGbIW08wsRM2Y+l+f9piyG9poNYDMmiky/UQoodp0qWK8
Lcr2PCthaHKEIawiwFEWfD2S6uxLQMo9aAeMXLL2Wtv8n/OhnMTlQPmROALn86Gp
M7LOgPr4kvIFDUZJmtqAyxpHRuXD1mI6CDW+obkolKqy1+yl73gC9XMNE0lY+OXi
XLx/9+6eAQf1NoyjqI2ZmRBp5eIg0ruskLi+DBZ5kdccsBKvDPp9Sowh8lI76/NI
JHhYwglVJForEZODKezyqV43ChdJbsTxIOvzt+x9ixy6MmScbvpY+u8ihrg10kyN
wJsj8LSnBN3NJ/+IyWeqUn6dp047FS6OpanesoEsGj1v9xwJO2yLBP649Ht1uHx3
WotLQjYuGOovJ7Bt8RBQZ1d2HgLKA/VQCBibf6ui+G2ZbR8dmWTbKprh77y4/9VG
z0W0cxvPpa2HoLzew7uWaMYxp2oPNErd/4zGKx4zli8Z+E5+XbskY6gdi20TOvDx
RIK+wOjzoBrG/tPONeoPuKrTFunbFX7f/lWxh3DZVCV/vrkVeIPc2tJeUchpMwGI
8owxc9w8LZBuWH+gPeiMAk7F2AGM0q4xX8NYwwouetmPVthw77oAfpwcyLeKsqak
ODWlBy3fO+yhPCc6orjh3Y6riIx/mH0qA8bbE+bAoFhJ2Vuktbwsuuhyut7JH/nd
06Q0mFVJ4Fiv6IXbEaToSq+Nt21d410LlLhBwk7FnGHPlcp7szTC+47UJdd+l9R2
GBI0+VHf0R5HtDzLO2wBwKXISDFmgsvtCeSJgMkwrhA1aDMUwoBHNOAlM6Telh5B
pneehoJkFCM+4RtV1QO0Iyk6O/FhaGd5dUaMm7H0SZWEmX4lyAVUcp1yaV+9/fWu
arSUCJUY2yEk53z72TPt2XRf6WG1cKD/ktcuCKUHFvRHPA6KziRI3ybL+Nu3JTvf
tvyJdAFJwA2Gqpiwl5C1eoLzxBhRCB8A19kw1+VN0xUgYJmpUvOJusfj4UmDyRH/
OZ8jSqawuQPp+sHOakGGnC8PYRqSUIFybqE7bl5QVWLYNZhYEtJSf2W3I/Ps+vup
jC7ATrAVdMcASWVVgBGGUpU9XWdX5KerjWZuHqUqFM3P0Ftr6Jxe3pI/BPQb5MNe
0YiezCYT1ZQcLskA74SX+vgxt7Z31JjqOwsEkmIxdCum9WFwwTJA4ZH1nsvOUkCG
WyDxLRb8hOkERNUG8y51C3a3KkbU3a1fzijfbNEa8d7QGxU4ggjYzNH1vuSIRcDu
+o1Qh7gLFyaxGH8TueIXBqj1DiTXSNhoro0+X7/oSlKf4atgxaAz0iZ0VuQoYRMD
tPAwTH3/MEqyX0V+2xAIAd6fFgsCiTxLiiGZncfCyGpgjcT4oWAUQYXf3duX/GxF
h0mBgOUay+cgJMSAV8JzyoKqvbfI/Fxfjxl9D5KxZH+yjDKoSZ5YnWmJqrAZXBHZ
QwW/EQZyMHZ4z6E8Tbw1VwmnBJ+f8xHVd5wxTtfb+KU92Hz7CWu4iZd8lEEFgUTT
PJJ8/VstXb3Ggm2k99L3nGaF8y8WlOTQTvbDxEXheniSuvDWjIhs4vl3nz0y+s8H
QVSRifxSbxr3TsGQlsyM9KeHsyodmHQM3t8YybPlgW57zfKXRl1CLUYXXVgIo8cu
LoqnLZCzgmEgPWcJoXAOKFQxJBUDcJGUWju7R6Ck4vLwES56WCIGNy1irkB4XGiY
G//n2T7Cs+BJ7Sr7htHcthhklBN6YVi/x4CeZQxSRQG+TAIGMuPFLFD4qv4hhYRT
3rcPNV3QCFaUtdh0MsPOsbcCOTA+0QEIlEYVw0wYDPsmde5Ddu9nO5Jt3mLsEYW5
dNc8kTXXoL8mC4EKWT3VLMtbozopkDJboeKzGFLWABbVamEoVA2j9+qUaAdW8uFi
CLfbppy081MKG0nv06eSHZsmyM0MqbUJA13VnjQe6ltXnX2XuOLHSngTE2T04AQF
FLqCWvnwERWnKs9MFjU6guMllHTuLHCZrevVpZln2/3amxdIt60m5e8CkUl9cWDn
NBsQ1YK66zq2cxJm5tMElrG5+hB7MwpuCSOLQezg511SewaoMcXO9JY70V+YdwDR
wJwAvNGywsZFXIensrrXd+LRvDBbMi+wkF1egCo07e75p7HI2xxrdjACu3efvAdt
5k3IM0yeE6wGeJnVtzEVIed14B2lzl6s89H4NptsZ7qrf6oqvqDsTh44kqvJHDwI
jMkNGTdN7T2bUNi86vqBHCY8uFw5B79AVheGtMghTvrARfBD7p4NY2+GttY7jtt7
S2uH/8jKfI4XAGIpKcHUXJh3j4EmDMhLpELAqag7tp2UqN0vALrtyMoTAh9Yu4qI
wYiFQ8wA4z9/zoMEZ/FY9FxO0pvUqwpnGhOPaYAyVLkyHs3vN81Dfuk6NIiQk2c+
40QUN0yGsHZxyEvJWI9FvrW0Z26lET6U3G986+GAfLnQsHrkyM00GJZa11BhYTJo
KSVSucWWDbrcg8jXhgtsiv5gGyOUzw9/K/A/+HOgQZOiThvv8Xkf29sgIeVKta7k
BfrsBqT5sD70zBaRPQvcxE+b1sOuP49iOg1jyYdZ1LCzDm7vaYem73goBub5wUYu
SHfcuz12v766VhfyAYR59LB2MH9X4TLxHCPQUbCVFugvReJCYsoKkHZtN+xWd/71
oN4O4IE74TGWVTZ1R2OWDVHzs5GoiQ7UVf42Gs+BE9f33E5YUxYTP/WD42dqn6Ic
bthH6dp4tAoDAKIqvgrZvtdOP3ovi8HyFbfU3CcqHSQ/B57ocsFPOsMwkYGWrNd1
uYVQEzDGbhEW8NvijUawp5bCwRbrIl/Qz/W/titbC75jT5UjDNA1vDOFh1hgNf/U
1Ql94wjqZ7YBj1pRC7Iwvt7aIkxCxStFxDCCrk3xVijeM5BwT//GvGPsfGWR3Oof
wq8MQ0EdgPd8vvmkTdudDNF8tvOQp8w82qVayYud8srots8Sat7Rrcuh06jPHvFL
YwR2g0p15bgC1bIzg7B3K/PExyh4Xk2slH1I6IpsiBEq3xzyIiYgLZjoNhUl7wss
Pp4EEv3uiAWsYVgJ8p99BnDp5RquMxQ4kFl5ioaLJhnldjonupJvNURoO2YBYVNJ
JBAt4uVuM8k4pvKh+QzlqEme+Atme5/Y4gr94ek1Fh4gBsBismxD6KlU1Rj8p2Mw
3CIwNNSDiXeRISTlFSGLuUGOQ5X196UyIV2VQYULBslk6PXxAVRDFMm1iLc1bVG+
9epCS7vTaej9VNiz2V8Dox3CK4euzeH3vGbKwNYJfDM+wTlFmgM0Ofg/yOYmPEyM
Ei9PRQ3ezYLjwSrHlhDty55TEPsAa/iGnnzWhYN35dy0J2QV67lf1ReRdJnAdwA8
MpTsPpbr0OMTI4qLwIvY4que2b8IQo9HL+splhREMdHiUzRSR1fc377F2WMX31RD
EJMOiJATTKTmHZSllcpcl5kAUTpgN9wyVy8+joEfkpTSfqfflDtviu/7OFC8mzO1
eK1saoCzIs9n5U0aTymZstvSIgRu+XYbNAzchVRCp3IqMMDpazZyYFdzn9y0QI84
M7kzKR3iLPrsSBBwQc7n6QcmyjS3aHrkfToZYnC0EE2HKRSnjLVJGmJoUMtcbSH7
xH++XTr5Zfp98nApf10WT57dWy5mevM6ktaCTfNlFTsJr+Ys6DrXwNkEWf2mbrsw
bVxgPYRx4pjeBP0058YPeSchHuRycX61+2QfqbQJkGjpta2W8ZsQMfFdOsD7IAzF
SDSEHzl//E8v7OZNz68XtAVnIM3S7uqaEHOeZ+CDlueh1+IbZQIgEWhbtILzYdix
sjEBKMAIZPikRDsbz9AgbIGqFn26BJESiyWENTHPSo78CU8Liu+d3pEr5qZ7N/zZ
rGohKeD5x2KQN+AvB0hS4x4H4fX3KpDLyHVWK7oR3hL0jZyWPnv+yyyBvwibaLgD
7X5WMAkD5bP3rH/oN0jgv6SDjWQPRZJRAOhsBFn0pwh5KndJdmb+dmMq0I9zA0MW
EBt9MMqFleB3UU38MLOQo6JJcGFVGfXx62EntbUa8W9n1redoTKekoGHs/ThA2tf
RO9FA6xBW+vaDauAPcP02pqYleR+VGB7OJTo5lNZSIHT90RNTB0QXvxWIrXw63NC
l/NbJKSu5v82hu05Hz+8jk4tamo4ahHgSaFwimJLzsammc6yGN1XNGOPg6a2iC9n
OYM5oSAO80xgYYbStxX0hyFvG4Lw7owNmsMPgDdGdaok5mgzxklZV09zc/U/waD2
ZaErYgkfixm04KWLMSb2ARu8dtueO6snFZU4fU+QUTqHbxcXQEnc7ppbmYEbJ1AP
qlCJeTuQmKSvYQghbkWN2/C/GYlH24SihgPXHiCRPiywYpUHWixmBNxq7lXtAYXg
ZHtUXWtMlKbGZt2LZz86ctNHTG1MPAHYyXdorvtdxgkEWkbibnGyk7PaHo9DEsx7
g9ZQLTvuqDLDLpAZIWYjq9B4HEqbMApGHTMtUFjC7UeEvZWBWD+VGpvrxD1ysNZl
WrZuqwbByAgM82SqWk+euIiHdXZwzKuZurai3hydOjAGGACW80tqaGgOqtq4RJME
tVA0lfSL9JGE/L0vNfZx0lEXCNKH6GEhDyGduOi7W+oi2dF1PtJ8sanY6VWJbRHN
NRnuU+VT01E807bgFl+a3adYp5FfYlW2FH15QIO8l0ex9W2gfcTo9A7swUwhOETe
LT40jnK+aRCMKSjHb/4OLP4229qVYvED8Z1TKjCXYdiNsDheoroXJfDjs+HNUivh
GP4FaV7VdPgc1aCcdq1MPjfVc1W2h8BG+tJKadowahy36ypAfFACVnk6G25ViZNn
Y2w6QTM5OWWeK2SgDvzlFJEvsizgNa1ftcUoskfZCLcUniPoEUKc9sSY0eME1RH3
6eq6NSX4LTVT2bh1Y2Nej6hn8bQ7pq+P5cnz2R/aSzno/w/lJp4rJ+N8CQiNOQT5
u5WB8WcNnknhjrVP4GxfV2sYiYy+2xOQcjhpgLbqHIQetxRhc3a/7Ilhk3S2QTkJ
Gy3XpZHGWwn+CntrFovVXPPX33SyMrUyUS9IneKmlmAElVRLJc8xBMPqVDwYBMwF
J67LzDD6OD+8sYd4Cn5f9zVxHFxUIJOUYrquCMQ8BvpqWfHo+0W96VInBS1DjndN
i/uMuwYj08vh3lUQCeNGpWce1jOil2zOPzMZwJw7UdaVGlwHEZjCMvaeeH1rrWgq
jEYokjtwxbQOHJ2zr4K8jzrMJSlPHViLm8385LzMj+hvqfcwhOb5+X1AqXagrTP2
Z246HF223RbCPYkSW3t+x6Smzq3ymSpADAHHHPcvF8ywsh/gmrTEV/awzt9ppv5F
fSqS5gQyewkmFoq3AiVF7NcKA0C4AcSLaCJawbPKXoW188x+LVg4IRFlE8U2lEST
h1DRaZWYgT8pnjImc9dpTjF2ufgqDFPT/EapkuQIL+vCG15ibDpTnLSV5qfFuFPN
0oI+XyA3ABEQ/akdtlYGVQhuOkn0uWexHNC/uR2u+QJj2zj1naT/IyoNYXrhnDlo
O2UZpTdnDjpkPdH30ETPsmRhs9onUXJrYShY6fjQzPZu+0h/aaPwINz/MNtkXLK/
BjyvbBWo+EcYQUj15pKj8pyNJL3ck6W5jCdiu1evOvhgDKtQWlpaWOXGbPyXfzfU
lhoTsLEdnrA3JOdxdXnQeOa4XioraLiayhe5kxldCA05At7M9uJWgOoYEHwCYbQN
ok1GJAe04/GfmJzjMWip+0Q0rCSgOxjIoBhC3D8vU/wXEiCvX8Jt8xsp9zzP8tNY
aiaQV4b2BHk/i3osgBKtNzgmd3z7idIsJ40MchC0NN4YFftSvJ9YVG6pmfmWlWY9
njbiU5Ypf6hqAA4opspiNBxrVpoQVod2+uHDqUla3XgbXw6ojx/VZUajmDwb2aqo
S2zPomOju0Pr24+pRBFjx5a0/MLLL+Bqy/+ZNULUHJDlyVZFvFP4qYyv0arrIBaf
cLcKDb1PoZrVt0z6+4a15suR5QTzwm7Q5DHM/jlYfTzPsihbJaE+rPIfYir8Ag8k
6/H1RWLbFa/+G3ZMFacZ360eGdRc1tFORYd4EQmNHr1MhO6atLo7X+oyrX94xRE8
8gyjqv2Dk0Z3Ld7LQk+fQOMLS7NIxTCr8+8U+omYzpBbZDTZh8ujaSZqkMR+RwDx
ow5Af48cLaurhlN9Rpsz6u0wRD278/2sDLzva2i9STjfU+grORW0NocIdXwfstNz
VpEzY6ZLI/TLOVRagF3bPDxCb+iclJXayXWbPnAWrOl3rck4uq0fNf/gPrQumnJo
w3QxIUiRNZvtMIgnL3gM7IfQI0N9Y+ar3spje79DJaUtnoC2C1DtuXBqfngll+I4
TooyE5lakKvX215If1xIfHBMsQnH9jXPFhGOPOeXOpj+UHiyqnBoumoOCJFCJPOg
BAH+Ve7SNoDP+IEvVOvmx6CCiK6SaqrNbRK0At4taHEioHZFJWP4BTmMd7NtJj7w
D7zpg+TRTCeZhStjmOIRJgzsjWDyWtC+k3TiQo5qyyS1ST7p9ubwe33ClD6KEum1
MRWFx7rV3/gtfCmnPrxwkMLCSujpzyfL3maozY/jVURslSxyWmzWScM8j5bV8OwP
dnAtP8rJTQh3h7MQ7lzhUV/MYH/99Z96ZGRtH6hHr2y4G3Hixry/E3D4hx/Q7WWO
mTehH25bABcvulBSmnwOX9QQpj8fpxEjWf0TOwlxBMrB5IxVdcsnHMSVDAsQ1NSi
r9VlLcr+bvEvpaxrNXLIz695FUKzG3Jn9HGb9gSSZrZLfNmcb5jdAITpSn4q0gDH
PtAWIBRUnwAQ6q/3NfFyTxuMXfRcmHnLnm5b5LJMDnhQx8jX2Gd1zwqmJ4MQ8B4E
OOJUhStF6rJmxvoQANA0MfjkOaQGSe1qKxSjPJ/+rhSMmonYb91VQxvN8TDI3l+g
pl0N0ZxKVHyQbvAG5GWfkjyuYvRC0BRq9kENNy1OP2K2sDUlo0twfh+091XGRbDR
5phRTbSTO2kgBRAcsFRVoZdXi0vcxgDcGAueGFmz/rxcGLy7hpXSF4SyUZqH0PJ8
oLCMpaO1IiHJoAqUeXkWgCJ3YXWcf2Hx+TLulJNW9Or++2EkDWW/EVR/Ub3k+bEt
bTh0prWX6UKD+y3av992D47iDdqM3h+hEWoJ/BPg9gm6NGNxMMLSE2/Q3t67yD8z
PPDaQp6nIVvWjQenSJ21++Oxz+dzUfYSr3qjovtMWCny8S1t3nAr6t9gTb+irTQb
y/HjCrT4EXKzx1Ib9EDcH9fshzzSipqTpUFY/jhtJZkmeL0i7izw00xYyn0wZYZv
D24ty/r2zLcihXqPefMlF1GyjFvwb4xBUhu9HQxmHpw5hM5I760HXNSTuHkAMIrL
5ATrohU3CH8AXDXSHGSwx8EM+nJymq4NPT9hgRnfTadUry7uCYzyHKi2P02IOGAV
l6i9QCKdJyIkvtFneAPoS9n8soztMjkH4LwrSWJs4sKq4M9QQFO9j/vS8SD/Md0f
RHX944KZoVos0Nja+jcsH87yIleqdf+ObUiXXv+5sXpv+tT6UMqZxktYrMXEECoC
P7FFQDQLSLieW+j0L8oOqZO6knkBZBhrw4wY42seFjJotC3glMCcoSdGHXC0kluJ
kTwrTeJ9WzySSvGVjSNdswrfOgZw5bVeKISvvXMXJHDmEGRAqTIpC/Flm/gSW9f+
ww1mK3QLi8skcjKVfhE2YaCEHmM1IgQiY6GYqZQKlom9p0/LUWt0o8NgXI0vxFXI
+nIkUMEKRDqMgLHiwRQ2GO8R5SfVTy2UKR00rrCWxRNaiJajaJs4U8YK2sP/PnRI
VS1Wj9MfkU01W/5XALIufoYi8fPcUZmxRVTt0xWzkKA0ReAF5Q+jarAl/7cb++aB
c6/ifk6+W81JqVlD+IksSZv4/kjcVEUyuMeRriGf4GyrnU/+tXXLJQFOlBcnhYlr
dNls2a/kY9Eisrsi2YYBI30hiS4ei10UNZVG91A6GsOondNiTH85Ybhb8XoIE2rz
cL/DwKGWcGauMiIkAAbxyVezouSwf09KidynlTnibJ/VBtOCspNY70L0UQWuSqYe
j5IJMwRUCZZvu2lgan2wyAOnhwijP9mhgaSPspLRWTQTpGZrbsplqg4uQP3HFLWd
xPpSp9ORt5p86tLxTVd/hcFOcyKL2Amrvqnn9Y2lRgQK1uBmyyVfo5tppr8vXpj9
rhG2CUrcD+pApxyjfAptExmGJTM6Ps3Mh0xVPRSMG0IgbKykXvXB7J30MGtercmv
MjpukgrGpH1QEmEby//IhKvM0npWVOVlCuiCNpz0ptxCYn2LHNPXtI7+U710Gd3O
ahPEZ5Ktrb0EoKu6eS9jT1EJViZ+AGKBv9ybSHVpRp1+27m9D/8bojscIwfBaPNT
f54PPv9YokuWS6/veGvNqTUAbY9tFHFyXqlSwaOLUVj/2j6R/BGzN0l9Xdw7PDta
g40mUsnNCcqDqtGrd8XzOFcJmIoe4W3hqC6DD3xK4TvyTugOwH7RMZnCOjHaeAVw
9/9U4UMOHZALl7paUoad7EWUKkiMoOS+IrZDJwwtxf2R2Kb1I2DAtSaMOcVmrtS3
7ddKmsa8QIOVi7h1bU7R7btxitPNew3Kzg6XGZv3vJELWiJlQCvp0Lp7bbk2Ayn4
hvNkJQL/+98u6QdSEQtf0ZAi/bJQ/z4HspAG7DRZti3YpF3Ni3hU9Y1ln3u8xe3d
tEIpjbF+SyZBxZjxrgJ8cgNRODxLrc77I/7TkYaVUwY7JPoCM/WZkD7OnqKK0AnT
soYB9NNRgvANF1g7XSsJEv53zUalF9xFl/qBuHQDoCqKdvueajRnUeZwFy0yri0+
eAZlAidloBuTOpODdfanK4Su/pt5hQJER+Lnrv6l4v0mIPKJ7pAgvsNgz+aFoN0m
F0C0l6DJxcgxXwz/pJe5A+eu1vyKOLikgmcbmkZ8gwEP4b4gv+2PRXhrFLmYFY4/
qwb1SOkDqEvWyKUziXEMHW2zXxbACQSqZUMwz3ih5RHVqwQB9MquAQIRjuMqoZpN
HABUBV0x+/OmGRQBBEVjfk+7q1e/qqfucouAtMYqgVTBTOYNblT4KS0PUFSMRuqw
1OuVgyJV+QZuxL202wEr4QyenCRQt6l04tvZsNsdGGKsNecoEhVVy1T+6Yz5F3mT
sGx1aZ/W1GDlZO/ElQvPXyNABO0A6yrvPNHDhO1SuUsbf/9+pJHDMPjK6Wzi0mOd
UG2eiDSMtEtj/u6lzf8TAGX5+zco+zsILKJ8/wnEbEpmjWWPYBEakr9Wrz61DOLN
DpGm5qb4zYtu7glRlwf0ndRrYjaTwvtWQqNVjUD49UhTC8zhrUOkehO0IajNMOD5
zu945ORTA13OU38nOrj7v3PaAduSpbMHrVBJz4r92JSEhdKqtBU+U7rWfatDGi6y
YRYfYg7cjOLCqxF6688o+hSn52/NTrS4hVIcxXb57Mnh39vkgDAAqpPJaYt/lcpI
xeXxkXOy8IxQVbHl7Ewml4oWOtf3mm5NjvuTfnHJDLOAXYhCx3Rg4acXUUoy9bBz
rE/L0w0XeHqbT2B6TWLcNMmJB1lYyGIAzDLWmSiUMye3wlju1TeupEMEgy6i5v+Z
8+wRe2uXXSoR7dnxNoWzlicTqCx4OIO11BSiDXYSv29OjRlqeDa8xVY7xvGkDCkQ
YrEuqwr3LWAK8Vaxz/SgkDS8DmfwaraRQGJ847Cr1sxqnN78lo8DY3Qx+R7tcgf9
9Xs8oeUeHdfhYKyt+kE2IXeDfqRoPw3IKXeB2BFWepvxSmAJqsyj4dEmvblHITNI
Lw9BdEhjYJMTv4E4dvw/sKCrmphEbi0D8rFMntUyAxAD1rJzB7MngKutc0ksfz3F
mwscro2YfROPSWg/AtwBVOu/DE38CjQ4L+dW1j9wfwS5Dyno71pZbe4yggAw2/Nk
bQfnK8ZR8eHhWnmnglteXVYuDvNukZ2PdWcdA5oFSRK0qBrqPSYC1GNObUZT54ql
zy+jAAKE70MQwptCXntz35HnPJFEQQD2eV554nfP1iQJeUEcAu7Ac4W+CkNZS8B0
5dGuk8szN1s6axtgPZVkdmKJHr5Q87GlUKZn2pBV+jMcn66Mrrw2qfMPYhUnUYxE
A0UKVGG7XD7ABQJi9JcpaI8C+DCtNwK2hmocXQhesxLObCZkSwFGWJa1YR/mUs6F
jlyustLGmDNbNARU7QKJd8WeXxrClwasDLkxticeMN4L3N9ko4HT8RBf6DEeG2Q7
wlQBq/EkPSDpidyyRWL9///grpokEMDzyZpBfAh/6dgFkrqGYP/jtd0fdvMGuyJh
K8dgOGKc8GOQlmJC3Oc15ESUFIkDhSKA0ho/0umR3jbb3mkWRmHC3AglYl+RFodV
o+odu/ycikliC99WycVpNhbZ6QFyVgQnJniwMJvhuAHkVkN8+yBZ7i72km+8JHJt
QNYhsky3HpUXDlJz3tFg64qHQ1YExblx7iIkhYAvLdBmDQBtogAb3RlgR0wcN8Ys
Na3jZPa60mz308c7pGanRmmfqXSdct5mw4WGyc2UgqX9kv6dNgr580/5AJIiwieX
Vh30ogoKu2pJjyXKmigRF4Z3pW3TNOXvFI4BHymgZakN5o5Sesm4bdSYCKjLkkg4
eer2q/XwEHODRi3QKbxlxNd3OismzfyEeiRDBjM0pFaESvleeORsgKYWvYFJ7CVN
a79OX2kNl7kvZ04jyV8TUgo6OMkBhRB0z2Ee6zqlnbWmX5e9lWNEy4vLPcJMthuu
gqQ4+bXg0MtlUDtJxsRUdmbvaE9LqHZzT8F3i/05AaSxAy4j0AEqN5gkf26TrFWL
NzVTkB0pa6Ew30oGNFy1KuxQ+BT53km7iXCde7cLe63AdcPU+yCRm+Ogd4UCgXca
NYBfWQ8BkrDMxi2wW/HPwLUizpMDQlTmHzPSxVlnjFM/d1NIurNbsEr7SVdDi3Uz
5wtMcsrDZDP1vPwMowv01ZlqEqfXMPQVaZo5WNvFYG/Cu8bVwqsKPGRSYKZrz90o
7uxReWiIuWhwOrPV3vWn97Ij5pTgkoQ278MenIIiL7WdvXChlVbOPflm1CpIzrKy
Lx/IrFivCdr4IMQK+1UVZwwVjfPHIFAlVRw1DHK1I9HmnOEDZ4ih8pwNaFP6RBQH
gS1JQXi7P4TQNG6E/a5khohxHejLJyDEAWjoRa0CDcq+unZk6y7P50eDqWqy1aYT
aJ/VrY9aDUBg5Ih6JRdBwqJIHSab3w9f+yeZ5i7l2xKSLNTe30GZKUC9vxSkmYtJ
+F5x0/g2ZHrMrT0kibIORkf8yp1s4QR7L2fUEkqXcRE+yTePhwV/uw7Sz9L4gBFB
ALweBTldOLwls8Jjtmw1v7tOqKo591DBPLZC+wyxSsr+4RG/J2I9VqpiJNEVRX9Y
3toUvb7aWdGMjBIKZgJRh9BKfr7HAa8pyCsrQwP2lW0B17Wll4EVb3+pMkXrf/Dj
yHJT1SJggOdC34fnAfurVoPeRiE8Pqhp4dDbLJjJgqShH8ysMpQohG32PuiM6DRn
D69nLfqfkUL214lFp7s9qCCPnn4J+J5N/1reaka5KCS4niQgZkr3Tvz/6RGzckU2
ibgLkOyZLmlNInk/ERzfnO4WxX7yiRfT69gUarDLnZfALlOYu+ZLJswe5nOG5YMN
4/xwE3AdT0s5holuvEU5EAHj2WOGQBzs+LJOGZCK621+2P3OkjcGKitpl3OC0NKl
Zr2D/D2mjkWH4bSbqipuWWv8MfGZdVAj1v3+E2jZmm/XG7zcaGiEaDBSpWYypHUn
KiF4Yi5AVppbboxwaiCsYmVQMuleoe4onTYr4OJctIRsceHKveXBdhY8bs9JSN8O
8/eaZK394TEY7izCq2JEL4oEbqK6kKGOwYpNadvCaTwGmgjf27x75NncpJpbdafr
yOWuL9CdevxlJbqVQzojqtqCDvFI1vsjprdsgqA9LYPdyqcBoivu8qg/eaAev5ct
bj74Yc8SS2kFla2G3scmKK4M7zugBD74jbuaRoYbAcVs/wD+XiTdb+l4y5hEpYPg
wYdQ6rfGXuJiSJZTYjLS7Pyak+GF4cJbyDEi9kvnk6BtVLzYHQhLnTwtPGGMw12j
uPYTbGfyoDovLyIOFdgiqDpUkApQTLuyhgLeRqV1/BJKwwVC9zhPPks5j9pFzrm1
62rAl1caZy/2wJE+uh/CthmdG/Munx1ObLdp7owHWnf/N2CJf90i0pgvAHnMPAmI
epqpbkUZLXrLQxRi9DQIXhOKXlwN5GpDfkbSuMDt9XX+tlkPQrLwPVRIBVWESvdZ
xwgCqxsyEiiB4LDeS0WwJ5EsNiyGFCAPAuk+2slCvRgDiMohE3akk0cyDgcRy+ql
L6yjqRxucjbrhLUMml6uJ6LwFAjZt8+AtgCODsXsTUEBnFGXqa3cnFa3mcq6h/oV
jqKQejX0Mu1C1wv0u65ZRAJZOx68Pya74Vb/WjRlrJ3CIBO62oZ1AkBw1Sicof7s
xYa7asKNDLWDjLhAtD97LiuEu9EIJVTwFgkNhayNM90bqY/3/olUjlcRlAJqb5et
mdvmzxJh3wSudKC6s5I8bmVe4kKXlPTrQS6Rl2/6KK1MgPduDF4rRFETLGGCWKqP
bzUm1XHi26geSobcSP78R/HczMsFYnK6V1+/94VHXruG+Bd4hND/e7vq8iIgRiUE
53RVvqQ5IJ9XBnZGXcYYhFBG2WT5i4OYVTRmujDfWEXb2YtLJr1vscYcSVp4PxqA
nglEoGyiL1V3/VKD7ZAw6Zn2pOV/bZ5qttPGyEq1i/RQ40T2zUrqzmGNz+DMpFgL
32vHXz8r2ZUSUSelh5joBE7/nNo6cw7Eyg7IHpdaGdWSoJ7tHnK4L6TYG8bbNifM
KFG9d6avo1zno9j4eK+uiz06WpFSpzkHG6+2zvg0RPDkmnY2Y7s8A3kP4uag2L8J
jubvKZf0i//JGc0H6SRHc+YACnO80QIbsjc/okiQ3KIObMkpFzIMjD0MhwgWq4Oa
3iNE6xUS0CHjLbMYQDqH8agR+hPD6wr1m9SAvfkiKIMHItH/qRK6rqfqvifgoq2S
zMe8vygtSZXhN7j1KEHTXFaXOTZ2cEv7Fv10iSF7DBHTWnyZc2kPc33BTUfP+fMI
XITkeN2WbdHYNBOfKMAuThcl52jkryBFtHYpqYiJeSkjDXX4I5M7U7uq5rP/u4Uc
IvNLHNceTwtxTEF5ATlbXPRGe45mcOejfCs45xm5ShGEouIt070QdadNI6PlvuXz
EF6X4P/X5du4VRBHacVGnAD54DUvbjpZLXGlK/g07ZAr6JfiEVEc4aPnCUkCHWh6
CX/fA/lQo6iApucdLmvZun0rzc9xAWikYDAj7CUZAqZncfFIZffLWQKQvcu2Y+FX
UZNMpGmqQufwWBVv/JarTB1yX4BnhEplKkgFkQ1d4A53miT3OT2LDT/c5EYL+F1K
LE+XxvNttpwV3L+ItSA3F684RO9wAfKs5LYIJv7vpPzHKVHDW4FyEHSQmBwG8MUI
zLI+5RFHPUoVzgQD0nKnMNdNHRd7+DfY1RBMBLow6eq5lmsoEGWmdo33oSNnm+Wk
XU7svJ9qOFD2carQ98kK6bW2bQ0s4bhqHmLShf8vS3zqNYpFM39EUKpDpQv/lysC
V5J+Em/P0CIYcanMJek7M6dVvGs5iO+YdpcFLyd4YfjFMyQWb2azr2wjEdzo6DZI
ELAg2rasTnlU7VTITjIDGaEosNMSCyI2uZQpCAOAFOXdIZe3s43ukqmaqOoUO5xh
uioQpUCNvr9WaoP+YATUzSdgqGpwgG/dvGfCSextplKYBvW0BKcfCga+VVwDLvvI
cD/ULxKCM29CGAPab67gm0JJIb5+HTVjJowZSTJQQs2wOfkpuicpQHWGEV4x6Dtt
PejnOpoeNMhb+yrkjHRE5M6fAfqXqN7BBJdj3ubaVNNNpsIh3FFQaXO8bSj00rAo
wYsbbOlJvfFSTCWRm8TCT7SXK8D6DCN1WOCD6/NA7RzcnnjxizxjHxWhogLgM5qB
HIQcDRN+yAwFAk/urUe3jMz/UtvCuQ5UTIFDcw96t99XZb0fVkY/WBUl4pz0zyan
f8xxOKt/QJ4Xwp+1Z3bPzbdsNRiwrkz1C+exOcx6W/GuQFpn99/fCh9tFYYYiI/s
UsBqPMdftuIgP3XZmG+ANBcygtqyIrJvydWLX5YJfchqZDnySaW9iysHMYIif52K
SfcuW8u7BKD3qCJzH06JgEBVStjnMGOK/oStQE8XaB2Db1NdubU7W7JY0uohFbLH
SRMqpdHpV2BlRwjc1SZD/5K3FA8ptQN880iz1xzBOlt7NQQq/jnTdQqouheJBRYV
VajpvqrTJReoPc56yFVk9AkTXPemssxBUzvzE/Gr5WqGib6tSMFrnsbCcVbhdx1B
8aevVr2r5UMecvxm6QNHFrm89MBpaUBSs1Yq9Nkwgs6msOTxE5FqHGuSBAqFpNqe
a07ka6z1yw6BcD2vXb4ezklS806fKKtcKDvMKRpoBgphrdqskl2/gX/Jkbp2KYx9
lbrA1wKj9DsFGRZCpEGAJhS/mSqU/Bhz6BB+DqS2lIX6xF5grixiHn235fs396FN
XCxNjYX5cgVITQ6JOjKCFY4RPp99ZIMvn9x/XMrsmcMo66sf2bPM3DiayQ0zJ1VU
dogTKo3HBZFmF4KREpEFphhTMhfpiY4ax1oULZCRWffq17mXDdR0uf/LUryXqFWJ
g9Xy82WcCVXoSfF1z+FAFFdVhAmhDlhIoB0I2kDlua8x4QoZQ+FwYKkbSNE9xCVM
7Vi/IfYf5JBFS6Ed0xfU+z4TzFMIqYdpqiKid1YJ3BihaJ2a1Hz0IkrHctdqvXCl
n73KUugMrKD4TC5tF+zal9Jz280awVV/t1hz5HvkYym56ff5Sx3yeBsymDDkVcT9
Oky1Ier2XRoK+PL4BNjU4kKvxc4ipUPX6lx3VOAOcnCzEkziIHv485yTYJi/2euU
M+ZlZaVQSXzWrzdVMpjprVNLYI5W/MFEWDztUrV1qd2EYVFmSVdbtcdF4AH3vFw4
19Vo0iRctIokatqOz3BhTpuXBXHNDKTZw4cIGfNXF1DsCKVcStTxIfOu51krKyn1
T9LNBcxB7D8J8a2IaR9Rrhe3bZYPHH++/+zKDNvRMNXExzWyEX43yUVrmGA/ZnxX
O/43PmYHRULP6FhsnjO7K8jxFQ0oVJHA4+v/AfKpRDfQsSSMYSd/+YE7AqVcDCKD
RZsrCAXjBSOrqi0kNgbSbV3Iisjg61mjhydPslfRDJHPy+MOkk82qScg2qieUyTl
jsqadW18m9pIVv/l02vy27Lyo5iub2kFszJMby+TdRD3tZa/bUWP/6wmg24k6fHu
jcKj1yCR2o0iRlWxZhCM0YBsUt01x9SDZgiRnFo9Sa8SPrB9smg+J+3Znc0bALmA
mMb4nqmaQVMmzIbV44r8o8KWVPaz/5MWhLHhUjC1fXJNiAt89tmZjqmYOAMWC/PO
O0kIYha7R6VEYeC7Cm2l81EgC792IsXysqCTvYykGVMDe8HP95ibDVjg4XT7LSdO
s7/05lshv0WnaGtE87Red/XJK9N5GDx/+Dl/6EeGUcbMKyYhTaMGqD3KW9zsfKC5
q2aBACAzxYSTiWVZ9TNWdzYQCBGU495n+ZjLOZLJ5/7cy5BKED/s3zYnnz4ROFJx
YwL6kp9gxM7uFbS9YCPGBDlijNFo8oI1C+duh1VjDg1xJo3wtm+RC6rbebTvirEg
3oFYVNtWn6V9njfdFEVi+5A1XOn1/7WwPVwh1YsjgQ/zEkqwBmzDng1K+IWp4xcP
qlVdMdPtBgFIkK7ddk2FGSJsZ1AnyxwsfhHWjg2Wcj/BxlZe8qhaVaMwpm0KUMB1
1bvQC2TkgEazYdthyIy86CVLfJZ/+X2Zt29CO3BqydGueyhxXdiOb5Pxge2mqci8
hhEfUJ+T2N7XI/2QqBAivkkwh+N9sfQCoA3CQtRc4qq0n0Rzzm2YKgjlYz0rcxOO
xTWPabblf8F6CjIga5j45nyWxHQfRoBiLXwiz2XxB7PO63AnQtv0jGdcPOwQXqmk
JzdqXO6B87ZL+EPd4ygbeAN2cSIVrfunYAcoCnj7ixYv/k0t/9r6YuI6Jm8eVvYT
4VBIU7LVvMfMHrgIlENLoXO39UQ3ZiMcC3p1LewjDe4+UaPmGmQGLujPw0sLpgAe
2YpUaVDvGqxFdyf7rldZ5K4zsw0cOuRiGCy09smnVGuYLC0D0LqzDmd4xPc6IrtU
KfHIDPf/xeqEND3ipGHZm4REySuW5PO4TejfsoyxlRPxP+KiGujzl4XHlVHY9LRh
v2eCWxqWu/E4OJMxeYtqsTUVnIWPdA2wLm6s/XU1k76W7czzRSUryvVxctBoRKyi
g/iSm8bx7yYw42t+a6QF82fSPYRP1emq6ikhpSFrhWcJ2duzPlXgsUUxqyNXCd55
W3lN4lyMSYTtRltPLCT21IQOnInWK+aIUEsP8pE6pFxGPtkIV7AcREOyQjPlXa3q
GKIOu1e2eglayXVf9Hsi6WgsC11mZ3C0hvA+tmFcxYivIgem9lcE3rFzv7qOkeCU
RDY4XRy4UT50LhqOfQkEG0nnX1jlt828Oj8lVsqYIIxR+tQAvzQJ4IwYFDDBYp1Z
G9Sp6TqDP2SADdm5u5MBN6FZTXtFq+D/v7EfA1kfoxsTymjR9GLfDdewd3fr+6Id
jDhC39urNG2GWc+7pWTDPPTQ0DkY3IS7ZjAgL7XYHPLog3EuAX/78WNV66s+UC/o
Lq4tQtQqPiJPk6b4lVAEMz6HcMDn99fToQ7E16CgoqNpYZ/bUwrZHeBNUWQabncL
s5cjMqj9fnw6aioQrbmJLLRkih4WIywpjW/peM3t8cBPMds/xDfQ7AlF57tjPlHI
YGMvkv001Zr1jOx6ykTzpdQv3UeqThtVwfb2wHqqWWt7VtUJjPR5UuujmW/2OVrY
ZrjvuMpwlWHuQ+9GxPcD1sQX4Ok2jgYsR23+z6iDA9i3jvuDF5AWOe82FJemaCrD
khCIPiEUiW61tt7eCro0LGdKitaXl+/UHHFb8KKad7FvNv1fx5+OpdKgpgQOf2II
dw//T+FNDqSg+HMg78Xs5EXUnYYT2LgSAwVmqEgBpr9UURnJFaubF5CALGF/xJGU
kpG6axzdYYxi68UHo9whRUdUSkvuXZTRoggvg9YOYSahVPfOwhA374JwInA4rOG6
jidwfJV0B+rWHsnKwilLh8BXtbQXLmBr6Ct/1PJtnb3qY26OBFCXjKQaK9uR/PlJ
bu5BhBIi4bXg0nRNL8Pt8Jic7+VEmTpT5lcB802yRMFHst8Gh6KL+50qJicKd+uH
TyZQyEnNjTVx5ZMcFBQJWuMubj/X4ABVw+EA4hHwH7g+sfwW50+2S/hsP0F/UQ/U
5Q53hFMXPPljjoNWvd2RP5SPIGoiUSdJrnmKd7qH8wlzm7501TRxIPSjsnVsflGO
CKgtR87xPo6YgvE08TYnbhd5aoPPP2eWf5N6oK/dszm5LkJakgNeIGRrlgGwAjI8
M8oQxpEl2XdECqbbDQ+8MgtJBGJdPw8D8byKFa+GRHbOhByd2PHwI46GlKyafmuf
nHHXd3hpHZpdjAr+oqP9sHkLfixl4rIG5mBuKH9V/ixR5B1aVlQkcuiFZaQ575vJ
AbyDGmpePvmmVEhdRNkFOijNtHQnjGanVRuAjTxjmUUxxn2NeK7YG7WaoRnxH3FF
7bBJhqCy4AbhHFgK4acKusgtNI73DwlrOjo30ceGYaYhQP0jn8kRuLzCTswP234k
ZOFZkecUogCy4fHTy6kRqka/0qvhGWC8o+EnlYHi6Es4NOTtbCuNvgoWm60QRYEU
4oD4T4cVmyVaNPG7keGONEQDmTr7AoLGrTwW12Nq5UmBqy8mNpDEEexJXknOcr9T
7EDiPHb9zK1XTXG6vk3DLw4GRh4rlY7IJdxqn+wHC5Y/qIg0ZH+XET83ZxoZQNab
9VwKdM557LU/GE38gmOaiyA6PG2tJfA00zJfVCMNd18XU2Y4GJHsx0fKtMKZLctq
GRzeLhfksVOlBnPHRUnE1Rws7SHOcjEDSp0mw4AmsTKP0WtSiljuo1znQUYrpjew
+9NgiKap2pWQY2qvDmxqVrsk6SR3DQWeSepuaVzch2C5PNchAnzOLJZqkNdMVrcL
dDV0wzpNiWltNZF25gFhnMkroCl0ZyIV1N2bcVIuDSyXxeuIkLCMRlDgd+7Ioa3t
2qcNwjP8hpH7BeVrYQR/YyrWLi982TKA3SkwyOuEexnRIwBJEVvkiK6NIauoIWzC
BMjakeaAbO1bdIO8d5lSurXiVHpBHmy6HweR04Lu47miCfq0hzFEzGPmm+O26UEo
xMMtOiayzlEecQ1zgcxHMaaf1ULb6h8uIVjBRmIgYnPcfQsQdTYyVEulTPJYdcg6
1Oz5ehXeV7YzWHJkkQ6TRLsG1cdgM5+eDdpzJASjszBRXOkdWFuvWxPZaOgAcJR4
rFNQcSp7eyloJi1e/8Mub+UJQ95iUucdmBjkNoP4PxRrSX9B7OHUz0Ujxf9eqVYh
XrkXF2H8pL372zfTR/lqmDjNRC8KtINaCS0M7zFdNZQ6mgqYbqf31pYz4wfd5nzx
ulp5e9Ct0REoAeAMvuWUR5rRzSEjl1TknkG9f3coI4uPEH5SqpzJo2fRuA9eMcfK
NmvqhOLgvndJsgLf/stykv3B+L3R5Q32ffaLPaoQCvSgLjhZwM8qSLunDrUIPAkA
rnslu2riFPWoWXGiwkwr1LgXaJCKDpLxlLNPcAR5eqAj8kxcyrbef7OwGcg6kkJR
xhF68bVu5tX8uRLRSmr1MAoXaxytgBDXfh6kQUEmOamJxAyzwVUplxjit4LYAkdT
hC/EwJiCVBXiIyzNujNSX4HmfjVpVoQANbrkIfKS8Bv9ZfKZ+QV7eWKWiBdiYKuF
OGhwRByq6LTfWoaJP00BaucVXtrtrXMcA349tDF7viJY8TO6uIYgXtZy6B7mUw63
qHHrHcuaDA0+iTCUbYkCtsLMOqLS/RJjOzvxIS9WAROCLjAaqN0GeM8Gc32XLtbU
3PlSbhTket2QclR1IT4z3rJu1T5NlvScfy/acsjzgCOfx+T1FI3wkxYjPU+ELQeH
PNiFMa9wACr1UEN7e0r8FMlJPH/7DPSzxJaZNFzopBZfqOnIGqQpC9TR+FjSMeH2
L+0ng8kcHuNyjpqpHFTihOVNwLXaSewTtf4Gi2EmsyomRtMOdLp0zoBNIcV1FJfc
2MPF+S3Nqx1bO1/rvp5LKk0lLluOdVmdBCXfaCFkXlEfvh0zVecYN0fbDvogG9DY
C4BFx7qFw+guhB8/6uWO4ORGukNLJ80Vxf6smUx0gBpXDL8vCbCqOheyyOQ2iZcJ
+bu7gaaUhjTsWG3WwwKhN1la0PXLu+atQwOF2AEKb7bAH5ly8aNNGiEBFgrdvPWn
EajJbZ+Ff7UXdj4ptC+49oDftkqDopTRquLVwZPozMue1TXTzkXby1c6LSFGiTUF
znGWzadLydA+HacZO+pzzn38BpzLOIVJjByesN1c0phdff087nXQ1ovPMe+Y7lwE
8A28esypdfxgzjvmi8rxQrEaGAhz58enDInIKcFyKha0zylvjWPlUqqpBRlBT5r8
z/Xk9N7ES0O0B9Y/T6+iUscKPuQMm7eN4K7+ropNvDoPcDcCWU+CHY9xqMaZgP96
GeW/+mE3dsIL3iuHXTzsAESsB7LDcOG86bF2Oy6b/VfE9tG0ldDt6tXlQa6RItsV
zI9m12eQlInd6xh1nZIgjSjmcMeAJcGl1m3BQ3iso8aVbVBErq9J2oZq7ZCTOxK5
1Dztznqo6vZs3pU32xIywDRrih70BtVnODNjFdwiKMhTGCKUMU6R30ZIAcyd/Ihb
UKmFx7hLQBkfHRSVnyqqom7/EsioKra0JLklCpe5F+SnlQElNKkde/SOoEbuXN5v
JdTihjFH+wjxVSw1szMVibbzY9laPeYKd5gJ3yQzsFnBmNDWQNeIl5kRmcnvRVL0
3yT5rEAo/vXucwHxyK5iCgEYX4Hz8aCHXheZDmiRd9oUrGO0VERDwiU7LbZ4e/iW
9c0EDigWIvAkElDerBvFX5XjNtah55rXgHi6HtVPyxG3eVS043ZBX06PHz08SC90
Afp0N+3+xDvisftn4p+cOHDzSce0sjopDM0hlDZu3QcfVUYcmZMslN61A1eBBUNu
JSaR8GiC8QtZ4rtT+TK/by2v7jkmcOXWJN9EMCeJSG0tVwG6kWZfrE+r6/Cw8RPO
FHFep/IXazR+GFhiGgG0f4rh0f7ItJoPHi/3CpmpMCj3VT3ZPrR21aaeJljYuOWL
ZI/hJhqGiodsgXPTFX1K9jVmWyDBdRG3DYkhSpXuZTI6OQGJivMlmO+vUBNarW1q
16pP25lIM4nixgBLxQ+Fyp8uC06dNI0W+8edf2/rZE2QsrK9624x/rLvoJvlombx
nX5Z2XEN2Dem6gKK3rgDsDAaRqU8amdBwFD+1BjZxY50mAk+nRfHyneT2k3A/ae9
O+021+PVqnul5Ddz2G4hlw0+0GxznlUu5VcPJuym1naTk2y1zAZPGiuu/aLBefL5
E11x0ohOwUl4XroCT/ukP0HCdRktISWNHLjjuGo8Qi4Ww1GySatL4Zmefyub8pAj
sgBvd8oCa7TfOXGtWzUEZT1FxuqXPORvEm1+DTlBF81aDaEaIXO/Pbe1x2HPFv/m
urHmlMRpGbe1/SEbg8gWCvSgSwJDvQPT8dFBs1RL5uRSIw2NOE2cdo3R0x1kiqnd
rIz7gGupkSnXj18XJwciUCZB+IFjhR5b+7D/aqN5JqfKBQVT5BfsrtAB453w6U08
iI4cbj8JBfaITvimOE86/ff8KA46uR3fqnriORMoVt6YpQL46RmZBlnKoREpUtD4
plcY23eXQxG9VMrE6rljNWv4KIiSnU3RIQnZmDlOaw4L8IwIfjhdLVgh3Hwf2n8E
5etQDlRtG54D3ytIwaLTaU3ISFDutGdys1FHzA7LqUI+FipTMtxAahMooiQJ64Ji
sLNphJBdn5/bNcUHEE4WwcisnOAYW+5neHF+LeKv4NoDQotV3RBH1w7Nhcp3ZBr4
pOaNkM0NuglwexmnL03UYdOh0n3G+A9LXbQ+ah3MWxm5ScDhphjf+PF1ywz/td86
uD+SF7FWXaRvaMRnVUs63C+pFkPBLsfDrUVmPZG+ajpMCUbu6RxMptvA8C/sGWQ0
0YVXAXNxRSLJHFFczWWZFmP/jbabzz1sXMwhdu+kavhnHGJS2v6RD+Mdaglkh6FY
woTHjgFSXv3AGHm9rdDYYC7O4QFeJ9NYwLb1rpHNGKkbmvrqgXjCZ8zhJRA71cDn
dqdRgSFoeaJdhvoTOwC47DZb9Nc2mVi/jhG7vyjzpZIVnMqrYxndqJ2bVCfQgYgk
onlvbogPNi59P9woTiI19HloFqzgPKeLjaYA4ygthOIYfwlbfOLAviXt1RDmUcVd
De43yTrQcTDaR4mTKgNnbmVaJV/MkuaIrFX8HTvoDdDy3ayBrLCtgvtz+AEFqmR5
IoNOH1+cg27vMxNiL7kKVOcA3F/DH/Tv+OUwPDY56ivb+UeIp+8ZS5nxoeN+NoO+
WrpLXBSbQDFnSLKjGjQihdiIGCfktFO3RjsmFwXyOZMH1E/vr12vBpnhqd4ImLQF
XKoC1tu/ifgPZ8IZVwy4gjd64RPcf6/m4yCmhWre4DYe4QHUDs1V3dj6OASCQPM6
gzSF1vBLWWaQjKir8sOR8WmEyC5YBEA/Jsf+hoWrEI9dqmU0fegJ/Q+40CnMb1z9
rQsq4jxqcTdKhoEgANkDbWdxnKD/f9jCqzW2SSgLSHz67YOOcdcryhqbz2LQ/JMs
lctFiRIIxRGgipmIwI1CbE+ndoOI73WHwmWOtmmGUSBo72BsxgoKTvvna22th0tl
JQ82UpYGepRjuGcaRkehhLHjKmdvyX2xIDdaSVWyYszFlQH3ord4BKh9mltqnMGp
Vo4wlERuzEOc7mLnQtKdBLIb3NBqHhcGROoUyfvfuDLrvY2xNYQp01xZipvTgYxl
SB6XhHiO1ZTfMxNDvElJvxB6mgoZZpXBSTla4cLDzo6dPDoYU5OMUul3b5O0r7Xo
PQzUKWPBtmFQLwgSqTeUx5+H41vr6ynYxLAgL+PYuh4ygt8Unp1TKga47/PeKOm1
UjGCHfN6sXcgViM/tE71bPwcTBKvtkYnTDCOTVdnMGpTIUXcjdjczAOnQKvCSdZm
OZqKlYdhekJ4XHdnUpZ6V6f99UXw/ypug/eQiUmbBvmie91iGkkzhq3dIQm2dZi7
KhMjdcHI1SC5zRbpssNGT9F36zW5pceHR7reyxrPfHZzCp4IEBEPk+awZgWfQAl0
mFO2tnvMn887R3/Uavv4Yy4m9FLdcpgmd2mFRrUCn9bHyP+wG7bjpr7nYqkrz7Qz
o/mu+yqq4mO+u7v50eRkt/Z4c0IIANLCj2FTUPvZ+BvX7bgufhwpEm8EiqR6uYMA
ULVvxnM0KIpSiVYVLcyXt7rzGkM6d2/BseMlzCum8ZaA45BM6TVDSLxNonjzJc5e
aiIzG9wq1WX47hS8k56GS/Suz6tmRMYd5MEzrqkJD/HlCbaT++PG5FDnJrjRA0Bw
UH+O00bVOJaGJYJaYHw1MZyiXiJ7GIvpWh1fDujFf7StjuvFEd928eOu5Ob8R11D
Knlve4l7X2sjjpnLifYEYUUw7nTp5QhqjjMvBFCuzIz8KB4oyJHRfbEVSp/JlidV
nPWS1spt5tQ4FKZkm2kUuc1KYc9CFxqsMDSHS6UDwk18LfgQVLkT0bV55bTu0SxQ
RVODaANMFFsqV5FYzIEqdEXmKD+AqGB8sf/e81Qrh7XfRZcqLR7i8oqQ/Y/+eEYj
O2hgE2DYV2AeAdh6x0nYGZhFUk6SnW9tLNZRZ63frMazU6MfqR0x+O4oE57JTyXk
8pamUrHA909oL3yNqWlrl/qxvn193dSVc7TrQKSUMEvTuvmyjUzanRe/bGvfsqUQ
fZW89Hc3HyNlWt4aBPHdC7TtBWVN1ZYvPAzORfVUdP70ItlFatWQXna0aB9KdBH8
WFEXAbg5x7mrti7uP2QvEWT/mSSlnXe6lcPyvr4BV4wyWwcf87rzhC+qJWTnSJCS
njivwxqQ0evK8WDZH277dL3gtxk/+ce6413iSqKmmYeqaIprJvuuaeh9de/1thKT
70dGoRKpxCvbfLnIwO7qcDopQ7QIGvMtp+ThjkeNLYSZUySTpdS17t7Aw7OQhhEZ
4TeYAdhDmtAAmGEAwn3EW0yEsYz6rr60v5OlU2BTbyyAuVHEZ6nt/Z8eo4cGOqh5
GVjEbOvgLhUAxnv8U4DawG6r0mJ30WIaShuLYsL/n9CXTWh+etK6XJC6CDgCRoo7
SVuAdEeHHDKNWkkWhZlzOt/7TFHq90TdVvf9r1LLAD6USBZ1CHCK36Y14aCthzaq
DfYOlozhaVTzIBnJnOxZEu9Yw2OKWcfYn6ciNvVAEA68tVE5Im4o0rnZRQ+y9YXh
eO8QkwjYS7N5QVqK3cL5MPXppIt99ohzumqeeLJ/LKYOkA9dGVK2MTOYUYzYL/Vi
9jkaYvowHyC9/4/26EhW9A6OeR+6A/u6ru/xLEBcpmsFKqkZhcR/2Iqvxsr0nxy2
RpUOmPqzGubMtcQ0ZxNMmriXKwk0mhdfE5DIzbEughiiODywkon135P3xrta+nmS
tZ8KFK82FY2lKNZWCA+esn5cHeAKHsK8HJWiZMx1ADFQhDK8w7ZjB1v84+GnGN+C
3k7zxogLnzjQT+6l9dCT5jSG0M1FFnkzD7cTcN1ZKZUR+Ss6XafpoMcZ+HnRfd0N
sQ++px5QG7fI7XtiXPCY9irIky/3P8FtqFTEcgly1smB9AVgWgt1BDpXCPDQjvL1
9zSUIrU/GVwhAUUUjY0cliYlDOeg2TZHBIkiREeU1SEjYAVXy9d9Iq9LWLtyYeJ3
NNiIjekijYX3zdnOauopy/b+PAMmGF39fR4zds2kAhNz7UEfU1VfKLnyRFDGwmrf
BVPT9bVH7rTUmutu3Ywhd26XtThzfNp/UaGx2RGi67XmH7sRvYJfj+TL4mpTRqGq
LaROHH7db/MOVRCChmYOcGJFa4YeJuf4wvkHApOHevWCp5KGwVCU8W+FnvOlWPrc
3j9BTWJs6hCfyhM/aKJLMLNwnGKVHkrVNBdM2ZgRncc/y72cbJwMbvxR2sItxDkH
ZbtKFPdDhe1MhqWYcxRgzNsbEFO1IYu0TL0646ce2/rGDA0/GunHx2kv4ixA1/Tw
buJRPd+8gHh4uDqbNZCgYjqIIejABjHS8XCDYGjuAgPd6R4VHUb7gQhYr5tiDBYM
7po7Da30a1lOj3X73lQi9N+3xI6JHrwTNLGCl10bqVCkjW+dE44Gwy76N5xyw7a9
6u74i7HbghxVjcgfhiPAhSNSyYGSXWQEaTNAQGwq8F6AcXAOX8vahcOvXc/kdetd
XP+HCeZCnH6EUCxs5cXEdBjvdQqJP/A5scol2iiswB5CTg2IwmxZ1CX6XTvuYcoT
3QPszgJ2loTLtAWxcQ86y7AguBRifUxN65Mx7hPy0KI6S5VvgqpdC3zgmqkWcoLv
GGE1rYiXRTbkrXwYCHm7zLVBzZAmAjx3eCIUJHHe/sKbftMQYRKga9+JKvQzgVf8
yQYH/O4PT5atlSp8zcVFmhyuQT/FyBIUvtTRJ+9SLx3BH24qyqGHbcjB1FM2CKDu
b8v3rFMcidUfETdKXt5+gcTqtxZ7XngVxdRdGbt72ReSiKxbnXrAd3KMRcaxPHn0
R6J1gqmhhNAwpX2wT6DXg4VxAS8NnV7PslSd9QpqI4lW0WG2XM8lQwDb4oRjz0cu
WLeq2xKGU0+r3CZPwm+CPktxZAAzB0oHE3fSbe4d9Uex3Tf9dOuPwHq4lY5hiU02
SRk4/954fFEZ6lbpi66LH3WnRphOdkqvecLYClB3WrnKH2jbkmXt05W5fEQbAsAj
Xp3Eb2t/4E3eXgDAdc8/dV5vvHGlt4+G0jygnW9KDDZT7S26EecOO2GMk5sHK2kA
/+jlQFmqe2GzTBlnxFGyvkoPxbdHXBBhDkmAHNhY2yUkpbbR+CTLB090zARAL9HC
5cy8Dj0AbUmVa4iv4PdFb8cgmUguNQCsDWwIVehK5KkU1N6etNb79FGQTENdx4vZ
ga6iAc4ZKgs9ufiNZVhh+taaNzYxwBGXt5Ime0UXpgmvtzjHd39Ml6Ej1DQiOIrl
pLV4XE5qnyoqsAy6lCJRCGBadtNdobBh1goc/Jr0Z1wIuxurDHE+xcUCUhXuInyy
TNFPBwtDsxdcTicbJTK8sUXgGSvFtwre4IUVS5C1RgP5MSGo5edEVcAZxq0oy52m
2Q9lfoATSHa3v5OSrPg+o/+pny3X/ucuyahvFAJnPCT06IjMDT8gF4Sa4xAPLJEC
r1x6L8DRxlgOUvuIInuWTMciT28ppa0y3ESf2n5QyVT4Y/57Ki/IUe5JIz4068Vh
yvIvVUdSKcRAM4pA/P0QSfJ20zrmrCc+ZjmfdsJlX9Zq4fsTEQzKVq53CyU7JNP9
qRQAsN5ufMQ5t7JWQz0UaLTvYH7LtJzgGXwGd1TgzCgdpT7OwpnMdXQfX/rpIurU
WpFkGqLkmQNmuVD8gR0028gCqMecDAXTzR8bA5dSnXGQRpJd0diglYhtcP/KG4h/
y3Gp9K81E9wZpFvEafKhrm6Hmuj+fW1uB4WMh6KgkMwND3rqsBjl+VcwBrjP+vaf
YqrkOVn22sy/udonmXxi/iBUY927snX3ATE9cI6BDGovoZU7+fOq05JCW7tfppYa
g/kNHrXRbBg1kfMrA6uq8kvQ0FTj+c1vyHOGjVzYpH6/lVGyzFZ8/1pNtNu9mmtK
aTB/vcDGmCgyLtdhoECFhKiXzqa2T8qtp2oe+TZc47odkgYsq9IM8mlyAIPvtCGQ
3JBRkDO9lv4a8ONoWU9QmvBGJQF1ouoFfC6TICL5QTN7/jdSqHUjoNb6xtfpBFwx
K0j8ML0vrh6F1RFGjoiVXsa3YZNWWsSwIArTlbhYDy+53i4kk9BXRNe5bijDfylF
ldEED0Qm2udQ6GQZS+2Nroc1w281CZxzRqIeCZSLAhj9yWAkDUzWryhIoJpMyM19
MK+rrW3DB3Br41A6VpSVkWj7jrN/GcGazCKTQSNnZExEB6k1A4OnK7TQJPG2STRp
C+lAUmNL6XxywaER+kanWY7ipAs9TOcoF8XbFeEZjPsBfAq540dBxZN7pPa41FZQ
Eaf65rsA/cp91pCRNL6ps2EWBOf8y8Pxxy3SrF9NJfzgisjjiIVNsRB4uk2b5Z9j
JCXTRnnWFPOqdYx392NeR+uBwsQyxhzlkRc3OuNBPBbKPb36sSukKO5skb/Q6vlW
rZlDwlhTgstLMzB/xqnMiS6Eev4ep0OatgpW77yedIDxTwNexCoVlPs3RY2MHquY
OH5OKMJnSjO1lEAStnCawHlM6vxhIj7J4SoC+hMrqzCBxc4zFm9PIY3jHLxYx06m
zx/924Trv2ZRNGBKBJxHFffRWuWMvmn0/P4BpYqqpHDbUPeqrr2qY/zNWe8Pd8n1
1RTcw+MwoWvouD581E9hQS8kKddC80NdqaEQ76rnRQSvdOxLNGk9GPc8AsG8ce4t
LCtoQmuC/Eu1TCaEWPc4+lb2LPnRPXTilL3au4r9D7EO9gYsUkAPvlKqWaQ5/v/o
/s7E6iMFlCZRTN/qvpD2iT9xV9fIvtjd6UEcTdP7uO04Z730i4hUMpbmOPMqr1l4
pv3B4QT2TxNm9bU2+mBjyObMq1tc1C4z59JEnzgrFeNBha0ULETwnYiepPf9OBo5
HXEN/UASbGDLJvhbZGDWIpV4iwQYO79OHdDrdkshlijU5ImS0OEEsHtwuG07HylN
Dat0HR5gh/EClxagsS3Dr5lCjzaiY9BDOduCn0bohykY3WOBmE51d++4Hoxm80Fv
e+TsER3a+/N5927mosRfMtO1GpG2Nr3etHkauYMXrQpb5Fs8EU4CuYrWtOZV/29C
8b+OTHQIst7VOCHWc/FCoi5bVsNjXxNFF5NsbG421X1ULWDe6Ay1zhaKFT5M0JIs
Zlb/qcLH9rOmkDmm883Hv/nQDzetQgwKF5qCC/SnLPycUHAzQ6jTP5l/jDRTLsrf
ki9oj2lSf/i2PybTO+gVLUY91aNkK2w9aENPvMw7F1aQzdwzd4NDw8uUL/T51BiY
dADjHB8Y942kRLdoMNB0KeZxCg2MVLSpyum9DGaZ5k86hO9gGENKLb50f8FqPlSs
fLMAn2h3XdHjMdcq7DXMNXzz+ohRDpR6fnx7O68DU0/fIf2sIsr4ZeKDgI9ctJaK
J8xFarg+JGS/P/FZfIYP1wQoGEg6n+doce4kWnqka5VJ1rHg5fGvRSmxrK6fczOW
hfamblGMoWDkpy1axPYMaXKGU94UZepXS76bCGwRZAS1ilhw16lP/fSLhD7rzA//
pTycZ2VPpgNmBF/M9lzCXY945x/S2LoUWWqwrp8DxKHAqW0HDfbT4HsIq0fwSgT7
zmt8fxNehVBZOn6GHLSJfcrCn3bbYlSAv82hiIBKNpguElJHotwgQBJDjxccZ+nY
rfOYNHEBUiKtcCSBUtbq3UVMiBI9hKS+Lt4+JT3E/7j36r+0ItpplgZkHYCdEH4w
CsBt8dzVDXY11I3LAtYXbIja247IZuXwC5KwdH9lOe+AlgZv7077uZ2rdTXkm8Ow
GwCSsWDpE/DTf0+y1l2xKDvbTJduU/zg5FqXbJPnMdUHRbQGzWg/JEwKab2YqUkn
gcJIeo1PrjoVdHhnxpQmwIklU5oHMKsJ5UFb90ad0Yn2NJs4ajh5zrF+lzu0T3TS
wSq19/YAI7iItvO+cpbEYkuOVdYZ65mnNPiCgUg1IuaainHmx5sXv8EpzxdDCzzy
VizSdibXjEJ6/ku1irjejQ6g1Kj35Hmlrzj/OrQJjjc0TGBxfbvyl1lC3ycpd7R2
AG5IJezNJSxLG5q7wDgTBTq6dyMEh7U+0cttDpPB1fxrCfh/wLDLpN0FNErOeOL7
+llmmOIy7qaPMKxsZ6Yh/8jQlBaAup0Xee7TXuRR0iZ6u6gpvQiG5QEzjShg7Hj9
QKVpnnKplRNCsLyZ73J97M8Ncu/0C/fAvuUQMCbpQkX3VCVKlLhPUZ3OIO1txFWW
sYEFFG0WfDERPfHWY6JiwRlJ2IkQPB26SvJzYS6uqdxQXSllEEsiZ5Ki25Q1gQJm
BrkdH6Q2QB487mKVvV4ZEkzLOAF364Jg2AYNmBxuWsPUF/yvJFNCmLC3T9hvSf7X
DTX2/qQvi1kHJBgUjZ5ZolCvLl5pqRILjjclg/h0tSCz+cG+bWU1p5y43CZTBt4M
z00SGGb1E4MTF+lDlPU4Jl/uoZ7ot7CNsJoZN2Tw4GnfQ0vSegcBdLlTTIdKYGsi
s0LzRIQHTECnmRYHikV0qOipOEKEtbJ/5e0zdjdf3rD+yRnSzWXYhrCNiAfAdCAr
zU2C9c2V1j8TC0+Z3esLGLu2T1/YoP4Bpc4Ju1an1mBAiiWewf3u3YfyiMxyAK4S
ACyjf2Xzd7ytrwiQ2gZskRAzsbOZbDqaNxGXIFvKoKfolPcOYUSQJriF+ok6LSEY
jo9lT63de+p7XQDeV+mlVLJtMW44OZBCu4sEnO57uy3AP6C1ErPJ8B8n3+rRl79E
k32QJ3KkykQPruBLexn+oJFLifJ4EuqjhzZS1oFwFVAC+0Fw4U/UUHMxjwuZB673
Fz9JcyysRThzNLRZKqaXtakoqf5fYVMWnQ+bMgqGsHLTdc3EooFyNHk+d2bPMR9n
s0Ay46xkYqti7OLUlF24yt9IIO0VPb66dG8OVbim4D7y/+OmZfwROrzJl2OYB5a6
h620zCEKEW15hSimJJMF7PBNi/XClew9QbG8aJqka1hMfscrF8KGhwPecAwJ8fv9
lzpzqS4gF51n4PSuiGelkbU21P59+16jqtkuvE5nilolSwfyoqGW7DBBC66GI4+E
tISqI8gFP5FKXNRNUpjzMjQp9xWccxmjRZJf+PnBf7OH7TwEBBAH53yovxgzvTfu
oIfhh0yA30WjJAQ/qlR45trLOjPlnyejIE3gpYNcTrminrxnqfki7MUcbm8j3XVV
2CKAo8A7mlpD0bwBUmtx0034lv7qMQVa36d+H9XzQLB8y/dChVyQeAdIfVCJQHVQ
7oReZDVLC6VtHWOHsFxjzmKkydFju33O/ZyRE+DR4wWaYyhtZo799/YeSNQYmOQ6
3M1EOrtvEzVGB6fJTq4EJEHHXoKv5px0dRpjCOAI0ITQCCzK3fLNVRPmPEa3/hyh
CJAQ6KK1SY7n1p1Nc+qI8lT3c7HjkxRUq9d0r6UihrXOJaveY7Tcmd+Uztr9/rO3
rw87ibzP+87LpMcYM1BmO90mVRDrM0OklKq5yJ2jPoV8mdnejTaXQ+g9vezlLuKc
I+VRehoc51EP6rUzUy+5g81UjAVv+W1xArB2vEaWsGCGymOULIz6OrZufZD4ojbx
8WXZQBs3OOQ47Hok/vPHSNiJH0gez3lEc5pEYIz6JoW7v03UApft9OZ+DSQ4941y
ma1utB+gF/vd0OWOu7FKfYbdHMVxvRx2/rF0KEHIZx6FNR1VaWvNjgMDUC7KYnpU
i9ruelZ35Nkv5e2KPsaeBnaAV9/hp7b7oou4GYSe2Llx0Ebo2x/+HOyVRKs8UpDR
E+iKnkfYVSDBV+1Xdf+h55UqYCbLaYWm11K0psvcAi4VrVmZn4Va3hkHGqw0P+p3
mxLDs2PrE1tn5i708kn9MbJEYexDkfoMSMbdik689O0mctG88vR2V0fSjI0BOXrE
BEu9js2wHa0hCD4zcShIvWfW1NVvsNvTZPalQzKryiwThgfkEb4L26O/C66L7jpu
1Ii6jVWLpDLYqcqBuN/jdTrnfSmqGIXQwBEKJcbivFu0ed9IstKx68lr1rHuJ2ei
IPuf4idBYjyZ5xD/z+L7fvB/FMoZ4r4XG2tDketXP2FPezArDbAAll3phkCOkPUA
AQrfb7x9Z/JqWmh0pXrSxtw6syI6pnhBusolqHy2gPlo3Y4J6ekjQx7M1mqWp2WM
/TaOJ4Kl2lArHNJgCmaCqnp9ZM13zkohxMFr1UbqiNgkWFC2Qp8fm5dbVOgIrNyB
2la4prbFhdTivks4q8IaiE7MS677W+Gyk2slqkrFEbx/UnB9aOfdPHS9HWi2vgLY
PsYWkPsRAlHsM3gE5VS9WFyz/EML0eF2gRjk40AymjP3MQJj2NjtuGMWvMEYvF9v
z3BYtrVQUz54ic3CZ3zYRETG5Z/xQiUNW2EpmrDZVyu6v0lT2gTzlKBtk1fkwR9r
R3OZslVpVr9IdQqwKg6ox8WKQBdI4cluwSY8u+XduHEKTQuPEXGT8mGBIHMotCzs
EM+eyZtIztAjy9+/dZhPFHvDiL8Tj5Ypc8D5sgVB0hHDYKxBXyv1hmQ/V6/j38BC
qd9NhPY+wok0P7iS6awzeTa1nCMRy4yoSKbXF7/jXqYerQcjhUjVfHelElRH8kJa
1vOlVyzTjtSjXesdS8v1Mpnz/XDn+WOxTA6oIqb6caMedHpD2pZ4gEDWk4JleZ6H
mDHUSbXrSTBEkNPE7X1Mmm9c54LTZTeXUJlYKWfjU/eE2oDWEf9lJoV0xMFOFfOy
D6oRvLwrn7RG1VE2TIe0DVhZlXm9Pq/W8pa8Usxpd6sCt8lhUjbR2p4CWb8Qpf5l
tgkEucX9O+H+jWA6sQW8eHrXl2210Ioz71FwX/5bSt5vPwUuof6uvXY6ARWiiMnr
abyNl5nEuZmfoc7iS8lZrqydrhwTYStC3xHmx0JVIzZ+rBa6IBR4LJ+xpd+IaIha
Ia30yri57/5Qi0A/eajzLOROe2maLkTj2/wlOr0LbyEHVV+jRTV0Z/4LzyUw9VaF
Hk+je2ivLIrnjPWlz3ubGsfiP69rR2nxSArAD8CH+6zMgX1JpRvJWFFfsI/cwStK
PNqGrhLxe4A71NWX77fPBDsOycB8D+di450qqF0sjgztYBcflB5v/3yNfAwA2cOA
vuz+RZ0ouUS4dAcx2P7nGOK+v0XjgTjDLw3GNpoKFa0ZIhk1jneEDIl6fshMcFvR
9SYd/mM7RlIRVGTioQ7sR8g2/F+5PGssN/H0DAadE6nFLR+ASyyfzRI9Xv8//DfW
Bp+XYsuuoXmOej5egH9zDjCPi6BJx3eNjqyHOb+LWNn8AO2JD1WBVzXy38laEMtU
BP9aABSrWVBv6zWOF2Gz/BgkyY34KbttRnTPKHjp3R9TtiRF6pn5IbCgCZIlSIQh
7HdhdJQ4r7d7emDImVi2F34dXfEtA5ko7Or8bDedGApwZaPWYJA0tsG1gnuX8k2J
5zcNbF+3Is0VBPd18a2qHiNXrER3DRCFIl6jimOD9VfERyyujU8KYF0WZSTWC5g0
jTAKtTEYvyjCaLKTmSlPfugG2prLTQ7ge+AluHFwL4BLy7Eyf5E2xugEpEf9fRb0
D7AGfKa9dJ4RJkvn/UMvoRNbKeRZchatSgJX8qDEafgG2DhjdVBZlrVdoJ5ioTAV
19U0gMnldDroASFJc7EeeVn8ZA+rBdx6Syp3+HX9VRh1z3iTRwee7iQs7xRX0iDY
GdjhJsRDunxtZOKT0YB8UBsxBSNKI2vd2HixFvQ+nqDzkIVxDrCUe4nuww9TbIPK
sWIstjMJHcvBfO4nn11vzXDRVhNUyXalj7/LZpBK6TtYJ20e1iaKuwYnPW8LTC3x
UpnYW6gaVggvqZMrP0KAwGXcq1cBulTE0W8sIsbkTRa/GTTltlyutbjo5bFgyaRx
Uy/ZvLPL5NRdKEMgj/UTjagCfZbF6SEj4Y0E4QXS/JrQrFSuPKZd9ByC/4dnbGFV
oc/KPCS7KCA6ULFw3VaMGTCzI80WT/YP+Ef1ZGOpn+ZwiSpjH0cGf2LNIFJ7ZbO3
vPTB8DJa9kgC7txKLNEKzAQIk/Dhm5X9E8UpJl3e7fYWRs2nEwy3rYedR8A7bNKF
kvhdEvMrX8/PLXnSwo4Ic2Lbf5iSYi3z+HKZqq9Ie2i+h3LKC33AngJNfx1hb/Lv
eOdr8D7LN954SGR3/fom7dG9fExq+8B7REXa9mmtK5U3xHSp56WgKeEE7X9yN2j1
LApJKfKH20MrW3bpqyvcMnm3+Rb44ddLiavxYo08ESELmwcOKfftUKoxVAfgG1CM
A9ZF8rUKs/XYA2IVu9hIlUJbxwBZ3TYMTzHYhoOxaxmdva00g1cNPmkJJEdG6F1c
VSGBSvIIDMb5nwLKw9zmMYpRXRA294bG1/YhBQTP55ZZ8f+KEKMSQy8HN1Jaq6FY
qv4dyr55XI+7346FbK5eCJ42LdwL16YMPONeKj++CQXXieNGBiv0uppCGeBuXXSN
tS8/Sx53uOE9qhBr5wHLVe0CIw4+o+slT63hiXbsrpFiJVd4bhHUQICdYCm0oS+/
QPYcTGFTZRWIYsSBVdvaWD2DkB5QOjcN3rB+sN9yH5z+O0ITsc/U4kuFHwcdAumv
9v8o4VPtFmkWnklZP3cdwEtDXTAyQn3f+u6hrW+obKsb6RwTqWVr0tIdFaOgQcHS
xtCWpc7w0aT0UBScjmjkaoMWHZX5friNyb/K8wdCP16rga96v9hOvN0wX/soFefg
E3120fUFxp6Lkokcp/n9XwZTcCzaByF2DPkZXjYvttd4bIWGt7XoqbtjGPswowlj
+J1CZ0QckMFU3vuVEilcQ58g0HXRTVnhv1gsBpiSivdOx1djlFNHz9LfGyuxMorc
1ZKVXNfdRRJeAqEd0Z4YUWoGcYWnGwkkzjn2yITRSnDlT5snIC/v74gYQt6fT+I6
ab/BtKzwyUpJiLUOXM3D3JV9JpMSNJHkvk7cRao0T4Zo7ehiijL0XBXEhZh/Mnf0
nNkS4pSY/Ml2imDlaJHvf3hmqYnAwBcEkOQ+FtkgEIAphfhpvSs9mcpoHjgaQnZo
1eNcyHDOVVTQ/6dD5lQgfkdZChrBjoYFM38jQMTo3/GCyE5aty38LIc8NFEAPmZD
BEpIoq0ZZ6RgkMa8KPmzfN3yPviToE0krOAhFIdujAj9WgL0MZN12m/Pi3uo6xne
R8gdMuoVFyXvzZQVL1Z211aEiXbBDhl1D7ai3NsveZUskS7QxDVVwcYe+mUDpLZK
HONbSvraHsyiiR5+I+00pB/vDBSW+LMKQhj0CTKpWvMf8OUnTGqIubDQPBlJVDSx
4d1qJm9Oi+GagoboW3dn6Kgrln2ZFDBywaEoZiRvSOO9CFdBsdnPc9V2+U8LD3CY
IMQK8bUOl+k79yLKAFltR6Y6kZ6FX5k7k/VJJgaj7IS31mOUTkiLLST5nqHg6Y+j
lnIhNLBrsX5FjH+xokjnp2HN+VetnGqRFMUaPdCHjxKZETKscHJkZM2jKM+TcLqw
NvXIcyDYuE8F/F/btO4Ph3hW8QkYFfRWOhf9hZJ0b9VaXYwOH/qgOeQFGk3dCgio
NQwJPka8oLag3+/mgle66oAUWVr3PqvtBF+qdRhFAqhiJTln57SgjNiPSndYT8gr
sVov2oBHfBfLHNVr1sWZ/XTC9LYWy9Kvg7VVzpb7Q+1znEiKSMvMWXSaBC+6ZfIH
3AMMCF2VoEneqv3dvmX4fUUYkOpdn+4EE6WN5DBugmWJMk3ckrYrX48dYk+okPf4
4QuQYgdwzznfvqbKllIFtvm8KBe1SitPnqTRjIiJ1KtNkEC4zrVKSSAfIQdLqsS7
DZkwCCuLfx+as9sA6+UF8GX25MCik+oA3GW+Ds9RVKSpXg6dAeTpfYbozm1LnCFR
2WyiFzUKbfJLc7ioH/gwXsE7CmemndpsiItN7NmGdgtHO4JucTtr4VRME/B3Qy0r
yODmRNY91dzN9nhhOzncj9tiltTnh57x2VcWHcj5+zVqJsFy0HSsvS89PwWbY30u
qShi25xNTyMMUZ5pocZadmhJoIGfywaCrhGwwS4WxvFkAPP0IasQualOC3QT7iAe
lAwokRdGgSXToQgk1IRjdEdQWowchyf4iTAx9o/0Lm7dtY2BcvWoFWFBRXH7M8d9
SWh4joHdnE6sMCrA8a9ZAwJjmNVWS9eqvezdv+E24gwahvmpJArZiuBy6pUmxCp0
ly6rVSDwnySDNb5/ob6KGQA0BRqvy3AlqqHrhccYy7DwvJOPGjcrsu+WHnM2dsfs
CJHt2OveMpewEsAjE938mOy39BNrXpOJRZ/3BBs+nBpb1+cV8lzvynX1fittmRwd
zrqzGM7wA24ec7ALEbTqioZ3EZfPfA1KDmcaDU+vnyzl5R7dU3CIVLoB33eNWgeh
CiQTD5I++lVm51bwDHxPqA8rvHcsnKRlvAQRn+40hmkTHCh6n/Sd4VVMj7lstRjj
NKssIeEAL84dkCbVb241OmBUjkM4gmoDJZ350C4WMW4KtpBQCxRdZQ5x0BxfagKO
hVXiGXK815a3jKWzA9Z++PIFeCg/pF4prm4VPyUmHDP31zCN4h66xAepJjmwhhgr
XLw10cVb2JTYoKJoCgz9PjhVqCIOkyab0AdWGTLnBFKYxoB30sANoFNnsGbouMc2
Wvp7/1zl13IhGxeUEPUoSJ+VFVR9YfgPtNbCGxTyf6N6XMnk6cd98y8RhTWcuXJL
eOlWIqBaIEqRWaCNsekAti7JZcuT+D4IppXvIqi+qI6oVqBR5FKEINsYMmko7ELS
Ax0hMPP3CDRsidkNQKI+tjeWsgskKFGzK6bR4VA7HBdZHx6ohCYaY5A+RFIGYfU1
RvvqG+UuUenHNX3mRri7J5Ec5D80hJSKz9CBqY8MDJRY3d3OHwW3xikpXAXEkioU
600NiD+TrVDTefpgFNFY1GKlRbe2i833j5+zwWCNnMgrplGayoBXM+RTQS0idGd3
MblUkMmWh0b9wpC6k+ygMnWeDklm84VPXLQPFEARxRdWEU2swRDZBAZsMbEdER3a
s64hDUg+jSjO3zOfcs3ywPAyDnNVdMVzIMGQIdR8G6jlWPDfBS9LCHUOpJxK/ydV
olg7t95rPggI/rbgLjtBRI3mm3ne0Qrh+ZokemEWGZtSBxOgb7oeE+nVe1pErmVF
qkDCsjZqfXCey9VwAak5NyaIeXzLQP+hEdWf4WfXlYAsbgUYjOGzLTu2UMX87HH/
c/y9J7An1TNWYvRY1OYa0lh4L5hXKkP8JQmrrz/pd9U6EqHZnq5k8TWDU153QyAc
/5z3H0oNbbnQzClxz6cQtOS6p4UJtpHfokzGpv525Y7Zfb3fl0TvGKGX0JnLfVBF
/w6TOYSVcAVMo/HJvU/ceohMMYjhJc34A1CZf9ek881LbGQZd/vvFwuIeaW3j1or
VC52Qjkt4A9LzIPq+o4Zg/r3rzRF3+4JoCSDHfq7QkWIkj5wYnwi7iqvQ9zc/mlM
+4stUiCCAnbN2gKikh+GghIZ1s5IcQ60vlYY1DeS6/MQ8TX2W1wMKK7iN4VLabpe
Q7Jma50QZ4OaAZTS8dj1yFBwb0GakDGV/uwVm4ZkQQtt79uVz4hRW5KuW6wZQXFs
F9WqDmmTFtwPLlIohmgPZyRCICQUpqFhInAAnV+NbKnXgWys3yXXuwm6eHTWgaLu
V42wJ0vvl36g5VknU8kDK0vVele/3M15gSxWz5JsPIU/74/WTzJ6UdTkfJ/B95bw
HPr+8VcItbjiW5xpK4wD82xnX0n+gu3wSyiIhdr6X2GyMNaZ+KKjyzY/GOyLYsGK
K9MqFQu3RBU1G8DqOhf0s0l4T2kj7PH9oREFZwgCUC1RdBwiXKnGvkmsOwk7pign
7ridZtzWWcwqMX7D2XXEhh+6A/yxZnOUJ+1yI0gpQFaO5pK0jFqKwuiJHf5lagj9
AEX49mdw+nsBJ4F3RnfM7BQqpnLaVXIqXhWDlKlCQ6CRblmvSxV6xS8OfflXneTG
SbZGAYthuYvWIP3CjGEsWo1Z7TJk6f1Im5QMkW1hjdNw0mW5W44oBNGGicLULx3Z
IUA3Rt/0vc/yuNv69JxwaWXMqQbMWRn+zWskA3dHc3VlwU8KozMCIhvkIcBqQpPl
TYNPuoMKca4QAK6uqmY/EmN1XsWVoB0qOK7K9MHj0sKzPLya1pOS3sRALVwvAHVn
m6BcTdG9w0Gceb3b4nIraDxHkto4bN7i883VIeDWfQL1JR7dmf1U8WJr1F6bXzM9
AIiUhW1Sxup2qook7bZqg/0C2RdNTNnO8DLp3IN0AGszzlSstgintNZeKbSZPWLj
IMPr0FGauWs1G/VhMkDvgwwzESiP++GSKNtoBtID/6cRe7kkdR4ZM8IWZlyu8ifW
rBXRJ6uAfpa8Ilq9ZDlWUUxvQjcAAi8eI7aFRTxplxy/CTTDcbYnhRa4ktZx3fBy
vvqj6XL8gc8iRiz23+P7xWewIFSeJNZk0GTqaYLxEpeqw+8bd6DqtUnkg3grYZXM
dTQwSEUMO1LfQdS/11Hb3Wkr18OP1zQvomuuJl51A/pM02F/o6fKtBU0IBy9ZQBi
tdGKMvrhifYRp47OqR82beQaKn/G2/A0AlLZs7ozOImWJ0dd8r3sWigv6YF0V863
g7mqUxnIhumsGXZ81QBgQfzgciUmzJ5KxJuhm9ODExu8gAOZHG93bbkAQv4RwWu7
N2hWq+LjtA2C9mbQfOA18yTnx1siNh2XthslSZBocBUYGGv7gTLQ/ZcJ3jBvZOz0
oiyvynA6zwJiG8up9kMcdbWGjoRWpDH9ami+H2x/NhSL/cG2qmu0pNj9/Xewaio2
aa0Igg2rTPK3YwmFgAldk/RgVqLsn3FBnqxhDx86yzoO8u7inpldVC+BrEy8Mvxc
x04TiTui9tdwfrpFBePRzpUKJrkfP6DILkxLed3LgLLVAIYOzQEZZm823KFe2akZ
NSVb3PzcdjBSM0ODLPsWy07PQ1up9ClWRkT3urrReldxYxHEKAjsZbzID30Xo1Xx
uX75yYECR4VfflBeHg273+i1RdBtwtDH6lcYMO6AXkE/HTn42zbp9I0L2axAhbf3
nTwgcTwwX/540HwGIuWTMgjwkIwHj0YzsLzxPHKCxZdQA/taWmCqzkD7XnKXDi4v
n5XSq0OMdaMPciFTlrwHK0lTGN8lSZ7wSlypd5Pinq218I3yAXT92Om7EWfWoP14
zE2fbt/9eQ9jub4ty2wRd28TTKqb0pgs2YZAYDm6v8pn0BAvVOTApnvUt9pB3est
nXYbtABgv2DY+sybpOO8CD/+HQBJj27U9zQVp7mH/7PRe+1P6Z4HtX+vuXCNCsKr
nny7iPJdvaOpdmrAacHX4gXTXVGgfocRqgQ1IiKEe50L1Sqag5SEdlxpHwTCkWmY
Mks9bPr+O5vmyoSYz/kPG8/Kn6U/Uv2xrpsbk2CKXjJcMUAOFLXBAUkpH4J0dQbV
i73VRdGapvJQWFFN+zzvyzxwagYuTjdYoI23bJAxmk8F5SxCq/eAoGyGvNUZzrzO
U6x/s11eCda4dD/QBLCDoJemVzIK3sKDyiJH4JIJYIx6ui4i5SVSsDNOcoUN/evy
pcccYL7J+WwrH8Yat/rtpba+iwWDqpPBotYZqdyRq/ygZJzLTpI+tWmnWwnnvqQ3
b0sdVMRHTD2WTC42watILjmqCwvD4PJlkouY0xL6B9Py3u/9L+fCQEMbnR11X1oc
HviAQgAOBNIXlKkeXZ/5e46AtPXfcFGrilOcripsAjJEWsiEJjd9UdwF8+WrtMtL
NSWCJjfU1M1Ko5Ou8u1H5CZDgd0ff1v4uQleYV8wRGPIub6AYCibmcK3OJ7SE2W+
rkBtmC753qRHuE26MYuwIgvSx+P8wWdReWkAfe2jWQyseAP/1QS2Xj0XpVCcczTm
9UXPxPPhSemJ2JQCuw9ol9JyNxfAiy3wCbn6V/lpAr4U0SrbJcL5rZw98gns6xm/
zHjP0K7n8ldL/7IAO7YWhoMp+eXR0+MAeBJSt6FBGqQmNShWQ12sd1QgwlxoNlSo
GZjYvMsF3OkRDyyTlnhq4VlK2ccMZXdVd5SZMdx/Mc6BUWrWivNND2KPll7fxBGE
DiyERS2CMVxBI+JNhhclcJL1avc/+kCI0RU2f0j/mRHKw7Mbi5fk7+Fkq+3Dv4bI
6V1oZn9q0gjUl2/3HTz16FQA9N0ljcI3Scm/vL8aFYY1TILTUbeml746J7Fp16QD
+P1wn5dEb4NLKWRFH6PAU59Hc1CFK9Nj84l6wWVoXTHePwBgWSKZSepenGlhK+5b
h/CiEwc4kjk40+9kNdNG8eeiiirRu/LctA9C94R0jlvfEDWtrt8OwvGHP9D1GDQl
DnzKa94JUk8Hf59inQkEyGTggya48FolFtifwvd4UEPzOLBLMp144SAaJ8RhFsfW
eGzhM9vHQDubYOmpDFJ1/1QSXuwRJn+f8L0UoCoy8cEDHvblMQtqXnNDC3qebJ4i
s0J8+Y9SqZMOcEqdsPqY07Kxyp8/MYnAkZXL6447O0mAsCF1G6cGWHiNQ/ADKcxH
3z81/Q3ZcO4v6+wyT/giOCHK65lya/WwWvaxOPDSj0UVluE/OjtIEeJmSKLvu8nr
OsMF/tai5Pv2NG9CudGPjGIPfWiOavoLjvOVNEfSiXswQRJnl3eudWqBrcSwERyW
1e7giwf3ctEtvp1mbTMew4TrANxTUyZY4crHqSgs/ifhuBTnybdRGhnqHx3V5KyL
PJlOy9EY7Q5Gx5JSjRLNY8FMMy64SRttn8n1oawQ2Y6cgWZKi1sFJdpzfLhfuFMG
DqybfYGUEhMclPD9p2OfwCBVk5k9BgU6VcGi5DjswuYFas5rhEnOUFfHlz3lbvfg
fyeqXnXL67+d7aQTBSK4O2tRrN86M+A79LdYxdD5kclKJCUYt/13IFxOIz4+g1ns
zsrGD5sL9zOLELiM1tgGndwl7jDvpvAE8wssz3UU0ZInAYMQYooa/kW2y67KR90K
AGDet0MAwNRDcld7flO44esrpo0M/TzVeUHQlmrHwj9wrCjO8nl/2vZoAZyBGVuo
NrCE1w4sYEJW2C1+IIfosyT7UumzSX8f3lD0oObluRnFGTHD7v7R1AmXVQ7opkgk
RkTO6m90OQx5t7k1TYKVIrmNwHe44aVO78b+lEU2ynJ4+GixClmabXaWU0riT4Mo
dls1wLoVbF2SIwEG3JQ7mL4CEnk4HfA7ISsjjE1SAkWu7yYAzuVE99v5gL2MJsfB
xIs7Pr91yuE7hjGu8h8AJEGiuo8vBTfu1EcIYmWE5RX9JQ2IAr1Y6y+7Byd5k862
Yy8MqDsF/lGSblCOKUnbFUFcxAhNvRa1qJA9sifvZBhEiOC54GxD0k6TOT0KeznJ
7Aa8p8hwhou682EvGhfisHT6IhvvgKmFaC9Rpia5pXyzsK1PCxc7EfVajVcL+7HE
03TBVhZpyqc+mYqvq70EDfXwnfBPTfR1OYMup+wKYM8vCCe60Mz+XfjGwObP8E2B
pSowU8UbIuHomxRcEspxZbar1sIURG9ZmhSAt9A0XGgg7S3mtL923E25BynE7AUS
nyJ4rwFv+5pK3nErxoBrJrutYN1tlUIagwrOCMifQJXb0oyig7JamMhdjd6awthy
ZlWvoUT3VF3qaON313mObf6KeUX0nDsJ0lGLjoUWiqQiNDS4lb1EQfDmTwFwJgm8
hUU2VtQqzZouj3kjQDaaqv84uKkJPHcpZIsqFyDMn71WmTdoJjQc/CaK/BIKYvsY
ASfCIPyC240dLAjPMpzZ8CTuxSq0dN1tpfha4ZY+gKIH/UuhhaxfVqW0v7hRUNHM
8W/srfv6OOEjOMulzer90jIKqBMsE228ZLYRh3FcnrvAxI/XPebac6JJd6RKrhyE
swKiD+yrYzMlWFHX3bCVX5m9m1YX9DA6uqlQwvtORyRmZ41BYcqZVtasQGE1ZoNd
lPC+SI3NLkr+6GThcKxq6KC7GLGEJ4DakCR9NNl+y9FFeynO0uQUX1OqmE5gD7Wa
H87mrJ9Kpu7zE2Fw59j6+n9W+8FmkaVMQ6sdIqISNuXY1ajo9ugDTpc538TbdpoP
IrEuFCaWJ13pcOR03DaoUogT2NyJSt9oMOa6NB2ZAw1vvTcEhnqGlsGzgfyBRh6c
2E7T3AM9knUfg9ILVbZWwfPrvkUpaLxNpGh420yYYCZqnRO/gy8g5XbSKb+YrtIz
/kSUpjBX1L0p4X1iMpcFfaTBrg6lcU/HgEeFZlFC1HxhA04ipwkl0yPAZR41HSC3
0sc/Vjj1/0h/m9WfeL17sQU3AbJJe+ENxuc1wVSJZlkHY6Hs3p7IWYZKsMXQT7ef
lEKIPgfoIDTJfsz203JOqKKWnibz8itLE47BvnAe2jjLg9BQLtec0nJe+J006Dxr
iCHok9flItRSp4CYDWvd5rXvcw0SRZ9Y5FNtdFOuPh4OJJ9dBXqdUIpq8wLj0L+Y
azKgC+/ClJ7QsLKlJZZeoSwVYtZLuOSBmoQHVFR8mHCx/LLoJuRzhbdZvAA8ww5e
EHZgvIVwiP5jEP8wqxvdwnHfSp7I7Ek/KZkGTQI1Y7kqhNhMDM138Djy38U8rOkf
s+6LFssieNgggw3ZNZlo5GpCz7F6RiEQ9DIlWFoYq1MYGzVsEprgWC9NOMNjHO4D
70+vVrfNLXxUVia6G7cEQzy9ryZlQtmXRCvTxpxp7HB0xKB1esBaJXAx7PAKDY7R
Dxx3TSv7ciyQvtYJziJqY0KPe6zftlZpMgza0TP6KqpKanARHkVtR/z9TIhya/FH
P+Rm2pe2OfuaMUGT1eubnYl5C7Z+0RasPRst0PigCM1fGhebQJnPb4bVjJC+A6bC
sVU0+xP0imWrUnNFrHJz/jSNaMuvGt9RtxTSjRAYH9up3ON+XKUJDkJ6kOPZxAay
Rx5M5ppcs5uxUkH+NKqLXDFshEY0elDS52yYV3Tcl3Y43Fck7myqZjdQkeuAv64D
0RIb+/tlrJpuIRJOSOMSe8lnUTIzVEJ3tVurTeWEl1iyYYRgk12ocE6LNYMaEb7X
RCXNIwnSxBsHOZk8gPg3Tr5hx8KLg5mr615/rgMXZxKOubmlYQAPKnAjeiqMbk4O
a3Y6z6Hgxs52qFqKwfLUKe9P3rWszqyQTgZTYkx73ftZ4cNS9CH+/wPgdhO1kJHQ
bueTGoUrfLk4gkOu2SF8LE6hu6zsoEh8I4mar9mPPg9yIp2m8OtCpZl+23GragjQ
5XxAkdDRImU/kfFDeom7BzwdRRg0/dHd6/xmwVo76+DYDBJpwzb2QgmvtlRQb7/q
tEymZ6gpdvz0pXfUiBokCKQzYR98Y3bjz4L7jR9xsMX9uKpmPXweXKRBzHoTnRL+
ii56cDdWnYTeuCFbab13PN2OnqRwCLNIbuAYnEgrhRs3ZgwlqwdHqK+rVZ9IVvxb
TatU4G2P+sJ3aXdpTXtyKYsj2QZph8wym/kVE8wNbJC7RXKSR6bWA8ZJzI4AUeer
VcwFafZuWGvHAlsyY3/XrNhtSO8VrgdvYu2Tn3tZoPmPgbcWE8U8GOxy0JT8quQW
MAbN2TQEHULnPg2hFHQYbImw8AqVqYAeEpSRWJw1gBPm6Wvu83mhc00IVX7OBitI
F0m4uexjNuFPPMWTPp1Ub57gZcpSUTbpRBAGY75MB3lGTjyL8MbKVIFbONOHaSNV
M9k8C1o78pULMsKrkKGp+3g6OPKb780n6GcuDHyNxaBAl7grcv29qkZk83Gcu7wi
qxIq6+JuXB/OnVm2oRL4PPxBnKd8cTustWkzdJ8bgNj+3HmI3TzJZikDC7XHRXqK
Z1/Hd2ggGorLpiON9Jrn66DxRLJgEIuET0GclWy99LWqOS1qiNqRezmeDUqb109V
wpq4ds6vzyElmwgDnjfDYgrB6FsMl3Pq9+Qs1B01KaL9v3c7vwHMsfh7smJ2r6Ia
qWuMqXQGdEVCTsfOPPXwEFRthDz96AjOQ3Ap7qDsjlYntYvUDTZJUzA0ILf3yA8f
HpPoQfx1M9+5y/HTzKJfPzWQoQkm7/rSxQibyRJ7007YfF7mM7O/4VGgOzNDb4Pl
oWM8N3XP2RE94xTHsiBtZrFGSMnbh+GMHCl8Cv3ys2UoU57t5LviakxTKXvN1tea
lXf1PT8Svd7wMBcbCPISvoyydIevI3mfuG/q6PU6FKCoPMI/LYgSJuS+zmJxWM8Y
QGcxBUkYdixmlOyARtFWpVmh+Cnfahkj7Tq/NNQeFNu9BkgAFbCp1iuRUmdDVUKO
cjBNgZT7SHTk5VSC9w1h1FqFBRPXfbx10rUv2xvYWKACYJY+xUb8TuVDs9I/Xgz8
tyVQCuDq3g11snxPMJNXCd0NyRYAbgMvzad/lV6bkFbR51LhDuVMUj0JXXdnLF2v
UdJSlASk2KWeCWAIQabKSyHqATXkT//LFrLKVnakV6kXX2+O7/jrL2vECYJp8k/r
taz2H1WeqcYjnQ6VgKIaU56gSPnodxkxqCRuP9Jq1KY/Q8iAXmrlN7wYQwXUOovx
U0cDctP0C6mURsEQ3CK2W6e+fWRn89t2kiTxBM45HfmEfjW+Om8Rk3v82j2l5esO
fpyY7vWv8n0hd/8hfVmYml+i3alGO4jgrHHA66i1TCqNeOQXbTbazrvxnG+ur9eh
q1em1LY3BIeozu/h/vRG9qcyBjgvepVAVuLmWHMmSG2oq8nRWuHmQ7yWhlzgwmHZ
bcUXHglSPDqFSdJZ6cweFb9HYPo4vrP3BOER9Hsq98uYO5wNyn4qO0lbea+cbAaT
iRgM4BYFbGO8SZAComZi8dseAnJn1x8Hyk/GF3wekIkpaSQWCxpwfN+GraP8oI41
naR4srEplZTnHrpgOWN8vEuHVEG1x0Kr8zjMI9iOmhuDpwGe9ZyqkCB0gO1HelDB
hhrJgSK/VO9+TYA6ORnPCS8V9yAvF9w6M64F3CUROveBNj+LjgKh08/xUvgeW2Lq
iqZdvTKBIrwR80s4EFb1BDcKCZKUBe9Nj5CcJRxQGvwMB5wLnenuCyOPyYFwOm8V
s2xYa94yx3SEQqbMuuvyQDCflY8RnGHufRfTl4XM4GAL2IsU8KhLMbSwqobi8NiK
gFXFKjxLAQIH5wqlqnG8O2SFJhBCyidnne5FLqfYUxj1nGWtu1WpKlRZW4DNpOht
ZHOMUkykSv+mbLKSh+JqNCwj3hFNKYk5toed5+5H5DOeTZwrpVOWOVIEB2pKIud1
alnTgCOQNjwXEXxGrgiQSTiPX1K9MUDqeE49BVplCR3SlzdIqP5pIV1OLL0EKFJl
k+KzGmI4Kk9OPkmJIFkdBIaIkrrm4HwX34dBJ3nO7pjn+nktNDAP0Th1z+GTh2QE
uCOBWZcoZ5upjVDCy3nr5lZg6X2Wqfr3j7Bh8PT7lAax2+aKNvtodubEzuH61cZ5
nhLgdFq6Vx39NlKMnLnjU906KRPd0C6uUE84oRST1/351aCYmg6MeLhTLGPVcJTP
/yOFlc8WmywKixjGraZxI3tf/Ky7qOxcIiMWtd3udKRGdkPtyFg3JPsziy77waGL
mDFsIJ/V1ZjyKZik4KOq8kK+fWowhBR15bfqLhH7aaJNUWzbqX90To9eP2PdjEX2
vFPEvj/OGNlju+ViAmrcZMqSPRDlYcht74zj8tzwgrrUCwfpAir1JEZFCE98TZ6Q
XD2BT9SMvb+4sQLn7PYOv3tyAWpS03+CHZ5iFO/+upULTaCTatTfTImhXprXHf2c
rI8vCY1kJasG1IRlJvf4afAtPJxrRFqf/E/CDqlCTszgGcx6xdHOKnglbMIiULwk
Br2TIPhtMExHNDR0f7CIdPdoBAePBL6sf29bhips0F0YB9Im6JM6hlS/+4a3xqeH
MOlpkYTfmESgBV4RthVeYLaZcihw+u0qXrg00mdE3kdYreYjHtTY1lxAkxozbi2W
r+PW2/xZ1zRUhj/ghDdOcqKL4dEcv6KHePzExrXt30E0x0aZoSM6W/47FFguwoRQ
u0d6I7f8vHCEwZcP/Upl87U6iVmF5mMTq5u53E3E2KnQ0Mto+mTX0+MteRveZHnZ
JlzIX7I9PKJsqkZKUlyy364nIyU4K6f7MvG+yLv3TeBzSauhXkcLuK9A1iSQE0Av
GwwPQ9GpTvP8PDZq2OW+067gZytX1Npx7gyn0lpkaanvvCJt9Vyrwh1pUB10lSA9
Q4/zoqzorIgNA+VoBgnA2F1TCoBRm/WhUsTJ05KUNULkW/cAcgDFp3Ad0d9E8WJ9
YCdhXOyZuP0DI1NOhQG9jKKvntBsL43EfZ+2pTIqeF0/s4b+eujNnhUsPLfytmaD
P4qpvjuDZG8R9382OGokgv0eor4BbpHVUd0e0Q8AAXivw7IcFwJ9SRgrs84/fYcJ
8oZYgkoghOP2lbN+HrQy49bKFNv5TIjXrvBhu68TTbpFN/Zax6Voo8xvezZwlbfB
kI9x6FF9+4F/XAyLO7wF3+ya9vWgqQKF3DAPJjqH5qNaSZzcaCm3ufs8RZsTe9sR
5kXXusoHm0xJuJJodXNF4SBf3SsaU2vpdu73IMA3Yvno+wEDyzN34iFoke8tEEG9
OwZytKkY75RokKdVgQcZuzhIBoiZtDI8yhRcdJbBecDCKgbfpAdMp+9oPk+kVN4D
RL/B0qjcaGnKcUk7SEEYVoJcKCZ5/yRNC86qcOhQI9c+iWrOSJH1xwLsp7XsmkQy
rhGn6+7ZKDGG4TnjgCuZBAY07TBeiVX3hhyt17Tt7iwrinHf/GVLI1F5YtTh2FLK
VPWFC37BYv5r/TgZ124KqQ3HSq4YxtZEfoUsUPIqW0PRgPaCsexsexiRSCVaT1tq
VjcUrATeVvP6NTYRAL9OlXKyR3g1uPEvldG6Hjrn1OuJ5sPE/D4zAy3HwVEqOsxW
9ebvE9RUSSRc1p9675PpfVBQDwDPPzu1WQGsE3NZ2nlXuxG+Uma20w/LPtBiMSyD
YMZHcI2MGHV8wHf2Q7RxRB4JrFpysKeFGkofqWOfFfjqrXVNKP5Jta1p+8OIg2ms
lP/vMgbrNz5gM2I6mgp0j+6ATTX26LUCJX1i5xpAxTe0LgXuyxmj6UV+JWYVIzch
4oNcChnhRUAOtzY5dB5S9D89x2CgIsAnR4PYyf1mXMGGAWuZnf7eH+nLHz6P0yCA
x6sZ1mekZXZvKtyz+2JWmJSzH2c9NOe+W/8ch1fTA02s5K2pKsI8REZduDd0kWR0
rI2XcUtB98XAM5+BmVmWHI4CBVGctMDLTT4gU9Nd9Kb1M2A4PIq7soK3IigqWZuD
LLPOUGythaIHyp/yIB2SDlG6CitAkQzOeX0jELKNTdQCSRAEeJ9Q9/K7jhniWglD
efbHRUmBDsgy6T177B2KoEFEXCfjzn0/wneLfy4vixpUc7Ohm4CHXS2FpXFYluv5
/LMaddLlP+4W8e820911pskEurSRYrtJEfPeCoX1XA/QnHydi/xOGKPP0QRGjFTC
op/ANONnxZY5XcSZjfKclPcMkdbydSQeW8IXLgaIf1k2OEEo49VUWCHZN1swNi9i
vHOYE/4+4vMdVl5MvArO+SK/9kKtTHbtPJZm3mK5HIiDtnw90v6QokMQYIjV9dGQ
GIvQg8oJfvz5f9RlzZMArg8QHm7uZnF0oUvENI141G+myuuPC8GjTThVD9HjyeW4
EOdnrVUgF1mR+o7VQxrFhap+U6XdlRO2XPtgvVhWmOIcsXDIIrvZ/UaKAdeLC3kq
4l1ZEGn6tTCWbdkuGDh2u+OHWyd3glNVVnkOIQKWMjn64tFWeg8O++tW2slRHAsI
K7vsyoTDjOa5qM37k2CH3G7mZUMyHSPsFhonJxQXFfQnThlN69xrs2pxLvP3hzz0
BbRsfMzG40+7o0b5JInXy8vS2yDURcS0fXJNRv9nM3x8MXhL5lePr0HuC4xi4Y71
nO49/Op7BuWwgE6v43XemWJViJpnNN3JefTpTIxIPOwnqZLsqiTlVMSghAoQgVgX
nIwQzjzq/0BC13lgnVXI4p+vBXSa2gmbYk1UO3vFYddYcT+3ptX5wnUyNS9Z3FUU
XdZpHy80oCLk5a7mkNC1uhij9HzB5KrsIWBH9+tleGH5Cv9Q0JfOTevwVTTnym7l
aEOockZDCQYffaltU8TQLNbZ93ZIU9Gv/c9joogfM8U2hUdZ1kJ/IYCaVvLfTCO8
5EqRu1vMN4LGG3GJ97/aiSAyUGqdau8jt030C4xCbew9iFIebmaSzObfmJD5mIph
Yw/O+VNUrgG6hLJcPwlofpOw5+QLIMZ/SRHOn+xbYFyUhm832JRlKMWjwF3muWdd
hOnYZzTDc8Uxj3LlctdBquHIxgig3Fm2/ZoClVgkJIXHm/Z2k3Qa2oIWZKyb9qVU
Q/LmEyBfH9Yj4v+T/rDxDQBDgpNOyx3XryPiPFFSj7wcfOFzbEvZoRnTlM4QiXE0
0E7LhZbHGqjDpN8EPgdAHhMaQk7/G4CreTWGnpunGwPMUDP5fHH5093l7gV07XyN
Lx6/xMO59RPOYJLmwC5aDsIpye9yBmr1m/hw8F8lTN5+FZzwlRCZp3Aw753Y1mRs
yxyOw7rBPIRYa7c91h7UngpUlRPTe7i4qxd4TAcI1V/Ja99BoxlDGj/TtBB5SoF0
XRQoMWfb42/ou/PptZG2/UDZD/OKCVuhrWEcfGGd9u0xGXH0S8WBVN0D3n/yvXmv
tQmRFmwPY3ZbdliplPVVN/ko1HK0YsxtE7whsmxeF44WaF8ZY2BP6tj6sx+SFiAn
SUfctcjmH/RL245WQ5DLILH4QvdyvCojGLiDnXQ5U4FkzLtgueS5lnH7YgAk1u+0
6mBLKfmp40f8BzUIua0Bj2DzjuxSkG7NnEykQgibdQZSv/NdbCOmt978sdNiVckZ
Fp6huV9EIk5+e3aYml5wJEVbnx4RQ4CAvb+ddSv2Fn4HlT+XXZhyqAU3m0JTsoTV
n86YiAvun5BE0qgVjTEJ4CFHtKQ/yO3wcl+vJvthLfliPKXwqOqAcH1ZGiruZ/tF
QZ4cgcBsm6lf47QA2y/0j/8Z5aCVz+nBtpuzsUgOArywAQQskDWtUIjLXhHIWuGd
srNt42qm/gYQoTCdablq2B7JDfU1jBro725Zb3bWuosR+KlMq1xrLRZZe8lBEj43
zXCxvNWnHBbEfR/rzj24iy7P8zzUIW5Q+K/TSPzujrobZReyvPmsiGJUydMm7WyJ
mcvkKyhgNXKnnm09MFi5/y5p6PgLNTcXbbB7VKZBb0VuhBcdsaRivSU/UqyU/77j
awORUJL8Slcnn3xtB//zrh04X73mHw8I4vsL0n9HuFe5x/njlTeEZIX1I6Q9efIV
1ogWjmoaQ3+c9CZh3JRruqHamvr6usHq+wqttIDkbl0WllfB+Ovd/x9kktGFyUTK
WzvnsNKZNdFa3IK9OLtakUmPXeqXG2NDki1meVRuD8doANqOgBiv354xYMMJtCVx
gc4Ldlgrvfjmwi008WBr88a56omxl4OAwuBJQP1Kax8hcE2esystAC0/p+uIxfYg
lopytquW7sLck3J/TwXn3qWilCEbZfirxP4EcAYceZBHNCvWP8olCQPKyX7zhqpp
PkYmNxURrCfGamZVWR60pFVIvKAdxnnRBooTLuEA4s25xGATvBn5O3Gp7wFNkwrB
Gcf637zFUJWF//yBZt1TbRjOWKDmchqJTQVqglhelqobaCi9MKGieQGvtuiWGx9D
uwhONJZLvRuRtjY4Q54QctyivpbUhpYuR5EGlLAoM3Vw5eIz6c/X5PhylSl//EdN
HgG0O4/mhn/l+ezjxGGNFeqzHl81KFvfI22n9GFnfsGE6lepfZbppeYIvSFPPv5T
MviRyNv0E4I4Dm8MwyOhNRmLLkjhB7anwID4EEjwXGS0lSUJgGN2rQfK44uo1vCH
Wkh975NAb8ivAVOhvAntLX0CBneYYfM2NHo6n6FuUUu8PzUSwKIAj44q3UFMlk6S
LNw6E4TDvklKaz+VYYWnGyMXk2gmPA/3JaEG1RrN9SQ0qvEs2CG0sr+gPcwzYpHO
V97fkDSh7bDDVJHJjHGW+TrrNNaVxNdDaR0OX4iy84N4Gf1B1E/GRvbkvB/qoeNU
SoH9B/ek2N+A5k36TtAG3cRRkYHmSfvBKR2qeTNPpSwsLBGuwUvD0XXJ+4aKIOpu
iKKE7M4Ed0XeCSx7Kkg1TM/TKk+DcXUDzhnHRSwRxVZ1MqPHtoL1cxH86zbuorJf
Fru7pYw1Og6n7FwC02V3guu41m469rWeZ8piH9BoZ7ToKIn5hWlzl3rU5wb5+jcI
rd9y+vpTMJENhZWYL516+d66Rw7aWxRMv7qhoYXf6UGrOZ5q01qetvngUpL3Fb+b
pqzNi5q/X51gWfF7qQv4qDa6ns2c9pgkqCs725Opi7k5XMwWqLCu5IbtSFcwD2hs
+0Xoi7LWObZyvcNyuDAQVfMJGz7QkQReZTkJE80czFC/Bz5h1LiK3Y1k7fRImr4b
gsn0e4byz7/CFl9di4ac/vl4BXcj6xQYZsLe31Yx88W+udMxsx0jsRgW6eYuwy2P
9jyDXR875T33Ra0I9mdlWILy4wTVNPCHfvZJKiTIyrk+hcKBiJoqKIU3rdJzfKw4
FTskddxKXPx9NIkNJodPTq9BE9Ba7xygPoF9dXq/LYtg3iQ8SLwFztaqv2jnd+hw
EP/owWPB0fVIWW8iBrxMwc7uTW3NBkmWFfOzV1sKtOQZHDKSxQARZaeHW2UgajBU
FAD8mGV+b1QLeXZQUSGUWXhF4MSDXskxQHSoB7WnS4TCNy71vIma7t0ELwsrbCiM
NVJMil4UXWngu497mBVseEdTjEDlxBifBaJ5EbPzo8S7JOopFsyQ9vwSZWsXwoXY
feSmDxBu0lR8/qLJlYknCJJOKCxFRnuGxEKu4kOlhUjE08hI3D5iFASOMfS1dFc5
4yjeZkGmSGgbP19aNYY0XDE/0Ai3XALdkPVJELy6hbnv9NxoCd9NbOhwChlp2Nbg
3xo88SZh8BuY7IBmEvUSzENA810bdJSXtuRt+gQC8nT8uj6C+fuJb4M1rP5M/JIX
O2sj27iYGGRRyuye4HFjKwP8TsMfCFt4eTGP40vi8jZJZXtS87rvmiHwsxnGLgYJ
1HqWGL7lZNCacTXu2F9toCYjUHMUba86RiNf9gAK/oUfO++JT4rFpsa6O8PnyAlk
FZNHHjzbUuxDYwhnHVap2/auMM19yTc2+HAjbyHMwQ0/GnvWfLhFTDxq3Wns9DR8
tEg1E0G6w9gi1GN77nK8CfOfwfaDAz06Mv39zVpqmpEXrIr01YEGL6kOPBJgrRgP
YCUl58xcO8jDJnGykj26Cb15UBA6f6nCda4S/7eodBADtO12ktWDb3oEAoDC6yqV
MEL906UpcuqG0qBA1O9QXKZ2VUvqDAOZF2l2wXI/wxM+ABKhP1SrdfSZ5SuPk6qp
k4ZJKWh17RtYQ9XTR4CL8aC6bulDCFFchWr2/UcD9mEBjYvvlx4NA9slO7LXMOj/
cdISqd5dbkl4d4fBRmv47OO1/MiE8v08JFMUbwyQsYfM+L6to55b2iE608mNz2y/
sccji8pcjmHrU85z4YtX4+DPX/2PymCfIUeOZmdrJ9YPihzrWE0tIPrsOSXI/bO+
DyB7kPoItOLq/uP7tzMbmRb+oRRtqrLRjgqFGDedqU58f9mzXocSxASp2g21/8dh
ZTdwaF+eDkP1v4WXY6l0FcW1KmR2FravEXA43b6wYEpHYRG8s08WH2aYGWFc+2Ra
M+Wvv6hO9BD/yCkmxsmdRWCVmIUvKdinKarkZLFOrskvdP3mAmJ61Q5n4CFrIOE7
2EbZWYvyCzzTCePe9UmWk1cmfuucqjMpRrzHJfpcTMXAX4PFeWlvKLOu/E4dq8yv
zSJxef+Iz/bFOPNS38EMsYKf/5MsnYX+BIwmILb3T80y4zSnjBvxW6GVvoDA/8Kw
///1zVfLvQ9TVVfK6MYdveSHxBS61GS61EdRZ3SJ3KbGWdxUZa5uqqAQxyGCM7T2
uTQdGRd/5GOFSLowg5sJGzRhJR+5UJYAK4sSjh8Xo547B4rbndJ37kaygcgCw3+1
pHhGAzf885KA2J6aScxx/yb1lH2m2YBwy+2yRUBoDZIAjGTVP5FyWmZElOmF9Nmy
kKFUYYocOCh4pmjHAZirzCmOed2Os0Lfdd7bSHsRlBffervYJ2ZURJ+Aec/uY1xk
kJcXA8Yn6y+9g9ezhTNZ31CpLuVVb6m5MMEGPwhD+RMfgaiuGg5lcyXIyeyoGmPw
ppjPs09LHzZLYOEw4G7X8FjXvmHI7FbbqO0kQTWEVvMkQh6myBRzaoSSb8X0bG1q
+YGkJeYMUeNMkohkaN30UpSsw+TMP1AjsyhAGwQgdotNMCKaqU4+nIjpUtU+uNQ5
OgCTOcMB9fCaTMEo4btiCbyvuLAYIohdwQMs/DS11K9Xo0H1thCjaWyKFkJfMWl5
uMbrpIBhZghGZjbMjeIULb18yi6+lakpIDIGpJGLv+aml7BEH5iOFqRilmWIJx4G
8XmKwcxGCK+/wkXCTHtKK+M3Igtgk1cl05GFsKWkfj9XGzwQl++VMA0lFOhQbKA3
FY/TZi091iKzN+A61GqFjQRY17bfX775eHid9dx3qPqgZjmLT7oSgYqN63LXft2u
Jo3eV1IpUtfVJAFk7dEmVRQx6aPE2rsue5p/BpIbqaxmSLCfwu1lmt6zJeFG8rrk
wtS/3HhA7Tt+TueQRXhUaJc7pDBNVZlu1rceSDntzCpVdYVmFUKeM17AEEatXLBy
B1N6jwxpzKb3wD2Hjfkpfpr4zc3bJw9IGXanpz1l69hwXmbqfyHNCPXDcxwoooeT
bxIkoQGButLt30ehNtiAk1LouWCb57j6nqJwxKtvnARkAwAZlhAiiglWlgvXPlkk
tJA3iMwcwIjA0hgV5Spi+aCQ92DbI9raZouusMbipXE2THlZrRfVlWqbbzwTPuZq
7igTd1m4m4kz78f+H+hr4KKKUkdMPDE6A3G2MXejltWN+dI8VOSVUsZg7jC+PaGi
e6v4zvKf77SKIjXTKUkcitkfXKnNG8KbW5ZHUBwelirQIVDxLTX5xWqZywux9/2y
qy60P3mWZkjSU8K2PuwTUZAIfyALEcT7TZkkekS9xVwzSI/evINTCZY/k7zii2fa
j0/1Eto/2BYd07U5anoPW3aQ/sKsYunE3qCdt97AjPpxelKrrsP1yw1XjfJWgwLe
1ZsAVtqfsLQilhSUZwSVw5dKV0z//ftV3BgaAp3/YGQJynphOJ34VoW/FiV9Dh/5
yKz1R4DrabRb7Pvkk036HOwX5qHxHAHk6E2PdBnRcWnIiK/YH9NdWH1TtzVMvWVE
1SkNBERSE8UQ5VymfAEuUhJVG5XwEMPDSwnIKq6VOzRuo5vw+m8+OC5bamy9OENI
OKhvuzEfx/NrWTTVeBtO1xqFV6B558AuSx0PNrBTCMUY8Ab9OaMhJ3TWT4xQ7Ppl
8BG0A4f6yC5j+CoAA/AvKEHG+rgXneH32WVh1i+JEm6lppi1Sft+HTojQyHLCVnb
ZKPK5vWYHoBUbKFoKvVbH3yBZ1IOJrvZ43y7p7lrnFJb5JQd2PA/tBMe5MDYUSHM
D/UmuLcNsvBnPotGtTX+4vFu0KdNTDYVb8BcTKzmJj2iRr1Vr02OrDmQN3bXLcY2
F+CapGh2K/rqzcnMQuX1B9LxPJAoRG4Ln8OtBEyjrSzcPSBV2N4sysoT2BQ+q/E7
8MZTRlZSXBhg+NSMOZRRNUJJERMSnyKLo5pQjJ2RydGsOhKhVSdmyj0HqgX+kYTd
eOcDSJfBZH42bs0Z9gr8aUzkua0l5FhQJl0Gkbi0qhbMfLJRsqC8uyikPWGjDiW5
g+69ieocdi3ujvZavffKWF+dv1jPlYArSz+SPfvRAneTt6tJF1r3liVf3HXjqeEL
FbmyQhUEFM4nVujGbmLsnqDozvAAuu+fTPWKlHNuo8dwHnTj4kmjEmo0pjafzAd9
gwBehR9Yq9jKbTLc+Ww6EfEackYZjLnPBq6Jxetv5V/lUEcFhY//2+kt3G78S+FC
bfv5VG3rjueEliyoZhoJ1mdkiYuEk6OuRVMc1LASHvF1W1OhVAngFtPeSZy6Ygaq
Pre+q7mTqHCNuefxS14Xdt+306coX3MQYxFy0lpF9pYMoKbIQo3ahWkvz0g24ZgH
ktwCnR1/yIZIy/db4zMejcZAO4ZZdQGWljbKyvmu5rGufg6csj+5vSw6F3cXWaR8
6KOgrsr6ttTxWLOaIRuapogUHsgnLIcOnZ2f+kxV8xMakwTkwwmp/RWT3+2w//pZ
rC5zZaaqqebbiHXbxjAdDw+4IE7dZcpDKSApJcUPwO9SMnOEIU2raiT7ibqjjXji
uo1jWKQZs3R/D/jZQv2tIt6bkVfVcj/oalfWOwCH4fHe4MJ/tOqVaUsKcy8WJc4o
A6XcEK3usS/XMWLPYBscd/Wx3/q22XIlxWYH9SITAgbaAR8C7l1OGfG91k06aje1
HjwMazhmcrUjTIBnPu8z54BedBz97CDyzpxxQPxifDp80HrdNIKHH9AW/gtfMmEB
g330TuS/hvB3MgHL+diy0Sole0GbRv6HvIVZ7/SxQdjggGBVv/ZspYS5f8Q2c25A
2OxbiQk1TxBtQMdfPJ/IvlUUCk4LCOdliLDIn1rylBwYxQ4blKLze5yJTnpIowb7
I7YoskXvRvCfxIA0mHYgItbWKSDv7lYvW7VqRqRJh+i/oAqMPWZTxQtBxwUbUIjA
mRD3qtpsUb4fAX9TDhZMo1Hixm2NcUg1G7xvqhvwTIAQncoIkjmQ9Mk2PVbfQcmX
vXc4OPHJLjQI+CVDywtC3gNNknyaYnnatY7atTDunLu+3GBdxtHXVksvxWmOoEnC
GcTHupVdVV/Dh3EXYcJUn9GjUcoTdd8/AZbsM7xKmWKJL5mHiR+U4P3xfTpcF9pS
3on0q5m863hLwHJJCRcwG7G6zH+O0W6U7vMYs+Mhc3+pGicZ8ivAFN7515dkSmCg
15j2/dxLm0JaU7YLQHMEEtICnIqs5BOFd4jXwO4iDBmqv19jqZCY8AdASEVDYkKo
vg08BYzeglEoD+NKLegF6oXIkO/faefU1WH9qOS2CCeu4B4KWgdmvjtuGU1p6b15
PIfjY5WkvHblwVdNQa1JMyfgp8qcRoAyfv7qrrCtmUnRArkoL8FfLMZiw/9A1ekb
UJg8SCglxErE9cAj9QLcqz4aQnWfxDCdVK3jqhJUK1/Jvpp/N7Cvie37W7SA7Msv
Kiez0h/pWnNadVpZYOJOU81O4g2xJM0ZOub0sChVZ4VtRIErINe7VK1FGsvjqvGg
x9BskK3uPRVqWpMHLu0F+Sdo3dRoAfti3ffnD/r8ugMgoZVSKIOjfJd/crfr7PkE
ypPYtGeMP+n0PcMS7YKMP6ESBiBcIEbA37/nxxVs6VXhLZnQokHs7GQAKkFiUvSA
07kqXABdN4xtdaDtwMKVwpCktj0momFGUA/92RDuzf41TSK5Y78IE1PgKOR1ZS/Z
NQ58ZuCSgQz9g7Rd3NjvNv0h3v04kadWqmD+UHQAb8J5erbtB7TB8tsTDfIE+pze
zkr6kmhK7/GWejcoO/SOVPT2SuxJgTBr9JLi4af5ZNf7m7e6mbK5EK5XvXm8paIQ
dNVUNTSOHJVOmccbYaX2x2Qy02UEm6l68j9AEkaYwm106xnw4kvP0GazndoSlF9g
CrRT/dvQ5Ry8FHaqrR02kGgjorsAcfBm7ova1f6IkBU/xeKR/Ub8AOnfx50QOamL
MZgzsgAsqhQnIg0ubRYbeFi7e0/B7VzSy60Bhso+RnAEbOzqEr2VRoPnIh5cnbNQ
d7aTrtLYXFKY+hFbFH6A+Hrd0Hmz+KiT7EqN9QUcFr6eC7NOVoieHHAwqfbs4Abk
hBz0U4yzwy9XVlj32oK3rctSOYW86db5AyRVqI/GuuFHOXgfAKaV+Op0759+NLFy
utTBCG7idlmcBI/OLTXlK7lHxZ6X5x4J9xOGQT0vxF3GYxFR4pVgbvIBqHSD2VoO
NQR/OzbiTTaLwopc8RfrU5s+opq5IFyW7TadFmSJdaMXvuIzXQ5G+aVtNzIsgSPL
C37/p1bLKignZYAbu+3l9NXgTz013HTT3lT/xyyO7yIo4Ujetm8ul7IT4RC7SoTU
dkEAr9J/jdDYYQVdbkNyXxG+7J97WGULJLYvILKSddwKhVYPLPGLMcZzXQ4YLW7N
A58nV+T8pPyvr2HC4mxRJcpT/XgGGZ3spS4TpgiiVZtfO5ERm5eU8cEHtZoLq9aN
nDjJUGAZUw7/t+4ocfQ0XXmbCd0HyVI5jic/icjgt1YE1iyE4o08m1kgEznRIlqc
mNnYiInVq334YxCdNowzXTUjztDIjb6vysi5ciePsnq5COUdkH/71H1nRLeKlv+U
puWXFnFm2wOJx+ESEp5GyxYxLcwltsczugDThIIMe0fX2J3wB6mxaWM74jocZHRK
wQs1oZxIbUG/03GyO/YdsAUvtnYhu8nSrhZvfd0DV8EKTX9dOI3WAiB/hiKqY/mV
NJO4zSPC0ykzqenkl8i+n3OnQQBDpINapmzF90M4veK0ZeWWQnyTvWCSnEDSIrv1
+NCYfaZFdVvVs7e1Dr9qPFYlAalGKfFjtoco85x2gfGke7EX905j5o8kBxB8s63Y
HtP3EjiXa2nRMZ2wTNu3dFuJ2Kpw/yRkW/Dnhav0qSldxgxvFLtE7s8V87bTQn9y
0vYoC1CAotllLwdEVFDWY8+zwH3+whgzbvfnVIHyHu8dcHhNBpGpJLnU51SrmLCj
kfQReICu/yitEFFC98PRSHdXtDSuBBRn74e0Ilap6a5aKNlrr9TPmDxdGjf7FXSp
qOJ2yjm0xS0cCWEqEjXkf9MDFEeqPsc71vPEuBqVUUCKu3hK5aCcxJhpxv9SBZVF
cZ5EtXRTbya3/8l4FM+/nffKHrJuNSz0HzT2XcOVWFEP/uhUxXtPCb0V0ah1pPez
yDvVhMoLYZb/U4yPUZ4mrF0wgF66pj3tQIU99JSUXDp8qITZgMVZmViAhzLkpTMc
RgcN4f7LRBQJwmkToQ/JH1vFTWGIps7qZb1QAskzUxQyuLIFZooWSfXNTpFbbk1x
PGPgXwyTkYG8e5qHmCoztTvoOPtTBsNzN2HYqBoXtWGWZcc6und1BugxeMoLLEI/
Y3WeHpZcugfcn187xj66knzq6elOI5wNj/rhtsEbVc+RgaMMPpuA2JSUGDI6HlBO
KahqGMjw4qPkR463SpplEpYraWT+JpbcCChxo4CqIpo7iCj85ghS9tzGVuedloGq
lO/1l8MJXBlb6zJy7gkZWay0PwqKZGLqURS6jE2yFgSaFTTxu1waSoTqGk2TuvFA
KI2sOJquI2WlMaQAwccPxrIc0QrtO9ieeQJTO3H1cWTB8MWn3bMrdfIRYTusQK4M
x+HxH2AiEkkQ4VgYBoNqKJrfUDLT68bGHo05arYlrNPW4D7wwFmXLfq2nd5f0xHK
x2wKL96yFu0mkYdy+6oDLjP+1bvsFOLW7AfcTibApJn8zP24vNNIeUZZOmidcyND
MGT1Shioe/0QJpMmK1pCbvo+0zsNpr5nH99xNHXxJYjOm7m36QG3gXUDS97ybHyR
5ghDIy5dCy3nkE1M0NSjQ6Vn/Wrn9uA38YMkHdBKAHZ8U/d8lx20927+MoygkreG
A26QlOwUUrVIljPiRU2fxemQ0UKt9aEUv9ICRjdLVrCYgtuX+uxd3wJhY9Uf5ldN
8644UB8+/vLPLB/JDD0ogiHMMOvKc5XHwYmc121b7HyopC2p9TTgsb6ujLKt3JtR
7uCAN/hnFJnhKKHrE8z66ZE4mk9CVaS7sEcUxhOY2a6cEXjv9JuxQ2idOBKm1fPK
NSh4KEG8+S9xr1eNoQJBlLGtFNb4pUvmhqwjJNErkUtfD4VAjhax2XyYzYvdLx/x
mJGHWx8HZ0NavC6Ms5c0U1AI29h8n+dF9sbqHcC3vQjNwUVxxaw+Yk/pmBZbyiGO
FdRnkRMlaihZ9TF5ML/la4s0dhCr+lFNAqG5WqXEV1JGbOsQse1bOSXtoj7o9RJg
Zke8eGdl4093tsXMTOF3i6fZWsUEQVNo7OeJEYen+Ka/lpglyJUQAaDuZM/r34/P
SiO18jcVHCzuhr9L7d6Ac68RWmJ+P9d8stSLv8/Htk1YAO3AyihYjM7UOlwSp0+9
GRlfVEJVM7bHRM7m1Ti3v6tTH1ZY6oLYEk8UsbYdM1oiOQTeT48AxY67uw1Sqsj6
Asjn6Pvlc5SOsS4kqJnLRJQTnKu7Io6Q3EVlXJ9V73fFRurjqFe27CrHB36fKzAO
A+2lEFVfFm32rfHxPfNdX8NFcmZqRjd/6MvoqtfnLzDg68s6QYfFAIBEYALI8mU9
frnQFIR6/pq92eOZp2iEDsLSYkhe9tuafL5YU3UlJ6IGPWMtnBoGeK4obwgBp7Ze
uvYAOWGQERoI8woF/a6ItAzIF7fu+Exh6kBO86hDN5c/vp46OBIsh5WrDdtfKGnv
ItbLJ+jWGpS+CjF3oFXhptOtUjZFZFklqm1crprPOspaQgeOVm/+j8UMqfZ9wxZH
G+tqr+G2Ye3nqe5D8Oz/sunrEIbTf6x7H6Lyc6xGgug63NJopTARHgNhXRe9K2sv
uYgUwplDYYoj7SD7v29Qumj/EKmF6LrY2iUoVpOIShxs5OBMegMUVGsAnu9Dun8+
Pr3VU/D+mc1DaiKGoRxreQ+TtJQurb7vvdFbHf4CMhwHizXQIj+QxS8+Gu9cZ0oa
ReoW0EiaDYTGFi+fx4LX08sUCmPUS5ZqgoC36Anlx0Q+PHvZQ6AgPhEiRZpHklxg
ehBCZAVq6JqlnIRXzRh4FbSECv/Gc75PHHbf4XDZNEfzmMJ4EFhS/ksuyt6Oi7jZ
6yS+b6cRUUXTxxz4YTv7qWpBcyed2HhPFqer9bSdLbUlXj/w1OKwLWDFhBZhmdQi
ewwsCvuw3SfA1/rmU4w3o04l8N89VUSp64b5rfkshgky6hj9Hh5roYC/p3bGRlNv
SDYQWV5tT9RZAGyjw5q5Q8ZbtQYUIMmYXAvYuljVe/I8MnVQZtkyx1JWfqnkJlHp
X6q/9O/LyKarg6GlRiJvwd3mNM1IBy6trGaSxOdCg0ouTipzd0lVzHIkUH6pQkGl
+Y0xnGHdprXqcRbtQCnYFeOuXTRWuMDfcgFB2sefH5ciVSDlckeynby5FAhjyzbw
Do9DxJlOuqj6gVPG+nzBF2gIX+wf8E//7JxO7+VF8JUSDgD845/c1lqMUw5mBEM7
uU1UI6r70V9JRrBuZieRwsDyQotiEQGiZvBFS8aXe4fPEMpaf6UTi/ROkPlpIt4N
767Au0qShfRsG4juAKcrY34eFqxsPjXLdb2Hj05QRmfk9nRHJIqh8PXbFfUW7zv8
Y86dj2vNNsNVUWg16rpyNE8V/9Xt6gNQYdWE+Ds0Jxz0hi+FFYtMwqmkNRih5l0C
A0rIi6a1WcajT8r+qUkXMp9YaGNFTtFH3J6EyO1FELmmsrzS7U1lud5F69uyKkxn
Z7DmLq4RF6CkAIT/1RXp5+LhNvukgD7EAshQM7CalqipQo4MrKC3gFIZgNt2ARMH
PBmTIpgcGljN/gvsof25YnoM/K30U1ln5xMOe6TUw3A8wrqIvFpiXqcuDU7eqpGN
yPaXBbTbFMDL0YhSqFzqFH6//WQoL6HcFz7n/19dTJ0TzT3ywh1mLjDAo+gyA1Uf
J9C70ZhBaiiyh9vw+XWSz5tfg9myta+ousXiXJkbc7kYwfPmfDOjDR+EvUztFAWn
w90klbdJrPytNSLdPCR9hiCC2MSvQ4Iw+ZNLPHUvDRouxm1ZdqxA3PNMd15mVyyZ
ky0Io5k4fAuuK8LeY8AJyUTpFnZQGHJTyA2W87OaUKPB+nv4JAHNQZT8TKyNv5hL
ZGFRBRY6TwTDNja02myeTgJlK3Cq00a8bP09KcvfJJHTWMql/TnNq8Eozo7XtKUE
W9Jtqe0UXI6zRh9hrF0ftt1fzIeNb+Q8kiPrw8z9IaJ5GhRBRyza7iJQp8r6WYQu
frCgW8mOPayTJwKUZ9rujsvYXFcMwqaiRz6ycUQ/k/CtksnNaB15xczRBU/COh3G
hVoZIsTCoHR49Dd4jEI9rchVRaJi6xpDZ1k58UQThs0fZVgLP3WQZYQQlatpw4YK
IwNskJly1X3VE4TIKMWPBClBqLnFE0fDfy8fRFuWobbDPPtqJcYskvMThLY3648B
u3AnClIIiecSJbHQWZAa+AoRtsvbYsdIg18DZhj4j+IZNrAVpfucuLS1pZT84xhu
27ttIUaYFqB7fNfMDuJ0q4MDt8nGdAfKjPu1UdpOZbE2E0vjjn6rkghNjUG1KB+Q
omFMGl/XPRZecSECmWTDXyq3QWGw5+qOPakJrtbIVzV/sS3JHVFhdz3r0hkBKaXq
mmV4GUMrVd1mvVcSijAAWx2nMX0sILvS6hf0/VwMj4V3GJRnVvUDKwV3bQnsg6EX
+FSOUm2WeTEuu5j6+GcrQEbynWxK64h5HsVO/SizNHva5N4ymjHSegUuffuWmKZE
jhnVmT93UHxOavnLwCaKsnYJ0wmF6lB4lwyt1SGyFXTpv0WOrdusWvyzavzxIKii
Uv+FKE7CsFX/1YqvTefY/z7Fmnr6BpV90r7eFa9qAIXPk9dS1DQx0OljgFVUKxpT
380Xw5XuWKD31qc73BSyHlixiEGZYfzVs5YhCOBweOWT25ld02N7iZv/4iWAo+3U
2u+JtJqgIqYwojQFZZSGP07B7wKDZX8zSP61GjD9KLkCkVAS0GKjEORAc7WuuLOo
KLx+KN2uPGe7Rga+6uGxuJHG8s4nENWSKuRlCW/GkS8qjCKSy5TrEiWuzs9faFZU
GYHvT0zsA+NSij5R+kUtboB84Dva5gWPMHgWHbOwVkY5/9TANvun5K5yS9FOQKHI
x5fk+hK+y2Aj4irOh4V1XRv/wUFrCgC8K7IYBKzTmGxXByvEiHlqc7t45wnsOcAw
6ktVJqk4oRz3XAW2YeUwvY9ZjjsUskPOlR9Wek+fFsN6wSxnNjZEOLY39gwxhne8
wRP/CYuBWVx2fKAoDibx5tkstiBj0Y1t73HKx7EMu1qX+/3yz+tG4elXWiCkJstv
r3QlNxv9V0CUOqx456BrYp1bI2r0EixyOYm+bY8Sdp9PNbwpGAmjpO022vipowQ0
p4sIYhc0BFEFzRQqYDtG36yqVnWCbJFWzqV3Ng7LAHwDXir8A3XgXuJm64owKhMw
3q+bu26oukSq+3fk9phNNAgj7BTHp14VrxE4ET6bcklT/4SAfMCKWvuJsqoKg01N
fLQ04Ax86xaR8guePt5Ir+HfhvSFDeI1JeGcxTICORm/weouXju5vfl5E4B5lj5m
0JmxQSasitul27ZiHF4Fv4G8cFJnHdJVOWN0Jnv9/dhh6WCiU2ik7VOxoQz9D4wt
KBt66fWB0ewLX6/rNdH+i+4d6dWdR50Ce7fMXT49lZilcEd1CCyz5D73ipq07q47
ZHdLhZ2PDr2cQGYKgahTTJX+SIKY7FweZetyZSwLZozoE1ReAd6vcR9xf64lMJsM
f6CbxEzceqf5MOM/XwExnYSXJzGjCZCE+EQa9GiXLqfrzypTkYRytS+kybEQEIO0
0WFH6aaXGjbNz63kT/6y8bdOOGfoI7eXdlk8X528QubJcAVqgBT7BY7NtqcuMsiC
JX32miGsQ0I4vRKFFnt1Cf1dqlhB1swyaXRdnZQUlkY1CpMUgsn26OZ9YZyO2UIe
6HNE+yOwA69Rit8LEBqXRsxQGEoDHBvSKWwlYfAJ6C5zYMYqePNCjBNyR6+Fp3fM
6AetTIilrTkHbIYjHgTP7DcS7FY+SCOOBhIr3aRIrcggS4kK87F2zQb4z+TixCCc
nRsppNf0xS94MT2bgNk7QLKgJdsKn40seRiUs1QgMSDZ4dNYQ8iU2pgvPujJXS0L
czGkEjKOuc+gSIP+vhz6RruvU6x0O5Q48E4/bJVTvEeuqKJTTTE/+Kj21a0pldiv
T7vMEyXY0+9gDgD38jV1uFCQGnJL0lX7btg9qrbUOjYAc4f3JcBs33Dhd0O1bJBz
pWiKbWidmzC7sIrKU6vJxMg0rjNhp9+jo1vidMNs92D37Y9wNfQlVHFQ+ARGsNiW
67x1DCGcPbBJdH6v1mcCZPqqq9Hak0rkSBGiYEEwaQgMmO7KYSEjZKZsnfvAdlB2
tIk/QntJHldtrjs5SzrVJPNDLywMtamznvqrvcv0R4jkOHPdm70BAMEJSyVm7c1X
DYXwUJ0gt/YG/4G0CUYylJJZu6RlPtkXRDr+SRsgYFF3s9vdyiCYkbzzgPg1RB6f
bmS3k5FjwwYZA5shpJgUEgyoQ5IqAH6IpTy1q9GxgIhkayYWS3GY/6nfFYrtdgqI
pYkn9O3tjRR2GopRChx/kI6mRaXDRXTkzdqzYXkISrdaBVyw/cUzGvlc+XcI9jDh
fF1EwUq5bcmjXUX6s7p+AhXFrdPTud1eNiSgs/dAvUFXrZUsXJSZexhsZ/rYzjRb
0tGuen4HflkTjVlIiKiZkd7WQo7NdkszyVjgu5KF6/hPN89rBBTLXjhfztvzt0ZX
mmRxBBxkyK6llH+uu48bTJCTxfvTbkQQ6tIzcSiJGglCg6MBq6kSAJ94IS6dEqpL
ruYJmsWm9iXNueXMfxrZt4j0cz7WbkXT76asvx4M7zn18jeQFOjKTT/Fjcp00QZj
UYSTshYICPSgmL5zOaJLFQ/EcnIWbxc7ODE76ULwnxCzkzVhizlveOhnCVON7bLn
gpv3upSWRm2qvsyVDl0vgAatzXlEdMu9wPWVl9+2iouJNNhp7YufpjmkVgQYE3WY
osAjCDBBwKtZMbvPQoRusqCHtfP8XhEAq2LAii1rNc7diQGXYfsViGe0E/UeR8d4
LxpCW+plKsk85/mSKzUOGtHxvwpv4hEiOpP54P/Up8Y7KVvyjWKtYW7NCKbGxDEn
738M99ep51f0eYE8X5iBNgWKD5U91Nyxm9ubYplw5hhPVSD4SV8VzmnU5WuMYZf3
xLrbvmXL2Pj3mUGsdm4o88CZRi7n016NWtUm+HCEL0irSSF5g3sa5vcKv0IUCh/d
ukKz/HyyNUBUYpXW1Qmi6Cq3SuOkAcLNDEhi6Yq+gRALv0Fb7vR5rQOgxrS1iO2E
Vrpb86pNGJfilGQx2JIKsvHLXNlW0FtYm1NRzefQnmADlI9TdFSWKWnW4CTBOIad
L6NnvD+psL3XKoGH4pygXbtvOZAz6n1MmcxIB7egmeB1593zBBUWDZd6LMNd1D46
LWIP1HOEJv0k/HoxnPvHDFuIWH8FRLfwbaowzPcId//x+c7IqVvi9YGA0GcbpXNT
qyrwVkl8Pbz6/BzkzA+XddaY1+bXc8CPCWBgMJQA5I8evjSA4iJm6UWnNhtavttH
XscTOeEPhsYV8cs1miCPiVLbBZzjy+CE9LoW5MmBJlZp0CZCkseAwkm41Hd08VD7
xH1B9LNipMhrugEO1BAAePswH9rGve/fKLzJwd5/mVPHzVbo0WqKZsMoc8vg0lLy
WLJ6EkyzxOyyzc7FbIIZk2VBOHsyV5s55v3WraYRRQylrCw/4J+pXbs93iNznDG9
KJhDcCUpvb4to5X3kDZu2HDYQX2jOb9B5r2NlllSrgV9wgWL89HWQeHPytDjnyEo
bCqiUy8l1dmRqkSwwcQTsHgutmB1zK3TM/A1ZNajyiHblmbufn5/j3DMo1tKrUw6
+5zJV7XD9Rs2AUpRg5mOoiczJHd7hSFwcuAnSyJAGhXFqZmOhDHbALG6GJxp7CG0
SycUhyVqbGjrmc2/o8w6UEdxlZS2H2RVjMhIWhGL8P+SUW4H8BJ6UwFQ3XcI+EeI
+KMIERkAE2Vq9gEn70xXArBahxEpmOK5RrmgvnBAiglMvgk77vvm0SbyxiovHBDm
PF0FFUsAbTacJm2CciqXEsDyq9olUYbV2DQc+/qyIF6BV1YMP8WWkxgFf8/n0JTc
t1frDxj8yRS+ir9SnYdI6zJH9UltvfkwrUT8vz6UEFmwEqdRtKbtS2OiQyHQkzfH
lpvq7MfdcIgTBJsDoCPeM4veSo2S2Vb/WM3aGMYG3CdqMWKzgrujhfjx9MAXpoy8
qX9IPTKdfx7AfB3cJ2BQ0MOsZFuzAO40fziLV3ouEuUPc3OHYAW4xSb2qPZ9QzJK
Q6uyorpQdFsZtDCFkECxDcQ+29lqfzi2ilELeLeve+IMFccHrecYcJLyb00YfWJr
i/+9UmeLsvdw/ZmsD1NAqVcEUYDMWTz0+TZ27jV5rdmz3gFsSfekrOPlFJ3OSEBi
P4yMXEegiNUyOCUnbkrBmiWqK3qMm4pBU7POx4vu9R06j6pzOVxi86igpREvSleo
hRP4YVociIM83h05lvFAIR81Bzbekq5auCol3fqvQ8KH+p9lgUzAgowfHMgNCoBP
2TICFc81yHGmJrJIA33kGYwm2UCo2vKlRIrzuarwUDVjvcwSqBYTRvpUm2Qc1rXg
z64ruUUuK9daeM+RGFIizt5tNSWWYbaf87w7VFb3yN0JuLwi9+njNOYew7BD44up
5t7co4ujTzRt2BjzmNzYjUFMgNC6A9pYfaSz69CTuGkwZOmRrQf5VR3tino9KFMS
luKNknhecjmt3z7Gj3+qTgdaEr6dzLG1h2u6to+VkD++EVsmT34eWmHoYu0YoyvU
EsN/WwOz+phw6OATV+t9j4f+sMVOzr0rAOtFj0xgpGf6LfkYI7CUrzNBLRZjLpuH
Si1NZTdxWXFTD7JNaqK2/9p9UUUXlN/GBDg3J8rWrKF6aIvU+ahTiaiKisRpw72H
sIXOBBM2NyPz9Y8S/mqLl0CWqb2pwqFYhnckX2rLe3M9FSLs3GARwiyWdtpiOkSj
tF0jF8+POne9ioeEHXtZ87EHp8Km3E7SJOJ8a+L+jNUSNkw0y9SlfdnWfN4pELrl
OBgnmTIMZ/oBlHUMkODxmM06XQ8n0mJ7JPTkmpFH21gkDyMGXQH0rYyFRFthTF9p
louoNw7HdCdnvhnaNykVuZrgiuhu5vb2MLgTPztj8SmNnIOD3WG/7EXH99A1shCw
/Ci+2Knm70Fxf00cdDgTdC9mjVAghOxHxHSFLnENx4Sc3mQcwYkHc2J1jICiBiwL
dDUFq/hThk5uY74up/MU1AqW0WWsbRAHYsJSehf9zjayuxME+sWeZFrTHE+11hZ5
6lXPJMbR3PUUUSsfFtGs++2r+pZthWXka0bf3vCO2BRTyQyzh89ZSllIvfGPnRqI
qB4BqYiF9RNF6TjszEF6pCRASGcPWxrNv+Q0kKURm3eblUeWk15ts3cHwMXnbOmv
ZDL7lz7/6aeciLF3l2eD41gAnAVNmj8SxrptflngNQs/CfcweBNCdZbiB/0AFaIa
bt6hxK4NwdUaroplIfqtQvLv0sDczU0O1py91s+SVTpTm/gvdNKDl8WHyqrK6xbp
CYhSjcLR2tzcKmib3Xu637ArRlMtC77v/xj47O9jDJRgRNHG8yzbO8nYko20BWWy
Y9px44Y2SP8OfOk/5Y9FLgGkHugCztnHx84Ch8G86SEfz1nFseQBJigRjbfT3wTp
noDU/XYn3dXERySt7s/Za39kLDFRZ1GVXynUcs+hta5qis9nH//bFRx6vWglNbGf
e7PTFxKZCQI/B43M5Vqn+AAATr5Mg29QXZxVTGY5WtOwLdQ2lmro17rQ8jAYnYiu
V0znsRct2EkcsQpnrlhRIUdr1y93XgycspYo/ypWSbdp621/rwK3kZBnYDmK2uQJ
CwN8WQOE2lJXWrmu5Gzl3A3QJ8CsuDEoWdj1AB110ItryDpEnW9CRcYLSGlqz1ZE
XP7yo+6YqKY6O6KknT4OrEJYRhcqEzCV14AQDpam9P1hWr4FZoCzF2HqwDXV1o9Z
4HsYaXp1J+00bF0a3P1tMrjOvBzR0vV8W7NKCGoM+clnZpla9S9Jp49Gk5+7NqMd
nEyZY6JSHbD/S6nmoQxyhu7ytSsEItgxwm3dVjUwz2lTd+2NmX2DPrriZZYm6JAl
OndoWcv3juvcQXkFicdjErVMstl1D8RKmOCaFAYs8bRL8r9jQhXgoCX40H1cL6fs
hffQGcu1ZQdmyknsHczw5eCdnwn+/CXjCwNVhSuErkEgfjJma0/xImoCucIheHvH
aUMgUW2eIWMz9pD3OSZcvlfnEaVayj9qZHj/Sp2Skpi2wfbb5Yi5qmwhDRb7r4h4
GYt1z/iYAYK1FOBqrJAlMO4zKwdtP4Sx7FP22ViIfXubsKWaGSVVYwV3JYwYyLOf
2xL0WvLCvYjh2YK6qxxXr48KAFE/3FHWNObYa8o4G9AZ+U0lQ6RuOh6NR5X53uHi
BAwjvB1N1ZHbdIHXa09nwXxolL04Qk0ZtQeEvWfKBI36OkPRV4LPvQVAf6+jF8HJ
FtRm1rxSBBCgpOP33/cpq/2JF9FGam49g51nk4l61eraHwMrYW5aFOoOEhjqxAI2
PHxPtuL0zQ+E9rUHCViZR0J8Z0CkmRpJxHzr1cJeFaaxU82IRlr7i/SKjLj8ZwAs
8zrtTHnhpnMhoEznbI0bDVtvo2tnEsfYr/J/Rk9D0a4ZbuzpiA1j09Qa+p/+a7ZL
DV5G9tnXUPj9+stqr6za8t6jS/VscGo89gdpCXbWy9wLgRrUTpbJbiWPYqEgB+Td
fjFFpPVFjLc39kKoL0kvyfgkQBW3D/AWTiPWDsIzulEFmB23SjHjvZ1Fo2EVo7C9
yaCtce1LzWT3wBrhKfopfYFxUo6zx1LleL/XNwWkdLVHr6Q2AZkQ6lf/URt39fbA
k98a4rM5ywTlQRVhBWSSHaByJUZmQzp3XXVPZ4KCQl11jDiIbFYo5+PAXqslB6yr
cMKbIrTTADZtXLc5OkEvaWEFv8nN3PTwUzpZ2wUilhe42ciRkx3iWX1tq/r5CntS
X4ki4+LC48/U6XF4z0a+OGjqe0rAqodXhgvk/wWDZSe5gLj8iO5l9NqvKqvosgy8
LgnyLk1Aif2wMqOtJHlCaSTHpQki9WTjzuzYD2p7Fnpg/y6/oq61DLF9MIQFllBP
qqTqwAvo3QzxRD5RnfynWgw4BHPpUPdX10lJaXTEKyC5+Fpp/IlMbUx0koKirQSj
ntPklcLjJ30SyqiVz3V5ET59IP9MGZ1vM5FwkZrZaYZIW+oFYfAISczJvB4z3C6d
zGQ2zMF7mj/q0gW4Lo1wcF/ZxyqQMr31zek1rzSM0ww9vXcfx7NF71aFZNL05dcZ
yY1Op5udo998ThwuR5CQj/Am8YfWcADS5uUkXP5L5j+pKPl6ZnvIljZ/Bcj9UxLm
ff7WUxf4OulNPu35Bi2qsiFV/eGZKV6gElHs++q1cMs9klMZTGhJpziIEMrnSniP
SeuMx5PGq//hoEddyQlgBSG1P+2iERdrQevWDhrr0JPbMphU1uZQl0Aactsp62mE
8sla8idWmZX5h5qW0HJ9hgTVzvM0YatGuIJns91t+E4gX4hvMjo15qKOhVZry9Pa
BpihSEiWOyTdTW1nZ2X/qCgbPU6DFNefbigFhX0UeOpR5XwV/GlZMXKVd1YZr34D
zBNtDwB7oo5UVeC1fStr7k2cy6491uigfBGzwQ3diQvZ/99FQcurXz9aOFJPBG4g
CzbHXSDyWPe1owU2CdlHr87vHFJnkW/5M47t14NDOmhch1YRsxjeMaN5y/KkK0g5
kzvZ9o7xyDl2BmpGeQ19DVzvEcpSTmIbVNbfBQeB24evBytqW1p/+AkwNfzeT09k
/lUUpfdn8y/DZfM3ozCAX8vbAL9vGP/A5tthgfQib61pnFeg7fXR9NDtBFuOp85j
BQ9RD6eimB6ZnqeFQORPirTaw6S0mc9CdEzEYcwmLN1ty2aBiogvHZ2XCsYFbYC0
vfkSOpgFO9LKL/BTlW/O02oNAQnyaX0YDllBm+Y0rPlrNZdFaAKmbREQIBzHq++/
gwITjbclgaZ49HMeASqhi8weIrEURjhOyAqFM/QfwcKS39FvxkMwc5rRubXyGGq1
uDdkS3E16p4cW08t/Z4UbEAmFBrYGWWFlcYjBUptHOWMfzHeQUY+Y70HYSNRxl/Z
WXGdRwLkLODYUNnXqqfXNWf4jO58KUPjZMTBYFyFRrrz9v4n7ZaoBTEMZvTdb3P9
oVpvF/Do5kjzQuoreBkbsAJKKmYYygrp39pRpkFgNHWFP8ssl4Xb1Itrzk4RoCNa
wxAjUUIA3259vtZ0qHg2WEkJ9NeGxEvembbHcNLu6pMFQSNOvVR0yUhbSdRPa9zm
9MR1z5su3izD0z76TzDPOL+ekBszxhiealno0sFH0GpVgmHjVGGdFQJKpfUUHpEY
unwjTtOOxmF2pGpOtG21lVja8lXLr7K9+QF+s7jpFsTWtyr2OT7LaaV28vOOClsl
brEVCg0vDcLfF5C8Xdk61jlFLhLE8mIp/ROoD0w62M1836ETHalqtvbkMAlyK11/
KEutYwcoMiemeHGQFmZVTXPdyDrrlKVXMAOAYlWCHeOhIusV46p92CZyvDsRqwwN
PvF0rYmf9WKmBnfPVpB5Qa/VZKEhc86jfqty231+IRPa74+rGsn0WmBsUVtSz8JH
mKw+e+y3HBQrHp7DR5F5ezM1v0XcOZvgJ3gQcLJj5n1DahQWVU9YKugFnGxCZjDS
AkSrrOV6TkbqBarJrVThkK6LsfOSnOyzsK7filuxtgPUYlIvqJyJOREkXs9r7LOp
dTg5MQI1kT/ps8G5ZUiovujEgafeDRNhStLcAbHVscVuz6U5qE5cFupbyfYvzkSf
Tj8FnWUzFTstQhKh017LU8BkZKdGd/jRuPLTQmcwhFo8swwbehVbWF1pH0Rjynig
nqw4LQWfQLLwt3v0p6SgxFn9FAJ37/epku0MXW8XGwY0Jx50J5gco7gzR10oE8Tw
M7EL6R9Ijbm7oY8MiryCPCbssOHQZ23zW8YCHRm3L2AEnBZtxt2P8GNXmrdiGSev
htv07hDNSqJ6+7sePSdJKjEHyDtC5Qnp2trEQ/qMARKoeBAfR4z4HfcD2LsqY0ar
5qbYw80b2oHEzGBmRvEHwgxxdw3sXGSAYXKgv5Gh22erKPeKs1UN/YNoF2u7awAT
OdF9GpKz3Q4slChc6zZHSyhv/jKUOr/H5ctV3AwuHxNDz2hu4dgHMT2me9SLDH+8
D9C1zsC8Q4FxkzGlPxzwMFQEZDl+MS3qiyZ8FvEboo2aU/vRpx4ntmyBj7JAGKxn
xxmrVh3eQuWzsccG5S+IwM31F/saFcoNUPfUugyT30Or3TOHD28pY0o/Xs9BIrUx
vUEfNOrZ4xDDAiG99p1ZdFIgf9T5MIJqmdZI+bAxq2EglcjEluEhLsovaQnDBfGr
7Nu5eUy18uq3h4O+Ri3fA6XAScdgVFO0sKBI1rDi1Sk9yiD0j1Mnid/TQGn1vzlo
odYP3aCgdR0L4RSWcnK1nZA+ZOTwFK5NpL/otQAEtOSX6t4LLEv8veKx5mBWYFOw
sR500p+3ZaKTPYcJKGqswQvrV9P5MJdcL56xqcH0oQ2AIIFvcv0rfLWHbCyO9/uM
90Z+qoUrkaiJgvkNqiRiWsNoAdEr//MDHcIeKS9YgVzXBcad8whcG1MHgVsDRPW1
22Z8aYsGJw4O9cDXR1ApdOQMt0ovZndnjVxBGpeNhNUzOZw0Q6IvXPOqPYC0quqp
KgiV5VMAb0qyzsThBTBl6sO2weU4hvr6rJcPq/+50wTf6S4EAs6gBW8nWCzuxC9X
743xXCdcQ2ttt1zoJVtMck1J9xTZljQhwCAYan2s9Y5snFLVqHpAR1A2FdK7cgVN
P7MpMXtLV+gKEK6LedyewpSYePY318vbSWKcFJtdX63EY+0qURpPeFPG9Lc1IpBh
aQJQ8CJgOSapk10elG1EjALT9sX3IkbZ7a/6HrKBIQgKBr6BhMoIOWodsNZGMrmc
cNBrUtqsjm5FLCQANr+iztOYMwWg6j2XfmWlW+KYfgTTZJNi8cloCEbRHI+XMUsA
8pHk2dZ03+VDsLn2bdMk/419hZFCIKkMyFzANJEweloZWjDE9LlZZSWlZB+tN93Y
bOIFbntKCfDMdA1/h1Et89AJTczmNcOLsmHIg88j38G2weCZXcsJsMDnxrXr3uMz
CNeMJZ1FOuImBCRgrFi6fNDcC+FXmfPxpny+H8LsEvhhdh4zryj7+jwp9cvyU/K3
l528O6g1QTHQHwvXo/3Sch/N6PbfICWIfpa60lSpUquHEAPBER1J9t5RRhKmKUk+
MDYgb86PZpm0XlNAl8GpldORDBB5ujd7iU1cGtzwaeThA6cFTP54vWYTb1//vefG
fNv1I1jBFMPR2ml70KtOFjOROequeFS5gpAzX/eJF2rV60jpmUxu5FZp2HXXRdFo
6ZSmqpsD6tTNIBylelq6gcFl/uZhjwsJbmuhPxzVfN7kdvUh3Cihixz9SHnZ82x+
yzqF3lVMcW3mj1ntXorfns49EXd7fVtLJHIfcNO05hyz1aNjfK/jNRablnFzAVGs
QtdUp6/Fa6Zfwz4OUnD87riz7BZnuuVW0B40ir8BQEt9MjbbcHkMOSzc38Q1AY4v
T33t9Z/8/P4e2d1UHYvU0AaT2u3MLlEb82mNxCzSsXRduBSb5ebWLJcIO3eYEzjb
pwNQHlyfpOom/KVyfqihlss+zH0NQRXj7GI+CIA4hJoXBfM6M+PWFo8T0l6MuERw
811C3HToe4Pc8rsBOdYhk7138odzPAlT6nnxk3rbVUo5Ule+DT/Dbg1zcN8od/M3
Okjlk7kXVPLYOWqKMOMDSIExRlP0SdCaORyNdemO+eG+ql7pDozWDvEJKctgjGEG
DjQ+/6CXCMmhRKdaAIMSXkMSlJH/LbDJzi7TYJoDF9NsgrICCviXhvY9Q5emgGh5
nh6mtGtUn6EFx+50wVhzVAEEp2Q5EzwB/Dj9L+631wF+JH8hL0OHFRJs6P0b01Xb
JFaAbbZGd/EPMFltDth83iW62G9uLG90L3Ym75av47adsDX5cZYIXmKgth5rxROU
4jwlSK0M2Rsp8FDaz4UdrzFksmoLdd5pP1dqzfYTjkbhY0jCBnTQ9THj6LZ8cfqw
4Zv4cuVGEFEvBaT9y8k5aAhCi5BTiY/W1SyPYdOd3EdAm25nUB6BvtMH7K7smwAY
cpD7cqE36QNLQcBE8KPAeD5OQ/6P7PbZjhyd0PIUTGziglCxYjDOVgbYAD+myRG0
IbI41++A+F27ErwvGtQKR8VB7zx2gs8WD4yB0kRYFo14adBrHIt6usQWQzS7L7jx
Qmz5AeSjQZmjb/mU7ja/j5vzLcJeTXXaV01++46hO0NOvyPjDE8RP/6A0SC2LL3j
uu4Poal0jLNLxc/vE6kgREVYAB7Ca6ZlsTtNII/j/pWmYtKvbTu2PpCIBjBJwb0P
AyYRgBRQit8OtlTa6dLnufJ6jWTMuC95kkZIsFeRpg1ICER1tnF8hKLPGV9wTnhj
g1xVTubWItNbg3cylOJlDAsAX59K8SCANAak6MGDLD4thqh+32fIJUMywuYLU6mV
+nDt6j7Mg4KJHsKViBoHVRKFLwV5GUKhSaXU4djmkG8naE5LynpLUZrfSN8lvW2P
7Bbsoy+5fQD128VVLb3snx12nXuINrvD3BcTAb93yYzXrPs3CihComCePxf1BBKi
4gR5anZV9D2qNbcbZzeTmURqO4wdiK5hY+cxfu6o/94y2pdEWPR1oQrpyhcVws9f
RJQf84sOfe6EA0fO+wBgT+Ovv1U5Prcqeh19KBB8BNhIdUHM3iXlPaJ70jWl9ro6
LWwz8XapDVajmdVDFZW4fP2QQCtcx9ShgD1wZp4BuxxfSNjORXNwYWAMT3ST1bk4
4+H8rzbwztnsnNicD379G62dk0amjty4DyQw73erbEaGAQQgVHac3Cr9Tu38ZQWg
mKpbEWui2rVG9p8+p9pxQ2sTLP2xjSQ4EdF78Yiav5evBxIT+sjmAA4Khvsn3NFD
4OnfyvOafMFw3Zp/eSsPpmwIYLTQ88iWfqJaCcfJtH8WxMS0dnyOoFSei6EXXIup
SMCK1w0W4JAUVdrZ0GalfKpmCIuO3Wmm9SBNStnvk1XBcqseTi03c/yxDCOEp9GR
M+QZKPXkLRHbzVcLN58LBTqsGSTuH7GVDt6s3vqN2qee99mKXlIU+J8o6/lGB9nd
8zJFavsPy5P5bejP75e8MAJnIBlGmbugxdRzJKbxif8O9wLiG9MmbXoD8smtmRUw
fjMdjw4TRVCsnZnVGXwtkd7lH+1vpc1u+i9+OMU3n8hsEjv06gSAJb7vsS3mCo2Y
HOSc1hPE/hV3DmaR5IkxvSTURxyF6NqGdg2sMmi07BLN7vLnAvAOXsAFrhFdpS8B
rlmtucc25RBh+IEemL/PQoO8Xya1hQFHKJce8k/pFU6W+OGBdCBcnqHsFJmCFzLd
vHANDdEkazbRz2W8UvBCTQWHLJDn2VdPxevSc0ePG1yNgBQB9KAb53wVVRMv7yqu
5itTgYY0g1HYVdKfbLwCX231jYYTFuT9UgZwrn0hKiLV9MdnEGl+yFwGpQPw4ZMk
PrUe44yppw6iZ9I/0yxhjEqpE8KMz/nGOCeRsI7tj1Knh/llyKNdX4JAG64H+0Ix
wKNK832IOS9YJvT7ZP6ou1w4NYa3O0M8zkwxoUiLxIhKxsSFE46g9XKBPemVo4FR
Tk1YM516unE4r2ObzHMcTr3pqwZn8gcmqMygPIIPbiGAm0PXKDlqoX2iA5yBmbkS
HM5rTtOERfbSNJ+FI2nADm7msb4HfhvKNy3SrXdA/n9PxGlyJnabMJvz1UzzHMIq
zbMzqAnpHSfNL9lYiGKblUPyV7IPyokpBYaFbVWtHQlfC+eVdoPa0MK3MA3DKE9v
TA5JAhKWjKpdAhrQR72p0QF2RDH7oXbvc6X/q64JZIKGiSB7VQO9gEWp/CfIT+48
Z2I+ZkS1Ddd22kSu8SK/Hr2jQ07YTnEg4pHy4a6ZDnpqGkiGi3x0wdzJ5aZfIYNk
q72Ke3fKs1mv1y4jVPdtWB6Hp3sBB+ZY8tYA5CsHQXiuKZUA6vZYU8GxHcSdkLcv
Y1S5Q4q081QRJUGFx1jI3fRFUKcHhnEBTMmKrPc8ftAWsKRR6mz7tj+jzYQGkDjR
RRRSvPyvLE2PICVK7Ggq+zrKrJHtaBwCnYvCyVdpJU+wJF+eCXbKHdAH/i8C4B32
zE7V3F2/zihC3dzA55gbB/nTWAwMlQK1i+0QMbB1/nVRVg+c/bfxLhWkLHle+uZe
anSpujdfujH4UhPCy/mXs9xsDDC8UrqDMIuRSU+pFYZPESJ+O+nk6tBE14ZxrBUL
lkLsOOQ3j8O1RgsS9pwK1xDFvLnUBFIT+7yWyNeUxLyTnxDi0tWHkSwlbJHMu6XR
TAt532lbUdMJySB8ztDDNYddF1V9u2qJhTvY9vPp5TRVlg9NcmwQ9vKCxtA1/6zg
0g54zKdTWDS7zFBgUkoUBMJL701py1CtsYLXgBOxXfTdkClS3Y0ju/h+QAQ+wS4x
Z84O5gQ5ez/u0ef0Jm1xH9VlIpogNzdph8Bj/AmuR16D+vWCPXeXHbcoZtMDmHhF
yTUBBaxdyvVuf+BePJtnLd5xffQyaCHtwrUOShvPq8idUQgPEcN8O3wPW43bzTW8
xEgnhtFUNhSjU+OCKGok3eG2fWYoJ+lA17AKCqh0mxsNMtl7Q9OkCv9gTu/lA5mT
R6a0plBmAwrvna7ixJizsrfJEi0RB8bycDxcPzz2VEYOldoot85s2GtYOgn5VEoW
DVG9LHN1rOjIInC5bRaaLiVtGaHS/dKdb8IBYwG4PWMpt/fxtqpjOdjb+DHUWPn6
Hrhqt1//B5XqeqXA3Aueff0rKlrPpI/ucKI8JPyCUwsJoq5+6W9st49N9HvEiBow
0GBErxrFGaOk2ehma56wjV/YjBzDGh3TbOlp+kpue9UMOtBg4Fe4LrYH08IXJO+G
c0+2nkyh4LqpJmIjJ6O7qSvg9NIpoAW5VbyR3s6Z9b8l/whTjFThEE3dGnugTiqB
CNCZBousL7rkCsKcHtonSzWnQmEtQwbwCX1fsx0lASMnYHsplMZqUJgq5mQ9rryF
vEz67nYkyQCdWMgYsNBuybHstHNsM2h24ScYfcopOSHMIxFkXUfHPv9PdAzPY3Eo
9+vOK0XWijeKA2TX2HdA2XBKSk8ryvtpvgBg/JFTNrHV5rEJDtyjsz1EaLsEw4mu
HH4M0XAQgWl7yoaXc3AZz6PiBc7OCpFfbgAttj5KY949gAs4nlSkMvYp0GMQNT8P
Frd1LhsY/DYz+zIwgD/9KVhPyPqcNiU4DWE9EjzlZWJbmQL2GnbiH4l3b4Fpf6/M
Ei2D43roJxGeI/KrARy0lIX7OotGe14hTqDGZ8XcK5v/uFtsghfIw66ILvyJOqe6
K56RKJ3dGb7VwpcWy4DlmZZOseH6pVT0f0t6Ao/mrXYp4+4EDU0jeO7TknWUrn/w
sHCARJZdc4xT0tLAkLE0zNZOWRY/1P7PnpStArip3qFrqLSr7Hd9BcEVJvHiVIAf
rjWid4KHE5jg3ob9oeE+W//oLc2FT3bak6DiwwoDJooQw8VHKqqkwtTGha628RuL
3iKYIbrgUno+AJhtuMv9CDMZDLewkN4g/F8ma792XKjnQU7VX6RRaU21tlL5u3h0
6RaQMGSwpiper5gA5rSVzXCthXvhEKOXVutu9U/9HfaKMKTtEbTGLbXRwgjqu+zc
RaLXd6+KG24xLflmoAyF2RSsxUeFpFe7FY4HZ1uY2G8SoEJfEBjO58Iv/E4nARSD
Mx2CLQ/ENJFRd6T9e40LlaqZm6xKwpJnJsZUAInJw3F5efexbCSZWFCdFI+Kupsy
GEYO7QxcwhUsoywhOOuaR8niKg107hgkIBu8y8YhyHEZTxBr2Cys2VnofoGM+UUd
kNq8HPxALTnl5uGXSC1iQ5wmn9aGHNxyCHAosY6vrKvl/LY735b/91Rtozj0zLJN
RGndU3xRiEVnVE7CQDtiP8fCfB2OW62WYW03lVlsTS/cQyQQNN23iET49iZ5HuZu
lAyZQuWBY4hxFlES/FjI27qgBQjxK13x3TeCI9FtEFFPRJwayo1X2EDTDf+NbN2s
EAopBIAiahKNyzbxbdAEbDDEvSZtnIgikwIlaaO7WNKtgM4q3WX2aSMaIZMnQdEO
n+KKWEMr6YHvwRFImcoVku8+YK9I8c1803ix+i+WE6PoaoJ5EjRaHhX5eqa5Sl2R
U6DYt/nieOdOGDy+gezh/msU6L/lDcBY31jSSRwmh3wOO8HWY733yWjKpnXVRcdF
hfgrmD8cDXgnD1Ie2ahyiRRAI/PoD69cYdlGlji6tIpnehG7qpy5LEZ2sK9nc2TR
V8XO/Dg3x2fXptByTDCGJqF/tJnmIshocGM7SkuaEUwVeFmLhNiCqGK97/EFixFT
a1130TQkf5JNvxhX4oHLodcO45Bvn2vMt7vaVDAwIRvPtZi2dB0U2I+KK0Dd7KGj
7sLBr4XobsqtKyZzI8SfX3UzWRzYLRb5Ck7N4A5wudQivx5+MJsDP/CrZudZSBBS
426+XUDv8aN5FDNP6HguvcTb6fGzBANtF0BC4YpDX6LJDeGDQTHSrqeiDmfiUy86
bcUrP9LbaZdlGtf2ZzyxmcZc9zhgk9/Z7ZfY8cxvepw78wuMDKA/SEFFHZnJbZVO
FlJ2V6xOnxsdzuIfmFgTDoIQ+80sVTPkGGh0AS0T/r7XADVbsnX3FGodppYo1krn
p+BLcAC/8bHYtdhPGlILSXrYUDCxs6BTgYpaXyMA8hM/dkRBxoGkkQQuu3x0wsVi
W435xLn/wuDApMCLW3knU7/RM8YmZRshWIDVULyMDOF/fC6eF8ifM/MZ2PURLdA8
JkQl+ZQHOuuv2lFEYaYRTTFdx3UALCeqeSo48CYPJg1B/6Lw1estOE3WM+YYOzB9
e5P0N74bRBrmg/4i/FOXPb4Xl6mBegBOSYQB0UcavCvE5OfQapP3W7ajdnliXYpQ
eal4oh6sy4IFbNVF1UtFDI4C4mdJ1qS39I9ViRgFVlDbtOuEuXKBeYg4P08pKrgA
osSDpUVfsrL/p5HD7xvhyS3em4TeKLFBz7vcgNQKMzstKr6uaQJAbtKYk1m/ejf6
LHl2YFkhIGM0A5TkXxdO/rJvvvWI2D+GmPDhW+b1CAiKyHqSFFn9jTrcnCl+zcoZ
VBPUCb892jS2G5uxohJL3KpOkBmCfFaIJDP5sqe1/uxdx7Tx2IbNbzp0k+YbSiVh
k88Aam1gguK33Qago87cv6JG8zQ8xnTdTd60+1UmNtsjNjDgxKaxnzKzUMSVIyxw
jqHx22hsKpfip0ccG21ABk3/kYG+6IVcP289w7HZq/lTOyCL48NgyVTFuxRCkXgU
EWr9lQTrbMtdsB8jXCizUJi5DNbhplWIP4bskJEZXta12rf0i1/6IwBb9cLGnfbl
Hon2LwL5xOJDdT4mmWrkbAs7xPvZeC4ZgIm33rQZweAXRZs6olhiw30Gjy181Ccg
H2uREwpWgCPTsCdIB02NUsyd2la1qq7ZbM63gq9P7Ndvg/tiRuEd/lPeDG9uwGXI
LgMkE+1eJYL2oojPK5k4u0tiIiB4axEyTjnz+e7S2JJ4ZNvD5A+h+kPfoSma33GW
oekaXtbZkkqajgqHt7SpOdUjPOlSKtSkGGwOH5tei2TnQDChzyB+JhKMcEaChJjO
QS0fuPL02KEtFoIRcJ8AAPP0hUO7m7WOYJ2V2H7BKUuu+43lcldX+mioGxuIAs/6
n6gYLaATlleLBmnId9osNusXd3tiXat97Om59CQIEIbK2mxpqAL5sGOIPzsMhjKC
JqKB0F/rtTQDjTmNhdzpUxZUv4rtjyffahTVumtaamW5KQIT0GXGx6MD1E82SGuJ
nubRmI9Ah9zi1VVpDjr1RdcJFKkuvudA0dV7Imf7QpPerC6xAmv7mhTBHRR02HX/
iA9lEYrN/gNCqzwqY6t08GLZrm2/fmiZNibjikVkrc5lQ9sFcOeu/vFbTFmOP8MM
T224dGzgFPXs9pYfY13LvQihoJkkX/RsA4XiuVpO7fyVJgwq7cqo14sIhYi3aRcS
BgO23fesL1lqqZMZTd3DiQIEPk8+XVaUBhSjjIDiJHP8BhwQ/HlUqsG9N4X0VT/q
RI3nsJuCw5667ym4N46x4wq3BqHJmv9BM9fDyZjqN5ggJXayWEpRbUEi1BhUlql+
K9bCLLokFqcxyB/LHlTQW1nOvD6ndXP9ULbEqPTPmExJHSXAh3Qy3KUHLdxuwk2+
QuFy/Rh3/cm7kzyJPPGxBDFJHT7bY71HtxNr4SGHt8shdnAe8He0iTGw/XsT16gW
4B3L1XPrmaIBdR/fKe99v7NL/pNtNmYwBCy/yfkWlzbhdE0NtvhPanilGJn5llhT
HYxZGh6wtWeoMd5jTFyDJhGcIkdUBr+kNO3c80QYx1SISDcP7sQ+D79qNTX4CJrc
gVmzL31gDNYz+rOn9th68g8hgBpNlGORqiizeD6vC+etcqdVZcCWVLcvNjfLmLQO
9fbSMhUvrVTK7BCCQVfMDH51rRuWvKF4m7R8iEwmCzHRgYjaavr2eJM/4OwdWAO/
CukPY3izKauZZycou/4/rTJHN0O+7BlzERRSY4laFhDBpxeNVgnE35sTOCjmn5rL
B72pNzITwveVkRpKC+jJ9Yjw428X/4iVEpOikinApUs0efDXdfl1v34I04GAtmYN
xx2Ql/tIDSvWxTUro0qGumLKCoF7VXZVV4WRExB9t29RPNx6Jx6YnPXb30lNdVj7
vBi3oNhdR5/peDESfeUQAshRLbSB5myc6zxxrsR+lDkuZQ8sOWIrvNSpURv9wQd1
WPcGXUIadmqrjAaP75hjrItjg5tYFr9zDENuEcVtxdv5KbjSH2iEt53FuNiJVvuH
HlfgaDwXmFDRBcLlTRnnMR5KVPRU0tBCNnvFpSV5fE1yGLdKOqsvPCttqTjMD4eq
kxj9l5fgSNJwgJZTiaKgipaB/Y5XAZ3jDRGlpC7S74vL7b9UVM/HlFVvpgING8HY
at+zQs590srGWvrQQbjzY67KICoBpFEJVNGOwT3LY5OwT/sExvqNoNLT2tc857tR
rIDIa2Y2eWRQHvMB8j2LET6mQt5j/A617Jd2/xbJVlcVeHtbflL2xL74sq6BtZP1
n8TMVz+C158WoKrMUovR5rJ8BZIGFjfSFLIwx47iO2gJNiXLMdabsJtm1BH+YzeR
PnYB391KNvxLhkbsCHalObEa7S2CsUZZ/r83fjQLJlMe/QtVYRP5xzeeCLrQD5Wt
tP423+i1H1Owly/tXBiKot5DdNqWuDx2GAiGc091e5YK62Ieb8RbHR4C07362+lD
Lbyf9YSmmXYPlm3tnHDyRPaLFqLrNyJx0KY0Lrlenty0XHYZ3cuJvTWbPcElvcz8
gmL5eo8ViklmYonPiBeFu7QZ4l7NQ8xfTkUiw3kMBBAfsOxcuY6LWtAaUFJGrutH
06LBTY18rJAwGzIN5p6HnQvTG2i0rmTcMJzIYjErt+VPZlc4Gzc+f+u42xrhujfX
/FrXKI2DMSQ2TvVN/D5oep8OHb71wQsNYRgX/jl29X95K/GEzpquDQeTB1YnBy8c
4GGzeyYPPTVogptfm4UcE+vjNjiSGMiiHIGPNtsp+p0zcthJZQbVNJZ3yOW2H0O+
kE8GG+Dava+3PwEQue5K/EZp2+cCDMGx21CHZmZqV6fe58fwuj6QFtIlHPFt8Xua
xDq7NROIjE1O8v8yv1KuA6ad3rd6HISgZZLcNqsgba1md3YYf708ZgW0jhbbjB/S
5PcTIVXTNx0+IfKxqsags3QLpfpwNUJWjk7XFmyjNlFNALdj/tfRocIGd+BQiE0s
8WRLQLY5VJjuv7aq/dEwIbjyiRG6E/gCc/JzpINxjR1Tr/lvNJagsLhP49VU/xsJ
KYS9aj1i95aIB+81bf7ztFArWgpPMBfuxFVTIGH1pAz/y1Xx01/Q1LCy3/KdRWt9
1HfIuFGf1Of5Km7hp6PyQVH9oNbK64wuQSVu5R9Ro+IjJtBLmT292BAZPpb1Aqso
k5RAlxSDoxLhRq3f4oauOCHUbcdjUYiirnTetCVIpyAIqzwWuVgueHfrYHPVh+J6
Rgwg+K7zXli4TFhH0RgxWCPhYLgXYsV1by0jZkj0r3MahWKYqq8J5i5hTNVquKAF
51nGl6fC+FWkslssrgasgq0kBMm+W6/Ly6/nLePy59wy48FQT9diLsOzqJ17aQsV
5mWB4yiWEx43q33w8LSJqTUAYd07Iqz8AwygDTNz0M/6Jaf1R/NE4Qd2midg2qb6
pmmN5aroYhJ8VAHCckhprdtoE6qZ0Vn5Piv7i2NYDj5DmmMbRNPnPu1j5eZEwek4
MF3viIs7MoxvB6/mOayi0VzRFx6eUZdZQRYt1xopJeSUo7rOgtdr+5CULwN5RDpY
pIdFLejPyYJq3xxBbeTNi6FLfxSy8N/jcufHClmj2ZcYep0EDfcIoCatgc8LiEmC
2SpUQ9S5bQ5AWQLO3JJoLdVdu07gFijRwztFb4Bxd6eWbQjdnUQXAj/4Rj4r9LfK
hZlfzE92ldbnV+I5k4/GKlVz8+z7eNA6q+eAiqUME/247bKwQ1Q1PRM7AvgXsfpg
vci9i3IvHSqPnpvVBdjSg3LnQt/44Qeg2ThliZZ/rqldWnPcJ4aDFTshqEt1tgYJ
/YJSH1k/Uf0nDckveSUVDU9oQBnKHQUutWcXYRsYhjnwdivlDISleYAvWGUeXXDa
Hn7fIMyQVpt9C/QXeG4alz7UmYDOX9d07ySj5cugUmWVr9wL/wIuTErqV73skQ3g
z5ZkWDaScrvCJkySOy6PxgIXLIaHpDDksinc9D0IJLzXbxlUupm9FJXKwCDQ/hnj
W/W6BiuqUBTb38/SebBMxEOvPB8V899/caIUDxjYfccBpeG8u6KR0kXNWzNETL5K
EqalgB1B2MiZkmA1KuSaJ2qf8x1KJ6zubcOO4BbiRhVAPMwPLaFuqsADHBv0zhy4
bdg+DMfaByBSpRSLV6U/uQ6e8q1MuAvy1E8yiIYP6rWspfQfGPcDqE0tE1Z5NLri
FQDgpzutPjn5C2MbfNDD0+8YOCVjtDwK56oVyKATV37stBpAa5AXE1d/yG4YJ4kZ
yaLKBWYCKcmv/sTU5VDFCTXa7HNjdNAeZO/os6CBhZ/wkgSmWKxTlnUPMTl011bL
mN8m2gTkVhbL273KuGbfOcegSLqWA2cRwAPoGh1V74ImEvekR3YbmGfe8LdRKMci
gqjzmXnm8eCKePq8eeIgv1Y51DoQI7IjBE44jSwKb5asb1Ree8fD2yJKMbIJ44XN
Prb964kri5NaTph5/QaJ+x7ljWTdQaZswD488ANgblxFjtNeQSMMWHe4cCfzexRL
v03T0TUQyRL1ApCIvEA7j1xS0RKKX3/UPM3vekFecbnvT7nd98ODwgU2G0qHUhfF
ZeECCXCGqGLlOaip1nWnPHe0MDJPjwfEDDn5Xjv43P5AyTHbyIJ/EL/1ESk04b4k
PSB2m/2MEpO0j9UGzo4Oro0p225cdtvBcwWsjhK3UHM0sW6N31RUD8aZYmTiZlYt
lrK8tiMS1BVXq6coE3faz4TJkKOPbsvSPzisanZoHdAPWYBYjDHn53u3V5GfzhFV
ldbcA0+Aueh2yoMQArvm4De9nMk3MmQqxB4dyzOtrdMHsmgOboKwQz+iRA8W/vaX
jb1AyqdmUOV9+N9rBN36CvO6eZaA6JaHqDXAaqbdxSx1N4nF+Gqa41/0tNZix7Ul
UHQOtU3xoZ9yZaMt03Gs9CRqL2bAnytPEmXWVLA5mazvAihNGckAVhFboD1ZbdAB
OZaPK1qNUYRLbcJhzes7rdDfqFFYETOTd63spLMkUPKBKRCVpiJUTuxUKUFOEoJZ
f5Iq4ulNwG787BbfpIJ69vjcEWg3N8fMgPsPngDdN252NvFY8I9445UP9vRYayoe
b84+AF2l4KmI7BeOOQ+7jLvNuvKpFnK8QsDPjf86l+wM8hIIcgtTN3YprPRuQr5t
nKB5IwPCWo6DYnYBT4OUFytij0BMxFiXSQewR7WtKK1R6/RJvIQnApsd8pxczMd3
o4iCCHV0TtkFTwWhneW3VbyAAEVF99GjL2KIvJFv6h+NSG9VEvhLgMsXAfjqGwPq
EfaFB7BiRD6FGUhTREtXq6vpPq4CgFF/NVOGG/ECUhZasdMLIy5GnxWacM2N/jvj
hUTtSNurRsVZVkQGaMj7zKv3+03ZeBdAv7gK0OrvicayWQuHp+ST6GJ5hxij+ZYq
b++x0zG8UjMcElyfRaLfDTXIYz4z7im5/gsBFznKCTPj05XJmiy7NUtwyjXqsJjW
SiTpe6ynVZ6OBITER2cqoH/I8vaaoeMOrSnWGLCSJlHZnWXv7IoXxvfGeZC5rsBU
uAVlgZHuIMd4cxPWx3D4A41mb8A3A7VTIwgMj9+lKk+TGSgfSkbjcy3rdCFmwO5U
AFY2/Kt242t1yDrDakcTWZTUbF0KN/k7AqvbgZy/g39Wd5gGDdQzH71W5jNlxfvE
x1QDsX5Fp+Iv8Pmd/DiJ82ORoDGmWKqVaxgBOzd8zc6iOwET6uLqgiJ1pskzxmSY
kk08YAAvfQdj/t24EeQNZngan67Wf7hZXp+y+rQcf7lBpJF1GR73vqlxvT9Q8VF4
tvL5zCBVvvRgcwBH/X5GgB77pLX6b/y+Pd85Q9bNXE2uL5s7MUWGwuW7OeAnn0Gh
KYJDs763+maM/Z/Lco5xcV2mIZadMt691uLc2awqbo58TrZNkyenRgSM9tqfLIEc
ty4ma45NP6so8paYRE2z7eUmq1jQE65uxwRGLkm0a/RkfT63ju1wMYq+EtlhprYH
xhUZ9GkGgiUre5ABk/RCDssyFzIeu1ZVoYVPzwbWLXKboh+U8NpDNVpaB/FxzXT0
yxpM0XW2PJzvRJ8Msn3/CBiW5e5KXOZAAc9h7gVNE5VnlWQGpYDXUqfqwrmnEz+E
m29mliHTDWw7rK1POjOB37hO7vwlNQGi/CqA7gdl5dQq2Cucch8ASeLg2acZ1YWC
84XZNAVD6ViBFeG0jUOXH8oi/HoMrtAza5YzLPGcOqpi4aO7OM2GNeHFG5Uf8fgB
bWDmOkXdkH6O3mXZQSyO2tlafndC2aHnUTlL+KOAEJnXe1A59dg2aY7qFfWjhDTb
qQMgt+exuzqynzz2n5ABHk8ptK9UQkoy/bkej6M095kbE3sfcPSpxmox4AufkvOi
y8vZgdX0SwiJr5VF1jtaC1IeAsItkHxOztID5dPg1aPzkeUvR2SAYYd4zGMmTcLo
q9dJYn7fBoDs/6+ojnc7c0YTbGrJWu6H8sjxw8kCdl4C6Yg1+sW+Lcea8RMxqOQt
XBLQBONhZfO5SvlF70x8E30hz1p+DIul5P5mf+Mhrp1JNVZ4TM4cWG7UMMdeLAhE
5Fu/6pU/TcsEmTHioWDJ3JjgFcfUnFmRglhkBwwMc0ioiI+tGVA6QC7xVxJEFD9c
srLacGEhYVgqdIO/Ellj6746RCvunblnZ/PDesuXF0UuTBy9fJSDy56yMd11y9mC
nK04nBxaCyaHZfMS75gqG6sIoDrU4QjUqihfoasN0w0xUaCpAHmz4lzRirw39tW/
uZ7u/mWEj2+3Bnot7bAmwZ2Z50sZu26k3FSuQmev1FXYuJerw1j857wt5GYMfe8F
kXx1QmAv4m1ZUsUJUirUK20e2VTnVXaiT7eMDbxgERVyOnYflb2RTPcxA6U/LwYW
jNOxcMA63LhVWZHQen+wstX9UGEo4NivBKXMvps0vSuuPUUeNVfzzToEt1apSmxI
0SydeAc3Zula95dQY2HcePsuCz5aZnuzf3ibrVKmTWuFMwEwik9Pc3l516zO+qaC
mQcVD1s1oyT9FyZ+i8UBZNOpRpHIyIa7P+iRKw3OdZHLyPpsOP2P9tExs0v2/iOa
7nLQFYCESiba7ccaJYK4QpEHf3PF7+eMrDK+8QHX9GBiHVeYx5ZJDE3BFgWxuQkv
Km0DRZd71h+eC9OoIEelfFjURVcjJItwfYgvWgRR/Bw6ZjVyrVIXRWWJNKvLHvr1
5bf8phTEnFQX7Hkj6yuH3LnU4neAxanSg5sTsiK5twcNXKQwqB79odRoDphHO8KN
6QkRgFO+MOgo9XeTXnukP+/o6OxbSmTyr8CocHXVV1i39g+AoponYJJJ1NfYUS9U
7SqnHMJnSnIJNYPX1EQGMZPdgkcf3IJbXJgDwXdNyLFXbro4+4nCWz2rduNuGrPL
JOAIRsHoS3LMxEGv9Mq3wX0YreaG6ccleLxMixj/j8mCGget01Pj/b9Ac0kfTofR
bBNYp17JJhXY1Xewq/bnzTl+zJN4nkeFpZilSaAzZbv34DR4A21zzFrrETlORV6G
tn1BUdwgqTRDa+x+c/ZmwnzEv7ZqeTV4nurhvyMEwZ5qbEqk8WrjAWqp+DXKWoHR
BLnouwUXs8Nw25m0k62vM8cn9cb4sd9xOEUcItCQSGW1ABu6sSIkIdYZVa4LvznC
d1pradw5Lwdo1oebG6sL/IzhGGODflc0+LNO6tIa/BYxVeSvz76SC5do9Sh7Lrwy
iXA9hK8icaC20MMe3sAS1iCvvOX00iQ2h+tCBsjNSYkxn4u8gXlpp1+GbEWioN4c
qWY/v+bGUG7SoKW+Kcz7I/UucBWqbPit1CKrClgTgRWbLeA4bXc3cTQfAPULgTbP
b+I9hMEbCZsnlnBWBchGxlt7FFENBphwzhVhgiZZqltzpZMF5sA4b1Vt1CAlQox1
DOf+DFaksBhgpqVydCV3am4ggCab1oMOjUxa2X/KHVyg4uYb4PGN3tLL23MJ8CKp
SIRpB2CiOVQvugTn41KBwOe6y1yXdO8ZKHaXq/yZjfN2tX+4YWaB2tazh7YvRBLw
Y9B7CY+G0qaM3JlCYuJLKXATUXBr3zdD+32eZ69Js1TxQC9brOxWmNvKiQaieMwv
C1wQsp0LqbZ3rpmpL0KKej4MzCjp89dxqTGPv25xruTd4wJsuAPnp8oNMleAqpbF
cjjzpcwV2udxlZ8k5wV637ENtmfhJDnQbnKsleoGQkl7qvP1Op5r9XFaN9WGvcWX
fZUxn3vZwX18/oVlWncg+J3/m0CGATIgYDH9gDTEsoVapH6vrmBkjMW8R9T8iLfk
xmhtW76K+xp1i78gASJZNtHTeVjKx7uREbvi5/g0SQt+BkeNmOwFhVJOXZHYEu8R
ig6RHUkvcCJufJHA4VYpjSHlAUzNj6N0SPmtMhG5EOgqXvY/SlmwiIMpmSd9co2H
nOLD4akoXmb7Bp4gqcAnUVBruRBpwXU3qBWlEu0EdxM5MMOu//eOzjtO4CuGJd6Q
11uia6bvOJETowSKf3oUuwnaoOZ/j55+307+KtRnOs00jc10g6kB33JkJED6IZ20
UzGtNiOr8+ZnvjBqbQDfEWKMtgoZtuIm7lyVyAq8ZfjTAM3OpbwWRlIk74voWjIa
64p36csjdV8yyzsOh7woQnfatBtpxr1V/omUFmED3kXPQrteTZb1QPGPAEd+hCPs
RjDcTVsVlXFq0lCVLp+kWe8x5HlHPZ6vwqKgRz0c3rrgdMAO6ieO+n43PveGYPNF
PG3OchS4WU9x2unBW3bEAzR+ZGuqyte1CQ2Yto2RalYuPoS08G5jx9GEJ6+baOXL
DM+NRLxGGJkOkqqsBqJe9s/plXUUF1YkSzIFfx5bjLPKcXxCv02LyJOwssVWqY6d
TIaHFI4QdH5aLCQGS8MKTqxbwoZTikcz9plu/AdeEGuSla6N7d20MVb6Tmeqnvi9
oujQJyi/Yb93c5u//3f8d2q1im39E3VeqLQmuehL0pvu7gx/dKvfzo7cxKN14kLP
7IXKChodUufB0Z85NGr4lqoLOER2ZcL2CYbtmAbR81l9V4Y3hBMpUgK4WLV983Mq
DWNvEJWJEtn3GpO4Y97v/d/dx3cDqSSA+/273PQgDziHXOmvKu3wSwPFfpvdB+GV
cAtnbWHEm9rCOMhnfpO8vNaHyFPBgx2Co7ZOnJh5LkfF00Bwxe43lRihorlzfblA
Gp0nTYKX7+oNz7O+EKmgGdszQqtTzyKzADO5+XKR0GmI7t1pLudLuWm6XE+DVrsY
3qbYobT+lbrSxPn4CK2HOxyamCBS7A588Z3SOHNKjIg4uiuOnW6xk25RfwrCaq5g
Fgxi06T8hJkl/z+p5lgMdef6KfDomGBCm+FkCrGB0+3lAeyd73A80Wn9XhFfnO7W
bucX8D7bBCtwLTnJymIHhPAfyg0HgW3msitIhXIXlf+Mllaoyv0X+kn/M3wLM095
G2C6U1RftHD4hcUi2nP+sRUgiC5q+szmEoDfZEi/ePNUAflJM3eIQ8WCksIfTxSz
956EDReO1PvDysYsgbKFXN1dIlXPpTSin8XjJrP14+Gu0Q9GF3DHtia51lCbXHq4
Jq6T3lNPkpooiKUfygFbeUGh6BQLuCU5BHBtopBwMHXPQEReDV/Yx6Go0REo2GNR
G41yxIAXbcR+XZeVMZO1NBu3MR9u8GM4ckFza/dzovfHxa7sbZhL1XsJc3n7HSx8
1MFKEwVCXrStSfCg2Jc0Qz1CBCFDlGz6IB+OiapIMDHnRQBXF7ZeFegYt8osQlwC
4ZMTePoU+RC4szX8s1yDlrBRrScz4wLwxcNf/yhJWXx7UweW4SPdpgl88gdDyaE2
12+iNOpJOfwJttAJYx6EGfnKqf8cffzI5FEFROhJSmSplrQVII9dKBXM9oLaKcoZ
EMZDiF89nbZrUlgFN0HhKV1T4O7zOX8zoPARVZE3/yW9YgjncAHIFsYuKhK43dCV
GHwMi8GZaI8VYIpYGRPdj4JqCt6UZGzNOJlxVpWBzbrIgtCvRQhMld2ZRZv1wEiO
xVHybn0MZt4h5jYIMb4ORrnX530o8yJO8UP0zzEZbjG60kv9l5CrWo9MLVbRo3Sm
EqHBi+4CdEmd/hwYchkG/Diy8tt/N1AVgg6muA9imKE8RCVnfT3jtfF2qLoh1Twc
Te+C6Go/1o/BvUDVzuVl1qdyz7OpPOmRcznhlZjm4IXniS9yKvZWRdlTndoFFdjH
bOf6H1U4JsOWBxgqMd6pwbVNpbECokK37K37lcPy2GgsD4zexHpKPcNWlFocdNFa
noIWIPPHWKjvVB8d3aUNmyoM1QHsvtTyMGFfL8INcG/0lSHpcEATSn9hnfLjyXav
cs8QmDJu5lXvUNVDGpHV1GJa3lrpW6fkw0R3jkNUkeuXqRYZbn5OF7iPkx1zCEdx
1N0xzu08iuRqYOKoCukkERO6ZtVtjkPO14mWa7Ie9KlimimSYzey8tUQLRfrLpFf
p4h4UgNSeTTZ6Dwu1rGhhWJZZZ8F6AbjbdhhCtG8IPzRupSWOzLY2+IRTDuMKeRU
uYJknj3bQMVRVD5cfIYpLxRMTDoNNCxmqLNAq6uYnwBrDOTNN/J89LdXc/5h9Dxg
sFMDEqE0hueP+0RPdnOzI8L474B1j104ANLG468MTT/2VDoLp6Smzra/RQzufwEB
v9EeNve/cZBAuq2AoLru2I4mAd0n9jr5iXHUS2vaq9Iv0nAOQJQrv/cRrx0abp2+
5HO4gCTi59yKV4+p4/waPIS5HOM2YOBc/paLayj3puDfqs1HwY8Ey62clGTH6oW/
kYSgqHWkngv6mgLfVpKOupJWtT8Hq8pKLbtdRhsdcBLq4xQ3IdyCwf+EZctgnlfp
/Irsg6yr7LJLpmNs/QA1/3BoA54gq2M7y5Nf+a0kBZoADqyOjDvFcQsYepoZqOxu
FqtYjHsksuutBF1EpoxfgHyiQ7P4gkON+iPqXpQ/dvUgHA7mTVjbCPzL3l9rWC1s
drXYs+MpGIcu8Lxor6z35NwavQD2wdikSqWVYa/E9gMlz2tVTPvpDs9Ih57XnLCh
Ov75cSPFCmsTJduqt+53XxmE5Kh/ZSAZXk91Bf1PU60vIyDRy9XrFgaXaghsVhsE
caHM5l0zLYMRhCg3eZ07XjlmGlR86Wq768+eYR4m6sX34CtTAbT5icGyzsRRh+b9
1CWL+UOm53WU7MX/Sbnr7xhHgIK8RQAMXJbepQgPHTprMXZHWDvvIouDoGqPHCmd
lYYAhBd7bRhz0MekokVaC8kiSjvmj5p1Vy+1D898Ljn8DcvEnlcf8fSJ4rDYz0ll
mke3zzteA8/UH5Y+dIq1wpXsKVGoufyMPdtI+ikfmqyCUUpp/rEW7PIpl5sREZKy
qHi/pqHT986SKMiedxuny4LO9dQMdlYf3aEK0ZsnI4C/XPIUR7GK3Vis3+CZXyqd
BQHDc27LJn9wtZBgm58QcQuuZwFJJiIN5Wa8qFThcAA6gJ3uAYyU0x1wbI6qQOey
PAHMBMSD1sZupxG04IHv5UKFEX4uPY4eT917fnHWxl0byAt+mrV7MSqr+zkF5UwM
EUwA5nvR/rZdqqgFxSqnF3RCJ3r8RO1l5fmhqm3+5G8eM/8XL09NWcaZvq2BjcRn
lhYwmFdKmMISJ0E2oHY/coAvIO5dvmVN7zTNomO6fuWqcxQPtkHs43gRSzmc42L5
pqdS08ruTUeJtUsSfIhzKuvSsD1xcJ6XsWNKFEQ4b19BA+9aaJ3LkgnK8H8iyZNq
7HKae1VfeZmK8QajpZ+dQxT62xyvAtZzSY796BVyp2/xai8gH54GHfNsH3bRAC4X
5N84zWaUgh4+rDEgBLMNPtxkLqO99Gp6p1gwR/8nBH8l14tI7+wERZTeTdmZB+8d
WvWBk5wQ1/Zz1vs/dUVLPZ3UfKMFxn0e/iQYULjDTJ5fAk+dQKKDXbTi0ScV8u1U
u6E4OmRSB9BB7YMlJZF0RT4y90NpWoXu5Y1ZF0t3kFJv06VNuLigbenDGtCre0x8
/AzzvQWejEhXawCsbVjdd94PaAQEx8moKM6Dxbh7kOqwdYYZX03DXBa1iGnzJezP
ByxeNT4SJabIZPxIH0CG31T7IyFpaGv2dwouXTDxXkcnNOAE7dcRFmf83Wzlvylk
m9iBxbKFQ+EMME6SJvDx8lK99gXO86XxX3RHyWBkT5KSMVNkoE+IYiKm27ZsyytE
LYF/7dis762w/zkLfSUElXJI0+7Yu0pBjlPGM5BX4md/dRLX9ZHBYJjJq4VzLbU2
MRT7NGO3SKpKZXXntJT9AeKmEiYyuCylKZAftZ1QzO9eulCHQxUAl78xOuk61Rcv
2zIuJSJbMd2B/PSreKr8369w59KaSHdyvrSPF7dxrPfSei0Lf2vL/Pf4NvgSQlQ/
tX7wu3AnNufBqAXHDkr4RvYCE7FmWeyKR90R1V6xOOSsg0U1o4ZyOrgEOVTdBMkZ
g8xPBKi9OdJ2viZ9/2thfCYrbUrcrCyXHGEK2qXIFG7G/orwcWab/aEuqRBmWUU1
qWqhaDAA8ZRpkuclGT9CnxOPcG5zDmPI6zxsLBw7KbW0jQ4kxVFHDXkxj4EhvsFe
ry/RD4DL/+bmBY4Z+awF/dH5hjz0DIx/Ng24caBt0I6vzV98RJi1//5V9Gp9b1WR
wQagFuFSszwgRIMnbhBuss9vt/KgdJYm8m2JNBT9Navjh5brhegSo/aRyKAi4VKQ
sP/cwObExtU0ZikBCqkFufJFlVOFoEMOXpM9BUY609ZdvEnkM/3aCa87rcgPPpcW
OpWeJf1r8BfC22OCPfM4MCCPLQLHGAWXfUbVq6+QQZb6ukxPjRATyh+Fkgkr2yCP
7RGjRp3RRS89XizQrL8/vhQ0X/FFtzvsBod4MP7k1f6/JBn9l9f8Xv1eKSd/ktcK
1LWxwe2m824LFv1JJH/pYH1WCCp0wROO2qu5izlIfPk7s49r5wcwfzjYQratzNLy
Juqsm1SOrNwYgMCsdZdsBqfCz8u89i0ylclciBbWmqNVlmbkEYvKSsKznvuLa6zc
o3sUPHLyUOEGHo9kvHEarP5bjoe0iAglLIjxllS1WJEy5ll2e8/+kj0gKgWukwJ/
cqQzyuYeZJZv0tlAsRMTLBeiM3tBwrCwUUhA5cechha5NGLO4MKuHaRFBo6xHzJz
ruGWu1d4MXruGu4Ri1Y6u++1iDks6Iky580zxIRTEtROUs6wDm9VVLqlMdwxg4Fr
LON4e3RJZtMEDzyvqHrRl8x8TgMW92X/IKRwc8p370IES0Il7cK/yB23gTo7fmZK
2lXF5NbYavgkfyBWriIw7NrWPC7AdXpm4KDmf3FqpkjtwWX3597Sd0ymzICVuLlv
k70y08mn9DcOHso5uMYoIXX/v+T8Cdy3aHSNPmgjS5qVxmibQzqvBAh33FEibG8t
A11l79TveBwWZL1fbG4FbeeRpsQa9vHMnrOSFS5cG5RAEBgIbZb+9uHg9GupaR/c
6WgpJYdEQyD31fSB1A64juW/VszYtq09up5B09+LSw1JEh3/qFoy2zgqLBNqStwm
UPeZEmMd+KvI6gPQqgRHVOLq45jrNNNwVQMiazF76HPBHiOaQubihNQmAOcv7Ddw
hkCMy2NPGXUcGExX+YhtN2wJSrecN8RUggRMFThoK9MeJX8THKOuVwtNjNbpmmt9
Bfx8EbDUYs7lBWD1KYuiJ1NRo2puF9Qdh2qbVz9Qycv3WOXBS4QT9Six2Wx7TeQk
17rbPt75CYU85w5RutThQHNNctb40GE8kta1JhdP4weYKTeGe5YUJ8f4QHk4d5F8
gXIbpRg/l3CQ4yb8HP+atkzzkzDLyhUVE8wQxpTv45zwmlS1WwXaXam/8Lr0k/nM
w24XmDXu26cZSM46Ks4A8pHgpEI3hVZvX64BfS+fzNj0nU0pO0kIXXH+y4TCT1ms
L6j0WTbHkcFEBzXO6WSMU4qLPIISMJHh/bwgcKceRYgJdIYMefIFji7asVpsvCO4
pIgA5mr+/coMX+itYp/c7gKkYYanzNEBA3/qd7EhdNN/oc3AkS4ASJz0aZDOTMg+
qhVDYvFrGwXVV7xS3yeE1S1CM5CQ31qa5eeo0ZYUb1XU3zdW1M04v13txFe8FaoZ
/GVmvIJ/gI/0VLugVh+cRdFjJDSLaqt+RWYLBjIyFH/Ys+HGTkfuXepel91RhcVX
+UexbZthgyTQlrhjYQ3HWx7JWPWG+5pQhm3eriBITkjOM3H8xvck/GO8PaqKNR8X
reHsRUB80C2kYE92ny5grnTpkPbK7mXVD72LVioc5k7VYdamFjJSW0T5PdquOtsK
MV8pEcngmvSgTFcBjbUmiPe5B9JF4tty3NykNN12dQAE4xM16V+LrX+nPQST4Fu8
Bz3jQRYKK9bI27Uigv60T9KJHi2h6PLVMAUgoAkKo124iP2qU21oYA+jNs7XyBec
/cTnQk8mBxJMUWkj8sUKHMtMxBgJSYu5wrvj/D82gMd1/GT93RqtnJIBJUFXpNfh
l2sCCReVEBqfShiq0gYADWN97QTkYlrO+/WLyKvdO54xB22PUSycp5o8FsYcOSzr
m7PYOfrQB6CwanCr20zI72TSr2YAhW85kwpM0CkeozEadmpGNhN/GvH9ggt1Pxwj
4fCgjAviNzeM7W54erEt3VlRsyysVjtTCm2PusjI8Rf5p9kjeTKa+YCfxCRz02c1
qAn667iRBcX8nzDcUktqpbO6GuocrsqsD7AAp4RNMxbfIo4wOdaaD8Nwz//+RR8o
CKhyAb4rpnn6C9pIz6Ql5n6IwkhBzBZARw9R2X+rWho1PiopF5snuRByiCWOZcM6
kGsOS2SmA0xwdqrVOENK12x/xlIcJyfF6MBXHWgMeeh9FZTuK8ZGY/0SJ+YZKcl9
RrpjnXWUMP+1B2+lHa60Dbo92FflJtWyu89KNTdD9bnGxYHQ7Z5RNJVseaSIM/rK
geDW+eqdz6GZwnP8gbm/tnqzGi5VxL+b4wZeSdf8xQfhr9l2mmAjvCEjF0ovrvQ/
kPGC6yIGYALCFU+iX5rrdrfIvnSvhtIWY5FNeFBLf6iUJinz4njSzixWsBpU59K6
9LnSstpv9rhWpeiNG4bA5vnPJTCHkSZiC8ZjBSAtomGhAWTgncSGFK8C9KePph4Q
1HITGm63sxN3LrzzPq81L9EVKfp2GCewIzft9gnd9mqsbuezhiqeQ6B4DKWLfACf
thffCr9ZFljfsQJmoCJj+cF3t/EHWqfrRsoTpFDsuG0DVAL6POZBnMZueT9YRRN1
dgj4eqQPQk0+e3qEO2aQkfkyxEkqxFsT2FK9cfdTvvL6lyyoXoBv1Y3/+DLaj6dM
sY/a8UZ4P6s3ki4Viv6SEgWRFO9/E6ug1WceHkCJqGfybbACdXZ9YxMliIdRf98f
pzygzklTU+Htsk2C1h15QtsUQyOkIu8xh1hmYQhmcsNXEdq4zPei6O46o/19MlYF
4qA8MmuXJTj8GF3UQ1hCITUUvv6N3KTpYaLRSNEl0G+NM4atSU9MIqAh3e4/jnm7
JCyiBjOVlzoXVUJXGPqZ2dy+sqvx0Fpaq0diM/cQFsJya6z5KVxNIdR4pX4P/yTt
2qiscZr1XHsaWIktMbteSfW6MDu5ECYPfhOkwtJpd4tXIzpmHB6an8R40QsW8tJ4
0nH9nAqIAS0pFRpbsLztA4fGfPNA3E32nahdgNjtE7o5n3z0YcGLGd7hekuVdyzq
Upb8X5Os7nUZTzwAyOIoijNjZqiy4N2fWRm4O2BbT2q+onDMEMHYE03095UPayo6
s2DOtmksDyTecWi2Lpy03eqI7Us4oliTUL9a/tXKLimaK+EFCpRN+YIT7CvcGdHs
A8RYL6x7mi0o5sevh399pLGDbhf/9h/Ip5fu0ORAd6Uqb6aW8OFTJZjWPuXmPhHy
zy44/o3QQPTewSJF6oHOxURG8dMRgHu7tWBhUIePtvzxbEJAMjCs3Lq4Z5FCqo89
mpjPez3cE//azROdZTzLIHW/t3TAP7TK4T/0HXPz8FjngP5SFkLW1yf7e26YaNz4
YBboB8ouIP1wNFfRnrFu88J8CWT/9J5ap/N/jclw0zay/0ukgVGRnyVlTlg5DeB2
JsPC62r+MqBUF8OIPmlRYY4iIDeu+qCu5YlH2QSw+NpMKJWKWJKY9c2yE8izgFgL
MWDaTUApzMfX6yCvk0oYEilxS/9Vduf4T3RQ6q8joWbDK69X5LBRSqgKaPtJ3tNC
AP4nbHc4Ykx4AI1FDh/1DIjxydgnHDEwVeBDjbdf0l84+t9QbalzG8Kvtl8+HTAv
CpPewtRfRh8jy0YKT9D2t0Dp+R0143XlT0BIeNR+fQPkuJUi2keCDnQX71G8tb/m
ClYUdAykRxKgJqOe17JSLb6ivp/g3+yFnuuE3fbAoiyUqphPmCVW0+YClSxcn4t9
dnt6IymTX+W5WMTj/GkdpYtlkqZzUxJSNhDe/4H3U9cExNamlTDauN0r9dKSwePX
e8kbe0VZ77OhjMtjaMeHsR2YQ8U5OdRYHOMsgE2AY0pYt2KyZhvwlPfbPUnhyyzL
PNHyGR0Q68LUmPEqOTFDCAEjcWWpQioa7kwwi7LXp+9tyh8x6E/MR3+m1gdCIeDP
YGSG8ZhmTwd+EaopLFu9O7p0agDGNgD+8nWJIKr5RXpJ9i9hxUKEN1HX9EmkhwQS
UJN+JVYj7zgipx3KgKkxvlLPvUYyhoK4f4jmfVm73nedusIuxKkHOo6KQwK2jMXp
H1WdJ0m5zWcAzuVrcOk+N/D2a9bMx4YTLjL+uHdANmCfGjYUmdoSE+TY3rIOL4X8
sA8e6+e/VMJFrbctwlr0LjF0Ptc4gC9CR/ouVIBHV8KqiP52BRMxTOi0uge07YQl
lS6CZsYrMe7RplD9QzxWuBQ8DMh+FkF7EHrcfxOYhe47m9gCpJNPVnu1p4L6ZaIh
SAqz6CqcAdWjrEotECesPSfbphutSfGSH8LWVKEw/rcXKi6e+jQe7MgZjWmBNXvt
Lfkc969XEH4MkKad3QcbkjP43bxpIc/PZetd8+g9fF9ZdGlx/5wpheDHQPB4VKZY
/NsV/EmAQvNZC/a2GBWPmJAIeZKoh1mRYbXaDfb1qds5rlrMQVQ/OzNts6UWVRp+
6qe91kyk2pG1ZQrinGXsh4xX4XPoGQ5+poa0QqtYzcbkuANJ/LCo8rbHgnlnHnB4
RppS+UiFCLDcXql8beY5Ow+TUfhoQDMPhV/eookj4E37ZmCIrYJYV0OsGq7h1M8q
nkVh6OXF9Tjh9PjMdCRCpdhoyIP1JwmkLmcgVbsehFl6CsXmrp+twDSns4YLjs+2
LpachtB85s/Pj+sGizGPDxV04CrF7UV4zOL2cu9aJZk9lLAwpljJExgYKVbVsjYA
4LdnIvMGCx+r/98aJBp+tjVEUth37l73rliPe+4c6rRAVKI3kr9IGXuIF7AaryIs
3euTDZ+VxzzbeZE2iiSDi8miHyx+QaPmqfUl5D8GwLXPQPCwhdyu8Vj2UHQT/oEj
CgQ5W6y8gW2fQk/5plrLHA1MR1CvW+mHn7NUhqQFrZXHznmtBO/DoDIFUoHd+m0R
Psg6D9UdEYDgTcNivcymajXNzPOhJbsjdXed+xVyk4coIXG4xvXrn+k+kdgLRuzX
ylaz4Wav85L7LVI+kKFY98QGgeIumdwhXLTXb8LCX5tALp8r+xPBZ9ghJCLwfdTr
r9qrYB1VrQbaM8BeteGj7XOOtLmAia2sSkxNH69ms9ySf8HAT+RnEE4Wg1Xr8QfH
iaXMxIm9qqgX/uAHc2XkO1f1mBZQuuYqJX334kR5Vycr1UaJ1dWo+CP78Iz7T6os
50+2C7SPiyog9i8Q7FjuRA/MKUeDbXk5ej6Jq2J/HbdP1UEQsIqdGlBROE68qipJ
s1pbFaFPvZRp8K9DIahSS1cpuLShW6ND8l4ELSuutx/70kYLCqlozDDH4JZLtDq8
mBEoQ7wA01ZpGV/gg9n1Aet0A2BXlIMw+PiPKbJLUrSfWMAk950aRekEon3o9t0L
9bI73O46XdGFUeY+ge4CPhSnyfDMdK9Q85o1pIrb2K3aZCeHaMLLH0q1y5Q05ViM
2dVhDJSQQeqraq4kJTyPZovLIV4huFZc1+xs6/NGFPQNVHGVvM+w6S9KLvSTd7Yl
ZNbN1e3WIzgfFeFwHrhLH7mZS1/AUemfDd+ObpWH2XHXBvJe3IB3uC5jXGx6UyJ4
kjZ/o1YQpqV68jJO62e7odezefirvf8r5p4GuMWqBEHyOAjCH4EN408lUrQyphCG
SKnHWKWvF8g6NU6EQUbou9/v/pWHz05qxOsjMsvNV4/MkoiLZPEQQZQ+YEcRCFyF
baB8iqiBN7S0bARQwVvhzLpgMKwWrVSB46tU1WKCmNA0VtiPi37Wosa/11Vaw3sG
56/VW+99QBuVAwII3gwePjhyzr4RZ/SJQ3ashS1qzl61VdmAnJJ443AwOox6BfmP
bxxm02qpXdpfd8ikvAKEL5R0vRvgwFIbdajn0Vv3ZUcv8S+2AivT+5WmUjNkM58s
1rrAJEmhPycd18Zkq7Q8gCuN2g/s+Z8gafmIXX4z1oDlctOYzvFJ4un2MNkKg4L6
UwtIhGlph3gEzO9sbmo67yy04dRadoeN8aGplWO+j92qxeu6pB2EBa95t/vQNMFH
u/1r+Gy18lfBex6rGBYjVLOQ0HOjZ6Wm3Ax3tvmjQHDBlbYGt4rPPNJNk6YojEjF
wtpRsNFzqn/h7OK9/FYnOT2IFnT6YlnKL1R+M618LvRP5iTxNHNGCxgYiaVzwu+M
5zTGkpN5lNI+/l6Ns6wvax2zlilWE28RiLLdXN8nmaL3Y3v79vjBesW7ubNhY0VB
/c0J0Xd9CeqRvcePR0IbPdK04apozlfYLhWRe6dTl6tAwD7gdhuVb2DzUBRDJ9TG
NFWXKWYXtAndspLLKnfmVtia2HfksyzLaNS76su3EXPr6vSZXgwsmtzx6Tvb7oYb
6FK/prLHQLrDv6QSDl8h99oXkExceZjgCooYQjCiOqgqFKfmlTLRR9mmFiU0YHkA
AV0T0Vv+DgUvlcUzdlYgKhQ+Rbq//C+9jFb14/ypwkxU+cWd0biBr/sJQJ2E7o6m
AL8WxWNDyBmnFQu5YzKsEqRvciSt2fn1gTpZkqDKxSoeqDdPqs4KZkq6LBWM5Nw+
EinokF8XrdXngBp4+aqdtOvCHnwpXOrCvtnveZ/tlF8ba5lHvSgtLNe02uI2LmEl
4vUmdS+zwJyBdew5h8cfIdXrl+xFHn/1vl3gTB0jbsskILpQOH5vN/sLEibcABod
JF3Jvw30lmjSeJMFEGR0Q1petb/gH3O90SXMjQC/PLvpDPT4PuC6BQAMzGgkFilE
4Ejzobgk/7JlqzoNN0iXY67a6mj5cBRqd1wtmuN+X7HTrRYslh10sth6D4amhfeK
19oCNzoit4hw+EJhViwmr1p+SLK8l7WQ1fJk4Z1fJUggxSutpC0SP3LHSRa4hOHs
Wa0JWMue5EQnQlGCxqQ6IdqTrVydDc9EK1zpWmxHOhB6IebIvFwGjrEYVxtl6enO
oIu61G5MzHGz0S5LB6U8TpRCB6xbcZfuPWBYOiMzcb3pZz9PXy2CJ925tp+wfQAu
UvFGa4h1UIgbNu/hFx56d4La3Mq02Sfz/W2luJgdee3KgEC6RxP3/iZZ0QYrq7U3
ossQXZ1Pjdj4oBevAUW5vyYjXO3TRllzUMjIyIRkqJiADLoVhJEKSmSF8vzTsAYs
oK24sW3iM0KfSwhmtVbgEdTofVI44OAmCBo7ayuht+RDGiOadhqi+PoUnuTojtaK
JnEWbCI0/SVKhgjokdQCdW6KLdyr/E4PzxwZyxLLpXGSapmHmeOtDj0ldDrEztYY
3LG+nzSCQ4hDYjpALVr90PNI1eQ8cd4pGaTWUNVpHnV7LUyDI5nLVsCGpPt8/qJ+
44WkvjjqjB17F2PCEyJ21qahSBnqvG+to9qP8ox8PN/bcLlz5XgdKaLMjstZjo+i
nDX+rdtUOyVFo2yi+pPz6teHZXXutLKhXX3rEUWpudzq4pafJeONr0WJ1Fms5JIs
bTIwGr40K6gNb6WJkmzmp/fykRyxxnUXMX1NTQzQuqzE3Ggpg+Qrh9ev2NcVWzci
z7wbF8FEvUTK7ZT0cdF31Ysdjm2mVvmV8/xTS0JvEiKv6qBdIy7gHJbwXrqyv/Fc
0/OYBapYRIamnlzdi5jpvwr7l+TjDb7LYS1ZJaFuSiiTpJS8ksjvblwTG3OnmZ24
BcWvfiviSuDrM2ZfDIFQ5Mu0fMePPgrnEtUae4/jqIobosMIbNhhOBHwfgu8RTC9
z7GgcMJgSIaTD6BaU90NLGF8u43CbHm/86ITy6sEcuIqYlE+BlKT01Pf7Wd43u4L
J/l8GZYrrHcoEyR+yD2yesowv75NuXqQrSItGwTci93nzOfMD1svpn93ttTtM+fy
yV6SX3GyI+xaRnsw/c9wLIi6ewGyy6DG0ktEiXmc4twtknCnn5VT18cU12QZ/S0m
OuRYTSailYAdyXU+79L3EjxsWIDPcW1KKqw/XFNcJ+ijzV+42oNMlIUUmUhYGnaR
QTHFpoM7mDtLnjHPD4pX8z8wArPpxcWAuZJX/yHjBaAke4LEA9NOQpP0SuR4y4nZ
fW9GC82DKmlPgB8vCFfaBJaSCxonulHU+xpgHwNQo/sYmNQTRYIxKMO5k9FcQy63
inNdKp9gFbLPkw360CmmXLjqRxhAGLipFOM4EkLyLqIVVd4RMx9MCXiqx/2VzOLM
6vvcZrHibJbLdWw5IZd4V2HXKhk4ljB3g9Rpl+eIDLMsrpROa1bguZgkSf5fAohS
BlnSKuNPA6Lh0bofugY0f+SGxc3pEpFdSeskvWcjktzbBBIvyEuPimqEEk4LF4rz
XOgIKfGk47GOf9zHsU7gUyExcp5br7txj5duLPKoExlv/goS4NBMQ8YHR3N2mXFB
iUi6VVxyTaonojsArieXPfTmPcUySSg5qKXSvR0NWPYLbFopChTglCztOm0w8HAX
USPrao5CCLVvyo1kmNW1saxdhsctDAxpzZPLlc4uI1MxeT9o1r8+Y0+VvfmfLPGk
QhtHpsYP36RtEkks19cVc0BHmJIJUCgJ9RpBLMpHHM0bQx60NoYjfGpoG4Y5It/S
s033i0QjB8YNTHuaE5udpW5yCFuCbzACyQEI6pee1btHT82oV8ICyLJRKZGPQFWQ
IXpPsmkLSESjFI6a08vO6+RCjBeLvOSTljxC8xsejaqARL9mlhPYyYG4Fu99lqt3
JWWRke0NJEtigfNHtqJ/Lhf3deUUCYf4/U+lmnub4ArX1mZoo2qde+mXdrRLjvh1
ojppVPVL9LDtY4gS6YLibiDBT2wdB85q4+AqrE6r7xsrz5rTLPU4PyZooEYRRahg
cTEoVk9+23dZV4kTFI43f4Dgmq/zw0lfQ5cUhluzidKSO3/R9gjD5nF/PrAJ/Adc
Q5shyq/VpURRR9VoH4HZx4DL4R7YwhFalirEIOOGDEYdGKjYiA/IAYI/m0xaR6FB
dYXtkiPQN7Nq8qlV3W6pAWGFYqu9qra3mhkRmwMWPaAuWA8EEnWP/GvsRK2qki7j
Qn5EHO00Q1ascz/v5t9LqE3sfu2D6GKuT+GsAUFu8kFWFq0HoHo9dDRIY0W5mSv5
YwQvxadyTb0xA90PkUU8sKCCl1X9B6ulMfWftfN2/Hpfqh1myGtA1Cf/NjotZpsg
rxFjX/1TB5F6SBgko0X1dgiki+rHk37JHJWMynG203L8N94BN2OOpKL1DWP/QyPx
nSYXlGomxow/II2Khaefz9YQGFQjjRxKnDfMExuXsF+byUOFOKO1jBA155/Vb8a+
Y8bTBcVb6lBtcrxzWfEJcBbqnY9pGHhI+qAmfbK+YWKtkOWxHAuMaQGm+DTb3vre
ReTS2yxRL/3AkuKndk6RZw7lesJq31bTKDXRwr/qHn0d7jbvk9vlRzDUbqRnol6a
3lctg3Soj+PYpjESHm5T/Ll9Nqvr83LQ8h3jMXNKzjLjHE72o8A+bqJODLYwJcsZ
mebZ48sPqOXJyg+hb2HYvmSm7TEZBF0pQ1wa0b8glCpWQcTP+KtV8kkkYa3p+Ilg
3dX13E9QgckL/SOf5LGobOiCJUeBUntx4zI6usA+CfRhNbDxXdJWjLBmZPMXH1QK
DLm4oejGrJ1R/ast8gVNeejY7uKrJ+imwEBHu8y+TB8vSrD65mj0nLzFrN/vbLh6
0UNUkBPcQC1ex+ZDo3RECR9XmWOaIgusNBRi7oepnIc6Z0mroaQmhrkGklZo9TmB
vNm2zgw90It/4sQmN47PIPugTc7v8WdX78KWYa7x758szaShbLN1hXmo0ycuLoUI
4lzgKLYHXi/lrOJ5P5PRRTLvbnwoHbdWzcwxQDgHlDKydwIDdfO6Tehp15U5Hsg6
8kzpOjae9FRncA6jHRwlFEZVX04FovkCROhPOFfQxkce0eOwWcye0R8TXGbCrAaW
xvA7stWIm0kidVcXCNLDX/apv+kHpiauQa/xRunzvsacffOPUk4KvzO2RuDcP+d5
9cjkwGIzVWqBoOUpzHrTMox61ImnEoIDLUfstLfYBT56yAkoiV9Q3g+IbaOd8/EH
pEoZGx3POXrdqHtid4yKzsZDAhLrgVqjRl6+yPMhG79ljU1HBUcH1uefpsX9giJO
H5VAUTu3Z2d+XqDCYiFCoTe+qjVvP0l2mgAEKhZCMqgRRJf4oziqGm4RdWNqPIEz
WZSQIf5FouSii3CjbxXY1EEmZ423iIG3rbyaVX20ovUZWdT8x3xEA8iB7OCUyJye
qC6AiiZWE/hmWxtt/ffPXqaNZGpr1b0hKZZlyWJUrpSRbhVWwFBLPHEEg97I0o5j
n8klvr2Xw4R98omsTNxkTb2mH6PbKlhGD9xkus+xL2YqTQj4KZVfcgnbCIKNKhkp
eVE5dUcKPZxEjmHn9N3OktNkm4afmMV8lTlGkIAJQAQohmqTN9pNZ81UoPrm8Hxj
RslcTsU0RN5sciRZZWgRa+sNSWhND+ZyYrlk0rz+NHoA9x1SV36eXwc1j5k/gmKz
mm7ZQMApABRMhli2GIe/w9oQT/lcGUBVVMVBLvHe2n3scVtByQL+MtgfxdHCynLi
vER1oR3fdZNGVkVSzCZ8l+1S2Iw7vlVMjaNmCzQhKT/ozdBthulLc/2dZz1e+w8r
2O7zvG5vwZTOUu4yKeo7y24zAooIImyknetaV22n434Wa5qwEoM1HM4VngO06Wuh
PqKHoSek2Dy9KjNcGAHyAZDAQ/tiWwOpU8vCdFhZJLi/ExTqMl7Kn6Nzk4hW+vw7
H8CzoRrrT283QEObDWupi06UX+P+uxm4oYWXeSHtZlKva85v4jWlEe7gjV1TSZXt
HEsErHSb5Bm3zMRfeBLHpM8oYW5C6LU/uuymXgZb5KP/I73/riNKlv04/qiNJrSH
xVzcxaFJnDRg7hXOT5FxRXtRykaKl+NO41tov1Sts/0S7B6oF7yC0V2NFUHygN2F
Aq3806tYaR9YA68OeYcNQpjqFurP8EsgOAmvSjp7OTmaRNQj0yI7sRn5egzGWVhO
zDNT2GU0Gz/ODA86P3FvhvcQKzQLF5oKsE8Vh8/zewXGcAn2MY939t1fh5i+B51m
qZiW7f49iHusxdViZmqkvsqD7wcevIeHVZ5aQ0A/Hm+bcEUupUNonYxQoucgfQpa
vOk8KwGKJ8tceK9o7MR9naCEOGHk1rQy3aNbzKHPUTTZsIkG7pZLua1VuuQpEX3z
D2J93Cyd6QIjHfYIVJN6g8SOkQb5TeOcpkfxcn6SSqAnYO1VgyAOwafdIbcWHgIT
wdvtKJKb6OuMy8v2+jGAAK9MCtLouxBJA9FKDSslqrAMF+si2Pca3/sqWt5vtV0N
fW18161sBVnnX26WLXlwzFsB4AiGeyzbXDXUTyC0jCs7xvw40427++G2nhhqiko1
XxSGe+jTB0YUjS1xNaFWHDb5FFcRcu5AxQo/LTlXrPkvd/QjeHI3P78FnBhheFF7
08CICCND13utW2mYjc+n4T3jUHKkCIz5947mVxkPG7jNV+XBjrDhBtqrC4C63EoA
F1qATAibU5tysDykORaxhFyFH3UeyYcTUUuY//Cjhmor38KevumXiWWLJTcFelDl
f+lFy+E7KZbD9pCrA0RtpRDZL4FZ3MamPAS+N28BwLPeu/bBLztUTSPUNefYeEIl
j1ZNY4xYzK5wCcKdZlBtNLUU7UJC+/Mmy3086/uABIqo+DOYdtUi8Ck5hcBSfrIU
TJ10PbLN8lWjYqp4JV/IwHHYA2BGzCfpvgN3qidRurCxq3BY5PHQiuB6oQrm8GxA
ohSn/KHGC1lgBqxC6A7x75y9GA1pq97bbs78I8ukgxn8bFqfcQC7uwHCX0OSTdQW
+pVZzNKN8ABkPCCPZcjTeKiH7/xG6LivIwt6f3xM2I/PzrrqY737Jq6SGMWzwmaZ
cBeHo1+W+xgZkQZCykdzmw/YY04lj6ljVsN8XjTxjVk3etwJIUirxf1oqgCogva3
IPBOaywmb9wmmzF+9ZTRsfu4AvijdKuRpBnwLfszt2qx9Q4q5EP0kOec4Nwilrn9
2weVmdRZaVm0o8RCG7y3UnPVerjTruSYIm2rwgVsWumSCZLqBw+Y8ltUlvEkj2xf
H/KFFEFogO4yxoe+CxkRO/5FgdalDmZwP93C7l9refiOdAzcKdhYD0uLgnL2bI4N
Fdbt0GP4VWpWEzbwH+PAiT5Awaq+69suC1ow1Rqul+Ab0f7M38AvI1RTf1uimQ71
IRRfrwb3aj0OLuW8TpU+4dWVUWHvMmighJ6kQhUXmCWgXrrvAZCBADC1re0GuCmO
pzYU87so/iQj5P58t/WeSVPowkWftpkvk262BddbsPb48xNo3RWMEUDChHgUy6WC
H/fbi29ioZs3UOlVSzz7FlWyUfssrq69gsfCEWIApOpHuNZ9G1hrZScf8CMSziW+
m406BU4oPUHZzrTzs4eDDfrYAjaz24W4Rc22unDQ1EmgF76zW2ZOfibbL9JbVhF6
8yx3VSoWL/WRjB/8cmcVB7ZfnrN8/mJ3ShRn2FmBItGcrKElwqmKZOtIWR+ZzLjS
KPdn44HrndIZrKh6wg4s4kmXlOvpWfPN1C0no3ljp+6qpWhkjxKL7MbDXE1QtEg0
cZznbOQS2YZurbdWN09GSFYElaRox3tR4ydNLMqcvb69NVywqVY8s1Tl1eTcllXY
k2qD/syMtm4XR4Iq+yKNmdQZSzyWXKPyWjMu7MTtUG3tNY7WGwQcNc+JTi98BgXE
wlhN/yxV0mEs42u4Z3+2BrBPXViPB2z6OKssUDMcJirfK25QK3Z72FJanotbzSye
yt7I3RE087K2Cki4+TmsiFHGMBGbj0+MYXFY0awA5neuVwSFKx/iXpPJqQQPp6rU
cqYuelHo7Sjb4xOgXz7hQfGpL3VOVjg/V70FiYMeR6wCUoEjV+w1IUgz4kZ0URaZ
HfXKk6e9ShZCgD+6Hn1vlhfVrdNIPRcikOfjqURAKdsyUZVvVn2IuAhVgRMlmVvP
JpHvdIiJsI5A0TF8wHZ+DyXfp+iUBN3dWp5I5Yh8i2PgPVDsXs1Dg+NUPT5bNr0r
Ng9G1qIeotSZb8GARhzVnXk4t4fhZgzs9mCYYAvn8pSGtAjAi53hXO3/Af32yjbW
dA0d3Itd4lfOd4gpKRj1Ab1cOxXo0bgSGJmm7gJAFDf1gyoubdCTa6qVFMvVISTS
jqF5+lXNDjvaErvMyEUXdyfwB0qZkouqF/znBpQof5YqX+ab2g403EDo02hnIKVb
lNeHLmwAMJ2oJbeoNvhy2BPFkifWIo9U6iaVu1Zz9ERbtx+BWBONqLZLx2hvThak
2bwXCIjuU0nj+jJ+6AA0eorzDAMnM+0hLqpCf9y936s+Z8FDV0IjAkSYGd+D2ETu
rjDurHd68O2Mb/eWI/ChskB/z9XPkMP3q+46Z6zm6+3CU4Z4OMFmqSDEGz80cmn0
Pt/3AxTCxx2Dsi987Gxx4weDEDiwdNB0bTbjXcc3YLF0Qb8Pf02xExHAaw3en/7U
KW4G8Rd5DWB0xGGaWoDt0cgnd0I9I6Nd0IDAT7akD6ptzDRNUcNkQ6lWpyrbodGo
sggY4lPoa4sImTyMWopTj7MN6RZY3vAy5VvjPR6Ne9lV3qkAi7bjy1fezf9Enj2c
UeAkBFk9Sb/0av6VO8XVPPeajW66P/BnPBztXKnjm+rA66MBYDzDjKT1h0GcHXNR
AmiFxiReDhPRIWKWiBH4lPD3GXwlepmOPnPoBlkzGiPnuzEsxzErNWbIkvz/fJvM
eMUgIYeCfPLS2tPZmefbNTlL6U/x3DVeD9onPC7iSPefSceIkontHFt6IafAtlgf
E9yEH29lqhjmzV/sfhDttZKOvwuuq2nrn8s1/gX1P+CMlYboUFvVuicwTS0m3G9a
PMZJecY08qfgrIp7qkZTOhGdWwTNSVEPR7x/Ym0C4EKZD0cMYm1LR2LIgxDhBnH9
zCMWYt4H92dp4FYt6M8XjVfrfp4x7akdzMKEJSzrudVRMk3d7WTcqFOhn7XBCikp
bmOJES6uMfA0nwO7U9ufbldrwT6MzH5D9+tb+paX75Kyi01OVpTISzZQlfGGTz7i
KcUwELDg+9Ex6xiaKZIMF2G6r7dkz0OPJkuXopWVp14n96/m554pyAiRYvagvzNE
2KzUs1eaAFRlp1cwnbPuvZ5WNb1opxFHmVQ7QmWWn6Du15aiXBKnCdeX2NHPzsGX
HgNRlGwYaj9EQlHoWIWkzqY74fZ0sw006jdMttOOltfqACYcGVKkbOzwnciF7Oyf
N4QwOhRX4ee3Gm8h8UQPU+xVqvQbswQsCXvF0VXpsrK5qJLHUbzRk8BITMCy+Uit
Ey18S0T1GXErymS6WyVXroC1HI4Au6QrXUMPcR6Nm3PdoxcqqtOVf1dWSKPqpRVD
1ElMHtW2U7xd7asf1Wcgm3ODrzf6QUE32qyzVc0EvxSfTPJMdCfiOVPKz0xc6KS/
zT30bVNMczKP0u5uXMdtw8Ckh9PYwtYqgqey5s76NP1DjOGQP8C1HOidpC7IVYEg
3cGOKqLla06zW82eF2UfBLXhQXZ9kkFIPfgCPX7afcZm9bsTHzgpmWbA+wG4lBrb
jWiVQhgm4XxiKxG7jqvFWZ1jlsUcX9ELA0L/0S5FyiM8809nVUM6DmDdU6rVmxMR
58GseT3d22jObNyZX+A8jaMLpOlD5UDZSz+aaBdrYDdqmgHcw3ACLnV7w1xZk/bl
KKhTrRGAmdl7iYLtSO1umXrJLhU/9tNJgGDomyB5kCHym119up6kPUdU4RxEuGw/
YXljy0D+oo53hycbNzla/EhMWdO9MvST6+4qccplhwoyeItxr8HYwxPVAO/secNM
5HvQp0qdTNZdNY2vH64aLGQW3m6O0N/INwAd+ZySuorjQQCa9CcOdz3OksfOi9km
sqoVt64OS/Bc06Ln08QmazwIErbOxbuUYanlHyYnHiBs/O/0uJf87Oj6ccXv3R/4
rWJm/U8ZSqLc/O68dvmimZGSFtG1XuQUNWt5HmjqJaSZTn+C9iYv1yQGNgahKwlC
vWuFGmYjTtJ3yjKK9gJRw0G4kuXsSWqtVYqRhQUly6H5i+6wvHh3AWaQ5lOPYSwb
qodgI9gEt9w/cyBSFNW0cofAS6ovpAdkZh/8lJWfgKuyj9JJfKMjFeP6UK2lctqL
dyb/xxCYmkx574dHCWXqhpwDsXdM71ZCbzquYaOUqEkLsk+Ex14Li7yK8n8QYMvN
mJiWfY4LmZxvCkFXpuXEBrPv/A0OCL2DRAw8P4oitT9EXsIpg9Gwp2IgnvZcd7da
ka0wuZFjIyM2uHKG4L4Ghnq5ReBJ5MnbzvrPai4c4WlEdR9cba5poUum0Mmzbyh4
kZMlm/ztnEL4PBcQAGT6WY+X1Kzc0s27TWifsBw0fcuGDY9eXspc/971WPRSn0yW
dHmvYL3LHU2E2Mth/LFee6q+pEPXlv9MEEQqS8fpS9+yxKzRuusD4e7jzdr037k+
d2SoNSxGeKPBL5ajjFAgn+nKSxs3Az7Wy+7pSQQ4aTQQrBxGXTuAEDFq0vnAj/YJ
T6wMG3KFiJfX/WZMGoUxhrCOdeIl+af5OflDnefwbFBJtooqcnOM6a6VoyPvHVS1
UESCoVW/DBSVAbEiDJTJ8DfWyAvcXjpwy7QdOwxuwKxewVem2B9gSqrpS7i16sqm
Qsz4mJ78wMhIDxmuQpdcYglsf62Si1CxjiWTX7cNpXxXzEhUOvaqYCOVJCKA2emd
UHKaUF5KUVx4i0K35Ng0dKAzgBPxSoZcei1w3Bx8uEP0sJapq7xb2y5bTTjKB6wL
8NZ5Uxo/uTxMoMgHGmq3eGpb1Dt2SCDXUrJqVyzHz68ri7w9w3z0qUTtUWkO55F5
6njb9+ruaxBz8IUmN75s8/vPDbDk8LhOWKC0jYfovCouH+4bk9JZb6Y/tFLtlgQA
GD5Hv5SKoK0y31AfsqoD0aoohgryFfbCUI4QIImwh2EjQkh/dMpxlFR67+A71ezD
4EVrp3h04xTqn+GZSExviMs9oj2Ql6AIIaSa8Gms8JRK30eh5Hv5Fti0PFTaUm8x
N1Rt/Z48eqVbPZdFC7Z3njMViW0YAgCjpS7kbKN6onKv7PPh5wI8/uYcHScVcYJG
iFKaeziMu0Rw5TOQ43me3MgWKBNq9uhgBK+Ddg77Lk/IQynai3yvOLmnBjX8Flts
GEMvt7Lt44shzx3gAuGVvwS/YHSHY/UJV8Ov0XnzKxdoWtBHEdXqCw5QTurkurzA
tQLFKhGHlegeS6Q3wv5DKC2rszS2PbFzVLSaGqhqvfHnj79Pc2qvOJaDnS1qXL1a
Os2WWmDNqmvtxK/qcQwXQoscz9034gZeO8Uv2fmOD5GXgZP2psvFRimo63inkgsi
EWaoU67noNkgDQFfeQQiN5JKgl0wUlxGQ4fCmRh7ivWeZqYrKHWpkSV+aT8Ewo64
8reWWz+fZsm6xzjpqlKryoB77DyU0WCGfMycEVUNi03KObMffVBHeSU/ZSqsBUkO
X5Tp+W3NJ3cj/2WqqPBng5R8APuPjUd1fex+f8AzFeXR1GUOFPCPhvHCTvpgd3CC
TAXFULdkssBGLw5boT0UD0nBQmCPDLx4H70Wdb1HpxRGWUMCeFbqPgBKk0c7VfK8
QBH1+iEnlSjsUlPoOLxXmSj2KBtBUVd03TSGfEnnHKW2BtjCUdoYrJ96CXExiR5w
Cu1hRrIOK3qxxK+tKyizPSacJw1VWWdiEo/qxtr3A6SxWkH74kKjHPwZk3FETzoZ
XQe/BzgnyflpNCGgPqZRkbXDOsbJhrIwOy7ilRNFxg33pG2W4uHc4+Dc3A6BQNOU
ZxbPTGsTC5LE4rVyAUg7h6CMuQDBd1Bv5zZC6EDl4cehAwC8bYng2hv9MPSuB1dD
7J7y8Rpout6mKzH4ZMhpk5Z38FJKy35QxGxxLTFy5JnHjbIJle+s+qj5YUy5CRLM
g2zS00VXhfp7zNIKAQPjrFkzifB5qxXNN3+Pu9RWx7VEDsMSJ9T/jM+xDBTYmRHe
X9bhnXaDfGisfuwBkA4MCgp2Ox/Rym/kFnJvCL5FFyXZnv/Q5jvbHjB6JTBMj1LX
U3Hk1+Q9b0ZPTO5obAxuBkefzfKU0GlXZw5Bl1+C0oEBVZeG1WwylFgoNH6wbaZC
S7fqEhgnYOGvDQUTYb3AUphfemDk4DQRxfRk5JAdW/4m/Y70Y1OYZqk7sTzOPxcp
O9jQ3hR94f/YYjVlDuSR/TNiHMYkNFr4cw6itL3C0jJNSsnDN87j+LGip/Wz2RE9
v6deg+QCqvHiTCxK2ySA95/I+8Os40lO9k0ZhaWlybWSDH9PavWDz0wnTlFO3eYx
VzUcPHWtsLpHwBkGVCWGSJOuGaI5rqoQ8r7ZhCZYuGk9QNIusNtW+fuxbITnMZV1
YSZhCjSTFjTgdWZ9/2eUrfHc8QgMKFKyegztqVZ97+XgcniCtN02rMNc+GzDXvJg
dxZMxdDrvBezTOoH4SKjTUpX61GORi6Cyt/muEUO+R1fGrFrP9JhJLOqZr1xVZUu
NlScQkwtG6JkGgmawepfiFWKCXgxEuCcDFW3+rYDrM70D7R1GI3B3UrWQ/DqdNXd
d+v0LWPiUmtRAuRpZaL2s0xe/W1X7iDXmdqEVQqfRB6+URM4eeu6CxntT5J+dhR5
fmZXcUH0TJDpNHQop2dj/qETParNrEbOSJdtMUxkv+ON5Io1w+ESLisreGvv7838
NZ4iXcaO6oMbITCIPB6X19Pw77EMOyAjFUz6vo2ariv9k8y3HxxoeAteDKl8OoIV
uP29HMh34Sfr5VPe1F3O5mW1Maa+dAxT65MM0UTJVcbhZHCzCS/slZnc0E+uU28Z
e0MzP2c0exeWjKLoPM4cBMz9vEksBsoR+VhOyL6EFGkV+9L1YLGgbeGLFgttuozH
HX1s41qm+E2GSd46RRmC7PBwW6o3m67qCS/0rRwceqNryTcipzvt89Hy9RKEjRkX
nGsnCFQWHkLrmo2yGNvAQMU4CSHIspOpTV3lWoMkSKyP7wRwAsHxQXmdt1hrXCpY
GdMcSK2jlaBYOuKbz0h3lylGNwfSHmpzoYCtNlvTX6/KyKfV3B0sjUPl55ZkA1pI
iz22qY5y5FrZ/+ichQpa6+z54fa58hXihM6deQuIW0svFfgfNtNyL7JpmCJ/Kwey
qov4MyOzZju0V9fr+zY1jilxCBW2kq3SWtTcMlwiK9Cwdd4b2ZMM1yMAC0qspDvl
VA4s4e1bXSv1we1qTdpGgVfIzFIZXnHNkN9/9aBlWCkrIFxYmoK4Rge0v9p9zQTE
s7baHfxycuz8BwEIiAYJq4j9eTW8ZNJrTlra0YhrV4Q+U6176YRhDKJSt1UT+0z9
9ndENa2bmP4FLKifr4VuNAPV0GTQnVwQuCvgRb3sGEGrwOLwi1MSFZlv3OgPIDsf
y9y3NnsY7DAAan2raUffZ6syFyUtzGIWVUGDcmEzLlQmnhP7PlGVaP0AnDG00YDJ
SQq91MWLJBofZ9Wn5iSHycxPus9ru8v8SPVGeteMC79WYuYtjRKamFqWze4T0DQa
0EfbPRHdVZ+0pCoCPB+MnOKFACzga/M/woCVqpHe+RvN+fu1tJxpuP1L4KFFf+zR
9RPZQhoqvEt0deNraWOBoBV4FhzDMzwl+ONQ2B7QIbSkKj6cjgfk7kRNzH8/UCT0
WtoHIuiuDnd5ot/fEvyXBdPi95S3MZoYLl8jI3vEPOJ6bl4O4LAP/mCPg2FdsEP+
vmk6WABb0xV77B/1OVAjlLkhaj0zru5h3K3L5kxXuwEe+Hnx5GAGD7hqLS+NkLf0
rePOvxZ9BeiNJ8RDTvS0iTUkpsFbcBiRMhLcGlcN2D62lldZpa0UeLqSDOSRJCYi
a7S/5dxRR5kiNqFnDzH9/LBUufpz1P/36guXQcRqJQ5Id67zWrw0iiadQ5Kjrrj9
1sYq/01iWBkGX5MnMWfhgEB49YSSSe1T4x+o4yQ1zEBVKqxHX1fHDw7GCWMmjZ8J
6R/iPFHXfiTGzdGi7DgHRLpQsYsoINQ7aiZp4cZPlxn4sFzaEpwOS5knESmVz7UU
KWXgSlOChada5p1BV1LjZG8JPaABc9pzQXQP7aU+saHn8cZDdmXB4Fvt2ItvqO7T
Ik7XAprurhi2gIskGNSd/U+JV/EzXG2wXSNLq3fW29DggpUJUDhvuovOOmEyZYlb
fJC/LwGdfY73o4RsMGgg1G60zgRgNsyh/bxul4V2E8Q79Q0rZvNTaA1Q9r3be4AP
/OHhqUXNpYYm5dId5QORIcQkhsd1Z49n98Rqr+L8dHZ8IsF/xtpyrr6mswI+ZT8n
gOdhi4aXZR8WU9mAzjTJMIX2cxC7I87Y231uVHEMM611n/jPqTG+ZoE5qLWIapoQ
MxzdhLGnP51+fUrPYCq5iwvHCSQ0siHc+eQHIswAJudidXnQnUiO5eTWvXwYtU1f
5I1zmOdtp0a8y0bmlC7NA4Zt6K+vHB0YNx8KvGwgso2uIjH45li0jd6ww3xkZV6F
Ex592cLszCM6YVTH2TmplNm5bys8KPzx6k5I1A8UBLkFLWNVPJmLYpzudxWafoAI
A/ylawij6gDEkJqUEMgJn/yWXlx2TlyKDPzbNd932gRsszskG1IuPZiQ61KoQZCB
pFvFnmtDnIxUEtg9g8TLG1YYd+vem8wwLVz/hMNzT0FAtl4ExxjH9Ip48RjhiBfc
Lt8aoQ0IboknX3f2TdA/zKgrd4h3Gd9Zq/Ehj7KQCMm49JHUzDVzb9W/Kh13rw2C
pvummfoZoX7LCY08rbumxUI1TMyDE50cU0pE3vzrNIV6b9pnjbu2RU8LFjpn6JEW
ucuUOZeHz6LXy/GQYJyHDKTCWK/Kmf433mae05suxvXQ2cNZXt/pnFjgoeq1ESTG
VQ5jB8t8+Wk2hmhRfrtJSVQZgYmZsaQW7Y46d/Hk5Wma5QNBo/2Cr585TrCj/9Fs
WmmIuo2ckADAHGD1ToG2CJVwp/7m9ji6FbDs6NI7SBfSjen8qNbCZWMWDGfYeflX
D7+nFUk7pRzAKmIbokwxhDg+0e/+wPgNXa8qyXt9M7CJ+UuRmz7HeRYrXl9g48e5
E5tflrHBR4P8KQbGPhSOhimUNVye/FWhasJdp7U2SNAqTY1uavwM/DOD4POv50HP
aocJsXTU9n1u0r035dNNNojHeySNljr9IBFI+ESltTVZKJC+lBcudHR5toCv13Px
M0LhEHMciniWOYJY5RmybjAP+FlqIC2hsLcSTIRbL+lWTw2CPyazH9TDCRIuhKle
hdhR8PLitr7v/P8MitQfvlBdaDeU91hFErZBfMlmkJ2UNzBhR/b4dQherz/Xuv77
gUczdH+T70OO/mVN+KOUwFaaf2IigtfZo1NbZQp+PPZY+1ovKzFZvpnNU1PKvmZr
1WH1cmS0h0neQcYa5VWoTMR3x3bHoYFgReSkJtQD0XJIH7x5deDTFH8Y+XACqQQw
Y8zdllAZJIIzL5Qh5OHZn9REUIrcZgAcUL3DaOXYASFAxhgifm6J+MmPPrkUEALW
800R5aeLtQB866E+rNAQvGYRV380P5HxdYszOV4mcXrxVJJnyoLRoqcxgQE/EdXu
fIIoWmcjQcqboi25Mkt8pWVeKy17wrqClZ9FAKZD/9C8W41WJX1m/zDczhFyx2UM
kwzEiB//lPdyPpvTPZm7CDCsTRE8muzKXd6KmUGMO1aTk1zNMEonruhev6V3FPK5
jtwa+XSLqCNpQVEXax4bra19rkkoFZgRkY7UggUHx/GS47ZRmKZmQMG0qL1ln1fB
HFzDpsgJB3HFtrOL6+dxrqNyAzJJzTUA+icakkB5SvLyQWQeczCqX1BexFVuKmSj
wb2Pm+Bleht9MWOJeYkY5jXiAAr1mjn6spKKUUVUqo8o8GgaN2RSErlmj1j9OqeB
bFJM5PCcsYBDygKf+rxjNoi6YQoMGVcQgkE2hZLeb1g+rLHZ1MD8zl6v0jJCSbSl
fInLz+i/bA8vROCIHjbGgNAGgw2L6292rMAo1e3sNHXBfLHwRu08ZI2uzD7d6oKO
jpxgsUwKpwmvVCbW9DX9oUXn2M2d9/LCjtfxN4yC2CNuUCDMCY0pPBnHs4LIdDo7
ctCGRPbwugmCTdg9v2sUyX8DlhBEKWaHpBOTGn1PU2CIOwbrWnB9UvokTz+tVfkl
RAp54QwyAnp4IhMrLRWDfADDSMlfGxmIQGKxJ2AzqalIfZfaPUtMdBNmMRb7+CG8
qrbTxr1C2XcG7Zo+1396l0M1RFWBxiyNFBjgQa0psc8sRW6UMDd7dzDAjUZdDmNd
dGIUXs8NG+L4xzMsYhFMV3vEIRFfSOz3eYkZ8opIRvGeCJp2/TQLuQ8NCf7WpI1D
DXBKhI+j3k4vS25OeENEwaSTEfGAxYDTycXwr6inIFNyt8H+udk2NLT6YNb4BchA
C8dx0nCBbHV1HvYetZP5qW0IcRzRgek52qpRqVMvc7W53tzNZPd/nICJcwq7YOfc
dHOUzjqgooEY1ZzuDYw/OjXUyRco3i1roAB0wylHLh3ErPWgSiPtbAnFlODgTEL8
uMBpypvGr5UL7Kj5y7AfMsDG8gAopdtqqcIJt4MRjc7TIInFS5RCes3CCVDNYcfU
HGU4WBNvDE/a9+Y91Xzw9ZKnXxNoKAp0QVgP/fn/glxEGfm8r3E2f0PhD24HXDYm
sRSNd1t47QCazZpROCgoZeWgBWYl9n8MQK+qm3Fm0egrI7QdVONA9e8mQK5B8V9w
sHyK/O73kl/V6w8OcIHNyaJ8sblTsjj7o4e5Yp/wGG6n8o1VKK7yapJvA1NQXYNJ
DJLYvhv3y1G+xDEEYNk1xOlL/EHTJMzpBxYCHEJFh8+YJX4o6fy8UEiGvNVzXkBT
yYr12fobu9zLLurIBeqH7l7BCvh6+3+43da1wy1SayMa9DGEJ8IEl+vRwYh4+Ml0
m/oz8z5zmJO2dhws1/id0tjg4gz0EckHW2+wcPC38K05VS7fPt+TpvwrMnAYTeQo
4NonujS1JD5jjAM/PthndPqAOrJweHc6cJMcLZBNkKbx7dAtEHgSVMAcJPanLR4l
kuY2UQUMUq7e003e9kVmAXOEp3KNICpotNUwH+UY2vP7wGKg1+1bVUfk19PjWyY/
+5iKiC+yYdsHmPTU0fx98ozt/pdfaf4xxyeHLK1dfeMGSNRKd/P05Pue0I+yJ3sI
1HfuQH4G/sLc6du51dUyuIdjxrdh1wJ4BfVACk6xWBJMxliJaxS5ftR/CIhDnIzq
ks45mICQBPqbttVdKY7sN86aKk6LBOMrHI45XEKVaIipKms6yGGeLf1UwsYVIfI0
phQavTDElOlXOM/UXvfWnZCeGrHcHOGMD4zElIdx4WuOIfChUMGCKurnDnGNufHA
jSC9qZaFJytqvFSepBRI5wxLC+ec/pNL8JHpONyRPqwmP+kNEZ7ETvGl4DSP3UsE
efw286Q7q4rE7v+qHpmTSPOMtJDKPnKn+hpIyAxm1ViWeHcHsl3ZftEekU7EoY7v
whXZ42Dy+GSvBxgmJG+YqJB3dFHMmA7iIma1MV3dJja5c/jxoJm9TGsDknwrow74
tNDF5NcTmGy7O/Ui0qdtw79Ah5qjCNWQO14HuoE05V7sWovOU1pMPmrFxsKBsbCn
kWndhelS8Tj0wNDPSz2k7Vj8248vGR92AV2FY7UV5z1nJ/AfG6yHpIOTHU12lAtd
j183htae3cHCO0KyPu48lzURvj3QqaHJfMUdBspCCf0mrgINe+X71gr5ZfCxpSCN
pqZU7hzhHNQ19pOOaV20Bk9jYyNnUXIEfjwnwoAPw75gVfsuQm1pJCjqEYbiR6gY
iKsjFCKP7qfr3h/8Wn0zCHu3xAyJXMu6Y3pjduB3A05K99IF6rT7oguhuc3h9Yvc
BMQsq+IucFOXB8vl+2TYUF2HD6w8GAUY28k4o0wqp7jCSWuXZnemiBs+phDiCI9c
dDSXFibF0r5BQSDoZ65t2ksfjsCmlMMIarG9yzBdWom1bowupQ5RuHcv68OF818U
oXytcr5cD+9cdva11vsM3bdx6Tdg/4oBxK7Ew3DS32ejR0pBYrZF+7aVTQUeTStH
dL8DMAD7buiw8NTLSDOZFcdtzgAprt92wUK8rqEZ+oDUdpfrAR7aUZT3uVwmVGse
bZNLQIk3Qsd7j9K6Aa8ho+3NDYDTnAvFn3TYOQvJfWl0gYG8/YKrhXS8YZz5Yxwj
C+PKlp/lR2TAI/B0eyxeR9U8msHZzIZMH6xy3a6k60K1Y7vrOGkL0Y91yWxhNwbh
aid73kdd07lWuq2P2mrnER3Y1qLz4I2HHKLqSMjxQF+rueJB1t3PBPKFF6yVrxKi
9okSGvgY85snjIOPktQnqfFex69KyZ/B6s8a/tGOmzkYn3xxxd475pQ0h7rYazFZ
6XcPKPDf1O1kKpKR6du+gVZxi2HpXKJ2HljaX9QvtN8Tn6MuCu/jdI+GT41Y6ZtT
HSIcqSH99i7m6OdWe4y8KsfFx+vKiEuRx5FMIJEPn3Ja5cBahQVCOX+hseuxrRm3
/Q6qj4Kos6Sz1imurUr5Ota/JtwchNT35kv0lM1UQ7Y4r4MzvMLu4tfnWyUNrAYO
ClG85raiSuesuvX23ABS5qsNN1pAV3pTYrpKknXp+9AdYajs7xMylZlCaTEy5mXL
WlUghSidKd/grFoeu2rqXYztVCfqrH/6cITMs8HqVOEXJll/wELx5NPlU5cD0XlQ
NJxqC1ZW6hP762ulpE4KheKc13RKcMzGm93IUTAgXl1X7wDJQltAWiYH2dXwNuhB
FqZ4TthzR47SikGQHvnwwb1zblb/h+03OhEjfgN3UgWMLyHutwOCT5vm9GwxJoU4
w9eRtMEnSvXYOs9hb4NmG71o842aCsmWj//ZEU9tH/FH67VRnFwuTcONQaV9H6W7
kncsJQ3o13MQsunSDZ1C+xFBhs58VJHJzKAB49A20pUW15G12/Zzhube6e7cLKzn
gCp+SFgEENmhxLfNDLCegK1cA8hIuPuiGwHEDZWqC1fWg5i8uWsD3Cj6EQQWFq18
K6spRd4Gf0lfzLEFR8TCjIdLqEEwtXNb8WhXe8C1IPTKtN1JNGB+d0jkKgoxL03n
q20bAa4U82phioS0vaeqMd7gG/DhUdRyHLvf07ES29o6v5hbUaraGEDPAVuTb8pp
woA7Wzn7nwbhI27gKgOi39l5tYEUjMkaUtsg1JbcGxCPBADLwf87j6BNi9kth7mb
EkW7w2yecGfiOTft1Q5cFBo3C26YrNrg6yD/wVoP6cB20U+DxH7hVKb5OSJt9K/p
1D6Pd4RrehBiDf3PxgKCHCSlsdYyYIcTYd9JKAlITpVYJVH6nQjAMRPb03uDflfv
ECbYGtkspxl0Bh8ZNATLkIhKPHzJUnGQrCxFsRCI30TIAnFa4Zh4ASRCHPERJ5nM
VzxOSuGMB2NXYnj3Szbyw008AIglZfvf1F2HbRShwTKZHIi1vOJyOG//EUvHrqkx
NbgK0IpEYXJLD3gKyfhoC+1n2jLsA/DZqHkJ7QhRdxMZ8BW6xf689FC9yBX40+i2
7IpeaHt60qgDgyR2gSk2lU7JLmyMmPLXJ1NtgGBb2TZ2cFWH/Icp9xgjou8Qm/7W
nKKS7yVlB/N/63WY8hTVmtJNXCQWd2TTQYeOVgCltv/9bSaPVf30kBmR3CmVFYtY
4q+SThOjWW+BVp2JFyGOAEo3SPBsid7FA42An39/NPsMWZr6IlgHmpPrhTHE3nG4
nxl16qFRuup3KnD4hd/g4plzkBy0qpZKYofuaY76PI2FNcXhKFkujumKt1UGOWFg
Fa8Z47u5L+7VOcUcyLS31QU+4sl/Dvq5DvN1h0AK17ddG7lDVyJ7skUTLtTPPyl9
kH4gGT8Xu/Ly2kxWI5W9zrz0om7J2Ueo+EgChalw5xvewdC+44A4PGLR/dywLGeH
mq9rl5st93I5ywcOLYC/GQkBz2/ykVHjCC27hPBozM7HJeE7ctxwKWZumbb1RK5F
wUo7dxQLsJ36Bj4/D/zF4q3GJqgLkJsTrpX3KG6BV4Hc7nyY4Lx8jUtCDeSo02am
j8CYtbMhSOabns45VUDDE00NcYYuv4EiMWFmLNXtgrG5CAM6QL+u5WYJB5qwJ1WL
H9MwIJwnyC9R/xamuoJYrFkdySgpdCORW3ky6g0ZaDW0xdotIeD1b8a3b3HihHUC
C7W8nUcul1gUjPSnK0ZEaDfbUnEx1yjLOYLSjkWhA1kGqirSTOfZ1hyHRhoOTxbn
x7oB7hZpzSFYbf6AGXxjOfj+QfWyFfOxRgep35SRGZvoPY7nz5pc8Ou+D/lAAknL
O7RXEMsV8u2CrnSVBipAsL458vrb5kutE0QV41h29Pz2bZ0gFE1G+j6o5hV76bI4
YjJXw+f1S/OPhd4yiil+4ZiSW21GM1QgjkBlXIu/EfFVbZDaTCYgmV7QabTohOeJ
mBr4LHU6XNxtGMwS8iD0uEFuXKnW0s/OeKFPOXI69gfwjCMhkDrGTh36s9OMnQMW
ar/7TdCWY8trPHREFHoVWsuKsnEjVkAOczEP7s/VBwdcpab0suBPAeNPwZ6lSMzc
06kgOKyCAv2wXRgyW7Xl3+kIPqEqHz0yqIDxLA23UQfgvX9ZDL8POZJ0ruIN6jJR
F7WGni65XMHIRdzCNZv5AJG5hyf5qcHJ75/XIiTapdIhYtCJkpmIVmepw2T3xG+D
b2PEeWpaiMIXPqc0KbfSj02agxWhWzHXmyigogjsXDtGM7Eas10d8ulNgLngg8At
3kePQRM0uwLlRU5PidFqV5qGqZMXkGFa/ZTm5+H4VhO90SubfXyqwa//m3hM480b
nlugad9E6owGpGEbe8nhJim4sF1i4C8DNgdBUamgESG+s2sZkPVD88NYa/lvIg+F
mWYtPXiMMaEQVJQMydXGCSeJlIdVeNw2MCkMVlaFQRv/xYDuLBKseWgbgpWn6EnF
pO8TVTdevLdO5BL9yZj1t49HVZQpGh7+HtvEKmGQez/1mIRubD8t2bB3lM/WW3jX
nW2o6QR1aviRVFL2O2qQI4uJ5IQ5ka0p3/pOB9PU0YX+D50IWsO9VYtqMiL4Qyws
rqpksjGs6PUYdw3Q157DvmtMUGnNU3ThoRBUW8icIGf5uonDarAsqpAiNoYYSddW
wFxDn0G8Z8r++tSk7YfcU12RYmhY1Mrn3mjcEuFOVv611lj0SO8uFKmOJw6PNWqc
FirmSN12M3RUzP4M5eObEzD9AKOvL9UcVQKcpSiI/cdgnvai6lzz4/FBjFBaIHej
3qGQodO8CDAi+hfib+af0+zTCyBhfT8vQYN5TQIFBlIdvvUadJ5KCi8y0eO1aIai
j934XFM6U7CpPysadORRVJDfSi6Dsv0PULJxIDWpNIWucEnEzQVZocovPv4EVs9b
1L2HyXeRDBPL3LqCIXmoch5ZnhWxa43OmMUqrlOowpE1SWWlsGiOUGM95MjRDcgn
RzGv43jsVkPSlSXZ7tT/LKvn+e3WgDJ4aFQQbvtKdOtMuTJ+xPO9DGD5Bv7j9SkN
fWbJGrqOHxk1XGM/bo/tZZiT3AfwTUxpYLCx6EVGZvUivfL3C9rScJxG+Fp0VtCA
dct5agTkgNi6M4+ba1vbNPWgpjmbJ4tBr0J5bWd+V+mMUoTY9AEj6+J4L21RSfNC
ShQZFOXa1FC6qOpshhAZZ6a9LbMmgx1O224+UP22s+h0hjRqX4b7h9QftkvrSDaa
1j0YP6hU+k8EVbGMu93YnwCj/ifSuakiIPz94EgeVUotRiWVvURr0Yw7yX6Qtb3y
aXNVtAkkvA/pVknicRxB5v1f8PBEIxQcheD0UwpcshyAYMLiCk94VR82inNjYTHJ
n3R6ItjHfZtt1hjDC06Ivm4yyn0zfTuuaHy1NadojNIHyv1LLbMXjrxcqN5yy8bh
fuKls+MeOzO1KHfFsAGH0JA27+5lpqUctzGHD9/dyf/qWPCxyv8U1//wNOxveY0N
389fAXLGlHJHAQeohyf868+ZDLmzaDfSRDM6gHJtrZcZ4J0aqJ69k93/isPPJXf6
ylcLBr2+OknOntMuKTTI45t48P3PTmDWKGIJ0UUantZhRaznOy6JtfoAiEHhro3X
DRuQVQO9wTTD9eq3J1sDGTrysS7J2w59oZsBzN9J4cAWNmuO7Ri2g808GH3aWVU6
ie54uZ6JCbH+ua7g0Lb69qPPVBN/raXxKjy1puIqVl2kKmOiGn+xM1WxXrfi8Sfq
Gvon4azvovpI2hUCTruk6UNDWAhKZuSqwWNvRNRzXBMQPun3LsfcxwbUyd+wAz2M
YegtLVWy+sIAoIFxUVo7yt/GLKA/JTsAM2wdyLAEhzEAsdb2xF/vNsu1mLonZtJW
WyIpy/tVkMmSIUQKrZMfBLulyVLJpvsvC3KyMzJIxltjuM0+nNZwry/RkMq9GVQt
6y14TeG2wo+96U6N0rGTb3mvAxXz94AFsFATyPaQqFHZjxJx65TUbvbe4hDYosoh
GYzQPmX3P4Jf/3VU7VSHlpT9HDs1LBnlPUBuu+pCCEsKCbeT/7Vt/cj6CbBaiA0p
BTw59hrURUxbBzBVQQ256Gv6JN/2/1TwKwVSXkpTXo56rENGzDoW1qkVAS2I3RLs
6w/hZjEYh9n0W30frYMhdoCRQdvRzCtk//84wjcjKNdnulrBKaa94A8HTn9ARzOF
LyEQtUXULyaPegzf0XrFoNPxspGaUvFZzVD4IQphonvNSJDVXHzseYvUISWuKnO1
qeK202pIvScb3vXtC6zk2+6Zl9DKxYJD1MpADYQZvJod9MVXOUkhBD3EPkfo3FAs
jjrihX20eomwIp4Dzl/h46mzUGaeMKF9Jz/w/DxMWR68KJ4WRE+njWAXbcgDnEtf
uQkU0bHuTjtWyQrTwsq6tNcr8Ljs04RXVjkltNrwucKAFtO8qf4t5MW8VY76QgJt
FiXyWA2C8kjgabTh3o9dipvw+ImBchKOipIP4i5D3YkIxpi+GVxnXnvktOrbXtLz
PoKffWJVjlSLVKNQls79olNCDIvTfon07QJ94Ggx++QL1sI20wJ+xpIM/xE7dTYg
+DCQ4CZTezYEha+D2MxhzPnF92ZcYE7xgoJqpEHK8lz24zzumhHglYFoMGA055UB
2O9iiw7gwyOtJfpwOMDt/JtaxtY8YjyvfbXzOxFb9MItA/NNbFYa7KudzoTkQfDn
O/U/jo+sROu58Cv0C/sNPKdesW0P5L4fbEcbKv9nRdFbiqzAxE20P0g8aJubz6M3
UTXeGDncdGf95azFWC4zEbxO9Q/djznHJKyeAYvS0PfHgjwgzv+NIGIqkSdltqPX
kSdEhRO+BILhfXzn0qMBOZce41RhpEjokw4ACr18fL38UrQZkEJ6Ez4S0/Vja6sg
ZmevGLDHJNo0tMd6FIMGSdqO24VNM5YTBWORS5h5f4FROzE1LyOxZO6AN121uO/K
e8JbteiZe01k5vSGbFI5LGqZMVuscPRGYVFqxa1Vilv2IcMuH1K77xvDYcaxki2o
Hm+3a9Y+Ab1ArwKfor1Q18OQ98CdM9RC+zLwfmo7KSKrPErPYdBCygM7aNkEPsMs
8tOUjDqoe/RBYsNeKpcYeqDTknAd7ohbMqBGWMe6UjXzy38OM01hEg3PLjFCTMrI
kqPsRVvMEHwuhR6x9mB6Lr8FE7hpDVjlJoFLYnlKoUMEI1VJyXCUkbUqJHBLte7o
7CJCctpDrfSoQVjmthZqmpXxxi+ossA1es2/qcz7z/gaX41QR1lncs4ZAFygA9T/
LzJhLYBg2CQk33eKNqu/W+QIy6ny8DZ7NmCa9Bq36FOugL851egr35DDCe9DUhlN
Ggiu7QSpa8ObXcFs1gcrxLNouUm5wCuMUYwqSOj30tejIY+Pw6UVX/Sg1hmz1t8D
EVB1IGPVEZ9evXvoo/9Rjhbu4qNE6wXBHX6jJDPSZwkrVSSJCmN7wHZ4SrIGSsGz
9OQTFrjCsWtPBlWit13FUfGFGYKLOZ5geVuapFYsSrXYXhE/uA90Z9ZzeJGcHtgy
lRV1GKNwrpllRCvY7nkG0ibVA/IbA9/OVK/Vzj5IRGCo1hjPAVp2j3M99jrETRHK
lXM0AX5/UhRyJFIVgWjXhy6yYUfGlwbE/bJTmIAo8VqFcsNLDUtUFT4udch9OD2v
c6na48swj8skyHKD/3fzV0DdIpn6+u10M6Bo/t9gT7TRKFyGg/RHq4OdWPbTri0C
POeeAyQTvifiYvr+SkRAraMSfpjrFdC7LakDFsWgpKY5xPxcSQq5T5+xHtxn4Aqt
XQQxUqvicXYSABONH5KbF9ksQHPcj3Mp7Rk3HKW4Zri3xwiHWkYRbwSGiuF4iTob
FM7Xiem3eHKfVpSYVl3uya7cdLgOkTAibdwmgiRddQw+osav4y1Qlc3URSp9zJ9T
ZM9OOz4CN67E9BWlX49Wex6E4iPI8YNRWckZkgWyjVJCNP5hTGPS+3alENNLW3Qx
AFrLikZtoWfRwUlq6Cz7WJgz+mL/U4qTczBMND96cpUHIUs9BpFVF2N7kkmMbWXl
UJ/ueBnNkXoEHdKJ1NQYj4hO4pN3DvyLJhpQAobjUew+IdryAOncZHrrbyP0gIBm
0u0Nt7qk4LREPCL2LGqmFncpQGBPPPWvz4Zr6+icLZsippnxqRLWaa0qLUACF9sY
aC2ewgnXqWYXDoVuFJL8ghaKD/ijP6YiPp0jWYKfVax6NQgl9szNJnGuHeMfa8vo
8FzJVBMk++Ye+EEXOG0ywoeZKg8bGC++pfo4A+opfB8C+mxa9KhcwsloV2WfvcFP
7t6lh8YgQjgK2aPjcyTW0o5+iEjEkyGDUzHqRtamEsugB/tdA8TzWWJ2+6cmz304
Hh/19z5q3j3J3ryrfB/jnk62LUjAbnxEtZMAy/cGAJkUcjagOW6t6qTH9ubnYHxD
T5FA1aQJZelCfNfJNpG7L3vE4fXxz8NUzf49StjAbFRUbmGrsVdisJvBNFteS7L/
7DcphEp5U89c1PPxEhj+3VosFCF9fbdRPv4bCSqhwHvkxiKLtNrgxSID3vXTK25D
u7yiN57pT4eh3a5YkLSHqQa7XcsJrB67GS+oqLdDjuHy7y5IrwtRgOadfixMeuML
gmcWi2F84Afaifx549lu0DoOc22iwXUd/yZ3UKE9NPI9CTp3dtAzF2KCkfEuGz/T
be6jcg5mJgO3IuRveEvjBTtaO2yXej+GjW/+RP+jkYw0ma33iLH/BGbJjW0Ky3Hx
jJMo8WaxFWXgtHPFf0YrWVvQrTfbkAmyPuNTFUE+AE5pJp5y3mFzjw1zVBd4CY6A
4JOWkvCqIwlMAUpEjozWfJHGxMju+wTulLGh6fRAQF1Ykclqq+m896JW1TXYVaOe
MSvDlFlDjQeequnSU3knNvywGkX/q+IL6Rq6h//h4dalDAEHRTHkpuNy/GA6+pmA
jtq7r2iIQLLSjZgCHZStjaa89KYcZjFX7Bx/4hV315NpXOMB7PKhnsI/J283eQae
15ko6ry1asqUczB2rcm6Zo5fo8EYkqAI2h0ZWPIWZo3MmA3UgzU+Xuj3OBxin6Ne
j6Iw4biEYnU2VfBZcFakOwh/FpsoS8HF7QAdKAwFHPm6GvdtmWR5hvcHt54Kaucz
JXq1n9GAN9bA4c5Su/a+A79VzxNd0NpsQeiiTJb6btLA4iXtnilzXHdm76tNITAa
n40f7PKj2i/Z+sE3kcyKCCLBE8Z8841JOm4wrL00JsXrQFibMnHrzG3I8U7+5zaV
ycP8a8luMGHJXhenx7+VOLyuf+3nJw5GC4dgw4yGxc/JTo02QrJyqGoY6Ff/66lp
amFb6lUG7nqDqXRxH82juNy3JNq5ufQxy4InnAkeweI1BtqbQlYpT/WQCCCe237F
gZ8xpFTqN7AOYrGqD3UDRfCQpIscB96RTIHzJmfqrhMW5mKAhCcdBaZJff+IrNox
M5dcIbCwhY8hgOjqxZPEN0Pnmb1814opaHOuHAdeGYFOybm1EbUBc8MY3fXlKk8p
UMjRI1+93GMrb02zZbSB9j9lYPoGoqXelrpX+0vVIJ4pY5mmyZ/xGLteGSMrc6YP
PGiPNoo0yNYzS/+fXYAa+BGSU4K6auyyKC+RL2IKOJgA4kOjtdXdrvrVwqLKDarO
QGnpP0/ChIhiLtdqVsWrF80emXlGBd90dXvmODntsqJFPGI7nxGBfjlLG4iPnsj7
4S7bhWhDsmNMy+INXxf7qtxktWuoM/SPuSDqCZkRZHekbndFVLaX3ubXqn9FoLHM
kcrI0BHFvjA+8DPV9jQ4NXFsznC1DQSAXRws8PlXJnJoI9ZFYyS4kouhfNzyips/
ppCyiwKxDWv01S6Vn+1NYzPzSpXtjYvRkUGvlFun8GTdzYDZ+2iDr25prAuE6SBl
gT6qu3zR15FjAxfkQrIpS5vuSW7HdtIeg4YLVTjp5TS8dQ6k7So0kScA0YoxLSOI
9qUe27EjucHT2pZiK9ksJkoqLmfx24r/mdq5z5jnq+BwkFmgwB396RTyx1TKdW1A
9eoNJmtKThC0ORn0GPZPptyH0sfgNBYBXxJNAPSFAhmM4TUNsmXslHop4L8hd2h6
ViOo65MibTK6OH+MwxJlKDYFLrhA0hhhOQvxAJgNOSETgpWohOU2/12Xabm51JGa
O7l2uCVoyMXBdZ8J4wr2I9cYJ2miJ5rRuGfe9wmLhMPB43Cgkqk9/TPbpRUPgeJE
PqjllG30FnfT6wM3NDXygjxwYjV9pXpgRMSn8QUc1rPu+7PI34z/9+NCmlFG1AaQ
7NQm2Y4gBj7R6nIkgHG1+1qi5Bu9Mc/fD4o5KYC+xjQwjjoTbAcqJLWvuSDeNSyh
MrGa99XBzs+e9EUFtjR4b66rHRQUZMGsPUcOuu7dxGnlOUgLawaut5KR1R73hrQl
HmcUkKq1xgu8RKhO4LMTZxWl3/AmO3ox1ZTskkmYyyk/0IsIM5lXD/yZ6eLcCtfA
76O5OnS32nBnfuqHg4ymM7DGVoVna4HvI+uHQ+X74TGAht9g1UM2qjT2oD/Q2fmL
6ZCVAjmBKKbpQE/DbRaa5jEm99hmlIs3k7o0Al5ych+npx+TgWfNNhALsHLxJdv5
pdKd0S1c1PMfhXPhe1MBmwrICsUZX1Cb68dxEpCO0Dl8ng2nOv9RSJlnG5xENNHZ
QLMYNVjvxYCmjYxxMUs6vYCuxy3LH7HXB8lKkx3JhvUpCFRPYmQPDC/ZT/ZIqevE
DMpWTZnJXVpbiLAiI4UuvEkHDY6FW+JC04i0qNrBXjNUWQQh53yBBfZcFnVNq4Th
ocLfoeoCnuD8fsOtw1ulwh1Cy84F9zezutkOv05AEbnfQ38+x2fo/edsRSexgDTS
DfVugLSAdFsxGHgr/3V62Kq01ctGoV5MCoNP5Iwzg9rdvKNSbZJjheFaln6Og5HF
a4acvbNzc2j8zLTVIVzx/WTP0b571eC1zHiO8nNdFyFAlKrAS/2sCgGkMf8aUdT5
kGzCLHDihqIS6SoAcIoI7CHQ+stw2+/0R9P0V96z1HB3xbbbgHRjRqZRRC4zybhn
LSUdC8eBWsyWv4A07/cu1UePxL16oNnqMS8rL5Fa9uDtZ6B+0Nyer+xi3tsIT/CS
PN/dieF0PFBHj/tdJerz+PZLx9z2jbwzUmsa1DVHT/Qc1kDuO4AAXKCBIG1HtWd7
msTxRGj1WGarlk7ngZsmKEufDRgnz6LsC40avfWbgrA2OJOYQ93l7T2x+LzmdaSb
M2vxQ4MMDWafBWakyXiWd9CpCgFCMDjihs069K9fNeSt4+pR5Sz2k7NlOWmICdEc
fsWhvHBSSTopv6mCt/6DXpkuHvpkBuuqJXd+05p+tCKiFEsA+9PRFNdpiLb/r2DG
Z66bzlT0BRHW5SyVjh3qJN5sgU5avz3fi5BHhIGzicSs52GgcU6y/8f7Y3wlbfGZ
MEksahGodMlYoMJLsy4LPMZtU2Ui9E9XIXxVtNhL49mNvfq7SrcQw7JtNuvB2qk/
4W0FwrJafH/2xGwvYyW7gucN9urBd3Z/hSKakJlaq7XcjQ8CWTvIbCfgHo3MZL41
2ypjzY3rGNs/uzJV0wsWef07S+XQx01eU16Q2kYTV0Gdof0wzFG093fIU6OcDkFr
Bv+oRb1lidO3UH4k0ZdwlxDH4v1P5WaQgBslGq+BLBC8eoZk3wvip6W9UB+GNWrT
UiZ28qlm86Vz9orTKttsdIvmPYmt8Iv5TocLOClwjE2Hm8eRZNoQmKPP9JdLkDQ3
zwdzPnlGAXCsSx2ZuVTA1Maz/A/AZHB35VBLloXxUPcT8KmBmUcQmhZidhcG/CAA
dBhVez19hVJJs25gKXNo2yFXNE6wmeW9KtDgBNmZ8++oK0P/wdhYARdkPYUn/4Bh
2p7mYbsx4BvRLIrGCsv2nnPZTAOvIH+Bg7q1kpJJDi/1n1WiOElwk4Y7GkkSsK4w
VTz7cRNThwwOpBty2KLhOMO9TRoPS/0G5B47it0SwgjVhXvT1OIb2f6rGhx3tWQa
AgnplW4tyLVGkS62dyKPMTw2yL9FNp4/SidveByqNaF51HRDR9QF7jnXR57Tu4tK
ZdvAbqwnYOwIryNyipm3/1VOj3thAAqcVl5kNrFlnxX7q7JqPn2VYJ6rIqv1u5Fe
TxBtNd55u8qymSIA6eB2WVeTUxVTVYOaWMr2GOCy5OFeXxssOYE/S7bTtOstxEJJ
vZOK0WzSU+7oFEClFCqHU+eKHCyGNLiebyFcDvQi4StfsW6XaQl3eAt2F5/fC0eu
Lj/UWyyCluY2qolBHogy2B7BgOYCiU/FhhUGcfBsYBSrf/wNRa8qgGutT88srCoR
mdLqp9yFLT89miUJ4ERRRjjU1iraQ+rpj4WwnXM73tfPvm8PJeoVWCfJAxiRv5uI
tv90vLsn8/PU6fxK6GkV57AdJP2Dif/FhJ2a6vJMfgotWltajYIh03/atKAVxUQO
ch3UOQ2DE9ct5jSzgwrb1tNncDRPPd6wB2qvMh3u5r7D6T5Egn+egQADN3gJLTHO
qakdtd6tYVIP3XD2ThVQ4jwL6LnlRw06vs5GZv60NbuzKnmewo77JXkwxe91Gu/v
O+nYdXdutzEANIaiHFWDVOQK7Ba314CwMIrcFqJpfmZT7GPzDiftEKyHvegR3RVQ
AEfw9WrvAEmKD9hva+vRiDMqV4HIkdevXGLgqIBaxSBiXv+OBRUCWwFgDs3lTSSr
oHZhut6uQrQeMEFbWdfhC2s4yj+arXH812Kb6yAHBkWbYgxfDV7AZFz4YNXDV7u+
jxs684cR5T8Vq97PD7kPmrJZ8Bsuc3ulXzho6PTU4+v5NKmWkONVYl7aN5X57HWQ
7ktFYjzP7C2e4HrtnjvxMdrsEH1fjN7xmhUQDJnlyr354rCeMtpjFsWRPVB/LItb
ETFScClGTVLCEdwnKpkoI8D8rzUU55WTqaicPWxH0H4FKZ8vm+b/37xCkMfZq3DA
I3j0SC6mVq6Ogzk74C1nqMsI03By9sCTGB9b0mB3wV322LBG0aTEHopPHUJXUffF
6dW4/tPt6QaSp0TxtPoEX301cG6WEmiMp5nVeJdo7hAY2uxqpruU5GJZFqNRh3BV
gwFvdEZT8XUKyl91LitRQoQ8gNy6a+lHg+DX1IIN9/FLTVF1RVnx3gDdKekqZpLW
HDK5MMOYhjkuYPeyEbuvj39V1tWIFhNw8iEAx11hYJE/cvxQ0UMtYzAQKKa75LmS
u/UrTAF1guur341AhudBPRtkS6MBAT7NMvmL9ZOYykqL6Ph71lhMmZ49o6Gjw9yV
tYj2aAGN7FJNiylSMYXXBF0PusyjEgczz3ABU3hSPo9PZ80ez0hlzYyw1EEaDxLj
59kUObRl17TWINxRfXLAd48JWTYGBSKzt7GHSkyKHtvIj8rs8/KrgIXprD4C5GUU
o2zUCdmY6KQcQ6+G4P/Apme6FupSvhWFTOhkeTdcJclDyBCvu389+wOhjlhJll9Z
RRB+VtQ+wzKjVW338cUOt6bNh8aoqmcchW7ys7VnAxH1Ph0BzCBjoaEW2g5LIYwi
Y0mqlX0z+27jeYbxGUDCJqQjH7pfeVsg6QY24D402rbyqvlK0/fFN1lwX15Vv4iu
Ib4SqTijpxmF47TvPD72GvzQi20rGLkn03cSFB48ftfUTU4ZwddXHUnbseH7hn7J
Sh4HjcgJtrnleTy2o506iTrLARTVHRccRufjHYQ0ZkUN1EiXDQ1er4q+DiJw5ixf
ckmyUJp3uz+SCjLLJas9zOtiPUtZAcu4sMV+2vY5yMqLdILPO3I2KTntyiliHW5Z
C+LquFJeTaCOq3FB2+mH28VNqQzlEUuMr/5CLdRVs0etoxYC0A8tH9zngrdc/rrC
3GNFIdmrc114J5orI0kY0us4QSzcvvTlyufQk+97H3AzkDExaSmicBg4ZGn8KBG7
qIAX/+MfWxY3xci5g2sYYvTxS8S17DXLWMqCZyqyXM1rko3wInY+Q7dWLDjqqo/w
RjvnCECURV5k4dUDtF3r30axy2vEABcf3mB22cqFRa3FFG7RDzPQ2Ab+1K7rytws
xzplBi7Q0ox6hbh/MLX09lPEV9OunmB44/rsXvY1XYUnbyiXX6c8YsOyK2dTas3A
EMbqbFoA3r7TQ8pCnkp+Uvha8HA2CCL3SSlot9TanG1spghe5B/NAx7xSaRSv9KU
HVnP47TXSPkkzjS5W9rX8rT514Av+GTVIYgE+STv/zxmjMl6bL4C1fvv3hYs9t/J
IlbFlDiFg+0jPQmoMzOK4CmfmXUlBXLg9gqaGH1elyXQq63IKgKF2mTJ5RS810uY
qNAIEBltFQpWsV4mfDE/wi3IoewvSySGJprT0r2S/xkpzQyd0Re+F2OMVadZ1vGS
OCPLc04LlzEWIHZRSlnvK/6ErxVn/L4xGS3zF4lXyeySa/OV/KVgF+TLsc+DiQ9K
yzSuQatuG4NwA8v7uBXWUY0G2QROYc/FALnjy2k2CEzu9vOzj1hA2w2nmZZs7lAO
UL/e2rsZRMyWTSoQt8rklI2ACxgnzQJnmsUwQxwZBfJ7IKgGK8BWlcS9XAsxwaz4
IaORQj+M81yzznY6do2yKtMl9BPJaPCt1ZPqxl213XIuLlMc2iJQAeIiFJqNnpSB
K7WeOl6gUZ0KeTEV/T+hDOcLXPSygu6u26cFWNWqEgH3Wf6d4uT3UWh64/JS1YWo
nQjbCwcEKWN/A5spwX+MucToK4tmndElX8hgIAFnHepAU61W4sbb4QymwLDTLg6h
R0d2ow4Z1qL4T3vugZK/ba4KfdcyAOv/Nst+22Z560blEJTK+CDXQb68xMwOm41Q
ldePOwt5u940R+d6QiJkgh2xuD/I0NSSENxcDr/Cew4YsAbwq7LsPBJkhurueNLS
nT2J1bci0fSouyuLJwtOSaUmWL70flgJDB8ROPtJl4sIyG0XzF/J7XaIKUr8COTS
ixNrNS+fB6OlGwZfzmVSGwt7i3tTimMsNohLxahc8LSfghL30fgK0L0YHBrTkwvw
hyuOG5coVg5ZvEahtMNIslmCrb2casKE9XTChyzjcxXds6EnzUB5/7OKGX3MdrcS
lVShJs7ctHTF5AfeC0B4OTy1E08+Ae/Qh0rIwG+g6HjEiXQFbedYbwzm60KGlg+7
QCSRrOi1JMHROPRSYzMHPZ46pK1YSjdEpz1N5NBfDcSt/Rf5b6y22uzKS14CCUed
835uOEaYOeTbum4fEXx/qpbIXScj+1+UIr/c64hM7rekOHxwGNYsMh5YsFsq/WQ5
3gQU+ZY+oVTaCY5Za6d9MiajZyK7pLdCwv7KvlkoBzzUcVzTYWoGnPZfXM2YzKLf
JUizUxE5mAOxZHs+y2PVy75crVWt9HtgCistcO17RhVxQAVoYXqPhyL8LnuuI4k5
gntz5AnLcEzDVuNqaOXABoGdpUZDVUveil0ctn2c9ijslGwX4tE/B3dqFCdF8JSi
NTX1vb7rujdzr6j2x3/WIxFnCd9Ld9GammfAwLCjohqClrq90urkzaHcFbBUzSFc
cOJVRrRhatTvdgxo6Wczb3O0nNsUCnu/e/DmGV5qnqaUSfNmiC4ofm6zhUd2Ztpu
sHmX/rTyTMx7amRtRWZabnkV97e8O6pbm85tWHBZ7sDEmbFEmnAuJVxsuCYL7YoJ
9SFEff7cld2yMW7MowRjbzHqCqr/lwfgGpaOTl/IlWnyH8sb8lJFVpVd6zh5EDew
UNK2FT8u2DhQOTJXUmVwg++95lDdKLur1DDyhTD2HmL/4IHL5gkbKjJhqNKkBtTS
n+7EFY6b/7oZucsAbC73bnbeRgQ9NEjkdGc/A/CX+PI94ruL5qVVUoS5iO18jan1
yYsDdLhrOxAQNWzxNEWkeGaIzsZKcWTM7EsmzTmIPsQHTGnstR2oa479QS8y/qA8
i9vREkeMmZCSSs/2AmRVA0HmYfxdSKqlVC48k2k7JQSB0UgMkAr10jQIqanmLaUn
jifSp4sHTjKhpLwi97mMUvuiAqTicwUALxio9dCgeU01SdYUbAdk35RCSorCP2ul
A4SKs4b18yw7/zVYH69MKaJvAgCbs8OrgPNqSNeENfyd+GXncz2QE39onHLLxGOu
PmxYziVD6EFq1N/TDXKSUxAen6+9X0mbLT+jcBVqk2O1SlvnT2Q2DItVq1FL8Whk
qSV4/bVMCoulb8MpH3snKmjQ6MzXl2NQwszoTeU2tksnwFmhly4pYJXblFrG971B
whYwGIAc+WaaIBw8AVNm7zB3uyyMQlVDFC7omzWqdKQaJEg3pZQFX36EUT+EorDV
LsYGnafmAivUnoCxOr85qVYkdspp/mWIQR9tfiOlWiES1GOD+iKoR2ytey5C5m2Z
GY6u8h4bZACOGx5LgXvqM+Io3jstqqi27ElkBAk5Y3scGzLU4xJ5fAi3J/0O24FK
iNDsNGVELZx41CUW29hLSSkXsqaFRP9tU9WY8SjxJ5rgWerBuGHe3JIcHegju4m9
FnM51imUTLmoyvXAR+OxHcM9Cxc3F/vdUjYMRRurcAXOf8k7iKB12qS3pOOQ6Yxe
mzZfugO/YyKfcOiukf1BzrYTO0IKqps6bRcUWR9JPDmYiW2DSfGPG6PiV6FnixlW
xhIx3bH1yDG+kEfIBS96CnlpM/HWfuj97zFS6DWiiQf6hNoq859Jj7X15D4cRnuV
7/VgvF8rDJnxHJRVNK/vTspPP57ujd9i+TEIgQfwHdGJeNzogOdgOXkC6mFUnwdU
eoKASK+/IzAot81J5To2rqnRConB2zrdM/UWss0kuQtpNTPdIpB9BYn1G42WDA6F
acS0cOjdZydQ73ATl1HqV6aSPB+5bgYMoECbX85q1DQ+OmYHHp/IAXZO1dLOIEiU
rXsiFfx7TWq5pv21utDa9fot4mfr03dYe2CUE7Dy3bTRHQ5aX4Vs2ZEaLtNz09PA
SUA+PS62JLwgqVIOcX2B/8igKJ+29VPU8q2S7N8obfgd8DMcR2sfWWTPWi/D7THC
0rppjX4z4ymSbfaXxlnPC42gWlHPOcAsHl3ifRYPStidE9+EOuEy74VPUUYI765N
qxe7gPdWwKmCn4sSNle6KEeRcmFOOWHlMFcyBK1gk6N//Xl8wISD+zE0OGvQCR5f
UDEJKetB8Eo4ZnmnGxz7RttUr58wxq9Bqw7XYPq5L235/vyy5LM3PfDOjl91rboq
/NJidABNu6mbcxj/VfcIdF56Sqem8Ea66z9Sa324nkwvY3qvU1Wivw4scdOPJh9v
ZJCBxGKt1uvmH6YNNhu+tdgpqNXHso1Q5tG0nV1NXjVppISUOtlkQpHkVNNLs0To
0ERG0+dvc88GrE/UGeR78ISatEuNCP+k7IKhKkqjxlWYryG3eJHvyL23xFndsPna
lFtvcgTwcIfx1cgBFL4EGazARigMk0I+jbw1C4l5O7pnZoZUy6Z26jPwZq4hr0Lg
3lPJDQ5xAIAl7MD4qL9771IL0Gpdx+NDT0ZbXMfE4EeTIRni/CS3TNBTShfdgS2S
EGjv6wL3mQ9vE017BOeTYzbGstAOZ1HGo35Z1dVXJnpRJfKXJ3SC+F9NpcoH/eBU
HTmeDcwlF15iscJltMNbUVX84kpgJZctaQ+YgV3Gy9z5Kmw3k3kJrdbD7wilkwxB
YtYqoU1lbYwIDtmEbVaKn4Ffwp8ZHrpybAPd1TjBH2o9kmZbcc03LISnYUHQRpnl
RDD1gOmeQ3otwAS2xy94QoHlimBJteB8LWJnLNZ9ceJ1zJnpn4sxE95nuszhkvmw
ou5q23hdWcus3Vmqd8ZaR2tfreZqoPiYkav8Yt7eF1yW6IBrMDzXGyaMR+mzf7se
mc2CEZ7L6rE2+kS+UhqyIEdVYTj9OGEZdYztoanRHOiogR2UFh7R41dEBaiJHI2H
yjfUvKbE3PflQ8KUyYmOSeg3SMvRXkuvQQ6OPpU4uOCn70Ls4c1C1zs7Qi2Qdkmr
4NQkZyLAOYI6+QAA16AZWO1cPVCEjRLXhxpbvql8DkPUz5/jK+dZZtwCJjGYcRiq
pfJAfNVi6VF/QA+19tEEhu2n5SVbPc51rgyKQEe9zajDG5MKWn4dRgyMeeTZeqbK
MTcVdtbMpt/cu1h2rsOtc7HIMvtLTrpDtpvqEuu7XD2uHUtqMSMA4hZo2oQB8jQw
mMO8QdFCe4Vr7gJgmnOqgi3snS8CFthg7BoB72mBZXMBbB3aFQ2UrV6A4l+b7Sp7
Ks+LTO36KqAIwVDY8hdsnCmdkH2rNQM87J1RNWt2Xl34OHyZtaWCvvBz6/i5KD9O
a/wpZWpx6BNxtQ+DGv2M7Bn2BVZTnS4sheAKzi8kc2nPoe/SgXI8q7pj3979Lkgw
VzRcrMF0Z4zNuEll5fUO6hqdSmKxzlsobUVcX24zkeDnxLkSohCjp9FY7jHwFawX
skpq3t3jO8ODbmgRNUzKum8NX8a4Gb4ADK6WZNyiZeomN2wijBd/z7SJowqo85ra
fBd/sPwIxGc8vuieGcO0VR+RYpeHvvzia951UwwG9OIpQdrqmVR3OMbwtPhLQXPD
Me+h9BCMtbB1Jx+EG0ZN3NazdB9LASD7SIfoXhdlKuafvM1UadTIh1U4obEHbJlM
KBMB+TY1wcBZBtufJfytl9gaQpRJLSL24EhkMXylq1dqfEmGdCWk3geAl/tPyuNT
moW+1EEEHlfVjfEH8o1Aa+74ZYgoi4j8CU6PfPmgfb9lcWP/Vx2tDngpHW8XCeEP
UprnkGEh/DgKqb1FBSA0zcYpAGVl9hzW1f0Pk1iXho7AI3rd4CBOStUUdZFui/fi
A5y6P6XGcOsfdWQ+/arH/C6AnEY5dX+vglndQpxAUT6oArxW0ZyK3NiyI5P3Z62A
a6T6Y7zEPoN27ekMGwNP1T+T70VHqoTaVkst4dEYp+jcUCqcOm9l2RNwoZvldQVK
75uP0W/iouj3M1bsfL0fDNc1MJ9Cei3RArnUaKg5GmgnRlX4WDN5LezbX9yn1Esd
2QPZuTskU+GwhYTCCDCCJT3Krv/d2toHe9a3CFWg5rIP+gSCT4BD4z7YYtNTbc4J
1m6zXdKYvFH5TBF2JKSr+1NODs6eABxK3cL2xNyHe0dBWm61izD0lk9CR1CCM3eU
RDUoHtyi5X1Muv/s6tuqMBIrFm65n02bZVNJQrAtYoNcVWGKkItcrTjizhO5ofGN
ByNm6JtZL/TyLu86jF6ksEvb+5Zi97JqbQnGrhu35r5SXPDPbMDbfTox/VB1Ss5W
+MsOy8vto5iW3e8Z+6OrV1pYohlhDSgSZ5VXyDAVnnh2NmNL+CpQnWJI8LGZdqYy
IrWyhWN8PE6++QxSUogsOtK7opuNabBwhIrmbRpqkeKjfEuWfhL9m6EQRtUrs5W/
dmGmMxwsAOmWe+s8LqEtzSha8CVsLEgRUbUkvdjV/CT1ZRPNizT9dG9RAucOeSiH
kfcum9ZNDTdr5LaKSnXkO6+T5/cltSMTwjZdHTOsTCCRi+XT2URDimzVHgbWVyKj
9JBk/UcfMS+YNOoJiOKbFG8cEki5mcafUXMZYUxtxxpHp87+1peEjtxmjFcAkFWO
uWleFJMpZ9k19Nr0mqKjGjpbPmRDOnD4xMsRkXqOakDqjJd+zjRKLMSfumP8ylIb
MlAy2RZfY1TCDtvJ3jK7RGUqdHNh3zXGpwudn1WQxaVrXecJZUop1XpYv+Gx5xSg
pVAywuA0O38nBZ7RDHUkieqRg6O3kqM7A8emn+A3Ykg94cShr5zCEDRgh/DKJiiH
31JmAyr4rmX+4OYxT9ykMm+CW3kgdq4V034lIOxb7cUFhRX9x0qeAaNBb9tOMCOi
xTpJP+OooJNCRjZgz3u4l9bEafOAKDNFUDAa4n+luxEuP0JIYDQXy2LYCFCN5upf
0954CKY4wfBiB+88RWdswmKXx/6IxVRkU6MdxFGwqRojPf0hYBR7HCMYyGl0iezl
PpjRx+pkJaWZwJyyOoj+zSjp+CqjIKDH6Yyln2CqGqDwwXsL7iQFbkg5+3dZEbYH
s7OP7maPjHTMD6a0DKx5eGjHy0R6V59qsTWWxTkLSqz7Aqo033MihoF2uZuasvOm
aN8+WuvGDvMO2oYAFJJ4x0cWIq1adkotRY8TJZWFLVcyHr98iu2vuCRCFnEGTK5P
45SbZpKKbfjZFgOerLoFEw4FKS+1T1VPSZ8wJrteCKdwhmxAeOkKPB4P/153RA5a
uSkHKLLlEHT6NQgB3sZ9TP8TVgh3VUHT16i5EWEU79Y8NVg1++ShwHBUiCTPRLV7
iVLK8Ub6apMIePzEFI71K8NTj8/8BGHJQiMMgr7H8zXCxYRTTKUw2l/jNEbNhPpk
1N0bg3OGQJWjT6U0zO1HIBHfXu/aed9bYXWphTTfsYyE0Pi+lI7SUi1q8Y4tS5xD
uTp1a8lRHHoeTUnZCWeqAEK59I60WvpGo6sTZuJegq0P6zMW//ZmnE1y11JvZUJ5
PqlX16D42itm8IfJbrXIC+ePTLD0ACrdxi8ls/vHt20nYxQaHvBuleG+yyhchY1R
b9pEsY8xUprlZT1304zdxTw+qcro5Mab+dqfLCghhbyoacWl8HavnAI9ntkLjOjo
4A3twJZDE4ttaMHtaXZGHM/hp8wGp7BvKPZfXlGCNUf0DpIKrkCq0+AtLetwEm1Z
q0aE92FlvCMmMlQhpyRUyLcEYur9114fFQUavbNLj99YfI44axh+beurVkuRRSAb
WeCbk3Fp0K6trzOMtne48Idxg+rV+Fi8z8xGpBi6bne/nd5/2BnOzb1sISkc1rUY
SqsiVcvVcHcDp9fNqDWtj16HugbEl8liA+8HZSteUpWTveUuIeHU3uYxrIms0YfS
mr79q7bsq95CLiFkcJ3osYPLDdkoCXx3Or2/vxaCWAK9lBJeGYZvy8ZyPjeFoMUZ
o2VeLXRdaZNU+Wi3rtdCZnYvVMZ52Mq3s6VvMhL1leDd7ALVDL/auwWqq8Wxo/Fg
PkleGJRbm5W5M9C9zLqI/68XnqsPvbJdkhT7nnMgFfxoiPwkQ6NY9VpWuW446jjq
CFoz8U/4aWuEM0mViKPk20siTby5LQ4GmFCRfC7iptuBBPsGOT5N4lSwz45M/kjt
cT/6z+JYm2l3SeK+YeEzaxCdXqY7/rDo70v59WNzZJSe04G6x2zH+09Q/X8t0zVk
YSyyJRVMexWKLjFPcCBMPA4eTDoFDqWD/V4X5JP5x2T6ykbZxBDFkRLVv6enc66x
vFPvdEUk3VKSTJgRa0R2ssuogniuYwya8E9RtjwXAypBPPK0S2MEGz9D4fmJW0Mt
fqeSbfYGLpPxc3IDpziOsEqbDguXvVCaGNzkewR7L9VmwvVkTwYO/Bn4uK6n+b2O
fHL1neRLqQ0WTqOABr/kNq6GEpEqslhDHg04iRADBv70suc/g590ubYxKKWaiin+
YWs5/bQMdEsuZxG6pRQfpqniBu6ae8GUy2nhAqpwiBL2WrIZCqSP4wsbKQFCg8Bx
0hhKFcGpQL/WlmqfAGRaS20kK3mNOxryM16DK1W+tmWytgaYJh88fMJEeKKD7bLO
UUsfgNlMdCkUJSd+kIHTYp8e/r6aVQP9ejoZcOQdVMZL/1j3Mllz1sQNTtBzDCcU
l1yYGBYG3PXRSHtb/ibLdQUuujnGA6oKhYHLNi1wKxSbTJkn9VTNoCkPOFQ6X7eV
/C9PTjrhGjHv3s6eJ37PMpx2bR6PCAmZj2484xUoX1llr8mJJqX9M5qXrb5GUgG/
IgFrEBJHukJnTB6C5FN0PVGhMlUfBbwSL9qcJR4YZgbUFLHTRmJOuhS9YeA8BWLs
MmkWwAvoPOasFFmfuTerZrCguUVVrv4PHfd4oc/rrqu3zkykZNbalAvkgpgmQMbC
EQmFmtuEkWSYWqq+qkyuWpQkfeYT8oJ1zVDhCqbcm6nYYvJXXiBoGothomTCBZxl
zh0vjG6H0u95SXrTs8aH9s+s5txxNy+lEGjUW+zvVPJkfM4iwtQ3ix+9KIzAx8yQ
3Bv4yB/tUziTko3idbMUXoEAK+3iX9Sd8oRevJnoF1z7jj/ZBV46MX0ADMEsUdnI
JyeED7BzAPpWFS2NXOqIi2E8qGFAwky9b9R9ZyQ9ySieqTD1fqWwWegaXnH2ejAG
XmxZbo5mjIC3PQc/6xz/SJQuejUMGMU/E/imSY1NUgGNqxnjy4bcQqvy6X4dT6AZ
vZw8HLKOaWMakmGIhIJ8TyBYJm6ICPApuIaB8zFsHLPA/WwQ6qaJOsIt9zipY2ZC
Sj4gdnkhoYiym1IoSI6jFMxC0zlCi93Fin++8lyI5byRTKKu7lvSu2iwPdPOJuC9
e3QVU/PV2iMQ3Bu3jDGIa6iC+cGSV7LmwouCIEThUVYm9pXyT+w19EXgATlz9X3R
S8/vLbIZCuEBQcSI82rM17edXqJHmIgKnw3R3On0iPK7XTZcSKfxKmFmMPtIDt/E
4lEgcvuP1hlRO2pszluWHh5dk1dh5ATXU0XkuIP18ZStgOrmesWl2nVaOCK3I5SR
ZW+us5bTRbvv47hOyEi+iciOEWMZMMRRw7JV//KebNG6NCoVkb79bdFxrfQcCUZf
iT7mFAvuZWNHdGYxtw7muMQg/cjJwCLzTD+DH2u1rz/mAGmfLg01b3VaLQebM6LP
wWXbAsNF+B/oww5KXKUyHvq35dEaHrxRWuDSkRJIeWC12GPK7bC8oEhb6UCvq/Pf
ngljMiIsd7OcoAAj50Hg8HDHWDJqCJWJxqzF030UPuFEuz5v9fjv5ONjHL/5/3vl
16LiEgMHaen7U6XRIsta2qiPrbd6J2bw/dMe+uPA57OuKmwZvLi/VzkwyvLzugMo
kkGSGsicc1pCaNxO3MKoxHKn7GmYZWLmexsOp2L8EysVZxF/VK+bQIyHptLaclCa
5uP0duPZhgUDC9ztwT+b9pMd9I0OQo/CC6Fe/SUVHqShRQxhz6obtYQOUFNRwTl2
IYN+3MeFzjsivTg583W4yk4pdOzV0r3ojUyyNJxKToGUZDFE4YNICShHwR7vjojw
xj56XacRUW7EzHr22eTQDg4ADq+YH59RLbBNa+uNYqOLuszz/uEhNmd59IZ5jNLC
4TLkw2Qgzk8sMRtPnLMA8tqKFrrhla34WJuRPsHrBzLGix0RaHWPHNp+G3lJRQ53
yYQ9EpfqwqDh2LcrlOmSTHDqLIJ54DyoD7OtwUSWTdB/N0J8f4DD4t5yOQr6+V65
FoTMPsxjznst206UJqr4GuZ5lIiLSf3HwuNT72zXjC9eaTo9+98Q98eSaRYmhxvt
lzg12jHmV9PmkdRYfBbAcSRywn9cUbSI9tAMB3jatBacaOskwAbXAgGXSd8HrV4a
1ueakOdPb3U1Ave4Ct4wXe5YHpRVAIxX85L9ijyCJRK8v/9CEDNNk10kdrz8yKvY
Xe+cjVMyfORxDouGYo6c+IPZUoacV1ucm7Ixktq1QMvNm/cDlBUV+nZJJp5/Z9/B
1SQoxNjqGZ4ckOYcJ5cAR3Epwjl4Y7MAqbGATq5rBM89leBL4dw/sY6MqNlNKvTj
H64jeC0swVxLM4yLITsUqFq/wyW6PlbPlVKdLOUmcxguv/ChHCQFYlHUgMXSSzkZ
UnBuyds0rysWpSxpJ384BtgAezS3N4wDHcIAh/tXvOsiCae5DToPfOKT62TIXCDn
SsM+i2opjrkWPkbsrCk8tT6Ug6VMfevqCka/ss5tZS3BMZzul1cQxrdoJ+VJSeym
oQ1chHclma5QEI16xbH6z1phFarlxgb81pwLlIiab+nH00Pl08d+6ebKeZ92doK3
AiHqZy4LZ0lCKhnYcCc8H+/RGFJPc98mCp4oMOyF91sjZhh+rkICFvuKS7V1JaKe
GKfC0xYiudU3Klui7T3pl306EYdpVBmDEL/ndIW9uHYeQOo8N5e9iNsnIUGF8vnV
xqCJ2ST8/YWKQ1TqTn95ShY+n9On7jDTLxcmAMP24FyxxpO0TzCo9+ntanZL1yv4
E6sU8+FMLdehxkjs331KNMY7GfYJDBLO3ui6ePb1v4l/LEmoHUFEd6spMptNrBXy
3SVy3WUEgkJPII4oFfQUgBeFbVE1xspj6t4Y+vwt+UWA42LMAGsq0yRt/Frqlfm7
tPhbB+GB101ohTjLVV7vK2w7J2Ca9AkJHxlFv/gMCxczKbwZb/anxTG2VK2zVCmE
s3c19o1Sw7lly+3jYpMQNsV0FZhdA6h3d/nG+qbImbpi1oz0ySVPSI+GdHNpHCcW
DHOEreuxEa2tl9VNZ7HFyZ4lmLp2+q9b21OSWoLdxKPR707KC5WeDHE9/gv24hAh
CDGPNNdcXdymxnW/7SLoaGa7RxPhH8RS0fNVifPFcoPDtaKBWVzTQKkWCmkWEeAk
/CwXPnij4hHYmNLsDzsvMIRPkrAXDTns3qcHNIbGOHAf87sHgDZ8kEvwWoOjg5+D
0LlH79Oll+pxU+LMjBFJcRNyXpnkvmOTNp6K8lccpuy3AtiKeCaxOxwJlHCx4dbb
AKorWIw7QoIobqDfqzWFMHq6owif7G1gl6hJf1T81BRx04hEwaBe8e1ZXJkdJIOc
d7qOzITL2FKsl/6DTVUX5uUBJxqS/oCs4K7vSLUNW/tdZdVAZZXg7rTgNKW6o0SJ
gB5Bae+WYGNHOamAxaFRHdCOTCuWYFOQGfxiWRsWtCVly6XZ3f+UoKyUxsK/9Qb/
sxavJg57r0KuEE6tfbxjDSoxbdrvUNlO6cGT+Qis3she/TQIbCh1G8IEvHbEhJJF
B0eCft7QDvJRKkOyYON21vUwtUVzLZ9HYSZ4rsRW0exsoZKH81wR357IGGFi/T03
CmibJGze9Poyrp9FPa4rRXgi+P7ePw1OPiNXYVeTInu3a2qhxUq4lIMphskmcnjV
hAzNVVMiO272Srp7KMOc3lLzBb+VdWlsNJ+8Z8mqYzHEElOmqD7HjhfJH3Fq/+Ms
2TJw+S2mjItcsL7bBmaH+tR3LeuTcQuCwDrWTy95lorffkOghgeEC2J3K6zxOlCP
ksK16Ps6vHjWytVyH+8ZlKrhCoQHMQmpSv1L68Jbe/fKJAMv5EKrENXTDXcQ89bQ
Zp9SUxDzpcY8W3VjOfFbGnH58xDgaL5/ko9lLhgmzU7GiYb6COsEXql12RDDi9Ap
fCcHEzneNc0prWAbekMV6FafVqc6agUl5Kpn5hqPeX3p8hbPK9ubQZnfR0jc6yJt
32pBHCl1DtWB5eOXvxWDufszA8Qm7AneNWVYT3yzAROkHT9/ckU+ozzUxx04QR70
E2Nka90UZObuFCl8s3IzCXZXaWeHOTrkJRDXlW2fVzokB0rj0XLzYuIZDMWRbKp2
xRGfrI3maasFsk4yBy+/+qPq2vzwipQgAD0OUGXjEsaRQwRfTYssZ7b9WpNNa2TS
IHgYM9VwC+y9MqpxefRZpTqjG4BSHDk+kU2GIaRqlNd2QV5HpmBD7VlpYCPyV6LZ
nJxPdGZY5OF/RME95MFOEto4Qokac35Dz5aHRCrS5iWt3ly0obYU7GkaSa4icI7N
zamOw6Q884XuxA8maBT8ZnW0cx4+tPTVo/hAUUO6lB4T+lYWGgvCjDwxvw2yKeOd
JssJQFV/4l21MriZgPv4csuswBdDDZMSB2ORxqoqoPLhCkCp67sbPi5/Lq8kJikh
1enqeQs9bZ96XKZED9fP5EHORFo7muHuEkfHhHG6uoG9B9A6R4twFX+VYPR10j59
3Btd4eR5vTrxKWg3hpKStySTHNAo5sntVLBWvW0OlWDNAa3nu/RHiSVm2ibM2YX8
lGuW/vAmpA2j/3WWuHVNjt0PC1lpSAWihXnoJZSWzhRG/5NpsVgJUKXc9PLGcL/M
l6diiZ9mPEpGHIyEcjU67NG1uPvN59wZne/Hfz9CGcnEjXUA9n+amTpZSezjCDUl
eUJVNewAb3gmTWI9pxYh9/96lWsbfM80CCJUY4DPRHo8FxDhKScYNwA8oAHuUPDi
lVkuYeLNO0QpaqFlLy1YsgTGl9d288a3gyvnKKm08GFw4lxO01JRXL0zuy+xhsAN
A1bjNQkIueOVhOWUwXuq0B6IVTak0EB3Ma9digagwCbThe+mV+7beeN6tL9y+3rp
jkcxli/nMb8SrlimDknEPeoy8BAj0udIHyMjc8dad4tdl7k3M/8IZiCwrNe7Jr76
Uc8i2jW/ooVzmVBa8b3tcbY2hKVXVF0eiX44ez0mYtpP4tK92t7ILdQvhxkCVNgl
dCYIsnVsqHKYPtji3bTF/fjiuKRVUknak3D/oj2JcS1srE3bBwuwEVQca65hnBHb
AoyCWayKPT/owTKdF6ga9k3E6GV5jC0rh2ExwuQmgPsIH2w9yiMYiypBLi9Eq49b
vrwM5Hi7GmZmnDIw8COt9Hu2KG98nPighieG4rjO/nElM6lHCFXGObk65nx6tJIT
JATfLu0vYNMohTX92hbGrssddEHpXi6tpV4Thv7KTS/pkidd6RQ106+Hf5DfQ+2K
M4SIhoZsgKvgRJO6YxPzaVhiU+vY2bftQ+w5qjtJhe0xdJGOzHlnv041MWri8qNs
QcPR8bwPAhCYiOo5T9DCxTvQ0Av0XnhYVMsKQ82K+D6K5u7kRU2MQiFNu5qJ5WCi
bGHwOEPnQg5W2nKNzbDgIe1FcLPgs1b+YTbj0P5NtdAn2DUdZEfqVKDVbpnXihyE
wDKISte/ouvoDkBf+Ap4/l8WLxkftaYND1Io1pXV0lMwwrZx+4zh+K+O5w/cNqWk
M0hoVrpnAgVvYtfILPX3gbb35YpDKJGy6fcvuwhu1seT8mpuTUH0SsKDE8EI/TCU
EMIvJ3uX+5tf7YNfj15Wy3UNf7TS1rjx0Zzj5hv1onM5LZvhuMq8Yp0bXs3K5Zzu
O01r49GG6JU0wyFemWZuL0JGkkxVKrEpZhcv2WG97CRTswskupgCD+x9azKOdtBo
zCmyzwSZw0zDCxChaQyLlSqoppG5V1O834ZMDmhL2TGgPV+GPfUe4IQgpSLTpvVc
y6EtsNv/R4hLu0rSGzvKEKLfuA/SdygAjp7O5vLpL6Eey1GfnFZYqZBW0xmIzZLH
X2/HK5b9OxP7s7OJk3M2gYSwiveNzmPm5bOdbCF7i/pf/6t/ha80CQrTsQR/Flbl
zgbOta4GS5xHlc4yu01DgiIdIWE+l2yxPAPO1qZegXm0BzScN7ZwDdPhs7d6QkPB
gcBCDBvOJ1i0gYP4TvN1TYqewTNH530x1a6RG1AtJNANeiO610zZboGGIxax4FXe
8A6dCS00QU8pKvQMgjpNm607toKTAphwAq6D95N3QAX4MsnCvNwJT5woqpWJ8AhQ
gA6sBfLqs8xe9Wme0kMHyU5DEDzPLRtbj+2qiOeRd6b4nPWe2XGwqtG2lHpZI17s
osH+RbdVzBtaHBw2Ya+Qaql27IzkqvA5NbFDDA1sKZDYto9sIIz9R3tRIRYAYl6P
4L/8Pzt7L55YkoI8ghyp6R57ICHJHkz2S+mPoH2fdUvs5h4rbphCfHvyd+4lhWsL
Zpqyf6T1eABHQlzur1PuaQ8UzkFylSAzl/y/eE7cKDLvONBL4713behnKZVkauNe
xXlY18qJ7ocTqz0g4b0En0M1BFWFDD+qiG423L4te/rgFotcFlqGdX/z/+Hs97am
4HplaHGpLK6hC184a3LoEhD3GiPy18ELjmPQsbKXeSMWNtnZVWPgPFifQzUHt/3/
qv53tuMNbSK2bbqRcX8M4oV82tHKDwsXpossAVVONNM8FtcZqTAa5HGg76qdTYIu
AY5y5P8z8n+Qj4DtPoaeaLSwWdm1pQw5qFyYxWtnxtK6tbX3KHNxAbmAIs/rVqUZ
OTCdZJVii+5smpqUa2b4qkLuQE1uNvPi2pC9HRdcOjB7bz5S9DTQvKbKc6OSCZ9G
/OgzBdkx3wZeTpv1xUrFPdjy4UyEzy9zZlGQ1KeRR+1KmD3gbbIDST8vvsWoi9LP
1/DXe2M0XfX8lnH2MCj0K3in9vDbCfqiglbGSgXYrODrDnTS+ebZ8Rc9spB6f683
I9t/dP0g7mdZZPGBGYt+FISx5r+JhjQZvp12R6zACkn/vtsalw48oXu6EammtFaW
Xub1fUo36mKSyyzkaX+XuKW5h+rDrgt9Qidms3GoEajaey/ovS+EEhes90BpMn7D
75o/6S2jBSXQokyTlOaLqgy6fMrdz5gLHOzp0i8IbrWujOVNBeLNQH7aBuUl7xyv
DFNOYf4eRthoG0g1K1LsuZ6wSV46CXnpYi7LYlPMtOrkEiJPirTkT//NH3iendML
7ht5ow39dxNKQRDExm+VgI4SklmcEeSruRHkpTrOG857utqJHtaiDj4ENxPsATZh
nyyrQ8Iyg0AO4KyW5mSF5a5wayxdqSPfjadD5E9jDNkiZBhhT0KGts1F6k1UAf7O
SbvVMnskrA7jqjWHVWMMOunMAhe3gj9z32aEjPlFTjR6qj2eRIKE3QYSCmO2yLLb
tWvptFFjckAsU34Zslx97Bj3oC2i/bHWply57dBr68bbvc0nxhNXyBEkQ270YUsC
yosbVw8ixbV26FtipOJBBuPK6+qHw3U/xZDD+zjPkCjJ8Vs1W9iM5mVUd0TjLiAG
Vk1pVc2W7+mXQD6CLGyxVFacaQr5UDjjU+0HUvHm8NX7ckpwLYRygehYcVgaj/hi
L4hXLqtwhQL049hToXtzvvW73WU2VfViPhvbhsIOuXiSamcZTjFoqoM7E/q3uXun
RM6fDkaQDEishfsoiH6cAYuUA3RVCXDt5yxQWj6Cr/tKjLqBTZWk2wQZs+xxPM6C
c0gnxSFsQzYnmZtG0/U7lJ9F9tv1VhB2G2X9CkExEIXE7Fl9d5CeEVEKe9dwVjk6
SaY7q48LpaJotlm2sUc0XLaMUVxv4ldsQtHqYhCrtmH8mTk6VvcXdOH7pYhR7rb3
ktljnUb34j9Xum6uz74OlCqCfPpo4IivkSC3LHTJWHwp/kA4mrUfvzRhe0DBHvd7
SLzq7VVpixDxSY1vpMbi7ch2Lp7taSMlLfZLmGv8oJrHQdDJiVbUbqx2naaBaalD
aT9lXLE4JcUTFYd+KQef6WtNj+SsNRJNRQd7Buqg5czmcjViX/SLZXqKvQOjNAbZ
OKwv+Vg9uI2BaMf4zMshK8sJxcFOi+D7QBhCAoetU/aLQYhACclr+qMYbvgRk/WI
w04PLHpC8M7c84Y8mpyUQJV1ORuknjxabMl8+FzLJsOz/ClBNgp5FLAEOyCuH4XF
O8yCU1NvjNMuqLczBW1QR9T/2+lTdQ9SW2j3QU8QMQaJ/fbVQfg3tsjWqk1RzDnB
9TVm69ixX5/RaLbHx8xSjQl1qTSy2BJz4SJpMKRuO6/9GlOxqDXF54wsvst+3OwK
xk6uYGKYqjCIPbkynzX0BMPdywKYwfJunpMUTqaCK8OIo8CBYtxzuqIb3V2sDYiW
qC6w5jsyweI68YegXtFid/JoTZrdZ2mzdrBHYxCcUvNDA0txSPGYq82fpKOeVjuD
gbL4d1zveXZdBeS0UcGOgbuauzu8ggIt9hKmcqVHrYnf4FAMqZ6BxjLy2KbpHfrj
9Pn6QlwxiEcbl31HDIYh3XJ9hjQIWkXfQriYb6CSF4/0yg1LTjE73o90ddHxrovn
H4DH7ilRgic07RSg4sbze+LSr9aEGa/sk4dBe/EvyWgv1eFisv3X2XypaXNhfI70
TR9SBgB1RrDycNcQYA8R8HIkI7wXBD8yhJ290Tnb/pcspCuUUMqxXtGT04bhcaXd
HyY8F4RtbKfuvgSc6gI01I26h8hIBL8JMsnFGJqtrs3qO4lCfrsY21an+EOGCl5I
VrrGOBkz/tjjrK/YIllgNQ1iafIypQSdj5h/OxGinoBAdjsylK1BV39OgUlQwaq4
X3E1SWlpIKpXTffw+0MGmFfkxBYSBF6wcV1FmyvoP0L5Zn/8slKTIt1m+AZH3qzK
EDfuy9H8D+xqDHNWc6JRNcFtCOSczmc2mIRlUlr5J2nTDiI7XtInWAJ3ccmW1rHJ
bNrTGogKwe3khk4l1QAHsal4livwY8Ni6cRUfZZ7M8gV6utbInZQD0vyNvL4Pfg+
1m63qzjfTCv0fsUtIrUTQjutVZlIH8PoLZcAk6nbnmNZtW9vjBsRQtT0qlIPvkJC
UzBB0CfNpUxl+iRgCMrjOTywwHjWa6GXzWPhIn8EO1aeNslCXWXZ5ZwOLJiXmcEa
jtCphrypV/aeKHKaGcSgFaOmoKe75Sf/NkOeaAxD16+tzVShyc7mZ8D4BQuiEMJ0
+B3WeGB+SJck0JtsgFE1oKqfynAoZkiRegWEC1i6ZZgAvH/bhn/Kiy6wAkphY9XL
Hboza0FPuUqkrr1gsxJJQV53ZFhe//dryKINqkURYNd0YpkMkCLUpiuegyPzRoBi
6aQUmHT3sly+Mz0boukxP6tIFYBMXxlixgfjjiI8uFe2EWDaAp9dWNMzetXSa64j
dSJkxewpDMQqZynl2gnmuN15wEqNxeCxBcMtwyNCP+cI4UhgqBwXrAiwFHdPGZsG
N6Ljfw4+Y5IixmPWcnYHaRPBu0uUrZuy7XaY/RuDtu4k5Qduue75GA1Uwg7X8idF
eUqXrgbstypeTgundmm50YuUU2yb0yNOXnnyRxL9NMy/SS0WKQmRTcGAIP31ukpZ
i1mY0DW5N8xM0ceAYcVp5Dufz/4TWPV5IzZ4EORopOD9Xqyl1lbJVM50kevnc+Mx
sX+jA20hdokgNlbGW4M+S9sSbgftiXarlKreBpy8jrXgTj7njoXjgzklb8bjeJBo
U532ejDNC1slTewXVobd8y7vbdV0XSoTgVso/R6oAE4j7kCL8NNXGEVpyw71NfIu
zdi/eov2U/I3m9oBUqeVJ6TstbFwqlsd6C6EFJm4iUzBcHnZt7vqUfvK1WZu5gN0
QTmvqhXie3Z6CppfbtdPE4P5oZqxfXwOW/uMFwz4TRX4kDgrUMR4t/xu6wVsvqTI
G8c8Fuf9F7sP+uG4Yx8sIahWwBtPn9bupe9djU6i5fB0N4nQuomPxnZvoxcPMPqo
SqqDQopNQuZVcVRuBLv3CuiSBYDvckRWEVUKhpIwVZIsKpevDeuc09cdbZI6blPP
73n+bWPDBHXMptsTiz+6w6PplpB0IhSv97eHX64E5RYAwF2rT0bahb/XqbGFsOh6
UYDrDiBEdpvqrwI29v79iIpwdOLFtTB+TX3uCbx7fUkkeXZb6iVpiNb0mYlgpIvD
tDBhc8rPapyz5FXDzX/p1omrEzdOClo1cP12ByWZjYc/vVq+42UCajjke+fWxjfJ
m9Yq915s6sZJUSaWQpf5heISrzWDF9llWF8Bh/rwMF3drD5TXFTJ3LLB7Omoovxw
P7d11Mu4YfCeKs26mxm2+FScicIFiKRMxKLTEA90viUu1xhCI0BLp2IahShSgaDn
QevdfLs22vnyvN3WV2L3yOEWt0n0uIgN7lHMpQksv8VmVVbAb8vGlsCt1gjivVej
UjndZXgzCjb631irz1AViPBCrd3Qqo/MMEXsLkBr+ozqD4851HhiZr8qJVaEWNyS
YGCEBHkreNpwKsEdLJy5/TJqGCvHUgHS7b/p40Kx2J8GTco0UhYnh9MRyzfGzG9A
MAl1NnQVciDuXSD8Mj/WpLRHuweYejobiUyu1fVz+zOIlrhC49H3hFd6Y7Dr1qT1
3Z0pk1tViKt6HZNIyQ3BfU01KLFvyPS+IKEK4PHzQ6oqxd61JDHdqC6Q345DyeUv
cDXf+c038auDkmUwUjW2e2PfK6aK+CivMhGkd3ZqozDdE4chfc3gIU8SJc5bqPg4
8dpDU3txgKBQ/C3duiFE0towug/nDIkhXa8lQo1XJFN/9tX+e9OFv2GITk9eNYTY
kedjxQRVXjo+3ye92NqxoIKeRw6q5bkMJLlIpmgQ4TqEvT8wd0l7YwQwntmpQ8hx
VMZSC4VqbBWqSD5yfKjWsCweykTgzN6VKdB4sho2yxqtxu8UODoF4ztF8ktEMmoR
Mgox8Cs+tTvbCdOMkZc28vcDZyEEAsLc4IropqG1wBsvxudgOoN7m1mAKhuL952i
flgc4AS+iRPhhyWTtazjPXkTm6l1yF2HphFWw+FEuGrqRl4tBzfxm+3H3km+uyHK
W0XpPX3rmQJfZ3kw4t2cr1mJyTXAbbsiwryjQOuzD6v5l0T3xjmFdDhOo+231FlC
02Su8hVxrO+xFNCknT0JAriEYgRaJJwMlcw1sw6j7UUgl+eQuiPWoEtAnPRDuept
yNeVZS+wL2uB3oFJdOwtFGeF4awfXbVK/er4OgCo2FyvlY7T9bs8bLAKttuvsNYq
I/IFD/GufMq4LZYJbri0cgXR9kgiBZEEsIQItYmjExkw+JVMmAztNSlfHDIu4ogE
YfYCwOwNljDEvfQSBK4g3yoQcuHBiU6IRkL55shG/NgwXtHSfw4CwQV3vQK/WpH9
bALsDLmUyRx8j8L3FKqjYXNsvECgwULu3jxCdhpARf/Q5r0RPbMS2y9N6hHdZLf/
N8KaKRwASlbO0PqHkZGSfd6h6JPQT/u78GoNIXmsqhk2WJtO2dYfshz7Fp5KDETV
UZGlaAHUaCnS1/EHqBCJv/e9fECgWZ2oRR2L7YyCI1oWEtmvmdTbkkVAOYuCcNjk
77D8bZsZpw20uGvLFMdKpDqUFnlOyWfY2Oil2KEN+UxYa7vZkWOs76XwCGOa61ii
pEaMOShjhOTQEP/mjpbef9vrRcjHAOAFVqa3aVjX9l7xSQwoi+HF5XXBAnisCtxC
HHO3RwbGJj2FYNy6hJYUD8TKZiDKCBmWhPHxIEMGC4fEdjFJCFIDGX1TB0/x+87x
PV7R1L1qS5WCgPpskpkMP5h/HXMvgKbmoN5dHqwz9R6w2NuRj6cH84MTA9LkL9B6
GvOv49Bi1zd6Ayze1nC+7Hn2nd3ePSazkNjQEFiwIz3bB3iAAIl8g+KD+Zb2gnhg
kEZ9N7AhFBVs4OEhPFDWRcS6DrtID03FLC3wJYJMRPElMwxOirLF+AU8hLUGpn+p
ygcrbVmob7KaFv+aoa5gCJihj2eDHD+f7ErPg3/+fY1oIP/C80/pNU0dhMALLRdJ
cPxmXCVeloBIaiVQcWPCr1dVlh65wk+ebgb1xkn3HPcTSx/83h0+mmGMYSzzob2j
TsMeCEyizYNa2yOPl4a2Q/36OfOS7Lnj/nH0uRCR+ufOB3bZNIXIYpdGO98jTLKj
DQP4zFAjMWAk4tOtSQfh6z0bO3FcMd0hkAKJDVabJBmKvTCjK3EcHBDXJZCab8yR
zgw3HeVrcwssBd4+/moFo5Q0HdcugmaabAgcNiXPoXYQ/64+dDtVIP1jAI6YDa8q
ghB83EtSyx1b09iIcIa/cqfu9DqwW0CSPQRVBgHVrLbu15q2O3CyrUnv7n0R2AUA
3+8geHPwBhXTi/dpKWTZlgv55opbz8p65ZWeuE0M8NxW/BDiWCYqTsrZE799LdTR
WCZ4jHuuLXR3c+xxaXJI5fq8Oz+hK0clf3gns1jJYKbKsU87VXroZmGjT0jopene
+BDkWBzyMmGTe2kCmsBo6CUITu1b8TTWGyNON/hcbkYznvQV8UDMehMca/5sdtU/
0sh77K8lLCJ3yf50KRlcNsjnXw9QDgE9ay5HSni/cQn6XtUFWnvqQxPMbxO9tdYr
5G+qxkFGorSfKblevztPKkoamcjODhlyYZU96qqy3JM5AovUDuw90GvkyQw1Ee5O
HdszRpgh8oI0J6fl5qA2gNFcw62syBEz8rUUrK6fDhgLDel+Rf2CCqbBh37LlaIg
AUZgGFnvACMhJFy+13C0Zskx7AuFI6FvdvWswg0XiLSvBlF6WS/Dnq9/KP/cOUv/
s0opffH8KEru0IssM+JnyumzS+0wMNqdyEqZrnizpDhF1IAfqqXaXoE9TV6lWD8L
QfXnqWN06hIhAj/+cqJipFebcQr58FAkXefkGD8NMIhSgntv8uPbHvQ/5oNcNVvu
zLd1+GNVM2jY8bC7yWDd16l0LyVmIQIMISmMnAS16b+vXIoFqQJOLTlnCI1Tftg0
Mrw9HKkGRr4QRpSgQz9vKTeFzn/rCFpoQY7bbLEvXzaCmSqHvYdW6cGkIKkHOhUB
we+g5EGIKyGtZmbasT2F+p8225hzCH6VGkvX8VLsXPJkHDhD5GnEmP17iNzIqikx
4FvIDN2F/l+B5BTsKB2EPh+WwYJlwyICEsKoyGNUGOKRC1YzIRpcb5WLalGjRwBB
pJnbQpafjPFmFYr0DAY6UROa0a8UN4oYOThCIxFtq65j+C5Rk2D3aBknn24RLggK
CrKI3rOkv7mpeFPDD5glZEURdA4CD1Y9biVb2W8+0acHmz4ZMRT50dDIcSx+LR1i
x88GDWRlwQRBM2OlZF0yYGM+3yyuUm41Fa+J3bQOVKEqREvG9Xu8evTSigsC93jz
uR9r7IuB0MvgNwkV/wH6GcPamn8n8E8EItj/e2HJbhqgaHtIDcLCWof3my7LJGsH
1y9ia6/hoRrTBFtzc2JuWod+6yHPs4DAse5XMq30NuANGFD7E0x/1rt/OOx964VT
bE4OgZRfHxaaiPSBMpRdGnpYBqBfhaxYVUFmYUcKIXhO2SKn0AhTqeXNlfvvpvbC
Jewyw2IZUyGhu34S/KhpuOYh/x0PEFf7rwIIVdN6KMMExKJW6q3dx+NnYankgbgB
Yu45I5hf8OxAe1mrirmud1lnrN2v4I5Aqf25hyvYrghq06A/u6o3dV3wxNHrnXZ3
aJXPxhhqkFOjMLk2QmM/sFDztFgkXgWRT/Xj4UG0i3d2K22EeaUq7nZUXQJqKVqP
zICsXvnnBzenpatBk1zc5z7lWgi8zs0Tmm6CnpFLECrPkkXtO2Ptdb2aru0DJm4w
bXr/Ji30t26VRaJ4XyKRcFaQDFbTooDc7GVnTeveeuY3vtG/2DgRdSPSWDobEScB
czYnTedXvjXceBItm1cY8Suk/ANMEAKMawvId6Mdd4P9QjQznVVQvsqFIdX5SSoL
GSgMA/6k5qqPu5adrdDQDlKR9Lln1Ranp0RfgUd9IgqlLkrFYhPkvRuXcaFI9b2w
yTOiboEV7esR+RcFsv6+GDFbPqzT/OdZuThVhOTGQa10ttXhSohHGlnwvy5sh1Oz
hN4j/Ibadx7DzxGll5I8FJrMss5YI5dVonm0isupKX9m4vYsnE/B8MfaNyHMtQbV
vcnnqyvHJrXrferKq/nPWHZoW+xpaAB90fVH/T71RDHAmrjt1yNLXin8x4ImRe7y
bwJaM0QRYmcrsNWbq+C0B7u/FOTTu4mFv6SQJapbAm7Dzw7fVfiqTI681NZ6d6WK
OeHPWerzrhpSpG4bMBjeKV7bF1fV++NqRqPzXyQ3h/RBnLvEWihnrgiW0m394A4A
fiWw/eMJ5KZcOn5DBgSfJIKEmQIdo6Q2YHqS8WMgRjP23+yzvQc+Slb3fAyv5lyJ
d1989hFZirsDmT+hx5pav+wPveT79RggXW2JnyesiIw/DO+S/Kc6++SDo25PuERs
m2ufbFkJF3ALH9O+WpNlrpJ7VlOyPN/87+8Pubpeiq6sClhogX68+yIExNWu+iLt
QqBM8KSDiMXoucx4u1uWiUACNZEzmb5HYBdE/TV1fEyrclleuHtjmjUXbSKxXoC4
j/zsmYzncy2Bl4X8oPRadEGxWeu6exM29QcjGmsxlnuoIS9nXFrHcSHWP6wb2QWC
GspcYmmbCzsPgbfPULzxIf577zE/ZduQYi6dhmoCxUT75pvxyASDWGaEKIHTCnKc
9zItrM6jI8Po3Tfzm3sZ13rDLVsLpDVVrnEoQZy0/vgHx6LwLj7cZN2U0wZK5W8z
16xwHk296jp5qEkGNLR1gxRX8tG/79uzvplayRhAyxQF6rKRNfLKvxtERbU4Ad/m
Jbe5S8RaHUq68ignYa3kTz4gp08Q25suaQBkzImCO172EGaQnmKvJTdtD+F34vpR
m2upgMamRGdZ0zOoj9tpru9OITgHg85PO8VBobHVb0fr2uTV+lYfgo8V9IZluVXP
szsC2AgW/1wxuHMNzH3ma/wDEoON5mVWFLvtg9ehf+zGwTF2KwjIEhdf6r8ay29t
RTjfUrAUKQqMACF+BUClF2ph5Q5kd4aU2CYy3XFGxQsU2pCSIjskDneGT/KeYPqQ
eJjBxWjtQuFrWVBbu/5PFJ3DznPolxssDx5laBjfUP7qF+wtIwuCfFNnfO3VJ1nv
0bU+D7wAC8Fm6O1k0+D+b2tAqTA+fRlB0eXh4teRLxKvzJOPlyMe33k12QNgAqPf
cA9n/Z15KP8QCNOkCyr1ZQ1fGaoa8pWqYjgRlKz93QsxJIV9cLV39KENeEzjgRBS
xKks5L4nHVxLicZlEHz3usdCRGslhEFK3kJOEYRpEHE5ZwCZ2mdxJr1V+DGQKGo5
3anzDfOuxee67/8tNXlApeuKWkfyT5n1yWy33UMLDee8QFC4nc76WOencLh1qkAc
NNdIRx7ODMKcVGU3bmJSSQNvwBuW6Nxyrk831ST3AQqHqknHq8xW4cJMVJBVmFjP
+CytumgJ/aPPVoLo5cR031ITMVr2UPje4y/ebCjB+xr4t7pz71n4JHOnuPRwd0Tg
ZDyhNknhjtgyIcJ0c2s0KFXO7Sa3RjdpZHxxJVNH+KXkUWFg3hBOTqrRtRX1Ns0l
H5SxJawMs+/1GHhkzx/OtfUcxjR/pF92CuIZLA2CluBq+veehxAElpA9RkAofzLP
yLwsl7ngJKDSbFpD4gUgboJ0A1byoKWghYEPdm/X0uw43bFMfVNVNOMwq9bZh/ng
fEjx6KK3vWlJKnDLo2tC77ldwgnzlc9ZxgjybdW2ebjPLSPrqtHtNCwMvhr5EKdR
IBeA36sh1SQ7IVlm8ozZMF57PtIo4wqeu+3qfhdi7LVC2wnL+rKzsrq1kSE4O1ez
xybx+PPd9IJ4MndvkV5Nm2BU+w6mxayLfAfuYIN32Z2Tarjwd8Bs0CXcAsASLiZt
cd02n9DQz2ReW5/CAZ3CMM32jXI9ZF770dD7CdTr6VpQTKWydsr490JVLEHXluE+
OP/JY6jv88z9e5a/c/Laa2pHhXVan0inUACkgOu4eMwiDTb6a/iOU1Qt52QowQRt
H2WypY9t2kktbDFXKDns0MrBQ8QZIcbEj8RxGa3dxgzeX2oVFq4jw4LR0tdMdlGo
L6RPd6N+1oeNHUbKX/gPb0QnoDyekd8IGIeL4UU1yx81neVZAlrc4tdDyC9LWYbT
WjoRMlxr1sPIDwbPCoug+JkcWe5cafCex/JALS1zAt2CQW1auxWd52A8243iaKXm
iaDtG+pxWRhH0x0jDwQxXZk39yPo35Db57O+lOxTqjQhalgk6V89t1DjsFwJMNQ8
1VYOW8gUzfA9hPl489Z2g9UTyIeKu4LEbGpNKyA/z2QEDTb7JCJpaNuk6OO1ii99
BmofmGCR7RzI9ijdYntxn7NWE1XJgsiZQ6d7JvieA0KIu5RjH4Dsl2eHMjdTUFVZ
OyivOiwr3qAgocFDJDAQrmCL4GduZTMM2FZNevCOk0rxphCpHeYwgF7NtN7Tc0g/
inWMtDDej8zH4N0Ukj8OCenEIC5XwMfKJz/rv8DMGJysX26owDlJJ8XuRzigVr9D
hMoRlvpdNJWy7BQSPLWwLPflJZf/5zha4EKwzwhODh3oGd4+OsDsdokFaE83cDlL
GNV4xac6Ul+o72Oxva0jmDao8R2Wvj4SyTrm+o9VhqaM4Vk+IEIW2Gf5ZTU8p5Xe
EzkmfNwDbdgdt8R/9gmZYOVedIUxaUOt412iANtx3xL1sOBBkTrb9k0GWeqDCjOI
fXH+SEWHeCjnE9YJAtjoHtpYQJmzxh9RvgQdTNeMURgruw3wbjipML7SLVnOsRif
wIFNtBOKZIUfQD2KLtavR7Fh0P9VpydgDGiOvkIpEXdTm22RKMRoKcQBq6zRZzx2
iTzlt3bDuPGcxjaYXd98TvFE9R/D8jyDzaYn5AEzjvO6LPbiT3PxZ2iuD/lsvNq0
LN8W0fa6CNofbBsVrAUtXjpqYhVgYoGanho5y0bmLHGeqhw9CsE5F8yFa4CIf6xQ
1DHDgqqvbI+j2Lkz2XVM+cCcwUgddy6TV+9xQosVaYfpo8tjqnbucjE99fxk43Tj
wvoOYUi/69NYtU9bDsZjwwOIZHbiQbTN3hGuIqkZOUZwUqYZSbGQGRAJ3j+avphK
m6Z40xkiE+8klk+YIxy0dqLnQ3vr7v4CPN/7ZdODvQ8airzY47KqfEk0n8+VWmbl
5cq3tKwqj/Cvl0IkeWFOCLQ41YNwz2Q2uDC9VqSppO/FWbgqYGrj0uLKgBEJszDi
+5VP5xK+dZKCUTWUBzFBeb3dYe2g4Q8kKETv3lyEUBEWnqBiiWLmSBc0PdTVwnyN
J0KBU54VMD7NrmL3LqoTIy8y4f1OzHm3QP/d5s2Rwqr945i5uT8xIdB8u/B1ljSY
Cxe2c98MBXZxKwC24IySqaI3u4VLWhF4KY6uJspMcbnzchMCBLDe37N2oLV7+GgD
25LwId0o+/soafiwpV0QfM7vqX81eLpuAM6MsYfgkGm4SRKM3ojQ23OcD/FlmWW6
66zW9CytG4HJ+SF/gNCAIjfZhmTgeRA6Ni+BkPrWv0W1LD7NP2iex3L37E0H6wH3
4bIGP1F8evA55ehUmzKHYm3LbdwXhiEV5yCjBD8dq3TkNSmbevcTQSTOWHNACZaB
/dmO0Mml6eytSDFAwSeOOAuXR8RXhFtivFazWhdWo4SsF7Wh2tFOn4x5D0BsKvaH
xYL1BqZIioZgY34KWbsEFzgZWP7H74medRKm+UbajUjlnutDAVBVa5rGJb4w/KH6
Ak4ony0U8G9xH8P8HLcNetmSm7MqVyL2kvReF64yYtImB6aSwQS/WhaXUiMwyusG
Gll1JhtKqHn4VyLWyc+7NorhotuaqrnyYj5zBRjH8/CHMkFyXVozFfL+j83+g7GD
kWuNMdtSixUJDIrAI9ajsdZU7IYmOyHqEA0DUxt4zYUE7ypC9aLv17vkI67T+6fP
/R4VQx63hvs+xmyRo1wHSdC9jP0JEBswonAdj26TrL7CoxzWGHKWpYNtjJatL17h
e732a6at2Pvs9grVELmNFpD1FlyqbGmyMVQD60wYxd5gnryEhVH4ZdqES3fM9C9K
8rwiZ+3UAXzWqxgpGdia+pO1fsOmwXNjTb/LhWA/+FLyAmWLTCxZmCpbExK4i8TT
bT3v+ZxqL1zvCIe+iDaaI0TOqhlbQufPUfA/bKe/zAwVYwrtS5npxCSF3n1kzpJR
Hb3qBftmrvmdzBNBg5bGyZZBnonezqjTYUoUkvCBnixCmjYJCMtCuTfLT8g6RVz0
UKhnFUXisLYvfgHum+rnfA1unalmcaN1Ww5A4SqPvLNPb+VdrpC6d8u/LDYEyubx
y4bhcNhPxIJNyLew890zhdf9SyTkkYoYvyhWMWz/7DsQW6vAi8FjIRp+AemlM5MN
4m5FcWwqYu++g5o8VVovUctvrJaK6cRCRS27hTVX/7uo/ehQGd4z6s3Ztcf3lzQI
y3FZaxmjyuBgpbuvp1VbekBqokhWGckzx0ip4H8jwr3aa0Tqb+y50QAwNkZSSHGK
WD7zEZJAslNFK70xyqrSEzUMbXvlRrJ25rIA7pYKdnumYnspitFURJUPOUwKyqxE
cmdqnLN9CIutVXjCs62VSbaAG4ckxwJD20XTIxdCNUhwURW1muIQRTDvvAgS9ngV
l667GRyS6rjTWIHdrEvxQN6WtpsdHCC5D/MwFdjJctTg99ZpInx1wcrZJtZiBKKV
SC9ajaonM/g8aXXzXH25aaUypGSWxnfIcMqxWjpR/Sqe6VPJaM0j2X/i+fy6FBQy
Ps1FlrSfvjjgmDkZ9e1P4N/qc6dF61EV9b5gk88VplADVDQLPDGxmz4tQN87itfA
HB2Iu6tQDz7q8StKf70nmg6VoydNvuxVRmg+PHWTDqi/j8K4qAqusqFoqC+zGclA
J36qUf+nBHJLjUqz19ggjcmEFlvD1o7f5DrST/4sFgrGTUXk1rHYgWonsR9ocIrw
UGw0Nh2xWBe30oXRT2qrVEPYLn9zsAY91g4KLc7RB6Aq6YjaVM5y/fObrQ2A1fIS
+SRE06XoTVyTyn95KRcPayoMhZIYYXXsMjhahsZu4rmGD0BYojUnod61b/eRQrmY
wLrcRk7kIxp+9BhA4Y9jlAEfqbfNqCu8gTfh+buC2Vb1vl1pQRepP784y6o8fSaX
IFsd+04ZzAkhymdA5DLiRYXaD4/F++KFXKW7yxnI4j57iqiYENs1KmqXB5hxbJSJ
U3bncdTkP9eecLcl8+LWhldU2OkyOxX9+f9XYZoJcId4vb5dLvBnt48zaO56jUOE
URP06jD7kpIuyClhqDd7G0fPPLGtZR9YYA7AzkMmIcSwXwtjS1FGpGMjQ9CK/gdS
rqnZ9kOrRtQbI7vARPrHtlUHz5qByv9tTrO9LoyXaGwt6lDD2WF2pwzh4ClfsEnn
cXQLF6lB9joLXKLut+ZTkkmGILkoAr1QlG+/88mwYrrVR3q/COXAbKyYfj8yJFNn
rXnUXtJWKynh31Fhuma/b6PJVbSW3I7XMxIG4abiuOEEi7pnDhQmZzXnNbnPL1aW
8XBh8bw1McN3bb8dA2MPzJxWBgIm9+xYVUaIHhaWAED1micsdeteBBLtdrvSWHeA
h7wFciGhaioHBY6Zl6XFAD+wUEGZqlb8ki5/Azr6YejJHTyVR00kcZrI9PCTYlil
tPuBnSM1C7Idcwa0Sbws/Bj8OR6O+QEwUaleNvPMLFlRwGROa2NHzIJXxgdfMbK/
LIdBBcwVedpXYEHdnVOL2JS6G2i8gzTVaXlLhvsZaqBkbG3KJ8d25GncIT5WAEHu
PYJYXmC3xfJsnSBqhJ3P5TAuibUcGRnp7o+ePiX1YnQjlJe27bmM+7uXfExE/KXr
PEcd4F9EoaebBTLeG1uw7SQZ9kqcvqwGCNEI8sZKWEA5zhunRXstYRlSsdxO9DQC
NFkf7BJI4xOeotik7LEf3bsuaIC9+IIamJ1a+0+rHkv/aPl/5bMvklHrvfIJXHn9
45StCr6MKOBYhlF2sCGQ+EQbRQd+x0WmAdI+DKVrTt0V6IXE+Cr4HHFrjNBQhuip
zYI4T7+50prNfDLa1iGr59GH6VUGfNEhm1KBt03++1TiiAdX5ssxE6UYz9JsLwvy
xSoYt4RxAP6hkY4a0Cp4q1RQKciZN7H328naFih6lyy1OcHiRBy3O3uRV+S/fNE2
SQ9orHDJ12Xr35TudvtEf1ph2JcyHQW/ma7/04r1CI11wMW2I66YHFke5ivLL1kO
C8T8mZYjS49nj2KJgVUspk0IZssLak4iahNy8dLDY/YSytdV2yxHa4s3aZkaZ7I2
Vetw2ZU8AZZoIeS141qRwCBZ+IIjntbfxK+4z2cPoSWZWEWB7MJrrphuI+FSy9Zr
OUd5v/qW+2rGwbfCMzShX7/GcKK327oZAeUbM+4onCEZ1Lq4fGKT/pAjFaW3LzpK
WgB/BalalvYYJ8YHA8dQYK4Vz5QItQPrKmQf2O5JgOQtwMVmNi2DgqjwaNeYjmo1
IIDizGRkJNJMgXG7GqChwNnVz5Xt1Yt4EEXOF/PkFpzmqYLodR5oeRM+yumvVYDu
vg3q9mofTU0/khIn0uxzEE9V1T8CWZBiC0txmrSVFuQTFPqsfUoMYSSBKV/qd9ig
TUupE8zkdJutFvbZWZb8uiBcSwUPkxIQOTbrjukjIKMCO0NxiXXJIF9eX+ikLbJv
F2tGgrZbWybH8kTLHBisYPcW94e1j1HZ6nEWPOiUia7ugiMIzLgDU6z1wXfaQKCB
oJ9JPITaK6YJ59MYFsNnBjrVGTZv0W1ikCEcrGq4oLAy+KMQQJSS0T8qNgmR/sqf
1yi7efYrF2RZYsi9bO5B3oU1JHqr4FtBivY1ioM2gE6Rw+AM9Xm/8Kg3/ShgaUQD
NjLT/YDhAUg0FfsikJ5wZjEqCHi7m/+58HLrAVzXlPqpW23cC8MkFLhkrrfcPg1G
lbWfVmpaYRQQpMxy/LiRqGQjKTH9xtCYkazgb2tvtKyebRIuOrXWvLSkdNhpFVKJ
KsF8TgUqbqu9J6pN7eqZfYT9j4RnVCL62WRO+GKmEYP6kw9Lyplb0YMgiIacPasw
nUyEOuG1MtWeD1vzjyYvoP2Qxwh/IqT5Q4uHmblqIDC6aGY+1w9eAKqc2oAA1twD
bT/M1ryyDabS6J2Ftn0UQdioJW+vKlfLBchh6QND6E9RhUts3+hZx+yTIO5EVoMe
MoAOqzw4FBZI+Y3P/y7HSEq9VD2J95dRNa8hLSvimckvVYnHe2gSbi995OMF7vLA
+Hqkff0ma5a6ECox7ZMU/iTfhbXUoRx8yVipzdP//0KDepgpjNuld9MlRtbhUhP9
tK3YctwYLwrSBZKKGmpuooNXEkTcqF0xxTxoqATfQu4xqEVgsnG9xj5PGda9DX3C
C+IZojA0CSJbOcKZwfBQOba/iwlygjAB67dsGHjUPecAmX0TfnVGTrhU1/jGjEO/
bJYI3GBfQlMIDae4IhnLQ38oulIHdohd3bk10W2qJpPkXL00CNw8v+N7dIuxti3v
yWkLFJlmG03ZNAp3hzQ3H/fBQYLAE7t+TNZfonP/QInXLEpUjU9JvGx8sRopRQXW
KBSGJPqDj99IrFus7HwIOcIg1V/VuKMbXh8p1mrF9HEOeZUS1f9WfhV8yxXpw0DQ
955QNDXqtbOZqTPacNzoLISiAYeYyRvarTCtTZBH7DaaE1UfIimwc7j4pUMkbWfT
rfdzbgHfgzIvtO+OsRsqX1AdoX2C4m1P0zUB/fBmgk4fc6AQNjcJZt+fPJdiPA6W
74NHXLQqbqFKVCa8Ofx0FNfJU8W3fEVnL9XCCtyeas9LEUTawyiON/QmHZEebG68
IKNShyupNi0i/oOI/7eoPJTM89sTUUp+ZHlay7pDLbffCoNt2jVDbV6WvJgdMNBc
PCp2xQtRs/tP/HSSLkgkAsgkV9DklD5YaNGSDoiTLNPlzQFB4fetPrbQmwgX0hxb
bI9OJ8eTLbdUecspoisHoCiyFGfaKYprB2P3WqgpOJ1idReJmrdNlqTpiQ7XtY3V
6LwrqRVped3SnUTwggootB2n5RRO3Ov6pYpD58lUYRrX90WSqP+LaA27QSC+IDUO
FtL/R0VWkbQjAdjHP0xhrkVl8NXZ9N9wwJSXWHwRcPMrBiuW19ffF3dgggbny58k
gpsLcevtG7nKxlmsKUqcFDHLi5GS7qW8YhjXCMchUJjjzdEREBYzGKKx9LcYF6cA
c6Sb6hXrDnwZ183vUa0b5d+3AqWW1Ov6tCQTh2k6olhWhWh+7hNg6QuFLxa3uPjW
if7Ca5BPL3y+f6GAygi+JO3Sq6eqDq1qIAGaElRdLxmbHuHTG0brYcpBLna9NdPl
TY98zEv3HnEBRIytO9ZTppqHdAYYJ9n2buUAy4ZTOzHglVUFou9K3IoDpq2wnkVd
Tt3UE8cAtcT0BS0ko2Vrek+WfnAwiw62m3VBHpVS38awfv47oAI9CuPPda3fxoUB
KXqq3/dORYSf/lwcXJxZQViWbwQO3KQ+iGnoRbkNsnqDKOm6h+tg7bHQawxk0t9F
3dx1zf6CWcOI9JxttQBjinjENbJVEJyeQEG5MrmaR6OOel4F7bTLYST+q+KEH8Ai
EZwV/jEXq9w/+EKY1g6DJlphpkdoDGvAriDIzibSy7rXfO3HeLBovHjEqwguoHy9
osANJG6Te3uaSCZszOCF2GkEL5TuAkFuRn5P/4gqivxp7gQp3QmBo9jjFGmKO/LA
wKKKQMV/l9gwb6kZSuhp8U2SqOO/Q7DoEN/7OE45N8z5Qw2BHLscjOcIAP22OXt7
mlgCTlzEF10C8vTybztFCW6A3/ACRimwXWGvyfUr7v/jDnjIaoj+dqomv3dnfGwz
Qz/ws1TEsjrfbcsOGY9Oyh/EHc0PanAJzwje7ZgYpgqjvZdK2wamsC+c/expJqtJ
kfOJTvVvipx9cgQVKMg2wEFQxzpCbj3PtwaJpBrmwtBhbQ0Y5IlHVj0bG7V0iW+5
sBRRAHt9DBMjEnRh2EnG3uCbsilDag7X6m3P0L/CyY+d0othQZI39RBW87s4QTT4
L2RIsanUyrMXDO7IinKC3+In0SAkz50aBQWp2/2eHM+o7P7BBDuZpVMzq2vpG6SN
WCIeDww/W0sP3ilCnOqpRNIcgHWj6/U5pSFSsJg8f/KIBY1Qx4AlqylzDfGCZUB0
WCh+qm382T/gyACD1nFLZDoPbx2FtVaPzdDCRjotdQw1Gjzb4I0+rQJZvdYC571X
WqmGBfJzw+BWOQPBYtj7ubkKjkGZxoPHRggrYMX5s/uPr4XIubsDWu5VxxqTVqDs
DFpS7a7w/0tfgiKFNb7xlr2t0NqkOTSPg+t0yC0vw9mi0IrrAzh+SQXLkZwZsGd0
OlX8U94x05afPq03kZxyT76m/Rxs7Rgqm9rsAi+c7Kzj6vCt7J2Ms3FXzPZcck1A
kMC2MZjdwQY72SDZrzn/NAjWal8kqCsToghhk7LfIOXr+ykDDtE55mGTpJwEKBx+
5vQpAgyU6qqr+O29mRJS3f8j9fsfncS8vOE+GQKE6BJZUj5ljolbkQIDkpUIS28I
pN9IoLwoefuijPp2C57eeKpVmpMoIL8YLwI5IE90sMck4fA7z5/NMRvX33N6sSPS
1bMR3K7t6N5LK7igaVbAN198znVzibRKHVCTqs5y0XuYPwAGB7H39L8Cn7wsjFTk
OzIgNhtAnByxvHTc2ggD9nj6UgBuq1EdqHnOsapvZGyN25GNv2aQy8SBSpEfn8XQ
Q14DRDesHkrWIq5xO9ePv9KZGi8rWWvAZuspPUugiUGWZP12emSQ1u6RBtgbpIVW
lz4EFiSSakSl0TsOaEDalBrm2UHHSJcqYv8LMvXfshoIArm/2bsFK4mm7OGjxW6D
aRlUSBEr0Xww8HgkDt0Y3914eI+5eC1SgeoeiNlqIuBsnI8Pe4ZaIfNkAji/zyuH
tCyX/ptRk9wBCt7vUfM34oOY4XpUGuMYU2p7QghFq0dG/vjVjqXPAFus2XbevPVs
J5XTl//ZbC/dg2Geg1ErBCGHf6LPxEm0N7b/xJR5gutuceZYVgnBqz99A4mJJ13x
4UbhWvIy049JspoFV35vP392G46TQTU+UEnB7JYUUPlRBYI9VD5n+9tD06XRH9wA
Q/tzEMtaKM9ZLFVsly2LmZq4j1YY3Rf/gseB294OP5zaEsuJQUHvD/0AGwarmsWo
zJdXjzJCXmkusLDkCVPvNZ2YDD1GS7/3T2T9SJNFRr12WzVIy5gRoRjmaktGXv+6
rYAHt9CenxxBvPPdiqUiDqj8wfJXHrHWSYX5vOTDkCteLWfCPl2Nq8l33yOEFVD+
iTVfgHxS0CEdx380GHqofchnLzGrIK1uehr33QmDbwgCuDjoG9tf2AQyrFbCnbW8
jAN4eo2T7cYZOi6tnyZgnROW3pmx5VA4jcWWFl0UHYMDsgGDT9MLTw3gz1aLji6Q
nU8cpR3KSHFYgJBahl0VUo48gyExNZHMAlaEP5/c+q4ydvxd3PvhCIOsD1l/7Dq3
KogvfXM+dYY8eq+MzqVceSOkQU6WP5Msnu3kOgkVL8AcR7LCt2PUYl2yAVYQ1PNF
JAty0Dn1VB0pvOxVDsfAlu8cNFraih0HyIL5qU/VlxYZ6t9PC/hyVTBKP80Yjdti
pF8G7xGCxYs57BnYwMPlZar+2p7X5uXCxrxsNshQeqOHAuaXJYabchCHzr3Blodk
/f6bu1C+ah02lOJPFvo+VtimQJpVUiHau91ii85DT9XWOP4TxypP9lCPSc1vBvZ0
hX+t0J1taz8Q0kq1AIbbA558QqE7eVl6aBeTguV+d631GcUAFBlbYL2c5uHT73yI
XWPFzAbIuFM9w1jAArwenWqy0TqGKUO2yvOElX1KP2fD9c3ZpQP75PN+j56KKO7F
kH/CjCkW+fii/rYiAjlMyV/1tZE1Zc7YAEL9lBffni7dtBP+M3IepgarJP/hLETI
vWedwy1PH6ZXI1oTHojDg911EEDO25PK0Zbdc9A4pRsJyjnxrJeWqJYk1Rj+fiGs
SV0z+ebDpdeBTJrvu9yRUpb7k6L/eiJ4hyTUNhq/YyqkSTyi2Rzrg8vokcAs1VP2
OSgRgfTlmfQL0ckJT+uhURhes3tfSDxAn7496232Mxsx2U61bKVNEgrvgaa9I0or
FEfcU0Hb8LFksOi8wzfZWWqM7yXO+iVwQeho87KQhXatmSkOUvTX+zAVTbGYZRJw
QWVVkvN0bO/R4fLwhP6p6TQ79VbN7ybcOuXK+v1zfZ8CiQok6MSn/l1CZ9Quc29S
ep2PgD8Wh0/BRP99kPVGJt9F4/jYJkte8fK8BP3eppdiuv1XdwqKLYmyFC7pUzIJ
eP9HRmHE/qkyAE2vSiyCdvVx8T46w1WilYNrtluoulbu4WpqLdwBa95343AP+/UI
EnP9kOFP2zl7z1p4mSQUGcy5PkeF0qmDQNCiHVDlVmOSx0ueXsSEz8I+gGqf+71t
M8DUfsz4OUmJxf1W7/Tl3QH7Q3XDFuHgKY4JRVgkSgJhzqiNDV9d0dTJiglqzKxN
DOm5ZuhZeF3It1bVMXW9N4DS0lM7bUBJokAx9XmmO79MxWvxmv5kNlyHRIPaNhQg
3oKIsY9aZvdyxPBgn+HNGqTQwEnRJ9zU+Wp+xWHW4GG6b0VrMQoBY/kjtjnGz+M+
UFJyrFjrIbTo6fVOac+tjKSehzuolKcAym0VmHyhWHqwi1kTZ3V93wOL2Xx09JLJ
xQ8CWDHZ73AETeWJlEtn5Azs6SEZvxYBXy6k1PtpLTNt4CuXkAjDZspvtXEhLWo3
86J60vhNhM2ud6KnsWP4roeHftBlrV5QR3fCRNYw9mNiK11k3eqX/GwvhRMFhbsz
PBHPAoO+frVlKfm96FWvMmDmJ2TcUmS2hqYPNIYoA5Rwm5EQHQA0xJ7MI7N8HzUq
OcARgq4BUQ/BpIlBRw5AmnIQHAcG8dfXFQzNSj925f+q7R1f2PSnKG5meCWE1a7J
XYxpC8of/BORaxE11Xk4g+TFddNTmnhriMsbybk0fjWcX9smjF62IXGMxBlfItZm
OWH0OSyzWy2aLjo92ilpM0KNxgIRx1Orgoyg92uD5Hh/MO69P38TgeLeolccnN30
y+zg9Y8eg8BdQiGH3Ss5ml4QlIKGloR+XnZZDJWgh6BYVr6Z+TxcikM53nGL+k0R
D+aYgv1GdpD9Pi0MbZZJ6uHCXXAaKgWxZ4wntEEKPqz+JPDDP4VOny+8PMXA11AQ
xNnrrZ1IvTGBrk5FTtN9353ynWHb+hOl+2j4IGo63uJXAZILH7fxEpvKAiA0tjyI
bZ/GiOkmtDD9rZ66/En8j8P8KFkvmBnK6B7/LIp6f6wuAi004NuyuvWOILgYEgfx
D5zOF9Oa+OCFmjAzPQdYPKI4rq1e3tZX8ce29UUmJfkNhnLdNdG5Fkrds6/zt6Gg
ypOALQFECsJ+2vZleY1IDIxOMU3smBQCK7tHMZrudVEcHTga/DG9jF66tPkYQEQF
k6iWLwZoGOUSt6YBqNuesWnp/YzEq/YlWThGTKN7FibDKjzSEGi7GEte0T9Y/ini
C8+u9I/7wSWw/U3HQHJ3XfVUhs1zHEWMbHIpG4gYC3+Rfu8HTrbx1KxbfzEhPTJM
aQltb21iNK/fjLWfwSVSj1JqLx2eEF+mT6rN1qRaFVKZO/p7zfrNzhOWP078r91k
dYO/1MrBSoolplI4OEXJLlwtwLqPo/C3Kpha0FqpzQce9Nomw8aSW2s/jmOWHH1I
xj93YBBoG8s52EzeiKXbjQdvfPUddGdGbiA3Nr7LlYkNbTlW4sepJryzjJeF5ej8
mB56U9CV9e1mMt7FIfCjzg/oFE5SF3g170zh26QCJbwCAZeMhkAKPYy7fs1WLSdp
w1j4FKQ/5ZBK5orm3LrpNRDZzsDo4dWCF+jwvphDPP2h1KMayY3YfWpZBKaMLa7e
H51/7vX0Ntu6wi5XZJPIClSvzN2CjpdRTuefJyywxloubaoNkCGXY24P7P237OcK
/JVREB/5bbU1n58QJRZKMbvYeT4bykaAfCZTpS07fJsdLaG5nfUvT0kLaLD5Iuu0
+AnsOxj3a9IfFLhh/GsQuZLPakYlXS20RLZvNlSq1NOmSjjrn1+Vd/BMEAm6l5kq
7VOWFxQITR1gkjHhUd7MpklKkbA/oF/WFnx5QG46I3uPyA2nXVNOMFhVBoS/JO3p
MCu106msxXSn1N2771Q1XzkQSN8KBSx3YWaaydSREacp4mYfMdQ5BA9S2rjM0m6l
4BsMdtKagZKIm9p9PcfoaWH5arlShYiQ+/zzIeRowUgzA4V88+YGyoe1/DHJ27Gl
tu0xi6TaeiZAi5ZW7EY0WUa4uzLBVzPZOqOVehdsk8ii2uWE0smMhjVA+ul3RGKU
fXiZM9YmCE+ItiUUZiwiGSqIKcNhi0nUDNV8oI5gbvVzRNngOojy7cCObZgSOiQW
w+Sb/0yy9JxnIAbl33vmNWRv53vaVocF/ZORkPY/Wllx14dbFGKnr1sMGZeyrTlm
i2E2CBlFNrGSAU8V+uZr0CFhTHcuYOFxj1OzvBznuIYge3WxlNHjBIk1sC7lvIpc
YzpBkBsg6zmzdIJfQkKzD7KYQDpvReUOoGbeiKiKrV+xpDqJLMxXSvfNYgQu4Jda
/N4L8hOTn09v7NlYNgCbQsgPNNnd9IJtDfSte7l9IbDuKQXKMg9Q85+VUJb+4nkx
9kwjJv+ewxmzIzFPXxUTw/8Sei/DjsqBkZvp/zxtH8hqtfCLrjFT0xAUZ5PCj/up
TlGag9PNOVeIDbKBL46pGi8XDzvA1UdzVb3zSHDC4PuQbzP9rNuPiQTTTbawDd3O
sYsvBuMoCVKcE5W6Vbs7PZNC0W0sjr51jh87TNvl/IZSbxGy77NiILdSDH1LsY22
TlBQnVnq8nQrM2TLoG94eV7YjpFQ+Yq0iZmtaq85GvKfcc1mqBDzGFNvtWv8hV8w
8+vDG15GucXnNbH6gRBfb4jrOaHqZB4ZeCNPvGO2cGsqeFb/h0clIQrA85V8P5i5
15ctNuDbIhVUmtootwYZs5pfVypADPYqL8cU4TRJ1Y9HRi6Mx8oQ5S9K1NXZuNLm
A+bRHE79KuyKUgVgiw9QKabjK7LaWvPJIMuU/bNW7N68xd39CYVNTo9lkMF9SKp+
CJ4nssn2gPoD/56pLemhxh+JYTHokdK2BtF7UGYVwtBw63CdKzd2T02xFq64RNvA
BCo5RPPlj2+tt4XeGJxUG/iQWS58MHk4JT2L0O3vS2bKaIJeXlyBVTDj8b60P9CJ
YhDQbLfkDsYsP9d4w66xot5D5rdMFZTEW9eQ/dn5UEYgvxbX2A12VsoJdu+1zOUB
b/vrwwi3STroqQFxR3yOL4T26bXDrr/XQWCpvpWasgQGRxecQTozUEgw1B3ZWB5b
i8BZCwZF4bjHy3LvdjgjkMAIhGE88ek0GTnJiYQo1CTJBjWdLydNGPRNBczY9aud
HZ8oa6OjSu8cx/Di0YzYkLFA0JOxWxCZaIf4w4t7rXT024FFaAtBJ0L+oCp5HM/D
y4zXdK13riv5QztTnGw5sOt2RAHaSOibwXxpm3Q7AvtqxHxLTo8gjUFZ06QNZ9Dp
HgNmPFqSh/IBDgQCwZQZfR5vjUHY8UZNux3nLJRrzIilMhVGnCmvLezwfBS+rNDD
tN7x9GcQ/5s9+uNNZPZrFqEzSSCkcwa0re0yeCq9GgxlLugip3e3R8AzIlwqWOg9
SgNKNIJgHkEEjbAIEO0RzRYmsXx/PkJ9TyMfUAte+ygqXk4kKwajaXRDerl8B/iV
XTyQfe+LulxtCIneBvKxUoQg+/m76fQLLgK2+h4Mw/YaOAPToZZR8uQu0VcIPCeK
vwotnBOjxEJ3exmkVUE+OoUbLhMewBccu2X/Y51w5SXHiK8T8x2haFdJwG29+9TJ
4lZc6aJ540BkDrpO2TypZEZrQh/IvJ6iEa7es4i+2FIBFKC4nO8MxOaVXMvFww7W
eEwRs+qOKyYJ0cQOmRceIx11stznShDY1njdm/Afe74qvCe2b/rWtcX5Q4u0W/G4
d69/Jj2WzHytubgQ+tzOyJ7m8gHJ06JDy1/Emu//hB4PY9/OMEg+YJ2INUTztJrw
U8zn7RuQ0iMVMdyueHki7OKBLsF/BpDllgC/ZTHq+O2CGgr/IfjDlpWTeDntIjM9
KxhaYfPFR3/eVCe8IbQjrmpNZUNlwrmMGOZcRrzW278uTAOn8zPSsIm0wObY6+Zy
CeZSLavKb6ldYk5uXui/celOdFp8npkAxLyzxYQUsbUdQWNWRkQieNkRI3amG1d5
wXwUJ9y+EurrTX4iw6d8hWdadXKo64nWLcbnq3pksqW7OQlAFUXbRyPVBkFMMwTK
vE+l8YqlVu6jot5BOR5X0NQgBWKE0XfoeXmw0YyaHTaBzoxB65hId7wjztAmiHAX
k/SBZj3ByZ4KZUCGDhWW7ecScnJ5mOl5YD1fGRnc8imxHhsVn9ry+X1RghyfMh7S
osFQbg4ztxmYL1uda0po5hgLOP1vB0tNArZtzRFEB7i7RVz1xtlcEzDr1pkVTh1w
Ia/6ScJDdh1qqMGQ4tvkXnnPy6uVEKWhz9bXlHze3mzhH1dqKCGXO5Mo2ujzF2ZG
0yHGVJ5xnFb11OZZNfSMWHQ3c7Btpewb+ojcMBGO7S19vnAVer6NCqVf4Bt/f8eC
Qrcol9l4TOVUonx34ZnK2cSRYGqd7P4x+SbjIDIYqRfHhQ+rq2z+dSGC23EJTzQW
YFz+L95koZb3dl89RF6gh8zwI5c5y1tzPP5/FKCfNAzoP4Ql/yOnbdpB3eGJeNjQ
pqzN8dQAvaf9LbxoD0LXD/sMQXztVHVynHZXyaElU2iK3SvXd0kSOzn+qryvepTZ
ONpc5/hvQ9zZTdQhFQGKVC79xhh4eqP5NHrF85g/E+wdgrmZviQ0R/67zmzNRSpg
PQbQot6vPrw7imyugmv6A2xpGthuhFVoujqsGfHBDKxRYxgZrETPQHbhs4dRnyUf
vT7AvkNIlyJKua1d48iwkEKQDZXRUOv5w7onQc/A4MLCxPxEUGwOPuTM7EUYyN5H
mIK2Fr82/Dh3+3laErTspbXz0HykJwhpBmkp2cd8ajsQNiB4ZhG7QKVVOzsC5aSQ
ioUyGy3vvXiB3AcgM4yp1PEdouvUaihMOS3kcMLye6b8O1Eb2EpiaIkHmOccLbC/
IXAeaEsB2mTTs4ADLBU37LYPM7EE0TusmLIcaxxqDyQ0kfeYbxqEZWfzp7DW/Hw9
KuNurY10mR6Jx7qc+oDqOun+LNngnx2V8SHy83IfZN16k8RpXO7tiBUi56f7JTk+
C7QKG0YZwcn1gokWpEDYprVZ+P+i6ScRRW/wO18aNKE+jr5AE9iaGCJGlpLT/v7Q
qsswDVaU3rKQAWPX2NLh0B+71b03ii+bHtgBL7z2fK93FDEuiWgSpVO4AETBRdLc
rM3gNSzp+RIhBN2uLeO13I7So9uHf/cGRvwbpTTAI/7hox+M1PdUErtxvLAxLAzf
yGOhaQayfKrHi2OT+RynQuoz8CCLxUhbHxyKrPcn8dsGIx5UeScj1l0FapI0pUqJ
QKUUO0NqEF8X3EWsVR9HytuqO3ke70eSLBKGuKPB3bfnMhh4+dtPwa4faB0BG8sb
1w6E5yPZsY8Q6vBBRjguYglrMMJp1Oz12QcaNySuibHf1/ba4C/RbRj9m4enGY5q
zNXKs4nC1Gn0CtdUirvXFVjshmdpxnl+d4Kyip8y8H6z7Vy7p/MtoAaBOY9OX/XA
n/SjiF8avt1tjfHjuR95E+MIy+i8XbI9JpLmakx3K+wMGlEe48AWtxRR0hRPKt2o
hp9UuKsyAqsDITNipm1K10KZihY9A8HR2AQtzh0MEs8IX/kLBQmuPw9rIZ3gCU9r
I0bXGYo5LPZmtU22XNIP4u/kv6UFz/Z/ktt8iH/lynW1ua6UihDEds8/RojliNVC
kqUjY42oyUaJ03lEyPv066OcQd1AOTCQ+NDm9WvjvKBvMS2QYhRy4expdkltakVq
Ni2pLXTu8wIXiD137gdg70A69bozwfNd693v8S6JVfFtNKPU5zkAqtJx5xaYLtF8
FfZGZPdwUz3mxPPI2Hc+Y1pMpHid0djZqUoL3JK6ZWFYjNZrYuIrd2NAX+0GjbIN
1SE3zyTjCKHPDX2RvvlO3yGSoL6ekJu/Q7Ye3sEDryANBL6h84J0HU35yYh3F6rR
WXwCB44ebi7tU9Xaa0JToSOvKAdtgs+UlIWPX5O+SFHuJOIVBw+t5fuTsADW9hTH
Ja9C+TTDnOZANm4Lcuon6wfTvrkv/2gK2a4qvuyOs4JiJW/u50qP0HrJJwxm9/92
ReVQPc5g2gJkjdJlbbiAllf7t0wIRkercL2RpmUNKiMeWprBGCM7xRBw9fxJzg5l
uyRjtd49L7b8OQMOUcPg2b++77lk9f0rkEGsL3ycV18/o3XMNAt/AvaTAoP40qkz
tcS56Wl5FDYrv+M3eGjalCckJBrqbS+1lRC+rwO2c0NI7WmoxLmPVgGx38Dniddt
yTA77aRAcgTpGsigOq/FSo39UXCmKGTk4+3V7GTuYxvwE1Ix+wHgR93KS51FD8xO
8yJejba2trseaQj9/5BzYBn/Anug7weTLOgKDhPHMxYHidkZCMuajDDNQ6M+i5Jz
PzJ//B3PgnRvV8lwHoLRji0hwFUopszmslszE/UxkU7nSnYv+UmKePzpN7zNRVJr
+H8KCwbzgx6tb/SEKz8hb0PYzmCT46ZHcAx/ovCaOxLf66wUfG1elwcec9WGRMeg
TOnDVHzJETMtvwRghf2q5wiCU252sRSO31JCyFyhlZpUyPZcOTv6H3I3EmFGc2kQ
2fgKXq7u5DZq49Sbhar1yhzWtJvYDPqP755Pupny3+1xQ83vlilHyKsDZqQGXZez
YNUOecEF3DDCP4qfU6fy0+8Vrkj0OuZVtw/I7mVj82H5La8cnoNl0MDAmmqio6ov
UlrQHp/5WYIciIsX59KN2OzjPlyr6OV+bG215zK73imrfIJqOsVDm7KaPisD98ER
kg+SGw/qt6I6bhjBtW8Jda/iI9qHIG6de23s4t0En1iNGG9+pp9WGqQL2T3dwnlZ
tbGfZcMSRnScIhNIrdrcWNoJrNdH6F7x6ffrKzjvfcYwEZZGwGHhc1NAtYAdcFZu
+gB7mCS2pWrnkNDD3uQRroeL9n+XVlPCjE3EUkgMWcbVwkhktjc9nnWy0lIs0KR8
nfJWKIQv3jstOC8O/a4XgllSlKNGGZpuNgmeh77d6PHFVBxRfbj7RZO3NMTHIOCI
goK5+/eQnkTpmeUcsTMgnNXJ8TfzxT6buwD7ZIZ8zTNls1XiUOJUdhYk8PhLIIEG
eJpePzc24SnZT3UpAHVs5hcTSRclT0dvmWTNNNPW4Be8Qthvolpg31BHc4RMaki6
POs9UozBO/m1H+NW8jJhMj7m9a/v7zZ9BQU5fbzedGZ938yk1XP02Y97w2S+lz6D
RGWBJGE5/AIOFRB6BI6GqKh1bnt88IxZVY8Ya4hXxOCbRi/a/see9kjfmEvizTzn
Sv8VFONOmvyaYwOjskkk4d0JJuCKDdyYgIlPuxZjETPy3wIUbN3CE/91CSW5J+5C
gaoAX1ka5GLyZbXiD9rsCNdvSKSvTVxZ36RkOb2lhO6N5vNl+daBxavPjwhbiV42
XAoTE8TFe556A8ydB4AtKEk47tMlLD0aFp/9IQduM/Qsfb1opJaBQwCFHSy2GZTE
5WbyCKKnVcBxEmB1MOe6me3eZYl2TMt+OJV6ClU8uwWxURgqPzfIEmv5U+Qlwo6J
V+qnX3PV/eOUvkWDw6GHDDdkOZsweYeMB3bR3xiPnpMMh/yA81hBIZf+LSfSYYDA
Pv7KAGhuMHO7tBfm2d+1rOW0LTh0drE6+uikc3OZ/r0lIl3qnMdzWHRMaoU6lNHz
X9CEUbtWNLinliqllt/KpKUQUT+xWrfA30PELFotrz3I+Yw11HTpV3xCSCXLqv42
Ieb/SsxBUJNkTR5hmyE0xJ5nrNTDOyjTOjetdBJgg/ABCj+WWzT9+aBYEXYgCp6l
ldkcItO4feyoS9xUfec0WrSNUvuQV1QU63CLMJw1sSevEJjWqcwNqCIHgVdGb9ho
gp1KfGGPwZ/6fTpI+o9TZ5fa0iWd1jrphGXh9BqG5irvVZcpwiok/n+btnEsfaR7
oywWOnw+8tsKbPAnhirqbi9Z7asxyeiNoqBESd3/xPzKK8tOZdgbNKZqlPGjDXVI
+wOcUH6sbR61WrVbEf8Ky3ocDlfX8h1xIjL5lKfxpROUEft2vec9JEUZ3mEU4bIT
qWLsU0pQTTYRXnPacpxmjN+LSTO734ecWzKLICwm3ioi12mGnjW4VcNvrdgOLafD
2R8BuF+XB9Mj6yDeKKsKwP7hV5cY5pEHSdqlN9DbAFMvqHGP/42lR1lTwHxXbHJm
EPcvTz52F04TJDnE5P5B9tNOW93BuQl4A2GVPPgItonL5QoKTUpkoxHegHz7OKmE
5aj5mLY3+K0YtXoTHEfSZLF3EnWta4yZkVqYrUVCXtbqWiNTYUil9M50dSCbRnjJ
aS1wzkrM5/c/JmbOmKAHK+T0eBECGk4dvEeXB838msCU1MqQfLy2Fq3DES8BfXqH
p3JD8IjiMBdwvOG5b3A3dNv56ilA3+rzpKH5z/E4jpPAfK8Wrxn3AVvkf9fjh5N2
xSAUr3MiVkLzc1Z7d171No+/XY/QPPGYn6S/ayD7EJWMaKhFUU1vReZDkwAf1XJQ
4Dbdv9l4gLwKgagwFK1K1ewbopCiaD34ooMTjgHKFg4V/22JL1I4Ymtq3Bp5Bbm2
kHnVdarD6B89czSWm75G511SanSVgRpRxdjb7+Spwm93YdtZnWRxj1/n+x0CGyzV
0n2laxIaFpOe5pFewH9dOrN8eZOKtx2ueIwaZKiystWlahZrKi0nmKhEmtZBr4DC
h0G3iSok6JR4GbMfD0NoM7/H6tNPOImvS+SvrA55DdVOCDnJqA4vufyo+qnDC9bm
eROBGOvMcRzS/UNWU60pEVkF7zo0i4aOX1Ofw7l2nyYIKlC706V1cyfvVeN0ajIK
zKA751OipHb2xEGeCSEoAadd+uKOEjGVbhDxTgndT2yXlJrHYHTi4jk1WszwzDjW
SD3H+KZqe/D2JS9JoXF6YQDb29z1Yr9/RXarbcPa7utAJHPXKqGS07P21X9HEcw2
D3XNfB4dXoTx+kmGxDWXom3EmiUBGLekdEBxq0mgP1FlswNmLMM4n+c6Qt/8IL28
1LZLwPnCEJ+/oVdUMKGyyNL/pqk00DiHiirkTuIcyQRkFtaNv6MpQgLD8l9nnuWL
GORWNIJAFrwXq5lkqtDRiPYYBsftxB4EPfbbXeCZX6d6OE3E+HNULragZVJu0UM+
Aqh25HVEVDNr3iCXp5iNydrcsbdygVO96Ym5bjUKgp8OfDmCDoKC8nPrri4aKjvM
zaD40tm8nqXvnFP4uxT5OAIlPggaIh5XXkbA88HxULansTzO+iMLwmjsVz1w3/F6
aNPkIU3IxkTBl5ldMLnO6pZyhMP0a17Grljmap7alCNmfkxXouTQtoJOYOXRFS0f
YP7jqCnVpCjuqqGEC5qiOxAHy3rWFi0f33N4o0Dw2JUQeUL29Ne9ceuBPQSRgX1v
vOCB6+NGoMUVKd5dQNyifcWHS8dS7bbgxdCw/43d/2Tgje6tHJDL3EToz1ES+eqd
uWuG7KrJ/FcwOWidmQzdL+NoFwf2FhaW3197BHxIRY34fnoaewHQsezp0ozMzhg2
hfD2OtsQLzdNa3N4ZXh9Ecs2Ii8+kG+g5ocfr4qbiqlyR9iiSVe9oqyVdl/leYes
8c61ja1ja54OjlxI3iwE/YWmm5Hwt9UUo+iwEekM9l0PHigylS8mEUL24lI+o5zV
7P6ubLH2BerfpB5ZOoha83GK64hzVXn+NlAv2T0Aa4+zCPPvaXbYhkUiWL9KStBg
eqgDfY622mANmE8z114ELMIvIMr28VqbenXIJMd2mZnoEd+JBNQ/l60sxxdKYv+V
TOah3FbbFyzJec9hogZM/YR5Wae/nJ37AJ2ApgndAGxmW37694qV8s+jCGMloiPz
Zx6rjokj0JNcP/a0MgtskIMlBFMMIIFwZrwwaBji56ZbVUw4uf5BfVdOBuCKHjqf
A/OKhClYL4PKffIGILXp+K6eMpCmZpJ9drJaun9XT/DKdIwiNKvSR7JlBPyHNQry
EErRr/b6ySHZ/VvDzkplV6MoAcG8/+MAlZZWSJg06j5qW5ItCenC9WI8epCWJbbQ
Jj01fK9ZvsUDIeJCFcp/mTBjLAPJhZo3URou/Jl82Yd1DZucXEMcW/v4FZ4XSaDA
lt1iTX6lQ9fud2fgczJCnW2jj/nHY7AQ9cCxavnDf+Vt2DdAJfp5iXG8a8BVSioO
SXsRR7CLBq7SBhUKe9fFkfYwYhO7f4kR3Le4q5mupfGioV/8pdM10IVmAUUqsYhM
1Vucig6tnL6TwDxXF7P5G8qx4Epo63sGLsSndOySD9uIn+FlkBHVLJZGFcAsjErD
sEjr+zKtacYJ6rupIGwTR/S8OL9W+PfFV7RY4ulF7SxYZgvlrMy3v+7vyW9FAb4g
HMVE3gfXpCkEjxql1FWMUH1AopqiJZxN183vYsZvNwrlS2mXAsNzI3MDDoMrq6PR
XixiPXdhOA///HRn9GhFrLEGG3KwKJ/DCzKUXseUIlbUATDCo+iPYPgjmZ/NdTpO
ixiCqIIWR1wTvQH98F11llv6K62z115MSrsgkYMs+qFmghZwVnI7GW801VmTW727
OUvxZOAKd8uemX6gH9Xr6zr4pGHmuJ2fQDJTB01JaZ3KY3kLDvky8jsXZDeA7d8s
gmGh4BzhMB2DBKhmafvYKqTePOs9Wt31O+abTGEw+PfYYhJC0hGCGKR9EZUCV0Tj
m/anOQDLMhH838W4vqxyFVcd8b7V2bRgyVFoX4RARoRo3GY8etzXoyrbUQJ6FPuC
4ssuDyKzhkBgBK7Lu/2NCC13hH7/UJ/axuVC13En+WPHgnEz16zCTIunSJeCB+ae
3kZ77P+gLZ2W8vVCu1fFo6lrBwhuq5oHw+ugx7S9KGiFOOiocnWjudITEEFVHxo3
pN/n2RhgmAHBtSzPjq30C6v1bgq15DaMeGZXlPbrl3s/2q8WohDcXUs7lwIjdTvh
F55KTS15ePb/uKOQTd0QNgoVBSqex2ViQevq3TbPNecS1s11+kGsMvER5ZwTcR+o
S+5RG9PICG0lVTcd5OqzYofjF1a//BWY5LLRZJNHVfWkqace7YMj6tGstUsGXxyj
bz5jXRLnxsMBdX8g4NsGas4EDSVOUnf9sJHQkZfzVX6KSTUNAUtv8vLdJTaixeg5
ewb1goroviUsX8SNLZcydyfvKI9NywTYibQr9ESViGt8UK47gpWDU8lQStfTc+wc
tPHsLwji+TsJNlj6aj8gN5RIqlsGYT8QzjOmVAR56929+z1g0iqUddN3riDspwQl
0TWJSSmE4Kz3o/3Fj81q6f1CDY2D8294zPVX88x/6hzeT6QZKB6oY+3e8rYF6v+U
9kaFbFFcVZb1DQdalw9uwMiDvLBOvm1tTO4IHGFt/SqaO1KI2oHMOY97In6vGtiB
vVAVi9KnmrGp7I0iYZX4lp+gXhsBqg5mesS/Yjzr/eYglq3scHEGrHNKTTeZ928J
ivLJUFAuXOq2QiPILXUc/3d+dT7FHg4hrd2HMEIH61GHwzXqW7p90QkH8FMhdyVz
5MFNfDPlsqbebP2JP2M4DiUfwpSms2v8j/Tg8tWu0WBXenRWDmJ66ID9WAY8+6E9
jiyG4guK0qkY8sXPiRmeJkndhhAVMbOahk7OogRYLLbGsC4IoCHCRxpllVeJywr9
2LtooExmCvCysonCk9qIAx1vDPfTFdQgVGspy+NWqz4qwAcyKSp+a6jy8Kp1cdG/
xf73nQpjKeqXvrLvIIKaWIOdIRDBGypqkB2c+md8vE8dNPVlAQ4UILk4zosp9CYa
V1C5dSCOYRcnfojbO5e3gaZg6bvhm0g8E1cr1dX4vHxvz/c4iWot5n4uvm/uY0c/
mD0/Puji1dhAemthxNprDemcLExfI5oeSSDgDMlUsE/Y61MfDOvX7f9g72ksdkQ4
XBIqCrURVQ0NmBWyqWfPrQjfbGA3Ji5SRkqlJdA3XRqvJpVWPlIFVCd1lsU2buts
4WMVN0QFTfuR7VkDOaccW0gUHedG0BM+gLW3jMt0FwRVJWlvugCyJ9LBYRUMKnWr
s1+aU97NTjSleg+mUHbrLxnAoEHShOzcwhuLMo3YGL7DtJ/wCvpf4hRGbzeREiBq
J6E/GlHFB+GOfGNZO2AFccpyERj1/UySgoMqFFq1Sg+xYuTqWzztQqCX1XGggL14
vHffa4yTL0AiHrADHPyT+7PqB51jHs/fd0H0ch+Hkx3hxcjp2a+m7/E9IN7XRq4V
85X3oPD6saUmzBm4tRFsv6N+EGCDNVWPFl2iiB0FTzTL4JhNHFh/WY6lm8tNUYK4
L2QXL1aVpV4hfzTw4G4LK0aQTzaUhAQ5U9jf/l7GCCyhvAxnUq2RBCBRur5+8Iti
uuaO468b8yeJKSyofOEdeN1cXKIpoMaloQc+SGGLAtOqdVHvQRg9sjKZ2tUIhEB6
lcPYei42LcfhLCw+AWohId6/WsgbsHc1C9RgcvvOhNHQpGzcOBzHb2/O21D9K9Sj
Lru0WfkZPCoYZ4lP/PhazEXLrNwtvOhwp1opbQ/zY6KSNJrr29Zjb3sf45GMiabv
XUGTHc5LJnp79+RjLaGd9E21ClvKYVuX8DiSd2npWxJfH1hoZJJe+YRwIp1dSy3v
1dgz+yq2tdD1WCfmD2DSV2bxIDdNvWLNG9cvn36lIYul70xatlpnBiZgbcvXQEzJ
5OXa/DSB67bbVC8yNgQy3a14x15/DSYwbJg9zVHG8Is1dt+vdxMfMia2TGb88e7V
fkzVR1UEZ66i/y/vFqGVbaU3ldzftr0aaRF4uKG7B8NJXwg2QF4ANbD+WJ50h0ww
sUXAAPmK/QhaSCQ8bpGBE28WAPb0wtMvDDNQBuOcw1qS8ApAEb8an1iC6o/uWn54
sjyCKFHzJc9BnTTQT2nD3gobsYBQGU4A90hHB9fzFR5jA7noKzI2UB8noLwtthoo
nLllf6XrMpgIXUTCMrRlEJGTcGG3awHvIMgAyg1z7HUtpCpEawo2B4xPSxAO5gX0
YLEnwJakWZoP/pGb1WxNq5bMdYxTl/UIAWfdLRMP7mH1Sz77UKs/T+Zp5nAJVhLB
Q0emWHHfu9zzWB9v3nd7yLLI+WgXWGbsRsf6NDtqivckHxONa5XeG7zwC3lVUrBS
NmVkBoqYb185Y6UhwAPB3S+AxzylUSBn4lidHyIffmqbBEha8Nh9xlm1hwVDEvbq
DwkPJ14rNvRFlvh2NuR/QeOwr5PsjD5vTDMRaPi60kJj1TxJU6hAfWSCZz/WXqk5
veM6tBYZbnbF4xs+gKsvUmDy9kADlA+eW1xHLfYVATrAwngOYu/nAuiKVCRxy5X8
r3UFBvnyeakwVV6l5jnH0kqeicAvA64NdQK4zQ7sXNDoQnJXDuqRbJvGRj+ZHtee
NYfkS2R4mWyz/76M/ZeqTV6V5xaEHkp2Xae4tpN+rcowLhn6+0+//BCY0VHMdQRU
JH1Rauq7rpNmZCXrKVCVHmAVp1bdZohdkKGc9Bg3hEfOZfkuaUS+W26V6Jq0gxYR
rxF4yGfyYwhUDasBl/SaMSh2UBe2qSIByYuUn6l/EuZJVMqTKNpVwaaJ3xwP86RP
iyWKlXOWmsM8cb2jO8TixYDmRN4F1hE319+TepZxt+8lNTz4+xiTNmHvSfQid4pH
0rm4u/4pxjjuLetxZr1yPHxfTDZN785611p+GiO3fiFhGJ9pweAu01wfu166uTX0
oGiLOemP5cVIg45GaUevoeLNSdOP3bn8BoDMH6b4mXQYhNph690gzHVNpFJwL0SS
h53VolbT5uZyCawUhXkBZEcS6I/f5It1nNtr5m1qW58gtatFaC2vyVp74PCy+Hgi
GkqtkF/mepqrbwNr885j7gOXMhgAaT15cDv0fTi/oZFj6nP6j3EfKcfHV/EY5eip
RHopiJem2o6MubfeShzyt0+SyfiXV2faViTtu1SbimJQ34H9oUEocrUiN1qOlz6b
kAPrynvw1o+VOAxVcP477Vq27l2vR/6zKXewo4XkRX8K5Cz7yHLD9wpZYShfQfHo
GQfDxEAh9jKopgW6DCmJwuN1PrcGD+OPDCwGfAcRhuUowNjo35a+a0WzyQvlOrtr
T5PqYBoNjnvWfphvjGqH2qWRYZqARt1Mt2sF6n/4GEJGN7RysXf0ryV9XbzMAuu7
9GS2Nb/SJ6+XRrHV5btaKfu3kDnCV++x+0i+NJjVKCn1eHv+rsay6Mo/ZyrneTOp
FsM564ygd3uNjjt7spvGUJwjV1U0ZSx0FD1eQl4DgWvCEchP8K6gcsGQbwoSYVZm
f3LoSbxDdNIFCAiGrcGee5kwDcobBOIwxpMtyYX/OuqFdJEYLshQc4L33wKN3zMb
FynlBLaiKhT2rfDCzg/Z9OzbxTMK64pypIQxWJXg++FLHC64WJapENQdi7UF1FqG
mMBD5lMEvnGhniC7UrTiy8aLLb1boJFkAiZ8HfHGBCXhtOq0JdqyPHI3LdAc8lGy
4j4yDgL4LiuVWpJaYVzzXmV09mpQgl92UobiqthbauuTWTzO156ngVkihRFcn++a
YS7EjDCiY6rtMzNu7vOAZx83Kb6/8YMyIxl3C6uE4CCCx0iXJVVSJJoHySURCosB
d0rlYFWSIWQCdL6nAuQfPjKylKbLcGJKtYh2LigRoOgwRVWZRJj6PqQ40QGd4xF1
AneLt5i1E68sCn9w2yllQ3sqspmvlvyghiJ3Hd5pwBGE3/Zif/Q3zOf3VL8GpoZ5
T+bvwA0eKaq6ZzQ+aXjfCZLysX8a7hoaBXWtb1GEClHwls0PRTPoi7UUx6VADB/P
yp2YDZov69LagbPa3jOma5jTa3kErJDR9yLzr0x4RexWaHWbPvNsgcxPjFllONto
rNTFAyV1YnvBKmiOl7R+Z927roSMk6ZHZoxdbEYx+whDc7bT2X5eTACetf15YiNE
HsRcUuIEekT5lE4uDtAjMvYKDH72WBm9D+6Be3LxMBDoRVifpLTSwVH/Fqarzx+w
nkVop/qOytnUUniX2CTbEsbpEf2igeiVZH1wgnyBBMWrs9rRv/J8U+pNZRuV3Ago
W1KWyPbnDiVLRoMAro2tluA89pJ9Bu+7edov4Q/i63HAo2dxlijCz/alOwKEokuN
mdLMVuj79l3cYZjMC7cIdvBG46ICiPN93z3Iq0asJ3mY8W2FhuYr36J1lg7cBin3
94S8GdobMA15k8w9Yfq6abwMJKkyCq43qhMy9Kaxsl/qhec+rC5x1yDwGLYOLg44
CClSKOQkv0RwmugowS35X0JlrsrZRLYuRjLFDPskN3ioT71zY+mnITTai+KjiyDK
nfoP2SxgRHh8//HfIW1m19xacN+xDRMyX1j6yU0IiyLSeTIqSvsMKQyy8uv3TPpo
iCkxu5tfdMbcTJ5WpDbnlmKy6zqh7nxoeXCpbZSSmpxR1in83BjbsrxDcfb/8dLD
AL/IW1QO297UVGsONRs3pWAmfNblkXNP+f+K7xbXYJzLreG8gdM1QXjyk8Ncu1gx
+nm41bJr77FYk7Y53WcNiGRdxhbVdKKTKKJlAgZ02xRT5OEof+wlKc/mRSrKW8cE
s2jr0uAUkZLf5/f6sTdpclVdFErOh9zJQWSoldNdxIvm0SznDUyLak169Q4ixhxK
Wh5CBKABY/FhWkXbWG7uYd3W0W/5ThYjyeESaIQ5S2oHYHkVjA/NccKBtG+9A834
E+fvWj/gtuZ3PAw1mujSm1G0KcO+8dlShu8BiSsZhWtxl+0lVfNV4G9Yr5UuG6t8
BDGUMBhj5JITJkc+QAmn3yO28RrFypfIQ2OeJN9wvfTAqJdaeSd0vd9I2YTuhh91
oCO6ATtLfdnCmKLW60P/s9YvUQ7I6rAsPQgwQ8DWiAbnwfVWxgQey5K4+fRnhhWh
UpZ2AIyuxwrAl0Wef9gYG7s7PxQzSKUJBgDt1XxYRuTC8gW+pcxb5SgUB5uTrG8p
yu7/VNanTKRrt+otjXQhtyI0JP0WA5IB8wonGqaixvfrh7iz14BlJ1ffVBS1X6KP
rp/KrkbFSsyxIE27diTa6ebQuWus8TzHxOqYKpowZB+uMk4iV8K6DTrb9xKwz1m+
to/QW9k7DaDiL1cr2EMDOsPquwpY1doFg/2HGLVR67rignqtWmSc9VmF0aafUNcF
cjm0wB56uARVw3SXbH9h8fkXhr3L050R1YN9ApWgmQBhPOx8PRVQzmzmYY02hsaE
s+cTGmmBRFLqvNklgmhO3qNwPxv+m91Nlqtb82sLEwnrRLul3kI3cZQDK2C/wbWk
ME9ZxNOZ8ORaJqpghm9Cf7XJ5amPJCJfe9ZvcN7sBYcXVafE1zg0RWJwmSwEF5wt
Z+gmnPwhy70YwEE9TGL9kljLTXm82a8ArY3XIGcPnGVgw/y/X2bs69YWGwp58L0F
1GCv2Fyh/s41QP1Gqaycs/Pm9hBWrWdvmqmcKIeYg3cpi9VcQJddxUt+pp62AoPl
zOR9VZVoWHTz5pq6nAM/G+fBPovBMJ1SqbCkWNWWbcGDgWirqSdsnqll4YVBmFnz
kvc/UAQe4YBw8Evjm2QghiboNMOLbmbKKIgJ7KUslAhdiv65aZ5OSZVPEHJ3FWFW
E5C1e/FusbIXfTcnCn8FqfGvXPYycNlt4ERCe69Pm1cBR5bvr9HaCRzlU6LMI5IS
5GMkx6YjtE4gydPPIY9OJmzeZsTweNxAbMHrHf1LY7Ei40c9FwKGjrpIXZApG5j/
Kl2Ys3Fv1kaUCaGL+F541vZaD8UMAW5/+zhb0A9Vm47JwV9PjwyyS66eHGdNjQTZ
LSycSTBgyEGxbBKCZ5VxsjkCGWw7LyPbHOZxVd1jZT5oo+d+/2JovDsgNs7j1ud2
uyyr82x2flOjgOQii/dLV0RbAZ23Aw6OeKTCS4Ix3b3w+6weeAi6uuhJg6H2727G
FEAYj5B10kVdizPWBc2QYh0qiqqKsyzPtdlgOli16FOyJxQIKcQqM/1RyJPZF7OA
DMKugII/AAaY1RNUHYVZWYN/wH1J3ue+mfoEHSZdypocHkkT61wWc5y4yeThITwV
YrQYu5TgnF3W5pqjyFqOSTJ6BLenMGBj63mQCtCOTMNa29P6I9RWP9w6M/NXpbLJ
AVoEByMuOxbdim078MG/HXv9+ECjqgSI8URtyRpFzTWgILyF25K4Y8AaVTUkyVX0
Oxr+uIYWodDLY5jwXW4hSa/hMtua2vQT4PLcGg/NEHJW6J9J6rGUXnQdDUVPIKcE
vDowvxRcVermzn90Q/RCYD0+qU192bKcrovDFlqFZhloijV2bohAUgS40uQ3a32+
5hbD7SzNg2Lnqfezljay/Thaste1XBKoT6+mD6RV+WH9VSadnY1E/8x0ezcDJnLw
+8nNnJsRN09ZIlQmlXKUi42v0oDWVT8Qt+arIJFswWNUSPAnGBKR9jWI3MPvMech
fW2qXrqDqnOhaUGX2oEnVrUvJteLBWsFfhm3S+GJUc3X4ln3fUBQuS+WNwzuH5xw
NWwqG38avSCNX1QGI3aaQgCC0x0FEheQ2tqjTq5nScTMUwoMoKwbEwbOJB3XSuwL
HngxCdBqoE1+Tdj7BECd8Cmnc/skJ8+2MFmFTDxdZNJ5oqZU+c4XxhtP0o9W+7jP
60aSC1htk7tc3uGMglksAkL4I9v9run8d3/eIsGsBt8dnbm65L1QriVdIhfunsOK
OTyzb4a8HD8RFhT1NuWDj7F9WKDKtJ5GSas+hcDHmGwsFqJyx68lXEFTA6TbcFgz
wcwlJmWDdfjB9qK911cGBh3ozCz2fSR3FQR1v6t79Hc0tWL8VhOVFzkELCBA9FrL
UngyFi4gCHvdwrz3m9NCWczilHPdmSIJkYrQS3WeDS/lHmpWtubzJ0b42dhqd5gF
4ZUFVC5ukwjLAShEvS2Fno+cVypjOXkC9R8CX21HM2K8LXdOvEGE/O6TYc7gGDKk
JJQnr88WI2ojseVe8lLlvF/cRjhUe2Lf6woseaF9d8bw7/4kN+orBBiCB9KoNZgH
9y2rng05z/DhpfCJ8vjELBERkgSCk1lfgXo6Nwgl00QOrO82r9gDPLC2+GslYAYq
S+XztLYcvVnDz7/VlDy/LlwYrVtyS+rUxPZXANoqqAE+Z7uSyhMUVf++Bb1MhXh8
4z12/SNH3pS/0Uj6TxBBWPhFFmJ/RVjwe/aMGHsMCuTpTgllW4EAGf7+Jqr0uf6F
8HWbJVLDucVE3llx/buwzsDL3BSIKbZqrXJxlQHNp7wim6QpyrnEcO+ybd9bzFuc
ZBklX1uETX3llHyF4ODi74g+2veXfPq40jQwkLNlWmjeq0uImFEVouxcWpqAMMra
DA/Js1XgZX0D3MqyXZxpz/tBG3TBabOUox83mBd4TBLVMR+vkEvEX/86KXzgcJYA
XizfYgDbVBpryJNRugOXAfEd92ttlUtlTkFv8tZka5Gn18B0afQtfVoNZdLdoTQh
tSUCIi5T/EA7ele/wCW5PyJRrbFJAFB1ApyjafYDyStUzKFhe81VpIueuTclvVXc
Sn/eDJuOw8U6TcKpQnTCC5vWxWSqZpRsH13PJ/XoezmfDV8UGpOm6des7kRig6nm
J/PAqPEZ/mH2NUyjMRJbbadvJikRgupEajZSDnkgLbh+BjNb/kg5ja8/LcmoMgA7
aKMDo/v/aV5K8F0Ta/pojSME4jrq5EkUEeY6EvjY/nzYpC3Q/n7mQfEVXT7Vpylo
re/4+Ds81kaUTUIFnEBZvZT5XFWHTZSmrghUp8OxSR8ctzO5p9M4Zmvj2s0i6DCt
DAi4dFdNaa2uTr3+CGqb7Fe5ON7OJTiA2rj+4lgZNbsriCVa6WBZj1ZDBCROCSv0
TpHxZgob7NNzoE0oLw7YDRw5qVJjYnu/cE71v0iOCdr5wZwsXV69koeBLtohYoiF
+FoxL7jxJPQx6s4zoBW043EtHenxVdRnEn6jDhlG0FGcAn550jAocGSQQ/scqAo7
2qGvmp9QHMF5SYjOM3djGYguJE5dFrQxvOQ0olSyaNdHlgUqKGwHtqRKDXjyCs1l
K7qjhQtVbEW/rpIT8BBsYmv5sQk+SK7U/LxrSA+9lcOF7Z2XzZTSuvlZjwNSm8o8
ZIbOFt0xZVesEw58MCL55xiAsrjPbhG7P6qNRU40uasLPPh6qsx8Lpr+u0ROOU/4
MswGC+Lp3m9Hm+Q0YX+s6v24v0cty4YczXZV/thZMIrCIjkKXwrzwJ/PATpBSN7/
nAZjX6/jKpioeJE61pumpGdHcEodaVNRofXDgPNIg1LCNjG53lrDEb2XVBXSr8sc
nk/cyog/6iyCVpqrtlJC7MzZgXrLlZ0AbqA0JpdQXyD0KRkodNQhEFzPI6EVpv9+
4cMpZHFeuovGpUxb/BCZwQA6kEwpDPg6vhXgcVWKnWXDnG1S3KFbxRhfHPJMg0mh
uUghYOOz0bZ42QcUPgEJpXo4cs2Z5rS7LcVxQKbbT9y/xU4iywH2OMHkmqYJ/rgO
Wqfb8RzPKtByIel76OkF0j7QGXiW7uCh0nY04IZb3Xl2P8Hpj9Jb1jsFQEmdHJXq
y/wYw1AlY2DOqn0CVVzLj7FaE2q829kf3CFtH/rt/vHlFa8f6x17DU+RNYeoa03N
fssfL5ZPbl9PHgZtIscmG6YLs4/gAQTDaLlLmwK17ia+W/HojXCCjOetOmfU/z+m
by4nEdePJI/VmSbzSw7UDkDtbjI35i2Lx5bSJL4mC15hF4ME9nLCoWO4ylPGwiCU
FKusGfHdSsbH/6izFATpLU1/pZrsl8XO94Pa6ITHOuPKKpVSgjBSmKCzlMT52zKL
rW+eToR1ACA6+J6aMG0DE2prCVBtO+VwlrjCOFn2zBkct9CI460NEKxUlsnX+KJT
SJNF2Fajc4xxBGzxVzqCZjRUb4kGn28ERuDmZETuCuVtQFEGGWo0/eZPNpee4Z9E
ko6fN2sKTMmpKaRVC7cN7zIxwRdfTAsrwxIdag7G3gBCcqnux59MrppZJ9ZJTiEW
C+NskjkHYxs5lw0fG3Vfk7L1kFR/6/8FFhb+oBgJ/g15kGl7trlb42YvEERxZXXB
C+GCUpNVSNmW5Gs8v5QAipnlFOhBNUhOsHH53eWwR7jDpQLdcuvPSwhiWGcifKwU
0Ez2B59bbyy8YovZwzqDAvslcsqsnvUZeeLmA0tiGzfaQVnbDtLcog1LimBA9e0z
Ob9EmZhCPERXwoQ+12p7AlLv+2jCusBnf2G66DAHbIHJq0byiK/4KuB7nui0iYt4
KmGxyhwQSgwRl2CpKbUh0WKDDKlSJ/syFWRzAb576cFpK+W1KgsRfvgUaXBNLqJQ
DZAciEb0rukSadvoIX+4ZAuGK08cfdMffyIBPcSc8V7ABUKzBBtHavfnDHQdbqCc
v/s2caj9+cTnbkClXsAGInA956Pf3eLYOBCtf/lDiYrjJEduk7w941m1gJl4/8po
Wm5oT+Xu6+OlFcydOkQHZmLemphidbAqMxBrxKjUgJ/rhqrIqz1hQkKJAbOxB7d9
cHEnA6DLo+HZgPUNFddjd/LNzCmPv9/xLlvzG95BSuib6kYQdFVa8jwR+I4aZHIc
A50uSPGnitKN00ubfSllrSF6IF1sX4qKEz89VguITkLX46WUbZs4z7kMogcwy8iS
91VNkdnSotzTKc5ZlnfGakG1pMounzxNdh2ieoif5ab+DfxdLghHbVgIPDl6vF1z
ELo+fyLY0xQRHgVpoir4fszA2SLIYePufFbCuc/7KQBJOhrO/dtyuyB5kpf9P79o
a7GBtHXZ2o14m1pMuL+ksAcckSNmHV4ZjV4MJ5cZx+ci6zKoHtOrsCWmzz7MnAHC
je91rjXBAkx/MCS4htpp8GrzDj3c81iJL1iunBp7lLRZ6FM5KbP0R4eFxzkOPDqh
WIEbrhRFPRJE9OVVVCVrxevFWXs/vOB6g1r0j5mUYFpg3UkpRmzErzAyjzii22bb
3WOpIuNhUgaDe3j2/w9V0Tp4R7L3pmwYOsfBGxQ6f9VE5Hi2yQ6h7uMjtZLIJ5J/
0nczB6F+lv8IgBpyV0wJW5J9//tN2bGIkeQYhcUyaeunk1fmQOyx5mg8EGvsx9h7
tf5uT5OzIc2OoHanUFNdLMzV4ZIwPNw0oNZTYt8vnzJ6cyympucGwhJVRyvAe96e
T/wrf8vZeKIGHsSW1Bqanfp1mb8EB0HRvtbdYE1f1lrLxYRF3W9k6I0tRTjkrzcF
RsSph40qA08x2rjPEr5LtAIUU4nxpQY6DCIZPJ8AM8Oj1kOxKkrJyyBHkHtsvOeq
FHUbmP8+hd7vHwLeEeX5PW7kkuawdt2fTrgls7en4uFOprOtD++bHnCbx/QonU3F
r4OGCwmOJmFTLLhpT6HzNiy9/g1QUIVlSIsk32nMEtBFzNE+KRtSYLrMnjFwhUjb
iuolHyV4TpkZ3jfliygy5Phq9GlK2bkOgoduwBeaiMMrlrklOlLvTVHIsKYXg6tE
H4VYehnuJMqkwgHBS93pTByr68O1d9sekuq9O/NBrTd4UKPKoe7hL0nAePKJqBrR
QUOGdNVEEcXpiSlapTv9OH/Oj7Or37vS3SC0KA2nb/BBNQ5jGavwzqJS3D9jQm8j
zwvpPtW2jCBUcbjd6s4mKCCNpRrqyJJ416ebPg9MESJr6eh7B1NN6b1jSYOrqSP8
qpZ4zWOv34PSGqke5vQYDOGe/ChjeAdRembC51Xbah+L10sc0zV4d4qKKDkEMI9f
Lo8hKSVJEvWozOVya1GYaowa9dHZNp6MC2E42CjUilnNHLjS1QclxL58BGk6TYa/
+pUXICLTy5lL6L7vXbnFVuQOUQRJhUkuzyRbpySUuTu1rn/70HcYH5JceNiaZrlZ
/3mqv859KN1pfYiufmw4VxybZrKjf8fh+5n2tQPfcyJMgaCiUA6fGtUzTHQNIjZs
gukrTyFnYH8V0yFmilje8b7RM4KFZioeKTyTRjqUpfPzpjSLXpIc9AL1cnsQcPbW
qNfYKyYpBt0DJ3TVi5xPp+7g5/8LryEwoUfwx4DulMS1KLf7gHfbqXsJgJiXut1h
mCb76HJhgHz6+7ap9IO2jxo0efs1wG+ZBjwIh+gYwAC4c9oRSvHE33FL/LHUD8hc
Dzd0XHREiEQ+8/KJug4qhaoqU71Q7DltuQHpBmhmLyXQvXSZ0LYkJ9R3e6Su65hn
bgwPZZfTSKT+LbXyygZJ4HyCLU7lidgcwvcOz+gf6o8GhIQw0QEMlG/vCCZX0fHk
d16iTjGO7vr9Yii6V5YbNtkhyoyO0fNAHW22dkw8eZ1U5S2qd2a9HMCYGhGsVA4V
G1t8/dyENKraWu8FRDF+A0W+bYcAROCzW2iIwU14vI1ITqAlp/sW1kF3m61+rqc/
jRgt8I041+cnln/3OoYHeXa+mjPfGTLJlhQrhf5xeW7FgrixjqseKX1W1mR5Ldv4
wo2wl3akmT9SM6SsvuPABlHb+FCdmwacVupOGJnfWk9hovm9m8NnL8dBvJ2BC1cs
uycx1hmzysuhtPvzHiqapl0ypoa6GGxhvp1RM4Ss75WECv2v0NEZUcNSJdkbJdV1
xI/cqbNrNegWzYoYrLiV5GvKwrkHIlgQhzHACzeOVHRZr567D6Cy6vPeUfyc2rh/
Asct2GeUCT3RXjh3oLaayaOqkx3xaxZ44SCC1C0nrByB4RrApKmf7z2TDx0oCUq0
ySjjr2GNN2GF4JGSZWiuSWiJjrds/Xi9625hT5dn765ADpCn+nAh/kdIYxZ62Bei
1kSqTapV89qX7bBgj+PTH+vI7Lh5JlZTGauymd9MrIBpY//sbzavMp9Kd8MfZpY6
wG0PjXEkRsFfi19h13AG15bSsrpOB9V+9sMyUUUNKjaCC+rKb+DIYfyGGfD3WqTu
mNBVUg3sAJCs7k8LUfk84CE3rJ1EM3SLEKRH+geQyFm7txA+oScVWQcp0+UsUfwj
s8XvZrTy4Y7CGHOCRuyZncjYlYwTJkwZJYAj7NgPU+dxputal9LRBwodEOoj1Nl7
iRsUpRutPwJsR/U8ZAkhLgzDdBOptASWfQJ+Xnv8FA87MBYMYsjyiuFkSBRxc0dp
qC2B4JbKJahwFxjoEhlg+IqVUpeYWOyp8ea1ULgTHVdslyv6qPqgHwiuabCWp5ed
nsGSacllcsHbUzS942UHkzRsRedrOwNix9yg8NEMqi4GreCI+65VdcufJmzb07c8
6ysWSbuHX5uz7aKpHSdGBL+It/ewRVXI6Vgx2aqQaXggv3mflgwN2TRVuXFm4fB9
gkb2iAlyhOTjTplYqMaNzgDBjTkjQkdPiVnnlkM8ZnTLzzMKJjksTFN9Tzh3zJ9T
Mbj2zq4d7tRznG61g0O+FN1c12KnZ8rNJN+jcfJES+qGUIVq7Lz1NSRvAcH+D1AQ
qEuZPmwTqbQCeLSPfQq0f3pBMeZ0UZpE/yWMjCyXQCFmjZnPqyJjuMt8C5iHjViH
1k8nImkuPVP8aLWW0z+deuYwZyKh7qk42cUa8llMPvkG6tMMMEyL7yQukzdywL0x
+cMsF5u9H0HXBZksgB289YA3EahPJF+Qso8+fPVPUMvHDy4KJ47qA0KR7m8exFyN
uenmIYdX/vpuGEt7DgLMEs1OmfWvIYvRIJr9AgKuqBf4BQ6GR6GVAJJ4EfZfT3EZ
eLEsZiVScCkjmINwH0GWXSBhBCqENHFgKpYs5WhaZTEXKxti85tgXNqsaP3k4X9A
/hClhF7WOIReTZdhGOm1BUIsMXuALlqvAWnTbByN20VCcljGwej9NDif9QmyemfZ
QdIm4WP1mebOEp/IamCUvdjs9Q7VHGjdvduVK1mKLBZ2fzd6/5zSA42wKQAqRwin
KM0Yvg8JBTj/Zr+XwYvXyPWixAqpQuUFZKxP57VL8h/9JxMmUurGIy+OAaQLClzn
uq2PRmuCmfc7kL4HzhNYoXbFT3yG96pwte1g45HWDf4epxbJXYaUVq/t09Em5JIN
ow8DxM8u8llKZFOgFXBLoxFFt1FM7GzyWux6LTBpdYI6NnqiYLd8xKyckIe5syA/
kHnq9rkGRN8Uy/gNx/xFOTsJkx9FZL8LjR+6r5AZreAdkH2Cpz17n0GIG/Mu1rxV
bGVmOjscAIps2K6h7sZ8pcQgUjFApS/+Z3ZXBmVqOu8l34OOO9eQRFAC4XgCU3iD
sHj6tisN6qCNuFye842isJnhG+3fYn8c7+O+VihZMbmS5rJAuRZ5qBHRSy8DmYCq
mK0ZhjvJRIMKOGEFf5Z5eRakKpao3d0tZofg2X0/GsSXByM1zV+edgcJSw3hGbHV
XelgAjakdTgE1UtMMldn1HfA1Wkqf0Gl77k/SdeLKUlQgxIeAK+WpSAH4dzad3/+
mLjNM+LKpqzcI8GhKrVmvXyksJNEM3sOwR1bucKM7daiWEhkVVTIzXxOO2cDIZ8s
qm26mFBe8F5fKR9M0yQPwjISNP5+M5ZctZmPQOZWX90fx7CRxMH3sCrQe5Nfx/WL
72/GOWTPMz/XbrcPqpwZP5J7uwONQ4lgNnf4NzzoIW33+CihcjA/mQcUp8cu13QM
5malQrdoO9DLHaDLgQI8SXHbvy9tx9nGbbKhJ7Zcmh3liyE0UoOnY3/rohvM6Ncr
qapTq0j+1/Jb2LRbo/zN4gJssxuZCJqwN4mJaH/WktKpElGzVtskZRTadiReOaMx
NDw6EWIiqd2FlgHGmeT65Wt3hXqYZHqq8zKAuOEbV2yu1tGJijjctOZwn7dvw24m
wg8PzfVAGmHU4mlp9ShNbSUz4iLx4/8IGzapDSendrFZcqYAauPV2NF+vAYGirc3
hBx5KrighstdFp7cgM7dWDsc1cugVEtLtaW3kFJ+i5ug0biW0q1B6zyw5Lj/wU77
xSG/BNFl2S4RNQwcfY1G5jEmuseb3CXLLD8/ubKXHwnBO4vIpUySVGLVjmTg8jp0
QHetlel2/V4VoXDRPXP1FKj+iyuGVAq1tM/zvl7+oeQ2HV2MgBCdrUB63DovQVAK
00dAnKba6qGxDuHO4oCnbeWp6RofhGg7wMjLNWS1NRE9gWcJ/VT9mKfFbleT6j86
hDcTp8YwasHBwrbhqhmxZrEN+c3mgWfTQQU77tLlhuM9rFff2+majl2gJBsPHKgL
ZyLnn2PLVA7yBChdbMXhV09eIC9VCjxIxQjEoHUR1T4o+FjpgG7I5YJbG3O3RTez
q0DP83GopUGGkFtq8QXAQqQsJYzineFpxdYLFAi++rvDW66qtMiPmlVt312nv5zw
V8J/EEYXcx4vs9xPJoBT2jml++LSTqIBxZU/yYji0ur5z8EtmU5HWGCV1fgMrcao
NB9CLdfFhljLcFFKk6HOdwgjiPMCrvDy43afxdwpNCsIp+rPbevv49h3v0N8Baxy
JEK7dFYGNERsVfp2ZZXsNPL58kp3mAEoatFn03u1c9YkPZOC8OvD/94yne2HHJwD
6RFJB2Oc3hzkUvW6lEtPiSjZCyC3EEkWnGGNiCv3gmeSZ3mnmzrEmud9NEzYb5NC
zTckNSF8Wdm8SpcwsyW0J2iaIaH2XNe9zql3gLErE5DlWyNezacVB8kfodPLQgtD
c70EGTDC9SxAQDwMdxJQwqEQEfu5oixe+GiiwwG7/j4YwQjMMxTsX7MIR3N9Dcd/
enbLj57ZUq2NCipswRFqm5QRGkap0tUbz0DxCHgJf05EcYOXk4K7wln6fG72qIcm
PszqEsJMkWTBJDlXhfgDw7nEiqsiLUfFvK45IQRkuEDrq1fpB7cEDdyqerokVYvV
DjZXX8tGXoZR9Arb7QgOH9gesyNP6fwJWMdTCBNTI7UZy7PWzInpyR1Li91lZxzt
PYPxukuK8c1z3Nk+j9Qijyofnzp59HdqR43qFzW5WpbpbM64fcOvhrtcaFGY0ZoJ
zGbGc2eYCYczZIzj45yssWqEBwqweD/84FzlzH2bwSjpGza24MO0AARLT1yWAsGP
DVOoxMRmdARflqW9zr+Qv9ylegjqbk6gWeX/dRfOf4a/gadt1BEhjxY0S7NtJ3rd
E0PVd4igdmobIYvl8XP+SRtPbcw+VS4s7kAj7qt61aAkW8NtAd6MWq5YalQe1Mgv
tcbdQJPENx2AqLbnVVMEWvbO+Wwwcr3zfEosK+0bKJcakFNmmBZ1Fn8+5M7CengF
Sgp11Mlue83mZacutsZrov2PKLYP4dIsLghWnNPGkMO1JgN6OlgIK6MxWfqQB8Py
o4eZ0LcOXtSo+bm4UXJ10Q2nw2udXHULlbuUQvn+9rP51pYcdLthvyTs6VNprzpc
1/1Bfz5VY4kjzoVFFIF/wbM+FjXTvwuHU27KtofHCM6uAo7W5ImcfkTXcYPUeLDC
/raK6LNfsmYNMQjt3Ui+ZfC/Zuil+F3h9Qy42D7YLRL/vPUn0nK7a7pCHPI18cvb
P7Qd+KpKar36G66cHCVPa7VvecmV8QG0qFF78xcsMj8PoPU/8CQRAZWe/5jaw8N4
LksLbCw12fWub2LEvVCliEjjMgpNL+Bn130ydDLSa+SvkG4GehHgOL9XQeSYeCcd
SUSf7x+0pxvahHKQ0/oLV2ZZenyPX089oA1hOe9mILJYBwHi5Cuk7y+3Vnaame3w
dtFEbxm9bL89CqbvLoGKvXBFgCMMhIIVYZX5+ytH3wpZoNBtxLtk6Dxd5gWbSOjj
rX2o3c/0Bn17zZPylxtDTOgvqhmQDESGm5dZI20KnizsT9FYsUXUdpga6oHLAuW4
+n5WOuP+IxFXGCmfDpe/fwzDuS0syFTqbo+6QWDhw9tCmRcrOwvGffe7l8Ok7FL9
/GI2qCefAiGXkSEJlgG0RVgLp0A/Y88DOervzF2whmQrs48DxjrWh8YyIfHy1BGA
2WfdNEmXPJKbRmlPgiTExJJPdMJuSJfkhancTNsoqYP3ZulefydyaLDIQBrF9Hkm
RaMJ4MfdNxtJkLScH6+ZzuucbQCVhFV1IGZL6+lg9OOgfdL2YKOxCUsCQDG/tA0k
KR5EC4a/vpjiIfuJhNFpb9J4Hkx9icONPlqPhEif5V26TuR/UqdoZTEw9YOxx3CA
jO6xWdATL/PfA8FI1MPMSAUZZItYW5Q/Kxk2QjD9eGklYIKMz8GFKatLj7Zg2NZg
rwFGhNn6MdOjW1W4/2lTxAPlIIjGeENS3t91OmRURZv73X4fYhhsMsLz0kvSwNjs
cYGQKrnPD41yr0CfrgoFC7v2Rlvt4c5BwIfdEbn8CPgMw5Io1mLYCA6VARGqWTFa
1iecmjVqypi3PJdZcTK5ihcrjKfTTHvHsyqUvUC4ynUy2C/lxiF/Qp7sRvHabQbv
s1fK4+aBf1/9DpjJFtcPVfyb1eyvGwFZx4lYwhxZ4PWd/AIHvwYlQ+kz4OJx2hmP
DZNYq+Geu1XF9lWvj0XzmTasJC8mzQoVPAcy1X1zr7IUjo/lQFofFLTeIxpbjP4X
zOyosYIwatQsr3kPCaheSheq/XG2MStwNXiwqhnivztQeUwocIYueWN/9Y6wdHaO
t+d20IF4eLiuS+qarRhILb8NsvEzZXzEqTKcn1pCkB7Co+HX/IwLcQLQNQ6DGN04
QoKt1yGJbEHUtIl23ycwR4qjHUWbm+ZuQjzWiKBkyQPer7XrXA3r8KEfkbKSCzOa
mfmYuPyHCu5NgdsDyCQcjhNny4ndwoMSNAU1Uyc0LM3P+dQkyYjO7QFnrdtjq8/C
OtwRTRds/NX97PgtjqOZIba1CJG5BKX9iOD6GfnfiNtga2qC6vAGnxXsScwEX+Lr
ZZxZLhFO6LWi8ZRfrEYT/o78HLAjr29ZYioXs1XZ2WjygXjRIV5EeTXFGR50gouo
I5n6074/HBAUQsBJXPKUqI+0JGxyVRvkUVJmQXfw6vuhbx5TeyhPTBBYBtXHOzVJ
8/zys1vQnZwopMoAp4LXo4k/HbeNoUx8SnHW3K3dC/fICOHzuEA1wUExhqETcAF5
lxXo1gKvNTaNuz+ApjzKO8DipXvwJ07H8DIp3Hk7YPo1u0Wi32pqq8hz5h4/s51t
0XA456wC400G1T9+CFy2bsTUYjj++6pKSi0i9bZwOj6HYq6gTmwmzmOkiot6Zn21
351WCPk8ugjCJssDuD3Wnvz6/LShJhThDieo5BdAt9NA4OZ/n/cKWyoy/YZjhde5
ViBspZzKenqtVAqkTxAsjRk5O7BdgdymRuyYLijkIsA2fwBO8wDaCf+tEgNOJm+g
ZZ7K7UU2lKYwfN3XAvuReINi8RQ49Rwk8qbivzWKOEsNnM+KDvh8ZAChiObArNWw
Zhx5tPh4XkaTQr60+ref8xvMqAKQaqrFjJQMuHNkJyTBTs6Uy3KwQW8TRGo/W9Lh
hjELWmVC7WqtRs5arRv7kqohdl8nhbuChgSD1Xyp92y+siDn2FcWv1qJP4HthmLg
RYEzBbXuPMlQW/hxKfJBnAtxaAXIf1lB6zM0xV2uFPnQa2SCphreMqmOlxwXAgyY
a1GHSNnjRVZn+5G3O2FPD5PvyfYM7PGcJ9/ecBPSgJ3OWUlzGRssMYl+zNGmxwIC
wiHhLali7gz8wE0CnTOfNCGEUvmg3s0QbUGU0oyQHLjtGlG75vQSnzwhbEJbXvaq
QQohiBoyfzKC+Yz18KE4ZtPq+RBBf649SrzufKuKmGcKi92StG2DOfc6v6ZcvpMv
5smlxkEGYK85MYGL867ZcMR/354Pj1aT5r4NIN/AnnAUawwFqsyQIu/wErptdQMT
BV4NaqlDEMdmax5gr8JLJCGdOY2q170vEY8SJcHnn/xN0WzZf2uYWWqtOA2jMoRs
GakxXoNoa+jQmlguaTggxWD5lujUCZZsT7l3Q3+Hb8y0YzRS+RgAqw7hCvezxcfy
Bc/rXPsgStZI0xJf5LQjYGJI3/r2bmV8E8Lu3oy/Wcwvike9ecxtFMUyNTTPVc9u
AIVBvoRz25JHaltEJfvo8mpMPwCf5hQVyNDMIh6oPOnG5I4ZW1uH2RdiHRx2BcUi
BqXVvKl3onWYU5tswlbKwOG+u9tELquqk4bWv+6aLNEZ+qixAMCw2BScwpj9PAlL
4AlUXugHpiFFJN6ewIHwVcvXyIMw2/+HqAwQbM7xcdkf73krfeRSXNN3oDXszfxR
zNp2uzbzxhSDAoTJThZGgM1IwgKSyVxfk+vdXj1/mTF9h8bMGnH5oDdMLTqveZBH
jys7JFfvuCLbSl6673kCUjV/JBBucSc3dhXEJvpmuWbW8GYNzID91/iNhnRcolNX
fJWbh48e/8wumn3i3O0fKLj5pRecTnlLAINoGXxWzwe40HmgYkJly4RoUhlqPSON
YjfVEnqtRP9DiD4f2amJ9SSIW7VslbH0F26rbLeWJiURd/e+vT1FIbztPXKx7bdw
2798PRsEGPhPHK9S+JLTAUBoe/Z/ofE4QV14fsAw6qA7Rd/cqjyQH8tOXNVPB4o/
gXEf5POb7Lis8Ul+FsAfrHLi1Bk6qIdyWjBI20XPVBZckL8/0qN2k++In/FrqblB
Y3w9mtgwREORRdlzhggNeflsORod06rWaKMhQQl1rVdHtmjhdbS+p7GGjovHvJ9B
J5VtAVnP/+M7cfBlB7dshncqMR+c5ZBmDyPC0ao+os2RdposMUgZg99bgxk4D8zD
ta6lsRD5qW/awYw+AmiTIAU0wIbyE5LKpYwehMSIWe02qEBoZcyFJygyv9qjgD7j
fcGZcExDdwSu29Y/m9GvZHClHiUusOrYPeaJS9/NzXcKiEy4BjgVZPaJADvuGBzw
+qLXf1fpt77eypslpi8n9LTusfjhwqiVH8nO7ToYQhB4w/SMc+hLbWvyAcsZa7oW
llm01TtS8QY3RVkHYzYTDEeJSs9iwvSlms3W2txUSjERvpnjNso/umTbVvlT20S1
PQHSQv+P/M1o5sYtMrhct0wVAQ5iG5ylreXe3BgWb3KruGNoDcsXkMwLCP6KDFiX
K0H/EvmJwuvSgS+7nIw0h257V3ZzmiLARsWANRIbmTITRXr/fO5T4/lg81sLFTsG
Nw59i1UHBuSll1Feq2eTSdBQ9gvUuPuL9InWOPSAVThwwak9kpAp7dffedANfXHv
ixsEtCeyVZL04IyGthduxG5bPaPePxvMbENf8Pt7gkHboCTPW5hbqBZmQGLDttQ8
VcsCkOFgroZ/JyyN43eaprKyoufTWa0Touvt7zYH2XHlyBiaaeMw45dOUprfHfMa
n6Piq4w4Pq33gyAAtBLfObFJk1MXCpA+vQvJwfxGuj+ijvdAEGHHWmClT/jj8Itz
oRLOLt7I1mAm8mBrCoKi3NkYK2ddQ3O4wzrsZdESNV0GqmD9vEOmNctsXeAg4gjU
7peJL6pc45WK2KHFm2f9vTVsV/rZ4kDDylUbZuIuih7IKJUYYvN+ID8ntf2KPovY
T5G1RfqtobMEjlKFMAZFVBAiRpffFIi+o1KlOmiZvukPHPbdOEOhtaexjckchZTl
Il0eA/UK0oPsvHcVMZtAtkQjPfNj/Dz2VeB7JL8hkeItFc/8FL/wDYocJ+lHnRX8
sj3B1Hc8iP46jU9OycOxIhY/Kw53FoyWLmY/7DoujYYBkltaxD4LPm+B+bLd3N6R
Tzw0e/HFYIIwUlptD/1BVKTJvpHp9P7umWzksnu/E67mycEDK4th1CU0xg1aHdfJ
RDE0E+kYCWGsDAibSaKAI/HkocIMaH33ozOXPOlvQPKVbJG7dTTPpDoaaHunqeS0
0SBIwab3NckO+cMf127Ibl9dOJxeJJJ0zF9qrrHiJlOXjlMksrH6m+EUlA4SA/8X
KTybmEfsXWXkwdZt8TDPbymu09BtkTvhkKM4M5tRv/0r2yN0pc7s/ODHCJARGzUd
H3A5JDS7wy9E8YqsIhW96Ao6sbTSRqUhnOPPlzAIihFGgPWIsuhpPaeh9FjQXPd/
LMIJUQ+/J3xxRXZuPUdzP1kKJ9FAi10AtyIo4y6Cgxi3we0kQFH32dg4SE+Feowz
KPzXzSxgjuB0BU9B5lc32OIclTcFvBv6nGZigoAUZM/i9Zm7MeT0NGNRglQadoXi
o1/RSkmY7+z1qV1vBMgc1lRVNSai96FP2vbIRh9rFe/0cn/lPQ/CMZoHNrxAnWRG
GMloqpVB+6keovJ+xADynYVesmoTyVdHuIAH3+Zly/b8kAQwgRYkK4c6MMTusqJB
1zNk0NPBWP4iv0WiK+yf7SfqDXE9Qm7QCeFW5eVVbItCZRW+jmFPi0S30XWJVmf6
ICHD522neyJJFCPnEadYnrSPT/F1ecF7zaj1XAFg7pNYtdjbC9g5lpQtdPXWx417
/WYM6SmLmbBhTM3Wjx1uq7vRgybtbOqg3VR8DUXZ1A8khphST8N/54CSKNAmWou8
XpOlOfDzhKRafQMHGkWahPs0WwntIgbro+mD2XGwKOukJldfBbgKegSeacrN/NhJ
koFVzhn5qLawexE0gTXNF0fBl5hchggtj5M4YqL212ST/P5b38Bsd1UURgPWdnoP
cyxNhPzkWgZ5eX4ckgrzCnelc6oze+bhiwxnMHW9elD8UtEV9TP9PakqqxK5P8yu
2yzU9zjkQiOddqw2sdHxUL87f177Mpf/iymnIO5C3bbYOoT1ukm+ZuitGc+Yd2C3
/JgpxwHINLFdGiqsGl2gTnUu1Of3T1if5L4paZ8O+A3m5VRZpzJBGd/sZ4hwc8yx
gHxu67bnVUC93YVjc+EhQwjpzp+QsoP8MLEvHejiEuIzHjU8D6q06xHv1gKocXPi
xTice3wEv1xqEpkVtAj2KqXngf0QhFehNjQAK8jU0Dy587AehYEACWCfIf41g9Xh
vMbmUa/w/NYgbzIn1H3WaXzZLVr6ZvnLRZirWIUFejSau8s+fyVbPQPJAlW/6zz/
h6vp+Bfv1kEOwGL1YN1WBRzy+bHkhGIhUV3G+tLM9+b9+1ClkNOzys1PhNxov6RU
FxXBlFCjcQfN4d9tvxR16JHhZReBwEQiaIDJKmEoYUGciB+lkhZi7RFUeaPmOK4s
sEyQ+2BVk6NPPLXrcbG/uzh8MQ9FidYsgSXHMT1e0ALIW4s0Ew9TktLqCtLMTWo7
Q/u0OX7YGVdK38CH/Q5iRcQ6P1vrMLnXffVW0XrC/BR0cmTeVA2XcXTmn+ppH5A/
l29ik3ntiA3iD9MymkiQs1MQrkIEoC5MNZipnKa3SM0JINTVjSxpWMLDYgHPlpBC
l8+vgZFfKBl28BNU2ZeMGuimWtbGRUBgycpHpL2wH3p5iHx8ekSC7pcVLlS6xoIa
vmOKIWjhZSFLpNs3iTCbeIi4j1/VGgXMA2l+pqUNe+Z/QAU0n2Jdy1DpXGxCBWCf
IC3iXvH2u1hLAft6e7iy5ekCDHKVdORic741BSQ3Ios2DbIxLwfjaqjSVUKvmDgq
P0QKwdNNwta7LF8imn2/waRLH4qGIIkh4J6EuyIb/Fsjk70tIJ9F4h4RZNqS8/mK
Kc7qywLhZzrOyrIyi44WlSbarZyBODUd0EQwaEJhb+VB/qcWQ5CA0Kz91DOnSCVo
bhPmiwlTKkh3+jz+5qbD0YMU74yNuV1+5785Mh+sSGb1ssWYjanQPPOV8EEDWLgS
Lq/ghyhANiudmYeYF0C/0euRUXpmSvRRhkAyf6iQV/GqReObU0orQ33DXsJerrJ9
iG/6nQH34QCs8D6ohV9XsjQCZ1kQY4JF8Hi+SvzOnPrZj/nfDmJD9AGVoOdhEb7b
c8YAOeG/2Hd6hCMauvpJW3yctp/J9bVAkLTD9kVvIN/jJtxiYCRE4uOt10oAmUrc
DQFcZ0eNXIgzWMyKKwXro3Uzl/+fjIXLTquIon4HU+WbbTo1Jbq/v6GyJIGIbcI3
8iBRyKL3Bhiu04/8i25gQJklKnloT1Uu3c8wkGdbC/OZqnyvLVicmq433IjpRWwm
WLmD9pmLTXDihzqCejLo4iwQfozfAsrJSNny1TvT/DA1iMlZrlCkMvOzcdFvZBm+
xPeOWZDeVhbRphQZMeCKY7pOY43px9+ckSO0W4Q4vqLaKr0sR7NZoJTRwr+t7KMr
e4Wqv8eHCZo21P/BCUd2WKdfvgUIQGa6+1v46XanJCbLhdOWNdz2Yf9u+WY7wsoS
vLCv+CykQkLCeyZvLQw85ko7ft0ND/Rs3HEFaGIUjits5vX8tr/Hs5cQA0W5a9yz
cjpm94VSo1j4NrnGAa48lrA2VTBRyyppBhsgfkWfpspNhVjMeHz22owlkwwe3Zbl
d1C67pU25OOewzSXVdfVUjKN4LmU1wkaNeH++mQsrZzfJkwyGx6q/mLNl/Oh8yNm
t2J5gmrk317uNLO+yr0hgVRNk3CJM6uGvMawlW5AoNixFlM44abG9oyjxOp8/TnA
Xkrcd24juwmx1V31quE+z1wbPYgqxWBmm5W3l4tV/r2mkfct/MNYGeMqcDwbyzK1
v/LPQy0SGnT6QYRWBYcxGT1ZUWa8yR7IyRz6ZYDjr6FO/xhhJlU9d9BTeba/ykyk
f71vqMMz0JCuFh2iJEyf8935DrgzDUyUoyeOUlrnS7AZDXxZZ/r5+jXS40XM/HZh
eWHrRLUT2SmzC3IOytSaA9wztWBa2JsxcFXnFIso+OTUQvFbVFHZvYvXq1M4hXkI
1XMKHVHLxste2KhcecCjwjLrFpIyavyx2OcSqCAHSrVI8SFLrofKNl/KBUkGo7Ed
VFM8Now92p2YVAEp+zNKcHOxBLm8Y+5ez88misFaiYaORYMrsnhs8YwN5z+399SC
I0KDM3sZLzMa7F4Qlk/i5p1Ft7E5/h/FiYJWp+nIpIfLUrdBLXt1a3SfsUiUxOcr
ovcFnbU4Tml+4N3A3pajikoY0AirgxYUGT7QcldFjC2k/2n//ImU4FKJWdJJHJAF
qxG06nhnZnQGalgSV6eLNY13v67ZgzEB4RbQilZDsTFv6cjOg0rQfqJNiXsxcyJ9
vWSmLxcxmKUnTlmPt5WTJvPV0Eftn6pvGi27BUkKYVJdUfBhT/vXcd0ImmdI3Aej
tVyeQ+aJ/4b8hkYylrZCbRu3sY7M1DhaOMRcVyxx4m5W3QmSCtWtYIXIuWANR3sw
i9aPah9Okp6ZyDYh1Yb7/Qp3WUfomdXgw3rzaTlxTwVQ3466+5+CxRD926dJKRIR
LP5Vg+TuEI5fTYtvA3Txixq+QyqCneVHPWaB3RdN41Qqcq88LW/yyevz71Z2beeH
Pfuqkbg6YCuyvoPihcumKXcxV7/ozI4v85IjRMT74b9cdphMVlLNeqQOqZz7QgQu
4lw57CIFrxtQy5th/IbQokvV2/iQiOzyhJ3GOFDrOWxXZvtqTrLKEFDME/UOe9Ec
535+SDSr5vuMim5Lhx8DMXUP8dL9gArbQhf8dcYLJCDJGK9LcRS0vJ2T4osPhU25
U9OSas286GWw/KInvt9Zt3EBRz0u0NiFZnSXdbZDnQgmf3stjY27+VkazUuMXESd
/1BM+VRy78sk/Aqs28OQftKWSF5e5OkdqORsZoi87pbqAwHwgcWztOplsUMHr5Mn
X8LEIvqTliq/fl51/jYFcfp4pXfvucZw+/AL58LDqJQJnW9KGFFkgfeWIoKO4QcN
/TPppxI5TZePDiObwsQlYaNbeNWU9bIv7QUd1Jjqz3zaEqQeKNzyHyQArVSVCSTg
PnbnO/CFPqQHDKux5S3lTAaVy+x7dG2L8DMHEMfPm3PJ/cJG/fF3aKnvanlxD/mY
t7TC2p6IRZW6g2oKKu4bEmSpUkX47FLKZVw5EcY7tNuryBFbWAzcKl4C/gsoAh9w
wl/kJl31mhvzCTE/3ManlS9y/0gd63/ficqxABEUOLD1hqsLGL4g7He59FiA6XKK
LkFzxMvnYpL7BTJqTmlbESCs84uYXKPaJS927R5hAFnxY/Z/UvGFxxktpzb2V+Mo
NiLVOH6kjtU3fjqaSnHCKYgP7mtAlyJ35LjB57O6+3l2IKN4kJOWbydXaLbbEi70
Die9rV/J0MVrRYh4z6frSBAGjVP9upPhmVUEdqi8PETDa41wyuNzkTMHelljH2N+
whBCBdFDc0HILc8Wmt0HoC6cGuUeliZDa1kNaNQNeybWWCEp20CiVFzxVmNo8sX9
YfKk9Fads+G4WcTVJgC60yUedwK+/V6i8z8wHHQSd6HY/NeK5Ve2kDANn9xqGOeh
jdUNkY6aSuxqv/hyzXmYMx0JySuFjm3kvY5EKH1QjJBJD507cxqvp22mjoJ/aAID
B6oKfMPEKnxLGNPtR4iEueNhUJlZMWSswiHaxAb28P6PSCTt9Fiv47FgLVArOcxB
V3AZZXp1qrLYCaonQxC1lXvxc6/ze7sOEpiw4VvF9c+sPWcPgoA5/o9KtegsP8ts
RLnmL9Dd8DXBxzgj4UMko7Ms0/FtSr64qiisvg8vdgkfcBpiEWQ7Fzr+aSV/cItT
EwsYLLwqXfmAe2Cbm4AFB80mcGraXbAXWZmpualnnYeug70RLybYHHQMUGmxfxj0
ayye/bhfYhV7DBgFQYWLEe4cIb3Yl5B0Z3zZ9uBxrQI1jm+RPOmTagrOEeqJFZim
dW463+Hy8P0guuXFxsMxvtThF4W3Iu7DOVItg0VksFHOjsRcfNnOWpNx7r7NK3Io
X5fa4KEWIUMMMGIdERosB0HXRYO5wJVbSWZk4cXTK/ZRirPIv9TmLYd1bM5J9491
d2UMc+AcZARz/k7eXaIPKA69ImabS9zMLQWwhmsrTuj1zl20NPiIkXz6FRV38Hie
lg9uJw41qzPxGjqsGz56WRMcZ0EnT6JWyTjv7Fo9eTFU2fx7xOKOydWBRlFlTNi7
3FPbKZp7mGz0b4PnVfoPjvtYzG89g9id3PvpKmN1OF/46oQNwi61/RMlUet+WFBs
z+RXfw6LFTAUz37L1Bjre5PCls/IC1Gh7Pi8DXbBS/NLMTNh64vkWC0Ph3+3ctjL
2CTd6nEE8iAxOz1XqaEHauM0O2ZNJqi3+986rxhVv5bwwrCz73M//V4MeKMtkGMf
+NEGw79ypFGY9ejnpWeMop4K13BSxxdtCID+ibY0Uk2QdX/J+gCInfOoNVm5isEO
ZSLgN+8g0zTPMnBN1cfzN/6I8agUclncQP+uWo/TAsrjkDUXsEk7q1TgrUDEhbXm
ObewYQ4nIXVE52oF244SMEMa2Hr7Q094Gtd3N2qyO8xz7Yt/g2HgogWEWGgc8hCY
AgA94Hd3JTIcxUaUTl3C0be6PqK3vCBd1d7/L20+HWyGFalUwesr8Kr+X2mLDkPB
9ir5USZvpOzLrRhkBlolo5igeh7MDXYK/u+8DcMaDZzYwFeGDmu6/aKtbi3RgYNM
RQvMkdIYDf6SSspIERb972RX0/cSyn+cTH4Wo6Fxh4OD1DHRvmUwCXXAuPn8P1+s
BVdydOoO4DWJEdqDJC9nvuxCDNlVYM8FYEo4tzwT8cvtO5oP/NSvKjexDpU4ScBQ
XBswyRVkN2JBgrPFD+JLbrV+l7YfI12+tuAeHaU+znaGrYlberDnN3JLW2wae9p6
C6oCHUETfd6O6wsyE4I5lYJ1ZJIFc4hCphpnbmZSsz7LTQ0l7TChC8HvXmmlchje
8/Wg37Hz1+Z3ms0/DZcHyYn3LPqkXxjw3LC6Nl3XXYTLTudwT/EprWReEx1brHeh
ceMCjbGTikEvjfNE5OWv2P23z11r63AnmLfKHbeJxJeB/u/7WPlfMmMu5dhfNo6a
kkKnb3A2EhYOuj+02avCv6Hk+HvAmCe8xCGx54Zui+MoljeHc9XlZ9M2fzyvCpR7
DJzXREMVysaRPY69yk1kAenwNw9+pxoTpKtsZaqC9wQRZeqtIcH/OAWbaGY58LZf
R/gqBG1Y2IuBCDQ3/Sxdk+XLircALaX0Cmcken+CCbbdVF9mNCFoVQYXpDhHmzm8
J85NnuZ/J+u47ynRyQuoNZ0lwLgD+GcQBFznstbeMCMA+GvEbagWBoS3z4cnGrp9
7sGCvqokjB7055P8nHHkyxuxQi1VAT7tXZqAPpIBCM7iErlKuvK+0AZL0s//Dmrb
djhSfGyE+NTvPHuyYXvOYa4kqtXSRS0zbd4zwI2TxWdPSdS1zJEZz5T59NEKwS7H
ACKhCgV7kG6AF+ewp81guqCH85xn/ve2ujI2zipVZOYVKfvlBYSDf33rK7+/DfR1
UMpCNY4Nbesgfcyt/xnnPE9+bDTkKQyHJ4O7ToVGBa2YeYI+7BdC/W0jrEdX2G/P
D01nrKmi1Ypo16+r5n3afYZTY6FTEQ3RAxlJxtD7eZF1AzzA1535iTtX/383tdmr
dCQ5e5Hrt6u+KlJmVcEbyu2ji3FXTtZyLlBMPTxMRnn5P5vduBfJbAzNXDIhkDAr
/f9QrUR6rxF3RiaRTPL2drT/1Dqlx93mqJgB6u/NETMvGpy1K0p9mq+az+yk+7vd
T2eTKfPSQ9CDVpVPkMrJ2Iu+4w00fI3zbFfbe6lfdh5T18cXm8ZHP3p3sIxGGRmB
B48+yhDztkLum+4ZBb6R9BmiJJvSIxX/UwIZXCF4juCXz5KCf84Kqn6eP2tyZJo9
1YinkhEM6rHw7wi+udTXn8yHC+9qFad2mC0VgYK9gbhQAUylf6G0x251s3ju1o5N
mdixGwGyaZz4505kbVEDdTddhGcC6W0L+QunMABUygiNQskGYJpXAQ4/yIjbkyZb
TQ+5L3keDYrgNQbMxINRJEGwYP88jgHNMqf3zOGUEYyndW7nogWIYjLy8010qR92
p9p4S6T6FWqq/C5+x6ucqOwYjSjaBwf+Ga94MnTymK40UYrx3MrUV/iaWm1S+oNK
Mp0+71HAguc+fnx1QHpyEwK0LbrzoyVyrXgvUR6zOfMglsdZQ9UgqX4D3F8GFvq3
6nRbGH4WqERR+immVTepl7x+NE3pMAb2cvuQDZIWzfAanvaqkA/+8lYCx6+2KdV+
dzhCN7P6aP6C02cLUbw/523NOBtdm5eX2Bc7mvEi/v4BX2SBJzeL+Cg5hW+Thl4B
dU89o46nAbSulF2oRR9bVwtyW0rWHBj+yxF4zEEs5eCkhiOzVsqIZ7tz4VEIa80D
36aMxF4mNXemCjMNCyVUtLpE2Ogx9kvBfZAVgLJ+47yjwZv2TntXQtkpca1cBfCa
jNf9nsB/Eyto4L4My/LLS4IIl8krMv6jKtC+g5+S73a+EsorVBwH5OmYW9zI9hav
EVwQx0leKTgD6VgmXPG40tjVZ/EX7h78jqIcqexkyO5XQlMt8wKcFUjTfue4+Oh8
Sn/tMFycU3jGtfP9b9gHoHZlpPczQYSRkaQPVQNOwlhwDcBYVz7jr/ZPog9mxRrl
jsJKdai/oXdhE5vKWPI0QaIfd03A+Dwnw6zbdXtZNCEXuFCPRBHHHdk3O9CZtC4x
cx+eg3wqeFHEhggaPby62Bb2mHzwdF6XIqoatwRA+rEqi2YLEvQOTHSXncrM0Wmr
kX2NUfM+E6J8VtToPhq8yqj3OAukj+SRC3sJaX+VeTup+HCbZ1Az0DtyRfXeWoyI
b5zoFQRoP8a4hnB7uKSDWquyEPKtYvaj4VoEHjFAGzeWfEW4TLDmTYMbp7TcGM2J
kkxhFM7kBkMEDgphB38zStjVVQE3gnHzz211aJB94yTZzvGPq/mWsMCEkKcps4ax
FOHMrrWoonXjZuykyAnsPfRoTfnUkpsHuiLkNi1KFzAxIy6V4x1XL6QOTVpvciIA
s0qGhrkWcmFa1yUbkKSGwcxicRUV8r1gUyGYduy8RpCdpdo9PwALV7KWvFq+JFT5
o0jlOmk9UT6eob+oi9yOEK5N1OUKmryZWfFDCaOE1GCOnS0iXhxYQwRdD3SyDW5w
jOhJsy7yIqEHbCpC4elUI7xDraoplqF7XyzxML+WqAHbCtI5DSjHery1Ah0TmQPW
0rKxh3fflcpmK0cE2z3W5Efeydw7aswxAsXg4NCLsUEkPLpzZgoR5vhHi0hp/vtd
ewzRPvw/JjTZhVU9MGENixxzYBG21FJT6ySEVIYCfbMeHbcLuDiyJfthBGqJp84Y
PBRdKSMyorkuGdyeBYhGRq7QSKFTdqubrjzzIwPCkoLo3Dv1qpZliyL9MeRZ7wkU
RjtHZgWaw+88b0IZ+hJ8K1KXe1jRnCjDL0jhv0vlaZGnOwP7+vxKmNcwndMqvogF
kZ/QPED2eJhPFqWpY89FFY2+HimD1YoopLgecTongCujhQlmgZxFHChuM5MQiV+3
jz+cCn+I7CmYQvyY/oy5DSzMxIWfliTR6cOu6tF3A2wOluA0n+hO8CiJvX88kcmU
Mpv0k/q0Rb+vdQgt/+DcDY2pvvpjca5Dq9onr/RE9/Xcf+YSz0mwtGQ2GtQV8c0k
1/o+MDHOeG/Aen8tP8Ip7RAskAMotNT/DN2/gCFLBlA6ZG8+5Y874YWLj8yLrLVn
ld0kG++E7yklXv5dd1DziW4sVzDGJJqi1QiokWwtbRm37dwJoe3aMoBEknYbAv8A
kbcklGtBXt5zzJcAAiavx4coK72NQzH0aPp4nU/tzIEo2bFHtQLgiFb8ocDZcf6o
Rxy520K1N1I9/CWrJuiaH7xyv9v/fmyQZucZmA7GBwfOg+8z/jde5YXXu0eVG2Qj
bR+QMt/ZjYGAoWpEhZeNR3wIJfLkjNouu9qfw3P0GaySXt55tWmfy8BbvKk/UUkE
qa4kvUG6bfyLCQb57254ujd6Jiv6mk7PDhkT7HGsbyeUpdYMi5UK57XsfUcHmUoh
XWkTBEWO6FxkZfZ7PeXbrz+SQyUrif20cAq0VE0Ap7bDrAxHP3UEpruIWqU8090K
7YTT9iIP9NqFCjcwFUhWpY4COccT6cUoVuMgzFuZlKHmr23Zz+Db8O14qNCVhlgo
WLVkoeNol/VdHUEeUEXqWh5roNozLsFkBkFsoKfwebPd6IbiXeZRAFNVwsVkynXJ
y5Fp8jPpzuCtmuvigJBtw2BfkPI3fKfVoF8jfFNM4d6gOt9l+0f2qUxEORgXNJVN
V9SoR9uw+sDppN0GDiDUodNGQ245NUzn6c+bRzCvTLsp7FyuWPAVTGH3yV8WKrBg
46M9axs+GzroaeeMwobVQxD4xhSzJI7tSRR/P5YZvbHkeC9QYq4HI/d5z4rFE1fA
ZgB3VHMyoejviL3y0aZXtEMciRmV7uBdWpEM//OOyWamlMtJBfguLc0Wkc5W7mDL
iUFvfKU6GTZUQqAY6TOravNeY9U5ohELIuGboa01t10ykwUHWySVjSYZsFWr7I40
HvzqTD0RLhAjO2uTGVmWcsJO/sNYA5GvzCUNkrKVpKnF+FRAl12X6Rs40y5nWKU+
g44FwEcjyL1/eOlRA/iZJEzDKW0wzWXeydLYrqLFMJphVn+vuIrMvlL8a6L/SxVO
DSXjTwtZ98b/BptL2v6VafBiZnfGC7GtmsvfHdm2JNzM73GpQDpif+YRmBdalBZY
WZIQCvMP972ymKwhBtM1TdmftaG2YZNw3x0Wf2ZsN5BuOEt4CcSyQxOb1HkGtST6
D4HJ/k6/3BsGmuMhs/GA7+Dtuzu2t3oW7IiRrPc46NmTPwdMIgKsnMODpmmpF+d3
t6rO/esmhNtnLOgllczWOaayAkSjw7SnTVdlNdawpHxWtJaEIwXsramj2/NuS+dd
Ixu7FuLPCKoTEg8x45ZpeeYX20dz8EMDl2JvbVdcHhwcFA7Y6J/GC8U2OK5O0D+h
rtxaC0/HlgUcxNo24qAkIzqvM75WLs+dVqYsa/311w/u9X1rFVzZjJBjXKHmLKfb
PTZYcTQFyBNzr/oxgH1I2KjTl8VZA24FBKPccGLLO4nN0iDcH5rpCV5D2YUY4Ds+
rgun8IXDXFE2RnH/xwmfx7rrbLGKB2sGFUplsV5kNLpsfFz5PPlc30+HNVsxSHJ7
QCG5tXvqMN2+UutKCw1Xd8N36W70G72MTlUTbfvk3QiazIBj+XGrrqr4blARiUDi
woADpVOsuBYe/Q5u6sNW/wd96LigUbjPeEmjMJdlNESw4zlWbiafEnvkPWRPLT3v
SDflmirH4pxSlEeYg6cOHh35QbpZUM3QqM7moU3JT3L003nN2eLdizsIpjk39GVv
NyWc1uLX3wVxIIoybK12fmgIVIxL/UATz4DsEv3rHUc7frM3/daVwAeHbrEjcPNN
/8Gtf4bmVpQmifo9U4cGE+YsFdhefF8a8Nxy5EN/34+IDMtxjyEceGbHOglBv1u3
i2nJUZj/72mVcsM19osZskwXNDqQtAVJXTC98O4w9CbfzKv7hUaMSXRfFUfeVP2P
yuBZk7gLSzHVT9Q9eU+oYKqFLCunNK64NB4c9tx7hqLVwxcoFCAagAU8WftS5E91
n7XxbV8dGSyYLRu2XDiqHTvJEXyvN+u6p5utC+aj+2pN3WYzcWn6CJ9iofyxRECn
MepkwhLBrAqfnaHuc0/pIzjm5kwZwTOleZnqqHEWbc8Yelr9aPGdJbw2W1dbwyU7
voHKU6OwBu56T8hrY+D+YCEW8ZwVD+p/Gq2aBiZqXvA+ZWFCe3KoBJPBGiKeuml7
dMHyy9mgA2zJ0YqCSoRb+U1hwvDQhDcNEqbaQaaUGqf4rxbv60tP+NyR1euqOfSw
7mNxEzcgNeamCxxvG4g3mbwMonsU2+ZcsXF7rpE33RbZKszt4TRiO6BFaLDPXETy
wq4pQhkzACp4bWaIelX65Z/bRSYUOfWJAppEEVRQc8VpDrG5gHUyZoQ2kyq7Qctb
WZn/lD08oGA3FxboPfY/lCRxLSHNb9HKhlvxPlRdRtXeFM7HV4z7X8JAVTNLoh4s
POejcYDpEmh+G327VIyWXk2cjcub47C8XbvvKpgOFFIRQ0JnGAu49IPRekBQVm/R
RpY6e4B6t1g+rh4PeHv5QWcUdz4skahqSvthdCKHli5yd1yY7aF8/vtdN9a4hcry
0OZJ8bPq3kFEtMurJHU1HAL2mOSSRzanzqpPvPggcg5JtNfK8kaFXjdjVeJahd3J
zaxGKSuIwMkJqo8LD4iXHLbpNx1jAjRudFAkS6tpgUtyLZFQpkgKWsvEmY9oNaQs
diU9fABaDE1K3rLYR86dOmU5VhEEjjY2XPts+zH4cCLn1zVti6spXBLTO20wh+5M
13W9D38vfkvcL6UIrXMKHsfe09lZXM+Ywg0xlWH3rXz51ZmDE2eiDn9AdI88/fZL
/zoUUJEg8d+ggAsJuRE6z6Qyt0NNL1IcKbTmks4v5tCzb8m/vAHTZ16Z54tLACPS
4nVpGH0u75DvnoW95C5Lr3yGby8cYUoxDJwBnHm6+K+DdPbD8H1SmC3bnB3Svq1g
obXrmLHxUtyvfuK0/XciVN1kIo77hmLGfeOcBHqPQmgOR2HkjIGGII6OZzIJJ4I+
LPgl/sUhfAu82QYzgyhcRyLGQqr6PQ6GypIrOUxj8Y8GtT7pUxI2lllbAWlcSNR2
I0ZK9NtU7XO2ONpaGFx+/XK2v8fuUE0Cp/m484djCJWa8iSOuhK50g+GtWOK0wqR
7r8zKMc3jo+MMJ81rLfQj8IUffZNMhlsMUmo/uu8bPEJiq9K/mI8cDwjf6B3gfEm
7f74UVdzAgbjkgxSJEazi5BfsNu31IQ3ytI+sOxLBkNKXfGaNzdUVvcp2JGfiJDy
sp3dRuJJdhOjEwd1jYGRmT4nVAfImVIL2Z1zfXpFMRH7ZmXFO2/yRzYqznnPHSxG
pqo/kOnjAdhCFKroOb/A0BvnOhiLXTUh+9MuN1j3HzhQIX7/EPKcbXazRMQowUgb
9RVNlnVUeLqVRpHrJVkL8G3fYMBWMdiLhjUSdMi8pj6a614UCkaY4UwRdiYmk5Yu
bgzr3qiiUM8mOKhzuVjsWhbC1Sbmwhl46v2r+cn1AQ4cQd2xlcRo43+hXr3Fog1W
bXWSy68ADRjiR5vIEQeb9/CxFvdi1w6q35hU4VQbaDXr990ArD76lLl8M/kyVBic
OX4pN2JaBN2HASp2LMrHdNzJOLTAMYVCfntG+aUZl/51jpLTdHxbAdkbbT2k5W8P
8NPg1F9EFhJTwobedRfSQaaEoODoDYRH9jyd/E+2YZG6IV+yJcaGX2y6HIEbSYit
kceHNsRb3nmEa0ebblNC5Mud2fh7Id5YIf1/nNW7DlbMFc7/Y0nIlLNw7zEAF+pF
/ekwORA6reQhA8gngEFBDDSHHvy0QIb0GUa3Kd828WMjcPS6WwVp7fI5KUifVEZq
JZI0Hc/fKcy7OIXtknunAhDhpGafQmbnFiY1eH/w6PB7yq/IZ02kzHJqUfNbXSd7
UJhRRvu4N3IoR43d9MhBp+Mn8awqxtQP+JLTRVajnOBZ0r3pKyMpFftBlxdHraXx
0uO2xDvyNYIVdOcFddA5NVMRt1Xur1vDH1OTGeabK/s6nL+7pISbehAZJNant8/i
zOKz57ut88viBI+3hknXmSe6Cme+kOBPKG7tSWoLcfZbpHfFnmdMwwYOVdj0tOSO
UFl7k+INgV+Y6WQMD9sBaTpjC0lZiszFoHI8cTXS8PDUTBfS7Y+s7QwYY5X+kpqy
uDAi3ZUfAFIA1aEJFibkyVItqtoAh7+vqgjSV/a1stSLorNC/DysbJHs0RQKIBNI
QbaZTC4L/Ezzfl9e5uj9WfAIxOgl3tH2anxm0bg5RyEVtkSHkhyADn1jNlve4kXG
/h4bV0urrFv/ozv94SyOFtGRupAQg96oa3fE7LASTWSv3mYVeZHi1QR6zMRpev9u
V28bbARVRS6t0ev0mP2cCJEDB2drozT4iSXhspkBN+Q2c/9RvU/vET3kbpoXNyrj
vzffOV0lHEx24vukoiGME/xNDOJpgkjzRxkxn+Guu6vdPVskfLBClAsm0TaAUWv9
bALcLesd80KDHB7NbVA+/IhBh5+w4DrCepoSHNDNtpWxJVb8ifEUt3mUG8Puxq0t
+IUA/6iPbj6zzclwzTGkAwQkBJYOq/YQLgJoRymhRh4NQH+f/YnQStiiK7zxYrIt
cdDNwDcPZtL4LCy4xHCOeL90koUtSXqKh16xc29KcnS69/H6XbZR6DZVIgp0Biic
Li8a0OQFPwstdC29AMduTnTKG/N6wNuwlyjoM8/zH2Z2txTBsVPBrQF3TRf5r6Xi
3+fSnbwPdydiGKzWwRXH0mborL06tdg8MEP6b71fM7nn0C3X+eWCuJG1bbvORoP7
yEBu3jJX1/47TUObU1IcQpnV/mFxwo8+f+QDvL85FG9meaEKXPxX03guiVV+bFct
wC0d2UnniXLt7RsiBu5KlgC6p0K8MtnRm3pUp/F/vSRwN3F1MfjDPPs5xeTpuBOI
x45H8DHwjrto9gVlG3B5c7rcrFOsyyUmLVw3dd9uPuYI/sGQrS+DYW0iWLigTP/f
yBl0htA22aWKLyUG/lLmAhsnzyEKREQBOcK8uThFp9RCabsVq82mts7lTGzG18VF
l1KkAPInJBbIztW88SMHQ6yi0rG3dh22YrLfAoBU4xREIU7dUUiXnNDm2lOo8SHQ
uyNaIxvPcaeb0KS9JnBLYzYVKF5N+TsZ/SqZN7nL0cnnS3K2WbDBp5f6FqxcPdVm
SnDJVbNauHVkUFy+oBNrnTNDk6hjc9T7hTh9F+Jm1NUPZeP0DeCBG3IEkrloxMkQ
KWj0rtxvz3QMzZ11Vet61e7RC6Kxfd8RYdGqQV8omLvmYIHPYaXCX8VqeEZIAfbD
eY+u4+k+NErgUD2XnyX90I6m3P3iekiJaxnCkOmkDg9P9mbIvt0nkHWFEMDhW8wQ
VDoGns2B7zW8NoX05xAeJ3ikntpCS4x2iz9CJDefOp3LHtXfZ0sHVExQRRCM8fM6
SLLn8YvjhGJ0WJBLZrcgJPBX8qVVee5zYvVHBOosmlP7WPM258mx2JiilUsIdTNE
RO+7qKoVZdxp63rS5OiWkRFDNzOPCksU22PycN11VYahd5Plr8NFEpKAtLXTT3GC
fO93UvUo9XfYnHNVWeKHdyhpqFD4uuHVokLj34S7YBu/kSHrnixU0PrX6pK18iu3
D7RFHfuJHPpJUzvMqsyfvAb9/KuLGb6BofotXsHPVfPw5ZpI8SX6dseAQu+GM+Dq
jHQqscgTtRosYksxkVBo8BUlXmqKJacgR8NIT0b8LWDHhv6a7iBO5YXSOvMaLQjh
B3HNjcWMIRP9xRjcyKHsy18QVaN65/pMIGDUNWDYqIVnfeHyCXiEWnuDWzYXW9U4
Z6iQmYdju/Ob9WVArE9owtggAtmU5hLAyWFKN1trJ7Ily6Yp8lxsMWWio91PY+bl
j27htR9AHmqfifWnu9bxc9OszezL0072PAdyoUVM5Xa9NPErO6LEqaPMiOpbdph9
xsQJioiOfYO1tV3WmsH9U1WZ8qrV3nmhajKwfpHWgMO8fBBp5Jqg9W1Uj9DP8ZYm
P/dm7qdPzkwEx0UXMc53wI8KOPIdlo/AAcv3/K859LM1BgRgrEnukixoiRRg4oWN
sMR5NlUMVhQoHBySV0xbkd7nnIyvFwVYWsMz86L3ZF5piSbUep/DNsYwZzN7KKR3
NizXIUkBlV8GuYxAARpG76UxsNPki9OSPRL1sIoT2wXvpmImiTGcR/n/8grZPoZA
UtwksTorJxbYKT6ZCQgB0dRXKM15AczIXZzCzuCPwzHGMkmsbSNchN4s4M3jDu7y
iEFkC4wTxah+RdgLK8tymd6gqgFz2s9xBXRzEqlvMM+6FvSdd9e69L7DRaP0CUlh
+fJ3xGTvySbMMIBXJvnub7Q2Nbi41c5nxs7x6XpxBeVwb6CcZKDTZOIXoGeecBhM
xQ9jxKRfVtv3nh8m9slJmWQvFUDlZWgvxoSyeWbBEhJ96mqq5DLnMm/twc2hel72
D9GIPC+RUJ+bDMn2E24L0uL1wXUkV+xZENpx6NMQR9QDhp/Hqhc2VD97A/qUn+od
CLphiXrvP0Qy7HhFFGGW7uRBICNQOgoVZOCAb2cDD3ZxRfgHDBLoewlxo2fTcwo9
RW9+l+VkPVhLdFIj/TO/xYbsGV3uJEWjSmOLk5IxPrRu20NT04jG4wGBHavXKjIU
Eugh4zL6lbRsoiVztPLKpz25JADqqSjo+u2eZU7sbbJoGgzZC5cbhDD58TM9BwDn
zr4Mkw+Q+Dcl3U/KFQzmipEL2MXvDWRqm1jyX+th9LsofEhgRIYCOkU5z5PNpdZw
WTkM9mgzfL2boviekDWywNqQWAc7m6BrS7NqbNC36tnozlWWHpFtGy/+KaCPf05e
6PfUYa0IFrcwMTep4rmtME0erJhHJ3FTTYafwxRTVPuJaDfl/ZpC9Vw7Nwm7ux/J
ZNVY7sYMKHz404PArYMmcs9gnoiK6G8IpA5xufcYw9/1RVks/F78032Toar0+ff5
boaM8hpeJTuy0q5YSqnAlj1SxP4hsWh7dvVhnKWo3OOxMDwSr3U8Kjnd7Xi26EV6
LA0+x4HNjY5wX5B5iGiKFbCxxpVcWNFVPOSf525jP2gqWD5KlfzJMpfu+ZehS0KK
plpPVolZrHr8bB+O6Fvuaop1I+3qpaF8CZtkdYuv2ygpHwu/DN65wpH5c7mzXkId
2U4j0lHLscX27hhKx1Gissxxm7o1tE4WSfHvD81u048Cs1WFvPWbFphjJ061SIAQ
SBys6XR3y3FXxi0hQxTuXJ7XWYj9th6+FGTBTdLfY3CnL/L/O9YnvzrK58rQLRRl
taER1NFmSywrLrUU4VoyjELJbQw6e/PGlqyKU/9bbDGop6jMwMB9IZB3NfIkh60i
c2o81HjBlQbXkMSWWhTPD+mkt0pUv0tIWXhZiTh7IgBKHnX/4MFJ6f/lKXEGgxI4
TtqMcQD54xtkc00SIUpoUK0a3hD7x3Ereobr4ic2XJ61um9Ydad56Yec9/Cq33rq
vi7pePSs9RX6nNb8mqxR7SKnKdRpi6uYWsimtoAZT3HQB5EZvZNZyRGnW0adB7Ca
FgkJInaz17asxm7pWE981pYF1AiBosPIENJqnddm1JEHZJSTwDU2akgZOyY8kSjD
8BG1M+ngclFuaPIisM+/1uKoN4YRZkTc8kRPs+xHo9bE/75Nj9Aoom638cLP5QFK
C1cljCSZrYMryLA/ZBlH3XdSNc+SsKk6NYl3J+BE3D5MoYu2J/JwOG4Ib10zuwrp
OuBvVrvh+3sOYM+9NL5/VoSrx/GMm7Uxfyy4gKo+GAzQTWvcecWfGpOFjY+qGAXj
j4gN9ThAAyRuCEZ1EoG6TqumcvFqZ7U7URfh4BTLgAKNFDmbOrnxpNY3aOxQG00N
jgAMz5KFJYIMGzG3nn42Tct5YEELAguwSFnqXWznWCkfwNVVlH5q8LLuphAfTaQe
02UJuWzJ/br9Lw8c7h00tHC93C8AwC4C37ZH72JcH61q8OUWJcEnzHS51p9QJjqL
oWp8IlZAOYU6rn56gqtMlPPr4EbuoauecIGzEGU8jGEUkTtfp8X54I9hH3Ivo8Pu
NNCgoNQHTMLmUUe36LguGSuKaZaCSBtEHpQBAQXBfHpzM3HEXuPukVv5GTkgWS4l
FvyARiGz7e2oTphf8YFKguu703wfpsxPvch/fDpM8pg2LCLmgQU0CYRbwVZiJZ1X
X7iimdKlinErmlqbzQL2nR/nBTCcBRokmioeSFDk4hiEdU1VIg7bS9a1BEI0vq5K
G2PABKSS5ip/3/6orEQT1fx3MBr30cw4z6myyE+p2A+hW/7QxoU6oxC0XV+QyL0m
4Xx0QMPV1b6hSu85HUbzYaHLVOaPIJD9bVoGdn3CKED6fIknk1m8gK4wXnHoaRsR
dJcwC4yuB0f2Bw/qn41S+qmshdMJYKRWZ7CWRRnMga0mTee/7JB3qANc2OgXWEDY
WPFt8FXotiLWzTYN4CmV6eYXm71I/OI3aYSdIkVcSel9P/gnAtGxPAPJI4sk+D/v
Nq/JbOUjwErWM1GIHwskhB6IMGbOqHuOJobjGDSpk/+OyZHZ94hButuPiUfkQL2n
XWCV5nDWh+NuhsPOOnCzVPOlIn27xv3KMMh0WkX5le2TbRN+wIwQVTVTcmnFOR3n
/ArJzuVvrGA9/43AL6L0L3rDrf6zXSodVErwRuDExxHI7pn/I9mVMVSqsB0X3CvS
elIJF8Mhr+fuSdUfGlEfxdPIDEe+qEPpo16+fbWpax4nkAe1QcamIRj8q+yAvcDV
QZQT+84TiFuegqr/csQXLtJJk7gzJmbH8C4vDMlzZs57LHNZFyOaV6NOjY40Qh1E
R9Sn3+yzsibxPltY0GnI8n9JdeaojAiCAULrgUJTQB0KRN37r6WptYIEB5M5nglu
uYtpGVj3DGirBxAb8fVQjmqYFb84Pvgu4wJntGlh5uXt0NLnnoRwwB9KIiC5rjwC
Omk28IAjeBLFcb5p2F7mYHpDIR8USqI2WwJJtQLu5ceR9BAoz+i9MicwLTVx1bCt
wLdDwSQbC9xIVGU0kyGWMY0zhWcavaFht9PhGgTHxh0A21C5fI1Wzqfysx3ExUPb
NacKcvyjEgfsiFyAki3AKK4o1nyrsaxpTj/Y6W2XUaca5h6D4K8wk6MXq2B6wv0o
DFm2wyyocHWZExCHmNasHoBL85Gw0VgDE/y5sR/MQfD3/fd+zCm+UVh+MwYMncHw
xjcxak9aUqxblJ3OL8VPzPyQmtZ2kryLX3ScBDG1PnJvFcP/PPXfL5eawniuEkjO
nP/NqW8zjCBtvA5H3MuMBVHFUeeRkneNv+W+X6D4O3d6fp/9JIlq8JLRlg3HsPOU
uVbdWSut8zzyOIKjhgBSFV7JCbjHsIaKmYzWjaN9ibzrZ5q5j5MDVJo0z73EuheF
yCrfa1THE/peF7wTTAbztvzYdu3avZzXKxjCvN6I1IiqfPo3k4A4ZA2Qv9pJYUKU
4Sl6S/xAG95dzp/YcMq/SbB5431LBbzex+IMbxEDWidLDuRWCCoRA9ofmp+pYQNa
IU3oIxIjn44PbIWhR3Nqn2B+VSea3+j0DHgAcRXFmJEKVAnIlHSvtfWLEH6D6U1x
XcngHtYGgFU/SHIMCo5mCU4J5aLNZrDD2ScNxm5bhrwyQdYA3Sy9kzszWmG3cuSN
dkNwfIg6MSwv3tinjqAQhTxEPXxqiiccnHexIwlvHpjqELhgaLlGPnjx+bFEIBwG
66ASvCV3FzfzFkGGi04WckhufbFAmftrPMiXQ+0EXJ0SuxlfY6VE4xzio6LUTQOk
z0v38ZiQMoQvVazKgHBq3XH581Wo5iok96dYofZi36/7wuFbSfu7XCX8Sf+s+BHo
2YmEuOiYMsENhoxT1q5WyD3AWRgxLT0/T5Wi45m/+xg1GAPg5O/978iWY9ZC0eqp
ZvsdvvXoUj0m5dHwl2iDfkQmbUjKcUV4Nv9/TkbbJSpE6gHNg2mK384nisrwJzq9
v6mrya1ADyCLJVg5IhvIO5zgOSyNIQ5EXUocnVu6ta/rT1Ae5ilKAp90h/aZrQS9
Hmc2hF9gitQ91qhLbWVhmIbjiidIB4elREBJkY8VuH2eLki6yr9Uyu8tJdsC7H10
168HjeOWAZIroaRCZxHakeZ96hyeOmiiixuKR4yok5MQz3LdU+3yK7deGfNvTtwE
dXruHzD5cUMBEkG9i/iwcl8/jH3GgXuhSpL+UDkf5j8EwUSrGbxPlTaBQyrWV4Nb
RwemxdVFDAtyld9BwTw0oAWYkv6sH0UjurU1zYDCIS6FqSwd72T80/oFnvOTm0/6
/4PBNFOykUeNdBfG3pis7mfYPzav+DqdzBW7R9HuCYhLih3cYIQOoiLAZLERUs47
det+xF3GeteCiOqu4oElW7TaCkROqt9PXI55wCywzKFaSazMwRZfR2OUTrcYYlUg
VydiDweJXRJ1bpQ3GCzWV3tetWaSM62O3Mh2uDFlRRM3f0mWyVJyWjhCUgygOJak
IS8gaayxf+UnG0Qw1MmyX41koFUuwMz1isooOkaEy99fFCdvSZiTH0BqmTL36v/p
g0RGvom7oT2YPM84WvaoQzYZxGrS6LKMOiE3suUYJPHZwo3OMWHSkq/H3FWKoxKY
2xUGKCvKk9cK+l1V5LsTjH0q8LZcx/+8VyK4b7Z6ClBidGeJBzwmC8LBIIr8Hx3C
d7om61PA9aoIo5CSh4DlYLxnhkMFIjPn9N0N+paLQd6Tw9yV5VNcBO7j3k2nxlr8
/pqGm9T2bAbzJlbq5E4SL5wqFEN2KbpGjv8zbTWklOGUJyzOvq7zCip7wi19mC1J
3NqyAJtAyoSNQlRbIo++uJGGJnTeSKdcHpDVY/aT/uLSZ7dIVIGAbF+YO6xg4QaA
AJW0BhUWUTSKShRe0VroyHegaSDhIiUHawyVNzJdUf+GtfRH41j5OylMidKWhSXI
LU7RiOknvM0yC8CI1cUQ9etqjsxHxFPEsnR+OyADQBeAkj1lqUlQKkxQecCCiqhm
agTXC6U/h1O4lV10azY2IXYWTPhQSnFk0wXTxykPb97ypEiRCO0WEP5lfJieTjPt
sqJi6Xhx/nIriJ/FT7FnMMjwQdaaoDSdVO8n8frkdvbWHzdSScJpVV8ui6BV5Sd7
aOvMiwkykN/8fkAOKATJuZMORbsQoFacPkIbpjikuS7VkdzwUC6q28dwMkjzWdEC
VxFxEWPn2HEt6M7qEW0HmOMnp6NEl4MW6fS4mziCBCvj7eLXE6z2G4fEznCeKU2z
r1LEYf6WdA6Khuw3BzDH25NLuN7Q6Sy3YFZ1DidC4eyYDEN4E+UQ7TfUhMsyMw37
AbhPFkdbfP2ZnE/q0tgmWgp5vQ+P24XgUtI5ukUFMr+KGlNUkMgSmZ6bYYdvI5XO
a1wQ/ollA99VPePjYwNQ5BJ3ro3ybdP0+XFxTzacInWDwZBtfxykdop/2DtJJSHQ
5YbV4n3QUoL2+Gh+nb7un9f5cn+qDPlpiwwoQv2rnNBSuPx7FISHs2y4LHFIEtzy
q513B65whZ3T11GFcA3bwhx+CKsJqMZr0sD7pLnwPKHIl8KlQLXsqR+wj6S48usS
yiGuLQPkLGtO3JLR8Za2RKbr3+8KBkiLG1qPK007LFxP07DX9NxLivQgd04x2blx
zYgIOiIeZX514+pxSIQhG8rt9w7WPLabtTBVsn6kNsG6QxigpmwGLj0p5gn0/8T7
2jTw0eytpXQSFDXO3jJuO2FaRy/s9p1WbG6m9+XCYvgqOb0gU2LTJ93GDxlq3dbo
Ue42Yr0dbCYTAHqDr3sCosgF7VctF/nvfqpwjTEjewZLuq+K3TdBPkeaw+qcFNdI
uhH0Zu1L1euRltEjBNiJdLermMn0CTC6SakOoZYES0/mzSZqyES2e4zOPnPrLx5M
Wj0nrAj8wyqsLRlyocJ1qwaBhbrd0t97CFqez28UR7nyCGLuiGXtQGulQVAmgN7g
HZGOY1G5pbzqme9bbgPXnpFHxwg17gmGEioa70aW7o0nL+v1m/2a/Gv1lDalmPgS
1TJNT8Ye1qrmJFi1sSLplbxNM2T8bfyT35I6HtNKyGu8v50jP+0FMwF6FNovFJCf
0EfXsixahYNJo/xOOY8BUJYuGXNp3EZUTeS8M2qCHdT3xdQyw0QUECOPR1j9Rvoj
eCkNKlPOnEqqZUbhQjfZLsWPq//U1HbKAh8PZl4/KAIDYzurx8x7BouJ0gB9lBSi
fW0OC2wGpZhF6U5qhCgN3FjzGAKa+MSCiuRjp/dCd77gi4vvhl5UjgoE9RcEXViy
1r5B2OOpV80wMrLSgR9idExRpBPW0PhTSgpFZl6iNiMPzqz64p1c1CksQ7vDyGo8
265EvswnruG5wHr87GgQFdM5mZBINOUQebWxRyFvGyzEKRYLZdA4Cr4hxPXvBgv4
6lCjY3SkExa1eq7vRX1uTlqv4HSwRdQ4ZOMmhgWCkJsUZ4sF9cYyxlGoQMe5wFY4
jPfK0pm0rCAsl74FF7KCUcQFcmLMtPUpMdfpJOZwWVwPJz0cjCQdjh4QqfVWupSj
u/Bp11F3V6C3cLoyp+6q/Fu+CfVvoyeTivgzQ5dyUVz3aL6V/XRgcuZEKOozi3/T
DCxM3WLP32posHPB9lCOFDxFSiq71wWcohDBpLzg8aJLPWoQFr1XllAzLFhf3vXD
efKWoTNWkm7CBpvR+6oaY1//ZoKjOjq0cWaYMErL19Y44o45fwi5pOARwizp6u0H
eF1XP9Bi5AIA6hF+LE4Q8GUrf1GtWwg31w2U9nsy1kfliu0mca+wXdZO/2HJFT64
kIQoPJrqr21VBCEKkhh03/TRMEOPUVUlrtr4ApOg+Jy6aH08eVjJhsMIh8tTJOyl
sI9V1iy/vzAsZeCRELbXrBc0/SPFjvo8h0ilk62m+XhU9/Yq8C2+wq6Kcedt4kut
OOkv41okJdNhePssNwHj4sXXmAnPjf7i4uRcMhuzcCtPM/7iHM13298PFsP+WrKQ
jZ6Wsd1a5FSl9KAUoieDDKRVYaKdJYO8qnkekwF6KvS2zW+DvDjgRTW6xekQ5XoY
a62Ge5ZO9AW7KBPEuaoL+e6ZGDuaoX+zE00zbtVflgM5w4UryfO1R31zMZZEV7th
bS+ncbXL7kXPwasOwxJbc7/bIedq7GPXL/4E2wpNqeMxAj5JtW541V07FRyE9b21
Tb2UzMzPwZyxK9/62Xi7vDSxCl0bvzVsxK5DR7/msaxRt7duw0iEIUF81k4Cx4PW
S6hQqtP5rf2VpI3Vl50wRctu/5zBiMWxydJjpSLnjP5/zem/tYIW9JhrQ2RA/iBp
GaqU0bPkn3Mo9LPFn/1rapPLcmAaGtn80g7N0X6rALXzue9Xrh5nMV8F7FZT0h3u
Oqr/I5JaLCWbGEHKocPHryKEzB2UP0IQ7MgGOxUS76RGJ+w5zmzGhMzwIEk6jjyE
H+V2UGISVTLvUyGvh4cvyPInSXJZ1AqPZiazFK4ugq4/vwW9TkLRc6Fis6EBOHaF
VRvFWyrBAHF4yw4nc9ELD9MZay6y5u+GfBMUrW6f3ZDgtSYVOLULsPiwSZGj+YLz
ahyQdimy9RFE7JglDEzsWg22GHGEn2m7ODW+4NXwXm4Dw5virGCNlKsOfPmsUF7/
P1BONXhL7Psi2Q4YQNBvU7F0m84SUXdrEzBonS+pMRzpq+P01RWdSTJkL+93dnlG
FYLUrp/WD0Yab1AkqKp596D1LcXed0KbsvvQbBah7r+RRXrArlnJSOhpv/dgGBvT
HymOQ5Fp6J78eaKKCCbsjM3YGm3RaQT17vA+hVB/hopSMgf7jyIVh6jUUiw98OYm
PVWSjVL0CROmt6lctI8XIFV9W80FXx3NLPqtzWPEvgTRDKDqPWh9NX17gaSaxGNM
FcqBxu424tQMpeqWPjEr3EazbxaZlKFWqn7SiPNqn163h+y5KXMJSBr17UKH8xW1
I+VYYsnGjB6fHkGeZgfLQm9KwCYggprn5kGEBfB/rnADazBhQe+WV5xLIuxo8f6I
Brl2586SqYf2XtgKK6/5no+PbzS1IvFSKZdVRD3obuCNDF65Y5a1kN4CLw+uLyYU
iOOEPxLJVwOnO4G7M0gZI/XALOpKGFVvSpbZ2qHO3TaR+8evFrSKpbDAcEkkOCY2
GniVs4b5QJFsJOOcneSVwJK+3+I6lnM9tTepxGQmzYtULqJK/oAtYGVRROFKdWnb
K+Mx0heyS/GOCM7ATvtY6alVuQb3u82ZopbQqfPCSjP98UeMZGCeBl8D2LYfVIXr
y6V4EH5gEk3AV7NArnFFWvxrotL71PF2khpDB3YQNM47LnUbFJFDVH646CjMbD+t
SkD943y8dc/PRcKv4JJIwjl8tdKgDjfGq2DlIPDWpmrz9AZDC3psK/q80Samg/L4
lKbvAcwKZa6l9lessRqSQJNEPXL9lTBWgf2wE8JcSb4J4JIcYhieajAsFpocxBtR
BswLPX8eLCzqprds6a6tUwcgmHW46+2fbrFF6HdXT60TKi6GKO7rrI0mvYo/92FC
M/TUbYwYUSaiicQUaLYGF5K3FfP4rxOA6quMOUPM0UNQupuy1ljpjbEvO5KAK/E3
C8701nb/ZXvO+6HWsrOWM0KCDdDzH2MAUKGTqQJCcRuxfoQetFL8J01d9oZx7HFr
Yaai5TUak9r+PmTy2ivUuiA8uU8xxAL+eC/fJkc9lcluyghEuuRpxZJWzQ7uMzvZ
Lj7+a54K+4B9sc0lvLg+uBEoHJTcPCxugfqptFJTNz3flpWJvccWn3IhvgQzePPQ
yGz7BimUz4n5D23Bv9IMedTpm5iGICgNciULOngo8ftXFm3aWhhF0vqn09fQvlXZ
oNfl6n0lXnnoOq3S2ZAOCXQKbFF+YVu64ez0oVJTvZ/DIxs9zCCV/5fiSoESX2js
2wbs/NX98F5PNrn1+gnIoyE/31TZI4S8Rw0jzriLHVQzaLsDh6SZzY6vsqWK0OnY
MLHAdlX9B+1zd5hMdRm95JKazwp1fSFalB00wsXmILMbga8PY9BGTeAWnwU+9UVA
mtGLBHs1YJLZelW8a+EjYqp1Xzt//lT7DFkeka3rn5yWAvaE5sSjJmuboGD5apK1
AnZFiEs9qvVLnphL0x4yAlE4U/SUGlCLoLAo11ZjD/HNZm4UNsxM+BN4yv9/pOF9
V09mTOeav6alSDng71AvoA2/nYEciFGqKkEkLCDxLAHIxWQgnl1rVSK7bAQslB2f
si6BU/4axSnCE2pyadt7ppUpPH5t0Fn1jxS6ZWXihAc8rotCCU6BBpVtP4hAQRwG
P4TIve4R02sb5FBXv59xlz7/cqeql7PMzdNbEDkL8k1LIGl0kqcYvL+ATyIAz3Ct
+h5ydvjdClqYUf92a9gQg2UnsbH2d+yMQC2w1fGAxsvpO7CAcF/e0FWWv9iUzmC+
um0yCPP/coSsODoTKlvV4Igui5fyD9a4ybVd7OmzRaGZ4Zx3hEkWGANwUccbJv8x
7JG2um2IHOiT8YYZCSpHdJteNzam6tEH92stAw5lgUIi72E/5xwrhnsR+7v3Rfqm
KuXCtgzZs7p5tKtyY5IDof70au308MU6kBRz7b52kD1edel1gPET5iwGoBUlwOC/
CzmVv2e0AacT4+ExulLI3K/qKaKzTUVVhAD6yBjEJda/RzlcUSsZoLCTI2p0d9X5
3RkGZSxIkDHsjc+paekEqC6ftMzCGw696qH1QnuWdevSvMr6QfQHWdvwXKe3H7uu
y0sZHGFWp/ZlbNBOvRvdHXCAtfTpzJe+V9abe13SeWfrChnJtzyqts9WaLaK1eGS
Da3FdjnU/q4wqFD93Ly2boq9ytILQUfBsHfHfQ2XONc522KfWT5RRGT/GZqzOme6
1UNfieorkUwIR9WDFlooWPz1iMm+oyF8GiBLzcMFwxV+s+FZCwSaSRk3qHBXh2j2
7zwjiwO2wEu8PlXODV1B4hcUtdm/hhmyHEhcfvOTG+Gqprlzn04sLTegsVK0Ci+P
MVc9jAuZSXtK6dgWLOMUuvvPtaCDFvzIWhzyo2/Zk9jYU8L0m1Zpu3LObUMKQjYu
6sad8dwivP0W8Rd+XtldrlQ/eZUox5HI5KuW0TGda7rftgDquoGkFXOKdIFyHgfZ
cAURh6IrZGYdGz3/Rx/cv5+eRraYDGoSgfwn3hVao83kiy0L7VNrjgfn1ykB09vR
O88U33rPj8YM7zBhBhHNwlQeGVithfvq7bIdp1YcGUYKlCWTnSvCo1VJhKg5f8kK
0DDLO5gUd6gXMK3Yldkvhu0Cr8YSj+EoSrS35zgWWrrVZLciUSiXRhAXbFfTbYRP
3hECWRk6waoU0wp1H8J+yOGUGicU8jMbyH7DfznKOR2EB/9vSH0e/OomewJPIYfw
N92ldqtn9Wgkz9EaYSEUxzabpbKZugZvJRkJ0EJhrBU5yh8yNxcXlPiNWqse//pu
RZX1HLNvr/Mbuv4P1SKBBrSIlKh+5Y0pyAoP2Sq5BOmrwLWdwdUKLxSR2qKs0x3g
P1Ff66jj3+a3JXUXRiAkVeLvx32zVA8ShnzLV+bvYsWflTjoPdxo9bI1b3+a2pTH
1YvLtNL5R9JOb2w73C1e9cRYNNh46ha+L2u9w50HfSn3ocfnQzfZzwvEkjGmUyY0
vJTMVdp1GZb5fpSwNlXSNsMnnKkB73EYqaie9itktFJVs/0CpKDKpM0WYxYfKTtA
MXED+ZfYMS7R9nWeXoGx8/erH6jKMaYKfyNFiF3pttxNOWpD+T37wW7o9QwSqBiE
rv2LbOxCgsVEQSrp5gRXRv5mc5zwsTlmekzX6GaK8DbRGkFcfUJoikb39RbiKRl+
LHH+9qaJZ9pTGSWL/KuayWCV+OIa8nL97pGQVao/wg9dhRguImuyYY9rARx0gDKY
eW46pswslB3pwaTCvcS0oLqpanVmoJ+UoGSRbRpmREq3KRIidqe0ugXgBWF5vpog
7Eiqqsfc1enYt0Fz1dMoJQBbKSTGL7xGYWWe7YGZCv1hUoxumeAsKubMzFHyqVHi
5h24TkjHBxcD5F4U5CnoGtyQoTzM1KLqV9/CNt42RJa8ipRBjTjNy7MgjWa5wPXr
qBaA+nfdAY8JoH23kOfNNz8ZalgQWtBsfy8lvXU/HKfP8mqppajukfk7GOn2f/2M
2rx9PD9iPMAt+cNG3vDHdTUxaVwFIqXA9zGmN17+YqhBbeQYqShllFi9UBRi02Vy
2B3JyDnUACNPH0JLxAkyr5EMfTt/EoZf+uxGXlNiqItpvzC7qXYjKGYpVUWhvvHT
ZiMGmR6wV1lg29cJC0ChXUH3a1bB/A2efduCC0k3QSuQHyU69z9rTq5jHXIksLiP
Bma8j/JzrIh0THy+vtatsZ4jwrLunU/WGEABYgWnVspfTjr2Yhxjgd/uGGCQ+YOh
CwmfZ0Nmg8BdvxxItA7PzG5dLio/2QO8Dw1wyoWFwlbjWDyohcxmQYEKOkw0N4cN
oHsJ0AaxV2C6LmsLk6LW8K+C3MPUUQiSZWKY27NHpMTOZG61zZsd0LkW/RXpOu7R
G6nnjGPaMalejWt7x5doTaw5wvW9s3YgOca8rXdmFS2mDUqxiiOLr2e2+CE2uSl5
JWZMT96MfqSpi/rjutU8WKSoiVgQUFT0bRiF88iVn4KjiFa0N5Sc9Gv2IXa2h4KU
j//KffaQZL5191lI5R84x6xD41hQeJQreDI4OGUNV0kbCZoWlwMSlcAEXwt6oUxj
31CUA6ByrSIT3MmgSrfWzrYytlxpEvvmSQBgLQ4JDVtQ+EFsIsu/wZ8JGBwjrBvc
Gfocqfj9pnL4LofBeCCRsVugnLENaQ6XKtS51KYle69JqyZ5mzqwdr77L73MhNt6
AjRMTe4OItXm9JRsx46RxUCxidusSrqG2RIoMRe1S1p4CoPDx9eTGbHhWNyRMdOs
GJFDmUS38Jkr/5ayNtj2UdgTtHvf0Xk0dAnrLJXf1QFyV0115GtCurtXn9sUswtI
QNCq6v3OvCRPFg+6Q2IjtobV++cSTnqky88pA5XpzCXcvPuiMJJ0QD5nHRiv8/G0
99SEHaEO0KE1HY6mTI6Roj14Ci7tKt7VBorxLvoEtDsnMYSeKurK6J/nnowpmI9d
dUw5pVIUGieYjKPJEQRKu/U4Omi33Lx4LruaHYldLOTjrFbkNqRGOBOtHG74Nyes
0D6uXGrlnySyHjbKtVDCrYk+gJb4TYgPQQcmpTV+CVzbj6tkmtwJUSyTifxa3oCa
BwZbI+QWzA/kEbllaAPeO48r5+Th8asAiUJxIi5YSSaYFfOQatTSxEwfCD657UL0
FEV+NM1Z3GHxdBtijW592PffYf2DONKhmBXNoRGzCLRKGGXTyzLHIznetVyh8k4I
A54B3BfPSULhoasEEC1uzAKZLzPUpE6c+M1byCfexvIiN0Aaz8k5J6MrnyhSc327
w7d6Xm5gJni+vWeGdaPuA2Zux5KtCnwW2h3oCjnHdhkYuFivnrPsI2daaS0iAPt5
lGeXh5BY2R+0+9xR4Cv8Mu0nDV9kC1KEoYt1CuyeZJefMcfsT3u+tmnFt3YcUwLb
HoY6e6luzNuTjwDXVyWRWxd7DgQBqqaD2iDUdVBK+ygdbtqP4W/xbVoqyfjtQVRb
4Ftd9c9oZwBfr2E4pqB7ho3YSDLzS4P/S206wnxF2e/9GBaL1u1xjsyk7vHJiPFk
O34t7G2zo3h5lJZ9erTqUeTAqd0gsDeGNamnLUmmoy0DV2tuCWFDKdJKlfFLWaqL
6phwzpY543lpJVLV3MPhJ40wY7wJWClkAMNbPTOhfku0ea+E7zC8JhzBcpeOesko
f1xDOrLD/WqJ2dlH2BVQD2FRV7wI1q+rtQQXOOzU1BVlVmQXXKawRMrKGnrvZobl
+mjCiV2zb9SxvArsqc96a+nX4ct3x+pJY1F68e+jeeeL/2rInwZi5HYcXlFGygyb
8paaXvkBPbWKnzsMPCW2fXQ9GwI9NftTJ3riWyHkB4pPYPUjWZlW8a+wKSvK4XfS
s+Bst6a6WW4cBY2ka65b4AgsgRPx4nyqDPvmu7FNt679I0HIZnEhwZLhKLpqV12B
VyLkSM20f+AAPZC/zqVuzBFRcuBy5ZHftWntv8A4NIkOFGu7nPP0CxMvSpo1DkhJ
+Qin0lNUBc9XF4BWQoSwjP3p5e+o/k0Z+dtBU+rFIkHZ5iuXjfIyy5WEs+LnUfLS
sWwp6z+tfuYJYelpTZ6vHAIyoIPT6ZQccyws3tTCDt6nm8u1ZfsDa+W8h/NgbSwe
35rZ7wZFCfhWm7VE+RT70W467oneVKV4rXphCNP4o9KEpvw9Xrkj+tb2GHYmnQAF
nO7XvmokBiO1ykFfbOaFflob+kfO9FhJyJR0A9q38i/CXHN6F4aRCqzzsQc2INzx
VzX76lcBtwjeiLKKNX8TvU//0SQlWDLQ+npbuld/nGPyZq1JOBoLrforu5FqdGHX
uyGikWanTuT+gChMXG3cI+//d+t23+JkEUNrQcCIRhPdT9VTEq6ejLUPwLzl0IIa
4dA3te0eGp70bBo8yKCHCw+RLWKg7+Y1UkrgyHgqCWfDLfMfmEu1VZPa6zeT5QkQ
LTJEBCYU9CRF0Hz2tt/MYsKPBTxUfzRUUG25SyWlB92Iup12O/bV8dvCeeopWWxX
L9/UXDuPtj9iRIEL3vu5IFB2bG6n7opi8nbioGj8w5JOt5KktJjJzuDnrgOEJmJN
+k4e9u/KFM4p8V5AsCGdxl1PyiWP8JYSWuT9YJI9Q2S1QOzIhtpgqB/247zAR9bW
Y9ygjQpK+wI5Vj2/m2dxieVuTvotiRZmPamP7TL/JVmvvyzS03L3lmplo5qIXrPU
xVDsNR6bf7VarD9V6LRppgU4RTA4U7LRP9KSkLMugavBH54tDQxbIi4R3wMu3IoW
1MVQ65UmXqNoeRv8GDWgJ4vq+YHJOMq6GdDKboiNDuSpv5DOjkMJgGuXpYMewtyg
bQVRIiZrntSOlHD58i4w8IbQFm3k3JGgEOMr2AJg013pGf6hqZfFg0KN+q9eakXI
g1M9dQnbB4Pzs/JHUNlZQyaN5P2yNVzTCeeHTKUhj5J03JTBtGF+HjwKcVhO/OzV
M381N+gMqOvbojKMUX5iBn9pFwbJjnlYY8YC48bI5ZEJiH7zRS//85iQkhX8M5wL
hic/t317rbBADVPWNbGCuIs4MgR3xazWG3DxIw8hqCIBeieujE/wvOEmhovUeyv/
NJX4V2sqln3uCHSkFnA91UGrzz6B2cJiuiNSxnBVpcPysahlndZgP2XgrGjJf75Q
o9dL7TDfyqzspJ6+A/l3Gj99QvTcXlV9VKxQ9GxJDciFOFQngi7wxA5U6YQd3ejz
pfUwQB5YaHx5ho7ChzfcdIK+rJgxT6pdo22QThzx2Jzxf4p5/45jecLJSnedrGwW
ayXCXlFqEvukMTug+RToQe5Q6V7UkfIOTYSLZnDrqXnN6n6wwHZ1VgfJKOX+CjP0
H0cc8pTNJU6zC6dPa5EhVMjECGTyvDrKo5T+DO916ufOOKSt4QArC4L1cV4t0uNm
gSBB8viwS3VgUCpBBzh3JzSltP9OLqCWF148DfWlt2zyXsfubS3HlNnu9gN1nHRR
hNIB4bJA5tFXzJAg/RBAKer0MBH8mM39rNpV2JADzMm2dbyF6H9nZaU/ka3JOWO8
iNzJEJah6m4r+mf83XiQb49PYDMpk8T61SEIYU7rApAoI2MCFg0hN2U4DChUQCys
frsyyII/kE0XpgU+ZE1h9O3BIBvP6CS8yq5FOK4NlMtwEwtS89pHiwpR6lXcdlC0
FbctyRYuSHkbD44MKA8IuBrnQgBWrvDQ5zceIe2AY86D7k2AYhtbtd+vNYw0iVtb
J7AmyTpMMphIOcuWxeT9C3t+2AOIpkrDBlSNRZGui3RsCotevJ1qZX3498U6InD6
0ENFjOvbbhzysavgMBwnIFa8pD/5NHoXfMZdjiZv5PjRbBLgnM6ZfBpeSp+ctbEB
4xFnA/NAkZNMo9BvmVNz8aiiy5DiEQe6wuRw2HYutU2GyeYqCARDnndVzoeCO9NB
9KbUm4DtDn0MXWO9RMfP3Dstj3Cr0RL2NylEwvPVjIEeLRwJro0+u3vz2Jgdszy0
GJURbOivYXFW4+ci+HyX+0hmgdTdtu3EI5RF7Lpwvrj3PU8jMr5NxWSeNSawD/1t
PUrPij4QpXxPHQnwmzCSVNH4vIkrSJA9AwQZYwVBvNuMayv7CGgpdyyKT+MABt3/
E5CtUPqIL1eETNdfZXkellBude7oxGzUC8lXVwQzGQfaV+YcozgNBTJMPicq9T2V
VnbkQuR0qSYZ5UFifN00hDufjB7FhA/L69clmtplUHSyLy4NgCE7vrun4+PIh6WA
dgIOV7R/FR1VhedLH0Eygb1zcS70WUFcwRMj2OJrXKQ7SCJoTw3TzI/6ZL5Qf5Bm
uyey0Ftn91FdhkpkF62rN6zTSYZYPA7eG91pZ90uQlxo9KMNajIJcS0VnAlVfQSO
BG2knrB/kh5ze+Q5nojo56csivm/wHfiNIuZcjC/wfPqVKVyi25cThtPYPijQaDd
l7e2YliWOSbPLM/qoA05fXJQzTErF99B6HnHr9kN740XAEfAynsI4I1ZEcKN5MVp
3s1d3/Se5BVLWd2/4yFiPTesTavgf2zPp3W91zRZw5985ljcKnTzMHDlGqFvc1p8
58adqg2hVekPyPwZ6er4aB6ksmhqtpZNk/IkKxNkDWz8c8s/OhE8G3C8r9N7Mg5K
NR2hpmg/Md2VR0oFJT5EF6cfIJbMj7cYp46z2STN6cODYahgZ3mo4ugtf19yOhUA
PgTjo1B1ub8Fzu116wgQpXbWK0heHumhWfV2fp7NHsq4ImTB0tCsC/54z8FI3HbY
sqUsZ8MP8gF4ujs+ZOx/kp1xK1iclwh18cH6/0a28R2ypn7uaQdzFTuGN79IXRXP
mIUqZkQxpln3U7TPgvmef/DTEKmdWRl/M3so2zS8cvF+KIC8AMiqxrrSotrN+vM8
sZ0N2Y6aEMBDP3ZZ/1I1AkHcBLltv27DgSofF8ZJqiBsQvpT0drd+yYop5SP+NQf
2ky4flV4U2MCj3wF/pGbUdqBvw4FsJbxoqEsPqyfA38D9m1YDIlZLstxyDYMNJMP
LMmWE8xWZ/Hcjd+ledILBH7RNXIBi+esDt8UTUJGTN/JVg9SFIQJrPg/7Liy/tJw
UcG9GD/O03UqRNgNsEWAliIOhICB5xk5rCZceaCfkPtaAaV8ky6J9KBsV67zQpED
X75meSeecStN51ymWzJnX2ktAvhU/uHQY6sDHcjDqCjvYuL6OZjBjz/uCYLsXAWf
lXZu1dY8Ua9ThiyxP8hGuYWTmZgGaM2hwVoa+JJ1iJb7LuaZeD5cJQD8pLQEy2GZ
tb7iIzzoCR3CjDVZZy6QEok0FW+vsp/yH9DXUiysiSzHGm4MzNs1FOO8c44h7V+V
y0j2SSJNXDTMYjSc41UMrbxVgSDksmo7axSMT2js/kiHHp+qxV3yhJ8IoHwHn23O
S5dIvMASxLW/+mIY7gCQtN6JTP7xHO7csvt+xESIJhGLTIJB66kmpQcbUer18WT5
4WjzcQHollnq9/oiloPzmR8TmYPaHqkEFFGz3oLzP5KQiNxTpneeA8aFH5jgzHna
CqzJ2TG6mpZHqoGSZE58Oqa1sKfB11hVaNF0Rg+32Gbpsvz8S7YAySu+NY0u90Mm
V+LqdBMfSOMBQ47Xk5EXEB4T/vTCmvmwEPQAEvR054XE+kowm7qwy2BNSDoO/din
vb9dwKnWoS4PrMP+K6I6DLPA9fzq5mH1wpl/YDOThzWKO4DT/qtk+i6CejDDOoVX
iLTCFNsTfgspQtx8n7DluDPcT6xJoiCKjzCkaHg9K9kkiURVNQjrUoLjReiqI4Dw
Za3tmoI4hlESGqej35w6+0WP5g1AaGfPLJ1RSwyxvi1VccwVAEfsaLnK0wuIqdVd
/WbJD7D/5Ng6m1quiE/vWTCeK8iz01qBRDbWs6N1vRugTkkSRNUM7eJ8MMtaCDL2
pYHLhFEJV6dEMWPxI5/R5FUKMMfMGVcSjjKD33d6htNkB1CoDcFcQPoSfFHI/EIz
17rbhioXruZoBhotyXiMtvBg3np1kaqB5p45Qkqdb4k+ox1m1FT8BxTN3UWtwxZb
CguWP/QSYph0h/SSgURQXAaijLC1lYOytQKI26U+zac89/dVD6jZjMkVMMfQmW4h
U7vYPjAEFBm7hDlAi9ItnMdda1r71Secjixq94+TaMHnIKu4HpT/bVWRM0UgjBe0
CHFLO6mrcAAe0hPamL0VsPIxOsBZlYrxIK/fNZEZTaro6KvcDstHfPObDgxbglhi
DYHEXiPOCFuy+PWNS9/I5Z9f5Z/QiYl49kTIdWgjVmyvK9SMpx5wLljKh+vHMdB1
X1wVv+K7wYUWNG3yHplsokE0uGZdG7MzbYapTatXIObUESKNn4Hn1+dAK0Ne1P3s
AK0IL1YnL5zFkNezoozdpi5oVAS5vXSenavBde/fR9oVQh2uKWePkkSelUIFP/Nv
ZwHYLalsRgu0M4T2Fh5BfnkvW5VfIChLS8BOxpmP/B+EPmGdzV04yWBBJdTaTqOc
tHR5wuzALtambAFy/sbcQe2hxOMqq/PJaz7O/1d8K3YT2nm7FXdfoSOsR3ZiCPRy
HQEbLRG4plKjJirDj4bHhWnw9wFL6oGkRySSumX6eziovmvjzTta4zinBwaDQDUr
lY5+48oJYpuUiWLBQL/uyz2a0VI2oE22Jo8u2AB6pxs9yaguZCFxF+iBmXMWID3z
Jg5YOsgr7lkabtwrnsK9DYMLEcgYZ+jMN+rrhjtbNVD/6NTn0Qq2p194yl9djcWx
fLEt+a+TMTphchve377OzotrS0YlSHiDel8jJOWd/ZZS4gG+uA+LPdrRkh5nLNcr
0hi3tSFdT+Na211LcsIA89C4u4NmH7LBL+2li007t3xLoSbn3KwKorvUOrFkVsvP
eYr7BokqC/htrU8uujEU+cbX4Ous9mgLhdeQqkGapBexy5/VMbVyWyMJF0mWGwpF
X5zEq0SPyu76Pwfyspz+SdiVI78/1Giru2K7QbjOmTn8AeMX3mgBo3uuDgHqr8gJ
OudJAf0Gyq0KadaCKe4tqzUqTTOiMal9AEYl7rWCueHuuom+5gqMRx3ytxr4v7Ma
nbydgw225vcngjGxX8rQvh9p6k0iktaIjq4fC8UbMAUWqOvazxnquEwHOXXiyfdf
Rnf6bgBk1jDc/eQNMcS6aHnINTxnzbEtZ5sPNi5CvmSU7tcHOOg2BkH9uaVFnaq2
YFwgU7jtjPzNo0H6ObyWE3SepwaNJ0FxfDYR4LK3iZGJQ/NOIOUxnhoGXWFAIviZ
2XDSrAj/gimtT7kSw6uUlP4XE/aK8YDRaicW2j0muegUNSCNb/5ExLz3pyI18g0f
9Hw/cGfPUx8p/w9NbN1kLavnmAvT23rvE7G9B+cvDzgaXOWC/K2g6o1W4NUq4djl
NSQafipfUZMbe+vSvm0lHXEKhfDgzAHwnVQyhETGgLblKjb9w+JQvFNZkr6w7KU4
E+8/hAe7szr380NoDWFn63TeECnBYVpk0GBBddCwSl6DPH01g7gdy0D+pJcQwh/2
tR7dQzeqBfIFM/EJ2cPeZvsE2ACMvS/QeZgtdAKT4JO/mqP6pZ4E4E7DBUVT1qRv
X2Mx+xrJtmg9iT9y+SJpwYPLo72QplLjl6KmejZxLxHi27/IBfpoBW9Jku9EvSl0
x+ffLKtr3z3PevsSCkmG0LYjYfnS7Ns6I5pzEs1hzARv7jq6R82cG37zdAH7mfI7
CpHaa8PrYft/gBOD6EKos8cXjik0azFJjkWvdTUJeCpskoBwS/hDraQ15/HvjTZ0
LS6VRB6Ze/iTEWODSPTUcO747mq7zLgwhjRTZdc8BxIneKtF1MxFo6sDa7cg3qfl
6lNC6X4fIaVzBcxKGHLz0FG3dzaBD2eopYxFGz7kp3/9YLcX9/YjaNjeaFPNAqPG
Y58BTTtR5tFBOQWiNs3N7nF8xbnB2Y/6P8xSxPHljUqVFGEZARsjnNVZ7uiaSfMS
h9GXVSumA6TwyEFwCWmtuoAD2kkr198rrtSud61p6dvQXm6XHay/84oqz1r4P/Ty
2cYkdNWrfycg731Vkf+MS3BIqQ05nc6J3g1/GKnTZERlSZX0JOh/ZvSAGofws9I1
VhBcBfWGKiFOFcfzK1kv8/kl1e9m7L+g/inCYK9llPdb1Uk5N28kvBvjv3luOJdX
UhBUpUSUSbhPDMdS3S/pGcikipKvFnoXI3fng4yTywE4c4nRPA/i2acsUG2dUeFk
pUIFlFF/YU8DfBV16cIeg0aynludoEWFHvpWYe1AJHQBsKpPpuhjwt+yxmcJ952t
FzOZ2rNgYE2MAZsj9Ny0EPeGXJeYlb3+zlPPQz2Wjxz2ksMDt3N1YYAoqmszcQ5A
XmhM7bHV8AumXA/ldH2HorB7GEYDyi6EDrygkmcrFJ/ckqiJocjR9kk/9b2v0WT2
v4Yir8SKmSVkQlB8tt3DmhkIb5hVaMisQMlLUbT0Y5TFPlJNAAeW0fnGk/zzqalR
svAtx8BGhyZCFLY5Dr5CtmqMtSjMfl872aqCDzgnH+BcJZtQfBFDpVyvyDXoaOQz
faMxESoR8Tq6y5xjHC4J8XZAEWCfAmpxZkx+XoC43YXi73boYyU+2VWEtF5V3nS0
3yajqKWefqdzMoQGkwCFrXBCJQQ7f0ftNwv+x1FpJplu07oIFR5WIqNpXywrJoAj
ANPNA3iuVDUvUDlurSXcnBin+saweyd+O7FV5luNxiXo50m5egARsDMh7gsjkUV7
VR9VbOvGEssUPBAjDEm24YNRCaGJFpU1M4Vojj+mHm9d180oiQ9GrNhrXsBuzEXe
MATdlMvk5svpftxWZAG/ub2rt/Mfi3W3jKudd9MejFqri9cK/rYRC4BkgNOmfs1R
v1CzOCcWdHgPgB1izdHBTq2GbRpCCA+KTjf72JWdzj/TrZdhtAug98Od/ivRG4Hj
jtkQ3LBcqd2exNuuUoPt7HbeVa3McK6GCj+KTmEc3+379yHqst+OwDIBq8BCuLOa
0RDQDsYNtSU4Iw6zUwZno4k9g7g8tewKIZ5QCDHyoBatpCbMDVFBk5yJ2W30zfHz
jBpUp0ywRhXfemnnndHzQlRNuhWOnoo9wNsgEW6+MK+34ST6qQJeidj4bAWk3E/4
bJ3yneoAdMrQk6pD4yzAUrdtG30YBKcAooV8vsknDDGdo/ZD0g1pwhGR98mYwvIn
p8AHcmY8Q7U4DyKXcL5pKJK+dIvTpDp2erYc5iZMvxBKyrh5dWqbcdT9bBaqyhHa
0Do+KLAx0flvNLswgMXAEo5veWp0ZhuKhE9DFZ4shKTo0ZBkJOUBfxn/BE/777Ap
DMxJB4auvLYOOYFiqvDENMXevzAxOtwZiA/BxQ7wivYgzvj8dUvj2N3ie1iX9rvC
ZoPMADAjAE4RIpjpMuIiZ/4Pd9ch9UqYkjqB+s84Vq7bRYP76y1wDD/ExAQpraD6
Ur5PsowgBvr/eBkAHkiQ2jyslD1fnaEpLtu3kWwyLDkKQxFSmFAfGgJOkBhUg2+x
5GjrjaiKI/EBzTcgip1SKhk6hQNB+hdOatcVOT3IPoJH+sv4dNrBrpEzV1ZcE/mN
3FWTZafBhm3+6c5yW+GK/SqP3fVVKMTedO7lZXC44FfgfwuDjv+THo+SOJXtcE/g
NbWfvKjdyitFppAh7BUyEQ6d64XcQYBhRCEe5J24fRa8Bt1iGT8yoMK+1ntTFhP9
6+5h1cCQ0d8cP8ZPt/NE18fdG6QdcC/FXYDL3PqZR2w5YIqXVnWipFUBb5ih5FYg
ixigApt5zAaa1o22QWqt4hFsnSxDxvVCufe1SSMRTpNRRnkAyhZ1wEH4Jzhdzvzb
3xJyL0wSZ5VBUXYLy43+FZEdekOKQuxxbxwjbb0ttPvqt2arNYjCv9CwgonyxR69
D9cPuqufKmsyYfZS2IDfqlEZylZ5mltRBGSKTpcc30hYvQBTNn/Ic20K92nQIypW
GN0cac+o9K3cxFF/gQ9FarBjj3uum4CMC2E/cXdfLcHSHNEzCYYaW8qLENS0saZP
20HvlktKmBD4w1gGWvoDn1KSD1zC7hsmhAh3AVl3IQJmw/yKFY3UnKs49B4DcM+j
nXqeADExbQiYlQZedI5e59jFSoCeBZQm3PaHtewJXYkO7d+gRSU1NqYVxVAupCPt
E6IYdbVsjOsjffbcpy2GQDioRa6rX1DXjS8raI4L55eqkIWZKr99V3dcIXGLfbHA
9xGgs61nc2C8RqMlhNEVvj1357MXNhfyFklWaeMqZXtqdM2ahKlUjZTy4fMwFtEj
gjzQXQ52WG9+V0RRUlI4xcrJsatwJCKg4RrHDwROFpg1+LmPbbc8aZyBxJ60pjE6
3fgOvet79IWmHmJrnCkqQ0Lds3fYN3bmvNj8IwFh3d+pUghIQ1Sso9MTA9GK6RSj
gh1nznm8mBHdYyrEWeGfeG/fgW55rfPiQwTnHjvxV6GXEPZcuudYe2rD6iINpZYy
LP1gmToVBYDnJB18jhf4mN9o3wbBtXq9tft/5UNt9Da+GXdA12aKZ7xfjpFraaRk
EyK66Q+UsUgUj/WU2EXSP9We7U/so7TLOPtaMlsOJUlR8Nrt3rOZ225STyySvk7R
vmgCDXJ5YSFTgUR68eB1MYM17QY3uEAC74P4K9/H34w3yn7EruItlS0CGHTdMYjw
inPN+3liYzksBAcp8ecskmNGAq6r7j9BFXUqBpOMoWDSV1B9GuEMR42pTcvwR0rJ
SEJytR72uL7YqyNfu+emu7zUgG4a4IxPAbG5hURhCTqLxfgecI1Ex0IW7vwbNsqH
1rI3ljiiiT9wtMorbE799WLFIMy8oEUoxtV/9lnu4VceVoVNhq68sVO8Ntn6R76F
jXd0aDk9fO17S75t+4PTNggR/W82296vuSC2s0GSlCtXdAVqNcpziTjwXUbZnXVx
X94JSTAilKerC6mUkpMv9CRp7u9g/idP/vK0Jg+RS4goP2ghVYJfLumJzC5AHp/w
hRhZJmHuN0gxlm4TYNIawKctn4ok2yIwW/x9hQbHdj0GzgPyHW2uvt5jhPyBCXQX
zAqcRXR5SrIWcWlts8zQB9SBf8E/rNPhUNSQmI/u8+9GSp+Zeskvtofcmh+rzrXn
phVeaWR7cqOSz/UFTPXzgBI0/ddhkHSiRfzd7S4l7LaIH5cEqL7wZJPG8Wtn/t9D
THEnTSZ1w5su8NpOROBkV4wk78ZFpDOOczvvlnph6kIOcd05XPgV8ouvk1voeMCD
IabDFWTZASyvx9Kg/PonsRrUky0uDctAbh4z6sEMHpoOq8Qtrzfw2Kacwf+l8eJt
frRqfC8Md7XyVVgfMKBslbQDZsgXzG0GngT7S40JUDloDsykgMpSwgTnqgcuq8yk
rGgk0fw8S3ZvY38NiuwzPKu36ICzDST4FrV/VYdHJm7oLsWF+jU2ezly+t5RV4mN
YViGA03zAzD0VcLQ81wUSaaywj3MhgtQbP31s4ddnZao02A7AevaaTQAKM+hklSY
fpJlPk3+/OGVr7DTnxAL7WWzZ10m0Kzy4U4JxMJWcLIHI04yxjbP4EzSu9hgWEes
KmpVQp0+CjsM7o4/1QAkt4DNcy5g62SZAsYLUAqlWUNIVJOxZlj899gJck61NP7W
HfQwNsB5tfdAIaNgES0WowYPunNekCnKKeVtZvTNR3tZlnvMa3/he13+ZHSRV/To
LoQ+0bqyyMyo+Y+jRlrFqWdKFpcYPYUQCn5h52ZL5VhndNHGgeh/vbzA3GIL+MKC
pcEOcQZuvB5yxQCXSM3RnEGCfsgQDly2S0akLkWPKtYeBe5fn36PKOKUNJ89uCq7
TzoPtktKn2RK5v4Wu9/07sjhMXRX8BHef+b31qVYFOW+7XXWyECMlKRzcFHI2Bcf
An9Xq6/AkDZyf6qcEYMEN9TEm36yx8nyQGUpVjOYnWZOWosiCxSQ/TVSPCaDlEEE
tjhrlBA84EssRIoZkvQSsPkP9iJSqTfH0NEohmzKjc6i50Xz8nfBwchCgvpn5h30
UMjonrRJgJvM0LbF2fMr1+1taDmJqa4/yFdkG1KwU748BH6mCccX7dfT6yiYSELo
KuhPx8FZ+IoS/NF6PwrdECPTtNlakmllyLbyDT7GJIvnz0L3PEJinJF+3E2iXVaJ
Ao5DWPFbzqDvWvMPOd6kCJWeE2jsY6IRk7Z4Mpd1ZlxQ5hSzCIGDzSHqOzLQ/HtU
sPePFPD5+yKi/LlWNK1gCYW94c9QBzTVhif9iMw/CrwjDw0mkCgY93Ddllz/Ne4+
vjmbUfbTbD7/2UD9N6KYRD0jp/RHAK8woEZvRiMZdk57XIqQYu8hiAdcSg1+euz3
kWrPFDo/ECYohxO2RPio8rWfddx/tCArKH7hby7aVTTPKdpr5wUMtfTkVlmeMgSd
pFaXR7HmqSknu7WEcBxurON32olrPuNG+FI2+f6CS3qKpAPJHdUFUW2D3W3dFgoq
OjD++rrt1D0kHI5RJlqDFMbjWHYUVuPulYXwIVE5LX1z3QVRN8gzxSCw1reK7kZW
CFJEvpid93TS6RbgBH+QcJkubUN4csGM2enf5x23AkAybE/osHMx+HgmBJ4LnT2i
8Ae7jJ5KrNos5PdXVT6cYg6seXfuoRmgkptyUIqO/DYOQSjKTimDwA2VuLwGrXhi
YqQ5wH6xMRWmpWzYUfofIkrDe/i0i8GRdTqsiJLyFjAAoh1FX9jO41ujT25aP2gQ
FN+CzQmKZHs4wMODNLo8uDvHmazPBn7Ef6Ao6TPf3Ni0YUMClbhtv1qZx4SbVLvS
LMa/DkKS55mnMOBrJWxWEyt81Coo0KSV6Ga8ThxDDSlTniVXv3ncP5FkYt8v6F7i
O+PG/CsexJ0DPxLy2K8j5PkIf2A97DZtBoCSzG+tliWtvrYLPXZ50xagU4lu+LOi
9efHEyF3Uq1sWgoSH7N8yB5T7pkuzNJH7w7oypzoAZrIoBQS8Uk74OGWZEBMEuja
7cDelTX9daOlYXZqldgTddgL9Mv3sVOEMxgH7UUvNDmrGm+dXfj1foWCxnppi8l9
T+9VLHcldf/SGTHLYkAMBg5MrIBk6diVLugvs2sJdENT1BxuOU6MlLYgb1G/L/DH
76i9nNap/+nUHpXoUjpgYWfOGOinjr73Nh7YOumUdVB9M4dTtRkHQznYoCLnSJcn
Tu+Sst7bu5BWHxo9sNv0qfHTwBQolge62O/XcaiQu5OmiXX+vqKfTe2peCr4tb3N
OkGsgVLCwoyAC6HpaGbtQCxoJnzyPLdgZHWK+gOeZ+AWBrnRh+WaYStXxSYqLE6t
j037DVMqQfdLx4EuLZn+Viwtrjw9SPB9yTfzhVBQazlg5ogF1azFfrFpEUCCKnnW
U7tIiQuXeUfX5AylC61b19X5G3zI7xlAwNvdv16JEF/9rbkoqgzjuBAELqOtnTKS
meltsAFE89bTdimaBsjJ8JCCI10iKVWdSr6DFynB1J+471vqLm69ZQ5TJ34QfjTH
GyR0bx2u7I6MPdztu9ia5yMXA85EF27Y7ybpUt2280+JQgbJwB8VoaCbe8HU436w
UjFKN11piUFfY3pXsqY0EXhXGYQordfA5htUqONBZu1A+eAkDZVKjCZ2rzFBn1kJ
XvBSoO1LGzqgHpVOZh0ZiqT5Z+Et5am7NnSqZppRBLNakuYM9z33bTvG84Ammby8
sSpijMtmLByeVbMLVHme8lp4aqoMGCAemHLZZOApsVMFGuBJRHHFqtc3UzQdn7oG
GaV/wuQB9AzVIImBVUr/nykcaMPV1JrxSLTyPvAoHHrLHnYBmvnwjhLNaPdlDzMV
rzJ0+r+NXICRhsPZYiQmsz3tJkiYzrRwLZS0EsOuDmdLGREnEMbyXK/HO/+bVZwt
DmpgBybgJPWxNMDhcDPqKL+Algcn/WtFdPxspg+uOoOpyib70oX7uyY4NbpWaos+
cljyY3SqNZz04vmTWHAcd5kKGtno7HxIIOnw9OKBGIBQ+G707E8VvLNEVbq6fUTE
CGP4DRw9ELzOEqaPYWnFeXmp/TaTPWdLii4902LykKWJO5wJcVfDlsPz+mCnJqz2
pVjsqUTuQfMzGpTPkNn0KNApWp1GZrYgDPpRiwhAElzJ56RjqPT1aUsgOPX+C76F
hy3l9ZYH5S6gG6RSSpvLIyKvs2rxjAlD8d3zqtySVIG+8BWp8nVqiSnYIxWtMPlH
7AcBsuYy7scMXKhskqoE1uIy0anpVgrmjFN7HWAQ1nen2c8oGmNls3bvMrDbQER0
tqaiDhGBVZB/v9K7nhz1Vollt1iq02k5+tM1YHA6umjs0NVtaHld9SCKwJZ4YoY7
LkqSHdHq11cFG1pQezW2DtqaTAQBN2SzGi05+u7s0Zp+tt4awAXlDoQzNEockWMj
KhhJNRjTDBifIbO+jQ9grbMFROIWl1s4MjaHok5Pu0TDnIPD/f5aJ3SdeltkrQIR
mZUjeMnzeRZ42O7yLPwdYA0rCItU/bZhAR86xtdbcdIyPCMQ+4TYzAQQwVCEj6Sr
/QZ96f+MymxagJhhi71/u8k6hGYyoMc3sLIwBfhQFaGEUTXCZNjHbbnfX9YPiMPh
sGG966oGfz+lNp3csHVi7O+Zb9twodh5bOMDCv7zrfHdoPlVpPn1edw8DuLgwrQY
jPj/3f0abVbRYc16LLvOkY5F1PHBbAzY/ARHI0+fAH8WYHnvjRnc+UnVVjDawE8K
VPCyuZc7bd6XtQ30kpSUkKNmVKBazSES8WuZjuBJkjXAWXeObPtWY14QFgUznEdv
/cl2cnmpv7VNsJm84LEh2ucAKjiWUJYELlgo1qf4RgWwycOeRWSdy1riWha1IiZl
Z+ybenRuc020SlcRM/TNIz6slRV+x8wpFISoGl6fKAQaniEuuFKN+BwpQsmd5Pcn
cqEZoHzB9mPIT+9JqL+WBlmtbStD7Gw6cohq3l8gy8VnuRV8pzNT9gOUzeDsKqr2
JixcV5ejsDbECCV4y/KbtoDVPHO0ww+456nEKykOCfeN+dglMRvA+XahK1PN1TzM
ZdRVFxv2FzcA7QN80flrNVCXH2Ep7C49gkKiqaSnME88KN7isoSlyGi+nnei55xB
wxolpbtbimurkam5zHvoXmXNvkesD9c09967PxQAw4yO0IYwXuwS3CuMGGBCvPIv
0YTBkjDE9v3Zc/7vJ0T8MZrsDKhoXqLFpCqVkldzVtOVBjsA5CVq+swkyvyjx5Nf
RVZeUrMJeh+ZOAKmzZfszFe9rjhChI022PfFOEaLD9at8fWPlt3BYf/vs3tygT4x
iXehy7wdPdwE5/h9y7XbwbIpoJ0CLOOLr/lXY482ib+jKINS/Gc0ANtm2bbUfIje
Rq0XNNSEAALFgr+RQj2VEbSggMgvmJ/2crYNLjPEeG+pL8g4czjqWEdpR7ePu06Q
sQ2Rknsq1fNv2vv8sn2gdKjgmHf04WdE8HC2cocDg7Sw7KkrhpnCwe02rnpPvXwi
YP+5kZ7To+g4ihaqmjag5HIlLvYu+4WcfiP1tN6SnrNQGCdwyj1r9BmCv8HKHeta
ISn7aYE6J6qLcL8+1NZOQI5cevh6xTGgC+xVhIbs/JD10t0hFmTZWr/rZzjsDcFn
GYvzbklEMPwXBHJ1AtM77nDCPT709GB4A/zNF2qrm89VSQRiFPOytlema05ANhWP
ylmwjw8SgxDC1zHcy0kxIWnYCWDsAWA9KPr8RPbus0FzQ5AsTj4ZM9yoUsu72qXg
yeNj4GAh50vrTA6OOrEMBodhxyiuLKjI36ureYZvrdB0V0suCCAl91O0OZjynops
SLvm9PH0vvyOOhIRZ+kfKIS0zXQlzvTRc0kssRAkPJWzr5D+zBfzo2yZdzleUUlm
/PK9VLdwuwpnMhfbvufU9p5QgMCwIvFN2vBtaIVt/8zaOUuO7T6KeBQFUt6FRZkH
xSomnRnxBZnh9Mif8zPktDE/6BvRPM647+VwsIhyzYC5zNxzgZVHR69BmUjMfaMQ
4ix69kTvm17qdfKg6aIIXirCa8vCfGk2E7wTdTOGA7tNGHnd7+4zZ4hnQuIwNgjM
5N+ljZ6rkPZQBZPfm3NjlmWmH2DzMaxX7OvXa4KpRIpbVSmz7t2m186avfNTngA3
nkzrb4ln4X1ryI4kCKJt8LY/bwP+d/2sJPMYlTgb4MTtr/A91xW6kldIpreTeKMa
KO0zW7/DjWPfjLXY02UFAsjYGW0cfa1e1fckskYYoYexdL0/Y9zyhPMoyx6Z45vx
rv02WyFvFH+JijM7kSM9RERRrSLEQXdNhEr4+V4OmVsOmAFglFh3PUXcGUHCxhpX
YxHRaAwBYzAlBw6yyS8LwS1kQdotKUSVq1F77Bk/VvnYpGPxhnpc25lugYe7lqbk
K/4ryccf4JBDG2oDNvc3rp96fQVObzoYN9+0DUq5NT2V7UCOq9AIEAp9fTlpWORZ
E+PMoLtn6nyVw4OOKmVdjtHwlAepwIXGCN8W3tcOF3upD6CAWqPpF1wQAn2aaWAC
O3PESptA4Dr8tfS4Gn3VupOYunXFDHmC0ph4zmpkHYKbI4Rr8ZHyLIMKoMey/0bZ
rAM2NkhD2NCTBnLoY5k2JmMb+tDTdtWMICWdWCrzlv2wRQkZCzhZFP77r0Y1u5r0
A17KKTfpBe4uaVEqwJuGIVVJ8BiBwjr0j1I0dfxdsXgQfL90JmsdXRH4g5/7JzR/
wcx3xSKa/K4tluqCSauBm01szNQe7y91qSpmqAOiE415n70i6dk75UKIUlCo9rYP
rToxVFU8F1yJyWQSu+EHmq2lm/mXJXNfhgA9tlT+LMMfpZ9mbbNdJ0xuamticGdb
sBUwCX95D6PxNVeO7QCIBOHVQfYHuxc4sysH9a6DSbLU8HUQJLnbe0IpxcLs7Ytv
HwR03fcECx7yy8C6THCr7bYITt/o/66g9F4zuhKD1NXUTXUoUIPK4bWY8ambc8cd
A2RlBU8CG5aTeTEP93JeAcsy75ZFz7n6uVe7KBgDJD62UEBe1rNIG0grFB+8uL5W
dl+8rgH10+iu2+8ouHnC/qZ3q+5LjplVFWq683G6egMkNzOr1ZUjrlgVIX2FeQfw
D+XncZu+kunfAKuf8b3FCaooZm5HzM4bEepq/4uxEvWkw02lVjxJuHtq93HVCpKl
uJJtw63dVb1+X0fIy8p1nfhpweMs2gljQS9M/0E8euNWauXwTVCy8UcPyddDKsUb
5XbopeqvBgwcoFoxHHwn8/jIaQfwpadFdkO8SFhmD8mOoZ0/8209UoSOHPnI4+v0
1OnBKDRXcqxB1QULrsjFYWxcryWAQUrsH6C7OOPLw+vrhn3qQtAcUJUCIEDCZeIS
fGlGe8+nevUkXtYHf+v08KlWIakP8Qp8bMg8P7MMxstCJzDu/7oQqzV5XfVhD71b
8/p2talyOCQUTKgr6tgDjnoNwmeGIAq735INN4zOFZQc7ldVCZ1A93S4Za47N8GW
Clx5fhkD+OJGon8miBORme1/5AYPiNwZZVoBMqiLjLNchjN0ZP68lJHi4eruI7me
ANKVAfOmiTRjW7ccUsa5IEqT800++06C4rRjV24NiCNIpnDzhegd0ceqNDGa2MKg
d7aGdQJxH3A05nTUKWMI880FjcXLWTUSJKncJF20SYF9hJnqN99t0lmdZnlq4V1W
WRI6DTC9yxSM6HYLThOXfwJR2LUaQlxQWp+ZCMU9nycX96TqI36KSt6Wqap1/sLH
JBGO9rluc6wulEB4IQCFgDtcFWPa+/AO4Mlp0R2QwkBJW4uTiiJxS7sip9GcxeuQ
coJ0WkQPRtIcOJjcrH5cz5MnB72R4yz/n0mkxQ7+SAlVC3mK8SPiEsp/7tPvvGKU
7445SqThzVgKOgUd5gcZrcgmggejbVblNfxUpvOloHCVyIhFVcYa4xw0mw0Cjwh7
iR3qzGWNpAz6LdnyC91O/5zBYGXJwFzp0Z3frzxAdg9QVT0y66tTyIvSmhxp5tft
fN/NhowKpD4J4LvbzC6t5WB9Re+FcqiE9f2cFk6LuWv/9k3OWxrWNZIFylChIOdS
AH+Duys9Iyw147dUIQNqUN5tLpVh0YH5ArQcjz+ppoXmtdtn1me3sVtpw25WA6+9
G+ORQEfKmuHsCbeBJiC9JugRvgsDCTLov8pHKhj2gigi/bkbY0eCcqXuO49i+oYp
wBg4fCA2Ue8ONv2AV+F9H2aWHbxjo5zdoZlqDQ5X2YK8yanpS60Nu0Kjh12TIERR
uJjCFspQPyEI+mi3zbm5Bh4heaXoDCrzUKGeX0JcUhIXF0CjV7ivnS1R2AoK5SWq
OsC+BI3xaihYYgRgF/JB7Irnp30aZdxvlUloFg9sN82I6bdCIQL8K0PCM+Lbis7/
HLwHbwknyDISP2lwhfhuUU0Xr4K0jIMIptlkQtDxT6RWadiQYBB0rp65i/Y1DYSO
D9fGHmFjVU5CEC+LsNeRCVA30u9XtY7OeGxboMtCVFAtUzzrOIihTjGAJOCaefdL
jPB1fGNUCjsFBsoo65BDVRN0Q60oR6Btf8GfZeKx7m21jezUzknspL2IEWK+/SG/
5GVggykEev9/Q++FpaJKR6wwS76yiB7ppbur6hK+c9s5md7hA9bzBqTo5xL4Hhe8
9dRl4wwd6aGFrV6CwWNqNgp/Owdwu5juNWQRXwjxGoKCfnbRAuSe47XkNGbxNBL8
50N4lTiAc27yk292/l0y+j0IS8e3ecU4LDYvUuPNrZzuoEVbNWTi3pv8l2PluqH5
Xpw84FGTb6j2RZZvF2LzelUijHEt2R67RRmD1a1NEQCtKPQrtYOEI3dCPVWkJDo1
kUiWyVczT+cx3ti7VyDSelLRGejyd5KAu2VCvLza5wl71r4Qah84g/3nMrVSWkVI
QfFWBEjWrTixojQndiJZvMuPB89UCaoQJGefP57BaUyYawqbL7IjUApOFq3mx8qP
DDD2XSCMxBCIUrEzdjbarGxBrlydcmuPu3VO4JYR53O/IavYVl2/c5wTJhbPpMSc
/1h64sX/SfQtJtRkOataHRdj9NmUMg0AHwVkxOSBHPDDV8KqYHrWvOTJoRVI2ujq
ifhwlOoYK/Ez22JtS/UPfr5WbxMgw6JQjfZPPMEycW7x5VuvNIKLlVFKEu2ZWAqf
xT+LjzoFAQinHUgSzl8BgnoQ3iEGnbLHSqqgWfObRvax5buaNuZip0oQb6EQgMtV
TXruvuZ5B3jNrxr4QKBWQ2VYhoAf/p3Bwo7x0ZzSjkP5xIMS2RmmoA+W6Pg9o0Oq
EWtkK6u1xG1zzo3P/O88zx1l9XgNJQ8vz143cQmmP+1MrSckMD7cuvuAwjh0MB1m
2LzFsCUtu81k6OnYQKsyn/26eWHZ6Q3iss6iOFY5J0SUaW5EXaRPvLk856bqAajM
h0Su4p7Zkg5AjvdWK02Zak0UHc9B4EuK90x88/TgZ7XrkpwNgdd7jTh0hD2PSHyv
xIp8SW8Guzk8wVU3ZHKiSP3NkGP+xZoOoiZVKNpSU4XQ0kOZg/uss1BZw6PRsX0v
vetYYSqWKgZyu6yO62vOw9fuT8T80e8HYAhQztBA0RkzG0scdL+pzgCU92LEc6hg
1HHJBCnWa5VPfjobgB5DYoVsquTVuqHb8qUdQ9TaRbQT7ouIeI8y31w1x2A3dVs4
WjdPoFxeCXGk47tYcNHJhosvqf6rUHzfl9ti155HUn1kDxgJ48tgwMwL0iEvOXhx
JYduLk7wcSFcwdei/tiiMUmfUCkGqwj1T9FC8zVCA/bAdUzhqT3rTfpocSbZtXna
vMxdRPttv72xbFbuRI4Pv5xSwqjpOASD1n81Bro3lgwgY7ddAPQTvRUgAabTY+WS
qVhm+p7EdzzqB2gOgZg1Ob3t0Ou1Zm12tUN9333E1eEfQE3itdfGqlG7qrmokXnc
OWLJs6lbOESTCAcI1U20H4YZ2Atp3oUOcuRuclcd24e7NwgtTw0sjnwowDSkHFqt
K6Vktkx0R1P5AZygsZqz2Q8QbTPjyl/IIWpYVtEp0aPJLcZOOa/WH9lXfmNl0BcA
LaoIAM2xh78J1Xtw8qoUdJ3WCAwIZx0TPrVZGeHMckR9RSAjXQeTLwitKsvuA7T9
Hpefx2GBrm2t1aesODfnxNPTJFJNd5PdOOmAqBd4LDtTO9av5UZz7SAJuAtIJoPZ
psSOHHh6+wKW6AVe5cQDwXMtZa5jxN2z/MnVDCI971NwXjs80OuLO/xi17gBRUvB
j7iIKA2KKmWNVDbJNXf5blAlKADCUFO7GLP6c3BIdLd+WiLg3Qsn1sF6odUf+e0O
XiK7quRbYC98uhl8UL8DYGXl1inOIZexHIoFx6mRSAWVFU+ArSYyALOvFeNhqx8G
pFJTPJxu2xDEkgJX2mH0BrInjTxCszuDsRMpC8qAh1xcJzBKnsTmpj94w921+LSM
b+LksbKo/toAYWLt7ux8dxAeb70WnxSkJD7G2IB0OA7HQu5fsqbhOFOt0ycDJZrC
Qfbu7kaZ2rOIwjJ4xj0OXd11vJIKqFyG8ZiXBcGeIseXwQZFzsttOU9+KWjIE1nY
Z19w2/BQgOO34oTS2QWzNdxcnJwd2FS2QfpcXTNuc9CWmbZ1hIdDVQP1BN+lHUl3
rirHymTQpHUBtavLqtV2bLX8Zr4NJ2vKAmCCfRJrPQOfVGsUgLy107S9jukrnz+5
9GBZuMC37t9ljdSBoGDpwdbe7t5BUUQLLPo9dPYBmQyemv3oGDgeaovDKoYNjdt6
eRZyMEk3r9AYFG8WC/0Vj0QStmdgdshLmp6q2sG3i1tQ8HWqKXt/xfLhCILoSSEt
nAP40Pa+V6DoSK00KHpSmkRNzDQGquxccAgIguuT5pALTh6wWJ9v8puDs+vL8YZg
0d4jJ9Qw04SEGcxVls3ZAytM5Bx5/AryoKruHV8JPa5Fhl1FFZX1GZ/VxwQNOjw4
r4eQBdUyeMWbo4vYjK2LLDxjSV9BOVE7PxAgNdpe82HlWKSYcT/Qi6S58quHRlHu
4SAJGC4WuiAx8LSW9d6b6gXY9auN5WM2gyOVcXKzaG2E/oFz7Kror9VwlUsqU+oV
tGXVH8YNSFDMwcCCxlRBgKZFo97GM5sfQauB/fGOp6XD/QrUVGtxYl8XkbMTZOFI
Zpnh2A+xRMWcR4c/eoYfkjESIFdrkMvHMjMRrM/VjSlVNrcKDRbNefdbLF/W/568
9rXBkWTADhYQV24mYqZEjBqeEzWrkzELJsFRxHRzHRNORk0dAb3ehDEUsHvE7yVW
rLRM4O2ndnRLf7Vpi8pfoTJ4QeYQcRCt8I5sLd5BVNUVnjG6H5hYACKK81i2AjN+
EX8z1qWzA6AwSBGu4RfmymGDhRgrzUxpzkZVMRpxC9JCsEP9XLB7HZraRlLAq6Y9
zqLsvyle6wPlgrqz+G2CXhTTV90kDwDpH9S3EUUrIrNCPLJuuEuIdOOGjhuca4MP
d6L4PMj9GEsWZkwhoRlAED+XFwuopqH1kjqkgCHPY86vB/DsJkdH2rOHlsJqrIrJ
9i4EKpHVOLawwHDcb0rO15nrgwZmPwroDCRBPp4voPlA7RuNjPfvuXWP9kceMSr4
btVl+JV2o4rvktD0aWl3EQ998sy1EnprryVH5LPM9q1ccSUHxM365jLzL7V0EIdn
nS8aYRUrgTay/kNVm5KxOHEyvgad7t5ioJt6C+2MskkRBAV3ffoVGdJcY4cYD/va
yuoUnLyCAH8CJtzmtwxB0rjtFjUbSyacFE9IqP2yw4vqJ2i22qWqMfbtgGfPNtMF
b6KYqcEHA0GMWXfSr6kgoRA3bB0rSHvj/vhAXK78ur5usi2vA2jX6kGkzjut1RC3
c1OKiWfnXLrHw/YNu2zI/t+bWykd7lDj5oWP4KOSz1dH5sbGtLMky25grH3Xw2Gk
aEURSF+5WbWKE33QeFEEswauUs5wBJvn0v7qtz2xHv3ZWz1YV5pOkgOPC0+BwOmw
lUdIYI0QHBMdUf5wwRZQtSrf5myO2XF8A4E7+KXq2ZVG2EMf6y/3WlUvCGkjGtJj
GoHiUrYv6/mf1GFJpfCVHX24i++9g7dtibn0IC79G3J7YiMmzDkMpQRgkVy1+GMc
RhBddH98ztabXDQiRRtEruoBSGLeQfA8NXIkibJTY/+R/ti48Z6IPkthWq6EEYa4
RRpGiLhuajtxwYSgLyiIzFu6BQ5FCPTMn8VTTc8Lx35l8TqhKC5zSbS7AGMJAGgy
ACU6UH4wGhmV8s0LDEbpKbLue+9R5yW971Fk9W0vVRm89iW9VKPv8rc6QoLDDSVZ
MSV/3PhI1/RUgDl1W31Lo/CVt496i00cxewprQ8SeIhPiVhAkzpgEJS+oFSg2vVJ
e600hEOFdsrVmGH/mawxOljszobJJsICbYGVs/EtDEpU1+jWZXfbnbkTTxaEIRmC
x7KzCtPwrbaNGxwILPpKAgHZgLx1Mr9hSiUVxAIqU01Yd+c8dnXLa2t6wGRSHISJ
SqhzbtLAwK9gRY+8IRGwWbmNdRMTLwFH9HI8clEu4rNg2Hh2k867sTKOtTmPJXm1
LLXeqhsYZwueh7r2HqbzIKT9aZGmU9wcL7R12h9TBzNRjc/xKtSVzZKWT3r3o62L
B0xYcUS/whJmtQztNljzfQj1Iy5M7DsavAdBdrOSrOqXiWHKkR2kkPxnDpI6VSxx
626Z2EREQ7uuek7I4C+xr14vJTyyjwGnD9dR/h9YYEjJvJXfXpz4BxNsssFmHcMC
YahxnJ99rCEyCqrVKb+C5GUCYg9fA+6HTe+ya+hZ5GrR41ellHLMtrYDcDcohwgX
ySSZuPKHaBdDo0zcaxLcZ1ABnQZ0Rtuwn6FdSI31ZMpLjP8o/kmgMxS/R1hwN8pq
jqh2H+TYZ9lVtYpl4nbBkm6txuFxqQSUL1OifWdYvzOXPqsyxPPqUbqEByHefUrl
GvWRrVE9FE8UBMRYpj6w9TGgGD/hITe8eR2Yaqa4juj07RjNc7zynI0xJCNIQGYL
bwiibYq+/wD4ri6UMglbZMGdtwKGUNVz//LVgTrCONH9F/a8VgdjeYTbPg6DPlF+
42u8IJ4/Q0fHwU6GM2kYwXEmMwrqBN3Fv1vV0vz6990V32qPrJLFsRShUUffIjpw
8T4BFzq7W0ZfmYwFWzjs9ZWJe7iMzIQhRWhECYCOG9DkM5t7FJNilBQ393lZJul9
7we4nxLenCaoYK7L3m9FGKhRZE8TPfSr4CvmgkuhvVVKp5m7nkzdReVNJFQiendA
Z7RSvstgpCbBpi+o81u3qAuLRqLcSea9KXnb23cdyhPrvYEvVhUV8k8cfIb7MjLg
fTuTL4+n9YKn1KXjTbZSSMQOvVdsmmOT6xiGuxcTia0YkEUu8GeG/PRTVlkiWyPK
QicsxwbEBsPpIjsYGyO08nfpSvRTpdhhgvlFn0SPiaOEqWmTn92cuPb2a/2fvEMP
EuZmHW2iA2Wg29AEkQCoDXH2/lQKROc9NPCA0DYBVl5f8gn0CfalC6CAoskjNTuq
izvqt7ZPTcwmBukad1s4jap7fvx5SQslMgu7+Jb+FTVTYrSx5kcItWNsnnZhvENu
uTAFPO7RxRksicnp8+BDignbL+UjRByKMd55+0nQhtmqLOdT8+IneG8J6LYH1hqI
CGH+SOA4G7UsU9cgNwqMn9QnYpspb/7opgZx8BITBQCnP/6p4IvutqkNGYfjRc4E
DiT4CCw3cS3wLXkgFAZ5ETuswxhQl+P6o3bzXzxkyIIU9+U8cWVK/JC+KzDaeWy5
/1F2SyPlZwR+ehl6g8ytWwbS/CrapNYTGm6H8eBStiBMOkdM6NlN6pZPCriA002w
7JuiMVxIEE6YDo4if0HNbPthOjkK8VszQyNuAmABK+rsM+xx985g15vZsBPWR2oa
AfG0WDafxYW8Z+j+P7Feq9s5vC5/iQnBETm1hjnCysRRThuyYj7mzhvkEkBlYwyb
Um5xNacdwzqmxECvF+j0jWXDWHb7OM6IaW3bN+S1YKAOdldD/MK1LpsVVFuYYVvx
ZCcXDefQKIkN4DD2XoA2ZDDMf9v5U14l7Bv7C91gXIe5GYsZMZBIUjkd07+lyOYr
EvyrbZH35Ix5fPU3yQ3hLrQWQsuM9izw9DGZl2vTfkVJkmcqDBengZIBwmgSR65G
f7G7s9rTHMTw7HHhg0K/i+0qqrsfjANQjDx7yUIc0tjXzBq8s52DU+uKomNn4RXq
lw66LMzxM6G9rDj0z3YuO0tWWyCacoCfb54+r4xxuVB/c/8ciXpgAWE9Bsj1jdym
11kRWDY9PPl0MNCN26CPNdQXj3ozko7kVYN/OvpVWBo8lcaDXW4Flq1GjA/WTjUI
n1mqyDizoc2Oy+hLnKNX6Y18uo/CguHOC6Iicl9BymrKyjTQOjpMM3DZFbFZxB3Y
HbgXTA7I8wgKqN0tGaJPAAGYC1ryJm51weGCuFvCD8cfnOACvjPDNvm2bE0K0cvL
x2/mjrT+dsRXpR3KsJF7DnYVsitgQ2UgHs4httoYWWAo1prFOr4Zv+Ah9G6e68Cr
8G0yXjNDa/vAcWa8oUl0fGYbhwlgCVJft/A5syZWrU6w7eq2hVRXr0A7jucAp7lV
wzCUccuRClvNLi/fnBVjQhNCc2Fd/2Pfh/W84SfofKJmiFAwf/JkRTLpGpovLT2a
phgA6Y9OYDdCuvvRqoeOieVjaqc1Wf/H0lPFDCOS75tBQCNLgcVxSgQT/Fj60GPf
SmpzZzY7aAIS+XWB4bycUa8mpA1OxjiE0UqbS9+mcekYGCheSKwMnFrkmFwtu7YJ
fFsDRgzNVIW6xtTZ7zz2u8/lkeZPvYo8MQzB510LPt2AzEV3L3FH1MlKqkEIn4Qw
RAuJwOIQDJZ7Mg1c8RVHmcezvbU6yn+TzehLr6ZDXSC3iaNZZR0+ftvp03C8npHz
10aI47Q/1PIdaOOCDZRlWQCOmiWP+Q1T8RXezR3vBG2Lh6AdMC1uXmxTftRFLzRl
CTdDgI0UCx2zFM7v0HfvWs+6oJgthUqNr1wXkb8mJm9TJEFxSi4qPOvOHC0EYlDR
QujSP6pGFHZDIDNiHeX/MpCfEab/7DCqC2sbJleBVvoYotiAKCE8g7Ew29S/4M0K
s1Mg4YVaHgZWFVNZiw8MV3grJtUcZtchfWFRYpcIF6NTGUGsQmmLCpEiDy+ffOOE
Wl5EdF2AYkUGi2ROG7CzDNUAQ5F5ezysjDJFDRB8NkT4ZEOi+Wdheg8H+SX+J0iK
YBgNxAuh4PnslMvh78maDzbjK9cttHaefqeEcXHxocX0Ki/bNQRF92xSyp42/dm8
SV1cypJPq2UQxODFfrHFR3ljtx9GSkYzbUUEdu4Bpl8y2Ku5T91Ro5X5OBaQbTrC
zFSVTaYz5wkCZ8hIvTsopUckWvp1MoDka6gEV+bNjFDAD7o+Q+jFRW1BCU1qAgnQ
Zt8QKcUOd/rlZisrKmouwVoaODgwwQ5lu4oEkMtqb8zz+9utqFXr/6MnPQ7wrgGv
+PnXNHMe022QCxBzLPIvhmHVjyPvUgR2IdEMStDT9iKx2aZUZ0UA7zJ8yI2tmdLC
1JdRQQFsZdz88mNKDlpy60vC2k7pS860dfgYp34TZQdQDbQvyTW1GdOgjq2iTiDi
SQRp5tF7p8oYFtkH1twDKNrsq8MVPMozcaD31fVRWWVXZ37gL4ApxGqmbczGfFMV
cnZRGWV2lYm8JtwpqDlDVCTNVl3No5dnf0LrhfJgpbvHubRFT73r6yBO5kdYs+S9
MOGDyU3lhf/0OWHS+4eyDiD72rfWE01/GqocamOeh+GqU/bt3IgtWRMPFjD2PiYc
rwGbLc70CnPTA315OGoiJc6G7RcCRpiM6ruNCtg+ZhGCN8QLUdLhCY6xUO/QqWSx
Xn49nayRJgyhhZtchfONlJ2NZJWMU2zkSxjS2c+/pkD5vyULNyjV9FaOI++MlM83
KAVnMpDO8yTE/NGl1dG6m0TGuAIoIaqg0Vv7SyFQz5zuCyjJW2N8JCD0Ai69d4DT
yzXDVHt1s5yx/3tv42PaC2RxGGpLFPWa5kG/im9hBRmdHq2ABx+P20W9rrlV8pI5
QkyxtZHEdrKNyuF+eNNUZaODKxMvhodHTQTtPQrvAQgfE58In0ZEcL3JexOYEg66
Hmhl1S7/8ocDbhc4k2c2TmHEI5D2YqczEv5fdvKamSU3ks0drYD8kiSZ4cAFx2tP
D5cdm0enHsH3iPoCn1J9P2vx+jYvs8qu70RMTy/HF17WAGgKpzLPABuibHbwYCpF
LGfOCzaOfxxal8uSnlkFUUCFZoCp/ZPxiPqb3sAinDcw/I5ffbR0PKSk9n2tzT1F
xa+ejMuTi+o44VyOtAfQfbM8GaFtyVRqN8qA1mi1AT8TOgtOHCTbj1QqjKr1K8ZV
vPbxNp7nRmTPpZINoV7YsrL2b6T/zZkEnSf5DcnGg3Ol7K81DBe3BxmkUI/GvMC0
uLJ9OEMSPDmkuJsgN+ysTKmUhMOHKpg+7s7pMp/GdxuEsfoeu/kgqaUnx9s4mF5o
2y92CUp2mijK5OKxKVPH5nVpcQ3mkskzjvV/L+MAI+9U5/k9wHNmqasfvO7TglXb
EUYUR+2v1ZDXvSrAaAp6VNjFEKcI05uc3d//v+HMmnqXOqhum3ljh2sre3pzq78/
A6bbwzHsNegNv575vbiR3fHv+OgXc1LJWoSCxFwUq80YYJ4b/kS4uOKKV7aDAnvz
1yvEmwgEea+iHqstDBB4ABut03dsJrYYmSaAR6JBQvQpGBKYlMp1HafYb8/00JxL
YN/f21RhYWXIpLnCrDInxD2uhDIBdZM9gDB8Jwa4qo4z8kol8+gcrLukNUo74jRb
6NjucRPxNzaMsAj7fpvjDiw9LNMnPyM+DYHBESKMgre/5ocaDRJxecnzjdAsDMtX
SwF9KB0gG+IbxpiRwym8trM3DJEEwRTRmljrbk+H162naNUJXT1uVc20EKmbrpOL
JZrPA3U39Xd1BXQKWvTgOviqCn/cCtEfcHIYmOC2XtL25h1WkW9GguEKOmxOOXHo
BRE/Zlbt14Qj5dp3eimS5czHJgr5hKf+hUIiglbP8kF006/3jajbZMrfWqP/iHz3
KzTFUT/89un6k4vJzPJF0WFMg/bhve/OANiUJYFvRviAkQlSABycoRAtSCfclaO0
0anHS9WD65FNKU+tUnvS3BkRNvq/HwiuwD2YOg4T3B0YepAxY+U21i1vB5OL2RRm
F9s+AKK4f4PaqXnrqyBiWz+O2tvphgKUY/1lEQ8irvODIcM6g79mlBOPp2/sElI8
GHDk2Jl3/QqV6b8QO/uGZ7RHcCO99R5+L180R4VBVJU0eDNX+5+gpasJcM9XBWI9
rBW0+9nMC/v1reQ0u8nvBx2dCNH6ybEeO8socM8glhuFjvNeMMVUsb+gDJpx1h/W
Q0CKjLsNiOA3fkvWfuLy8Bn7lOXsBAAevEGxjW1GekrtJ1sy9J1KiRGsAqd42Kdz
omaZYgQklAC1GgL3NMdcIrnNFjxECVRgsylGHsrDAKAZxlJK7ICuDOjxA01JUwLj
Pp6Ys5pz4xrsFb57lIgxNH/4xB9DH/fJVdQIIcVNDs8PfwEwCLQOCYB/xgmViaav
e8ogsD4RaJAa42PgaRfcF2tbs1gDJZiKoVMui6+lBinbpvbDYi78QC2qM+CAcMts
dR1f7nmV+aU1LCB71I4Drfn8sMYt4dF6Ve2mcCPXzZ7WEl+cHw2ZOh3LQFFPSYhT
W7m6dUw7OyoiW0Ui0WsnyaSr21/i4dYmNJ/C2oCq6pcCCRozom5uKQDyhmU//m2l
PjI3QmiG2+Yj402t8oDACrrzz1mXrquyHW5wMcrj6wYUpQnnBqque0r8CCJsWSHv
6K3UwIcLt9eejFur3RAbwU+bxpjbHvazUPvgli0V+axWOfTpqFlDo7JsAq+Y0fh9
+TUYe6tZ6EQWy/D0AwklKYiH24YaEfznXbRxvZSdYfOtptEYwpN8k1gs7CZtngJX
LimwSvZ3UK7mUALzgKwh/z7EC+iDz3Jvi9yCSGHA4uPGgHmGhPAogZgY/kOflU94
5Jb1CMeqh/EYPtd35hZUjCEu0bPI3D62p4ilqv9VkpLhl5btNvcEbG6AET5i+ccz
AuOv+fLNbiYy6/ib3JbMY83Fn9hb67QyaO9lr2xyQIl3af9Qvay8VR5+oXOKivSy
DlBWn1rOXhcC7NdiQyreYgGN3zt+AJA9EEI8fje5okiScMEkitDI+9pzdBaXmEI9
feOHMJ5hhx91KH3fRljShGRDkShXdsy0kocJy3ymT0C/YJ7n73APtAPBISBrR90u
/BRbqPc61cZ4+kkJmlIG+gZg8L8wpsrjX7yDvwsafJwrNH+/mCp0Oa6peDUiAvMj
xwNF6rY6MzNfCQPpWCF6XneovqVdOM3tqdbN8m26e03taQBtzkHLKmqgfxc5ofJF
IypBxGUpD7i9VNDzQmKE6p4h+rtj8rs4giZj/2y4F6+lDS/lHnyp3uX4fHL9lbX3
KFDxBuZqdG1CHpxe+BkvGaZg+OKla/BLYgENRPNxUCCuXzMbOq8iqEeotxJIHjMj
agnQnWq+16COIPBLVrmHN5lgT1t4ZZGZUByGMyp4XxOQKKpriJ6BgYCuhdWWIej3
IfoyH/Xfm+ckda5nLm1bnKRtkkPGoZUJhtuxhtsy2aCshIoParkNV6aYCGPkIYFk
6LXtC9U8dGVUXlhj6kEgJ2f5rmtOliyY3yh8lTHk0o91XycPIYxQwnu9J7cGq24Q
VuPjFT3aGkXusj+n9Y6Do1ZNASG0JKyngXlrbKOnnpg1oCbgp8cF0xigbBHrLEyn
66GsR/fKPJkyVe3vEzzW57gzCOwBP9SLvjNJ3n92J6QMEMt0ojeMZqV0TISArNOG
tjU6PtUKv0TfYk0+Wfe5zbZbN2T98hxrIip8CELZF4wkas430BMoVNEAaDKgB4V+
YYjsE3Pu7k1djsro0L+e0rnpwQS6DlxDGiiaLKAWYujqgYfJZ6Ld1rxHurlLtJX5
GcNQDh+xlOv5RLc7BNCnBs+DkpPUCoOfndDa5NCiywpEyP2+gJhXZqH+69EvYSni
IWdfD/z/o7Ur+XZPV+i52vum1wzbjReQA+tAJfT1J4EokoYwzM1oCq03Jfh20o3T
vaq95KcjelSpmcvXxElWMAFT5usSROdRsuRzyuevwXUPnPLWYTwl6dCyO2+E5ddt
R/CYgE6kBawF4iMgaERfqX38vCqqHFO/kLIKLrobbiL+o/sTj8+NBJJXjEJvDGNq
cQFoiwhfF4LCx8faH+mYG2l5RIRZRoWIdSS+C5E7x363FHJFqRHVC75aUbRONMe8
S1svywQlrP/BNdFDBLiGDGjsMvUlCTqULoK2XppFkETfTNoSVcrcBgrMxUsAyr0K
YzJFXVaoQHCg4GLGrVqyqX0ijRVpi08mDUe6tT48bQXVkD3UZkib0VBGWWP2fopq
C6HbGdjlbkUsbcVeEpwAMFQPWcXiAep/7R0r2SacCoY8aPf/3grw8JnRdN2ohtrd
Iz3l7nYp89I4cwDFN2feDT+IUNuPYXczAVqPRE/xra3jkEfXI+uh82TohJsBJEZs
OzcWmruhsrbQWpryEd1+AidAq7btq2RgC/rUEl0Q4ftE6Jj6ikXUU0V7AkXEigPD
AnNgbNdLJMSWPsRzySX1zTdK99JTNbwhGLeI7NCfIqrhGFKSqtAcDQ/KJKCv9RZf
QgZziXSN7ydMTB+ObHdRXFHp80ygFMn4wPLx/iC4sY2FFftSTU2JpBWkz5h8ynqm
JkQC9bUlCZ3xm/xHMobpOtpg2Q7rR2hyizGm9/rIwDzAfnuoDL0troeJ14K2mggq
iIg3YDxxiyVofWl4nW0tkIpFXlSd2DKPruzfO/v/bj305EYveTzaqxIPy0x46FaK
CVa5vCTMpgxSX+xy8ycao69uvOM+eNVPT426OdVrQsNMghY0u7UKupJ9+yAhx0WS
VJKkwZvKItgLnautlXMfN4UHMYDDbcSf48bQG+D4CYWl81u7Bjo5OUSPyg7rDWTm
94OpywhP4mx4coXuWtjmSrKvdJYeoIu5M/WatRJTRQI48fJ6m3jwAghmDddxVfSi
Z+6vM0kt1NLH21DKftCtniP7qK4vxpfp+teft9u4IyIOAd2jwpniuYbNXRVC3dD3
WS7Y600l9exbgNBx6HQNvp0iiuaSadlAPuhe1wcn+TCgpIKPOdbdxF3K0h3UdM7t
csx8YPnck6giw5QkxDFw/3PH9FIrhpXpLMVbPZCzd6K7bcoH9+boU1d0LwrgL4dp
dJgMUHb2Yb5DDHY6utbX6+uRSj/Au6TwnBACHI33F9wey5TeJs4Y7SCN7pJmLMza
dFwCkdgua8hexltsn7amDr1RhtWvULLG7B5o6FP9noyCPZDbNlVtLttzKAxaZBTG
AORjzhfTQ7s/RN7+xFFgURfjJK6wHhTxGoXd4hSMqcr6wgR+22DCb6Q9uiGaOAJy
V9eaRgcOumr8Fl0PtAMa6mJvpRBGPOqM5EPF7pV3zU/GjDDA+SyTvfLfQnqvR7NX
Q+XjRVRq1FIQNrrhTsNQFCPBV+Xukib0i8ZgfQrsuwMttEDrEjSkA1Ruq6Tvzu3h
OqXR4Z0QebAWagj9wuQ1TeF2VRHdLRDs9NK1YM3ZUiPVqj7iY6xmswRvkvDKb1x2
q23yeqirhT/RqktAAnOBQpavxGntJOzS3Ruvlwy5cWChxJdXrPKenBzDxcxcjkyz
aswzZBHHGQkl7W8Qps1m5ta/oXErlphC//BWesjIhSiMevAs6kjKkFgnnIeXEv+J
NYds8XRKN0R9zuFqgQGd8YZWY3ik8Ajmg/D91hWB81wqxGpzghCpjbYAuaLa0645
2BS/R35o4OiTgJz0ZpDkyqG+lAgOD8rW804dDF6DtvmL0nCeVCIVwoiVot3Mg8zB
G53chtq/5Kt7tBxlraarNvmPRCOU/Qv5ROvCw69Bn67q0fgYqwCUWlOWZPl+fOUW
hK//fCdzNBJpJso75WjJ+P+M/DaF3HjYimcjcPvqXgQIBq3+jiWbX/x6phGJadtY
AQSQyEB2q8inf2tz2aMYvQPOXE+SoNDrfe6pO9qVQhJfq9nNV7cwXdq7TBh7C5TS
u9btMtSfFUb/5mYv9uc+rYxDjkFNY+4l42w4p4QHh9zSk07oZXCCCYTEDbuHr/a3
7GtHzbcZWHAvY+RTSsmWRHOcbULQWD9dBU55r6LW0aUSKqPRe6TlSZ8r2wg6nEpG
e63SF/pfXwWJbqNAcdnOZIUaUZ9yxNgw1d0+C0/q7AYbAQVz2XjW4COodXol5l4c
jNDrEo84MkgRr9XQpcgR+GD7IgOZ0fZnY43wBQgl07SFg33W1uEAxQND2+vBEvs+
iwPOCKkfy9iszD/xrguutzmBnwKkvWmbRV/Kw7Q4tIWw5/uLVfJyZaZTgA5/NX71
LJ2td9sX61g0RMmRvt9MSkDFqz9XcoeK8qxWNxXU94icaHvWpYbLAt5d8pqTKDzL
bOj8vKS2QLvAr77cYZVVS173UH+YIiLCq1LCOZIquvnmDxY/RZ9axm/uHxib2KGg
XbDsa8yxKb6HzBXrR5DYwk/FRbYzMMKD+JitYeDyGfVrRiNtPo8jJrxWC9CBqn5p
46A0OdAFXYui4ttPXiMVVc8Hu17Oa9YfhHwZChPGy0x7XO6cOSaslOioi9EgqysR
29hUDYF9cc27hIN3qwO4IuOc982uHqye3MwlUzrqMs3MkNqsBcU20S4p6QMcSkwq
FZT1p/8kM7fDJhvm7BIiuICl0MkTEe8/Hk7xDKAqOB8RQZTRX4QlTRh8NL/Ckvqk
inQhUGh/nsh/qWbvUdqx7iNnVmjXyc4GiLA9OtPZ10nJW1jNYxibpUgzHAlQyXWs
PUiAnAeXAiA7LzqRsm190lcgLLK1PJfKp+KQh+MI3sWVXRc4JNM+GYFN5xPbI4t7
jRTVdkeP/ucwjTXPO1Ibi36H1zpukEwIe0diqS/HjgCXgnjoD8MoA1w1kL+jj262
ZavTqq+2oC3Nlo6Ath7rrQ9oHviVbPhZcKnhPR3PU2GgHKatdXWZ2+MoDrnpm2PW
y8WSg6I1P60FaB5k23wZaSd/jL0ZqyEF0WIx4Vejg4bbdTeW+4WKZOjFj8DB2vT3
HpMyVARBMf1a+gvngMLO0xDWfIipU6CokKalIHW3guqKoFyfs2HA1Q2xjfCiTM/z
FMU+LMFGJ+nl1AZH/hvCRtxsayBeDE9qlOOuEOQGdEi0kSByybo9ZhvLpjOZAcAW
KU2ZcNUbBmVBfKpUmYNHhGPpp3/5nlpvYRlva11qx4WGf0yr7FnzDQ9t+O277kcx
T2PSW7283QhG8Xj8PAa4HytbhMnaxxu8bZjzbh60teTaFeOOVpDV4TVbhCRrJvuc
AmmhW95TP80D68gyCWy2zmI3Eo55/TIkoScaFjd8rk0ai8Itj4WCcLqwl2YFk9RE
Vfj1E5b2hMKTkFsVIAnO2elBNgGGrFqTsAaz+quUgSJtrpiqZ+li2yMnEPz99iXr
KzF3eVSSE4ctCqRrwnvOTiGoROPISsKFBGUfO0uX3v7A2Q7OwsMP3SX+XuW8fOXO
w6VuTJNCCbkX/4M27VCpFAPPHecG1kM3Iyn1bPXnbjPhJAkWxrR6oRseHVl9EC2B
13L8uiI30X6LieIYT0LQuyxnRiM9ca/DIjo8jVQ8T5V1Ky8Je2m6MumewRPlfmBr
qs3O4HI47Ah1TUEGmftsoiA/iod2CDXaC2ru6xIrvUHjhToa0aUSljBGwhP3gURB
xZOFtcBMQfZ5h/n8c27X/gJOVxzA2robsnK5gdBs6eiycexza8/wWoIdF///r+wI
EqyZggkdViPbYWNYRrMqO2LgkZ4VzbMaDuvEr7131l7HyY/a9jU1DvFO/uGx7xOJ
0PF6dvH+WE7UCGQarr9W3z2PPKuXMq5oLw03al880NBCGeOXqdEOg+RIirRZhHGS
8WHmmg9s/+IT07MZ8yTVLyDM01KeNPlNs40/u6X9QqyCdEt/Pq7o2XF/GUfMyKX8
r+YO471dYvi8wrog+QCpIfhfIVk6Khz6Eja4QcCIdyyiDq/pY+o5Kc9U7HFh6R2U
TYWEywpIqEVWvx8EeJoY15lTCaid+uTiAw4vHNiTKVlDmpqdx46BMu1i9gaN1zXq
WotyxoR18sGcjt3snlEQ7X2CMy1KGib8aRjiSllp1gHR703w8/f6ohZdUbRirRYE
bpaQkDJZtgqraHW0RUgDWpgrqsAp/g//M6m1P6mAm9/5KN4Bhk/aSUXNq8M0zGk4
R78PdUupVYctTCKIO7hQpvViPQXdvsI2za3Ss9ZOjC69M1GQxX1CiheQpGamd0Nf
PFNsPl+3iYFfcOH4Ml8pVNU6z6gU5i8td+mDPAyG5qbxH6FOkQqGdfcPRkTBqi+w
RMyBCRsjrawik7cDpFoqNu3R2KCQjYW30m82Dm2L3yFY0eMQf1T80ugEdgxRdq2g
FYPkA6UzY2V8MsDOoj3ZCFmGMfDP89Ct4TP0tgTEYnfkpqQpC5u0ZIT+IT2BpI6z
p8Woe6tTBae4/8mT7py23BLm+d8+Su9Jxdk8c3mYdDYC32Pw13+tlNSD9nVxRpdf
dGAqzzjXO2Wl2iMugTzomlO/FqTemCKX7KznCAWl82a+Gs+Nyj/GP+QqdjC1QI2T
2OTnNMGe6pHJaeaSNhSsqwPnPoWeDTTMftz+pIgbkG7wNssJSaF5bB5Te+GlVAWy
MBdQhOmrp4EvT4XoZt2D2/lbOuT2R3fsfDc/bmCjy55nMK35dHi4hlutyFX6Uz51
wzfFDsh43L/BRFblkUXmqQUZE4mj81t81rxepzPiaj003xDG7ZnyEg18L7Q6ZZzL
EFEsjvn5x42lQ4ZubvsvnogG2+UWTsIEWkTNM2KkXYvz3+dIhlLOn64DRMUJobnM
qG+jB8bW1TEtp/1mqmTcYIXNKDQqiplgQh5A3AGHoGZ/0jdQhsE2Mpy/xbyyE2C4
CYU68nnxlFBlHmXHeUIxvp3cx82jp8AjimAHLV3mgImjv85eMSEiUk8MCnfGVdb5
UDAsEpaxK4IZ18M02iKvCEseRYCNMJkCI4V6NX0mxIqtxVDMGyl19fZowl9B3MNF
pjlMF46vaBMq7JK5b3LfFyBP1j7rinO/eIfyE2rNXeIQCZwtNV3Sp9ejGBPMDLrp
F0Sxfyu3uNtHAf3zuf6g/gk6IhHTxXoi1BOCSeS2ijTB8jopH3sXSPDka5oXXz17
BmJEhNHp1+Gbp2xnFQOZLuCvb+rUU11E3Gsyl43kXHjYPsVGHQrssUYKA8wxItmn
/Uy28E/9+VVlr+Gual7EH7c+I19A2x7CY4JiPgU7w5YbsZLue6e+g4XA10Th+MKa
X+qUIlGZpQTedts+zpH+fYgBC1CaYZst41lWkLLbYpSnljDPOYPdXPVgV4RSBJVH
qyH87cIz1fioGDZeYNYHzj0DEXj764SMlgn2A39KSV3J+cg1HmwCslHhKF0Vb67u
knfhK0hNNfmeleQBsCJre3ga6pwgXUudztSjwhnT94XYlBl0+xHwWRK8SjxHBAL9
4W7IlsmHxih+rL8We8lD4QlvXsaNlKUy7Z45/DYJQavKUJBecBaogq756m4YSKaJ
GJg5nTPZblV/xFsuOV+h1tFHoEuk86ci79zUi57snKAXrlrTxCnCVOuueiJp+fLd
Kb93AaGhdsBGYFL8qzC1xjtM3WS9XTnGdcQZ7h9bcszp0w3ewmHwETENKpcVEkXn
70cVhu9Z5UlZs7LGngLYxhE/srbDA7/1gnt6kHqt6EXADaSvJbF5yVjMbpgEqaP7
jReFK/4+iD1Qi3GMiI2mlb4YMNNaQVESJKqNTCekpEAmquHWhV96Bb5wjZxk4ytY
1dEbAosRbMjaFFWCl3KajK1/aXGpBGGy4Y+DyzPvD3rsiIbht1NGQiSKofMRlOL9
TomdmE98xFbOdttkB472OaBI86Jl6DeGYoEunEMUHtpy8JT7oHno+fR8mXn4A5ll
oHOh216Yfa9k7RGgmdDR2l1dZnU185Jmvvfb5xJUMG+zHrQCKtkmHqb2jeIjjTIK
3dzeXBkpFJh6r6LDBOqZ4l6aFVCBLMuc4qR2u3XRY/RFeNEiXLWhRRwx8UVREWBb
iIu0vmpGmk5AAvtBSL6EjJUYucsZsTUUA7pOBmHOWrRBMjXIkGSoitdKEOsv7ecF
miPetBgQwU4aKxFmS3JUErAS/s80j1hj5DkZqJ7VOsEUdqiczVeqCzufHzO1k9sR
dhRjPD4roWd8HopheU4s5g0dn3ZdAAb9wyFJP7vq+w82YZVjRe3q38VclSF45Esc
bK05CJ2+slfm5gyzmINB0Neri04c8ZHX61vcMj3+Q7A2lMeEJI0GY2hKSMqTbqg3
oDZOND9MMTKqOUfTdaSoJw3fwmZNeK1PAdAaHWEmBRxmoV9KkSQ0ZpgNKH+MYR+i
oY+wQjIUr5x2lGT9gdZ31URVzwgAlT/H/6JC35JOs6rroPURhZZUQis28skhv7Uv
0FzpGYBuSwB9DU9ua7SuvdL/uuANalQmb6Gg4AjslwGsFwsPt2w5kcyfvBNl5/ZN
p7xqXytG0s9D4XF8rBWsEP5aZ2LUnQpp25NA3QTDqyB33jAF+NxwWnWKtE6yvXga
tjnu16aQz48cix5vXdhxu67GHHuUlTHFhL7K6jIRsZgyFAeU1j7bifxS0SufR6p9
oz+nSvSnO0Yo239U7EtLjjpAGF4kvP8adqhEiVQM0EqoZcUCQz/zuzzZ6fPOA9Tz
HcbsGd8kBsVUifNQdYxegqSNxUEY/1C5H8HD8uL0jtO95/8339qj9qgZ+9j2fZk+
ZbpvuiAkNDXoIFD9ezFYZPZvInRIWBGrF0DZcYXn7XHuFaNIfYdgFq/DXhlL4f3i
hZRur36fNU3VcfHtgIYChnC74Il/UjakNcDy0PelPdfE7yLet+UyVC1WOsyXcjVw
kbjF24TUhVXqbdnRYA5gpF05GKP63coaBTFJE6kHv3C1Z7kx/uN0cg3RusNiXe9y
9eAeLp6+3P8y+lN8Vv1SFEd1jBzlyqMaLgUWWIKC2B8WgVOJjwZDEseyayxRgQTf
3X2g9Z0FL18Bw2Y5/T/vjxMCPSe/InzXmIgw5+S6ggSoEzLVxJphXuCaHeoYWpYL
SqVRcy5WKHBb86GzFqmGrFPNgtaBvtoM+xRuOJWVUK2DCH1Z7UfTHhaeCCctMYtZ
v6WAPUwaX59hk6Gb6g7rcUUuYcQgtVZYOY0t96x69plociLPaMrAbGVAZbJG3rMW
PeiR8+efBCZMZOyfa0c88zuuuYmW9WhFZtH+osTM6CwQoKacuNEX4PCu+rLlPfi6
UQnWHY6vpoGz8g0G2vOaWLUK2DKA++YGuFKOL8w/cVSk0h+15BsTkTnR2tHMjzGt
zTpBiXJ1lI/S8vDhnxJBmZcMPDIV9wXPduvcHT0yxwFERDyyp/OMUOtS+NJVMXPu
ka0YCPrWscyqckE7ztacINI+0QEEq2aDc3lonufuxRANFCEGYyq1B9KhQVAeF2gT
q4K+SOE0xDgOQSmzl+oZlgl3ErzlbqHALw1wsvizmN1Jd6qUF+ra3ZYdW7iskV82
Jg9qkZDrykQO8I/Kb7IRQmz6dzyBhshtyzbbWwaeiDw4U6RBl0IXaPwLYNO9iJFa
P/iyhzzkPW4GFcIOG5yxC3SRNLx19oAn0yp/KwPetxNQ0MMCcWrxyBdDTB0dwmJ/
tyDojHaqtoeJU4F7elZef2LjTyBqlOLkT2FrzH6RhOBcPVMy7/t4fqPg0M4qzSNn
EjuTDThQsazcndB9BQ4eppB/iZYBU1hqHKDcLTV7dQLS+MoKXMUm+eGPkDTqPSZi
7chTmoKkf0qBtBw3+DTx9U9bsaHeh2enRaq1J4zc20Rd2nOE7Wc4JstPmvvrdIGf
GsZUwTEJa3D+Wkmil/v60S8yYxuKHRCBRUO59/KkpZuXhbLCP6xxM2MaJXYaXo6n
n9jWuq3NvvogDQBnsBra8Obusr5kHby0WdU+NXWYsvKx3070mpni8cg02jT6EAGy
x36oSngGivwoa1oXwbwKkGC3V+vlPEP3TkXeGwXMyUKYRxMARIqLBll/e+oatZHg
d5olOZn1UepwiRGJpvnMtT8ce39cIKqKj2M6a5BKYbIo6EjrxF3GdtPSbxA39Ldm
TlByYA0Nb8ntLdRissouYlP8BIhFVNM6PjOUzghntEexsYZ3khh3poyw5U7sGo7T
NuK7C0oryuGWvrOE1/sj5maUqGogzAXP7UCjovqqvQXHG+ZEUr9j9iv9JAClFA+W
saQ5Jhq0E69BR8QVxp0Yelt9+E5+IMEjvB6QwcuYpF+6GIensCo+1VSVSDv95faG
mq7MWtJ5c6T9xfQWLtvZph4lgKp7DQBNUtyNyroROMHsdr2lfMSf28o2EsrZF/+B
kqipYeXWfpytxSnQqAOXBFfIhkB8Y3upa75GlyCj8KKlpV9iNDeWKTFbigOfNdsd
pnQIyDMosamcd8iKn1szXo/JhQSf2XqgrgfyYvCqOdcDkZutKIUy1fVyfPvlYE/t
nCKeadbNKUQG0hdYQZ1h+rTD3GhI0E4cmECZJ2z2gXdiS9/NFLYKNshU37j38N8H
tg8sqL6Tkn4SM1DKGcHsmEfJPc1I5f6DbxzIi5qqxGlrYzFW9GDOe+gOAVQcDbcK
voutueIue73PMpWXTaSfsSi0IlV47dUSBGLkDbYP4JdGVgp3KjhJc+Qsw9lBCV1d
FCGeHD8qhVAg3JuFNnbdUKy6opyUqrOn5t1K0PIgGgZrX5uYsE2UNOFTksr4FePj
R9CK0HMU1WlYJ3+wMx8pYAr9PfooW7yHnH2x3zx+0ZlBLshNCxowI0zNfZYhjN64
UNC+F/7OU7ap6Wg8U+SJSwZ0xWdXznPrRdcVxhs55XksYRx0wUuQG4sL3biaLvyM
moSNAM1sMI7OH4T/CmCNMxuJZQr7L2OxgqUd6Q9eUy1HLkmBzrNUtMwpDmjTqi4s
corg84PbSVXK7Y74HF9P+UugYFTLoWcwBkomHJxHx/gSbx/RSNK25h87kGhfhmP+
yMdM2N3MI8mNtLueCsaIrtzChTT4dEVvpyDNj/iW1Ni6maWbC6fKIi7KtMoZs4ML
vY6qbde00dJsqDgdQUH6JoLA8E63XlM4y1MVcrdNXRqdFNlDKPlMSAS76mWNtI9m
dzE7VmhuncQYwm9Rkrk6cSr3/WOFX/NR84BOwOf+LR0+l6NtSpK08L5Pl1rBwidV
uVQmZmryQ/XXmu0nvoDkpwxMj1Ihj1D9lI0R0mKJnPn7Yn6y2KseL4yt8JSFpcYv
b3p8ZUL3N4wr9qT5xc3JDEXkus5T4nJbkQbCoj7Qzl/9NF1f0DuqjoWrBjxU8ioB
CXulnkeEDLg93arZBk+iS+/9N5jxUNqUtAtXp8IWQY/pph6UbEN9K1TC28NSEvP6
vot0WfZFeh1mPrNVmdYYkbzNwYOZNjIUVTvNTOYUQNkzjXCtsVP9R0Y/Ktro5PGu
ROOYN3t/UInGh77DmEWPXpqXykL7JwWybh9mfp0XYCxiWbQPcDSAhWFhHE2xFCyj
pibJJBfbwnSRd7GdcTHKup+EN82OME4a5kSVLweBYBqS+amW4hpavwzRn5qANL96
PHsxwoC68hcr4CI5p5eD8Wo92zlgUe1kMCyjKu9NchPtWHbVAVQ5dk6rPiGTaJhD
sxxeStt9db+eCZ+ZPxYzGpRipBBuUrYn6SCEAupAQnQ+gtfiRNfp20wNAqhl8llq
9hkNIuNHNWqBu+ZXCohwn1v7hR3A2GGUQOENRzJuuFQzNg9MD+tUURx6FfbSqZkw
Xr9iCRvsRXBL/I5vKP8Ur+y+tFUC0kZKgCpiiBHZGP59vDj0BCuCsoWCgQqd0uV8
j+lZRkM3ZOi0uUFzOKB2bvNoyNUIPwnUaYGBiTi7+ReIo9HBoRRHZq5g530yJ0hc
4PLRqmb76ZZpVvrulOyso41fWRdua4zl1qatHHw9by+0ODcnAwt6jVJM8d+VOv7q
AlhVISCWOM1VnAN80nBUyo20DcIludHNBbAO7uBGCfeRBydAqpmTM7WS0KJQr44f
vwcOMgsVO1N5IsFiDKBOo6pJRAoZGCg5ZW99o+CyteuoJfV5vdZPuJ5GvCoOe9Hq
9S7V3b2zxCt8oLa/TRhxKd3aar/caisOrIFjCjStZpH3wgvtypRHOAdtuMyzROr7
0MD1nObiTJoJh+cXFkZVS31SGX565LR+r+SpSWnTQNPO8VwBVMyfY//5DHYpUpZk
/uO9FV4I/cQ+/8EMAUjzck/mrSqJXZrxTk6emjE4iYxRg+u3BW6G9xF8nV74/bWh
VTN7WG/vpi7oCkVO0LfmGoaSrQmM2LmDf9H9yaPQA2rMCqqp+hLShv1msozpbYFq
pdDS8w+C2aPZMPTChaeLLEH0iVJIqKa6cPiN9+dXCMTzNipA/bAs1w+ynDZ8gklr
X/CBMyd+Omy6oR75h+fe7pLa/N1vPJCTh2vK07dXyxfNDvqv2W2afkTt/jAjbZkl
nCssod7nvqIRvdlAfd2EeuTex7P7d9zl45Kvm8wJfC/r2T77sV5newzLsEfsbccK
SUtoC7r0CLQg9tcnbPArW0wOmnokfREzUsnuuLLeQBXuky2mEckq+TBLFQbyEHf+
19ZEvFp0NKKghkdSJah21N1W7k08aCbrU9CdHmDaJ3EakQdKPtjdhnYqfxztET02
l9AZY1ew+0SHnZC2E87ytvIQBs2r0YwpOCi+j+UMn1W+w7k9we5B+aeUr06DqXmT
s5CRqe0vYoU+I2WEG9YsHwI79zGaTSJjFNVYJl5QXraKFaBufXo8ybtX8usQ7tKE
ZHzDMLSYVu8va/DaZQToOILfS9qrBKVnVAktYRW2iuMb0N+G99mIkNCULPtDwGJE
U7bqYZnVZGHmauTaMAldSX1r/kjlElTZDlx7jUAmE8jfXQLZPFYw/hHrg8pLskc3
8cxF50Ii4Z7BOr4nTylMh3t08vH4nIxURMzlPXn8a6A1cMwXh2SaShV2KuZW8HqY
9EdSV32eJXO14c9uaSIH/kh8wgBGgdQQPhD5cB9khhToRAaZM1XiEYKFJrxIr7iK
QbMDAYSNS5DDuiJocdwknCG45UoDFMsK2gaLglhDWsDG2E/mK4hCOQCp9e9Ok9LZ
8RBJApMfGGuL4nak+wdlWHvzI20LEZN/eQJ3ebWSyU98VEOeXFUqwDsMaT2Fe9yQ
XKt7QLcG0FjgS4+BStqQoNcIzV2+mOOtCVmtYk4EJtrWLHkMuTrdEwtspE0t7+Tm
gHAaDA5+bg7HyhQcRx5QBdQE97en1mBLvIhlgdsDXE7WoOSXiu2EFX80gy+GFvwd
63yLz+C+Nca3UnJYpspxHWwjP1K7CyIvbJj/FbUY7cS1C8kksg8k/Q+ucOEPtVFi
0jKMEmXXFedmPT1QK6WDfcbi2GTeBqCaW1B2dMae8ou2kLA7upQ/xCftCsKERhcN
IXWA0zKmiHQjXFeTltrMsf7TyFlsTWrC9IyYo8KtBoIB4rewQRnTDrsakMOYhyxS
bQACfvxe6iUmGYZ/2XWDN4ZB1MNbFQIvio0qJdCVQStlGMMiWiMkjUOlVRn+2h2P
cu+MjcwTQKZDQK8N2/8ndQbq/Nr6jvqu6lY+JJZEAsX/9wP6hMz37wjwNRPhOH0u
yktp533BTzGBi32QitIN3WC2S7ztJpOlHqY/imCgSgdew2i/SSYD4dA6O0XcfmKK
Sl4EFa/SJC5XJtQZrofrVEz2VhkwuLKxDEO06NIk7jUic0WvSDQaPl27HBcbG4Ly
4sjzPOA7ZnhuS5E57mxhzKpezxI+5znpKxItz5ixw2Iab6Ax1qoDfKsiJqBYTUnt
w01CefSGJ+hE68FbYf1TJvaooa8mU8802C7VOA/uVTdiPS80vbWevhR8ZqNg/Gro
B/0UOgEGxEpKNmQOiBdakfU4ywdsQLMxis1RfDzlA268XenxjHCkMKolkJAEf67q
oWcRMplvGQ1uG5V9Wj1i4S8yWz9N+1y1gyznMH9hpQzfd8LBMmo1OC9mFl0iuMfz
lB3oNsh9qzv74nfZ3FCQ8XjsaerdD+08EIKVH/ioizCqkHq9u/+1R1cTX4ycxhmB
3r4SiYH+XyfnPCMfkADYSEyUPvGznUHg3qUKcc36MUBjqMAC5wW+g1+tepaDsuYa
1+FgJb9znZlr5HVQa269rrSThNKHYymwcXSuOp3v5iA+sz8lptMahE1R3mer46N0
+cM/zgKEIL8wrxVh2annuq7ttDwi7Bg1G7yL1lXgaDRNDxpJ3/PttS+Uq9KlPJDR
mzG9dQY+NtB9gg0Afz+Kwe0kxYj8LFnqWww0bmG6yKZh5UPZbqqIF/lpIdS3Bbo/
BKokrvGyr3IGeT3WsNvUQe59P7EqaHe9Z6S2J2tZ2uK7DMFsrB3Ykt99UIlSL7o1
m/vLpJfQ5GiTMYR/mWyeR8tSzfv00UPwZIuQAqX3k4zcuCt7UC5QMOCV++auKtw3
4siHk+IkbA0M0SNcZRbaUri5YiicL9/YEUJpX8qIpERfLCEPxVvlw9Q8Axh9oQ2q
OL76hRamDsElGXfvtJ69gWVDbH749aAA0c9AGS6xgANPBjACQFAUw1Qnas1Ggr1T
8oQrsX+1+3bG/VPRfPIIhZKK6Iill7dNTsMHkW2whGf/nnq4rhvkWylWDNfy53EP
cAkU5pbTCcYmOnccp4b303ebml014lxDJY8jFwjFzv7DwtxLHI2+3L3iAE/LgQA8
6cv22SSy3EhJHSejgWraCOwF7kNjtFSW/OUDJtHch7+6R1x1ldoPyl+eE/n+9Xm8
3S3UvSs4RQ6bOKhspAEsPxLi1Vv9FdXhUCe0M8sTFA0q3W7+Lb+tjRU66eRj3OzR
eZGzkJg1gux7dGoO4+fHa3y1DokxVrCiv5N3qu3QZXq8RcLqozO72unhqPFwV8xd
dZZK3TS1YB/W9coWrwGF3jBvX+aoCc1hwpikS3WQ05j60FomZJkRSHBh6uyVowmz
MRzqXtmK1eLrPzBHY8bTZ5oSE1dY2nEmrq/o2w4oDKsC8UY8HrumIbJOq4B35/D2
mY50TzNCbzyOt9UurQK89vdyp8wNhtnX2CzGNtZ1Y5kv+7oBDG7KxVa6NaB5ADIO
mkYnfv9hb2xRXRgEyKYr2D4HrLgBTeTrQyIvetYkSXRnvrl7DfOrxvXMz/dzT402
Xji1v/UMn824qs6GHJTBGQURvMMVmjh7LzvPK82g7Z3g8ft34uPMfonKIrHUZTYf
sXp4Ocw7T66qHjcMkTAxffXXlA4Rs4u/PXF4k0/QClXRRktHFKVtkCg1jPIBgZKW
NIM67NKpkmdAzd502atXVUsNCQYpHDXNE0CKsrFTxLJagaKx/fYjdYKqSfL6vdZW
XMbUvFSRmdT/NzkQo3MeyfjD9i4eYC3QV3lpLwywfwyFZOr3I8W19MH51d5T14nC
NcS358+a3MoOSN9o+EVxM+nzdbBXJnn11C5o7aOoBi//mGlY2+JTck//xIDMzKP9
SaMs+4Nw3x5rYjjiqDXAB4T+fTAujWuASfsoHbBwqH9XcLcsdXi/6pyZlOARJoEK
Sf8/pJCoZv4h9YtF+Idf9OR940uVotyY6Rf/Wrzyeu8XwPI888UXKXJbXwEBce60
kgJDPu/YRPmkxGtaXg8b5Z8aGCDQO99RSXj0IJt4AOOO5+kZccM/xLj15tqEltqZ
ueBBdtOegSZsGufXyYyRa06cb+6wIMh+JAEjKoP9ccOkI4/MZmopP6IoWpPoVq/t
txPUs91AW6Xe+WjS1R3uDwtV6g0C09AfiOW7HfGtgH+zjmMJpPCFsnFUgevFmDj6
Z8x07o0I//8Ai36otinpv4TNGZdHnkP/08QXWRsnGtjhj2tRSMO1Fj6lV6QjhBty
R+RgkSmuvhbeIHBNeqkbKFZCEeL4GpYs9CkJ/krR4rN6u6D/dN0gfqOd7jjaGpOk
NlVg2I2825UaByHnpJclIyoYH+izrf5qveAsRD4dw2WWHCqpIk2wZNY5WgBlrTKE
TLDBMmL2D0glEBpEg9ruBoPH/6Ly61xdrc9liiS+MJZuOorT2/6FtfTqOl04NnQ2
vwEAQgMHJZQN+0v1SkHTl6CsQbdacpZb+P2p3USfamADs7Q2yuYPlMgbtPNkc8ip
Z+Vvmw3s2nar7H3ki/UG0SLmM6cZlsaYS6fGqFCA6UIGj7AV4P6PoQgSV8stwTeJ
a1OQM5lPVS8sXRK+ugQjfzWZBCFvMUA5FDrBSyRvk9Qs9IdDd62/yf605L6ETjhn
i0nkp/vRM/FK76V06b1UF5OENBGjkS3CTNbm19IdaEgXirxxtk2rkjuq0Ux9lFzX
HATcx3GVVtfVXgPM2h91qnWfcsbk4297x1HdAPevSmej1nS1EhIL1sU1UzvkvB+g
iRrOg8AgOOdZbCES8cWtZP5F0g4JyIabLucCwzkYDp5w+5iNaAhzVwQD4WnfLyC5
WWfO/G2sU0Lpurt3rPyTX+PttCmjnSfNA5sMfxxMtK6C7EzsqqNJ8ZUTTxxIP3yO
aks3qp+xrNYDWcJNXuMn1vgl8ln7seY5RAkJTU8VeGiu0giw2k/PENF8nbLHqN+M
e1VjdJezZ5NNfoe8KDGBFCF39W6st21Xb5DwkLJnyLUbgbBqb55BdJQbKGnSL3pp
l3JdoHWsQh83Zome4SpNVUGNekz3aB5bBEYGXWVyMzWnJSub/f776qlrQP1Mitqg
hYaDSxFKKpM2UVpapXKLh3Zt4iwwn4Kx+G7VCiSv84dU3kDhKRgq5yDavXpU7kLz
9mohiLji60ytQMx02GaF788e2uyvcTVksRu79bKA1H2XhGvVrLOsPmTAgPy4Baeg
/LYT2v9xzVxrXUcpA1nY6DPbDvXWTb8/UUEGWsx3pAWRFjvMpfxR/22rJKOFrojn
JhbjR0yZP8SC9qoRleq/YbZFa3G1QW2iXt5X8LAeIqHS8228VGY3zASrK9QagR14
z9Z8B26Dx5BM1MIbDj7Qh81czTwy2+Xg+4tbiyw5GI7YhCwrmEd4nWt1fMor43ls
9nwoa+yAxX5CMRTSiZOtGJ+bGNndUjwKQSiwX62XjFvRZQQExbANVnHA6Jq4YrhH
yCvFQSjgPV7Cqre3CaJgZptekf1zcgghzCvagkQcSWNbg2eF2wgHpjYQT8XMxj/A
x/KSBqR6j4c20xf1TKJf9kTs53krMUc7ObzKWcfBNXubnTBNm66NAamWxXQ8MzMW
ETrtiKLbjolOs9L3m6VYKNeTiOVy6Ov5cPWDB01dHhGicvy++aaGAR83Fb88BF8f
uEC+jMzICniFAp4PB1EjJN1GQctAGI5UU71iA1IpEPYnliNRbpcoiLRkLyACaEOB
mk/sVydWY8pOkoBqqyHruqIe3vonHG7rsKhM9CtvDJ9ldO8q7HzedHL5UZ0swZRu
qjSUJDKfj3/vLo2FTAlDyR5n6E2GwGZU+MW+jUnyh1aoLTsOKWOlgg+5f5OHLlyf
ovHRvyF1nVnqqlKkI2pZxXyH9uzQR33u65jb7KMsQqp2azsYVVaqsibpHIEfO0a6
7w90rqaf5pdiBMNOo8lyu/NnmXPE2Giad+4vUnptCJp2RqlpszqacjqHsXVbeSON
+UMjtbnnaiLvhZ9C1ggdamV4ToTeS/B0e0pjqhxngWGQPTb33oZ/u7tBDVTn9dxB
8hI7R4UKH26mxhJJvWzA7K4n+FT8FhkSNQBzDh3mDSC71GoWq/5CmsgwGTKldrlB
tMC7R4cNk2kUXlMdbLtbvZi8Q5rhHA2e0itPD7qQRFjlSjIerzCHUyArvKW/Et4w
f+Tlv++0doRJYLVkby8V4pHQuZwPaHHrEjJBvAiHqyzNDWo+kPYnhgkDg2JlA4fg
PT+ERP47unOv/FisAn0ZQOCP0fkafBlfVzu/qjiOKb4pUU9otdIlbYCvdWZi+3JL
iPSp5xnPvnaX2mejNe3EF+WUQhp2Yj27rr0upec+6MkZJekrJrNbxZpq347DXHTO
2XiubSqyiesTuJSueigBYTRVs2fY1/BaKMy1XWkF55Ogb/gZIXoc9AwXmz4bafbZ
RYikTrws9KhiKeJHCTX7YIen1r6JBhzIZD2gicamRY0wC7Pv5s3sopgfvY9gn54N
OeQtuzfd8ds0kcCSilPIPrb5DLI9wBRGNbhgOVRAMRcZdP0QNFqa+G6Muce8Mr8a
ixlFJBeYluWIPUf6Mxns+7yxn/VZ3FxLV64LS3eHOtSGCoXQRFWai2FboES0JY0+
7qDGSpBUrK/jApkefHZZTsmG6ddWNoHs9RkkOsBR1wOG5lvEAlcvJ7XcNr9KcTgW
my4ErvYHptviCnNBy6vFmgwoOuSFRzNSOdPJAijFgYQApLDghLRIRWuyDeRYvm5S
PNEyAHjf5Tz6t7RqGVZTHhz8d3IM2TkFTUn8yducBieiO4MD0iwDX1ApkAmQGZ4M
tKZQwdZ61eLkG1ze9iKOcFMC4fsdcLSZrrNJsbsWVZRfLYIHGBkqDPed84Rvmjee
IA0wS2WAhR2XukzgAd9+oaR0LNjSP/YEIwvkjM9NCpglxPyw7vRw2gcwExAGZni6
58MguOPNtj+0An3hpO5VJ5HoH2GyoD1b5ckHcBTpcmOGCfu6xUZPzcPChguTdqyo
yxP1yhzURZ2aTyLpS/YpSfQJx/DYUQYK1PM3TP2XWpPl2mhZkbHrmNE9T1/MOGsE
uq4Bqdw0o/RnaV0i4ijxfG7/8VU1sEadcXnUSwqbruc+gBRpAepQxqsrZp3jfs3f
42imW4GZ8U9mOw9JhGdRbbtj632NLoP583vW1kRmvmEr0e3HIFGSBeIRCZKIEaWL
EEHDnwrqcKHqd4eENV3AeFJjI+K5NtSdqP4vLPRyGo950lsdnxT8AmRb2bu9VyZv
nR6Za+VzBSHilvssDUdHC0dDl7AfqVc1uyScEY628VqQZduEDZQrRST3cIXaLEHX
CvyzJDkGTZcAK5lcl30uiU30ICEXx0T8935LZuWoMEZdrqO2392l43Ik6xHrKleW
zLUhFTWshW6TUsdvVwjTmN5+ALGY/ku1Y5SFSMBfHqMywSqf2QONQ6O7Rm2XWXAc
ZPlP4s6R5ZgVbaFS/fwCiGO1sFvvDGF/2DinAod393Y18YaqrKZNPitrL27VJxXL
P0gQdg+vmpJaIO+g+xvdAz2SYNBg+AeG605LRolq7f97HjcxtWjFG2UHL2HLHCJo
1dScvy49kOYMtYKqDEyfYqQmq9kfIh/wm98HF1dufrWY6FM7I9qOEhkbLcwRF3Kl
ffNkMiotDEzmfLSWcdhC7ZPzBThuqysZAaKIyDCML0xl/YtVblO699YvCOI96gHJ
zOYtwc3SWXsO2vepbdT5L3xDeO1WF6GExVmwqKUpnmtNgjkOR7S1AbC7UornW1fF
AyfR6dqpFH0xL6Je9HyRR95lKGUT7dJCKKAEGsXPOTBRCIIGqdPLfER/PWZ/KSdX
MWY6HVyHC/0XPawcZ2mNmq1rGZmgoGSI09xLyND0MQ04FnK9+XaRyEU4OWE958wc
oIt0pVFRS0QOV4uf80AGyJeS8OA5fbtA6b/4TlrjwPLE8ToLiE1W4DIDqDtavX7h
84nzslzEMEAH6PIAaRAFaWBXaLcJTkETSvoHO1qckRP/X6pAE3pYrcMXx4Qq7xM7
STJhcy5Jl6gYYOl9Msdh9PvHPMly4DyFwYt0IVJyhHT9M58sCy2oNE9FIhwhqqBk
9BV2c5xywgv0yedv2oJjoylmRK9KVciqFQDBxClsVjHxeTclisse43squ+vyoekV
ZyJoDrOiiQxLROje4HOYhVM5QAqynnhEoMJjvOjWGaRzuuWOvg2V3V48W/YS/ovW
AitgY/qFk0Y4zvwYgAk/o8R9PHcLfWZcsmhsUIUfbxkfIs/U7PrqWNOv1rokzrrc
uSUgARIGbYNQShToKfZI570WHvWYQr/cnqfx5B3fvP/YB158M/+zr9KLDOcCC2u9
00sF1Wpz1ccB2Aza53GUPKvhRIsJk9Y24PD/HUh8bYFwVw3Ip8FRPc8MZN54KHCG
ZcHhsfi9Ze4MSD2hiRcDlE1gc7dAFCHoMIrTVJu/drKNNxbDemaZ9QK+9tXgAlMF
jHs0xZrqqnoOZAwKzMBS3z/iBHLgJHFRIcobpzfMuKKzxjawUkjK07z7AgiHWIf+
WLO3brrpToJt5LcHy2lM4UekbikPS+uVIoUeGwa+bp6XiIXvuDWrOkg6ax9y31d8
BU1AToCNvS9pjlLg9EqLAsC97/2dClPSy2cK5ELcBc/tzhi5EHhf7wKG5LIYLObZ
u0JJ7TM0mG2du+Wbxf6OUno81L7r64Pi/YROXOqTGBxVluqZq/iVGkdpBbG5Csm5
6c38zddw9cBtyoeduieRfaVHWw3Gd3bEUCXrynz1SXInq6degR9pc5j2bDTwIcMh
Z8Vwt4WObe4ZC+qVXXObSlaFlW+DYZCubl3cxl3L8E27zGuAAG65uRIcKjfimSXm
HkRv3KH1LxTmnCoVOilNtBPDy2avDlpqF5oXml6y1NLdLVQSKjXYxm1xnNm+aPZY
JtYl35BVSgPIGUx1yp4/zoGwYb0CE2PxYwvxAIp1cu7TKRWdO05w1frpPKFb0/w4
RRzRss6qSRwCvOVklreQRdnI0v0oxE7leEIUk23UvwPQbMwZx8dvp6WbRVrp48U4
CwfvhwzBvGN8qlfJDRVI5+QvFzL8la3iukVhUIcWymQidc2D9SSgHVs654U7xI1F
lEKzfPkhrXcadaHfK/6B3rrSnvgzz9KSw9GitYOm3zqLHpsbikhM5F0KD1n8TYKe
UvCH6950e+t9i9mFY2Pbrp8ZfZQ++4Rxq8QdR09BeWpbvs/AnRBh33HDldeh6/5c
6C7prnaDQFKvwaOmld/9Y5kn14NiG0vUS3aL4am7IogTvhPbcQTpY+4FJmfdEhLd
B/80Zakd93zz4+UGBLO8flcH8zmstS9iYpap6DH9AsVmcAWf60/YpxFe8yMlnVOK
4KJTMC0+AG2K4HMHumnzZNdZHMKbXMJBo88pMLFipbCEwYEA6LnXs37UXbHyOqE/
uuYrFTOM8cXuff6Dfmg1ZdQtWuxm1MNG8fqLL4yrTMrIRGHWjAOQRcunop31DOfd
PP87jUzzpktyYQGzC9feibIacJJJPBgaNxpTFyNG4BuyHL01fOnuI1wyp7M/w+t1
H4eDlgV947OTnXAC0aWwRg7TXjf1l4PhGE3uqhuvzruXMEKE0jlbT/VRNfliyHDJ
17//L+ob+h4xhdjCYpdsyVFMj6yqlqTsDjVTkTr5H24c1h0h3dKHYQCAanYndh+c
nhkJ2PkXJXIwwm/WC5N/GwsE9HRcirW1cQDxUYlkYjoi69b+gUUx0D/UCQLmMXez
D4PWvn3/tq8es9hIItbGXTtFzPR9+nPmEhixnh0CarQc9VC+FWAbleo8d0IntCpU
isU95c7Q6T52zN0WkVfBEOZqmRm0Pgg/mGBiWZQFPWwySBEndDrJtMT9cy8T0bkz
Pa2eka4dhjrKyvaOqBRmuzSQwN/6LmLGyObpjUVIYPuTqUgxXavZEL8zR/qnA/FX
BEGjOLDDqZnm467v8bDcjMFehse+SKE/TtEuzlxhwLTaGZZJSQ6sTNqBuh1cNBD8
J0NvblkXV14ohYKYGdy3XBSKxx3NLv/xT+CxGKZOT1hJlHK4NX2RHk+YmJx9jc4f
YBiTdTwThqyqISbnrwK2UAyoYGAcZDYra8R9uroLEdLLfsuxfhDSXhlKg72ZKMv4
zED/2ZWzoFd1l33AjTqm0beBSRTpN5HseXUSA58sk7BYClCMrj7p23r1ZMt8InoQ
v9tKMJcQBjwedF1m5wD1JCLxjWfPNGJrPJsxIXd3WQRlLKl74LP34YisP+cWXXVj
CcRMgm/tScDc4RDuspYE2XJwwMOsVn/JL068coWj1WJxx+bQMxNQhbZgBdFZnPlz
EgAyMtJba/4QutCilSTiEGGS8JgxTBH6RnntH9NenodzpQnKgvnXE/rlcgGUuaQi
psuQpgEbtoY3zVS+0u4uYAwujuMZk42yCd13JDcPFIBKviG+65FJD5YRC4ui6UQB
SLAFlaxAMOAujeSijNtzs7ZZqfjH7XDzYKgr6TZsGNuHBDb2pcjovTpAMUNzXmX9
M6PIqcKnD/OtVdAKTAgEsVBeieVMPpfWAkrqyRDNCtnqDdT1jS8Ac8tvTqZwIZIv
W8jS9Pak786Y8jbAkDlevYxByWZqw4g2auFZzh6cLtWMOQQ4AIuDiQp9pe4Nbksq
ChvvQ7GKCfoynRL+kE7yUaV+vNei1bfZFEbXGlS+w15Cs4fzge/VlQDVFFHOQBn2
vCZ1t2KbL8ytAt5CTcM/86jkltq4YxochtRk29Zq7pTRTfAkX9cwXskPvBSZ/PhC
usuQ5W79NTV2JNutdxLGEkE8jFFJrVagrxZqDsXKiXrHeecNhz/U9z5LYGj6nTkB
iRMNV8UurAw1gHq3QEL6bC+WP+x7rxFZcHjnAIYL2fOZVjC4RUdbzVrgyFfEFn/y
Apiywk/clmaseqyqSpK4QgJdrqTgNDC6IOX+F3Sg0EFfrJfQN0KMESS5wOP3hmsj
Q32aVCdE0bHDeZiTcJiSR6MZ9p+BUSBKH1mGFYXJmLge2tOZyErACIpMzRmL2PXA
3OarTdKGXk2jhudcblqcoIK7Gvu+CRX0mxHUEf8hPQZ90EB6OGldoIJDrJ4UKs58
Kgnxauz4KeK0nE9pvQ5/v90ILJfuVNdZWuVHMPt+hmZLF5y+GTV3LIRlNj8L3MWr
RrH/TjeW+m9grhhDKGofLfWQbsFSdiprA5Hpe/JOsYmYS34ZOZZVZXOiyHpWFso4
wMbKIhUzAEmmQYpXLl0Xsoc4wQz5JpgnQ0fPwYCEcrTDtlQNJLaJhCKuDHpGwdNC
rjn+7qgsjZTOuicOxsQ8X1I2/sTl0pDnNv//AVrEJqnWlmlP49XTYr1/fXuLoxo0
Ui6BTxMRiz8EwDSysf3j5Fc/Wpk8NMdSl0Wt8kjLiiPYlskPzqdnHZIMOa9ox89F
pJ/QcvUZ0XSbBWPvpxb/z+/lDhH4nfNeuxOeIBjTDeb8GP6g53SfkBu16p3FFnUs
UQjMVRItWAT/mQaimxsLmohCjjNjG3/Bx5nYgSEFwvo6OzzkMSsl5kI5gjqf7SU0
n6+dGUk7xkvZOHtQm+3PGL32VRJdZS2xSA6GPsbUEjqGPVdpxagceEG4nb38x2Pe
zchV9BOxaBxd94QgWC6Clvqs1TP5w/8yN2WvSGgmosIjlg3bRbVMVE6n7/JlnTb5
u/BmLiMh9FbhkA7YQWV6xf1jRaRdrdk/soQw71Nm292P/kgM3uhhF00Ty4Pv2Wyu
eFu2/FA/XEuW4VhLwBpzDURGV6/ULaFTqTYah/LcI9hpAOHUfYsxGZyq5l5PLNdb
qecKr9YkdQLoo+HxTlIbTdLTiPTs3OQPTE0Z6NWQxZxTH5rxgi1LoOVguCMhotyb
BgeooFj7DOOvsMmd9sLUCvrI/d6D3ozjzuLrqgeTrOiwDhaCxzhDLI7xbxTgvjdY
bJV7cCif1ynQz5UMNdoQd+k1uBT6wYKBVNSEpgtCiw6mqNW9a7lESXM2xHdsYyKd
CXBQUhepTR+TUGxiHcrkHHgvmrysFehZfFC1f/fLMZUj28SSFY0WbWtvUMEGU60w
tezkAWm2p8d0hFztm7RMK12wvkH1IPSeHa4dbTyK3oxB1CQW02iGUEv2Ip4U/HUJ
rSBpc7iDSzBTOSrfZ+yHP21pS2C0+xMJD08TpZVmd42LMpPHy5fZYybtzTbKoZ9L
qk4NWEctxHHKIyZAlydSQom65P8syHTIrVD9CaAoPOJ0mzxm7KTxESK8x1Ub9Kb9
6FUd1AwLDE5eFLsYGdzUnhvxKQm3vSgbq92V75tG5KDtiO4+SvVAHF8CrwxNJ0Xe
ApXiftW18BfCU8fA42YecyyFSjSfFr0N6c8H4WW/TDoL5oeYDSHZCDxFcYkmdsPu
V66BRIuqXkyZrd7+GM+dgE5PNMZskPq9k/5JwaX42nocYaXX8Hl/YAXj1WgH9G8d
51VMIs6LdYsTW1qNT/JX4y0Tmy4HHvLuY8Umz2kQ/fy3VjLY19pZYmJalIeQVDQD
AcL+OAJ+OAnmuhUin3QnkYD6oA0olGYPZvptmq/mRMIASdPKzo+NQM0GB8mr8Hhv
HqMRLfgaDJEnQfnl/iY2GsxyLsK79IlHf22jerI4DFhiRhd9kH9gXA+tWDLgoQWW
cA5CauDy5rs12GNnZNUVNCdSoe6pkwkneQorPk/pcN+yXYidAhyaVPg7uCA/FdJ2
Yhk1v8XVggsi2cvjHpBZgpo4B8xoWJxo0gTtaTHiPBbYWYVeXK8JpiDFEbU4JydX
dJ2BfwO4RziE9lc/16GE2uIqWBXoZcrwyWw8y4T+mi4OFfOW8JBl2W+J0OEfaIgD
hqZwH6bHqRAByMkz1ppSN9K+WxOWKBJyJfdClsJt5ZQqcgf60Ppkh0SaszVQDR81
wLdRMsmd3s2YJffSOdOpHDy9fsyDwz/iVXjFYpBLp6z9sZgfvIaBJnmN4rmuRI5M
Mncc4WgO+GMTb7wvEJiQmrC1a26bIuw+acLrCEFfOXSqL9Kh3PItwKpyXrLOKNKG
E2i64ub3kEUlJM0YI/zDwIZel0GBspq+WHdSIrZDtxAgNDuJWPtc3H3EfGkvFKnq
WTbxFfhNU669McvoDr4YZk44sPLoRKD2uOenXWbryHqclT/U89rcXhN57stycDSZ
Z2wj79Vbm9rLVFXGiEXg3hmDNIYEino12kn1eKyBuabnvhmeEzSJoYk7r5frWjMC
M4NktU1PIFk/oa/aIFPFNs/xydyIRPJcMfetOGcA+Hr7veOcAj66CugYhsUcyow5
26D8mQ6QYdcerCPEy/KUMGiZ8ghUMLg3qJjgHaaPw+k3NBInuAiPZbgC/JUJXHc+
CYiz1Pq7QdPrXoT3rNMN8TDqZtbiSZniUF2b3C+PNofVbxtnj6fDwXZFH+XeKPhh
bq2OnYsWpmJyj6tv3WUpvVVqKyUJQD5oQxsbBUR0MiWHasLaI0SZEKrGmE4kvkoa
1xN3aPEjX2oGYsWF9OJ0bRnsmBU4USb1xJrlyMFOpUtANq1RWHEsBI0oI9DoYFhN
n6Qer2EYfPw6nNbWDGdOF2n8gRkMCWifMMk+bLk462iYRtRltQbsmzyML/PMbFDS
HNrbj7MA5eEQpJgpczqlON0JZN82XMvvOq2GJ6QfHjbw9ih9HVTGU34F8FNVifJ9
UmMbQYM9FrpHRBL+7tHgKZ5JF/MiTj1TV/EPVehKs+0Facxmayn51ONxNzaaQTGd
6KymATl1+lnU8WYuIB1eEaX/INIDYxllPlRf32upYPyWGPxsak/pp7IbMqHNXoTq
UIj8r7JMozGVwmRtmdSi09yEwQhtiaugjWqUJehWd15SXUC/3xFBXi90WQqWJIIf
y4JHPEzhao50tOqdW9BGkTxYRw9kYDjWw9eRl5ku4ags80n6fSh3TsHRxK9UW0Wg
gRpA2kPamWDECVWFbYpcWfCpQ+yogT6Jev7dd9RSioxcESi2h5AEEqxqE+/oT2iF
JyQvm7kRkExQFdQIjYcZ0plUJzKE3KU6fTcTaCI3cFNfPp+LgDA6EaVT6529/oo/
GSBjEZ2HZa59qAcFPvCIf02YSZfj1e2iOLws22NSHTxkkZji2VGY6bjDB7ulj9Io
COTFDQ4/MvdySxz81tWdwPVAl0jVOlIbOzIPy2dUK0ShTrUpiCSTFh3v0RY2K+IN
+2n69L7ObusLmjJiacLKfykhfsqseUiay423G2zduViv/XgyUZfLfzxyq+MtBjIW
H+zTTyF3Nee07V2uAZDyna7L1N7CKslOeCQmDJcO6jKMrqk+dJI8WhM6af8gcOCu
J+XR1XQhhrV+xJ0HzZmwQcQnGS8wTDMItwQAZw3UCQS+65KAgPS+lC3dIayEwBar
vmmQFd6TFmK+I9g7r1Rg2DG5AWnCX8/r8oUJppXRFLYl8Gxm2ebHNPfLjtFoJgkU
rGxISaPBax1Oys0GI3SjdV9/svqrHvCNvRq/Vb/PRrzRKKWLt3LT2pxRZQM70BUe
VDgrtFOxtc7rMnHB/nyY6j0DgyqsjS/BkpmkyycbGYG2tJjztqNR963tWsZaBf1b
tcnokddD0xmjgPHXVIPxXVx44sWWtnh1xBk594YMJfYnaVgn+Xc96TYv8P6bhjrN
sOgNbeXHmm6eXxsLPeXso5+TuOLQrBflbYty/6DX7RG44kFlHsdpPv2/PfamIvlm
5WeT3yT5VlNBSjzbIy4pYDtTckwppvyVY4HGf48hO7QYOjm7mtit2BAhf+3oUjba
Af3EaI+jdzUtzEoF88EZy73kfN/JNgJed78dcTwlklPQR86GsPik42jrvGvvYJOX
ohQJkWyeY2v6ukCNcXSZ8ZXT4fg9lkCCzKw73dHR1ZH0vxVNQzMThZazOWQdfI8h
8AoTnuqZeI4EZIlWPlzrED2ROVnH1oO9oWaXKBm64RdiFq6ZLWiQ8n0jnrYh8fAD
l7t9shVZhxloih08U1Ry5sr/jscTcmbxKLmSbJaB2nIfrNMczb73y3RqDpLWrWTS
APkssMjoO7ffnMJx9MNnb7IZfF09q6TGLpN+5EbHalc6Bqmcyv8hqFVf5to0kO2t
ewm7QmQNpy83GzQNJ1QHHnmn13DW2txu8OTU4E9+gVXmtYIAIA7deE/SWt6nAuun
DTl5V8hUs779lsqi3FK9h6VIxh4hM/t4F003rFhnBwdTPmiR2Nn7iItj9fC69NM7
0Q1MW/bfBN63SEtVy3YPvVbIefZPBAnVeqT4xGe+uFcOKYsZR0dcQaC/jnJoZk+u
tCo4wqzEP0kV1wlKzqumfRX9r17k/jcZqidj9KjpMY0ToaAgKgBgNJ9CvKc+PkO8
ZP9IcGi9iTlWR9St0McoF4MQMRXN7kHay1PaDKXvl5qau6QkLKIghlbPDNJeaOZR
HMJvV2DqZQNv1qKy+9CwXa1MffpmkyWQsDNMO1QOLA3zhJz7Xb2CWSWR2fySVjYr
S1WVIpj0LBiQBYIwyKIuju90zoq+/WtT2IpjpMfAFYRHqg8b4/oPGONrenmq3sIl
Ba3OB+B/rMWZo7DOivD/JALd3QuH2gNTjGQ7+LBfg9NV+ZlKQTlpYKpz2jAGOVYK
umBlSfVvcVykKJj43zs7i2hivFyjfpZRKdGHNjLnQ1WoSFe4LhYNzdWN8m7AtRwv
Wj4JTSIwSfgBxAgz73OMknYDUpji480uh01AvbcESZrUPwyRkhSqIxMy1WSv3l97
buoNFvJznF3czKBi27utphVI1V+yYbEmoRxdVAi2qaiGJp7jePnx0LZasoijRVVM
AfwuQYiY2PbW5JcA2RJptpECPiOuUzc7ABZEL/CFybQCgwLuTzpl+ATgKNbHfIzx
7LN0GIgmRIO08M1C0qD4fho/B1+dc4uwWrlNI2Z8ay3p9NfzZ0lH98mg/tj3t7sB
77+cwJH6LeRX/pj2Kmg0Qht/zhcup1H1+7rqsg2wsJTHNqXwzZVy47XFHmiuSVjB
q/ZU9iJ1JdYUPFaNGdqcN8vebNRn4n6G5wMpjfHNA2IFKtBZeJZpchhjvXMgn2Q6
XR/JCGaL7cAJOyhJpjlPo81iLq+dHbNl+j5RGMailKO6dE5+cjjXqweCSBhwHXu5
rqV5vYpz5ZGQ9wuL76+bQpJovdY2ga9SyUG1N/YBvXOMuMaax/kuhcWdiKK2HOMW
8XutS9Q8c+VQh2a1ba/7eFLlYmTdNPUxa74WYoJcSdiP8+l8aRc5axhCh6yUqJLQ
63fGcsFSpEoihAHifyzBL3OvTZf8iqFOy4nTJcogzpIH3M9GA7++z8K3bk0KguO6
T5bPTjxhBzlWcW0VCnopzdRIwpajKqYctEZT8kZ/Z+MoQOYFydnlGCrJahdcrAmd
mpzBNwSEy4ImkbL4FOTK4FhnArPEzjuNmsOi21qi8opnuOo/VISv2rWS0TIKsn5e
G3yccmIrmUPpyjwvs9qYz+gd9u3FIKAxdWmUZx7ShkLPmCr5wzvx5zpvqQX/NEsK
fejsEsHIx/5rmNHpgveTjJyo8PaorvxvDup05DmZecKL1a0iHue3HWjOvl6wSnCK
yFAd36nkhTfnY9I/4tZyKg6sO79BRgXJjH4old61JsHzNJarpm+ce0RfndNPmnxj
t8Fb09ue7xaMmzgSsKWXbxLRutRRHxym9G6lhfIMVADE7sZoizX0lR2KJoRl26yE
TovgbK8sFUC3TuKVrNL5OOhXHXKSlXgqgcpIYKzqw6mKu9TWDa2k4f5xxKKZZWW+
THQaH6JBPqZvG/x1EPmJNNwLejoKsgvsJ62BuwuioyWwVEv/EUdWP4bWzmgllhDd
OOZbfmcaL3TKV+2LRvnrnJ/wRLG6ZEUggJkfU14b/lR48joWB7WzAlcEzMor/GKY
uWkZ90XXtMypnliSi62+W6K9CQq99w7GEsr76G/K8gxEG+kKvt81O2JMxNd0CrSm
Yhu8ntdDmoIER4oS4XgxfJifkQmPO3fDck0peyhzFzPNXVzbogocfFNhiZ3QZpZC
bOgFDkDhl/Cw8KIwBtdKEv8+ijBYPC4Y4rsi68YliVxROXC0h0pYWSZqVeCb/Qa8
DFIY/bTb46VwqrFHlfwVlMP2qT36gqeI2TXePNgnwNWnQkpreJiUJ9h4cUWhox/q
U7OxT3bU7J+DN0q4OwjprdvxFDtLDzEuKVT9TdSwuF6eF/wqFAB7Ay5/5XykRsxD
uQFKQaokz8LhMRTHhP//wjv6pZFUOcq1mL7ko8rxWBys9zjvSm1+OAlZEi/QGZFg
U0XrNxzp9dNWdW7MsyevA/kyUDK0F2y1ku6DAGJ2eA2niQpIfs6ZKNIkDb+GzFwp
InP+3jNlCXZNQ4hnG/hNFLWwrO6hXwreNLYcFzRrmSstTibH432OnwErEj0Ih/hc
yjLg+IaOJctS2PrE9gjHc0cyt9pRA+9Cga2lzrdiJ+ZgWtiptW0omGVMJcDOsGbH
SktZZ4InNnrdBIYV30XRQSAjZ0w0DgdVdMTdZEZkSEHjIhJajRnijjiM02dZmrVQ
j+BCl8y/RXoVvSmmKtExyy5OQWX0CKQX8db0NA7NWYt3/LT9ZQqY8nEjDGxCw4uj
dUhXMjkRqZBjUZLyguf3lSdIjxDNWSUtj5WL7tEGg6MMfCIYI+Gm/BpjRY1pbfjS
GmuXKDvJ8vxAoPFyDP5Zu1ehjAKEXp6cjdhOvhV0YSxkUv5lLiYdyuGLEne9c62V
uy6STFyY5HvkTJ0ISRzxucJHbv3/h1VfeltKLAZLfP/kYTtiK2cXmwgXlK1BL9/3
Fn3nUJ7vEg2pTyv2dTlh/6bcLRw6NDdFka5Rc6uHm0gt+tGWwVx5bOncRtltbU29
ijqxR5lwPe598CV23EH+He39v2McXVkEFsoMvPrCOMjYkfN3Ay07hO6neCVyH9iH
2x79UwomZdyxHg6teGUDi+izcJQfqdqRr9b6OxqO0hx1OTPmb6ABobqfGfiVjVVy
YPn5BxiwqF7kfZAk+HqnTdZpLXJT0/0cDl5JREW8mK76azM/H040/cknL7g2wxRN
rvQ+hFuD9ywG2bXjW/DvuhwnC2wMmUlOQYGBmRPozpGgfLtIlrremgbn0SdLIpD8
RO62qi2TTefgz98ZnCDVhU0K+9vAKbe81e5nyXQRtuqfoKbjxJ/bcZVioKDQMzJ2
susf+cqjj2e1BfRc9fhBlBIOvUE8nrm8X4ARvbleNskZQyeritR1a+VxlqaFOiLH
ns55WHd9KCJq/Eut71AAppqcljMltwL4CMI/iwU+NisbEAfda8j2oxK5esRwk/3q
bn6m2HWlO83chIRrTc6wRduil7wI4fY3Arb3/gZMPzJQVWwSgI/kg9HM86At/mCH
cm5sHf7w/tdCIW/hGOwBwbPgVUGuEb4JY9ZNGFkjzTwJ445+ln3Z+TEwhyx1WEpy
zSCP3mDB/FOCT+SeiHdBC9vpD+ZX29Dma2zpBHLawaTAzg1Z93Dtt+OXVcfhszwz
4SGExTOFTa0Vv4VKZgx8Go/U2hUj4XY/JTPkUAhT3tjHG2y6we6O9aiHpQ6JCu+f
b81gCYYJJVvyz7vCy1ahHORE8rvCKZf4NvQrzQDLeztpa6BgKlGHhcwr1Ib7E7Gl
PqBr9uOY1OPm5g3+Kv2StzFD6rWp6N8oOoY2gYYPcAxFAlVls934HFNONOGk6V1/
njb/sb2CVUw/MoSC9U1c0U+ycf4ixt729BRnOZCaxLNV6+1YsGequGhLJhCYoVmR
vnK1fi72cB4XYqsMJKXZB72HotCAb8oGd9woqNEJCSZt3Yyld3/oztjZR2kLsagY
u4Ym6kJCb2CONJzjO7WjwxLVXSC5O9NQhKu8iRLbj0z364IGTow7awf3Yy2adYdj
QP/Ef8ldKjB8bmfyElToNd0OGlgdpsrQptz96PTye5nCOAAsgslos9vdxwgbOWul
k26Hb0f3U3uN4uTrP009WpXEyxyVPf2/XORlsozrQRNM/WGYaqqrzjWOaX6o34lI
xY/sHdPdnGBtKT8rlKCuyqpvOV4v3K5yevxWpG/FGyo+SkIt8iuY5oagi83jPjXh
Ol3zB7PFoWv0UD5H9wOBa3BUW+M+x+0QYuvmq8dAGD7lAOZ/0jxvRT1UbNvk3Q9q
sZCIcX5ihJmMgkevy2XRro22+0MbDlgTc4W0jKl6yJNDoXnA2tzuYrikm9LTVy9X
TXNlfPYP7HaxbdoscxX7sWdd6s6fz/x1ntrPIQF222ZPYmcFUw5Zhq8aICuFq0Zy
9nrRmTGiCpIsBy4dCFZiu5LRSw+5iQkuXCeND3/kioIsRT4JxbUwr7Uft9RNkAzt
4DvNqN+vfLqYyJ7ORn1ZCpnh2qLn/HIHx6D91/SNI34LReb69D9b+JVXqOWMCDU3
y8HXDrn3f42BBZ7mi8rfIJ8YW3TuccdZwCqyDJenSN+azMOERt0z6Pc4saovYgTA
3TyAiJrfeF1sFG39sGuHJi+7ujxUAuNJq0WIaHwWmpoaXl09O/qgJ/lUw5L91Wjw
NGqiOkzXOBH4BLgTGSCDA2Q62Mj3LbBxPWTgmQcUvXDxvTmXkj08Cq0pS8F1A4Ya
D59YAquEMWA92UVSUEoreHcdqIBU5b4FJ68xVA80imcMb5dguaWpA4rA/xLXH0Jq
GXBx5r/Nv6DF9M5/fiVcKEKLsHpBdV5tBxAKZTlmClhZzMnCvz0/I8SUP4cNemdb
AuO/RmP94mpXgq6mIaRcF67l4p4IHSUab5jtdxcfTfnLg2N1/Np31D+oJsJficuB
6jL6L0FtCnMfYng8x03S6EElhjs/6OAxI9IuH5OpZNlGr8NuEkF+oK8OxuGoHqf2
2B1CJvJ+FW9BkFML9sBkg5docEXvK7lDQjQQ0PW6+GVYsErVQcsPxUI7/1WmZmaP
hf1hNxFLlef9108YHi2FZFmV1BwMxzxVYDwKevZ/AoDbv/Rd3herkFU9M+sAD0DV
VnrskJQP8SElzwxz5ipODcOp2p4tFkqtpHcU749Vh5M+1C8DIkM9MdiVwygciBsN
XZ6HRle26kXZFjfVeGuXTPm/Y2MsPN10xbxucsYBC7zXvrrEjtX/9n0mMv0rRTxD
LuLiUFG7F7BRtvPs3BQUBEg7VqmRq/NrPCcADz8Wo4gBchxJ4UECPC6va7t/i3ft
bQNjMuAhcDEql657c++NKexIhGTzU06sGBUQeKip14+BUu4p5NVtc//5N9spsSuT
K3rHzIra3JGHwFmxM+POQbf1V1/hOYPxfAZO6ACnSQN5e24Rf4rArsU5TyYX+tdW
K3zN6CnZeRzt/LxoG8OiUDuXwYsz/tD6lnS5aGiu9hn/8eiyHBNnVRiIDz2gSwLC
HV810JOEWezozOCRbuP3mbvVG8LakC1iBbO+ioP+bUl+LMZrxJUV9D+luq91hQv8
hdYQWZRmJK/ixTVHM1yKR/YOBtjFGXlYkWYCsybNsQ5YHBAj/b2lHK/TzPwvoIc4
Wx5nxszC1+bC/F+M7kTZcysb4bby2yV9I5jlGPRPfE7xkfI9sfYLejLANLoKx+Q7
v4AZOjjdQhlzrtzwIdjEpdYu6aYbQih6l6rS0PgkHg5GPWyHKaNlPyjH4yfSEIhx
C5pbnRDeYbcgd4DX5EnhKOEiLTJgiLW/0i8H57wnYysqk59JMKeIACykqytDMMnR
5hQfZT5ubf/j+4OPpurFOWLjyIs8EKITklDZvaqAQ+yaQKlwnb3BixPGEatqtiHg
vBI9KB9EaWDJCELdB8gOpKpvCxo/iw+TmPIfNICi2N3D4uxd+E9EADQpKx/K/jCS
l6cAbe6tD6D35G+PcHeHkwKA6Mtd7GOU3e4x+eOJ4wGqrAXJk0OIjR5RR1D3IyT1
SWRC/fL5a3aZmwHn7HDJglK6GFJwMT2EdEQ8TyNAvbmutoUIjEa1XqojESWBHskH
LTxCluxd7NSY+MvX+FJd13f9biAnOEP8VbzaTuudwWEvRIrP7Ktsx4BCNH1z/arl
yp8GPA68q3AienkhCQgi2V94GPL+G6liEOwmMcN4p/ZlRy+WV4CSpK9mZ+k+ubQX
wgjd5b8QrUKf1DtCZhS2xVCL8FMNbidTfUmYhGyVcuI91fk/kd9imS+QvtzvrkyI
YKj36Rbk+1MKXZkfSD6fle50xGp2y5WJYDD1S/boIJN4BR/4gKoVboSFORr99rFt
aGum9fGx48hByQKp+tx1uamgL6T5ju1maxdxH+DQ52eStB10t8mqTmL7ujDQAPTT
mp4qoWNagLVdunHe5dMqqKMgbEendbaGhQXeQWfSQUoI8WYoAaIYAQGGBYRyHB62
UEpCPkHntXqePGyyh2B2Bna0Q0odDfPiM3G4ZMiJ9dgCVKcU1V+BxRqxCqrtYkCp
qEmghoNU9NDbP0pUSc6mtpG6ArU6hy9QAYW0xsHDhukiWAROe6bQs2cUHdfQYOHi
wtuAxqdl5was6hEMlosKB6r89GQpNFuX+1vueFpey/Y2faJ37Mn/Mb6wuYzs/tnh
ciOuSYvqewewuZZwwykLiOojqoEyaRdoyfrcqvJKv2qNYG1QDWzVE6DmTveADrxO
Tb8dBxStC9FbL9mR1kJh7O0PfLZ47CbeSevX2dx4vsfcv+lSmwLlWeuLDiNiic3X
/tCExDonD15bQ1x3Mdy8U8MOdHEGpXcR67Bwd74HHArQDrOWT8udn7leu13vlVkC
TJg7JWeYkc4MsW50q94jV1fvlMKnvQRHazJgyzGT3CkaBfTI0VshNgEC/Z3yxw/Q
lGxSJ+tr/Rt4ZzXeWbZggX2vSg8/Wi1GFMTbQSMbE6JEmVyepSb0EV11YnER+XmS
qMNQS38hKZ7BNJlfiaqaNPClfjiekkmmTAznbgAmHPglfSHy3z/tzsQPDZXnPeD8
cDko1G9RDEaduZ/zoqXOQ0XkeR/i+rrbe+aJI51+XApeE6LCMB+33qn2VnOXdMVU
I6UxNbF6nqt7Zp3OGlMReLQhiXl3ruzBN+bamrahgBnIaIWIdXCpVGIbRvm87xsm
/W6OAcbgtKRUg+y8ai/dY0B9xVUFX+x4EqaNvGoEE5nwOVKpBYtiQ0bUbaJBNMVx
s05VAID76zUQQGxriiXbla84hp5MazV2g9PH8XUlVUCdork19/CNfvewrrBTIyrt
/eIpeaGz0VYueSc87ti/SwGWxEDkAJvejDGnkpjAmNInyzOTXElaFpTi8nz2tRN/
2+k3bQKSe+G1HRFlfvR2XA8LBTyG4IljaHR/1Pfbh270lc476bhxxDxPmlQsYK+U
McjK9rN+yAHEa3SgBQQvENU9ZiPV4/0B4lHG83CaeeVItX7cJ/5PF57s7I6UNlvY
bqnYNv87DSn6nYR8VTs00hV3WsjSKoF8FUt0ajTa9BhvAtnEXfs/f1MKOI0CQnE3
foNPXTfKBN6NyCD5u+hM7NNAbCIuqCNo5lK32t1HzGYitZfO9RsDVQTHKb07jGNv
PkQw6EXL341Cfb6egbqUqvyjSjdTlQQuFyxMeXi5Ynpe6pY+fX080zrjajNzPaKZ
GbosFMkNXXqygLOPfFdi5GtcsutJmArIG6/jgdHS1Ut9lzMdJiXXvyacvG6mwOlP
hRvwbPZ76Fm/WucvWawH8XskFLisyCAN3yIt0iQO3U0GkY+5Iaug6/CKCVnFF5nH
9+DHLy4TO88Je5zL1KPpf67/C5FGhVyyHBDNopltZJ0T7N29AKjaQvwdvCqQgYGY
xaPau72mCNrt+oMFNoLOCaWznkpTU2WyCK5nKOuIGcgnKqdtYs4jKKorwZs2ucZy
6iyNIC5x3psWUEFeBkDqDSfuDiCdRSXlKbGrA1PP5vPBTegnTZG5N2TGW90hEQCN
75g3NymiEhO4+P0pQ2qNj9lmeJI+K50ERUGM2qNq85h6C5ob9KMYVaQQt3xRm2V8
EVM5apBcIjp2zOl/1ErpVKMztx9s7XtjUoaF0e0C0Si0ac/j2S4PqWjs4WPuv/cS
SRxclAi7elKwYAa6v3qze4SKHuu1+F9//hNqu9+x7L9Q48JzhDWKDe19QpznAi4W
S77rWp3dON8Etx43cssS3DLq9GdGkX+v+2pBWcKQGaeLDTV4Bnbb1bPOI8a/ViLQ
v05ulYsX5PRsNy2KEGCkPf/X63Fg4KqHBGHImIMYZ4gCnNjsiNMuZmiMRH2wrKBm
qOwdxmvQZkAWr/ezZ+8BC34jJDyWkAfcdio4o6unYQRioZY9MGjJMl3iz6E1Onfa
Uzcqzw9L7EM3LFrVuBNWndHDYdhVW2RR4Qh+aDGzVoz3I49jnRUI98Y6fNYC57mA
1hrq0soo2nOEya+sV9TDEI7euuJGptCq+85Sz2NCG7lohDjJX7AxhjPM8nqmCPwO
Z2+P9/WqIuPHHlrouVZ9epsnUEs67C0QqiolxzSJFH6VCIW/3BboNlXHajoTOcNH
5JBnnYiqzRw+IkxV3gzziIPlQvguUy8TVgfYT/DM3xflELCw1GnTP7tYfTi69kyu
IkeAmtqOT91Wp859lds7wWSVt6bStmkVsHdpTBw/pU4Q7FepWfYcks8TQRtaZvjC
Kqto4C67Vf6PzPDokpPqFmj2rfUbUh/ecXhuQNeMs5V6wOMhffpMuS1h8db3Tazn
A1cMqjEYG7SRDeNkCWGaEiJVftrC9cq2ISgDpd7DBk11GZx3WFYQAAJPuamf2RmD
JwQhfyBoCTLOPwIQPrzN/uoQ7koM/XLZhIoNXjR2l76M07f8pb6Hzi9OETqXO+ae
n5i/iQNHF/LDTmGSVD/0RV0yALewKx3HOBuW2NYLVfJnY7Nu8Ng24yi5Cxp/bpRO
Z5E2pBcDb7cTSyOHPvsbXGES5kCTO5pFz4TU5ioUIyCSZfegaxmmu3ceegSwyz3v
zh43FnwZse9jo806w5nKIV24DOoIOfvTmVsDREz4V0WK2LOGPgYlYu3ePgVaf8Fr
GbxcV+MFDanXsH7hIH6CCHBwVdih7qtMtMoAfOIW0kffq1dh3biCP7gA9CPrco0P
7ixGIhNgNgJv49uKhIaXzl4Tki7z8T0d/J75X+02LQG9ZcdDH/bz5VYcsomV6/xK
YeZpVFGenphHTaodAztXqe8SKLGyfukUNuBrMynegawSrRPoDerfa8GO9oBfq5g5
6PaQs7I/2lGYTewBCagk6cNH9NveOSiUjr7a7m0ekAqRwf5tq8jlTIjuzx0yWW7L
sxpbLT7ODWWOv2zkwetCnR67OEgwX1LkIdoo8gUQFQNY8ZN47yiN3gZOc5xOkUJR
2JJQjUtrIQP4nQ+imEudfVNB1OomkuoroDu9V3BhggWOQv6q8ScFkgCqe+dPoMIG
1bhzHblWdaxxTvQErWjVh/yqhQIpkBHgDkQYBT8frVmi6FFv05ELrmiTwHrhfNpF
8BzM2PPqr/eyTFjv5qG3+nFr5jFX54j2tOqpL3FWB5yXNNLqfSLpob3Nd2SZADUw
8nxd1dfJJqli7pI419dLtHGhSjSy/FhWGZi/jgRhHB4K5pdYGq5wYDEADA/Uj8W1
g82w6FA6fOZPm1jY8pzdcf0Z59CbFREJmqVv8Xj7ybM5OVAn9yAqeuY+S1822EIe
JvOu2A9zRdbr+PM3a1Xh3n72hLpzgiNOJkT+OMo0iy7z/qOS2Wh4ANPODe7BBkEB
3nQmycJa935hHATpH788mPPyzcTPg0drl7/4i0/eaXs8bmHit42YgsJ7qRPrlxhu
eajbk7DltsW2e+c5rEae5FdQ2I0LqrkVOwUNTFweJxmVhLWVJzxgpnL9dOHHiWxE
X9N281s4igkEuvwJ1p1jQf+TCPT56mV1GSQ/tUnhYzZx0Em17GMrRgTeh1zteV81
SURc9zImAMEfkSI42WTCeggIfnjG7UwL+2tlHzMJLpVEjHKCDO4IN3U88Q/rKsU7
W1EoYHoiwHDgUh5q8bBp0sbPpD57AzxRFh+Ascef9PSmGjhitIzF+V1NqnW84ov6
beYnE+hk2KJqkKK2PapokNqIfAadmjQ2tc6+PqtYhPKr107VQ9bTLSbXUtPQVVhJ
gNpP4MoGDxVJ05VyYRFaKLfq97zO4Hrx+y6XHA0T5NgXi4IQjYpFuROWGJtpq3pk
DXjHDo3sLzU1I9oIsPefBKMx9eMsneOhm1nHudvmNOv4XDkXkTlNFZFDoBrIG0pw
RDKdWtrsx5HQFq4P1eyu1bhMkwh1vevtTrWf1/GalMwvvu0nIHjhP2zgcKpnABZ4
VmgSs2zwAC/QAMqcz1h1EG7jkq4dTTYQrTSRHWr5Z7dhD/xtnCAg8CKEY+CtnMwr
nwDrXqDGuk+CtT4frPjyjAuZ+GKue+uQoc9oy9fU0MBbY0aN+s6xtvw7ApzsHKdX
3E4M9nZs4yh65hCG7RH3Me/+21QqWOrw22SeqYXhWMS6hwVLZ/xw67IMkvFBI/TL
YYt8nqTeNIk4MjbAgUES22k4he3EjQTw9EwJurzMPGa7/gll86olswLkESZc5tmr
k3j3Fqbpq2aVRPLw72yjoPDqMxRZQEEa4NXAAKZlG/aWvuuRMwcnsPN5/KN7CvUK
hy4zxWm4GDm2TuwfDG85aoHj5SR87B1Pub8tEX5gI2DNpqFUbn3fh8sSRkco996+
4XEzSleWFLwK4Xd8a2AEihNVF3AkZwnzEcsyNS/c7C+mPCIID7Df4z2T74928a3y
jJoAXB9RBiwWK+vOl19WPRaoIPVniCEngBLBsCfRQ4s0NUCISnX0d4LYTD+4IxKx
HXmCl5kKkc7/nhd0EZiKRmrATKQEd0gBlbvIepxDfC0KoTftIOAymK2nlX2J9wIf
JqpfSrCt0YrFPozU086lK0yV4PfEkircGpxCYYbGFbjgY609whtIUcRBvg0iCxUU
QLOLghQ+C+xP7zZNXgyRhaV4rx8OqA2CSyahqZGcJv6SI+FqvYJYec7xxFI4octK
881D7bPuBe0aJKtHKk4OX7DLzPoAd2cVdIDeunwX7lrUTZ6kcYwlITehz/ILOX6S
+UQYmbv8mteZxPSafivD08/ioQ77k5y800y9ZnF6JvdTk7VyaT3n2I2wxiQRC86S
OhjBh+J0F7k3/9Q0WQzg1v2APPCV49wguq6Om0V9Qj+h+6ftI3+130Vk2w9g1dqC
2YLNnsOvHI1N73f/biYwgR3i437uAYOEcGNFgyc3XRKO/MQe8dC2luVSwwmlc3ZJ
S1xntqz1GQdt1Z0gFqgV4ubjiKY7cquyZv3+JuFcM/nHQRKdrpZdF2feI9Th0IoE
LEoqVA/bToXqC04ahVj0j/Qko1vr7AMKpc+muDcZRk2v9AAhe8GsbL6CrtBo088M
lEfx90z/yZUkelklcqIXLYb7AWFmVYHEaZbLQqvWSpgfI7u6ifGCxbaVtvCamW3Q
7o540eqggdMirTna7bqizecNmE77XZWa3F1Jz7zYj1TtmZIn31nk4xObsILQM6K3
7wnSXHLNsMERpd7uOgR1eycTvm97VI5vj4cET9yhZY8ViB2yLoJrnqzsjG3QV1NS
3TKQsEzGVx1GryC/IZKLi9UJvfUwid8LImIcVkkYhSL86n8WsCTuGeH5/64CZufv
MQWY0j2oQ+5LJ2tlRRhblxZAPPrFqiDfGuLsnj+bQUyhGSGrjH9aUS84c+4S/8qf
8oFsPtVL+QdK8axPxhtlTKaq1Q1hE8VBHcHaY4LI3EKgzpey881EeqZEt8fxN+aw
NFGrLa6rfK90ctgxjIqJfqI0cP+iP3LZ0xJ0BkDKHyQmxqNOfrkCbIHK9BqqXPqx
e13BVMYB2LrD0GZqt9+n4aXN4O7aCjnKehxgunNKVnBWB4OP8PVxlJwnGKYcenrE
mL2mtANrAaIgGnmwWurHfmXZMs+skthp+XzeDHNRWYkd/3tuZvWvFe6IKNu/+aAa
zmBA7ne3nzBaJEc1qGEYh00GCTj0wXSJBQ2ByHc29i5/ALu12iVfbYCjFyAU8d/x
zw8du+AjN9efZ9lOPJ9rDzt0iRHovKeV5Mnv7EidzPkGmgbob6/lI1B2VG1TYpxZ
EKixZj7TeK7qJ/vsj7FbOidiC1GxX5YUMocWZu4sU3PtQCISGhBUFkgku7HpiOFT
b5TEBgHgKhGjIok18KFQ6uEvB72zP5EtTbUEjfJvU3XwjXXVaeu8HA0iYylb8ysm
km7HOi55FahPeXb9miGGqnvkj9cTeU5/gcN3d2/HN4KyBHS4rdv6wJYRCdiS8kc9
lWRxxucY6oSsZUu9wdgAa0t5KRr9tTHVbTj5QoOc7oqgxvf0/ANo77NVqkwcKBVb
fVv3JHnC593ikZzGC3p/PveJre7GB+Voxjm4Z8RhOQR27spPxogtfSfkJfbz9ySZ
Lz9s4HJRI4lhMcHRL/cwvVfJcDxE5PhdDRD8sqS4gRzQJ9O3DjBzkrOClPbio8jy
4T1vwv/x7JbXoSfblEKFDaVg5Utnhc3ZzNuHL7eG7lFLkMUqjucGU9eyoJIM6Xwh
aCZbv0vZfFBziuXUNfXZkGeY1GiVEOxmyLy6B16RuPwQ38RTXRs13H2/zk3gPP2r
sU76DA55zaF1ku0EM2fW0c0KRKCME1FfPmwFP3Sf37Vx1/fRX2Ie3aIoygGdKHCu
2qkeMm2xPjZbu3r/1KxX1z8Y0fn9zyD6eJuZgOxMFthlogr8JZsQxhHmJyJqNaV8
q6Iz1UN0NhWKv3fu/sbkY7PPKsHqryETc4LzrKzX0NJh/p4rXARrsb4bPynpIsuK
QGgq/soeNkfeOzwn04y91trjxHSAF//7I4tM2HsFFRktkMToJsjBwjjtvt5+nYGn
QjDpXhgLiawSlw1fzvnDziQ8RLFFFYiX/TM3FcXQRMlJpqESJcI9sVIVXuE18tmQ
lPK1s3C17iBas3MGwz9Ubr/I/ypBr8QGuFYmpOY5IY0ZTgGQDqtAevXQvM32JFWh
nUsqozZnOfcKoB9UIw843f+0Lo1GpcEfI37CErWM9OFzPtQDdY0c/GY9daABmxC1
6rwr/TrxaZk8Uyww9rUBThf4kcQCNRm3tV7vMKE+RBM0Pxyu7k3kxMQQO0uM+aL2
xSzwbfvRXWtqixFysjtiI2DWdnxlRRIqHx2jNd9zTPcurwOA7SyALm3oj1wghHmY
2gJPzEB/qOQs2fF1rIWWYP7jCUuCodFufRqqoo9wTyucV67/0U4EXSGrBCi779nl
iNRn34EmfwfW/HZvs/ayOcwnd1sAS2rp8kmCobQ2ZUPJSC0ckaj9QgKLbsOHhkei
HgPkKONfi744Cp/ifFOwOb5oioo2Ay9zyFkkO+9BnRpwJkEFjuwjEkTqzFgZpOK1
j6Q1gdwCPZvs4x4FjUoIXZULot3Wn0ng/MbkF9wvx6KqwSgyVoyzgv4hVXP8eYpJ
wTOQaKokW6dfV975i3c4tQ5aiMFTLIeuRH4818VQLcxNMERDwJH6EkMbZxmCu+Hs
XeKggX1go2DYW4U25pS3Tvs3rGBuhzHSAr48cqCxaGiTCOBpcpcEs6FVSS80gGM2
hKUszMBjOIovjCT7R2SaznYkExh9Buvw3ZTvtb9Cf6dr6Cwp03dvRFxmy0e4sgnz
wdwUGEiehMmlnLYaxkA/2RixOP05YbpDz6SJP6g1uP3LqzIXrlnro5jL/DuVezKI
Kwm4RPj+5s44cgfBhNXOK3PRs/ow52lOPvSWSj4OaYBRXTFQzyY0hnW+SuczoIzV
t9SRlcIw4YvqXMP3nHq4tx3WVMVlVl0w10TuFt+D9KSiXvwgXzsXswYJJK1caW9r
/1ticzkHSBTFxSOLbw6FMTnbGRncF7oaAAa8rWxDFaQNiMOVs4qmm00meDZqWauL
Y+rVU257pYsoNNFHuj4rhXY0tN2SfbJOZjWexNavtb3uzUoVizLvzcT97uJUlQ8u
jU4PJg17/AXzAgHd1ImQQ2Lp/vmQHQsPoEnamMUyfiqtAejykjxZzVmIM3JYKj+/
M7UCTnqeyDiVnvrewqVFOxgOO9KdSfkUgYRvx70tMt/etsL2IWiC5vBKpAOhL5Ai
ULbRZputiVXsIwfJdxQB3Ti96/GPTduj1AAOoK2wrCdW47M2oPXWGkAkJcQ+bZp2
EiXD7OA8ypw2rb4MzMxAtaZwJ0zUOpb5OHtO0TNv+hJr/Jh9U4TS7i6Y8R0iPvpW
RYg0BjxriZOKGugjZAOss8ZhOwqAdK3P1qopEpnqGTD+dFmm20XyB2zT5ojZx3nG
V4lkLO3+GHfGGYIjd9DC79zx14EgrqPcc6pBcHp7ZcasOeqNS7Os+R0uGt276Uf9
31+E8YgsuEzQMrkPH+3UDJbyMNMy4jb3SXkVjwwRkRGAAreqx9md4BfqP/GM5Bpj
nN7t4W5zHdj8K7Cfoiodaje9YAN5hFGwOu0aZ4BtPtHW4o+BNsId9pm23oye8S1j
s9l1Ma8Nkyf4XWRcs0leXjjGMg/OL7LWduV/oQ+nOCR7wue08FDxkatiVirA/2yv
IZMrwXCagsL7v/vkYo9c5nwNBiNxT/DQJx0FgRgBieD71omnFH6kFOk3ocL5jMCI
6yMDr8iJVcqqJ+Bq+HfA1SzLsudwjrQvZSeVSH33jGDKU3hhT71uJiP0H4eNyjmO
SvM/lrcfXGSil/2rQEdWSm9OwC3t2+tdQWdW4VxoxuZQa1fK6+5S6FPfotrq9bwN
Lbo3q4GnwksbjtR1hr89g2mT48UW3MoDOROsMyYXagPWVfMHVFVLk15JS0pRGPXF
O37oygyaORgXQ9qMrQnTeQ7uDvCnoQMbSGdW5oNuKzOj2CNrYO3FjQQ2HIwOIErn
eKKlbpbF1ANnJ5r1MKk2kGmvXRKSUUCrKIqQ8m2Hdi6wRyIcw7ADTpqmADZpHXnB
sowJG6YR7gNo0bsAGg/lVfXy7q8wbQ6s/iiZGmsdc0vJ2FtCHCVmIIKc1pY5F+zU
Q7wcv6jAvGGkHznZ9NPl1+DED4mz82R0bzh9tG0q3sTruQpwWW4ffXpJsBgGHU7K
AWzOJjPVzjkjNmSKKO6I41sFNLmX0Kizxw2Y9oJS/1ce/ht7YdYwrkojlNcVL3C1
rOlzQa6JMEpIHtYs1JaiNlXLgokM82wie+o4xjlwlGs8lPvyYbb1PaSu08yADcWY
pWLj3Lz5dbjXF1TNIqXhi9bopH99uYYh7mrK+9hgNQ4Pd5rSMx/RVtSaPt0nv4Yt
I2aHswmDlMExb4Dc6Iq7fCHEsOdUk4kJzbUaoSKamL6pvuOaiWB8JoK06Lef9d4b
cz5oSJ1gquEtIzZ3i/FDyf5lcMaT1LpGdS8Eg6OnFTcwSuDM2bCHuE1LQbtOL8vQ
WGEGjRAC1b5HHGJLMe8ru6mkMsSEHd80/nooiESMBDHGxdKL8e+Wa9vyfFKReQFS
2kR5Mh8QBuBgB+cIuce8EOMKWFbUh7VAGqpx6d7CL6O5MKkaBScq6kNdX+2+ZCph
AFBTSmr7iIrzR+ga/krC3BFZR/SaffBtXUzOh0MFrayQ+4dBYLpV5RB6axZ2x2Mu
aoDcyjRBxcOyLG7wd1fwOiL1wS4rPE3KzkckJIdgHJ1u/MyqvCWKZMBAYyZyl6sj
Z4S035URZDjcGq7WRKr79yIq23DTZnnaXvrRIL9k1c0RVdZ/iF/DYTJ/zIXkPE8K
PCPJCKUW/vx+qkG2UEkbiAiHpDIM96IiGm19ostS+gqyXuRVgJNvSN27pSenGUxt
t1Nx41dEkXzvnQqO96ZRfDriXY/dY/l0TIVmWTj/NgAoE3tdcX3VdQGuNjR2JK78
g66SaoSjelwiwJBOz2XEZarPrQcUZGO9eTM32uQWKV45IfpFJeoxQ05jfjbgutiM
8JQF7Rf3aJU1991Cxv7CilAB5RomWLc59SIWQsxGofY092G04P7oqFm8WXQbRcXA
GNt7osXKhFCGR8javAWh3UDHToAni8b3Wi6pit26qasC4Ak9RJKh1VZ2X5xroJhK
wHkRlj8zirMqyvYjP8zlf9EJQ9vu7PEkihfKDCIm6U0qyRgBpcEoOcLsrtCs1JEh
3aiTTSi9fAJWNDjZ4h99DQTvBC9c4BJ2P3gF05Y++MqwQ8+EGmxqv+61wGrNN06C
r9082IKf5CipGK9eybAmaODXBipQb5XqMYnFhIa9klUPG3ndT27iI+OgraH4YO1Y
6uHTu5xdQl6Cnb0Snwk4WVt4eH1EPh3KP2fgj4vcgIIF115HoVPc0ODJkpiA5wnK
O0FikElMxmpZVSBb3wvowt1xtgMg1q+0cfs0+SRmDyzChEVMwNIY7bK3pQzVAVBo
RTV3PGgMABXmjtw2jGcqp/CCmnd7eCra24u9U8RYletr5Ku6n9O/na+F2B3F+Dv1
sZd5vgAjJbP/YXEE/fOgkwvauKIJieP7Y9XYBNlaYy7j12pxL03Y0r5GQPzSVPOF
2Re3wBBvsz5ZNvrmWMeqI604m4LsimPCKxLRe1AVHgUrltVJV94B6tILIi1FJ6OQ
s4m6EPhfasqAry42qufFk3uA2di8bYid4PHfQJgvhxAFtTtoQC3vjzu9Zjxy0+JG
WyjPXLh1/xC8pcAWyfOg+1XgajezBm/PvpK/1pv0PYRvA7ZB5MNTlBUQvoHC8XKc
9qpjQ0uuodpF6WTjYUIFc/j8zngPVTXYB82dpJ0fDHSy1x70XFeSRKlZGiP7jQQL
gaw7eNTNr5JGPkMOeRxqNhQDITATwwglzyjcShStiD7mXG8laVixc8cBS/VpMzUT
hjz6ZXK3qgK+bWskzyDr+3/6ugpOI3VL6n1sdrjfSnCHNcOIXvdne8naPMO26RcR
kYg/VirFYdYvFeqMHf6KnKAjIxA+Z3gZGNfnf86EKe1wOEM7n6rnHtk/z5IMVvfD
BjTY40D1MdbYvXyqfQRuwlHML1124g6x+latCsQcNBF41zIcL9Jq8KBTCbJWtxSY
Y6hINeTs/b+seJKMsjmWF1isAAc+ixmmxVJDQr7BXF8WrXfnkEWC3+ybEzMw6lnF
Ep7n+EQxt8r6Fnft6vIXZZHdhIK/yrx8Ox3SNJ+OSxx1SmJXbHh/NDQYuqR++hpl
H8E9gGSO3z7l1/9uisDE3AQ0PmgghNk7+0hThNCNNxVKsH5F1zDCF5XHPMmoTmaT
TK7hNYoLCdTpyKJncezoRAZWNPoAgNJ71JLt311TolYR1akIbasquDrOK1ktMipG
TjiuZv7SNYskPufRat/kX4FJIsikCvjkgHGaQ0gdRC6PaZj+rjJ6mrj9sXFAIfWj
bbWXevuv1plE8QqG8mYyPZWIqOgl0LCiFmJ2HzmJXloig/WaGGvkKx8/6NK5K5FJ
co//ep0wo9FSZfAuvFakBxY0+gTv7QkO9W3okGpqBvlAvxuKPCwNbx/o0nMOGHWU
ObLkwdVDcwk4xRU5KY40mJmYkMrQfpg/sXlBi//WLwYHdMWMQaTi+vFlZr439bs+
6cjCD7K0hCmseqiGr3AIYlIym/YelBYLce4FGniOR7xnMoXRhvMl9vU35gOHyGBj
IegEsGDdePO6pQI9ne/lLGk6u4zdPf4C8N9g0WTI2F6LxuSi+IxPYwwWdXayUm6d
1oOy1UowS39naTlPNOPnx2sfb4lD9uv7L7xHAWRW40yu40ThfsYkIpWhhVbx/mk7
kaCCWiAYBw3UPaiWOE2N52EHZHbPCMi4mIDs3/CDu1QnjDhUnpFeYTrsEgwLYXEi
N57OjZ53+xuCQ7OqV4HqNQoqj6al2QNI4tCBB/rZu8Qzvv2JSQdZSdNClJb02pDD
e/euHSU6G3UTO/pjSRbl3CEp55Ow7mDNw06b8krsyQXCXjVqUncFTf3OU3OWajRP
dgjAsXtB6n8YEcyqB8J3T+iE6LqZ7FQ91sHTzFPMZRMBElNZfHS6kxiVYCu3rHhs
6XBAtDG2UPuiFb/z0i4W1dHUXNGuxMxPG/ZZF8o+d0pwmPFz+QSI+yZkGU6rIIJg
lEK7+X7wd2rqILkdcmqNoiYy57v15l20MlV9WfoDP1fVxstd7TQZK8++b/8qXDGb
12vLavgyRYS2Y6qxHIjwra2AITA5awYyadkhzoovkcohvxH3oiffV4HJECgKkFdl
UeT9175iMNMBFYzCJ8IldXwUdw+VDHiu/fXlbrfsu/Q9wAxkN5bf9TYWsgPLY2Tn
R4R8TDzI4AND2KblVCgGL872xnP1oofCcd0g30BCfR80AnnurnaOMXEIN11gGqdh
2uV6OdlRsopDlrrjoO+7BOspy4AchQEaAZqi2+Apq5fC4yFCQdSpKwmMW5eRaTO5
Wb0w4yeiJBpBQkl7/436GIiVBpQ/gBGI+U3V1bQTTGgmEigynHRK62SuAsGsjWZh
y8x8i64Qwh5ap6RcXYFqIlkPO2D2GlDZPc7Sir1RaBq9UzQTLGlrSmRgyoSwRBG5
Oj4ymWqB7XJ3HQ+i6UfNwmhbw/yTFMkKa7cg3WJH95di5lhcro7ZGJRhkFzMRH/j
I8Psp0/kMDl35PMMI0wHzCM0osSDkqO/SvybID0MM9V99brSKhjgJuLbIjtKzRDV
kK+cfT3oZI9VObIEUolazPJJxqB9n5WhI8VwEC7rt3E/SYrC8V0pMThUOhfWQk+6
0IbdbMxZPJhUiDqn6z059xnt5Q2aTNMOoY3Rp1de4rzKElJTBXYmLpDxWzQ6/Qnh
/LneZ0fshPnSgvG+pPpC/hV9ydUemQsfYRuRm0kAwtDIswOIa12up9YZTkj5e73z
uMDw8yna5AVb8CfozVRYvHh0ECTniz42p385lg8CjWelukCmv29VL73/Giex49Ne
PR87DJ/CKuq50pqf/viF1P4twYkLcsxtbnTGEfjR5LFbKtXmn8kkR4volDTtRqRn
p5ZIE7lmH2GcjlKeiQgflCbSyW6+DhQNTle3G/S5R7ODiVeeKyl7O34oHTt28nJN
N8y9pp9O6fOlYOWH6SgRMEEiIr6z3hi1ku0I4wcWv8jvH6F/c46lwekR4NP+WaJL
+eGUU0nPuNEVAFzH287+8pM+HN3WD4XcId3oQR056Z7VWchjgfWJlLWL+6y+Uz1O
/UnirCloI+oHzhge+/tjlazaAeUBSl9K5b3EFPtRwvxCLOH04bXzIUEvKfvLUh9v
ji+k8Twtqvq9WCU3dULAKPbuP/oSfBgPccTZF4OT30qG2RY1lprSrFCX+KEhCWzI
LZDrf0LQ47OHvH31DDTZPkWVD0U8qKai1aUtMfOKGP7spgPMyr7FB9/ZlEOxJyNy
rd6DY7Co9rr6mK5gB6OGMEVr18b/xYfRp3RT5o8NfHCpQOcH6C7wT+wg9/EaT0zq
RLQrZZdK1y4XDac7e8VSyV7GMdhehe+9BUwwYcozXHu261IEOGieMGR1608GC+Pa
lJ2XDLI9wTo3QsoocZejdOArfOFLOuZVZHpiv/KCDiTZkNxDnkxnH5cs08edZCRJ
1SuXlLPlK5S4+amJ0jORzzqwqfAD+7Ewh3Qo+3+IUsd/cTVmtclHJzvDvWfsNnWE
NArBZrP1qqiCC2XSjmx89qHFMZQ8JpfScqQk0R2DG+3zY+f9i+Gohs5yQGFfW3m6
71SolzHJNEs0QyhxtIuh06NHB6ARKsEt2/DHoLXypd/0WETJt3co8Y+q7V2TjKVt
adzRt7eXPtZbU30r3f65aAcjFuNzrP9JI2xtqIZ/K/242ydPLEv60QSPgDsXzEZ1
zhmeD+zm7Xe5u11z01GmunYOcqOWC2zxgqfHeVxw/dMKlDyHAX0wXflObhnmRMmB
zvuCoVGtOv8BggqNIBwty+wGVTcwDNUKVLGmqoIsR2pYb8piBsrcsWpFokn8n94z
l6iB0SmVpNx0NXir/ZgkCzvsXQApvD0haXB3XfcBCnriEDJzrFnx/XXMPOA6rMNj
coW77i6GittSMnUwmPuO42FCQAXwoqf5E4knKGQ86/UO+3TZWSzuCtUnRoi1hyPP
AkX2rTDQ7r1Y5SLwmsZWnLayZ4MhwMNWPq+lssAU+U1ZK+Smwy2Lfy+kZ7Mprwgt
VLCNBzYr5BZtbLlUoqDBFIvLxILDhGBIxc1o7OnDXrargJeFWQJng84CRNhPJRfH
WfjDypMKfpm7s/j0CUrsBONmQac5f5xMYvgnBlSWEkUzeNokVbNK98laSsK1a1sP
hifUqc4QKNjAXQg1yAmYtcYydcwZPc2Y3j2ubdVjO3dvDKKlhHTC//kCK9D+8x9B
U4lCNmXapRHNQthNMd+ZniqxZ/NYtAZl9dLzsv9Tes3PjXT0r7LR+TY/Oqic0U6u
dkO46AB795wlfCXKoLPj1aOOu2FSH35VWGs7Ho/KwG/7D3yKqgAo0o0htJSivjRK
hs+7SUxZJZGnPLf3qfyih/QzfUio9CE2+RU2TP6p2ZI54WfxRrzc6ztyczVlHVFm
vIiEmNhfe66PeNTSjD/f6m3+7zGxG9I2/uloRHYlwoWuQ9ulUf60G634j7y3YLP/
YMuss1FUyCOx872KeWdXM7m/mQBsHbVRoZqffhQTdp7XuHPkuzSj/PijUXl6m3hv
7OmFsA7mICqiuFl843/HHDbojoaDrHZThEb17kmrsXY6pnuhY0t0zk5z331xTLBw
UVqhs6BC+5WcCpKsOlwTpEgTIMPoizLzriAX0VkGcNoKM8RrkGuKfHF+OykhM3Lp
TELRG+xQcouun8FlOTVaUKvldBjd4rs6/drBDMC6HKFQaWUKZjyXP3aUzzterTZr
mKqRTnRIVyDR6ogdNu4hMSbCtUQ3hTnNm9AyjLLaiJTywSxtYQFzTkBetWoptEso
n2DYcKULEhRCjn7Oyl6l98+drTRRGeeZbHNhD7HVgNAL2vmMZllPm7aISSVZ5Liy
yqv+hPwxQkv8v35hK9cBE8TtdIJjUrSkePmeZsDKrneX3eyu3GbQ/1JoD4cn2WDt
eH+LFOyEBaV4gnNZcX/cqxpcFCB2zsO2bzJ2R9QPueNSAMlRu99pGLP1wijMTwqW
kN/z0noZ8KvZJbwtuq/uzI5tM8sopuf99Gy12Wo6NWMnNGt2TbmXKp3t1squlnNT
9Fs0mPXpBuf0pJYaYol2XHxRVepHHqal8N6pzTLmm6y6fwCBU5DLaOOjEECAWkzt
pV3S7lPDq+fkWlBztKY+lXKtJu2x1NA7hTPK7ok6+6BHb3o9AloT83sBuc7YNJpX
KT6aD2ZE3OaD5gQqEhys9sNFoS2oHjCMIhDU44JyCYqShmPuviVKCVlEoDvZBGlh
pqibDEIpvtQZW+zHDmZsUY7NRp50ItWHRAcYG8u/9IwgCVcKdz0WpZ2aSX35Ghy+
SJ3BmWxpBwbz4HlrTn9y7/h8/gN8DGAPzouDPQ0A0jZrdn5Qmxr1gg0ugGb27zQ1
IzHWDS2kPb6Zc6rlkPjDncsW+DHMznsIj7+a1R6FPw3QToW+0shrmBkMuKDh7rm0
egROLfK7J7KuFeCzyUI3dQbRXmXzQdM6LtHAOcbtqD5xu2O+XonGj6QARIbYCTFC
s1PgZooiFeB4Zl8A+QShdiFIqgDuRpi9VBTueYeEU/a40QmT4yeQY7QRiNVA+wSX
YLQialzuIvdCrsSAc4hZlWEpytJTHFq8Svu+S8O3Jm10tY2MCA/xrF0YZUC+vvWA
AQUpa++IhS4A366At8BZVynomN3YL3cveJQiutQroxSsYukCjVXkEqZ5UV3Hw53r
HRzvvpaDowKm3Rx/V+5/1Gvo792tiahPikE+QV43s8AaPiP+jUj6FH6sXaZnzZLd
w+0Wet4QimFgYCsuOcSvXMi4ErILdq6C2kbxOQOLsK0Pjq8h8jce1clcQodpE/0S
yikGSYnuBRH1GD49K7PvH24cvOERbkWp517PSro45jDGchkPtpcpx0Bqo5QVE6iO
5esmQAD3hWoweuZi7Nz3ujJPFel797uKJUbXJgZ+uWP7enSQJCcwu0JaB/No8q4L
euzIwo452XogIKY4c9Tpoj6Oua92Q3sgQPtuNZhc8pmbEItNsjjH6+4m7PYF2JlG
QSkrcgUIuzpupwpRQcmbHTJOqclIyrzIA8fFvG0B7xlOfgYpldkCJOmXm4zqp9FG
ntxv7CSJC45xmiSNIBS2E4155zDsbc5fY7w2qKbog1pfQpSZCbHZ0GB4DJRXQcsd
vtJ2/7SiTLNeBKvplt87kquUzFivxAhKFELa4yB4zEvOlyWUK6g80ivHIBq+VGtK
+RG1HPdM/ZctHvKp5K8IZdBNyEJSkht77uTJyLjr2TuGzIodg/Iam5HT28jYYSma
xQtK/eqhrOUkVa00JjV0cMHswD+ws7Omu7lQZEFAV2KfNshfNj+S07y8IEgehQWZ
iTQA85jlm8L5ZRxZZY2kEYJmlAzCdPzFJ6hWNtYBM9Etc52yf8ln1BRqa9IDLVJU
0U5p5YgoO6kvlinLDbC+BhwhjKeW7nNDcntv+sx/pFYKMK9IcWG5gHY5rQj+R4ww
GfpWZFwE42N5jqKyu6akuQbRo7xphMmoTc5rQV8+oSLP6+MYaHFdDBEeWq2USrP4
YVriCbNTHm6Rv2KG41AhSxQMWNDf150UpIJTnkiyQ4KkqUxBbKYzMmG4VZ0VhuIq
Zzqx18RL5hXaVoXrORx78FrVnAsNKWO8tU9WlqEdt5k9PVXah8RGHBv/cZAZci+B
YguYZSJqkuhqJT3TEteMyUbo/VBpXnR0lSLNb7dsDd+rTxUEcZ55WoaaDmZbo3bG
EigyoPkLz7dQ7sAtUxcB+SOa6n5rk0UHi/zyMDUOXSTTIhxEjorXViZJSendPFwq
3grXih3GOrk/VjMt5wm+77+TbZCby9Mfx5INILIfryUrw9y2b0F1twIJNPs6f6sG
rtWNEVEiTwvjZOYSQwEbX9rFrNVTCE45PcJGIdYaJrLxj2jretHPadgB6wsb7uo6
qtNqtI5OABAhUiL6dyzoxtqOE//MIOUA8b1bSx77tAmCjKxaUiHexJlOyJzYhCz1
9GI41pWUsOoHo0r+gHoUzcEbZW6D+721cmNBkxLAUXCeT8KOFpuZs+M3zPJ3kyVq
A9ggm4/ka5auKRzmU/xqJBxqxy+yoUe8Iu2nXiw7FpI8OdUCH2y38fVjsl2MLYA9
DVsxbToWXp1Sn6UQppe8lqHpkNyiSUusXXW1srM7uvBMUPlsoTCh7oDt+nfGjJay
T4MOTL9Taop/UIzHW5Q4zsmDKkXFDoHyD7mKUyzotmDNrtFygLZmzMtub168aiTu
VdHQ5GVrL7XZRl4QqAxB4WPMSQZvyBsjCMuTQfY/6405dGW5ab0O5o/ovZ4Ni0qD
XwGIte8Cd3Ixz4rABVsD2SYUh5Og18ASFRqhTjpKxZxTHkYXoRFWWsDwEVUGb+3T
H4gFl6GVmMOHCfCfc+Dy0+Xke5jXV3GOqF/k5Z/8ql6usz2GJqfDNzDKa/dPfWts
bAjGoa504QBsm/6OFoyTEBdbYHwRL/5mvjmNcpeVvxFaNCHTq++lXmr4wSDzPowa
Oczkkm78oAtnKAX39itLPQQ8PZf8NitaMxEIhXjeU5wh8NvN39ZTQv+Sa1Vssr+6
8bCfi5wQwiVK1/ua7Hn4kaQIZFSp46TjviGJX8N6WC8AdtUv9RUYdeWbZqVPbyaR
T6rSowGZR8q6ezrMY0L6IOFATaDoTr+aPGYb37OG2q4IZFIfXIHbOwdkd/+xe0f4
+VPrUi0x/kHCsVwRLfVylXtq8aift5M844UcOBO/Sb4x+ORNJafhlbfKA2G64EHc
Gmuf1dTd6NmYtEVPa1XtStdNR8qCP0yDhlXtv2sdOiulL/XdE4PGA7yRHblniIf4
w/cX/rWtX3vYt1TeRDXD1fm43j3QzqHbkvnbURduoG13Y3qaAYaPlRUt1CCFcAY3
cq2zLMcRmcX1Ixdu09m2CH2IGf9JopQ9EsdOfrYC1VYXUgY8U+WgVhYNIGu9e2qA
BT4q3j35kVC7/oniLlFFqLnpg894mGZhwgDxGwMsM39ZZN9N9Vb61ajDI4OVJCB0
HQWl+9Uu/cDOI5na+nrD6+EyTogxabXfdgw+mTMPbxqKwJr2k56j0a9qbkGgcbaD
wG9HUF4vQSmQyx1EGFmJYTl9Ul5qVQUam3WkDrRQfGfQ9P4iT9DIrkDhPAv+eiCn
arDQ48dVEZbw61UONw/fSWh7DnQ/7ItSqVKM0QZzp0KELTU0bm2YlaZNVm5jafQr
HSt27rAehGzwyCOseAhA+cAqU1QGRZgyvzIn2IxxjN9yg7Igt/NKhopHVRMTssmf
WP/8hnypohP6H93B4RtL0BOUgQkJ1pWdXi0eMmCOril+7DxtBl5QtZfFfLq2ypFn
WCNmDg4Gk/xbPt3Pf+30rSMHUQ9q0U+sl973Vl84VdpqvHl/zBWoYnQ5VNVSecOa
zMhHPltrulbrNj+hiftx+iX9akRkTFtxAOGIcF98ybuUaQYxQYExwFNGDWxv1ClX
I68uT+BrU2tIsQTIsYoAz4HE1L1cNF9MjPg1O/cfklwnXOkLfvgc6+z7tE/jSwi3
FDNJkOFrs/R+znkJfK5Ol3Uz63gGzhaXaM/Y85Ks5eehYvAHOTwMWa5uz7BRfrBw
z9fHt2PdUo470SvHTf+UxBppn9f8SoFUphfEGpdXiuw8YTh/e0bl5uCEB3HJQdZg
kxoH2dGLWupotylvBLrmwdUWwg9B6Zz/ZNqEHBUsw+iEjAQ9jxPGh1B/iLa4FS9j
8isHY1FuMMFwps08L5hAMTyuds9bFgVp5nYqHqgOUMkAThFJTUYRg9um1AscGik5
23IovdE1zu9Weq+1tYAYJgqCyP12Sol0Y19RpUEmFEjcgC0tnjmTVIQ+bEjcHZlv
oWa1uVbB/XEo5ZCUyASTIqAv3kdxZh09Lt19b1sTB5Vp4T6psilQlJ13V/niWr1i
9gF2HQrhqme3zgIIWRhPpfCq5mVEDoGSSxPn3qR8tRKuDwUCr5H1EOSCNwIhiU/q
FJQdeQG83Jfzh2iTO75qnV2Wro+ZvCGzyEx1FeiFHXzn6uJ5Of/Tm3tQSRC1ckKm
TNwZ9rNRZo5Gp6OpgKipyVHXNdUCvfZikmmQPYJ5Y8GqZS0ruv/hxMecYShVD5dO
KZByff1eQOAbcz7ur2YHlS8iqDSC7NAapOvxEQQWaXhDiU2BocmHs41DU0382H5x
waPEz4EFpEQibDb0w1wP+dhEj2A/My2dmU4b4iqw20y+rK+6TtieXIGqmTlwhgAT
ubWlmSykO04tZfhs52OPX5goFOuAk8i4moPY0vyXq7cTB8ZdO7xpZu9aqZ6CvoGB
mvrRsorEbKbYl2wpc3KV4wekkgNNNj4QWRSyufJBbUq/oOT/xR+UYqfLPWHbdwFX
nbGlhSkiODgdun6w35VG61/ZIJH4SlZvjUKYjjv76ZfsWVrOZKWCfAiEbKPs5g7C
RheNqFLLxF3uvEzGS0zCz1IrAsULA+w0JS1b79LQeGOxhPbEg2nfzqJyHtrj8QLJ
lnbRYnkWqvAjj3vL5keRLWs5xwPUN0+La9/nxchMeMf/TD46tQhhcSsSMYrazWdW
SyJ0rayNm8sPUOASF4pMpc4QALCM7JlayLUHkd9rYpq4/vt6/YZhzQ8uGmiF+wkq
tD+4eOHLEdzifndvYrEuxh4sOPCTp33yJOZUQ+iaLDAoe+9OzIcUssIKyHLYugPC
5xJ2iaXu2raTYDICk75pierYKJUPINb0+uM4JcQcRjFMXvasyR8fumjR9wQDa2bL
5QPRcCiasTQRBEWtMfd2rjU+YxIOr3Wuc66FO1CRA2HDKfjf/XUS7SbLbf/X8TcD
laAaFyvAmxRwgfVegdoTSotU6VYjQCxjf+dFAdNrjH6Z3E9SYVN8oa00Ox/ltXoi
Td0XiNbbY0K+Sq3g8w3fB9zc39Wwrjf2kUIFD3vIncrRUui47GXZskDSy603L6ZS
fB52zXwLJLqnlCV3f726baxXyKaPJIOOPTEjxajtj2LzinmaDUaMJ8nAloKxYoPL
opKkZ9DjFytHTk87FkzQBE5pkAP8QV20WuumrgPRgiJkKHUvBYSDhl+v09oimSVK
JdkbPaxgBf/AFsdxm2VmZ0Gzuv9ghymLaTlNw5lxECestAsKagRNc4xQgT8+5Sal
zbMdPOfWVZc4wIn1zwUWDtteP9Ojc+BqCuPHb8eNJKDZoUuJtrG9cLAanPxEFEF3
kq+65tWrXe6L2GM2jlPzj67MmKja59octay4JPA6gDl6Da7/AO63RGd1cZNdAPNF
fYuDt9uuY1YKzrB7kTPmG3U8+j8Q26zI1V2jqg85Z7/1m6xRIUcqk8DFQJMVd//n
vC5F07Q9A7OVuvI2bGoxrhgLZvjTnKtR7NaPPuhh2ezOPQ8HLKGkmK9nxVKsG2cI
dpSthCLlrZ6GuJxrUU8GP44pRvLnwpuHorCCMRp06f96KV6OeYGzaAlI2HgSPxCJ
hvyUTt3LCwGGxKD5Oftm2y/ggXHTSVUN4y81dZEY4516EwwVYQT546FEi2YkyUE2
rcQAKmavBCgaV38w1i+cJgjRFYwApuRn9p5b3JvH00b6DxfdjHV1Bk/N6YLYf+t3
HUjAbp2ZtaHVusxlMgZZNjISkCpUfMiGsOiu+4Cea+Q4RdkXJPRhZ8GXHql23gfE
0KE85Q2xYajdaiyUeIY60KcCseZJqehVk0C2PGuQbZh7ddc8jZ8MZWejM+ADFdV3
EKLFdl63GDoSjcv/4txPPZ/HoaXURtktbCyIXgN+my3aekEV8EcAwz7fRrVtNsb0
H5XCsjzNF5xLXuczXPU9ptRiXP0W6xsFma+NBjA1sdGLMlHvEDTbrQMocoqfgteU
XDfrlRydPoYfgcAQ8XEILSlGe2gNoUjNligdIb4guDKmu/HPpQHDqyv/CT7fC2N/
ay1DKvjstFX15y80QOhkDM4FsoSvg/qpIE947Hlg3ez/uoHdEDrzuIvXTSJ4epyn
3eTsp+kFqP60/QlUtL1Kz962aCRZMT0uOuqCf35GiptXNZ9k5YDb2AVOoIoWGuyl
kHvfmJlTG3fnT4iSZT+5hiBv955KUDxZ8/F0arQKbYEcJyx6rRBn3fJvco+4jhuS
6xH+1/xKbTvfC/G+7GW+0PiowOJU53K/6ZkTb56Z3HpaPYKW3nlPdWwxwTgp6LT1
T2v38w0chkPLl+iJLiPv1kMbhWF1d/TXk7AEqOsbb0hpa11lgp/iUtB2AzmEYb/a
TE2QqUoCGp/baUrieAZiLUCFAm39m3vnXI9Y1C/dUBU9pBcRWRkoQm64jems1H5W
p6CPRUKdONPL9jXFG39yokD1S7uLp/XvctAKxqQyreVGmbBr44/9WxY8rtsbCbJ/
c9V37sIZXfNDB5J2oFtzMnNEn2G73auPX9ZjoL73WPKSLbsvtPGkAAbuB6dJgvhQ
4pGLbwdovsANG0YmUceR2wyhOy9NEOoldFUFmoEApcWe/Z5FBgEk9xw8yXrVH1Kz
e5Nqo67OgVBU2SeEGXxz/WeBt8HvQN/vA42K9l6N5c6SxanxiJrpWwj2nHLQGEeB
Z69pHn+TxVHI7LCcyVWeWEAgtwuKAHiGcP66Om9FTAunnK7BhBYRtAtSMQrOeAA3
K5E8cy6UAjVK9jO9S8T7Dacy3TIjuDZyt2QkJmn/R6fZzdsecF3Zmia6o1At25Ua
MMy1W/HqfdvQxh+pcqqbpq8jQ4dAxFub+KBqrN0YKZbJ49+MscYqblzwRZlvSVC3
6kxVc1yvk6PGSEiwL1UfcAzm/VZaHeQ3K9fYCA2wTyN9iHAgimddqLwEeW60Lj+T
rb5uXzbKhv1Lj9+G9rSBvEo2zMKzOVOGFjUK8twnUJcFtFd2uPpw+BVCHsn2x8i8
wN2XpjpBGTmDjoFMLzkDgEZi9xWk5l49/KFllYpscE+EOke4IvU4dHMt7yqMWNZn
grEq4lWGWmpjunpNrXtqxlsUIMjneOiGMMav8bH8Id5enQBR4lioVtWIhYl+zskP
P2IPo91Dg0qXLchZkN50/lqE1f34tWeusIIhwMJo/+dXiSmqZSYSilm0knALWC+V
GGCCGvPRYgzYswNu7bnEU799e1IHU6k5SHN78enssYc5eoo7mTPyKxO4yEQ2Vret
Iz9I1gzwz+yObArAj6cfScXH0UwW8NX6mYpXxzkrlOrqBNo3DAVWERMGn3/1Th3d
Y3N0RsVjm+e39I5Bzr2TqbSCSy9aW2QvuaVjLEiP+5VKJeHx1pZk5HKADq14xQiQ
KePqhUElMZcgAhfBLeK7jFQhyhVfkoxHQFHb1H9eSJ4CUYvvB1+H07U4uGqq+m7S
gpVjQu0vD06+sT0G0b0QTsEaUAN2slG+lPxn7rnpgwKVi0W8K8SPxsvsYi0QvntR
PpD3JIBGyJSBqUqsMomvGyWKC5T/ci7uZRzCChaeWlBXI+SClKHplipuSjvx5pUV
tITP76/Ow4bqf6GIfG/W8JaVJy9eihVTHyzPncwrYmTYZW70Qc33FEBA8lhudlRc
3sv+QlJD2FLIjVVOKURj8GqBP4l9DQyCOEFTTEof7iUE4BRhMwIvRNqFG6O5Y7db
MLN7ezs+U2bDe1TB8T6Nk+GewM4HUZ21FxAdZbvTsHG07eWSQvAhgCYDvW6uICEs
pfGWanvEuF9Ikn8/Fnhyn61ZEEwFl++I3jauQRVSy6mb4k01fF+mtfujuEdqtNy5
h6cc3FDU1pVTyr6XniD0wGjwgzkJPJxT+7HBeJP5W5FLW+hNId7JRSUJuLcDxfFY
2t/FvmmxFGe9DbkqB2kP1FYglikjjl7JiWiGlYwWeENHIB9JCNWRo0288tvTiqst
EbBnheQBJSjyO5oQIU3D2ncLsLvKHvTw16q2RwyHQ+n+eawihIkJUq21ICBcDMRA
2hx6WY60/9QAanLCI7KauoOcL9cIlwkJgrzox+Fe8YbAyS3Pu0rhuGeXwltFPqfx
qxyAkMx/eqMdxLKb+o1PVrrBKenmxGRjC1BVPwZL2QocndL30YW1D3AFJ1bKSaah
eOThEkfdkFUf2ZLZfLdY2CS6K2TyOeFsBbXOdyeOFuhcFWaqsJo1o0AGce5AkoHZ
+Sm/XuHsxGaJCPApIrt2vGEzW4EVRLy2YsJIwm94HIj78FfBo61slS6bmkMfVmWW
52FtV9cNllmwBEsbc2sFOEmzpmIQR+Kio2GKZQJEObg1AXcI48KjxeGj1TyIf9bl
CyP464sukRrY33bVAbvgqk7wTO5yo05GY8puHVLoKdrCxmKVkNh2xi3HEdjC5dtw
QWTWI06Glhvhyb6TKF+a9Qpx7ceeeBmnB6CFco9Nkumd7G4sHXKH+JIDlqsMve/l
waL3SCGEvyh3lmP8vSYWspM9Yj0Qm7Dzdu+kTu1dXDFnsHMr3TGmrS6lSxxvxQtO
SBeAdM1vmic0wsbXpwFSVgv5kEmaUCtnW4VD6clICXnIjD/fbT5XBL4dG3OusdWB
G7uEqIV6d42aUpXlyPE9K6ZBJFG9S6O49mzIKR0hrgy8ck7WEFSVAlaH/YsSnrCF
alHZXgxuG+8NN3dqCDWXmNJdXxft2KenFMquLQ75BgohN1fJqaXaDLuGc+z7E91G
rtnt7w4V8FM7Nkz3nBflJ2BjmuHPkG3Q9WlFUmre5nlNeh1ht58hIh9QiWDrrLFV
PgWjXm03YCZRV7VDBMGHIHmOE8i5HIIo32QtMcw3GlbLqXRetqf9iRpYQm5oHFSb
VuR2sHXexAojSdqoEwDz9cSDRu3JuIHqngbmLZKlGgQj3FD8j53Sbd8s3ltLx20C
HN8Q5dhSieZT1bBCoN2ctyjJABj5Yep79bHtexMtkpUKFm2fjImImM3lMkszv4XD
Cm/oyKVCdlTp/ontjcbHfCJEGX15CB9PsWanc8TrTpWdCg89YtMYcgcU+bBSbu7+
GjswQkZpvby7+s6SrMCf9+vwT5QJulPogHeF3fNkuZiFvI49VlIUv1+jFSnQaxn1
1VxavODABFPwHefNGiiUrCOxW0hYjgysCZ+LxcEclruDp6N0nGoAnk5bG0eKGmAi
velOIn+b8JwPMdC5ULN5DDWjFwzdF88a0xKG8V+an34XeCWjITBoBZ8a31jpEX7Y
HvYAw0uFsxwADhDBHwyBwSfshnC8+ob4+QiVT97oYzghJYweeYlnXH0dj4Q0XzeN
1XFYBJVXSpaqcGSJGo9GIyV+mTXVMPq0dJP9kc/wyqSH3MVWwS5kFCc5Xr/eVuw3
AIGdD6ry99wqtHvapALK9EcfuMesFnH59Q0dsYBNWUpVTjqnEEm7bmxKZPyEMyj7
Z/NbTfRKTtl6L5gJkvo0jVcw7wTBWQPw7vJTg4M1UVDpKozYXdgMVx0/2Q/AeGLm
Kwla9JwcSVYs5R5v9QANSRnHPU/Ypsq6sB3jbTc+QAAEhWw77lVLly8/9Jm+w1Cy
KaoZszftzJCC3AtsJ9B5qWWdGRY6WPpmX7CSlCO+zahfyi6e1JGLz7k2nW7GcWKR
bOoFOxTtYiuBwSwNpyvyrwTy6N2s8A8/Skx01wZvXZmHI526H2vSa3vjMvkxwMoz
ZapVJoEZgHiV0wAc/tp7HQiwAZmrRuwDdsQAyo8VtxTmSvDEDuYb4PDoetcfkh5j
Tm5Ubwt3gvxCN6xhYcs2vsZmog+tT7gfSwJQzR686n0vIR4g69F3fwK/G0RmzGT/
aVSXCJ9iqz/BxRbaGCZ2he4Owlq6OOXltrWsFyMXy1VoTGBWyyMSp/vPTNkBtLJw
Ykib3StUeLOfFK/esuHyqomIm4LMZR20D78BDGQuXs1rIpZSZqZEpZ+yqnrF6VDK
xMy2if9A7lNMPyH3EfqfZ/y7Bjf6gLBnscDAtX6E+KR2T9gToColUolarc1oTMJd
l93MEYcIZiYxlQ4zAolZWf95w/vwFjzPo1sVIluRUplDQczmTteD5rv+zrSvm5+I
kE9iVBe/JfQU8nFTG6U+gcbkmxDTBJVTgvhgXR9JrQKkqqt7tutmsqPO6IoDv6pH
qa0oUnY1HNDYa++3UAGXqajsIDTkS1XLjTUen1cUckJvsxhhGaKXpZKMN3qFA1/R
Vv4YZjrsg3iefwHhvaqOT33UVXIhRTjvlcJPb/qnDL7hx8wIjo7CKS2y95FvRAuK
CzhdfV0AbuzumLuSd3mcZLS9gZJV1LJAAUVKaEocsh7V1Mq1w1j9WuxlbSUVajjx
5O23W6z7wYMkkuIMvlIQQaMutuxf8g8Czx5z3tR0xLnyYDrP/sgPtBWfHMlb1mae
2+51TXka9bwNa3f/RTO6r3OdOnLmKCwjbcB7O9UG4oLC6shaedHS0c27LOrESR4w
YprySswVXroDT04T0xFsyofod9aMchTwkXugxQ/4+WnYrbtzQJQybDYO9byv+kx3
4g3WLxwI2DEgvO6hANKQWNMhbcXvNPBAn4vNrAb9cm2tYFj5nn6AklaV94SbIbfz
U2BQOgzSFyOb+ureeB+CyuLZCaqR7ZOz1DI7WHYzfCV0MVm/F4kjKJy4IOUWJBhP
BP+sl8RPxJ8PmIKWgiUSpuu+RrUWgFO/3knd582JKI5hpvtdnK+Fm9NURgmkMxEB
bcl++nBE1cCdTH8v/gk9pPFU9DoAaWc3oQz6xHX+jJiCJZLMyhhAf0WJwbZmiRp3
lxSnoQVD6oyh7NGoyLBQrmUBbkXtQShp9hy7sZZMjHZuZz1g5dcYFN2ckXNFQT/l
U+NTHvqxuw7wDEDpjBgRgAIDRzBWnRw9XBW+kS7gM2s02VQnFbJnnSjItKLaGtlu
QU7QCMBXkC+6uZl2XXKl4yL7nzhe/2ovhEe9z73nnlAQYpHSP78vTddXMfxw/AIQ
aXW9hk0qmpuv2ZXpb6GS94VSnBs5GNwm5NBAxP7fCV3gccM/nba1uXq77jot+sAl
H9nwRmrq3gjeyNSlbUzv+7D7NIuLVBG7Bw+V2AaKXQugLJ/BcUWlEQOjjIz6hulT
5LQlGLwLh2fVJ88EcpOMkWYk1bmw5bSwsRA18D38UEDLDEcTYhnGMDHzzZkJFOgI
6k5YkOWoMJhvYFe82wzY4BOX/IdZ/yj1RjxOxjiC4GUDrhu1d0rWu5icEv8U6yGT
byuav1SFWQdb+fTHsZjzay3IGQYo454rkPqugxFdFaDg0gdqiAgfIay9tjIO/CyM
uWFZFu5ZS+mbczUbsFIjpaICtlyfbeFkD6ssZqxxVnNICc8GjlGKCXqlO4MkRpqV
dNa5ZxUbmxRsuRl6R8WkgoecbAijZkx/9a0dar2gT3uLBXVZWJsZQJ483YO95gwj
LFNsd3b8YITfvxdbcxHHY6hu8s+IPyuS7ycjpO/w1mllYd95UkBcgMZku9vq7URR
zF4E4sGrjR5+iieCxObsQept+SaKb06u+KI0LIY/iJoPLiYWNvE6idqJVMDG7vXR
xnaAtZbF3yyJFCio/dnAHp3MNfkIYvO9QgE4mDold1+BhW+FoHBP6Nh6jIcBgG95
I739pVItWIvorjMm9GhyssQ5Ftp17hiILJGXsQXC+yFpIoZfXyqHukEXfDjfeWQF
MoEkfN4GvwyNvSqShLEKy+ygAWrRX01o3xPekboLfVoH0TXfSUdCbq0fqhOeY/o8
LXycvtnekaZhHhy9x+9VTyVkiHs9wZZ7DZaLF0ft0lKV5U2FYoARyb1nTXR/TPTE
o8VCzoqWkG5lEoKOJIkLltX48CHC1Sq68/2GiMuSjB+15xm0EAQ7ZV6No8G35XcS
H7csJPC1UXFi4sZoitP+8xIWg8X+zURvLRFSWHUGc7vQmuJ9OO4qo81gJfWBVvzs
Mm4Zyi4DywkM1L7IFgNiVP4nIcmcJw0DDnNgQaAFsCYj+0U/j3PBRZJ2/FGAuc2O
FRIHGf+Ytgm+PelKLuyyhCDTo22l3y/dlJ5EskUkeB6SdTGWj07nDlGi4+2/WUo0
dDPoeTi6YWTxzhLhqJAOvXTNz9qj9UmrjaXhrJ+PFz/UFN98+QNEp4oWtptRCN4h
Cqy+xZl/cdJ1rndZV913tvv5QV3MIGN+Cm73FT4kEgnyIwtJOSC1sSklxQ2sgMwm
znW9BGtcgVYJZOX/ufkgVP65/X2xi2SHoc7bmwyy0h/q6xPXVziD4egAaxJMp8tX
kXuek8u+4EPwQYqSad/8MkanqvDitRlOIr6ARx9NrzuJV/GCMC0z4j+D8kijvG1J
Jh7LNDl+a38JoebDFiejAUv1KtLtIWzAcb+kJloV68hzodgO0WNsjheSd75MtPoF
Fklzb3XgTWMb7xVsmYK//T8dj6H3Lro47HL16p0lNPi4NSD+tdyeiiUiiDgyk00W
sshWMoARzKXnV9iDAndFdqOiR3n/8FLT3tzB1urQO4CSpRqEs5CBctCayaY+EG1r
TAIcZheJvkDJBCfAK4D7M6Pf7JrrHpDcITiCMnN7b3+JeMdh2x7RPaBxksERIf06
FABowTDAg92vYiBXTEQS1RqTBaAfzeC2yoPLtUVmy218UEARwmQ3Lo5nBUhT+2w4
OKWi4++7Ehf2ezAqAoGwLnITTrSiDIZRfTcLfiIdOSdzVQC7/tbgMOVLygG1CZbT
LmGlgQWGnZ18ICXpNd6t5URLBYZ7p7Kee8H0EWw4Li6LjieE5IG2LeHjNGejvzdz
lo6Z2nC/Ok+e+A/6sMcAHKuK5wPI7jXz/fJHYqg4wBVRD93EtzzIZvculhgNqaAm
sBbKPeyz4I4Of1KYVradwWadhOrwF8LC1n9HVM+ngYDHG/w23df6vFCkPBUtKLfc
+EYtlBhPXFg/GiWAFrggqUrVOfh11BpjfcAeKDhYUmrhk1nRCBJPqtDLYBoex2nT
t/8r3RftTGcz/AY1xO0g0Q4UcHUd95lA/D6OLZR1wuMZbqJvo6AabKgtic9w/5rI
QhSWXmdCmBylW+t8t5GyOtgvYTQSYKV/rwFpR7DmY5BKH+kJcN/f3kZutwPGdkp2
MukCax73U7PMfxCv8WSq+vCT4daijBjB97gKvy7G7KzjuQSACWG6sstH65JLrQ+c
bIuenVPYFLj7kyqa0KpCDBrGbYX0imTZe+QXTkFR167Ob09fpKStiQ1Lce3aJvTA
D5JkF/wM+LyrckrmE++v9oOSdcJgAh7h3heonqoiuHzZY967EABMT/jOMwhdM/mN
qZPGW36SLTgKewQap37ryt0QPtBWnosYpsdu8IUFsa1zYqgjIl2Sbmj17WFRrew/
gMKAojMzaBxaaLsLOdVKQ+wvnIAcyAccA4AWPXfVTrfx3PfQi0ZTPNwYYonosYdX
ixkib2x1P0y+vOUNU6Prg0qYm0bAe41zKwjTtbBk+aKHPb56s6NDwgyXP/wmgX7N
XaK9LYEPugp5VAkp4dtXc9T6wjeVMGr1iEJl261ZhD9ATQsaRG9/eRF8QjgC2++O
hmZBxZvcFM2YlkyXnG9v2QVNxhRoVLIYTK0gmzmbaxu2YPQE3E3o3J6slrz8okXN
h1LmRD3JXxf/KNWAAQ9HkRV8LerD3Kqs2jXPf816ts9rwC2dokRTtm5ApPbOYQs6
+8o+UDzvxhaAYL4tGGBzlhA1LnGMMCvOY6q6CX2jNIIgOtF0EMciB/RNayl0FUpK
0SUC4trg5azEvKw5/Vv39V1FvtLw//n9lySPJZt03gRToP/zI3A38BrYf1KRLHLg
SoU2EyJ3bNHJeAtn60MtCgh4T8a2Y9uxwTXFMRduOqZeSlTErqn/PVcyzBBKgz6S
TAXkg5/KsZlrNtpb2qeiRR7/4Z7xd97UQNKo6Dqj39+8XcTKtmOCDuNKIwK180c8
Gr1iJppMsSJgoGRk7P3nwOUxheDhwXDlR7SWVXshAWfOYCh1T78pSIxfrAlFNUk8
zcFf8HmKVzlwMLTT7EOCT4kYChv1tKb84ocLZ+3//10pNJwF5IMQRMsyPwxgpgaV
CojFLj8+A0yl/UjGj5O4hA49An0RjNtjN/qlGeZKuKW1+to28+HQirP1aOtGJSfN
iv0MbyZ9yriiSNOya1dY1JRQ6P+pSeLByENCaVY0WyR0CDQ7bPgwbQxku2tc3TLH
jD9fX0loXNhtiRMU1Sh1r7ktFE/ANLMDuowNOWXFTH/KWWkeQIB1tNvl9o3gSSNS
pvu69wSUDelVT6SFNQewh58mtBWUIHNGrJND/OU+b4tk0HE+H0V9zcjamXLhIZ7M
zay24b6FHmK2hU7tlbMc4j5xBgoYx6s8BbZojidhgazoJYRDjJzSyCvauiVqkahe
L2bqg0yM7okzuRA/h/yvo/WIlCqkGBM9wn+AzSWrEIhHlD4PFLjPj1lBt0j4W384
A+xI0hwP2LP8yYdx6v0jnWUqH8XGXvUj45dj3X6vLK0QqpBOqD2xOr9rWuojOi1J
Au5+JTyd2pdpMNAVcFTaUc5BB/vMBLNawA/zqIQgObIUG9BVgahjk/ZZZ1d0jKFy
c3hqd27iIcF9kuwrouOJhFh+psCcrJx5QhkqjQLMEwnRM95zQI/0l2m6oUwgQH7a
g3NaScCdAF1dm40EEQEU9u9zpoFRf7uWLwcFJ7sfoOjFrd20hLaXiQm64ZQQAZr6
aJFI+9ZHscHNQ+HoNJZNatvR0gECoT+HeBwM4nTQRl3E4/jt9BMkmf1aokRl2sfN
x132/pBGD89c8GzYf3Kz7GO+grzvggZAtmgxipHpVq6hjioYyKqZBTxkh4wkpBO3
FuNNuk+dttzyXy8WrtUyHkegdK7em7vCV7wBHFTm3xeac3AO7DWyYh2hec/Fs2+S
wY1FR0ueHGc4+XzS7axw/vLdRew7ZEM/o2wzUBeoDpRuUEXDG0dyURB4F0fOsIue
bgDDcqdG433Geq6XoAGR3qeuuycCTNgXaozJWw4VoZGUSTvHDizqLUQSXzvbUEsW
Kb7h3UPQfJi2JIY9K6uTRog6hxOgSSbDmFOPuxdkZFmPs/nWK1wd83q8SuXNReEs
oUqI8Bsd5uXPFH4TABK1NP/q3XhjOD9As95ldNcW//yLrEVRthGFLT5IIyNJKpie
yVdLvnmT1ATdSpqhDU91ET8pOZgJVyGy4VKnhFkQq2NtKlYiKvW42sp4BnoY7AIp
1tik6P5JtgNMHv3t6vNG/K4fRxGsHZsfSQjCauXddRu5AuQrN0VRcYNN/uPKUUI0
JkO5EJA1Gw8AARGRdBCq+wqnawXB1kKaS2Ngp9+oNko/eR1Z9BzxtVPZWLLsRoDP
NaZOP5i/juPkquM59skGJxOdJ+c6NlMg1TYxcf2qiJd3BqlolHK83r/oFga2ca06
JJgw+aSpBW7+VB2esNHozFgkzYKzwr6ar8No0+5yiDav5DlfnNk4JQ5PcFIC+iuX
2ukdBHFRE2V3ozpIMvWxcKOy9gQgvP8K6n7JiRtRZ/6FkT3N8MPpjUzSfakV8ES1
w93Kd3CCCyQ5iupAnvxgI2CFtTZD+F+r73NJNh1XN+aRqoQxmA89ACpZHO19ap6w
qm4rnkRAgUAeTrhAKQ2K9YKU9+vr1WlPEW/cK2AtYGJIGGVkfYRyOwBQHJMabvRj
cGIHlTaCvAb1YWcxQkLwMh1VP7fZ0wd1p9g28fiG28U9/VpZJC2aObmZf2bv8H9v
E47Rm/uVmZBO2ZcPmHlP1TZp7XYoQVYbAv+QOdMkc1gYSP0rSTNSd0eXH4skjFjM
spO6IiB57vEEjrQHilaraqysuhmpDAPCbrymCOkgy+YOXd4KxQfbHiyUmXn+aO6n
MBB69J1vaPknrbx1NdeqIidG5BilTxTIA/VozvS34CvWXALrRpj1/O8vzxhjDgz5
XMnCKi1sfd1mIMxNxEKtgxOB2xqjVKlUE+AhmeU+xbeop7l9RFV+xJkz98LoLqUv
5nqSLOu0C+nXOsfd/CNVfJ9DlWoKWqtLq5gupiY68X0049xRf+A7RWYiISWjPQQo
GX63eLsT9qepEutLTPm9en09SSr8zLW1P0h9lKmSDixWQgBTsgJalCemU/kpE+Uu
UhtZkUNtYLLs3lzMe3i8ZPEKbPBp1EKChChYx7lh/0ZfdkDdzv5BQWs4Pihetcwm
Ue7E7oIr3Qo6WrcyT9NuEBv5oKS9+vIgYeUBfuK93X1JURpV0wP2NW/j+NpsFqBi
I/Ze+mpB8oQ6LNdUUCJQmgYlP08Wu+HZflNsmzRRD/UINEtLghO007wszMYWOjq5
JHrvmQCoxFdU+JwpAE7mkCWenbs3XtKVt2ILS6uDdn/izd170l4aLkjf0kwO+rz5
iX2S8p9/LsEcmnBWIMk/THtvSdus/ayqthssXlm0ubEerqZbM0uLtplRYr2qvq8Y
8FRa/I5lsthP9q0MZ37tBRgaUQPq/KlILFQfRXl4MZVNjrfwKLnTOkqljgmE0mpz
oNeKSqLq3LP1Or9Yw916Eaasdd8f9twe6DkgyGjiWnEKP6nZ/v9A8qx/emgYbG2s
hRj4KmNQZWAaFlXk7hEpC+7HdZj+d4IMwpuvUvxBQdcfF9CmPCa8V7NRXqiT2pFd
VeqKuUbqzv4hanbTuGOb9I+5D55yZSL04RVrSPrqp2toRrklX+nVy7AxCO9cyOjl
wi+eLUjrzgynwXs1r1ixZkXFB42vpgu7A2dQUNyrFbYXEo37KPth/fjBQenlz94N
IzalLsqWCbD5a06HD+2ruTPQ5RZtVIShv3PFPu2GvoiMayMSuPGCZZTdf8WFqDh/
BxBNhZEELGGSgGVkHHyPbjhVPT7GYXQCniHvl+gM5jPnheXZWOgmzI3mbQkSaAt1
YHvPtdWSgqdU2HRiGqd8TaJcPAh8KLL8y3QyeyxeADZ5Hrm3T6bhsDXTwenjcWI1
cYjZZWyh9Tn1NFmhdrIO0zz0BbkVrsQZLP/c+M9aKF74MWqi3pLOap4xDmF4bP8r
gtyh4WpX3FY36FTu0Y7cwkyrzgJazu4t35MIP7uy+XsqrihJU60Y7JiPR7U7vIDB
/Qo0CobUgid38F9OQoB0ryJ9BYRT8frJLXkp8N09oVuGdGpwtcRlZbKh25s+YZO+
b9IHDdi8qjvo9lH2Bs3mxy5VtAJS5m2uPWqE0cmpNn2hGwSzLI0s1Oa4wmrNUaQj
9sQgoFXmIVjQDgu/36idefVLagI7rGJagdrhhQOVMGWWmuM0/op3reJv/J2LiCnC
Zo3U9+aJ64MuZU9k0Gzg/av2SK0WQfwjmuOeILJ2JOfWcy9zGo4wrCMc5Knog3/q
PjoB5UvYPaIze6c/4CfjEG4u7P5u8YufmguAaL9Pgk8VZkSX3Usp7FrjpTsecEMO
dFVelW6QbV80oz+IjNYnV7Z9FMNY8Q4h3Gqw7Uz37JdgMHbSgOJeaZzfZsf2qTQs
g0jP5k4v65k49+BM6F65a5oqnvII3pkh6oOV6njGP6RHjr5kmOk56HyNMo4Rr0SP
yWex2k5HunGPd9fkj9Pq3Y7/RDUiRWclr5+0VlvimsSW2fgGQZiWfFSXcB1miC6Z
ym85ZsUc5/3o6YLcC58r8nYEZNKGu5LEIcv+w6MnkdZ+IIxfhasIYxhQnGZf52pZ
BrXVNMKKzF50fToZWAe/s6dfdY6ImDmxKV6oujrQ4ezr+5A7shW9tj25/VNdYPfx
51UYztky8Z6OS0J6NXqBrMECHr58liTMZoQKD8s+NJ3W0EPslCljcwDxW36SadVX
guQHUK6Jk+tD94noXr1u8zWbk2nF3TZTdRHJxQHIRRnxYuqBy5x6Q7n2/W/spNf4
/tWpj9YvBSQhqhf4IYPLBXNn6JVhyQ10ZzwI7whPUhjTQ1UFc4S4Gfs+yq8jiBlT
cftfIGinrxKKvxFMpi9PlYhu0+KqJTeh6c4Dxt+wiSiU7VzvF7LVieUvsvQ2Mqt+
Fd4KivKMXW/NgHBHIUUhuk8tAixDCwaE7FDKZVQfTrvZv8Egba/7Mj1aLoSieDbC
y/YirXtTjnfg8c2EcGRRFijPuWWuSjT9bWs/q+QiiVPFvMhAk8wh3N04LkvKDEa9
srP+fWaXqTjWyR48FlRbkag8DMJqIfdULSQqTRBbnG+c0Peqt/IMCvhu3oslzTLb
Hgz0I20Fe9nnq+wZtZMtCUtFlP9JD9yE+MvUYfA7RIzBCZUaj4clZT1G47CWqUSt
QRb7Qqvud5wTPkDgQLFanJpeiaUmUwXdJNvRoqJ4orTcMO5TlkRzTqD510TFFoqj
BFRTnw3/wWsZQhnyN9LUeSra/qKav3fDjcbfBM9fHdmRvJYJQGUIq9UL8kbqIa/U
w547OFLlTK2tCCpDdHwGy+pBdy12LfNCDUI6O2MfTNdKSK5g9n7gSuxqR9d7W4W6
OBCDPyig719KTos2LS2AI3XeAMMLnoCEr/9vGCOZL/Yp7OCO/NUyqlm0Dn7/WHZ6
1Qp08/+kf+Jkf10ZRjgwJcH2jm/IdVDCdDB5yRHOmk7+q2pF9nZYuf03u4GL/i5p
8A8PFyamTmxTNuUPnXBhUXzX16LBiiQNQ50Esom6bFDRm84KDYffDiuk4mTpnIcm
P0GxPzl4Jgnve3z1CMJ/LX/WL9jUPssdHfywm+SPGkJU5gBlPuLZy8H+MQKSyMel
Mb0mo+OcLOrFm7tqTITYUD0TavzwQb7ucULItmihlmFmEXseUDfDi9u7jmRKpjz/
WMyq/23M9H9q9dfGHJcR7rlhuN30J57Y4bORWsakW3Qqu1y5yv66XknxMtIC/LxF
OOGU9OKffVCw5bA3Q7MzPptiacOwaKSiKF/dQFoDN52EUCs3uR4HgapkwDLy3nu2
AykPcN1K0NwBhJdkiwhAbjR5XCBvgQhTYOmWkAxcndY0G6OhmKBRlOxkrioLYBb/
XFNl+qdacFld4T86CETY6qS8Ysp2VkBTQav8cClL/nUuEPL50xZ2xlzFP2gBrkvc
B2bph4UUKSdCX71t5liasqWw7sw0hhYriH3l9+R12lY4KCBlv5pfeXk7z1P7KZ5W
6TUvCpLJGDi0+00ZSwFdskL33uYOY+0VCRvwmeoJYUGxcGNE/f2psLCjhPr4qqfi
tqUVuR22bBploUTVYpVIVBcqcS7NU6TVDcQxsuAfXafs7M6G54VF0RJnf77VBuH3
3yUXqkhKsvxW3cPWre/gFOdbFufxwbJ4bGQDYSqrKbhUGCBkuDX9mKPPc6GdHokx
3ei50cucH2mVy8MAmOccBIjTVlv6BpFDGfnvX9QUTwsznek3ZAdxulKFOvD5IC9a
j7sgVMo7HpcK24a9sge+eru/RLTcFVkVbpNqdWPK6lox8mruO6E9A2M33bhWY5t6
5tWw3oFQG/I+wFE+Di2lnztLBLZmAF7Uh7rpVWErBPPOeoI7sAzfel+aZqiLABQp
imLx+hnzyMQI4Naj6V45SfY6+gAveEokhk6t6NeHtKFWpUzk9uMZsv07mo5hsqde
qNJFOIFGshx0NSgJYuAGL687pon+e0SwRDCR4dm3av+ONDTsKs+XCxo0ZGn/aDvW
KRNHOuyxjv7YivUk/WE1eArQ9nAPv+/DQXgICArY9mP+lL4lvxG04yAHaG4zdbNP
nvF2SMS7yZi3A5gTX3jmmwBLIT7ksCxCilzFbC+HWRqCQZEJSLVUs7AqTl/V4EqX
yoGmgxXP46SkgHZ+cPMzx4p1MLVPncdPwwAPmDEWqw7JnptdRsfMst0f4qW1j0zS
0WAtaDI3dSHQ7iOmEirHHzIxBjfQZdNntOUSWWEVTbv0VwfDzJQixfaVb2BYZamN
Vc9nwJE/WG3S0CsgQaypGVEVz85Jx6tv5HKceU8DX5GJe1qbkDyLLsebZdqGfKuZ
U+ksR7EfcW3eKwv29LIcbQ3+mZI74Ju0d9S7l8y6p3DdZd1eVpLutExDdFvoqjhY
CUWsmU5gA1ClAEEdMDU/UFTiiytSxxMkmfZOvL6ZwwmnbGWPqgCPhGWvTKYQaS8e
7VovI05kS+HAtnONa9+bXivXKzZ9bJ+AjY49hCVUHi4ft2vWVBBnGTBNfIpDICJc
lPNXYMrKd9zSj/Nlrts48CbOYBg3Y7EiJ6Yi+80XtdwcQC7xUFfcVjhBFCkbu0om
W5ldmNnBXko9YlHBMCpDqnPziu7rxk8reJptyFQsDa4s6Imrvto9M5TJhFmnGdAm
ERBgAldRrSSg8KBKxaRpvMQr8grVAmwEV3NtfjqJ7VZTEhvYnWDsHTy8BIwh/waR
5R9gtxYGCxQTmFaQLepPbDGQvdcPU77gThpTpzp/Y9FNfigWi/oYM7hmCWrIpSHc
Hm8KHl4pWislyycLmqu77MHhCxzDAlteEOd5JhNPuTmtbu1QbdsT9qXJgsISfP4e
T/m0G8dUGNoFk4zSVg6jNcQO8m9t9WXsNC1YyhPzey6N/q4rRU+qTSgIq2F8NEgx
4zs/ngfYFwissiWM+qVR9iqYSAEQ/Db8zCro+QZ27sAoMn1MjiKm/8KENxrkVC+0
Mdd1fnL7u+ubjFEJ6sDV5B3dbHTO00YOYlwSB7GD0BF9RAUNEoqReXU/VGK2RCh3
YeInUBYtfMxIGmTFwAWgMNFyDfiArcP0Vx4i0vcxzIsPTtZR11Ndps6dSBWKnB07
w+AujD+QkLQZbi/WIce0kKjuJeeU2XRrFEiIHPMdrlQNYkcpZ4l4g7Vhc7wIxD0p
W+AgvXIlD7giRxnzcS+WDT2dg+QBzSbsH1J5cTMyaS0gdvvrq/Jr2hV7VqUi2kwQ
JcXU2qrpScIRiLLKkI1S3kBL9YuEOC4jkvtntb3qQe8vVqn4U4aEa5b/swapCEde
2aueIFH1EP5l/b82eZ9IHfyoHzfSVVWGYwmSN7sJcDbHs0fUS2a7MTRDb9PqMWmE
Ilv5p10l29JfrguGpy50akhgGFq4ba/4zbjaAzpK2SrL8D7gtNwuUXWfYdNQKqEa
Slpt2IAjClD2X1IwnASbf1oVChTHUCUbjoiv/JSIWXxA4YXXm/R4+x5GhGsDl9+F
3or14T3vTvdss0wyI8OirJuTCRZihh/JTSmkU0R3n/Df04nL2Cg0rRr1tfafQh+v
Q3OqxLYG9I6y+PAFmbtmEaODytmWFDKLDdhylD2UZUPCrLTHGhIQHVvzMuzjl5V/
mKq+24oKtpIj1EiXkKEHcbQlDWc33NVi953R5fAbAeUMaUJZQKkq0a7vwtki3/9d
BPb/WRf14cHRKWWyoGD6sTFOjcPkv3BL3ikWq/P+yCmw3+fcvnbprA1Lo2WVHUzP
PQO380fwXNvAWkF1X+gexVOH4QXx/jFoOMutRCVexTjfOFCBynYuIpgr5vQI92yW
mQJxW0+gI3rhat39QhcHHLV8KAc8FCnWAKKsG3YzJzfOmC9Zt6/iyIDg680B/A0o
VcFUPoiSJiRGRq5QlAZltDywKmjQsD4O0JPfMeOWOmcaZAYL0nFu830tgoGvQehO
jc9Ji//tyIdBYUY8JF7C1sIzXLWgIBX790NMSwfjej2uS6ALCxvst3VLLnXZo5s6
XgsTFb7XkMk9+vI+fG6WkXDJEJROI8HlmOenu/cGCJPYNzb9rOndb8M3F5x99mIC
sYHjKuEP7rnWs//XJ969pquCRLxnZjoO0bUW5504WC+qSeI+nPwS1GeBzMVfzpKH
r6ZFfxJeFd57Ah+kHatLTRGKUUq8RMn2NLBGp740XXvb+ZdFj3RkQwQp3M+ymJ0E
2LmH0WE6yLyq6jBietijxooukOg6lLXR103MIsPOJbGaw2eCgrpHvWqGTcm9URx9
VAYgp//6pLMcUyYHTJL+l8ieddK/Zxp4ZJLNZ4XJOlTscZ72VLXIioleVMxeyBU1
hw+k4JjWuQXfNulogpI3ft39q2fZcmAlMxR1AuzELCM5iy8ovJ/oQI+w8gzR61iA
r1Z3REbrn12QB3TzWdr67fIB4fN4eCY3P1PJISakU7IRVUL9iAq7KrPtQHti1STC
pnyDxdEucX3Pg2Tp7VXLcKLjl+jJAs1rKPtk/qKCkEMgf7wi0NDYdWdI7oGwkwZR
/Jve8uAViwz3nrMwt2ZtWFcFZFYAyaEekboDS3XTFAH7dEf+Ps706V8y2ls1sFiM
SP0SYg34S8e9pE64NOir94ZvbEQoRk+8nfpv3H93B6OZIs/qVVAAadHgs184RAF0
BkL2d/5jWxfgdI6kinG8aCK+3VyIHyAtCmLWRWp+Vb0lCYHTr07BFkwGn897c1H5
vY/Q7YKuIt8syYig/gQ/a3FZdxQqnEkt810T07X2FLW2IXuQlATOTBDUri9SU+0b
fGhASgXWRWFhYfmIsXIbRb6vGDI1IZ+ZZjhu7bHJPhHXu/u+X60CpJSOIZnflcac
DUEQPNsRYVWwC8kX2CboTPuJjuPGHmDzvLrlRZzOh4RYBHeng53bAecv1YAq2yqg
B8BXa4sMpnEBuu2mLfzt4Pf0LtqPXWGXTlLPJbIdNUWflcY62gJ7PZkR9cJC1tve
7VuPyONUHUfPIcrgi/HRJOfCeG4quNKU+HlZy8FZqw1nYo7ejcLkYuLBeygkZlOm
w1c4kb0kPQVa4pPSuVhjujNkQmyDqDRK28+zT8+fPC0IdcXO/Y7t4emKzANg0NA6
WhsppAe+5nTsiTu/AOn+r0JsuxpAkCus2uH+IrWbtLJX/rj00ucmiPOmEELkPgep
R5kunb2aGYpHNgRxE3GfKLu6zdvvsWnfm07cnX7vVg/Yg80D+cC1CLS4TZ59NyhG
hHtZKd/Vyz6brL7WPtRxnbFDePAv4SuU1GsaAmy15TMhALsxR86BmkL0OuIEfo6F
w53B96Sg4j4fS4J215R2miV5lXhJEhXp/Usc+wgDuOPnH+KQnO5KEVKlblPvM2ne
2h/DVAcqluMX6KQS5ycee5p4wIIn4XyGt4Rw2VOS06kaKWlYT3qGdpN+uFvR9haH
LaR4BAF85/yYdg5YBumNC9h2rLWhZl6aSt4AXgLRAwKYn9TA5+nXL+1CxkskYQHv
of03+v1U2YDa1WIMl1Burt/C2Bpul5ERFRZRtO/x0MifWV8c6OAAIl18kH7iRnHF
XICmIOH1IueQMKo5dBvkYXxTYSz4Btjji5Za6aj1yChSoWbtlc9iC7TIMJGEtYzp
33pnOgT19LS04AEiXPofyZFLhgcnmQNPSXebLN9U+CnKItJbTELU4v2hFJfC/Ef4
bhKbDSzwPdcqtaABj1bExxt020e6zpL82WaafpIpBmsnGaCIFV+T/Lgiqe3dtzyu
BNyitVcq5mANJdY35xoJjHIe+h8NvXqw0Qy1erlGcv/MKiBzEy+V4LZUr29VhnJY
wBazagJs8K84zgD8u5ZU7APlIfbbDYboLDXPHp0K6lc9Q0BtsO+FNLzCwm0viRcN
sWfi1p87zm7DPpDkqHJNX3GALBmViW8vgGPAAqqbKVFGMX+TS+Je/jiuIPndCWBI
lxkNDOHYjeFmcXcbO5LLIHk8xjLiRQ2svrlXTQKgQkMqT0rIVtjlX/wzsgw7aaQt
VTisGDT7LvtCk+wJbCcwbmNZNchyzWfX8JrB/KJZ8uZJkOGmsKiM7BrIoWYH8M6u
we+/mbU4bg3oIl2+IMPRvknE6ofNwnRuk9TdigItGpRHrlSL26uhv/uY5hTGckrQ
JUJMEFIUDgUSu0W/6Oo+lA8Tx/XzM/ti5IYEcaZVD/KWqvLTyy8AEx1tOofaP5TN
dlxZGz4KW4jJ6iwSHL32c0OnrAdn9Fopv6XE6NszANWZB5mDB2a2clDdAmkNbl6+
HedKCbAFDURLLD3xhO7w1aSMgo5/IlVd+lfFaIvSYqTqPmir7/XxVT5Ty9Ix26ou
JDeBe2PSpCuHLwX0HUP22l4xUJrfERnTKOVSn3/mb6K7JdoYxsHXIuseVcQeGCst
cmiEVoDSbvLs4r8jD6Q9KtJNOtQZsKIOKgvHwe1b/Siuy3upa6det4BUv7M0xj5/
q5RpbJliagvSlj4cPQcErg4/7rR+12IgjX1b8V5TbJJ9b2wLHfWZjdhXshY2UIdZ
CvKBmUv2OCKKhZ4nOM/MuZacTCScybLr74W9kj15M2Ii5XQ9AJpySxXOdkRV9VaD
NMkubCIiF6DTzOEVKQ3UzFYifZzewXGhp4hMl45payquD3AYclPhDzP+/nofklMt
/XVnk5b6qdvuFyXUEREqPuUlCC4goVDgIkQFvqEJxl/OCnKn7M1J/s50vtHpunM1
YD9p5cWdxbFUwllrWd3Wh9MJ+Fs7sJ224CPeVjBf6M5oTqK4KZBO5BRzVQImE0s4
ZL9aNJAR0MhmFpA5tsidZIcGMWRnhayPLFIwfulkN5706xstuw0N4h118Ym4ZxIS
PjYDYQChdZeQKF33zFZa0pIXwnFj6xwzv7u1O1coA/3iUrm6LIbWuiqAQrUqoYCO
2b5PCxzARokoYvPxGGm48H/bxJqV1HZKE3BwseyhS759qHo+2Pnl43xjg8GaHwuc
Zsg4D8PNplH6M6gioNvY9IcBTzxQ36qpUkVDjb0Nz5wY53z3o1xIaveNWKjJUl9R
yYrqUokA6/WNpb57xQr6mmZC2uWBKL9hDunSgO1ufc4C7S4pf35z2/oK2aMhzSnI
RC7WkBUwxTK7hkB3/ZS50n7+W+1ccUFhb+7lYYmA9+lT4cRxjFS3+gqtz33G5jy3
wlanSVPYZ2zQHVaRwQK4M5O67JpJWMIhMgqPxw8MQiGGEa53T/WTsOmzIpogGi1/
Dwa02sj0BK7Zr6VvA0DTbiQ4IxW54DGDfUUj97eM1F+yloM8usU+YH49EU78qngu
EorJklnsDMwcY+yxf6kMPisfr+c9GTxxr4w/G2Uo8HaEP3FdulFHmSF+7nDIDFTf
lghBVbb6PeWXgdAQrbf4T713vWb2JSJKng7tg1x5QYHTXEH6u/YyLdtNzp5XeEsH
tWOyeqCFFyaJckG03YcNJEQhRQMxbtn8d6KfT1sYGa5wPdd/FUtK/DKgXaD9Qf6U
0dkfALB79ZoqFYSKCAj+cKF2fJcwa4J7FODJF/4JMrffifxDiGbRlIX7W4siB4wi
rJmPswMeaXBr8Ni1g631wmaB9E5eQzuZUbzFjrr+ombUReCNPViKXjQIs/YnUSOp
Zj07xexiaD/KP2nvOG9HYopZ9jliLu4gOeNHXOnBXNeIVKHRwVrFc5WWiq8fgtzp
ys1s4ASE/M9ReIR6dtmPBkbAaY8AbuSp73kXGmVmJw3w+QzVlXNgs743cSLNnlrb
k2PhiO4ayErQWq0z4xet5RIPv5pQwvt+ZPM9XxfesHZKn8TJclUJsuH2A+VX4eFz
XexVppnLhN7m/lWPVRLUMGWeyfOSeQnPmT4vcIRmKkHoptE5PMvsweT3W7H7NDR+
T5+o5g6wZGGaQlO45drsgBPcAlVzxJ3TcQonJcvYHGs+9Nhc4YHC9VSKjvGMo9F0
/hhwpMtPsf1B9fIr6Iwk3zjICAYWTIxxjRRlWOEIUVPZnReR+y3wSt7PbnCA7yr1
gpaDKkjMWJlx+ma9bxdJwujRFXmOPrUBLVCaRrTFDGmOGXxUx2ygMzbT52A3Dvr6
fJ7oLTfNOid5T5n/VJCJDEzaTL4yo8Y807pN2IJMpKyn6+lrq9AoTa+KTVq8RGom
GSscGLIlGtRPhmmeq6kpgpvtT8WHNmfPa7TR06Dxmg5t6WQ/zrsQHzCf4VmyX97S
stjgf8TgcXbi56gg4i2KgjlR5/1p+sIoaMvIBV2J8w9XIXxgw/STPkaYGs6OcwWq
BKh00QMxaOHsPij5P9gRQPcFI6CyiJTnRIF8G25TIlu7PBpGRYxAzKWleEOhGZfU
+YdZ8vxzmZh5zN3JA+VCL1dsgxwJu3nFhRXdGy2NYiM4xAHlKukczh2O+WKuadpo
qBLxNt07snBBjyMo2Nw+qNnPZmdrWJ+99XLyr2aO7QWHkERrTVxuXwUlxozxwmC/
JGVVgfpjLrSxZHrw4QA5SRJ/S082pgZ+U7RicN0QIa8REHbC2EG5zAD5IL3H/93P
vHge+rBTPlRZe+5Gj30J1WYsg9Q2AFImxIMpdFyVtTRO0qzYLuVJfkrZw1HX9q/o
whMSEhVH/vILPk13jRG89nYH3zG26371st0Uf4Fd9H/CJPuPFfTahFaiRmMWda5q
j5c/vCsAAzTQ8Jd4Ercu2RdUIEUnFVHN6F9zQuXi5pYIlf5V6ks8V4Ys0me4hOfE
soaXBboPc4a36pl53WHg/JT5aPpQOkBKJze8H02/RY58769TIQDVsoA4kggbyKYJ
Vj9zh1JncMH+DMCiAKTFlEhw7KAQN19of/5zJvPU+zyGZpom/6zaGx3LbjqUZSi0
SuN3fbLLIUZMzHVUuwpIjpKmP4jjo73aWkGhF+OPIFoKDqMEh3IT8TZ2r+R5e5BX
VRihm3hzI8TI7kbXFozzDqvaJHGHvjIPbKCis+M1u8qC3clDOJa5o70folFmmRzw
mZOws+YUsMJEuEIoIlJTXzlfGy2ipQPHlN+58JMpN1icKNYxFzzzs46DMJUD0Xxv
ahRGN986euLgop7cRXg1AQwrqUJhbbD/KfewQnIt8nG5TwE5fpFFRENCH0+5xr/p
YqewAdcPQT7hBsVa5eGQvRPMuOuqmLLAH48HVd2tnwtQPDuDigloLsom97ODZjcp
93r1mWJ8Wbd6K+JGtSb0nw9hKuXSI54F/Cj/oQb7LE/AKNFN+pjPExG7OrJHZwUm
nlg0ge1iMyOuvVYiacWcrOL8FbeOQcdMb7jHTjA1b12TEAviVjPuiHuFl7L9SPCy
6vhaojs8xEnjRg1b/H8wVZwZaCIQSrmGNdE9DFFq80NiHrGLQONK8LW7LKJNtiKy
/BUqal5sOR7xkqek5cwe+HEvYvxqjZVDINqt9n2oYe1IQdtCHkZMvUvP5+kDkZPQ
hyKqdpF/PG6Yg2KQAJNqTlxAGQu6/gnQQJrEpFl8pj43ofP+tkZSWSp+08EdXlbH
pAH3U8ZhB+eTr9Dqem8bvCoTGzvTPfwJ+iTdPP1DvusY8a9LmwjzV9JwyRKeUvu5
MHJcED4PTiTiDpgq0BTOG0Ifm+MWjaAfnE4/KpwEryaiezykfhWoDbPD2CxNq2Rp
vusaL5ZzWwwUcB62rG53GcNInii8fSjL5XRWQs+cKjyNZW/90pcT+k6iYykpNeb0
MwsVF0sGBLjd7z1UE7sW2CmqE2JkDq/fdbl9g6eHRww3kn5d/ck0yyDZEXX8YAOd
B5MCH+buxjCqaCdh1OlZ+eeEP+aStvtQuZEyvYY8fyv2ysoNkuogqinepRt+RFaT
l+VaSngfCj7KwHEUGxHpDAVvzC8VZHbUODwWoq782GNEYTaOuOcNjbnraGnASMze
xO473RKVJLpG6RhgmmEuN2H0qpADKeERH2c0hgaKZSikfBpv6N4xKQAuOped0BvM
f0Ap5DdbMlvDLYf3m67zoNoejppffMxbd4JuSalte5fgGtImT0NTlZIZwkEf3P9+
npu3Wz4Lf8Ab5aqE6NJhI/3L/2v3vuFPYRtSbBtKg0ZAT/JVm5DClyprghmQUvYy
ND5qi0Da6A7kORadrTmdFyqlXvmcp0AsdOwqHas+OY2Xoy9Tzc+GNMYC6CfDs+13
hOo9TnvxPV0nKWcAFKMK3eqpaCzqP8LFRZYvw98fA7YHm8Ze2Wo5T8gLJrWvvyTQ
mpeYgyJOI+f1beRgwP7Jo2I7QR84w6W8+o4SeyUeyvQP8GkgP/DEab+kAiSw7n/e
8W37GA73rS+H08ICtdGXIwjzzxGvknTOpF2GSFQH1+WxIoJk9DIUzt4GisWgGxgI
EI2k1TjH5zvDapGQvNzkSa0L+oUKvopX7SCFWUZwpBlqmrGHCpwrEXkAP3U1YwrL
X5ho7c5X7OB8Jw9eG2gS0ETZBxAzQul8RUMvm2ymx9IXAF8Emn1AwwTgjd/UyLcv
YJLPHOi4UY7T+l48fbXDWMIzEZNoBDE+i7Q5vqPgfUZ06nNVrTmjYwCdTRxD2Heb
Q67JzGYZPkf6EKxk12fVHWVPMup2O/vjXqtVdcZcYln061ha02D5jKLU6RuN13yO
4GBU2Qs2legKmG8eoIL8IzPYcNWf3jqNvrwVFuaVCOtx+ec6ODy/Q69StUHp7lko
QybfKYLRHeiN8Mhk5fbwvkQ+26wxEn+Bx7lzn85MhHD+/NcPWmPvGvpv88DuJnCu
mQKFhEWJOhmFsgZWzUUyUippoVPtI68fiEeq2JZxqvfT/TrYD6Rc49xiu52t5586
bq+5eYOOhi6/kTlvndJO6NPaLsc09Cq8etgi7EZlARo+Erw3zYdbrlu2DxI4XMTX
Qw6QIetMvF3TqbSYQi5caYHUy4jm7iuzQuPEWpMuH/0qDHwiJ5Mhn7OQvOvY9Mn/
bUKjk1MZecUHPcL0ZMEljLWu8XR6F/0Sw+Yhc1ukikPvo/GJJXXHsjKod27W1/zg
dYoY7Bd2rjJpgBIxpdjpQbBttN7lUYRYDV9FIS2rSw7zNWodCQy0/KnJIN9cWn0V
BwWKfwt0VY0mnKkxeHoOw5K9h1TZFXtUSmAc4Yb91rXEBeLEiM6m+M1VXxMvVjjF
1Vbi5rPqxPX1SAd9Jz1C1X1o5bKNj85eKzQd85RWngBAHixotnFkIt6Z5ZbKVTxU
UH1YdZMe+VgMGBip1HfPUqjZ8IcyySW0tHQRGer8GQn+fvuyL0dKK/OtQUjE+LRN
PCWGRaJHUk020ylSUVlkbwrJ9BRc7hvUVwND+ng3hCq6J7GnVkh42itCjS8CRGxf
Utha3ZU3wy90D4j7+zB20fL4oVfSNZzPQU+ws8SVxj2gwwQEr4QsIqVyrethPxbU
aqg50cTHRdtRh8Gx1R8aDTcTVJoSy9xI7rqM48wiYapiE86fyPa+f6OYiGl3V/im
FRKzdtI7FFGoFcReNiKbtp4rihvE6SNxjrTvMkSS438fgN3weotf29dbGZm8a5ow
D6SAzPQ1dS9SbG8ZICcXeuuvoOwHYQALkDygBHkx2DVmDb5tGBY9NCJJhczUl+WO
2B0nvCBcaFta8vJggeilo9I+AWdEREpXeaOdUTPuWJuVd/KGX98VD6riQR4a9/7q
e8R988es6Y+n4lqDU3Hw86V4n3XiO6+HSGsU+HjSCxhd0yLrnSoorqDUe7UrYqtd
t/yLD5qKbscB7YrHVuxHQXSBsRN+QQ/7Vtj60yWiK9yEWp5dyjx4js+d3Qw4utLK
Y9D5jPyxxlL6CLYX2vjOGyaEnGimt0Id1d+v8XPbvwE/RtSIsGjLKHCIPUMDhHUl
z5vAPrGqdNDxMcLk8Wd3x3JPwOuKLDuJXmmx0cpzRhfhflvBjGiFljKSYKgey+ht
uewrZR2JWOc/d6OOICzORaWgH+jFZw8MaOnTY15rXPv61E8RkKm7vEr3iHMbK03n
vjfYWyf+OUNlPezCnSmTtToEOZVQWlbvAKF8cczwWPCQPJpYrvy2fRPADwqxKwWX
W+xgFNB9rXpRUM22jjECFfRlTllDlpLvmLhy5BFzcXsWoBbwhMOQQwly0n83RD00
diz/qgdIllDh+/bZzj2tRNa+5mPSCOya+UbZAZ5+BgNiVbQAZIKF0NdabkR6l5NV
RBBFqmBZXCEIjmfygwUjIssp/RjRFeU9LdAQyyrV1EpzZmOaghNh0jELmQ2LNV1N
zsOLoCX0RaNXj9VztZIFLZ/WV+FCsYcfrl5MPdSCFJWzRI7P9vEs1ors86Aq7eXh
7odpIMFpFAN/39d4kUkxtLFroAQLKymjE25pqnFTRFlcWLrrpXcvc57YnVcon3lv
zg32gQiAnrjxRyMxwqTWJIMY04+JkHj9HOLyJUNlB1RjVtNqEzbt733jg5hznV2n
hF4bwc98qRjfq5tKvF+jtVaSl+T7aUwGa888T78aNYium1Jzn21lX9Sfe3/iUYyV
VzhFrpR25NqHXwyPgiZ0gey9jTNFf6656Tqd+3W0B0B3xO4nJVimFgjpvFsuXrMU
tRrQ2jheIubjyuXYMk500h3hSIwO1UdP+c8QXinX9N8fzAL2PmgnKabSrR0dR73R
Et9xZA0Pzg7+056Tu5mGwVx2mDMjiOUncgBayXVyyr8DH8jI9sSqxeERuYKezfaL
RIUuHT6skL5JzSWSlJei9OrggOKBUGVXvgK5VgmhEZShjZOhOZyezKtZfZHzDMWU
0+X5tfr5sw8LhwEJiMoLyajDYkmd067RXCkoYFU6bzPI9Pe74Whhumdv5P/lnIhO
p4Tlr9a2LzfVEfDBXHGooF3HlqbRnmVDmwC1RYfQO0ZgnRKn7kW5lSpUsDhlAS+S
sEKiPZj3JpFoyLAJBhzpMILCpxXuh2sUlHt8+I0498k7Z1gldsIdn90sT3cd0MC5
9xRAxcqPLWcXT/3wGDkHo6mTO3s4HCdb0ZHOdBvPoKPNS+gpqqqJOtXxGjFcoMRg
Ell3vSOjjIN9303HihnpK6ySHZlm/h+vBoQsamDqLSQ0kJu07+sXv1cvg9AoW6jh
vukmuxWOKNajKR7PvKK8oppf35nGzKpIC0CJCwCiN8bGm9iMJu/rJtlYDeU1Qjn9
/yexk6xMl/AWu5/FiMZcoxDJy0Y3UyZuY73B5BvDQBHVROLO+26Q1IdTyQaq1N1+
Bq2/5T5/5DyRafcVzRW4edf3uYyKVXFauNV9Jedf/MxMVkbFHPB3hW/DFy5WwQ03
a4fjhlpKTu9ZFVd62kqw2EkujmeBPOmxmam71jwgVz4XwprxOwIHKgwu9pSupanw
xxRdr5Ha0J9C3zTWbI7T4zU5/a9BfmF1NO/xuK7MrSzZI4NrBTumFiBfrFtUrw57
JTIyYudBFbRqvx6cdBShzIe3cPUcKi731e7USEQeUYZpktMX8cd/bF5itrtvWjwh
mXGeQzrhy2RU/L/r9dGzklhSUXWTfNs9J1KhKEKupJ0m7nasCvQjf40davo1uWxF
c0UEEL7HFk4kkh0LiLFDwR90A07550cciOQog+ccHmccytlSkLqlYg7lcvjjtHJO
8w2hSiz6l5+pCSYUdbxvHgNCjsg91ZG1znba25e6xU3yKmInFR2juvsTC6UTzxWO
ZQP48aiBZuQXGyWn2LTFX8mxx5hW1dWESa1UcgTP1xgC9GXQNM2pUexZquuBcyW+
RxxVVKoMl/SYPnYLi1vl8/Bj8y2Y7bxUSgdfCJTANLDNOi3PEnqKPwuY4LayZZI4
oii4P8RFlNcPeR3A/a39spdsQcBKGts+Z1JT4DctYVoubS0tLT/LzOE35cDpBTcH
Nygkw/mljDB60K39RkwYJIh2b8VA1sQvjLholQKxuQzzjwv5MXB5ArjhUJaVPqnr
WCdUuLlETUO5cho7+q38vrUS6p9XHsmhRJTpZNGSlKK6a2GqJ4mUqKasY2v71kha
BCbLSpxcctvLBxhEaIQ5GtYZJIxjJjGssfWlc/xX5rtzw+63NlTZMv5fs1x8GmuQ
tGAgu5FnUy9D8WmDZ/jzpcueKYXERBseRh8UKz0me5m7bUVIb+80fW0vIkMOah+x
LhMyQwLNhfEsClutwsNySdv1ibb7rujk0Cqc4KSTVN6yCAaDWWt2r0YlWe+V/c7Q
WoeQwayHEEOKMzOKHuX461Y3Sy2ye5Pdh9SuYiL/0L8XtGPOFSzrCPaeSapOeJ1Z
7ktZYN9PJaGTrjclqVFVZxDFs2SVPJNrWTmCwYvMKlOpCY6PAfTvFO+cx7WF9jpD
lXE/rtx1v6iuQ00fuAIYvINjGc6c+OTSffr/Ah5J4pNBuyOk6tTwzlaXTckmPBDq
TpV7ksS4t5ePCqCa4Qz9OGVaNO5Kg++R955oWdhRgvxelOk/VRkxFNEGpNCcOV/l
VSPxfrfYSAMEE4yBBfnazKyMuY/eN+elAhXneGL2tOdCu7GsMOKmS5faMkGlGMUR
qIc0+bJVqw3MoRFsoCls25kfh3Wje2tZr4A/Xyu0uuOb+u5KzNHzNtS2WJfgu6Sv
pf6VhUjwb5JE4va/6Eem9+DHekvDktYeTfQZjLlB8iaeUxbVuDt2bl4uIwRg92xe
lLkwkbbxXNX87hz5dBQh6PErTo6KWHwan37NNmsPshPyxUn0uSHd8OB/yI1jCshx
UtA461heFkInV78H3aCF629rxKx0rDT801whpgEWqtOSzRHdNUI3F9NkGAIKJuG5
anamhOHhlMXVvGcC8+zfROj91Xl4ecjzv6TXTYCz1xoTvKTXUFfKMbXFfNpFLs2O
Ow0gDwovxskXzFoTbVE6+eZSU8TRyLID/i3znRVM+UIHKVVqjO/BmlscrC4y59V8
MGy/MsmCDH7PfdOvbQ33SK5iQ/8UIfMwLP5dNt9Ziuq1mSWDKe0NzRuroAnI5uUc
L3bR/sUfYcqcukqWb1mza5avpDwhcdEwxuE5TeVX3kdy2MXaFuGupEtoqNAO/T+R
cbOtqy0XNpLCT2ysCPN6GHl5DLQ2yonKdTcNteOS8hlBHHPd+QNrbhTcNdK+Egv+
F+4MR+93n6AzVPy30dUJL67G6oIo3SbECbGzxs3P9XTnBmll+yI/pKitqBAefHpa
PE9Sc/GZE1Be9Wkw5N6dJ2/rIlI5ZoeeHL8qvAzimyoyr1yPhNrn6W8ZNH5sTklc
W+Hl+7ltqb8qxpfAOIaLYkYJJuCaY4YjcU35fkXiZSWx8Y3ETNKEAfzb84VhzGla
6Q9vNL9LkkSLkiu0pqgmlEBY1FP+yn23P6OTBIgFP/ZaTTtjub6bLuLAQt4XUoqP
7Z+uvhalkZx3r/LJCWeQiC/BqqMyTY9MCPYb+WqcgGSikI0eKTvePcMx/ILlFKjl
X5Ndasrw602KRxR9/AhZ029BbmhqxwmueB+AsI2rl2oze5OmrcCwHYsZL3FWbycg
a2K3TKnxsR99ygXQNN+mSGvZF0kGIhmMuOIWDak77LSssVqnAgSzxD8sbDT0eStt
Tf54QO2j4e6hHzSUhA6/pGt9i+SASLTufQdvi994OW+7vfSndp4r44UeQhoSz/HH
brLffVzps81N7OCr4JPyxcm26E3Tl9bhlmbU7+nElU1YORwVwtJ3twBQl2Vt5CWy
SWDgJC2+nUCjF/xDXIZj85KXAXeCk/Q5j+jET8ANgnSePFFZFrSQkyjRTWIVOT8q
oGMxKpMLPNzDQTHxVfhgbanEh+gwidcf9TXMKm7CItbthvDmnXEUoC2QCFXCx8p9
HUL4m8h6Z5Ggrk48Z5M55zPM98OOlkC4dYM+cElCb9bNEMyj1o757RABtOupgPFX
qhd8AAB4uQcrUufGo2dTSZISoIpFyWB+iK9fKqisHO+IXQlXAid5BmR3Yj5m3hIO
ZXUkKaRPlYLjFh1Nxur6Z0e3xIaCIpzyoH0h6gyMJ8Lf34ZkxJJmnbdlAzYc1+uf
y/xtGSy/vXqxAGdz+hdpwr8yuZkLq5fUGS1B1bOZT9q5VUsmb64X55dWCYU00hnE
BsrV1IxkVJm6iT5CTyMOyh3mleToU/63SGDXUap6NhCX6fP6kudXRb/ZBWrv8cCq
s/ml+Fj5J9X1/6ezPyHrOplYJ6EKWkr5XMK9wNMclv6IwEkAwBQg+xFY/3+gIOhV
kSR8FzzFBY30Ovb6mY6IMMFNOUNvPSKInxiIKqYvBAqtQzLGGRhR2hnOMP8dEZVi
HQroRF1TAvDXoepDYBqL1iyBMfhiYt6+NwX7OZys+H5kV43YVuqWKBJSvnUHhdxZ
iBOiY6QbE9aHbRBG0qxyPl234iLULc8J2vY8QnOnwJn5n4E/BnTsKRBzk97kMceU
7dzpGvaCdV5E3mdkN8nqYyEuzqq/+vLq3++vknmeJlOH2/cdpUUb2G598mp1W9f3
U8M+1GqRtOsM7KXYBFMVoTo69ugpxipBTmNtIZc6RbfUJAr02wHf6F4/gTWkpday
NMaP1NjEEVHhd7HTk9U1u+7joWvNvbmU7JOXCYr8TzoL6/apB2lAE1GFSNceKAbu
1mfh2d9R1+75SAmjLySwmHSXC44U4+VScHWkglAp92t2catMcEc16Zm9x4lom58A
uqHGBAkYHLREHHcds/pTSz5yA559vfAK3woNKsUJjNvXClv4VvQUkdtQTqwrCbYd
jiqCmswDV1fPbH+k5TBvwZn7N9xHcfSQOEj3ujMZg1C4CG2a0R9nh8cAcQO2P79Z
peQry2fssh/X0cyQbdHz7O18Qz5vcsni1By0XG6b96FQUcdacLHJkuwaXrHRR5Zl
M+sthj7/NmPFadyJfSxCBBWmrISO0wRhlNa4+RArDJbq6nJpWvYdqUiIGEY/W0fS
YLDkn4TEJR2ZUc8yAPRKtAOSt6v/72P3Kf786xr//adceXa57ZgoXrHtC9c8vZ4x
ibFDIPjo+z9OtoTvWvZJY0y0echacTUizWoBjpJwmxjt43aLsXm6k9twzJegWYp3
voKaPC4yetp2GkduzQEUjoqGM73v96j1VU+OcZWe3e3tJmP8nqcqKhWsHDwPs887
STH8JnOWqQVQ1TRgn3mSJzKUWUivEYqc+gvqzxXC9bDtabdS9fdOcr+NS5bSq8pI
pFMG2iicEiAKaTpZ/wUrnpOy/WE5FZBxivn7v7D4LRW93ObAJQOVmDM52FEWYS4b
BzgpLITVn80b0GMIfwRXw6Vpr3O6zSSXIayMwg6w24GF8T1q93f3AC7q4hQfmiBo
f9RJchdhWbsQBaWSH09uonV+IiIVlMaga9Ji+EmnqWL95oXORK05ANugnX43qeI1
nMEd9P4JxP9DvVi4QlazcKI/09EJhIi6XaIDtekoJeZ/NwHwUIAh9sgKNsr0MpIB
jeC2J3Xsqr/iR2TgxxL2t2kt0KE8kxLBNcrit5BY2J31giuyLLXrYMapn4NcIbU+
R9rf+UoA/W24R8foLPbEvFBedG0O3vtLmV9g6yuaopTyqYsecqW5EOR0savGLYrn
loTs/5mQbjLFXZM8IrC0oCwaqmKdfTXctog/tnHcp7mXkbLCeIKlaAEIoqIs/Cs8
6ESvJ+WM/LoXGm9pUrHcPGTfLx7nh9PLbPa8bcLlPzaVn87R5DTLr6f+5pWt/lnz
AtzBwrjq6OYb5XNXeg2itaXQ6L/cuXRQZ6YmBXuMk27KkT3qf92Lf2QNynFDnKMX
9hCdOp5pQaCO34acE79CLQjF9hX0p2rNflUenm29LbDJJL/Vbjqa2AybcVPaXBb8
S6jsdOiDcgX3zAi2vjuawGMjWFyuvevHwV/Kmqlndc5fJdcR9RMIgOZHCpsoASvL
Q86r4H44sfPiHe/InrX+Z0PGmgO5Kqcw6AGzLhRYZwUUgBF1bSCdR89IHU4vdsd8
1gPHQ76u6Bhz4bj9tq4z081sezhyKuqRfL/m1RXHZYCwaJYzn/PUri/BXUG3+5f0
EE4Wl6SQzNkAGAhFuRUZdrjBY+KHTBy0pqB+WSWHlmxpcI4fDnoDE5pv2+W5EZTP
C68j6gKxz0ZKRW0LGVs8J7BfSLBo7K7pOHwveMYI9p0+8qf7VhE6bBbYBUYy9Kjl
Z4QQJjzVyJqhCut7JqqtXuZtYrq985PR0CGVlnvjjp/1AfFD+WqChIZXCmL3U5DM
ZUL/lrqc1AR44esCvM97CLBDSQ0VGJv2/PQxZkCu01HuSzokTlahAIR4EiYSk91Z
PsFYiOFcTIU6AOZE7qip2cx6ar4x1g5p+BkHhdaQGf4ebSEvUgbgp9/TvJg/6WkA
59+io6F0ObBUheL18KI4E1tWFGbOG9lJsJuXJ4qX6zbMM1r1jHlr6raRPbgJADsG
mkLDbB0dQMbZkj9YpQG3YtW8L2ShQR/N9oNUOK3t4LWLxR/EIMmXc8u5iNi45jga
OgFQ4gCxx9dIMt8EIDMDf60AVlNs83vGvnIVs07yNSbAzai5W1DeSKCZR1NXXl81
WHv31ghYPmFLL5onreKhurdVJLKqkmZpwxLzP6VpP/Bh6CkCYEG1/5RO8n1JSPfW
jLV70hAZp9ucBvF2thhZ91tio9OwbFmLrzw4goHu933jFbdQv2de5oLs51XqwuW6
YOAdEY1dq5X85Qmz0j5KClVtPw0SkAXXUAb3xiBPZaIPpUiYBA88Iwuuog1J6uUW
ftH7eKUMXLNJBv9xR0MstvoOqb8jp6n6awBP5NY2fbujbRytJ4UDfuCRc2i4A0gk
SMKB2AfKedMp6qW5RDD/gimHbV38HPSNC6Xh/+HMgRtLCAnA/oXZQ8/C19Uquzcq
IRHAorNr1gCArOXktH58xV67eNThgpuxmyOtVDtLFgFd/d0dLsVy/176w8kxBIR3
0Uiu2uWrjPXUun4KmbECm7zMDzzGN3+z9eNrCbO9ckfdNNdCff+laIdze7d3uB5O
AlYSNvCfo/a186sgWU44VHsv1OkDDi2vtrZDVv9gpNiYm9t8bSCgLHWN1DBiZ7xb
uM+R8gaU1JJ9c9qFcO2tDsqSmshv4hHIHQ6Re0SVNBR+epCSMBcL2AjbUQWj73mj
oUMNo639DBxCuZexrTdftLglsOn37OGVC+rrJtNb4J5qw4ie18pgIA+VJ8MzM7O8
91KGXFdjhy6xWeFVsVPZDRyoUyG6XXH+MweQwulCyoILuNh1Hn6Q3b8PrRtLr60L
FMltRg5FEB03veYyo5M/weFqk6bg7sc/O7paBZbHW4tzJYvA0g1G0a65yV82/5nb
A73s77Ln1XXiPblthPsivmUt5Ut6loa0k6XKEDbaSkGKvXzkg5aDdqu+9pRgMgli
Q/OgoR5ZpMMS5rJb3FhVMTp7ySI4L8LdOc2vbgzUedcMi8/AwZ8uo4AFk3LZBAQh
NWQr1XDXn6AquOytZs8MDgzZfMNyCIBv2W9il8t8GxT+MmE9LMtqwzTXVzH+4ki0
ed1kOlGXN3sbW6tfAO8lKZ2r5rQdwVTelJB88acRymGDMed9x5GV/jQgT/UHaz1B
XhNSdGVFBivtkFk86OKGk0DzYBHwFDGjYXGB6vyLkF7Jm9UpzG3sMA1lajPCUSmm
Zicv7b5d4ZQIpSGk/iSggRZgI2AEnttjQUTiMqZlQOKV7lDx8y5Vk+MQe5ujDO4/
paiDB7V7IyztUKvaG7GUwDzVEMhbbpuja53cYiPwlHm0L1UVUNKbBPN5UF37Ku2m
ONLL0Ma5VN0HGSJlDadIiQiacYKgVgPK6os+wyxN2ouwMQAUq2qwOJW++e3b8Vje
0PGCTk3xPrRaMYhKNPcNxDVvJQCcry0HDV4pHDQylm1pApE8es/rIb/5W2e7hDpP
hQUn86bIkDhGRIU3c6cnyXWb6YmjdEXMA9N/mOu4F0bS8jmetNEnjJ/LqJ+yRr2e
2tejxAYkBXzVnfShE8dYFsJRevLahG1ppow8xDFCkE1ScNfYq/Pcff2ug6fgd2BO
X3LUY7KH5W2GqahysddKnmWMUtWJXyBf2rXnVX8QI7OxxzuWDdQ2bzReXWTQllLv
tMFlYKgPf6r/qU3X3CgynEUceoT8+tEfoSmNlN+wSTaJIHR6C9I0+1mmU9BJbWzX
2UxxgcBb6KoKoZaPAEQiGEtX05ZcLie8nKq5JauDT5M6xSxoJnqoPCRH9qsGStHP
gkDfFiFaa9QpEfZRxVe6Jlb8HQ2B/m7RDWiFJjujfP2WMXA17fb2kWclupchF3r0
K8dSCetT1UlC5u9AGmZZ2I8AKX/MHzAJAwiQD0b7c524oNE4ukvWfY/DpQDkZz7V
TsnK6DRYFv6nky/HaLEriPyNRPconFZXKrFxh8Lj1rVSwANV+STl7F0e3yMlOCi9
LFSUH6Bv1BTjmRM5bVYZraFdi5RvoU6Tv/KEpnOKWA9dRpFLgPKCsJgmC9WYthr7
0ItN4566BYVgz9evEQsGdkkSFzJ3mniTRWvC3g1wLMag1KXN/+sKgC77vTPTkABf
xqlWFLON3dV3kFzW7pdcUybFxGyE1oGYFfPH1ZF4k+YbBsFwNUEWk/ZW0lFHqDmN
QwONj9C4zDP17aviQGa/EMt0olZ+tAD5MWU1pGyv4pioX1U1l4MUimoHPy+u0s0+
ue8yW3g7xwBD5EEVQupsEJaPY3yvhZn9nsAj1gLa/qHS22F2WtBSGypFaP4Dztmp
fgwcId/wNVPN8o1Iv1btJJxIEnwhj0EOsm2xCR1mkMSB19L5DMIrReOlr0IIPf4O
zT7fKReL3T6spMEE+5YTpLu/nfuDFB+5gtS21tYDGdf76688k7nO3PN/5DBw+8O4
z1xhjcrYoy5kJoxOx6Y3FDNlc8+dpOQEf1ep4dEUxdhGZvOMf2rYTUcmFT9EBat7
5459AFk2/mSD/RvTtviTZ1F9A3kBLd0eU/i4ci3szdUXxhvvSQkkFD9R6mUBkuqG
aLbO6tUjIRo1GrLEN/0A5yTP6fDjJDijsy8MrwWUpspfVfSYxlSf4eOIEsDah8IS
edKmOwp/QHriTzErD8wEEYKJUIAaxViOiMGXg0eB3xCCDI1nsurXcVYlTfn9cu+0
ftwnPV2K2Rvxqcuga/f7U66nVsvk30zS9wrFfofNtkUybbzHkzPLGKvvc6jIVCQx
7UjxcbdogRl3F9r9KbtIWudvxzTk0vs31IMCzu0YYTIVyXLNhQJzKzUz6Rl9Of+e
9w6lTz70rh6BXAZm//kZK7x8DbOfmtoUvrTfWAfL9XlWI6O2ZThQ+ntCmw6TZbzN
LzBirRkRLNl6OwwAfIiBVni4rK3bTvm1yPYhqbIm5zs5gocJE1u195lZ2Ix6Boyn
S9zRw7x/3+bbmBltOVZGL/LkWcL2N00jvBP3RAB/RYc/YRwJnAjWjFR2dSB+OcpJ
RLcCmbIMkA3oHLjmQkeIfgy2225U4MHfF19rfrMqbjisc0siNyfwmnet0g4mt6l6
3p005SsZKge37coHgyyqoXnnFYN4PWsOqQiiJJIsyTzGghtVbk+5T0dN2n8kev4B
a1/+dIrlQ19eoxOZYVoeBcHyS6qySM0A7jh1cetTfTWnixETAyArUw1xootfdlpC
Sq2gjUk7WRJ2bi0u6vfAybUhJsKsJLIcsh9tqz/b24hIyNpJP45k2bdmWIS3a4LK
lzNhjZ9sZj4jqPk8FTw7F/L5Ik1f+0HGzQ5yGmxlSFThaQHEVt/DmkfXhNUevDww
Uvkd/D/jXPZ2rqrarj+yMyK6G17obyktYlcz7d2yWHHS8rw7ju83uEMTdEn+3fmf
QM9A5gEEQro7COO0cc+l+E5QLMy5yLiZzjyVgm6T3CjzGSaMcAQN+WY48SpruH6N
BnXGznmHuNkDFccjoK160o2TkX+wBruiFb9MJsxuUj9jvmTsUkmcGPOLW0iwg/R2
SZ5TpZrR/20kHGAamJWzQQurj8ZXVSjej9qFplCuvnXYdzxjtupR3yHKAeIGhLHJ
+Lu/ZXaXqMHsK24qwz5Vxa/YylYFfMVa+5/tr0aNFEfRKk1kK4rpNDgp2Jh5N72R
Rz8foQeTOUcwFLEQnesy2tZgdFAT1CIXlpBsiWlgvCH5VJxBwh7bXzb/F5mIlRvi
5KjSiw2jxQ1mo2ZHQjZWlVlAuKtBjR+Dd4SyIdDov2fT0xphJDx+6Hc5qf4GpJwu
X8/JhdADH8mnmiiURfTYkKBSAjkWBbduaI7xQ966U284hPQsEzx3GGEpZjTxdhl5
T/YWjWQkE4c0S2JL6/N72IWXe9LDXQCmXVNvQhaGrzsbOqfA4zWF/0PboGUuUdsG
3TpJR3IRLQhbL6R5TKg1m5SzAVWYR7n1St4I9ODgtE5uUv8lRO9KgHIntn9tzDnW
d0FjttRB+xBKRaC0kCiQ/DNA0wP1RnhiadScPVD09l+oaIj8X4zC2cUHjj/6GaGl
u4lAKDVQ+hXG3XV/CFxajgjWpw9AqUVhgK4imT0kvFUTWzFojND16at6QmlQRIhB
H7q7P7ztdQQQNW74ZWlsYPGnnYIoZyvGgRWAg26BhCzX0H+8soiqb6G8OW+7AXp5
G/tEJDAwzOCIbmkUb836HBXqIdMjg861irrplsEQBmonlGTEDSzqG3q5C4RRAbsp
EorP+9Fi3sj1w+rOdF0NeW3jpIJ1p3w9xrSxORyounf6WRKXr05HuUnbG6KfwZf6
JOj1Ja/czWVyelRLqXbCPgBj6z7C/E1jBCCI47Xe3Gk4rHBq7qTPfHZq2sDPjWru
dsfUNgnl6X4Y4CND1RkdeSwQcjllty7Lw1hqx3q0mKdyoIZxsmiI6Brq+InVEDj/
eKRKDgSLBkx2RO3D2qfwo0Lvj9yrNpJTnmmQ93Yv9x4WahCV+qCi2LpFQFnGnTjo
Ggu9SGbTDxSTcyt9grK2fzZxxW1gAPGGq0jD9gyfW14tTq/6VFuwb0DOsGj5IL7D
cBVeYjc9xrkbJtHZh3gJWki26ZRcBJIEk6g0d8wXCExsCSj6Ma4XgiunSC1CHY3S
5O2cSCCEwj5W/+T70uG7g3dcpBPE4SMAgbhubWOsDHW1EG0zO2iO4Em935ZGCFXM
n3NOePJ0AnyBpybRY70uD3iOPhIkLA+m85x4rcoAvcdSsrymYHnTsre3bwLgSM/n
pxNRFEps1F0lrIZmoofTP8u0YGfmlAif64En6V2zLhDM6sLrumsISLo87vdf8Z9T
LiyWsLURZc1/ieOZlJ38F+em+PkzJ4i+ji7J7mR2P9VOu6LGi8MqMtr5DApGIMkU
9015oI7JaglLt8aeL+R6/XYexk7O5A60qgs4rRVvLVLqnCIeFsR5ATB4OuiakEo1
f2dqrT7sle/3RVUgKMrML7AnX7vqpGy3z6DCANd6G+GQz2cNwB/Oi5UYQBuQKsyR
vKIyrVvHX6pwqF9irLuayRGvi/hvFxaXjA3vf+NTJfDZTpaWvhBDcKgaGm4m0f8v
ht9pCVo9+AX/GiLV+0trnPyu8dvXhuFHAcnLB4FpTCR28uOT/HYWOyNZ6ioyJfLS
JpV3wM/zzSVt/tzBCYz21P2IIflZ5mNpj/P5iJu4P7Oh+icSRcrmhGnKjvtUPeed
UQ/3nqA95t6xKxzwq/xy1rkw3tNudvj6Q+q1ROmZTUo1GOFyVRci/vYF3jVxJJHQ
I0t8DzrTJOZDkR3f+9mQJTt2R0zR9kCruXPMC50E0tkbwtzsbCvGZpsKEeMArH41
/z31qmj0tTwRSCj3EnacwooLSAwp8DnyUlb5XU5quIK2XcG2PM0Uu1gynagJgSjH
TRQZJZ1yTQu0IdPFKtGjmvn/gXhdJ6va5A1IXemEzX2HTSvrHwmDGPGUMlPDRcsH
tHz1SR5KqrQV16yjSVhyewFgDPbnCjqvOTyAbOdTSjWBk9fGELLdV2bSJ+j0qd+a
RilaWQkk1M5RsvC9p6dDyQD/TdAl1oTiIVeDj6YQoqvRO0XbimvYvZ8JQq+414a3
Y54T+sM20K1isGsK1foTLTymTkpFoX+mdpELWTIe5euqfHLVHz/ktpngo5IUPYp9
q8TS+sfNORwDQiZKwTqEUzyMYUvxDXB0jPoZwn5hQfLqmwAL99ZJxLjMQXLzc3D3
MQ8Tyrthnz3bIJCvY9baAfFJpHFWodidbp7U10FwWG9y06o4JAggHodhymNt25Js
GZ9nytzjk/S1hkoKYixtmKutlMC2hVeL2uUWlBEC8b/bf/wHaug0NkzRZa3TLNrk
vwSRkfgDNRdIYc+1MzGtlgdNswGHHZWX/t6nkD5PIqWfAoISiGYiyapfujr6Ccut
smUJClU/qDg7cduhPoaXrFrO5wPL7YpJqEOR2JfNhrfvpvlqM+CVEAFbj4qbAMWD
EqlxOJjPctB0Zcuflrcc3UamLqOwyF+lvIF15B1gNh/oZ0AKFJ5m5wqa4o/Knlrb
ON+/QesArQvKHmSd6YXD0WSC9M+QnvFfwDdsqacTyWFzh6ysVYUp9oHyLqfGESi6
7L39Np4/FumFHVtWX/PUdqiFCQ5Rwx6taBbCAK96VZyRvIfBg88IkeYbP6OheLvL
JM9OQMCAGp/DpXQ/8y6yE1KhroMrTPiWDD8NN2IshMECC7NPfNg9KENWIQbHysaW
w0zrL5OXevh9vPXnyhwNU8UgEVCeHc5xJWjD4W6I6KiFgHthn0JivJFzhkUhl5au
zfUhXmfRols0M87rsdvGdwdT/7/NsHpNW62OV5jJA/yv9Ymq61+HlI3F6lqWDVis
3wvyLz5QDjfTtnDFRqOxe1AnYgXgMRqjFKQe75nPLb+7OhlmZvfw1lw248KSVecg
Bc3YMqBruggR/AAloEfujdng4mtJ1/wG92dIvfH2yu/2tnHhhgmtgdUCVMjK5Dir
so6N/LjOuXsobOvKAJv8i6djDIX2TFI8nXuwsi4dId1pXX3dtbiHDP1RsYukgn2w
bdOB2ZE3bGaWHiihvfCGeCeDjzvpQQrX1vJa2s8NZSEAhPaLrSGpJljjDovqijYW
bJZrqsIRwRDBvFx3zipk7hnePuGYS6aiz4QNn4gk4mercMMwJNJhhG4AL1OYdeN6
jmDNdNplCSv8j/fGi1SAgRW4x4F9MGsCDvsJHOKmAOu+MJ+6JRyP0+zScd1Nw8bb
ggHvWUMCue0fzD2Mn+q2nElmeLGgmB4I0rtSA3IM916We+acOjuZfC7WTjIx14TR
swmd8xafbcnJhdpKYWPunS2f6soTrP9WeZ/1GMlwysXwFzfVt3oVNqBKx5Uw5TPT
N6T7vVIhcu4vS5xoB6GDhxGnvQ9ePXhfw5kzZpGdL/OV8XVHhXUYDDMslD1Eg7sR
Ku3194O6fkX/YkXAarb3FLvBxwSpk7qwen5/JGJZ5AVoyJto+TK7hQ4KwV5rxvBj
3N6zeSjEg4iP6luXedUg0q21XY+DFtnXU4fb+RswMw3kCwxYnzuwSbQpm85E8+pS
Oxndv2og3ILZUe8XBqkK5WPtLM6yozOpXllTyC/Kg010ANyb76s1LmC4reaGYLEE
QdR21tnwdtUoVe/PyQBhg2CtBNpEiJkVnz/dFDNuBjLK4eE8pKdtUHmh4ESCTduP
DihsvRY8a+TytUoitFlCf7lMcfEWQu3h/r0RGKX2NhWA4HOsn2ZtAaS5afDs3UJj
bMu2vW1/NzI6Ffhmd5Qy4JOGs1oShXVO0o1/FtRzLcN0NuOHliY8789svsiyyLUd
UV2yvJB1Y8wockExjITYBsoxc/FOooYJDsB4a1JIU+U8/VbtYMrtVIlsWNyVftlM
BeOOcp7ilFxSu9rJLowdEAcwpPaYLnL7oUB0NvWHV/e1IbzQ/cT2ga0Lqy6FI0LP
HAQs+GSBhjRMOYgMzyEabjLrGne6+2mCnlNwlE5etE04eRS2yZvbNIMJk46nZu3R
iHS7JS3HmJLdvyEsENhkjPj1VSQWBhKQZWd85yrwKej2c2zb5U0tOLrUsfoeph2A
FYa+TAOSqM5jglHzUAhr5C3+FAGaiQVPSQTKIF1GYWs6J/0EyYObVxwhRjOacMuS
6Z3HB2xz61k+dVFhoOGHXrC/s38Wv184mw0OLU1mRIppJAl8oNmQH4AlV38+/6al
wABqweytvPXUPafgtIHrSf6vQ6B2ifRl3Ha6/WDH80uhrYoRk4rKxbkm4DxKV/r+
DX0qOrBA53K/AgiVInIOjWe2wh5+FRCmILYVKmN3RE8GnS8YcixrPcz/K7bz/1nf
wT4MKKyCA7VWWaE+x0R4BurTBSB//mTohkIc30Arv74Gf5L1ekhDNnwqJaXAHt0n
Q1E9XYR28FdXYqmpsLwfnk7pDmjudBIcV/c41/eKXvM+2MGrl0r+VXGsGTwte791
NMmLtxHlAC4cTlDB5EpEAITYbdG5jmXnE8ckv3UxuMW0G0ZkuSsnck099C0oeT9R
u5VkRZfTuSmJekEucvIZjXsmS66ZeoN1GHma9UEFvjm0YKns4Wn2RpVYp8tJL4LB
rON87kPVLOMOK02AWQKd5alxObyQJ8iwiVd2TA5xdkur2lYhMIKTQDVLqo3hJkxP
Qjg/kGGDCjKNlRGQycavvu1LXrqii5xeUvMxkPYLSHElIq81a6XPCkOo0VdCM5F2
7yVBg+vGEIqOFZJ/O5oV0mXoKXMIw/joGTzyvfldw1OuJ9zqzPnkoX57nDfJGZGl
KN3wcZCMbgLF5P3ZcQp9cvqgd8G5kw0Dl0cPESyXHVKIUb9LY/fINIEgzc4Tx5jQ
OoOEq18JZ4Hkj1FBVwLhvwFPeYwghE84LDxpVRb+DpIuZmgFfNY8EdqQS9dY3VhA
l57hXJhw6toeDZsxEENEk+gAghsD8V59tdtlvukZ5VCaLWpGMnR/Y87vbtuFoBJG
1Mz6GlozOa4EPuhU43A9RM0jpyLcxZSTd8aUcinf7W39CFhJgML1vB3X98Lwgnj2
OBurbjm0ptT8O4SOSk/Cjh42kt1/Z7SPtJ4a7/Imfb9CNu2C9UlPcxKQSqMtcL/b
2xzHr/K631NbhayFlIsPX4n429eCVvs3lN6/hVCZeqWlG1GnYWWcSRlx++hhRkxe
qF100M9zqaUvkeMsKhcQpfPE/sI19ZQEptr0D2Sl0L3TW14KHiwHUQDI4ZeT16pQ
l+ezYpaelpX1bJuWfiwTKkPFiT0HJifUzJqX3ijjfoQx1Jg/IFcF1id37/xlVKVC
hFRa7Q6LcoeT8eGOviQCLD/8Jsvz1tzM9UEtjyrQdEUO6T3bMiu1YdAxVpnG9mfQ
XyFoNHoyUUQbi1hKf2BE6goBZSUwwCzboyKGzqKzPL5GrnwWIhO/b4YRo95/383U
uRfSrx0FLLEdnG9tkVs89c3roGnXETf0CbX4WENHfKjDMWjbxGl74gDZxPTPruOd
n9osDCBMxCaYxHiHMscqZNoN4h3UvKSQgsmK0iHQX8y0w5M8J1lss2ttvq9LRKl5
ocvI3wYzbDdWyFUewQWK5C+AgGovIl5Kkf1Xd6JHWI5Y88sVN+nYPozW+dpN6ADT
7FisMUczgBNPpoWK2CqJrJOlsMQFO9OuCtBWQnFQXR46UGAlVdu7V43EVw4PIk5V
8mByvf27a2q5kwQuzgsgDGRynjFwQ4VVmoQfg9NfFbJDSo19bYtZ/TC8CqbpImGS
vh9kVBC0SKFZ3m0Ojs+ARnnCOlLt391ssFLwF061UqSqi5ZqL6XRBznMvxbOurvJ
5KA+phf1i4mSc21v08fB4KLg/7PbsMcaOSWz3YdKXPkh4rN8JQAsri8tWUf11eZM
q+csCm4hnICdk5P4Auss7I0TYrbc14xkaa4QQDDF+389RIZkgIE4NRkDyKKX+SdA
1+N0oIydOXShpz+5lF/BWBojquGbRbKzQaEmG2D9Kfq+7Ca2WVLsTA+PqDYUm3m6
1qvRpzSY0MHypf6lKij16lH+vQexgfOmpTUJJiL62KXTEDk37O9FWecoW2OBHX/H
5Dk2p41ppUhppk98ihuAWesWmdN8wqz9o+YyvVKqFexnBMgxGdqvd3T7Di2HcuFR
q272b3y+S3yvaufIFc2cbXj8b8Q2zPFJlazrF+CXcer8+tH33Jg4bfOal1NVthae
MQhasqqbwbJRIweqTpif3cP+YtomNXnRHzCXyHde3lbo60IqieKtw+gB+89mJCja
HwTpXal2/59B8pLkxr0o+MpVMKZxZQN4rc6rtdnndBc0+gEmCWNUTxa7MUBndSAO
B/HqlXaItwbxvMTUOAXCy4M6lISqyPNvdghrqoK+hcibZ+dMiL2pHL/Jgp5JZ+90
NAjCQ5uFB5yQiTDOiDv6hZLKCUyLrGeMC1hZ2AgUYBcTjhSX/0sN6slZIbvtniyj
GDcMZI1tNG/VmChiIBNrg6oaAX7KzaKl83j2DRBDdPZxXvYRZzdgwPKUbjTHsw3w
nJM+GInX+qHuKUv7n9ncRKuNg59teWFJ648Czm3P8+hnjmqEPJyzNEXulqGYSZxR
tlTM74sut3CbK6Uy0Bx8prunuOdRadF8lMXMKLrqchmBgD6ey0DqzS/Bgotqy5u1
/lgspWj91gXmJ2V3+4a7I4HFMPqpJ8MCeCHiplfN3rr9GqHFpcaofZkEUakpcqg0
wpOrsVoMlOmCERydnim/37D3WpYPirJ4/iEssMml1Lq33pzYcYT/XZSyVm9aysqW
G2BxrtQDNYwIveqQlIqfAjLbd8/G2QNZVA9SvZTkAUgFpoNloaQ6mtGevQzlOyKD
kP0pbDDh86+D0WcHEMYahes7ZWY5zPOpdImSN/gDKwGdGR1s9MJB5i9Av0QmT8ty
WtAlGnBQF7C0fkW/bGDbnaOVvyZoC+dMARGSpj1X/GdGmTJJKg0eFu0xmim1oeU+
dyZl+2SzqYoWatFJGvj3iOklxI4lGxwxNVT2EayKhYKFjoLWWkEW0ZUmvYDADFKe
WnklECrKQIP/mqXGvtKuBc3I38zztGf2WBT6uaIJYXToNdPwNLKtFmyomdUYmgue
6JU8h1mZD190CJo+R4Vu/h6kAmhTU/sHCY4jBsbYHrXErRKctP7DczXUzreNc62G
hKee1eL8o2ZqUE92upTJembwG0VZPujKxmXarE1i0WNmBDG4GFK8naCVz/21LFGJ
HP8qjDvKeOBPqhYIVhcAJ74NUkETYLJOU69Cn2x5fAiTI2sp6OFMcPFHZU0K5aip
FzvVw6K5ZByF5OKz3CkPnK+6DOENAV6BV3PEEsCfGJ3E3QFUb9XWl1TeGgKRLRfH
MAo+3Zqh9OHGRgOijD1H9i/17C1Gg/EccqCwC0u/ZRnohxre/vQ0LuF36X635hXz
83bjDtBe4whZmfE+cJw3z3mUGwkm2RQBns9CkMDwAaZL7LD1vpADH8Zeb1IKUEOL
jxnK7x2I5HRDe6UaZsyPgHyn7PDgGkX6XKMPOyLh3yAkIQmG6uFu4lEGYkuVSBi5
cVMoQsKNb2SmNlgsuOzMa1zJCVDtRoozcWMORl9gZErX718MgEd4grpZGn/9aSca
rVHxB4OHO5q3esicWaGxZez4kfcyytIyCTTBjNxJNUcE+759J4i/jccKCjltN9vo
g4zEsqRVyKoV2ODZmHCObFH82YXqYlB1lAtRuqqGWVSucBpRfSbF7VPKyOprZnk9
TWBnFUDRQVEHfIavjW3AM+Pvi4MFpxR6so1iYqK2qHT/WhCvMb6vT92DA05zUWzz
/4vMph6m2bEnI964qyR/UwqnsKeM7wUKIDDVtK3sX8yeokmA2E/tf+CtWUslV4XD
8+qt4hTcfMk2VumAotpBWHa59XceCr2tt3DMoW9O7MvwD/qOxjzQ6Qy1M61rlf1c
QC9JfifJhqy3AczkWANfg8AytnBguR5U1ilMYWY4w840iQ6dY2y/DJ0ASCHGvdTg
4fqrOqwK40VAK3gKfMXN02ZW66DCyTEnQ42zV91IQp+HxA6Y7blyweB34EMf6UHN
MHI5vz2XHFyAo91IpgBhh99lkO9SMrI27DbfJeismpE7mVTZUwMC2sJ/8RTtaWpR
uzd7s12UNfI6NlSt7I1FvAuYscy8BgHh6WDZiDCx/NInSc0IxDtesD3td1HOAt6p
6FvH6hFho1dK4LNbpC898WABr1mKXCapcDdqwcJ+VU1Z9+ZpdZasNWzQm5fzQWEF
drHbhV3ydZ1Amt2lDKzduHZ2N3VOJlzNTFShW3dMGyk8GfNVXc4Vv9a8dkHwooAf
4aSoMNgGBGehcD6HdJZEjEunUqTmJuaGxE18nBQz7Gk0M8Ls7cf5oO1QegkYYHql
Fr1Qw+9qqwmkgZosiVp2Y+8yrmpKfgd4YsPWQcJZ/uT9axQ1f24rEETZXZ/LTOLv
wpWPBR7L3ADQRk+giBlGWcSqrBzTWSteiQsbEVN4YMCOWJ76Z+7GLYXmVNXrUjHg
F7TNj+p5s6TlwWilcVbvrJEoKa6uqokVEjNOdidDJzUSnWM9n4uVJWK15z+HDi3j
qn0wn5gVtUzcNY/jX05KkOje14BcEa0Dd1O786pWLrzFBze5Azjr8rvhzsbfZgAh
wO2zNgg93CnVtvtbEip8mWOHvizfdgcbzGTgxdXO5L0oDUWvEYYat9q3pvL3y5CZ
EELQbo4nxPIteIaW3VQGcTcmRv1DDKR14lqFi1MXzKSWz1xEftdTP1MJT5TG8Yiy
3DhNZ8nefP1T7G26B7nKjDn88/oBItq6u5x3a/vk43c3K5idxW+u+JEcWf+TRBzN
L7xDoOMN1V5iZfY5I7VPhIGWK4Od2u1AzLCevjFNI3G8LkekiTzCi4HDOwF3SPt8
nWGLkcmpqTNjY5s/oKEm3o62fGbku7n3LK3iLRVD3cURxfZWaTym4lP7FXg+Rbpt
JIrq58dfQcWVktu1MKRbFuiiCFiHytyfDwD17KbMi6AheNyBCx8/x+ctfquFsQjg
eQnqCb0Bo5UGHdUuXrIUzZZAAyIsEf3MzNki8jbUu7l3vbk/UAtpa3GWMfBzPJZk
MGsFtV2f056tvU3SD7hgQ/3XTaQvRdSCNmuwOIWjA6ojE+kVr9L1/NB/ZZfoy/bY
9ukQfvFG/dLOn5FkMsK2Ok1THiMcMOFF8oalK14VFYhTZ96SkMmpnGy/1OgBihbq
jSYrKd8ARQP+wh6TY/eu7AzJg8+VJDWVQmEdeIpKzejk9iAxPterhdOJwA+tzrD5
xI6S3O99mMYDLWnh7UbDeMJIQ8fir5Qv0k+U9tj7nbRxRh+nZAf/M1Mz/L3H5urP
f/TmmC9V03Y3Vf5fc2KzIzD0d/m4Y92HAPJY5Cz/w1649EDzBA49qnsp1qNcU366
aO/fclBOjfeDzXlUBbHWUegRmAgG6KcwF0/q13XpSvIVGRcnCKttRn00m+q44anp
KL4HzZmyPOlF3zTMbH8C9ftKNID9L5SCHmAQycWaw9J9tcQ8E+cZ0dq/XlwQRd6N
jKriJfb8A+251JAaRRAJGN9MTg0gEgndaB7oyXvjE6kxCYkNTy5sw96Q2SVXIbPk
YRW/4rnB4BMb/LggiC+mzKdr+wweQwFxc8YZQ7W/DcAczo7CABAAW1nPd9ky9FFK
dvbJ/QYR2DN8GNWzo7Dvm90GXLHXqhbiRv4FMkGks0HYiv/R+n2cRxFwvPTjzcNO
864hdZJjrE5rXQXFPMj4ncWwEfYwmLwSHqxDg3LdFHDyOfM9IfTAn0+hannQjeLg
Lq0j19qG/enB0K0MvVT7DAgC1fWT+xRAhrJQGceIkgcFjalVoCo4RBOM0bpXlvPX
HhLSIGqzMpjJMrsQy4EB20r2sH/4urID8Yqg28hiPeed9Or7Tc7thnHvsZBecanz
AI6SR6dhpQX63x1Aelk8lyWxTQChUjuO+gsFvImYVbqDZecPY593+1XHISsLLdte
ANQM7I+9pYfDgH8JoLn524Z3W6d99MDfaGl0sWHv8z2qp92cnpEWg0Ix66n90B5V
9BoHLWWmy3Zof5FnqSNY0hzfqhvT195vPh9zzOQ664/+ZdDc7qrOytga6vmObpI5
1m3RVARHip48INfKsdDth/o4gzeaAzQEcWoaLsVIopYKZmodbPcJHz7yEYXCSvRN
qjuK1qFkAhCfWBGRA3D6Fnz8ay7vTOAkt609l3nkOzrRtBiPbffxcpU4bnJ5kfTk
8aULdcMo3DODmh7oj30367gjSTBAWSMEMl5I3UrGVZmJHLNH/Kz+hbTTogIwtBa0
b5NpkaZ46k14SUrvGQLX0TDUx67k+5H2gKJJzxWBiAG4HeLl9HaMO8WuLEbWm8Z4
B1QIEdMkEY/A4UZm3k3OFrwrFk0JPAqtXmNQrQrPZ59Qzv0C6RLa9s0pSjdsgL/E
LDe/W35mp2BlIMWBmwGT2JF+PDy03XOuM3Eb7ye0IUcq+vipFJfEW4hoSCi69Ffy
1CTJsdG6vqQ6bxODsemFj6g8AASYgPMyztA938K/WsDolTxRGZyWOIrldHAM1cpd
ex2s/dMbU6zZNSQwiLhb601eBt0gI+BRMZJUCjnP58a6S5FVTS6DvBOwuHBOHkYh
tVs7rs+fRl+6zpEkM0r1m4htD4F9/uNM6LrgIfZS2HzCPftEtytFYFxBx5A2k40o
zOjTeWKMZwErvQgf9Jg7siicPMWK8CI+/EUXl1DeK2LIL8TpRfHydHk9wyk98kzi
mOMSafsGOmxhMnCCnLDWgJvZczCU9dgg+a6qHK08lVR3Z9cv/51J+2enDnzepQbA
f5xNMHswyxn873tmimBG9SYXBVwbRIK8Ppisb/e4XPD4gi9ivUI3qbClTNVwCtdT
shnejvFhCB1G8tm0m8FO0sQzHAHl60MW7J9JKAvho1+umba5y7W11+P1VDOom0Ui
ZXQHfJNVBty3Tbhre1lGDVlapoIQAIMmjChNqbhL9dpVZOhGgIJdsqtQvv68I7Nt
rVN2SBGaKX4Dl2gjq2i+njnbImJhFEp5PqVv5Bd0UfKKQydznZRJXykGBjSQvwyc
9vckoGhhARK6ZzjZujR0cmvdq4yHIjiAALgwgzGRe3Nv6LknxfzE9nrxTS9a0TZe
d3WrUOeFByP7c0FQyv9CBgqhnow6L3vBSOWuQYVsr1DWtD76KR5CHww08o4QX5RW
W3MYWn7Dmti0Bo/gNituf33cgFUBOP82w4YxQcr55+3+VsMMumL3C/0yYQZp5+zk
+sgKV14e+TEavCxo7ZUA1jqKCt9xoJQIQVpq+a3nwkYjiUFbOv0nvlkMSxUUqJwu
wQ/HVWLnsrx/IDuwuK17EzqxjvkpHjwikGd9TzrenVqXgW12pgjiasK7Ppp+qO4S
7X9e/XOJpyphZHlq5o2EpzHf3OqWqx64gpp+2GvpqyBHe9zjaeh3VHK3ThFYAff0
QyD0Noz3CDM4xmQtPp3nwWcl3PW5hDg0fF8xiYnqYlCi5Ls134adhWLqGmtsu1Ti
QmhcMF2fQrckiqeYVxgYFiS6Hd+KxAG4/ESGuoqwEpYOZZe9hFk+QkOKiB7J+Zmz
dlma0HToNrGrDgE2dOgqxJJb077W/9PoSewHadEyCUIzTyQyWQXPqPohRx6dCNz4
nkai++b5/GL2IZ3dxeb1vPt9Mc/SmIZbbLJ5Nd+LwamYRUYX/9J0ydtFk3XWOLBr
CP8SXVWgPD5rO8PmV0Rrs0OSSvMOupeisOlHkeu7MSpbDe/RaIJrjKC6IYKKMvGR
9XXnbJzz9pqVl7MX8zDFVOsvcZyHoSinNum59GlVySlzX9CVK9AvEvIxc64sdbVS
cnNsbX27a2HAhiNH0MRegaiAL5APZNma2gpeDkiAdtCFpiNeqscmdT+i9fYD2ZHA
XOoz5DHixRaHvtktU29qjjHWWcS0Cdi7Z52TO866cmb++av1SWzrTbUb1LBp2FZv
X/Ymlk+g3ym7LvQi4VlufioeQ/newZNUhJM5MQLE+dQPh/xnaMxuG+WkIDA0pvSq
CmpYkjYamvvUPNpMYTEMH9L4ij0xddWUN7H8lnx4JGnTKg/5YhVedpmQogtZoTw0
0nDUuczl3SkWaHzZMse++9B7IF7Z1w9ldGT547VAgAMUPqAraETxp5EJUpZG2GRG
GlWkrDoMchJezQtQF/JezGqRYNS7My3NIYWUTqreiEXuEx2dTLV1w3XwwYA79yex
8WASVkoOBcuu5rM5nrxprzJ25msCPsTfeMkkfP2knMQ/YMNU87KyKaNHRvY5/26c
fb4Ddnz2KlKDVdGC8bza+sPxBZWk4XZkXv4ZS9RNFQOfNqu0VDy8j5VoqUhCZx3v
wiZoIgDGplx81nLbjGQxrFBcR2kl4B+WrgyJ5TJRFdGxjuG5mJIciZFi/KahTrDx
OWuH9YQ/VWtCTppGGNM98ced5PKNywe/PvMjChrWCg2+YGAp2fz3anLE08sWbZpi
dZQhUrqKu5BGHRJ1RYBXVffPoUCBg7q0vokZP6dWPaArIH0qz3Hqw+JwBAexzywn
zGQkgQ4NMb+C9Hg8xQiyGmKajmK44E6zYBxHl9R8EPMGVL8ZbHCiS0IG0QIKdafw
Icyo89mu9ie5X67zrChMgoRkaRgT6JzAb0g77NrFnSkYyaqbe5PlXhEr706DGNTd
Ou9QRp+K9QcUrhdrlBGGLhCsX/H1Mvh4704nwlqDBpU3wZgKoF8gWsZY5F5eNHjx
0rBpxo9J5Lkc8VFbgUyoGsIH4ojupfiawxACgFKWZ1OiFi4eaQOWqvHYrcMq2ePe
EmxMoXY4YGDAcNhIGZf7FBlVpYvYwm5QUirKMIEeDik9BqHvH0Gu163ou776AxSE
pyH81r4JnAjq35c5xZRhB0xShbs0gsbZq2KEadmVBDk7csRGjpQQRNDAK88Ssevv
TN5OQlRxWWJTuWXyLXLbkMK81qbOvL6tVbTLkBWPyr9BwNEEO0XsfQfmSsvBJlra
S0OstzDQx0Kmgy9oSuw8jxeDBfnia+bgnW9b3i1inuQDHpzyLEKlwY7NI51r2NKZ
xworIA8fGOUl+YtlZADVAug3kKplrvHgsHssieQQO4i/WJV+kR/8MMhK/ph/tXPg
ut+ji/+Fe90MI7VdE7g19evQ8HEWlP339qYgCpaGSa0P1ze9aB9TbeVn+DqxEbqL
+4Wg8yJluQOFvpVjJONFnlEhLQbAoY8oj/2VZEOYb11sVO6esoJhjdvAk3969T8p
iLVjNUqF/leBZxIuoG58I7K+8ZrbZDo3nSJ4GAWRR4iq0rOsCg4InAD43i3CRS95
GfsqKYhqRRllGtcQ3uZo5FDgcWCXLJFBw2JpZKYLoPLdLUGT4bdWMGFajIret9WF
kD7+SPDDsT0fIw61OHmckOa8MCSSzmjkr22xwJIlEsibzICyG+t2QR8amAxUSd96
nOad02+IwzxYr1FLFK5i8ok20SFwuoguNqQKCosxJwNSzUyNt8Qbu8iCkPuOl5yj
aEq9TSBn/mK1uP0AJQ3Mp0XGJfm4qHSgt+wMBp9yNAuLS7eB/hMR8cEaDU8sO03P
rre2EKyNC/q4W+2emnP7yNkL0ny82p6VD0BKssHj4SsvdNw8Ilpl6dSfInlmHlTJ
YprPcJS6qTxi5k/po4PZH7bf6vPXBDr4ulvtV2lcNTUqCEAFEF7TX2bQTeq0/e+U
E13+73ftbmWSWHJ3ybEuuAxW2eZuw1Xrx2rnVI/MUMprJSm1n0+sbvtkoWle1XhH
WCL+Hmhe+6BLD8QF074KypYDJJSmVUFvbul1LL3Ta6rS2p93oazqrGoFrCQNzgPh
XOv9h726j4p18jEvbrIP8ySdRY8Y3RyPShRvBN8dhlWdJQCQ+d3tlTbnOe9Op+eF
zV6tNmMh4kAz8kOEcUEjt/whIUONiEyVX6KlZiHusrDC7mEHkSEr+v7ADqME1emv
99S7Kr6KDtsBQRzJIBBkNcwnd5y06NSyr86WlVlTXqMvs8AQ8irfFUwoMe/AWaOm
m6dylntuIV4pDxftFgUkAyoZ2w7eYErnL3Qc5XCh02FtTiDGV5Xfkv1Za+XNSJG2
/P/+imAK7snxH2cT0KglbYrSRLxfHiUqU2SaZB7erm5nThYINMmGYPE/3AVE1t+8
jcCkaeIpP7kEUDPLlefpE9G2NGT9qoOcW3czhCMA8Ob58f3NegiMZnU85ZGxhfFb
92tcgeuhhxMgkCMcW7jAycvftkEHYwUGgcQwg5g3imLnOcx+d5sb1Rn9BcaI7Y3Y
0abLxt+siTuHnJhlo0R/bvHuN6thKQpeIvIC6rWU9UYOuxNMLEL9oeuJhhVk/V6a
gSYQhKOlEEbzDh9bENe9QwIRIpn1syzHMFrgo6EJEiYOknM02WR5MZgPYNLI7nuu
4q7gS+vxI0jCWml5tIk3PImawimZBtHE0uaaLUpCGdroLoHZWqECwe9TEdXerMjO
zgI4ldIOWqqsGKR94+X63WHmFOLTkl/tcgK4sTgUhNhJspUXe9jbZKCheCtFlyya
4gFmcIx6dI/CVqNKn2o1pm+iVvxmm5VVZlRDkKKZQXNJAevvbypajExaQGl9wW9x
v/WZeAzDZ81zW4JtpBiwH+wWIHfQl6jxQEuRTjVg44QXtdka6q9aRpns1d2OZjR9
MX3Zx/KYSX6DIpp242R4m/8ki3uq01PUSvMWxDdFBR07Qe0+6CITHJ02dD1dLfwk
fHxK+2lluk/9CXJsbkwkC0tF+2RL4g/hfmVIq3O2ChkT2uCqznFH4bXSlN6CgRFF
9nF6crxOTp/jkiiubX6Fe7mxdc7iYXc+hlNGEdQZUTUM+RvgP6ODtYcOTVOaZtCE
TiDNWelGfpYTtvkKxFYxNtd5VSguQ41Qxr7k5GI0EM1n1Km6eQffAupuh3FrzkUO
hXuXFSM7nO+VeyPoOwgZO5+fDK4VMrLl91rif3MbTalR+N6qA62M+w89K7SpmtZP
WkOHNvnPb1tXOMNfD7c/bRupif7Mrdd/VWxNz14q1x+YY4WNiVcMdqNAou8f8vi+
N9IkmPUGCFb3og+Kf2cSUdQSW+7Vt1VWzsizXpBFX+oBAQiRY3s7PqJtFciNhNSS
8s+83CQa7YNQDjquR48pVDKXiI7YYKIRU3WFnrlSX48IO8pAzzLv7QPmfhHhb+9u
WfkvTRLX2I/fePjj9pcjg2WrVpOBijM1AQZD9l7aeUzPo2TH66AtE0XSFtz6P57U
A538kEuUCrfzCUAoE3/3OTH5lkVKfBIATnT5MwzoWcTR6QtPcmLf8nBRKKbzIyQx
wHdUYn7rebOVv2YSMz0m6dD7m7MKGO2W5h21T0dYzSjXvLu23lRFIo+cWBiUIRZ9
bIC8lwcQrz2Tov7nmhWI+emMqyT6Gi1IlfiyNzQuekkaA+/fbvC/xP7wjoSAbcIJ
VzxvDEOFoCQY3xGZgQBH9efyRgwkndG/S8dOc3PtMRVFbY9j9ENtJGnPJ6LOExlc
eN2RWa1Z+E9QE1dACRueyd9QOQ/iVNj/pQ/g4T7AKa9Rs7gDu0nM1vCv6JWqfCh6
42LrrAK0t937xu8SQUJWhgTjad3bC4HKu0cL2ZclglioqLRtQMFzcLT8Y5VFEYL1
CeDSCD3zPRuWAy0XD95r1CV+DadZfZgLDA/LIClduCHKypToAND68sifRRLiGYZo
IfBj6+etl8GwFlFej1VLpNdx9jhZxjEk9t+T7SkqB35Yb1G9nRgS+xsHFzsil92m
rXsDclp2tYx6nk5h2vlJKbxOp0T9fo/p+Yf9VSSLKIbK4UUn8TUCV2kRCztek0pm
cEPEFpBpi7F/b/KOHWOM4PBK6D410Onacr3lBD2Pt/M4p1IyMoxzHUHVgaL3l7Ih
/6AnGq1C88/D6U+lxuUyD/cThW41HkzLD+eJJf5mOi0FZtIZyE6I4oaQwBDrbB+0
KfKkftlVrMSat9uYYyf2q4gBFE2PEHIoZc68P5EzvJfq8RSK3SYpfclj8eSs9ORc
H4vWujicljpFb9WgDXZnVDG5o7+fOfLJ49dn7Bw/Wq+x8LAH3yOFxrXF9CX12T3X
SY/8fVLVyslHj57KELMFla/xCWo+E6r8pjWatBbrGFrkgWV23Tll2WNgeaNHXoMX
nn79pvyoGwoOP3CYue3zapLH13N9k1sB2uIw5NO4qT9nhlEd9ZuL8zC1Y5Xih27m
JJdXA+K6JfH82ljIVY6oFRFwK8VUJXFJJftWu67PCCKfAl+X5DXbiJNR88rmu+TT
Ex6JuyL/XK2Uy5a1uTxEYTGwq5EZDEBNXHqY4Uso1jjXBhIHtlJDcD6itCVwfKCs
iJSLVSdpzi10TiX/PCP14h8fClSgzU3d7SFFxO0o11gHVHHQQAz3NCwy1jvkJBOf
m95ytA+sSkonYh7PQaTZKEqyOpkIGxb/pXehIySMrnhj7pcSffRxzZ+mM/jrOuP1
a/pxxCcT2e5qRJkQWMB/eOIoS/klYezdsCCaUnZuE4gQBSn2tt0P6i1Yf3kFa+ja
UHZRQWRv4yoh5Tn+tKVkT5W0tvwBaCr/ZubTmqe4h2Hn6SKPTGqB2E2QBE7c8lDi
AevCg/XzsVHdZhwgUqyO9ew4dKoJ8O4P4sGwnPD6T7EaUTajwCdiT7mYgA+XMArc
33FBUp1tp5slT2JQ34+59GjF8xPICZSJt2wit+T7sPqSxjcngVCur8xMEgyBqcC/
LI4kDgxGnNq77TbbQNAKOAlg67/0bZhP6VvUBxj42RoikJpPE9KIwNHY2hs3dhAL
JY3ksy45cCp4z2VdtywsmDpredd2iqU7DSPrFmeITknuAlClLuXjZKnMIOuxk5rb
Ll1p0ZEfH6g7C9yQu9bPua3mbzohzoi9VVN2ZE24B2LmNUeII8R0VnXhYYhaaEPY
ZcuGgy2f2IvouNHTSyEaCIvgBudou2jCsUghhp9rRqROUGpsppo/+qCAMKesM6Af
qJMdDAaLr1LAgMWPnVUy6Yoh1JUw6jPareGonA8gpcsPe9EwNtxrOWpICYI7X5aY
G8IJrsjC4wCaOYdxfpchW6ELIFHt8qQN9Gj6gCRMeEu/YSgfuSHTCwpiCfKCH5hx
aAGzvvAlEUZu1A8df2tOCixBZkXIkbat0t/sIrVmTt468BsDygCyJFNacno3TakE
KHTe8DX+OzEJdPRNowDkQ/UHvOODtD76CJmBmXqN91h+qrAnGQMyhs30pW7Q9368
AGPohA2Wy0kLohcgOnjd/zU6oPjwMpPAw9eB5xTuvRNDXJzUsF2K5Z/cvN6UyUzl
g3jnkhJ6VVB/DWj4fBG11XsalU9/JOlCQgHWrtPX7fcFuwXxbioOuxG1lDr7/dnd
ESy26RXKA3lmijACXHJRD4S3V+TtT7dytSAKf4vZCzVbP98s7WEiUz4IAc76HeD9
e/XeiYDKhGw9dykw6JOGaOTqz3O3G/8FGiUqdO/EfIzcbIb3/dBTsOlSJvrgFxTm
bbDHSscJ67M3AMge97lSkuAVvhBt/FaVXutdPVzU3KfCKYazykui2IZY/en3F87h
twMgJf7SBZPzlvEg8z98ljDwB7q3DH65ccCE7cv2gTJv8JNiPswJutmOJzQq08LK
q1BgHqRmzPV2SMuTEg9dUIAVWoOB7LU1KrcDTbsgoLRwWWW623uvS6nAf6G8wlfD
BtTRcTF7gUtlF8mEx47Xa5fQQ7PjBN1AOqCaIsTPeuHv3Rah7+4fWDE5DqUrBfwL
3VRfa7MLR76wj9A224X0wQn7B5BcN+UzRzks1O3fGL0awqYFmv6NnUnCQUjLIaC8
7FiUkhh4hgWxtmcFPa0m8oTckbwv25XLIzvsBa6iLrDCdnkoPiBEs6hkSWQYYuDO
g7v9Lraa6Y41ahhhoxJ0sSF6VcfpYRc5KHWyLUNNXvOM5nnoCdroUJRyF2hkiFkr
+ajqmo7Z9ZuWLP2SwBZEwdvs+pzpbeaMeqAzCbkIBQK8FwVJLEza78jo/fyKFIp+
ol6+1qfaCqVxpFPoeY/tT670DwrF67NWheo4TC1/5Jq0WuMYQG5h6bt+rgJTjoeE
2d9H+Ww0wZziWF5S6amswV+kWAcf5c+Vpw4tP2jQXzpWAX+HuzZ17Z/SehUJ42tO
wVjK9nYLgaHCUPVIx/dxUBVCJSGVF9LHZP1wBV25iwQqmLxg6uGwKm59fcctpN4z
1rUPif45tA1eUiKBUty9CGUZ0uDfskX+ogHGUDtly+93vV8lcgFRIZVbBDbUv3tN
mgqShZpYlpzTu+Y1zVD3uisUtMOTTAOpS+40oXntKfy48JKTfYIqzbV979yvXltv
1WNge38GICzFlBPhlZMUgBnEkru3DhwvXz56FW3S4Pvt+7lON98NcbbIBlAlydTB
XPxAkBrnNZQbD3O36rTXOjQMn6GLVZ0syNr6SrUCyLkmv9ZQ5/QcgXMIgGUIYusm
opDaTnCuLvZXVDGpUF4qnNB1Z+THbZPC9YvTwl/kYobi2GvN0h4JP+vcqOm5Kb55
rTnN1fdkK4sEqRdDQob0ZOfy1nU5849oI272nxpZRk41C/U+c82k2qkj0P2SHxkV
582POEhRrLLVjWzCZ3WAg8g6S/yh1aqH7Orqc/omkiB9JeyMES4mucSRgAOVq/CS
NiVQNoPhkZqsSusnWcrDTGrmyDCpbBgIV6RHJn5266koKWD6YKG1PX6UgKUM7AEP
/eARnwZgw5ZXTzWUwTeTvMIKQU9tYc/2q3S5Ov8EJUzJiPUJugonTPYr+7Nh2Bd2
bcF8n/Lo+mt8A4LJPqw05SFAlsCjlntCiPRWr8L0/2BD7G2S7sKN0qXf25gkACbr
DT+vGC7ubGU0imZi8rEkOWWwpIyrHgfFND7+lCR2fMUMODTSVGZ27qjwiAK0jfmD
GRCKrObPyJrBaqJYzNySIijzd9rl4gylqjncUgKUzsBgcyt3TVM3ZT/y32CJHQnU
8zuNTkanpHoKpr9RWXVm47tCUvaQwjRm963ItOrIBwb5vKt4/zrgKX09/HOHxHR+
7M8Q0J7wAhnpm1jQ8Knefh93DbIHBho3oBn+8Me6jhn83kSEKK3pE4h6QqTwWPs9
ZRD5yeowbCqChdSS+CaoDcc2faTi3f8/xT0lvX/LADtnnyUgEdYAInikJtcXyU+y
6cHcpdq+flYbmvTbVzYcyi/1TDols/EFNzTldVxa/vNYp4E+eWPH1UxX42BRAXJ2
x2Mb5OtcuJt6I8i6TQP+U5lNcVetHuXJzlzssx1CpZmPBh2DYA70A9M4wysWGGe0
XPiLrodhpoSSFZgOa/d1Kb/FkYSDGw6q1JOQXzlEEm7poKwzgK5VtvFqvyn9aTfu
7i0hs8ajZKEXNCPO4EIxJ0SfmQDhi6KQaH46nObcdYQH6Mo9a9GNJJrEdOuA9Hsx
7uvW4BoZ8rFcrFD0vRuUUxaXI7Ktquv8rwL0AGlG0j57GgCf0WWeTFc6WcaJFOhW
ybqm0ND/+q2Hdk2d32u/O7T+nYn4fGJs49UVf1BJJlxr0SDWTGj9pICu3gjgMWDQ
7H/gnRSftAn9L1oGqFUc3vY7gXhXdgliSfm8QhW+WPHfCtLgIEpJ+80NWzCNmGaS
8/d3fTHKYzKv/9/4GVkgDJhCzmg7sI19FRsGCtyX53aw/HtajcNQ2ZtLeOQsLQo8
K/gpD4qK+R/z3yKxZ5EEhSGrp4ifTpHpCdb0ltvdyGguqqTMel7+ofn0plCPJFXx
OSX7KdvPIus8wSrUQWzijfctOpWDHeTCiiE66Ns4cMG5dBPhypWFA4ZfpxFtvui9
+aInPPKs6sMMxrMG0FXKgiQvcr7lhIX0R8LFf3sqzyYB9FKcPWyb3mCM8jEyeO6p
dRY/4ayGeNAx1UQY+jsexwRXkGDHAS2+DTIIXyvIIJoeKZUxUhkvUTd1F3PV9YZE
4MPmM1lGlXghGbfrcCsXxfqmARZCwQnTJOkfoOtrcamguhri0f3UNs58QgzCmsXB
CBsJtS+ZMfsoStBBOkEPpH2j79f48SWyzrLY/ZSEXNUpatEg5/IRTeYwE+FOIjQI
70DOq/js1dZTjNypqgufvCjCz9wLIYzpx2nq0BEMnbGQ3GodGX2UdNpE1mQ1t6J6
rStNvz+4vdzpZK46C24BphE0xq0Q7bFYX8Ad5me8eHpyGpdk4sCd/WugKUWWfH8N
nOuEiXHoN8ovFBZI6nM767j/ARzTosUTKF+PQ4SvhisC7R9JB4q43tiCWXGH5z0a
Yl8aopFeX4oCNeiuNY1w3H5esg4/kfiW290TDSx9RKhK7GWD7F94Ruu9qEHbGTdL
S73s3ncXhgYipWKuwSiFyEQtMhkm0atLr6DgpNZQ7qlDIiZH3rCUq+vM0yyKEQo5
YMWHuGXJz6J4mqBGfWU4cnzmYwcjcHT1Sl+8+v9bOUPChSMiDSyZDfdTUiKcYEND
aLbbbUIdHOpXRgFLHuJr9IKpUdYEii7ouumY83LcnMqbkh/ViCMF5iawFqOWwHYt
T3MvgsBIJyGi2UKTwHpuMbcqdVHNQT9FbQd9a2UrAqQFkIYvm7eZf0ehmMPWLexv
z6FLLTz1pBrapKAKzOvn0Fs2l3Tio0U8K9bEIh8B+S5Ww2eL6/LX1K/2NSbARGL9
ToNS+zPMIey9sYZQuhQY0dlvMbU/g/NBovpEJRb2e7XqXqS4B3kt67ARj9PIzvsL
MQhr0Q+eak6eCDqhmpjZfA6MIRrV/bLZd9eJ/biOyvgdxx5Q28ieEyeKUUB1xOQp
F2sSQoUnLfsm8lDSgY+IQT3fNO0JVqbfNqCsuICYeEuACcgUb1oHyESb5QQAR6PB
dw8gk4xDH4aT8m/HiLzh/yy4vNH8OjHQwOPOEa/q7W9ddEbVy/Hzuots8uEc0tPz
W4SO+iQe0HK6ZUbmDgSyciNSxUDiXSnmX7KeW8SZCgrQlahHUdMFBZBVA4LdCOgp
WmRfv2bA9o5depPtF5hsPNa2VvArAGOZ3SAofQxYcDl2QEmQi9jikr2BcIfnkgvP
mWWZLZSoB1/2+hAHLb97ForR1DRoo+8GrPtqfCSNoZdTiN9QDWfpHFUy8RH2/nVw
DSs0LJqzlw3eFWBg/h58WyOyE1QQPHuzSqBxyOPdnVWQ3ZfO0+14q9G7PPsOuVD1
HL9HTET82XsIdVTN+ylGzWLuqhpY5+ypmVsmCnqXl+/A3m/6BBCjOWbfb+NLELRl
OPlb2c14cjM9YcEGFRJ1RKfFzVdrDVuofohnEEZBA9kHwVbcYJPNtbBkh3Dyi5wd
XgNFNdWG3aWOhUnYUCGZrCT1S4kclrNAY2YTLanK46sekwY7jQSxCd+oBnE8PGoa
ZUGxgIDDk19k9jRKzDSoylgVWhmgNbWSuJCX5pQN+oCRLCh0fzyb1SX9Q9sxakOY
88MRRVeNppmxpf1EfF8JQC8CiEYiwyK6ojvBKpRvxxKF9FfJpQp9Nh/ECBAAapgC
pugk9HQ5GzHSzsm4XiDYSAJK6sUTgQq7dMTInJcZaoz8RvgeZb4BuBZTTDwBylzl
Eu4P1aU1Xzmywh/9n5qx01eECaad+zAXaMJI5OhX5QeOlXVVJurZRyvYAKjqsIqG
4M3JZFvAbdrTw8uGnaPm57q/jtG3LFa2O8sAw67NtXezxLWwtAEzwzGQG9g2wmws
m9dvpRX/X1gYS3G5lgzSonrnxzVlPt+NUdf/k2feqoRiJgKJQE6nCOYg+IXkJPuM
J+qVXFleA4tjYsAOxJ448m04A5wL1HMy1ErZx656IZBV4+jEd0Knb7eepplpcAKg
sjEVFwXH2ykHxUxJGRrR5CPqYEdcsNBuhg8TK9DZkLiJFRpyUobwpOJJFfAIYURu
6uXGp+dN2t+kaPGeHZZrmyWEP23oryV4cvqOHzGQsA6pS9hPRYBrmBNXTq+8hl3U
imuIdafUI7HZbOuor05aMFFE3aYb58XXHmu7QDEOvDcnn17LDZQkC74yhY2iK+S+
laHUngIaJab0O2ty8gzV1BnGzxMu4J2P211Prx9V8hnKOnpjR7Gpo+U/CyaR/AcA
/EcY4lweUME6ulMFq/LMfXIp76hJkZ4xe67LiKnBkIZ6M+opWEdbkQabmGkYQr+O
AnhqjlcoR+fS/fEbUMQotWXgnE0Jl3N0kAVdHJCFBi58+CsZtIrlFHApnRhwS3zQ
Hj7WxhoNJtKqGguijkUlgOjKI4nlkuh7aWX7vLchF7IwBJQumEHLTTIP8mZcKGOx
nAxxDQNhmfLxaaZlJhNx5EZ0uaqVqoiTOtQoyYtl6DraiOz08BGyRABLNgOQIrsJ
NrAjoXZR5R9JO10ogeIpNTHuci1RCEHe7dqJnydu34PysX0E6uxevTTQvgXMN6hc
Kb9cq1ERP43uTSSeG40Wjyf1kjs7c3kShOcU+HNiuihbELAKulN0fvEgbTdOpMhr
KZr3dhqpZ4SWziRU+mrcaL8Obwtl9GDIbigImPsQV7fTn5Sckad7hKhJuprwRZqJ
8zAjX2xZWGsQCA9ZrqI0dPMr4lumRcpLrO2rXkgC8nEbl4uNVjEiYF6e5F4HxzlB
dz9m3TbwxYyh2nFI4G8k4a4h4cs0Hj++lgC+90qHvzKENEYEAU/ABndJX+xIW+Ea
1nurhR0Kts6kJTG3b7GOtZSNL4kz2CAsuaA0I3hGPlVvpyi4ukFFzPxTkgc5rpdh
vOTWHlssBGq3D75tZGavW1Mzzh3KhpMAGTkeoh4F3BYOVyu20u8aw1/1MrlwNRXc
i89MFs8gnkRTjof/e+hBaJxn3BNv+IlkjZyzL86t1VwB9Hdt1NsxdJDVAOvWCSrS
Db5RROieCaQY02pebp/ZPAnnkFPbDbJxhs+L+AEObQILbSxFk2FXxXGuyXQDiR71
CkkPBlZyYOvukgy6++Q0CgFGUwcglFVlMemaSc/T9Zv2SM+sdX2C4v2qN255PODk
TUYvV/ypOfoH51ofONSRSXE0B91whFsTqE4bmZR/j9J71CngQPu0yFvYPj7mLPfG
9YirwdfOv09Tq5aXMYWDLPk9KicOVOe734sxs0rCnx9F7AA3NLA6c7qan9dz1gKY
K3nACvPGjv9yHGQOWgAr9tDu8oV9nVFRGKrOFGyk+KXlHTxAzQgRLQ8mZLVUeu9A
AYhSfbEW6btGp1vunYSAuhMMrNeg8ah0+O8VxLg5lRJB+EG0K/LizN6PzRkGsaWz
+nR6te8F9Kq+FgoAeW7JF+T40ud1eEgH67Xaxqp1RSSIKcTu4LA6aQo5mAUweV/L
o7q0Sm0lZgFwuX26wy7rRGq2Sa1XfH3y8rUu3/PvsKDtKClt4YiELvN15W+YJFVH
G7pZuQoI7ZOubAKXmc599D5nyqu7GbeKuo2AojlhIWhtl8+G7UdAiJx37EI+qJDw
UPZse0BIZb+gtpv7nZJOQt7Mw6/NJgare3Lv2/FzGywHqjdpDDUUUn6MLUYY3MTt
wRAMWLpDjOfkMIUD6AQwvaLq71nUrO+y+GZjqsJUjfZ/baDMg24YQK4XPfK8G5O5
+CwEB0Lksg2hgCPCUmiRnKGCKbJh8CbGBD3plaKmBvoZ1F9h9gEYYB6oacDsa/RW
yp7VVxc/kY/F/IS0qFv9zAiYCJzgg0t8cnGEGPFSCf85lqU9u3HCwVASx1lD/VWS
kKJ7HTdKv1Fjil79DTPBWzGhhbOceTKDnhqsBKe5I0vHHtpGfToX9eFA75ud2rf3
M5fpR0Tqkk8ipguZ/plk48UnSFy2AEzj4aFC9Jxulg6ZH1He9ePj61i5wsDVkgsC
yY2+ZK/liTrqM8kSH+NfbzfCzMVAxFsm05ttb1Igy9/58yCHtU2RnEYG2wGkeT06
2KL7bmq3TUPEleYXeIO5by0NhRAuIwN00CBEQxaMNZl8sRxfejpNbukj6C9+MrEn
hLvMplWw0MhMwxyxOM630H6E0vr2aI3y+oCw0kBoLiFIJDQqGIPUHii7UyQUnDna
p/H5lD0NZ1AV5zbLmziK/e1wgmOCZUaTAqoRGqY8FqHCLmq99XwaQbHLTpHB+NGr
7qGyLZ4HJ69AtG1sP/Y71wNE5mp48/wYyrt46UgXInqrY4HhRkw+ThiJHIYRlntL
L7oSiBQPZXKOUwEH9wAqHOo+U+B/k7cg3CtWlEigtEBagS6BavwFAV86KvYS5Vdv
RES6Q0qNgU8EZCpccMpjpSbmYpdLxUO0VFjNa0tE8+R9IyFhhErzP7URpmYavo1Y
EheJgft7a6g9GC1fNId1B9UDsYsjMvCLG/EPTJlJV3enjCRrj5Rq7TRGki/OQAWo
+9lYmDl/uz/H0tcM3EgOQYFk0yHI2G9fTaWp/iWRD0ZgIXDjmdNK8DKfXQchaiib
E76gWfOQZtZ6i5+WX7yarHcbAlhQTItYugY3vYyXiPXMVAbqZur2k/FNsN2e/XEI
0v3f9aLVlhGl0o31i81QAUg9DT52v5Fkifpd9jMfdlKERDO9hfEyK9gr69CqZbZk
G17/kJ2s0NbEwMYzyREpFBF16tqlkB3Vyrz20CUkTj9jwyU3OcUbw4KJLbNesyRW
VgR+rwG58zry698IJhtH8SVuQSATiTNORuAI8Sap/n5xgEPQNQfQ+CVOBT7+2Nk7
fyrqU2POtRlLOdby0+LPUIFWHG8ezV56zpcaKVjT3lHLqgNGipY8Jx04aCPjABys
9cuINFx9SQw9EIN4VKA2TsVEMdSHtSrX7t6qXk+KiXdVAbmtGfN5mvlphbgnlS5o
DQWx8DC6X7egThDl28NYuRO2TcAyhpyiMOCNih/chROpRTTlocX6MMAp4v9jbIhB
//lqLqKvhLzMGuQ4w9tUpJzF/bav/hpzcYl52i4QcBbR8ZLNfgS1n4lQBacfJajy
XyxxTf0Z9otL5TKban9BOaUhvXBGnwBEZT0Gy+1E3JY05z45nwdUUXJwG3sL/t89
+BggRTWZ5Z6qmLLxGthXwujZW8PAlQVmgLZ0W9XvQyHV+VYYPjC7cRlliDq7MZc4
Uy368tVGDU7izTtTPYgvRiuFQYpP6KG/oCMO1TVqEVE5UBIHAxkUyIYpYNsEHW5T
P/yyP3b4WKpFF3avyxapm4tzR9PE3+4OJkYlGkmWfJ0q3d1rhR4/pIoJfbMXTWIi
W8Pnh8nW11ciJK6NGUgm2EGQ8yqcz7kYInLGyYN+DzB4JZrWycHQoiFUvLF0h1pq
P5bqQ34hU/0Qk54XS8EzotQIbCnHaNFrtLlngpcYABog5imYrOwvj4C3WMtWnRte
BvmlLRZT8OETq7dAEKITMYBHqoU12TggJlT448NimtEZoY/DOtN4RAuN+YB5xjS4
Vf178fCbt+Vybtol6glw0O7EPYzk68MS/3Xd0aK/r9wwNyrxkGZnaHoog1WD++nQ
rZ+oiWLNU78nn4jLHKaCpkvDokSz/Sz4pA2WJYeEPbRXqrS5D7V5THLq9EWPD4tB
2Q9lsA7MH2nMBNgIADifqgDvvAANJNbDQpW024/mSPkjIAORoPgxlHVERNjSzgt6
xPVEr/9AYqYn6iyqoJjAhpeYTeC6Qverj8dAArRJWrq7sASlHgXs6J58nzZIwCzO
Uldb2ckbLgH4M5espDMfDLmrr+35f/SOfG4bBdN0suyTu/FMOBCCyC96zIF1Tls7
Fi4YwQJad3P34ZykrojLiWJush680NiW4fbK7YxDwsepHImdAXWyOmPr74MgECSs
dhkmLuC1ef/x+YfUzyNRxLdWUHofamdzqBcWu2MU0l8UqC90dz0OygnYbbhHsqrp
bJVg9gvCjUE0xP3IIP2py2auZrvPUPsTf5g7Q7+82AqykMQoboC9/eNiZKdBYu5c
fEWOP533HUsPfWRCe7kv8j8WydKlTYxaDzbu04XcVaoj+TodpvtYvbYEZ5hqfKOm
GrT+EVChy0BP8hyBxbwwym7wngNYRlytfgjJIIU7KhT6zoFh/2S/gsmWxwqUWhC/
pN32Q28a2PTgBLRviVj0v+R4sjLuFc7Ot8W7ZvUHpf9Ya2nEUfmKyRaCES2dyUgh
Poz5aODRfIAbaVgfRH1Ai1r0ndhM34tIqyV4KgbL5oMlsDTi64rov2Be1RExbr2Q
oOUGgY0E4YR58ZTruPflY/O6SdTeE5Jo+ILkTjJRr3x2Ns2idL/pKuZ7e0adzqDH
DlxZA3JlQ+lWbZTMTJRpsqfS4Ou5OYaQGp+IJUFAGgLEB9Be1SWspBjptdfyF1vj
VS8R9gSZf+BzqBZTzfwhkV1leF6LKrGkg7Ws4CxpMHyXHb0udg9wlekR0jZYM9x0
fFp7h6hgc26gISK+dbw5JZRQ6D+/cZeiw50I+/UB7GbcMTAgM2+QhoAEc9+1u+R1
q/8eoq3U4WS86grWoWdK5ThtvvjmtPF0qGev4NqlFkM/FWStdMLJ0lyxdHQS7JRi
QrH5V5q0JvxCG7WfLGapHhyoKO+pwVOzNeMupQ5+ZLsmFN4hEf7aGrwqvZjd7cxK
ngt2i0NFhwAFGCmMPqhemWXLxeKXoE60F31Yx874VcEJG5Ke0uIV2tKfioik8Qd2
IJND5W/35x0swwQHgGBxejqnUiNR14arvHRD86H4aTkd1Ozcs4MzlIucUaq3cOwC
eeyNr04I+h9/VZOeO43/VpmZtglZqNopdI3lLtiYLp/cvKQvG7H1Hpis6E0mEfOe
S0XLp5J8Ck0aFBujAhFsvKyJpdUxY3/VIqIK68Yv+bAzRDW5bQCZbGdLn7GbM8So
PiryKMsWhiisOu5gVfufkxeOSMhcatOeO2xvWBJRepEC0XJTSmhQq3VPkxgoI1Gl
WHFwGOS2uuiyj1TrVMmWIePtasxvM93wzcZxKd8R1IUMhz/XAiAY5uGW70gio7+0
FO/CWgGqAdhB1RfnMi30oInFrPYoZlmkSxqJKkVC2nGEsPu07AlwRqoxvxd6+lsd
1LXkaTFJq8QdfdjgHGpP8HQvcqGYwgE/Uo9pmZKX+TRa4jPMAEySxOIwFcHc8x9C
Juca0EifxvVMFX3ZBzUQ3dzd8Ag3Pn7qCZYGUkyPbmf7LrmN8/BRShuwx0v6lsgs
AXZmrHdYdBC4IWMNwudmNKj6LQJdIV043hqeIe/84sjDB72Sxx48M4Sp15iKsBcp
bnJifESOj0BbtTDHhK7wnOKstrh/pa9O5/RgHcN0js1w94ecfMx2EHfNGbWGLjKK
lYySyK4jWfKad7SRs+wwGOZ7Zcx37El7v8MZm0JAdLjQAN14PYQSGqzRDBAOav23
4MucRxbM/0pp8jqREB3nG6jBcdbXmlFB14Ck9c5Dz0MCwAKBjoy4aA1FlIJpS1X1
ISq5EMFVFc4XZyBWGygj/9mgUJQmel5LgxUgw3828dwSpwTfbsG1a4N/s9YgAjsc
oKSIalNMZDLgbDcQQrQU62EnubDc9lz2AqNr+rkt8V2UVZLG0Duu6ipL4x7Wl8k0
JEbzW/6piO8JpBRKJ8n6KSnrsLYrFGSZaMoDlf9JEnncbvxBva+SFLsDjqmSpRrC
c/UEFDjx/EchxXv5GjfTUdDMvC89EgPDuAZgos0Jn/fH5fgzxXieCrG0xQLOTwkO
W6kEZxXItlrbSBo7DKBLLZ4slArzizfF5qoJwy6G5kAWe883ySOcjfltEfbVi4Ad
++y9rkbEW2ECTgYQYUarpNIA25yYqRB26vqmm9P2d15kx2WLPT80+dG/UcylMq4L
c2p2xvHyjgeDJ+a98nZtROUbMrcdmT9xczu0i4YHfOR71VUMWbO3GawGR4ld2YvR
qpZ6tYBCd6cwe95+av97y6UfpPfWFjh6nsJ4U+IxZx0aDSunrxiL1412cjPo89lQ
0eagvknYR9dT+dLDoeScLY8HEut/QeiPq8xStSOz78i74SeKDxyeK0XH/Cswg26F
HdirYcrjH8cZFq4nPtY8KwdC131yB6i47+2GbQ6fSO+qaC+Ignh4eYBQ9o9UYhY7
bCvcdpEOAILhUVVNF4lsQN7PY94qkdIYl7q0xj22UaGvmqyRHIDNh2QT2ZH5mgdp
3NToZwmxAdpnmmzlwO7MdhMR0v3FkWx5pQpsGlMuS7WKQ38nYZTz3QL+jteJGNiw
U8Ud1WvhAYWp9hJu+96iv2wHbqUdD8EJBU5u21B/O9EzVlChP75oT9dPjgL1EDjZ
elzah44E/oIkUr+rYi4HKZFWEpsN96gZfd0V6gO1taigzmZjoded1j3OU2g8d52n
In4/UDkEg65G1r/vGxvejPF3g82Q3QhjRyT01124DrWovPiMJZschfMwaYnFfOby
sk3iwNbglXnzfvepT3MLRTgtx9UwemLDnZJOGQH3axMlywoT8tqFJqfEVi2Pyv8u
ex4FdRU5VVrdX068Y7wFBv9JrOGIuYgkz13Y6UE25GT0QIuKJAvq+usPWxv2/tFR
lZJKsRCebpQOdiN4DZfob7PYKzc9fsxkLzFlMBlZx3KX8uztXuYr9wWweA8yRv7T
ieJu7DCC4/2n8YyzZWaclGg+AINPvKUHwp0zOKmHYjGlm+UT0ItNg3k8eQSShGW6
VjhDv8U5dmSukc+Ru96i5Vqcqc/wUikHVs02Lp/vxa/UMR74152C9QjGALk6rU99
gM0nhYNozcBspFXkKoNoQdoG/wvimnab/lLMK9icUMhaUnPfIGJCIGVFo147au9Q
V2tq+jdRXyxaAb6JtzJcvbu8dEj5KmS1NSyDvSclW607DnQL0ZxS2ji0rxpgMf+i
gX1WacdGIprdy4RfFWEuUjY9ksz1fvmxfVyiEcJSZ2DU8C3RNyTqV4dtHtaR/mtH
jMwMw07XdhMwJzF+S92NfB/BDft5gA0SULsmshfLa5mODmFzibwuOMI0oCPU30CB
mSNLZIy1mMF0NHmG6s3igMt1QIBbl0JrU3P0v0jFHOKGCujRh3QENsdUB9V6Jhni
VnV9ATShcAu6Mzzo0ntNE5u394jV3nZHdItMP1OlOkZOD/3wtvEux5JhAZ6HCJQm
aJS4aAk06XM8HERnvSRpwhIaHJH408nnDIfqqyNyu23V1hJOVvi5RazPhAAdr48u
Nv5IJETeclPycmrjcWEPEJmGHIvz06y5545d0cuscCC2fT7RR6RognV+YyT6b62r
sFSwnvKbqzwxNkzE/a3jE7RoZF5nGPnls0gKzOteLXL+yfChEMShS8AXewVJS6Yj
I9FHKFO9IxR+1KR8955MvUhVrsyrXF06ryhXqofv5FqZXweL6ob/jTFzHvaKMUSD
YG9efB8MdwGUwwwc0DCO4D1RhR9u7quMTcX1vRm5HF9Hasg5Fn9DQYdRBFzl+TVv
84RZjw6SwSfED/6TkvUo+gb+banCLkG9iQaH8CVK6x/u8M1MMXhvAhG/MPQHB2Nh
VnYh27B7IDiYq/xa7C+t0Z2uOvs417r17OESpI6ubLUo22dKjOms3mGz/Ib94xTP
wPBaMe9CTwADLqIqxiFFSXQOWxc5YlRU0Pg5yPwitYmAndaHi3u11wiNLDYEd2Hm
pXBNHu1OUiv6+HC47Po8hFnnX0k76jqpKLn6tmGFjujoDMQJ6dD8OG9gcGDff2v2
fbdauPQyX0YUe7+2b4ndMMEMw+3sml2ladeNSOS/Fxk9eMNdc4Vw2Lu+CNwJDhaz
iZPQYLCAgAnSEhkSRzTOB/ZQ5LBVlyn1/pZjPGEWmrJQhrJVaupZIBku1YAiaXRj
dpO8xLZhJaRHKUO5ik6rMouQ6b0xMGP6xKXXLc/XzhzSWwBS4m/yNw374AdjpokK
JYHWjgpFpLuUy5mcBg8Bs0nb2i+tJz9bc3oRYy99IK5DGiuD762tG4ZcUHDWs7mL
+iDpAgmFgjAXbR4dVu9kh22K0/SrAn0GVwgXdbCZcj8TlDrfi3lw938Kp4P3Uiwv
ADQMXg3UAN0fZG1WvgwCilPWvQ0anzP7wBSg9VeonEpyf0LfsuN7oR1fJlDiO0Hh
wAbNPP2JlNtgSFrF9X+6ad1vhhGfG1GQw0RNJkrm6HROl27W6rN6BrVstYe85zuv
CVUdjyBgnlz8+Ac5wFCw6pW2oLtA1PaiiSElJX2dyP86oEMpogXXM0BVBxQdpqg8
TOfC+qqvYm50Mquvp7mSOqFxblqQifmQ8dKWJyEC0fpztWmOrwgvoI07EvhjQ6YM
ARjQXRG65eBS3WqHoi3I7V7m6WMQjudw/VThh2KuFUvxy3DG00CNyAtcH+mn8ecB
ZaIO3gZF9BvF1qFN33NP9fvbCa21rrpRIhgw+Udvpe8rQ2I8xus+E96RHe6pNYI4
iFZEfRGeIwPkznsAHsJvgMhIZbLLfU4RxZXj7g4oDx94TRdIIJTVKm2gZUIrLfkR
0GdMkxskefLY+LLZGQ2OSkfLDqhK6gpMtl7tEGmdcFNJpL9jL1Tsbfvrq+bjRl45
wS0HBtsGcBxYJAbY1fBRa00KrcAflwuTqb/Ol2WNXhPR87W/CEn+6Q3VLwmjB/0I
1GNQYJ3KBajdxHVVszCUsLWBhW6q1WO4fyPch+EA6VWLg6ot3KumRHar59G0s5Ag
uCeDfR5yiAFaWioTG7AfyUsD1Co4lSCjwm8lnS+fmMQbEuRWqDJGqQ9Wj9sir0+6
jurCaF7nS/NAKz+kfqO6QiOw7hqzFMPYFeZceUT3fAEfjx4tn4a/vumZCPg3pntj
UiCVUWYgH0K2X+OhUZp0T97Nli8PqD5iVoZVwv+Wq0Ew4qeoOmGIMAjx9bmqBxSu
m/nArBtv8JEKr9DLDfPZIf0uQQAMK/4Jh/+Fo2624adSB4LTkf2xGkLtSnLEm5kM
g+mn2wNkz1xqmEw4zM6AU8Hrp72xXwOiyiayo65H0BXzadbFsfnJ8Ty1QV2EkTt1
dNvuHg5es+UUb89yTOUG49yNGnM9lOI2t3KZc68Cecm7ewzbkvD2f6Bh8L3vsnl2
uoP8IdQzjNA53SVsX1T7If/7U4LUOsY++gPDpy9FAjpbj5bPJKz0KUVJ8lMD99u+
KICgKSL3bkQwxRgNG6m8/c7RQT2pB18IZHg2/Ch53D6dF3AJE0Ykk0ffCMY2KhSc
jNdzTMn4ISbBURfRZQo75c3DXL14K5cnj0e8SSe/I7D5hsDR45yViZCRrQ08v7VZ
tUdx7XQV0530VE+ZMZYy+Ppqc2aUL48bdzRQ8t4eF2enh79vuoru7uCy2suaWRJK
NWEr673cnuC+ijaC+QqPc3RVdmso4B+Qs+TJ1EnuypQ9v5V5Lnat0qcQijZ+U3oU
M1V0CkuTO6Hh1slJM8AtbZkTSbiyJXX4hTdNlLK0+pw2fXb48WSE/q6YU/x7Qw+q
m11Yv3FK5J8Et1KSYxxVX/aVDShlXsFPGeFryxhxm5t6JPgmZOrkzIQqiakCJwnN
6gRitm9sMduIYz0pfMEzwGZaqtr88M6Gio4EZXaRzG3xow1GVm35fUaym/D/szj/
FLuZRl90nfAfDbRs0O6ODwXHaGaxxakkf5Q03EJ4hxcPX62NhJmQw6LoTyytjHaU
trg42xLJRl6RvW1/AJfIDYZ+FSPe+gwjWe5xrOYYBQpdYu7Tf5DvKkTGHw/ILgE/
cxtKm4yqY219X6Cs0L1uKT4EFUGR2wSQH07DPw3mXgYmUyALcxIIYuQQ3di/P8my
nNWIzZgW76LgRoO8bk8+1Ls7J4E5O21PGdOj+y5JgJDY6hAuUrBivSQUl64xpNIC
rbNEXG/JKvkkeBIKJrPHQWfS4j3ULUvyzLXF7ZgVX/tZaoyzUUyrsa9NF0BXm6FJ
ZPKPY1S9B54b1X5WuS9QZvin0TYlaDLBbqq2pcNjtxCLCu7LUyq8ORbHJfxp9+b+
z/KMAB6GqYxbgrRHb2p1g4E6yGSQ41JO3XqhYppe2nog/qeQIRP3K+S2d/OMMzJh
xUvrYLPtGx9rQSrXNJUuoqLTsUNVxhHmcmp4Zev+cI6qg4eWwaBS+Sv2yqBoFvJT
vHvqaiW4hrBJNqeVrseDBVz/73U8juqhgkffk2EbUoDjnTEzy8OQTwwGuBzh/5Je
cnPNg/wqSULt7Em+9sHa2Akk+1XoPz5alsGJVSz548tiF4UEZUg+Ing5O3AQ1ZVM
eWVVEMm7swvHLQvl0OhhMhxzNUByb+RsmzbeC7+3x1JvMry3XTUjVFx4EqPiTuDc
gZ/sl8xkRX7crEz3vWhrfd2N0Q5V5XAd7wdEjCq2H7K//Gmf7xZfniR6ZrdhjWlR
r/aXjDa9etuLE0by6xEB5GFYZgCOcy0+rAl8JPe149MbWtSPhAmKCh84rjVctVRL
CBKNU6LX542yAt2Ww+FUXSTIkZcHFmwefsxfeL0L71k5xNuA8aB1uEPrBE8gqtfE
3Yy+Tzy1ZIPDszMSCytMYx2ceqdzt8CtybX3ibtJmFMGRCqMg2Fc3h3g1qWNSGm8
h0H9yK06nk6Y7KZw6qYYT/Y7qgebUKBS5CNHZ40GLzZR6l7fq3ciZXpRFhDybBGm
6KVZN7PN0ZlmT5EH8M+mzs1u6wDjMEuBaWGsLWy1qQYVN4K20gK5jOLbXmqjbcxw
z9fcJ//upgXXxBp7AdNeFxyA7subilRJGvo3rJKlWPktJI47B9m8VCVs8V4TEPDn
c8DFYjeJlTPF2yWf0EYaY6E+wQYDndeasFH9V3VIjUJttu5+q5wAtb9v2jDKXLxv
Ah6lt7uZiaTBHFFR1RT8V7XexcU6TdR6ioqAHz0mgvOwWRK19Xwm2yfg7DqpZJwf
jiMbhp/2WLpAH7xg9k/CEmUYlpddbSyabIPUnTKGZ+diJXrkr+W4I53+Zsp9dL5C
a6/esIegcNlb19r+uxpE18rQ+NJINkUUeeCWvF0eVFNH+4lYBficsRaFDbWVkGwf
U057zVrzDY77ccOe9+DtXekGjDyMeVQqYscPO0Khd28A3mCzhzsDKgSC/j2OFIXj
5gayQh2k8mZcIoQ8RjcskxlpsESuYIZZABX+1rZs2M9AKFpTaqjcX03ee/soAGd2
/Zjk9Jc6H3RegUFB3STEozbLJjwIjD5U/ebYiRdCVllylVWfW+gs4decoCJRF7pS
kcgWcGic8Txl0z9HSaz7jPzfxcIip/MMg4pv8lCmE/Xe6RhTM5DYlQc0F6fyF7In
NjKlmbGaSz2NMn7pOc3fLTXjIO8/V5cr3JzwHHEzQGroLwVEso0QCUk45JH/iFIc
sZJByyVEKmw4ZZM7fashEC3rhIt2T+4jxXLhjgWCMN0dnYvaFYAau43+Fstv36kI
mduqWi+KTVmOWDEor+5C5wHKnPa6C8dZkMChmTqsR0Hzi3uMSLNNTaqgxbyb0f3Q
2jddcvflEgjFPFIBD+nRib1l8M/LTPnPmboOvzEx4Su7rTydhp+9rQ/c+EVYfbxw
e4B/b4X2QlZEjC5fAJZmlikVj05xMOGreegNQplywGlCdQBbKkWChdFnT2Srm9ar
c4hhZE8QAgtrpImf3V+dU4PxAxp6wpMNpkIDxyc8yeCsTy/xLgOSINmdvmYXpSFg
6stpeFzUc8eXzxn+D9pAJZoCmPEIzDGmmWenB6vOUS4w3L+OInwDrXWXuPvqJHbT
+45FPYuD4qL+WOd3QfP02ot6E9JLUd8kTcmsMB7ppMu/f4g4lREBbkm6iZDYxB8V
3aOhXuUETk9EA9rW9KLzaSIeFkrFbJPwdXvqIBJErPR6jSCL8FQEXo6sCpPYXVn4
wtcExGUfeCjWU8ljCrzBIRVJfj0kfpGAhU5EH6B/UcvFa3Em0rKY9jy4DEsLQSgf
QmgloVhm8pvPfphsLWkqiFt9wqbuOPRhbWSKkAeXOhAE0xx2Du7FSRc+/CP2GNG9
mmi1xAeGsXt7Ep0/NLvZJaY/DH/7Yv8y7i6H2Vpo2Ekk0MAd9JIEEN1KB3BhzjaN
v0zBwW7ytv2ZpxxPEDruJQrz5kcOQMSVCwuTo6yA3+E939JEG3cErY3360wFIHeM
qPQCbwX9gfwdJBDaTjsyDPgtQ8H1k4yJoTWY8OzJp6uBbfLotJ0r7+42ZQZgPqYg
ssbMyBA+/C9HgmIepz+Gr5aok/jK2UA1m+fMM7ELDcR35G2yAlP3f+/m0nxYP0VP
9x7z36bIKDWtkDNQ8iJWEEo21P9wkejHTYZ3J0pYMgi3dRhrBQBcOqr1uCkz8f6d
FrysIgq38dxyAEWTikb8ZVXMUoBTje4YgwRiZG6Yiv+/VRxVaNvxcRMcKnyGNzi1
1Byj1POIFodZKCtU+yXAXiTTsSh38ZTcyhS/BxmEZxJtlwelIf4H7KseHVMcTttl
vSotoCUf8tXUvxwRUkK4fNOdGHLtqbVxQcXQrDn8S2Pt9waYarU9tOCy3aS9mxzY
o+nmNOgK/TAAHw8nxbGgVg07mK9/4k0Z0TqJscmdR1ppb1biqNWVBGrftyjo8Ikw
4hA0d3dQHmrRO06fR4b1myWhMY9LOXJodvPX34fv7Iy0O9wHmkrpeuhngzsOEDPr
X0Bf/B0GcmCHTDmgiURhOdxW+65N7mZMv015B6NCSGBspR2ZfAzRCjGjkBVap1q4
b0OyuyUFiSIJRce2HyPZ1fApuDtJCQ8D3GFHSH1/+Ua7G5AFC/vqF9phTW9lfT+L
Y4QlrNWj5MziyD+dm3SguXddeDsH3WGOyvfteUp4FJXLkvoTZP4kNlqjIgx5iwtD
lahKyr3gd7+VrZabDM0J7gVtUcxRiF+YSVV69KxQpPU429p39XTkP+WA5kPm1MXo
JYL1F8qxmSzatbgvLwv9hC6Jf6uEtnrdKSGBc/ivv6Zh7uKTfzs5gwd5SrgFMOFz
uIW8IyYDmJvA+IlOqKs9ap9Dst79xNNA9uaLu+PwBVJG1EQcMXSX/jMUFLZfeKEZ
zQQcSL5EB439ze15KDqRc4+htjJfG5gj5OHrHrzxmOcyotEm8K3k1ilBFp0wUFA2
txbN4amkhT7r+eqxtVcBJieuggSctrkzAsoqUyNZg3BP34ghKC01DnKcColLI62D
/cq+nbDCyPCbvMTRhyh2QijB/fG0a9wbMv8FJMTLeAe/4KnoFscbtYI6x+zfLFDT
ti7QZImgMWzvo4RTyNfx/8T1OoUdruB5YEkGMc1IP+uuTovldk5feskuh7Gxc5p4
RN/AKIpZeBE6hTuhv3tg3FM2dUZ51BNhSK7be66UBH2v2T20od3cEN+8m/GTK2Bt
Vqbc9wZ3SIjBp9vLaB3btk00Nh7MDanQzuWzQr1eT+COgGFcPdkFeiJ6fIU9zyPU
hyfHbEKHZ2nNN3mkMwUe9kEN7mYABoSDwoDlP3wWqFLdDKxqBKL27MUg4fQPDlLH
CYip/QYHrm4rWRQGRmto/zO4vMaoHItXo5pMZQ757/u2kpziUdllUDEyZriv3Ln+
/iOZJMNhm/OSHhZBreXpram48r5uKYPYBQlTEnkk8j1lrUh275oA2SioudVpNt9V
p1jXqgrjZWyJDBNInbueAL0h1tm1J/W3GegVzKQFhy5zgFCJz6qhKSECGWDQ08cp
0hDDfZBZc1b+Tb2NuUP6RQT8y94fJ2wFvSKZUc2t6a3mGiaqCViGVmptmtfkH66j
fPe1Bd/v4fkeJK+uVaG0l/dxcUa1xVlVIZfKikRIWTNVoy0feMwd8QgIIDrZ204S
flGHMvL1ptXkNM5HqBg+CdSwfhRGmkL7FRJUI9d75/7ElK04jvml/jnapFi09301
4DZRRb9w4Sr1Pbu/5vIKZDN5LbLDadg6K2Fdvlyaa/+tBHvtwyGrdjp2qfekt88r
gcX3AopxH/uSKtGUQxpgQgw0W3I+iviFfQdD9Atn2+oQ66LN/GQlitte90MRLs4N
cMLxQyWb76ig3+IpG5dq59/fx6MlMVV0O69e/oQJrxvfVdkA9FuhiNomUsz2Qu12
5fUwJ7D/j7QU9+hvIMgvZg+7ytHeb2MyM2FplRYbyUaN2er/vTzR61h/EE7oI8Cw
KzxHXbO+j3qwM1cgqYBGy/kdG+Eydfmua4oKp5oFb094JPN2/MSrycJv6YakKotc
PwbUk1nBm2AyHAyhiOG76xszI1JgUYmSSLiEug3sd5OrlsbhL2n8WBlni2kaltDK
eh5Dhj62qxJrL2JI42RkG/iFi666h/c7qov2aPLeYdtiYsGtN2gg/ygg84H7ooZf
JSuaWlImbDwMWQWgyH2U+zEK8KRp/T5PijhLK7HoAsxMBzg1uwuN8xK+OWedR+uO
e30fd0wVJ+hh2JD9b8SInlNlVegal91TXUPYBOd4wXDhBTejySzxXoz+e8PqLtdQ
vG1M8ynjj6OMPWhLJl8gMIcVdzvSb0F+oufYW8vDvMlVwn5JEW/McgIVlEP8cIUI
TdzljR6SMUdT6grx5/PisuBFEWsD8jckbvMf2mEetjFZOmhGnGgrNqMGbNT4UfVB
Y26+VRKTzAZx+haanOZYKZJLEJzSiYrQNZnctOksBGu7nrTSMJ6ChSMoChDXP4RO
nifQWsEpWHilPTqWw1SXyfTwJZSA3FLCSaT6rptJMi/OduINrnXuu3MLWrrX9xKu
vHMlFs0N5Chv1Mjwz6fPrAyj+bk/8zzSJqOydz/lqSrjz15SBxpoQQDJAPlvkGzS
soyFLsjjLUG428A5V8qFib+5UkYr4YOyleS75JeHzt8zpFwYnLg3tnzrQ4skSJpn
UXr35NnIuzUGC0/vbDt6KEUs+7P0tSHZdz3/LfIX0RCLEMlGDBR9tpUpsJpQkIvh
3TCmW6OHNnvPLBsviADzV4h+cg4LTLG0q2kNUkjlQ+WVbwUhBSCOtlOsccBjRPq5
auQZs9XEfGR7YQW1ntgCF3vvktsQzrAEcA2pSbq+mE6xUWATA+kMKqdcvLPAta6N
q0n2YtDuUpgEzq90YpzAlQ/ckn5IFM67Ij79BIiJ9xIecf1maJL/EDGBcfCfM4+3
EAzCcT6csP+WVdZbYcGSMJRSz264M9UmuMh2Eugao67gdSo15yReZMtACrjveRJQ
e+1xHyzHdJqsuvZSB93KS9MPm1KLpscllwVw9PfGllbDB52M5wwSA30O/Li07g/7
hZCBEAEU0I+DmmsCeY6CtMABYfCthbHhvv4+Fe2mZ/QCmx9a4qdPIR4O0bm3kL1N
nLWu4U+dK0Pw5lIAmU9qxVsD90QorvWsJdTdljLDXJVEZrSbddv9+riHn3c44fMo
Er50i/nfZhjkOEcnEQNdKFNyO9qbSQaHwpiUCohcWi5v2Tq3jICRS7RlaXBzI90V
l9xQDAE1PM8KpSk6EwGOiAfsvy32tZ98Gzm9GOQ7SjMPI6lGOOPRYHQP7a40UpKb
mR0FvxTAh+QovPTYnyMh0IwRVlwX1ugyqFEGGqNUyNgwINih5fC8Wx+UN3LYCxsT
X467JBIvachTxkexPo4sZaZHWFmuBQcWCsCz23uXTF3pK4gV1g2ZxSEMBWsRCeGA
pYcJ6r4P83cCDH8Y5CL2ZtvaUntG1UDdlSjg5iyc6XvMZ6ugqVSHGQB70daY1c4o
qxsb88QDib8lgiR0EPdZJt18BrwlhJFj8zO2Qjk7DB2O3opAqASb91zwF1do84NJ
/GXq5BGR5Z0fM05+7wj5Crx2iYL63A4lyb/2aleQKPp1ERACn5BMI3GanixBad4R
8C4Zh0Hzcdo5kadVsOAhdeS22+Rrmri/I/ZJZMpc1asgnw6KZ7MMLKU2sZWSlbb3
085BThS8mC1aZKn1k5Eltj2V1/5Wg3UUmeVgjVA0h2pOvYcIXdoZo8nL35EvaBQz
D28dA8rheQRmJc3O00HTq4ERi75FXt7Ra3ORVcNe4MWNNOlrO0el2RjPhksaJogj
z9Ie4g2gG+UJXGZrPyAXw221pGpf0LbCCaRoLhCJIokzJtPYCkNiDAyZG49WnVE1
sBcI8lGCoPKAHdsiiOqDWBspDAV6B/joLbwIviJ8WCFlxtUvkOGimm3sKkNImMa4
NcHT0hL9cYx1BcIZvuD7HuiMPy+Cw5c1N5B714m6xL+BxBAEGNFZZeVLg1CWgaYu
TEDr0U9qBQx+cr+hQTPKVQYJPpHRGANKPNu+YpyGIwaNgLTzuzvC2FFXWkJ1dh2l
9fGZDLEd6Lapti82EBsyAZpMbtNN+skWqCGThJ4yPQDZLuBKk3F12CxOX9Awtp0j
KTPs+K4SwKOIc5w01KSUuJldklHzbqmLH+PxxIsS+YixMyFZafuKJS1ESVZtww2r
DY8T/+692T13zMk8x6LoqpDfnENeLzOLwajsYykyl4BMP1qQJRBZhRbysBifPYQn
zdIo9dMN4OSAL7aL4Nt3iOXy2SADAp+FVYz7QHskG9u0s7jBOAamZNo4zV1oxq1k
C0ubR+nQygcKHTY0gi4q0dtcRSXxbDFQTwTBtzna9AOKSl8x59x8/rLbCj7Eny6Z
pfrx6nm/R8aRhuj1Nym1w5UDymXj9cJwhBSkKBxXeuvDsGcEUIsNP+aVwGXANaGM
WlVg+ZhKj/jFc6NVJFqUixMGRKxxqkeS2/LFe5GtlqvF6NiIvcHl1CZbbMnQznuA
PkANk6ORW/GAraCrmdGpMpjafyu8wagpFt7LVYMLwfLgbVsBOhWtZHDg203KpYDT
OjqPRCGePuQa0qQg6upr2owRQLdKX+3VLXHIfJcqQdSAnzeUX4PH6qgJLPbSizOt
09qhlEr6Uvwzj2KJ74FSLH35xEkRxDRfJ6O15399zGdCDy+taJr988HkHsSp6bFQ
YsIXZLEYK70CJ/Ivlh8TjqMbTkhXGjPS8fS84Ed6vhlWS4nn5c00kx2Qebgz/hMG
0gld8LX1zkK4PlZD2ks7M91rNYKsh3JjEX3YD8oYq7Wy44G6Rnbghuh7LyF33dix
ieNVX0BUmoZzXuZLen1GLKKUXBquRbzuZBbCAtvWZvMlJ3QirVx6dgMIvdpErLDT
WYnEx7N+ryz50tpFPxKv70R3eYlA7E4kpV23cyFSM3L1IJe5WqmXGfjgdCWu4Kqk
q0+s1Ybbtr9JwzvKJLGkAniHVuwMwyCvGHBq+BsPjvSFwiwD0AhEFOpI2AOr9ApP
9GqcmpoQGl9BULmW6CAS6t6zu55qQvkO8Z5uUpjPQIXnzC+y9Zo5k6UAr8SRuWcD
x3EYS631QHBTPy3GDelq13BvjoXillM+/RucoEGkWX0ON/9x+35S8kXmHjavaSrd
Q1Lr05392oNLONHZdsjLhXkykHTTj6gyI1N4PaW12iOz8pgBrB4XeKHkFlDmZDHM
1sLi0WQdmp3qvr4lS6aBSz+bUycUiN3AhVRLLgvsaB4Y+z1jF9h9/cMPojLfvfH2
8CdibwFd2F43u32Z9vrRfARx6HuqroNjveat/d5phWMp1IgkL9Q3FCqDHCGnchHH
i/8avlPu3LM9jZxwUnlw4kGwpTjaM05o7hZYrsNoSPSy4rpJ6F3Tx6jIIHNO82es
5XS/2MrPONPw6vnn7E7+RF+hPuxAKqfjw6lgctTP5ElQ+Omc2nCKQRgQfe6yu1wI
3ZYD1P77w3t/JNpTqom0eAcCmN11dYECuPIYP19xxRIBkbMtv9OPBLCUBF71952R
4ZhMWwBQmbTaViM+MicHDCWcPDgoZ1UGX0NcHFFGdxrPHIPKtMsPGRxozCMn4Ohu
OVq91MEyjC2VTAVBey7nuCZAlogmuCzFy7MA/9/tT0ZqMP78TEr+QrPTN92SFcqV
QwpwGB/d5T9mYT67lL67CmiCRNr7Ir5zYJptbzSwpDAbuNuB+6qVQ6WHahQzNwAr
ZMPmcO2QAdfWHhPqIcd4PfAXp3BwSca3lpgO3bZ2w0lMis/gAMVMidD/n8RV2Rkt
phWLwlq3vhf9/JCQCJPLsy6ZcuzRHaIrU2yN2XNrJz4gKlbtVdUGI8PMqBTq9d+T
2SmwYTo0aGX9E0UXxGdbl/E5KGqs3OT8xEjZDIjgaLJaD/03kGaqjYJYc4DBrCYe
KuNckTYBor1ySb2ahQ6V8TiAiPNRpvb3D07oRGC0vTrCNDaxi8VS9J7VZlDfl21T
koGj+answrn1joD3x3gW+RWRBoE8M1pIGrs2+1i3oG4kuiEJNi02pL1bD4EMwPm+
AfGg4OFg6qPiko7RRp3tOhur9uj4fTPddlvrbVVnveaxiXGn1z8TWWsqJlq9blVt
bGX03HzBJOJKYNHLpuvZeVBpGYkt2jibc7p8tGTSMg3xOn7B7k529Fxk069H11jQ
VObB0e3GkUyGdTg37Q0kbj2CyTM3GdzbBB62/Q6MauE3NbNKgZ+Hsc0ODdJNKhio
oPCQItzhss0lc9gp2Hr9AKEBAfEGRyQo3B91GAfoJeAx97QQst0hTbXEsV3YP8+W
QBWPtUQKesXGCThCB62WafRXipb3Dwci99z+27xPMG11MnLcUnaClzFPXTFJWWuB
jB/YOYIQrzsbE17NDT0Yh2fTeo7EkFV51fneL6tPjCTmw14xHSwnyWua0yw1FKu4
D0f2zugrjcplcKvF2iFoxnVN8qM7gvSgOsKBBpmjY5ym1HTXdT4D8jEibjmNobXb
i7EKfhF2NoPa+WAjm6Gbn+BFgUsMb8GFYfpYMl52ktlKDpFTovmFQp9IGtVr+gtq
eArcV8yq1kbHVAiQ+Fe+0m+xnxCLd4JFtfUrC/UQbqNszMd46JdQqsEfxND2umuc
Dx343LDqEYfTilTg3Qi90xllE6XT3aPSeea/ivxRguDZW3U4oo9CIkErPyDcW3b8
1ko7zoKGRHYgyrawAGMgWjUlXrw0HluWmoYd7UNOSp2FB8eDIKeAel82Zi5+/GMx
XIj/DhtqEGVE5PIWT0cg75dVXmtWRZJ5mUk8jgS/TYGDQ5pVR3E9z3vBYHIw1kMd
jBbQ2iA/oS/valWuST/rIQHuZ1a8O0WKKbjlx/pH2P3NTbrOua42GjmCpQHkeXA0
4Zn+4Wrxs7aZcd4391YrLZ7u6YwE2WH5sPXumIj4iJLes9Dj8qXx73amaCW/jg5+
DKvMjUoibPvaR9EQ1hKT4tfzqiBDE2jvvjPl0DpkMoIzSQuyPpJEVm4zVJEJsL/u
qvZF3Kes5swXh1W7OlTTQgydqKxNFoMTKDuifJISSnv8LJBV7BKWmsxrQZpxsjpC
gqY6NlOUu7Ss4eOP3wp06ZcHFgBAAsHP1BDLR9nEa2UvAsNXbtryoAgeypdtuq0H
+MIl0D7LTDXjBcusSJy769gIB4W5T3w2SODAbxvqGba4KcOwsOwdQMc0jZlCXJN+
fw4YBw0KLRcjRPOEBEQIxIDxIxigrI81mCAyH6L15mRsv3AgMytwCnaXK16v0l0Y
XeZnlvqJcVYmvltZYHIevG2zugRbuL5JR7U2qGDW6nakfUIC3/FvLBkQO4gxgi+U
Lzx9qCoAGPqvpp60ZvkxgA/SmhWjR0+b/E3n9gLI0XY9tOrMztLvctjDYTqvyd9u
GdwwM6/yHosE0Byugzum1sf172v5K8YfK37Sr507/fUZiLdfLXOYlR0ax3Xacqb/
OCOcD0SVjUfrSe6vseBEcnTOWHybvVNvoMgyA1SHUgKHgLsOVPy467KGeTR7kauw
z3h8uhMGPNacX3yW+KuhK+sR0mAQogD9waepgSnyf9/1gRn3efT9jtQEpSR3oUji
Ehy+tWe93oINoZI0GIZHsKLxx1xieVNR3Sua+SU26a6g3F9IlJLhJ1XgU0zp7u+P
6+XThEqSO3cNNqqy9dWp8xbopUKO2HCabc3sD1MpOrqJNh31LzoOuCOL1cenXA3i
UjnqFpL9PpkG0F1Orymmys2FUPQL0xB7xt+HZIXRkKha+kd0e370CMk6xtRDGiNv
tQ6GOwUv3FYHypl1SFx13ioobOyRz5V22XB+sKp5QepDBn01Oq5SauxoBq2b3DH+
LTThDJVEVeEYU8gZumLBXs1ZdIOdJJAZFqIcPbAb959AV4eoz3NHimVLCGuTZD6P
VroOOOpkrNw2ZNGzpHqsAxg+c+nhyvwVaECuWvO3nFaIBqaUz3gnyNKTz8XihiDS
csHRDadzJ5/AS/Z76ZUSLjqfXEIgvyQ8YwAZykF20QwqkHat82XDAJjvYkqqJtfn
fuBgbEvsjcTpj1rkd3hMhk7TNlpPxDCEDrxpFnDcZpE/LD2Pj9eLasxo9ZCLViul
NsEsnZzaVwpcKM9UQDZWK6hRbx3lcX8nhtNOSKimaaSUBtPphr5RGr4da5Pe2Ifl
MzNowDSvyJexjL3PnTBCwmJmcjBN9vQXNNs0WhI0li6webfUd4P70ovC/ZqDQTMt
VJdxn5fPvxD4H5maidotq6WB/mAqDzm8cSRQmYrg7zI4ukk4nAUGxvVd9f6uZDNF
uupegW9+l/4DCPevQOs3rwtOcUCToh7VLYzzEmDgqZrxa+jRcg7yazF/hlLzo6Mx
XwkKJiPkiQGgvBv2pbjrkFPpqwhtdAznUjVwmVXLpL8dub4g31ZSHaaQ497BDaJY
d1pUs3t/7Ri84/z1SU20aoegjGjnQhSZCIDwLrZpiO+laiMSnj2CRqyLpGIw5nPI
9GLFK5l3e/ARnPDceT/QHBzgpMfLz+xlU3GJeSf9Ox/os9KxkE+KKf3rXun7BUaW
xSJYbSTEh6Jijiibcxs4iXwI8sv/QPiuls/XSCFkHfRdHKoyi6bR7OiTKfEMtCdo
LbavnQtR6wpJA6ldMoVU4SQ70QG7x3nKUZ7ifGVhMTeZTtbu+IesPWlqpTbTXYHq
lVIL5dGSluoILDaa+EMEgKZ28lM+CqcsxcpC/jSzLhDqY5/BwgbyVGyllIQJWQ+w
0YYKd/VpoiQ04P+q45XFKtUVt8rP0/yTfK1hlrqlKYF+95i2vtMlAEXbbG0y0Cec
AHwlF4iV/dQ9A/3x3cDWBBxkfxObfmtMx6mJYSCscno/ZYz6NzqRavnIDm1tkVWo
JkwdW/t/vXLhr6EFgb+z0P5BiqU2FJVn1k7p6JH+jd91eQENXEVZ6mwiZ30os3zD
Sq0LIiY5WsF7HnASM7S5zuu3dNmCS0hOL4CKWCpOTZK82w20NPgf07EszBOgfniC
x78Jszozk6f7arEM/3doc923azFGutvlMY8BsOSFowOSQ/mg1/xgdnrgMisxkixu
oM0IJbhBwg6qZAagC0ym1LLguhHpVVDoPWMqTYBWKlwA9C2hMFq3m0AZtZ+YgU12
YVYtdEWf5JDx/FdMEp0flMlBhgWeIdnRd+An3nOVfTRWEkFV399gIbRk3L739myI
tuZ7wNP5BSxAqXz3LXoZ6HZBFhC77WxWTwGtGp3IfXN13AhK4midSimIXkALS2kI
k/s+T+JcNDgo9WFlSpc2qbc0s+RXBBXX94sFGkGoBB6bqJGkutpuOTiRcZ+ATQkB
un103f5bKljpcRsY3Zo6ed0yGinis7Pb7/TBl2YJhc+k7Szw7I5TXLcfAPoGfcPQ
Csmh/BaDRo/T0WUMUpiAHEaAjZI8Kj07PAq9QfsUL+OhdJ1Hbiys1cagktpryr+V
ZwjPxzKta0KZdxf+Q3RaG3GLa2yrM3MAOvCZJW84yW3I8Q+zT9pJsKKsf+LK7gHP
nQwqyX1h3vroFQHJKf39nHi3MoeqsT57SR6FeWjhTBX8ToFYEqN65kfYIsXu4S9l
t/vmlnWAKTJHy42S6DzxEZXvHxyAjZVhtwhZ+7xcjEFBzZcdiXlJfGB2dTB19ZRv
WBumjkMQph6KNLOSIRzGggQY11HgzqKUjdw0T+O5xqOX4zKX5rwUUtshTCx+nBQd
1xo5SzCF+OXggynRzD79KCP16SGzgH0DI7ePNMd+XXXie/xVi6A2bEkb94KkAkxK
nelDMwJPnBPpBOcSnX7JBKHK+qVoeIstHn8UbD3dJF6WoFuih1SEDIP3xx0qPPoI
I4FTWuYfVIO7CKFGPhKSmCkEkQFprqnS8cPNjYl3KC1vwZbdHVp0NjnNfysMHcwT
zOv5H6ah91QIOE3fNeJ03iTVqwgY6uaoKiUf1L+WCBVlxx6bpOxzmyV7wzH1Tt6X
8Ho5dFgsoFB49fozWjp6TgsDw5TDWAx5s86uJEWO2g1SgxFTN4ZTMpM7sh354wO4
bRuW2BUd37FlNexIMhG86I7uO5JBGs8WQ2xWiT60iHvAw11bBUJhvLZleL5EVBIX
KbWoQtO4T0HtBd8fL97kHg6uLaMJuEjo5q/FXPqA2p04hR1vhjQ45k4XexYdyMuA
NxbB5LNzlqDixNxHF82zB9GPMQHmMdxHFn0GZo/GGn9XHI42ZQudSOyegFpAUXyP
SVMHyRXHGJDbGBmR0wngcDB3/IsIjCR7jTwEG+t9xf5Az1BX9LGxR8CdlshIjxvP
+acbaEgCqEiYjPWRStliNATIOXTEWcfNXiJj2oXIRqWKgcF26gipZ1oVcDYzlUOz
y4puEHELDpbPmb7TwUlH0ISK8hbZKTV4B1PpXpDnd8zfzHzI84epThzyVuYYdpSr
/WyK0UvdxEoOO/qxTvKgFKntzMIK3vQsQi0SwI33vrZts29JxX0BzFqQDhOsIPmy
n4ivRKzf8YalNSxsQvFtghWWqsBPZ/ep/kE5O8+R6Vdwxm/SR0cLN9MwSxqHI8kA
3hR/li0bxxA9d6X0la8uO8VbU04Tz7Jq64Jk4dyMBg/icPgUuuYSZmSRevqrP+MT
/TiCvfn/EJCwYbMOfqqJyA04r/bpiWo4yiblvn4FPxHZ7VnutAWaB3bCwffz6i9Z
rp2+dpcqNthHRECedItDBtcXB/MzgFQTiJYPvGFl4Y7SDe4OPQYUe8sFhPDZbP3Q
rTU212UlEjp5dhruc5+SW4nxOTaWb2cDl9lx5K9vME4P8UHfwAtmQLIUCD5E6ETv
huJ16C2cL9NvdrilzwXcHCP68KBH6NPDmY7jz89QVjAW7/wRaKLOss8pSBNr3QKe
R3p55lzx0MiUB++0F237+VnRipL5An0hfxXwVdo7/+aMGcE53nMwX1o8+B214xNp
f9b874bSDCcfD8uhxlcjGMIoMoEnn2NFs//zkLpYOxORmWeuf3qKj1apgYpNA/CJ
gKDnTW6UyPfNPoIw33m8MHi/NWKQBcRY6jNuJBxTp5MUN6kwK9bHW7Uh2m7oqcxO
kEhDmHbg0vnvlmagNMuV7oPJJVsXm9o7Rve3gZTV1kx/fR1mTHreRQOQHEBCgdMw
YbKigwbiJlot5U4NVdkJ6jVVKpX1s9L1YqGkODAEzsgdJQqbJBFZEPER9CO3XKHQ
jy9302f5yqf+LWchhRYLBwHw4Vyuxhfr+VEckyH7KjWY3ptVEwxvI0IcdIfyv/Mf
FHQcnczwRYVrEoTuek9O4ezULU7duvMANoe4iLwzMQtJTwMtnrkuSYhbEStU+WXj
N705xML0oBWK9WhItr/K0q9Qfn0HRpvRLs9bIJMhvY11uikiEDPPIzRXNygS7ha/
9qRtfEx9i3oaTm7XeMd3RC9MxB/0gD62ZUr8z7Q+LuOKQ062EHXt+gvDZHqVsGmV
XCytkoi+K0rcY5iGm2meS8qCSgK7cmvx4WEAYK2roqMgeARBeLip+fzLkPkvcsS5
YeWcVz56f6pWgOmQGAeU6zoil0zLmfOl4nMj8h3WvIUH5M+/NAfL4eKVzzEf+2/B
o67OggWcZsMggNenkdxXUnkF63yK3LD+yFyVi+OwL/qtrZYNX9yZgLDIto2xxcVK
y8mDnRn/BicrxXWechwMRSbBYQE7gZB3MSp4WEcFi00t1TXIBBth2/pN6T45or7G
M4mDxrQhZdwhAvjmNFm/B0ClD8hCdDqvrGOufD6unm8kezk3ynW1WlhE/3XYu8JB
NzG7CHDSnlIrOMIxMXaNxWlye1gc3wTRUom3Wd/zG4qE6vMfaRsElLQoNOHwu406
mGFvhlNsIAYB/lAF8ekPm7BI1t25Qjv0BIdd2h7t5eiN0kxJmIjO5DnS5QGD486X
luR7L07Wsvi6P8+zNn9KG9vy1um2l3IIPdkLOECj7pQzYvgsdDTyKukwA++j+qEL
3c4cJ7oWj7rJY2tv6k9bajifaIC9NQzgUitYC4REw9nacE9/Y+WKX5/kTWRl9QJR
7YlwJsuhXBKzCB8maJJuTwual3hj9jfFs5PT7L0uHHKaEu/85o7sGQ6f6Pdqe18a
qyaqVJI6i8j9mX30c0aW//OWSADlGOBY/oLGOhIwLHiO/hRkC5jgK+zs8VzxSs/R
fMFqIHjWWr7dhhiUxWtA4XhR+t4a8XPV09Dpyrsmoaa49kgCDNqXh55YsTXAQu9e
maOJH0gho/XXxDJ5TqBz9fQIoz68Tw0z4OY1rn2d4OyVWkMSz1xTnvxcYKZneeAG
loS0e9UAKHGSKSX2c2ZVyob2IfKPHuVolZMrTRTdRUj3374UlCm2R0DJturQxx4y
OBTTjg6twx+OWrGluaB8IOkj6EKdoAIzijLKkxW5SIfRxk+o8rpWZCyPuB8IpQj7
wxRyE4dlugUqw7il0nswY9GFWVStIXjn88hKuLbQyW3mQ37vbAXNOier6B8cnIe5
n1cAGdSi9r1uhdfZ3C4nNGWz+bUT+SmcXiuA+v8XIz8hpvcuPyZ5Pal4zJ9kLMaR
yLzouTxUkJmXuALc0aKxHL+lY0KoFN63E9ErD45L26v+TWlR/321lBLJgzSAu1VC
st602B+tNMdMnjmhUb/a71RmosrkzcXUA9Rp5zm8POR0zgP35B21f7kBC2VA2ovT
Vf5wNPKvlfpTGBjnB9a4uzSwMGP0Naa6yWCBa5Mc4fdY60fQF4bAUOu7ASwYay6w
FQEkvB0WQvtG6Cx9qTL+JXKcYx8IWKvkTsPTt7SDXoa4wlUwJGw0rIFcj86HBkPi
fzEyXmCw1sYs7NnX+2mM4Ku4VIe6UNKSXtfWkP6zInTCmO77wm4SA3n/vVPAbvvP
FmIwbQIw4CRm5WoVt1+RJfbR1HdzXoPPJv3lsZwn/GaHExyQ567F/NN6GFjHM/p5
r+rWjMF6vRCIHmMU8Vl+SRFRkxG8UqyIgdqClxwsquUShu3/xyZyYb+b0Hg8CZYx
j1rd9Krq5Pl6tM62+JzJIn02YbYIIioZ2ptNXNu/hZ79Da3nxVDrOz2BuqD5c2p1
wNUmsvXJBhD9GEsOxEbfoVmxHmisM2lzhB5Pr9Rlj+fQDO1jo0myhaJxTWaSsm2d
PyaToujuOZar8uy4GoynN7hdW0xGlbZP3rKWiIH7eBU9FxHfUYgZqBzxqNq+/j54
Z54UKM74ml7hTt++HVp1zftsU9O710NP9wKpStsqbezwzS5GAUMg77FIedfbz5OC
ss6MaJEc6rzudc9LHSjosXKDJGEBePW2bPJRdezcrZWNrrH4TXiZc7gSiA0F8q8F
RcIXytvkI3JqgRK5DOfqrZ+31QbSadKyOMZVfFXl2VaK0aV766oZjQE/lOF9Eq1M
iskrIz4h4LcQqdoo/6m46/MI6v9lnMqPy6wUKVM+i9qMLCoWSItxysHcYWbp5AjI
x5Zbw+ktV1l1Fx5dJT2vFC/c0l4rS8T2y/S8JBitGcqWNilYdMNGsG9O1T01N3gc
2lsipj3CRlBHkf2VE/TsqH+B+rog4orcuNyfevVzrwhUUEdsWs65RfGsD61Wok0D
QpELEc/2oHqBeEvJ/z54l/JK5wyXQE0F9qNP5oMrXxSjK32nc11xz/XCCGLkA4L9
meXGZLSfFkt820LHh/+xoD5oo/klaK5XBPUM6xzXIJdqDWP5iwJKm0AzUsa3fBJI
8XikDtuy+yzsfn+cqQdo9X2/qDiw/dG4I5a9ibfM46k0+/olxUhFg8LVnEWBr7hb
ombZtx2wcks5VBt5ad6kHEjx0YfR0gGqkXUlU6i8644yOZCT9azUyxJ44idiejv/
hNQNUgeoBTx9EpVnPD0voj1TpbxHDwIVwVbydLFWYJenKezMOucEejnG66qgMVOi
6lqJbwfEjgvdMAJ+b+rUmfTw2kvooxxUFEQw0ld4Y5appqLmdtjxsduIPOTCl7we
U+MXQqI7ecXqgjmU3E/vsyrhpzo1S67c8OUggkkry933V9y1+HuglIWKSwSYnbA5
OtVt88vaIsS9+yfgIz7xtToF1aCW+H0/VHH2IZnH1HTLG4X523lT0iMh9FL82kH9
8hsMKyIF8p/qofL7ZD216nawgH8BXI78wLLLGto/3A8ClaCDS1oupttcNudL36eL
R8TViX8QeR6BC8Kc1G5fGyG/q3hv0qEw2a0SvXOqyezV5XwCiIpIO8QQafkF1v5c
kNyirb60IuYQUQyftF2G/Q9ImuW7kpJlimpiWtL/blyBXAxdBJSOIJezfkyQzUoF
AUP9HKLHkJnYdgagpUIvwCwt+5NcluVs2Th2kT/To1TcHypc4XWB4MF9qth7Ar9w
K9tzzM+j+EpH+XfottNM5DyzkAXKUjS+LkF0QsGQ/QPeiGwiAtAwR3+ZrRHSF5h5
nrrkRE8F974ZUtLMpsK3QiiAASEr04F7U+SCN5jbW9Soqap4Up+CsfCSZqAOv9SX
+uUmBC+ct2HfHUWAaoFUivGTjFOq4DrjXp1+z205yWuaywNqmruLeSH4U0pKa+5U
BndeffCVfXe2a32w8ZiARbMv43AKidNwF+VJNzxhFtrQ/EvsuSJB6OmdQ6UphKUF
1VX4jDgMGvc0S3GNBENpUHfAleIoSWrAdO5mD3PgtnmRdPpyD3VmMuI7csliOEpx
5O7XBXk6OhpG9bXAQbE55cqTbH9r8eonhbH0QTgNb23WC48H/j+ag4l/yIyRY0VZ
Cq81KAsRbEmE89LYoGSZSrRPY2pJxZf5iToK6wzXx7oqc4F1WaqoN5R3neznI0r1
fYHb30H6v+dTUxbOH5yz3B+okFp7dnbyrPJNKbmk94umARJ3UB8DAxytXkPwjC0u
JeUDsSlVYZo9fOsu2+BSUvUe40okU4Jr+7D41vDg5K6hiFt+0B163lVyVNtaqUOT
KSyKJnT7eDedsbIJ1dVzkPym3vtd4/jBBgs3AMOX9NbDDgjJytqWtgLjpBqYSJ8V
Hun9LARuiyPA3rYixH7OqGtqy8q5bY74KWmHIwLjOicZuOceVjyukR3H1DIkP6Uk
YSGiQNlzr6Zh0onf8f8iYr//gGJU3siXa97rqXQxYYf6nJevaGcVbu73/6NBYWvX
HlvAMzV1fVk8WiogUiq2Ro2w7daIIefnThoYKMBToc1nV0gVgqL9LV0J1sQpdMFd
hT7tdN8UZ+1uygzqYnGUoCjbt3i2MrgP6OHCZNkC5KlGeBWZJ504bhkNHb3XIidN
HuaS6A08cTKKBSFHh3uEwc+vlEFmoO3JNvU2rstLYh4urZnXB1cmFXiLtZGP8tuP
BOCHA/53SkwjB4IMfUAum+BZzSsGz1tlqsGUB/sVJht3caPyRn7loP4ZTo7apaEc
/K14d3heFAm6Yt0AVjBSNy2duRhy9EayenxfK7StrHo3UBWQhViy0Wes9oAqlSIi
RvZgVyoAsaHM++cDrx4ANI7sHXJjqd21WWcfB8A6RDv1xuRnDPF/2Asoe2YETKP4
iTRQi+lOQrH3pogTRyxAYz5bHzE/yDpthUGgNb85OKz8Bl21LCOE72Znk1VlAB/8
RvpOnjHYRkzgcBXJz67pHZ8YEV8z1iGi4/WLaRLrfJlBGTITSm9qq/O9MSrVTEGW
g5HKDH/ASirRlRJFE9Y0HEGHBd7+bB3IH+w0qXBl7YlQGPbQm1nm4KVvnmYNjmFs
U4aTmEbE/ykSYjkHALEMtJ3mg31hn2HvVTBC6+OI6wua5OTMwmetlcwD/r50xV0T
uMT0fpXT/oxxLjyfeslkmwCBt5BntJAbiiKfPZkCs9SQwYJFTqaN00cyJWpj2Q9F
MGttWVke6RAjCUZN4tf1mXTUXDDbn0eT2u45EaZtRItHif7N5VysZngsUVBuuPND
XCR2Qlbfqir3hqZkP3KdLvjzXFXL75NXBGEFfVA/W/byMNf7d0x4KR+9cdLQIt/Z
2IVw2gMLqDHiUoDHgYCcEXkxsevd3LhbkBfN5b27W/juP/3LuKt3CBBLCMEOz6yJ
V+8zYqwTV49XST4/KCV5jZM1S/1MzPMyIF/QtM83JzCc0clnxsUFa8bvOCzkP3DE
/Acx4yvlRwWxiCWQqa6mTGaV7ggAHhtRhO5ffpKEpKoK0RsRJhu0ZImCgWrQzKdb
Bpba7kM7neGS8IhaQ5UFC72EXAkT670tWB7sxSapfG9QGSGkOhy0q3sm4O0O6Ia6
1OtJACyCJzo1H918IxMOn4eIruwx9x+og4yWdXDS07h/o4LQ2w6qGpYpn0fuhcZu
nYGTTpJRmelV4/mFDUOwFxmXOtHSdWWnDKdIdaHpa6CvFFdfiALqZDjgFZYd6egs
yNNoCXfB/HptaIklDHwiJYur4ZiIejw8D0eRpxg+E8lo3Cc7apBkFu3IdYcgRNuF
y7wK9G3lTMV9mnkrFbl+1fp/zA1BE3MdBZW22B59DysA5VkM6LtEd4/4m/7DtiNa
spO36Abo0ttjIEW+dFiNZM5v++GYhVNtzjbqaZJC4AyAJPGT/OyFMSHEslNRObLw
Eee8G5tEpOac360tzzkywU+UGMbLn5+oYbTEYmJ6cE1U3cqLPdU675BzMMx2Km3C
5+tSaV1fKVIMKC2n96e3gmmf2xMqQVJZpCrIB1uTRSB0tEW9lkomeRPqEIgW1mdj
IcEDDVsGwIU3EFIiLpq5uzTNe9ALuQbX0QwSR5s7XJdu8IotG97MqI5VThi0EPMH
PoMD9xW/g5zEtu3ifPtmZ8E6/vYTmKwq0HfIJzSlUi88/0V++H3KV3oM73PTxfGi
yjDSL+uUXVZpI3lgCU1HMhUWHJLA02GhQV1a97ElLz1GfJFTAsb/tKyXp8Ua4zw/
HBv7RfTYYujtDG6M9euj8bZC7LtueA2vNGM3hMeN6KMD0LFD2MYOJ+XQ7aHVDT3J
DJoz/ajwFI/TJLdSMvtMrU0IgQlWMpZNWeIDctr/k5Vw9Ph4fnXQH4laWcPrcYkh
W1fhqV0aWNScbyhQQY0r/qalyVFXjsq/Na75h8Oi1JSTZsmF0/DzSqBEn55hgotT
Swf45PdKvBLYst4B2OORuSyt0lOM+r1rPChR0GGPC24Q8gOVq97DqLC+2M1iP2CE
0KO8ILPehwpHN6HUPrGPw9bemK3LSmcB3XRA8QplFII/MY4yWHG06k7w+6AP0L7J
wB1gAcAyLsWKkVD5HdBbx8+dCT+IuUeoBsbcHqcMtvEJNYE7YzBNnL483K0fTnr1
ljnWJk+Fgefjv5ryQ2KiLPbHt9qeVCBLdUry2mJ6kDpXOBilSsiwalLvEqgGz4Ee
gx01LAiuSUQf9pfHbqsFMicKeqUvQWQ/lu4DmTzmYmHM0hqoBFHYbVzw4rgYs4/2
3KNve10d7cpvHupzHOE3RrhbNsZO6ybtHOoWasVAD+0zYoRa3TTGmLyRN8HI+Edm
rskP9Ds6pEQpCw498pzwG40Hau+6NOcIiQ1GwPHmpNtrsseQTNHX6zPDA5D7BEnr
6SZ62kGx6Bqrarz+7zz2DS7IWjFe6iXyshCouzzKqXGDO2MS6A2cNW3i2WfevTs7
+6ka7hDSaWDbzlNe8I7L+sBaVTzF93HER9PypWT2V0+OtaMskRtd7OZT47FbY/cx
fWg/v6GCiTUCZ28SNlji961nPwtwYyYDEyRU/BaPZWzgI182KWWcYLksrJKTYaaG
To3MoCooreQYgw4GB9XF8NY9AJ6Dvr5WgGxCYGu+CCj23qfu22TxXc3JyHgQSLzn
gkBv21SY/SPC66rr6AXz7SUnSn6tX7sUdnNdLSokbEQEtkSAhr9HSmy1uZQJNtnk
goO3W5l0XBQF/ma2me60+Gx8CjQ5fmatKM44Y1z0+ehCxrxgHXepZDR/PCN8dYAM
eIJXvH7f7mTnjaEtNV/dAaqdUme9XmSGP1RRfl7LbDrqgNOyVbTu4SZv9o0o55nV
YwnG+h8aFRYipg+aL1SOaXMQUbtjuzbbX5d9h2q6NhWQz4z7DGO3SybM9cca2yWV
xCYkHKF7OvAavRLlmT7jJbgk4BI0DFDuFWaglnqtMOJscmxkl79O3TxYZW1w17xE
k1NkXlulaNlyaPZx/0h+ac7OZ+t3gdRfWuM7+qJS3f+GDw6jo5Yp5X+n3JnwHn5A
1TCAtmJmTz6AwZoQ6LKe5LSTgJ2HwPYkU2th6DRaktZfXbrAUYVG6akamh/3S8Il
ZyhbrRBUAW2XKZAeMElzuSrR/VwbU9s9YuqHvhUY1/8y9BdzxBog/ORcfCFRA+wx
EG4se19B1ZH3TmPokHAJeEoyJ2osJpYcg6E9U3B6KFt2Jbdxxc76M/XD/Tx1uQuV
SGAxWOgNQBO+3T5KYOzplADl4rAKP2jT38LqBPr4OWnudIx1jhzQRCjvq8xIndWk
bAMFbEcDTrKfhtqhaZvegEv7eqZ7ADVo7tGUHC/LZRSwgt7Tjz+uk7blXOe1TV0Y
ae8kqs4ehkwTj8OVhW93oGmqC7/mCbheCcoURDgn9VzxAKknXzsdV7T4S77OcKJi
ZzNXjeqcOqLE4ltJGWc2nK1AhlU1YkVxD85t3NlfQgO9XCta3kNLmq8Zo/PxTy05
Nwdj8gUDer0kCXk7a2AwLkvxruJyegiMuTHzSjOrjLwkPZ/54cOMqafbECrYTWEX
/EvmpEz9k0aEezXhY8KPfUvWsxqUgDlop3ck/G8jF/VyTooA+hZPy/uGCO1FaxEX
NaGQZSy3JmpvWBnzMw5YQtPqYYHuR0B5imZP8uQ4Bp6ZRrfWEdOYyyHGvZzsB0Zo
vXryLUC4LQthrwbReUD2QTwV3fGYaUfXW5dUqy/g4uVMaRep8x3ABkbgt9DT2l4K
VXhW3cdLbESgoszQo9e4Ds/ftjkBgUlRl/ssrfiEM++oqfSvEx5FyCn9DXYq3qBO
Z2YxPmtksLFm5ztydTv0tkIWA423KlZqndFktE04F1v31segRzhUxbt8Z/6YUsac
WsB5ipn+YTK9txCnAiFSuDOjzFgEuNgV/CokcuECPfutqdy1WlXUsBBs4RQ/6pFz
pexkEfGFzAEy6Ri76d33pfKMOBe0QOP3Jy9w27HqcTaFnPSw6kUmw633oJ3+jrBw
yle2HirnRBay15m38rO5kUuCkuXgDKsPk9lx/of1lji++/Iu6LPaWSEB5ni/Ud/Q
5D8CEpko75KC/TkFqtzA2CnavIlu2vRo51EAPr5lmFCG2a4/US97Xfi1Yy+TYDrY
/OFyln+crNRN+K4+ExvdvpKmIKCFdENIWpqxg0EcclRb2zvlAOaZVnwW6RNMZdsx
rVfIMcn+V148R1++ZhuKFoEozT7s74tJFcnWRwLumSMpcfGpnw4reofwtTK4ycma
2LuV5+LMqQzAxtD3H231AAH3wPrnQ934yTdZFscMNvYYHEUz4lV+i2ygCXPCArW/
ZJzUMWFRkbm8SdSakVXtTzHPOHG8VKEN7TSGChA5x7ikoZfM2lGegESjbBB47prN
qs0oKBoIPUWQOgBzkvOzMN2Hf6EF7FaML/QwHx12GVs6CcHy4cqF7RQR+F/JvAdA
AYbK18p4PsOEFC0jhFKY4J31OznMOJx+tgAp5ss4+qTIEXQ/p7W9Dd8zsr66AcTU
/dJAA38NuF7mrUVOtd6sDTb+iIwi6bnE5A2lB51Ltrj0MHpC2KB/DOy9oM8yMkOH
OIjp4hXYfiev+NOYUNM/CtdgnnK2w03OdF5Z4Z9aNkhz4W1NI/qUAhSbbUoVHvAh
aKI65ooQS01JaLBaKae3koxRM+jy71lWIMbMiySd0a0OR7pZMQwYTQfjjMprdwa1
xlU4nkuNMKiEyt82M1+ufWpDBoM9ZDBybi/d7kHDWsz6rwtJBwWsqnu4RV8Pehpg
IYBQALuYaQ6EOR6rK+1hi0MHm+ARAX1eSF5zlzIcjDlNCeC11Gz0ZyYDv0YzquEy
iIBnTYp5YQtHlOReI/EAFsJ8zojVyO3cYGViFevLil5x8DOMFi7FbmQuezbTflIM
Iddv/3gjA0Mf0rMv5Cf1g4ymVAKMW8ia5iFGlSaFKqmxRGFxA65dfdi7riCASg5H
Ulk3qiwai3oiSe/MWmMf+JScQscul9KmsRtycp2qutojUOqLVljH3tdoc83sRd95
gorewP5nP9tM3uqTq3ew0E5dUv7OECn5oBOqUZPislBfx6m3kLkgWouSsZXeKrkF
OEcgnPHVMaPAQzHuKWrGWLeCP2tV4KSQIbALw4V11TsdV46DcW4aCasuZrB+HO9p
UV2N0URaU0TQYRkkeIoCtLyJGgCggATW6vWAez5jk+FnoBnBIiokgT21JkPBQXcn
SjdypdtR9O2aK7doyZ5bfGJsyLZ9zAStWmSvw64P7k5pAAQeSA6yDBcrxLFKkjHq
vhgXYtQuXobBiT5gd+ca2gwoHkUywO0cRprO9XEQCiEM8HsrKunthz8m/VNLGjHj
o4KMbDowP1eQKRbh7STcm0Q0me5yUq4X49v8tdqGCEEbycnUjDacLj0v9KvHNlj7
baSaRQeP0hsZlc7TzDoKsKq1EVgxIUtdvC4N+qzRx2OZvuxwT309m++aCLLw9fAO
JlomuI1PV8+83WY9Vfi+74HC+e8/aEanSP/CsKgrVAafMdErQ03OK5kve2gBTOlq
esy8KIDRonXWp3X1BBmKREIIn/Gu4rh87l6FhLunocn66mmcoPuZbt6g+1SMn9kX
+MTPfqVL+DrR03AsSSPj2R4GhPOSOgItXvWxbdJ9hnM0DkjlGpyiZqjiLL7mlIaH
nzgXCkd/bi9q1+3qvAz453HNYnHXLK1O9KgTheOVvEPM9iYN7kzSxnDy1nZ3GX2J
r2O8VmunIhhh5R0hA0q2kZ+VbA7M7NfUEucoO4BB94SEc4khKUjcsktffd3TeRgo
W6CXN+rT4gGrMDZarzqU/I6UfJK8Ts9XlEpxB+9XFnSCARG3zmVktgMVCVWSncIs
ng8zYsVbwYH9RGRxKRqaFekCUvu/34nszHxHoUoybeN4Cxm26nPXvt/RWxRaeUiH
1rao6Gov1Y4FZAL/dKw1Ps1OV9OfMbllkg7UGfBL0AA0AF10WW6g/El7xcSbi/sw
Mt83Mz2oVO6kOiF2DLlWxxyGhFnzeO3dJ/e1NX9c9yFmbR9I5ia21OuDVPBL+AT8
NCstbov1KtBo80c/FiAIFS4Q9qr/ia1drEJ0r4E6ogNd+l8gAxROyW3iebjzcqxn
C4lN3sPFfd0j2QFgnX9vqp5hV0IcCYvjq/hu/qUtiDAElpdJc3M2TzJPTTTNKJVx
Xrf/nxwRxXM0XCRwxqgGLhDYwvyo2biQHN/kCtICi3ruB1VBR8lIUxem/QlFH5xe
/tGcfX2X6JFlzpfmQWGlc40Fz3eMt+8P5jgDoPpPzNSINr1ZRcRuN8Uk4z50RrYP
TTABZfHYFen7fkEcWjOClFC8qZav/bIfHKQmmQfHYGGhDVlG6vjAcEDD+r2j7wHC
dsgpcdagV+nlUB+9qa6Q471kBj3ESzg/2eNK+1IyduFGziri2SRsghbNQhpfFurp
LMPhKyCUH1970drbupZIKjO/kwXxV/o1zmHLneFfiDaZ8L2dMT9rVlCt8pMtXbRY
TFa4OVEl1cvf297AreaqTWUQ0iE4we2x/bAivjnhlfOnnvFUKXKs8lrdH9mgK93P
bfXXFeSHsllit04zzqp/3WN0hkqsDBV5ZSw8EVUBy3IOlCKvWIJdiHxcSMYF1YBI
WUU/SBJ+9sDl2AIi5FGaoGPDMXlIiGlkdacw53WBGwX+xP3pSftnCKxQIw2JAdCb
rELJ3NDHt3CNVvept4H8pQSfAi8vGAuBqVEUCdj02VSaWPcjm1bmdhnXK/N8S1tu
OwybBjqIzyyQp/2s9TO5y5qMCA4mCtUktOjWmoK65FHdIdW5nh0rKs/aE+jGaiSI
Ww8soemjyVPDzu5CdC4DAChkeIMDxjQGihVmZ4fOEq8GuASw6S7TELJE/k2yHjTD
GMAUlWcW66Ylv0bSXgejdpfjcrfrSeMR1Pknjs8BrcdRKEXdtI5/TfYxzVanllAl
hXQqNc+ThPVygmLBtY6nmXqIGCv8fz1HdcPdQfv+1Pricvuiysst4vuCQNM4NhJA
vLisICdhj7lfgGX7HRvpdXd9CA2e2zw4D/OjteJRMSITiZ4T3skNT8jgeFqMQnDn
EKjE/6cKG8EZ4pMnpZ3PXdH8ZNY+DHdOgjHDmUDgTrWKe+dMmB7cbA24GTM4q9is
UQIogza63fjrIGBzDfgpsyHK7gwnV/iUBnnVhwNfqZz1Vgq/EZqMRmlq/hUR5Nsz
dEY3blohAuAdQ1D8zhzHKOv6e5n3rEpqWw+FocYGITSQL7wQ7rgtUKfE6IZ9D6vQ
6xEzZK4oCeCbqZr32oV9xkZ5z3QjxMdDkkcWqpurrhk/31/pb8zt/XkI88ILhX8G
jkkCWlIyRJDh+yXcPw3g34us2bI0JPIjg6wpVzFigThliSlmPkDv7SsUK6JIhomX
fewKIwFopnhQFXWAxxzQ27ChzOKF1YeabW5yRqE+pmeeLQszEep27G7yQRuxVSLa
vEh8LzywV1R7IchD4b/gRccDmsRlpX9dTrWISRxCuB3KLurvNwgFq5KZH7Qx/B4P
V/nKKrAdtomEeP4pEGh1GFGg1/Xnhn50Yjcb1sRye7hcxxMfZpUxw7GYZK3SrSIN
gLwvyTJ3amFcvXUWbM+0crsvK3X57FSV80Czq4IPZWDOIXFBBKrrE8uocTj6op9I
dJpr8NC3/Y7S3lJbRG4+Ry3ZTYbhwrn1UdBXRc++D0H7NTplpE+iucEkvX1NuYxB
P/Hqy8HsKkSJRWJjWfJKKhd0WtnmwN9efbY/U1mFjc9DIxpFWrOoUKuZzs/3Ah/y
31cSR3FHQbasYq4hUicdk0nUm2lcH3U762YL6Nf4OSoF2ToBXY37/z9JIZ+1c+s2
2IxsLcKfunxt5gfzLht4Z8YpXqNh10XDAh3LM8GaQ7wVUzlID+nPP70bnh2pA7Mq
GfRaN3h2dLnQv3Tu/bk37QY2OoR6vmWpSDmTxGGHU1mJ4Wrvd7Oz9fHoCfbh6dLR
LDBIiEWsFXTY3UyP98aEbdkcTmiOzkCeXMB/UgdN1ZqbkJV1qfNSrOZSjVPSde1D
VGGivrTFmbnUBeoZct996DPtViS9tg2zU4XOqlFDnmYtbitSu9Q3XGArgHdb0V7H
RQBnonUaG9kdsWBBqVRMKnBuzY5gV/5r6r5jqQsoB4I2aJNK3Xie4X++ECuv3Ymk
hVnsEVmsnzKE7fVs8gKAQH7zRegfX0/aBkjK0DyTNWdTxkNeHvcJTf7VItTZn2/K
ApOb9SpQ6a3HDGPmC1CCmOCOMu8z/QO5fpVye7OY17l0p8MEe44oyiV13nkXZqLM
URQ6WlJPie8zZ5ZL++vwXokNQSuosVet4nuC7OKi3HpaHj60bqkF16SfjyvXJej2
Dk7uKFtvp9cE5kVyMh38i/PBq3cVa2o4HVSkU0qBUcP2aeLNHylEPBYX1ba69Tve
WL2qqaKxvZ9BQMchD/1lY+AGrZnafCZmoPICeGbeuY5t6XyLeQTLP53eipTfkkGa
iLvd/hUTSBV6zS5T3JewPX3yIUPv7Wg0NZ5gcIKx1/V3KzPBywMAOvr/v/PK2DoK
w4G7AYXczQrB1OjIQS18tNPCQCCwQcdhak/EFtsoZlv2qW6VbqIim+POU07wnl1o
fCT1TpC9DRExr0N3UASAiBfq6M3m6aaJ02yNI2XaKU/mGaW6wLlwEspSuu6kGyzR
lyaKpWlYRx5mSKYH31S1suhfcwj8wxq+74fUc+6othiQcxUz7RIgasYrbpjTfMX6
E2M3jX/Emhe3EZPFUvSUKrdwHI+v+QN6uuwFNXDcRuYLCGW70JN0nVJev1dGrQic
luEODjbD+I6skS7loR9t9zfzO9A2eYglTiE0KpFRdIN0NVGUIpnpJIuXtydLZfIm
V7kaZuTKOjFE/h6958WwGNZdWZkFUNUFJ3rwWhgZZc0YJXaF56FKU55za+JtupX0
OCnXhE/KT4Sglw8fF9t8tRCuhpMffk5KEtjKS2HUJhO/RlWRHzGAEIkubsAsZrFN
DlUJaunvf1LVeBN42IrxXL6y/nFLiKG3UU1wJQP1StvyOSjetpHXWVH+U2NSNq/E
PdUxbHsOO9r+t3Y1AiZvgDNu/oZuCjkZINOe6I+8i+U9SyRJyrFSkvdX83bmhr9u
TVfg1fmiLYkElVWOUz0P7VHE4GX1DAn1eBpgCWrqiFHK3IlUgln3Z0D3BVexark8
3pJhoVv2Itov0b7//n1I+ctwuW1VlHklQ2CzaIDY17254v2WzlW4Jcnf5+r1h2+o
EjsmzEBT2NVf5a2sveCv1/6zV0sJkfj864CRqaKaU+G8a89i4mMq538mw3+B/itC
Zt7ALg1PfWlTeSn+upCJSzuIM62LgdDsjFQ4BAnZTDn84JyqdMS0yQHK4mPC2g4G
uk2LG0Cuh1qk+uV4MTLCmKaHE9g48sn5aPlUhEQyc9es5oOi8Tos/BWj00+zbouC
MwRsZ7ilLA3L7wI0h6QTE8tsX07JzotJ2/N1gUmwf189WAjOPsDVRivyXkWu2WER
bqirvj7dzosD3PjOVl07ZCglmlrWWUiH152GebqAUVNL1LWoCPCW6nGJO/Ro2XHR
p+kmtAO5sjfADFxq7fL+N/4bqQ0QnBostrNmJP7SISiCpI9LtU1+bqKYjqh/4YK1
NzhFeaReakOJU4ZLDRC4aYYecZZ0aN5N5y0XboNrQ2ezwmhrfauqm6jWhVRYMNcQ
ZkmR+TK3beo0U4UZFf4u+2tfPCNE/h+GgeGNvFBaB7R9pYgMbex0EI/nkvdPInT6
QQO+rwDsL5dYtpgmFFW09kLHqpvQ4UsP1wfsJzdD9LGVGSbfD3UHEEdICjllV8pr
7nLdRX7nX39UA6HgoGNHOpPmhpB0RQGrkJa41zGHA8+r9U/On0t5R4XV+0yV/rNj
AXCw1UiX0hu9x1KPejvC0Tp0jJaQb1kuZEFQPhXiwlRIH2yTdvKXm53m0fmQUbfr
QPxRGs9hnt0Y+VeYF92Y4HoRPhSeUaQzpwer2PLURFcGhhW0MHrtIRD4py3wiXTG
+2EjhTSiyULkoR9cYV/4mXF5noWBggrKq+xi2FCRvFVR6hYqWcY5ClqWkOIZRQQP
RzMD2SXKgg38kifLclDT1suIz3ZS4mX6Y0Gy2eil2keIDznL+DNbNI5xhCQ1pt/D
Yf+iOhmLg1pIjfJG32xhW495QyRlFqAv71CwlfYGr9GSZYCH0K9nv59dSS9YI/pD
jr5JJpDr/AMAKo27Q6Lbz1mGMy82cX+6R1ANWJWz5TGxWI/IKX1sMUxddhI1E3rz
DhfAFR53ZF+kE1kZGkugZR4BCJbmBuxoXu+oBna9yMsZJkLx2gw5DN6LL2+TciMG
WR+0xl4/LNHOvx0GW+zSF240OB9vvBq/bp7+FHUr+KyLFSIz59PDJWIOxocKwenQ
vcgGDGy7Pf0j92yyFfHBzyQfbfETyGq+9O6pT0Y0td1w2O8VfvEVwqMFGfVa8HB+
gg94rxd4LGK5OP61N1hl35q6oNmYT4UY0W5pKANTSueq0/o9hVhW1AXxzdwvhoMP
IdWTtfg4XiyYqaYXgwFFfUwnHi1yetHSvUC8bC40lN1Ta+pE93AUsTTcbHb2t910
vURfwTs6kv/7oktohYWsMRNWQUOvw3DxW60sYLa606hzWG2yhcA6AIt71VY5J6Ur
b9bYBk22IUYCOH2jFWVd2sZFfuNuJaxPtF62PDzw15iVA6qWYOD6qXyDf7z+c8JP
eXknMru8k967zesBTdDI7+gVTWcLibR8z+9flS3Vd8459ldkBI26Ze6U5dil8nEG
d/hDgyjRoX+KNeQP3i4HcDQ4tb3GdOd9vAolFRldD7YxcIoBmYrsfwmcXHbJeE5s
36M/AnR2rhrWhqAJO2mW7TFnQkaVPA7GWsGr5Q96lGf1UUwRWjwQ0Oo9dB/sdm8M
VUnnm69ltMwCCyhUVyBD7t+mMM14pfRfDPiD7gQkW4YYE5+xI2oKL1oda5B8k0wf
k2XsRekwEU3v/EZJklS0pRHUHCNkMZ19uamekkwpFwld4vvmdvFZ2po4d0CkeiMw
aqORlV1AZsE2T8CKM/+IR/WntIoTxV4lUmTXYRIu1mFz87AU+VplGiTxwFnJOUgf
GpJ82VKU/ZdAUmzEFms4ZvwzVbNa9hVP/6RiBbJ+QCWcJHt/k8KzoIvAr+QKPYmD
D+3hi0PM0LBIRge4evQzFoRR9qUcdNqO8EZFpdLV84wSo15VOBqwLEBgmF6C500R
W+svkR78RlXJmfRmKgAv4+DWpjMAYefe4yvhdyWw2amr2ekg+ET8d3GHjAk+3JbO
RITqyCanViVLivKi6Dg9GH2zBCYRQx5B5gyiNr3IqYL19oycW7YYsaXJ0Yu4bY2d
Lgw2iZE9nqdyZHLO1nBZ+xvpAyKlMHR+PLy5FtbeNgmgZABE4/DhjdUf8n9zZSdf
VVYwe5H6qBE1TXcE+f2IUI62BeIHbZtUXv7pf4MH8Ut/IsmlHq4ZEHelLEwTVjPL
Bs7e9et9NyEhfNLFAhmr+ROosF54fpxuYGJOy/5ZzcaXUe96k/pRL8wY+mdCJ+1g
GgsRUc7klg5dlmS7YIQNLrBoUR+S3UKdyrGZNDkabGc26fzUjJJ2L9taQ/iAXl3V
HRaKlJ3JbUx02b/iNSeXg1rtdM46JzCEWld+Il/wHrs24rp0bgBpFPqdcy1hN0Nk
mUQcHdJfYt/9+5lZx5Yk4Zm2EaKkxkYEjEeVV7m9c45m4hhoflJnMymt6vO3izB0
+DFeaOCTQPG5CWdHRUsgTzkW+flyXPSjqpaAOPjHwtAE4gA/p27xGwBU7TYRz89F
QKu+QLDjko8ZSGDfh5BnU9I5IHkg7fq2OphbKJiJY+qdiZpyikDhJ0BsjFjK/+PI
UdWp4QAhV3UsOkOfvUAWPnrvkii5QxkPCIBleNHLaDUPzhovY8mKaZGBSgMDXrmH
teAE+6DuDaGxSPBghdxho9VBA2J0PVPzyiDnUbulKcSmOJP0Wd6iTRPVSCYk6M3h
8gJQJgtcQ/2HXVaoBhHyOHg8sRrTe3XzWZr9eazJa9GHphmkDveupUesyF4ggELP
FOaxrq7b327kaog2Mj+e0/B91y0H/Ld7rthpmkLvspyfxqXnqW/XsVEf87Eg914K
LhCvLvjzBzBE+WiNIWyqbEslXiWf9bAz/mc+vLWn/avbd+5SzKYdeYPbb3E2CJjX
mTLYjTGhmqV5Im5vEqipx/u9OHOfGLxvic/3axiPnruXLWT5p0FeQGlLAdMoWn6+
48LSiGP5wnLk7JCeT+8zWWdKsGJprEy4KGBv+BDd6wDJ7vkzCbxOuCDoXeReOU69
1jB7c4EQEGocHAo/hrhIEjoYVnV9UpyDIIHkhyrPu6UF3wAVEkKJKleAFTr4PNyE
vMQF2ntKu2F9VvES2WcnJwXsDEygDp/EgNAK84/wMZDX12JP8xzudiowL/s4nRd9
Cu+1E0f/wEyp3wS2PW6x+T9v/Nt0E+Eqkr6xFdYim3kYCf9KyQM+9Q0AY5K1KOf0
cVnGajMEIrzVM/1gsJqcIAxevtPtUDJfVPfoucNFdd3VxfNaI1dz/aBNC1Cqxr7T
KDDSTaPA3QfbkGRIxad/9e5UGpBg9tjfCz9YsWPVtRAApatADyN9e7eB8+1xtp8R
VX1SCpW4Boi+rg6nwbQiUDY7OIDXdbPCF2Qyoa6BM1YgCZ1/59fXLGqvPRoBwz6e
ckZxqBIcBxOPsE1ZT9oB2TkdyIgBUiOY+08hchEmTnbn0/qT46nagUziCXvfpjl7
PhJmbWJT+N3jMBMcd5Ek0liavl6kpToGMSFRb8fypHXwEbocBBrj8FGuCh6X2/+i
HfG+6P9XP7GZ8AM8eAiBVkkn8+MJyp5xDjFyu3o9VbDX6fDWuM4NAxCmTKlVg6Ll
GiqmIaSjwTa4GPNeA5sMyQbFWFThZWlgexVUfbfAIo/SaH9jp8sDVlJDy0MKJ5zi
CkcNAPvpF1aFoar5h6UFE8Ee6CNRuBNQTSuj+3+nzCrTsVZ1jiqkg4zR6uk1avrq
IrqY7sFGVeYEdHV3tyq6s3Ei0HTuIqsJsgi2OBvty3V+WZBOmhxeiQF0TRJvfRuN
x0bKG8xVVfJazylQUAoDWnYgUtIr75c/AAnzoPtta30wvlU7heKQuaSrcq3zGhkp
I2BMvbhLv1VeJOUnIFErKt2+8pjSbJgxqjTJK0zxWuKKnYc9oKijPQfuoefAa/mB
CXj5ma6+XfRqhi4qGJb7g82PdXegLUMYqAwd5HHnERDZMThdX4JKqB53Id7c25Mr
WWS09dwG1DrtDY9jcryMj31fPEli9eZVhgbdrSvNWIusAYaK4WxIUv5QhgVGrqcq
Kntxy/SfNNgbC/Gv9intYDGFBN3uWh8kgH262g0ToU6oVuMR40d45qlpNd6qS/x+
vYbYnYXJiF39/jD4CKUN8UcSBIaC/YLvsgddRO79aYI4RnqGXU6sbSvve1A/qNch
zgONLDqG7pS8iMcslBis6ayKaVHCblMX5KaPn8qG43l1Xl40NtQWK9Y51uzE5FDj
E8cSRvjH72ZLOvdEz3ftZI34TLaVK3eCCjcnNTRor9dTza24bRtuWnnz8BTsL3zb
Hy51sd2f25lsnAQVmpEzKp0oAzycLRJuandvPX8dHsj4xf0kiM6VgIZD/6ySMT1J
3s7w4kEdODYGKEdpURHdjB9OaD6vbvwHv9SuL6logwc409tR8ivE+R1lQ/IYaDku
aSThSts/dXlSSAlrPCHn5oJ+hduTfr77g4kofkZZfNjCHqaUTRyotSH7AQhcV1eK
WmEmIJpYK6inStDRvtxuGXZkxbxmVpYOffyG31PIQZfyivaANP5gng1SKWE7NAiB
PFoPYkttLYQTNiZI3zdtpNfYviCPaS6BrXMKCiJLWDjoksusxsnsYAUjMgPjQyw3
skgjt1780puvPRwrSJqNWeUnu3igiWO73I/EKJuqRufIplurLezVsiOn9tuaTR9U
VxXiFcEP9RqvN8MmcCadoKxI6tQ7Ix15mO4dn/yZpScTyLC03g0YRBr0o9RgBgsX
biXjwpQ7W2FCcNNvVmY/ytvzOYyRbcWaTdukazO/jg0xU6TwxMT/bNdMgLFuc/8W
HtT+f/kzzL6UV9KE0Wp2suISSXcjv1uJsJ/9OpEoQFELOxsV62sX8oE1fqtwFoAY
CIa3HN71UCR2maCHTqiWizKcTohQR8nIjTZkLh7aj/cYGiji2yqA0JWZEx112nEK
3xmsAYDVlF9risfOd22uc0mPj8RebwNnxy+gOC47QjjmVbwpGkxWmKq+/IxWiyMx
gbWbg/ebyvYpnlITVcx6wtvZjpunYRERyrvRy1h0wEIgyoPT+RfNj6y6qPE1Wu1z
UQrVoLU9LCElRi2F+vkm4hfga6I5q/OunCo1vSzM0+nfOn7C31MXTMuWEnPAyCx/
tQh16tIunK1HXSn/Hg3keAmtSAZ1qhLq1+ncRAM0kzjFllxbYNKMuBRkIIRMKsbE
feo1DqESiP9sH9h05LhH0di/lB3Ka4f2ZDQhaAEYEsLO4mvYCzuGUkmgFSbISrLM
EBuz2OhmsP2K3isf27zlSHl3EqoDF05zhpQBYRCrKDxgczIc5vHm799helpKryBv
jxIaSnjNhL1OdR3UGecA2fhy1dNKsSdZoloBzpbwySym+V54JNAFuySyUCeNHmTU
x6Hiq+F53n+4ZpPycvX89KvocJ/jcF0uc86M4gd0+5VZfzcFxb+hOSJLp2nnJUIG
RJ/UXDlzBVxjvk7UX1VwPOXds668xk1U88x0JougNMU+3MT/+r9Sddovbu90GH+y
2L7HVxYMUPTtxZeVSt62US2MPgY2MxGgsWJGS3ruOO0iYS2rvZKvzASPKaEm9aLq
VRT62XmyPbQk9tglsoOxTITtm7Awi4lp4QBCsERTZN4UD0AGXRjsmeqME1Qp7hch
nNnfT49+LfvDvajIaFN25SE+uNEneIbkGaL/ytbgGAP/js4ZNgFD/vT45uc2TQP4
/eaVx/nTPhDPuKiH6/l0YBpYRDBz4TKyQpwB5w16OjV7/e7vpKUXg5+P4GdZ9uk6
3j9A05JIzzlVx2AeHZCVF/tQ+cx/iIXoso/TulA0VTtfNKOujP+wo1MO/XiOmAoY
+oO9B5wkgFHbAH4nxeY8s0xSK9GMqknLc0b0mXB2ts8vjndGVvi4/W9eq1FTBlbY
xkXZgrZb3y7/zWJLtw+BFMb01tO1OTK86MwuK/gY0ESJkKB7BhTUJBIVb7fEpDsD
LfBK5HCAZBLZi93ApmaTpGnjFUWSo3wd+nTgbwBA3GLPnRa18IqvnVkU9h9VvQoQ
FyWnDJRKFwm1OvN+jiHZKKkFPbuP1VB64fJxk5Qj9bVDUOEytuCsgcrS7u2TKbZf
9QHZYk9DIL73Y9ItlIH0ICk2g7dBhFThylowC9vJFtvNxJ5wxh5IbWAWayfjcHyZ
BuAWKPHPnpl7Cp5DTPq6I0YGYEY68YhE6l6BkMoG7z4MZGgT26tyUnJvFKgoJsqt
5HxmVcGHAaUGNFf8PmTxv2H1kcSx462I9yoRNwKB2cnvqitLwB2v/2oOLUHH7kwy
06qK+Qo+P8DWLt6TJnvrGmly07S5NOONDv3gaF9PBa959VEgiteNpvLXR/TAbl0R
u8z1dOkvd2v/jUDfgdfHfY9sYWeBsk+dqra9OoV1E5YtIry4sNTxA5lhasy3zwAJ
KfiCjj1LNG/vkq0eG5dqWa0eZHxwsVl9Way0TL+Ar6/naBMbrZhFA6waxfw0H2b4
gFzP/HO+fa0XgkRXzqlXseiU7sUuAdTD0TpdTBuyKtmPAEM0UzEoVQ3JbQJa0sdx
q1tidvy4gkt7EebwBB5BVGhKdb1z5aH2pAwcp8C2mAg6TNqZ1PZRy6PQfTIh1Gnm
LnLBfHppGQy/4Qrt+jY7+OtsjZLterrppqDq+6PL5H1q+2UXGr/2X+O+x62MpWP6
Wz0PX/KJVocg/ZUSVfKD5R+bueA4gRpmV4GfdM4Uu1uRy7WeMjlHieifozzZR6Cv
1mcNh2dbrjGaRrsdIVrm5xBUXtS/WUxb/U89i3qG6ROu4Aft/WeSsjKnIREtH1Pf
/Yy9GVgXgA72cmd4DfiSerWpuGxZLqGt5e8wOiG7vflY3e12TzEtGjV6+j3eQ173
Lb4c2yTanRBYvtz8mdFHp8D2P+VFZsPRR5mZbNbNLtV5mk+PPhFMtHk86TkoRTno
E4DaTu0hAc5D6JnsLigHDtgUGWkR1TClIzwAJ/DXNuwfWHi66ydE7ZY/DMzcAgnO
z4dlD52NO1hVjmBFFFD2AtgiX2ymva3OizXXD9si4AYTUWTCFH94QiIj3n+Pvzm+
SYLXkoHOj2ihiRoX1UTIkLqirM9IRkeO5yxZFiVclE/PFQmcVUHkgFxoRoBxelDs
yh0Kk0czvYqWIJefXd/QjM4rcbUP71AMhCMMA9kbzGKuuXZM9Ec1df5TZGlzfrO+
DkPig9xx7JjO6lcJxRg2Ny+VKGRB2F7bNEFfQcgG9JF+XWO3miQtTzHFIJ5AEs/Y
obIMCOEzTNHSw1ppCXUCupbCZ6f7MdqjUTmyxUF3DGu/4xyiCFzFLW/0SEBO380X
xiAxE1nUNGLnM1/id+uk4JLaCe7yDa+zVt6kRYKlK//FfMdj9SM81lZs9aUolios
FWEbehqzPixPwtktnzG7ISJSRtYWmnQFVBfAk2GXD3+rtMae3LBOUrK271ocycsJ
VE+fZoUs1+Jb2Ho2klGJQA0W+tBX/0WOFwgE5a/YVyZgeEVxVkIekh8XEDV1sPr0
gC/wF1bFKXl4V5qJhv2PebtNF/H9E3S4d/JLBhVdvAsOToJUBqHTbrdyHVDk4Dbr
ADyFr9NKKTkEi5KFQ+pmpdZHUrsBYA0qZNnMMKempt/2e1KGS9qEXrnDpiQSi2zJ
1laP8nzwpav8/6r8Eoifd1UQMDL2B3R0+tQO7clZ44iEt5bw2xHRxtmit0EmhG6o
eK7uACNH2UB742h1bEedzK0AgLgooT8Wen3U1eZ75NTUrsJx+dMB9GEh+diPanob
7sIpgMNkFZ0mhsVtbANpOKtUCxMbKgSfx//a6jPFgWa9fvtHFQcKouEi+XMDnXCq
79QG0KvZyuAi3JqbiMlHKasSxbuJ9DOJbgZ2UN9nCUNBtQN0HSOMjo9VbS07TNpc
uxlimn968Z5RFvmw2euKhFyZ/0yBhXj1wqUACb40ukwHvaq70+A+WNa+CyCZuxPL
0ZLvf2szFF/ZdXRgxzA4CtII6WBD92vfFOl7b4o4j43/tkv53heT9VsQZJhzRZ/p
PmM9aa5KCkhs02tYBSEWYVYF1RDcNBeH/fVx6cKrQZAYF638K5EhjWmQFrSIyiDh
qi1XyH1Bq7n0PAakaDKuA4kfiAL+MaB5dMGK5ybhPinlQpORVQ7BSEsPT1tKMlmN
gjwfY6EgvcYkjN3HJczEiBvpPmbysY95/x1FCXTN4UkRRuruqrOdCL9dZH2iKhIP
IR9cZ0Acx9Agr/XyJ5+QKX+8nkPnrWd3Z6N2jfKLSk0hALNnCItH11EFVl7qMXJd
Kf7F8jvIV9x4TukiFZqjaiepe4PdLTB78xWnZHy7tq2fC9Vb5CgYU00iYTnV5Uf8
5Bu2fUCzwMmSJgyQqSDkZE8aKmgXuZ8e2dVyGuIVMhXwH9tshOgo/cuIUP9Px827
9o6Rwkx3y1PFHioYLp98KhxnNwUhdBMAjR38jDK9q9eKsWn6PzZUIhzWiXYY1t2s
XJS8Fzh0MzzWuxVBaOEg+NXE/QYml+Wqw/Tf3eB16Wd1dgZCyPlTVw0rGmDiLufr
oAwtN+q7TfW6UfYQ+hoHvj2IqB175mRG7lH4o2TZIifYpIQSilnD3KLozMlOtMrV
GP3kKXv3/f+hmirh43BfgCJHdoHsi5/poGErxaDr16F4Wh5TG4GLeGJFMG9Ugh6o
JMlVmF5ZHeULNe/pWX9I9iQYTY23qrXDyZixAhAeTdF0zW75AlSwQCuFpm6vJGSE
RI/ZAJEfqzIAdsr84Vi3cyomdCmxE7Msf3rGpTtkbE7Rb8aPvVSQLjuj3r7xvelA
i4B2joE9+jNmFOz62sOj7p0xJDlaoe5vrgcvoagMp8MmZATnDqfClFG5you8kGXd
AMCoE9KvKU9NNW+AdHTlbOjhMK+C1BpaQarU49FrJt4C9ETNLB8Q4FiPNHcBtFk3
/vYyMYvPUPUyJcv05Fzw8WLfG47+1bO9RypfLhhO91OD261NrkqpDQho8UZUfV/z
lBb9O+K+x0GIlIpKqperzhq5DkKj53vWiGxZovtavDALp5J8mxqwNlYZBrIVaM8r
0nAFS/gecU9MYkz0E/c1pAsh0P7Nc8sW1VRgTfF7ZvGnqI1wn+dDFrJF/57hpH2g
vvqfXAU8SLc02D41p7bn6XAZ+YWt6dzhpKZ+5pPHSbJd9gkJKIJOHL2g3JVSgYsK
91kUJci6p6P44I1ugtP+GcbrsM+PtVe5ajzl2c0xyqFcG8FY/mavw+Fi3hwRBv+8
ZGAZPhWoM4QtaBVV6SxgsADTliGmlMWrNB7AQrXj7tMImg6LvvCv6umlRoTdPkU9
nYwKkhOA0Cfrz4AsCLYwvlydEc/dzolELM2W7rxYlCm3Kf9MhLGYxEVBtxOvLuPk
TEBbYmFGnv7W949j+GCwQnZgHx0KbgqpVWKPRpM6ePCIglinMNY8If6P6Sh1UpeV
g9eE9vO7n2P5qLhu+1jElWGYtoulFpb8ctq6fj7leOU6DiOYRPI3daINNmdBqbB/
aOHdvpYTm7JZE2b7fHG2ztD8CrMjKWJ+rHmkrcY9T+MgNsAuN6GEN4ayNwKdNbcW
bSQ9TcPKrL/q4XCxvqhVokQtA1IbSIeqBgeycYy5mMmF38T0JqE62RbYr4kc0eDW
hw6L0r2ltrkeNk8s1PpkphD6KmKeYWYp5FIgFA/Fe8U3eio2L3l0igJqHXMXuRJz
GV2w+N/qv3Mm8m4aT59M+3Qxu2k309CB578sKZGajDAQcDeIEpgixnSPraqHgu9e
vT1jaVcDuz5CngLQuWXUE3qm1bHdsGDG6Tr1x7jJQLPGezwchQqpWNxdGZvutDux
Wq7L9fkbcexJ7XxrzStbOIBdZfVy9wMJKlgwxqwNBX9UfdhH+6kYslMyaNYkOBpG
ZNVCJ5MroJjGLwqocEecxRa3mS71pbwuegwToH2DIPL2By1Ti9F2OlE6nlz7/0Q5
qYzdFfT233o+eyTBB6zYMzDJqJ/RLXHn2UbwKXgM+7/U9Rzpox0nWlQjRshFMbgr
o3rG+vB8jG3GGZD4Y4gKD7V2d3bcDMPDOvr7RtRTuiakF6P94kQetLRPaKRHzQZn
9WH479aZKG32gJr2UvfmTwQTLkuP4YbmdOjpiMyh3H05NccRyTVQQmOAkwPVinRi
XBYYFcOiki5E5LaV1jw/ToSUOwXdfKC9BSddfDqkjag2wvsl+TaK7jzJYLsKv3Rf
sSy/G9g/eMuIfxaOazketUQ6N0oqI/+5ynWkt1/gHSEQNbUZyYQOS23SyT4VMmKZ
PMN/QnZNPPp+CZvVAm3SboFHppIY+IhiNo/J/zqFSPLYXDXXCrFRYIrG4JBu8sid
SzuR1DzVMVifQiAlUrsU+wo/we1rwRqB9WOA7mirp8wJwO3d40Iln10aCW2oCWuG
TnA8wFpK5Jbh+M8OKQwF1MjAbwp3FzTBkG1dmU46931ZKNisue/IaeyDkUqcZXHz
ggo/g7EDv3laCt3KZF7cl4HW8JRwSWjSwfiCkyFnb1EBR5ke9QF6N3a/7x5qgF4T
LHPbf/fy4pzyZt74uOLEL0ZwQ8aPNl562eny6brojmTSICW56oRBe5xKGOIVFp6p
hfMgAASm1Dwo+svBG7saAU0rvOHuImsVERATVhdeksIc24uLLKB3CS+pD/fU6lex
VJmn9d/KSGXOOalgJJbP7xbik08l9FOAJiw0395IIa48ZdeRIS1FhQUZ91cbSh+q
6GOr0GIluMHQGK06Pa98uRNB10Rf4L6CcsU4L/Hui9fl85ro0mCmoZ4DeXgwdXus
uSZYatwByKtQnKgko+FGU94cDZJWiLtqXPiKtK7FWU8WutQqN0BTmDGoYLzcIuz9
9q/tJ5pPg1YCjsiW+1bVvxiAJPsB+K2ML4P8tNcRmCQGiUNfz6tX8cLciiuYSt5p
KzpxJa/xVn7DMESeU++uwk0TCxrFEhIJ32KIFxt+LnbEADbNTTnYbSRmZciYABBu
T1+TQAhT/dqUm4aHgZniP74Gif4jJSCbELKWYSroJwLyJ+ASY/wHGZwwb19nDkT3
wfyOqIu9S+z0dG3fCFlxsp0Xo818+IA65iDO3Vq3aQO3fGj+E3bMrIiV47R3gmK+
Kqc3rU81XER/sHR41VB0yeHpBUH0UZ9Xzsq8BXG9euxg/zzXw5x+tvytVDyt+L9J
bmMBDyV0BgXUaWzwUI4AN193992dYIZdxDtZlgIt+uIPu1jhGfTMoZqxRQRxxHrd
vAwJZe6DfRMj6qXLp/goXqsRSD67vCckzew12FYphkezg2PEbkfkJw8yi2KfhdHK
zIKhsNvHg/rC3tGrqoMyhY4j02w/tsQ+VWjV014CBZ7XF/euOh5C24fDfWqceci2
9NZCrppEg7TkAB/FrvPvQK/kXia6rPXgskToYJS0hsNmN1THWO07TdsFiBFmV3f1
uJoL4GKxs+nU2BlIGJA2qupvmLuj4A7dMFLZKdOjemvSnbSiKuP8nEW9UYSIertu
wsyoulMhAAzZ79SWHd95VfkDIpcNFHEBI72aAgj7v9dTU3hUwdCbilcoOHWug1XU
S+GUljU52DrF4dWG84vedvEWbgjbtZ4Gp0GqGwexy8JbJOsjKkmhctMismuesbVE
aqoCpK/PtZyS+XB0ZSxzUkJ9tldCdgful9BYhmTuKfBfVCeHAVIgoVfqWWWeh9xa
4IPHq34N+dDgiQ4cosIx/Cyte+9HT1F44KQKFNdOOwa70w1jZRueZRTwXbXrb1lj
prTlCyC/p2nsYAAy2ovpuUxbXDVLSSK7Ql5ep8BELQtYDPegpptfMLRrD2g+plUs
QpjsndRnqEqTkWm7B1LngqvtHxcSW3NxYL4wYW6GL4V9G21KoDgAKPUBeRScLWfR
wE4GnWLBRUa9mGsQbx5tx93zcIfaVg0SdYV/54nxoQYzA+2Zbtl4NLmMC7//zV93
UMb7LwYHdqaYggPhlQOLuyNtG4p2ibqyu7MP4lBCRa4YHeb5FZbDY1l/536wtXds
BMwfnzcN8xko+DCEY+Z7jLog0rFJnrCEYFN5NBhkPNl+fiKGvrpdC+gysAq52MT4
nD5iyKXD6yNiumr3OS8IBtwXtXvHBys8DO76x/ZoImidp0OVhsYQgZBngJFe1XIi
PEBIZs6oRgwkiRVLIqmv2JKwpn0NlvgMrZseFSe7w0zOb/pu7kZHHDeaBcq+2vXB
8olw1BRwE36qh3Br+Yh8RzFhJHc+YQFcokYyQ1MwB8YOcNxcl1BgWvfC88D0scL0
ArhjdgsDtaYO4Q9HzPoTYvE8rfayhmNNESPkuseNe+9kWtyeCU14KepcWYeBSMLi
Vt8vO5NzCDYSXo687gdMiC8v5Gj/lQUq2URhM5mAUCY4fb2FMHtjK1SzSbNT71Os
p3VGOMRewkrfVwbxBwPp1GBNsMZERS/Kfq7IkVyq+IGmkzMb3vZtomSMYlusRdIE
tv4FeHs+vx00iNn6WR+CLCBmSKnatcE/YL4HD7wUa07bBKqyzSt7lguxTGU/fPQg
qf8gVtsjWMfLzV1wALkHqjBVL3N3yfYe5sg71hdrM+bK3ApfrJrfe2/xbjczNbTO
Y6yI/zTj/cyewuic65EJ0LcmA7ggeOeOTM0EeL4AT3fZwVzsUoopBdglkb14JKBn
QxKtt1aZkfP6e+hkPDXOQOA+79FndYbP/6AF/ezIGQ2aMUJft5Ku8SlYjojMs2iV
llfiF5rCGy/tVB4wA7L7332OmqPwNfyUO3yRl6Qhqhr8SSfYgPXIX2tVWivmo4Hg
6mZt3wFA6bm4oYr2+bjuTbTpzO2zc+bDpUWNL0Nzpn+y6+MWwdLwOeguuHHIh77Z
09dPyZMJRihIOG17VqROlrMvFofHJV95uVqO6aiX2OHSZ2sFdZfDVG7ieY8XgckM
G6kawyQgXJxmVb8ba1IpagENUWomhpzo3Y2tsB9l5J1vb0/hwnFqaYTXNKxL/6nn
GkhMXq6RXDKYFA6YBP+JSugmwGbaiCGyAlXAABhdwqFS+aTENJWKvcTAwo61zJvj
aQQzZHCiLEzaUTuy+rLcy+hsO4wtJ1xLvESC8dLRifH3/r+YiVXuBwLf4fud2m4I
5FqfgOfhOzkK/hsbJov7s8N4fbKAVlMounvq0+Vh4GzB2HxgNxfFwpNTDr90zh2H
ejmVHN3BiBL7SK4CsOYk4/MO2d/sBCaV7DcK1UHOWWjE1OfdSi+u2pN5cXn1/Rpn
iKRNsHcgeAQTu/zWgEOPMbvYsy7LA+Idht7qHDG49/TPxHHNhYwT7eHIKquVbE8j
t0bLhLBvh6rBNrmpBlh+XSLWUCFz0gNsX4MHgslP/WSaC6wMx1FJH8vl+ct0Lf+f
u9fyC1Wn6eaUnfUi4FU/cJYtl4nHnVUSdo87OeTGozc/WIHuVneGawI0+XtUXtEl
tlJZY64cIabI5nIrKnY7wiQixAPcSwkvGWyaSsWsxN7SV8NdxmDtnVUg7tD27BUu
toBt/tqushk7Re2isaUF2TSh5tP8E3TYko8OpuTn4Gl6SOeZr7BtXSulNmgxAHJU
1zY2gNUD4S3q6uzOsbohgVn4TR+1iMbm4+DYXI5amQnEWr58e1Nofa71N5ISEP+d
Z9N+rpWivkBxveBtSr9KB6yxv8MDZNmDw/BNg9s6jezwTGA8hFfXrXnrWmdBbf+X
C9p6riXEpNclDNWAH3qGJD7X+lP7qr2SB4O+9C8/pRln1Ot/z7fmakGIk7VGWksM
/bL5ZmEEGa+JwFuRHliVXlhxQBr24OR6E4GStfzwpG4UapYh5x4iFN1yRBNt1wTP
lVg3pCWo1fvUkGlaoD6wluMhIb5n+iLML9s30KoK7SOI9vNiDpO9yxqNc4kEyUq6
SnRM01WzgchPaK9KDY9H6stJcX+Jf3sGN0Ln4Wv86s5nPKMobewAV9vNW5rkcIZV
pvEJJQskPuDfUHnimAHa7RsMfBmbhzwtcCrYVO8HWaLz4893Bg2OaO8JOO1PV7Eu
C7LGRR1u/Lx0cNS1PvyMKcH+wOpel99KM4pMUwvs0pFRq5NDj6/m2m65IhL8Heh/
lReZei9wrWhPz5hoeohpM7e6t3/nPtYQ0nLQRu8hMbbpcnw6zNSEVy6SIeC5K/Ga
kuTO/gr1ujAbOPzK/faJJ0RxU1qelxEBgiCs5CgPGd2pq+aqC3123UUUT5H+7GdS
P7BjuB72BYm6VlMMBVZ53wMwMlZz1XKp05ayXo0aqzNLR88dLZzyCOTelVXP3upJ
BI0UlbQ26pas+yz7PGnQsqn7VhluKURBWQaYZQnITeULR078hmL+iPx9xXqtNsqX
s9o/TYnYLUDkd6vfYnH5GNysHlANEgqyBHcOFkbpKnF5edF75M0TAEPewUxqi3SK
1wqsnObbjYdLLNd2EGJaQNsyLEQIaI3NXYcIV7lXICJ4xcOP5Mt5vgK2efg/oRnm
D4zBfh32sQPXvO0ekpWm3LAvOEpW+9BQlCvkAQ5nBa/qsm2+9XxJw7bqp9opdN/I
hoL6FoXtkRUpxFgeHqlCtT1ZtoXMP9GBLr1KDjKxZKjMLiqAR/rJw18K1YdrAI9u
1TrAIoxMilq4UZlFZ2EqK39GorAd1AdTCcDNsJxPV+wx4iz/ELmdF/ErODYWyFzB
q5/UOmFOke6nUSStDT7iDiOOq6Fhc+DGkcEeFGtPLhfN3J/ZxtGKa1wcafzGUPBH
WBq3g/oEegrXrYzDJ9StzXNq/RkW7LaVqvnAkd1a860itRnlUfODmV3KCR03p6qY
t+6Z9cYd8PE5fYA0g1MjVf3dQQdRIEzPqtUkbLYikMl4v7dvTtBNSgRsHYc6plub
DrrIqCJpIqxPt44jbCSX9JxebQk1LqvOwGmIIRG1RbVrr0/bXNnLQW1UIckDcBcY
7qfk6XVmLZPyFbJ5PyA2YdhgmEs/c5C8i0s36Q/rxP2qFpdwojGzZz4rZnYDpK+O
hRmUrwK/4lZXsqj8rcKFuIvAK5HoQr1iAk+TKBN+4PwBGJrri9sUiU4QTNA4jota
fNs0Eb8LTTgnUMKEV0/tecKoGUrOw4rqqPVGo2GqQj5lkBJ/xUyjbBYVMVSjKSeI
Vdttb7kYgJPDUjT3koNvA37Sn27g0/ArU2NFMd2QrvU3gcl5N0LK3RQJ36fB/zyT
b5M1ceMOUdtVSFcN+kohI5JpGCmoet4ZGEdVJ0Y003fA2ct1pG4On7mUj2C9NMev
H/QoCxILUtw6u3Upss8VuNxny8DsWWMoDoKsB/t6GNVNz4HjmYrx9uvEJXn4ieSh
cQO1Mc92xUpQznLT7XWCQ35B+AOliHI1ZrPqjPef9seP6V/VOTxut39jyKx12uFD
kAn6gewooRXaCoyR2ya0PD41ABAjbmi6hGgfpi8Tulw+Ye6GcS5Vzu57yjU1ZwVb
5j/TB/ubu7N4MuTcYXfsZs1qAJqGptBqtanGpEl8vRal+NpVIeS5V6V0iZP2RzEG
RiiLysr34IKUqAsDj/ni83RYAxXHRMp3XUpQhA2JM3bXkQrPfXChV9xI1bRV50hl
3evlQIinY2jmF+6PWgZ2uRRAWP0joOfWN9uoez/atoaCwD2QAYWoT7h5rK6uk0cK
aT4k5ikYsGOf/s6L8RWS151jFtBIH+T0bnymX6PBlqr2+4WLz6NzuvK+wKgWNBTW
LGQDuIwDWz1U3jRHQQVLzUX3xBuj2/m2BC9q9GkUMDTgscD0THoxxmUYt7uatQpk
KJNkIpjAAX8EblBPkmOLQhDUiuMoAnKTWN7bAyvtMUgNJh0fRB1aiYhNzVMwkiCG
jhpf9SapVmEvwfFTAaSHkbu8EGJ+ytLViiAVd70pu3HDjFkcIlKhsciFJwu6PX6X
DWA3SRxqWpR4sPR9DU4iUyYY/BZnAI0+OzDQ194sCA2DGcMZJUPr7s6IAvk37W/D
w/u4jD5sWL7isdUXFtqkteuDjIqCHRiKKG0V2NZ82eRnNyzDMjRto1HNfjH0m3yJ
5pE6n6Ulk37hzWWJDCmSFtSs9w3X/OWm6JpRrIf3EWAI3oD5AlQtu/KGvANRjD5F
Eg1zN0lV5YxCPbWySwfJ3impTKCB4JZKmVBK6/CSUmthRyt+YAxO6zx4lTuGYEV/
TIlOTRuZZPmWTHm6kSTxq6il2nDKnbLET86aFlEuEJP6RCUUIEV4oe5PyDQGDJZp
SzVv055TCnalO/Tto26qM4glCDn8dDHhpcXc8IdvSYaXyU15miMl2oiqPNYu3xlK
yQV4/pPiIyatrWX2coBC5rZMNa6Vbda1XcYC/v7XKyfYGH4wyBFHAQJgeQPlyqZy
gsucKb1x5nowPOqTcmEuEzKcCOGbcDM3JAeGzk4ObjZLaaCvNsYZKsKV0IhVRBwf
TT9adsBNf8FUCvZMdOyfBCl2ItlCbFuS2hlghZDzPkuPJA1zbJN9CLq7yB+fmLN5
1Ta5wqj+DoEdrFsc/P/aIbgYjgAvdU8v08Dk9L0qyyH2Kx/TbhfaLXa8SGSjJtGp
+/ANQxF6n2vBzGT87GEq5ndCHsZUfZwmoey2EgZOqhNM/x1Bmn1f+f5WGurEpzuH
DPa6YyKvFt7c6tLTMO+6evmtMrHlvihDsc3xc79+NVz0WWW6O/mme9elqDCebBy1
oD+8O8Iv6fNT6zeuHmoG5z0mPqaynd6+IRZGhLfdpmoEhYbhhX4tAXoy6egocUSW
buK8pzxpdjSLmqDwbY7obIE6oJQ3z6qU1r/18+mlgvpYpb7tPHvstkM82lZa+dfO
JuNiInWCxWLojfzWSLEQ4oyM0hXIAoMzyMYWDt8gDcgRaNdvVuOZEaoCb5D0i7Px
hapzKFTva/7k0K2A6SKhqWZ5zDnDIIeuATxyUbsIcVjKpkKWKUzi+HTy1B00lQlw
d65NsEEXYL8K7GVaTu0F7hlnphaSaJVLV+JFb0G6qfSvmVnDzUdBblLP+LNL4oB/
S6MilDqHgfCiDBipgR1Hb8dSUGdzgIjjjQVD4rfKOc7QPuuaAcfmlpge+kjtrj1c
uCOOB9KvCLAK5bpCbFEG0C+jngX5v9IspwQdzJcr+hBXkNsG09qVqfns/ZJ/K1P7
LoSE3Oz/LN7HW+Ui/EGPgXvr+CNb73U/JDMQF3ALQurQlXEmj2u2rcDhwb8oGI2U
d5asACV/cyKKllOnfYwP9PFZqQ1+7m9tenLgoYag60jkLmWCM9s0QItRrH1ireJ7
BpJvy7B2JuOn0k8KKtktwVyxXWd2SmyNT1qPJsZnPrsltGdC9gqDFJaVsIkZO9Tq
XNoJOZiV4v8sdCrJhtf3TcGISCr1IgHj+KSSkxFPyxLotJ2iof3OUrit5VRgFYFN
Os0VW/PweDgnQCAFXCMAZfV6vVLVkaSCEMOzYzEtNOSs7MIS5zK6bBTcjki4N+UW
Jh2RXM6UNJbFgah6/mU6bwdPtpndDvw3lGsUGw2pUC9x97I/f1bYiLFLNdrAMhSa
cTOGqkGwlgwoHtjTZ98XO6j3aji7c4AyWVwQvYFz8bHObqtPTv3LURGb1STYjsQK
+8+56i/IXIDanpTOeq65iiz1JlU4eem9KSxjIHQusWTHrvw6u3iLwGZ5B29+bbUg
QPu6PtdJkTMpmHRABdP7oJHIgEMH8641CiwOq+bKgAz0tcOAzGlbKh86Kh8A8uSW
dvAUjURrDaF4eZfovVVR4wwOEZl28oPWPlpUFgYwFU7IxR129M0tbTKNi4I7KAoo
sfQiRZPJmP+S1nr5piLaGzuoY3arPVENxQ+EFwq7IgZhpF12BF7QmjzEPplbvOQB
ZYlQpePzgRCjuyGdO3Bn9HEEk7SGuVoak0R1YRvHFZVXctjI/Kxc+Y0aFoH9vDES
R/xxvALIpxE/v0mxFYExexF4bJXmXqSxe8mPxWWkkPm2QeFGbd3OOoPNDsD+8FEQ
tno5b27JHBiQb/P7FrEV89BjFaOVv56lDh4EMA5mmnZZA+Khj7qZzJNPP5yBxKvP
CqPFZBtnyaSElZHTjB+42NnHvBj4pWhCGqI10LDJqA3voAorAEGV7igtwb0f/jD9
ege7V91MyVSCucPWX0PhHhg2koCAbUY7QBq5Fradf8M006CmX5wYiPAAMA8hEYxM
QifEJXCF4cTa1sVn9VcmldS9xD6fPCKnvicdfFhwmurKfC9J8EMfxEvi83VbVJNd
FpLtSKONUIrtxp8v/iXE3hNTJhctGicI8FHiWWaXWoCGfnbKTP5Ta58T/PA8x6jm
tTV/JZ5SzFIwbGJjo5r4i4MOD7pLYltDTpwBhHE3zJkYZxb2zU/MsmuJEbDSrulG
ScWGWNcnEVFNcfwgTFYRV1JbLjE2KezJgGsmfOuwzOQVB04GO/uyj+H/Ri/UcMBM
0r1CZk4QQbuLOdhfJeWt2+eJrP+V1/eY4Zb3LQQ5mzh8j3OB4R5ESn8w5HyZZ1lL
S87NggoE3bFkNW77JC+7BKCAaMw+0i4Cu2ymHUD6XEtP0p58juFHB7DKBjQC0snV
ysyC6jS6iFq6Vyfoe3RjyIl+ormFbbkN1i16GvRUa1LuZEDfbwQ+n0YmDHyQ/+qq
GZM9REOk5m9c9CDWtoq5xbo6FvPYrTmYczxRqXnbgO1XLwCoLHXXYzzbqJULDzuq
leG+CjRs/prcgWeJFA7/ETwGMr1rUwvIPILqHfuVwQyYgoRuEqQAdw5TP1uQ0hzO
0wX8X7t4TwyXifeIZ9zzT0pRpck85XocXvEdBENjbqy6lpZIF681prorqQXeUcfn
NXZNHyUangFBc/ApG/a53aiMMXs17cP0YKXNBpij1vGtkgUJ1bJhvAdIHR3LFcJR
9VXKDvo7h3tnOF1KAEbClA/KkBRcdEkYqIovCmHLJocaTFHD819OEU7Goiq4IIgn
Q71UECiVHJZbbvSLL9Oa9qFQ5LMx9TINzW2ejpzTCbN0HSUCaqT1LhRAJc9lHl/q
oqCfSFSBm8/AQ01D4snxPFiPOPxREBtEOh+Lw3y9fQbPMfvZ/AvyIwVwxbN7x2+Z
Ictf/X/oqamGz7PneqCn95NEvHNaTjp79BhxIXThqOD8Mn/hSTBjFyB8Wfc8fj86
ZdzADv52lawMUdBWnaPEOZ/7HVA6iXrXd/eQGLSZlyMCerrIOR8sc6TSE3bF+Orq
UKD18V+EuFkyyIl6Phx0aGO0IkYRQk4FF/tqpcA49AXtC1E0B0fgS73NhieNfrBf
bTD0Ya96dvkGqsntasLrkTu6soL6exq4EQSlPAsom69wli5SM5ZV1NCLsOHfTNVm
z/6zeWVeJvgWoa3Q0uMsrr12F9XkgqiVaVtA2AEsqpWyzNmjYwK3jvCmHlHV6n58
ST0ckpTDiGARh200ztMmbj8sKmNfs4rjgZCmei05DhJLKzs9ogh6mK7SaG3ZJFIh
jCj7p0cB5PssNls/HHBQ7NK3PJobtygJOXvEK3BKD7Yxg8F2iYObIO1Qo9kTCuYz
Xxt0YOyYsm1XP4vWmyeue5FkmD2EAq3//mbicFfo4Qw01ou2Gg6OH7mnyWYx8MPZ
BIKLLz8NV3K38FkFjMOACiL06CeCogos+o3CmasE0S9379h5lq44Thh4/RVA1bXC
39lnTbGof133Qo0uOm8gCBHB5bfvGjue6G4SsmKfuJvdlVC9knK4apzA/bL8JQo+
446KE0mC0PXqUyVQscUzlGU5M/dDO87iGh9J6zdlpnumTkI3HRlIXCZxTYBQfhPn
15flHe9SavmuE2bXF7+xr3THw4YcEliKfeV1TlrGld3L4czfbSY/umqvOq+i54AG
r1S44KEkCrOXxZI0u0UOsBiCBQaRwG5NAXmkIh6rLzCm7oUYXHWEmqMjHqWw4Wh3
CSjSB4i8z8EWkBBGzL2BOavNyCAjf/mvmioUyRLbX+F0t806pyPOHlCWr9/+nkjE
+FpAEyMsql5uMIKDWZeZp7NDZDdUfps0pzLQZQ5S6bpFraeW02I+t7zYCJJl1STk
k+0XktgUxPqWrELXlOPVoaLLquBhesBmry0aRgP/OICahji+zNzJF5Ya0DqxpPwV
0mLwCdPR1R6io4q2NILrnYK1uZoSmRWa11uh6luyVFdj3wVHu2leGzCVFmEokmU1
xSlsxOSD4QHf4dC8TyqbsjFUe53+6cSS1gQ4dBWzK0gLwfTgWK+RHuG7EUjm6kFl
HmaMvgLBNBkelw87hiur0pPcl/LZeT7x/qX2wFE/Mqc70wxRzeBL4akkDo3aETMv
2/61VpauXfV7XOluxhZlfdc77nI6raXgH6ztPx09WzMC3sP4ma5lBDN/I3vKoslM
Gn9YPZiydIcUF+Xq2nboHz0zcuGFw3UFSA8LcCFEwnMT+eBdaJhdEdPGMVN41tpr
vfqXVOYMg0m4cGuB2i3JL44t2b6ny7HGocENUecyCSHqxR7Fcm202B8HBM5SRBQp
xQij42nQFT3Mq1C3wX6J9h+JatCuH8mtDHCQZuhoTOhKHELvwe6DmI9osZQJRJMw
sMBN07yONhkXZU8zNIV3sWvjW1ecKjVb9wmH4sx6P+fy/B71V1i2JIxvqamaSh1u
EQNXywV9Omqji78TYLincA6qIyc/DZaDSsh8XBBfEvscsULi299tv8Cib9VKCiF2
En6VduMXR0HpHCtrRHXMpaRnoJ+ifoTKhNmCqf79uUlKCPA2pGODRZaDNDTl+UUj
UtIlLDkokGeP1G3W5bQm9EHjEsVapuY0Oc3rkJQlbO+tKgbND7nafp+xfFmu0Icf
Y6s7AkqvmQJH/OkXvetraBRDCXx1mKrL7HKtlA9HrqvF5JzAWWR7czIFwaNzfDeJ
BrBT0+BdFHxwM+xX76xeK2kSTAY+DHySTGrYfwuOb1vSBqwzcZpG2/J1h06g+lj3
l0ue8mO0G8mqNtu2Zw+KV+/nfv6RI9ovG0/HElyOESvMz85gOlT8FpNsYWE6jEXy
jV8x7VxccN73NdvSY2rRc8GJLkTQlTJb+IprQ+3uVIfy10HqTFhGq+wmMWxUiYr7
rgeW/0avIysgALWiGzvfHOS71GGs75K19oOh7S0Fl8s8FQvV1JS5McOyyxr5DksA
FV9RGSLVxmPUuyUPZ7ZHLMzmRjkwWO0YpCQXvXlB8/bZLLlTBhRZTOj8QfOVRco7
hFmVOJqltQRZWPNR7aKN7Cj3AGRdzuedWDjJUBP2pKjlpFU4b2pRW9lhuvq3N6bE
tWAFoSvHC4Or87N/Acjd9bJT6NF/Mm8xQIjbv7XKofqGn2FPH8q99kfAuaNnbf1J
RO1lt1r9AwEdE2o/Z0ZIrzPMU3Ry8NaoOeT6MNBvazC74KPnEG5AnpI1VzONu8TP
ug1lBvF69lcwfMWSHs76QeDfjH/4avYgoqOMnWNCkYb91OmoauKfjm4Na0w6lnT0
ZABCgnmVqVRQd86NprAMBF7yTkQLvYY10yuhlyVrub22rUkP7Dkvm1diXemiFT1C
G37DYdntGbwinMGnrmwAyCvJw+zu7YO6AkbP6byd2hUJ5A6lNXndFk24WLVpbQnm
mAHRqrO7zPCogLXSGDmArrdS1AmUgJFtJs2j5mHrorPwonXOaz2HjubZJPQM5K63
MdeM8JurEefyIu+yLOtlT5ZjLVJkbw0n6xWWKZxYiWwRRv6rO/wTr9/JqKIIHT8w
lErKbiB4vYCJhSOcz8Va1CusBApM5yYcuQAYsuJHLRW7SwJUvC8mdSdWZCfbGHC8
TumETtOCClMNMEb+ZVQ2f+thF6cZ3R8Z6blhzvxakMnXu/2uz8AaGh8ljJspc+aR
6WF36zXJZSJ6Jz/xu/ef0iJTtCuSPjERLSxbXiTlaXdxF+/Huu6I+JgOWc2OShMY
hAzHiccxfHbOkqsDBptEIW+ip6NLln78kcMdFWHL8ciy4e5hFflW4dFB7sxF97W5
3LMWyZ9sxgwj2+W29sqRrK+sedcx6ZGt+Rz4IG4aB/LDvn7G91OG3/Plu936Pi9g
RxZkvf+GWzq5wjPwQOoeW/Fr/S2hkliY5xUflQlXV7Rv444Bi9dZAoAbwF1eQimb
F1LxhQ7N+3Z0EIBsqk46QsoF68s0+hZzyPju8fWMAGB+5fi/4U7cxSiyPFE8fQ+T
S5nA3kKl93/l9lAwTBnVujoAM/6Cam7/y1w5yYLcEkuC9uiHmxSspv5Glcg9svdj
dBGzL8yhV0NspHYXftY4pGWuZGikO85wprm2JNwfWLYGmrFcAPqEl4caHoAKBKE7
Sqm6hstUZkprdkfZVqOVJS/aoGQRjh3XhHcqCz5kgb9XyQ8biyNqxZWfd8sBKO/N
iWM15rk1TGbTy12Iye/GVRNt+NRwVkenEd1B7F+scrvOkcJUw/xrFke+wniobDzI
0b6H1qF9tq+k+ttj0RNwoUcBhf+KcJRTXykk3/7GtbCOHjLBPUhJes3ZNxuD8jC5
q+iX2dhzt+Zqf1P7WlbCYlWZyFV++h/RkWt47+Q+yA6JcCrsMf/dn6t2s2yzffDy
8LY6HI7qXJiE7ViSuZll3A2zD1nuwDhyHV83MSrmeJTuc1M0n1Wo1C1lAuz7DisL
RC2ByGcec2QbIhgFfW3tepsL0THJQUtdnWJQX5cmtSSPHObDMym5a1bTvkftNgQn
PrCPNE2/dKJkRocabPKaVH29x5mPz9QcrZNDv/9p3PpLYODg+O4fzR20FRMD7x9f
77LSuQFTAmihygqWitpfGzlwr7PQFcgruTcj+VE6hEU1W0NQjBIc3ZlJ7r3Bjlb5
gEOg7Cg0tNcLFmkZC665XPP7A7fKt+4gYIKDkBLqdcyJtadlnu7ubORTG7p+S2IK
w1NFlZeeL1yZmZc+bZe5CJbWF2IKEe78QOSHsvM2hBOmbr+z6fBN++jicjCEB8NI
/ti5QVS+wuGTh5D6gJmrtuGFV6fxlpXQzaraKHfHIfdM8/l0SV7zUUkCqZL2DjRI
cLrM20kt6nk4YACpBP5koAtZRItYMMg2bC2lbgc4b4KteQWpPFzj+tCCvKRFbHmj
LldS7PseOw/6xg5cLE7y1QvPHPsEpXc+Y693ymoJi4DwkOAp4PQ2Ojb8JqcMDQIv
coQ6TeVumHSG9uNtwfwOY/gGFUt9pPQgXgDu+e9ixQzirW+cDnh7NcWwQOO1ukTC
xzqGb+I3xxq95UGig05QKZoIMYEWtDJVeKAtRoP185ReClwaBFToVvpSMgaPg/fm
llMyYj8TxPmntdB6vT+29cvK3j6yt8+Aq3yejaGzeuJj12cguhKC4oltsenD9cR/
iTMg0sW9CDMEsX/BD21L+/564XqsfT7Ljg8D/QvPWgSLoRL/BwBcpwJl0YWY+v1x
pm1DS58L0JcYMKceJgfIvde1kM6sRlo8CJ3hin/3ImyFmx17FSSMIiQ4oY9g/0EM
0t5Xu64uS+UaXePcGI2UZZMmSDs0dXa84ltFju4+lxOZZqwq90m0nVBCFPCubxoZ
HosxSqObXfhbk4wXwrULnf9VY1AnZG1BICPMtRaswrqEne3rGI6eH676Z25j6nQm
i+yEKr112ZP4jJZrur6JsGvlPcV6rpfvhqG5Qvp28KKlmeGzF/SsW9OGXM5JZZ/a
aD3XEDDZsGTnHSDMNaZdOYg8X0OWvBFe4GlSCi35GIBF/VSOLnpEIKBcYUmGYywR
PUMRYexLuGuUoYAmuWNClUQlLxHbKzKI+DiwzMWjiOkJdBBn4wZS4doWMGMEl3Da
5zTrGcbzs29Hiz3W3X1aixstN74NrrkGwKouBy0OKsUySMEYMlMPmYs/nQ1UTnsc
sMMwdHd9eau0VQXUOVWRe6LoJ2O4bOwRe3cUA+HHiQSFQ/FnwDkDJCEGBLfO1eco
bhZ55CwwLsPPyp+fWmukqX/g+AIBEqpqvy52JwGYhSo8x/PB4cTzYtlZa18H4hQQ
pFdQuORRNQzIi+DtEwBZTnkBtgZXOuCVn9lxZiOL9KtpdaxOynCKbgY1mBZjNH6f
JSX8qRroppRGwvGrZ0ZSXIiHtLUui4nKVe+02J/mmjUBZHbjDihgKL+8AORj6UgG
DrWNCPtMW8juIPIoRfg5QAUGyXrIXMTxu8FL01Dc2EuXEi9msedtZwlDpX2XAplF
7kxBvDqTYCRvdXrs5KVd2g8IOHq7ab/88mWp5XpIQCIBrZmF4IxhtoFlf0eID4lP
7rfy/MwlCaOVLqAw/mas9oWCM/TfEiQ3pgUUJVZNs9FzzcHqxWVNWjvHugK/0lgC
6H6nRhxeqJGQ0J7SAlNiRZBxMI/rLjYv3DIzn3W++E2GKqC6UXnfIAP8hq+mg+NS
nkY+//5G6P28RD5J6ZisSmAbrwZweuiopBky6r/Pg0JxV3CvZ9Z/FBdKr77ceh1I
/Ghf126uKk5whKXJ8btztYylgpdfJZSw5KsGwUe6qJ4nKfwPkibxYKD2hkrb6tZp
UosXx8lOZTKorfz/zgDsSnM7M7hajvRzm6pxMjWnNayAZ1+ohDFOdoFVzA0f0cra
4h+L/Q+cQH5DXYoMzCgaod4fADDHRcxUfxUAHyq1onJFyJ/A4syoWNX+Ip6Klacy
nHnnJ0oqXExGODspuCe+B6tt6SJs+1PJpOUb/bZpSGiZ14R0aCd3GfL8eOGIiS8p
QL8wcew6EE0apOWZWP2iFSD7uflwanK/p+jHtK3j45cZVpHqRxsN5UztIcPAibFq
21dCGupExPBt5pXABPv6hlRr1YzuRx2OMXYrqJ2j35AWK47ZcT9gRrRrXjalzZwr
RwCyGWxESfpfYFxWTi/OPgXy+hzkKD204U9QTYIamN37d36oVlkb1fA+h2jnq4pJ
hcxhsC/db1QHFzKhtk4CSW8YOctMy+vwAy5+7sUDUR0bx74+2UELFh6FUscTx7NM
t8Sg5iIp5jNwR/MQSjR4Rd/a0EnekTddnS0hNeTZqzr8SGq9lYYneOIYaJ/I/uZf
yVwqYk4/CEQSVkLU3yoo6LBxnMj1N2dub7ljASp+zPgyctftw0qJg/TivtsxZHpN
PhlbSjFwRf/qZ6r9W63sSTrDOiN+AWyL94aC52xFdLQTCGplmmGBtyecTzAUOj2c
CDwbB8OsI9eO7lRb8W7ePPF3VnwdorYf2BznDsCtF9ppwrCq4sJnUgrdLQGax3G9
OmxyeekOGRDVP/H47h33obWu6dcw7T1MRSYOP1/Ngfh+5esGlnRnxvlnVqtO7wKu
ZzaC7xiYi3um1gd6+kZNZlPnAZTND18TJpiKg7SgVrWrbtTJQFRsLS71ZDsFvKGB
eyeAki87V46jvxfw7uGmTHCnAZp3yiqh9BJVadgtRZ7dRMCvVbQauHWTYZcgpy56
rl6IPRachmXSb2kT9hWJ23evbMjEMom6VNjQw2Zxom7Y7Gwv7O+bI/gl82GWRbq8
0XYTBFT62MfOF5ClG2bzqoUI/JGjstRnb5d3vNRTu2wOcAkjEtTZyOtOeIQ8fIu7
jMNtNA5a+I9DUPpj0U3RUqhCLNrOLI1mnYMkjmfI8aderwIATd8UWoCcqC66lprl
+KCtV2keAXfC3Hgpijd+0t/r8SCIObxrbFDcN+h2uWj+Tiu+BYi49ahaYb14P6L3
TNQmH394DUYRZnyc9G1l3jnAzHknjrsJbblYSZBi/mimKC/EEQ7WAw4/DOfk3XGL
8NLTWZJicNB+MxalVVtNBJrwIkMMFGWbPo+PcROrK/qyYc9eMrWX+oYWkP8Ripyo
u4k9sHozVvHG+9vhkKK/QbzSSphs6Mxw7O9fe1WAQGRt8BHZXjt7aT2SX2Tg0WdV
+xQAsEQw0aB6rT9TONhBEW+mTSD+HHWYFO/3z+IPxzkhDuBkSXqpjGj5hy8D88Kz
y3NTVPJroo9tswSENSbH/UOGSUdyQP9X7SRtQUCDN10WZH496cyt9Hv33Cc3AA4D
11FCcKtCWXWc9pcmDwnRIhWF8fH9QO5jrdJ1qDRyAZ4KvfwVYQASWKcQQyT51dYK
Rof01dZ7dTqRjiLAPvDkONismve0PNQbOnUCrydObbIIsjHBluCryiYp/Jq8x1s4
fQJCwVzWyofWOKmauYAffLxYIKr82hLxh2AuwdPOCKJEUqfF6BrWBnxAKUHTs758
cpoVmd78LSwK5qUX7URHL0QxmxJ2mJFntPCA/guJO0p3oPnYESRkvmcfopeL12OG
enddCv26qVikkf72hjISELgPeBTKe7ArBoWCH5/HcG/ropFRLq9IAjgCNAHnqiVW
aMApVOK6ZJCr7VfaUMF9HdtJYc/uG4ttNAzUbN164GXOUESwn08nLrcinwbuCjWZ
nZjxV8Xc2Q5Ub7UN0D8kiciPyQJeGEAmUbQbgMZkTTYW7LUdkjQ3ygQLzXM6Dp83
BPhTXjdzo/MPNo+CEHkeSwz6iGF96CDDkSpm2llxUw4F7LISICohqPgJBaouWOGR
L1GD8UQFqOKIWUIiiNb+zfq9CYmhTDgJuqarGh7KbrZHwgkUcRdro8N3mU6fjLtJ
eSdDGNWJ0h8CkHPr48iyc0aREhEmYawjEgHmCUPHMaNdiAD0uEpVIhpcSJj1InN9
GpKFHMDAsMtgOWepBu8fZAJnPyopq4nz2alIgkJDnzxXxAFSG/D+COvofAdSczK2
Mr0+NQmGp4VAv98bTsaI1Wh9NhEMlPIpAx2lqCEg6xU0azcM4aGEsepzRTC7WZKj
qWRSb9GI2xsgNWLQRtrNGM9vfBfvpuf3RyaTMCb3HJlrAKRtUfatLTO+K7hZfM0W
xJjaLQizKhiukKJN8ZMKxMy8L5n45bichcZksmMC41VN2Lo77tafDt+rCnQRI8iQ
JLYpZbF2baKbX7Uq+kjcxqQywKs0VJGgLuouSVTDm0rvn5f9+UMoJ9+1tk3GwRMx
9oFCaS+4OS+yXTAHvyVMpE1iCXPkzSE905a8tqUvOpm6T93uIxD1CKDRjtka2VN1
37zaQMXsXqMyHceEkAGpHbCP5XfcJKfs/npdMy2CH2YUDXh8etiithfbL9fPvNil
YD3mBEna528c5NzuH7NUNdaWPfhLP7eXIakEfqPij52t84qNFthljpEsV0J2Ctnz
dLSTrZOdjX7V4xZ2Z1MARkMa/jJ23wlC/kACOo6pjSfcx35h+os0kyo/Kmx1Ei7D
udVwx0SVgbTkZyUYmFmz1UOULVba89VbOGmDfkDPNJQdJeIcsot//cV52tlS8qYQ
0YEnRoaxxMTGKLEvRUF5iZ9okEOj8O+2azgf+sKZ0LKxhrlwMfGgzJxh3RATHVEX
hbm8Gtln8/EZQYw6mN55j0qSfAmD2GpoEeBEkfJut8DOR8cURDlNVhEUGoWrZnXj
mNh65bvufWvV16IkwXg51F/tRespwypvmXuITIQGCO9iu8/8W/AcSAiSYEDxgL+f
jHqj+JF6l3Cqz3ERkWadkLmYoiZLhW1cZILDHbgmEF2oPUEimxoBp++lOxJC/l00
oKNdHMyFWT8Sc9UIlHL/LgnKOHaRT8uD1ek2FSSU/XDVoYn3+L46E9bMYPDqpEXv
iXLh1RZdx/97scZVEY1vXhrPvcyQm8617ry5bbZaEPEnxP6m3KVfaB55/oKaB8f5
BGbfqw1oYwzNNFtmbz9U05dDSd8TN/qgajui3etfgGNplErjGv6UwSReASAcd8mX
/Px4Ids3lM7pjzqDPe2sDy2cfH5+ypNn/ybvcLOGc/IACM/WbDvUbbm18eiH23BQ
80GazhxnOIfdsRLEGUGbTZb3RoTlFYptM+LhZWejbQcGDpN6yengRF1hMJiCDMEQ
iwVKJTLmBkZUSt2TCPB3N2w5ellWuB/iWFPD9lxQgVStJQLXlMX7pun7+Q1fM88Z
HMC3s9QktikSm+BT9ymxQ9/484dx3TUKFPEnIUtDwqzvGIDBsUlTmRK83SU6rhWM
lKrfydgoL6qhjaC2YKUja+w+7/FC8CWx+1Pat9Uoq1gjMnO+L7vKc2Dlbm+eioN+
PI7d3Z0VIei+hie4L4NNvXCSkd2xI5HjnUdLx7gk+6lv5dI+o63BmEif5nJDMx/Z
KKc7M3qbI9NbeDzV0LurfH1cOLxc4yXypW013Ml/lG1KxwT8+Yc3Xdq2aLsnEqer
kwBXFyGZPsCHLWjDHAZtZxju4E0rX327aV9MZbujXut4TW+E0Q+d14Eb41nUcdnK
5FWdAWY0u1Gwe9njY5r7VGeSuGPJaj/y+0Tr5n838RrbkxJuSBR4sZtJBoaXLKi3
nBpL6LrPvnlf189eZeBeyXNYx4L4IR9pwp2IVUyDOkq7MARPJOlOUqTQocZFLJgU
YQGM+lStY3mBgjc0XZ4eVtquTTLzjU0IOvZKh7KQrGAO45t2Vx7Q6Vu754dRVdT2
8y4WoAfyVThjDT6fx2Hyw74Y40TY3a15gRxrCZol8FMlKxbK6X3hQNQbjrEb2wRn
486cLIEi7NAWohaEbTFKXWzdOiQdcr5/lMYyyBOwEMMVp/CYCQzYPfIo1ATGUsEW
O4Pm3lfmm7jCLNAKcWwIeM5cVrr4fTBieUSOv/tjDRpsvuCtEeSolKeywSnAfzJE
Q6xuIvXfuySWdfJvfv6x/cGJOP3OthLOKRZ6aJPHzUwWACS95VBuy9yRvEW8gJeO
ffe5JufOGl9oxGVKMXknawwvsYG3dtAoJjetvaqxwQnmsvYBsWl0n/gYtq1vHcZ9
QSaZSkVXd8eKq6dPc3Ut4f1ADHcFcClohcicNwaOBu3F/ufb1V5Fz6ebggr5pcXm
Er+hwHnYpyLGgB9RiUR0Jrd9e7p3+VA31n0OZF0shS878p4wTvOvaNNy6jCp53yI
PMOicFjK686oE7ELjCo7WUcjHnGwOTJ++nJne+J7Fy1yZ91ZGfQ5Q4e2zZ2xM2kO
GZyHYDTevYYWjC/PSgypvaGAVANrsHB43a4+4hBYn7i4enP/LlcWHthoOtd73OyT
bwxVArAjnm+1RNqVn/SbbL4G3r2h4JBuILmjwvaNacqeECL83qr91eX3ZBRfju2Y
ciMiIacZkE5fwfLf5UGpPwfY5KGDYxzhhfjFnTXg4nWv7MJdr0cHhJO3X9bKt4KG
5R9ItgyMgUI6deXRwYuL8IYcWbp3psmmAAdk6xiSMontgmjieWsaRFF92kGCRlCB
lqC6iYiIU3H40mnVcMi/z2F7F6USey8rVy2bTpaERE3I6bPhTGZJDxr4Cjs834uc
bDky2W46yJcVu0vETxig7YEpYXu4SZ1fcUdxxnO6IXMUBWOzcvh46UaV0qwyUvLO
LcPQPER16jpEQhvFG+6q41Lk++lL5xRCjgLZdrnqag/6mktiVc71gkU2rpAn5b2w
c81ZYX7QYqgsP3oE7WoHgWzYMPiaqoC3VoTGh1MpqhD2Gtr0LBCtdUKjomOOUBV1
wO8ol3G8t2JhSrqQhYkXL7C1RPYM1Jq5g7Y+4KDo4AOe9VRVl88meBjUOrAaeHAX
7TOevrxqZZpEpfKx6NFmRLNo3Uw8Anrr2iOHSo6nywI9G+pz0xctMitsISI9175J
KVRMhYi+QSnCd+lf0+b+Li13MAZgKbpVsgRHKF4nLyJye/HNxClMbLH91+L/7wSA
Pb7ATKG3pdjp681dGWi7j2sC3SH24wFwE2qMtxfPpXe+t8i39EcaIrkjizublDr/
isCXwAIkIPIaWbi8B5M1EKbT/hB7Q9n1VgUzttwGAtad3+F6sCHkiEJpeq2iES79
YHKe8+8e5UwvaLoSO7sgNZ0tTrm9/zTG42UjcPU8YSBYxOe5Ewx77VcJ9/z4PSzC
3CdbbS9VkZYqXHlwF3+V9vunq5/DBVPKR4+fg4W6MwEyXewS322K5T4MrfUuli/U
SoqVBDDEJTXemaX+7tGdk9c4KL1t4E6c8ingDs3ielAWf0Y7k5Te6dF0u9etv8Cc
zmbIFIfa6/WNVEJIQo/31T24CvfKbsBm0O1sBJFpPTjRH+6Ep6pPicH2pMDgrk52
dHPNf/H0LFDJcYZgf7LUNDLrD8NnqDmPHHNpToIGY95n5SRo9n7NreZqMVLnI2NB
clkLCeb9y2lb/lcpD6KuUClZMqY16wG5pvf1wUsyIqAwVX/RwsEE3dj04gwjy8L+
lC+4SegdqjvrzlwambWmmxcRCUnLVCng06ertmH8pWy/w58E+fy61VJlbI8MQFZq
Zqii7bofK4SPfl3dvpR+WbgFgf+RtHSPIuQ4QchEZXdpg65WgWLwbBEKcDpgL83B
bN1GycFhuPF+kspgqBRWmlL0/CgFiaCEK7IDjRx6xTUWc8WNX6OQpwMErEi0V3ok
g3pJN1ZexWenc3XFglOOYSpSMfZTUAVFWGk8Rf24/Fe6xRrapR3kSJGkVsGTiIYX
IlOBFK7F0G2bOn444hjF5JC0L29eqNqHN9ycX5AupKcW/Ds2gwSrCoyOAuKE0MZI
bQ0w4hFFxjjquw0/3MT6Twqd85Daxx81G5/TLwhPLv5ek/L0X/C9zVvjgKrojpaU
50qxIUjIrH+dmZ+3lzSjs1Wr7fFQ4j5Xv9mJKld+IfSmQHxuuO1vJpS7sx+YrXF+
Y3ss+eY9FzSZnFGd4ur+kMQOJBUFShynBkyYgGkL+9Es7ewAHh6zJ88/gr5MxIGx
hFgNC6+GOFryM/xw+5dQcK6M4nyDohorixAoHCFkf8VN08hHjuMZsGa6UmJxsvAL
a/+JUPVF2ItnHPH2z77S3Leef+bv9zZmCUMnxeWvKedyQEqg8XkyPNNfpQspCshj
kCmgWjS3K5ky9WXe8/0UrQ/svcY18seGaeuwX+wCRG3wBuTiHhi50SFphBKsXKic
V4IArutbfKmDVEsOy88ZZurkhrIiW6878g78Lp3YKxV+ZWlDcPxhwmoN8VTYo6Yn
HZPgjX7z8RNbqNUA/Uu0yb3/rFC0LAcNgghPX+tx+00s8NkBwHK3Kyhf6CISV4Fr
yHDHrlrn/boANuybn/j3l3846wNMOoNsyjQBxH+oMkPCdUlisYr57Z2v8nfZDYyT
+BdBH4IZ7iZz0LLKGNOkYEc8M1bXm5j1Kx51tzV68x/9zwxlibuyrOYKLDxpDYAw
+WLQJ/497DANhIyWm8bwJQj2ZQktbAIvborYFXrgtb/aWLyNxXXMqWzy8ShOxHHv
qZwOy/PfLHSiM3gAix3T2VM19ewce0BGOCQJEhngdK/tKEyrKU/aRRRV1nuEjOs9
qMokDMpXELYgt1r9SVm4LzrB1MKLso8Ssz4McM5Tya44ydgh5m29hDxfF5XzSJ5P
swPR3Hpg2jGZ1AFT8IAkUELwZZa9sAnM+RZkKsjUqi1s1mNR+fPerx4W5U/kCK9Q
DkxrcqYt523LCGU6pjLQ8aSbjNoK+zoV6wP0TWcFRJ3MHOt/uesgClH2ydfIAg/F
I6TG3s328eFSBGNrwNGWBIZwoEB1gkDbClPiCw+XugpWRT7cJ5z5dmXka93nli29
AsDio4afGrsh1eIxORmIaAl0oeOZDIaIzpwSlNjznRfsgounrhkeE3zBIfg69WKs
yx19WIpX6aVktVaSY4WzpcjtlMgs4oDuCXvs79lXw7CJ3oO2gHxegQA7DUmNvgPm
NpTkixJxlST/gzONwC18T//E56QyGL2kdPaLPyRbQBo570KTsd0bXo+KUiQz5ouf
fHWnWP+jzh7GmDmLdbO+oIoQtDmy3Afo2F/gb3YvHx2zPyeJfy/m0KzHI+Jl6mMr
A9oRSP1phkJ8toLDaEFLF7FnPWwyMWbT1l+bnFfFF7NaQPPzRRaZ2v4Jb1eLRQAD
jvgqfSYggVDnTbGEutg3fikm0Rl/JQRWR8Msw9pej7MhZ0BI03pSoj5dc7vBuAOZ
k/+FPntCVMhFy86PGcGXT+oE53IETqm6+oNY9CMEHVXIBSkoQOzTmLpot9tyFtcc
cefVhxboPBXOa+YovLcltgYXe5SLy1HHRi8sxOMORi/bD5yUbnMM7NFflpBoEOwB
gkxwBfmZEwIAd2Up1fN/Qwh0l3nM8Ffc9MPQh2CSnhKJ+DlIK+IUjIm85sb5xogu
Fzgv/LCcMHZR2OYuQtXhF/3LHti2xZURyKNFmHg7LpivmpbhCfWzifAI4hcvm3yf
hbQI8P0YrR51MKXuc6WrENM6Ja9/LBuKxYWtqM+TE6k3ILAt0lv9SA2aPJ09HwEi
Bt0e/pvpUvc2ZqTBYMZTEsTDrZqkfzXR9GajOp1IuDYphHN8pvKhDUUkuQsLNeVR
I8ibz+2jPF3r6yLjsoBlyUvM0UZCWut0MbZ4kzZg4ooz335VrM0JKf2iSoZwM2Ac
kUNi1SzxQiBJK3IuOliQniac/XYDno5igAH4eKAkca381QpFLRJmND2QK5h6Aous
0clgYIh7h1CYwLys3ZOvhl0g0ScwVb+CKaT2qDqYPQWXV5Y4J5CRBSvDTsz0sf/M
Kyfqubi3WPrCtOdZarKK1rHEWLJNoFxOMeLUowZnnkk1n4xoVzSlKOwkbLqHsMPm
wjAN8L0S6wSdugI9VUyqV+mGVm5T6JC9/6nEVIv/XXdmegijwWULc552SWKNYFLE
9zyMn/qCKnXkA7yEcPOt2e02Xsbjeiq4zWQ+qLso+wo7XGOaxQViIxe2B6fa8bv8
q1gUzM0Sl+7bWGSCDdjNLJjXfmWfDTehWQF2oBV43MHp65oBVg2HDfm5fPxhG+dB
7+uHH3ktbROAT1/at/ui6lEsTEZXoH9Uy9qXxudvl5/g/h1oG1PMGmz6sMbWhuOn
PrIGqLpReN3MumvAPg/8Rf59Ou61FIg/I0ecCIEgifCLiPcTNNHwYxPI1UWPxd93
f1HExOlnD2WyGSr5QLuTFTN7XqJaqG6hcZkln8O2BYviIUF39PJwTI5QyJrezoCg
wJucWT+IRhOEyqWpnXO388njc437qNho3vCjiwOi7G+IlD9ZqjJNPm3P0KhRbJJf
WrNodwMqPPvCnZIifgdLTGvX+YOCq6zMDRYVkyKu0LwaYihLVQa5XluxQP9SEMxm
y2tjzArvF62jbFOCvtbVhisko75IN7LtDG12G5FrE2pwTq/sRIfV9I0/yVlfWnEP
6N1nZxkZwsKAphM2cFw9BV2uQvLiDgNKK+Jw74h00Mb9OobKCLgyjVzPR29C4XCl
Qd70zIvVWo5ZlR/aBwfCRW8M8NbK/V8NFT0yOjKZkCHovXnoNpPz5Qgrq3Mz2X1/
hC01KbupymXfR9h9Ig7YWay6PfZvWKe2fY2zv+MBlNor6N/uzXOPMnJyCu4DvrtO
LUztuMTAG8xMCliJXzIQuHnDSq8gGbmWu4mkneSg3SFRXB9cbh1p2kp1oAywuABS
AR3xHsIMAhKETbejYV5lvszh7K6WMvUnxzmlhbVVDT/QSX6ue59jyrxmauKvHP0D
jF0++Qb/znrgGCmspjzMblVZMlx+1/13eLZ6UixEkXVxS9XrHevepz7ytonm3BoS
3H3WniRjFbGY09vzcPHDavJ5hFXSS7ms70GPu1aT+bJogFLseqzCtTz1joyPrhP8
xyuvOsDxkw6KTaNJofOlvXVQoPLGureWpVl0WM59kIB3iGwu8gU7Kz7XvNm8kIFg
CarDIgtprCSqS8LKeqIX1hRWxupe+y+28/G9yZEghv8YeDtmq+mF1Felfq0xJSWQ
hScL/ZHAEDrxz26dbnFiz6+uOrdYbgdV5Gx1mrQkVCWtaZuA/JtHneQAK+lecVt2
JOwq4dInVurdpZRYSCiSuNAkfR/A1/56wKozmK7HP4IJGUDSxIcN9ojFNjuVDnVR
KDjwVTEftUXF+EfQeEOJQN+mDgh7lFP8Kb+msZzatk4eZ03KCOq89NA6A6VjmyRi
B55rTM4t3jZstods0170yV1jti+KL0q5Tq8BjaoDWd7jhkM/87s4eXiL4Vs6+Px5
44J4zAWM8jNAERmmUQ7O1JSGcT98DlWSKOWPlt+lvbeojWBl4Cx6uTfBHIbfQytn
V/DFcgsy86cZDB31l1ZuH2zwNjl6TtLjAvyLYZGQLYwggoXsLZnMIfi6Jcrr/Khp
kdHQFxb8CgkYhSa8ZKRnHPDEseowizQXUxShD2ARfJ7hD0HalnLqy9c2DxtqV5Dw
VlyZa17eA2MFYtqhIlUSL3VgKa9y8ODV1/HrD+gL885Qw4R+IId7AiEOcCoXsgKb
2CL/0HQBRqEX2yA0Dvzaigw+0Tko+wnGyxMtXw2mWlkw16BJBal8NnLMIsHsBPvq
wEwjwISkJqKNfMd070+yiw68ZJCn+YyyuOqqJkF+FAcCqCCgnymBDFSymegRFFHW
pdUPAkOqufiw0csMLNCZy71wTKirniqK2U+Qg76IOMFWqIphauigeGuR1l90F+H7
et8c7js/zV43QJtN9IXS5lDtnDAyE7rVXJNDKwh5pkEoTEOb9AOIfnSpxOUBRKEB
NixYE4N40Uznuep9YvsjKMsIawUsvCTAt2ebN00C1e8zPzU97Ec7riGIB/AqY74m
VN1d5EclhWHKjTETfdkfqeiqGlBMO57eTfDBgVy7C4k6ar95NNS5dX8M+wFlrwDx
/UOog7aJD6O8rvPQrTJQq1Ar/GbyzG++fInGcCrhblxgfR9AfOrnxMacquXT7Rh3
nSrTf0ZrDJLScYIjvR9ekT8TVotxxOEA5SC77Sz+ofd4ItMPMV77u+VyQYiFrSjY
uN4fWghhVdkqtssaegL2hy2fZh3QmKvTcxbStWaM0UZHAx/nDNBnswFwpwI5tpof
NfSvJ3M4fYwyd29balgqXLM/brn3IpJWWxcA1G9nXM+AKKf/hUfO47JzG3k86INp
B1hKjnTVOoCfpIsyTUMRFpAC1+bn506kZsXhOwjBdqaypNHUc4a6H1So6UQTI9bA
sqUMxpg+p5w5N1IQZYJf30XTI9dAEz92OuGthBx1tus1aFtwhB2eNy2IPVeBOpb6
I6P9g4hJgZDucu8Bn/fxgQquIbKDlrY3ymGu+A+58uIFMW+MZcIalEllwvFNxLoE
BKyIQL8OcUF+oFw6buTispSsSMBOaSd+rU3lTBA+9Tcyx3nzgcq5QP3dfpkDtAys
6x4Av+pmoHvuL9glN8CKRcMB+If2R5BzWZqkA06PT65N1aS1zQewvk+OX0CgLv2X
iR7UxW3wYqgidIrtJPuFsv/rHSTidRIenzETwiXLM32BUjjr69RBPn2w1D4ezay6
bOVbbDopXZPr7yu9ISWV9noXsMmMQo2WB+2F0E9dl2pKyC8EVruNCj645YXGWMmM
RC+4BiAKPfwY+4+1CiB9V07Z+kgHTkug0AvBjE5VKMJaRHjB4qBgn80rQa8wZX2w
Z9GWgq/jiP6omF+wd5j1rHlmPp+MAvBm1X5dAzXQvtC3ceRVHJDkVp48DAcoGpGq
5lKQzjemnxyIaQqG2waJ+86EO5JQTgKfEQgt9zmUfTJC6gzaYNcS/yoCWUi5mDu/
YAYBbFRT2T/VcwO/XQwKRy+02sq5ez+dDYSG4ue2RWoNsgwskfodMSLeV0r9ATEB
0vEpIaAiBakIk885VDECApuwHRLdglzKJivJKsSaAQJsMeUduvHNGoUpmEJOlRB6
hfoycYqXZOFh+rsAjzsgu8t05w68Keiva9juLbyxbhXFMABLdiFK4F/50NyoMqZQ
RN25HO6FaaXdu4XNYF09JRS4jMym4dHLJ3s002fnX4RQ6d2SKoP0f1KGVQubS2JQ
P7PT/lC5eQ3aHOrJLcYw8y/xefqIKL4oDTsQDXvL592YVe+kz8eclnOieZF6iJ4K
RO6E1uK7puT2zerFLdaG9bokxLZWYlVepJx9vPah2nobljl7z7sSPtsw1FFThqDN
E0e102AZ6CTVhaBX2YoLzyYvt271jMIYoWcjLL75bJOyOO9hcCQkLv5Zgq/pGqQZ
JVIQoKzk5669nb3rHJmmJEiRqg3otK3mN59VcKAWM7/OqRxCjDw14ivkbbQeCurk
8p9uy5KsLr8DbwfPom9vfWlomodKlzC7E6royh5G+VjhHm2keq+dF157pJrBSYio
UPRiyfTYinUyYcYjwIWJFi/2QvRoZqnbKUbzwHXTSMM1rLCI7wku8O2LI7yb1Owq
cUJEjE7WxZ2/fucfwW60ysk9pIOKYR1fgbG/EOJ6OfEp/8+75K+Tzpr4YxeZ0elQ
f5fOfcdlJ/ZdZsGy9weCYxIUuhyctm08zeosan4de1BqGaIWTsk1wq+d6MWb3Hfm
VJ4m7opW5IqKzP6n2Dcj6CbTyklaTDKscQn2IjaOOOrWrRYCCYAu76EcpOdTAwpX
8YcdwnLEJ+5j3DCpCk1NGMYcnup7f0VhRys0Bph3FvJW1iKIUg6V6su7CzQ2lHTN
BU+s5rFiV5aioxe3EIsOnjnxAqBVLdAy4T67wIZxCYqwKfymNUOHbirS76wAj6tl
pQfmbz3gq5aw3us7vqQqi5jyi6B/U5aLMY6zvMlyRc102MRD7ttmaFtcdVsspyS2
242aJak+tr9DKO57e2Yajk1sbM8ecqMtFtYd1p1W5bnl6hcVyTG5oIm3du3aHIuj
MZOLmTmaTp7Ype4fRRTGNwgpdi0mlBtJzOwGnSxY4M5dTCipHGqFMIKckv8G81Qh
nkVbzNlT7+eEQferNWfI1hBqlTMZVOHaolYmr9cIPYiXT8hWtstu39UMjV3X/bJx
b07eRrNIyUe2z09g8y38tgVxXSUpzji9HZVg/3U+u55a2xeCrwHCHk6li/A36MWM
8ieoazaTW4vJvsNWXrN0Y35eNxAMvxfIz6NEHeIOLBVvrlKzNAlVeWigqd5izKkB
gUBoeirY6uLmhZsaLsV2hm+iZI242sb+IuXBwO7Y2MgtQR0WtQNNabhOMSn08mhO
0qdNyWTJY7P7M84mHmA5SfbclScAHc2S84QRJEbnFAtX1dTYRH+C2uJ5N69moa9V
npe2D6b9V5gnwivLjHOg3TVHJEu4O2mI0sERLB6q/YQD6AhzRfSfk/vjNSnlCrUH
LYEDDiPJtEecUYgoAYOcOHjKiOw3C+nEDc6wImQfpPxBpPiTEYYlADDnrJrPOacj
aa7RNjqCSsoVL59Q8JpghceEaQZib3EjtuxgaIoBjjszVU2oUTRrjxQxVsXsMFPz
pSUKWiMBFqtLgECpPyx22CFB6xkElCIVk71S0nItiHiBctBeRZZRR4fDQQTzVcDo
u6wj3hFiByzCUaYPqHs5PQBufz78etA8Ph9ma29ejSTGTVTgyn2EGDmYnXqowKji
1YQfa1s0URw6ohrK3QYU/Q7b9UU8kDhmUwQYvERMiuTBEGOaXLs9Rrr7DHGt/fWp
Y2shl4ToNPv3y5iRd416bkhtcAZ5MkVGFcmJEgY1fMRWjrXrwAw9V0V6qPxK80Jw
37F4PRhoM/NWKtNXAiDWQdpLz6i09eCvuHWeU+06RyqbX3c9NZLBjg4GgH8MSxy4
aqnnjCDptFgDurn62m/IkJvd9KlEYDghR8jPOuvqO67w5/Fw2dyCjrl0N96Hc/Op
lc+OvLQ4NESrMaYzpIlmPE+AOklpH4RKj4XePoFoTbZ4RFYosv0Dc2qV9hH7yuT5
aO3JKzt+ySYfZ48B9z4NwPmS4ecgOBRTDW0uNIKHYOlribIfdw5/DdC1iiDKit4G
Q5Khkkf0bEoQnYDNsGcubxTc3Vt3z3UJEr9R2wKTlXww2LLAKeEU0yeBbj98ucTw
RhPN77Bl1lJZBfSkJk1mFQ3a0UIGC6bnDXFAH92878TcrrKH/JHKHNNpv84z5iCg
bazkv4O81bFXc6nX3+0XI+EgjFbDUnnBHaKwNlqC1NhSrNv7F1B2ZMbqy+8DWKfu
KRCdB0jXBCndopqipLiUY59Foh/oqarqJrc2o5pZeZ3kUExgHVLWvFn8pE6jgwR3
67BdeAtOXGg9NhYpvqqx56PX/Yn3a2l0BkEF39qdnDOcMbcE5bUZNFM+PktbBTda
5ZHWWuoYXQFBm8N/8h06ozOTYGLfGVEXQ0AfIIzQNOunRRaqCW3iyW/nElsDg8ki
Z4VQMtz7gUs4cbukIvTafqqkJUG5LHrC5HB5e+rzJnrOoHpAHw2u7rsnPcW5bl/Z
9qrvejBc+5RNHdg7KovOBGPu4Jy4il/nWsqT6dj25zcKFnbuH7Xlpyu2TdDB8raK
3Qv5HRRabnNLugZO0AY2ssOrhQeWYfSE6fqaVgWhqXirepaIEy1AMXL/737hqzyM
HFZ+sOuIArOPKflWbHfiBIK+C9xakocGuynQ77JBbsuHvapTGIYL2FDN2ubOXnJh
tbXjCbHYr8xxj+g2QDIGM8HFXmOcCLiMKmxXCMIMj9Wkv+zIRpsKj44A6dJdMm/7
a42sX4Jv7TVF9FeVVezC+CvAcyZvz9HTr2PQ29eb+x2UEwoZo2G8h1y1kYWtqiNu
IAzIXJb1kq2q2GFrImeOXaWphrmnxJR3Zp2sQt4fdSFttwe5wX62xhbBbk0pu10I
GCj7xzmUcnFggn4vJ05rwjvNKo8gDULSJ+mdgmElZyayL/G2qt3FkbBUcKua+Gl4
BSPdf2pv+3L2Wjqj+Z5/GK8yNk8U+s9m5j4knWTRnuk+6Gk7sjs2XG3t+Fx/nZOi
zajny770vDOQsuWvNCnwoZGHgB0nyUb0uLMM5EATXRMDunpt6tXmwyAjPu8e4MU4
nB37QTFEI128YVnoLDRo7ydi525FgO1H6EVmKQ4vc6KSPMfbfnzATJdZMWv5jhr8
rJycRHbuQCRFHLEF/pIQPmAOF36VTW6CKIh33CnAtt7RhH/4yB+/5PBmjwp80WsR
NkNlTfrD6CRsPY4d44svm5GxYujEAv8inHZTgS7vOepLiC60xdnX5xQVBVMPRh0d
iACy0hv0Amgxepp0VOqp2swb0qZAHnnXpLjO+Z4zh4uHRIh+Qfdv+y8oWUXwuoZY
eIxHIHueQJBZjubX4hne9QX7FV33fc6y6hk5/IjzmhBZ3N/suE+AAvI7Hq79XoOB
UOLY+iKjj9p05mpc0K2InvWNVWjfTM/r4Df5RIobt+JvP0pJk7dM0fkTGbQBsfEi
ahz5/xoF7wXEabkKqN6kNIa7kBofOJ99+eAzx7TmRSLZaLNiO7XJTyWYcrJY4Jb9
WqPpggIkONIvLN0eRmLmCnfeiMxS0nIpYQT38Ey1lyGGM7PECu7IrE2VYN2ZhiZE
v78X3BTB4erkZsUVuQPgz1OqJIdx2+O3HKmeiMimRBMV7aE6O/In94Ym02m36sBI
k222i2FchPNGJC9I+wCgxKUVtyvcRwzDy2jKhScswHU/kjYaDmDYiOfo8y2BIzzb
KtIzF2t0WFb1qim4yQtc9gUOtyURtmCcidVU8bdfuTYyqN+6QelWrPjlB5B3GSR1
T+2DggcIpXpZRCUNiuoBG40ZRQ0bwrod3OKMQxnBOdMGxnmWnWwdNoXlvgV7D4Sw
vunzBgo03DTwaZN/IHsXYrunHIgArc3YG1SEh2R59w0TFs/fOT6h6MbVJyAn2rbs
GmA/gWXK1Z6NbCvOormk7MTENjpR/U+K0p2sJLURcx9QXj3nA7an5Lg3Ahc6u5uL
sRGhA6nRJmtgYJn84xEe2+XPQkAwycuDsetZgOBZiepvQHZddPCZ7k/kcQizmmI9
/GG9L6fU+mruAuunQcmm/IzCHgRD/9fcg9ebQXEb+9tp62lmSxzdn8niZciVgHiY
WVQVGH313Vwxq1Ib1FSSqhW0nUwR+XICmMfZ8+o5DHbCiIZeoxAtIihxh10MSeqD
aespXiVSbZGMjM6itGrA6wZU6BindabS3wC1HAOmnw85lVVhEKFIw65DCoK3qsBx
pb9y54U7em6TKennRiMp9JWA70BVJyLZ4lZs98dsiFyBwB/kHHcjStP0fL5+9fjC
qBrlPeDSnDbdmvwWM2YPxkgL+xl4R+fdgCjhXBwHU1hh1n+MnGU2UQxND9UE8c2o
AVfi4s1q10YCeWQABthhef5oUxyRas8lDVzmP/nTorNj5JHsW5yPOkvHMrdFuJkP
lltsZq1pCxdyag5jqJ1pqW/NRo+JLY9UudiwfT5iGFkgNi7Ix6kmW1ZXQJAK4t9d
vggAot7fV8BnmA9WIb7wNDM5R1dbS/tFFyhZbG0rdXZEmudf7lWQmlY+ORNO5fEH
wLy984ygyuaomp9OeEhE8rkSk7efnSzLUsGOhkGOJzB9bYfNy63MztEbfZ7ziY+6
OgX2Ku4MfD69/maUgc9F7HvUf1MMAfD7yyoiNVeX1N0/lY3miLTbH/2yv5imQ/gx
xwzM6t4nX3Xw7dyfksJY8StIxic9OBny6w0gf8bEj717m/fBYr/uZtFy+YVcrRgn
vor1PErPahEYR+uduI0IBt+XaCn/KWtY9ZhrwM4Hsn8vR4eVevuXnfS0Wu8tGxwS
lEwO55Qa8wGO8Sfy25SCcXORMy9gdivVixe6fsom8u+VhFx/54+Y0YpiA3KmbE2z
/A6OHolNyNuWVeAhbOZQTViZAiouSWLhMKFZ3IdWkDgLewgpf1Zl23FPPl+WGWkY
LmAM4XIZIaadraudGI0I8JggrUAO2TM8u8qDr7grkux8isH2W5ZXdoHDXso4cHPo
20ZbJtOFNm2qOFxfMnA+u0s02xE8csl8QFnAQWTDNPiQbLfqh4Vu1dTqK0VYyAO/
czanP2ZJEY2FmDU5OlJcwAG53ydS+wRUKxcQL3p76xfZX3uF4wb0Kt/jRy89Fpas
q2X9FPMa1OmbGySNspmIVvKQoHGblTs2CaIP6p53Svmg5zB+FX9sa5ESyqTsBhKv
n/vr90zBcfUg1CH0mxoN+XFGM36YwD4Zhsx6zlPcBje/Tzc+R6r2xfG6RdwSjjdP
uPe019qi5k3WAgEWL7kdQGqIx1dkqcbeFxWbGaCm2hL80qRIEToVlmvzjOGThtEC
n8Z7KqD8ldJWljIsYKMRS8ODn1PLF+kXcs2lrTQqVREz5TBnoh8BGG6WslrW8DRc
txYcQAlUldZ8IiRuVl2b9421oLowYpstrmESvqaXx1Dnw++mDJhh1hK74nJmFaLa
kBOd7bhMrRXQ/sj0tQIT0cIGqKsvNrul72LXKz7JX/kdvO0iFDPYe88uXvgiMsDX
a+YLlk1ao62v1s2iq+pO++7FATvByIbMGVClSJeFQW5YP7lvqSss6E0ujQYvHygN
3dieNiKRVft/gQ5Qi8Znx9BXiRTuEZLyK6Ix7I/ZxPuXaaQN/CybxMuK+JA+W4FJ
d2nIZJDN+aQeTkG9TZKx6dHddGlu32P4G50dDB86groemCFTlHzceH/9dyXi+fNP
yVZUFluvAO2jV0ULy0ctskOFNEEhXG99g18/lkYcZSAyWQORoAMC3u3WW/Lghiv4
5H6+GEIkjDhQTl30grmZiM58Lro2uzR9dITwSyt8sVc60No5crCTzqg02t/am+mA
QRmqz2lRmNDxe/BfMTVZARCMPIhf1NsDLwEIAY2r6ctzK9qh7Hv+XHi5Xv1jSuXj
1UcMgEgX+xJ0kKoM7JQuSCsouWjl51EFpc9HIGTni/IuUb4pb44CJCjX0C1AjwzO
czggLfCQyaMvfrCojASzBICdWkFpyJdqI2FE3yfIeRktMOfdC0fqmbe27zt6fQm5
obFkfEtTs0cHodFhawn2pUcq0VVKNXTgqK/7O0RtybP75jk84TkZX/jk/Hw8BWy0
Zkxc3lgxdNQ0m8yMQqOnn33Lq5QH7QU29UP0fVdRL0BYa5LZ+hN6jGoU+aQRd3jI
Vr+4pteQ3TlXcCoozBGUfpPpRNZhRjY8ymy34ubvXGwb5ddVXyhbvyPWRVENRoY4
hyGIilwQBW3m8s23mNgv8sLml+/Zalry7IEIvrKe2BCT4I3ZHBW+rKJdF2yvDKLa
v6tnj84STDjiTXcyTKrJOR37jH+xzvBJ7fqHAaL63qI7Xqi2vq+K2SaOW6GFiGNB
2C/myWJKtx/xxuE2jFJrWFOvod7Fix6KJz+5ItTByq4bKkGkcIZYONhxlpNjb7ob
ZZ5gg1leJq1RlEgjLc9NiKTfXUbuhGoVy3ykFbcpZRjLe2N+2Ce85QieWIoKcUlF
NH2ujUU/JzDMNscBD96xS0FiqJVbED7Mhpf1Shg/hdtYEvqvKm3g6Ez1kLNZigUY
KNfPC0mvhOBzj3if0HwZag90UMfbhZD80nC2aptKYU2Z+2pX/iTQJwS79UAmQk8s
74gaX3Otm+sYmfCUQfqRLHN9DlBrxp5S07UHduaVhXIBil0YJ3JmeW3Zh5VZbDoM
TrqvrKzYtGkeeLfTu+poyfdJUv7i9r5AE8S8ZA7rnyeqCm8T3FyGo/RL/VH8WyGI
NF9eMF+Pfq+ABW1HJDTi9ExcEocH12s++oBe5fazlTPNe76HTB7BUnXIlUDXM78R
F8lHpPLC3fmZkJ/wjCackSgg43dgtDMwa4TnLou5eNRjyq6hBUpWRChKgbSIpyri
R6HkA3bakdGIXIYMOFREwhaC9h8oa4563Ihw6IjqGXLVkMKqX5nmSXz3CIktcsOZ
LcU9PBID1fcYikdbz3YQCIc9Ka9+s7V/X/RqnM+Fiy8oS4DmVDXlX5b/yW39HV/9
wYQeo1UkDHd5X90UqNZOm+cORJS1dY6z3x9NZKEIVm5zIgQJZlJeZSrGMO6Zk4fK
YjfLkRyGdXG7k5mUZ+ylu3EEewiYLQDknIJZVgxkwXL36csoi8OGBRKIrrmAhV12
5zqXXIGxoZFv74orZhFpWdzZXPzDuD37JP1sRJ4lPcK74F1gLLgdzeYcs4QMPQwA
Ue4M2NaakIFs9+Y8NsCa/WkTA/Gx77LsYKMrEVdhvB0eoL6ecWtOyzVWZfIlxXhT
bX4pHRwesLBRPM0AMSltNQ8XNOI5+rMw1zznYJJ+NKjMN3HIIUO9RyihihofoZb0
/6cFbiqB2jt+fPfFnsIO1q034cuGoGdtmmtU5b7IGf2PJuKy96AEiYX/rP/2Nmy+
sqyNIrWl4Gpw4yqjrS7obfXhQ0dt6M84oZI+zGIcIFRFIhzAar/1ci5GHENI229J
h7BOvetL+hGTwkwn6H1KPHPpz9PJj4M3of1jGF1pncC0RtEISsVfI2TZ7GYIoLST
+UtfOGw8y5VGkUSoLH+W9HetTSuii8xiYwY+TVOjlFjiE706MXa3YLnM8Oao/75h
I3yIH/21UoiW2n03h83oh5rRqL1ERmQJ40d4LR9A2onsmaz0kTzNjx589ojWy4my
rUuKRIQCZzOYPCN5MvMkv6ZaX2fP0YSd2YdM4rbAOFutpear+14VfdzwK851tYKH
525Qn/kwGtR3tYtSn5UXg/nL50ktE4RGp9YV1zi/X+lTvL9blJdyXrvX7B4A/Gwr
Z6dz/sTTt+WYxDaZgfjoZLeZ4c2xYp4+jfAYeySiuY3+gIXioqNfSN/TP9y09zVa
nRyqEgkuXg4GJYn3GbzBC7BPtGVzKxxloLQ8I4SVQ7763ADBQIwjJxBkaGYoCrhs
0LdMI8El5ilAT/ogMVkj11jdsEE/msEoE+CRmIJbI7reU+nkBv1RaxBZCwztm3e5
A4BgBGNzKS4lnJGDJzLNnQdh+Gjz5UK7qIUdbYGdVSz0Nip90EP0rcWLXMTVD9kV
+c6xf2tmqTkxpq219fskgeBOM967VXAkwDfKe7xbi5S8sMvqW+V3Gfm+OazrelE0
jK84U9J/jRBh3FxfWXwvNgVhirF0YTMTyHki8osiIKAppY9ywp6Ggy7CIKGzOSGI
lr5FiAujUb/fRj2VeCytcztcqZta0bhmaqu4PlLWYpGvoLFtHZXsFVh8k6u2HLw0
MHVFPWQc4m5HKLDaBvQ485moHtLPgI/YP/1jeO+bk006lL6NUkYd61VLmOAOudfa
5pFcCbQQQpPxfoQexqOpc6VspbqDQZrj9wwKmFsTmblb0enbzQ5VLbeweJVBydGx
s0ERwZNwTDcbGS8tmz/2mYoxgRRKLZ0RDuWwfsN7jFNYjqJa+nICiY9eI9Gl5Ccl
/W4BLqKJB9DqIuLiZJpaeTmTJnAjGZ52gxctgfQc3RdMNF8JY1jqse3bxixfql2j
sL50DktehJxGG4+nwp6JxDgiGn5ata+jvJpGvDwe2UsC33xvkBWH2mSlZU23EXqT
DqOEfFkcSiaCuOl2dOX5JpTfEpgxn0em020N7Qxo5WtSZ+4ITz2+XbziO5lcLaQ2
1f9FJeVhx+eIs+BrdLBH/iPJkMQa3bOj6VgnU5qJbCE8vYte0/TFPMrzjdB8ILBI
ekAeHVjM2znnmXelUACp+gnjHkCPMpwx3E9qjeIS90zEBsN/hVAsi4wu4w7XQuU8
e7LSwLveOjBkYiiE3gJk2ZeHukb5gry51OjOfc8O9kEGJnZSjKzl0CQ+OsdrirRq
vyqUo1AO1Khw+qr57kLKPDDPT2kHWXksbO4Di4wEFyXw2YXHKmrwsp5tqqeI/bou
98uuRpSU+vdnRBvqwl9LBSgLnzWNyhgYPqJKnx73OomWplbkBQsAQmQAvsoYdQIR
C6jsvsVlRziVZFio/cPAjr1pUY8aFks6bI/pqpedr99jKoHd9KT85zMpEIQDJ2Ag
uo00CKGGfdvPUZXcmtwpTVOMd4jeHqa9mxs/JQDtoPkxC9ogmc3r0hOTzE6EXBTk
/zshuCEtKjx2s4K09sjjzwhTzHbVfsfGIiFpfj6XsStLiJMATkj5g3XD34zES+Sm
F1jOWo5tSVnmMDJCDRnLxm4qvvB5XaMHwhypoR0DhXMEQhJzXCOKzi3DN6OkmSJw
o9glOHUbZcqUidGHXQSSUOTxT70MQeHCtbz/MX1UPZJjA3R7Ry35uaWWQKAnyVb5
Jv9GdBbQLXWbr52rAEExH9jDypX5xFrfLoFJHI3rfpvCm5W2DjhU/3qNHKKtfcRi
mUCqdpvVuzYVA+LN9aGLeSs811gJAC0V73OYc3Bt0XKnJYI8inLZCf6lmhXIii6h
Uji8ySAW79HJ1HUK7+9/2KWlVhLzbiDVmE2Gi7hOagwoF+9TOEY0DM0I3EAEMcWn
RGTAB0dp77At0k6XMf6UrEHcCdovuTAhrSuX+KHdEMuwl73nQ5B5RuGPuwn67EBI
7N7PqLxUgIQPd4BmiTX7s9YyBsIbX1+o2dhPYxaEhTZgXWeCcPA65SGqiz0Tybc2
upax303SvNp4CplrMUBLMhUKTizwyfJTO+wIHjgUVvaPE3xQgQtgBnZgHlM1bQ17
sZ2t5gYPaZqUudpGx/kbCpPygF+qEboeqsxVYbT7j0IQytH4NmzcFH2aXNB/0O9J
hy5SLpG8KTNznRCbS+A77l+C0OL6wM2nHbqH/WcB6In35ZVUD5kLtdyJVVoqeAKk
cnmO5NhaXxo7IOW5PUoM3loE7w6DE99ihn//zwXz8wPO/Vj9ecbduUr6HMt5DHP9
y87zZvtpCXKbcbRffA1LNhfwL9rgZjPbZeqgtXLMJsZyhqLJ+Cjkav0wT4S3fqkI
mJCACPLFsC8XxfvF/ehsKC78112htueDlFFqMeFvFVtGQOuemeoz/RMQ6+xEs4ix
NYEJSTUxjGOztPjillNKHa3r9MG1aqAtq1ht39uzkR0DjVk8N1uzg1pmrdsPg3dX
QYsSSF6H8M/JDbv4er8xjRAzUxtjyqWXlmOp8sWPpS2Q5sWQ1Gv8ezeSjyK+Vc+G
E8LFGsT643RtHDR94FN5QfYEM+x2CPr5o/wn1dhbLCTKm6n+z59Yb2JXF7iAQ0ni
aChyaf5dC8BaaqdE3cTeBbIB9u9LRS04RN+F9eIDo0jeN4lIPJC0QoNHBONSIRNN
YapS3vR7/ayTE4hc8PPz0KI3FAhKbo6CVFt4oRfVIIsZfIAjM7PfOssfrPQUIRPo
VwO1R9Tf2g3Ostwjye1K8Nhv1JpBWyUXt+U1qwNzHKjK6wGc8hDUDOFIPUTbHSmh
GYpHB9x+D6lNu/4i4arEMGz9lqqa74Rdhld8Qv3UunivVrLgzlITxym2FUecYwGV
hkvKyfA6FuJUdHar+0OdTlJh96pDVt/fjydzrCzRVJ6mRN+m8PCcOghVyYT0j6cV
fHOoFLwrQ0INfXBQepPXPhA5g2tQDeQbQPExWfpWI0gRoYZSdwlSN99SHOH7KCY5
1JVCaElDmZn00+xYbGXlUlxlAM2QF4AqErLdMwtbiGb5a3vNUH6D9sj+I8/8Vq9k
oedIZ+J/fNRSQf+XXZYVPIxE1bkSk3FED4pinKsDqelMuOWypZ54JYAvZrYKtBq+
Nk7m6dLdHW7aHAWhQWOhgTIaKfhEeP5f12uLGLtpSlshosSowkXPS+nQRLGBIBEc
a1rf2+szpsqLB5kuThjMQsc4lO0n+co4E4mAw2MpKAET4QpjMTMjHhl0gsOAMU9B
sET0g7Tf8y6Tw08wgs3iQIGIAZCwzmYYSUiu9LJkHbajI2pKQBi3aJNCR7U1IH/w
3OxFC9XSruNEqF2J5eLshEpgEYR/kTJy0P9MU++57Rm9l7TjPxIaylfGI+n1v00l
YEeJ3YW5Ki9alvGTB++sSACpS7gMly6IsAA2We0hPrZOMVqzSplhxWj3etaQU13y
1srSE0aN4/ktBfgJn+PxSA4G2bnSgUCk9SnM1FQ10VO7qILLVjRqQ4YjT5uWCmOi
YeNNM1CN9FlXjUgwGbJ7oNu8NCSBDzns8yVzzwHCVl0dw/uH8oT1yBBw4h1T4eOs
J3usIe989Bm1AiWQ46AXVJHvfqZEFMVX5VbLHZ+bViJo9ZNyCAuEYSfYWs1yfL9P
rJbTXlPuiQRN/1p1k1CpX+YKv1zAvcLGzxkJMj11hVC17QLpbqMKj+liY3ex5Vxa
Q6v5ndFThCgAQwMOJDP0Hvr4dnKZAxrYxRLAz+1W8bUOSOhUvdH47XRK2CZqeKY3
vnysnZ1z6MXmx1NWHSXY6Sy8oJjv1IdEFL1qJEyUTqrS2uibf8NSPsvba0t0kzyW
uSdNpke1wwb47t1HH6WyiD7Iutm2CsU4RiGFSq7sIfVKaF6f5baX55Gg0t9wvh1R
rmvfJNRwUIMEN/Mv+dVvE+k1rbl9awHdQUaRhy8meABJ/ZDdPmckCUimX5ZhaUKF
89gVd/YgDwNnbWLoYjujzFHSe2pbnAE27ULbEE1u4pMaEXraUxLSckbeqVTI3BWk
JHGy5PRy1qSa26JeS2gujOy7t95P0YJRBk8NT5vvnLBcp06Pl7JR9KqhgxxMm52G
3E8NMCGPEvNoWU80srFUJTMywe3VYd1dBhzlzdxTxRPXWshHQyGMOBpuNpaaUxLv
TkXASbMi9mik9OL03oASA9xFquffP/n4mmj6Z5eaIOl2FqABA7p88W6XAWhAqTFp
lsZa5AX+tPeMG5cG5YkX5ltYfhnHM1W+z00+01YkU2yhVrmoa4+1P3ihQ3Q3NLl/
SKomB3NDjIwodDm13kW9TIOWIAGcaMswJF4TBHZn9wwcW5lQlqEMZy9m0CFvRqr7
w8eg9nORzLfDBuNB7J6X/qLDev9EAgQ2j4WC6256tLDyhtjRghwXI6WtzoWHEAKM
GxMiFznlvtLG4UtzHLFHxb0y+DoLp3StiSjT85KlM8Sy5RqhsGwQNSOh27sO/xTf
c7rz+cOCa3fEb7vaIjgeTghO3GDSYrLhdkHJE2vliMh+Uxt/9WrS2FjURyZPZctb
TjLaPPUEvimhMooY+wLmWkp+DHtWziSdEbc4hn117OPGX/ez6aiZMUtgTLpcoWfE
0d9IpI8GFsNuXTRTOHTg4YJLsiEkh5XHrBwId+VOSg+8qVgUWcTnlI7KZeiGPSuI
LRzT5AohZzP9R/uHI9ir4nVxHsxD7S9Vbpy41FeLReSDCKNxfBP/5Be93K5D3lob
fwDMGEpyE+JFcfQOPT6U2NdIbvRziQ73xF+3Sqs30Cb5z/aA2JfDg48IwC9q0wwC
GcboWf6gBrAAYK7UCglp8WraFnBDN+pyN+pfSPjf8wbJphQRJAoNP2NeFYQ7nanc
kuvwHnx9u0D/bPAulvR64kSWOYbVde33XVV2LRRtNSf7jKstEJ4kAp8nM6o1AiDN
6Xe4LLVoGI2JS1K83HXq7XRRPBwobsA4qVKrZ1ZqudLJev9/A0+ecW2BhZ2RwCls
M2YtJf9qtHRjfR8H1Quk6J/ldPxjLSoWntllWnHW0SbdjJEP6buA9G4Zra6XzA7r
cRb2ht3+g6OrB3XPN+AgfD5Bpjzq8Zp8oyqyeD4xw0PI/41lZfbssvSV502ZWR0X
v80tgT4iZkei6Yg/+OtRomOfGsxrtdXZsJLYRZ3mcSXjefLSbeIoNKXgj54/xyUD
A8ChEvZohWGN4Bh4tMipuJvaw3J8tFiYc2HH+AbYcnsKNGfehnL0SxK91sVuApwE
gSi9waEoVNA/CL2vaAzD0DqAFM4yT8FYrP9ydGPAOmVa6LIuwWJbMwGL3nlA5XS7
i8rbyaJNDsrrBKy+TVc2Yo8Onm0DO3r84N7myyfWSZuoQfIgaOCoTojSfXmgXXTW
BlDRuBRRq6k03k7CqSFRZucKbYXxMMspmUdap6wIj8XQkLazCNOzAzpCLwQ4mIyu
xa/ovFwsKUxuY4fHmApq2I15X6pPTb7AbXOFTMlY2qjbcG6cyuV1VIK5Mu7iNoGU
5waMpwDUfhh0V9QPU/rbQ8gj+7qUb21yr7OsZJu+ViBAMd39lUAR5Q8U5wfNeeQ1
5przWbgg7RRXjPYwn4JlLsf+y/vZQE28KQZYlLYIUthUjTtymo1QbV5N6z2dk7a4
EzCENxiEZ92IfVc9EusUavUtmHYkKwnWAdPnnmwVmFOab0fMeXA8QwY/XWDgvfqm
G7dJ5JdfcL1peWdfzU9T6/URnMeWi+LCRvZMLoJjrHkzH6BcS0pXqqMimN/ppGZE
lHb72ZMrS/hkSainumv0YTAmAWg5whEOyspOvgj9yGuKA/MkKEEadlaYlp5Y/4o0
JSLs7jSUlUa2+pChxaoz2hgKN0w1E7LPsOhTQQHZgDeMwik5O3Bjplt31buwKC9n
ikH3wAOCPiym7nLMLCLV9VNo98pQ5t0J5UMw0JyUgBC+WKR89N8UN64BDmuylwTw
Ub1jeXR6UFxHbND5n1D4VK1T+T425YoObtBNJ7ZMjYjBosxQYtecreeODZSDP3+p
DMdWC2VA4+iB4e9+p+q1N3O3XkrnrN8bdM76VJZxPZ1VPUZ2TML3+kR3nPE0X9SE
Sbs+u8MMCsXa6pe3U/cI3b0vdlDw+3TghSjkOUlkPm0foAbEQcAo+EUxN2XeO6Lk
0reR0vRXiKCfSN+QxMxyffUD2fzfRFwNyUPQSG6IEwnlLAFWhi2MGMGFoRr8HsQC
+Hk6ZZe3v1Yg3QIUgfcQ3mhSpZUZ+gevw/4vCWOVsF452RFdwxoDjWy1gJqWg9+5
ozZZSBisMICwvKJEb0WEUyio5PmhdF5OQhXF1ncoFZ5UqWiFHDvX9Ir5I8DCsxA4
Sk1jxc2W8A4/Ti2BmZnhYopvFIHwGVTil0mMSeEYkca0Gqsrw9e6AsDD6y1HMcL7
rcJZ7SmKYc7Q0BUddSLiEi/pMWD7cd06u9sdXD6v02vaHi5fjg0o2KmsylbJ678E
CnR6eSjlyySQ/4JVyq7d33t5KCPpz9+dhuWITEu/msOOxo3Gjd4XKBrwXIZNtsbW
Bg4gnB9nfJdpBe7ZL7H1k+/2MWpDPctNtPXLnPf8HX45ybweJmWb+/Go5LS53uHq
+ifNNfdlF3RlNCfBrX4THjLQQVPakoHugKMNJZ8axmrujzZpgKisMV2XgI13+uMe
Wth0QV3TTzWkCPMyQG6CCStaqAz5QxA4+PMn+f/0TLno1ORdKfDT/2yQPuV7EgZO
MtuY5SHzxsYyvyMjQja7CxATa4k/yFY+Qorqw9KqWEzpQwlFEMjN9rc8aKiHSyQ7
FlnmUkBHqdH2HI8Mx/6OoPhx79CxQfmyAQzmbrMkrx3Nf7jUorybdcpltZuPeFJi
cDIGIfi2QwYoK81iULNWAWKtaZu656ZVOle9KYTieQBVra9+wCxymcYDSSHtxWLv
kDic9HkupV3Uj+MfhyW59/XXV3ANCE0VqHlh0v8bAM36kVXGgNHFG3EZ22c15JNV
8t5b+OM8qszCJ33vn/G04Xso+3jAnC435j/B7Ogd7pwNSec8HaQt73y6A8Dl1SHN
cUVszSQ3v8SEO+kWodJPNuMtmAhQCwchHjoGrFP03ey2ijfvVHbUKqlOKKzb0Fvc
TUqYrtPNGhBbFO02upJ7my443woPoIGQN/RM+XIop3XwXphiHh4tYxpWzez91z0k
EJTJ6Q9E1MqCKnMLHju671UedmFdi1GUUZqtOhWXThCHKZmESn5zOkWTBM12raRD
e6RbhstHleRsIK8K2DCgvMWGAgIoDaqsVHqO7Z6n0yQoeytCqOxLNTilRQcyi1IV
CHSJOFKltC1xMdikCEBPKbKP1doRsX5TTln9pmc2VVFBsNwOaIvw61PsGz0Pn7sj
fyHs0SPHK1BseKMQMIGPV6PTJtF/E8+6oEhLKVsYZAioQs2P5ltPF1OGMnQ49SEw
Bms7CqQyEUkoOmvTsdk6t8KL8/B4PFWv6YD0Zdmbub8+jgbxeNhVGLghwGLReHlu
lORAze4NGdVl43Z0stgqZFuiBfc4UP+6MGYJNL/H4hp+dt/x9H/yF2B5DVJsZzVf
bQppy01/Uf/+SQ6nUNHkNMDSPLK23qCzABgwcWCZWPDUkiv0o3nwc98bdiqpIzZa
KT39tI83bW0UNkxGIJN5qYIIl5XnlxeMtqQneLIvKqvU13mkzhi8TKB9+FaFFJnI
WStLt0ZDOi6gFdZDlj92fPLRE/oGWEasm9iNgMroLdmjjBHsSUpRPKSgthGFmqnr
s8AeOIsIQ0amWrGpO8OxJW/aHUMiUjD4hOVz7b5JPVdwVpGNNIPc9q3D9iH6pmOX
Dz9Rjm82ZBd3GtR3g6/gWk4nQlaNb7n333AHLoqWjZJ7m5cutGEOGKbDSV/duzCC
Llr6ZeQQaWUmimNKtQEXsGnCU6Zaz653DTxlRqkbGyGkgbKYoDtuF8EsGrxG6CB3
CRNo2VH/Yu89yJ0txMpTBmv9JurwecK5FMz9OGJ/w8+IjhkNNXvIHC6omlyLE0I8
hQ2CqE480/5NkaQn8mWa7KXqnAd70C4WkuiQkd36g8CGwayUbTXB8mP8G0geMjuu
w3ztlsEnFhwBJzxpQztcmpAY3leWcmG1bqnUvojveGZZLwhoJKl7cZeR7GI7Oc5l
fzyapwZCctqZy9/SxorHQeefbna1djQZfMeBLt9+XDjmYZ/zgOyAJ+vvPTdHZYxn
a3tnj8vDhTR6jbCCA2M/t7wRjwZr1alCFKpjUBpRvRfNTTKBk3hmolXGom2uTWEm
XakQzxvDJ8k9TebEciLwF9+to8+1oA+at2MrFw5ZI7O79leLNpOWBnaSlG58BKR5
XcYifX+3JqT3ws3VeNLVu6LWVl3vPE5TXirp/jYGr8iAgmXcbHWq4gBnem4qw6L3
ld42/6uMYcICXMNxFOTJA50RfikDG+9TvN+PtMydCs3CU5L3oEAM8kFRTzJqjnak
/qMKF4tKNSThm6reTt7eA4rmGUx45Vx7lhQIrt8+bl/AgQpCx3XBjzrTaP5XuJEr
uGe2pfTbVtflLDCzL+IRyfKAc/Vqq4XoXNwszFgzefVVFUaE63+9pV+WFPNoqMYI
XRFA1ZnOCuWPPGvx9oh28wrflCxpvBnGS5Qb5RZtdFm8euYQd13xXtubJrmS+egM
W7O4spvoa6roo0LDuWLw43Z3tsZf3IezH2vhzmK2yKsG8McOBjHmCCTl3/lyC7uh
6pjJ5UOqYyYthgTpW1atig+MghC/AM0dWjLkeu92fcC0usJmss219YvosxbGLLgK
8xrhkvFKdyT+kA0RRZAAOppYHPhgkBiQ4FIciYfsPqw7k6IH3X8nn1r99lM9TE6G
6jhap6Ag/bEchirgvaOgZ1ucv4fFji4GOCx9FAARunftiB6E7JuhhTNUOf9/w0HN
tVJ363k4H05dupxkKwP553S2mjZehS6ust0boLQoDKk6qUIMkrOWMlAPfFRbDnd+
wBQr7qVQfftajiqSC8oOn0hUw/vvweS/34R9mHa7pxRBZQ6gZZ+z6Uqv0I4Wyn+O
dGoN2XubSQGyjfir/Oymse2StibCgTazB9kaWIBIq4gdpJkXfY9jhqZ91alQPewY
t0VfJbw1RGKVvCna1L75Bsy8+djKQzHfgv8ecZbv/yE2HCXhoJXZ82KcEsKOICng
TvXU1mvGm1XsEs7tRJhVR2Ln4/KbERiE41ueToKmaw2vafPLPPwQ3sG7XHSc1agu
8KFW+nv488Mxiy3BvY18XPfJZMwUAaqDcTXzxvK2niy3il6ao1fnOPY4p2Tg/wKl
4WlE0UErV7yxlqJd7Fh5oVr5N8JI/APVH1GcBXWT/L6iJGyRWkn4m1uvFBrl9mMc
IyDsg1fHBynextYT2IpXnPTdmy+C55dMWAVMy+KkeI9mGk7oXr9dKV8iFNnTYGQ6
/Li0nVY6S+auhpUlndYYx9EINzGyfeX/AMrU7CTvYhn/WsnRaQj6HbVh4Vk/BVld
5gY44dCNYFMdHCm4NgSU0ts9RBx5d1sT8zNybqZiV4NfUatu9BIyZaNDhDzkwqaA
4zUjSuBstdsJXEGF4I7tP42h+T7Dhnum6+gfbXHEF7IDdvgPB8nBh/zY+Kp52ZhB
rqfQrkhr7t3k7zhRL+5A1n0FKcngk/s5NWQvrElLROmjzbVcDw8/cd60B9Cm2Fcs
iQjKiMEllOLjFtrpDGnAQXuAqcFZMQBu76SbCHcXnYuOKKvc179Lw8haO322xe/V
cqoq5zMAYbJudGXH8LRb4FKYwzUqKUC/7NH0mV9LsWDlKOM6w4CEpJT1fQB06P8g
jXVZ/VX4ickv73xEB3D8hsPWe1tjr90rvzUH6ib2HLhGBN+r1fNWeawonaf9fJzZ
awtG/4sQQzmaLL9jt7JXJtgiMRR7B0YtknRdriKsXY0lZXTi/ZoDRjFSSnwoZ/fg
Sev37qp8JO5Q7eG8JEcbp4voPtKlGOpjM7QI78Xhnt/NuSWoEZ+gi0n/tr/3wBUz
G79We/d+27kStJ0o+aFI7luJNigfRxkjzmFHdILEp7rbNAKfW7Mw9ksnY/prDRB8
MIdS27QeCbOjN6z3dL1YdZGci41B/VqCWhpQagNc3DqAfKLdq9idvgGHhBtcg1uK
sBfPgP6zc2S4cR1y4BhdBqQp1ykxOsMs/RhIvzzyv+3hspr+8N0dyfjuWPo19DVY
4rf8bsRsbV+qShiM069cdohTL+V4/WiJJAtR+l5f4ufyX6iy6S93pJYRoYRoopds
D1sxzw4YFEjAxlyrn7dLw2epC4LwtUCfpB4fmKcbkq9gNpteQ0WuHpwfvJvotlaG
2VljjvRCIwjJHTUtZvFwHlWVbyEReM1Nc4ojyqnfMViEnKYVDnrJ9Gt+/1AnG1Pv
W4jEWNhjh3mB1fpArId5I0NX3A4aBVGvufDc3e3k6Qbkzbbe5JypxR72zxIHCqIP
WTqiub4OqkgvMVLfuWsFxNb2ulIUqdax2T7Uvb/srP6rbAc4AHyTu1e7XRaqRnXu
pHZWDX0rYA5IhQReUN7qArUbOmD10PICxSFFy36iltDxHR/vyssoC64KpN9T4bMJ
6N30FKjOMuuBsR20YoXzklbRptqb9O7cEleieu1/7OjMaqea6CdUEJy936ziQ9mq
mRmueDdFR22TB5o3O1gCeTzdyhkBdjAhmodrDw9n+ChMVzf4qSnd/dKPKyJGLV+M
OjTqmmjx3mvp5fNc/QiQSJcmM4dhE8CKg3cGReonINCRPD+OGiCeO8UgdQw1nElS
6agMqlfn/W8vzTKAARdmCDnaXWeZ+mYgFic4nguwhi8nVz+KPneKqJR03zSnxLXI
horlir9LDC6wbTVkQ8YQcI6MpQRR6yrYibrV2neYNOHb8NGTQJLpqJ7mA7boBigX
lazrL0QwBKWWE2ST5jCQb125iMTZLlJyq+WPwUEBik9I6tT+Z7pibIuthxJq9B7X
J38fZCmh4INw2iG/dHs49ELJstt81RPneZHyvHxK3n6yIWQWEWzjdE64mqhb1hVY
tjkRKAx9qZFk/80swIKHGNEcapnyYPyfmzJ9ZsCIwgGkv7ztGxIO6RbWFZFEAkPt
5wi8xQvLFpVJYxRv6yAVuriDz1okyCV7cn26+A76UGT587YERGVjp0ePysb1HRzt
RbCi5R0SyUMHFf9MDiwaX4iclGEypiMv7YrYTiuX8kt3i1NZFIvbIu/NXTE4DlYm
cHPqk7N2XmwlWQostedruCFMc9ppuzZgIe7EYqomdr/lJ/QXlsBIJJ/NkfHz6iBr
k/gG8GUDpKu6QTswQVeWXrooxL+Kx04L8BAYzFhXleMcUjDDa4Bkp697ppNsxfUb
jqxYxWGBG5k++0EoPgpm+/RIDjlcE/Kqik+vemKbky/44vqs5XWAJBHxQ7XxGr6b
WnnY478/nS0GX8ph8dmLfIgO9i91063P2CepBSSzYJsp8YM7rkJh2aipr6S5+5yB
k1yWJOLGPpy7mRc5ESgk9L0Q4Yzv4p3v5yPdxAll6y/L2Llk0OCP5WPH1mStaY7Y
Wrp37Kw6AMWna47LLTFDzN/mREtIDA+FjQNDpCKjeUMji6uouBD7OUhrbrR9B9Er
YAvtPs6222vE5JcGL1o3kfkYYzo8jLO8e6vrRl1+13yGcIje6rV2qTXVARVeB/7A
fwyz6OnIf8WTtZMc57IfMD46vdIUTFea6WmNbj2G15N10s5mVr83adMFT11gXk2n
ycGn9v48jjCSf2t4O0dmyOGP6NPCX7CtgKF5W8ImoirsnMhVDzGT7qNg2GiKg+DA
EBJsPZNqqQv9VWVBjXHsoyuWfTa/6NBEhbxY+uTsHnAVw7BgIaXw+a5SJfwCWQU6
GlHUMKn0C3oCKvK87FkPjZiDxEYozKP7B7ke+OmkvdEfTSRtqByPVMLWLfJrREnw
GQOK1nFjDe4JWHuTgNj46IzCJUSu5+qZnAowf7WiRnZvkmZmNoyf0hH66VzSEh9F
wwmLwOEkpKgussTC/obBf135NDAJSjdQGa6W4yrsdZtr7IH3MSJVKA3VfuyP79NF
qJZ2FstPFmdEckuTd6vfYMCPQPxqUDqSFoTP88fsRJJPeRbt+mz0r6mP0qF4Oona
dFvWhQ17yYlPcxkhXVpyx6Jhqvri0UYr4V5bKQUMH0GLoErwgVLowKvCTe52DRMc
7g4zj1jjRMZSNSoBcNw4rfn6CeE0mE9WrQCp8uUSpCPz9pGsu9rQw/uDiGClletR
FOK4O2s7iEpVYHmvPA3E47Wc5woQUkm14pS4cX3f7VbN3X+aQBf9/rzhMIWNLAtn
m0kOyfzQBtazcVyA4hNFnazwGVV1YT1DKC+rC1Usowt8vRaPkJkQgtdk7sFnQ+pH
KTO7ErerDBPjnJAzZqZQCKoHuYdY6r+9VdwwQFoFTC4D/vBhSEa1kkp03uz0SdEr
+ku5xWhXSDYVxuiftJz8vrRHw3UcNaJmTMPpP9ngV5DzIEWVOKudmwhF4+KuNtiJ
X3AQxNSIUdQIe8mI57Z922DEjrcif+OVDg8I+y+vITYg32KgbWf9HXo2cxNajfdK
bG7TfSOFz5iM3iUPsjVlmw5CHTtOZeoexGCJz5HdTU6xStNcN9viigdDfIgBwELY
9q0ej0gvE0GiQ7zeH1Q4j1SLBSc7ippuejrH9rUsrneNuDWmTfsCJNEPknv7/niD
IS2P8mRbF53Qq46cRDF3qlqrCzZcPUE1RRFvX2demqLVav/n6vXses4+oWi0Pj4F
Brf0nM8J6fBa6b0yQr+7igRrb2nJ+ZxRGiFnYb7wvxZmcxFsJ4MAK/ETrpO0mUKZ
4h0CoQngYfCkjShObqehYaFkG/0DrSZJk68BIeMinW6h/6PCpEtApsVD1RXOHbOp
t949QoXfMwqy6I0yD6ltLfESPTbjIUQTUZZpFrteWAiW8l4tZFRqAwhFtfJaCtF+
sEQeJQxGthSHczniwlOw5Hgpr0zFZejgmyFoarOa9h5BeabixsUKfFO8l06dTKGM
8RIPZ5eLahRBiLyZEwqvd3+lGNFFgK0qnZT/VnF/nCoZHxzaFO2hDXqR855EUcDE
6JvV+XRIYK0rW5ZdQBz+xoXhBck8C5rn+CShO6YPZR7qIsVjxtsYUB4pAUUDVFVK
gvZn0mzb+vRWuIUQO6AOzs316jK/KTNHMiwMHBCmly3JRfZHINxFJ0tJ/MyYeCEj
0bcMCDvC9tI9nhH/cbGkbaDrrHHzzncAFXqITxqMG2Qb4XUx+Q1scEGBLurbAZWg
2Nr4YBpFraPYjJ8MVAVxj6BkCmNqv2vH2txiAYlX7o69z2T2FdA1rmd//6yLj0Fj
pbRK+EAMNW6kH6UQYaLh/X2Y5LSp4YHqqZkLNnpZzGhhLEAolgotmzPvKXMqx0Kj
XMaO9oSlneEO72u2ME9qE9TrIxBuG0BpEd0VqguQPsPs880P3cGzmFdrDF48LWV1
IRgrUDneMih/LFM63wGZd/qRYwtz0qS0XW3hXKZuSd2nJ4iuwR28S0qW29Qz03Zu
xAU01hUudb+LCmU+rMfddg/IBXUDYBLxXXu6AGi7RFr0ZLYD5fQBcqavNzpFyvhQ
zTbdCTmuv8AJAfk5muKUIDiwmhyRm5Ik4Bky8sO7c1MbnQlA7lZNPaMtGGm+SfCn
Nfos0fGQsfaUF7dPazC53+vsVgAiZAc+fgDtfEzIb05mV/jUA9nst7XDvYF2Avl2
zKrIMywMlr/dLfY92KIGSAzLF8b17HtLenxSnYBhj9frBjCu68SKHhm5OMUPMePE
qEjrRgIpwi+llXvG0KPkfImqNqHrPKmy5bo9GPkeSz1Tw3qpJ3kn7I0WuaJNB1ht
wQ6mBw5nfHAlSfa+b0GLfQu7GNxN0tvCbiut3NYo1rizHHXKhH98zaz2TO7b9TJT
BBtarX6pNPBkvCmq+fTTdMgWDaoMODlYcxYzybrddugnEMRMqsgzIc/icRSuU3JN
ay02WxHnxx2RvXz2i6OeKls6ymyOCqydpcSnD9aeLVpclkvdvSa2TXrZG0feZO5p
/kt2xgSmTpMGorWvUFdG+cs0bmWMVbWCVyA6IAVVNrAP3HP5StsbbQCgrt9Pb1gq
pB25+RDNe+Mh9vSaDL0nJ8cz4+/liXgokvSQEtOCN2bXZKrDV6C7DBVYNhMtbkhA
idDTn9jE3zgrZfCLbhxBLaJ3SbYfeysEde//ivmGbJS6RBUssTQIthFQGz/kSPtO
ZTvBGqyBaqD1zmbvJLJHZI+TwuPjG/BV23xxO7kJo/S8q6TI16+UAJR9geYvbTSc
D11zOgiU6HstUIj329zTg3YU4adF5htyz+Og7/yEP6jVOT5wc9MUL2Ael5sDYaWg
PYFMklWqPasncZb04G3xBTmKo0FMkb+FL8JFPjE/Dpg+8pk1z9fXXzHeX1piFpmI
2EZ8QpPcB6MJ/PWwDt3v1XNm01uu1U/xu8n+c27u2rrNhBW/Uk97V2mxpGUTVSM3
YcwdxkZMmTNnwvdqpptEOnovEzgZjbYEkmrxiuvEijW/rnSKHIxTiRuvBpLcxI9e
9MGccXdZ93RPcCdgpaCVIqqx4qdhH0AF1bRSeSqV0l7bzeqJ1MQKbMBG6wnKFoDr
pLtaBPxj7IK07cVoAR7MTcps4WTLhMvG7m+ckQfuYGQFy+82rn6wFrwGGQ3q0YuS
DKSnH6ZWfbKGr0Zmo01U8xNgu7xOcJDvQFgOSGcLUAiaFfo/Uubr3944AAoZe43V
CiXlJ9z30cBWnl2+GkjZ7jiVXWrfuCLnhcWAUjYmAOby5oWbp3jx+FCPP8JaU4NM
YFhSMcz+gPUHFwN+eSquqE8CBodeA3eOdewBJCIpPGTVOGjWIzbOgZ47ILwIeQJo
9oUFb1oXWA8lQViIXjqu7sR5DPXDiVPC4qz+XCx06uGEEgJ4ghreYfsl8CZFRMYZ
jaauAKlBJffY+2aE9p76zz5pupvbbvEZOHNDciBHiew0S3h9+RlrHLmdBe3BRg9b
wPSNn3CmBrfNMjHaWSy/3xhEATc2xDSMMajd334s2sJX0BP1T5tKJaclQ4vy5SKL
UYWm+nMy44j14ySg+3rZUWjTMUpibsSa5FWYrLxsqtzNMbVgnV4HD+kWFCY2Lyyi
txHhTuxzxCgzJ8MDIUhpgKmWYjBd5uHkTtrWdKExaw0uxRfgsl7Pw2VORT52ho2n
UK8S+rGkm7x+LIWFfIElbtHuCg24ES5S2IeUMwp7QgeQVLMpVlJsBXVv/eaYCUtu
ygjizHQeWKF2C+Rvb/2onpC2+VwN6yB5iGrNoURE+vC0REFiM0HwW2HVCp358Qgj
QdSCryuGqzXasPpuOvA4PcTUS8a8N2F3CN6yZPR/7EPNT/H5392/jxydRS0g2mwD
NFsM4J7q2gEzILfGcgbptXQz7O0pplmDNfg/xvdgwkg/fT/MPTCfwsgmajBz3juZ
O4e/nk61L/J6AE+Q5ISN4YXbJ3Xt/BfEQlnPyghaBWGTfIs2zK7LnFMDxLOg5BMO
Ma8pM2HKp/mHhWVfG00+YuT9rKPlfPuPWsBPgnPXmNtu5SVhDfYumhvFm7rd7sB4
ZLlSvercmnBwKxel9avv1M1nLw4NiNehBtjoKdxky4nc6eCUA90UL/qr4kbr1pOD
wKIyCdOqm4iFNlZSJO4/GFnTVsQmZWr4mtpA8+thclmxKaqXyWllEkF0q7hBfjhT
r/5LgFW0GbwpYKOk4pgQDrtagTjwGdQXAFzJ11pUnzf/O4lYo1bU0O84HOY7M5bC
US71XcSFKEdmC4PiRCNk3UoheMa+/3oJOTbt/yWzz4e5r3lbU4pfIG6wbue7tdwe
JTO+4FpARreIbpaZdY1VPSEe1rZCcstzs3T3aqNkxl/1cVdPiUisEXXYPK6y9eWj
c/g/YGqCu9nK1yf+me3r47riixhus2QSXRi9OkSCCFSj/bBohEsKUs+PBCbVcw8J
sxVazGVoGWJpvWpWskhdDdCGoI1vDgxTy1kKu2w6Si3grxmcPkOemBbIIf1qfNhy
mjFaKOtZRIgct/vVX8yerM5LKx24KGGHf41uM2//YhTcy11g5waq/TMvhGIwMuZZ
z9oCWjlj4LKm+SwVGlvzrYWzCrg7otCSIL8kf/kWelAvckgMo3vSrkbDcmrG0FB7
p7OxJBODnVps5g431Hg1Sii+b7jnlRlcDOPlT44L3JxiOEceaZqDzpYldef0/MpX
ArfcoEdWmlBHYQuZYASlJOPmmVn96ROFWRHw55r4t/sFVv/tFSRjGvtQRzby4blc
lJhRkQ0EHY2tw2LO9E5ujpkbc8h9k04uMjAYNevK75JAFgdBMO/OPKCjGY8GXDC6
S2+LSTWY+rhsyOS32v2Qm+K9Y9akhBrmdCiRSRqazwmvRDVvHWBmpyfdJBz72ydc
QL0R+7WPEL3b+Yp2obsnTJVUur8tCiW4q4OjMPzxqIY+xDcRDDXxXC7I5e0UvwVX
7nzqStoWNzZ7k0u3wntSE6mi9rv4nGT+BrjotphIlXPj332Xs/ZEkJfvD91MUWmR
R9i3OT+rO4huhcL6kDg8xaVQErnVkm0NZAPSHAQG6y2AlMJFo6WX/0hbAYRoEwRu
jG+AaNoiaibhp3J90ijFF9EzJJk38eSqKCC1yIq1hunDUXC2DNmBImAwdx9g0QQC
7CBgpP+ViCrIyVQjWuD1uhoYUjon1Ij8vyBYxFQK3hr2QUQSAGnJrZ9OElCyoWZq
vhx6bsBUhEK/s7A5uyMm0RNv0A5WHmsPyDLWxxtZXxeAGcLCW8gXDEJ7kuzMlRcF
AQKqtJgmLCvenvt6+np1DCAHlwNee8XqgVCK4xHJf3f1u4z2bLkDNlr0mxxhy3GU
zzbPucUHoi8zAHPZxEPJU7D8JxHASSpVOnu2OQtDLdCSSbrm/x8WqpCB4jI9XLae
B6X8p456tbfbXB0wPpxR6C7tVI6tn1gZ0er37hF2EMTPf42P6GEyNTtsBvEqzWew
ZalYptSTZPNtDWglQU6vhgrbGcnHmnn/3FAaVhzlfR1UcvlMU0Ku/AI6k8d3IMXu
efFNJchA1Yc1SMEg7VvcMEVotQVVrFbZ3t7qOFt1aYcEItWBOuwigZixWbJvZNJW
sh8e90mfZ21Sw6+4WKauBh2dUjU1kbSB1C5u7Dd9KEDkVnwF1ITNx7i595hig5aF
fcBNimNWvZLtgG31MmQ2bs9ziuVzxeQt00AW5uoWJD26HzvxXnZ4wo2Rrf/yYTOF
Fyd4I9NkwZq9jbSeqkw7naRMpUpPRZTVglueaC1niAg02OUUM2eyfr/p8+CKMao2
VbqvIyvc0hbbmyiuzINaZfhIxqDT/fj4Ohszz/BNB5auZZZH9VwGw3mFx4iavWJm
4c1B0ESmc3iraXcjKJXuV0UIdxcYxF03s46b3//EnWZWOEsJS7kg3evlFP8jeDro
7JsMjwlKXNnP62a9x3akbp1ScPYIqGoRaGsMoCQBh4Uk3c/T838IUj5m5AOS3OJm
oVgRjtG0tQni0pARsl96cutHan255tysIHlGfn+WYK8f7cs5scVVfgI0vCK8o8Bw
Vu0RK4vZmC7GCwD6ae8jTxi1dGy4ZrwVYtPoJO0teD4FwR1CsyF0HTWQekmxMZ8x
xZn7C3DQ2VnP5c8a7dLoRse9vFCYAsmwWagljSFqqicFu1kYF7ecozgaFkWb8nqt
3L1xcNYSSweZ7PTzU+bevF5hSQ554gEKM2HrKh2ggTZUdMzn58OLwctPsMRBdyVG
yrQRQ9UJnm13BGHRL99W0F3J3Bgz9OrV5vMaaqtzj1A2mOzzIfx4HNl4PL098m/0
wERZe3+g/R+fFpV/AHZnLTgsKBK/eNKc+rG/5XOjEQsScgL8hcl2Jizt1+H6An/a
xJkMaBMsZghSIhIPuR5trcpta01mLejgfdfqIs1xwExR8jF4j9dmUg4iR6tcLGao
Z4uc51l7de+I0PlC2WH93fBPN/UWDDbHQB8hjq013006NzfVopES/uZUt6W6/isP
f9X/wlOPp3sL02me4rZ7+SPCG7DJUBJUFnXFrlzyBE3/rDtgD5aEkFrYFM4tDpU6
FZh/wl1fySs7ZYo4c4d2aEiW0rzfNzkkRySirywE89XCFZGN54sudvhqFHLFUuxF
28ttVob8PASkXJ9HQ2LBX08jRbdGomzw77M8Wc8ZRhIRjuVN+EHdessgRYG5IUnW
cQNR3Fy2kKryV3N2qG7LPMRuUuCW5ogRiSsBjdAGSAEGnRMbDWvLfAVIBzER9R3q
FPk42HEs97lWknEe+hTUz3vyyySlA4nWhI17Mn/rQ6hENHlW+Noj2WxuSQ+1w1DR
yDVHG3WS/Kl8dCiYn+U6Jhp+rxY8PZtcb8YfjxvqQOqEUxG1Tn8xO0ki4acy3tt8
pSJ8mUA0bge1AzWnBAUbUC/1YuRnjWnIwo8akJVeEbf4VEqqy2MCz71P62VpyEXy
Xc7JBvCoBpsAgiukPcZZtsSof2QXnssbxUGXZF6tX7d3ZIp9vCJ4M4LZ26ZDJpY9
f06+TFTVxSi9B7+DCK5XwjlJ5haPYdLx4B040hNAX3ogG7Lc9d+hLNVbxPaZka/4
cIRNU4GK1uRKbLZ8mA1jbQJRt7+yUnrbdlROxuIe0HeCqdEMY8cVFXzzhWS+/yVb
tzPZ49opIufs2X+RnY1pCkw+GxRVfqHKJq11q8f7GuZxNMgMiafyHlY/rH+0hALm
ILMQ7aZPCUtY4OXtJdQUqf8KYrUPK4YrW+VOG6yl9MJD6khc8/F9lxr5DOUbL85V
mdfOnkVkgL7fR67/PGihQAjqRMyJ4gWcoRK9j+zLu9wtvCmgA9Yr7K79PzREjtRT
I7BGEe+JhPx7rHQ7lVIG9fL1IcQB7Zq67LjYLy98W1pIqZZmT69T+5B25fU/ZY4U
DOSQUAhfaI3e7GIxBzcQ9jNSyUpnjugafGg0iUylL5p0jFoRhlQM5+Hemlnlzl92
FEJY4ZCKaAQ9+6NOz4JSl79YYEeqLLafEc96IrCkCdofhEYdeAfBSqyhSG5I2txw
BDpq0WHsxbUPW2P9mPjuSmthhXNcffQQnoQCyMFhkUcxge3LXGp7rwcaI7t2YQlu
cWa9djhq5Lpz7Humtj3MpYYCoKPoFRlkL7a4dXH9InOLOU4jzBeaT0AJ4/Slu9wi
5mB74grQDPyFFuVzJLcnHBHnUDLMrkcloEt4ux4jNT1MUcjkfXVWOIv8/Ehq+hPR
n3hN3EDquaKjE8eqRzz8CinL07allQ4zqSiYgpi/dk+nd3J+TvbuTMqTFQ22i4oT
BB2Ij5P4/kLOpO6662oVvTroa8f05tSDUoP1VZEou5xqZD1jXakjWxlKHV/g5cF7
eIwBMAmvnHmi5zqefA58x7n0hX4s1m65Efg1BTwX+IZMQyNAl4iE8vt0HM870yTv
Ho9/soi0y6ISjIBI2AygE7OwghTiIkLjYYwJkVKY+Vt/qP4vco1HGDzrr5INWL3/
xeuA6ct6rxFLsqh7841jBMAH9jHGF7w2n4w58d1ahXK5ZDT5ZnttfC8CTzt49pmp
ZDNp27+YqsmeT/wyggN/4RdNBJpTbDwsAAPybVSxbGPlcxaonxM4MbnudF0uV6qg
MW6dzi6e722V04zDjDEwDT1mqnKM1uKFcKHeOMfP4CPnRD6pvOeffQiznk5zHnyl
PbfrMSbaPHO83s1f75NJs3XpELaJNGP18MhkgArc/PrWji83Ki/1RL5BtpufjVtp
/Fs7ATLjMSX+ky/OIs5BeUXKzHggzm8xCwPQ9vHsaXBGOoiQ0BeXwRParhri8Ieu
9Mty4YOmQ/h+MhMe75nnBSO619/Pf7wsVvWbtZeNzMD1HaQlnImGwAsG1bXaV22S
m1iLPbpvo6yeQoMCqanktLmh0TSi9PjwyOSDR6j/IAJAwotTDxPHZI4fY/aK3PS+
lcBvUhQDe331CYAJ9dqHVFe7Bbh8q0dPcoSVRQLbkO4Ffjr7aXQ+ezPmQrjuYU+C
db5yt2F/DcJoM3hPwMN/MSmhGlNyY79qSx07DBxtGq5IO6h4Hj7H/5y3p3Q4vkJv
xksVuMlxBjdYzMRtPYIITSJjgCW0sLnnp9qdEQmn6PwPsz8Y6GhwnNs++Ziv/9IS
8Ijjovy59oaNNPKfcWvkFOclJjMTxsNnFTh3ekJLmd8T2BUzq4372fIk9q9le1of
/xSKhZq4zdmJ0DInW97aZfw4BBhP5bqZXVT0hXWm/IKxcWjyfab/VR/kjNGGLuk2
v8zJFS8tJkPWiDwS7kgyW72C9p213rPtGAI0wddRDTKNThXYUT21quX4Sm7HnuN6
jxrERTDW3CDwdcfgQzvvuksmrzkvCyYuvCdQRNJmu/agjqqBZsrM7rC183MtOugE
k6cySlNYcVXjn8uWuH2cQ27y1MzstE4ht5+ENF5+TelS3aquSN6CzfJTn+QCjFDr
B2zN6qWeieDqpXFRGiwgNlkm9zubNjKmhXOwFK0O0nuT0E39A3bMrrolTRxtg+tE
gfFJEjdIrYrl29GzPwV+SjVrf9D/kGypEZF3vE69MhUGCLd1DfsAVCiDMcQiZMB8
R3IDhtmce5GZkZ3o/kgqWPwsl9rnKkNpI7NCFjbmBYr1rlQ0GRgF21d6vX9u7yQT
HN5ZCYjR/GoUdezLRmC6RIDdEfqHIerfO+93kqVUTv2l+MwTLknVJWhv7nrRAxgO
RmluEeuOGXZj7spyADWFm/mNk7PEnwZ2qt4jdH+GsNoA8uWGi9AHgW7+hrRvzMq7
KhLuUITBu3p8fc88a271GHwvHcIxqhLcRcWIJ5zfY+Bqphtovt3Yez6ckT/GRUu7
2T3p9iAEoyMl+W2y+Eibb7hKAJ6MI62KjBkc9bH/Qt2UqcpP8QGQZ7h/IiXBBmEq
bcCJoAvoosqV+RMytaWDSWqeYGWbneqYJa+kqtw3zeUuLBns8u7QurY4ma4e+fg8
TnS6yWSEbYD3AGhCuhUKibzs4XMDy8Wn9xq0aFsINHiIyFKZFFY1+kGyCHD6OmIo
kY6O7ysGAJhd+4M6Pe1+XzjT2VZw4UCj4s7w/8wNmLSgG2Q6gbCyrZ4t9RBicApG
btqIFIYvBqT5Ig8do/PAwg+PDQuNLQid9OVFtvKL2mKF5JDAS4FkpvxW6b8etE6i
d2yhSSUAOVq8Mo017YmLDEeBRbYXJikgPEbVAv+dQAIerskWUWxbKmzcB1ROwlwf
Q2FUvNpgwcneNKyVDxrsTsXTDDKuYI55SyZDEebTrIc27YJNFOaz3Nr4xTuxXzYe
KJMK2jRjuLLiWWJw8tt2gzM66IIQgIRLkNhdSzSlMRLKB3we1vPcqlzRY7bwPWpX
RlzE6+qcut0yzuxOmusZAnvh50bVw3p5qbvFc2ZQ6HpSNjbBqPxyLtvS3JdmouJm
CxrNkItUnwiBTvm5O2ngKiAVSGvb6fMT28QDmHNDZw8KgjD7qvRVjIZUlVlLeUxP
NgRHNOgOZOacw3gR3/RjYb/ctgF9tBL0q+0/UaQoWyfuQ67pwfyYNj5NTVfVQkPm
i8GLvbIEE9oXtm3OU/GvivTo+wW+HS7avdHZlrwtXVNPw/2BQ32I+83oUoauzVsf
CBSQyri4bljZ2mtkmXSsIrSHldUu/JQ603iH9JVP3vwLwwuSl37RhyDILIUXROWe
rLm+QMVXIru3igTfXh5MOPYnsOmTKIlVB5rI8KxS5510pknOb4hfQ9VofeQ4x3ul
N4om8LU6h0y6DYabE/yMVUeqWO8ZyYdCEfMsN9hihfSjl5QeWHIhyJ9CfOS/SrM7
XMgKRJGFqRIz+9WJtd06vbkpK/2+puG93jf/75AZUbYurEm9vLdbWbKkLuP6XCJB
JDa6B3b0+0bxQ5748k4td7cmlEZAcx1NSxvblDiNmb2VJ4GdFR6Nry5idwcqE41D
lWUoRmQ3Ou5AgHdD69waGyI03O2uf+PSvRmyYysaCTmWgSxXGRm4UmcKfhB9OWI5
ab814Idbu4fR7UxmFl5iiHkKg8xFUXD2bYcSbSiuz/jHt35/E5vp+sMqsM1gRjC1
ur/xYYWSPfc8LnSXQ/xOsoqsjyfVwvrIhMArWuMTv82hCTKP5w9YcwSm5PM1yjCD
4SX+ZQx+iOHZynbUWg1N9CpJEWAbkeI+UGgsEZmGHupEto1eLjjaI1SUe0HK87dn
UfHiU0nC2141ChknKF4W/a+mFPplIGTz4RqG8j+a48AIbjWT7l6cAI+IItPOfrol
Glra5LA3ASiBCxkNztUrA9ql3L0blTbBRHLXD1k5xlYOZnBiAidX3xdbpEizqkyN
2GblTr3JvqBcSHUI60yeN7Z3xPn53/6ZyQjK+bWkYupZszouNYi/FLKVD+tS5d3W
X5rmYcIe344/whpY592ZYrZRVh+by06IPl7T1TcDVp/g0J3JRkgCOe2iSpxaP4O2
WYnqFXohZHl7v/y4wFlrpZXOUW4otu/VWweFwqaniapfB1DTY71tIihFxc063dz7
r0M0h/CLoKEQVmJMHoiRNsTuffzrCuy8tTSOMM19bGeXi7ZV8ivd34QAC6zMi7/e
6ryYJV4pgrL/YuYysfS7e5gnW+etGn4WbZHie1DJeIXdEttM2bHfeXP90psnh0qP
f4aCL2zcnY3zHx8ktW9TckywOYD5MUqoKubbhPYhNPEnlE/Z03i6w6lXlyQ5WN11
DEW4JHp3wl5QoQ9AtP+1PnYXkhseiP2S3PJNVPro68mdR85JOks0AXvV2jHwaQPP
ddVOVKF0DeXmZE81MXqAM4hN2wYYDjn2WgXBe8HzjcZ3xH0jAHa5w/p7s76yIUiP
RRutKG9PPmACJ8ZDWkgHedGGCbzeCIchirBY63hrz7vqTZSxuSyxRicHaFdqpx/j
gUNHz0phvFgPmlbCoRvjGA6p45It3gZp6Pe3WDfb0fNE+hcCPeRfeIVrFim2e88m
bC7F1yGSY+KzsobrMKiAIrGb4OjUhwLLbwLAHLFYM5J5OgxecHB6jypyatDxmeYb
HGV6Kz5bRqkAmS/mUMbPo2eCtbCCkz96NmNQI79kyWcZs+Ls3nYDr9jIqQj+ZksJ
dE+dURFOAZHpn4pckvGcWWX2zQZT+PXuW76w+VbD8k8p+pCx9q1eg13pHfZR7Z8H
K9TkLpifdjrxoaYGeJseDdO7LFwEn4J/Bzjda4FrgA2qkAY6ncPTmoNJNaY/5C6K
6l8ngHamsqQSuzxLbjCfw/ToxNuAOYqjeDbaZ39VjD4QNoY3ndVmlkImhMzrmJ7Q
df9RQMdAxYAuyHBLYo0DsMUxon+NdbG+MailzFPxKD65Jt0IdRPSNHwe43rAbi0n
bm1ly+XkJTLrMiYeyb8w6m5BjZX9/H5Ivjjf5d7fmUCCDz9Zo1YFV2KHB9r1YI+O
zdEXyyg22o2EIjnlmBvAvNk7odAbmBjn3giV/bbts9lXfm+o7Z+7R+oXjy/B+HrP
BaMpzH8tpimu9/yrpkgk3legPnU37SjDKowL4HQs4Ic82PDDYvV4XcSioDqRO6qN
jCeOj3TEBXG4TIzRlEq7K/ZKzJ13icgO1BDFaxZxkanVsWcwoYwWWWxmKPoRDQ/R
U0yTpUUKmpevRZsfTK62nOg+fvSSPkB2ThmUm+IYjI8lDFBWjhZtTwGSO92neWcU
WtDcXYzT4wJY3+F8GPyXJPX62wOOo7XOMjToluCGcVZjL5vVqc/329YvqyCPgH09
YUmXeqyuCjVBAmNWChoiw2ZCqisOdj/qqUN4wvYc4auEKcaiEVGwceZTCNZGYy74
QlUznPV8GM69Rc/VPRJLsfvRQgSsf5qd1SxREiEeoGB02pRdN7brn5h4do86Ejl7
EOBqgZnQgXWSgNQaDkLJwekyyZ+lmbuWXPt7ti6URoUsZXUvT7myYSAigf5mt+FP
5q0TVMDE15SJVGo90ve5HP71cc93Bg/Hx+o5jb4XR3+GBuujPIX3lkBCVaj3Rr29
kvgLlemjpGZc0QgxMLSRCcI5GHzXnIUjVScFNW1VmtX0n7g62GZn5vB+aXaTtZAG
HmlkqZyqrb8VQ8rTI1JSfhUdYJiowOtIavERrm6llbX+TOOnj1ijW5Hp82b6DjEE
t1LaMrPCW0SVHITC6Ro08HqP+8NXC93Xb9ND1vZRee4ceK/+ywK52rpC+4JOoJ4S
mqIxp4QhmBzvbUHhGSIyzXcdEU45guRYNyl0PlNkfRiEw7pD0BmIqlE2GYmD4/oe
j/6RZWS14SwGxCIQ2FVSPsw12RYdvZkz52AIh7G/BxVjHZv9q8zZGQDhicNl2Ojt
6W3jAQw51lurTCbgfXd6BSRUDJQ6DpxhIAbsPvb37uBQYKO4ZVr4Od5A98xRvgVp
xgEEayQqe/qNoPZ46cAcwZcKjJo4nI1fagXEc2OZ7/CIc2PU1CjJ3Qov7u5BSi0/
dYXq2uVe49FQhMm2+C+gl/k19Wf2OQIf1sjdtChrf1Jk6HIcY5J7wCGQ5j3FQKp/
VpMiB4CQiwidWJ/SNBNm6QyAgFGEePQd2jUPPMRHTMCcMjlodZl7d90NcJowzZ6Z
fsFQd+0kEpG6cIpVquUh45zR8Qe9xBlEUj2R6dXqNvJDRdi/sBTJoHEIkYwb72t9
57ljsPIA4MRBGLEK9wkSBffyEMroj5PsJgGrK1k8189FYIYbaFETUWjqd5tvxZoB
kgSCd1xoLiEoIgui/YNMyeK2xtaYtNYeA8v7jhViah5nvWyB3zI3MpU9DbB+DW3e
up+q6vB4TmgwpedkqcFuo7GCJArnvFk7GtEvFxp0SpMVYgIZVeifYYstjKKylFZ2
nJGtI0tPlqg2nlUBxR6/IUNCxIUxARAVVrrRW+PDgU9P84lfz0+I9P+MIjrYIN/k
Zk3lC92HMUHfYsNoRvgjMQOvPSPKu6dcEpzzKX708EMqm69FftWQTkTzm7Uv+++Q
UU6NQ2nRfF36ivZ/x7ZzrTHoKlTgoLYNHABSJioFZS8QgjWwn3QcBfG9eKa1iP36
bAkOMHdJeY8hl03EJkklHE7yjPrfmMICH6YnVr7PP5eNKvsWrTZminYKKtCiscuD
dhSE58CRS4jI6hbeunDf8ec0s020WJBKBb0DO7TExjGi+kDWPo4gDcmm3h60jFZM
vSbSAS8aMVUkIppe8CNN9AOQ/czsvDDB5iv+eX6NkT9pNEiJkdUlMK8Nbwo/IGkI
rq1HFeHJpeAphSTfwmnQJbZ+3jHqlonsQ+Jr6Z/wSXTMOtMwyiv1kY0xaLBKsSAp
MfP7UjliXjDxtQrADQGCON3SGon4kpFtdpk0y6fGkeuDqsHCO9LnN2Y9KliQ63vw
zL3GSD+ZbaclClGMk4VNEKkhXTcGG5ub1Ev1l542rVn4dFuUZEOUdYBDKu6uIRDf
rA3zpJvfWkjEbaBtpbHiQsJEpxEpB0GvnCRz2U5jEW46t62XiLPzqzHaakrl2dsH
+XF91tODQsFQJVhXUBmp7dQwdH0N2qbQt6mcqP4HnDgT/451Drd5SsCol7YIsOB2
YF25AeDfAqf4TzXJRpl9zYRoZ+DOtV/FCq6/gdOhfS/SRfBeg2Mvgd/9qGHrTHcT
6nraFNZZSk8MSxrtrB4qu+ZE0LPHrOx4+OxglH1E6d8QwDGFAbXz1+T2Y3PiNQ6H
gXwO0CYs0bmN2Um3E2IBdD6JI4PhsgSbYguC8gVHjhge3isjoOr4lUnZ6yzaZ/QQ
6WlUrxBZWRF/zuggETXRjXyjblMHOH4tDjfOSU8IJR2z4+vzkaBDY8L/teBOO8VQ
Rp29Bk7rrLRiL6tC7k9KLXMZ8e3RzBWBWbOstK1vOGEPFU5++UkSo3SyqkuiwP8l
2PentehZlAxCX9tLH9ckAZM9YCLJWF14QjeMnx5wRY2WG3RyywyhnjyOQ/wkt9ae
DTrxzZK4tMFtg/YbbXNAJD2UxXVHSS3ZD4lsgxnlM5fFpaWgelcr3Pm05G3wBOWz
Om6NGycQpVRMR1I3mx/aD17zh4c6iPWHbUeeMDQLx/oACWPknAJnmrgD+CFzHwFv
9Miuui9P7cxE7MS/aQBag+Ey2LkavSH/sBvTjHNOEXlSaClhdIHcQiFAS09W3RdM
Ca/Nk7vrSnosAXYBKPoI8U4Xv4Yu6sSUR98yvK02+aIThYRaWJ50JvzOL4Imt9sg
llIQYYEZf8oH6CMD9MZH0EjY9hLMdgaOsj7jelQIsgjENJdt0CQ9P38yDre+1gHH
3r+vyODs9ynkm1Dw2O4k+LUElgF9uiIR4s7FexaVibNsyxkkyrQKrrTgSwDbtNts
1RtGJ6Z9cYA7k3Z1tKxrH5ioiFF21o0A338lYNhmosr6sKGoIyXmhgkf4Ld/0UgJ
G+eFHy9i7tKx8v6oG4MUFJeNuN3vAgSKDtQ7M3DkVBRBy4+15R3iXi4FKumP9CSw
1BeQFjJDHIcv5fIrROdarAkQOuPJ6EB5KMlVB4ze/juqQZm+785yUQAaGp4YrwpU
zYD2STHUqTSUd3gywwjyLeMG8OOX4pe1Osh8qW1V8NSNc5KpznPkxJPSTn7VnK6z
YnW17L0hgLefwJKeFf4fnSkrDqI66HpMHzmP+3pcfFROM9+e5yrHxCy7vE+PVa+u
nwf4M8KUNhRO2A40H1aRR1YGIb7WOQgm1IvYFE6eyIq2gloSqPU9iutFyPRGWfea
SI9jaQ+/+2pKV9qsUgCRHD0sI6IsuzDzNrD/meeNB1Eel9Dd/EqGApGdi6gkgNwa
fLzKFIk7Zh9FupG9B4Rsp3x+0osQ/1F/PW+ZypjJWiGI8egyQUt9f3i6fR/IsUeN
lsNY24Q3A76dFXXkfqcBxGDkHbGVghxfyoLsXqrNgVuXs3aK/5U6uLN7uXYED3PS
6J/ZyjX/lC5R4buohLGD1YZRQcYSxFaRqWfnPLHqecyVGa0XRLoGkBxawuRtHVFX
hSKjL26aEW7hyJmIZS4xSW8rxoKMAYnAADI64A961pO66D8ZVIvjbIdVusAwyllE
aVgVuxijNWHXK6vlxQ73+JdxYHSuzrYjL2YF7cn3t6QPqEWcBhEP6OFSZ/ZVwVVj
xxGGA5ymgj2hCdB1SB+YMh1gvgZBi9QyCyJLCMpKNxXkzRUhYFSpMMFRlQrTT837
bOeob3QT8bGLL1IZq+jmWdl9CNWWy/PSmv1wO7QCxSdlqpcMYHgEKnWrtRBZ1tuW
bM1Of6Q70AUuUeGjRSdh0xAops9tglCS8TLbfazhMZKGCrSNmKjXnlzP9mOCMov2
t23PZEa4A7mwf71d2/agaAXbbY5iIQ8QCzFs6KuwhqF0emneqdSSzrFYLaRXy95g
wmmnJ33C1Yl8UxQ35v9fE/KrGP/KPdfd63sEl5l7MLzYwvACgQDHvH1JzG6Ep9HC
oxSwTjSY3zXTSC+jN8QUT+jLY6BlGecO1M+nZbyTxBkth8xt3ARGtMLfx6x/82Ok
dfXSzCVNjLNpgVrKyLKBExmsVO2bhlw1a//ZAlE46uCcEIeLNVVxjVToHerQ6w8D
GB/VApUvDlyHPUIAWni2bgODCeFzZTJ2xxPVEiQB6olb7biqny8SEilCOrMkfpuv
i7yis0qCB1IgOc4v0CCDtbWidSQlkT0Ybvf/5DxOA6V90goCRspIbU/rZOdUn31P
BmgE17q3ctVapB/97lVg2GugFl18My29NQ24+B4QO0XHwGwWCZK2AIAXihqAghzN
5orwvi+tWFNUVTvlIk+sP4mYXlRfe7AXF/G0A42N6B9tpIppLqJgflXTVRq1+t3e
fbDU2FJPW1W1mQ+mpqrJ3JYkaRWOQ7+QiUX8LYbyIl4q7c0mg5n2FOmp0rsYw5h7
L5KjxGTE0UIvFZTjze1IfNlz+qN3Ek3dgvG4aYBYBFw85IwigqvUclunIoPUM68k
qTIkW6bulOCI3Eq0tdcoNGOPNbp20QNZMrZdZOo1Lj4lH9RU5Qwmgh9PWGHdfcx7
idmCNHoHf1pS5UFPcru1gRuEdQZmRlMXWgt8rzVf9J/hmkRYKBnr2vDzLpCTPWrd
beaNDf3xvT1oV63sSjg5PRs+XWxIJEx2yq4qSMJGNavPKQVJeDCzXDsFxzPqLmS4
DvqXHyxofTBI7ylKAzTEiT4g3Y7oe+IawjiNw3pVNNDIrKTQPxjEw+Q3uWnPKn+q
LXrg2jx5FFaOtr/b0xD/IMpXiVz+Wt1jn60arncgWypNwloFjOuTMhUVaZeFny8E
IYyuCp5pDDST7UnNn4o18XKUuX0h/qRVSgrNLCIxyDVxgIHDPwKN1mxcy4lnL8lT
6yJWvplrO/x64zOvBC6HBQI6VMzZTA4wwPVMg+LSWaOqufY4f02dc5hL4gt9Pwb3
dk01cjrjkIHEs8b3NMMSQqqkGw1+0RuTRC0PX6CGDWEAT9cyiTrSfHDH3VOUVOo+
KdPAOMd4wm7wsrYL+zVdmOWqadh062PUNg0Jg3nctkNQTW4Bt1c6ginwldgeNeDP
0CCUs3oAyQLjOc5OYF8B17Ai9uIyDUJ0nnlZo0zPPnd8paOtSIstddHC8QhaEIgj
iOelMo041jO/GIUTLTXVZ4bp5pTBRDbRkBwGXBNDuDRSb+6y2vAKo11ecQnhM8Xg
Q3NLKHvUTzOCdW3zwIEQui0YwSXs5FBB2wtd5UdOHmK5uIfEkFYdMcjVIk5pRg0V
H43u1xnB+dBmT+XtJRyiNHYlzUVWXLS3xn4Z3PM7PMF0Tkfiqpe33sfb64h9voGw
Sbw8XtqlqR+ZgaPW6OOtPYg1XF3AouKW2um7hMgY8IL9VBtZH31x8vVlB37hOyBz
cU6dKGa0nbPXDdZO997cYzy0lQVK2kjy+8NZ3GIpnTbLs/mM+IsNB5HNRl9XLVNJ
UtUZsDcfAShc8sOI4tGtY9C4wAbU/hZdPBXzDcYR7xs/uGQO+EATcN0FQ44nPswI
fc9VDKU24Bm8sPQ2sFRykU87ndg2X09v1QsHVLeLp/Mdq6nnNoMGPSpmJtPezKDb
tTnSBJmzLS9BwEl3sQ8KSlSxTM8phcR1K0bcvBtQ/WE3YHmQxbUXHjKq8/sODJt6
jg8SKPOuCwGMDBdadgYlaJYxAZnjNM85m/e77M3oBz2ohXExk66tAur65ZHklXAm
sh2JOUmMTLUAK4zjgnvCiji/KG8sIQ1VhO4CXJ1gzT1iZGwHmNaqNtZMNzEQA7pP
eYvWgGpCHdOQXpjSCyz0v+7neOihPnUNO9spI1kjtQTgKK+oKispNIa17SdWKobS
IDDgQwp+jhTQNgCtMhmT8LfKTvGhC64hfFK8ZVaD+Q3X1jevgJjRwKBeP7eh11yS
LIT5D1uPdg6KiMSzNYCtmBchnSYYKLE6ZNHAqF62rVC8qVU9OK+k+eaZvLhiqLVp
vqsmxYobQ2B7uEGwTcBUZBLKP4OmgAJNbLvYdx0HKwyGGhjp3V2hB5b6DHtaMO3y
2rIpsMizuOSap0Y5bJSwWjVDMM60Xn6NZGD7rU75Yybg70IQO1ayOJ6xjUD2rUVR
I7vKyxh+JGgq4EiYK6soaa2Gpjlh69xsaRRP5PMhsFzoHFHWpWmM8e+i4kfgZJL8
ba2ApDyYo6i84dHwJrYtzUeH8J3oK/XHdzDDaxaMRJJkidfj3ipI3dzz+wsnS7V9
X6jeMkAgGzBg/QF9sNN2fQWmhpnprAdlwsKVBo7KCMDLL8wvR99k2iGCYQ7FQ41c
E9EpBgkTK1uP5f7j4wt3przZ42QrsuBJKpvBtf0G5K/fp9SYSzsN9wtX2Lp1Xg+H
VCBlYYk2zN9bq+MRY75EDH7tYHPA1DWgxD9EhptuV4ISwArLsAtD6nlR7FUCEP4y
P2R6uN3HuVO+gIesEO/Idc7r4djprt2C/JZ94DkfBJnDAYjMYfBILSaTZI13lYp5
r3S6lriLw4J9Ph62NNHdjWhJBOHEGaE8q/H7OLbyotx/o/DqktYUt1yBCFPoGHFw
o3AjChIklYOlo2O/b18n68142Ik/+HmTKGLmesH/i3fE3vZs8FsKWxIgwxQ4YSUy
ABD7UjwYlE/E7GAX+wdBAp5uO9ILb1+1nOpkrUIt+a2j328P4adaI/rVIhEZ6drw
m+20iuAkzG99UnxdMpiD8yA1pRTXy91pLOYb4ra1nB0ZjSvKtfDL+BW9VdA4tdpQ
n9AK+2fzojW25nhDQ/A2mtL4FY5wBG5mO7XAT05c8P35sOPjLYay9xaj8oOJhDEE
LY56cyDt1Efb/+SFClCR0y7p6LcH3fZvQdFrhheNfpgmByDKejkn0BwOCAU5Vx3n
SfjNOn1+vsBEUKgfStdoA0r6ROOoIjfhAvkrESG5xEAEAoOLgGAT72LVsLhyw5NY
3zBZfBeMCMu4PVEGc9Y3RlpRLervebUN2HJo//7Aipv+kFbPa60s1MfoelV6t+CO
PDn//XO/Lg3r891WRRnHWqbNNrYTzk0MVnfMQC9aqgTMXLIsHX1M2L2F94T/71vv
IPIkSv10t/d88F8rcB2pkoTL/r+84PLIWwCmb0G7SFMpDnO7O3TuXjyaLiRAe9Ut
f4Xp2E9ftsjQfW5PLmPfsc1NvNb+irKTGAZDFX+2l5M/0qF81W21IhEw67AMiOEV
mfKhvvMpLyOJS6ouG/I4beBMbWY2R/j7F0DIzaei2grnCDdDlYefbVs7BQSEWVGH
jM5Y2IEDNZxhoNSIEqH48CLorE/gWdpWVoclr7Zz+Yt15QpqL77KH8VPkRzeatga
pKlmD1rpbqRjKpLsoE4s/w0Txx29QsMfXygGAMptiJ7iZX5PhbM50EVSojR9vsXX
6L6tUyJYHv8GttWrganWz3A9cgRjXpAliB2tcWHNEEgVd2QSW4EfaFDOQfHol668
W6oerXxiBV8iLH5LbtF1YpFPe32n01GmTnuaDKZZ7Zp1n/PPHhM3LiIOAnaIo+l/
U9a3YsycZnGT7tuuYavlFfKaQfOMavXT0DJraHPzW7ND2U8dd3bTn8UstFYINEAY
AN2mwb56rRdRS/ipeHYv8H/5KvOWVvLNi60+7V0k1QH/QdzHKRSmKaWby7D7FvmD
G9uDmSIYVWRHUKLuJi0Pw+cxw21+92NqE+10uE5U7aQKoBAmQNgCNKjY2mRDW36i
nzt5xS4xZYgqE8V7ETsROhgDJiYbous3VpMtMgMbMuU9M3qfLobq1LlWh3S78A2V
3f/S9jHPhU3lcHIDMUwEC14aXTnxqd7dg8oANuk1GhWKWKBd3FdrL4/5Twtjpbsw
T2vy/SmzUUeeaE9vfGVK/vXpfCSVu92fMfObOmTUc2us9RrLNORQK8A7vUFZli//
Pp1qKKohQL6zmkiHBAE/2hWovIZqXLmOMOxbRrx/tKqW0hnS/qNaiBNyToY8qu6+
gmXDinzOq2YThncq4AjWRHp7MZm0B807uG+HDNabCJv8TOYXL9vgEs2du+7dXOkm
JIJsCl08a/JiuwVtHj84h4/h0vqNameS1KvaOk5FCOx+80bg/K+ekQWpmUC97+UA
eqlkmxu20KTkB94Mk3AmDt9kvd9baOROMc09TC02IRyoCyZvo/+WmVTZffOtPqNo
uDtrFxlidiTUD63YD8D/HrIYu0Rc9HMBInvqT1DG5Wj0CSkcofbriGTUkOJqwwW2
n0rtFW7KY4VSDrKxCB6Qq9PV7nzrKPCz2yzLhdz+Jy9Hhk6MGvT1Q/NsMDY5W5SR
iWE+6yZWjn2lkPh+aXvkDtuPwDhNiEMzANNaP3g3zM+T2OD1yYWQ9RQ6Wcimig7D
eDHGUpnBNiN+2vA04VuOUks6WFQNp75Ldp1PZw+76M/TIuK3TsfB03KhjkhSZ7CB
WGxTZw1uLqVJ7BVouQdw486MDJRd2TBnyMbUh2hQy+XMzdXrFM4tQe32OqLildpQ
Yha6+02tNKZQOFgcR+jsINfb4pqLiYv+9aiqKUxD9qVtrfDAsfwrekzyuya/MRdr
dMSH3ut75AAKln8aevg0MHaNgJjKxVrAuoRyZ18oytF+o/ya8N/SvY0UxWYnYE4G
hQ3jHJIky1m0MfKRd9Fe3Y8ZnmLJbmvuC/20PoTvYqNgSvfk4tsmB93V6uAxf5HE
0R+wwGx1trz3Bf2eVKgu+t6hGr1eVbcnfK+WZ7e8VtTMxiGgFjVj3nANgmHZqZk0
8Th1wkJGMju1T1w/LG81sewvn1Pq6JRe76yrrmnnlByDyHrixPKq2xmuCm0K2z9m
P5MukiXR6DIYH9jx68bgLApjX9B1B7Q1DsLtxKWnvTl7nv33YUGBOzuWo2tbuzbZ
iXcgPrBrbsovSlITdDZFztKK65t8d3pXHlfjV4sT4htsGx79sPNTjWFFtlXAWkfB
Qy5kANQt6DDg8B8E9NFLY/SAk6q/CfLV7LG0ArJkQNSTSUcsI4bDq3X+L8v/vTYS
/S48GPnMI+5OFt8YtX1noOYoxsEjq3Itg1aC9KQVRHnlt7lc4AxyQmzxR6fIu5eJ
N8G/fQa2Yvi466GmuCDdTty/smNkBTBAgNOluQndC5/t4Hc+wwxfAfUDFLYvzJkm
l/OmA2r8MoBOc5BzxLLSAbxQ2HcMO4/ByvcRhDpK3ujIQMPJ3ugLoprzcU4uKbhB
N648XiSR4CIA7kRA4aVhxdBSfu4PqaT58lLpxoFNIzzFZi4ThsxSukkhAUy5Lu7c
ZbkQra+0YdFnmmHXezdPt6nsPXsJOopoiR04j//MRlq9CKtB0ZO8MT7L1IVuxsOv
K4DF6UxnvtlojNHslzChIVjgHz3BzR+AS819iEFP/T0V16s2vHRrc2eMCnPia+/c
8b/CbfFX+sI4P+6lQkAD0cWyI/OkOXF0d9ogxnOKoa20DxLTfqk5jE2fTgTMHsrv
DE7mDQqsewc1bHSmJymRGsjNQGmSyxfiHETx3+KaEzju/nqL2cV5mNKy1dTPAwRi
P+EVjzbArhhc1Gu0g8vYOOkEnZO4SCxTy+uay+b/e//kI7odNkst8H0y8YAMloep
dicz7zKX0COseGsOUG4onSOasYkL/4GluuXLrFGnotsxbi0G7+TWPy2ceD6uYBs0
zQ/bgOXsVKCPxy7OOLHqBHPRfkfCn/1Mc4i6JY7VJkXYzmRYB7IPSQqPHHrgo9Bd
4A3QF48YNBorw6EvVXzQvISufKKZSJyF42q6jfmYmIr3kpC42Y16Uw9V8ZhvQgL5
/HduSfLS2/FpEXnO/V19w46G8qd+RLPThPwFSDkIYTvl0oTz/gACFRBuSi9XGPQ2
8mubzRdk7uUkUNfGWhd8kLJHu74b1KzkYYPD1huOwoEfbG9vAUgYGziQZ7RuvlPq
faD1aGmZGROcOghkaTlnj6vBhICAsgQKtfFzeDXQb2OQAekmOgXswTMz4ormdOWP
cpgcm6VnXCiV49v5AZvtqAG6FF0LHvDMy/UKP3hEW6WRMC3N/+4MnMLRcc+tOHNb
ljDEqnjCvozRskHX/Sbd3519TnW9unjSZZpLBHqvEjbNOj1V3skwx2OqWMhPNbZC
Q+RbbXIh1NkvAhvV85IvmQVzkqhRlatPfNbYEPx84JKl0/FPjTUmz2nTqP6s7Aff
PSsDBwieAkLxfHvRZakLB8y5+tAV6Bo2TilZ+66aQYZ1AN8AG2X20z0ndUSoMQDM
oJUVjfT553VAr67Xdvp9ckvP7qP5qXPcrGX/D7pc4jD/G3b1D/Wr/hqLCy/gb4l9
bRpsH6wn85Q40LO+sV2zaIAgw1C/LcGcXK0RVSkMmfsnl4B7y7Ca6NmyXiAAo4dB
YsTFVhewzTGRkUylKsNfc72N5yUen9QhSmhhtSEbIBJh+Z8lHxKUAvW9HtLrOgkA
PomozHk4q5OfDd5K6mh5KgfNweBI1CAAywBDJrnQOx4Ia9p8XrcgXqGrqUt7wJ4m
47ld6asmIXzuqxZDm33/CI6d+652dHUjkwJF04wWK17diwIH20yrkR5+jmm+dXZ0
CLh5TTVGoYmUthsuII6fz1JvW9nN41ifRh+M8KJHNvt/HaPvkMvc3MhVnuxddUfK
NgS17FFqLFtZ7e25B95qF8r67k6ZbTcTElI91GYMEvpIDCqMd0q6cPO9xgzLishF
FI8fAEzFd8M1yyqfcautIJ13vm7L1+y9itg67tZf6Y+ZDhA1KRPs36oHiA0X7G++
Crg4JI2RXy4Y1tL9boPnODFcw9r+/gUXV0K8gG1trhuqQDqrDPAIlRfPwVH+X3jv
7FJSdpgnvmwvnDZWs+Tatf0+2W4NyxL/59YNbzIaaXfkswRIP7qK1mrSL/b7jYDd
Hr6ZoMPV6RkgMqUxiPLpzdMvIgZ423X0/vBspAl1qICJ5cIdx1y/yroa4PeOqgXY
WLE499DppAafHGEKEChXx2rymTQUpbBAxz7ohmbxQhd6nO7M9l9NsaAJDlLSJEWb
jfAsZE0YP/+fMSI9BQ9CECfaEcASujHcXoeg8I7ESiNAoMlT9QTU3yXXo8twlJ46
SCm83V4VveDH5u0ogf7WtVHA5eDAwvhp71u9yO8kNd74Rl4B83byoxj8m8rHH63V
LbLGl8zmsoNJtNeWKz0/mh/fYCKWa3jzbR2cHRME2mqDtdheKe2++1/j2AZ/ELji
DcKrVeDq8lNqF7NCu72wGOJHH75r2NSnSBP8dde6Z/7RDadE6+jpdQ3QVkFXHykE
ysgvq356BPiIBZhg4SyMJz6Zxc7Au9YDmumKZmrwbu5jyxOQWN5kYrS+dJJl/UTu
uBG/QIMZjvzx6lAxJM9YOV4K9k1ZCZeBythZycegWRirQKF4uPEpJA0CURM+6cE8
tJPaGj9lMgLnWxttInTWzDkHtqrNuNs0PnKYTQCWmgJnuJ+2JRoJBJ+o5PfLuqBH
9LsTDXRJie1Z97s9S1Pb2yTyVqMSGdnmS9+mOW+gQlyr0esbRLT0rVXnDofZHNXf
GD2T4hPkVtwfFg8jx0uGe2tZMJ7lOy4fkCTRBSucfNSRA/vLbU8+ZmSGeApYAsFH
voa766IYiY5gkm0OxGxCOVOQYGmY67P4/B9YhwuOa4vSZGP/1KBVGc1pPXTGTShu
9lLmEwP9xSpt+dPjbEN78rnMl6NUcFjYYhIQvG5gc2vRT/99hE5QV5srRnHrJlp6
uuFpumjd2ug83t2D56AzhEwFp8qAgzb91lU4v5V2N1KpbyzDKi1WDpABTwg8/l4v
VMIgq7byIamg87bBKd74UXIOulnfUcIGlfeopyFAJCywh6FAgUKUx9SwYBH0n76n
nk3MmyBlygOYOoESzsOTsgiwUvaMZK3xFp92LgUxXbDut14mWGQO0xklcETMOTxu
hYHWDut7hmodD2FLUQyCaR4vuUPU2Jfq+o7IccIdQc0m07bQH8mkk7HgAZv0L5c0
JR+RhUxi7wHN7kyUe1XBw9LGI9kfDnnBBGCY67MSUQcH7XjCpJy/YMQHkm2L9E0K
FCwCXhycqsNyGvt1agsTEMHBIxsblOn2Zsskn+POCoY7DudKauQ/Gf6slexZSKq6
2cUEnj6M/epl+7If60oDJCPZn9tZduCA35fjfujdtSgJ5hvvhtn3LRo9kLOnDxAt
UcWDgBrSreoCXPMRtyiEHxtd/5TqJy7e28O+jLUVrSbjy4ZcVpuwBf5qwWD87QYU
PUIj2dG+Iwtmj/gYbmNQVVY3XYHKt+J6gk8/WBGAfW60/VOlUzeCKuxEpXiYcZIw
qi9LENa2Vn0TjpuoNpx5Kvg0QaytGcvfUEZrnpHVm5yce7UiA2uuuM1QaVkptBqC
WG0jYOPPxVLceW89zklFOtbfouCiZs+dH76y63nkahmR5uOC0Sofw6Gx9l7/7RvR
5F2/o09sLIcxXmZ4G7/7BEaBXKKKBIa2K0+4PUKQSaqmm1qFYtSnaARywlYlzV0q
E3dXkVgsBVf2UYXjhZBdn9eP12AN+/1n75dV26y3FVSlArsk5kt0nBdj6yeqR+F7
ddPZC8CiExa2PU5YPfQwSlstHc6G0MuUkP8IHXFdBmOMupTnZwwQdH9FD68vUWMu
vIawlTekBPW8vvCMmWvboPKMou3MqM2gMmkJhpt+WveGiApQsW4DwSrV6OWcvpt4
XjICKPAUSMg4W5UP1+fB2M6qQNBRXeayuXrPd5KNOt4xbPcafywVoHI1zLpl40Pp
iIwQtdSyw8BCz3a+uNDf3DJcYoZQ16DCfxNLlJXsQ9xP4R2DT70KOvwWdqdFlLOn
21HT9vhcGOvrdN1MgRv0Soi0cmyrzZnxw8QTM5+VjoXuto0CCU+veYFF/4gTzIwo
ABOE2KjgEfVWkHV8d6UKb3Xh8cmk3liwov0rUfKIEhUwUVPHijfmujZQMpG13KhM
1fxJDtp/JPw5F7XQB+XryDSSW9M9zKukxo3ws64E0I/7AO46e2PLyyM46ATIDLE2
ZWZxtLvJrpwLIgye8QO9HdAjMl0srEDrwhDMM0jw0brlH7sWSaCPgJaEtLXmkhOb
K8iQJ0eOod1vAFiqii2XGQS1927XIlUcz9oTnVmCNjxU6VhJEASEpCKd/C+f+OmD
9B49h8i75bPveQQr/wI548mOR5sTyiqSQCQBZBBPKNPSxY/q3+B4YiGqQs9ELYzw
CP7bCFrnKUR46CACsRDPu9JnovQSytIms6M0l7YYOKbzExJ9lU9/pPLqQa8erEOT
8PmvQ5wsKl+2FKYwLEMUx4jnl0BS70MCiJ6nwalpAELxWRUCl+xDIXcsce+qPKIt
MXQAEiWNkV89dmQAeFPJh+3pfUGfrh2YuHdasjfYOwubOKA+p7yazJEoeSuK9e3L
nMm3WAmBlSA9dhEl4GtmCQ/a6UyG573SoG0/7WTLAkGaavE5kVz5ugut8AeyDpc3
MgaLB0l4/YnzA0mEdNwIe0w5zm2Sj3TtlPH+kDwYHrhiMzeBYtFcUZtX99MlQb3T
nvVHvkCoTlVrTTQMtRsKCbhpIfj1wfMVeZG3LKmz/RLYCAkKd+f2G+Xk0TlmASfh
zQGFNt1UQCTZJF3aKwV6mR0EeCVsy6M8CI/lb7x5DNXmaWJjxRqL5iPzY/KSbZRW
7l5kVGnJxY858WwCvFiZ0jBgod3wBvpj2ABuLBWn+5z2lQCqXQQR7pInNN4+b8Fa
kPFAVnjuVwrCCvbJG9uUQZJSRNgTujgYvFkgTlZq59GNYHm0YlpeHq4eQRd2zN8j
c3/C6FfIrjfbDuoTCJAwfCQRZT0MslvFbLHLPKgEYPTNcwyodzBwRsz6+U/2uVdi
EO+kQDdpKhCntMPzsq+kDPWGJrMH5KGTdwpYKAzdgqXiXXIfObA1eEz7UWgTVoPA
uZMpcyg/WKN6ypLTbGpK4J0tPM0aI4z7Kf9sgX3JnM8Gfk+MNJFV14AKS1J13M4D
bl51Kx82jzk1s8XZPteV7eWQtIs67aoZ4sqN2DLoat89RiEiIRGIG9Hipdfo3UgF
vIk+F6etVNSYn26qVTQ4w9CmJ0jiu5FYs+1mgPo12dNj+1SYSPZani7UijcUIx5D
hQqHGIGPMBZzMT4/NDDEYaQF/fwkjzHI/BnPVRSjXE/WNvztKnEMu2uYo9v9gLlp
KpH8ptDwbxAdZKrOwSMsXqUv9dFJlJtjRGCkzPCUiT+Bs4xmzCc16R+2u+2nzhm9
q7VbOg3BJrMNEqXUOMlPnjkBozPhV6pd3YAw5ili3VstPp9BEjZScCD5cfZLMsJ5
ESAydZNKWiHwtnN5fYp4QR+ynaS0wOLqay239oOC4b7yzguUkYAkx6l0HK0mG7DI
5rChrbUbWqFbvhu7PaFCIAHpni2GPu9emPeGLR77bnaXKCWIQKjvpdebU8/rJbg8
8x8XHebX6SIhWSyGG1TO79MRbZZF5CZJMjjNKjYV82YlxSpCwKAv6n5Vq52A7Qhn
kCirmpKD+zItx9jW2Kk0YPpHCF5hmKufAh/BheSbweqStLQdK95LIZYvF6D1R2MK
DLSUHMnyWa3+rdMawul/jyW65SYJdra2QCXZBxPLu28CBMPqfNG0tQAFzmV5paCS
tHJSCL9vT8Vg+ydXYH0jo+JBrDK0S9VXhefRBTaUB3jRO0ld0HmIjWi1dorBOFNX
F5FxnR1irodp2Wz/RTYeAOy0sMWSpanHj6m+6cAQiFG9bRyZxL9k7OdfzTPcrP6I
KzY3s3N1TqIH/33JXMbrVNAVJ0gc+bce4DEO/c8xMIN4tjimCZNtTu4SG/meNJj5
3MQ7FANFPr4wkcP/OlUHQUYbEvut0NpLnpxd2a4ztffxPm6rbdIzUltHutexn63E
ypsJXpzkViEEznhAQyFpnMHFEsp/GsY/gqNdVzW+3/Op4a1FNOmynR1mcU0TIq5I
q+H/jA190Rs9gfqe7nuxGRvtCeBpL1JQGKe3R3HxQ0nLGbVKvDcxE9/lOeUQSpKQ
+s8cJP0cY9BgKH0oZNUzVExD0OjcRGSpiitPARATEo/NLyKmyH17u0XvvsNZVPC7
EsXUFDq5XN9kdf2LvHpVv90g+CMsRYHvvo/bNId5PCv0/vnJRL27W7upUUkziBC2
tOUatK5JNa1VTu4GHzqKGqwNzQRrSsvActkHoFJMYnOgTft+cHBSSJDZVGyCABV2
yfVwntcOy4/4XDBkCBBBXnaQZ5pG6xLgU0sycqPYO1tMOODCwwWwwyIwvIxB/RaM
QPzeCoosDNLSfcSI0uOvG7Vf0liEn5xMs7qgkFJY+fetA54DEqDO3FbDMEZzaWnK
qvF2SBRPvJRFVlVl3sUUwZwPmy0kwO7LlrCgEXIzWmWtmgbQ78N87Av0ChwnpdeL
UfJ14plCv/LjOT3nc8GZzBoVwAwq5vv4k4Beyio91GFXq54uew6+D4mElMgEebKp
A3HVAob+KJmJXFoBMN/5B8tTwM78Wj7trSPhqBiCuqNcLVFMiebZOhT+Rjln5ttv
fCtB68+x/xMbHTpHz2kiEjJARJCy7qkceHlcAcB1Jd2guQflE3JMiOqAZ1Zu9IgQ
SWMuiwfjHl4noetRYo2e8X5UPsqs0WSHRtnmYBCrfYxLEQiwOIbHF5QsiNobCUQC
4v55esOw3oj9ZLBrJWkORieiiwpUKxlXYVLjwDngCf9J4yBAd7TQEsfFgig2hGEF
pUbUMa9HeuPsK8dHRH40zjl3UiiwRRN7SL8XPFRWJmU27E9+tYhS2cMzyb/mDvSg
SMS2fYrox/WRD2dByLJ/N3w/QgyEvIlaTj24bXH1dbrYuRYqiOsTS4vGL5D2GRij
Qrf9vemoVbPM2lsFWnz7pxLJX6h55DChT7j6J9KolWYOrnQwgQtfFvMaii7pDldI
DHOGtSmArm0nxfD0WEVIKWSR6LbUN+d+qniTluSuIzRGQFO/UjQSqKDqTVJZqS33
6fdwneZIioSZRF3gAMsS8e6MY+hjnR3y8tkhl7fxc5bLMGhRabQwLD5ZuEfNwjOs
GdchyQ/0UcaXr22yTbk+xDsQng3fc1iyxH+q3kymIBQJ6w0OtZMaTrWL9UTZ4zSy
oYYNYyfV0cjgq+mInLGOuzJLLea8hLHPncjK4BQLbTDrMwXFv2HLWZDMrA/MtnKP
5n4zOs8XZptw3giaiiOl1eFJ916wZ0T66XZ8NB9IcgzIsR0auBNLQfACfxxYXZFQ
7wPApZy9nXbDX+6htc6aHI67Z3ghoWEPQ/JIs2xE6m7oAHHReGAhNQGbaASAQskD
cbmngXLc6ZXVo6nOxwi8ShxnH7nRtw4gI6M2c0tLJmF6i8ol5J4tsN1U1fh++NzU
RluSQ3iGT43139I1ztw11rFmUd/9MvdOnVw9N/CUiDSeBoyzZQkAoKIk23JXp+2C
z2b+QY499O+e2MV/BzMKNrkIHxGAVmdNmKrhpT5hI4vU24/eVJeYfQ8bgy/EXWg3
sY/EZlSxlrJOYcpAmSzwQjLXMZuQrb/SY1lNlnBQdnZ62JOYdSePf7D0wyqTQV7s
L3D3TvztAsJKUHwB8ae7swDMovFz/nrV7Fv/m/V3vK54fCdPJHxJUZHDJxAA7neQ
5LFVMRvuvW+9wXa9h1ldRVBY6WRUxQii9gc8Tdk4wKFwygCuVPOIJB2gXlcQXCSd
aCelZOpGr/tCyDVgYAo8bfLd63niTZrMy+xH7By38r6vB5r+N7k4DOYpdSCRA5I8
LxYcAxoL6Fg2LZpr0XhWUquU+D66EbOa9+VOucUUsmIpXBEV+WPeucHpky6V51hp
zKy3acAuiK8JKwb4zlPB66gZMXJIjXEeQfZ3B0w9HghISV8birwmNwykfGtM9quc
22pN99Of36vTtZwj0FkjIkWQupqmcWeXEwYu8LEPhdufkmEcnYaGGOW6VOTvYQZ/
uSt8Mau3rnEfAzdwRnei8HM9P4fxXnggQqahXtS0+Q2fzbw3S4bsX2U7RmYf1rZX
NmkncOXFHbBXaYDUQQDINYkR1ZfTcnUC2aZqF1WU8h5VCyHgzQ0sgA+7lgl85g2U
Yk/oqBPXDZdeXoiEHuCVseHy+/hi6niX+YT0GAzB0KGg8EQbVh7xYt0pUmob65YW
Ioc2fPSLvY7WMapYPq/2ms5+5yqdtEcfwtIod2rf2xtoIBXONDLnF08PIwMcreQC
t5/8YBMtjgt58DtVNIfR15EYpJybS2dzVL9ifRS2wve643zwtwEQbpKPgREY0STd
7+vfyxu6J7FgdXSyPwPu9Ml3CMtdAx/4+R7jwlGcW/uVXyCdik8r+R7NqKn4//hf
DtNU/gwRMIHIszQsYp7FuVlsjkbGSno5ev0ku6ApO0A9OSXdM899fLJU+sXhmno+
4kjbToVi948MrkDaCxh9vam82mCL/wAZIIYSfy9evTEIL9Vf6U0H1wc4wyDE7uT6
2+lsd40WvIN83u/cuppO7y6KbFceOcr/T4ElzJFbO0G4oXs9Jr8CFRPk6gQc2boR
xkopFMZh1EGE2QNmRi1qFw1UZJXfke/29NJL11da//gnI6XgclZInD0xtnMSgBkQ
eAdarEQ376dDJDLSJZhssSSmcCVupZnVTYiz6speITBRm5k3/xK5SCSn9Webq/uT
2RTyXCd9V5d9Wwbhtyqeg+jj6UR9+uu8C3cwcp0G/QvR6zUrb51vgQN7YgFe7hQT
xrFRTZ+Vhhpcuj32Xvyc9W3ubgWT1hS4VTg+HDXC39Oky+GC4CzqIil35n3tY7yj
+ZphEHpHE5E167AK/GUFbi0IAKwUVWwKNwZpKiKKq64HxlmcNGzH8F+2j2GVpJGV
Llt5Ta6KyV/8wClZP7MyZ5amZMcLOjuM6/wclzzHu0syScnjuHjerbkGsx47EotS
5wjGSFGCslE2dDVkj8bVjoT6USS7Sulcp3990wcI/qaWTp9Rpsv9Mosgw8cUyZ6H
kMXbG7hrxdHW+sLqp6r37zB0ltM/AAlNI8BrVkPlG6S2D2epe37rrZXAG9bHk1fq
blTFF//kL0hK3A/02D9CcE3HtDvAuPIl9dLUYqFN0GtsDaobrSZUglx1VOUiJ1TV
m6WXy+wuaNuGC/Gnhs/slRANOvGBSJRzLBWWeM6XxfaXXPCRMcouf0JHUGSWhdZB
LOflCLl+ck/RtvUAD+FU4RIrBzRpoMtHBlNGeblDoukBQ7ZXhH9/5+aHhHdp6Kug
TZSwsGLoyMFEoDuZ6ra1PhdGQ9kXM5T/U3xeuETjMbG3H83PvoWrQGqN6UT08C0Z
9qtGXu0VfK1V3jgXw63bvK00wYGopvA5bV+KZKuW+wE/CkU3hG6wIsJRdR+gw5K7
pSsIpaGxSRSb/u8f7/jrjSo1osFwtKX1aoxKGETu6jGo6NrLxbOT6e3M8joLjGAu
ATb4pxdgzcCBvm1C+cTd3tfJmJjfjs5zYa45Zf92M8GnAkOOH71Bf5Br8UPslgyf
1vGjZXA3EUAFMRkOqmdFGmQVDAVdRZ2w+YZvW9PRVk6Pczv/EjnE8vxAqH/pgupv
nwKS+FkGzASkF2COVRPOxJIJvEodXl3OTcnIs6vSpkWrXVlUW6ReahttHvjdaKli
CZmAxynz8gxfHZdk4fema0QgDCWaImpYXwzf1Mdau69kMps7J/N3hbR6k4E81bQ5
UvszMrYCmk5w3qk9mF2PFeMJyONP4VM50nLy+4XLl6w+mDzjbtmxYCcdSXjSq8M6
Vcwo+CX5/Soog+Rr1C+Do4VHTBPqE5D7/cJtrtcKAYm4O9saAlkIAN79LNlrHii9
+r2+jDdDmig0pp6ohn0tMrDH40JSpxzF7pK51NZhot5ScEQd8x9MM4/ya8XbGVTK
JoHmnU4HYlKksQxHmn1aXWDW2Px6jz5XMeYTC8iDjynlVom6e1O47VtCTFrlFdyT
t7Y0by5KFkDi6DtfNDJFrt8W0hWp9p0Zqq/F3p/y9R2GAMocik/xXMGjA1PUGKcV
KKvsbR9KXlDPWR/07QgyR0ilNSzu7CN9O5A9KD4nLLdJA4UT1vOpU6E/aGc04KFA
UPzlBEtg8JjXkwnsQrXM+1XU+Sk8sTYn91Ie6/y8/tdfbXY2aQB7qJkxxUEvLBwy
fnXLTb5s/x9qD5cHOiHNmQnDL8w/APJmeAIrVemvz6yniaPDgnQe8A1C0g1xKoIN
ixKHsQPJm3nwSwy8jXwmAnylzbusE5HaI35TYlVTXnJiDzy5RwDPW9a2Qew8/Lmx
pNPVw8SmeEUpeBcU378keSarGqODqngXrm7/MYhl+mSNr4xJ6HY1Mdas5pLavrnt
Gh3F0BuuO6IO2nY2JxsXV9jFdqsqLoQwtfPaIVKqFeFhENkIw9lSxvQi/ob+odGT
HnY77heaskMzC/dHRoGguE+gvXFbtREShspDvzdIasmJ/Xy2tnQQU8PYqKZt/clO
hVecSVfvBzoCeVaxnGxORlbLemJBYqjzfCa+QTcZ/Bv497IqbQB2xxUakpcevrbk
kT74hit3efs9WwRFYYTOjyJRrUWf60CcaVHd0P5ZUYf4dI1vdmloAhY7gf6Af4C7
Ox/Ex9MFHg/m86BW2hkrTpVcHqz1ZKsIfDPHDlUV7HkRczOQxL9/OBo8Q4Otn6vD
3BUoBUvBTfheLLgAg0M5d6UcRLRw28pE7mEzLpcs6UC5GkSAIK6AMp1trPRM7LKn
f1fCnfei45R8x+pErdEGoMXZlzpWVL7CXV+LmkJzULLx/u3XVK5+itEinxlWb8ud
ECMDTzshHWKjutcjQnqO/BiC1kSAODkv1b5V1fWiOLW7qeRcxpn3qWEw0PQo+Lgk
miGoZ7TkSpnL4GlTjW5xhtNdbaouX9Q0AvS5Ie/O7LbCusw2WaCGZmCWx+tynQGr
UIlUJJFeRnbHYiF6T6isvlL9yfW9Lhm6c9pj3dqTzo0aMeVrsXHAxMsaNtZR+j6Y
Ye6Dl+o2JaNhQd0+uWg8O5kmsZI+FrxVgQK80q2xPhNl3DrGx5DNZpKWGAOLbWzT
YSsKvp/IagL0ABHzSbg1pExXsWK315UFJ64EOCz/yifTerxW8/OL7xkz+mCj8Qea
0aY5c3n/Qf/Y/wA8zlBHqs0evJ1f6uTks1t1gVqNbZm73aQTsMMc4rIpkx6x38tx
EmXmDj0H/rlfyVx8qr2bRWYwJeWHCwq5Jo4G7WUlUf976Ul2+YeeGqsl+3QGNgsz
D2B8gJvj4cBfX3eBBSEbuL7GCZD4Wm6TUVMNwperzR26nuuNIlhv6vTuQR+LNJge
vENTBovTcUIGLhum0LarTr9LSIpaQ0EyWsUWIb52zVNUxGa+34Po7pfsrbveZvia
gcB2Jqxqjmru25ko0XlFSVQEnt+Bp9QI7WWiwE9e87vHBFucOKFbt4WBAjNHJmmx
Y3Tp4T7hpzptA99cnfm8wWjlRGKbK+/qIMBMXpPUpFloga/IlD0Z7Dzx7k0jzsaT
+S86/FVGNpGVYm5KDF9Przk9sQeTcxfM04EjxAS2z2fRAKRKuccHyPEged2D2yRV
RYg+gXwp6PdCbcV81am0RVeVj0KVIYDAqm+nFq9x38v+kMhs2qcFZWIUaDd9P5A3
wkGjrAFZfQIwj38ZN2HlM/sp8C6DroptENCAMuewrRmAQzsJN8vHZOLJLuxGzYYG
ykBj1Cw3lsOeJ27gYXckc2jX5g2IUiOPFM8m8n92Bz+VnnSIZep40V8x8Z4MlRto
oTYzLD1aXf2HdZCwODJZe6JLTOknvxBxsk9KWmcMQHGJUfxVd4gpTFendV+hZ6xc
+IR4rmHOWKrCFQFT9tWQtCMJesYuqhvrHjC8CK4dpjM7mc6B7Ws5zaiv4H6Rc2wC
+LAXoK3A3IeoyfKwvcYC3VPR5Xv5CwAak0rkIhBqEype4e7S07YZCCVh0Bz53MIM
1n+x4Lgs3erAqT+g5UwdtegNAgN/nwYg+2RV1BDkvPtKXhoDfrWuFwnrmNwfn8l4
o9nTOz2TN8XLMNGHg7kOJElN+okFAW2MbESuHuVd/UC/G1Iq93v9a4r4fcFJq/dw
KL6cqcUB9EYPTfIWxVicZjx930MPdB0NQ+vGzRyIq0B83OY9XIJpkaMMLCJby41J
WPMM4yG7r6w7wXqRHfcNfhn/aRiE4tzpoX9ZJlTu9aJUV9By6nAT8jtK/r3ZHKRp
JhSjuO746MDh+yigD2L5MGxLS2fQysgAWceAyxcbsiTyIG96KRxnYqwK4nM7B4oB
zW8oowpGNEyThap1FuUCeWjRf90iYCqUAvgFRKknIF/bM0maRMz4LjfuwnckMVlr
tNbI5A8VY0FGOLpQ42Q7dYiqBEHwGBVxB0MMr3mvBJtTZCFtdJWruP/urpj+q7UO
LU0K3v8A6fb7Pbots2l5ycYbBNXaELxzShBpMm2MBDlyTQ/4+sw0CEDG1vb3i2/V
itahPfCEmTKa6uidSuhWlRfqyEUXQyDFtA7V1kEwJmuaZbNWcvYEBif5f6l5k+iP
1NkqRyVFg+jzVtTxt/9t0hq8ckQm0uOJkmvOQIsvQQoiDNoVaRieMU72GPJ3hAm/
wCyRVKYrYBEfMHfTXEJkYx1kJ5dgCWEBBpkVzX6sWb8/Pw6N8/2oqq2V+e1PY3ru
tQvczNTmFyF1rVToYb1ig02BiVQ+2YSc2d8CqKsgk1IB0n5cCJmXk34qkJeHYqcL
9iSyt3fspaBBCo28VvyPqd+WFBu7QOuaS741FRwwseAcyELXSF55u45cUwUeGi2e
H9SKl5vqYXWtiSEm9gQpSammpTZLtCfBX0l/FBvXs49843/XGOVkuqJ2rps+QOft
xF/zTZiy+/STz/xyCLVe+eJyqhrXcD7Apq75NYm+nf8UQm50wBBlEe0gl/gB+/7M
lRvNJbxEeYjwly0aXhNBKFqDbErGJaBtSUaz9SifD4CDu3a5C/fBokcMLZXwzrJU
JdUQSOQ05TIBAWE8opCURF/NFmQT69Ng28ry6IE97KtzmIv1HHfmGzxLzreyQ8cP
TM7PsiOsVLmCPKChgMh1F4Nda7IO9ff2K775eI+9I2g/wtdBR0FITdyJS1SdmBf+
MdWFS6HcuVOjeh7+VbcLrsMj3LFLw5LlX8a6HFytxGejIne2R/bV3Bu7w7MyHdRE
YcZ3shZFppmO/u+Y+OOlYdN+EEi5WfD0hSJfqOdSlt1elIUwB6p7tgHVnOnypn0/
MUXng1tfGStRg90/4xN7g8kibaRvyrjWrs/KXi0Cv4Yj0QTVmvkUMf9+TZjbhiGs
toduy4slM1/sRd7HdIYTx/s5BIcHGZqEbfD24AL9ebc2Mxwrt601Qme5Pn8zeZwS
/ZDI6ZMFh1aMLnDF44nC8SogDH8EmDIC/NSZ2/wsy0DOryKfP9Si1AzOjXh0erA7
pXHoY+RH2Y/WulIJUf4vh3LJDhHWZfMJFNU93e8tvsJoNHR95h3N3kjFHqNqeY0V
7RThs2DhU5GPegDXsa5YAwAvac1g7VhDblVpf7xZbxQYIzECWauGfzszvSSeZp/B
3QQ9haS19sDZ8kZxv3mGKQdl1JUblXaNuFlCFKlQdZ+OWiczzD/pcTnnjM2mUQSz
DzGMH3nwyrEfX10EDJ7CymbDVqms5yOt0BabS+GpH7aevzwpiWmCOh+TdmI0VtKZ
sbylDLlrQ/VysDUw+CN1I7PYncNgHEYboV9gM4lapgW2GubiluG+B/SBLEAsNdhy
wrJPWmztaGtro3SQYAUCFvnGvAnz3yAodhClVEn5IYz4S/ntL/wdNt3oZmkenaIB
PTGrKSzrkZ+m3JH9kiBic2FJUicI1MaiyXPpz7Wg4VWHzrtbJjaDHEZ/d8dyGjAN
uXdbyYnvAtaU4CsClWia2958AJ+Qmoi3zcKkkn56kIbpSLDhoMRgaHmlSAjaHOeZ
ZHV5rLRrtS73xls3CouxQUL/TRxHjYT5/F6n09EkBn9UMNL/viC7DU3UnbFrCunY
tvfCdH8qF+H7qrt9Ct2hOGWfJnmvVf2t+GaLttAvboB7n/luxtP1XLMY1n6PUimy
jj8OABSx+XC79nmdkTp6z14RBpOU7F8LQPqCoJvH5vg4h5emeb0C+9wupwq/4wuQ
2MnVNuLt2O94fsFi8VsAPOUnBpXwC8bz6FO+QVjOr6i5jP59400e05F1i6OOQD3b
OoTdm8/VcRxAqkEtQOv93Wc7a7DTzJrS3sit5rMcg+bJQhTRfCalxN26edWEpDvl
kNK+R2rWyC2YwcFjvKW6vXGADto+XEue18owkVxTwY3BpG351v+BL/jLyfQoGWGQ
kZdPEgcTIIwTG6t0lKQoASKq/Y/3d6l6PJaYUGoNmj6tIINwwa28jcK4bAKDewh5
oqCoqbIKL0AjExs/7NgMkkYqxuTUXOSjZSSHlIniBtBaCKnQeAJmPlbp8bapXVcA
r/nZKNUqDJ3D5wa/GzrEz01b2q9CGSNpaO1O3px8GxjYS6i8nYJDGfMBJjEOI5Ga
U+M71oa0vBa3tvLe31hJec7ed8hoGtnUS90b4FjUVNDNQs1Tv7cteNyrcH3K5Z4E
sk/hglFw8BfMwPJdNYMQ24qY77WlyC7OVnzlnadDQXy3UXY85jS3EAtvFvSwJgzw
PyBoq3snMS8PaCPIAVfp03DjFXEjGQA+/c8EGvOY3b/yCLtaE9N27QHg7IPyvEJG
+l4CYu9GCXfQ1deJIRRnW/tkCibJ6Ia/pmuo2rpbT/kVNU4jhO8Sd+sQ29NfWy42
UUJu1Pu7+qcPawN/RZJy3zohrK2GfKVWkqNcAp0Cpi/YIECgEEslXTdcWWkCoBAk
L2ZKuBUrETF14eRlNAv6q7y5IuewdJsDAFilUgpjuqmzJFlVjVHy6TngZTmdwVdZ
D/ueL3qumk0qQvZUCoOqUIv802D+m3aLdunU+X3ZWtT3j7SXbN8X7gMQi2oVgNaK
3zWfupSVtWF5LsnRVR451c7adNqrUGLa8vTzp09BbTZiUa0ExdXG6LgW4iIu4ELp
KJjJ1L+aPOluH5iyZw5S66CCgJhqLmtOR9S+DiUhwaa3UTMFDmBMZIbMDQginYD7
H6ZepQg5tBV36QKf96lVwtNwcTIRThiS0BUvE3qHWKFObvSd4+QH5HoWlg+wMi+9
5SZtrETnIOAQFa49UeKb99/I2WxVSqQgd0jJBGggpyz+7Hfn2Poucaj+cVvh30Z6
4FIWhX+4VrSoePGEq8TOPt9Gmj7xo7KBsA9VTFOv2d/esHu6vvi4/5i5pA7kWNID
gW3/jetotTtDLa+WPlsc2OtRYJ/5GmkxAZmz2fpviPnR5ulROiKzgp29RFGhdJmm
TB9ZU5aIHJHmBpD0Jx636Ip+hMcENMkLD9rFL0UbFBtAxjjo5oObEQ+V0kiEoNPa
VHD69Cbspf/ft6XHYAPhvVz3gBWyhC5YDb3bora4rwMGUMYLs6ES4JtaZOpS/J9k
D6E6uCz4lp1GGROfRWC8pxoQ0gDcYsxAmsu2jfDo2mo3aRMwjzDPgiddmV16cNBW
Pgn9VOG2/SUImJmpV+n4/l0vbq7p1h1QlNx5KxQwe7SiYM2aIEOlhtzN1v/GH7nt
0GU2t181jLoL2S5ThkfbQlJYDR+QbSXFNqsm5Hwza8HKODC0NQYyPJRtnpVf08+7
4sHvLj9h5u1OQpHpO9/VRmTvMuz8y7gD7wt51WYCSq9cP0GcLGMuq7w6wsscLOF9
sqyDfWls7bVTnA0leSWgR52h/Ssgggq+0pFWOqC12YsoqpQuPtp/qSrKLEcCd8IE
A5JxRQ+DEURqNBC+e+oCHNhizIRJ/yMxXJfrqMnVz6Cmj43sFMfow+4aydGWXQtr
EN0k6/NqxL1QGfLYECatey2vmYBrRhng6c4e8fJzSv8++DZw8/R4+bwZdC5H2fqD
KYJF84KyBDZ8FzLrhqXwu8Hwarhz0fYVSqQAVEL3862cs/yIe8QDvYxjuq7uOI2d
2MRvMGonLJJNKqlJQ7b16svLfIdRWChf4nfasCWhKI20p/t90Pt1hQ4Fb9NuIAQa
K4ccMo1hi4AJyD6+++6HC0JdLLoaUe+ghWj+P8x0W35mONFUZ/tqS4xZQ+XtH5T+
Gavb1TulIYxMt32eFOcC/3XzPqGEpctgVaAOBqtCh8U/A4RIok+wi48RiNJTnLvw
VJkUJFoOKXbxD/SA5pD/TNOb9b7zBz5LycYgwIzhiROg5SaITCdy0ilTBrIBd5/l
yRtHZaykPw3/L3W8jb4YK/jYbHtlL64XmqzbKtpzgBCPC7r/1zO8q1XjzWMexFVB
hEkzT4yg3Xjm5vD+VVqOEvY9HRH5I9t/yxNDg+r3Zm7nVtMo+NUQ/svNch1r7gia
oeBBtj/bX31vl3HUT4xlXJT69b8XMPIoVd39FJgEciVHkSW2XesZ7E8R0ZvMef0n
BArkJYVVfN9MVJegUpRGB2qvb1zEXQgRIV4giAQwDSZ6j680M9/Y7G8NO926L99E
vAwOYrvl0Ahq7HJbCDcN9jXf7NbQg96yu2IagJDt5MYHfZlz0xMQk424Sk5LNWDO
F6c5PGD8qe4ouFZZ82NdY6x/qxlcYrJ3YprlAYf/yztHwmXCX0LvlvdVrfVtUW0F
A7ew+P+4Vay8op/RezoroflA2uKnSHm5C8qvBDiWoTcXUVKtC1jtK2QC0Xz8K32C
piIRM9SNT6rhO+ToH7XFoTfDRsOdqwcwNlfZtnv0IK20R6Dskc8uJAD+sj87Qmb/
J+Z+OxisYqunqnFekq+xWJVw/gvK4Ha7pHXfU/Am37uh12IItUu2msdAsLqWyCx1
3Sg+1x9Q45sRbIEwPBR28L1MhUz0eFYhNit3dvAmT0acJ+Ey8wGXV3ePZTwqUey/
S9i25yd68LK0n9j7WAdGXNXRdWS2UYpdd+DDjGgCFpvSsWy2LoxyLr3kdTnIVeeI
glCWzSS5nGNIq+xphfWrJiFxkctCRoJmqbYbFJ+7WCq35HT/RM/sr4ALi2tE7XWh
HTJmubmGxpTlGLrBWi23Ia6d2mAYXAnEmCkoO0im+L0HxPf9zD0qem0oVXo86Ail
nOK6IGLVMBERwlupEN0aiJLbRe/IRUyyYnbqTvo6aqiNyg5XvrXJ8UwZO2u/cah3
fA1ByNodH/aI1s+KimkWT5TGog7ILylvXU8T2NKgtSdT7l4Ivq7LOva18EdU7wrT
+yJE1JtkzqnYuggqrtoZdjfTzTReHS6pvksYHt4naGCXcqZ9vM7s7S/SInYed5qA
wiK4xbycBR4E8Wi1F59+ljRu6ZxKIH/ysk5k02K3Z+finEdPQHaA28L4to17xrar
3YiHR3hkQeAw2M2Tu2A9LcBFrgSUVdYNM7NRLIRssGj/RJ+9SiH/U5j0bt29TJvD
JRrpPN8DAoWlCUlF36F0141AMaPS91PJ2MK0NdVTkCp9iaes8MSJzXnNS3iCAk23
N1q7UBUS2vbzqIlg4E9Ndf8qe7o8lD14EAm793B0eNzoIXUPXr/aYwaCD5rn4Zeh
hJNZEkH0LIUihraS+E5+wLiA4jLqgZ2qZgo3fGJ6CAJXteDcAv8yyYcvuI8sjVSa
30DJmGgXq1HjxqhBvkh5rpjIblQjOubcimY+mfQU3P+BW5glRl4/eJ4K3v3vsWoS
cXw3faF8Qk2z6L8Nmt5kwVyVFpFCr3O6Q9DV+Z33m8mnbWMt2lnKmF1JacMy5TB4
fkTaFLuq1M/O0mT5ch5RiEuqZdzZXo6PkyxHro7AnxPN2Tn6OAmw+DufLOiby5Ah
MlsW9NOej3qKFvxs72pejkFR5njFm7p/w1mGwz2nD9z8Kq42cWfjO9RQUx8HPpvz
5nt5TQG2j6qUj3THNaUXaYZ0fA7hVYvZBAj9tOpeE9WOWZyAymBCfMvnM/rbYhJW
JUeu5CH70/WLdOC9HA3ynIAxpjUKjqjnMdGdn+T1kyQPDjGmOxl7+nykfYrjJk6A
8cG9Z5aJ+hQz9SEvxvtEcG1gGAhvd25UbozLg+xr+EVwyWc2Vx++TMoLrGKV5NPG
4RJGnMgEg5qLkVmhzEspLR/VvjkWgfX/mFaEbnwqlh9JHpWPfSIoAVpxwX5EDXVd
S7Aipa9r/3MfJDYfKbGRubyb6j8Tph3ZieUOK3CDdMlFT+HbtsA8OK1rI60vyFeT
3O75dPx9bZU9t5IV38YkgF/yLI/ETIhWOO5vmN2myf1LpSkgKY1CY/x6pqCNXhTh
KXc4eRpBFs6B2jVHdYoAjkEaJ9JskJBGaucCtQM9aRLk4J27B/w5BrIfhiyrSLOu
HuFnxiIqAWV2PIr3NTnjLCoutZr2k0K6CWK5OrA9Yh0pOcpUQpY9xcAbJRr3G6Hn
mQsdZW2BYhBSoioi0XTVOqUSuK2rc5g1J+nrToo+YOK65PhRXtrWhva5D7nRdFzr
i1OQ0cHUduXYYljZyGdNJmZ1e+wnurCrSVzaaaE14dN3AK18qe4bI3ZvwZjczBP5
WqTph33Prg5aKq8PaWKME+3pDzJVZnkjeNbOcUzZYr6slFAaa4pZ+Jwg709SpuiI
1lNrHNqWARdVqdgbSNAaBANhSSc1WzZ8A7XGaLrgNO/71UDerPPUr+0ul4Q4bv9h
NFe+MDtZ1mtZrixixMmIYx/5mHP9haONit4BqBXw5BD7dhpB+KJfqJl8DFh8uKLL
MrpCscaiEToIzgOU7ljqWmjY4yuJ/N8AYs2kx9VHVeZ4tqzMjurJtf2nzzT+ZOX1
sqJk/o2CNBz3qyhC1WxMB9cOTTBst0k/bp2YnLP/1xgzyYImsGB3fobnIrM/WuCF
eDouvF3xZ1OTmy831QBdWMaa+jQzE/UOir9Q/e1Z+9uYEGrdWMpZQUamOrsJMETX
47Jlrc84a0+VaA7BWFzW8cX+3+TbYD2amGy0F3SCLSZyW2H8nQhZK8GVcY5/tiL6
/owK0W8nMeGy4DiZRTAjjn29ai3dW5ShbV1gNhOu7hyiovOlNSOOZKZs/cJRS/Ho
BA/5fauLw6CiYJSOLL+KnAwwl8Kt/yk4uFiJqLNodegEZu4VghUnQitRzYwbAjt6
PxcKV6QCWlGtq2VJcqCPPVUFflY0P9dcWKLyZJoGT2G0usxTi2MYXPhV0rnPYqax
ShZA8FH7hPnDSZxmjP9u/owFRSeRl3eo/DxP7zpLnE29xcVhc9hTidaaFyxfE57w
D+DS76bkZzJByA4EHOPnwCjiK/gjT9cJu1q8W8TaKXolsmOEFGLpOeBdt4hxxpyw
kVHl8bnx7GHajVKp+2onHM7ZC6vABlpyAuvMrOZolXwJUuF5k7F9Agjs6nCbanwq
x4GR3ud+uho+d/oEg5Bfn8IGQgFnZWy6hZT3Wbu/jJ4IsN0lmci9CWlV6oWncmT8
L3ejxifiPKb+tixErRbyaNPgPF3a554W8acNCiHs37bsLSJyGXFrypu53UYDraYY
NZWjtV4zlkXoI/ddXAoIdPMBQkCDuiiwPEyJpxFSaTtdJEpNsKs7dIpEiaKcwrdQ
K4wdICxxbmVlNS7wpLSFV901sYrRZoaFJw49Ykf16ccXqIgo1DwuAHXAAKgXu6q1
dYG4Xs2lP5fSXrrKLSWh6QgnV6cnl9TOJfAVsq1YXui3nToOrJXnd9T+0wxK1IQh
Yz6OLnUy+wnm4OIyq8sm04P/mLBGZwoqvVaygKvSLotYG/Ve+bYpWZi2xcKryM5+
YqQjHPNSu8vda0FD92L6M0emuJ7NcyumXGWtnf5d7A715Z1pWHpDKgohTYLvPt+b
3cDDYjthafxQVUIoM3KC6mvY/Zz9dizUrLnNNsnHjAqaJ9E7N38w3Q5Ezw1NgZWz
zrtGaLfExSh/YmkHn7sOXIfO2Zu6R8lTtIlYF7i3yQy1rTgcwLzWuNSjo6w9vNIj
FJV0uoKHRmgxuWEKlmKcO8yDU+COHgNsmw+JRjrzOGKWRISSnapoyzh0XfiAIVTZ
vRG7yqJQKE+CCurueTnPqSpGbbdRh/3KYZi/1U2wbuxm/3RHMv1hk91LPvi0lPFr
AkVNHfRQG+wsj/PMbcL88GU/9P3fRrEeWn6pl1/vLhQmSSU8HdQg7lELQEsSVx5i
dexmhdsnPbAqWj8WFOhgN+OlBLlbiAP7kTiu1IJm6Ayau5h6KHZ8ol4qnDBmRQWk
8klWpfyUe52zTuhjzluUL8xuFJrClhK1CTcVUcVNnfbAtjYivnczWjNC8l7/m1rj
+ZmCdGkvdZ94Q6Ky66ZXhWS+B41zznHCCKCp3egddmX2DnHG5fUMlrTxf0Z1d7FZ
0995dl+ySyw+i4pd0tQbmPGVBfCbGnowqCKZ68kzmyH5c68mkCvYGhYyLBxBbYCy
wXO4HwQS36nADQXEbivNvxo/15Np8XFYQJ/R0xbn72F4SkL9JXEWxFY7Bah2zY4Z
ti+PquNmCL2ioeVm1EHmBP/dKMf/2J/1M7qNLtXY0TSzo7h5KAN6epE1QxBLUGIa
9ckRVD/y1YvH/RJspc/QJGmHD9+Rxy93eMyueZBRZSff+0oajTtgyDwje7/Wa1ax
wa39ygXp1hrbES8sWYlv1vu9Aet3wV3VttsUpxoNKAuAE4PfQPxhPVhia3U6iU6k
xQlHEHa+s+v77V/WQ/j5J7WgHnNjPGSWQbuVTyVtLUBvix7HBtqeSIPxD7gBjjkM
AZvAPAYqNKY7E0I6hu/IE640pv1i4YYpZObOlGxfPSrBGt7m9VS5J4oQPDBfjp2/
2RKgsri6oDO5k9wFW8hJIzzM0vLtSrtmDvM1Qkc1TcgIyxumFiPUwRRWULDldu3C
qkqG4utrMKS8Ztl6LRs5Ai6AQlJFzxVwbgIGjSRCU3uKhsFAPfBQxjY90n/Vo7Bf
DvhmEWM3nZo7+Cpx0AdgbKLodrZ3vrFn7C1I3tcBfBrG9ikDQIVxxWa7adbPnnd/
sc3n0gKPiIot1863/AcYcq1XJDIw/Z2hJGoUp7JpqyWb6J9vPmwik8T/7fvXzBfU
nl0v97NeWeq7JWveorEJwJnnMk5bHQNUwbUGrvIPo//+ChcwY+R+GONEypZWJmRt
+zn/FswzZOBqBaijmfMynOkfeoHsvRmq6YwtJJC8Jtdkynmgj1lmmrDqG1gBql79
HV9X8kIEAr3O2LPFCZLQ5dUt3WooCvc90K210m+B1lp9mQIRh3ZqZDCF9bUyc5DF
xZ9HBBv/rAI6yReVlAkGB3WLwkMukAgkYG/S01RDRuRkTvUISu3GpdxXS2uMhdw8
m4ZpFRepieELGJQvB1RvdHxrL5ay7vB3Db2fhfWE4FXAXFjLs73/2HyiHFl3xBiz
jOv8XW+01V7ZBcietqHuKtoL+wOCe41swP6YGHbLd7FWfbJSQtecX6Cjp3gSJHGH
RYPCMh+vlwt1b3stiM8t/cwV1nFSvh0OtDk3s2/keafl4BD7CQFQ33BkCyz/Gh2u
tjzdFhGvSXPiqpZMPec4QMtOC5lXZT1xbyE2FMcLzTejpF1bvod0W3k9+S5ikY/4
hKtCbURWejL+Ty/1aBRx4f4zl+Xx6NrunPMO3EzFJTiMMAa7wf2LtaPNRGZsXfWk
hzKknypq88TZJ6NfnvnbEHNi/cQ1ka3DJfTH5QTMEV81guRzuYR/qdKHnLJxsvRG
TzQHNg732TZ88t5rZPw06nkNfzem261Z1SPK82JeblcEo+Oilk7R7CF3WLPou0JF
oNNrG1vVovyFTMsYEn5JXuEEQ+CteBI7FnhbuY7GhRP5ID7XZC1K3IkoA1a5DNwf
p7zKysbVc3PzhnqWaXqdd9hXFQ7cqWRQrejCwmoxJlxyoQedDhb1BwA3KkAdRhPU
fOCysZiVujsVShrOMhoBRlVhE5zibCVitx6Lj7r7kaX6PK0rw8SPdGOIsUfqBv52
LRyxvetNVjoNP+PlqbTjJOhBvr4981bhxukFre/n6xizX5XaYzPikS0YLsKg0I5F
jGMZZ/MaOm6cS4niZ+OfDhktK6j23Vpbu94RtjbQc4g0xWUtg7KJ/w7/J+OIUiOH
QQ/3VbB0GsCow5Ik2qGy3hm3Zev2ktWbVvI6cABF/B0FQOYu+97nWRn3dqnnUFUC
G9sVkXHSnfvUTBzYFtI+fLZh3dVvxWQbyH6uvEEZniNO9xsxi3enKWG2rScy0rw7
DKXP7S8bZ2DnCIDrEKlyZoCfdMoDGEQOe1UjDk5/hIbQRJQwgJY6VDdOMtl5Zp95
dnwB2h0xQ/3bRfr491SBppGocAt8HnL4Pi78GPUwKNJ5gZodWaEfPhDHvmp6Z5nB
Yq+1izTeqtPZhci6yfBy6s1rcIISDU8Wl8fsKZ1bAsp3bu/w1FJkb7KymBDzQhzd
EHTk8xqW/6qHjJGujWoK7/PxOn7/N2wZ0P0BjysDrRDAfxio4kBHoKRdELfnLN3c
pHklnacwSdZzjQL9++jmY7vAxlggw+6/ExxznQBjHEYcaHDu+622d92daDzLdrZz
JQIKmYyoVpL0WrJtzyBsAdonF3wW4Z+KPoUyqSk+EdKl1ctF5KGMMS4Grwyu+Juc
2c9yQe1rkEvkkuZfzj0g2xO/2n29MJgtj6r7mn70KEM6CISzmzrIBHnPZ+UPfHst
PBQaB0u9uLYWstOma/Wws8/NaJVk/Jw4F4RDPkC3ZLzaf7yl08eptfvupZ4ZOxLC
W2PuInKK9UW/1v8wsD/ED4YFoDwJb27fD6slDa7eity2cDkqD+Z7ghXIWbH5K0Tx
6vgSWxcbsBvlnUdZMd+ed8UjXycxPLG6d1hM6C4q/OaFBgKRE0/Zwl9HqJQjJiGm
uIQOfFrCNUDVsyUW4IKkEwuNgbxE9ePe2PuAo3iqnhDJzIPeHsvaC2hEAyJ+v63O
CO3+1dY8uXFqqtBEr0dJ/ycPxrHj8d+RyaLp2XxQcjKDVSMkbkyCCh6TE/b8e4k4
mPntw/nZHmXQ2U310S1PwJScebnvXNjIRYEPlickUaHqal2tfGM6DZ5IKg/VLjuP
SPzj7ub2hJRY7wxJ2tbmOUkxDagZQMxAoh5MpbZOxJZw9ujka7FIkNs99v/tj/aC
RqHCctxThJ34kttI/ozrHKujObp+Y7VjGQz1PEmZKdbeUOHNrwKOb6zRrNIf0LWG
p6pMUYLwbZrszs/8eWbrIp6p9twjsLL2DDwz+sHKtYcGJ3I4vfREcc8MdUPaHd1j
ntODB/PxUiEbwLWSyRSVC6C54uuIN+ETYIigfj1Wt5PI+Bz2jDP1NJUj3CAZ1tBZ
PuSinxCIUXApXjL9h/ibbINf1Xdu2PernQIIalP5WXiptTuPKHqKo8Tfbo+T2TYK
kgX4SN6/+SY1mZx1G4cm6Dl0qenTktyPZfktzjlRG8RlDzgivEpoqK9szMPUJXtw
F9GlZDyLEOm8Jz168/8YFYfD2FNX9qSaiRACKXfHqLSrYIk5nLRaUyi1fj7LThwC
K/XfPjDe903GdML23BXfN12IxEJ8DryzuYLSftnDPMD5qBwikk6aEOgybvzOcIcR
mCq1E3JoHs1MLxfcOSdFiSl4x2e+plHaiN6w+dIkmvv/KasoMTx0taLAIKXVTQdq
AbpINcbNFyBTtFa3Fj2PRD5nwZc/QPwu0NxygthRwRCR3AyxkJWmBAm022tCYY4L
MRwk+XTg/OBCNTAlroCEvlBL0PmhDPCfy+1imh+nIXaJgWh4jefwA+3AAJkXadn/
30xgb7B5iNQbHNXIHMvLBuhWDjvWAHtnJz37iSagSDJm5y7kye5hTSaNY62PdprP
fEe0bkiJeLd5fvdSCcoHc6fgpT+ZMce4lsyjAR/J/E8Uj2zRARGJxlXthBizdP0X
MqV9R1In+Z5xmQwoZiYCiApc76xxpnLi+WDXdHOzeygILl8xaHpFbFZ79QWrEmyZ
AKLKIGkrXODJz270tcQi1ZVoYZbfM5SE9g+uKu/POi+mTO9Y4n2wus0RuDcVuil0
TiXW6twdXwiTn0cY/CVIBpmO13W4pDjS4ZBLIq7q/ma8Aj8ZHCr1YWqRFmINdgfD
O3gqswBqf1MWh7dnm2Eja8u0/kMDq4TJy/eI0OdPB7RgtPEL4KSp2fzzSl5cTDi4
sDTJTznBx0SJOBVstJpHZlvm8Py3MPFo6VGg70Ofy45YlyzmfMEHeQCH/rsWohLg
6ug7kVbwX9QVvcZ7XvN2vXVfM83OITlQsnZjSiKmN/JV+B2vWKEkNZUpe2LblryH
H+RIoVaQ90mFRGr7FvgwyTD+6o8UwyseMv8QrItdO/MQ8ZozHdOdGGaFbgsvKv5p
f+DgGF+Kzs/0Lletr4TD1aiRt+QG0ggqF9CQ79iWI/GgjWiYOMMYI05r95ZoD4iS
yKP3suMVsG4qPAStS7FbsDhQwi/rYCM8LS6ax89T5kv++W96fi0lfI4cBR8JT++x
edWsRrWf6lo5IZeckOQjPEghZ+zA57e3NoZhnPbJTW0Ms3jCAX6d5LHV+7S0d3RL
CjL3tk2QZnK++iiaPt1Hbba31wRbwcfpSyjYxk3UIqkgTNu2NVfxQUoFXlJOwTMj
EoXcDudQ0RTP2Xr3H1LhxwzE/Qe+6R1OhyLfKXVX2OAoHJ7qOQLXtdGpFhmHIyRO
/kUMHeTa4BzXwrPvRWTjGNE5XieL/AWOTysr2qC74UPVTqWdoum20T7ejBheh4oM
nIyo6vHx0qx3pDDsrEsFAV1o7yfQmZ7ocxxG6wudkszMt1WN4BFJa1nWpkeIuFpq
vNc5kBv/+RKA/234Krgz+8OCfLP6O+VKqaOuapLo0ls+yZCeIHmWjSf0P6qgeXss
OyR69jQsfLivYyWSxEBzysDlGdyFkGLIkg78VYokYEfYBK6uPCzDA81Hu0DyqrSV
UpQ7a7V8AxZdWu/SYFTPeeINgBrAWcgeIfGROHQs1VBjKPVBJVs20Qwvz55gbMGI
zmlMAcMEjfjOEt7aU/CnVee46Kiq/HBjhVKoVAB+CDL/9QfdLAuMyNzVwibeb1Xs
ZdKTh8AfUwnkqdYazOExV2EWL/zELdn3Ji/tTeWDfa2hMFfp78yd7j1aVH0B8f2P
qCLUqMUbBUZ0nGGqG8pgk2GAx9AKJrDGa+gzoam6qdxLMxi5O01t+k6RP7Q6iV3D
RVKejJJVhz2ulasdgyS1+/dEHIPqz6U/wzhaFNYF07LevvH17EFyn1RbAG9XMbip
JQaxbCQa2zwnkP58O/8DlbFuLczpz6ay3wnjcRV5o5qDiHirS7EiM35qTvX0qWBy
s/r6STima1+LNozwR3WG+Ezshu/go9v502EvsNJx0WaGl1bdZbxxqhzoNNQtqOv1
coWoRC2CXCt2WItGU2o4LVs8xkPF518XrU0QINoYUcFZA0C4t94tcm3E/7rMR3U9
/pmYr3nlyivqdiCeFjqS2Jg2Qo+ZhrYW1COtl0y9wq2S+VWgcU1D9+AruLqnLib1
2fGgl4mTICwNN7rP9Ra+DnWu90Coh84fu5hETGCYKCvHpO7dLJLM9Icq7dBhSap4
SRaipalSfCHCgQmv4S+JLSpZR6YA3Jr5MU4b7qP4aZ/5uz3YnfW2Yf0Ma8frv5B/
94hczkjQTpPcdHSys99ebJESPyTdH7br/+mIN506G4SgMIVG+bIYaB+HSWLtPjg3
AnkMr7U03wOQE5zumOgMgRzaKLZma/yuKdLK5c+V9KcW1IRqRc37/A9iIlxyF9Xv
nYbQ9cyFf6IKyGKimGvInKF0nNzObNTkPDNG2nrtCyY1oXcTWr8t9msWTAD8thip
X9QaZLPpjXFsRuSqYXz54mb9qxTmedDvzXiM2w60VuEcPGTHiXpMA9ry11Skb4+E
QNde9stF2qYAt+RyorRo8LtmnoAeQA77gJBzUCHk6FYBNblcazWudUYBXJIp2/0M
GAROirO4ky6000w9dGWA846Dc0E3Zgl8bezWXxeGgh8mi98D+McgWhHIxZnj7wsA
lw2hWqRMVAQ3btrQ1sdX9jbBOBJitBDi1N/eMNB/Td26OSbNj8B6EgE/JXtHL+OM
KWqZ1jC30fGN08tXaUoWRQhnUgRv5uu6003xvnD3QWZcrHfA99LWW9dmw4XrDxpI
FdMsAawBSjPGQZgTriBRVLasBVyP3nCMq3FntTYtoia7ugW3Ge8UFEe64KlRMNCd
hSBEJDv7NJMJtTIjkNQ5aEwxpwKQO6Gze/w5mbELq7dYjtSXy7pzxBPILbwpcJWd
grAep7W/GbgtFFhO2yTzzdq+9GCFNMZ1qoVmAPATnbbl/aSB7dLfJ+79kWKuuzWU
aRBcYXrdba6IGj0GBdaSIaQU4TiBW8HV98kiz0Tsi1qmIn4Xn/ffDtGh1yxC37Uc
2kHp2dMhVGUuKxBu8UbA5OOBXifPpYJau5KZoMQVXPrUoyHQkwu54MX9cXqHiTAK
aITsttESEvRi4QtjP225+Z9MOq1h42Pcth4dZf5G3jsMK2deFJPvr9c/OgcG5W9V
WAi57Qxx7lEJiLsSHWJKj1OnyZm6XJpG/ajVjKb6GvVo0rU581CA0CM+i4B+qwKr
ApX1LtdtzCGJwemVuHuvmzA3L+ru5NWspgh37NcIphRia4JuTp1TlzGnuIxC39Ps
9kqTXDx6Vzep182LyDgV6wJei1B2dO9KQT3PquWkIP7L49wzp+oYC74D1UYVqvQF
IuQm1oxg4hLbYSuJXkjsfjtwnXYity/PvLhLhwJ4zVudV61X1L6u8kc5yYht2X//
x+NTSHJM83L/XOVlN/K0SwLi5eJoj/q+9NVpEuwUF9wQSOsH2GZEUFA4XfELxd03
ANtp9jVc/Or3u05C5jh82JM1YvmwmXsFsKhyRhaXHOubdL9M9Dl8Z5itXiEaW0U7
xvgokM8n7L5fBG7VJPrYt180y4q5S47yHKS14PqzSzmOZYA7JiUzfF1DDI4lkJod
KEgDboolcoV6sA0Ekm7IXEgrp0RGBkQ2M907fLtOL/+Cwzd0GlA0fXtiDXKKSV2A
/Bily2MXzN7pxEPgzpOFsAhmRuDjwGmAQPvSnZJxS0JUblF5T0GYsQw1CwuHqAZ9
Z0d6WDQRmItbW4qocD6+GmfmlYSQ6ZvW9UtZyajomXRkw8orbZBemFtgHHhElQ05
R9x/kh1KEuLdN1SUrLohHWfCQn3z/mA3J2+XaCqz6D+Yo1xfxzGDL5mo3uaaVAVJ
XBfAGMaFGHtVPyIzzjWohRtmzpOrobvfO4KBRFXRC9Rf30QcTgnSpGh4ti+qcwD+
59LLvsw/YtZ9O82u5s26ZCOKwkU8pyM/yjrB0g1aHoCk2LGzTJ0MomHRjQulce6Z
JCPG/XBUWH47aAoFWHuFUNAor8T5N6ISjoPm9NsgeCXU3bjXENlBZ03wWPJ3rHtu
BnmaFckG2aRRA6OlxTKrRwDCgDCAbtKsF1b0l7GL9Ckh6y9S2/m4svqHMFqbvSrd
B8HkqCSD+uo+UvesQGAJlDP3PD4M1aGejW/0cDusV9SGcb2AWifORvrkwAFjpOQB
K8NmROPbYy8Whmo5F6X1W/rwkOi/BVMuMY6tcd6UOlPVX/aFykf8qdG01bN3loru
lharcdIvHV4kLr1PfGT/Oh6CukU1b0k700NsnoRnMerd4+sI2fNES/qU6p8T28ar
u5vh/aA55dFvtzb7KzFUKVcz2m3uvam9TQtZaWTMjOhKXu4KWGBd+3zY3gxmZyz5
OQyZFV3G6YLFW0YJSZycFgwCfZo0M9VCX+cHNPMFso4rrUqlqrNPPXDx7drOM6VI
h2iM3ySanXbkT38qz18SW2xLIfAdZo/tKyLXYoajb+NIRp042oBYZUIneE49KfEP
ANLFiSMHi+jkMQ/KbiA5I+vrAzaUAYWm0mk84fodd6tOJE5pN8sjL6BTCthBV1wz
9JHBVTTyC6RTgPpMlRQB4+4AShFoK3p5ZbHHwFJ+6vCZp71BU+vJX5TpMH3EIMWP
EmA//OS9tpVxBlxhZ/unUcHdAu1gmKATcMJ1mAMx7vBVsXukjoBygHlVOdFKZUDj
NbllRcaAxpapio06zUH87cCaN7Lji8w7crDvFPp7c1UynrzLWrX0PqeAwsrIqVP4
PsgABTO94nI5T2ACXQZ6XMJZ9yBYtxfEeshzDkxIn8WTNWQofT6JQUTBHyYn9JX9
xdRH19/Ulj4wUx4tEsmloD2kzyWAewQZQPOmNj39e8NFeKX0583xvqikVHCCFSzU
wYDAv7rZryKFwfUVTiF1kAurjl2MinoIFxzQp7PE4qYKN8nzl7apPvczSCLz8hIk
1+K6gun4HbP+iEdrpliyF6rfsZT58oxHbPrNQaEcbQ6gGam42b+zm4HplT+PFf/2
WWY7k6ZKCu7f5Pqe51bGDABZ3oMETMCqAVfMhAzq7gFuOVPOac4ENMRTFIWbaQbN
+5y2RcOdLBk+Lk5aXUr61Mq+gjG0wpf56FfCjr0tUN3TZWjGHaVE3KzSJ5iR+UVH
aTAduGfjdM0WMdSiYUS22fjHpdMgDT0ZJhDS1WnkZOSYbZHP+yjUPdqKk86mKuFl
7xLMJ0f4oCdmwqNKOK8bHsQbRLoGa3B9AenZH9txF4CXVvDkB+RUWE6BB6xUA29h
vNKxLfZF9qzvoRy9ap0awTibJNBQzf6ivT7aP5VJA3CmRVEsp5VEoGevC3j+yQWX
tjhfXKgdYVmQuo+5Lo8kv1fLMecTanlR4ZXNtoALs8m42JaIJIWPXEON/UxKiZtV
Ene999+Ntd3VWVyA/2drt1HOZHn3NB9nAOL56Ywk9DezSrdY75L1vH/IPKmZqkWJ
wVKdKOmpCsgeOmpGVbhTZTU03bJE2zZEPwp++4xDumiIRh852zrqN2TO5ikwEqoC
G6E/S1/OoYnczam6JqAe1v0NCg7fOvFlTMOTd3pNUZ1FxuBBLUrhmrAUIrJM0p/e
wZcNPnSx9JiAK/D+iQW6O2JSzf8BwMdZPpBYihRwKQdtWwhEp6FVc5C9wcxQevjS
TuyeRUBEtIVmBtdoUaeh/W62Z+sDj/x4a9kosrYdCB4Y38wG939ensUXee4vzz88
oUlYz3BoJifTCKklLKOLF4C6mxTWinnT8VRgBvTfORRC94IPRsPYCJgQA1OEyQiC
3D64twCLws8hlPkxpxDMjpXYRk7ec1NIw0OsHmdNh1cDjr2lOtIPFa6+uLXgLpSr
Lsr1DvhiqeD41sgLFlSrJU9zdH4KyKGntUb0+Yuo17yZau5NdU/NcrkVBBUh8Bzu
BsrAHyUKi/0t/aj+Q8YLK1nKCtzHWJY8wo4I2+bVZZALf0FXQ3D+BLev4C5H5kJ2
TbsOfDKANCu+h03rKSRmjskkDpxBua2N8fFfVN9lFvehJlwdpij4H4X1URy5TvO+
Bfap5h4dDpUrxMVootbXVkoCJJFjlN6pMRDLlWSuWAm9TOuX+E6DwKk1dqCeCKHW
xghBZVnb1r1cAsQcrUjAzJVenUWXhuyHLzLgHWhFqyuoWSk2R59UXUOi5E3zYhMd
ew/nH28sPkp6eE3WlfHgw0XnykJvC5m34aTgXZEVcBDZ9IClPCYa4FXW6x/Top2T
ShKcP1i4G18N8IdUAGAza+21EL8+TmGSAA6nrOAROcawm/eT9742qOsYbYADTyOT
TcddhqVpd6J+bC5ptKtta0pWLGcWGbJhNIWWQmlyHIOhf8tKdq3G0ormbVGi67Wh
144COTE1ld6cO4AjAkA5VvSfJ53HFN91JQeq/5neoY/x6ljMNH22h1psZpJ4b25H
M9MgEwtnSzP01rDcLtSP4/BSTKeioTCFQM+qOmJ1XByV3m6nK5mswDEp+hv4VDZj
S0ZvERvkxA3xKBxMdNOOpu1kPY0PdHTsvzXl5EidxZv3+Gge6Hfs/B46dYIprnkO
9u7pPslKd/CnO9vwZtKoUzNKQCKATCKSQC75+t6iWKwgdgwCjPkfGpLKwDJttJGy
+qFQHLr6kFsPIZevoUAOGuyztKarUYE7VcbtHVROatDnzLbHXJFv2WhWdEEeB1Xe
v2uO2kT1ayD4Ihy/gJBYCS5DPC0X2JNTohjNF5pwL1UloMjhv0+iqLnsJIHrZOhk
HecFqVxpvMdveWp/yP6VQAhdgfJaYzRxkqOx0ReL1nlUi437Vu9sgT9XKfsp0IB2
mCn0BxD731s0F2WkS0eGTEGFUrjWGAKa45bCH2WdIb6vRafXKua3wygBcX0rVyIr
w1dWCTmfbTqhEgJQN7xbpK4kGZEQ2UKctW1ALeHY6Rhql28cQrW9JsibVE6Pz4Lq
bodKFCO9Q/5OG2jnL0e5rO2uvw11Ck8Su1uD/dou0iYmK7a+enBGr7PaqdfMr1cb
MMXIP+TxtRuwGQYLtSLfAQxc6qgbFX363owgHH+X8VaOYDXm/URsNUj95U3QOgf0
5SErq8Bw3DTi7pBCtecQiMFMdRkAjyg0E6n9de3Gg2K0muxf+Z0DV2wqQ0+GGZnp
Gw8HoeiMen3QI7ESv6cyn1Lc63MGpz4LKORBLY+Nf8TluIhWBFEtgrvtJmRvc0qK
MqJ8bL5bA/uDQjjJyMwvMM2WyTcmVnQdR33LirtALKHOVv3VURSDeKaGm2nlG91y
OSsD6lqQIbOKm8QD6rsskmSvi85kINHCnWOg5JuRUE68GZD+P+OtA3JwxDZTiu4K
mCvyv+8PCNXB/bzPQTt0Ds98pNpB3oOUBPV88O6i/3g9NW8Sdc41hq2EDtjmdmUe
nTFlRKFBPbvvmsmmcq6uSnd7HyRslQHOFRFShAU2vgxaEwFgvoEPenIehVNyOHjD
FBDuRgXWZr39D4FeOMNsIfLsxbHmNPObAyFHDUbWGI8/89u6IDagWJdBhm6xNPWe
Jhpt86lHczbTtNlSoHP5q2sONeInohy5QjJOK5VVlSFaMC5VImwUuGr3dHtRoTZK
pe1Tb7WbXXK+p7mgYw2EViy6vX4qcbSvgvEy6nKrsKbSGsJm8le3LAzimxXumaeg
AQQLWYtBKq3TTiAolX4ZNsPewNseyv/pTQJs1jH/7SscwaYfuwd9oeQiDzECPdzQ
TpQdZqDWo0tY5Am4Na4QZ3tpJC6cuF4mHOPN2SKUvQlrvHAb0IdBuIe8xnEXunfg
EIKMFQEjmnphmC+U+e7YfCWz4b6XqfcMcJv3GAZd7f4MXpaZeBg+TfAg1Zg8cs97
pQJak73nOZISG2JIydRYUDGMhjEiXgt5lfKGpAcZWbqFimX572/UDpp9YEghZb6Z
tauKTFWIEngIh4DT6SHdvp+CeCa/CQ7Grs8JfapB905QC41oSiR5TqjuD9hK+AJy
1Xg/lFntmBd+RNy0UWBcd7HoRTyLacjw49lidx01OP9qPwQXVtay4SKkCiBeq84u
BqdSfcUxcaCYGXis8SZ3mlkT4KwffymDEPaABoOSIkgS5lHzjTcGfuEPulpzXkfI
aXGPThFE8WjvILBfqHVhXnFDbXf0Nar1a7YvM32xLDrXaCIBnXNHYaB/YcvTG2m1
GmdnJg2jhrGxOMGpIA1eU/82TK89znZgEuTlwSCpOkYQu7XB2APkze1bTaWU1TFG
O57yBHzRBxaKku78g50KFsqPgaqqwQGAK8fr2BQN8huUIuOJmgf1QVC9+iHL+Lr2
jbtRPYFPPrBbl82q0p1ULNm3xmrwiMMkUpzRXD2sZKD4yBfyHtERqlLLVeAwVQ6T
6vojJNBYv+ZQOChupDICrjXV7W8gYlvHWUgAAJ2EQTtJOwhc8WCyy15E+v/2rn9E
pIxecWqTJeTpjx0dXX6QFUdsBDDDrMsAPmoak60Mp7tOTRstIKG252P1KyeLL/Ct
h1yf+p6t7FFHoFW4qr0Kb6tQ5rSRfsMLzK66jpvpaceZT5XhDln6Qlu3/hGyLBlW
+aGve8oNIWMpomai99rN1uoGGREqQ3RKCOtQ2KHGn/oXz/lf5osN8l0MpywE5ZQd
CONlskz0ZNBUEtcY8vwpaqUSpxNZe/gL3PYVPj/ZWF+9sp3NeKKZlPEMzyykKkr0
94F7HDiADfyYmeW5jTQdNV1JqRQWNPUf7P9NfKrWkxQ3F7Txd9bppLvFOZ+fhF/Z
KOOgxrxvaUQdGwhChCo7mK58ZDTg9tI1VJoWwcseXOthfK13/jCOtP1DSGWx5v8K
OGlpKQDbOkO07pOiHyVune3QziQvuZ7I5471OqevcCx9gRo8B7oIqt+Fsp8Vn6Hh
jOkbrqTqq4TtNkjQna7DiC3cLVglzG1maXWUURgogx8frleE7daYFWGLbLoLlldC
bjN/E9sYwpneLzr/Wb6ZnRaggf6n4CTpeSNGKZHTVPcGSohRLG+B0vcyPFlrt5if
EssNS53+aGZpE7op4I1i2zIdI9MSLMQta9rXU79Y+G314OOqwUwKoe/gVAbWlAqK
5Iw5bTGpWqMneZd6BEnoE0zoHEhwg4uKO4lt7bxBzhaatvFGvQhZd8h0CM13fkt3
fVcxddzQ0zqMBxOncpzUJe7OiEBP4RtocVOnjg6uHSu37yzC4R9tpBvNp91FA3kO
+uCAbj1wTxNqx0oH7TUBM0gbJkyZUi0SJyyAmKDskijSrF+fFBOBLeCfuNU0UZ0K
Bl0q4TQmtSdg454b66rTWC9m5RgT2ChsQY939YNsktDogFlARR/Qe0NPz+nlfkJJ
BDPB6urZHxIH17yLOhT/4oUHqJmVrixgJNSSwq8PYthkZWr73ybim9NyBXRUgpYR
RH4ETpQRad+7ELTPtHnD9i358MFoDOw3jsnzbriu/T7Xl0PA7Fl2YYWuYGlvA5nC
VGPGslwjUV8fm4ZfdDhVtshmVWdv6neIeeJXVIJ6dihtvpTBWQ0tC+yQUTdd4e5z
tYlsMey6rRx0sIHRIPqYe08sh9AFVqno6vh685i9129gv2csVrnODuu8KV8j+goy
3EqJPOT1p7ds2HM3cgB5+OU+DFFrvSfaCk+NopbQJxLkjb3IG05B39z9gUZwUBWA
7ooiPWpXDJqE06QAYXWmhtQGHxagNY2O2lNUSrB1cuIHDsGI/Uy57TQU7mdm0Vnh
3uCbOyI2yto8DIWq3TLFXnDeLjExTXx0FqBCFlWdz2oe0v8XGv1UN3gGc8X9+LxR
CdQkU8gcA7B1gDoI7/Ee8Cref3XI3/Qx0u8zb57K2I4fG2cWP8CqCwzsr5DGEf8j
4wnezn/FJIRs4EmQIvf3tlMoDMBvjwj34A2jp0NHzMV2yJJGVjkv7905FWWpmSmT
1eLS6ZQdXPmoaaSFqIdlogs1uO/xfJW9L89W29Qur7lPAa56PklvVpntHggbXZEV
EWJpWVxXhXkwwTi84hjWJrCHyD3wO1efQ3XJxpOtIHaAKa6jYjNj9Uqc17gwsvBD
MkTKlVUI74J6vvdqsiP7xpDhEiIbcDHbMHwFkVBtiMmTfu2yHn+Wmtw5Wf9cFMTZ
+rc5BZIe3F1vICFEaF2FetoMMcBXYJQRNgxbXywVPOLVro4fsj/961IsRPJpqUGW
LazMkgpHi1aib9IoMgqOCR8Nu6gK2jSVvn8rIcHUJCMpMh9M5KhAoOI7gvU1cv4I
fM8AbdYyyf9w7yFoOw0zrkGajjINLn/GiPH6hmmy/o82e2p5EDMM2c5SQ6bTGwh/
pm0b/1/HFW9CCYqm5E6GZh8SsN2YQNsp92swK4LPtdeUnzU4QmiOif8nOb7Qdiid
uuzgNkrMsbR0hC0/xZuiTQxi6C2ET3fuCWvRAi8E4maTVCc6H1tl0yHyCtg48Ozr
88a2gEESh0M5QLuIbowTQ4ExWh2joS8NJVzzdS37+VhpB/7lUMMguTm2JwYY+v93
XHGN48r9miIx764QYnR0uWStn4PtZFUpVyRndMCWbC/uLIYJmx49OcWC1meB8cp4
x+Uce9bt2dSPNRPOj2hB0Osm7PxlGjLiowwO08BOfPES3z60ObZykBVzdix0y04l
VacOWqGUP6oYCE3bRmZpmL0YgvEkKHIZhd8g4Kjc5lIhptzEIbNQRAmQR/zuklSk
NMIVL68iomKXsbcCh5482V7TQiYf2N+M5jk7OvDNlyuDHXh0qxy1JfS0kG+3q2L2
vtXXZkI6qGADbHI4Crvkc3i4oo7l+lphuU09z3t0hCP8DI+pH3hJ/OgUSp4g38dp
OXKUTs0B+sElO6/IWQ2DqmElUwbJtE57D1LK0oSIA2iIwEdl1HsZRixurrb6VoOq
RoygeuiUCM9dbuvLuXHl5KR1mKfjdOV1X4jIVd79/I5RJzj++BKdCqz90LnvVVd9
I9E6aKzfgfmVizubU+vMKGPrwu9Lt8I9aEsVzr0QKQr+Ztg3EugC4pskEL8g3sUt
1UcY5l2EwR1mGIOcAkNr8ikBf1G00dt0Kz820YEwILCpcYeIO0wtXRks1mlv7wIx
ii0dqfFC92GYcp7gPwmU/eGplyyCAKqLpFuk02LQkFtmC7e8BuTf/Ka0nX/dDFpq
LY8SIDV/L0Wn+J392k6qm39Xsq4IqXc7hlwyO0GFz+8Ul16lfKrkrUTA8d9Upy/S
c1d8/dzmMFGrR1IBRI8A/Ijn4Q2PSK0Uup9d5rVZsHp/Oaw+uvbCZrt/Okls4b+a
YApJfS2ColVMJyDwCb+Ka3CKORrfNThZ3+ktcDn/0vssO0Tzq4vP96JumiajFoIE
/k51igfCI2nEttlOWuimkIUfV1WKyKtKmoDGAyU9IfhMbN4N+wITWMBwhSTXXkiJ
f9XBGjO13BarjRxzTsCHwez66/FyLvReEMnpxNIx5BDo5kdM1MjpQgkFRyycjn0N
/4macUeLBl9/rTM/np3obxTm/Dp5FZkx+kWWRGS1QYIOpfz5R3ElzsI6Kmt9ohGj
AOwez9BMXxaEX1upROV3L+ekABrt61nB8NXpvdr1UKHJJD8cToKtaFZ0K0EkYDhX
BPzsRMGz3oP/Z7YJ6lzLLP+ksZCWEZCvtq07i4AIaty7U1HFAHRxt1dPeNMARGDS
MOA5CC+CKPbUTpzRl8MwHtzgSn3vw8ZodoQIA3zTgJIoiIrw/vmTCKHn3Z9O0sSI
URntKoEAR8xTCphOZf45lkAwHh1zvfqHYkzfocbeWiAMLBbxJqYYAKvfVsxdyZQc
vqEUI6JSPUFfuxKMrOsA/7WXKMJ3zpcB4p85vH21PsqD5Bs6AMrtpzu2AhgewjIG
t6CRw6+5VWJat4AiNUXiLffYKUHrcXhbh7l/1ME6kOlG9DMBUsGMGC9ndVlSeOMh
RI9PXLWX/JPbszNDAnNVtg1ClxKmmQNA5fsA4tTc2ERPPkrx2+GSsC2K/WQgUwGQ
nmSjMwvbyQ5p4LAiwJQ7iJ/XPYISjAH67UJev5fhtODWpXuwxn/ua0wOjgSvhNpP
LArARs3CiqQiiXQgAiQg3UnlMc3oZKzwuV4KuhpQIc9L31algoKnYyZWmB/Dxfpf
VeUk/S0Hzc46ojoHs5T5xvgNoXzrBq50Kj4nuy+1pClNgJ6M7uEcvZJTttqLBZgZ
h4GscE5+B08KpV0wEKncfl/NxZjZJP3feh4ngzKlTdaFNjJKRCSMzU2bxt4SKqX7
3Y82OO0pN319YLDDDVpiiDKcnllH+SCWqVSFnZrQshOIUXQkHJ+CS3+AvfALque4
SBEJaEERQE8yu2fOFsLQeuHE+ahbJPuQuiywnJczybianH6PkGNlDbCLbfusyp8c
cfntE4qLZNrPQ8CIdy0//eavEcfDwd046rmaSW3Wa4IufjHCFNuBLKVQ714rurhr
UrZZtNeCf0eb5qIL433AvgTfUbdNg1tBa1qjH75O0UGS+SDlj734PlteLjqPIahV
FW7WgS+aSGx5jQ0/MUOdUINJjNbVTmHtLvUtL9A6pY8K336box5GmyTkx0/OpKDt
ha6uFcOmr2iTEAZtF4vXZAOqu6SIyvy40o3S07Ya4iz6YeD/g3HZ21yZSSoef2N5
bIdyjrw5dacQ1G4SDazJiE1R7h5faQG+sXImFTK2cuDerb2wLkyfqxe7EztBWlse
//vCL68/fajnrBjboXAc0TsglRa5hPq8hMJTBV4UwhCm1Cdtffz7y2KXK0FCojuX
eZSDgTiQ4ERhLncRtptD6EfEpGO9ZWMvrtf/LlEENih5REoVcwvsi8FPTz0h0T6R
2UB866SEQMaVKnGH4lLmiWdLG5MYFEJdnA1Rz63ShAGrWP3cJhMc5xFcFQ0QV1td
A+tk00HyWCAFtT4cIXx86Kl2UEVVcZ2If0782tA7ew5LIuiRPqH5SoxIFjPiXkRu
6OrrmyyMfs0zFsdf4r0DMXfLcRZZPmYNrwueaZB688Gk58od3HTcJzdatVBJxDVP
uXwBNNhmy4EBN7MNkCv+TA61Wuv6F/VlmKpFV/efNJsM5Nv+sg/5WKaJfDGflp8v
0KCyRC63MnnccYDqrXMTRJXTG8rwiVF4XPD+AlNASeXfiF7Rkravs7xF/fpTkORG
uUJFjrVFrD7Fg0K8fb1Fu96yIung4bE9UnvTVPAv8BpT6/du0EI9n2sEtPJgKLsn
LduM/CWO5q1EwSbgBFV5MXO+0b8HrCOZamCNaCI55tdGQRrS4zniwQpZ0mgDOGM2
9OnCqaOe1PE2hV7LWYmdy31KyT5RxMHJqghyJU/U+TFGArC0kltM1R2FkeVo7SMB
vSrpVnbILETHqcS+C9AgXzNchMmkdClO8bf2fRmmY4Eb+3l9eIxnx7SyxWopw267
r1GGLWlkaNdl/XxTJtggTCAPlxSB00scJmkWBundb9NJ4CCsjpQWbfuf1xYUxIxC
lHXdPX51/IM4iY2QZ1nAlvJqkhZV6dz52f07P4RRKrtjCNoOjCIUAVQVpfD4J0eO
5heu3Brb7qHmWGgcaXqIEmKLF1pLRwzR2vmH28nNW84agjijZsUjOvw+ob22lHDv
mONop4/TFA3uINfofy9wzKeCFrzj3zVCTgPy1x2jSnbK/nxZ+xHqXytniM5SSo2Z
MsmdDaHmf6f1BCicoGwpoBiPJ8Xlh6Assjm60TSMrXSFsZmRU1w736/jIQds+vwv
8s3o3zUsjjh2ZkA58NfrnrY0sWAGnymH4Lan2XfMqsYcOtAJlmI6D5kyfGLnUC8L
odmT/Eppa2671ajsYHI55rqDDd4q8Qj/s/f6N9NWd/s4bHMG3NGkDpGgYmm8xcCj
viVOF+lxlQQLu6BcfXOl946cFfdOtEUSeWhc1Lgqp7w5lEeZVA21LbBAlyAxZDaI
38iDV9bhZjgzS3FkS9m6r0jW7oA1cvHhRxeX6emdQPqvT8qeKehgxceKg7iIbXNV
w1Y48XTfCQMTf5t5F9F2Ra60M/WFCtjJxxC3BkJktjbfQT3YZqIG93iWMmG3qeLC
bwakYvGlB4KlSHk2PB6yJi4P2L8Y/WeLB4KiCxL0cqycfS2lZxfSEl4tREItGQIi
qWXpmgSKHekV8wW8XNFPHYv5hqgYiKtIKNhFTgTNCl4SSHoIvI/ckQ/GmIq1TX/w
hq5i+UqizppA7GgBnVPWaGMFMDwoQVwJKnIdPDLk/eyRklPFskPoucmNiBpszHHL
kHQxZtL8hkr/+2DNfts4q/rSK5FyilHGiJfDAvXq/EKLo/9IdTYRVxE9OBLwzqIp
RR6HUDB4VAu2BOwbeRirhWDx+SN/DzmyfO6LGPKG0yk584fV0scR4uYaZYGSsnj+
bplQV8NMyJu0Z3W88ml6vctXVLVO49wDHvrsk6VAWEP7l57CR15eyBU0Qck0pab3
mOWSGP516lUp2J7c+SzjZTr4btNPZM1CbhSltIcCpzCz9L8E5+tHrG7Jydgu5k1w
bsHOP2QkqqD3z9VxfQUiGB3yxbpvZGQOEBYIb8MVhRCVRYq3fVdpeyUH2xesSFjo
OrBIC2eCdAQ4Bj0URgAxHWEJeh74icKzjuHtMdttHya9D+82GNnz130CevdEWg0B
LqZ+rxir34esk3PZDjahTq85bxaCgdgCDl+2gajI1G0XvScyxyJ3mVPu0DlWsfkE
ZJ6S4nBKTfF46RpJN8al3o2fHIQwDYNlp0Ce/mjzP8GRxIWPannMfI5bD4rtBpbr
Sv03NA5ayXpOLoYu+gpfmXLFRhoAnFrc0VS4f9h6UHRbbxPEaqwDLMoP9aaM6x8N
glE9DVn7p58qFBshUhbE/GJzDT8tc3Uq+Z353I8zmenMcMTrJ0yZU49D+1i94rdA
+l2HidGq7a3uj13RxpzA+ury7Q+AKbalnE+7/ivnJrCus+w3kJL72Lnjp1BTXEI3
qMR7e40fEiuJ8LV5Y54xqFlsP1/wKpK2q3IN38rkvCtVybGhXuEbHLMJlr3Mdipc
vyfI9BnhK+lG9189G+M3EDriMzFlLqyG3E+2hYHbjOkmDzXhz7jDhHlPCmPMj2T7
c6cnEsmtcDXyLS4ukrW1i8lj4EHf2K4eVzyhM/ftUqDAtQYMoSo2doVWAlgaawzs
L8jVeJQYrzA0aUzNs4k34QcEOAlkb6LQI9cPicNeX+CjTQZZsYtyX9/OIW/SJFBD
acv30sGl5de327Z9nMM5t8kt1pP2aAfidktexhoRv0R5PyK47d7YB0ezITpomKM6
MGoURTTpTFbHd1d7rzS/5UfV0CcfCvR+EybjcMQF4H77sxiUFz9LL7SQ6nx2zakH
BNjOCOYc01CckgzgoQGHRADFh2WAgWwjJbdpSMPxaCegZ2+/YVLLeLDdqVMKB+uo
bSaMi/ACMDQ+/UJMVQEEWdKSZ9bPW5E17u0xEjPfJYTEe5ZyedRIOWebYfsdBFdS
+apzRoRPiK4U8RN5OEStT1aSP0QildyTBEKxoqcZiooPbGFluP6hjEcZnHQ+EMG4
cGPieaNx3sutmP2/ztDOMN0T0ik6GqblLGZiYqzvA9eUhQG3erbSlwtbNl81V53o
jOky32nuYc6sAwAHLoM4kz/f7NJ+OAlgnA6viZw3CP/0ChDxwQXG+fdsQ5O718Ps
3/caQ3RfoDbPIFEmkzHXGquLQJ/ZLiD4js4TPUxc8CgROsAbvUOklJu8dVgN/pWU
RFHTru2MK+Pqk7yRr0mzssgpZpDrA2twJ1cKd/Th2TmMmGs8BCZpGIOg8NxIPYFw
rqqnv6jmn83Ovicb9ZU9LvrTvhM9hwN2VSlp4dFch/1qYhzMAI95ljaPE9W7tMc4
zQavHZlXRibPDCpIrecROSu6+nNDBtlJsBRsYAUL8UDQUdNpOG000mAn3eqHs5ZS
Xh252RSWPlObMoNhuuaJ6vl8/mWrYGcQP1UkQE93QTp2RcTPTeCqTpTsq7u8e19Z
HC/WZWIp7D0jfJfn1jd441+Ml6cmSUuImAu5FuD7t0EW5rRBwMRrltuNltOMLF42
wGlXTHuf2EGaIGP05IgoPQ5ImzA+pLTF0Sf6sodYHzBUUWP2FpJwWHZvJWlZT/5g
K4e1ZnGK2LT7odOSw1S2lbv74W9QxKXmc3/8T//mPF6fMF1uWpFWI8foyvoRrDV6
J/UiwR9sloV0CgGMF5VLXE7SDnsItSi+qj/glksAKZENQzJUj9Ipvi9PxZZ7JSmy
rYyAlJULUBRim7o+2EvL1c0UQhzI2EDShN0rZCqj1SOCh2H8quWgIcwrtAFbUsNZ
qcaV6haU4JjcnmTTlHu5nvmv5LEd1QNjadurPSagTLTp92XPJ+D+DKx/FqI8Uxvy
r0cJkmS/sefdpJp6od+kbfkoipSQZ1QrGjGcOWG7vrl0EYczZ2kna5EPJwCDn2to
12f7aJGkEvuLDxbGGbNd7/DdzUnr8m7qwAW5u6hj8LZitbqctgZmakU6CLpBEiMP
rtCqYXM5bgayfehestXqUyXZ86m8eNFOXBbq0P7vSBcG4wzLAWp9KwDtDpDmbVQW
Yknk087zM40cxTvpgikBP551G8B5KBR4tCqipmuhjvYzxb/R06oJWVBcM88by25b
+Rf4CyUlRXrwiEWemHIOJXRk4Lw0NDBrcnwtCVbAZCb6G9hxQuvAv3KzAJ/pP3NS
a0f53hfWAM1vd4a2eeMXtB+l+c8pE33nvZv0hQtPV+yXBWAy5wu1qAdayaBhSdxN
qh9VC/j6r4Hz16BQTPO50CSfcm1Ue0cVSpvEIE+giGb7ygGTABxMhX9BIkuEFCUR
2qGAgqTN052JbBvlBXM/OXZQN1xAm8Zwly7RV3DKnPa16TgZ+xgUr49M3io/i/VR
thVxT90Knb40G+pGABqxf33zBwRoX9KvkOrxCMptGpWRudZVozvmeJ3oecLp9ML+
xS8qxQfw8r/KQBv64g3VibWVuoETE7LkscsUPSMHxGXhS1/zrH2TcRexHPKDGYQ2
3HMsJO60uKz7c0sG0ZRlNkOQuJ/ntgxvaUYiYxvCmYUJs8x5ZxvDW3hkUIQx4Qy8
jMAm2JEoeyBzryf0yM8dSPiG8rJovsMXvFcnxvl7knXuumPMarVThcxoXWsg1aRc
5qWrPu1U0V0Oxwhv4EaAgKGPaOd3oihzZBALquhyw3mDFZKcXiB4oXCURo9ns6PJ
ENL0BGr9pWpWkq6IY81G1z7yYJd0UFatwjy2g2jIFG/cS/47Ah6rt3JNax6zQrim
crKEUdIH+budjDNQh1iXhfw4RPMK3dDaZ6WbdEXftjwp5lTzwj4auatXKUhL3OGe
d2MBi56zCMl1eUNuqr963tg3PBRDDoG9MrLWCedowc5McfcUU8wo+I58VW86T+xs
DvPTVmd6sHOYJh7IlLAOeerbPURPzskMxDm0Er04r4fI4oT08rskDSZKDpKJDV9U
774NPDSnsV7kRkGcSx9bqOrnf2H2pFT+PbBCbJs3bmebCJ6sVc56xgwUE273CtKq
ZaR8Kg2vK9rZHCVk2jbQCFEOK3vTidXh5MptYwneEb9gsncTPNkZQ7n2qg2iiazE
uQKaOrtOvhh6eX81i0mygq4I3JhpXIw9xyXfxDKChCzEo6vOHyP4MV+bCa1Bw5Sw
hOk2xDtPddvKjbZG/pLLXrb/NZhtUnKnwdYUovEbMrnyDfdqwepwM4xE/S9ir1TC
OMrzTynCJm1JRoytHqc4SpZpUffS7AYLXoXRnGfqP+RI/bIxP5EyT2MNYatKOvdz
n4rZEH2NIh57copFT0yL+bdlhZcokd3Pbm9CFSUsHOvu5T8+1VJrceO3YGYoGj8R
DLOrI3AsUmw5BPMI8j7Gl1R+BlNT9L3O1J+7ipvKtlQZmuBeBac9NtB3z6A8UCvL
YbwDNQ8aI+olIsyATuOzj8lzSpbmSJ6KeEROAOmpye1oSaMC3DrBmKMx5T97gjwY
JZm6csXZDoNv3z7CEmvwfAUZtdZEv+bxQZ0bRXR16t4ukCbdyzslzx143aavkPZK
pBQId8QHkcZhsx7yHIUwgF300pwVJBXo0EMRjDW5oMU4zi4Bg5LHbIGdGLuJ/eiW
+6Yb4ZKxSCG+QeAtR7+TYzUgyO4V6fCKVBOM1ckn+KmenIEBzeHsG+g4Okt7Nm46
XTzBFobewHWGZf8XIleYyUv2FaLjGAsLVTBCQbbMtkvuzRsXUJn8yvk1X7wZXIqJ
qkoYmOtV6dYCWns8ktqj6Dupq74j7iJm2q1snPU++6KP5ox4KXfS4OWp5nXUQrR9
nOjIkwJ9WNffkCj/gLE+G5v74Zl3HY1Ku7/zXXW5+lzizXS0cPSzFpGTij6PWtB5
fEXtVdoc7T7iRyeG3tX4c37GsCy9RpgNGUPkvnOTZb6X27oBitw+tDByR8RymF37
2xWNP+Twttl5XodaDDQxU/9PfWr2oQatjckcSsHcgf6ue+xSvO4anVMYLkSr6fb5
j3eXQ9CbftVksdvKnymtr0KjW7Yzc0pufyO4F2PIwkH9D5+Kn5Cgpmc78W4MAzy/
dqO2Sqvi69umlYTwkJCE8TQIr25BOx8i6QnMpi5N7OCRbIu5ELhtuwhKvRTwNhtL
Jn0PD88NZWXis+Rf3gCAxP2ybOhYlbabaQVHeFYd5bBnpLcLU+SgM1bef2a5gBCU
UPSxPelDR8goCNN/chx/RJL3WijEPQgmzTG6xlYSqdPBOlO7IYUUa2HpP6uYjaJ6
cQg8nBImFoCv/4orVgZTvBww8TwqkFoBHlPwFEALTKjTHMVZemd4nJ0XdMDdikAv
Y/xJR56jJmQu8kYXPW0Y/CuwsaUWE65qxJrOT3m1z8lhG37UsAPO1xBSVSXI0RzY
smvvRYlySsaUvG2f21Ku4yPp20mx1mXhMuUd21OY+dcxmES+zORKxj60jBkPuM1+
J7KYXO700IdJcWKWZ8cH2A0z02tnNIBIKUeCu/SeG3eGpeWOSNbsaN5s4oOjrud8
pTc+8SReEd5OhstV58Va4JpfNmFjEPjSUMqJyOwVPeVS0PakRXH0Vcoi4IR485Qx
i2MQz0mdLmnFdU+OSvKa2rWTMnWK3gPoO4i3rYbdHRXdJDesPmlUbbn81JYg0mvj
NFIgQW4GZ6emBex9WzD3vk6JCPqBXfHBoMOXsE+PGfaLK+4CIa8NE249PpNkuX89
8Z0Wmoy4CbYOcU6e4SKuZtbcdghRZwBP0a81SIeatc4hlbA9LSS5wXWlcL2rDIQ0
RSRD35uBdvsa6BRQYBf3IaxRmCoHnrKjQjxRiPPpxS6bQphA3b0vNdSAYXCGL/7D
TZvE7pdz+WHOep/9LUyMZma1lHM3zqQgfdXmzCdieK/qOJDqv0VylEzcJWAcH/h5
WnFirWImyqypzUbqtpefRxhK12XM9imHvqgk0Ob25/MMUuX98lGjJF4ePkXugAJo
ovcUBdB+vSd0oV/8ZG3Xx05IBb8wBZYOHbG8z0Rimo6MfFYf5yKR50dr/5eq7NH1
jHEuLpobbZ5k/pIS0nrl3wBNNSetZc2cK3Y47tgsYtoW533WVCxlUKlnDo3dNOZh
rVBuK7TX+b0YFMB9u/9LDlQLDc19/6iccacHCeyLvKeg4XMzK5yJU2j+ZxNSWrN1
hbXbFsVT8OBXPCoGj8NsmVReAoccL7AazXHAAiezhVn4BW0HpDbQ4B4AWMwoIaqa
Gr4nZ9yg+Xmyct7sztZDRHyzYrpJUUKmvFZ6hUWU7E1+wX/UWi9d4PqOM7rEjqTu
CPZjIoszS1bVQ5xKcafzjf/qhXPAslDHvx5Xpc+SjRGZKSBSTz3D6fVaPIwKX+RK
erHvU1thLrM6J8N96dQ89zKfiKL7wC4dIZoYO3ZYQ6U9oNnX2X0n/Xubrl4iwqVJ
ET0a79QbueeAtwsCxRojYCWs8yaokmyEX2Eqo9RE1OFpcCwBKNbb13xC+6GzZrBy
FOszN4+nKZVnk80CviZjW9mAdBxcOl2YgoI2Fr2XeVRgpef0luRPp0XKPHcimlwa
zI6PBLUKy/l1mj6Z+N5q/mtoJOasOEjr6HqDddFGWj07hMjXUAMd1NAB7jt4pzmF
HN6YbnHcw47fyKEp6OGPTmmRCLUrSlspQjH+sbN8zmrkXWxPHNq43siyEFFa7t4e
hS2rITHQg8p1QLXgZqS7cNscjsLz2QEUVReIdVpg7r1hf2ISPeo+i6ydreShOn7u
D69TCt6vuOn/ZKsvI1X+BGCTaAyMVOcfGcK7bNJsBw+wO3HvOEJ7h1ye1HHd4O1D
f8nSfVIaB120WXCtNWf/A0F3426fCgvTEE5z+buFBM4Kp6uNO9ywM0WMouiQqHWa
95B5TqhKFHMKpEmp4Eu6opLbIyqi636j7DeYjdD9kq0XN0ipgqM73+knwUIxcqiL
xGZx95FnrnThEltjtccnSVk4zhgr1peQI2EDHyzhnjzeT+n4/i5S21Ye0rgPX/yw
kljvGBWJt5FKsrJyGiupgdDaXMYkDxBnlzpwdOuFBkWBruRFJGHsqqpJm/nAndnO
/7TsAeBDcEtOjVJ58H3NqkPQwGZNlJVmr9Glcq1gqm5su/c7ASxPETmXGE/OSMcr
5EMpZ5ZEVastjChy0DqS7EhuZMjOU2JLz0b29qAIbXmoWydEODb4zCNmuD1RM9D+
rqrNS7zgr1Lo1wdwCv1vr35qUZNy+NjZ8EpkxIPnn06PgZoS8i0YPo/W1F0q7XMx
Q1NFtngARRC6tjouHGrQyljPifsuFdJSsj8xa3MinDUb3yYp98MvMTXthsKuIlJM
LJO7oVPYNDgOvo1j9mIgRbRxbpanjbJPHq9FoFQ2kPd6oQps0focmya0aQqjpv4a
gibjRnk0qtyAOEf5tZMrD+eVvUhQTikgtSYrWhvhuiCGQ9CD4irjPej22U2HxpEk
FD+GG0QrQ1zZQ/rXeSU7Sm5VX6XsWx4s4OX4FyPKR+4LwptfFh277Etfbk7/hT3+
bwGAv35xNSwOjNfDx0UYVdndAAsM/I/CQ/YU1BXErIk/pk1QT176G6DafC6Ggc4J
3gASeGSj8jhvmE/U0MaJgoYtGXsZ4WSeh7CTfxgenoyNr8EAOgl7rQnvwhXwUtKP
6fstjxYVwA62Jwy6oZ1v3cb8RFoMAEGf2RUPOLpk50KBxi/M/Wom+8rIO+PBI2kz
HtdHLaKJ4yr90BFjyH277u1raES/mHKxFAtOArw8AVoH1hRZKY+vDCyaGhKfDvX1
pm62IpOqx56AJV+S19Fv5W7eSmSdHr4k0KNBjMleIDO2TDqbOcgnCSZdKAyERp9e
H+lJ3jDG3ByB69O00f8Rn1YZoi0fukgWL5Du2CjEVYANEHTtRvsKA3iKY/ZmSF5n
6LTybkvZhJP0paH28ReOUyShwFoor8Gykemeiwt16jVY9S4PEvstFiyrlGHk6PoQ
DGXQSMRHWZSMAsx3XlN4z0INyV4BfRSriR/FLvLEFp70X/3Jfjdt94HdzPNxiVJY
0kF1ExMFjKLWo1E+EXglf2nR5oi7RmyLS2wwh29SW3WRM9XYuv0FAy7ZVCb1ReR2
LRZ1ezgs4yUZ/A7CvDOwh5Y2uqioch4/5fKbT8HyRky9D2lGVzOPnlsKa4lmOgu5
SZQ9gGQpPoeSV1CXCLNJYXvaO3Uu8XupXtdsDD/5yej951Vpb5elysa8rR2jKndX
13/fAiQi7XlHny/4yOWe+tyD2i0vJ/0CwxTmGaZNXAmD9vJYr+UchIGO7iMnpQjI
GsnLznz6gxuiiVALWN0FNWfydaTIXL7s/1eYQSajo/7DUnlHpX/FW9/8QtG73vBd
C9Lz/WMya/ICu+TbBa77BkuhZfir1ufftnQKYiy44QlEliZZnRT/SoqQpqLA6FAF
3hS4KzJ2X3RzxKmnlSAd8eukBIPZpw44YNVVevaY4SqK1x/BOhHC1jVs5ORwRYn0
nbPhM27Za76CEtANTkpw/1j6kxsy1Co5xGh6pOK3NVUarA62h0Du51NZ9yvuk1mE
Y32XS/C26GwQPsSDvmJAkwv2/j3330y7vPiOLpxrelsLubZjU7JnuQTAbHAarKLQ
Tktv+SGXA1CNwYyCm4BVM/Vv/TQI1U14EnfQKOOQpph6BTs7RFrkB05uD3bkLM65
er8zOqVTW1HhtjCcrFFDB3bilfQ8AHox2kSk2CclDre+AwAM3U1gd1/YMQMeknJH
E4z96yc0yodHKDPBzlla9ziNGiJLKkCKN3Lg6lE1kW1vBuZYVTHsTK6+PTuZua4E
J7nwuWrhVgdY7cdmmiRbJJAUQJfLO+OtLHYpvWPwVUPvRzFHrE+1P9K7V3+GG0S5
njRFRg1rQvyzCEd4yP1pR4K6M/XgEBrCkIPQE4RXDfJOgVWAveLM9qpHh0o6BM5L
j23t6wdGFabIi+ox5z2+KV4vgFleYxuN2uD1rxLxda/oOjMmpefHwBgjPMKt1ALk
DUI0KfUzTgpb0Gl6fomenzgSB5VIhHIftHz/NmgJ/bExajewJ65/Wdldl37bDQcs
ZjmdvXd87h6lfXxMhK8b+jGqMwqVfgm1Feu0JQntmqueRzWtSgB9AWiaQY4W76Q4
mniihttsybislxaTCvEK2KbxJu86JWvMx+2pEzySXMDWG4NtmCYJQI57Q25Lf/vk
neSzVC0+DyfvA/aBEuvqXAc+Aj4x4j0XTyw42h0wuvSD21fhUDGVEVdh36lx+sKU
gYcYEow5fRKHWq5IcCyR5ieBqtBN43Zwu3Uoi49mWWCygesHF+x1nSSLdhWWga1W
cevteP4j57ff6OjKVNv5BtA1i1sq+cOhvD/t2VuWbu2NK//ZQuJnxEdl0Z6RsQYH
fbAoJhLypm9vZTbnOqcOPSmr9yeiM7OLMlNRuJhdLtg8MbhFMqSsJdtCpJejLXNw
FsZ16Q3bBG+cDBuyy2pyiBN743FrEhTapz2qSwnxcUBoP1QryMo5/dKVLxPJLqME
9OlBAUSoGOJX74v4fe7nFkv6kW8Iv3HHmsqg+p3m2onVmzTd2Y6VDHCev43GxIpr
+To3Nh+dMeiALNff0PW8P+3OAQ12eS2vkZoN6n/cVVZdDQZhdixS5J1wbAFFhnaq
Seo1bEMfzk4o1xiHwUI7O6F8Gde0cpzw4ubiJUG0GFFsw7YrfSQXASiEa7jW+D/i
GStE3djHwtIyc5FZk5H2o5DU1ihXpNO/fh2wyna9Y1OjpIe51BRyW0hiMbNpymT7
bYpbJmJ+B+fLqV8vMkaB7pVRaeBdKPlqmGehu/Zj4XNK0NT7eNzG9FkAu2NJrawX
Ay0Z47l+84u7S9fi9EXVBjnE+Qiucf+RgbElIPN3VW2NWUxVFOEUSX12BsaefQXB
qL6IBzV7GZ5QRolfvkv2/+FGBMXkfXvaYhV5tP3slaOB/v7Wc9kkoZdvmkzQCMnP
tQrM+ib0HGKv6KrKksBrZUOYQISpT5WNyKjtzd0KqR3dvAUWdfHmZEDxCoDMKL34
PILE04FyD6ae0i+q3vX3iqHlI2FbkyN9qL9SNtzujLLo8bWcORPKLIn5spfNOI/i
G/w1sFXIrczVYOneCqzxheqTG/uJmLWiOGmeMvle825CDqQPcAOwKl4mLw+wK4Ql
qLB3hUxhy9UpLiVEMZKwyru1S9fvxXhWMQrNb+C2j5ZkIQyrLygUwpYzXZffqle8
BzVyEpavfJp6OpQgt8PnjEGy60pQ/qdqGPye8SAzvbsf0WShU3xDjjrd9JT0DSY7
AgH/hcwspUmsqRQ8LXrow2cKsy0y18GwXcqBykVypOLsFHiv3UZBaHCYwAAopdFx
2zsTsSad4tZ4rPMLzlH8OTB8nC8g+cjCDnF/QZddjXdaayS6hMtx+pwmbwGV0Al1
dGOXApHzlOWtc7sPwkr4RUAoRKu/mn/SHTQ6fGa4DBNQT5HiiZ1KOoEfaEg54aE4
+6v5S8jB7EyWcgn8I0YMzKIHSeD53xbMfBwt8q3wxXc3YPJD02ZqhAj4LfBwFyWy
RgRF6nGJj9BqmhkVypUEqVTdttnJiX9a9DP+cRW6jfDdWfHNheN5kEincWuXCVs8
9tZRHZi6hWA/kuV+gOsqpLIEm1JlrfGB9F3k8LTuN0Uw/t8PbNdwxmGaNgI6jn2C
rKLc9Ocdzrbbj60QbP3RO0PJ140LZGWU0e4D//tk+S3FSnRATPLnlhezsJcfTZ6m
6aM6WlkIRDDMC6mQlW3oLM1jcgVChyX4NvB+oVoRIVyTkP+9GdzaXnNre57NyixU
Sli10J/K7V1oJ+gtKY/4Dwnou2ntQSSgOiaDUiUqZ6nss01+S+QjOQDkJyc9viaj
zT6aLLWdVqUAa4gtFk1S7zkkI8SyEMSid9YZuI+aDMNMD2IJATLtculoUI18PT/Q
PTXedQVGJ80LQj46WjlVqbtqQf/2rMHYBE/+Q106i1U44+CiFnIdKRJQxk2WCtYm
f358apGPB+b1NrvXam+luIrMNEHb1PstxSxwq64/9c5t4a+gHU4YtVTBor/52B+j
XVMS62RFdU6dhcBGOgKyqpeTrBQgS3GEUxmL2FdGa6Xvt9SV6hAkROiCFNdkanUf
ki9H3l7cUV9bDZAj3Rgo1k6wiBe/cPo8Tm3DT5iGF35esDYGEJiE6/AP/d2qqufN
SXAfL2VwfoOw4VInq7XsUayjJOaR2Cbpk38MHsEziEaTScd38ryf7be+v/xDh+RG
ea+qP9HrgJ25qT9RGsEdNe2McZBiXzoxTxIca0OhC89ysmkznVQL4otxRL+cnrWB
jX23s+05Cuxu2ntMIs1sMucTkV/iczERgiAvxkyymMx2eT0jfkiV4sXh4x0qNP5A
jH0TyMu/x1rGxzRIVWnho+zGQ8GxyM4RXJUkQpKmvVF0cyS1VGkI3DMN5yTpjVTC
yj05IarQYbjx2GKPP+lkF/rtwknc+0wT7vcntFfLjLn50WgI1JTBuR62EHaq5U0k
MSbP6WZqtrphElL53zndUgHC+ZYppu2ZMRrksuctpXzgCrZYKTb1xjbd0eFZW8h9
YAZ97XIlfX3tHd6EpUeTmA+I3mUho3Q8lvrXshAyb1a47aL8606wTUiG3Q0y62Wi
Pu8WyLIzt8K8wugXsSDuFRT2+/3zLkuSFAnxkpTov4BhrTrR/OaWRXt3XNOstIcG
s3gXsoKysbDrh0mPUt7G/o5m8mDI2eyBTmiM78mOaqouimn9bavt3F2Wuu/ZsOpE
4sKHh0anZy1BkzaY27c+b8lQHLp56A/0lRaTNee1rRsRnXSOVZAHILpG3+M5/F8g
t0NS+5aaP/sUxEkshR2r1Z6JVlC3XqhJOzAPJqTHQBtVs4BtpWzlouPja98T95Iy
AvRbQ0Q1G9zS0tK4WT+Vn+s/pToOIFPTfdq3VLZY+ZZyS+ND8HHJID0QrbzrB442
aNP6GC7LLUrzkuRZwuWI//iCOzQR10PU4eT8FpLpTY0ymexHgSnXZX3IyKZcMEkE
xQTOMiS994eEIdtaFRw+Uw6w+/zVRTls0P6uyzIHIcJy4EeeSvgFAeqqlSKu/oyC
JcXQJA4jn46MABDv5xL1LJGJr2Ki0WSh+MqtyvqSBzNEXuXH0FoHLIEueCKIigyb
cB/uXOcDD6m70vy2wp1uzYxdT5ibPQCh0Uu9CTHBc//F5bnEVz2HwfRZvy5nlxdq
I04onB0AcfP0ujL/KczcpLQ3e1lC2YUGUGy9WsFbVFF1ABtVurw/Cb7RsTaEn9FF
oph1BuREIt+y0k2mtAmAPh7lL+dz0+DWOUP7ZdInBWM9c4H3I6E1NcbvPpbIrjyT
qnN76wfEdPtWOBD1S/CpjtI4MJs3pul/J94rj1XMjBJ+nvn/E5dWBFk5J7qsnw8y
YhJVH0CHdng1aDMlIQnNEtJOcvJY8LEt3MZ8SuTXi7f3QiQA2cqjcUefOC299s93
BU+rvqtvrq0/TF4XF3d3mpWfqlqMxY9QX0YaC+FQPkPUMKNvyyiYuPlk4qOnh8UL
7BhqyzOvC4/WgBK1qUUcPO6bRLmgJcC2l3Y4CmUlx7HTRhRSdbiKDxf3Q6laax17
hASLdMXuzdRqbWgHvnklmjtpDeoa8kPOiv/Ej56KBVA9WXEe6tyHk0FlR5ZU+qCX
UJ2mJZERyYYywBBcHH5tblHJ86Ylt72aEJFFxrAIaUkjEmclrDZQOyiukg6DsO4b
gEP9YDXum2lZJZRXIFqPawYqow2KGp9ODlk2dridOCc1xPcYhSefPibUb11JAMJL
dA9Iq5ioUvnWSx1jr75afb3IEzVrQqjRCS3F7WKY+Nw2yN9RKTvIuq27yvCRx4a0
5dY7g3KphkY+J1JCfNhuiZdcjYQ7Gdoro15jCf67rQJQ2xjbWragZaVBVtLok+z5
YdJaRZbAHc/lkibaXKV3WVP0Qu1C35YpWo5TiVVaxf0uAmajuA1c5lM5JZ+IbKpR
BjiRbS1ZF8htdNiFHT80y4MrDNYXyQUBZxsa/OCfXmhxHbUslXCmYqvsLJ7MEbQv
ele473lsfV0j+0wzdHu/bgj/1/G49L6DEzq5AdL1584kWDq7Bsa0Qe49MKRvkUQo
Qhsq9TbnXdNwwcT4ZiTMpNw//4PkwG8tuyZgZTZ3MEDD0EtdjMeFoBdQQzHea7ls
0ki3eDHLouOPYzFMGI15NSvChZcnxIBOTP83tK1fpkI4rj3XrEo0oMBdfUvQeVWW
oZ8/K02b+iFOtmyizTY1goU6ZDGnPnW6RY0G07+mflvin1ni/pFuifohn0h/zP37
bdL6hw8ME4ymIovi2e4HozP0a3jbnZ145uVq6StqXPd/NUyW7V6YX8ZlQOsx2rgh
KTOOaPqr6JCBi1g2jx15gaG5uuu5PP3gCoxcNfa/QEAbDhnGYBFGXZmSAB1yikfj
ysukE4n8xrljFrjtrtggoU2Av+O2YApFgR1kIvTYbDt20tnHKMVJ3DMbZEXaNE2b
ftRX0Fj+C2jkvCN+kNksgt9LHj0En40Uwmgzp3fy513r3TBdawfaEXjxOJOZ+kLu
TNOX/X82keduvlUynoFe7IwqqCbOOz8jmaBtKEvSPkjieLnsyPIYW043QKeAcfgg
kjFcsHf3A6FoMZhBpImu7bxOxuQWV+MXJK0BA75Gb1vWHtoaoXY6IJ+/4X7eDUuh
DAUM4xH38dQHngGIJ+3TDs5miXNISBU4NW7jRnAos9Na1JK8bE+nNTq4wLUFr1F5
9SLNEVHrcJ+YRSSbRIuq6z08KI+GhQplch7w47hqebZ8vyA/RNI7n1XV1YGq3RST
rblukZ4F5fl8fFYjW2Mk23QrG/V5O+c4esBFVwSyh3Cb1g0Ns6bj42Md7swYdLAT
CxxWy3pCqe1Q281Du3wm39JxAXciOIL3mzvDo6XQjv9GDEoNVO5jawk00XBuHuvo
JWzN2lxieJvxHILX1Slm3gIpTzwtFrtx7rgeezmSf4FQjWQels9SYVifwEHe5gdk
gBb7YERl+3H8fLmn0KghKhSdvXW/oam8wQaQM7MSJsER4+0EXuiH9JoTde9lsesg
ZHUP12ko1wZy5HBeTZG1msm5uFjtwNFCIIDWCz1LyM9k/3VxLxcR2hK+HAWXYudi
1wE4+xAUMEMhq/igVPuy8/a7IasmyXMVInyN38Sg77JRoOgLdw5C9HBQoeZPWWVC
mQ3KnAXZ4oWGkaSnEUdCMut/T69kbIXYNFuV5ASrfgkrznadZiKd9ygh+bv087Fh
ntBLlj0d8fKlGwdK/ZAaMGp8G+0nM1CedDx96WlrDhHgoef4F/3xKtW9je4SBQkd
G+9P/vWMg7TuLOsk3bbTRaz1++nNagvtVpgnHg52+SLNfx95e2HqxtobfQvtikmI
rURgj+Pm989lXdecRjrQw+p88ySMgJdw05n83Qk6hrqNBExahvYBY9zpVsxIZhqA
IOiO+ifXkDaNgSPHEeA5XrdI52NpDiiu4K/eu4iv6dlkVl2u40iQfwia4CUl0DB9
iVSCbKVgv8nm17ZYN1eRsusF893ZL+inzvQ/quWNVe6k0G8+lhgHICVoBWQ1xB92
RInLCDIxV2LmkvHeXeMVenz85pPv6DeP5EAXGBZwgNBTSMAJ+Is646p+cbqqFM87
dAkR1lszgaZFi1uGBphwmEew5XL0Gmzpa8fzDkfGZvCiB+9F31i9fLlgeaTRaLjb
X3efnE0J7cu8DAcPozcpUl32SlhSix5cM3bJLRp4FA559IiWN+7g0kHpKnOcLdDB
azvIEMa/ys+Eu6ucSGfagoVGqPf6xDO97/WfBAWnCbya1WJ5ugjqZUOpJv1M8kQV
7COhpDogG6w731mMcCFnvsx5e3dNdwfGhqbTKtpuEte7Qum37CoGJ/HuPehGKJUb
wBO3/jKGZFOEO1qKqdPn/LTRsb3XZug2rrvO4fwMMIl0oFbgLMsK/H2PSWBpK+B0
X78c5SWC0rXzjN86GjLTf+itJ38vhUNKVkLlJjDAueMF0BGLXB/l722s69hVJIsW
L8plUlhYxGrHlRVtc9KDxTqEbEozFPkSytpNbmCONHQuMSirUCaC9o/+CkT0/9PU
8tcb3IaGzlLBr8uYX28atvTxjD3aEycuP+6SAUY5SBiT8fFeyCjSJnZR+cMZGLpi
LE8eZOx3Yyhlj7GiocUKf6asp7eE0YR86+dZLAHIk8EGqMOQ/HHJ0D4eQamAr5Cg
dgUT3ZtUgSuZCGp3bIz6bu0/dYgWTESVTB/CXt9bu1eVBSu50iDzR1qZqsV3Fjyr
Z7B92fv9Af5j6EI6BFVAh4+HZDMIs7oq81T0PXQRlpVIdlsiDnYkfd4tKaxAoXek
DVxyUTjfACtEVKqIKI9o9zOZWWBtLyhWzPi7b9CAguQjXDLabM4LFbsECL8mHfbz
p6CPttUhjnpQqpFebOTGhPGN8h+sMIdyLhCHskkZT07wut8froxQPkXRkboAoMdg
IOgJrUg36OKTxND0Q2BifZOKRYTujnAMyH68I3xxu75ncFH2WCynQffuKATSwPly
AQllg9+9lim0Al2v6UhHBQ/cmoTwfSwlQqwRGl9MRQpePwEcr6vQaC41/YGBaCOt
/gbR02/Fr7VmQa4QwNIZtZvtSvLbFnJLFoPVfT7cBYcQwst2WRc6h3orWoZgS/7J
vinI1oJXu7fhmlv8dxZp8VyF/FBz61KlcI3epoN6bu5zQMmSIL4Y1Kd7bWyDX6u4
oy0LVet2o5M/Er7mz0VGWeaQ6wKyz2aUlY3f8uTEKSi6/JHrOBRoLGu8ZNPAXGnK
ZvverMwA8azefGenEuVLV9noTvY7Zx9ve3L1GiRcXanomQnvnqINQ4mHJahsCTVC
X5NZ+mTk+u+VdYQzJOA8vX57/S/f+uXkpKu7ylzl/v4RXHIcrhKogmrjetLP5Jzy
DytXWyCvdCCaFpfSGzXfdgLlMoR+CyzGP1giubYco7dzG+85drflMCa/TJOkJAuM
JGWIavQ78KkI/i/QCqWp6dZjNW3QhERuHN0Jvut7FfIIGFoFin8LmrcaMxA9oOeC
JYAanohKP5Ibc8yI8c/BlngIigERKST7rOZh3xN+D6/YPbnA7zc7t2fY2RZf/+x7
tcck5zXHyTRz3mbcIA+JB501VVRJGJmq/vhO/PJK44VnNRKyyoc8Luj3WKOOaWwy
1zL417DZc0cIvzHTlJcvvDeSPyw35AuAKV5xtY8uPVxo2H5tfvjmFRCcQUc8SXP9
Uiq5tLRr63kvEdfj3uof11J17QhY6RL7TfmBF7gHWDP2SoPY3KIcY4aoT6TOr5Q5
PCINNdt5QqZGqNTNPYBJpgVATtLx3L8fTrHnz4ipa5D5EiVKP/kOa2XIVGingQXr
6LYL2QCejVLd8ekS5ozZm/XdsB2GgSL/kzNMTAk0LsB3D0A4PmR4BR5gmk+4/s4J
BvG5OOkI/p4NsD4yJ9tItFXH32y7SsNzGSPWQgT1G4mt2VwMo/yaH3uQdvJvz/Vn
4Sat2OSE2BSVtjVjpTN7Ils/EJay2dsd/iyyt1HVqWCSmsTGQ1wd1cnz7L7cZCOH
Mmr0/Db+5MfctXFZ+WGfV28MqjT7Y13ibxdR55LVo4vOfRBUYbK/mb8qj9Oqs247
iCBt8QaaUa5/ddKkB0fqn4BK4wo2S0YrC0MHpbmFDQ/f2K73sHm2kpYznjPmBhOs
HQVGmET9QHKP1f2AXQ9oYVJ2iwPiB026rp7yZimCHMsosLKtjjOVXJg27hJ8SW9M
XNR8ndEacXmbq6bxEDz1Wr8mHJWfKo3TCM7H9vj7XTMSotUc9VEE6I2zvGQ7lqEi
b+voJV8VsRpay2czW3p/1R5t1nUcmBs6CEsDyUjXGcmh9F7tL77Pjs85FEBvcOiw
d7cis0HeXVLkbUs8cbi31T3tg9FyhZGAwPmM+JPnLij3Gv8TBFnfwGSkbZeKd04M
MQKG9vLYG0kBXqsvKT+gtXFJ5dkrY0RsZUTxWXTqTY2473wHVUqjQgMEcbbUBMYl
XnGVdi5TLjrUO1WSG7j1n83+OYp4nkwPQXzI9svCkOqy667OzWDFhaS2zu4A9v8F
gR7rwIYt8xtsNJjCkyQpZ+vXqz3pjyqqBNV4OZ1t4kcddv3mR+FF6JCPwM8xxJ1h
AcKhuX0JGc0gUZ9+upXdxLH+vowXBWcJQkoMa9ljIfpir+GcsXKDP5m2lq70WmGJ
mmnr6PLFV4SEwlDLzJGvnegRwe0N4AUXP3Z9pLRT8xUwNjiMPyPmbwTGYNn5r6Ze
RNJvDygz3TIwQfsLS+kazZm4YBjNB82tD7LWVCAsHXFd+0j6w4Wzmx6VnqSa6a2s
vKql8ryy1AMho0AnTwYyIF4UWcYpX8vCW/FYHUgKoeih6LrIzaWOEZQf9m/toWxt
aPPaT/dIexm/5BZfXcWdEH6kHVd5YVVHuXKrmRTBvTMWUDOzAY2BeH1OfpD7jWK6
UYi/YYqESgXyGOaNts9q/F2tYnIFmUjQa0iRXP7dWeMH0nYpIzdtdsLn6/KDSID0
F7rw0UkghCmokyvNZ0B4/X/yZAYk3rcsC5RfmStdCtlGwVKQRffJ+KhHcW/yN9jO
9cgsWmi/uTdtQyGc6Y7AZA0Bll2fqWdSEdAZiXhvtLV2UVvkwUHpz6fPcHrPN1d6
Uvu+YUDowHwSPO+IEoYw2ZV5HWqlIWzPgL0R1jrrTrcqSNI1s1Ti+1CVxXT7aaN4
69LUUxHe1AxDlH7BeAj8rQvuDk5mQ6AzxfklbrzZPWmSXTdHJgHtmNl03pHU3SOC
C4zd/WclqgE2DpvWXj+l2s1B0Ocx3Gm1q9mbSA7K0V3ntcpugZeXBfVQ9JB91/rl
/93akgbhQg5dYxV/CpzPmQthAXtVRFwM/EqklWmr6+tdjVKyef0tY314pEgXCRKq
X8MyniEzejfoASDf3awE/MlJpsataPEsuIT4j9GmE8W727I62qj9eIUNfjPz+Kv6
WrQgkTVrNo5vxOgm1DxjXtSF5itoks0UfXPfGs1pnuutyEYRF/0rvXJbnmHNUWR8
yD4qQsmzcqYmy77tnADo2EquX+tcGNfurQHq30xak+t1RXbUiNCtM9qL7ampcRuf
bCnAJhEDVfRGDdKiBZmLrOl1WVhwk+lkBJFShhsumo2jVkiIld71hEwtbPX8K/1t
cN5nB34d/wgEOKBGRoRfO5h5LRMo/P/Lft4JEfiFmSKXNcRZ9RaK9XbOhtjHR75c
VbyuWUIIjTlq8enoI9N5bUmTX/yV2PHkMYrTL9r4FGo1dTfGaQ0CLuhPyNb15tjQ
Rqb0G71+6eq1XICl0Y3jOX969fdHkE/zwjuBtQSGzAf6RdyNGhTixqUBrH6/PpeE
MzSDdJOwYIaWlJfKKAqcE2KLtmwgwY5XaMzlaOIHoDAx3QWoG59ck3MPcOnOIo8t
27lVDgv2L0XevgHbvLu2GurJpVyWEsArIGLCBFtZBaC6CXwLkAz/zujNm/n0VXS5
nvls/rpenTri6QCo26D9raqQkPk7PItBI3dIuG4DMFyZ6oMp/tbxhBi8SgxFoQDV
tvugHyCKK1o7oTSn/Po9lX5YNTFf+i+PfA+zqlorQqzz9kkeADWU8jEl60wSLnrj
LkZHOy+FtZsigDkSKV0KN+6LiDiCD/gFnIwAMLOHL99etctcA3I86kdNUFzONsi6
fNiy4EcuwKTG2KKpv/SmL1uutnruBjiFZBnCodj7s7sjljXeFCvGTBueSggngQ5R
gy2QTgw1PLFpzMPKZ3fmvGTFHHS8YeIrE/iufH8zAxUn/yxx66o6JHMtsTrrVnYk
Yn7y158Dhorko5pfmTBcryV/Gv6IcfU3VBvpJv8A0b2VctqDkOHhEwX/FfFLzdsG
/fQDptutTW6K1+7aGM9osRlEmSPmq5lVbu8lO1RWEf7SALRTQpkkgzAdch4AH0fw
uYdKQOn7lx1mGZGGLbXg16jPhpfJln8EG0crWc2Ebk5Sr5r5KutQ+crxZ3IU5BO8
THbSMcBnUS8WbnxjATnoykemG7czkeDaQzALUfQyFbSmKD09xFp/TlpmgT0zz8Sx
ptQcEw2XBATGMxBJePaxVnqHFnOUHuvRsCq5tAF0a8PQ4PHBhgvcjjuROmGBSj71
sxduBKUrZpExDtMRcSACMU6d6L9kpeLK9gspfIxvCnA3k5Weg8Ovnlfl62K4axis
jJ98krIPuubsmGl4/+oNLasWBRe6HYC+em9nc9g2tdtaEH/zhcqQmTBKF7TwrMyX
p/TDWYME8u4vqwAIIymdbCSefbvD2TznaEbt08rbF7y9MRX0E9r6I22U/1g+TazO
oKUnqIauQsfQ67LQYTE6C8JfOFdiKYmQfWxCA5z9cnsoB+7Hljz0iFB3Ssdbufhr
LJ6LNUYVw24zLvUfQ5dLCfjhgZDnAeELVE3gP8XVneOoymIMXIqttCCzBYdjzj5v
su442u+4TmO/xDEaJPlBhCiivWaupQIJKfpwan8jtfXYl9H98xum/fg11fOFRcpa
kkeV799NhL+Oe01lVQ9b1V/7o7iYmWt+PeFtzTSBpxBFeMJ7u7kFci44lsL49eE4
c8Xdh3qnT9Kh5SHLM98CSbCiEi41DOrgs80bhxMnt4RyP8+Ejaul1kdq2xf29eSx
6tjxcIVG1kRcU9/Hms0LeAvXUfNKIdcxr7jJ/wnECB9LOaqr1bDE5+1Txj7zqoZS
fxnd5ijMHX8wsTfD5W8pnzQ487JBte+7r3b2Tgwlgaed019oWxVlSrJmv3wfdqZF
b6Q43YtGF+uSq7Zpt3JS4R5aInnP6Obs9bAqxuzd0hZTui796U2gIJH6SgVhhPkn
zGQFIzXwcFYHS8YwznDDH6IJpKQA+iWlOd6bv8Tj43yT2U1AIZVG3ricTDOCow/6
l/zmzXnjZBSD59BFnvNatm+COWNJTBDHfX1czqlGGJRorTo5/AOk5MPW9sq4fSW4
5M0H3JJql8QGeMYYrxBnA/82mtGrVCrUCzkCgm4hpOFsP1XM3t65hH6on4msM2ij
HOE3vkF6gvtGq0KvWPhyMZepyZ05qBO2xacoTMXrZ9OJ0SjLH1tHIG+wI72+i6zq
Cb+xdQHLe5p8OkS4pUz9441W+OMV25QCEXNuJ1qvjqTe3RRFeyF7ABK+AcotzalP
otTQilgFnjq3mPJ5HDTYdFI0ZiAC7SvvN6i7gdX1kFEB6Ga4OIgXK7XZDvCp8RXB
qhdZ+EiKc68H6xbTcIHsQfJYc7ajKX2P6ppVupw1KclIgvXSCH0Qk351MZBm+VIU
R2M5oaV1K9InWGghJQJIvtEyZ9FL2bmfPUknss9aYdhZrt1PnmVoWvcplt5lihAy
a1nrk0Km7Sshm4HTka04fW09opEmpAIEhKRAw5+HBy+lnkmzPPW87vJDf26EQC+P
gSm+B52WcgT2rY5rn5gUDG/4UT3DO1mv8BpopmhwPtyPf5iJ3xUz+MaO+rdFCAnK
4flvCVT+r0LbEVuuvUrXWOixHgyd+wupwudo/oh3vr7D0kC0V8Bsjld9nSv6ZXC9
u1yxtF2nKSA7rMeksXtgFbTqNVmtIdbAWhBU8+k8DxWGgoaUNLCTHa7yTARlggdy
tj7qvwBjxYLOaKnL574FlRIDMXPg7t6TKLMkXbQkY1txOzBrsL/hLQHXhf/6U4LB
h7HwfYwa1EC1upDPp3S4aR47PyjcC3vO2UDynjTsGknOXwFSXP+i+X5rgRLODojJ
4i79vvaRnws9MKx0s6XvF5Jti6odKde4zZCvXckVatqpv5pYaj+/0OvkpNFagJI2
rjuRwACy/ZiAuamuwpxTunWjQNxid57T3rZgxatlrU9s0Sadzq1PeNmj1pLj4kZc
DrkhKMI5bJYf9xVL39AZR1ofBB1zYNbV2nrQcAvf1vh5EoRfQzRDgYeGYzADIvRS
cjpiR99S9lT8hDRsVrdgn7VnlOd2NlPlEYstd89VUSo0/IJj6+aqaSdlh9c+rU3v
9Xl32Rb1PB3ZVhxOz41BDao8F81Iv4tNfJ+FO1DJf5GBB+ND+r9QCZH3oPkVZse8
hZ1cucB6BBOHsbusmmhziQAgQKHbktCJbMh1rqqxGZPUFkYvenRSk4uuxSE2VdwD
opQaNSB9HQYQqHaH0KPCENVlCUtLkO5G9HElqBowAKEZKKVepeUGmrsXb6dANDPz
1MEk3oZzwZXcmVvMJmO3VzmO7vUF9cCGmCUaHv02C8Qc/xQcEYLObsHF4++Ki85e
k3/DPNM9SCgLgHByg7m/C/52GGtSUe/tmDDgeLihrTP0HcRlo02BFYqyrzdnMboB
bM5a6+A/G+G0B8v0PTeWCMYPdiqHa+GCb9nnrORejsgFSuZTsyJAaCClwZ6W96ng
1jwt1onheLHZjFuCJhVVhNdxFJCrXcEhooe8iURDaYnsoZTJSvKcPs4h62dwAW2e
EmYY1UNcQhodUa2UYHwbfv8Bz0Mq10llTceDR9Ulzef4pvDZmiUUwgnl/ixlTFrS
n/Ik7ef18XIDomWR0tse3/9VzJ7sU8eAypJAPalq57hsIaOFsNKsB8c9/Vr174vR
A3qM57A1d6FVrotcQUQPvYqaMZNhWeu695AJsilQ8Cmk8lJffwpO3oTx2Mf9yEp9
T9M2aikccvdl5bOtQoPYEiZB1kllB5prplQfXmwE/82xc++U+UlKhmFgP3o+BrW1
GG4omUmsGvG8GUm2Mx80esBDiBSp2fNrMpEp1pNMAW4P5Dqjogp299kTj5oFRTIp
RaYid6ijwe/d1oDgGz9sBtQE/gMQTMJcW1FmtZ6Go9txi+R0c0il9iHnVl7pmOji
MhvS/WkHWFwVv+ecFWmJCvmiZwvoVykghRqbWQGx3CXaGagPEExKa44IOiqD7snF
NWcq0c/KtQL9W3Q/OZX04/6JqZx7Ih5GFCH6TVIOEQvDoaoXToCa3sclomNMKheC
TxUq1svdrXSEaGQJyIOeqGuA6iy+GEtzOhwesqHTR4mJSLyg0HQYaELUNJ5jzoII
rpYQTeRqnwLyXxM0iGzL9eh5rUgQ71o9Cd7Y9ka8gLIuVKNPj33XItbh58JBYwYM
udCOiZMcOWyG8YOwJHqH+5N4K8NZoz8j+MFgLyzJLSGLCJ70rXUb0CsvAigVTPLA
m3NBTL5duTpZtjKRMWYHgRmhGpwBvrFMEqYDb84Q7nDX6ee717ksokGSF67DvN/W
sXZzj+BfM6gzS6716JZ+1HgkZcjrCFtVS3Dw0nVjPyVk0aeMidt2WLOlyhW5HRoa
+m5s09CFoRpMT2s39jGpvZyTqSR5guZzyIC3tPcvkCubZwUu5cOsh6OEIhwzb6TF
p8y7izPmoQfw2WfYKm5wovDVm9sMeEHhpUCitJ0LRzHJuyuLCwvffnLs8dyq4E7g
BzObI5Q6KOTOJ/YtcqBNPJQpD2kFF1UgIoLJlotmPJHuKAX3oAx3lwgPpEj1v7zp
jBIU10IDG162hnfOzxxBf/k/kmx9r/w/9ZdsDYq0cmlBBCPORQf862Va70eTh6qo
VsSdvi8YrvYzAPrfq3gL+kgDMO4tv9++bn84ClSk0fEwGJ3UahuTUCbeEWjiAl7A
VVxNXdWTttD2usEPj/ZwSNAryjno7X30jFb32vXNRB0npo7kM6+PdD0yIEC/XfNy
v7tZ0+jSOzKU2h7eqL5pLdAVmneWX8LwePjToa4dFde9cU8XK7t/j9U/1m3sycJZ
P9zjmzOREngvl+ZDs9wZEVRyBnnNoR/1ya+eZbEUUU+IO9YQcRXDQDphHUylxiE8
gqsazIZsceDmhVgr1G0f1qYEUYIwIJwoGAShea2GcIBncRtPOnBmZUsGv1iD00qK
eLRsucvVLNgfXXsCG9CTWfBYY0cyQkCksBGRDigmjXPYMG8EjYfSERBdyMeszITA
d3v7KrG1sYQE8/QJG71V8ukapSKm21b5xrsk1834Qv6rGVWTnavbr3cUisMBp4zM
t9d4ESEEpj98hEOBgeoxMJ9P83wR36YNS4yJl2FVvddYLFJektStfrhhWEgvw1uU
rPU1sxcs8YKV3GZPjjMDtl+TNLqmlsq7M10OggxWu1t8yuwfJcq378yg7iLiTbhb
cnP0plhN02xAZN1SN/nNGSdUFU52bAQeyyeDqx5nkiVUsGx3KBS8Sex2P14MJNm6
zdll3jAH2DfxeMR0HG2CXLYgYlk416OtSFpuexlvDTU7imHm0UIeclq+mAlFNJyy
RXw0mJH9BoH7Fcjq5ye7k/pDsSs7bq8Zkvhjzy7dCAIt8DncFCIYn5+EEySwjmWu
9hCn9tF7jvpsBiYilDuTBGLIbLGTtNYwskKQgm8F5tXeTIBXrWWw3eiy2YibOsUF
UwULSCDFGrg0pvdYZpJOmGnS5HU0fMPpWsn9tKwNb0GLGgcgbRi66KjzuNCVVH/a
jXaKypmP/qFtviUeewg84isrKzHez/zgXO1nTCw4GHxJwnTB9vpgd2eWaAkZ5xUm
qWFMzIhKjARI6hHhbG4/UsGN0/ICNVRXYJ8s8hmRBt3pUIIP8U6LtzMABjoPOqSL
Gx6gOpNa330sN30XVgC25lGlNPi5RozX5Z/zHASA9+FI6nWQ5jBG6Qm40268a+LM
4nYYJGWfRdpcvzrnnGtLoXO3vvtpz8laiTIJMuw7E1jP4DPBB1mbLpll3cvxmhqk
sBybw0XGXTtCDm3BPT5jJkAADJGBkqH5aELnDgYLRIx4rG+lw+ur43PwwCAvAXUf
vrYvlHL9RIPYNSI+udZJaJbvRp2LpIsGXKGNVEsz5iGW9zqQ1tVTNOCEAGzQ1PJf
87iO3gkrltphblQtOe4fb/M0SVr/M4s2lW7CscYHM6VQT0ndN2H+KPw5h1RjSav4
NGnq5FV21DxWiYPafa8BhrTnySookvMAu/bx3U4UE7/Scw/1/t233Y8AcIpFcZhy
lx/1EpCBVH0WMIbxTqmT8VinXn7S5Yau6rsyaciiq2mXYxBhs9XCuJVKWpLdY8Wj
tAv3p6KYppAVKkTPNsBctsOSIzyp3ts5vpgkst/rvYkttRG1hsl/nOBzstITlBnz
YtVWjCOCtkXlUxT7vuSQMeVVfe8L812XAbBtBu4adOKKJH1u4/SWSIt7MFVqOCGi
R29t9zVuvkipf5aPcO2vnQV9VolQDHTOzqsH142++lF+y157KH9iAU2wsyZWRdBk
kqos6z8njtGEo2IvA4HHhJEv7eAAyyUqsiHGx81uLcIAqvOfEpgtycFu7oGPVlVl
AWaWKVe01M73ughceW965IwH53SJ2JNl2VuNNbKd/DtX8hNgf2dd3k22O2ZvsLfv
+DGQgREm/ktvDSwtqBNsHUdeBicnKu3CrWb1Z0SHLKHiq6OrpyWyc0eRmcgWTuPK
PF1MnzZpByH1tbKMHDOQVBDNi99z8wZyZJ4x6OqVnhncxKLnzuIe5+MuZaYg+9qA
bWtJFIxId6wHv7t0C+yAZ5gssSAENKTPAfuZV1FZCMeOvwMysXj942Pe+tILI5+8
JVUqyJfslXkKIRaNXBlx9piOm0VXacKLewnSsFndbXffw3w+M+AmPSKTr5IEvvx3
1+9f3XXQbVVR8+pE+eZ2MjaItB2TwBIul2E8/vKZ2vg4ws+WaxNu59fpng8FmyAM
qkOsoOnXr57co2NciJHfb4SKJKkwqYySUTgjNbUtIzaDSmHirb89LxKvTEo2IiXH
xNVXpUjNUEi7dvpRY22TpwKGUCmUynWiNHzcBQmDZlrWZVeolsvxA/34xZXSkT2/
D4U/31zQQDhn5RwJuE4HERpBPko4SUB0Buzgryt2kqkTYJbfsC+4ctwE04PaX0Zj
tHozgi4LSy89tnB1H8/jCl4Wi5skKwduk8obZgsRc91ZNbk9cBrwcNn8kJIJRPqc
ZwsBEBtSmbel3J5Hyk8oSZwzkZLHaJEXdpYs4ffowWGRQGOFRblA2avsYPyUZepg
Ff3MJIa3oHnVUnLqT2qSRMV6NLtX3seX/WTy/RcoFcFKiixbxEOofFTTEzvuhzr+
pV5Len/DIBbRP5B9CPb7yytS68tiifXkUP5tLuW0fm3U7PnWp/mWilvFgMXUrjpv
JhQDQqTrkZoEtu59cG21Qaf795y1a21s444molipe2pBpL8cqKTXtFnR7f3hdbBP
o8AMFfA00XzkNAtsuYn9HN0jTt47uth09/Bxf0DrH1t4PmQyV75fkqHat/+j5Qt5
vrZmdFrl1RQP/UjTaL7p8FK8U/hjw/hbQI3xTgqwwoeHgNKEyxcl//JPcX6MXUD3
02jMBpIhgtDKllApXk4QVH+cYmiQBQlTO4UEHNo1sP++HsKnPFt77itfYOrMT33E
1AO+oDbDoR6/74XmmEso9ZKfYsf74Kq+3SUX604hyWVV+sAPccs21xLmcWA0yHQp
DOXFFZ3eoLBCr19HBvuUaGCHIH4LrKc4HiNcLC3xkpjhobye2751u0lytVFld7yZ
7jO6UlFhi9YTqprZkJJQNzmMBQA1mdadZXZ/A+HiEKitypsX7L4XjXXd9Ofx3NyH
2v7+lcTUyktDxf3Yedge2Qr+NV6AEF7L5IzkIoC5W+YPKMKJUxDkTRqkwxC3WRzz
9hrhZgTVMvYgIfrHvY0N3GuzEg5Evy8967GW9KC0APGt20Rd6OxalseCmdMS9vd1
9m/KdlvIZ8i4o2sxNsFrO0kEgq9akUO7W/KSEhYXPTB6clGO8MzyRElq1X+eAtnV
9BxoM96b6QthDA7E3F7F1X++G3s3fjUvmaSpmD6Yqp06k5O6CPFaTQRYveRT2/Gm
vOPsdX52Y1ijgytm+rBdvYrhRgykVojIk68KVO+RQV5QduDccCvFWAaSvnt4xyQm
MhSomNv+T8bkZ4EcgC9uW+OS5bmb2uo4PVY0ZBblboCMDoyuCrxbJkiO7W8y2xXd
EP94SZZtrkp849ShwrU682N+8jyIZ+7xk91aDUUgry2S++2cER/8/wT34HI7PEa5
y9rj17tCwoMEX3b8Gy23YOFoJ4PHqw0Dn0E9B0YxQmehBHBU61Vv2TCsemYIJg7A
HDCukG+QLTmT0q92ifyCr/6RcLEzMBk7iGiE2X4gKp3CVYp3/ecJaxlp6G5nlKYW
Br2Bdp6ct8JxVx5PJPNqyKNC3VRtk1hejCWxPzk7AsYErvRsdD7gvSU6XVqANb2R
e0ZbYrOS/239GUvu7Gg8Y9HhXP+l7gUX3DLbKpDQPloTrTL91QQ2gu+L6/YteOJM
Vxfpz24W6xmxIvOwXJX52b+NrjqYcH0xcWtMSx2AYbGmTpKp7e+ptpWD6FHiMsd0
p6HQtRSpT7H83quhzXyMkfjS21jZj74LDwnpQonoKHOAn0faum/EXqeQv0MmWal1
AnaScGcJhbGfQvTPXgR2NUduqLFwvXZWWgmh3GMagShxtruUXysUi/n3dwqC6Pj/
HqAGqZHDbtzu22u6vN3yWfCT5GB2GQEvDFiVX4ZksVeCTgzw045y7gI2H24skRZx
7XOJNY1WarrBEkI4IlwoyKhV8tUdV476Vx/PGOMx11Vzvez525jJxteEjhA8jqc7
XLM7p/VmS8U8jlWoiZoevwWToc53hDGw+hSF8QCxizlkUrOf2E7TFfnskGTPCTER
ue2bR5aNVNO+ka6NpaO5ktJF6RhaTSrB8VAxZbjEXGLYsH/6jUdqYKXGuFDHQ5Pw
BAqd+Cc7OmvgsyHBSLGKlGjPY66FIA+8UDMqC1aY47WAcOb7U8YPJkEaiBfVWlPJ
YGj7HIl3ize8oi6uyEtNOki6nX6XW4bW41JfMy+KIYkhIU28aykP2iWqjmVo6k0G
dwW7+xy3fJpFc6jm5RbWJ1FhbUqqp6xwTLOmAEeW8jakE4vc8bjqmqIRqR4kqxKA
trwVZxddPfIopWvaCT45GQiI9WZ5gSLlHHOpT8ZR0oPyH+6E7bTEpFSfu3aCR8Hf
gWncQ6g6xl4OoTxCziCg+pnvz0DPOGo/eecE2KdGD0pitIz29boeTV5WBB24p1Ft
XyORMKUuHedyJp3RpfiIonST1/kwr+dL0gfcB2Q2f9fmGuMs+39L2A36NzHYoSV8
LDarOHmy7ziQvhRjO7rwchR9dVUUo1HRwCTRQjBkxesPWWZZ5ypPirj3XVMDUQ4n
7EHMjQp8zdEvH4WbkFexQVXAI7Sz+OlF856cUMa967sRMj1gMZKBbQLh/vVOq/BU
wHeiz5fglgyEPIEewdLsRCUyZCIafZAoZ/NtHJKP0RSJSWaORjdMmtjlMlFuXBTy
erBaHHC4hZWxCtOyTdW8f60XwqzS6BPXcF+F6fqPsk2YAUdyYmpCWZwCKG8sa0Ih
Iu8cfuMs5Iyws1gRDFiUs4tMVu5qF+PqNkDZADicgLkemKjd+O9ODGVbdbtYx6yj
TdHZZXrvWApD+hDbylP0cCUXJNBckp7XYRl6kfLRctN3vS02mBuSs8F1+Sn3awy3
kYm/O/OPKRoWx7fDsoljyq1EzBYM5Zg1yFJ8jaeBX/YhuklGyvZ8ZTHkultiNvIO
8HcNhaQbFm0ayZf4AiHLAl/DG9eKglfcx63K6GL84ARqleV9eis/enarjluxmB0h
ZHhHTy1NFnE6CSmDUCrpNG2/o8jBM/Z/w0RWuMGH77FGcOhD0EnkpPlH5VFrvI/I
T/vIfJQholULscQJ1gImlGOqblKr5aFQxbbJlhFdn2yd4UXuJ0x3ovmh4R2kDU/+
KlbKSgtiCkIE6sCY+ZNMfiyzhFu/xO5a/k/ErRMyDlrJlmAMLroM/EdrfGLfjOzD
DC19DLRfV/TVIUVINLySd039eUJazgQ5XYQ21sNoqgQsYR2EA2FQ8ekYsfZdC1rA
yso6cvxcUjd6SALp+igaltxzFcxyyrdymD7tlPsVYTc2y0xVY+4Rh20evY/1mJ8q
rR9VGY58/LC9clRV33ZRXtgF40HTZirZGVOhjhVampz7lNVybmGaYL+Qy/sM1swc
sOtjoaT22y6n4wCADezF8DU7TiOOEoxJ1EpZmCm2sUCvaAetOZ7LBeXT6uEldNnX
muIRfMKj0eWxURCDjcqFlgTyQ6S/fnJVImN/ZFIF2WxmWfDLxfq3Zdd4R5I3T9bp
cFLfXtBSSTqfZQGXBhopwyNNklg4kxWgKOoSDMtAaHm0pQiYY8w3Acy98pRIPVCn
2OvBR05jmLsNHp5DZr6Isq1Dx+HMfn9qpQfwYyhb3Vq9xt1jziDriccs+10j8MJc
mqgEVVclz6FX3E6OTZofeOdbVQQBs7SrEDzaDSuZuVzF/zpzG1qBykKnBbmAyEhD
bSCNO3vQyMEMs//iPSwy8zt9Qo3aNIecvdLIMsxM7TbavqGJld75WPAHseFWakjC
3XwSn/4MCYgF9qM0ETI4JwWxoArD9WC9/n9NqMB56x1hPxNPFSk8ESUDy5TlV1+R
F0rJrF6NVIc4uf8evYLY5K9DI6z00ih6nNMAEw0XGYR7fDC1wO3fiseHrTmGIyJV
9ZWIAbdPXL4WAOYx+XvrKWtAJr4/8y2m8qbNfGxlK47adw4cUKqgCnxBAC6K9wHZ
1bep0k81GUTeg5v948apeGK+2CmXPL1Hu6UpWGoDzfAHeovL+j8C7VNWLWd0yG/8
vykGF2gzyEjMgTZMeZCKuCVC2dSuwmmTdG7IeO0YvySqi9O9rJ3kZCbbFDNJ7hvU
FeTPH7AjXhzbcmlNrgJVI195HJOaUUhQDuILs3lRn/914Xvxlb7+HL+suAQOU+WS
MHUiWeq1W/qao4mwmJOAWNiemwYTRdQNS8pPaWp5K5cGc9FZQlBhU1X0MAIPDpY0
UPPp8yqsm9guB1jflIo8umi2xIoa8QdRFklYDEnQ3FfqscTnwAPjz1j4qod7vvL3
5/P3yx0RrTHGaegL9d1zIbV38Q/old8Du3BaO+DlHOmyOCSeXchgraHA/R4EF6JF
h3wuCE/ueu+LEvLEXRGcDS5qypl/SR14odaBrzipPdxIpe303kpLuXRmxBsUm5DL
41w8j/o9rUR3mG7WfLM/++IyB1TKgcjN3qEmOKScSGMceA2yyf7xBqnHYbzulzgr
DWRvHYws+btMEtmq2N+fsGxgyASmrHlOu98gmFG1uqmSB31fruzbsFkBEazrSzd/
WzSUgXguOtcbhyMlOq4DmQWJ5Cj81DNihlNAYA05Pw05sozmyU5MSr5EpKaL89/Z
Qtc8ZrNHfcBznwZDmk0mX7w/11enK7u3xPx1Sg02h7FN3TeO8MLJRAkp2Hy0+7DS
QFIpK3XLxk0PG7VzNC8FM2gFtLc7YHIdzQBPJn3fRBVW+q/SoT9etMkk4CyLd1/8
wvYA1mTsNHdO+y4i9kfjJvzjaOefT9+nzmxYRlK4GziEXozd8IO15NhClsBjE7ow
8NRJRRvDP17dCbmFkR3TO+kZWa3dYoLj92NznLG6Nsuj01h4vKGlNvHX7h6imjTg
F25/6Ds8uP6TmrJ8z+bsxZK9IObKIJ1l9qSmfBQFpxxv79efq6J50iCUv+4qjkcf
m38cZsY4aadlBFNXo2f9EOfP8VJy498COQ4eOs9VWLb8CB5LD3OS9NuavDKAQM3u
ulzldu9zhd83Z7LYvNxZD43cyvVT5n9U3gJ8TWIvqTz+vt72oYxCwSddZUClxR97
lFf9mF0Nr0T3lpritvcp2SrrXxoEyNT8qvBCWtJM6EUTAa7DA3BQZIJhudWV5Bt2
DTjf5B5CKSACopA4lW4m16fcKv5JoHA9IbKPa7jOS0QZ2gkTiOas1dNicFvTiN1q
QU+dtJPEzEbNpcjOt7aenkhzlBcgZLpBZI3OUNjnNbGGycd1hDhCtaKcCXuIGQAt
7DTdku5T6B5V5RG+FuAlMxwBqMIXrlNzfCJIZVluPjhCNf+RA7ijIX4Z6QhRhK+M
/g+sDUMoM73kY2q09ZwK23u234yUp7tS7ZeXpYiElYX18GRQzNykxz9TD+DCeNfR
PUTRASkDOBgqqZuenedoB5i8kBiz5UQLlPGobziUyrU5f74gy9DDNTT6+MelT03Z
9Ez0G3H6vg7UdJRMazjkoKc6ez9/ioV/TvpOsEO0gEZCzJgUKlZ3ipKpCWGaREKF
scZuJ70clC4/XtGWeY1cEyJs+Mx1Bl2iWe3CAhIg4q1z/HaXL32rnjCc9FNRIdMB
rGDVn/8kG3qzHPXAzRwRzdXAywETo6GMuT1MB8v0CuBffgImOz8L2yPAziOF7Rxc
x2zkolGXzDzXDZPOGJM7a2j/CK0rhm0McDVpoIPt3nvJ8xX3mNscn/LObmksYe5C
1o8XnUn2/8QJnzDqq+mZsyL3xB6wAKozRdGHUQNMkAg+7ejtxUvrJctPCoUI87X7
xppj8BBo8hA5r7GEQcf6GIp76J8UFtcNI/XvBY102vC2MbmrlbbM56Hz7uz0Wrsa
tokBVCZVZeTLEQgMo+G9cxR1IJQvQIFJtfur2vYxWPzwDsDY6oI71Kg43Dwuc9bS
WaTR+Z5uEkkdwO7KEnL75E75JFr3fS1u6YyVZOqZ1a4dFEjyauK8SocYJNOELq15
5OnxMyll4Ws9/412lo1blJUi/2IOyxS2rGtZT2pBRNJJ8SU1mZlwxq5j3I1vBxto
SAUpwcvEWnI1h/D2EPIybc0deGoKW/wYkMwxjF2UEZ9Yy9qAOKmjrnSBQZY7Dg8W
Pvcw3rUeIMHiAslPpLGoqaaUL+7vD8jgA9DMkvs/uVRDdq+KjfrgMVwiNrQc9ASK
PlINgXlU+1DcCYTrpvHZ9YeKUuHJoqG/1Wy6dtZ3Hl67UryDb4P3znBfwQ9NYHCV
q5lPA8cd+KATJNGbAywRR0sZrVk79ZVbP5bkqe9y+cZWDRa2zI/WAqzGuDGOcjY4
5FW3GHiC4LuTP2d1Ge7quy5K4QlnEzzi0xrZt4JdN6K4Mlf6+GYRO+M/zv4cE1rK
cSw1jtTOVkXGdKPXp5135Mb3rpUq/YPM9uk0N4FWgfow8hnd5su0QwzUssyFhpeT
RXoj9Dw5vF7+Mv/uHCGa5T4tLHB7+lFoyUxZaFGbJK1YVG7vNCFZkiKqowobl4ez
ynCZEfcsFQsaaBww1O0CWTMq+bP9iYaUSsW7lXtytF5CsXpxSgyqSrUPSRmqWBhy
YGyTTLDgdlAgxZRTfEMqxyuyDhhO3dP7+io4BWNMnnRYSnvbSvfTVxIDQn0+9abO
beH7a/sw5rZ8riuKMeYqAyZ7C7HPxdb0V+NyzgWx0NCPxu7pDMeGI0dvVGapDMdM
2fpqyxp8fR9eJ4GZZDRciYRhT6zkUKulc58eQntqakKxbHpM8dbCc/4E50gZPiO2
eHUrJpYTBoahLHNsb1iqvdvrKXUzXzIq4vIE9CVHKXSr8dLiORkHpPrWHhMYHOic
9euNww5dUcSV9C0RRty6hAmBKK1goqCERagTLfRILTNtywmiMpHUT02TlrEwHpZL
kIAE/vjDj//JzEPazCxHM3U8ydww79nzYf0FuQscABNwCjzaHr4+niFGVO9BCEYv
W8z1vgglpnKsUh9uobk6KCgQkv6vD7tY8ELiJqs7GfHuFtuYhB73LV6ldL9stLAr
TGlWWRnF9bgCnDLkCroxDZNWqag1XpB8M7z8JvVICrk3j7c6Uzd+/bQWJzYwmICd
RET+3fHxCJ7mT6lt296I84YNXkEjLdsayV3Kn+KUOq23wORFqTxT9bkc7WIp2aoR
J4PqjUylp3IeRCG0XPsjl+ZpLSJwlCIrTn4eIQXJNGw39f5oAceQiAL1pVGN9j25
FK6sO3ywJjVLlr8T1gXahHpHMhb9xXsI5D5gk9y+Wd946JDd2d/Sw1QCvAVEkY73
3Sr3CghikBNDESWuUlj3qNfLX+OVV+14fYjV7zuCIX8xBghikfOHlP6J8S2177VA
7CrxdF99LDBEyaef4oZR4m9+xRpqKUwZG1bBhBzOGFkRRXQD+FH+TODyfMOe2SIW
N0m9PGwjjcdsheUU+U/Kx9cJw1tZzOaTHxSQGjjOXZmcsMps+MBYsvTg50iCpLY5
yAuM2iRz4xXHb+OxrqOGYctdrK5JU9OQ9Kdx1IhHZuVQ0Wa1Fk2GcIFwerZdzTVx
q2ukACwcwc1pXymchsw1XsWy+dEmoZG2T6d08YkXbtp/7b6kO9J2fDsYOrKoZ+oE
MmulmDQXcFcCmz/DTrjtzNs6ASSIhFw0y8XoW2OE6GzibUr7EVFkx62R5Xr+7bsw
sM4wZVU1dRvkz0asOs+4vtGCBln5T4e5WnpEfdCz2qAk3W1aieSs5TuoHOW4sA/U
ceYSOH7ROHKwKPlzNW7Z3ta0ZWCSFde9XZpKwqhsXNX6Fw2IURay0mhzZAtk9yUK
/TlwyH46OuZLFEzTFjT9AyfGpy2f0c4n3POKtF8clRRI+ToFFYlyr8SKKYhUaJVL
GZ0aIfUPZkixiJH5joCLtrh6S5UX0NfyVqq+Kzz7+x0pJ9ulaKwqf2721LSwDLhF
3j+qe1qESWEuqPPYjHNEXVi3gGA8U4i2thCHgPl32vaaOHAq2oHs6x+Ae2cfS2wD
27VmoulnhA7ablXy7kuSdhebaKT/3NN0Bjl1/0ppYsa2msGXbF+OnoKHUfjWluJ7
YyuVEASQE8aeJzojeAslIfYrzpEqQgZWWi+WRbHnKT2/miGam3CGfK8GwKMouATf
jDI6KDAZpTxIuyUUT7oPydcHhYefLAM8ulAwRwY1uQDDJOwwf5X+6Kwx3VbZLbLJ
BZ1voVwlXSuh6L0MPswULOxuS5fQQpfpf/I1UugED/8SWTy+1sNOL+/GZJvFFRmZ
oAtvPJ1X6UN0EGGVzVgSIJ3C6tyorYLle9Z3Yl7OGg0EUuE8tSk6ajO6SFvndt/A
0zI3wFjOseeMoY05pL+MGInPSdRXIgz5TkjQBhfgvjGsLLHskysMrBBE/peIol2D
yTWhQpvpZ+icQ7vsB7L0R8ohWixV1K/z3ZGOXK2MOJZ/h1nviMbCCjTYe5ivR9Ds
YGIJNfR5SVRmtny7T67pSbk1Twqwg+YSVB9N6QfGjve43Lc2mDyXaY2lqS4VbYEG
LkZvABHDKKHMaKHyEkGvTmfeS+V+xW/K73MggtTcbGaOzOzwja7TFcoU/snyb/tt
qp2qFWHdALm8IXgGSIT8q6NDM82Ubg3d1jmHz9yc0oPgvEt6dFTg4hrUZDW0J//I
dOcJGFRLTtoiHg8xGgM0W5WQvU+D+tOIv2xcqAZt34aIKnftZMe5nOGkwq64pMIr
YN7iVLpRmyZbp5awVR7FTYTB+FmECmIqT3Mtahr9pLhVCl7zT5yr11nPD1E44KG+
k8Hys/4NygDIikC1y9F4qYH6FKZc0YmLT3NucJRCk28L9vGPT/1mzsNG1imCVKRf
WvOQjqq6wu9bX4tS+SUsIffOMvgZ2ArtpJgkOfMYbGx4dR7HIU7+bbBlTE+weyyq
k+0QXlNPbhndbK49Xb2V+SMJZeaaQxvIrxzXNVJqu7aPMJGdORkZkJBzbe46ZbvM
Wn6hcZvCV0n94CQP7V2hatPyEFd9lAa5n4hWdLdtFfDFUEZXb/C24cEp3TgV5o5/
cs50Pi/7+cx7E0an3ARpN0wC+DNfphUX2smnGjGbUkuB3MSnVOFTmMFDqsqNFwXA
TOfwuSCskQClajwuUkLGoDLtrBCt78msZq5HPHRPZxUDoHqMD1pPiPIqIxoRuiYB
OOawGMa1g/CgbsUGRX23t4gaBAOPlYkeHT6xl3btnXoPJq9M/iexB3Eh82rFcYI2
4FS/hKWZ93fe9+Xc/mNpZdhVarx2OYNisr7d1cd2QZ28LEYO2yNGkJGtlzykrxoy
X/Qa2JcJQ6KUcoINGjBX8JJXrx/C60rmcd23beRco4MngCKtKGtU4PdxrfPg2UuQ
Dfuu5aLP22BJ5k+enAhoU3CeFXDhzPoboRLbbwty7B2QyyLeznIPcQNKOncrf6QK
+EbauoJCcmcHfumm7qMr9FYit3xlOuT6T4U4U6maHBfXFRlPfVBme6kBH7eT5rCM
3KILvUB9XKHw+HvzQ4VUxgGf0Wej8xt34W1B+52qdJ9ViBygEeFjYiW5gB1wsj7W
m5O2rxCv6JxPhLUVK3gjQNKUX6v9J6m0cMgZXCgl1YGLJiX92Y0BtRJvk6nnn4WN
nYgagdFgWdwGGV1uJW9igRwFruqdZL3ofs4mOjYjLEGNsq9WP1VUPfIf45928n9V
YJe2OZwdPilymRh2MxPVa+T+xNCIFe0W4d1h9XI2Cou43vgmR3ifcIMSbkD4TulG
ZdB+44rhXefX06RsXexeYXRLcQ1XRIpRNCOGSjpxHU3wOMZhyJbA7fzbDNiV8rI0
76PEcfgxsybfQXBgC3wtAOsQbyhPVL038xr/GqGaGmiveBouEQeZexnRWeBSc+gO
CsJlpSC/TSpjf8rWqLvZbFXeEmzULHuko6WGiaKlK2IEaVWwmTkcx7yhUGjiAhHZ
/Qbtw7fCpgcA6DjIObWqPtpVkwmC8d0mRk6jKS5/782M1t/lmLCxN+nKBLie3moZ
kRcw3JHdQHb4NaC+Fl/G3ldkSA6tBGS97T7LLhIybZg7HSPNw/+5T4s15JwNAoNh
AcQsV3i19pnR3qsisiVSxODHBKWEmQx0xdZPdsn/xveELmrUlSDi5scZC0UC4qJW
5bxs8ant4eeMp8dUQCxZvsK3bfv4MgrkN9E34T1aPC1JBx+EOr6Vm9PmozxYdW0m
AEL3ZbkC+omn6wWBC5yBh/cIG5ODKO8lwxlUy9fO/zkq2IH38Ag6msf6kXe7GWWD
tQKSEPvCRXFGZC01KW81fWI4ElOotpE7fGPXzwyMsfByTriq8vgQy0wXdhb7uhbI
RKDqjCgig8XLDazTPN/WdltjK3hrPnn7nBXSE8Rpi1uoe5wiy276O6D0D/iA5K0S
tBSY49eT7ZTmjxuio+Z6DsGfC7RPNRAjPLQGucIt+hkaeSiLWfW2sT5PqYHGGtMR
IuaVwYmhGwrCSrIppHFoVlC9avW06fV/hhDty45CTtN0mEh/J+IOoY31pzdLGW/h
l0Rx/90m0TZH8xBNYys4gjc/XD/RWiFu9LPH9UINVT60YWfPtDPlS+Fb0EbCrngf
P2q99turH9/Md5T69kQqRbH5nQwnTqk4BiChyH6p0Ieeshl/6GcegYDqyMwXBak6
a2tZjiuxkcqqY04I5jmkoUyDjnOBR5svVPLZOvWM5eoiw9Is+O2LA8x2egbGHoAs
quyY1+/tFlVGTQDj9MKSfFMlB0EfGG8YAc1ODn6anSI+YSanaFafge0SRqAsFk4I
f8wUbcdo47n/fvEiIqinC6vWo6o3noY45HEjQB78nSmT+5fRnP28z32xJ2wNdywu
VS+tAnxtGYEtJ126HsZv5W2WAZrgoACxrrL1Y/oXoFzzT/LNWDjOjMvUMtam3U4n
ijmQ8nSNalx889LNbUFK+nv8bDGiPjV+jyHJwuxbX2gtGUv0mwCkb5pQH7IJ/tQk
Xxu2Iv+BlAWRld9K6IaS6WtLdDfwicaR0pvCgNE0yA8EBskCG4lZr905DUO45dTb
UfZSvudAEz1+OEu849HlHE+V0i6XolcF9HN7LI4NoZM/s2xFmtJhljiN1QMIrpkp
HwCzHy+P/A0NhFU2WDIny2pq9/w8VAFr5dEnD4bZJ0iiiHIisbwbYI0ciicq5HYe
bB9/3qeJHaGGUeaFO9KZOQ+bpTbwd51iQz2hcp5HfzduSieP4Tdj6xTLlgIvikLp
cT93WB+IHI788uXmqQYjUZzf+WOq8/YnZuoJMynRfneMR0Gph2jjp0JBnAajLq28
WoDHDv0lmLenEJ5JVcqVl/opTTYOAekOYuop+B7xpGGCmJISe8x3dzuGw5uag2Lx
xr0xW4G6ECurMBLo6mYPeCnKLcKv7k6+ofYswJdE63II1p401e4JtyW6f5W+cXj3
dWBuo0yuxTzPTf4g7FqRnqfiiQCXJ/NRnDqm1Mff6wZ3Q/gOON7pIb8DJOMOkrMl
UZ1upJrO+6l3ZMImPXwD8cqppP6EfnajmeMJ2LolkAakBpqMQuEMTi6EqbaFyEWe
qmxTc/vUsrjumDecVOAwmg5h62and1KjmlkQtyR76ka2G7e/TTGIfTNcrmxFi2f5
NxhtCIqtN6SVme48b68jxgFkLQc3h1N0KLjEiG4K6Qks+92nM+H3T96R83/JmO9+
WBv0R++1MoCTOMWUHcqVr5L3EmMthGENbCrmog7D1O7wdc0W/S1haPpU7eodmxOc
i+/MdEntnjlMr2UDT6ADmxw43+gVBCzdnVTU68uNQ3rflKqWz7IOON71eKeUk8oO
UCHnnJKx4QKzboSM77oXgmxJCNF/omHsgSjBJHt0bcGdW85gwW1p6xCZA0edk6SO
0EssshDH6jNV6ubP/O0hYYlqxKA4uWE2NG+TzR8bpKA36FJrF2m/iqmB+187uMoB
BdU2037jkn4ajSOVDphKWjusxg1j3FKk9jkiGRHXC4v/xR9jVngzUZyRdGrtW9vI
l7oPfis/Uk1VmnZP2CyCveCwPhj6/Ln8HX3355kJxtmaq7kEScmVpJzBmbGztxvJ
sFdI8eNgLPL1avLN9P3jGSBPCcAS/6x4ITAYdfz/2NOD3zxMdcCBINqxiAAQ1Buu
CmM0oe/hmHcJByp6RDGPsiM9V1ZoLV3fQ0W4MyWm1xvjk5Ploc7uXm1Z5zOTERSA
mOeqidls6PI+8qyr6dWh3qrYLzHrFXqbq/NdoiLQ6QcxRTUATHh6Za9/5zJR3t3j
5CzN1P3CiLYW191jNvkGRU6RllavZcOfpwi10Tuay40onRsSDNz6sxwazKUJ8Obz
dJwtTh57TjTTaMp0T1TdhRZ4IJW7E5WamWVp8t+qeP+EJKq0XbpyV+vhozFKPRyf
y2L45Qbm1RT49rB4FVGyEyWv4WaUzi2mytJAFs1+mFWt3cZaeRKDTW6TUuyiu8+2
V2ANylKTbe6WQWhb7SkzKCagne9YaOydqXHC/qsBzJJVa6wx1wO0IhTm4b8fw0YQ
wfPDwO8mn/EsfMq2KK13QiGZ1Uu+XMs5gySi2c4JYbWWVB3ElRQkaGUvjuqlu5rm
GuCOEOMPAYnEEty3aF8k4nXjXP07vRC8DpaiIh7/vibzptui5KlT1ov68a/5rQmW
dZww87yIX146FnrQ76aoJIstJWvmauIQs6IhJHzLm62FLe1kIQIeMvBPj3r4SE6s
rFq4cZyQQKJVIx8zzmAK6HNjyuaytNZW2Db31hAOy/ct4Ao8WwpC5d8WRowCtXMR
nSeMU8J1h4jp0esQ+7i7Wq28TUdig92663x/U5Xec5d3hqw9444k6ZospoOOKn0z
Jwq/BUCKFhg3Ng8dBZM1kTqBNB+X8Cpo7urRVCIqA4xn6UsMxXCSxsAtIb4GpGH+
huBIkh1IdjEePKjAPJ4FhGYLHB+6GRIYGW+srrP8uI1ndqK5nDO7cqxYPVwn1E1h
HEYPzuFfihCek/5zXzAV0QXYHiNtECg3VvDbToyoJl/qtBeeEYKglMDgcfSzzlCR
4HtBJi6rddTO2pl+Qc6t0bAPHz5y/mCZHYjN8tnIWmg+6LgxmJ81aScMBrMfYcH6
LUelR9SIs6i9IodESCr0ow+3ZnyXbrY7OK2DpzMhiJkZvhtpoVsISD8m00cCJu0a
HvujATRRXDB5c1iEwP1wPq4R4hB7WA7M3L4eX7h1VR3l7xZp37JMePl2A0vA3qsB
5eUwveUt1imqv8dapHN0sNEhqwzh87NOrB8eGge4wySncX0LL5iV1urvwsWKXazr
mLg3mmxKPoIXADEGFxT8KB5jzSVmxFMsIILleTCklkE8v05Y15YlPAX6wNCFAiJK
F70K2Pn/nq+dQRXO80g1/gB5PO3nXt1bQRqeJtCloXAsBj2N+Blvs5C0sOPyc8vT
AUL7bQiK+vd7Io6m9Mqe/lT1USH2cff/YgCzo4cQYMdfYdvzM0CILQFPZ6AvEWIo
WIhwFuZ6rNKEu9l1VUC0B3/kEn3FW3qSyI17ipJPSfmte1E0RpYd/1/inCzE5A3u
oWiI9Rfd3C0z1kwKrEXP3j9qq2ZbUZSqnDqkjhUGm/yjnuVkHRM7oICemg4Om7LR
Z1PjVYjrtbvZS86NKn71X9TiX3bADjs/jWHgOQm6gdAC3/bJpljZpf66ydqgm9D1
ydzZT0AD5XYtoZySaoosItK9OlMY+G9XG9mGnMTOwO4O7lUrY70mDstl859fKsOz
sesfgBh3nDbwwShnpZ4RxVKHrY1Dvztm+89nBbuOsiFP3vYCX4kG60UAplEYDi4J
l0JADKlMT7RQX9sCZjL9IIbTzyf5+ePHaGN43vWbsqArUYH0og+U0QSjOPFBY/rK
Kh6UNsJntFSQSqsoTUUFG8OQOtIUOdMCAelvVKf3JK81L1gKMMhgmmbUG36ns/pO
0kBZ/AgrekbwZHwHsqfwCG11oIy3SSY9N9K5WcfTUF2p3UVlm8RPbe03vTnINwnR
JUt+0DFomwSYk/PBkuoj8MXTBuHFhYUs+rRPsqW1q7RW1EHsc52wBL/QymcnOK2h
kNXv6E6kFLEqXeRnZliKYyldx4lag0dieqQvzTJnsXQsjEu4swHi6HBMoDRx3trL
GrOGpvlIkA6kt0L+KbcYmaY77p5eMprLLHivICPTpf4wXLiMSnT+pjqQLdD2MMNh
jHJ42jCejBy7ieTxXJCYiG9CXunaamailObYFG9Af9jY48zsEMwQU15+3GaSF1r3
upIZARe9tAOw3Z6bu75xMFBqZU5ov0NqtAvIdS6cfHl2kEyPhaXlsmBJGPgsd0S/
k5tmrsPzqJAwkQj/xjBaqnoSxciDJmhk9vJNxjXVGeM+NMdRk8Osri9qouOyACFT
brEUPTp0xhsLzRoH3BQ//WPdH8iAvoW3HgdG3FqQAL5EY5mrHDDWT1aQEyjMfJdy
hwN6Joj/hwJloz8H0qbI6xmYOlFVCXbqXup59DRST9KRtUMiJnQXOFrA4JLQbWYf
wwsoOat+9e6Iyp4yilkPQsE63p/D5fQANTKsXTIiIMrd52poyPo1ib0jRd4PBIWV
D+O8H9mISYy/IwZc770OnnayyOxm1gS5LLMP6nJ3Z+36j9jRSdJk8Tprh6TjVxy2
YAONRN4Qv+lxH2UdzGrHpZFUCHYUNa+QKUqJvahsM43ApDTYV+E3CbUWUlaTDeZn
A6aNTPgRq0Owih4+IMBIUugCBaZozsfUwunKZf0dgrQyNjjfYynu8/ce/AMGi9Fg
QjNPB1IjP3JDK4Dmx8dYoNlY9w8gqUVEfJ0gd2WdePaMyDtw0wZ+T16wEbuN5moT
EYLUBvZxJHnsTl+BqD5ToeSf5tTUCHhyO2v0CW1ec8sQNf/of7PhG0oSZu5yPTHf
VgxayF+cDgdqGVqSoXEeY2dMQBVH9wmIsEYnHVi22nTdaUnEDhjAzm2R+ClzoQg8
6Dbp0vx0/6vXXd9Vru1RhH5kATEHdEZvGjnELZKV9DViUSbkMq/dAvIRwXz1yKM0
d9AiTEHpXTEEtj4WIEhs/8YC6l+mqTDHQf+CXdwo4j32mun7ePwOoa5ArOUIfBBU
b0oH+wosNydp9ECxodyjktQ75bU9c+XTnkk4Giu02uhjQgyENhljem3JwIjWgzn4
COcHVlMTkAU0+q6WQIR39iBjC/Njr75R0BspRKuGIw9ExFRF/Tp/AtqvO9CoDLMQ
N1qPJ0aQqvKRNohfZgnpIchhTy11bEV7rrHLD8zhUV8PuXhHGhYQCwNBVOQc52Yv
iwQSqahoC0o2jF81WCbmMUsd0zYrQhESSTS4qEU6b3BmJvoG/mlOTn2fL7wDZxvS
NEiaohCcHIMQmbiJOYCnCCzkZqsMZvJm5KN6JzJoEI4wq5BuxQR4+VLh3bZvo6uc
qcBqZXbZpp1qdkIk0ATFqabw+w8sMyQMGnJwaN1xFobeaZfnQcQtRSVrawmaXe7s
d/9uiqC38WObWVHf11TTrlOYcwL2eGWSwrjnTFjg7X8/sraLpdpNZddfuugstO7M
RDC3XFVGX5ncCeKTmtcV9shVbxD2qfEsJPgY43m0oZmGhKY6iKQHIDa+nvu2UtZU
cjVRGCideNk2MDRuLwpjo7vBoQWn9bXS+oQOj27O9KAVId5MvC1Kjt8xE6OctLhL
UrKUH7RK98a7VC7hHS/MDuLk5azP1un/VPllszKEKjdeBeVl9k3GP9Y/jeEIqIgy
UsDlPrivjD3EDQaFt8i/2/kHVYIvSFyQYbpbjFg50/pDcUbM20fPxQKu6TDqKZ7+
HlUnU887usezed1gguGGLezi3UEhReDPgnUQRvGTYvbBxy9MLZl97vklsoXLQZmZ
S/uk+9gWcXKlvy7DMOK9GEyji08XvDcNk61DzEFIoQJ2pKQYGKx+g9NWP+yb5g5g
cMemNSlESzFMIPIIoO31HPZYikMTLnkC6nkPY3s+Pgx0lKuh3I0QUY2qH5vwQTc8
o80Knzr/d/P7hMpgJR8RthLPZ7MWLBZNI34l1nWxWLSOFGmtITPa/+HB/z5q8cKC
vgKlO00HdaZIPPLfjvXQzSodo8j+y8R0JiOJJ3AdN+gTnvH06dhuKIHPQzXa+v8z
jHSC/WTFa6kz/ifiikacFrNnPfNDuHtDek7fPoV+6XQJFtxw82P2AwziMlQ/bdcw
V3e60v3X/rcmfr9ZpobFN0usvCtb6JJ9uqaNB+fcfk1v3D85JdsxqrypZqczG87O
0k4slJQ+lRmzXEsh5pxKklP7s0HwYVpGx2dS2MmWEsvNZ/xBlEVArewsA+VTIX5A
ESSm8l097iF3OkojbARWxhjWsRQynLIROsgCufE3nzUA06OSPjQ6t1I0wHLagCH8
EIGbT0oAJ33Z/ZpQQKPr2W/cl7XoTkcXQLaNW3Bvr2KqeLk6iKdhFeGEYTM79YjR
htyUyJRaomZyfpFgNu1tqPdFxfdU1xFFzP3TrwyagDcpIp2RC+PfcdZJYYKY5vCk
4KCPzjh6G6PxlZk52hT/hIJRe+HJxZjbeZSiPEMpQzemcErKD+J9yDsunDGqwDGk
Y0qT0GJKRJz6/CnG2rJaWtTtxfhM4WIMVy/xTc5uvZmWDFKjiC1KSUS9k+YOm4OX
T2KVev+0pFfwkmED4DMGinFBRwgAFbEzAvui9Bv7wtnTem6v1dteRvOQfRjn0dIA
0e0HxIZjE+qCy3ZjmujC2d6e86/tj/i+1l1U7sWPNFFAFVo5993aECBecbdi26Pf
Tr6P6GP3VlRRORPdctdvzoO7ScgrOd5+xy6GltR+ttUjP8ZkqlrxWJxpodc2GiDj
hhnVW5+0N/oaxmVffHKYmuddfMYqgAo6ueE2xTicjGO9kDyDA3YoO1mVdkworQ8r
tvaJMalYHWW5YiCy0BivR0kmPkm+Gh5ggQ2x2oIUQmL166oHqYcc7Mswt8H5iayN
owDrXANOM7IGPJ1b8igDJ75KOwHOD3qbkw8X7B1NsGD6/BHOzpVHMPlrVPpZ3TS3
etFA+gmi9MQnGjxQlKqX5V+y1kBIj7szK/ymeElGdZmmNbwHMP+2eMHmKODQ4N+s
dLrOIMhkWWiLJPVmnKkdWSeRp5p7esRhUHEEhcJuwiC6TyY0Xl+KhDhnxzMwgHNO
U4sFGTqeXWbZdKzD8LWtWVFWcrnwXPvU2DvafSH074oRtb34gkvwlc95KiFyjS/E
5d7gjIEuB5CNVvwXoFd8EtwaP3erNs26KVipwRW4tlaBoPJ3CaGN5LaIkE/uOe8v
gTP6nACFWJAGhc1r3qzqm3plZk+j5UgtTDQeBHXhcxN1Pd7evlN2z4lCZBrwCqBp
HRUVOHcuf7EODOAN7qIuagBTwBOCXVFH5NQ5+2N9Tg8Swpizxnnve0UA6MKTXhxA
Rtbx4mn/GrMgDEKcJ4GAmN9oi9TWMqo7FxJ60J9sjgVyhwASgA8/Y4ASfb9ZQyI8
/3UNCCMAhBXYc9AjmmGesWMN+MU/1hfBTcnjMMossIsFRTvKghurTX+yP9gRFG45
+N/L9lBgGGh1SFTEgq2qc9JHsvcDkpXsOl+2EOHxj8MUzoK28/vhFcqEaHy6wy2/
Ld3KYtuTvRth57HfDPGNT4ZZfcRSR8WjMam0w60exoZ36U0hzlDPflvTamnBhraR
Ux2mD4+3Oyoy8hYBvX+CJWD7PEoZOTrN/d8+l8wmx4AWMjdsRpPHOqztoFWQQhB3
E14x9YOi1ZlFh4/0RKsGfgKyddLu29Mm1HYS6st+6mp8jouAQFit1Dm/4YbTVvvs
L2tglWNuahV7Dl3kdbrY3MzdIu0tHfUwDkkEARN7kAtN101fN9V47JF+fwcjQfcB
8aXZNdrxiHEZchQ6goyTSlW56qvtZItsJVEim1A4WcB9YbCUKfdQ038UKZSrpRFJ
jSxzAQBR05VLPvS/3CJb//ln9R2p/HcgpoVp+2MU4UnBwCouujXNLEdx8PJj3FM2
VgIajhM6MpBDPS3okRJmX8UD7cNKreANLFsHFguQoHkOuKp4AVHBvbARe1qDzalj
1dZjltASCw8EzKlFmEJ1nC3Xu3xbcf/ahmmVk+nOOMxHqFeIxyaE7M3DfgnQLrdY
TV9iPpUKKfaubMxUioPmQ+4JAONbsvruhHDy8w7x5mnWXYClyr+jTV77Yxu7AtEW
XfB8QZ3MNE9de/s7Ek7ziayix1k+8Bjl52t8IDINtE646SGQpmR7x3WA60XhWxe6
ufFnkLZTZ5ONuR4nERiNeGla/sHWnmoJh+MQ7/kUgBQrZV2AFRR3FW23XJsqioSL
j5UOOlloSFZvkpKR7ln0cTuQK20fofH4cHY1XZmIJB68md2JWumPbaxJbEViFg7L
teurip29WS+0xoEDF59/Sdik6r3XbY1upk9JEpAIs3gFJkRMoOX43pqfz4EXJ7PG
LMrozlHkqqXsLMvfLalXKt3SZTFwufYNFdB1fkh7+mKJcpd0tSeMnWVS6wLN29Mw
gn0hEFOYrbbFruMn3s2XMCxiAcngghVY8eciYDfmSEgXY1QoFA2Z7ratDAPScbQY
FuLzoABEEIliEvXUx6xm9x+ZbyleaHhpYEJPVVbOFiiATreagyB6VK2cFZotpBTE
voZA8QjRmBNutXxH9uKiezpWk4apDCFH6cnhgC1R1ak2yE4e13HSndztw/wDyJ9E
EAjsteNr7u38jhTgd1hBX8tbu1HeSeYIkmRxTenv2/TgVrtdegysrtQ/VAfkTVF4
JFkF6HQxMtljKyKQooSr4uy9yHZOTcMG95IaNkAAmckLLg0OOUiWjSuZCQdZ9vbT
ms6DKukGdJZJkD6fE8Drh+0z2m2dq3cXfuxWqG6qUxkaOCNeXrH/7ZeZaQ1hyVQQ
X5TQ/JG7GkNhErb+yggxCmQO2OOa/VXHMek+LajItQt5a656x41nUPnsgzvvbOVb
kT3dM8nev/9DU26NfyJCxltTGF0PQ3fADO4pPRAyKzcKtTtWqEuu4sfYP95PXwND
q1qYmt+QlOYzTQcab+A1TtcNsnPu7EDrxz4Hz03CvjjWZlXQa0oP3HMcIhbA4nOP
oJkS2EMZwTnxe7EjEVEPZCBkd0ZDjnQhiGI9EFWkyDVSNYbgPjfdGdSxUZ3tSQFj
1wLIfXw3lIxs6hIk8mfzfZShpXcSH3g9dyMDsu2EJJo/eDI+Fun0VLafeKKguPCu
xLhQXQNrnDou+hm1HU9kAcYoiCKnUXI5OVPhnny5ryiMOZL43K5CONWD/+9WB8El
NhirOV3UH/3eS2NRiRCtMgZIlPgeeci6NBZXKeyr0dMNn95dxvlXcBZ3Io0JbBeb
GYkhA/fu7utaBTO4h/arVrf0fMnUVTfbb40QcZl4oEXTDqPptLmB20bifopi8qrr
pGb1ApZA6USFGIqM6PoBKCFavuixhlw2dSwV1Q1ZBUK9fWJYycw8S9j+s1ifDlYR
hQyGDhoCu2MXg1Sz/kUDKgCUYoJCR62mCeCbAHmt/0T3xq0eeNN/fn0PZ5MazuPj
KVYMlWcVKSapqLsDRX+5/12bQ2PVbJwTJKV+hA3ii/f40uPqQFf0f1r3Hgj0oLBg
8INCGF8C4ptqvVYRJEl51d73LfM/UsA/AekwBvNw9gzjt1sgvzqGxflBje5+qRgV
wk19tNSp6EKVZTbpaJox1Wa/S8/p/ooLbs/hza5TdWO+yVgZFcL4yZ8zRvsokoGE
sT5bFVryQgs5vCCUpCbtaepnNDum9Lj6iD6iW3uC+GYpX+yw6O/ad/GG0wMFBU8c
0wSQL0cO2ceh2sD3I9L6VZqeBQlicSRFjcZThyy3b5k8gsP6MHh/T+tm6HRAWvpP
bvEH3OrIPOzgwrIfwawLhNrjfnLknicNzyRd3NFEc0je4Y/qC7fxDkkLiQFiJt0N
rGk+BN1jWLK80ZEnDutDkl3Xq9Xdk3wfihBwbaW94UmO20BWxz2xFmxt573MD8aq
kygWNHupjx5WcvcR+nQpC7Ku08qTJDQXix17yblkdHh8zaEnIxhRTeY6TklwUXKL
zDnnUEGaC0vXrXc2C2waZRj5fz7d9kt7Y1NNsY14eKMiSeNeUW3SEr1yVX+58hbj
+DTdIJZQBobCwP3ihzRuiOugpG7DE6wA3dQEvzRgGbdvienLk8UiRmKDV2t2HKAP
ajm/S1CoERgg4XgA6Dye1N71rUVhRf3TcfXR53Sm7Mp5DTy0M2WU5jlyVdFJMTfx
/2yyQcQJz3chlDl0nCXrmwWHj/sKpkLzMjhVqKiF1RmTG/u/0VX5F+RSTPSuG0xo
y6nGi4Z5ysBCsH4686fq0kXitVDZbgA0eyHQKzY+sbTNxq8UM2h8JzcUabry/nJT
/va4DBWi1IxNkivWzEby1HjYvJsst79aWFaSyQ+MHrd4+pcd39x/GYn6jkbOTKPm
yCwmXGy8kpoj8idtGgLqQ5DE79QSdmlimodHCoBDCv8xvE79PfgMf5qcBxAjZBig
VJ4xcxIVEQ/ikLhzrhV4edoAxF7YaUPeo1mFonP276XfYEnnSEVMAKviuBa35aBJ
sPgpjgeTlbs6E+42tszVbeOuCGy7VjI6jyBS9RvxxVTKxkGg3Okes5ezSmldQPZA
gm+B2QU5aVmYq3jKDA4p6FW46wVS1jydEUja6NahXipTdkdzLtFZjzJwyPp6Z312
UJW+PI6uLe1/1a2eD+bP1nkxZJK2QWA+0jwruoelY6da1XP4nC808wQzDTJX52yI
2yUUSsKaF4sx+qF0fIBHGH2fcB/soOrG8fuZa5DD3HYOcJA0jUoYgynbgRLiKJ8j
oDu0QnfcXxBDRFE7T0F9Zj9NzMbRxL6kW9aabAdIkWR95Nd+dGIRbs3QNcHnztos
sa8B8LjeAkyJ/lqPPeF8jWy02Lf3zpjV8IRjPgtsu/0PRvyMUkOoFSRJsl11UtHR
cKYta2SX6Q4P0bKDwq4ARaXZ/WPv9+k23XMCqOB9JAzrOrq+1bvtqS/UK5UZWXvE
7QfmaiCzqfAFZy/+nbwwGCujPpezRBIjAozlzUgCabI5OELTO2oQh/0zAsMaBG5f
Fkg5jn9uGOQEhCJMecb+r2AwYayWF/JlCpTWi6k+5JzkjEeG1UatbpHi2Eu8TJ0p
CLVROb3z/UVzV+7hDv+UJkZP66cIXgq6WKBW/oK2XVCQd7RDaBpjoQFYDAB2Umqp
WnjGkaVH5eroQ/0JO3TH6d46p6zQQnTqLPEzOMju1Lyph6mD4MLfe2rgjnFVdn5R
6Tno2wD+Hf20bqD3/qcqDFPj8GU4dIYXk0+DR8vEBFszetu8Mx0vW0O0Q3OYCvOl
7FLpWREXAfEYotCVXhwUiR1n49tFil7KYoF6LXX8psvw2qjSPMLDm25V0Qe7BEbC
pMM3RIB//citZmn9gt5w19KiwxwGKi7EAClyO4EG3vkc5XRI9GdmoCirly0TWowq
+SUarXL5o7LyxztkQ5C6JrViUa62aMBRqvtkjdtHshUVPWPXVfUKLJ7ZU2abSNfH
jbw4doUvwZ51vTY79DZaHP7gmtgaTjPdPXhMeXA52i8vjML9caJPHDeBy5SbtUs2
DnR68yvL5Kt9rctGVsir8pORfaBdDriL3HuujuGoKVQA+sGmK4dEUjYmBZQHHvkc
KEzYt20S0BVNuA2e4acDwe46gZhjBRklJij2Lwe24UV052G9aS7dWUxJVDbjrmY4
tt/2zGYThw1WD6pd0eUa+2uYOp0Y/fayzj7TuCzK8ZVaCwF2nab79Lbt9NlSphAp
h5D6nQhdbB5ltCVbNQSb3sBgCPMDNVd59ISRLLMX12EWkM9pnAdeb5hRfKwYub2W
wf1XQZyMEuvJAnC/pZbGeGlyLSfdcx5dSwzGNPIpkzAuHC4qo1jCDaSU2FM3Jgx7
MDysc9HUElsUSerVZ8X99qyeJqukZQXZrP/jMddwYAyOhuXYXFnLwC1Prhmt/oC9
wZet144xrDSA7j4SsXCK0FqQ0F9HziDSfwGMv62JxwBTyKp5QWMKH8FBRQ9SfFag
WcxzdO/Kl5dljKFXzZa3k6PhsNuJaO4BUDSvhgdmdoIepjk5wJSDppqo17uHgw5g
NT472XaopQWxnqOsys2prAIiirvZ80TV3K6v8kDgvIf9RHrpKPaM9GkmOUlCRa8Q
/jpvXIWue5vkTlceMq9l2HETsEDpGQmbWMUvbfgemA3QN8i+tDIYGKyQ2vP3nNJO
UJHRzE53vIzUE20Yt/jtJ10IEr4J/IMBpQsRjdiC4fUdV72uKiwMX6C9Pyqtsod2
BFxGvUkBPmGiacmF/41+nFOo1rvh6ocjjMxP56Aq5/Jz+n/OVOzidQR/lOLgzANS
dpeUjB1jKFHsP13ftVXdthG6N2BiujVDH+P2/IITCQjFisHG9DdP7gFp1i/bOrci
+VlV6tF6Ocrg5AQntXQzrt0ETEYsE4iefoJjX24JVtjFAsdIAjoK9JvposqBkMjn
GwcewDuLtGpLcBeRm/hQIaEZ09FkCChZiDlPMlj9sXcaHy7fSOEfhyt70Y5bUjLj
Oign7eQ+bhDhyjwCCzA+HHxIner/1Ppbys/mv29OIOA6YpFKqXJlZQu3ROQWA5On
0PE0QWx31EZMHjJKUwqG/z7YLjymjEova2WirA4Fzq6hnQLZlEPFaCSGvTxHEXYC
7ZvxNUeRMWdn2FIagC0ntn7fK9r5ahD4VMg3FlvQtaj/39Fes+JfaLfDNgX8eqc4
IjRnhNek+VKDwwRenQi2UZhXLRh/YXuzZDO4rppzSC+iZrBiItYgIz5ZPf5TAeHN
8d2T/WUhUcWYrQHcBPO7axMphROc2bHTnxvX9dTsuFw/BtJekN40azEn87WQf9k3
yaQ1z6wjcgL+hC8sAZNXd7UWgWHHVdyHoSZ1B+KgP83Axp9hJuxEEh3q+i2G4Gyt
lm7khggKfwILHFz2SfLcYUezUBvur6rP+gYq0Wqv2LBoPPa2sMA5RKTtrvSDY9w2
bWIXQ5qxX6Ck1XkaXMhSm44j//JRMur5UtQua3qI7cz342pRpOr5Nvo+q1z2d6zE
kNljjKzDhiKSWCYH4udtVBj9MNk/kvlIXBWwAv7Jn4e3sz617v0X89lnbWYQPvOZ
ZyeN5hXzF3d9ePJwO1hC3FC7ifv+BnF7VjFKTXKxIYAAZalYy9bUwORAPT3Er9YU
CBuDj1/HQDULgoHiIMj0EwoAtlJuNz9hpDktjQ0UpV+vGUw8qAniHzHV9lGUCpm+
JJ1zRE6QgWLMTeFjZfuO3Twpl3NfLg7xaoGtUnfc8D2hyPHCEQSXxFVT4iZ/OlRT
LQRpYMCdPTbfBf1+QIl4G+CrxIRkGs9bq8+IX13r/EIxodE1ve+EZlXj7f0AYAqm
nzgC8XiTfQTJ8GSxEfaeEZ/5B006R67HPB8gvFxxBkIpqoj8qKDPdd885H95aJdU
akDFdy7ORaNp+bqEWbsCVycO5IKsSD55TKj7AxpOrFPwZCXV9jBd6MN9cQ3QG/ZD
8OSijTCcdxWNe2r57kw1h6MhCmgUhTKr5BlU3bfuV5SAiCkqJufLACTfYBBJJkjT
JMe1sL02TxmygcvMEv+QNLnueg9cXE9jbr59v+cRszyUlOScqBdSvnclX0TcGVkh
soSafDyrKSu4Y3t3/PGp55GiYcJ/PU9sENZ+5iK1BRrI4Tnh3VnLMw/edOjpliJv
pCw30ng65PBYjEuRty/5mXSrAHwKUO0v70KdqjQVyezrP2q1SNoF1HY1DSyAvNAW
UVYvjt81/kg2XUYWk0rsaP98kpqvwBi7JpR72LabQKhbsPJrANk4+rJspGqn8VKx
+UYdXZAjc44puz7qm3QggW551gOmq2gZUyHMXsJ5OEzVtkRF6uP9ChMIXpE7yG7t
VEQYlp8RNB/mUj8fn9v/LUwgLSJjkmfRENT2B5SPzlnmnQ36tDVfe7/HgKEGpYbG
qh35/bSqkEVIcFJLmkEBbjOtHdkPvYOfm27ASyKuefITcMBI4nMDzMIyt8udzZpl
Aqbe9wIOvkCYgwsxxz94oFh1xF74HF4LcEO01y/IExRGFRZJPT2zlMi1nwLQMAMs
hYfj4vS/NfreIUwh7p4S34SAVFxW4cWY6NrO1o+Npd5YbU5G3zjRwQwAWQZ0ulJ7
ZkvyY95xRaAGx37aY6SIlZekG21F9SHsDrPzFNMhaNNw43/SPufAVFWBksdAtBol
n9QvtZUjB7xC3Vz6qq8ciHSde2bVnjS7J1GPbKnC1WjFLlen7trl31w+yEGjrjsO
zzMGlAcl6UGsrHEBYVy9NyQva+TvITqb8qN9uT4bAD4ZO3hLXD6pQmmJdTpye/9W
7wOnmDnf+r/LSlHK2sNdQ/IQMoKH3Rv+jo6yvEyNkiwbCQ+xXRdZEfHZojLH7InL
zOm/z73xYyRIrdGrkmHbsAiT1DhjY1YOEvhxjVdGKck88h1JJeDOxVy37DDPpyrO
eS5t2pZ2AmuodU/35SXvYVFmTZfm+XOYW7J0grUFOLjE2XZt4S+wyA0Mtz2dSRoK
qitlxKlJE2uG1p7UWoQe2e7/aeNz7tzkdqKAmr40lGZHcF1aWx5xVM0JJIBcnzgv
8/WleezXIoYfpW3Zy6zmyBVu1cfY5Gv26qkYxyAt1hi2eolHaLW4wI7dKIE6qPz5
5nneRuw9RZdZo2gQje5TL052m0j2n3CLppsLVOxdNe1tAf6HYhxnQELPu1VrN6J5
uL0xTlZx+tPJi+RAuLQ6bsYDfAG9l9p/BSP5fc6t4G66sGd3svWMi42t6ONwVZG6
2qNLlK2bhug2QBsTPYKA+vxK3av9Ajj1nQYaK3WoH6ovsTWhsl+7hMXEg3p2NKIP
oK/Q8X9VqhtdslICRoMb59yHzMZR6f/han26+unDYeCk1fmmv8lQo4fkNihOBQR2
5GT2Vb6umbSHXVmERt3iItRSrHtm1RYjt95kSczIP0z3V+CIqJLIAd+PVJbg2i1h
XAHASCTac0Ha2Wt50HkZfh7XJ3KvHEgSDsPBz4GWW5eD3UOXlMOSC3wW+H2AxZND
fwEMhDCBGMTnee/0YxNhEnPy7bBlQNOppxqI0A1GaPc+xPT79GntM7LrwvK+T1VP
ayUgVjVY2M6eTNKe6K3wvgm82bC43sulLP2qRhmeHBeaqRftHh8cfr2OaRsZe1HQ
PQFl3fPvgyi65a4mFKxNzR+Avu3DPaMEISxi8Q1wcbsdI7B7a91Lq0+bVYZbkpde
i2sK1mb+y9RQGsEKKJgD8ULGhH+FP4M6WMABEHAAKNAUpIZI/iaH/T9gbEkXygVa
I5tpskJY9zYiMMXxCnkAywekv4MnWpTmwb8W+a6jeTDY7DtjwMs3NR0SM/MLryWz
usAdgtyJGhAX98DmLCZ5tIqPNXlgB35PgsD5bQDXhLNctuCtbgu9ZcBsYe1yHZoP
qVdmb+EXeKMp0N2Zvzaq/kuycDtX+7chhcb0tjCPKVHbRH50TdZCVRqw/KzCUjpq
sMSoR5n+QGSgp0BeIc/vigugzuw6VFgHiQ75y5VMM5yZdjIT6xlUf8hAinaTMr9Q
Zp6VoEPSR+QhGyr/DCWKY+8Biphopqh27Ij6mh14v20dvWRDDBUcrdAuLrJfdZQb
A5bEDR08AW0hPEDshWP4FTz9vlw62QeacOMTfsmNX83kmcFNiOOG28JeVjq7L/Wl
gyO9eM9/nxJkh8eFD7Rl45DgRPgBN+u6Kir5IS1JWn7P8uI9AVFQ0/DNwmLsERFd
aQAxdVYWGYoioAfuHhm6YxK2ag6Vt0r1vFS/uAkT51HnhqPXAmkFJCFTP7w4g4ha
KgwOKjh5w+FjRswNMDA2edEOb83fcJfWLeWGgc/8fjBQewuSDUDsCWwn0AWUIUUL
RPlZ0YwFelWIqJEcNAY/Zqmn44hQBMwmqmFJ2g9BFDxAazvTNI8DP+mnh0wDYpjd
wA4T8grXcluS24PBLxlNYLrvVYIJhmEYhV9ze0TsIlKKXKkR1kg4snN/u1Py/yvq
iofk/t4tATaj6aW/eXN18EDuJA+LAE8husncinNQ5W7G99qjo7PJKYlkvXgTksSj
03OvhKtUB/ELyo1icONO2xzakHdPWBwjz0GW6D/23RD4qYKQgZS0bfy73pNXJDkS
ayCF1r7UsjBEPCrqUw84A5rYdU6VGW0YGI4g6CwIEdM+QZD76d3UkVnsdXefY5LA
8eXL1PJFPrVdU+Rdq0bpI+60UTxyX9pHSzlqXcLPC5Np5PZlZggRTSJQZGZ8J+wY
F7gkMXMSXKAQsv4JoMs6R49FTEVkgZH3T9o6qenRUMdBJ/0YJlHSjUgVrjKtVHOa
NaSdZTtvtb/eWq7BT4/BFmhckkRKTl21Prq4XDbvVA15xKdCy/gcYg33kIqnIeo8
jKu+2hWaM6lQpZbVGffhGu6wx6oeOBF5GEqyYl08zBLbAYol4m2SmTUHbm1Om5hV
rSR7vdS7Ebe41HiBNxTaOQFAgvsMPGL6Us9RF7gmkBPCrlh47k9sxFV0lCnJzO9f
apMkCPE1FTueydI9sO8gsd/p/ALzBPxuuqlMm/SarM0dVR68kSf8C7C5eJRjYqPv
nziQr06a1U0VHfk+y8hU891JqBXSy2cwj3bJdv4a7aH0h6UJzu8Hm+WZKP5WIIQ+
/dRIm84e5RmCmg+P2B0bTzp3n/oYXvXs9mFsaU2EVGiHhlBQ3zdnOxmls8b61tIj
UMD8QuqNRuC8GQytL6pqyJSpz/QRHvGIvIVuVSUXEAlz1wq5jCiBTL/JankVxJ1w
sNILWxa2Tt2Hlx4yzKD0s3zX7jFXrGmU1Q4XJSHr78sRkuYBmynyLbwOs1QR9w6u
6vIQq4q7KcwIZXUdxH6WesBnypTdecHbS5xw8vciaIeTHwr52qENJB3TGtvJoGpA
LKdsSFABLHi5VVRhmiHstw5eaOTtDlC/KdE8ign1gWbbqMygquegECBwXYerIhgN
CkyH24tFN2AMwa8adYCIJt7KXsE/Mq01718ynp3sezV32ndyx9dqx7A1Ge4h63lJ
pzLrA2dEuFo6iQoJREg2wLscM61JmUoza3hVh1mF2saV9FbHDkHCgheA0UhI+Nws
f5vE6SIHVMxJYe7uTEBrNpj2aIw/zPDMW97O7cQqVLZ63GQo9yIl128oACuKFbW1
0Pb0mUA5dsAy492HACDK44oWrZKqjfG3vf15vApsOGPzyjYzUdMIjlCOWJQgn1G3
ySy0+KMIQHWqUY79Ozs3dbEHsBLXweRlZ9az/Ubxlu4W94w379rdKTD5PyCT9mMb
q/GRAxFKaDI6TsCYve6ZmPX4Ds8dCKLpjJj1AXMtJV03teEEFhbGeP5/d2U/Ae5f
JDIOh3G+AWvb3DqSjlXhmCkELiEKv17xka7GUMbYgKin1j8SkejgmvNJ8CDEThuV
yNS60f2pGUS7gRGrO5SvRSSX6canwUWO4pAOVkB7g7eWV0926wBqK3TLBoBwbYfV
RLsDumPE4wS3yg1M38uvLEV+lYlmUZiJCnPcPb+465FPYRvQfUUoh6330BuB+1hy
ri+vUN55oJ38EmyYtjdbRghniUPzhrIB3fMprVXU4KNh2GkrmrsfTE1huiNOVAp/
z2oFdkHTxVO/SkBOPU7a86ulVlMYjk46DOyWDCXb6r0EC6jh7BlIORd/9l3jhNpz
Ou2OgoHvBBDGzIgCKZf2Kawpb/lmkTzt4a4sxwwNmijv9lNGAO4Zb35RurgmOHae
7QQ68oqJKNHHDX5L9BNs3jaLeQ6Aen7SQYqlr2XJ7G8MD7/0xIGnnmFEeGDJxcbk
EdpLdLr5xax1lESm0uK0NW3VZkjUzrnFtdqG6a+6zkFli/L6R/lwiKQJLgyougC0
OTA2XctAY0bFUhVWY2WU8UKfH+1+YfdU4VCDmSFUqeYNPw0h1YTd/ll8yicCwOMV
GXoqv5co8HB7sYQ6zsvrY4zSiCk6CRXwVNqjSI4NdowJNgF6mPF49F4HLZ5zxSsW
hHVGO47E6hSuuaqLQRTMnai+AN87S4y4wAqAPcJI/+FVfPdXP3Wa/IXgE1xvd6GP
5jF5YgkB7y7WjEnPi34dlrtK0TCIv7qnt5yYe+j5ndPYJJkezqiC3eASGpi3ZQ5Q
VJ5rW7X6nyuhXMw3l2pGMnvooPbIWeCEuwPWpIGxAHd8lZXFM/AKYOdL/p+ZtZbr
FRu1xaRyKogb1nSsdrua9D6SFFxueQScDpR2mCJeZ4Vu/YiuOHh7MC8b9ucvWA2J
XBmAWWwpGqv/NQ8HM+LpPxX2KravrFsjAuC9sV3rMKTocdcmm108/iGMe0yJKIX4
6h/2aPjMz4U32Ika9f5QCI5Cnpv8iYbq7I5EBuZZwAc5xQOZ6W2UuygyWa3hm/fp
DYS7ID6yqCumtc1ReRWbJ9T/5A5xSwndQb4JxeipG9kfVf8U63YP3j4INsOkBMXZ
/FRrwLTdPPsEx2Ii8POxWcU8MX2YBOtHEA5QckxLg0a9/FilxGi8s6/JVefOk8QE
kHRrz3NATkXFeUdwqTJ2YI23KWOPOSrGx4fRXmZBepKt3aZRs0No56DVjPbD74IU
3SUlTqEByQwUU74ptYicFDi4PXzhfehvAqMSuWwXVL2ZzmpQaKMUIAUSimvn0OYm
7FRPJM4HmtjwLQ3t/wRM0hGYIyU5j1EodusaUIEY3NrH8LG+wR9yTMYKsxRCJuwT
lURscaCJC4y20bgqhYwnj1pxb5d+ra/qNfOnPOX9oCTfknfO5Ty9neC8bP2XE2X1
6a6q5TWQWybcmuVLV66McIA4FxfaO+z/7wa/Laid3rQP6oIrexS1c5fy4yOzsV6p
0RpJqtzFmfOQ49HCpXE9NFpHCqpGgqnZtDmU0BzHX2Ty8aUlCgGtXJ+TcPasqXtQ
wYdmuqycnvZfyhc5F7Me/U177TuOAS07y3jx4K1cNh0DthsCO075voyIf2P6LVu6
s6RMMcbSLg05Cz5n8vhW7LRXj95Bkgq+EYKrnBw3f0TUMkC7EPZZLo+4+f14RVkE
B0yLucSwJdKktnY35pAVjdKiE3HXWajwnlYmOV4isAqJF/8JqNGJ+CDWTzTsfh0F
D3NlnT+8QE4fXP2oxtKILgKHvpMjp6sSNy3jgSm2gz/duXyCZb+0LKArtikJEMSw
CjyEIATD1mG6sQRRLKoeQQ5sK04pIgM582LvR6HPdTatGY4bqaG8J/nKOfnzNGbx
GTjAvyurXufBfvcic2D1KXR5fE5FsujI+85RytPRqui2yvBcJRH4i5G1j8cYkE9D
LzI2ZpRHPclXRonIClbCfbrbI6g+RyL2jP7prBrusYZlZaLH0GR6lCMSwdCOtJKN
0TFhbzmckkSu7lgO4XqDKvp8a4h0Cc3ooLXXfPxM4SiwWBnRSrd0l7eAx+/dfeVL
tLSJE2gAc3VgyUoToejfaYFuEigDTD/7dlJm93qnjGWLMNceOvC/edrVEOft4DUI
JUWk4xirvynA55RHUhZPOQX/8+GfQD/1X7XHLDd0JvH+OYAxYO9mCMnw+pc7TYkW
qn3YUydjsku2W91NJ/bJ75p063/0qoCt5TBnjOgUhBZ9Q/eLeKDbSGOXFcwBGdzt
6Cp1C7C1PObtBXj3JBaTzumlNTmGyxB1Sj1FfrnDxmeiNzs4dh6+IrVP1Kpm1nKY
ZxuXXHHIFqCM+YXl7Lp0R5R9UImk27PP4zFhliSsSeNIm3WIQSKNfM6e/jYYfZ/8
zeutmbHnkbIysrGEf7S0Vw7x+L/7Jl5fS+w/J8flspFW22SPaoYdCtFnaIDYQAQi
t76ZdSZvcR5N2ZGc28tbuY3irUzYNpO0/rTOEWJd6dHMV0tKyfF3bqzZkgnMjKny
+GAmPX3/ASGVzZm+44J7n58D1RmLg8EZWdAiy570YV0QLeFKH1GzgpkjbjWPEBR9
l6Vjq55CkE5V9Sm6r2bT+6E3tRWXr5S6LoF9iDagb08jvKnTGJ1PZ4syOeGlie5G
g36upDVuGqcILJqM4WihLVC/CJ5Z+wPQtjWBVQXMTmjkOviBt9IXT2YxGHMdTS1C
QMufK/7CDwmEe40AWU3WTrjycTFUAVYPQmHLqtW1V+jj/zrWMabAGVbYbyWfVLwk
6RU653oxe5HS6udCKXmjiOTgW9QLhak4WzlmbWU1Yxn+G+khJcN6EMg35Khk03WZ
gcMtfzaWhX8AFveT2pxHNG10n+HWhaqlsXoH1ynGnyisG8pbaL2OfWFpFFzw8GVt
P7z9uM+E6s/Bw5s7ipOyZHZAiBV6duD+Ot3ebOz/5Epho86CYWsj9SGibECPIlfi
jJMy1PKUaYMindbEhObKDoLhcwLCsQtU3/qSdCilElWaYH6chYUiK1zqu02dWPKc
Qi8yTrQc3T1poqGcRW3gYWolq2qnBH7h6FzpqBuF0GXbRaGq6KeA5pXDNFZE+HKt
bz2CcEursvV5P4adrgorAMyqYT2fSK/OYGdKDup2gOIeN7M+zsr+qXqRhWJoctUL
JRYKUNCz4dNp7OZYhLeyg7PkMCrzPkiqJNKkRuMbO/sqYK67k63p/JsoeivrcHwo
WqVKFmPDFART6Mhxvur+E+FXT8jf2Gre4n50vj/Mqr27bBQsTpm8BP6oSmvFQnOl
3Q9WQwMkJOiCyGm7cZEHa1xgtfDBn/EQYdK/eTackeNtMS9aMQTTxtns562xPSAL
baXL+X7lL/lYSTzSAgGeyvcjqIOfeZeAzHPtRn58kKFBdvk5PhMNVpCBpClqd0n3
vcPHWuA/EC8Iiu+ON5cSkMZO+diRNll/QUjSmU4vZG6M3KByKoeORjfBdjDXCz0Z
0b1cSJs71K1WlIeNuYSaSsZAeg/4ny1M8QiRAFILJS4+7VrfAtcX3wV9mwyAYEdo
bK8KHqbuQDyTIivfK4D+DRkNL7joqYCxqIG3JJ++UIyGTOAsXF4UV2n9eNmzGrjF
QRNlgjDKdZ/L5F5tp3GhuP4MASHvwKy9E5/vjRhuMFnihjsmCBOwNm0DaOGx/z2D
7yM2TTcw00+9RyX2DfHoe86xfSvxGtj9EbtrxDrc8YP/kXZfx2wKOf9rwzfMep8w
9WFMcLpNPKUxJ3cvKEZFFXGP2ssS0fB95JuoHJfraYj5i6y9tawRJp0AgdPyRBJ1
/Bb7LZVsPvjCBeEXKSkM0cqckuQZaknhc8qvkDPlQy3/6QY1xIqdXKsaBNbiDKly
jlpqlsv/YIGDNvuPZsQRRYAaS5hsg24FQn7YhHRFnp+4IDphsKZ7uHRkJU70BXqC
1ppJ/vSnKadCI9cW2rRFPw/vZEzL7UctioDw2+8ZlBhAn96OcnVgT4Zb2EWoKFcv
1D87/WVviZGwCshwSY2JWXNdxuCRXkzg8Q4GGE7NNZQSM+gfotWjP87UtH/9osrl
jKsJJ9XkFjaFoJN02a8oO+4L/drAwrAJDSyivbf+EsgT8RXtqwPRDnmbRLSnshKS
kMW3lBkV5yaIEnyS6N1m4sme/WbHiR4kxzE8+gQEkUAzlsCxQEQAcwNLJ6VVZOlx
2XiQwx5JsyPQ2hOteEsEhAlUEBGzoWRtfrhXNeOd+IXscU84OZuzn9rBV16Zte9z
2MQ502cnjunIPMEZeLwbR55RdOBD4AldspPaRFe+LE5urI80ei9K7S5yoHHDMwuJ
7j6uUdojQEyr3jyORRlssOJEin0QcO/WzIi/JKb0rQbUkM0Mo4pGcD+WJ56Ot1Hf
OGMRJdDqyijswkZzN9mH646lX79Q/+V1CC55Eb7VvbuuwGguMx1oYL08sSWQHntT
RVVJCeh29nNPWXaVRXN4BLS+33P4KP7Jurfjvkoj4VP7zjf51CsMInZEOZqUbzbf
6GLgqWS3Q7fn7OlyQnlBP+od7l+r1dGDUZIlF9kxaSb6pfQ5J741igPnfiTNvnk2
Yz9RVDC8RnDbijsVo5sEeHZPHxmCH0buMFemmEVrSf6kHihPrc3qJOOKYurXXXcE
kDNoyARm954VUHlichIef5hwK2t8LGRg4QiKG515fShcrFXnShvwiqNL3OQz9kMn
57eU/glVO7SHhn5Swly5p8Gidp8Q1+sh3jVnaMQw9EpYuMEvo9OppeSmHbY+jdut
NtPUAYGeIjfsdSgIthFev5a0CeBgi8n4aNfX1VoiO0CAnJUQadNzFJWaSjKGezSe
NboJBwaOXsc/oibvSLrbOxDfsarUIaNistK26TW+/cF0hmK44R4AEiWE99gYU/qb
ROcGiLweXTuenAVy/o20kEMLhStN3j1wCXE9OvhRn4Gytdhd1oEdh/3LTduHKYLe
XnWNwHkAyMhhFiAhuqA+gy0MjIfZH/nh28lcwcV8E0aJ35LnoKMy58Vq6ZwqNNxp
Ib5964JhQlXhgEwyEn2lPohr/04wLIN4QvEWzY1P2JEuKMp7AEh26DYbqykhDj2B
5PeA/dR4sGkmWNEIzokPFL6Qw9ZYHioO5gf2l1LbccKaDlR2/iZ9ZXdieHRPVTpb
cJk/ABRSBjU/4ZbIbA5rWdaoHwZCXhjZxaEnMUOHmwr730jI/4yBOL0OuPnR29mJ
B6HgCnaUT7kzG3kQ4GOUZK/dWIwmM92YznXjMqj7hWrwdgnbjtbaT+0EGo45XsFs
Bck8aK6oI/W98MNViF85g9lsub3hoakC5fmhTS6ZKJuYyopDa3I/GkJhQyt0lCE8
4iZvRd7OF4kbsb5yq8NdngTW+KhE64ZyFLXT6qKTmo3ThYXx/gfGsnUlibn1eLhl
HU6S4TkBfQy16PXJhuD8n4/7UXAZT3VhIg+u7bvyUDJByxfNuqeoijvTm9YgVmmS
+tBYnQy2kpbV7D2MpiA7zLJCbzSQoMtqeO/sVMzVa6me2CFJH1+cpvmdNGJcK1e7
vRm09mBWEJQqSNuoQ9kufFoen9yPmLxWx2dy4Mbekysy2rw2VjVork/8FHlSbldi
cg04gv65551a+fhZCtQIJd27OBW5uf0K/ITrK7Lcx/mg7BFVMvPIvCxAfJZ9hUKm
ju3oxT02/Fi8hzusfYjFuhK52c4HNUGunaV2lg/gRGhAeFa7alxa/D1rey97fb5i
Jz8mo+MwjEsDAPJzMQwS0Qd3/wA4G3vUu5DR2ThUz8lEJpGU8AWY3k7pR4HUlrJ4
hZ9+1FWk2bnxXWwfcgyhud6VvySqGw31toxVVY9aif1lgyrCcVqxNtQ5C4ueUzaJ
dRbWgQK9kNNWWk7EjDtqVsUlVal5jYL4B1alJpV+Dr4G8a1/io6IWj5uozehNZ3q
qZ2Aae8iAKxBF2KNL+ExkD0ciCgXLK62JAtiQwi0xtiOTreAEyHIT269PRlzrdXx
TaDXBYXn8sfkDLRypxoBBWb7RVr9Wh/O268dgBqhzkJsFhBRHeyR9DGJE6nFYiTe
NxON12MXOdbJhAcLo7BanxKu95DB0JMxXPtU9gli9sx8vaKMpv+wCNsPCnmMA7ST
/dDc9gopy4QOccoQVPB58AbU3AShDk3TZSKupRBvJkfwCy5peg0p8n7of/WS+ljn
BUW/9nHX8jOlh21+0kuKvYss0tF0jyuWgS5yJuazUPIoOzYjsfBg4navjatXTVXQ
M+HHUAa5AhIhDGwsWe2cigPsM8+CsaQZ61VuzglLMA3j1kUbXQ5PNdO4FyA+B97j
77w7glQuks33j8C6RWOWPmPDoROkJhO0s8v+Oc7hUf9uBXv3wnc13PlNAS4BMO84
PnIO4Wm4lybqkl6vrEGeq1Va7wQkRLdOy5j8oOPY8sdzH6rXDc+sxCxKXQRTiJfz
QkWgXNTZYpFQD3H8JJPTtYQOrkdabjX3QglL8xQissA1dNGVtZbVUB88s7J4/0os
zDemOtPptfen36DtA3D1WuyNW+gvessRyXtUoZtxBoSc75O9Z/4n5RLK/SNcJrE2
HUqxSrIVf2qU4ETfu5pnH2tDlpIwWVQqusCBN3U699b9VBdSqquuOQV2ImNbTu0T
mA4Ed+IyFN5QOU1lUOCNRuBjwBss7awIF6IExmWxX+3HTX3XIQMt+Ywwuv+l1GWH
UtPZIqfebn+uGDcKRXAAAAIZzTUdqiitFHRp9eCN2WCclr/rc/80//gk8w16IiD6
7B0UtYH4Gq6llKeZlV4DJbwOHZ/MYnkMA5j8y/eH8LhZQO7zyzNvJpQMRNfvK7FA
xRRyRwZ2yfxHcz1cHNyln504uH+SQr6BRetoB+1vMUc+zd+clhyLWAVQJH8FhnvP
piuZCWvSjgtW63c3qCUUSqzjp45kAGScF2c6omdbHv8nf2ibH4t59go/n4yu4TPL
tJ2rBXM8Z10sePv64YonrF0rXevsKpvGxh3OYwt+tXRYK1Zd5V+eHZ0VDTQbM3U/
JsSrO2lxjSUlww/eh0n589YtCe0ZakEqhSIx/TXEiVz6XkruUkqXlUPj18M3MLcN
31lMLvGCWy3LGeS94OCASDiCHj7qSZLhoak5ePmNCFY66AwDE40av9Z4S1mDBXm3
O+WeT/NpFfTQLe9aIP8+jDmFThQGBFRxk/JlWfm6BZqcqZSGMHDSsgLCvk+H9dHY
xtNisOME73mQS2eOu01z84NsB+GMdJauOU/MbvP53IZV4L6/xryhfDGYUbf5VBq6
SOiss/hRU8M/rWhaxxlzz7x53VHkp70CCXA8CojyrYvh2EPdtIRXRxHQuM6kZgr8
C91PJyK64N34aJSbOSJI+7GWWpLYUMYT8llhMNUYsO+KOvGBnHY7lXYoWWYDKECY
3I7J9fVmKsxM0ebeLwQbgP28hHbvoI4Xru0+Y9a7BgXhKSyEh42rYTaqgBf1e8P7
ZvnkG2b0vx5WkAEcdvQraAMzHVSw2zy9X39uioQVDMS162ei036RvbrgRR6g2lIB
D/OPd7UoqGK7KoPe3yYuOPXNHpD1Il/OQ7HPBZmlRBAnvWIyFzYP3ouf5+yT2WZG
OwQl4PWBfU46zKO0ibyEU7cDcOcyM99GhFFtjUGI1atFCE336Rc0w7emp+nl47Xw
LQYb61sqhRB/WVJ96Z8fWR63IGXxlMzFxzPoFXWy3UdEdS1tPH/MlDaeD/VYsTfO
/sDN4TneShUaSmx85gvSyHs3e4wi1z6mUOaR/oKnNHrAOYsnLoEBA3EnQg1IHCjL
Xu7TbaTZGJj5L5B/1u1bwakuC0SYDVwOa5+G6mGwKYOiWQOVcKrIe1jOsBFnfg4x
A1nNt1YXT4VSy0bLTcXVnwhfufYTHUliHgitwjzV2czel51ib8kH/CVMDVqZ5EvU
s35BElUyEYXTQzfyognjPima61eRc5vFa+cydMkvqQ1ndlx9nEypHTzJD7t7BCmV
XMTTGUsGqd45IjCGMSr2dJ0AtvNSXCVEY3Rav7xOfALjTPTLZmUvQRASV+CdlDKo
kVt0WN010fziH4ilMPtJlqxcDgUjKtJxOJ5kP4alYFbp07Ogn2NBEH3x5168eM7w
NIqmhCFnp7wqYotLmcMsn7BeK31fSlCjX5Bou7n1vfY56P+4OMO9hwV6l1OP8W2L
I/FENW2qLnalqvDiMe0N/pQksvG4lmpp2u5hcfY3wtud58M0V+QivnW1A101QZpK
Z2EIfPxJAVhdvRriSu9byfFZu0T9ts/9E1IT7H2xMgkBDZiyxT1+RiaE5uSoab+r
rhmbUgdel5ThND3BFT9XFiEQRBTIBjkOoM27rp1Jgy58ri4utEz2I1GCnVK55iJY
CEVTZfzryE8CjKCU+1JSzgUeZK1LSuV8iqdvqa6zD55XjdVt2q/GewVyMEewc6/d
JpAvH/k96T+P+tB7FZoCuMme4sqyboI+d+8B/WlvGaujDeQxk7w8NEGQHSDED875
JQ0gKmy2k3c8ZnpLCR2aCvrNK+sqUw6j7bYmb6h8Ldc2/8IVjZaWL9EtuqHFQ/7r
T+g7NKA4FoCFbNB6cBMxCGfc5JUPwl086OF6/CwSmxhyQY5r3NMNrtMop1q0q1A7
5tCqatodKVmXProf8t/L0GwogcET+KGdCF9DSiJ/DdQe+64A/Jo4+nT+AIcx10tP
aRMy8cJcy4DcRz9/zJWe+Ggy1rzVy6ab0Z0YKUyncfmsOJw0mrEPPKD9RS71mY9E
dclOtrRoL7b1rykMEHAzJdIH5k37j/uPRFCxPhCH6whXyt2JgoBnCPne+hs9MPt6
/VeDqygBRyLXK+cFj3GEHM7WthB+bQjUEvIn0rVeWnRebpZtCs1nFEAYTF2fH2Yy
/lQWsvo2rimEiGzXeTQtQh06fSCGAeNCg57B44B/Agr/4WJbLBp66o7Pn7bg8Xc6
NcYUe+hUPShp81NRVqzKhtj/o4IWnmyaxIA26yboTpV7RuxYN411ZOulE/svSagm
P04RfTubGPZg8P2y2t+44iGZJsiE0drLnIkGeYjt72puWSb5zjQuOB6dpca8teko
ttcvz3+SnKCQYNMe9hncj9tcGNr8S0kRAh38s2thM/CcUaZ17TM1zsgTbTiw66Ih
YM6fusdg9XOXdcp9weT4HgoK77qLz+d+4FatTAUmsrUq+6jjYLD/rFGXfpf9XWSM
ew57v9OWoz6OrkiEr9eNhOgKg58YjJEEMXYVLOXEksKX1/K58AmFvFXzl3RSttcu
s33yqkqwq4aDy2b6osW5bn7iFpfY1T/flwQJQ9xUgpQQb2bDAGqJ3s/tHlP4WUsw
sLHZiEs7L5asyXDkEYEW91kxwHMRXxkVLkQ+W9QkMvStNsTlifLGMWnucREd2pag
NVWa2La8zilFWyYbLAHkmNOur+Xeor+b7NZ2zSyrrpGT46StGdHfMCwi3l+53nYy
Ym79ST3IpdFb32IgjGNLnqN26V+k1Sleb6i19am+C4tvw+FuLhd7m9qDFDvo4JGi
iUl2qwN6zAicTcpbsR9E68BIj8qw+I69kGMZFylhbHP6RKz48Ej7dOULCFjUPuxx
8kQNN0nomj2h8QsnDtUB5Fhs7EDH8wmyFqxJB3dutThiyIzsZ4Vjhrr5B0wcts4d
fnIn4f+yNTEisQs1QVfzZUsgL8BV4T5BbdWMdb8O5/xZAQLFgIBJKzxQnD4s0uIj
fZAm6yRabLyLy39A7kkGaY17BgoTDxKC5PcgCLjRO9SARn54W0ugwUcQY/y6xHOd
v3D36cKnol610aHjQQ43SbwBOKUbD2rFkRzDu5B1iimuegyF/zj+ach6s33jaOa6
BZg5xWUrWqCZeuSZdY+7JNQ7q2hnMuRte8iBb5N5CxvU8LGMaEE6MJSRApmQFsvP
FPneA0AOuLpUKwZEtb+E/rYl6jC+J1Ty+jhNEdXHRglvPUq2aKcGaf//rWJ61kZy
b4Pgvada76MXO6xHPomyG8J097yizWiCrAqvBj2A1P6zbLT/LUy7eqa7w5cMRa/4
+KZzH+2oR47BE5H+ocogA9tDLRBA18zU4xu1QTJu23Stx+nuTv7T7VFEVcr2O4vc
hc9IU4lR49zrBCNRItuoDy/LxZQhbSgDNAspLet985mov1TZ/DdVPCHb1Wja861b
q2o3RoTWXONagrgHKUVHRYlYrNSOy/S8291b4g+NqEkYV9XaEB0EKhpzN/NGtjtP
c9qMdD4dU/GSNcif4dOhQXB2UgmqPQo+UhDKbMFF4OoD0E+IsXVesZ1EoDgcw+1z
hA3DaBUzsQXMB358dyUBYil9x7GVX7S5WhU+WNwIWlXdF5v4qCptna+9rcZeW2Jg
/KyvNBCZcTKJ/tqFap5NfKjmgKhLnFtwBBJx2E2HQ0gNGag4lk9qd4yFJQM8UkEq
j+SUeO2eIbi2+8OpfdrufQ2WUNA8pAXN9gtq4LtMqD8WEtUrUdraGXkm0OApZ+KC
qYzBON5enzRqXn8CtQ7YON8Ca8A2yqfT+p6x//gm69DinVDj7ODH1E2hMlQthXRi
H4ENY0a4gOvXxYafKMbylYf6lRm63jL1DhUaVsz0o5DkS09j8Gk6FffaOzD5m/Os
1qPGNqIT448T0g9i9oLQTSsaXfCT2Ao/Ia8Fur3OvmO3zmlzQi+xtreEwRcFUxpG
7Foj0Fy1yvPf3xMDjDkGU18WkXt+yMPJBjLq4Hnxg6oUei91NyHoYS2+6BnSVuOC
gvr7dNHMlz3PEGNC95PLQkPYBid9q1Mb6ciwXSSCQDKuNi1/yFs2y6RjgOIPxUg3
Nd4fw8Fh5Ga1e/hPSzDORZTxTwNbLK6f5LX1z6OL9EfZrVsKQV9tRs9TDCCbFPdQ
ng2WX50ZGQsYiOgH7vSKDPHYSlqTqtdZX5a55LC8pdfCPMFfD2OeFfW9Ie+L/e7d
9+uh3DOjB0mofstO/z0pQD+3u9X2ldRr1prGMYIAFyKPAIKpfdXvKVGfYd+y6sA3
jQN9b7I5wqc95bkz1gQz6dcKYaUueIQ6vFPTpftqnhPBA9Ew5rsohmT1ynbcbhLe
NWuDoB7UDe3oiRXrHowv1a+OswqiKMvDFgfMOJct6BvSTtVo6ssdAKkl0lvGYZBb
lzSWsAXhhuDI1Mjlc9q/OzGegulr+QPebpJ9wMN4GGYepT96QV2mpnp3b+NLe899
eXDPLb0fiAVPAc8cCp+DViN6Ms4nCrhXXFZQmlVd7F4sZrZaMk+bcsZVlSzyA1U9
qX2SXnagbTD8bCUiw+0cbiIevz1z+TlxPKyQy9neaiD3cWLDi+XCdEHZKd5a9Hwd
xzAzFIvXICYZtacySR73OrFmFeBZ5gQeiCa2vXpqevzGKduSL21sZct0Q53IJ50k
hTCn/t2i3HoLWszHW1RlXJeQTEfC8+tPtwtG1q+PkwFM9ySf2xkdDTU8+e0OQLIS
DcfyioXUp3Y+4EQi1lAqr7iPNqBVbfJxZrV+MBizy3YP2tAj7zblxkAngDWcXwHv
SrdZ9Lzuezw5tVf+bXNvvvVPtuXEXdq+aVTDAbfr9pE9uZlcWEDK4ebcG7Hp6CGu
EDaTyzUdc8t4yF6R1T7qHO/3vuBKxkQqaPIBbRnZ5+QfSo472bD2krCdYyt0TR6R
x3HJitNAbFJTbZyfD1NSR9jJQLSLHQ4zdyeiKpXAzuXcglHSTshTuULM8a5Nbl9x
ysbRY8dmdho9BC+Uoa9k6HOS2C3ewxI7Ue+B0NOZ0CaVmSnX/H4PF2qFdC+Qkvco
l5ApVG8CbgYv+Ex6BI8Y2Sti/8pQi+jYlbqE6pQK9KGrZc1bQvB/IZqWO3aQ5Ncl
RsWkbp9xTE/Qajrs7U+o2+dFZWbeJKSHI/ICmV/H6RQDDs7ip1Tmw3B1mU8Nil4k
/7rn0uRRVRVB9yWnDfiN2aCWEhDvxm6SQvznZ3tNawPEeDoyr6Q23APydnuvqNtm
dZgE2P50OSRnTOApKnt+fMF1Wf/bJ9SJsxbxPel3AXJPYuqXuB10O+E9+h8n+ClM
aaVwzyQPiozDQcgZUoGktb8aBgUDmcE0fIqiHRAAiTzRO8OD6BM3wWJGuMtmlvzx
hfYqUXCpl/qoeWCNkEfSQnsI+AjlXAuQAzqErUV5i0SIHgawKwH/FQ5tsDV79wu7
oJoWUMwNi8fPsM2oMtKNQcX+j+W7MfGHVY7xdZnBEqIg6iOjvmgALlcI10S0lTHS
a9qNRC5/aCgZxm/UQW6qSI/WM09fP0HcmT7wxwZ6eCMu8rGWo02jZTPToI0z2qhR
q6FWUCaWSDCAdsNJunQctBDyyH88Kih+MlfrslesjF49mNiZIzDRqA/WbxJK1Rqt
ZZue1WO0DzvvVrj9kaQ5I8f+ybDgRkIbjdXlzC+Iy7ietDgPauZPX16x7lwEsWfc
9w7HxpjW+XFpCDbqmrqEGLt00s7LZKC3wuuXx41spDOoIQu5WKSBRednlTVl7sf5
qH/jglLxMYSFknipahULC0BBK/SLiMaQRFJYehZc87bV8/gje1OtzjSY1/mPZO7p
VHCf/ouu9RaKjJmu7EhCXzW0i+C//5bb3SO3IFi6e8uj59MoHJFxhZi3aqzzaQly
vSnCwR53KT5xHqruQ4P0SLtnIguMSoiI3uLce+pD/eUezgiLNOTXnyzlzubfFeeF
jNmvg2q4Zvpf9l7PHuh9vl+aUIxh+MXq+6W1MfgNitlWDoQpC1ze51vtNV//IfK+
NYlaQZ5Xjjq+fNPdHopVRWaBeTl+ugo140fyfAv7RvrLtpej1KzXTi6VNE63Rtm+
/tgNys9BpR/9ZmkiBe7aaSQVFsCSKvku31zfg0UzYs6sqbv7SQHeP7r5u5lo0Ccm
BOEelypRXYY8un8+OfmJijG4yYK+IDK4Qqji0U6KVx1lxTuFKT/dWvLTs2XolQov
OxuW/oH8QX7KYJOdD/wT+21rmfr/WKEuPv7dBzXdBZmPGL5Ow9oLK5Wfb6FuLfvc
4+R82cUPp46PLjejZTAT/sw7IUu6a1VlLfIVbrYZ6//AfbVUkZFRC5L0RjpNvphA
SPNf7QXMuaP4OdWghxp3ro7itF6gzPoeq5pvU1lgGDLC0UIn5oU8vis4RrRqaUnL
t1yg7h2ZGd3ABllilIRHkSHkbOfd8s88K98tQkJBDmzOkim2IoukwHRV9CAVdCCq
9mOpO9gr/uJyJWJxrZ/dKA5YbYNzhU9GDOvY9aRqlJreVyVGXMUiSvCt/VtQhwwS
6o/YOuD+IY+Hugp+uP61xW3AK4IBTiM5v8bOLH/38omXRHADdPTK/j7keJePrH+z
l/JyPUgeBqf0vU9N92ssTgSAek2wks1T57i4owFdYXtKBruqu2KkImBsNvSUhE/R
UWxnK82yCRGDkhZpb8Ckk88/lebBZNMt0AC4hRR9ODuExmpulIt1F9EsfmZranWZ
BW34o8gnYGgV4/0cTHeoTKYnI8BbrNJCUOD7AqxiG2YtvHNaXVRPhAEeKy5K8ZBV
MZ3ndeZ3cc0NjtiRG07kvKQ7QpslVV5dqJI89+HnjrzyFAFEKz+HENkduck4Pmon
qaEhPsOaAYV7QoN+sWBeTboB5vooVuMbTzU+hFGDiiXOqvbk1FCsbglvIr2fVoBP
it3+kSRd8WncAbXwcM50AXLfU/Rxi7VkLQRv+HEgz4Kpweu/7cOmOFmRxXlkFRMH
L6Jnva9vKeTV+ntCSpgq/kldMTzlNMjkAs87bIq01hXoz19gu4Lf/vlYD8zZf+g6
bgztFsysJI2wA7/v4CiO9RV3F+VECeQtYOM6DWdH8jRTUt+WTlZ+NW+xC2JFyH4j
3qZ+RYT18BgSSus/PbOoDBQXJTWCng3B+7owLSckfR5XxVp7evI5Pqagsla5tZjU
isOlKVbdJWNk0lG4x63xTcFfLuBPt+cADmwr14rDbLcdq0ofka1PAkrwOtJrBpYg
sCVaQfO8QojW64td6bK5Jd6vDd2eI4ci48a4tFxNJBQhm6BAYo+KQLCNQfHpHVJr
uinOBVHTte87GWcpDNzU6HVTk0jBrSpcMU9K9o8LJXE7jAehx0cLoc/OOdM4x0yt
qtNUN410y6dacpfMpQQlKDLn/lEIXlnbXXprxtuKj6nwE+AVEi0DYee+WJrmj/nv
6Jk4uizdZUbo6HOeaFgNagFQdj/UxL91d2YnkctHw/D/wCS0muDRJOdjOTuSrHlM
rckwFoJm13kbUAWMgwYNidacypuP2FbiipYmZNkUDTCchXllyRS+4lpEHBXTBGYG
Mg8JCSNd47pS3/UIV+afmiKmWTmr7P/9lVFeITfNiHSNGSSDrC7VYEAB5gi0wozk
8Ws004VYzox9dgBW3liTadwS5/03C2xhkfqSJ5w/8spDmd6tfKPsJG2MvBgmV6ff
vjNs1Gw4pUPRksNpm4DgZQTvtrpampR5OzeQefIVnfmB4cl7bKhAkrdDui0azWB3
Fi7j7aYIj1dsW3zs7ncWF2bN7sYlCwNRD6vdLkM6bU5mndFwyO9b7B5hyuKMR1hb
XeJl+WMR4rEB9ic2U6slGMnM68yGisPuhc4Zh2UvECelUsCPzfHr0dQ0YiYI76tv
kXVtucrPFWRjO62BUa8CvsLgHvIM9qdqfr+7wOD601b838OKOkBYRYJu8MMaqf7K
D0OQHLOC20XqzH1qRbJQo8p68qGHutq5ufaszXM99W0GEASWqS5sojIclm0EWYTd
eortlt4Er/b6mlueZwyh5tsbr95ERzZxa/XzMKKYYKRRW0quQ82H23CtTyA5tKjO
NAGg/V0meitO4HhVEwzsGPEaVaDYPl6ZZ2cUOHSwhBN691PI5H+/XfY2qMEsBv+y
DjAZUqZtjr6ExrYCYKmr1OT+yT9AmRPprTiNwtc2FeaS1RyfTvUnQEzCjj/gM7K/
0LYO5n4T6fA3GS0XrRRK0gplDPWZNwn1+ZyJfuJTgkUXCP8F0dDSapXwMYBOuAML
0/SIurZfFhja99VY9sA9ykEnD4mfOkcnuA+EGpHMw0kZfRz3fOjMnR8sZwH8tUBg
B2n727fYx0IHbqXxn5ERpjMHH0HEaeXLYjgMYyevaVbFvbZfjnAWGFroJSwPznyD
Y0uN+4yIMFLMEvjVMwrpuNmLg+uEFWeUi1xyR4g35A2K8MgNKdNZHtIG4h34oPWW
BgcKmMXoAh7aondyZUjxy3iYAoIgS0ckud2PVTrPLLC6DMWJgEeFuE094anIn4my
doSCw5CWTvel5f1TDEBrv5TWCaMhXfjPDQgT5SMnCDfB4UhXhVXIRP3wOC/8CJ53
IBr10T9vGwvrIQGKFpI3etf5vBt8p6T8L/8TkQGe2IfLkUY/YwWqXiiMVBnVHTrk
zHRGogGal09Yhvrps8mgu7vx+d98FLPUkhEB0CECuxOHQMDQWcmD1HS3t0TecjPf
Yl5vYJis3DIEt/3EAM8sIazpNRC8/BflaTeaGwUGmAzopXHkR8eTcqkVwBLD7aGI
V1qlvB99+4s9F1Ef2lG6kwYb1PZnc6jC1CqNk0ALJNulcfZwmp2upjayN/jNV8Gb
qMJ1N3iQQkbF9TMH1Hm8Xo2WBnSDnVFeTrfyNFWceKLXGmZUpkg4NI17QXEB2qI0
y2hevqmV/Pk/UcMf+TPv2ZBn/ycTuQlp6UdFLGnd+GwHLC+14GFV5GRHM50ihBYz
R8HMt2eOEAvcT6F40pCtKW5hrCvhFoF+uwfANFzgk3QytpdxTyVYMrqYcEwGRNUR
uMJYrMQp4teYL6Id+DrGk4fvvbQoxyNZG+S//xkR+NiphWTADoFsIVIPvZCPs15h
7zXe1tljpn8Fj4E6j99kdRSUhe4O6jWd+/iYojFoYAi8wZren/lpCmXZ5R42bTpA
FZfgFGrcnH8OiB+h1yOvklg2S2eQh1UOrwl1mHhVeiIk5Xz1pKN7CfQwrRzLSooQ
F4BdIgrvH/csW7qzsJKsHFj4TBI8VIq5j9RjeWDtjUJSdlhxGsBRn9toVpreszM0
X4VCgx7ldaosANJKj46G7MOclM7o+jbNvnCecXkeQXmj0jkfb0wHLd8SDC3Q6IlP
Wn4oREEz2pL3tI4SashcHrHTmcLPufgyZPCehuGcjIsS/WAuI3FkdNiXGQ+yH3Qa
pYd7woNIBxBtZaIMpLmHzrT1j7bVSZcnQWVMvgV52SbHnlAyTiZkwpv2NliQprG7
1Df0uJC6OH/Y9XESVyEA1EL8VHi7AsYmhViAspiYya52zy77brbSF/2dbTMHBgTP
n5gjiN5T3j6yOfb4V7wLE8iPwxdtH3tLwtKjyCrD75J2IZ25pNc4kG5SlI2nRMEO
bmoSIByJgM44AHCYU6OhsL9GQ2XHV6UGJYsaNhnkRbYmN1KHEH/EerUeF2JWex3j
0T5kTUidOuKX5ijVHdBElljchy8NnnnBJE4F+v81cE4p0LU43y+VecBACHJEyA32
Rj0Zo7GIRZiwqM2SecC21JlvkI8uVTmOOCX+wFAzLRUunzin1rZQ3GYDPFTtrBVV
KnXbDDumm8b+AOcNhr410wTG/e7AdSaqOufbZk34EmtLyOewucPfngq2vf78MSkI
73v9VChPG+eTYDs2AXnqOueH/3CasiePiA0+G7Wql7RALXr8cp+YsVTo3MiVFtDn
Rdbv3F82IMVnGb0E6IPaUC0I0zaMkhqdv8FR6wlkyKjZQpy67YA0KxJYYm9XhBU/
3uOjEX3w+Mt6iCWQxvqFrf8RO80Fq2rm+9MYuLcpiixQIe9mr0SvF3Vt1V2bJlHt
uqUWDklZ4wMjt1kJe5ziSRFMH0VbD+aAJPY7oBUPlhURruPOvfaPztG9Z5Wj1Hqr
KU9Nwi3SFPkDI7TZeDR7IaYr56C9Qg/RI/EL308nTUKqf6ugEMGkbtokl36G/JJa
p3rmfHvWyq1W9gLMMZzy4mHyi9exQ0y+1ULo3babKRYMp/fYnjGXzPfMPh5c0RU1
H/cl0/Lk5mmK0EXfSFmAAsX7mFFw2RR32laHgjCCW/xVehzDiv8dbzOFiJcUZdjB
CDef7sWXwNbsg8hw9NiohMd8gAdqXqHcKziwY13oBeeZj/+S94OWdZkQeEhiNkN3
12LaLzIAV8RBsDY0xvF8IFoGzpYN4BWZ0boxg7ZCBBlOtOZMzKfKTJ2XAFlxcxlW
OeDYfgkisnryKeOe3do54KYrhffxFvgvJ4ZXHL2Zzyk4GmXaXL7mPRas2fQ7+DR6
DxqV5JBxUv3s/zXp41Gx9r21AV12W83dDKrSoCx+ugxwcZZKssFKonPd0RTOLkCA
FB2W/uDPk2Y534nAfhm7GWCOIQ3qKf68mdOHV3RH4mKxCdBDpKYLYHWYycUyvBST
CwtQD41r8Rb+vP264weRTWKRgLFovGaZYw5tbR7zAJPIMRxyhwTarjPRwokYWEDZ
KD6RRbSFF+1mZqFNwL0q28YTMT7AaLy44M/q6ef+SuBkGPOeIopC3yiYy8dRx1pC
bLf4+cy2UJg9L88Dte29OG+fOJsHNfo8zQVspBERGG2gjlyr8LzbJ5FYXxr7pQYk
7kI03sXp7xv0/QnkKG42X0Cm3YtB4HIYqsGFxw+ug1E91H+e6fwFc2aC2VRl43ti
TvNiD3TGd9Byw540KOVPyf0jhkqk6VBVdJJx8Bwz7+2zllg2pmdULUyZXcU1HnB2
m8LmeDjL1ZWxradM6aIU5AMm8eD4mSGHatDnskK9AIHEuy1uCDKO5OVQHaFzDqkv
BpyiwjXqdf+yCxtqyljcCJswVXm0oQCDNIzRgBRJY4OEDbZ0AHaPC2QMnGhO/vJ+
LSyznmCZDZGw0gPGQbadgDvVpAlEIHbwpjMdd5nDhVgkHdFETdnbnO8fxDZ6QY/o
Cl8j8J1Z+k3CZKcRtXnabHq7Xnji+Z3EAz5JeH+YGN7PQ9XoFfkrvWXygIfhIpKq
xWB0K05vEJ9d2WQXmhaZucFDY5FJR7wxeqinXrkOHxUEza/B1S/o7lec2vNl7iUj
blwU3c8FM2uQiSDxOJg/vgpBQARjKIM4hlAwY6zFpkKG51SKkyx+6SlkI77XlUdM
zCydbuqJVgHIjjjn0JzpMgTkYJmtCtpfSFUTobK9tWByIpABW5GYR94/6pqG5hO+
m3esGIsH4Dcn0eIaxnXUjDrfeV9P3YN68/W39vuIhENZCfNXCILyGi8rzskghByV
0QNWt7KyEdZe3W/q7pN78wed7xXJ61jzY15DSiFEaTtc2VH6fBULmXmkcPL/GcDO
uttglOBsKCvPpdoK7OrW43CqfwKFlMTe5rhU2En3AGPNGl8JmchlKg6YutoW3klp
ilEneBQnpHkbWiVKSGXJHJgOoAS0BNJAWOD/h/AJd5NoYo/uMKey9cwrs4V9tTvq
MjWY3bt40ylU5lZTEvc6M4fqHrrY7uZPn5LoZiDFCGuiMDB8txeZqKS3/8f/9igz
EoTpP/1myzugkXoyM0BGJichXkcyjcPQAHYt9TSYG78M5ZtrV68dfzUjE/c3Smb4
223hYem3F9pQfcykA4pf+b3GxBRfxIyuwGufZrohx0LMK+zKlwEAvzS7qRZNjq4h
ex8qkhubFYmT8EQusGqKdPH7I38wcfYxWcXbeEjPysUHoUI36k1qu6PYrmR5xajS
3vd3iFvd6OTGmz1EpLuAZBEPHSDPUcpNf14Y+uPyBS46FqOEmau0NuKwdUg/wSp/
EAUE64BoQXCMDHNWLtdVlqw2jcapyfJrWYhVEbt0taGcK/smF4zycmmN4ZOPVpps
ZVuHBkRGUyScF6HKaahIxwL6zI2J+0PBJJ8uZJZ3yYRuhXy/AiqPKhoJ+22WB6aD
Dl/kJVm8JV2B1a2Sf9yIgCA2AaTZkOWiNeKMa04krMcVQBCWMFql9uQEKSwJPZ+e
EvJouvWvynoUhqHjtAwxsStIt7HZfw0s5Y+jgPlwvYnjBsqf9V6UaYNfMilsJKrP
Uj/beiG4pF2RU62Hr6Cdyvdqf01EZr+z9ZEagWWCBdzDh+ypg3lL4baQWHvOMzAR
jwU6PUa5MrG1t3Qu7Wxkr5sw6Jvnf0beWe7R/NdIL0xyURlQY8oK1ConWhXobba1
L7C2RNb0ZSNX1gC7ElmV6q0KA8bcx5zdZBswsDyVRSTWzIn3ayv+jI5qQMpV8/FH
+izNt2kbiOiZDUVTS50yx5+O0GavyXo7NKsbIEfbmJdKJoyLQiiRxQEHUCN/YG7Z
8e6mOgJD1zxZGf9MzkMMML8AUO3+1ZY8bfyE2bV3C8B0BB2N0exwLYMzePD9dVPA
04Y2OmzjqaP4+KtfDHUP5spqHTM4LyTMnPU8xlgb9zpbSw+LzUHtv41G0GfChumW
UzXU92qHhyDgh7EB2kzrbHrUccwwKnV/YRT8miN8zEEWhRNv1KfzwQ0T7wNtKcRy
biv0jDqbUPiDvRDIVHBlkRwZEzl4FadNu2pU5TTYyHBJ8dJqx74sOqNZaMK4vYJI
ipAAeBnrw3yQHDWDVDW4rclaz74sp6ifF1CbJwEhd8MpZMJp1OxtdKmIKZP2OVv1
RCMS4WSQSuUNGp4nGRoV4GlnVW56K43OB+xJGcUKSf9fPBE+Z1jL2uLSqYfbULVe
AbkJCpmbwWdPH0eCqIiw//9KojyX5e9dhybePtbEVTfzJVpjwhWBbaqsMG1zMMmw
RheAya6N16rZoZGXJWy5kO7Fkpb+dbm3LiiZ5a6+uDo2l/to19rp5gjNWOKNVBRt
3jo7vk2yDOcd+yau1fIKisH0T+P3xJLua90oXz1STOwjkpWPvjdtM04ilRRktWPh
a5QExIdjM2ygM2dHMsrhe51cPyPPGtVZGvEjFaC5yv7Go/OYiw7r7DnGmVQQDTXO
ZCiXPJ1I5gpLachiqUyI7CQ8U+1KPF/MKRZQc83Js+EEbdE4/yisKUwifbt7tmRk
RXgWbNO/laTwW+2PVi+sPUQ8U67kWwkPtqptKvLhD+duMxMc+khwWSCl539Zg+1+
T2VDFO79meflA/6e03tsNCJmOnkX6muKJMOCh6vFCgtkWoBHY6u37punshTbHoYA
fgoLH0PcXHfvOUkC4U4IuzYeYohkaZ1/zByg+bfsgec1YOoZWQrfE7vKsF3p5hy2
SNnJ7soXVMMrsaB45vB+R2BSs1I3a+sytKyqODxpNN4HP30ifso+9nNqJrJvqvBL
y/ONT8XzlxJHXK3rClPKRBKncXwu0GcWrf1n5JNaLOgog4W054pc7taNJJBg8VkV
uHM26YnrgxHb9wgU8K1RXb8oXdAl234eNrq5gyUPan8WWG4d+ctkxpjDT6gV4LnH
u659DkxLQ6GDZV1mW4Zi2MhqMpj37keRzOWDTzzC/1oT/tGMASrF5Getsd7T4R+l
uMzF7Lm2fVTnVzxVoC8NbtnguSbo+seBHMdX2b3wf/F92T43E4533UheqbgXFh8x
k002UFFeKu+e/DURdGZKS6BeMv9hBNhnyDlL7MH2LQxwZpj3QJ8cl3Di651BQXbR
qvZGU5J6i9zsChdo+TotES1OQvnlDYjcHF0m8kOxjwEjsrRSjGiOR2BcKn76mBiy
L/u7nqW6Qv0vtvJxbgf61/s85LDGZKzV6OgOzC6WqRsZNW/cineOQH3r5EEkkdH7
B7bB5+LYBF7jxARPIZ0dfyVJATYD/TcylB5H4H6R6N9L3erQMwgBFhZXFFTXpnO4
x3Zn9x100MGcUQ9iMJ+jG1/642XL8LkiiAKdJ6ekc2VpokCQNWU/et+ePw9BRUge
nkbId493M3S3o3ehG1UmGIZPUKtQ7laWyw8+fQvuGfiV/+UI8XrhOFObbzVkfYbt
jYjzXd7alSvbUBlctskngh2yR6RANNgE3TVQH7v+8tBnuX8vGzJNRueP2w6U6WBM
pGQy5gX+8fVWPP2PLWIYrANdBgs/bZN7fQY+5sKsWKG8POmoUTGQpjrR3mLskuf/
4dMS/clyxVx2K8Q1QHpNpPpEojno12J+yvqB9kfBo4uzr9bY6xsaPa4A+4c4dX9o
kfuxiru8ZYfMC0daTOcIex/fBego90wTrBe66+EW3hA7EW8kigIVoFMKSexQ4AXc
1jeIjfeqWUyzTaiFZpwJpk/ijimF5mSwXDgKFG9d2KyT+98Yadpr3xqW0bdmj2rK
YUaUWp4nPMgnQon6JRB+sICukTvAsymecOA5tz+M8n+g6HL2jqdNaL6A2S/PiBL6
E0OS9CraLDeP/S2pszsTKBhlxLDwzBmxT/QgTSLEOfeuaQFtLdC31MmInSDLUNfR
rp0dY0Qyx6xv+6/+/GGtbhOzwbFOv++nrOSOa67gt93qskWJi3OAIqWcZDT76qIi
WjMrf+ZLEd3SAMbwMwqq/kwVkGZZgtT7nbN4Lup2O1UtC/Pva0vmBxYKem+Vovr1
EV49Vrx0VzC+sepciDiMrgNYkhmw30g19s3ZcNXCnC/OBQQ/9HdmQoh7CaPIZT5U
SCqLAsMy5hHt2ZvsikTHXmKqjc+tUITEeoZ++oQC1j+nbSCmI7veBroeX5OPyNts
ElR2Jy3uhvj28NQ91Zr4gTYOssWZcp45fkOgYFNLBqiqP1eRvVlyslQM4DU0yS4y
8RYjf6MucOKrwpu8rhrAP4HRC7qorQZ3BOo9YICbIJ2FdciY3i9gYFFBDCHrRtyP
A6Dw/3LodSOZkLMImCo7JNGecblQfZyh1+GqoQmYj0fY5lI2C7LzDRD1ctFtHOd5
OwbLNG/QgfH0qT6F4GDcyRthc6vRUOJ236gSj+gp1LgCZA/0cLrIkB7ZBXiBOAS3
e2DS4hTmlj7f/R3CHq5KfCIpOkE2NxKIP10izNny5bFGL9Q/klxtmv6WIQgsPkcE
020obeQlCvMzePfWvyS/3C4gHLkHkKJ9WAmQlfNA8OnOo7rCdG4oaqd7HlJztsf4
3GM1I4PLJdXs+tFp4Sy6FoH0ywPY8GC6gFsueABZX1Cpl6LkZvzVLlxA5MdcG+Yn
TNrtrOFC4UtCNSJrQYfTGJxvvtIwfNN1nKf5UQgrs8DkUNBYeCg/qvfFmqsTUEIP
t0FE3AASE1Jm5W1qTuyxqrrqXfJsp9J/O6V1Ag3VjjjWaUNjMgavItCVAfN002rT
J6dBaGZcknSeS3dbINsbejmOQAcZ/BqvTKbuR9c7x08lhfKlO/UUOz4661ni3fJk
rY9epZaEGQY3HDDrChgJoOnXDVImZHwjTmt8WH1PyHvwxi9YvyyAJZC4wdzbkbif
tbtLFkLWmTROZoqg8gMgt3FRkIr4Lhty2yIF5L/7uQEJ7zwV6vLC11vDDTi7wEJX
sqeK712eSdvieZXYaZgDx6a9terbyjzP78DImafdzyBdxrruOhWXsgb2ydyL9lK7
Ds2deVXb8B34uujet+5wYfMyBQ5rwqfUP43uDj55JFnLG/Q2BkpzdlaVwMLNWl1v
xJg+8yDfnPbFDfT9iTAZEY3GuRBm4AB5NwSMmRYxBezazxK27rDqIitwL+tSA+s4
14OViOkxMko4r5SXbedDnnY6EtQK3T2gY2JVhWRycx2Fh7TbE0v0xIGtzvOVeQtu
LQJ7sYx2ZZFSv4d0ODQ1pAE6UBc5XYxqTQ5ZyahBek10TOFaJi9hTjGLqhYX+gqR
4W0o4Rtmxpk7YvsZ3qeaZTLBmfjZ3XhyNKYwEp9aK/iDg19VIi9MPnsPOe3EgHz3
huPpJ9MPFQM/ZncFBZTqpu0qvjytc9GGILU6iL4VZx42MgqovVmiXalI3AQnAqHZ
LPylaYfN99BpgDJiPeubBosFEkyVv8baJ/3UhvvseDFGV73NXna7Sl2HaVvxcZqT
wFMMstrUiuvMqDIFSYAjJHVxDBdIRQLKL4Nwo92c52CUd77VbzT67Y1UqCF08W2R
R5fIsr9VqG0YwyE7a+74vVO9So4LMaW2D11M/oZ7qtGa3ysgMt4KsBzrCz1YYpA3
hduPcRoO/kZYmiI9aHtnxz1/kHjAkmWh0R3msLicIj8oQ4PZ1UgjdE40uWIQ+lPw
OD62wmVsvKNGWSLr6KtDPZBo+lHCE4gAw2CnWg5kj4RrnTT8jwTRPQ1w/AxexrD5
4xDCZg6Xojj6IaIVkCyeh3RGA3CmUa+67gGyLdKd5aPnBkpuusCzGZnKGLOCWtpg
zaLLHXIeudst0u6CDP7JWP4i+tcsa4OIhr0VV7d6o9RcMAp8x6RyajbtqykSa5Hc
jBhAjvT+hLQelFRYRQ+CC44pwz40AhTauVvd5x+Sxo6fcaJencNztr5kRhS7RrbT
Q3hFldzEgv7ocwBsEonvpffKy9LJqJkI+o60tIJgaTmAaURsTm0WZpsrNBd2QHv+
YOvALTNyq7Q5su6PVgmKSNw4N7KwdnLjUJxNqcN3hQjRIhMk2/usWebUMNadsaPB
axG16cZGjIYQfAMJX0CxuGctEZDBByGH33FKTSteRejLiq5B2K2jSRpAsUj2W8SF
DQ0sOFYm7xNhfKzU38Qu40QTTuaqCx4G/ytazNWWKRhFCdHH4sTc7+/opea5/8IX
O1xFv9FWfnSsRJtaYiPdSXsY6U6e7Xjh9YfX/ejnURrA+wDfjs/mWMq1BrwChlx+
Hmd+j0PN3K/4aET9unGic2FWRAv4sUx/VGBb8SQZdt5KySOJ/eBqfy4b6oNaNnB2
qyqcjKpN5LrudVmvYdy/o79OgomyNcy5bwCKZ4HqjGeo4JkCTBwgeDbP4utDKh7w
U76yn3C56HPvrz3k2VgIsYW7MOTgYtFSy5tHlW//XDGOhlzNyUWd4NYM8BpVF7Kv
7V0YCtI8jIEZWDp54VypMKDW5NeF4a4/bDRs9mesbOFRWQr63sWPfNFhqe451hSU
C4KNYTwcD5gjgs5GaX8bsrcaKGnyFP4dxLYUor+rUJ7UIAo+ajXQkezo82rpsqkg
zXmerr1fgeIRIkfR3i/NFrrCyDnWhQ39BN7RfQ+R/eEHrQyuuIJ/SZMXL2jB7Sry
GIBJZVSHb1nUWrV/wbk85msew0lpANx+I8txptJYmZ8tDhKbNlJEzkEVUHqrs/Uo
Q/twf7DTl1kDRa32L4opGxBjNzNme4COz75fhrMqpJEZOHN9O5s1BPe5L+zgHPgi
PaMdAGEEY0VOAzbMdmzoXJDP7UWp6W8XAd4+hJz7k5f4TIhrD6n2AYES3+1Bk0ri
zP+q9ZD93/XXJ6zjk6m0sqkU8SZDdFruDIy9Zb5oBpVNTTxbCAm6SCCrzXF3j4SK
mVUYezj3KRaTEtCctC/mGYx6LuCJuzSpJMjbP6FlL2KkpGAjyu4N13wQ9ju2Pbfr
vb3QJga94sljdyhb/SQjMb0oso3LPll+it+rRCtarYW5UTUxE2AyWd3UCej37lSf
PFbpvEZ4SNFChSNUQe7/md08dFkah7pPm9FJCGTqyTUv5yRf7sxlQIliaFIkHGyj
8dYsjf4Rq6XQQ6EAuaKMsYMOwAyhtcdpmA8brf9sGkJgWbRoz9dUVRqkSBEC0djC
lR5xATGG9hM8KmqPxiQ8GH+U/TQoVwKO9bc0IIFmcdXcJvpBTeL9bFCNdGnYKvo3
EajwF4V8sr6YnXmpkfRES78tlH8Obx4acFvuxLLSOTLREK+DGBRjEQSuwkev8C+h
a9AmnOedNLI3/tYYhx2UPNFay36j1Y0dptweL+5c7fKK7EoMZ5Kkd4G8p4/uyOJ2
pYWSoTq2Lh0P+XQ0vwxIeAxdcIM0Ajg0z/byj6dMdpb0DBgttvxl8Lm/gWXX6Cqw
QqF4L7KTqf1zMb8cHfij3xOoKv0vOPLPJ+w41tniaizKg7qBNw7u//CjmpK8xCwC
X4h4n9U2Fs8PqD95BplBRiH5qlCCDFLUiOB5wraXH8gb/5h3V/0a2sWAW8RQmYSa
iuHSnWcTlKkf94IzR+Wblr8Yp7pybomu7vRRMZ3on4eFgDjyBowQ9DfIlbLqUl2/
8kkb4FxCAhxsqAqriHuUaMqzzlvW+lR97gaE7xEMuwt/7Zt/DUoPAP2I4wPA54Ib
G+CCoLy4INTwZJ9V+Cx+AM5FzG84dIjIvZIHILVwyd6VDOsRmqNOx93+a7EdiG/4
D3VopVwBKeJKBFpr8IGHJOxWE4TyEIl9n3Yk/n+BzTq6AP5UUnG3F9s6ay8WLgsG
IvmUvaPZhTN1TL/0UUtlhmBnB8emvTaw7Qtz8bLK4THowuj2no4LOU8gect8PWx6
mEWMuPoFH+r484C/1SrU3kij91MhrlnL+e2xcMMGQMYgFIc+FR1sZtXlq8gBXi28
ukUmQYKrLRUW12IInaxBBfuoNmVfai2RmDIBzLJHXMre4s3MQ8IS2FtQg1/Zaw9U
6D7qetWKw2f+oQ3vMqa/avmk/5FnI/lWb/6vlCKqRSbZFKxzajmWrer1c8AlPGoP
Wiyj+qUf8otmALW/+21lGqawWSqyrwPnw9j53wYxQoxEThG/UAasgpbrWBhwuXa5
y2F8GX0g8PU+Sjgut4cczHBgHw2+3K4JcheJ5gqO3JXd9L491jsHmG0CFr5Qs3N3
1Wca5mYZp+7SwniyuMrcC599kUsbmxyNoY7gzSMeEA3g/7FtunYqfYCxsCUrkdtR
JVmD0b1n5c94hACS8l7gYkAYvHApFcozfIxZnygri3jKtXtCC5qbY7zMcB8dONM0
IINtdudjnvd7TvWpOkSSA7f7Niicr92JeXJA5/GLIg9M0vLZl06VvLct/w0su2aE
IUuxLKDzst7T+XdQTb5ma9vVjijkaxRZ/dfKLL0cbHHcZLENOjPpTy6TL0suJmQw
Vf1bfKlcC/sfRMPQzbU+xEpnFbHr4IFq2WhSyEOhXZIABV7ZOfr4b1Xi966zL4VX
VDvUa+ZSCMbG6w+W/B09mmtzGqtK8sP1VyThxZPpjsUHSJYfk5nUR28Qx6UrR+C3
iAp/AeugXsMNfWocZgVW61m7JXeAkKmgSuIViIrBzkIpWhPuC0URQK7974AjqG4M
KOdX3uLWIkNz0ZGNdHNITEH50anRnUxewjATUdBGaugP+qzSN8EM9vxSlHTfI93S
0Q8DaN2tM/kdKe/3kuSmhzUu6LqIxKzRhCnihnPyqAOwI2kthy/3BHRUac++aWAP
GlyuF35xvERj7wPnu3Tc30/3LCCFpFVznz0azr8eDw5OnoYH8zvgGL5odspnwaDp
/UvRlvtnYYw04wX58qq5idzQKjxiQGBQWa05O2YzxoH0jmsRSBMWeF4S7dMEXB2Q
vXRwJ/lhCf3038h9J+/aDtHKNTqpxe4GMz7jrONsIiac8lpDAl8J6JgUJH60yZyX
2u6x6sYGOMzhQFN1/VtMhDS9ABlBpJ9FNB0bEc2ALC1wjO3kYWJ3XyHggXzBlyRm
PrgeqtwCf0yz95qPKpy6CW5JmnSHJFah3gx345HfB7fP5Vz4OIQhy1EpPtvlgtfH
5+N3xlpcwzXixqaEPBXgb1P1e78sUzzs+H7/p6eP+DZNfBCsE6r71xol2LYA8mfm
t6W9cbbwmlJ8qh/nFDATzSe5fuWJzr9xzSU3owGZBUNLy9Q4u11KLVxHNl6WNi6G
dus/IhpGNCyTdgC8D51Am76GdWTJUupZh16cRoYl9LgTPqeD4oeRemRgdAdfp4b7
j5HO3V8sLc/tftuo0Ei9ICD4n4nAKtlYY+Yo39eGmBEGHT/g8mMWPs5CtEWPntpF
UdNLxd4jGgFJ4BgJHUg6v7SpR42ogrAs3GPJ993gjXJeCkuKmhiggEbYEC3GPE/S
pTQBc2grex4X69rsnTMdUSIkQ+qEPjBurg12nyisbC/jLqE79ke8Nd2AyKrzZKJ5
ei8EuUfuLHZjUDdch8INGHpQr3ZKKScXSL7n/+bHSDD3TtKSLXjllYSt2OWPyhQ4
+gkLncfqwcCzRrBGkktH8rL2FqncsU4TWwQTSedYow4BY0SaKmuzfrQqhqYzIAOp
HIrR+ZfDBa+Y+4qEf2HV5ejzhtPTo2l/Qddlsekb53p0p+XBTwYk6HVGolZcisUj
dL5yS+7/IzF6IBobbAPNaUwe4x5Valpr4gzDVOXpl9K7v3XEtnpi/HBked1CP9wH
V2OLB8cksnLogsFgmMH37ZtUeGv0rwqeUTeTBiKLdEzULtO8/iB5kxuhzxQoGX3G
LrOBDwOA/k5P10hG3Ek9WRai8OTBIdocAaXQ8aLLuurt3Kxg04VAHvdpRuYGQ3xW
UCNY+ywcrpaWraAeE1SxaZvxsOPl02yVnSz8fl6HDLgLbtPBqkQ7+Y7hzjcrWxOz
I3rnwJsxVx6lLtvUqQejyO1R9YuBPfmREKqG+VEWf0ny1aOvEJD5x0JMldK9pzyr
W2BqOXnGj/bvDfNSZfZvqeOPSBx92DYDx1LBz3GZQeXqC+l2IcVWzaG9IOSI5K3A
T89AiYdJQm8q83krz7kaGjXJeM1tqdahyIvMR0BGuhdzJSMmEjPPaM3InpkwCNOM
O1j9TqFKr4eYB0Pi3xnGZk2T98byZL+KDQo1Youmo1J4WeAYfvshje194KE7BA7W
oW0oHzgCWNF3EE2Bq75ae/ta2FqKe2nId0ar+9ntS0oCmt6ogJzU1RtRvKwOrNy5
c33kfEzJ1VvaNdL/L3zkZ7FKi/pW77JOOMe/EU8087oYLd4NoYVv2GSMYyStSaOb
Kxdgj2xRifgvxriopOVMzGh4An66MrJu3a0jq8rDbksXio8A+jAfhrk1MdGPXqxv
9h+xHXcuNkc2dAI/BQ/oI50Z/bjq63NZdcUdSVpFb3h4lYdhYnI424QZVGRQqcJZ
DIJpIJRI4LoPfjC5ZTCvaE9BtvelE8vnWpCoW1Ld+zBF5cAW3q9z0Qvfb28xsyiL
kpWqenCqfPlNPTBt2uaswmUUVYuCzXJf2BrqburO7VwCiHZnO8JyqHc9Ib/1pEmd
ttryP5K56PhNR6sS6tTtEr+xt1ItjgdgRxoz0tdGbKK0pIbyWLGUoJTLEFTRMZ9c
m5Mop8LPHBnLWh/F9vcbSIiBIwc+93lTyIBRvEquuWnnd35mMwlzt4p9HqXfjkMv
IqC51vTE+nh3wPs4aDBlEqvqeNjcMerHb02WRMHL2UDTAkpet6J4DgtffgkOuzPH
MeMFvb491WwtZUXYNi5oGNRbAjkZneDTQSvJoRIMuHoJbAUVYSHCw9Y21Ff9ngET
MpX8WBzmADDKXqVh6iwjjAp/4F/dttMwQ0fx0fPeUHqOi5qK2CYP08ZzpS4yExsn
68mS2RBvk5YSiz2SJTH8ETkVoJMsKtYokGwZk761EssGfoaCktygbxNS+2Vz0Ryc
8Js+2n9LJcY9lRB37UuIcBnMlCvF2ImHB4BQ7q+/LuPDGBM6y4luQikMb64ZcM+J
fskIKqpQvAgpQi8zVTTb2gdYyxNU4wLbh1pFCMJclB0d4b3QlgX5OME4BkegnYTx
zhYRdZoUY/mZrOKfFKJfazFF+PqOH7noxIvhiVRm8LBWO5sB+nxhkMB2V0jynSSy
9zAv2ksWY9Xe7yHIp+MVQsMjpup8heardBl9jaUhQSMtJRjc7J+hlFosJ3hVHhNl
eIKmrqRtqxRf6YpT4OXzvh2kWjUz8dR/pGSwsoA0pYO8+ZWQ2ltkExneplzQ0WpI
9uYT7xe9ajtAOBZT7/9Jtv9mIJojNP5UeN5zWKhDwcmtXqnxybwxqqJdsI47jxoB
orOhUOX8L9+8esl2WKwOC6+9B9qVlgW1WUCxdWy5EH2clX+dHsNCFoLntQMzB7CY
Zu3kiWW013f+n9kJd9Yp27miSwEeIyVyYMiNNoGNVnWFkvfqvDeyi5O5sWgosjc9
X0sV3CZFGM4ptCkiqfUDTFSTGnjUPhGGtZayj4XEHAoH0cHD5uGG2tiN2qPxL5ip
yo8sJ0zj6BXhDuzcfzgi3g0v4qXCj+RZ6CpsqMmPWwS3kmlTNOyT3PhvZdHyZ9+n
fxi4QgyteytM4pKDq6ifCm3MguQ+VqkW8PTwtXafuDjoonNxIEyxSMruuDdq1Kur
1IEc7PvliCExDHSXDCvPNqLz3f9yoo7pLrh9u7IBKvaoKUG9KcX7j3VfJqwXaxQ8
WgRpKVA7vL3GEtCr0exrdt5RtmfulMTtn4tvmBTyF1sAktmuWKziVYLPZxfaEJ9u
QUd4Hy0f8UIOdp4GUyH5VOuE82/Nrw86tCSs3WhuIPgC/Tg/Bs1IAyz59ky5hfBm
2t5IGjVhDjNefvt03M2Pplwr1c0rKVFPGl/tlyrZzXJnQazbB619mofOnzmcIZdk
7KB1+UTYLpWb91LTJjYVju/Hqf/V+hytJhFewfugO4DD8mKuXxaCcDkYVA7KVJFb
lAMWdz2N5XTHf31ahcp0e/W/qRoI6uYx9xZsttNS0JxZQwUuLmL1Lv6VBdVM3+cO
9RSend2mm6m+HPKdVsBfEUAo/Yzhi5H0X4J2S/x0XQEMyHdYqDJaZc9qj5cjywPK
TkqhBf7emCY9WXMBZ8rFBmnvWy1ImkYiTlXqDH6fqlMMzER0Tk72T4n8MeIxSYp/
6PzBP+KnM41yB0+E5+QBr7v8ctgo+C7WYJNQmF1PJ5q49oQbqCluuqP/1JslGYxI
RxvpChWi8ZgZ35RDO54ksw8sLIT8jI7o4/ksF5iId8nikJ8nJWkI75obfxuH8U61
C4SiJXDwdVgbMt0HBjdhVqX567EUVtw2TzQI4Be3PUy53N8U60OTSS5roEPt/BD2
kSjEyTLaZCgSDYMNDAOJKSvpf9ZspbEP96zsxTBRnApJwEqU4d0cDsoxUsfhSVRq
biLrJcs4BTMkW0sldFWyLtOeZlGCdJXa/gHliKMCHNJXXr46YPj69uJKRzbSFd/a
zb2C8l1TVmFVfunD9EDRd9TF24JqdObynhLs2FgYKRxNwc/h+ddlwrSHRZKC44YM
5vYCJqZQuYkb6fRjF4fH+l6Arl949p7syyBee/enyXUFYmn5wrqAJkxHZjIAuvp2
49qpwIeKasc9tm8ux8bJYwnNbjSBZxpvLeNpiuVO5Rsep+lXknf9vR830hLUR7OL
81GGlEBSnnqzyEQibXB45teQq2413i8aJLReD09cHW9d2lNgq5lHzZpS6wf7tfhf
JF++upZ0jixo2WHGdp1Ns40jiK8/M5BRowuMN4wLveQpnqk+HC27BR/IjqT/+FCs
MNK0wUOblSROYET3BFZkoDJpgeNmjFI+wjfQPipkFFb9IUqhLjIzG7mdbaPRcc2F
2N48i/UyddFSRaICqs4aXU5bUTLvM7R1nxIVyvlYq/OvaIV3wg9qKB5LdrQM3zsn
vNkyyx28mhutHVPrieTWnlMiOJmxyCa18oNv4P1o2sccKNY7BW6wWAdzUO/Cl92Q
lqepG+scJtnFDYFZcy3HhNWBQiA8xBh7QE/rR5ODvtjkskJHdBuFfLnd7YlBoC54
PfNCutg47QJ5x2eRHG+K0K/tDqc6FfBXyknElpwY+NMWHjBxdSXh0xaxWfpfqxnN
VPervOz/R4JvJ7YP8TjhFPhLR1GHdhGQEsko2ia5P8eLXu3ZzxZ6SrBRvsm1MUie
RxDnT2llSfNzgb/2NKh7SzUfZGhKzV9eXMQDU7Cr5fETZfMO+WUSmCUsPDIme/nR
X4+opciVd2NX0c8DI5OVNT+P7uj1Y6KoEXgrgapTO5lDmWOYLuEr9H7em7g8ghOO
cR7WUfyG68T1auVvsJ/p4GIDKWqGqxlAzmO64aBjEcq8LDVsIcGBaiIoi9qPhgXj
GniyPq0EduBcQKpWAPopWniZXE4yBrjiHlJKBZqQTH1r7VVV2/GD4mzSW72vW5ri
vv4wMCSEuYmX3jNhZ80VIwYJv5owksNPQsLjWNe+yZBOKN7C7gfQRjzj78ZAV8Wz
tJuhVK8cte1N4G5lNgBFW3cAs3gQaUuVlX4AcMe+hXMKRUWXeMGmffhgXrOeQWZg
ktqiZfXY2IFJpgHB0ejx2g37wYrKOGoDjAVBHEx6SaPeAh9PHPBF2Idf3hp+TBUq
xTq5wza/Rgje+jMSYfCEUKwNfzYUMCVJI0qASB/WPz2jsSSFls64wZiLAPlnMT7T
E7J1LSD/XDz0/Z8AcIunpyk6tYYM4UF+uRVMmD5czOSYbTqoLR2CY237zRHaZTRK
wkWduq6+KMocnqkB0CIFWcvyITKUuKGRcCz4xYB+5Z9sV+vifjVrnyQQ0K0bWPC6
JBbQmbE2du/+pclpanGYjFsubQdxfIX4spXl3Ik04CkAUL8Se75cqT51SlsZ4/1w
toC6tb7EXNRvnNgRmnUBpRDoX0Z3oHqYyaTqrGYzq6eJnhDjB6CQ1YX30fumlBvR
Yn5ghnc654z+8cn6cttUGH8IlU2O16om0Gg60VM4ah+kHPcWWa8wa0bdJV6RlHRm
lucrQM8WVM5OJzoXxzMIsH/HvKzXEtQzCpTk8rxv5lv0MsPjf+ya5mBA45DcACMI
0WKmtEUPJZczktxIxCntjdrLIXfjRDeeh4/detjCVwKjs2aJpc+tab0nXM7iKUre
JHrh6dSkCemZhsB2U39+ji9s/Agfk9QDnjIjal2n9kvYDdhp0YsZaNIzF5sf6qHK
7woY9BRq+UZedVrPzEhozjnzoiXhd+gaWmwCJC4b4RT8LtwLARcWCGLDu2VxUlj0
NvL+7J5hPJ9r0lPyyJ+o2XJTPYhnFNcLGcqOHcVAqNaqR5B3Q0zXo7ORkkySpiwT
8AbfaT9XPK5B3epUJcBMz4YdIv/lHIycHf1dhFp3/9tSP63mAgXUAuRzZXRG1QFY
v54RhrTygHQBJ7UFvsHQ1b1Xqr4z3nY7ogtb/9pcCmOWDES1iXV4oGJ2K+9oLeET
y+Sehemvbyy9MpCocw+79PUQVn+mluZkUzSaio2AyEDJrwwtNaNf39UInKAt+R7a
GdjCusrS3E2p3euIR/2pAvhE5NVr2Rkk/dlx2AtkVwGl4DQDL7eFWX5qv1gVXV2s
NDbu7jFgdRapMxtUev+yhFx0B+eirndevfM5YZntUensVifqJ6XLi3l7sE6idJbl
sh96561qxTD+hChmmrNMtzJBmnxDsboDHKkeqCxcdqGnkBY/YTBw6vKcVAj+qsmO
gcWfAtqwBnX9YZunVtQa+0ndPzHSUbUNgea+FNxT206Z+PTO3tBDjFjhwOJHJJOY
YZNnFqJtYp5SLfG3V0W9V1N2cjPR7EYP9bA6VMg9Kv824EQVgIaeeGZ4YQBLbb5m
vkQI0aWdaex+8vF8aFk+yA6AichIpSkrrTOcQfGobVevYDYoz/YnT/hcMCanipbs
0IRnHoPGWb0eOEnmEWcCLYCbkDn+q59ct/D4OjAMJ2KBoMFpDmcSNOZv8QyOby6j
Ps5MCEwnKj0SFxsp8BAx9ZmeYY4uEzr2SshR9vGU70WwY7NYQNeY/Vxp9KC+anBA
p+233qfERksPN/l/q1cRVWrBGn+ltahMVFMgBofIT8KnwpJAr8a3YnvA/Krrh7Mc
et9dyMpwiNUmjJGkkBAOARzawk490DdbmfeGTLWQhJuudmyFvNCSu9Mb/yd8NymU
EMLclSyOSOu4G0HmP62AHy0F5B5AX34V3G8ub4wIoDm69Ozsz4Hq/wp2iMjHaxec
E/F+/vyI/3UNgqOy6BSxKmiPhhaWkt4xKSywRdvYAMRZVltdrhaZtutBqJETq1FJ
B+J+K3DA0A/ap8UIK8D24r30suc18Lj8PcPOOlXfYtCRxO7YWvGCyrZ0tfEq1cJ8
WEBti0jkEb9SLVcbo0oUPQObajuKCp88QF/qZkoiCFlpG8sdkwVXzEs8V4Ve6HKq
yV1Zkba4mVLVj/HuZB2up0hfZmveMLxFWuWf4LsyDeTtp+NbxeD7OJWOlDob4dox
Tc56zmsIqjlwFmb0+H+qVKk6fcYCPmAOe9e+KbX2Hzd4fbzLHJghVEghb5ucuoqH
iwzxKwbHqm7bswbXeClJMMEsRv+O6dqYtzhckSSAT1A1eZii+1F0xcnl1j/xG+BW
wVC9KKdHYT0WJdrCPyBXLwhulz+wwofECgm8N9X15qs50B54zh5sXnjRIFYe+1Yb
scsoeTThbRJkACS5OLsM/jzVMOU4hXndT26wL6zcu2ICKSBN9bMTaC7aprYXzOtG
yZdIRCUfvuekMNDnPu1KB8V6AxpTxiJ6QRPSVh7kJmkQB9KtLG0Zp2B+NtPyg7hP
F8y97jRsvuzsR3ZcNyt1IouC7A18l2ORgbW46nAAa2/54/gC76ZQT3nbCW/yyK/y
qcfSs9dSFXySdhHBaBrh0lJFw549gBxCztnTb0PkADWA0CkZABKvK+R7ok04Y94u
KohKKdk8lU1xjmoT/K2nP8ZvHj73DciT7HNMRTxZ3PzXwR3P/m/rvuMvB1a5ZBZh
mojY7MG+CZA8L0Vra5W5vU10KjzGM+DQnFIfjEkk1KcoiLWp2xTKu3/paEXjfXGY
5j2Lg0h3oT3qyVHspQELSyE+CdNwXwEoP2BENHrMFBHczWlXalTqQzDZoqQH2RtN
LOnauTgCwbUc1EV3bFkyVD+EE0y/nxsHvcXyhqyOHPHErDG0hWXHSBLCx+QrIgZM
EDuoSJYLe68ZMLai+4O0af6Vjbe3eIw9FOI/uPniOnPl1geHfQrANZHqAnngHeZU
QjUmCfctOfk5N9NV+wgHnCJhOGSMJnY2gXWo2+DH7vKNBpC4ID71ERVB2rZ+IOX+
ZchAjyX0S8iw2q53qKCRUVyEvXjks4e//7fZuTozc9R/idAIWPXJuZrZh317MccH
9r4clQ9WKOPzBWGLI45HfDuc4iFsty2ZwIuj2cmRGdP8YycSPVpNDS8B9+9GdJr2
OL1dhxxx2NZIK2cmTTbX1VQzXSbUkl5YLHO4tHU6Cqk/Q/+ijRZm9jH0f/dm3NI6
u5DKCB2+cy5D52Uz/rUvTxLmf06LT3ub8smSojqN9bYzr/XNo4TvxY3FeBwHiEzX
D2vqglLPHDzDdhTnb3Jt3PWFFwoE4iKVC5c6fz36GCcoYpMIDvgwLLFKm4Yu52Hh
mrRSGHvX1kuNw/kCc1LFrg+Zbr6VJy3LFsCaLi3cCBEK/Xw1sMVQ0I4VmOqg345/
tZfYJp93uRGz3Osu6ecRT5EiFI+YwPgOmYrzS0ahJOMSAYD6rQXesWhAUpQwKzHu
2lNxOCsprJAgB2Lfq01wR9XE0+yjGJMHOnkl/Z8q1VydeZHcjpGUIXqOgdRGaaY4
si00OZiz+2+YDTZG7Fr18hW8NCYbA4TqoasITaOyDk+6T3QXA4AqXyduRfhbOtUy
kHvqYGtFYDFdIuD1lyT3hxZkBjxNa95dKEiLgnXn4Qz2QXkL7pWv7wzwtUSkT4uI
1szMam0/I3jvijbaQiP9IOYfWgv0olmYNyzBZdmrbHqCeJmpaPVceAbegBG6eANP
b/YbVFMJgqRUkQZRDl6wbmxDCx6VNUmlIRfTToTcx44jCBWuaaZRSnl5tKGl6SoH
/KZokLLLkxyz2DWUq0SwfDEWowFy/OYmrPIrDnOl2Rz/v9dshgXDvH86MZdJnMZk
Tovi8RoUx9lnsX/fMq9Hh4WejJ6VHZhg66jJqx6JvFjgUwqfflbbI55Tzeu6TH09
AHOd588CRQQjdSmsgG9Y8uB5e1mlw476yzd8S2mFG+NZebHxcmXY5529N4jfHUB9
aAoctC5Jo7RXcCXKymd2tgjIxDbTsGxuvJXGO9uIm9YC31+hT4N9iq2aH/L5YZ6M
TXn+JOmxQSTubslEWn7ocC8f4bpgdbk1svGC1PTP1cHodRSPBEeDW28QHy936frP
UsY//SK5h6qzuv/5lhjLIf+hCJjROWFELt3PcLZQZ2qgstKI2KgH1nrrq3dEIwn3
baUl9XyMH5L50KVgoaiPkG46WcXQoHSz8SvZ/breGwuiZ6y50wTJ95NIM3fwAZjY
sl8DTT0bL7tqvVUZ8fEwHWaVw0Y7UtNQXSGbD8zY6SY3YLvWKI4O3R9C75f1Bt7i
kwyFb1Na33QDOKpYksiVnIfYqqMLJmqrb0mCwSstbeBEwsco2iRPBgt1c+3v5HGH
XbY8zma6nFLTxemGrTlQApdc8Cfxsi7HtUgTBMtpVVOAz4q0LqYuXWx3XR/95ITP
anSpK3t9MAR0MJL8GGXfRMBS0SPpqzivjxVp7fi6QTz3/hTix4LP/GoFi93VOIUQ
xtyUjUbztVm9Wyt9+Q3HgaL4ZECF0lEoeQlvp1ZxoRJfnYoR4IkCYmlpTyHle0K7
dphvyrj8RNBmRuI7Prh+srikhJOYDbKF95AjMfX8y1w3LqgLE2/qAFfgvvd4Bjx3
whcdocRRfACmCFcyu4L9P77RCN3JarMn2gfv+GqReQO138m/q/e+2VLx2HSDoj6g
rZVyF6FAUXBY1+aBBxsXU1MwCzT88pCUAEDwYy40KHqHIR9/0VnLXJqtuzSnpke+
5EZPh+jpwSwL9lbbk0dlJomn6RRLPvUA8i5uU48uDDANvypdPedtApKePxEX21sJ
Rk9+9hg0iqO2C8chK8JccpEQGu5JfFJfSaJuUO2vwrqqnJLsewhwrmx8KoWm2GIA
Gk00cAITpssK9I/gTB+0UNexAYa2BNrrOR8gQLd9Py3Fvnb6gru0GSOPCcZWG8s0
UBCkHLQq7F56BiEHZ9YSRIWt1gPGM8M8kf+1sves5QIT3GPUr14+f+WefogfaOje
PWBhheTeGeycX3H1iuiG3lz5HzxaflJaQG8NiazXwWv9kWsdlPkoyf9B5RscUWGz
E8huysroWX5vjuI9tFp3sGVpyVlLvFgmgvgCQ3cKYXhe+eBu95XlWchKyG/gsPap
tyC7gIBrtCsv5GVD+xyfgdtA4M33ARI34sLhxwZmrdpgrpKl+vLLaRqsGSCVIKE7
tavGmpT5/bXXheJruHC2jdO9Kmhd6elzME07DrtEj9odvwhE1UosABXGgDL8V8qQ
tJqUz77MfsyTe2y2zMULAUG4uzoQBSXDxHON16+QCnqgPLB0YPpNUTdEl+t7wRx/
VkDgJVNycB2WQQxJfxFwMJ2PpDXDNQAlm7WxB1G9swdVjd4vYImvNLXrI6xcrTnX
TWSxK0JbS2w7RDFziigxldceaZ6+rrQ/B/L24GVPGg19iJjzxCNSRgrFLFPZ9Pzp
7A6mbKZI82xpV4n/R3JEkE83U//HohBcnxk+sg6ozjdscFKlo6uDWi0wfopDXLnM
iVV810WXDjUuKc2Dm+sLttGRw4UmQbnxFlmYFMenKUof9QUCbwSw0UW0VvRw7WW0
dt15OCdPVip1qkceP92qOfzoYWoUN6o+EEhbTisiOU54ZFdfb9hqOfoXSC+8Dl9W
n2zQagSqk6fMkLLydmKBeOYBM9MLF8LPHobn1ekeWMAk6v6y5BRm5LRBuiIiI9Hn
edtEU+MF4LpcgFkTjc7dfSdhWKyjoeh+hRj2rHb4h7CYMZNT5ctKHUV0Uao8GxiN
hA1sFIPN5tC/whuURcV/BfnBqaEbcAaFEO9Dig9w46w2xw8yx0bDarPY4Xg06Rv8
anLk1vI3QI6eqUHQAwDLD7znFXcUm9jlWLYg0L+rzImBd1GJgeMAyhjInKMa+zrj
XCHO0SUVF9ktS7X+XyyJIAhkH+D4vGjDKiEck/eV/hcChdQOfyRbTsFPZ+0dYeP/
G6RUMRcyvJ1/eacHCsKWr5iXjJzaqoMiVrbAFdd61JT4bpDRMD3ccv83BStiwfow
ZLqy6NPlrA9ZeA9IVh6mw7hYD/B0GIlCeiIJQGl/iaIFVsToW7Zyz5Im88pR2r4p
cTD1a+Z0saEpkcpG9kMHl7AZwhdW38Ysn9gsWTTAUm0eEVZJ570SA5DC9KOrgPsw
wTTD6JPqDLXJ49R96mqVAqtrs4/738rcfh20fGHE1v9VL7Gma29oTZH5aFbycTBP
if72hbdFgVgksfJqVdXq7AFTPv/V6J5UDySMr7aPBD9NM58xrNwFnmPJnfMZuXBt
vwBVPRxetWZ27t3/fLTSNjSmubEgJQNKcSS+cGK0x9rEqWpinRjQYLSAl0uTvuLs
ORjuSnd6IPZU78NWtRasto63b8zKJMXGThRkQtrqSvh7BA/VZ/g1XIAnVbSZJp3Z
4OEr4CM5BcFPDh4W/em97vvQBIPRtmfcMWOG8PRxiWnXQyrYGNsL4lePyb/NatQG
JM2U5VXvjOcE+X4Zw3PQU7Cz+/fkaQ8HszzbonWR6QX1O1o6PeUW5WXSsB6O/vDJ
wROu8f2lbXhQBogdDrwwS3A0+p8ckbuRXHayqf2jfAia9H62K/T8ONsotA9/ABGP
Bz+ILYQWcIp9Fu+EgbiBXHe/eZs62uR3cFJNHii2Okpb+2g4klnCMjpt+CnQ66d5
FnwXZjf7nN9nbgWVmUkV+2jCDYzHDtyqSb29pgA2IKgtPlyJh9i9RNejjI6he2NQ
mwLlA5YB8JMnfvKKMLWEBKf95ROtNQLv3gc1msNw5zPlhW9Eo/1wy0H+Zcfg8KvA
gTcYtMBc7zP3UCul+jT40ZvJXo5cFUUb//qlyKd8Q29ZHJDwMoO4Fy7MedjH6zcm
TwjwL/sGrcoG5lDNAgkvr53bC3O268ryF4CyKJ5TQTRkteJhywZj1Ux+LlpVsPZZ
skDuOoKR1CJNrh9knsYkz7pOV2lixNWxfugDdEuwetHI/5/hZhutwO3T6QqOLZuw
+fkT9A/3cWkCvu1WOm20zFA9bzn3n11e/aUhhwCc6dtuvIqd60hzwo01O7TwNU2C
OXy4Y1nlvJ2VGwUZXukGtMxbOrOtmHHX7UxUMHcIPRF4qCpBeiKbbCmyYxIq3iUr
BBXE72gWil7Xai9x7CWXg9rjj9wzpHPLul5+sTHNuxyp3gjWRWYXNlE4n3G193z6
icm/BKN/2m6xAWtfB/oB9hSK6UtPCzsOA7ASnX/+QZftV85GiNCqSl3Qb13VJY0U
refvZ/DBxvEkqpb5Ib17SpwWNH2ke9grUPsWKg46fhfVGzl6uoJor0ZMCfNxvED7
HZ8rKGCa6bENElNepnsCEh5YZ70RcTnpRqefWPM++YZQQsY0vcXc0JbLCe1srW3R
oYUKypOHmCLczpOtbceDNQq60sUH1KiYJyCSm+X01VoUMgtuCfzFx2rUI1XmLfJi
qdH8qBiUlY5ieZrLALPEVsi10To422oWwX1NhMuCuSxVb35zC9FQyWRu+k9zkDeu
sY98DbOCM0QSmhfv7K7Pvzq3afLl0GgWcQ1fWLkwKR7R0nF2hxwNvYN93fz9xt9v
nKiD2Pu05+F4Dvugeg2urdfc5wnfphcM5g1gC9cfSq7NgAEjse4L9AZq/rEcXYo8
D4NkXTPTKCdRCwesj2E5+gUNXJySOfRVuIYzjgwPceDpuaDPhaxbJpU4VgVvg+EG
qkKkPcCEOUdkPBRi3B/FEKNQcveuIWgFmB7WIPM7DB6lFVVhREHHhSSB0mAcq0B1
10M2+S8KS/lm8uulrdVU7yebasGuDXodgJnXSkkOy065fMNjQtclN0IUmqKPatEb
C+27j75qZABsxuHAitQyHpqQtmD3QqEwM9G/EiJadYXcD68cKnvnBQvZ6FfcQp7I
N4I8twwNcTK5NspUJKPM8mA9jPDvAsG9MLkpZBh+j9q+6PKqBEIX5gsA7PTedkYu
fPg/s3gznJ5i0SCGeJoqbQ2M3H2/LORhZ3XqRMK2tOnaLTEgZLQ1qyJa3xlHKlUo
gJoFsWNmWJs0qXyLk8VvipFH7otZzjA33VbPcdO0oL6Xy4CFlxmWZDJuJCLG8JF4
5kiPNdoJaPnaYDb5lAqJz8yBNJskaoIQYrAfbmoo97DgvXjKAj6WoqPqVwya23mo
C2MpnWWHltpatYt388srNm/Yt2SCrFcs1FH+cVM5O144Ateld5cmlL+n249ouSr9
tHGmtuXYDb99jsCXDDMlwE8Su0FN8JoY+swtIy4qbimCdC2axtyEBnujPOwajgzt
qNrqs86g3i7ClgDh5swxOI0VzIp5orlbTvPVCVKvI45Dhx+AhsXK7MSlQ7yBl8fs
MYOQlbO0y/y/IbYLhDsbQSbnCAKR1tRETg2TY8KPyz7a87l7YmpOz6S1U/IalWy/
9p413o8Rh7lO8U88vr7QMqsVF66O7fPSwvLQ9t3owlAwJhcnkpak9/QKra/olmbP
GMkwLIJ2FgpZT6YlGmQh8nov93NoNFHwFROCJnsG7v/WVGLR7dtR5SpMMvlmzdDK
EOl5zJiyJGQMB1yO+qMQecxD2KRTwrBgAb7haU5wrGm+K88wLJf8UhOgvapto3xl
rEAF47+5NoZvxEE+CfBUSu82W2ki9NHvymP1mbsHvsmORI//XK0txQoQC1EHmsah
lSuXjxSHYxG1XO2FoNxADcU7gbX/PqdH84lzUombec4ZaVzpPJD51xlq8Pms1+LB
kylHQkjCrYamGdRllI3bzIiknRv4X7Gt+fS4urIsHoGar1vfqWE2UmyZ3BSGkjdF
44vj+xKhwXYv15MoSxjkw3N3Atnn9MTMPMveZ302WKJ6fd7mklaBheDoUPAJbJ7U
ZX9JIxL+HvPkP0mA3q/zz5CPZScKc6Kwv5+xQgaT0ZPCzDAlMv6uKxfgPL3MB0Z2
tlPAOFbDXDPaoMHmrUVBVfzs4Pg28zE13NqRlXDc3Cu2DC4ovncG5VMIqGsScq57
0Fq/L3UNdmIF50N0vjUVZj/R92ExknZo4jQzvWspweuGJOxvGz8AyB4N8sLv1WrZ
4QcGdW3lV5ObGxr2SqqU+2T5m74Mr3RPGjKAYGY6bzGXNpjTKr+QdpAms5ZhwFS5
nT9h8L+t87L+wsxE09cODXY6eKCERwPGDlnQBgV9hNzIP6uxcSJrvqEOnhbPWrCQ
wq8vzuKHyFazo7VMkan3f14ja2SxJPH9u+xqIPGah0VvODggZkKZ4/rndAjGMxxJ
hlMks84AP8aj85PGTaV1bl16/PQyxa9KKt/2sJblNifdFEFTbivAOkkRMfKpF4yX
tNhx0rR/03cEdYo0uX9aPlKDwH2SAP6gJdjlI8/l1nQuFUxzPq/BBHNev24gP56t
8yQR7fsLxlTzdcc25tdUgSbbx98komXQ9Xrt5Yg8thCnak5QEMy9rc2+/Y4/WuJf
PYta8ZhJ3UnKUeqbFdk3MCLhCa4+K1ZLbucoSddJkOipIL9FRiC7GvxQ07MpWLnR
U8S73Urn5sNfmaNTVh0NCDnAgISZnNb9eRB7yyO/WeGg3LJR5el3towM9zQJCX4w
nsfNFtETPDpsg42tuPrNT20V/l2XdkxiZuCVfhFSHiheX6oh1pv1SdJOEYHQQ9xX
dtXkBTCXVXq1FGloU1wOMtEMqOfqZcUfQVjQnZ13oi+ly7w5BA7tkNsLC6cdkkRM
E6y8qdkrG4P1fnUmU7ICioVY7bv57Fp14YG8iEQRZ/ij5wHy+CDsgo8pL7X1xiLr
A9h6zmQO+TghUqHdSo5+VU99Oekle7vSBWH8o5dutKcSCQIoISQF68WVWWYqFJsD
1nmyaVygcHOWT3IcCZi7mvh77zLakp+VyuI5JKlpcsFC3xNJHj76yRI9ytxXh/Y8
BX6TktOwHCyF4oBULhSIVV3r3hLpBqAYb+DWDVEJJZ3RVISztUL85URackx11W0T
aqonKvYWYWnRva0mEhhBsQNY/qJG5t8/xOdzMZ19mnlYgos9D6HhMuFYZvh2bLCp
7UJIWj+HmPRdyejSFrXRKz/Bh3TJtVFAc1EOvJV1rM8izsMvoiDBijUcCF3Y0X+U
80CfxICcFYtoJ9LaOTz+Qjk3LFukofkGtLCSkAGILk7YMhWsQ/zD4O2kXMcwP1ne
XrrMOhtnwjuXZlse3ofWD2n30uJg48T6mUPInfjCywAJ55bEQC4/1JFaH7vQyem4
XJGxM7cKmfVuh40rLm4N4HvRO9Kz34gW25aqNIbkX8HuTurv6MhuWK5LZXYI79iI
ebKAMNCjh7si/lDpW43NdIzBvb+2NdWl5R97e18E7Ed34Rl1qq4vtvxxGtldu/30
/fxs1wNiUiaU+Fp9EKCdBp2hPCImvbmsElIOTiBxJlQB28bbIKxFkCfO5FM4s2KY
t80h3Rd3U30I8GUVuVDncLxFNwil5WWSitb3gMtKdEcNhhpji8dnDoc+6yENRxJM
a2D7Z3LqRw8ThlnDv1T8rsj/V5iqOwSPn/qmKtO/t0rMUe/+rR4MRzawW4OKipaN
mB28DlTAoK2N36laMv8y9WDc89yn1g5mp6phLVapofj1EaqOGZUn5vE9NHyt2Pec
YcVx/k6AE9SLzzKdu6SEiE+f92DYV6VmmWn/6j2B9gw9qMZ7SLw1LccvO+rbCjPW
OE2j1GjijPqlG5wnymIZ4ZwR47bvmUgUex3urIz4wHkIt3Vty5qfa+bdUfgvuRPZ
+CHhU0sVeDkCOxEw0FTd/ZMnavNEkSbY72heL+DjhCPMjQyT807pa59UbUG+1WUK
11tbIkfG82i0R8oyY85qhmuDpsaxwTqVnTYHyH/XxOE3MVWtBfclEbJxQj0udXX2
v3pFeB9YuC1rzk8N2uSFS2RTpwxTzC6hiv1CI/4eGWyV+jAIq89G2cYB2B+PBMQj
kM5LCdZcklUbnadmrMHKzCc1MAe3mxbfaeExjE1UeR6FvJqxRs/qVmb9XXrklZ1Q
80kTFFeMAG/rQwSHTsetRuA0ZJw3Jr8xbQL4jsB5nS+Wm0ARHIt2nyCJ3ZoBtclT
NV6qwl6Q6YivkcgOkUhX8U1j91PCRBDq2zH2doRcDXgPT2zhTkfNDiMd8LpmaPeg
jzvyxj8JZD6lMumukLKvFegxSn4fGu+7523ykedvl7kPssRxjtiQUh4YvWQX0W9Z
3UuCeQUkdcLkfP33D422QD732EA5FgbfdMpvpzl29bCK3YyxfPIbJcQiyBHcZ247
YG4iZmvrmya3fTWYjmIMCDg25yOLS3wLua6kWnEH6nXSnxDToTOKyto9nV1H7qev
R2BFNUhb9mRYZPhuOA/00nGTKHVrD3oOo+KjPgB2vG6vH9HnB1yQponS8Ejnr3qc
tJ3CLY5HvP3mJCcrv0ThDtnsml22WBvpUKtX1DtpCt4ICNssWsVRhWoLwlKfanpF
oRapXa1aB/4BQkT8VwZazpBCTkvHCT+HC01g/8UCMnMei2K8Ik7JJOHb5sCu6Cp6
UQTyiF6XElLrbH8aK4yrwSC0RNMN5Nyia8Oy3ObvtJMiCMMyWLulhBN6vlOcvjy/
UokLzdAh2PYlTzHlP/WD61PjeaziCPcws09/r4vaB4pb6tERuI/gZeS6RoVoGfM1
mH2/TSFSKQXYC5PBxpqMFUaSCc8RK31CyR61u53mxygSr3kpbpT29NdyWsXGptd5
YE9D17gh3QqxojSRBH3/EZm3ZwkzFDh6iB8lzlBxuzFNR54iaFtGH9ovDSATCRES
O/sEB1DgaOFZYTkKmhahrJJ0eYTf3Zu0tTsHUYhH4j8YzrjrXP5KRQKvOGPY/iFZ
L0cdGgL+4SAvZxTFRRwZifE+y5bvjPEEyE8ohh1ihdI2kW4UtvIqhwe+2IHoN1XX
deMoRTXk0Ok7opbGWNI+9mJ65Bb1Q6QdKBTvm7Xll4oBpqXOeNjtFpFFM4J/v/tP
l7I159gxLwwBVCs0D6kE6R4y/24VCi3tI02pjf6nk3i99ngIiTiTmFE7Cq1z3gYE
ZKDiMHvX+hSq/gS7/06UP1tpoNN9iDrA3gKBS3YRarBL8zWyTdzZdq8llLFfv12i
KGcLqF7dxebMqanaUphks4qUICMSYjByB5JOSHM24iSESw7+ZysQLIq4ID0q+5F1
qtJA9NihTC550aCedN06t9c3lkcJR9YyuV01Q0mt++jQ2efstD3YsCLvqu3q5F9a
36kVCz4F2a2r4riw3Bkome63EH/xJPsvrKipUV6FpCiDsUbwfaBzGMIuMuxOYUjB
VTnopqWyP97rqpdthU+0N4FmykvU5jk6AuF3fI7O+Xg0/3kZ3OsvmQxXK6WlWncL
jHkG2qXEAftbUzvCPaSMvvkbUJBv/WYn23pqhEFdSIx8yzpv2AAtIeEIwPRC+Ywn
rjkQ+ISYfBiG1EEA0mLF0QHzAWahg46d0m7rbnv6NI2+74JsI0o3PqeblhRv0WAO
H0w7k3A8XoaJvy0FsoMVb5h73aWOBYVHKwpX0B2KIrNLk39fSqvtml+Nbq89alRR
kW8AFrel0y7sDksfzYUVojteiuoV9T6GFvIllLJdx/wKbYxnglBBASfSzDCwXxdT
4SsB1ds9/m+Dv+FrEfQ2fMGx/redhPppc+QVexKG+VgHtWn0iub0JgjOvkclnSl1
f+fjAiB60Jc06e8x4LGUy/ocJ9DoUg0JvYUOtbfTA16tZ7xASbHAWxhxAGC9YIJP
Btn9Xmm2rT0y4KXUqkKkQJZhcU3xd4/DZGOujjp5cjOw/bioBCJ1uCY4V1Qo5p30
/Am4nWxqMJ7+kugD2jSzuRlhJdwkMl/282Yuec2AiK5lLqm2W7v3S+bn5y7sPs/C
m2/+v92t7zQZD50RyOaNFztQjN0b1C39vIz9tftIt38ajnXeymRt40UNJeaPLC2h
N5KlotcxObKA5aUGE6Qxy6s9ghwpWboI/6MglGW5P7Xz2+2d4s0FauEb/AFR50hu
olYrRddaxBM4YYf72NmcMMs0NJKyrvRBqFSUHu7r2ieHPPYLMF3jX9i7JLllsxzB
ke85QhQvs0yLf/upKATT/xGgVYUwg71EcnrgsxnVmj6HcEfWMkn8TJvDwy2rm7pj
mgAFcsbp1OIK6J3ja3bRgaXSEgVumStAmmaTGKuTivTDH11xGGUH1FYnCNQKQgB7
z6NYc7kRv4OSAtZGS/0UVnJjGmBJLrpZ36TEfX/ojvH8FJ9kLILnW7THSG/VHgKu
VkYAjmV4RxVVvwjeITORIif2+LoyvweLiTKpJNVrk9Ca2yr/6Nozn/+O9B0Vz4ch
K1nTm9C5LNIHKaf+PLKKSdmyzRp7ewH6GM3sBZbkWSwfdYTy0dVdTM90CVvEBEgo
a4EPOxh6/mI0QkQXLKG1f+Wn65UhOJgD/5ok0A33C9GKHD7t4rA9gvgYk2IqdYlk
hkfVjpAKOistVNSbjkJiuWV/E1QmQae+juqL9GsJF/k11zGYMY+pRdM8rnFC6JpZ
m7MTS5wMzYroULfL2wHdJtxfj/0AtgYotwZZJdxk3h4DgP1YpOr3NZP03rztoqsd
zHov3GB4lXLAStL6LCln70ETlu8iBi2R/X7TcRQELITvM1kunaLGj1arLO5ndMw/
/Tf8PhRsV8MSSfjods/h42Kz7a1Kncj6Fjz/brCv9B1wLrjz4LuvslUcAVwZxEvJ
HWOqczADYsBQDGXGqD34NPAC+8VP/Yic4PNdu6iZNNhdpm1zs2bGKFYZfpUrt+DD
yY8ol+7m+xPQFGeVnPjKzxOBZeoUFhbpMY+LoqsYBAXr57x90dq3WIEgE4a5tDNg
5roJVlQ43GxSF0pe2d8C0eruSqQ20q3KncTnbiV4amLZrGBgKMdlCgkpU8AaAPGn
U8TDLXoLJq9gML2vfcJbWy7qpqlQaNIc3nYPiUN8wjoMWvfSkWz7afSqo4aAS/EV
hIsPJJsy4qdgT9AmdKBFMEI+DLNbP3EjWplJ2kdKDeO+kJl/xdYX8srqElXpeBO9
1yswiSi3BRLPWjuqAIsK28zaU1uygYt74Ebv2g/HrUxTrOP4CQFzgXLNY8Ko5PH/
fL0p+Gw+0q4dmvZUuYjUbuhU/KPo+euAtPaPFzoFoXJoz113fFPXsmXFXMoc6Yyu
lO5z3sXmP1WtS4JTyRyH705mTXUnlQL2HjyFzarmT8JeRMF0PaA2mvRPfdne8Uh9
UCvEv0QGwSgnBz2BgHQwCsKIViphwokAKoIgmbVpjoQ9k/07y4WKLoJ5vnzLAepk
Rwg+PnEAyDYucO9KgydEQpMRGEuLxB0eGeBFZvteIkxEM3PE8GTCGkNVIA0QPghx
ZDJr7RyiA0pVUWFrCFf+GcO709pMSxIfqbzvr5FIdsjd5AAAhjtfEuRJvDiYF6SU
S855aYUSUGBmEeNzaMccQfVyae9HV2WgXiuZR9XS4IM508FrpSgkyu/fZNy1/WS3
d61Hx6RK9eZGkNhXp7UbRJ4t4Ovczp36k3LKjPDT2/t0uweOIYyDeCAbS0HzaaUj
fKnhfwPbswbPiOEBBpw8UYvfcs+wBMrhd8Ic+Xf7WCXPE9bKlz6Fn1rbh+g6oTnn
npjpxQwnCRcSwIXvljO6pQyNpLKAc9lvJb4TX7sMz5k4wRzd/cK386ayy8rClO/P
GaCZ3IWE3qDBkWezi67mZOMHnmdFElYCXL+Y42z5aFska6JxzoFdxvEkZ/CdCqw2
85lYOAWy1chNUB8t6ODuH5D1F/ej/pG7Gt9NwQlXrcwnoiYrBNDJfaHsRc0+yZgR
cko47RNAyqIetY/ZUeULrIYl6iahQ2uhHpIdK3LVQ4LBo7HFDZXITOCr3saVB1m9
RINmxMHpqm5fVM41n8wFdxH6aJUZM+mq/foLARI8X6L2/gRCHuouPRBbWChAVL4m
uWwfJq20l03yA4D9vIiy2fPiY/M0xlC9B1mcxbxnVkMUD1q0ndDhCi71G9EHfhog
2xwLiakaEsOAH4nYVMZE2j9MRVeQU8zH03hEJxMq80IfpFeYfL7sx420mv3oOnVf
4f4mKzmEl1GRvecoC/64XiFid12djOsjqV2jLgq4gEC64+/ITcQKlAjfP20KgIme
msvMbPa84ZU3VRQgBWXDG5ZTHzI1BiCjBc8JGdkLqq8Ey6AKxtjtB8B79zEVKHxU
AvRCDekY1yuhpdMOB3oE7NCjQD+ZVhhefZx2NJCMdZvz6Ouvvr/SdE3du8OwrCDk
SRZ2xBfgnwexI2NrVyycX/oiAjKN+SrDbcgwy5B79OAPsmD2+mapXB1jzzSCXRvw
Bf4+qpKRoy+MuxolVmkTQnNOMHodLgxV6P4+S1JVo4j2/lMXqmOl+KFAI1iCDAtk
+EjMDYum9/DRhE8ntDt+YB61nasVBkyYIN02V6sd1GIfRW/UVNpqt3AlWHUazJoH
Sl3U5kj/YSgsssbEkVY/X7o37GXV7l88aLVoa8FjmwrbN7LnZdhxDfzdlFbUGaAj
ZhKg0Vjmj6mLcOblCOjAU0x762NXW/E1I6mjPoJDFAcXlZrSycDSX4DW8rtpsUPl
hyhQtAnoJHxKTd913xBF4X1HvVlmiwtT7J/sJPT/pu393QSOR+gy1gK0pbZzbpYB
zVB1LT4V+UKP4QdVFl7tPxPyVXjbatntbG9RKC+wmMJNUCDHDQRm2vWTdf6lkcDS
7sfVspEV5ZZk+uVImt51BxfA+bCW/FI4C6MkFI8SWvD7ivMbROmqurJjKIZh/dzq
+/CUYrTwawwr7r3aJbdoV94QD//V1KoU2zdWuMA2NHAjU2ATS6W6m7a4BjDgQbn4
S+9qYCQsH8zoT39TgBLaH/Cs1TGCZXChKcvmxFNqf7Jcwhom/pk8VLNcbEh3ZLC2
gWZx8cIPQJBeuxZANKOLRRC8Zt7n72c5Q8v1MP7MUb0gIS4a99fPiypDXbKEbA4z
rar0++nVzwZktLafFX004lruwL2upkuIoO6OiGcgU230i7iuYlAQqwEXrpW0VVGc
5Npn4NVJqY66pJGGZtS/kkhxrBUw3DQFAvLrydfT8SPJ//t3z0KJeQA8rF2nQx6F
3dep8zSIan+TuVP16QDyaXH7YdpwafUMgW6edYdRdAHmWkRgy1MCkZd/wIx79F2H
GWPd6SZMxgrM7YTFCxReeDBcguDH5y+9CQdnAEsqI0M/6o2p8MoBoF69WN3dopqV
iZcqWEb80nJuaMtWOH8wcB1iBehhFlKQXDveHFNVennnUynnByHBUj8qA8Mnmjbp
tpB19y5OJHA02b8RcRSVXdhxCFmkLsQW1S0U1ta+h5FzxN2zERniTZwYG1lP1RPo
2I7ciBwCFi6xqHLZr5mkf3ee6YhCAXi00xBcWNkkSVmIKtgQYsmuoBCVMCEmkkt6
fYqd+XSV9mC+Xa2WHN8iwmZf2aVsZPMC/wv+I+0v7Bz+ouFxI+rTNmmdKaHchAXc
+zX7Z6v5qHJassCT3bBMD/5VRLjVGiDR+9NrWyGKcHq2Ypr/3pE/qs1jsFQFoUZ/
D7faAvXYmuWbFC7inrFALkskjT/3P8S4du7cD6FxB8Nmhi7YMGonzyRR8zITeUSs
Q7NT0G3/iWRMxxxLH8zX6CbkSKik/65xfZwUzE0+SSWNOmr8mWBE5KdIZ1SOjcpw
JrM6cMOB1I4XnCig0E4K3nEw0vNyMYR4vt7hUk3ef3CVUjfL0ZQJpmY/C/MqXPLd
58v2w9qfSG2qUaXPEJjzZt4QFczEpPqJmI7MHu0XeKsC0egNS7lQkrdIGEAlWciF
O5bET6lfiAAUG2u4k+cPkn0p04KcIclF7te9RKaHc/tdrcLn+TkR/5Z198YVme5D
mYhm1pnUFaART0RIE0UnI6zaeFyHTpF3MxmsH2kLdxr9kGM8+Nd87k5eCdHdFbD4
E6A7EqXMnMuUf6uA0JcGUWOdESQc/19Y0OZfaTqd9c0HFRfGBDQjBBYqvyrUnhgJ
jPDvMfyxn0f7t8kzkcyk+J207KPI0BxHhiuNsKq91gHOmRaesSjlcB4PTFaj9sLD
oT8SNKRhDz2es3HHPYr8DE2UqNFBuGgPWavJlUz8e0TAWVGSKfWX8AGG9MpLNHqd
9qbI3wrkcpAeYARGwkvwFZ8cTGPsX59QI13YuCJklSvcwTUA44SJrwoMWYeR6CgB
RmatWn8zSPEAGr5UhCPgt5m9ibkvvAEAeJtGr5FHEOeTZGPux5OILrRAQNyKJ4Mh
l7P1AB/qIiFKGQu+KxT97YuH1A+/l5He6nijqBnDrzbFWlJN+TEMQzClo8WJF0F5
lMaCJq7SfpcTiMDhqIdyk/GXwN/2eCFWWahwmr7chsC3fb8opjqF5Ir3aOxyuiII
Fvh+/R67G8i+XXoBPBpqBWjQfNqy/JQsHv5rB6rYt2SiovGV+eyKtMPtAKuawG+O
L9tbmsMWEqpAAEtcKLDNby3mCQP2n5/8Oi8dVjX18r3uZM2yz38A6h2u0SBlUoZH
d/k0BAd+/pb5s7p7EPqc/SiSdb8+oncO8bAA3ci5bczn5hZqRtHgOQQsZieVL0m+
Ubd6BGmQ4t2aAeOA0LxgIH/Vh6NHa4SX0dOEs8q8W4ReEkWY+FUoSJ1FIzyP+/98
4xyI3a+yyKLVEtWRmMJVd0fqObrgkQ3t6WCYEArIZqdpHI/cpPtp7AzqxwCA6tpb
MOpNHdhlcb/P0df0cJiKgD4MOWEU0rdQbTTUIhgl8gjxqA5UBiUz81i7fFfPwIQk
ODuVp/ssYPgHc0CswBl9kIkIHj1qMIONN2z5DQahCppdv0LqsxSakdHPVCeFMroy
POA8avmMO1+MR1HG0W/4dIpLDln8ikNA1LDwdH/qy3sY7gDLYkQSuaVLMLycVWht
ldUFdvjwQVyn5toZlBCKt4itwcVhhpb0C2phrpWdLhWn4jAA+jzw8Os3+dPN43Pp
5RMT0Xd1OaB0n1BzLWRuHDGGAGbyP1AY6Q3JFuPk+5lGj0bcfvcogHk8NHY+P3Cs
xYXGOWeDsbodXrcpf07MAcYR2vv9lvUL3wzS3T8IU4nWKRDJ5qy/o28Of9rhtD7f
dmtF6WVIblX/bOY56z2ljogsbOluYA7uw+RhdXr+0+Tlr3vLWQvCHqlbeEcqo9X1
lYzhvjmEALy6nK3+uRsa7ZLmxy32dnvURxdrLQCk6884pFjuoL8Qnfu1ItbzW4Su
4R3jjurdrlHPVuYD+TDQbiy+WkEVPCrjNNJEU6t/6ozfzJrVwoeWl0hUj4krC+FO
BhCsk0Y3HJLzbJUxKk2UvbDLSSFuAL84w+jTOzLFqNcipdPDUEb8uSuzt35EnsEz
U9Pe6How331NPukQc1twyxz2aJBSXVo9HXbZpc3JTRHQtzljNyAxsqXlJtSPcs/R
YYWaxEY2b1F6GfYkUcpgxUO2UQwEZdlLciVn8oQq3OIrBZADxPN9NKdTAvyLffWd
S98OtJBiptiu23MiL8tcYHHi4v6m3fg0ZnpaSXZejPipUrl7AATOQI2h4UjK3zVu
W5DSyQ1YnR4x58/jnBZL+QZarUm/wTEUDK+N0+S0c56sRzvqwDYGhjkcG8+gnJ5S
a2NRIVJuPg6rQItwJG3Zc7/yeYr/jzcSv7GP80aO9hYgHTGSvJ+KXWxN0FUaeERM
qLc1/iBFtxLo38qOu1J+lzlNkhoU5Icd/+BNIJl0JIlBVDcPM2Ccab1wOMmqBYNe
SkH4BDttTJ646+t62lwXs/fRw+NxaLGttKydklWrr6BzHr98T0w4r/2foDMIkiB6
xqNGngf8f9a4RJuzut+hgozKosErx1Ku9ODUF+stmJeBFSiQrFpzoSMU3FkLnCtn
nQ/MwDL3aoDb2rZxjdnqmbODCOx/6oQtJEq2iqO0XHOL+vounDPb7F/diniMUJ7v
QSG0PV+jlnTtyk+3U5KH2oS/rk/2sfXn6nB2RAJGMXBE8ytBsAIK/Xj/Mtj8vco4
XQ83Cq7+N9zMCNddQqaBlfD5iW12LdpSF6KljAvmQD/F3cnsATaIvGo4np9yEHb/
Nnc4D6MNpxG3GsPGLIRRh1XOQfW834m5b0tRUw4HmRYRnSuv3pu4ciZ0Cs5MoXYC
DsZ0S2sMOQxTpi55XvNkhyf1h2hI8Mi8ItvzJpI/omxNG7slP7xy8NCUKuBI0enB
CXu0mMxa0Yz7E9q7ggf1wdi5WiTnv3jYBpPAtfiDbS7LnLBOHsUMim/NErd0uh8M
kbN5lqyTblHd1qmV+D0nwyvrTOXsxupIupyhUoBjBIdu+5Ykji0O1392ROYKCaWt
kl2W2FpYKzqG1Z4cN9d2hh4NTOW8jghM3kBNZZFAA6Nmif6maPARRhYJvH7HdILU
UmTZxM8XuIWa+5EWRSp2MszHLgfM1vpsVS2xyl55UkYRU3cQNwQEqByJ1sBFjtuK
blXLm6qwcf5/FRLcN3/mVhh66E01TtKA/PNiCpUP19Ozl8439dEcacQZ0GvQvaaG
9SjeJuaduH2H5RUxkqj5/tedM+WVLlJiOnAeEKUAsV/z4OqiBGe39elPs+Melj9b
K3ibtr+4TEDLis4m08GMthLkKWQsIAL2cM8bAZKXJZ8EgZBtCGcBN20DPvR3xrcW
7546MjRhY92cibKIqFqzJcSUd6s0iXThOGp7UeEpRLzJc6uOKZYMYlcAJw7mQmXl
MHg+qYeX4YAXVeG98M7jq8b3DxrpBQ3ZVjgIt4SXVGkWezG7N1yzgAfXbZ0D3EWz
+llbfCQ0w9TaGMj5U8nDRL6alKRBOZeBaEochEVrX4N9SezUc/y071F18jL/fRPF
adNNxWKhBQWBNehiVqM5t/q0s+qgMbYysMI8ua/TOu39+KQ5xJYISP1qXvcFuoS5
MGk2F2OJggx0Ev8wnq+MA72QSOGAFBzNrV35xc0sIpLacUm0JpyUJcLHok042GL3
Frak3lVCxGwEQROo/RAjRC7BodcNX9rHY6d1zTXFrsyhMio2z0lBQztHOP/uXRmp
Ot+uZ7WZ1RnS+4mklh7sPo5sgtBgqvY8TWHI3SjDRBEuTx21oVQ2NJKR5UbHmmvp
a/zsR4GCQIphPyiQj3/BLJFLoUk75PxYk3a5THCR+DEDEZa0KaoacgVOw9OB+hr7
8rSk44K9nFLO6BrF5JSSUQJWNxQTgVWx5LTqVGbJhyPtYKUangGHxVVIVOXxSSK5
p+ZD/AKf8WZf2C1eA7X0SoC2VSdEZEMBTfDEaG8+s7LNtuoDEYRfirtsX+P40HNO
XLQkgpnzuk9R8iXmdhouypCzcUJxgmNkS8AYDZkpjOSekz68mbLdPOHV8myjGtlO
Vsy6JMnw+Cmfm5LX1RIYx/LRNPfVaAZgQWoESuujzmtThx8Wb4uwGlWTB04zJkVv
CuZkbqQxIB2+0yIY7k6FfWY2srcOG/zLvnFi+ZK5yTysKEJ9qHhvOIj7HmzhDr/s
UCQ67PKyS68E7vyjCr0gmqAeKl+o/qXHOQW6s5G/LFPct3rDkZNYpbAhpgDg9vhI
f0TZ7t78fJEfN3EZ2sUhHk4/cyLkIb7B0UqsMaZ31V4GRplRjV06gknru4EOd1BE
4fLsO/4mhGVK46om0Gdh57Rs0+w0iwGRP3/Pv5j9G2xFsl/tHeF1AlglknXKzp2R
4VG2nIpmZyJlC8phALkuRLnKtl5ICG/GDpY5FetOX8h5AZPx6SdvxoRdDmHaLvSU
4S966pzQMgP4vjoM+Ul93EHgzOjqh8aR2bCtw3QxJeBOYfRM+8mqAXmAI6NWhzyh
Jufi8p4bbsMMULXrdC7mQGbKYRM7ixXfhHaQnfd2CNUVGOUQgXRwws+Gn/18fiwB
Jk/2ytTwR+2dGsha6BIZN59EIi2f25MCxRi89z0KhXiDERv25+dxXc2UEFtXitj+
42CcnWrUjV5rzD6s5mRhNs3J/CAelt8XS17Sqz5HYs1pny5kaltNEkKpVneYxdfC
kIzRf1Yr5bCI0GQCdnLO1Ce+LpegiIYB2ij2KdLUXUroDyiTMcz/chCovipKKLzU
9iPRia1JMrNUmaR89a4qg/et8Mo2PnTuzhXUSXAYlCbqVUwZ745XoBo7gzkrOuce
JzisDH/cWtxe7mvXo/2lAwON3F/IYitf/ijPBvy0JMJvP8uPvLT4u7SOeRJBclFT
g9TpeMnmPT5y8dX8M916/K6sL1vdwSJOFPjqHuKW99tiMFK0S4+aJtQu7z8tC7iB
VhzjSSzmJ59LmPxDhDDjiMyAQeU6zqXfhn/U2t5HuOdwGfk0xD/F7rXm/RPloIdJ
TKk4Jcdds4BMoIDT7MslTXPmXt6ex/CuKjQB+pE7MufhxMvBlYR7c4uKjDuBo8PN
fYv8+okYMqKheC13zDYjmIrEVd6fmF0TbuB9o3csK2tAsJMgNMjzq2nOLYYYJGHK
RWH32EXID7e75EbZQDf47FW+0vPxBjwd4yvMUX5FegrEFXo8LMcvJ8eGZ8L491jC
VcBuzv7LbKSoxusOVldnKTle8Bi9CBEb/kj0xT7YmfzGsbAQqMKUbTQomIWTWBAY
BNr5lz8wmvmRSaHAs+10QjMBrLOVJOez6Zpy7387YqHatIA1IiKdOTZ+iIdwi1oA
w0e+gjkoW6vuf/NRARf8OOWYjNyuZK9G2FN7nH2TDcZ7iWayczheHTt6QcDvQCVz
ypjBLnXeARL+/Ug0vD/blRgeMfq3kxmu55MRkw+skmWi3Z3Yi3cG7kiVBtSMBUNX
xBuDiEYpsTaeZfdui6+vbwWi2IM62Yizy0jqLP6JHHeluTJ0JW/MONoaY2qSFpdH
MnobXqV5JXl6FFV9Ax0VbeD39kWgh01z5CM/7T8EzVGsCXT/dG40jZ7woK1lC3Hv
m0tv9+57L5Tf5BUV0r7G1+DHE/OWCxqV021YkduWLZhDqRUAoHq74lK25MgUhVYr
giKq21O98ZvASYrwp6F0HLc5yrn2Iv1l5NiMdFXfFDKNy7H7PvyO5wWvB8/qAETL
mrdqcK8I3mLRrH7e+lrtpPVspQihTY8cH4qWaWirpNKNO/zA+XSRudxNNYGdPvN7
XuA4uRzGFh1Tegg/m2wjlv/kSDlszLKFGryp/Jz36DYRSBi1QnAihfmG3XfUT3dl
SUepDtvZrP5raejyqY+7i52RxCaUa0Lwaofy/40F4KdM7UcnrUUykToDCjZqKmOw
wOdUFd+gLVEtvuhr5ZSoJgdUNJ5dINk3CvbicWnmHx65iKoTbSqSbLf3PhrswO64
NCCnIr+Q7fnulrHovATMfRDw+SiLW5ORxyNd2ZxpFeP203gvWYdPUylBBUq9QFy0
PxEVkWP0UdUKMd0Ol+afli83aDx7WFBV9dPg9UflmH4t1SBNdNxJozYl5iE4Argl
sikyu11269/y7gGimo31cOa3o0HKmtBszQ1VihbLXMLDE5RIb+kKwRLvtUSFiQvm
o9oNTJ2J6H/WfUYPY2aVhBDaCDu5gcfFveYC1sKWOfSdIYGeYO9Gpco1rS7Smeu9
kxP1PMM7BrA22iE+3ZaV91urBL7S/Oomr4G9rpR12lNob6LvdGC6Pa2jS/Xb3zF7
/xYAXUmpYF2/xVKHCzb+WIGwMTqlSrPJqEhtkVnVBaqDaSEvDRVKdKdvNTYA5Hf/
MnguijSDUfoexdfTaUMkm3ZDwUANfJIZfjPGhPBz5UAtg8bLE4NQ/Z6I9SoA4VZn
txpN5cO5axOV+Q0oXlzzTAP+nc7zWHsG4oxn+L0LPlFERLD+3oXplmjqA1ZNfPOZ
7tT3V8O/5Gc5LI5XnoqHkCOrVu8tKgLa/R4B/L65XDga5ppWK6q15MVognRRWbsW
fj9a+T4XfbBl5Is7JUoXjet9cw1PQo3qWWeD/uTvlCx8vZbcV57hGSVMypjk6IkA
9p0bjQYls0R17zowlgSnQt8cap1loCPy0vntqgIgdaVP2Wu1BKqX1xqgT0jllARL
j212UvBz0bpEXSuE2JYFhmiYterWW4WVao06pC0a/iw2ZASzWV0saNpBQi5jmIRC
1ytIdb+nmCHWdWp4sZ52rC5fIKW6NahF+Yi/ZxwvCdtWVhqMeUFBgOrG3yxSaXYY
/gXvaZ7b29b+0gygZRbgaLRBmZnbE+0BukfniB77aiUqJfqd/D/vmU8UdbcvcJ15
wpPczzq4NTXzlaQHm3XwJM8n+2q+lrQf2CTlATfeIRi95pYdBd0xBHEbG1fzqqej
O8jR/KyCYHKIeedeLzf501YluqKWz+7J5cAf04QOzIpvTdPjY1svBK2UD4LuW0oK
o2WkAybO1k0iyg2HTaOfbYhpvGmHR96hoRm2mjhv80RCVcW4X5YIJRmh6sLnbJbh
g0f6PlTf8PGn9ZsGoXis54gTYTzxIZe/kq1qof6713VGJc8f4Jq0QdVyZcEzWe0Y
FzXJpMCAPMClGcvXGb7APBBRk2yFghghHbqyLNAS7KgviGEdnHB4HrloO/kSYu3q
+nWLrdVEGUGX4X1jqNmVozB8SYH2jx4jZ0emOhcqd547PDOpVK5DiRmlyA2TBVBd
Sc8viDN6WLHbzVcQgYCxnjoGiXRzjTK6y45yIl8qMyZFbByZg9QAZKMnkFJFTijW
F4G7BiQTl9/Kd6SF/Ex13TDdv0tiWcU29hTGj1iOV6StqhIVQMUlW894XEVHSaGY
xhYn0CAhftInWJN0FwLEwyMji62qiUXSYj5yrlkC4vPrqnvOAU0XmD0eHe2S33fZ
VsKkoZK9kyt3q8kIrEvhDBv0/VtStpTec2OsDfWulVn7QhB/ZLW7qDR1p9atPSfq
m9r2qAH4SQMvbLqhmvWY6t2KyUw9bcXNrmMtH11BSnMwk1aeo4D3Y8S9MKFoGMxn
owE2UzzHbVsmpE4eVTJuo89N59Bi51Wg3wMXFALv9xZAv+5VGFCZPYCm+casABwy
lMN0tPVS2ZWlrRW3wm+4d+VgwYtV87sZH1H/jHd+ERg4C9CYAirQ3LtZT6T/u/fB
ttZ1KWwrUsvz1rblsIxAILlQTXg8738mppusXHqPvMwHpGnf9R3NcFSfMzJrdfLm
syIJJpZsQOCiB+QhMsRYcY4T44us5yOpL2gCUvlBkqEnaOIxTOV6i0u9PPExW6TR
LnBS8alSsq6HeQUnQxffNXJZFFuI28MLzUiL5ePrv+JU2KHBvm9tTaf0GqfgzIPO
6yaXCCYdhbqfdTdEZ56KxWt+kjtapeDxoKWQ2qqQvUtRNDA+S9+ZA0iIPz5eTvry
NWeoWEsJGEE9y5VQD1Rc19AmrXOjEf7Ezs5FrjFwe5d3HFTGHyfSOWId6yGRHjaz
/VySoJvwMXSmcitLxZFHnw0cIOlW1jBvjjxAy2H8DlCwXTyZpNH2gHgP5QoLJc0Y
BUQLjQVzdfMSKzPcnbnpJo/ftc/0ypJPvM/kHM80J8xMjC231B8qk3qOzZDRY0bJ
3pbOgSE4+dMtm6J41LOqH/jrWA0VHWWjBRNxNjJQx81rRUJKqPRjThbgY6GpLuEh
dpBQe5KGmxzVEHd8Dus2AHydR7tTUCP/4L2Lk5dh48UyaCTvnqD5BXERZ4c3qf9W
zWcWEPKVrnQ2mgxABIf5HFGeyBOm6DvzLGK1AJd/TH2evaIS6ZsqJ+6psx6QzQV8
+vMg9weVk17wtxw96J3H5jAGzGGxdjMU4PKFFlYLo4dP5pH//cm0xyjPNC+TyNLt
uZ+KLMpQGvDRWSfIVmSowvgHOzPmZsA/k8lVuEzgsc5lCRTy4Nbxzu3v0f4Qe7QP
l1wRYpNZqlbA0oa0uacPjdVHyg8hnCWCEnhiT6he5QJ4Q8IRreVK6Akv5B3oWMu/
8yIgRnv8VvGvxYaJIHSfLHE6RNcD18Brg2Cq2Lq7IbFrFjQ6mwy78NwUzl2CTG3p
R9uaBsvhzU6zUZlkny4SgfPdfCXZOXQyXutml8iN7rsTDsasAmG0BKsHbp/EodrP
KXqkOKgXQm0pzLPp5gUEZB7lEodhmcFjwh+x4nXjp4VJkFV8r1m1WdYHpwjvh+4J
+iRk/Qi3UXe/NXyN0f9eggCFrJVOZoAj4aGj2d4MwS1i4wRNwwhPAor3uH6YqnZH
6VtLIItK6QgvaA9mJShb46tMklARSb/4AqNoHN47w/RgVZdGYw8rSKMl1HZHgOeG
liFOd8GH3J9QJp/VgCiDjpvBxp2ncoAqGL0sBCZ10e+I7K8vQxYgHJk+iU0e+0I5
A9ALOg+Ted0x7MT+Xh87HqOeibExiidNgjr37Kq3kSgxYtVOs0YLiYEEv6wbqmhL
FoFjWVaYnd1ef8iLYyTsGSU4mP5DzBkpcg1Dj7XKLLQRIvJW2kaoAiSpd7HqUhI6
DlRT9DdsI6cpj22diMGP30m0OdVvDgQEBLDIuIgX+SEwtlMMTz58qEVKZntqeq2C
PjgXSV/gtCFHEMVX6mruVPM0H5ndgqJSJzXlZZZ6QC5aP2G3B12/DLSR0YpE9LGf
UHjxf4FdwIHYHia08gnflfS2zDX1M6GzJ8aT/x+A9LtA6koVXsw8nqF1rCqgWSFz
KiktyZscms6uqrZuUIZ+FZV0msLMTyNJF8dDF52+g8EoLomvmEZfB3COFUB6Lwgy
4HMpnh8UCqVCF0ZRVGRCKu/UVX5P13Udwjo3h4jntIDVcHs6MywKMwfE6P2hPT/e
84HhwCRZi4fE/61JC4FQ9QvISSxbcyfTXRyQBZCTZxbYbaJN2S6u2UPDT1gOl1dw
kKGHu9k8xt3ZZXuh2IfYdZFMXxPEM+TNiFg6tQj44tKFBEumN2MQ20J1saS4eD4q
VBYWF6VwZ9m6z77nsB6jkQYjGX8s/BGaPbLLbvPMA8vt0/ZzAOJ3TR2h2nm3RAB5
Rle1Vbbx1msQ+7wkME0Q7iavkEsX9EzILZOnQuBDBGzXzAvnRZ7SlDmVUimKkRXC
prkAVccZbMeo0xTJTFuhwqQOam8clQ9GpQlIfQg3eUJugL3hFqAFFF2bs9EIe3Dj
P4Q07xhMUy1sMj6/6GndTFz1pJCSOjkq3he9AqPrqjFgUpYk1sLlj1G/LCEjqqyj
eZjWin3dwygNTVou8Rr1vq/MOyO6OJpq+vGtJYbdvg/nZ342yT1+P3XT9ISxfCQY
HgwXoDua3d5JrPy2389tNdjDTb33dTsKId/fmD7y4zU/1hLK+ueJFlU/1iRuYCGP
UivcEdtrBWAvm+K8P3fJGuXlVdNajMIZ/PbYLTsDewmAUBrtuPwuPYah8MgXlxl7
t4DpED0uXtr12Im25df36jpQF7CYZTXHAW4Ow5XwZUvw/rbT+D/dtoOe7YozwEQq
vAkCbJvV1KMy7fN/3DdYXCbHUB6M1HRNk2v6B23NcYQF2P5j28nonI43tZ6+cdgs
AuYVXeoKYTTAK7LgkGOW464q7yqrQQrFPTQzQB7s94A0QH2eMmhY5SeEctY6QvBY
So8p1tBi678ErHjLMuAm+5Os51xjqDU4Iwlo4aQvY3iH56tBUfX/wZQqTJN5wt71
bA78/hksrt9Wet8Lt1ocW1AoXmFyqIf1+Q/TybZqd6Wq2q0uGwdVEU3nVZz0gafx
Pkm9KuSPzHq2zsKOdwOqQ+mUBR/7o3TGK9vPflpsmcjKxvFhglGuN3JgmJIJS20X
JWrBSR9UQTjircGDqM5sA+VttfKT8vTTqFGFqCim2o5HPijYvwGsE9f2bjks90tV
mWYFDNRZUZ81VwWEMmLQE68V59fjHVUpingBnqrCXQJmYETpYKtqjA9iIooXK6em
iIysCcfhdk4GKQwGSYil9Dsx9t74/F/tpeAIo1i9dG3EbhU/X/WeSLDcVX3/xjjt
70pd5FPySyd47YosCxaS0ghn0KnZmgGyEXfhROgEw4YRvh7LRbre0CYnvIn5cerf
hMQ+6me5bkNOTwa0ILTeujkaSZNtmf5TvaO3CWo9aEvCjqSA1p4xk26oJXfsjenS
sVATt8SpipFkBxaOl+W02xUVsFeuxr6v3o0Gm9HerL5v7CYJJ3HiMaDUm7EA9qKG
AjQFlT0X+1LEM0XqBjyIAjX8t4cGBUka46MigMpltCT2fYaqnKJm+ySCkgpna72J
iRna87n0Cc0a1xn814P/S+VYLjPW+7XNV19mKDHL4yE/MSXNgTC59Y/3MQlJFSIw
vjjFgceLO7LzuVS94QaO3C10mHCz8faVqrPGOJzUpPL6nh1BDyHB9ry2bspiUeWp
+Qk6w46iRNDnRV48IrWj40cbKUJ8HM7oQTadVBZjE6w/bm2ObIUESTnX2UGbf8sS
+SIhzDngV5+rfjMmIePlttGmNRjvS0IhxtpMZTZOU2il6+KOc51BT8OkOS9Dm8jv
YCIDf7tO1bkzuyBZxbrvCMC5fBP1tIyyZhRW3/cz+cB0hsAUAvNuZWPMXO2qXYQf
XHjfapkpMlmUA5oSBWP2sd4+JirCvXfe+OwjIcbiLbwDSd2mSfXxbx+T2+4MhNMl
ks+I+waYyS6+xgBlU16EEBqK3S/oTc5bYRTzLiI6v6roGvGCWyV9EAmU/dsl2fgP
qaeoV4jyy4Ro4fx6r1jPzwdJmAqzehwcrh6kNV5beQW1/VjRmuJoaq4vwkbMs8rk
YhTvCLULpex2ZR0tSbp41rVhORwrFMiBjytx7FOTb0wou+PqQveevXv4grqYulYo
Tk+R7ffeFGl0sHO2qAcoH42BeHIyHc1EbcbyXDEhwo+/caOhMmHBjRWfEa4DCEve
aW2oSx0DJYEKePYGrcpOYd3maM6g8YKafs8B1IB1NsdW+hWLUnagtyUVdlGj1bsh
eIB9HbHleUWxWgKiH4u7h998g3+h90232bV+69vOX3ZASF/phDIyoT9Wd8YBd4QL
eIlK5sc+EYTIasuewTHRM8N70FWYY+qrwBnzcUkdc67+7rUgw/N/uZR9HeyhraMZ
MSpVYRH0UbrIgnsDZP5RNkIYeAauvfDm/mRTjJ8lvFyRkGD81cr+/o6bD3ISx6hI
xNfFLoW+3ek22kxt2LVJ8rYhNtJAZuR+j93u7QMGqUcoyH4rZ0V7DcQKg4y6/+Yu
UamBoQGGqupJC+V+wJ9uBWm1uaBABipQ7Sw9EZazJjpa7qCjg9Dv6xfBqr11/qwE
xWKlSN/lXM61GxX3mEPLW/E3Jbp7YiFoTycyY8v3YjriuQaCXmsawjqEa3vlkrX/
5W4rrGC/bBkSNgFCGElnElJMRmaw9SbEVGfXi2n5hnMFsvUhNgYTD89PpYLCcWRe
Oo/46FSOTfMeuYTsMJElUgeORyVaNtmt8jxTsCmRHFsZf7pLaXIFKhoQEQIgLVxT
+FKMmJtMjTalCBuJr2whDOFEBwnbmtE/Y1ZrTwTlUn/M55Trbh9vVNIFlGtc5Syw
K0+onJ+1C6IT7zvQTCKFLlEKg+wJn3v5XV23NHaQYliY4Rgy2AeGRY/0ugkRYQ6Y
hGktKaavokOEMezNxBXDlAmC0FykxtuSwfhJ0SCReLN5PXxmfUqiif0oJ+2liEIb
B/Snv3fYPB3bmo7M+huujzpVWwJcvbuOui6vB4GOt4Mja6OuvIcjbu52/QTzxEXn
NXL4q/JxdJtVHJTm5Op7CzOdyLQH9E72NjmzAkb0TwuUx7rOULjWFuq79wsFuCcr
Zkp/MqJAAETkCuc7fchBOdpwuHZbpgcOf5keCYIOYs8jrC6zAFQ+HWEGM99BE7Uc
+t1XwWBFRkAIU0hYPFtZJF4Uhrc1bKtFrUE+5oO5MNBAjgdPMP7afKNUeNvN4I3q
0hxNreO2qfyPKfh9f1Dq0QMNwVpCvC4OGHAGAeK0Ca7rnDBmUkCBaByDBz0emtyI
Lb348JvOdE21FaSjd/umbAaX0ZhBewcudNOscDeNGMr00qVvCcHuOTcLN8SagS/6
Zgsg8r/RZBwYQlXKdsHJfmV5Ia9QFKaQiZwpDzA/YZDWErSGl/rZVTdQESfMSJdF
EDGm+VW26YCWjncIubvFSYlyclnFS2dpsSNgoPnTmqOa3Z1V4SUsU64hz0G18vaj
xhbQcLtl2QAYlzb1MAHigK8Zq6zpOmBlWNkoomyiKNYdsXJRzvs5ykv/MJKwDwwK
D3v2Kg+1N6SVZ1DBmHGkxZwV0zPMM+CtezfNV29PsT4empsB9oJWKAZ87s89SnEW
k+QELjnzoWY3tBujypVCr+AmNvzWzx/VKhNZGGs800QzuuFWQn59Zm/lStVnSXot
cGek03u1y4XSXfi1tSsQp6l/rbBYpmY0rLR/qyZpBynNf9nbK5I2OlNzZxjWlM+O
JSVlC2gJAFU7EhlG8ZYo32YQgHA5Iiil/ZOR/nG1EPJdjQTmZhnGyOX5XNQfVRiA
DNRxnuHqfFiKLZiF1EHvP3QjVdKWjrPMTUTQd85dlEipREqHJ6EIVkxnv4sER0LG
YOT9HJ54RrX8A0PKE8QVpP0xYVaS5RIaArXhse8AZApd0MdchLaondpoq+igbxAU
/gRmStnC6PAZAAlyO64M7shTL3DZOa1B8LwnPvX5a4uzYtSK3DnBEQqMrlt+iE5U
7OnAHTKD7r9t4b+78C5Ig5CrcDNyveIneF6JH1k+b9jlFySW5WJiQHxZo9G7oK/d
6k13w4xE8qBVo18dlWEcBJlPLjjnqR8/eqi0JBuLOQ6QItgjhOdvoICfXiVdK0Zx
xUfGGu5zqngW0GR1nCKFbIcweYts/THddVIl70A99yjRY/GXKLEI5i9q6wiAyyNk
s04KiG+p28QBQXayURw8DdqyixBzs/SXua5XFK0b5SoIFRjneElo/9gCi61AicVJ
oZppHlzdJcqKXJiZ7R0zrS1a9qh6ZlifSYunqucowgpEnU/9ZH4BW33QqTTN2npV
UBYcAMB6dAFwfqtcP6q1nHw6iVGtWn8tlifyOHghHy/HmfzP9uP6sLMyIvLTlUxw
Si2k+E1OuBYf4qJy3S66htfHOmiOOMLrmtVJAI9Gpp59x1Du2cSx9YkHRQOJoMsf
mJ9LsndfpID0buIcK53LMX2aQ0Oc81EmJ5GkBhGIGe3m/vlZyRdQpVPw2JQVwdWg
6+VipssL4iknovRfCTSyqejTCB3extFdemc018f4yvA36+NLWcn4sV9JVPXlmMVe
W1MswpHYd86TeKP4flhuqNyAxeedpSAltm61l2XVOQVpRUaExRc/yHqqwNc4O3aW
jqHs50lTdNUMCB/4CUQxq4M40+FLy7jvntHi5qaksWaMZpM9u8ZV9hHMq/uAuA+y
Lv3uGYH7YBxi4bgGD7PUFZeMCcJcm30LTYwAtDmQyzBALsfHVFpy1YD5J4/YHDrS
OeR0UGcL419YStt+8pA8+6cH72qjdSD/hHp+5z3NrkMmCtnltpArLvhSTZKRVD69
tfB0f1ge64/M6bbABH5/wzcBhsmzA2OvMUdfjRaljqyF0rAbMxa6QXnfNaBusSGO
vKKIdhYvz7JZZvTozhB/Bom/xVdKJtWUR5t4dUXucvEb0ArqFUYV/IFEF3ESC6OB
1vnHqvBbcX/uaRmyMhEDRfKiTjLNM9wsB3A2Dnno+XrWIbLNdWt1SKLzMuO4KTeq
c0SdDXeCzecTsbqcO9yQ/V3fgxFfPs8bTJaHoLdK9ZaYHQjetR6eFPA62LMtkuCi
EDu//3fNl0Gf/P3rPi0ctIRlo9TIJ9pZ1YAdEXYHslufHogWUrltY5AVP10SGXAC
tefM9Dhge8qYB/7iah+ks6HiPtxYA2lapdfjsubXMMIMNEcoZWNYagL5E0UGtU5d
LmckG2I/M5lMQccXgkMxSBEmFiP33WhX4xI0zzBU+jqKbtlAw+CdtqHGtYfbNtPm
xMtZAcnWfI486HvQ1vRBVHkTIeH1sP2OG4MFPmHV9QZ7XhHS9okxtMKT/oZ/JYSb
bo0uXoDngaZ6OCTOzt6oL72KSF0ytlz6ex3VwpMu80vHIFsqt9Gp/Ena4NJmVnX3
b/MAWD8NESpwDRsR1dG/Bq12/hntLZGmse4pfEoZBN6u55U1r0dvC1kZRodO9yFK
n40blsz3BtsUgjkEISr+fhKotJL1E7PgNrwkNYKlX+nxd3O8e7hYKFa24YmNrYlg
I5VM2HWn0YFF39Nb3Lpc2E8oofyv2V5rZ4hkodeH64uAc5gVohp69HFpKuBO+sB4
U59rPqoGjD7QiDds1IJvTJFswCfWJ7CUZ3EF8W1kbBdSzkfIZT9tn2I4yFiiL/tZ
Mp8pJqQ4pnJikiY5kqC+tMRqmj8U3iKfqS7da/dHJFewN+McIDR7rxlVSvZN+GJi
Qxq9jk+5OQaQ5qdb4m6HMW6meCmqQUJUcZ3hdPAfHbheMXF2ccgWMS5JozkgWK/E
MbIYt35Lvrehl9Q9atBpalsNiu5MKuRMvJf3LhmImmHDYsiXLjOW6eqi7wKbcLuT
L1DaeAFrjHDszFkefzfUyoNBdXl6BK3MKObFLyZiJ4oGT6mauI4FkLUBNWsX8Bkw
UlKvYWWHCoOi1ZJdWF5dusB+fWqm68eXFPFt5SVVs1sZm+tzFrmiHau8ZmTd+51z
+NrStq1gFsKNVcSMR4ZSYVC9SmU+do2COBZfhVhaYr6bLWRCvNLUJ6HhizSft/DI
icIQyVU3OypcOPAwPZIZr2wC2Oqp+llk7nhAgIVKV4YozfI7CoDp8ujQgcTAah+9
jQdmm4Vk4rEkglZNCASqOTxkZ3pb2EeCdLfmhF+8X4QrBk0HNC2WLUCYEuieC9CE
3jDAsLrm/c2jtumb2huLVKazMCk4GSMRixGK5OIXKcHw2FVPquvHCVqSETaSJ6zc
IG3ODdKoe1c60WuM0dGWkn+BW+b1+0ToVl9pCGcvj2zhYVpCFmXF6jYAPrI4FAL/
QwuqReG/0S2CLIlUN9UtEWbKdDO22RaizMgTBBQ33HZ2iE4q7lawoUYlgL6MGPJv
eVP2GcTiVrM9OhUDSx62pzJXc+uwNRYvzvtHKKc2etUv7VjVbfRnp+JVGhZov2Jl
gYuabeuLWWukmfTz014lzNaQ19KzBmRVbNJu6+2yGxLDhZQL4SUXVpbmT2W8c2tI
FAqaar0PE/5s5GFXaY9wlR/CHFrxobgKC0ohl33t4sJvLLkyaXzqdctvUK8lFwb4
MPe5reBumwk0sb06LBqIpRtzNOiEEgXzCUw4elPu93tg3NZyRXdUi/9rMM8AqjGJ
6MIIE8jyCdCHteewEmpUc936bareHTxxaJb9lXZSjwMcONAGrZS48K6v9X8RRRE3
3JEEYjPwacyhiDXS/D02VQmO4+Ggr2YNArjucazin7y9xZXl1tmUc4hQMjF0aJOM
3I4qoGXiohZRBtuAKN9NCUikBzLyiJwDw3DYr45lAtFWxrLw/g9KMCapmk5MBTXX
M19q27FdbMGI1TQ4OsmXMrVlsbSt8Zb2+AbV4tB9TQwZvSHjxL9cZ8LuiYMP8g9N
bMTJpUXSM0OaiQx+pLNaGYL8eBcDyMVoie3YjL5KdQcGtnBA4etYgLWcZedkqdJy
rC2A+5e1rkHhhlpklaiwduskGHSaIuxhLn4cF1oa2Pi0Nuhho/OF1CyBPkQ6mudT
ihpI+GCd4rFfH8rYTLidpJTLvw1Rq6znLa9DuUpYlYuOnHlGGpbwdB6dacCj0tEa
1SycadZpBrXAGlGG31IHsKNjNTnvRA1znzvnrYkcHfhQIsqPMDpukbl+oTDGmV7P
cd6oIv4HMCesKyW2FF5TLxc/SA7Eh9s74oy4vYUOxg0+Q5eC23GngFOmb+2hZNlg
Arklj+ZTVTPJTDLzDzFrppUcrxJRFLYplDlt9/1cm6nn2R9b2DE65teM9U4dJP5Y
XE6WdnXYtkcVjsHgY1sVyxeE58i9UkxhmulV9PPYciZqoIVmK47CObhEZuzL4lHS
npTGTU5yDftsLo7pPI+1Z2aazcwrPp7g16z6ZaC+gZe1/yMkp5DArCF2/vmbiSgL
vzP6ZB1m3htGhPEi/1RxNzqeRdRGIvYiK/ZGuZ3rXdT9CYh7cYc2MZfVfOHpyROR
7pwuY/7OtYye4oRg6sV4BkErH+eQHIgi5XKaEN04mSdz3P5cMquWf49RiCCw1ea0
3V6IFMLZ5hO38kLDai4SnIJxVzxJmhrBpHDRtfG9ODo75UMODN6kEU8t3j02WwB1
qR5LqokS+3OzguBPLQBnD7fQ0xDU/vYNjaUkgea1fHSSsjGsre8xpBBS+oO8GhF+
uhIo3nALSdurGkmOsUqQoeI7CF6ueyX7nghB3rr+h3JTzfWwGZNP7qX8oZSsz7Zl
6WwO0gfzO449PUSi1u807tvZKEC6V1iugG+PnZOH98qKo70wNxCaku0nwaA13Oqk
osdmAdk0ez7TTz962Q6cgGNGLovgCigVZ+jUh4MlHg56AEK5fhAfutjs+bdfWRIj
5nI5AcKw5qTpR0kvPuqhXeCT3TBsXCgvR3Ui6qxy3g7dhpilp1aR8mjyuTZ6r8Yy
NDcxbQPiMenjvBcr7XhJ5d2I3UF3qpVd6aEPoSo5gNglc4e6qZYq8kuvOB4YstCu
If4ZT6ATULfFaIxQ40aUic05DZyNAKAScUJ6l+kdeJiEREBUR9zin+2XDQmQ6bQ/
fOzIvNbyJ3tP4BYb5Z1o65y0gquC+mrA8JDK4jIvzVBIkNsAm2sN+HzGBbeWXlNL
KlhoubILN8hNcXIgIXpMGZTaIvO3h1PSy2SqSKMXAKBBpmz+gtXTszVboYBC7eUQ
gFx6+IL8yhxanI9NCuH6zWRx44xnb8mJ9I7sZPhukXruc6LKL0JkHGkic0p5lPIL
slfgltZVXOa1E2FkDKR2Zb8KLZdvUv+fXD5E54eiEpk2BWUkCACU7yQjpEO29moj
F2c4KEev60yNQm3naEZlcW2DCfXl3gwe4uBUd2l2isGkVlawiS5Q5rW9Tee1Rjwr
JC5xB0Lk7AUmeJtl0TVfJo0YWKWsLEAqeCQzXak98V3EhikGICf7fEkkynS/pVbE
23Qgz4zHsBzSUs7gypWPhrt5OVL4RBCqvgFBGbsrLviObQFR7Xwq2OEe0eu73YmO
tXMJ3QszA2zqYdKruzIeogbVevTQyl/HlVxKIdCOcSvEQtNE+HZVdwoDGtBxWk9h
Q20AvleKoaV3wqy5u7mHbcNjKPCxCj3rGopYIjRuhSLYHipFhP5oWIZjkGIk91dL
QL1hFqxVpQY7zsiqFKdbzZ6Zd05dllmCjte+0scOy+efXm/fr+1C7xN6UwCM0R39
wc6u+2le+p55icLmND/uPh/rLWUfUL17XbpwZFyL0q1nOKRJKnXtbNur4IFQEqs2
s/wjIsu7/nbGw0D2JR2br7hl6ixFHtcbq3akC1dyU5iQdfuVUGx7SrUhi2hqEj1Q
WXKEQUGu4vDEnDTetPjti+Ck1X4qxr8X6bdX2c+Lh56E26baeY7qsqDSBGHmwcT5
JwBNqzNR46OUa2wB++/Z/ZqHLnWA9GRxPGZf+1Qm8oG21UNFOBHBUjuNujgblDCI
DmklFZ7+Is1RAswWI3nRMbKy04LWH2YEYYn2FOzpcyx4pkc/xpHSp5W4HNLKB6n/
9un23hX15apT7cid/sxrBcMhU5WIGUfwQRsyKaHB4yWrsexKPNmXSeXgzLfcnK4o
LeQ2Bt0Re+cDOhYkvlLFBZuuxWePpYb/04Xz5x6mTcyLoJGWeBCKmEuhbdqnz0wu
jVYUXTPQhoEdIUxs61gtWUuAsyKByqcXpOz00P0i5K4QNjgmtwjMpFZSPrYyRgPd
ca8UE8XNd6ETQxV9xiCjybFi9l0dj/08kBRjqqIBA3EpbAJrsiKlaHjNrl/LSmnc
AdFjqEX0+/SkstjFGE6M0xXa2hJG0evBYDqHr60aCQFFoRATa60yVTdmrSPTWfot
N9/80jgclDrexmptw/r6+KhTJ9WVkD/yTEQhbZxrJQoNmmkmYY5+xD/JHK3FxkOB
fK4sudhs2Z+uXLnJCpNo3A/KuPFXuQgX0p3Rc3Un03jK50+Z+vrHAdEsMayBcUR+
SmV5FQs0q3mKQvqeJrX+CYk3F8rzXEahEGRKM7HbQ0YJ91/I5czbyLY3RoqyVtzu
WfEVYK0ETJ0ueuEcD8/hgo3VhW2LxKpYm4leKZ0ZxFAQRpEhlcIB5bA1GCxMEaA0
Jk3/5ISNKML5klSsgs04YwMoMj7C2vS2hhGwFRTHcqY9UrkeXTmxSEuZaVsgLZSj
gfAfhnq51Dy0wEMDKVOoWH8+XPPJ03tt87rJieNmbaF9V4nIN3J5m6EH6oDNm30m
Bu1d8l5BzK/OozleRYmZYz8ShV9FNqdaEA0cAaazGkP3MtoTieaW3Bf6h8K2WLzX
4XdYgtCSI6A0hNOi4a84PzNuqcaR/9gbclAsan0N+FS0hGnkJWR41dbSFOD9ryaD
yt7yMZkeHoMWtF1avL+yUNZZ/cpzydstOQIU5XaKtP7MnK0O7XAGcjSxP6F9b7yN
JXuuZcU5eDzCTrxbeW0LeGBPyJsi0rHZ6xfCpzulDZEXWaxPLPT7jMLOZyMYsr4S
DZo8L+dOFHiaWabkssliAULaVDilMsglG5hhgg6KhYRKGEeZ2tDGMzAlJAHyIFOl
Cs8Zlg5ghOQUJaA9evVCzOl6hvhnigSMsUe8fvSdCYMRAqCr7nJUMMJ3MGSausvx
XHYFmbw+gKuHEAsom2LwhCiA6RLtDsH5X9IAZzP4c3Kg0aKeXo317d/f566Wzt0q
ARHUF0QgbELoYiKm0e1t2pHjMnW/KhsippRlrfeFTKCPw11ysTKjTeSuM39GAQ96
FxuK9icsC+IQCW/67/F5E4gwZkmBrWDi5r5AMVzjnEV5xRyOf7aadADBFwL2v0EY
UMNYttsTbkzLTugSS+nzNkBtiB+vXNVZkHUTNfRmbZMFKpnd4FgLDXMpgNkzgT8H
TXTCWz0ArKJfiGLuxTBCDHSDNiVnSNaaSLt/ajZ4xRI1KXEcl460MW7rvMG3X+gw
U6PDBqa/OureZ4soAxMFZZbAVMV7DHfDyvdIXRNGcmilehgMDEaPIadbgG4z6j1K
m9gmO2ivnHRg/H3yOEQDDHNLsqhwJcV2GfwnBFOv39d4xp1ZyFeMbOn5mTB5h4VG
R3SMmq6Fe3f1dLLyFFOXfo8EOWlk5bqjE1Ih4c/mkEs6JuVku1T5f00eRQhwOXAM
IT6Q4CaVizB7S+eGzWoVrxBeT6/78caaN3Fl37DIvwIn+HZ+rWrA+mxRdUay6XdN
S/IEEQSMK4Gce4QQSupBtxxCqPwt5qvnB7rB2BLqC+9CVY/l3Z2qx+Huxoo2NOrj
+tTgWJeaIIimdmJZEAZVtbZy56hiTQeg93eI0QOy+rWhdprcLqTFOpJZunLIef2Q
oYZZ6337d6oN4favT5Kkwok8dgQo0hRezojR2j/gg2covVhBzrGn1Go4LXkOc/Gv
GRcaxnn1MFy4Ot4KP+BZnNfJ4gs4bRxO3Tqd2LzJYVzcw+lKyB01ioGrer5unpiJ
1HxpiRYpfJ0pkVruHQhqB873x44heQ6fiUiGjTsVRTq+xo4SpOwJCGzGlx4bC05j
uxnRxH3d4vNW3j860zyBDYeM5G0aRnGwMmvfYlIFVQpA+t7TBO9g9y4iu+HngUZ9
sm7OZnc/116H7g3WzPSFDon8Ql0Gh5BpuDCI6e+BmD4KkO7eVlkT9S/wdVJYy3P+
tKnV7gLo7khrUIfLtx/Eh0jJDj+OWHoNXQ5u8yjSYg3eUDj+4FlTx+aSpEocnBjh
dLWtRCrvfZiS/oTSF29hX6y3469VYkOqSI3BqTklYhgGmSIYgX+ZabejCfMurcW6
uaREFfJXHDYJO2sJLcUonu/5BYHQ2+jUYgroEp3kD2eCII1wui7uEaPGblnCUafg
AcHltILeoZATQ9DH/6sdGHkz0ewTkcMZHjvzGyJsZp0m7zMfgTT9KpJTp60ybzSR
D34zSrstxQFRDknof5ABPjxWPMEXwEPbdpFzU7xlaCddm2AVQISdSMp8gC6ACMyV
EY1XfMJk+1Y9SRxT68LpPkzbdFMaRfftqnDd6I2o+y3BbRSKCKD8nQGx2f4Tht8e
HGFd6fy5SAFmhp5IqeH+6Q6YYWIPG1/TpSSNOVn9iN7OcxR96svbL1/iqFEkct0m
YcGr9TdpJAtxVSuBtZvDNBsdRUSJSIBp0EqwNA6XG0Vq6tC8ZneIS9iKmlZcNFBA
Kt39xCckTZ2r3xbO1fKbiWNwP0QRyowE4s9Rw0/mr5vH39hOahHAXuNOvngi9Aub
os3QGablEEWMkX87Vscyqy/qjuelxvPYM/OhuhXPLf+HA39JGu9JOSufRsOg7/8J
dkTmLyEl8vTQ2LL90VVTjQtrkA6lLv6iq5RLNld5Hx3H6J9eCLFGT2T7B/uqhFOj
aobK+r9SFj3HKNsBIAa9OnyOOfeDTqis8U3NVrTLXadjRKnLsYgUU7w7nIS4eiIa
J1wXb1Kp5rOoTTmW3cQx+UuFLecRy5QpsXBlRbuq5cUwsuwyYJm6PwPCKMZ/eTcL
1meexIBX+C/w4zR2tQkz2IhbwZNEOfd8npuIRylR3/OPOjvJo3jg/jNYewfNKZ/v
JJkOin4dpsFtC9OC0CIxayRmhkslkkw24YZP4HZ6Ngq/Eo1IjM4Q/0pwQT9Ov2Er
tdUdWVf/Mv+KLboEknMFFq9MQr51KJliT2A1M7FDAysOTbmANYHAxnXGsbml+AOI
MzYdVVjgx4eWTtTJvkUHdvst9mA11dSb+fWmW8fGafbZC5JMcKrmloh2NJndITrA
x0XgQIPa4iFE+LA0QgFcBp3IVUPY/TivFgLuBaw6eHqSm7ZbWE11+P/382rdqPvA
vAW4P4OGnn8TNEzfyDKPkbbiZI4MbCrkpYYyzzwOi3QS9KbGMc1W+HE+uXHlhNLr
64Vv6iEyHijpzk8xDkK8Pzn+D0iv46gOC4zP+H2EtUZeC4Xi6rxUdBJFqGZfFFJQ
yP024E5LHhIdW22a1vSSQm2m1J3khHF37Wo3QMtDRKpQ3pEzaZcjOWJvBaQlNH9T
KA9Pr45ZbDEadjEWeVEK1usyDS3RMkGkNGxD7F9jcb4lcHafoEb3pQ5TRFpI54x1
W7MoWgdA+DvRzdyeHMf/YF+4DV5NSlsyP6CclIp2gQG+Dvbf6SUKu+t3/sHMQKrS
bzijVYlYusg2qbUPLsTKp6pDD1xHptetche75dXPVIs9g6aDHsO0F3uWYJIa+lJ9
XLN/QOTc9gJsqZIUDdqhaC6r+QtbwBp+tz9lyVjA1T+LqjoxCakU9NOHeAx6DcnI
xrQW4Q0isEgp1aVZW2ADDslxMLM/jlwhaUzXvviehANIMDwc+6ZdpcoDpah21d7x
SGz/zdjdOPgsO8xEFzClR8W3i3I3w/xRKzv0TjbrIr1Q78duuYHjPtbGlwygF5dr
dAGCQTbGMXQcTplYgQnECQXBLScV+FYrwCs1/pjIcj1eaG3mW0FsOztfCcWIUfFl
EaF7ETIihY4fQGyKuMdCtl2aprFSvZEMpVuJU5FvQQsUoC+FjbNYOMJPggI5+cLb
d3H+I+fZe7Be17cRBCJfRUWaH1xQW1vUPZ0DyfNcEUmZf/YXJ2Sh/3hG8hqK1NGD
0PQh+ayVc1r8iZAT5SUzYa0cnJYGPsWdSaaE5E3gzWKOMBtFFQQN2NiVD9OnVSJJ
FZ+uP7DPvEVE5OYDJyf/NVIFScFAwfYNe2a/89ecmqA3nwBMRwYI4wOZFoOlBVeO
TLtd6XVTsnuFr/fSbjuweZxYirpu8SzbnJLzTbRfhgGQ7JoLNF2/19FLSiBQZJ1u
FJSQKshgA5d01gmoPuYXg0lE9LItZsW+Lt25k8YU5/iay8/vjKJO4ZeTUN1hDSkl
cGPrSMbydzFyRlFd+MswE7Da2tp3aZQK4CDPmpdHyNVJBSL1iJH+0hOpRMVRLTem
Cc7O+C1YgXJV+YhtxyW+8Qr1lealmZ15d8zTKH6hneqSJuEsFuBdCiUU8xlXZArF
oD9yaXPED9qnkSJDSa1rPAZ3MjbzPKrUpfAaCX5Y89IsfSsmP9kkzl6UrwEhNBGn
VR5r1GPmS2ECoS9mSQdxtEvurrGHggczGKOoGIuEb2ReRosppaQ7AdwELDFZ6+8O
wz0rzkvwqJXXKDdvK1TKR1jL+H9DMbJ229HJoCRkK6DPcGAWEl6KIZuVqgUC9FNh
HmarAN9n9qBJRmtZbK7+pP3bfxdt8CLB2vba2l8O2y/zYFFT9WxUfkmHEmAuCqRz
VWFAIyT5NbgOs62OIYI6aa1xAMhNjr+oV4HihYdJBgVGOFv5kXchE3czjqmsK57S
GW8OmK09XlJZgA0gnPxhSjyHeBXYGDb/DCTY4a8R77Im7LHeEYCgn3m2C8zTfC+s
t60UZrLaoob4DzHCT2g/OAUs7J8kI3iirEhwvCdJgNIeoKiZp89rO15PFIlFRKJN
WnfHTjHWAC+6qaSmKHHrvcGadzcVukL+FfZgO7PMbfboCh4NCN9ekFGfzPo0l0GF
7CWHAGYWms8JreJCAR0LzvyRu5mh04wF20flEPoNzd8FvKVPUReFqQPBf1f9I1MF
tRpLFwUWoKHY4l5rP3wij5Q1bvC7Mhl+EQHMZzlm5VvZl0oB7NirUSR57kMG1GGM
pz7DBy04TBzVQTS2p7yW6oAXrARZuJ6X29Wlp0EAse1SQ0FSrPjjb3k+pg9Lf1MV
z6mCvELfFQ4xJt+pNxIl9aBKKwOA0kYOxKGpYGIUXS7NzijJ4coludODv1IJvC+o
w3SqpMMX0bUFpXfaTvbAV54ediyBscjLvk6YXRKK4agUoJOdfvkt73pIx4SNh5Ho
yWlum4uTUWKYEqu1O5JX0sO7bXP2ZNrf7m408xuZQLrvMFnil0iIgPV+SBPL6uWl
7Ur55Gy2BlG/REU9BGncq1dcr+Zcmd2KIM8avUKt/9LpjdXo+HGm7TvMlA/DO55v
3VNLyzzg5dBP2w+qIIVJ8/J1fK+GPupVMdRZ7W5WG1AGk2BYUVXUxcv7MwPVJ73a
RK2dVOHz63LAIQ/+3TRaskn9fhY8hu1Vq9GbISuiIDfRw5sBFKI8I7r/S1TWAMFu
uU3WZXcP1yyfoyFwcTQaDIFUIqjWeRcZYwqRt3hGRZC/epTooeYrtNKsxzQWOTaY
Xr7ger83Y0YaHjQul+stCKTJIrsuDDrQdsyaz9BfVXciAOK0PVkiA0PgtrcyJFOK
GGGhqKmXP0HBmd//JKzTWxXI+pVswgPg7WNr31+EBC9zzW/E2t/tU6vH5IbRFjuk
HEUxJYyLlB8+RI+v2o+gMPgLhFRtqaA1y6VhHcdVys9DdH9cycLW3t34MivV3PaA
/73C9LfxzAaj4P0k30BqsDXZ5v25qKTfpUNXXWV8bHBFdRSjYazEGOjqCiQzoXb5
dbjlldygeVLTB7ILUrSylhATmv7sHt4/jGTRAO6NyPIM8m8p1t3JFHEslnNlPbwC
iJeTFUH3/s1Dyu8FgegaeYO+OucKZC0rKHmrGZ4NcEnIeh7a96OzsIpFJPlw8Qvf
l1Y6CwmPsp4zJ7XVUSx0Zv16xLUVHtIma5WgALp9H6Zj9d450hta23jAmCyI+C4a
znfB7cwpPttGSX+StHKwLbw+tnQnnZu9ihmrlOl4a8FESkfGhLk/RGPa+6BQrL5m
dbJ3XTIDEVBIJhpDri5g6TSw5+1wXmBMBAo6bGSTCqW9QgA/IOWsfPWYIBSg4rSr
GqhCmMlBbTHDMMN5mWJC1LMGL4k3bt05v8Tx/TkD2WzMDZhH0SoVGVK7ZxsAJDN3
GfuQ8j4klvDhxaJ6xvUFYTHUKI3mXzcZ+up6FijIYg1kXZSZ8ssAvPkxG7609mqH
DfOHVvEulEYwcVj9Rn0NON0RBjpmQo4xxRCJn4hsAuGCLfhEKP4z0LPvpbgwZ2+z
csDW8rJ0bp/qCIIiYLTr1Ef+NWnbntK6PssGc7dJIoqA5x+S5Y+QLxk4FDVer7c5
eGgY17dI99IHFJFITd0OPm/6X1dng6Ljf2h0vUzxlyAz79cmL5PC31bgUK0ShUhe
a0ZJjqVPOJ9IJ64mMRYSxKV+aRUsxpeJupszfj+nSpwuHK5IvDf9O17sAXCuynOy
11Ie2+NWuhqLPnknfUyRENriKdWqoVVl8xO4IA0tuforbVeMyA4v5N2bExZc8rMz
qHcj3ufj4vSgKpC0kSHRKFXkbkoQLg1QAIzCaBeDKztq7D6svkbG5vvxXYZCUFEw
kOd7zCPEf/LGFxpDalpsgmdh6+7Jvc6bxN8cL0K6iqmRfYWgWAkjRVYp0GOEj4VP
fWr9iyMWYGpS7+yc7mHEhVqVkWOM0My8Ywl0PSyq41TstIJCGAGdqWvUpxW8cn1P
DibXf3A7oLsfa58YPYqxr3JBtEuhzTamMujSe4CPFwqZLMxpIpzncan+OKvKY0ed
tkMklgmnwArey3X9m5Oft/k4UMexI17lTGVKN0Jc7TCWctnEwJX11S8HLg4lWHY7
PLAt8sw46f/rxRYTMNc0f5oVo8gYTVRiVex2zoNO9hu2RsUe09hO7mTs69jew//n
jSUeRVCNRUvOKVh1ACzfDTXmuem1OE34iHqNsGr4cYyKAtr6YHbQGSIUFuxO0Rij
tpTrTACbHJ6IOwbte34vNQZ9LOvREUXDrTIA1/HEh+pHYOOBJ/sExtiweo1g4Ter
JqFoWBtXSu9miUW0IZJtQ2rNE7wQph5SrgWk/blaqwaUEYGVUpYg7NmjlBw7GnH8
97QxV6MwelEe6EGRw5xcrf4GvRFMDc5OWQLRgO+PRP0VNnwnM64r5KXXT9Jq0Rd6
8CQfwEznKJVK1Gvfv8mI7JtqhOXrzM1CY+oQ1t+Pk/SbJvLLhFk7grm0J8EDaFbK
SlmqLeKYRRrqqS9XV6CXWZqN6iiKdl4pGASv8Sut2uy8tGwo5osccnjP3uSLlQ58
l77oiDM0PME6JxAkYHWJFtQUvSkDdMBwKb8X8U07CikOYUC/X7MPS9pmx4RYh4c9
nJqkaPIDI7JQXMptZAk55rEN5Pp7DpYGU0pus46+W270m4ahJ66McFZeYSQSzOIz
xzERQdB5YIrsHz2O8D48a0ppte8Ivk13lX/S5aPpWrq0zm1B18FzfKFzSbShh7/w
Xayj29MQgDSdyJSA6zCxyR/5AGAfEetJTTznBMkXY8874KcNrt8zM2lX8CdPR9U5
oLOHEEKDnmA7Zdyl1n9ybTwO09mRPSits+hiQqVmvIIpWUVoidW6VJD/bbW7Vw+W
V4jv2eU3rxiDly0vkZt8FKFgLiJxrFhfp/iEwlAbLMW2GWC+Y5VrKcMzyKuOOvZ+
WQHugJ9THawCaWLf0sqiHaITeoeulAhv/Ug3LyxIFxIRZr+K7lWshUmnOn6RP4Qq
TtSjpeE/5plyVcfKFfr2sdiMdC6b5Yps54R8a2YboeP2rO7s5RbSDE+P5DNDdBt6
8CWJMCMnTBkg3GAjWuuD9MJ384Avxm58OuXP3PSD5tWLLKcjd0+nYwkengJr3kmp
14qP1HN+qxFNeGtbBey+WJi1yR5J/XGLmqUzpT6231u/OSFNfS8wljzBEuZmtufc
3VYi+LgYYgZClO63AWqJVIU/cgXSIwQruQWmGhh63wgJ7gVdv7pw3CllHidNA3h/
at/Z9GzTYLUI2q5Vz/WX5ovHTZ6wvOImfZXAN5jfP24M82mNjHZ+M+6APsxpBn07
PBr5eU3e7dEZ4oF0TcLt+zebfuXEvZr+wTyIDfXE+ryNVSL+BAI6LH+p0w43HVEx
Bc9g21ztsgTzlvnmjBZyxmJ9mhtD8VAW9/RVaR+wGCYAqiHpANtKPla89okKtK06
TNBLPm+onImcIBoIBFIJgfg8+1VAqdYj7QR5jHdfOHk/Twf04Ep0SOYw1n/shcXc
p5kjAUTlkrfUU/1lHo1n1Nr8h2j8P6L+FUpdEGrEY7iJ3slB+M6d4X9MJGFi4kFr
kJejc1oTXf0Zg2YhMY/zXcVy21/dN0pLJUTlol9aejT109TaseXUAfB1kcwghiqV
MIT2xx37k5g+6xiW3n7wVqddREM8fB/lFgaNz/D6DwsOPKZCSDseeoQVsDCe5nX4
RjUlKiSoKB9HB3zHXBxeDzMZYnuqNvrTz1n0K145PYAol3z75rSkO5latJQPtRdt
v8kmZ39IpJvU9xX6vY1XjXzWnjdDUX1JW5u/PLpSWd4RDNpcgXghA5RP3BmEDNEJ
DbmQYR1w2/ClfEzopNQTB97ox7lg8JwVJIwP7C3hRV+ojqbcJBO85m6R5qhBPCMw
UtEQgyV5l65KOBo/ydnjlK+LQpRZfy3BylW4XyXyQfdOZTHlNvAOQ6O2oDpqKBu3
tmlBM068ZPxVC7WfAlohFoHlqdhSjYOK4nI+cPAF0AoPMucXOWdTnPqiez38phtX
wwZaypFtZC+iQOWNvYidztWzQmIJxfioIeaPN38oo4zqLZr8QCLcNBFZYYTXFtgz
01WoEEAsZPsRkYm3V8gQY9/QnD7jfQuv96iV3UnhwThvrJUej9xw+Ok4P8k6mZTh
vRDqsjFMwKokRPVbEJWGSQnppYLHKXzkL9Y9vqDHaike1q6URKMgNrXzpuR1VGVu
/FgS/V7G1iKMOB1a4tDXvliFhB3DVm67DteyCzi+sxl5bi4TbNIPf7avD641gQgL
2gqCorsxrT0c+IEp3bR7viwJE9xcis+JXbsHaFL46+ixkgAzxv6/Hj2qK31wyqnj
RUNxCSeuPxRZEGbd/+QlzfgseV9RpUH+8IpV9MeYZMG0DNiDIeUUzIYAn959ZLou
i0qKHX5Ifmp1CfgLPBDX8ovTp94eWqQX03AELHJuYf8MabeK1wzIgKmZvJNnU1AX
HfoXqH8/XPq5Bhs0d4JO4fQih9aOLYmYVwr/CkmDQA4jfbS/4xhiOPh+1/ju0QZX
8DFYDXGt7BJhYuGHqp8Six4yZhD3sh3NlZ4g951Vtd3+8AuyabWO6yJ1v0c8TZtq
I392Z9fa+rT4/BJ0Vrfwf2tlq25gS8a2qDBrKbvcz/wTbDrvhobYmOKnSEDFIa5C
lIFQsGhrSHUFy5+FXvlK2P8bhXPfHLcld7PUEoStynMHeMBI/JH54vgQu3+AsGlk
eW6DDF1plSKTf1vdqtSePp8J5a+NgNT00AcUAw39yGwlCw8ICuwMaNfZqjfiiOY4
wqahAZqYTFdIRj9G+kik5fGG7fiA7lztngP6m8vKERG/6SHO3QaOYKPwOAayhRgl
/+N7xyM6BnSZgHDGNWPXJ3IEjVOfyBdzGBsaFOY0QafHhCVqrI/jGMMQvMTE5mlJ
zMjVi+xbfZgJwK2xocM0pl7HBwcHqyzLAcqPiHHOXWuG4o9XJ5V8jl9smHcmxGaT
z1sXDkL8NEwBOxbQqVkvf5QxVKFUbkUhO24UnstNSYqEuQG20sWqqbwiv/wucHf8
Aa/6Z6m6gMZyd6C94AwgU6Leu+0KyWnrhWtQZ3BKi0kG77/KzT3FFwi4onB8/s/a
EMhhZC4VvfwL7pO13j9zt0fSV2kfdfymWQEEBxHR0lHj4k9sE28ayiiDnAtvgghA
9lpQxhza7TkOiaD6Va+UWKPECi2DfHfTqgkhUT5HXxOsLBtuCeIjqP2jmoUiroMr
Ahfah7XNwHWuiMij8HGWIW32j887a49uQSneB+JvlU4RoD2p6I/GBfZ0TDosT9vc
LIkN6HaJAL08ARw0qnGeXStA5rEZ+khftRpRv6TCfiT6vjKQq25KLrHiJP8xtzio
wAGgCoOx5ovGFWbU1p6E2y5b371BrAo9SA2MjLhyuOJ7mJvD0R2DSl2sQMji2B5I
REmzLphoDxXavd97dgbskzoLrdhGZO2dMrQRvxD4qWnX9B6fvRuyFi99MmBzoyce
qv9dCuG0IX5gAMSmS6FOOrLJo5gNep9sHbqP2Xe0wraHzZ7tG8/NPB/+NazdAmC4
MapYUBpSc+WN2LucFkP19e6SCmW3yQeDmoyNgLesurIKqFdGplW/GkmnQ4ZC+Ezj
A52K0KKc2rQOt4bDBrEtpuSk6XmaH0YjkF715k2aINt20QYZ5H7+sQElLAb5Scb2
yDqiyBEuBlJ1k5TnWbjRhF0Td3e17iXfGrIlkz6NjPVBTsiLQqVhWcSXNDo5BkKv
5mgiR2jyL5/BV0CVJ9JvBXj7HOqfMQ/Pi8eudo6EOQ2/ftoTBZucicX6XcaWXfpZ
v2p6oXkfEpjhUYE6rYwczdeNtGUMKk1U0e5EXOdt7UiGq2LGajk7hjnmU7KdaDbj
1o6TY+vqqCkoiXpByUMdvVaBLk6lqytZ22Zg+xIAOra/uUBBgTa+Nfpk5fePKuwv
TBRb9BESFU70rZZbztfcOdpBQlw8qD3up+/fyB+lkPfBAHQg1X9qf3yNp98dkuNq
q2+HZVdXl3huOpiqy9Sv242NRk43NJfknXByWXN1FlEfpT2fyt7s1msR2HPr7Hod
QiBTqE/HszXiwywySVpiUf7lJ7vQFIghM1zC7jEnLwk9SWrCpLQrCQe0z1irW5DY
KsKYMECHYPSLsPh0P08n59v7bp8selZrmK4YeFz3MGJ8Yw9m7i9ECoPBqDDMOpZL
2uXc9lQVgLpOZYudSosQEXI35JaCCmHK+v9ZWey+2qKjVM9QcG5fLBl1R6o+bitM
2t0BDYtn8X+bpDJq/LU6BUY8tmOBumK/t+BTsM3JYaCvIisVp13tu/CNnyVBAxZJ
U8/C1CgCFgjiggYcEU4vJ3DPPICDdeQ8a2mqgfUBijlI5HC+fCKuJrPNQa8PrlyC
3jvR7L8gNrAFjXSea3N8NWTijXdugAcI5guZv7FDaLHoHvti9nI5P8MeQ6ymUdAG
cgC6W5fUuCOi3iFvRKDosygjdttHVskDEVi54IwemWbWxVF2RgkzTNi/iprF32uQ
8OQ6POBYdpyNy+2uRgzm+6heXBxwGWO7qZ3yQabnQ31MatQt4vq3i+bUZVI27cic
bV44O5omFziWQXweG3i8XkHa6R9EBedzVNEz0dNVNOrQSAC+MhDT0hreSjiDDOvE
+ubYivbMjnjQ1Sg7RC90UUsSAokCYFieY2VZWblb1cAuQriHYeaT+9trpsfAVt2E
myy+vJCec9K8UnpoOYknMXB1lyAK/G+9CiOYOUDhairDkH3l2f1Atbxd3D0H1ds6
Y/V3Gg+N+FWQ7Xzi+m0dAxpwpHlbEcNUMerK3dG0vPueVMmkfQ+G6WysXmpAkRoV
sAxYm/qF4M/B0kbMthtNpDR+necVaGYctEchFxjYdCSjdzR4KrFYwAcu6F3LNjrW
ET27Mx1jX/udZcex0hRXNOuytgCFoBdpudQOIDj+9LcxnBP+/8bh6+PxqTVQa+Jm
nujS2ZXxFf8nPOyQPUz0KUMa3ENK6oCILkZg+5Ool3cphOhX4cuwbQvfnDEZPA4s
5Zu96nmwyP+eFsKCOvdBQfsVHFRgi7yft4siKZrj8OnWpe2DsbArAE4evj41NUQl
g71Tsb5gNfYS03jnxc/AP887CfRb1V/nePhT3u6hsBh0App3DAzztohZ3ioMpmir
8OsGoh2ptML3FkLUbrIGg0eTQ3eUCrl1goHvztXwQPhAzjtZIk5qCmMR6ZhKS3DE
N9JqiWuOjAWEAfstq8/OV5xZM9gO8uOd4bHfEVJSlLGkhYqZjVC26SAC4qMRWkY9
L66AzFuX0ikcv6t/QxHfpmxbfhjZ7dpAb11PfuR2kKTzUtmOAKYzN3A456kDwZc6
Nfdi27tltkAC6zAdNhk+fnu23HjvXfu49N4PLOn91uBkOlKZRAudWpZmoIk3P8sx
I/vPrvddc14QtHW+9GJkFNWH966geabNo3Vvbp0SMJ3TAC0C8XhD3vVZYzW9s+NB
Y/I/v5e0APDauh5We2gf9YUBKh3qRlUJYB9FxoU8exuzuZxdPytl/UwJshhTZEu8
/JERTcZqJOmApZ0/QlfTOG2XGVoHzW5QSgDApZRkfLLac3Soavn77Hm+HA/0CXha
5yJSo3xobDvF+V04ByXQvXIUcBW0sBg29y8c4bjlEtcs4U9I7y7hM5a3StMHr8Il
em06r/jL7D9KnRnmnrflV8lS6dxYzY7tl2zgIuE6yDCFjsNCtA4zsSdylSaEAUPw
rjqvKL65RuyFHgbayVaGmwMt+JEQyzMs6kS3zKWQPUNkAr/26CNroo223WZsNnNO
y4K4iSAxOdwGooJ/hEs8qE9sejbVLq1m9Y6zHBosnl+URF5cFxtMxtu6q3noTyUm
q+uCokVANKWLP5YTJlGrgki95kK/ExQXJVG92LocaI50q21WmGC8FHtu7yoNTLUj
YsvT2kxlMS9iGau/AUWXxjCLO+Ek2iZ90qG7bboUANXDYlQxJt/K5AuD9jhRtr8R
8QK+Ibp3ZDd6CDBwqssIMCjP840KhLmjLuoINn3eFSKyWxjefrscQtSRkdUhgNut
Nh0mQ5FwZMk3cTPYiaNL0gDj7ueCDsTNCrsI5TKGi3LkWCsxDWEpENyzwkTSqmqX
T4wF5UAvY2IcHBrikbPm5yco8vvgoNmLoUw52YBDqQK5bH0NaHlba75M0ldcH/Na
eyZOg3wvRUuLHMpk0ysudhRvetDVm5hI5nNuCv6jo4XSOs+2cpg7rdHaojEc8cDj
oSC10h4FO1WN9ZSbt6PajFY13kapYsk4EZhkz4y3CSMnnwYUKb4ZaL4UV6k+Za0u
QriMWNmbBBm4F4T1Nv3mmcC34PAf6mnWQ9KTywhxNGs1Yn+R2a17fO//8ZET9pl6
jBY+LpItNbIm1Gcs6FxpADsZrCqSwZFD1yhrdpCK5kikRaR95u+/sON/N3bjuBeb
X6Gix5Ah4QnoJ0gTRA5siLp7GAFeerG/9EVtSLfPhhbkyXlLCAmCFY3jGE5VvoQc
f1RdfE+M4L0bKBCTNJpBlZs+OWqz7ASB9ViFNADBPhKO7QJEIwVmu7B1/glbK7sS
8AXhjRLH5mrI/OLOvIQi5hHFHpeI2CA71QyhO+NMUOjA0Py1iR9QAQ9seEaVhgTt
S7DKdeQNIVXcFx+ga69lDsnS8gbx1H4W3rqR0qu1H/sd8z79JRVfR2LX+Fqsk+6O
8eYWLYtWAsnYcYfbTfdYyy0+bbQpBZGJGde4USiprakD6uBBGUwITs3/LWbsTQWo
RAlU5A4bS4IXpADy+tVTPg83XwcCsM4og+05/fVF7+NC32+OSctHJ7JPpYDyparv
yT1I+EgH5PQ8sp9eou8b5HspRt2cfUFZ9HmVaHUJA0DyS8z0/GZbyOzeP2bqBb3X
0xkCIBKhoZZU/lHUqssClBEE7hZI8Z6BcQGhlDOCaT9JEwar2I0rEQDCBempsLmz
HxFi4A20CrgxMYl19XyeyHR4zHjf/8PgWlUvuOhmIQ+7UT0+SLmTnBt8bVfRpL+T
id20qJ02Gg84tFpD/WN/2dJlwgPZInaJrz+jNx5G0Cb5u86P6vpQ6XjdHDvaalmx
6qgUFKZO+fNjASWkoNYVNPA0sl0QA35OYR+YR7y3dq4meYs0Z+k+DafhN3IRk+6A
5TXGRzqOCTp3qumf1yCEpbdIpA49IEqfgL/N/owTWzcLB2cXix3gSACJQOnmaF4c
Dyg8x7BGjion8eqizVnvenAsMAGAP5nz2y5DHbZOFWhZh3GaaFwttJg0A25hJiFe
i0PSxTVwsrVd0yOZo5IrHolp/yEwNzUvGDThq6U7RCbzqL0HsJWQPqOIjjAL7ItT
mwH45CiAGKA0l2piJ5SwqlV+NAsZaexQ0HD7txWlYmgdRY+vK5tZ6pI2xKVcb4sA
ihYDHRDQjrAO/JoNKuW4G+JE80an7y0vmwWkv8gRPVxazZucbPDja9umUQ63yDrm
4aKiRWpvH3dk113gxu8xu4LBMN3bWgSVGZq2q/jrHFz0cqSgsD6w/BGHLYyqzVWv
VqhzoDDcy0U4zWYec6npmV6ADaTcY/eiXwf0cpJTUk1K21at5VkPn4SNE1b8uJ3s
z8vPGaUBBPGG2OmJEWsodBfvo79kqB94ALizG04623nGchRy89HUPcRkHMONnotc
rZfoyoM1pMng7NiTPc6wOHFC2w3jobSh3/1DNRjbFfRabzrnDOcCCxwNSeeh3xtF
era0TAantD2+lKdObDPiYomzyBydkzX7MxgslSyqsHLJYZEyXCl3m+SKx9ilsLPZ
MdFfwYYOV/40z99dLxNN3jeaPd1CnHkQeEOzQoII4u3fkrDh1lYNNlVMAb5h/mUi
4En04RfDvRP1zrRU+frdG0AxN9S1sN3jnjlUzs1H96ppe6YaV5f6X2afoJ4Wmdc5
7TwFKoAS/C1Fjk7Hzy60lJBqieAQ6e8IfhCO6It5pc6Mm9aYVEVjeH5H53A5+ENJ
9lY6icBNhN7oeeRdA2bCspbACl3dhm2ImhmVnpE/Iresy0e4LJoqx9667IT6rzg5
IGd5fkotJbRCTxR03XUdoVKGO5G3LNU65WCECS0chB0yY79J16zFlIvnz26QRIMo
YFNA8naS0HAAiLfPb5MT8QFpTcbx3F5BB9fRLn5UfpFieSnRARzzDnMY41yeTv+M
4bV6Z7N9okxn5neK51vnJiz0vDpNYroRjl+6WHB+HzM58T7KWYcF2wE0W8GtJQs0
M1BbZaB7pkiq3HxRxXrQTx/gqCSPanmYToub1CSq0mw6whNcs/j4rMpuAx7zjq2a
dNhEKGnkALjkZXA9Ibu2zWDk6KlMxLsSupHsrnYxuwT6c9gjpjLqD+yO1KFranfY
dYXfF4stZQ9F2Mdnw9TZU48Fb4/6gwRHS5RU/wMaEISVLTib+067FvJ89vh6HrzE
27/FXWRrX/ffy2e9pNLz78SToZbqT8CiB7LoM25OgCh9l//GLR/ObKoJq47vYvfo
hRiow+8Y195suxLjq3SA2JIxKwjJVEqZnmd45e/85cy9ADIX4SmPi/1+Ikd4Clit
yv9AiBT/b5qD/TJj3b75X4soP4RyD4dYz1htZfqUO8CjfKEmMhLSKq8M/lNNpECZ
AU0TA3mKzZINB45jVDNpwWnggdWbKafEcHyN6NZBkOU1gnZUQ8WaY+3/zlNLBFap
57+ILuDC47iwnJV5aAME2vIi93p0CNvsqgaGNd4gZGdk7FCQ39lJPzPdPcTL9OWR
OItUTPR2WF2vxmFjDbmMY5x7rG7rDGJnajmGA9Fmj4sK6pzqVaAYcZ8wk6Rg3gt0
luElyrAkh9Sb/EYVVCHYx9eRV0YhOZjijgj7iwDue6zM6xSvA04z3azWs9JzFHDx
PmBTF5jLdaneeJNowAtIN2hMJlTXEvGCHBfaghogoyKEleqaWp7/5vBAT6k0K6Ta
3tlmL+cPTJw1KS2vutK9/m9lAhbZXDSXmlAbWJuyseq4L26xJskuSI6+c/YsvTT0
yJSRF4h8fItwnrm+yUiW97rSLcccJAjt1Iv7lCPTtADCt16bLouFk0NsX1MdtWx8
SwnQi7CUgzqUvZsXh8FGECci6wtdkrFiM7M1KZXOX40WkXhl/siTcXDhHLqiws0s
nHGqrPK8Qjk6ebTYo2i42xc7mH0C/y767VqWhyWeKNVL0NS+SFp9DdAcXKXGvrlM
KVl7xDqkVSrHv2bXeIZ4ynrRo5WROO1b54J2i/9meX+Ky3HFMKRHUATHkP2XFLsb
vQS2T0xGpAf6o+9qXvWRHDd5GYBSOeVQuAJo3Jjoxa/wcsAndDnd8gvSGR/wUI85
eVM+DJZbemRAtv29UJ2W8BLr6oyS0twaf+ZHs9Xlk4nGBXpjO9ldqSjwWU0DF2LT
v/1Iwyc8yJXPwlCdoHRncD0fXIwvU6QlosXU5Nt1v4zEkZ4GFQiJR0nCt0lKrc6/
8WcGplAZ98ZmzEnA+5Z8i5H2ZhWcqr+uIFiazqw5zMKNMCSwoPi8XgkWUNuf8yJi
0KhagaRbacZmOXQr5j/J7PqGAmGyhI5S8Lj9H9/ua6qeaAOBl4uMMD4CtSREeAHL
d0yUQnrYnivugWRkZxT3QXPK23+IFaaBY9Lv0FEzop35kgxyiN37EyzEpiKTP5Nj
5UReUy0709sC6QrsYLx11rxAgBp2MADcYTKh52O/Z2uBonqMHnxq3FowajBbYsSS
sFoS8wVoWKtx8NvBS74wP+Lbjjr29l9JdfkHS0ncNwpy8GJYet1rHhUq7ZGa8CCW
8Mavu3Q+noRSpDsmhb0/zQ14nCfY8Sr+nJH04HuyaCAVgA69blW7AW7DevjiSs+y
nwLC6ny1SSD9NBliWtE0hzDU7LxHPz3+XdyoBNDNFIYE0be9U1VZ+bKKz9OB9wF3
4HGLvij93jKaFfXsNS90MgjHWl7mRuMDdAViyBXYnSwfe6e1bacnJI11Kg5fGpHT
GoMrzMxTNxQfupDzkd0+E08+vd+ez3/uFhpI7XaG2a2sAT9d4WzVTpjpsE9PuqVi
v8doLerEcdTiq9LPlX139eORO1CRPAzuokti6efJmSNDdK613JVl9P5xBYl603FS
Wvap1wfq5q6UktTN6WK5mm9pYC6UajQiUoMzWnOl3paIAN68kMZ99ItfrhMhxY0U
RC5bi/KCYrpB1QVVZJ+oJpHMdkaybK5T5MmgQSo/CzlB78Pp7BHTBbKPFin+/fwH
DG9b1K4zDzabyPyBSezeNqcXS7VlOKW71OODrEaaa1SCNmb49zxahnAHYLSQmCF6
FG2KmN4jrIa4YPN94fu1d73OjmjIkdmLXLD2YC8/6YjsirSVCk+hi6r0UoV+gbNo
yvcWAY6Uo5WwbIvreJr2jWUuGFvstW4FGK3NPNXvkzIzNkJOm2ny/0urQ3bYfu6h
uosUb1o71ihaABN+YDoKbvhX1oFgNoE58MoSm0VowLVfGTlLB6z+5M2RR8pY9wbv
KCuEHBUWzXfAXEUDMXEXUOMI+UsLugmUFBvp7Sn/upcIhdl1i5hE1z/6hc5TnKfl
jZoND7n2weF6O9bQqqw+OlG/S03MZiux0bwt6HxxYIEn6mhMfkYJ+cv0tyKRmkjp
bzZKkGHI+c6qnzLgIlIW8PI/rU2ybWur7vxue3muDkDZQU3FkY6732qwLXCWTkqz
08+ugA0iHw/SH2cHUV7cDUhrRrOG7TzhvZbVGqiO3xTLAhl/0XTA2aavIeagfsno
gYl+myL2HWkHheCyGMST0BfdjYgVcuKt5ohQ+vvjGvLEAVU6sUvEjUGRwBOi1Yrz
dMNHtlG0jhKT+cD29TEqDkuutCzBuJtboUe39lUGbLicqV33N114rMB0hh4n8WDn
uI80X1grE/MWQ/ZAXW9koLtq1x1wrgETaJcEdNy63BOxzidkV5y/3tbNzwXOQHNV
f/rCvDQfIfzvJjgkED6tjtHdcYx8TtUFiPF/zj4RNGHvXAKo9FZ/f4fusS8LBPPi
w+Vn5XuQgrD2ukuFIvcgCBg6ljO0eeeMfsvtJ8k1So2q22+1GgCx1oPmJPJAef5m
z5hlFEONH5m7Sdg3ttZD93/6xB4+QhW376GtjrxdzsL7CMqZz8Y1Px+oJ1bVi5Cn
TiRijwx2bydQXREIKkBrylCnRa50rW5tt2BbFuAwAU5Wu6eHgeNwL7Pl1yTrJjj2
fdzzCuRqet3NK6TS6FWTyCx6PxvidILkPzKMhUWWFfMF1mm+6EiOYptPdYxVRvFD
eFqye+nFEHOyqJUbPMZCO2maUCZxRmOkaNFAJJeiio6D7HmW7/dFeS867yRCmp66
vxj7aEYD/mHqJpcPDdWjBz07ryIz4OR2oLmYkHtvQVW6q384c+20kI5iR0sBg7mE
AitFZ1fW4kRPSgL6nGdTa2bXS43alEoSSsV3a+kTBL9o2qPs5NltUpz4SPPZYwH9
YxzxFeZU/iI4s+Y8c8RIIovJVK/bMlJamxg6mxhw/2TLNGAkxqk1DzCEAwwc2aGR
NIMd4bRPu7rFyQF0j/1kEI75SkpS/60ioo9gFK4JJwBC8Y+f+YFWCDCN3eWwo7AT
KB8/D3bKv7pCzGXku/lTUQFQza+nOWzPxLJtmnDHLIVE43zZ1ZzCjzGgnR7oBZ3v
JcKKpaK2fvma8CU1dokgAvT3FuhJhdZZwCbePrOY0C0cFZY8qKBGQB1Wu4piAbbb
uA61+tRhTX3zJ7NgIxGtL/2fi2eJof0rd+/52H778XR0ELxyUzLskw+lWsKG7JNR
5eKZxO/InL0BzurhQ2BQ5BECbewUbum99eLUmxupEfsCuE73WbQFn+xsY4ihRrq5
XkFAhHu6PvzmRpjWgLaDj/AChIMsXXT/Cx0W49CHOptOimcTkN9eZDVKV9RMoZv0
+2hEeRkfBqtUCkSjy5Avqpel8BpP2VT7Wl3zNtkYsbNZRfOLYPceCjKemOkGU1Fa
BFHvQJ6gIGOBhdsnkcT6ct6mFq+EGiiCPAcy7i0o8xUmMoPXZ8Hf+LkzMCzpWNyu
84gzLG8zwY6fpJpaSKr0gctYiFY9cM/j17otBFAEIpkPyKDE5NiKkzWMtbKOy1+y
9hwr97zOfa3c4fGlCrR/Nato1GRacajYjIWTbGQj+t/703JBbXEQydFLxhZSeDrr
phyeCezKdF6dU+VTjHnG8TQEtDOt9P9xm1p+ProoKchvJ4caipaJ8p5m/c54BGPA
wrU6Pzlxg4Thx7aWYW4OOVxuthpaGLOn8xsSrYm/KBb4YC9VjbrifC7A3ZaQRDnk
4BbY93il4D3zH5b5B19NBKeq7MDud1dXrabyGLtJO9maFGM2r104ZCTLEEUENQ4S
X2GyKmIfkmwV0kyCIhNX2hHOrgGwFHTtxhpMAA/MiazACu+8wYLVj1brW2q1SbGS
heVUodRln2As0wikpYdYrUUvYRgB8kCmpHmqtnc8Y9Bb9MSunyUCQnwZ6tJzSso+
Wbku+fg7SxFFWpYtl0vsFN4x0m97dfDm4gBmbPhaOtimpkOwfoY71hT+gylwggQi
FW/wdTjkZsXzFxZQPQqquQRslUao8wNuUTtybSoCc3NKkMwo4Xggj8s2pK4BiRyz
Sl0TcDnCsF6AAlTg5OWQRnekjgu5+3uuLTjTYKajXXGDVXD1YTZS+x9UkgUTGQyf
yToUvgr+p7q4HI7peQOKyX7svyIUHkYvHDL/ooastm67o+l2KE6woycJVJJO35BU
aE0JYTSUPmNk7HofCFLYhHp2dVM7WV7GPRdwcyqX9lYxxfaFzjcQrAPIk1GU1AAT
OuFw6+IcdYc0fFFyQCdK1asKg0ZfuU27pYm2XZgG2zvKmJgRjgiyL5/5+8RmQH0J
XdmgLu2rxbAllCgYV89P3iHgQA2cjXIXQT3N06WlNHsSLY7jqtkLcBYihjB2zFDp
ciSTbEwu0Un7BNY9LbuV6Vy5X6M5RwM+TQOK5icGMTlE74MrJisbszcwMYEohbi4
YoWodqmdgeJh3w+c9Gqw7NM7WUcwitcpKELmvaoNB7yHyl+vl+pDWePshFI2YSlG
cxZMoRNfB333dLolaZ5MYyVz0iVIPl8efUpuPxWfnDYN2eZftX4UZvDqM+d39Thv
o9oqD0rGyGBE7FQkIn/lPC6KQnRkXek+KJ9jI8RKA3G5lySS6CiRprVvQJqB1nGM
O6QgCAMdLP3ty3GejYxrr+HZl+Ef3oe2GY8+uBjsS0H6v2w/tD94Dzb8ZmngT9oM
uL3M8adlFjvtTVOLiPCps5Kp7Q80aHCZafG94Ld7M5CjmzFNbOwLpAKetku7LodJ
J9ws7Rnm2QNUjvxgfBcCiM0t5PnFIlbfm/e6jlvlbmc9PVj+U1DsecRJxXMRU7D0
AnnIt9p3AWscx78nOS0ypy4xTtTEAUaeTrPOykr6kjrTkcSpI33O+EiAlaEXpYzC
D8LGKt7JtDPJn9AKAJSSw1fr1qAo38nUGHA9rBJYLvVRFo5p0S73F2xRTeu1+bda
eHrFnN29qcHcUibiJ8yNe75FjahxMYInLcHa3btsWbBppXBPFPGp4hUb5fk190KK
oNpo7D8iW9IkMYiGYWyEfX1iCtrd7j796WE8NGiCGBajce7e60CoHv1xHAtzDcP4
zeiin9CNlea1mhxBeH1VveZzZgFZsvpXTF9ym0SQGdio+cO+qDr9vR9rTKsxeWUu
B3KL07/KpV1EX78nX17IbYzXL54p/yc813Y9mGgkaFUz/Mk6rZRbDwUTHK+iewde
RM11dKYYyCaCv0XdLXG6bzvTPWdEwuXvWHzMY0zy/k5TUEGVicFtnoJI2RT3NZ/z
WFCfwyKlC+H5ZEiODzy6KiwCe9V+37Gcw6SbmwFnvrVWQcxm1wv7R9FX+Fxzprxg
+C27taZiaXfaqiXuI510mFh2CKmZh/VXlo2dg1a9YnNQR8ZExnhaC7CsYVgKDUgo
2VlxoRM1dQlvzXcUlxmJJzjVIMKSIncqfKSJDciz5w+jrk18oG0kscE6rCA8D5Z2
HwUA0QZMvOS/QjigEFZKkNFK9DSwiQu4tCLtlJX2OU+dVx9PfHc2NhCch6EV4Ywe
xtFpqhXdaFwQSTvbBDL6ClfaHWeOwpioyJB9SuZiAQBdspbsjQyV8VXFpooLR3pn
NCXZeiT0Qr+Izsv2R4ALNizyjhrYj4fkuhWwdbXq10XOLVB8XHtXvusRVZQaQiMm
AnRxJ4CTMBv6eQkjHB0YlntX5juBT2vMobhs1+jTwCLcs3Lxxb6Gh7FLHrg5fLvZ
88XtS5to8dFcCiZatg/iIRQ5M2VZx0u9q5juBNezJFp3y4quDGZY8P1Omxs6ilKS
N6yk07zjPRtk6RoMZvdwN00rdtzGr0QwLxO9DydofitFyoMdm6GvU9GYvd2tPWvo
OnpP+mngzLQNVgkwKlUYsvt/17sH7LBZ7SgGnVKfRyWxlVtk8v1T/JqHwcp/MQqe
sP3ObFmiR8s4JYV/04BC+eqLG3mCg6vLvR8fnfWCuVCSWGMZ13PhyEMFdSew9TgV
RjPU23iqhg2doBya48CRQhfKQfDx8xQanm4l4N1M9Lfxo8VHUPBNJExj2TqKbfRm
dUnhOhM6+gYxLite3EK7G61HNZBWQY01t7+Svzxh68VmQSRMOLeE5ASftGPiBgOs
wXtGKQZ+XoXyTgdPydPPrISzsDJ8O7FpM9i0z1GP2zPngihO+K2utS1mQdAkIuSB
L9H7Ob5qr7Q1wVXxsvNxwf4DtyiU/1FYnvQABGYIl576Bnw5FxwuJxtrM+crFQsG
l6E4ouJskoztwgWFXEg+GVlvjRni2BdFaONyilcq+32ek0VR04HJgZlKpxj2uEB6
cbUupMteoAMXfoZ/ra/3eLAVUUQ1l6Rah5fiR5ri8LXN2Rms8bDoKlrvP/UPw0et
fLAKdwFZ07du1bo7KJGJzeR/PHpDD9RmsHimNQzG8aulC4Or75RaTeIL5XaNFYO8
R19USdp/u7JOzQn8f9WyxUvhHk/Q4KZPifeXJM+ZfgR8rXPdjiKv8LzKQcL+OLmq
f5sQGZuoSVJ/0ydxf1q6RH6dY4eFp6swNAiDC/D/T4DN9usaw5ZcM21KA1j15dZT
hJJI6O6nXRVXP/jz3Ii8MRdrMPomny/31lZxrC7PAxecwM477lngkSykM/CLDuwn
LjIV7pUkUJWQ+vBCaA/s7noinBFhkxyn+Qiomcre64JZqj8912Pe1+Dwu0BW0fme
aAWeEgRSeR4NIUT515b+tb67NjRGYUlStdoI7/3UoFSsb/CPDjQkSoSBqPHRdEJn
1HXn6QIu1s+zesPO+/NplaZfCJWcaYHzxBH5N2gF1rt2+h4cgT1RvhpV813/aO2Y
sIn2WiY8OK+2wAuF1tdnIA2OS7b/jje7sM4jZqUcPZr6wY1EnYpC40mRmdy7OdoL
Fc0L4/JZbHXBOmUxO2lvyXKto0c5e/2MeYBlQ6UV6yrUsVht5mt5ntcfhzCjL+6C
G9oIwzvE8QXig5jKfv0C4UZ9X4DiADuE8uuD+Pw0x9ryAPYmYgJvYaUuJtCXrj7b
ayneUU6YVVJzk4zHYrmsUASUiJFRNqaz0PIk60YEguC3kxVeaqpynAy4UmPNhZtR
3Nl5+XUnz5Wb9FiUNBsrTp4t0PRS63etgAUwZtoqiw7YQa0znah1dZYOhkNN0rNt
DujDBGO0SD3DkreJxH1xDIPjWtbxtmRiEXPJosRZf7UFpJHkUyhiLeIKgn66A81W
QfwUIs1BzQUjL0LdpEXMB5bkxCc55FsW1T5H2yM7zkVJ7M6D8fOF1gkEhCE7IkJt
LtwPnOvu3d7rWrLVij42/vlVvs3kSTAbwfbqT1xLfgj/o5FVRFBgxA85SGtvriw+
Wi1z+NhRDqYKQlcHg0QlK4b9U+/Eiqpk6XdlsxPVH210tHFuLfqDVpNs+Yg5EuR8
kHboh99KbX+tgLd48WOSy4GWDLDczeTkDdWV/GbP9XqBEB5Vi+U1GrE3CFNWeTiZ
tvBsYPCmrkP9j+tH5z2xcZ+hbyoTz/pHF53/kSrGKVD4yfF3aLcoK7qb0yTpu4Mu
TFLQPs0StNIToSFHOWWuqi9xGiBOip8Ltgh8ZE8h4nst1FkFI5pC2TuDpVXvLRfe
7tNqhEhZmWmEhRbZzWP5Iwj8OAEHlgTroa8apuqxtId2BN4qzuAFbQYMbX5hWv6j
zn6Ydmb0QsmBLeC6V/0ipRVWJ0bwjKKV6XtXh1XkxFqKSNeMoKoQDRdMZZMvh0Lq
Tq/MUUhU+J+MHc5hYO6Cg0Vu027MJTRW3zM3aXry6P0fiFVMD4yAZXirNTL0nqSc
1eQGjmld1heBlhIj8lQaqKDYraQ8c5LeFbURtybKcoIqV+aa8AqVaxUqAdOhK0CH
az7KbVClJt17rdezAlro+WV3BMXgJyWGQ5hvi/EDtBnUGE3GuCUpCUOqveZT8BfT
uddN9vtsJjkDu4hlyifCjkD4FmZXjkUJZ9SEmhwwZitKIMAIvhwf4YSc4nzqOl3E
3FTqHeoTipIEFc7JuP+MRpzvAOHshkIzfmGHGh/eFtCm1T56LAP4IsMHtxmrFLwq
lmXNugtKCYpw+Ri8oRQDUHBbuQMLAa+K/SXqt6VUwYRDYuJZUUCioMzttAhom/nf
lNJ/pT0IhaoIh4JttPyXRlXHBk82itc60Az+vdUKLh4eEHWP4r6eW/3KbmbcIkzP
Udrz1WRi9XjyZ1shcNTpMefH60N8SYRW/fAnic0CkfmFSNE30AmX74RGsCTi/xnf
9DLirL0OqMtem4wUKLakXUOmW3W7YJX59I0b7MYl9MoKjS5EkLWPG1LeX8g0cr2m
Oa5KfoWlc7+y9iYiOQ9ZYLnhe7HdnYt9i78xuO0QHnUJGgtNH45wtfdHdAMT8A54
uitjS6s+oN9iiIo9u2kRKjJysBZxUDDHA+Q7ObkSLMOeDrL8u4NhjPec6F1atKmZ
gFn5wSCgsp/ZwJo+Axg7AiSn0RWF7RaxmgucNAJX+dfITxGIoYHHnaHvmnZBLFmr
bD32Z7L6Pm5gUgvufKPiJJCRz3VjwR0s49A9eFYbVy6WLaSTsurnbREN5jxO633T
Eoy0+qobvBp0/pesOpHvbpn/MisD9Nnb92dqCbB4Yk0AU4Pw84nJUb8+ECV6Ffp8
wD1T5Fo0QL6YIJR0+MbKgmYxBRM+WpthPhdg07VjvYa6RQUxnAHu8XgTiWOpw0vN
dHXqpsQ5a1N2S6kugr1g1mKMPLtYQn/QLke22uACQYvwERF1ep1i/kADlLNrAg10
SDh0sCuDnGDDpcZ+1zslscirIPaZ3oNy6f/W/HSXAkW2Ca7s0Ilztsrgpxx+J/bu
wAZDi3hVre06nHg9DzQtCKsRx0wq7KZJr5G7GbFIGQLIEnujl1NKdyyMHftRITT5
tMPk/QwVqy7r9RltvH51cJrdaCkiAgN9fIFwatRflXYB9D6P06rLTS9FT5Pz3Tv/
+PGg4zE1qCPNa+5KCmEg1VDO4yTvYP7TkKfGx/S8yhUAd47spcgZMD/ne4Nv9eUI
2C7SUQcoQlGkJeWKNo2MST6Y3mbwoaTZ2zl1Zmipz1HqkF2O//vqTOKqOlGRZrLC
/TPCAqIFImM30gG4koOq7y7IS3EzG5IInFtcu/mfwb9DRGuSqa9frsS1TO21UllZ
ow2QXKFuTrdFD2OTXIoK/+BLlR6SvCjPHn2l/arX/SXLTnyHSayvlk6RO8GfZZ9M
jtGMwng8SGiKQ2Gphn3VWLaXqEnYLbHhVQysz8o+wPqtnh9UVchC5AjbBi/axjmP
Nk2pxGdiiBQIDln/jV8Mr3Km0kPnfS/Wn58pktZCU/5XGLzsKSMBFVGFS+i34ysv
Hn5YozM8H9zA+i7e9/vD7Cw7lQh36wMyHTb0sz87k/PlPuyMsQxKpWfu/7QLwKX+
2x9MJJ/bXIpcHqICS7WJiLxzwfgs7rCMXFF0V7Se8Xd6LHQt87+ITCoo0Ac90/zF
HYBmEu7zfJcxlSwUqSUdoY1cJGIoBNUh1QlNtdg4vcUlqk2vmi3CG9i30GDDdtsy
LVWN4ZlXush67w5HSWIyp+Rxz8UHtwsCQPSiuQ7OZ2+sIG7gLxJAQBSf8jofoWVx
Po8qLyeRCHVsfguFDviVoyJX5JLPVpAU5mdDArFh6q0h1fRCVPAEvJdzwhZwP2v5
ktmWjn9J2R2dfO8Oa6ROxI0CLAs6jIWbXTQyBn9b/MvF2iIYaPCUixfP4F+6M5ju
kbhSuKdx377or5MN4y6N7TXVVlEKVqV8bR9c9QTk/l7yzjuq0kpqc2KSCwq6QsyO
w7d4a23nsApnhnrmRsVjpD0MzUhzubBehmFfTF1hw7eiyE/tzUEBp7OEEhdu1H86
9pkjhDZj4wXYfXIQh6fqPpJaVcyAvn50ir9a4mK9cg/StuI8+/Mih/k48KHZdjBf
fH5cNVb9wS3q+EOi24sWcm8L5fGDWGts9h7d907UlNRQTm5l0CTWzH74+t6tKS1I
ZuC0Sw4tZy11f3Lyu/BiHUc6Uo5GfTWi0dUo74aPllx+YDQMOdxNPRERbvAUX/VD
KDQPWAiGxCHFQ1yHTv4fuK80EM8eIRRkzMObAeSa6KQcUcI+Iv7vz9aHYmstIrm2
aCNlKUxXzAloNtKB+3X8c6C2PK6VpqX7UEpfMe1jtCMesZjyKoCYoA+ZcwQ1Bh8k
jFo92yUlqHSoQ3PW8ITlaQXQfFgdlrJrX9Ox1UOXx6p2z9ZdglWXx0Thcw+NM+G3
en5kw49ILoq7UzDT1TSR+DXMBDiB6eZTOWM79VAYe+wQVXkUokmOGIP6xhnPUtpu
i9o3XL5OLC0OKbuZfxWRdv811Pqp7QlNCjc9jt2O22j9M01l+lMlpeZmZ7ZmZnY/
ZTdB05nTKTPbiPcGdj7dbtsDZ5rpp5t7kMndQVJOGzZWzJANU8GR3TjJXyTJqbu2
oS/75dtxlBNf4Q50Qt+oWacjUfygiLgltVXTtUp4eiyWwN8A8kcl9oRm1T476r8U
Ug/GRFMVOah3SS4WLCGNJCLKwdiJgx80lxApeiGFIgMKKa3fVQX1wnvo+V8DVM1l
7D5zuoEuqxFd2sfzNYE6JSNAvVTBBtvRtCJIkJ/HJJvUs9hSTxRwInos60ZEnRZx
X1yXnF7bXw/cbzLsQZiXZvRE+I6RrngA+LobJujfocy3gATqd8LpCY/G6I5eRzhn
damJJHnknokekH1KnOrzQkY9ZbQ9ttkvuYBh1Vl7YG/sLhH+1cr9L5KNDBctwC2i
WnX5HruvFb/XPvIp7F5Aw/79zbLET1YS2GERb6u4eYMME9MXPJWmHrx+smZDB8iI
eN7gyRUbsojx5v7osglsh1rdKElG8G2U/p/b0Vl+bDtk7Ag38S5HhSUupMeBxyx/
X5jwjIku57GpGTfkkhkZgf1o8b5ruGusR55B67gZNb9KcB4GNJ6rdmh1tJzsqhT1
pIA9a/ELDdVVlPVL8yI7YWlsRTksNRL/M1R8enzqsjZPWzY54lSV9N8MmhYEZwLl
lBzkT+q4yTyN+g7zCfm+JPu8iBvG7KiY/P/7McpiXian2fqitGH8T/he7IuQouUK
h+rafrfTCDQFEIMl5iXMK012Lf4sKP3sqztwj6MJopHn2x3beeAAyDDy6kSU7+A+
HQXS5NZzIaIEJraUlHc/zzLV0sh9mt/LZwd0nJD4RMzZKr0Egy0gtmRJ3iFWB4sh
WYYuGlblijniA4aOHVDfzh121DKEdUm7iQxbMk6CQC4K/ase5eZu6R5NSh8dpmQJ
qZLEYVd1wyzLEsHzpumv0IWxt5T7UIKbWsMsXT9HCXahVIJ6aNtXd8sIiwg9oWKo
8TDHXAI1szEZDxr63MyIaYav7Gd0w1iU+LoBrD8NnKQ9m8aBGduegmTD34ygb76P
g164fWHS66quKP9oG7f4CCD6/fA05340EDk0cIvCM9ByhquOTYTOuR+d2RtGG0k2
ySDakEuHQOZcI9SKrgb0IGAbM/GraTQ68YLucQgya9YECy+KY0rHLAzjztk1meTp
Svvy+17NT/5PuCNZvQ4ZJxXaH8H2ybZ+Eq7n3A1tFbrbwAjTbks34cHj0PC7MUwo
4cv2kPkY+tt/OmSch2IuhnSD2md4om8zI0VSDSFAJAehXcWUnTVdSooP0HOwAiFo
4DSOWHNt6h3igkrQ/2GtNLF3dxlgjYZZnvBUUMzqUKX6QS1Vgcq39/aFSQlLyohy
SDAblFGua/YTEBiBVzjL+AP5pZOKuX4R4td9kAjsYyNhtDFmIz0XsynxvDqVUnhz
R6u+kRFRynFZ6MfHyA66K2n0KCI2JHeOR4u6AfVYolO99Ncc8wBwxwHDJXDp0oeS
A3I1G9s5Ovs9iIQI+HVes6ZeIfC3nbEePLdG7h9wG3D/sWXGlzJAVbqxessWMyNL
vlMobAkfZw2s2B6QEyMlZBbbm6cwI9gW2uokGbtc0+7wof5FFPZ/v5xUaf/N7FQm
vfsnmSeyUKqKCQ/+xP1kOR8e5vqfGy9IXCzGoqP97C1Te502hrAnZtIOzzqeLt//
/r2PFspOTwHuQq6ZKPSVRnlDzoBf2ZdzBqwOrsKMvlyI2SPgixVPs8/yEiTSo1Lv
RTJvuMUiz6v86/3XItbb6rUPLp0QqMppP4f/a6gfw0+uxsF6kiZs9Ku3JxEvzcd5
0ZyQ50yi9J7JzxAj+jSVTAYkzXZ0B7IBUlPmMLKP42X5elcPyirjA6fCOIHtNbBs
AaQ2lA9qydRu9AIvGXVdZ6VvFqCTbXHJoxqTVh9sld+FPM4f6s7/yeDs3AT1Ordj
W1Jkh3cs0g1ZGPCovNlemN8nA8yPxzNacvCeMY3+Ci42ZaPC263ILbuP/I972E9s
LNK4WyPpYQZcEFGEDsIoajxN0GFg4si+J8LSveYdVGJWOZLAsHbx78tRQrNxwuhH
TiyM7fada7VZMsJEGZbQ4j6qO0rhakPxFhnda9vqS5A9wRR39Fkimw2nmphmoGoJ
0xWPIljoCalMXLi2d9vVrNzU2olmj3I72QoO7Mie98gHF1WEySZu4ml387E0Np7M
unXVdy/2Kab+bIt4aIRU6qZf9veKg+xGMBKQh0I5ziORdaFUrJnAkAOtjvna6FpQ
OUDy42Aqr+fcEWyVdRnzQw3JOrCERDBPFjNQh8RpneqA7LTMiyg+SxpnVWk9jLU/
5A7cUi0dnH+vD8Z+Q22pF824LOQSwgig6QWbvwE2WrEUnpCEF5AfyLF7twE3zTdI
x7fqRVbUTuM49K9AZEFeODblE12SRWEvAwNqvbJ1ThaumYBE97J6r+5kdMz7Jc7P
+4ZgqMXXfUbRADSKTwX1jveCtKxTzF/zaxSh8gU2SRFUT0ye1BTWrH6KNOjFPiZ6
7b6ASrqJ5OQ1dkOsdeeHsrpPGvtNoYUGRGdNQUD86VEzDA4ONY4NtkY+C+CnRRbc
RTwLezolNRtLMTtymBMMiZNe5jV9e8pIlbaInucQPMWA++k6sL6q2K5M/uShMrzR
/YKvcf9qCj76GsEIfrkuz6Asmg8fOIJo5hwjEYI+kPZuT/jyXvltxI559Qc30cxi
SCo57Qc9i84Qh6y255APE1A2LKfhGi+YKupK7kXGfCY4NFmw0rZR1yHAQtzgxQVX
tnSOxYWCTjPUrkcvrmU1eAbluue0kpIRkLJJgNW40YGh+m2kaSBtm+X/N90X6NEY
MnkahYrJKXr4/5tD8U0GgftSZujIFANGNbgcUtPh7az6QiWlzTAnuxCCwS4kDpy2
+dQDzPUhz7oFmMwWSc+SJCGFgl9A8ceAbGA9fQ24FZvafzPwRk3Ok6HQrhLAi67L
AfJkNq+EAn55nwW/8mj9c//bn3V9NZBh8rRzgfLUbM/NZ5HUG/9pvsx3QkCCdVtn
SiZc4n+TrP6CaESecA9U4/qXb3RPlE5NrkZtxm6Hw9NqyedeY77640NaSNf0L0OP
wkXB9O5LW2JppD64l6tT/v30ht813YThgZtoMeD5OUFHn9opBuI2AvGKplKD1fAz
XXz/mcsBcFNmop/kXKxGpil4MvHuCLKvy6H1T0ztAiPUQOf745yQQZcAh935jtnD
a/u6498fN62RAPCehx1JpnIvfjlNQbJM3B0bV3TKX4EEfB57KZhf3JG8mdiU8owo
KI/1eTFz+UKptds3FndaAXjO2d6LEHVxLJotZ/4lWNbsT1eHztKNgmoSdsUsYaoz
hI0D6vXMmoD6S8wh1lxRYB0bFSCwvWVEe4uGegWO6GVbNoBRpFynbFvsyTBZBMkN
sEXZpSD57YNaPOaf2v1mcVUHpzOE947n2SRzwY3kyUzvP67w5ijVhxPlg/iLyqB9
vRSBSBpDwYgY7ADus893nhtvw3nKa1zgUhPcvsOnFxY5Z+i5ZcHLx0RPXVAVOjeW
MX0yb4SozBIu1O16cj8D0+u5QvyA+cZ9olKOmmRcBYMLmiwSnpDpcMnAHto2XmuA
w/NHi/6gHBqsMpqECBRROvXFb9Cc6swafwNIIwBhl3EX/R2CjhBcv9zShDSbnGrL
vvQZn17hthfUEroPzs561TlpMAlpsDwxFk+8mSAaErBts5NOaAIImJA+ByNYR5re
q/ApSjsEdqtYKl+nRhhNqRaqF4Rlzopf3D1uI7DPhkh8cO7Bs3HkFJCbWGbzbPd9
ITnRSQ8pl0pjfSV0vgswTjPwD6PJh36zZA61c/gNLOdJ9yIPiUFWM3klTKNRK+IS
OXM+LHNTE88Fbi7tVRnNeO7E0HD8q5DdfkBs98wAzxmd1WyrdFYzLchd5S3mk2Ii
dR1G+Ms/JQa5ugQ3yerRtgf9iNIaHfm1DYMpVpGCAbt1+EYkRAXKxB0b7sxTa2mS
Pu0U4aXEp91Gd58zt32Rb52xwKkQu9kvbkv2Rg8xpfT/P+Wv5H10AlT7WnKfE+Kb
pRV59aizqoiZFMErg3Dg3YKZpt4x7j1F4a0DWjnjOdswY1l16YKIbnPJqH3HSUQ7
OA7AvpgywWB223sKvazFvt6yDD3edYeSqJTZMV7o9W6ldpqELQzOu9PEqahFc31F
71l9ft4FhNc/JPyGFuJAz332Ib4xP1YV9wlubZyE//rQ8D5zstXlkVhymlpKPtwV
28FxG5noyjkbiepI2wVekueRX5CkLaT1HxFZEFwMnjDywwdk7ERnf9VBfBvklJYS
3isyi09AY/isThODUvKkeZXj/2zondq7cd0wG4Dhfe/HP2jgVQrJOJ+Ozgz7x88D
0Z6vsYzVd4m1gAn5Q0YIxuZBFa5OB+RDasP3vkpV7ewl6EBJGcGPcdmtD77FEh18
QTQVXDcqfcxCvoikCqaftuN91j2lQ9OlNoedr14Ea6Bmc4xxnhVgTr2eVmYYscge
C0oQB77wShrB0XHQjBAGuy/YZxwGx2XAdsJRu3TvDbePafxiRysAbjJh+Y52l/jz
i+uVLVZdN9xXCHPlbxsdnCn5dxKilBVOoIWFKT4HRpERS6SsW27EoFrRet0bP4zv
7wcv04/dk4y1/Q5HCGDmvFZqNxNteHxXaq/NgN8MpYL/LNDAj7tAcNASMk1fgOI1
okRsYhWY5BEbpC7kYvna9wXk+PTSyIkQ/m/xruX5MfchNmIFrnr4vzqkERdmGo+J
bgAiV7aYFN+5ygsiIefIwqpRphx76pSZhZyIa5u0RYlb+EM7PNOfnp4jTNz3eBTA
pd679ulPUzCwzh7QsxUbewAKSu88pF4yxmRcE5jsxypOQcf11gJrVTvTjlluPrs+
/Bi4n7oxv8R2lac0v2ZWO+zOpG9hASEFm/aj4cUkR6uiOxA+n/0/F1h+eK4h4NvT
S9hTzCAWug76czsIADA32X1ilCUl+gSPu5RIEGkw0X6Dd7fy8sMGkpsVSbOfwYlw
EvWQ4aRzv+CYDmQh0p/CKff3QB5i1GrAdeoHsVChn+ge2QGLTY1OvRlDd/AC3rrS
8yTQXHloKjGMUAqoof+eLgdhrRpyr607x20reLcVEo/R/6tQfEIVhxG7zC+1QKPR
6sZYSXeT3VgOcQypH5+5fxI4ELtM/CyQB4CpKUafiNZSO8GmqqIT34HBNi2l75O4
xPVoMovON10nTQr4IfHwl9EQRZZKLVoUJBckKNbLIL3YLdjyHSN+UawfQEjR1sJV
uTFezSJ9hU8YoBMnrr3hWC/6sGqn6SQuUMxAgBW3j8ACVyc/VRDsMoc9JUREXTqa
UjnZYjA7WsPWBZElzSHrGW+fN1jiTaZkuLAavxOdQA11/gMmzQ+6P7xLrCu7xEgD
xGM9Y/LWRhDz5cVe73KebUAxyhWco4tzb8an9orTF+6Z/+q1eHIN+tVkFi+7XW5t
l6mLZkyEdgCkIFQRmOSDv9tK7uzxRVxin/VHu9PxVKDZfi2hSKPkzGQ7e0YCNkt9
Q9yDRwhAiXIkRnVYUHr/cDipCa/Cst9Cjj6keRXK9opOlyeBF2Tiiecgaug6HWqh
c6PFMCQMPiVIIUQ7WhH//yH9Yy7cLXFOCICH2J08bKMEMWO5+shm3FTQtipuQGCZ
b8u0zZnMKVKEEZGojZHJSQuHzsE3/iix+6IinCUWfQ4gxJvsHLl2XcVC6/5+cisz
Ev1qch2JQYuXx3iJpxlwfB4oTEeS+vmNipoHuUK7VgCYubTvbuikYowmjtqiceBD
bbvZ40FTI2LhOHAFRGJfEKqLgOI8/8434Yaw8H7GXk1Syer0BmFSYDl+4beOkyy2
JdZ9fqix0JQUneM7dl2brcgPfuJZhbXBHZfsdr4/Z8IlpkJgOafXYYFNPvXiMink
sVj8gpXCe26Vu3DUvkU8W62sPMs19eJuJ8dW9FNzmsQhGqkeXD1m64k5u5co2GWE
z3AC2tMbOyoROgyWNbogImKkvSdK3hA3KRBgqxPldy83uW7xwEG+fyizU+LfquXO
1DsRZcpcmx8RjrAXHr2WHWNs9bKEkvLY8CKphQPN760P5rPBo2BB7xm3pSY/D9v+
Y7WmVnH7U4SgZ2WQnJPmvpQbsdjOYvh7/DLw75MLQfTOrjNSYo+jHw3XyJIgnUey
vfmfLx0Pb8c6b/+bWWrxDnk9iaq0+GWjJHeWq/BJrFsDVGojX8AeE6e+DW6qyYRV
tWZXBaNzihoijhwmLV49pPRq0NiO0PR1gDT8CNqoNWSgn1xWpC5OBr8YwT7mwokW
vcvBRkRuVfT7hK0T16ViulM9VIchETWwO8ja/0bQfOwCYTUwMWpCQ3iHY9YNOppQ
xcV+G4ssKSRwb62ixTO4jvq3TkBb6F6QDbw0JRpx6kk+/VlpTurCtONA67q+BFx5
fIBiSgsQUJHb+WoBKOsgErD9ELyQGxWCcWJNy+X02FMK/64oibGN/6kadCtpNavv
oZGng1sIl+Z3UpUd+bMpbSgkn3oBX7claklYcK0chbDDphb/hwA1fa0yDEW5QV6f
gqv1ef+//zRBciWL27uOHGEH/cXf2e2LEOThjQbMaHeQ0IiqS2vYfJtkSqEXs5rG
Ru/VK+LCWE4Bzq0oGFOF6+cx9x6kjCBjkaPE5K1J5P9dT0HzMCFeTMVT1AoNAKgq
OYbtVC63pcTqVsn3J6YOTH1yZ2x52xmNGHhmMjksKxT3tFDZ4SijaOPUG+nQYjFo
/nVfypxgjsfIOVAPs5/DVTYts3l7AiaJdeK4+sM8UEXP7G4jf6wxJYBoeEFkk6yv
9NEWFREnEXD6UOVSc6q61sJfTK8n4FxHIFI6hJtCx1oV/4cUredmrzKBtfaUv1d/
zcRiQP1lzgS8Z3UA2QPhkf+4k7G9o4XBpwUbP3RDpKnS+1VQ4oPK3dAMIR7J5al/
hFQNzquZQRe1chGqdRTcpMp+BxcTzFiUpBL+tIV5DlBFwbaBCEB4d5wnm+m0TnWM
f7zBF8Fu5HGCuLlfoq/tyZRrgzGMC+S/91rhP89D/A3+sscBpgOgmfL3Cgn35qSe
PnXA/244g/NSG6P5DwinkCleEraknT9986XjwmvcNXO0grthdYcu+mHjDU4lBgkt
HwNLKj9VPd4JyrJUsUj+AaRMnYQw61EHVr0q09KU7m1JEN4Mm4Lo9jKvXwcwBLeP
HU1sOVNTzXh/azt/eW/J01hr+9Goxltf2SO/douYH9U/cL+tkq3L2JRiv4kzDQV4
uZIJXnBqCp7zT37PD8O4BN21t2DBiGdNUNNzKpM7s0lScEv0RUUzsk39KAET3wvs
lJxQgM2NFWcPBxWG3WPChYUGaKpwqv3kpUqs08xpY3XTC4SVwUp/qkcB7IOvXZX0
nyOF9nzGCWJREQYDgd3Tia4ru9eDZUo5RR9O7oM0YWHDI2h4AL9g5pKmAm5Yz9Ni
OsQ9/zcSznhNhSnBvAeNrPXCHVuAW1zDYIVAzWq2X38osbCTghut73tG5ltJcvPl
bOqdvsgZcrEseM+q1+LTCQ6fgXEiL47fRM8ccQGe/6r/8eCE9VxulLCMawYVZD5I
YABfXt5hJrMvJMWpLbyvrnky0auwpEAhrh/ji+/TUTzKj9IGPjaMoNRMrJQ9XQQz
N4SHoaQUe6rAHBSQaC91tE+sBtuDHbhtRPmj22Eth++wjzQSTMYpCvTEUFWodpgx
JLo3ZBwBve4E0LXrGTdmTo3lB0kQ2YM54Vc+TFjeQkrcyzgt/GCpCPzMzPALAF6D
r/Ok4/ool7X/ZCkkzlNNoNeDNGBpJGaWYY3bvtlo7t3GGdFhQ0mNtHK6oBktputx
bpmbUnEEHq9p7rvQdgO6hjHOw+HiEoZLLK7XFb2cZ3eMvzF6m29QZzdDmfODoeD6
TzVseYk6tpQ9/8ftN2QTruFE+a6F4g2Uo3g4px3nVabqQ6B0Rd6G3ZWiCKDxbQRF
wbyx89o+gzs95DWzE1EOfp1Y8dMMK/dX1bLy2fOUsQeIXtxj1zZ1tqQhA4QMYBu7
ysq0CAbZesHSteQ89xLEKGKNaPrOoWG5S55HVAIDJ98JVPeXL43x+pkyUEUS1bEe
v5M/wCQok9xBrG1n0B4BcqNh5zpoAk1fltMsrHz0cg5oky1IbKvsrquZhinzDwm5
W+fULnn5pfs/6NZe9Y1uF29A0TNqeI28FFhYJuSWRELGtp8qbjI9v9antJA3a5iX
E6bgp3WxoJqu1dQHYacjzMnC6EtyTQn7WxS/ENV0WiqTF3m6+IU5b9vTyUg6SbM8
zhPBOhIRMZYZM1t95xuwibMD0/Nz1DC8p8hAzV8PbXoyZ/3K/EX/Tugb6rdQw13P
GhbVNiloEUugs5re1J4/EHEitcQz39hjdhzLSDdUVVAKmyL3N33Pl9dawtmTivWS
r2kjugXzPbrV4TFa+0lTM2WMRv7eyr1hAZ89UEb+2mW45XUQa5cxT3Ea3iFJ0ydl
/MjH+95CYqrUaS6wHlxkWk4cT2i5wbiWgCdx6CdrNLzTFG4epSsE5GLOYTSDg1AL
JdfhuMVu8PDyTtTVvj9GI1O0sEhbsnV6q6zA+iaUOWGAw3cNNkrGnoj0cvZr67Ju
VQtJlisIpI2gdGfGGjdz4rUEdcmNIPJooQ2wmCgHV2V+rROw9DTwVbsEL09JqcnN
XQ0rLL33KC3iac7BFtkdgv7jSoFVL64EfHEGrwaxRLHnFSkV8CtYNXhqOJq9iwhy
NIyqEmOUIBlgR9yg4ytRNwA3IKLjKGn5uv/zjN9Qo60a/R/pW8ozEX6esPiRxwxv
Vv9pj/OfS2fHaKsFNaKnm5Bpu+X4vAsQUDsaZ4yfYBXLkGO6NeWkIK9fTc/t/F6F
sfC3Xkt7Nly2e07jaZoN4UMRtICMvXQn3YgicJPWZRIAAS1Mf71JHreyAG6kRT01
TkIWUKyTaKh2FgGNKEYrtp7drE1RFIDWdrUt6R77PZ5xCAhvgX2skE2tlQK6BxoR
x963G8rNR/UkUPSKcYf9J4THQvX7eXaGtjRVVbOACWXPrQp7xCSnf98yV1lDHYuq
gINu71rKzwLcU8Z2xja9R5EugWhE1M6n0fqw2ROYJRLYnLtV5zcPFURVtsbY+3x3
ZUX9aUuDXIg7rFU4sSBHJpRzyvlY+KfplLtY9zlV2Nx4uPG0fs0R3UpjaZ6xAf0m
cptQ+WX4yqnV+pLEMEqwXTQVkE//5UGAoIOEx1opIDrcFrKpoFcYhsyu7ydMIgaw
iOaAacG6PGsG4XzTXkcJH0vEnJaS+eYO4tBHmcCQsP/7+dcexj6XqCufh04ETZQ2
IyUWVRFITfJ/pyszvLPStM/BJDKjqkLhxteUvO8024Hm8m2lNxOgSow2W234F8Ql
6dtrqrriNJSHU+5792cuX9Y1kcG3E9GQNfdJ/vYuhv5HhckDtBl6VfUM+Y6wwDQU
WnPke9xB4zwGnIIF/6mlqmxif8XRZoku7qNL2zVZ1uTwuxZPAeM6GPGA0DDDykY8
OBJHVVM6qnnSHKCvdI6fgbemPXcZ3GVcEJmfvZSAosKk0Cji8sd8qUnWfx16tIjZ
LE71CB71PaxA6PADegh1AiZG2ci6aaS3yfku1oXBL+1nPMZkCOA6dyRzEkBDG21Y
ULVU5u7fHgCghS2f0KsN7btdfGTBZlEMNO7BIWJlNQ8OJItA+sge8+RSvqJzafbr
i8Mab0uunYJEMLVLn0Vrh2q02xnqQRCe8RlDAXCRlyCbe4/lsdfnRbNbaZN1zk0w
NZ0b0hlz3bMRBrRZWM0Fs2lsEri/kCS6DAhhlitaR+/rChgekXwcZ/mOFz9CJVTv
GvWOk+Fug8hTCwocILrvR6zG294uMZ1GG8RcfkqF7JLZ7XyokBmNP3HypzXR3OKS
upCi3ztTD9agbv4ryZ6SIupAyU5ETj7E4fGs62wn8kxSz0vebyWfRvXBfagZP+vN
JTJm85re1rfm0RgtG0mhg6wIUe2eDbFuqORSO1qqADwEnsVJHM51jy1nDkAyo/vI
iQlwUL3nb0IVlmbcmP6c8CHLJHPmhJtVy8HzFMZe8ttauFekxJPASNWrhfnEnMtY
xT05lt7GYJ4SJaguXuU8l+Cx9ovl+WfLwBSGdGSHFvPhQLHl7UQh6hjruM+2BqlH
GfDSGGwLA8O1CaeZsuK0faDbcLqgVN7WYO0Kk6cBf9BLgYJXYAThxgHHk2ElgKeg
ec1DxLeTGQHMDvfSml8B0PflLd/CD6i000FSMFRQukhWXRT00meRHbJHuPNk/u7g
V90CNqc/Krliu0PdatmapbaCXx1sWz5QOMG/kwaI/pESzUDUw6rhZDwJWUpmy/+x
4CRVc+yLvLe38f6Gk6KuUr6oXYnxoZhpFWQ2cXm15QjpI7DHz59WRJrp6MKXDitb
CDTYIcFODksbqqUTKh1d2PU/Fo74NTHO9By9y8H1VMlKyEy3B5HqLB7a3MY4iCom
0JVW0q8qZseqmujka287YIoYz/3IojtIwGPyxMR+9vRzosvvEppKTm5HnRObFMie
jZQF6uG/Zrc2816IpeAla0CwrKUP0Wm/oxLCeOhcSCPkeAt7O7w08Qlw5M5rxVFj
fsm3S3hKNzyXfXUIL3TqFhNRL/IjfIMwhtErXjjZcdw0tPRa3y+WlI6MrbTh+uEA
QsEdh9Tor+AddZMw2Wq0hhTtolC68Rs3eAdHhtGQ0U5YNY98LZeYYVtPpctVWGU6
46uvQiUR1Ir4eMGpAsXMOcBxQuHDSVZbvl329LITXnXKYKByWHDIn/BHdydW0ASD
O5wZd+bH6TE6ixAtJU2gVr7HKlwmjeJQZdwBjDkDIpww15s+feZck21Gh2m+KMRE
NdNQVmG59uWk6EHYdYIi4H8eIJGtIAKcEkTb827mziu5PuwSxWyfpSIGZY2xu/YL
/mfx6u0u470v5o+PfFL4TrOSw/VjEKf+/X3HBdDsfH0vSCVcc6YitJW7lA2NJuWU
ys68FPkpkJc5yUzSUn8IexwfxwzVdd4xNkEXulLkWhRkuKUUXX3LMeR/vsd7Efpq
a2WywRJhbeWvPVwmcjBc1OzlhD3jmRgF9T01EDRQys61QDGeZLlNF12qFFDBypSX
3qKq1Bqx2fzL79IE932pijSQaOR4pStqoUiI2I8skqlmYKJ7fN2Rn4swzRzucWyP
ZSARLYSjAvt/+aV8IkgehmJp1a2xej0kHzxpkugYob0XxRiYelNyJTK+lj56ncUd
NlSaS6oDbGM/FsvmwXIF+EvbsmYUmKsRauA5Wv1MnQAqeV+apvyq3ZxX19meV/+w
HMrxt+tZ4WGJg/MtQJpZD4xQERFtmsZhJl/C3B5U/j45zkkrlFaGg14l7qW26fh7
0eOaVddmx1GjNTwMRwRBv43iklDiYgEbnbP8TSC6GLwT6qKBRg2xLNLSVOhUzGnO
u0mroBS0LOwoW9X1NuxihnVBDLg1DVUMBBPdspcZnWzdYMK44BBgtQt2XuAI8Yw3
P039Tgxkboq1oUHZvJXsiF36hp+XiwP0lErdeyjaSuCFMLqFRbp5s8k0ueIunu5M
mTH9Es3X0xucpU1zD1vWDPpWHbPsvuqpH7uhoO0i2nTN7b0saGsWLyKBO/U+TXKa
GtXmAV97oex1Wew1gQqwaBpZi7nQYWWiXM5cMDGbtXDVTcyI1kONPOpPji88IgWU
G5HjprJ/h31Zpfb7ECHh6j9GFOooAuYzRgu1hkSvphM8S+hgK8HIu5RsSTd0HKYG
/t5Qwyoac7azvIXzUpCw5uHOnW/ak8pjjnh/WuJZxDfSv8tVZJRihcNOGvbY0phc
mlfsHUod0O4A8cE491j3d1ztdWb58TLrUB4n8tBycKbxBXOW6/zMTCFAwOM0J5lX
V8P5jFPQBHURoKOTosz1d5lRZcluTkbfh3XsbOyGHJ3tx23eKYXpRFFXYJLMkWFi
KEDiKeIh/OvSB63aCqLXWytunmx79Z5NXDXf4GRCsw+l1Vzr364h4VuUqcmBffUt
HuaFZQ4QspGfiV1VjbCLw7OisxAd+WtDeGemSuOl2qQvT+G/kioifkFpVkT/1bMo
c9g1gw1uWNL+dOdbjezPGvBtA/Au3XX4EM+Os4ergUj1Ui82Oj8j3TAnwqTITXMF
ROIyW8sHeijEMNiM/rbgfG7FUTQZc7gv7mlF7TmvPdys1J2eTsdVAna76y7rFMZF
3H4Iq/6nVKG3U5XisisA3QHYxyqMa9t0cch7MDXrLu5SbgJ58KfGN80A0ZIEpKpc
ez0n5+Jr31l9fnb//k+syRKOg7hLAfkjQVxBtgoDR17up6mTJjphqiU/PejgIjmV
V8/ICmikhBuBqgh+Z5GSAZJgrj+GEWvSIriAslJ7T4Y3fpm3LisN20v6wbnTP4oN
U5MEXl2iOjjjVuJvn2R/nzTNIsJAhe+v8KMde32r0NxP1yhFJw5iL2BWKMebQ6jm
g6wOHIdDhncoBJoZItkTPUcQMtIiKk7ciIxYIL+BcNKHBjUU/vZtOnZVFgjpTuL2
jL/OQaAw4Stg/LKb/pcAsGwi6feAlMUq8DfZ8TxRxpopnZdZdXXZ1+0ODxv7aW7h
4iv69VqYjtBbFSj/vDhn0bZfpNYrM+ffQSxdm3MxK5wxDLW8mSlIxjChzZ8sV1Oo
6+ZIt+oATOwSTe9Vq9xTCd831wa0ZzSFljFMY9TAnyv4M4dSWcewmjagZ/BmYoKR
IJzktOXaJfNkmzzLmXE3XJUruy3oxViq3trOCGpsUhgjO75xCB0yLLc+dyhcja3Q
j/haqY/7ZhpHlW3+iAXqHRBxcOoBCEoRaiiFBJuRWgF+s2FQeuyUBPQI9FkXsheU
FeSkA06qD8B8bbQ1aJa/mplGmdpgSyEJZcE/5Sx4RRWPm/aHRK5vXPncrNoUxZ8u
L7RCQBuCCjyemLzIcjj5ugIdD2aJj2VSCJ6vTV0MafQrgiKX0J4zNpQH1L3PZn7h
8a8s+jNicOnU2QbiZlTK0R4frP/9rvpPphCgzxYEoQEeIuuHLSZzlID89Mq+6cbc
CWxp5nyDuMVIU2/prfwGd1p256kwc9FIvFQ7C36zjJyM13S74N2wt/BmFF3B76VY
6v5o82sYfveScGCSwjQ1lGwUJcdgaiaO3dbQwTF860ha5OQ/o1PTZ4Lh1KNzduMu
vocS9P2bbyU84BcIW/ZmM3Opc1Abmv6kyD1PZ+wV+82HQcy7EpI0XXlaTvpHaUiq
v+9H2UYLUAEmxPf7FS/wcQy52ChMkJLq6JgRkWm2xRBjLBgJNZaLkgUVpzovb04/
UR4F4Ra1TQFr+w44X08i/cS9KhDMXjAwKLy2XqVPNZ7E367ktpb+zUhz0cExeMGz
Pn+YGmPWs+ptx+SX0aIymxDK8lguq6nPkQy131i4zzVDgykL5n3zw4ORRVxp0CB1
VneWxna615tpCCxPPaDQNUvVv71+RC9ATRudgG6iCYqfcI1nBlIRDWq+D4Eq7WWv
hSlyzQKeyNid6YXH2SDkGiXwOSGVNqqyoz8Qcdq/4Qj1M9U7Fa1uFs7Cz33OmGnr
JPuRZUPZq1p64hCMccRqZI5qg8WShLCYo+Cm/5WAzPM0IPp+6/Qow7qoLjvKWvSS
qozteVRmOS/YTrp/ApcHm3d48DbeHrPOqMSdi+0/bw3C0zSPghWNMlI74u17glbl
ZawSRPxwo/JF7QGNuckk8tXq6O39EyKzS80M8HSjFPhsJFudH23kPoz24aV2bt9c
Ajy1JVMiLCH90CcNVKfj3erdLUIxLfEcb7Jl0sH2SzXrGE9Lz3SXqX21a69l0SDB
t9CiDuWDz+Am4+O4ht9k2Bmp6ZQD2rBFjl9w/VHPdJCJ0frS8R5a1OiACRxbTsFz
Ntl0Ui/VnIBAs2+kN5iF1IIy5RKj3etf1IxPsFN3uPTHPfwE/aoagqCHdLeEVqol
7eoCto3lGb4T6xadV9ImWE5BVQMRlr3pHw+qqjC2yRc/FFE3i8rG5s+2e/iPAlj4
LL693xTC0Mi7rp1L7K0L4Z3PmjDJiN6Py5+T5x88o/UrKCeA23Y6exgXMlXyqRke
Y3A0KVQXrqr98MGscjMG4b6h9JheAX4NdEVBuflUC7tfnzQ7HIFvdjzp8w3BdiAZ
Spt/ATdOzMQjzPdTEXCXai92nIGUBOoe/KS0rd2v56zFJaVU3RwL5YHIS0Tj8guC
E0raL2YLzeUkz+zKZLb6pv2xWFJ3aoyjHGsDOnJF6wnFO4k8K3iKx9TgnJYgyukY
NtaFRt2bowhKFrPoPdQWOsN7Ks0wCJCtbDSgdi6UDZc7X6foiyWrumEKeNFt8N2h
B+KccBe15asDEaubB9zl3KiCBNBdG8nnxPOqnEsVzJSkkJ7+0eXz6NV3n/k04efK
ZyAkGZkMRAyYjADQL0vS1x3dxyexO48yVS5o4/bFjYttRO8RzzpYy3pVXKLiA0OU
zdsK7n9lVvzFPDzi8QWwaPGitdY4mvXC+7yOpZihtc7EnmYMUxWDv5P7HtAiBT7Y
0sHJNqyw2XsYW8+QfKa95jYsEbPESf037xLRkNLElC7wY8q4cQdyFRD+7wZk0w+x
uUVRy7g4g0Lrc8+JVgglvdgzT5PuQ4Ngqewx5bZYykYekyBUp4fJA5kFj/d1NN25
VZqgvb+HmBTCNmX9UIxn/9bDJpF2ONyoVXGVkq3b+3IflvtSLvuG4iPoXGJuXinj
9/JhLBH7+EIm5/pCkORq50MxUgi4q6iigoMsn9aIDBoJDvCaQ9WWTvJf8Twzd+Fw
es1RjCf7XZSx5Xq1JlcSAjaVzNi3BR54nOW9dIB1OV2ILCjykqIy0AUWi5wGs2yX
rSdD3ER2GMEyNHhpkinp3HWX6b2AkaDm4WUvVBaBctnuwxmumrcvu8C25BtxmUrS
Mhbz6IUB9yJRsjCH5Cbfa/1Hz34J/LZlrojqsu+3l8yZXcgKjX65DfzlBaHyY4eK
n/wsN/PxLhAz6Kvhoh6Ckjufk8KCOyUmpsZNhjdKs+topc0viPqsNpB08MT4fbl6
7kYFLA9J9giM102glxJaDBTA1rNqJpY82PTsdZCUOV/tAfoh3Bkh9G47G66eF+vC
YJBPPYnVtRJvEZHwFpqVTOMwa8fnB2Frgqq0xk7U+yXruyhRAhu8ciQ/UWtEBSap
8LAPBih1qKxwu3CpM/CScpuvFl/4YavtNila+LXUcEe8BC7TZKi5EoM/hMk/Mpy4
LqeZVYAeDEAqQ8IUqiuju/peEKUbAKKJFur6AGA+93wBFoYSVDdBbjSP5rQzhMjF
G+SMCn2DAhXcH9PAeqa6MEBrzTNQ20Wkex5yyv/UY+LMBUFKbjp3mA1FQZdfxM3m
hb9kHItqeFxEj6rbeKyspoOZSNce3djATTWmPEr31mIulTVGO3WLawwDKPiRBwIm
J+v4iTbz79T9IyGdyhbxTBkiAsw2ww7/WY4W5oAiHun6j0uBndA98+7DAihOxxIf
rv1RT0T/HXRCEh5ih8qpJ6/xV6xui8i+KLO7cfG/zuhOZhNo9Iy+gk+9cr8F6qzc
zjf6ITZcmEwH2UEnivyXLWiCs7Tdp/OCc5iJIO5LfQxhe4q7cACQohCqZnvA891R
+I5T+vZvJmuDTWIBoPNsTYO++D18zZqCAjD/vJkdisyAqJkNFakeNGKc43K51zGd
OqncgwsN0qZgQZGl0u9+CzCfLVzsgktqv1wJn0oFIR/PkODP+kwfGoJHUdHUSKr+
7DvQ2IlSQINa15/+TzzhhB6TTtegrbSCKv4wAbbZRpWu8usIz1rkWq1MUhJvpTmh
oIaaWUtesJSQ26X2bsp0ilAPUGz1R9R6BPchEqnddfU/5Z8ELa1Zmv1fKr6PXOPJ
6lNyuv/2kzf7vZ2GYEkdu1IWiiHy1zecv2c1mfZgssRF++yLw20U2z4x3OYr8zQP
QZ5fsu1JONg+PA5GCngymLJEfPzKQjXow6kX34vPVLQHt4LwOMoToWPIb2JGj1RU
gpTQ8A4mZVW6tx3MLPxyL9V8eh8p9OdYSkEcLfIbN/+CQyfziXxoiSE0ILtKE6HQ
pRuPoLrbb6uFfEYPv+/QeH9ho60V8+3rn9rVUc4RIKlUqk6bjeaAL/PWcCmLItlp
/9FwsCvoN26j9h8Eh0yRCBKLNpou/Z7JE+tQY9BesUuSV2ayaw1+27n/MFYFV1Rs
M4jgdPLoue4EztNKxpeA35aGha17gSUiBCw/jmLLHwZIjt+ipnk2bdseGetRs+QU
y4HxXEFeiKERqwg0LG0VMvnHGngAtdnIci9EkHRayqNe8h+fIpvUwDqcfphSHwZn
JXk3YekmkY/nnjvn3v8BHfTWw4qdvBbc24mRtUputUbbwW7+ZrMU3YjCBT0dfg6F
yjrgIga5AVAiYfZayJaS+t+cTj7ftwnl+rRiqetdyMq18jgCqyZroRjYTbRwQ+Pn
q9LUPH9JaC7y1N/GPda7wgCNhjcX2N9Rpna37JH+2I+CrdDXjhBjVIfcrscY4ze/
GE3aYBhGUKuCvJIPnopDrzrjZvakhoHVLzsI/ygCwwgQA65o0yK9Vczq8p5949AE
Pk9OPn2ie7ccb1u0ghO8u2Ln+lGjoPjmcaiAMUk5CAja1h/LyOxRPtl7ev+Ud+QX
W6gPjycTxm/Dp/Lf5prO9AQv6jDwajrFu7YZytfur42JZ9jUBULVAELemOA67BQX
cZv5uVOpV4epKSPY7n8s/1Fj8dCmoRkIuwlBxbuJfIt/FdWJwtYBxGXcn9o2ZuZl
6V3YExtUDY3cikS75iagVvWFLLIOsNApEn2tCqeXHC6CXwPFQQPnoR/8EvLdj3jB
bZbG/lFgTkSPEWQohdE1k6KZWsv009wXqlCt1pe6KO0Cvc/pIn2mNEMbahudJQqy
IAra2JYfkkpUhkX4UUhFJLHCYPQSBrKKa4u/ZypLBTVOMLNRGep4aHPJAeZ8KYtO
5yOvePwfalGdoN5qWQx8Knv51J2Ejgi9CW3ms0M9lZ7ysjBMXPm2LD4OtC6U+YQg
Z1mgTYbz0v0iQBPhD/ZYLllxdIDXbVr1f3vpukSjs22IUsuV9SZwaskNCyhPKwlO
rECAJRjKKJ3q6eJKAN+cSo4cJM44gt8X/1oMm/K/XmgF++F1LKC8z+tXGYAx4shh
EWQgla6PYaRWd+CyhDl+uplROzJsa78Rg/z+DrJ4QcYSWpKInUwh9kLBayfKvom/
aZPQVHXKQLvH0BJR3tSAlA6BZWI3UOOvI3ISI9Eo3wsDh0veTK1pQZSTFkoxfWq9
b/Xt9R2jQas/M7w7JILExBczxR/jctZklEkckbuSD52yvdJ7BnxUKSprGABnjziW
Ynin+55HvsNnVPIqGLbmYdFIiNcVe+2tBH0zB3LAN+ybikqIObAfjpH8k9Z91fvJ
dQuqHV1yPh5r8q+TEWYbvUYdgWKI12uWRCASXiA8O16OWJhS7W1j9V1mFRf7iIjL
n2Y6PiuwaExq6AS/nmOPyBSSLP4MChNxhkWPppEbiY9KNw3y5fXrheBNSeO5SPnA
T5FaOs94HDt9kqa4UR7mlbrCko7adqpGMdaKWV+i6NhM/X4kroxIg82pVHqxUxKM
2lBt8c0D2CgrrB/azGyWmjjl6AzJ5Xl0fvVtLbw5RgoL0ElLADI+MogOOT99UxFX
RW0ItKduVId+O5C4KWHg5gWbqZ6O7p3NKyxtir4CNzHoWHnpG0MB8MxUp/vUMmXA
NPNL5lnjhxRwUUXZ95zrt/iHIsxkfLT4MyVyvIHGZ0eSfwR8CadKCXlwJuGQBE2W
rcmLY7MjcJ4NEgClUaUX1xsCy7j8AD9nryRZAkPpfcc5fe9awFTECc1Z0nbBPbKa
y/w4lPiJNjHDO0Yqr6gYlB6qjpOtwZM6FZQyTClZT1FndyrwZyZjSKF89rd/5UuY
DkqGZJ6KSAVPOGUABZXoh8TPdrKkzzmZwUiEhCMV/STvhMqy8cxfxYN0tqeTEFto
WKnclF3a9Og5pVih2Q7MWfVlqFgxXYf18JhT7eqw70+Jm+Uoiz3LyKTpTpHc/uz4
1K71C/FPfS/7g17YLZ2RV5jqZTe1TiNqW9VqMV2in0L0gl43ED6Yidj5TUTorh6z
6bE149CoFw7EFXD2ePQTbSzCsawyWjmos1bC5kUSiKe7jVoatI3P9L7dLC9TCGTk
iwx5DV5lbBbX9skcTKskCEV1kDBPMbfZ1Qk6JUr+6JWnXHNcx8aXe6EYGkkidT80
NOM6/B6y350xRyu3fraEIWgzwfqoMuBnPySZewLu3kHZc3jTjfH6GYYgE6upHUfY
jw+rHCg2L1sDhKNyKKhtmVYcVBw3GCYItSCSanhuKrGY2jEYyF8jEOg37nLPhXOs
e5fwqIMsoT4mGoiXsyLNXvfV+VGhPIb4lD4lHg72kHfy2w7Eft6p+oR5HZzJnc70
YuFAoVoaHVL6YtEYzo8inGOLCr4zWrPkNKDH5Hm+jehrrK+eNDu5t0GnDWeTEGQB
w77aA5u2S2Miicmc7kJ5Klxm4Wcn+pu0msgE8v9c/uokTmmiVF72GzYTD+hv8Owu
81eQyfEV2XMPfl6fH0abOG33lRetIS7rwL6UC/OE6jqTYWObnXALASRYRJLOco0r
mjI8fPVl84KyXvzmGCoVa18H5kJ7PMcjAurAfuu2nRUkFfOGEfxdSa0+YhbvP+n+
bczQLIyrk32kQeDl6ZkokNn35whqdkXZ0u54o2+rO0NA80xUXhNM7iLFCj7YtuoO
JTKH7h4Q7DbiHzM0ITdTDf7xQK1JnYne8tQ4+QSh112/9+cOtX9sEbtGEFbvbOAt
SVgF26XJ2QCVw06cbTi1SHFdBfXMK9mkGtrWmANLJequHRWECFelp3SKDSDceHJf
10RV87cjWvkm0tfowxIW8pkT4ekBVzlAQ2jI7r0W7b9MnB20RUQUhOi0E/YNcry2
8//Vw9fXv7BGF65N7+vrfDKnn6P5J7TBG3NviMkSJnPRi97huC0O5EwuM5om4w6O
pInyiNf7F1B3Twsv07z5ZDyLmll5H0Bc8i/fUOCpBocMZs4Jys/vEPNe4MTIZx3c
jAlSJz1B8PUq6oFLUWM3AchDsoOqn08Y4jPM4PNROYBEK+F9hLAJzbpb1pcuESJE
1K8zvy9LO6hL2xtx4imn6c/q2TB9o9PerHG+b09vWHG9vo/6c5yk/9gvOjRKkmgZ
GfG4FMjXJlKSa68DFXn6GQq6TaH4m2niy6KRyes5Yp+tVFN+pH0w03E/TsMlF+TH
W9sEYvmuAsZk8wWln7hUEL63ZvAXec9f9yS3UYSsG183ONb9jOLju0lynascDIzx
K3t9DZe2GHxPYq/hVOxQ83KffM9G+97o3TW3y9DQ5iGVWZMCj8zet/yfazKD62eg
nI58IBpMytOw4xxTJeXSKtVaiXwOn4Y9GxL77NmK4KjHI8bp4PR5bOtfUc5uxSQ+
x3UyOIr1YiZ0PIWF7YeFlF2wZtBWcrbNpkH9S44MwWwiAOiQEQbzPjQx9f+lav5n
cnpmCWmMAJ3lT6n4wqaEyVx1nEvce+kyxmkkdpL6bCh1/3NrbN4Pu7D2SYkkTPSR
SP8CacxnP3D7Xllisp1tfYPzdBg1y9px95qjMaFyNEiqgjPUb9+KtjfT+qbf8Eav
QVthM1AtruptpubGhIUMevW6KNUbxE4MjVxhHZI6CQrFZZ5MLOgUVnjGZfvEQmhN
Mq3DXyoW5Osqf0IkzkJxskc4pmNUGDh8qurioL5Cwhi/8/cwvuc3WNFOqWj1263o
UwTHRUyED83rfUxWsXh1ivB6SacktWK4nfsH0TA4mUrV2FF9C7V/SxftLSCMqH2N
neNB/SmuTUGCBZxSs8CeA+txcQDdd1P7CqmhRyEAN9FwuOz/Rmow7Dzi/HByTKnT
IIMvJ3ISrBLm9VmwxSvq0FIrdmkOvOM8myN13qV9n2LG1dUkCqB4VdAf7O959xWS
IuIpiUST9/BnFQpxtCuEb6+bVdHUwe7F+OoU11H/nyFo9WpgJPq7i1BqH95sIXFf
j7YTiOzsn0EE7Thl77ceqhBs0jSnxlnj25kVRolKCa3LVYNMUhFoESfdK6xpMuVR
2BKeD9HDE8DEVV0jEffrEO4IRvEW3O4Rf4xamlnReCUSOdnJZ7qfi4bKhNo4WZ1f
GwP4XI6gCAXCEdJEeLLMCbLswP8X5kzS4j9ractLNy33cnc6QXaA3aank8brkP4/
a1moIdTLDIiXb7/nDiZ1xA900rBr59XIGQfXSHo3WrF+/ulsx8DCmS/BGZtx9Wup
TINi5Tft48105gh59JzlG87RQUndqmJoSLTPwaNKUkgQ1jpyjOq+EiVhDQWCLgWx
7YllT+8cL+YWdD+NpYYK62e504FpeAXdACJ1qB96GkEzeATwaHSo2/oEN7BEbEI/
OCT+Gh0g3iVYpmDN970qqZJbo/X50/a0GrDpJKkiiBrkrRTYyhR7uP+XIQ/ozjQT
Ip9p1el6N9AR9qYQ4FZiRF+emQXk9H5uOp8WHa7NjI1T0xLAvwce+/djewa4if3v
yESgi1GuHUO3Pj5rlg1AL+84reeruJ7g1VSV38m42eNjcXZPdgdikoefD90rXelD
xJrtXT9WzTwPPBVDU2fHj+9ZzMmjXOk9bVKl5fQkZ7MtcgVRsnSv8YR/UBxMvCuc
iWypnzeVwFuRnCbDqMQCHzeMSCupLg6skS9r0jZAO5Y+jAyQOk5MPlf4ajR7LO90
VOjv70ndN38z77h4jAxeJMlSctKjmfhV7Jom44ifuJmy1SuALYlzDfjjHnGBr72i
gy0XA6GgHRWsBg5jNPgOAqMpoYxqd7b1/Z/ek5yI2iwpdchUlYUgyRt/TfSSnVh5
h2wE/SZ2v2u7vgoBBt7aQEOUbECxgOG0H96OlmEplsVXfEoEELjF/w6IXZbvHCaE
/JRtg7ztjznj3lUz0wJxkPLnBbU8EEVqbduFWGjO0bMLJ2i4O1P+8GRERUYaQkPJ
jKJQP925NbT0DbSivFd/QpfktITd3dN47tKdlR/92MC2p8uF2DbjYc8bGr4r4Wdd
NvgQsKfH9Ff+T0YnZuhgfuy4FQIYhKe2m4UzD5bZUIFXJ9/HK/hRYuQx1kuTztM4
i9iXytfX3fxtgWmwtfc5kfvWcAfcARjQ0BYlQFzLspMRqGWw9sy9wLyzOBqqSN59
k+t0N1zLr24tN5n19+tsESSwVZSPrrbNVsMLG95tLhWFBEplK+VWKS7ItGd3+EWB
D0ifRHsq3jABRfJxzWQHnSmD2nwutdoVEjMV/TzE5x0pDxzMpt5xWghwhCPuLsU6
NMlsvR8Bu365BWg8AJ98vq6NOv0w/pKXpZvsz5XQ+L8O5bL1YSUdPxQhrONSW86j
Z3lsCFB5zYZiBVeWt68yKWZnLnH4YBT69D0+OsPbcw+8Ld/1aZhHS8jzPLd9S4IU
f/rhQX0mghEASmyHcBgrei9xqYWiElxgeBYVU+J3lWefnaeiZwzPdbjPF1xqzH0M
x+md0e8O7lBEQX37vg1a7y1wJJvsOPCX0naVqF9Pu370A62UzUCF8bu/rSfStqR1
sWat69VUV/H5D+gj8W2sNmn7vwZisjxibNEHyH+G3jysjyeAseOib+XHU9kw94Vz
FmgMSF3K9VRs2QJhIpLuql91/SY7qHNTQvfQJIT7wt79QmQJk3VeropBkNaVWa8R
UOu1mjebmiybZxKTIFjWQVg5OLZW5oCZY12UnUVqHiMRd4x4fvL+Hp8x0zOL56kC
lSBQUSfiXobgorjFopcd+Y7yTRvaRY7U76DyF8lU0IlvgZD83gleyBNjpMo5h2kd
lchUkhMcENPPaBWiSwMgGyrGF7heJk3pOX5p2lY6IXvS835/gg0MLAUHIk1Koh1b
esPHslBWdl2zn7r6HXk0fRuTsioa6fJdfjp5aoxkAi+Mw2LA0Tc/kuOxnRnkCcjU
4gQDkm9k0I6zcFxPoqgmNEtQAX/VSdNriShBA39mBh9H8yTP/sF8u/EdbVH9vovd
XvyU0cpumbWmIEtDU33fX3WppqLYjHVZiWa2zitAEV14bV/bXRU4kPHqUwgLpmXZ
TpJwngTIMJTW79z1gnHj+TDXriP5sqgweoCHqWRzFAl8flwkUYQT11MqJgAZ+ag1
W8ynjNoWuWUGLMYuknt5ytAPmIztaTQhzWaEpa4U25PwySG0TCjIeLG+vIzSy918
UO7CA2YqHp2963jkwL7Em3vFILUOZ6Snqd1bH666HC4xy+P6y0BTysU1hLQZNpWL
oj2HkL331T5X+4newAxyS0P/ITDYlJhUPRjFDJ8MRgw1Vj65GofVMfqanRfKYmWp
xkKwuBoLnPD3NQPT7/20LYSHTyzFoTHHV4KV7qTiExCPvLOsVJIjKcrofQRiTlOf
QWuS2antFflOGeExZOvUN6oP5hK+4nhbsS/DOkVRrntUrzSUM86AlKW1MF4nzvCh
4RPZJ49ESCg/srNjzpKnPlx3v68DJXlvsNGP+AhlMvpsaPK1ZdXGxh4buXLjWSaG
dyKC3eX4ZvUpWmu/5hMMYD/sN0rmky9uQRqOfsQGIBZp0kvnkPa25a+BtZag0AR4
x5XRpCPKSZF2uDU+jRmQnM1OhJ9qF637XwtGLU/JiW0aDbVH8iaiDsRMSjvT2Ggb
whaS9/UbrA6YMGN2GqtUmGbl7GUbnLCiNs6b+8U+dxXImHFVa5nrqPAw3qnHi06b
0N5AuqLX40kCDHZvQ6iKi6e0GybYNg1vEUMg7HvqU3lQiF0DOhjoctVOyRDuBhbF
JvdrzNrcqa0xyWCbc0Ku/YyQkiks6wbbygsExEvr5jWxfXgI2JFgn53YON+cXyjv
8c2L/AHqbtlw1l9U0d7He3WUxgUeEPcsOxGETveB3JrjfxWEfxjW10Mr5GKbvmvO
7E6PjBWn34ImgFU2orT7tH7ZbPb/vK1E2cBAMNwnVfFFjHGskX+kQX5nanF9UDzt
9SazqDyJgT9TKuvv+JvNWi7Rus/YPZaNp7XEtTUTMY+ZMYV0MtYe04eYz3YKvPcG
b/S9hbVq5befxpUMfifIfgEa3C5doIWbYJTOesu0YH5U2JugSdOLWtp2rlsX4Alc
ZioCrwAs1aGwEasJu/oXGk1DdN9Y/vwZn4IwjSB5J+AJeADrjadLV/VPz8lW/gIW
SPJ2nkRT+3o99cgZUR52dRRTu1yKag2Ux4X19F2rQV93j6AVap2OzqPsjdBIPzds
AqFLiBY+bhQRnclOI4K/zbt7/0ruWzH7dud8xSjqRS6xnpX6uj3Acr/rxgGE+MG8
AD1aCesSRBaY3rfALT/hjzYY1A2tdEM3k6cHAYjdpzYInU7u3AbUOhmA4eDr8LC2
lTdRTsPMvm9DzRh+97mf+jlDm3iaVE4HNqtKn7gZySYgcHJxNRUtdUQr8EhwZkZ6
7sDWA2ZH/Tw95C/34Qup6JfRVqIgY7ThXLNdosykG8anA0QuLtIcyEcY2UyMasuX
BIFORDe2p86HWn3T/7M8Kz+Uqe9Hu2AT3RvN2KK0/8VPALJb/Oa9m4dIylwYqxSh
9vw6JLlALEItPinOCh67+e0HJ05HFfilpx8HLOlq4dDpyBjU1QbT28pV0nIDxdpk
FH69EgaNjuJd3zU5NP+Ka+oex467gJuFoa9XNiCYLRKnJy2enZvH6JvCnzrvXlTH
IrCPDsdBSyB5eYM1GumBafpITJeGACMsNOxcy6xymSPb5Qt+IaApap1zgMzWchmP
68DS/gtWfPlazpl5tHTzLVnU4y68YkzQznPc5J/ZL8HBxHuGCRYm2pLoasRiYU8Q
pENQgNUdXfPXGsqFCVXhFz8gd37159DZiCJVJ+vFasvSb1cJITUJEb4dKHu/SSyo
3g6SC7lcP4ny3LtQRFFWKhXBtXxqAw0VI9dGcHgEFt/oA2m3uUQE6S/d2rEgU0SR
PGyJujVpP5N53gHgrKR77HY+jHYYpfHafBNKugq2l6qc8DgaBoX5eI1R0Svb9PdY
rzMUDpbWa/rEpJNUvc2i3QwdFRZNGQCbz5YIvgrtm+AMPV2G6uVt1u5Jpl53D7qD
AFPvKKDnarvEdcSVSE8ox6EX96EHT+bB0Wpgqe9+PyXdWcvIQs++p/sBztImZrWp
wedRVJD/pwTA1zealyp6dFk3iRGt1R1/IbNHMjOtm3tmfr4QAqnuqnZL62iVyDLA
qJCoYtDzVyl4ep7hIU1/7Czy+2lxvNx+decmf0Szk6tzxhaeGf23iRK/dUpEqJwZ
kR0tBqpEV3cIHUhpl8B4qQ55xg/FeV+NfWUoyTDlqFH8AuXnrlApDi/6OKV/A7rY
QRLuvABl68CQGdTU3j8JX8nX0SwbvYBZEEJHsOIonIcqS0jTjIntPqX3BK8uNAhj
jgx0lU0CrNP6JV6B5l1tZyb/L4APIJhnIFjDH16HaHWyst+Q4itVhHI5UBKZfTlg
sqHjWMAAZZOQsmocZhJU30Nts8RP6UnN7mw1TbKPowNtf+DlP0UFas2jVtuSLiM3
tu1ndTMy/NEDcGkx6Zth4nWX5cDYA9yUEQ/6hszUaeR/Gz5WRI/MUY+EuUIto/+M
ddAllZWFCDkjvCP+0o0zCv1wa1Y/vk61pJJTLiVbodroKmulTQr1b2bSxzeyY1M1
JOu0rYqEuJTFBBdm3yixIfzASHMSy5pYpIrgqZGb8x9Z94kFUf93l8JOVg1CQn9B
f06wJX1dI88uze8BcM76++eKZdiB71TVwqdPBsjvx4Jw9Mz3vKYLkaSpLjU0WQ6v
zx+N+WoLI4mUkuc/JJY/XecenApVGb7h5r97hH91pPkUDGa9ik3biuY5gmV+uB3m
3Dgw3JEVVTYFp7GcR2ZWQB4cUI1AZWGoSQjB4PuUF+6vod4DnLmHdyjj3BVwgFPm
FT7FV8ZhdDWEB6FU+INuwvDTsb7HHQ8vexk45iFajX74Y9MRmr7qEJ8/KR99C81M
PJ+bzmR9RHXHkOoBvVJg/UOWvwnSQu5wGBst52jouGBuhpXyJnDuftxDC0DNf1hX
udR7QcWnL2WX4F0Gfu7Dsi+8GFOS4jnmcQpu0YfUWgz9064SCw11w2evM0jr3vvS
6gBQYWg0xUqwWhxK3134Tk1GFm/xISet7fj/lXxuQICkabnfGLy7u7HR5FO5ox34
8aevD9Hl1g0UFEDHzg+cNl3AT9nIiY53upGiphSGEMP0giAa8dr58yfbLkzVXem9
LJtt8q3Ig8ymuQ1lftAFu+OAZzaqPVnRqJd3xW4fWimEWD9sBkoPgcczu1b4W5hQ
v4T9HT+NHc3TaGXblzTeBFzUZr9udZq5B3uQuyLpwvDh3A5ey2gdB5ANSM3cWeJX
VU8uza3VILxVGEk5PjxXy0v3f3khaKrvry72LqrxnxhM06P3lLS1ZzlQx06OK4V/
RcPVwb2Vtz3QnfoQQ7rhIAWVrVEQmLv+6aejLbThYkgbSYscwupY2Td58ymD3UG7
Vchu9nWzVMmTMx7LSExaeRP3X/TaOGodHzejpLTtd80LO0oQRonghTNngd12JVDT
t5EN/DEJ79KOvOE+Cp2XzEXc2mGIs63hZzQZXNJ/DGz+nvosjtwooS4HuRZJjnuf
pGnaTCCOA6PUaKwP5Fjsw7eo1FxoU6y4qVo6RC+NxGEDE0KKMDWneDL+3/G1Q/2j
qw4Yu8DOXaSfvxvlUldJYQsAYt7CcEO3RjvR2IMniayS0YJTonHE3M3slrSklfQy
43vzomFeaM/8RzW1pW2dHlgtD2LWYruRHdxGlFwpyns1Umy+SDtsmBseGI23WY2I
fIcvG00pQb2+fh3qOaOlazufZQBGhyl8fNfpSS0z1bnZKmgK0Nrqq68mBNrT3I4I
0T6uNMjMvuS1c6vqitKGxma0vr+Q70KlbYHmS8MarY4Yz7OSJ03ggGgX9rs2GtBp
jE/MXQKMHGnZFS5GkHh1cofKv/iC/9MXA2werkJBZUiHtlKK8WzKnyT/4uKLkCNk
+uwboa0EcV58pPlKnePlJYd6NFE6GpbY0q9e3WZeCfGgylqXQ7z9L5241Ww5yd+s
wQAAbJV2KzuqImnlx1M0Z9oNHQoRxrzyphUAK5VJPAY10TxH3uAgLFOUn2iELjvA
Tk2rfjBJWqXlGbW/m6Z+1uH0QJM7XqLqCpb9540BTMePVuGU1MNpLpMRHzcSOSu2
PGn6rZs1brnHcFOAfglmPjSoYTla7hIUgF/Y6FueWD2QuxZQBdoS6t108sesbyd0
F3aD7UquDQvjju3QIV6+jM4LyimMV9Qc8Z8nikfucBGiLARdY/uriLu4k/FJ8hUY
HB6FJ9VI2cn32fV5KkERfRwjPe+nAbWUZTFp9myvxV+KHMGzenuo7EHSWInoMyqa
otGbN66+n3M9XyigTPILYeoPu9Evp2SaN1mq3W5pB7cLrF79kDHqj5I/rqBhgqZQ
CEAkdMzGzGWSwf+1xN53fmVkbX0R0istt2XAVoZWakgCrjL+zvMEeY8xjH2gQpuk
SP09+wVudsHUdQfrFLoEeqSH7rJh3yDKQUzTzVPBvXjPC1LgAcCTsoO6zDS0DsWr
Zb9ITfzZCKVEEwc74CTaus/GOo/70YuxWjI+CGH/uYTuwtpfnQuLEI4KO1jOi6zx
s9DJrQb6Oum7zBbKTO0KOzRQTVyCmJmxKLuyHbUUtWybqTESUY7mO1K7tmvpH44a
005GzG2uBr2cB1iaX4/wAMz/SIexOcfte6z4JkQiJgG51arcvmEP3Gd3I69kY7B2
89SRx7rMYS7g3NdJq4lZhWFzXn2i74ZX37zLNua/Nrw/wa9mYjdpt4Y7U+wK3jB/
Qsc7lUl2Wm0/J0IgcXqRxMh2KECmpTUjZj6QlA1/g/EMRD3mFEH8RUFldhpntABW
78GhbmrXZw9Yx9mdLFUZG+dD8QRl1NLNB3iIZ56RWJo7ghDwlh8PVIbNVSU11VEo
OBmSYmJC4P8QQ5foHeHCCZrf3XzC3eD2cShFDKlrtWazoFQCocVqzbNBEBNjNzHE
CszzS7Wkaed1ooD3eerV5zWajNB5Jt47WrpJu2TGqYXKhZ72SB38WDzOWwiPs5i+
6/MkgLn6QsFOvRjUjmeFEa+OqpFoBXM5ci6j57IsQkae1y11qyqfjvsQSQBidzV0
Qgx8AnbG2TeuHA10qEHxyl5ulBF547ug5q7tuuqgfGmFBdpnyNpAU/7+iyVAQWLh
iOQs10iHW87qmk5p1tHETgftxJb3qpaNJlXBc/VHkwkaZbIEXXmBcdeg3FYXdYwE
qRSJXbcCQAcKvMJd7L5hPC7XtR2ikzJCKefEanGDnG00QsjMuEl3dSiaqmfw+wTE
CJqd/umjeggOC+XWt13QneVfVjQKCAHbyNEde6ZU9edtLj+iG4UUlVoBOcTeqw3e
36oTt+X33Ky3d2KnZpzLrM4oplcrJhnUkTyNCTTLrQ5JE23IOFzqdhPR5lUO+KcA
F/NKBqbamn4t/ITRX0DQfJveIpM+KRhxHqr+l4oV5Nvx8jabcVApqBME7HPvTLYk
AszcioaPt6yiIViSDN0L18s0yIp3eX9YV55ovU7jB1Au0v0+zaAKeS6viE6/bWmp
TDAjgsNHY5aPzR6+KV0uZFMuhxHfb9ySvkQHHVZxTHQtBWJdk7NxzihEwGadoLXe
tHIxJweA+iqKZSOlGjwm3JTjBUE4blyHBeOMq4sYf044joc9jwRZP1haKYUEUNii
ZYC4kM3bY/+l6UjmEi1+GFmncEt27B5kiDX6/bzJuHZs22TRNLpQbnCjWPUJ0xY6
suFOkIQM/beLS026LN3gx9T/dCw8cyeb5K2xMyaSil6Oky/tz4h1J3lOZgsJ8FB1
UoWbkId+Q3C3eMLey09BrtmgxeW/Db75RbjHdoCDJRW9hqaKPR65YVfUjhsxfjM8
CqJqRsJMifucUUeRBXsosTu2h8gdwi6hy5r9n9SPmdGSO7NVzmI23JAtN9VBUAJP
CxJ3jJmi81BJt1WK5xytoicxLSvyGGIDaZetRHBGhEf3YPkIWNAcmHh53AocF/mv
kC4EbCCbqSp44eg6nF/kUIprN/JRB3iGsI0FZc96jmr6wQ5G56AugQQuW3cN9fIe
mYACNUUcrGFxUb2t3lH5OcBz4HigCubKGQfKKZM+ntBWeZRXDYcTthlW+T5QcoKf
jWm3SPkSYfA7NgzbUTTDy8XHNmPHjH3Z6hegS8SjmfHBCiHURJ0LJWk+D0QphtPy
tv6XG6vekRlKQ8o59YBxvbrhKj1wqTLaO1ghtHQEJPbjfZKIuep9ThuD5L8jNtdK
T8ncZsAxq1/AW57UbKmJdJ5o1cNZXNHbIgraC1kxF9SX63negliU0STwt9A+sCi+
BVR6luG+pw+1r/ETmkS4x11VbkD8z9ox1cgfYBhtej2NbPSxBv7MipKo7fd0Hued
F4kxwMFP2pUV8cDd/gvlXxD2qiw/Rpmsb3HC+mvVU3FJl+f0NWhtr9rtMeCjZE2W
MCRk6gyNkqZP/Eq9IfhoThJ6mcfATFADUSJD1bwEWf0tzSz0y9n/p3W2Q2YKvisv
lTcHo+/p3Jo19MEmcx+/Cwg+YgLUZGQ7KSFJANolYpiT2jjR7RkznAVT00QtW1II
U2qSfELrzkFiANew3speGVBrfHnehIbmWJz5YbxKAj1B0RQbzc5dzL0B+tNC0YCY
F5RCFO/jdL82+OmyRDZvRktmW7q/0HMNXEsAQxNhoEs9pSoZm9Ula2F+TrHCdjyj
UvkY+ODfZeISbPqUnD7QOg90pr99+f/okL3h1DlLut8VhrjGvaXgvvnflwfx1nGd
Y6WPEbPsLC6xtB4QndX7/tHaWQmIWt0/DwAqNmTCNKv8pSimxd5yMSjaGnW4ptZ0
JSNjm+qVo7SBXwfBgAU4KXEJOtiPavg6Wwp+PlxexM7SBXRyyhl8qjGEa8Qh/KUJ
0H+dE0v65bdc1NeA1sjyza9pQPsxiVHbN5cI680b5aSnsFujlkQseGqCm+D4Q2p7
9jrd06YGTVRA8xSa4UsN9PtkCZxsO1eQ95K8oc3DhfW1SawImZAKqv01HOfiJDe8
xM+5rvAipFXkzocidWJj1sOCPH+4wsGdfwF0HmlRSdkqoCdl/ii0tU55vxrbivYT
C6sF7yGWx198vY4CrJOqugqcJDRBOKt4DMizlPo2FLmtXz/7zg1Ecm7ZAQEgiIw2
FX75Zse62f4aogAYclzt9F6TtItxN1NHPlQgeziWgpX5ng8NJqSNBulrk97P2Q0b
LYF2BM/AvgtvxqdyXjmZFdWSiuUVcwzFmnpBvimNv/Rpr6Og0bQ+lHAs0OiyiSIB
dQaY9yZprkd7H1L41V/bg0IqdvVJxrHCaEt5BDBLEY5w5i+gccAgxWzH5avLCROT
TUgn6xCzPWd4D807dSJcv3iFTA99bwJakNxPBI/cmoiQXAR7CmSZE3bLycX2KXFN
nUhUui+L2he1blkEXY5449GdBJPHJjiSzPl7Ig8NHMLHqGeUhdolmdZqCGv1m8Kq
M4371tkSh82pN2Gon6vL5Bcq4eO4SvB+rcKMdqnpV28O6QMFgi0FNEXcgSlTYnCA
uo26AejG2IuC13Wg9RKdFSIme2EvKqq39bJaxT+RvlaR4sSYBe4Jmvt0IXEvO/Ej
+CpF+/R1MSvJ7NeJcO6QgF56h+f1v2PMUgcEzshRV6KsKajJjCDgTnsC8b0SRV9d
in1sCHO/xFWVrWjMwO0g2j4idPpLXQVPVwaXblwQuQYFb+BBziPSMEPJjFm4ND2u
7x5W7ic4BeG+E91aiVsMmvRg/8Su6NAGVtCNQSGzMOU52Xko/3PUsMZuDgkKVutG
aU6f1exAyeYruAvqmirO8a3CKjVgTbCZJkCDE6DkPyit3i44acVpZYA/s5DYBDPF
wlK86pCPzbMj/iuMu4B2scr/WWBVDavbyT+remUL7nOoymxi9xq2gkyrrKgV0wy7
4k/8u8qogRZLksXIvnie0HGZtLrxz0R6bWfookpnd1Dbmt5daQcwX+EPHzcDAOPO
Q2V0eh9+dtwO9ebJcEdhdgIN4mzmXOEeIPt5U3xCdBMxivy828ng4KiIPaAD6wh4
N6/Lpw/WjzFDQLz0Jp85gXlb8cDbE60eQRCSK89qMm0oDJ1kIwyu6BKeiVlZQEQX
dEk6eun3YfbMdlDZZ4eJGMEozWTQkGDfg92yl0m2M2SxK/odmDDSNjvKOHjPHCw+
RxJumjIWpHM8AiFDxbhgmIcN2F/oFlRTNWs5qSRQrpsxDgO5HJ/2zSHBOVR/2FIP
dVAVD4x4DrMf60RaiCW9jE5BTpFH5YAjKSmzrGF1SJOz3A0Vmzc6l/+4uaEZL3xH
/KRGJe43IGgkP8BQE7HTTvZCdKc4bbQQYgSExgYRlUFnkVdyBrA96BX2kJoHuWyI
PQY2APdjpCtSm3Woo27p/VnBKnR6LhqPHtCyxFm1tOUsYIk4/Zib1qVErDBLR1C3
Xlpl1hfnkevsG8EqLy/N+FCx2LBPB9tx394gPNir8fHz5jPD+z7eSbNAyGJTUQ2J
uVSyb8jJczidcWCg8QSEGheb/0n026OJg+0TzYaNZFsqo7+0xc9dynmvdXXv90lv
O/XYIyGKZPkWyJjcUn1R9ru2HG+qJ7gw03SKk7ZydXMDN6nKFtOxNdfO9fg6w3pb
XjEAJmIkBHcM5LLraTceTVohdPNIySBgT3/uT2AMobe9JvnybOV4koXbXIHTiYOf
cXVuOfVem8KXzfGZW1COafCRKw2k7gQc8Cy9KNa9H53fg6u/z67lsOv6i/UhFbp0
pgibgUZaatPUq1TWpCYI9Z0pOIEDRpn58GGGtRP9rnuD+0rYAj/i3R+pR3s9WgWE
/35jpcIYjAEGkwRQm608qGP4062E7cnu4cO1+TwtvgbdIGgG8AMHO7Tx+lLdzCkT
sdCHSoBndgn3wxVlx46+7mkMQH6TJhwS11sFltkGnCMBcVhtjDaDBKJXKouUHOg6
geHksoybYNFNK6IsKloBJi1gbc3e2aZilwRj5DdHCVOVXZoKIswZm0pz2VGHAeQI
nDSPNIpj7SNXA8Wzjapi7Os0plc+lbsEKfDBAujlL9RFBNoIOLjsMUzwDcYZYTUk
Bex62xrLyjVIsa58ySDwXLcDkruziyE2RswYOtdPgMkVBHsKyS99U4H5yVfIUdPT
MDZT8UR+fGsZyTwhVWkeS8h4FbY0xE34fRdWUBzzETGLtlUUC+bX5BJegjYhovY1
YmwQNVRrcSU+yUCrPN+4U13d3fLSTtqYKtUCnO/zLTzosl66Ra2VBfCyXVv0nB95
NFo8te/z2iZroPHo4MO6RfwP0tcm2weL+bMtvmOKV4LN89mDDwpnu6efffU2EHqQ
wjFGE7Td82ZFOrk9X14zr4uSSgeX0KmSiOcakcwwKXXame8i1iQiQQyu0Av/4Id3
tr438e6FSfo4SYkY0wqcwC6WCKEwiye6HDZElUXw+B77HfEzwT3WETQcecqvuh+r
QqQZrLZQA/rHtiwBqC8nI7AKI90hezxhTHuXcttl3TW4tZ/B5TFpILsMgTAuTkGp
quVKeEd30fEcqmHRlMg2ag5EP21dTh69rabwRF9OlKSHmycGJfBPzxTQQP/u3OJE
LA8Rb2FZ7F2e4AwmCoQ5/qsWDlb/VqqcKSjiAMiNcM7sbBu03AnadHWK3bRBw+L5
bP4NLMMKx5TVGTZ8pCqwI7aFAX+uP0tbGIYaGLIX1/WixHDFuRe8KcmSQldBMpmC
pgac9G5xvhOU+Up+mSIBQC8rzlH2aQxVue1dGHiSzP7+yFEtWRFvKnl2oJxmKq9d
lPg2w6FnUl2LZClwBCguafu5zscg04+9xE3HracNkOjH6Jm6IZYJaPoBB1NQhJl9
bgU0zs4Q/uVJrcykxwnxrRkPHYxMyiVRuCe0cTb6FZE3TosyfO8cErywmoean8YU
RYJZ/mayZm9xag1rRnzW2q1+j8QWlXE2S/pUZpr+O0euVv1VBopfB3wB3PPtW3H/
Qy7fhD0+26X51I44zoDA9xGlAEq6kDSVacEs+70X+pvTLfKMTLE/E3KKEZF/Ygao
jqgZ+0kTq1FtSKCI1cAWx5BHq/S3kxg84ZlB+X45o9PyVwI4sHPHRWFdXHUbg9iL
Uq/Y/aOWITby1QO0makkkh3KT8MYCc0yV+4+UP3HRZhh1otahuJbEC05X0o4lweb
S9HcOdJoh1o9i5UPCND2TMRrSEI/Qrh6TyGCNDxk7KCQnAFl/y+Olu0xpQl8LfQh
5TBNnFLTzz7suZyBPDR16Jgdzk2VL0GMkHcwdnDMVnjIyvG/ez2pkXYZyTuXD3io
uLLN83Di9cfRiIqihGuedVFe6/Ub/xc0F59794Y1r01vN0cCh9kawZGCj6j/7fri
OyVsR1dje+NoN/Fxrx+HUb6EIu7wMOiN8uOfSwyKW8g4RtbRGGcLdi5F3MEXTOsC
ofv8LJURIORvYGqxiJ+87HFhG38opShynijxT6GMh8WyUIfMoKFtzogI/JIcNkLq
UWr2HDpQ9pI2IoldsUVFN/laCVTNDWLcUcnh9jmruK4a5mBeaqIHET15ceZ6ZNDL
+Lnm9X70ubxbDaC1uuDOEaBCZDUMwCzBHm5K4976mE+gHOJqVv/o3izi3YPdwPRa
IRjDPIKg/9NLgCkYr+j774uDz95fXZ8+Y/Dzg52tMqLN7jbbf7YgbAR0K77FeJUz
6C7TlfHBtAg+2Hh25++JfGEcUGzIS6XUfkD+fFtkw/6H3wNgXU/DwQf3QQ8fxbQw
qMoVrd5yQU8rRvxYrMaE0TOiqtjJpHKiqaLN3mMxhnYRJihn6t1XK9qEb7YZ/DMb
rjGRV9pJb7WZRotds1GOCEEi36IhN7/oxtSqpKgcNpItyACl0koATPFpAxugYnGm
BUBE0E9O92pTnFmXQZN3pCtG0OBDLkk8KAhiPjT/o98T5MqQ4Bw2ACeBd7Sw1n/A
fGUQrWTII3J+SgQ83qerSp4hhou6C4vKWVyhj5/ugf3o+D2q5W23YpT9uY288OJl
HcnmFoj2XfO+yeVLVT+yYF1Ieuo8T4s41D/AttzeUD3s/y6y0RUGcpt65PXACmuY
xS8MqDrgtU2VwaSmVtsL2HDuSEQL1vW5PYmxw/1YnTek/bT0gfjW7L7XuCXT8e71
guOA2jFFYH5jN9sCF0HbhrYckBlKXVNRCX6c/SX1cX/Py98HLbZnjnXUPbyg/3sm
r2y4C4EY+UL2TX5VTOj9nBwhS8X7l884VXEkhsktjRatwSDdW1YOIbZ+iG1R7Dlu
NZU0obmzz365bY2mmRoSZXwG3O+a2Ce1D2YKOZkSywZ/wFi/OTMnFCqmh/+8JKN9
yHRG4Mx33EwbCMBJ+9Qjf9qBGYm8NFHyJm53x1PwCEDEjgo/1h0m2tlSnKO4W7AK
t77kak1GRfyqTEBeeVUAihpQKddhfeFA2WQp613ULIRbYttSLTIQA1AHuwC/ogGR
y3aBBmarVjDkynzmQVEaCJQW8HLKaMp21KUcpo5qo4gJATVq1busjG+Y8Kld92Ga
E+aJtKLN5tTeEI5w2X7C2nyUsX0YUJ8bBx+Qji0fb6hT9g47Pi0v6xNlBc7UpZOy
oS5FXX0exU/EN2aFohEmbV9lqA3FaEZQfZ3jyRsPgOBYZ1hvUHdXZuhVV2mi3JyJ
l7gope9lwrhI2EkQu5q1iVvCBJxdxrGusYehCEwJNJlyr67gUiQAlMjs85mBKWAv
ezFTpjRt2S1njK0iaHNVPG1XtJUHaT8a6ZP84LHn6YipBDPipe0Pr4DZvOOw94xo
XD0gRr5jWUfauFYw6K3Q8d5h7P1EaMaICQCScWfexnwo93JY7JcNz/Ek4O1dE619
7MyWDPbu7q4HqusghhF0twOTVJSDp+eL5cHmXBy4xepEnlsP4+w97aQArj3IMvSe
p9UM0fh4IO3Q+3iGTpH+cl+PF7os1lGvgeQptv4Mc3iULvjolVfe8Xu+kliUNMvi
Xc4NnC04Cntv6kNH7PczBKbSQa8buHkpBX0zZtfta/p5N1BLIbYyu/7Lcnsf9dAb
2j6tWkqUirU2qmT5sFtMVNAu1fw+gCQ/TxETTNF/FAnjLjpvn34a1mxVnbNIKX+4
shzQwVq/ASYDbApcQCWly/Ga9qauDh1o1rgk/b2+HpGbDW7GZWTi0l5xtCdhdvK5
dx3CwcFWeLZydnJSACerxowZ8I//vIjab0g43BAuH86WnznpcCRbkmvJx/AGPGW/
9PORZV1SlyTJBrRy6juuLscCh51mCWFfaT1LwTmFc5mANJfSDSCQ6OX1ST2/lbmI
SkbBZI8wuKgfINwPwMAqbyxYHg0weea4kt9iYIko6x0J/uQOdrNeFbBjs4pAxhp0
pU8KvNvWtsErnocWTdU4RSMOzxjg3mWU0n+xm5ItnMJy8x1lS2T4GGL6bGSGzzu1
3F2qbbRbaT6UPKIkFwiDDY4dfw/tQQ6wzAE+LrWtoS9QDERkrA0m5AIP3CKcJEE4
rcHs6+UI1uNupKTFo39M4aBG6OV6alUIRFWgispDIufy7YOnpTiBHpzqG3lR3N1Z
Uej3AyMSChIozREDKVvHMUMebzkdPBewe8m5SmHwVxBQ7ZNj2oMtvmC+fj1NYEjn
O+JsbTzds9LqUwFEL6lahiTotoWuII6lQ2KmcGf+ysFG3LIL5rz3KLg7qd7SAa7H
WjZjAqN+EqeZ4kyBH0CPsQv7Hx+/SH4oSwTaW9vMjdfeiyttcOAYdSWimpfIHVK7
CcW4uJS//f7llR7JMOmSFPl5L9WD+cf16Lv4xwLpWNyjDTkvRnbwPKQBmQM/6iHF
eMe67Shoz8VSqD++55hDkXF+dF8fbe13zGhvC2VqABrof3Lkmmv17HtXuCd4QS1I
xnQ+A+TsJYPGxY5g1oAQI7Zh4SL8NVCsaRTQji97Up/0fVLvS0uZzwDIBQgbHzfk
jF2ENw4f4AhVsc7dxDD+On9XWRc8nI3di3Aips4r6vlQ49RFBp+fC7j9V2u76icK
osjY8JdJR1BniV2pDJwjjJ8pCHlRa5JCJcG6ZYq958kLUAU/dXGM+JA7/0nonw0Q
ZD/scMGON8lIKnvsfnf+dB6RFPAYxirOdrqaR/ieuhzhtaRXYHXQwmL/rcf+xcv2
tgtC3U1Xe50PAvlQHeJ7bmRp0jY54P2a4j2sbqmaYrj3gFstFmPLE22EKVJYx7cR
kS+IZ+OKJ9EoWMNohlEepm6xSC9U9EDtk6klHdRS1xH9RyQ21URSls6TMYEmgUvK
gaHXAmrnnoVKncrBeY9T4O9Fo/gGBc7bO113pziNsuVxB5LGhPGCezQKb7khtRNG
l6t8d5JxRGGfHkX4XVNijtJLqY3QG7QTBSUCsaGP6unBBNx81PFVYl6jBVO1Ge4s
528xYwU9Wul0MWHDcb14RDheaofbKODSFnDrf8/Jczqj7qghXyDnuAxVi+2cwAh4
5KBEECMRCcllmCj9QlDrYyfpUhoD7cPFPDdAASbyW6xjCADVSp03JDyTrx7DZTZj
XcWgfPVEgRguAvVlgImq7OXv52wfrNJWuUFi9NNZMPWaNwSnHIthASB6kGqb5IOy
Z3Gsq4jafC99UY8jPKEodXKNMkYl8k26tw2Tiijrc/44fwLAjotRyHbAwQibbqls
Opcs7L9llqe93qtyQoEbX6dtB4Y3+eC5+VpPCnrTihB8bYWM8KNJj8fewIZipzOM
n1fhOUVQAAaJ8rlvm8Sw4JN8gGLiMzbxzLvb/e7R1QWjlyySTvhHXAwySQJnxHla
ehbj+zWk192zi5rIgmQ1U63NUNRFe7m8/X2qAeC9IjBP4ZAw3smCsLO6SuHQ/vSO
anslkIdqX34QnvnHG+2oNNl/VrBcYM7WTn2IdiH3+j/SyvIvVvTMgAIWyw+3Ii0A
tjfTN++1zH9GTz59wD6q0Vek1RMBEWJrNTRrW9slFwfOyhYvIN+kcdfkPwIwAlE3
3PBFUXxT9B1bTnlepzXhQb4enIgFTHWMgrPq0zAl48LMWMho1RL/k0YIho5vRjvv
kydvR6tf/+n8BgOXm4rrHo2VaMxuN3tsfNqgy76Ki0heCymVqziRDjLtVJadtp8A
bii+UGg/jrMOn+eeq/X2m6rIUDNCLErdD/YtzQs07DCRXin/smXQjzcTxC13JnkS
BvkmPWYiW/0g1V5o2ciD8immWrK9/q3U4adJzbU9A18vEfSFiqxPRW7t98X3f3lW
7AnJa4qkWmON2Gudsm2i8OrgWdjpmdTWyef/ysFlFlEXIJsviX48JW8p7X31+WAs
PN1oAr6+aXxKzAdC/903p32S+TpIe8QTbtZ+4UC1T1zEvhgbvPoJIvNUGWfmghmB
jrxPu+CCf93RprNyaPh6iP/D2HgtEAEKDwFMSVXyozEaEiQfMAQXzDbsiJ+FHn7f
EgYZQlFBiWs0GYzuocKYx9UamU7IeCqoaD2zwu7QUbdBXZ+0eQ7KLn0g4Qg5sPBm
dtE/ES7K5g/2zSW4ovCPZUzisr9Pp7wV9qermNkXuIzJIDWGpqhPELpSrQ071nXg
He45bgU+UXcscI/yFDxCJr9nmD41J4qE/P8GSljjA0lL8SZ4KqVBRsg+oANtWc5w
IpV9UfmN7Eng1XLsr/+1xySxMwULDA9w38biiYYHLRwTkEx28PFuKhBmF+Lkc0vW
xhmnVdb+MUvXfLgFj+K+PC+PT5ffDojJPzI1VXnyCnUPNKboZMDe8JrLEXudDLD3
kU72nmxFBJgXhZV77OsnUBfGzkGK/yxds4uPZ8KYczUagVLOyQOjy0xYnFsCZAM0
nDngQJgNlsXxdjWXI/7ysiGhLGwGmEu8mkSTtQgWT6F38b9mdDwYS3BuTBxH79rn
uwmm4WjjkiQD4tfuOd/yTV3MzrSHhDejQKLG6YOac2TBNgQRQhnkOPoZkCAteZt2
9d53OjHzkZuavA1DDLs4FmO5VY6uPDPoxf+xY4BDRDQh2fAfHmHgbSjoHlIYIYqQ
DPfxJbwvdWXj8Uoz5aj3/DyOG8BuadjOc+Frh69ny5brWkHkhN8cUi48K01ecL5O
HNnfKHKgV27iJnixgq1JB2hYMpBPzARmuTUrQMgEvswMVSm/iblMnXxlGgDtN8Ln
E30EOXOjyUN4+kboxBqUlxjdhtZ5jLonw4UEcuYPDxac5Aj1p6UK/ZaRbZeuisnn
3zmOCOHzU3oN4M1YhNA9CEkRgMJ2lIda47pzxgsw42W7NbQrwnkZ7S17ycGtC8tc
a8/iXkyS4LrTEassDmzeCd/LqwkUPofUYqwqCBcckgVFQX1VuzGsWTDgBwpbe4/6
s7nGrLRSh1MCE1P3MBVqiyM2ATeT0UhkeDtsFgLGK5E8ishPu/Q+kWXVwXkTRb0I
i9dEUuc7RXppyMiS+t/XTCggy2XMjZIcmk5YeYWeKNn63hWRh320CMuF4nRjkWwc
Fn4TwIFvpMsBo/n4hV2riamGU7oUi5SG2z1dRFOK9qaUhCL6XqmmwxywMay2dybQ
M3hXqJZucfaPyRsxseGugZRITLG/aX553Y4YnKo0TjgwWyaZibDc1GS8JkoiRuYh
0Mr0bQfkZ9kv+l0zK2d8dx+LEeltH9a/ID/yrIM61o2cKs1g6LCI4+FurHgQi0Cs
PXbF9mpmZcbIj+2mB1t4hVnRmfHJhSwcav8VDiIyw1PKMkrJpgCz9/VGR+Lw4EPh
/doaKvrStxLJpORbyZhzOJb5GjFl6Toz5A/EnbZTgdRRAxtSIRfXkO8FuavRa89M
NHj3K9rgak5iPSTQwPtJ4Nbuib5CO1dWhadeNHLy/eqXvg6nvKpRXhA9nx++L5R8
w0ggdnmlWYIFYhPiHh/0Afhcm9aIWPY/uEoqUFL1M2FwOX7Xy1rMS4i8ugVX7qbb
V/Pb7o07DRh4kkgXkCMgEon//a4bMm818obfQ+RaU7R3fPN6s+K8KcpILXqoqQRc
VAP1jQSIBQPRenNI7xBaB4x42lu8sqZcnE5qnPqOJdgGWlDHdbuhvItKf8aLrukS
bRfigjUL0eWaLOWrYL/3RGNVMHZFIKh+LRhXViD3p8EnyuLx9gBqgCSyxD2iisD3
aqeHBNVh/ERiuc+A1m1MylsBq59I1wae8ctznncyK6LFvZiDUHd88fFfmusZz4Da
ZDs/If758xvJonpv6YtNnxBQi3unF8kC1jcwEnMQYR1u8Ti7AlYGV6F9A44MdBZy
apa6HxXtLmgX1YH4GMVkeKJoe0qnbF/fhSVzTjWvwT4AF+1IWFfEkdWTnwJRI3zC
gJM5AdCIwlT15EO67woguWacC/9a82TVNfRPWt9sdgZlncPoN+cJc2h+pSrnj7T8
xnkgNmwchFCAtNTV/UHnHFoDINk1hUvwulnnnFr0rTcONm/P2+UVnJ60eO43UhDK
rUE7f67Q2lYRy+RQWkJNBwDtnqUoDLzswXHqsccusMZCiuNuOydFaudFW2OzCMXt
v4ni3AkXKKdZxr4TjTzufeFMyarGjt0GC7Wo671vy5dknf1tvmt++lBMZVH4YA0m
GIy9F/+AMmbrA5jbiTYcjUOyAeBTuY8h8TU+tUUXDlS/6mcg9Vdx0FKuiQrjFNul
g1ODS34K3itthTcNgRZpRfzS56ZlyE++aznOYrstwg7KS9axIWfaZPq289pcSRNy
EBl5oG7KuQWuAKc1wboqKnsHBcWMu4iiivGNfHwu22+Iko1zHjzdrfya926WwUOi
CaM6ECnOHb+gtNmulQFRLsg8PRnLnxQSP7xfjOvpg4JVlSSfyWR7KNycxs6PAyeq
xsoYWSelW2SOsGvXg0Zjz/HOmwVIjBXKmHakXS6EWEPXdOZ7Va/WF8F/g8ADATVq
COKF+FxW4Npm7w+7bORVdDOq3095MvQsg6hhd2TFjZGQBrvprLAb/e0mS/LApg0Q
cjzIxAZ+C2Ue9EZ5W2CZgFC7WM8Kiq0gR5QJVx+lkGP3sywJVQO24CQe5Dzi8hcd
PESjdbyQGBOPD4OwNYATx9CsmJW0Q9+Vg0uKMORN4IrOSZJIr7fRZb6EW8DoRlrj
ZOtUy58xooYXCZEonJ9qxL+LrJT2jjxFyGk3FYq0Z6JavzluIJAJM3w4k2wCapvg
5PcGimLGKVO+mAKqQaFRc0vOJjJK2SZq15QLS1PLRpuZ2N/8J3OIzjC2ZqJHefvJ
TPaynVuNKOmlzQ+0mDcnVP3GQ8lDfNBL2CQM6yQC0CpaGiNNiLQqv5P/wfwhepHe
BhP+EHGGa2+dhYe6SKw2cDjynPPLNZDff2a1c6F5e6nyNF5gfHykp7ERZ04n1H4C
xMWO0HC/FO+iMoBfRaYW+sOgUfZfR+HzF/DnQlTISiwWKxcHfPZazUivw9nK2p3K
m5WEmijyyzn5IJHb92Bv363xhhQuAmck1LrHt9VDoumg/W3mZcv+/IiZER8iJ1z6
7O/QqZ3aBqGSMqd51nHb38VhjHQF0n9R6j0BEvf3gP5bQh3qkSUyB4BsgGTLshDj
YZoQermPCVGqyPOakHS3foknwe8dfXdTCOms1WEy0xn0hNVug4d4Wa+FPk65t/IS
BPGvVOTIWo3gxpTG16YbrR4weh+NjWXH91iNFIK++aT9aaHHRE+98DUBp7SZnvhz
9AkWuszSR2X8XS4X9kcgspSPbjX8mfz8q4hRH505Z/mrmjjtniEYyuxA3+533dkk
Mr68quCSVGfoAkQrrm6bjlE/h0uyxAt7DZ8QemqBPfUWpJbSPlIUhnmS03/9vzcZ
SkdEQTNRkbxa9x9AzFzdOcGKAEqw4IbQFGh5LlupLs3+rIkRJqoGW+/9C9mZLmCA
27j5S1NNp+i3mgguFdsrqqyCiB+7PWzR2MwGPld3qck4gsQdv0oDLv34smbCBXmx
sa7crTtVCTmlt7MOWCiP9XPOMVt4kuzgz5igpNFGZ3YJxDSViAXVyovzW+B7MFBv
cDmqkfWwiYoNCGXLrYDfKbJLMHy520zKb75P9Wb/EdWYmXokUbtJQwRr+nJMMu1f
S5WUvsQH0Hujszd5PD0Micy22evldYkQhAvqeA2IpOaQjrBvYzuCfBnDvyUTRFDt
Wv628gi/1KRMRDIbzu+euWMCez/P8S16R5CQXLiC/0zbEjvyM7BqYmags2TpWeUG
b1l/7roPpBjG0b1iI+Dec6u/c+rEDinaXKKWo6YpGl5Bn0v9N9xFFt2DwGHrZsKY
VhdPZVpglLQ7xVGUj//9U0T8ClsHDlIkMjN+I7LUqxdvBOl3o1ucpUXwNGXo7hTO
fyuUyDpB3qwpbRPul9F8vuujFmEfiVAFY5REK82If8IaM9mWdVUtw4X57GrieHgE
3GxXX5bkh6uM+yX29e6XzrxYNDR3SJLw2c+f5+Hj85BWNILkVt794rRz1Y3fP+hn
Xmkyd+SG/Q1HR6DbQtKZ4gOrMLNZRYrn59qjjkUIbENXUiL3SitF5ebHMXSGRrgr
m+GkDvFCuo43NTqhwvZpXFDyq6tF/W1DzuXS74OYUW+YwTgwzTvOVoNLMC9SP9Nt
SYl/Ce677g4qlM9QFqtmwGjux1LXogtNDmdvLIPWMv2ZLbU5ldcccHG00KQZdMoy
vl4OR7Wl0RmrQLZTQO6wHOmP8PRnUDhpaCUE74nAiVjSfZ5kU+cPCchBcvn5ZGWF
g1gUGnw3lSBFScNmKur8efG2YPyxzbGdnhsYtByvdYSVCScycUr1v7wchw4jYsB8
bdfHEnh3OwXRozWlAJioK/gBzWsNdCjUlV/mdo8uE1Q1Qg/hoaJLpEn6H0nKRaIn
K9WuL2Bfz1BU43CZ7xlOgW9UlHZSnOAWgRE2Z+q0pHcETf9KZ7FWswLyIIeDW0Tt
Vrk+RmJQOPZ1cOMn3tLNv/8nWS8qdgt+0TrxuVRq54UTMXTsTw+jI8f3/8GZOFz8
beNNv3PC4q8Bj0vO3zwZ4N7gN4Cyo0HT3qzwZegjIfc/ZnQHLcokMe7o4QaxT8CS
vZgKXXxcvgsv7qHMQX8J9xs27aY1wzoq6JEezo1RmH/3nD/NRcPxg3pEsDwPeGeu
1ekHKNs8//8bKmG7J2NCSI2Mehh8DtYRP8kPSm8aLlLBHTJiaNM4w3wBkeMLoBW+
MrKrrmQcxqcwbq0yART3Wu4MIqDzN+BZnjCcJi2p1FZor8Ik8OUn7wTnqTSG3Ij3
TnnTEo6QaoP/25qUKknfvLTl199yeWUD7zkBUBatd6txoS36ZZHEmLcL78cAVJUd
pu0SDWfkgWxSAZAm8cDmRLXzi8MFUkuqbFBoW6NNweSLNa4VdaWkkxLIbtZw+RE6
u/ZhkG7GKHl3KZgME2SjFF3HlC/jbUxfreSahwugCNnFtYHQd6kdcWWYmvnoKxQR
ebxR235tmwVQ/c9rSQpAtw7QWOcf+mQpJevhRhC898/HtEjVB8LDlqNfj7vJV/jt
Ykir7z4g94HRSD41cgPhN5KP11Ln3/HRN0BkYPyW4IPYcaRbMOWoRbLTubRPN9rn
AAksMRHEQgQfFreJcMBm+dk5se4/572Tf3ik1lvJw68gvkjH25B26u3L6dp3uktb
5pnF/4kpqwb4WggFuStgnUobYGbcESAgoV2a38BzsLcMoKdkLaZjLkiMqVliS6c+
uD/p0FlvUsrSJ5XIEAiBhGcPCxqWL8WWW3+O0mwlSMDNLkvIoiFeGA1Mrm2HNSI/
MmNonUu/GfekIvUHeIUM2urxdLHBqauFw5rhB01i7XfO1TMDznUNIwWRrTc33ZbS
A/NJSLPUQ0W1chHJAjQ31Q6MySE/yBEKB6BoJulaiNTPYyKV/kNndybidvkbXVHU
SdS9EkYZ6dR9OVbYcV8biDDaC/B37J+LfdmmkvrGb+y3xJFYDFXRsphVwC3PjjZc
1O1zQZd8t2x+hIiI/W6xFY3eEaI3OmFQY0KWenA1FtwmHcJDOvU3O6fIa4ovY04k
u5jhMkaLwCjsGXv6Iv6BUQgPVND2LTZ0M1E93tDh//LXKjG7Q88SP3JHczZYT7ZS
bmQlUUps/a+fZnQfSr0CWQO23jQ1tHoWaO2ivywrSXn0hLqCBo7zFbZqif0gLjgR
7twcdEUrAyj4hzHEDQNejRPm4IopK9Y5lfKYObTiYegQ0aWvGDCMWY0U8pzpFuat
5uOo9snRbsThOAHOjSFMOeGpBQYLAkblp/yjbrDM95fyoXxMQ91JlhCY1GlW/GO/
5nUPT+vmwZuk6/QMVZw0Nan8Dt6Ber8WrjkplUZuRLD1yORQ16VSg59nR4hpdnIn
MWVpzPxEmFsqYeU7yIixWu3HPsZ9OK7314OJc2+W2qK9hWhwkzSxD08IcEtlqyJE
q1oUpAdX7AckPpMpeTxOgJqFlhLoQAkIGB7mai32+XcJ2+5k3x6+t8Rq+PP6Dg4s
WHASeNcWOuwK6nZP5RJsWijk7ltS3DVJIzoAHZT6tS4sMm8+QXCoF2ks1+u0mOAx
XcYyeF2M80QIPlGVFwXt1l1n1G1slciRqwKc/nhC9TtKDP2hgXvKBsh0sCsVHqWl
Nu8B+ROQYEchR7Yapi0mwTL1RMQAhCuRjPrLDjZyT/WGpAzHfUB5+Qd6J5UC8+sp
R26A1IDK6qJsGfUYaOcp3F12f+fpPg1EH/LYJxReTpmlWRr6NcDIXkoLvsBeo9jz
bff1vQOhRaltAMxGfyC97kYk+/520uBS0lWxL2mZZ3EJisEK9+4UTLoudjVec9IP
yWjY25rwxHAMtJwd2Nu2xNGLQwhLM2dXPnzhadbndQVvx4PA1Hg+eo6wFNXjTxo1
Zt5XBx+ZZok6x5EeV3A5CX1I6WyZaGI7+MQQ7ty+F9S1MrGH1eaXgFpEifHOlHhj
WFfx2J13aZPOSbKtziY6RMLmNL4cKrQfu5maSduvVCxsaQwx1PBJ4omWaVDYHP1o
SXMBuMpzRkrZ7W/q/rsWKaCVXDi3M76yIce6v9y2nwNbumQK5qkFi3XjfeFfcX5M
JeaTwQyrYBk6x6vtdxM8iKeaw2TVZBfkXXHCLMbD4B1natb6H/NUBJHycNNN4WO9
Enz88Zm7mEKITRinoug6NSxav0bBcKZg4o3XKySIw/+Pqnx0H6PsTH48ew15E3qv
7pWxM146JuyXqeNcr3HGXeB3i0RFxd0YWo6ii3nL3lGxbrzl3X6Ot3PK93ibygCP
ppjAlXRQJX3fcEc6i3P/JPYtx5J0SJcwJOqVUfy1w/veiScNkQp+zzY0Hg0okh4j
+zFvQTigVdsi/rsGak3yb7c2GxU93M1ycC8x476vOk1WdYBV0mOBEd9pnb7kOhq1
9icmj63S/xF7kjjd5xXhY89NhEVpVyDviMvWFtqjAFP3/KNkJ2teherZN8Z1ZTtc
y2YTwqlMwy3I2R+mxUEjLtfhK5HTtrfEMEhHVCKxh/dWDj1gS38PxRCqLlUQzV9V
ZGSx4lyhJifGvfIz8We5ayJaohRFn5hT4sboBTXSJCwt8Dz4Yuq3Sqd5qTmTfkXR
TbuWImufzmgiMMIWgzIrVSEQu0kxmpxXj1bl+mgRbzzmjROpi3RGIvLgkqCEGVHD
gtIuYI1b/Cb7oZxTILyhmToSdNWcDdwrrbhx3t3sNVWYEIkjlfC8zy5etVO3sHQn
PyZ3a/08ktacMTaTpRO556odXZtdmDvnm9eLrxSti4Ky0onz5NgLTuSsxrompHuX
QOmz6FAe9K7gkMl12gslmsSb8ypydl1pJFAV+Yip3HWuLo5O1rrYEO0qRPMBTYwH
m6JPtLRoXjdPhdGbk9bhBCPBYipWd/MP8h+f4iUJfbhwTknJTJYfX8nn5mqBKbU6
PatW4FnGS0RpKSZVhZK6I8MXGJlxpLA6d/NbEna9GFt8dzkKhmt9BE7XLPOR/hkT
FC6airYVsX7WZyp2xdxEwhl2iDrRYgfjJyLBnRdzMvIyrLTT44njwAE34NIl9ToF
9ANohV282Q/44uzyVdBdW2rC2ceIm7NqW2Vu9irG6O1waooTZ7gVm+3PdASF3jFT
WUTATemJz8ilq3z2XYjqbcX+zSbe87c5eSJBRjvgNgoqISM212DZjWdIgax9SvNg
iXTFcJrMFP8LlRFEP8NBjzDmlxnaisRmjrES7qcJYBbSgf51U/PjT2BtTebnyIeL
FkGk7EHFBXQZCh0Cgp6qcM1UCADO269gxMywJWHGXM9CP+XNkO3Yct4tyepxWjLN
R3SwC5yuVskLzNjJyzl7qUIgzA065a16wPQOv9ZnjlMm/FN4Al6I1de6LbaT+x3X
62Wv1CKqq6/D86/W466vaAg7JFNSC014uEg5yEiqRrjtZ/SdMkOBPxzDb0X8+4cs
AZOAGDkhDmybZAWx/9TLox7WHZM5BTXPpHbKpGPge9QUSqG7bqa6GF0HoDvZMI7O
PwakRHqF3zAhYQAPMRgTB/Hmx8JFL7WbXuSPCtoRhjtk4hAy5u6Vprfcljit+buw
AP/nTW+AvNpycwoLQY5CNP6K/fqlBnGV0Gcf/FIjhFyUeSiWN1/aPLiCmxXLw3WV
/g8y+JsZBZf6niv9mxakJjN5HsTrGTMcnEupSlvXHNdU+4883yiuCe+3Qc79FvSJ
lkLbeUqPLZifqrPyC2AKA2iClIL5MDc4qQQ+flfIIj4Nc7gi7cFiURe3OvuHrHbU
T1tr41BVNcrm1uAkxK0SNox0+VYmuftZ4SOtyMhgncoiNanrYxF15reXf+dCbvAG
KA2pSmT7uMQmhwg6R/X3JWjM4xjz7/vIdaaV85hYq/91x/a8VqKOUNHiadRWnr6v
zJ76gD2IQUdsxxeoR15pCHz9vm0Jxpmb9DjP1hT+jFZ8z+68EyHS4D+1MzUrJNPP
nd4v4fmSHKgLctHcdpFDpBJDD0NW+jgZDqUh2i/+NkiP/+Pbnjr9+FHV7U/2MDn1
hpsUGfayNQZ+WGQI4x5I5X4S68+X0hrzeTL2+jdnDhi3yKX0sj8qCOpemBY8X3pI
2uHBBbp32pOOBWEqug1mrcgWcbQBktMSX221uQcO0oYv1OR5Hlr1IFK0OR5Sowmr
VnLudmN3uAOaHQnFfx3M9Uv9b9iwE29D9Gi+Lr4Auo0FezGi3BcuMW30RgqwSY7o
oP0v3SLMnevpiydc/CaGd7J2WY5x+KPQVneJLJJ3Bewbc/rSUWqxAgHzDjoj5F13
X2zUv1lzMNLSiRe7Zb3EaefHt4h8xeOYYgqvGnXuQxzVp/W7dijTfkA2TWZ0AL1c
NnATWb0YNufeNB0D6mWhMDkJ78cnvDCz/K13t/jIJgAp0uCVtQes5ICPkZXU0lrL
D9TJqMfHmSVyAWlXwLvhcaO0afAO4q/8miVuHFqUe4RilWx1Y70K+LG9/+LHMbWQ
7lN12Y6JLmwH3KEmgMcBAziGzdwHwMfa7V4PPSq0f30cNEU8qDmyXmO33qtCgsNU
lBK/FXoXisPMwWPqCjov8TgRGx4r1oB+2rmQ3bes0/kk5AAwYErOmeS0lVilGfnJ
yERkVzlMpjN8kbw2pguinXqo124NgsurfdU6IIl7E78kkE/HhB1NEW7PZCsH4H67
DBvEDuCtmJQftkCpphuByc3EkozgXjuX9j37P56xPO3D+GGl90w+MOagwb1GD5+6
BbaOWO/hic28OIoSwBlZjNqQvnnjP75VqMWehv1gmbiYizbSfdN3xnjWAfoQBBEB
mqk50YeFWpltMbfgulJDl7DGwGPjU+oeMyYjWG3rmqwfU9eo65LhNsZsgMY4hc9C
zOv7GylYpq79mAxoDHwmDgjdK1LiMU7KFhPUsR1zgC7yag/J/7mpOoZTytuPTGgW
5Wz79TI1w6WreFtEXQN07Za2DgNi0AezPasStMo8LTaTWwDVQhgI4ooJqP7WOCI9
vEQZGmTcy8cAdzvNKZ++Z7PDaEKoFzAImSGlU67hRzkqTsORxrVGdBzoKTxQtW2Z
cZDL4sP/UE4K7E/zwnX9iyteOzg9Y06y9swXHw6DTs7onczK3phh6DhBjWFehZca
cJJZLYhgPavohxhAvC9SEhbEcAht+QSYxnhYw7BdQ93WcXUEIVxpWplMmkYzAN5Q
y7n+OZ034FZZ12+AAOAoIAZJlgtjsJt1FvGAgDzYG8VvwggBAQjkDQi4uHSv5vCN
/K+LT0uf7eHA67c62B6T5J2iEyahzebChnVAsKKbXLQ5vMbJZdPjL/HbuzKCJ21B
DKR3pm4wmILeHajmSCV2l+XaMB4cLpJiIHTm3L22LpqDOBlKtrhF6+nbB+ZZGyXx
EVXjmanALVmNl+8cmVFHQ30to5fOKnjcqmaSWBQzgx4krnMfosFOF9MXKC1ebkq0
vT3k4zF26JJFiA8w1W+zPWkpX1cpTPcTwmjMj7SIOQuIH9/jLArOXdQy3GKmSDhz
NrAWH7zbSd+RHZxilvx/VtqFv0y8l1OZXL/bt/LVFkqdqc5Bte0lOBUVUjL6gT4p
Z1D8BSjFeOM+VOGZUDBWLxmM5u2T23O6XjSKDbnN16XCYFOa0dAia5XBP4h9D3Jd
QLGh/IcYcaH6IY41s6rijLyMSrjfB426qPgXpIyoR9FmbyVLAAsbBxSvt5oaLxFn
ixgbbSXlotT00Ai+UlEp2OgtNR20lUSYx9citSBkLVRq5lTaEooeuwj3ywjtj8jV
ADr8zVyvah09RkmYixF85qBuQ/u3GBGAIHd8Kk3w5JNwWJbo2WInNwbk7VbwIYPN
/XfLoG0yoz13I7istExf46ku14BKnZ5ZOGjFtlwW5xMX/aLFMSrZxxc4ko04AazM
0a7v2D/+K+me2Ptbyxq2qGnYK2XJcsNIJ5EQBiiwQrFumEhZwcWp6neyLKioJJ2E
4MyvcYiXflb/ktmWoqEPCbAssOte24jgOEL5YK1a6o5+HtsFSB0FI43YMc0SW98P
cYQw6wXvQ+qsC9E71rxeyDtW6rxT/YWHdP3R6Yp3Lfhnz+TMChCM+s9U292qc/2Y
d8iUCBweiHxjTF9UZc4G0CuUomB2RpH4Uf3giX4VHM0ldb5NQvcdAPqhMBgz0aFc
WYJpLxtGJJEiYxaaFoRuKwPtSM1BwH6U/SIsQjtze8pyiq9RrgNGN22QpxGx4mHk
42zisvd44xP0GGsi5CqZezqPy/yYHJx8a40w3vszdC1JlgHpCgBoFDHsLKVESgaC
E9JPGtZB+HxrlDJqydcfwWBfYiSDpoDelKa8/awOtThp686h+sV0FOUVm6jwmaOP
dO3SSEfIdfxNIhvEYPmzSvsKRwdU2TRUx1XdQnFVc2HkjyHlVHuATCF4pgEuu7hk
N7oNad2fUgwNRwtvYF/xSYLUrR0HtlDEHJu5oyFHTskscCqupmO6KRjoypVan9FW
zcgmlEe2V8bc+MhL2xVYrekDpQWZqr3GR1H2pyOrKYrM65wOWQvksxHm09oiq+jR
+Nwb0c/r5qR5vpqzNJquZ78wITcA2GFhi7iirh6QMuZQeEBiHlyWBGRkslc3KPXw
u9LFgbUOGP4ZbohCcroff+ddJKm/sPFFFTqOMwAEEZ2FA5/H42mb4tCMc1cBATVs
Qj1KgeAE2UwpvNX3yk+5TwewPAWJbE/cWFVfqV07m8XKWdqF1QAz92uLOhR5HBS/
x4myv23bKs9ASMYRAQUqmwCJHX+RheXm8URK2y9qyXZc92Gp0M1NSQ65QWXyb3yg
v1PRBtw7PzO6Wtdx0ha5FBlsf2rJH7ZNg2NebhoarYoElmzHho91LpObE+0npS0w
n6awZx9fhNF0bk/PVLctdyn1arFdJt2DrKiGo6OuymFeZl6yQOtpPDwMpIYisEzJ
1K+hozw/GpxuWIaS8lyz/Lz7l5qCX+tGhFAWANvKB29S1a9eMrjfxsmCrk4ANO5u
BhZcNSCox211bH+/IS9o3+58WcjTXxAxtwPgZJMnf9vIFeVJFq+aA+snr69De/Ev
hCvDV0hUdjSzolUq0MAPbBKe5oFrFiLldj62JM9OvaD4KSeYmNQvfspT95tj61xw
E7pfDWmcU7qmG0kiZH5v+LrOXEHLLGvdawX6w/D4t2FsowiY8XVISzt7QtWiSVh4
lrsYFTHlKSltOeESOchgAnkmzuyLUDz5joAcqwHpszQa/iMV3CtymMJpCAEgwEq5
dDIrn/lKLgK1NGlLEcn7cdwrOENdEC2tM8zRGvlCwwwlNLJtGztG6gPbOwfk93/u
ibIDDDLmmMSnieZwQL3LBvWR2b7F1ogvGMDlOVMdObArIGzgXf+2hlrO8ALbH93S
HCypuxxIa8QSW7NHoBcFHiJmC64ODUajnkx+BcAuxgkfz+vewAv/EBeKWiUj9xNo
/aJAP/xt5T1KS+sYP/xE95yLgWwNpXR/Ok4QZfxCRgV9rI9afdwtgnWsBz9N/1+k
meTtzD+fo7kkqMhblOtDIPhdVgbcn2dpQw69Oc8T6hSAjlZNk9K/1CAFXKje5QLy
7LiZrY7ulbwy69cW+zDz2nQD64Uzn2rwPuDBYlbCzds8Mth3wHNand9aL3a4akGf
IQ3bJyyw+R93/KjMBhhXAQ/zH9Y7DZgGuQvS9RqH2h7RC0ayj33WER9t8nVBrkXT
5tYDK2Gc0sKQEbuwA/R6hdgRr8cpIaG92Suj3aSIWtATuPQ8OUnkbyDI471ynT6k
tQzupaYwdf+VRkigD5PD6utOtHggiMON1jl0G4KxVr189hzao4ZIkFKdF98WUul+
eePzks9vcV9fJINMfXNmK9ijRP5YCNEuY7d124BPBqYIqqtlFHHJz7jTUURHBK7T
6QEqBTiXwfyBnLgrgzvBatv/0DC6Uh65tWLdI06PdzXFrl7+4y7DAnmxnJY9R/2I
/bcRaSxtYIVeA/2lG6mJR+oM3C48MzSUGXY7CAsx2AfkehvamK+wUirbsYup2wbW
zQnOVhbTuU7H1hOxY8z91FsSsnUoUr9GsmZPVPjWwLiq+biYagK6Vrh9GS4yUMAv
fI+UC0D5Qmsm7P9G/zw2nHAWcXQrNAK6lRqUh/UtfEivN9BaPl/2z3fiH1v4eypi
BqPv7iJgS9EHgpknHxq1ajE+tnNbForDzQZ3QPh1ZG2mwWLNWax8L1qOZs8AizT8
m4nwttieplTddI9ucEqyX2gq0poFKH/AgZuBaLB60AIxpmB3tNiSI32EXJHSrZCL
7/pDLeuYDtKb7d4ExGwFXhMtDQnZjZ1UywI0ZNZ6tvWDDE6cpjjbzQlRcJ+Wb+tg
F47hOAlcYAoTBU1HPTonzA4hdtMBthS8i6j4Lg+cEuKiBeuCXtOhyC9qx2UuOFP+
sQS+N5RmBeOOGwN/Wbw9ddVF8EmVucFOevLN+4/PetF5PR2MGIj+Kgo0RXZTBvbO
tLk+ap0qHLam0xRp0xFFunHXArYMvc+I8XUBeJ104vlIzCCCPSRNf26XyRbdZm1A
lIY0bFTFhULYJexdSVdhiBNRnU6puJ7D5kpLIxd09zgo09o3fNrgUJ0oKEneJA43
w0Tt8b4B4irLyic5BLDlbS2QHM6r6Wj1GZI+qLTlySPd5nZqQgwpjjPUeqFi4PRe
ylv0xQXtefpcw0R/rwdeXz/ChuhWFTP+HRgSNbaK0Fg6ktRDAg5Vn4svG4Etfh8Q
h/yayhGpRjVc0JR0k4mCy+Liacv1fivW+OH1E+i3xEsPjnEeNRZYNTFOh37bMNwb
uvrJKPNdIGe9yRS1NzBMWeCQwD5mysFW7ZGWNkPeAnb9hYO4fIqtpeNCIyAkILyM
Uz0lozpV0ukuTqrzdsVjdO5N/9PcxsHFL3vSIwfy1I2I7tJq7aXeiI7FO4n7mSfc
uJLQhRx9PoRIJOpKUt+JjTZPrwhuLf/eHFypEFmrvACeLSuPEKgsBIfewKBlPrCk
wuWBZ+Wj921dzYFdKR/Pp9PHmQr9Ke4+YSChpUB/RCbpYwSbdKOZKfWIIpJSuzhf
hPWPtoIwG8kNUde+CF6cxRwq54Sm8OErvcFNLMlCPzehBFBzFSQ5mt7OsyNL6YWx
25bVy1tgNqBMJHWo9hc2u115e4V2I2IHUCoASAJs3eR7Fj/KfVrJtXMvwPOShHGz
VUAZXZBw5lVQI5/+MiLOJBEoczdcWkLTjAKSb69sGOdacuOckcIaUywCaKgWfum3
E9F6vVldaRyqp/btOUOsK1eBfDQPMvHl5rPtRdQ3t1cy+CtJnsPfIqiPErJ0o8VA
fs2dEqTYQqqkzUO99qvR+y2bpTl20L/s+KwgJzwEv27lDVcjiePNoUU00ejcbPIU
VSXNqx7twBy8xos0T8/Oc3ORQ1ly6zmA5VNCoeRPTJYv78khliugph4mbj6Z7XDE
B0gSGy7kQH+c72s6r2gm2hhsXYztrQYFsvC0srvHItODwoOTIl8q5NpUa4crxybc
UTrPqq21Mza2xwTXhUwudIcGPsRO7hhtoTw/xw8ouvdmrMbO9z5K1Wr0Lvs6j/XJ
XAYFDP6VHZf1z4LTiBjsiM1NdJYInXHQ+D3lxlCV3FeOaibQREtlrk9iNbY1mfYt
Be3besRra1+b7Dq09zZRHnVSxfXq3ryirdg+CVWWZElsDS+fpiIj5K7hbg5Zg6La
Oe2YDs2pb6wJwrQNDYO8muCNXrTFbJwahSZwFR11KGFN7Ff1F0C0CDYzxDgQsXbq
s4my6lJHXXGVinJkcL0dRaqgy/kqrg4Yy+233vo59kRisz4U/oxw2DEmj+XHw2tN
5ZI9o6wZwip0VaWv8ygQOP3l+DywH28pdBoS2Dt+PmZBwTRjdJcjolFra/HT5OTq
zUUaG05m5tUCYvwylVXqbtEPQn2dHz4J3tGiCpd3Ikr6CkukIdskJbzLiF42bw+Q
KT+l+Tn6n54oO3SHSo1Fq7qeyZwp/D4bjsw6FX2gbqzlC6ucyl1gMDKDYMWadw/6
yBBAq6NAZdt3xl1Iyg2Y9WBv6DKMlbVlYTXWJxD7TM2PARHOsw88ryFloGe9ft9H
m2rveK7FMmU/pw3LuaeOUqhW16WLcpUekR8J7I3Le2BjiTwqD+vz5Xdx83w3w92t
PURYEKS4gXn2l0b2Rl7rmvI4tY985tiuP5tfG+T0bM+nKctaIuP8gunGmcS7I4Lg
Xo3+STwFD+8tbltbhGWQekaK4CVWgMO9JmdCvQilBNR0h/glNmiOH/1LttwMe/Aj
bBGyIgGJzIMh8ytD8E7IPtUHjx/knuMFGES4gVR/5hkOixHX1F85Tmcjua27UjT3
aJdic6PDHF6LC4ERCjXsac2BewEcSuz9tOtrLA0Y1KFa3y69Q/p3uXy4nRAPvOMp
7y/c5nV2E6wanShdakrEzwd/Dr2SgWZZIJo5QH3PfPpkSgUdrDI03zC32yA5rXcE
IP9c5teYF5HgBp1+8a/xZtyLMBw5fOIXz98xpCi02T2jFdP8sTjoWD3NW6VLJ++3
NfSBUEy0mRYI3P24Mji3nWtMSn5CLajc3Dm3ymsp8u56XuwffHimz+wW5E1P+0Oa
VdBV9FcrVZjE6a1BDMyomS3FufSnOmmtdaBAnbjWCmW+c4Gug1iRInDyZcm0BMNq
q/hFqsIuhBxq4oIYo/Ns8dTijOYljp/9fPbb1m3A+8raNIVnfGVzVlVnsxaFMJKe
eb0z4pR0zSAxLY5jf8C0FTjRiB15lo4Oo8jTtTsGmJnK/ooxenC4VkhyItbO+qk7
b63mp6DQ78zWa3QGxraR09cC/EbBZIQsRI4vJDLJLD8Ls5UCGHWSE0mkkvmOLFsu
7pxRinhB7ROz+iamKp68hG6Yc4tTmKh9QirQeHlF6SGd9JDKWs7/FENuXSv6Ahvb
e5LYNzJ9VDRtqNennahl+pV74uBz98tCAisEqAqYbCMU0jL515SCf4/FaTfPuZ2y
xbyv+d34a+VhbA2uPx9Ck7dTTR7VQfLATS+JgwaWf8Usw3o3mgXixJnPMeJ2Nh2n
T2qgN2GT2IrP1EtYb0fNYTGRZKWAHtTMuYIf99mRv0oHvLdQvHczuveN50G8rYfi
ub8c8tJXjmysi152jp2/NmdFVp/EgV+39wxCCepY6rsHrBCIiVFMZEFrckl6HQi4
/4wUms44Po5e8Rn0V4FpWmxkF1kRS/GVMfEryRECXMU2Eqi072xia5pcVcpII1MX
/OfIgFV9AaS2TQ4ATaqqRQr0Uw8BP4m2gVOFI55enrJjwGVjmtIux4KbnCYGi5OD
rhsGFIX0TzKVuRpXnHlV2owbKWTsUIyRX+6sRsIm2ptzn1tnF71mVPZ/QT5dLnHK
8nGDElM290Lm8DDFWVqSnPso4wSaGjHqS78KGz2iVZxGiyturzqq8932C9GlKC+Y
bASoYdqG4T0novvgJIXfbufv9nSjn6KstLoqH1lrCSK+DN3Pb426Tn3OG8092GLH
n2V33RFOptpJTF2FBcs6n/A7ozHWFq+ekrUf62XbdOx2b7wXfUE7WMlqVL5vfgLs
NWxrqJEmOJ8m40kEuq1D29B2UcKulJCTbtS8OImXuqxtghr5w9VqYBk9VOKcf4Xg
xQNnWX77W+6b1Zrjp1TWZ/7bdqTj7XbYggNxdl5hKu/k5ZJ/qjs2/BwEYmsqXN6S
PGH7bOSqChWHdhy2PjGTn5YJCkbSk/WrroeL467yXBOXwfwldiQ2nGUntdIx+BjN
wmfJlgtesMTjAIRXZocUOJgAyuRp9u2FueFxa6B9usbfT8DHGsdAI90v1n8bqksM
FGyg9DvZafH9ecOZL18258Prb4TgdxUlFwFaTYnTgPdiJUqhVKY/i6Ikde14NqPG
M17UoT6Mr4P/5Vs2IrI2zm34k5ndTPOI2gxwbu3hT5luWc8hj681EbxJugDC994j
ZdbC/qn/DBYvtKom8fWuX6iqA8j5AW9OXRdLzpaLHbNjnO6IxCNsEYI/l0AKw1Jk
7lVZs0Fs+GRDRCvhKn4jQRGLTgxAQgGUAaf1hh3puB2+jzIM4n8EgO4P4YFNOAZU
7XiKmBSt7rwkZYWDLSG4rCtKDZ7FAGtBeS5KwJxMUOD3X/98xKTnZTOWN0UAzAGZ
iMYz9OKPs0xgOln2Hf6rexH8fM8Z5n+Sp6yxgL6WLWNb/b8G4NNEwL7wnDTgZ11C
3nsxmWC9ezgbNnnuZPdb07sZogIgqzVWUk0eMu6+nzm0iMz38zvnt3OjZ5iTpynS
NIeluxw8T+nnwrDB8nlt7JaUJqJitSZJjr9NxOY0i6iK9dP6iYTnk2+18mqqLiX+
k56FNPtkEPDLnGhZfvKVEnxA+HfxbZgF1+M7Sqa2gsN56//x56Yvml+DrFl4uTsl
cJQkpBbQj3JZZOvqzuIHY349iw9kiXBY/fjk4EtPoTnq+tcj1R5XI1pgkQagyhmH
xrAJLidFdQQAn1eLONkVDlyY2dfA3bcJbBz3P5r+rAwr22Gr6ZAlhmEZsrG/JMoK
9xqRFy6/JncjvIt0PuMWWojlJ70TsdwM5lDiSBKHSk0T8itEofcb5+Ld5qDPeFf6
E5LzarwDf3x1AznnAwMTz4KkyyeCQJC5JJr42M1mujwAd21c9noX3ZmcjKk0GQNX
gRTDJ+keu2atZRE4Mysviqa0vv+RX5PmgYCweIEPWLGHluH5s2JA9dikz5WXuCGR
RTkg4nccBZl4lEuxRnR+YlEPZCf6AYpp/gIQvq5vPnKophkn7e4z6834Iz67BeRv
WtbD2NlkASQVwr/pETcatYSHWj1LovQpCUU9Co4e4abqdpURT+5JDTAUkpQGmAJ2
y6KLAkMXMNdf7NpgEtnTk/RVIlBiGR/3thXE2/pBwofU9a1FBQKzHgAv2MmhZaV1
u68xHCIxVf23w+s3wWjumsPzUl5PtgT7KGAa2VDOCLv1n6JV1QTFVjNk4FL6N0VJ
bd6cVJS9QXiFi1+TX7cDxcN9R5x+4j0UN5KEhq9lDwZspM7KPZQSODZUWYlTrRAQ
yLEKCR+ooKxZTtUteJMXh46GzeQDXew8ynePqplaUqIq0UaGIHUaHO7psso21J6w
11KGFc1k8OQIjQdumFlP4WnK11+HBlYHmZ0lH5cEBgQb+/J+c4dFqXZ8+vjkVyFn
RZiRx75nK+gdvpnE5aIBOOrupT6/XKuZkJxLIxs2h1IS5rn2E6o3j0t5pYIYHBO2
c0z2mqY76fHgiedLHDZIsxjJmMWcGHTE+5ONWLICjZBa3DSBimn57E7SBquleRNA
2CUFJpzF5XeJ73lN6UrFyORru5zgPDDI77JKBKqWmHXiSPq4ITzMkrR4zKaVcB89
SqtxDgfBvWfY7a1FKUmt1Z1EJRaK1gaqjhWSgl9zJBRELuaYy+RD4V3Q9ZV2SLUQ
/thoM2gjrmEJzazAiI5oSyi9yjMoA2BCeOxFKRy/gBy2t3Yk7+pXWb6KmVF3jB68
rLceeDMSJMCfdF+7dRQnP069P1jsUb6blwk2nhR+vPT40D7CPa2giAHT9QWk8Z/Y
9hyjI5SdBAfu/GUijqwJa0PaeR+5KIuT/CI2yRSJEvaYwz3P4yZ5ZfKCIV9FYhTn
E6YUs8W9YUwK3COPDyJy0HdytuNlddJra9aOAUkL2+B4hYCRTWeTl4MfwxEEk9E7
NgmVzN8/Rgf7wcNRbkV1cCRGG+3h+KPZ4fHSaYdHP+WpcET7Kr9ahL6I5X71+C5a
qbB8JohG8atXjqAvGnYeYXKJxeQquNqq0sC0e2fntKUkpknbXcJ/5mdPrlh7tWfq
WvUYzM+IHQVVVosqc+EhdhH/95PkvpNCUctxUT3nP/uPTznhxAPt89kg5CjnHDDb
OIxkyihCRAhYnISJMVMyC/N8Nm+Lkbq9Ds8mJBQFDquXXZ4ba2kHXUaDqA5txjck
8VDjuCjS/gZIlsjuQ43iXdYwAmB6dvMkV7er4PG3EgwmdayWH8iS8+YnN06q8fH9
IQyJccXMsDGTywzyLIvrScRyE3MbOu+LhxkqpuqSfA3TBcOp9N0ZaWaAVJO7fZd6
kDHoKrXgn5Ghbq8s53/5Xskza9ght/VejuZIHrtJOIWScAloBGfXzilcCq2XGQ/K
CWwO4hZ2SIVN02x/36puQJrK+Hn49pseGgKlDq3oq5bhZohm+MYdyHs1iFql85gS
20B+xOycBsGDrr2mUdgmvo/KM7TxiyLk6pym8ADApZBSn4bjIL4yvUYQzf5yBvqE
QjAmBNZ0xRjjfY+Hncn7Vd2QS3o5mUFb3uMxO6KuBhZtc1Pv/MeGnPutA5QNfY/1
+hDR0NMPfb7NuOXFeBSKEnhIqBPMF/o/GVcLUo+UaEpxF3xK0hTyBgc43xbOBBZD
ZioGyl9YCuZn9zlZoy+pC6kEsm0Hk9lwn2CZmTF0+ae1ChY4y40tESdu6HDm7OdK
507oYSvDL8WC4iNZW53WU0Q3FNFgTTSoNpT7ymGO5H5AEt0Hk36zapAusvepsM4k
1fGmz97vzePiHiwyzUgoGV7lCnXnymgkyjU2EmfVsn73MgjL/6mLYMRcXj9YuaUe
tElqh3laMzyQze8UJa5Vg4EH6sc1Lv+XLmD1kzsMSdeokJssgyxdLd6kdqffKnjz
Aa2WIVYnKuGTkgIvkleTA7wqJ972kfhSGXUwxPEKv/d7Yz3/xiNuE9owfUVmxNBF
9xT+Swo2kYqs8OXfM8J58uuRP3csRW0TWSoEZlSxymJ41du49zvNsGig7uC+n8xW
Wy14qHB00oDiPhp8MpEGa7f5UXKMhcu7+Ybw08pBnDfFen970RDO6XlCn5yIZiXK
kz/4fVsE/3+aRPYo0zWZsV0bIm6Q/tuW/D4sSyVVxPSdcyjV/1ABwb7BWC4SvcfT
75y05VoE1eQ5zhXSaa5//XYXfyg8qBsep3YCh/JiZAieTc6WsniK+yM0XhKa8p4t
j/+87rPjMtWiFI8Y9nidUgxgs2FExXVH6ts0G66/eBKafdSgasEf3QYAHcObZnaa
K2FHbReGjxkZB1F5clly5E+XBjsnSRxIvExKRqb+7sqUHkRB2Jv0I1RMFTz3NV3U
3Wh/jKm0S7I1e7x7TA8XwSnmCzyYrzLia9OLxdfw+lAz8sDilfZRlQ2kAOgFo0eK
5ogxDT74MyEgmiLBK6WbM9JiFQdkMq/3tq3wULgVPC5LOQVpX1oYd58RFWvsANmc
S90ODgziEhvK2VsVT4aSU7MsEcFqF8sk20rp25nZ4gURYmSc4gi/dm+GsV+JSOfq
7xv5zTZFAftSq55I9pukyAQRUtte+xgoU/3w9qJqV4SWzuLqXPetbQbESBbGWhda
N89zB+i/1f7L4GR6STQj+udbUsyBUpY6hzjiXR9aDJTHl+khppo1bnZuZizz0S2X
HZ7M/KXkHCwDQFGc2hJB1ftOrpvsfxuYABH93Qz4Bh6MFPn9BWey7a3lFO27iVYe
srmGIRaBA5jl8XTV8TXpPyWXCo6NxBQoQpNw+ijEY6LWJNbjhdfX+19/+7NzDXtu
AQpH5/wLday2TpmY+At3h6OqbtnAGAYF6+WmIIpuEwLVbcraI56+esCgbjT4ZLWQ
uYBJ3A80j0kCL1Ju0k+49Fp+D0CUV4MG8pbtJRdqWcNVpUI07i1Bd1Dp7vh1Ixdb
8Rhrpg93GvnKKDEQ3K0kfaLkxoHUxRL5BvvR3HQ9cdTiILFiSLjSc47FsYtmJScf
BNNwnPK4FHHdJsxGDG49LmCjOGd9xCe6XLepPMc1+IOjq9zsC4hSmWMWZQ8Ol1BG
rFopcX/bywGLPlfJ03ZvQeqSJXcLn1Av2zwLZBkK+FDQEy3RMsXS4mhgiA2Xom+/
+a54Bqm2L4z7kchopLlP3+lbCLreLp81zqOGWrSpNZ4RDqul3S/4fp3znDp/xOf9
AX9GjRa2QrjsjwbI4lMWvHmFvf8+7UsgBptWDtTloPRrK5QpeyMcC9qMcnoOFVbL
vbz6vLXIo4eXEaHSSts5IkLzzVWiOIDt07kfJ5HhH0qk09B7465gwpynxmKO8sMg
Nveui3wQCX+3reMjKraZHO6diJVYfCM8luFbfqeeiiYm25MhcZVbAakZYbzhKQfS
tqWvuHjluFWAaESMTfJRtCPMqkhzHg/cqPcuy8Z/q8j5xBx6GjC2caJT5M5T3fvm
JfoYqvbWevPnuS7aJKa74uQ/7Mqn6m7z7yRt+5/At8Il042m1oZMvDs9zM1Kl253
yC7ti/BbJKdhf3iCaVkaHEp5F0YPg9UaHzFXJIhDt1kjRB5ozWDL127uRuEb6B1S
8MKtoCtK4LLwfczdiQ8xWNtlY0Re3AwwQeYg/V/6eg5ad5INk7Mo/98SIcFpTDmX
RE5dRvySzSsXg4CMqqfeAZtWBMi9UusORIAHIS8mrXR4ZtLHjP0BWgqGyF8I5lXH
RYJuFhTstXRTJfJDld6B7ajuoDTZvu0uvDH/MAOZ5CnIjAMwCYlktdfH+FnDPxNj
gT5jzeTXD8cogV4Ygbikn7Y/s/BpuEb0L/c2kpsqaWM5jUAzVD9w6JTJJinpBkUF
JGHu3rzhfKaRun99SaUYoHrg6nP+8PhdRppfEi/gdF2GZ0T1UTCoJ2HY4rUR8MIJ
46QCdynCuLgI7KjvYXxYskHJ7fMj6/7jr1V+FE0UsTw5Znu9w462iVGYEgolyx3T
6788LQX7DPGFS7tEuqNpRhIfLaS/cNl5el0EA0+nMQIk2Rn53XlJktOJbqikENdS
PUA8npkTbB2yw9gk9VtfvLj3Qxs6TQAzvtgeqSias1sQ0V7O06ywa6EQgu4nQqKb
JIakWYON6n1RB6l98KSWLgj/Q4E7PyfYRIq1mqbOXMIuuFVpfvu7mmuPa/2kfdt4
zw0ZTuBXP519OWmXkwFoFUpaxuKFe62hOULlBywbQe73dYvpcMHET3VGWI80nU7H
RLeiIiSHD3fM2jc2VRBnXqcavgF6xZqwwuaYR/zn+AU6hcnclCFbmLWxH5Nd1Nur
8l5QeWZ/GefMkw6HXL6Y5eiGLWUWHvBqaMIdjKZy5OUH4HCbwcRUDU1/QW8ROugN
6R5RDXsEdlzBOQXMrUvox9rOIkZDUkze50byxE9CQhTcC1l5wkSPe7DmSy9VV8Vn
a5ZdKcTVATkIEyIJLXcAV58fr8EviccQ/fnrDz1Pq9OLjs0UB7FI7B2viyfLFp1s
8ST9YTgJx2jOBsWDFA3Z9w+c8vT3WzaGDPRhBcfSSNac79BxRiBgqa1AObuKfcho
0vdIXWtu5CjeBi8qvAtszK65rHPufSV5vnDYN1EVArRBGnOmlXkr1/KxP90nQ6wP
pdIyrMoCUo+xndMX+WmTLlnWvUpwGMtzb45+nJnbYgsQabT2b9nCUV4KBGFQu9Pg
SdiIFfubHYvAqqCK2xmXIyd8vu08nhWbu3Sce2WEywjcWHhPokSu1vGDJjTOitUh
tTwE5oNj/Ze3d2cdp0Gh179Uru/5mfO+FmBv1Aqt7dRwlYE0NoCBg54HCRQn3a91
hfN3KH/IzkNb1aw7S5V+ndD5YEl1iQP2/lrMNsWkbQ7cXRhSIzO/AE6buFtkufql
Fi5kYHpCMM43ZTRGRENBkLpGhwYkgjQSNVjvInyF0SV9cyStJNDxIYBLa1zdsZQX
YgeGrJQxjPEUqkSH3dser3W2UGga7VJtGBogp7lKwOU2ybk9RJYGhtqIawD1cIjS
Nzf3Bxh6GzWrFL3ZoFeaAhMq06oqMcS+TN4WuJ//bwRtOZnz4OHdrsAaAlYpZBxo
YBuAK/VZlmeC9NeEjdLmsy/b7j4dXPzoFT+i3nRXUMtB/0LUljoqHR5339JudcWB
NR9q/Y2U1wcB6zLLkM55qT2SFj6KED14CovPoCN5c0ptA1JDRWGQVLEXaRXQxXkz
K3zlkBwcnCFLL/I2NyIP6P6lB5NoZtHIxryVtRVKgdRIipe07uBK7dcCZliuGDv0
sxlJQ0sUtS/u1h/RiJG1g7Y09+nhHKTX8lKiLoMg/0THwQorLP8hXMgeQ16O27Ut
vippKhyM3TdbsiLGhJBGRT83y93y126NOVfuqMn/+tU4aFKaupCSJCavo9R2AFll
C5XO8HiifYT48qjZY2/fsrXSmltDhZ0/6FoG0hhWTjEMITh8i6SQKPkzfchB3fRN
e5PGUxTz5AZmvoLc7F5UIBQut3qLAcXu1B+W0Aq97sEUggybU154qmO9IS2k7MqN
XTxgPRjbiIjz17ZmkkDnCewpdL1RHDzKmCpfk9M5VJpQ2AWCqdFo+7Mx51YAOkpv
k5o3wQ0Np+hyn8WNuq/0IU5ZSx6JJShtY3tyhWzZfHzM0V5PWEl9AE4/rqOSInEJ
hboCsAAfHxkk4WqMOsLeo9ZCVHF0Sv8e5fdG8NXos8as6URGYyIe6dE6P2ePqkMv
kKzdEiIg/zt4HIsE+ryLTOBCVoom5hmnfGAeqK8xcuV85kGT3uvtsntmtNGcBXBI
NhZYUAufWU/Rot7wgwFZratJsubHy+VU3n+sm2IU0W1AVC1XVNL8Boage+agEBpa
g9Ys3qrT3QfYYt9XsJ2mKzt4L3NF9gDdKHv4mDr7xSpPrb04ZUOck7n3l/ZP06F+
eHmlNNy+JIF2k+VP1uDi0sB4wHpISMbRh5jCKUrxejc9Fa8FuwOqeCV7KUM9+Kcf
w/WRN9xCwHCW8PRROvXLEE2j1RkUdrli1/79x0VToP0UhxNt0YMfAkUfCNY+DfAR
In7UfPP2Ypv1ic/QRWwG1ki7uUapYJdRp/kOoVdwTcrU5lPYt4Vuxeuiw4XXo3XD
/6gB8d9lCTudznhDOoizgxEdMTvqNbtvkJn96w0kuhP6WFWXx4IT2jZwPqiYl4gk
2rkoBXoPswUZXflRvbZ14C4iAejk7k5EfihoitACSRcGsTjRPw4coaVoiWSxrsn5
MGLZVXGLM/Iov50Y39Oc4n+Mq5fGNSJj7jA373yAuhbh1ku1zvzAJaS5mPEi0sqn
aszC4yMZqnzuDOwU5v5spG7iHSxPgVCabQI1UmMDBN/cdZciqOhQzoJK1SDTT5lE
5xCS/NAoed2aEp7DviNq5DGW1KLb0nydXSOwrKrDxtEc6Ih+Dqs7n3uviX5pDzb/
lKVoBntHMFvW5s3gMLrzWuQbVi8NndyzXUQ+SziGhIsm2fDYyABvI42/Qxl9EZh5
SdKxxJBzSdtv2FtaNZja2Iwt2laXJcWKFkVFNJ0grQFz6vFIlrxU7Etx/NWptBjq
OeFsvLcPVdN359OTNcHkUDuAFSjEsUuSoA8B17+kvn5vwXtXF+PK+OvRLNpylH6c
3LPWVyx0iec8Ys/YgJJHPjY5SyTK2CduLfBpllzq96Po05DObLP+tv4dS5ozZHjE
yREUXYUk5PerJKBH86/AZ/ijMx69BHqfNu9TmZDvMibEx7m3iBqyf3NOOhRS4BJi
o7GXQIOTag9MLcMGC+F6DGPJrYuhtJ+4CTfh1SWAXZIn62GVGQcd3MucHdtyRzTn
NdhQO6hP3Q+Jmg6ePDTPQPJhgIF1iVVhalUl6HA8Jk/iudIupjczH8ay5b78OTv2
UM7ucEsbt/u1jnagz5FSu1vcjcpY7aOFATVMmmEQo31F88bTRGXfUy+H7531LoIa
yrBwyo9OkQB5Oc1QTMslb0u/7Y86GuVanR+WtbEuDWSFEHiSWfJhAcF5hRAv1QFw
FUZXH4/iqv69Agl8iuRUGM4op9lF+mBARN+FXOGgsvUCehwKpmdEM5glH1Rnt4ek
Ip6xYM55D9XDj2lmPTdabl6eLKagIMySU0NQHSJTF3lFlzAE+XH0I22gYPvT4hm3
i6nVDdqdYPQNsjTRcMV6G1xzAw94PT+RmbfdneyALAOtfdHW7eD5qGkx2penfYLI
3GdjbRUjop4G/6tV8yvsKTQSe7S4Nk9gvv5ne0BEoMNcp7NIJVT6pIEEN8t0DiuN
JQhyhsFEvcVhBzRYosgjXNv70DCBbg9wbJ0xfN41y6I4LQEYdseKrEF0fWv9Qf0l
cxqqlfR/15jlpLIM9mW2vs71zTrXvY4700mnyXIQPFPH5H78kr09ICY5h7JyE5P0
QjvxJ3tse1XiH7HhhzTQX9X2/o+olXMcNowxRJ9ag5ZDOAWh4wZFdgbgm1QP/Tk/
zdZnq83uDZZtDD5wCnuodx85KfT0mCVRpkFGHFu/9o3vu50FEsGEE4a0v+3QmCvi
UPKi6Dx5LPlfYZZZIMDRnOpModDCT4RndMdGYZafpXzK13E/+egeX5KH7Cj52fbN
8yj9fcKDINUCXVwWnUVA74Tp6Q/MJXtoO5tNBawo1tZ1l/OJhwroXGb5BGSN3GjU
R/e1cyQIyhxeEwo6sPvpk9CYLCuQAYV94nQo84v263rmL7bItvuLfiASHWcdv2Tg
CYqSyHooEDulEcgj9buz8h05i6rYNAWtFPVtzqWWCqTPVSklAe0MqarnDMSVlius
B/1S80Cccft7cmjLsGoZaZN82SnZ0Sb0M43AdAtdeoCp8MJdaW2tzQ8IWDFApKW8
3aiWOFMgeEyZltlBGD1A0n+1rqYYUe76mH0mF1Mze0Su71WVPzBHLmJqvy+zMqzr
DcKSyCD3S1YvgdSGjm+ufMUQVtT/haTY/a8hGT6+uvoZFXZBDeRjG+v5HEwiUTyH
dmye5gCGAXSDwHaIAA9LibzcWZh2ceWgb9xPkTwfPXbgbne741AqPykDoy3LhPCe
qwRAMIjl/LEI9FPOFTeQ2GlkGuV/dtDA8GDJMlVznltsPHZVbid4dv1/Ox944FGe
QCCBNwCu5g2kGQ1AQ3rmsrvthGn6wnt9jIqv1DTkVXd2F5caFxuaxkKfSqhDsPh5
yq/xS5vj7eOzfjzqgFB9qojvfRxBnld5tbkUgjw2k5DGndYg40NGoVSj1Kfl3GfY
uRNirG2WbxZJW27xsXi44jWddcYJaJeXGPRg/waLJ6pldg2bkmKnZBJWvmNjBBsv
mO683UtNylb10IgUGS8m0+X/NsG8fb8/Kh42PFIDZNwWxLdW77s6ajq9zdF/ud5f
dIMZw691TDybq5AliyppBlx9DQCVnRg/YK4SmytRpU7z8wCTaagdQwSOAovzEyKh
7r5ruG10IG9mghV8igGnHhQaKja4awJmcTQ5Z7xYGKVX1/fOt9pFWrOtCQdmYTxx
7w33tgrc6s2UcbJV/mfdCu2suTR9CE70PtT6n9sxzGasiJmjk7PtLj43e82xzkRW
GgsORpzIm+2PopLMnQQQdsPaOILxfZYtRbQrtE9GuZ2+od1s3XtRfVv/dYGFY3NP
Hvktp7fdeiVc78tc9fUa8ewMTc8tIGXhhgul8VYNOUDOQ4gcejRK9e0RkuqbEfPx
qDQxzqZyvLywnjpQpN6GKuHQdfuOQsgfxrh/49Pe2r53woFioO152u9AalYorKNH
I5uFAFngrz913CaVLqlEnZCT2kR8UOKyu7FZdk7fCPk0h6O5H7NT8aRZ5GfSjfeb
cfmQCT1ZJT7n/laF0PsGfZeTDRfxtbYO7/WqU0erescTFwsaPQvhIGj4BCu02z7w
1wjoLInNhynDYHd68NC1YrZVSgUluFH17AQ2I7PfWAmDzYkt4ZwiXNMfkEMOlc9T
THZBqg5pbAzhBcxTn5WlmVgtB5ZBFfb91eISS8hhymQABXdslpr0kSGEFIwziv6K
obIXTO5APxw95/mLbgTMKCUg7t3+WS6oXyryrjcpgL87nZeSMbFpOPt9BBjzW8+7
BCNHyVDZzZ8+0xRoN5JPLzwUpMmJGryfc/kJ6GNQEU/PhXAb0ByqTcy9IOya/0BW
pSuL+PVYHBDktTo1C1mpco6qydX1qQujp9Lz1vmOcTCpos4rgx63VGKYr2DSX1eb
nWV+RXr3RZf7DYBO3lLb1dMlawYnR04CBhE3J/lOtKBXdNtwrlz+Vw5BgBL/HvTE
4ZxAPjkI+onU5fSDu7JpowNAepYFBVqM8cInPjKQfnr6KnzZ6Uwqt1tD3cmec6Rb
fUQ4e5FFHkXQ6XPCmjAPQ437Epohjt9L3J1LwA9GxKNhxTvxtrEIeEA7ta36iGy2
n9KV1AKJQ3Wd7HUx3T4m/HI6/ZIz1x1WOwOLHGvIfCRgm1DR69jCPnIkPhLXiaZS
fMj3OQ9ReqLAfQqfiRidaOPxZmxgNlJDKCFVMv1fYrVEyJjmr/SSznWFXvYLOKvG
Rf1qa0zxCdClApOwrJoZ7z/3PEvPvslrZvn7T/YKjqvBQcExeQJ/KyoPImorGatq
t+oA4yV/ww+AjLTiw3/rcvUPqm68mas1O9eWCfvrNnpB25RRgIredSM3Fw8TdnCt
359klOUkxhP2H7cDL65qitl+NCSUZMVqSlmaYXOyi4PqZIiszf3BCV51AzP4KRrH
ewyRPEyZ+z7l93nPh4G0sVXWzCTp8sapyLANVwRTgsvI9RTqaW0KPDNNPUbRLPqA
KCoV+pNJMZ7+Cg2/84rIlfuUp41HRktN7/L2tB+i9FFZVjo9qg0UIyMJSzRmix8C
T5tLo+a+TkmWCicOAjO/K7QcqBpY1+FHnFBoYAZMa4fzT+KbF9Oi8i9iQ1SYdU3b
XLrGwI++9oS4x7HeykSpaWktr07SAOS5ZFZv0Qo3oRtZwfFIK0FXYXqbRZuW0XjW
SauqnnaJYTuDkcDdNS9Nq4MCs8nK3G33qDPN80YxVn11Hn/rkjTL8Slc7jT1Sg1I
0Kw+6XC9ZwrN0kHbBX+0Rkj/O7X41tvZNBwZ4x5syQX4izf/WywZWchP0EU0pkyV
9VTfKaEtU8A3imwlrtl9m0jc5Mb9jLVXKYCzNu2bjrBXdBjInmbVQMK5hZe/Lx3p
6GMEMpKr7FHi/aDPBzK9DOksX2CUpp95IJ0/U3UNx69sLQQlZb669k+OFgNPXZiq
S9I9fEyS+XJWx6NODK3TfH1fLGwyAYIq+oV2NpGy09dyp7t/R364aHDD2Uy6+gca
tv/DZMoWapkRoeqYZYr0nv+zHMsIENlpFB23P1DQiyNO3ncvaPR/XwMjV+yECsmB
MisVDx25tu2TtSIk9Jr5sy/HAD9ug1MwrYxPOxHcypxDYNWSCQY2XGi9JyUEwYMw
tJivyBFQYDqcqQbf5MBYKAIOe22GuIi/P/A3EcidcGvzqWMISVIiC2CKoTUKRKR+
+o0nAYGKyJqInBTFobNbWDe1UOlU+eFdttgkMSB7ZrfI8nv6Nml8BMLdRfS3cEKg
HCu9i7Up9nTBOv96h2OKZ6LCh7RMhQkQu3aVwCGGsYgArFKoDk5lH0WuzSaXmXq2
eCxVuiTQEDplZmPcO3215TGNIewK62bVn46D4Gmg/Qb6jMI/2waLiPEoc4PRTWiB
FyL008fDhh6ZScKTwUzCjxjSikp3Yp4XXRSXV7q7BobHY359sf7tG8Ad/OApbZK5
SxI1yzO5m6F/oGeWqLlqBbIBHhHqdPKy3+lvkRfezRm85z6TbcQ9WGmaOQ/oHBVx
8o/uIsupUCWk7jl1+6T93CYNiZhtjMJkcCel4rsBenGTaw7BOL0ER7uK6ySF/hzC
kxNfFmLEDazE8Gi3sJGK+wxZFyBgzqWBirNEz630Xa5nt6d/6kraYjQ2HAsm3NA/
VHpptd85xhFtLi4aGh7KB7TXCWnXfl7rbWkR3rUZJEhFZ3mmu1aCObjnS3Sw+skH
xW9bkCfl7LR5TcFGIAJd7+gifH9cmjR5cAZqcI7T5M3UMYJyP9kl256UaplRgmB1
JLBoMo4z9C54yOF/BBp3nqRDgUH/0qWjyNattTyYfKx4i4TpA3N7gN8LJKSBHcCD
V5vZXfKQYSmmxCsAct3sOtgxLqwvnQjijEMFImC3PUjbxYSbG+3cD7nWXag343io
rNNQjD561cuzeV8sVWTN+OkJPdiqRu2mZDIgdPKdtNfBqvJvHQz88l5PSRFQVNCW
026uanNA02wWk7+psnH5junM/wnS7xwpC/USkro9+z65qN7ST0L5oEg1uW3mXgpy
nhGQjkWwHBHjYq8j75n/PZjnP0Kb/w04dMPNVMd8GRywwnRQsiaUFypkBbzA6SXT
kwnu58S5p/kGvq+Jdi/mAOnMTK4jXYx0oWIKG+eUGGUYu42jv9ujpL8uFZkA0V/C
uWGQQSUIEpmKKM2xub2ocIqC2/eIK0eAd6PuJe3HcMxO2t5PLJZI7xlkOXdPW4To
3dUnuzD9gWMxJ/sLjxzGNuYAqam4w13q+JCy3m52yP0ud1WibjASAhL8c1X1WNKD
oa0QnNMG/YknQmnnqVi2fx0NQ95sHrji80xUDlkDvd5ylR6JCGpAHktlJMVBobtX
mn8NT83bTKc2Igi30328HHbtkS8G6tYypJUboVsSoarqq8FYFttmzQ6r32JzfVtj
Ay88ytDYT8iJUDXbHieiWWrV2SqgbDbVym88i+dO0FhkQvJty51n/8O4vgH/OEFg
kvQJUa06v9C6K/ZzYScZHxCIo2RCwhOPQo5OyzLoGxO5dbo8PPcACmIVGB24THDF
JGwGb1wEcyGJXnUsIVDMCIXgh6z09lvAge64Of2XwqC0v+NtF/ubHa3dxFu/yJLf
loSRiRKbFCB+XIviVrwLs87w7II34SiJdcdH4VT2dhkudO8UxOtmM+g1yYUL3EyS
xX5k09DdG6pkNyWv5QYNzK9nigCM0aIH40RqNy2WS6zGOTlD8qmKm+J2S2MFP9Hg
nVjnvLnLE+wt0G9DyIzm/yWk1t1bYQCLYTD3agsHoXbeTd8M6G4h2Fa+vNx2+75U
WaShjTZjCN8ptrCjXi2kQjJ6M0Om83lKYJ764T6NxSWjAiI2+DPm6Tp3lkbW7+H+
qaKO/v+z7+1wIvFCTxjJXhe+0XNmCZd1pJK0dezBylvMfdfD0OykHfH9TAmVqery
SumbMo5OfdZ8Z4xaBs2Sy9KUO2PpecKAeK/iRiVyUzz0/reZgClY54LbKOaJY9aj
sUx7eoO64PCeUJW6mMpXzBT/xFOd5yzIv1QOcT6ZhZ/3GQB09KP67tbZG+WfZwIy
lf97jIdLCF6TxVHWorqR7wJClmQ8YkPFTRCW63QAVpap9TUF07vm9UE+uHmo1qXk
AOpfBLtspRxv9/57LbY5nZfhep1TBy0SHtVy9afDsvfr1K8xJOHtwXX3HNUXb4rj
YDJXaaB1kTfMZlxsK0CmgGopqQKKX77q6GgarWFMqYnjcjXqBHZrhwK02MuvF5hI
RVfZo83aFrIOdg9Rd/u3cjcWCNiPQ1XuRJHlUeKjhOsVs3MXFdDCdw3PiwfP+9ug
OatqJ3yM4S9HOrV2/nEzaPSntClLW1Cdv/5yazu0obKoXAcdjMsT5ExNwU73dekD
Ncz+o/2GPIK6IZRale7qPWxTHh1/wmJNmRDHOOPyQuJglIOzHqbt6SnSDU68/93t
+Olvbj8/HAy772CTj9cA4OalosKknMJ6gm5RrlbYcs9F/PgUt+Xgaie91+Lv98hV
YTQkSqgF96VXqcsqrFrppcJ/HbWqksaCe8GDC6q4BsaZYg48qibpiNZ16d6VGzuY
XSvQeblvhOo1GZBeA0LHkVVIYJBwBxKBmoE9fIzVIe60RnB522SJXoyQTD5cAiRa
6tCCh0eGh4oSAS7qS9Garpl+gZMEVJqBF2f+P0aU1SqU2tw7rUFyv9DhIlXHPfAq
1OKIa1b5WiSGThxFm7lcWTEKrlg7lv1yT679/wX3YzmFcWg4GocLN3zoDFbjhMEp
jB/qi484RBMu0KVrB2PB5qpvAvZ5s9fA5TrjB4HzXc1AcIUoKQsLPj0j//u6RqnI
1Lg9gPSvkD08nad7tyZi7lC8oGFVRBOiodxjw/B4rm5xMBa9egItH23nn9YVzmxx
SEfoxBlD6Ly004v5AhDte9XYY042U+BK91TkQvVjsz4oHj89cz7z8telWi/6EnDH
isWwHFGNpADtEQIYbb8GC1lQDfLdt+qjokc/Giix/ERFY9eIfxZCTm/juV19MB8e
ju0PYwEFDz2izU/mdsMVowDuf5eFWUbBCh1WFp5YpNPPoub7Ixqo4NLQUKKSDIlv
nf+E0m26RlrG/nvEYTBUma4XFMZ4kFXxC+38HUv/Zh5wDohhjChK+4kjk9wCVOMt
v0MyMIesQHxqRUespotF4GnLJv1BdBSoggarqdvFyTjC3dipEkWSwfIcgtaWoQpD
yV1N7Nn6CUg1iptOk6ioyscfO08yJZk87+6/Palp/nqBcKjIUmvXhXdxWigxR52M
w32J/HaEoL6Q57VVrHJ5wxjfdyK7wuu1SDQKVfXRztcsaO55wbhbvxLqnRe02sF8
5bm1LR461Q/CGdNre3SabT7PeKjL0RsozHFmCUZhQsOmgbsYDBrudVDe+XbNTh2N
QCHPYR6GMeqoP8/DlULvQySpvlh0mNyuM3EdhzWtNme1R7J3HdHPUTuIqhcK0gdP
ygHQHSBwHRr/m/9ZN++dXtGypQbonewGyHDzZTXvjvQD7bjLqmGclItM31FyiPaq
uZTZunUzal54PHAG0sQhdk7tIRSVZ+2strr/OALIXjEE2wXoxb88y1OOBKWPcIqA
XunBpKeEAzd7x8qJHm76I9wfqhdme1FVnCRa4WGWBVP0XpT2dpNFb6ROl7kCkhlh
iJLuQdCej5cC8MlkWnVs3xZ99pC1WqwqwXv0o3uV9x48A43/Kgzd4hU0dEjDBn7A
MfePyRyA2UhlaPNgmXw5b6xylHLXGVWSl5k9Cvsl+2BUa5ZQ9kiRRmSs/bGyV1/G
rQs05c66T2z86KoMDGzLmcq68+7pM+HQwyo4hsR+2OgSetzWJHjxijYAUvheMUNe
TmXQLCOhh5QAm7rSvgVizg7nKeT/O+WrpnQdID68nCRJE5BwABX86HjuEem115hS
EvXiYFaO3PW6NxCTijQsuk2+IFQff5T+3aZjIZme1UUcVOObaLBIES5FKu4ph4Z1
xQf1fGPRQQ74nE193z/UOqVOXgKJ5zq++47PB6xh4ARVunYV/VL+1JaLw51G9wxT
VhVLr6vZFIiKCfS1njPkvSoV9B/EPr8wVMR3Fjj/7voWc6v6h1Ja4c7QoX1M69iB
lKMbpB/0/Twc74H/PXRDZplxpmC0L/0z21WjTHDyZTSNk9h+yW6Ro1KBPxEVdi5+
A7/cTCIA/JRscP00ZDK0UiD6eVCxgNQsApSdQtVBE66EWhWOen6QSiDfdaaqEeOV
cBKXbzYaAfXYvR5kjqhHPqyQbNv3+9/IQb8FTfVC4P6qgoeUTd7npFy2G9B7L3kH
/Swl7MoTgzmbLsGp8KeSSEcNPwJHMa9xb0b6F0UsCa8s5DE/PmklKXgve5LMN35r
y/2ktc947j2WmeBaxYMWUPeh6z/ZqLlSY+AS9FRU/qgTw1Hq2iWxzUtg9rE4dFcQ
2yBt8CreZYkSg41dybfFHP8cdCCyQaRyF8KL6qNlfwkBs8skGBENxyKUKglaB3aT
VPvboPjQFkmSF7ycvmSaFaB6rZtgf4BGwOMDKGcFGeAdqNuw5LEXkSYmjbMoUPl5
HSGBNePxFBVwHyPfVFPeNfNdGboWlZ+a/lTvGKEQcNacArSx++Q3So5bprkRmMec
ocwlCBZX0pHLLnfP+OH8SUpzkybpVh2UJDte5C4xWY1M0v828O/oT5HSVpHmFNe/
EpwV/gDU3vM4EKObCYKmSWEKvdp9umqsCHLx0ouMX3MbfAANHXOSq7nOBQBFP6N6
laUzAsfPvaT2tVAB+5cw0d9kbEb2f7BspnKt0MfVgErdlj+QOSaNB42V/OolgTgl
6rqOv8G48RKcZPZIPNMLeOdun/IaMYTsUWPmjbFW7MGQpv1duRs5THohHAz56K48
IGMqNjDdPz4wPtBvd7eQvJPvXA/9Ax+yv/CnmKh9ZksMGYzPdrchAlrc2hdg9EXS
3jVP//ejzdaizS/YQMsfrTUOXHLM6bJM8p26TGzF4dKZUG0c4Dbd46pazUZvzU36
Hi+8YJPal9vDw+FPTHC9ba5MZJAAEHYH26FKLdVV6StgQBq7VZcmfiBYCraMRaD9
PU9694Lt3zEPirOYbeb5YFRCn5zEAoiMDZvzPP9DbsLwoltvAUDSH9MjAfD88Uit
Zp5Z80DoNWK8UHTazN5KMIG+jFd+tpk55didPSqxPo+OveIT4utUC7jtnZ+Z60Dy
hG0eJ0PXY8rnDesei8RkzSPxZjtErzKhW1jSYfIpgWqfZZYgo0nDw6eOjAbsQmQy
SP30gSEjYoWld32eVVhYgLc3rV6W2j49RFExmI6mEVUKL3NiMKGN78M7vqQihf7D
rwXHNOqyW/jCtejzsAy80KYS3PeBPjumpGpp+j1Mxv8vk+aLrhEZfMP+I1CNuFuC
cJnOYFFNBgTnsY2fFdvKq2oYbEQQMFGG5Yog32bAMzJKgmG6lJxOO4cXbIeyv5ID
Zlfu0lp1dkr/3Fdm6mGxrCSLKbg4m8EgqbOx1XFR5BtgXaYOEFGo9OWpe1TsV5P7
aTtisIzWkrWDG5jTl0fNErCmgfz37GvnNvqwT44RKyxiMw+xLfqJbL0OWr5yQdlb
aBxTfwN8hjmoLN7bjjiHvE8wGkFxiSVaEexIhiSsmUh9wFbLlmk9gab7quTzkav9
nuaXGQeieISHQf86DnBkjctpbiHRGKrYW6tSCPzHRz/fqv2ge8zibpqifwhpKiaj
vpS8cHCzEtV2FWfIm+2HeZ+ra6jBHbeP2cO9bJ79IiUG0UPupFgnL+M9MMQjn/1O
/zrV5xbxsgkXlZvNg38ZAByratNYjMcH+9pRiPFxwQQu/pU5X6OdUoFKJ6s7I4id
db8Sjz6mgVMjaYV0ciVAtGhhf8l+L3N7W3rOfXF5w4Zf2No9ajjboqj28mskskiP
uwdK8VnEmLt6WIi4j63Aw1lfHuYlhIKawVMh8+p+17GzZrzfEmsqPJyeO6OdWUR2
3pcw3KTZlwNd7W+Os0YWDFvxRmstXIXjztOs9A3YR1x8VsR4RblCsfZZHB9hIIzn
ekZydHykgH/gKeNVYtj4Wolkd69m84VuH7DYfuQOBwLVi7AomoKJsx0FhdYxnzg5
quLSQVaSMRjka9k0BlsFeki2vLrED+gkngKAXre7axZmv6wjkgh2tGk/UPKR3Rvo
m1XifwR9gXg+ROiukgYVDgiff8VVPuyyAacUr+4CwwTCz5D/6eiiU4d+/CJGrYwW
JttRQOrR1NSPbNtTkeC6BEj+8WH6TSjWEzH3OjKngY6Is1ysOfNjpTP27yYlVc89
H0lZ/2USOO27XA0DTnxom7uuiHA91CVJNa7QM/gSVCdKOyh0Psgtb9iDhsW77aGs
3XyAlHHCiPXPkPgETVbj6fQ00GI+ulpws+7W5pr1xirSne63qTvO0JUXUt6zTx/s
vtTpj+jFBrUeplKu1mWJcw0l+N7Ha4mr5+es+Qyq6V5eXQz2kfVkp9UfAnoinHgk
Y/Eth77O54oGkaLrzzSAPAsH//4zSObRUVGVZ8ZxrIMmOf9S86mxFTigGcffKVOr
eL97ygy0OJbCctwotCIXDsGAKGFAWazO0e0TSBn7DLC3W4l/38v17fa7OE5sg7rq
ScGwaijSLEuoW6FqY7gjJzrebBm5+6BENAai9Zl9VSBh4v5TVqwT4eAJKK4ZDMZ0
UUjSNUI+QXtPI/bORSNa0Z0SAN7BOneh9Zm6a/MUlweXHQSCNsBjKG9hr5IVKsne
GHkkr9U+fm9jXQsjQGZ1IWCZwSUsYeIJvZamFcRZyAaoaLm25Ksd+3geWcOIR+rQ
KMLISwjUq2YSMhariTsEoTML1/ZbpBnJE3aBAYs8cJy6edchtvuIFKlswBpxFvC0
2XmK3uYqYzudgq27Hec4Uy42AyjUjfTmWuQp2OhryhHjf8JvQF7YA+Oo0PHdC1r2
PPA+v4fRp6CNKz1CdG0OYTQ14F5bBCiZ9OznaMaagrrHTCAwKJC0rWsQFvCPmE0Z
wbioiqO99/0Wk8Jf/+/HzV1nmOxl7414m2xJtUYLn7OcJP8FjwK8VQXMPotDJMPM
tAUUfZ67jk7c8O/F+LiJMRiJqypRiP78KbLIM4SljMo0jtfDVYE6yCOKhpk0roVz
kKrQQlm7fRDlrZ9L/H6nGC9SM4S/UGDSnddCRU+VyRcbk0wVaUF+KA9yhVym4Emz
DqRQXZnacA+HkhoAT+pG+uTKgBfS8Q1nKzYg2yOSQ1ke0QJ0iYxmxB7eHO7YPF58
eEu8EvzxfQIEXBtpi6MVVH3kMAcIdVX0pA5a/1V/70KMge/vHKSV3/cuaT3Ddygi
1dXJ154rJwHxa1yiuufzcrAL79zN0U2jWa1vHSo2Y/CBR1skBpcskJ3I+I9jBFCW
E+HIHVp5ZvYSnR5w+eLKeoRigkNSLNYNe2N/7jtJcQoRSsVxFqkvC9kqncUGQWA+
mNWSAevYWNrvkrtp0Kd8om+kRbnNrEOSnsvbzc1h4WVeQfu698lTe3mYqwOzNJ7B
lWSZJ23ab1OFMcRzhpiorLKprAtaPmzWzOfcdGuqZH52PYphfdV+QZoeAOcZNxeJ
fB+B13xm1Rk8TCaZdUJ2y6QMJVIqff1oHiY28Imfw7sBVhKvrMyz5NpEOGCFMPUg
R7bAvlSMyOaFYycTaGmPi9RZ1D9Ny2Gob+iIl71WYGcUttAW0Cvqr5kZcscjsEoO
+OIbbtF3p8dKn6mRNUgQIkk0aCSQ/Ggg/GbBQXI85Vzn57BlqZdQRayRgrD8iGRL
LTjNyRs74oR7QcPvG8paO+vmBvO0XmP0NXHWsHPaFfCbprTQrDSbqtQJtdEMqQoP
sobhnxck1GLY0JF/IprPeTQmjZ5isJxq92galQoT9Y/SO0TAi3iwEoNjEW5JDtWc
TTKUipVfOxLeSTgnMRjcMmlnUSczPnfTwktAnCrfBHr48h/W4HdymvjNnkyHZuid
0fDIKo0wWouSAGld4myRoR478hhAmjpxLGOCYPqwCJCTciVJ3mca1s2I8oyYDk7U
MXCD5akO8F6HHdalMvlnsfu5yL1KkCJ3BD9QWkHxAHZmKiWc3aJ0BYECXxI/p02O
owXZZKlKZ9Wdg5s2E+/NHUfee0qXF6zu9PPxz3z3Jf/nAOZPEsh0gsNoXOheJmK+
OBgWc91Zv26YNkIK5Ly4pQPLhzxrErnywsAow8IdnVoNIwhEU6FvJKeeHJ+unzTz
iGKBlmrkYMvQNg8IaKe9yNvrwWib7lgy51N7CUQHRbKUG46ZS/kg3MUFz0uo/qCP
X5T9VNlzoeQkUw3VOxU/Pq6l/WEQujCQN0FgmbXvoj+PEAcnHsjLOXiXl+93DuXp
9zkSJxevdANRORvRfLt8cM5KOEGXMiZqXwuwTwEHSDxqT+s15nfpP1kGICky0dYx
zIPxBnijcqHrklQ/hrL+s2UbgsnFT8pTE8OrwVFYT+04YTLKFCpvMZn1F0353zSS
r+xke5psYEdggJw8SiZp0bJepBBgd/B7J3xenT8aqjWGPGnOVljak0/Qmb7zd/Yp
dATp+9Bbg4a/9EYEEc51C1VamsL61JxaqOQsTNocglZZ+Vc9NHM3CemxYZqTuzfF
UGqtR72KMbgQMV6S9R18nUjDT1VzZXeWdUlm8wP8vbXqRohfK83s1Z6JpZPfTHwN
sMptw/A3JgNQr/VZVwXA42SfWE+S+yXIsPmI/Fz1/jFVNj4J42+feueb6h86sp/B
jup1gBKGrOn4ALReW1hiZTB+6S/0EfROqF0Et3mSOLreltF5UakJsRyNMCGyGlUQ
Qur3MqcsZWkLh3aULzDVl0AKoJEYz6D5yrMoAcToPsVEP2GsO+Vgsz7rz3gCEXUA
4sva54pM1hw+qnj5lGQrE4nIwkJTaNMrxWOVOUd4nniJkV5CouK/sAgLQi6qacL9
9Y328eGDq85p9KLiOEOoNLNvVZ9XtciG7kcLtW+m37i57y7RcnKVdG0Qjr4W8A0A
lMyrTR1d/gcUCMbH5GNQvEEfjC3aw2e1RAp53oisbVnrbjuJCup63sCbAWIMOMNL
Xbgl7MUEj/nUquUCM9QF9IG3b9vuQ0LMXPmXsTMJMzjjM73N9JpI17ArssDMY6TF
CdstbIU4PApqIjiHKRib9E75+hf5iK7XR5PxRHGIjSVX21QwesIWIoMptnGgUv1/
CPPS5dcgV5d+osUkrf0sQ2msv8+rgXr/B5cacyEjMe06M6bHNUCc7WKNJNPJhZft
MKWqcx6Me3gViDp4qzZ2qJ8AQy9vww3Jc/wFADwmcBg82FH8QAb0rMNIfU14zX9Z
zg98vlN5/27Symd5E1rmBjH3+F2QWOv3+xo0o2CgNVLNyHtkRyQnSHvbvzNHKcp8
DsgaHmuxE3go8WlBqQQmW4il9h+Us2JBdIfZZO1JI4r8vzzKN+AeFceNOsuCojR4
IKkkJnPYrNULa/O3hSnLjWxy87RsDo6X6sFcFsEvoHSDasj7H/5bLiwYCUXANoub
vf1jf3jZDVUMMUreneK+E7FZQ6TkypvAMO9nMEVROR59HjG74se9f+NBBIHf9F6e
AU8QvAzpJmDEFYwLdwg9Q/GGoDFJ3663ehHUu+ovpmcSebghPDvUt/DZdQ+/MrMq
7pt+on9z7MhNTb0vjeeFAzQ2XRFX5f/p+entKd+yV/Bj2KOlTFl57XDz+bZrnaiU
VAyaEvLm1BRmK+mjBQhjZxpnjtN+tf1aS0yry+I4XBrNsh1YcM4HhI3fW7MAKqX+
xU04FiZbvfh0S3qD+JaidssbnKB/sV9LbZ8yxESAhumibcxaDEIdeTppcm9vjlHu
DP54IQ3Vd1hvkQRgXoUmFSaOqBSzTEyeI4bh6pfWOUkPgdOd2dz2sA401aCH0N5j
dzTEX3Bgv1pNDmjf34vq6rpNd9c5j4VCPqNrWIu6ie4jFT+o2N01TmY0B5t211uq
AND1UzrlwNfo6e7IHV7rGxbhgdGAvZQLM1TKZXAs2D4FjADZ935ToFe37jIIMCzG
gwCl8ycrY0WPCVXsTr9n9Pe+TTzMbEnMwj9uaLlxobN3t4La9EySxxQ9lBmCDoRg
eXVqnP+9NkPdt90v36aP7mFXQaivzK+RIfJOMeaBo7CJxUtR7ee0aRG/jLZanliZ
sOwC10Cq0eZk5vEt9qaf0qlSGIBAY9WbSX124qlfcu2ri7zQWlBDeFe1VP/w9yP+
BqQsRwpRoN44Gxe3+/LMP3YanIX/S0ppb3afH6OYe4zzg+gDnYtMbNnwbMaTpUrG
FSLhFOGVVmV+UnpONePmE+g2lbmhYBZeqgUIEf6y6WhM8qBLEM2RxRr+l1Qk7hkg
ZtL9AUkU1EUUVd4XiUsRcGSVs3xooZSNdXqE3zH19BpP2L2BHH9IWd55sa2YY4Kz
53GMfF9K49dtz3bQ5qEPc0EIK2k3/ySynPB2HCBCGODV2HUgxQB2mgwXNvRYl9z9
/mrKqD6OYA3GAhURjlJpqhku2TPMYIPiNJOp/aiOVPIqVbKk8lIr7hGNJPf4vOHX
3RSTB3Ec7b/+m5m8FyovPhBVkxZXpR6PMt4sia28f9nC7DWhCiLTOQMOS1E/a3Ca
NpEjLXgvTevCjhDJ2vGQ80G3jHaiu89rhzkZAghx0F+aVPp0qZrDnzn+vkZGJi6F
o1faaKCScwQ7hpIwsWGfxRNTN3Up9Lb0MRthZqFWimXsqonsLzmvS1w6UEN+WhXj
irO50g0mQR5GZpK04v3g8ycjXMha/utR2K7N07mst/afCNU8tKghXnsRGRxHGlUp
WHiAlmM+Q+oCKyc6MbqQh50mtitxSjaRYkAh59KOqRHgzphz3JbdyLS3fdsJinkl
GlAhJE0y7L4xq5FxM77vduCWBPNPuEaOY2Q8G8u3N0dqnL8F4uXrsU8/tgbCVxw4
lgFmULY3VyCkZVYoAxnqnIrzKvhjIH1d7ZwhpC4a4zwTcwpG45w5kRgh9+eYJkrm
o+flPik6QChQ0fNERy9Tfgl8h13fQL47pr2eT9486gA7tA8oe03TIIQBzBouMHn+
5QQkkJZpsXj6L58ks+plNSR2X0g+95m1Z2902/bQcyWlyA65qZcVIX5etX/cLbHB
UvbX9ZPmsGz6bEhtmiFzdWN/cjHsUiTH1vKluSBDeEdbLRuaDa9P7cPkx1cBwXBU
SYP4kYBCON4vZeJDM/5pMmL/3TyqFn9AJ9HSvQR9pyU7oWDSbBY2hBsHiFDtzWPk
IcC3RS7TEHi/CqjDumQr7z18stGhCHdQeSGc7X4sLSGlsLnVyxYwTR7EzmPs3wZH
FevG9kMpghVsywH32XenRuuEF6Pfklz7xToYTySjXLqf5S6t6HzJZ+LnblLh3/IP
WNlW32GNCYyD8qd6P91sDS9pLnV7GycgXB44QQZ6Jcs/oWdOEMSVXBtqJTRZ1aeT
qEBat2fO6YfiXqboJKY2KI83wBrxv0uqJp6Ccv72vmi5y6tbP3KN+X8wbx/+Xpda
6HdukREfju+sUVnm4024uGYdEcF04eVNlz7xtLHJUdB6CEWaf0VGgYArii2ULA/p
+jo+kaXj5gPrQSrecvcemHLgYFWhy+c2zsmwY2Mk+hUQAWLKvsUaw9vcbPmG9C5s
DuiR+RwJeBDMknhnkau4gA+di7zCUcm63fb7wBOMZizRZcbShFkpw/wLsa4/nbCg
VSgvio9wNXzIm24Ajyln8B7gkrYDSgDLrup3CNF8/Nz6YF+bS3/RJStCiZV6M6TP
TGB8rpuCTxCkm6A3G74Ed4pd8ihwbfPEAuueRzqQg23vcDwoyEOb/gQlhNNdeLx/
YGrzeL5xxKNN/9IzVd67HuUdM1CsVwXWtz6H5GgxF9n7wMvswrfpJdBi6YAcL+Vk
Q0j+xxLxsvJS0UjWB8h9FzrlhlQxPDxWe9mZvp1ovEyDWf23QemSxTs3xY7LJRCp
+4IBIPMWErjtsTWOPHNEiV4AwCG/EHzVgzxTaBgqq0Hna5ZE1DhPd6b/GRBJBiCw
pvnb/WkCmR4WSEwWWPc4xFxwIKfdqdQtUKd/hopzqCR4EqDzJUn13ekKvlZD2oTD
HqR3Ola+BDvylMuLqXdFYQ9vB8qhn0ApuwhtuRYSAGyP2lWEnPSzPejwYENaaFhp
rQpkWlvrZgUGNy1EXfDzmlSCXm3HDvnUHHob3JGjFduBpojttCL5GzbW0A50Armg
Ji/JyZLh/YaRL5vHyEy8PLKZWwTDJIsCsGy2VY9Evtz7B8SHBMPQ9sP4dgkFuzlq
VCCkBVdyz/Qe5hWWo2G2f+NmxIRX6yBxPxEpznJOy/iUjz4vcDY7Du2rQINMZ6Rk
GuojiH44jAul60+ea+Sv9QbUFqt6eNAn65wlqm3JG1DTjO02YE9MgwcYjV3UPHU/
7BjNMDj6tOisb0Hw5Ho4uuBQn2hW5g58H6+yL4GcsKd6fh+XkTfMfNQa7PERV17R
0x46vnjjIG+iRLbjv5QuMrNR7zi2feTOsX6DBHzPu9TmMx9LlRem48btZURvyu69
Q5h+6o0UGLRgfi7opnBsv/n5eduNCczELtK/nPM40AJ9a3k/wXDOZ4wyOvfsNyxH
czFs4z99lUhqjLLYEwsjj4KHtpx6V2FHNc3xKyARXrDahtDtcmk1AbWTk+LnxCDE
uzhy5ah6sqIBgG1a2Qq+NP9KfzBTpL15597+czs6NEluhm1IwQnWb1OyZXCtGVW+
wxjLqqwzc6aoO/iQ+VH1FeAWNRhJyh+60mdPMqbDKYoVZj7fzeay2wZdXrzhfS/I
3JMB5VN/cz7nrT3yYXLCkVOUY0P4KOc4LT9bfwDp3QfV3UDJ+maeB2YugTQsqJx2
YflhxKx/RYHWzzkxCSFjK8b9ccVyHv69tIpCYe7AZCPGyUWliiWPnnC98FeOj+gS
2O2pdoKYhLWeSGla4VjH3RddICSXEbHt1NqULHenQ6mDKMisUmjXEtgcCr6Eq8Te
6Z+hTh2hSKFQwjDwdPhkjGzmpaVvwFG3Zx4fEJjQQdUAojow0QfFPCMd+DUXIccs
KCuoqEgJobdG/qKbaPsH1x7aIC4Nw49dawxaQu1tOxIwr2AS4TeWGfol9oR/NHgV
OPrkRt4cnvE0Fr5F1z0JO9BEUF2242noJbVPplX0TCHGcUzM0ZpR1EppCSINBQQv
1HoQQjpY539cA+5Yr0RwrH6Bb5PzDJfaYBeirlGKpbeoHlGP2xF16hQWZkxLwCys
kAeaKiUv3PgY0KtD7Ua2sxNbUc1KPpoBkzXFysC/pg0iZdL3NlC5afZcFfcPJExT
T3KwRX+47uOud/pcdYy4WH4bSxMuYGvypeiItTfUBCnM3NbUw2kP3tTsSAKMiXuz
pls5ub6eVDu0oXI/mbkrs+6jKd+6dj7VgSo8jk1O8cRSXTd/tMz5IGY9CLw5wS1A
c4UzrfeSXR/5668AgeO7oPE3SNRifkG3s/6stBYu3XgKEjOKa+hh8Tp7c17uAyJA
QuZNKSpvDfUSGPBDeqHLR6SqCEE7V6ghP2WccZ8m37m+uw8CmjarX3UqY4P1gBPb
sqUgDSdU8U0PYlkmte3IpeQVzYiHEz3/QabnTsJVpmyl6b0p4TLas45uwZYCHUTQ
fLFYK5/33K8mRpLUz0OoM/ziHtznJKRlhIeZmkrjTEDxK1286Ae0MHvRGbpw5hgU
SN0A1GVOjhvzQoLPNWF0m3jBxqSKNuzAC30YpKQy0NimRiuPWNTrH6mlSDWMqNrS
k7fxbNHX+R+raxO8o30wRqMksc4PP8h4DcyzfclfVOCceNryvlN5j9HUOOoHS4sZ
6vdnmcgjBn9wUYHAqYeqNbp3u2gfHYLvvxz0NZVio73+fR/n3NeVSX1IFfkEPWQ8
uMTgiOS/TFpiGOFUUJFNL8T8IT8sglJKahVLkfFca8KHXICD07EZNzdFwCj23XdO
EN/fJJkULIzHyOOu2a5l8d+bFYzcDhOfVhztKTp9Q3vYvNQhqcxOlLIFtkNszSrV
vsab381NtJY1+N+M2Heq3g44ojg5KAt7ERRxZIqJThI0uqIh0CyX4SBvstko3DQ1
RCKZbDHbrIAu+61cD9M89t0Qmjr+90CU1P6nV8EBBEqUNbFI/RaNNOrgTg26M6Ud
8uzcbIBYtlRekwCV7G8FH0ZGAeG5g+BpWS0WMd646Ri9SAirNfHUB9YBqAsqcxAT
64tYX40WF/Mwrvrm1WPJVebPVnnw4pSQuZC1cR4cFLVWniz0mQZFSrMr1M4A5Yxl
wPXPcqxsTIRxmyqJWL3/QPtD04RU3/KwQU/KZ+hiChfHFU3eyNT6mRvwKcvjclno
KdosOMxa86PhiVOQkj2MVzexhvNDWObw8oeiSE0Ij6R2f+RcXBbwglEyp8rGJ9HJ
VWOhlrigknG1BVR9uib8oxCS0eQH8n6c92VuHgzuuAVamE+DT4cN2OXMCY7HnoG8
bfU6cy95F0v/emXVDAOXl2GQZh+DhdxPBMoiRgk1OICpDe73aEYHfkeuK30LXltc
uZd2qSiBD7NQvLWRh9VHDykGktyymMd+UTAqOGeCuEiNj2NqIAIRWwJnlegE/3XL
Mbk4OM85FOcMWe6xWU+dnux669fFgUZf1Xt1XUviUdcNIDFY0CllxVvfFq/MZ6JO
KLDrG/JYCGgAlZMRlsNFk7enlPRCPD4Zwq9/T6jkTNulpc032bNbtOddhND+1gCk
hUfqtR/1Rbd+clZQ+g/bY0Z00eB8uqQP2YCcqUxRXKwzAB49AJJ2QVwPz4DbmEpr
3whNw7cPlW5ht8tOh0oDp4Gbb1EsdWaxxKy1KCuuuZaMoa03apz9UdtmE7FL6LyH
sguiSWSBqJRCLdcX1BhPNaGhTaINHi16QRpHcOLUr1Q6neiFwPADLrMsTNtHRXOg
3Xle9r2aAaLGqhXbCQ8+TuHRJmapW4JG8CH1F8xutrozPcJiLYpj27Ky8wggFt7z
4YKx+dU93+DvttGYn5C7fkCJIujSDoxTzPLHK3/X90d5/+r/LU3UqJaToZxQNROV
MO0wfAjmWP6u9IQcjBqLi7wpQnhpKwmKqapZyyHyTBJgeSgPV3kGfy+Cug7OSLw4
+rBcW6hH0vPw4CU6QjRLhBR+lRmfHh2gHF/ZY5XzZat5W1uRoixhYDCNhMpIL9Jg
9r7BfNqDNVt6tvZVkdcnpPx5qrY7iUUg5IS6qdj5Rr1L0M2uUXaatyCHyjvXXzE7
B07PVCCqOd+5Y9ElLUnlrO31CMjgndP3cTtZa6E4gbiKS8pzSeFenUkHia+xAJlB
2TLvQtD55Lacu6y9RfrTKrg58yZ1SKImRwIO8hG8SYuVUMjdhAY63wvZj+EcLfyj
AbaGQivGjQgwyefYDzWotBY38I7HhWE1WT5v3cnWS0AMy0IbXn5mXGRZ8CJlSEw+
DBxkC6KItJnC/tHRKbjrnXQrIjGtI71BnkQHIpf0MISusA8XsA0tGRfrLhCBGkKF
kaYuBTAJAN34lyDOaot4Z7vzud/xmpGQDzZK1NnwadMtnt3nbvhxLYyYp7sWfdnk
8Q7LapqkLfh5f0WAZdu/e/ViZCFKWsokP9tSFYFe41Meu5JDUbS6uWQVKUNyPFYM
sH6div7PqGjMEz1Ra3jMMrBstDcYrTqsBSYKVYrc/GT1b+45JFIU4tQn03OeeSVG
dKVthWBejokXKYgc7+uGRCrkZVjoNU52vTzi4X/CW+GfwBbKxCVIxgWas7Q8eRFD
UCBe3vvu6hLxDCwX+DjYHaOZb8MI8ikJ3RuLOvgouOFO1s6iujUFJxF/gmgORl3Z
Y4qEEPpb4Kb5mkJKq/TU55exL27gopqCRGxaeJSfCC2tlUBmGtNWz6213uwu2btX
1Hxwnz+CKpGyXf6/rjU0warFmJhikLSIiWgoEBDyoKBCfhebiel4f81deEB0HzTT
vCVEMjewEySXGQ0UDKXaeFe4WZ1LpNaqhdwh+LXaD+0TG7jPsgrxsEg3D1pcFh1q
nshoNdbnitlpcG1j6qh2GW0Erhy0IWAbZuOiX6CogO65yDbi/hcHqwB/tlfbgLM8
uKR9m7UGtzuSZYr8z6ydyUruDmDyBSb1kmwE5gVbuwdbevf2praGe2XFgYrg4Gnv
te3oDm5PA4EIm05Sxdc1U4BaaP6j0WlUiRZcx9dIlk3OcB9EWhII0bwQYjkouK+l
yWoP+QESaaLuJjDesxt2JlIkRHGRAX7CyHXDTd/5rg38c2dqjZYuJStvaZJma+na
+4Byl4MSOTb98yeXthHoTywwa1Q64nTp3c+6XeoxJYiHA6+rei1Mf5W+ERRuRf3u
YhorYrZP1qSmccecHUeqBCE1f/gFsOWZLxrFCp/DNJDMSmCpzlhIvodCnq70oTtL
PQ1Po0YqKZBmRSeXBYBL1/DpOfQuKDU/P5p75WZWSGEQbU4QoqzawAdN3zkIa+wI
r4QJFsZFMHOVWY3ufen7uqDmJZ6jXx12nI96w/C6Fz+ViuxK2Yv5OKNE+kVQQzeE
WUFTWqD5gOvUYQb4QJmncVHqF7kQE5te0V9yB7WjJ4F7IEhaUYV0jldlawIv8Ww5
VxfMB2HmV1wpTqoxfgydmtmnqd2I0yPjX6TIcL63KUKQ/Bq1SzNRHZ7WkiIP313h
LBfIxiwmgjK2yBqC5xWh0P3R7EzS6eb3yUM3csqro06u5ia2s6CLOgZJYsCtdoXH
gNpnouGsnAS65OPSJnkv9rsoXRatBfV0pqCH0z0jAOsTjHfai7/tvvIuv1M5415G
RRcTTrM2HxQXmapMB847o+uh6WgFQSM592eqw6bg4uVe7EeeeN8skPT+7opPGzik
lMK3zq8lOblCiS1VE3QuS3twdNtnYJhXs/Uo7bACfKRxjmHN0WFHGGZcpyanGCDJ
T+ddF6jPdssuhXOi4/pdThTa9Jp/xNOAmcgUOb3wdhQy3himbKiDWbDk8CK8YXU/
SHsUhNFbPhMjIAkyFS1UauOsMQnMWgrG4cor2NcKBMIEPrOKE3KzwygW7yHZARD0
Cb/rXq0xfyRP2MeAUpDSVILf6+8f+ec5nfXBvviRy6t6XcEYsvC7qFueYbFNvszH
FUJ5Yp6+5XmQwII1SKInk9O51qWXoTfgZ2Zpboaf8hbAxKKapQ/h54JV39JUi1id
MVJoW+NZ2Tj+rU4sOg46/9lztoAe3KUvVH1v56pR/rpRINe2CQ3VpSeAGOY/XbOf
h2zO9E8Y1/vHcJUU57Zh9QTT/qFQt2bVj1rjLgny53taYHfVDF8tCNfZ4f697f4s
iNHx+3rS5JZRJBvEnScl5Gkk+R9jIGOj7pmRLH32Tm7kE55VDted5Fei94haeGsw
xZdx2rOMPl3NCFA8kJ/kFQko2IrGf3Wy5XJGQG38+Co7Fbs8wYbr3BnDYhQNZBsQ
SasSZEDXTXkdeRBEV4G7MuNXFZhHu9A5+2ClLDXiYkMfcWshdpwCkCy2+Q3O5sGK
yjx2luAJWCOn17Cik5UZNSgqyQT/ssY0FXLRPUwHz8ig87SR6iAbaIZ6X2TLB1Re
aa9VD+oOXM1X2EUsznkJLH8NEhiTN/Q4VtdL/QjSCXquom1c3oPuT+d0FdNAuMwI
Bfo8VWQ0S5Ze4SpsVEe1O5WNpAKPvOZnLmW7oM/0a6uS7HoP1+mKhf6qq0V175+s
gqarIbyfTetuFjgqctomPl09N/AU2xN4ruB8S4Z99jSuVtGK97DSD0DYLorwwTq3
B3Fmjrz7tyeMIIppOFUYJiFpUPIZql7QJtFECiYViS7Y6ez6jsnjrruX8IW4SR/L
Bp7qN66znzLre3mn5DSSk9M3hbHNzjyJDK2gaCSGrWwLRdb8HEt66QVsmTEpoa/S
AnOr1COXNfvh3V4zzX4B5TvXBzdFyR9N46IB67aFggupVuwBHPv6G/nZIk7JrUuP
ETOtiCcnR5Sjrmuwcd45/fxeQiul3v5I+iSRVYL637X46Fm7kN2YabKLsp4Dodf8
FFsWz4rtECiQny5SdWmQiuu5mZF7rlQDwmRw3gyKjAHmko2/yuYRlcl2XaQ4a+NF
ZKpev+inu5c0lFd49M0DaNyD5ITLWjeRlhgxY8gaTiHuQJUi1VKuS7QKEEaDtbA/
Znbw1aI9RDvF/n4CB5lnrGErdNKx2tHrfmf4RR0XkRto7C3Vk3tHV7i3y7mDLmoZ
hxpaIC3F/wlpJKGst3aCU3gl2Z6CIsytkqaEGh6F1qk12mPSzmJL8qfronG2QhFa
EqndljKPas8KHuc3ynwDwrUAceKYe6ZdPiqUb0U8NP2Y+osMOLgUKUCo8tGeHtu9
KBaKocfuEk+Jmi3+7hyvkm39laQKF12MqOfdNedH33/GnsTXIxFdoKhMz9JjPSWc
lk731T7XTh2HwNinNdVWQc3kFhjvWzXI3KRu+jNGn6GvxSvP5Zmz7SSW7zLdashu
k/iJFf9YuM6iZj9yiTb4cMVqMRR0tA02uEIobpLhXGxBwwfbJ8JJmWLEgyrplMa1
ppuooJ8VTkgLyVOodw5aNmjR2tLIf77R/ROFSG07taWufvrpT+UJthdxHiNSJlZ8
S9HMwr8NhlBXPtwGrjPq9hQo9y4IyEp2qt51V/PbHDU2vDAHAFKBtW7l45RU59Ex
Hx6XsMBF9gJDkLFbhNjN6ULFEwHZxOKJtRlnw7XtYcrhjNZYXGBmWztHOxBie6qb
3PNvk/xTy+0u92L9fNhjp6lLY4KZSWbDQSFHbt+tzaYCff6Z9uKp8zsAEBF1gcwH
fpQVKa5/C5fzo17jk6yabuVv4rt+lvPXbSCT0T0oDRBWihSctaQI2bfYHncD52GX
yNHBiDdmYQl4xLr2FX8a7x2cL0MnJERY3z3O4Jx6CMN8TTKZDRSYOHaVTJmw9yx4
6c2YEER3DSYd8l+J2mfQFfIQB/FUcGHY2PJUSm1AmlOSCrCoNi/1OPZw7KGOrP0X
HSQhsBd909DJSYD7L364OtEAyJgUfMHLnE05T9ZfWYpIv2usvvZZnmjVKIYTOnC3
imGRny5UBCjL/7y0GG+VenVTHZ7VxtrOq60nsSLhCHBwz4gOtaLQRrXZsZDxScAw
V2kjT7E0Z5EQAqi7tSBCG57Uq7ZZ67WScm21UTYRLWVoooZ6J6aLn+Qi2lqa1E27
FSWXfqXL1abCES8vIrrBguaylgqNoAzO4I45UUWWO20Fhy2p80WHp9I8Fnqf+v/r
eP5RZ07jc4lLXJwjKYIma3R8PS/Ux6aHYGIzG4uplNFhxgVAnFqY8kdYY91GLeUo
ASa7o1TyvZmEnZn/iJufphvC/24r4Z0FxxJqh4UjpQ38YzNrCNdYaTp4xv79cO+H
04q8rCBzSElbCaCsZ8FV2YBZm/f+bP0CzyX5VGsJwZs6NRBvh6Z2YKikC/+I7QIx
TiyMXHO+NjAvs5N1Ens0sPG34bACzAy7lz7HGmg3qONqAtimoZ5YZBKxzlBsEkW5
Q8R1kTlpqa8yNe/QsY5mKUtIGJ52fbBVdBm4kT4qol77n1XIBaBroGpM3VAO2req
cNHk6OlOcehgrvlhU54TWg9aY8pqF6IYWa6hDmjNX9WhTggpMEOotgnP8JraCuoH
7kOGirDeSLRn4uY2UyUerVwW7Bvw8/vgGN4yTQHyEFawBFiFp7424TzeE0vBfnHQ
2izdujNWAku1tLIWrPqmUG4SKVG0kYDrR/O7xpLgHk9w+pOcJUZTDAwtPCn/WOUV
6kYdaMJPpRtdqonBVZVzAWi0DH6c/QDANvC6ksSl3o6o5ltlWwq3gYWkRJ/e+FjB
O2dJc358LdWeQLKt8kvLF8Q22O/rJhHXvBB9GVKO/ZUGVXUU69LfqMXbSrTYqOsC
6ie9n85aSV4rpR3n2mEvheMRh1Fqom3XLlzUawv8M/ORTdyVyPMrjTkaSPnSg7ul
FwDQtl2pzU+jsFNmNprWYXFYppPcM7HM6bauiO2g9VMR+V7Vz1bzUxY1JaWnq5+L
1yDEVKYTRWhZdUI1VSFCLqH9Z/SArdZCl9cDJt/MU+A/vz0rhYu5/Duc+aibY/fV
pYjcTDrG7WFRe2BnL/4TWRb4sVYYf5cOhNqbb2muGT1X+7h+KvhVAegcPKn1n8Nh
VL1PhkyVuPqPNGCjPkSt6yyV8KOQZlVc8JucjGGZ1HNeTfcb6JYePYbOoELtqb8o
I7NNbM3X+Jks11TaQGWNEHNUraVj4HkiNZy7EdxAhljyh/PzBQwcxnlR7lkFyo+1
Ebb7eSocxjRyxT6eRsaRXaPbOpEm4AnohLbVuMWc1kS7Rswb7NwouuSBi/gQOjfS
je30f/5zHVnxdvjmRfLEoGJK6s3Gffgy5wNZ570CKa4VxhVPs1sYtQsdaHdEqwkB
9CkuPrCoNb20w+DZxprzJHuT52475cWvq7SugeFZkNLIhYPA07w2iWL4fvQUII6G
7NwpIIU1ie0uFdlutMtRqTA22p72ARLp/kVDCA1k2QPWIJlaoKtWRhZUge8rhEOC
/qdf50MidkkXtDf2dI2Jdgo93CYP9ZPI+Na89pU5N02YKtyAGbsxF8d6nCHOxlqg
q43mroxcWSwUMIotTuHk7+gSvarpT7Tq07xsKCyAkpqGrP+zWXR5ewjebUkk5hbT
/OsuYOoOQVhoLI5WwK53aZ8OMqV6vDpQoYegaEPCn8AsoBjbZAWWGA7AoX45htPX
7iX+ykrIqKeJ7f+CT8oGXUalnNRT9tnZUJWphEvrFvsKCzfN2f6SWbhPLjs1mNSz
m18M6Cq4z2TUdyCHPxE6ftY8QOL9btRK9FlxDw83Q54endrp9LDGalnK+e8CofB4
1p+mMVK9hLgVJ4LVtXlkD2t1tcFNN3WJdW7gs0arP0Jk9xdPb8BVwux3sJvuvF6N
bC3DzbiEaD6w8FYRsVRjiZmtv7q9ToL5rIMdRwMAOgEnz3xQB8M9OE3CtBTuZfaE
vA/Gmcu7zaQg22/aojARfB7OTmn4YVXXff3A4pPevgXOblCIFjwCP+lK/gbzqUvc
xx7CeZsVp5VW9UpmVPCgF+8DY+e+gAWMwYxP7xj8Z+PgxZJvMOah9w+kJBPmBPoC
bUjr666dKgz8oGzDQpzucvlR02JewH2GOeSaVhlbCl/eVwjGSbBnSNG7YbJyGz87
WwNLpNbE7wD+gnW/wq0cSLO0EXDbQBVnJquNeHIbMJDbR7ShzWRQK2v1a0jFOCkt
wfHRvT/4o/JeNI6XnzwFTJZvuxG+CyAFsayI2Py7NhEJ6HrhF6t98a9yt7rcLn63
9ytwKWeCHpyXhwdKnwSo4jEktgsmeTeV7qsWVTzENmylG6vFkVhZa+ldZqCnryXR
GucHajIuvGvDxpNLCuFECbIhyhC+03tF7+05vzAHZjm8HbdwTdmzF4IBJD2R/iuk
v/uAvhBJeoeqeY7wrzF4o5g32z9usXyzN9tcdPZg0ILF3Em0Iq2KQ7ktxkUL9y6A
hMu+u5PXc51mmsUwLbDP3QrpKNo6P3/uGeipNaki2WWo84hHalDd+HaD31571Yts
WI468taGneNLjSmBVmw6jF+rKj2NjTs7kCRA6S9d4/Fsaw60IHTkp6HHE26SFD6s
aP7C8m4VMi7sG+LIrMtmBjK8H0EVfXhe52VMD2bpKt/2mVrmBG33rABONH4ErajZ
Wrlr1c4/tClPtPI5meQEFBEm9muXqH3ueaP1tUwbYfdgYVE4XQpqXk/8HdGIZJ/q
BVDZMYMgsDFvtnVG+VkeHx51SJLEJ60JchrJdp7DdeEAYwex9b9faL7Qtaja+4Cr
DPa3mZL238P3DC6Wdk/N+vGWed+cYa4seKjugHXIPSe1P6CXMrFIOwxronWPGZgi
Rj+iVjRbVnwgBPPgonuVq5fTi8C0ya8tZRPpuEeScl0QT9+4iHpbO6drM6ztb7AT
+kmbW4YwLu5uCpFAjqCzVh/THS40x0IV15fPTUDCdIpc3pMjP2UDsKpAo2Q1dv13
tDXDrw03yuu7XZ6/WqTXx/ghzKGTdZfXivP1OTd1Ru/EmPVt42qHUIrpRuQH2ufQ
w6x6jxWMPEiZMRbnfC4oIEEfQ3urHKaCPLbnaG6MbIYziAB5iDRBYDXw0Z3NoQi/
9ufce9QMY/sqF7o5YgMhuLSt+vyUYCZNqAyLd8M0yQiwG9lNtOTAQ/UsiExaPgPm
N/CRd4MjCCl3rP/xFC31OzFsxt4tpd+laupPnYM3Utg+CmUFS6iWLOxL2HdDx/sy
1HyEH8Lc6+Pf0NYLCc0SmDvrf8PTHo8NX7C92MbOs+MOdsEil8I5F3smk079Mpgu
vTzwJBOZ3OnA4Mb8X90YixRrI9AB4N811CMuQMQtozCH/j2MkzjClVJG/w3yvH5o
8scR+svjKuOkkqCkXddMYSG1LcplmPiSs2B1NlNdYK87Us05K79uWBOgkAs+sbMA
kpGxvWS6icVNhT79bBDVs//5b+XCmRpXXamJoO+VX1hP3h6ZbhZf58X22XQFD5JU
SlriBARSdXzyY5fcgAVRznkmR3MdumjGm20wzE2L/t011YKWkeLL9OJY0Yuyjbnw
wcoZbh8jTfb42zM0DbsZzf9pV53AmOUAa7Wwdu8PIUn8+YpKJzQ2KZE2yVxRTZNc
Pa5GIVdAX6waJqnoYBlPQsq++VrllmEHe4ZdvHhQFcQwaQ7mYcVl0EDG1DYRrqn+
mbD0uJN+cjeDVxydtShVnq3M4pWJFPToSQ1nP2DFOB+c9uc5K2ya5KRDqFV/1+SP
6YfuMdYg03cxptEBQoKsz52whzYQ/TYkYabigYEP8E4SYP2FawGeJnAYT2sj+U/+
XxYhwBF7wBSUnWr1+OYOf07nzZmuaGgDUoA4sTtyUiAGnzIU2p44o1FSn6f33Wq3
E5MjduXt03tioBa8ukhIlOwhXSW7yY5xN5HL5A35bVptIXzS21/OU9tM1f3ARcxN
XloJUJ5seBIHyBvo70BNbh2qagIa0E1IQWRVkxNa2pSLzo/Cg46THiUP5joSpcda
1fnWefRXhD1o3Pe/rkjGpYVTec95JkElMCAqVWTxuvDAPCj0A7/47O7fjNJ6af0i
YaezZYrR65Yu6sfUmRhIcOBVT50MLcdzZhSzYXeH8Z2/yQ1UnyLrFElnjfcGpq4k
57Ihqo4ayF51q54Hb7jHuzta2oosnPnfOYwZe+l1x5rCTxolntbPOORTieoce625
RL7XOaS5d7SHGRp5y2mssTYjWe+rnPl1QTrQMlWzCaed1eUP/whrlIy+1GycWNDj
0tr4icoau2auDNhX9lXRW48TCBxx+J3fZeVI8yQXE2GCDUpFM04q6XO4CLrDqkIy
SAOHMp7M+9Gd6q3+NBo9RswTguRlJ6Vb7x67pZvDizpFI1/PhsJ2GY5jVvqsjbm2
uTijHKZ7zn083Ms+mYEN/rZtu7zluRcOX5nWiJklWfrz1x9RD9ZPRXhM/KVAzD0Y
6wh/uVFDXFHKvfpBagntGtWQmn2FUKiexU+QdOsOKeBmvOoMTJ1VdflRkZYyN+Qx
mqUKfGLnA5+Dew3xMqObKM5uR/Fu2G/QQ5aIaEFi9Vn8xLqsAwJPLmG9PNop6qGa
M0MsT2wXGXSV+udzQnpdECuge/V+MvJUy6LpvpgpwR7EpMXbPOrUmIaqINq17nl9
UrralHMx1xlFOd/NBQ8aanqsfSmJfw310a3juAwomuDOttIe+5GGsE/Nj6GRzv6H
Whlxi9xHdXIE/JnPnm9L+hseFUuW1ps4rIHM9xzRkz+Iuyl2nP86Bje5PNuyanx9
g2knpkI8pTOBJbUKTmUhX1VVmjfK5Z5qL6dPnL0F2jhooQZ2d6kjp08yD2Vl2wCD
qo/o2lI9jP48iuhdnL5WiS0V7ERDmcHjUpxP9f2Q9nmn7uYieS1DdCcmQbrZuIfA
dbIiJ1MpNHpo7CXmNpQbn7LmRjeU9HyL9MLLMYlYNYLaWf32s1j1kGdNO9NAoUxz
efe5Ekx0t54/BsrQCGzKMc5aA3Kx6NJQfNu8+r9mhDwGBCfTzYywhlEUjf9oXsw7
IVa6pmDrI0hjX7UyaYO1Bbf2aXP2WseGczuO2CFuIixzlq54bTkIJ5gpe0/Hw4ZG
aSvnFM7BN+xQLvtxMZk6zDhzECL2s7OqR/TgNVgSxXY2heCsyj+1ECM7oHpS4QTq
glLFgXtr0LwYPMLdhK4HcVXuZ1wMcW3u2gotfoQw9klmbhrpk7LL1VUwnxwlJmiC
VzmZpzVxaEHE+Gv0RovTbEcH0fp4iqy7WxDkH+WpiRAXvEZBwiqBlZiKWs63E0cw
4bMgZ7+Bg0MOilNMtdZbk8Vzglr0+GzSDQ09ykvt81rigXy+kAwCV04N36k/ricJ
JuFIF0gsw32CgTvaOq/q1UgJ70S5Oh0OgXHWE9arOsKAPvWRIdWKQLRZYs2O0PRH
ydgLUuVzh3otesdwMc2MzCCNU5ELDfQJjg1Od9HEXuAcry2blKqKK8dYxR91RNpV
xf3H+veCIpwY/exeDq6oDSLiQa0BfOdaC3b2h9XE4M4xHeE7iL4J/EPM6HpJWysG
ZQE8OpYBDZzXctYusO3hHKlhwZvQmlutfUn1gRLzN65dvMuSiRSfAB6HcDB46auO
F3Yscp8jqYmcaSGJImoyU9WImwdBskEvCimqRlKp/DxkZkRWjXeecQkEQxqsk+97
kbeRai7wkL6weTYIJNCIlL2aiOjhe/Mj9NVAzYTuTFRa2LipgHKsPW+kZk39GJM9
R6P2vW9270+kMSh671SsAZGha8fMNOiKzKl7sDyjgpeDLt4Tj//T80u3L7F0LoT9
calLl4RY2gomIb6c4fhElMaVSfoS2t87jgljpm4+AKlZ7yEsyGVPmnIrwFyPX4HH
Lm1IqVYQjABFRhHRf7/CVzaeyvZQc9xpN/L5cOdoNL304GixuwQPzCcTgBPUjZYS
kWZMNf81o+K4F/ixNBNE82XadFvfAlaVeirqdMgJVsuEWT4w1U8IH8gpt6MXLMEG
/bxp0SCHBeSf+CAaxrclGN98oI3flgvIB9ur8mDMc8RKz3ZKZOXTR0cZD3WTQ5lo
W22QPkirxcf1XmcEn9L3fIOAnKoQb7iQ3SUUpJn6sNzWgSU2AljoLhpZFhrupTlG
Iel8BsXXWvwxuB6P2nlu1bRDq5EVYMVwl2DtKN/d/ZtYhS06Szp+XHow/DIS0gjI
Kt4f0b6SsauTZfMMxYy5z3jpoAnkz58n1GxtgATUEVyhVO4nFtBerIDg7toolTDm
TpKiOUdrN5Q9IolDS238T6bMrfZBtFn723MDA6mSjUjdzy/WwR83ayi0vr7fQf5R
4IQUlrElcpZy4dXvx28/AyIiCIaE2suDttly9V1ooMvUkjMKLDKKIszqbDwQUF4B
yeK3W9IIK3KAyIpu3yXPLAzkC34EIi5cJzvSGEMcvVSLXqyud7bn9qvZFvps1mm5
M8fgChdcF9FTe8DrP4SWmFSegxUeO+Om+556SbrQU9pKUrjXj2I9m6yECwgua09T
d8QeBvJz4BtGINopjBidArhzA0KG56ij2VQR9VcjYTP3gg89cS2R3KMGImjWwVAP
ghBz6lBs4iuvB+KuOC5Sr0PonPdGjntDDi2Xt2Haxc/inaPTaXY63jliyQHGNjSX
q5HnxDOtcM2AJ1evQbJw1IACIqK2q16m20XXGwgxV0rfSPoghK17jNbHcAmU1WMO
B9S51IPjr8fOE3dOUrZTPQGgqmpmHtfx8q06fEwabx3myQwFqz3MYdaKlDEsPBoU
/tyQYd4F6d2hojBWT5liUPOGcFjc+7OD7c+3kL1NZ89vuX8xqZWjw8yQLdt3ZRAC
ibkwMQfWayM0RFfs9RoA2Jvw8N+dr+LsIu+1IewP0cSs8j03+oklBrz8Ej8ryJlx
1HYm2ksO8BbkeMfwJwymaoODlu5QMxcP7angVR7X4QyvQo3veeEPbz63CkiO1JmH
WImmNi+EIBfU/aBSQzd04njR7uzEiJIgMEIsn5lLqPUD0MhTwCubUUQCbO7BwkEb
SsAov1fzJtJJmiF/Lm38eEddvTulJFD89eqPUjs6YAIZWAtSQ7WbJb/hDXwYwUfV
WZPD31O327GxiCuSy3YPJixUk3iokZeDWujIgiG2EJEp2QvZO+H5BnM9lb77iIK4
wFFZxJ97v7YnSr+lvusflImKLq/FxzWH3z3mlcEE/eIZll3majsSgxPp4cXa7E87
GEsaId+tXiugegukv10YrIjP1C+kHZ2MpfkENbMgSJjCbOGKLEymGojilh5roFdw
3Gcw2GfoTMsX/GNYSHniSxvjuufrhuM5Q1pc8R5qPw90O8palpCQgx/qSsGvxRaK
kxeq8r7mTJmHGg7e/FmsS8gbK8a0JWjO5uLjgLXplVE/miyS+rWCMZZUN44nxj0u
d8YNgiThm/rB4HXPWJ/IJJD+7ljopUuC2fDe6y+X3cvO8OsJWJsPnYARaj3qSjeh
wnxFhkiR2Yzdg66CUMYqIljT35HT/sshF5RLyYDwY4klg0eLgM6e7UU7Srk1HaKt
X+/g3c5TXhoX0pxs89zAGHYXxTfUvgDPNm42qOzZVXJ1bgNhtV7qnGeosXGFgKoj
+xd8eKgQGzVV0m/aJkobC8N6rOmX2aDM1ymau5y+6c9EjbMlg/WYYOqO+3Z20ea9
CHpkLzmMTeOxnVtDJhmQQRc8fsyQwqoQuZ4iK82lQOnYvvzfit4hvcH1tJvk+9uk
DwlmVPLg2V+tqMhQWLDgYL3h1+fQDvAWLpdphDrGjXtlTf7Hx4kXZHx4703TfV69
WovlTHgSsReSZ2RwVTNuAoUgSQR2DFnZnf68nXJhBt6LNJNB0AUbR/6xvhVxFYXr
Zl2gpmIIpLR4jT62jkh6l6YzRTFs8qfBT3GBOjqwEZQpWttuS/n4LHkP0ogqSSuo
2jrK9EWmWAYbuaMyllwkoP4MHUROc17rptG3LuU/LLZlO9bMn0wMzpOFkpeIblW/
XP2WMwuJADKbB/OUbaD+eobA8ihJlwZAb8fqp1tfoCUVCYV2RPA4lpTKjBwDtsUP
kxTSVYSN1NqXj8j1wfSHXlUhqeDnAmKfsSvLRdW+daHhqaCrreGUlgyuUvfEa1VI
h+6GHeVRpRGWmpAZwmO+gwqOYxgRwAR9SYwv/8kx11H8das7A/4i1ufpHHzQB74U
SaXwJSaRGrulRmZSYUXUOW86cu4hPOVd5czQIMfQqxWw00L0y+D4sZhHZYxSV7CM
dXcjj2s1DVbu9DSAF6Nc1zteRoXrwo9h65PFqkCVoyNHr5SuLbuRzpmypnKSkdsu
SVm2R0YldIh41fUa+btntXncF1RzzRH6Nyuu60VK9eabSQZYbHvJ9Y8ZzvNq85Vu
VQMkL8cBuvBVTTdc7UMjlWh7G0t89hQLoTLFbbgp4OlRoaJATKbwY32tBszF9pWE
dcekw5srzBDwgKivAzontIPC99abG0cSjinBs98rSDUcXUrm7wNgytSL64qqtIw4
660x6xXh32F6xMGhkwl7FBtBJvpwwYzneYPbfZFnklOM2gbvBHJ0q0NFRTGWCfUs
kGeWFT8XX/MiPPb4HTbt2z8MIxFrz0rG+b8sH42nJR4+2IFJZ+BnZRk6yPkRKTPx
4WnhlDvcSp0HAj6Qpi+kb4vDqjXpo+ETwCpLFs/nou03PvJofWYjQII+FdVtsYt4
GOg0P+YBAMNbbdt5PYRNvN3IWZOdCy2BtRNdcGdyvPywpZPcrj2w4gntrM7ui+te
RQ1BZZH1ir1PuPg1dRv5pXOpc5KFW2CMF9uatX9rv4/6iYjDoGbv94QmfQfGN0Gc
FLgTUvbtqbwGun8N5xzlVz+Cwzy7U4aHV76Fzn9JgojxuuWmmN5h3TPo0s3XlOwz
lBJtRFhEm0TK6EmpFZ1WNwSXWZYwopuP5rYyCNFsZbM26fD7NhkQvqKmfZg/k4OG
Swsl5pII9WGP6cG8zJS7fO8+yeeVHpFQJWlk3If+Uy5H1qIGhC0qO/v6Rb57YtHS
4wlENgx/cvu5Ma/N561we3JdgtRbK+Fb3Q2dWyB5rtGtO2QtamH78orl/WW9UulG
KECLtYURsugf54QFB+olwThs/cQAyVHRPworYadG8ema5b9cgOx8cMbCIpVOfdLZ
L/oA/c1dAgrttF/oxc6uuE5A6bYJ+1BVN4IbMsJ4PNiT/q4I3sFbGl9W7HCjJx+t
nJLO1+tBTGbPzW44HSD+f6vimCyl0wCj8kLJWJSvwsFw3+fKPW6pTRFlVsBudbq9
qwIGSw+xnfTKzF6j6bZOcCOJqDtnt+NFcy+GkKr6WOgsqwrNOX+mEGHoYU8Wt3eQ
4gN/oigFaLpMEMs/IlMlY8RvmrC94LDq9zkQc14eSW+SAxoDfzvq7Ky/52jV75Ek
HSAlUkxBbT7QK9BYWInDYr4Q1F2Kh+DHkJIe0mwOyQYklPXW9jfN1pQd+6nqcBAz
lDcgeGIQnql0rluG4BjNTSNuqAVXwDkZ1akz4U7rWn40xJrihbyGNkph4BcwezWF
NisbZaYq/FoBKXrFSYAYcT9hRmPIqxcsdCoFA8ViS+gPALu12OdOBca5GxaqqN9r
M+V42BGQrC1Q8R6gEURU0AtpU4SIFHrmkA5toih6e19G5UKzhHk20dJLX3hbWBgf
3u7CB5kp26hGC7kOWD+qAr5YnPtktT3EkpxJxoNJ/d4gRGmnKlNp/B9wANVUvho2
7swBvTAFvKK1idjGzBdhhKQMwln2Zi3RvnvKtk631BjzlLKWsATM6xsVfqcaZDm6
LyFaMqhRVyc1IZrhWypgRaD+Ns1a78mBcHncIAO+9YdvDxk0WRUJ3aOtq5zz83/8
GS/b8+Of4xHyEzjbcvKwPYTOqct32lTAIloAo9z2H2Mo04Ywfr4LwAFoYun+MiV+
Ew/ca+RegAcC3k8pXAIpkXoEGsH9KA2VVTdxeL7P7GZ8LP6KLtlYdhhrh9nWfDYX
tjflbhKS//JYDsb+pg6D3ST+Mr8G6WTp2lHZtT6GPeRlCD91gv0gTlvOj8rC0t6y
7mA97YBzJjRnIEDaruE1RDY4ba8azSZFtSBlYkzfASatGCpzwvgXtYTY6eja9IrN
oaKOD3GbnIgHR8+bnUhMYZros2J3H6MLs71CAu5MREAImRvUyqhwJ1OQ/MWh5Qqx
qF4+2Dk501Db2oOv15euM4nlsfPGKFiok7HFyD1VSx+RgOSLmmx5etJ2srBeNWxW
fhqHzPDtBhT4VmbQlmXWyYn+yChqim9KFYf6sIGvoUCkilHTp2eDC5Smempfovkh
yWH90QNOKjtEtRlvRU7PSo2k2dpm93EhDylSpRFxnTV8nuoS4xiWWBo5Q3BpDSo1
/2LsDsQbsbofmSIv1in+aUwziXJOyGc3SbJ1BB0qZn1PSFC89LXmNzP4DvtLzknO
oja80+wZFK3fLjg03gqNeJww8YLR8sVnRSLk1h7GhTNYBGtVOZ7MIN+kjV+MND6C
tB1iJ4EAWjE7lPsqBespAsCzkRgW8TBj4res14brt1GDoQbvyoQRPzJwCIxKUONG
AMNyERU6XH6Dvf4nTv3dEvZVQoNWb/Iq5ny6tic9xF55xrLykrlkbLQs9MbGWkJH
nzsvtrHJv2v/I4dizNV555aOnxoBZKxoVhF/ymQLcfxI8A2lwUz2Jn7AaJ8HySo1
HfX6T5OMqeYw55Hp+htuY51fFm6NvzaNwB8m0KnLHHASfAphDh9+D/VCXxYjVJFC
5J1e8MvrlIJ0p7PXs1+9iB6jiSaiTXyA6643AKZ7j8Y/r5QGoQx6XKGU0m2ThQuL
RwY3PxSEmocGRjwTsP+WLVbA00Eh+jbote53btu50DE3qYF614A1F0ojNKTljbhj
wyKmRzc1GopGQE4Xc81x0+Bqx6FEwHCvh8sX+w7n6L7KO+h168k8Fy6aV+FZ5RO/
gcN+roZCf1CGDOnh0rGGyJvim5ms2dkKLG3ogFOVIJdJ3gn6tobEo2m29iUJ+gCa
KpWt7o/WzC05jnxxvuX/igrqz+IDAgPuHljMx3a8oc/sa2+YbYo3HjMzTDw7bHZJ
CRcmOPQ33nXdGco+PGyBIAC3CRngYtxv3aBXdVkAXrzEzY1IMwJX6I66Wim6Vdc3
gfVgW6oXxZwIygzRDwflf0s/awMpPmLcbmGIbJWsPbrVK57zdPwWK5vmKMaQatrB
7/6LoNqWgbPtiFVO2CFDdr24Xnn0s1ff+jg+tBtT8AW2j08dt2OOZt2sQoq5np8o
MNGiM7AJLBhDqmItlo2ZBM9I8+qeHUuJK3qmTKa9h5FKUOr6VLZVvThmgHDtjSHQ
u2rGpO5mLfzxQUXAWJ1jF98M2V1NJ1TdTJncO8ME1Pb6Y7HeDX/NVABzSWZTMCs4
G3MKr0tIm0MN3oVigTcS550otpASKiBaiAw+F43fve02b4eiQlyZoRgkbs922Qsl
XWT2tlU/D1XdSR4Yf9uEId2/2LVOXsHQf40NqaV9VmGrztKTsbg8CQMC9mKOf3Za
mx8idn3q4CvMP55dLeEpm2+7JqubGp437B2vJI4wiAbvMsVZumZdgK5WRRC3TS0f
hewNImA7gogdg8jmAoAKFd5CQQHIm89SfUy7y9uu8SAtMXwor7KA0IqPVRNjwsV0
ZV8CbOKGA6XS5srN3pUCe2yHG9/XDPG71uMwjCHfR2kQkCluVHFMrQDrdMHSCAku
1sTYGQ+AP0u06NJwo8asXbQhUe4/ehIryXQQru92gmL6b1KP55dImv+ATyh1pvRP
L3pn714/jGIF8si8Lgb2Y8TfiyCH4H1cQf3DXmBsJ5+7W5nEvahzU5D7DRdme/EQ
o24LD7UAH4g9xNzBUMLdgOxuT8PngA78tfkDqGVsnDaEvtd/W79WTCanye/awLvq
L9/CPzg6Ye8z0WmJQT6RNWK9AOCibuAtY2stW+lHX1Ys/aIEg6lnzxa5wxEkiL4z
QXl1l2IQpLQGaJV/LTeD+3ZryhOJNcFR3DN7du4enGUmtUmDkNicaKnRie8Z15K6
YwX1O6TKbimMq/r50hySNYsndtC+82xFSOBTt5IPfEn/XN3RVKJu12ypP544mz07
A3+L5X71VF+oIdJtSD+vywPaXlbTV4kkPfbebVz+Z50d+zZD/lPPwDN4KMsFcdZT
TkOti+OtAZ+3hNuptf6QcGAktg5dqFzqMQHsvff+LtR3tzLgapuDn8gwg0zXfbaE
T8SVop0Bar+mqMm55Gl2s6GLmxUcKz3XHUj+ThscghDIOz/bwOKrOIOBMQHgL4yT
6pDm923LOrKdb7/CYq1BvsKHWc6A5LCsVPVkfIKx0gqEjNxE3FiO3x5toU3jjfM5
LKGffTbFi3X/4T0UvJmhSJS029o0UBW+TgMv0PegePALc6hVTzelr0UJzdNimAdU
ra8TicvqM9PbYXaeq+YIQFvekjh2qfPG5DNrVPlqaVEvoZggvQ/eEUTaxXenaIvu
EwJNmcM9x7adbPn/Og5RmbbFLzsR+Og9TX43yX49LlHMY3QQOAj26BTslkizsopC
f+booNFVyxDBh3x07zhxcjory+8rbg5a1aRWy8Nq4a7RPFI723hEI0XB1MzbSKgc
CPxO3ZKXHR/R3pCCudBs6Io5WDQPj/+L/1CdEMZx04ftX3d6nCLZhK0Fb5z1c5EJ
3FtWZB7IYCtplnic/Lpy0X1MCDzutYx6nyLJ/pJ9Q+GNxQxnVlvY6npZtSEQzLPl
TX3CTvHmQVnj1+G0yapUkzt2IW2V6Ry4ueSFWSaLcuzVXuoTEnfv8VFMVyWSRiGL
FMii+tK5KdUDbfUBhO9i8OVH3g2DjIIUYAymzKuUqp8AP//E7jS5241TcHu1ARSS
FDJh9uHF8wlMkM4d9acRabrEyyW1b10cGF8+hsNvnLgg23PDoyqkK+y8Mx86PiF4
TCLhCsaK7+azXBtoSXtsR/xrRyWKXP9GJGyRItb5Oaw/GLm6e8Pc6WAMhDUqppKH
YnuNSqjO4bmvtwfhsO76+LycpQDLxHWq7UB4BU60IWGiCYqyBaPhmJtJE0AUxSyM
C731g7juTxhpebB6lynAhZ/8aJaVdlq5u/6i6lgSjfITCx+f6BxgcSp2oVgYTXY8
nSur30toLQlBNsd92eoKQ2heNndiAlKRCKurmuqahG3CeZ0VBUFVcSFQU87vpJFO
+JeapkV+kYV+8r3V0c4weimC6BOEngqdzYRC8D8JmrFDf0BHfPEKungkrwBKKQKl
lhKos5li16hs1fWSsonMo3VXNBYjTqMVEz+5vaR7SFnJ85UFaMSgBSSTGc5u1vqA
YFJFo0/e00lWNE319XTA640ypI11uBWR4Ub45oLd62tHltrhimzAWOpzhzYYfztX
+LdaIHIoLrC51oxMKFnm/anaZhvFCa3Bmns4Sbdt6EbojC9BuhwoPxixfmJTn2fI
JD6aFceWWcN48ydjUEm2FvrwG6BLn2+DuwwigIlHeExHEt4z/Z1rN5bdTjRBg2wj
vOc0m5NmRdVrGpKExhfILJAVj58YnvnglWFC1goUzwwR4DbFzQ33hnIRsUc1uTL3
t29ey2EXGv/ZVNNvSscvhzz6ZvdfYXre2tYCXcPLl3fq5sO0cc1kE3rkqXpqOtox
NARX4e+4g2AwBCUlon+zGqzTCAhSFAzeUM0utVg0RmU0rJIFfNj0nTthgctUa4bE
is/X9UHoO5u9Et4qY663IAAQVWs/ydzByFH/VJ9HWHgfrtbucdFWkUzdlNk16SJu
nsfge1Pev9Fbdv9ZkcYqsQMmXfHeynzFSbqgLBljGYxlmY0MAnibq+02tIjRmjWC
vFceQzAeAvD4l1hvuL+4i7wVtz+0S6OBdTmwRVz4+hHtqALpXqVEIrFWnAA8OBDf
0I+AjiBDwk6ZdgInIp+ffghN1lnQmuxzqMHlGBb9g6m4K0f7SMTLLPWMztuIrCT+
LJKZH0BicM++H2O5WT5YaUfx/ACnQpe+iWwwz2l3AhrQP4Z/jo0XhpSolq9HX3hI
t/NRdOk+ON9exgdqB5hlIOOdnNu6cbUSf0eUg/9R7XsUkZqb+MX9rxF5btuPgRlB
DzyTQ/3RN1IcXy4OOCfEY6uMihNdqQNuMDE7YWNpMOJZfdeD5Q/fdzsRIZxEVFCF
/nkgQow1mIWnClwdn8l3g3zJl9iaQuDCuWORE3bYpX3UOK9i031KOytZ1/0qcoee
DW3xhDa5xhd8JQxnOlQvdIyVbzg7lo4yaQc3A/jYfAtPC7hZBIh6ghpjlw1t5lrR
2VV5J5d/Gbfm8Ed7c/mx2zRA1u79ynl8mQnEdflcQBah5Sxo8B72AxJh/ZD+joaX
7vCRzBpSFgdc7m4KEE48q3BnUeGcSqxnzDRMfLy+rz//4p35s0We3sGXjWS3d06K
eZg24AtcA392X8mz0N+ADpKzY6uEgB2ipC2nh+S2nVi9ZjWGDtg9v+BxIVlfgj4b
05tA9XlC9o4HTMhJLAHED0aKEUO71JjcFZT7aEMlhiB4N4p1WRB8uvit+TrXUbRv
MeTupJX6ory/prKKM2UXeNBTuctaGUCCsUfAxZrxZsfQr8+5liCmJyweJJfT3W50
zjgBDpx4DKzUthV4Jjk1d2q7zh/Ajohc96AxlWXbGKaXzSHvBP/vSryUEKUXkOX+
5vaJPZ72GXdrVqRO3TZfXxmNWGmyNAkEqsyz/zjtP9xytfCRDvmkjnB/7Vv1l/im
m8eMLqczAv6WwBe9jMAleOiNHIFDh+NQiyiVIp9e0zzKbZPu/ftL2MbDTX7GK3ae
9UtsS4z9tdsnSOCOtEZdYawkdPs5oJVrIe8WUbCTjXdb45+e6h9KpslmqbQ6nGDZ
kTullxoH3iUE4Eg9Otu86XJEd8RADUaLKWGzdRSUHzhdmT5qFISq95UPX4s3a6Hr
sVPl3OV6OqFX6QAGkNmxxZ/TNUFtoH1BJO6DadWUc5oNiIm/UJIb43tDtolJSxhh
58dCZIH9FFeyN1CBll+OevHJCPH5NwTzsEKO8+SAywAIQjQms0RIjcy1rvl+/By3
bh8TgY6xMnFEfmOsx985L9qNPIGoI6SDzOSqyTwZHt81AEwgSd+XffbzpHn1k2vn
SZmZ4cWCBHawtX5LT2Zgb8ZrfUxKkJsLmZDIxhHzlXqfL0yNKgQcHVdPUbqcKLKu
3mGSWWqyAX1fq/zuj8J3kPHn/o7qgxKsOe0+a2FRV8GMwUutFvjc4SkuPHKvkkAn
JI+axNdXSLmcU/z4kFEeDUn8wrQxeRl9j1bSjgBzkbLKEmjMA68ddEMn6XLqn/1A
hjbJfo8Cstg4pb03GXofh+Gu1qqD57SST3z3emSuYSePgtqjeWVCE1Jbzv7pFv7v
GPwMOZSh4MC/vd4n5S3Rr506y+bTIeOecGCuybWilBcs1mCyOYgQCE26eeHYkgi3
ovp0SZJ0Z8obrPfyYLgu4+znRZVbt3LeUEHdrXxeF0nkYpCGpYvWZOQD97zzA2Jk
526Eu4N8p12J14QeImz3lNb8Nn5PSNnsH55WWRWYyG279yyBPtkdLLTWcIrYt9I+
0WY4NsbBNwKCAX76PZYczse9jJS/WLLLr4P5LaTU5a+leSEZKORq/J2QUQBeU96I
ETEKRQMa1ZUuwqE7K7+35XDae3mjaODN/A7YrnILhQUWS5mFq8+HqDv5+f+eAubA
8mig79mpDKndL27R1eE053rh/bkmSVYuyd9Pw1tGVLq0Z2+v9bebgqUmXMAoQDey
Pqkqtw5FEWgCM33C27xseDYiAvkZsU7/bgfgNFPITRI89EPJmcuimhQYlgilpujb
rx3SmpfxKiCHJYVYKSBVPmMm6rUIrrMN1mc1r0cKYKJdG4zqSpOz2hMrx88hmj40
KAwt6YrYoO8J/Vmlk/lDIIfjnoTVk2xlUcHo3Z/Rhg3QinGd8TLJyldIuQa5YntB
r7E7H78I2Fu8Y7p7QqgOsV57hw38gNDwiOdljUGN4C78tVtGhGTRvfuVWkWChhbC
vXyYXgsmZ+dAGufFMNlGarMCZiA4pECncfucipkCMS3HGbZuJFcaHhyeeQQ97Nd0
W1BgKxdTkqAIj7UYMjL2CZwpr9ZaBiP2boGN1SBZb2SQrfsmMVaU4Z2BnPTR3XdQ
LYyqp5PKqHlXHl9684FR1cOrln/KUXXFcTy3pQbcW93YFyLxZ00H81L7JBLyTC6Z
4uaJMRojzoCHldNLMhLMSLDtNTBvZF0WOjHLmQGzm92SiiVd+K4x2hjQeCNodBwF
TzH4oqO8Afy7BprrnxQNrDbkpz/aJivbZruO/jIYr9aF16BXsC8r11ZmExy6+XYV
CbZFs7tWnV6hJ5rrWBhBejoGE4cEv3FmLO/+CSZQOVkPAOqr03ZKWWOewSGBsStH
y79F22JCcgkXSn6VR3OX/2QS62zJYhAqKOpXYZ4+xlnzReDYQsXaTHMZlD658YlS
oPYjnyop+BtRmuSEsokNPdN7l57MxZ1+VpCnIvgJPXEXj6rPEkC/ndfEPqAcF7br
bSA06YzQVyXXyyVhgmG6tRWEFo+h5MfSFNCJEL5aKLW/6g8CrpMsOoHGMcuoLzu1
R14DLO4uPm9KrXjVviKdiDPTL7B67MgLtCVIU/eFuZIpwUnkLQ2L++4GLcVE/Bhu
d30xleeqqtoyMAECncfuJkxJmj25ITV/L3v0hKeiQeHnRZR+9ULurUO0e4Ntkw3j
0HFIuwEbVFGGbFmG6nJ3PnDZq4Nmv0ROYF5JMF2QKTEWMrcKD5dxK0hDd8sUWfbx
+llp/DX18gEIzN1OjqZCnlFr00ouoUYQ4Qi+CLdEvfgLD3aLfM7uLBQYCRh+0Pos
RWIBbF29dYVUktWaRcComJOcDcSJlT0bEBhOfdrv0wINs55YuOMxyDWOy2UmJYK1
f0SExlA00ZivupBj+08c7fbqO19YADWBa/Q4iOcEGfEtuHmQbOMUbnaorbp4edKa
CVWvpQJPlgOAzoBcwvjpUGz1Qc0D350N65dJonK8++4b0dbkIRbVYwIt9JDSQJGC
ur54nNZUKFsIU/9q2wKFRia0AO1/uUZGIx34g7EgdupWWxWH734JPnhya+MI+uUv
tpTfzfkMsjSu468WPmJtaIdMAUGW1jqTxHtdW+cBqUIEbuEcx+5BcVlTpb51wB+U
F5WTesrmrALB+8q+7qMIWxLxD2G99425w8w5SoGoNI9UzQMXJUAmfOSlYfyUxV+J
e0aHXs8zKgvT2GXuON87ILOUKWCTsvxOemUPWhPBqSpojgvUZE6xwKAJ8Z0U1HPU
do01ZPd/lZIKlyX0e9jzgur3xFIq6zO6U0pFxwjwkb/BNHfpx9vJuN6onG12duLX
ynggI8Vb+q7UqCs7L79taip0mXFL86cGvT8oH7OPdar1dFG2Von+CXIFYwbBU1nm
GLWzTR+4UIxZKL/Y/am2l/z/CVhUbpInJU19HsfM5yhowU5Db+8ejPrCpHeDMxhh
MbNRTMk7e9yJR3nGzUwnnfUerpYpJh9jxtsJL8hMv9+ndpGwN6/803dgMHq/Udbd
00KUMqfNnvThmistOWOppZOxrMppfWuDEF+2i78lx/x3Iv/8xuTpGWWWpRWpSNQ+
w3zTASYVR19BDO2BmyPZXGzei4Ja9oeCXzGwb4k5dThlda9/BAZeeTY0Q0Dh+2ZZ
EAmegRGb865J47N4baRqFKUERACkIy/hYSVu6IUbJGwH+yYO0UUIoHouxUYeGJIp
qvEe2PqNsvfNC8+G2LNkxK21CA0VqbVyhhY/3Pe+lKajoh4a5a4EMfQ6pWXPc6DC
itcUlZCbNvqtjys4t6EvusoB7aEhaxFTw+6aVrlWDEKMRIH8EhXcab1ZnOk4XCZr
15rUotD9ZYArudOL/MyCI6oJE6pvuo6rXshpxs/ULLUKviVWAatrFinpGEw+tuZj
lIlaeUqOCxUahOTY7+2NrLiuvZcHzn+dIN+w5VKF6JwQ8d7Qz/1DEh7K5BpgmlDu
aBsTLKsICVOCCkNh7lmkbew1hrhG7koMdnNAhulkpQ+LzZZrheNm9/NomAUu69qS
28lm5I0bR0TYEsq7+UyebWj8+gB+4tvbKbwW4mCcb6taF5Ex321vPmRkYpwavIkL
hnSzwIH0ShkMbqo8PCQNwydAE2BIpN06glPmTPOihWZICv4FtslzwDnh3U1pmR21
4ZiA68HMtqRRhuurg6IJvDRCxj0RLigt+JW9r8sfx94l+gSaOf4PwaXyK7tYiBzF
BI6Q4lZ/FSFNX0Tb/w3twH0OS4rC77FLRH1sptbqN04OFFKxdmDpeLX+Xqh3f4Wr
OooulsUcT18foJ/mw2SI+KL0hxj/uQs2EAcHU4/gzkclebGfR3KUZgjvEW8/9b06
14zC6FiFlNBxsQXt2drYpXIIG9Xlyi6DkypiJsWlQRbHLq0t6h+gm8YXbSxw5R8X
uy5F9+fmIEUc1SUU9tllA2l5cbenyblkn6BJHBB/reeQQmVL7jWSbhRnNfZQre8O
4mP0LIXb6edvFVnKUH4BEYP3vi85oXgw0ky8ozEcERP+E6u70Tng5Zlr8s/et9Lu
RL8xVa6VQuTSAQfDt1emYRaPqbhz/EXAUE/3arw4deKkpPbauRMJXgT5RbPoZ1IT
dVZTHi3b7tr6rNnZeWQ3cDw/ckKfG4HnxJwtb7eWs734mvJxj0lznKw4WGAbNIa2
n97bULhz12B0Pb0XkxLz2N5VBTC+WK9LeYgemK6J4Mlx2JbJZn+iozqEc2qly283
depjfyqzupQgARuDCsbBptdvhUtahZMc5e0A+ZbILA5L2Pbqy8jsU3fUEzYVsyVa
bJHy3xPx2Hi+Ra1qcznh1v8K0Pk0z5a8ZCY9f9ao7/ifk3boL7a91jJMWHFTNeXG
why9QZM0pqCYDgSIj5kr/Xw7K1XbRLRKSwy2ZBeVQTbuHCOK9L45UKB9xbjoPAdY
tF4IvABxGPt0gl1783w4YRt5c5QPtTIbdZ+JHu4hh0YfqtjG7RUfXzen0el6QBVE
jVwlLGvu5Y4qFz0nvo+2AaVgQppBUe50l41KkBxeGiuJBGVqDhWu1M2bE4jNSNVg
w/vlSPfLXPf5ZYfomHI7E3MnciFSQY6VMXYewfb3wbyV/MfbKWLX+DiENhknCTJT
Gout3n7kuha67UHkrmT+t5SRDfrNFUcEOQTr05qXd4FJbgwwXjGrGuzPC8Wh8Mxg
XTkJ8cA5EkghROwU9UeeYcPsVX4RF4+2/5rWX5fgAPOCZKunrQJBSbWUsGDzCRdE
xr2Sl73EgMNEB4+/gBSlE7Rk/u/aHXawzSZ76YJmNfG18NzfjchfAcvG04LKtlyw
OwSzU/y1DtnmlxMik1g/173olkEnyXt4fRhME/+j4g58rrQjtCrRqADoPeWIOonW
CGNHnXt2vgsH8aKsgZqjRMHJIXPR4THwWrSEE+8BrjtXcjen4gpERjctJBN0Hv7R
AuUCZWyJ5ih5Bxe4HAOdcNz5fFJ9VYw/4kOuqseHj5zr9Yd2Bece2Xlib43H1W2q
LhjQcqvGbw0t2m0hkHjY22Qdx3vZGXNsUe5eeRCKH56P87wlM5WsIcs1VIzVbv40
kI0d7JvIRgzkISItHJem+SUnFZDibGw782A3LKUwklQA7Nf6LVgp97AfS+SxIvdn
CS6lw6XkJbuU9vGXoMR/9KaAXtyNd+y0ED2TwVD8yPzQ/omq/X332tjSGQV56b3M
LwMn9jjnGxix3IrY5bpwcIx67QddfaMWVDxTMNd0A5YdCvCTglw0FtmCf4W0iZvM
KSlR07DN2TwFueooc6Nn0KRTCnYXxx4s8y+aYVme9ckyS+PahyCfhgxnB8n0UT2j
fJwsXVw/o/YE6FupaToviiOlDnzB0fiX5LD7Bd28YicgrTfPJ8QwTHtbLHjc3Xgg
nq5qSKB6p8EZj7xexUd7z2nr5LuPK4RgwOd8G2FojkBHxKAAxVP+5Y2sAReoFO/T
fA13DiwK7K0BTqqYV9t4xEn/jHiO+K4YqgAv0UMIMsMDg8TbWAmmRymOhnG44Ydt
bj7bqB5fEFZ9ePqRxkS4CiQ//bx0Hvo3Ylfew5p0AHh9cIaw9ZNZDiOPvkhTaayo
30jCnzmXh44LT5w7iNEKCCD39Z2bbeNZgeqiiaepl/sWmuY03BLyI7eN96ZifcJM
iknEjCu1eyndaVUNyHHV0Ootr0x26R/4ofNRr5qRGSS3LpEwlMtVJE5pjnJuYRVF
m7NklohA0aOtSgBu0ohzsRiKKP7eMtBYIRx6IcF9qFrv0mkkfry9K8FwnQc6/oOo
JFKTXxSt9wrZDDZ78IIyB/2S16cUH18xfD5YJxFHaOB6vUc5a/4zrbzisEvKv1Fo
PxAa6LU4N5uiaJU3u4LHI3G9sm4Wdx85LOuca5yfYoP3f7MujiEQCB+iqmG+Gg5o
Em7kB//g5sbzaSMGlWaVcjtTmIoqdLYph3gu7U52cklAfwhAtLIWiqaBFIkaDk+P
ITEsG5Qpw4fPZPBGaPoGr0k7GEg02jyDDXin8WYIPWOsQq6s/zW8ZosgL0iJ6mho
cq6WBWktxLspWuGdmsrs/rMF8F45gcJ7Ps2QxM2yWyEX0c1t8R9kuF6G2jAYbExA
SdjteGPHyiakgqFCZfGlK5H4v1DhZKhuKpzdR61u2U409tvo73HJTX2yD8j/5nIU
dIkkgTk2WsrVAvrWCOzp6DmDG4JIEm/+5HVJLPzeb5wFe1nNH9sIHDKe6UbOX/qe
idxxejgeuc3tFNwHV/gceO+TFHIFTjie68MCXg/lC3GOxeETjNwjozvuDgUa09VN
QmEOpV44bphNOfFJYLBsXATDpMB4ICPNSQj0pX256aiTwYQlvlo3ffKAXmyy3Uz8
Vs8rQCW+3UP3NIJad51Ynezhc4WTrrcx0u7uW4xO3drhvVC7PSvjePeHMP0WKhst
hUCS9UabIWhR5AOPLym6b1ljRvNszIgt30xdYYOOWFwO1WMFd8pKiuygc80E9rl+
DyJrBaFNKQbXPnPvrOvoeGXS+BEcMtiYMT8Qbnc04fIOHPLcaepbgesAVX5nKkqu
AtAGn1jL4RnQuGkGsFCn0kc2RbminTSAD492T9Jjas99zH9SgrAh2r27C7KxY9Ao
C0iGvbIsrJAka2Gdu9T8E8s9FkKdRISx6wpubfTeg06CjQO2+lSUfOGITHLbGUs2
pCugYrwh+kWt3XC609pB289hlnhsH/8kJOCgktDI3f0M7W/WGX2G+mF1EGDg00jp
17yRAIA7hMypa3Cbmsn6Z05KteUSLN/0Fyz/xg7WCAtakdI/ZpuP1q2ja6tWFqgV
sYmBd36wzQdGVB3ohaq/eMQGpg4smBFOdB1LKhAibBTlDnh6WjB1b82kDjam4QKA
8p556/ScbpLqrNGNmR64ULG8wAlGuV2lipz14OPxiPks6HWDJ9Ff8YkTRoS5UbwL
Ii254rLGN9RmEM3+2RgevI/a18ziF2I9XvxsXZT0sQ8BGoWuxlyRjQ/PdIZB58pv
MNhaQFMOsqhns5+8DvAgRgtTvujxyvbKLSfHaIw8q1upxwkRo/GCoYX+1THo6C2T
Y0Tz24w7r1OAdzkSlEdLeJ65sK+n2cjGiFIVXvrFw4Uh7YpCr0hQagWDG6Q6rA1h
uVtuLlsvFluhjcBrP3zYAbyGXSGOMAFm0UWHSlBZ519BudpyK1h4WfNZW1D9LNWb
iJdWEJ6XlnHMujOf2XsIU9xX0tJuZkOSO1KyS+g2c9tlWeO/GlGiJiTInz0UqDJB
4T2FrBIIqtgvfthB2jfsBH+4KD7qGtMFh6sry2Gb3Y9mdj18XU88gZjTP0IlxMtk
qD33xRRYUNQ36nJHMIihQUqQRgqrMxGNgguCrSoMntNdxemM9sJwcJT7yaEa/+Zw
y1k4p4WpDfrpA/d8H6EBS6eSmIo6CnkwW29mhdYr9UR5KWSM024TDZWS3ssfk0Wv
GZjCKfTFLhJnIyiFo0KyNQr8hlwW2u63oOOBEiwJowo6BWLHMZqyIn9LjNLRokRK
UX26tvhf1uaEDTcva2RSHNeQJ8Ba6iOFQCd7x7MKZNmK7MCIncklePOzLHaFZVb6
6e2atl62BJygXd0ODQMgikCgomVPqDJDVyihCqeb+SjY8AhdL6AYjbaog0zLo4wD
p3u2tqgUOCwHho2rYpgk0IpkhApe/hbYURZCK8a0oij1LVk41IjQDLLbgR+LFvz0
MBJkW4DLKlcMw05SNTknjm6cGW1YxVWKn8m6ls0nNuu7fo22NqrIlPZyqSj1lSdO
SWExeYSd4CI+jfn+WRcgyt5bZyakZwV2T9t/vmUjVaqM93O+iisI2nC4G/mcDrKN
AgFc1K/Ys+AXBGLD64QCn1DMbBIb9IhJ/WEdmblDYVaUVb+wfBVmGtENzX2MTbkS
TDYgXbKJx/mFnMwElQqIPVkknczIyV2Rc2LbBqAQlAgbsSziohp0s+r6CcPJUw3I
pUEeAaxeY3EKmOl1QlwoDtqvZaXy7Zui7fAUoAl4z8q+slWhmN4y7G8G6eFlAsWL
gKiZYjWZWtOjSj81KBLvdUfn45qlxinnDdJuoCEo3mNNLd7Xnl1uRWfR0LeInbKq
QStqtfcQFpxb0hwP9dh7RwwsZcm9NJm7v35iyJgpTj4eOXgBVS3ciFM18Qg89G6V
sPKPoLTUyPFeA48QhnDDEQtZd1mIzcH/DVKmDjPVhDRXy5Mu/wbIm9jSJxpIwBL8
rHSDoP0z/IIiHILEO2yJm1gtvO0NQl6HWt3Ttf9D9cvpO9yd7qqApaCNnx+Dq5cd
Rgca9Y9ulwIa82isXxDVXvLFBFD9Qu32h4rsNuDMIY66xMibZF1I8Iik9PA5GfVe
Zlk4RInqBKmXSik+Sf9/jQFU4O7zCQCKeV2c6GTKkPlif/m5nXzVdnp0AojOEh6y
4AHpOiQmS2TfWmcE1aKdXlayBvucxe1502jOuiIRWzAtP225pJOTtSCEJU5IpTpn
jNR/Ih4hWU7FyOZpnIPI5raAxnRF5idr1hf6Xirtu8l8SwGsagrnVk+7kAdnveGb
Hgx51bv2ygjUQxHoSZdridtAHNZk49+lGQd13scoUzT1c0JUVAdYSxJhTW6+RdqX
aP8HPPEhnLuM5A/YaZCOOk0YQJoU0qPW71I3OKwCgXRuBaceegkHLiTnxz/ACfOU
TXIEQJUDS1YzFUr0eMhaz0MW6OHuRQdUZ+QszfvAgQ1/vWFqt1M44UcyRqPw5TtA
U+SWGdt19+kAKHzrUvhvDz+mk7BOt6fyrD+BLUQiwQcPXX5Zd/G0BEGXFeU6hSSW
muw+Ktv9+zGlR1CozB5LKDvcnhJta07aEnD8QzzjGj4GlvAnihugQozjac1qSGab
zCQdTi0g1bgpMpekMk3/XgFCpflyLiy0t36iStilsOUxd3BUMoxtG3r+FjSqtdmw
wdGKTCD/6ZDnWLGrJ+ENYUYd/OLgO2/R2S8/adnFcbF/321kNOQujZMub8HKu9Sa
GQBKjRloN0grJ25kQ/ou7pNTQwt3ua0fHmx4IxmJVtcHTDfm1Wz985iP4goY6iFc
6jP5qAwzluwnGzX6I+iV7Cm36IDDsj7LIOrimQF0ft6pKO7lRiOVM6OZbWxeKr5s
EPS2ETcAYzQmMxAUiPueTwZsShWxNETDrAKi38/ORYLd0HVh85vDlRVfOYf/I8ES
G+04zUMg2amdd4e+K/44r2JSAu9jDhAOcJGs+vsoRnmqM+PsqcMz4l3Fo/ZQ/G8U
o3mS3feNJsbNdYDjlzVFkz91yuq0u+81TcBERK0TCw4e041xnbBZBzhhbCRNQdsn
U9Jhwtqbmz/dXwR3dV9Enu9tzsBXMsFH/pCLdIPKocln6NlkVFNdax36S5GkWS5X
ogflsX1R+cm84WcsIDAXO/C4ZPS7w8FTIIdu5Mx03I2wlDoPnmt4zA3atiLdD9AS
B5e9rppswOQ3IP1vacI+Ifg3z1EN182l9Fczgx0K5IJdouaJMTQ+FVcCUcRo/Dcb
cQL69UN+7ltnRegl0ZMbxlIHj2P2ZD/CEWUu31EXIRgO0GGp2Rymh6rETnJG+SDL
yXKHV2p+HBawwpS7S/8+8gsz7seH/dm7/wli7lUgMWarlzdOUajEsCXfqwHpgYJi
C+JtIRLlUbUHoeVE3oNQ6I6oxZto04twh42fm0lEdQoTopudPGCMlzcdjtClqZFw
wzAgytbhhV6n3fX9QRJ5WEFguFG4qQsa+Eykrgls18Ev17Yhqzd+HjK825WdEFyE
osKEEcoxUawSAuVsMNttH7HYeyEzwIdXKeI4bYvxBDNqYfdG03EE1KdaEgHiM76C
5zrBlVFVXKHzzt/UiDeD8Wl+PKbeePDMnTqpMEMQA0++hDavsOoiK349mA8zY/sy
4LDsBl7OLuAEQ7CoZs9BlD240QcnQbydohdEkfFWaXhwIWfGPBdtLVdd+HgvCc1x
Sdl6xlz1OC3+6eFwROQ5lY95oSRAkgtD98hATFOqzOJkIfSz2PMiZOjYHnUjtHQK
yAG1WMWgjZjIiDhRuXuL4yeSG4cP8ExIzLO82HEQXo4ogJdIAt71d0FI1sggexmJ
A7xYroc0wSOyRa81r4imzGUg3/xs7cTGJyrzscU71hErXOGnFGMR/70rcj0YaRN/
4bGIl6mTqXyxWSpZKDijkBMx5ve+sff4NBuY2XSXlb1RaNljyFA/xeUXtRZjdc+6
0qK20uSLTSeSPVXUA4tzc0PS9i0YRFtMLUxJ/4QuO68V1XhyE8gWtg2gF+RpIUEv
AlQTJ/ub2xftkZEmvAVahqV7HEeZE4SS1BVAHzTP7+Ol+xQgK2q3QCPOE2Wp9X9i
YvubaMNlvuYnh4qFrPc29rYPFmqQrGo1WXRYDdyq7SOSP4ky+OTaPpGti6rl/LRU
iL3pFDCHTllgrtrDizccU9gg3xlk0tltZHPPkYPofNSWTcQDsL0YGoOHrc/uW7uW
owcGwaiy9EkrD4HQhPnIMLp6Y01dhAon7OQXPqPf7u2pBMqI2LO8qUJ0XjNt+baH
vhFdG+fV5q0JVdOTubJSr482921wAVdV9szYmuC/3twjmd+8JO3tsaHBKQYEgpns
BFmHTjuvXPteXggJ8L1nzyHsE7vtGMP2BNxDELEeyIGATm5VadM/cOhJ80Tmzh+T
Pzh4Skhb7gJ6cOPfIv+/JsRdtwT/6hdLh2NHxClhKxsJVY6IXiTD2rJY6nl8fr4/
KDYntB9R/l2V3fDNCvIya/7E9HCu3786/C+H9RlokVOYg27EbSvtIfxhfzfhYZBA
87D5h+QOhVXcycU3HDz/24Hm4wzIMbVAFsiyoKZnZpGl3UI4CPQ5yaqJBTGkA1NS
1Ts8dZhFkGrhVt3CtQ9ekzefFZzHH3m7tle0iL8K9MyxtTWPIm0dB8+FifcsW18T
+CdVwUNPmkakDvNJUnruICvmajc3ctIMxcuJrfJQO/onbCsyO64Ucqumz5eVKknX
NnnJj4ktq/FfcC2n6o9vfcBCgTLY4hSUuDbCyTgzRjdjHoYma8XYsUOfr1d0LhM3
6wDl09Blkg8VwYxjsOMLiZ47wY+KhbzGo5ec6QjJfYzjTXazHXTIW+FPcYSoUvxx
xVtvszEtq6Ev82JOrP7UAa0XP6uGDaI1ZP9mYv6cJ9879fvCZY8UE/Z7ayBg/Efr
NilDtboxCwLA0U+NYLRPsMuadmLIbh/EM/ffqyAg6/Mt62BpaCkRKvnyf2omwmxN
SKLEPj2m5o65OT1y2o/eQgjsAXHDpVzbwkBfLTwBFaTmG5KcZPjNFXioq2FhVln6
4CqUIsl8blTIsggKzasQr0UBh4pmlisKVsEBBfh6IYShNCgUb4m1I86BsnRSHakZ
wExtwNLtHsaQaZj+Xd2+aD7/Q3mBGp4stQZmSy9GJ9ukvU2puJIaJmNsgEexVsT5
DACwm3EOHsCkU6gXL98ftUcgqAoHct6QGDO7ATQnozzUdEv7KL0l1PQyQySia03O
3UrLDZ8kBH3hB5IF7U2dKb3mNRRPe4bksABbu6r3RRdrqXknYPe0Yq2hzbl3qo0U
rd+1JZ0PAC8ZUuAHKIMBDSqXRwjcuEhxj+UwPq9T2cBrWmxnZYQXtgLVJYSi/Jra
RmuhAJFkZKyPy+aSkCCpQ45kf25u1cqu7rIcXeIAOCeslNHKP7D0z4GW2Kgt4a4O
a9LK/thTHEtQbVGdr0v3h06XM1z9FgG4V7vnhdKcK5CJXEwlIXfhKU5XwvNGl1FZ
OUyRYZ1np2OjsnJLQI+w2EHoP0xDWFSDW8Z2bLU6vXX/b2Jqof22XE0KSD6Dj25k
DtHSVduDuGEtPmbtTo4PHDobDKDpEB2aOv2JPA9FZKjzzzSiHb5vrZqr4X0++xCI
2+I/pIpQl4XgsRLkPJF/4v0wPPrP5P4TwT9ErsM3jmoAKk3cNlZiror5dLs/Kkdc
2EqUlvR0f1UIHAe4JKfJrI8gOMM7+tNm1fdd246i+q634EZqqb5N6kwGIb0Hcp9H
/3bnM7QQFqapqnJnWZ4Kex4QfyzKQqz39BwmOhXfELpl/yefo0Qs+VSmVJZFZm3F
3l1a/BowwdOPaMR967w1SfGdKHpnGEKD5DZk1S0tiKf13mHI9IePAbrVgsS7pAsw
6lg8rBIupXmKzUAGVDw+1WFcH5LXYgyxSSbCRD7UD85y5JErEtV8oJsEooz1Tk2O
DErMM0mJgA79Y2q51XE4BV67rhY1ZF535Bc8Dv8SC+z15Zj9Hxpljh+C4iLMv8M2
9esDcdTCAhkwD3vba6Ua3FL1NaIMQGh5eTIrjXVK1cFtuZOtijy0JJLA4Ri60Roe
C4i6SscRqifIjjBKbjSWn72486r6yTYFmEXqtAdL4PwbG7tM0RXyusQlJEZPJT3G
V5XmGJPyXrHTw+xZ8ZNdLK8G6195D0e1SfDkei79NvTB0XGl8HEmdBgWwYZR3hFz
ruieLlBO77lRidAZcanpt2WKazZn2zNqG1KL50PIpEXyneKX/1VMyVvOkdE0xQXW
uDdb23gHftGfuv4leAsdPWCgUUCrAA/LEJgmOHRMcJdlmOyhacWCzL45DdI4wdHB
fnJ1b662xx6ZeIjyum20uZKc6RL8wfao6nPPTqCDFVu7t0UdSbKH/mUiYAadcdbg
O/Q1L+b2+o0zifh25sZ62hAXZD/gf0Iuv/MEz3ZXEFcqC6a0DlgcJTEeLvRAoahu
j+P+HFFUXEiGEuJgWA3ydFv/5PFul1Vv98j7xdcelKSHISuhwVAHGnK3zi5MbGWV
96mKVrZMTUud2l1dtCmpudyyH8CAwxRpXBBLEaBFihar65IwCgZrshMZlLgijQ60
n8JwKcyYktwnhAsO0Qe04A4QYCa75OsUE+sm/vy6qyT3DeiAQThMmJKT9tDNNZ8v
oqPNAoXXrWLMnbnEWKgirs4AK2OW9LHmZTfBMwSsnlIxTObvmVNRZr7qi/Sn41Qn
/ZQHKJ4X8kaHYJ3WS5li8YowtOU5PCFltn/vhcQ91nCMZ+kdneC/BSudepm2xK4/
fS8N+qluzKuN3CpgSN9YIyrt6TiiRGK/0hhevLB16HlNlwy8riwAacXgyWVUXoC4
ESg6q4QW2ffyBuvc+zsGpoTavMRzzdj4cnsOQmWhUi8SeKthEJldYZU39b1Ovz1D
ZL//tVuH8OQuPWGbtsB8ZSV30CfAauSjmk/e5LqQ7BOWNwnWq5dPGo5pHHbwsSOD
guwV3w3/uGKfGIVg2vjHqo1Y4v/kAgWAgR0laHklUw3TKPs2fhm5QTVWyHfm7ryA
CHvXtj5oM+BvgPZ6S22DUvPbwb0ou7rlosiWDjGaopAC4p5x7QacHQfwccz7249b
m0iD3kBBh7v30zHpHr5MvKhkRAPKBDLR2D5N4hG8hyWbrJhYRkz42IB80bBv+Ue6
2tV2fVYxHJHCqurr4yyfb6JFiA/7zVPSZJ0j62wObO2rXneKuyPCamCA2/kNff9D
g4zLqrFJoF9gs+vsYd1jw4TBPO/Wl1Oc1qt5wcW+DR+f0Aju+mWD/NsfLCiNiO4S
MzZcZ1BVIvDLKKLWedM5hxlp0RWTUt51foQauursn3ccpMybrh+wLUQrJ0khWH92
e25IxaDnTjnsIM7L9gHd5KLO9ah9kOR+4kOjOuqWAH1xibx5L32nZoqZ9FyASE7k
J1SyjrQzsMgfukcjFmKvY2d/KYosk5rq+WggD6zCgB2u/ItVrQhP5IqxJSezpYbZ
yidApndEciXehuKY1ZC7bp/K6d26fqBJ/3IcSjsLOTB0w8gOGuoPSL8wjbGbjjKU
o+SqynF7NQwP6h58B0tp/l9aT0pdOT5+7+Hz+wdy09krJ4Eqzv22QniANhgdjlcD
CfBKE2qvEyqXscsrAh1s2P/r9wuIiLnDLxUZ2XRzv/lPSVXI0n7zDsxLqEj7mISp
4bBmjy29Y1fSqYmFC3lKRemajheg/i77I2YSX5/MQ1K778NPQwS/i5MY3dSUg36Z
BwldPQYDieTCXVePl0UJhA8wR7s7c/L25g+J8p8z/g3ds2s2Kyh/n03U3VrN23YL
/MRGrA34PhbpQfi/8ZvyOwSDNA/ydYqurtujI7SW05Y9Xmfm5CU7QdveT8r+wVhn
A20F8P2pw2HQNPaKQ6QD4BPR+DuWvzne9wl38eZzFoGxy3sgAYlxBIxjrSi6vVCo
NPuaOnvGgBh333QB1OHgSalozQ+rGqZavLlKrniGCtYirhJ94Ydqk2jau7KxtvKN
niDdXprtA4SjDp94cGn5v0p/dQcdMJ4ErfvwCXWqN3EhNL9KT4ay5AYrklH17EHp
hLOR6zxquJTrGtogVdjeSUohA6OdQ1e5cBqxj4S/IJ5n83I6apwNzu1oy64obT4E
Mkoqpe/Qcub6e6pi+ozKnWZRlUAQZMP4ctmuhP8A9lfvMUqNAONre71r+/FC7haa
FRQflOG1R7uyFLeObE/+3lNCZnXnVeSOzByre15VEeoFrX72zb8FwLmbjJzL9RHR
++qyZj31MwE/SWV193MxUsrb6v9fMGsExOALyM3IAQIObMOf8x9sLfp0kG83a16o
S0+96yjqHP/mtZe5t/1uSqj7zQCfC6LfpdXcgONmd2HPcprwLgZp/9ufCiTQJ3uG
x3vL5QauJOzQiu1M+d3OdR3llUgSA2jijv0tqiO2zNbmpahZd41ohjeW/s5LfaM7
ZLUdOg1XXuXiPt24RVWnSuWapsFdm27Ux7RVmvQDT15zUaK80kq8Bqffp7HrFygP
ILkcabufVVNb+eKTm13Lsp4pzVNDPDRFiGWSj+BmFqg6PEvegGpl5xLgLXWEJUFU
SzCCYGc9UY+7mAcWdefRkLzMdqXdpPCQ+Ks5iRyY1/6iT0k9fkXR/U6RtUeXxJp0
Hkxugdt/xtioJ3qncS+hGkhgGXfj6Z5mTBgSvB2NXBOiLuew8uSwTXLr2CJb2PFr
L2EFzO4rGP/HkIeGAh1V++aau+O46CeIBbTT7JuUJutLxMBYeIYHOscvwfoi12os
fNt1eJLRkZvvUoqQRkxBeSoM9mcs8DP6F48c61lEVvFbPhIN9GOjDg7sB9UUzb1H
EqVGwa8XNrN+mg9XYo2PgP2yfb0nAXoC+H5VMte5t3gIAWFqYFojQI0VhF6+6EOb
fiI6le5bQnZ5kV6HTpDOU8jvajhdTs4Ch4tOMCoeuuS/y3DDlIsN/Ifi6yTreCt3
qRu5WLhOVnUy9RYxfDfw8cgy5pPampj9K9vW5XDn0oUPDP4W2H/5nPYkG4ddC+I/
b8cunJN3Bag6ZvLCFaFLNhCoBcJUPxAJS/A+BdrAPtqoTEOFaaMZQzrFyXAoB+Xb
nwYWkjYXRIGevSOgrJgusFJ8e+fqOYBPjmr8GjS8qi1KNz7D6dkUS48ajcNhUvsf
WYWUYsPg9/C0CfYb7so4h0RmOuCD30C5/7M5olzH8zc8BvtMY5hq1vRTDFfgaTdW
u5hG0lBNQCSzi8JGndbyJ7zW50L1oZIZZKxKZ+JbtuEQowQCPQW/Nj6/OQboXUk3
V2McRidMJ6SGUluIcgyHFlWFQIRgNd1TC+XFs0jidCTofuYKy52x86OVey55zXB4
QZnf2yJP89oto6xDNj8sAniFsv88kP8I83B/qNaSBBGoMTYTBhYT98ZeCT/anjOa
WwXL8TPMFwlI5udn8a8Ujuc/kCIi1B9Wu7cGOWhv5mWO4oquPgXTlylDBkk95liI
jvbTVYAz0USToe6nd3bqOHIiH3K+4YIaVhyEkYhTShM2lFofGB1QkdqO5CshxRnk
QeW5yL5yUgvnxgx/CIVQmDQkR/AvywUwD2OtzYs/fnhOUCLCdGM5DvjP6+hjcSPN
zD7zNU2wM9GPcUcpxVjeaoHb7xCClu9/fpWTi1vyLpoRMtTNo6opsKXfBxHg4X09
Ix02IuP4eqTs2GhPE/dM6odexlKvDvZCXLN25jB7srkx5/sj9V9L54rpaQYBpeJL
+LbP0Phfb1eKxFYFZRLSBpwuzr9Pxq+WvV/bAYFnrvI99vP/fgnoNefJ6sU068LR
z9mq6Gd7f9eOOod1vFNRsE5haGo/VU6AKES/C14XyyxfomgWfK8RUHattwI/Uxrp
Y0kj90vBfWtK/N2VitiWnK2MVygIY0I6aC9DpsIz8WHAUHhqK/nbDFAiM/ahNGIY
DkWXL57/kp94t3zStLDqjUo++PrCRgdMW/f1zKVFvq7kmhDetbcd/9wa+iHC6sMj
gwtiuJ8fu3gmdSv5rnhIMUgVDQxeJNKNX2d6JtNgfj+31pzaIyCdnF5k28fEfvJA
GZJ3C2nR7x087uhZeXE5HHSHPr6+HaQ4cMJwAlD50IPvkEbzonlHSC/4GANqnZFz
t/Eo4/0cxItusIp9NDjO2Z6XLTKyx6UM8pn/+8Sw9RTY0ssHHBSvY2TdDrNefz7w
yhghzVz1AfE+qF2lyqvHxdUFIg3o17nfTtU+iIfQhRPBREjqMPg2DbBmwRDZBhAn
Sahw2SpIF+DhITcTuYydso4BGyKoLMT/EqQ1EzxvF5xjGkIgQaiRTsyI1rSXX1rN
ax3AYfM0BNY96pycZAuW1pvmc1JW49C5jX0VL+zqRyB087SA8sIJ7l/8c0A3h100
Kh1soUYRB5NsJXpyp7nBEPlbqvkKyBaBDhOyWJKFRi3QWxpwxI14sWGr+12Se2eE
XItRSvWcWIrqBK9kuvejI9K7EvseK1SJiqbTeNY1Yl+WqteOiXWWJH+A0DWUaoiy
qZPYdc7e9AqLsVFwdyvv61hHaweIEoizq4G/lDsWrbbQfileu9zbiioh1S7GKNfg
O6vafvNoW0nUB6psrBM4WApEJpYxz39S7UbAc6T+n8A+e9mEVHS4v93nIZvqS4Hv
VlJrp33KujmiheuGjprkNhZcWR+zcxKzj6ozxoN+m/53GCyJjxP5jzj+RQWFuBo2
DPjcS0hAWaicWOJnaqvAbCnQVeQOA/M8m618rz4Oh3Z06SnYxZfTn5Hpx3G0WQWL
Na89zDAmP2+BYwSFIEEpzA0cNpFUpDDDTjSdzNy55O4mqsuIyzXiqdtcUsGzhmgU
yNzAM4rcdbXdBX4kdBa7BaSvliEovnBXYVWzpdiOplt6tuc/dcLTswBYhFiwNgh1
kzGXv8VxicWeilQpmHTBltbdsztD1SJuTW4SK3ItLsPsQEcuE948T8J/NLkPfvW0
lxw0LbltNObIwbjZYFm81YIPWA+rRHkrm6GiK6rml1/WzmFSPWi4iTEe+exNkK+L
PfPtei2YjYtguX1j40UvZ5Io+qygpS0ikTWvo9FANwTLbI90Y9mYdyDu0Y49BeTY
Sz3BYggA51HtFuf5zR8xAGGlFzbVpSyT8LrCyvdX/9qCJckEwjst+agrmFl0LyTx
Y3ZJtPyKVyMF3w+fTDEGLfg7h4Qi4vBJgR1zVA64JmUUb8mRaTEBBgJxoZvbpi/Z
5y3sx9Uwwl93Y0GeXMGs3T18GiYvoQqnNAIyUQDBoCEeOVXc/neQhd2oSMDEiheM
mJI7/n4a0aK4cAcyOp0Bn8+CL5/YpC9TqHvrJNFuuMWWY8nBJhR3ekHGzLJWVrF8
NCY1riCFO4+hT1WTAitPwgRt77uv9VbcOcF8dThKu1WBffgHb9KRKxFVN6WJwEbY
/URZRZNBUAIVRRuPEt5hlOf1UuVWzRXzs6W1pvmuIuNIrIRf49uFrQ1JVCTRHPLI
XJ1iW2UXfT6746myk1or/C+SqJPYP034zHusbYwyRZNk0FUhpWVTz9eKjyKI1rKB
DJexO/dWQiwHhEfL9wFKDcHSV0y4FVgeQzVrfulN0+EqZD8cuQt06PlKSHw6l2oO
AtLsWqzb8CUAw9onsQIqLp7dq5vEtvilyOa5WoitD6MHwzNF2HH2cOwYVM+S5f7C
CIlUu9FfW4FQCLg3Azz4+iIXJx5CnQXRd2grDYPdc1wB7g3UYMCsnj/20oNgHz9C
IZMaBbsFvTTxXCa0+i2XwWyR4Lu2+P/xpcn+eitaGbo7p3+C5OvFoaku6q+0TX90
tb0YORSN6ASMpJLlV484qRDe3tULVGj0f0Dg8j+1Bu+wVUiKDGV74W7dn40YFDIs
wX5AA94zelC0V+j1ZqS+cvVQ17ol/3azuh2tRHl7XLCZWD8xha59FI6pkU4inrK4
7dNVJ2IFIXP86UHL/c2ujGlKN4iriX9WxS+v72Wwwcv7paIhy8UvJlxJQVP5tIUq
et/GlpGdo91GPQLo8bHr3gO3c3WF0rxm1UPZLRjDqmYS6nVZTxerAw5O70MTF2GQ
QPvlnEZMzorx2mx86GPBbDFqR7dQknNT6RYCLD/wTztqqX7pNKY8Jb2QxpWflX8k
OYU2j7cysBmUYJ0m1ZNyGQi5IEaDutDW55abzW/lsUVAQT6MoTOt8tBbaS7Yt1jN
VEfiLRFju3jMMgvXDTR537cQb4tQpIsDFFHuKZbo2A6IUE2qDjrlkGMRAoGgnEQu
9Q0WuqhqHPQOIcmzm82ruPYdH5iiLzbnDTX9ZxQau75DKklhbimed9p/+n2yDc5C
MF7Mo6RpYEjTOMu5cAyywggKQKFujqUHV67c+F/7ei+MKz2sgpXJlSu5BkfNfFFI
tTU3Hd2xJvhPr4mgS/HYdu64mnG98Y7FKQyu+06WGGuBw3N/tDOOoESNP4+4XaVx
+DcmA+MEGbD9R5kqxpLg0PXN6x1T+lTgv7eEHYphwArSIVeCPLVIcmlxsXwPyMzz
dpYKJRl6yZdWu4iJYAquG2LSTaQeHAZVn/vTUjDZUyO4hZVJOjxaFkgM6jG2OQFM
ZVGbKGlnGYB6CcYufg/wRGPJdEnjXEsKVwA7CCxEfjrT5GePYUehhylZes/COeWX
Z8sVPGdoafgaoOnbzAQZg5+z6WRr1ZZsSh98nYspxMScVOwOQa2+MTKeeX8wT0u4
YOTcnuyFjqBIXbEO2BFHHxmW28+/bI206koc4kBTjybBZTDwUufiZ22VvzWZgvgy
LCsCScueL6mpizgcdEB66ECAxDr3qtq/U4XTmCzIuTt1adaRjbgLPt9br98uPNoa
vt+kLYdwrqTqS19mdE4s9Aa3drxkpi/kf1lcohkKqf619oI5pn6NiBUZ/3P/iNGu
DdYglo9K2K8/VkDAEI1D8NAuBfHexbJ8xsc7cbumkbIoW83Gr1cqXyECGOIAH/7H
BZnSLt5kOfvYd7MushgrDvEwW14WlcXdsz3a5JMtQSLPAf7BQEvQeFGXH6cuFc2y
ZALSVYr5et+lpi4Hybehk9HZntbB/mmY/4NuFaBZYBOLfXXOmRlX3p+QmV5/KxjG
Qung8BGKRLX88EBb1qLJRBwgfsZ1DV1WP0b2aiKlBSKBq45P6w16qhyqbKzlGepE
W2cKIdX2or6W6bcLfbPV9DhAgKCJBFOxefim1kSlbSoIVW14W/Ob3twoUIh+5200
56u8P3Ao2rybK3cvG+5rFI2eBhvDnzFbOEBmoxEgj/kxeeApL3gQk7cZUvxYOzOD
0Wi+5fuAffQN9jGOhk/Xc5dBtTvnoMxOV+8onQYIXO6aJ1BuSFM/e0NbG5bmwKp5
RCcI1VQBVnQAQ5+DlDjb+/3mofWpnIGsgoIdldvtyZjx8ttXOTWxlZ9n/GZxxxb5
cshkkQxPM/m95sAXLDPcK9rGYU4higgEMUCaOVMGkPGOTGvcCUA8BP8xTBICICP6
f+j+PwO7hbjNDtgPEhITByqkiOQ9t4UiLU6+ClUaaKXxAANM7bBe75CUijzUveDR
XFh9LqDV6Xhh50KVVaoaddFVOvD7vyoZX+W7GioFyLbG0JfmLyHB4XnFDNCKoOT/
rlQs0ZGB1/sxIKxB5qJ0AIUcTtNEMT6UKlFsJGKDag/kMFSLty+nFLuGdD7r7aW7
VBrS8CzEJlJP3Y1W8jnwRNbvjpkCaUw3N6jm40i3HrlLs9ibVtf1m9BZpmU4ulbT
rkjcKam3LYWXCqc652u3W7kWABKf6GBsT4vSTqhC83OU/TF+sMU6NqE9AVp/Q0M3
YyX4SwUtuD5pCSK3CGhO/9/hFXDhU3pm/0LB2kX/gS7ujJjcn9Y5xs4puyseONhn
8ZVyfaQcLMKPAzt5hPLRXrO2ns4lefEU8IIGnDnyDEw5p3CRDxVYTM3Pvum5hktV
0W6DDR9gTn56kB8NjzYYJoLMj7qJx7ixEWIbGoWHty1BEOzk6s6Na6uCDM6fDF+m
e5VFqQNdGGQFIW1GPrINXyV1uvLCrStU9z+hj1UGjOdkzpVIL0jzZUfuP2m58Hd4
ULYF2hosLyNrQ5xqzbAAQpZbreJ2crvZCFbUCOazl+UoMteWAWzOQ6hA7O1nj3Dx
2f+ZJWVNYTmdQoJ9kzezk7Ok9woNLaLJKbEa+dvr8HCExNf7QOiOWSYWiwU80o+F
r9cSWu/nmWh2hrmoVqQWt/837Lw7n+O+o+bodp8X7SEP0YrPllH6NZ5uAVJUsD9T
ph1639OtFE/fEKCNPk1z74RnEttIrMbXag4cIN+xazn7yKG7PWviF8qaC9CNu6wn
PLFz2dl6/Qg6gnj8osYBSDjyKS4kaZ0yJGuYqUmOUp68F4aD91Tlk5yYcvTXNTuO
e4QqFm77+8HtQ5C18tq9xKl0azrIJ07JRKfxeyNdfeWOdb6RUi2Ee2R1N6Cm/SqN
2/It40Lx53TmzYQMupCCifZhilIJ9E9Ip1lSGqwQnJJu5acGegvszexjAUd05Gpk
dOD1Rv1NGmRYckItj4wnGItBLTH2ASqzl1jk9nWEWma7+NtOirOIP77Xa4u+hyRL
+1kWa31GQd4iqV+MZFAed7KxDUp3A+pED5pOjSuqe/RluXFpWEpi2iM8jPahRctv
wcUUrr7KV3vXf76aawiAyDxR4ySPKwew91DETMmNv5wrLNZHhkomQBvaMPl5nImr
mi4ohNBHRzQx4I56K7Hw937b2cY73Sz6s0Qq9EKq0QeaklNa6lAJ/8rOhkqeqIsa
ftHknvL89TsfiDbeiN42pVe+OC0Cd9FkvwsTGi2CpgXQ6KIVFyPMz5+g9BX5fvNO
kBElxnXKIMrIebERJObBCtfm5uO9dR11RqKucTrmA6tMz/rAefi02l893PZkkdpX
TefPAL4rT8I8x2V1kRF43C8HV7x6USAbdBXaovHF26URB8ofIVyK1liWbL1cYyl5
MZsM+pbynFOT/Q4kyBnvRoIGTG5S1s+lvRDyobpvOZEAxziBbMUin2N9BgFtF85l
CBQemQqIMUen9cEosXkp57xC9c5vDCFgw+RthcFJ6YLsegQX08iPcAODHbrGvGJL
+V91IcCQi+qIW0yHYTjxqIJh6fDD+67R9Q19Pq2BCCb7Ruu3Y2qCQTP3LI7gAZ+B
okKkj2LSX8G7vvhcZ/NZRMmIzhvbEJJ/DsG/IOhs84wfZX5+wBlYF2pi6OUE5DDA
qQpc3r/JRc3JKO8NNJf9eWsX1JekiGJjGUbuUwLC8PFlFQtRcOyrE2anTUWBnGfa
xdbEJPs1K58fUYPqVX3MJSy+FgvtrPAGFHJsQDeLrxvwDZX+BCxUJDmB9Y9fkq0o
r71U4TCL44fnv2/BXCYdrQyJ/BifGyZrdjXxowBgo1EpI7gO0e4TJ2seTINHMByH
QfH2lgKw4dGe1tfNjnHGS4GhzLKryIC6oOootyZMMgrjiwG25o9bEYu2RzdgpVZI
uyh+22uX+EOsoIniqPbfhrNoNO9R6BFAAFY/DW5AS09pw0oxmjdx0Z5PC/sutjaJ
HTDRrzexN+wVCuhoUBDIBBcyt/xXaSj97RAUlvHthhnlzzh7hQFE5XbeKOFgDEtE
p4c/CJJ6tmYF/DI1vwzO5SE1cWmqIHFPqQqQ0d4U9Tw5fv64Zg5QDUc8D0Glv6sd
XMzSEOR+v9dOLNRhk1OclSmZ7f3eeOx9GHY6i4j2yyILixAY7YmyqAhP16rwm+w7
lKOj+volRzLeZB8WgMIUKXsG3sqgalfpIEU50ArYOCi4x8KVmpyjl0xiqb8HapC8
Knba8DqULRnWSKBvMyB+RrU0bBDjfMEewiWZ0Ws7z6JAzL5WkcLl6xwuftuHGV0U
aOGdHJuBbSIL83pHgeBBBQXcbAxiBhJgSZl6bFNVmxkn59TqtY/Z5UjW0eQuuj+g
ruOy3fqDhc31T5qyqI1U9RBxRgOlz4Eg/3Qm2oG+lWx4UBgTBkjyK16y9zTEMhB6
4DFgBHF/N5YFa3aVh7CH3n4h84dY1sbamm3zttFlTzXy+r/CWeTj65+d0lLTG1Ye
05VsRxwxknk3AmsWyBAdAr9OelDrdQzSL84heZ2eiVCsby0pHWUX3LUfNue5OWCa
lNdt47SlHXY/C3lpNjkunWRVXk1P+Pjp3EhriMhHczbA6UwRUL3mzicdkrQqXzyU
Kb7u2UOhEuCZs9e0o3Dfe/P8YjIlrrZudPXskb1o3KcF3FxkYRxDtoshUPzplLQ9
uVaI5p+IWx6g6f2i/nAh8zSUJ6AwZzn/wKxj9UsBmCCWnVlIcwqdRrAeQGIH9SAA
309vey7nY74u+vEtDvvhLYfX6sNYy8xJQUF0uNHXCPAm5K2mRmYcpUml4hnb15a3
XHxo3f2o+KNKi5XA7fvjcbcg8+rxpLMEz3gK/3XjEZ4R2mX0JwXtCqPp+WntuBsa
601ZWE7ponf1r+mA4zz4pZXlvbSIXagb5qre14Gb60KtoxuHUnFZT7W5MYz92dUJ
hpGIjzkHfKnDMLME38vnDAv9kbsVL2P+BJbILmJwG8Kk8oovnKP/mgMIpCONSW9e
gI3RXO7MhRK71EAHpqWu1dmlNT9po8x3ulRbjjB99go/nTg8yBcNVG+zGjX2Z/i6
NpVYjbFq4V4OoB1dqrs0zXwKezZ9VasVDh3uA7+yNozl0RqzkSzidaQ/kOiMRqQf
YHB8qjezPQSQU9x91L7xPPk7c1sPyLpqywNJmWuX7ortE/fS3eJ1SJp08yvqR1v9
fRKWF0fa46Cv9Xn+jtDkWc2PSiEUkXP28GGMDwsA8uy6VnvDbTno/uHrV5brzcdQ
dQB1tObOJkP4lx/govWf1Qx5KmDm8ALobcck75CHf0j+6jnsTWa2FgAo6zCpaAcd
zitV/lQQFjyZASUXKjddDzUqM1kvJrj35kChzuSORQ5AhiPJLbB111yoTiBGd1aG
qTZNR8DTVcQ/ZgZDjgkcko60qT2bLpOGuGjVSaVm2tMquI8U64C7hsoLRZoz4j2N
x6+NMRnzDvMmUPhbveI7pQ4QIv+CtM+9yyROBABj/FE+Tixj4ozzWO71m2wptNNG
YCG1+l3DifF3snyBHUyQ+V1gnOgKx4dA7jkzTr18mdUB58pbKvY1fIZysisABxLN
gx7bSmcGjxsxr6mKujlyppLaWOMbe59zM3qR82ErCePI9/xLnfz4Nmj2OEnUrfQi
+BnkcuCIEHytTd5jlVRj+CwRIfnmFaNSw7eSiZBIsHaGIbhYyrSpPJvvP92X8Vbq
+L6Zw6FM58UFJewWPQ4BwBQzaOarYlX8gHJnnzZuQIYPaGEdn2eE0USIYRYBZCvG
gjtH++s9mfH0K8TG8R0kbmBHXPJ5Dic4HOe8QlDvLvcnCVguOfS2mYL9DRqNP35t
RoYvSZiN0zAhPcENJFdCDnrKar/PeDStPZM/WIJNviZsQR92Up/qmG02Jm4kjlf5
J4kS7CB/+FRQ5XHGrwQkjuR1M3IC6tT//0nZxrydeSOXTndFBzSbU20+XjQd148q
qKUH5hBOo3k440ifbUUR7hVmz4MSnXR5KskdWFnwDcOFTMrt0ibWJFtYoMWKf4BG
1QoUgyXTTBmE4TvGz4EeuIkZJ4BMpollrtPOQtR+SmKnmHKoG4ZQKFwDgY+px3Ax
/RKnoddWAZI0w2GyPzMitQgmSmiYdtmhAVX9JFNp5jyyseO3630ij6mMH2RGmU0j
s4TTZQa47IBhd1rNRWByIvy+aRvUqRBw/DhomtQifBomBLVRu3qxdVTAjMF09+m5
UIxIzOj7ez5kldFFVLai+WtDFHY4udF9UvFuav//WwEIAb6flDAbNRRTDyB2yy1Z
+QLjpKzhwQXHROVRAhIZ0kHVM2SegP4ip1sxRGK2bRStE5RR738aepdOLtYk7Fpb
h/qTmbAgaX7Qi1gjnWREQdi9PLLGiXYbAR0OBNV0DHB+hGTAOvFhjux0ITfFfvXO
XUdCtF+4SXZngyQI7M0dkiF3uxqJwrxdDkmCGP2Xk5oCfDVAx0Aait+98msPPXWZ
hHo5YoJ1kZPk8ywJefyPKZvXcl97Pe+VxexETWWCwXWZLQFBXarmpmMpMWZn8Cqt
6R/NHpzAwuS9lCKesTb/FGqNZNbKsGWQPGEvN8JiAiU+PxG5D5LTU/LYzjpwg8A1
7gTJCsYNHAj1uayow88bxBdnuly1ANKWBQy3S9WGTKHjOVej4ahQ95Z49EIavBTF
jwuLzFmCb3HWD5aE90aZVsU+EPvNOtW4CfQFveHnHtYUxLUSb+0ZCT01Pj+yEZ8G
617k5SORkTFH6tpupCjOE2P3LQQsAh5+FDkacDZjodMpHRnbo9BkwYL6eQB74aWY
pxEjpvdK258b22ghvQqMPc85i2rwlSkuI4bgUZOKnVQMkICcEBmzf5kY5Iy9amwU
D3BHkJUa58hYiin6vw9evPW+r30dRxgaJNsyt9169ue1ffUt+j9HXkwg6fAxEV1k
BYSkoM+za3rUvPMoI3XCJnRvBCxVCEIzB+Io8NmSN1H7XuRSnpKKmg1HiGj6P40W
7OOc1FeoWwAmzCXO6ormoSChgldztCgohAHMxVzGBaS8WJbjNHrQkAcAzwyqFmLH
irTI9EalIbhaYERJOROEVHzj+9MQx0xWtJN5Ue7W/9gBAmWa3Q4dpzzl/UU4ciNc
tPBVvy5ViUY8lmbOcURgYJL6BxsvryjL2rDpEp9lT6buuTbpnn1RtMKkMKGYxgIK
1TVPKihFtvf6VSfd6+04iPzU9jfrzTB9slT3qLWFnnSCnZF9w/4gxiK0mHlOcnNR
G0mEJlBjrDpJsM4+TCesuxKdWj993jVO1/Xymz/gn8G/FTp+BW8Hm0c538A3+dpu
WGWCoIeIvstng+FpFKizW1ZgfXIttppmoogAEbZ/1+5jpLsefwuD+gQ0Sf+AvWAb
gCNid2A0bbkBZfbozec3OLI0bjSD6iXqhQn7uvaYkVfrqD7PxPIGXooDABmgt/1s
SCKZRNcNOH4jW3dVJkQY1E5JGJRcXm50HJHTZLy7LhLSD2SB5kRhizQX2AxUMNVd
jpcMPvlcvx7MZApBgxXu7QUSsF/2JYiJqm1ltkm/6ju6JXCkYtM3G36NEwrSOgnx
PEWvgEdfuR/p1ee5cZ9ZpZlVTvF9KyGFJPz/nIiVjw4fnzB7KEMld4DONkdQR1UV
h2e+v8rgFwIhfEpdWjtVPOpdrjIa+G5k8VT8zsztTtXXP/INcIinAF5gUJEyVIWy
uBajvcSGoemVNdaXKfTlLHsp3/YGZv8f+NzV4p3qt0pgcBLrWGn1KBE7TfSOKkHW
xtRJu1WsVtuCygvWM+3mPnyV7dJ//Wcl4siGQtzzyjIlIo3OIOsOAq90T6ac5abc
DX/eq8fhnnyPqx05Z+fC44e8UWLk5kA01DxDXV6XwyzVUmbnM3gmdqPewUuFkPgQ
bVpltir5i8ac8rl6eel4O6xE4ssFkyUoykMZOQJj3la+MYW//Mwk7DuwUKt0OsCB
tZp1w8bSBRSlyh99PZxqrD3uXGgmkkytidz6sBsVyccaQy9qj7PtfqEYawZqiRTU
kTtuhS9RmQSbPIEJ4QQ7H+MAdKvr3j0TtJnDbX96UEDVCqWQvCy1LXGUfKAw4DCw
/v3cF3JeqfCOxFzxZN6mYKSU02N6VoPv0h6HZg5W9OkKXpgXR//u5UVl3CzpUM8N
Je2NIQQpgYLl1/upY/b7PMW78bQ/QjmhNKoWytkhnF7lrx40P7dF88K7N8LNql1r
9MBIIL2jx8akhIIL/p6vWTkPfNBA9j7tiT2kluKdjcXK5h5g+O20qSFzfetvXWf1
b6zV7mqJnJes50HRh4NH/H2Dls0qqjExJopZ4lAUtbcii3+YSaGMNgJW4Q9lJwi6
S8aCagJ0DsTuy356eUg7SW33PjdBdGRU0w1aePP1J5aiCYErJAc8KM3iJTTzZN90
hmKF9wIU7T9cCQ15UwDFt4/2LKBmAr9R6IlHk7mNaSKAyCHGCM+2bmq0M9ifsDig
ETqlMmMjydcDn+kYB/pP4UoykzFLZDGnt2+Iq4nX6S+lSAnF1BvKo/fLijddauYI
TJgxHg/9B+1YlrABIXTXOTYV7YWlLKRJvRazFUm6caUJ7FiG/0Psi5bHm+8dlxSy
Iq93Z7IkAzH6ciBAGK38n5Asi23uRBZ1oRtB3umMlLYfcW7H5mvRmK3Om3lDTvBX
SNr9JBB2+Q9TPWYlPZpYJDJrH4tGFNC4o8nv1JEzWYi6FkJWW3WemSqB9Xwjqpp6
kNfBtre5n2u9jhbsjZgDP46k3haQl2iGoJexpCvoBAM4Y3WDzCQ+7IZ1qlNivcZR
O72n36pBVTf6KtbsK00GrRov9oF6ELyIgvTycO7sTYAdbnuT9IHBBsg9xO/sSPRZ
sRZdZs7Cd6q7eeYUhOy377ZHHgLD9UJ07E+2HaT9XXYyo6PlFK8bFtU+85RE6Mtw
K5N3/HGwq0hd+9M3JHFjSpiQuD/kf9LadpAMyG6BCigw7z6ix/7xjyodKDBg2ZAN
1PsnIiiIS0/RU+ngVkayoraamxQDhQhWiovikZp0spHmUMBkLLBdt0/d6rNWddNt
ZcfSbKkOLuKCjBc1xwVvFmBgij604u1zVLijFIjDoCSyqdw/DHhB3AyKzYIZPSB6
jN/EbvfTvCF6VcLYjYp1r+iaLF/Bz15J3cgAf8HbG7V2SkO8hJHRKC6ASF8T+Td9
qTSorR2KWSyhfYAh5/jbS55VJ4mF4EYOVYvdIDtAwfLqcPCeCv5K+ZJheCICPDKm
nFi4VFF+VqxmHKfpwUghqZLthvsfxUV0Bxc3ZhhnJZrXpxR4XlVJ21nSchnxBlxw
odSsRzsck0auftiiN3SAm2AE0kI6NeugtplLbABUBSWS+BM6SRKLSfBCpFKxEct8
MfVPLhuUJgkdzKrVoEYNPJDjCNXXLLQgfQt1LoMa6kVkk5M/M/bU161IXE29BZFq
OOvqwRcqrASkQCzDHvV2bGLbVNpJMdkffBvNWyq2jOP0DiXnZGl7+TIDaXN9zgG3
zD4P7WlOwlAugLy3B7PKMsy5oYxoUahnAErrNHycLB7rldSgezA17/97kGX0GTT8
kz6bi/mzMSj4J2C8I2ufeAHKMMK72vd5wN4tEBDaJ0bLxXKx38AzPo+C5XYJLNWb
wK+Hs8LLKzr3JXTmLRBGLnZQBVvvCd+1bk4nuE4JIyXZh0I10ioWyjlALChbwg44
uHRDhhAhV0jdwI9nUaAYgQijMkmwR2dqBK2jQWf9dAb9MPh3/UxtYd6dV/YQ/rDL
ZUr7o0cBcup6NgAEWe0VfvS4+MYAdFzOLI555inrxXEHUZI2kse5pqatXRdRVet+
4s1d5enV1EguSsZgCPTVpg9rjG6aDuK1DIEiB2KWJlHO3cv6zHfPf4sh7TVYgnFF
OLYvUDlYeiOj6iJMBGTE9vwRXDFhuynytK9GQeVljUNha2wXVUdZWAJtCNMgKnNk
SVwzEVFXFDU2PHm3az5pn1MMOO3unZVB1CxG+3dp7RXcw4YtWnHCfBbh7ePe+Am2
aHzHeCQk3mKxVvAElZYCUlbJLjN20SI7KTW5nmGGyMoq3bspnsdKCe9Vp5YRVTWy
6uLGewzSButmPaZ9ZYdXqw5kpYDFAzl+MiLo9CGk0WWOapFscC52Mj5npIg2SzBQ
VwJdkZNoD/SVESY6QondExRpq6FbNo4TMgE2tIVV4o+y6J1glUhVTfVa/nNzZCdB
ZTCi+WCufuUJtvMxO4akpr10tXqj0gahG+LNAFYVeAcnpNiZJVDdWRvsqQTW6yFJ
OyXK75ygcq5tJWV809oH1mUhz+ZXaGctFkJ1OJuPa0EpY8xEV1QHuiqMtZHVmpkl
c7Dki37/yjueLe9M9vS+ZHYbn08zx/Rm7C45FUdSDFzuGxJNnAj3UpOcBJEjl55w
fJnoxj4dK6FeBb0b5vokOWYbVtTJXA8GmMhtvKlpM1r18fxSCEgxPcpJuzpvbIWf
kGcZFAhamcZbBw4CX3hVYr12p2wrkPCPdl5aZQ/AMnzW2GOPtYehw/WAvLatHfzk
q4Ljwt89ByJrBSbWLHOx4a39B+IbIsTuHgplMWHG/M2ZjHlT+un1tjFIVz+ntNd/
T3yJmggx6nxyUG5aZNOI22OiKKSFAY5UawBf+QIHAg6NJNlT845y6TIX7NbI4euK
v8frWKf9+85CpXFf6fEBIU9GIAXn6FaaUlrWLJ7oEROnb992RsLYsBWAXprHHr1y
eiId1JnjmX/RIzd2NV5XzUV102O/RP4KfZ06QsbGl8i5WmER7OJMnLxo3UIehnVX
CxKHt253tdsgpcJq5VjGrR1qFhAXcTApe5OJsmotT7/VLauSmok3vtqKuFjIs7oY
/mClIuY52VtQNXStxAoUF9LGpSppG5ushuvnkksslP/mXeBF6GlCL1phLgJPRsNM
LxxROjhzNqHpKYYfJ70/mcoG7NcyeBvi45PPjns0ixIdLxtHRY7KzEb/jGpjySXy
l91m2DTDHdtur/BJ8sf8zQSE1Imy5hA3/bMIziuBs2MSABFNpJiKVmAsodPTSQXb
FAS2zAZeE9494iAn+4DPzN7n8+zWf5q+CVoIHTAL1KEuKodVmCeuFXZsKt0AMeuT
zEfXY4civrHK7iNvcK76/+/TUBftQORwXj/gixwmILXrgB6j+kY2stwkcyaRCdOd
s3WsZSpYpJNwWq8D3jP2jGim+6ljBtHYzxS5PaKoYD7FfmNhDh7jx7aXBtAlr03W
Nl71+dijIadb6wrOuMA+PJc8rvIl0/t8lkyyLj6bVuOuMbD/vs8AbXhVuNOuugSx
+OU6cDgrWDPjFGO0oUkUhGWtIhqA3kip10tcRU1wq9Z2GWVc5XXiXT4whQn1MnAw
ttOFOrD2ZGZc0N+VPNlhhTajEfPDCf0jHvxwFfwSo0qgiSOXIOSc6Yzt0osKcwty
tV4ItAO5IeNrrkWhFsKKm4Hpwr+Kt/s6TEQUWCRdwAQoWs0TV2BUZGmXz+SHsvLt
eRsSi9KNKoMkS2wpgXLYAthJXvbKBg9a0p9gzd+DS1WMMmFEWyJR1rvhETHrZX8N
+o7Wj0p61nXs/rQsmnJJfMvkc4B3Z4ogoLHrcz9I4KlFFZxXRYbD9X+DC2Mhzngi
E4Xj9tuYGXqOAJaaKMz/CnV3nNukLhN+DONqQhV0w3DUNsRX073/ikxyIe3jVSHd
LdQC64jGaNLXppnBeMLG16BMo7V1EZsYYB4tMNCZ90H36TfpNNlgoP5UJA8SvZRS
qJWAXLUDVmBC3PIZSDA+h9oUC0R5BQ1OMNjkpF41MxNn2buCdbQjAAo1niIL/1vd
iOM5zgAISpt14uDZ8+oxPQP1JnarIhT6xXm4PdrV8zuoY+LvpaSFDbrS7F354lA8
8dXbFOCerJPGxTt4ks471fLxbt5Odcyu47XCOOSkAcG0WTQ2TGB4wfbEmh0FBhdz
x4TjNizSbvPMuOeaVYsqc2SxI8G0fJnK3kByDh/asYHYNUY4S5e0sRTIsgQexj+i
WVrHkaBUQ2gRY4GQkvrY4GqvfLe2glwjqdl2IKHX68d3hduleXdkIo1HmPMrq9Vh
KSageGvmBMZq75tl3togWfzXG4bA5YMKCBZkNPqKagrrEwnZPb5xJW0VhFj1M3H+
NAwwnvjUCAOiTqvLJx9rXfYkgroDGilHCZfbppI6jOnOUCpygd10GRJsiw6jXRSq
FO4eb4Fmz80UOp/IkDYrohCUqinhlSHZkQiqrGqDBVA3X2JUaoBpvRkDmoA4/gcY
MTa+EayFpBwG3mWrw4fkIOpy2PE02InbzH2C1E7MtmLDsz6zem2h+60KjepgMyBw
pNlUH0wkn7fsL9+wnBgTq++MWfhxIcvn1mS1CjASKbdDGrL6pf4vDrWvHnqFT6ko
igyXnNS6DKN+WUBGtf2tSCGZpW0XIF0ynJbaE05uGQsYADKvWa/nvSfLkraO7sD9
Mb8UP3a4WREilqqLMtG4vzbkXFTcsCHeuHWCrF7UKYec0lycyOha6VJklbhY5Zi5
wCt5IBXeU0U44WqAp9zBP0kwANE4QBVFS5PqkEMQcDSS5E7HPlY9cE0VXKGmrsVw
KGFpyLZ9Aar+hXawK0qe6u1z0tHrqG0yhnxizKRrGYEalCbNVPDYYRtFY78RUIPr
+6Rd/Y6QWJzMhJK3bZ0LfBX4e6ChGz975RGmibZIixZrvFptEy15JA60zEIjZ3ty
a5QjRHXpRcgw9Uf4tF+AqBG6L4MXadBMLl6GXHDbkGvwvniBruPKr4euJpMNshez
ePCZr18M16knuTD9YPotZjMnyY3yNgd40KBzK+Yw3bRbAICwDj8k6ncRc2B+6Xwf
wjngIGvl0HLAICzBLGBz35i/JJa2+2tnJkGYl3Owt4sTtZl/0OwNiZ0m5S7Q7KwX
RMVmynC1c4drxiZcKWsUV/6vLyHLRZ7sALHSNSnlfBz1AvkBpG+yyc7VELWg7hdj
TEA0FUtIoIsQJZVwxn5VKBH+k0m63QodWsS0LFi1RcBcMNpNBMFTlpZvdALh/C2K
QOyERclqeoh6IsPQy9xPxLVA4x67vh4q1sry2xEd3/zfcqoHBbeS3WTK9Pxi/nlY
9aNg+xj+4LDJVUhbKK2ZCvyP6qBJMmDO4EMKze0+P7ntMa9aYzh/r861vJVpmSXH
4U85ANj/EOYukJ395zcPgliwGnPpPyvOMDAPPtVfnEMtqqbeZcrqAIn3ZOJx9Iqa
CAOUDg64OfORQQ314uwxKfIKQLq5uesl2tH1WEZbcC9W9wfdV1mKenF6ffttkQ+h
yBN+/S4fAU0pSWhAb+v3SztbJr5K41D4y2pUQYVaFccVIvs1iDxrvqNt8QLCtgHd
Q9/iMukwhDPH+VbSZ2x27pVFuqT60r+K/Ist8JEfGieO3UEwu7fRejcByZkFcls8
/puxtUOAn6mPqdSJb2dGrW8PTrVkAXWcHMBIYfMMRuBp+hkKwOcA/+Fbe5hWQWgC
k13phGnA48eaKOulXxa25FCAVsbSa0DyPU3gutVuGAZnZipnzfCD45LgrROzhV+3
IgIJuJ+yTxDk1ckyrcEkXYwj2qkXk7u2Rcgj3NxqlqvaxUrSzdjtelhqiRLPCkes
pxF16jKmbXviCbU3ETb1hD0QxdSsOFCwpCzMlBZdM0xwl7Zq72hbW3YoxjPjvCpi
qxA+Y50/3qOdW/xShsFHv7+oj5x7UyyORa4n3zJAlzZqtDHVRtidPZ2zriyLdnms
5LJH45ByRkon603BNNnIZjM2TUxJk0jWXKIMleilzcJMRqYS3POKusU+pmPTKJd5
W2RI5p+ZTW6EezBU/1VhkKKHxp/SEGkLCJjBTJBl9Zd+JUYtrboJD1FI7swKJ7or
ZejEEG6UNJEGJ5lQg1OkntcItNcDb8tcnuybU9acNndDEYnCZtrCPyoBUc+RnU/i
Ba/HJyxHiAV/UWnfL6vXbtfKLmvzz/EF3sxEDwgm4Y9P6VtilOKY/pLw5mAMX3FE
UEtxOimKzx8SQ/5s89hCyZR1gmHdcjegSUWfZeUNKgkFE7ijmpdyzc08dBhdXamv
AEwFYJXlBUTBin5L1jq5rm45xpYIUIqSwKXyajWKntK0GF1ygu+qIg6YPNJxF3ZT
mUdSXt0ALz2YZLK5Li74wmeaGOnNxLGtGko3fH7wpIIWE4r69+DtWmYYLF6i/qrR
Oh4J8xQh+M+PVeit+LbP30DJaq6C5BnPfshLVvg0L/w9eemZt0UZ4evu8d4gtTj0
XQZe9h6AUEoXL2I8GgoQYw1lqmPyqsLKkiYclKFii3v6xVA5C3BSFBxmju/KS9Tw
fwOlFUkGRGn6sJcYyeJ+e0s1g/F7YA2EXOTy0pJuL8I8NmgeVlf/WWxHuCyLJBPV
7KoG9AeAhp2nkFGb2TrKsC+GjtjEo/JlI6NGpLXh9Sl3Me75Y+WwyNfQlL+4l0ao
qMFc+3Wft71EjbtBczTyipw1tasPVWPDuugciKIcKTmY2x9ezhKtykC9TfYnYYk6
p2AAXAQZKpV04PVIzN7Ib90accp/U8P9bbPGsj6Ukjall0+wu73PVMfSK3/MH3g1
lsmQlbfTOs33XD7xwJUfF0m+yjIIc7wNdQSrGsHvgvkIKufJQAfY7NKr+vFZIpmO
G3ssqswRylzRvyVTlN9Ba5VUSLfngjLVTB5YQ7xGkdmXyyJJMtBnZIFx9X+auNQx
tHkg9fbEr5pdPnm7NJrnEWebxnNg/AMpXsw32xC0JJl03npy/BrQb7Pr3JVFIxBx
S4UAbMY4iEsDoYlvBYfsJs9Xjlsd1CvMlw7qH36VfiiKoLYjlLYUyPgiYc9hf3iE
J996kfuMqtZ1CYroVvQ4kn30E4ShRzlA/Gk2/2PDAizigkXrMF+4wZ0QLIGz/S2G
60e96Thum7XG2vOBhHC1Jv3zy3cVm2voXltzQ2eOlwUoZAHLm6Q9ShiA3WmkTRd8
2fhnTBGxY3BJHXt6rWHNrKrtIqTMa7PSTBN3fA8UuBYoHgVcNrVSvnTP0U47J+a5
dXF6pYxoS0yx6dvBsoW9RbGbgCgSwbDZfA4SGnKyyEr0hazqceqqBmq8K6ILGOOU
rFtSGLftR5nUH3pdaybCtSo0oSvyOENKq41n4zN06xEmpJMG5Ah5D9v/+0DlVhSa
m/wkVOONfyPIYHnNiculxknoepzbAhIde3hNNXqpQ618q0RE+Tt45xrj4XG9Zh3R
L8/wCI8KdV5HklV4jxnqIgR6SCBk9VT4dyCBaUeZODNtfEa/XFQbxKUkCYxCqcxY
WVgwD+zQPbW3PxiP13L31c1uk+6QyV9wOvnrofMyC2aS3LOmd9a70pZdSxAyOrmK
JRqPNbgyWueHXWKo+lnrlFMqq0y2Lp111OnfRh403ZtOdlwydBY2KJyxFAaARt76
cFXvMW9CxSgCs/Z2l6vSySwplLE3v0Rlgm8sag9YJfuBxCKXLeWWEK5RyGTicUm7
0pqqB1H4bk/tW1Y1XMoEBkX/3z/0HVSV3iDUnnf5bXwsaBlPxNeOP/upIIl2SL6V
DrvengBe+dvpnEcowHW51ktQ7lR8pAJoEZ4qemZX3WMljJ3mjhdbSPc7kb7kvGir
0ZkqB/70zAlZmC8UUEXVtE3Yss6syGz4ShPWtKpMA+tv4Vt3tK8iaaGDyn9JqGur
hcYxdBKYDUJ6X/F6XxLLhKvNAzKUURm4tbBvbz5bcCTPvPD/TzJOkO6w+ZShn9Sg
NCN3KyhMK3mNog9AuHn6eDruHQtHUrS/Uv9QX4d+Yk3VBrQc5HSZwEcgj2gzojZY
PPjzBG92RLn4rYYOjFDRxkG3DTK/uNFUlU8+2/hCh14zqeM97IyR9EE1SeYjeyfG
bYfc2z3VE+xxGMjDliAfaZFg+C1hkUfzfE8eq8XgKUIfyBfYzpQ/cXqgkDl07w9J
2m+4LmGSfnw/gi/wcJSExMh+noNFl7FgT4xIa/ldtL4fcCE/VHY94WmeM6Mquo/q
HN30r4UQo+31KppHqbKnOCj0a3vVbs3pb4jKiqqCkyZSmXeuoTj4L5d0M6AFsSdW
NExuLm1m41XK3SdRL4Sll3n7iLEgGcZBHFsnLVw6VsHr7FYWp7BzzTjrMqmgPb6p
igRmfuSLxq8kVPKzpZRsj2722qiCHnS9qRkfZKnufyHpDLx7XR24/jZFjR+09WJX
hW5pjrGyBqPy0wId08PHfE0+P+qDo5/PEf5zgFUFMPoNiQY16MdPma0G82rrIekx
cOjr28yeHI4B7el/Nyc0YBc6n8tHv252d9FXzDI+RffymcrTknThZzhi0EcfuNJo
aTdURRWnvtgwc5ujn+N1rs29oiG3OYvSmCAp9msIPDpbAn7iL152I2JTK5ocKjwk
z1AHgDX5Mic5aeivx1Ox+GC1QKPYp5QnvJU8AfykZLTpYPpXJD0PaJ/YrlTpMiNr
xzihwJhaRrg8X/FuO3KxCDRQ6Mkfi0bEO+UlPHQn48t7GxgKK5JR4W0MhH041upq
/SmuXRAQT84mm6ArMB9zgMFhsUbIqhse6uMoJzQazBNTSjUJqB/IG4U5N/Fl147v
Iuk4DbnSLtv9OGysiPV4eUZKamym8n5MiUyx12ehIa3dwIePW3ADxfTbVf7iG23K
ATQiEKJxcxRRFHkD1f6cvF6Z+046gcOi/Ksgni37+h6fhCYEIgxgYaMA1J5ayGdi
ua7C3CCxlSvPmJx4AyPzOfalPU2Gte5g1GvYht2mct+fSTV+E2UsYR+yCC1FSG6k
lXO7a6BLVDgdfSh+tWuG07dnlp1Ad0GH6sZ2xuFq8OvBS1GNxbgQzD3c7ftAd5sG
2wXPEA+prHB50yw67fljfgPkVUP5yAu1qJGR+t9OoTbaoh/r+Yg4pj3lLa1ElzVV
gYgc9/NZa/rSfvjZewew8slwH61xZ2zHvWAAifpoLigxKwsBnSdX8twjP2iHZx5X
HpCIb/wnxHp4o54OwpkqLvwkJr8QrVb8vJ7H9TqFjFEi0d5izJ6Zsw5uOGdWk7JX
2cJcttV/ENpvpizEn4yeSlr9x4gVZ2+RNilMFKddXMMH3ti+YfqCZkLAPQrkQRoK
z1g44WMxcy4hchGm1AQFj+/fqExar65B8aaxVRa4wo38CSsgf3tj1suR7RPdH+hK
7cwelDMyyp8ecvMp4m96Mk+mmeIi1URNV8//5M8w/4F5h9jRdBQcd1fDo1BrZV0w
26n2Ha+XIfWLWveFsn3tIC7nvGzNcqR210gReU5eaY1pr3KUYKTZX3McZaCJ2bql
/cC+x+32QQO3IQL9UFlHJQ13pBo9RAJCXjU0qEDf+Yokjvs9URz2rwrr4J93fyJq
k39yu2nFBllDtg6BdEjvcU/0maGfdPjt8GD14iBLTwpAFHxtML5gkjVsY6IlN2iu
OFZ4/Aa+gKXIfLdJsOFKgiirj+gb5PYML2Nq446jCifUlZyRHBy9Kbabfa1bdSv/
PNZCbv7u4rmKPpaiJWMa3zmVjtfHn4tJWm7VzF9KdLzkOv/xF9TZ3vyhwvucNoK8
mz9LgnQzZW9COyTuE4T6r7rGeVFG2Sh+YFj2qn8uWBLVuVxcZPXA+xpGcVdxNB2/
Rf2pP1GIYlNb0Zh0LbutgkteCPCeawFGaJGNnIdE+E4lpvkSluGrYryr7N323jf2
EArCviU4ns6aGwDv/LUBksNebJaPV7cz1UAGsHsZaQA51jE3yWefZVCtms7iNlxW
R1W+I+aCAX4mnLbWKe0v8AxFYs+zJiMiHUFEDOrRlOrBPBSKuC0v7Yl9wl2zGSgt
QlbUNRCfGIyU4BTEHUFp6CMoFrF1fNk65vsDNXZbb54Xu14SdMHJxDDKXEdR4+Dj
6iYJPvxj5dNSX81i0Hi0qCszV6hB4aLFwKEP+UoP3Ef0uP0U74lYom2Edvi6Zp2E
SouGuaasKh4MQ4aH/NPmK9sIASY+uPmqO16BWCDA694np4K5hb1ZOVf0Saeb/F5T
3mGR75DfVO1GHa8rMGmyC2hZOkbkUy3FN8Zy7ur7bH7HHgOOCg00kSSuRPUHGiUo
s4bTVAMrykpewc16icdGl3F1BudkKLk4K99JFD3bmay0oCaftJxXe1655iuL4KzD
H0tQCQgN9+Hsott3RzpB7mtdJZ8LN0OBqrA3KNbBaceebdyibI2dUauiwYTR6JIW
XvHrDk67zY5hOI2w6thjw4pkDEAsi37OGotFzeEhvaAG5XHfLLumgy/bhMJYcGWa
6Nw13ixNWeQND/hmEkbdMRcZLRabz/X4swPz2NQQqspMI7EJPz1ot/U4KTsJvIob
Ot96tvM4uosDAitR7HVghn0i2fR44BgI03zkTKPnwpbkLJF6PMChlh8A4Jvb+Zjy
X7CcjxtXyGMRr2IoSrDDHN00RGMW24l4zUITHHtfvrNhndWChFclxq0hUtusNQhX
FIYAMgyxF2+fb7wk8BCk0oJK4lFVCAaSIOyhFwVZz64OgJq6dg8VluWL80rG9002
xpK8k9yvQyMxqIFYPZmjx2+Xj/2dYYQzqkRoaEe0yFHxXO3xb5e/f8OVqDzmjAjo
adN6eAARFWyQzzNskxg3l9hSwuD9F2aSr1ng6r7jZyNwCosBgG6OXC24WIXPJko9
iKLOB9FaLpLDpacxi+k0igUBcpSy/sI3s1KvWyASS333zeITeCfdh93TELzf4CcK
L00vTS7of7fM2Zr9+pLP1lKWGTHbanD1tkW0GvaRwYt4YHJQrschdvQvmqvTAnAR
1t3C9hOwb6BHFfUwXJCUPo9SkmUknPja4klvwDVD12kUq0tyqXOD9eHV3NaNJ38y
0v/NU2vmVzZJJEdTv1bOeS1EANiJDoE0sNb5VZtiuLqSlRtc2jLI7XKy6azdP9sr
vsjPHk8oczA6ujDqENI5OUOwf+hCdIDmw+HK1jfEsxOnMfKZ4TgNVwW0jOQ81IYd
cYA3Rjz7PVzbNpS9LM2XuBMB5MiYKt1IXq1CzWbQfn+NuuUEraT9r6u+OcRz32r7
cruTqv4AOSf9qodegetPpTrD1irGcET2vph9o/VxxgL1T1ulTHKpTZRzYaTex11/
T75lQrHL+f8KLKdosLwuCsUtB9mwx7b/EsetpXK0BoBOQIGKPAmC2OeV5BbPgEZS
m5G/xpkuRDckBN1QVBt+5Ncu0x1xS81I+Fu13jLzTPWcIpuKI91laV91+AT4gliw
VV1Ft4yD6UjJCx865+zsvmgWt723Gcl4vDhj38g4JE1AVLIMzd2YCzAAyORNuv3t
B530wGmQosMrOCz+oMbxDDbiaE5Ey/CTIexx7uI1RqHrBf6ieDkI6Z3QJThpEC+j
o/pINmySQWe9NXSxtYmx1Hy9/EN5AP19iTZhbDcrahXCsghv0N3fqdcDwvHEFgJ3
q+WK3GD/kU6cke0Qg8C1dGv9SeJb8gonZpJtNK1xrYrt8tbSeJ11G3J+TYsEQiIG
HtWeaz4wsq0i19+Lchw/40sTqnEJ+sS8PZPRxBbctj7+TeLJRBHlPu/a58IrDyiQ
phQZ4npfUd/jVfBi0UQW/No3V4vrKgkAljX1y+RCjodlk7ESwldEHjd8ZEr2nnm2
u9RSO1AYVrpb2uB7BtgyIsiMj2u6xxeYppMgfYhVtwWvkIayp+5pD9nn3i3F2M13
zxS5yZLh9qzmIKlPSqL0zOLMSlkCGDVYECx8FEo/21mAfVYyOhslPPEMkFHFKtYA
VmTD71GkjFqGkyyiwjVyJKPyGKRvhfbp3HpX1xBKtpRRT5fQoSvS0N6n78Zbplko
hMwgoa/+NJhzHuybNV8VYP1sjdNNKty5k2cLzdMMKSpT7l6eg74+PwJ9nK9Tr0WU
CtHZUa9dp43RLnEz3ltBEbz4s2f3OLZSpmzPT+1XhjT2BG1X6JP5gUx/5gAM0x4r
wvpMeC3acd2h9biQ0t/RWfX80xqVHfXiGVXxBnvIwp3YnPNS2dbenfQMVeB3LQie
zjmlQLcSJueMs152QA/QW2L56hu0Ny+rzIN87So26X9Ah9U/SIIvBNQ+D15GKK+h
UPUn3dwKpcTzO9XoxB3K8X0MgE9Cr5oA8XgEUvXKXyvcRPO13S1KrNqW9de1wyPo
mQIsREpp9J6MaM8HJ0So5e5jpRXUPoxJAOn5t5vAGlLGVD6PRB+KVtjwaVQJ8/VK
XrWj445DsJWPGNivWKmIZosZeeuiHxGQwWF5lgha1urwvuKNntb34jEFjueoKjKG
aC1s5z5Qvewwk/lXD35jYGahE/DcmAtjz6paqFwu11ZFgt4mzGT9+AKJLCTjeBgL
kr+9C91B2QPjupgDba5drIGpS4G9r69dN1UP1MwLx3v9dL/7UyRrEI1Yu14Zmnk8
Fo2MQp1ph+rv/pmxQHOs+1rfi2mnyRxwoefkETBRk2omDXPXdqJm4fhVDbAgYKT5
5qH076NKBNcrO9uE9td0tdhB+JxIb2MpsVIHLvP0Zapk+tLPUqaWdzUw4veI10j4
ydXNNPqMO31HEADEHInNrQNl1c0qIyclMVBJioYGQK+7CHqH0abfJcVQJXRtHmWW
qXMuX9LnBeAmJ0/0dY/+RRdP9vZ6eI474Vu+1tEDWcXpgs4087zMBuk/din2+uZb
roCZSwzi93jId9d/S+xSxR7awakHNL9sXaCq7v4i8JkmW8/kqg1cTITPUKCSnMJ6
XY8MXGo1EXBkWpz42rNyxF+55CS2mGF6bfBizzyLJ3BAHmAoefM6Dwi7gNH7GFUg
K/COI2+Pcsy1mUjDv0shZ6RnCeVSy2AMymE/1fsvOzpNbV6kwelswICgC/sJl4rN
J1Go92jCFZu3AdmbB4aIy2YTpB2AC5UoavsL/AAAq1qnWCxV89eAQhrdz/8D7Dbm
VG7U+r8KvMy/fDtWs7DCsetEPQVP2j6HOSPLCUJRkkqr+8+jXHAHlo1579OCwbzY
ST9gdER6VSgmXSW37f4KLujprZP0F13Bt2ADGz1uh+w/gGmEoNBw4c2DdK4idhGp
Y9AFT5g89DwwxGApM6dahFn8yJbPF1sijZAEy5pkSBuxDvSUfTNWeD6NbSPyCSKO
Db9msEjxJUM6q9HtTP4aqudE7nD/sytiU5EHn4CHMHQE8FGHg5fF6KEbMg5lntzn
DmqDaoJbGPtp5KuF47ToHT0eDTbyWrNcGwHtvGmDFUXqslQ1pD2VY9W4smBafb6m
9yvou4KPB50Bf4HBHoc4oeO4Ka2jP9l0XHmuzVoSQ1eb8CrR6AzlUriq+XOpdjRA
xm+heQ/pf0CpDkpBTgMaJoaVdjygcjlV6LcrfByn37n6V59SR0h23Gh0c3x7C4bV
vli6WBohoCF86HVp8mZ8VP6RiLAykqAJmZpOyuRpPr0R+RIZI8BrlmM3rjUOqWfh
oGjPH1ZPE4nK2gd+fzlHu4prmn+F3hM/Gzj5AiOShOw85lIBtsCnsJFw7pWuMdn0
IDC9qPQsW15drJwssdQnyWeFFW1sZ6TTOfanL62frrOGa89Xgk1WZ8+bfcAhx87p
GukP1wJNcjSSoOoDSFK3MStrqh1B1iiyMPDP9Tn6q1Ccki5G0ZBNf+oYk5kXM3Kw
VqtgY2ahO2jjoAArnC2a5QEF/vyBCNN68fQcvLVDSSmnrUb7N2jNkP8QzRVkZbrw
beVC+Y9zH2PIseOw/EA09NLLuMJ0/Fz7yLflqV/JnCkwwrO64Boi6Co8ggERCrr6
y3ChXoKP9UMr/cocT3wM2Ff/Vm4J9/iJaLITvKAa21cZH4ACnnpEM43JLRqJ1FrA
6KB/ZV1jhyPil1tdiwVVN+HG1xDi+meABvkc3+tp5UdvxmzYLsWwIdESy94q6U86
0Qk1hnl4AffOa5ebZQIu63G6qYtX56H0oiqsgQFHJe8fZmN5uqRpBPX8hqcqT4QR
tDb3UEltD7AsHnh2epMFe88CPOdQJRwrRxRSqZp9WIFuL1IWj4PlwP/p4ylWQ/Ka
FmVjojiLejbHbRrRCH4UMGAE9wOg0NqJrrbcwPUNNIUBhgmVGLzaNLwfMUf/k8+b
jhBWZPUM0hKjSIq9jxZF2NvURA93H+/jzKSrYDWngbFiBiF5n/7qmoR26gfmjLUd
knUNcByeOPAr/ocCTlowPXWISScWjercveqFon/BmR3ZLSfyIK3om9bibzrGC2bn
aLnTPk4nsnTJAKtLOB+sV+Au/AVS3NmoltQllPA+EipcIMFnxCP39JmZg5br8NTj
3XUHP+ZNa4rRat7qSfKHBvoykNYux6q+jhhbcxzVGPiu4oxPkKhgTVZ8uDfNNf2n
XOgEEtZkK2pL2ohpo3Bp7JpMxR4DmqYZQGqNuCPsPVm8aSzqwrX3QGfnIPhBh6om
+HqFjq5lvvN6DeHBpPJaUVAU/mBMlanHo7Ggk2iRdQAZzSuvQ+DkBD9bDj1WIzs+
MGWCdZ0etseP/xl1hiPXdD6Fvw3QvVNGfAtuVwodKtB6wuqUn2xhpqsAMwjbz6X7
wi2823Jruvn1mELTkinmczeVplOq9YGQq0V7VvQVyeFST5Da02G+O/hlsdry9MBv
KBRgJ1RRe81Tj+u2UarVeJ0ObFDFl8C/ggvYOoEVawKr5JA8XGnV1nDNQUjGVQkF
X7sELWRpkwXXrzdnmJZXX35EqcZ9hRiqbmhYoU1DOL2Vf5gtTvHCaZocq2JCvhHQ
oFh7+HNNy2KXljNWl0T4xscY31tQUVNnU76sKA0QsACsJ1AHPM2/7OkqXtbFiwri
dTUA8oY3v6wDgALjkASe9YkAvEqOAliYRVt1lFn+uL5JjmGgfYjLaH+dFG9y34Ia
suO0rLLxu+iS96Ho3hPAw8A1W9c9LiPFfS5N6D3c+BeDngRkS+WIuMnnf/CrOxZT
IaiiAxD79AJ8NzPybjDSj02yOke+3la0rxSi0SaAqB435Cr1oH5lskNjHBfE2Nq9
Gg2uo0I36xyJM37fI2kPSmjibMMNlmSqf5r2JdEAP0WP4Jspy/0yFBZUPULUNz3s
kseTY3lt/4KgH6KHHi2tnl4jh8eCsjOEARVgso/2HFWqGE3hHU/caMV5gYAnM95D
dDt738c9eGlOOE/3CkHMKWQsVyxGaQanzDyBvJ5UMakYMMpleHpzJCQVzUbQh7Dd
pslpf4x7ovjuYM4FFVY407lEinCErbfbffsstDT1vWxX2QmGXPtnuEIIvIEDgffq
gDzcKDDI8fPxUSeN0Gbz/mMFG1XIKDEjXu2KduQlEYLgrwkTRAiQrRLvFe4OnM3q
cbXmTnNZFofhiwFz9kfQvoWkhFeci++SMGFW6DortTG5fIK1e3nH6zNq08+x+H93
upMgc1Q8ZU2HjoSQHgRjp2a5YUbHnPLLmTija8gG04R6wYM9TZSBHY530ZUJQxzP
IemDalniGoMD1C1Hp397hGMMV2gk/VAKjww5ZA5esXV2Wl3Wl0VF50MTJigs5f7b
RHDDUq4daj8hTpKPmotOrhu+WJDgWXhujD5VwtNWFTE+IuVgOnoZpQ5+Bc4/XVd7
Dl/l4oo+5fK/pTYsG1uuHfN4t6eEFGAB4G9sfGX66uRJxQCUC94Nos1R/DD1xUJB
3Gxsu+Y7c3hdkqfRwmJb3usALk2sWdQbbWtXLutcKCmTn/epetNMpk5LBm5aLhy9
byv+oJl7sTjyXiFrEuEfFomPP8rYBc1xDtiFlkG9/uf5dnNnOv+/mX0bPzoLhBgF
fYxdhVzDw49zR1rTqDeGc4htT4pF49esjPZFD7+icipkSLiluW8fXn5raL9qiv+r
YhMWI+qW2uZCk1eYhNqAjRWK1ZvmZRrEe+4taHtPSi2Ez+Rt29MvriZgmflp6nM2
BGEnbnJID3zFfmalZdtED57B+FZp69Mon6d+3YDoTo0ywWNvg1EI3zpTeOGkp8hF
lqwDIdT/f5whBdqP7FB0hW79Hf9Z2UA3EzyeLmvaK740F2W8Zj2Cf7WIDzI7S8gZ
b8qO3WzllcJlW5R9NNp/Ss6MCY6XAR5pVjCN42RKKaDDCvlkJvLne0b6pdqMpao1
FkKVgKswo/V4Z90DpXktpCSrCtkByKDnEyquKk4HXge4jmeEbRAa4bGxaeB0QQH8
Y9idcq9dKgYJFwb/hQLoyVHTkgdo21atRBkJuId8IMghPMruTA8mA8LUuszil945
5advIKW1QCwVruzXjokO2SLPVEZ3K/IoeTXhthPtx77oT9LbwohmGWLrSiZkMrT8
XjkRE8cljPe9G17l0toqio9TJbRFfeFlaRIgWUIj3nFfLz4fBiXdJwdlu9edTPdZ
OAlwBVAq+WRuhHgTIhE55Ww2vuqula5Xz8MUhq9ybor+n5x7HZ0Pnog9EpwNUYvA
2sApNPYqQ1hUpKytYp2a7NbU+Ztw2PQQn1lc7IlpalW8J8Qi1riA7reL1J67IX+J
AsvEyeMAzj1lzAlDAvkEtwkpx+NasialjllOlyaUQJjpmfX7eUHv82tA7Xl987aY
0r0YWxN8kF9yueeD1R6SBifobmVJsjCOIMlWz6vNbtAMno6nUVpebsRtPYLNbKvd
E0csgsGwCwlIOKmp0/cmSypWQBqjKpP9CB4MhMJBhoP2Nc2IsTNBnVgFEAE9/ZUY
sKRcblUTe7+5YjsWMsqAtvPvyfl3OPr4loUMSoK2CkOPWEzzras31u+TB6ItyP7W
Q+RGc3+pNFOdaVM4Imhm5pn5GvFP0sPdVK6aV4bsnvu44/HgQAf01QZpsTz9iEOr
XNKt126kdUlL6gD0MnzRQ6Rf+j7X3GN63VAPqB9QnhVvWk/4wFarD2OxdEJWyuZI
ZfXozPzcv9ZK/BpGan+ICP+bcjnNvAc7bVvMqsshlWagfCpc4Pe8Uc9Wdf+RoyMc
IVvsaD78lNiJ68FSqnfcJlD7S8H0g5KunKIIYTWbGBTr0xNLRPFBq7hGvT/uu6Uz
byulivPvdBOhCFC86L8IjdAVraMxerTGP9b9xTWElatoNn6XjCk9Z+N9t33IukcP
geKlrwJez6h+u4XankEIPL9OJkiNJOWCYPzGJGhKl+mkGPsmEZeebKU+WgR0JfM8
M++YgpQEElemF2skr8WwLqiEHdIxb12ZclQiJrXRdDWN8hv+RJdjaChUp0leqAeD
bx6ZtrG8pyf5WAacWjEjsQagSlaS6AL9eDORKUrk7dM1Swh+lqLbJskp9SInBO94
nozEj5i8vT91F+N4ljnDCzerFdZ19hSwtxweIVynTFm0aoUlNDM5Pyoywl+w/oIE
xX65aSWagXH4WO9YnT625KWzRJztZkGxt5NFfL+DTpmWEfCZ09dX2SsBChzYTEiv
K0U0oJgNBfw1xVUFrCpkZlcWmRqBNLAVPPV7YJ5rkxJANDHNpgHw6lyDpEdue8cS
u+jJ0oyFe2JE6Cm/7EvGSRS6X/OzaHFoN2WK4ofdKGgarJUHXtNn2d0e+w1VlGn6
Uvf4gDa+xsvvSFvTRHUrgEhgzztkwOMPG+u/NTcxy+cLb8/5iylFWmSO9QfOVWGl
3wP4B/eBYPDotefz+Tz6O3wjRhY4q0scN7cj4yHPTo+gOLNmDhL66J/d0Q53ayUC
bWHi6K9E3U74g4pMjsfP0IJTuR0ZRi8ZGbMvYMsUy5VVXcqGi+sIauNRV7pjaDn9
qsi4/YOpmZr4seI+aNM3lhUldL57Hss2ry8tlRLOazjEVIDv72teYGmP7ha3HyOE
qJLW5OvWJUUP3/P7TzEcAoVAnDX5rDVQwUEQgKS5G8q9DtEibMd/m9DviFMTl58C
WrDT/X/O57BfI2qyYZy7lbvAWq4DT6Hiou6Hy6HmqfEjdSMFVZjbbKXjZ5uwZr2G
1QVm4oZZBlyjuBE5quZnn84dsMf+4PZ9TiEtNmg3I+VuIPYd6yXyg3hacPgVyt0m
2CIirN0zzcHoU6g8Jdqn/X6x8lQRjkGwl9YtaZQQzJKIxzbLniWLvkrWeuNdK4ve
rWw1eivif2ADwYZaFPqjCc0uc6C2FM2+Gb0qHkL4P6xi9i2GdQgRocqqYQG+hl/c
/duS9VxIfQCStJw7EFzm0DM+iqUqm98n44V0rAWn5bidS+NvQ030wvJyRRFUyNu4
K4QAipJ3BmE/JFbc0JTIPraPRXME/gSlzio8j/F2GaNMr23euQMzSXoB88J+cJh0
RfAeSsfQSEAInCLrxuXj+uVu6b/5Nl9dlBbn17hk6uBc0XHuazbiBv45H34zJoSB
TNxTHGkpRhVT48m1tpu9VCXhY2KODsH8KZF3UgzyxCs/pjWl0FPZDIl7kNUIbAFh
SInAw+OJ4JmSjKI9CTjh5HG2hqPoWcg72D3uTpvXtr4/8lCtlUUkX3XtBQV3CQln
qN9FyXD19/9MWCJeltRcjC87GzSPjQBA6YvFzSvQGOBK0ItkH1O9YB20LNp9usen
uqdbMeVIqRplY6lrEriGSFrDhG81LREfvF8zxKj6qkwg/6dZ1xrG/DkO+FfUH6d2
l1H36jYSo1jsPKdLrJ/+2g8MFVYMvzZ6DFTiHzT1u400/DaF4sKbcArkEgM55K4+
ac7dMwP6XqqP79W6d15TFEaINmlQ+c//pjp85sGyIJGgCp96KNwDDa7xk2hzTWnF
etVPJ0+8gsoZ3Oe5BYA2zvhLoD8L08SHIVylrp6uZqo0PdqTkwjvmP0JJLSnh5r3
PCfU9TcTo2UtK3lNYgiqxCZdlNcqrVLNoRlFZBfVn1QTeDSfLhm8pWDABZYnJGYe
HgidMLmPskn3dR9WZAoKHDN2Q4pNmBg25WBNCAxZzxmONDgJ5KRr2HAa2t1xS0F7
32DFwyccKm5D4eleQWnmnfDOlHu5Dz91InE54YCj3ae+3qFnReVW9baOtvf4NXKk
m45yZHXTYZCBGajAFX7b89ax41Cmk6ekG/+5CQfsy8CF43J1T5/+q3cyTwejkyqu
vgMmYS9CI9WLZsureMUOGmWUbssKNePosTUG8eb9nb/u6DjgjCPRdrtkyjNRNNPF
6x2Twzq1mGDKcdRoeV1LzVYrA2Wa5OM08U0M43GJOBFskbnR2qet1hmZUg/Nv+Mh
ULwzPuQJ8xFi9cc2Y4KhHHJuWEaUGd5a19iuUYm4ST/kHEyt8hyYb/MsiyYfgK6h
y6avRtG9CrtvkAWBJHUVYJsia4+Gbm6OBjx9p3ERo9jfeizupfVabpxpLbi2f4LH
LszpHXok0SKMovFd61GDf+8eDF5Z2L9H51y58DKNeDplFBWCBlKSp2V/bM3ZNOhw
Ih4OCaY0WIjNGyOAG3JRjlGiYYV0mipBIHAzkvQFsbLJdYR0RoPc0G28TbbK/0D0
4kaw+z+Q4TYmvBaUhYOjvnw+70CsB7KsW12O5Nt05+NIQxogyGAmK5DkdqiZh3WC
UAgF9XEN0Cjg1Oeved5z/XSUWiTzyPkquG3FQxSzFOt6DDifikO+5uEol2xFojxC
6Pjf548Q5gbI1bbQcWaBX5/WfD3ag2TebWyzK6JDxmdQvvg+GSii9V3cMhSx8/sf
TZu/ELip4LukiOQyL2V9BEz084UJXjpYwLg23jHr2vqm/HzLnD7Z4e9fQdkF21qN
8jlM1WpoLyH4/jMmJChH9J1zUJ50bF4QrwmP7+UnPp09m2AY3LFldAe6P9+Qir9x
ScbQ1CKSwxa4BTVzCbNy5E94tsEFAkwXAhasKLbWzTm+ymag3VXpIeh079TDozqC
Oly6zDC3S97QtulnUKlSjQA4Q1YhREkEuncnjVSdHsvruIt+BEeF+etYNYTTgQow
9J4ctZHXucDUxqkuztEuz0q/dY5K4z9a6rC/FN8I9U/osMziaxn7L1yA3Vp0IHUp
9ukj9hyFkPTrSTR4979EYzH+/QSZlhWZcVcdOYoDnABB4jbGm2RSp1TCApDBwHyJ
Ho2JR9vvEf0LD5wI3ZxkxUqmkHl9FKvG9OW+pd0JEpXcxrE+Z0iBeUVICtCGirUS
kCMk89YyN0jXpG3P3ht8/67Gqg+QsO3avaYiBGK5AiIbNGnPnazV57fane1A8pSo
MAuu04Djuyv123Qh6vTYwroS9+/cNROG9ihNzdVshNDq5nZ2jS5Mn0/BUZ5GIq3o
f4n8KJ8F6ci4nvnMgSIszodjKMD22AOPUB75tRXQsIsqwoQkPnoZsHzwjm9l2dpI
M4LCISMRpuMRHIY+nqtswMhqBVDJ+zCs5+uHWnYTFILPo8opwJ18QOre/Lm49sap
MBw3Ke96Qo43M1uRSMGOrBA+i3CEr6hktrlQ2gRkW5ZsxCitjfhoLufedciDyxcW
LscBVjj6GukDLgfQLvmBqYkm9SXdP1lluxcXQOLBDB6oABH9TyPDeTj1fsZuICxj
FRBiZvuRhEB0/3T4ZmCNpHOxk7+hbeoFcrUfRgVD8SUkLUsZp5vmruyvD8d3H6XI
OlouPamDpBaVOJNUNVtxDZNgokjbKG7DX42L9cHSA5hRSxbZ4rjkBrTBuQDasdtN
xjh3dYa41XOIkdgIHnG42z3SmjSq9yeQKZzW/SnDyBzZRJsz1AFoss0odcUF5PW7
ujRJDzLujQyYUZnNq/ywYRNFyLyjAhIyM/QpAW15y7SoMecrluNbIHJceFSSl4YF
wf7payBA4AzQPb5xhC0ggsRUzCzfebX0sdI9nz3abHVWoya0jsLVcQOXqMdezc8N
K8Um3rCSxwm7b9YYApY2sKQKa/zwqKydp1z04AcR1kvHY/cwgNviKn0oqwNLVCAa
gEothHIlBIAGAPmDzVQ7cBdvOf2Gdo2TlxXe4BBcNLUmMcxFZ83EV4FSJ8clevi6
erFgSsk4H4NVBjJnrutB/vgakhQ4lnNVyPsrw4GVQIWRjgzTVw/WTUH2hIiugcH6
AI1NGB/nPBFnwheX/pfdMmvyzzMow5IW4U/32XBLTVFHsD8oAJPLQcRqDuQHF/9p
jNSdOyysq0swLgSz9nm9ety2/6TgxOQWkDG9KYHQTU3BM+/N6laWroVKLwp9l6aY
btIcVO3Dy7F5lp4Eq0GgC78zicshLaXEDUE1XqF5VAgFKeF3NfZ9YT83l8F8HDrD
wQXWTU+xdpq9oE7lPNCk9MTz3u09upmEW61u9NbDnB2CqymoT7QF8L/XV4TmD0Wj
SsgW/mml2bEWXOXnw70YHhjcdMKpBnU5q4fO61W/mro+nRp5JLd5SqEMy4rxOTAC
bYHwIRB/AFY8QquUwlBu/TIGZCf9jL8zt5+E6Odhv3MTpXAI3Zv+dqfJdmML+XNj
3WIZ8Vc+7+jffCq+TDvCtuqbKYB6jxP3WNvxCD9iifh0gE4y9y3o+GQZU+BMQ1e9
CaQE+NxA0PMLqBmvhd8+igcUxoCExn2BzVT52KXYW9fAYVdInXgsppLU0sp8hcyk
uHmbAeGfG8qQAIg+Gly1RSJWJMqwX8bwEZGf/F8IRKOvY/z5wAiL+AeIRnORApHv
Kij2P0lddb5dtmw/ylYY+YM6yMzDKz4kBmP9GnJn7UzbxyeWctX4KtY0QS9hSQVB
EzxOTUeaDnEvHXD1n30y3JT8dDQgNpPyP1RQ4VksibF5VBXbaop25RNYrvwkXrzv
XSrzPWojgCLNMNkYxhpT/KWrIidPvBAxZ5E8NthR/qmo/blKPnW2EPMAkmU5f+sz
PQZjIahoHkdXSECdD+YxzZaqIpYwSdQOgGvnNOUbpR7o6JTFUfG6aKsmnYAD91hu
K7Oo3F3LjXSk4OUvRSzioj0viLnfqBn6G+OgBJ94uEKA6gYrSgcR2rurmL3h8VF+
lAnkxnrTtzq3/9IgcG2mN7gHeRR8k5ZtMcXk3wPOqkWH8HkvxusahapI4B5PL81o
h16fjLd0lIXOIDuXd2paybzC36fEc048EfxCaBP592dBGPWKg7UILU1G3dnbd1If
4SALxHD4AluZGhASNbEfKcdkuNUiWer5kyEVyEgXIHKgndSWYgBCo9RIiUX9xyMc
QbX2X/O1Y3CD8I3g7jGuF5IMVqPYPsK8haYuofgU5qV9Law1SVf5hJJvtZcJ2eI7
ZdrYYrccFtlvuD2npxIoAL3czY9BQ46US2u4u6MgcUQXlXNIT9GfPkkdIPNi/mrZ
S24K21VBWMyRDa1ygCDq7Z419TGUqk0+gpL44+KaovKvy9cSGZjo3uPDjr5KE4EE
9TG6oAwv8thKpwspJMku7meFjEDUCUYTFXGrY7dVxYRtBAGuXz0L4MvSgn+bh9Fx
97fxLF8bHpcl8/pK262z0HKoIzMXBXS+hDtyekLc+t4VPeHW/ilLvEOna9HSAQMr
+IHclv25kKhNwroiVyLPIQA4jpn+crKH4JkL89ffTzKOIdo3LtQn2TB/bRWrLX2e
B5FUG6/baTI8cQdTgvxl4+SVPqmKDOW+OAXMfZwo0cAtWAHiff5L2izzYPoUlgy7
sIHe9O6EX3724SJy9/42qAHeyeLbPBibIyDqYJwW1IsJs03XRM1izF0owccjEYrn
HuHiWUA5MXTbXN4TyEejRQ2xJ1Z1vIgmYN2Tv3RJwoLnKB8VXKfvCzbBexN9AoJL
mxcyfVmsYJgZytA+gsbdEHeK8OSHibvYzenTl8RNAOvEN019t5V/2FCXjI/YS7m4
SXr5xsX5wRn0YHgJ8uLOTVK20Vx4Lv1NB0XPMGHyF2wAjmt+eLumcsHQd+e0xuF8
iund3KKGiOaEHAwQgEBQ7sKE8URGfPQQUGBGRWP0owS0gfMrgai56uBCcjF0IYs1
wmn4yBr0qb0lJAM79YiTOcYSuW2/APhCD/iXHO47bAko0EswqAK9ACKMbGLAT1Wf
vr3O1MIteCfZ2fQoH/r5TtMoAss0aGMgqAZsz1cux/YfSuWDUrsBgUe/QcTolJMm
iHulzb+YkOFk46aoXsQlzDYGamehNwYesDvzaiVzRWU+NqQ1LCA6xcscPs0wgVZa
YRqSPCKoy8DSAUWbszR9ho5n1E8ZiEVhx/KvtLvORsw+IuLzf+sgTVJIMQfOtFa/
7J6EfXdtxnGW2G2tLW8EuhvcXlHS3NGG6kVp55+KLhXIb66qaWytpwZSEa3sFRUC
V1tY3eDZnAMvW/UNJHc6VYhVFFnyKrvgN4/xNEL8CnLmykY9nkt9r71IbiqznkvM
wDf6mCn4VAVG6bB4gQO5yMuYsfguIvDBbGb4uyyIWBS4//M6i2vKLHdDX54SyDW8
3070ewn7oRNjEalv7V/jisGQdeBNfLvIKPNsfiO3hBDOGrZSPhByTO0dMLOxXrlQ
VNUmxQ0GALG1oWYu9c18lPtN12ivghcS/YAoAfYXfODsUf+E59DtWTgndesNQMvm
OzNLsq5pu6P4FypP8n9wJBBYkci8vEwr6vDHn6Jg1W8D4REUCTPRan+A/QFb7dhL
l3Bm2cpuS91OIKfjxIqKMY2Pke2eYRBaoSqAqsxNx2Wt9LJ56sRVPyozGpdeiNQf
htBfET2iJQ9jn4O0jFywFHQFSPhv+CMbqn6XO773tk6Nl4PoHZASU2yLQK1vQy51
nwgx6DymkpzTqcQ6oWr0/G7xkZ2u3sA7RQwmIxJ3j24S3rVUPXs+vLVRpZ3OgLyE
govrSGriB8WBaB058uv4bqfRzAO8ulcp4ZO6ib858VjY60MNyDb5rj7D3A+3nYQP
Zva/O/BvWkGeBtoV5EZElrmybIfBOVOds5+ACmGf6Bd+Efbk+q34tx0gHpjDuSAD
ouwZsqhDr/wMpGHuy3O4lrG9Il0sHcURG6e6yOsjdmVzweFQyc81h3JumM1rHQt0
SveMjcwrbUMd8Xbf2LOVPYNzbLsZVk5tZyVWiRAFxjU/loEri1r8DoDPeYlSip3C
c3l4Noaqd0xpQxTV2DRhypVkJcMQYHqggmXXrUWaIStSWks7xw7NUaTypc4bsh7A
tEaQjSCR+AsrzLmpE2ULsMnGYyPIgd21ekQdXo0D2caQ1d3UlEwB5SkhBVN7rwtF
nOXH+rln3sGqLBkrndrpZ5mcCfqrR+2L7z1Zk6CsIeP+MY6NE6MxoFUzTm5ec+MF
UBSeA7mneVFROrg/p392gDHGYfpY1gjyk1MxvAsRNsWP8JQKHUa7mkTNwviAParz
rby7iTk0WapMWEVp9j4w6GVv2v6ZK2mAfIqUZmQGAN/Mr2tQmbwgfMecegMVzkqS
nH+WzykqiTjm++yTmMvlGYOcqGW2yLrSbZeON2QEOpU30cH81xc6aK2Epr1RHeeV
ERICA/lfqXpUrFkrvubTcJxBTO7DF+PTXv7fG+xKPgTA0Y4509OneHIt6T32xvI5
zvdR6uANfaAwAfD9WKdD/NM2sRrlOslKP1A3klJLhAcZm4LxbhJ6iYEqby307baQ
q1bSCKZSBbL/C1eejCQYdyOhGuf220G02e0gFy4wBSwNYSVe9wqIwHsmJSNTayj2
uEKuwvVhKrvlzW2NJ47BrGLtNC7pDGGQXB/vEWVWnRlkYVJIqqFkQg8j4HaKLDWd
kUR8eDREseaGi2WOSxxeBnUuA1PleinB3GIaOrhqkJkpb/W5TNYp4S5V0sCX1oVg
IgXwQzR1HuhD6MkzZE/eVD2QZefEEpT4jvQSDbyo971GMIXuKNwrc1QvLfmrIK9j
1dWPHomTy3YSuohHCnJpVT+5fc9Uxa0WJcgMJcuIM8J5iWv+qEoMVny6ptrOFxm4
EwC8aoa2tDssO+3hw0jv6a9yaPUGtDpP6fxOMzzgll+PFYWPoMb6MkupePA2fR1I
iYJ2JY8Lkg0dONDkkL19GqJ7MfkFqhoNoyQFxgDbAerqxLbcnHDPUI/6qaauvS8g
SZ2jgkT7TSKNHN7tykJZv7c4Ob3AHlmy1v796TJKcqUzVhQAf8Ktd1A3t15DYBEC
nWkFmyReI4NUATnUpVmtrkAhzPCTV5FsNHRfVGxG2H4WYT0bOQFd0SvDB7shHkOT
cZPuiZmNPETbJvZYerFalCBYA5sc01Hm++Zy9+koIBZyeKaOF/J1hSUshvM2Cy9D
iQ9Tu5F5U9ZVxSaR1gtVGEFNbCGjkaxRlHRZdYfhSFdfcSqbD7IeihOM34wEd9RR
BS0i64vBarCUrd8T0XvFj26c/nX5ngGGoWZMlVJz6PBhmP3mtJWqRmOgj60TBLpK
qspoOh1idhSwkehc3ROECRQJPHytiquCkPpOKm3+KS16ntZz1q2rvqZW6UL0RbKN
b5gkRN1Ba8Js5+m4cZ/IAkxWcA3FqfIKH1hU0D8Ao+aMthuAOMTKgTecXlcbYICc
B/DKDVuIK5O9ALdi4vtl2NjSLaIZB8sbJD6+NMThhv6zT6eMOETgeoScp83OpF8g
AFWjd6C26AINuP+euFLDd1NZow3Kmfi0YushYFy40O5eJBWdBdG9NkFr9wkKsfwt
EjKeNyosyPKTwbuU1JyuberkCqwDwGFoyQ0c1gx6nq+q7xnTKrB1Of54iDi9y4Kh
i9XdcXl/8TIbqYPQSN2FZL2aXd/XMmvDpWI4+cpMbWIVN44zuaFsM4gyYDeeMqs2
jPIUpJ09auKm1d+v7tEHYWrr97mrNM8QV0VUFfgVLaZp8ib6pdzv1Wyq8/h6WFre
5Mq8YcF9eqbtpT0PFQSILDsYE0vZlaj8+nhgbxjYvi0mEKUaPi/5WOigSG0+b4hY
WIfwJtz/hmMmlyzX2Bn6Eg13SVACL0xxm+E8vd+8wcwovugLTBi42iqjvI6GD95x
CV6NJLzDpHcez3Oa8zSVyebZNTZzCZ0KEZtZPg4XapOFmOs0BC8VnZ+jnLYdnXss
TczCCDNcDJp/sljrmnrb2uJ4IS0bOzCq/OgLnYtDfSQ5isI2uEizS/9wtPqDD8cw
8DEvREQnjxJzsgHkSCBs+MPftkFKuaKNp4DA6Zu2IbPDGVWHZejpH4UsruUFNXoC
J3gtkanen0Fg48l79BcrOzt+BQ0rUCoS+0+CKU3AsZY0waQVShru+AV3HhwnTDzl
WPRX0gPp8CdYUGl/0RBj7nfYFkGjBnmJF/SBR9qP3N8mnaVfElPtlFMSpRgkNRMf
8xJR2pusQKFbo6yvEe2lxiQv+s3oiRQFlAzB31j9YkqkGwXxjdyewUtNK34e5TSh
Fs5LOymwhj2Fdzbr6K2GF0SEBJHY8VyuGToSKMCvM0QEjTwWtNfxAECcv6dmgzCL
e9RUGnwo3stNxJhEW4DUpmNcQbP9XPnuFBzPjhOhCKjEAsdWF+d5HhJhZwwidDHJ
mb777tFhLQjM24i6JuMkXxgGtWHkys7yjwYhCO79MI82dlDEBEy5SgBqw1A8zV02
VSicn4Rc3S48+hUgsyutHTcF8jUuvpl5JSaff5EcUp2lUCBc00amNPbuKFlI+w+N
qDritKTsBJSDQ1mWAbr1LkQ381Vxuhqcdu3wPP5umrgTzv4wDDBvujaZMCJQnEBF
mu+ZjN+f6AIFaCKzIxZNP0+TcCUXhn8HhMZp2LgG8FXz99/ojDih73qDJVXPerXo
0frjY7dJOPRLoeqpU1mhs/ut+sSZM01Ce4p7vzdNi0aPmDlbSMagdje9tOLRvAa0
55uCiGExUeFukJLHMN/+xYuMTlpicKZ+tzEMdw7rhbbvWLYpZBFKWVh5bd+/iFvx
7tuR2LJnTeZqg/MZUYpNcE64SNbyqhbF2vYiSXe2ALq5ahRwEhwiCNK5rUVEJ608
/8yWfzlv9peJV6RUYY4ozBkFLI9RUTSs4uaztvxim3uu3Fe+VU2pJ6Y75t0DNUVa
JvDkKlSQ1so1LuO0njN8r1CeMhZTzfryfGqDgOpBRxXaMRuU0MYIi88nYVG8267i
0J3XpJmPnrbv28wIQzyGvceOyLljq1S+qeoBs3SsHPYRh2X3RmL962nfEd8rtKhb
MF1XSrIYX7rF3dOgmatMeeJpCMffZGqfxKR3iB/TPH2qzwk3QoEN7ROMuWOLLQY2
gCkr9PjQvbsg3RH6H9obH1eoGxIccm42xgLdnk9vH1yUvH6+ouNA5Gfde/YU/zHU
MjQJqt/ArFfHAX16Tr/dD2BcJfktCf1/KUEb87ZIlBDb1DHo9q5cGI71xl9Hii8A
F4OcSiIr0zXT9zZmeMpAYCUDsaZ6FaZC2kKVfII333fpSfQlPIMeizX0Hm1uaNdf
wNQVwHKLU2u8XdTJlP4GAA7OF6GFBL57sjIJkWBFcWotWXwiFWn1MJiNdr/p7MF2
lf+gfXw3KHAVRp3n82l5e08TfZQdzcYdRHC++mTtsUzdy6qy2Ut/YB8MSPE1c42o
b6Qcq+3zmFTAScsVevhnVIIOjOVBjfysoIinJbJBTbMLu1MJqusO7XASdgM3w6iH
dKCFOx2bmKUs+UC1WArT8eRwO873BfFzW7ovzFtolwrk/UCtPkySQgtomh7Xv36d
mhD89eR+IWDrrEpc0qrgEe7Mksh8Ea+GlCGZTKlU+cjNLOWbisF7Eh8NbbCQ69DP
NgLKPJU4MHpcH2Ho3lAbcKc59IOHGpSPEFTxugETJepbj38IgH4v2I4ZWcF/nj+P
rauHO0PsWtWBC1+NwhS1hF9Ah8er7YUYnkCCwaICHOg2sMSVEMuJ4dLAc3Mrot4D
KqlcNswNRJeaof39PkcvEzQz38efn2Hg1cmoQkWzNEVRaHTrZdLMMGbzP6I8Ng6p
IlwBPqWQyClnFAWEQ30WjHRGZq6kCjt/BVDflKYM+h14e+u50qB1TsimSWzmjpcu
xcf2Wo5QlVwoDGk1wWsFCBAFv7b/LKe9rtJW2McoOK9yg7Kd+jNKo+aAzAOmQVxQ
ovswoxHN3+iBveYM05Uhi4Zl3AeUv0zVgi4Y9hVko+Zgvecbf6iaqEW3XX7OwBCn
oP8j2d3q3QBeu6OggIK+92LETfkvg6ufKo7ZdPhBMBoabhvFYOofv5SVwUQKglna
eGVkYEIgvbaDdhhgQNwYPeBOpPJ0BP3lkOa96sZoYKOorulhN/en+JHGWJ1f+32R
A0EWJ2oVmy0LPYs8FmtSjpqBCoV22zOsFvUM32tSiAMmQ+xqhARE3ifbhLStcL5m
UWYSRPnA6BC5dNx6TkxtFtV7HR8KjFiK+jGfdbfx7CrYFjkov8uLIi+TTZMz24rF
ADbvIZy87HrMzNOt+xyGUwADZ7FLW5aHRVCHy2OL/WJqorMV8jZEbZrWVIGfkVXL
VBSUfDUPgj7RRsgJDqlpogk+ORLmrKwdGSyEQDdmcBHGtYu+NhQm0EvicUDPU7Xl
HnShZTWjEIAOJMQwj2GH0S8uHiD6Y2pM6GJm/EPdbvU+g2p3VtnQIrOQSRJjMQz+
kdCJcd/qGcETYwziWKMt4r4t2UJIf+4dltQMaJkyOeoOXYwRXiRMBqF3vixT8iWb
zA+lju2ZRowtCcf9wzoIO5RrNAsWJOp/LKSRlrGMcTtCPFfocWZ3FsIT6mlXev8W
KcoZeg17oXeU4W59jwdaEW7HjfA1rzGoqzwGL+LIyl2fG2te1zyzepU9rHXkvwTo
RdkdXpqA93GpGwvzxmUw4kjrEV4jGf8mGTuISjRzPHmf3OFZMXqlj1OUo2bcqPfG
L1omn6o8Eb+t9BdouqAKPgUWFH1U75x9Z0BxfPoCPKDIbn+mbsXfZ/SXX5hL92L+
QTI5cB0KzuxE/NY++8mXv0bvjhTZXIvi7DUN99hVoF758bJ8kZ9Jwo0syJ1tCBim
HPqKOB5biYA6qL6sdTP0mpPyHE/JkbfkxP/0Sq+bai9k6aFTDKO45k+aPHN+GAoJ
2G2Hbf7v4n0W1sIby/QgpjpEcGj3WcxLBQz8Sc2fnJ5G7pI30Dj7HyLWe9IfQ2yL
IBubTWFcz+nu6kOBDwdisDU8/vGB8GCrdtC9GRTjj7Jfw2HJ3fHjxeOqiUDwBtV2
6awcPpOgDfWyWpdbKsuPtG5Llh3/M85AGCJcCZd4GPRMzdeidhFuXrg5dS3I/Lb+
uo9XqU0kckyoDQQVOVGq1M+MvCw1tEogXKKlNG0eoC4f8b/nZDuz9iUrAVRppLfE
HseIOUhYwjCJzrz3kE2nhdNwqJ7sQDsRp5k4xJRdt3RpQNEnSx9Y+0sDJf7/K8jz
pwlG4He4O0cQSqhi07fo7PdTMWgky8V/WfAY5WeIWnjqnk3NqJmaAGazk2GfeWyh
ROBIEL/LHPetS71gsrqdUvZ45LXx0QzJ+HTFCKcvZjNzJYZgtI5s6BvY5Dp7AIrC
QCh92/V44/HGEWfPXzzOAwLt+MXojmX19kthCygUfn2n/Z55uFsGpCKI16cufrj8
8HbORuCzuSwrEIG83NordW/mtLkID9mj1xgLrPEZ5EsRWKbrOSYWRKKbHwRv112p
zzmkZpXqHNfiGt0jRvWsDYiIJdpZV0EYOfAIJj4PFWcJLZiXjaubcMPQaFyG7iN5
78UYeu+X+iicwWM+msOkWPDDKzjSs75lLs34qGZhbHW45ULLrdbjFTj3nBfZ39N0
+09yzqXg1wpeAQi7rNT+ft0qzdHIhiPbIBBGhsmQzHlVBaWYQ9Io3SCtgiY4fjPB
tJFvCcQ3D1NyOtZDEUXoc5Egj3QL9d4lPXuwyBtA7Xkb9M0ciXwzEvypwgNwRi6l
jcMdMvnjGvzRg7MJTntM7SbxC10q+z6jvfJ5dqO/95k3wA4nVGQB1z25o0w5lHVo
Qu/8RZ1jfZjgQxVbQqukQINDhmnah6JkIQBqQ8VoUsBNYKEH9Gp9oEWQwwZ+N9Mh
d9zfdr4stSpBopLvyDyw3W2vC8T4AhmktVGDiK7knONg89DX+Dj1mNYeDwKgXh54
sEuv/grFP/zO7x2H202JJwpheIeh47W+vt3K4cLl3HBKiHCqxX7tPhD/JrDl1Blh
9IVHYHWFXiXkS3SqUvx0pRF15+CNmSoaDUPUgRVxgojxgEWPOE9ECKoR9dVTNrp0
hxnaZJyyrhqKl+FMhSMUIgvB2v8fWuAzzgrlFemvwlTNQqufGrGV1UFpJgxhs/xc
ZAKEahADPuUu8VTnOnSjzW49BoSNLIyvpLUj3C8dNchiuSvIrrkL/K7ncbgCOI0V
JffTZIqSNDFGVyV6IXsFeSxPEiGibwFbwIiqIO5zjlOO21uVfo5wzs4D6B5g9bkb
uhDTGDVgxfG2SwJg2UtM4nuRyPS/E/kxsy3Zz5ukpzwLTPTFM22SM8WdHNChKHtd
DPRfdgQ9x7j6I4ExkvQmnGIr09JhytYXnPGB+ySkVy2l/xFoxolwillJd+70BumO
WfDMhat8H5ZNxtDr05/Py1aheeZMMwIk+fLrjukUaWYjsyb20JhQL+PEwCp8Pg2g
76ySy1zSrSk6Ked7EDItP5swDlHXdiQee6iOmUYDzdIvPtCFnF3qd5+Z1uIFEs3G
J9COO6jt5czoyBESpVnz3gX/HL8MICLoPOVWRuyivHlHikGCC2Z+bfpRohOAcCEq
/yOj6+cSVOU4CLiK3+epifi7juMgE7GBwBdjMMk9/dR2TtGLfaDakqKOcsTj1/FG
sEy8Zpv1djqJuuox5ap1PNIZuyq/KmJkYdKvkc4gitoLManWfz9+IBzJccvt0VNx
2kfIQ1hag5OG+RdHH0Qi+ighKaYH5Syb1kz6zsN/JVYKNKOM83Fm/LC0Tb4qtgqG
yWwuhZFguCE9Ni3cUsk40Py+cHuoy9f7yzVML4ZX//rngUhsMQzzgEzOmluKs7pH
Tw1G7ocsmptCU0c+Aj+3//SBfwSfrFl7sCEkOAgYfI4ZdR226SnmiK9duVymz7Gt
HrzgVISpHIOLKtnL7vmTF503KqS3Ngk0fzvPwSwZ22k5tFpoehLHLL7JX+Fe3VLT
DK/LQrCbZ+5Zgtrn+ma/51GTP9hbj1uR9A1b8I3NAN9l0+5aKnnaqywBDHEFDifS
b5v9XtJ8CTQrHBHjW0nkBI4z8584bTeP+xKHSN1UtWu5Aj1OSLA4vxFR37Y0M3vZ
nRm/L9a1pFJ1n1RrUuDvwiKXC5vi/BkSUbS6pP0sZhr1G/ZH1hqor0yQqbByqW+3
xWcrYGADaEDPsUpsWQwWj1hvO7Kw1+TqDE3vLoJVc8Q3tUo6VxsEHu2Pu/Oz0r5W
LEp06ENTuzXwrcyXOWex2d+kh+DskfGMkwqInYjd8xe7LmfEguEstTOSz31vZ8kU
l9jo/4Kaf4tHyTtKi/4nG2CeG5qsoFL2CIVxSd4zvQxSQL1uXi54M+fpCiaTX8um
lhQKsSmeKEkqxIDkEh6U3rc248VNWKeVSfuqP/3Lb+OME/C/69+R6BwQoHuLRGcC
AslkF0LY3iqIJVR4b0zvTcADZrq3aDZlFWlnOyb3e7N0IQ+83WRybL3FGFmYwb+7
Opdq3MzPoDdns88PgzKW5pxER+v1+olfiksLK20c2zOHjnbvKOeCMQKBOhfa7n/H
AeDbwXsGMjBl4tl5NaK5ZHutjmuhn1V9aDVdfZ/mWF8mSe6HxWOj6EFXk6DJ1Mxl
yf8Lqh8AuCSig+KQjjjy0ijLo2W6t0XGuI6HuEWteIcjb2dnlcfuHXPTVrD7KbD3
bsX6FXZuYVuCKc3AihgS6bMH/DNPxcEwdHLYgGI3wEA6wXq73Rz+q3/sreJbQta4
zFmM48IcYNISQmxmKpY4ADGQLuzn4zsf7WVz8TLRE1aYkJkSyA9xTZhnKPlvgT4B
fzCzAEsHCwVU5puU5TLoNJBlAgGJezZM1P1uyOtZJ22lESdyDK00jZwEy/32CEm3
mSkKcKe0F632rWww4Dx5sE7qgdJ5MpkM7g9NUICiiiXH3v+z7XObfwa3WmUlve7N
8Pu3nEq6W8QbjitZIhfFBhXPUwYbDeS/Pz53GeYpQySBwlV/jcaNB5cwVGGdhoWD
qguiI/1Ol86Oy+oeXqIzzdjaByHC9zsuzhpDV0eKg/y09cMMDqf4ClNKyWqEGaB9
oZO7ivEsgD7ietu53Wcx2beFqS7FeVpL7OwQzZ7E2g2BCBdi6zDnvRKyyKdGJWS6
kEGkXmNM7szROznz2kyi4ddfO/7HeLImKTA4xiszqQxbN5P/h7uLIarwtTupNaGy
A2AVd8Jxg37L+DD4q4o2Aht/U4FLFlccpS9Wlg2FFGtshq2Cfhc1S86K0hnrygVu
26L6CzPYYhpXDgTY+VPS2mhNDCUHUHKq04nRq8Ov4BZx8ZlzxHR2I6GTasWCf/lH
zKUwdGarafXoLCvMrq4Td5AAaV15cqLsaFVwaGgfLvTyHp2FwAvpbbx1R8EBBKrZ
n19CTqvt4CHv2m1sj6ptI6QWPouJEWqs361oPlDIAc4JmzNnO/A9MccVPbN8HStv
d91tzElP/fUjZBOqvskabuNtUPmXBY0A8YQW3HrBJoIsNwGjuKoQkoP6RZn3BOa7
pWMQ+HtpF/O25/EUgrApw34GEo9tg+9o/hgvsMl+o6PGkN23C4vo21fDqYE2cb8f
v1/nGRfFlxO7qEKeXLTx4E8mfiXLcdRxNmtoFKqkJKG2CvWOKBJwO9JLkY/7BbCz
UHl9gRweZZ7g2PvJflpbEPw2RGP34AjQx2rGouUlo5wDb6Olkv4i9uTLBRIgu6A3
yYrt9787vmmLr4int6XP7GuEEe9MUtL3KUrlMVR1QvXKQ6bolOYsIghzWsUAVSkO
SQzqboYEtCs4Z/Dzjk+M75moo8naxOmtMBpskUGmWqFJaRYSI5VDHDpMWUXoJWP+
aUmbq4cD2/Lenm/7iIE3mZkfFoItvpzAyujTKG/+duAE1Xo0a33/DjzKf461xpZI
yRLFA/mi2atrh6u2X70pB72/7CJba43BgSBGXbhl4WmS/tGXo6M2CYG/dqK8xcP/
YXnQrL59GNjhAl6pKlWJWlK9tJ8vcEYM23fe1ITq3ziowIUGKeNp/r7g6dPyYEXv
ZhlbjTIk/EQsSAz/wTYGIsdjGZ7E/NgFe3UtzqP9VnII/ug1WcoR5vvUSQ5APF49
VzGHOQ/3eUAiSOFMxciiOVxk7UA9CXRxoX+4JF8ZXRvxUVRWqcYBbeNYrt6fEIdG
o1EZUuK0jorbdffbb+B/cjONMjmtG2vLeN5TDiRWaH/DYD59x1/8k91Ous6fGlFI
ndraLSGLqWqMhYI/eQcnvb7YJ4q3ltZaYtgA6LA8g2cu/uEkZOiELUmTPTKxABek
t4wZYK9MqePW6XPdosdJFaHzYPxJwwIDCVphnJnK06EnWEkUPS7cRYZ3vRwPbBLH
0XWHmaUzMK6uGifQwx9Pl/Rj3uXAnR5dF0mHXr/FmqEwAi9xYy37ev3M42rSflFY
CRtks6ZIVbP+wkst/IKBnCmt0ed58W+REjdXZYtIcbYSHIiAnW1rm7L9udJ3QX9V
DYniltRsu5IPhXVQuPPdyIXsYkW6/dCX0v8ZI7YT4cERvXjUT1+xTNF2XJs9e8um
tOPP6t9yCu3YvEOURReYZLs4L8K3nQM1goqqGKW90fPJ7mCQqjV6jUN6cceajx/9
sKw4wLv6gUXFHwTiii2qw34GiME6gcbuG9m6h8Of3S19v9JugdvsMMT2tTTY42y1
SaxDSN9plA3kj08kO0D6dK/9m3YlC69MpOhJIWFPyLfCW5TPT2SA4B/f+P7NLs1r
eUrpMF3IYtsi9/up2PffYhalz2GyxFWzpq91PTeUWWRCRkBe08NMu0FmBsg0o6GK
3T2yl5ovWV7I18VyK1dq2D4cs05nqua5t1gV6zrVHaiv9b2JLRSS9yn+5I4m/xRC
Uzec7YsJKCxWfUlQ5Rdxuw0KjbdhLQD0F0oOTkhOVcokugVzQpMof3/EXVG2eVsK
ybhKpXNup45gxNLiQAm7Jt+Q61Sx6rLx5k7PY5KxapGsrJMD+qFBvpGzdkKg2Rk0
4x5wexpD2AQfr1sKOrvFphojk0qNKxwWT79jNuXwB9x2DC87Nt2bulIKk8rJwP7k
o0BSUNoBXMQEa2ufu2VEYSF5wxSxOw7ksqb5Eq3LaduNT2lPonUCFw2zA/URvFGN
iSJm6gBUXQCyMSYgvCHZL0FC5zTW+T1J9NU40XzZCYiHL8mIsKfNF+xK7g8LLHsF
xq/1dNDGBqx9eW/iEo02C6WJOyvtx+3ctiV72WUC8Q0GEbtfssQSFlFhQXQbBSPg
BTu7Tr9q9+tVxDlBNFsSNBsBKrTRGGLMo+Vc4OsEFm1X+Wl/ttGiAATVnXs9OUN6
9+GbJC/j7sCPNh+B/1Xf3rYqR2fzck04VsolyeyPYMJab/2q/enNexp7LCXuVVc3
PsW2NFX6QdXhUj+5ri4dtN1uMP6EuAfBmoNhEXjn55WBlVPQzL3An0/aTsSzzezz
Teu1KDkQWsRxNJHU34eE4v4daKq0/nkVRh5+fYci2cWabbfzSzJZdQow217x873I
2t9K2RTDqB4u/z48FYIh7zk0VpwNICGL0pU5wCnLuos64erdKXMk+QXWxmfm/k1Q
yn4TL6Ok2lLLC37chmiVJCkl/xgjtdslQ+LV6lA2J7Ar+tilwagACT79zrSy2imV
4fNUAojZJBRxYXgJR/0Zl+zIqpbVSXmsIBFHoM+DuZBnV/Md/qPKepKJx+kJ+R/r
hBOLpQeg+iY0q2frUKBN5tdRNz/IzVdMkGKfyQ4c7msw9BmXcMBbWDEQTTZ4mKcX
leAErS9cV3vnW0+wHYoILSxgJYxp46JejdOr5+l2JyXjx4IZuIO1r4yXUYlO5jyX
QtBTEGcMiGtuq5mdupIiFn7UpwiRMDMZwl2j0bXzpo1yyqvTyWdpnnd/ijzLc1La
RySs5KwVB9IR14SI4dYNQqdPJy4Q0KtycyPeHEUtT6tVRqXBBJg3vgjKtLYJYXpZ
VbqkiuvvVwFy/8BBigNupq1pz+Q1Jt0uxS00eE3TPVWaDCdyuhkmTw2ErLJr8Rsh
AocHdoyf566YERYzNQ2BLTpnDSFoRcYGRrtCq5yXjVrbhpn/ja58CTOjHhkXawIL
K8Gn1h7Q2pFVlfmlYzNtS2omvlsl/yINmMKNpcKndU5aDdA+DY3YHEW6NYOqbSqz
PrlFYazlRO9OkrmO7KnGAvrrX8AbpRH5yUlPBlc2duopvB6LK74j4W0CVXXUmiY9
/ri9Su5iUpxzaT/onCCruKe5O5jZTT4a1C81Yj/g75T+KedguuCcOl574GEeWGuX
0+Vau0J+FSxQrrUhcAF+SZqAZqqSDg8U/ICZ5398Z7cG+raVmQziq+LaUQhdwS+1
xpDseolaklCA/+LBa5xruZjGmNnEcwLzN4D6ecIHpvIcdHhEy2Gpc4hf9ee1LVgg
iul3RFkhMyDqs93s/P+aKRZPntazahq94tqW3nB+pj1VryW+i4m0flj9S30M1C8L
lbvL12GOVcT5xXc0DG3eOwLWPV2eIfGN/Kp033aSx7HMzNUeUf0y4nkjpsmQKFsI
xSCH1m8ZoPv/GU7NsWv5UZUCJW2WkuwP0skzADz7JDxbmhnJV4L0XicIbMuRxAuF
aunWLd1d1FUEbw8t1rdPeFkGW94J7S12CCDVin6svk0snumVaf3E4IrsV/eQoIgv
tBf4yrcIvCzBRnuvjumImUQ6nxrsWlNXtMxbUPeAHp5oG2Y+1rzv8s9Xvmj68QE3
LOoNS0K9CwLx59cJpW98OhhYoX6r7oB8rfiqQW/JyCjghQE6rIaYL+5s+UjpdNeI
+5wouJovrmM0qrVsrEz8RQLRT+YemwM0+e26i0YrlfvXx/cKN2JlCLFVtc+FY/3D
oifBxbYUuCZfmfGypkuiqYueR6u6ZVI1R5UpUf88/f5zreT6FSkNgmid7h4J8doW
6dY6TmzkrM/4THi4wBeNGM7JFJGMYMNKopLsyFaE4YerCP/GXldNAQ7Og0Cx77kE
ItOxR1W83az9KDuf0jNU7N6hkFSpbZ5xFIj7bkTKiSawo3q68pltO8s9sOxII/xn
GGbdIDME5axsYZKG4i+kms71VFSeF1U1ozmQjlWJMZy5RXbolKvt7I+7gl4Wzq39
ZFcpq4PAVjbwKP89yvzXBR60cX1iFfL0wNggxcvQq46Tykyajr0FmJYqrCFAIT2p
sYN9jvau6vhV0pT10k8vq+aMwbt276MXtnwIvZR3V8MZ2TF3xBqYVMrrXSKPRYyT
yy18eReKo4pA0HyOffDjRPtqn0D4+HbIBC4LYPC2u04v0h7/kkZcsyl2Opffc4dq
B9gAh/nw+PvsYqP90YsB7WESkAVYqbXrCVElNkKMt6XDqXjXr5RrHAZAuOgjgSsA
EMptt/tALrGfEUVPygOPXN/EcgZqFI844uwlX6RZrCy/AsFVBByJlGn6RykzMXPY
E9Vqs++Y9cF72BNHgXfVgvEz0Fo56sDFQar8+IPTy9F0xDNCSFA75y9Z5gKWuN1P
RkybVDSmxrN/bR4igSx8Q1Nr4XWK8sJEGTZ8H4jtXflLzI7fYBfBRJ7gOpMgqELH
TJtkAbTFL7BaHzgNWTN908jIsaGcaQV5SOSpBxhacU/35twQlIsWq/sE1bDQRcYg
iiZyvzNzjNuHiml3bRdLMguEmFvhCzKeBteHk1Yx3fuzj5eK9/QX1MOjGLP/KgQR
73+el/jx8RgSKrcDzXBd4qKDPCVZOYUea1uNgITLapKWqWjYfmpPlY6/FWIIvWEb
Xs5/TDvmr3komJBifcsSZYOrHg/FDmTTx5VrdWRZr1kyAGHJgco73Twt4rj4C4EY
CAOeP0kNBI7mkFwJVb0dhVBqTlJUspfBpbyMtz5Od2d9nadkoqPUVgk5LoFkASK/
lZxbvSRmRWL3QsxNqENQS79MIItZ8q3UUsSCPS4RVefeKDUurOnhF2hldiulFDuS
XehKgi3EqL2mO0lzfDm8uPyJGUTnfuoJtxASU++K0SI+GV0AWrPPSu6AV0146u/I
4TDMsmpu9h0UZqoeugnw/S8lyfEELI+hVc0/ROcwD8hGFKGKC23A5JjcrOgOF4lM
lxs4ANvq1zzJfgKkNcDzqLS0CmIU8RpAtm7b67TaQIBFp4DGvSprP7aAaMeV+nEK
8291nCC2+ZgJwb4ltK2NEsHm2tZpJLIJiXrkLMU7wzdPEWYaXVOM5D5TU+j//K9Z
Y03TAFaQNy89wQryPQAt2GpPcAfwQlgaAml33NzvxcmbT/Rj4Xrww+WjFCjRZZVv
a+gnSrONjrdkCu0yrK2UjVkczlR9glW5dM1WcCcix0DJoOxGH66FRUw1ncSHGEvH
OHRwEmD2r2Cev71LrZ1Bl13wz2ltVYDvgc62f9Q2UsPKORE76Dd+/XPBMOPER/Re
ED+ddtoQdSl9VPPtP7NhoP2xGGiFMzvJCPjeiy/tlIZ9lY0D/il6Lk+AAK6+qH21
fJ4NR0Oe1Uap3YNH7qxOrgVSqnufb/OAvRKNGIPhXeVk4uAL/J7VyzhqZpXTSxFV
dU0+OUv+buKO6Mx3XAQcWfG5a/kEi61EZ8oim4cZrmeGHGG0NrM25EbSyCMjr7jp
/BeAP+gcacyhx6PFB0aRBfn1N6NMWOQ+kV2Od1aPfzPedm/801R3yHKOir6A5ZFe
L0RjKYmw6uVTkoDcBeusJQlzQTcsMRafHTcSGcNVOdVCC/XOHBS2Cy4vWGrcOe8N
sh9Ywm09Jh+eMlQMFlBx7o8AC8qC+OyExPrFAE+6kRm3Msa1htSQgJ84JVM3Weqy
G12k69xYVt/dpUElV/wbDQxoDiyM2i0OM3QA8q4d91c9UdZIfGA3baQKn+WMhF1f
jaQRLgzANhRbW8w9o/XiYqiGWcUZqwnwUpebRroBjUvY1VdjkpPrTGySfwXhE1NQ
HB0+EBcx01dIyY8cXd3YPICpZq66YXV7050M+WUMQyR1PhN5lwPV+kyv/nuWkao8
XazqoWgpyYtlvsk2FCpKOBvXMJMPaUP6aYq6mR/1ccISmiLF3mo1bllm/ncDPha3
CiCgaZgu+i600uoTDsUTWLLdLyLoBsXddFm3BUceDQfHjG43JcupVzD3SnBfcKJc
uDHDpEtiyC3LCbtU2OyMrUN4vn6wZ5GzRKutQVn7CHTmt82CpT9XU5PCXh642EZf
7S3oNiuqTGwMP0TOhBsctbMdOX93MXnBec3fbESblp/WrD2ojAcfSW1nDHmZIUvP
xWiO/L4P5g0r6VDyCcR0Gc76nlJ56okPyzHOdzpOM++/H4w34d2unDlES9eZbqbe
/AhBqkvouobDRr3aR3q/zOyUkupyKNoqlI6CP+KKPBXkX9SaT2uf3X/DoALu1FDB
7ByOiSGGkPibmUQyaf16fK58SlOI07/nG0PrfqzT+6mCWvHppjJ3MX9sEndFrg0S
lqwIMAC5TYdB9Ok8ZE7Aeyp+QxN4ZFRmRIqg69kgeErTkPAnBA0/3HqaAaomWH36
UHSIhBSiwmSOzQVKS9OwbfJv9i84kDfflnCDhOOhTTSUI7xwNxCpT0em57faR4o/
aXD8teyp0r7wqRa5FFVSeW24y6XB03+gg8nAKJ6574jH1cEmh5VFQyj1Ekho8lpI
FsottsT6PzVmiSE0QR1VwUAOdghX1h5UzUdcQrh3hiZyfdx5mDqXEQotPulCkiL0
t6LHlFNm0Q3HO+xsWSADxtpxMPImxcDM0VxaKdnC7xxWBj9pycGoZWsxlQDEdXWI
707dxNWjhXJkOl1sm219INwLk5Js7IuRRK6fTSlk8Vj47t8SoXBzQHF4OfsiMcBd
OS+2FsK2KbTo3I4yZbykjlvoUVWZkt7wJ4O3upqVP/6b5IzWFBxIiEwFUQ5/qzah
+TvclLMviVuLj7zWzpwvaONp98VCU2pu3vNMEIKd71303/ANardAdDpwrP1x4r6F
RchY0qf0ti6zAne33lHGjjSgNWHQf6EqrIE2nr6xI9WbdxYGEUtgwTHGitp68/Yi
VhDaEjnit+qrM+UASjaxOLhOrzxcfys7lig8vXmRmomnzCxJkBuyJVOEJ8uX4wd+
WgLInlRDn5b5s/1r5ilYLutfG0St4uWWD3MY/NcHg14MX6deP+cKlq9VEIK3zNWw
C4zY/xTSLoesAmaKBFk4rtwe6qJfgYFzyxpyqxDgrJ4r+ZtMNfX4teubKtlDzD4O
+R+KxIK7v/56y21s1YoFbsksYhK5BptQmT8UzgxvIMnCNnIMOaAH6h+ENLsNpXfP
Mvn2h1X9eT4ZqfJ+TV5pxG/k0v/idOD/r1olzGGufNK3zHnRFGRnA9dOxhAQVmd7
oIrevWKVCsPQTn83ZF0OnYKuB5186H5XWDiDU8SJXgoSRwmCqi/5nLmnhhMnQqNP
bPilJJnXgdZSIGAL1dNlOfsBpWJagCli+h09qomMEA/sp2pz0d7WTqMe7vJAgs7C
vVsu9lixUIO9PSstdEzDC7DiBCS/YSDzCD/PVw/62rNLQyeTQa01Rr5UQHSho/JD
mvT5Iat+4E7ajFvjnG5ZXSYIAuFaapqbv7wP9HjbbXn8p8zjuF7QGehFauFUlqdZ
yiEE7MtwI2JFYkMa2OirtecHA0OcUM/J2kiXYEtb9ukxtIE/yI2x2etkxoXuxiJC
6yNsp1c1sIu6xmgSLuWFCWwFmoXHIrGHn2o2YfpXynxi/twmL+eFjCyWq/guZzEZ
BeRAt0X9OF+9fFWaPPw4DQqr+Mul7sJYIOPfV4NyzTKwD2lbdGso9Mb04cM/nsXO
xbJyh1yP5PC8d3zGXuDIUVdQEu7nK/4XP+dW8Nas3Dbxqp5VrjgtCv0zamys4G4z
cL8q2Rk0Zswa/KD8++s06BRQODLNEHctxPyfi+NcG/uRdRq4CnvJtYx/kpw+rXDo
ZHgybh51P8kNDohYfkSTSG4V32uqFpqyk7RnHKdeOJzGErTWzodE24Igl/7G7fXa
iI5UMu0RYup0sauBTTDnyuSwaVS/nD2XX3yw5XzttAHjDbMYIF4wVEdegit/aGkh
BHqcuZtdYw/grD/IRDUUqMP2xJd4L2lzhBhs9Jcx8Y8eslQG4MlzGRk43QrPUmEw
9kqH3iu3v7MF2asTT6+Dck84nbRqFQ4Fa9M9nnXZZGM1ETykdeStbtjBbl3WJK/d
zrv5xhNll+HClakqjgwU8uvzat7OqZ+Is7ClIMnG65JGJe+ioOTqxiUQxfjctxjA
CoZLVv6kKG5O/McMubE0xl/EG7pWFMwyWHx/LM2CNaZuHhru1e1i3D/Q+vbtN9cm
o70FUbtPmMfLbScOqCUDuTPkzDI3ANhRVcwgZ49VKJXctVidXstCsglZcLtJLd62
ghuAhqUZu9kHQ2My8aGqzYsOBopvOxikC/+NByChAPjheho8iGth6rJGdpqjCQq9
v0kelZ+zghoFPq8uorS7bT86fWhEvLMkQ4qaIskk0XUxImWC/Sq6fK/N2/LoukNW
pVsmJ4NhojB4Qql2yw5T7ufajSBX9p41TlqH9u7l0L5zJa6kpz1yai95eyWqiG+r
rj9HQuo1WK6mwABSkC30tfUTb4fbzGktvwbKG2wiktnkFH9q0Avu1YWlizWwlm89
9AsPPfJYL65WEd0bVudFT8m2iYfBsRZgnaKQ53mJ8CXw7NyxiDvqaag7jJ/N7NvB
OEtCzSkr0i/HIVuzJ1vLZwHlHnUbFEO4B5wZoyQ/SEXsCGCTHJUealUDi0y4kR1A
4l5LZSUN9tBh9skaLOnYPA64GHaeb2V80qpGK297O7noMkFpKmtyfc5ZUwmpQqt9
IZX8dz0LVpxCcumPixT5x4DU/ykJbxUSxn18PS7eP+Wl4Y95NsWQ+m9XQwinToVn
mlU9xIfqoaB+liEFvoXaqoOBxX1FgJJjfr7wF47kw7r/xB3+bxxE58+nh24u2dd7
aNZWirV75GgRHSlml/La/EnsVzNq+5Vy0Ju9CXNprLn+z4BQGxN9TBm8cFwAf9Pe
bhB8Of2hcOKiAGuw3ze7XpBfn71/l9uEWOqpvhPfIt5+8fA5k0a9KgxHkq0xvz/L
flu+a/BzDJ61sHrwSK9jfeNfyS/FNQYOAXqHyen8JXwNgNHjEuoNMwd0oX1wuERq
xo+En6KIGsUrf94mY7JcLxVnnmZjcVJ/73Jqe6b/Nrs/6JtGhhVAnCFNWdoFug4L
UXzlgsx1qbqZZPvyRlgmHxhcaLi7womOeQXyuhflY9abl/6Nod4J7JK7kMYhxErr
hP2na5ePOmMBPYMfz+I3t8RG5vfT1hDYwgJowrZIxoAYll4ziFU8wvH9Ps7qeiBZ
YaNDSc2mYQB9Chz98kEvaz0/A7zu22czlpnJaVf+prU2Jx7DhGlz5hWnraa9iWib
H+hAN7o0qwH/loThuCdlpqbsjwDWxzqa9MIDd+/+YFnMzZzInz310jFOihabY2ms
AvfN9P4cemj66DOB8h5vVGk3SKX/Y1ZPS4o7aV5bW3WtfmCOFzRhmKN1e0BbqU97
KiUk2qIrBF37kfudWJ8FHDqMgcthoxD7zO4B7rvzQO3Rnvp7l9gqv7R3xi0bNvz5
N98akXGN6BcwTgt4U7MG2PzU6ZrQ+4GMuWGVMUTRHOnv1dNfxtXFWZc6WPhnvV4u
3A46ggXXl99xZ6pgIH14vn0fFhlJlXxkk5p5wEWhbsZh+MSb2aBDuXudoL7QCiID
ibKjGpEiuhhuxU5SNAsuCA/ooQUtviZFx9ZU4GZSdC3bL8wHJUcl+dLbjBK4rfoJ
bhMogU+4YIL5PBNMxGb3PQ9036y6PdPQpTLcpU1DC1N87cPoRMj3xUQhI56XtL41
EPpiKowvtBuoTyfUGVEXbcTJC0xpc6JjKfzwHk51Qt5pgaAPpLk6GH09TOCdZXep
NCQYpX+PydlhqjQx8UyGJc0VX331WI12d3qCXF+hsAoSMzJkd7ruPXsLjFNQKo9F
cZkaH6199bJy5P9SoxRCU4KdGwneEv22gU2ShQrJlmr09P762eWplyjaB+fdGsMh
4lq+6sNprEnJLjfZqm/AWFkJTNYClc8EkPmeyPRlWA4nPR8XGPqKZ2pRLAGVBqUm
ZwBoxia5jxEk1cKHRA7jYy5jHxH/p1eIt3LHVN5tj2FFTY4kR1GvnxopHYl+4oes
RTjlPagtC+13zzDPrCdmmYqAOPFIXso/bZX3+HMJugWe6f16iJDimB+heDYXpaS/
4Q4PNxLHXz8LGdUYeu78OChcCwiAyID/b1EaoMhgAZdmQs20WaLMlTzqqoKbtjGu
ROoxfFvg0A6TTefvcUZL88P12Or/nnvhMNR3vIlhVZTGwNztwOaMD/9xq/B9RpwJ
q7KEWQSbGjkkKRWgCiDmtcUQvoqcywORLGCRpn7Q5IRYPEnNGbnvgEUzpVt2NDII
5rvqwMEXRrUkJWzkNQnSv5ic8R6nDSJyLRAyFtY9m0tpELP7zrU0bCAEHbHy5tGr
E1kXLhLeflsYX18Ff5utJ+g5JuGm31mVHB4MnII/1dxmooVkuqgneBarIDYvh8JS
jcQ1wa5eVkok9T5jDTdeqqEjXUUFHTTe15+m+uydjKfN82+dcAmOvqgHWb/eTPpA
h7QhKgIMAIA/8rWaUSbeMEQ5Z9D6LpWZ/lqWDlb5ilQXi8pKTz+Iev5DwwrRbbxQ
HDZqT4fN5Nj+fLvtk/lLs1L9lzYfrqdWKi2VkGZDs4wWf8JpfZEWp2YD+Q6odSSz
yic5X6oDakWiDw6ARF7ZoZdHqyUAU8I1V6GdNzmOMVwsFbjyOrjzI1E6gw38oCCH
JRehYCeIxHsEoWmkBJ3reoW27Ik/d2a+Mq/VY/d42tNSyxTN4oMk6RRdlV1H8cIl
LWf7f7Tz+OcCOy7Ok52NyiwlE0cetWGDDtjgv+pdpODdhuxhkZV4KA2771k+FOHc
VBlZLIdN00K8f9QCQQtCOqupSDdhysEnWJL+cfongkRp75HQY7XzIPJouBN+GI67
uNliER3ywY++4nZXAKkc6mklFoBYi9CIlQ7QavX32laP2dHamyvpj3lEMj1An1dK
yFCqKi15OGJbuxezzDuK2S1iPo40JjTeGP6qwkHYZ490+8HAGj8yrfK0v5lqdKRM
zFw8ajAvzWQgaebd227QW1lRhrQ/Rgsg+BzIL3qcxcgLTKW5LD7JlQL27Ef5OdbU
y3SibKYqGMp3LJJVRkcAXG3pYZqPxQ/dnxCZ4SDMMtvLpdd49oC6uEZP5Mx5oNJK
Ov1QxLVYx+3kffcR0r9Wby28dJitBQxZmR3TurPiOFAsPqekeAGtQy5pgXJR9tbD
Ufqlp49kUMU1y9tD2JUH3PoQkRruq44QlEa1708zNe3s/zHiMC7hTmZrh0Fy/o+0
mCOpjSU63ckR5JXEt+L7lqeevlgisF9v/F7R0pBfaUqBnBbqsc97o0kaanVzRJte
DgVWKjAAJKxdpGDpbJXCD8zIHV3wM1se8+zuxQ0+2zPi6uoz5BH53M8/W7tNTT/K
6foQZtviJsjnN+47TLjzADvGj0riuJYAonqSlDU38L9etOUtGBv2hcJ0nzEzQOIS
+pHkZ/0uOEzns4QiOPeVCFW7vUA/bc7zlC+KIFBzfZdpYNTifZCRlJ4GI76WCYxU
7H50AMvJW6eczutuihsZglVgYplhBnxla111SwBrdRJBv/wffdvUbocDKft7+mqu
1NVjo1nMgrS52nUSFHbYIH4WJna+6uoBmipRhUsjvrqljCeB8G54bCy5lPiQexyg
vL4k5JvR7EtTjrAANmLCEiuJL0rz7gv2NFMFiLgU3gaBSppkSr0fqCOlFyQtO1ss
Jkb7l9tEkr3EcEPtJyOtOkVZpFN3/ocapPiuojb2Myf3NN/lT71OKwPOFxtZGhvz
Rg4cjYY/hhLusTw5Q11ie5c7YpzZhgKLIuW5rRSI79ESofRthQPl6SjkrIoNYt88
DsVMFMyxBjs3TACetZXGSpKDCXFuPlXqGYr8KRQHKw6hj0Qeq80P7k9614mOW18y
6eyAgr8JB9v0RebaC/OOYGPapM01aJygb85GId7MiO1OXRdIRhlB89O1RZjW5A9e
BSCT4alUiGr/R9kktdZ4HxMWc0VcsxGWm50VObZG0/mAf4CxqD5iLP5QDps7wFFX
tf0NeVK/odtY4iBc5sdaye2PlpSIx/bz5IiZuoNtNcduJATZMfhIwo+LJ/R302k5
EZuusxI4tH2pmhVgckBSWFApuoVuNkt6UcMWGzmmyhc5fOsXhVu/eQ35iHzlJRmM
bMzRBGuq4TpgTFFa+oN3DCquRG6OPWu4fsuxDgcG8EdtOxFP96aqYcr1Pv3ZBRm3
Bo4l1xy6E8X5rucwtopy/wU4qjof8QOUVx4o0se7xKQ2+G54wCoSQQyIsWPyq49j
Yx1WlaXxVlrSVp4SPwIjJqb5M8CBiZV3Y3ZDGnZTLG6y5jtuv+W/2AkJ5VPnmpDS
6I+vU/7SMlQ6F9lXBfrz81cbBqqkG0MRJ5X8Q3LYEG9Sn92fjs+dL3PDYV3TMBuT
EFx2j/QgjAO9dRdtqp3Dud5tKw4cTYox927YIJKO92d85LbPDOqxxb/q16NzTAul
oUH1m8sTVNdAX1qsmdVVGOgB4/kp9RC4n+IctHAE3No6tl7lWmcnzn0JZRfOpMJR
eLZtd1CB9vqjS1ozRL45RMmIZmhfDWgwFQxE35Rob8UFw9jWahZvbbRdG8D9q3Z/
zVfFAh62FssczOn/jbTjQ6C7RbsheaXmkYEBQHA7vmsUnZ/MtlJ4Y1Ka5r6Y5/bv
QREcEyXwW8RB9m4QXHVtv0sAd94xB649t0ai0Ol8Mz1pmG3REUtGA4udCtVfDfZc
9Yhg5Ti5xb5brHtHPo49QnWuE6p+9b5Qy4JJ55ziy1ok6tp0ab+xwc8Hr8HtBp+H
r0Bu/1VbYoOCR9oSbLBgpWlB9MpVBz70Ra35KxS4IJ5vrSCjePzjta5kwOGmm6MN
ZzLDCKrFRw0XX5Ly9X7pN2VlPLL5Ma40JR3EiTSdUJv71yZ7/K1qmpfLTpPLp9h3
SO/DLYmiQ34qQr/nI6YVKNAIL1s+T19tb7BH9FonmWBSie9lilB6tQgNPzV9JUrg
j3c4jYImNuaxs5CrNgGLi/que5HppIX9SHo5fry3p5+d7uA7gzQhq04E9lHCLLr1
YV+xKRq9AHgVBeIsmkR7m7RbxqH7GOeOaSrzN1oifGlh2v0dCoEQszrUK0muQ3LB
JvrfSvfJW8chsf6hFV/f1Zp5UmsmkKIWCbUzy1VyaBtZxAP77RXaKn8gy2TAkbR5
tixjN3PG+mEK6Okj1leyZbUVRfvvsUZJpMiKTpLKG/Stgmds1WsmfNzU7rEUdoUI
seLZ24D9kAfzob86oukYVieVTf4WJFDCVX49aTP6WpWNDBGGpWJI+sekx4+xddpt
2Kd3MT2X+Sr32mmIBB6M1ikm3doZQtiwYu0gnbcXLc5p2XWNEbbC6ETOmOiT7s2M
lLMM0zALlwVzURLn/vKpi8nwbQqO50M83qiJuKEbVTxzZRMA9etCatx4qslmgmNq
zfqaB7rxaEwUXDobSS3z8MhS2w4/b4Yf9pJYe9oVXpIqn9IbNnSEroxPePQ3T/sp
hn8hYMKmhiImAPnqoVBaZZ7UitFHnFX8tTSWfL/0k33PjBnJ7yg24NL+5jAkx/nk
WeamqD78f4NkuljhmZQuDJv9tvQ8dJKqis/6QADljkbdy96T2bB5kX2rBsnNOXa9
W1Wsm4xIvU9nNNwE0SHdpO+3px4tWFSY97mRKcPHgx4145CH9us1zjI7o1coMU8D
9XuysoJCte2qMDhvrZCAldpnjCbyX7Cz34Dvo+fjevtKXjOZcTkF7cO5dWCMCOLE
YFTdbQ8i6HzlIk334U2tk2Fe8v9NRrEGDVF8jUvplzq9BZxmbI+lpIbMjBGzs6oc
4yqDPsWQUxqhQz1YrJJ6Ewfgb049nvVyvdaWXP9RgWPgdpQLUwCajEsvr6/5G0fr
DEeMN5Rlsn6RbyrgNPt+WokN1709nze3c2VTSx08rxHu4LOZnnISFuGo0ua4caRx
tYa0sEW9K6qJEEpit3SgwSGj8/TuxnulVx/SOif0/3AXJvJyWunYzEKxQ3FPDSWV
c2mwnilzPHYVHSpOjRqc6tNwM3YlELkc0R77i2jCjNXuTpya+IKf+QhZGkN2NBCL
OBFI1dGxQ122uaf9Jdt8UOxQh8GM5GImnNYM0cSDbZHk0pCUVDHxuCwQGh/aLESw
m/sImKmFIUEcSZBSZFPgvwmkJFq+/VJBloakfetefiV+gGFYkvZTF18qkm5OKdKS
/SZQaw1m9pbYQxR6HN6H9u8nLnhiqJ4XldjNhKBvNUMkqiGYvDeUYbSVZV4pb/Ye
jhFLSHQqbFzsbccSO0p7XKGu+vq7D4fZVmA4VUIR2PzY/rWlMW0Z4VnRpUwiRSo2
AKbVplYlNtTz0UxSNK1YcQ0fhxgqWs0qkV3BADDVoYB47xwdizG1VHY8IEJbrHQO
2NREZ9cc1aF7j/J/xMvxvul69SsTWJngW0D/Tq0YCnq2XADowADRJXycxQaTT90R
Pnm9RaUvOgr9cb/mcfhsN2xqpxWL9mV5UdaAr/alCg907Sg9u/1rWXjfnX9J1X9w
7TaxSOwv3PeHyT6ggwafpbQJ40ZjyUQl1a+JvxTOPO54JpcIKUNzYYULmtebNky7
7bjpIb7f1QSf24sxYUyOIawyyK5VFkr9ulTW4vAkAijob4CZFAZvVOV5N1lMkjSn
b9Lcz7bieCIzPflKmcsKli+UhZ8aQ7spUN3spP0ivDYu1oCFT4GWcHpIKaF5a3lK
HrvYN9cqcvongdgcPyEzcDQQa5H4zF16Td6fzRYMTjYrSiRw10pXrZCj8M9MM8YK
gQ1wOdWUrmG9H3Jfg54B0FQxpYt6bhwDVPPdZsVK2zV/dV5411x4Cxu3ls5O/w1f
bJZ+pTdU2RERgBrVMI629ucXZmrw8IaRui99+IVb8ilZYi+H/XJ0NOexTRczyNzn
VoLbuKQiqKV93QoK7Nz7eXVCHQUPvvwv0B+x3bNUNAvQ3ee5NU7kzsYiTtLAte4M
KIh903hrv/E94DRA1aEMlUNseFEVablodBWlZ5jBGgrrKzr2NicH1CqiKY0I9lEL
u+SBqTGvPgKCv1EzF64uG3bRN2nY3R+FyRpKqtshOKGmpIZh1WIK/HQmEW6hcnjG
Nkf3sab9+GK42b+46WC7xVMksyaWpZiqMFiTMud/w8Z6rEX79VzhqUZ9YVT425nw
Rd03r7OdxOpDWCJQrS8Iab4ny1t4y4TsWr0nSKNIAT6B0ZmMEXaqLDl+F05o1OBK
x+VC90Vhu2IyVkhNLBSeQwdUMvQctlZfL6vLh0oouxrBVj+SwlSGQcrCopz8jwq3
cgp5YRzJGLbId/R2vJZi6jNAsk1U+qi+AmUbcRUhZ841PlJlvBLeJONwxsDHCJLL
QJd7ILJ8vJW+FGdLikdJi37WDYI+1R2T4LDe3kbvhQb6w+h/WQpD1fvIbrUwHKAh
qjfzAxKQLLA3f+syZdD6WJpC1OepUhXOGbpqVC0kN6AUoDNHMLWgzs4fcsg4QFfJ
qP+yWkVtCGdp9JYr5GtbbeCGHZc3bMLSEZebWtQ7g8VQ/8c6YXkO3UziSnfW/sxH
ScTK2RzEj8lFV9v39M68hcTAszsUu42DUofPw6TVEWZjURzKJQFgFbEn5bP1qt/5
8KbHAxvZyzMXt5o80SrL0YkdUB3l7qcowAG5zmKt19gGIlTh195FYODN5q/F25ld
71MHGZX5BasAAhKUiq0AgPlNBAD3KXXY9s3sCVVXFEUSXsOhBEUC0HNYYn/p/X0D
GQR76PBbuumUiRPe9cMQjaiyunOrm5HCQc0QI64nXbIjrDP+fIFJjuYqIYcTXOkR
XRoqub8MF9K1/3CgoWtOM/XVIZXkECfxao3wdwZB+N9q3IlVDJ+6+kFAD7pL1Hez
kA57YMO7VOPsTCIPZyQhNN/kBhgYNXz1sfYFVbtTw8tnaMa7gVaqtgg4lzP6hoq4
xxuNF8V6A9J10uZ84Qk5aIHcGNgHv7axHTYRf4qhm05EvzkbmUB5hicycJZvcSD2
43w2fDfcxQQHvY5KOemVMGUnossVygyhN9NyEEUbgI65/Hkg2JO3l005PumKxKpK
2Y70GT7zEDl3eG2YKT0h34NTpVJmJLq+oHTY63L+ADpcbvH+hOKavP+cUzIxIGLK
KlnD6Wc6W11KVRngeO03fzt/iOkDenCdIPs/Vm/Zmh1xO6jR53iYXv+jLqhbGLwu
sUvjPGh3RvbaPlBpeidmqCs3NW884zX/O0S1igMejg6SQDyV3fEpwzmn+vgMVKd+
Z2rYn8Q9JrO82WaZFeN9kIiKdkoKN2z1m2abW+op5SJIFYt8ac4Nr3I6YABsjrNI
yqGKS/Er3cukBENqiSb0Cj8nhoSr94QGjbKkx5GpqPCcMgDcn1cFTvkS/a9y4iIx
jiIcwkOtL8bwgDIv64BMGhTuTJS7mrvNRL1BwmZ0TYAjItpriEhOwI/bzqpmHy11
UbeX4OSkFpdUxCBx8olRYrodOi9JtwogB9J26SPguW34g0PTtHUH4Pka3LfLKbnN
d9+zBLLbnxYxRv1qk/3lxa1t89uH/8zA6B7amRO48z+apHysSBdlY207lux6cPdQ
MVJe2FJxkclH0XR+ZXyzZbtGKWI2I0ICcchRDGuVHPitFUlsxJGg5upvmwoNGZAX
4RtwuqJ6Mh3IkT7goxOQ/Ndyg/J/y0QuRzJ0ueo6CeWShb520Lft8T8JuP/+/IgT
JUqwHEFXsG4aeW9K1BTQWvBubz4Rf6xd5i+uG8wIdGOxSsqGuqwfGN59ib9ciWCa
WK0zM4FlqWWkaA1j3NikHxVmgVKOihGu3VrEPUWtJzYoQSElHFF2QmyuByZqBDx+
UtbJ2ZQSIMl5OfR5u9u8RcoMiKXN+rMDPViuuHagq9Gi1529LypjulISmn7x1YOU
R8HkoGkcpzTrmy0YE1G6csWJHT2qAIpYNzaSWDiZkkyi9FGO3yrS74omkvTnld39
XpLLKGOm/lQ0WmqECRBf//67YNluFDYtEqRJaN7HF8M7mU1jbWpl8/w96f5/KZBz
MXgF5TeO4wwn3tOEyoq8SuZvj+55FsaYzyJWXCfgxMJDNO29xKreg7LKRTjQ1hdM
Tv5tbBcy1tLAEnCGnjy537Ex0x4JM367V7VyD0U8ovyFmQ33jtAg2LyG7D8/fFAh
Ojvsn0SGbUsjpiREwi2Kz/EDCgO7iWtOyU9Na70p015oMK+bIbpoWXAJ4bMLQbhC
wAv9E99FLagjw3MVANB0fnCms5w+TZEhXdG5AsDvFru3R5mnGB7MDi/Fmpz/vT6V
dWIFrZ0CL2m2d0Qioo6c5pp13RZa3njnfSWflFi4BB2maLdt5B5cfR+Uj+Rb+ajv
1unEXdDjc22KD/PMKJ0dCg4aD9mK+WMV4usurubqWKnMb8YATT8bL/zA8PLMapAO
c1h2VLufU/9f1XL/IjvNOmfQf7elzkLe4Wx25rwTMssbFINiCLaQp+NsPczDB43r
6FS6SY1TTgTICWk2yFe3CSuEL1J73t9TDFfAWtYDUgLShs4rPwqJbQLKpuDwGlIq
jznwSV3AksxPB+ly7EB30y7AYCzSZitVbi/wjbTIPnoG9bzGem5Vdx4D6jTVOk/o
mRfNr4UnNl8pekI2BzJdVBconoeI+O/9/fwp0rth2OgsAWgJlCAlT07ul7V0E5vL
NN2eX/5xuY5XUL/ZgYEcOkX0oCT1a/zHaHa9qeMgm4/+SPJWvULHJa+28gbf4dnd
UB14wsIzeaub9rU/CYRv5/42W3MzrooJB0i2FaW4J7rjA6hZK2o9r9SMsgbvZEXS
LzDszo2/7s5IDMjMUyKbwDHYAzytQ0G7mJXPTDrmHTu5/kBDV+ecV4NIkNTp6nwX
Uy5E/CCETbqckZcbx/DbxdEM8HxlWzjwKQfiw8uprrvXKCkfw+VuQcsFXNYaMmcf
qWbz+rl44T7sqeUccKgyhHsw9G79cztQG9pgp2kDRagy1c3AEdr/PmnXSOM2simW
o6Fmgnar0rrSxrQLfQEnjR002cKgzsv3W0fH/O9syk8AYDj7B48Ef/qieokH9M7J
mhFG/iCLVhjEWxVa+tKHHMh14fPw1Ush3PautVxrMqpWfweLJclIKltDqK02cSVa
Qr94sHqppdcxeaRy78mQR8XeH9RFvMEmmz+SpmZBy2ZBdkjBd5ySHmGMdLdmW2gi
VLum5k+TB7lr/tgrCsNOXtmufEcNsMEPCdaJBphxGeiUlvUtAkLZBaWJnUN5GLag
qVG74wSG7lL3dnZuVd9lgzRQQJjHY1+JR/+Q2yP+tfOkP/pwVU0zmkT6krBf0idt
NIRBJgyV6SFPLFVm/XvGfhziSxOx4aEKrlwmQUVkQkqDNfnudaX4HO7jgNT30lMF
FW5xCE1X8z11B+KOY6CCc8F3VpZ5kujihuwB22Z1d8WLdbMtTevl1v3lLxOpyHXd
5ssxTWXeqIVjb8HvnUH5OUAvuwqWsXLGDcosKpMACmLjCpFpCJGFhuPP976P3BtG
6WLonXdTJ9JCcdMXYuEF1fE/uGj/zo3wrnpaGE427aC43fhCepVPtBcmajiBTrHw
U15bd6aV4dSXD4UQxTr7gZZaXboX+9HzTAlUyMTcf92LOrAh2wMC++gDXdLkWZ0T
GeLPCHkzBqcsQch24Zhb5grc3jyF2Bj8NpeiG0tsmkIjZPpv5T5pfzjlbWJ0f24M
pJ3BcqcPHwCBT+q5rI51walbrrSufwBcqah4a+XxF9k9nWJP1GbKFrtiK5XyIWwN
1/Hjvin8lec38T+ZRL1Ds+1N37aWeMVLJZZnZ1pWRjuNaGbj21werwzrgkM70xCV
b3vrxnb3F6h6RkplOhOzh8AUEGGhQ6GZhr+0LU76qFiD1oCSiQpScJYv7lQD29Ff
/dhyv1B9Cjrb4SphDogUo+b+z1atGFVAJHRuumBMvbciT/vWXwD6Oh/7NyjLASL+
1dqT583cH/4TxS8rKawk9V9LZIG/Nq0JKkHVi8LtzEKFiocOZYUfPsYCay0sMmcA
RAyVFcpv5S+5U93FgFnfOwfHPLXhbpxRwSo7NUOWKPOrTJ/n8zxowZ08+8fmp0uU
la36BMmU6F3zWvmcd/jK4pslbZSxYbkjewpy9GQIVB6yfhYjK2xlTmyeQkosMJnJ
Cv50SJg/gfZHYEMO8J+U7AqWzBzGBbi9n8IGxxpk6vE3wFs+2d3wctS8c8DEm6DZ
vucCNsfgcJ6XV5rGMSY0w/PEn6h1AoqSKRYgaR2vWsrlhl2oLiQEXU57il/woHrL
FqR7R6KloMRXqi/aA3p8UfrDzEJOGdAj0GXuTvZ6E9mnlDEup9ctpVQFGg4topHK
4KnUiA5jcGxDw2//49WCPwrgb1nlmd5YbWqLcGItcvdgZTDZ6MxFvaBwiRdzTm0X
wVXNS6Z9JPdXsS7H+VxF62UFt15Qlkn4/6ps+2/8ofMRzTYmyk9J3Dj4cL9dVi09
Ug4s7ZLuzogR2R/MjqlPn1JiTpUL3apISjK3uhuTmPh7OoSV2A1yr7MjputnmLST
q4A4lf7aRj36crxfHNbMN1q+8EMKsdqHaokqZpOCkWXwT7VaZApoMdp66P5rfVlw
Ago+oMarYWC24hpP03u0SuFEQKmlfAoDmKWEy7sspYZ3D2QZ/sS4MdDwm12NgkGD
J8jtmkvXvQrHkUxkPrQSfDIrJ9dNuIdICLay5k+oKCciuB5FpnqNyJsxKEkXdqDM
7DCHJSrHH+nBwfoLcqThVceQOpM/aynyiC7nqFcagL+2HpkFplrrhiC5E8QD7a1I
VNDBCtcg7KFsHT3/2mLyuzBdql9n92JgIJA7jKksNN+59D0Mvm8BjnrKAZpMCbRk
eSK72PhYh/2lfUCgLCTuzUEit9ih8pvHZGZYT3KG6qHOVAaP2RU0er6RT7gbNvBA
zFW/KOTWwNkNYN/6hpDliT8iIsc/w4J86EKcbAhhfi15e0FyvzswcT5EnCNL00Nx
Vb/NtHtp+i9d0AHE1Y9UnLWG0zcBmuyhVc9BP9nzrytfJuSuIwvGodZVvP9gUNfa
6bG7QU4LNSA1dbdw/B98Knevu4347Ei6ZbmQHx+KXY1oGW8fBsJ4gRwVny4bqAly
19xv1IV1y+jDLjxRqedQwDLUIsoQP4o2H0PYx++9QD9EQ/7b2smB3XckzoVWmlmq
86EfQFI69CWbozyXvnsLzCg86jWtZ+w89tJOTruvlC/azSWcReg9LAmsCqILCxEf
tEH1YhhXXm59MoVT8cgVWIgKv66A2mZHXt7MAVay83O8wBhOvs7jFuibMeVYobK1
rs55/Zd5bUo/Lc9mrbWOf0HcnFPNXYBmfYLaZ8e1esZ7ncuC+HGp2e/NMvwKIxx0
SCm0FdGVVriXjAYh4k7FyGbIXGPxAUS4Qi0cg/py1EokghD6yLHAOFUbHa/FXcfE
WJ/k5VH7cUz32L7QE+RAmO4CcsjH4ftQ8yzaVsMH6IdiDIPK+5yFkb/jNALTghfZ
OoHom1DhYjLAbKN5CYyOLVoaLkLJP+YezvQ0m1XcSiRhKgVJjueEyo6wenlZCqjR
URIldtEbBmT8ACjpi3Qn7a/QiWvRGPTtqWjlFLUHHI9Z4IytRfSWq14fTvKbDyer
/GuWzwLN2hkQCzAzCe7wFp7amYVmpg4qHmOGrw/k0MuuLK3bhWjrv6uR1q9nqE4A
HwYv5uBWwGIO5YRFfSw5FdFjQBtUfaOPMMMu9+ZI/qivYn0gH+Sx08sbdTstUUs6
wbzn2bWMcH1d1/bBKxfrBf1I/TmdhVfttu7n4itPzeryOO+lxJ10pZ5NRUX3MY+O
UKBtLDuzg4E/q5HgKfkknwkQvFhPpbSkFLecGvrVNqOavhmTEzyF3zmXi3HeNtji
juRdUnZtivPASc8EzrTGeo0PoG7uk2o0+4Gt8Bu/9iYs/Q1AN4lUUR6cl0Rk3ZVr
kigaeG0WuJ8reqCUxFUE9o29qpCDi7ExqC2YspdsI3sk2ajvPf+KZv3G8i23TkNT
s0QbjU3yHrNRoTeotA2TMHiCF1uobbZbQwhnP9FlRTpQuNAm4xveo31XM/fR52s2
iH+UiYDlHl+VYOwnGKKEquUBm7KJFEdMoGyyjlkUAjW3i8Hpfh2F/rXKpWxIgeaF
lZedin8QG2YMCC4TTPA8MkST8EelB41rbyerBSHZbI1XxksXmxuOA/lmoxrdX0IY
dSUjeEMoQZEA6a2ZPrVHMJ3o7A3RHISSvEAp1MIgCWh1wvfgnp17ucEeSXoB+1gT
fXGiP1dA3K4Rbjj1QRdftRqQT/WpMag/JbKc9zrPDmviqHjuPU2bo/UWEsfSC17A
nGkKG+QQreN2QdB0C5CW9nrV71tNJcU7I2bipsZCNKrH+DNihBt9o+KqQNCXyTmn
N5PeqKVCgGKffNZpITBrsNXO3wV8v6WkPHPwBhDkavVTeVK2BiBaoWJvuwN0sp7g
HHvGe7W2jk9vJNIK6UB0LSo1tFqOFXGAaU51IEGWL7kX+95Jxzij+kr9ScsLVS0z
Ey0YuVRcPPnmxHYGhIlNUwJP8hxjwkTR7WXx0Xld1UuLs8vqurZXE1zCh0ywRGue
LFFheqTzTNWXIJC89OSxOLRf/gtcrI/PWyGiAzrQnsBYUa0MJC40qel2YBrsox84
0oNkZ0zciyNvgC0wLFV0uZ64ueLq1mt2Hs8YnlQZJvpqjIE1uYijjL2gFGVeoksd
dtEbtKDTt+cV5/w1oSpP9E/14mTJW6diz1Parzf4hGMmIdE77mWaQSS/bHzYL6U8
FTjVqEUlDXGhXyCLiVRy/ikQu+A2lwnJ5huCCuoS4B5MvbcUKCc2OZDIQssKJt7w
j3yPfMybO40a+234xkVSU0l8JjmLO5GK9NSwvwakgJlXWpZ6ghK0VcNlo7aVWF72
SBs+Y3cSNNc8nXfZVPeR58rbQRhKReRPBFQS/8VR1V/rgE5cQzY51h/o0x/cs9Ul
fKRblZHWcUlmGNaV1pxC1lQNuFakMydAcGF4fIW4YoonQ11qj6m7MjqMxIzk7N/l
YdULKH3rkrRtLp6KWaG4QhamYsvSiPvrmq9xOxZepZinmjCJeSU97ir38TkfoO+H
H3DUxhz+B2wbs7UCKrgNaOR1qdi8LrAqSuj+PZFhrHU3wfS5+/tf8J3HGk4FXwwj
eviZ/BFRk6z6PpVLti0sTkXz4ZGhKBffzxNOTegJ70flTk7H9Eryc2H7ZE4GszGt
OcoZTVpyBHX28zv2tNHg9Bpsdu2N8bSzjLQ4+0QQfdi7AJDQ7deLc/+UaWw7TlIO
QCyMV6cELNTWaw+02Nenh3UVsTl9f2UyRo4gBpb5q46PArE4ZZBg09/yAU+u+ZBZ
oxIh0Hmm5waSjWgzl8MTkOlpZZJmjvh0DLKnY7pIjFgsAjGp9gs0Txb9LGziwVyt
qcrbrDJqAd+S1lynIYCZsxHKy+WPX4gO16BNdEYakTe9T6XpyURc/S8x7Bc5usnt
zT6NdhcxqnljjGi9Cc4GWAERY8qJEY8RxJ/zor6AX/JPKT02vewImCysN2OAkxjF
Os03/+HJvvwwnFQM8W2hPmjYOQLW/TB4jCL38midM2SnrMxP7GjPk0wzxKQ1uuuV
Dbtnop8D6GSfIOuogR7bKnPxZ3xWjq3mmeS71eiA/4z27NxdJ9gSK6fDOfZXTFKq
y2xUG4st7Hx38lCnUOHFNO9INxkLqdoqlQj+8LEkprd1M2wyM8v/Kuauu3tJ2LnA
ga4AxlDWbse5LoTMSlFmGFgfkxRbvYDxRj+OH2b2YKqqvTzWFGmuSFOmXmj1XKvm
XykE77PW6MkvFRzQSVfoGk2KDv62tm72+uHb12ZR/lrJWCO15jo6TuaSpHld8jBY
e/5ilO3PDCCY/E67VMN1AoQ/V29TRw+wwCYmCm14VQthAo1Xd1z4m4kXG72uVF+B
ORJTbYWgkLvP13HIAYouswMu35FlmwbuCbhAZXgp+Qi/6vHphyEsbyxJzywzgGWm
GGVPpRqqQ2Gkv51c1r28K2LhlAklsl1Flw7qzb6eYod9J33D4+BtAQd1yyrGJEQQ
W6rKTEkSWF1jwGMStFSbJZ8Xu0TCQk2z7DdMXrKMu/VCtIpTLd7yduFnxYHmkCo8
wGE/Yre9eL5iyVxp2SvRrtNsPQ0UP9kzEpFoGBSQqdaFwhtugoOx4h1WJNBNhTaf
lo8XG3CFKzvGymgDHRMOq89fxEY1pRRNjyN9Nw49513smGMjg+RDecIssZPAdVcz
mKaYwpJRmrQAVkVYwn0uPy+wCI7JCLKie6S+VsCwbB7HYLpjIJjsIDuUb0+kc/Bu
bpekeTl3Cfsf6rIjJ1DIieuXu+mDiIdQYuZS0Fp9TSMsl1IKrY/VkWDbSyAzAJu3
bAHL7Di1IApavYDCdw5/eurOEkeljQk3O6LqdUGLeKqycgdwFN/20c/H1G99HOK+
hxGHuBbh/ovBERL1R5LslgUZk/f2tUQmPT4FCvp+WsWiMbPGCfKLd+yIS53WLXt1
/ifMPxAzmkASq/jKAZmWRJzpJncnH1n2pfj8AcrYL7jPSM/nzfoTgdA0mTDrarUN
OfBzQpzm+Nx7MsoGoGEwafko1Jr5vX7ovWk9zPDVqUU/y3TDhgqmki+zDeowkJeL
tviDtpiuR4JXGcOnYDPu8U+3e45E+b5SjJQZIRxVOeVf6NjYQrx9+I0t4Y8gbdXC
qZysO7qEU8AMVZ83ZA5rtxD5au95E2LyI2s6rnAZZ0GeAsViBqxcDP4lsb47G1h/
Z/3PWXzXjBltuhdIKOyhSKKypBNV1F/VSMx7lwtgJgJ9EIxVRrpM7bK0PktHuJLB
vqQtxKtj0i+g4Xhc0bPGRsHefEOqT7ejca5sg3wt0mXsp1dfuFHgDUXpRJVii7u8
b792Px9L3RZuFSwLpH6YUQqKFWjnMr50JbQxdTKXzQ8Fdj73pZCluHZ9yg4w+B71
1Sruq4t9i4YS1QxYJvXxT4BHlHbBiG4XSSVxMElBWtJTlPYDhq3rmq4+D6KPLKjv
FayhbnKfWLtPmZR0q+AoFZbL1YERN+POWsuj92xlBWPwIGqglhfhvbEuTnxKb848
4H3W7YefTZHYMIk1jZbJ3IpdA/gw8Hf1451nASqRnm+9flTSeWUR84QeBTq0/YY9
p5RPK5UMxcGi2eE/2aDGgCNCad4G6VFvWu2nyMN16wjY6ILaAuweMlTLyOrerpuf
6wlEnqHqdT2esxLDu7zBtUVWOncLCLp9D/GhkIlfCj+4ODNSgXIIt2HEbFQwuHgy
WD4qt4Q0nEb52OQQtaE7X5/o2axoCIjypBhGybcA7bZSxkdDqtyu/LIi9Y2dkbp3
PtlOP9/kzY7Gljg4j9V19mnmgYUHATSgrcTIrfDVMnUIY+dBJLhBrK4TXcwvZJB+
fJRaTJZDWAkLL6Qlqsb/Ik+INd7e8gQd/287px2rZF6vZPTJSOkuEJP9pZRMgHGh
NOZafFVhRp79LomSoXhZI7usvLmIQMQ60ko3yfM2nYH0oP0U3XPypv2ao4NTd6Na
lR7n5tn5O5i0dXCW4WoY8IHEG4Hyqx3DlDedIHYeoRDDIiBWkrc2hCd1pJFGJPXW
BBl57i/BV9zslscFL1JnZh6SWTkCc7S+Pf5DeJRG7d1DDbnoBHa79/0WT750vutX
BcWUlB1tZY/FdmBbdeQAE1uF5aQxFdd21OOkdRFUg0uI/odoSMhyGO6ZtlOSD5LD
2dcNSSP62jK9rBnkn0pbn6sGSPAdzeUAuxxI/skGQ+eJsOgg7YeNi1iuzN8IH48I
b/W0AgU7ESLNM9nNP/8IhtZg7jTsXywX94P2zzjN0yDY4jqEYH06edxf3sd+DRUL
WkkX4zOkYBcSNIR2Ec6UhCH7JiZSMYxu3DAEsP3wBBR6l9bnZ/atnUdrLdidrbBw
i1iCW3kddJlIa4xYWfTi6+Kk1xjHBn1afIWwTSdSww5SEbZKC2JFEumH1lAqIapa
ZcVqJXDNHejYTFE8o6grqPPZlRwII5EacGfpV56P7Tp6Z5RyOtdfpNr9wYLawghT
AyNrQuieTpYILZIHssPjYEViQUyE32NQWDwQ+0Oa1uHz29TLTup8hTyjUEQmyL71
3SmUXGMC5l2zYFKSslkFN9UGNojQx422zTvURWWDOMOGpK/sN2NOa56F0olTD6S0
fm3HZ/1mdeKleKm38c42mZ0gmkz43lxDBX9dlaVXSVFIT3mlzdqm7DFkCC4cBzRF
rkep006KlpNUFHpwvZifaFfNSBjt+bm5qvsleY/GI1h48mCBahhGcqFCrBR2xHpm
fvT8Gk58d9zv2KZ0c5t1p7OxEOFR0CP/ko11UlsuNdFUaFP5yK+Q90tKBtRQHTkt
B8HxPn3hTFRWTT6a/KDCk7HXCm2uZD5EOGZLOvxnh3IXP2cQmXxG+b1Dyq8Q+iHT
877xZkVcaAKCnn1pNoSgDYKfKCmLxLqDzMs2HgaRxutsiEaDHZhv52nc82qUaWko
MNLxQIeeX1KjpdMM+ecNaP8qDckiqiPakwlo2OQ6QC62QOCpmWn6TYn/CBYetzMj
GBPppV6wAxMjpWaV7yUalPA3p5WtrohBNkH9wvpk6zTadt7gEpWHsLJy6exaoatl
Q46rlf7OH8Z2iBX+0m8o6lYCMQNtmBuqBBTrxLfBgskqpqKTIDZjFQCDDqIMIg1h
zQuFSgbxzir4AzevsmiJ/uNEfwGEmm2gzzaMDUpMVpv24m4LCd5Z76+MUa/U+oQB
ai+UDcrZJTynS+EiZm3293Ys5eK65ZNlcWt7whzBNPshmCcwOQAPnAzVjNlDs5Qn
CSQahjdQGWRdhmxnkuPg5Xi+tr7+KZEIEObusnqPFZ/4GFbr0DqHjH/b1uc1g0+c
p4QTXEp0T9ascBoNv2FMMQeew38O2cS/OdFHPKikXrpc7/Z7ek1iKTQDfWvqX1ji
BKuKO+eG3mBlMlt2zIn9FHriPmItCPXJCUqxLcsDFJ3awQB/uc9znxF55hYnF989
KF/MhDxzOEIcW5MjrqiWi+Ridvzteski4tWpUX0hcwNUgt5KzWCbY00z6L2OzeUC
8qyLN/8aB7Y1hbpZQSkMeh70h5US2Acs+IBj9sox/JqZtVzrSsahm9LkYRG/DnfN
LVrKEOYM1wGxlQyjxY7dzBfwHG8H/OSyEQw6GCTtfpsJTEbYRGAsz/GQsh2N4jEX
CbDVeZZdC+83MfxRgTiQM8EOU32IgP8tb+E3O7CZh4NooYuScSTHiv3YGIfFHYL/
8PdRMibWIsKgIMym30oTU4QJDe/C+KJdLKZEFvEtLEA1HxtMMzjFaUb784y4Gxyv
G0qcBbaZocnlQSXmNxemzYUrNuYT31k94vKtzfKTORXCzXyAtCgacF69QEEFAvMF
FeBYirD37Gz2DYSbBZ2mGy5zMykcRYf7vpmtH2WX1ncL4CvSYoOxqSlNEC0ExYtB
i6vhkIVnScl353eSdZbf6ka0R4Wn0sGYf/kvTDmTJjalQxN85dosEKgU3p7sfPTV
imsOfiiorTL8aFJvPt2Qwpt6aYe99cJvVhG6qo0CWig5rdcWYm+LqGAqnYkTs6oG
TFYD+KwYCgqn4qSKWWXWLtrmQ39jblvdzRB7HFfzl/1CQu8cQcte697kkEaTZub8
MhSuRs91BjKFhRyB+4vvc8r0Qv6y1DJWZj3jqXbGnkv8hMy3N5PXZic52j6Na3Jo
D9Ox/BfAZlOuW+b/yiRM5JNqc4VOCIrWUaE8iKdVwtNGtP82H6YwKgU+c7XYk07a
KGXA9ZmGcDEWHExXGT3ugzOqgt1XQHk/Obs2MRNDl2IDW2mIM2ZH3IfGtglJgo9Z
qvsI0zDV+7YsUKQmgRZrlAdwT0wiMKo1/U8xbSb5C6i6kwARU2vlgprcK7wHLcNX
vmwfAzIG0ACr00cd4ZTJhJe3IlOKuM7Rqh0tRXxA+p/yNpeoEFjguIo64YmOJDPf
h0fe2T2U0TnE0dOMTeOVyuxBd4/FTZ7y0XEVY4FXV6pQu655L03Oh7gJkybVhT9U
jSWGkLwXCUxGYZd4t5XdA+gy/C82n6kWKxIK8IHcwdXlY5fll9+Q780UJgjIPZ+8
aOHEUQdiA6j3jR2jYMvq0QTpf5153tbvlRgldqjiYj/1qvTzOeODFatLXzMGa7CZ
SzeLmm9B9XQ8JC91gKa/bwyCYJScdBARn/NqZC40ZRrtOhtE/5FVXNlaXdXn+o94
5fcfrpqVxzHrgzoftvogd1P4lglC2eFLi7RCRpDEojcwvp1niMZZFbqxkXZCEiQu
XVdSIy8kqB5Z2/fqMlx3pSv9MzWR+sTf9K09LaF8VZngjLz7h6nibHrk/KcmbdTU
0pSB0ExWfzNYGlrOOLpCBUdgK9IBeASIlHnFJnF7MfUnGUUnI6UADXRGfxyasoSo
NWEgoHrz56NSYdZrmAnbkpRIppCtdW1vv0GEyJcSrMqVKL4PcJz0HAN5mOdOqi6Y
Tc+UIbb8NAlovxQysB/TPU/kmZbcIESB1P0bWOBLhE50tMw6FdMXJcdJKbHS0GYz
a2rSpc9xNigCauXNmL1TpOnZZboy85xCyIXrOLIZSUszIReB5SFpIY4caFJ30PgQ
SZvLnVmSB6lCmh5yBTZvkx2M6ILzkmnPnMAWST4OvzG5LHF5wz+O9iPS2xSBE6BR
PM92C9epY2BXYwx7fYRcnUjCoPMWBHsjXz7N2h1R8Q1aLjhMdxwkjzZUiB/+hm6p
UDgNSscs1AsiAUb33GPjbJ4IMKg5O5XLB91HGj8soxGI/hLeNnJPo2eTLIVqqZdR
1enmsC174n/aWWQz0BMwvt+RGFWBglA3VigVEW28uT8dbadUEF/Y8nySegsll2bH
s+iFS/OdwkZGGFf4QQbnbkGzb4LP9ReNL1JrhccH7KZ89UptoWupJDvR1wEB+jdr
1vNO4NqB8zqC+dc2R8R8vCL6Q5vL7HIiI9MrdiE9kmppxpyzH2gcofTdEzrT/YiN
fbSjChnHt19aHYYEo9wbMI92TZuFELvtxgTWycSqkCPvwWfY9aapMGqzzWlfv4jF
sXzveYy/7xm1y4E/KKsjcjYwKoSzMbm04qAkeK4vLrj2pna3tV9+EtNG5e3O+COo
bPYjNuKFfZkcd8wZ3D2AQU9WvsOpx6z7wpoPs0UTzl6AU5hWuskpS4P1sUdVFzaL
IcMC4ycJEqSzBI9d5W3N/g5O3z+oXmE1dD97Vsd/0Lraqd94OICRgJ5oJrv6Adqf
om655ISlmfvyshhmeUhwDzcFuA90Pn/zafph4iwIeWYkGcFRNMpu1NaQtsPhekQ7
L5LjsT3gh2W2YosWtiZF4962nDkjD5ZpFIbilKjGxQz0rW28rSsKi8MwWXcBmLwc
OI0oRwQDxXYUErZ/3YN9y3OoG/mC399KZJuSb/K3whJJSPaOQTvyy6LcfipxjYFw
DvN9V+P/yLgATfdbGzyQdUWN8U3NEoMIawsntuMOUSRhYAqMGAqgWlpon9dZrL78
y815pmcyNuqdeDEowgLw4Q827btIWn+oBjuVhFLBKn7DxsoqqLnPrxmNkDzMWfZk
vVJSQZCZVigtDqpNHrg3IW+I/HWwveyfWVF7KgCE6gw3Ju8J7cux+K16p1r1yeMR
mEWVD5nVkH3X9WWpt5IlY6v0FjRF0JyYnhTS1vyywu578TE0Y0tMa/Esi8RgHqW5
fYON4CSVQmYdR8BQaeHeUOaYb0Z8nkZ983uSZBiPyfHOYvH5vBm/hWigpDfblDNR
Lmv7tqGI8suP6Gv1XVVO6dwDiBbTgIJNaVv4tJy43DzIrgzffePATGjuh8ALyrCQ
huwua/QGVD28T8GC+2Vq+QO2c85LYDAYsgBe38JcDDAg//dN2D2eSckOpBymcgBx
zXe0up63y4B+GA6wPrKh+Hldm6Gtc4A6YROTwtOkbAzTINY6VE78hMGQlU9mHBq2
g+nhyGRMGxxO6eZq8Xw+x8nVpQnEph/cU63xCP6kCQmmM39YPkagDgy7PQ7TyAE3
/uUUizwpIgDLrj+pEddQve1982zvpJ/xxpPmoLrz8IQLcpegBOKiYiPdLNkzvJ8h
AAxJX2uN07nBiF8OUzrTBIEeMPjQ+rwqVAW/DoTjlPNXa1Xs+WB5LdFXZTpt6LId
PhGMqiJi5Z2/Kc6E01fRyPWTy8/OfPdJwXqObhuEQaZXq0YZYsSFVhheldurYd43
B6ahIrsY6gyBmP/Gnn0Cr+QiBJutm+FFMetVO5ylSIChFCgH5ozGn3iKCeVGhrVf
Q8Qke+2gordMNyNsF4kIxNIijCHyAaWWqUVdAmWwjYuBDRyT1TbqfFeecXkh51zi
sxt11gILUUNuZ/Fj7bhw2dqo9uUWByjUI/rn723PykctfohAAHFwXNljnUNZJN9l
Ob1rmDEKtq5MviLEvF+ys+Q36JoRyqdENbaT6O3phnVtQYWGNDTsX9VhtgXLtQ8G
yU8VnHMzz0QbH0xlZA/QI7bZx0YQAISMOublMcBe+VM7NlFohDQLV0TOJdaCeK4l
NfbwpmY4c3xQYJA8aeyxtlc6t3d94FK+X4P/LD70H1SljmVrcnus5vBL0rF3SSek
FFpYcPfLlyNd51FiXkwE5CxBBucK4CuZo/q4iM/KTlLbAvpLr5TwOc+kU38JhY8G
aK3vXiaTe3O4IWtWFAfVpoeU31L+aqNiuWdlrJQGQfGGfm4+ViikoARn8Dp1grhR
797fN993wvkIZ4A68KUvSlBAN/k3WyrphfZdnoXpVdURtvM6kwhXH6X6iByMgOt/
+vI/WyOYSbsdo2sNYJW00v1ptQfWZA+V2eV+Vu6TSLkFCmgGrAHj7E6ZeEH9Mer0
vPqn//NgoqVJmeeJmddYd5uB94XOF5awo9CKMIKz3zWGzDMiUcdl5oUWtuxB+f8B
R+DTrwyeVY+xvBP2lnEHAFQuyp65wuw2st0tjOeOqJ/bfPHl6L8GIZRzpXyYTLr5
s8tzTIWVbfCKyb3OdTr9c02IgQdSmHhWNgSOXn2M3YWcLEMr+9QiGdJTU+um9gaZ
2n8/e997/gVAeafuiNwgR85oKtQ8d8KgqHbuqhJG4DPl4aTZ4pSfsdUwE+GCKNom
S6wFK/w1H7QUBBxcU68nIOMQ6B+Pcj/klbdFHbe5rIcK/hI5wvsRryofbaDQHCnu
RAzz67m9UHxoM5gdimoc43JiWIRgUIp02sLM7BuW7vKcuB22VuYxDFkfmfMfyjZZ
SVcInT0yqupjrOZ6RlWK+o/oJ/KQdShjmz060IwoceHBEnL4xOQxOg0415jbUZrF
cJXQyWilN5rB8CTT6EDGQNEqZNV2NTF0gE3wkb3ZeP5jmqorBfvhujdRvjmRLN17
R9bTFe5TqsCOxuvNCASkZMeQhVrb07Dw+oHZkkTgfEsDzU168MDr6kQ7x8h0CUrL
1mQi4ouoeP9ECo9zx28MRAL0w3x8nQ00r1jsyQA8eCCa8Zuf144OHoNiE0Hlg8Ab
/wV31nRuOT/ffKN3WCRhLhx9Zj+iIoW5VtTCovi7Psx7FtSdc+dL8JOBHXd+SBxr
VJYUyztLTWPiV1aycNsHIgT0jkaQivPoBGw8Cw5BTCAbsDSE3BJvoiI/dKqPM13n
bWheouTRCIid94q43k6UamLyolACuT6oog0MKQYc1NateIaKLM49YMrl3ARZ6TBD
wfqwKCLBnr5LqHyTZ+OqSrFWa65IwLoi7FyihMPI/dgYUcStb/BOAzUKAuIdEu4c
esQV2ZIV28eo/PW3riybfyyZZ7Q/BgAeCGMfoLfK3uNabQlwga1e/kK1Uf35XDCM
wNRbL1NRb2Qa0C7EYNwpoiGEF8AKuCQRfqSRuB8FWFc+PEMVXr5BQ05uj+G4NaoT
WcaiE5vvEg5J6tSRmZ9uI5oyyQZY+T/jDmh5L4aqynMDYfr17yGFFERvLnawAqOu
VKDikqVHsEtW8Q+M8XDUcabDBYM1cxxyCBzIBk0odU9WudpwAHpurC/PLbQTbPvz
VKe83LuE09ZbZkQEl7QMYQxDSkKPxx7+2TWvyS5UhNtnn4vYnqgGydl/E1ZNUKlo
xqsHC7fOR1ZXqbZ45GGe4oiZBwVuSEVZtrrSW6UrG56nRXgU9j2R1AI8+etJ8/1Z
zmiL2NYob+DqSrfyhRv0FatZ6LQB01Odwe9gv9Z5nnIlxQ1weOqQICij+MjFvYg0
piwYPFxfFiL40rggWnwi7tf6FfJ6GTANxitnEGBAApLJjGgIgsEiKFD+J1RUcHzp
T1tL6JZgZg4dEbkvsB4shY5REWY+X/zTol8CzzKqTia9ZDMmkIM7KbVt1QQhnp67
LhFhygjzjM9Uu/g4WIXhBsGUbRRtiHjoP7qH4sW8zdLhz47owDHH/Nht0I7l9TIy
tSNGGtJmLl/HdRlfK93yK52gNudxo+sGsYV4QXu5kOeMvgqphU7gDvP4zVgWZErP
VJyDvT6AulEHcRFGN8nI2CTmHeB/RN4GDioDQB6Q4HFH5aZh4GHgXNzmlfODhgsh
IlUTcX3Hx4WnEiDcNx1lTgO4dMSxk+Bmax6UDOnSmFvtMCLNzETbA2arn321i5AL
gRSkp3fWypo/vhGGTk0oFRzuiEo5XfG4QztzHFxIDWmdFMHKBEAz1uN0vRbF6acN
Kki5krNZwVJthjAfjGrx3HbZSUaZ8LujUsuPc9sOXBlcI2HQ4dIlCP5BqiJHzcyP
34OyvQGRc9a4UkhuGqMBLvJcgypdRCd59zS+9YKPJKpKU5dqjv+arl1Tn94Ms/Yl
0C85QVvqWA9+xRGIIpjSBsvI0LLBoNE2iBXQ/8uyJ84iOOIX5de0YHEwOBbcY4h2
pXoVg1SZd9NibwLVLTv7WXMC8Y6u4cP/uekaYuPltDlJXY1QnROChLk8YLjlrwmQ
dOfWFQDPBqnQvNAwzSm22PsuiP2CLNQauQ++OURYU/F8OSlZjBO0pWHX+c41cPQz
pvTWilZzkvMqCScUfLmo2vzU+hPRD91KGWBpHPt9F9qeLGbsuKmNJFdZUqZh+AQP
hv7/BeUkSBhJA2eXTH8vWn+y0y8W/ma7k0GR07NuJ3ridtX7H3DhyWhkYKUx/WM5
HRVDOY0wElrW0zJqWeL4R7KfH0StPvHc/yWEwdMiq4iwhx7Bxv8SGPnN0pPysBCp
/DVTdAm5TM/4BAstoQteCdtlxHw6Pn+xS4XDnP4+k3AAY0bpdxFSrzeOISHHez1w
0B2kHyg3WvbuiWYMDHUhUiX7Wjqyu+W1BZ7ZRdYQiHtzER+NrfSNnh8rWY7NIhqH
fkRjJaeFE6hmOmmBaQ63M8U1QXk6wupClXpWwLt3gT5X+2PxF/DAjhGzcS6UOlNm
DWD9c7IvBlrlF4RpGWswWd2mMB8YCbB3jOwOhj6BcAPTlsB9glON3KKEeP+SgZYp
Y6w3GHC+IrjDdxH2ZJbYwxJ+F3QJ5O9Y9Jny5/fVNhCsqHYyicMK3tFpco+z+F4S
HT+h/iqUqzsxw56IQ+eQP9ARqEHRxzibKQJaAPssynq38bHh5YDdbZdhFQvEjLlF
GPEUoksL7BZW4EoNwufWklGp9Sd3a71EQExdtQJszS2NT4nQXYoBVt4FH1QZZOia
fHlNE+N+Q7O1j02fa4Thqn2wLbOqq41ImwJB33jDEVgwZyroEyaZUZkjpYS69cI2
zwAMcr1o3GK13Q0sBVFMK+nJmjBgoe+y1FVmKUKSC8heDaXVnHfPMXnp+xG39cVZ
V7+0/qRDbl7G33EuaOgMt3GVHR2FwMWGRYDZXxeP5TEKYW0J2OqltZiYaes8F0hJ
c4yMU8bfkmijWI3Q/oOcJtM+XBOry0TWHux7SiJXTQO8TvylywX/WJqEYFNoCuoI
ksP9BVOg1+CQGxj8LFndnc73Cm+h1XPTa+imeTXvAc4a97IaUrYzBLEcAhT9c8+U
p634O472Q4kBDdfFeevDVfOQrpvKIGQJVDsEnBJQHInsYIKziAbGqgGXYrk1Jlae
vZhWqL9GU9qLPEP2SmZZrSy09uUKqOlXDZpv9/UyUAt2hrEQkN9X/BQF3PiwNBBa
3p3TRPXI8RDtdkMDysw2o5GfmtrvT70UBUBbzvkXtSWHsZhI1vjIFOJZh5lHGFdA
5p05OI5ard7arKSX2yyqixth1ukblBKjiVfFVGltGWnU2A51PmuTvgXqACHuqvQJ
jN/I8/lcsUpOijmXdZRFlrkw+SBA/qh9fUkgnphul6oa7K4TG6Slxp6p8fNl3ri+
CuDDzPl3tyS4hUKdy8Y8Khbcy42By95ydOCep2nzxJotKnyMIjCGeifAyOU/XFAQ
iSCXn2t418cCs+e+wsG2C79ewRTjd7dgF56MA34TvHELtfOBMG4P+Kj3tFciKWOk
8N9DN0fL5FGctnwCB/onEIQpqsv0XcSSWolxUKRgMDtbug2HX6aDix7bRyMKdoig
hgDlGZNh+g5rrvIQ//Hxyv6SiOirolIFZ318eqUtHpN9EFscW+X3b7xsLc2ObrzC
iHESfw9agKS5ZSHC4vd/ZO3tsREsL7JLVjr4FIo8X/b5+1njOAITKoAsBCEQOSa4
ejcGFyKXQv9haKkdDKTbuk87jXLhSh5GMO0XB2UAtp3bDC4ePLbmaIxt4XQ7AiGJ
OF0oyyo3dvHaOAtu/2uzcVzHCpAhj8lGIecCRsI4hZvL66kr5uay0Cx/HiYxrXjO
6oCTwjTnDMKK56g4NO3dveMGNyybM4n5RxFKzc3LFYi55uTREry8Gv+0kKyR/aHi
JOXtTLD3FGOylQEOVS+BxlXANPeBq1LBMQ+HTcT9a1HvTXznzYlAJ4unzCMjul4d
m/bYIwS5zrCU67X57/+mtOiOkChJgYhzX2XwaC52S07rUswIMZgbuEVHMDcguY7t
xg14jqtQuisqE3/lIqJ6hgM7cn4a+N+MAx5jWByuNKAEBN44OkvjTYIKEHGQRxUj
8sAEq35H0Ri+0CMeAQ2RsVahwtm1f/ZTZuymH1pb35cn+eHWQMrMgLGN+2LNdZX7
Je0FjfPuGceVTro0wnNOd+iIn90Jd/IgNfNt08FmLa9iZwwTDcbM4QLwqWBNsFi9
JpOapx++SFQagphvQ5VD1xGg1HVbi6St0eDfyjXXsESqmr1lRR2JXI7uiPsNs05H
SlKmlgZQXsu4DJ858NIBk4An1WeVPivKQ3IP5HKZPMZimD+sF/p90iOfjTVjWkmz
hDPc+1jqwr9a5mjdv/uCS0Lt+zRfBvc+UJ6pxdXrAGkY9buhew5EfoCB0XQftXLm
HoEusoTkj8hanSezAKpFci1CzJcLvCqnFI2DYNqg7IX90pdVek8wyNWm5lfYxzXn
4i5Yimx06H2Dn7LCxESiXGnE0EakAH/DDznTYBYUMAIACBpShmYK5P/i+Y9PlhQp
cY+piwmrVtpNSAQfdQEojfbS5cd0+Ff9cpOiyW+yucfaqTlm73X2xQ/Xx9vkvwqp
MLYHVqsaWUW5p1aRupdRvmEKvVooDM0XwzwXD1W8vK8XRxkZ3FYo8KwTRZfgZ6rx
cjkrJZuoUaOLX71Wbf6Mhok1HeEMGHc13lVf3PoeGMhuuaikkxgicHJMoYJuA+3O
WUb2kq1dtiWt3z67dxbxLB/S336XyIeBUx8y3/LsVpHmztg8E4lom2z0x1fQ/0RV
XUJ+pW5pmnXBwwVO9mMt/v9cQt0DIm/jtP4I6V/hKwKJ4GvduY3IN3dwwvsciyzA
VBvpUj5d0NouH+t1oaIN/vGn4TwBIRx0oqkNPOSuviyM7vQMVra4xZlQ3aaji2K5
R/eyqLosd9aRTd8WRXZTrWPMxab+xEYoJR+MgzaZUpKGMKOendRaLax4dI2g9oLC
nPKCzD1JIrJCFe9j0z0GuW6TfWMqCJ3PGCtGq1B39nQ677Wqga3/RiHG0nrF7bH4
hfB0lcVQAhVBheBXgqGAoc7rkl0y813wIWSiJEVCnm+T6hzPR5rx/l8cnjXtFvsq
pemCPqthFhlVzpxVnjGYgUUVLll7EuHEYTkH/LyGMVRAKtvBmzCLfrdYDPnMv7QY
UIJFUhLZJdHQDXsXopCpA6Hr50ARHDv8ZDoiq0Ymsd/xPl9lGRVAI0AoOrnwm9T5
NoleVNbw466aNJQmvzi/iZc3jiDHlxEUdmY/sH8lIboPHTEYEedqNZvog4dtUF1H
XwoPPBFDZ6RqM4KUORG2kcKQlBw2ulWpPM7Ate4bPPjJsS5zl4oROxRuTTEoYDdS
6kwqfJZ1n9v6y3s558drONugPhMmfXt+qLxte1Jd+dX5RSbbSezaYDCpCghx8CIE
2wvZJwURp5gB7uDDuVb8bt936ua6AiCmmtTQkKup3sbWsE8iwUXwq778ph1YMMOL
GLRF8ivujg0TCgufcYuy+hvaCNE4outwmE9DJnSA1H1BAwnRsQ/rdsCgLuTe3cXA
oYJCtn/v6HR9ydqB0spfdajw01sZhJ83+Gybw1YTWyo9MooKCoFDKGOiG9OMEITe
6iw0Tp7AT+KJC1YcY/Gj7a4Ak1HCYvfqDCKg95a3QKigLOCDdNA0xsS6vkO8q+/s
t+awf2I1uB0kpPnlsChquE9hzYMb4F0QZtmOafnU5MKsTCgLURYKFc3ehrpLuayT
POeJiL79I8w1urWNuuW18VdCpOfFkNSKh8SCJJY6GDktWWWCpb0O3AfJMBvCs2vA
OCHGnCdh1bQMnrtppE5I/mHRu/31e21WN49PmsiBuK8skRyCfoaqW63LK+YD8Eh1
f4BF0BiPIM/ouqZBMUdLraLhnT8V9SN4aO1vV3Y7/GZyJ/NvYlmQZVhUw1xIzCD0
QvqOTNhhHEvWn5AnUm4cCv6MqflwToKd8wrK1Roz4SAdhu4t1UEsxbdzu3g2JgVE
T8BCSTq6mhX0rovnXS28j0zcTCcJilf4hz6+J3Jl9qUxfiel4/eVfFgrl7icQTuj
818poWukdjYe+RROrZy+5WkaFSxnBfX6rZuL+IJ0EhsDiVn43czoyVXn1BIwBLN+
TsUSLigB27tfu5cHcjxoAbGA+X5ujXPt6P/PN5iC+EVEmSIFREhahd8p2dxqdPA+
uPkLTQ6pASIxWqjoy4qvm2Gso7gmRim01O80reN1jGC/jBHwkwxMtzQdvtArvBtP
FS1cjKZtGJkiQyBq9XJOno3bss6S3Y6MVi3g13rsl6ZUA3eEUOyk9s1OoIEiaZYq
9bZESXC1ILw2okYyjGSG/4Ii8pupKHhlFhGsAKSkA3IpElAoOrIAITmGwf4XrkCL
WVF3QkFNa00529aatJA8EiH925C5Ikx+yMgdockRASL8m5K+VtHK8TYid22Z7dRb
J/yfxIQXZPhBY3BgC7iwWiMejBS47YNjtwrWltgbbrl1hBc+flcvfadpMvmQNtnw
AF+EZiS/7iP++ccBIbd5eyaSB6naIIOuex5xx9R+d+iEjUu6vwjyvU/jUbXwcdps
GOqLZL6wEMC9hkVtMteMiJL6SW4KXBSgJmxdKr66ybPTNJQUQWwaoZa/a6bdjrjB
lcEfCrbw+lihwKrpyWk9mtvrdu4DSy/qukD3QlS75Z0uRiMDoNTlaufCzstF8/Y9
dwrH7FVyDdzjQE1CL5n/YyuPXB89u6HfMQRi2JJNjxFoQN3tQW5ozvwOm+4nYm+x
Z7ry6z2ancDy4kbBoZIyBHBkGzjVmOXxvIjO401GabSe5+MllNUUOo9imcwmruXy
I8mjupvqacgzlixKBLWNYvooJFyhNf10N9RBFbknfnnbz5UccAsHSxsPsdcbb+3o
oJ3yDLx5Q0jc0BdAERBWf2O1dxd4Am5owGwsCIR+gkXyXA6XPOq5VNRU7G8Rw3Ij
+Awaf8dSEkaM2YtT4dL+mQDrXd2MAqzI6Ir+QPhSR/5cc89Uj1LvYHgRbvq1GVNQ
ogEHojh+uI7XVOvYJN5wbJQyvy48n8xAHU1BlyoD9dnrG49Go5fprt4/ctO5EGN+
8f7ZpH3detawIdOhlZH/z0KCXqhcWxa50YDNRR7H29Pfjgf95XaIv6uboukxkHPl
78AD7IQI6kf11oHUV2o6YvCtCdJQ3rEk1jFma2bFhb/ms1u+vFDds3k3vJhITsa9
pFoIMTGTpnvZaM7wLQM3kJ7J+74kY+QuLLR9EG65rg2VKqEW7pxffhk26ebMzWMo
OxKZaesFLq8c+RBE19DNvO3vfPJw4sLSN4Ns328UIn/FezxgqaOzDcSN9HB/mPIN
FiiNYcNgH93/EofOv80qMToSketDY+gQ8Qfl+UEaLp12k+OwJis0OZWiTZNnKHoq
ZI9UDPHGVt0jVcbd2pcjooNVnMCfZ6I8p9GNw9qaCozCdmP3VbSs2pQHPNCRzZHB
dfdyhJC4arpXhv4Sp7C3ZntFIJbncjExNA02Mqu6RIWMggRcR07CtL7WgIvTB9xo
b2I5ce/1wSQSXGAKWp0T2JhNnA4Xc2MZ40TyNeBbdlaYM/8rW4dKzPezutrySnZ0
W9x0l13q4u87DIJ7u7zjfDVvFW4g26I3zYQdjO110y7M0aH33N/b3qt4BmUMEXk9
ilzx+jnEUfKboBlTEomF040z/HfIUows4DOC1jgPxlmx7vwEzZSHpfQtehtRnFQg
3IHhp/QrsbuIbxY8ugSVpMNhNnc1g5lbawyq/fD0vPyKf27rjYdCC4qh8wIMA0Tw
o+nNKa4nNuo5GG5p9Q8DquVq1s1ujJdLKi5VUbl5Eul15R4wGRoas0xk4+NhL7+v
Raekjx93Hx1J1YDkuO/VBz4PuRG3JTKioS7SVRUi4p7DMUzGyrFJMzELk7XJFeUh
0iQZ5ow53o6wkBYJdThPUdim862RCfu7W8c9EsKgelvWkM7x6h1ALrs/Zpfpfb2u
n1WFHEVqnfunKmxtEL2NhDF2h0YF4RZSf02csUiiy8NSRltifoQQANphTW37zDT1
cFZl5xvKU0JbhM+xZ1WbS7fyVsW5ljIBIykcegvwJSzFoQouTLEpJA11nSsmn1gq
04P9DlkGJUKivVQX/tUsb0VZL+fzVQnNLpgk9HQrn8kFtkQ4Qjng/1B8GrCUDp8Y
93+UUAlN4ZhYNti/KqTmVU8XXxSioI4WyxshW5FF9gcCzNysOcNRQUCiwmHu+kmy
I2hCrkWFcRjxETk5mkD8MMig97JPFcAX13mYlIGqJxZpxm8FTi+P92mxV1pc+X0W
byiyxFRiotm/6FsZGXTU+llFJFNxdkcJ1l342+gBeP25lYZpkMWVmXIGMBbsBLWl
NYTdHM4CYSNLbKZbFWiBJOvUx22VpeOBzZSny9Wc7siEKuLqHNKdCyHc0vMdtg4b
9Ubk2rxeEUgXSRJoCkaZWjNtnD4AL2dCsOmNjopvDClPS0t0k2mHRO2BZzvUnWdJ
o/FMSBFqq6J2JuWRijzIjfkjPEa3WGRhpQzUaUkpd6xYWaJdkF4HjFjA0KNp8We8
wl/fZFnbg0QZu3unV9rPsD96YgAJyqlL9UVdfamfoo2ieb/VQK2XQD3Biapj9fTx
zjSs5HEZuhMtKUTWcuNGJm9osvPp0qmY9xnz1mn/+iKStrnyz+Ef+tQ57J8m20VE
49VFTPZrFB98y3uXgRqPzYzorlIm2Uisd2nhqhoPkUcrt3J40U8vlfw7jyfG7KZ4
AUY9VlQNtW5awgvlOa7S2IJ24z2g+UiT5Ee4bvGl0z+EiPA242EhtYWyGllt4LYY
zCdXPheKd6LTP+YnCxDtXtcKjcsdzF2FIh6XIJ5t0+IOKeXmgtvN2hnlrLU/dD4M
KTTOB0BNnOPxK52tR7x5FWXM+fJ51HrEr4ge9ZwJ7hMA8pt3rEaFZFBQ6oTxjWdU
04pqelb3x0d/0/a7Y4AnU5pMHUsPqKlFmxI0wvh9RqhFhmEASkTFseZTrZW/1JIF
WFs27GLIaVp/fOAz6bcV714XgekE9bSgitqeR4iGudCALNeC5Jlk4eihCnx59Vgz
8TkO6WRFejpBLob67aPhR8zLnrmSer3ZEa7gizX7Mf79xGNKrK65US6b+eFQL6Nm
T5j7t9/XE8n90jxTlxBTMIcPAd6eDPyzHOyn2z/6UrxjjvYCGRLGt+4wfV7GMJSu
IPmdi3Sy/uiLr0s9fuc8m4JlH7CxJgQdxvUvzHMRb4PudB+nGX/zjnrb65KYtA6O
05cAhf5bv8bXK6xVI6/zR+GtxRaeA6hqM6u9InoLUaODClRTqRe588HGz9dektj7
uK5f8mOLnPuOyUNb4Bf1BixkOU4VM+MP0T47RFS2lXuS+hrhDdeEsMsQMFnnC2ec
Hc+s5fvKUvCYOHYt9NlrR9ADh6BXUhKguTgRr+QOLJCU4dTOuv0KJTSYpKLBzY2E
Wnz4y81+EeTJybQkyeNnUjL9Eq1rnbboGlthFeLDNzWVhiJQ8YMHnxcLB1ktnL0n
1HSHwuUW2c6G6JsSM1nljTUgFPtXnSOYmO/rDHmA5R8nHcpeAQKSDH7yWU6hHzCl
wh3DLNBulBeAYtBKxycwCi0YjvrFUBKQZxWpxCcyXMJwXSygHcdYI62Ur6P6BunV
mIMjG1sJVTmww4EL0BV6mSxl1BZvabI4gMnJhAjBqqpPwac180U5C7YIq11OyeHE
/71e1Ap45SzvyyyHqq/YAevowQAYfJoJBHmjFcTwBNo02V3eNZ66a4BZxiofLDFd
rK9i0QmHkYRm+vn+AQfXQDWGdjMHnHpnBuNGa6376ZXSAa7XZFPJqK5ImYs+cbt4
tjm0lRd14CCnn7fo+bDN3ICySafV/o4RjUSuQTLOQfohS2yvEtgyif7EwBaa9cLS
gdYaOKQYJDq9mjs/fjx/qBJJmpDjXE6FY5brV5qxuv/V8p3JJeY3T4JllgJIHyj/
xqgg+YTYieQe60In3klQDxPY+d8PftPQqaNDRE4kYNb431u8U+3k/PkL03zDm5U9
0hY9WqTPWcNEMTYVnJoCeRqXAu+o+2p1z/gz6TxdAaGsOrAkhsBfLNjObhqMf+Sq
F7cOaE70VPgl2XJZPkqRMhpfo3YLbzhBf7OvkVzhEB0JHG8YaMdju5dxOQXA+5BX
DUlfd4kj1Klj6XG+qv9fJCvyGGUvZRWFAyIQlmCuG11JkzOaQuxCrHdxdVg+xVZ1
+Y9rE6/8PR4qypcUbimSBLgCINGDILsRl53OAQ7sGDvrfVO9cm3/ORgvb3GP/At+
+rwIFOoE66XTcOzmLVls/l4cd2s8+g25iPXty05kovCM794ebir18r8SNbT9MQyE
1QXs4yV/R3mpnuxFp0HAptgqTPmss14HUVEspUtGqHcG9ZOFgSwuJpaMiq4Lymx3
EW/ohZe3tcZl3fFUHrMURdNW24SLImTunjNefBwYaCfoSlSX7AVzDNPpSqzAMZVq
8/Kenj0+t/yPEIhqqJ0/Vt2q1LhcvjpR/QZj3nSTrLZJvH5YW+eBAnWLZzzFDEvG
kkJsBqMVA1eCzXMPqM//Rz36kjSTF7bkK/tiKOQEoap2Ttj/OxQaAxpQwbhSoqQW
IF7S77FNyFUyYkxO6XjO7IxJn6uR8QRAROFgNxOEiBpa1+EHLFuYzISC3sZACU1L
F2gCss/nm4ioDNnpPGNN4clpLKZxIBHYWZ7FnvwkmORuiLJURpPuvxl6bDll+9B0
H0MlxIsxqdIRrr1Z1nzuanHP4B6hsR/22QgGqxxH7wsLs8MdBk1ruNfUo5QXqGmB
vvapoemGai0qeQB8trxXPJG/AoXjh7rcTi0Yjsamvw6PrgIKeYxiZh86ECWDX9LS
Bs0M1l/4ugyv1/Kd+Bns77NMpYW548QfF08q7DnLc+36/c64n3ab7U/oAdTipTTi
Xv13rXvYUrt5Sn/4EVnMHvWpggMcUorz9EbYiLWEi+e9xukhJP9ezb6RKM0yhpAE
0+Ftk2blVzTvst4rW90sLnJe9+97/M1OrSi/R7x+VQZg3xIwVYqc4S5sHKy/6oJp
R5+ERXEw8uWTdVkwf9LWdzybw6KTr3e5qIFpkF7FrUJBTpQJpNuLtFmN9tgA/5OT
WJb/FTY5Ar6B51iqo0d8YulJvzAQHHGh4dsVOEZyU9yxWD1W1jahY9iWf/3DMqmn
MizowLz+3iSSzenk/A/xkZI77xrtw6+PVtkRCPXA+FSLQevSQ8UKV77ogTZhJEof
1QuQ7JB/gVkIT+5vPJMgLsfLv/fO7TQDp9ao+Dm9KrSE7Wimqyixy1GcybNAZMVx
UJ0J+YaGhgW+ZSGf8Z8uoBJ3eGViE+meq3GFfJPwtmUp+npU1Ewg6an1VD2M4Bmp
l2IH5m9LrA6sG3h7Eus1FPQEcNlw8Q345nqEkV5JFXgQfjpKPWyl4PXFr1cdA1RM
v5H4GM5ICDp+cS0fJbykKzNUdPaE04XvY3kjnzcWBa/XvkKQ0VozOXG+ZYjtK0wB
04sFwnC2U/AuV3qGRe5nrzUd6HGS8EMAogPuLXviv364ytltMYv36dlVJLDuQSlc
3MAR89u/+c9nfhszfYvej6cgB1NRiLwcDNHDqXwMqNfHx0Lunl7HwVBRUEqBBwj9
XvBlpMgbXX4M8aCEx4ePzJYQynwfyxlN9Kg3SDXmsZHUDTq1/B30XzESfOshz1rd
3A2PR8XOGNvuNHEbh127rNsflk6UKeA5JUlaydvIBn3PXepnFZeEP1QwgJGa/OP4
BWQ+LgQWl64v1ZZuBPmry/jfBFvMDOjr7s6ZzxPeD3kNeNXXTOIJacHmttSOyg3W
wL+88WCVchKI9HSMxvAuCDwJ5mulXzDz9nUA742rnIAhENaDiPh2X6IRh7gA5Yme
HHelqmq3bEDszTeIyRMrd0ffTYIL+xn5341wfuF7E/4PALftExe4q8CsXnYz/zPP
GLvHquuumxFIn+XxBbk7RvEzlMli0Y5yyoWVXPaUacOgddaZYZVbFpH51nrvK4k/
4sDmmHUU5FgDs4PbESMpap63Noss9yJav/rBdWteankLZ6rpYjtxPE8zNMcthB9h
R9pwYaJa+cVAIMExQBBhytjd6P+TNz46ZUX1Z3LIYgwpwloj9u/vHm4SjQkY8fw7
rP59+1F+1IbOHktu23XhlW+PGlvXXb2AR3HXLcy+LOFzkR+gJe3/+D/pbA91O0v/
k+l+5QiqriGONNdRNr2ZGIHHj7eOZVadOmhAmpJBc+qZnxb1/n7XyogUNLxSvEwP
q4ckr2CMA0aT3RfiyUtX5lfiNnAvDaEpbcNHKSDTxV/0cYZPogPgRgcCNH7utwtf
O3m1hm9DOKTtLmxvsKOGa9JuJtiXKbv/caQ8zDTwGXLWQR0Cb3hqeNy++oZLhzvv
RDXWGI+brCT9AHTk5kFjH/ea7FSsCVZC3EXOwGo939gf4POm3G+msVia6kjcaEqA
li+jI3gt2PmjxRqFHRt23fXBW4BmgRUDD2aI22B/+p2Kx019ioLhvPw9tel3z3yD
YuqRZZKKg5rsZF3Znu1HOJI4rj0SfxGD29A95rDnhsB4IiJBWbL2fgdEqDfnfDcw
yStIA/2a/dPq6eSpFSWhUgOXVpHao+Ltdysjcx264aLJi7hYp4D5lCKzFzzbIdTy
EPGVQsNBwx9zXQqSBR/Cl7bBrYuVy+tgmpxlYYEsATSxpshY5M/8v95RaJi3yO2X
mPLLozgemb5vKKsDSwDYnTnIxRPW2aKr15D/AhPPYkk49xpT6Z7Ixq8RVgZ3cPNw
dN2I+YgJgAISKNBdUIA9ZlA4bYL0vy98wTWINlJqUtzXdBHVPCJnfEJg4q/MbD3t
ZQ/zjHQBlf+VnOTx9IkmTz75mFm1Np+0AdJgc5HOpcKkf3YoAxjj2GxlWLuHrN1o
l9V+Hkwh8Vg+vvVU4ZtlPhvIuHMn61TYGZm98pJld1Zzjf2s1KR7kBJ/gyzL5QYV
hv+/cvDHimxRPRrrJUOeqtyfQA48OObHETHvIbqN7KiafvWYQ2niVXCBSDKKyBiw
F9rJI26/JJCVBIM5dSHKSh/3WP0dYZZ58ZT93Rrb34wYMT3u2PNGa2IDRVQiMn+C
49sMQ4IWbIiQBoAwEQvrdzhOsCxPTFhkmyWLiOWV4HM1yZaR3rZVCrs8+fjV5Z1Y
YTS9ZjTLphh9BJua0LaftpWVQH/m0QoIMaODh0ocPK6grd/roA6kkln3JF52cZdU
Q0lID5JcavQUDHh24fNmIcP6qec51jP1/b+bYd0sSut2LIgxykXQMaagjl4eNsCs
EJhmWLxIpHUtD5VEuL7QIGlYAAzvJh6UXJujD2bTK5P+il+yWjbhvj5n/KjwJi0d
emWhotlDciFsvfxqIgarVvOeZMcnwmTiSVYKHjEtecDvcG+mnLWW8fvq1kJ3tdk7
c0QHURekifVqRWtfHZ0zJenwIIM3PMDtrcKJQMTou8cjyDeagnpyq+k0Qcdjyxyr
ngNok0F9i0KF10jB4Z3eCHy4CxVKjtTcvXsYo5AeKHyTM9yHeJWGlPk5fe1g5m8V
/wlFIEUvorYIu74885jmDcC09tc4QJkpm2M/cQnjI1ZUfcTO4r0H95wq68UBheap
TVMPOD55W6KyluKfgEOlBR6HpR01MQHKhFAM4uX0cjL6ewt4QRr6AmevuT0KHEWF
YEOqDVfWJM2cJtGUpZ1BugTOjSSrGGCBZ+ZHVdTVPyWbP78ajLYBR3lNV4f6FbwR
iuRYe6k8+zrhCrw4XnURKw2HJkQaOexJQ5qv4QfnVhXr5N0jlmwf2xX6Spjx7jGu
JGTAZLaUpaFWuqKI6ofXyq/+ieOW7vpwU1RppircPr/jqCb7UuXh3TRRz2laE6Pa
cHOzFvt3jGVMMJa+k7Vj0IXnRCG+7DgDIJWq1RC1wVib4lSLYd6R5JPHtX+6FxZK
H2XFyNzc0pd/kJdRcdy3KHuG9p3EkIPO4D/MXrpW00Pi93rQE++wQMcIgjZCykT5
3Rwdw6bBBCU3UlPxWaozM/hStJspypyXoglv/zYybaUpHC0udUWmuCuNzy3Smblz
rp6rAZ4gRgyDMrdJKKHNgf1I8kv8ciyvQYyA5ryamPGSxKUxgzQF3cOs3xlrjSAs
VYH0+PuHiXCg2/UP8/y6B+47uKLsdEJpu2eYkmMF3juZtNZqP7fQuIawryLPCkYm
OPLH3c49d0Ix2rQPm9mdbkiEn91eBIVUye2BWIirkZ0+uhi5GUkErwdxmx9v0RE5
UcUtuWz/aYkt9JZDXKw8jqx12GUyXjuGksdg7TddsY1sbJIazIsiEjNBGhi6SMck
D72UooVRKFumFeYm1gDnU3f5IRawU8JXzokfWNJnRYIbwKXFQLVIAhlZxNZ24Bor
zktzwvGJ9BxPvq2da7WStda5Z8bqhYiRXbtpmpqvSzjpt/mve9/fRcGqvMPXdMZ2
sSkt0XidPGBmG2MNIJgn+dhnKDS/0AhJrdwdr7hCkehF4EcLzpMcilAo5jrn9q+q
pCfjjPxGgw100mJ30+l/QvOmduYYGFD1jpEyGvZy7NnVvxR3PR8EJJXkKJUzr0qA
nIli7qUbfRi4JmCMMNONPwXRn1qzJOwvKzSR2kH78ZptwAsrWZnKNyCup2ntKz9O
JpIcS8BpwIYNt0VfeogLxV/v9J0FOVpAr2iTexiUFS/NdRw68S2VZNda8zgEMlcQ
FiJdgCTbIncXmBbfjXiZNFttSZe/4j5bgNu2TzoXaAJXff/vZ18X9e+fqX1DOLt0
uFYsMST8/NzgnMyl3m4w7Y+aLN5jqtabTAMbhnc2FSwxT20g0p6ZiEKaiA8mdfW8
VmL1m/C+/tDqs8MLUGNdkkSitaZjBCqm/4DUSxnvqXQTsNnOyRdyvnL8bSyYGUMS
PIddgggVNpHdNWw249CbMR3rXZDwpwvTr0YqlsdDSGAFMh7ClDMPX3wt9WvIlh5K
t2ZGu2sHKQIMFh6E24WNGm+ARR0/yFlYHea5+ByJjUi7/lTVIE4g5PvvhjD/2ElI
EDYggHmUayPCeKgiNILSuFPEiNmsIOqcTkPscv9aQAin1my7zbWUCxiu0CmcjSsg
Dt0C2TX5YPE/KLqletuJWvv5UEqNtyojwT/OQ2CDhy3iv+pi4t5xfaWeLo+Fa5zj
XGuMjsTkzabYMlQt6tUoobPbsC3QBDen+giDnx3lQ20mWa4PQrfXN293REecrOzg
/ZY46MFlikPinBO9hrfG05hmKNVLzCl7sPDTOAOTScIFQ7LHM2w7QIg7KRNM2lFZ
vWRHJRg4EKHKxbak5fmJcalzWdmkD1HNvqBK3rFSNFXl8rLhythopDeh8DqrQA5D
n/sm+mKZ0uVWWQh/NsQ2fKlgjU+uNCiuXekw1GXNzB1Q0OF+raK1pH70HxZwsXOQ
SfXFitGGY9Mfe4/MVoq8kucqXInVgkXfVpQ25vO6kho7Jxz7coO8tQ8ThSlrZVdB
yUDKaBXskwb0KaBqbfZjren0r0Pb+BWWqdrJTLt4DxQJWoCP3/T9+2kXp73VHIHr
BNYexOYQglpHlFT/PbpBXXWVlaKkCcr+Viu0BXCQt+8doKpjeIL1WhdOusqNDEJX
STBSKIL1tJc/WkzjjyqJcPyWsBMX8sH0hyFGt8Z5Kt9iNfVvjR+I82Vw+cdBlJic
tloscfyUmqwztcpzb2I3pK72siwDdhjRVYPG9gVxbmML/43OpeY4CCK+bMgo/qWV
L0RmxEOp6fOBmhacWqsAL34INQoSGm/kv7KNQITTwfYbE+65+R47O5plAjKYKtgD
XpFcFRZJ4yrhMRt7OKI/9J4ka30LRBlgY0rfUr69YJ3z7A9YGOZ0ON8zHoS2klFr
k5mvl8qGghJTA/ulUOWEbg145qcPK8FiqTzcH0md8amjYnxo0pUEOcPoVWEJoM5i
YNiav8qDWuqzJHnLyJzu89Iuz4ruSbMzojGzr2Eel4tpSfTHyD7/AFDw/8ndsdfc
SqeCyUvVVULFLsaTZ/dAmeT7MCc5HecFf5wH8LTVGlFH55/Pt1ro3Bor3zrv+9/u
FFM60AWVeBw/rb13mtejGXHkZF1o0B5ewcCs4XhHSs/imA88xh4AS/z9XbTu/g36
cYE1nqPTCLi9YRRZuwL+0kdXTMKRaaNVvFkRi2sFo8PXmOqVPCImBP4jgQ7TFzU8
fdmnMCxErtUj8b7kvtBgn6sR+0JHtEI8s47NGCq7qu/cZmZ/eS14lZ+Ma/fCvIUk
rPbqaUnwaAQyOywB2gnKqBfNptkM4OhVfLYjGTbLmtAUSHIgPVRAG/46kEE/2M/X
D90SGT6C/A18jiLmH6mc49S8dk6SNZnIaEtIQ5yAiE/gU9JQYE+soqz7RXnBTqh0
f6+4XsGto218ueEKl9CI6BHIU7Y39tbC2aaD/5qG4f2kb9wLwE7qIXiHtWJqWPZi
HHGeuEa++LfQNsVXLfjFIYk/LDdPfYgHD6MuXsA0XCIQipQ/HhaYCIqcy5+JUmF+
c0n7hXb28Yups5wzEfU1Wdkcq9RoxwiWgNk7+GlnNPF27yXvl8yVyk/4O59XLuv2
FMq9P95kvUjFRcaFCNo6nzDPNbuLJj+uJdddRSsse5iYsj+JpW8l7zIfGAMxo+gR
undmzGs+h99by8uepNJKI9dlhf0pTL1IbM+QeVYgZvW6dbVXYyOLDsvZn77Ij0ay
s+9i2/W8gRM9CozuDEcmBOyvyByOsEMWpnBaRLek0HW4cNDG3JIA8CcH2EWQ29eO
vt0DJx1e1EnU3u417Bb+mVMmtAUj7G83EmYMfVpcOCKp0BWYhMxCBMPPSE6O5Ej4
5vOTPD8ZLCVPCPS/3KghJOlGT1LDvh+hwDNLTZH3egvkUksQHsWLnSmiuXQUMNez
CLxVsVYCL+xRwxYhWBGiqGWfg56q6NQHy0Q/rkMrcJJmRoaHzFEfwDjkpuT1LNcO
QGAMasqggJDztbLIVShZLVQ6U8Gq9IvZpFiqP0K/7IGx2y6LGIEpDrQhCSaAGku/
7GwG0RfjcpVmDKVtF1BhVgXAsxTUZbr19dUJ/C4zUuL9KKvLa5JF69FP2oNsdoRQ
7kv/qF7SOl+Q7YQqmEGlDhP2lGCtM/mdTTXWJotbed+ls6pvDK20Xmbx+63eC7Ec
cp/++FySKBD0FtUhrmwp/4NWKC/PsC44gVRY1FgJjlQWwSBsw55gKO6aDTjdwZgV
UsqUhVjhDYOvbEHXYevxsq3yrj43Q99a1BxAIUyb5DRzFxXoqO+/a+F/2cvrmYEa
8kES0Y1WfxeMFFg5nqDLTYg1Rmq59Or4ykA5wkFEEkKfuNrF1JU+6aRTKNqDFyR3
ss8WZr4ESNgl2GLpYeTZpC1QZc06G2KfTS8qs3qOVxOvFLhV7y8XQ5DMolgnXIAg
pkIt1+NmemgBJIrXHW7ngNzmquobcqJ4eZW7loNDZ6TlMlrs/lsnOP3g9+1d6PQG
MK4UBukFutkiRZ4UUJAg6BwNk157Nws2KJX94bh6P0OSZp/tsJao9UwQRz8k5puY
pnVQFi6trNmWftZnO0bXg/um8exJEDuOGMA/FbQ6gFO8qQYSXBKeDfN8/ao8uCZf
+PZZYf2oNgeG1iRaKA3ZL1L3wY6uzr3WW3Filkn497BwWznGNuo8dcfhylcp4ka9
8NcYdufddUtMQZOdcBaB6AI9bVMAKeBKMQHiWYwYIlFpP1fg4e5/MrPLV0KU/Xyb
UeEsBqz3oQWeeW7RR+0VKz6ZJmou71wpbgqPid5vDxySQNBUDPPvPlfq3AgrC+P1
1tlimL7472T9oNRVC3SrFCZQN0g6ZpwxdMFXEWvos3d0qyItJUO8GSoMoE3rDypj
x42jE7RxrXaO9wjkKSiHtlB6gENbqHKFuGDls0keaTAaOw9sPEGBfP0emelHOT8i
PV2eEDVtHCzCtzIvSfmnNJCpXHPh23O1k/2lBMBsLQKKdqlLXx1absL6LQtrjqMX
jvXPS8+QiLdAflbu+PQs/HN2/lbD27tmchS6TxvoV77AO606qNEqgQs/juwkb5FO
WhASW+s/xmepS/6xkSc6r9Eh933GNXylE0Lw8N8nZMbOlpGNHLWOQy/RIjPOo/te
+B87N2v9lyiYs+20n1ATFpz5hutFzqRpihjldp+2uYHjXq0iREseXa52jb7/nxgz
MXMCGo2+RkbLrpZHNLiOzwZURatEOzsx28WIc4yiLNIQV9ng3MOpXPu3ZgXCGl8f
JVPUtXQkNrC4r8uooEjhm28V5AMLjZdfB/Bz7cH+XQ1ROhsn3J5lF5Qyfx9gYYc3
UQpZ/PFZl1BlcBqWuC8mjwBg3nCf5ppM9XcyBp7PTpv9xijygeWU/oI0f25BbejI
MduSl4a07zOJiu2ID6ZyMp9ocoaR4w/j1gZ3rPrx5f9uyFSqQbh2x04qz74TOm7R
myPtS3htNm80oH/BlcilmvBbc5GLYOd8MFdj3G3GYdcWoo1LGhMilyGjPgNlXWZi
ta0TpQiOXSTTfJTtcw8OT4UMbyjOFUf1ewZWQMySWYDcwnpRvx0yGftCumSJc7Wq
I8t2ol9kBLNMCqb1VkfTtIStWYeAv2YNwCis74i/q1Vc1hiu984/BDG0uHPMU2F0
ZxP8r2TIHX7611lRb171aeHmFEeSuQSb8a2do4wjIRzWR33BVNWXgtFnh0OD+RRm
YvePfCg1NJg1GHPeCYCzY5tpK9q42jNiq9lMJ3vaQGJuiUiMG2XMh2P7UTD1ehYY
9hkoXxMY8bZbZD1MVLt3/w1m3sjX0BLQ1e8N0yhryWGfLJA7uW2/gLvJKR9sb4rZ
T2/Uo1iW0SXlg6VxdmMjf8h0JU8R6NkfcerxDeY2+RLN3XzjTUNpkeWXlgwI9eB1
vC0cQu3V522OwJ599mhZELuiinfjmM0lTACSIAdouBG9xnrWfdikyf/WIKW0y4Xf
kNY8AD+FvqP12KrAtlgDPD9v/MLLexiaiTaMFDBHkVLLGIJ1rPOcvkBs6sXaYOUG
zIFi/8vPuEXp7R+M7XcW2W5Aczvbwvir/UCvCERO8/RCHKDHAt4RPAhqzKkoIhCC
oj43F13+E0TyJl3TuR1wjcAO9lOHvgMjbwzCU4WOAp3lSc7EejdZPQ/0adyS2Zao
oT91Qj16yJynKnkhaQD2fQUOYQeqJ72Oq9L/t7KqimTZGF1zq6ulBLfE8O7XQzND
u4GNOPV/E1bjzBWORJrs4x8LGsYcZs6ayxitWZnSAIZ/u6hpauL+gg35kmGdR/fr
AyBj1MYeCgL3spkcV1rFuS5aK6nlmalqCjw1aWy9Ox2HZAHwEMz/jWvBb9jZ5NGD
UvlHsU1YhhSf2cHCTGXzLzFhqN4pd/I0nJX3YwvoA/fLAystMVbUHb0+1+Hk20ct
jAUAff8qHvXLrCAXM9qAr+kPJdXvcvPGF1+gL7iWqscj6FAurselhzxEiPZBKGP5
T+CM6ro0rPkWBakw+iDl/8aaeQXvFnbMT0mxdCddObtnYvIfT04jKvxr3d83d+24
o7VLAtHYGFotL07JTsawq6jUoWgnRy9IVmVY/iv6X1hwVRTNi9yr2Q4UcfuAeqzu
V8imchVUU2fW0WEMGpYitjO7ltTe46i/iKMU6VU30VLd4zMPRZhNiuO9adDKtwR3
U/k3bvgD2vFPXOMNZUgxilHD8687ZPp71QFCrKEu+xoVCWczjDVzG12EXPCUFEEp
MNC5TcxnTscZZu7pSdpmB5BtaZLjn20Updut3ms1AZEVMt9uvScaJcvmQraYfi4D
Nb3GwEKClRu+og2shU9/cEZ8oAGwTllWO97+ylzp9zqv32MSM6qZOfPOMY3Bywsq
F5ZUcZtpJxakHjYRCo3qZCrU0imV4B573RUV1ASZbVZK1TCvpV/IzYAFs/63cLui
O188+erGWuxD5dgTtwstMQb5vSBEbx+p3rd+HIDucE5Ct2M1rqRBSLJT04Ln6ToS
8gi2Ss3XECLOJQYSr9qxz9PrjqUob1Rnemm3p7UquzPZlp1uTJfHZz9ZUxYIOotk
tzIYrfsGcvLSgQRpAa7i5TxNl147KjjwP6h4XIq/E45N7WrGWw9jzG+zxryvTxhZ
sox+pJtIghRyeqQdUXttERjeGO8QO4GTlep3lXPJI4Oe5NgwMfAFjRwNa/6kdJPL
8yUZeECRgX1eQX+czccsiT14YLXOy0fig7Vcpb6eZH8f+MHGyyXl5Cu5jKF9pRIw
sxNZcGxJxAOsqlZCrNwN3W8CoedM4o2UAGwtmawb6Aa2AcOAKdfNL+zp59ip6H0K
oSjrZdNPHJm7zg+zCVu/iA6XckjdSGgYqLQeFiC1NXU4aVc2cm+x2i+X4lNARlaw
4xLg7eiqVTSMpxFnN1h8ASSfT/WLAid8Z6E8PhAtli/i5dp6BhdvPgOcWDH49Io9
/GLeYBoa3SPz6opqVO7KB3EBI1XdzOSMfhVWG5du36KF7zqOSk7K9Nan4gpFcqLn
mqa9mWKaUjj3wtWj6j9IOGQzSmizAjLUa+R8BZ11Q6HKgeDbQpRx+2YaTmWrpFqy
Pk+2tuLt09RwVpphkPkT/Xg+Rkm8CwqNhw2OvaDAMb0lnRiarkbiGxrX4gETRL2Q
RGYi5Jd/eUlbtG9uyZ6rUeAhc+fG0GYhjhl3WlasUTUB4ZnbX9S2aH/Sso3+omIY
bCdbsXGpDs0KY35m2vkdKNaOhdgFeGzML3DHy+Ql273HJt+5x18M0kA0UWNLqTyn
MAZoJkZHoBBZMJEN9jl/Kkgdmc7Buram4aH/nXyn7GYmahI1Gh1W5snzGHw5yXNZ
llXc2fNX6GEZKaCfcPJA7Kf4ovbEqrQEqbnzJ8JsTUiTegt1ZWPW8n8OgRMx8PEE
qVpha3jXJ5/yI1ae4a0zfUEcWahQMvFa+i36eYK4ZqeKHlPwpVVDo+lPOihBcc6m
wGcnek3sNgfO/FjwYzvMyDer0T+MIdSl3vMX6L1O8H91SLqUN0Ane3E0oMG2zqus
lrll0KsReSbfCf3Uw+2fdxux+jjwslH19hDoXzkK+l9PLJgB+e8Eo4GTW9h9AHbp
0JElDhlI5qca0RFHASSaSGzBWLx1uJCjp20gMH5N9uh+Shm4ErcoUSZ5X8TmYWcP
U5A2i2DQHlLz5OyysL5hTmr7KLP9X9fu+RZLO0ZeC1HlU/Ev75O84CcmscPlmIWX
Zz80vGcwdgX+iIJ2qOPB4NjhQ3Y4oJtHbAMq13f0gkhPBqjK1k/xGyHBKsiNC01+
AliTwNDjOurL2ProNJLIejJx+jWNPT7CGcFYtNzWbtITXiyHDRK65t2rZhM37i17
c+bWc9kVHwZIsfTTmqkFirsFQ/QFE6mtT/RgXGc3Cs1WTLZMY9zE1qZZTTxtjQ86
NKcSeyQbDXk4q55CG55EWhpMrN7JKRpUT3lR1c3iMlnwo3B+s0/MrHE8Z16ANRXG
0BbgvBQETL93B+Mh0jxiIQXp+KEbTq+QUKuqWg7m12KE0ysM/gTbq8xmajykClrA
zHRhnwh69OJmzp+ppd7/yBqiMiL4HWtWaxWfJCT2lpeUUGDUgIpsg/qnk+t13pBN
qXvOHhmxS/iCdUYKzVPw2GfcP2ZSy8jQ+Ao+Ty8AookkFNzrrLIe6gh1L2LdeeaS
eDs6Zk0+vqg4UwFoOUPj3dfyCMFws9vtibXqaiJQezw6Z7iRQJuVc9oDaOfbUrXG
u0Xd26MQcjxL9J0kXptSwjMs22OuiNDrFfJSYBv7u4//00Yoo2HfsWyoo8DvBlEV
2sgK0xbITMrNYnjPvYOecJUrQJ4JiQ2lCQodR1EKy7HolntcpMPKIyoDEBr2QgAI
nJHt5u70Pkh22Sw7goQAQcwHDNk/8JxG1kedxIUcd4uTMBDxvexxCQx5WxX9AwpW
WOlmuN/9BfTGMHjMkQ53YJULejZjodjiYg8mumyBrhuZzYl7bAeBTS6knQxUqKGx
Gq635pYwSwqDRn9L4N+CVb9IkVDhwcM50+tneYHeUH+MQTtHrc5ezAPeztoJ9i88
7m2cEJalTAKY/DkKXEvyWP19fATQTgCn5zqBsHk3UX8Nc5oSwXXWdjB3T/r8XPYG
8fjSe/K8I31QkWIAw/X8S24qlabysmFcbxD6keDs3cxHHF4zTxOEfHoHXL9IgYql
LJeIxVSVNAo+eeok9tuUQubi7qcZBLl8T6B55IGl7CWtW3lFGbVF/9sLP9ZtZODd
UvxwlzaudzNgtDAuKgIE8s8HiZEzun0mrTWiVMDUNbXFBIXxRCBKsN/NjcEaLIMs
qversCJVW2AmmDrXnib1tF2n8Eig5Q9hNIyxuqlgqIc8+YtLMyYZu1xjxBMMmkuq
AHEedSrdIeiJTmhh1V4PxdDdvdb/sVhtoDyWPqES8KDQiMNtxleE4EE9HFx5pPRc
BaWnFDTPtyNhTMblSzUmmzMDTby/hg+N42SAYe/IBIJR4y7EThFGO5c06zEPQP3+
g6xe2ZFVAzpAP1MaA0MHuYQ6we6YlciTWbn06E5G6ylkBt3R1ZeiYk9XpP6TeNM4
vltMn789+pm/U1GAd8hUMnmlTiiRcwzDsC/esGgN2hsSkNzaA+10XaseM7POCeC5
PpPXePgZCEe7MaNN0GABQT8Re2XVThLHPoq4L7++MbukoFYO4xD5Pi2Lm2zVRk9C
45vf1Ya053a0b+79imCKG9L0YaFXve6vQwBP6RKri3OmZOKjmP+k47Y7viGjaqRF
VPpwoFemmrWB05o8KKuHYXFGEyeCBRImY074MTLesL6Dsw7Ata7AvqIO3+GGXfyo
y+JToJ+1VSMHVsl54I0mMtgrok1uvK8KZiC9ezYq60D/RtyV6FCw8ddthIXfngAY
Yc9IIkqjKE9rjKFtMEPiJcRUzM7lQBSOe4dyqgYvXLnU2aXwUIMqNjFzEY/i1YAT
MtXaPYzbNZGm0QFs7+eeOtseJrvtgBJ9Glm/syQ2UY9FHWGTWnkKPEsdp9OZDNY1
Nj34gkrkIeLNFBhOlG0Sx9tDWC36BjEpkMFAOiabZM3yUPzTBcbZKA3zssWeW34f
eov/pXQ33L9vtxwzj1LWAxjk9kXsrwctIw4hE7u4AyFqEXl9Ag4sflIJRXS4rjma
AUMp3vXNN7Cs1l00ZIdtHxkV2RjOzLAFuCNlda7M9Tt84UiukDSxM5rfRaOZnld9
zB6AJYLShJDSYJD9kccEU74wb8h+HM7aiOedqHhgJ0U2MjvN9jYmrVHMnwQXo9i6
AKHW97zxmkT1bTmSO2BabJgZBqJyPel3IBp2nKQ/R/iqHKpav/fpluUSH50Qmk1j
DU51ZKoTsvT+t65VEu9gCxaY1J131pSC628nJMm2dyBWl2Y+amaRD/K+gqRN0pKZ
Lr0pXnIfOJ7bxr9r2grXdSEvVSpilsbsdiLDkZ37uol9h9gA4C9eu+M00OGhrEhw
+w8DpUE/8zu4kcBHIVlv+uZ0sXKMXmcJ1Uoth2lZG3pg8OXe7bpGve6/vb9/bNOy
Jyh2J9vZSYC/hesnomFeEfVEkeIxY56x7S2t/c2x4G7dk5Zmxp/cVhNddRyJyR4u
UhHVJGpS/JV/Ofrjn/z2DHyPS9OndslD4EFC2+Vr/5tcmWZPZZMM17dnQImQIsLz
UpamYHh4h9EUMLaApD1sXPaS+04WJYOcQ/IVNvM3c2ZyYhVyPo/cxVbj/K/2HtF9
dKotFLxinasZSvF0/jItS8um5zdydKUl2IwFO1sJoUOkiRsYcbrbCCUd2l3ZQ2Pu
eDciZv5+VY5VqKxdawlBkKJ/fF8GzR19m3GnA/coa8PRXJ/n3YHkrJOuuhDHkYV+
rAi4+oYAlu0V8huHDsbO7RcTuCwQTLCRUvdXvjFv5Y8i4Ji4KvjUUSuAk2OPrg5/
fJ0z2zIqOTIChbcHf+KSunml7DsvouQ52Ws4W/3LDKALTDD0s1GnH3dqY3yPUUt/
8b3xQcu0lZ9OD3di3C2PQDyviYlMQKl1l/BUQUMDTFsvsw04RkPpsGPOoBTI2PV9
PpLLb2x/2jGTVRLVmew0dDGWQB5rcp6w4Ne64TFFysjI92kEDH0fI9fG0xclR96n
OlC5BFAV/xPYR3uyEp7tiApKVH7X/ggyVzFQYIWiZStxto62avyYU9j7ZQ8fxuT8
Rx0bw3Z2gXU3KaOzrCLEnUOUzMcgriYAW9qH9C/JgNpMkGI+KgZOhoWgWVh/CGgS
0lNGOBFvjl6ozcZh/iShlsHC+AoaPbCo2F6+EuJLwlDEVicPRp228lRQEUC/ubwu
ahuEXF1AuWis/q6qSqO34fX8ieRNyl5v4V9rajcjI6dSTuT5z9hDBccF7pAtS76j
jxFOWaXFh7r3Z5LB0y/Yw3gF7iy2rDquN6paJkUg3aZHIJ9fTI6R/1QFcGLKLn5g
Sh4qZuOhMC4Y+iEtOSEXf2000IGxG0qaYUG80eXohUvRuTHBSOcW7f+GZQMozwQ+
jspCAJUdKfDNL6xEksJaaj108VIZny+YbC2cOED604qqnbwYzvWC5Vt5zYIp43E6
RpRPTmW+uj/hr6aPJ8J1DSIUV5m0xyBbhFIixEOnM61RoHhmr1we03EhvZOokPmq
UzxJPni6nGZ7ZPNgcBE9ecNU+m7noMs935Mjhr0hlR89xgkbJDKfkNPUidLw6fhI
rSQn9M6x/WQQKt+LGKPQT8nce36JEHEhKg8P4IZgC1rch+VwTVa75OGlZCTb7ZaV
MP/9o+I1msB/GfCgOeO4cqRU41F+aXRhbM76L22AXKZkl6c8B12Tvz+fOBLrDhOf
AK7+q66zVBlxjHywf/leeZmX5XJAmExPRpRCiodp+y0o4p/Yn2CSAR/17AKQlW0D
vzpMU6oEz2ya+nclZaMDxdwrT5J93niyL488T7qC3t/9m1k6G5RNJ+gfxEbV45oY
WDBR6qSz/Vq07tZhCNdawBnTGBktsnkpyWxoNe76e1L1ED3bvgo+IUxNfsEIa4Pb
nRyclqCVricdlRIsJC3Yqe1hZodTMfB0iAu837ozqkebQYNQWEwcpcU5klSUs68M
s/6TX7+WdgwVojCWLHLx788duC7piZUVdIMrfz6tjzckbwpIuW+LNo0pDrM170H3
Z7qsIFBi/R3ejxVAUwrL5a5uvggSp+QYhqOerhAnl+xA5TxQ3v4YguUH2EevVXjv
MSAWIo+zkB78/2/asfWw1pTRfMfGLeeAhqVj/2opA8mIgSJVKD41bHiYlycIX+tT
8mELNrLsx/0KbcHi9hQ/sfoHR2sWz7aaTTB0FhyWUHF+4U9REc+CZuuCo9AAyXlh
Nz3tIR6tGec3jXPvPTn7jwsh9S1s4AzerOL6MxigmaDS6u/IYEWDfUynuLJ6HuGl
XPcItZhj2s3i3sE5afrolPuWFBQ3L6CBUlkHRJ0RNmCU3CnUjOIlgyg58UsyCghV
BBJxjRVQOiXVQ8QNE7eUZglhgDoEXVrdPTzboK4ktckzA9tnsmRcQ9LSyq7Cb2nd
++X2juHgJK0TFS/JAWL3+XDIvJGmHCVP1QefzsoNtHiu8xtgP7ODzNcMhL3baQep
rnSnLsTJhLziSLwjX9EdB09GBzbG0tnrPhBlN6g9fwI/yJotCOdvgH7yfCO68oWa
mdNnT9wGrsCEoMtWQAsOwjBhYxvoNF9cDA8yPFQdbMvMymwORBPzIqWJLt4P027q
7CD87MUOAk1wdMnLG2soO6uvfYYGKx0EH2mdyPxROvfMo4lo6KU8QsabSHS2C+gE
tqCy7rw4m2/9imTUz609k6gbXAUte3PC4hhKMFbPiWuOZhM9fpMWahclgRh1BI3g
xa5YhOP1IjKxRZhAcVn2qkBaUGkvDHJVc3ejOpsnXsCBZjazt+X7786cbkaSdq7i
DSshoa9JP/yWL61JTjhKScJfLdr9XQ67YxFzPCVFGDywmZrijR3VnCLexbXS5iSl
OxX737mQDXmi/fp+41czeeB5e7VhKLy6CmYoC+8PEW6MdeWGFsgDzLzXxyIqHxrq
7r8niga3tcG4aEMaNJIoBlCuU0rx6RX2MCmzLxWp6dSYwlBmxH/tw3vKf932jEw2
hPFo9Gu/+hmA42ePC4EMNNgqwlK7Q84mrp6/og2nJ0f8aaacGXR+t3+X4eskGGFa
PPywaqs3auHkw3XaHrCUvBD0p06daJBGvsfpaul67+wTDD1PLtBtBAOGByP4DfQQ
muchZAhM6opR58N/ciRX4TkLKDBWh1pwznREYXLqb8Z38Eb7FUE6HWmyrUkRC1aF
izUNQJsmeudrkp7nqJK0dv5TLp/920n2x2YKYTBT42n5ZnaT5lsFeWsej5dj2Jli
X+ISQlH2NsjJ0iUWmOD5MDEZNa6/GaH6q5w1IcIFwIUul8cVdlkiUvaggysvh79F
xOzFvD/XQtS73VNxvqKxmpMazQT//OqB6jmgSdpYUBZgrDIejs6QOv1vX0DzPTTu
diA/KJfxoLB5vVvDAeid70OI55sxWwkIaO9gcDvruC9kAq2+WMAh4XSkBKg0g+Cw
L+1AHFrKO/Hbqw8Z7z1rSmUdrM6+SiikCBAgLl/cR5GTu58ppi1A+61Hdjxr26Oa
LWzN+XOBH7Kvm6EXF0WCOuYoG+dqe8Wg/owv3S9VIClPw73T8MkgaXvW32SNzS57
lrO50j4OQAM/kzoIQh+D4+0v/LIqE444UZ4vGaqO+WRSe7jbszwy9RNZ98m7DFyY
Q8WQamqg5uBrm75NZ4HifNuS9lmi4VjY1OVOkTw/Qalj8OisR7tIM7poBGMXcXTZ
xkWW64j39Asc7SsUt66rnuN0eaGY+DoLAdEmPZroXt6Sn+xuQzDbYNxXISck1+Mu
UDBp3BruOJYRtn/yjaiN6pmkJ3BI3f8oTJ1de5pPPwFNKNlAw1JQhoItKdgBPgQR
88brWaVF4Xd0UmdgzlTTbZau80FSK/vs5mMIT5A+VvFltBjwLHkm9iCG5skXaVui
vDmf0lTEDXBrCQm8gHfZSO7sfdk9GWom+N4lONth8XDaqvWsu0uSHBUxx7ttfj1F
dzZs5CYD849XVoWjn3Sxp8ym7LcAjUGI5s0iy6fbB5dq6aS2DI3hPHo8PT7HfgoG
vS5bShcqHlbQDydj4jq7HU62AO55B9Dy+MwKvelzGc/yLV2dHfgBJDzrkTXwU9H2
GF555+h7iY+qLKxVU+QJ/eptTKmBqk4RMtUFly0I4TU45vFOIgxK5qqY2rM9fY1h
dVAIlBitzlucDUNkUGowom1bcW0PlTDHXF+6ImmOBoMFcarSag/FbjVIWfgtLukr
XHbKu1MZT23+j9ukgzZYxu+zbloCoCrt38oC4BqoHi6pew8aQEva4O3y1AVDTWzN
RhkwWNcH4nvDN0zugpbc4e2aoEXyjLg0PDDyTAgnQWtReBFq+4ywKQgeFq5UgwjA
NV22o41td9Eu/0tN1iC3h/YUBiaso/h/Cyxs+7weBoVSMLTzSaKPOIhKD6tvZqVu
GOh641K7iUqZXO8xZg2LfWy+r697Zr9ijvFCDUcwz+b+v6t/eOZ+b8qTkLB/4RSY
pmmhVb8Kq4+wpHYx72QG46UYRJe6Tqu/HQmISZ6dKS4z5tZVpEgDzHshzMiN6FbY
JJhFJ0n9hixOcW43XcH3wNRWFtYr1TuZBsUvshSRXjqTAmGYm13Zp/Ov2qWAl85i
JZQD0UkgT+/HM9T/J1Jd9ZOhCXKYtpUzEpM1N0B77eR73xB++LI8uTAb9AENvxPg
lwGNr8Vc4avi8aCxmOEUqc4/0KvFBgPqwZSwvq9fNAPWmWiRvkOzrYVcW0DRZ9rt
0+TaozY78PPLadEUhlvEL8K8jDULOMnuXnvCVo4Lat9OxlSfC/X7AMPxk0aRxH6D
x3A5A5oBPH4MYVWMPqzXOiGgt55Uc0qnuhnTtHUWSxLrnfo0YHHVt6pTfQJoWlcR
mCBfw6GT3UqIb0Ie8t5U+BFHOzt29xyNNtSSRRiDipb6GZ85EQJBym6wa7sgvzeW
XsGTdNxHmYlGdyXmObYpjk11YLpeSB2VmaHjwreY4/yMtnIXP7tyHM4B81XjmPQp
HPerXTmzb5Dmk7z7XIrVl12NOH7Sj5uBwt1zXG5R8EdAcnOjxnSDy8WCvsfWly1K
VxjM2E87r7fvOPPVHW3sTrlmYNlD+MYMmjwsJCTpPmxtbkfkGOKqEySTc0KoY4e9
iEKh1QTNqUHHLyih9axy8JBtQFGi2dPeEnDy8NrSwwn4yTFco6t04uCefYGBwPJj
scpREWE/FEuMNAe94+e3Q/MshLm0ea5vm+RRw0haNYtxxxSLdcGZMpwoBvcx/Z0B
s717RWaTTT1bNR/6xKAUPjKj9+v55ed4NZ5878fwbsmzYpnD7HyS+WZ29Fw8BrlZ
WOZOo4lS7tms9hamJzcwJiqhYdOyEchtCGfp2a6XAWg9Zbjg7fkRAIdJ6hlfK5xc
Fi8gYCjMZMF31HBveKR0mxodDNwJqVLfCvqJDtR/Bt9t1JIHflY6NxnKtVL0Nzug
9isu2Ribr0gXvfc6To5nmVsu1chWrN83xFIdjdNU0CmfvevwhejwUHyLkh7RC/GZ
IwWQLZVNJMcRC+K7XZRpDgzPx3JaR7/V73sJqku9YcLYMjmToIbio8h82ECkuD5K
VkLobrM+YT7OGfbXCZPLxKyz5zaaD0a6ZTRQrkswEZTmz3v3Zsurk5tmCKtE1LA7
iVHNVruPsV+PShqqvzxmvhUKpa4dZfk+lzGzjnggt2Q1olUJV2ARnMvn39uheM/8
K+vRtaCQt9v8gJMHhgY2gDMb+5MVC/UQ24gZpnapEutOWnC/Qb2pnnt0783azQDO
Oo68/uu73cPhlt7TqRBVbA/qyrjSmzYuPlDDCwwWx+bjUkVBbim14auu90Iyrrd2
VmgDfrLExUYR8bz4gH0lP0AHtRjbpESvlX0alR3IToTgNPaQ9PZSwGDT5Ksm2wFJ
gt4xzzHHGLshk+9NFx8nS3WB28mivgZVh/j8jEo0R2QQ4lw1d5IhGB6j9jszrC2n
okKGsC0ZuwqgkJZWMfTL3yQO5z0mNL9/76ZNPshRRjkpS9bUgbWAOPI3Why8NMs3
2zxaHUblSF70M/UQmJ5TBk+cZVUW20tZQj8z516ObVHlw5mACxKQ1xQ/02Tmkr47
hm7snEjC5qIWJH8yA6Y+mcIVs3LRjsTtUIMUhqIolCYWejQEr2VZTSrYmIOt9mUM
Ab531SZv7/zYlzZaxaxFYbQqahU9GBCM1lvq22BAWQDci3eFKuuAUT7wsbA9wXEm
Knq2w1CBKuSaLF1Egn7ZLb0us84pZJyAG8YFwpt5e471squ4Kd0rvKoGRzKFpv9y
P64elV4cc7MDcbTrm4GjIwClSY35fWjclilLDy6eR4hWatQ5IPG43O65Bk+NHygb
ZkTsnRqJ/WA1OHdNFGgV1sJ5iU1Et139pM//d9MGz55x0+DcsYdnUgvziWrcxqfd
LxEPDx6pAhG0zUaGcedcPHXPf5/864Azhy3lIEaiCtE+IGqImyYvnXsNKudAIVZo
RVW8zOwwPb4kZjLa5pB//CgNIN0LbR6QVLgZ2VzTMa4gipYcyx3MpKPHuw9T75ND
R3I+gas6el9TJxxz0q/CAbPJnvNE6U54xmZNFh/Idh6QYfIofdhnr+UBnZ9ozYna
E94AI/b8KqcwNcnn69belIKn2CnKZQ3YhDrAmG+DXML75c16qYccne4iVDRFm+sl
O3nPDfj54vmkau5gr9cIJNW9n9NsUQY7WN5TwGHTpZ84tOpayd0NDZ1r0KN9avTo
R/GngzHn09JeuDGa9wIAo/jBBs//vrSxss40OhtvQzx7T4Ydd/tOd2EhMAcbpZwm
QbOuPzHaIoPfgeE3+LP+scFCOUSqsuD1ICYb8G8lQ+k7+d43I1XwC57KlNwXqQQ3
4NdmPqOFBXpjJ+1dOgw7fzrOAcL3NjhfDVhvgyZoandT10pyGEPilJ7t/+pzMh6L
Gw/oKgDrJOlX5qLsCfkveuD2+gQTgVBpgT7bpn3nRKlF1qEkE25da8uxxHB5EymY
YPshmEhNowa3YBWo9uiC4A01J+CG7GfLPd7DPntRFulBZV+euJLB29l8w8n7vFss
Cila2MydLtoaNgTPocHc4a1AlhfhOYHw5t1rNkkP0smPyFpWX93DDTpUx8/Lpk+5
Js9BIMdLtdcQeKThJ8eKHPIqTUqhB9fTUZppr0vQs36WWRfTXEvAbMZ7aLdWZPqV
y21huHB9QCAYfC71MIdrGpy5TMCxq4ptmKdqWJ41Z3seFOPz2a3p6Uhq1Un55qzo
NGAToIJtub2mowybBIl8eqIm7B55Zbtf4nq9cuHvnNFFr8O4wTUwy93Z/rP1vmCR
lS18svk86uaNE7ZxAZzhih1MTRm/zRarOkBtzkfTxYCSQ+T9kdmRHTjAy0owpgV0
pCMHpeSbSiE4FLoodfWBShha/cu7Z0l9v6xyZX7gbDFLjgghxIcXnUNoDa82TdQP
h18HfF4mtXe62/BV5IG1LS4dZw8nIbiJkA2s7ycNVj01uRNIEfRYTtew00yVbjUE
TdKTfovirZhG4XmQFriGKcCkE8HHqaQ/9QTIH58pu0GK67+Ke03A7fz9AeQfp0dy
SrjqMf1cA9DQ9Dkh6pefXErggoh0pfNCjP+GnHUg1tNZIUB2cvUveHGh1SgQebrk
4xyVQMwZVl2idERezYjTnUU3BTG29l74uY7Md2QQC3bN/vJwKb2p0itMWpcWkePR
gYjfyBCmCKiIxX2iSLIBzJzZs/1IeTeLuoe28AnMfIyR4MkZECJ8vZuExQqQJMKe
EGJTDSuUcES8RHKg0mvz2TnT2/TXjoL3nyjCvx39qFTJ3YU/6wGyCMttTEkhBvvI
WAXFRaSUmBw8tMYjk8mlYGVa0OftvJju/UegGLGHBVT8SVZ+m5vPCCFGj/dU8XCK
gFXsijsSzIOJ5n5lGc0+ODTYupZDNJJC3P+fXmSXpD2sHJifE206OTCOg2al6Kuv
lrgD4asoZ0oVoAAltwsgmGrKHIIRQUxjteqUwUA/WOXC7tfw+xmCE4683itRDxlG
dWZIR8kDP64p7wyjGR+Aq574BIS1k0wtLfL2Xd9Vmk0YcxWhW/NLIY+VVTS5ugRu
P9Pr6uBGOX8eLcUhq6MfdwiCqcNM0O8lEve5Ru47uXRpoWV5IrwKwwM677/wHSHc
ZA9LdsCOVmAWR5MrpFbA4eZQCTZmUK/5wYpNNCFDEAWHpmCVPZQoWYckNVb++03S
0t+SIiihzQUvkfqEmVH7sYe1btMAntqMd7RFst9UjQSPIJh+UACJNK3bXvQU2XPl
7zVjXnRt/pH2+sm/ataPx4RJKgJSQWFrE/cW1PR6R74hUeIq6SnDxUoHf12eC65+
PCkGMqaEoTTL8+8my3zLWUYypzDbtyrD0Wn1mMNsZQggqg2exNpQlvvcKPzyiW75
CE1EWpv5ghH6gl4R1YMf5ganQN/woCCOxUrxuhSQ9+2OZaZYKNC//1jFQOwP5ioZ
J/ZOFyvrgX7giZZiD+zPYYYLFfkBU/Yuwk7fZcMJJ2gh75S7Zp8no2slpeaHT560
E3k5u2RfR49CrXJPwLHrdoGemLC+2i4iJ/eg8UxIEjrM87Hdw0m+WWI/9prSDNlZ
eamzmlWXWqp7VgJe51FvQVv9hINPYWXq4HqxOU8c8lVh+7py/lNO15bjBtSOUWM7
AJ/9gbtB0UVkldwsGuCDqQx/yBbKQy84lHdlgfMpNnjnh/maQmZmh4y/tteAf9my
nl30Zm7ruVOjzy4RQmwaqkpr61kUaeaByXJQozR/8ALJ0XeCvR63KiCc20hcm9Qc
rbH72MR8Jt1nNMkrpxFqlKWapTgaIIXygrX8FjYEiBT3dXb5xIcjLZXis3am7TO0
WcnvY18dpdzHWILxurxrS+GyJxPWCPQtqZQyCoIEK4/hVDpYIzuY2Yx+P4KlmvWM
/CI+69Xxpg2VCAdHnctzdGP8Aqc1ytiSTbQ+sbrF9ngS6iUjGAY2OEYi+OI1Q+bE
jymW/RJXeZwHwOM3YP8C93vqOkvZqoz7ilyJmjGLAA/CU2xklycCBdVfjT8uBlBJ
0mN3OluOluyTPaz8+e/cAPmOjhM6h3ntbPdEYCIHOxDb4UW7h91oBhFE0df6Nu1y
rqTJ+BwNc/Q0yvrV/Gs1ZH7zFIVPAItTT0RlKy2xJsD+zGgvr3hLuk0k4ls/6FFl
qMtVXDuzUXkdf0kd7MgZNZHk41F7eYdX8vRLn7vfo5VzvyvfDoNOpZQro8ivKcvF
ahRxRHbszL5sBwflM/jhjHRRkWWW/oXDVp2PFgDOJZuBFJDQy6npMx9+8uMs7m5P
cazzi1HxeLtThbgK31hLymOD4ZL1ZsrEU+TO2YUh1qaAKV54RfwkOXkxpNIv4yMg
o1nJej5CbX2NH5WCJ9YTPPNgVZ6aN7dY0x7JKexDsVjh0e8uztdP7VpXz5XaCQIg
KoENyIHDy93E7bp0RLgUgQTXMpdKhJzhk778FKsFfL8y029a2mEPjdqZpGUq8ZXH
NuIbRde4I1VNX2N4ssjSqse6RinkJfx40J2h6vbfdYLUF4xZFpQ/tdBobRAVrk+P
5IH8or/YcqBiFW0dl8lYcWrnWZ/htaQVGu83S1zBPBUM/mFl9xGvU+W6EzPLE2Jt
kmmkr9VCmL7kxtp2Vt5nbVF9YEULXIxFHcQkCrPyy0jaQCa/v2lfT/1h5k53pRJi
tyEm9Zrk3oF3o13xOZxT9pligr6J2k7d81ol2sewGik5T7jsniRw33Ul4tR5f2Ec
aVa0pp7oe5XhVi358cj65spC8w7E6dE/O0LX2ZgpBNYNYpP8Ia6YE8lqdxrl2kWO
yvk1R1AJdyrUH8GAJo4WJIneGrW6wX+AhFI8QlfmbHRBskz1NlhZieChyk2naPQv
2IcZ2AXcc6TgEOxOde9/42mvLTMQOgWSQimKVXPymMCj9Xw0F0N9rYPeo8JBqNCO
Q22kEU8d5vBm3PU9DeXRqQ2Q1z7s9f98QlSR9xxFkwqpdZR8IOq449iUjYJb8c03
JmWR6JTqmkrr3bxJ3mOUziWBuE4ZQTwrKaAXq3O79P5609Cmg20mho0zcSudyreD
iIyN9HNjrx5Kz3VVK4/I4u1L5dDewjKd771KpKXqV1l+n1eOgOA86zhT6eTx2rn1
toygKbY7juJOOlfYeRLT3d8YdBi9Y5ADDKSGvMTQET2/RMZmnhtLWdTU05fH0OVY
2WuLZQde5EG0wlA1REHfntNwifw37pFmvdPGnnzjXYnuQ3vjvKHuhD9lRVUwWYs1
qhhJuY73iOsXhDUvwRc+GiNKVLTUK5Px2hnDVQC9IJ27UGAppsb0VDf/wP9KrDC+
xPYZ7fbI/jMeU+TDTjibuIR2oG6IB3FwJHbHLGK8BcYsX8LejT7NMVp8Eai+u/P5
idsdjfv8Hw0goNkPIK3TgZP/L3YePPRr2qCRcrGdzCYfJY733IsKxIrhhChG0RJ9
O/UWNeUmvDOIWoEmMd7p/LKXb5v9mfAhMHGrcEf9HoCEfASaG8bHjKa8xAhQY2A8
zatwONHBhtpw5N2RIgkyzX9cmAbEEWzWpCHTwbiMLLPY+vSPWkBDwYnnolCXrNmF
gFNQMkpY1uTl18eY5ja/lhr94mor3GQBR5ZVi2avdL1hKIN0se8eDOiWy4Q66vpJ
XrWauaTkKxesHbekGsd+x901ArVPCxzXvFDM+WClFDyZW6kv8mB2gL//CUx3rKu1
roJPEF/eyymjRnxmtPdEghQYMVRpcBkkHwwimYNi1uRPkmgy4JJyioVzT3i69UnA
Yc38TrPw+1yqNm7h46BYr/2KDY0fDmV6FooKBSSfzd3M1Rx4RjAv9OUyFRnGuclB
wqV6H64IfCWZfIAqCohL/UqlbSjs+32tVQ80yjFRYQDIIXuD3Tge3vDQ2A+FqMoR
r22Btot9PXc3VMMrE3S+zJZiWfrX1XeY+kHxxReD/xnCv1Pfjfvb9SR0Rfv5lk6/
vC26YxLy0oD9GgQAu6K1nVcS86HnWxK5Wp6t9/QJ+nrBbAxmDgmdK36So/lIEIkR
16C73ZAjLbStMfHFB5oMqhQFKydDvkFkZXx/QM/94NAfs4LnMY7O0krvrAnzoKSF
RzJzSo/U5jQ2/v53PmTR0GNCgf/i4waMpvGb6jDrWvGeqfZpcf8nzx6oN7WBjl/T
nhiHa5m8Bln4HeflLaLX2Y/gbvVU10MxfEzNfjNwD9GizFtpQWJw0ZWuo5zZiG8M
c7CbrfixM01m+LYoYKolZNemY7SWkjkYRXrTS04gaDUzGCa0Xi76sNNGfJcqCR6i
yny6aFPHKZ6W9yHqc+RHa6uJiB+Qobt3kQALXVS95i4eUN2WehFUQyaMl+3emDkQ
SenyKhK1TbWKnsIks4GfQI/EsUJzsi729M3gmCbq3BoRt60jPDlktVQq0xN1QImb
OFKMV684OB+pu2iRaXm3Dl2YgxIUNRui2+sSX4gPyUWfuHl0IhFSiB4RXAB/v1vg
HbCRjuMjPXogUrFD3tpzpddNGt3Dhqc081wxwYP0ksljU4mhSfLRLxJEqDAQR+wF
ue/5D5/RvJoun8IwOfDuDbpF64+ZJO+RSUNXUElGMr7mR4REH1d2Tii6pfGqmYkU
jYu/s6lnEZoNhUO5DuqN/8t3o44vfeFcjusE++kkFbcdLD5ec4fuf969xRF4MZcz
Pl3pADX6pqG3cKU0DaQIlib+wkv+rqYyAUGIiCJlitSux3a6vgL60kvjwBmZCsCA
F9PSlPo32lbENLo0w54Rc9bcqlVQBEd3s5IqkJ5vLdG7uJHAnndNLPTfn2NT4IH3
Zb6Z8I1eoyqppM0zwrCwL+nb4D4eIDIQf3T8rZGHNhKh8Mijej1pA1Xe+fUs9tuf
RCuun/a4hyXJYtdN1d+vDeFycJb4bbIg+4bkm+kO2xg0WqVReLBBZecY1jELQFzP
o/n/kggJyXZkqX/B5vsqaNyDuhGTH+D0UH51Mo+h+w7v4jW4UaVp6wxymnRUevCQ
VlqiP7LG1Y8o+Bq02F9xwcndK/Csxap/wE3Vkmv6OLKMSz+CspfG0kxHeZtc32Io
l+IOiEVt1hxgHjO27/BnSKOcpSl7VcwbmHVIJgM5NykatE8WFLE61G3Eo10ObmGN
FGHH9AMXk99yKX+r4YHHlgM/7PywUqF1fxWeFTE/LVxvcnyI+K43MbL3+xYX8VMe
BkMWqLjNgFP4mMECL4nxK8pLMJ+Z1APXIpxg3i93eGfZE7iqozTw6j9EDoNMKOVJ
iVpZs79/yr3ZDBx1tgxELsLPBabzsD2gdmlugd1r9zDmyrbXwxjCG9XWwpZ82cgu
BXCzIZuEaHcDxYfqDts6O4H7uHyf2Krr6Ky4QKdKzNgw9j8CPDcpFriEnycfoCJT
dnywRNnmAMsnxefbGOquS7iUbto5vkq7XQXk1HkbflyzYGV5v0Q4hb3RrewJlEsM
yX6rOn9fYeP+I9wWXouysRIHBG0XCHa16tnHI2vuyWk8IMImgguGK9Zup8HsfoNq
NfuR0ywsMBAFUXZe+rSASGeAm5x5jj0KqtMg66AYRotMPOzlpiNVy4F1owJBjuKC
SRnLzOKjmvZaKKHE0TTTjVUhTbX/1+v5qQiTN4+wlA6MtpnhNuh4M1RmFh3ZKOYS
q+mS3kOaYWlI9BEjQpQ8nihh+xDRPYmOXHtSD0sJ/FyARWIZNxRjSDDHJPDA2qQr
YWr+by01nuo+gfiFJ3ubfvBe6La1wqvhyGO94JPr0iWiXGzIgu3jEVcZl/bLmYo7
dlpaYdBQbwFx8ZswXa+cqw3o2PCup4L7kKwN/hu933ttggki6Els/J49X3Naqf6F
opS5Y54UlUbmy16Gy3ebaG6VmYKbkGAKIvFoY5N2K0vlW/HxoIO0qtcla3mMotb5
pMtMSfhN8+bnA86WG6bpC5Fo8oY8McNmO6DDWEbEo4ld3VndbFKLFup+3mkoWOx6
0lf5ZpZrpW86/SQUVvE7Y4JKBEwu4xU8uNX0BiW/RCRzMtAHqTojHY/zFxOZdF/D
0lU7lGyrrmiXaNzCTY055Bxa46QfdM0tOsyDvd/QcBlR/CM2U5NJIuIAITMO8Nxl
B4s8t1t5CXSY69ZN04QQOptUf00FutqaZKYK9ZrI87SxSOU++j7OkXccQXcaUihw
yWIZvOvxB/PcxTC1EIRP1xywVDQW20X2dM8vyQYWmO5zXPGgjGkMHZP4HfvIH92c
0YMnQ47bDvtf9qU+kTkCvzrx1wesfEle10klcb9E7xTFlYGhMT8gG8WFwIVOaPhR
shDWVHNj1pjYlCqvgnbsCQBKtLKdYXYaIvGQCgnEHFCKieTaBI1Ecx3vmSlgjiMv
ZIvPAC1UrpBuEBqwKlqcYgz7VZ60dL+mNR/a0qcU1sypbbAcgddTt9y+05LWzMOX
Jfi7adoKALODhdkVZfbe+RTKNGiCGdBNZay663ERfdOcpNXIi0bWzrY9vV5gF69F
aKDVreewaHmQyCUnwh65Z933TTj/lx00ckAsf+n+J3QjBCQvYnY5HjrrJJPGqK0X
7hIBIA/Djh7jJ8vRmMWajCBwLHjOpfxoJgdPdPrYUccvL7ksM9Ge2JclMMqNhraG
0yX46X4D4TZVWTjfXhOUW3JlSeFL06D9XdR+ycTT7o7T7P0JwMP00fXc/lhmWBon
axB0OX+BH9RNP4boBY24YPTxGT50X04R0WddFDEPA5GwdZfWej9wiAaOs8A6sStX
eWf+rppLzexy7gjkQ9nZ3INqXWDA4fW8rqmvlZsmMlZBdaca9dCWAgbQiKIgNnHL
Edii94QvNu7WZjYc5DLFfY7XtZerKE60oKucO+OwGcLhw6V0b6knJU+2Do8qJz0V
mDMr/h7B+3dJRGtA+BpvsNHx9cctAUYtV99uD3+FWZOeJVSHNGpJHOkG1NKX0cAE
ogZ2+JZVE/SwRUwDMRJglw2lP+MvHEskFo0mRMawy/HuRSio8b73fXuwT5FGWbmo
SkV6vbeOXPrMhJLCW+Jc5sGlT0iC2vqxcK/sPbfAWl5nDumafWRSXtFVvzgHE63K
DetMRmt9Z31qio6wE5+LX/wLqLIAGA0vSz/Wye+LNBLmerQvY/InE6L5+2iYT4em
3Ebr/WWG5TKz1aZf9Toe2oL3p5BrVxSty8FEO5HumpOSmPGd++ZWp9Ge16VEykwK
//CrvIuk8yiYnQB5oHJZcF4XS3AAjmPprXWosGTW9W4/dQmM4GnIpDDB/yxU16fJ
LcvQTjZA35COb7eS1ALCX/d4FVw3jTnN21KZwOF5Yx5xZ9MXfuW+/LLxN8VdTyNA
vlVmha2n3x3JBXYHUFddYE513Wk30y+954+hrXJ8KJtQYWIKioautQWKNLY4Fl0u
RpfBUkWv2yB6SPjeWlHaNTBCPpsIAtzYjb2u+pGQ1FoX8z1JGVvP6TXWrlOT29Tz
RlW8btVuvtT9QDCBG3ShI3R9mqhE6pOIan/D3e3sbrDKhDEnexbhtk8biSXDZkgT
R8ZhPctMAr9V3jmBEFYkl3c8PGDWntV8WmY+Y7uyHu+RJyA7YIZvwIb4pjI9Eg2H
l8GuF0V+a/ndChaBYdx66/JTHIdnbrOzBuLtJDBv/5w0ScLalPOO74YrTkmvJJ4J
b46sM5xSLVJP40WX98dLKCYqwL4NZs05Caflb8ufPZ53BN0YubcM9C2/Eqgcxcmx
WuePU1xosI9uOZOYnnVBvbDJG5Lww5cePcDzYVPhGEm9TJNbzyvmLY0g/QiaJQwA
/O1jLL7IgYbxs+mT71IWESxe1Oe7Gzf7+okVetrrd5RrATKdOhCK3VW4nWKDzKAQ
8nUgvKH1PqS91LUVSlJbUbKXD48h9BnQuVbSSyxIfG/1dbHIC8/XENw/SEp/UJDx
FZ3rYZ/KwoRbGCPVrrNwA8V/FS/SFDdFs4vQb6vNmZe0njQaw4mlps/kTz3oQNTo
oM7nKFEtkClPZjwbGAp124WOyAnWPfCFcKsXkOOPC98X/CpukUOfmuFzbCbmCLHY
b7RqjnCubano8IkKr3/pfmkNxaZpdrezDurjb6dlcxO5iMTtuzfB4Qce5GIAATqE
tDy/+4OgoEEHkGUkY+CsLUqsJsGnbbGqCNYLEUKhOtTHWg3xsCql/RZysnqFqWgz
kFwiG97bquSrDM4y6tH3S5Vrd/lzDtJluxqkyj0VGtfVEJxEjnwdzByXXOjMSdlS
cHqs/OCZKfKbp03SDGY0+YDr6aJplejCeALrWXbtEbVUlOhJl0657j3t08mTbBKy
bUeR0zaDEXxWUcyOlPFLdS7BUgvaJzRw6Tv/u7o1QMSHZxBTrF7GwmsHhQRCAsuc
+f02j957PXCBi14D030h7tyGgLiPE5MpJoFj8F4pY5eqzQY/1c4rPF0QMOCK0OwM
TqrJ8bt9K/tunPErXCEbg6butOuIaSoqAYjVvvWG8W8VAhDq94Ln3RFYHA0GjOHE
+VW5yBQxqbdhuKqwGLSFJ8weQJCkcYSbezg+IHHELaHUg62qzFWAP6j+eETCo/cV
2X+d/W+vkojb4iPntnEFItdnNm3OhV6B+4joGaHs2uUAlZD5aNI2dUmuOXcFpwxP
X06pic80ut6LaBZo0MbNS11FEvpuvRkqqcbcXWG8gOTTfEqYitVkrXFuZvkw31iy
JhZgqTttesuHBPUcrr7WCRE/ZUG1kDPcBJ//3ZkTQXja5MsJgsizP904/O4nCMYV
XRH0jyOAAfsHI6ICPdGiYHvGyxsnXK0fEIt/bu261cGzsLXdj5bF+WLTRYuw+Qmc
XeKnVHVCW8jab3wj6cTYAnYhJNLvKOA0phf94coA4olOWmBXiJOqTw86zfnfRHSv
Qi6648svjnPcX5f+0BUUZrGZy3RE0ep/m8jmmHM3F1+b/bgHg/XtgEQot+d1fPDm
9blB51MoVKs8i+CpUa2ew8cgN9i4bb2SWxjgvM3KRAa+uUzEsL4OV9fu7MXTuJVb
YCyAOam9/wHvUlZ0Cf8iaxxoQaI07SBDfd/UXTm8jn33KJldjW3tO4HULFYuIX7r
skoEe9B+seM5xkL7bKwedankzTPN7rhsaehkRuqototWD/EDoZq3zSEp7g7wScKD
97KkfaTbJoBL39+Jqo8uPwmkWeF716inbX3Quu6lZV2AfHObenmXLTGTnZnZe07u
5nNAZ2lMMYiMXZu6/zqjIwJ2IvRFfkMI1t0pUTYq0H4Tr6Q7R9YhlK+MkemNy9rN
dIPIK1t+AxR67QqWRebRXVCbYBzemgN8cIt2vT6Q7YG0/Ll7rTGRAAoiv9zGUdUu
ephqYOYUHupZW2yei9Ocl3oXjt7v8g2BZYejneSbv82iHRr0rpFkJjAcuZch58WP
4uGv/2opXfS4wEBzInILEV5dl2pW5D/+1niuDtANqZKSOQXYY/S5zXB2Ds+L8cqu
sEhucMn9DzVBLpPkd+oQ7uzptuTCjTLSL+KqsCXx51rXuvjuUTTfK3m+Jt8eMPlh
lBAUPo4C+1LQxWQjY3rMDrTZ581U0gpgJgMQmEsLkkmpgDX2+Y1NzYlUxwXx9lzT
0SZM9QZVJdiouOTtt++il1WpPoZlQJG8und5Jj0uwhGMbMDNJhj0sU0+P0VY4w1o
FQ5aV3XBaWVW3Rxd6B+vRdih29xsHQvZjgkSoKKhTd70CBHFZxAQ0CUN9DFrHzJF
yprwBRRE3hwjUoHgcoDjyDuAfAUw9qNJrd1Pbop7EkJB5qTeByGOO058ql2IyD2q
bOpNK6ITQs6vdQWeftvn0f+Y9o0hDfk3ER88G7H1ei6cnIBciEoCtzIbs4SRtxYW
gsn5Lb7TMLeSsRgEoP4aiaOj09zD4oOawZnhTpOhc3j1zE+ITiuTa9wGaPHb0196
XEeuCmHqNBXke3PJzdr2c8y94eAnrN3EWKAZC9ImHwFyM7YSW6QfHMm/KDTSfGuf
IMHpz7E5mvz9C7FcJkXTuS2MTnTub4c2+wxVmvqZrZg2Oxx4SF1Eg8c+zEs6PwnE
rtols9LgPGUElPWcKj5JfML4vom+HQnGwxa2NXVchzb4HEdR9wlBo6bXqhQGPAkX
v0XyrGj3ksHVgOIVFSnoIfo4QX6Hji5hAu902nq3TfXfJ0sEqjR1JhenXvqdRO4i
fWZ1BQiLKD7gnNB8yBzHZjL9ENkDfUgDmfTdMIzhfKP9/TeFDnsfaRLL7Ud/McG8
QV9E072TiHko8kQJoMBFWSP0BsfVpVOQfDElP24l7jdACtL0PhBfnfuw3RxcTBwy
pzKuQniQpKkZrJyImkzW2MzkkkX6pNqvLw3yaKg95dprlvZ64bM8CGBc1bAzWjBr
0B+EP12o/uEUm9F1W4JU3jbJ17Uikoc4hR5rlbSP/VHEQZz0OULmFyBUja8FOtD7
SYxZeQxaOvlfjZ4WlSszp7SQ5aI1JfGa+q6mNv9rIIQci0kds5cBf2BD6Qmopj/s
kT8UHZJG1GzbMcvTnz0/RUUDRUF8s+deRPjk64Rw5vX2B8Q2s5s+86uCzgMnrjr6
5OqmS+ePM1G1gVr0u+cLc80oIYzSbjqbVBnMfJE+ZEIuBeMlTVt27I4gMBIvgAcD
3dl/nQjXe0GS+lOwWEMXKLOd42pqeYSc8i9SfMHQsyr/A8Q6OvGN5b6rZKlMLXJn
OQFCdmMnFHX0FporRUv5HimAyQ8aBb1t4DbRVvWH5XnlALv03k3Ky//tDDklJH9V
Ab67y7FspkHaV3QDKnjWC4YglA2P4zTDZF69ruC9mGiyp3wT/C5qB/ieAbjCU6ER
pqyJV5PFAD92SkM1BTRJ5U2xujozsq7aQKWkESBDk1pNtOsOaqc+vxbFUtGn2/px
BLzCLOEYQBhIE9uEMYjND8ZkwGX0Ek6qs/6/S9fUPwZTiD5OvCU+vToaU0fjHzuW
R+ntbF4obnay2O0yESSrahkM6cubzC6/jumfbd+YPzS3a4ihazgUlrn9UF9iFxd7
UnBBYvL9WoMWxd6HF+bRzoGQQgjREJnDIiyRlMon5iJDv3iiX9FKuxf0PjdJd8KB
hG4H4asazM9olFkNxeONHDd7j85wDa6qJT6TJeX62m/mnvFYwhcrxutZbicRWEss
2mnQGnX3jeWAI1GvtcUAssyr3mpVVWTKrdKErc8h+eL2ekl2W7DCR1QyO6h4mqv9
AgWH4DqLHE9xKXe6J/2LR2U9XmRDn4rfAhtTGAvqNZmRgvh9wMp8AVTpXSD/DYPe
4K7Dw4dZIKnGK727XiK2z/HMy2Udr9svXQ8IBqXM9lpun/Xx1BkOj6tOQODXSVJt
f8WwXsI+Vvk5v5DpggLBEtNeoLsCjZqxMzCYsnbbyro7Fvh0qxO24o+SoLn3eMaZ
ehwAPU+07qmY2JFNJL41vBxuVQM3StaFZHkOqs4EvwjzlLdYDRK2btgjv5aC5/uS
Bz+9riE5tG0Li0QLwxnVA0IrdZiyKATaoITTILYcXJPqhByAo4r+qgI5JqAKLBVg
1Xtcn66Ulq2hwBX+ndHQ7FwgqRzNVQI0cs8Vq0JcpupgAhu4QD/oME1TkJlzSxxA
+L5yA+yn8kh88pRE4PG6oHZN2V6+4iG3lXGSEF/LOxA8NkCsrQIXIzfRJJF7llv9
0iNRa23G8kP8yx7iontZ3UkNvUNJxqV5gKJZCyYGzXWRA/QpHmHju9u+xrDuBlyO
XWRLJXClzAdi2S0iJTX7ZDta6UrsSPvlNo0D35NwLjUmvo5Ipx3JX2ITTAVh3j+x
F3M+oAdgM4jKSjkH8vHvepmTZAjsxOxUap31716944ItsNQ82Q0C8P0i8xk8Xyv4
qnzfCN1hLI3mrxGoSFN/5ZFfe7XcuZlvRfIzhpzBBA08OZFWk74c2SIVraife8iU
WNfTo59+jQnJKXop+BLd86sSvEBrhw8bm/LKByTgwhL8SXIgVZkN80DhQD8eMfu6
iY8hr22aM0nt7l+6sxzLpLBECZDfUaHch4UQ89Z99xJ8BTo2dO9J95cRPueamR/X
x5+Yzrx0y+Ho8F5CK5VDiveITI66hWV1DW6qHnAURM5/vBNkx2x/wtu308v/ldIZ
iy8l7U2FBnxivY3wm61omW4xRI0wezQYGz6HvKqxekdRfkK0gMM8JtJNB5Ko5e+i
A+og75eBZLohd/O9TeAhMttkMHNCJ4WfFufREunTEvAhINuQQMXwrcBsinjv7aKw
mHoFMcEJPYOZR5lmblyVMu4iJDC8KLfyyJH1qpj4MuAedUlhFSSk7NFQcuqcgdrM
kBTjfofyKx1koEaW93xgphs+Acy3q2waNNlQphHPF2V2Teb+5Mkr9vdgoudyx+xL
PiM/fp6IglobG3d2N9Pewi4HbO6Dsgmf/l9jKe8e6I78kvpfQCaJutWXv6px+h5D
AuajitlIpMlOurOjk5IQwt3dz+j5yybo/1wPZXS4OH5wfl6xvHJjlT3Ti+XsvA6j
1l14WEqEeuhL64N3/s7loORjlcW3ZIZI6kjNySMdiAQTS4Zb/FOEGKQ/uJCMfYWn
COza3sHyw7hGlcEXC1jVtFpwf5UaxSLVgj1ZhKWWNENQi1WuopqAz97rLsWSufrT
OCt3FzqUMkRIYJf2Q7fXBkbSyP9O5cX6HMQfFF2j5kCC6jHmclFuBNDVAIgVdb82
fxDt5rVdZHPlZ++dTgjFxVo+V0Mo9bonn6mlc/1kUAsYWMY6Uu2zZQSQGiO98Moz
G88Df97e0nAo+lHTM3ZVMV7eCdMJs10q5ALrk0tnMorVlHDZRLjI0mX3i8pZL+d2
KEi+YE0mdi/OB4pT8xGzIB6fRy9znzLPgdj51OvXhr6QdQfykShy9L5pVyqXR9fj
153JY2pqeknTRB9q6eOCVhPaNlu7vJEVYdc01XRoTh7MgDIuKEnCSWBsrRgU7mDD
qvFe558N//ilv2ODae5yUYArA6jemm/M2iF9no4WqfD7KVo6xfaWxd0rD0eZNXJS
kH3YA9KLfD8+E5Mgvm8kKnXycL5+xU+C45Dj9VGYTAwlubNMGt2As1CAhy7nKljr
uwQoo0eQm0YqJzrkO+zmVTNAwCPm9zJjVcpAAHDuq2TLpRVzhw29QN/+NiM7SiVX
GpposYsntaA+uaJs0lIHHL9u7jVx2uO8wDhalqVzssK+ypKNk0fZiwSatPVnIpiI
5Z0JRqytxMYX7HJ4pNqsdEYXsWD6rOz6taSbNfW0Slt7DC33mn6utjoWokpI4YeO
kjojL9K6faBfNH5SsMY+kC8oYIhGg6lWM+U9AUFOshRpg0qrX6VZFrxG7HibrO7u
3G7fkJ+lUThkJjM7IwLedLt9hvA7MrkMxwGCpPpLUuc2w3Lp42To2ENfYzeV/K7z
NIyxZkWk8G6KjMKOgiT8Gir/HsuDfOryRGE2sGSRfkcll6wE4m7mqo3bB7KyBchy
ijyTIMngfvQXPyKX/Ox09aYk4z/XbyHesZCeEErNeq21yZ5NXt6JT93HGuphvoIF
h7H1q2nhmlC4RLjxyPlgJ3HDBy2F8HdY3RpT7xF0dfJhnGpCbG661XC6mP0TeoSR
CKj2+qpjgUR/HpXlpCjWqPj9qGuzBXEuzP2SyxbnrIUd2ZUMS3u3JIOCunaHEirC
4jRJP5/w8FHaHcQVikFZ2bcgnPL8mv6usoVyQe52Lzk5hgJFZNld7XcTC1O2VSxy
T/wgIUdj0EaTpDJ8xcH559brm0NRe0F8XGw6JqEFmNonVQmn5JLLmmSifW8Ufd7F
fMb2Hvhn1fmFVIMvlHz90UnhM9OJKvnuPBSyio0cU0muO37cUriDJHF6a3hg6Qqf
slUG+KyFQAytG7pxT8iFNnrwth7X0br9oJlEHla7xDbRpLXZBi0FE1VZCwEMPDP1
sW126OMSTAeSL96rSmPrCBpGLoumjpHuaMOC83LSXQ1TPRSylqSEr1JJg6B21XsC
bcj7YoHOfCPXxezWVEVFOBOIwTctgle9fisyyAq0dx9eB3Jhh0PuZpkzyQTeebe9
e4KnBx8Lm5CkO4RzliBiDXI7jM4EZNSYboCFqb4mcvRn72ZlXK9rI8+nAvJTjmlB
9p1F2MjJsxsTrKxrj6Z0qr5F+cmH/sW9z4uXMVxUci594ukCBjLdfFPoQZiFLpZ/
9YVfQYbZ4kgf5Vmh7qfBVYGjpAaxHulkq1ICiWI36GNlNC3a0JA1TMd1VBWnJIgL
q0zNtE9BOKfwVdvOKgJQyYPqnotcI47/bgkJXgJgOHSPrFcUqPH08QAmKcRiP/eR
vwy7CmlukPFu4QHe5uRf7oC/7Jw9IOqx38J2AEzz4ONki2y/FqSmw6zTEekH8EjM
23OgNVWyqDLJMatJ9wKFaIzoaljTRfjV/aXPtUQcKq2KB+rgvFdZBjPXuoSZJ+fw
toMmBJ8i50bkG+FY3vCR7997G9D6oNUhkSwRyLoJbvDtvjzhQyl4rQCiGsHQSEK/
7qGwjqBRE6ykk3I1SFN0aYwxvEhVdSWk6DXTjC0AcqiLYCpAccHznwlVdITsc/kT
vXO9c5Fjqh3saz/CgCXjmPdk+8p/J/R0569aKREN53YdODo7N+3d24PYk4R0JmU2
HszxARe/tW0B90hvVopZ4F+HEYcsCJoo2bsyTPdRG4L04PscdQwMupye9Oe0P60+
6pwTcDQxV1vPcuh9scw8+T91pxZ2f97htIcbLuHIpQ9hQav/3kWpZHePubycPWoI
CRjPTdYZ9+z3ue825VR8Iv2dD36u96beLorgpoirEQoAXbZSW85Hf1t1l0IAJBZw
MCgGZo0XYZkfupSOTQrsNIpbdkOAwx/414BMvS84VyO8ZimPHptkRiSVmk8IpxGt
XgMxtv6QDfWFWXVjTkBx5sX+t5jidS8cKxlqv/HXiR0nz7OrfVmuZ3H++Dsi+LoT
BUSFk2a3hIFxuhr+CEgVrvqss7mbhSzBQ7pM0PJ4pIx2noMYlwT2MES0tvbglnNt
L15RV6EI350G70Fzr3BsauzlgrASwmeq60AqIaYUCQFX17ZWcy88q6jmUKxlQqAe
P56sJJuPmJxNDd3VnaU6AHHKgvDr2cIyCwnLB0QLacaGs2Q4aOUiaLaMbALqxdP/
pdqA+dlb8s7cW13fjfKWuEetu6lAbMdBg1zo6oaUcjDY3grFmfJHfZbOY8xCgIOV
tPZ/RsnOiR9BdRRuaMuq/z2tmBxbFWIAKj+i59FJ+h5hdXZJI2JX62Bst1kd7Vc2
J/AMH5S/EILiJ8I6IOFKIEkD9dhQcQPdu+N9MF55k15wYGWjkAY/VS9YE7l/PvAm
qFge7SACCItOHa4Qmmir5rhAPcfWrbe5JRFvdhuC5KoLDioBsn0jO6gtIoz7KalR
BXbtQncWXz0k5ETJYdi5nxY1KTV5sw4VYFuK5FMHeFomMsNKYkBgT18Wb71MxaXI
D4e+YxPYbec/2i7UlUTSBU1mgD0whk1lJicln8wmcWYwQiZL9UrKZrpYNARpykep
GRXu2ZR/tkR5341S2Ab4EswtsO/RRvp5FM1kSQYED/Gxxfv0M7vNTW8Hjl2y1zaz
u5f5tiuhlgFRuQWR+vmvEUe2e/uOgCXuuTHizDv1EI7QPk01Bg+5KsR6JQl3xuIu
33DUbMBOX2dcypU/HEujuT6EHaqd1QjejrREaKqB/Aiujndl4SdM6qTewccptTCX
ZC3lIOuTigmN3PVSisfHn4iOaFJLtph7dN1o9oj6o4QU+w/ZB18wjy+Npb0hqbO0
JcwHA6FEUkmGPCtiMCTIwUfTVAyVBLQOZCE6GDjriKTcvvscJHNy5KlUC3zWm9C5
61LSKYQw07uRat4LVdyzNljMUPo3HBUJ9r28eeWtdWZkZB1rlbFYWb7/DN+3kbIm
27NmP0VufsCjc7S0F03spQgkz2TvARvZQNPZYSNtbZ3pIlE/3L/REKI888Pb3Eea
lzu6ULXCiUkWzjtOPLwbB5yzNtkY946pU57NXUWNfgEVjEUFZCaHZDc83z3wym1t
pAmuoMEzcjm00RffCZOQEb6sqbt3zXvS29XCXqzOk6RnCq20jFHBHhlgh0QLIENj
N4HMiKUzE1qeWaC8AEzfYedBkBzdm+CoNO0r8U8H+WmBGHy0RUnvMjMN0yCy0v1H
6hyurUaw6U2+5heZIW9ve2ThUHHA1R4Z/dsHnA6DKwXvhYTbHQJklcua7eTzh8dt
IvZTIO+85zgcbfa4bDolbZbgV18ggde1PI3gBblU3heIpvEDX6dB590515Nft5V8
UK+jGq8mDmMx7ygYif4whAoc635eqSSuoffBRcfw3wkajd0+YhvtWkuSTZkcreQb
3NFAZXohZyXKaARsfRUT7xSTvqZrBKr0Lmp7pjVxgjC6gvJoFj6b9iHrKWG0cQGo
Afz7HDJXVJnpjdak3xh5NKjcRdHsP5MENy1g3ANm8EfX09Qyhm2Q0pTVQDOL4otM
lTM6pvPb9y6YtGg1FYCEUya3b2I4bFXX3TUUe/DYIsnGsaXo4PWiLYBYZtkoVSn7
H1whYQx+vo5zkyB17wk4ho4ll8UiVsNIZugVz6aLjyko6Pt9GhqxFUEFpiqQF1eI
Gtw1a2gJk6S5peNdcv+HolINucry23Bu7ZQtoMch8nfGuwcJUUUnxDc5AuErao/4
YL1cJEFpvAVZx7A8HnFC+jKUyr4MC8SLe95bNQFMEIyfHwhxeleFJKQyaXdfpK36
SfQUZzoJJkgYL9iATjuvHS538v/IYAuq5uDs+rwQD+rY6KHVq+2oa9WeM3aJF/X+
p7/iXh9wX4rTGZrGwsc23yo2+g0t2XXw980AGF4ofW8ZDpWVrO+H96mxls3npr0T
BET6nbOfBNcwY9MY9gSekoq+rUGuzQwKfIkA++p1B0q2DitBJ3dD9PhFDD6FMIy8
+qptxshxNjZnSM5ensPNjVlSBhx7Vn+ONLKjgTu6ZbDOy0HROL/IGf8OMUM4iyqP
28sSRRwUHw1gZNMeesAMSPVMX8Bo+ijXm/63PDD5YSvPO31jslIp8+kN5QDhe2Mb
72WDTn9H90Fw4f7tWA/60cIV/UyXKD4j0Vp0qg8Amg7U/DtpHYLUI8pwKfTmiZi+
pSlpm1UUGHXteAb3Uvt0n0ku8+76Rpg6ldqJAK5Byd8habUdiMP+728P1/mY3PVj
nib2WxB2lzLMKs0uxL3qFGZl5AeOMLZFc/c/CZunXObNzA2kmhbKGt0hktmWT2VB
FIModTU0kEyEEyK1zY3vzA7F9L30TJKKRBdeygsoDCAzQkreEgYMKMiMxQvnWb6Z
kIAp6ljNw7eYI+u2l/rHhs9PKCuRjWT+/ICkeeH/JimSelGSjfFJNE15q+u7CEsQ
xrc3ZN9dBSMMsKuhz9AxBe1N6LLhKJfqg8eGSVW1wkPUaQdV8cSYiYTKVG0AcTZT
hZy1OzaTQdxONwO/M/o++3+yTtXrn1zsi/Bv69kPVBu6GBLnsoERyZ1apZOMUpO+
FHaI06TIwTgUajZ2E8n/R9KNXSurq+k7jFyLJ/hbcx4Q0y2zakpG/A6gVwlqB/CQ
xk2VJ8G3ZhgWk1Udsoa9TxxdlPzFYOOar/4F+sF5sRIkKNfYLgYReFN8+Ssh2Jm7
xpU9c0Fe71n6yZsnUAfyvfkOodaJF3hHOwVpaR64sOssdf+71l6d/e1P0dmDuT3C
ll1qiy7m9hwtz2e6X0aN0/n0MhS9d1oOYzVeGCbuJr1+6NeN0wR3k8aCs7LnIqaC
65aHZZ6Z7W3po2A+1sgQuegTbP8MbQ9xUzDSEdrtb8WIXZgz+nu0zZTui//OuNUl
mLhXIGrcol1/4wU5QC6V68EuubnNkK7CX5yJtmTlUSFtswIH9VfGUO4oVHuKXEr7
uv0IA+iqT275FP8AbaPfN7Ic2YOP/Ct9F4CiWm7Ir8APqWqk5LoxXf+1ivj/hF2T
Ljkx2ij4PC1lDVYnePJxOQX+st9sO1nY2wFrlGBEEnqMDftHeTEKTb1zd7bMfJbv
zBnCNpemuXdEkGNMR+pY7GHlhGl0/Fr9w+syq8x5WiNIhyWqq3YvA1JssqVulKB3
p7gOMqC9uVGvW4C3wQpvXcjqOGVH0qT6lBTkKP3LIIJBg94mowaTH7MC9SUq5Trq
LFkgRfuq4hiT5UGav6d+rgZ0IfJfLiagDfRSUMbz9s/QJgg55rAD6t6++MZdlnDy
3i2MXTRJ22i4bMzzTBXx7kc6Mr0OAptwQ7lC1AFsCozdg2wb4itOhaBibwp0c2We
oDEcH/+RQwY/TJRjT7osFn/sOVsJF8opm3jORWPcyJyPXhnDJOab+esamESJjwFK
f9bLoDQyjL+XB+DH2+1SEYBhE+HhIqZ1oQWNA0ptJEkMGhyjC1yHdAHsGa9pfShA
Ff7CeRMQ1ShXxeucodFqIGgjA3tlOhAeAr0GGsxQzRlft3KmmYbt1TjY14hduirl
s2VL/sPTGn9UwMMYUwu85FE+gR6YyMJw7FnQ8YPlSUQ9qzvmxBWWpIVolDjUOOR8
R52PksCbhNLh5IPr0KVIW7yweYn6tthnUKoocWzOMcLEJhNE2MArQWmS7CekkRYm
scTpjcKrU2Kmj/ybQKuJU+0vNbbzQkggvRl1hfXDig/sNeR0nuaVw06yfg5u75wc
wAbBES9MOK+FggdxLeH7nkMc33WuZQn4S5kc6b4Y8YgdPNq+V2wh9U7dygoSp3Eu
oTNr9YG54isiGd7ji+oCrWSXZYcFUTfAn4nTcvQPvI55gg9ktENtkaJkeS0yjEZc
UACc8bpQYJvh3mRUi74ueFul3YsDAUeNiMWVZH0mmeoyyBQQ93aioaPrajxyEEyL
j2I341tU7l7F4aRJ4NQlusNOz8BIZM5vBlztNaNncMkvfwSjOSvw25jbrQBG43yw
O4ElV1dKvaHDkk8zF8so3A+kFqeh7IIHbLg6X89hF3p8ZUp4JloJk2h/huJOVFA5
zYtBrPKfUuyIgmqscP5FXVlxjQRjDK2I+HOq6EELfZze9bfLMyibzvUkG6zXHQLt
Jafc6jtU5w3yvecsr7BRlObAWwo9A2LZDJDWDsQAa+/rFSI2LVrvPStKFjqi432a
dVO6OKq7h/0umbmOK9WC17gAYvsp7g7GUNLdqAhWnkRL6dgWmo7r1HmOh/7W6V3I
y9yYMdQTQI6VLp6AdQxvvtE1o2EsZk7OFpk4YwTq1d3E/VWs8J8YiJAtjyTRNPxf
JkCskLWoUp4BMDpCGbzgg8ycMBahTlCKj836eIMLU4ylyuITD8PAGqlIUjM2DMjH
RA5u8aRrhZ1kCuqkUuY0hDRjkyK+WtahIIWSOXHaFeIREAQG0aATyezJhY4SXaSo
XbsiwVF0oxRBrW08kADdeO2LqutbAFuIrjlFUw4f1ZDkWTBMI4dCLysA58WASgPp
p7BJQ/7+Y+krgNFkaBkaxym52mx0fOda6ZHJFRL7ckjUtlnAuRhHlR1XPkV3o/BO
/rE65tqTnWlMBffsmxqdAxftE7pDyPeHZLiHGsL0XUHi80S23Eu/ktP0Xv2zGSzc
DqaZhkQGYqe7nAuGALsIvJkko0bI4gZ55RLSf9aT1deEPujp88G7flhq/59o6ET1
jDmhU0nb6Yc4sihapS+Yifgv/6f3XekWRt6IIAvPRA4dcnV8J97zh7swFJVYwYoA
mZ9khqXoMiwgUWlllUhUOzoTIlb9y67PknpBQpxURWf0SqfhVw63gEDYIku4Vv6h
QWhyiKJuvSWNeWlMylZXwkFWdBXWqpgHVbosCphvxxr4Yaew8n9LydeJEE0joan8
K57mDo1dbk6nJf5FhDveVQ4aZSJTHAWg0tjmMWcZSCQd8RGGISxjGBp+JFDMFs/0
c5kSCeuMWsfJZJ5MIUnA5G5ikNnfVBghdBSIz4ckc+KbbbYNJZPNtYFEmN9t4At4
T6s0BA6wdGDk2+p10363krN0rYIKK6j8jLUMbvl5D6bqsyWEYeQ7sNO7juUzLh23
0pRsa4nDUABGNzxjy+0lhmhbd/J6KL/76k800AvALjEUqjs10F2oSE7KdYa/VowB
iY2uqynDql3J9OgiWn0u6BxjhmHrh917EI9QTcKBRaPUHO6XZVaISr7Pep4SplKZ
QjWGzmPUN1VRKkcttCiMPi94brwXiwKkshCaFa9J9Ft5gIk+MdwVcBBGVdpzIqO/
FRhtbah2r5KEro7wRpqiDcZNNVBjEAhyDeoudd0Ipocg7bjJgFGkU+tx78DICgbq
AKJb3UZQpOZBpo226DT9ApCeZJB/x93bkJWGbcVj+eItikeF/YhJH3V9hOCVx1N0
kYTfV2x11Znw4n+6ZGs5x5MD6nX36iJvJGCjZ4ZafWhUwJqEOPir2bDNeNEVp//W
I52Fr3ZACX1M0UtC48xEZ2LTkgc3hp4kZ3petEh9bGu1EWNWv+50cBzx7jgMdDsN
MzV+s3o1P2hSuA+gWbNqEvpCXOTP3tEepnxabiDKpb9CDfTRnbVikZdfcbgbMTXa
pVAAA1AA+RRrsEXwy3T/sETJMlQKXJGitP76cKnnb/BShww4zNBVTqKhpMcq1Hq3
4KV9Jsenz2TfSuHgac5Kjg0M2PMNjdXgyWtrbaISRnccnbFLfWm3Ytz8g3fQBJkp
/7Bzbop+twEJMqC0DP0mkgP0czFroX5a9dLvFCcgPEDyosCelXvKYkljKi5LyWH5
8HjJMSN2SmuY9s6EAYVqg4UMWztKBrNf2MwaCuByDeAaEGb0LaLR/FlhuNI7dY4H
KmoxQky5y0hbdYpGJSGHj1oLGAVXKjmNj3NfV22r5pBZNy2AAKUK4ah7xTYPeXpV
NF1EiWO6mAPV6T/g3OnuGXqfB6/jkH2a4MDV+ypLNN47WrdSjl31GoRC58trDyE5
AoYagCZwNAqPB8rEMk2ev5D8h0NbdXhifhCZCocY2SmlPJAHD4NicGbPhNaw2QCI
+3txXZDCYD9vc09jIcvOz/uADvuQoVK2NX5WPizljsI1keXRdJhyDvcCxvBeOhWH
idYNgxDFN+fbFK1+Bav30ThrjnAgfi8iuxqEemmp9ZyvCl/j/LEUAw6RemVXrB42
lD56vNlkyuhV84t4sKLMtfUzCer2Bdb/55Z/74WqxRt1vrgzhU9a0TUdZfe5zrIQ
s0mmWMP3Oq832XhXSq36LHZBJH8eoySLWBZANEyBzsKnKRR7OFTJ8eU2ut5Y9t57
5bdQeOeltwl4GSSdc8a9hvzIILbOWwz5hZj+gvQ8QC9odJxiq4aYirookv/2NTU4
h7ZyIU+/PP2bjUx/5/5vBZeiJTolJSkDAj0giQXiP375y57McTShUoFVa9hvOb3O
49VsnFKv0tg1ahO5WIINzSAV8rbQAx7oI5S5Tgaok3er286rVfi2bsOPygW6r4Sz
5huXk+9Krry71smQe6gC3jLEVm33liIhQFjt0LKVIkk95ned066Hoa+EGc0HfnuW
IRns45cmPhJ+ACNb1LtpAnIKMZjkVCLhbtp6Yz8WXjKVWQ6HgIBiQJ97wT9g19/7
8DFQxP+66GubU3xaoPFhhhQ/TrQCUiOHTxnoD928QOMqkR59JOTBifR36KsQjFDS
gz+7rmxN5NyRKtFC+Xl7Pt/9jcLWkS4Pl/MbhoH9ITF+XCxr9DynR8c5EaP3Bd9R
4izFkQxaMusCsg0Wi0Q2F2R+RkzSra1t/kwjsmeRjNCsA61sawqnO71QpFSzFyoy
2vd5Nr1hvdPMFRUdDE7UGPpMr10S3YZxMa7lZNogOIKO9X7J7SCS7ym+L712ysPs
z7ye5b3kORyLTv9SaNbIs5rOJ80aFzt1i3iLHieoqdsa34rHuEfGZf7Gydv6mYC/
1gax5+0Tvsa9p+GR9DHa0THrA75gEmsIf4fNE/HwB9JQPupOmBHeNUxApLyitrXJ
GEo2H43StjNnth7Pn2AjCiy4vsx2nUgoHTWzs5sMVaeioxrBE2mfo9onvgq6YgSh
pfYf8dGWqxEamhnRt4ZMPgyIeTNRpH/5Y1uuBH2TfIK6UHGy1dnFozNK+tOMqvnB
dq1p4Qexovxs64OuVXSm24Kg+43EmvaKxeIvhmhDGfWdMJ3Tf1hRKgSkEWdNaZ98
qGkYCVRwj0ox/1xCvQjVTQw+VA0bijsJIQVCeXKNoo3oB/F+BI+axq6wYdh+0+2j
1KuTIWTFAuaWP3mRliRo7z74Obj8qCxMcQvEbieSiLcGKeeApfPQ3/FNcNloQTQJ
yl//xtRot84z+B6kZGHz4CRidgGZ1sbMcFt+tR7hswOf0vzp9GpJXe8eETDUOK/N
IYqaK4Obvgwy8x86qFMmKALPVPJzJxHVAjx2WssYa/DAEYQBZR4FOJh1Pu50gUv4
cSalGpmNH1mvze5H5Z6nZM0uoODHzO/aEgDb/+/NeUMQi6WJy0AJ8Y1Rm+b8z1AU
u3Xf/I9UTMo74ZmT8GIgMBPapePdiFSfNzlUmMcNl3ME/tTqJsh4+m1sM9I68CNa
TtiZ9G7JJ7fDtU5Ue8xC3Uo4tyUlOKJXsc6O3kaCxcEsLLWo1yNSyyu06/Tqu5VM
ngCoD1PKwgCVsjrvpC4EA343nc9toCGKryy886LjIGtbLEkaqYmz+TnZc7AN7mYS
d7xDXJjUnHsMI7vYX2+3+3ApKt9wcyN8aPAPMorSUG1JtQGJtyna27b5evmbv7jD
ha7UQUoEEAN3tqI/cCG795gMWBrRVA9fdeRp/IfnX7NkP3+Loc6uVdLKu1qZ6SIL
8wo8ffYsfjqHrcQvf22OmC9nwc9/LtDNhsrs+gyLT4Ax5ntEi6aQzmgSo534mkJW
A1Eg/N1wflh8fZK9Zx+DhKCRtVTwmRzihedsNTiPkj4AVgBsOsCqmXWluN/tjuGw
GK/je+vZSTMroFszMGKi4SHFOa4lBcPARspd60P7pTnGzw0skRIuc1K821OllsbY
11sl91wZUJOouF63twYd13xE9T2S+xzJxRnco1XMPA6+YyP0kKrRUNZmAzT1cWvh
y2lWFC1I3sv7zSvtt0zPgDiK8SVQdRMokIckq2QmGyPENZT1rUUkEn2CKxpOtmNX
lFIlNhlCwwl+dpLpPjdiPavRmhS0yQ89RNGdUwXBGntTZ/2PFHw2jD2Nfef4gKyI
8ZXsDa4om1pkiVY/00Wkd6LgzVHS48jZZ1deoUmotWMeein1rNebCq3Xm5LXHgVh
K0iUtNAKvOqL2AAtYjIlZov4sxGlgHFXKS3PsrwEQAgcHA0PcL42n5mcduGPIf78
TFDfclOZoAH9HDuQVCUYSpgAB8i2uqT3n8PuW4noto7E4G3b9UpRy/FEdiFftNCZ
o1veeCsOoC/Y62E9vfuyUW960XBflk17+4yTesVbfEpOuY7fEco/wWkTK9JbLIu6
8ArGXMGv/PW5Vg6kstcbM8RPBgOkXm+MmTeAtY+BKbOozQYo8xv2ST/OUYdy8lG7
Q9K8IdF07ax6TE2SHlpEkYys7VIpZardTD8R8PnIMbMJjVbImbpZt5K7bxjgd6lT
u0y3Q5Cken7OvwZm2aRHBr3CNQC4uqB13DRMG0v6YF959l9vuvQaVw1FnCEqEe2e
LdWgFGh6WKSTgnqz6ZnlNMCKT1l78wCg4xo2YY6gAkmuFi9/IkGh03inuVdXMh3q
FIh+ZNKvmqV2E8SCdVWfA9DgRZrMfpQE8mog6uSzY2X7wMEL4ItzBGVt294B86sw
hj6tci0rZ/KSXxlxSDjaJ3ld5qN/6Ut0C6/8HAtjC9sfP8/BCK5GJxJZfonDTyl7
dNrjfACsSkvO0rdE9hB4XN02iWLBBC5k6hyNVPR6igOpEnwJQ5VfvTl1fGWAA8iD
9rui10YXNGRkG0DxxwCR9gn8rDyFzSQjSY5XZdZwORWCJ2D/h6JolLiI3I1bA3HH
/BJRX7pcA39F+J3aur33dplnyu/BjwDnscJ2P8T4oom7PVQPJ0Yg+KDZReDvHORE
pTLWIhHsAuJNJAhCeZsmRl0ir6bwYzS8oef0JpTKekoWFIU4QUTGdnVCeutsKlsF
9ohk73wHKVeb4s+wSZYC+gTbVJ2tJCgUZzgid0RfJ0TmuF0p1WG/1R0Yh70KQH8u
C9b+7fMNXvOPDL4fuXBKznYzml2N60eFitZ13efZUrbRr6veQT3hOr1PLiggPvzI
3j5clk6mw+d8pYvcjRNvxwCGwMxgA8W+wlwLyILzzQW/ipBUs7GUFaUYUNr/0iHW
tghiB3FUfLgSD+jDvg+kPrGLMW6V0qMSumbFWkPfqshlLz+whCEfEV1IPs7w0jyI
ME2XMy3/0ZjFAMIk7gwBSNIjNBfUAkcbtvDhXA45+vTvspIo1BRneE8xWIo3d38w
7/X70cMXjUVsR2FLN0U64j+xA+jL8AtIC7OcciVFcLn1IkyOj1wNv3JcQr/GwcFR
/wMOCwCyT0iRvzWjwxuY0MQ7XKm66s+H98Td9PThOh2ifQFR2jqbm76dQtmwL1fk
LZ1khrppaWF2LX+TBvBXaGIzCsBoMdEhkxh5wH+40UrcHtStDPmQqTIopkcpFvCE
bV0Fg+aMYR+i/tAf6YM2RsH7mSPCFrCRko+jcsYy0vG6ok8NKC+m1Anpj7OG66/4
FsKUe4xa9j/QAv9m6yJmYeSXJn30i+wcyxTTwn0OO8cBnh2mYHzeP4TSG92dc/ML
J9iBaNhJPYafZvAi/PUbdpfKp34ScJhwTVYUTB2kSfqTT4KZ1Eyn1I2JS5HNh1Nm
MRtq6quGxg15gzJ7SGNK49tjut9K9FyEZRqVJJI+/6ajfB0Jyz6GdNR4PxpMcS1O
oQpR17a+hf58NVEaVRO0jybjJZsMO5rloNJE17kXGOMQgdCErCZDb7CqS5KSMZDF
YZp/FRLm1wam+JawtNtctAaN6QkrarMpU7Ly4Eo4va9xAlspHpwf/8A8qEVfTkJ8
k+O6OVQ4UTYJeKH5h4Z1bBdLVMi2d5ONWMXVuJQI9oxrHiIGGabHuA8lJoruwhYY
8WomQEYrRfAAdvI8WIObMy72201mECufONNvcEjzTZfGBWBJkSlw2lDjfInf2/QT
KuXQTBDcJAdUGHpAK3+3g8X0Uc1VplaNIMgdo+tpxeSwVqOYhCMMtmJnwr8F8AeX
BUgwQL7COZ+QVtBnXVYSt6KvGaWuurWOiO+v1zyHvLuF+nN7j3F0BsbYBx7Hma27
gmXUu48WXEIhlMcNtYGfPDqsTsknk8/5evr30sGIY+IzS0Uo7bMKWcgpjQG0PRej
yFzfWAigsjxfzFcM7TrV/uD7iPwmg6Udpd9oX1BVStMQvi/xv7upv3+dX/uw6P+x
ieRf1SClZlBtdWgiv+IIpvDb3YK/sOqxlLQaqOP7nK+o8ZZJmOB65wQ766TtuLKn
mHM1PDD0VOL6XVttNX35fe1fYtoqoKsDlmoTG4C+f+8IV1dh1xuhlyRqaT/C8/Ox
/CiyRjnKYW9bgB4svI1Zal61d4/48bdTsYZXwAEU0PAcYItP1K+p2HZ/JtDifVjF
n6k3NHPwUj1fqWMTZF+6W6ITCbBTBQiGV28LWG34iHT7Prr76xGFQpCHczCOYRZQ
d39IMwonIj5GHzhBnsst2WZOqilHRisBX6xbvB0UTo5at6i8SoEaTt/2S4NxhQSB
SJThlgczkJsp7hR2rX2EbTXnmKtIin0n0Jm6rufPUcoA/tq5//XR+e/oxAEO13Qb
Jg/eW0HdQJOnCYSHJKWE4c1a/UPmQJ8RmzXsaKGhaFzdUl1FBXqRe9aHFmFmRFZp
N/0UN3h63q6eD1Lggz4FjS6Rc9o4rBMvfULFPDAsf6sM0DPDQv6R5+Z7fDLV5ZCK
ioJaTR9TW541ZGd037fDJPK5EQFB9FORkf1YvdAMch4NxpcKeCPt/aQqgj/gAm+z
CSVOz7vbjnwYHX68bxhbUdR/HxrmP0LfONrtnLD1Z07RbjNuFteVH6vrgvGvLDB3
GXKyiWDrdsha5y/dwj6WIUUgrQe4kq1If4mlBZJokkdf5w+6gk5s2fv8BO0Zx89c
lnTSIhhWYOAQD0lmCvr16dAZ6bFi/2YVazPVikYTgkiNF6HgKjsTm+voGu/Yb9NT
UI0RdmNi9WpdNolescq6gDQHr6V1CDINfKMWZz4cvvAP8T0KMtCCVlr3UOjTAdcN
0yyhZJMdDrdi+aqne8L7sg6RmxLEBtcLrk1Cvm5imxUvgorSaMfa8vCMFPJHCST/
4xxMc4UWNL+o+nH7bwmmLxVTU5Bvt+MOoZ2RoZHuSw0ulS2sKFCXgn8JPPXdE9UQ
pxBuIdsMDv6liAg4mtlcHnruQ4RxdxzZE1QXjmiLPn9n1CbjMGlpBqL1x8hhTq3C
8HgkOBhNye4XcJ0ptZ9Bxkm89xRRibB9KZR14w4MARcF50dfw+LlSJXW7DYkI41s
ofxOiWs7xkXdmN/aAMFa41aqtytp1uqLTPTtJ0f0mC+RQ4qnT/nItSax4BU+DdD3
jm/2xSYCihOUprT2bYI5H5tmcNGrd38fEJukBYhc0rwGY68dwi8OK35so+Q5AcNa
2UVYvsWtYhltLjv8q7TepmBE8ULsnuINd39CjrEQ1au/wKjxbvxltGAV/9CYVz4Q
RP+l5VG0Us8NHCh5RwigkvGjS4pqk32Omr9wjGItI1HLxWX83sP/ukVKDDhC3bvk
7/Hg03NsUMYmSwlSz1QwVGPVOe02j2+wwcgxOUCcynVoX90iQrhM9oYS7g2hJoYn
UNk2wIAlvMBmgfQhOlQeoQG6M5r2uJvSHi4/RxUOipWYrp7jaUaOOvxHC6y9qkuW
EMqej8YpflIhT31fIGy0cqRHL0cQ+IZcB9tkN/l/vE2wCsweYy7omMwuNRMmwvLP
xyFGBSc77fH5xTHZSdv/aDbkZF1RwS5r10DdDTfGP4tWJTGLcXdIXkBsVC6XqVvp
MYRs8JRM9iJQDMXLrbFFuyQpJcaEpoLL8of4TarQ+mCg3tSQxc66+o/zgio4aLxq
Di3RVtf9lVyD8d0KhotH3DTsE6woqll1zX8r+7r1Z85SIGYeHq4KOI2U3an63Zee
3HyHYwwO6CnDdJJKeD7kH1FhnzKP5xNC6PyjiMM/14B33mIbI6GpQSXZqfJiUfJ3
wrZ2MoQkMjqfDygoMCBcRaQ+PrVzJUFys4qD83jjlxvgCVc8ECa7DlO0k578gh3v
vn5PBwrl6nz2GnAgiDRmdFdSDmjyCZPuSj/Ik1MUGn663ZdSc0C2Eoy3Wr2XYdas
mhjRCoclOk3uJ6TOh147onhcMmX0SEAZHbR2D8Czr0lXX2DVwTKBoani+6iKospD
YwlQgu9gXgVcq/a91eLOXTOHdPrB1dBTeZ1hwnviSndw5wLFB1BerC37VX4GPnL4
XaxoQsafU3jzsV8rM+xfvRpJAEQK+/vEziBux/YYob44dZc01uQDpa5l7uMbktyq
e10ioyHzwNf2xLFf6rRCNVPvEhR+SAvDNgnA+55Sqg0iMGvrMJZi8iE4N1X8/vGL
Ql7T2MtFIwtce2Go1GAZN3mzCEopUfGg8Urt12V2prSzSGG248Bc7mTbv5/3MQGa
37ywpv0BzmBbAobYVS1h8jRphipnur1CZBV2Yspg/PFdmIsHGzzTYVO32rIj1H5s
GtYIR/+qxDzBEQJpozS1Qnd9y8j1Ek/FjQQFnHM2qptoTVCVO2gXd1NH+6r88znJ
mEOOs/Bmf6M8rCwqt0EPlSzuMd4Kr6Puyn6bnyJAz8Z+nohwiftyck/Qcj0aO8iS
2s5BrnO2yBUQPSGVat/CqkmqkK7YavhhmQDgPEzV2vC2lU/47lI9Ka8DC9qDnlaC
YPyTR0vBRcrmanD9VC7NRFmn5fzaUbXKc6DtA6H3YpXWXjAOL6QZcSr0hQy5L6f4
P3YXR7pvkHMOtlIrjneISnoLPbxxRyNqnoxMvfLDcZMaKbWwL/l6gLiGqoCFYziB
3JXF777El6BLg2wyuOF/WuKye8Srm55qGfOZnEYUNOnMJLvwziRFSUsc9YIOQawJ
DmPPpC4YG4tZUrnVLT9ujsxqidVT2wuVPYr56E+UN5W+M3FtDJUvbreKz6M2xIWg
MBBVLMeDFzqNnc08DbW1U/uS5WcJcxbZYqiIdnY9zrvT/wtahnwTJSVOi+PCFxch
ZjPZhCrRHBqNI8G9YSvRBscQAg99opHEXR4mL+T2P2W/DUc3igKen2SFBzgAcLNf
vhApKL1xU1r1mrCXuXcDI9ye4qQ51YQ/88+4HKvlu4NfQfAI0Qd0011EmqGN9FzO
dneQlXoOMpoN/tegcq45TKxmNkq6RFLPFzhuDp3NVriER5Exk3xp3U33lSL9/eqI
GlP1cZEoWHqbOOgQH4/EIQ5jXAWtvyQBsayyVhCvX4eNQ5PC1D0NtpBUThmJJ8Qq
ZtdZlcLdxIckeYxivYN3ofnWCuWVy+VTnwta+WiuHbsLfdpE2bRRSmEyH4yaOAWr
W2akyJ5N40sLehimpqfbFeXkmLfSfkY2g/sVOAo8s4g2zxHLlnyLsth4XHkGOd/V
YXoVBfgscU9g4tuCd+Aedlt+uGdKq7VezuqR0zsPfYOG4rFuZaRtZ1SXSitulg1c
nCi0KnaUva0gKCA3r6F72Fx5aeFzscgIdr1SuWOfytBvQhbF+nhaxCsff/8XCdUG
QpFHvLOx6EQBVZqryt3OjKWHD3gpeMrzOlJfUmwmF+U8+1OmFrW4Z+jitZtXNgrd
198vXhowmkQ0lfiXQ0mhoCxd1jbqMM9qdYHaTGBUk7xmbQ8HuVIgeDFCjxE5cdec
CtH6rrV2blBtn0sJ0Iax5wl6UgGILifFf3B0Nk2mERiBWeOa+Y1Tolqs2cxTUTjk
1Y/hPNQXZsPn3ilj64fIzpKza13hPA86TJP8+jhrfGCPicHhQ9ZEs2sb3W3I/IvO
Xwldqd7xJm7uZbwXUhwbRgsJEIUZIqi/qcXuIVthi2l93nLp1cSySM40l3RJruPf
jIG6dpx75uKkmRGsNaFYtG9JpgLEmPci1HJqDEEywMhSzoyVuVEkA3DMSiRMRLgo
0N2F7jleyG03KMbgsNcsbYUGnHmYpQjvVftheSOIAypeAvCIPLWqVUbrK1HZAYu6
2Ld0nQX+E4admJNqXv/sKh1xRL8yuv4ylRLaOCYEckgzz333ISXohj9NJIDqXCYt
UqMNF1i9YiJmvcgrymPKGAb722sUboCT7yQxaaAcf1n9nSqnY6dzwuUz8llOWeQy
2aLeadyuAA04n8RiPGO9iez5sC+g4Q9BFF/RV6a44W41QhNiLg5w/WCnNrvIJFrr
J0+s8lEbjKL6myL1Q8Ib9AglChXHV8bZhPhQxUmtW+HbSurYPt/+czDLho36lI5O
SPcyyKUT5tTbbEXWMtqm+srVScDbb2MwSkmrTYYj/vhCTjnBLiyCZIDAEEekWFS3
YP3SE47hcTbfV84p87fWOYogNZ9YxU9KDfSkdi7uJTnpdCfnoHvqJHxEzul8btv0
55QilOIQ+u0SM8QtYf2P3Sej6R1s3TdU9nZbND60z3l9FXE493nkl51ngbyucz2A
sLT0bLekZXIrAEcVYwNk2boE5VLb2j+IUJRMmTsinfZRxXVKC1kRK9+tQ1mMCx1l
5+rV90EhaYVaKIPzCghL7pGtqEwNXmoAHvzjIuMWHmSqlqjKKTZIM4YTarV52xLW
wUQObP64NY314zlOlVJwXF1hwUNYwVU8t9JGhWDWq3Znq/v0fBviKd3G2TNbMhqE
FPQnOk/KL4MNyLbJrC1L+z0327wo8blO2n3xWgOK9I97bH4J69Ylqvha14maDro0
1WlOmIb7bpkkjDmpWBxLcfg8PLKPdEM1Rsb11/Qp8vx28n2MmXhklQEsoKNBGdz2
91kdpZXv+OzDy5YIHSyOF677JVOIZ36e6oW+a9OJbsdQ6PWBER5RYaeYsM2ej1M6
q0x6x1/EK+vWylLBI44DlTnBp//wQWbfKAiV2Zan6d2N2upTSyl3MPMNivzCTGaW
QmIkhxcmtSGSioYgtaoFfn9xLfS4ZidVg+wMO+jKO+GkKw1LCYIh70dxJ10F7TgR
qf4NYOJDylWtsAgvAF5m+254nRD4kn54UxLnIMEF4ftu8YfxeR4hbHPn43xjW8fP
s3XbKQ/INo8fRryaxftDLJFx7ZETuEedAGMCNGYjjPDbJFejx+Flk1OHRvtEystl
qRNgdNxMBAFRliuCq6HHO3+99dJXowUili6FPc31+NLnW7f6dB5v2nbKd4Cf5/s8
JQOMOrdTJco8Daw5/hQkL1G8tACnog6jjRPY6pqW1YZO1XH6PGwjNBoFT12NeyyU
NU7QFbaUASqFoAbQdApyLRFHyZnuXSTo8BFU82NybX/9u2cxPVFWm3JwrFkvH+VB
uL4XKD5WFEcv5YkIycywZ/9/tTE7Ky1YISrq08YARfK2Af+VXxNNFRMMzkyqJU2y
/IsPZOmFwbVzPKiqQZzi0q0ynOi0spyV7qGD9L/LtcjkmTb7sV3zR4odxqxABMaR
lfrruRKRaDoiH4OjulIBFz+jgWtS+F6plKFSZDWJUIvCJaBKWLrhhmV8eOoSCqZ1
dssivdVwtJFDOXDqbE0kZ8IIfWaItBUdK7WlOTvcmjU+hkZv53EKX7Pj1kDBTXc/
O5i8QqqLHcebczS6mZBkZS/mAxWk9h4+9cF8aoG7AfvrCpEjTIiuucaSCaNZGibS
7wUvEEDNtj5oCIfD+33Fwi0Ky6xEMj+n35BuMLp+5X22W3f08TVCtIX2OxVjD8Yq
WvVGu/lR1/+EajVGX9oo9Q28U4jJO4t4a7OJEtZzdUq5apwRbGjH8o7/rdY7Zpr/
Ak/AOLzSt78sCdyPNftX0hdZa8ctzly4k971PNpw+95e5mQDZhvGiYEi8S2a2QvK
1QfeWw8/BZoWELWGyOmvaT+xIDGV+g4i+uKPA1zCqqCffDQwmoNSMMJizdr5Gc3d
Jm480cJaVP7uPri4toNN9/o/f8YhZZ9TtEzqJh7NP0zQNxvL2V149FDRM7+ix78J
40N79kCIKXMO8+lKbLSRrKWYprNidNw40UxfNU+e0hnMdHPJ5Upz527ccAi17r/8
hM+4TH7EsTW3iCbInIRsiAtoPizVHo8L9P0BE9BHveb4VrjaowNKpv7bMwoTd6U2
00VXMkUZahwxr1IBsnxw41WXGYt9K8Ly778EHf5nz4/Ap4YU7fIdzXNKIYtT7u8g
AWff5NuqMPwd6wbpGwQ76pSadgMTZtO4MaCYrFIJj/J80HesfNNeDVwdIF13fk2+
TOt+1nswVfzTelQ6KdmZv5envJHcwABKZLdb4vnLt12EbyIdHVV7dGJQBI+akoK7
t8uiP8uGgWUL6l14ScTmkqoi8VE1aq8TcdsbS8TD8GHa6rgSOhzEWIsd/PkVjqg1
s30QLkoYQf9aPeGGq8c73+3rR+XpKJ+52Oue+XjFZVoORpjL0cZ+L/Balf79ZYRu
DRobkpT3AlNpCcUx48ISKBQpWPvggeu7b5XmwlAdJAt9KuSTpGAlqJtiy6lZMTAc
DfdK592L+iteQ1iOZjoXzYWhgGpOKt3C/OJ4f5G21guHfTZl/vos3/PQsGOPgTsl
USCaJ3UHCZXlYhjyGB6xqJKxgj3lIDrAIzCMU34lvevHxWtXbLUuz8BDSeoRONjR
mizh/UuZwQZnibTUmvrx14vtGzeTW2OcB0wQQ0A/I3gUP1qxpHNArvF2OOv8PGla
638BB/hWLMAvi0Fgy2xPFrniK63F0F/9HoOpTPvrPFV4R650YVHyal8THCyD4UeA
+4TH/9CyX3jmHVMqhdYafhbuiHFLfbZFwiUrR3hOqddXeScdJbf1ZAkAXf0Dah9a
JBtyjwGsQuggDukZJECFNtMqUurld4B0hhY9KRk56XEO6gs3l5Jf9gcEUdK9hnR4
BQ+n5tB7Qcs9mKetPPQqI557H6+WXBoAJAYs1p00qDszgqYdMYbU2mN2Mbg3GviX
QGwRQ0E4Jguu9UUuT2DKKbLwlPhHSUe0bz0FB2pKck2KuJavXRNSPot+h+aNuPRB
c2xbIAg0M22e4yHv8BDBAlB6IcYL7IM8HYVa8x9s5tlVZiq57B4FQH1P3M8//4cf
ZMoNot3xkeTNwRxkfPgXXwlY8sydl8VrjKTJbY2GZECmZKRGPeLi9x+CijZd/gJG
tX3qffaV803sRlMJmw8LTOpAd973npuAFKa1UI2GTVGWFSzjafKIqjARot1VxzjR
4rcIDTXHDS/lg4nLsfkrKNTPWpNMo3oNZkIEUrctLfbY6nHRTrLm6sI9iJG4VdyL
FXNHb65MbOrGI1pCUq77+Z9Y4DmpIGvqT+BgDw/301sv7MAUpH8I1B5DX4KUvCyU
YrjsgNwHxF/pRXzhKA/lNQoaN++4J8cwNePho4+NiydAVdIahs8dhpmR8GSvdRM1
OJM99f07hc3EhSnPp+W4GA5CEjBVsxX9u2BP5l2Xj8ymbG9ThadQVsaekw7BQFXL
Ny/sUWUgDgxwRZnri69rMU2ifra7PxZSc4UPdvp2xaykpjpKQetxEO2U/yKlxm0u
Sbcd79NOl8G0bUN6U1oGfqqEh5N7lx7tOpWd4BJiEzA3wkSpO10UVf1BAA32Q5h6
O3FozCQzbRPICUoTiGf8cGcQQV6pfUQ06+OUEgl1g0zspoAPH/kjAxbWAAyUt/Hc
fA1Ca1EDWz/elmY9KLVZY2kVe3CUZ/VJQX3pXLkDZwKq3YSNpx7DbizK+9sZMzws
b8Ag4dTNNqu1eQxfFyotks3EA17mi2CncZTwFwmi6haKeX8uy4O5sFvq803CbL7c
TaFLSrbqDY/XGzvAEj8HweFAkWpPr6bIVaWbyVNSpIl01wL75N4B8Fu13AFQJE29
irCJb7kl60gX4UOAFkndZToqNl6stnsR4fw9ZPxXcBrICEgPdXObVKdfM1Qn5wK0
yyZRwFAYNUWljpNXq8SqctPyX9A9xIApzjBJmLu6zYWc0jwxNwhcYYQM50GmDAaa
LOgPL/TDeYyl3XPcB6xXAKmsyEB88hixdRKzWX06/kOMCN/AiAbLhYv3+nN3SmTD
26YfiX6PP14+MbvvvndKQFwsbb6tPGoiK6BRlv3e+Ec29V9M7rnUFSyQTbWkO+0j
dixGXoXAB8zY98K3BcJu8BtyPCRuvKhKFaRBcKf2siqA2xOXMGPlGO3ffQ0QWfQt
HULK8XECTLAhqqOIPZeJ/KGeVbBBbDAbwT+1WFCBlNybywA68icbUTPIyTSDBORD
ory3NQllHIPJvufUiqoxjY0W3dD1nKLtKiMwjozxDzyOxoU6IasCoKZ9ZmihrBis
yvz6lboQlYhvF4AM+bzXYsAsIH/yvESW8Lk6k4O12A4xDzeqYovbSw04jU22uXG/
tZb6WVmQn4gIZiqJ1Vt5bZ52ore8CP7tBgKazUFsjmFx+nelrnFg06FaM6AVfzDj
Niy+mikV7qjnIx105zoUphbCzA569qLiDbfGe27gxZ68yDsvD1QJVQmMLfgmU7k2
Tm8Y1waI8cOHYx8tKXWPNcrUPdJSqFcF6/sOJ6PinXGSK3CL92ZYKIIrf/wuikSW
g8f2tD9Piflr1fk+OdHzU0VRrPw4u9tUAXxx3kUFamJ1uNN7wkU6VyaVKQVCYIfs
ZXeXXr1EB1jsZgibQAQLXpRLq6CMYOp8puhGm4jsVDECJHGBJI7oQ0QSsoI2Su3v
BdJo8ESV6UcM6ZUF43/VO3LTMxuysJXhohdMvN7MkbEQItNwRrYoubW2pthB5Iro
THDPpuBz9Mv6DMvL7Y90YBruBMibl91RaItUTL42jkYlo38vHj5U+DOBeg9i6Xwb
7RYRjbtCZf4oQrpi3hmQJlYp6DlOKuUbQa8qM8V16TNS6aCirDXgbg/BGUXW2uCr
klu4IwPaEAeN1eRKFNct1+klzXnQLElWOqxcUXEaWhV1tLDZnlJ7GM9VP0nt5MDz
Sf9qt19ApWNcTEtFK9wBN2p1NiFeZRLshatFSBVRE96AxvUj9H0Cww/o2pvtW9Ft
hWafxwZrEIZVQOI0RrSva0cECp6/nn5An1NIXIq1cJnX/ORldL5xMiTN8BGiG9Dx
akKsOcXKywkm/EeSYLMQ5f/Ahp4AYc5l7YGKLFO9I+y0uLCDvZlbB95b+C3IJG79
c+7/df/ZxTGUyxoBrRAq9sPth7Z0XPDDqOQlwApwCozVR74yWNtl3qHRSFOjGYba
oLYo6CzAZnzil02LMomh7Dh+HCKKAVd1JWSnn02kmUEfOne59HEo09h+aASuBv0D
uIQfSkf2Y0PgbFuAe+5jw+O329L+TiP/Ki/Vn1eoEBG8zgdJ95llOE9bQw9DAJg1
dCnxLEunvdJtx3jNg/OPPUwg6SdIeOTbZL+SVUgqqe4gAnWNIyW/V+V2rgJ2+r8m
YFW6MYQM8Fq4CRh+cT8krDMEoq/TatWpPFpzoIeTdNTa7xk70qJacYuNZ58DK687
ygc8t59difDN25DG78sTdLl5MNk4iEMwkKcFK4gTW+YQg4OP/4JEOJ+UaQMvHUf6
WGLvVtAgJf2JU4rZglajP6LuZ8q4ih4Khpv7OAmHk3k0DQJakYXprlUj+zOy8Xbt
1+iJxIm9UPnHoMRf1QZpURbw6RbaQ676zqJfNfuazBPrpV1lY1P2RvNREPs5jnyT
HrXvYREyRJ93rOcgura6PwJBx95t2YAEpdltDr8MB1A4uVQR6h+Sv80fHfulGfPG
IEr+ln65WCOVDgMEhMtkso/d4HDU3BZKmPcW32vVll4kcTCedLhDUvw+uQ5f9slL
gQDLT/pCO3ExzxAutIbT9jWHzC03XEpmB5lCcnV21ikI5K/SreeUD7LRXZ7Xm0Fn
NLyuoqLT7FxPPueA5dRcI1wwxeERqUaDELJ6SkranUcAGhYhWN4I6dwXfKYOcJBr
NiMKPl5wR8WhEyeJy777r0CoeNWcE1otJ6feVbV+LBpwI9MvkLJ93dDo1bnmlTXs
9U6Yrnq+qJ9de7+GUxM+0cWk1VSPKOL5zPbjjSJDBED+Qfy1L9BroC6I6Hg9AhNe
BYkpPeb+/uJz4vUfpW1gO3lywVxC0Xe5I2bPgtWkPKe0yZS0J0I7BNYD6w2htQJZ
pqZOfAsgeat9IUbK1PNRxpx20MPEZeMOT5LsVD7bjbc4NZkWwX5WlaaeSI/4YTg2
KRO4OAqE8SJs3Ubq/2IMCahbMwgKx6C7nsb/qexuYu/+2ZnPutvGoxf9fdVj/0fg
/ItKTcCuDt9z7iYaXjCLSm2bZgr4xLR6sXrPFJGs+x2hevhGFRNuoksTlg7AHlPw
8mRJ30j3vjdZKeAxnkcN1sxilz8QpsxoRpJY7WQEih1Z1sSPv2ilWP0qKzx2z0oB
BM5dvacr3CnjZumRYFtaAhmLnGfPKIvuKn78L5b0xejbOXIP1q5+9UZ4HEcdeSlE
zcbPA3I4rq0HiWr3UqZknx9p7fHo0mcLOyH34BjB6SBKuKBcFXwEhWh/n6GzMLt4
DoIb7KtTtkPrvC2eVmJ6hG/JuF553UxYqtEkru2xfv4xkbOzHUKZA6gC/g26JhcH
5NqPcuT7pMapFhtvTGogi3GD6ZjItEJsEs8+26Dy/HFM55mF/jp5MjW+b+W0BRUY
dHZV1npp5/sxXyl3ncceCoQNb/cZoauxmOWm7Z4Ai9EorJG06NBVITv7lk8qF0MB
CPK0pFuqw/v+c1Y8JuOIOrCbfS7EksgGIr05OyR7ayxRUiJkQX9MT/rqQpAxiS3M
PQ+eCbqHz3mWr7xBy7QfRBPXK0QefdXjrUe+e62Y7WazGYFhcQsUjvoo798cD7rc
5CE5cE4YliGCZcwOLl3ZEMp4UblG0BkpS2n+nbO7s3DtOXhOtSUCmgKqcSLV3YE3
/f0BkEOcxRcAKCTqDk+UxupOcUJKt5HVrrWbma0rO+JzUZLZCRdggEfuNpo8+SBJ
sFJ3tIvufrrlhx/yiP7avmtlDLlYy3Opmjlu/yc6yKdBV4oIDj0dyyUMumgcmWyV
n4Nv1paO8OIes2e1ro9SAOYnFrAZvoFpKwGPmYGQJexWI4yNZV9s/OU4nqMMVYZS
290Qt61Vu7kHHK4dt5se+tEDmZQqKwzdOcTloPkebZFZgV7QDYh+wQ9s2e8hO/ei
luE/PbKs1TeHrT/JnqbIPRgGOD9qDoPFwwm4vV8Kmrfyp4zgLksgi/oCuzO20Iew
WqtadAw/wFlkjgWkbTTwEf4sC2MhuU7yykP8cUulzDDrBYk9qkWngNi8aVrDjcAP
8a7IuXBQ35GgfFL5YxmoNzhznHQKJd2A2oquAk0hzuPp3iW0g29EV0LSRA16CTr9
hwuR0/B8Ly6BTrIxWwCF/oO5EIuwY/vH/3nTNxZGjLDLJSMcCZDpKPH2iYAIlNvg
gngTHtIVNdFDTv0cbaziuAQOZEED+MfS5iEFuhcU1VB++Bl/BUJPoE2dT5eFmGPB
Dd1gNH5y1dSwMxnPz9yFrAQqw53bQvc//d5ATUbbQ92Njj2UGI5jDY9ZqoqQ6S7h
8JJJXk9UrR0FghOXD8AGGDyxLZmODqhyCNPm6moHQSaGLZ1mx87rAP9/cAtyE1Z2
zaYg1SP8dZU7Fgud+Dafn3HC95sxID2aA0t4PhK/te3o+t2noHs1drChsw7BJnmp
Y/bxqFw5fUc0hkiJwL+djh+AXBeaIdOt9AXJ+VV7rR4MGIt2UuXmcHL7Xc5t176D
f4w1cSNgfd54nS5ZAPO8VPfgHWFhCg7v2wIGhYd+UoZrIwjiHd6XHPNL2+TTGBEQ
AYNq6lbu8A3lS1suPbjeN9dpWbDxNsHK2hD/Ex+15Y3dBTMLBmpT/fR8N+SOHtDH
Zj3ZAolqxEZerEBFVG9+bfcR+ktArxnC8Q5M6W2Rkq/4ZVBUEKnybR+ZIQZOM6/b
33FMsWcQ+QKeJ/S03o0lPcYT5T/8dVSCP+zeAeYzgJs237rbtSUL3NuW8kp2BQoi
D5P67iljn/BDSW+PfGsD+gtYDUI+E5qHS6f/SvxyUCk7Oio7TeiYrEOnFFaEg3fV
/AY9ZgXBtYmkPMqMkLa0XutcjV6FH1Sdn05eAKsPXFawzSZQnWUFNiqfDt4ZvpLy
5V7jUu9eSkwcMAkNiGXHBvV5Q9W9hVcp5/W75nZLFxc/G6WfN6ssqX5hU0qiyYA+
mklbEe6K6Q0wBO7Kvw4YiYafJKdbZH7R+CsyebxVvaj8S7uYT1HOjjNH71yEyybR
QL0AlfXmZRmUwYtLt4WkTd4209qZnYxIAE5wiAWhdrYT6w6ZpyHUBNenHiS23Vyl
VXYbaZN6RRiEO92KKeO81bXW1k76VQs3XR7izJGdwe7GuhMlb02C2Rr8MNl7NfG6
3INETuO1XcyS2LRG1S37aiBGOsenQo767iUB0cTDcLwT/Yr9vmUVs10ybAYhexMS
ifVMZMjJd3Of4mpD6OobMaYqaD+m79kUxLgm2OzWfORj2VinWpxqhJTMa4aURHgu
yowxRkcn4YjXsDAy6aiBt1whl1CZmALyYzMfbe8er8S9YGyBmHO5E/E39i2f699V
KKUPd5Nn2Jn0Bwi12ggq3Bz0YJfjvP7HnVnb57ek6xIZuDEJkjLX9rHZmSNzmw8k
J8Z6N4BqBoqDcey9hH+2rGXvRFoOrGJk/Bq+v+foNoebKbhxPNz4mCBavN+Yb2Cv
xv2ccEYuTwK2fWsDNntme7NVVxScGSofMHo3Mk7NyKOSQa/SHo6dYk8B6A5rvsEd
xNFEoSTKCoC46jVbUmFCwm+7q0qddz2/OZ9PgmexKl8xnTNip4zl0DHaQ05jBQVj
LvYhlU5LXqGRE7DKj85nx6yJSZ8Zjlm9vugLrbyEbMvWzdWWFimPfjEfpOAHbGNg
J5uvVQiRnIfx9YQZFeEDU+fLjeBRTHqmC13Eq+oX/PtfpCYuS5J7LtG4UU/PX6dI
mKVYM4IFixZ+wfQQq0hk6O+3T3CGUgtiHAUjR0fJzLjbcDdD+2im3tlPTgHhS6VL
vqs71VU3FUmjntSiH2H2O8TUmDDljwTmwJ/r7uFpjd59oTyXvjqbnaqoHRB62yE+
du46U39t8SLprQJJYUyLvTnmpQLxFm3r0KwG0vFZ9zaoeOwieulLKark9QNTV29m
RQR0NUobYYyD0UUGoJ7q1466qiumYYQtfdKszgueDudDmzqqTmS2vKlIIRD8/nBm
6o1rCmcTe8L58nUhYTrsv6Kq5A8fGXLKycYWVk3gOFXFKyXg+KXpqOKIJIMTkWOS
n0gZZApfyVhTlLimo7hbB+ELAqzi3z/MOTRhyTPf7HU2UywugYmjLXLpjhqB+2X1
QF4Fzu/+cWUICpUxouYNdhBEarh8pGbjsAb7qv+q6/jnCxrYWczlF14pe2Bk/rwE
wztYqiwkQtXz2OhovZ1XkeKdxKA8m3vXAoPPdoNays2hRg22HCKMBDtCo/DCyY2w
VNgxrCMG8AYDsfGdHXeJsThluHFa3FH3ar3Ddif7+2o77StahI+DyV9x+5Z7iCl+
lYVlt2EExtP5jlV6VY/geBPlz0EMv3+kopcQtLaqIF+jlRIydWO6pcWKXfTXl5cl
Zxt4mmIEU+gtNd9xL2ygc49OPiJEb/yWaPNDDf2Izxprjim9s8+6LEiOKgq6thCV
VLkRh7R470j0yJ5HIK61hm0YTC7EDQ5HOjXnoYVf1gAqRC5IRBwDr7o/4vQUCVFu
1BrSGTn0TxZ93a/Zi2aLLYaV4pJLXSzNJCJOVraHLLyesCIDSn08U5TnL20Fvf2z
a0b4UHOglCNaFeiukBkZmhsCVXTxo+V8Lk1j6LDpSMY+GGLDDjL/HcBUZIjiyE+g
UAh4oC1feSo1ZZ9UqzjoH2AnC9KMnUyJ+GrN14ZQuleDaPEQmG8DpipuTzI9ynxE
58nqIrhRnMRNh6j5NI8uK7uMKRK+LaRk3vgqhePBtcHFAc7CVR+RY3cR6ykB8QvI
+cQaM8DAJ32JBCwTahE1NzgPz4JHms4McmYwyW/HFEvvyqUX1qrMspspIpsvLqaT
2wvzf8DbZCXIByOUmCCKE6fg3ituOi9nTANNp6yNjvNgK4/uXY0Df0OKnaZUJyzD
Z+S3n64BhTNhWYDVC3jGTjOaYUr33YZLiZSb6BvSm75YVGujE0oWdh0NgGztkTMI
yEIHC/BUN0W+2DrIKa/otxIRW5fMAuPNK1qeLWzTbhI9DoklHB5mu/zTBx+XfGcn
MTC6VxvZuDZsyAnXVBfPgfrBkiKA66nj8m44caVrB9TD6VVkYAEpUG7Ae7C8tjTe
XwKkkixdQEZdQf+CZ4ybmdbMJtFpw5c6ZyN2W/NFRB9aoYpg3ybpNwqf3o+5Izwt
uKUpvIk31QuNMGsgqV9QGizu6N64HcQmDH1U9lO1+F0OLKp9I4KjpGrT2i/VCm0b
mFcQnb/yaPM3ChITG3w1KrbXDFZfesVxDAhXaCc3DxMRyNwwDX8YJ7Q0iRYEB/BT
t7tEMu3HkkC0KTYUlXXTJJYahpccZSAr2TQN3a4wGTKTvftG0rHLRUWTl4N+rfqx
QVZDrfrxnT+atzkGX22vxVtmFB+XVYq/9xYPDvFCDy84CPepECgCTFYrfDdRQMOW
IwwqGI4s7KPqrJTDMd2BaOhUeMfTPit0MO+UlCerk0SeT8/wK0JHr18quIBEqk8F
kRvBKKJP5fvkMHC8+fAgStCErA3N+Mh7ZIdS0EL+3G+hXKoJwMVHVsOs0ldjcJ3u
lHAn3ymJpRnzwYvKYrr9A94rXZBXMq+ghfX+uqXUAuU0/XZpLORQvkhFVde2aa4z
GJtYAF+jQ5WFyF9lwrFOw1nzLAJ4BFqv/wN4CrOi/MQ6vxIW4p3vhbs0krcqPhmD
xLrfeaDrtkyrkbgtiKMjxF1xaLzaxlYcxg+M7x9yBl7yCrlcYyo48hXNtIGUzkR1
cHOZMIfYHOawcNxMz+xztCQN2C3x+m1DsJJqWpDkHXMDxPvYRvb9+Bl0XnKnUJ+h
BQgfee1IqgQd9/TlAZh9+nRQ+hqeg9hgQg9+q1pEMWjwZmVlEryEGl9yjYGlw7zr
+sWkyq/CBmRjDuimOGce2GQfO5MTpJi79K5qHNa7PMlHr8PUAjNiN+nD5henHO7b
SWFuaOS6gfipvvnP6Dp/YZy6suBgC0Z/GTPdSsHsozN5UW3kN05chbM9yUJWR7nI
WqtljpRVxijXqPEE8iildpVS8SBVyZuYeVu9HyuIqPT51/0lSL8OhkFpbVRYHSjG
b+2kmuNWdzTLYkW15E5t8dLhD4oTR5EsGccUq2uVyZq8W2q6/XSXukzNPhbAsrye
2FbFBJQxynNrR+/J5AxBE9P7Udg+icbwozQ+V6ceMYl9IxaO7bCdR2w4w6woND2+
FGAN1DCnNeEk40l+wOTuoYr7mo4EXeb1ED4OUiIfUkSC8SyLriHni+P9VSVHAkZ7
DGB1iOv8ztmDK1zAc0Zrml/zLgssNc2XlEFvYDxd/v6wCNrA4grVOJ3PNoyI+jWX
OY3gJF+Oh2QMUVN5SASNY1qNvYooMaOw9eDkYZGm8WyUJ+Hj/l96XsYMUnyB5j8c
UsF3d7HTjhgmS8iG+NiuuqOQjus9nxKZNxO8O7TXn410+nmw8C7Y/bYXXizHykM6
mYjNdC9h64Ng7gQmZy4ERrKNb3XQtjRkdJAow6VzIpYefwRhAuBohKTEutL0Q2Gb
/CfY1XKNEY4ypfMxZ2d711Z3VEYaUBwVJA0mJd6sYWQR6bYqmlVTIxKHDtsRwRfR
8W8F809/T8X9yw2uAc9QeIl+xa8gGVga6d1WqOG6So+XUR/NebLevBI4rwlSQJ3K
wwuUtlTmsTEDae164dd2Wwv8/2QCJ1KVJzH5SqiBWloJa4S1mmC01ejedRntQSuO
uyyaybGUycAXZmHyCGO5VTH/jKFODP2bs7V3IVn69O0imKEuviCPfqUCit8JfpAF
+8lSi0glvjYYNgU6bzTauF8Bjm2gYg5hq7clcGxG1ZuerKeygS6nJvwANRraCuo+
yWQruQzbGfRkRo8MxBKmjz2JSfXGj+z4beRPH3kryq+aSTHHtto23cVaLUHenWai
2XK8xq8DdM+mDX5dYIy4LWu6xAjnYA7kW41icXFrtzSh97SFX2VM568OWMPAjK/S
Jgnu6lafGRgKJKF6t/cx9RMhZLRog//uz17vdc2r9yiCKTp4xRWKM+FxOXZbNNjY
PZyX1kSkpOunDP/5Hgqq58x82JVGgZRtu9Wsw6GJdtOwKiRiDLS4cEu/+jgJXDpP
abQjlYeWN9nhRsdbaj5hVuyhHfQ/yhBwJaf6lATExyAgGOsxYxHlIhYa1Md0GzRX
/nusayUEvLi1XSA1/foOZ7Hbx/2qit9ur8vDbolxodbf9UeL5R01DuwrHWgA03OR
8eVtAM0PEAx94nFMKc/yD+6URALEYLntuq52RShGBtqLEodhoJ+raVGCi3YgKAJ0
yvT+CtrSLfDkil6b0C8+S/Tpda3/dtyRn/nEkxuRJelP1r4QSX5nXpjc9oIx46O4
wO1W6UdULysZwXXu0dOhqUpX/7G5DlupaaNDBvHRU5gXEHkj8ilTS7mn1DZXAL2k
7L9EV5YKipD23b6CXPrlgJElFe8gOeXbm9ErRgZqLgl/Sx2jIRVAoYmS/nEe82Vs
Mjab6Z9cSkG/8O8HL4yNKb+1FYm3tRNTyUUj2my2Qbl2ECbsQocYam8wV0vtNfxG
1oUiIQ+U2HT/1xt3Xwr1K4AglBxHVb3CRoqt9IYsfvGbGjffYd6v16Nm2D9k2Mfk
SuqJimmvQlsVMIXnomOO3htLleV/IMFFGNS+/XzG/1Z0hokRFlWF20plE/d5kWia
n4fn1th1tqV/d0wJzBsZgQlrld5lh5eHo2aH8t/7PAPmZkN9kourEkVrQM2W7/cV
ZW/whI8ui+47EHo3qS4G1abc2nSE0zw7SVFa+4ZNx+Y88d+9YA2OgRB98ODFFDKB
eAEkWmBljZfHUGjIhuMuWDAapdmlL0uzEWHOnR3oyhjgN3xPEtf3zFdJVfhsoek8
RJW69bzK3p8lnm78iRemvX6OXBGH+KjNBTO0Kt1AnZrR6M9p5OYyjGrSx0e0gxrQ
5Bf4lUkjvi8einMx+OiafrEgRxXC3g8gu0Tw4MmlsQVh5TPEe7Y8Tay5HTzXLWyK
x22PCSqW90jAGyMe69waHdiLIHVd92eDk1k2QB6HNuE7uc0yb1A9nzzSAkCF418m
NLJ2NBsnIoB2S2EpPmWQOvonZ2Ci2jVKXE/sHJhltcbMD5o/xoIt4Ga8wLRKEh/j
HQMqHGnO2QrTbaT9cXwDl9gcaIlLWMfa3BYWsfP5MSUg9Z8iYcc4bhluWfl6G9DF
VYAKKs8T//JeiPs0spMyISUiK9YfKotac0qU0ajmX3Rcdl4IDp05o+HPxcDXYU0S
boVyzCggUahTzleoQBi1PuB8MiNy5YYkB2P2N0E5iBVAlORuwxVzLBDpM3kQUAel
SRirdSaIndnXzlbpsh8R8mvBwDbeW/bZFUUtO9kc6nPuQOFceN6n4sdNUzwYWmjg
QyCJ3tY1w9Yc3dRJbVqVLS9I2O3x/4I1pHcTNPZqVsCIW1u4Qj2mx2RFbUvkxoPH
wN+nAHu25B0rhz/Jyp1mKmArErSGMGeqwLlXQWmxvl2MXvSRAjO/YBYggqo3p41U
s0xrAjuA/AibHlwHtI09oL7wEiLRWzWgbx63BHWXsqd5KWxoNGAIaQr5aGw0D239
9ca2I5lprNmwDBWgPJ9oXdljjvpvjbmJiazxHLoC/yjytAV2qmkZ/mOOOuWVQOMX
MpR5E8nx4/OCwya9sJtm7n1cOP7yrtPpkznVegU5osaPosruzidzW52e724FMttD
aAYot3RX0VSWdtKCGSdSZWwj/m2GXMueZiAqQrS3FdxovSn/bLH9t3pJ8qwz3gXB
pdydK3PkLzuAo8aas/M00f1MaEzZS8aPC/N1mWEjjWK1EaZ6skH9LQISuYqObeZj
ogu5NT/4rkRKOiDKxYQChS/kwgsCaSGQDq+xNwuSb7RdE1kTxcqPx9jQOqAwWPrU
O9tqp7RWs8bFK2KF+q3Qvu18oxFKOYaipPDHinsxlmPSvzlGXSAN4ag8ZHGju23l
WVgA0nSqC6GGm7mpZ/OQABVt5NLLyW7vGWOmD7woLwBTjCnmMj2C/QldSgf8hpJs
qTlJH7ATIBRj7sZ4kBEZL0Xeor4vuk4XdVYKzrzHjTl1Nb/5ANpiJYLe8x9M6UUl
mRrRJZV3C2AGj04GutZtBVpWtE4pUVL+ReXu5CnMVOUnU7yVP4j40R7NQsj8BgR0
n74GoFJ76L2vRCqUFP85KvOIGwehA3ep08vdqOuAJ68KBlo6G7l2gci9WN9acAA8
mg8nqq4OkAddv5V4OmWPe7mL8xt8S6Bdaongq4wffkgm7RnZQQJGw/oxEtO6jMFM
JgIpxMDRvaaU/6XOAphYvbNa0+qQNJPXt9vnkl5IO/c9HLYNM0c6r1Kmp81oeU86
/iq0hN5dBcWTl/sqnqi59b/pQ3VsyJXQsnoC77DBSDkdEDaKdk4sMKhI1MmYpEfb
77y3YCLc9734ksnnwh135PwI4moiZxYdR3fN+uZIWbMJvUEj7iW0zTjQZNu835+8
wO4jsKWqF6o/jD2xyc1/oYkrAThMjBpXGOmrkHTW+lyR/ciGbb5jcO4JfTaoAquw
aT+IqbjMwRdMJ+GkQT7v6iHHcaAjULcWRYiDicwSElhJoCHjeNWcwUk6vwUCa1Ou
eVvrBfGyE1IlWLd80cM+LEPFsOcbs/vIn3MMnibc9939rcjByYVYCk4AIKL5HupB
9Ikqb9a0hiKfDcjkucZ2BzDVBHoDM+tix8hyWBb/K0rkyUTT7YINMpuN+ypXmETp
LcFZCwb2WMLTD3vmzgi0x9MhO60jXDxueCu9H6CdM1m4XLIVOrfL50dn1DgbS9xG
ZP5zZYcpruoeI/h8Eoy4eANL5ddbpJj+oSbVAXfz8qpJ7aHvJdvVQv9e1bbs9SXH
rBip4bJYn+YaCXmAaMcpdvXonFyUZcEBoQunXXFwk2Ddcj/zYcH5EJkO8DWXwDE0
5IGxymfiKuRIbAsF1P1BC5DnfRErp5WDJSbwex4+VysjM9Vg5Yw/IPhfOyDQqHr+
ZkW3WzHp2KMBuxZDHPjgS+wiqiXC89G51xRwglOWqNAekN9TClq/If7xQ0U0eMj7
GuLgks8BU9m91kLjgDqtmD+XAtaKbLrbjhxnagwRRglasnVXg811QsiFWCIvx4o0
0EYDSIKfi6y4cQHJmQ6yKssSNM5epWkEfrpu5BL11S0GPZ0ibGLKs/WYTljS1x3a
euQEchGDaE87ABqYWq9c1rbJ24YqLII2kUGY/dQyV/r8lt2+I+/CWr7rVk8LImjY
V2rZdGRdsUr4vNEfikHF2AlfYZ/p+0hFSxRowF4MlCD1uf/aTqQ2MMA7SaQ/lYpZ
j5c2yRIcmJwQ9gv2wKCo2phcV9PUlAr7OGmkQlK7Cw7cJV5pbKHYJYKFP8JuPnXY
GhuMRzQKaBWp3g8IlLHooT0/1XeJpVaniTeuGztqPJ7zHsrxvlGlUGlK+r0JHnOg
KlSVH7CuVw3jlhgl0HtZV8ggGIUEpqWDVj4rWXNjsuxrXz0x9aglfJEGQab+grb7
4292WjjNd6gx5rxxwyjVlKAP4rGZLXpnQ1n41ws5nRqQv3KPfh2NLG2j58WTBBZY
OBpWhpRLpvErd8R6qNJxNazKUXmDatMtRR+ruWHL/HoIQwLGLgpIHsBCz6LI6c7t
cNB7DipOgeD9vhUKx3mXQs9UlKfCa6lGSDkIGjRM5cQ3r7fD9nR9IsMvELwh68eP
h2JY4nLL8RjNIgBeQrRRtsScuB1IqltR5pgLm7OrjxjkWNYSl5WdqowQT96b2qMO
wIZSuUeYwuUU4a+83GboSJZdafd6Tybptnq/788SVkrmUEgdwSknJ3GLJMy8BA9c
hiZ1YzLmZZdWLMJ8hA6PJlglaVYi+MLU8D4Q6yPAxu/hvjoD+rtmse3hPs+bSHKb
8vFfElJO1VoqqoybAokiKYObD81yJu9NT+WaaV3c/QaAOnNdn2JgRjgDlQ5WYBPC
2LxFGS4tZ9eKU48PIVnOaWsPm+fEOduqo6o/7R+vmg3d9rqFmD4sstkVzE1vIOdO
fGKl4Zq8L8Uj6nKWRpWEundOvlyne77km2gxukspDKIYhcW+VoPlq3/KFGLFRv4B
R/dXJdjiwFmiFiwQXJzdu9i0iHdQwgEKv6zgmdDZ7ysr6ZgMj/zkq9jBWCQBp/wF
89+kDtNuH0pxDq2XusLZ//4Oax6uXoPo6YlHVN0ruIgO0K8NF5CW+xOziuCfK7VG
loC3tc2Buz11VcEPpgZ2MhhoN1nQHgce6blYr7fLgBU+UFxItn330CQCdSmvzMq7
uIh+uhPoQdWMCD9wIIvBh3hBrXLyegp46Gt0rt/CglUKdfI1xnETPGABWFdQyDpN
CflXFSZPVqX0E19nQij8yBQA9lfSMauBckhwzTAyoAPrpkWw45W+CMmU5ATiYR7q
xg+VWbUvwJwwYRq1pggU/e9nyacN2BpEKncHnOgPhfzxKa5TlSHa4L1coU5Ah7gw
fvp1RFwyD9Wf99GgS26TclQarkqM1jVCvtl+dxOYCJU7IKQ1R6++l8OhypH8C9MP
yPBrb2bygw81QMOaNMhBRhY1YjqH1I2TQ/F0Gnzutc4C5K/E6S/r155imomYdtay
AnzPUOxUC1uK0de2ttUrlUwkonhPhGGaf4vEhFCqowlXJ8j0yp3Fk/PCoEHKyJd9
ahf48yiNkpzjflh2Dm4ZMLmXHZI+ZSdd8EA1aYUM1UmJHTFIFvttZoiKrwuru9vx
PNkTtvb1nqZKcm1iPz+xj1fj9lKHpxTUimsQGJwJIvu7a0uC6g9py8UE/Vq0ay5+
W8xFmdCUUwKdNLpLMsHJZOSkHRRMP+NBTPqQWt8Z+4HmqxaFVPk7AtogWPA55264
xSUA5VDvcTWZDPpNAYNOqbBfi/vYVUp3NCiMdx/ObOmSs+QC8PN3IKdJOFO5yNLV
MrHOfF7kRnaTzO0OMs6MHWbLmmO4FW2EtYh/Y3IyPBJQm7WDuNzv1eL6fU96OgsI
395d8spIahyMpO2j+C+FKxQZODFLD3dqNjJoDmFyWQVUKilPHKta/FuGO+pPRv8c
j34PeiC5h77QOapenfUUrT6VaxltEiD80zxQ1cKzxTY6ZUhcsTDbOQeAv3CtOyZU
PkihdonciOW3gssibNtB/NgBfhFp2YiE410gDbaOU541eAQQGWhtgykNe7dMAi6Z
kn1ws6PMahshPp98TpY95dNvcsQHPPpAbC9EKo0V/z8BZDyh2Q7pLJn1NFtYZmul
XP1qOJ8vN2hIIjptRe4r71xjv/MeaZ3eUHkgV1d1PU3zeuw9DsBr70lnRvHiOPLM
yv8Z9T1dHXMjG2ecEZSR3LBZbbzNbOa1vWeYOq6zCkGcikZttw4cFLSL8m3CZIhV
ZF3loZKoJnpHeX2Je/gf5iZge5iWHJBGTwA3dQn9HwrZvMfGkGhi81/7dTGKfH/K
VQXBzaC8aqNU4emkP2u7pgMbVrwvoYcLM+qj9To3ueycGkheT0nekCh/i5kK5EUU
NiwFoBNX2/fhIzBx7eZjhpQaOMtDKHbDMTSt7Bd9vJDtc0lSjwXYF0E95vVxJp30
m/UZWXkTLOxODZ+6ziO8KDKTGem9brFKjmFbqQUDgcNgrqWhENnYDGEs+yjRRmBi
WMMSBA2skLCXwyb10cIJbchk9/pTFy7hDlNKR7Ravn0l9s5O75AHxyW0le2n1zIm
s+Ijq74NS888L/SZ0FnlFEgFRFwr6NvFfUhe8sup4xQD4Sn7yganvbFR4lEz0c50
LW5jXGFH6D3w2J8lG81EedhZvWJk4NzfTBsEFyF9Sd/BonEoRmbWsp1N6Lv/eLfP
yMwjHeGABYJUWX5gmHo1C0NDvbbC6GIKtZLZuXOvxgD83hgd/Eu8dM3bFhzEDdsO
Hetxwx6jWAqQ7MfiPslIhjoYepBDlWOaY4jN1RXKZJkSpVL9An89B0o2SPc5j+T6
g0PTOdoJXbouAsATrQm0vdnoUzKoR2wPf6/Vc27Cmjon9isPm7v5UuVeXIQqIvKK
9kbyanZX5XEhHjFIBIGGSviM2iIfUHiuCKGnCQ5yKTy40FsGW8f5+keBvOXQ4zF2
xp8XmS6QkeXN19TedWfxU3N7iBQV3ctavGG/qXHqrPKCB1gXmaX6CdOs842bAueq
u040zjNeIyHFq5PlJxRW36ENh3icPNc89xIByd0k1IPPgyun/KZ/3owY+B+9I8Sv
O3nhq6I1SIJA+6uXskcRmzcVe0aeJ40BPGzDa6XAkjLQAEbTJYGZEq2RRhaDOPD7
+etLaSn40K/FfVA3DGKy1m++97fTvkfW505mWcjzPi0wPtg5kG8E+oou8aACQFjZ
TBzO1KVY7QcPubpsO+XhQP7oEMssUp9Du2I/4NVJdAe7pXqNuew1Mc5e6Iyg+DI9
P5IZ7pKGSVR7UuRmBzB553Ufhu3u+yAzqOxS1z3XTXpXV1zS56spDPpVlOzit0pf
B9DzvRbmaSZUx41C9hwpzKg75Jm2OcEf6hdHALllzG0dKZvQjm0o1QrtQlR62En2
7QyGTOAlPjjqn7/O0kBq55c/8PFLKu0HjAQG2tK7JExui92A0UpEBYrPpoDjepD8
hMyfq0LlswhC9c8JrKpZXHsHat+ve2dzNguohDVv+8etH06XmfQJpwNRJNd97n0O
KuIDaTho4bA4WRNdN3I22EbpLhnkYGd0H5hLI/TZ6Ioa0ODsu2VhJSepOTMNQ+4A
E5fZIYGFgLSPMeVy7hGKvd84LEl+aqu48sxnM06HXZi5jliosrd43HFtFupCq15x
/kPGmhBtn/wxLHy+llqNe0BFormzXCu3bPdliMrIscHrBODcy3H/hWJSc1kOVCJV
BvmuJfxY/2JW/7R5TbooKcB+e9VlNxSpxYI+lZGbwrCK9/GpKIGW8fwk3PlOwesD
im0APnUHF50r0/WMiEx3W1tGi/FOR2fqqAQ2hI0a03cr93VF8saLa5ytezQCtx8u
UlLInv8qawSgvxyhFzkvA93DBX8ESeNuAXlLo6cTE5VGCHUshLKJOW0PTKGgFvFJ
1Ll8U6iE9xuE3QTBgUVaB9tEral8C++65WKzmSUcvqSFiYGGflqhIDbGxEi0FifA
2ISOTXmVkgccn/Q73YSibMbNhLF3fLUVwzd7YgRr/AYerse0Envw1sDMHn18ptDH
1gPCNGC4ysvBiQwUCVvoH8TO6bbBVQvsiiZnIF8dvmghe+6Nt6PX/6eyC7B2MbAW
Hyd5peU0mfiohVSeNsbY80tbPGbZFwOHkS86yYqMZ54j3VgmvY20MXPVHreGEDCP
D7x69Hnky4Af4itcHV+d26XKzjmvTQ+gGSohfRxEBhXa9vN1OEtqe43XBjoqXkYn
x/p/76UrfjrFP6Kya3x8hm/2mgX1NiiJv02WLa05EW8IfPVaNQ31bZ6urAKnmaSj
0z8LqyZpuEt31/pg634oFVKkF68sF5YizDopor2+5sNYp/xtqE3vyAJeatF7NWfQ
Bp+qbGV1kxJ0pCToHWG6ZV5OkpScMpjwR2CR599viMoQBIYhBOUtU6t/St744VFK
xeSFOuUUr5URLdE7GYc9qtL8O2xlAwaMoM1ckYgZr3VwkHCV1hGPkLBQmGn9Q0mC
iusklnVVjAktoZejrSLhkAgt1kvpbYd6nSujlda01+EvKXtpuvEWNqCCNQrut9WU
lzQ6ZYKpY+r5/EacLB9Gtv20gMgYL9RLIKMDwNYtvu7OWIoTpV+urYACDZaHQywE
icOJueCW5kSIAIQ1/LloPIhSTzMNwFRK81pXEiLO7Sy4XfjoqIS0GM1gvpj7z4dj
omZN7JFZWxQo0CJFxCRy/XWZ8KpZzj7zH3biUbzWCxoZ/zVLqeylS3X90B2ViZ7O
SUNQN75OUkzysuT2woUI/PpIgj+jTceYa5Gw3YESsDJ+Dh9ZzteqspD2drut68sm
qoMTu1uzK+qWfe9qWABTJS1xCSEhekeS5cvSvMbmo4egQ/vTplmm39ZDpHnNCT7K
CmSae5tY1/L5tnbgVXla3jdR4UBpzZAFUuiyUTR1YnG3YlUDV7iNzp+ZPntYJLQX
W9HPEb9+D5KFXW8dP9p16+aKzHs4EmFD9FQpWA5Gh8DfiAA6aENLIcCuUtDTCp/i
N9Geu/uBh9frC4E0zoG8O3GUfT9bHt15kABfM41u65uyMjrtgsDRcvvSJcet047L
mhotieJMMNn1XMeWbXD2/Mo9bqlGKZyXfnRJFpStuBbBRi6ZJoYooakL6Q5Hzvi5
cLCpCJNIMttQ3CeUXAnJ730JZjvGUIuA5rNTfvTVN71zQ0v4Am0STxdJFqW7QqMK
KBTpsElcRVV5g4YdnUCrlAcNSB7jG5RstX0ubojDFTm7pzFNoZcXdHGcpEqAERYw
xTPUtnoxev9VmARN4XXVYt/0nL/I8itK4TYMhneLN1OzhmBRAYrp+WO0Lj5Rva40
VmaLeW25S7Y0PupPWiBUqsPT7tGkhSr7b4JKCa5Xr3NslqKuoyqCaiXfVpul2mhH
fxjcdUM1xIrEfzvP1WwFX0jcexkQ/IXd9CtQOBDqvyg1CrJl96/bwMv1t2D1/hrw
6QgsgTp1TYKn07cpsa8vyylQDvqsOrPnzj1Z3SN65lTgZMwmHqCUlNTvDyVkJUf2
XLzRpdQjAb5hbZTH82TtxezspHFYz4Iis5CpzorNkhmOY6KCXcMX0gKPuMRCK7og
uDZVJt1LwYSX+fEcgrqYtDYjMwOpAL9z2pPBvM5Fqthkry9Vf+x+PgcPT58lWGgk
9xwR/3EjdIkaQODZGDRiSY0dAMjbtFJahlXAFcUU4j4ORpAmnU27g3cv0cTPf51c
3V1xJU61q9GDsstS9PHw7aWXP5g9J9JJOOiPQk2BuoaISWkrHCZcPh4psc4FPdPd
1eik5C6l4xL/9RPKGF/Ox1y1UjeRZ2+30JseOx3qkU7S7V2WA3X3rA4CCEpPeiV5
xEgZDIEX8yvFQa9r4f4L1evlr/myDchktsmm/BARxWhY6Wm07YmI4j1hXl4aDW/Q
kgHzyn56FGvub01wSsusKR0OteSzn+9NeDx2ao+sVKp/fuv7ClvxqjaltLMkaKuf
73i18jjE1oxYN9Th8o3DVlAxkGXdQeORrUeGbgyI7BYa3teaXC1xILFdCti09kDb
tlJYMIZ2nfmpll48HWeBsdcjl3LZz2e8VDCmtQ8sYJQAHpgXRAGW3aTIBbh3krKy
0JsVTf0VY3NATLgPbhSoguQBpKiuftMZ5cJWhIVAFbh9oKvwIXSnXq+AublEscHm
h70pU1FMuYhSG0O8jzTTUwOx+DUQWinDnr3Ul7bwWtfarcL+gNleVZPJo1vjuZxd
Cn/7IYEk4W4QyY9gHvydU7BOviLzQBVt51OWv+T2MXfYvECtSIVXV6sRXcK7k+94
35NiWY9ViKIb57Xof3kr1hifWd061AbaXHC0JpT1zeExIFakLYGPaR53jUwZOYr6
8jCuMLuKdhAk03+ioxe1x54azmlZG+xBbGd0/M/vu+m4hNm5AiIEGP5rAy+R2J9A
cIa5UBBj84PNG9YtigltZ+EoYRftt/m/xukzBreOFl19vsMTf9+55AyP409g01fI
PMFxXESLhIqpsqjdN18WwYqiLr3nMN/g+Dtcy8ARmg2olMZ4O0kL89GsaU7CStUO
3AmW1GD0Dnq+yMedrJWIVcFaqG42EQclaFUP3+ITkgoPUuMC2UaFhgvXcytv38+y
glZOJq2imuynpzDO65NUAtOur+jUILRU7NyRuih1bJUJE+KsUqvCe68mJF00S67I
ELT/nWFNK4qZOn8htctqDCbJzHIBzJYKx7oDnO4TZ8lbDlP+NxuxvyteeXhKjQS+
KK32JDS4IzGUXQIbn8FE1QkLZrHrkA2SX1W5aeYL2xtIyFw4SKAGP8/HDARETpzI
C/BthsbwRSxcpsgZP2+NurW9BitAkwHWrL7Zx/9gZBEp/4ZlgrmEqD97OZ6sdHQH
rpUOgi0Y5OTvJ0kGD/LIj71gPkrofPsvgIbOsuhyhLupUjjskSCqTAze7cAi3E3j
EoYCRq0DwSCbwl3CSyMOMrs2AlbXLbZZKDck6XntFe7rhjWo1U/4c+Jv2AaABODk
TawRn6M6HZuvw0izoqMR9INOFm3kTToGO753ucKNe44u6/Hcv3yctg+xnQ2cspib
bndfVyOLFflPbxbwSrcXNlFL7Jsxo0VLXzQrI1NiDiZDv/O10BM38IcEzIlsMsqO
xIQJQy+Vk+/Ztj55RqBz+N8CI78HpTfOamvyWSLV3RNCj4n1WOEMrm0VAAn2ZNJt
lTSeC1sbjpxMi2FmFNqDDUFVxwivycGegPfspRm9DNDt/d7yeQgIXg3v4l96maGl
cG6GiegBttr+bQBN+5MBjwg+U461MdXhl1WkODxadMEFlgw4uWwxMIOuk05p2Evm
zvdNzj7jdead23Ac7f+SkoJ2JvpAc5Fr1saYe4+wDY+bYyvA6FmY1EgUvwTxoZ0I
/lvh6PJO3C/r4exDATuuunN+ZCuLt0Nw91HFX6jByhGwPn4RQb/U91d/k8VO29U6
8jhYfJGAsvzz0onEffY3dimWDTdgxNNvH+4UsjBGg5IxmEoPy1RyIpejGSjZ309j
RGeLAR/qm2KPMHU8dXLMJkMHEYUU2B4ZEcPOXQi7xdWR3oZ+VZ2v1ATbvd4pdXBO
qF2tAmQcXO3IwJ+vzwBMmOlKjOnir4zFVzalCmtai4K2ac2Yv2ARHyQ2by8vde7W
aD+5+Wf2Hf72uacufPimmoVK/kPUqi1vvMVScSnAOg+CGcck5brLLTz1RbaoOFN4
ZIXLrOAew66lAPbfvt+VAahywYxSUcvbH0NQda1bv73wDa3fySLSa5ye8Ufs9Aea
p6N+K6NRMEQXg2TFGZOEp57bB/NIUzYoq/VLEKGSLof7KG8+UBvl0znFQLM9z4Tj
0aWDn8jv4YwIiTrUOxiaLYPbPt8EMMp2oqj9tkcQYDcOeB9okozjNFw7gCkMZGF7
BXh2gJdHMK8A2twHd3kapk/NtH+O7KAuBItSa7j6LS2dNS5msBvLbI/rFG+qLhh1
KLwd1RNkRCjwE67xvrJSMWzX7tKm8TPXDrEA1wOIMgWnMqtPx+mg3lMANu3roe6i
Ivgpg3YC5etqo+XuXhbx5wX9zkqtg9ekgROadSX4rir7T7MWkI0RJkMeeLF5UpXE
M84hY9O05Q+zlPfcDuTj6zim7wwCUrS7euJW50pEDFUjzaO/KH7ZRavWFJsbLYSh
5NicrSi6/qRIs5/iU22nwbUyGLu9lac21bW58VfuqTDK4to6mAMc5a4cKcrXAEyD
Jl86zNH1jT+zBYPtIhJLLPVGi2oJUHYpr5Pka3MVQ8G4GQ2sPTIvZ3L2yiKZRaCJ
4mH7IOBTyWH/l+54YxNXKMkBdRQeREuoNUzfVdq6K/T3+BMOrYqAYROD95G972O8
YuZ06L01XQ4+2JPipYzO4uNvRi3z6ucMmp0UL35kFVTyDEn5/HeTE24uRjMtl0V7
4/ygnYWueM5iCeDuZ6yoZD5bfPd2YshJVWouNmNifFReG5dm+7JQK17ubeZZ6pwt
bP8fPljeS9Ef4OJwGJtSp5iYnw6LVBFciRXThmPyDH1DduMhXO+bj5RZMx+pbPoK
bE78yTgWZp8QUq3gvfMyK3DcJZVinL6aK/mhCYc6/V0UPjTRleKY4KSU/WF7i/0i
6rG1fQExtLP4kYgVM4VEDYOp9+kVd7LouTe8wdvWWctg8ieyEtLhLzPF65pgqJpT
BKgS+DPM8ok0lo9Cf+nRvgCWrOhcXRos+cVXIqijEuSDQtsylGI0NEUKui5czlVx
gmMHe3jxl0M1sedw5Tkk8YMtJLrCetSUBWkoyybJkZzcTW6HcMOg8pdrNWnoy3e8
JaLrSREt9/FZyk6d8kB/iJhxfmEIG1+2ko3FCRrHya0lMoRXywMGRG75xbZHLEGk
5KgB40P9R4dbPQyq8LndFgh2BSNH5z8GJhcJIm+tE3XaEBjf+nNuTXyX4b/PjgaE
eQWxn0bkjcvgZTrc3HklEH9lKTEGzH5W6a3KIS3CdwnKgyRuwjew6kk2Z3J1hili
f+Py/vQZuHNvt0xn2NZNMXqRP2akdk8QZOWaG48DsN3yB/wbdPN20vhtQBL0F2zR
Qg6x8q9gD2TTr7lYC1/DuVodwrM1FSl6cJ9HR2rhpHhBWquLJkY2M5BeGPiJWTyV
sX3G47P005VpkIPOo7nlyMOpnDMCBpN1FYU31uyZ7pWFR2VgtUW7LRCZq+AZdFN3
QvNc/MeC0fAqtlaSsQH3p6ILzecLIvm1hvbxambqwfSYHuWkrJrU1ifTGciJG0s0
51f8K9aui1xeOegO4cvpvG86EW6O5uFcBgagoFnas8GsBNtT7CAuObpsDA5FUVHq
ffYiSiCvy5hFcxNf9ck3BF4PCGZYSz/nh0d7ZROUOdjWq++WfKJSA19W56ZZSowo
E95gF/H8zUgtJZ+94Z7YhL+uhPnmtC5NboHHqYku5Z/VdQ1vLmoO/e4dWTGDiMts
N8vl4qyUFJD0l4IucCjj07W0T3mq20eKFMQ9+gM3gawaAOZw/MHQcvjhbn/j1obP
moQwb9W+2nvrmmYnZG171uidYKShOWLWkni35cZnBiE/ZKnf+riQGkmNZhXOp8n2
PxjPn7cN4CN7/R6UPy5HtgPRkw3nXi2u8LNkNfVyRM1iDrMi+YY/N7U3bhp+80Lo
qgjNQWcIzaFXukyjZosWmdB16CC5i1aZFxiWQRpDrf8MXNVbG6cpEQ2UbqxoAvaU
nxlBsHuWsAuPRojrTSOd2baWo7AfyFhaCWoPuOsUmpCS/rfQOotv4IS4uxHoui19
rTDkj0nsjOQpQMWdPpMa5P54MTknPgAmLOUioO9ZVO2X2VEi4rq/wMnL0uQOQup/
Mnf0GfU5wqkHcP/Uc+HSPUAMRE2UYr+IeSSam7uJhcEPdnLSWfGYc5BsOY7gZ6bm
FSsvuAUY/v4xz1NrPRhZTeJSNp0CV1Pq+SVhRAj2wSqOhQ/mGP14xgmlYUFnx6t0
v1p6vUjjx6FLW15E06NicemGB0lsUT9ft0ro7p4ryFjeNnTL2KXBlL6TMl1IQv9Y
fYSGNNNUIZPkIg46V3hCbUDjRfQ/DqP9vhbR0tP0rguE1r9znpWsAUGvRk6IzKoi
A9aKEVE/OpHx+YUwdrUxPQ3sflHaLOS8CAUiP1+w87uSL2YJgPs7V+URayN4eVcS
cCa8T4AlUMozOpbg8Z33dluPe82tO1O5Wl6Z+3kX9tRkGfMpj/iABLL80PDWeMxJ
KrUbTOZAa0+ANBhva4tHyZz3fg48nLoDhOKlaye7aXOnmOHrGvhKY2QyWJRCA7bn
JzUZfgk+Rflxyn+AQGXrZPV3/jcbXGKwS13P5fS1/D6E81t3nDS29hYu6LJahXW9
6OO8EmfUAhzzJJJPyAR4hmdVZc/3YgjDOdLgP+4QdGXNwf5vIdyBrBr3eZmdD+dW
G2X+cqF4XAAHrkbipKilinw2fC34uVZyxiUoxVT2E7mulL2nDgh7tkoOXp7lNm5T
LdDB7/PlCXfIoziBaM3//+kxB4TG+rVXnSdsccnRUWNwl83B61dcCPkIzbPtNNZH
Hr89QUnNEtJWVf7mdz+2o+khAUBXBU6BS+gD9EHToQzud1f1utGn7XUcJRAospHH
hNbJ0RYPx7Rf8mhWfKO+Nmuti9w/DhzwhK36Bvd8ZPUkRhkX/hk5KMgc8SaFCwHP
Bd3cgI6I7J8woRjv80mSFf0IvteVOhiQ3gHKCltBqWeuJ2MRmLDYl3mvwWvDnJgl
8rTrgEvmfVJDqJ5z1smUWh4nzmbFj19rQgIaHqpLGUWgG1K9oDDobxIR7a5uDwqg
Q+8G6Cgf3mjMGC+B4kMEIL0xd9k8lyfs29mGu1oZvNvK4LsFiklWwIddRizSfhMD
NAgyRUBLmyZZFLdlGXqFgeUiIVDjdILaEs9FiMVHzt3gg2LTP+BX4qG0XMAL/mjc
Xj7ak4f4zmNRiwfbXIOdNLPbJKQZhn9XmZsKBoOaQNHzrvqzoWEzrOVTVUjdJXif
2MC/yiGtYQU362v1r1a9f3/apYRwhYwLnN1ZqEALC6RTGsNo4UCFP0ZoqGHTyqT9
C/0RSCzJQ3uW2T2aSJyDUsIXqcXQNIfoJ6zV3zTdjvXtAzl/aAt5Y4MEClujqCs8
6O30b3H7ONBZw9jUeQOy1USlLQsDP6GL8T3mhLY3KnCUmjPRaRZ03Ydlgtsh2awK
02cagnOEhuNeH2Uxm9swjhgu2hCoBxa9TJJLb4fw4WIXSGhj369fi5tGXcj3tZY1
5jSsmoOHQ4gI/HAOTaJGVMPY6qVVsaGTOlO0IQ2kAiZDlgyGn6mEqE8b/T/kAFVO
eK/klM3KWCXwB2dHl8QulsaafTWNMn7/LGCSStLvax3PJljij+BzIPpK7QkaesiI
JOC0C5TJmcMjsJZTVC3J8kfonpSMQ/BYIO5e10d7Cvv2dPUHXqrL0TvlnoLzS2Hc
rShyP9Z0g3II6caiiRmp1/YG3aU3JxWcgyyiDvIjriuxm3lt3/2Hd9FO94gPFtsR
HHj1fCT6sSmsQr8uhK4KKF8c6s0ZJ1On7YtD4E0IoNSR03vyKPYnMhcMh5l7eGhB
2wmBaLda/uO/2b+1egQrRozL0lRivb4SZjMcFfLi0Ug7yxw+THDWxDWZspzQsChQ
3tdaE4vsrBu41RHOHkpEgXWMCjjO+IyeclI5KShufu49dNRglkhigQl4VTDyDTck
BVgizPU1c1U7okR5yES74p2oYBTmDeoQ6cKsg7Z4lVw/Gqp9oqUl6RdIG/pIhUyU
C/IBXM6Yvt/esLhbNcJda5g8M1QTCUSVeDH0ABcKY8rVyaPD7wChf4TMneAFqjxL
hKXPT+ETrcVWGot2ukJGkeDXyRbL42U0vI21ewSUZIHlvJ4k4VskwtQ5NO76T8tJ
H67z08uozD+mbcg1QLCnZ2ZtxLiNObjCxKBJEPByWnHp61krLG4yyVRdqCIDmg/z
wtJ+8qZJvDRcRQX4+Sg0XYV/xwSLWyDoBHMp54twmRpJp0Ytw137Rwuglu5QCRM+
sOahhMCRfFLhh9NibhkU10uHz9N6Ow6rruWgpG2C3YBvoDEP5cpt9pNnLAwRLvvq
L7zdiwfHjUhZx+GlxZaTKg7mPnb4570G2lTEmFjNZpkN1tRb4GPnclMPC155dkEY
95j6jRMJ3w7SCgJJ0YgMJPL+jYKvXtv9kSjFQAobDeEqkF6to56K1osV+2nKJCag
TkRH5xsEN9AKmxSO4xuDNx7n9c2LGJlkIEGiIsEMMn9WwdIyjHyq8TZvcN4zcq+O
T2OkT26W39djbU0Q11/lLApPN3KoMK7vh6Js7lrgiW6APa8LL8mMFoaIYwT2kdqb
M1vyHrIPAo7VJBHWCjklkh0Hq8Sg7PfVUD1y0BuvIPlr0IpCHY8vh/D8lQhXN/Fe
lv1DbCddH5f6UMtzKC8TkJa0o4vBhINxCAYQIiJJ6IhHNWWCr9pgk4sep4rCvj/r
zjy7naGPZdauW7Sk4h6yOXo2nX35vHJDwt18OKesWfUeDDPkiHVZk64D1/sK1pXx
5+CqMsHz9tlEf8YLTVdidv7ZASGspJQ+weFBTtSFH5SMTge+/77+zPAwRl1P7a7w
Y2DBQsk5zvDmHaAtZir33u4Geze9QzIS6lyb/d9nhWUjhcH2kP/DhMA6CBi/EPl/
gJluF/VY94GpAIkeRS8LJ2R1waoca1z0XGMK7VenPZSs+oYuRfU7553FAoFj4WQu
hxWtVx+3yv/CIv5wIcitYBSJ1d0ytlpqUH8Gr2H9KBDTCKGIEqw7EFOjXx5SbCyJ
MwOWZ9h6q9V8QkdzYW3gYwmmjIqchI0xCMfWwQCRMY64eg+IQcvuzjtrCqxI68YP
Tq2rRcIFcSI1+1CA0HUGQ9ZYKdRkS4utzMA2y5qE5GX9cXyYsqaOkYyx2QzCI9JE
ojWDKpDjffETI/gZumfHxRby6a83I/3gajKuGjFAwW7hzeR7iI2zOzlE6Kd0Nx0E
MxpdV8BYq+jt++JYsRohFWSljRI7GPnjhOSRMEfuLDFbV8ONPkWTmda6duFnxFbA
yG4vSeC20o9TQa2h/h2LHf1zkhy77xtcr009fWHpy0Gq7I3/cD8/B/AYbfIhVSWf
Hm+f7T8QZ3X2kqPtGtf6G035FtUT/yIk+2IFvs4mU6uDvh7fhyx1WkyoVoif+vBd
b0IKlwjXNlPxWBptV3u0cqqzwXbRwvsfTyrb7qBwjGyx412YpuwNdj0BKGHwhtAA
J14HUPKWbJKPCxszD7mGgpx9nNYN28ufopxIEM952msUj4Q/87b72NW9Zz/M2RUi
UV2bVq62z9hs0ajsWq+nyapUQcxW3FtosXgI8s2qss+NFHa+XRg7+hXmqEPAYn0O
oFJ05IY3uzXNi6cSvQVT4C+vg3kBQuTuwrUGdswOnTJUD8y2F1F6MRMsU0hb7Ory
yy9V+xNWI5OYLVYIzcAFIrKBh4Yqx+E4GjrweS41hA+9mTFH3AnlvhBm7cNPEXlz
F2o3dhf99b2z7Z7Pd6+UTsvIENSVoPY11sBtwkaY/4qQM92/7Is8KlA9jqAIASH5
VPcg1YdoxI52fdgc/s4rv0D0wrdZDewFGbZNccW/U1xyyjuWwPL7UcHy2cEddzR9
zNChU9qFiqWiptcKBTSTOK9zAZ3ZVqf4u1FY+r9Ecpk/cefE77BWRMGfXXKKG4ck
RyhHAv3tdVEDhuc8o2agjVjGgAZzWiiulCmFopf62uW8+IoOBecT0dVmERuRv6ng
hfMufivtMwA+E4zFl1czmL88PClXCJL1bSKCZVV+5Cj0rGQ8RQClpnQRG/7VQARC
g/6HJODFeF6kmWrBtssbs91jj5Rdu0mkzZherznLlS47bv73VN2xo8HR4WRmTsWN
q5Yr2eGyIkXKYZi0yLtlFGVzzCM7F9lURBnVABqGRAttvqb0WHmbBk+fgujdLjK+
isAOg3rQ1clZPcflWgO+q8LV+HMwdsyj1xWOhEhDIp6ibCupN7C6UInU6nYGxw4D
fWz6+O4TvF1I/e3yQKaVWeJ8wqzwdm7qwF4pARtDEQO81MBXnuVEZj3uYQMubzAq
7ddJOKYijvyrgUgNeyq6NGU1aq/dSiMW8LSVu4EH8U+BXz+tZqcDIRsZTk27ic76
sNf9QhbyhxkW/vP4f514YQTVe8Kzm+3twVsicO/60kMsFttLAB9dRmzP8Ign7lBy
KD3Xo1Ntwnaq4t2TV+ZUbFVwNixsr5EouspfuuXRXHRSzVPssNK12FpKrXs/chNd
HRJc5aIRigs2twc9LSBb4D6CIbnJm6n/6fQkInR5II8FfmAf6cDS1Kk9ZLrV9k82
Imgxj1bDupz/8yRYVmbU936s8IuM4ETFFMU2Fr7fX0gPIN11wXXdl1bsMpDippsJ
fbG8VZzjdJXhTGMT3SvQSlR+m1ztMk9LtAdD3V29vRmV3YAuyZj9fIENtmihLj8g
j1CYMUc/SZdtEoKwzWbWQDv3RfALPOR9ynDXhLb/4WWx2Zh0ihg2oosA43xUPif+
/uUXJOanCPEV2nSt5d1G/fabO6EEwseM880oVyeZvGoF3cnEwd5YF0VDcxvy4LnU
eyYhrxaz24YZPJieTOd3k3FOxZT8DJ9kIFQSOD4MBIosx6WM9S7uXY+h0fJetKve
I07vXcdQu+nhJEzCcVQmee6Basn+f3w0OecqwV9DQoykLpQEl9ASAUPoiJcTqv3j
wVlI9zHhd2YzENsBFEo80iZDKVMpCn1B+gNflcaW+tvU3yIiZsOHJj3sHNv0fU/y
cK+wDvWY8Fa+LxhGNOItBtB5wGtQJVIi883pA4mQRpyy72w2+EEui0jLGGYlxKFw
1HnBzoNlpoPW5C1/lGmGp8uke4COn9PfWVIil+UgEDk/pUWOOxaIGt6PY2fmhsCu
0QmgE1/zUbsqL/yEPJH1ho+sQ2cG9FoYHH0V/egxb3/OL/iEEQwO3y1XzwMJziXM
5YUF6LFNbKswVPA2Dg6ygC5NK1F1K7vcLnQtPOkhk/slCJ4Pth7epQJ63FMn2v3M
yn9eW0Ry6slrVskQcXay6qrzqgVWTp9kHkq8B4fDX8iD/9PiDpdrdOSRsO8/Bm56
M0KaJ1toRCPPGrVZkX3sjc70cAh1LPoAXgIXN7GCs8oCvKRz+bP7XYFv7kcEP1bn
RxMpV1TAs9/8rfRiOnYTfmUOr3OiLMuuNJbmUnQILtrIIrKwKDZLa1PHwOul5MXt
ConBLdzA4PfQJAPOxWK9foklRc71YAkPslwPDogkBfCz26a87rLY3aKyud5YlijU
Rj+qVi1BfZhFf96+EYXdOyGfJ6Pj1OQdcfOYIcUJCiMavqly1uIrq6MSZZeIIcVk
wZyOyQrXS+XeKRbQouKftUMs/rkqHlFnDXsPemgs2CqVNOQ+oqN1zwoV7P3FglVM
oVQXRTkVRW740es3830xVkaFFhqyULtjr/AnefK8DvwTxJ4avSoGV5tC9sTiXZGU
Zs9grQGCdQzo/bQszo14CgFQD++lUV8xmd6P+Pn49gVYjZVYg2jCG4lVY+eIMwuM
0ltAwKJ+zuo1ucgI5629Qt0qGfCSzVfVx1T1J7Lv09KBWjlLlkhPrQS+BRXUfGW0
QEpgGmBzL+Wc4GtB7iPrTAA02uevJjYON/Upze2BGMdF9hwwWTRGKT+2JZMiw5Vk
StnGLNl5ep0wkzT+UOl4X0FQwjbCwmMA9VrrnMUQpAGpejl31DbKeZON37UyCgpE
j894kkQzyjsCJ+mv0N/0ha2O+DLlvrErXdBe2dI6NZVFV90BA5E9raqitKUBytfL
2bOIHlMnVnnbPSr475htwMbltH0QcXC9vs21ROYTeLwt3qFGO7Uxk9/YqTECqxil
UBs22ph44gaqZ+kymfQ9MqUp0vN6zIHZO61r1CU1+yySSjY07manCSVMBYO7MPS+
SMfyFForgegvdP3ukYpvGlUFwgpwihZuLefn3XrmnOKfBj6wqAlr7jj8NPEWEY+i
U2Mu1YRgXdwC/uUmtyl1r6gZ2CLapPp7DHUZqzGUlsfAjfIVIKHptP83MBg5Bzfa
2N7GU0TO9Hi7AiFcPWS537xgw+tF3DMFfNzDetkBr7BCrhgcuXp1xMIU36rwYtW2
XP1+rjeASBAo3YMohp1y9OCyafuT0gqwm/cUX/qCQ3Xx2NdNywG81WeZQQcUP4DE
zWhsT48DJyEhrIcrDIAx7lNxfYCDfmmOBSh9fPoQhbhuPKQeUcjU6WfgiRSQgdJs
+CTqykqfGpWAGAinmj8N/ZDlVZHM33IRZf9dznGc/O/+Ui+xuveskGBQBq9v6YBj
+fvEb+zv9kU99RDvoFA9tvCJmd7xx3SAxwrZN37psPyPovYt8MJ3nYaHL+oA5j/l
0Y3Bwu6iYXTK0zaNsu4aOUbyYVdnDu0PYbGOlF3QryZre7BaRHvRscCtaICGEcml
HVqlseBsPficE47womF9GOCBezwPkjlbJYxShj9NhKxxb3Waar3VAMZVBmgZ8SxU
8FxdMgQq3yT+iKIvIQJ8+ArzETLp/UK3XLSGA/Q2WKaL4FEFpcCiMNBVpHdmE/ht
hqV65iUjDnuitJbynVbgogmQy1yQFAK70Xrx68J7C8uZQJA5FChPbHtiktYg99LO
LtDl1MqxKJZiDqOQruQCq9pmXUcP/ZSfEhrvvDIojIsOeBwKezEdUKqUjQ065c3q
8uc6C1BfQ+pNxbcVT/flKx5wnUuoqjsehnGFqtWyt0lJfwJH0/apbliCh0dSeXpx
ZG0jhXcPHmSP6aNNS4KDUhHDpnhRZoFDt28ObIeEEMYComCGFhR/VWPo231APPvf
94wsq+z31VfGwBwBnkQH08RzXWMIqStCm0uaeiB6liMn8Dm1yY99X+mrdysHc3vV
MRTbDqSw1uHH+it2VpnUxaQMm3cp81UdA9jiMh0bnZxYuzSEYBIojJ5WO8pIWs67
JrjsN/278BHFSZtqbeVk+rE31hQH6x8zEgd/PKU0cuzv2S3DYEcCQaC3Oi8EsVj1
qDWYI8IcsryNmxF1zq3MsEj5UQRolKRg224yxC1TH9t8d6YKWIcOn6DsIJWilbWh
PmnPEVp1nD2+NORfbdKTceTWP3vnu5mH5y8t8EldB/3jSi9NiyyBM7ZHrSqH54PD
S5NUbps23aqLoRNllI61/txgSyCbdLRofAF49B64PDBPtfY7e88oij0u6MV5UXeX
EYoWtnFCVF6pHhgvFU3MBZrfZANEmKbp+gUS91zxDGnRRfwbLsssE2wLFFQXBIMP
y5oiC4+bxprtqC+O/zaXPMZjM1Jls6nR0kM4vF8/PraDLJMHRjxpbWReeROSjCk8
+OHwG3Icx6CHSvlMW5rNh0S5wv1pubQY3hdGE4Roz8C0SMuk4CCQOAY5sFHy+woD
SPjVX9m4XKIRS5sGiLRHKbNae8z22RI5yzTI1DiaNL2Up/xd67LbDFtcNa0sw0dv
a+33evSbIAqGBtcnJCKF6wxRt9HRoLBbKsehoAY88udK+S+EXrDCTE91yKrgq3uH
zVktpK8DliCY/iewsi8EzbHA9FE9mFaG68DgCNDJbn+tp5V3siAM1BlTOc1ws6TX
wJg3oLjmtHqATjvjg//TiB3xI4wDrk6y6GKyXAUKQOv6R4Mfe5IUIKjpoM1IdN6/
1K+ycZ7KIzuiBZ89A9zIpoTsBtIvWJB0uR5oSfDCxPjik0ZuCJl6EMSHhNSOb/BD
A2K/MR6u0hP3pZsltiBT8/ivVuZuPFQJhq5BxzDVOCnsEjkbMSKC0DLboCUimvEN
DpI+kVACU6khRSMIDDI7ZBaSh2v8FTC+7fBluterFGn9gk8BAUvJHaOWMVDTT8tu
y3muk9s6uEzRqQ6l2ir7WgWlwOItmRPth5q88Llgvraj1PZUuAC3e0ZMh6/rpJm7
yjmpw6LC14y1Y9EAG9mHq+MXn//zHFVYMOcjT6ZoCABjtryS8B8j38i1q7XsLhWH
GEbx38QL+xXrnp0efeFqcDL6V8BW6tdSvcNYP1GsqOYgeGjek1Yjyr0JmeCRcx0b
MXW+t0HTRIxjlAfVpb+up8Nj8C5BE2ul+JoXhLj1FGzjnMsvHbG5eRhhz/ZJKp4O
I1jb6PEb14WuMaBY6/nfD6meWg7D+7v07aze85zDADhL7d3m5Ol9v+w+ZeA1jqf8
tQBlFG51Wxp7AqUKoZ5u2bisuMIJ7fJlGFv5rakreUgVI/cTewZ5pX7LcRYCRnrV
q+gUlstu2c4QMDuuEwkcT4rs3p6JJnhHF4MaB9BPZDU6FTNP52aJOJ/T0U15OfHN
dZGGu3h8AlAOzki801kgVSMUWsTVUDm9/6J0xpt4CCdhmn7rbeYUs9pg+0vrqjy3
oW4ayoSK7BHQw00nt3YRDBUYHtwVANu9Sb63+Oow5QPErkuEoZCcYK8PXzcTgprd
9ZWsKGlN/Tf7dhOBFN4uIPXZtQA2VpwISDslEf/kpeu534gIxNe1CKZRquTd12iL
x0xK6rFjW8lwMEjTePqA16601uR8HwDM4IVoAvy/LLdBKjFO58pYXRBiBhTYsuAQ
zZyeKVnBB0C2DUgcDOhjO4O0aeOTS9SZJ4wB436H40BdSscktWgmaK29YIJeMbLb
5j9Z3tVwgeAvy+wVHL6T3V+D8wbfPI7EJlv2p8kWTfsWePJfqpKz4ymxFAOh5Ws4
QW/hGULw9ruXJY/Xj7lF1YW0lByVi4SmcNnFH7Dr4THYrHTdRCfMaTwGFRS6mwMU
WHq+rOfuPEIK2exhYyOgECU87nvtJR/07E16YGJgSHCSax7V1fjpJqVC5CZVW9hk
vlifmqVxao2HkAv2Y8PwgMbiB9TciR9b5z3n3ITj8bIK9fqmV5SGq7QQpEmE8vSB
rZhTSRIH5jqdMXHKL0oi4crDFfK8Urosn5TKKUNdX3JmwzVeQcTNcbFuLf0Y3c5L
GcyQO6u62awIseNAg72OYml3Xmh7CzyJgvL7FsAt98Av0T03lcRVEf6En7wlPbBg
94U21Dst6n+MKebOMeZdOn99dc39VxUWSsa6hKvPAX7Fx5qRM9hjMef2YgrX2XV0
YlmmtYF7lhxzpp8amba4reqmAkzSWe0txUObGom0T1TrWLgZ1fMlP4es6ox2U10i
8WYDekNdw+kzR90OxbFSiIsu5KH95QQRlSRKcETajK6qFbHsMJoIHdIzKNX1TWK1
IC5E6mu0PcROVDcYVJsYLmLxBT8iSAN/7gbPWlrRyaksQgoXVNfAj/88Mz2DVh4O
qkl5j2D53Jhpqa9jclWxq0/KfaRG+S7a83tveOR0EboZUS8shGji1gRU/tI0lVl2
3pgrEpZ6l6vfbE+Arga13VPz42uXTTlbxc3bu8LDovKuC5yrZCr+7asfPHHg7K9m
wuu6e5wgYNbtu7QIk0bq8dy8dmQVfA30gJsDaC42bvJZzt6oPyYJCoWsxloOvC5S
40kvJZlHGgEQDyLTsASNQRVUlKLO09+5Jjf6KtR/uWjnM/A4SeGgKJPCJ7Q2ahow
uY/gc4mcSXp+eCM7KYcTrmlzpFiVsuYDyMG52Hz7Y8VAs0qec6XgDVpBPpcUoC4g
kQiPNbgVc0AZoI1T1Zyg/5iWPONSWUbJHqvY+mIv72LEWz62iPglfjcezw3O+v1h
7jS/33dbox2eSA3rtDWE5rAavvLwWzm8mZCtMl/1uoiAanDaAn7QfOT2ARCUuWiP
07AWvzE6nkn9tj4S9zjOyxkwSgvf7Y0RqA8m+hMN59v9Ch3zeEPApekA0p99/ze1
ZJL72wiE8Kj71spHyCpMa2N9leC19v6x6+DiYFzAWPrPGyqI+toZXb7bkwlwA8Ei
mkSIfHx8MfqNUYNliZtsULIHmpoTIH+gY17bGzKyyqgcEXmDdbjTHg9Cc/6f7oop
HVtytfUdEtHF3yUekzRF01DPpfrmAK176Slet/udA6rws9rqN36ZSb0f4VXpHNFf
b1xhHO0EIdFKvddZtWHDnI0+3DQ0u4fhC02FdEhb42an+hdAzxMaiX5T2NKcwBtJ
P1JBqyW9ZUXjbSIekcRvbPXa8HNJ0oxHheT0tRZPegDzyRMJpa2GebJ9udt0/0j7
9uLVHXU92Byw3tf6WWhgudbqYEmQyq+mJWvtKZkioZ1Ez2oKEr+hyIhXQBxg2OKe
X3QX5rVkalyfhyIbDQ6qWJNWe0jt3VraSTLRjatzmQVXaedQ/rTky98vUfGAw+G0
nnSmygTWG8NgQXlhVtI41nr8PpF3AuT9PGEhQaYy5aJkzdTd7DjCdSazjmSfDClC
HcPcxDOswZtnb5JwAzhaHwzr9+beLHuRJiGZJGMExVh21bz8/JjFd8/8tkunZFHC
iH2SlCN0KKCSJMmmEgjhkymMa5l99goimvlL5wiwJluHYjnIuhFeO8TqxLZr8ozH
EUxtnPgX+7ffmLFSIEeUMPOvJPEsSppjanWKlGU6lnXuIgDoVaFNjaKq9eYPino2
SJaWT2HV9Z8TwpRkxbgHxq3xRDZEZfvqtLhXxof8xzpwpImmp5uuJdxSPdlAiecU
8R/f8JXt9ts2jpWNA381VI6mPZJ4aACB9Q0Qfsv5fjDPpw2+cysHnSajhnt39lgT
Dn6CNiaTdOT4Djv4F6egpKIOLMmx5zfO8dRMX4EcJXP3DODTpPTfIvyraPGgHEJp
jcS6d2BbQhEyJUf+dtyHkVPkkgP/VVYfuLe+jSlUcJeIuGJjn1+j1wk6npEkAzTp
7jhldW/bJEFW0Qsz/08CQQj7mzJkrb4MtWRQYHV0kZX6kzgiAqmVhRI3TE3Y9prJ
bqtgPl7N45EC5E0CeOt34fmimPAFEgMkJLB430BbOJ/6y9uvNhj49waaszvHaOOC
7kbTwc+HE/JItq8nX44PDTCKH8L/og4HF2X0aYKC0dAr0Yco58NbFgzt6Dbwb+zQ
8gv2DyDVeCsmEjbmmQgh+yvw76aAQiiYWycgiiUo4l9OgAlX8qgFrOo0kzOHJANb
ptw4nAiK/PEJOSqtBT/8xWh0T3WUkFcwA+67kDY6t/l2wukl1G8gn+SyIUQnb/5B
nEzR1zFj0+3d50fCkpiDvSLM6RBpMRmoKLNENdGU0FrwvifSx/XQOjJSvdz4RgeO
3MOtxEPU0u2A42NwG6mFVMGlbUHHo3rxOIT2O1WwNM/s9/vxDgfTNUcBRm0Fz0AD
ZjssFYYF+pSQ2WSy+Ajk6B3tTm4ueZdanHkW5/QpEBJgRu/etnf1rFXf7duW8v5K
lASoF2YfXacWN4d7QqCwAQCuWWfERvMYktYGPXWmnQyw0iUJ25SRf59lCzm4MBpa
bMcLbHHhrAsvqmAtfGsOdseSDKCEDvqnnpU++T745RmikGW+FCY+GzQ/jIW/9QIQ
R+2gpL7bPnbf9vFel/0l4CK5pYUMGK+w/isn+v3NAw/s3qfo4SVZOOez84PGm7xr
s7XmG6D465F533ARp9eNkAG4aoqtK4eKhiTobZq8PBEjPGVMLOK3CC7maIbm6z+P
2SaQnXtal7Jgd3vVQhOx8EComLQUf0MUKLRvMH3M24fUIpPldZX5rmplA7yyUINt
raHl9jAGq+0KgNCOi1CY1s3AHdrWTl6L78Sged0k5awGbQ39GV4lCFkl4lD6hjfn
66bn5u51NMOnkgbw6moZXakc+Z06TMv0TLHpuGIdviyDaq1XJNicZuU/kolhhKH+
lAII1D9e1IBNhJGJt/w96Uq3OSkj5UcUo7nJsQ6Jq8iZtRtqpbnpljy0NTOama32
u5gdO+pPWTD/iMByNronsOO00QcdpKGna4dj/vU6bT3CnQB81u90rLZ91/PRCQEO
VjvoxmgOv+T4ZiJVNdgODP2zhI78UbQl69a4gUQcLEdBJvAr7lNgdMZ3MXkZR6lv
A6eSdJzwrBW/LIDVsBZiAgQhGVefAtYwMZO5JPYHlMBFkEwsdpcJl2asFzxgfdX1
URkksvVSlKWvgkb2x6nxM5ZG5zoXMllsMGPMv/l6x1M6X8zBd1IGAOOR/jmXcdUI
2lZTVLkZtGiGNKS56M1lGkMk1cRGU/6U+/nrRdbPhKvs7NxKhCFtwBI/Y6YZyHF0
jn0HleH3/R+SnJtAwEcnxzUbYwGI1HDnAnQWyiC/9N79PxtYUn89ojMHL13p0wQG
iDKwdarq+FWX3RnDJCOwC2WVNnlswpd4Cq+VMfXE0UO2rPlXWVrD0zH1Ea/9zTUQ
gveKhg7Xu48loxgUAqz22gqwHLB2C4LleFjUl+pMn+HI6RCoQl9UZ4xNlR8bu270
v/uqKAZIeXkmmgSrdVZ1sV0qDF8fNYTiYTY7XEgkUOfO90jRUpd8Ec4w4Dv1w6eP
LR8HaO/k2Ng1571oPF1PHxMmjrfLg23amn/o7/Yr9e5mVNV0HkUrStOgiCW3kBjN
UeN3i0Itxplyd4IGYfmTHqcfOnUeayVgDsEcqfFPMJHqc1yHFonQrKHeQsSGOOe9
OktloMjn7PNljhgyT4Kdh70hdpsVE3CAo0eK8526X8TWf+zgjZ07Q5HDDez5MN0q
BRIs9EroVlhWKw3ZV95pvlX0uNxyNcO6YWDdlEf+1DdkG5wj6UYzzUAxU6fwTao8
RYh3qZA53Fcu4+IohFAQwmc0onGQsvnlMn3j19AZR5cWq6p2s1SuR84HKbIIFSNN
NFfwK1aWZnzAYQgfZEos+AOzSw6uex7xHPwPxTSWGIl/iTXr19OTVBG4s5cbb8ai
mj6c16EKfeABb1Obp8Zl0GYKid2Ky0p7qoGJLrZCuNotp5UsOTfOiW5jiu/+Puy4
o/BiqRPQm1Wb04nTsfQ+HtVL1zWT4dl+ZHOrHQCAHM9II9cVSgSuhJKKGOWd50/w
Njs5XJwZ+nVUU4O/uw+vl1lxmtO7I//OqIr9u+uJhlF1CJTvV4K2f1OHg+SqqtD5
tarRTi7xHrPzsklvZ8ho2sSsMMY7jpuZRBKMECNRAzBzztuJFTlHq9DB/TM06t5e
gl1JI9ycBrH/YJn0yYLXKMlFxV7kqYUa6RJdAWOnGK10KI4vTtjOLRBXEyx5X9tg
Xct/h0Gh1O/LX0QCFykvu67YMrYz7MVsYkyWq4aq6U+FvyrTb74jdXdNuCq7wnbd
e38vGWnAHO0rKkOfFKdDRGOjUmSTJuOZgOuXG6SV0T3Zw3g1c3gce9MU1IYZM9nT
sQCpA7e4M8pVdWbH7klAU1XHWl7MMAC+ispSRdZhw4czHjmLvxlkLMteHzFALlmY
Kfci2/lBF6Uwr/LjC2zJwHvkt49QR9F0KrbzoBDt+f+BkboX+z99Vv+dbQHm/gPF
aJd3ZCeO/yQfFtnr5Nra8OL7MZR3V7znMBys0xxxljewRVojtJY2a5GERSLYzng3
4K0EU8HYab9rnx60lszqc2C3CaHEmPDMqCwiVfBpz1YC0cCCUJUwETWpvX5TftZp
MH5vEhrQlxtWzcXWxmoVTcgR309c4Q3vt7jckkNA0FR4k89QAMZ88mk8svtPVAHC
bAAGpLPYHDpfYjb/qSMcnH5J6aADXyozTBQkwTDx6CNmpCDzfD7dExaHijXazFf1
T98BspCWABrJ7VgDR9a/vBKhpBb4GvzdM5GwhW1m+zQYLW25a11V/ORyo3xHwRVv
cWD3XhudUJk7tOgZAZByqeUB9J3ofdi5jlLY5RdPYAaoF3GkZ3yE97K2zIdUXIJP
0bP9ehDOFN+RVhWwJrL4bW1KS9mS+Wg3FBwmcBau0I/ZhjjA8J6x74HMk+ctT3nz
5sW2Vdgd2MleGyKvvNhUrRVHc+XbPvS++ZnLWjhiIAKLEztcSlnuCCTfG2yyQeZH
50SHBx6RWq3LcL7DixPODDEajsJdk0feC6ThrqD8J1sAQlBb5Ll6GIKvb1CAPOZf
Bz70M5A2NttFZp4KOfdWP9mfF2qEF+7NsHwHnD3EP7EPUYzGwMNVi3Uh2y+iv8VZ
FZWUH78ikpK3N7m8Zsxq1Ao6vaSE7T7TckCXpRSyMNXk2E7kP9zgU/cnfTn+dzSp
18WZWT+OR1teMgiydDDPVVEUr19hDylH82FsNuOtr/8Vq5kMS8IqTsR0unmcAzrI
R2X7lfZyhesNWahh5DnH32pHgXBKSz5Qeqj7LBGEIc7EK4Uc5D4iNhNZDK2pHLT1
ueUddu7jlV+g6ZnVo8b3+n+Caf+svxa0GS0TiHLqfxZ/CSlZ8puwBSwIOHY9+qyT
onpB4uBgjTKzNHZj7134jh3EBL+mbkixh2WD6adI4qSN0I+UdEceHLJCsurjMSSf
BmdT0MlpTVFZA34QkYlX1DDlzOCOS9oUx7tVMMR3h9FfrAPlESSoCaxKZ8KQ4eLd
GmTSb54tzS80Gy2Frr/i5kKqMlvO/8nvDvDAFylvmd8luktqCfcYJ2ER1M2fbO4G
f436JDbNH0S3VzFadk6QWkOfD5DiE9/ec9t3huM8anLHWRhp4TM9u26eJRTdS2t8
hyybBxFZp4F/ZJMK2LhhA2sxUjQtx9k4sansM7yCUHZ9EI/GUpnVhL+WRw7VEnBk
Lx2JcXuUBGN7Vx1tdGQ/u7c1TI6SiFRjploKVfdluIdnCsrVbfpd4oEEIoXQ2KcD
c8aT1S4YD7lFpIp5aK3QiRrRRMc8wesnF07m7S8nhemnM3mTW6IMNY4huHsw6VLy
6u1fuYHgcM4SXoUAgk/OWqW0fKlEYkQGXBg8RnE2Iuo6B4jJFEC/Uiocc92nJnIE
bFIyz8OhJIQMuvJjyFqiirRYmHbBCseiZ9cgfF1M30vPKC/ekg5s9woUjP8N19dS
h1q7VSv2HMCewzV3LOrn1lL8eOd1oYIo20Ohm8K/o/2GxCT6Te35oi1VtKC1ue4R
DALKqH5N7gGZnDvDr7pDmC+ShshI+KURaFZIGW7mk2/R7CIR5J8il/Scyui/+4/w
nA6L4sxbUX3HykF+CSn7yJq96r/rmB0hcLU9dK5zLOEP5mE1sCMFnE4BPtGf8Hdj
uW9gXgP1IyIy+ebZpzFN8p5dETkf+r2PfUVv2KfCnaw3UCH8CtFSFUSUsMUYJrBO
vMtN11BgT9NCsD9u/o0zNiSwnEBTrMvd4ciP7M8tqDc0iiaa5QCRTdSLlJ7NBRSL
KjfOfazDC4Dab8a+KftbrEv6PK2pmJUBsfLWtL+uboypGjEj0m8vCFPT5HiWbcRa
0voaOjXI4CTNiAXdmlD4GAL4Djo/TXeb8oClOR7VHkj2IpIL10BlMzZDBDnjlcHk
LDuZnM4oc95RbPv9h9L9Og0SqTIvWHg9R0gvaQ3Gd5eHSKFEorsL4Xcb1vaNYefT
P7NyHEYwEH0TRfw8nzNg2lJLd3NMCiDLJXHV6G0L+qeUV35+Kgs4csDjezQkkIOT
HdAdUGdRhXQsc/HGHzOO4mGBww9ENQ6hvjop9No4i2qXe6mRhs1FHNaSh1CscmQ9
Ld5aei63tVjyxrjGdLUPNGAKr2nBkU38tMjIG4nQfZP4O8y/AquO/SO9JdP4i/Tv
cDn4qgUwZ5X7G/ET2RE24zQAwVJXTDNiGdebpJYwlsHZkyq/r/fw/WaN2vIhqs8C
10vNj+F87vT5aeF7DWk25+fOubckZr6+jWq6ShAsARwuuicAgrbyI6ScFyhFu3ff
ezzGXkiUO3tutrxm/IhU/bvOzK0DmbGnsw1p4f4OhT+BefzeutlEodiv1UiVZ1ei
84jVJGBOS74a3rXJ546jn83IrYxbF/fQiymRXVKxKUjeI5OCdavTtx4F+UF0mmOf
8EdyWYCq8yIRkh32jAX9/kYcASfM+NIYr6b6DcQs2c9pbBw18fre1MQVphbdBYYN
0d9hQNOk8tifdkOTP1U23oMF6xJLKWmzs8S7kYfj974xaOClGidq4aHQUeBYhkvR
PMOQwN8d1FGA3aZy8c/66MmLRISKTzxLFYC5gb59WFffQC0+W/e9wWsIfc9zYG3N
HhVP4Uw3/cseZ5zE5nYWzQL7J1FjLYdd/dk4UrKmfc/G0KxG60OCJyosWTtJkSbT
cXmVPNL6g3UNMilQq2YXi6Ew3GN5/isrrvBolUKZyim7KSiqGnHew81EyOK16LXQ
4kLe7Mety/r776MCJEsdI4m6BK+8aABGAkFwhAjyjdjQ1SjVg65+RWCMfHPdfoE9
+8ZKsnhJbZX1y0XY57fLHRiNeiFXUh6QkutJJub5Hyi4Aivgs4e2ZV/w2D5V7z9f
EyOI9YfpSUzDH24FByfC5C3ICr9o0SBxBfMDMEpP9hf3xo6Xt5CBxaIr4bIW4TuV
9bqvNmg/SiIttxp7oNwOliQmL6Np19+lv8TduB1YYBO88h8O0HJiZ0CrZfAoD52C
+ZaQLrp1JtDE/oLHORbX3sHfHoqreZqN0Cwc0N1WhUpqX8knfeorp7CW1tpPCxw9
+BxfHUXSnrm1pZ+IGr9ITzf7GT1UfD79HGmbJtGYr2FzuDpHIfruH/agilnWIQCL
cY7dGvL8Fsqb1yA2hKlmGoT2yhWdbmQ/nyoauNmzfYKdFYqYIqskk+et4xSgSRcm
lQhy3XtBDv15L3T1FiVxFaqk2unLW549HLzE4HNeD327PA5WC0m7KvAhJ+oDY6Sj
GGvHlVgtSdy8xjkvAK8g1LhKOMgNmVoMsoOJmxcWPNxDv1uFWr5r5fsuyQShPfAz
kNtulFuulRhneIZY/D9H/Kq7i9i1/eqqFaHAGbc3kHb3FKpUhqyn168BcmX8QAyV
UkEX6/ARsRWfIqV4OSnewmMq1f0NAjAQMag/WXaPheg0t6CC4BlfNzYG89WcrsLd
g1edVsOrRrgzKKeT4FY1suJgznMiu9Ina+vO4OENxG+tCxXH8SD7RBB6xMVS904F
lE3DTpVLicmGVpKdQWZrFrIeetk0zpdobOdgDqDcm/j/TLUbytV7Q5XqHklPMujn
X7eQpBUSkUt+ksHZCE7V89H+ltQpSeEZBHncqDvrTVHXFEVuKI0OiYAiu0bwC+vh
4RlX0Z/KQ5CGffiDNAaMGt94OiZxmuQUBjPWXFEWXXPsDBAnWlvyzYSK/ApqexX9
DpRaOeXBgd+5i6Ot/TZ5GxeTHIy0Fsy1i3jz+PW7UCt2vk4IuRMDZl1rZnh6bzlk
U1a6Izu24SsePgEhgdaE4sd6GA7hQ5wMMcEj4a4PSz7IK4Uk5ladVr4NLCzZl/Gp
TfIqK2WN3SRwy2erpN26ROsQp59Wq12AKjNty9QO7Kbta0S3cgLbTzOZmfDdMUiE
RWig4YimquULSqKhU6XHn2udfdihv2PFhLVezfPKaNe4rzFLGmpUSjWa+Wc5LcW+
WQxJs+xVJ7NTmeFd1poz44JcYDkayEvuDQ4mnnyeirxPB78LSfTx+KWpUb0UxFTU
mliG+KGE1Bn/xIwDKHgcY1eQObBptzFVCtT0c/lHMUv3iaEfYzBQjPATe6A+jQJd
AyQvUZskd8dafdihsUveCH8IRX0jHho1AdrcqL9c50V7b93CyCejp9J8/LQ6z1A2
Ck5pbqDHYck558V25IpZyJAOdQhchDUMUzoSP4W6QpOTAyUnYyBy4IJ0rKgm5ViE
OnMlJwz2SYWLR/tCanHBgph2zd2h+m109QQxuGuzgUzi+iCtj1SW9oAIcgC7mYwO
U/3n/BUNG7FvSx1u1d6MWvEcnDH4q7w9dyXxVB0bOLegP20agz9UdbvF43jnqKxS
oOcWxZeGlSfP1UWPUbueVlvamf1zhJoT77Qq0RVe2qfSSyxemJVGjg6J7UQyahES
+GqZz43tWbLNH/hPZQS+mG85Fwh2b+MjxffCIgVx+pvTnwdJ/DmkR5VFyt8+MTzb
g0w4VI5XYA7hk+StKiiXTY5VnUZtp9D4l65fHxvR3VNiOo5niqkHSud3JkE4THWl
Gf7KqNXK9NmVTNzdPPXEJSaoN/zNxMPky9uBKTx70x6Ig6xkp11TtZflmG61kV8v
hAxRYgf9kTh8U9ZEVmlQ2crt39rT5MsyRj/dkfCVw0T+0J+TFkF71Nhfc5+7knJj
LnG2RN/k8cHhocvzX2pZ5Nu1mTchr6EHzP5vbGfR4MtwlA3PsogvEHXtcmCai47M
xc3bqw4xD7kxky4+wPsNSiBXwCI60I+M5TXGDTPFvVleykR0zc1/F8yhey9N0j1C
YGc9b0N/+V5fzca/jIgpSSRgwurTA5dHezSwKxLynQ4SS4eTje7pHLq3KLvphlwJ
fA7p68oilsJULQYyrQdVEI6m01U5IqpPGHayIoETp+RWEzK8pTHSeca3PmYG6aTm
LRv3xV2UVCdFNvfAu6QEQM+og5Vn1RYUX1sKBIsggvPh+45zcJGwdILqyl9HDTbi
oLpR7MTobFC7KrkrLwmsh/XSHgiAnMABfD1O0Sesm0XQaeNrUVyRznejNiH/v938
DrmshzEZirczz+N41w7/MlbbBGlVvL6gmis4bGVyDa9HfR4ApNcCJFqhh1QZiFwy
22nsH1Q+YR7uSLLNWTQkTJeo6ndVzgvfLayzN7y9qcsRJXstK/BjBgM4KIOUxYi4
OHU+u7TaUvDa+u1xC0CzY/DoJFoJftrj1x5jcilL/wi3kfFb95OV0Cml99LPS9jv
K4GZqcVbZl+dlKb5Nv4s402hB0R1UdYSwSyO1J8tYinKJSNsVXMUH7DtibbTjF+h
pU8DIsdsJnRsupvpeSV/qpATWXwXgRE9JcUhssf6tAclbsDfSGH1kNCxQFa+BsJg
pK0/sOAZRKhpDDyX7CPr9qN9ISlJR82M0eyLcJGnCpQWvgYKX2zqYhLdMlUq/Spr
SntTwwa1pPm26gJKn3GsHmVWHUmQlxfz9vEKsnDl20pQN7Deou316x9LY+SzRIPg
p3dLfVfbALxPOKmkG1aHSMLFDpEOV7W3ebOomzcKlYWZ20i0uTbNvwXfziD9fPxn
Mr8wbkLUbUGV8hfKz3PEF5PaZWTVDg5Y2pLa9a9zWeUAzt84dLMKRoX57GllzYtw
t8P8Mnjx1V+chShHDu0WEM0gcR15mQ5vqlN7VOPafacl9N+5QOBMLaZB1xPqz/fx
ykyIWgp9nhpHnV252NKw48dbVY/91l4yukOjULP4t06IgJTffxFmmHfdNvKhCPZF
JUDyLkgdT12OUzIPaJF9ZFe7t3/aGeFnvcjJo8O1w7EWRKzzg4EaPNQGLvW1sh3o
y1+ta+g6le4bFIh1NL3eSQ3HWj4TerRmaH5W+AHINkYrbujJdwm8sB7f6JQ256lj
H74n00SIu7kTDSWC0r8+Ql8TBZyPR95co0UVOXzVyXBjkcQxCDVSLNLoQdY4triy
1kNF7tbT3a5DZpjGU1b0/lHZN+6s7go8PBfh/YTZwvc6OrDcLpCSR7kEde1oMXv5
r2xUYA3S6dRMErqj20CrfZM6MVGndBRjJqhadVEhnNrfKrMH8WNLqePG3e1I3dCd
170LCyxuBEjAlQ3rSp/wiNdGNrvE8iLz9Ee5h7PX55pyUA559A9z29N1RXOUmwnq
yrJHUS8jcfHUhxMkg9AQWCuYGar1N2sGSh87HBJ9ae43pMO28tdEL2MGXxDO0a00
G93EeZihZPc34SPizmMcgtJyhE01qHe9sPGAKvPeo2Ak45Eb1GWYM9nSIR5Wm+yj
ICC24pNn1XlJHRop4k0fjBSZYaQon0PFftpBeuTE2feUoa06vUcPUpy3xRXY+ZF4
aaun70bEGsPteVMJVPUmOjvfpdiJNdaXW3o9VL90JZuVfl5t+usOZsZntn/tiK5J
mMOSULXrEy7S+2hY0jc8pV4TJ21OUd4q8+TLf6bv1LUiF/mTIGgWe0EcKwaTqhqX
LdX6QIo+PE4imgyiGsaBfjOrWZ9iHcJ+Qo0q/F9WSCz8fxKFwaB6GdoSAPYBZeU2
FPLaafPHFRGnuxXqxqyh/KROcB0zxOdaAcgZabi51H6KeMbGY6/rnouvF1JkWIcI
0z8FKn6l9g2ZctnoBc3W2HRROyMCstCf0OkoWSxMRpFFdAOTICATDYornr+qTHFp
UzJ3taUQSslMbpiJytQjYVsGXkRG9S/9CZyujVv8/wXQ1F6ThRmkZHKq2xYh4LPK
eJOJUzplVmGQOkiYOqBYZTFA+IdkxUKLt+eBnPpDUmgRyxC+B9e1RiaWef2Dz1/t
vgMsLocvoalaBju/ASj/xGo4uLNu1zAJoB3ufsO2fr2B0SiiSTpA2+8Rt4qWLIPb
Zzvki1dku3MsvmGujbpSSx2aGaf5UwHa+XZqoMR4jMoqzABsb7j8MSt4eGV1Vb2T
Lbc7s6fPs12U3p6FtCfzJm7X3f1whjmMrMgpzFtJUS+7+WDjdwTaxV7+6KIVFynX
h/oJcxXc1cm6vojy3r0xbl9Gx3KYqqF2xwExetBdvQVtI5LqlBS5mjK/doBDJ20L
kwC7AI2rA8sBzb0JQcgi3qagfAZBQ8wsszR3RnqRNtTLyTOuSr2eoPKJEkVDkV1m
/QXJDld8EJp2X5qzgKKE6vsjnTg1YqJP2ARum3UKAcgl1TUIXJapTnD3HDYBg5ii
ZSlsm84s5sS+FDqXSWWsWz6QNw3RZm5ljz0GYPCHernac0P+kr8Omgxnrex6Bszd
jPXidjOXYj2CxdvWO3NaSVozsYRZ/4Zin9sM1F1q+t1jG6mJDT2HjbzWPHAvxepA
MJpbn2CHybViQQbf3qchOOJfQYgMtlV7/rLmvIk/wzyEybO8TI5oMdv+lzY5Md4r
FP3JCu7tmW4wVwFvD653XUaeKBs5enMFyEMRanBZvMbOZMiXBbNwrYbSu6UQ1kbs
hhBRQh0v5fszF5LBEodXkKDI61W9vtZJ2180/Q5GKDK1TjJKi0d7zygKlr5J0P5q
DYo1DT7mNx9Y08xxeq6cHYQiFCJ2KOhTHjA1/Wkdhm+sJAdtz6b8Sifo78KNKCgf
fdHJZrm9Z+ZXAD7g266a0VeIlccSVHAdVpsNc1Du5yg0+mDZZrfTtQvSNhg/wAHX
7NF+Y7/MmQBe5KPqb0qOhfwIZ1my3fzwHj1z0JmQo7pJ/bK261/n1iG+jC5NdZdH
OY176GXH8BuM7MD+ooMI0rKC5JsIAXi4N/3gXyKomVGiua1DUX2FzkYPl6WV/RQ3
ANUcqufIeUEpTYxx6Lq9WKUBMq5eAkIc7ZnBAWQAAO/yDQsH+LDRMeTleFiYYAN/
TtA444Epz8ELSsxzpJESiJUzaihsiEgclFX+cYN28h7/m4AeNr9gcYDVzDkHeSvf
XclC1szeh+HvsHluz7Cskc0lieSi/5FI8OAyVTMLWqNwGN+uFFeTyZiT1RrZT9XJ
Zw+Zege8kTP9tpZSj+dAJJmyPYm45SVjr5Gyf6cyPPDErS5xOs5n1NgSoJjMN9yU
O/5ILTJA1hRvzOTxFsAAeUCRmQgNaQIQ7W2KijMp+7uS1pGm4NjNSzYz3tnjUEZZ
TgccScQ9bOB3TwnvvUw+4MR23qyBlEJ3Udu0MK9foiblDupFR3jqLVLRF3coeh2M
1iXAsk/YvOA+MwBLEtJvq9Z0HI2COsx0Kk4AeWlhxaSXhNrGcQeFUlsgXJJVdxql
notHhxszOBEJA9N4qBFYSdrY/dx8NRmNR5XXEwGAeoOkPi61ha6Fjkpbr5FEC3eM
BfvVcpxFVveIU4sN9AJCsUH0O3sscOkCIy2XgrU4PpNRbUgahBWGz+b/cPIQdDH8
Axenir4aH7Deqqlv2bnqVNLnIWQqQyd4TEB3P0fE+ffuAKeL63LqN5D3dEYfqJrB
tKOhPLxNuM5YDykU+oAGJKukZG+A9y9WKCOo6JOSA7xLNJ3fDhrmd8j0Y/3C+Gyp
BnfnzuDNmuKqCph4+3bggcvIlEEyUGEO94XI97r+U4MSySTAWjivqNQGmh/J+1nW
037UR4WUS9tWYyNzlZ48ZjkiglAywicj0dkTfVRZZD44tHD/9W+idDlxS9Pr5n2u
C15kjGHpUT1CPD/AqKLnphsXM7ufVmgIvaMxkZpKxuuExpEeIoiwl1oVF5T6GiST
RO5+DdCgzkhZ01h5jQePJZZlHPu2mNxbLaFeb23J9VPFiYy97m/iIC54EQOREy7Q
b/rugn8TEyzjAa9y5D+o3ktkqDh44ucRhLTXxCHZMBWgMT4SRJz4w/Iy46GhZZdq
R/o29CpiO/MMlSg5qqTA7dVNk9NfYDTvhiOezFal5woHEyZBJwDn9BI1pz6bUET7
DI/7Z4Jz/VhkY2UPG5iPpvRQ1vihnMUxJjGNPDy3cjXABm5eL2dFHIBWtNEiH1a3
LFMnt0bxROaAfyiQyoc/QdKqQX7M9sIiZtg7lFIZPZgzMHo0GapIsmW1iwDNl8aA
9AXTNyxXZoqtWnQzdSvKlyE6KwY1dev58QzbqPwGhPXZlcre+AtY7RhWPu8+cd8n
XyecqajBTDys1kwriqwjoy5UOtIPFuevVhSa69F0MW34x/tMnGVXG+8Rb9YMREu2
BQP+F5cfhB4d++zp+2ocUaMU6XMw3J38mgVHg9KOayQY5RcUkjvSrkgnmz4/UVpC
kCCq6r/A69fyLLsgO0xn96BCy62tqqhhdTEJHbMlNJlcOly0eCcy8jGnrcM2h5kH
T2rbErO3+mrLiAsP2rnvtreCD0Sk+RHBgdqlHfGn2J0lT8twzigWpNbToiXLzJfi
MRVLsQMa5K/HoujkXk2v7zq5VxQPE5VIbolnAmv8fApiQrJW4NKN93iwgrFVl14G
ThfX/okuBY2nF6/2OmAZavQKaTM8Q20ZiILAdfhMTHr4nkMRnUssg/jZJy68Zc9a
l8A4/9Uuz1qS7kVSGbLNemqctSbnuvP0ndU6Csho2Z9r27f/QdYNqzYNXLjekGMU
GyDiyzeVYBweHco8XxYEWevmP2ikXGIaYsE2kHk0Ym7evAiPtQCQMZg0lbb5oO2T
tsDokk2RdNZNv/h6qihQzHsyd3vV7c9agfmBXhHc5cOrhuPczQe5/LjndyBrxDZ6
QJi11lZCv5nc/IMoy5lW4A33m636xgNr5PHlwT+0whQPDOMmJvpGG49gcsm+Aniq
XSv+Z2pa5Onpx2gK9Qp5upO4XuaPMjbi306LIyFqBn/1fHnJP1bcDOKw7h5BSOGy
H6kPLKn8yNKXbr1YQ/eUlq5NLOcOHeo8fph9+kBk6mtucssgwcjWw+EBPFahH4Mg
Akh3DcqblZvGA/8kb2UEISTpNQLO8vpfTCkdFtTUg5ux/JyBmYOmVfDyCxAfCLDC
PwktW8OMtGaOxW+vrnF4K8B7j5BWIrLSsA9F/rsYAO7+F/cxLl3Wy8t8riYRz9d5
Ry89nrtMHoRWaSp5mzuOozdwBStBbs1kCBI9PMS4/ZQL4RoulaXf/wMF80z3MVAr
qJJ1ct4FitTdoon0NSOy6QlkSmY237MfsZZX1C/U5Je860CQaEBKk6kroMhYYatU
M8TQLxA1EUZ4txT4QjhAW97OiBpQ+PrPdC/f5muyj0Z0gpENeFgChbHQZ4fIE46N
ET4oSvWbEVKdAE40sE3tOLgi2si2TfpSFNosmv55UEEEm7OEymfK4bn1fer/oi/U
VmDQVIWsbIEGa+0VE+vLo51YT0KBFtbO9S9AQDXqgkjCtWeaRzn4uQ3sOs8k5bEf
5Az8rs6V6DIEy3j7DPMV6MisQhg8fyvT0pfy6R8Va4snbduF9KmupxhlGhQ3ZbnX
3s+AYmn6TmYBdK/wdMimXj16f6Bk6SJnRBnPk/PHyE0lpW+OtBZLnoqvPMeT6Vmk
tMdmS+bDh1b6NaEAAtvSDYhe6W0Rvy3B+yI0NAWY1gcoPDRdYA7xucx4MldvVsAC
eVH9VwXLxXAhEr2+ErjmgDpLid87NjoRWk4ZxcOB/po+bTb0XIvIBheY5fW94vVO
J1EoYCBEYBKPm7zRFeg/G+n+3qm13Go4uHPi+RK9BWQSftF7F0sFbROI86X4N2Kj
6rAKOnyn6QWiylhpMY+gSb1kSxPC3FN8agYwKTqcjnVX581Janypb402+ZumZ7iD
UTOfSpdh4BSluL7YFx8yEE7wNi28CznbyFZT/IfHK11Ykue3cq0wVPtPnV9EMOy9
W3AcUe432IgOj/nUDLcvscYiYnKFVOR5WphdGbtFd4Upv1frYbgnfNvAqCaVL6pL
PLAnUDwa9NSn8fdWb33kJkferKNaEAzfy7maVXaMSS4rPpkGt9r8Ry4kBeAuBNZ7
LtdVJXNJEbeWb7C4U6JrWeb+lQVd3iuas2o1ctnyfnhUXeGWeWuFARRAXYw333Qe
JRyP9EiDn1lUdXt2aTS7VgJIKBew/ksU0C7BmCeg8Z2Lxc4cDLzh9vbAOOFWyRL5
S+5YmtmTtASnp9LiwFzAcHYNQCu+Ph7XEEW288Ug5CrQwvPxw3k6zWfHnmMn2P5y
GTCN/AcShctr8nOD8iIf/Xu4XApKaji1S0ni2lnWAD3P84fLw9JnBhJv9MpwnYOu
zchWLMfX3dKELNIWsOxI7/JG/2najmqPjJ4sQfV5bGMv/KlaLDPhMqpe6TNEuj3j
FEOSxf01Ro/ARjwuDDeTpjxrLpgDr/jFxavN6E/BHKZ0IZB977OCTZbZEEz8/Ycq
SANd1cGAjINemk1W2hJM9mWl7b/Y2Ifrzi4IJiYm6Xs/Ony88aoCNJBoYx4HxHTU
r9qrjYtjO43vL+w0v3dTJSC/UyuedrCWX2bIb2eoKcgpum9xNJrDb3YdWUtBUyjy
rrBz0eXd12tboXzxsXyuT6r5FuVuc9OX/mpG/1sPz3QNv5YX8F/VagzgfAHxbbfK
nlZ5jdZwK3g16fUXOuBSTuC06wyoJOZK0LLzKCyEBDgzrloiNBiSjopSve9SHcM2
fCu6RyoydnsNDUMoCYyw++JmT4a7M9+fVODnJg8Dr7CjEEsS+sIT10idBceAUO2n
hmJU+RhZQ0NKhafPfGm4NIh6bdlYy+qkMCk3XWouaaYSVLX5WatZ0YXXYvbTzYnq
HTLmMlGkJeYuSDzQz2JCKP+wRoSCroEiC5WpBgcucjOEn5gjpNTQwfT9oehQmQhS
qypQ2O1IA+wNKPeljc3PiXoqFYs2nOsmCGFrDMoZb1iXWtCWSpS1D7+bPrXZVHBr
VALDrQpNMrG2kTC6dHk47Nl/WBRuAKMJ1Q93kG+wfpKJnHSWbqECfMuspPNco9YB
3Vd1SYPUiEwEcWbeK3KWNTZLWAtKdvQM/QcI2Btr/zTGRvw0puHCjvzDd8swDHyW
LH/8oNNaF9mpTsijilWwh2KML5z4YjP6NxlGyPLYwPl/0DypEDR9TcspXbc14zLY
K4mb9nFMvMglU5abp5i013YJsTjGvKBxwMbhpCw8ZtErF/RyQJf40EyUWti2VnL5
jfmAOmCUdpetBPl54H3b7jKdG0p23OBqNA+SXzZ1l44S37GjDudb8cvuYECuRL8/
Xgydk6DB2I48Yjd4gV90MgWzvVJVaN9U6Mt8Detu4HjV4imaXMtmLRANBL1RPvAG
gnAakAlugyHGDQAYVVpq1BQzjg/b7Cw7JoQ49NJLXfeYMiKowEyTPc4Veh3nuIIm
AA1jt0anqxOAip1yG1CuJX2UCEX0rq2KJEZqiurooSHP5wOe4BGiQOgxVUSHDpLe
pPYsPYaIb5gWyOOJBGg1qnkmmgMJhR6Hxz6weNhysCRPzPYleJMnn8AAze6XC5RS
96sVMbodmlt/IsfA1IOsFHxlmLnx3sfvAD0PBKm0ljqR2kG9dacyujUaDTZjeG3q
EsqCLxb850gbmdVoO77RaiY9NXVPG5rm3Ke4wy31j+qdhjMd0iQZXq8DElLgHdTU
eTWFnmFB48I6nLuB5qf/Op1VaUdry1Wud3kSJDsWl6ncsHuePc0H5R2a6RBNIUFM
4o2QW3wGrhTxpGqDdGU9aVEP3QTBNJXMZBMlmlCQYroz7NGuAy+R4Yk4wKik1GpJ
ySV/yOncUl+bi1wNFkbFt+W9+Pu3vGOEGE6GzU6rETEP+jSpmKTgvLfBoJ7kdkDo
7XJF2HLXsyzZQYcLKYJeI7orclL8GidlJ8MJKVojv9RgemrVb+l8v93PsGP4EwG/
yyo+fTJ7dbbCddKlUDpRzpVv13g1HiHsv9jIxbtg2t8tL8E9jesddr755VBk6HbA
hO2T/PJIn4KEZsyCjb0T/0OkzNitGKfjR1D7BVv6q5N9XISv8w2Q/CVoNczUNybB
n3pAQj+U28fScov5TQfoQJbIYbd5KZ8sFN9U9AtT15/h/ejk3x9uJekwfghU/ejz
GWc8aNPNJfBDRqYBBZZhEQof08BsL/S7dnVLcj36keanEypnkBKjlwxVJbWsEQvh
81IE4GGizb8b8j5cRw8T0+HwUGBm1VM021JrKIFipNyuerKndAOXMfTQ2r0xHPLV
qnlmUCD+J4mJjesaM1Ss65JwRqzldEh8MOEv1HeNHAC5zjh1Ms5sFWkp2mn6fSsB
o2me15gdufD5k+Vrd7lB+QMk10cvgThokwCfpwYoZ7q1g/I/ozZ9Afbf/RfnmV33
Vj1hw3KCWUyMMNDvvQnnUag8IUz2J7d7+G+arLnzawbIQfkm2an/7XDxG8byQMTX
3NKS2p5pV1Ojy7iXw1Ezx4FApVuJZeH55goJLS9c6WbrLPY3I5HD17/heRWJvL/N
yLF/dIwNkfRufIHeJhqcfgneR5Kb7IoKOmKkCKgOoVmTRovPalxyLGZGFDV6WkDf
2bqdfXq31clgB3jzbkoNb6fjhjJ8SNBn6l62LUBzvSctuEkYh8SAFDJ35IVH36pz
vt5b7ciMBDwEKJnn7TOvu+YEwX7m3uXYkAGB9TB1EPxhdgwMLumpXyGf7zchVsqF
NIj8Vfl41yYi5MsIm0ko58AD4UMbpgZ/st51hVnkCOKpnIFLQauYyFnalpKvFVSd
8hv/SJJ6qLUFWL/mZtIj/4XtYjOAsAX2TkwS+eoWUUHM3+4FnhgPObrgMwzJ1Obg
p+twECBrHv5dbiYknZQS1bo0u8GgtXehQByxEyJlylmoy9oRzNQT9dUGpozEHfaL
Bvrz7ilzSgtUHGWDe5ZrBvzOYHO6tiqfco40+fXGO7RylxPJYjC2czTgTHV7T2wx
b/E8rTQUquJJ00MQO+ESHXc9drWs4A+FexY0i9mwTmKcyHrQvTea95pKTFl8UkUk
jbJvLaX/ht66Uy+9FWwpfHnSmJUakjy79J65mRtHyRN618VYu8Bj55rG46+xRL7Q
GX0R9KhYvIruyMsA9+tLzTWhdI4uXcgdd1SHoTRIx8DdZzm18I0mQjO9jDaSRGqw
68FevbyS2TaHn0geOgKe1Ygd1bvUsbBgnDfjcqKkKJQcCrxdjBbX7pAyR6W1xm5U
HWDX7zmaqyD1fxtPzE4pEBegm1U2Phn/BzSWg8Wq9o3avH6fLi1omu61tp1SrdZS
uee/PhwY8la9CHlrdapCfeqhVYqFpifBBsR234aeBBuw9aVGsT9fZKQqfWGhASYx
H25U7cdjLm5+IvICXLHys2ats2CNFq9z9n51HB+ZAmmGbzvFlRIWBD2bnpPYAPsV
aq4E/Qk8lJ+Lqh05so3Ogvh0bVPDSSUJUvlj6LRdjZurj/L5l/Yz9zE50moZxMAv
aoBTNK9uNWhfl8Sb5KIQyNH5SsG5Jf3Cu0K5k/jWURHl9+OV/jkirWzw+8xjdcZK
vIguBz2vVnsnbOpitdYxaPn6IFJMOlH6qRA81K9bvpqPEAUg6aXrL7f8fT1aAVGT
IyvBYJ4q3skbUvHSvbfYprWjpP+m5Sqi3e8/mYh3hzfWKZuaJrQQERba2/xEaNGz
u9XhJcyYb5cek5W2JZsA4nOJAZYwB4RCklcA9RKgGPDUUmfKwK5Y/+WZA8bqeXpE
3hVCj+7j2Ja2a9tfWbZ1HI2WKmntu6dF2pUErHe4jXgcGKtrmvGMfy1RxMtiCMdN
G3FT97N1VNOLrnRxcy1+zjybNtOvQPggE9TT+FCJyx+w4K7JF6w15opnSmOSQlqe
jU2FfmvnpuhBFkUs9KZZWPnEH2uECEgd530QToY2YKl/lD7POkoVk/PSByeWS89V
6PETk1Sq7znrFLFOIpGK1ZJ0OErZI6Fw9tQPSIQm2vNOxBwWu15+UZav5HXvmnSp
4/6nMfNhq/uu7G6/3Z+h/bIpiZo+5+3PqyIWwkGpaOMA0LAX5sA8VKYVepWOhoLK
lgJmAUmd36ICS1XEiMATiN03A9d8kQoI8tQ40fXg9f8g4SJwgXAdHEwLsHcw3vb/
HQ24CzBKfq4blE4pqup0s14O2SHIAkV9MznvahKEQeV136iHfV03RmiH7QTurKUb
lGEiPDj/LhOVFGORf7gtbOcQsqY0oHweO7cQmERnCROhiEFgn1zG8dF1hYsv4G24
7eLrapScIta1xGUVtSQzm5u/nEcjBseeRY5kT2D4rXEFZIorsd6NV4FwJOnm7wyB
1xKEstlDCOOi7WQumQzh/FBTIi0E0FRi+unil48ycfoLoa/VctKY/N/Qq/pEkj42
qjVf/PU37FLO1Rr2xISUSV/D0Konmk1hmjxf+cmG4g+HrmkLCSANV2pA5EjqzsFb
52E3F1S5L6h4WXS4ecmMu3TaPx3EJdgAGSigu+ttyyRzxmzlTFUcJCujqREf2xYm
kEP/AC7L19ebwP8vGE0TIPjhBJ1e6AZ+sHfzh/6+ASRJpIQ+RMrknBqiz88ElvNy
2dQTbJUGoRqBgkn8zHUa6BC/HKryOqIR2OLl/Hv8IVwaHb9kh3ej6t4PkjnH7H1W
zT1vrKzn+QUPaObh5TeT7UUVc8MSRIc8hyLioqv12yz8LeJybb2Wxaogg9Ge8t7i
/VPkbzAHL87rS8AAGtSHm/vsaPsWJqBBQ7HexFO7p2c63H2q64JwhCV29S/jxHtN
QbfK8kM1QNjHuXBf1GpqsE0+9tJxkN4YsHdX4209ovBYIIWt581dr1iAVaxpTLTQ
4RSYrDtMnfOhU3ieanpRnbucoTDIRSuQudOD/9czkxi1iedhNd9rLPiM+Mjwqtgq
dZ4tdwaAQJMxCsZe9a4kE+5g+1lpNhthunOv0jZHChewQR7d08g3Dc6n4tWUUgzM
03Ew28tafo2+vYq1MzsCbe+w0DrXhasZAEtIiMYaFmA/Z9UATETsCvzs6IAX5lAx
K040hRnb1cLnztauipy3lrZ6jPcuSRZZvUJbpYzRfrbyegQ7cwvvIDrw4XwFHtUx
fq82OepCzdhTKvS7f5mp4+FCPBo4A8fMVm/iBWxTe3M05+4Hp6sVq2hV+BKYVT/v
rjPe0ZsZ1koKDfoTBbq41BgRJAvB4g5NZih/9gClTNfRBfxerYphOfWHWOdgXA/t
PhIUop1Wy+d3ZCBpvCHOOMYrFrRb+fjBebC0wvFB1JQxSy3H1QptXC9T4aRnV/st
ys58nX2IWn+ybkJ8igfxJUfviIYwvnaXZhSiqAc3HQffsI8D6lZHn1repfU4ZSKu
i1mpNQiA28rDYE8rUUOUVPcUlnjNBVztwJhVNd9hc5DH7UaZ5CugcVqQ7pIb5FRp
mw5waxdSJx6vIEBSQzQTqTByoDhIlDrQALDvRZa/mOA6nHLLM8unlvt8GVauzYkW
/rlhmwYZOkEKO1vr+FhaBjYGyrMRNmkehGckrwSTN7hmTNxTJmbskrVx97vKRISF
T+zZeGe0M/Qmg3d+haEhA8Meu6hAFlhMyin20T8nuO9YrnU94GgDLdKaWWPn0NSg
XY9AkkMj1IJyV3GA4MnYSCEZl/svuR81F8asMYTeHsBP2OJ6/ugkyKuH4zOHf8iB
V0cjAv09Wh7tfKBdq5XlLshDWFoe1p0tpZgyEDa0r0GfPgbBQVYeE3E0Rm+gO7SE
7rTT+el+AjwY9RiKFjebRLKjMj1ljgDhCXC7bZ/kIjpQhVmW8Xv6Tha3SA3Q8GW3
qA0ImVsvnC/YZYoi7fA2KTyhw1s1O05/xQIqYFJWWqQLwsBv6jPa7RVhjF5RQbI4
aXS742MJM+NgshdQDgP/ovLvP97Crkfc9YehrVzM2kYKmRnGLc82lgbsly5ehGbd
p7BU1K43xZsyXfjvJVn5YwONN3jFL3xVaQTeGWh2TiH90O8RXW6Qp4Bl9vHVLYiw
SkuI9RszxnEAeKpqNviB1iWiwcnqRUamen3fH48BNKHWajO7cc7eIrqaUmkRJREg
bnHHOn9uZcCdlhGeuyXvScSf6EIsANtdy5BDem0ogOqUjZ07wPm64Tvr11T6hlxc
fE/N1zAP5ebclS3F6aHqIoyZ3SYokRl/Hi76JJdq7Vf51XYxPugOf/0JRMx+VAQq
nzhfqMh5IVUA8uVIGwoUvdCNcirdSgXCvJ1XBBKG7NFpAH/Jt2laTFq40JMutK/O
6Frfgana0ULn/mGJuLTTD7imT7emULkkgqR2D81VCx6hQUTq6lSmaDdsetK469+o
/2oPMaajZ7mw5bpYRGaPri6STc1KIfZKzLFGKCywWEr3RTHAEk9cClB+Gie/dDwq
ZLF27zEHzL4D3Okz6NBPAzL4zWpt7uaHEcNhRVlHOFiVZ0mTavN+FqCAJK4a10bT
UuOFiXZBrCv2EUfkDv+WR++hQ2r8TTVJlsWZMUlHap/3sFMW0zqtN206LIV5E9SG
yDMoVXfYZCPpFfQ/KRr9IaeW+auRBG+kLMVTOpI7B0Yc/OcYga+OnLZoK7Ghm1Md
7QFgQDS6Y6+4cu2rDRiQg6nz4l2aRcFeKl1KRLpFhIBlJ+30gg4+1U4NKOvsORfC
1p6qraXhSN1jKz8KxUUTsyVybK4iuoWEn1Vhz5EP5RzvTA9WNTictmwaIaFVgU/c
Vftkng+IN3VY0NKihd0eA3fvqGwvnZmwRI5NP99vsXG506bjI37dKW/FD69FVN4H
YJT6CONd37z2lC+jVxn0MfhEWEdPX+kx4j5nn+fK2UjwVSxuDA2pbL/Gdpt+IYow
/pewi4G48t4PCtQ4TJcX1CiULUULB90qmoo3Z+SP0vNXITE3/GgmJJFGPUbQJJe0
BoxKj5NilwCbqKssx9qT+b+Hpm4fQyYmCWGEL0dywXkhlZwiDmgSIXm2eEJcSxNB
NV5Wj6xF3wCZT9NRDTbCTWfViXrvYeKnYcBf07PydH6erpN0opHnOooasUQhLbNx
K9uyvwkZTzNhhd/3f2ACfyRjiK51/RchgUD/24/mJO1uKwqsfMXJSKl91pyuBbCj
rd6CesSllUoduVuOH4GOGCbL6SbrXmv3VPE7Q8aNbwQiVMjXQxXPgu/kR7Y75zq8
6Yemi2X1qRaSZzpKWxYiN1Wdum+5oox3s7wSlTSqJWQNorKhG9N94/LtVFrqkYgs
9bfs74CB5yaAWDwFLUzxsaPEXWGRQb7x09Udy1l7DsfyFE7ly+8LFB3Lv75P6n4W
2KWR9KIt0ZFkXvG++xAxK0fvj0hHGzlVi/zEskHzSMH6WGJLyZa/ma/co/IzYkAy
9O8tZ6iUhUedJ6osG8DrZwmd6PzaHRMTWD6YymMxT97qka2/02sses4LdlcosHnO
DltePFJE2/9PLbi6zwEklEWVGPAAMufrnXwN2fBGF8SpBMzEUnSDXaR/jjQA22oW
AQo5215PTscmVnT/TBnjy75vIsp0PVLZXHgjeUo1QkgzrnyQcy6vx0zDVRlwUfwU
cv5Ft6Fe1eGApe9XA6rC8dnLtHUuAjGr/lUHKTuHrbVrt8TL7qXvXRA5wCBzuFao
2NTavlVlSkh7fbM7bHSMzcNqdX7nA6ek6qRNLZiVgrrpPo1zXcFwY9w4ZQeBVOkj
EO63wUuVSfyletJdoPqA+6B7dhsnKY9moNr5fwRBEPELtxoU5fYRjYbwxhFaE7p4
t4pD6wWSvrB6yhru0+01SGgs9N9UniBNymR9H4X/n1j8JM3+bui8omr2bSNopF2B
2iv2b1+96J772nmrcq/Boiu93TPcg7fwV0BI5SusOenZxt4kUnaW/T3Nywm9Ck49
874uLeN7W5hg0WPkBp+TJCZjYFcbPnPfLCSY044FNYV9wmIDOUKQGOUhmshTUs3e
O5hAjr3rs0Gp1qZxwDElumdFEwLTcGBToWR3vP1oNV8aOw215lHdgW0THa1VlDLF
/HUWrrc41l4EyKePU1cP40XzvvUSTGn0kgcLgN6W4ZOsUmDnatYV4nOLWr4OZF6d
79kVyH7J30qgtkp+MlBiFq93gY/ebrHbaleqbxVSSjkcnZd/rBvbNudXl/bn/sEP
pAY5IzMQSDsXyZeUYdJqrUAlkRelWYll4rND/wDttAT3KC8vUklgLlO/4tPxLZPb
/yeyBbSC/X9ZVZEHphfcR0rsrC9NxgGfegJn7TrHU5zPxaMImPmz0ajegDQM6FgG
ayQMT/Dpq+SPsezeOOxOq0D1BDqetfYlHrEB1Cet6DVsZV4al5qYjh5wYc+W/fIJ
MiOzEfgEl7vh9+nxwLrzEqosn+DVayjnHKDCkb0RLYTbjOxx5tshsETnh2u2yW8J
wGvx88Kai9/LGOPlkOPdx43u/DGmfdStM+2EBncRUaMDF79zBVFKM6nt+o3IjOKc
P2+F4NlZQIzdMCGqTIjyQa8PBRRjIugFcm1g2stiwJjBrq7aB/CFNYfPFlFDChu/
CBZElLTYQt18mLUUbWec6foeHWZ+0dAV0+djUkPNdMrggb9NE76GBxSssjBEVyDN
0yZvX7MUcaHb05ldzHIpnAWvO96iKM6wmBjh1gY3kurnMw+8RR/X71EpnjenEpw4
7YyI76kzVuak7jt05IyuFfs5Wx+K5ZZ54KBE5A1/aBUAzXqs0kwPfFALEbyS1fiB
U7UrRL79nS+bKNdquj0mnj8IFg/pC6tEz3x7g3WhNGJPCxILjhJrM6AUn1O+jrCw
5YlpywFLfKlOtwTIGcLfDE3es8xOkc4qRO1RKZVZzsbQgcfwt/qAHP3mMzopKQ3b
Fwd65XYLFpE5y4Pu08sjeT0H9E0lH6GVvqD+5epo/RHvynJUG46EM8LPEuLq0SMB
7MSsVF2Kp3k6UuIjMUSKCUp8Wc6ThhWym3BTgVo/9VZ8fdSnu1LuxI2XEwds8km0
tH0KVsr3YMVDxoqrHEPA3HrFqphN/nwHkR16faJjk/DQxfI+HrRNI0njSYgDqbqh
W+aX1VHKeTo07dtJlIuffKd+Rn102uH2PobhyDm1G5dmYVTpIUAMRVRxVrXl5PDp
ommx26/0a1HYwm/QB6CYaUSFaWWSU/sUzEAOQzw3WGjXnxaQEkQiI+ZwblRq6HUv
iGl99YMGvpQioVVou1UkgjGQmphb700SvO7LI8PV9LJVfEzt0OashFmQ3U1so3GZ
+/1+hx5X6mhu0Gy3o1dzKnH1A0ExLQU8jTOedWA1OkJRBovsN7aK95RjLkbkcRNe
kvpTVQe6wqyUvi9JkZ17V3tZUJPtCOpfAdukTOnoxeMOwNroD+RB4mHnr8HfjS1B
Ep4lCm8ac2U+K2hbIbUU9pIdXID7PWUgmOXl3dcjD7SgTeEFhOQ5GKYNfyAjGWKJ
VqGwBjgiG306w3B7l+KjJjKh53dPxSvODPPlRAuSTc9pcHHwHh9LO9XkYXB2PHo8
86p9AciJJCUNOjcSZXyTVWy939CiZ5GJm3WjVt5YQvu20m2vSsw9t/o3L6KQYnqf
JD2kBLeXm41elJPH4264UvoHRCRc9VgEan6Ri+z+6SjsScPAUBF9k1GeC/3ipc95
IVcrZUQNRGbTEXfjnOoRzZnWKEASSrYIpSkjlwLhvPg9qqXrDmTHVYvEwsCxB6d3
XHacDikbuXB9ZglBoGOiI+QGnB4+cPEvsLZNr2o7VTuipPKGflY7AK20cwXdZFXK
kPZ04H2lg0QrOGhb6FUPcnnvrCDNJSJgpL1Q1AU5hS/158m/rfeZrgjfaJUv2Z8+
uNMv7K08k+ydtK4Ujg8shOyzW3E6A6G5joLBbd9TK2QLp4700EWsG6FzdqeF3INo
njVHu5FXkn8GrQs+dJbYA7sbjpkMUNmgPS3UzNh2Sl24dNu+ywCvd/CwZVGJTiAj
xvF/IheZI/vAPx0TPxLaZWKrgzmqZyni0535M7l1Dl9U2JNapzDuq6d0f7kTE02t
zp8Bm6lbvkKvb6Na2k/l7JxYKDZWSEGLrwmzMVMtSBgl32fXgJn3FRUNFMML+SEb
np+MQyRtKpzvjLHbvBfF576Nvd2CqKBmnMkOjUm84+9Nxv29hd7SonAHQXx79mg0
omCNAmxjgCr1VtmmgbmRyAJgQcxsajsw9QIFLwuq4Dcs7l82XTgsUKBBnzSVYLCP
NuNlrMRNIN70rGWDW/UnhAi6UndexpdI6eGksXMuwPiaIVBmn1WPh6u0ncOemOa9
ckuITTXQSngfWnPiBtkOeP55w2tS8GDdRqbV17vzGj92cJ1tupQOjJpcnaUp+AT4
CSZlRXwau7BBvyO9cANjsm4YPS58r6d1ENpvTIPnLE/vbgSJSDuILk2Z7RN37HMs
Qk67J3GfReagSTj6BUFAw4rV5fzZvQu+VAen/HWX6VSMgSuZzNlo2fiiVvTGAGqY
q2s9BP2PYHY4ihy8rjr/XJNbgdaZ7SRzAPRhh7gcAsAzFVTu4XJKPypPjZVBYu9d
KB7pkd8QvotTr3oJPXHq2Xk+nrswg/VREjMrCaBaY9kZ3TG60+NsR4Hn0gvWFwg4
kYbt8Gdn+5h3bUi0Uq1ItEkGUK1aF8rIlHwmwGAaF0ClNUFJGU6S9qMxWw4f2PHd
7ayiTk3GXHRtRu3PcoQZMc5rEXT4gxGAN/cIqaddWUvhKsXqJigs2ge33AhMISqG
5kqIuEeD3kz45Ko4vcpKehjFBWlitEQt2rVyYLSM9ziHiElfdIyBLxwICkBGGXi/
rKevk7pFZtDVTcs/lIAuAcX3vDhfCqMDzw0brXbzFiEfE+mc2g0NEJ/pUq65Hp0J
lFjBZu5PVN71PAVs+f4UdQvTtBJxDGv0nMae5ms4s4llzliR9RYpHg/r0rvF0eu7
+gbnGl6kG2o7bkuIY22M8Kf7zIjUrQVsf40z+HeIU/S4N/TbDzYLOlTKU8apqEjO
I6njpMf+MNEz0GyBW1DsP4lyBaNvSoNLDSz+tLzNGQUPc2KNnrBBP9k6ig93JNeX
oZGB0vD62soAjnrt/xRZ7x5N3+YZy/ms+3mCDn3MWqRdbsD+wMNnd2jEucHwH/F8
DdA141kGdbZGXFT1ZVTTGg7Ywsptlu0qrsdn/tKMoO11sGVr/g+FBMmb2cohwjK/
fGiCJyYmiJNhWi3A1hvwXTRxJHPvMHhWnNsCg/LjxvLq3BbkbufoOCdcQkGZ92Cy
jRMX8NT6Zcch4fk73kLIFklCPrerDQ9qILbaC3XM8UDMAFJ4kQLqhPFFEzYR1UZH
sMMemqmNWWQPgfol9rH3Uyx2jcKrKJGoBiy1d9rKaYotiXVKptimJaI0eoNgx7cC
HNAb5wRGJODZPEgtl4dT5Ma5l57n8+3Pv8LfIcxiWX3nLAUQxI4AiRyUgFJWb+M6
frCBxHUFrS+LheLASutzxMgtB4XuFj+/uE+/UxZdZhm36Y8nkRh+MroA7wAc/OTG
MHdY3R02/rfK/qHkTlNgh2nfw1AEBQg6PuBBZbZDFNt48Ug4fP/rxOZZH+nAh50i
6YUi6vS8aorUvVf1cZbNYh7qHT/Rnre2XYjfJL8S7w6nDIlVJU04hEPk5cCqqgaH
XHYG85XDljvczuWSyphH8FoAgDh2Y7qSwrDYDI++UBphmbt4XtDbOzUYQ8cUYH6W
FpIe3cZAPMs5HmYaZIyYmCZOS4Ul8jW1o4LNSkMBaTv3/fI4SAMXctUctCyX/LT+
gCdaj1slPmaqiSPqFJhXkDXt1Y49ZOOFXZ8IBodBnmi+TZvru37EDtSV7bkrIRJE
94pv6AmTyAkSq/nIAYj6fZknEofvZQy84zbDUb1apOHVouZ66XlWxDbgCKrklooL
6lpOBY9533kloHxcbuqfJwqkIgtYpr1dwt40IW/V1W8AJVUqNVybxwqFYndF+S7f
fgOmGoydIk+f6VCT5Q0/q1zWU2lU6vgsPqIoxzNLwyzHsnyjN//07ocYzdzKew4G
2Kr6eJgWeNNVmkWu0ZAYp5mLZeaivMs07Q6Q1ECCn3clCVK4WHgCdjDLNxDDmghS
aqOSha0zGZTpI4kxEot099abbJgJUPkpKY/dhzdOVM9+3rc3l64VwI3aADxKFHhH
FlTwftuK1W9OF4ugWKTwX5N8D6/oEao17i0jCZGXgiZ5gv6CI9DStnjn4cwFCq6q
Ml0oCbKLI81jxjh7GOH068j8FWeRpwlDh0HG43TylZvD/uwPq1REUYlKPRFA0GQb
h4db36wRLmrHoJWYWnDR65kMZLFfA4MyyDU/dB95ku04VnG+jPyKmKNO1kjECvpk
nr55Bo4Ee3jX+CZ39lgW5gXUPy5HLt5+Zught72QonHi0EbpEf+iKL3Em0EODyW3
x/0MVu6fPSy3rkUU59nDzr7cYVHdlLE2+m6rHV5egVp0LMhHmiQhjpqw6khD96AH
JT5gwjp4dyYX5uGIkT/xqs6nC3rRW5r7dfAMQgYST+bGvKo1+5j+RkqRGIWhrRAt
7F67NzER+gCMaNmDC54EFONp6V/1UoqbyOkX/UKTeFINTO6YaM3GMKaz0V6UjclU
VJkZItrUDmBVCvok4tP6sDumzCeGDomQV5t2fxMKJRwIOzeINLRJgasQrnHKwS7W
tRIvExA8U2podw0F/R/HZg8OzuYu023Ph6/Fjg+4UJY0Qq8lxcIbG+K4YZs0cc8a
1wd1CYNZMZndrKObyJXD5WY1+2BAzS8J37iGroUrF28MqPz371n+9OkLC6kyaeI3
Z6sXGkFIClDhgLXhWXA4dIjQLIBSP3nNww8zfN74jyuT5gAVL8No83s7Q11i9bqU
ETf45JsaVIWE6k9deGYWmAsZ0R6ZAESyOxBQ6/3Sob0irEGPJfwa4eBHAw93kw/s
Ewf0/7gF1s+zcQjbhCESUslhPHRTx2t6T+9ZAmFShOu7fAKIpLeOLEbQENT7kAQ4
L+sLdmiZLr+OFf0bfAOJKbeDpX/11xENDyAxmQObqb550CnvKwrj0xdGAD44wFgM
SOI7N/sbiweDp6wbwwt2jW0wvzkDBmeEG9ii8u9Az1yZyKoNj1tstdHmaWcuhUvF
hSWJU59TSZi/h9zzc8xhAmTSaCE9jUxY+w2+JvvVjF4+aiHFut6BYrYBe2lGgb4H
Do26kZx9UOD8UFoIOS4tzGIqURpE8QMHhfMLRGPfALoiIZSQRmgqoI8FJKc5MxWw
Mc3HUPj8sKwAvclBuuFrjgBiFPSGtZZv/Z2jKQJOee9MFkmoMfG2kgBkB8p7PE73
kkSwAFr2srLIOLlxkpqIC9Sms1jT03Qdu31EgA7mpHkUwPteAhwKJT3Z1V5YB4H/
BVryJ8m7J8XKtbrmJzp21mCYy096/+0E6YG2t6PVHsG3uZeYMMD471g/8pg4lg2A
l4ZQwIm3lLrWS2Xe1MZn6sQopSjDV3E4QKAi3PkZLxAyMJpytWjagcUYE3Ft+04w
TvL8dzhduH2oTZqweclbuAVSK/k5oJWq6JiHrl3atyRLsKQNZmv4A8x31vuFHTcz
WKHyGJvv4Wmyv5f84qslNXyELp+C8yWmrP1MQJOdofivyJgvmFJP3kCHjY5bpmdI
jNwCodDXKtWz69AloiH3gKrCJTpqQbOcrF3IB0myoTSKz8rfL0sTD24UKj6m4xV0
7E8IPzFq3SE741lrlewYIip27wXlRdyPE6oxidsZPboD89Ng5kA/gKl1aYfwfNmu
LwA7EW7BdRexaKuv+nRlmRGVExwDpAveyIiMMFOTYTxsM2IEEd2sSz3Q5iGrp3Gs
QklibhdWVfgh1a+i37RyB9YDiUUpc4+G1NXF+IjcJ/d4vlg4LuziURiHnCFiCyMC
qLeFi+QiDXw0MqH323P4XBIcSjKixejhO7DnXtAJxPurLl3fDEzYDnCubyhC6pWg
vnR+OHou8s5YRSTfZ9RV8rmWOfV/oXamgKTQvihVtCjIBCTjl9r9FzWPp4/IZVDG
huwNl1iN07HG0pvVhjomLZvL0ddeiKTN5M91bzhk5FaGW/LBq0eu184GbJkzEWG3
aeoEEC4RWZPEnz/LGdmKdy1KYSAMj+5v66Zmx+JIa7h9lZRh3IDqRMy5BDEppN+t
aB49L7KeySmkYp82UGhy/SWRBWb19MRAoTfcXH2gsnQgBKwxzlFWh+DyEe70DAH4
uD/mb3MLfKMThGvYtv05uj1tedE0l4NAcBIYRdyqP71rz6u9rq49jwDs2EpPcu6X
hscrgpjYnS8VdiAqk8p8Jhx9MoOMOotD0DEWsoxXYEAAzaa8y9iQ+qlMsrjAD+cq
PDHshFQet0XPmlH/Nlba1Uicpc68Wt9bDa9lIGmkwJfwSYDKx5p6eZdzf1OTSjJC
fnH8XKW2QcgSAi8k+Vk7ASR5DedPFFU5PVOknwP6R8ahj0qbm7flm1eSQQWsIbMz
//z0W/0NO1gQSwA4R/uCBLn1GZj9TkZLls1MrbOtlKUzyqxtD6y77ADL+y1eXgZi
Uloc9NcOsea7cEAjb6yIzVa5QAOVBimWae+GXguDv7MKIM1EjZjo04PI+2TnuM9p
HQuR/ZXzTxqLZczpishytEBxcCSlSmcRU0lrZ/46irfEBe8LNslDNJEv1atFteqi
mtR35qs7Ayou2KmowgpKSzH0XqEKDhGuMILfHQ7erVsUGz3k8E4DXfYZg3OquKYG
0vEFm/XHo2rjGZHFwtXRHFT3WlSkQ6YMkAagQPeRTSL/nPvAxfQKs+CXvtJmD6wC
oNM6niH+yCvul+GzQ2BW3BK6wP4EPhBt11OTp+2T8+0+ejiUBXjozW3tbGKbVE+7
arPLxWq/Iast5qxxxCazEhDZ92s6cY9POhBr1c7FuiIZDLL1sUIWL6jv4I1nj0Me
ZVu5YTp9l7rl3rJmfzTJsirOoyBu8lgg0PJnpeJVl47xnubT0Sk4vvUkat7IyUpp
MgHcfvoMh2pfkA6bcnyZWjFOcIpNtf7jJ3q+IbbEbNEe0ZQoo6O3oFK0cY11pqGs
RAlNecSZHPMxjMfPK4saE1dVDE2YyHHDoXnpI8bWn9LNZ3h6ARDnf6zkGaN1CXfh
FjKprdmXYJlFJ7aGg+HSPiFbEurG2oA91EBR1sTASTgQpIpSX6S8GQSZdltkZVBA
NS4n+5X9j1r3qZ6qlVGHUI5YXS5/TpO8C9WsKv+CZ8wYy0O37r4M5eOpHL1I4ks1
huuspNlTHR8hXCdkkAx8nBjkK4ksfuXcy9kfXGgVlkHVMFX6U0aKYhoLGVTy2cbG
TZ7Rp+hYaUBOZYAlLBq32jbnhpjK+0kvzr6UP0wHc9v+geWtYAfCUbSXaEFl/K6q
JO3heLey/Ycz0pJlXxH0oQdbG01tNStHhhuCoCmkFyyEdGSRRqk712OvQZ++YPF8
op+y4w/fnksedflD2NcFDRGiM2B5VmbgUxYhRa95SZtWhZIbrGE98eRl1jLC6ep2
iWgX/3cHK5HNFoZtOKF0f3OuUzqkC+Ypqv+j2XZYUM0CdbfWO2x8bbAmVLGGt/vp
ZHOvj5+R1WudKFUSRsfw26ZNuzPn+IhLVJNLMTNDRcUeHEkEstxqGjdueqNLt265
WM9dRBRTgR0snxli3O2XzC0pTZyihFGQKbvWUrqHdsHgB0rzg7Cfl3D7IOsw3ew1
S1OuO81Zt6xroL59XuCZLOttrKN2zhIULuiOGQ/F8RrI2nuhP8vp47ezQizmnMp/
Ht2YSJfzlwhIrqY76SjNZwsVpTpQWBJpAPmhtN7gn/P00PVHNmM6ktvIpO6rsynr
j/LWvwKENW2MuwstB48yA1OIcdhFZSO/ZCkZjeCfYOvMxDMvufSvasSYlixCFxIB
ESR4eZrz7dl7CF6AO4+aP2Jwq/I5/WHma9yTONwqSQjbQTNfquQykEEQDnF6jQuv
JCF8Un3Kk/opFaHVyLPGYX3tGBa+7nvziRM+x3CIWr9MZfiy0K+b0o4qNHk/f074
ABz7odeDAx52qcL37Ar/KWjNB+bxdcv86EJlcOBNChxMC49Rq/lsfAD1vns3Gltg
Lr2IPjt35mpLi/cAkK9/LxVkJb9u9ZTJIENIOm4/om9upvNHwnptjWY/KYda9Zqh
eeW47dOAsbrmqGJN50rvRCCXYO/cIZBeNT+ZW/i1GWiZwTz/9r+hsLGV5tkmHc4q
9B9zXj0FQjLiPGC4u0ijXNB1zLT9JVZo/d7sXMK+uIIP4weyHAyWs8AHzc03mS7O
3L/Lt3JZfkkS4SrMLLqzrIoGuTirFIGbze12x/MTAl6dDkphnouYUvHeP/GlP94e
gPEpYkKMJz0iMaN8vzfFFp4qhmptALccGXhPES+O4rQfMaFn3l+FJNbatlkrVgNF
Immi7MWmkGrbo3BMh5XCjD/+qMXds4IWKygLY1fExD+gkfmCCw8w6FeoJg5YBKIZ
TXe3fMKNV2NZvNhNbBMJfcEsz4SdS8mEI+sscwIBi9cuttIdRlDORjzXsDdTdpbT
0/+HBeYUULXV2Mof9AQLB9Si6xx5MTcIzDEdnr0kUDrIUJ6DrdPG8m/K3/wV+24C
nPilZauXnkAWx8JvZUAYIX0OatzA4QXtpecGYVCuh4J4Ryk0LNCLuCp3hjldqr2G
603hQ8ECbrHL94eAl9kKohkhKD7HPuyadIgyWFwAeTkyV3LCNj7mjoO/mrv3Mho+
xoGDCS9MGqfCciRVJ+w6xd/t8xcf9DYqiqC4r04gL3TLA9zW3R2idoLx8rkTMz19
5ZQTrYqESLiI2cewmhKuuPivzQ79+91A1Qt9V6DYLJi2TsnNUWUV2cb6y6GwZyDY
vwaaI0tOvrvjFNNYXUsv4wn1OydWISjY2qwXLZaYYqNODjvEyoZNKpkulYakpJ20
h0hXp0PhpTJLN/wcG9gj6bmfnr5ME4A/GE7WGjKIPN4qgB/63GXTtiqnCEYNaimT
IZyN/Pe5IPAHxwSQJp3db1/VB9/hTOpa9lja76Uh8ZVHHvgbdttWyQeYA2T8G2Uw
Vyv18bJrtDVPz5xnC/quwJ9+la86EYBgrpakwLuo5FXpZMC5q4ElstaO1CR9JkXG
tYaGeaobnMDM9421TqJAJuQp45BEEL1F6CiwDQ2rm1alxZ4lbjBS4vMTJh+S/3rQ
yQI76vK3t55kTLnzqqFrY3Q2YJ78+dstVYOqQx5yiDpYctYKtl3DTdRgjXPv1cDK
cRXMhTKG//+Xk3s1m5ODdSZeVPJ0gL99wACqDKz48C7bInovGWXcHumletcqpqC4
flSrRwSPft3Jsd6w0pR6TScWGmdsrHf8Tg4/xB8I22ZDG6zqVmIhrlxNhb/2apdb
7Az71bHbHon9kGms0enzOzVtot4D/6EY1sQzRdco22bK97b3NUtLK0xDwBlMErgA
TfKBA7QgBJcL4QqjURL3SQDkM4AC9AWTdihFcqSXyeB0D52FRfUiHmF+eUi1FFYs
yzi6yrJBEWlAG95gU8LwbA9NWvRqSb3xiypR0E9POk+CU8jK7FvAema/XBBemtBL
Ft2NdwjeFnu4duRzYowbmDCDQsm7JmW1TwBtOvMkYiVP1qv9KgSY19E8rf81zA4q
WYYz3DpvPSub2d7jLYwHi37f7kqi8hyjl6RBfzDmnrTd4WFtD1J4BCSBTqcJ3Qct
8DN9zbtre3wr+BeMgOl00B6SLEOZBApQPfwwcK8eP7EfVbNTpNdxbl104smth0C4
q5sLOW7GBJzPskYcbr0OE5NOuaXaz/QmWTbcdIKACTfUl74nP4lkv87ObaySr1tW
MEC16pPDELHfTcx/0aW/DsF3hgvwxq6M6GQJ3ZzyyfSxsETfI/Cf2/dGDLQwU3C1
rb8xgfuR/VhoM/hvK92M/zSuomaAPFlRcSUfTJYh0emIwupJ1jX95FSHDy1oGFNt
u/jblLR6PZivxen1b5gsqyTofA114OdfI0m/fMzd15G9DIgQEV7NJlU5KBk9PeP1
WKfM/LuTs3Ka26YIHDknyvWePeZY52RxIMH02PcjsaUGv97UozT4xtn3DyQqGFnJ
Q7QNwA0a08x+EeAFpfFK2dkRx++lsNva0PJHNcaCCCZCFSZP+nGMSUPK47eLHC/+
4nUi9hDq4MsDsbrQglTgXyP5gPPZwHUz0owlQmV8VBV3gZ6E0PwCGHCUkN/MKtpF
RjqzRAj5ZFLQuaNpK/XvgBjKjBG8T+Fv7qlWlhylzpm1PlFo57FRKGj6P0axjGZt
59D2xapv8oErhT92TQZGYU9MpuAinwfqHToekQCAKCK5RNqGUsAtt+sWaenJiQQo
ik0rCepZtzb7WfGqBh7ZWOwDkGKEFeQr4jW52KDGSf8Fb95a7SHkYvHlO8zSmw8A
yOereYnTdI0201y2DGePnZlyF7VKCUETLKicLouniKEBOjH/Z1rxaIY36YtGM/6/
+s9g7rlgmiKlNwH8bOn6Yulwialf7/rWFnCobTp8GbSbDA3CClHlZ2s27jzYDYCH
dqcuM0Rr+l/9wfSe0Pt2wNEcMPPGYMqlTptiN84GfGuMC5Xm9UI+hHPXAmKvti2B
j8QF938moSUr3YFVEaf/SR+YX4kASBrAEFk0CmAb79hByONnVLjsYMicjanTKS1L
OtchWNaPVRaXjrl7ppcxGIkEQAICN34pcBZ28A7ZEaOUyfKcb3FlBtJKRFLym2MG
zR5bOdWZm46c4SVsFyYVhKl5yfx5NTrtlw8PqVzRNJkPUSy1hSzLMh8nhebKg2db
iJ4N3IKL3KKNruHByVXPd0Q9cQjPHActPqCOxlNXAkuMg08C3bD6zsdB1aUOaZSD
wEQXw1aBYO0O5phZgUXv1Ul9OrbHWvYBWFrzSFgcK4RDIAmxwMqSGZbQAGiWFTfm
/b9SBhxnzQXLLDwutuGbGT7sVXxry9Wh72CMAfwOZ0r7VIP47CMyxLl/IszqaEZK
hY9AnR+JExs9AXo3daZ9A51w02BNEgvgLvCKP/GcTQNuHm69qVJW6pWmBJSazJaA
TY4JFNJpUBoQzba/etvGwO3yVtk4k2dFgLc8T035Eyby8kfYMrSCvoQ68EHCb4Kw
dPjqTOVLyFcGZCHJb87Kl1lQHnOADtRWJIW1X+FqdiCiIGgMrM3ySUZdl8LPipPX
HlWq7iI259MTIBVsIP7nd5C0DVQa5wd1b0T3yYs6Jr8VFQj1HYjOU0ONW8kt3Jbf
T079/uhMy/K+bu6rVxn9yYuWp9qNV89xGED8Zb8iBbHRx9/CMKkShdyvRhOfosBy
z73hUdJ2ZFp/osrrfmAwMs/MehIX3SFylyq3xsVpAVG8FSHM7YIPtWO/Tc+o2jWC
RHEaFf9c3I+pAECJdgQP1rVXdXwXQakn3jXK+kcqWt6tE8ELoD2O7ySHaomkTFK1
za27FZJtbJ11umoGXPZ01wAPDbybHbZ8j9wMIZNlKtkOG95G0TcpqU03XOeepy+L
46W9i3AZZbZ3/FThe+Lh2OfH88o5oWYs3qW4Z4Iu/6d2ryQOwkrL1gzZdbcJjtLe
lOTRhFTjigyrT6VFo4YsBcJ3WmxdoWsfZwwO1p4TSc537zlZ2TTNcc86t06GlWCZ
DLb3s2xlC+69xqYQStq5v7jF7LR7OQloFdOKCvMfSBI1doM6rR94kQ3QbP0roMFR
MTc0tH9X9MxHjkXnxjBhQWnkaUbsg9xxTndXj1gKl7uW6dTxeSg23fFSwa3Cs2Sc
WJk7OB8QOenONlntJIVam62G/0Uuy7JvdsGEC3C+7kkX0XnRbXkKZsOV0vqy9cAs
jYlFctbODmy+0spQ9gz5gsSkpJivjo/nTwNEv3JOUzLmMSsmBuPetvh5VUzYQEpU
tC8rXyajvtKj8Oklq05NtbY0kO0F6k2YJzcbJ/lc7beVKC/1zgpuiMCgsSAtik6F
v8N0k0H4abABOYKcaBpbH7N5x2SmEfcc+wnhA8G6Li0V4nWH0Uf5yxmeq9NHzLon
cyQnNkGF+xEL3LDGKp5LHoYl5uGL891G9y0zyy5g1SMJkqy1cu13cRlVgS5Q1wLQ
UjFvS37PX+CPdsyPec7+l1clrcMJEGD9aCXWBJ3n38dQdDlzgYV+vfRi2MHgtOoZ
9OS6Tdo4FjRGObRG7+Ay2caksmkxxhLJc2WkD1SlfVtqVHWTZ1tLIp/RqK4DtPH9
gDpJ/JkCd6CcPGiFrvt2YTP9AZWwGR7USVyh4BxLy4rXCNHa+6Ci5oMbp/lpFLQ+
7LyfYmH9ahyD/OAPC/daFeW5HLF4TpTJ4aBCuiAYySAez8pio30ZVZ0jFTaQhTRI
rBYw4b5UOXGwDti8h6Ymbpt/62FCRtMLY3vzZ7OSzC8lWqTAiFL7gaYJXCLVGjfc
XvBcUQm+sMPTM/ZPlKPpIjYHhVvmht4pkmkvDWie8aHwO7Dft0Ue942qPQJ287Yu
PFzAoJmWBrMF/nDhQyydx3Ix2iOQRmYDhz9DuGhoG44jQt+AvYQuxRegGk6uHfOV
wyiOwsNO907jirjUdNugv0VU14Xw3ksOReDTh4GSrijcaxIOhU1hoH4WWlbD4bU8
6SYh4GlUFK4XSdnjEaj1jxNQQfgnKchz5Mh2aTQvitVQxc7JvJ0QH9hUYVK2Qka9
+Q5iR9JaQF5a7b2Osv4QEoggaSF3wRK87eJiv2blCrkNJA1p0pk+fuJeThb2dRKe
WbVw6nOzzf9Y8zSmLS19XzM5khng9EgfYf2QTUXvDFsQEgsdAEmSyimITwS/LhIU
DWNduCj+0ElBQZhQ/yLtu2erxB0t2Ny81b9AGlhGEN4dlqw56K3/EgOlW9Dc785B
XvjgUVNmyEUVleeqcNJ7eqpCklfTh0A3RDhVqgfPobIL4z4dNGptpCM7cXGUc9Gq
mEdOjEpnk4s70UwDQ1Wt8TwL3hKxrpFTVLRg3rbGBQu5Esw328P6+umaPGt2h7/H
HdIUPqTWKHeCASDjZUgRF8zpyp0/OLmiEFIWKgKrT8XABGGYPGHaZ8BI1Nt9QyxL
lVoot2YGwsYXEH0t5EqbQOVPaC1wRbCM3qvHGOa8S+NbIonL5djkF0z1ytP5tD7a
wa7Tvge2DcVBtAmADi7vBWDySPVfbqx1OGTZg3AxhFDrei/BA0uVw89tPJG4ybx0
+fbm2UestEUOek7psayiHwdckDxE1GQBIJH+otRiFoO3L+Qvkj6x+sGTlgadPayD
EUm6EZQ3nxqnYRwWBggTDsUZHZCQVLkWiGLvM7x4Kwfjqvh6ZJARbpIGRtyiJaOQ
XgT54b3J6DASVwYUwIu2i8jDdkxUai5rBKzYK/A0oOoCQksgvGcE/3cO0eekdG/a
vm2zh4YrYpjazXXNlYcKAI2R0l4v8EYyYnBB61chmIZNAmlQuv55JfflH+xKT+4L
g2zirTx/v1+fyi++fCY3TkjyuUQqva9ypKtKwmehGurEzeSSanKU2Z9JieTKFq1A
W8QmPdZ3PUcQg5WPBcbYQpSZMWLJ4j4r1BstwGBjFPWJul5NTV2r9PSSW0U+WSrs
Qtok7yQdw8huj4uZYjDFgDWy/oW0bf4gg2WYRGuCaess/6hK4ZtnoUr8xvJgRHgh
x7LfZZVpKF6kGRxU45fQNK0oUFkGZLZkJCsiCFOsKhrliEiCr3zJ4e4e5AK57zj/
PLv6/TCIsDud0LhrlFOFSzcA023+5SMeoJYBX8h6oQiG87aY55IghjvUKOC+05BS
Cn6gcNiBxwnYCqKj0rDgnQ6f1p0uH6x9z5VdLzHP8xW1FopZHaURmKUIX+qoaoYc
PraXPIiydPkZB28d59ypP/40El4DGuPQSv4BsEhtircJAktf10qBS7WYyF4npb48
3FcIWoA662u/XjsjXv5OYMUYzl1Xe2OJ6uGtJ/mKWvBoEKNyDOHIrDzy6hfcNxTI
9KObWF1aWaIavo9rdsjbNArVx3fVr+tELMgnBZMd/YW55MiXsbRkoRYho1UjQnxX
itvqKbDcD5w3WGu5+RlnlDbn+oKCK63wzi8RxgLaQ3+6ysEpmmXayAASUGIYA8MF
DAQutXp+N/9h5itxMQn2gyo4sQicf06ZYJqTUP3brARGrlu9LFujPCM6UxgGzzLJ
OJdB4e0wustKjmzZZuumBf67Xd0HFQZ/wgv4m00450NZWdw5kdT1h7IDVG7GG1db
HydSf6Js06UZaU5R9AAF8fQtYeekPQ72R9rhJWMJAZaFcu3d4WF4oXCCpZuc4v91
/+m4UjmyoO3SVLvyI7VKm4sUKDXq8p2r+1EGtX61xNM2ZERWBOKBwpS2pAbdsE67
ka0qKlBLTvdo13Hu5d0MXuujnUPSUhJxLh8QQzs86z9c9z0On3DNMWLaqBvWhoLO
HofVAnFZOzmQlqfFVn/0GGioB8F2kiYr7okz2uNYDRsqLwVDeB+vx7nqWXvTZyK4
PlO+rDdD8pnESBb+b4W1LTTBLTeRouJYjOZYKRVdBHqYWArAF1veT0tMlnsodH2T
9+3BWwIgbkshQag+GRH4CkWd3gaCAkXRqOiZhenmbLTbb0Vrn49lpwx+oO5DYAn5
zDZ/kpGQbX4Kd/C2uOJ6JQVmy7NwbTi3wAKIXWAOLifMcp39lNT0M5VdCUQoXLgn
RBu12+FN/vFmVkp88hiLKiUQeYvvU+OzxxFgwq7LCGQjuzpkCbJnWRG3gBN7wyiD
1gwhVtwLexR7n4GI1Pxk99hC57yLrKYZI+MkWw9C8KuAhh79xeOplUzgGrCZjj5U
IvFuSqB32GeaarVB0DSyrr7plKhqEVU1NEixUyMkaIcZ6PVKy7IWEXD+ghfcXWB0
UZEbc0bMZHSNZjpR44jGSAMJTYVUfKNfakS15BZinskK0X4YwsvVyBIK15xy7pww
HgNgTn9kI7XNGoa445jjy8sCiOdz87TTv7t7BgMEf5nwbUTcfFoRXmdQrXZ7ToKT
anOXMb9lB5xSVg1wnxiER9IIWzXEeHHY+mHti5V4bLk+rtO7w5rAtbwxFMxvg+jh
A9NRmgagBwRynk6VGBiyIOInSGX+UumGAcP8zhnUNh5cJ3VskXB0WARqe5JIvXNG
p1DyIkfa/WaCyNDYeNe1Fqk4y/SGHS8Ew8zRAU+8a+vRHdMR0T5mnaaxCZpzDo2R
ft23TkOgdAUIabQdJo3WVcMR+A8Lx88pKAYnU8bJjqA6nPSORmeWZFjZ0o5gNCQj
dqKTaJ5BYeHNIuTgmN8qLVK7zLiff34y9V/DUeKLAyA5Wt7NiRWing2ov4w6v73c
lOezZ+E+j85dhmq7ebffVB2uKC3WmlEp1KL8vp0myfjkpAX5Kk9APgt7oqSZ2l15
6QkTkhXx6i2kppfGBSu0w9YXGBFHRqzmMQG3qSTg1MhvrxxoQGFmCzbWKDmch5f0
4nqgrfAQVpmuX83GZTc8PmGiCdcxCM4OZqhGAAxaou4EXA7ZQNjKQGHjEaU1ePoO
Prz49Yn9Vb497u9JJy/JR5omxZOTmWg8lMwmc/wlnqmdUIYxnguZmqpncjJaAq7O
v6MMdgfQpAS1EHpdmwPytFDIj30Og+feXtyzZPRE2rx2I6s3+PqPjm+a7MWTEc40
W4Yy2w8QvTGTbgRX+ija331k+gft86OcyDTd7MsFy00IWjeA749rk2NKzvhKravr
MB004bU3REIyBLrd+nw7zLuxsKMxpWLdtat4L+5zFTUfBH/Vhsyuggo9+UnnjGy0
8Z2iHaztNsNGonXJQx8Hdh0QOHnhZpHh6lacrqiGmA4gUZ4g4yPV4FX7u5yvdCer
pldEJYmYYG1QzwqJlc4xZMmYMqVmFbUthiJnTFjOOyx8549ojZzslSv0Vr6xf/gD
bGK1pdG9zx/CCGHyj2fzzL39ayjKQ2Azx6eEiu0m470IzYwrixzQoPumP2hMmNG0
ZYP1mci3ZX21uieJgRflA8CrqVRIbn1tDl5Ac3UnrrWX5LKmFOXxWbOvqzrpfUEt
Vh04m+/+0mg0TPoiWe61hmEyVXuVYNSyT5zF8gF5x0JhflA2DlfQp4DTUddqBL18
ezFjq9xirIr/WgIFf/lu0ZC/ukA9A9oZ2amepNc9ej8vpg+7lsDLzCfvS+tXeUFq
UF19LtdbK3j+9H+Y8sqa7k21OD8HalxjhLtx44z2Ebu8SIKRrUXJJETvmt0qJ9po
q65xDwEbRsazmQ55/T+v17qTIz1AkN5Av8M1t/B+pq7FjJK1wGKScxPmI2RvRnm6
E78WTD5gXie9p/5PK+1xkUBPakUvPM2+bOU2FWby168TG6jw2kC7zJOB+3GxlE/b
ccNrust5yFuMcCo4R1wzP1mqPqALcpi4/yNpNdzDMwQhvsOvo1w6pn0k0RRKtvQ/
79FczFxcDB6vAZCujyYA5I0sgZIvo+Q/UDh0F/TSdyGzgMzhF9uFvE6zos1TjiFN
GVj+uUBXaeR9xDZG8k51P7W5lA+Qj+y9F6C7t7YdDGCVc4CYygo1Kmt7CXg0s+Sm
Z5nLLYKxSPw+4883mthz+NvMaJyMDrgvBSWkGR/kDSI4UzcWO6fX2j9KiGE4gc1b
N37dkZisl4AbQfy7xo596mnU9i1tbdP70BWbjPSIgl9935IY9Wc8RIvbn8IIeM3P
0iXVI3pYgjOXDnflGivOeUjK4g9kWAVzGL9PTJnPZ6qL22GmOQxkIOWPY+OXLsaI
Y/Hbpp6TJ+HKg4Lr3urTJvmBiZOq8mYxgvCDcTbv8jQD01jxmVCLQUg+EB6XWl0o
nhkN2ObIG/NvCZg4M5VOugTrpPdsP7o22+HmO5kWjFzWOApwFoVvkchgSoaeMDm+
iIAwPc4eGF7BlhrmahCpKczyokQ4mU7UfzBE7R1sN0DrQCNYX/6FqT9LlntVgVGI
p+L+Fo10qM8Byb1YMBUiKcKvkQPwpZxuBVNUXZFDqN6D4WLf343k0+PrXE/Tj62j
eRILeF6Ieewwb+LYnBg36E1W9QPThzZDyNwPebc/vXHMceQBOAT5OlI8saa5TnVI
JUe7hFXB0HrJnfkTXb5c19lvKoJEK2EQDLhtzeeEAT6jJojRvRnc8EVklMQRvBsh
l4zlsftzpkAbilpDxgEVaGKxhxaIwI2uSgJED6gVgFxW6sQC4wdTEh+2DvdbPhNg
/rlbMPsLaN3e6zuJynjhRdL2RnS+Mq4iDTRrAv0YEOqYt9vo5MQAHZvaHs7M/L3Y
uFnYFt8vGs1s9ZwJeJPjI5oVPtt2pMnZx+FZPLz+jdbiuzNrdfJB8qIC9XPeVck4
RFDS5BLLqylWBGTVBsXMdI9UXIOvR0KSF4XNvi14vwwBp1DNw85Odie7/D3XPXoi
sAW56Y8IKeymlp3Vw+jRmZIKrP6Dtk9gDJBTBe4JJrbdxgHajBmFyWovfb2IST5b
wmtkoDFSDhJ+tyT9IMOaX+R/phTz6vAKyjmkkiELicbBa8iA1m6QXe2vl0cfJDo1
lecBpZ0kDVnV7DaZmFnU8hZVpiMj6+8pcDfU+6hgaV2gNus/q+/RqR1Y742JlFsK
0hjI3vDHav0ZDsIUw/wglVh1N45gUkVDE7s4SZGR82dMzJTsZceBPS9zgmXfdQFs
uRayIMG4sEzMqC/HCVReabt/lWfGo4+sYG8AvP+1d2r5fr1rsfVy7ikCPT1ziqJ3
7y3fmyntPV4BeRo22e2MrH4huNwLhaXFHIvQsDoZWbuWbbxoMC2q1MU2HGdWmimx
Yh9NkZnFWNRXwl2h7E2+ZeiiKe+C3ReFFwPO27lp2Akncd7nh9Xfj6QWDM+CszSV
PtR8fUGNq0dep5RzQ80yuayx7XoC/0TANh7s/ff5/mcCviK4Vi4SZoOc1jKZDlnM
4HSdBPdSCvQqzRw0R/Zf24IGKwSv20uFK9zxniWmVWfu1TOzlAr6a7uVTBj/w9dQ
4yEWtWITuG00d6d6PXzo0pfPEHb2ORDxNB3XYBfwAbpIe3/o4roF0RUby4WFCx8u
cH+Ext3wW+UXncJz4pIRF5Zr0xevmVInnDmkNPxykVWvXiuKv6G1IVEPfiGfWxb5
bANVL19tWgGAWTUArizECIXQK3qYim1IqMRTvmJIQ5L6ypJ5+HYdY/Uhg64mJ99/
EdVLN8veL2Kobir89b8zjacWwNbVT94+OQ2Xi5jWh9H363fX93BMAJV/t1pA6D2v
4vqQxKsr4LsH8AwxtRzmHERe0PrtXGjZKnOqvV+kKHB3fVCDTfZooRyastVep3OC
yKzNl5FhoEdkFv4bieP5svOrg/bmEz9K/EMe1FC+gLerijIAEr3vObe6bk5DNVE9
vu50V9wjjoDKis1Gu0XRSVPe8mqcXPS1keucwR6RDB64qV70tSy6D4NomyHcC/VD
vM4c79kEcs959bUjNhPIUopkfffcrGEpnrb6Jdaw8dXUT3/xi/ykCY3LqvbLCw4Q
51B4Q4CW1Vq8A+oOOtVawoCDRN/BG6TAvc2HlpCcvH0NeZ2NMNixHUceM3pALLom
Tnqgq+XTulhgWZU/iCxTBUPH+ON1wTVqaW81pw4KAC7t51MiVNVqvKzi/xgFvfaJ
1jinSiMnWqYlHkqaZ+6xq+qCwpYQ2sqkkHRT5yfcHDrthfAaxpB5UHDaUsQf616h
1apWBn8NVcjs37peTyVTok57b10U1cSqOTJacVGj3euu8T5c+rWrMG1/W+0SbXgI
adfxznc/pvBhZF7BFkODe24g2WVo6F1fH3j/F6FDOiI7GxopsHyrVv+ker+hkWtM
o7YBibBbAIbv4zAykKoKocg3It9Rhc8iBA1PutnexkaxsMlaB4eoyO6+kLK8pOLB
ktfxSSDjBdvS/yLwWUhMg2AKNLuTwS9Wd2FFtIZdx37cFuhdAxypW5dJOZGyzHZX
t7UsSzo9Nn42348KMoilmk78GadGWQpo190wXZSz38ufoyCWRZaFcioNXCcGeMhT
ZrcFSYK/SjgQ5fB2fYGqPGrLzaPIXgn1VXSIvH/WK4Vy4lnocvV2hxFTGhgTKY6P
qWiFQdS4/QJn8QgueLTwA59gOEu1NbeIvr2Oatj92bRnah5mGybWwpPQPKjusa2M
C7CV1vYZwS8To75KXNxGLUOgUeS/0mY0gST7IL3Z5AfHLb7dalyxbVzrWTEBh0RZ
ZL/YtDajaQgUeOtYpcYiKomNko32HLNA+/VN0m9m63rJzOAgJEka5d0w1UztLZU3
akI9ApWpgGShUSYDypwbla2QFIPPlGqhOIQmWiJ3+6un5IjjyK70biMYho6Bju8U
pbwfL1smZMN9aHx50FVbcXnm89TM0BlgmfftgRdVbYE2+09/ZgeZ1NWO8hkDs/bT
eBapl8VzvSIcku1b+/HwSm5CIC4xRBiUth7thgd3zpc5Kagq3PMfjmfDlKyHeD8q
YyUqJz2HAjIcf0CP1NOQyCTQJCUv2TOjAwn15OK/r0Qk+7xYUikUXyS16G90YdLy
JrNxiKBR+2+fV/bAWjKQ8iQFWrVb287Kx1p5vYdv2Vj9AOrMmlssMUhgKJoVFijd
AxRfGAEUMPcoGNPxLOK8tKHyX0Jqmtr3NuexGKQrMYEJEYwIlig69tFLW+B2HBHf
9BspKvBH0Wzc7f0o5lErSiqPpxvjFLpYbY2l9VEY79weanxD1H6ioNSa4U2cmxaZ
rN9E6L2xvHYUU4M0z0iVhlT3dtz4g9AhzlN2x8uJh6d0tn5Rh4nrNCcOyDiX1Dkr
vlFxFEFr3Rb/CwWkCv75kW+90V41IMYo2ppDxSmlMwwTUPqHF/W4LSOL3osacJqz
S3Pv+fXaGljwQLfCNwJHDMJ37PYfzq0+5Z4HPQC/OZehBKjYBpI2a7eLx82JhMHJ
0FvYQc3+EXn2/rxHENm8QakvEpLD4KZ+BaEtltu1+OmzZ1WvLaj4+ZlfCR3X2ICX
tHgWA76U/nHicBYb4BSzBzzKMODCH/PRc0w0BR3F2Yw1hCNDFTEWFD/ma6tUeYev
IuyTC6dU8VgltE8WXgP2vHUBtKZmR7j2oTz70wJbGMFpfqH26RqFYcg9y1a1X/ca
rWVAbJPHR7iBDEeXEnYDvLZgLgxD8yJoLaCqYzJDurqtGEyMSIRhIWiGHCmPzJYC
5Tm/PYrUf8uMNnF0GXOySkcLcqVC74EWWKZVwyeD/wAGabyDktt0bUUGNu4ZWxel
62KRQeD1LvPVPWdsj99Z2Tm1lJpFlLQxTo73/HoKpvba7gie6LfPkcC0HwIhgNvp
d0PlmeGRqVO/akfvyslneD0WfcAjR30fVXFRQfg/L9rQAE8qAIhus/w7Tw/sjrSo
h7kC2dkeEnz/lkK3ZDtbjR4b2Wpy1FVWtiyreYWtZppF8znt9ODjN3SKipKTI904
cNdLifaFPCFldr30tsqdRdXfT4/AwYuel/Sh+JKkBuOxbH3rrRGQ1SPqzXiUA0BC
o515dwm21dpUdm/er88tfJpThBcukIdNDGSofChsn/VxdGyadXKG134TPjYmD+ZU
Isicm+Es9zKM39tcTAIpin0FKHpgN+3EEk/86LWDorHkOB6Llz5hiwGuoCHFweW7
nHTqNZXmZB8z7ywRKl5ybU4DG0jdW1O6VmdyLOt+wJE4wRwYPn7onLPo6+BcB0Dy
Tu6o0NGN4t8w8XVFIItIaiaKpw1XGcoF+trhsxFkp+eX94CTMHDstR7LK/b0hFxO
PoZ9owZssb2idBUdyUkepVHarOschWFY7eoiT4CK8LKfiDsX/C0HjQymxh9a1U3p
fU1q5EisOfSsYoSaHJy7H+e6W5V+FCGXdM6usmSQat8IDRC2+Mi8eOVmdL2LUs2B
cfTtgKgLha4O4KmTx/o0Q/feSHuw/bEjA39SZMc3UNm1fXrI8pn7YVGS/A5MDs7n
FM2hpnKHyny2WF8/8P+fTW2fcNRWtO3T9HPPGUKp978NGHnMPmwRnQek74a9dz4G
mVOugO19gFLBhKlM+hDYLn7Z/GCcRssKtEUFGvGZUioyEF8D2MfwufFVW6HgZwZz
UBGL/ZotPxltVW0ozh63sBAJGYvWqmQwYZtk+yAB4CsWJ92msJpSqH7KU3S80cnq
rdN7Nma89aWRQXzUDrn7bWhaVUzxhyk8vs+4vF/hvdrFd1JB804MuVCH3R96BSAq
NVqRwWw4Ne0RAnBuRUvpohu7xkpPSdVUwuTbhwEGhVpr4AqhN6LytIhW4V1PAkQo
fGCH87Ul4BZv4wDebBRKDNh8hMPcmb9wmrU/Uw1PdGbiln5z2I3Uh6IocMpcBJJn
FQ/rbP7hnSbOzk+ioct3VfKREN8xLS3n98whDYvMTP6dCf+bP6xz7vBAcbvgfns1
v2MJUYAd9tHGjnLACtiqcDa/VE2Bft5+/MZb4IJ4frjOTBlAYRWujjuU/Y7r6ulF
6tR1Gt3aNV8ybI4l+U03LNCfBDeKVxPL6cZRQPFZqPS8sJqZ825onsRmzmBdbehK
b8JG0t4C98phcJO3big3LZFjcE9/ZY8aguOa7NOfETlo4qdaGzSIT4gWNQuuGuq6
7VuhCrEcML+LzCkeS3Lj8AZNM5jbjuD1nsQ/XfLfSQg72Beeks5Bvz/H+Q6DXZJe
//190xmPiMe2TN7nghX0sIDzqMptVBpmfkvNxuAALWgY2G0kOi6Q0DObhNz0mAtg
DqeCOVD+H2sJhU1sr3nNnhcEd9OH8zy7byYz82OqcQ6hpFwC0NIvBo0ONp1WiKDr
V5/IzE/LPEV/r1F3UrAOa1BFls+LaMOwEm/1migkq17d5c3UAqY4+mCvoMGkZ4/S
aAlKqeogj4PeTSxUkH+ydAUxAgUW7ATvVftnsCTKk0uBcEeeh6JJW4McjZLQaQKL
9RvKI9Ax0rkkdYKP9nYEw3EaMXx5ReZr+BBxnkZ0F4fA0H4bxnTYJsqcXNcQRJr9
ep1+TNFH37coy58rhxMwUTNvZ9i03eCAo608rDdZkI4gRlCChpZEUETDwTjcXctX
78FOZLeb6k902ykK9zoCI+40AOzrM5wwFKcN6XyikeRZDakXAcn1+H/6GoEd0dEm
+d0LqwH0npl6QDTBSH6R1mDluaqFvcUXkMiwA0EkqmpYIUIeU1tPutPZqdv7OKOX
UCHDQWlECW0qM42TeoKaSK2r1s5MpKaEok5G82eTx0y7yYPoBKoQcuUkMPuCpd3w
BkL21WvAvima39NRyORoWOpHy/jMk8SYTR/ADJrSchPvl3e34wkip6oyYUjvlgSx
mWENN4X0mecv9hMxFFjUbYZFzTZ79FLLsksopsgYmbokDQ3p0b2vo8C5piDEzLHK
l++KhwDNqKXGkX7Wi9ZB00uX1xRhwqp5MgptF/xadon7KPzaOdkmwPOeQ4u3OLCn
oZCIjxx2L/+V2Ki5hu0sd5seAGVfmSu8i2KzzihzwsupVWFChwaAojSy11+QwWVO
fci0uSei1liuwL6bNCwu23P0VSF/Bk6pzD25eyT1xfth5EyGVQ/a2BdkIzG9vhEa
42MAh7kqFN6Yh6F3Yt/KUoFANQMtCwO0isISp2SXKhYoXZ9eTw9nntTlIOu2qn0J
KLVxlzhrd6YtKktY4xJQ4uKGQYaUG41tjT2LrTLe8g6fNo/FGIOZz3bkwmQ9mo3s
RWOqkLWgtvA4KA5SI1eL4bKKFfsauFUwj548YjH0LrkRX6nUWb60+H1LG+8gXznk
Zs5NMsv+oVynorJr5UNP9T3GvkqEu78ZCso4c7fA+DakAvETGB3EF8Jqr3JhVKDS
AIgXjlqC1inXAw0lQm8H1qXQ9iSg6tEfYA6Tvz0HeRBB6wxTJoojRYj+HTUAxLhB
0AoonA2aAoxaqVX1B2WV4xCcwMSLjgIq3Y51D23I4oqOAmIC0rvRsgGHZlWG6x2y
i9goES44YfhvUy1b4cUNFRIDpzcmsrV6tHhvEamQYCiVAIJrmL053woyDtTZF382
Bcr3W4jRVnL+vHMv2eBvllqV5Imz6oWv0ER10B34Wu2m1laMMVVi0Gx801X7K0Wm
TI/YqK7c58WacrumyWMVYsYEJ1VcyPXMvaQ7YHzVEZ73nlx82CBgcPpRf2Mtql/Q
mwpZu9swLCgcg4/arDJ0a0C7j40kwpU2SoM2unn2S3DhfYWxJ0DdiYYJMzeoa2dW
k2xmNEbYOSt5Fh+m5ev7UFZSTpOOlspRZBr7cxHNgpCydOLwNUVDxFzn5tH+yXPZ
OCbo8+xgRrCpB5DfT7jfQI8ApTrVmihb7HCz14OsMhfZpWQt0cxZxw5pB79EfPZn
My26uRHNVrDXDitWYbI0dZgFexLJb9o2f/30S328jyNrHBkiTbm+LO0Y16CGJFd6
GzPZNCiG+pgnBfvz0KVK3Tra2QUmANHcqo+kfrR4Ei1ag73K1j46tJeTXsrGFpaO
/YHkK3A2cgv0QZ/ZMdwl/Z9ZnpT1X0OYOYuG4/tpDu2QxZ+ElYCyFvochgFenOuo
gpjqyslboM0u8Q30NMLv2RXz8OAGNiTDitp1tdWuPKQ8AtcVNJhfinjUEMe0JKKg
cfOJ9IDYgLAvf0QCTKhfC/fxKqgOUUJjN9bejZN3rMAAK4DV/U8GM7TwDM7ZSkHe
m4MMIbEAaM9Ee6TIzqibl62rVRzUssbCoitG815ericv5pR4jxWOLpYUaLBOwh40
SJH5tmJFuxuGmtrhsmUzo+PHNfeZF3duDwUTInWoKhv9Cv1trCsswWQxiThyZ+Q/
XXHubT25oc0aR9AIfqNFo+POzkTzNs96ZRD1diX6M5AvkKXj1jkyxLtMKWYr/pvO
SAb0S8onGtkJN5tgZhCLT2fK5twZzSltBHzS84mM1pyiO9EPyqoBCZrjM4FXCbEN
hcNhiupROJk9rahkHU2qlFTetilncHz9XX9eyLRtMy4qewYMt5jazItGNe4q6Fc3
t5zjggLS8K+ZZkWfZzsguu++xtYPzFJPeGx+8VGZ0dhaV4VrTyx1mXe4WEgaDy7y
hVTXWAoNwirb2ICOn0ux9+IqfDTq1CdDhR/X//9bU7DixyKrwATHeRF2HKhlEo0e
qkadYnEWq/Q7lvqVZx8zoQeyoIpZoiWzWx/9IJAfdRq+8AWyL/BDlnenNKJMPjQI
vHFRjpTIdRzIajY3oS2uLQVwwBGKBoYtltqsMahwS52Iogzp/5nqooObYfPfT+yV
J4d3UBlJCi7zEkmhyorCEMBqqdCs33jrC9vYNbpzuvUJ9ijuXwxvcZVVhT4bcGO3
CNWlXRl/0+SU2cSQoMybqY+lCJkeykCsVp8kFgWJsYkYkFmqlQ7LsxZ0/d++mVvu
RVb0GvMC4w3dl/C/j4EMA+p5df0DPznHW5Atd3dphDy7U04HXHC12Pd55a7JIsAr
/LNhNw1VFRo5XgX77hlB5fIwuPJTVDrluZivmGvm+eCVIXHQEf8JlYurOqrVnjue
XypP1bt0C6p4+kqiNb7K4JltFS0gZncUzFba+RieYxhbXYBG65+PEzrUuyriqT/g
xDCrHw7cYa7HpnSk0xCoCChYzaDrpDB6sOJwUADTtz8IzpxnjD7ho5tfd2TCk8tZ
eaZ1DDn23X8eDNvtV9ds4DvS2JGuNnJmoFCx9+m4waSGhhoACfoIAffA4Y4CNNnX
2ZfhNxfchz3qC7qFdsq2gcPVQC03tJjFkB+i/XrP5aZ+0PzJRGYiOG/sRShQiIqC
JslH/e0Q9HW/UccMZr4cl2aCtKiOAo8s2Mw8/5cZh5gTcGx1zt7SGua7hHH13d3g
M+rkCqjy3NGcsfa+Y81kaxy3CTVm/OvOjmmyQYFMo+M6PT5tTepl394IydX1qc9l
Yi9xj5+iZULluYpozWuP7hSt/cE4kqllHQPfLg+pcFbMMGHaqVdZiRMVpNi0Bhs8
T/swfBHnCjP1yw8hFvz2I21iYSvQ8796DHaIdwYC+PGk0i7bc2XtsjZcgyWg1Wu9
0k9y0/6dUCru5u4JucvNd0gH+eCjr04mkfsX7b+487HSq5d03UWASSg5q9xMDJM/
PAqTj0JHd9nnwbEMgysVb6qhqZcrCPRLxHhG4qwiX/y+lUq3IOaQ1MrdnLXC8Huf
d7wlw4w0T43xKnyW7tHGoe0IygDOuON1+P8FUPX7rl52ZfFeKZoXWolPlgylxxd4
BJVxCJ3yF+tmkgHnGWllVrUNB4GFu1XGi4Nf4XRO7l7YIDyZjYThTN7RsqFUNWYG
uIgvIu0r3qZyeF0+W2BskOD1vcBQW4tWTI56egPb/BSy0jfPglUZDA3KeLgaPzGZ
+ZUINDIlXPTxqhxkf9fAUQhEmbfp7Y6b2orYDQ0LKpfnSUtBe/qz/7mbk1mXqlIv
wKPG1R35QIub7pHYprUHRAS4BYoSmJgXj7hpcP/Y2lkrpv+d976n33GrxyrkQheE
0RzyCe0/8ya7t0u5ZAm19yg60AefX2IyD/sIa2q7mU+42q7WLKCJ/sSdOWPyhe51
JZoQmnad8etnSOdSxKWTqBc7LXJDnGUNhsaM51po7oBYaZKYJibMsOx8fPsviIU4
ZaDr81TBF9vPhoNZEwsLra/vGVXAeytCmzVg1dlBjz16uj8OhkuYHTfUQwOiByoy
FY8PWiKkMtWJXI2xsu82OW5TcYMsk6yPk6YdsXrCX9/y+Do2s0d2FzWgq+NZ/z/e
Bgynr59LAyVEgYrf0SqDtqFKEmagp76HwGYO75m5L/06AT6+qi9tKEQEB3h3fkol
MTsLW6N8ROmJuWSp7vn08WzuEG7lBkY0g2DdRrvTQOeqXHdrWpcOFH2Reair1KGa
/VZbS5xadeWz+LeisbBMi8en6+FwnCAf+RPuTSEUM5Nu8XISLHbWK6Yd1dWLjmDG
p4k9k6SlGSxyETan42HGSrCt2+cXLrY5avjJlHBqlUxHd76N1J5C1dSAb1bO6Ro5
FQJBOs0vw+Z6Izpy15Orq858rPKrLu77/M3Zt17GtXtJvjluzQ0My6n7erwCxOKR
NWgSmVNNyao2SoPJc0zcy7OfauWXocwzG5FpnkHidFWCBBXQw6GmuZJJkae+bxiq
ijLk4LP7YhqpAH7jsX1Fi9jnAyhsjIfU5Le2B1P8MhtwGdX8PoS94fKhgarH4abb
F0y6F+oIrVQevVb7ejy/IXLd+9NDqFoR3ZAcEnaZuAZcanDzgaOpxyxTIFFEmkDQ
crHdkWnjzw9uYjvxZm/N9TPov7hGKapEdfBdtuyUrSrzV9xiev33clonYzAI4P8J
ZKC7WgmHjXbpvvct2ZlUo9OzRqXkXuwCYMvbPr897KNS000GFl25VinRf961dk4W
dmhNMAd7a+tT9zm8s3BjFnJRgz8Ic2lIJtGIEIQIx4BIcHA5kQK2caTSy6QA6QEz
7+bkmuVImneYp9hcqrUmoyCm0oac35kU4U6mMyMZ2cH+GSehcBk+xvoZ/EWky8oj
HXDZHYmseWhc7r41i343gA9zjJPsDazpjz1HNVuPfIfVcKNDNzBfA1f1cZUAgs9f
tAFLZDnBTVXwocScl7YbVgwmlhQl7NfH/8eNp9eAvvkBYHHhYuQlUCXyqYRrNIZ0
fAW3V0vj//nEUItj76YJDT1A4a8w9U2NqVLfjnksdST/UphO3t/US0wYHWh/eN9A
6b/OyJ9m9lf6pNvRHqKmLUY47fcvm9BHfQG+tYBf7y8KgzHxoUPPbk3a+XT+ObXR
pqNRS4GVF7GlkmE7zT3eJBv9JJ+3kAX4epLp8vq76BU6WCi6ph7csyX14eL45WMn
hVN5GNbs3FpzS0n+L21t4zgef4b+80gelYUUK0S8pA8TQR5CZC/M+zByX/6sDahX
4InL2l7NDtvJjLRDtPCqeFWxKz6yHLUGj5G0NcCTahKawgWySEVLe02pGM9oh+h5
6OocH+hxFbheZqhW4uzK/Ot7rNLH/ITr3FFkDtJqKAkuG7Y/WQyD5L2ngl7O3ANX
vuvL3fsjkLNUb+Lo1LsWQqACXdRUWFsNM+MTKkjZ5HsXar81BaseCkHBMC86EPBO
S92Z6id3t/zoMaGR/WFmIYd0udGMEB2aXlqe3Da4DP6wjq17I4qLpGyXV83kvKgP
f9NIANYM4pUtdwthMQz5dkYXp4K1b2sP/0O/MVI4CD2jp1tcjml/rPH7y7wKRjx4
YB3SSmRufKVFUMDOD+wuaAuQ0YUybW+V1C2RVT0U3zHtqav91KWXPTT064IQd6cY
WRXql/h+bG6ecT50e7K8WQ2yh3ZMR7nYiF5HzALbDqU1aRxLzotMDeUnvvlQLXIz
W+QFzbnuEclLdFOA6wa1NKNgNtx8BhJn8dUzUikd25YTLsbA4vSxd4GJL+7Zdk+O
DFXOzjLChuqHDKmHHFx9qtqAKiwWU8UllKxBtQ9EvHtIUJZ4rrxJNL0u/XFSdzd+
TPyRAk/YOwCHt/sTOeaszKJQ586c/25kvdquRNiPTXovUopOl/CdxDsIqfK5RB20
8c4EQyfF2FYzAxWZH1c4wyg8UPHTkKcb3XAuNKvESwdd8DU2oFzlMbJ2KBqCGEn/
T77dCeGffcPVsSUKCR6T+R086U++Ys8tPhoUjKqoaBhsCF2tRpLaavYXfJXKHMNs
gm3YYiLolwqFJcTuC3d4u4vQmENulljrbUmSJElPhkXJaerIp6H0o5PIyFJqndDE
wr2S7fThg9NicUmy3YgqZ5cxzRa04D3J5NWw/j8KeswhGMJkTeH5lbK0dvTp7z+D
ryNhnjUyxycuDKiJuPec+4IhcVyJZD6yFCakUdgUBs11++QlOcP5j78yfDH/GiG+
MBzbTHeeY0x7IFaL80irI/9GkShbo4H5HVXqG7YwZbhPfY0vAPVWyhzEHZWwKocS
h93M7/qaRnMFG580J8v1LCPhEfsqxDfLz/z5nL5OmWAsf1ByWo8NUm8IXmAr4fP2
1EyuE2cuaPz3MP4z6/n2zHfCgjcm9U0B+r6RJgOjD3HdkEP6h5UasnpaljWN6j9U
wTOVD0AZHWz2kHCouczMFueTzPq7F9VDZlAsZicqRpHvjSqRsy+SurTnjBLGP8zY
hLSsMf+gOV+AHWV6M9v6z43CN1NZhKyGEKENtxx6//waGRf/1HuPt4S+dg2Q/qPO
VQGXHAGNbXG0aqM/fNRcvoUl8uIxT4OKdR251K9tlvv+vbeHjVzumF3g6ZQNZoFd
L5jb2cxbWN4FNowQROY1/wHYx7HbFo4u+IP1/lEoh/3ePXqSET++BlsQkrfIXbGa
/PxZrj3ahCBXylD978pApil82XGSWQ90ur/PC8KKeZrQOMKq9vOmc4wFSaUCNwBh
c9Jtrua56S7C2sLR3wUxy3k1lmU5HQb+kge0M+CllTTFkTZl23VNRGL9sPK9Xy/k
tC1Peez91Y1skDfThEv8YT1Sek3/BAOUfl42/ldMLy/7F/qTMw94s059U+ZPlXEG
QzCJqgVsdFvxYLouhwVQpalVvHGGoWxAIuWvDSCyGEyylkmkGcyW4k1AjJDWrVtx
V97kHY2lXXun7x1XOz65vT4fyNYhjKFa8phgV4NPxpsFaIGk0h5vUdfjmDzevfv/
OxKMIhRMcN0w+rNdD4wBYKM2yBFJMrp2RqCaYVs1ObQM0BmG/0BQMobl7xrFC5ZL
d7jeRyfUZKlJRoHKWaK7PL87+7hO3IQUpT4GhYQNvIVs3uIZ3CEmeXEHiJrF6IlH
rJu4B61kM7RAkgQJenxMl1/MGLTnWOMKubpGVWeyZ9s23hVg4/uKdnDVRKG0gNso
Qwdjczj25WCtHw+S7uHroTizYWL7/05jkdnqF9XnHUxU9sbLtAmEzX4hViDV0O1s
RYch83TeXVz23s9B0Iv/RlG9SbI41LJfaULoDpNWbhR7jJI3T3GU04BZT1mdndk7
Knq7gLLfr6vym728xRC8545gUJUVtl2SIwTBNWWu6GCR5of1aTztaHSDPE5N94Vc
u6GDW9i9GOgz87P5Oyh/MafYctv26Sv7a+Fa9RROA1UZIb1yBiIUAlJfaqckYfMM
naWO+ricF2E5oZHNlxsxoOld5JCWfYCaP4PnLKytPNSfsUCaLaNF2hMQGsUymbA1
mURLjFohyPY7xfXviiSt1Ej5IzsIYij5QA27AQWXsfGC99rCgKCRd5bpmYQiV56+
MqbnFL/zpFtbJWA5POnxgBe902nr6ki8G/BZWyqwvG358yZnxI5tkXVXHB3VTGv2
EHWLxEkYNf2CL3J69QuGUYoBizYONDoyKf6PNIwvSc8MWoUnHtAw8oN2URuN6TtY
0DI3o9XmTyQakhKzrCTs9BeK2vGoJFVMYwPl7ZblAv+/T3OFb6lPN+J/3EzPSOx3
MV5K7ODBn504+SHuuu3Uqu3A8Y0lzRcdxX9u6rMt3T49irqO8u8sqXsV+NzqX9T4
Mqpvn3hHwiS2xIF+adNFkKy5kkcnxQZr9bZo6S1j6Yw7cTd7eQRIvKoe8HnfrRLN
zbLBRL8aUlUnCL5Axzjomi1I8D0gXWXFMxnlasU7Pjo5hga05d/YbEYG654HXCjp
jog9vEsPpM7vCsJhhOUXAi3ThQDiXV+Szut6wSgOtwmHSXLYZ0M7uuuEyBl2TlXu
vCKeIUOZ6FCEaQC8bnDNAbUWfKt2HX9va6DS6Qf5h162G1+wEGwGQshTpI3VWWx5
QK3CCMKpxhgX11eblAJ1/2uTAmEChV77t/F+EahG2wFayDxi8pOmLq0jal/jUzUX
gBvt73iTzXjIaOPzTWCCMkTc0R+27qXTyxRqEDe0I0DD9+GaZM6wuV+jQgVp01gL
AdheBQqqVaZbjQi/1pHwesLywKzbkydt+Bf47d5JPKEesvu5ylLWG307oqcHGXkh
Ip1uBjSBLpcH7ZYbrLa6aA62wmX+qzYqt6Q+V6SCDDnUQGLYbLzoI1wUdkQuQJd/
77rP4/p+y4U8Uj1faltDTpi107JjaZYMpkQu6W0QjPp06VbcR0iKe1+8lI4w0JMy
3U3HwZG04TEE2s50CVTN6+IYsyPFg3Yd3qmw9Zz4OYWGOfy9QP+f9i9oc6ppJ3Wa
AJLGBNPvDL+VLdJc29nTP2UsTAtIiI3iBJKwgmMa0rxoZXLWHHEtvdLKaoc+Q9Cp
zhgKlJL7RSdKHveYurA1XsDzb0XOWgR3giCe2UaUEzzMmWUWnvEkr9nid47770U1
MZoI43unW5bkD/1hmXIWJeEA73ucoasXvlGl33FMUQTNlDbMmDtAIb1qeeL/k3R/
N6D2RGzv1p7voTvfRwmjb43ra58U787R+1d7i1XKbjX8rAqOft6UYVZEd8/fOJxR
164lwCqZDozy54g+HyB/RsdNLs/x5a02oOYHjbHSWObqefjt/BPoongpG17CBHIO
nhL8GQLCgPoZ1ux47klheE/F6OWo6UAFbgpnSaBXj2LGA3V4JzMMOLX9h4o8iCAw
AOi2560NM9HOVqzHBTKKlcfhC0g9x4omMAKKgYH/4USWgHTVOLuDBmkO4acH+8UJ
cpRpoL9IW4WUU1plYRq47phV0Ud/Q1yJuxjGEzN42bPqMNeMivJVm2oUlu0hiSMH
GYqjeDgqDx1POV3X95zGoG65At3yl5cjyW/Kkhy7RZ9CmxV4uwIIf4cvYuwO7kDy
GppM5+8FRWJ67ojKxIjo9IP3U8l9rJkb+OOekPjXY2wUcTTdPjzV6+DhBeC1wT3X
/TkNQNhbjQdoMAQLMYwz2XqswchZKCN6ig7plZQfepJhmjQiK1S8xiMkK0495IrL
DNmH/f3YS5YohEYRGNrYVoVApNSA6nM/VULxzzoV8uvpFxUnx4fywUqsJPlVat6e
plmg3omTWqDoXf8BoNcFO+zD3Ad8AHScvHN2eO2qTpBM0EJMYDgtQq9iIp0cRO7C
ItKsMGZe3/netq8W13zbwtDolccmOBXkOUEbWKHF0uuL3zEiiePbWOm7F9m5l3dn
wRK97lualxwqG5mbERhMgcNQel1hxdj2IH5ZkB9h9hsAB2aVP3xD2yznl2oOt1Fu
6CQze6DKWAW0DlyO8VlrsY6iUP75UFS1By9OehkiyduXNySzlPHNEeo22VQ80vZZ
ykOcV06C+cBTd6/jbw93+d2iUVliQbUcOADdobbsiLJRDEStcnLBBrFDvbwYmzx7
Ws6lSRIKHig/HavT4dJcShYz1yFq5p5Vl83Q5e5Agqp84F4McgnbPVNWsExfdQfe
6EC0Wv7P7VbWxRin8XNNkSbb8rzLHiDrEeWPuq4aO7jzi268bLJxbpl09rQiPv5o
XbHzb2K8QjB8/i4V8UweA/uyaHUl0luKOfsN6fKurf70rPhZtex2/QLtplAXGYJj
+3M9m+dcoPD4fPRWjFM9a4omXTxEkUeBWFKa8uw1QG2nGCiSDXjoRcR6KOdmLHRH
52kWouX/3p7a7BzUB3YZvf+VqNCFNE4vGNma+LqRzrsmKvDKDNjv9pSSLzhUPaCs
sfobs1Y7h2BFg2imXjGIf4AIOrDV4wTQI5tPjt6xtOCdQKAgbHW6xrYAfxKDdsYk
iNVcujM5W7B/Lu3QyCwdZOSDJOoB+oj1yujdvf3fFkCkNQacuNC/f840yTU5kUtQ
4bxA1j/ouVwa6G9zsvxh432v9aMw6Un6wotnQg79X7AexG9rVqPX4Wt38Et8a0qG
GteneL5JX36wf80UP86Kt1JCzKn8oyyHsv0J1LXvcmkY3um+QLkBVoCc44SPFUfn
8cmPXdx/6XJieDjaT1TTE5uk++lBhjDZCKpbQ9ktD/lTLU9ely5U2qUbThEi6P5J
sMfotG8wdBkYUu3syB6Bg83shWT2zuo22OWe2hDUMcKEkep8D93UEU7iJNNIPUTh
iYkUvFJOzpIfwHzwSH6QG3eNC0XA7+LH4EdjHfz2ehtjsF7xdhmjhoUSWEMrGddH
A2LlzpOBjp7nQO0SPpfG0n5YjnWQ3KaJZt7vhYsVMbSD5vGEnftWIsfL5Sa2QUhl
PhSfngix23CkOBXq5+S9DbkEzG0LshMJTa+nu6ff2rs+WupKYvS6oxcxPlO+wvXf
SNwXJLUnjPct48v/paE0VaZqiy47VTB6lSefXGrdxPTj+tnVJDqdHbwii4va/hUR
07aRmFgTt3HG89AgenryUhUREBjDgdQ/YVujSD7EC+jvc4n/31nnU1usM5PBH2iv
ne0JAMunXOr4uVmfXM+hqWplgmJDKKTw30FNbzp95TW1EazBLGowbZy3gYZTYYlM
GFLckDQeo2jmXnRIJmNlzsijRskJ6KOfL8lHoTlGQOtcLBzSA82VWVl+wx/pAx92
Rz6lM/nSJj4wKKtP7YJLwQmpB45TY4Gpnvg5HJ4y7EiotZ7T1ykWJ4CA5mddLZhr
9iLPfPI4A4UJgWFn7WqYhTBkw5Yx2yO6w+XpxQ3/gP3APPXJjir5BgHGYbTmsoSy
GAzwJwna33tgiOpF9ynIkNjKrKcgPDDUAzOYjemxQY8MKRIK9I71aDssTXTQ5w1U
vjPEO9i7cua5hMzAEjpNiOICywstcKCn0vwvRh/CZ/MbwK1eSprTEd81RpkRZQEh
5eDrpR/wr6nOEf1sGANfyZgMi4fqPAq5u++lkQQUSK1ar92jxanmnVurlLDCEh7z
wmstiqxvU4jAO5Xly/txpztzU1ZxcG0RiQN9dXwj0X+eWsO2kxtb2BcgybkwoPwz
uA6N6K5sPJiB6qxFa1Cn+I83y3kgN1NbyNiQYcv0GLvOpTOW0FqPiCVW2QnexmSF
ycY9HbMFrNaBE5bdnAxkYTreM7smDrzmIZ/V/HV3A8kuW5sHs85bK6Hyv9aLl4f5
MC52mdqhJIGDDYut8SqnQFvkvlmv9YC0W5HuP37ovvFOTAiGHjWedAh/vS1X4xKT
Bbr45EpozWSN6u1OhJZVp5WR2P3Gy1DDQCue7VZ0JH0Qk8fuk5k7SI8fJ/ypn5GC
Tm0zemr5BJwgrHWtJyzzl9UShKkmxwLjsFrP7KrFJx+IskrRLZDDY9jbiqCKr5e7
gDNYWS1TWY33Hfl/XHcJfIvE7K1XaCB9XOusWaE7nfq5AeMG53zAdcXH8AoSNixG
79unlMH+AMCdFVnPoqfN8bSagK7xcM6JaH7AoD6IM/t/NciX4k96ZjhIcxR+sT17
XblY9+bVeJSgUZImsFHECrsaXRkF3dlQE9x7lzn6oiQWpcGojAheHzKIpJ9wNpdq
Yo0aHPPvmYL65bpngMrnpyxWHZVEcNQ3tvLoLgocjsQyYLcXiQmi93FelxhEQHV6
042rLVQyTKGM0z38SnKWMwPpJxATKCQay9vk+/dHS6UEzEGVDVeQTc9nC6q19NPc
lDzu6iO19JZFiT4u1MpUohFFAs51LUCAut3TDM7Oooj8Q7lWKUAzO40J7YRGC7vy
7NZRwe0VbVyWET7JdLYjbYpwXjMNrG1er1SfQ/bgeR+eK3sCaORiCVH3jNXLDfVg
oRakWAd0yCVtcPUS1wEKpY2HGlfxFGcvyo/VSEtlqxOsosmHDR3UUTLO4kf2Gdxk
prqhiiHM3H7yQKKQVa6836lXsV4JX2qPWZubXpadLbNbY2C0Gax2Be0lgK1ny2bM
tQiJIRp+tLw3Y2PL2CPba8xkzPO65h6JYIHjgDEq71kjYLFxtzPyAWDsTHCHqpBP
TChSVwrDOymKLwkDgBQ3wBEsE5Z0sYpTahXXk1RMiy97MsuvOqtlEf708wyqnybg
K7mi1u2XTd4FjnNoxI5iPivSl5t/wlzlK9V3Ou96Dgz27+fY/cOiEoi5RKiSPwk+
hNounbkLly27d9YDhFE0yd2YolUIWV0ULkI4WV9L/K8Jx/AF9bm3WOan8iZSm5JF
wfVQ29P4OAw4OX+xL197jjMNTppY1k6Ii27/nbc+0dEDJz0P3SYLBj1FQ5LDu4Ve
01W00lo12J0gFnI1Rd6eUqk8oZGhUrZDWZLF8cSPZ7Hn+2evxudy9dw0cktvHF7I
FIW7EOBqxFwx1MdMIgVs6cc/sro3rid7bxnnh3VjR6nlwVBMGZIee88cTPZbTrvJ
Nofvw5R9fmu1QeTecYvb8huY7kU1IyaGIdkCb5Q4ctU6U8lrHh9GZmgA2Fp2tzDe
7KkCR4GWzg2RCKxKqXaQatduz6pwbRr/DFeGjlqFKocF052AONAxrg0ry1UOr8o0
/fXd/bGs/0F2+PQEgPKvKR7uXFuu4hcw06k4r4PxYEl1OZbZBNTfFElEMIBQtayT
Q/byDPHLxd6zuYa6JRstFJI+QvryKk7enIRqr/qIc65lxu5UC50fgh0/yMjFEkgK
6aXJuiLXd1Nua7MDKbINSr5r+od8f4QHGvTUBBhOvySfrJv5e9GuexkbGBwkyu/G
yiBje2hrYOEohB3FBHlGNSZ51Boc4TNQNgymFOwW+dZK3VOGbJqzch1Y2rmgVSeu
zL8iAC1zTttk609yH5WJt+KNgt8RMh5Ye5aOTcjFLPRIuUmRLUkhnKALptJdA5PB
ZHcdwQNBbo8CIW5GdD9QWcYPxEXMXvRC8CHeYIg7PdhNi7JJKWYYYu2o5Ay52uPT
7Nbt4OjOS87FRSGg+4CGwD/1Simy7gYH/jt+R5uM17hb19DNUENyA+Yw4YVnaOyP
91Jn9b0liMDS87pgD+/R/qs2AqugN1V6XBaMgSbo/D2esMtz2ZiUy9IJ+Ads+aFY
kCucrTSPMh5UZ678Q4IOdF/ppQ80C3utvTHOudTo5QQL8Zzpr2Y6oVkf8LR9LweG
LqO7dI9/Ce75xNxB1u7PAd/JhTXQWch/4EkHE95iamztm4fS+ab+fSWF3e9JfYbE
/6JhcFp4Wlb4tWig0GdLDS3nP/L5qUtQNxWHe2bQfzbMk1bytw2hw9xg/ETeW0xF
WhIiWkpqtfkUxcKuUty+AnbFfmRp5v8IlnaPSjKm738Yhp7OQdcwN+RBkCnP2gXG
lZGzXxBb0oxI+wdYrD4FPvzrx5/0UgjpemhJneBIxKA7LsYP66c1+5UUam9Xn0Jn
4EDcS558OgjtYjivDrDz9nyghIARSdNPKKZjhcIbJmmS5BHH1zKhmeGPg8beIcGt
hlRHywm0/PBrxk1KwUwbFCsOfBaFb8r08K0EdaygoLE/L/kDI22qS6y/rGjZrxgv
YV4gMjARKz9TXgOfcallmuBBCg0IrTvgJ2jy17v/6nXYDSDE/ca0Jf44aHs2RQMU
0bUY4wXgfHzEnKFIn3KgeKbvT/rYUMlRkf34Hz/i9WgdeeJ1mVLh8GWZYMDwofZL
j87xmZ0aADkm9nugWGnUhyoCPvnFVSb5behUgtEDsgTDcNVGWdsyNC09c9T8pJDL
agTI84lyaadTj7R+MCjtbasu44bZtyLWI0Km0JUiBCbpeq3aPI/qwVCEVZoXKXb6
BUj4kSJrNZZQWQ+K7qx2TCEB8w1ziOON31mkmE70XjfKElf7jBren1RmHJiLt761
XWYd/k0KyIoMq6ZdkLRJHtv/YdbOqXXjqg0zhn4bqXHI7Ahy+JNVhHBed3ZxqSBB
f6kHwLdG3sItfk/WlDEbYz5de/xWm06iB+W+dvtwgh5EbFFTWbQu2skHr6oc5LZs
LC100ad/5C832YbVc3JbYSOt/OagX7fTR+VcPPYAlStOLD/M0lMR5/9JtQJDlRXe
NwleiL0yD5VVzxdHGexb850XpwZslwNjhRkB270wgbVvOUl2bWw1nY7Cx7kVNb8Y
Tt4VF8BcyjvLqq+f9bFjqxDdljUg27jsnEAJTa4jy0fX3gHi4nQKJNGdZ6qG1WvL
6B7TQ6H2my2xnZLwb9QpX0+3XAhmpdJ/uxqbFIfEwCwJC8nfNwBDkCtM/OP7WPXp
k+bFoQA4LMfBGSiLA0IH/2zitwG+RllRXlsHUBLIN/ZyOeOibvu5tU/L6/wfXmX1
0tRx0Fn9aIpJpvw7ldi7wML5qOayL9Pk91/Td1MnCC+JlxlkWT+iNrV6St7qYLAm
t0QiclzTUDfK1Q0FHHbrKBtfJXxzhadPtUVgrdkLxwuQ3XfQL8ugaER+dKytPNhQ
07ubbGvM570U6EZiIQiENNfaoHKJu7tY15SnfwHE+5ssNsmVIvUAK7NBosb6wH+W
/Fz0DTPSan1L8oKIPMDkqonAS4MCu1+IXEPaRNb/YFvx7rMR9nt6+uFQrmPeo3dW
Cpt6xs31EOUKCW18MakQh4JHGAUmJSwzWVUGIS5ozpQGsBI+l6QD5ElN00ePRSSk
bFlNYyCVhEWqy2aQ1QEZxc3e6xZBZJcelLFVL40ZP2pf4a07mpNNTjv8RvDHDeT2
aLqUIOd5NTxSz1V9vIhT+1fxgS9uIPE96M2gR+cvyCnUzM7Gw2jW45/xB6ju4SO0
AzV4/fi164xAB2Jdld0FX/vnZHh9G4OKMu3HU2jvy59JCVarEdTjDsMUoLHDc+fH
k3Y781j0DMBW+mgp/ExcQRC1KZjzVPwymdMMqp7s5lFhDTgJ0NH2RCkrX4Kb70b/
52jXBn9eEED0sR9TGDMTUA1EAsehdM+DsTTrqi3F91V+SOTrKFqM+rpp+qkhgHQI
+oDowPE6ONJw1bkdTV2TK9OJXdxxTBpbkrAMkfXk2esnEfmL74xV1q0qReOmzT+/
zHPtN8oeis9IDSvdF9HeH/p/+C+h01N374tia355a1CrbO+IYh68E2NZNDYdt3NJ
jUNd79NLXGafs2eQMwC5nO7+KfAd6a8GHMG90zY3doa/VO5zOgJQL3h679mKQzQJ
1jHyUikTVNZGUZY/2Oyq8Jid4G/GKUNRcFJD+qIVxTc+NPxYw7s67PMbLyLrqH5g
xTPcjZb0QPidDgx7HZ+SG+Oo98bLgPPSYZ3nAfQOJzwWUX+cZMLrs8WMqZ2cP4JV
xELIjxcjBSLL0P7/51GM6O8mST/9OWNaQTkG5BlofCGxgCwiq4dgGoKhGsRh2LJV
TO2mstH5TOuKgzqchb4nzp6nNGimBOMOohXoGEKEamCM4R89RlO1GOpUYkDnUC7E
a12wn6lgVrMDwiuvx1VzyW+QpYoZRfIwcm1Jb5bwqJH2DBSZlMOgVZL9hZRVjG+A
dzR/21ENBxtSf0bmFcAo5gdqDHBc7MMAaUgj0l8zfxHD5TWwgwfyEny6/J5DLtnD
/hX8lcU4eydMA9vOfGXNFEX24G8KedxlQXgWvsvUKamhpAAIUjsemWs97EVQlTSV
gw4XKhV2rsHHeVHFadHSwAQS1tL0D918bJ3G0RuRxlRKgt0/xaJJ2cL2sgx2Bxqj
VmRziK7ScsokvvyVJoduvr38spW0CAIZImUnhd6fJL2irqXGoPXXOHHxmO0pZ9jQ
tGe6drjBwnvr278rhE8uQS+bgTTKB2VG08Ec1zXYJ28UpJE5N84fYdIXQgnfhHWE
hf57ecSpb9jx9ng+NMNN9tko73R8W+QYFcIcw/kOP3bK55LzTmTlEWXdGVS0ZoWZ
+lXtu1SBd/LY99BnFUYbfoLuD7E7qZsRWz50E8OVBNmTTSg2W0Ga4G7lY6n1QzUi
Hb371z0cvUxYAzWyPco4Wn9Ymv4QhWYnt3lu0ovoNQiOcLQvNKKuPhKKChun4NsR
Xfcf3dLngxhQISV2M9Y9zt2ThP0xPPvock/ZdB0jT6CRPisi7wueYVwk9YM9j35R
fbM6I7vWMG1XBRYZe0axEHfi/xiT2FeW4bf5irvtHyr0499CpTQj+8zryZs3+/4f
en5UpijhwYnpGUfCIEqNT9XKX+i7K1C9sUY7z+fWJSr+NS9NH6ft4BOsFVK9yjyb
vfRpVlMHivhwtMz2o/GIMQmzR+rZDKV0FqJ8BFNxAxzdRXBj6b248Yn/vWTlIp7E
H7nJrWVMr5Kcf4qPV/SfJBxH97RLQ4OofEdHw02d6dewIUf4Ju9CwJhrNdONyYVg
2nQIiPoLhO+qfDyom0hXvHR1CmWCe8j/QueGwQ7xFfc9q60Mtnxk/x05uvQ5pRUj
bNDJhQZBe5CvEviDF2BLj1gz5LjdOg1TY5K8uv+5ZRfaZEdYHGp0zCuXFT74xXvU
mLirOhNN3fNn0cs4j2zS3OVedng8dX8PvedvfNm9seO7NRZBD8ObobgUMKZkA1dn
GIoUJzE2kAKrI4Ilan1N3hnjVUSVrRiel9YjW09phkoeZ4eTW4roxPjQ77fOKiQ5
AWBBMw385jiILAuvC0aStUu7vtcJLdgle+k8WGa7cMTzq3A9U2f8HYl7qWfCcbtI
/IR+Rllj6DWKZPNtf5TpYFpMed5UcPNm2TGor0FSX2FmLKwIT7Ppnil+0fyam0JI
b2HPgepJkgW/kjT2RNUjF1kXd8KHt2O6fex3Z3exe1XDyYbw4s7XKeTA8Dj/+ZiG
k9f0hxReks85vSR6h7JWcqUbIdeWlIWUnXnr/tVqsQlo4I0ejyBI0ag/ryxuN60n
Jp8LmIX+UPWGQQ/2ed8B8uZvH05eO9tWYjN9Pj8vl+TZ0StXU7zmacUBiCV50Jxb
2tJocZYLzliyPlDu3wAWJ6irbd1kh/dbc8dnUnIiBzAWBCeTvyQzU5UYlI0l5KhL
ldtYW8I8quCkqbL0ozMwqX6+sHHGJuvx1VVhWaOuB5OvHU0XerPOYcspIsbyKS1w
TV9y7ELTTR2B6bchDtk+4pOcyVLxuJ8i51MG03uv0qDEzO+1vYJA88LMqicIl+Dj
IGs8TN5G6gRkcwdWlHZQ6vSpUykIHuLtOOoU6TyOWoAhcoelqRgFO34eLtW6upgu
4XDhBTgNdlGH7SzdlG5I8YlwMDtZ9oxeWKXb6lkodxLrgEM98ASU7Vq8mgjRu7kE
m0oy09vzyeWUUtD1oHimjoYU8UxRlobslBauMi8nwztnHEgfvfsd6I532xgddUPH
nQ6SZp9IocJlR+JhhZZuH+yrNfoSe5k+L3fTB1HpAUFRH/rWgYUFx9+YlN1FgkGp
g2/5CDwVdXf0wDWh+rBTlRGhe2dnIPMC+morisJ7txjVM6+vN6Qv1yqY/40ZcmoJ
zEQ+JlrXaGeJ+a6u6L0NDdLtMizo7HicHbfzDSnSnDwepdafSXc2uDE2Hc+jxfrx
YiExr7BSGms/9vWXiahwDY44VECm6tjqIpliXhhnCG+jXVrGNG/oCM/ruZPT95pj
BdFCyCq1uGX4eybrSn3D1vRmViB8NhDj8SianxKrJSIq4w7UaY9XK1K72N7P9JhB
xj/12mmBUjlvbBcAxkgI16e6Rn1ucx+4znAG+JT/s0KY4W5xpmTKiVQe1Bo7vXyl
Jo6NkTkZP1tMa6Pkzqa+ZpPbSd4isHun3WV3BWeiZ3LMR8tugWZADc4U3CRbM+j8
tDyQzb0KrehMtDrQ/bdyjUvKFDR8H+dsUuD+/VK7q3dNnFHC7s/yk6BoZ2yi8Sc8
5BJESnwUPbplzYfB2uG4cwT+p6iEzjUgguW9NfNXmwtAL30OO67nuhdXyGxX3rv+
ejXaT+kIM1SWyIAMP42hHKyj9vgyzHgIQnh+tErxG9omUpKAd3XmicQ69cDHelEo
errEi+d76R6homQwwUQXR/CE7RRogPFKOatBjamjxSWhARY+GrkHIbOn6Xa1tKPQ
oqkbCskFW3VrcCTr0PGVR9GA6CoLoC8M7YwGXco3Cn8908tu+2h/loi96YencWMs
j4wtfprUXHxQmHSnFDZIXoSmbaxoRULX2BmON1Wjh4r8Mwm5XktRHktXu+ZHIIfv
82qIJB7Uj9mM2qkEhSf44toXnavyPeiZ5Blb88iNNE1vJVMuXileHVggo0do8hds
+1phz34zTBUo8UPY7nLu9nTx2pzgmt0SVkUx4xPilszyRmFD+QdZRaRxB70XWS16
RlrgOkb1Gupw9ChR0Jyo00VyI6w64oabq6lVqO8HszOE8Nl8bhuc3MMU9a2J275F
inEQ05kSen7LD3xjW31p3T5fnp0ASPP82WFkeRWB+75pUuo93ZwsEAUqTbblSvZ9
a7/+sYwTxR1PlQDMO6xjN/fAwNVc8A3YqjroopxkOrQKLgat05bbiYvdM4v3aRZi
S/BvgUBruVOSmWJ7AF7b5i+xHn8i2QXJERyFHW1cBMRPANoJYo5xLVVwuOtdttpg
ii94jDXrvfUnH/WphLJY+e0KXsgoBKlarP8mXjdQKh6RXagOVsaJRsL4ffbivSJB
AsVuiQ8q8JJfmwQU+15Gninf7OIOfk8ai35HlUkGN1m5I7kiHDdhpgWscvcJXWIv
+fQlG23Hr/BlMyJo/OREoYjXpxE1cC7tPV5X2thklf1ibTeeKAe3y4fukd5tEqWt
2rMEZzc8KRop8C3Z1g/lV0ehDNNgvPY1BRq4VC+Cf3P4QrE6YOP4a7lIwKgeSrOj
SShCbd5Hg9814ArcU7QS8KSTx5R6TpqDcdrfrMrrp67YzFfUYQPyErkO6rKewL60
b/oMBVorqt61AQtN3TaTfCruC62hPITW2E4WgRiIBXvmp4v8hdONCUoPQcPld1hV
rfqnHYuqrtCPEJmbbsJIajgHTFEc5jEx2kAmd7l1QjpMYMrJwJShxTyrkggnpwj/
+iIn4IXidboJFMve6KhNI4U08NAfIDd0zIlZwV58SY4X9u3I6pGLi7yOsouajnjW
XLbeGAahp+bIspXfJzjnPupQvOuPNyY6gHQO2XcCFqZtIUgR0PgqhCUseQCGZEd0
KazIWWN4AnANtJW429Q1R9yugcfC0KvcurUk/ADLn5bb67BIobEPktdnp+nU9Cbc
PD0ZXdnLc2EbLqOtFEO4q7qawIHcXTtj4lAmwzAYyewjNlxYH+d8Ddbl+NCdKpDM
rMqkjwZ8r6YPYz9i8UqMjmycT3xUR5eu1v6viEyQyaI3XDZPKFbheqcwYQCcFhoI
qWL9w2CQiFyNLUFB0/tZXVkAULwq17hrA5GfovGHgoPCz2l6CnZL3ShgNzkvBUdr
0yx1fsJyp4kv1Hu5UPxKnzmFCce9nvi+0LtZYd4EJvSkR4POWsvsGW6JgAAm7D+9
cWraf8oFFsJTiOBxXiXoIPQl08lMLc2+TN0ldkH24u+JL9bevpnpEMwmDxcJoVzM
ezvpX0H73iQuFNNORNPDJPwU0mOudb7U1+AFLXn9zIJdFtmgAC4mSoOS+YlB9PTD
Ld+nr6L+XKH/v7AODo/3Zb29PRWxYBoWa1JULI5B8fTlZ9vd3ug58+7rxNs1T7it
q5OICzXaZQxC2UBe8TIZNY534RRZKAejqZ07BN0aMsoliqQ7QSYciJEs2kieZJNo
iD1lRltKUtnNxbzTUfraJEoBMiCHxi35OxaFbhvGU69PWFTMhgl8GlH9AStyVC67
jv95CDmAiVdmWy1QcRIi1KhQRuSIS+Nj5Ug5x4hspVXjZ6ziNxgpCFOo4GIdt4hm
NMSQe9yVLAqkhz0cH+otuEDLThJQogxPfbJemyK/jjbeUtHFPyFY5lGvheGMI9RB
utPFfFZa1fTWOSdnwLyZSX/z2BQ04ASfF4zG+cohwfL76Mm5O8AlkPv1pf4TdFyy
QHP2j0UJ5G6H5DWWFWztfMy+Ut6Ks8HbLED1lc4vl8SDUgieCQqZnB6PMoYNPxte
y60VAfiKN5UtQq4t4A5XJqzL1kwjevsQeUxFn10I84tPerGPa637Jm2RzIne7niE
fCSU41K6cVEmmmdkwD0aTN87I21CkEwVEkbIQ2BmgYmx3IgfV9qYat3hXvF3UoAL
X9X1HBfqrJJyX8If2aQt207+WTRSYwbOP9jbjNVmJdNWcBi0fDwENpFf0GpKt8di
/HsYeOBNmTPwFhbI8Qm5iJEU0MXbOixRfoyqi1yLC3psHSlqxWFyNfb1aCITOaWl
fuipEQzoRDHbN3ZYrX/jVaM2eJjwIOQVXyPL/mKWo+VNRP3hqXFwyipa3I7JSmIM
8SH0mt/b1JH8mQR9RFEh9LwsXb/jmr/cfM3QDjDQNBCFIRz/3RVpbR4XCUSyZX6m
e7sJKX2V1rXJehfTzp14+hTjW6cEEojINLN0VfiUMrToU2YnDH2AzRqsg/ALpEuY
xITtXJtqMj5BcSqpI7jKIJqcWTMolNRTXvSbEOJX/VkKW+LNItLQlNoPi7Qr1Bvy
MtlOa82YuTxu0YnOl0rOYUPmCNb/zx5XPIOpzbq54LJ9egytADov32WI/aq35ISn
xgrtlSEun9PL8MOja0ozKYe/SMWwejTwYINMStzRmWaTAdbmjuP71JA19CX9IgQ3
f+Zq6dthMBzMWG68+xDSXHTx5qw06p1ZwtKuoFE90s3Gzl8s+mmprlfZc/YPKdgk
BjcAnmRazj7ydOHwVR1Dp0nAwtKOc2xKUfAnD5qt58qFL/mvEdGVA28h/tZv3dzo
zfiZgdDNY1NF6VeA30YkXp/tpNt4scwYREKGCZIE8fqyST/3TjBFvnR/OzNDJCuG
N5tPQTKCq/0pEZZ4bEb/fcVF+dX2p4p4XkREUu5Qxq3IG0qpzZFyu2YzPbBCWToz
y2eRfcDUdyOKhIk/PrrkmlD5kkWzDfpj+Vz7ZNugQeRt9VP/TzFFWBPSzNZytnKR
0J3v3B/Lxi3+09rPcQ3aytnylpoMEkmA1IFU0kkivkNrv/pRo6/diK5M1gadCixF
XUV6avhEpRpoSAoNmRKw6xDsVKCTij9pEKA6SOB1IV5oej0paBbu4MI+wv/XZYbl
d2dULl2XcBiTh6CClIVfXP9zmcUnNip+3OgTCWp1401CHorPkXww/3uxYqseDOks
0oCjasIsdRTi3QeWaob7KsSqQj44gw9rnqJEIxQXaqmzNl8/JedR4kjmM2tHowaC
o/paWWNaRStJ9hbh1E6Kgq/NzPNBumFO8EzV7hJW/WrFjss+ZfzwjtWGNMdM547f
7R622zxZQ2BapdDjeuUGqJDWnWGrnxFoIMxqUgFShvZPBJQEfw3olxr9dnLAVBQK
C5xsjYjAldRzRK46otJrHN654fclMz/xWancCiGg4JFNlIuqMr5j3OAW4gyOqQBR
XYbJxCZWDA6thshdqpOs1PCV5sv045fT2BidzMgQZPVXYQEOxrH9xoRJWhMOQzvs
7gx/+HxssaBv7tA6t38PZrn8bPjDyQR8Z89htkJbCMcEZl4qL2Ns6c84QzR8/fnA
/qDkNtl9GdD6kKILqCcEJoBtVYnantMWOfNytyM++NvS2ktY5UQeeVPyVxSkwii2
HKurP8Lbja3QBJeeW5G6107DYwocrN1uxQdQdukfv3s13p9qgoHdt3+oWnXD5ddv
Q0CPyJBPdkAcUchsySGeYPYLqfTcg6Q6jraY2jEq+4cOtE45JxGJ0B/QqjVsa76I
RqEZrP5rKriwRJIO4XxRYuj/LJcruZU3R0w/a7RzAZDf5on27spP2oFZuUxeUVR/
lcc+U4uLQrj1ir2e/eC0zmPaKfgYoAf20ORtitrnXakPiwM7vBW6aOt7nTkYn4y6
+U2Z2w/J5STxyN0Tms7mGwqMgU+msx74N97hAeXwCPuuVPyay2N7FWyQ2mdYqiy5
tHcyLrwcGxG8LYpb9sv7eW9ji0QDASwk/vBpRu+cBnWi5HiK+ZYy3DL8qka/Jalx
O5dTY3YaAjNeKuG3ngPCCYeAOXfrhiN8K3RVVPMoYRAKtWJak3BnJ7Rddv9+9UAQ
HswWm0ShMovToZq3+CAFPxx3+Ox8CME/iTT6aoguQruZJ8BzKBAoZQTmZJhtcfuz
I9BEW3Y3kAWqVK0uJtDI8jefOwgCuShtQlROP7oR4FrDH6J77K+oGHWOIOqvgkys
gYQfFYBcmXs8ao3sCh9o/eZSsJSy5EvyJD3U6TpsDkKF08wIRgLk7cROp3rggfau
xGdbSinwg9c1Loux694tKX/9D1m1cna/YW/CC+SFAf3ZvmG/eOpKlU7jxwPOizsl
m7SaRsW0kuPFhJ7xpGDI/rQEgXzJzA1T8m8pwtiJDuLzkvPd1Eup0hrJUg+Ls0LH
vSyjKPJ5IP+fQHP7nNhfE+XKjH2AwdU1ADApAfsbgy5otLB4nDmhMom1V+z5VGs9
sznHp1OOOMwywlOmOaxu1SCkr9FLjo0i2LsJxrEAww4+eNhQtfBqPoTtrqn3HvI5
qZ/yi0QdOBRf0hKJWhUZ8/lzJq+DOpX7vjnMOxPyHa5d6xJZhKkoXfXT3Ilxd/7D
2gvJlm8O8TCdNNk68BH9loHMj2ZrkiBZjyZHci04GHCkNKUswhiy8flLuROo4i+K
sQoLHO8ujC+YsR140z3sfLBE4Br0aR9eWERrYKmmdkuhjonpJwCd5tmukLJsccxI
s2WhIkm+mL3ZsBThu/zj0bMcJ41MjdEQ6wvlfAvTWsjPO29fqks+w5p4bsrCjJaO
XCVDeEW+Tgx3mJqQooIdxuq2vf3YgAhCvaSmvJX6soXt+XL3/XyuL9As7S00wnxl
vlG8rV0D6M310AM+3Y+WVeCnMOUoqxNXzfhdpAKsxiAm8OLgnel0g8kzT8sgJU7p
v1SMmfWH85+rxWOIp/k8Nt/ESU4XArKJJh9hXsCQ41KTLLwD98J/0cxRSzAjSbj1
NA7md13ts0MSgvSGrlxRS1t+Ndr6ezGTAOP4D3aZ2DxKrse6IzpcL022pYT2KgT/
+ECVh3akkjyIv3sSRNk1GsYoMxXfrB3RrvAj8zTgGKd6ki0zZlpahTMQf1NTFO9g
x8+Q4+/9hZo4Ay/sQTOHKZEy74x6vbSAKIbnALW3a+i7dpZEv8EO/ikJ20m8TrjN
FTWz1L/tMuvP+0thqgju0WrbNXWb87U5DwXV15f0MWSvSeeRQS0Qf5hWrKjcieCv
thNu3pc7fQxyRHLdFQ95KgeayNLF443cDySIgN1k2AUKCF4qqdJDuhrCkk7EiSX2
2LyWxGzAjEitwjNlWrApC7OIetUBuVXfndDP0gRupeq+P2uDk7GqYvRj46qD300E
wt7d58zK7EZDOvqwFnLYjrc/LnNJ3ZCJttlDBrNnL41zghY42mcaMoobsHvQIWgk
GEIum4ItFs9MVvphl4jQCHDlM8MszEMzWnj8Sn+o98Bu6WgM8s4fTE/hkHaTp+ip
UpDE234+mGxLdX5Uw8U6FV92wP9PcpuebZOYSfdTiSraiiIgoeqwKkrdW6usHpGr
A3trNNfJkhhBLIZe2fiKqjb5dlDJ6cSFTMESxamIC3kMXXQ3vEz01DW/jJ/AxhEQ
LOn7fauj0Nl0TrlQOTNHm/PojuJj3euASXfu7o34XmIlDI4ZLXmnrXMm7+FoylGt
TSC9R3BN/Vw221DDI9bhFUtrVfu0d8LjGgOj4zqwDcJCLbsYMg4JMjUG3/fhHBRp
UCjqW76Dm9Vrh0VrFhNKolMiZ5XSBtjLTA5RBDGQlM9VuYauhlUG+F9COgkMsgfa
OriLZ7quCJ4yjZumH9uOSpEiaP7R0CjbVLJUQZ2Caxynw/Gilgfj2kydRaH6i41d
at8+UJn5jdxDPxO+EgqtyUQu5U8Nft8r0UmweagRBIU9hCAez3tTeLOEi4eUUJiZ
1Us+6LnhjNqbPyezmtlcu2PZsfx71apkEFf6PkciIYUKM13s/ncZdTS3Dmq82FyA
oAvHIuYBNICoNn+0lSJb6Flpsrba7QARrt3Ofq+XuvyY8bXaIT1AgfWAUlUjj7RY
cQJKps6pbek1zQzVXAY442L+QXDkhXpCYwOD2ku9mCk3gtjI+ioYO5me606ruEry
M/GBFVGvCt9rnPTTcUohx+JvuTroXagdTwi52xtFgImabwKbCRvIb/DtT0CN5jdx
R73Itq8HQvN6o4zWAcOgcT7Kx+8fjAGO8aqhh4Eol27FH6ZyAfBp0SNhns02kvvY
xSyaGJK2w3C0N6z0JRouWVEcYVfP456UqcY1TUf2EPO0o3A4O4tvF4H3xlmkgCi3
SSe/2awKgl0yWFYKh3k8Sk4DPwsAAPW3HimHf9jPWSKESl9WzjYwlfBq70Iia5H1
ZBCnYgebEXd+3Fs3GGlJDvdoSL07OhR8L0FxO8zIx4mF1ILdTrl/pM8Es+oIRjVm
7Dk0ECZw/qSjWBsTe4BUjnf++m7/lW7I0yjMzArCe3z9kr2DhFFaO3D+hsWC1rl6
617kZ/5+tVn6yHl+YSpbVXfqPSmjmnTAXmWga9OWqocd1zKDOCktqgDgww9PNJxw
ek1szyviT+a2z9d9ZOFbCTEWYwCIXujJ2EITSuRSTnhcJTFNKtGXYnMe8fKNP6Ss
rzyYehD859AgILfGncdJA8NAK+iNI/bouFImork0ocl7R4Hp6MpcgaT6QZ4ty0iD
M9KPA/tJxtoDhtUElT/jlTl4IbEUt6ueyh8njO5cuD5jxS8cq0PBzT+A8N7iixBt
d2w9IYrZdGeezegeYXU5Kw0d57ZsgiqnRZu03z9C8T8RuspyzAMWfeLTPOJQ2c0T
zfxQ4xLVzA1a8KieCiUO7s1mQNtRuv3W3JvhQfV3uBpy51RyqOl74phg7gDica+g
rXIl/AqnN4L5TxptqJeccue0qzKAA3D5zjvq6KBv1tlIMY5f2Bn2WdJAiuzJELGw
IH+mYY9AGX1BzwSN0TarHzXV/M6CXjbAsbF7X2UYctIoWpLi7qKhW0X2mBOJ2cH7
BccFiWqJshTs46buJkRF28YJM96YnTz/DiE4YLVTyGriyJfVYM8fwm/mArUEzudf
2EVlWt8WGCeSVeBVNxmEa0plZH5BenrgCwslEg7nnDebzEeObagPMDM5QNwKntnv
vDl23sYw0Y/tQQF61wMHSMc+ZGqbFhkl7rFECfL9nhfEKoAdwlXTHj0SYi+1XDkk
v4hIZOkm0cx0eAa2YYKKh4XzXG4/Yef/87wxgxtpUG2LA4mC3AqAvfJtTFyF7s5L
HCc1KM41kgKxMxtnfdku5HNBM0fOMwbyAjbJJ59BHOUGtmRI6Gy0zv2aMQFuNKcV
AjaodbpfzmX7Lak9MgWtALNfA+4GIiBs/eVd/mM4vZARm2rfvHYXtZBZgSCqCMXg
jJznjaNCTSvo+d9+AziF0ANGik2xbzij/mYttce7/cqU4vDJ8/zhy+f9k6geTGOH
rAuk0FIybJ654DY8bDTHmALV1VShF6o+XXX4GhAjrcPy47Y9nHLBCVf44q0Hk6CW
f6d2d9p0R4KwKbtp7svzW7p81Jo9StvoP5dn7kZeTCAmyIEKkeQ8DNSCiQ+caoaM
0coGPRVlKqD/PiPIXF7qx/+DAqP3T4gWsorVOdqQ9TgEHY2GG6+Fqsal3/ZQPMDi
IHexJpPb6aA99NewGWAglmcyGBhgkLWlbz91lqRgV7Cft/16LVW4+ZzdEdG2CUBb
4aj4lKht/Jh3nnPPTBvjlvguXqvxlGKjMC/h/GMnVI2Y1bMb21SKNoYr62ITZX1Q
b5Br7xqx/HFts5E2CUqmTxJBkd3xxW3Tfazz0jiwTAqCo6baewRyZhKRmJf0aYd3
lP6Ah1xOutlaM3xdE2jrJSf+ysa4ipM+rJC4Q8fvtall82i+BX1HjBQdFL6fB6Uy
s/sTekE4d2xM1QARL+erO8qsyonatjy1GAdtBO8BaZZOWZRB9xUH8sm/cy8qJ+Tt
W3V7Cys41aQQLBtMeE/+HHDVVtfU1LcN7pC4PNDyuISJKa8oUA7cI/GK0i+eS8jY
/wtc3HLYaQ+h4dHwNU/15GmoMV9c8+vYBXfS4cVdAj1Ew+lZxk2A2qRS318/nDZz
R1JRoseQ64oRGlyVJdopgB2IrCQAm9ZH07FqvAGkCxDkTBE/zjNDdRoIPVV25Jsu
gtXMFLS48awPpSkqv4ENz4bUuZq88hgtqRJVmSrfAyvR4o/EswKTKhcRIiJ14g1W
7BqOW14KMsHTyXYHI+WvfAjuAZvNU8fIAt8MtrjRdVasfcIkFHAxDQlkUDZdjff4
NMDr5k8atN4LJNYSJNb17Er4tbw0N8QMXIcPYeHSIoaW7GW/LjNvbk4yQvkm23r1
DjPBNcyEpoSxH0TGOb7Tj1kTXZrl0i9d1NMv7YfxCjM92+IDT+TZKtktx/UKDSs6
n3eBUChrq0md/enXmjhCxpk+DXTfzAmz+C+Ju4FOM/GpVifnFF02hQrtYXLNHp1r
NdYPXzeZnvaHvTexqpk3aMXFIext/jxE9LkHQIox5zV4ns6hfLzFwHOI/OxzDNpz
RbwdUZ+ZM85hlLPFuuYhA2DScioLNb9YZhZAGpZxWkrtVzf7ttR5r++pfpoFHTbE
oPyQoFIFUX9M9OlrNnPCLmILg5xeUiVq4BHHHHzZJSqaN3nOSBC+VD2+YagKIMXU
dOm+RGhPrPoRcbN/gnCDNk2Lb+7dXMO82AVl13TlcMVhCOHqPGD4cDiBEyfkvHDc
tQt6j2FIERMFKWVijklhBOFK2XGi8zl3qto3vdNtlT1NAjjT/wf2u3Y/csSmzHsw
uIgv4oaj/RwtQ625B2pgwpFQelnv69dRvK/PE9x3k7BYFKpNlJIETn00F0lCbbaa
2pkJJgWiDolo31B6SS43did6AUDGBieRgm3g0dzw77G+tiFBuvKBcIG5g2WlutkM
3na5UYyXeoi6OQhLbvFVeRIECoC4XOwu8RrNdP19yrmce33a97/7JDZ3Anyq7DCs
4GhCzQ8GPzqn+HE+iepU7Dq71wZsHhXSSadcvRiZQw1Xxz4VvtaYXSFqPT41nxS0
jRrcSNFgZ9IxYUOSX8uoXPuzXB77OrqwQalDG9BsfTgyxZQ+i0lFxxSrtFhvlu8E
usJPZOoWdv/BOvun6OxCa+2f71lnpRogZeZ5rnrkUUCNH/uKPxT5309k41yJoXtb
9XRLJdeTQh3cylb/sCPFszVSwerX23N55aCDbQ0IFrKtqkXgbHo29c/Se5m+kcwg
/ifDgEBtSUnhHF9aMuC5kpw6qPi5FlrFAmb3LAdW3eYpA3eAV6PPAXkrRptOD6ld
gshzgjposYi8FBHal15SLkVo/lsXJ+Oa8JONz/IO9ViYk0p0wQxotLiUrpxYtCHB
DDXSD131WVwYPCjhXmdeszaeXeQzc8I/fnlpgMCZ5tYADSghgRxVO3Mx6dhrfgT5
M9UTDxv/ZLXH8Ar2BTr+Ht8wjPPQkh1OGJm3zQqqHepGRkhOCpXAiulwYGJYE9E1
duLvE5OL1AYkvbjH7nT/U3arVcMXe1Ia1q/hTxjoR+vguY0QoElHPC4zxfp+OO0s
L8tWLSy7E1xk8448ksK+rOXHfrlubWyEpETC7Y+h6BY74D1m2yIFpsGKdj5eZ4at
P+c2F9YPXG2kwweGBmpLBo9sB7/mQGiKe8djjUI3iN84xDSNHzCayi02GTsaB2Xb
tO2iszn1hEs1QX7e3qlaETAlKBXv1pm6uKeQYptCDkyEM5KokvFEZQw3TWCFNoaI
7jFWpTDvDL2TuF/S1WwJpdIbLaFELR7aFfZsGzxHL6YQgVacwlA9bwb+EOpzqcgR
0Qgoq+QmZcrZwwzeIsWZI7rXVT/xtqVO72EK+Heui7PK8dONstTyVJagIJAoqXei
jaLMKZkVdrCJs57O7iHMQUUIeNAhn1a+hA3/XP/DxNQ19MtEpQ+nPrspQEi0QYX7
je+wThz8JnL6rlRiFfnHeKYUF+D5KWL0TRFO4UrNzK+kMxtKhNlGGKoMCxm0WdcS
mxcH+kZzM6uqiQcm2AOuvnES0ys7VOIl20sMrDXLX65UI160o4x2d9QNR9osOAUk
KoScWHfPBBU7BOlTtftsRjqSpLv2XOdN8K+5Ru3ty5FJDwQlka0Zj4NNV5LrTEkc
emzOzDemKRuB3qrGI3QVI7dyHeWeQ5OIJl6xYUdPNMFtOI9SJfVBhy1Ucv4iQDAD
bpU8p+9vLfHHhTpynkgGivd/XNLS2CxEABDPt7CM6f/7BecDpOravzoHm+tHTt9g
ApM5wfkkWM9+B/wFh8Z5GKNWrYDdD+FL/GEyrluFgp0s3z5X8Hhq4NjxU3kkkzss
kQw4XRVuix0IedOYcPnLVgyy2xW+1f1JyTEWOkfbMo5pjPzVxuFbOoIuZEYJ05vA
CVGz0jrtZE6zqSNiAajq2uK1QktBrs+naAyKuvbnvn3T3783qpg2WP2+Q39D7zaJ
xkEQHeciYGwkxdaHHko/qM/fk4FZvwz7xkcqkmbpS20ITSIKVLfji3ZjSfC8Qbq/
IyVuca3A3qHo39oq+EgXzggNHPFKqHlup8PluSv8cwVOZlgrcg5XbEIl3+WjmRDx
wpZH+5Ya/KNOmpnf1kulLQl2XaJrNkg3H4XmABug59Mde1i0pqovagCXG1Kt92iZ
FvTGVm/nYSQreYQyKlIGS9FtkvWavvx4eTxYGncbXD8psk6q2ZRE6YfOskaTZneN
I/vNZ8N4Ej8JMXsZJC/2JHwxuO29+nHofE6LlLza2jmwlFM2xCG0qLmlgwPdV1aM
JtlPUXWRrq+WnTs4K95Xo76NEw04Lkly7wPK5KzsUvQzrRYJJMJZQxjF5tmhjkBA
uQmabwDBsM/InFR0tuYuU0rgMcAx+SYZthorxyzaYCsBtKH8NfJq30exmS3+L6Pw
zlvWaDAbN6/wQv4iv5xEQI2hy9rPPw7Oy4diiFWFKeZ3nrqdcREbDWOfCeO8q3jr
02TQxurdEfQgauKvO/5orp+g5G3mRI5q122HTugHgfiJi2Gof00jnwUlHKp4IA/p
2UcmL+GsBHeDRAc0Y2Mlq1Q8Sda+6L5V2zlBGdPHtoi37bo7gZup/xWr8U9DgTig
A6WasDxxhDDJfmMHod80uVW5Kj6Rxl7IP4otJms9cojrlNrsTROUQvoi+wM0ZBoG
bIqmosOoAyu+2O83ogZ7HYsnaehdhvNuLxBBk/ylp6E/8WyEfMLOvPfQucgGTfw0
hVBHPz9r17Ae77IrExUHhOZmUG09OXXIMnxIilYI5NquJONmIXUYPZ5ai3NO1E8g
px/5Ip+5XSHAVVjnXH64LjWbkZJjkhKGUvCAd5wUTFTFfkHVjGcB/wx6fAVRg+CJ
9y6p8qUx2ssAAS1AYNw+ZpwgI7h3o2Tq1qfWRzotRQNNIhnLUBf3hcOHT2z4QzrH
V5U2L1ZjlmOz3ADSFo6TBg6WeJn6aDOHCUMc+TpumPJ4KLXyyHMIco2mi/boK+Sa
HMT26ZXs9skZerla2kJQ0McaALV5wXolemXNttNQu92cqhTcq+de/3Zi13A2Jxwx
rY0siN9Uha3WJi2TatgGGGlRmk/qDHR0EGegQkRsGizPQFxXShtIeWSu3ti46nVN
2E1M03wFggr8is9gI3d6nvedsdqUXl6jJIzFUB1zIh4L682jERBoFSeX3kUr6bel
5dwQdqzroH24QH863458GI7ao8U3iGvgwihBLKX+Mp94ERVmyeXyIBe43hswFWYl
HcFYfM+RlQPe6O57UzfUhrUaPG99UnEif4dXyu0dCiJnYiXpzRVKMc4D3mtaEM7I
mdTXN3GgkHIQPmjyxfBlKRHAVvZZzH1vwRwZF+hjfz/6h8MqfH+JQlZV8X1Vlaxy
aNIn19SBExAbKIujqJwSMGLU982Q5Rkh20R6AlxckmSiual0bC2q3y+emDvKuZUo
LDDiLNlSrFHNogAmGEFrkMLGYP6p9FGlw2iS4nzBW1bglY/w9nOiMKX3V+iveTtJ
3aji2UOfjp98n0HfkQVZmKAa8KTgL529uEwkQhU7FDqPRTlZkrYnMjRLPFfS7uuh
2r1e+nawkBvai9LAV1SC3Rbyd9NxqejGfQI5gzD4qcZ7bf7De4t2jIpVJ2ObL50v
nsI07nMdUEv5KET8IFB8FeeQyoxxxc/zXOud1VLzGa3lOvOab5STGvMRhp5/puAj
PLlh6YaCQR8C86YkuqewKpgY+BNGYYna5BJSOdIUwWb8aDuDzpr72Vgq3S6xXMJL
YP/ypFhT5YJJFQgoTinFQGMejz9tLPHZvMnWDZ8eCEs6Ql5SOH5rqqosur2FwFpP
AnmAraIOvb6XYRqoC7eHLF2THPMMaY3t4/Kj76NG7E5NqCjK2/ncIiAtv/iMQOGg
gmkMRJOEA/RID0i/U3IHiA6JNMHAoYhBMRZxiyFG+a8ssKoF4CSqJ7AbXMwhIpXe
nlxDVaM5gnj1BwsXc1eMroCEDVkdIbLqfhyO5qoV8c67i0J4uA3rd9elNICiBROI
bxewq7RvzbHeCn3uuLlvwZ9LBqQM3fFVSnOkqq+Gzy5JsFdEADwBAMZImkAImTor
TLQ3546So1Jgvs23et7C+lPjz/wzod8ph+K2gKNXv2UaVD25PlRD1ZrQfvQt9C/O
JYKDuBIIzbzeSYQAz5mDNyigBmGxmQP+JRpK+GTzKpEWreZJzar0GkyJQ8VPqT97
cSe7RyuTeDYFy/T4hwTh2/cks5C+MP4YbwoAVS+/kplqHMWkI7AjJ40vGCe/f5+s
Z8r9i9OQ/gwqJPTO5X7XrB8G8amoTmTNGTTELHrMTtcLijQBK3fAulIdUBo5YBFR
7qWipy5VpWikQxrIofGKvKSGubz0IJV8kApigHxEv0mtmIYXtdmNjGPlwHajKw90
326yihcrvuhZ2ml5ESMlE2Hh+UxMlSGieAG8gdEkr+z/jXYvgpHo9Cs06Ccm/hrx
JLu+c9HAPMHM+OsIzYOtZhdofi+aDrIaLirBmRJl8dCLwIaUBQ/6xXXhp253KP5F
wpTaCoQeUmbOjv7KllyLsTgL2EfmFzMTElRUhKn3qDyrXwGuHvmgZvenkvk7vq42
xkvtvw2mNTLiw95NRTiv1DKHdDf7nyhv3gw/VyZv2qgR+5+EFR5cDYCas3t0hO6l
itcJVtjkYf6v0PRX+3NE2qhz0neT8vt7+sbvQI2tC/rfj3E44QdQFfZ1EQh+SIfv
FgtdYo0gAeo5RIPIk7m4xFYcERc5p92iSHKhSMT6VLEe3aYkrYRKeK0zgXSO2W7w
VCnV3zojwuKzt6WGnREJOkbL6ZKrvJmBqrh8+OcNEJzSBVd+FATHabWXkhj0iLra
0N9mi1rebkOpWFEHN5yAVB7/Rzh3k2EQ8lrXtEL7mqCFASaAgJw9hQnyvw3dfC4C
gz7vAXNVgDwCq1HyxiBeFAHUQGh+SeGoNJf3pOuRVPyqdfV0e81eZ/yIxULskNmy
uOLBbkndsaYA5lrenr02tjvtxPeXzIlGgbCe3HheEBm3tseXFAdQxpuJSALehqDJ
CUFztl6Bzm1BLiAtyKJAONZsb4024coaQe+s60rFQd7ehWAM4cKvOq+sL6vmrRTO
NfHolYCMeZk71k+YpGtoDfz9WQRc/gxxXHiI4t5R7r5bvgnqkVylKjc8z/YSXa+v
w3jK/qQOksmY8d5gBmpBAJeD371Doi48Tl86ufTZjgEgg/PXfz5Nu2c4ZMIiBYp+
z/ZG4/2FNlQkC7v6ZBpItCw+3+nsJtqlR60QTXVDvPsA1rJrkIxtdoV9kMeTlsXt
rqAJInYUHojGL1il0l+A7dZZrD4ZjIn1cJPHWyvmyG2v0kLoxrGWPFQs0anw5fxF
m5qddqXFgS380wO5nVfl7KNi4gpONg/rtKWKKSO75DgOel1re8ZBxNGBX4WVW1GS
ASFtfJ1qWXwDE2Yz1OBG8mJCn5J5g0myi1+wlxykpVz/uCXLokEB4jSpJ0zg2fbQ
vMBv5plStYYnobrcWT24Jk9CcUQlGUuQ1QHtCuoT0XOuBNON2RxERnl5+xwc0tgI
3/fzhjT2Zr673nIBSVzM/ngK/C45VRmBnf8qrqkM+/Z4/JdlyB9ayUM4fqB+Yvji
mVM2JRoSWqqcjHMXuv9ixF5qjyKhSh67sb0rh0kR9BY4aelxQACkLyyMK9Nq+f0O
Tpd0pCHVR6E1uBtkT2R4fFjR2dKWiGOSsrCwNIw5+db879dDC+CFy7Jh8TsyrQGY
Ij0tBqyAhrsojN9QLPtVDUoqtcH3SGjk8EDXmXJH1cQEY5dx/u7Lr6vcLjg7w9DF
ya5JX2YmjJ1EwYNHkhtyaaoSN3UlulkJt4Zzdh068vDlo/90/JuDPII56z8lnNNZ
/PyB8Ah2ad/WsqCOELROqnzBctC5qeDkopMkiCm9GNMExC1lUpnHW7gvVdvVTgap
TWUvfkBZktkjQZuSAcuxyc35LVK56KHkMIjgfoNDc3MrpeBKQ373sx3MyS77y+rp
tkLUMSzYFh0dbncGcODYpea01yiSu1L/ckttKUn9xM3aKsEY0ISXHo9WNps+3YZb
qK5IN6MAprSgd70BX/z00vHqrEASRvr1BjwPZ3OQ2/hcv83vwUUAUeGoR6gb50GS
IZha1vEXKL1zp113YfJZmPmJ6qnNHEMZQp1GUJUMqgjF64tISuNGVIY/zSgXtA7a
++NiuC0yldPf2ebOU798BygNgjDdAoVMz39i+TykxeEfB7UI6+fqWoc+UtizM4QY
bBq8PhosWW/PwncoO3M83DG0eveVz3BBWkyrQRBit+vsh7/pHqCFinpDZLnb/NZT
XPiAElB/ifZyFHrcvhvZSdvOJ1mgBgaZlQGNoNU0bUW73lOh56XQrlko30THJz/e
SN2TU1nyJQ/5MuYMaTi8rqMWBSfMnQWoF2o/NzVkpF0iboCD+DoxJWT3fXiraKjc
5/akkvWSRtsEsyueqPIugRSw7OfsYrGf2VKKxLo1eZuZh+XkOubIHTixN5iLOu79
+yFc4f6Bb0tJYZiWTCkHyyvfMv0JnP5uNO4eI/yahkRYG/7POzwAhIjkCKSK21Ky
0olbWzvQKGFYgP01MaitcwbxjKBJMiqMjf2XoU4O1FBu85+m67zoCqBFGIAcYrO2
GM6mwg719BBnV1vGZe2KJ2KDKRFh72BCAFHQfJPxEiYe9/8aV0rUd19TaHTf5EWR
bvuPVDUal1nP7iDDoKDSgFsNRHrpc4pGdoDMB+U8k3/6bOoj84R+iMA/GVPyl3el
Ir3Eaf1dL1MP5bs3Z2UAWfL1qUyglbImGD6HWtdxRDd8XPyaaduuo01aJ7U3/A9x
mn95Wma08XVQMwwfh6oNY3SAkagEd2DDj37XDqxvkEBlmVWsLpack3PUjqwYZNqi
kE8J3BL2gT+0a7LROs2gDEpP3IVDMyYlVCGFgbaFZOlCtxUrkheNMgssnFxnNWPz
KmLHkZ56Fd6ECzGHnUe33udHFVj2Zo5DFdDtO2Vxxj071l9sQKVVPpzS+7ktVhJ8
qDI9c4JHrM+mNl+Lvz9d7pZ8lFhV585UBJH8wFYBI7/mxVeQDpgVnLWCiJhrzpMe
fiLcQN4r39vxuH6E3sK7F9L4czQQvE7GDPYyvAk04PByUmhFp37G/KwadrfO7MvC
uOJ/WbqE1i1j4qAm18WXs8eysVBhQUaRrzRjgrRzL3Jw1j9sTsaKXQtJUXtufY2A
gzMP2CECTVhUlqnYDC+HJ5PxZwtDZHSpb5sgAztsHG9BRyxxfAYblbjKfxGIpNmC
jPEZXK1uUYlso2RT0I+AguXdt+jhbUsGU687QL8vbmuGBif3YBB/ZMmoEEd1TwaR
wqNXsCwqObfwSRS8fJpGfdrsMqAnbZYmMj16IQLqN6Gv9BzKw1QV1rLCw+tn62WV
CM6aTTrVdLJmCdBApxBnHEaxz7VUbj7eTGOVCELhjFl+EwND905fZ7A8zeF1YR7i
KFJ2is+wKmHKDKBlma5+RC3YOZQcqlpPDmCed8IpHy0Z6+8mmr2dYruZmWoz4EyA
TxtYFzKYABLg3woknDgZdcFtM6i9bfi9UU+cTriNoTkDTuX7kiuDiXpspSJx9llC
bwnJIuOxK6bJolOqwzBTQYuZSPNS4uy9ObO/gcAZLk+PQypgYHeiz7IRVM4GHYHT
EAIv+tUYwRwZ/orNHg/YOjhIwQiiBTrdxYlWVy922OIiRjHgEyLTKSQlEOxPjOrX
8+KHwKNGAL+bm6PFRMY4RL/UmAIgi+ox0dJytwqzHXnrD/N/6lKjU/RroZRThZ+u
nAqBcsqkKOjgwl7nCDa18xrCNx5H86tHEPXDIWdsu81IYaNuiMzCSZtcOqBYukUt
EgF4A7FH1sjxAnvO9/w2t5QrleN9Z+pLRwqdixwG5FKfq0YKJ0BHw3QgFu/GMC0o
WXIoOiSrTMUTEENoQOxL6kBQ3lKAQ5FgJ6TPGYcRVNk0JdThQjdjweM3Kohy7DOL
WdipBvmb5Anvo9bO9XbEZU2CxIx8fche/EH1lnwruUgF1X/ABSzS6c9mPQ4v8mPp
ZlgNhhr55fVa5XeAM+Wcm4x1FHf1r35eedj3YdwLu/blWTL4tG/1D8jew2G3X/vL
N5BPpAduveW2AW8+kAE+rJWUQVDCYGnXzWYNWtM7VQNVYWo2ffUhcqcNPhf9jpgD
ffCMFePrDm+Jw85nK+ijjYcq/vDH8Jr9L5sEyFiqZew4EyXOcMLT7mZnY8qNrG9T
mchpecHjUPZOl50+f3ZSOZ6f1czUQ9CLAANujWsS7ed6BPyTfk7iQ3xY9QubSm3A
+Hh44v8lgrqqUfQ7BYzDZwcpLZBp66AkEueCVHE4/qDoImQWAfgr1yaWvxE3GKYW
4YWo5L9rTJEJJ998aAoukYtlDeSOygvXjHx+8ry2ilflj1OVa5M5ENpAGkaqeQEy
tHSTWsCgiGfRPOtqecp/10UqzJP/GTV+YkkooiGt4oVt6heNf7dKb1iQ/l5LHxpM
9ad6BkxoBafUSOkuUei2dSHfKAkN+hJbgJV7F1V0kfwkVU0lYGxycTZ9EHidku2u
21L2y6xu+J05gd0Y0KDXMnyiUKIbMQ4Am1WDwY7PAjdrV8xdfZP/qFcqcdAD68fu
9YXWHq4BXjuJFvQjsOf2K/wcq5K11IHHSxSllrfwiTCg6BsEKx9behbjnk78XaV0
qDghcUDrZOA7TSiUywvIyU8zafk4cQhKRjrupyZQKissUe20odVADDi6WAs7LIkj
oVB9TiMBc5H1Bx/AhRytRtGRA/qW6j53CMgMQA+mhgZv5CVrkkbvoXm53QDAWZ+F
B24QOU/9r/RCB0oFB8K6ltdln2kizqxI5fB8MAFfyEq41I53VfOqRVFg29vPkqGi
REyBVdfWcZNthNJRqEFki7nIkWHb3nJ688xN1GfQ2d6uFfsp4JV8aTWH0xXFSMi7
2Pe0iIhZy++/kR0+KGRPkCDGuyy+udMXDeXRwUEo4IQFKBHL24T66rG5+KsZsJQ7
WHzgcPcPlXYPyI/4lwefXcykj+0o2ML7JnDeCiuNkWs0ib66QoP5IN1JpV2JWPBn
/zvB/Dggnt52y0fIgEk82HPQdZjgtCvqQyliVqmxty+vekjO3Ts0Olsz9xQGi/OO
1bHAQb5M/MY4xTRhhKXuVB1iz/Vig6e1N9CoEBXHw32KWqP1xDGVZwKEZ8hxCaWi
ntW5vjvFUpS+VD9B7D6SaWLX2gyHKAKPJ1Mi3mig3EVhtPkiXIRB/AMAWLDtvNT4
GqQRE7kPGGBXniGEFht2wTQjvMZLmOeIX/8q/Cmkeejw9o1eUARmrvA07S31ZOlA
JARzRF6d/6kGvx1nvKloYoOu1cTaE6HUari51BqxZErldxxUKq6I4rmo7tKPAy0R
4xeZGM2LKVLewIIj7EGHwLJmREYkld5oyPbeDfxQ2RXD9AnQqUTzd5RoFtWG9ILM
5eNPRCvEwlOSWM9LCeMRD1kN5PWUgLVXb0m0vbJ1f1z70pDIAhYtM8FxAUp1l2Nj
M0HMil8gs+NWBVI9bZPD3kdtQGrWzt8U0dqHVp4F87F8kaW/ApU1kno8jOwr3mPb
vIVdZOyNf8XuBPAimxBy5T/4/3mxxHNDp7IpviZxfFe59Q2Ttg73GDYaZOHbZrdC
kzXlifBrf4Z7WHNnz5ojpCJYJtw5i093+rt+rN/kW2Zhlv0Lex7fwRrrcakFO5Hr
YvG9uyLMDTvkBvGu1tAqOzCl6m7nna7ytYaS8s4R+1172LoYCJEvSBQ9pTjqPysq
H7dMBr42+fqqg9SM4rqjKEQmdsvY4EtcMNowU7XiOqp82V/oXpQc8zPjt7+xUjMe
RwaucP38P2w7G2PyL+XSVO1eUZtEi1rp7yzdFaAvnwD+ah27ADX1mEFi4NSQ3IcW
ae8S/LYP/s5tTIS9/YzMC54gIAcROXCj2ytUrbOL3k85dEjrVpB8LYswccJ8js1H
UaklBJeFKfDc3/1UStcqrp6bKVeHeF6c6R+Si74kFIBX0oTxugfl2lG0N6LzfXhU
tSb03AsxkkeZr4q4sly6ak6RVfHCqpzntTAqjfjvPecgRTQdf+qpsa6YaaC9kDFN
d6QAlgN30xLZZJlXGX4smLey44NYYa8xoRoSJsFuTBWDnUCLQ1OgT0ZdIwI+7cwn
IQJZzd5FFEAuOBRvAWGNScDvgcMW+NrJcuWy+t+qtFxoqrGZiSwVOBi+1RzV/Kk6
oW0dU96b9GUBsLT9NInyOB8Pdhpo6jzl2S+Mp0fFOIxg+LCsZD15ZA99Ba7Qbqx1
9/Oxd8Nx/hN5CHp84ilUF0Nna9n6mu1YDspbl7gii8A+E+FeoGr6ZXykMLTx4O2k
rfrhvIRblYUHkwZjIxgFCkw8GDBG0dXZPONzbleG9wyLU2OFmDA9qLPxz1LvVs7i
LafvF26cYzaQPeQh5LThKqDdUM9Ft48caHHyPylr5YuTgAQWhVRwBkUIUBPpc0Ip
WG0stI950SxKGXcUJtkXDvysX5e3hdwc2L/4IURplJ6iyRsuJ5Q2KJia9QKyXGFn
Str7aWOWaFNBATqaoK0KNZ3DO/Lmx81ERP+VFqh601leHw3+QwD6mgmrUnq6M7ce
Oihkh27UCgDeKHF+9YBHFBbsa9ouZ/04BhorL9XvQMPCduTGgBW9nX+q0PSZSJk2
sbX1Xvo9kY+7KTSFAuWx40hfVju13QPX9T8eLIC8Vn9tNosBTOvwmRv2DfUSOj/6
WXZdWf+mXKHCSoWJSvI2F3Pn89IZhZZnH0N3Q//LLWp6Jd5XU+N5ZxScXQ79oNIZ
41hcuama2dNWgKhwEjpUlSZw9gVw1/CxX46PXzdAicqfdqV648ZEIjkRXaUkzhP6
//w3pBcizJatbo+nHRPN8i9LiE1cypH8T1IQX4+SVPgTmceeXRupCOfe2nlnBnQp
fxpcFkcD8tDcImr1mbCJtW+K3dW9lrlT2t3gxv/4XXwKErqbhhMyVVNNqNll2BBy
P9YQrZ96dvOpgocRBNT05mXtjNnZHD0bKgNqBCcMIZbI+fkq4QnVueJbn0GKAltp
+IyGNg0TS3fl3KN/AGR6drogyOVQVyziojZJ9q2tdTfzcGCKeJ67zsgQeB1iRKWV
jqxErZF/Ga6jxVj3a60U/164ECERINJTOjsFfJodkjSoTFKSKfHMa9my+mHg0PTM
5QhjYgr501DtViV9ROwttib0OhVCndleO7YGkeQnhFnwkC6lRaanHXI5+Bsn6mlx
xVsZgXFQ5lqoFQSlwys9Gr1xqHIUXwo1eCGBa1FtAYvGRjIXzbTEzAYkjZuNk4uw
qMY0bIfLg9dL8XK0gE8D7v68LigeK+a/iH9QxYCpGsqIMrvQigYRJEQ+GioyLZne
Q/oGU1pcbju9T7SNxXBJILe/wu837S2GjJfrm6+X3jV685G0NWlK1QfWzksYiX1c
CiD8IWrC/GbsdArj7/W2TeX5g8WWK5Jg0gJjn+WzNHPs5J+fQwP63aDK3Ha51t0u
EpoxbwfC9cOX79GDrnAoKHWRWXfmXg0G2Nq/dm2e1mB1q7TMlaXhAeNdXKiI60bf
cSF90LD7ceatiK/1d5N1G21qEd+yM0sGE6atdVggjSwkvd0e+kuMEJ57miZZ38jM
g6TgBghT8iO5iDYl900fxpcu3UzAjTQnoN4CqWT+K7KgOefd/HHJSkjhnZZKFnVL
yeS8OEras6kK9tHOjzbNfQDkYTvQxQ4UqnxiDpB1QYjM2adv/WmsCRw5cqx8W+El
ndAwSM857TyJziV/UacWdbeUfP1wCvVpHjZ/AJDxjqJzFZejzx8Aa8poaxEv2h2A
PbE+h7BAfFdj7z9Iy2SUorn2aML7q++LLiWXZtJWH5kwx2TMkLzxXgJ3qFAzx0qu
y63JFySsyDWoD/9ISSNBROyAvcFYlPl4etUrW4mZPAb0PEbTm4SheppQxJQaazJm
zhOSAOPETL4viJSWqyG5TEKlep3fSm/t/thGL68opFwpSVT2jjkrI7NZmhEzasuQ
JkRH5ECFw/DWhn5m00fQV/CBwH6zumkzqyyanl+8eAC83yvT6Jyax4IwHe42KvBV
8XzwzI9am+KFLszKoGtz/ELcaQmMa2NrN1e2mqu8Ap+ujj6Qg4i7yrG5VY5v91lH
hlgNmyjExVw2S1doUeQAk+4d2s9cCROTItDDaMnG6NnOiLkPPAKaGzkT1FNhaC5f
Tpc00Cs6pYpZ+HTYDGZvRHsZNcYC70k00tb9BCwvxdAJK/Jfi3DEw07vKW8+2g6V
MH4r5YTOoa9w4hjJX7jg4vSMRfhe/uSltvh2Az0ulZG+eI6seieGSmEL6oWp01NI
NV00Pk+rkm6h8zs9c4MniO6FwsOBwjjAxgOkD/88pUUorxyX05nrOM5gDP+Id/oe
V4xXyLhw799lT2YhYndCZcIHRsmcoP1KbgcO5UWod40CDIK4w6isnJ2ls/o5VBkR
6vtRghXMndGKNaZuT6h9T+W43emfAFxYx56fO1CpZM9DH8vRHDPzKJLU/ogn1PQB
R46zb7Wjcg1tODeJSHNMA7LZ3RDvhN5NTWtAwz+w3+kiM5ynj90d+Sy5Zka6BjTV
4f76m3USuwUXBFtgskWZ/NvlmH1WND+N8KiEfmwYbqZ8aw5qPSlpMh4rGg59H/kB
RGhMdcz7qiKonlE8qqg9cfiuLDi8O2mu/GUSA9zvOhrUOUlQkCK3ZgxKcOTX5QRJ
iuc4Oj2eJick3zQp5d5yQdnzcGxNsL5+DUdRB3v3Gwd2pfxFezOnjEhELjTp0YW0
qHqJtuS/PcE5UFvz2uwcWfUq0ePyvNGIiC4mSb+e5pcPmROunCIwxsfUnWTc53gp
wY0SmqMBOBczO1tWsMnO9UPMQZ8tMS52e219C5/6+IUaakb+iaxePa8ASy1PabWV
Zoh+9kWa+x7SNIt1DM0xNy3sMBcWCOC1ll0G62ZPcM5ZdjkHHgBdYleIc8T2YbOK
mFT++ew7cyqfSQz9NijIUdhmHvAhzfEFmLUS1dgVp0233/qoY0suixjN0t+JVKR1
Srwqtn+DUxsb2kORfk44sLSMsA10yC5Bj2WC5+dcZEELAMovPoCykPD8K8mZj6+y
to+fVyMkPJQ9+LnX+yzXkVSDyiz3b/9qvI8G6dv1+dx7WAwWRe17xxVQnMOhOJ8/
LURUgwGI3SXkmmbxn0nFH1Ln6IYCkFO+6BCC4yxhltjeQSks88pG5gxMIVrmlAB2
Zd/+h8zbj1zq7y0subQP0o8E5E7u1NJcSnOSE1m01JJm5nWz6OB/5L1bvN38CtcJ
elO8Vkt/2QgVT0b8ewsq4GN3utX5lKUUztnO90U4y0Nwhfn7xWXYy/S0pQ9xEWdP
gVXzFeMpUW1XLrqYWL02fP1yJmjIf/kI+6pgWF1AK3P99B7Q1X2M5ZBtzKrSY4Au
Lgfb/G+8DyNBFHh8rWP4J8hGkEyfMwd9IyU266g9bYU2agJWKZ8gUPZCaEKfl/S3
TQYNFUFB6fbMETM1WSwqbidscaM6st+jIn3BwVH2M+4WITGPdqx171nKddWLCcrk
BfxXdmu7niNTzgUHUjoACWDv0UiZNmBmWziAF0yRvbCo0556RW+Wszm0UFlKkbfJ
NQh6RIvlbdNZIvgBzVJ7mSuZCtDewoj5OxfGZU1ti5ikBCXXJ0x+/ExbyzZUB7+7
Z2IHib9EBDeTrXJmCz63Cu8IxmLqiQRxfvgHrSNOLiWck7eAhJnimGbnWP7cmYhX
XijPlzLB88KW4Yj3V5aslK+NH5jgrrbeJV7v8Yr0Ev0KXUGffdnpESr54pcfA6AA
4v8+QcE/7jGzwKrlAM7EYJIyqLNPHd0mmIRJaIzh6fNbZ8Xu0ljDRfq/Oph3/o3p
EAAI9RdFdguQ+gEPl49oCoR8n7iN7QZfSjp13wJARyHksqarEFQHeZdGiodcAYtc
DUFRwE6xyDHgRhPFyTNb1GzraNVaSGO3nmLLlpkOvkLP74lCJOgmhqnGfVwAmbvQ
yb5i4KS8Rlws3vmg/ODm4+cvf3IQUK3/EkWdhr0UjIVULLeWTryEGd4mOsjYxLJ7
+4MylB/4CY6XVxuQo7xB/cS5ccB0UCDxvTu+rcNX2RxUR8nZkH7lCXHHO88nR0R+
vdPaXnS1oORDI2+hV+5itK0KV/axANSPvy+ZicMC4gp5s0jg4ciBBG6cUCydrY2A
agaD1bre0FOr6xmZRTP0+mhHUJEf0gojHgMlBSsOSgABFBgHl/l6qkrdcvLElIJ6
VNSyUynCP6XZZEWOqOYIsKR4I2Yc88BDyab6j7h7iDpVFzc3ljPLmpMc53s7awvL
BOtoLBgz3gtI0fRjVBomyUx2ztPEb8dLva/Wdx+vuvUEflUiIsUmvtArwj10p38Q
5NbgcCGnDxVjoSjVykH66Dz2XP+HY8PzNZnijgwQPMtZF4e67UXRfg/iejZV0TbO
vFvGRd38PxEWN5JkW9vACqXGW9o4P8dwJ2tl5Prjs2PZn5inOe1Tsnoxmj1KWZT9
PiFt1z3i0U+EYGSu83FNIKYSHxuCVl0r//I724lsGwyyzikoEdlkPw0X6UmzsxBa
xI1ft3OoVcoaQ1mNiXBQTXz1OzO+RGRQ2dJNaZasUVz8W1cLfrStzKQmarmM9qI4
FU/QIXnE9IE8am6sCgYR5JJkPRdkSkwX2jgJ7h+G95li+yzLnss5h+7g8iMlQAJ8
fvMBO/caxeV6tKx+/nTmVSlokwDx5sO1FmPwO89hwvWicDkV3PgepkrFa2IoRIZd
sAUVzp56x3Dj6cBQYMlbvUe2N7xnhLDIFQ6wLEm7OvZneEWClp2Sy0KaVxV7Of5r
b3NLFhfZtEtruTsMBuhc27EilieW4ZICtJC76hqIFwA5b113YRcgxC8kFBUNoC4w
qNhaPwrtxyh7N6wZwAHWebaeAWMTN4wZoGzLsGhQzqiWH3k8WfjQPAV4aJ7uf1T/
hA+ijNyN/GK6D4bmHcgD4Dag+JxW+KU4LezBd5d9KWqyQxpQVtflFzGGFFdPolu9
Oa7UCunSDoU/ePRKXhi3sZDjaAvTPt+EGrWiWBJQdJAyJbONylwlLZcMPIGKtLn5
Vo6PehRwXHFCECVLpuRGklDAkOkwiqLN26/eg7SFpOT4tl9nZtjKxJ6c6Av0pa8x
cn6+HYW7MHhxoOPVat+MbavkABGFoi8gSRtkc89qX4TysZOXwKzfJitBwkILtZxb
DjbngKxayYTFS0PWtmwubuG/cR837PRK7nyVsrGxrBK471owIbhZOhqs+XzIhUI2
7XUDMXvL8thDHvIuUdeNjuD9Mew+x3l2l1AFWvj6HSHaAL1Ke+nFNYpa2sazMcZl
bndazif1XClHhH51WHTW87Te1pEAOaa2Pth1z+7Wo0E5zV1yynR4u8anN2GSsfO0
e8FSukt8LesiSvA7xcbcR7YKBy1/sStAbnhCkvaYcRZXfInx+4wKVuDUygzoKm+7
022pkbtXVpozdvB9zZTV569um3wTQHJAOqwfqfGeNkhbR3XDwk+xIqFHpoUvAIdj
jMLJerm1oCa4h6NY/Lt7p6fZKus023uvXEVsboNzD3R2OdmIzS+89YfWqm9kN46n
20l7LxkeIcUlHwhsb/S0H8ZOrAJbsHtc2spR8hwoe89ZRgs8U1PQ+3W2y4txtdRA
cTOQBmZGmTyM3QO1ZVqJW4o/i2MZcJO3H28HLtMueBGez+9F7IpUTChx8STYdRut
j3GYQp/tbmlMUV1JuGFBdPIt3o1bcmO98xg+zyF5pjHNHLT6D1FWO4tKxv1TFpiV
FhicaBFkALMkmfufAjPRK5q39tutoyE9arPeNwnERCarR1KNBOkl3kiAzJaMv26E
2MVAF6Y3w1436MSTbX9eOFaHqQxDRvL0CApdB+sI0lReti5if3goPO910EBgISqb
heoBSoK6q2ULEhaMKqrRHdwjZRNjKjM3VYSbogJ8ImANB9S0Zf/dmK6IksY/Jz8N
JbOF56JxWwETD3lWb9/wrbCLYOlYwMbkH2D7E9gtJ4Orz1Qo5mZGGbaOZvVX8wq2
tFCQ8FjhE6Z67PmlhnHxu+aXYop1mFno/qOj58rmX/+qJ22HMypCiC3a+L3NSNkr
0NFl7rrsB6HscYZkK9EAgILoH9eIIix9VutCv6lAt4Yj9e35B6pFR19m+NHiGLlX
YJcLCy5j1O/iiao4OqvlVhsh9c+qPalmyz6RKlwgzwfzJliR50YT2/YnZzLesr8f
i9UDnUq3XvgOiPLaHlUOEaC7+I9gk40ZE/cjzRZV17RZHRKVMJXpUQ+/47YR2j13
+A0oPrnwljxea3GmGimBUrjz14zRrU9mFpTI0yapE3oquH0gYqBXUABGGhpueoIo
MkZdyLjC0StxAcwB+zYlZF5QM+m30TW+O80TJ4Yg9KPKzRYHcr3RfS5saIt+IyZU
vK8g36w3GbdlvZxgHZGuNjw56tV5ZNWwvnEq1GQRYRwpbTrA9OQLHxCn+DAkd/Jr
f1QKar456hlZ/yrUkggLAQvchVc/9gUo33Wq9BRX6B/ZxwuUk6/O2RcpGMWf1QE/
Cty8Dc0gbjVAuTmOCP9fFu+Sl9JZ4ODC2H9F3ZIpnC+cTJWggebLPCU4td25LVKd
DG2/p9sw9nkcXTajuJ2OiXtte0Gphb+DalGyR4/xxEkyuFqX9giyppWGMuQupxeb
2fq7T9Ql8T6GFTctf0Gut3abBu+RUFuLlTrEP0fMo4hfOqjsVs2FiPK4ssWMvX+f
bThELqqpDQnTk3MW48nb3SYRmLkmtmDUbV7XAXER7m68ZbFp4NpIgkYnVBr1Ht3+
276qyEN7HfETWmVOH8F1KyuYtceYaOcrsbIQNTXUIF1HtnVjb4fqLOcya4UXDfDh
VDJ/su6/doI69jwWCtMb8dIgp01AsKT7Kr8b9E9i3RtqnZIz8+yDSSUzO+Iwx2e/
4mPafzN345JH5NS1qo4V62GyjdfaV/qTAQnjJYeZo5ddLQx8YevLT4nQYRayciWA
JhHyKkXsuF1IsxyQIlvs/hRGtVLV3o8oSdjZfyebYfLwb7UAjFKR/E5MOIhKLAWC
AqkOqWusF/wbIV+EHttIU1LjeFmT2Oj6mGAuutSeovEMR779DWaBTy+hvVWRDsdb
12xpurYbaDOn96j855eTfNP82FmATFe+U8mjUpPT+Idqpt9ylCJrII5nIu+fB59y
oeAtjz61GGA6G2bz3+6WxIg336Cd96GGOB8ypazgbYPPtRnm87C7qypLcgiuKhob
Qul2b8ri2i70ZGCC+z2nHmZOTU9DS/torcPzqrHh0CtNwI9cLmXDE4DEoWG4H5yw
NqyY4qBoSZXxa0330h9lJMUprA5FiD3OnA1LeXgAwaixTIihmDBqdgYgeK4Dwg5s
hgd8R+ieNN9ioVYdde/Ya2dLYDJuIUES6pLH/CYKU4QcbC2OXY1VjQFjPBmCMQwA
sB3qQQzMwzRTrMa/5XCOfMb1nnYzDyyS12qSSEn0njaNf9dzd/EXAKMNX3aVCa9U
ung4a4DJ6GDdmHPNAjIGsbXXLFJGduAaIjWMlRHWBV6R/oiH1SI0OgJbtQrBxTxE
ukLmE6rP+COGcYcmW7TnNHTIDRA7laykOHysIlJdb+gX1oBBIuQoetv02+X2VQSa
1KdOEP5ZxcRoqI1mSQ0mm/LzQJIQtrU77kO7bi+MpmyOAEgml9pcf4va5IkHeUWn
XQyasPBIDUt5QQb9ZzGgC0OZ+KNiKxS3EzB0pPDsfNvUqDEI7ZVbtjBISUHLXg9z
+mo1vVbGcKxmTsqtZFz420VXqEBynLI1updjgPcZhu5+53jIFGlspYJuHlpTAchq
DN0IYhvzBss+EhAcr4WT6GbG40UvyZNTK9OIJDYRFTSXyZRGkJM9i25fAUpKMz4J
FZcPPhOqXcUl/In8hYuldMwSP7itFoq9g+17A+iWv3eGkwTdL8SUaHQUwsm8NIKx
sxpC5eBzybDPMID+gV4mgWNERIz4ien3oo1ZmGXP4hHwfKvMk3Obvh9yhzqG9VVS
A+0aoPx0Qa+WoRb+21NgXQTzgd6n3cL100DQyWhZ1X0Un2Cz0lX2EupIDaLAO/vO
F3v9WSGkOM4my3TLh8XCKOq5aVFoCLHOs//JI0hq3aPzruT4GQ5Z1Y0SrfSFS9G2
JMt5toubsWKCIiOHSqcIpaAQeiIYLSuk5z0N4gD2nimpPVztfjkzc8NNTTymxAmp
kvLGTJJxn08l7c3cdiu7YTj1EzV/PDRSuIfNN7qQi7xr//bt7N/vPbd59lzCo9sd
CZ0Q+GkKfjL1WQC7o6hNJSbSf4xFxjUFkPE4J6DjYe2DCkyLuxLWOWe+Mrwx2D10
9YjhqW4dJOVqQ4DAztZwAPHCiG0BuHC5TFDr4L3UEsC34UgMAdpYz3TQE+pNm8tO
JDo8dJ7AbxIhPWg9vNH7mHa4DR0bpqhK8RT+OiuUSYafHqyI5jC42I8+rPhBS4oo
DOZZHRzFUqlrX7idITxF/4qq04jndf/imhgvDDgNv/JzaKMTIeFdV35JEfZPYADR
uQEgR04cD+qIibhiYSZPI7VEytUNoqlYHe/AvpLgacc88Dkfurx69pRvp56Z8uFA
jX7b9C8qRzw2Wjtdf/2VCOoIq/w4mtp0VM7jb5k7538lp7hMJmhpwfGmw8Tw9br8
odD+O7eqgNNUez1vL4FySwQ0kQjB5Hvv0sWKjhfymwRkM9/9FT+HjKNCGwFe2qvs
TO+j0E3WQoOaVbr15pZymc8UPyB7PVDVg35AUZR/Vspgx5+UEvB/e61dSCqS2gTC
Ji37Q+pgYo8Gw4pxjB+G1DKzuyB2wLHO45y7EScK0r078Od6WazKLGSuK4Qsj4KH
TZTRJBlEOpejJKQ9BVWSYTYgtBnhYfEp5fMsYZLNxduhnLe7YcwZ91ra1x0A2YZv
ZG6lLLTPArtWdqFeHz6h80KUcNvqdR02Xs0XWPWIIzCErhjqa96WCfuceWJQ/fUw
KioXxvLWMG8sbGx+8m3/yF8ZzbNCtSvnTjW0PPVc/PWYgI/IIqRutHkaYDPCJdtQ
tdTd04V0faD9IsF4M9ivcNze2kmYRKkw3Hzd9NwhuWJJtwyWntQhTjYv+41b0F9C
igYYLgBWYxKM7a23+fkz68lwhWFmXed94c5gApD2V0g0u1Y4vu+HqoE0PhiGQYbr
9FReRdPUU7LYwRYfI1udiFMdQv5V0TGeTimffCnIP3/27Wpq3zB2JD/Bs3MvXaDq
Yk+uq8Z/uSVH6Ec3xVe/lqsZO8MfMozxB6kRWYVLveJX+4VNcdjzDoAu5SzRvXmR
t81yKLFrnNffiIe1pGUp5Fx8U44g0WYBDMe1Beq+LgBic3Js947l62VwoUEXqtmW
twV2cFTBpKb6NM68itRqP3tVV/L8CVFmN/+4hKgXvZWPepRXbnFW7VHrJ7sUzAui
4YIjJBf0sHpP/0HQLbBcKa4rpdAlIePSWnDIvPLvkJrqzEYjas1fMruSBbDjQb8T
+J7F7EaDOe3UNigIVJlPxJzsvCp3uz4e7vgbnKNi6JVPwuK4Mj3D6IW2Wa9LqgU1
8481BQo+LKmb7xiswzGciXNKewR3qi/7nyI68nhi+QOn8SgjmcGhbeIJmnpXXqWv
QJ4sTwvAJr02Mk5AENX3/zHVSsiN+yXdmAh+T8xt4xOy9pphieAMqUN3JjAiEd15
BeFggqF8mqvYsLJOW6omlY57T3ZZJ6Mj/3X3U58cBAhVEyVBQ1si6cIxyeLt5pvz
sd110x97SQi97cQ3meoZLLUvctJvofNV3msJd1VqEYB+2CKZbUHarFjqy4acnm2V
91sqMC1dvgznUc5TwH9sGERbVFgsuFY614OMWCZ8QEkLvdo9LqkfDODOPzXRQZ6I
H5YLmizHULxuD7NwvQh3Ig+T4ItpmuooVPnt7/v6dC6Ivw23rBYNvgrRw8e+miln
rVDOCMaU9gYMDjWa3BVtvUPuNC0Gd/wMpTD5lewTqvqN7O5krDVZ5YSIGWX3sgEm
TROZOFU5tVvegSfpIEQ4W0VXlb1z77fnq1ZleMPmMKUjhYApw/rr32HoMiF/AvbK
Phcm99BKSR+fiyaGRrmNT7ed9t+TrxfjAS84ditbPIKu0SM8cxnweLckXxCtQHtW
/DGFEx1f7Xv+Rd+JdQ4u06ym6xq2HfpiRz2N1/dv44iXI+Ue3r9bS+xRlwJ0/LBD
iK4o/v1U9p7hvq1icrP8c3MEzPxiy1zZ17NNAiE8OXtaT9E1MSD9/id/tvx4MmHq
dN2VjRskeP89iUP8b9bT8hVdYCkme4PY2RCdQkzucnBYKOuDXLt323EF7JB34EyE
/xnGoZ7YpWLxRYYIY/vyPLkB+jSZ0ZeQx03djWDJO3LPhLp5fsUf9bg/xu/HACdA
a30GyfEqk23Z38Mt0H+um6U+c6MChQrnbUbL/dqfX8xlr5AUY/aYz4w8dqMeLi78
Dho9DBM0DKSxtAviPoiKrfCnhKP4o90HC97EcYae/jLubqFtUq2NKmQEDExZsXRI
gVT9KkWT4EdPxLnUjbFUn8lRmSqYi4XUJp81rRPrbVOyWjS0QVX1yqmvNalZ+vCc
nhH+bX2NYVS8BeNnHiW3KvV01g3E6gQAvGkbbuX8rSHxkTjZAuYpy08osPWZHWUP
1PHYqk2I9halJsKvuT/PvZHOnVyeUg1tfacsuySEFM1WtkYKfmdqR73cFpiA8u2O
kwH3etFX8ablpYiRZ0jrnJLrb7baYEnNA/MjjtcoY/fCOI7GPUSbvQoWakdkthPB
4O+KtUTJpXj7PA5tOG5OUk+Qr2Vvfc/8Jg0SYJF90amfp/hMH1I7vClg5IV2CHH8
H8wt1dbBkry/vEO7p6XmM2SLdI9PK31ASxrptmSgUJNLvrTpw4Rks430ZMhohV+7
PaeFflxPvpdXTLzK7Yyh0AKBGWqM7WTvwYwiYNWhT3dnM9rkU0+LXwDp3XZoNvdg
AEcwoDers7Z3rmJjnWH8VD3JxHYJbwd6IPr+S3VY7MvvkG1cdIQ0ltMVVIi07I1d
ad4m8bAmc0a2OMyCvnKoakEAfrB/OgHAYyE9LLGtje1z+KomtLzISEvduo/NSI9M
sCsR6O8TzH3SYZaYdbfZitzI+C4PJbPFqmZqIPstaF8ooNh+eyUCSorAP3EzBMHI
SSzSbALAAg6aowy1JpiOBS/idGv++VKlCpvWMtWKvxlm8fWY6vOK15I+5UUOG+rb
sUiTLeoYdrwZHBhll0lwvIp2SQVvIYGYD4OUO0xHEbuNWDNAgvzShcxQTAso7hjm
51FQ4suYNv0bnm+AGBS0oDpUh7ybzvgPdNuS8EJwjHBBcC3F4KKuxPdFgCvK13lV
GvaKGLTb8PPGSOr+42XCXXI5lNjqP6e35UdksVhaeGuiWVxyUF9DGy9A0hutFOEJ
zOCWkkZoM1rxeb2w11etn88mlBf6S69G8zZ1NCzeemcK9iFaQBBNOWpBxiTctEi8
byE9AivM5/53vXe8S5Aee9CmuJ87VYjaPIfNnJLuOFtkoMY4WnETYLfzpkCQeN9W
dhPs5456vi9oal8KGOIe1CSY5nK/FWgKZK1C1j2wnCQygY2WSEv548Wc5SLiBlWx
OVvieyB0+ty0CmAvmQRsbhc+x2zWNFeYb18TKj/Ev5J2SDcWnsQszgpl2EBnn8i9
O9SKObwM+b8DVr/3sYrKHJJCHMnDCFRM2kskKTPZuD1GgxaYbeCJgVi+zFiTukQQ
SkXBk3PlgirfprZeqTpd6mXShBAu9QNgoO+Yb+y+mRWiONoQZs301Y2noIYwkCUV
iLFAQHgxxHB0qYc6BOzfjGqO6iayrPljSviDdNbOH80DM0aqV0yiLcRObK3LydPr
8kfq8qrhjI7VR8tpFQhctboRpZkau43my61KRGWTKG2Rd4Mcn5PtH1OU8VyKMOyp
KvMoIATcBih8UbcsjJiRChcZd9DIhziCn+iu7CRUlpsTPvxSmCf+804xxZBi7dJn
+9/9VaMYf+myO9vX6AszMelt7lsICJbhY+u71sqzEEtOOwyvM+k+Kw8cyXx+VAwc
6ZTlAbpiSuR44KcXv6WB95jMqeArSIESz2/HZsvTH7qFObVO4Sc6NRNMZjefjjM7
iwyXCltAfyjmDrZpd6bdSci5nZdnhkpLFWfx2TV36KXYGjwBtAsVXhVKK9d8dnbM
zx1nhB0FKtUBul/B4vugaoRXgUtKv1SMi/lEIic3WW2ft1LsWgErtQ3XwNwhjEhx
NGdmjT2nBCe5b+4rh7OL73GId4cDDBaCfkibO7gHEYYpyVeqswa9kxOgc5F3iDxE
Q6NWK8ILxxCxHLNXsBBB0rPYtenE5bKSS/PNCSB32M4Sno8mA+di8mViqRBuk84P
AVhd00Ezy2Ndx/L2boWTdegs5SBqQqcOhn2HjUvrgL23QMMUYej29vme6QCbmXJV
FTSmIfMe+LgrFdrn8uTPlBffccoxsbUCsLjtVIg7q2S8UzO24HX+55XIBklJRB8S
pBkjHxSV/mjfHjQqw8vO4kNDN5MeWK3BiJsp99jt6gadej23Kj9QkB0gWkhU6Lau
1syOWvtgg2xx7+B+RWc1OLxpbtvZpKytyQp7Ex9G0jc8pwNu4rq2o+uL20MA1sfS
98tDRnrDThaIu4LudWv+rb/offdlc+ICaVdMPGWCkIwNMV9QMb6xdc16viSBTKFd
X0zNgFSqDkqnPGJGlMFXiYUo3kM+qr7HpH2lKsk8sWmpftIBt4qD/RAENHr6+fIw
Y0B8O3LCGC2hilck8pB3pwhu3ioo9HAgCWClp6EvIu/khrcQi2JFZO2YdWyBKLoA
XM57kh4fndlMlpP6ipaqtnWHH68fSzr2MRGfnV6aHDlOMHD8UQRfqpydxZOWk1V2
IZWt86MEK2cf1Mj4e5CqKHdRVN87LHkOpXq+syc66CyUj4DfQ0PILXY7nOnPITvb
Fbr5B8AlidVS3DlAJdr3nEzmVuFFVtx4PA4cst7bpWP6qQ9OZ43xQ7Yr3Oe6HjFO
8/TuAM4GjvYU9VShQ7TPym+pEGAwSt6DZotNIr6tM+5LgbTqxTEO6P/P6VrDBFEH
oz0kxiRsAnpNDOvMdq1SBJ+owb/rjYpexTyE60F+KGYDf6YT9ystXh/8PW8OAUNM
2S3vKOGOSwo3o0oRbrXtV6vmurkCPerhSMIiCTr6NTPWjJet+QbaIkSp6O9HQSSH
Alsla3WFSaBhhplgpo832Ew8F9TzcQvSELGas8BhnKiHkdfJgij4r0dCmsJ1jZXI
tl74XXGBVfh1to9zhSnvGmRi6eiPtisVC0wUKB7l0V0O33MlgBGvWo7hEIsXVa4F
dIjsZ05BCc+Par50Fwv1EWTDlaAaf6bIdks6oV/mPjuwIAtKPybbO74ieR6NrTEy
5CT9Ybm9S/il39/2xLvh5QEeazbrAWMz2NTD8MxVYhBEd1ICEBOkkWVUF9D7tAb8
Eu2gnFpxhLYKIfrUSOfkInGaSASq/SQ3/38tkc8WILtSI+dh+uX2zFsZkfU9UEeG
WEYvobzzhCDT6L8qqPeVenl8Hx8xtxnfvr/awiuaCSiM11dGVGtMBrThj9vB5X5P
aMvukGBsb2pzLSOI0Nhwq0S1cjL0ZZFOB85jI7yaf05OTMaKG6C2E+CxfofDA9zt
lMwJXZ+jM9jYuFSPX4/+qICaaFwGG6oNnX+c7ZmJuCJAGx2+ruwNpClMcLtj1Y/I
LtblpgDzADYIL8AfrsxC9qLOnP0a2adSg3UgWjlN1MUsmOvFAFywWVwKvUIxpiq4
2+jQO2vLoS0G0WTCMBCwq8CJ9UkxZLCxcY6fpKCSoDdHdwlXiblntgFiEpypHm4z
/pbD1x9dXsaf4lX26IcoZmlqvXEefROS0nC0r48aC9jamPdqab6otnt29wcRYNs4
1H1le1zsNwJC3dAX6bQ93U/fKj0kG/oZhIIcxhbF0Dzhg2/QnhrbDrV9fDCSB8GC
6RdRm2Fpx/fsSebVLPG1JYX4XU4HYMzyL3/temCvAqdL34GoBZ3Gdtu9iWsTyHFa
Z5J4eGpEVMywegBqGN8Tt+hl2OsI9Q4pEiUvuofQBSz/iV7W9mx6Rq1cIRPtYItj
O9oMW7+yDdh7muU7vNTyCUGiqPsoYp3GT9Ho0+5w7JInRgqKMN0S00MaCdFR1Pvg
/r+wTduRP0pMvsYuTZqcrEY8Ch+DV5wNmTlGZ9eP0SqAwvDOenVSP+88L/HyVi/6
+JCFQKTsQp6mrRwLMrDKSrS4THI4JBMZCJV+EVef1J6yj9AeGRSwxgu7M92idWFa
RZiMf4nYU8cR5fbO4hel/xojrCaDi9f78CqYXMbRW2eKbGdKjVs6C/pgMRovMoUT
YuBOXju5zmX+nCa+uff2brCeVeNxvIE0wTqeMDkrg7rFSQpd7s1dIW2h6fmVvEjB
cUNVr2CdwRdjnAptXHjQLScqVrgB73ZdREqj1lhLUNeM0PeDRKhGDKMnRfTnRG/4
BQAslR5pbh0lvRzmqDCX8q5hMRhgSI1LNPCmkqClHyd6Rq8kvsYw7E3TR9T8/sIv
EwFuXNKF2YslI59Ds9Ql8Xi25wmuWhMVZ7JYuRHQ2dlpU4JKZG9+F7rO4yF2kMvf
9jU+rTfgxh7Vh9RHaZCQAHjnWvC+NnO3txvUCTQfMC+NLI16rBW+50y5jzur1v0Q
hL4S4rAiS5HjZf928RSof2MlvhVLvf/PePwytvk500WNiK4g0aAunmUhkTCyQaoL
agivnYmyZdb1LDZ0Ove9d6IHTnL6JyPmVhPXfUOVCT7N4pi/ET1RMrm4IP85Xs4t
EzbjBh0Z9yRaSJ/x3U5v1VijCZQG9px84i3YoRerwowWJCQekgnS1lsPpTDnXpDN
tnjswSsUQ8XIwYjXcXEap0RZRn2dstQjlpfAssLRiIZ3Bgs0WDGrm+DmIvZ13fYe
MCE4LUDXs8K3tnmEI5i0+LjILr24LLLvGmfR0K0KfwuXL4+g7S47wey1N2gKk1qP
Zifmm3c3vZqYaYDdRbCMcl+ayk/m85Y3/TP586q7WXdOwCrG9f3Wczmnu6UwD4qK
x/LH6+3n6P+sIM6KdHTCxO4Pxaa/KZqBFwtp8n1Ilzp2wu1fuYHacv5ugQvH3dPO
V1WN8ZXHsGpRQsqNF7bTsE4g+XT7W4n6p1xCkoC+QHYICV86I0BrdIfoQShnQ9uN
cn+LUCJfc8DTBKa9GDpZjX52Gn+kFRsMmM+W2BH58/SgBUpO0q5IOtlKWak2xrK5
+CnS4ehPj/MpDmhBXnGCDrrgST9Eqr36ZefWH3RKpTcAXb+615HtG76P7kwc0WCo
tXagZg/ImaMGo8trAaQc2C+x3e6AGguabT485dJTthJCXbhj/PwCQaq1X58+3C+T
OuEmwSvLoYPS28eqnXrG2X5+6a/YGTknsLPw9Xic2j5sf6Er1GLIL7tPXSlNOLx0
s32Cn7BdQ98RDJ44d5tckzIBP5zee0/0YrDlWYmmZHAh6lHRz/PkLuIWWry8ITX0
dGZQk6ugo0R99ReBTsM+tGQargU3vDu2LVquAEKAan/jsbL4L/Xzb4DLrpICln9f
EuYTUaUaVZwDPBsfIDCs3ezovBcaBtkbYBdZ9kYMb32/XvKOIwvUwSBnPC20bh1m
hleg74uQ2ZYUEUaZerIbvddqhMNH7YMh3kW5TV8YcvPIJ/T+eO9Vt8Yh7LP5D+/1
BZd1Z6HPDA67gZD6Ha+NnPd6zLIwtGl7RGQzWXf6Y+fD5dVNDFKl7W7/dndoAd4+
cyeO7Q86oLgj8B4sfzC7KsDhy1JcI6HoJ4KYtRKUWAJixoocbDiL3hjUU7pBQHxN
KqBnqtBSojQ/leqL39Gnxi2SVy8SU4zU6qRW9ztRZNntqEQCBlC0Kw2QZGZ1a4Xs
WeDCbtTGYvR5Aj2pilLuiIpnvxM05+9cPG6R0BZFkVonVhjjAlKnjsYzxY1XpWUB
qGba9EkfVEek6mxg7mR4RJo0YCdfA4pkWeRRbvg12RRWj4A2/L/7g8BmMCYTjM/P
HQt0DrMCG37BTe0GxKtwBuXD7BVn+M5lgRNmsKmaUySyYTElnBvy38z7oJi5cCWU
6ZP/HO/li+urXTuMWLIyZCeXb3QA8gfKcUX0CoxL6i2h6azuDho61USGR6O5u4fD
X78LM3Q4IbR+YwJlN1jf4BMI3hFkixmUAWurtL3oe2tfZgOAVJsCL8Uk1aYhfpt9
MS07hs/i4jGz2fbYKdS6VpSMR+6c/Mh2NXN6ZaPgPmY1asGcCKGJus15JVzcDRuE
EnwsP2xJFz3zhlDxfu7+w5rmQUpJEXefi3rcgcahHbNrGPRWK7XTybYjsSztY59k
nIRBnCUJyhvlYl+ff/EclbOh7phv1IQhlxn5sXubUHCd0u3v6psYIfKWHbSs2CdF
CE/6lO2R/Ot6HZPjuLMLqX4oNKvJYM8gzuZsFb7FrcD9XDBIh1HmggFRsdYMRg+A
JofnHlRWN4A3bY0NI7QOvzR3L76RWAn2JnNKq46z3UIjHEcolERvlzbkE3Qnm44l
Id2yVeuyVswIiaxSBePorDC96kdZajNYjsV7xSp+0w9OgEqa4UxTtItVgoRPRGAF
aiW5nlLKe/uOrlqRwrBU9jQ9e1isxv+3Jh0MvuJomVoOlGNlPUyNPZ961WsFYsEp
o2G8X2DTyG154GL7c1QD6ZBPZZLAmv2vAq7Ysm4Olul3JlcH2879ZN8uq3zHHY1T
p7AGLvETcpJncs8MTTuTZmnltzc2pAClwYoTXi4S9ohZ+h7ZzTGmKJUzoUosIJF9
rpASz8To//OcsVGWm2n5V3MeA2IFaSmYo6qzv5cL/qg/2T656V/k1hDbTmUp4vjq
FqxRx7SpUQhUksN3g2uRH4e5XgDzc6YUf2wQQnp7VwtbvDkpLY9GFbSxYGMOsKws
va/GwOhhzadmluPnRZAEoeQk8ZY6q19PwcijFeK0PM79CK3x5r+Kb4xq/RwENKM7
II01GTm8dKyE+oRhZuo7uPD0X/AoSm5Jj9IP/Zbxk+o7PdbHsttv48SajSlj9rAD
4wyQHu87B8EXcw9pje9AbZGXQmA6NmtkQArvJeOsi7sW7FCDp4ZeZkTRI/2kpxAU
oVj5tDTJmOPGyu9BJxiS8llfIVmGQHDIEKvBZIvvwHzOjiiqDl9DvhpkgeNpega3
won2yLRlI2g+3h3K6agkWicN2T0IFSFnrvxHNEDI6SWDVwI3rqzw+op1sY3t+Xh1
jux1RxtBJYxXTw/i2duo4x/BfPugQaUlyg1Kvo7mTQ1O0uE8gjjQOXQUG2MdfQ1u
erW5NZTSYYFFJcJ/E+YkuAGjIVwXK5SaqhkSHi1nJQ4ZWo1bSXn1O71f0AkEBa5X
8QXfW42e8s7xFyWf6fHr59oqd8qPRXazOwAmzn55pDagtwmWcI3vNrsEeh2bE4dL
fu9Kzz9DCu+JinAGLl0U+fLe/MZm9s/SsNNFuniPinI01ASkIcht1EPJe+4QjfE7
bOFkwUempEHwbILSuzXwX5MiksYMKY4r+u9j8hRGy5yWywYYbKvy/nHLOYxXOfQb
lEMLb8/XaVcp2EwTqZmK073GR7gTFB6tvLsK1kgLdoEra25fyiKvnG4w3VBSQPte
EI+nzrRXRunA5Qb+xdRVk7n6glf7bglcvfc1gxEvVQmskyN6Z4xZQ+h70CdAOYoB
3K+4lcAsA62pF73Xw2pIw4y2deDc2oL8CuybFf4THdzJtyWbfJzx9RAbdRDmaG0/
QLbc6/hAVUFSKF0PwfIPQViBxlrKPD4V354QtaeEj3q/ZXR3IL/uOr182NDkt7Rm
NPGuFyVWbuPo5HZACuwDrYdKgMG8UZwslu5yc51Ip+E97edp1eMRYOHwBpAC5vEY
/RU7FJijCC8rflc4m1HXsxJuE3PRbSp8vFHI3E+HOFXHTmqi3ftvhWNNwVWYAHR4
rfagi13LGDWwu9krctuMmLLFWkNHgDItS8Dn6dvha9y5QwKtkn7whX94MlrwD3W0
9Aql/8ALIqHdQHyf5jWQb2fNAepO/WQdo1npHeVOdIBs5u7uRONJADxEmQe/Nexv
B0J7h16S6/vM5WdPPovkAwdVEWGu5IpermX/HBWtzjhdWPH0cs7tI5POf2Jsf2Qk
oodKXB7rPC3ouqlEXfID9BTxONwaWjWSbHNqF7vmkPGInhchDuiq1YfgS+4RKBMv
GjgHtR//sHyKmziG4bAHfB2ymTnZeTHMU80bTWddxHJLavvHDgV0WKBzJgiDNS/l
8g2dDN8i0RjyqCMkfBqDeZCSiLi/DWhQ3AZHOBpknS57rbrH42RYaRBDjNTknGVq
M/K1L2dvjvSuFYQVNgXKSPIEQnrbI3u/WrwcgZ8AhZ+gkeO2aJRtL4rwjuOsC6lg
4nON0MpCrb0djpAenB5476lXfYVFXT5wAXfFTpU16EO1xTayICbWyCqB9N9BwnVD
O8cKh4yxNFmmMI2jsX26uxXD/+e8wq5wLE4sHgbJsL3VSwdU0khwT8svaZRC+rF3
0tF4dB8QohFW06KwdgrYLeWbPHZZKo2wJVu1qhq/J9tmH7+4L3JeDxKyZIsEnImx
F79IQ7S4CE7ne48si/x4O+I/i7czdhsB1CJMAeV9cKLExHmtehQ4HPIf7Bq9/cEa
HBGFX3Dk9Gi4BiIjJ52MCBAjY5X19WzUW4i3CLWJrdbL0+xo5BEWJuW3Y0fZ4m26
xEj68HN9OeAxzNC4YqsH6AzKJ36zi6bK10mLkBjDFSjvZyBdZqc32akBXSGcgJyA
YxZYCGAsvjc4m4sMNRzJI7Rsu+E1B7mtwbBJfWK9D0KOto1042bsiK88P5R+NsOO
LOU1DT9h9hv9AaqiZ4l6KuXfmnCCyTqYOw1nMvTevBFlFfcu0dp2O4r2dpiyZOJq
tB/K2rMDbZPtGQE9VM5+H04ltygDe6zue2pekSVSyNzTZdrx5t7wbp+vcd0Cxfpz
WVUFX0cmSUV0tCFey/hafchXVCnASKWycmHt+BdI+MZ60MLPk1ZPYWZ7bfSeGnn0
Mhqrk+btKisVCErjAQ9BxK6S1X1x2HjqZWm7PZgwY5NOO4Wo7BSvVNQJXA8yq2iu
g8eENJidsBKTP4nwQi0PvhfcX73BdpvE2uRHplWdYdjpx/ow/ZKzghJCEUwsvxY7
cwu9ZIexN61u3sAeyJgJmZu5n8FBFgVQFN3ToC2sYXTIN36dgbkKWd3Z69xni2d8
hlH45SdP6wUnhXHcxfCU0u6pD1zANfP4v0yyYtaOV38adF4cMz74qwQ1G9QOJL0u
TKmuFVzTTktQFyIq9BRebVmpY59WhClX6kz43s5BjsPNeDsTRK3MjCGxmobujGuD
8oSuB3OkJe+72BIHfife2ZKDHR/X8HMksH09KIPE9g0PAWA/R4qjncesoYnfAgsx
eqK7gf/CE9kcLEV6PbApjRDZ848xNc5hON0da7OATaQYqB6ShUCVEqROzzNAePgD
xgohINivNSnw6p3J9IAJLhP0PSgCujD9jT6zrA2asJv+cjtJ86A63cFZ+RUYYwWg
7I9GrQb10mPPc5e7nGDZf+HV9tzpLmsjPTvr6vZ89eXKR2FmHEAaB1dMg8rGLozN
dKvE2tRq3DV9vwQGn5aJ2NS2lJjJsBwDak+kBBHrQLDVccX5JsZnrIQordqn/fA9
7TZGFf2QYAxhgP3TB0iAHnk1qcEKaAoWCMpOqa7+CY6s2rmA1jI9EMxLDJSrGm35
h29HSS2xZlET4v7HGJKCN24U0xYzdz7Bx7hhWBTyv3ctj8RblVc36lrpewZKbx7i
Mh7eKW59DxpICuMK3N4PaA08QWTAH/V/ddLE0SDZ8LvaGo9ViigoE5Kae0o5wbBp
3sYIHvOGbJsj7bO/u/wCy6EhVmU3aWu07MDvH1uxT9VEwoFy9vBIe4BRWX8BCkpL
nKBo1Dww+8mfv79+zfWyrwJAyjDQpFJR7DLMyPpv6yGYQPAk5uJI7nOtU3qzSi8U
Ab9FSZVSdC3lz55c4/Rm626Hg5k5xZdlkFn9Wbddo6R2YdxEQfakEQR5J7+Nolkk
BXWmoa9WdvT1oGDO+xLyiFq1EokCy2XzpQecZ2Xcg3LIUjy6mUMEiF4KOl8Vv2a8
Jpu2p1lyq7Zhx3JmElknbavm47Ain+QOISn1MXDmFSlZtmBvpmhyLs61l1E5qqyz
tE29rm7uOliX67PsAENPyTrOPsZJVwu74I9FlHyek0uxvmpOdALI3o30sUxaQ9Zh
v02aqw9f9fKoUI35mbmg+dQNxSj4Vm0d9sXLAcmyno9aTQEdfPmgcvRAknOASL3R
khW0coS7nZMYLLuasZj+ts00kVq0qHZ7M2UOM6jFpKdRsgiJU8e5bT6+1lh/HbEf
pNZyrtxzI4bd7wkv7lPUfImTYGcne5eOpuOKl4Wi/PFgwGRBgaISplK3KwyeXEbM
gbO2nVwJtzB/zStBD1A/Sg9vgtqS0LLkFRT7Oot8uSRRjwLoKDqsJQhMBK4X+fN/
nPPDNpusegJ/UUaBthrgW8eIL2IpzY0AbOYo75yDkAtRkU/46JwhIoAIGqwJdSeE
xCncmzc7ZuXdAE0EYYvxZs+Z7UU4RkYa1qyws1YlSi/wOyjmT/snEsXQY1A2YV08
awSg/gT30LgCmmhN/9YTKWCmYVPLCFUaHW+VNKYJ6LMAse2XhUicpeWczybdPvDO
owgB3E6JzUodAiCRs1VWBDyDuMlciMqx0ReBtWPURA9ukkv3nj3dZD/GD6jLIn9/
ONg8eqQAiAip5KVkEQIXoRHoXqgqaEGOT9XsBf9tvcOk+V7NW5y5HBZ/GJXLdKdG
CjLtxNBLYRqWnf8hc3v4aIYGRyYxybRnfqNGc1897m+gz5zY0LURmkQuwQgZYX21
ry6de9j6VDR8rLOpq7N41s4fMTu24gD+/vKioby9Dpt4hIChAxuH4H+wFPS2ybPl
3wkNGM4GIvcWeWl+4ezS9S1+CfzyL3kPtwVB9hklUuJo4991cYF8r94l49bNvMAA
tgWzod2Un4pwojNR52Tx9ztfiXXAvX3VG4nPiRhykboR+nyAy+W77wk4fPTu73QP
1siCcLNen14uOTtfVIpqi3O/ftAz61q6v7Ha+7ux+YVDKwh1dKjKfX06WFQ9vcqA
sWD7/8S4e/aWF7AYT+ZgOqAgkINoyCBKk6GE41Pn+HGaKlo8u0p7TuzlQ5YdjnE4
WgA4CiEvZ4xnQdNNltvoWFDhaIB90Ms/ec3hIl2kW1QZKWyD1+odMnYMX/6YgYKW
nGmoimJgWkZ4EJm6kyfnnMZlxgYuU0pwDiYhkfjs8gEOhC8mqfKs1Tpdm2mqq4E3
9owj/2oEDpLD2gM05zICrPlLRimtVj/seH9XgiSquKIGk7BSHn4TmCZUyNbQCKdT
4TjA5+gBXGav+UptIeKwi6ePCZgtpCH5UPc0eH/fK9vz94Cq5w9PUEuEra3/V0g3
4yJe+7G8YtE6eiUSfhgHAKUCZewQ7kJLogmFhbjqD2wfoY+J3vbP4BTQZ7hCOEdV
qcGibS2P6nqoe8HUK+zrGrYKAlyFKW5D+iXjUZCpnBP0NbrY/DSnQ0Iu7qTiFSPL
qP4YVCOPV343U0HeFS9xAR55H2rGE7DPpGUPDhn5Hab2meHcjRxnE/vY3C9kDLn7
9h5+o/+k7xLGTLOl1bD283OZ2Kfmkus2aKRMrVPdSHW2PGb/1pZe0V6ebViJsV+K
1f2ZzDejC1kaQzJIdL9W4KXQUYFrOi6Iclb9JmdkRfvcKl/Sh1KzSISJXkTLC4U1
7DqusLeuCyX2swwn9CoLgD22F2skW+XOFONKRimLHO6O0YH4rsMu6+1CKdQbGKdw
2ej7Xac3DJWIRXFgShyb9d0pimGa60lg02ZRW0nbwX8klSmGsJ1H1GM9e5Y4MYRA
2GQ8aMn8xiT6pqkM1EiDAbyABlgxFwasd1mhjaz1tKiVZNYvKTb/Dgn4cVJCCbjW
KFlEXaWQ5HbWq6GLWG50YICWBpE19Wec4A/IF0rixmfweAoXY3vd8Aul9bANtlcB
nhtCZ5dJ+keGdoWIj1Z73uG1kNb0Qn/5BNTY8zQxIp2xJpdycghYdiKF9W3ga8KZ
aPm/xRG2ghtyMqSsAl6XWbW1XMD6Qu3VmcTzsWXU+ZAuTepbO05JUYN0Y1LY53MN
65fW1lepAk7RQTMFPXB08acE4Ow9sdW6qHHfu7EyQlEMPUvIH/UT/3Fj0nlRK0FZ
Sglq39KX3qt69YnxoxO8V9GHEccFSpdcgR1Bb+6F0xmP+4Ny5fckEiGahjJ5x4mA
lJy00tlHDxthl9e7iv2+Ajc9opvwe0zdUI4o6ELBSnzNSuROZCtEsDlMSaV2bkgo
E8d0ivxLVNkSXp721H7vL1rohq9P5Yhxcp5czrrq6+GY1hOqcxzavkBusLnHdzlh
sT/S4KYBYXtEnBDb2jvhDXtewBCOK8/3rjaQvDKqP2RkN/ig4FyXsWQyKmggUf6c
39jLJ2Uk8hUYUdZ9XZ6eu46Y+1O2D3FjIGNBKvfuEF4eBglIMzrB7LSvjVl3dpAW
or/D/lyIAEKaJwSZTDPJ483WUfVq+uxkDrFL6xMiOg8bkYG8jpgQXTbYNrVjIaRH
7thuCP5mh+lY2sbj+PMfFce4lLeWSJ9Z5zxIKnkQLlv1S82U9KSPLvhfowR9OFee
AQdPnZT104lwhEACmPMQ6OJjjRa9+Iqzl8hH2n9fPfEAHR+wpVtjw3Qch11AJ3mm
ozF+4tFg+tdUPp91zw9HoTHOyDJvFSOSk9vrnGPZDM44imIrtAq0AkydHx7RA7a7
XyETOOiNdcV4QOmFx4uthXf8N6DOm2YMaHwOx+EnBioo5NDrJk90ppDgnF3GNSET
FGOAso3SZRSp8Xbbqflxts69MZaUfmU/tpcEjj65vj/n1m0EEygpXz60s3SqLD2Z
dgC6IewEMJvpsoaxmbD2Mr6xp/nFiqEPVYQ6AtAmG9NeD9x0JxVO2z9yM+AB3SlA
rKZwTIBHjrAzd31rBSm7cMp/la/iIUPT7y1uX6MmiEaREljhsrUYy9pxndd1aD7T
BLM+3Mdz8eWTD2iRP9Cw1pagXQIy8wjJtzC1EZMxdSQ7kxHZ6P1KM5wS44DkADya
SBFHqUvKPoThvUpiQ0IF1X8nMotcuzO/vM3dy4ku3hzQHFKKkFfriSpo6pzzgUV9
jr52yXoedg48vpGS4RT405bFIFzMf1vq0HNxSVW/ZXEXBd1q5TmbzD03psLQmX0p
uZbDvWZ5JoYuYVJ7hpxGlhYJL4IXOGpyyvmhg5oXZT/akycPh31IRKG86Gg3D98N
FFtePwD8gHD9TLK3AXVkcYPuoRiBZC1BKccfqxsGoenrAmfpyYmKh9o4KsifqHLk
g38ex7VBNGYJWvqAIOBLPjG58Dx3O4a3k2VuPTY49mDAje6Ap3RpyHyEWOFHB0yM
difZUu3DjkXem49QUid7FEuOB4NPC4I12rPKndbf4QmRRIIx/49CpjGoml7bG/aU
zXIWbEZhZUBzbxLH5kUi1Zj40hzsY3Ftqk7KXDdtj40hESr8d7KnONovEAAX1uJz
CT1lqvwEHu4bFSNkesXA6dSB1VggyGtXkZIDA4GS32SNGw500wl6PqxNcWONP2xj
fhU3v3IEAKO2bgYilgh6yAapCichDrjx+0H6rJmeg9BAt4HiXx5yM31i8JXiFBNV
9iCPDjK3jEyBW4OQB+wzzXqvETyvBMx6KJDpnMEUU8AhqByqH3e3njdagrxt2XFT
gJpGGS6/Sf40ZUum2icCT+QtG8yqB0fuadxQ0WjvAvSfaIFOTxZh+jHM8pnPehcs
z9k0O2r9+JSJiEI+eMuM2PA5axmnR+XFR0wEeyqD8pD3ED115RaYdRKFYfHXR7hd
XcxmDJlBrTnAT0wA8vtNR2PWIHrTJYXgXm5M5d8IKEiSGWwzPv05QFR6BDsxIcW6
iCmxncdhqKWo3K2stqvRNPzkslHehy7y3B/LtPNCH7v3amyYyXn/4nJ5pU0BIW+s
ed/8loJPHy7a12/3A0JHFg+iEtiuuA+uU7fT4JV1V4Q40gas1JKKmHl2+9gaA84x
7VNd/RWtNN57OsjIX+RKmOTui3MVwsotxkcj8e1GqfGDzUduAWP0JMrR2QM56ipC
ixvFhedPrjDOk5p2rywejLQp5KWI0rf6u/V7qeGRH79qErLUs2kAh+Ik38NMvqzu
T+QRiyOVyBw24wDam7/1ecCy2b6QBeYK8+qCWBsvWSQyFd5SU1F4YeH9VU6ODB1a
dA2GgjD8m/NK4yI4Wh2HrYufUgVTrusFLvDpTu42NMfTqkwBnqqK7U+C8v9Kr+fS
5hlVYSREcy+l2docGo99+kkdGP5DpNfjSIWAZWLp9pI9iZVE6il3cXGXIArurjDY
4lMzfG05n2r6mQYD+OJ4LrOHHiUgMsXkue1IJmi4xT04W7TytnEJQkfJ+Eg/h487
p4EBc7heM9q4N4gFXMakbPhFHOCnOtF/7SI+LXO3wA3JtFihbjteCjMWYYVnNQqm
0JCgludxJknt04rfjRToSKOWiLQs1ugl77zR8GQva4QJUChriTfwchxblFUx1wvM
hAHl8BlUXX538UEJaSpPLb+tVRhi2XRyRBLR7WkRacG0hRfuq22SP1g2JA0Dg76a
/Uo5Eug6XkIplSZnnfL+fqdRip9rOIiJhJSxzus9xY8a9b/UkIipM9dIvw3ltPH0
rHXxWi5ofb28rXw4COnSS7AaMjsForPvaKcuWGfuMgzaOs7KSscx9+jfoxUUuDYk
EIcV/IhV9Yf29gB74f98wZZG/gSvq4WDyB13lCHB8A7yoI5O3q2klULkeg04LlVa
g/4JNvCQMFA4uLDMWPTFHgXEHuMGyMRCGEuqvQ8jjiCRh0d0wdstx4k09/MhnRPv
sdQNEarj8aHinucZWmW1tt+lwMLtviBfB0pl+ebuGwuyaSUzRwUxEYlappacTrRa
VS5+T6NYpnIGwBSXsUwuaWrlkph75beY36rnYsKoLFHp0kcnHnJzPIU32sRzw2bB
RLnTE2uXfIpgS4G9xDYDsDxiYW2igbOdmK26V0jGSuufikro94auCWu1IWIsNNKT
+A82EbgcytP8kyyEDohxgcAH4LoYrQOJnrma6ZAoD8NmabbcQse761PaDKm68OHc
CwmozdXWT59xyVFrPO12kU6yOY5PRBV9o1wZKf6wBYbYmgJEfbrQFKbgHn6ZRVfW
nTIE84IsWiZQFYuhcAE1LgfaTGZY/SEoZoYnhpykwdhGUYfuToSP8Y4JcGLdaJkv
n/zhz1M3iwG45ZA52KJ+nZn8+K4vAj9wxjQUYgXBDliIyy7XlTuisR/GZ5QFQAyn
Nk/KarCo4QoZPq7ohAP/1IoMrGK92PCzSNt6n1P6tRNs6WzdIBaitzg3rbEXBrX1
U2EU+eTVwdmuu1Y9U0AO0qQi1G3bboha9B9cfC817ptDR2ArUVvs3m1DwpqjQb5M
vMby5f4/gloUpBHDJz51jtVnQazyOa5+ofwGGgSo0tKuloBvj1XA/XAZwCP5j5hn
9+B8RZnMd/bu+vYd4zplzN41BHo+UfwHdtsMUeoLg8HHuRtTgjAhyxU14Wm9qRhS
tdAdJBpPDRLBqofnE3DH6+oR8sExmK3oQnMikitQNBAB2e9Tb/ImGfYlBlW1caET
uaOyyMIuZOltBDS7C6gdImhFRoiiwJg8fqKlyEzepWN15EEq421Efh6KbzLqn1rp
hCc8ZHFI2LngMGhOCo5bs7skIMxvTPNW8nt1RXqDizEEquWYFFvRKolmz96qctRm
JPmXDipyK5Y6YTSAlwMsY+vpotpkofzlKx7zrQxQEy8AvEdZ47/pqMzAe/xBGjqV
WO6l1+QnrAZX01lDSveiQtEfDgy0e5jvKmBEoogsAs05Z3gyI8lyaOBWhbDtsYQx
WXTl+6vGYc3lzyDcgtX87s6lHfSHp9VlalVHKNtyb0mhk7fn+QfbxL0H3XOv7X4h
a1TbuRLZUfc36fsaK8RjMtQ+FOXjAvT+jjr1wATinrb5WybHImjrgfJsGJJCfkbw
A+CQ0Wx0Bw7u9RVO5GJB0JDcFwLnO6yJrFxIBFS4Qi6E6Pj7s93tOvEZBzJKdqyE
fmO9PfVpbUpr9f6awuyekcI/bX3zPX26JLhIcgLiEetun0ZB86GwJLQXbI8rOXze
5n9+LlZaovXwrXjPYBQimuARo4nOskGzyeKaSP7DCGdQN5ez8s/WLm5y+Xt/VOqV
zhiRNI542exDaSV4odKKAoZLkXlwZPesGaV1psc4bRXVgzjDXCtQZghlgst4Sl8g
qkQf9/4hNV+B7Fy3Pn8keOVj1ry7q4V8t6EQgCo+rp3X532fKxHkCxuO7vWXSWfZ
z3V5gzTWiUoKDUrc4OA1Q2f1/QqEO4qiTQr1gs7icfnOZMSCmTffe7I6HtIuis0i
aBcBh+qaCT55Aiq7rq1kQ7UgduvIhwRqKQ/2UNGsS7+OW9G94sOXLMyzukJAvN9p
XBM5sOWJuuXpqD9QtHelw463JFUZPZppwqLVlOScbjx5XrP4vNmFc3H/kh6ZTH43
rxIiEicak1BDsi2YmVFDLcycG/IKCdhaeqrnZ2ubrK1K+fBCw6TVoqBPDApD+foA
dRww5eStoPBC4antc8HTZsBZucls6DGVVw4ODo1Oa/TDz+4HK910B1QAP/kxee4s
l4DCthxIX6sVdS7bsUEGpUki01/valddcE44wbqdL+RJgppPOSTG5kvh8AfNIAk1
q4ZSIVtTe3l1Ri7TMhY1UnB1cU2HzLU4r7BFMO6K3pBCCIp46h0gH2p5e87831sJ
iQTHF7wuHUI1hhXWbe3BrFhgGYHIr8LPqQTlfszeH7RgX1S7eB3dBg98aTi8D0at
u4k1JyrtIXBwkPQ4Y6F4Nprh8jcyjyp01gJ5wNxMQQQEcsCjEvDOFuy30lqgIAtc
zEhYKvPPIy9MVYCM8cPjABrWL5n1GJlXKu6IRz7b9s7mCKqlZY5VEBq3oLzeQh59
aMnzV1RZgUdD1/e6rctm4T/m2+71Ss2Spv1Db1P9T+Ne0/1u4E3v+Z0+eOncgZLg
Y4v/1BQObDY3zJ0QcIOWkQ/cHXTm80GRdfHcDNQV6zzUJPNOjsxFi4jSEcg/kC9A
7CgspvfLmYCchmQXJtXJYNrBT6bwyznf2WJTyChU2E/HRnDP8y/CHsTzpUIuOblm
m//M+1ujKYW3mCMdHSAulsUZOrxLQn6raPeCtVnUOZE+1arCbNjLUZjOZTfbXaEZ
W1mbOzhdeSb1r2uWwhHH6ceoF7N9HiFs7ZnUOAd3oZYGXLS5sR/UBFde1AicHVLU
33rzWV4xaySTRF//OIW7GBaKO/y4zBOb7cUJj0JHLQSzu4SRfcC3EiVtsVv4URKg
REVmp1Zvq4ZdqdGVfGj37pdwn2v4QldK9ViCfvSLIQ0iaT+MgUKmyCv2dtJNIXC+
9Hk5aSMueSW2eJH9qB3mtufM9+//9ddKscUWmHY82tfgNtEfGOhJsph/HL66qiAa
iHy7TinWTxIo21Nk0GvhYNzkRzcEy0tjb8HadqC4cvubY+aFQR6VwJLbLOMztdDT
nbdNHAi3uUH2SXIro3YVgPPDNCZ4cRoDt2nwsQkt+C6onBj/jUSwmuZhRNpNQj1D
7tuRzqBtOHozJUyCHdkUizG2NZs98xCLIJ3h6Qy3SKvcR96OuL8B/iaoyJiWZBIU
MmOt4K86HJecyqUTHABYe+htIMt8wDgTqYcEBi3/Lo0Tmg1WADEhvLqAbLL6DSN/
iJc+oK6zI0yq3I0PvtkUZ1ieP44wT+GiKYcqff8LkL+oiRwCsgy1dDqDd2tWc1Uk
eoWfwonGXIW3lTegHV0BO9OKsVYxBKmnQKqWSI7TgWzzwpcTQHdAPeBvUUNMr6sy
ofPGIDKYOcvV8V00sGxj7Aqt0lgfvy5iB6s5Hzdoi1yHuna4Ee6E0fv6tHL2psvm
mQf+ZxCEgQw+iQ2NykCJCqTgIWjBH9ZPuQpEKGYE1V8inMD53IikoRQHkTR/6BFM
irYCgLhf8wadlDOCTdLhrGZjFjO3ma8nuL5JE0DTkDswAeKA7LbgtlqndDahgP86
cpWSrt9D9Chf4pUSLdz9jMUQk1KO6K9vQgIXVHBMPb5iO49r8gRmae+3BE0TuEZN
P10u3/CN/WMyaK3+8lhHhHCdxJECkuj5SIzpkBvBEKNyKCC6QR9jJtSCQaK4Ujtw
a85/Bd4YLfj0OGzMq+E+OwVYMBOSfbTJOQpN4q1y9RAek0D4JLHNtMV8JswHKBmQ
RXXpVRhINPoBmXSudakDZ++Uoawh5UnxNOgxOm1ishT8RV9vkxu9kRUzQhGUKSSw
Yd0dOXd9CDIPC2y7n2xZGgKIjQdnCsLOy0UgRlL5eOM1LoIigW19WDHtQe8al6hA
II2uTY48ZrMYdwFB4Cqxdcz56w8mBaWLzE95IPTVM++GIqHuZ1v5Ijz3rK7tk5Rn
P6ZCa0o+mv+2i+ecvLup0A5zQJCFozddiMTULMrvwVGGA3i44XSDa904o6+73gRz
Qk1KQWcisGjjFBekg/fFVYhgJ+OIymLAA9BvrM773AWs7dwu0fkCD4wEFK6qJDaX
ZMHb8ql/cGL/0mHi1V3n58w+XJsEf/RAlqgrG5zo1sDGFJezpvemW4AcDJHeXSqE
5FXbFTBzokeX0JvpB77QhI9HcRrUfGH8Q0kOurBb/c9okS1Muqz7fvABt9W+li3Y
HJybCuw5L12Uj43KUXAr/SXjeO/eiBn/1Yds1kceYdcPLSgqqioPh6crPPQWwh+C
hdd8eC5HLXkAIVtCytSmNYIBd9iENEMCLhp91G/4oFKtUoseMyIt/61NhkoK07Sk
UvVR1PDfe3928fgwpjYMC6yscjRwjF0Wp6oUqk3MLIBg1EfZySiLt19bnG7fO2h4
ILpHpj/o9JxzIFiRWR5PN5xMC4eWEt3rFKFUijhas75v3AUjpJLe6MEJniWafkeO
KVMSgj/ExreIOhPLmIfwtBIy0fiEhSEENhvj7tp4KcT+PDihV/teMsDGsnr9PlnO
V7WjtWrL2wOGEHxvdc15t5QRAH0+30AGwWqcu4qmPnWhLQ5a8dJCYZJeR5vsbV+7
hAnA5tFUoYTbVRs/xzLz3ZzWDcdhMaVUTEG8be7zUmRo9HCRyMLCWgXW22lg/LD6
gofaYbQVw2D0lNY8CmCbOj4XsHqook5GLc9WI93e7XTSPTPqi3N+emqXile3dFfV
0pP1wSX6QHXTwkyEW7d2S2Mn67v+95U34WjLbmFGp857H1pzf5PD8vNzpgp8GEB+
Njh7UWup/kxyAdWB6fqc0jEXehyzAAnTBuRwV8GxuRO27ZBnCcJ2C+QdKoWObj/2
DjCvGXmSAM7SGboETTi9Pgz+laq6z7+JLFy7698N52zKoQnEvmXGl8PbDn4tPRJw
qhBsje3ix1yhXVyyNNDFIyE88QmDmjG4xINg9OqOzmvd87Iv5ju3f2q8fIiuaFh/
en20WzCDA3bzWwkvljzu2cD2T41uVCk+XUf2t/rxei1jqgRez9TCDyvMr+qobjVo
rFR0OqlX3BAdMO/GHCnAiXspinBpYBj8sfMnqlCaIgBXNAWYE52YhJ5LYX03/UVP
fNpRXeDnYfRHZudpbnfQjPAcRS8wGbpd9CSdP5EUr1ekskIhl6ndcamRcBscXaS2
kL4+YeF4D5BdvxXlcyfR/TNgFIT680wOWJ4uUuDw88CbP3rBzVjgtTuAXyp0r6HY
l5NzvrvvM0PMdhN9QGxczvy/Q7ushGV42KGItR92J1f22VD8bpfWCb/eJ6yWH0Gk
jLg1B4qR4iQOcnqBoR5VwZ56F6i6/YQEzc+Av7WpIYcaKRdaiGnwRfkkc1Fc7mFV
ZC6qHibMdglTpG7uquQ06PC4eDmj6T5VJj4lbsfl6aAjeiZjV+y2jyJ2bNQRxBi+
t3PaB6GqNxSrPTgLSWGNgcixrNo2DGSpBgwn4voCZtq1MbV6e68iKZmQiVxfan5H
RS0EFvwzyzvuWXHuV+MpmxpsGu1/Hmcx6VXo3gdjGbs4lVCIa/Dq5MHIzSeIOStF
4BIfHDacdT4xF2xee7D1uGLv4tlWmFljfgSR0uJE0BqbpXwUt1DK0ExJg/FN708g
Eakjb5BVdTdNLRUGyG8SchFzYInDX1I3ud+14YktMyfH42m7tKWvTztdgwfESl6O
DXFJMKSezJ/XQzfjNod5JQ5hlMzTCQuEFbsTINEXd5fV+3nFiXxElEYYH8oHWpbo
n+ctaCJbAv1VP5Ci/wJFLbmvm4UEvmld+oVmZKltRUpG30kwM5L3cDv1LUun9WEd
EbzYFtgBdrc8wg27UWhu75A2Q7dJbcckVdYg3uD4N1RWuNSqOpokKgRBxr9XEte/
UTp/feZuMrLT97iYTfHoNMa9AgEfyDMlcFrr4EnYCIpOxI8r+KK/lqv/cD6QIBwt
qIb9XDizY8rxjiUcDmvxzbTXS0YvjV0q1AryOul3GFa7u+0TDk0zJh8MZNdVHyc+
7PRQRGYjoDm9bhCBqUJ0XGlJ245X3waJdYJuMFS6ieHkzc4jcjj+LNOpY0BZfLo2
jyVvRjwKNLQkALA50mWjyjQREj5ewT3blSneZRCol8iFBPOSLSxB3+8I6VmtGs4q
i4mrSMA2DU5wKGecV1Xkq8ZXNlqF/HEX58xMiqsb91DtCoNxd45HJmqJnimQMzDT
QINt8QFbBPnLv4LWAwgrhjNMMCfrgTdTt5kgB3t5zy1hdch4MDIcJ2jqNThohxae
YrDxi8fFguWo2z27oQswj/HQ/NmdynYSx0nBFc6IHPlrZ5GcHNRL6MIprRCjwdNL
qUq5/NK5jeNOfX+USIhc8FZaLRYKQCodP029oEyXZO0YLhwBJggJ4ogI7ZSfhoNn
tcaibSjqp/QmqVjcjAs4tk9oNPfvYnILIi1wRY1i+N7ucObFF/3Fwz73wTJsspwF
dVQiJdo/VCN1OTKLs/fMQYszKVibEo79o4cpARZE91g4u5vZfw7A8+6WWGlEGFbV
aFs6rq0dHHIFuawKgH+grF+fWaaYyt8WdkcqngRtvmro2+3t4zYuBKW5GiQ6CrIQ
u2jFCVjcST0LK/rbzQa0sbCrdaCtIZLFSYsiICXaCNzW+jQk1Fy50xMShBciVAZq
f/es+B9IMP+6lOv7/DIXMmNxrdIT4h82E1CeJNRxMAYAgRXwoyQiAUgZWF/rvygS
cKvjSmHDmcPVHuenWFzpnuQJx2oiHqDSVrL5ApzwqegAgjILBmAdiL3/5Yijj05L
pSObi6ICHFoksqXu1ELYkwUTdvb3SEhuXET0RQ4TfpPT9+nWoVAjAws+akO+f42T
bZ0RXJihpueo8uJiyR0zpRQEcnhXAr4iAmOM4h+vZORsOdVsG7+DxXmpfl88ipkD
NsyHOkXv4XanUpA3Dk9SQLdCaMBAafewWgFpGFtQsIFOk2rvztn6/+MF/60qRkug
T1hh84PhkC3nrbFqUXLBuUiyRYXZvCfVp8DA4U3RDgJ2ukno1LdsBFHavSyLWPye
A5hzz0aE6fL+iG52xwYncC6T3Tqv/iLO9/MksxyMpCh2fq238WvklVSs4x0vYQFL
eKA4UWjl4Tr4+7lqDfAadRCWIPQH6ZA7+uVzq4sQe9ciEPmbo5QkgWKc8mjc1F/6
glG5nTrBVc0O+g5+OPgzLMQLxKku73qXQhiAkmpRIPFalondhocXpLfJbLi6MVR6
ZSIDNLX5wNyK8fBBCPjbnN8BLdDQEpArj3NerjltL637A3rfCmh/IBB7SUlMk3ZR
Q7OC21DYfcNMUQDMGeF0W3AKklE3q7h4gREg5947DclT/BVrZ8oNBmuXtkwmdMzk
Cpqu4B7KVfTSEX/zzwrWxqWmQEiP8zNtAeJvS2X4Gt2RP26dzNhArALwHlqDpngG
KpPG1jOwEIgvT94li2dcIoQMI966uUD/jSwKxllpubPp/cZCeF3OSOTqXKEBS2ge
aaeM7mEcet1AscLaTIGxvi/eAa5ce2raF5yXBjYquvDC2449km+/M6hEcWd2UUvQ
GTJZsAOsOH2sXHO0WEfTGADQ8UdahO+z1iP/PyIFp3/BaFV2dxovhiLNDcfTWRa3
4EjrI+Z4cbaHy60cLN3XK1siDp/uIIyvY5AXzV9/vkwu9gEBdjvksFke05GLkKCk
foFtsRwQll4S1P7S80dU8hH26QxJOTjoF7VH0HpBq6zcYaOt4sX4p3Fe1nk8MBcm
EKFjV6yLs0U8AAlG4LhWXYrbRTyqPWpYw+/fXAmV6TfGPJuK9cOkOF1xZFwF2tWT
he+2eXcHiT/PuyuiQZy4Zs55VUWwa7vUbRNecgnHmDO6XfGXyJsw9uT0X9dE4EYR
c/hQcM0Q/qK/FZfUYluHyEJiON6X8ZuymVegJbLqQdtDDkXlZ+nwL6ZNRLWEK1AB
9e11ryW+kgNVfISpu6ZftmbwugvxKeKRBWW6Cfy2qgKgCJnsomuX0MMnP9cFTqR2
XyWM1ltYahgA0+b/M/aUckW1RYb3vcu+7RHhhcrtQjNEE+p48pE16hz8qkq9BkPb
dmaZmiGyREBZ3ZVTy4P9f1inayxWJDHFV9uZ+X+Ef71clFIBB9siPcwmhMbh/VmX
80/PNHpG0D1lCCErkd6nxFZc7cICgYU2hwFjkLKbVobEk58i9/orurC4uAApRg+v
m8J1855oRBzks6DsWHdoH/DLfcImCoPeE1n6q2v7eaJWBfI0HfNA3vxcDYJ2HQbu
gLMk00k9q2lN7jh3eu4xfl8/khACYFpGHisixNeJwb0tzvZrREERUZ5vEmLQPGAi
vHBkrWF777vnJm93N68Ofweddq6VYLGkdPrLlPUHWfphKIA1Yo7jlV3i0OQ4DkDZ
tUVCBU2b8n9IyWSAuhlxx51l6IKChNsycpkfjnlST3UeJRZmO1bxwIZAy9t6G5KJ
HBywW1fJ1HuBX1PRYCpTcOukZNaRwQdvnBVI/eSqBAiAfdqccHi9m56G8mGii4nq
AgBa0tvR/PmHSxYvr2dT8mZNOsudTY31Sm3pEh9mVh5izFFazarcWBlS2W45gr/c
/1eKIpBhUsXz0GpocTF2sPBRrCHbHGaVMKpRcCypM2crwjaxNZOFEd3kuaydsgvs
YhgFjn1Tx0XBMeDQKTEG2z/FTNXXW1caSmjMho9FKMLgY/OtDLMvRmIIIGkVCIET
GRW5tp6TLccIUnW8doXgirutYV5d2SP6/oFHfmhRSMfN6d0dFs4xGD0wfDOr/ii8
sS1T4A2XEAe+vE1aMbOKlDwRrTSzVHeoaeu1DR24puO2QOeteHIVMhTn70YyfKGl
WrgF8/7YDC708CNlnHSpS3Cd9MRV2eWfwdDOnIAwbe+UKBx+gImS9/v8EJ+uFRcx
J/W5ymZclHicpKhVtQQ1RoPdgZUbpv8VTZfKWpcbtNKWb2QzJvEbSZanFQvO1Ink
eSd/IJACGSV2dOL4fi3lsg407LBLM+e7oMTlqJJ3T9IGWcMM0mchosBfF4YLnmDR
0/I/CYnTaOB/oMdHNkuMsUmrVnYuZ9lNuivFbYC/jZyFppew5Tx0NJ0g6V6FTc6o
sPGEQnLnQo7gBsNXJsZ7hie4weEsq2dr7s926w0l5o5KEt9oYpFp/mvpflytUhKV
20FT/gK8xAQcdrxucI43huP+kjvy4x28fv/2qOIcmMDmq8RpRKxvfXzHG28mDtiD
ahGHGjdx+SYovwdELXMa1HG9v67gUvYgWT8pEB7Xky6PyGZMToVwwbUQLJWKTUAc
JNShfN2ob2YFMc45LOMqvAcrlTeXgj5UrSFbEvBbxgCuYGJLJ7mYTIBUnxXVdQLz
okencUUlgq1/mcHA94K0LeHV1Se/BI8/Uuth428JYQqvy9Rd+oi99QgRxxEsgO1I
J8o+7hvEoOey/JUPCcJtZibRTAiq+YL7OMHlXpb++1jgmSl6N217Q+sBUHt+/NbB
D4ijDy8HHc49KSr7SssMumd3QJ8IVLLHASM9ogb9mxJ3qN5rQcp4jrqnUqu9hX8d
IIeI7BJd1EoVEYNKTXiCgbVkAvR8JF7r+cmRWMr2BOxL/YWa5VAPLxXTWrOiueqY
nb0od3XG5QU+Nd0O8S/qMUT6MO1nwgAYyPs3dutiPnUt78ZvbIUjCfCR7pxOZ916
5kRsXXI92Hzz+qm96kDuFF3hnuKCG6W5OOff2GrtWkHqJzgMIZk1uIOdQcQ0w0Dd
2FuezxL6ilZrYdrdcIagR+3Hz6FfgPEgcMcGwd+ocTfGzpUUva9VlUsnVytwR114
Owd9KvyIVv2koySxz2r+EYR6aNHsNTTSuHIhEakoTteZmpYE6I8bGn5m7nKyv5vn
3rjwdJxFg6/FLOfmnmGp2Doxprwuc45qLhMLOH/xHpR+qCjmCwdu9qcP+hZwUCeh
tKX6GFCvHTOb5dD7L/rv+oPMHaI8cOA0IHM++HxZgdWY7MpC1v1AS0iYZoESpuZb
clkgUuoSAAuvDrE9kvi0d4w277Q8F/e65UGTkIkrg7phAqsHXHwjL/RnTSXW92I1
qsmEnNZGXH+G+qKXg8ToVZ+QtCe8xbvkZIOsHCYz1c/MMYpb9qcabYMUh2aedoxs
GyO6+Sm5SX2dCxLU/1tU9Ysn5J/ZJY9t+Knm830WbxaxPtbfQsEkpmvZ2gLvlaZm
4J4HaajLqVe+qrfgM5KEEKELWy7DSVwuWFOq7iR7vTos2/aa9N/uonoiL6ySAYOB
DWEmpagw5+K6W+Ja3u80egPUoHxb1zopdM8V/LLr0Tk9r705EMU1aJUcDtcjvsIb
EwgFSguUovgjzui0djj9fN3bnEDq+uVZ07y7bCISpz83GuNBfLrfUnhquFUNq5ZB
T7sFbr9z6C8weRWSX5KVMIoWzfUpYKY8B0F5XZGObLXW41bvVfJSZhM1rRVSINLU
AEoxQP23pCglCZ09pvSPw8AerSPFWQSER24fzm2iS3DZ18NbW0CD4aUA3mq9JNUO
odsi0Rs0Z7lvLV7rgp7ds5LIbLt1POmktzvQXx0RVw/LkV55y+8qt20TLv6SGlg9
5XZaWCoMMo5hLhGDp3JcMELd8/lDnSGXeI5evmurRdw7oKecI7DfGjXSPfxd120t
p74N92ZflilexJeEGCto4UnruHcrLHB5i6mUW7fjva9hDzzlL2rEV2QkwRIJu8BN
PMshbPGuPj8Qoqurq+1NMQn2fL3H54kwOQaK8VyBkj1SzcjJRTgjnptJDIg5M5lo
mjG5+Kd2jdBxUOyOc7VLk8D5V6srvW6ckdklRSyPuDSrR6PeCjdHss7Mwb6dlTtV
I9oysYv1aYAuqHWZ2FwBGGDz2u1iHQTHYcLPIrlfOXVNDjDuVsrkf6W83l546iyN
B/3kqaIAESvcalpEQg/wSK8GlSmGGmg1JM2VVWIg0SuGGYaFjV1TQE0UG6jh+az4
T9LL0I7H59xeRCSfDBOqDHPklkqwxLhezUT9dxFIfVbWjl7TPcj7k35yyDyQaw+0
tj6Ku6NlMCId3QdcPxeYitHUeWgBC/y8MfQljM7weSk59bCbauqHjqqnZC1jTsLn
nHgIatdJNwDqWOglO4p1g/G4A1QfYVS0V4JKni4bq6loneQZDBQvWy/LKbNvExAd
iOApc+RvKehSlRhkp7M/uL6NYmU5R2khcf8N/MYPruw0liA+ubdMma8knoyIH6KV
kkTWgbdazMeQGGBT0DhXsBnASqFfpCySQ+CyRhP+xxJ/Hy+lCWt21r3yjo8qVPUx
aDpJdcS5z//9qPm8P+JPLZUD317I3I6XK4HurF27gHo7cytJ5UbzDP2xe25OVojw
aStEh6RRgYUr2K4NIKRsanM174u3eWy45uym6FjWMCRCHJImjku0e561rYrof+qg
PcpCLuUPmq3I1aRAANz7m38WWKpcp4RJ4od2axWCRNL95e/bJW+8TiQlhah0Pxhg
Iq7XOQ/QqnUPmxc9mh5FZGYMtnJ4M6B514JWyyaEuC636kptUaA2nvV4WPRS3Mm4
EyMqGht/r5W6Xr2Vj4+fI+BB/7zWAF+mlWS3HSXQS3yQ3oL4Q90F8H13h++mWaoo
X0Zi9ahKROfB5vjEIHnb+u0EAjopKpnk0UAu/MxBwMpuX06vOMhpXY+RrUVVsIfE
WhctIhJhMPlGxu7lYoyErX/gP8f7408eG1Z8UH2o+Gy+2xAza0GZX3QT4MijtnJl
X3ud7dFjzmWMg7WT02DGNyIH0D5FfxAP90GyRa/mFF5OEZWW98ioR2nhnCqn9ZaD
1OJK1Yaeh7+wnJ3ssIO+dDTiC0GXbgY93sDZhsQYMCsM8apHXPi+vrkBEl8dwLm/
if2f056OGvFPkRlmHGeWA6eBjIXj7xhWO7Xc9EXQEWtCXEBpIzIWqOjotg1Bd0QL
J2YZMu6QThU+NtKAkhvM1sr6DxmquzVpenQ2wEyi/Zioy3GzXOK4u/mTDZzilhTh
lOLxEE9L6l75g93MXQL4xKXqI1BDl1GcLQFBDu+emHUvhg661FfI/62CcwHB6U1W
DqOez82Epg63mjJV10zKZDVIWJQQZUFhDzl6b/vL+CLUPDMkXszGE0d6Z8YpI4eq
+f7Fr+z1u2grq0rNrpPvfjLL9V7TpCmXa1ns6QZBUHFluGUOQPhzmQgyOwFpGMM1
+X19BkxkGgZ2TeTjC+5Y4Ay3ctyaYVJfhtH+KCjhijxpntzRt7akwOhCtrGYhFQY
0ve8Inzs6isTCUOvyTkBLg26FLlXrx5RjwApexWVQOOS64GiPAogspx3Zb1ipoAl
P1jdVWsLiucVHuREvsBxnJN8rY0FFMa4cADgY6SEBHrsg1t7Tt4fiAS22gi+NAgV
z5cUgM3O61B9ZIwIaFplxH9tyd4e9kuCDTyGyC4zaAEd+yW/lNtrnhL4Jx5i8a8V
4H3fd3JfrAKnN+w2um4q8C2BEs5jMvut+kcs7llfySX1LtKrtzgzw84hJ69JbtdL
epxMT4GdMOmO250Zgs4FmbWHI4zRWMi//i8LHQH/PkwK7SIynzmqcVwFpE22D6QU
EegzRnm4qVdsYgvlFdqWESfU+22rc7gqSmPYA9rbst+XjwZwHZMSMAj4QzJW9w+5
vT0I3LqcJ33Jb+MuyPL4EibUowtKZ5J+PyGyojURUlUXU3myT7KmtOLCPYJUiVZR
XZU3/vvGMA3gGt74R8LQu9QA8YQ9m9vFwZMiaMdAPzGOieYUrOCHujOfyT1CQcID
HdD7OazCeL4kk1Aj55xMVQIpFdmjTxf1LJ/p4eGpH/Zu3MCYAZZW2z8XwCZSgcq1
TffTft7btAVLrBnE6gqUKCOae7B5pCpRxOGKygfiStchFu035lB0zrjdevwoS0kO
vTaj0ezT6slMUSZ9ti15ZB2tWoRRTObEc2QNPk2dxsKQ9q6m0I0Q2oXcLTTIWAzr
leBkXO/XG+kwtGDeGVQCZxvCOgqsXZYRMWjIXRGqYoabkLXUTXyTJAFEUB7PXynm
MoVVm+l+GypL2lO4qZ8QvtWdCOseUsC5kRuVaROghkUPsZ+0oWduBL/4FksC0eQz
no1imFjpzV+J7rHofn+/UrqtT6jylN1tKkYKggPa+zCi/zaWk6htJ8AWFCOPUZnA
5uwDTVqd9j+FVybi74+beHp8x8IWTx5A3Ns9QGRuWaPag/KrhkUENoL/tU+O5xGq
+YVdDV4KjSCPAnoJEWW4zFgQ5gPw40tHgW29ewPTIDk1g9u5FKKSNv/W2LneQBsQ
l5CgdRyrdcfU/12gfwsMWlaxmVog96fztejUAN80ab917NrADyOPa4NJDLItVGL/
wCKOrFaPc5d/K3hioj/sKIaHErlEZ0GYHbejVLALNXqdjYbCvZ0fKUbwZ3NwOQi9
Ssk1VRBYsMJCF4xJKbiiBE5kwBt8dcfIt+MHkioZESo8z1BdkPvnp2K1GAHhoqvD
f3Ipjg5AyOlZMTaChZsC1bDthUCSI73dOfBLuvCVqlVlX328A48S5z3m6wz4i9+3
sYhT7Xyh8+MQP+qaRQtXEro40yvBmarrOyAvoTVPLjC8jFx3k6ap6vlqhIEbxgjt
6SPEYKmJGqxCf3dKjWiUGOIBT3f13nEvPhHJQGPy5fcZxNERkZW9bawtio7N5dUO
2QnnyWA/N377E2XQ/k7HD2NVFaH8xVjQGf3fcXS4+lCwPp9LFIlKf9dmBR8kJRQK
3x5w9JwtXyqWOTO+e06MMUtA12unHH1QGVqVrhL5wGko2PVH22hb8V4lxpMZR5ej
ZBL7G7orOjFBw3TvAgd7nPohdZuTjcrmGLyJG3fOVhiUZPuRzOJE8Y2EHcNAc+Or
oobo/if9GDdnErvXhTMfYf4I7qpLO02s/isqUteUHp9SaUQqfiuMwR1w6L1rBKTt
sh0LiaLq063DGXISaFS//KBNVeP39fnpCI+hSPBAKD+p0+G+VuDn2mT0f9zFXiSg
UacV1F+OsdNhYOlqfbiijGAm3+rlQ0P3WDMrxFHhz71WHjvuZNgvb7s1p+6uMt4f
wT2jF8+UkBS+9I+fRjEUApEzCZ8zo9SuaPJubNl6J/DIXzslSuvtz+wu18OD8IqE
M/VfYeorNCeDg6YIjxYa0O/wYxfDYcaX9KcGtmUuEIA53sYrmsZ204GjmyWHlM45
iJOE+O88QC9gJz0AGLldtEah9yPzUG64aht0e0po23RuNrb+bCCffUCtfulC2jj1
IbQ0mCIF7W0+aBvnuIK43yR/HBGVTeGs4IViAzq24q2h1ysjMcOYlXGoHIJ5dRp9
sUYQCx+vjsDO1tohEimfrAmNO4mnOpHeBY+zaWzQ/l0JDl8E2TwE81Sy20ASrI2r
eBZbj/b9ES3Opbi90M/vZTdkEpYV5YO9kyaj/QnhW/wVmNLSho2y3GhUDxqzmvnL
iH0jPiui+XMBGh/rvNCRb/a2T/euZISjn4/8KAi3RwD2fro9a0jL8fPpFPjx+F/j
5mNthbszeLya4bZiWlKzlvIISorG6Cr+k6nCDrh47bvlMsmUSIt59/IqvBNeNW91
xve3CMFfiHajCJ+TnK3slUYpAYEp2ydQlfMkm4ZZHzXMjpm0nVy1e4PnddPlVX3U
Ds2qmXTb/RarM2UI9YwJTtrwyUeoGHlJBOTpOLak4cdCzBGaXwub/sNwo0lXKRU6
yYQKe7p3Ix7c8x67WHmcFAfbVAiJl5T7WJcqs3G96JH6p7eIb8LnDzwF+xO9jodE
HdwnRPbBnW9Gu0sRUUYwdd1Bu19hWfNQRAGeZ13hR9fO4etNXzpvE5QXKNKdtrAt
HQerJ1+izikfYXsIHosrE6N+JW50J3pgB00U7qQU4abab9uLR1OWklsRdhuT7VJ0
+Dsz/a9MSTe0Tye26CHv2hRd24aMW3lZp7HiZi6tWrym4+sJiLGvkQ6aKHxAp6aN
1OSM7LPVlXFCpvlj27Y9s+cU3T5y1QqaSwAcciR6XIcrum5alqSTpOmqr96iJHyA
pS6jyCuRzDsiK/RlGu+Zc6jdfqArH8UuIKoffl9N8fRU+5OyqNUkIC33k1PAKmEQ
7O/l5RnlDJwyHPnXPy8wKs+CifGvt6d3hl+afBMJ4oQI06LEHsCC0bk2e3FW87AK
/4JJctwwjNtHRqMvubZJYaTcqnDaM03OdC240c2NufqT1U4ZadCAlCyBxw5j8eRk
wKy1nfy82DyM6+4+C3sfLIlSJWv3iLgjc8OA5Jmv46xomfppI22jViPhSKNqpRIr
PHBuZdpuhTgyYI4diqU3BBL0eqdaKYn3s5vpaTuLrwXx/avnpJ1PRVZAAtnrrMye
tiW+l8I6vDSYjdDLVN0bH0593yN/9H/nYOLpA49E0/U3I00QoK0z8/NC82DqHL00
X/5aCRJnPgsHEmYDqu+iBZn0gBEM6XFW6smVYoxcH80mSvcMyYH4YB1yoOsPwVSd
8VnkLBf3uAaCE9wcvrZI+gXSFOBA9qIauWmO/OtFjo2TD5AtmdyNBebps0taY2S2
HrypX4zNz2OAt/j/PDJifbsnqHQQMKnLoCPa9WrRBeCOttQOCuRM4KhLrpn+d7l/
hoIlFHSYEqBvSdGVxFBnTWpAqoMN4gOdXX6syqdwwXrefHYhmoW/fUMOkSVokssm
4Q04meIoow1/8MShTsPGOxX3Ib/dEeMqgZuhiWmDzVYKA1zhlANXH6RwHmcxG+cR
TJRVK5lPhKl8M9qMMfww8JnLfFcEjUJnzT3zi9PSVQGaU52UaT42FtSyYSfyacQ8
F/jpJTc07NYQBbc8Ph+tYo1EY9g1TJbnIrdvzVr5s8SkO0a7TbbeJ1PdM1atqEZx
gp2roCeK3iWCYAGxzPfAvYyAFunqwTbtetB7Inv/qsBdnbQG4QyG3QFOFBEVkhxO
aHL1ixfORUHOdtpcmoMP5RDtL3f1b4069kTnlF2pmOyRlntyNJvz2cFu9LdhpVxS
nzW1Qzm8G4pRR8elIqTKqdVNLnp74TZpdQ/nSsqzropYCP24QZM+vSg7+beaWTy+
tl/OyseBR8BNXSUsVy3+hoIybNlE2zHSL7qHv/Ilm95jWrdzKA0HzPar2AIf3ksw
rGhDR17Nd2UEhaNpW/KYq/0IvIRi2dHc5/x8RPws+fO/5UTJUo+rdjTrr6hBE8nD
7Qeo6GhQBNASBdwz1gIt3JikGYqIp6oi+VN3tLnTRyz6dpChNOLyiTXz3wvg11kK
YbFG16fpw5XUsad74VqEduye23KS2hq6GPqaR6jCZSeMBXLVaK0kcmnnsow8cRsN
mrJ21Tmzao20S7edd6QdaW2AEw+A27UTU7Zvo5+ne+0t4JJ0Nr1mOxjKs5L8PNTI
fpptHnY1lkIlGy2FCC4o9MfnpQYi/0E7nnVXrCcxjRCBDs1hQj1GUsg/liXRXNjq
EUrv2xNZdR4dSUNIJiVgrKh1ZPk9JNCrd0rlYRxlF8MFGfmn+M1CmUz5SEjGP3wc
MyFGYPIDbSPz/lcEyycfucNc3kiViGO9uQZ6BsDrcm911b6SQTD5b9kb/NUbGWUc
QcQDqQD94DZcqOo5zgZ6I2dtk8nx7+bHDHC6dQ34u4c4maQDcCHU97t9xg1dENlw
1JXo3uATe/YTDMdCnq2N82P7d+sEICRH0Yce/uTh1GSKwpuuJfB6N6TzuMbwm5ud
di57b2M7n3b84f9/GDLmqxf1WVP8619yXCWMj8ySLFQRq9gCTI3yrGg4IduDLvNX
MmXnnkg50E5D3yCYb/vmcH4XpINgRRXmcVJ0kDulmdRDQNAoBUlRwgEJCPhEryP4
PWkD4yP5H7wJvq8QUfMhxmWC2jHZRnJya5D1QJykieMD7/jlHL21z+OtLQCQfxzA
YdV/r5sl1d4UkLq9I6YiB7387FTiRCB00Bc2uQhVlEuiF2qyxiSFmujptctxgklb
y7XkL9Tf8Cs7y4uIygTkae2CYYTAtAwYXx6blUHF0ewtejnISbti7uGEOH+GgPty
DzWuU7zPFfm2A+egnIw+4R0DgGeiyiVFwgtDJXg85SmoFYNoXWPe8PdvzcA0ZFVS
CnYv7ga+zd8sqXLk+Vwt4/Qet/Z43HGdtW1VSmU2v466XVWSNAblnSM7DUtuaZj1
cuzpc8PTuAl8n3FWbZ6DbhBrmogYar/fh9KZJ1csNBKgfPNgJRVy48XVJneQpTRT
rkZVMIwjC9Nb76jWyM+YWIu+DZfsjegCK3D4xRLcs3LopuTiEmo65ivt0r7zCjOn
i4l949FbCSVpMYf/WdzszJXkHQpQB1Ks+YRyAo+889tG188n82Pji7jAFvsJXiei
4vvnjAnfsrSlkNSbAC7e7+5uA0ttz6TtPbSd3sRFkY0bbzAci99sdWEhTVGSm1uX
60ifQNEGemGCZ/aOnJ772kG6aYtaudsBmgJDV9fyy5+fH8Dyt4OHOutJIMOgKLpL
iEAy/O2VmuBfAUNFVFZzIn/lqF5RbVhkAMTVhAQKHzQBtahuiY3nARsa5ouarLeR
Z1vUCkwU2lplbtksP/E4rPHBTXxy1sL3q1ELlwvo2FTMEI7UP+q5wT8/E+vXzxRy
w89QjTlnDLRXDtAYAeYHnivplksQRtzlXARVKR9PilmftuiK1Z4wjnkW+Vkf1KeQ
YOssm/T+l0t/KQaQSe1PGgke/QlFoPLZXceAXKpQxiGtExtZskipBKmv2bPS9qbF
dJD2nXB6usAyg3WGlalFhO8IMziWSLPPtg4fkLo1mZVll9zmQhjo0RdKAgQ8Q/lC
Yly9/oFM3Oc/o2U3i0cXdWb5u10ogsuRxmItj+fdrkIaCPhDB2kCpSxmEzyy31Xg
YAOCDKmWXHmjx/mgTXGKHc2JoxGMI3iz3/gw08jC1pXGIZevv8wi+U8sN+W0Ar29
uYHYVlNCATTXsv+HCbtRZHroDTma5ke2aZsXWtkEaQyogIKxSumc4QKC52iU6n62
iQgo0FOvPwZeKWvJwIEgSNkqro/ys+5YZKr9EcPnsIM+DKcIAjM3Y/VyHuLLSKej
RO8w05duQoBFfxBVhTkU06QLIqUN0YGkUzImcIzMDEoej9RyiWCuQFgCE/zr39Ed
wGnvsRyFPez2b5gWyanT5jOpfd5XjVzHSpzbTBPPYUwpGwQas0zYJYbkzLArO37B
x9pFX/pmBDm/4dAhZKzi+yqUwfgmT/sa+MN7DQ9kGEYm+leYHnwZP9NcLjDGjoRl
D3QOJujkUulmFkoN3SHJstd2ogvWOe9G5mcSHx4kokiwLnN+QQIjZ/Nmhbn1WEts
J/Hc7STFi4gvkFgy83Jitc7V5ebrnpD32ENLj7lmZfK2Loggb8T53ck9dp4NxG5E
5VmwKxAZDdysU++QJuRnjmdlZ2hjQs1Q5yuRb2udGHC/S9dToERajDZ7Jj6NAwg3
ael65Nb4dX+iwP8yYEaIGgf4Dj9PbrRYplhW36LxCof8U1u3oHsuaCd7VUcM2nPi
tBH3Ky5ZhGw8vEv/2TyHxiuu3P5X0XQcO+8nOJAEx3RMwPaVN+ixp9pm6xewWZ9r
ReEOm2NiNbtIn5n2kISUCmf1rvf4jHA8QLPOp6Il8eaADr3Xy20V3uXKcNuCuiCr
vJz1BVhsAq6Mpw3vW3glYxVXPmi7Qxz+hkAa8ovjZ1e/WlJ8UArb5Pm7KiYuvGL9
oFWnR9+H3X7NegY8JCVzzttrO8GMYmO4opmtZ4N+teavC8cvAyJl0thei50KUmYn
jGKXDxOoNPUo4hLUf9Q+cfOUtVWXJRI2IjDM5LBwdTayEKs8+dZKNKxsE7OCINUF
aNRswW4fx16e4HvD4LS6V15MnJX476WbIkVuLtkjrak8rQh0L5BlLrzZ1Bcbv6VA
lzJMx/1/8Db6+xqJBdvBX5V6jzwerImcwGvRRdajkHgKwnxw5hkgv6DhBEZRBq+E
JzabMgw/YZgwByK6782bEVj4j40HLr+f7hd07ohl1tpAAnlNHX+VbFuEHNBxruvI
mcFKHbVP3bFWf2+PJU4X2XL+bePYvS7iqUAPop2gaL3MHBW1ex+q+bbH5t1KUUrk
+0ItKJSNDrobJhXgVaE0XkTDa0s7uSxOHTt3v7d5JwAZOJaPZ0LU5iXAH+eCM+pi
DujsTfPVN7KR9uBfOHL1O16ndM2cNA0Dn3OGD5NSF3rcm4bHciawUBnXTeCvi25w
wttb1CjMy1i30BrZGsQh3C5hXExl5KbEQzpJ2r7Dno0p+JzfHhMk1PeOUjU85dY7
T5yidEfvNlRMNvjNIwqiI5DyZRPazefFk7bGIw9TMC9QwIHD9ONxwXaWLTqWE0Ic
/AJZjUIOBC0agSzOAgtOxeV/sSMvqnFMgkoz0bE4UkHeSzpQ7y/Dw8SpUbF88Djh
04LQ5gXETLCUulLoag5ZzLukmBEMeLfT1U9Yz0KWciZsPxeHw777/m0pgTLsy0Jd
EHIwNQnEmcxZVhueiPvBeTu/AoBtN7rBSol9btH51d09mRMwqc8n/PJ1wTEjzpKi
oUWJ14nVoEIr0GI/c67HzA==

`pragma protect end_protected
