// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
Rkt8CGkOd7kSMutAt9iy2560Vao5BqscgF++tSTqvcrfemfEoH652QtXR+LvZW/56uICcrjhm1TW
DYPaJtfyxKQ9WW3Qt/UihEgWyQeu2zW2kTwhhudvWXVgS4sLIKfH4GneSxEVlM/JBiJO7OiR795S
0DDQbjqJjkwW2NVnrUByTMm400QV5h30BLSBCO92A3vzi08hL8JoaGAJ3j6TsQITi1NipgIMyd90
/gzuHgFjEEcZVNg46PG6+wb5CYkJrYZuzGrsrF3eHK/9qJfTneF5FK8hMWqqQqP5QfA2JAfJZhNK
F6X/jv7D4/IvxVZcNiO95kQ6MKj3YqfkbFrtYg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 44848)
dMYBjNaTU81RKxDbmhg0b4R+xkYMI6DihS40oOu/ZyqJOMtdVqV1RWS5GmaeW7pfnk3SBBqc5DbW
mUY2PEXQVU7IBepTdtUOmMCw/Y54fg49289B32/Ueon8oTu44pC5qvGFXkuTZB5C7GKRzAnIzUQy
AbUYGpx+x0je0Saj6ugUfYA4QxLUlolD7J9v8MbWuvjAw/mjYw8d7kDsxBqnFd8YvP1KOXKIFY4V
HbVYbQJJymAGRM13Feb780OvhoTsG5CvdXpPz8tGmIiJ+aKbFjmVMxwKle3p+RSKmBUORHFRXuFC
aeFmkf47Ath1wlXrSHM/eLB6EedvT5M3yczyuxooziqU+BaPhoYOa+F1TkGlqJljMemVNgYn0sLD
jel3dMEkyyduyWQOA72ChA9Pje8ZQr/982QVqQmtwVCKjeMbtXxyQ2K0DYvXtTZXIOjmXXawKF7j
Y5yR/k3hRlfkeaUN7C3AoBFsZ+unEraJIksibmdN+Pi29pTMiY3CZznirl1834MOwATbpy/Z5Srz
D1/aD0H3wG+SDzDIW1yM5DrrB5amNH/An+7PwqrhVXoRr6uchPabYSzjrBcx/HLxb5hAmOW1bWA0
7kJczcCiHE/WxnUNudWH4u0pqmAufKvoGultnreIDJAtD/9uw69KJiB254xtmcw4rWcuQ30NtMFs
ZpcIN1PEwhJWvSGbecX+l/BX/kN6FLkJHQKGN9XVGRv/knCUDOskPthHJNNTUYMB9sqP7UZa3yvh
376mIqFu9gTTZuR/3VB1QulPHlLXYeqGkkeG6IfYSKBlwebZX7AO4F2Q5JHx0E0FFPF9fHFUFfSo
g5eA5YSR+OhB0NenxD0V1q1Sf1VkBN4fokVsfG9nH6iZ0gcLbQFPeHWRJlwQcus+hde63e8Z1BA+
r1AYluznfwgqlgHMVQ2kqiojJRjI/fjsPjJSI/e4PKjDEJeEXL8minyglwXm9i7qJ7TnYycMAQ88
qLIayTVNQf/kJmZI/XSvidZU3vOKK7uWETdFUC8jFuMl8m927LnLvXhhz4+3W+2ZZlKe8QYJeL1G
m46sReb46fiLuIZsmhzxkUjztCQCHpYFLMCZ6x4QybJ+nntGlzcJAHCEjSnlRUXc9UwV4TqxxKDD
UshcN2AHqsBTB1uR3n2SMFcTVf82/pB/G1LAK11uZ9kNMx3Mlhn1UM7vY+AHm4wBOWZTiSYmvjxT
Mf6tySMOZmgz33P2qac1p7A7VVvjU3+xdmoUnMi77Kx4Rb1Frbif/7IDyIOCpGvE0Tbeug+Cjwha
MH+UwGy3kckKm5cqPduJrJvmdAkjx/X+2JmbJb6Ksm9VZZMnHmsxGi+DLvnGNfhcxdvrwX9hgUDh
pkOrxgJ4tf41Wgg2KhyWopfY7mm30k4zYlq5Jqxjk98XOICyhZLhtWNbVunx3/eREgrf5g2x+opD
I6yvThnBFqAIgewuDkho3kHOIWPRD4lW52zi9r9VTwUoUpklbGcAPfFLXcN7V3KNKTOT1DmIL0rh
IgENGGS4EZT4yihyoIlvlonxK8c+lFHQsfwzApM2gxLcrmd1qWh8mBsu6pdhkNvQCxeWvdKxqMf7
3rcaudvAe3TuimLARKycYbqJklNBJDRHw264rkQMSJcRRjmOVyiI/MvJF7nl1dOOL8ucZQQSyXd+
RZ11PB9OgmI2qpDVoOwo7OQK/p5Rg3guKbOg0W/4Fx6a0mS+TXs5TErlmxrW6CfaI6iZtmHFxVVe
Q4nMWdNgNd2CfXImeWldHXCl2S6z3RNncA0KvsKEDrvNR+eOBeOZEVgNvWsiwSJurZTE8H3Wmmm5
S0FmX13JC4NfDyMrX9t+om6DfdQuWTctkfEG42+6Ps2kdJfCcJ5zEQyO1ieu7wwBrSe3dWxSxZqO
kDIlmvrgig1JK37FOQfvYq0TmITlFSV+RMoAugtlKd7eoRS4ia841HW0k8JSLh7LkLvOodI4kKnh
arNNEF6m0nfIwII4SgBc8ar8l4NAS0EI5sPzG1mwpH6kzhZoqestZLDwn2uI5BbRlIFkOZZD58ll
WowYEjrpsJnm/gnZc+qhEBC1BBcce5x1JgNZrAUlQpzwNJSpuZOXEgH2s4PMSP9f/XFe13zY6/2f
JE6SnIqeudXVeNMgC6vK3FC0FKcMffJ+KRD+5Wr9zltrpV7OV5UhJisDwhFaqKdn4QTqvBUJwy+a
tzLQX4ZnPv/IUJezoYCiQzvtKxhH6X2xDepjpARJ9ttE/+MoQtMoKz6ExM08kkP7Vhe3rmiP9wF8
9qEnvJCE03Y9p1R6ewcBVfYWeWwpAS8icFGbSQl+YGIEJSAPdJV6fBkssAJTvwcQI8AYh3uituQX
nf5sU0L5QfZGJSgrQTXI42td9XcbnXqYWDDaxez5/3k3T7PyOcdK2I48T3cmtDE5oDzVzAxHHTKi
JF+seo+1vMDc4Dj0KS6LnaLEtyLhni5e+5Ho5P5hXJW4UCmVYyPFUJS2IXhk7GvY1nzXEKOosent
cWEeLbEQSnhaFWDcW3i/nWG+QTRB5Cpmb5Lg3SIHF7E12svoz0G0VXLaBZoxz12Y50T1y0flsnZ/
rcSmTuCNQ2IIzRjxRzOlOJsjtdQxvOdPQwClkSifZXm9mPLm681dsPe0QuvSt8FK7bJGFg+M2sui
GVxlr24WFgmMPbVuYIsRuZvL51Qai6QapgaGpbhzL7ijcmXHNfakwQ38sAjK5SUFg/kmZJ1eqgGV
MpP6EPC3sdE6dIUk5XMriaDpazFI+0qTgKJWvJ8xnkwh0Glf8ShD7W5bJy7Ym3VsUu2PeVmD0BAd
9A1TzcnsDSFqYFOKLLS3Jt3MKScLLPBMAV2ZYctaRcMvbQRcfhWOc1JQtKo19mQdwXjQtLFWnvcp
tWEZAZaQbxfAugcBsY+qA2JpKWVZsYnIjUDGTe1USpVEBAaiIgbRMhULBN2JqfrIXrSC+FVfUe85
J8pk0yOwWTh1VNpdEelmrHQRHjEQpW4S+R2NoTpCd9pPj1JkOzn9ANirJwiV9giwnrFgx/zYQYON
gEnC8PiimzeKozjK0aKo0fvYybZ6ye5TkmAwEZ059AyQy088hdrCHBwPll8rkb2qgkQQ9GmZyQhl
vZ5e3UDUXsqnREgPTzytu5ihXK5xcmoJ2UBENw/5yJBteOO+gbvZc1fo2YhGG28J8pmhlPfq9bCd
0Rtv0UdiWhGIG/c7KPrkILb9yzYia4UYrs4L/HOxaBPyHX4CfhzhvN8OngdP+KxJIe023iSN1UPT
y11mBgJDAtH5E7AruhDuHxWCK2qwCsUNNxGuScz/L6e0OOOiLPNz3pjaMtJqzbgwCTu7rFXpLK8Y
vdAdrVKRxr6TE6SYHeWURJcxvZp2ABOYTr20MtNw+oapNARFkhxgC9IwhiLzOe83n2fG0SlQvQ7r
AsjewOhHaZTtQyiYksyPf41YvHXQza3AcbEu+P38SllaUYc1H1NhJPXa+ht16XO6i1F7a7mjwElD
PoQgGdAlAdyWen9gJdMPAsBMWoc+nszIPTncaHc4vv18VhL53qZnOY+zaHiapVgi8xnv/UkaxkwC
e4OsowAxj6RqneCjFhLWo9g7g2i1tmhYnK4a33i5ue4zFKbU+EFgAikiRn6q6devJ6cKoAocDDaU
v812J0l2xxH0J+VvIyciygCdpGaDp03dfxk5xpAjvB6Eq1wAgCoseS1PVchZZF7n/c/oMc63qBxP
l4eKM5qoSVvwqf3PNf56fRJJRfB/EvUwGwkGDiepk2hNWpOC0YR6AjPm0vW1G8mZnaJAbAB7kSnZ
QDJsGDEypebOSP5mnm0yNP0X3MbRkhss3FkMNtw/eI/XWEgDIF3fvMUGp1aZtvXYN9SyI3G2AW/w
+RN8aQVOV83UeEH+syXirel96heIn8294tgj6W0wxmJoggjsapM/TpppnkwtIiBB49ssYayH7SIt
Lnbb8NIlOjYvubu/uHr9R4f+tdXs3imDDjASCWfQ+H1e9+MtFY3TjSsR5eY8T+7uGdOt4lPbHwCk
xcdAE5vJHvOAxr4bGOT5BrRqLE1fcXVOOQWBqMCupNv7M21l1sKpFw28dsp3htSCV2fH9lEoZyFo
GrAQolAlw0BBuFAda3Ek2YmgJDCfV5140VQk3miKbFokvbE7kCNJLFMEsfnajMcyTfIFmio9QyAC
R9yCzAIqD7mIL5AX8UUBQP/E4FrwEw3iCNGKBLRa5QvEUV/n822VPqMFLlrjYwPXsIGcI3G4mIxt
BFWEld0JSEXreIXCIQFpLDhvidJxl1pCIVXeqHg0rrOXTO+6++KwD0MFeCk7n04GpDesPORY9ezN
yeEFxOHyMxwC0vWKHlI8zEJCuWmvlsLyq2Oip+pZ7N2is1teIjHdUfGbkSQqO/2OhE0oFh3jRSEF
/eHJq61j0Pq3x0cx+Fz4Ij1gHmkjzq0xXOnXNds0soH9WLfavY1XMgBlBbbIQsbIZCJRwt6fz5LS
P41KvPuda1U4+rS/29oUUejWjD4Mom32hNZoOAqzN8FfjEWRnJkROoChFsskz59UM+vFO1DL5VgV
sCG4+nbKGdD1TVAByrVHica5PvxR5J9aJUDfatBPyEehWzl3wj5ef2Of5HqcdRAM2ZOniTkr1tSG
NtFR98QiG26A1vk4hpJZYy0Pb/8YUN7EBARQs8ltVfwfRT1uFEhWqjurUoHtyu9udUm6PBB/nPu+
FgFM9ale+s78/lAAiBqomdS942KSDKNRvMIcZS5AMAD7xL2yNvAnCdez3vnKwSPdwZtaRQEifit8
zXokSTegpzveMTigEDzbcyXjluT4wXwTD9k6SG6UV1qiTxA95SWFdZwkd/pRC9rqvvU3TPEQxP2Q
ccuXmV1xd9WbTLab7//tWalhuzHVCGnu3De+Q/wNtM8EzPUAcitH/67cLiu437ANfKmJAD1JU094
DOt+MzqoRRBI8MTtIv17oio6eF3OvhKi5W88rUxvwjwpKsvcVjzFpDbF0wKBgQI/L/ckNJ21n/iQ
Cm2UHWHm0jgBolbcAiImcOtwr0SFexdkH6XjRfl1XZTRfYI0DpV/KjiyKWrU0+mXKex7nXmUOMIC
fTjOeJYBH8HoNjLnYo1vsZQ69cpRc2OzJ9oY1UWdoprrLs6Qerhy6sOpUbNQbF5BxHjpp9Xb1uoy
t9Z3LnUV/fDbj4ZQTEJOoalm6W6vSYizHxdqNoJPbeUNVfJRnRxXfNVskdMl+mFTqpmgfXs7ZYvk
zdl+kdztiNJVYanPdv5SxR/LTzURXKpVnUR7OLCT4yNQboKrDGNqj4/8wV31Xqz2tEl1vqr+p3IN
1xQTqVtaUvI7uBmNjk2zmRAnwSDEfOMK/QEqcHYw2yAB5OieRa+MwJBMobHmFgMlbCtVPX39PZju
93M+Et1lt7WzkZFWrh5P4+V92qLFJGdfuw0nv29F2lcFHupxP1b1Ocphi9iivvKqoMz4fiImksIj
0Na0jl0QQPqbG24qD+6G2NoHhzZhDjAuscSuv82Sdo1yAmwyO/EcUEzEONXN/yh/Uz4q9Un/AXWx
CJEsPixxOIkVoii4pY86cvWkUyZW+EHnGLIuqF02vT6SnjIcHPxKEMcnLgOUQ7xBA/gCiFuuF/D0
663P5NxsIIT8oRANfFx+hPUqFmvG2SGjqXh/7TDk6dJ/0C/y3KK3UOXWLJg4u8lTL5eiyxNGT9So
o5h9d3HbjFnSIDDEzq3UWxB7aD75k886ijxAOGQ6dKpwMESbKQLvdewsk1r0LUX5T/+TvrVphYdX
HAup45enisUkpg591OHud6ScIAYNR39+VFxplD8v/p8NOR2jGAoNs2bxknaP7evwmHiZHkidsrfW
YdGBtfPF0Jsk8VJBxxb0bJe38lYwi3BIefCQkW3weJfXf+iMYhZLz1AM4zGCXjHkUIxJ2Ro+IRML
9NpcD6T8n5hnp+8Zl42FhyYF6o+yP/L3lcb1a2drmp4sWkoQcudmEq5YWOgmO6tr72iUWFuvjJ2l
/sfU0fMbfXApiuTWmGfuTR9/ChEBPleYVIytUdPxg2wumVNI3TmgvdaIzqE6T5F0vSzGc5cwMUp+
a/CsSb6qi16IMy9D4r6SruNZEvPqJKuGsEZTONerYX4J64+lOi1abtWGK7ZWz9wq5+yZmCKDVpoL
uiHTZ3KJ2ZLT9fbk64TRLLOi/wsnsh3SOUB6mgr6X+IQb0NNmGJc3GaeIU+1ZSYQoFxf8Usa7kVC
xIC6nr3L1DTiohwJTzfDiPNaZV/Sgder/RBDsVmB+pzTg2jwv+cbyf20YJU3+QGghvWDM71Qy1gn
Jp3OAkTluqC7Ed8gX8xFSRYG7kZvCZtqBbedEcKG9dzfVAEte0SRL8OPNua+KrU5zsY7hDpGTjOy
LdH+O4hVXCCMjUC2/7cNKpYyPC4CeUKKGerCdoZXd6JL0wm1RyngxDrvEW32apXjFJTsz+r8f3In
/waOyUa/cJQVa3ySY5YZeC3cCwJygzpVI4tqy0+BI4iO+8uF59EUv5v5V8D4jPanVZoz8+K9JqSa
5D4f3iVPNhBZNGyTCn87Jt6f2DBG1ES3YUlmQkOTE324ekvjeLa49s2sqMgHMPeHM7EYzXuz7655
/Xd+ykMLvR6zdjfPuxGmcsxxnWaJGs0FVKZ91xmpUVV2wBNwDZW9pkpEXHa4n2Emm3mwkz+b8KQm
KVqH4luMJh7ssZzJjtT6HP9S5Hnww1fzxL4mR8jY9MN/iFvD/mwf3bLaUDcrixuCTqDRd8vmSOLu
DvJIsY/PlWSq64JjEI4JghBMD10GRyFWbuB0mFUQ6pmrjfuVJtxTem1yfwQCSuyhlJEWcI7CuH1e
TLsZJd9/kP1OgHgKXX3JwYg2+l6gduhjn4+frRpkd71IsIbEk6VsQfzvhusPhA8EhAne5HrzKqeQ
7/uet63JRkx1FVKR4GhcfhdlxSGPQDp9UCuZK3v+AeG270wnlLDqeF8Q93JFMhbiYz96KoAqdJqP
i6TaJDlqyPAE6Uc2Xp2eSfZSr/Xq7yV+yy5kyRYtPa34mrsypndqdb+0Vxxe2X0ljWBGwK7LRR5w
ONPvqrdb0Uq1KcZeYnEof/0iQTg5zEFEUI9ArGj5fqNbuNKG7uOHl2ZKuiTiQRHbd2Mb+1GnRVsi
C1TNqoYn5DE2yxOgbRWq0t5d2SEQ6472wx2xXd6NwAeOSEJfbygY5hztD4yK8iMlumONfX5oZ5R+
dNHGlWBKLGO61GxK3ExxfAZwSQ4umT+oB9wexlAiNWgYQufxN/aIlQDcPcUTWQqsNNxtvlizeqyX
YD3bGASPyRWIcXMFLnulhGIgPelwvuHEKrPQPeFviOmB1iLr6WOMgqleZ5Z/WmEg+TN3HGPD3i7K
Rs9afrq+LDfSY2sXfw0cX/gvH/sWuGcwUqQTrJvMKAAsWAtYU2vskyRLLmLQu8qBNYqfgKoLGQjC
UXnEeLv9/tK2CrnehrPkJhhDAfYiAtIS41cOMG+uxqpLXWmbNRXrRGrt1NtGTIhdQWJj/z7McBiF
4FsOvckcQvn7pZ9mf62/jKFDgnBO8VApat+Y/Z3B2jIqDYa7apmV10E0Omrim8X6K7CIladsilmd
+/qOcFiBbmv3oywkcgbOFsL+OfP+ABYaumlaryFRHbO1Dx09RZix/w4ckN+7xAYalpHaZSrIQxNm
ff2H2dVw9WStUqK+4jcgc+ulX7bdtnlG1Xw1n+CoM0xF8vUBJiLFbFX77h+Qb3YOlXpn/N49pjLw
teXQHpZpHEhUYNNnBtVu0zIfpeaYXroyFDDejt2yC4L4/zcPVIZC23Np2vc/7Gqvv6knvzacJMeg
K376Z5jcBlys5Gtx2tausBfoh8aPbbQqM2wFapOngJPxum3Y7OjKHxfRwmuBGPtviHNVuRSpDY/W
VqqhL3TLJscUe965yxwRbllEiyTXz2SNBtUKfgQAC4oOQFa6s+whF/IEpHpdk3Mne53pGeXhJpp7
L6n6qR30USu4wAwsFO6R64m6TNllc/tQ480UC9YYhln/qrcvpG9StE7H5Qi1riE44z+H/T/W91Ed
QhMeyDtkxmEcuSlAytKGYNv0w71CKlrffVFPA92u5nFdldqml2I23OF8+XKDNu1HHa0ELqDhzdyc
DtAGhzAD0i+o0/NkYcu0URg7xoJjvAVew7HJGICfjzzIGzjowz4xp+K+/LpXy750WfZO9u3FWH6f
GNypI+SeAI2/kt7dwAXFSqA6SUho4P3kjbdyTbixo4n9dt+CmsUe67cLHkzsDJzJXRJRUAAkYSYt
JgMSWAtFOlRemBGlTfJLtChcq9laeAjLgzlQlmNe8jZtbFxaqEEgYiBjOKks9nvm6EYNjluXnL05
PDHdG9lv0DtFKO4Pe344Hj1Crv62H7xA14JxGVjb1y3xJuGOk+DtIesUtu/8HPNm2vuQL2kpQbBy
s6yzUqQwfuN1Zv3dKeajQk0B6AzO+3pooJcZos2ZYcuQvpb+xRf+3SRJQi2oeM8G3C0LqMurOVx2
DASYyRp0IP5u23IHDFI5NHMLNcjMNUbaWpFe+m23xyXBJiaciUwWao/Pj+1qrM2RsJjs+R9xOmxF
sRdBAGI4sMjacZyzNk0fUN7ugXghNACQegG8mujBNX0KWZfdrJ0YwD3kChssVnT+zRtSz8igDItg
namCaEn6MKq0nvTRmT12FYifMupGNrxULn2zUioJkEQu612PgZrPauVNgyZfn+PISkpOqZKHvhh4
5EKZSQ+zmSEDp5fYbCsXoEa//UniLr7MJWn3ZP6rmRUyp/QdffNn69bqUlM0/EnA028ccyi5NzB0
ADRHpe6l0jx5nLgHUhFLXzqVL6f/uK74rq4LQci/d4vuIndVlZkwXehLOXHv2S8NjvICtYV/0zeN
/QHp1mFkRJFRq5XMawHJQEZq9UsdOhjFVdEr+bXBTI4e2QRuxATI7UScSu5ywbmCq3P9Yo8iiSPW
AmTh4PK76wjWg8GPtEtldm6Ymwf/T43JvmHHoj7Tcl3Z06f6hIWAFcgw9qIZMn13wR+PfPThlmCv
cL/5PK5hIfYzC/axeXyUzDpYwHygR1XZJCF6dKYbj+eVvfyhcENm2w3LhrUzMOL7RWVUJjJhSftO
LcFeddcs7GaxXdT0T6RbF6m+3nsmB0BQQuMUeksd2QEWRJ3rTHSLBT0RTDknUxVfu2I5PCRyhyMH
gBQApv6s5ccamIPZ7XYTVceP29pee0ds3ATZcfyBxOM4INlL8XDtxGETVJMkrexqWZ4ilXx2iprM
CcM7TuGIQHoGMGdYLwTMP80i9AWKD3t+C2lnFWS3GOdWrMTewGmIoo4uZxmmPeOTannf38l3jsYZ
tbHMklYQVb01h7kGa9WATWACyx9WREssKMREtLvl+WdqV8vX48wVQTMjj+x8rcQIG6Bk1aG+AIAr
wov6K6S+hE8YLrKIM+THN11e86Y5NrAKQxx7Cd6PZFKbxATpJSMZKWfUzZVoOFjJpus45jzxh9Oj
zy1AVWpz3iRi0QePumOeXgLGI+TPDAYneQNKKWWlMUvjnERe7KikJsRIq2FQdycnXyxRQrEYzT62
f28ENp9t3Bwk7lkSzvpFKTYPz68h6A8h48P3mmo/chota1YONl/GD6EulEeoXgeJ0lHwZhb7wlRu
zUsLZzb7/XGWDERZedgOcr6W9vyG15Vk7BHD2erkQ7wJOg8WXqSkutSbwSD2ql4/Xn94DYp7WSEr
curaDDKtjjnB3MUb3gbsH3oSoBGHfjsTXKqHsQQmYtBZVcEbpGhsNxJ27pDSzOxHtSJ9vNMZtS8J
eoCgrFckzN0hYTNdEtJ6EACI8V2W9FGtSi7002uk+gexeUmXkP6a/4V40KFw4KVIswWDTLKp/DRd
ndtHVN5d1HTGxKvNF5Moum3DuNs15VJmAZNvl/MkbpNrTstg3ybrs0EKGxcQbdobZg6mYedFsPmj
ENSgmTmNi6fueQQvOyMvGTdLO9lHv472WjYmsIJB/VWQOuNx95GBSW91PYAY7XCVt6xJATI2nmJn
kLUyW/6JWFqcWL/vZ0Z5h7jJ2phVU6NxJZb2QpmA3oYC5oZzxtLV1XhhTnr4TP+Ooxow+CLuxbSG
LcPnc73HKgTtRcLrzNP+iomCWyYj2qBf5ikROlmwos1bmY7Xt7hMCJy/VqJyoxq64Iosh1eC8NDk
bWrWXAKySP91QwtYnKHyX7YShURjp0dcOHObXHOCrs01Yiez/35f/SEaUB5CNZy/5S4Lrd0CPT/Q
N+rtkoUP8KIVDKryW35b2mm9kB8SRPOEHluLScldlvy+mtEhinFTvtskpVrZ57cpm4W4rdnIvjTm
Z/OqYjw0QGq6NawNC5+o1tneBv4pCsEWwikvZ3l/KBqHVdrnD5VsQCAkedwnUt1b1eeGwpH2LlJi
KhT1yXsBhtGi+SnWhm1NokukufzFCvogE6DceMP3SQDCsNAnnuVwPvsRfScV7DV5hr2RRT9AkR/i
7tA009/MQHOZYpXIB8kSNHyIEIBLDzQwnUvRIMuJBD8Wmx7GYA1ddTNqUyJZf8OXZi5eBuEA9Uz7
ng33ZCiPc1xnXVfjpl6rqLKGrYdyYD9ViKMdAHcj63DRWK8Ruhb9YlV8B86yBKqx2uB334Enybsm
aL+Q3jgW7JwcPePyUxG8ExyoKy04BOZURXez4keSssUooxra2EtdcDw+Q86ZA7i/vrE6FrBsZc7m
UV9rQ3jtIeqWxNvFy0o3RjYgdzwy4krRWmL1nEoTbM3HfvnoEnAF/c4KCjzsYWRQZ+0s3M8cMOLC
fx6fuPBevQCtdItSdu9tGLgY9+I6GOPwY/62kdid45GjYNu9Ki79L4j4h/4IKKFNpGd06ClF+SN+
AUizvmOrVopFNvUKkb8t/Dueuto7dlxTMGdSZSxtQqXCGzhwjaavBGH81SqvoeHd3cZw4pqqdunY
0FMRCoxmAr+MvzTnN6Kk57lr/zRyrC+KBHIyt+0yPgY+8lei9oOq0juM9h24+9C4L65PLpliUR2j
0JMtA9Cm8tvmIv/AprQibglD3uD+7RiSeh9jb/5L7NOkEro8LG5YIaVkFCzhcxu4K5x5ZH6aeOBn
iSY2lMzR6L0XqeMN+jop779HLMZqR6IYgxbRkdubVL3mlnYXsFA2a4RmHZj+wLka353cA1XM97sX
xdzCEbiCZ1k5ieFPo+8p/sNvnAGAzhUr7rav4qrrk1d8lYkrvKCusSo9XqsFYNguBRoUQ4OowziW
YryLFvDh6a+38CjdPXJyIvGxw4T7k9v2cjTF4o19QkKG20aMQtIKDMxWucUoixStiOsOCgbwzW+S
GTD54n0lapP7nFptR75YvD1iFQ+t2Qo7D+cGm0egq+ddJ5LzISIfzu71re1t8UuoAfJdr4HoI+5N
DfVSQSVCw4MP1N1u1KlSaHk+ukP0plHJ5u182vfilSF/ZZxgcJVV17rpgiuCInPbDMSjlNrWpt/W
bTHwacwTNSn4oJZ+lHKG9DzXiF72zE5H3zOBi5ScxCMWvx+Q1ah5VeIrZylQCUhpDq45ThcC446E
4SMl7hncLzhPLRM2nniV6ywbgtyGY+5gjWxA409dsi9ZcuKR0upweRYxFiYD2FiauecxtO7W8SSt
Is1y+ryt1ahhwzM4jgpL1LIxCR4teWBhO/yZYjsnHgBAXx6oqDqJgcooTnxRuP2P/l/5Z3NUDLR2
2DZD/GdIfYRkiefsKy4Vgi4aDXBef8VbBuPth5H7z2957yDQclBJePyr1RTPSkxiwgGk0XPXH8xk
oA5SH3LAVGQVKaYjjCogF2mkOFdCdLH3w+jfOHQH/tPG3uTZUVI+sD06/pLI2w+d9FyIU+LMkEjn
oWyizzlWNwtslU3mETGAk8BjtN7PnZlowPXCr0/y477dAhzNalrMByhHxF3HtExWei6q5p903MA0
WC984J12XN2MeK04nFk+4+CjHBx6gH5Ox8Q2M6xntYZjFyO9MhEcUuEd2h2L0NSfwS70/tbhoNaa
7B9aovgRsZdBSEQmxVw+8Oiqk6VIu2h7YMjtaHPOntoKINVM4hSEo0AA9v3j2KVRrfYSZSXxk1g+
A/PYxTl+VDIyYob7z3P2lfgW5IX4oxv9J91PDnQgrD6ZAgyuvv7GC4MB++jwfTGEsYwZ87vqot9Q
L4ACRMSY3oLT/RJ2rIAa8w+qI2n3uHZetkT6CnJXUS3h25+1MbI5urKryL2PR39fvaLF9VyJ2Fre
FpqFuon3HmIcpK3mAF41A9cxblyhNeRC7+GgOE8WKL7tyQ9xMRPm/MfrT5qex3+fsTuKLZX2sWS/
dLT9yj14Z9m57j6Vxe1Eha2RjSrQp8FXUf1l9JPcytOjByTArGYaoVj+QTPVeV5gfCCKl7xo76wM
AZBho996+qIpQVC45dK2wgv0FWI7pUOau3IfMQE1idzftAq4yrTsMAiItgHQSJDzA4wff379SwEy
ZrN6DlZvGWHFYvsaw7T1Q7wgwQ3X7PnbmzmQUJIPmKkHJD38OArT8K++GbMSWSWgBV+QlXgijAc/
I6N1FM2/C1AzoRNUh3bpCoQ+Qn4t9E83ynYjuEPB9CpSRyv6V1Zof9KC3nD0WECMQC7u3r+X1n45
t2v33L6as3wvCdMUXoLghZ8llAciLhXiOVKVZpYe70nS1ty9L1OsutN4B1rAo5cHhcmDlWOykPNZ
LNgdI/EkI6grF34oa+3YGUlFjUo8VRMLk6w4rr1E1f5DUHUItmUx7rP9n4G9l/6Li1SIE90gruIX
Fn8tO4lX/8FX2AJ+M8/dcyvjDNLerW5lHV7NixsLbK94S4bHJ9kfnB3dlfZuIjvyp4Uc7dBUon+i
qss5RDWDTCu1uW9p7u9UR3kjg9fULGMYMEhMuOCByp/P8ClGqiIzRHgG9RIUC5q5I8KOyDL8gH2F
g3rU9vG6ETljA7ZTVXUq6+Y93smpci6rqo3wYb4ELCRdmcBKnbsUZudXmcbXQha5dvzTkIvuLfbX
udGTomtwBK8Vyjz8XN3fJNU+mJ8ufhcUvtHCI83GlTH7tr7i4+7qXXgvPpoBAvzMOC1yZQ01OSTY
N5UzrHkMZOnRMGwFC6SNTBmYt1F1hypyoK07oM2+ZwWf+2K3xH1esj9+W2Sx3vUN5r51ig5Ca71M
8AlCEsHcNgYQmhqS5Cno+BNEJaSFVgu/frD/EnwEt94/VXEBrOo62obD1GT7K4ZUIiuB+4MNZC1N
3TSuq7hT83xY6C6HqOZQKC/ZSGgSGzPZQ/85q5/2a6JAlmZUoMdjdQZdCMhKJmqvJj0yvVdp96m3
/MnGNAbBLP7+gJPNDgtMjJtPNWFJVLl1ho8WZdZet5u4RcylFw1OFaIxLDZWXpj7ZMnT4VqAmK2E
5FAZi2nXV7SFWQ8IPvF2LSmKGYMRj7RMntO34fK1a2ezKmgwrU+4m7yw7RD/SvRt6CXrQfiiKwE5
/Zva3XFMFGnzucwhQcLE+gHj3/J/dN0mLw81t8+QgKrzOWE4mMKeBZaXueE25WTqu3uChUYMCqFl
q/KbdCbucgrAjZ7FiyRTCwZF+c9Wcr/Nzl0tPmWhj5jJNNTt9m+8lbyVvR0d+QPsMRhB7kRS+ptl
xSTdexplyUpiNVxc1skL5bNx1mfhB1QDwlNX0bXgCEG/hnoHxIkq9IOQbJhx+VRlfHmm0tP/K1kb
nvbrmG7/arCEM81tjdKHyUaPaqzQpK16uJHMn/JVJMQ3S5OUoJVfk9QvhMZ7hTgUf/alsmY5mVcf
7NsxSzAdutfp0CwucKMJmdLaZc+Q5YU2bbrsV7hCYNoj+U9IpNhYmcUORioculENMfaqqmn7Py4B
hPa5n3XsEODPRDgjn7aJYcL37iIoCNO+IFzjrUtPHHwBiK6oIbUijcKnuPH7daAh21PLW6q9XIUI
0yduFwgOP3jMHeyYBd9qYo6+5XIrIDs+jJkVVa+1+2Bv6DOi554yrv4eyi55llo7v3gxKON/jUsR
vdWNLr0dfL3Kai2eEBlESWEPZqcuokairgjPLpl2dhbDY2e/06RqiPiw9U+aUWu/pE39xWtADlmN
3pFBU3DOC1jTB9nxg3Oin10BaRZDl4QwSXyb8X/hD1w3kxEk6coP/YNdSuBhToK4hOdCR94NoAKc
FrUABl+egqI6nqsh/iKJwE9yH/Uyw1dxc5OgDhRFSml7qX/U20pC88btQNV4H3jX1s0ABMQsA+0k
Jc0v+Nczskk4b5bJOg5jadg5oKyWmoBQcESI4qhlSa7Oul8PIaQMWuHag/xfmoAdpeT9iZ4dpk0T
4+cvTGVMowtg0ZSi7T94pyYIPLdfLSuLQAMMVMml9p+wB7dYyRKyy6d5nrrCkq2ks/MrlEKKT/m9
MIGrArMOxsLRofCHFQIz5YstVLw5D7zTlD8lBb1kNz5p/5UjR5wPTDrbkIf2jdqvs/0tJprcJFc2
CPPhHkxex7qPD9rITTcRCBMjpa+v4VxBjG4csAuIamDkMB6QDASfHJGiXd8dC2dnpfajxD1+/M70
yj6TFYZwYYfuCnyFDkAcZbWQOMMVTL8R9uRGqBzq1Rp2HSPRuxRJ/pJ2qgoGZS4ueAsES2sp0+FI
rqxSmDaxjl+s6T3qd+Qd6QNOR7itslp5XpERlaeRb6Oejx3b2NILfyg8kGcsysUf4/fKad4m8YMI
3MYIhhMYva/9szhaXVuWtMnEw589xGiFYh8scU81JMykv7Z26eFTyEC0qqDL1qquqYFxy7siqfN8
y7jJT87Q+7bIWUFqiFcC4nyR3sxEpJyDzZqBZ/BhbwMn+Hd/OliRaM0j4QatfH8Mn6Nlv2RQFZJP
XFvfHlbRZAalUVwxLVSlNCDwl5KOQdIGC3kRdZeb4m5fPzuf8hiydQyPlanry4gdNEXthmdrFam1
J1Sp4tQ3id3+8owwI+vbVD9vskuPd+sIevYDrqnWbMySkBhbsTSNDUixodw/PrCpzR4xX6vLFlwh
VTW6Umyo2Ic9gkCogGMBig7Iprh79iDt0NdM4g0/4IapycGoB7mDybeudb/DcqfM84awBmV9ozQ3
Vre7FE2xaqp0SCgXZ/WnxtJJc7JfIF88Q0Qc00fbKDBZOLneMRZOD8+ISZ2YpB9rg2QfUvSPsq3m
UxIDnK9PMHkowQrBuR9HTU2+AP4vRy41hQAE7FZ//2P41UGlYUrFl0lBjxD01piRs4QPn809wqBY
Iu1MiJsE1ZlMgS81P8Mh9C71jFcLJ3K3Hh1jV9CAiYRsIzh1XXjUlS9BNZdV4G7zSqP1RrBU0rb/
E/holz/OrUYBvMgIiWUPHCg1BGCEIiWJGFdaZG5lE5KZ4nLCon5nhAaAoQ3OUnKkm3Pd/AkaA63z
iFammddtlkRa1ZXnjAjBs2IUXjEzrrVtn2ZN+Mwp+/98iZdg8SVoatwmRR6eDlxeuwJ5EhzzyWV5
4W3nWmgAy4VCH15P6YcJdfH+VB5ohR2+YHQXM2pYx4N+XvADF1Eu1n3MXWaP7U4eoIlDELLvnBPU
Cqf9Iphj/Gj5UhAB+iR+YX9mQdWLWcQs8qz56xJrahSnZHUr7lJsv/bmW2wE4D3sSn6VXXi2hQGR
YLtQ0ksuibk8FKBjYvZ0icLQ8+JcxuTy13kU8ZNuE9DLB3dLvMt0hsrS7aNikbFiKoqKF6nkeTv7
86f4DTwOSpGba/FOAwP6hX2x+4MAkSrxpPM+9QqsnXBt9dGFp5wbtxjDbXhIU+VKgIcIvUDDO8ge
hMvOvWaI0rQiYQwoGk6lRoNUuMmTqSywRunGlSbwUvRrefZTDVuWzl2A/9lJuRwuKkJECtJo73k6
59AGBDUu8IjsfL08sXEXfAfpO89DJCQRMZb59RGM6Ckgtl6OaLfwfb1M43KKsf9rdzklugEVMZ59
D5z/Hfmp4Yogk8VMgBKe1+H2atmdk8LSPQ+/Nn9BO+vUpUY+So5xS2CxYeF3VRHy242iitYultmU
eRvH3VedTSbzYqv1LeSKUT1bg/Cbzb8XG7iDkwJwDaU/es8Tti0/g7nJAZOhYIiN6ozFG9lHx6L+
bKZUV6oPOxuHET54G7UJJ43gMjhs3NEbgD5GCFMiMcnTB5192KO3apuBYyXkhQ1FMrf81rzhwgsX
0Ud1Nh3UfePt4gpPr6kbxE/QLzX3SfkO/zHSN2TgbppOUxcw0BrOAtVft+gfuypntZgwpwcmP105
PE/wJu4qLj6eogDzguH9UA1g8XeSZu0bmyCldp850XJ2C9kNSf8y1BgpeEZ03xPQ4Dfl8rAxVusL
bGb+ggyaV8tlzDxX61cTQM4VhzKGiTcqPMUdydzuusz4JkwPrli5Z12om0PppeAbPMREV7EliKJy
TVC+yy1jrv8qokGWdJJXrm6eik9Rj3mhD8vnuSaRTVWw4G/WthkoUAMke+lk4yaMDmFZP/QSsW5x
kLIZbKvsc9opQLMMEYLLIM2jt0fPUE3SA5ZeNVj8xm/7lJnw0jbpFrQ8RFhBsdle48NlpV/E8YC2
0B4MAZjemu3MZ7zOayUQ1Gix11RsHTXyM1w5NieG8Ljkgoa8K5Ej/Q74lKa///RPDYQN5YIv4DSb
jpmykz4XLfmukOAUUhmZCf8ig3k0fnDyrfT70EoqGowrlDfi2QX1qIInWGG+VJp3AFg3JWOgYG92
XyP6n2oKeXZoWE1T/Le37ir554CcaUFfnMsJETbP13tzzdQKPFg1Rr0Jpmys85EH9EYqRi9imklb
3Qomc5/6qNF+HQaPM08szavzApBit+Ze4aNTItkpS1YsBdHcszV4JdRPeSp7iC3f4SolUYAwGyum
10NAKgDxybo+uFxUwkTPL5yrmdVQsmTkJ15jhaV/EigfF6AaO/effAG1MF+gJAaE4+a11ZBspvEf
znc+/hCJUemRerz/k+ztJDFgXKzGLIexM78hSVl7SAoF9CUjxvDCOFW1WuyJT5ZsCgb0QrVsVn6f
U95ZV0a7Elq1N8y3gX4XzbPGzQzASyeLbPQJO4VaZf+EYuvNQhmvaWfOwRYL5i6qBifUeDbgfPNc
9cS68a2s1Jp2lBhiATq2ODl4OUE6s28khntqhAiJCWtzQ2d1BzUiVS4W9b1ZUxaN+5IIoZdl9D0J
EIly6q1e/7VVQNEsFS1P0DiJyZT+CR7bPK0uN6VYoC9xfHFRGlSbsuBkegJzhCFULAPLdju6XtDN
iDuDwYzGC+QNV7rMIPsKwR0RFU6nEgnF7LdR32SaDslwRZQ1szNYlc8El+234w/Gga+pSdEYH69W
yIkoVuLh6Rku4O0Nu2peaa4g3yjYgI/oFTG5p3RiDVNdRdrJ4sDDTSAAS8VrVp2tZEP+CoX1xqpr
WNQrawxNLl9a4uwYDz1V9s8ohrGhpyl2fIKRObaR1rWervnIe9U0Mt134MyWpWIwXZDZiINifPOd
6XfnfWKcdKEPBcilFLLBGQb3WznGpAKhEgHfsjs6V2rueacSujZ843fPLUrhvqfcGz1upB85gY0y
giFa5j8OCmTsJPAXn+BavXlLZIU6ZvJe4nnVKTbAVtc3hL67X2RhD63tz86Q30w9eJFI+Uel+yX2
qJk52MhV4QG9saq8/oClAV9VU+8uawk3XLy8Yl6qhqnBapqwqUHPtVg6G8puqRHvpnAKymOlo6Z+
2L9KRlfI4Y70YPLi4bJ/KVUl2fu/JSeco9KF6UJhdybYJqM8tmSDPTtH1ikB02vvShc2uyEC9Y0c
1RKPvzx/wBVCZIOtTMmhNqC3H25kS2oQOv9jOIgZvgMdLktJPHXKPKfjAN6f+ubjTlN1j6kyaiBU
BSUfwSUKC1Sa1k4h+JPf0OFjduOqJLj8mamPFe8l6jOx3BQqbZJC5LeYmy59+TROlIgU2aM/D1B5
LZNaC3cv1tQAwRV3zghb4jKOU2iR5jETozA6nznvs+6qnb8UyZ2nV15WfqDAhv6E+eTojYO8ylkW
UkRnSUgWTE2HOxKeT40x4e2RgRuh9nZIr/l/8TtTYMLMAq+0K5RGsHkwQTE9ZtujQi96cipFSSCR
IpAFDnlvlNvi1sRIU8wuVxLG1QGo5+6jdMqKiudsFi+g7ZsJMIeyxyoRijQwe5k7ghz1LXOhGIn7
6YvBq64XbxD60xcfto4NS+w/U/5Grdxcz3HzUXW1hNtPHZdWYmXBmDpCgvACgNUZhkBN2H2yJeoQ
F6PqxOnd9sY+rEr3nC++0MV1O8PsP/02D+4+Ie32ubTMU75S646MpIIeqbKTpGuKxF73t4WNhxJR
Z3r2ZXmqRnRLgZ37Wyy/wgyJ1MLjrctxUtIjQNcGS7U/Fhx6YyGX4CUeGTdsVf+TzpMOuKtOJEEZ
SCdMbRXSrqU9Tz00PcAvKJXHycG7CA6Nyc/MIubU9bXvnBuwrJqcgiJ1/li2VUrEuGXQJGdbOC1G
aXvgVVscK3PrzmOEnbIXazPCRc6XP8mtHzBuGFj1FeH967knzTpkYx3GwXzsMiE9ziVQWypLyJkA
Lzt855Oj0+yHYElZyjn7v8NTBTcJW/4cxZ8xPgcX740L/vUMsodYIsjdjhX79/vrFFUIeIZzemcu
O/6JXrl+xtSJPbOOb4UFF9Kdh5+s8UmWuMd9i8ibCg7F66/uxLjgexcJ8L41F5Gw6KDe8dSO8KHe
KLxneZOsmWut31A9p/KQZyGz7YUY1D6LRJUj1NinA5XDOlLWZx6Lu827HoOf79sxxprViBUvALAT
DSVcByLLfhJfArY8Q42pPtrZ7tbuL5+tKktdS5UqH4CgjfO3cu+x/ezqIqaenMKYLd0t+Dku+EYy
AR8Rzs9+OHE25RxKen3Ezi/srRiKomZ2AKvtaiZWvY9icoMjHQ3xE38ehmoSiEQRMOglL/ZE9BdG
czcliPWuW9XyQ8MsneAJdQHWWHN13CVPfSz3ad7Jgq5V2n2OMQGz2WdJJjiUcy7Cvd0lNcXhqzYc
e81p3DNQEAbTxI2aMCh7jRNrHgLVtqbJ8PyfjOWO4ghSqEu+134+itungBZGssm4QHrjixAXprZD
s15sUuSKNSJ8UmoStcYgEXNmg5ri1iK7Z7l/y1rSEwhks0s4SJllwu7zJBNQUZhFINUa94TzIAkH
JFcElRc8D67YAAiShQd7Xi8WNzKROTme204+k5opOZ+C7ef1sWw6MMb6YgJ1yZAl2DgkHAxAaGHl
CgYuvYwq0b9u0Nh7/dQIIlb7FuJLyWTlHA5OjTMkNZDoHUi8scufrUorjh5Drg2IVKv0yqD7ZVKl
rE7tSY0dQr9zZO/2TS+CoDFmCQuSHuVtun9PNVKqs18tF+8HXobY7hTuX1ssxn3oKNTIUwG28zO1
cOSUmiJswFOMFXi2p+HooTKVumUhc3gjGwH6V+/xHqV/88QIRSvtO39VQUejqdHznexIIyJoFBNj
4+A/WazE8k65LGzHeWxFJQ1IfHy3S2bnfTy27idsRFNe1pe882XlbfBt4uV2IbvnbJSZcJINnUbA
Y/SUQahyK/7d0k6rUxnX33ux1/SQgE+LjUJieEhynQ3l0A+7/cvPnsK6lXIeJlzOrgUXeAwqqnbv
WvQO6XuCg5S+H6zfLSuq7i2Tr7p3VKPus8uKQn6Em81dbmk5HEhTxx+ACkBE+eHJnFOpK+HOtP9S
8AeN2ponyP/zz4iR1d7V2vBbOuPWrLRmF9Vj0x7AbFaI6EPEC6DxhgtDMgVMwgus2hEIx90wDA2g
5PVC6sEr45PHN5IPLu2/g8rK4W0HOC4FuFPgwWkRdQ40WZ41+UL9vxjaz7Tnv1UEtmy1BcqrFyc/
CQA493U7jhZGecTsAhDf1PEk7IRxsLDRg0hNnTxUmAs3Cc1q5+5tcZ41eHA9U1qFaU8HY6MNr8Bk
wZG2GZZfu+DNAo64uXSa38wZtwKWIdGQrx3sy4MoZBt7HX4PTO3bxcI7NnS16Nk6WakINwge0h1m
88ZaHD22AZxnX6ng80bJd8lirUeehYH6B6AvDX94B3BYcoFcDnQ/Xx4lwjAYVuixSq9gVlhSKLuG
/uzDiSFzxvEZvqSvkX9MHgCejVDw6tjZUlr4Lo0mPKxEvxvHGMxv5WSjoVnSfL8i0CUrvA3qIh/g
VBiYTTRRPYr/l1ymnizO30yUMOpsZeAorG+FTHZYBRwt/zvRRTz58oYnuVG6OLkTHemAn7qB8u5c
xWYHHNGla2X4qTIFpql7g3Nt2QmkL6R3is+l3/HcHhsfOKlbEY3g4oJFmsGE1uJAc96eQBTrnfch
yNNu/Rb5/7Q28if3gZy4aYOys0zj6E/tIzRuPXkxrNqOq4tmuttPqSI5CsebLO0zdWOJt8XlyDBI
iA42XNWyK/9W7W8V0SVpCi/whf1MjbyS+2rRhZbqGgEmQCL9qgXz90nnvVW+m6DWekobSHhbW/3P
HQ5Y0xqrXjLstULd7vd77PbMaICoZqI9jpSirCppXvXCk98yFEJJ3vetQTcl3xcDnSDv7FnlgfJI
/26JnSnbdmHqJK5veF3FHvryuEBQcjcUhaww1KlRmJFjdwtvkNAtvZvcaJH8HpyQpmG71UeFm7HW
NDKcTguSEMm2LlMqnseKgnacFKDqnBgmRT3MTQgJs469KNI6jzsgX5xVRRH1vV5jFR9ttmOAimXe
4ixxhIBPRpRyG1LOeRr1vlkxIXzpjpMSZ+cFJS4JVYflBfmBtoVn2RC2fdAdBYe4kuvP47Xc2xNn
VSllG9nF/elwbtk4b5x4IHLVJMApZY0r4Qm22IW2DScXE3Lpu8cMGHQeIPUwNdHkLxHDb4nyshDj
wJKGgJUdkrOdyZ9gK3euLamg3Fix6YJQo7JFisM58cmJltYg/nA4pMDPi7Yi0EycCtc8Uu4F96oD
7bVTQtub1zp6HO9CUeStEooHS7UFBQOnuHDjlHUDG1fQT3T1bp2dB0+0HAGYNWYn9NWkpFU37GyS
cpixgV5Lia1Almh0fba7LmQFU0A+NICGq7rMPXbYEfAR2xYfqU7P8QFPpgpm3E7rYW04YAszk2aN
CYSRP17YWrUwUpE51jfdO9duQjM9n1hbBHuuwKOop5xtYHWBFs7mZbJRE7a9JSxFmuK9r0cMMe7u
qJ2S8yqUTVNlcyHwwYIhP8gxx714865RpicARWb2MZjW/3hVtsreQqHRSr8+5lAfBNrIng+TvFxO
jyZnSrKJa+n5w4rYldn0z8sQM2vLl4Pbs8AXi0u/ALjdDI8l1ic4zVZCtwjE+lQrwD+fxcYx+lFa
UCGtVgC/TYU7ZftROrZU3EkVT2nzy7IwZKC/uEt9Vgj2kECoWVp94z84uAlBAUonIoBqBbooXWHp
wWB7jGy0+NB90NwzEsQD5m64wZ51+yTfCUfkzad7ltPo8Z6PSDdQC62o45gHbPmUvcj3vXj1PQUj
wvyopCRSNkkOsomkK7mydMp+kOcuBpAfjgzMuhbfGUlw/ryKyp1TtOlmKIgpazQzqsSFGZBGB9wc
vCTEyK5pcMl90BQYYlmjcJmhZsLDVb3mKAUprVCWCCt2nqifGEaWFs9qA6AnzoHz8oOuUPpkMLrN
LGnstUa2Ka6cUTJNT+8JH9BuPPcdwhIeSJVfRW6p0AWiOp6/FM6Hl5ZRdn7N2L4I8bAZq3rdMvPh
r82ktoPjBtdgowSqAMO7LtPm2QMgn8eA6Gtg3v1vbFD3/s0YvuKb/4BxYz9TJsMuj5iWuO4+9QMC
rZ7jTUHUJrCkFaQzD4o39SIdzSXZB0CfC1NiquOK3AsDE0Z0RNbFTOdC57XhFEAxHe0rVXPtDM9U
KNPFmEwQXSJm6XFwBp+QNlRWsk93T3wkEJzvt+14IxYzSD107SzzBX5ScdDED3n8zaXfOZuuwfu9
u/WTggZPFgH9G17dlk0KY3iL9ZC1Vy9vkhjOnDYWvczpkQy+vs8gMl4aPGEkW+O6IFdVY/cNSCGo
8d77TU283B9jgFlsws752extCuAkSBHoK5w+3byA0xL8/T+A1iSzpRWsqNPTTZMPXzyBjM0x5lrq
nb+DCHufsKMidI5tFm96V7dxjm9Z9/0gjt2odM3G68P4oON0mZIU6e/SuQ8rdmWdbPswIf3aG1vD
PiR28xYBc9McQBJyN40LEWjNeiNXEdfOu3Nq75m5KqsLMSgd9pW96VYa3NjIprF3jI4H2bD11IC9
ftJHZUkKZMusk7rwJ9Zt+yQ5Nr5VsSve4T7A+EQSQgWS3TfvsCoET/SurBHOVjhzcI3aMqQAe9mH
4cVV2VPPd2cr2YnNFjRAd7mQFY3MVNtT3iSOAARqvSmpKZeiFPN4zPkQte9EooWnuQhk579cKs/n
dFjS/qZMoUy3WfYOQdfz7YcAh8K5fmR5v9mBpfKao0S3hiKEKeg631+EGAI9pSCF/4VdfqZiMvaJ
ixwxk4h2jwlnssOmzBxygDyOe09dMMNta/YulLXpUXrj+Gx9uDlwA0q9Jjskf3ieBn0BkvahR5MO
lwJ5MWQcGRZ0yL0U5YNi1UcCICHJKQw3VKoEiWMroYdZEH17qg0KZKv74JW3FAVt+PiNEqya9ItK
WZHUCeqxxD2w1X0U+cVcZ+14vxFZQeOkkixEoxEjKhCHUobWrSJmqHG9R3FQjVnZRX8zy2hmFSUm
Uwta68ET1MsFgXZLkEypgucL2KkXfiKOcG64DMSXTg9fRhaf/ybzGB6Uf7BCQetbBGozd/cV5c1D
nxMB2MOjoKZZs/cPIaGt3ChmDrAHvlalC8LFNBy7KAEDOKOfGhDz8nesrGk0nV273D2nv4BaUYEd
Vzhz5BvPdafDN1Que5sJHluaOENbm/t5iA/SZ5VoolH+B9iAbf95ejYXeK6dD1ZcOPMxak96Sf0F
NwLhUBABvAAichqHVcRWvNaxxBVRb3keK/ndk+ZVpwz0ARIfKYYjUzkp928UvNLkw2wdxJ7ZzBJA
c98yQoiPOyvjktZ1zqPcUfvQ5lcqEKu14y+13uEus5cQwTQbR5jTRNMp8jcREY23Qc+Y8O2CJ1TW
23nBGUyjoIMQ9ZNHNlLGL17JV3UKIKhlq09/oG1JBca8tuIWIIo43uSszwcAzpwa6qX6WvZmG4YE
J8WOlhjpqlz4TbhkwnQLe9j1HSM7MCH4dljOoG9mNPlxf3vwdq5LrlgsudffUHnkU9u4T9jjhTHn
vejJPrCHHe13mtLc3LweFbi2wDcNzlxd2wFQJFMcBu1dMejqXCwx+vD1kuhWRtEUVeaPG+QS3jqZ
VEL8rnAk0dbqiW6910KrtfkyPdr6IJbrp9PMx9chMAL8tAT14zWo5l6B2M32b/054nQDayACDQZx
r6ACh9999wUVRw1avvK/plAtSaceN9VhAIdKpu/xqzeGQLaSFdLFJg78bOaGVey9QU+Brq4ewbFp
rX5/cnGWSWhlFt677f7noZ5CJfgGcLSAMvghkTX7S48ZgiMGjCcdaWTP2N5ojxflp4MamLAV/58R
6MvryiIchRkuxJEOb5nMI/UUWEKpShwPFUZrWSotWugboFmxIVIQMVaNLf7NNTIHO0joedhcMqUA
rUbY/2ZsjhaJkh9NLF51w5QWpxObLSHxbRG+mQo9iJBt38QeMw3TS1jy4hbglMWS+VaHSljo0q21
yTUW52/7FrNwWJNxGUm3mo20JqPpnF3unuUJzWRtRcfgXrd6w3QY4fwuMrGATHkSY/9OMU4sgqRM
b5Kox+9zVM+dQNzLEnEYcfiZ0XfUDlhD95sVilF0D+mxYB/A++Z83tcFfgrhYTTREcswf33JjKjl
9+K2FipmGygPLOCDegg+fRFur86jpQkhlQB/BO+m3lvUPtRSNo4zI5pJVqSYomQ0ls63OSkZbV/8
0jHzelKLFNpcs+NPNKaphgUlkLc2EKlB9FgcAAVQbst58vP7qzga+NmwfCAa03choEfOkKWS56cJ
WI+FPxNp1SIHcV17FRZhBCBgRL4rF1Ihwvlk+/dMa7riZ6PBhU+7T6rOxQ6HvXW1oly48sXb+9uk
AjWatnm5WOSyd15ERsGvuNijP+Q2Uc/RbnNUUCRqh1I+XaUKnGZaXL/mFkQ6LMy3FDSg8hGn5/xN
2EKbH6sgX2+MAbKH+N7V3md6rRCeS88LjOG56uAkljV3zJYDuK5KbIb5xtXrxUIK5iel21GxusDe
kkL2IBAqa4E86NwQYO+BA4mZKoaOyov7rtuw/du9rtOMs912u36A0JUC3Fjj8wHcF6uA3nyMlvaB
ZMeDBNCYZCrpi6NxB66xGqYfGH8QkiylFlmHpgwknwSep1BIhn3mcRZN/b8AEDDQyaqeVjS2eTQe
zG6G8/IwLfWf3g/4NNdWCxaI00865F5xeIUHfOlieBWXvJIJB9UaWiDBAlfaaktnAcbFe3brvPnU
L9fLt/p1ZnZ1n6YNtxaKOK+OY8dEKvwXzZZ1QqHRXOVFJ9bNAAxuBFsJB8afBfKw3zgDibMG3Xe7
XDdhY5AXTbR5+2dhQ2HrjSM9KE8F+0dRzE4P5p+GTZHYvRIFoK2AwtM5u966+ZvFnaWeGKTk5+Dy
AsqVhiCef8dLnyzUwzRuIWIATL57GfeDY6WY5nwzpXZc1WMtY5BvecgbEbgvnfE6Rklt0U3ArsyA
X0axmsetOuxMwZJ8Y2kvKXNFWbuFZE53Q50yWVl50sGeVFAiIsBjgjrX6x79YnuJaQg5XxPDBrYi
sbEVRy+fQ3ZCWe2ORXIm1Sorc+0B6dqD+RTwmsSGM6PLu0ZTIAjFkh2WaYXq9BT2w7H+e4HJUlly
3DytskSLufJ3yQ5YcsbPmr+D1HVfcNQuT42JiHnJ8sZeii79ZTQCEdcL/RIUKq1ObCXJpaHqrzlq
li+AORrAS/hBjyxe853S28X51jmSkylQf65UwSZdJkJxDPv4RlFnzhRubAbRHdtV4EVBbWdCKrZn
f2oHd2S+19rAR/BKkfH6csJXJKQle2oHf8Vpcmtrivcsg2lotD1cGJIhWR/c18o4CEDdYuqOTkIo
Ck0V6FfwOiXg2+PnurEJkgLvsKIR3MQYmz0oc91kwT6SovKiH+HZnznIl7JjXuK4iCbpwraTYM0y
OHXfIRgJsLKijEX7gnWBFYaukevwGEV4E4sdS2pFaKibjIoxxNt6HXMyqBm003lj/VbGUq5uCy7o
XZappjBYIUmv75sujXC/sXbpZhIC3JIrRDu1chP9n4Wp7XmrhqT9xyq1yKTPUmY0aY+X4L/QQq/g
fmY2yV1U/LxORFwvMxnuuOdO2mGORrDWtcOgL4RAA2pVGlD+/9/hnpUzZylYtyCbNZUHUWKgGXpy
CAt0MAIRnypS/bMCVikvmW4qe+pIR81oR8aQicWa0lPavSSj/CBgW+pamIVJ1Gkn8dzjAz5y+fbr
AfYz+qoaK/hJfVbT3KPzUir8CLUDqheUYU41+3lzryliDrx1qMWUgxy+ENokTJlZ9my5wNKCiJPK
qrhuHlNLmyAPOh4yZGvWm7sce/seyci4IFAC/B+QxsDaDJlMPSst6zj1rs/oRQZPWS5NNb1V8phg
snAwKSAQM2b/LRv5ve734GwI5oF3KuXKFvO++2DGRFLDnID4UlnIOEcVN+TyjYc89PH9rdVca0z6
/hL0QW/qhUmOFiO8M80fI8cTdSUEHmNNt2iNGUzqGsmHoK1OLGmc6L4OAIMjP4Zi4nA/5Bhq6BEB
/LPjAoOecJ2GVGREJNesHLh0vjkpOJE1sCqtqF3xtUvuCyIL33gW2yEZmDQKwSkq8/TEXmh6NMb/
zOXcYAVnDwvPiNnScuxTp05YAzU1SHSTF4cSjGHpCr9pvOKNnrqAMD5tFpFs2GRedKYy9Y/HbC93
AYtgzJel/gZlHDEqUUcjqB9y0O39Czo9tMeRZZUsv5CR/aWFd58wELSjSNjTtJY9Javk8n8+r+x7
fuxR0gZrsf5v2mDTMEiMOxuIrd3CTDDxWinzC06YNZOXqDurZljnvgluITzRcom4SAXWCZ0iai18
9U1GzcSZhUv+nwmYTz2QjmjIvgiUjxQJN8PupA3lznmaSzZU5WTdM7fkDoEaXx+wR+O9SS5dvC1Q
SeozCYOZM+5zfNt/Y4fcaIaO8L6589yfWqs0hJiZWK+7xL5gG3045l/99N3RAXAou49Qvvnnp4uE
JfQrGwYmgPetsPw40tPYABJgA+IFX84aiDy8/Ha42NTv3Rtgj0c7sO10erGdMLp71ee/35JOEGzr
6KboRqCtDJyvq26bBg/x9RLp0zTolsNbRGNMSPEMijPuIXxyrgJBVLw1iv/IneElOT2w0zpc3cMT
iFmb1dyA02DI0Q111BIJ4TEdz4wy/kQPnrWepiMxPPyLAvdYQv88/Xk/UHuFCs1ydSIMwFbLeFvL
BMvmgea1OY6gNSijY2devdCtB1wQqltHg91LQbg3OUVk6FlRD9UFKltvzU+hY3Kfeakwii3kgRHT
wSfAEy4y1w/P4wxd91yRsMoX1QxR/a8jA3FD3NvwV8X/vmRrwiMrHsnM9tlXvAslHOYwqHjO0sjb
6qpc6UX+JhPfyjwgzXpaORPDaGrRp/4XjmCfrjxJHSJMuF/8nIPWu+D8nUlqDg3Ls+wVfOA9yzUb
diVW46aAUzMEm7WQWSy5nrPzR3S/CWPgXx5kxvPPJCX3B0iNjjiTtaexcn7j2o/5RKWHy3CBjwCu
tVxrQuQg/3BepNqCJR+EcagBUSuZsHbm9zjsA2bRRmiOKI8YZ1/sgUk+AngQV+AgAJqpwQPbUmZG
ZbHPXQLaUV78NnyTpafRwn+Kk/Q6C4NtnLxAlfJOZY7YUXIPnHypnVM9TPNEpQKyzRgrNIo9GFH1
naWfklFS8x4qsa9e3uuydDoG5tWNaZrkFsklUONmUn3azS0dQ8o4YZxFBR4xTG9BVqbuqJKBw5SP
KqLQ3pFhp1Gftndso0Z2VuL4IlFU0dZENDmtuOFXHkDaCdLqTZk++xn7N5ZRaIEWwBeE9Vcr1rQt
99TGQHCZ7EaD4Ibz23JKA1e4iqzHYsIJNWhBsIz49Vwkfsf353dp0qg10s/s+a+a7ZbV2HMuFwZD
E6CbXmiPNeh0kPll86iFh4NRyIs+X7bg8BxJGCFPH5yxBj0DCGQb8IZvGab6mcC2Xdx4HPbMekcQ
6Ir/nE185LUCJxyEUq2KlWOK/Pr2gf8AX5YL9zp3hVjNBYHq627Zstin94Kbupn0kSgIhdbLi9e7
D/rWWlOqakPEOm8fl+KMXNWfRQ/fXdoA6r780xtHMCuS1Zf+4EDJkCZAV+0BjDKtdDmWuCP9BKHQ
jI9xMz283rI5eMhwn1uLCowduJzTMVWBnJwpVybE5rdUr4mGkaGALL9hLnD5oQEl+dkww51l3uzZ
wpH2BLIQtbHv+uUN/LowTklXo18gNsdlr4yf7xwef7pYnpPPRmvEEeZYQMWiJdiY58oi2qOl0rbq
1UlTd99rQKc+IveUOWxBaGxKV91JuAMj//Qup2XJsq5w+YOyYa7d4t4y/yGIp4DaNcK7BUjxaz/Y
MKOME8Bl15nMoEwA7tq7csoiB8usmsdFsoQtUAnGW10y0uYJ+MSPMITVcSnedQIflxYkwXXnt+Rb
sCS70pBtWw0ebbkpMsLZm+KsvGZTFhSMliMShMKsbwA3Z3sV0YcFjof0C5U8wSJL6Ym1Jglv6X6t
6nyR5/cmRtKn32W6t6YKbwwTzv6hHIwhSnPHYknHuCqqrOAaW6GUQTak0pYxKEItGKNMAWohpYkx
r07EZ9xH8pCBNEhHIdwiOkL5GhC96Rjl/dqTeYnaBn/s7bGOC42igyGQ6hfxiiY56k3+LIBny1yf
nmYJm2yYsDHzeS5f7IAH9V66IkYhT+rP0RAEV7/mCObRxg4yBzPKcihwC9VtMb8IEY1NacrMypn8
ab21prGpsPlSXWsB1tiw7StMoG9yRBAL3lRBU7psFtfL7WELUb2dlWR6JI+JWj4NMXMFwBaCZswP
u8OAp+w1DxmuS8TyExNCdyN+9zpS/9RYM7VgQRC46MwBtZE42lN6HdF1F4M4gPvkC8AXt5+hmojo
IuZUeHzaDLZ5GYTLWkTjqfubGDdVG+txL5DOo0t4XbeXegU/4FsxjDKoicfXW/fcfR2n9eyZOuzr
uMMhXqheatpnZo+t8Q686Tg2777KnQUzrr6YR9VC2BQUtpT6WTSEJFgrXKY9rftNjlGJpeV5H8LP
bHbSnKpu+tlmFiBvJ1CwZi/I8ZAlTUO5uO4L/SR64kon8ViKWdxMkJuuj6tdYBwif3UikbUf2btK
52VwO61ZNxMrNYCbUmhe6+UDI3Re9ligGccy0ojPCL7XBp9sXhliamRKkbS13ugMBfbhdnL/+tzd
Pr43n5LXdPtCL4FDzP5ucosRebaYy/45qJm1eEBKFphS6Dj166RaWt2D6BUzZLSrv2X21Z4ou2q4
IFx46wIMnvbp7CSKNCB0WyGWBophJVFBoewNB0Ph0wFJ/O2XMGBT0ZXP7gqOee6YNd79nBGdbaQm
KkgWvSM8+D+P2ToRTSx53u/xx+khQEOmZFOtjZBWJcXs2441N9341S3tmTqKQNraUxNdzt/XndUj
4tt4Y52FHhVB7hMfVmj9xuOWLGhqjj403q1PxDi3jAZzqxqFgFehvtvezz3yM9CAOrFCMNp8nQhS
jbaIk3IovxvAbfZz0ayIufIDfjx3XYB6GSulCrcrEAgM2fNcvA1YqG3N6KIUMyBCwluElAGbNYW1
8F9T9CxGYPwHdTQ0ZM/IEML8tbRmuKs1Y/UtJtj8YrvPGf2WzlEr3fKe5NyiHTQvTaJ4Bloi1oGi
STO+4UyY7ABxxB+xPZYqob1MzqaP6y1VK0oV7621QP0hg0/NDozTmI7HwhghKQIXYu+S9C1Wn/MR
M2Ly4FMdenb97xd2r5qbeRc3GiiIl4pfwS6nWK6AnTFq/IThRFB40n3EsXwWZnk4gUFbgGK91irU
fNvQd5jZSfLr/Vwn5zODUaaHOButaeJuIT9nfHv5L0rk8HQpLJqon0G0iAFdojyTaWGW+iknmymk
niDAt9q799rPRz+/vSwLDr9cUEhRIHee7QVcnGsMQESOngvhA1wa3DOUZWQk6Tal6qY4jsJxH3gQ
DhFMcmNLXRPLM3Mr/3Pr8JOcxkZyjYn5xSpoIPBegk1Kw9kpESeMlzC8xpHHbb40lbRLy9/qvKhb
hOvkFuzVMGwmaW4cI4bbMHClxBsxw0GcqYxQaik6lPSdoz4KgXpDV8nK/IuCByd5eS7ZxqSPHIND
VTPnvVdowJH1G9Xuplt2Guoyb5R1l7Hq73ynlstfBt0anIBBcN9wlEOpEBLzDEs49zesXIh40fWB
4uhAJUNacS+Py8tIWfXF3aK/2z+lBY5sKuyGul40pWqPsTh/cuJXr+OuzSbss9/N+gQ5rYnGp1EG
sEMbCqQ3is9m25p7jeKvlst4Fq0G2J/pqdTr62I4M1wUZ4IhDsos7rywNEeN/nb+X1VHAq23YX3t
U1jf+Miq42CVZZNUOLldsMFppAAN9sr4xX7OFRTC/z28J+SuUBnJaXBqqHKaLUVVQoNWUtAGxexc
/Nbuj0pv2sTcfd15698JFP632VTLNH4tikSi48NOTl6xQhbSW9PB1OhaECHx46UoV9y6wPktosAk
g+Y5A7lVCcdbavJeucCs2JyeXlHqpsYqgjHSCrVapQH3XKdFeHxDr4m576d/JH7uzh1NnxGehUlJ
eT1/v+4gmb/3VHWEH+SA7RoBOh4SzkSpupi5LX/ECNiWzfLiUPWM9igds/qRIACg9ZTnEJadd2sU
H85ua2992TsqRTfWYaNk0irJBLXwwKwxcUXPyP8mH+id0b9j8XBEaJ0tLgD1uYBQe17V1O+gTMOp
wxFpq0BinzzgyNiIWHJf1rXl9PFiJFBq6K5czD7G2uoD5w1Ip7KQhXjpTt0wd5/mppeOiEA+P7tv
yIdSDSdra0PKRNuWOwbdBiNkn8NAMdqB4ohz0mHI5m98Ej9bpA3LP1+pz+sBWYcNSFuFedaB9bdU
MVYFYRqOD2PMVRZRHxACsRzBXH97f6+Z2DtZsYmylMzbPBhkKGk0eMmf1FKM1Xm9KEnKzL9Gg9O3
3HxfOhb8ejl+8gmQn3MPidFj6nVDn6DF5cTZpgXpdlgZugFzPLH3M51ZgcBMG0jAPQj+qsAg/EOx
ypgoqSz6oJRGJqhrqlEqMd5G/G1scpo7t686kYfHXlZU/FTYEK41YvyMCG6enK/lqyC2yVUboTkR
/xRzUwSRgoz04pwQIr8RCD+RJcXyvTTZjz2GiGSHzvLlgYaCtW1zBgJX50Hr92FqqE15DaAmCbn6
Ut6M2A//JI/78eIGwfQ5esTzgO81Mb6ovK6qi7UAJI/eIaf3ElaUGvCJ4VUz01Hrs3oyPGP80Ewd
tBqIE/Vz4YYnl5ND2x9RmZsztbd65ylaWnCpGg+7mbkUWXPN2loVNnzDcS2w3MIW2Hhgf4UZR8IJ
RKXcHZUGTxAmOFGzOalvE7TyMZLGo/oXM9jhX3WRQdnDZR1N+zUHrkRq1coZVurwPeLeikq+ECgS
gJodhJcfD1qgg/fqkTkwXMUO9KqYo/elvyBwItBSyV8jOocaqLE0V3DwOELeUpSetPN4cNLejHTe
9WEJN7AiJWrvmY01/FuYRwATC/gUl9X++J+I648ZnWGHi1LI9VKSQ36ew7ut0aiRx4cnNTwzJskA
htTBh9sbG0znCH8ppizlNzZVVn3Fgz+9chs3LWBfPo6hMrcgLGdzok8omjWM/fMAm1L0CarYoMh1
UtHUWJTK1LIj4tc3LwaMZGhleiIuBUgeP74JBsB248r+8dT5NB8KdoeMGXFF5LMESHcGiPGbnsHV
hbSXpfBW8r7WBJ7Agrz/UMkQMOJSgtmvK7qykFnoGK3XbSQ5c76vl1wNP8t3bVMD7kWdzJV/I8Vh
m4/2TyqgmR0if3bR6CmX7Gafncwr3AAx9XmQ1Ea0YSO1Lvk6EZ34ByP6aIhZ+sH2dWVhFcK2qkX9
WxYLDbXchvnZu5mFPxcFS1Vg5o1+8wKunrrGROdi1krpofjm7Z6Y9yyVKx/+rfaGVjlPR6jMpqWz
AKbVYZXsJ0ZfUKaHzZiIRgwkm7jRYG0hE6UWj7SJGxZQuDmhjAmugfcaBQ0OaWl8qjWpRZb6fSFw
JEjqoE8N3ikH2NKBAk2MjQ3DT2nhUTcoWSjiIDWVi4jHQce0Xuvdcf9tHCO5mSdHJ3XOYBs4zKVR
DQCHkCapQu9/fXqYZ0FM8uXeb+YTpsOCNBAoIvlDAnjGaHM5w+/jn7FZc0nWyMaTK4t7U7JimN8v
sxRL2Rb+MnPIWxiRuVxAjwJe3V0GCsuSwP7JPDU/xAtHa8C+nNxdaTwXdBG39DqXX1p/byef12+m
s0+++xuyjfuEUg+7MSLzePZ47IKjXoWOFLptBgkXszOlQ4POx3nAqej6VVuag0KNvJL8hIY9Vzxu
YlwXxSvwYhCjz9r9zXShiQkC4MhGF/Hrw/hmG2kZP/KFaWMx+6bPw2oqm8EREmaLalTL63A1r+YU
CqsyC8m/SPQ225KJjtSsVhTAwesIIO2izz3/so/zu/H4lGgF3Fg6FZsh/WDJjrvv+omgMyq92E3O
ZlduQUJXysxufoNPlP7NIHhzW5QbjuaaMwakbW/yAy4ukgYQ/S3pPmPphSIL4jlCcoBd/oHsHBrj
r1ha5/G/4xG/KCv7ajHlrSYTEUK83liH0tLwiuR8SPsqq8i+5WoZtBvmB1o3SBbV9V7AZ5n5h25A
LDvQMJccBYTGxSrBiwLUAgybgmCOEi6s9Sm/CpRaDu0QYpGInc/dpavTs/wkIZ5S5h93fWmgQlvc
BpGDP1ZdcvciRWbiHoC1fXkMAaaN6Rk2StBhk/9JXpc2l/8es/CTWlopnnnGrXymYvy5vNzQBAIB
WS4uZ591kTz2vtNv5sr+dw/YUl/I0uyLY2JSNLyBHsDPPBZGKrSzhJLYT4LwqVuzPZW5edmuahdr
br8+9c3LDT/SiLp/oQKPsHpQVYO/Fe+aWyIfVFjWX6eytwDQ1Rmeqhwtpph6sgLOWSOm7NiZmVb7
zi5z6Glj5JFxGrGT0BAxJnp3VNCV/+ikQrfHD32nqtJeWPiJ38KZvBgNyh+m/+p0otA2Bl2qXOEp
TvQ7Ri8D9masCAEbeTXhP19l1c/Q628Wp/UGjfaWZrahW9reWtUEHlUYukUARs91Jeh1RfYsZVbx
hak5Jru3lQ/v+a4Q8Oo7EaNIa1pZAFaxvic9XYTOh0LslixNZIwOA9u46hq0deEWAjO5N14yB+By
6SKVKrYvke0qAn8UehtoP6IZQiD6xPCEj6CxmrHvfH3DyG6OeflUtOlK1sO8//G9rkqDUxIEDAx4
dv+x6F68qNBvr+amoTEwTCJCYOJ2lDnkWPDGdGONV16i/1heq0IK3KDkIIa4IDjKcDQIhLRDoOn1
qWrOJMhM3Wop7UuEnm2Hk7aRwzH8+yomIfnC5V2OXIRIEhpJofPWr9uXPqBrEw7LS0inU5B1i5WM
6nCVXcBf1ctWGcyBHbBnvaI8aGwFDXfYmH7oFb2op0qLdYX8sReTXfh5Zktxxb2IvX8w9k8kmrMS
3PibGaXa+JKFMw54iP5u6S2/PHy82Z2FwCemr/YOC7cyzid6KA9L+xzO2KGFJCEgkoq7VK8bqK+2
XF2XMWZrQfRRmjRr56wsVzOHLtZ2XtoehpDpW9PgfqjYpkjdAK+JcSVXxhWydo/xn9lHQCGaLK4t
BEk0rzdVcxR/GPPzZItExrnVFr4XdWQ3QPs+eeRrVHMnZi5CTShHXLZ4V9CZHlQMTTtwBGV3odLX
WjHM0XEWfWUmInJPrCeSb7AdxGKI6J+FkY1Loc0qptBd6mxb5Uz6LJEhOnxVJGLAFIdFyfw/utMe
FktdaKmxbPIQsEdzIRm+ySIjgzkskP1mJZaqM7gybGogJqyvl+nqsAvyDbsjR9PpPUfU2KHz0iIR
XOW+Lj2Zk1gZuZegt+3Ur5M7UBH3ZQ9IGk/zEeac1bBdic+Ude/yUvZVWXQR5WIY1AtEKXX3PbiY
MWuHOp2aoZuDEx4Pa9tVXQ6hliItLFQ5341NCVvB6fydrMWGzt9XS8TjQPiaUfdpGMKbxUkopx5g
3OPHdy89WYk3wYlJRBZX/Vx5mm9ikgZhjPIeHO870euKvM3Em4QRCp5lyTJHXVIGlfUzqD+PXh0q
PZhpr1c+VYu65QGveoDfGc02+5wKbRW65+vcv8UZXw/A8wCpL1DXDJxJ48LGR/0zVVMJQ9BcrFT1
2a0/gafxO0BI3MeNsUfYgPmhsNtrdP2x3vEyazAd2r3h560DfuGI9znRgacAOkl5uCOTUVHtmGsl
+1b03xS1N4es3d2YtuMtFSTUo0NEt4vajyhhUqZokChb71U8BWpKAre/V67M5tMBSeCVZxSdiNxL
Wrk8wVX3qsx39cuphjO6R3g4O/sawtP9frNZMeWQPRTmBaCtrATcqYB8jZ1BOHqYBtDHjsnLgjH8
paxKJoci2ok/eCrgsL2HRFB+EL9kdhRQocP3XkxPrhz0DJ+lRP86dvx4ik6amqneo35OuHyUfUlX
DcrMRwZuVrag5fC6nFolFnb7axgdMem5AS3Fv4ORFWvVXynPUdaB9U4i+K0sLMCPFJ/1vEEq41c8
f9dFL1nDw2jwuOW1vo6QLJPkS+qCrvXLaGYbV3TvYFUEjSeezkveDhP0pjHx3L8Yt36viw45Z2fB
KMTABavNI4kPHd+mpmORIAIms6KHOdU5hOKAEU3pjCMQELIIfb0pgk34YfntTksm9pWkpt0CWpHn
+6+R3/z6/L/PVpfxRfGg9QYvstLK1y/DF4oksU4g8GGKCCjh52Uv1VnaNzQp+yGWRf3d461gUnhc
CD+Wn12XClpFO0Q75U4C4irg8HIMlW3bMgDOUFrCYOyh5rbHp7gRvvP9slTGGLKNcbFTyFa8TyLx
17F4nKPT8QwlDP3OOHJL378WIUSfcFhM1QsGuT8HWcbQVR62uEBEtw3XY90qonaAcWezNRp0vlMd
ByR/Snur0Sat1WWNsSMPF6omRBTmhtQ5avZt8eTt/sCTvfasy4EvWcVl00Hsl3yts/mWJt0p0lwU
OP5TNHyVAjt73EJEkeAndcfNAbZBtEsDbA0HvF3EmD1+Q5k7Az9D9NIIClj8ovwsUiC/1RK3L/Nt
JiyLAXOJ4lBeZN0sRlVmnQYS5TPYGh6LH825g1tAKTHOmsdpnFlaWmGQCoWH499v0ef3zlSymj5N
DWgOSkXtYukYSVEDRMpaKGqTYU+N++rPneojU7TW1z3BLszONhxlMMBNnlX9aOk2BGA+5hHThtpe
QOpUQ18cYMPpHWLWUwFsgexy555J4q8xKCaDxO4OKfi6cQZlDNgsapuM+nG/f/zp5QwGFWdfyl30
zOM3HJcQ3515mnjFdCusNiin5L7KbF9EDAkWlbcWZoBD7C5A+Bm7we5oZ4aaKM4mu2IFvScvoeGg
XhW6y6khJu/+usBI0yMVjMBrZX0imJSbEjM7t58ZMsHWyAfZSE7jncDueDSQaPVlT6eqNdVmF69+
2emUY65No+iPr2Oqjw3P676pxqZT2dMTd5T+XZTxCoAPw75+rUq2uqolkf/n5AsEWbSbgn7jPzNh
3vnXHIEIQH/ZJU+MlUZWRKmPYZ+JTldGY8SEoUpurVa1kqHvbXecEoDIBlmgO7n3J6U23tIS7fvW
pdtzqJfDQuAYE0uoDb5PfBL0zTJc/27bXhx0mlzKqac0OmYxvclD5b9G9dqPTaoJ7hIMbgcY/9t+
takHqM65ip29I1M8jXqJMMLB6nFPCu8fxx9XHfNSfCP1iRcw9aVhsUo+9hlEgQ0FByHfH+rvdwp7
yb5qXCJC3lKmpFR1qVxvUd/Oqf+Wr1ladkKdKQzBTQDDtHyBQ80VreyPBx4rDSnueeKdDLzF2CYm
qH6WIf1JV9mR82quzJY6CD7EC0ifKMpT90f1TKBcmwlcb8kbofNn1WJGbOLA92i4IROEa7V8g3tQ
zMHg60nqw+OwxgBxGoJOpxsA4T3iBZsC684ddcy0GWw/qMUNwOOKP26ki+LQAJBbC433SxbRKk6X
3Q2hyNNnqxqWBXkl6jtUxvcvoiZM98NFi+95x/GbCYkd/HcQsAQf0y3IDZhCGn8pCTWWvNClwjSv
S0vXdV/P6L3i0xqGZchvy57ALRAFv1CA8QHWy3M4kFS0wG1XPPHlHaIcz9597TY5YjVHscF3pCx4
4R70/lXBKhwZ78QmtbMtbcZH80/WCkRSdUwjZLh0V7YeDyffUrBmaLpJgQq+5E5GVZ5NQ69j9qRA
SPa64vbAc9eJIcLdaj0ApMZHuE/ZUjlm2slYpOmF/oXyOez/aBJErj7tvkvCwN9FcPFM1gTJm6VW
6xWaKSRLi7Jc+S/o8PuatPP4QSUMqvBSpj4C0rj0y0lg/RT5xpevlnhC4PU2Qcd5rQ5ccRc2lBja
xtRxmBLcGs9VLUC+/8jrWXwoMtuMkX/63pVHfINDqaeXSspORAsHZUwi6bRuu9EvjIBrNejCdca9
7gsWKbUDahnLXp/5l7zEd1KdxASfqp6TUexA65I6GRsUffjWfvTrAw/2aUzsE5yA5EpuEwp+wJgq
KG1Dt/SRqQhXBKzR8pV31rEBKmmK/hAy79DhZ1GeSlt+KfbUSlZzf4B1LqueYlVKAMN4hd5I8xKY
WTEHEqDmM82PQJmRDgu1BqepR1gizrKcFFS6eBJqI76OsNmExFog6RBtqSUTESEu2IX3hW5ScGYe
UpxEwg5SFxeakGVVU1ZZaUzqaVw2UnhPD0d9lyFwa2Negaw58sOtvcj256h/SjnkFrT6BwZdXHEQ
7FUApLS8ZJH9mAYmq2vl3nnwuV0XjC375KeiuFDj8VMCmCDnoINB4uWbLXpMpQuq8aCuMs7C1t3D
gM1LPlnrvLzYJqWt4tXnevC8pBYKklZjNr7P9jcYAlt14UsT0XCJ5m4DgqtfDLmWHPKO2KfnhMHa
/D98CML6bKfW1hvm2wYfJAzSD9SbBTl9FpQX2qWYPPP5gehj5aqIC+2MsMaW4AEQl3J6n/M418hZ
PPjcfNgdGh29ZwI5bZWt+spJCrAOJa+6VEdy75dBNZcX0pHy5vAp1SmvOogzFgbTtoHqXY1nI6S6
YLns7XcdY5DV5DOeN38S0jjXcC8CgCaSrsFFNTYTHDCRjH4A6+NSuhx30coXWjtBhSNpYMcGKsMI
Y5EMyIdF8d5WEq6+2wnHUDnGtC27g0i9qFx9MI52krY6ASmq3pzuufnpDdgu3D1GWsyuEvhr9K0P
GYR/+u0Z1bYoJE4VJaW7bD6H27ASEw5iVDe+7IJLmny2QUM9kNUXDIiD/SCdFzGSQubVOOWAj8n9
pB4Hp4jzrmjy8K2plaM5KWRgKixzB76IG5zm3ApRFouvMt34T5tF0DJQ9ZHe9IpU+WKN+mF5Xkdv
oXqlQYwRxWCDJIbNBI6xS0vlZexg/NFEYh/p9O0yU8JK2ZxLku+Rsuhn5vRoivyg6v7s7aV0+V4t
vgt1wA70nLAa5pSn5AOA13oRhvxt3lHo218QPfKPs+1fk+iot4YeaHw8ZRJrWnqkhpECG+y2rmjB
LWPEN8FgGBMrbDHZmicjxmH3LxNcGBjPHJgcFZXSCY6tTF2z6vPJ0qR/RDoTGAM/KdOa2rWZ9DFH
S1rpPWDwTYEdDkR4bQMgPdrUQz+IuUaynNLgrv9QxJ6RGThgUM/aQSX3WLcR6/ZkRBs5wJuZfsyq
jUWATr/AHj/p2R9q9qEtzucKH6aOCSHhIB9evs8uZTJt/7BqAUhIYXAAoxHpFfbnIBWMHcZ2/ioX
E8Xpsd8ZgDkSivOMl3mHbvmiRNOp4OHcShb4/U/n++TsplgVJepAbNp9ebM+pJeoaO2HM3x449PM
EbbsKr/fW89z/eICOtgcKDKRlwS7jSPfj2iwfveS+U9T46Km48HZEB/Pho54FNNddeOEBh+lI4zX
/mjMEAa2JsMw12Gqj+kOx0kEyrio5MDkLCDEDxNCq+ICJFGiHUtDm3bmR389bmIsiLNlPEwvxYV4
F6AaclGnChwsGvuiS2tex0LHEvW/2TkwFVJeAk30Kk+8+sm9ejEISD9TfKQZLVKU4bTYcwxL/oRT
F3YndGHGBQZ3JTH5JUp8gq0NBW+IttaPpA7eGigLCuSfFWw8wk0Hj/iac3FPAEiMGrnVfpn99gXP
6YiUxvUd94Oe0ypEVYyEua+psS9/DfcDcHM2aNIjXCSuxE5O4stZt8b1+168S7crVO/8UOvq7KVw
5jglEYaKPQbxlZfz9bEpoV7koM/MiznFfWKvKbADAW307p3D8wLCiVQT0gpQizyudkS4goKZm6xz
zbKkZiyI9g24arvjEoljUMw+M0VSTGSmmwqz7x9vp1uvXC9DraF5btgM3SsLMwMKIss/uBC4iSuM
zJK93myTiNvMLUSUOFr1nQNsqp/RlDdXuACMTu/NCNF1wD+7f+1Jr6/bZFO3Up2sCP0asDJpNpd1
f67a8JPpLrrPvBCeI8HfKkfAXAZjrGi5HUgTZNI0svSYCbnOXIfiLELCC/wOZPcyyWEH7aHr1IlD
DLk2/o4FuA7pTxFRPvQMChlcJV8ei6YBsERy8wlIunAYG+2OdHNL7nqF6OFgiDW2uaLaONgrHKLZ
GH6wB5gNlk5tfoLEcLdda7Zipcx62HRIilOZ51rV55ZWhYE0Fu0gnt8DKSwh9S1Ni3BQ5+stTNmt
o6Ndfoqo4mgia0yOzv/k1sQ2kY3eMygqGa4DwNFoGrmOGNyeYMQW1ApWzNrsgaCKeRqLAUaSLeex
LoRlcRHkgvzqiPMY4vWBlHljtznNrLn05dBKBcy7BaRB9prENT/Q2KHmfhISPtt3BYrYivJZX9Sz
7NLKzi7BciMSJXTFxC9slWOHymupG+jQ9Z/xeRro+BBUKJh/ygz6v5STmWw1tme7zSOXfO6q0Mrh
NwwWumPKysXlBm3oUWvhI5bmY2N3JCjBJXlkSB42uaUtuYENioBHqc3xiPwiamQuuTSq2Gp2/GEN
imfm6B+RH46nzDtzCK9afMigOGijFM8rz+81i2b/9OPUUL1AX06dN6V77pUIimo7MGKcb0bZaOft
JlOWfNq3OSEV7VYs+g7YmnF80DKDmkdTKDxHAW3iTh4Vcjp9x1z1Y71wvBpm7v67Kbht6MNXQDvU
99nigxbt7bp6GjgA/64XncVrnKn/rjXf94GWC3Inl8Uv9HSvv0b/hG809Cg7DhuoE0xCwocXvuR9
KoBHSwcOhM9mH/A9XP23a8TsagmIJ/qGx89x+EReqU69GL11mNlsnSQOz9M+AkZqIkFBWMUNfe4r
CAXGvKwF3qaLUAki5qlMoVmZWaOSTj2vGSqTGhtkrHDjAVIwxfwxrm7MuOwLe2HQGUEtDz/ykQxy
aSSmj4LPJR6xb0ZT5Nnkzreiyddw1r4GNm0NSGbAy37dsMPVwd238aYelJRUITpm6jwO9xaY5po6
TtpasrWmzqLwbxMJePfXSrUinvktkR872EutXulaL0vGRkLusfvDnwjQdyBdev3wCfmOb7gRth/i
y2ueBdJy+q+ZMPAp9s12roTVbKkGvQFcAjO21oEZ7Qg6RWh7TnlWVNK9qI1Dq8tp5sJPGPViTGUU
ROn4wBLHM4sNANossXjXuMQ6PKoPRWNnEK7iwbWKeAyvfhwStNpniDNYvEqhHdydfdjEFzecVerE
+6l7K4H4EFKLzUihQmw1Q+/QmJDXcCgXWjA7bE/P9x6kng1xx5qCNO7IvsR2gLsBNrc2E5q6WT0p
9hIkg/1jCLU7KhPt6pW7ordUqP67avsd1V/GkQOVemsvCgbvpkq90CShTtAeVa055/I60PiwIeam
VRO4kuJST4oem3+quwBRCu/vmANB68JU+y6RcCXM3SXFlV8SO9knOU2Go/mkoC8euyuX9ce9l0S3
eHOCwKaja3mbBmjg0WJKFRvQX5GK/NMgm4Ex2dGcWbJuPqSQ62O7v1OvHk00PHuce+5qsii4hCWj
osZ0D9fZTEOr8td4m1aweO23/WuwiYmp91AhX/6WgXeYwZika6Bj13C1p/U6tRqUWUBbdVlxyQ3D
IkZh6Sn2zOswyIqDiLeHEHPXJ6UrJmSVSDpYaZGlsuuTWJ8J0bwO1gAzf6jVbAsQUlQCJCeIyus9
+v774HxuCBSC+K5oeBV6sXZxBbiab/biHJFQFE08y+4xVLL990KWE8LUIXukVRUErfiheybhr8CW
+Zv18JIV6h5p3iZdSvGlhi/ygY0BKLXfWVIx9BXsLwIwdv1zJtIaz75qU2OgW13gvHhgUJN0G9qB
3oZWXVFtStGYvpbcAZCNCJgZxp45sl/xVrGq4gQcTqGCsgHBnPWXTMM6QerJXAMddUdwGLhLJQUf
vEtdeMNn/pZtqudvc93MqEAgjbiTS2p3Q1ZOaB1NyDQD6RxdPhyhQw3UwqYy/LSv7t0NMfuUfcI3
7Y7xa/G6X1wvItMJGrApgPcYmZQ0itb8ilMDNrhnHHxhEmAtskRtPKQ/onrYgNXtq7ZMvpOYEEoU
vyYW30zvNWtHnXFQr2WroU4u7CTKKmgbWU2OCAoC3qYC2eQZhAiAP2EGl7WMLCrCCqUs9DYyOeHZ
dTwiyTbyHjdsPx0N61YNVriUKYLBZKC36u+GrmNHButEVENuZC2zniiLBJCnN9grmqxYUbo2Euj9
FJX3et2O9Ul3S1Yea6+XCofxr/981t4d98iR+iUuJnGsOU2kgVwGkPH/HP7KyhU13hSyPw7ndl8g
xe8oT/RfPPI5cF/EKUYtlt9oL5BinBWRbYaeywC3xWUfZ2L4ZYfP9CQyThmUvpFNEyZ40v7O9HiJ
Q8l2MGZ1JUoJWjrfB2fW2PI1PHdOim52JPqDIp0z+mEUT74OeuU446G6s4a03+YKveIcTkhgKXNP
lnygIsfY9vT6bPtSW2KG360lbdJqhB/3IXuDlghq9ucZF9bV8c9mmxLOhTCLXI24nMbMm9lStjoG
9UdrhXPcHrFPM+i+V5X/qXd3dW8h3uv21O5U1Un2OyGbMt6tHrBquy/90vwQR8GTVgijLXVVuGxh
Ut4rOy9yfBn2NFT9ik7vkZBnYkjmLeN2L4rCK2Dp0zfEQNILSXL+kC0kJpPREzyeZ2RXaJfCrv7X
1Ybbg/xScpc37NNLfCFZW792V7nNjTVvgDnKXwKnq9OYr6BIsJjui1zKRrh/g2QpSyk25WIOlU+2
BzeiMpyrbQgGafAXQjhfAP15fBqZeeq/EwxBjVCf0v1JKcG6k1mEIlRtzT8dObMWPt+VT3gBF3F0
2LNqJWS9/l/Cgd/+VPe1E1ZEm+2v7igeXacKcLrdp05kIcpgkW3XKnYQz6NLocIzlZilFn6KDSzk
eWp7LqDuOWN9iglQkP3MMCIKULX2iKSnLhS0HLqCF+VhueHsFDWMlNFBRXPnM0OhhJ6hgffWQJZz
DEDAMbYS+Gkx5RSjI129QWCJVgXmFVNz/4PtYhjqTTiw+cZ1TReonxh96Gz0N+FkzowcNuLW4zS+
XM2Wq9PNo/3YI1DLZ0Iqd7U6w1e+1c7RQfZaBYl8EY8WaSiA8vTGdjYEZUgZo6owr7cTdSEN1RJh
dSkwPdDBQ5nruD4fuc5CGthaf873fbEPjjj+k0/DjSIcOOF/93GQE6lR7lRsAlhxekl6/+ZwTLQK
XJinD8gM7dco4eLIuCtfPRf1J9snwqM2w5lIj9ls6GKtTDx+WmmgfPS7Hp4QXkMRu/ZvvAjpfbIc
pobch7QtT/p5kBXevhQBUdIhroPbvZ8fR+zMW/TpRThyzWAxs/ukUVzuxW7lg9KUxSdQIGcR2Bgz
lnsmoqQYuYsq9JnukAR2ceoJp5kgtOUajXNuZhvAb/9Kfe5/SjG8TojfgxaZffJMGG+GNjPpgapG
yguzq51/SVIeGMO6lco+8dRdmegNxARefc7zSr//FKlzpxbjgqBUfdQfVMexTqBdAfWc08zJyP/3
4fIJOyvur9YrdNmPDjJxb+gGU+DPD3jUtb5lNcqEZ5/xZnRZvCazf64SP/PiXZ+R3rH3n2+jxEWf
nA4ve2EmWhr6wW70/IhQ8TXBipVvc+Gubq0dmI0f8V/guuMEEmpwyaNhMLUmBFmb6zul97rqOQto
BOeH8gzSdY1JPQECro+zBBDbuRQtWRzi4ZFDI6TehpgKU/0xF/pjrErHgLAKOM/xh2WEFCI2KrB8
0oUmhuNYPZraM2E+edGUbwYLwibcpYz+D3/tgkowWjBILqoGKKSf0h1mMB0HdMWT04bn/3HkH9sj
g5Dg8xh3FSgQvGF7MLTLoyeOVA+I+O47u7wWlFRaJL5mAoa4jMAgaabtQDdwYVGuxSixbLN++Bhe
1eTJ9aqG7odbGh90zYw6KCNPgIwDO1X24FgSnEv2shDP1eVbD0iOpnCdt8q+Qv15uhRCwTBwuie1
hLHEXfM0bEzgha/vKRFdeSQfTZMGcTwmn5QK+R3T3khytm0Q50FSnEgNKkq6xTG5ahfUr0Rceb4x
4THsYkniHGroYFSAITYW3OgcRAQi+EWWJLYjVqulDgDUL+sf1UFynKA6qaGuCYrAPx+FxekqugTq
v7GrhSD7tObaUz13AYkaQvy9YRzsK1AbH+IpjuEdnjTOWAhbWP/bWiSGoXe84KcaUW9fBX7GTfEN
VbLOnP0LjZNtB7vnnFY+BIq2ONe0zhVOX+DtJVU+xPq0n2RF10PjI5MGaFHrCCbrLKMMo+sGEkOo
N5vp384LmZsWWyRT/7R2Uj5dHnkMtukf5wZkjgUGdT5tl67g2T6iiOYCiCjPsqwiIFOF5JsePHCE
tw09BRkfxh0rMNA/gkS0BUoyKKOsFzV7rgU+6Vw0yRXgKU4LnC3s4DbDzqs2yolTPj4IIaqqj4yj
l6kdxayE4DBvbadEjTNSCNKb4ZM5RgXcFPpegR3uMwVv7ygkJDUwKlL9KRjla1etpZMUWVyGAxSH
j0koZ8J5IvdwaL2nn0IFStn7tFwhbeqBDgTCn6yX0U4NAH5YUthQJCL3RLs/jbUwOQBHx8a70Zbt
1TOmmfTRnJcV7oGyjB4fjvKDrqkheqA3+uFYmPm1tqFVXLpK4sh2c8Ks+Ffx8Qt0jFbUqYPe5GPa
pDnG5h4h7ijcfmiO8eX5R619nhprNIoQHnSVMUOsCA/3qPHV3R1q3XHRPCqgXfoEGEDVodUup5Xt
6LazO8Csb7UWTJ7PaWc2bpykl5l50yNlcjUTuG0OBuSIgkY94oSFDKa3L7Y9iDR7Xx19cdD1tW38
REBkM15ADa8ScvO4Q76L7sN4PBM8xJ2reGKScl+4oQvXw6BpVZjS9W4W5sN8hAUgj9q6LWpnYteS
WPRX90WDWOuiPmaqH02eHYeAt9OqGyEnrbwDhJQvldnRQIihgv2UfkYbs61iOPgCesijSMQGVxK2
dO9za4IoJhZdi8YI0KObjswhG6plxeNyAWI/vxV3kXVFcm8XQtHK79Sa3jMRwFg9W+FeyMkgMsVa
Ll+8fdzLZtkozBDfKBZts8VaG7QrUsn6qFBfYZ9uhuWIygp2xO/dH7CcmdvrWWWnTFMdJ//j3b3P
2An4K0yfmo5zQBMOUCetRk3B5E9k//8blqmllKDKqPVY11BOH+PCRIXFkACmIfARuVUfxH9O9CbO
9RgFzwT/K9uu1LxD4/rNWkcmjTpj57MYVWeAya/G/Dcq2SBUAFtoV+NyjNqAzyIKXsAywZTdnKk/
Ne22gs/bDY4HTzQdeLlSQys458S+Oe+ilxc3uGYZDO/jc2dYe1AOa2VjzDkeb65iqtMF+boAUuj3
fjT+9ma0qUHl0G7kh+Phi/jhmDfxMhekefRiRmHCDyc7MQgVMNIwrBP5SlFRVna2sPfSUBbhm5Z2
C9xLxKACqGrGHiyRRLKMoap2fk45PJfY4wsqjB32Xp8XsGHnwl5FXRyKpNmapoaTNTp/ZXy740Hp
y9jU9u6nq4//qCEsY0DQABq5ZT5ICpI6MUqYiIp2BQo+pS1I8f+q/7xmBB8RYd3w5/ZKPKj40jbK
8Nx7TkoGfContYtHmKf3UGmv1iBryhU4kLXfyX3RwUqZ/aoMYidmVAJ2bFnxNT5nNCS4bwyhQZB2
GZp/kSKcwiLTJKJXxA2DQKrLyCiHZyC1xoGTd5rFPcWT1LL5IMNGveFNL5BeWWxbYX3PaWsvNrrU
Opz4On4u98TYBvj60dUmI4stZLTYSUFquQc44dsYeJPGnpwu5DfeOXLeRV5L0XiX8d7CyIVHe5k7
TO7kCeEQgaKn4UeBNPuUm6P+q7XVDjG4LNeZGY0dSrRU2KzA/WkAh6rqu1JRP+z7n5IP6r0flyP5
2vD30lQS5Z+tronZF/Anjxuk0MgF0jKzxlfy//ChIQoJDoUmzra/M2Sid0EGim1qgzYOdqJL12Wi
CEq+SiwFXGuUkFlh2TqgAb4Yx1gp6f+ridWN0x56AVDphV9cOXHCgBm5vABhHlSKGauQD1ph9PED
clmS27k7CX2wEWeJGhPTnkPjIw/s3Calg0Bbab8T2F8mOghT792ZrkZzr1TczqvP56XxK1nQaIXc
yQ3+wKjVolL+rNGSHZWDMNtk83dhi/g+G5XwmWRzMxBo5whzhY5q+UxkfVxQ2f/P4hD3tm0P8aW9
48dRoAuDB6OG4rKpN5H5/moP8GpTIpXWYjxoOJqAUvkXGLABWgE3raYXyIsZh0I9h+xakhDopgja
HhWj/Ip58Rrs7dMLoOsuu4Eysgh2cebSp+6fL3BC6aChOK5XSDPMIL9+KwgGnY/q/TVv5Vz39rG6
/Ke6JZBWZjaQxGee2r4J8uOGY1YOYBhbZLO2NCJOd0zboHUhb3IBxl183B7iiunay/K425vUylnh
H2VDXjKZkyaDvSRBdAn4zaWHNrXPFQPeFKo7SxRtIKyM0Ze2egGic1TBUyi22Cu0i9F4ZBmvwffb
3c2wOeN/g7GZ8f/SDJWZMWRqYaj/Xkc9bWiuE0jOZcbXXoFN8zOUsuc0yf/JFYR7DPTJ//QaI9kb
FKPdO3rZ1sIoG213N+JgwBkBNSBmnZkp6d5i1vlUs3WC+JWRh2mVHO6Tq+x6g8+nOEfSo22c2TxI
VsP9RX9NGGSmMP877Syd2/goZpij733g0bYPQ+o3tqBeLi8xLpPQPQBO09uWozMv8dtjRvi82aXV
/ZxNGXjQSFJo3diZaeKTHW54+kKcvzlfN7bsVlriiZftDBu1wU0eCKuyIPbfMddVWq6IWKCpW7ft
moLuOeL1xEixUC7UeES53dbTvFARGHeIhfr0FPXmKJiK/iimSMGLByn2LFnikEBHP7kgycW7iK8M
Qn3PWRTfWS8dlbRgXGE8FRY8WVG1X0dfdcMSDmPMgCx9WTGdTPXS+URJ0MEVzfD2tMdNSh6492vY
BC3RN9pnkFBUWel8zLin3CQEBYu9xpPNITQP4Kkbn5howJoIrnm0OhsV9/9fVaUg33O+Y/6bkHbE
M8dhYgxIrINs/xUQsie4X4XbbPvTs5vX0IYCHd9geToMJVnZtJCIRopCxr6eIABcGdjKRgTtKL8x
iqVkXVkzG52mhZlpcGJzdTXSsCJrPGwi+/3EdOCrm3zJLzfGI28hGLmSIq9Xe8FM7km+Kkwgp9MJ
mA9TKZtc3KzflpunldYlqQY8Xk+cvun1Nf7vxYZOqLkRyRFF/sjUNR6mVad8xTWxAzaNkl1DwbzN
anS24HO3REc71D8ppcVxdKfeVLmbsmxTSqN3mx5NtrtPa1bal6yjyRVpGhocU9B2eU1VgHFB+unn
7dQOlY4kS6BzndF4qAJbYyDti65rvxW0TXXxM5V0CAigCBYRcZ2UaixvF2ZfuVZ7H34vU/py3noc
hE8AmPcZrrdm7vyqLpMUXSZFixl+yGJCcsYptacG9Yu4z0Sxmbdisy1+BYZ1BTFT94ZReKqh0Y3W
rcACh1Sg8CakahupzRwo0AiU34sPBj/bTHGLGEPdW0xAlItcp8Sk5IM7M4lmt3oVADu6JGmCdTLT
gNeHlTlVF1F23Ih9JYjVrWGetl1/Xsi7PY3a5NwOCmZDIFbGZxfs2rfKDQ127fQYXt3JqCuc1uaH
3u+VUR56jkvM1QG831ubaclygKZ26a4qHUBVq/kCd21/UYkgElkb2Q3PJY1UtZna6BNlbSZLEd0+
NFKR6aCexzqbprJ0Jo8UzgMdN4lq5OUZeyhnAABktIjBAPtjHVvfcQW6/4cDyyfmJ40Pcretl3oX
vSe3fHIGYTPQmOlM0cd3GGCgSItNTyf+6XEbwmJt2Vs8UyYX7G9taMLWo69KpMvrsTEE7MNnvAsX
ZHYc+6IIy7TFBMwqs8DG/1qLno+KeB4LBhqyYmBc+xOqXkdDUBSDPEiZfWBY1tggJqHrXs/xJ0qz
5sxL00m+2GvTuAt1Gh3JEyi3DZO74FaVDnQ1698aQCnQCwulCF93v2mBYOAAar3c4CsOBLdcwrJJ
pmKVuBWytwWOsCgq/AxJnvbk/hxRGjAsH5svlkIRkcpJ+uNK9cJEaqGUXRs+44NJeXad2X7oGj4P
Pjwj+4WGSc2nNfMYGV1YW1Y0C5qf/6uMUvzA70e2pquksZf/XVnJLqCKBMN14onlhdLpNubdXhCW
O7GQEL+kGFZJfckTTC0xGaXHo8Oe8eOINld0hgdPbOkd5LBisFw1E7GkEkE10k+78Yzs0vOC7A/K
YQFQiyZzkrvJV+QpdZ6YSWG71ZeiwQ6KhIlpsV6/VlRDu5t/Xaz/sb5/MV+YzbJIViTU0YQERsWW
M+R49SGE4aeFEFUCWWLsTSS+MqBJZTOTACg5OhDfRjy+FjPaHg0E0ORxgAH4wDDxhtEIXRTax9Sm
ancf9DAXZ0Y4K1Em+iWFBTsnx8+dErR15UulAHt6aZB64/w0B6+wSABXgT+qW5rIRZG9rKiUGKsk
Nzy4VfPpX6V2KgdmXmuiSlUaZqWrCcXaETdnobCCyKFRoco3c66xRD61kIpDC10Yk3XK56EbedRS
25GpY/oTVPhIYPf+Yi9ZYtcXqOGzM1Rpf5oY3QE929FyGaKBn41UIoPszTTU7tsnFkIeu7z1TNrk
/hy84bygTU8/duLXb5OPTA/5XVMknZ/WJf7to43jnhKXZmS46ZSXOfFcPONWFsdjZi4Oihh+vvap
MvMPcZ/Ley0mJPrFnjsBOvMC/SY3/gdCGqXVZ8Blds4Uer0dnJFLpFoV/zq61fiAcrs4KVry6NZl
9Luq2alM+A2P+5l27GbtoFF5kseE9bepN9oW3Z3QF4LRnLLUnaQg5XwzGtOoC1fAdoZNFzacux43
0k/pBhIgTL/8eXUP1ao4yorBUariUEyX7mVljBSXYY183iLOEybUlaK+UY15PIgV3zMbSN57fB4D
ejQk11AJ4q38jEZewH8yFxZrlJYifqA5MYfF4ulczDuQda7dXhT1Q/8SW/UnqNDZO8tLGGPOymSD
6RjDQr5k1w7bpz/LdeuKprNjlxsPgqIeWcmwA0AdI4WclFAH0zU09MxtdnxxJt//9QTbHrSJAZ2l
OCkIhAD+CC9zHVHLymj4/nZoeSbatf35MqUwypEheoMUZcRv2TpXCXd0g6eHvOXsgYPILpKAgyP6
luIOZaoI6f84TsTpOFfPG93E8iPC6gQ7q7hanRUJsC6Airh/tSeyNQHERn3QrBZZ7/SvD3IZ7F4G
wZTKLbjHq8gEGNBBWd33XbK0I9fQC/wrANwelPAbRTBgw2e9Sr8sSeGHJxocfaXlcUjo43sl8PCk
tSAMabzZkz2CIJIHTZYsv9RO4Y2TZKd40i1ROHc2wvU3tzTCnC1Z3/m6ytqbsNPdyhE13VSnqeSa
YPXWmFs1FjCwElGblMPZajL23F8zfd9Zw2XOofyv6OGuBh8RqOVxMPTS0bM/19OnPVOioAQiKvu7
1hupcBvPIxhL7HgQF7YEAnrYVIqDgevqAgI/jPx2AlUUTGqeHDxedzQAb7O8RG7Sknm8X+3F6CTQ
W1AvWisb450faJ5Asee8VmjEHPuE29vkp1HDbkfS+65laSX7F5sUg9VRGM2rrXtieJADZX8zBS3S
tVP6whoe/SnjSw6sKzvLbTAK2LRlq1B1cFfb3f4ynkZqQKIHlTfSqTOJYPoKE3cwXaldSKbWEwhb
+d1/GgavNqcMLk6wEl0Mpo0mhxQx802jK57jEpDcdhyef1vNnchF6Imlq74O7Tv6t4UU3x6GfNJf
n3gnggJYs1ztXTVSWtx35v3LMnZVv5YVZAjG6oWE9LYXz67URT/uXdLg4XJ5OMfpT4av/CxTvoqs
5V7Dyc5eYubwVhJHUXlHt71Cxc2nEUa/2Wm2qoUeYd5/dVBAUx+BY9jR87JV96cHRn5GQcqkr5xO
mVWt7/Qg56YOKRaKbJHlpL2xdq9o4Sa1ZiYslFk8VoxBrZKdbfquT9zVRLkak1gf3wORxbM+srPx
jtmURsoEd03ZVvL732RtuJidYwdH5l7j46eYDHeizGFcSVWfZLEZGOLavTrapI0dq+PJZwApejH2
Egl+XA0w3Ufr/RUsgrlmQsl+x9rDmjsvtbCK54x9vHc7TtS8dDZ6uqk1DKx8L2sfVawTcTI23Oze
Onvu0CgFqdwSoFoa75DBVkoSsbZbp9mC7TrdFMp6uKBoK6dNYlS7I7znTXxBk8gY7wdnoSIq5ng3
lZS2R7rq+9B4HDELFSgPp08DWlUHZidxUTmD3JRAvn7rs0gikkqJoGXT22Ui17G25Q+kxk7JPacI
coAcZXTiUPt5wshsTf0kI/SKCviMdF7/I5GBCm3DbP5MiFMrtyrecA4j45pWBbhHMbcw3PajVmbU
CffqhudlFFkeIWOpZucYYOw1Y0Zmm5BOnyAShHesRWzpmVX188WfgMUbBUHRL5eY/4zzPhKQXifI
GO/ujauyycZBMq0ouJlRmcCbI4EfwfwqPYKdpn1Ulu/LdmXW/IpJtae8OjxGPlRVaddVN0fVDXqw
QJGuUkSDBTWM7mIFOAqsbnPTwdkjpRy5emGuVsOx7O6e/FmycSbTzD+E6Z8GHTMp002wUr752T0J
IJiZfOUOlXXjMpxJVobv0V473rtKBy6K6cZL0l8gZ9BuOWvICoKQFnrn4EBJL2PG2beFYD0qJ7+j
HpOFmEiKaHaS19MUCvTQBkfqGdpCblcNAQyb5vQE68ggTT81tlL4sSqkgBnBOwqY2MGvXoE2K92s
gH84mIUUfJ6KxqNkEmv0zhPy36DxrdVroAJjZkg00RwyZ6sgFwL2NdvDdKCqP0kFlI8akgcQ1nbS
PcTAXwpjzONckpsfUTqLR73V3Xup4D+Gyta+dFaJB3TViFlrIGPzUdLxORmroft1tJJwh4A3c71v
nc93tSA0Te0ZYKuNBhVpwwjvKJY/JPAluIzHcwfreULA/XtbKopkdbgknNn2tmzm7nQG3idWI5J2
L3IKPDH9ZLCE3E+ECGGRD0h8NUjl7kF6STr0cXkTAGv0UkSzooCooL7dTnx5OOC6rn776n29jATH
NEwHaGQ59KK1OqQQ6FiD7DCM+FDtcyxsNR68hS95Zr0lJCxgWpG7dakZZDlyhhl4PZcybI/r6W0I
Fi5q3icsl9PT/p92I+j7lyQlGJPiZrXEFUpT67CFNZ64dhdmrWWJpgFj31FgluLZzmcD8E/wa+gI
nDxqkgMEmhDuS+N/GDgIyshMbOjNjOBLQRikfeMzaJxnqpTAomv0RiRMkV7qsOSKhkQtzXy7Y8Sn
eB8+5FIIS76TiWzNP+lpuuD7RSXsbCdk8wFNMz4r801M4nm00kGIbl/8goPvFMGyIY21lU53ubuu
l5SigF09f7J+aAbnbLsHNFw8Uc/TTFsLXD4gOzJ4DsDGNOADVbu6fVBWWU7bFtcEMD/IuqkpCSiX
89vD1KeC+qVFlnMVESZCrw6t/nxvd4IDi5DVARxaMGeYmYx9wBLyfd81HOLoSwQnj7C85rmEjcg0
cAJzOjytAOwW8XsujkkriVTM/t5KJ9jx+waWHoSPAlt4HMnD+75w4J7wMsFDiPxz/wFJGGVngq9v
shvrrbhYM2dSsqXRI0HPYleW3MfvRVpSPBtzpWOAQv6vDvQqmCGC9mhxsE16beS31EsZ9rQU36yd
bIObnF9XpYCn2dd4IW12uSlInl4mO1RO7mQqVzr4ZXERqQv8+FYfO4pZ4aEsjo3JiMxEFR9NufXF
arSOWvibj3CJKEQZSD1NB97XOQW0B2KljmITD8KPwkQiHQSH1SYOiNE15Bn0SDuD/6tA6vMSvY93
EX4yWGHfALKE3Yjlj9MgCifV9GX7NI4zmK2Szm64Kglh+xNjFVAFBHZ4YiqmSuCmt4tjI4t/NeEx
kck/Q3esXxXzvOcaV5uhvWQ4cAMEJqdny2EK8Ta0JQdLXJs6wfv4TV3y524VFJMbOLeeic+XU4Fu
AvP7IEc57TnJgCRR5U/Jx+P4fhwFbUsztN3dUhTpRX5CuWYz7Hw2MKkYOSda/z4QqYOb5rgeSFL1
vFh1B5xrig5DENE55rKD0WwvKuP5a4SzsQ8oo9MQ1vBDzQbyE0LufCSQbaDfYkiR8KiWGgvGSyjY
aHiVHWTxtuk0o+LPCP641tLdt8q1mWChole5E5irEtueWlDOt8Xjhbyq3OgmN+tNVXYzAMkPGAYE
a9nTEDTvAZHTaCyk9119I+QDGDlh6QnYidcKgVbGWJwzj9HSn9bquufVlhkAIb895h1H7rmwQLOc
DHZydLygzRw6HVgZCyJ3aiAjbnPMKEAgaWCwRz7KUFnAZRVGCX7UcMx6Mx0q4Rnmdvfc1y/unZPs
0Ol2YUJSpemV65NXS4sAOiiU4VpO0+HJ3xQ0+CBkVFbKeF69fesz3DjGA8Z/M5oEx2YLcUNbVlJh
PrWH7PWfmN5RIpyFReJSWn+wph6snojMoqYok0YUcbrYNjlw6PdD+lPNKgm0pGKn8NPq5oiiwlJw
ea4PaLhpWZJdR8xOcy0Kjc9IZSD8320uqQMyydMKcisLjEUcLbnWqh095EsqFwPNRARBMMQUVqE0
+baY+2GuwS1762iVPfbnrBSxVMDbbS0dTn+ElPZ9uhzV1RY47kvmkYeMpEZT4crjCcXkch4H2DND
JAJ2JIPs1Gm8AvNdap+eg4PBXV/1oY1986wH3PtDwq0AL0jcWlpz82dr3OdqQcu2C3AbYSbTWVg4
rmzU+l/Cs31p8M36UBoUvQzN2vJ3FfFkinDVOTLBWELSrVzgBGcu1hjIk4QtRDG0itaEJbO1LtmF
+Hz7keZowcl471cIouuNsQJTARR5Z9bZrEb4IRD+I9c1Qb/tzroAr+IbZ9vFjsAQgpoJj3petQ12
yvmRvr/EekY1syMzR/YhjiGoFOEvt7Ws3GmCnqnKysOHUSnJ+UXJ5ic7xWd6F6Yasw0NDRLNmf6q
D4yLk0w1CAQk8m32fX1iXlW0qbuFF4BauLYf9hzw7SZWXGOTreWQvzAjJ1z/gqgn7e5bwZUbohsb
M1+A1KruakSood6S2xzZGYuWP5fZUL8mtfD9h+P6B7XY6nndeM0nl4ypuTPlhiOQbe4++GnJIX40
3xy1aqDHnI/6tTI0cV2i48roGWrnAR/oNquSFWlPchO4VK71TonfixvyqxaPDa+zKdZoQh/tsFgu
5vhRlKYv4sqoPW2fs64M4FezV/nFxjWbd1iQkcokZRzWcsnvkafqhwqVFRu/5WEtSrVamQiMbe7n
m68lop+DzUgsjy9XfvTEsS5bGXS5yNU1P6QGgiS0X4dSn9biKM96qPk//e9S6vZMAiaQoF4OIQPR
B/l3+BZqBzAljWOwnS2oXgBtGp1QNWysnOpGWjAiUqmKBJi+PuaVm+vO8VyiQXh6C5N/QUFXkYHC
d7CZ64EJP3+fGfLClvZwKBBXc9bXT5ndeMnIhMaJ3EiQBASy3p9N7pk2afHOPdw8eUL30XPqrQww
tEgNyGM76WEOJUKg0hvGjWkkHPnNKVagcDQwVswIZrT45fpJgVFvKGE+QA+OcSwijDw3+4Re9HJo
c4EiVqQtFNR3yqAOIYTmh9OzAhvbaEkYrlW93fWiYCV+XVSnCdHo43Hu5pHsmNyqUJqAhCTPEslW
XzR3+crKvzDcf/DIk3B2VicFp6nfwoPN12BxZ5DORswJrBCFHjtUUVQO1nIzL9yfwXdOTwS8tyqc
/UBCj130M7J7eFFPaVJU7OOEUfI5mBHG6xzRMjZ9kq2dYGrs09L70nJLTkkpneWQTZHMfYTrhsg4
HJvJTN/1NpQPvit0s4IXaSEwCyvPJ9+Xdu58mid6pN7XPZAfJW1MKsGPOH1MbTqG4hhTC8WJVbjn
PT3OWitFaD+i/wriTxqYLPU6aItRgi05VwKbNhHA+FrA48W+HrsQHEXYiaFlSeQpdr2qK5gtHSxK
E7GembkwkoSz9ZAq0r1XHEtpk6ifhuVqeX9KS8g48nhGvKg6f22HfX4Qbe8VmFEwnuD0EFxUWhGp
tJ5KFLzeMM7nu2rbke0/a8dYHoJSaiWCZ9rnKzIDcfEAljZ8QR2TBp+6RBUYROrw7le6cbKkjBgd
ccpzXQ1UPwQwBS/1ZB4YJrffScDDDCmTII8i7Y2Z4t9bWOzzqb0LBO5T5v/GhdQYewe8mXHE4Cvk
awXJTzVgMG3nT+PdqrEPCrSDdHalIYI3TA3nUrDkD/YG/pkhH4+a1eoBemq+HS7iVhoT28ZXVWg0
i3460fxOnXmmKOgwWfsn0329wgqakelgVxefg7541vT7s4+odntTjJgABVs6qvU7/105OGVdEJZ6
IIffao3xfUe+TRjxFnI/GwV7iD2EQvRFkSBSBufhSHguaoHAZbZi7Bnt3qU5vAaFr/UiOsMTJiQn
n+uHgw+YQVvukFZrXaDN5rSHN3IFoKklUnNB405gpZMF7Whj5iRyKr/f2ibhwk0zLRBM/TBurNlK
3XMndriIZOyfVFU1ueEPFIp4D25I5buCKdJ3OIZ/xGjp0D7FcE3jjPyNvqcTe3tQ1GN+aUdwrZhO
CtgbwdmUCPl19za7ZVo767Rui7fxazTzKtmdvYi0Zz3Tr4klEd9PgbkQQWlk3bbpLKtROL8cBpCW
zgxpT+TSsmO05HzbZyMYQ0ZJau4K2UwIaadZca4aXFlZBE+fB9rNSsfKP+rjfJyHFfKAKwd1jPK/
WK+v7lk8Gi9UWWMOOk0UktZqRNEqjtN5moABOKJbvLeFVRkkBguYdIH2wXQgpUm9HTvncCk9iWrs
jidxiY9n7GyOOsS4wFQRNCVySzlIuJVKqMJTezOPxI2SFiGsLntKLBtL/lGwjPkJdTWZ0ZmyIAA8
Oblrn8ZBjPpEzAutgHck7RoebncBwvMak1gpDIqejWpk49eCE2vgmwsUh7xP2YggfXMfcLLxs++7
GHka1lotWR+vi8+P3RP76M6nrcmAJx7055FW9xY8xGIIIOhMYkvF6bRZQNuWQ1kK2emXET7+mFST
ih1gZk3euCEevuM4WJ6voqzHJzkZICcHCbpu0PxmblWnzpilzhol5ZUwOxQO8JyYk3Du2huiKX8Z
WxtgpV2iY8z2XlywUT2jKd1UlTZA0zh7DHKL99RwBvuHkzrxdlgst2FSiaabjWahFEHPjJ5PWF0n
ab7w8Ht1hNYR4MZplJqpUiGqAcy78X8a/gF6qLI4WgWYRTypipaumehdUxYKT45rJfjILEhKVgne
pnvuKo8AzOAIkIc/dLtyYLZPLtVoPiF3On4iR34JFLI+sremgb0X8WqUg1GRxtSwd1wk/SQxtca6
ke5zf6tbf15JJuOK8vvXPSW+f4Vx4yHCdlONE/qElp/EXkcJz7Kd7xKSAq6cFNdHDK6Xk1W4NvMY
yGSdiBpax3EDbOZaaL3SQrEstiQLqwYWq0D3gjT4AHnuFFxHpdJSnY11WcdKcVAv/bsnU/eWkOD7
w3k4YeKvEuCoC/dR5FrZsMWcIEzjmcNZvEzanYS52pahicL1EasRF+azcpvf0HImcE+MLPPJ66fe
H2Ybvl/c9Ntxm/W8VbdXrDptpKfedSaXKhjTEmdZInHjQX/8QdT7NpAbtOtP1yh6+R8K1htvq6Kq
SZCszEV51LYHXMopyLuMz43CY8DAfV6lIVKZJbeZhjkHH8Qy4Pi9c6xvmAJmd6Rk+ItrCq+OIuFh
92UmxsOt52fwbVOimPXdFtfOwlGOGxO7X18nv8Mboh3/kyUUiKM6/W6QJCcP1TqQvNtdled1WH2l
iHQZN7lGU4mJFvUNpVDd+MOH+16W7r0FHGFQkfcH5/71ItCg4tBlBVuwyRTCO+nuYo+4QbO1JFa3
frffv5Jh873oHLMx2yCQGDn1A4dX+rivOpRMw4/txyRlz8fS/hwDWXLqEMpi74EgRCflR8EJjR4+
z9dEjPm2Uf2oUlpmq06iOgY7MNXhFm5BLJ7kBscAjekJ9HXPdWUrMVmMbdv+KSko/yBVZ8to/7Ig
BnqFMdOMLSEJzLzHWBxdvWyGtQZHxE3x7Ar1ndUZCc6IPYOZcMpnFxcVEs0+z/p53SXAVhQiKhVq
Ru0F6UgNunXZGplvNn6Wu0oOZXfuCfjRvjWcGz+L97HUt2GAYmuGdSBqPt3OhUuRK4O0GNUwFe/F
6HTK5sOYhvQqYeTIJvYneX7O4HlHzG2SdVyO8OA44sqvwuxlcPJGVzwH88FthedZDL+sfp1+pRkY
OXCu8VGKhJYSJMz29R+Hwa7knldEJz1R8Aua8pscsEumiYB2NAo5PHXPOioNEbzx6PJYEfksnUPN
4tFYD8Uq9gFBHqCWgxSjFiSAJwUdYdisjscSULMsFcF8EW7xy47oUFIy3oJ6MBUmgkoc2Wzitq9w
Kc40+nZ81PZgaAaOtEDkD213xsWvrjW8k+9wu2qTzXUFZHsQIZ2XeWH1gY6OfKgU5InRYU+Tlmc4
sjHA+vGwv64RwHCwvwigyOl4iV0VrKlcuXRj/KjU91QS0EvoLzt3LiwLpB0Nv1yDd3O+LbSBI4pt
ahXRiHzrsjcx0+iQvLgJIKRJQEAWYyHxxgfyMPXs/s+hrEb8VgjGXyVYMF1fZxUCWBycfdqvluE0
7vxGerzvKjJXG6nzl/MyZ2hAcsMaVzgwi6bygrtFv2zycSVDeRnfY8VUDVqirodL7JO61XG+nNN3
7XdFTDx+r+JrQLscR1/v2Dj7JhSdfWcz5VjuGDTHLPz3kYMdT+0kDY8TQAIezXTtLrYqhVfwnxnX
JaLsvZk6DgiU9FzHU/+IMNZMlueOWrLPt1EnOAiuGlasuZjgoOz+As+iuEGiojuCvR85cbbuZpxm
2EepG3VytDXKbG8KFdDtUUWCHdCISqmDVy3E8cS6Fng6lM/4xWYSUtpttGK6FR0FACXmeOgDHNvU
m5A2f1Bcj0b2h5aCbiYRzPgFnLhVQk7KxTQnBE54hMOBDWfcrMQZJcGB8foaxg0yvmJfA0l7TSFA
H549f9F+8zXdEHL2og5g+P8I8d2JTF2whWcQ8FD7VlU092ntL+teaJ9Ap+5nXtKXWn1D8vAYcwwF
Uy7Wl5wsC4JT6QAwu+KYQUALslmK2c9byXSKTKv7ZVoouxzU2TAO6yry94EdcdueFzkLbVAZxgfx
XBnh1eUyBcVUZBZOWoaV2EZWJUOijfh3Erb8Fg/e+sXAUwCKl+HyqAtXlosEnkAkoHTFYuEi7ai6
q+iHn0WpcyyFweqF9C7EXrSWu5rAObVAZMUwq+JPuzrTPxqsi74Z3VdpF7eB2WIQGsfCZdPi5B2C
djwFSDZpvBzMqfC1c7AUOq4bbIczIWeop1BYUOOQgX02HXrx3hdpAs88x2UJwibre/wKJ66yvlL4
tcQ975PKSBtiL1tlBW7kofYCfpFaoAiYTuxR1BsMUHUeTFOaCQHM6nTx8ZLPPzKhMWCGSGCBM+1c
qoNxZkWZQNIHhLSIpBh6dzsyXm7x5Wp5T3LRJZaUYz0u2S7RigpUUoPgSBQJxCIeECOvAklb8+yO
UzadDPlI3R/W0GzxcUxAvW5etBDjvzFflb6OUeiOJP/IIZCoJUlbFMiekz8R16yIgwsebcBBILcP
GAg3tnzsrPxee138VX9LhTDAw10b5GIJymOr9bMPNQ8RxMLx8MpgIKvcVfrR5E1ODGkd+mZveupt
9Ml/wMK7P4d5gt5C891CsuYND7KUnMbx7KIuJ15zVFqsi5Nab8Om4jvtlQ2Ta/50r1H9KFKUg60e
kRYCHOLISZdN2JwI/Pyt7JoxSmcI0SypOak3gyTXezCp5oazEytv5SXOFA3Xblq9L22F+KkQEvPx
1Bt1Nl3Z/rQ/JoTG8tW+eZYy5P67AlBntikFj2dLAm4h4EK/vZ8AaOiUBhE6EGYpkSvv7mfpilIe
m8zXAW1XTLonaxHqbcApACqpqcVKIgxPbkFh5QQlgMoZdf3r8bbhNsqbzFLUZyQE9hHCMamtTTQG
PkgvVTlfavA8fJqYVitjvOuz/F/UCKCNBwOfZFQtOuYPSyM/NPgRjZFH7HqNk7fKMpeCWkblkT3t
gw9c+uk+uLsvhU3yAk3vg/F6pC+LiK+4V9rTru3nSQV94uliCbtuIb0m678GkpGsibIzzU2V+Sm+
TcsMeqDSQvoDEMsXZWleOJpDKgGW3NBWoY65gdf4X4E2ppopv4cLsq242fBE5WG0+P45ign4q15i
WbIqN8ZF+R+t9CA5vO86ryFEJYnpjNQZTh34RI8ZvmkR/abGn6/jw7m1IaJ7iNXnAiXjr2MdgYhU
WT9t+5ppGXCbI+W79L2oa8cttp5Tt1FsT/AIuOrRfn1hiffqIX7y1ONWTKhiBqs2n5040Y/+DsOH
FEx7Jh4tB3jPh35jwb0VOm99eYAYCTFSgb0eYndeHjWHDQkVcIy584E8L0QYCdU5w6hHHTHqL6gj
UP59XVM5uSXP/faAkot/q8J0jPmMftypuH/vJLw7OpndxddmQsq43Mxnz/tLpaBKLdaJk+1CGXLG
kIaxM0pDp6E3At1VsxfwiqzuReywwNhEwRGQkgnQjIuGhbeYJq138syI1zzAuiNyT9dtpn5WtR5N
tm/QQ1rOAEpsXQgHZOT+qVS3whoHH0xDHRGgTkh06FxDPdMjX6P6Jzxo5kq7QEfE/Hf2zOCFzG+7
p4oAaDdAo4AnN1WRILWa5zlWky3U+s01z8+Uqk/zIFT+YlBSC00HOHPm/wGiOvPygnQAEGQyqUbQ
7t4LlkgI2XhobzNl1DvtIHmDQlLrAzo+nNcsiIJCeyH5InN3+rl641ylFZaA6dQXaUwIO7hK+sTE
2o+WM6nuTgFIaHgsNSPmu1mN8REOmZyqbWlfiga6WCv6TRPX3iQ0Tgy7dTSWkv8nUfsjH1KcuU3q
4YjVPOYxg9uc/z3N2IH9Jy/RHS24VY66YfcRhw+WXNoyxFxfF2K/NtPRJsbuZYYO5URjz3oWb0gP
ELIlIThgj6ciqyCoubpLfXNmGP7iHfEZqXIBMZ6C6kryDn0Qum7AOvpMCRtKkckRZYpXknnDuok1
eIRbbh42/BVR1OrQ9Uj4L3sk6YYou6SsPVvOYinfiQeHpvrmWNqZSB5YuYoxHtxM1cLkwb5IWTnR
dMxhIqIDtdyFeypq4T98ku/BmeBeO8oCndTy/hIKVwAgh7ZvNal0XdnQULEm5i7nZW0cgZ7+6jBO
61ZR0GEU4gy5C1sxMjvy2tYVtJXEYrDLc/FrM4wBVpzja3LluGDVbPyuYzJMppLSjQDJtBB53VS+
+zzZglf52gNW5npIodKE8p/razGc7XpuQgh8YMppjXKXgJjMMSCxGSMHUM1CpzXth8gwd+6TmFZF
EhfKZ+RXCO+QqsZkdUw1hu3fbxCiAAvWUaRNft0oOJYoep3uoEQe9vvORqRNd9BEwOolFcw04ISp
v4AvZy/YIkS8XR+z0FkOec1uLrilx0n1HB3wun7C53R4PvGoOVqAsLnOy6rwiiuuYVBxf6meid6F
bvUl7EsIVxOA/pm2AfRM9jMbIWDby+yX00WvqI2Kh3lZ9P9om8+uZolJnj6CySMfj9NBUbNSX+wZ
7K/m8tc/s8N1N1sQYA2aFzu19fY8WPqb51ms3cLutIjB4htyTOKxZeD+dBOwD7EAkJotsVhlz1JG
gt7JEfXYvAE8LviOTvH7Cuzn/189CtradD+4FeRBpK3v8pEuiCiRvxXsnL766enrZr2foZ6FAZ7F
OU5cYx7C4M9viUBpfEk4moEKNSDXz6BGZvd9dt0ZO9JsBok71gwcANzGGdFPUbbNxTdzSrvIb4lD
nhw4rGMeiHBaBNEPb7qHYL/xtyK9c14EhBvZmPNmSZ9PZb4YmHucJ/MOfEfAM/F+qkKkme3nWx4R
eZ6uGUcagLEdWL3N81OKK3TbDFowgiSkqMc8Sf/mxm/TvC68mKPI14kVFjvvhp1sThQ+Y3A+2fqG
mgAcWrYmoK7NvrD3aecG3t8Y4XSIt+eaBQoXxTeCgetLzngKJ6cL9Aexfe9mQgjTU79OedjzQFmP
WFeCqezP7/XVI297ed8I8wfDFlNu0a3WrmKVlNAeT+R+ppV4xrotSYfLOkZZX8aN1c1jCx2fDFno
tnl9TNPsgGDfjWcr+1i6J4wrOw+ha6MG1VNyYl4KJ7jAEubJ1ShcbYu8czcjc7qpx3w4LjR7w+Mu
0UgD2kZAK+86WZeJwMg6Gv5G7ruHwoC10GkFdnEaTb6z6sAUNp5Ye/1wxv8+LKPueJroOiAhcsQC
sg765+QbhJzCBee/6SpJQ+HgkzZj0fRjFKtjJW7bhmilsWJvbm/siD3BI7Gj2NbDRP1X46SPf0Ui
rtTUHZDCnxEss60208gAjY4Fl4lWOYE/hu9SphL0b4evvWm54H4/KoeIpX7kD/TkyfbllAY197H8
la+qzFyYctxUn+0Oa4vU8P1aumzobeCwJ66M+wfWZPDi0cca6kR0YE9LvMxFKLfh4+Lkk//D7iBa
NNQLo/pbZBv//SxhHOAGJPRotPimfqdVKu1fVQg3Xwx2WiokPsKz5r/LLq/o47sQHiDUBbOgwF1v
7y6Sk7/SWxv78L72JDvmqQYegiYzgQYN+Iq/ZgPfcnUryKTeLnNyXwnEdTWzKK0ejCiiEIh6dy0k
Dasrw37mt2w+ogVTGMQcTMGIAAyNAajx+yxkrwTfKNCPRAgcoQdYQwXqmAt3GvrY4lia26Yl5Mau
bTVjHk2vXqpVcTpl/ta7d3NjRmEr+bQyD9JmGQ7ttpMzqVsUdkfyLxZ1zql6gMWSXUHg6Rcwzc9j
G+NiUsVHhNMT0fMB9kykpOS4Xv/0gV77UZnjOSihAqZY5HfQS9gtm0KEhN98KpV7CS6rBaPjoN2w
UjNqU2YeBY2E5h79ZO9WeWtojBBxMR07+GxjRlqsR6s/xE1U44abTfG1l2wgJ6xftfwsLYbidilk
HuSsiH57Q/BkTj5LwXBVVygNVNXJiyazISzT4H4zC+4C5d11Nx7uXmtsLiyp7XE7dg2XZ9j+OT6R
Lf273FNlg5mnkachC2b6r1ciopuyOsyBV21rGMu1rvZMsDeQ13FgNQR6v99hY7LYMkXAp6bTaPMW
c2AuZNaAhst7XeHK/aPojpXiuVqhH8qwexlZANgyWxX1tHrYvMzaCwyoJ/Fvb6M8Fv0h4AQU5cjk
DQVfzNYV95XzpQqTauueNZ9yQjnvis8lROfFKreIX97kHvXbr/yyWQftkbksglKU/8TOk2y6mxlE
Pq3IrlQj4aW0ekcHfS/AlywcwTZ5udmnV9ZZLfzV7GDzoZAOU4HGIKnQZGkGXfPgL+yGQer5SOqJ
tCBUa5eM0i1KuFMxOh7mA5XFD/KFi3gjK2bQNo42BSrGuFBPYstAWNTTbzcZ8UrXI9bH4v5hCxQz
PlRy2dMmKwslLEAoeAjphGwEDf26grPrRQoaBjcPLlaK6TEDfNF0g9lhRh8xJSJoVT9oe8LX9e4E
bXcevDPvztUhDYLhSrRIOyjNxqACG28CpbrD9NtS4kyy+wDxD2zukQ5zeMBXzLM6apwIsqiFlp7z
VY2UdsBM5GV7BzC8MEs+cWxoEDC3Y1ZacL26kdGLzyTA0pFUU3pBjPs350G2dZj7K5U6V7gAgI17
1zNOYci2G3EFa2SPJMjGfmOZ9Qy+/5fzJyqeeI8yafA6JSydRU/ONBef9KJWfd3WFb2Kdm3bIQev
C4nLvxbRm7PQxLsDnRzJWN+tHAXBguBzyh6/T0nKHxX5OGyM4Y1eOiIcOFJqapta+Y5o7GBcvQkw
G9R5nLfMoGcR8PB+twFNS6wco2JKIgegVuy4dzw8Rwtlb1XrUoMR32MBxB0cjD/z17RRi4CyKrqt
50HeBDcxqFM87yExQsLroEuQvSQbEa7SvF0LmIPbHf8d2nY9c9FHmGHq99hCoBbwFCCnln3cBHz0
9SaqNLFsVp3mRc8DykalXzxP4uTQhJvc/ejZZZIUnFb5Ma0Aj729I8MrWG0D3e5qngUoNQ61nBep
urrfmntl/oRaSKx/giHQNq9fQRapUNCPpVAaDwUZzAEKuGIcNQS4XzStPDyxcQVT3AHenCwG0fSC
R31MSmbWvytw2xOBqcPADxlm8NrwsRZCvJ2v9zzK51W+P5S+2Eew2WFSBq6LX31phLhfTHCsh1HH
/g2SWOf7o6fl5AwrViFcYzXjbraIolvZa85o0Q8vY6Q3r6O4nviv4K5RUEUvgcSkRSxQerg6pMrA
2nnHwOWhpE/yv5vJtGfpgUUgnzGSXLRupeI4TOIEWxuNQJFNvD2NRDZ6493OnyW0i/aXq/DoHbIz
/121J6KK6ZCvsbed1PEhPP/XU0Ip9DMGf594pIii2n8oqRGn9FSRpslvBQ9Jkg==
`pragma protect end_protected
