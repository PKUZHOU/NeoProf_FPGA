// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
PbMeMGmc+GPj8+Ny8hyn8EWbKzfnQHZ6I9hg3vULAV5GFqcQx1q6+xkcfm+U
wZVU0TP9PAyjvnlo2dfcXd55Gc0lijf+vjKDOtDIbHMshnhIutkSJmg3bgCE
0oMNxjTdWtGZ41tHSach8vY5BCQ3FmM4ArmmIaQrqLTP6oNP63/VaNi/Dhi5
6hvlODaJWZMq2QBzLpfbFN1PuCKyQZQVT1YnA8KocMzphdYvx65lL0iltsNX
kajFfQHk99TSC5z3jUCODLoSIj0K6IxXP3ZNJZSQuxfEVH43rfY/wgbwI46c
HciFH6NEsORaWxDOw910Z+7VJqoWaCPrF3nKgQoR/Q==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
jz4lRi8/NuPxP0bATDBtT4g0YiD5w0CM26wnVp810hETNU1RbDnWAFzU9MJx
s/A2lEThx1AeGu+aYzMcQogNGb1oetYEL+iOAnZdk4KxmMkQyaARXEljinu4
db1rpSAhw3UXsEybeymK3waHeSezkskvc/mahRO6XPP2w+tNu9b0YoFSW2QG
fGH+63VQ1fDQ6ukm+9QAa2PO2ivKXtwHDad/rl5RLMXGpYhUUZ5iB2uhL2XS
56B/v8p9ZbnKaZso1pMzGVOjyZMk3NvLDz7gd4XwYCzFA6hwf64drW42aWRe
9wq4OEOJxAhfwU1zbGMQZzHO2NO5BxNPHAyaUyjkbA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Jhc4j7/0SAmrV62fcV+0aZgxaomYPFIrE70kZYLzs8Mt5r/bmXs+z6+UsHvy
bO6Vi1u72u3fzOafoiwHhj5xgpGyYhOyIyiaKyQGIwayw4FlGLuN/MoDIayE
YgZmsaqezRs0AlwMWxlQQjmeeYWTGFcx2LHm3KFVoDdhjnn3DUWXm1X0FVsE
QILLa563PB8gsYVL4mgMRN6tbib6b5DD/4a3RgvYuKS4tvQJ98TYYfUN5A/0
hoNMPstR7qthHlvBFWstnK5t5gLYFp+o/T9f9IcdcK+55PwaUQ3smlnqI3MQ
T+VUtOIrchp6pCGDKoOBilJTc0q8HLuCodmu7g9pgQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Ke9bkAuPdIijvAHOXaaCwCy9TjFgQ11lcrob1Oo4pBh+MGz+wSYXZrEPrzlF
6VD8Xy9zdFKVcS0+qolVqqIM5mqIIwN7zssDN0ARO9H8mYY2zDx1CdSh0Hs7
pCFaYaTigsuj8NRrsEr3Od4+N4N7XT0+vwIEbqRN0RRcgNuNKck=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
d6eGmb2NhLcE3HiVUC43r4rhJKIQcDzR32+zSUsOOENENgxWsKOZDhNwBiTS
NLnK3lHfoRkWdQ0dV3PR2kfslwXcvtUuTHbOYb7WqJeLgjNSXT/MPWoKmxpY
/i5/F5Hp9a4x785jk5MKw61st7bJN02F2DF17fDyMCkRsU2X+JosfiJ0lQiq
7EswKpvHFdox0AQunGYOtfT0Q/MaoBokTvVAKizFZkkGwtjet5QCXGmtSYoG
Edi0cXHl43M7Kxy/GHPBYbiPNjMMZNibQFrp+QPm/Lx6tN8CgRWs3jSn1jdY
r3EB8EGlHCv2uw8GrGMkkHy1L+THReJOzzwLZXONeDFeERV56kaAqTniqOHA
K29LGzH00AS14DURtlyvEKpXlAnKiAnY3usNms2dr+eJuigHZbwgm3t8KYvC
OcLfOIDq7UuC/6vL6bmidjDtxEEcSDNSMypGSDUvn9W9j8948F3GWoOjc/p4
VPaFqAig92NrUSdJZXvMqEK8rkGl7z6L


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
EC0PjBw/xBKMRwKkYXblouxQNxsLplV+8WpRBU/NUhcaZCgpKwknydxPMan/
/WxwSvTkBMxcdFK6kNHbVl+3stcS68dZBNPXGc9aXTx5uHCSl3rL4ivGsie5
drtXm2JN/CigDiHc0VdJwrnjb1xA72wANKCzwBdxSbNy+vFafwA=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
od+2d+KUTZYCrKMjhgjAUeUaNVf+8kq50T3BEQTdQnBmMUrnpHy6Lh5Z0eoH
vkd1ar0YSeeQfOHm/kV8YuU7syVpWds8q7I0zcpCl2Tvbf1SaGixlm2LOxjU
UnIP6pvFZaHXwjP5UY1FRgdtzGyx2xjs6/Tfvc74bI+NPVb9nKE=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8192)
`pragma protect data_block
xczv1elPFOTA0iFkeWCnKB/c1MqqMHmLbdknW48d/1r4sKvfeH5HCvwBbaLD
OPNKnCfd6GrmHJCOtQhT31RjVmdJqUkL+sJdgqLfap6pFRPTy7g6ax0vzNvi
jptJEoF5dsNtDBL3nZtk9Y6q8KlZmkd2fI2Ljaot7N+5UQAMcXr9RLwd6Izy
Tmd5g10UEF8R0gsJ7yQna71vEtxenQdtOQ5oFdzXSl5QrpNS8tRIs0T6Qymr
EENC4zlDmbl6K9ocN3EaWYfsQQpwpSuO9UdZB/aQbgHTcyTR1LbYHyCauDXu
dq5B/6qf/Na1go4axpxanIRNZ2sSVb+k1kzHiOXgj/AZR1OUJwo0iXfD48ha
PZoPhKtT1qmnmOACLYC/O0INUURGp8d3TL95ZSFr34xx7fEw6E3fs506H0sl
IDhwrBcewZVieuADYeV1KbQ9LaUZkK6HLt+tlpm8shz9Xar+d2yod1TsKlNc
TZzm9qmTL2MM04LmkeNM8qvYrJ5MrJad0dZ/FcFxn3FFpnBk1NMjPrmuFHCY
E51iDkwar3ys1SdTnhUG8TQwG7Kzks+ApUVkjG+RDSEfiUft4uNlP30FvTrH
FSIuGA60g0JDXisvXzJuea/ud5PH2LNeygQbN+vCS/myC3TJRD9zgD3mkUmg
+n39Mdo2yq7uiVLB6R/eyrfpPoCtsf8+eSZSB6mU5K9zTy51fMJnv9af3wwV
11nFyV8oCStaK9RDJHjoX9uJbk2arDPMQ/Zn16NTv8OkzdAjaBqZdam65MC2
cNVFV6RSmv0w1XJAxAkwHGR2P5LlxFPfSQG2qGpJX4/cTSwewUL9qJCPXn6M
a9iouLzVFq0hO5dC24EXCPklRilg84WDNBizHxG4Trimtbb8RtR4pfNyD+xv
StABaqULxT8BZ+O0BVDQLh13op8WMK94jdPhy7uigkdWbyBBcitWI32umQJo
24UAk4kVZTUrcIB3i3UzflljMzdrCFLjcyDiWDt1MfUtuAXza6sy2qnYKsya
ipoSeUa0xFzSL58Ufe05H/PDWJw1H1RYGkVdn4zLji7CBN1ei6M65TFut4sM
vmf2S0gKclSzA61xTci+g4KJrlV6MG/nGbn+CPbGjg7pQkMbMy6hTN2M0zl2
F4SGghFbPrq9ZQgg6TsFd3ytQvLb5M2tzakGUQXWKPDLhG1ZtCX/M6SQEWTm
KDknoY5HiHSfCLYPu+A91nB9U/4IvD3/ct8CQGcEHuGwfGALZTS/s5FcN02R
Texxr5Y6qYGdU8LslrlP9oKc+bfGriClfY72/zVDPUA/P6yrMSbbZijXl8cm
BkNtV0VUPMn2XBwyQ38ahcc2mcRPDocH2SjXu0rxjHGaZdq/jTsIhb+9oXmu
5s6FGsfws5qEQIPK5wq1Qhqybj60c0Ap9IcFuRDG6CgeYCW/lQPBVFVHkb/9
TxXg0Z7K3gqDA8aBCLQoIFDK1Th4aQ1n4rVizQ0o1Y9D2pCpMujW/B55cVTk
8lMD87ceMFJa+OprLMfFihlxvgxx88XJlRD3sJTSD/GGiheU02JgEmQ5f1Vk
hRbPM+Q5m1qzx5G7QrCVszXCEu0kllNK391SryesrEXdvEjSVokUq6qX6VA1
ZTo+3r7iHx3Xn+S1kgGJ1b3IFN7X7xHVd3TFHY3V1/q6GHTqwRz0VaMgEJkn
zcjnnI/604bJAwUxPsJPDW54uJ3JA9Omld2lzaha0sOOBpFMm8C5i1vZWuaf
MNzYAygi6+CJD8MWPwoeRxr/LNxNMsS/JSCU1swz1DFxLIaKu0gbFWFoqdjz
XC94UpSZz4FQz6sCcaoGGFQRFwiSZFD8AMZUXduq9fLg3lNYwq8bIKzZTwhr
sRp03d8pam+AJ/JIc9YWjqjWCn7C4evSZPKx4jlBMrLKcpYcIP+JmlnByLQd
DusoFcljkD6Y3dGLJW11YII7wXTXmXHcLBby2upvjk8rKDghAteGW2xFiHmB
SgmuT9Z6kD7Jga9nKi0o2b+y83havjhKH+Yb3CUD/BnyrfVYKoBTKOLuhzdz
6pzcM9HGC+z62sQfnHmaPc31Zb1ZkXglgTU6erF40g0L0vXu2T6u32KU/wg0
8CW8oXTkVLUIUGMXYXsFxiDbFLpBKJV9/gKe7wJ84trCpkjSpsuEqr6aIM5x
lTjf9yfZkZ5JSB0rZHmj1cZJvegIXlh7GAZGoHZUzlOeSX+p8GzUd18o5kXS
IgQxnsscmkGjt63L7GqPfLx1qWnTBggn6hp/WQ9PRnhGaTBsDdcCOZ+iuVX7
NtZRTxsSRPgqUozX7Ax07QbHAYg4OseixbzOULnuIO+dmawD1+3u1LvHllc0
TYdP9GV486qYp/EZQmzuXj5ziOQDWVvz2cXjd3dUhAaOy+n/cG38RWtpvXK0
xOyZnCv8OZgbNSGhihf8H4Ya/RjHs8jUwucPJ/dH7OhlYTBai+RgqjvKzSn3
cdZid1tNVJz1aOX9w29WCJ5jfzAs2W+t845kdFpEGX9oq3blJhv6mbJ3mWc4
ZEBJ1BUug6imTt1zgfES+LCcQH5wBA9Y/62wdKK8TJFLfuu0nMm9gF6Sw5jZ
8U9dwtLJ7ptcnV+RvCGrtqw1f18nKqPy9ByLWehwZrlW1Z/kZvHI0eADSGnj
TGrAN+8arAPFMcOn0sQylZ7zjSht/aqw1ZD48obtdEt6heQmNicMxRuJCqMc
N9HLTj9mnQZRR7s+onSGa0VUZNadsNfH/KM59NCkihE2xjo0tEsH8EdSzA/N
igh8A311IiJd/Ih5YR/F24DO9GSmbI6KdgBvjrKmkl47lVF4i8OQMmVOmrT1
74fKdGdwIR0/vNBfR9+zA8tmNihLT/DXCAw8K6jjrBTOZf1XdscnME5VuV3b
vMk8/aBVWgRPmRrpDBLTUUGW3RAVoeVY8SQTj78La+AxZVPTTEJ32peYKkZD
My87dzZbST2co2vKqG4e+AedX/GbxCINP9837/Jo8LzXo0C3vDeJnwD0dLPS
zFMVqOWj90azmx54prFeZ5F6ca12zw0crGZhdcppDbgfGTx0YU2bk6KcWXTn
XdCXE8+sJS8gpEGh10kRLVr7Ab+K/RLxReGFSK5UnnrL86CbS2Mrfgp80SCc
k2VMzr11niPUtvdb1czDu+jxkWiRXy8FFfpc1t2g4BVStUTQmaR/GjhmuH9T
kqK4/6V05vsyKfP/JIkHETN5M+m7cqiYaxt8rPg06ra74dpJW6kxWGvP7Q6B
8DH0TjoOkzD3TTmq1tZEX9A3X4ZLZFYq1L1RAujMg7dhAOymLhAIK8ad1ZyY
inKvEq3M/w7rv5vaduNxKZh4bNxBdfNc2/koyDPzMHBY75ogSD/7e2SrQHm4
zLGpWDy42uPgGsbEfXgA2FSIAj0XFOVQjyLjEtqNC0Rta4V7sFpKSvNvCiZg
Uf81G+xRfvKAF7pIXF12XYGiU7fvk0qwuuK4KopOijq0HTyWFbgj4YFBHCsd
ubVa6c+IjtWrQzUeHvcVhjSoFRzlrE8a3hbmA6w8LcCj+uh4OLEy6yOk3z5L
JyyqDmX1Xat11K0NzQC2wbXG3IylnSctV//jRs7P71YEPGn/KMWbIcOsZcjL
/ujffGfGXNkb8WFA00kOA0n1ehFzqebdsPJDEBbcIZHXf08l/CC5s6OBytlM
PLcLoakrPC0XWcv5m0Kms2l6kNLZ3k/E7zRTYids4hPBiDdWCtXxIsGhOZfv
oJda3vZHU9s874tCI6rB7Uo3OUFLOxnH/b0NeOJu/v1pr4uPphgddAOPGaMk
A9apKj/356ND7pbiLRYLKTqYBsQHdpOt6H5Sc/P+Plawxw4smgEgAUvlz+ax
0J0bh9SpcF2Kf6HpjGXpMqoH1Wk+BIkGWBJl3J+Xxr4XBNWrDk5uSfREL6vr
TLzfCNY9zFhYHO9TodYxTd1bZXB2JLD7x29oo/ALq2OabbRgwukZIiHgWeNy
P4QMhd4unbijjVzyfYOOhPAaOhFvnsxqOqL9ojsi3HQeZNvZ2qXXlBiaOC5X
vDUJo/zbIbRPmfabuTDC8AC5Yd1tEGW5/PpZYtL+eom7YN+1ZnY0H+pbYcWJ
wVHX9n5in1tBZtGogpWVQzeRSXEtlO39cAL813sB+IYe9+zVHbd13RDZuPeG
otNv7IscXHMvWu5hiYkaRCMbVjjP+qRt/do8RFS+omdYmLplJ96s4wmPMYwx
9HacvuL93ebaFRmqeuXDzGpH6WsRJQVrQhcTsBNT84YABxMUtKKalVs3HOAd
QEL9eCcPaVEOUCYNOm7N/hxpBQXa7qR0Sv8H13fOEUWvzEP8asmRrWf/82HZ
TpN2iSi9oqCW41lPmHPv7dCXGgtWQAxtXnga9e1zSQNv+VMRYf6yMIMwj4K5
f9ahNjb8WHtCpC91DIwCakDA8eGmHG4TIbGqbNzpvcDh596qCPCkxixgy10+
D34TX1MErhNROHE8DACpkFi2yaXAsoA0Khb/n/6BgB4PcBSw9QwFp1jVSw7w
XXfy62nsrJA7IUnK8t2WupqUirhvFqZFoD7v4bLENpusl+IPLZ0+AqPdQ+0j
OR/MaGb/CdIo8SH9qwGOL88/PYqadnhfG0tO+EQ+pNwfCdMl/cnY8ZT/lWGj
gPED/ZfnUgVLiYIjuxRRoW7i+thjhnQxhcuTsWS2ICc6hBayGYiak+qmywY9
tzp8WjJGF599jPyplkcZavbSABmXdNV1YYzmysS11rm/BhFwI5jKjXo7qJ6O
TgTK2CRAfsUJPMsod6TxBb3Q5weqMXoDLxSKGUAmH57Sxu2cIlKAFUf7xwjk
sUVarlZQfNWCQyK/3fj0M0eZryBPOTp+PABhHpluBPcBcCVl1n2A17NR9GhF
rdiz4O0PPQfGr8yr8DumarNbiVkNQfq08TT1hnc1Y5FV2AxLSILp2yqxlvQY
BcQxxpYxQPzb9TgkYbj9ZRnXFvhOqOKVU7J6L3xhBt5RqRIf/i1uFt+SfJVr
hmvelOLY5EwpDAXH44y+N/i+gNBijR8k3bqi9VWIOEjBe0ykE6oGuAOUt3Yr
PCjBnxPkbZHHR0GAz/t6Re4pFA1iGTD7BYC3VbnZTZw7Mt53IpiWhAtkTMMX
m7kl2iUPlhvONNorCLw8m278VDxVHLNbFpt4orMoZIKR9IDcDSIH3+Y83rGl
htAPe1fX3pwAsK1N6FFdM3vmpz0bRgrxtnlIgq+S9fopImCW+ut6URmGANXZ
iZ7g+OlMF2LUm6Om63gRE1UoP27SYkZqmAI+PSlrP4ZujaI8DayWPGL8tU60
nqOkJehkDVjDz3wAevEx0EQB5XRffMsQHlof0ujfE2C7wi/KH86lZRt/83WX
243gwt87JYLuGkVrWVTmwcYGO+HArpOndWvJOMcRwrnA82pJoaW50+9q9y36
eS15agpS5/zRBCaH3rN/YpzyS66cqrGa/Ii3QfNfL19FDqfpQAz4SD58E2qA
TDfMA8XqApRckH6+G99fqiipojvka95v7SUpCwnzIRnTVP9kdDo0pgtb8e8g
vTWHuwa/wcU4UShKgljPsr25Tg3F2zIjFOWyNu9QvIGURz8fmfqDGB1etcmT
P0vScM6Ec3D9tI/gn8cc3UscAU0zjAoRPty+8e3pZfdqeCHsXRXFJ91R4+U5
xxKlioW2eMN0u4BSS6ccos6tGn921BQpMTpmx3wyh/muL0faJT6zZJCTxPGt
pu4ip/5K9+qJXIIDOysCfnR14TykYjsvZYXYZvb9UdXkts2pTFq18+BCdADa
q8AGnx4XAiX2H/1PLYe97I/raBSwAQSItwHwFixxY/djyEGa4PgDEslB1Xi3
5LcSSM0OYq+0p7XwMQOmUSyCK53iN35i1mpyEs4GdDohff5dDu3ScGpdlrTF
gVs9QNxPgudTLWLAZgwIXDSpWOz5oXPqq6uUlCWZ/hhJOVkrtQ17ikE4DO2F
sq1BSygZm3UFcDPODy5BfJNGphZ3KmvpIwqQILmt6EW5pRPLYfrES0ryMOpZ
3RaolwpKIAj55pckcMr8pabjp7B4XZe+CyFVRg9RkWWrFbva+dpIMTrvRVmK
TsVyiV5/joL+jg/X294QDxWPatmNgSWEevnru4Zsxup11ExuFke3H5WoHn4E
pYnqRGlJ2Jn5MjYntkPp5IPE1dDSHjT3TrCCa+MBUVvooSfQIBC8+GGme2K/
BoOAf/5ZVTLuvF+WFUXJmjiHbZIMAFW7CCZp6zO0aYTwp26Q+BLiPPeqrSbV
WAWIHlCMZ+PmH40p6eNqhZFzmeBPLClq3kbusI2KQYVBCqgpFo7itcJZJEsT
YqM+F5e1kmsBmHjUNaTyFTlZL4ZasJ8IWLzy+5OZX9qucHUd1deI/OVyOikQ
um/JHptEacVaLe7zqKS3adBB58nQ7w9yOyFQmM/OIw47hWGG6KafKSxIXD3B
KhAXnc1qwJhfZYPy6zeC1oSYWhdqIH+7haDX4CDiIDvNbWugrk2l/+dP1nEd
5Hcie3Qgyw/yy702hWs71WunwwOlNP9y7MNfnPTtUwVKxyvNbphYOPSupO4m
umaBBJxJJH8XJrh+KQS6pZL4ehbEmw7wekGAQYDFH26dH2UcKvJR9+qBjP2g
/2AYACB5AUMs3jyXfXkTWtSpICsDRiqq2JK8WB2WWkhbhvve7IbKI9nks1MX
6OVhb6eW48J633SGj7qwxOhqeaL9//vEA6lozcFXIzaSogLgP6o2q32eEWG6
bmnvlmxrK5+9romV1QkXuLUvlP0gcVVwTgKzSQhn5xvd9oXmiOqwzJ7zJPta
aSYdUP0TgjBltuW4vS38a+hFFkuu+xVuGULj5Zam3fKgsBVM/4N+FVBHZfvm
P942JjMlHzA57LGpa9ugH/paRSk9CZYyxqM6dEO2TF8vmMpdMtGxhctPW4H3
FSLS8hGg9ahtp26rCAkpGIjToHScSTXDpBSq4TVomVg7ZHhQMtUIusevhPS0
w1DBY28XeOPk+J2foaUdTz/FAO3jiMlzHuncXJelltCl7RrTf1GiSuYwYJMY
88b0s4mJg1DL387X6MUxVe2u8RS04+Cecd5XIDrfM5gxdJ2qasjL2/zPMfzy
jzbZ8QVBsqedYr+kKf3LwIEZ560rNrjhzOEOCMxoKrD/Z5B/IIRrdt66bS88
cpWMuB5TRDYxyauRjd6czW7DFLWN2ZI6vu8906ngHV/VptJxqDGSsVYIkEt1
nYH9MZAP+DTmYwd+puC7dbTy2CviT+caNh6uYq1QvtN0ilY9wyUfHgKeHOws
72Qw4NfxkVmHN6f5k/rKBnizfOOI17sjYR0pP8ju4NwU1lxyKNa0IXXTqTnq
xWO22d6WDSIP2qSyHnKO4nurGaffNHSBx146fLOGcVN+ShdG3ZXcGQOXJX8P
fFn78MSTAA1sTJGjz7aQpFqMiBULhyXf9suMlL3hgVT+N/p4GYfT/3QPoerV
VgYHIg2IJOwgQg5ObCDo/Ij9+EBrrYkf4sDFRI5fqqDcoGyBMthwaEtBHYJY
EopJCQdSrkSP0NJ+dRADYgj2m0dJb4z3XTdm5aSDrHp1gebdrZucYyrxa0bq
y+wRtaTekaB456ahFdW8QwoN/OI6SlVGbCd30Rkvp7kUPIfcqf1lNB8W9iNE
2ctw6YOTJmF+PysYnVVOd396odWfnGMxSeMCYMKOgenCiMiZ3wxZaBL7LrNg
hLq97z1wbBp3lMu600H7AqGl33Rid9nvJy3FiD0tCNFdhv96sXeeMf0/kO1a
/P6Y2+TRChLq+LMXIvzvCOI2bmH4NmTyAGUX8KYmafk6FlAOrCcmsV/E9mgM
TlVAPmcdP81NNpir6ZspvYdICUxkDOdFTzqeXFmNuHNTN7lytIvuOH8AMUCl
GeeYasvliZnIDYIHzE89NAwsOcPLjz+rXmukF3FqcweTQDdYiZqlJrYa5nU4
80DWoSSNOhZzyMk7Ylk+xkE1RB6FI9RjL1D26jtLN6MWezztyF1EMr6YVJ6m
Tivx6bkXXkkRYoqXiJoeNbxBW8Gurz+CcW5UbL0HQD2j1V6AM2F7lqOiYjd9
NLqOIatKtvDAH2Qr8QwfnELXuuj6lXeIJImDOAULzeYnvIq0A9+e5W3i3Bxh
ET0gjiHdpDQpiDoeFi3b7ipVRHQR9YO+wsOcGyNNMOxukadxBYXO4E2pFrVl
j1aLT4yQB/f3Q71N1AW5S03fB1UT8uoU3ipfVJd5IiiekDhQxwoUKpIoVzLc
61RK5qX/i6MXK/JagpTC+50NKrV/7uW8BJZD19HZA5yEFZ6GSztafCYOP8N8
CtD1ovvJtNky6bqorT07Xw/5e4HOynkEd1M9OYACUQKyU3rP6Ko2mpGUFk2y
9ZjIbbYVzK2Pk/ffmgArbsZn+xfJ8eitf+WtvxKqZ8Z5yBivNYxa5lYpPnta
WU/Tj5i81QO2h0d6rvV4aFpSjYXKB+Pujkvld2vnIiWIs+X0ibHTd92K4Tf5
+R29aB9P7ZDq9fJg3D7bntedqqEB2YheX/dn2ooQxdjc5YIxSRoc9mDOxFS9
IfSaJesNnpjB/ymW+7EMWeo3WSGPLtIRIq7p5zoWSbiMzXgn2BV/OQ5n4js3
DhuPq3aJf9+L6D688t2Yqo5tLf/NPB5+B89Ny+zeJ2P9EwBIum/raAJyXgbs
gIVV6HhVGv8w9uQ1LX0y1jvTg5hLKnbV4gCaT+fcMgxq0AhOp9TGPHkxbnTR
QmcFYMcl43Ex9ikVDy/37NkEnqgzhQ72DxcCwM8Vg7t4fQG9MBtYHGvL17ya
2p9d7+QKUOUE7LCAfbpkGhP7p346SXdxgYtumbJHdhh8qQUBDNMLxOq0+Cr1
5hnXnydVYYxMiNYctnDwW0XZ10kAZenAe81lOPALzDdxTysoPPOwUA+2YWNK
fGm9lxojqDLTr9h74hh+rL/Oxp62EFx9d+sy8Tz3Gx7QCd9JqVGeB9Cw/hX4
zPwiz/uOXpZA+HAWokBS+SOp1i2/E2Hl2FKfIF0sw3UwEY+r+bIHMB7MgzVs
z1PmWkpG69o1erCUynZYNbnZK2tubyIYOK3LL4J5CYNBVv8cEPMLGu6eKNE6
uXWuoMPycLCaSKQGr2ehCxE/9J/4Ulv9/yFSSPBA15ckfItI8Y74ZfRcPP3v
qb2ioZLYAJXiQ/nhYoMARvSP0wpsxhn90rfjpPjM2LETJXMokEe64Invczub
WTKEj7HdiIiM0oE3brhWmQ2rz/kD8b3R2oYlKM9DlsJaVbZ0zLoWw0Zr0yct
f5E8RfOrSNWQRzyMenfdXNvjcxh8QUHMRsY1+c1aksfIsF7w1vwt9oUPinUy
V6NymEytz2xdwWfR99KFAWvufWNFJk1nuLkb3m+NrBBTPXy54Es/26D1efyp
WezAEXCgnw77qH6ZKTejGz2OwP1I9K6RiALSXaMyAO0jlWjzyKHTBSFM0Oby
pUo2hi0+jt4Kh0SLPqdasa/E3CCPYhfCgtfLr+64U4doNtAeUdDZnlIWvmNS
juSURH75NY3IsAJoNXQDlrbXOFDBTWqkBAchliflOzoJljl3xm2N5Ppfngaz
y5dA6hdsVqgLmq1Z/sZQUWTSel7NxNPqemKEdMMrFeuokncX0IGjDwLejCzH
UHPI8261dDIAlt/+4toDGqYuGkl9RRG9BW50D/C77l4gsF3bpE+GcV7iWOfi
j/KlT6brr2kkvSm+ZywZ5NMYqb4ug+FJRCBBmMfq7HZIusYuabzBevcB/H5C
9YQQvC43zOr/es7uPXTYUsisLk4FYh7y4t8d6PlmSNU0WfpuAZPgaGJXu0XL
BdFIxRspodt4eZbVLBsmS0kOYbYWZcbzkGKH3S2i7DfhvKMWEkvfXV7dmrA+
RySgtrdLmmbF9sjmzaXct8Z3emzoAM3VW3vjjQAW4gzVlf9HK+HKmIv55X6x
9B+y3QOXtU51TNBLc2lGlQoZ8rgypYZy8DqQQ+vEnDL3FXRS7RjLy92zNCvb
t6bRpk3uV8YmrLZBohz6mAJdtzbQ9vEvefTfFiXyG2I38w7OmceEqwFmkJCN
VHj41iDq+39Kh6OozymnPjnu0NLivGiLlO7z07FF50mKyPDH+Ey4jxyn4G8G
NjAnCK8JJL4lX18LJKaHweS03a1mI77bS+Y6wmx0SaN9XsP5TnWC5qoYkL4Z
Lxke8te6dYN+IUU2iRqEGl957zUl8T/WfMtLXb9B/wsnJpm/IgsFopHTZ+pO
lBjH4pvViuDI2ZnUpVO6ckzHiT8QYw/KyZE9T8Y2/U8N89KF1NVaBft+ALl9
HSCeK5nmgOy65rxj+GOMEuKATEUk9WJrFaLtwjYyG2+SDzehxe4eJdPchNAs
p1g0llkiumvA3wPlWo/GpzCNPzNDpH4yjUs/jIzH7iY4ncRznbcCULNq2c5t
Czt+vO/qxr1Zza1wtS3PKIzjGjumxTPysPPbKRW3a1+UevZ27mXQDZ5AvTdf
h6qyAdiwphXaS1Oz1k89ZLvwq/tvGNNlKJBdwtl6GeQ2SXMDJIIZYcv2s41C
mj1wNNvPRywIlJ0nU2/eqbCb5OPiA631o5us7GVqAI0azuqoV4+hfl3nor2c
TUlfHLuDrYbcJJoUsO6YYuanl8cTc503oLmS4e0mP713NXMLcXVq1BezhCkr
+G41Bz6CVmXXk9FnfR3AYi/j0jVUH8HFSk0z6/pV3DasFUXU6DrYEZnUdR7i
jSrq1AVyJxfZtEAnlyaVQmVqzn7FNDDQLxINzkgLvzPpxoHYQ+xb/OlkCoM2
D7duq/BJ3+S/nL0kGaIJmDv0s2bHDnnHhHVr28EiaE1MlOllmmRyauYyNp2O
zM38hEyKCtZyuxkOVm3DOCTAFwD2kUvFflKFutzsWexUinfESwvuxZkuV7Pm
7SiKVedoQl4bslBTdkLDvNyIYH7pQleqI0/vTV3DlXo6NCl4UwGLahi8BgGv
SlA=

`pragma protect end_protected
