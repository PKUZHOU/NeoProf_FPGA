// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
WPPddj/HOcrlUuGPrhTudg6NUIvxaBJWrSr76GzUZA4DaEZUDHOdKP+iyf8eNZv0
J0YidRuzYVguRZb+DQeKPCsVL13iIsXkPxW5cCVtdzl6Yx1mBZWWOtyrTuO2KJau
D0Q3726fJGk6BVFuzCXVanWOCs4S8+qSZ4oZnblUXU0=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 8496 )
`pragma protect data_block
Ba3IJ0tg3Z/a5eCY1V40KTOGV9r26cpLjTCOQepFh815YlQ1N/IlE/rhmuij4SL0
rzMLRKWiz3Nv2phrniDn9UKjRM7XOvzeSXiG6jaHMJmM9g+iCQ0WOiTe4ZhNHKqQ
5VwgEUdrutiBNQWN1InCVy7FuOB7HZvjzSxRG33XzTkcEbONkCWzPDUEhOc9BvGX
/bXcWtmlbq0cbAHX67bEU0ER9NuXlSeklnuXrc6lUh21aAjeMwG9QtjmVTS9q/6r
WpEhQbybhwB04rjyt70K+rF/vf4Xh/uAqqtrFqFMPVkDZzLxryvozZ6BPjQzI/kk
Z9L775jEgqRaBqLcL6rB9BUCDXoCV8pWVsJhyTyZFj2nmwDPnhT3l+CTn67Po8t2
Qg92Qb0oDrxAKRDwLaGmlPCkClzTXMHYRRlTM2yvp1bxiQ5U6CUqV9qNwkza51rH
AWWjBSNyl4UBe0wY3nYYw6kAI+9y+bpT96v+ZluS+nj4n3kRNDM5sLORkg+qKgZ4
fIU5MWjC46X9bcFRbrsHftRq/upjHO/Yc5Z5XeIQbn4LuzkllzhgprScRk4z5pTw
Oji0r80epkx6lIP9mSpyXslCnTfPpDIHaezh6mb4eAPvfqg72T3GxZEVse/GsJYA
8LQCUOcjdl7KsjJFYwITrEjzNCgx9mMXrRCCmnEO6NRlpSiYIKT5vCobLnqlFO27
MPHaO18AFv83/9WFjJBddRn82xBWOVaa2H16ySVu+HLG9Qi5iZIKW1e8Qp8AMn2J
/9zRGxCx7hmPxoH50ZK+1EPn0Kx78Mh8vY+81zFnVz5ZKyCCBf5DU3wVdBZfcCtK
AJsr/M74lyROdUcd0EJumAqEhsHiVz5mrA43ldmrJ52UkWspBa6DMdyn7PBVomYc
G9PV72nzlWTfulCuRAXkMLhueSV/7+bgdBVFBDnODVH0hXNme+Ka+AVkG78FSA20
VB5Zp+A3WPPQTNiiHAIfDNTFj01umAXKduTSn517qD3cJ1kC9Nq+gRMoftR1W6Et
BpAC4NaE8RkQo2Kt5hXfHYD4XauiC0fZprnLNZJ3eHMdgOul6kVEPSVCHSUPhxzg
X09KR2lvdnSjNva4vcNtoHa4MU4k6TI5/TMu3BlhIMhAuK8WGP9qr5Uogtbw5FFR
NI4YlCIPDao2TLD+RkKbWe+CI7qAbT2mVCMjr+GJgUJo57XDHnlmj3/GdzJpCAc0
1fpXC+0YpXdpTV1W/GA6ZUNN+awIeShpjZxxk1JxpYJobON9iyThcE5K5xWV0VjH
8NHAQ9PJiNWr7EJtfI8+dtT1fNjTJDtI6mruB2EVGFnsKJ/LjSiBCrxlhstlneEh
4XKRi0DRfjeAnj69sk7E1GHHqrBfMRm/rGBAT0HEMInm89x1pJz3xdmJE1DomipI
455bHBNCTEnDn5xmTY6gTQapKiequJ6rP0oqt5BQr0PWvlBRuSUFY6+w2CbygMc5
NhPcKsStXIW76iYybJEDxAmeldc7DrSkcTAL4UPvIGfl/BsxVwICyflU9+AHiZUl
qjYB/KJi7Ju171lIMs4WvVTjQiCmOJtnfniMsnwcpUse2MWialPgOgn8RMaPHmrY
kEhk7rJZUhABxrkQ68zBpWxh7awCx+KDX2AwhJBec04zvJ7Sbt9fRzZKZq+ucLSM
euhHX7oe1FotFelDjGtGfi7pGik8Mqgu3EwWACfPNyvgRCZJvoD/pfwqCnu0frjO
wswvwFvSEneLU5hi0h/nCgFwYZEbf+aD/JVCD5u64jglqd2f1caAUincx06B2wDC
Ces+eyYRFDJXNyLMuLbxwlq0+KbNm/c7o3KLO/KQfHN2+doCQgA6/AGqknnlnaXz
hKsXOcn/UfTGpAeshvzBtpBIXNSatE70WxxKlKOi7aLbWpcdnKXvOtlTJW5AAy/i
ZY4vDVTH4UggR/iAx14QAnX1ClVNaQyfE5QeD2QiN4izuRNxa8CGYgQNxqNvtveR
p2gb8HgGKUjeUHELD7fwHYZg0lW6x23DDGXbpOkvklCDgz1+KBwdIVtyTvoMIC3w
ivWfTcq5us0QE38u1xWKHI+SpGZFLJASeml9Zj4yWnkgBW4eM4W67Cq3KXhXt2VG
xwgpsaOkfhl+mG7LxWQUaQPK0lz4f/QACY1VIO62CniID+5yhPRe+Dc1ej7jWEmU
5282uJUEFeD15mBzLB3C5POD8Cf8PGjwSSJ9N88hhi+ZJHblBeFNPNuau+Fvtoo0
oeeHRc71fiwJRTCkwgKTmiL+g6EjKCQ/RqDXQQhsN0q80QikUYYnIp0wDsfte0z4
9IC3qBsUTuUanlWDWUyPHNv7GN5Fion58IU8XI8F4T1/sFRASFjHTvQ/OcS1AFY2
Y4QG8GC07Bs1b6Ji+bXIoSMiN1iKheGoHrHtvURk3QaTYa+Pwd6w1bXBxaNuAtm0
l076Woe29NeGlEBXKLTOZeh77Ryu8pevUtJ6IXa2LWCpR5Wn2hpswK5Ycqo6ppID
R9EKGoLrm4bBZ3D/ExGfmRX3c22G+hrfqHH+EgvzUYaDk0ceMh/ALaWzZnk3w6U9
OP2mXrkLpQuIhAIzxbq1aC5tzqPEn6ZjoAxyz7JDrFAmfrg2dMV3nPlgH9FuX91D
ymy9I0JOk3J7bstAYnezlcdIsppRuSexj4pyE2OXjAEO/i81GaMiV7EsrRMEOr8S
I3u/81yqFlvl1kdUIdSmYX+DS7Idg162XQEiXnPA6ODdoLp6I3+OkbL35FLhLjwC
jzY//dbVnrJQuHebE49GLJ0KLHv+OzRVg5dBQeMcIdkurSBTjxXQcgCfj2pMkxPe
dUuAZBRF+WhGAJRf9iU55RTZl5Jx8HaRWTT6OmCDStDw+xDAQfNtEkboqPKGJCEJ
a/z9EP01WtznEVV82IZeDCOVOktHFdNBqr5P16j245FFJm9SbZH8zoYmP7IrYvcN
rYfiVWYmkF2kNvyhKb7CjOAOO0Joq4dsstG+iGhUF0f6Rh3o9HENoNwyfJEpbxuO
Unn9FMnaHWhaGflGEZ/79zYzpFGlKxsLKkA4ZJfCIJr7bvuUte0roXVX98q1vud0
gTsGgZ3uhLpCFiQOm7ibwQgDSajpUMDfQXF2VyqvEuXFv9WVKAVTToxnawizHiqc
6Jl3h47QL/+sPVKdcNrdx5Cp/Jj4yt3Wz0Dn5XOy3Ub006klw35POSWuiqUua3NA
wFRljk+RvNFPEyxrP+sqCAgk6lAD9ljgq/1EhTSSpwNuEXiajBlEmODwPkYc6L+8
J6i1lapgxVS5Cl2eIsnVF0KkHrn27mZRX+WLChUecWAY5gAMWOhxTYbRuSQp+tWt
L+tCtPQRqaGPXD2oYJEYjEY9OAIygyPcgy4YLOvenBjpfVt2R/I5XbxcLu76deNk
+jiN/3tm8kCko7Exa0mPz6iKvQv3LfpPwZlhWZ24UAqSF+1TonhXO7e7jii7l5Xo
RjBcSsUo1hgfKWn5u7/cFdoiNiKTjIlhBpenxqL4cra7LA2OOseZaGfmb/uSrSUk
aHu6g0hGeREmYofdjQJPronpuVlYZrkcyUyRIQ6WbPMtQWkwqA0+0/km/ISBQy2P
sUG4kajP0SKdQUCjR5YlICslnuqsST/YVtGs8pDuVl6TJraqbbp+aLccxl2EQiIO
E+KIy0xLLiMnTkY1bvm11Oog9eLw88HWPmss2gjRRNwHCD19dYgBqCrwgbXF6Gb1
SHzvMgiYMvaN58zrGclnB1aGsOpQHtyZDDGpC6jkQ78Csk7Ofp+AqSqQDC45R9De
0d2E48YUBVyHZ/XA4SAlwqwX++TOQzLMWdmWpvPUFRvSLcJurBhTeBWHK0HTAgcX
1Z5S1oM2tCYlSG5b933mlMyKJMX2QHRw91GpXCyL+1aJ8a5M2V55T8O8RUgLdNNx
lnKI0S6doszxc4AIIxv7hNAJEjxdJLrALVKRwT1oxz/7lU0yn2M/tCQKvDsUqYwN
oT7x1MO+K+jN3lc5aV2+qIyg5yaxcgduBYurN+9rId54s08a7HB5cOhkUd3eO/KE
f8O2FCU7E0+mEvWQd4DFAJvF+mHtSCX0C7Ij1zuwPw39kSlAw8U0L3C1tg6T/ZBA
dcJL7w8VyT/tqrsZEPxtWyJ5w8413Z34SZU/GbH6iUgOGdZh9jLAgw59WTpA1kyp
I0tVNWy7ooLfEBOPKSYcKww0n3cCL1hSUm0SEGB3r8NNydMMxh1Sq432GCSY3mn8
NstIsWygJGLFhYP2/u5pxNUKFq06NxcK7Bsr4oT0F4aKDB2L3x324BriYpLJLpl2
P3jYwwJ9qQuh+CRVjenIi1Skl2fj/cP2EbmiuaC+jKoxsT24Y0n+E8X1VsO/VJN4
xMhelEpJBRczZpYCtQpvnvNiOatITJJc6RI7PBhyUUkYZ+FGrr5kjnmXdqNtbjEX
/wl0G944U2CyBwFsB9ysj0OM9lDxzVV1uZnam7Q7P/5XLLUSqWg47k8Dx4626aX3
FlYCGM3a3WjG2R8XteQtOB+kGzTt9cpFmg3JAGfU/Yd6TWvkzVa4J87dm9KGIrc2
SElQsg4AnEEDqvsmyNfkQbbcSfOZ7472VGioXcl4h1vj2oPPcBcZaB/RoLLojhye
2JTk7zcWKX2gTmE2dIsmaJ6e6rYfa2JKA2iXgbHJloT4DNB/dsdFE6uU3HgNpv42
kbk9wIeNqL4VKBDQMPY9lLmBEWWgPzXAC14pgstkRM7QWIbkB1qlcGF/5o5vYd8o
5xQmcz+9sKnm8y8RL0EiuKYncYuqCsH0+zj+YmmP/SH/xEYECz5MQttyFNihqDUO
XVm3l2V6a66DN0GQtwfuQTSxm9tzydhOKoLSkuZBGZRE1f5o1VY5j5ATrRsLFzs+
jGIcHtApVTOxlR8DVysjHboOSsBvawB+ns6Q2itJjThWEd9/uixm5lzSsVFv5tDp
7UnTqZRS02SyoHyHBlMFmCAW0OfRnCKOVXznlUMoEUQ9fGbpxQ5sWisy205UwDgx
OLLjWtKSeTCnftv1gV+u4sn1tm1GvB9SZ4p6pqSCweBeoA/zI82/y7CIK0+PV8/t
AkqAwAMCYX07v5U8A86c8fDs0UKwRfMpzH0bxTKd89nC9gFXmWUmP/nAul8OK+qr
mAAwI0BRXQYHT3e7qO69evjs+kK0J/qBxHz5utpr4f/JSoV9Q235qJQB1wQVDDCK
LXRy88mRH8iPMX5vZD2t94muEQ10G4qSFGi5TCoDDe+wQO6HO9uSaIPzTFhRZGdf
bIpFfaY7lau6yrfYaGpq/+eJRJHG8WWlW4vwXKP0Hzmo0Nd7y7IsI9TXGaL9vDGN
iq+qIv1qJSsSonWOqijqcfbOdzpYR6fMs0tRPBnmh2mT1ecW4Lg0ffOzJIr9SOSK
I+p003XFplHILbV+t7kgOnLyeWihaRjp3h7dOEmoh8wEWAia1PUS3m4US0BywjNf
Kf/dgCIk/Fq2gvTlgP1xb+11mLbUCoPlBADpyIAe7hy+j/pLqhqYZEP27tsBEiuE
ASWCYvLuuwYArhKI0SCakcIRyoE2HLUJlXOhxhIjF+fyO7Nf1IJId2AntRudPzo5
Fpdbg1ZJbIzYz6OY4YCLxV00CvvXx77n8WoSz1uBNoklj0lsz6YhxoLXs5fOU9VK
rFd+2YJBuwJGyIELEaHQaBTVEW+WDDgBEjKep9xxeq39UPI5n1VKRH4CdKTs5S+z
EI3Il6nRd5jVlYJkJc80bazK0kEnNxr5edcShYUlp/IDNx2TEleB3n4q7U7Rttfi
pxz12dzeWyczaGZy3Ab0D6raPlbqISkg4ZVm45H9Tl5TxwEVC8hHO2VxSg7MSbTx
DmSBKbVA+ZftDZnBNj3t1XjY8sH0cJGftmnJeuRpXuIIHPTj+wHFZW087+ENKjD9
KtXM+0NcTMAodsCwcZtbaV8FKzNjxrZIsI9AnyO6ZcCKe8+HIVJ0u6OJmrgRIYOO
mzUOx23j/3pkEJvWrna8iW+okLAKv2NoQXA0bWiGQo8QbjFtmPkOOYMMHFBaoO7h
QQs6pdBBcbAh6s7SEGqzKZJ4VMEaSW+4NCLw1wOPvLXWl8Ql4XY/127Ztn/ZDW6O
TOgA9DQj19wLiRLpyMCkUwH3Fr/jgKIU8cH/y+3w8V40JKmocyWoePyFL5WGBpCn
qUGj8elEU4m5VEdvrsJGoBqoKbJMhuhwbcuHnwqX025V6PMuC+LfrZKH3gYLKSDY
uu9xjEyNoR5U7hS3tEdmGgVFJXsy+8zUDirgGeDidbcdGquIc7XKIa7NfOZ2RNx6
2LcTzHqiekawY+IYPqS2zvKPaY5efauZSAiPDWR6iadEfmt/ZOY3Yd7iJ+tcNPpC
BEdjOVOnCqBBBeQ1CXwY5sarPl9vtCu1ZPsED9fwwFzDIaic2wYlvE7JVOx1cKtf
hBh7pWKHXkEC8NEqKU3EAhPa5NFW1VrxvMRW3NGNffUTbFDguo52+MkyJ22Nx/y+
oLeEd9eMsBMGuCwtsk62y3xB7AHGWhyOXl8gUWSpYBLRBK3+l5It8gd0zNQMkBf5
EQk8CqOxtqOUgaGyCySh1bFrW9nPSh4mrEBRW+qusSG+P5GRtbw1JdrLqhbkEVrv
7AqQS5/p62/cyRLgl1XHYkNKt3GUZdtFHL56GKG23fuHZhkOKOgjOhBGyy+9QjCI
8Xfb2alJPMMb8R/RCzTR8GYrh1TiPERwDppyZbjlfUNbvnHX/VQ0RuLc5VRGPxmn
CQFpZKDRZOOEHwrsJ1iia8SevrMdvN1+BGxqyFAy+/iJiFFV12lFBODaikrNK/CK
By4g8RlCnmlzztIYLNCUuEeX4l667QHkvk8Phfxz8/k9/KIltZCJGPUKnHBjWkPj
xgyQkZnDxWHm4qT9l3eW0wtb+bH6aaz0NkcEyNGgZi0jOTT5LRdD343Pg7PZT1Tt
Xq1DI6wj/0TXlIEka1NUNwfGgR/wMrDne0pYNXd4utJW48Lz0vJV9YhOTjVnb6Fr
hH7Qf720iTjBIjIK58pbjNOb5JABW5fe0ESU+SnQ6RD3pStAuLyzCZtffF9FB34U
K9oUajughCJnnQyPdi5IJ8wjg8n5Ayn0DF17EtbwCUadn2rb4etfgON5pv93/6JP
DYX3I8J9bsxYbzw13U7aDIo5D9ZpW6qLIoEdef+7s1KnpiO32mc9DaLtD0rzJ0Na
fZg0HRJEC080JjKxs+fsxqILaRapI7corBqUTWN8BVeTqe1WnqBX5ljpB7iawQal
gPiWwK5BAUME99L5rgfhkUGLGhVWf2dLIRR3wrL/XLvaTiDujFE+PVg/FZ4GJs1z
E4gwJXpFV1E/FAfMR9BiHPHhGfKQwKwijEuLGWdyTjDQ9js4eeZAdsQG7R+VqJt2
rzNFFpovYCOngNPV/IaMJn0dZdXqfAt4+L5doY2w5sf9RWjLbSXwbHrtoeHG06ad
+Uvf+Q0L7FgHfoRWpfmVMiiCezGZoEM3FkYl06a6+cSnVCa+z9Uy7J+eR77lSJ9r
7Nh7D30/NSC3OKBds2LktLZRuPJDoEIeFrFzTYGZBhKllqQFndbrQG4aQObG/80i
cj1CV6VTtTMuZaY8wskpv6mGlDu5eqeEZyKW/rt5MdSehz1gegGeOIjw5w5kOBcY
6I/PZiuUjtAo8u768gyg7Nol91kgCBcGST+BZBn7XDi5egT6AhOcWoBmG4OEYBU8
iS10veYe+XfLNXzCswrflVaaNInzLT6ymXvGVOyu0PPXpFy8+4AvheuAmMhRDlrk
HGNkoMlrtCS8wNZbqAIJXh/i7Nevr4T7T6N6jzKoly6vqfOXLZp1KM9gqNFSRdr4
Pwe+rCLHQmpsGIY/voik8BQzWnKe8AbyvZfR9DwKj4DBM7Pj9igqMpiNJ5tYaf+A
Dhd7EoHqTYNTZNwsUyZrovWbXarF9rUpcWfj4h2cQgj0W8H/fGiH7qj5N5Y+J/DY
EDx160db6wgGrXpe2MzXK/a8gFMIynVJSdQS5rYg6TccJr8AuSfDpiGCx9ozX7Cu
bAjxVijqmdqz1QuygXou+sXZ+QfMM9NxvItoG14iEuPY+3f0BphIY9rp0CUH/SPM
xcw/ORz26KDWPbxJYR83DNF5ilbKeynXjj7l4KEsWROlnNEJniPmPpymhMG0E5Rk
CE0gP/yM3so7JhSkf6cLCxTAIq+ns+hRv9D27Db7w9GHkCKpola0f0kXaACll5zF
ZjkPvGlhUKNHKuddhBN0ftyYSLZS4g47uBJiYPeuxF+7N5sg+dQkP4EGR3qkafZe
8M8eOPZfmJuf14PYInyXxh2LNnDBIRNL93ITVcFjbhq7BJJ0/dVExIpm1KSEkBiR
1ZLcNMQiH46gXB1RH2/6zhIsMa3MQB7VgA2avJaQ0BxdLMMnEiK600Pfgv5/lJYY
MHaak1Inaw6sceAtOY/8jbh+WAu+CxZqY/hWr4aCvLvayvCGgEcZElVioQM4EYf+
iBuQneZ72ktbbGpNO15LkJnSiM8BDJ+QFQHk+uBweRQg8qlxI/7X5DdqJ97YHZpE
LYQ+qng6g1oiHE4BktHCsLv9UL4kYVuHQMecZxj0wFsq1ubrY62hirAEsF0nh0P3
0MinBMCco6Y04TtzWTJ53fH3ah28xOPq9i0lTB7Czts5C7H7htmStMpHNyd0KJvU
vozVwNdruA8tIqupI2N2LuNxMH14I2Ek2ubKTlfJJR/kH/eoguyIJi1ZNRgk1Mtw
4egk3JnG+g2k6iSbSX0Yt3jEH887+sGTFi0cvHGhvF+ypTlZJA0atHvvoPPxm46n
lCS4Y9IrJGrWmq1/9uPJELlbW2TTm1jn6gPcZYdoJ6fUxjBb+GQoLdpW0yzY/dEj
GfZrfWw1mLMdSF2Yx8DRyh5tY+5vp3v3XEUTe7Insvg8f71NfSL5OJj9r2CySKdA
kqYr+LNqHAEUhOCjrb0DFWN2Xt2+vqQPgFz1CMTe3jkXnL6FyO0v+xino8oGGoJV
tyO6qWp/eA6lw51BFwKeJKI+ZfZfH5yb9AM7w70LLK2BSFg4QvtxTcoeR7kT6lvt
qTczgGwSb5udUZ83kEa44OXsAWOniMsJF6BkqISC1XIRKM/uP15nZyOYKkyCRlzz
OY4IzpCRdHDYePO7fAjyHUTQoBtm8J2nFZN8zLl+CK/EIsXIcK//oN6n8BpswDUT
oaUyhOVOxdaPRp5Tnk5U65ZLk/hRDWhF/LRE3Uj43W2gW9CsBpL7mYzw8OZbv4PX
/LT+YPh5nInMQKum40tqxMMQKClciu36bwqUw4M1phM5bhlUV6B1mXsxkbTNIKvk
PTtYgJ3VB8p5n1NogYSUXw7CoFUC/2mJoegUZIrqZxItTzWEnYTBI1RIrqnrrz2C
x3r7zdnbYMVVAgSfK3pnOYKclVZHpS/NHJof/B/PKFLwPHnf9e7lptRrS9Y+M1ZU
IBomLQIg6gV2MQmcG/fW7Ji7YxtKE9nPMY0zKWh2opravXDFxtM6WUZTBemVuCCD
2459N3jdYPX5ZcFP62WWusRZq1bCtr3HqgMaETXwtqV0hKHDZjvCRggjgwLtmEIT
nKLu40QWIQW2u9s/WMskbvZ7H5v4daHDe1Yp+r8C/w08uCcCSFZDJEJNCxtkbvCy
yIY+je+dDl0GYFjv4dzQZCNtzwjyvYIzXAfC3UUO1Ieg61P0lxjSXSfGWRlfCXJp
xPsgck0JhSngP0kwyISvPrWhD+U25EA9Vz2OrLh/rQIthNAAvhYQaEF4ftLSJRg7
Ixn5D8E4zB/EPrReX61P2V2nE0/jWn7NzJSkjBjVMyzxdE3LD8VjeyylomHXxdm+
e36XFXEZyc5YVV/kDPGoBuuhEF8f3YD44SQA50IPWMbBY0jSKDKegKaOoj+A4YLG
jGNeXPA/r/GNt+0jTLPnBS3yK4eX36npNOV2wCgGNh6oG0vw2Z40qy6MZRwN63mS
t1Zw1v3OEoQ/5KUCPF5Fi+VejK6uxsTxnnY8kAjJgT8fEjhyVVIMWQl2DdQ1slc1
2idYTfyKymA/4O4tHvyqoDB+s4dWLSnCUaRXRu/Yfm36v89lQqGem8WLpDKelft/
WKbKmMkaBeBBeoqqTMwkS3dHk6GSX//tyZyD+ynNhj5LIl7FURqVBG1mHUhikbOJ
+HHU5e5sft0Nq5/p54og9rBpQ0krSfz6f8k2QnOgDMVvDSvH3db4MVcSG2IPyCvT
OvkEekrJr7Ls21Ph4gUvApSjIG3Gu17zlF79oc3Cl3m1VqfcYRdc8mF1eqxO3Phn
m0Qeo8dVPTm7aREFz0HrdFW4YZVz0KGH/+Y2YSsFEv4yw9K/TbouW0KAb6olmc4f
4d8c5wx1yPtxRzNyXCac73G689PgEVUcLId5/bBYXv+ps7Mpxw9ksGeyjkPHoTJu
nSSUNxq2CF5+wIqKQDe9744ceMOUZzMnwDn4NMZgqzUm1AYAYzkOsk1wD/yuX3VR
RytO8e52/tGQV7mlCj54sVgzqAOzHNuJHkEDZSDr1Z8JWHlDiCmQ+YCEB42/+YU6
f3s6GFkVOKLO2ocj82DcUrBGClZufaRYns1SWOiWh4WIAmIogq/kH4EDSU472ipt
6jerqsxHaDj7cL2GlLGTwk/PH1TWJqrM/pvgoBHhUipTOa/ODI8OoFlTEYNa5L31
KyS0+zHNdrXMpyYw6jPNEhwMYMZrT0Ok6XuPZa2kzzMRLMXJgyiyChTJ5btYt70r
zbYDOc3HhxUa5oXK1IMBSEFrX75PAgmWl/BmIpHFVGp8/zz/R48nfcLs0gAK6Ct9
bnCD1VIxUgM1L7eeNDFhCxykVOLd+z2UpgNOFZbKZ1hxu12rWHAigVNaVnJh996Z
0dkXUUAlHMuo34qd2tOPwNmg8eReD09638iKlKhxox0GxSp2I6eJUG1b9XdGJrpE
QN8UwnYOtcJ3RyT2ZIHj0LpxGfs/dwbm37zJfPSXkzXctzWFGm9wK5UmNONDIRwb
UIKbjGZ22kSKrpAZNvNaJM9xKAhhwtLs3lkJWG2w5GSS1kKg+4PJdiZibBNPvCeN
1VGg/BCeaw3dC1/b9NnsIrD9/HjyaMBvdMaY2d4OSpadR4LsHFk2xAkSXvWE8CtK
dkW5CkiQrJlTlPx+Zn1Ta06xisWSsygd0SObeQQY8BC4j9yv85QQ9/Lz/2JUjXCX
i00m0J3ww+YmFpxKvSSXwjskWUtn72EDZKn4//gARFRK3UK+eUwkOZ5eBdReDH9t
jlAAUc2iM10iAHiSeldw6i8PrUUuqaqLL4qxajf//oOF+TGe96o4HZpt8FvI6gCh
ZXG4dH51YcWSyQkTeXDyIDmw6qy2c/l7ze7T/qAvEMQZzy1rIZntRSir4L+3yiK5

`pragma protect end_protected
