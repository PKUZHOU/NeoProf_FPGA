// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
3nblXt5gi8M96+dvYuVvDTLvxZCvbA2IYH9TSnf+zUZomhxg6aNhvjHIEqFByu9I
dpNmGps4f2uG6vOqprLPAiVxtodme3ON4p5c2VuYmYeLAHunSmp0meArvlpKvhYE
zWMtUE9Xpa/bv3O8BQ9jX5kBvENmIyXvoTirerubcFw=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 18624 )
`pragma protect data_block
I35usFb6I53D7nfouHSfjTLW7LQ4CatsTFY+bk5cR3n/035Eeo7j8KAENWSijSxZ
GGBVNmLyLL4LLGz6BWmbkZYjTjkzUnVJWBByXobLg8gRbNsQ7jBrfnYABUUoUt+2
FvPIVNfho6Mirv9v/JENlsE6ukxaIdq2j/p4lUZQ62CnNxtaCnArb9YgKYyN8ZRz
YTxo345X4ObWUeOTFBVTXLBvAZZFTVe9DlWp78/cYlk/wgBkLSjCGauxBJM4DhTV
Nv6ZRAHYSpAkd1IesaXGJVbzPRHi7WsvNSTKeLCjgkh2RakH2HIYeCPTtdlWZ7aG
pTqrhIYj2pMECJrIDxTEhWzNMZO0B8nDgnwfpIYjqwp0DDtM+WqjZ5yL+MqnLiGa
0SJLYqNnQq1fSSE+Up2yx4yYrMVfcY+cj+BcrYqabip11XVKtn/kVW/pwckaYyUi
dHcS3c4TGE/tSrGeujs8sZmQ0b0x69T/JGRdDgLs5ioGJmiYZJ5az/1dEp5M6mFz
PXASRX0INzmGnr+INRtQENtDOdikj/fyKiJ8Ja4Bnikj/x6KrHYtZCFHRVaHyyyh
KOs6E8uxRH+SsfNKiJq3MJwHT6oxqHOT7oJKOPHEUgIn2sYHhSFK1Qv0l91DczTl
h3gwaNSapvnGMiVNdjKK+gMZL2lqjcaEY57iw3xPXERLYMsGgIx08Hm+4+OEUf/K
kwTejG0Fb8RUum8zZskWedjirxb9ByqEpZxFYSfMoz70Duy1n+Bv6OGlg3FdkRcB
uIsv0MVzH5R6aA+I2t2brNqUnm7HRazztJvbrV77KqRQeSzG+B4wLCwa4540slzJ
fQBBvVwA7/N77kQg65ABeJGYai5tmhVSAc+Ywo4aX8csMUH9Rp61pb/VuFRjfsZ9
HZPEPbf7ncO9t46vLDQHs80nbfaBRavKHnBYnPPfj9AWGWcC1SVu6QHxQprWgpx3
Y53rETjYb9AuUjZJXjmIdNUcMTTK31jzfrM4O6RBKsi8EpoJkAufRNIj865T0RZA
X27DaFnDgysgsQV0HByaT5NLPGS1N4eaERuDm+cb5MjFjwmJJs1M2QiOHYVJStcY
HN826AbHbA18BzbkTWX6rpfv9YvSxQVFQfF2r9lhQoLFZC0wKAg91hO9Z+FlV3Iz
QG2DRDlQBWU9xQc++1plTeGiJK0LknoJnjXCJatyyAGY1RCTNCK3eNQbTe65e2F4
KQzXPsYGwBku113LAmyKoMyRwu6ToGg12a+TK/O0GvXkJkaZSzaGRyGlY9gQt8eW
HQPOX7pduu3xa9PoWzurwgdWXkB+w9m+R8MKq/i5UJOKfHlTRHxMkIh/7VwRrNqA
7vAhFLrfb/V6+eqZY2+euz4FeRFCOUuxLZ8W8Ly7qKApGqdpL3d3XzBOdn4sVKf9
Xh1xJ199JKjIAOGiu02a0l8/A+qxtph4QnqqNxfqPsVoDQTlefaGUftWU5OoIviZ
1ngS0mwcrvrvcnjZq3ogDtAtDIo4l/u4riMk/Z1lVEFTj497dWcNXod+XzOOuxUt
MSfWXOghuCyHE2mmqTSUlf/jMnBB+TlMdlQiZ3KeU7axnJYccepQfoQcaepUrvzE
1iYaWPpBYeTmcIlxtDekFG46I31XNO/eFt2GlgqbUotTf5pBSc9xC0Ri+eIJM4eT
tJYu7PR1UF+Ur0+JXdtVcMViDhhNzZehglnzUfN+49KKYK7M+DCG7A7xPHbhC0Dr
fnGqsVqJIVUcLVEZXWJmRAXwdlslLSA7eAwFl7TjUVQj7vtQGjJm3zCONN/xaDQu
Ba8GLEpNveEynyou10mulyElW4lKBwmjkBT4q9CckO+uSW/OEzCp0Vnoh+zm9Oq/
M+txQcUooYA3+5WxUjISElTJuIs6OahsrzbL+r41imsbQjQFLWvJiEhrxRlhBKTU
Yyk/n2g/sQ9vAIBsUigxE4sP+aDTgEXHBniTHQ4Qs4WDvmy/JAMc5OvMBrO9xUUz
/KOkEd3sqghR5Xxro92S2kCCAC2UkmslhRjTd96+G185hY9oSugjPs0tcoNcg1KY
4QqyRw11OAMdXkARKpynBLgwtam69C69N7TMqCAsPsNIEmlBK3sMFxaRF+wZUHfi
bx2FQ15dI4tMqEyXeEl9HbSCH6hXaVqCaBxvC/A1F4sQ9XoTrVFfA5AAzlkg8a21
bZD93EHA5Knjy3wgOFsXxjlxgkhp/4y17WOolskL6KFz9zV7YwuTzLAmAZHp9SI0
l1IHrsH0eJqzeIPrf9wP7aZi8OUPGoTI0viY4Ef7pX3tbnFzlzodqoEHIZ8T/dIp
seuUYR4cMQu4yZ+KExGfXjCO1VYCfK7ec/IJc7MT+5LDkNxWIMc7n89ux1VYCvRZ
m/lbzY+P4KglbeoXMIzLbZbtBgZYL8qsMJbFKrEHWfZd71TgSIpWzIkqJ6peiFKO
IxoHzrGVT2KfAsYwviDdWj4EIzXfmwaDW81GEeYf0vcaG7X16jRdHog+R0hVDh/9
H6wHq+sEtK6BfyUQr2j1/sceLXadz0J8qQiSJisJHo/svTYXHqUq/amNblPLkEd5
hcYKPuNGrhLxc8H92eQr61+xBFRsm07n5VvCeO2F8x3GebbFcQyYB+1juh4LJhWB
fQl4lSTyMSQeInzSeaTrM4P7Morl5UxU50Cxl0QZX9l41eX0plyUc7oujWjFXifa
lfU4Hr8vrDDrFkIT4DNYlg3vgbAHYPHpPf1jyj8qKoU7ddVRW+pkx/VLEPFW1gzj
XGBxhbigTfQAyknkjfqhC91OLYnR1Hup43zo/Yk7HgirqRKtHR89QdGSz2t1Ls3Y
ac8gUSqd67EANcWqYGP6ahj+/eTGuHgf9o2o1gv7ohU9/4fRM+z3RAuCQ3ECDuus
gJzMoeZrjG93LG0EwK8y09GYTKO2P3sx7h2g2EpSnB3pOi9NHv+vrSR9cZzoZDfS
vIJ2KOmyytNQEb1aiFFbshpX7qHFJlDXXMCRtGyw/Mk7rGiv7EYBpf8uvEv7Qm9K
33k0/+oz6As3BEWUGZDidjMXkatcWg5JbCbTgmrET/7DmrHDfZiX9Ne9ADjJpdN5
bm1dJUpR0uk3BH/qR3Hyx6eJII4VKIJXhPpWqDfgUQc2IF44lMsHUwbhZBZ+wGbz
pC7jWv22y4XONxbfGKlHFge4cpgFQxSgvaBFhZqlLVopzIkV3pwqjVB9jYDYXzsA
qQ7LA1aaV5l11VapTImVAWdzSM5ch2fvykRcbuIkjNQh/haoWFuXTNcxZOkNPMxm
yMtDypkRVRnd/B1BlL8G81MrE0jZOrOaeTUjbF6KVOZyMArLx9ni1h1bqZ8DU5XX
WAjv3faOJS/w67Nd1nIwCBVlOkJ4kpz5q5ljYRVkZE7IR4zO1Jw4X/HnqYRo5abJ
EGKfQeh5rZ4K7/yQywJa5YDlQ85YwA7K+2WeO2k78BlkzxUUOrRSbtiBBtRp4Vbx
/oSunWASO3QwRtNvX6Nv7HpleTIAUQLZBveZ8U1GSAxA5uM3tMeq/ITezUhC5Ivz
cLewpVvjxTxCyvTcUqk7faIfvzXnm1BK5DtRF/dMOLEFb/K6FqUR5m8hqGi7K0K0
hU9F6Kh+Zp9ZxJpTM0r+hFyhQWWkGHrf9ctOuduW/It272bkr2wIThZCsASaWq4G
aH2qhvfI/wxEGoZf0o8QJwStQeL9qFNt3bzC/nJ3RVLT34n4A/v3sKnWHzLHeNSm
4F/KeP5Fmg3Xkwv8HAU1lnhbbkbCnYoyWfxdSm0R04e2wD7gKI/cQl0UhZy3nLaa
I613wpoZwFRQrKuje6+BpZP5eND88ALpN1MJsm1QgjRltwLY7HZ5rARgDsZMg2ME
gGRJ9o2tf3+2etpayf55d8FntpN+QAQ2fyE/8clsuqONcmGtOicsl/fPhmkAZs/G
N5EOdoweLnexugQE5rciB4tBgVO8/eZdKNwpS80bTQKva7XiKXSxuk4DZ55Mq/EZ
ODsie2yMJtFiKGhJU7hP8qi/pcjNqdKGUs4yv7YVMEjz/8zdzRt3bWaBkru8OogP
PXE42Q9xhBlftdAm0bq9NarcpgXi1WGLEQi3y4o4An4RqSr+IgccRYHz48qJTLaj
29ZKGf+LuvVLVFR/UMWBQJuHaiJ4HQFxoMsnLNxw5gA5gJm2urpWOvPCo/4Pn6IU
vuJU+UAd3zq3ydDNpR3VbolsIyAlqGGpPGxGLAlyH41lnVrMWupzQN6lNMUUd/YI
LM2bMA9DpMkcPD+I3E+529VPeUHQ+PkDYCY03NllRUk1n7wH/y0ZydZJG1pQ4XXl
6kXnHqbAIo2IdLypcCT8qHvmlRDXetoxDpjYlpb3hVoxPfbU7TBT2SLzmdTkpHoJ
+M7uJtQtpa7KZq65n10Fii4eXFZgucHMjsJYmInjjSt3Sa28Q29vBEytvlSTcSen
BSgcy74YvZT6UcGOG3Se37nPPmdwhEYCatbI5GX0K9EVRjnHGt9eanaStsfQpuyE
jnpTvgCR59lEiLOQu6UtF6qAEsNGA5Mg0uVeOMg1SLb8SVGm1e8C84V6XfhGgYki
W5OAUg72pTClX4gpNa+CbVFFlGzP08fZdxhTPdb7740BEYile8y2aTI0pUZlbT25
+FbCQZnFEJ8/zFS6Gt65ZBTo92vKGbF/D0o4rG6hNkoBLyQ6K01c3p+fB7Yqj3AN
v4NDppvOCDSmhjD65sybh/pb2PB1JNQ5wY1zNmzjpSfAnmeKJaSJrP7Qd6qhLbJj
JtN5CVaRIlfDnJU+fgpEyMkukMDUhcyBqDtCbRUujpORip8lieplCPHdik2c9vHD
9q3MhmlSJKNxP301T+x8naMWsteaKFcStPRP61mu4T34xoYofzGE8K8GxYvkJbnZ
oDbbLc6IPBHijLmRx9xAIssLspFFVPA8nxG5S/UZFgbnEKjwZabZgvRxphDfgs30
gDEBM454gAdzPtbZ2NqKyHi54iebpvLtT1hJcv1HhOJnBmchEt0WpD48wSW20+91
R8M3z0jFJXZ5iJrJwTsIqFfED79PagAIFtA1MrWnZqGZDpSVWB8JMxBHUiwlbmxs
QOL/fyomZ1skcFC12V7ayEujVEgoc6wwC9mL4tRzZeNEQz1GYoFfvetHRCW4aKyd
fCQkqzPFP1OIm1i9yIj2fz7UU3MFinMrN/4UjjIc+i1QUKUVXMErAll6NhPEFADb
MEtuTCDeusrkIg01MG5s37bJZbZuNuUlaRqn3Vt+x3OjPP68n4Ehsqa6BVRse0sG
JDTxiU06nJ2JfLTZ1xwsW+L3SSd2GQQu/1Og2gaaNYdN6mNCjJXLYdp4ortycjj2
VDALq20xhl67j265nye5a8tgNW1D1a2F/Pn9qtKBE+eDcoN/dK9aj7WAekPuaW45
O8Z4ip7S37gQEZH28ezFbCYU7NdNjihsg6CoUz1cYtdX7rVcoi+7chi1iwWZtOFD
i6omfj2jEoymya1pVpzSaIXr/CBioHM7zFkmn6GR1Io9l4EsG6o2tNF+H5+YNP/+
oCwoVnH9GxqExCtvdRMhsdKTqD3nH6HrhOchSjsk85M6ZqMk7ZcnNXnssBbzVDKW
14LUV7OmBidWx7bB5SoQQG7rKjFN3BwGc6F63A2Q+K0CKimIAAUuchJe2BU9RPmd
btGAyOle7bJrQT8ktA4wMzsqlyXDlZ31Mn6DNWbuFEvEKQ5suu0EzrEWV5Q9ZytJ
TfEbtDZu+gZQGbbAaLr6dzKHA1h29yg22bCOgRg9O6mBI8HS5W1yrlXcyS40TZw9
54Qi+pvP1hyulqz89ZpgoXZuQ9AzlHM6zPjkJbnIQZ/3MQ9wEiLhEvElVF0Kaj3V
TsjM+TKnZ4Rg8rUrwXGoVkp3NUj0U/DOkaADsmZwaSc3nLxaTJwstuDBAw8BEAqO
87S/pesaXP9HO+ZDRr/9rtVGPikZsRXggk1pGoOFnI9jwRRv3uZIZPpNJ3ilWgeM
TvZXASBABZp0IomsClT9vNVXE3T37aMvC/XDVxSK3u2Skb+q2EpFUkqKkSPCvXGS
fmzYtUzE391xHZngYjOoNsj8VNYI0k766TGw2XJk5Qml/u/1KdvjOzJCStHjMVWW
jvVlxm1wUd7RLJbRSJUkoq7jtUygmG9sxJRxC7BdDzoNgqBrOHPi4GDZ27WVLEOM
lIOMTAWqhIXmGx+EIljedX2QiNQiIjFSbmVaM/x6igKOJdzrQrkO68WbzPvtvbeD
xU98L/AmUhTy6vfNDGpEWpvqi60FAgtyN1AxVjA5iRD+GJfomtq/PB1dlI9hX8TF
MY9NqEL+J43s/z/ME8TTUew5eWMSzme9K1sBQ2hhtaYA7t2I+tC6K6qFSDvtZrrR
pIvGveAj0u3pV5YVvh5YUXVR7iT7EFluYmBRRPAMBg/k+MeSRDOjXfq71OMFx8Mg
QnWSwpJMnGES3kDFli+SbVlI/lrhX5I7tKsSdjKrfoI8KtMdaEkLr1L0qr+l7MyR
iYUSMbVfKufkRMkI4+1zuNRPQTl6lf8rteV6LmKmH0WKG//+Rsj9xFrMHZwlGUiP
7bUNq8CPuZVFwM8TN5Vq3Utm5MvHyTbJGa600tEV7+DjDdkkmZ058nhlOrCtN7gF
1iPhYTi/FmjMrw5d24dTNH4QzbnOOfSj/zZzXgzK5P4FtGlkGxEmrHiEFltHCKC5
kSUZ+BbA5DZ9f27ab/mxrDAUJ/e4s0gyd+oEsbAwbu1ipsOGkmDx+g2i6w1OgMyM
llHXCZLiFCtv1Athyri7wjQm2gPZ+wmFR1vDviOtKIznTkj10Xwa4pJ/drqFTG5h
ND1GkJbm/VPfAX0A3VQ8qBvAzes8nT0SNz6pae3tSA2QB4kaXuoZZjdJyyL28Wu8
VBr7OhzDLUBQamwbRT36EM9NJH7d1R4dQe2+wUFpeRUABFgs1s4lZkvgtXlv0+4x
ygWgKI4o83jJzLjNl3VHR3tvFH20C22rvteTtxuyqTeYU2cXzi1dKoRFWn1KLSav
YSv22H8NVrpRS9A2n5GE0ZtY3wzoflzRx6e7asiD9jVCZ8fx3O3v6yVv8jrZQuK5
nFV7PL26yoCVHcbk4Owz9VQZ4605M8Lj5ble3ZdlH/2BwZoM00lS/ZQpmU3Agaj0
2OOud5ViwkVpfkk5/ZwDUmO9XpBh5Xc2p7KXnBAIH3VhcDOt2Jd/BWuPU1ovCrhU
yQ5PC+R6HMPdQ0Et/qGp0hL76Us7hAP51V2uUayrPI9Lwd198tMkzYcPRiWK29GF
Dv168Yw+Nd829mHFecTQeujibce8oHBVEPhqqEQ2RyH3akL8KpsAfSKQKHILIrHu
kgf7430Wt8p4CBE4WfJK1dEK4x8Jx/cfO0qePcgjMR+u8YbPhprnFDM6lmueMvmW
mEibOp76BJM3A0aDa3irc7S0oK/DkKYpz12S9saBgOurWr7GCJHQ36n4XrAQmjwT
nFDaCqZoXcQz0Xt21Q3eEhgN3xR+GFUfKv8clNzn8QQASMABfrGsFxF0ZgfMIfrY
QmimC4PvsxTWfX1u49V6RLbNowUWi7hNVDhQ/YZ4HAdzXlKVOBrYlixHrUGpxmvl
P+EdbS1w7UXiI2NGZI+3EthghTd4qjvES4OpPAFmlo8TP+pBy9DPye3HGfWW6vIe
3Pt/MrS/Cjyfmo59UtwRhnnJeFX2cJ42VYkA+U2/tEjQ7RyrbvUEqnrYNd6wrLF4
RFQbE4jSeuSe0NUW0rn6F2RUJRqi8l8mqxxPmZrbRmc98BGGMC3jG0n3y2i9OEhR
UtUVshx8+qMDG/VDPVYHcHr/b49ZqJwJkOdjogvrJLZA7dYDoQFCuKevQmmJ5a9g
KjbNZrkXXC6Af1hL3Fp1k07Q2gw1bZbxhJNsEFWgM+w9ufncTMK4ooexl3rXgfnl
As81qGjZeO9cTEg8H7ZbrT1Mr45Dlggs1nery4nzQK21vVZ1OUblqyz2znqVE4cz
k7Z1VZNs/9gWz1TQ2UbU4HAfq0NWOdGPaC5LFiqk3FVxqEHyJ0vKy9NLb59RzO7R
FJeGpat30SN3i8W5CmLNHDqa4t9t+oa4RZ1g7WzBjxcr2k0Xm+Ifqp0wql2njTi8
kE51ji/VleVYVIMfaGkBveeXBkEtdq8LcC+45MvCGHwZX52+KN9i5kinKw3OL34k
9ewk81+yFnMXQNVrgbmN7aKYq8getYq576BVRW/JVmwb2MZtQdAUny30/5Zq4yoT
s3pB0TpS9o8kCrUc5+EyPvgQpJ1n6RwYAbN/xLo2J/XmNJgU2FbY7S4KvFCV2UOM
qHFE4wc3C/Kjz6fLizJgSbil+rQ9ib158wclC1Boq3J0VAI40kpAa88gBOI7yfmS
NQ+pERvXyWOOumTH9Q9sU/6EFiyF2OmYXzkTRgM1P9fcq6E/BWEH0gcCgul2WXhZ
z+Yc8VhVibH06X6PbPjiubH1I8y63JA4zvQHiDW1NyIQ8g/Bn0Zy9bGe+GWpUhJO
ip2e+KX7Hkwkew9W2DfyTyRgrAk3m/dmc2ob78Y0VgzZSs6tO2cciF39dplIZDtX
Ve5xktYmQ5M/EmlClx3AyVd107AOvTp7NUCl83777inHy7vKF1QXqIv90BK+b+2W
mEABu5bgY2Abs3+PMrLLgDYVYoMyogIz8C4SSgH4+XBXgKVw32LvXGp6Fz1g4tTQ
6s+oN0xwzv7ZSh7MuYnKifobcFP9yH4T2GmxXAojM9FjdSAV3Bir7MpSKsQKzmWF
yhc0+mQpY56IxntPwvfkbR2iOCcdzxXjA7eBZaUQXSWEvXT4Q6nmrHIciVo892F5
g7wxTK3b0xzb8zascYwxFdIQYxWQUp9D1iqk08GnJN9a+wgqQVYcanscjrSiXNcN
d6TgQXgobiiVVGyBhywi+YneiybS7VpJnRuC4okDMwf0WjSmLjldT89+5YMGUNXP
5GQ1dRGK6LNF7Yo/t7Nw7N8a1OJ9OgKUQkyMzfQl3bdim4hORV1X7R3HVTBrMAk8
FF8uY8HOBwvkJ/9CM3529pACcvxIflb660idBFKyWEiQat9PvIOKhw8Uivfo/LM2
GHi5BnzLDJ4LOZFZJh5pRTjMLcaURVjEgYaK8Gl/I3GTwFsTkasoGyRC2eiMZ1/A
yMVUk41jiJepEzOrLru/FfNaXw7s96wsVfZE9JH8nyFrJTexf0tEwLB6L92H330l
E8f1f1nzRTDZ4T8tgHziVCIjitcsoRh1AQJZFhiY75l/zTtXJIxQF/LgpGP0RUwb
STpgpKTknrGo0JpYvFv+QT4YY9jWMVJ34S0UbC5/OXnRckE+HWAKss4FU6u+4Ph9
Wtvp2m4uyOMRtfEU7ekTdUCYaB7VV/PFrVZgkvobC5JqsVXLTnZWoCluI782VQ+F
DZuqML/UkgECRUGSnvQTzPOWzldc6FezblZQ4LbHliqRBUJXcxsgkXtwMUPfaLAJ
MjgMTSTJ7pTU70qAI9imumYyjm68xl1J2joAKUOF1ypsfQmBKx6w/WrmmtgiEiXr
ffXRZlZBBOCmGV+5iecxRVRNFJJiCKBU/bPaymHxRFhhCj4/yVuUxt1YXjNsVJEW
IIwqSG/DVv4eNxwzdXlztbiJOpnbnhNTpIeru/PxhbtIA2crOTJAX6ZFeOifHK1u
y4KDkoGY3ckRQ1TbE2p03g0yDM5gvekzhRTHbviKNCtUi11RYTo8rnUY5ml0VqNa
1yoKJ2QTACzn+TW1I4qTLJ07+0W8w0thphHwWAKPMH21qpSjOa0hoIugGnkgdvzM
YROAkR7jbm6iRNv9XV8vp+6nQjzVpTMrdnfcArb6zSTMbidxi9+iw7/TXT9zseqT
i21DavdnRqQgIIcEVT+kz33ZSsiKP7Zb4REKzkbzX1w7TMQ5MxUDUMP2aDckoyQi
B+w2L+lVqB9OIMqt7GjIwtg5hQEyChrLNb58mOvzWvsy4aveDUC68n81vYUllOuS
/3lf3kel5CTQ5fWbCbXOnOemskfzfYRyYm8lTmabRdjI2eJHOm15eqGZodiKxf6z
dQMau/DwzLdmLKkZb6e43Y17W8U6vSaRWbPJsqEtK/droA/yHJR5Vg3q4EMdArAz
vYb0k0iJqoBTKnrRlJ3pfIKuotDnyn9WRAWbvMsbzvP8L2e74SvNCFkZ0PPXHqP5
ixIr+Olx25uow5qe/0KrVnqsd29XX/2PLXmItKgyMyFCns9Mc3XM6qVMTAgRBt2T
Ai4CrGWd960LjGZ5NkAguxPiLKSW3Sti8WsOFuHiIAd4etfyXjsI5Fy/SPVlkwR8
053HznlTvc8i0wuPpJTF6j5KwAeQoiy/hpudLUJNThW7WubJLqOn0ge58tpC1Fz2
979pVCLwnwm4+v4rWwPaQX6jvYoaG6n8V9U0y7Bb6jRR3Brlb5KUj8pzwe118U04
1sJDNLkFRTM5ZF+R7BedEx72kBhh2UbfQQ2uvIOILsoa4z0vwiAEjC31kHCvtR+j
UdI8Hc7B5QcA6s3BqmoLsgoB3fmHyi5Zgv41/tvwJwATFRTZxFvxx55rwYgxknyD
UT4iVcHb3h2pNe0fBOgy7dtmKVVKIMLVW/vWOCSkVKLj07l/bnmhcVrmVydwj05k
Ak58yIAQGzYRyQJzYqaZ6y7Qumz5lRMlUf1N3aaN4JLbcHzkH8SOZ7p6PeQQRUQr
36NcXx4O+qsQFTACKeqFdFHPek6CxXCY6cPohx6KXD2DVJvMUeeJV7N+92bH/KNC
ALX7QgxG2qt7twMZlGKrrnBTGNwKN8EXCLMA737P7KFYS08dLXpQhPN/IAqMSuvw
edAE3LaP1CfFzHLj0uaceWZicQpP6jZn6hdj9xa4cRq1nG7JIA2FBcSJcC/dFdK4
gqHBMHlLmCYhPYWb6oH9GddUEJzFGSXX8ElOK07Zd8I6FUykWvyTWOFliarM8j5T
QWkmfjwLAMW8nx5kq27uJ4tT7/n5WBeXJvTw0e17GEK1kvwhqg3xR1tAPmI3pwMU
JlCSmVmy+2GmUX5XZl4NxlS/glbH1a9yyuqVukkJNqldZuJVmv7cTiXICyNQBU55
z0iYaWIdLO8+3Jdbp18v6aWKJgqcCRdCExJe6xFxIwL/If1t0Ldk3uQDZ7rVKDqU
TVvFAWH41pzX/k3aSu3h/Q3cYHdxhUQFl1XRL58lcozpFy7t0QRHCu3z3kUJJbba
NIaAWghWAQHKn4BmamgfGciN42TdDufVmQrrEPrsdstwn2AUt47nDNT2oEgi079T
I6WQagj1Q3cWFU5BQRqQRD9+F8DSDZftJG8PC4Yh2peLLz31BaqyVjA9T7c32dhi
L3u7VhDLn6PcudBCfyuMO5ALx5uXk3ex3Y1KXd34SZRAEt4KSCo3rcAxWUF6BukA
i2fxhy7SUCVffsB2dw6c3b6y02nGvF6eH8n6KR8AuD08a1sawY8U+OhdqV/4FFP6
vRlrfsyrAK4hCz019gQnj4BWnFC8hlekIwcj0Ulpt1H0G9vy9WQF/iACHR0F07l9
n39bcr7hIYLDoUc73twHdVxVHEVaaSpDbmft2moiq1ttcQIaBkOscaj8uXO2aGlk
PYUOtnuNwkumSF3aUTpwexL46389lPaLk22WUubFyIWaxskgDy78MkFi6FOZa4Hz
j/hvDiSI9E4D9S/b+LlIldBGXdZYXG/xLH6sVryu3FiWx3lKb7GuXAI6HINVFaw6
rY2S51dq13NKoXMYqDh2YZ2G3++gEmKvaIa8VHk8vFE/VMrlctJpDTa9pqlibmxZ
HRNs1rCadVHexOmsIGzbF9qKiIIPiNgtElPhPxEDIDwpcrJ4TKcKoexLltSMZ1Gp
AmYVlo8Cr9Ukh05wSFXa1vajGvfOHzanp8hPfzrHr3Zk+KmO+4lwbKoWzWpilsid
+D4me0Qacuy1oMIZ+KgU4L/B6X1dhxC7YWXLs/ervehQsOX8g5CnRa7/flwMKFcU
KdqO7WKaB7g2e/iWj3Lq4iLlsIUOwZ22n/bfLmNQfgLunnJgYE2OdPHN0aXcFkHU
EibMYA3dJHXnXHeTAzmTRHGrjlFiPerQTXB3zwUJm2LXqBljK0QCpvRznsfzZQ3h
axxPRhqc86x68J0uiav7cwJvjc1Ww42/NnMHSlOSZAshHFDseGblUgOiWE+c/FTt
MS6nuD7lG0C+MzXAdAoe9YKP9D1zoy2I30OPl8pbytP2ZxHOFMYcAwIDox1R96sD
7cIusFQtk9PKXnlhQgJPud75IP/+g6Ah2FPtQJdC82/ZQNqlgQV4TmTFvUZEElem
yhaVokCrfexkBbH7nblilcdVnXgNfWtPsIA9EWjLBO/24mljVT98BQyHS8xSGIpk
iBUdcnNKzutVkAFDTeYV6uUdbOmI1RCsUBU+99URouoXT1ZMZ9D7y8gS6ag2ocSP
XcMa4bhtOB2nu8RcuF9ICaFCGpxckWojs8rnWwiqUvo07M0myqSukdJc8RzndJXJ
yO/ka5kT8U4oBy5//WydxE8Z0JIrwEed/LmEF7UzKds84WIYaJdPmRDKm+EdGbEO
80ek6Hs0zJgA40NQfVOHp9KHO8YdkRbrXW7bDw+tfOPtzvgJMRY28d0faVAUS+Sg
S9uPxyAMn1piFaiBo2+Fs9SlHsD1V2WYSraBxdDPbNlhCYuJ2W9h48vEQ/RypKv4
wiNAaOzGaQ+5r9/BwwAE0BNFeH6Q2BLuHDUouUpTNUTqCFgrS4VoBty24ThaVERh
V+k2HJxmUkJ7XjfqfTDTkO3UAG6np2+71JbL4DE4WBpRb0iZlRZsM/Bl0Xkz0Xp0
1UjYSorv20CFoo1uh1NYdZl8/PCrD8JlXgskOqhkvFc2X/wMpG8wxes42KhBxTV8
sJ7hBqOOvfCxvg30bbF0ssxL3h0GpBtRCmg/YhI9HwfktS/kPu8h5LXqJfUpD4AG
um3F3VkLvna7XrOICTunfty3ThuUY11NapHt8hgFg0hrk/AEqXo5l246Dm7kko5L
KhbRsk8RmVsTE96nhVIA4dvn7IvsG52aBBRtkH5hKOqGUOMlwZ0ZyZ6ZuFn8Awub
VQgrND9x7EvWTwsHfCwmxsDkFwXoruJCLj6Yi1nceSAP9apMeEQ8EHq4UD9rTN/t
OqJHSAmmn/OQqeWJOnmHM1ZPxdHN44d8MC6lsdMcM9WTGUKaZWl0Y7LVPn1eN8f6
yHd4c7j73Wy6Z7yRBi7aOudPTZTJY1Dj0NFhIvcuVHD8WIjnoiSEXJN7yrMkwMTz
ky7Qe95X/Jf8tI4h5VLPT1UJHeLcMEe6X9evGCnGFJ7fU7V0KpGlVCw3CwtJaCL7
ZMG9o6mxAWGI6ZU2p5xcm66e9IkrrKA32N7PFjbsM79yEzCh1Hv1WkgpZTCMJRet
w1vmq1MCxA7yeI173zGwDVLD6cSugcB2fvgf9WfQOD9tkDnhQf5mL2SejrIr88Le
Ib4HQx6ms9QaZDc+6cMKgtzL7DI8vaWjR1rja1CuIXO6V3ESUAbrVZ70WrRS80d9
t6RPy6dLqqShXTHzHUpzl1FeWGfZpLi+w4xWhLHfVXCIODHjs6SKlKn6oDAut+v+
qjafF+San4+DEgnivuILIsQmXEBBLqsAyybndh0cUkA1bSQg6rZAl0FIdekJG8ah
bQKCo11G7hEaWmdM7gF8Xj8uxKy/WciPiVrrEIpia9Zt+7ywdEkQx5IX62ko+/RY
w358gf/2Om11CXfhXTpWFvBk19zB8X8Uv3mm9Kdd+XPM9gMEzNECDi+gCA9KNSML
VlS6JGD2u4i4ugUO0MLYHmc2G3l8d1luFSiecAndgb0BnUDlU68GTkv2OrN0bX/p
KC0LuYnevlyxeBaYSvXJWngskvZQK4J1WXn3TOzuFmscO+4zgr1wnvE3Z7OhWjlw
i7xEyOQHnDr0DXGCdJPfyxUP6j2rzoGe8vKHqGcaVjDVtQJKayT1muurkQ19E1JG
PKsSBzFydrFSjl4xHVsP4VnRXMuBGcPpOhSgKWIzWoYwE5udezFgwwNfaHTYDLDd
0szQPIbnMViGN2eoqFLOTlHxlfEYot3m01JA9rsvNHPfwiTs8Id0fN7gAJ2auQ8H
4knmGlq832vYjw8h+yVWVw0wV3w9j7Y1efPFoOmbnznYWN6CY8uQbhia4++8NVQ3
8wvK5l/nq/2MTTszojSRYJf/k4L1kEcW1rIvyXQEoGCwLxjgjoUvNuQcnfkikoU4
YdgXv7Q+AFnquyPy6vQT7ZTIVMRJcvADjaESTWlsJnrvrSWopA8zfc7PT2MSO8E9
JZW0nbHMYRZu3qvSryshq+VxK9ZOaCWmjHwnU0pVJUeKrcfROACEaLRtbwEZ2BWH
+ZWQicmoG8z9g/P14DDHdILBAOcZXK8VG4ERAF3r1CLKkIWCK7d4IwZHGgZlI/aT
tCklw0odewaSw3mKxH/qdL5gKs5WGAX4gyZT/HgZUwU4+rPM4ssjPQqj1kRUfAjY
56qpy4b4vREmKJuykyLPMam3dP/KumS3GE6IfIZknmzHIvl839zJh78eDF+gMveQ
Wm7uDEGUfhN1FWjDW/ZIB5hP2YRJx5EQ+kT2rIzp1nTBxkOaCodkZRRakOPg/+P0
dVNr0/VamXQZupz2SB3Kd0DRGzoeE+4KWeCdXszbgVzjk6Rd0XRZDEsxwM2Z7Kpf
MFIQin4fMX/3pLoq2QTfM+NNIpo13RXsLb9CW6ixxwM7ZjYD5F94HdyjRZyZjdpV
xEsm3LjbE9STU2ZFxL6dgfNogUSopAIa5wHfBbyyCpJCyCGKXzpybFBQ7C4wQlQX
8kbhQX+9b1fwD2OVwsgdwRil050WoOjC+rPIRQAvaISOo1IKup7qCnKhGQ3XYoL6
J5EEJ3fiop6oKBObluz6VTDuZIwDJ7wjoCCxkSm8XiDz+hDUU3PQ0de5ltwp0DE4
ibTiqREtbdc++yCLBwojfWh/+qrhXpEFQlK3QREjuRaWAdTknvS/yLJJ9Hiyp7pT
Gijxl2j1G1XyHwB9sNOLiPb98KnwbsOJxZRyxXutb8ObDhVcAvl5t5fhBl9Fk34/
mwKaMuECvMlQMSK5s+5SJX0USJOPo4w0emAcSE4fUBYYCJLnfLlHQttoKYcgrYRI
e6wd49uZCBWlenDrnZZzWxBirIsiPy+5ui7iQKWFhoGnWXwDb9U7jChs63SMWwhK
UpCr/+FPrCMagQ/P4k0xJNdF/JHCjTucBKT9EmhBrQMAj+iy7LY8mVJEWQMT5Pd7
TsPvcoDPH/98r82MVZlzypLDEm4ZI15URUHTxaii+BdMzCT9pMDpql+IYLK7gRGA
e5Y0SVlKC05jLUnCqXNR4Tv3Uv7Ktx8YBHdyr8FAxp57McncN6kFsGCjyS4YfC9r
14VFhzyX0XeQrIHyxRYsuKjWUAl10aizKSOQWKjisz26/m06dt3SbP8q4k0yfHEm
SaNycQnoUMyURQ39Z152qQsY9ioSIWJwvGd4aRJKZejbfxX8z4KPqtDNcB6UGWQV
MUy+rxmzN+vAZ8ALqspB93sNIp0uY/MhdMu5LC0P06YEQmQyKNGbE7dvbMI85wzu
Dcx6yPSGJUZl5H0KW0Kry0zVn9Vu0uBfkqEREWPbUxZO6RK6fyGVenEAX/PhKgLq
f6IXfnCE39M7sr2jXdg/D20kAynM0hvFG9bnIlNBJu1R6bM9wUZ68aFDW0ZcLSvp
0MjMNibUKUlVmVrbJck5G2k30kuAR9QZWL/f6sZ514CIi/HMfnGghKx3VOQCdIbW
7D2SQ/l6WA9SZ51oKRBs3Pf0bi4Ki9QKsbmQCEUu32nwUC2p/lC/Iw2p6Zjrubjg
rdp2fKyWqT6Is9RsGaEMWwopH1hkEqYm10IYI2ldPuDf/Y7e/yLS7fhami4rRxEB
8T2ugQxMyXq2kWJ3YjuP4hhE7owXg2I3BVFXL/nTXRj5ANnJUliw+JEtHpuhwuB1
vgGkuRhWng6gqVUzx11FyOCJcnuFLNo4tQ/ih15/SflCO3qBL8WUc7t8T+793rFt
nNptw7yrYXUnZVu6sv9uXLZIcA+aEg5c3cW0HzJSQiwQCf3i7c1ul8fpT7vJ8ay2
kIHlCdaKXzngDUFNpk6ZHdrv4c3eShrew7sMV/anZuPey1lni1g1tVGcwA1w0lk1
IQTFC1pnNZpB7yf1/t317wa7uXeyePle/RQmLafs6SY3PhNhGKBCc/RXzXueX3oo
U8S04xuFtONfju+TuuHYi2juNGtfcJe56uteU9Xv+W5UOOH6n8GoMMh6SteI8LZO
CZMLlgUiB+pUuhwLhXqWxKAJ7cdxarnv+fUYBBhu7XNc0eTFrq8RC3kwTG7lCFUj
DYczXB2qkGa8jibR0IQupQYHL+cyR9aVoL2FyFMXK89IrEIAJSgQuXTocY5ZG4HY
zelXDcqWRQ3Kq/7lVYs78eFVaLA+gRphTtDWKGzPmApNJPocQygR1ZY/TwC1OUeH
p4oW+6j/TB9w7QQelJ7Zgkeq6E2xDb4YbKbhLcgy1s+88WEDxG/ynINX3x2JAAGa
9R6EiLRwhViRUZhezhaxIcWVyz7zbEynJj5Rck8AAj2RQxnOFxSyqaahqGDqb/X1
WPzsOZG+aJK5KzmITsMFwFPV+DGpmbZuObMWtm+JURh/f7Nt600K142B9y6AOqS1
pXurmpAfRfjCAyArJKe3alhDCPaehddvD4p9bKHIoCMJVoAI1KsIRvlxdBNil3NA
nbJGxoYJgkJeLvN7DnIO02he/e8JutlxzN6mofnVZSA8pODs/WR9zapRjdVPgTu4
memzJ2B5vNPfrlfqvTPytqBnFJOoSUHUwV7wTKfZX9UaVaaS6pjIhxLcGGtQ9745
CNWPv/F3POmVGg96O3+QkPHZ7C3qFNNYSX1rPsFdJRiOCHMtdoxIGHwZLB5E8dsw
+hcHdGh/PFQssDW68xQLJyjdzicXax3zZs/CUJCke32fWpUskBJKsA8l25Nil49C
vZmkWBlGgQrc70AVN2G58PVsqbpTePS8H6LfRVsQOWYbCglBku1anMPJfcumPrK0
OaMtdKHQOB/BYQo/pH3GNWZx+/0zbv9aT285CAf+kYX7koDb+xxivCe8ED4GBiaO
s4qBPoFiiHFNwKtaZsnvUpi3sm201WM+PFv9hNWprfLY2mhItlLkoyZqiZc4KTWh
gclu11qIZk3Xt+Z+CXSEX4CxF9CJ0CmbltpERMLiJ5+wLMWK/PyszS6kQrPnD1ae
H9vGo+j/Sl1bTpkLWNcEfPtHSmHp1mlesKn8ZgyrtuU37SKzmbRdtC3NxOgyJgmL
4T+qZw5CnZIiDBJzT0cwx5vs9ft606R+/RJQEa5XbOAnIwAHecGzh5v2bpVN3JLt
kFcah6j34Ixb8P8mBcMxFWH9EObMeyzTKGDIE6u+zdqEKRyT6g2u+JC6T2+le6QU
tNXIqD6fiNsS0ERECXRJTIo26XDTUwnixDgu4OjefXZEc9SLoQ7UldJPbRQL5Tnk
BBVnvkedxgnDnXx8403n1BTaLmwn4eN0NEeQzW07+YSArt+ebglWuEsX0x4fmCgD
34aL1huiHoa1HcWCeAHk9fh2BNcs5I16agMmPRLD2mp4uLegV3hIc3iMzMJRyUKh
rLbyNMugwAo7oPEPTE5eEQnvyLl0xi89rHuYUQJsznKnprHk4bWOzjbRhAxaJ8iV
hKEQ5j5fJ2HXeNHQcA5GMtZB5NaI15nuZnHaf/4o/KCrVPXeK1XACbM/4VgHcYur
u9zlEeVGeE62D7VN20W86gZKR7ARGM0i4/oRNUU7Wjpb3cizbjsW/DkiPaLCySuC
r4ez4MSO+h2s0Z3a4c/Nb6V7sXn9eORheoeZGd9DGYsKPHGgCFU9hnnB/CcIEk9Y
wOCl17wz0SMCOLTs1on5EMxwevDeXDZaAbPNxkVx5kGVG0hJkuLdCo7vCVpq92te
ZLtZ1FIgx8geCzAfTPvtxjtYpixecS7tibuZKKrgQfeFDIvTiJYONGCPtMo/PyQp
dF3Vhm/ZTBPDuOv/DHboBQHWL8hWjWAMpFOWgacAl+CEcWDlHRPP1dLpSx8ttoRl
zf/Ogc3VCJ364RXqQOdaIhJd3qWmL3eXj7h5Kkv9P1o3hmlZ5Q3468AH08SHS9lI
/ov66vvqPaPSfN5r+ivRKwGKJ1KrnaQwm4j+StGEr8AvhHm/xiijlZOtd+tPvE9W
APBmOIPWVY+0Cj3SkHYHBnYos2HLEXJU+Y8YZnkp5zAkG95m9OPGYhVJnR8E2/5U
Meyc5auR4nh3CoiQOfABM8Q5FXGoa+ObmJ1XBN8MgDv9UTY1OCuuA+b59rj6I2Wr
dG43Y5r2AP67agO5Xpb6/jOd9du/S0JnzClZIioGPPrFFvFsBN/YxJK1HGlfGYRC
k7Ttgrg7F+Ji559A8I5reMTOJA4P1tqbBo56xqEzDgEJNvFCkY2b8o9TIHEGSWwV
92j8Ye+W1RHWz/ky7YESkVxHmpqU7lV1aOfy59fPzxfmb7MIvcu0ffTRX4A4VMKF
rPzb2ViPEE0c9zpZYe+/cziJ6GRn60nF9UcxpijYKUEpzBHo1x5wlkggR711GX10
KX1fJGb5nwO85vmKPIGI44dWjAbpKVjcBSk7JNJV1yczyXIlWxC3sE2jiPGBASti
bS3Sea5EHvNXdZs+VTP1AE937rG6nBegf+F3/1ZIqHUSK9gPRdA9lislVwhCUwtF
u+bqiRWh1JCEa+bMiGZQmFp5ZlstUPfBKYp5XDV/3q4ysOk70XtD1W8fDsiT0YwQ
GC409PIEIsHSGFARlEH5UvIh4kxvn+WSfIT7mK+Mq+hzItSw7/SF9qfo1ugBfPHK
4bxlfjf9oQ6W+n8v0W6kxggSjiILQjcWYqWWdi5FPw9EEhJHgqLBE8FRw2re5cZE
HGrEzPXuvaMGc1PLp0806oPMRymhCyTgAfa4bP+f7QJovpOu8xh97barTJZSBMdp
SY2/kFgjWd5DXu4fwsASnE9gnO1U8FXLCjjwy7uIQLwDIMjyw6hXm/boRZuIhWi/
qlvF50mJY4el3VD2hwhpa99AVU3V8bXMcjwF+cxIxK/kqpUWvSb22YHNXaOmgbQR
t2FjIzWOm15i2jLfHW6ItVhYMFXW10/CDMYIaXPLF3oUJixYhsMZYVMI+OS870Pv
ALQM60c9HnIRZ7auOrW96/F3u7s3fO0IXvxqXJEyeJxEk7XuJtNz0GJ6NLJwLMy7
JqfBvqYa0TszfuWHcDAZ//Rvl3lX/fy/WhpGOAo2HgEAYs+bmyRMhEFSfsHM7hDF
FN023pQCHXHQ7Uq7cKqQlF9hzS1MJ8/7zoVyDFtJLETRhP6trcNJLzIi1zqRtVib
BiBYrzu/s4edklhmAwMzAPl39rdQFdxJwg1H588M1TGjjFkSKOoltXTdTuDzRvjq
Er1/E8KHhuAhpLq9uYo6ONtsZzJok651DJOZf/SPBIZro9GncHkiGMsUfYE4E2iH
Ktez1ptFoorU8qo+dVhBCEETwO8vJzpA5/ksHGTGaEkHBgoXKPQk/uAEH6gD2hvG
UpV+NTuqUvn/zse2H0gG87ZuZerZSeuM99uVCP6h/0pCKTZfVV+aaUL8YgR2k8P/
WB9rmuySsydxdHmVKwBhPtsJaSh0yZXlGNmppVEv6YUZ1MV2ANJstnBcqy6cel6g
7qqbl/EA+Qd8tUDpn66Z8tFTGfNWFsmdDpiqu/jW3zSRlQ6rFcALGA9XIMMiUi0F
dwctYjLmVam2YD8BBQz7c9xDsULXL2Kf9CyaRD8y38Kn43vuEaJdWz47/I+eLl3k
6CBtsaZTG3hTDq+tA4/1lwSUtG8plFpgdNRxBY5J0FMhgi/oT2YB6U/J008ChoLb
m7TN7DJmzsiM8GjrfN2Q/VrB6kwREJ5/lGXyB1FSOvHrHsBBIewD6KT78quK9z5h
AcXp4uc5SyZNwOFd6BlvwdHcozKciDZXyjgChGySaNCNbXegS2jl2Vdcv73VTpJ3
P3ma3/PDF+AAbJgyGsMxDFBkB3SHSs8MhMr3CbwgAE4F6ls6j0ngAOaiKAMTwBTp
3nIZb4P+6B4E8+VL+XINhxrzyPWHVRb51M2GA5Lwlf4SvFdiLBH6gvl6PNL2hH7N
Pt9asRzFaICIYoaCt3ENfRFJ8hfW+2Vvb8DS/tIcZb4fwvTYspwYJk4/u4H0rx+F
IOBGYR5pKsNxcuu1boIz13sRAmX2vm/PrG9EAcVA/vJMW137XPvWINcFWZPwUd0/
uf7HBmJwRSVjT85KmZYyLnG5pZM4GX++eng76Aa6llHqtNd7L94/itTHYEK/zCT4
ToTiIoLcAIgvlYeUYmttco5LVjd2U5m9tIGpz3M2wxT8M+vWaEqgZVzlgtTkjv1n
rPughBFplHPQRgk7yVGWAbDVzlsV+qyco2HjOpDQkfCvbRZ5BZTecnK0ueV2ogz7
Ekx3uuEDD3o8o9Eu+ydaYu2cHHkrsKjjwZwRhAFs/vLO3D+zm0j3wP6/+m+uyHYI
XuzxSWaMRl7nUuz2SicVjzcMMWdYIcCKUQTHNNV03BNhMcWrSxRfCbsuZ0TcRzyX
mWOtevZEyk46cjEoP7rokhQ7SYjSUoI5LyealxLVR1ZqHnlPgoXa3F2p5I8DQhrN
UuI+JBLELH/L7u9fWqPmX4wToPLBfeTC5Ml8oQiMgmr2qWZ7HO3poS7RRrblk1ph
qBSzH/gZKNAvHRPM9/4veNerkckzzaQcYJ2x9urjUJ6NA5bueFQoC9CwRhb333jr
8m5e5yaylOkdIe9XxOZR1KGGQnIYZDcGNvARLeDImjZjzvuEY2sup50wmgVFwEvt
WsUwzovICt77gNtNrQQfzhZgHSgIUcr/JBlaCgsXXaHbbaGHZ7CZnQCxNpE0Z39G
u6aWE4h/pMCBXKIFpN6dtZfDBkaYKxBYE8qkBlEprPBvvM2KOlJJt2px4Mgo/5mb
r/L1+9WRVFzbalG3OHHYfIJ574wz5uQtgYg58ewIpEd5lYMkl6msx0vjJD+mtLGl
x+k/AlHEJeBRCkXy/eZqRdn8MVUaPCZ8ZmTBBEHiL5g7s4ttMuSkNXoGZRJxrzZJ
scABEJ/WAuHfZeWUgm2iDxnWJjHs56IkqBzizVfCQjZqu7l7ij0diOguv6YzlJBk
ajDcEHIQ7gpYCHmAxCyVbF/m7P8rAftcip0IARKk4qH1i5Owc0tRiV0RU95kXxaM
9D3Av7oFeMtX2/3/IyinmxGBKRsknV6PLwq/I5LFqlJNwHpk7m7IlmWUkSZcCl5a
7y7xSd5Pr35Ms3fkCwj7u31JBQkPzQ4aUtT72niqBRSgp1iWQOWo4dnT5Z4WSW0W
azy28HDCxTFBvKdukpjCph34Xm1Rqm9Z6eygVOXfiOOnGkYddc0W26bi5M02VHq5
+UzV3KET4FZKVhO25oI0olAIVLy1MXifuncghNsvaTFmlIdC55T/F4HlsF2Bdk52
jre9H37dCa+rZM4FaNzrn2vj86fM3meKQfjSekr9E4tSa6sgYyR/CWlc0wR8Fnh7
e8Qxc+c1tevo5N7klzEiJcWdlI71XwX8knTUGStSQeYjv+dNVK27JrcabQMqsnAJ
afnkk1U6eFspSOSEisUSFJlx/kA4aFeJKmIGaeZQ4CyDwaaHpp4CbT667AKcJF/L
Q4VXHlAImAKM6QDY2iwCkCdHrWjH45z667zL/VlUdD+SdHgYrGvZnXbTov5onEYa
IPnfTifbj+Nnluw9e49vo0d3kZQUaYeigk42zr9OJDhVL8v++XNYahpDJzkld97h
b/QwWFBGBXgaWFpe83uOWrHNuGKnFzf74Q6QrmZE3/qMRagkfYg/ah3ZCY++Aj73
6sUaFcbBNyK/Ngtxfnvrx6OptKbti1/j/aW/uy0jEsr8IQ3rla8RbODOK4FMG/rq
uWdMnm1lxZZtCbL6zuJTJ6ymeZ3TShaZEqRrDoknC6vAeB9akl7ScMNDcOEvJpEu
kY/JR1cGJFDiYuRoDFOKWcJVnsb1ITEMIRRC4Pysp6536BKJw+IQiLNZYXIgWYVY
jg+8rIt7B/cQV/nzfbbUB9PBP0t+mM5dVchvaosKvbVvzK+wvpYxLZV1G8DYs8MT
PXCxrlceMJnRWGl+3CiKXD2OCKNrewAVbpAlIAGvPBlddnhpbNucrUtILbqz8iU0
01TYuSl2TO5Al0OA6UxjTPdXuB0Mm8uJfPESwWJsKO1tlpcooZv/jZ7m0mQWIP/r
lvfYca+5vpQfcV+PvNoh4++v3C+erJ10Zlt2FNZsdI/0MTc1/r7HfFKaA8M4idGs
ICLZJEEuYxUxCIPeWm9itlNibX9cc4RquVoDmcamd/R0DHDzKu9uRQrMiQ08H4S1
b2PFm+digcTZGqpO1O3XozqnroyfWIg/ZgCJsx7KudcHsSSkwGJthk5BcJSJEGka
E0QDQQyAZdI2yVdruJIIc5G38C1xh35FMOs67F9mGTOg3ow/PbHTt6VtdtdXlTcr
V+OhhUhh4N06wrF8kbJuZ2fsfea8/vIyqmuNJMK782MS0XDx2GSwNs4GAtRr4Cq6
TpPZTFQ3lU6tyb9DiTgEzoJecAi3Y6/i6Jv1HRD+h2DJ2CwPptj6Tz4RCwWLBbuH
6mcWzEnWPPu5t4Lvkn3xdKkfkkEXwh4nYYH+zlZFtoyl4HJJ01WRBR4sShMNM4dU
fTdPkPWi1ynDXSHhZX8bruusdtjVMW9x0hEAYglfxQYxS0K5N+q5g5FlLA3ybxW4
0LcRc3mMBoj0mNNVFzqNt1dQ0R8UJHIEO81SOzmIjGGbLyRTJoRJFiF+MuUMb3Fx
AaVbV90cvZFOVo9J78q/DWNX9Ni7rOpXZ3ZeaSNzsAUYQ2IU/1zxzCWojovXIjF/
WyIOyxZ0iikQGcSFp1ffRqH+cZUpETXxJ2wiZA9D3TQTcl2oGFJZXCiph9W/BAbM
71mSVUARYhvmlDIQOs16H+vdDYqnI7qq9TPPbekgsNSdYFRJv6o9IZWNiQVvBKb9
b5Qt3dlFHCiTynsD0By97WmhkNL3RavUre1i7gLunOAtZMGDAtDi+J0vqCZ3e/Zo
1kh5hE6Z15zW+lj/IWh6RDpgYPbhFKCrL1zc/u0EHtjUVCe0iLN4+2X0zwwfW6Ng
0dgAC350F7wgEIa2KLd9zO6nOGRtGsfxuO///ohP0ox41sFLCD/C7scazGq1VW8g
YmlhvVzs4pG1tUhyxMCLK+I8aEP1C0go8dpbMDRghKhL/W5m9dw0P0ybNFgbc9D+
Z5QRgztExxdo4DpJ8i/T+/fTytTDNlGUSJFzRWVp3bqtS/t1YrmWZDfKe8qRYKVy
Syojo/SxqnZMP7+GXY6IOee6S912UQxPOTKbeX/iXY7XxKwjpIOupriSLm0D87sD
ne04LYDJFFixBptof9aCULqT2LiGIw4u2Eq8QmztwK1vUuTVK7MPkAzrcuCkLHIk
+rI6gk+vAJDPSrauqRyj9SeB3SDz72vRm9AaZ/jZ5UXjn0UW6AbxKFv7ehLV8+KD
/IfbGcdy1HgqRgeZrNYul2S/Lx9O272VGAqXMiXMHIxZnlkDrnRM5vK2ar4qG0fu
h52a62D2BRWuuEezRZbMiCQh93yb/DMDuWpI52cI8wJBbYUOl75G6DeJBIGfWKE2
xRLBGO1DAImY0JdmGZkCWf0xUUAwKoNRJsh/VnhUy8FSlklQPwe9orNgWoSr6CIU
EeWBTSTSRUuUWaL2W7bVJP6MDYlxFdOkwDBh14uDkRb2jdtUledD+WVBM7JcGl3E
weouRzf5qJTn72DKIB9J6OYXkQifqassvFN+tGdW+pa5vHkm5zCi0UAlHB1dL4Oc
fnHgEn6ET7NknHyGNyhCDAkIdfKCnRggL3HI2WEymdRAlYcgQzHyT9uon7cmBmN8
S9lH33kK/X6TxAy3iN+4180GWmlnrph+xrzZlkcY3HAvE/W4lP6mjvI4HFf/Jd92
G5acKGNHofpBnlue8t5cbmGmFQSZLYd49TF4tTfXduV6EzHy+l17GCHQjEKerchk
WY12zhwxw+NhEhhqnFiBAv5jVVk36eo3Oa0ijVGUiJokRNwlgx8DNWtJ9iu2Tb8+
mqLF2m1dQxJpWYFVXu0ZUl4/+tjlM+aljUzKeOSu7xInLpkzOI20JX1rRpUg3T+Z
r6l5HerbeW2NJSJI8MEZSQ/eUDMnWSQ+bpMbhVLzqYdFGxEGRPUozklGrnrl6Wc+
GbeQyn1kFOJ3pUPygcFyqhxw7j8c6V3P2J7JjJ9VxvHvijV1l8JpJN8nk3mLGPbj
dwvrSCmv2ze/XjFAvzY9kLwqtnF75iXaOvd1CaBPiwClsoCqF+3Z9RUjbASmh7bR
TJSslm5eNVWdV/MR7wljYSfgxjRvtLnyCdjtJHzRZR+aMxNt+i+2mjpy3NSDT5Lm
AgLz9ykmlswAossMY7SQ6u6qJdYltfN+8lsOhRFKpFDgWno82CQ0DIkLuloe82FP
xO7yguJkx+PwvRiOjY8Hqi6U9cCVMoh0cUYq52Uq+goPiqgyyHszDlzrEF8ro4ki
f8RlfHZWbeqFreSNvKAsYunPyclY33LVRTemqwQo6PuF4MBtCchy7UomxQaLGBar
wemmfILv6EA0bvoKU/4ZZvQf2+0UWmfl6wsD9o1dq1dLL7ztxUr32lrvF4pjsOlW
woWO6d41c0yYjXDEdO9R0D4b/dSuziZucS0CyT3+TwKrnrs/RgBa4Akdm82CFuL5
Tq9BB7CcNDr/2xfTPfgINR5ulS3v/HOnSJqwVsRrD1oi/NXlT/aV/ueOGbJCmsHK
3cVjY0JQ7cahFiOr+Kv+35iD9/ZQ9kefb3Cz9RjMoROUUVNQYuNYGlQE0rxgvJX+
vBNLWPpcBdW4VkJqtGpeilcZZ+46ZI2ii8rjrXoRDH5C2F0RPjfLkD5UOVNhB1p6

`pragma protect end_protected
