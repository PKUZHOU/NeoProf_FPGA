// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
LRjZqN08aRtLNLBfxHQnOGApjcD4i11qXVNLdvvo/NCnspqz+ouwiRYzIeWX
9GCrlsKM+Qrt8kcvsEnm0RvhvJQ2ObSU0j7o/oMZ97/IjBhRrUqbQMDeKvn9
hqtpij2IB2vFDzDxARDX1CIdgMYvOzupphaf2wOhEPg0xbESfuO3RjvDPbw/
6MPt2Kf+DPFCw7qEaM1G9E0YKm+5GF/re9xnA93QvLDo1fXX+mIoOSuz4QTA
WqtylEfbWfuIooPurMG8Hy67TnNk+GJWDK8475xq1eRQTNRHf1pVpVhIEDX/
/OBcqhiLS1AzWs0S6G+BO/s2thw9YVdAU7d2CVl6ew==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
X1Lh/k/GLDIFTBlSlQYbLrmmC+o5lUCAQaUG9zect9i+PKW1ToDeVjWItHwp
T3WqLUlw8nBqIOosL23AmPkffnam2CFow4AcjVrE3OsWYOqCQ5cQUTqGCq3z
0Zw5LRzh0HhvMwHMLEAt1IljqaKI907Sd30hlPx7C2sibFSp3A4x7x/QzN2x
ECoUGVhDZQ9jYmnmsgcjQ1XwD8wt/b9h4Yij7rmOkqh3J5KTxtjWx6BmiPyb
88AFArfMnByxO4nmpF/i8BkWFmHkdSATjhvhTwJazjDMPSh2LfRjVT+ZIIWi
7GrwToX+hW9QTyd2iZCWNa194+YT/2PfUANX3My/og==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
m1H0XI6DUJsMTvM8bPE4zdSZ6qGqmojY4usCia6f3kM1PL4IIiLZtOF90Lrg
5nsCCn+zbsXiZd28eUOV7gKSQlP4d2sLMKTpzRpLYgb4DVGCIta8DHxHtvAn
2TOe0hKcabSsPGEbJEpa43I7Zyg7xGW4MzKscDLJDN4neL7/yqolzHLqMZBq
7b/iM+XyRyjcrJaUmDBmet+4vUNYyo5X/f1jDvsQDqGIHa2ICSXgljqd+ScO
d88ywQJbDz+tsFd4y7p3A/DMBlAOsLpDYM72NeG5s3JY8TTPK74pce5Q/O1X
cSSLKwG7kLUiWVeKWHzQ+JgGCKHeNb8coRMpAL37Nw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
eU5+hC9c/xHWyu//aSjrf10K4HyEXKFV23Yz6gCGQ1pDPvfK7SbvWrXc+4uV
ymuGAOokp6WCiuvLtCwSvWTchlIVmBHLhwsXS0RGoqpXcS1sjwr0gNqPYcsc
271XkKnhW3AOQm8J3CZGiuEkqiFPu/PTyXfUdv8/AtDrbKFQAok=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Tq2FP69yeusaoWCCissqsIjB4zBB9eys3yS+SevfhjjXISCzwmLXA/msCgB7
VdQW22scyWu7nNSOF5TSm8JvJIfsx4z0lxG8oDq1J3WivxSkUY5uyMajXubA
TKq2a3xge6Ah8yMBhWsHpvE/K3niKbPsUyweKfNCZEmUCWHj0LssPoi5GA2j
Vttdj9sBOIhizwGHJFYxKUmKaSu69Wf6G3m2Mjmj3JrfvzmuhspOVRdDXQR/
TwwAV9SfBlFIlt4rREukXNBdolFd2O9R+MQaE2UnAtenvfKkxuNhrHaTfXQ8
SzzdQIfbtWOyFD8kQVMvF7cQqoV8Nwwrnbtn7DFuQT5wzwT8dxbMKDRT1VqX
y7FQRUbRJvb52Kfng+UOPE4t6lZ4Wf8sBAgsq8hLYrCDHylOMcTJDwXh9sEW
YOvaxyHsqzkqKwSbBfvPCOzSXN+l/x/e8ArkRCqHNDloHZP52wXYbuAm1kIZ
l5EIvigSlDV7wBK+J6nsWB87uuoR5a//


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
fXlmmRjoUWoC+oWqwPXPxQ8U2l2v8zpzXqsIdsBNReegwW5SjSI99wR9WCEh
4mO4Jbhocmp4q8/wsJslADm0p7H3fH5R1DEq7Ppw4nKoYMHrvm3mlXE5xNjL
+W0PPZr3+Kb7Bsmy0ZS9Rhkm4/cMyZopv6/Q/oMxBv3nSdOvItI=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
b//2SaAVMrANasHTY2hE11NkqyruoDHEe1/PNdu6fRrFUjoCXTxHupiGwBPY
g0mukT6Ff/Ktte9UJFA1VukkkX1lYYfSrjrkDSLmhlng/lQ48GzjoaCleU+O
VqXj7yDt43l1eSBknAQ8RdwA+DcpbMFpJlheNALF+p5A5VhoDOY=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 10112)
`pragma protect data_block
oZoGuLCfy2Du8PpT/H8Rdm/ulsoQkA0yO0AJ+rkXQJc8hY4fZ0yR1chNIcgD
mczuImbulF/w2P/WW8XKkae2eRrHPXWx8APxkN2DfAMHmfoZh9XgUMuHQT5/
7XM52REyfMWSv9ePGE23589uZ+2e161Z5AZ6Hp7442nnwEmv0GfACK9CEz8I
3KUqw8V1b+H/8sRGETZbW6dkSrIQq6RUvhSD4zgnj9fpNIskgFUcb4/t5E5q
4nGvnU8jEhmDI/+7XXf3AsJT1ltz2iM1oT1JV8WVeygr4t+OcOkbCVkGL1pr
WPWnhCysezECpy9nMTfNdWAqK9wvEEFN+22JS5xJcjV7r+6njiwHTD0S2XO/
NhQ2ELE7okFvscMspeE3bO5mGtHZ/cb8t141s4ObCpuntMKA5sucXNBchQG/
MYlN4k2buI/zqkFNb3rzJu7Ka/KjTEERKNo/ftn4914NCMHtc05hy7mTu0wL
obETS1r6sdpW+GIkxXppK8EtHkl3IrarUsjG72PnjyV+4zGIIiGa3DKPHTpX
ASpoTh4hVSN63SQUvm7mSHYH3Z8ROa0FqQaEyfDPkmeZmz4s7fsXmTy1Rf79
CN57vn9HOX72GTSPg7eJ3lFhZISzS7OUJy7Okt7aKdDOVk7T4o3w07w153SD
TcnI+Cl6EAw9IAQv6KnLy0cdVhVU/rDO+yj/phplJrQWrPvkq2qwhPgln0Qs
rFOlf2wYN4hcmCHje1IXzXobV2gTOt2Suuc9dg/Mvip/T3KAmrl4x04SKiqy
jXaXXOfiKdNZyIz1mWpGTyXWD5J81yamf5pz/XjOQOcGRsTVp25c6SZ5G5Hb
yqGm6GYJCN5ND/IQUgAdhmClakPFj6c0KGRg2wTY4iweaTFhBqyQzUBp3IwX
mNTskOwWpmJkYcu76mrNNPfVpeOk1G63r1Ma4ybh57cTQxt2k8I21Oc3+sFe
xYVkCUq5/SYCakqwTudQu6OgqKtwy5oVyjHhpveO7natM9ED+Z2XVRdHpnVd
0rq2Ppkuu+UXZlgHOJlD1jVWYzK36Pn3Tba/3kJsoU8IuumLnKbP3o0PXexI
cP5TToHjYRDPHV4IbVwt4N1KlOXhbWCpX1nQtnQAfmcxqaU5xLjxzWOhSbiw
AF9T1pOA5BdZQD9MsPigpi0SrJSb3QSLnncrbydxSW+T0GNRGQyRvYohqiPH
kuOzjauw5KXZ0MwWSpbBfwhLwFQZ7UP9nl/10FqO4K9tHfiUrWNGlXTVg4lC
z1hl65vm1XowCvzX0oGQjHbKxAQrYSsCQ5XH6W4wBfcz2OWYsCIT2WYcYJoP
QPCUbk7JzwIs0l/nz/1mLnv6VHM7eri1x7UNsMvAplhcQ369FCGrFx3JUAh3
K5UNAgoaBamea23nPchrHtQh3Ms2W9QPPbUskqJde8yJ+YH2sEZ4RPEanAdU
c/NtROJp56L6Z0XIOQifJ08LMoAvSkim5C+7UotK7Zt267BxC4UewIDJXsvi
MgOMC6bpwm7TqP8ODbxQsKpDqEM/ZFjjbKjE0bK/viA48A9ZtpvXBwXgP1aA
34Oww10nu3Ma4HzoHGGkDzffQTGYEPql4kPhp62MWzvUfgL0TmCuAIXPXC3Y
spHmFzIoOjAUOG9qd1ihGHpeikBq86XniOVTv2vrKliNiFB5EUDw7b1XLeVb
QX0A9USX+jfqAf0yMu006XhbTFSNb3IipNicQ9APn/Sp4G1BpFJKb3+H225A
DxdbVe5GC7XKw5IW75/zntF9/BJOXWtThOJ3LngtKyMLE5uFyrusFahDzFxo
KRHrbkkZj4kfGVWk7J3KYJfLiE1aIe1O4yB1jlEZF1LB0080hsQbgeS6thji
9YN8yv8fgk404RCouMNyvDOtYD004hODan75qefA+PmaPCrtqLdgrufcOz74
1MMoZHpuvjeGzT2ROjTclanWdDYCYnO3nU/25HAAPRdo9J/A4ISEfPrCKm78
ecAjotDPuSan33hwyWbb/d8+nZRQOpKJ9qdgdBJNz0Cz0Tyb28LrnteoXljk
3Nlqj2xz4JtvXrQTNqIZJrnx3kl/mz2RpMuMmSmYU5QT35hJnpAg6Yt0VCb9
23YhhxgKiHADi8hJg2wsb0CbR7wEnL93S6Mm58tWT+Uyswg1FTIGineUYww1
QBJ2yfgQdACLXOIajQG2hJaNnjssUd0ORKgdT9gm3QY9fWLIqmwHFS1L2/fI
WV9pS4IHi4v3FY3yXYLgUDfaxAPkCnPvIM/8YugMg2y1S22DNkwiwsfFY91D
7+2f3pqn4X7SpbVdqRewKn/HW+v1PxCV7vwOsMi8AcQeAh20Mh5vdcyG1Cjf
Usb3Nwfb/jcUIs020Sv+XrN0xX2wyZbJDEOuzos2/Wwo3JonBPDQS0Sfncg8
vB5zqjLLgE3qCW+9mkNhsL84km9orMlUvugoMIje/4Q9NYWmVPwCy/JLZxLf
TR8PuF48C6vAzQIa1VgYSQoIZc1aqgbpajVI4Klo45Fyz2IWUluQfSoTXTRW
XJHCkVLf3Em7idew8hUNzTro6SIfxWABnsv3AbSb4WurGvOhHigcbDLAmxQY
q8MU2O1QIGmh0QK3H+GAZ7wlFXEp6YJmXH5yt0QGobIJpabQXGOTYWt93Zd7
xaB1Eh1sGhVIA3d8IHq8tyMcmEL1c6iDHd0/TrzbhlSlAvs/LoMX9H8mL68m
in1bt5bLwHuadUFIe4CkZpBsj8yxhZVMnlQ+QNoGUGRKflgFI3ngZXiRsW/3
ZKVZA9XrJdNF4rVlG4iUCmblEDmJf8tr6ewDEmOC9c+eKoZHle8GeCd//l1+
Sw2gqdJXMiDICh7+aWhqqCillIsS4lOvc1dmOuInEqlxap06+8nagfY5nGNw
teoxBvHWGM154xMTIj+R/W9nTNKiw4w5zkyRwCe5cMPVHmu53ue87clcmE+W
+P7qDqncBeUUJd1hLuNrKOfCKsZgFmZ7TsKK9DEkfHsrxrctssVRLU8FMjn6
qMaJRS7Tt49BCTTcKq8qlntblNlZl7AlkN3a+tYLtieMtWibNf5ag/L8hGWu
sE+Ld9aDYwsu6VEjxEW0FQz26may//9zGSYWSgvi+HGb77OI2lgtgSg76Pyf
wZMJnG1R7/6D46R2VNV0q3j1takQ+Dv1j/u88UpxK/OQptqT6PvTo5Q091rE
vRoluEJm4MPXp6Q0dxFq/Ux8kU9om3g9HFqGa3ABNtJoojOaoDLEaWS0o/J1
awca9FE8qvV8YqNRkRq7ySUz8JIHEvztRIvMij0AH7CIe7m3CIZj0nt4d1z3
tOE5E6/bk4MjnxZv5XpzIp3uJ+mrOStctFW3mv6/GuqAhuKW7atPoJ+mjxGU
fbCMfnlP4Gy4DtPJrkLuI19uII7CCtmsyFYktf2VD3HzaOS7cTJL7xDupxES
hpsEBxConXKWrfIAabvsjULaA/D9wmaimvcwoezWBlJOpnbNQHLd5X/3p369
iYQ3xwD36v9SQY1ykZkrAgFtHABQPXXARgNjBn55fmOKbjq+dmwfN9hS5UME
HnRecoDKl/JOw/t4WQ8wyJ5acFQlv+SBolrO9ZHf9BlESllAOIDbPB8fK411
+DE92vSzwlSLPWh1D4/1yGAErcpNYa/VA8Mv8kURmgzw6AEgiY8aVh4Q0ree
zaRbPOpr9lrt452WInM8v3UbggP0h3R/BTk9WWvoEPBT81QF3ztYANMZSZFh
DXxT0HyqqXHgEJtO+I1mmOMECDmJEfZkpj5RFDNPV1edh4zgvNSUjOgWSHFZ
wyuVvSLq6GO0tFAlUBA6NkDBL8jKzeUWrPv0LQi3Ys2Cr43fiZf537tjBhj6
besALOzzMLU58IHAVXKNGvqc9TJ+cmPLhhdNT4ZgYpwfRBINE1U5ZUYzj9/C
EIWCCodudOzxslJFB9UcjQtPOXUyVXwIbtL1ttS0pBhyWoYh4k6eIbzWZDjo
7y4zHy51hmF07VdBzcHhQH5CRvqk9j3lqxjzXuwGtvC0dwYVnrrFfn3tHKVu
dbYleE93eozbb33rP91SlOHhG1Io7g+UQdJcgZXNl1ftQ1e4Pb7MezfJaQwn
w32A70/2alP3IJpWfsd01/FT2+Rc8iF0GjVo41xH2M6z80WFPrNgrrFLcX0Y
mnJOClyIS3j/ETj0ZK3/ikRx+ROcYKANOEXAkmhP5Lzd8cWXgEatVifQsU2d
mZUhbG0GY6jiEj/6Tvb2BRFy79jt/0sjwqSsB1b3vPiZDQzJc6x1qbaT01Rx
bWYef3M03qhGCIYbc2/EhVIK1321EsxyCPOe5p/UdVspec7sRQnP5fSodXgY
XNuvT7MVkcmvmEc2IWwZf/9sfrVCeXUoemXyoU3IL66fsfYTYTXaHCYf14YS
D0gOcl6c+nSncGKcv6rDo9JNSQXxlee2DO0QvsLmIzpL1am/vbeYHM46HXYj
7TPIGJTx2RSWgBsBQ5drJiBZ7CzrOLyhDyG7MZXJhNvzWaWn8WKd7/mwX/6v
4/1zZ0JaFJ0tHfLVq6ynMz56MaGDuAzNSAi9qMxKIAgPCtKTmh1r/EXd2PF9
WWWrqV2i0X2nIeIgsGGVl1Z2Kie4NtiQ6n2hOZJCUeFALZSC5kpadzoKkCpm
umfn9RriNeJjTiid90x7pLylV9Ew4KRQe3vvhRvcWLsWLe+ejrGm3dpOqZ8+
1xPcNyQ04Q3z6OowAktr74UtuCua9bB1LDf8h0xCaDRqraEHqNakXtPNtoWB
W60+JaawZs6+ccd4FUh4SmgzsWQoz2p6XNZURBUQ9ZJtXrxyRLX2x5IWraNM
BGLnMXqZpz/+kSebNA9Vcc25hiW9xciquY/XbW8ZbcCpc8eK8C9hQAXDWihX
fnIZiNe/3woZaqar9emg2/0VXDywi297NE3i99a+jKi4mOMeWeT2XzSmpoTb
eIXsdgepKnNBN4ymKqGyAn/joUhXl2PEAZLAvac95vMo4R0xM8hUNgcCRXrJ
5Plk+5q1vnhipHPztgtr5eM7XrP1QB9pbTSg01boMTx/gWqFqVwxahA2A5Ng
pSgNRJkjHasNVCVynXsmYKGDJeHEpAMjE9Z7Pkz9dsO24nKIdHW+lK4Baxrl
AnWS191xoMKeYenj8BVy04QTdRjbuC4ibkshBxFeTJmNxm5T6VKzbRz4nX2C
GIlI6kNo3/HNIJPiG54bXudMcM/kWGQUUmDoAEintnH4RbpxoySnudhQ4JtH
fpKPe0tg/OOVoSczXxJ+Lv8WrWvXid2R9i66XCj1OQgtRF5QJaKhhxUJIQj0
vimoqIT6/bk40h4Mi53kZetIT3sc9/FGyDwJARTRuglaCTjcFK+K8xMii5HX
kZPw+q7jopVqC+EQc+18lDgzGRxRZucdFjcGBOeSVqu2ai0lwJtqUarG2WJX
dfJlp5g3OEdBo3i89F8LhQwqolczd2u3uD4I9Qcawvg2v2Dia/SqcZVplimD
/BdCvly8B9ifpf3HlINCwXfCwsBvAOzvDgWspvkCYMmX2C7Eniad3RD18zA1
fiXaoNznpJ/xsbt/3PlUUlNCgRyCt183IQb+tTvOq6lx53r8MmRgUVyqv/ZI
utB6onU6vfVdJLK1TE7WeCRrVME2oLI7qiT1qxRfuiDwEjEdhRf+Uxxnzypo
rLeqq/LYW2+lVe2hlcX4aQmwEZywxg2MmZpPj3gX1zLX4MJ9Ry/rMvcbyhxN
j3BR6jOjfDde/Sf/KMmJwCk0pFntUQ+uayouUT65+Bgmay0rVmb4KoOsT8nA
qbO76K3sbmANYEDDkfwry5sC7SVEFwAgJLV2PNskYPtJL+fe/4VEBsjuBbtq
1FUEFKkcoGxG95Kyv4B0PugGTfZT2zt3Y/s9Es1uB0r3BgY9Pxt/ph0T5EqL
IZqw9vyQvjTyKLfF79zq222crPXdzxXJiltvg1rE3gwbvHmPKvg7VtuqzHqU
pwa24Dq1228g6EFnbCsQWYljfCnHlM0W54jpcgCwpIZge+Jqh9Sj2BaR9V9S
a8q2zkAS+OwWQ/6C4GQIv4ZBdUS1mXY667vwmlOqpkApGgwC668Ii9Fl36TZ
Z39ZuQwkx09ccP7K7sbr7m6mXKoxzPfLXTZojSMR0DWG0/5VRCUly1QN1xGz
0opWTLeYxz9iCbh/FjIrbuQBG5PhEUBMPYB+Q+voXfo3jA3iQQ7x7VBbGiMl
gq1pJ8QuuqkO7ABlI0nGTt53PuksYPayTs13kryNxyqkkNHRs6D0NHrFtQf9
jBd0dSQoSBdb34KFFNZj1HuscN/iPY6O5Gls94rGqZZ+mv+WCF4uhnFLeXNO
XmGYhtAvp+q08U5JB+whrySl7CPYA/g7zzwCgW4B3gnjHvfa8sALFHml+5lh
qIbWT6R85Dg1lGUlKk3Kk519PvM77KbOG8jV3lU7RlZsIKWfOrPJwUcp0YP2
VrlvJKAuN1RCDTsjce62IfIKjz4FvHCg+AwIbQLkfq5UZ+st6aLDq7viPSat
f8Sel3egJ9vneAUXTXBv4+d2g01s/scIy1VkOuBK3uQtegWI8Bw2V83vhBWA
YW8oIaTkXwZzcmfOa4c7Vi1XBJBOibyRJRxh4AfaCtkWVAnLJRwkgiG53yR1
wHPfpBGXYlsZdV7X+XQOJ7iYgM1hyGG1JsNamkOqlouIGItR6t1QeCwtCwwa
pzFVmAbrANhDWivbVzI2R6+sz6s03H+ckmdlLu898hyAl1DccTqm2hyY9gl5
5EI+uy6c4LFE21C7Y9+4R6nbt56daZ72nJhmJWZWYy7UzrFsIJvzZ3/4of8B
hijA8+iJ3wDa/RYdQQ8/fltWI3EnL0rlQJeCKVPH96FWVDMimnVIX1vk2X39
JcSNX3gTPpwfcRIcnxtE3C2D1uHGewShpEYmsDyulyVVRLmWRKgtAPUp12Wm
F5F/+IPn7pLvWZDbcvnmnf3XT1Tjc8PuyUNs9+PwNbmKvHFEaY8EGv6U5pYE
gu3al/cGWfUkUAfuBN7NJ4QXy/DHlVOvpNaqTTztzxFFttJHaUOZjATBl4ZL
44IVc1/IxDZgWG9+s+OVsBZY835YheUY3Gemb9vSFB9/ioyFZwXniS7ufojF
YfcvRXrHlruiKCiqjqpGj3TanZ4bwSWluw6uVgZU8e0tU5K6PPB/Io+1m+Pt
rIdazCIiZLKaX6haSgiMmGw9/SGPB0dVJVym1apGpFt1lIrmosPVpOSckfrO
bh3YlRg9fseMKS5G/LDJQxkswqtygBtSNhiM2SVrMguueLVtRgf1Z+MJYPxr
nVhg85SJMPclojaYZ/p8F2DdV+eM3bQlSZGqFH086aUfuauG09FKD7NOaEIz
i/vTH649CFHXSU9R7EqyEqZC8hlo6a72GwqgsJ6uwKpOy3wc2Bnc3cu6B7tv
0p65ytqRxZUzAsrDE2ET1+aRWf2lc2nZbYVckWF4pj9ptBRta5XvRlUpTurN
4eV0DzUuBla0zybmMLpSj+lpuXxoSs2xePToQRsqOj/ZPoMCJ4j8RNXh7MqZ
FlG1aWlQatMnUk8ZLh9LeN+0HnlfOy9t9mig9oj2TOtQ7dxIVx0dnPAkDhl0
Pwj+b6cAGOQ/Cfz0SbayfvikTIGo/o3Eua+mUoxFg+YRhpFOmYCxuNZhVKJg
fSr64lWJBfbPK/hNtT/GWdTDPjc9ulkAFmuGT4unl8JYvzCcUrxT4eMJ8f0V
qlLz5DVrFr4JNEPk42cvHnDsdk+1E1obad16Jq+dj0Q6etFPrWKaQcZGyzmD
H4Q4zFzjkDELhejI6Q3bmhv2bSEBjj53rrUCc3xiUkv2pjvAA7qcaQ0Stbz0
WQA+rT4Z3ogb3cO6rH+j1s2g6u3ZKbrMMLZvydgpSk1KpmtpYBbawEh5cW6p
fXURkQz/EkE6oykcr401d12AtGgBU7k+1CBcKByKRejmAPsTToFSqxl5uC8d
FI7/CljsvtInJ8hFl5fB3Dott4FbLvyMHYtpa/35xUutq3VIjdPNaDDevTXA
HQ6cQDhllAXYOMmTBRYVTmVrcnHLFRu1+5Rer5F5Nd9Bx7j83e9jkbWSTTEd
rGO8mvdoGiy0z6QOtHmAW9u8eIG/5bxK3aVW1ZHrxj4Zze3FsBDtt6cmrS8W
pzOQV4LeAFHLXl1+Pv18uvZnMDEhQTm6oFrVOy6Y3YYVtZIZoaJ5YsirdyI8
FsO8cK5+vn+gF4ENUdAe+aB+DJAcEXK0UBuPJDUwePRnboQPeBVVdW67WuBZ
NfQf2BgnZKhWp2AkbDAh8s/9ldhkXb4B0jwY1hNMewRBBeVffxE6EmQW+2Sg
9s0l/DEY7IMRdwMcB8Ni/xwG7s8HdYvAMP6fjQ16Cmro9eq5e3gIDWitmO/q
ZEMgpQVpSIV1BKyuZm1vm8fRvcXmjD678sPv54azN2n6+O9eb0t7OKF5rWvY
oEu1lV/kL/SqtatPkfuzre0fW76S959gHxnaVh/g9CQ84du7wqL0cxcgYy5H
mc4/tJXGJwT4l3m5TIbNVeRBmmDr/bCQY9OuJJSbR4Cf00wV3zN6/uy+94Rx
jDnDj0jQn+4PgtbgBAypHBgiB2wgKgZxtjIDCH4rYuaRAxy1Yv4rFHE5MFgb
cNNdLE5rzjBZZa6QeV6FEvhMWkJxfJiVaJzcc8Hv8XJK8AUzCUbsgZ5LAd4Q
Cof9fkNo1CW7j/v66me04wJPJf9VH3kaOiiZjOtQ+i2QfcsKB4yQECdLpFei
F1S06b4PxXXBXUIvuWqNqQL9ERWIqOTKqdcS3+R4pTAF9zquU0oWEbuHaZ1S
xRFTiJyQin+cslaZGLUeDXUh8f/qOLhySKEkU7TB3XDwB60JMrcJmssWEyle
vu3jLcUJIwhF+mp0pFO5iPf29BFm7fW85KdSY6QS4moi/NlJLcHpl9tEFXpP
y6c5xRnoT9QKpk6PcMJ8g1opqxnOkrWnX4w7U/2FcQhldEGJ89/iK0yw0IFM
ZrZbiA7yk/J3ox41OxEJ/3G4zpnbrYYNj5V2SB0jF7686lAtrn/3hxL0jBih
aPKdrutG2ykMDKc6/qQ9XufDBzGJN3jEBW3f+/DS14ojNx3nmkEyfe60kskw
gWiDd/O7VyYu1JxEWNiLJIL53MU9aEc5RJNpnqaZmKSQPWT9Cy0TwxdIiLTG
RKnmfyLcUpbh5zojnW9q2JBO9563E5rezwjko7nup4NnXEVjc/EhDbuoiUcL
N5yhrY/yOmxjA7i7ji52TI40boi0RIcWK/iE0ymi4kadg33a45AR7wgyXvKx
QJtvRFkL1xcvkw5tiXYEmvCEBV/z5R0XU40klFSuY7zDuBpBP6gdnjD7/S3N
SfG3KYhUp7VvQwev55h/y8n5VbPFLNoBbmFFvdR0O+Jz566/KQwfP4XTRuo1
H9wvS0dTzlHudLmeRPgFmlhuB6qj3KeinOGiNGUf93rPrUW8/Yz8ufMfLbPX
BEn0lZTHmPVfDnmV/tUPJWrZIU9hZ0J6Mm5Ktwk6slxAXwa/Fo+IgsoWeYxc
pemQ6BdhyKnN62qX3PPYd5kav78SdcxMvh/Gi36pqKy5LyXC/vVm8lnOnUWd
/0dMAGnglnpdt1ke7f9CjQuzT96Q+711Nngz//JAQU4NwV/pEaJ+MSME9prS
D5vLW+EhdUaUDyXrokURbndNFyykUfdimV6A+FZf5hVjx4/ylOllDNvZGD9M
WTobx/GXd/QGumZxoBSvpx0aosyMzwJZRNyi0xIdmswbtyJz0fTlw/IvMt+E
codd956r4fVUwRDa+EEiOg48S0jx2DcQfpotZLA3B8tawLXb/30mGcfmTOd2
abqUJiDtp3/IuGwRwKeUNYNE03ludgVtnBYKAvzk/XaQy16Kg26shv7pLyBc
+267LKn0IOz42LfUMDtoxBHUy371wlHi82ER4RXehjnwI10kDjly1yuoYx3A
MC59wi1LxTaBW0WWjcfNleHFEH9moSGjqVInkG1z1B1MLdChyzfMPqkj9fSZ
EGp4Ggft7O9gUNCJ1ay5OGJ7fpoO2oLaqF7/74wlmUSz1OKCSJ/30pY5J8hm
dxDOM32va87kqlzuBqMGMdwwKl99C5qROlTZFRP4RshoYO0TKC6TaWgeao6W
ppKIpRWPLE8cbaJCFmRjW7RUaI6Dj+xsRU4AZu/sQym4CZj2RKEXft5AO8Ve
i+BKfho2nT0JPkSD9Iin/QiAQuMtBP3cJcNXUbNmnk3x2pT7K5OyxMBBeYOa
i2ygncQm8XmuevSenhrivKJjtrGR/XsflO/Yax2ciBdpxy4FmM3pCP9RuppV
ylFvYh3ZKNjBImBbAYkfnUvX4XuDvcjz5WV29UwH2AVdHzGF9LKpOz+nUduU
DV9Ih+2rweFxGufMEz5S192bcZeTm0inuDaEuv5URkJQgJyvWpmOq+NGb/xT
tFBVdbRdpUB5vceBPSJLKSLx7Qz+N6h/zCLVpcUbubWtGdH2HYU/FepFrMcF
Ipp3gqhTOZKcJ16Zj9Pv8bLCCGveAQxn0/5kl3Fuiou0GUEl9SsBxDsdJEDP
tFZ0ivy0EU8HpTWxvHvSB8mshgjPK6mBfHRrywBbu5Cux1/yOQi2UAL3WKjY
n0czxWQ8gpoZUrj2kkZFnQaa5cEypVJk2M46lLFzMV+jn1JPhw/pVGekbjhq
cv/Rvukdibse6JrjVcG/35ZS0Ggyy4F7W88TZcY9aU3Bg0q9gFizWWPZywvE
vLPbV4+EqrMgCmLaXqVO9R1cnug8DO7MBFANluqQ/YTc9Ct1R3D6GWXN0c81
uTnX2++5niAOxtYWhzprRV5xtrfd1TL6WLZ44kL34vNvM7w8XEHd7V7OFIWU
m9yKdD/ny6fc7PlvKmxhoA3yFQ/m/eCFxuX70fibUOe+sEZ+EeS3GrgHW5eF
lHvmGJLEHRxRDdGWKAQgo7QvYwEF8eAKk83liqQRBgFvggAtUc0zVnlJiyo4
61/YkjfNcBWUcy/Z6lxFr1eqpLVsaGXrpaPHc7aXdlEFnCWnjLaTetXeTtrG
c/k8N2pfMjINxfLLFJPPKH8T7u5ZCcWXnjelbMpyvA5wYF7m4vGcjuKUS/vJ
QUeVd8R4O+BSU/u1zJElh4uS1c9x0RPY6RbokHOy25HEZvq98yNEKPlXE+XN
HNT/bUD6ZInU5Q6jdT3rUEHX++sVKC1990r6bw+l39Q8Fz0yEMkTYvpjUMNT
ycEHi+h/RamXEBuUT8rziqcklMcTNMM9aTidIp0/8ayA37CD9f7b+vEv/+Fq
UaONcPZJUJYrgPxTEpsBFKWqdj1oUbcgLl3PJDEFUS4psU7SOj7YU4V95wW+
ZDbN4QQLS1/qqx8OYQWTCXcpWYubekbBhRq8KfFKo7v+ugI2eOmeZmX6/h6G
asl+Fgz28ptVSrM8G74pEwBdWNtiF+f/E/oncGHi1lPgOJQeS/PWn2KCTVSb
2LZNiF4YHEnI/NHdAferWQbp36gPEYa90ZrHY8DVkCgRf33HpsmdgN9J1nfk
lb+HOC/XLGgiW4xgiSmplGCiAIL9t/fu9TG8Ffj+csLrINhkFP04tL3QYAVN
2tyXv22SOvh6WGjmNoQYuBjEOl+3sgih8ty1llEoQX5yxNDuVm28CbiDglwg
9xsx3oBHffLOrGrjRgAW5Z3VQA3Hh3bHHbo1qtuYyW7YzTygBbqsWqvpf+RX
KKV5VMcqtyZRbpxDN946R9cFvipkmmlk/0gSqWW9CXwLw1zD8MxkjPX2K2bl
lOlcYD0evnKR7/QNso9AzTDrd1O+sxg7ud1BmTfAr3UEuSeGQgHCx8oz/ntg
CCDJ/YV+ujiqbuTKtYf88zyeNG50joLKs5tbs04qJhQll/AluEYmKCh3Ho4u
2im3nV3NLyrX3HrpI1wSDjIr8+zwDWKU4XeT/OHonVOm9FIXQ8Sp+NMa9cAf
6DUFqgOEUIelJxtn+CGqi8EsIC3E6m88Zm5PbD8p2OKda+HpV01LCBboZTJ3
V9hujeVXO66TSJc0+UsVKFo9IXCVAir/3OuVnnUYqXNUZJeDw7J7CQleUqpk
9KUUjLsQ+h13s2KG6wJf1sUXobmd/+jpBk38B5pRZEooN08Xvm3ksKnMXS3E
+4HP4KKSCfpHvZ6SyBCNDlglKs8HK44a7sbX8EL2lmHAyTvi+pU7u6uGtRkJ
VYIvgyRUMFdUd8b4Yw9EmQRFjFOUwrmbXFtg7muntbu/puuQrdutoG2lJK/s
ww+z8OLsNKlLkfa47iRAjGWkmlcT181TpIF/GxmT/XcYr+SHMr5hVzDk9A9o
fAe52TBpx7DOAbfzqixU+vg5o5bIX1eUiRrpIwO0pbzGSn9KuPeJ3xfeMUAj
J7EglPZH4+DgZecoioPyk+FaUekStMEjvXQHBxHbDfFo9kh7Q5q7hzYvZmbU
Y6YpzpUN65j+qbFCApzzsodsFoJsDcRyCDBZgB+PVt289AypDsSqX/4wM84u
iLlDokRQYTag5AyC8z7ORk64bdjgGBEajwsFF8u4hrWrI+13QNxLFpgUsTuN
u4cgfmR3sS21t+zZN606cxoZ8uCCBbJJsXtFx88RJ7GO0h28oW/f5BJvLYVZ
1ad3m5tOOltLYIQwfVntIHGe8T1GpailR8VJ9XnWAOfPLsimS7R1Vjg7F0wh
twbLaKaOEn+8ccKqEU0YuYVbfSZIv/wCet3w+HoVxNCmbXDLyJRN4wGohvHx
JMXPXn7R4PfTXKWLeBRXy5oAbie6L61Fo54bRdUJkAx16H7yENTZxmHI5sls
vcZvO4lp4J8DJ7h2TgrZqjTXKRXJWobn1ILrb1g2+QS4tWBu8jrCb0XRmHXt
ztH0pdFWD+enOajDWTP4VIsr4DOEnriPr+x04h7VKUach8CiBXFwtbHx3f9F
9O1qsR8JTqOR+KxhCR9bq4nXvLZL6TmAD41qGbu44jdVFuwDRsWH0+vRvVlt
AokTnBE26sSRy5f1U/lLd+ayuv/710G0QiDCprXWEyDYYyW7cruXC18LrBVG
jB0o818HjPGk0HoaGMFwulJWwg4HTXrL+jg1VnX7Xpm9DXqD5S68A+P+mVZ1
CTUyqp/cJyXKJCFO6uJ+4299ZBFWWadDmm3oDmimY70PtoWhdoyPAnzFyZqa
aSC/bBDET5EFVXa24HcyR3wnHLvTN49O4KEhQTHvzrEr0lZFx87XU9oPNofe
BXzMT/awYHAQkFgIzPhi1eXB+b+svRG46/Sa3XAAHmNs2JyYCWKjUNc46VWP
6dPIyuc79bfwQrrdOMEZWDLpoYgXyTVcbBQq7grSNsCexRIH/x6qKiFyugwr
e4qdqpsLU95L4zZ0HmWiEltai/lLc4/XMtzwmXk1sHmqqSMuYeWsBbIJ3CcC
sQ9n9xkVLtcpTolOEJNeXHVPYJYUNE0bJAh3wygczzM9C2D/++6GEVgkpqaF
XrZeKbgfFf0D/jUh+PJ6/2e/TobY5mTRCO+uTC9pwlCxzE1GdzfEVRHq6ccU
L+5+M47kZFaCCCtq+3fGrs8Rg+S2NBhSTz5osaoIM50=

`pragma protect end_protected
