// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Fk2sznS9UrkopNF0PdR6excatMPYiKw+00egtz5npyN0ucHscNOoVJjUQPvK
EmxY0NTfrk7mP1imzFisAWp2MEZQhEXkBxOPUaftg+eU+AURtp+J0HE6ijii
9UpZ+FsGQ4q11h/KDuaheJyTEosdtyENYw3CHPF/GQ+ZivWhQCmhBJq3hPjf
jiTSCn+4ugzLKbcxBKcYR/atkfDtbBMXUSeqYZ/f8lgCgchz/1gjDMfmH+aC
cJTwuJ4irPHUPR1kqXAzX5LNzb10hocMc1/DeDMVQp1NiMKRJnJZRifhwDwA
Vh3lHWQqMRgGi9lNHtk2aUqaMW4tBST6bNknbLfLaA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
dDa5dqSQ26kA7+tmnoheykPKgANshawgtmue2CdpjhJO+a/nWpuyoC4BkA0x
YgShoSGKrxAAJdZnzqpRcjZsnMArTuGXJVSZlULqmZZi2zctHFkWvMJT8o49
+no75VgDXw7viTYV5/QGAKoZPtJSOl+QwZ4IBmuRAW7EJRtULCeb4wyJpwNI
lNb1UbEDRcE1Zl8WZMXzerfCMA4xi6O3Y7T0UjQbyf5R4Hw+oPkstJ9DAYW5
ZNV/hmMXG76D6fLEQZxCQa35S/npm8rnhJDpASAh91P2tvi50vxIozpgEBZc
4sEHwcd6BwUXx+qAb30xaJ/Xd8CY+z/hJjhfh9NWTg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KbZYgrGQwPKIDEW3hhNNi9IGGSXH7NCJTorfU+Sir7Hm10qI9otegFvlOb72
k1LCeZ4bW+1pMyTMnewL1ZJt9FxXGwENg1rzpVGdMQ6KiFs37ielRLhomI1d
cPFuw/1/uREgEld7j+hrYWwAgQ4eWBrhZ1CRdmlvfx81RHigUMHr/plpXXE+
30OnbqCT+cLCJ1M0ZynmhMXTFaF/5D6APFZya15TqSEDc6/PCS2w6orAB9w3
sHHxaw/WRKixIHKorIdz8fpNJBC1GYcMPXyEpbjaXkeC61Dsr9X6JH8uILx3
IDFRNL6hHYETZJcE8u7pCa3U+kgTAcSVb34BBIJhmw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FOEjUCCzquTiNUuwKgGzLI/qwnM9ll1xP6ST86Sgp/bJLkJ5LcZUCx7i/IgW
PK/En1F718o7K2XLfyCAcVcwWH5mbZXBVDUcybHxuRk9PONOdXKEZmJgLr5V
+bM9yaKeD2UFIh7MLF46cIQChaHAh8Ll1QmyDOPCsMWGvylMO/k=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
bBBvTL211nXTx7Yvc4vjVvVB1o9ax/FHV32NUDGVofauISuepLJeoFK1NAR6
GCPuui77E0Tmbi6Kef9SS0OUlzvNwmQ2O8BHh3CY2YUpQAREZ+nPt59WtZ7C
Pk2SPNIJ3FPNQ60JFAGc6y+uMz1qdIHK65lWNvrNSwXNkQG94HyQR6WPCHzD
aPPhp3T0sjjKR1+M9vtZPNVcAltiIyjcH/p+O9MCyu7sya9Eb+YcwGfo5j2H
luPlLeUS06PK2Z/vGp3ruY1UrTxFwy6F4xs96rEiwBw5XLx3dc9bMPj+mcgb
8T4IgMSSFyZRjZt8blDkn7xeWRYERCARn81hT8je5x5eIzyHl+0HZbHba2ZD
HDw3Md7g/dMsiuNN+9l62VYK40zydQtoLqEU9AKM2RZVBkTbOAd6K15tmNtz
hA6PDUnjgcKXwevgfAn7GLEa3CR1lkNLabr9E9OTpmCadJR/esOPhJmbb4LA
UHsUkVBajrttqCGjlFVjd4pUUcLK/FNU


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
uUPoT2ZhPdZ/koBWWsNyWIo2ikPLWCo+fQY4JLtKUUigLRr7RjQF6ufyCRQY
MN5l47uJxD9amt/SZ6JPTfcC8KcWplU+qafdz0HuuXRp6eAII3ev7vLi5wmF
el1ZCuGD5dGB0q8CkSJDj0kXmdnedoGaCEZJegjTqdN2V86/2c4=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
fE+qV4qNVJjK6iO+Vvuf5K0i1R4Is7V6a6UukMCU32wDCIel3U/s54afviEL
4y9GtKibRKMxzv/fMhF4cyz1eDfGWjteuQpvN+NUtNqa0UxO4hTXbQcZd0Aq
uoAdSYtP5emFrJLdhK/XZhWJ/cL4Me0i8wvuyt87yfwLy9euZaQ=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 37072)
`pragma protect data_block
SpCxzyw8cKZd5t7na2UfRDCqLbo8qfEwvrp7Ck/UAFhAK3fDxEjddW/hkgeu
KMTih0IkTNSJRNHMtOR2Nlbcff9TqQXr5RRwch00ZwRIg14uUywQuGARtM+W
Y9+JYeKzDOSIqk8KOGdZVKk0I4PHrTv5ap2b5p4Vi4AhEiUSAqcsHfrTd4DG
bQ9Dnef74Y203loi+I/FVw8mUytXHYOZ5Ln/2nFwT0V1JlAYJQ1YWpFjESNN
9XVbdoz7X2mLCrcfv/PCtUv8Uo/LIu/qNbmuiz53XZhr6CG0+MCJ+cKL29bR
FuOND9qwgMCGKRerdYViXvqPB7y/MhaHBhm+fmjM21ke+xwjEFADO7VP3AX9
4xhGnBQnw6izGu7zND9bK3UMWeGIE5VNxk3ipFcdL3VvU5TcOlP2CrZ0dXCE
XDpIA+TmCLwHdTfNd5Jx4g+t9gdJd04iP52qLy2tX55rTYEHayMwIrLFDbzr
nZ9jkdrJJ41t4cvRucQ02TbVqs4qHltvEOOLSqsHHAK07W0/Gt3HNysn4ip4
edcCLVPLfbifK73BdxcPhN0M+8bSqTjl2atVGK6EmcYjdqrx81KQWYOKQtFM
tMeGrX1zpW0HI33rjpQkQpEkumqN8cvQo2H0Zfvnjii2E7fX3FxFHxZL516c
7zMfbfmlgWbINL9XwtfxkdxzX41WAQdDdKaOXIQGIF1gFhQ3N1kC7Ob0wvjr
m6lxysexCI8LItXXFkIHRTc2Yf0BF2DAxSlVKI9g+myxXb2CSByrFqWa9jQm
z15mZAHtL9xqRbrvOzKCve5xX6SKyZJBCUysO/MqxngvAZy/uTu2Vz8TxJ+1
Q4Hltfq15tfLve5z5EiF946/TfyjYxn6W+RPcu3UYSL5AjUfe1tqits36LxX
uUvIlEGYIE1x1ehZsqbmEE+MbLnJVnolDrD1Mm3bQR3N+jxEe++M5wJ3ZxwW
dlePQn8TPutZLj5lscYVyWKOVDHb0fjWvhdIXm9c4eanHtRvvPflV/W9sGGH
jMZq6R1BwLGMD4arIKZye83glQiXDzmtvGZfnFz/Z2Pv7YPqd4LFryPp9tFk
DafQoRyDadg1gPcwE0zVCH29muM0jij4on3uueQTNx9Yb8a36Wee4i81Yhzz
k0Xnxvd1UuFrRO3UQZWGjLe1CLOGU1208Rg5zO2QTOmtOAWyriEqynTzHlsT
vBBOm+0bDxSMFLhezMSk+Gk4RZjd0fB8doQm6taI5girQWtr4TcUJ7S5u7kA
3r70jwIpuh3qNt7p+ehmP0LsOSDvzGY/9GwiztwD09MdJWwdISRLcBLUSrZ4
XHqGVH1Gl6Dkjz8758ySiIjbreWSh1nJdsl718W8ALy/F1+QyAnOnedJ5D7Y
O6LjWFswH2BsQpDSxSJv91vsIiAJ9fNzJ2jfIQYA3LF47ZDV3Z+kr9IvWxwe
J871ZZU1S2WsSmcmHKVIRe7Sf5mk9zo17UFDCkCItk8oTsSuHEwIToxqHMrU
yvADXwlYSCHJzCOBEO9uv5JlFB4t1rdkDCmDSvKurIAvhzlmRb3U8U9QmbPA
xOltziGMytlMuUoKNHbPBsUftT0hiJgqzaym9OHnZUCEUVbwhJXjwT0kNz2f
WtTIoZR5pd3+P6lVP1yI6L4dD/+FbaG8eD9Rn71zXI2r+JNajMIIDFwwRgt6
Dt+V3d4Sv7KFXuXah9nGQMNK6gC5WUPizUImjdqTErPjzEL79d2yMPO0bK2f
ADxD1DUXvKe0s/BcagSxIQfJLs9GXnqxhoIYYDKcB5QOqIYtABlfSIlIP+Jm
Kt4dAeGAXKa+unA3iEp69JwVVQOIIEJVgSFIuGrxUcVCsU4Vwk7sX9xvzYKm
I2RuGYziyNHsOgmA9/Wv8L6vea/OWRzqpu34Dq21trQR5xDg1LrseswZHaMN
6CmZUx7x7mKerLaK8hngpElte1p2XdTq482jyH0pFDOfEJ61QS+cJlplj4g3
HRnWYgbxaLblr4IdzH4biGLPUQ4cNV26mpG/v5YWaGQfSymwN4aMubGaMxbU
oo8Iexg95NuxUjB5BC5ob1achbScMOy4fTyx2dNLNootUb/RKNf4voj66/Zs
z0uN7CWns248NA1fSpY/0RJTd2OFqsAhYWZk3ta/9aMOFwVZAzNWlh3rml0X
0ZRDS2JaR+n69RM/QUdhnrjwn52Ua1jiznDIxkPkzCcHCWcUWDFAs/Mm4ZCC
l4QQeiNDYKnxIdFhSOjUjyXkHn48qsABLRqgfZk09th9N8LOEUKqCSBFlUd0
lRxehRB1mS7V9m0VNkMdg1FUrhDxHo9m42yQRp/JgT7mexhCTLXiXSpCSKXS
MT+KwSiZZS4tdNbPMOWf3F7RXd1dwS5h7auKs+QVQxOAcaCQZYqm1SJm9qKA
CCUZ15aW3o6RZnsxyTiOBWBN+xme7tVFJBwBegBLBLEI29Qnaw9M+Ws8qhEu
ZHJqs+7mhd20W9C/dtKEuvAPbVG+VTwPWry1quLT3uS71l3VYUOCcEU/55qg
pBe/d59FP6k+XxQOs906Uql/Xx6hhXLjLnb900QVWiIo3JtIry9fpMZbos63
YbRSSdLVOSmPm8tPiR8363K4y/qPWm7wriFKNJsmxZPtXcwhnN+wYjzGfBYG
J78IjX4WWu1p4It39p7thVms6kGviP3NQj3TVZpRBVh5Xrbf04rN1uO8SzFE
vdaa1d5uaDQPhoSt2ebTPPTv15hZPl/FkwhMzaOeZVTBJ3KQ+mBYxciWpRyA
d/VjQOSJaC9DUOMd27pK8HBbM0fY8tBG797gCWlSVFe1q89zc6PIBFphXh5R
S76gJWoboTCLFFc5cQB3paZb+1WrPOvegRkxN9ZX8VYksjWlaHlbzwAFo37X
AqnFNs0XesqePnenidyR5cRhkNzes5UIicnz1BCQUHQ5WNt3Hs2t0MBbs1jY
/7F6GmjCkm9HvndLTfwkQUdNEdCiFUaDbnxCLJbNZYN05/HZB6aYQT00Cv/C
rDhNGMbY4lrvzsFXTBCwtBR+j0sul29QPlVe4h6rBh5jsluy/4/zTeXgvEli
6RWLo36ej9A6Z6f9jokgCrunJ6JuSPfU0riCnoSA8hYf4yjVYfW2zWJSoiW/
PmwnKl4Pi5LbLIvYRxZ1tLoGYPdG2gUucHV/Hlm7txm6dInOvqfuC5v2Pccu
XE0N8OHazECV8LLvHUr29NB140D9qfo6d5pE90t4ykAB2dZQHsMPvUeRZwEm
VOzcqWzKUG6qocVoIBki/oPSQ7qielLUa/v6kMM9L0qVKxJn0NogVekPihv/
61PVdN1ZUfO5+YvwQiGWvOhdGRWGNIyBkUOVcNYMzZ9Zg1U8gVMPrEOV53jx
effUGo2mu+TrISwEcFGQmJVRuwPqzfHrx7ekVlgFoUXeB4St5C7WOapU7o03
WFWEGkOk0wslqA54gJpMLPxr+wnHxV9+bB7Z9/dHUjoc48HPVrc0CdLQUzNf
JX9VTR7GMxpPm09ebvTroakUS8vzQZ2eVQ2LoIp1fz+3A+i5kFjnFR6Teu8N
aDbbGNRVz4KmybypHdddX3gU6QgA7Wu2ivNVpxGT9MEvqkIYt1ZjrHlbzorl
7Z7FiIrK08dZSOvz6rpoS8C2RHJhdizSijbxYSkAaGSsZeKI2qa734iO0xud
6C/KZFbdV56PG4ldpFvxWVj1UIl50A9HvbRFqL2AhijRhF62Arm5XYmRiRy2
RG0H7LlrhGu9si8pYrtD2jeqNykLBFb4O9itLJP9vPfkN5B/LZsxj4OPBxJ0
DcutM2n6tjyPMGddBjMB+rH9d1eXX8sP94kaeQG+fdNuMeXLT3EN+4gbvDBp
soeTvpI4eBmId9T6PrTmHjAG9G5TezYIzBXBORpTuIWFPtMYgwURqXZsAJZc
qybYKyj0oYjauQVlR0y2pfstbmsfeKe7mFT+eeCMIPkFpaziVXHaFsgpM51D
qWoxH0BR2iZUVzKYMGBhpI9UhIjHzVDKvRv2MIhzMufQp9pQ9d/AWJpe0vop
y2eS0Of4GDy6IbyLQbiwimD9xr10JVMa1prlZf9up1E6h6j/7u9tM0D/0nhw
5OqeIVk2LSPV+adEKBKbdbp3vG1oxkc+3Q2rvWj5UB/QAmpycllmftXlls3f
L0CDD2onpv3MYIskS6pwSMN8JnQgtYEqvB9OPRVUK5fM+s7n5MOiyDhsK0Ul
Si95TKZG/herkG32Ib0HCXm3crZjbk4epuP8QPLGzJxZzgJPZkQHMTr9la4O
X+9WSGubMwETHlb/xiVjyw30Ho1fNTtvnvjOI3k34A72SwiGBmMgwOQOX91P
ynAYDf08gzHeqPIA9AwtNSdDQmfUTHuQOgDBDHbCb7ZcRGfWnNpcxxQrqyEX
5UZlopXgw64HdTAb8e3ZxFsr71vccbEAtnRKOWC8OKjKz71WDw79KYSjIFmE
JJQn11fBpjc4fBEk9IfbMdhkiMyK48/tT6nGmrv2vTn9+Sf7YXhee6QxQXsU
3luSGEBOiiajUDuxTo3va194euZzPEqQvwUnyZ7+cKtr8NitK5h7QaZYBrci
/zXAmHN+M3afu+6hxyBfgJ0b/SDSelmSdAzFsEbqtuI2nEIOOHsZxwldUell
+zz0nx9X92kk82H3WMsA7h3OkJv859aorjVSZfTmTKHYY4m1KD9K/GQg6SDc
8YR3TBl7YqlA0FnExs2+lR5smZ0WDWJCpaXGyVv/JqLzFBIwNdUcEUfXM8l0
qbSKsNmxJlEeMS7YkUlh+tpgTJChJZ8A9WUoVpvgd9V44irVrkriG3k5Dais
iYLL7BRkqQCHWOPe6NoRWoMJB+9gRm+nL2g7Yg32E/ls1eKYlOx4N5wPi2Ac
HC7kvk5qD0jk2sR2NxZzXPJB0jjwnnR+rwg5MKPJUWeDgrFNBpM/ytuG2iFu
aj892BKgJTJRROfvRH3TwJH1Q/m4puYRlYeRKETcseJKAexmtkiCpVDN1YNr
kc1+k2SmVckWohYX1FmUnmin9vThixfYPcN3nY5yjm9zmMgRBLoXaACZPJwJ
8JCs2qXX4ol7FCFJ8GhwMYEbafbq/oas97OCZ7gGLZQk6JxmbUNjbJ9CuRh+
3lwh1XvFzWYHlqylawfktXT5NfJCjziDiJumeMn4DVQelLcDHqfB1I2kgIq4
V+L1i4XNq6iTm1IYa6UrZCQGFb91tViuGs3kt48tWGS05UQYcOciIX2a8o4Q
koQQiKoL1AyTmhBb8IIdpLCu6Fu1a1Ot1fdiiOT6/OGHw+DXUrWwHNl4iwYz
OtYv3Nyeo7bf2pvyGqZtTw72Oe/Uyxnw7vpYSEtnGTjj9bd0NwIz91KDUbv2
8xb8RWeU64jBbiJD3qIpuRiCYsSqsA9YEUbRJqtXQVMeLZ9XwK5BCfeQuhm1
j5W3SCpS4vABO6zACuqj2Ss42D5lBCVdKkf0e8W4495YHiGcRog4dYU9SBAd
ICHob/iay98vlvi3AMn7xn1m7FC65DQ0EIE5nSzLRrPq8KPxtkiX9v/zb2tU
DBU6Ebdb2vTss+B+7bbAOhd3m2jPnle8KsT1SAMLGonyx7mu0aDz2vX+vwrV
rv34yInKuefAUcCmqdgwkYeTlEkhnALDPQRS12+uTmP/mAQTE4vG98Ali4Lu
kb2uPfN16fCG5Ew/mu82OZRXd4yapLihRSJzUePM3NkuxW6SX9jfiUFKe1x+
osyaqniCnl1gc0Od9x1/OLPZ8Xo63N+eKE1gPr/svFc9KYsktuJBpWZEMevX
FBktnXq8zEmoNpOoX6xtVfFYZjiAr/dU2fH+gGLfHEJheihkaFHS8/5UZZ3z
g+cju6H2Je1KZ0HEwIXORyWRbgvfpM6o+d4pBAXbsi7Guw/e0vIaMvW/l2MK
iDA8Mm65xKAQkcpL2bQBg/n0jAG+HsMhLUwlREpA8RQKaiQGV8Hzu7Z9dA8A
RqYeHrgN3CJnX1eMh4hGpz55Yy7Y5nfObCGtM4qREjBBzxT1CDTbG1ZTTqlJ
FgproWyYCdjMw02O4datRemvOBOkJjp1j87LVidmJX6y2GURLBCGw/jt/FRC
vCTd5zw58kMluR5btXI5kSO0XBv4IcTr2ewo5xIQJXFmd7XdvclDJ7QbscN9
EQu2wcRcytRaKLpmdvvhjC4r56BBwooieBaIFPdt9IV47CJIXZGdQH8uHWwk
BgkAmGAr+r1ctv8PWCf9t0JIv8TQyKB9i6yHJIpRBt4D26CcSpkD7CrIbfH2
jLaAk8+oqnKDj4vEDUwYU2iOhyHZgp1pAmPl3B1NK/lkFP8wnmTqXCgFbYtV
jVMghLFdb5+8wIrvKiyE5sFDyfiY2HFA1HqBSwXA5KZIaIxdc/3bTBt/57yt
SlLpTtvEejfb18yIbHT7ojRJ2M6lJNkdfjcMymgbQYA8rv+VJLKOpE7YNzeG
l7gK3ycwZUd3UBHfw2ytbDdSirKFlq4jaLwLAjvJEnxnuUDGhbK7z9YToRRC
7DnHIVqoJYtJao1FaeNUQS8+8XyPmYf6bLvbRPZPrpYTcm/0/7xkbSXobCFQ
oAIMS3pwb5VOOXFwQA/ay50NZ01prv+8Yk/AgeDPvs2axKOQocOBqTV4IsTF
l3vmDRiulqtg5dkflbyjK8uIHZ0TrwjF/RHY36emT+er0XdUjmvpHumnuvVQ
qB0Zwmq0GJIfe06i4otoJFlToPz3A+7zVHVlUPOIuWkumsADd4WzvyjyZcOL
Y+fWu+LP/AYxq53RpRugCaZBv8Gx8K0YPrzE6lrG5yvn4YyfRIGF89GJYnTg
Ryug8TWEQ44Xf6c/afzNVVGoWuElAfq5PYl87ArGppmmVagwJ1CCOMC+VMrs
SLN7lAhpi9HIdXcPtD8Tvl4EEcElEw0vE72D6xhsxnCdNCi4PCraPhP+zH1L
4ghfpcWmDNrd15DQaavlH/EwvXndaqpkKd8/A3REQf3JpwhpTZVDfpzPvgQ3
8jp82GhgNB3pKhpU5LumqGjJdES6gD9w5ZLEr53YcTesOv7eVX7BPTopwfN9
myTImokHxENWh2/v+BCAdn4kJewDpZSi5V13P/mpqH3Q3jrwyB7rEwF9f+F9
mmh0DrXIhRWxec/jj1fcKuZKI2YeQr28PLa+eoLPAM2RN2kRDM+f1i1p9Ry2
41G37WRdNzyAacYBSx1Gj9W8hlxMPrWIL7MOVszSmAqSUl6EEUSLWBkwI0uT
B0s3uUSA3FdwewNCNm1JmWD+kbBgEkrvoJNPJcXNVrPazwjC3iZVBq2kmEQG
iy/7OeR9NMc0OY6iJV1mPf+hdqibrQsl8jbO6EcIhqForEa31spJLFYWRe6m
zqPDj3y6c/w+i801DSKFjzQlExI19DTWoRANWhDgB4E6ThxS1uF0UfSLN6Y2
jOzepuc5DS5JU8oWFE/XHneUQ7x96tJPwfMgnvSGxM8Vzk86UFG9xlwXaj7f
zQQxKV0zcKmW2ENSir+IkgeQnAmW0UhVLZ1uXHzIOIXURNfKhR8kPsaPEpDe
ntr4x25tBM4TCfmaODUTfP9aXY07KTaMOxlnqqW6TePUfPUYo+4Ws+A5z8Oi
nwegCZie4Mv4Ly4erHYFcltYtwqQhLhMQbpFWiwpmgFQj6G9xHKjCG+1q3X2
4ll51PCJ8Mk8E+iEOBBCzclyEBDI5noIb1Qjk+8G1VKMZPwEJy/TmlQM8okO
K2GH8XsS8xvvt9dFS8oXVR3RReNtIy1ew1BUKqgoaq/jPSLtj+AJeo8eYhBv
zU+gc8xMe8lmza9DKVZ5mF92jk2w1qkEhjGLflAOokzdka+KdN+CL8mGmEDK
PiCEItn6gDa+NYAXvDk6quWG6unAe22o7TfJW8fVf1nWnk7i7FMe8HBXAkAL
2e5slOae0wabLHMWXogGkyBXX1jRTwq22h+Jgqog/wLZgcgq8JdupdyF1Vz0
ai7NNcuoOR/Tu8TxpJWrT9HR+lB3pJkbDgp/V2cnsmgZs5iA7JMBDyYDhroN
/4OoBgh6mAHqnvafYyXrHaaE9VZKUg7TEdAbfkuIxJtXTulQxlGNxBUJCXr/
rECDt7+XRqnFZQ4G3qb9O6pYPCx44ImYTjK2PCruWZM0XxWC18kL+WP6T1io
Jg6Q3ijc2onZtE3KJiWN2s1POGdzUEyekZauTOtvWlxcKkfuvj3YtIk6XrWC
VHVSQ9KjgtYekP7+yrCRu9f2xygLQVHgzU8dbUFlz87By1bfgWPI++dK1I3b
Y0f3QvphI0lRv+7o9Ps8yonD2YXkuDlD3Ap9BxVd66suJR1KmCLmJhZRnsTA
BSD1eXIVcrlj9Lyd0tUolWwRPukPN4rUUWAc6NX6gk1UOl4fqvirhZKTQBea
uj8zpypljovKryrrx1hZ9yMUjOwBnuzs4mkC4sZ3sXOKFKPuemtYNx6qSEAD
0p03ZMeNGujU+Zalwai2vyv9pKI93DjI7zAafIVNNzwcTuY+47uTDJQDWinQ
kosfI2RE56xfvjE7RLQQJzwqvweXPG8AKcMxeWj25p+9Z5hZZtka00c/2e6Y
tsjHoItPF7WhVPvsAP0icVePTmfDlTcIiOb1ESC240B+sYyMidNYdrwlDzNU
lwTEqwpos8h9QpExIs9NXkmk7OQKlw2TUADgNuZsUl9tySs+4KFvkTNfrcf0
sLsnf9/j7t16iVMilUE+dYNagFSM6K+ZlXC7J2dU04/ZGsG++Mz1KgP6yXqT
vAjDeQoID2ts+gZ2fb8VxblFsrhGOYLspBDpwHSaN9nN03fn5b3bDCFux+YE
LUcnO4pVl8RL2Xu1lgAyFsK/xwCHpUcdomgCapPJAazDY5SVJ63SPqmCFEYV
0FC3kFbWNUQxfMFmTfokyEYNjCCIwXemML92rzUujyICOM3ULs24aVOnz4FC
ASLlTcTp3hPmZdX8PweJCAw8qtyTJEiZ1nNivUB8eApa3vM3p4Fosa4lR3Ix
q2YpvKFX58NPrp4ilUp3LISnTWnB6hwvp3rr3wFCUp+AG9KzBjM+lIvpNo+d
KPSk2NfiqS2ojyM2eQtR+e442AUmimPCCts4i9znU7IrMCxCGDsdTeRuBwYQ
qGXS3de85BdRQcic5+vDAlcq1MxI8JF+KtBjMPTjdUAE411h5eN8KBHNNkCl
CynSZd/2ysCaitfEcGfx/94IPM5gBZFoxfgybDZcO+7fY0gHoMS+FNDnB1Zb
doA3t2MvW9vLC24MSuxXp4Jo0ESjQ6z35451l8VnjHCeqDpsQNza1GBuM2TC
DGJCVXVxpFW4TswM0dsDRkpKC8s+nZDxoxZyIIz09a98vd1vNW801zYUlqGv
Ex/+ftCyXLgzj2GPpq3ZuNNYAFKSsXfOeq3ZJ3DWnjHbW8L/VeFtuWwT6B8+
EvXq93t4mWxDBt6aZdHHPb7cMKpLG8zqrmC9YMoCABAZqpTuoRPCynMvwv1e
7E5Ftn0344UkgnJjiA7GrdMdCpBQycJGRM8g6L8KlgVvNTxF6OSsss/l/K9H
lJ6CKAIqCsqmWkGpuCyGzLxM0JZWBaKiOzNCaCY3U0Gxd4j6v6g3HLWGAA1l
vGTnNDOou5Fb9Vh5aR1S0z+HoDkDFd1ufAVmMyqeXVbEj0rAcFT3WJUHTL7D
LzQy4AKXQxWm7zJjn4nAd7Ww3NPy97Ds8qsSI/ZhHgsjLTZDXNreomojT6rz
+PmeCjfzBaBtImcWSqji9xHGvnVWWupc9VlLffICTA3mvbOBd6vcQhidmBln
Ujq4eGUFtNc0D9MWDAGQ8SSK6rIWytT0MfuOLPkUVY23fT9mMG8UHToL0ZTt
X3uFCll33RLGbR6iDq1YYbbGOJtl2EuKy0XGqEhYuZMY/SxQbK3z5s+PaUvn
OB/Il1dk4ai55L0BDsTrhbNwpjAUiCwAxLoQHDYXIpVUIQj3qHflFcLXYfhv
6fUyAhbhu3rkaE6lmERLXjHE4UH5Y8q240AslCFi9USIeOKIhMAUyUlXFA/q
e3UmcAi+togOxLV/56SzWrYg1C1rl7nsYRb6sVeZoUsmX5asAF9o3edCmk9x
wtBnUpRzAg/vjEg/C5sMpITrNhcQa2fFkecLPZPBfNe/EZfQ7ekFIKuS8Qqf
QA6uAF6QRUnTe5+I2eUeGD3s3soAyAxmFQ0HdDatN6zU0Qu8YcPGUw51QA6T
czivaWtlRQWpfMZtdTfGD8GGNJGGw2NluLshBecMkPq+4ilzohfHidxdRCCX
rv9hi/D5O6Xrg0mXPOPfg1f7RocWZPx7L8Ag5Isj02IDd2aLKjgBtAJm4cqG
jPwOw8CSOhckBffr1Ggi+sj7XOeLTBrNtiYDhw9LHIWe95yO3j/dD6YZaEWi
rDUfOSq3PQf8eptxMfqCP5nZZdA/yrFXRcG/W7mEc5dmSHGshmdbRWTztuwB
SKTDZCDyApUZ9WDMha6KjdGnwH3mFfNd4DmZdgILuMN09YPGYn3m5mGoB4lC
AkVeYLfNJil+5IWp61Jwx5uWHa5cSH8HqDO0HbZ+xrZuw87YeSHRLGWbth+C
kSsKP5tnJhOcZaBYoQ7ake25dT+vMaqtMQdL8r+opTOCZmDcvpB28Akf1stL
bQ5EJqTmEda5QYHJ8enEnoDaGLzxV3BgP7BT1iydBoV4B3ODu8V3Cb9JB15F
2rHAraXPscVZ6OGzMKBavH7vqWapvBj8YAoJUBXz4iiaCfvVnD+fG0Cr4NlE
nkykR60q3zc3RpBH1GTLM8++oSiQ4VQ9JPk/gR7XE31wxHrZrXV1pQd/W8qM
jpkRkZIjp73Q1c4NpwlmDByhGSd8daPF2JyjOurQt2nVJZ43shU02aAdqoKj
4RODsClN9HfILPKQHN+KPOqH3gmNFqWBuBNtpPES35sr8DBiotBUF72oDcvf
bMP9jmZuFYyu46Q4AgWL3XEfQkH4WK9Mqzz6eNzRUC3kJ2gdqhMZxBsfcTZk
SJDanzq/QmxAVUvTziouaGkIbkoziJadpB3+jIb2Iub9bm3EHp2k98pMQVZX
WTr0RWH0YWI8DQ9NiaegrlxxOv3Lx1Hj0ZO4pK1aOAhGwjvrr+RX1Pw/JRAo
GxgwbZXTizecijRC3z7jfWQ4AsqPm2m12gfgx6hG/mMv3MYN9lw0ofN0RFJE
or8rGnXqDttLjNi2HQQnholYDzvP8yQK+yMUDrKV4XUr6z04yMXzdT1HxOjr
sXmtq3iJO1zO2T76LAGm57YZAmaHb1EfT1rkwez7EU+62d6PKYYKFcQEPHF2
uLRihu9wapdGyJnKmyjL0AorfPR9GffGq/NdCdKbCi302Ailo74RBwmrZPR1
0tbhcPn3Z5/J5A+AatQU6igsuXsN7Gqow/PxP+RJfFnNx7ob3aK99GrVQZuD
yxwkhWLo9zbG4oYHVd7bpsJ2tB529RG/Ps2PGPogk7l+tvpIcX5S8ODvvpvD
JiYpClFrJ+rPlWHMS30hThcDxOOxa37YcjTO2M+FOqAQgyNPoWJanfebbD9G
9jI5apqAK67zr/cNMwWqOI4Vom89wmOnYldxqjAeuZXlOioSWUU5b+6nOzP4
yG0WJU74TPJcneocHlXh3PcSdLZr/Y7Insdmuw0YARgkhRnv+qpdb42IuT3c
tJYngflYCdt8t9cBixj7tXoOWvLg280tfWhZkdYW/FKv929KB//hD+zKw5fE
JlSoUTRfA1tuJYzyoStP6HhQjGbV0uTnUWzzEdl3xB+cdhDuBPLmC66VmlOC
Zns8jcZ9+sOS2QNmJwzku/DKqNr95xVkzw426gD87IgmJ41E2RWCx5la/M3l
ZY2mion5jtX+Fy5uLMoT6UkLT6jxwYJJ4ibEKhv2nSb94XzTXdm1mQ+C/a/0
xR2j1sZndtpdBMbNP5/SB35WdXFmLfSIaJIESrobE2M1N0XGSJfF4Qa25LMI
UP2DpUgMFCOd+xsQPRn7aiivPSaWfC7xM+4/LJBOeq/2xdwQyuqd9PGUnP+W
oqBsERq+nh2BRPtua9R1zNV6DUr2HrVMZos8YP+87fm9LDI9DrEIeepjtXss
kXcuMdIs6+3EvL4ebtqw5b+x0uPgKkE4ir5aqfoscuLk622zIioLZVputikc
YYMtPehSMQ9A+aFzIEzjdCKIX2fgCXBZpL9H2LsK3LofDCo50m43US+oj8GM
6wxsESD3DCl9VOI0yMk94/9EEXKq+0ge6FVGS8jkgChhgtBoVxKhOmGrVF9+
yXJfOcyaboF0M/PQ9s6J6rAa3l4WtgEapankzPE1Xbp2onALhp3VOD4SqtA1
Uw2RfYMqIdvtXOBxGIBL/DRMWqh3PLwa6NP55NvH3y0rsL6qXENRhaCTuXEw
OSCJbgtelEB/WplvPFZdBa3r+eqUoYmgl1OzRmppXD5DNnEasfjrC4+3KZj6
7LGXo0A+RHcrDRdYQdySy+c1ZHX1CaLlJAjF+dlOViNjfl9duiuVDctIq5Os
DI49UousL91V0Vk5GIZVk9qr66fdOOaWEhSNnpKaFH82836boe/yxUZmneAB
EiRuuFISXgRDhcghWnWf6mBxHPQzkjCTDYimz1UgWUkH4baf9TC3O3MV1kZK
CH/Ur95638xKY4YVPbOd4L2P88CZnrBA0hOEoEqUbtXRJVgOj1EV6cW4cUPS
PKk5R3o7lD1W222pzm0atXxANol8Z4monO+3KO9+4LCh9FGK32oWcudawZo6
Jp+Syr4QvMQEKosq4eEP5aGQqMaW4lqADvSMjCQOqQKrefmmrZHlv3BZsHkh
mb/WCs5AZt1n+R4M7sIqJkeQCuYsEdVuapAUIq9MNzyZ3d0Xka9djgvQYDFG
HAxuMk1ke4xHOR/Zwe8wxpcw5+zSW4cTMVMWd4YtECq9uMaI66kWYCQzOTVq
wqMSUkSJHYiVUQ7Z+gsaz49AcibBH92wNJejmj4HXr1B4kYyOZpESXk0f1LK
GXHlFpkhCrpYvzSBLJsmTfzK51Mq+ME7kBwNbe4UXC3PZTOfTw6mgVxZiBqw
/q18xQesmJu9jblOtUOIu/CIOpnj8ikmg863ahWRCXZca3thxtC3g9IwVebE
1BJ4LGCuP38mPLg5s0aA2JkS7iRZJGvvIDNuZpdiO8ueXDCeU62a7Ia9XftX
wqrc0Ojq4ntSSKqWwAdFj+p9dIGax4gVg3exGwtURb4x/HRuHn8ZmZigN2at
QBWu9p8M3BlzJ85CNrSnrfq+ipqKLkqH1wS7pzFDIJRNBjqYzuQTbJyAb7/K
MDoradzQ720jvcK3SQzQFDSZ5fYuz8L3q4U5pIIOiSn4/MEk2nQtOYfkMhgF
yOLopsi4aOhwSRI31HwlCdGq5U/iQYC6byFa/VCYtjmMIeVIGAzGkEln04ON
Mt9ioqH0SLsbaAiKQBVagX5fBz4j+wQnWx2Bm0ys6mqiZvZ/tTeWKs2fr2IL
97Hr4h9LANN5O6BLRdSFoYN4TTbg7ATeq6c6SX8CHSK3nEJ1/VxOCqSa23P/
kuLqhVGyQ5qBTGlwwbxWW59Vqt8r+EUVCaW7O+XM3wZAwqAM/cwK4TA5xxLb
qDYwi+F8MsV40v/0fvogohWfrS+wbELAdhHn8/whYR/8sV9VWuy0Zqv1xEUl
M9R+TMbgcMjd1JRtjW766iqH+tR+mQjDLEyo69f+CCCldiIWhgSBXaTNB8WI
HeL/PvZy1t8U5QwMaGR/d+frWoe++Yp2qklxbY5MUivx/4Z/PG5F0K5Xn9dt
cNGMP/0Cj0EoQiMyy1YksEWkzasaKVkVUwz1AsAYs0S8jpZ3uYlqDMNOV4Pu
0NA5OJ2UJpBmHwgvJTOwQXnInMRWY634GwXZGY+tZg6kelV4pB3OJUONkOQQ
nQhkX4iNiPLjV3RgHj0FaVmzGbmg8SubIG5h7rbIuEbQfwd9s8Q9xn3Cw2Rw
0LLMIHHy3arpm/r/VqbM7GEgTnWZBzpS1Ew58ryNLMlIzb1zUU4WDxCxba8+
v0qlbaLZjkaCJmzNkdcOR7rM5/F7DxLvTBMjChLE5jifiGglf4ZjcewMuNZQ
+8TToYEoFtr9Idapc0ufuJG2hLWx7cZMkIrTM3JtEqX5rP5byLQZhdu8kHzt
RbsaiZIjixqxfTV/QqYE44/AtzY5ro+5Oycxzm1HBLrLXw141RkcJrdCbtNi
Ikedp4P86O/iU6xvEmion3PEQpFkJbw2KyHKWvZ2nMjQ67Ozu3bk7jhHWLUK
Z4I6z49lxr+ILRm16VYX3TbUlkRp9Otds0OPp7vLafc1e5lb4E4XXuBD0UhV
HdoVJYXdkMd9XaVJV/LvCRQ5DPQz2EfkYsIR2/f5TE5qDFtZBNb76Y7+8Qjf
uIQmFrUglMh+JQ3ULSdhjrXhNrZYxx9B1szH89h+Yx1f0qNc2Mugw8U0LxJb
vFMx+cYn5DFVRuHIc0gsnza2exXkRarLt3lXdPXdlTNRV9XYtW3qF/IMb2+0
w81b9cs8zSc/i2jR3/Tn/supXqXpy05weR0PrdJo6fZe0PXFp5eLoRV9E4wa
h3/fZV7HEl0y8/1YPDU4q39FmuOJyBP+gQt3jGK99hKKR3wOsqnH2dZ057bY
piXviDO0IMk5iNo9dzMqanVbUQCKkEvEW4J33CTV7+fFKYLVqLUFPahlOmX0
W45MDH1lMeijzKJdUkGgNdG0g+UIy5VbAOM7TWPKYRx5+zG3d+5vMh+sIkA7
ZbjNR7C3V6XzhEbAkTXiBzyC2rUZ6Sof1vtCcRZvH6ZYOAf+nxaSERYaBOlb
zElVfwvLjvBWYU4VleIjUYoi9m+3Dq4VJ7gcRKYsLoWtwPJw0ROTLtb07ruB
2PhO7OmTgrycugGkqPq6H8jUfjGVE6wGtZfEjqkq9dCEurTp55L/2lvVRr1y
hv/R1IMs/IMzjJGv9CI9150g7WZRJA5+KG89rWPK4bwvZmxmtDk/n7dDVhn9
IdO+CUCdZUiXUlixyM+RnhpP7nOdh/0Qh2e7jQYaWLkh6XOZWcPGtJWeFgQD
2+pSsdEPrdI5+fJCJ0/UUyix46av7y/ijtCck9ds2eFC0ZgtUiE87BkTyaUH
0HwNTtaMq5LriA9RU5CE9pBQ0xGPFWfYqBnzKrYFUNDWHUhM+zTEPs3wlt+8
GN3e3xVG995L981AmVrIq8CMaQAGmTWnp8wXf+Op0U/Cd7B8P1BS5ZjNu6cY
E82+X4q4A2rGeFCzEKM8poVhx8+YZt575u9fqXQ2wNBCULl4G5d1LWgPVGsd
LNTf9xw+ZOD0vao766B2bo8gFTLXkSn0QgqFRYvsStsrGeBlSz2ak9bXIXFh
TduoA/uGCfX9nhD4MR1um6vUOYUDwLgCfIhvT0Hz8SX+LJDH+jhvZwurBrYp
QFpa5nOaU6SZm0qd5EnPgYriq6hXW7tzQ9Bdb89Nlx2CZxq955JvdF16Jt96
Xjuglom15R4dbczor9gRYdsqa3Ug1c4Uvd0QZ/Gc4WR9jcojdxEuxuIBebdP
Q3Nn9rdU62YexkjFBsKLtXa4gqMoQgt/qwJp16rHTPfN/Muhc2W4FLWCByXg
A+xTEcw5B5dkeut1Xsxrdm0NzFjPj/ynYlzVhHn6DV2HICBwlbYFdWWJKjFc
kbCNsg61JeKTRltie6JT/qzjqHqyg2mV/jpp/r/DsO6nghUwDfAODZafBBCy
hULtumSuP1u8k5UOqrhT/fnycGSMbLrm8uKpSXVmXgI+yOd2n/zzjAxDHC2m
s47RwYAGYm/bm15RilvmOfjz+OA4p6/hu1uxl9xLExwAIhskWHPYysH8Z8G/
xC2UnP+4G6BIBEYGZEZ1IlgfoXITIsBwMRI0ae5TzGnaVkccGfMWI8FuvmV8
JgfFHla0odWBhf/9fNhkeq3B/5EZJNaDnd/hNvqftD/TGzYOdNqvhJW0vJYM
ZUx2MNCBHcj14JdJJnA06ZngLQEn3CAgwsYl4H1vrwloiZdGGbL9aDTfgoxA
4wMpBoxceVTqRQsRlxb+NsIfuz26mACm4XLq3JHajL9A6HAXy1ipkF4CmHZH
Pa0BHkoQV8dBTgmPWt8BKS/IaFPa6OPm89Tvq8CEKt89d0JD78EKKuj305Dd
BYh4wCNDa0kVlYS9uf0X/c4+Sqp+hvEkDe5qgL+jUR2gj/Dq1+pbDa/DGJ/7
AGiwqWhJLslLXqgdr5PfRDChNBAUTIyAleZU4ERgxYUJ+/jxKijr7yY/ZoOx
pB++DPpMDjAd3eUVafYkFyNm0yXgRcW87chep7mIEKSGcEAnPWN7AkrPDgQ6
fDa4SRxepZy97QPN6GG/vtl4yp5h/D+W4FBCUmWEspI2htQsZZs4hYghLikS
vKdS66tad4Yhq82MmJhfl6vt4E+api+/7w0Nt5YAmHqoGE/QS5GNzdejtp81
cdZd0OoZVGxS4il9bS86avNvQSbebShFgVtcOOXETnN3TFE081dGKYryFLV9
VeQkjJ1EbqMreXqS/+fL6Bo+zevFbqFAhKTJ/yTtM+60P+qKmhgxoMxsDgd+
CzYWx94JTmXZAnyfJLTBWyoEaXFKMCFNhlgmFHCg4TuBPyBEUy62qpBfzRSA
750CFNKe9XwwVUXe6xmZJp/WIXc5e6mzFBTtkZFIeyvofbWi0TPvu9KLsfVs
6W64H2SSW8v16r2xV1T/pWqBsIvSd87atO1WOSSbMnZqT8xkF7cbzaqmdc9D
++fbtpIV63dIlwQMg7YnkSh7FXuu8i7vr2y3MZaZkgq5kuzr61KVE5l4yZPq
0DsdsTFX1a2GQmNUaMh6RpSXcR4HshPNiDyZgx5b8ctR1UeB21DY2TUpGLcN
7qh127az+y1WvIeEdcZqG6phw4jipKBqb2osXCJtCsTnslNd93hlad4BQLTC
OMZY8rjxtqdaGsrNg/nSwITfscJyJYNsNaSgDmUvw0nOQq+HNQCNSnVZQIpO
DNiLrO1Qw/Y/hBddANFuDBELkjDoeQFIUCc56MylqxX4cCR0fbaHGowlkvlo
q56keBJzXoLPTxJSiEQtna6fYy7p8tCAVfj8VYQH5XVoh7MtBMYftncFVM+d
uhPbVSX9jrH2CwKdZpflv+9u6Zgq5YvWhAIMzZ9xECwh5xhk9qpbsloqmPBt
l5D7Qdvr4Sbi1Ea/ZYyZ+O7uPLxISDZiFSco2Beu/Q+ob73in+pMq4lY56hn
3o2HtJWrzBJ44MNBVLHEsaS2J8MhCfxF2M/qNSyxZu6/nNBLEs/W/FTqB1Fa
Adv+JoVJatM0bSlNJFa8R7Iox0n23nPKIzy5O6xMPk4TFP7POwQyF1x+bD2m
8oFB8jN43ShDMi3RVuX20TjdHAqrkYB0k0sUIVoIbrUfDhUYgnc1K+2hb5HG
w7LS6RefxbBG6EfCV7PV+ggRhbhM5c+C1u60nC7QrDiVzEKk+6h4qOy6E+Ur
gnogprLV8Uawe9KI4LAYTHV01s+Q3RfQedqGicW8R2nNs1xJVL0BxrJ61R67
VlM3OsF/3o/MXexPFZNuFd59mVptCSF6KFC07Y5Sw6AY6sKQ9R0LiQ92WKlr
J7Nx7NIBmB1KjyMtnKtnW+eUfKUjJyDvSBPhB94fZfzkv7qmsPpYG/8H45iz
fssjQqmLjJhEml5U7Z/ysEq+rM9VlXJOsipkDC2uzZ2sp6EMMmptLuLhSxEt
maIMJ0RvHB17eEk6NXyszWFa5vzD2gRUfFV80znaGvT7a04Yp4pIDSrTvwRe
y2bxJLE2bzn4vHuEUm30VYpBIbdCcDy8v7C+mks1GpfFMrsYFHoNuTS6zcyi
dscsgE0y7/c3EATeu3ksbAPUZsqZ2YS3Gya5VA9t+8OrWH4myFjVbVPiK1RY
AC5D3lJE9y8WOmO2KmvkFAT6tYACJsVrejia6A452/yqb0djZ9y9vIwy5tv/
+OiM4U9pSH65hEmGx+jxl8I0iyX0m1MM/H0Y8iMEoQVEbcofDVD+5Il5z5Zu
GNRZhXqzeztyySqj7LOnmjcB7w3N7UThPzLsxJO3KwVSyae/Bd+dtMMC2mU5
j2fMs412qgAQC7TbHqQtdnBZgKu22poIe4WZKVdEnSvwjAlYJDmXkeo6QmhG
C9FFE7njXsiN9QxZrBb55m2FaPaiziQ+UoOVDGaAQznixAs7Iz5paW6Un730
T8kOQW8Ai/h1usEhkoFvPKQs20ud1Ipc5jhB7DpKSwy/Qgdq5aXNfQ3V5v6m
G25qE7mOese5R0M0aZVR5RfqY7u0XIoZkNp4sxWTyfNNXPAke6LgmbLd3yKd
SSMnSg321/80b8MT4RMVyVaiHLlsR7wv17MhFKviF55cclxSD9+2KIhjb5HN
wYWuKhrwrD7MT5zypsEn2asDUDUKMZPz8BNKkW/xTFiObiDcoRFUscR3OT5X
KvoPZ0YxUAvho1flOnxZnze1vwyRIcOtgiQkuGjOSN9Xop2iq2mUWmt5Qw8V
2XrY9esmmz+UXg+mNyzkgIoo7kSNkWl7xdXkhFfZvGzPf9X/dFcYYCOcQkw6
MNIDVT1e5Ei5lMOBSR2Go8U8qY+LFKjd7OLKQouy4Awc4Rwf0D8LAoyjZ1L5
7ymawya198MrbPqU01Dfmx3JObCu4TR8W4a9BpgpD5hURwalUua0ASYoyjNd
jdhz1DU/pyP/ZKVshrjugkmuJx2hLGNTo5xCGTEj8sKb4yx/azEnT36RshwP
m7pjx8vjkOeNuYnyhblACVJMqf1fo3v15gAbqoQc1LAc/gz0oOAmtynFeA1c
IWpqiNlCx+/wDj/67lkBuFzIHorn1cP88JLRlhdSEzHOtH87gzNdCHlxNH36
g1oPjv0gkxxq8QQrNy/vDxtL1bpMJQFccULb+WI+j/iMFgkmsDKAzoSi8LbK
VO5QGBHyEKqvkl0R2C/nRg0cyQ/ILWeDWVgSsX2AjeqovW81ynaK1dT0Q41C
1BSEjZ4b6a6OKGHoriXHR3xRMskWeJejQuDlEdTNwPX/aauZIyRMwxbD5vlz
K0XV7OR9qXKhOTDTazWqp6CwXrS5+DDZJtuXMH+62IrP872BN2ZmmRbI1ugX
Kron/q1gMZi1frGBqgau/8Gq7uvZYNMlYwO9J0sG+uj+E5zbmyUIyyzpfXzZ
SQBbs+ERFFwXrUNzm6AsR5x2amzILih+hwf21/qOg1ojrgrMm3GWqYVbYb94
LywkJ+YpC6QURm/yieNXomH+PLG2Eb1ZJrtJIIjuXLgtSHhJnmb7nJ5EB76a
dMIpz9lilRWVI1inxmX2GQHRMEqjhoOSTxocPDANwPr9K1NsgjbtQazCYx4d
ZwWkSHenOsnQutnLpk9aaIT1MeHjBwNA5cXWew9IcYFJvTyw9Oy+uPgCDSDK
FEXXN+Pz5IsjliNikCCCrUwh6Vo5kwRs/gfFLb/tRSs+Q+08RnfDGecHFKdj
KBJ1CAzkjwWkSUKA9j54u7eTVNe2cM/lL8jU+b3HZt6md7f46h6CLUhfyke1
tOdYEGzgm+AqQagahaNK2sbUyqZuT1mS/UHSOu+8t5hKRvLJGeQ0yHlp0jz3
u46uHYXjKnm2js4cnpOnFUN6422IN/IHBtxc/NRTsucPrio6yOfRuQ94paaY
Jsgb7W+DusxvjoeehtRF7jBJKst9R9X8BdIQtqHVao2ObVDRj1b1wnwXS67C
ljrqutqJVMubFzy3R+1js7Je0j+x1NNBr4y7Z+Df9wSK06FAOlP3BJNx5UNW
+dEVgjEZTnIJWNef4vuf3a2i8IYL4OPQj/jWh84tR0o/xDpK1CD8K4PenHAL
g/Brzhl5ISmo80Dpxl4ZAEgcPBPnoM6wysOs30wI5Ler2NetpED7l7UByWRu
WwctWt+ZKHNamGk0u5ddkm5zqb7/8X2XaVFbRJ+Z4B2uBXZYkmYOhBtntqT9
ySaIrMIcYLWB3gHiW3GiurY/OkcmA8Q8ccLQR9OrBrta4/8Gh9IrEIldjT/p
9Xy9ma5/fPyE25M0b1ORpxKdSCuqZplBZjchEHBRigjtWHAGGw7Wj1obtICe
Fz7JLHJO2jKmRXqiV2cpfEnlPpEWCoYuvT0O+HZ5uZBpTCVaKF7STONIch2k
2E8PRxFuM6BoQg2wlrbqpwayi4xU5J09cvdvviioYIXfBgSRVCG/+rlsSSSq
S0+BStkfGDQUpRJGNNAhnLZ/jDzWRGOMC0342BP8nsRsQ3BZNai3LiUn7n7w
r26IZ/MwaPtxlysxnEup+y8w2qDc9K2d94zxFq4cA5sM7tXKqhNbHOfbv4JO
xcVkA0oe+AzNGiPMK4aewZmEE6zvpRrn070pWmHUCzLKdndllj9JdFRP7jEi
qockkd8mkpxsMcApqeK3x7zKHCfbiU0yiBx3aGwTxzhyiGDE/QbDXOIXUZRv
MvAzBDexuv3i1rmHUDeiXATWVYVD1Wg4omPONjgKNxKkID2Aq47jDc/Qmtwx
pnilPfdX3Bok0qHP+UcvHk18TOEmmX/3W7dgQPXoA0gwhEsGVnRN7pRM7vWg
cFFys6/Mb8i9j1A0b/AVW/P/vY4Adfr4omlVfh2Dq120MpRzveWGVVcJpVuo
QoPsZqNbqq+19URf2wnYk27RAWo4vI8nkFsJqiwhoXq3O6K85TvVq5YM7npB
yte9f9+aNW/Zel7JUYuaKi0ZqbcLAhEn95MPAK2GqEJm9HtaGOMZZt6P1l23
QCOlavgcJwot4Mw/S33FiPuxWwLg6cGTHA+/lXseanVSFDG+vlpb8FqGXqn+
WoFrfF3NIKAl0D0+kwZos07KB8vAxVpZ4PIzgLJ9h+T5ncRSXhs00/u71quu
+lcJ9nqaSx36Ag5ZIeh2DfUdJis2kEcGmwWtrMHYjUbUnBAEUI/imK+e+dTe
lrDjITbxcrFhCuIf5bshz9Y+kN6RJkdcb+2RDe2QAWFU3uTLOkhtcF0Gq9Fi
yNu5r0QzHGwcjPM6bar3rQHaYFs013vYj5Pq6SSaW/Dr6DoBIWwbrkIocuqE
1kbgJaeBaTbFmfdwZRhCbrFnMEX7jD5l/hAVPK8Ecq0AP63bexdg1tlUECd2
Y4orsi1R/lJP+cnLf8AL4EeB+iIEaAf5zjofTW9ddilBLmVEBC7wDZf0/BHV
/iLH+IqJRqAUBrwGJPz+9gpR+PElal1ZIY3FphBhxs4PHzeZQ+zmDkIBxTGZ
DPZlQNZlKLbFpo5YYqXzsVqGtjqjuWVjw4yXMUQv8GGJaUtJS/6VChT7EANq
TUTLy3JNMcnmG56blB52RMqazgY412/vpOI/DY/IG3zoI7gCPiwsSn9xZC06
CU0iA25SKoWbDM4kaZmaEYhp2E+p1BmvhMkCxZM5/wV3Na14MNqDSYYIfN17
LXt41icVo2gApk3sBtNJvRLb8teWwghqK1fCmxfcumfqVOMl+Wsdccc1JhE4
DI2vh4mQkX2Y7th9VVPgr173Om+ykKis7KUg6kRyOdh0uaDnUSyW/7nx8Ypm
harjH3H7DVpoPotzjpUDoTPWG5fL52dypO/pfOb2eDSltC1gIPNNzUcy7LnL
QdHVCymJb26GmEQCBXecm0akIG+b8FuukTyEk9/XNITe9D2bzMhzVnFVatJL
CZH9beW5XEoFtyXM2TFc+JfsdHJAV7O7H+GY39wwxi/lbEm3I8dLbz1Y1sIY
jxQmMFKB9iqR1Mjzo5zY9hBzyKhSXzqhLqyhcwwiKwUad+bzOXiw46z5cmO2
HdAof1HTujmqCO5TBC+1/nq7ESkOSIYfn/jOI3jAgq+JxN4NpqyZwjXGBx2m
zVE0SqEue++JjZKTaYLZXvOVXB3z0mQXg+Wxksi5BvOF9AyjYe+MQqppMCrx
V4hJxg0TdYWKNKhojcm901efd+UBoXnkNaTdNrpJLz52Sxrsl3LaECADb6Pg
RqFaISkGiPN+ozTZi5VCo+oDRI/4BX1O4Knzmb9QMazkT5QSoL80Z8P1ONp/
W1h2SDTkUVJ3Hr6R1YkD7eHpvKpE9eWbwi0eWopzjcIMBqSgT07e1ZUU/vcx
HkdO+8gulDjSt3f2UIoBjQqlV1MkG4C2eaIvIuuzifIvmNgxKv22H5hZnSK/
wbbXJ7Do3p/Eq0CW69yZXupISZvud41WWsf71omjbfldb9B7a3yoXgPhCHt8
9xjcvPsbb1Y7PpXEtumMWvOKN8AcQhNoHXCaNmTLiE7Bo2iCTFOgl/dgCFVL
O+fFDOMqQRUwwqRvgGGHL3Xo+wn24XaVER0iQ90Mh09JJiZaPoVegodFpeIY
ZB+SpJ1td/p3pAKOHbuoCtLIAiBG88ogtDEY0Bl7nnbLYVWd2w434M0xg6Pz
/U8AdVCjaIxn1ZOKZfqtSxs5jxleyT53zE2kRUdu33Q1+p1AQXEtFFsz+oQu
nfH6DBOqbs314yyKPmnGRles1lkfcSXmyinvmkl3iLuQ1Epji4ZIugkYWk1S
AsRGjIFg+jP7LMq+q2AHeyzPWEpmXwRSWRiPHpn/Pfh+bt/Wh6DnCpNl5vG1
MM40ZuOjMMPivPzIVscV7KfaZ1UNHhf1bwKUtrXDtM47IVBG5ULh7a5eHNZQ
GlXkVIxBlongeo9Mz6r7Ps51EBjOybEuUzWGmbxQPhwtnbwymCytd7z1HCrb
cbe+l9sZeM9ENGcXooOi0Y0b3rGJggJVQCiD4jf9dQxBg+xAhiSqoa0HUZ6a
Nr4HW+IFSPVmnHQ7l17PpaAw40WGmG6rxbiL3cQslhlmdq7wzQHr2K5M9UPk
Mk3fI1Y3E43Z+CnEQ4qchZl6dJbCSlvN90SfFZ2yqXpeVUUxWEhZ/u/L+pxl
zxCo5Zgs2s63m7iVoRBRCq0PzjMegizHKIlqyojW47F+WvAfwNK9PaQn+dpE
CchMPyQ1JAFA6Q3CNMzP+S9VVOLAlrAYk9uE/Y1Z3LSusnX4gZY2Xfk4yfCu
t18t9S7J6oqi5cwrywfBhj9Mnff/E2WEQRB8Sal+EJo9JUV5RLEA1HXDzxBT
uj/wByb3Ua6QuFYpeit05VKvto1f1Xy+816XRKRKyF9WkQLlZElNXxhOBwxH
TWuQ20ORgYPWmBCnZkuWaSC6vsSAzdO05Ff5uFK7WC7FH2EZZnU3Q7fkxisB
m6r6U+sz+hKI4QAP2GscnF28GZKTqoIf7j/vD5DwLrTQze6KJuFzFqqfyeX+
7QsmewzLKp2+r3MDWnDFoq9tfaPoPveOhgge+WAQRojwE9ok7j9nxBErL1RT
EpV/h7DbQB3CY41Ehf2OpdxK217S37wjI3ci5/uTV+3fgZbnAoMXUJisiPaf
mGcdtMzrfV4lGSGWNNDxzNT7NjfLwC3tJ1IQ6T0C7N6jlFlHmkXU/9umroeu
rWWEFoLYqPhmcSx91ieCPGG16okDDglR56fTaLjoD+pgI3SvIrrfrsBncl7W
6WLQYkOM4veB1/BcmHpeWas55IVelJaZDIiys/idbjsrL8k845B3vAueEfHo
Sh5JGa3zwRLwYtbZyt4mBCZNpNjhlb3RieXXEjYdPBjzQpCc/sTyvUmW91UY
emwBq3EyCdO39tntVnPeiFG2UB/yxIO5u1B19I6TMY/XUST3YVEPENha+VkA
0FuX3cYgG9sVNquR/TuparC3407Q6qjJSgKU+iOQbyLra1B8+9JFjstqgCGz
HYRqJACTQrwgFWD2rTm+WcuwqhnNiWLXYkk+w7DybCG5H1vpR1doBuxCx0GL
WrGr5EkFldgZ9MufQSld2z3itGDt9ikPJzyyOBA9675UPk8s0FSF/ddk0p+B
Ji30sZ3liGE1TCnyEkTFi1cvP8UxkFO9BVhUVqZ94pVZQZ/kxc8GSRYp1BlW
03NuijoE4ny8ptBfTnx99J2Jj91kGfcsuYbLsxChAeOWMZUBoh9u4ruS9R0+
jTO7S+bjbs9WfoiaMiUc0k/OaXe3qO+mCQYVQ8MLhNpa5U12+dg1ob8NmABJ
dzvwwoxBI+ytixGX0xtjRYHovUCnCU/8g6ROTNpfUyYxwvsXOmLmlMlnB+QM
MccDjLLCfWfBjx65vjLZdGepXN1//o7etLqrrymfoayZfAt7efTYbeGojKeE
ppo4H5eDRvMZjmqVEi31EKLwEKiEsGeHFN2UyW1rodqp4qpwaOzpjY07cdaQ
W2p6YCYzRj1ofOKREsP9Hg0pzOhXu9BpUDNJKzeg90HmwBjS5zZ0XxDDbl0Q
XBZZahHxS2YVpgzRZApp+RBsxLoNz4DAv5dOaIJjo6zvWHfk1IP+oVBaAHul
liY3HAU3utXgq+cfAreUsyFvNVnZPCLOaGR0DC2E15R2+H/6hUUGC3++brKm
g8pIsTSUPp/a9f2/gkvfF+JELulO28WftMmDEzktr4Mx22pr/qcOIcIo0neY
gZSavhNlLmTlLl9GeTt0zYaCw0SFmAOYoqqsItnfkp1xoJbg/tPw9oNQ1ko7
a7rUbERJ9CbdbkI7qxMtJFpPJ6f0HNUKToVooQHCet75knx+om7JQrQkAxzV
3MSNQ63G5eQyj82vE9PcegWGzZEG1EL4xhPlv7Pj8k/69d45g81nx6AKz6Kl
LF2U32i/7lKAdH9lSNxL1LKQc3sQrV8Q+EeIdyREdzHgYLoJpaSN6uPcO9X9
kp8e500b2DNRjlTKJusN5nizFJo0ILgNJvr9jgNdlDXBaYxm7qMY8OUZaxwG
cLfUpn4SHxgXLzzaYVpeeSfGh96rLymiQ/3MF7D1dbqpH3V0A3urJUwtUbVr
8IgxmZIqM7rT3pB7bhZPSm8v5uv26jtN2IjCbVoZpJLSZfF8HFPSS5hV5nXO
OJt8M+2dFO4fuKQI0NWgOh9UoxqympK/yHFOxZs4Lw+ZHD7zzX/K79VQ/a3E
tIfpYkd/mYB7Pk9yOUl4U+V7xLZNSf1RI7cQAV2GP4naLKOdehw2YepXViku
IEphrMy9iVl5Kz+KlvKD5GsJchFmjiyMAxAJVJ2yJaZdNnhbhITpgPYTAdEu
L+8prLjGWWguYnwmC2wUxeXQYlFGuQ/v3cEv6/S94OKlELz2aUSWzVFbYfoa
1kw7GdarT0QcFTsvWKzutJD/yOFFB8zg1UetghXc7TKKwYmm3sMKnxwD3C7a
nZlFBWuiMSmMVkpwucf/g1PHWaQ7fYyOvECNFJUY/dvc3S7+vy3acPQ8Yqdf
g9BWmpO5Z2JINHKrJ8NeEx1qXnyzjMoqfNJqtAFPjs9dp32bmQV9VX+mawEI
pVESxnOfEvfgLlXei0Ek7re+6XB/TwBnLcL5RcJhkGRgEwAHZ+ros6Fpodwv
nyOm/N9qDk3CuFAUWk4q9U0fuIf+xdMGZ8Ga+qQCqHkG7utoskOfEdDeTqU6
zhcHk0s2VY3R9rQe88UkYfm29MWTuJVrOIZVrAigksKBpDKaiNUwCBttpYMe
k5MlN9lMV45rbNzqjil/cpa85sTQF5Q55LXh9zRzEZOrg+opUpKacnpKuSsH
TGHTFKzTGCJe0jCyEfmJ5tkmG7yY1Lcxw1TmwryJ47AQg+L4O7oc8XrKci/F
qenKBuFrb7g5HHKQABOwx793YuNrnIRlMPwViTr3Tude6UtMadK/kaVWQOpo
W6Iotes2DAPOCU+0rHJWVcc7krai3ua7M1If1KCuFOPIYf4SxOOofLnG/h8Q
VimUHF5bbwHEend9vi14jmbjXIe0FWZx2siJpdYGfw2OANRQBlF8Tdtqld5h
F9HkSDbUafy0gJLsNPk3vrFj51shP7ujFMuS5ZX+AkUCSqGF1tGdaFwSkOC2
l0npYD5eTaV7QAKiUntDOjprl1ZFHRHTsykfaxxtuoaYDbbbFFk74a6pQ4Gv
i/7hIAgH0z3Fx9afMl3MxwVdZFxlqHj+PbaXquFvtVYq9uHhDMHlhG7f0M1t
T2mALIVLAhElaSqfchSZES8lRHJFURs6DcNtcVFKgW4QIoYpLLw4L7efLYfb
sU8q0BUngtlFPCo0pBuTtDQmCq3TMtYQKososzsZFVqQ+vijsGZF+krTVQFF
6gC4EdIvpwvQk7Fej2Itx7V+s/ClqywzBoCwaJHZshz8+YrR226hhXSVbucS
HzMka/RjPzUSlT+4R68invewMOnpf92H/5Zu2LpgtAc72zgIlMSWHqbxnp5q
fwZGM5TdbeWdCbfSeS9wSJ0faEB3bXOeGatoZmEKNG9pYh02GNxLiDQ5BL+K
yaPuaYznXzqwSLV+SxpKiZb0kD8q84hwBkIAQvuoGfyzFZWMEKz4WI2yuaoG
zgE26oreFNVCnTJWU0vOoh+UouZ/qB7hzdtISWT1OzPr+VE7HaLlzBd0rJ/S
d6gABnrJfKnooraTXVQqa5FBvRpL2kjieSHOWMy2TOn457PigthRIUGC/Lpz
2r9rzWWnO94kxCXyYzg/XEDnMp8rrk1re69sgPY4feh82kcxbvRtBEaXH8Yq
rjSAyW0Zq4qIeZShZKZDA5kllCWgffsOGWYvSFn8G+5dy4doKSBoTkaSvwqV
GjILo8VEoftu8aW05FK7N6+35YGRYwcYMbt3dvcUWLkf+bva/4LyLjQtHkkm
TIiSjQcowv4mEm3D2AEnTFcGY17H5Wvm9cjoiOi0OVhUuJpXPKRNVvI+OQuk
bx8qWnM48r21LngBKaY9pVHk/EowkrJGIrZ9rUZYVh5iMB2BmQfG+RI+V5Kr
o4HepvNoNQQrjzvv3LqTGUrli5Hv0kn186/CFGjVusPk2HxtNmHOujYA9gwT
QS8yxIKBqHGASwE8341ah7Lek19DV8XDH7GIyYCbXxp7ljzel3Gqe/qhdj8k
UOU7OJz10Pw064Q493e2oIdeTZFg0Gc4q4O20D+b+r2jvYPe5t/w5SyATEZ8
hlbvkjU2qjqfotm7TFnVRb62ABrfc6VDgvzfppd89Uu9NDzUeLNHrU9AxC88
RAsD4MbkPo4ER72hgBGUbnVo0xwwpdMw4kPJHy/VtTGFRSIqfBwov6epTpgR
I72Ujk4p6Y9f7I03xNxjfE4JrORcMnv04So7Rm36FHqm6aENkSeS30X/fXQk
kdOYJs8EWoEYnIMFrugm+tLuBD21HtmAMjMrFxQKV/gzVjMKCpqkGBaA/d5B
ZXxajMkNym03LoXpYL0XbOgrXEfGpTTYDLMQDWNPSDsG/MhCAx/IB7oumz+/
5AyK3+S3hbQyCIogzvYsD1148NNJkksolv4g8DvizsfsV7T89kFbSDxdvxLY
7bWG0x9P0U4Jhun7VhmVm9HaZhwwhu6P/n2Wpl0UxW0g4kiHayUzJvzAhlAz
ICLIyZ+DSdinvT8wED6e7IBDQ9WgYAMcfwAxcQ21UqsdliJ71CEOIIekE+DJ
w9azorTMa6mfl+kIN9jmXAqq9TqirACwfTe6R3pC5fxqM4ntonnhyDo/TfxT
9NPPxIpzRoGbw7ST0KVp9gOS4ZjKu6xjBIE3lt3j3MjNs3ZcZagIEa/h76bv
Hc5Ui2FXzgaRmUq+WsBxLab3FFVlk7jzKw/LOZY6Gi+ckEJoze/KvriBt9tx
jsAOAUFxlkXzbe/Ni/HMDW28C47XKEmhXB+/E/4od8yqcUNdQ6/lnO7p0zYQ
LFJT1gqGZ9fH2GTeizENjgUkBjyrb4ftXOlWSUWyZMeapJla/98eabpx3KRA
vn4xj4ajJtALhCaAWbaRX1BN7pnDcaeFngl6q7uqQwo9bVU/bWWLlK5ZxdOM
WP6VUG5uusc7dL1/XTp8gsw3Ev26CeP93S2Ej1H7rjSUB+jfF2/RXyFlvH7z
1QkJ0uHlQ1cnyMEF9DbparqBSRiejq0mjDWz/0cAOJnfkvnvsR+Ytw5eoG97
76Elm8mU5JhWbGUXu6h0d/fKsW8vcivF7xvFcPKZD1Bft4s8RM4JhimphrFS
scCQuo6KQZXpCzQ0+s1xkr7BS/Wit+nno1JssEJFqpcXWGeP2lIUazPEG7MZ
KMuDx8eolOAYJ+YwoFJrBoYPqsBcccONVHCP0J0Vcii0qH/SNcZ44fsTk6gM
76e1veQSrMirZw3HOWVYcp+RAexYbn1HXndObTTpOI7yqCKlXFDxN3nsNyr0
C5jptvqVHdh1biORBXD2BJDmaKhZ6+E1ET5qmKTJRmWqRlpk/+P0CkEwOoXw
HL0OftbTVXIU+pA22PraAylL8qElTaMXYzvvahQfUSLkDxp/SV5zfzArRL/F
9YbdPEqeYIz1dxGwUhHc3eysE1XYmsEISz9B3nahF9dxPZ48WAaLTE12/8Ge
bMzZBZRzSNqY+GKrr0v4BsnCWumFkP4+vovJ9Lky+2PkcINPHtLVFH8X4PfP
pVB5Wrfs7Xb8A1uVqt7VBDPoV0GpWslGNlNiRbU3idEyo7etoEDDYph6EfQb
WkNh5g8RKsjSew4s6KCKxZTwU7I6Ywz/rH4fJRP8kwybdXXySnpwBs9YBkZI
BVrAPQCA3mFQ2wGSGrTAZ2r6fZVD+bGB/GpVW4PLIvuAlAXmiE22mMSy6qlF
67i7ZwPlVmGOqcy39ffbQB02ee7f+0v41dlZ/YGmYPLmr7i2g48HWDAqKyjl
jo9ROeqhsOtDH0tB70fj+scBIJxKsqUtGYZ25uqEGfDx0OSfmNLxnIY9l2uX
QUoPAF+HGtxUqIDYFMYkSotuWp4bAcLwNPY7PDACnXrtOrWNG6y/C7BKCOA8
y7WJrdcU+sARZUd2Bz98ch2Dkl9N9N3roSxi4lwU8L/+Nkkz8OCxxrNUhUUC
HNld5lmaURRs/G77X0+0hqeDGtuzQLFpewaMO3PG5SJxAEhSopxC+uWzL2nD
h7zHIqOoKgI+XBQHCjSIuuRqrnoigCHvQaw6ZS0q3vchhqjdqEQVDh/AEwFG
wGbPt6cCieo9UBl0lqa5XGif+gWl+iAUmkvDVII4tT2xsNx0ce73NxVT12hq
aB1dyTZnd6uaZDVtPm9Cg4InA5x26sPXCLY0v3+pShjqsQ9wLlmXE8febHjH
jA3b9yfMas5qkjWHKHw8UosINcXTR8HCDT768XaVTQbi7FekVnA8oYX35VKF
SQycboM71XDaUWXlcH6shqKEGYU/8+Li9cZOFVPxj4joq5RyB//RnNJuaKba
5S3nt179WzuGfAI95yQuYciGocvIjjA3BQi5zHGLd/7oXwzrudtLtV+ROdR3
C5iQPdt0fiJYWVaEWRR9DujCV6yIOJzKc552Sd+VyUxhWQrkECD2p2VVdQ7r
JARq2/4jeEJLsMkWeODDPF+V3OGSyuyodW7SJfuZJn/la5xe6250eJtsliy1
wEFFhsMHsFEB9VKCKhNLrY8hhzV07ZPssPFAWAgN2Jt/dsoJEV8iKVHAYK+v
z647xrNDfR18Lggxb/nA3saZhZGmxb0vOUIbL36HOlVXrwEf+0DLjWLkeztL
siLCHizhir0vOSlHDOGE5x2Oiu+H6Us2x/8W0vKpO2uXHC1n3kSP/dyKmJAh
2RSd8J/+AkVP23RLUtJrh/dx6kSg63z+ZWGARhU/z5dVvhkhLEwxAtsm7uFQ
9wQriaTapZCz4S57szKY+vcohnF8FImXYG0hupCIqxpI6M91gxlWUKFSTYZI
64BU7xe27DPBBVxzxewanC2F2J2Q5sdBcu0kVc7eYnYO4F8oa1NBHA7Y1iEb
QWgBfqRQeaH9YPMqnSo8SZ2xyJXTBYVxh7XqAB95e7Do82xRQsfgM7LXNq1/
pwdAVc0dsASDzWefMcCm3nTN8YIczef3Hd635uG3gjpVup597wApwr9ybA9d
ITZiy3vXqUCl7wCrb040vE5lIFtaG63Q8AvQ5blVILjQsYfVc1yxjG0ANqFV
R6WqcI7NSvtRjZWYI/zJxWLHH7XXRy+tZQTlrCX8c2PBdKVXVR5WqaZSBKjw
sp1G+wZVqShC54idHh3BvMVKNlRfRnnKb8/dpyeDOhkLR5lXO2P3WxvPUTRT
8KFJEJ1RJCuZhNv3rY7TkFqhCYs2JRV3Gda46whgLt+p9SMkxWI9DF+5k0y8
BvOXFVbR479aMdIc44voKCjrtZIjtpRYkdtCM+bnsmDF/cpQ9yGeI8D1/a0R
q+FtyNyZAoYLY9GptU8gyB0jwWntQb686rwVGfAJVWBgYFYWklztvNZZykyM
BmeHmhDilq4vLfF+vf2U3zvoitnwV5ZPUGAOJ7EERmhuwvCrR67mZx4eSXzK
+14UR1MsIZdh7SLlP6NJiHB7XWqwirYVRS2XRfhXjwPqlStp/dj64cEsJeLF
ISjyS1LS1bjs+j2GrRx5+u4yPrccNmQwc+uW3kRMY2VVO654UAYwiBSRBUxj
pkFE2oUho2S1Gdsk2nrdcf84JdjuAPK3PobMfvHKNEbL+xj1F+C7V14Djww7
3+Ip/EeUDDnPxnrL1Z83gFXlDQPmtigvgFG0FRSG7EhPskYrGRx7zRAkGF/l
sQsGY+74qgz5vNkS1+1Xwsyi+H6v8q0KXfpj6xOFZ6V3FOF8L2qgOxkA3kSl
DyJia8Wpm0/bwC27Hizr/JwHnq6h/DT/H2hSGsYXqUsbK5hcXJRAyQi+tb6b
tDSHE7Vd4+kVaFoOE/dsoJGcUyDTEoWfBElIejVv0Donu2VOcEIPMpQu/cmi
KUnAIcul/csYJ7o4CLybYvQBha8aBjbp/AHNdCaCaoylefl6e/2lzj8j2aQR
FZv67rwNXmsFgYyjwTM3/A3FVvFCZjeCd8v0aU5dCDDGkSpVyOKn07lCETp9
To9PQlnQOJvDfVonDD0F3zfovaqvTw7lNitPr+y/bnp2zfBmNGT05TGIrI38
MVqvYfuOAb+coo2Ni6tfRxdEXGcdzsb5+fYYnBvez1UmnqjevrsElUgzJYcv
DuOWpHL47HUH8cC/93mX3058Mp4wWadJddUOeBOcOvSLk+3U8QjHxRcOhu52
rJj9xn11raxoom8akSd2xqLM6Kjy2ohWuaxS3U6z6DbOBtCBwGhk7JaEa8OJ
qetzk/kAjOHJBv7MQtAS18J3zyNtYk5MV6G2TiOHha+tNEicJ4A2wtNLeQED
MLN5/ZTYrlkWAE8SW9VbsBddeRh2hkA3vmfRRamd6olb1YjaN6WKf5zUquHm
m7DwbfYkAJE4tx1yCQmuMN5V6QkRZyduMgL10tUDabjvBNa9zYog0in/z6F4
qxV0CM+PV8YrwVFlh8r560Wgm12temNS+qoQMH2fFtNBqVkpcyPGC1sN3PS5
c2WDf4C9JY2R+TT2Y82K69nlH/E6bbHQ4qQV2MfnP7jiIWCrmr8sJhRXe7JK
jUy6La8ebDVDNQqyEgIB6P3hqscXScaZ6jN7BbkthMKy3pQutyj9SicInPRb
liNxsaMju0Y3gJq6ggnoMIkwOuO9JiszcM9AzWPZGCv2VvwoJtKvwmsGQoeC
SKpZf66lgkzj84a5zVasB8INMqIkuVmQA1AXQFWtphnq3WYQTrNYV4iCmFRZ
AgCX13gqQZTihsZrU2VqtfPDJsL7BhnUJ/cGWpqXllYJqQRVXlzL+rrDbdzz
11AShN0/yjcKM47eDr88SdODu9u0bjGZHp7/flR3UGOnh0epO2+oLYZLM2CT
G/OOmuWA2iznZK8W338Cy63l7VS4hkuXkZk+N/a/DqBhJtr39cOHxgoDC0DN
jHkMvplW8MW662+Q4SowtTmvd43jLOR3GSW6JVdpHVbdK1pg5g/4tpedVV/2
BVXlQf4eG9jDKgTVHUXkzK/xvcmEv5f7CHgs9yvqN53PPXes5/347RcHEvsf
5ef3VvfNWdWdNM8io1YsI42/OapqWAOoKOtLut77Qe/+M73QynLtSbI4h1k1
TsFsVlrBwNY/sxajtpXyw2EWQSxuDaiUTcQrtK9WCPi79hny2WrQdzfRvskh
GLuh9xLzhn6/tBULwdO7fFP/2m/rj70ICb/f55zpJlbzS8uhwn/qyvspUYxA
tHFKqZLWGkxQ8WLZwC9KaPuS27Ejri4Iw5V6d2vlHId7Z1+wOB2ADYbfCEau
tnV5L2WioT5ARCSb0yujGb9lydTObTF10vAh6bcKTlpX1A7TCxtYV/jLn8iv
cT4WoHaTE+mLbeahMuyeKo9EMvgnWscWfFlAseq7D5v8IpFVfIzQqCG6ElHg
BvezKcnoAi2qENK98xtEZ5Iw5gkb3mDRHw4SQNcLxqxkhjKHsewwfi8Ql3zJ
hdtC2IDA4avTdwdRLzTMnAUMChx3w43fhEO/7+jGxGt+GdHXwFD2KdKyo1lO
8iteCb3yDESKiY/Jvpd+Ugs4R7I/am7qjwUJKThd5OcSfttJyXclZRXBqy8O
/3+Qn020CEXLUIYTWfKEOgNg/5uhAyf/qPvvxQ5PLyMEXLilUCRAXOX/2k0T
/Aw0hWQKnw0DPhGz7v5nMShgmesrAcZqjsq7JJrGG3QRx2erBhzMDGpa9zre
7UI2gGpU0CRwZptkzznzBTnZH3YjVT1apTmEJbuYhhmydX8d8t6CiFuR4U/2
XQSygCjmTqAOpBOB5LdXdscjwE/HTONPGoIbDbFAr1CH0nnR7wSllgLD/bjV
NWsUomqGIpdDHrJlCZ61BTy6wWAjX3H0Rj/Z8AtZ8w0vIr0dyTtVmhmUwUEE
WriangI4eupP70U/GYThkysOBq+0oGFump3BDvsrlLANslSEQyqBcr6FApsM
KwJjm7BYmnsD1Xl6QUljEu6Zqv4l1QkmlpTCMiwEXDZj+Pau1Rv3KawrxF9P
oVyWK1oeBPlguqGG6xu1LaWiyHJ9grrX6M5XyB0GoH5OtKl+to1XBbgLcmfe
YM2XkOmfIatu4okWrJdT7ibf0e7hoN6H4iD4Zg/Zaok8kd9G/ks7X9/ertqt
ytUEnmzcrXxPYhXMhWh9C36vnE9qhDGxDITbfXkwDGwt7zQxFIPe4Iynr2a5
1cvNEcT7gpXKd/LpfxyifxP22AC5yfMHnmMpwonbhlyCZBx6cTZF//qwvec4
o303bK6cmUs92kEf24mJNzd5a9B0NXyDH514iY4HHWfmJKIbP/dRwtj3vOGv
Y15zXtQscfl+Pb0Y6clkGLhf7G68E0hvDHn3hWUgxiNniWW8W+aYgEh+fiu+
g9UjCkEQBEsQrrFJK54gKwpJd3LD1dSbvTxh/WDLScAGg4fNaTwfFKCFH8N+
ilAEWZIM3XVEtcKdqPdjFz5sltqkR6kF2CxjNKmBLbHRbl/wqAWHz0pUcc0d
6IONTkTmO65vckHyOWjQOGs3xPcEOBeor8GwZ/wXy+0PdS9gPmICrWWJ1wWY
cX08FUZzrjnXXcs33DKaz9S5ZQZmFVoUVVbdi65T8AzfW//oL/4l/9eliTuE
13EyOSRHaEJiBKu3ZHbYUPhtWAhDqFtPRe86N7J7FD4c13G+8RELR/e1fTCC
665UffUou6cmdH50dZahuXJ/v10XNrSynj6LEcn3OrugUKjd0300Ghi297wk
8Jw2ZpZ888NBn5XhLvHpB3yZbJ2VdfhwHgSIHxwd+mB4a9RbnQo0elpM6gLP
3sksH09qnEwk0mFnfPu6Lj0wIFBhCNfVcR9aXOg02Z1hHZbfeWak8ciGSl62
ck69O3a7uQPdGnhVhi4Dw1ELd5zYVvyNJETBnTfyExnKj3BME6Brz3/8i1M9
qbXgPaa5iK4I4/rYlT0h1QbJMIqqYBosWH+kQyoBoHjHLm0DF0c9IkLqOKEV
zd+51NUC+93dN7Do/eGN7nX1noCyCb52LYiW+AT2QTr8nwD76EERgZQ8LeQx
PDUSAEIN1CsWuiMaZ26QwZhGEb6KqU2C7LyPhs59AuV3hk2b1oHfSmrrturm
vX/97n11Sfy9wTxz9S6UmFRJEdGKS4zJZc74kpaBYlGU3k2jVIgZTr3dQcR1
3Yl9x23mAFmpsrxTpXuAg35lKsgvDt2NoRGEd6bsZARzCYAHIub0LqlZOkNM
Ol1mDKZHAxBfnMtWsFsYkTuKBLnkgOqLVwdr1qHMPg4tuFpH36LZx212zZFl
bjsviDfr+nYX7NbO1NHeKp4XdeIwY4QZyBe9s4gnEpg4SsafBw/z+4M96auG
QUQF4FUZLJe+CJgRT/FarO2gGaNfF864xVjYvM7MPvPptrpagTJgUVf4JEBb
RMQDfnn7LDIk/Xv9gdDTI+PD0O2Db//QGHGDw1eAq4+cUgMrpljwFqymR9Lj
JalG7T2xs9PpllRZWdVz8jwskQUUzsiZJAv+ewELan8KRwo1CNeFC7jD9bfn
PVei0ASW1KY81V36No7zEwaaPPtxEt426gusSNxddTKUHN0Mk07C6EtJjtlz
P8YtzIZ7I3TZuztE9CbRYXOylnGajAA1eTgOpMvCLUMA+2uMi9gdbu/6PIwn
PYYmvRW5RAwVgRI9Wr2SSbarWQLJ9ofCI3Cmn0Mqhk5A7U2shR43UN8Seo/a
azQpUo86msnInREWFqwf5QEeqkzMuT0GfkeIxqHtIxu/G4tVzZlpFL14Zumz
71djjjfewHKF7zkAh7s0RVzxCod1VXG2bz/z/KDO3QlX0S6kolfgNvt5NrgB
leS3klnouR7cbfIIG6MnFqr0IbK+axaRp7D0W4eQ89eJwWo2o/RQoQoe4DMM
zJqxb3aFmyxKkC5CNokoUUlryyfdw1GatHDArkOjkOdc4MufIf4LjtjAKcbv
DNHI+l8FUdBg9DmArZ9xSQFLsxN0Dp0lWIXwm2Y8Bxwkkytc9gq2p33BZzx3
IhSW6ctwJwe6+nivJJJ1e+80T8DeY/eK8oFXrYE2DxIYQD7ngJPuvX0hdDEI
jT2kCrDFopkG9yKHrT9xCgsVXNSvUTOKHFye5dNDtKy1i7M0DU3xgnTF1N9Z
HGXAN+y6mQE0oNfb/ThxAOeRNHA+reG78epSmbaBnsp/WBI2MvqLmVNg9suq
VpmIuc1vUI3hid+ZPl94/dmRDFZ3kwng3gI6x+NWO9zexhBgyktAh4n/USxO
FuC7d5jn/Y6Iwj+ruGZF4FqRj0ob/B+ETR9o0WXM9eHR0ukQlFVeLEJ6lZmn
29XBLlpwXcjrVfRJSP25J+5laJSmfZdFgG0yLa2KW5E0uyQwS03DPCtMcdkP
TwvaxenXZIdVbTh7vPa5j2G7b/yPCuiWZH7CsCVX2T3r/tIRJzF4BHGvU6Gk
dffLEwEY12HPScodZnsURla5wWpK+cIvqyQ12C8GZErQl01UBIMvnv6RVIdI
Unlov/UoZoGIvbbDXzArFwPVghRA51SAayE7Zs+hs2MmYjQux5Zq0pPvslBE
7liQ26eL0ViWghqcjzVJHlb5gcoHMXNbAjd7v6qIVtdqou04BtIksAIwJLXi
CthKkcxmbbWI+FTW1/K12JM1Yzci+0r5NxkgLvai0pcZQBVBEG9ztQbtFgHE
w1nOkTpL631rgJNd90muhskoo9TzYdxjyNp0NIiSFo2fH5xjAbeJTn/UJjnX
IktXR6HNXEEx8J4gqWtfJrGlncwnd6V8SJM40pUv3XRyeAwLlYmS8UEyZNgw
8jL1T3ESCgFNZnnwtu+u4uL8B73llaKDAjB1gAHH6rbrDzo4Gq/wfUpfgyJa
vMYajzVAmojM5W1AEPcAo/p39LkLu4up8/aqOKqRC8GpXk3vko3hlJQBY5AA
pMppN/mx0p70YfsoeL88R0h6hZiw+7VZRzOiFT7IjaYawgYOlzx+4Hca5QcN
pelNnuGoiZBOERF4bpvKSY10HwQFDodwdGaAS/TVnfYfB1c1O2e8oyPcBE1e
cvJZEC7ujzj5DDOYu36LfsZmsoe+v/Xi53MzAnS4UingPbbWxV1s3UgM/r+s
OLKyDZ4M2lNuDPVvPXPAnywOHMdUY9cce+RCXV5YE79+9qL+tW1rKapFnbiS
IixWOjWgmgiMuiy7dhCHecsao6Fx1oA5YFunbARU2lJKobWwrmj+8Seiy3Lh
bUCBgebEXiOgRBtZYtVX4LvK9aynSwjwQHLkj3+xm/a5zh1hTi5esbguwBTx
FuWUPL+spsPOdujB+maZOqE14/2P2sjUw5OjG+2BvkR8/5+3zecUdkGga6Xz
G1OVfD8dDuoT8gYArGjYDER1iKUwHeHQa0LAzzV0wENuwCqDCnt1oXPCTyAA
jdkW7P27OHIureB+Jb5yKRDRAkoSr7iM3rPRGsOIE/agH7RoTl1v/mbQu4Eq
NdFC2winfoIC4bR0U5X6O3j0S4EZEdrAiicLUNrjmjjDjRiTQhpoO/IuMLRN
3FyGX6JUNM/f2CGFSap4NXPPiEUx2M+khAk4ypYvBy/IC36sjIEwv/2na0KK
1Go2lhclH7beYHxGtih0C2nUQzCt2ak0CrHEd8AQxPdvoboEm86PjAvx232f
UcIp3AzVafVGRuwi4Ww8wY2gj8ZTEkm4p+G+IOW6v45F2IryOzcn+BnPQ7/V
Tay4/LpabsotFaAp5WFSzwT9irQUaUL9e5p2UPiUYq+5f7h0FZJevVw7aJWV
FYUbRm2bxqHC/j9jIQR1X+yo722th3RTNvb2q/YpXK4m/tAw2X4pFmBMLHyz
WnK0Aj21Ol8O8RusF5PbhKIqdf1k3vSaZqygMEX0jAwxMR2JtbCfVXxs5sv4
13qY8DjtPBQUNdhD9nMedzKs8ig6AEXedM1S4QZkoesrluFS3J+ydjxpdTZN
hyLhrknwHOJQanm4sKbZwKXhZhORLVeVvpPvGYuTOh0omw1teTH5szZTVNCe
4zc0XqkSfTKfKDR7J2v6PaMMhhU2/7j/qA/7DVlHazq8S/drscgaq2eWXv9i
TtyosxOQZlPAFWk5e3aAoPgrqHXUN0FIMsyeTLPDMphTXhgF66EE+Qh4N0Ia
UDeFr5eCQSBrDf7Morf3s++Rty0Vz7p3/i4AhrcO4req9Vs0g6e+4zvZKd45
bIPPGGXXqndjvaFOqaOPutcBOjOySBVArby/o01NvCcOb9NWKZk4cRt9CvY+
00UvGYSLH+ztfvku7qkEwdienRABe0TFxKFzJYh4W5lk9lhoSQxUB/Qjuhsb
jHO2vIO76LnMW98vOdTlStkkhzpPSwT3xKFDY+WizB8j21sMNNArxrzR10Es
744F1VFA3Mnna+30zIgIGiqZM0EZJPE3+m2+U34w9xn7t+VUSoAIcRe1NIgY
4Sjv9vetbDTVKTHAbs+BhhngBk33goZtJrg/6qCCHR98xg+bfJBBeXOntTdH
aTlu358pBxDuFK7y6NHXEF2ek89nOJQlShp/0jfDgyjepbxMSCRSE8PO8eG/
8hFWX37bYEmIxSsKJhwC3pkqnJc7cZ+I2Goq7pu0GlK59UlKtUZvdcar36Bk
LsC3UcsnnfTvbD1KJTBXQCYnt3vzwJYmhu4lgbxENlOV7uA3XvEhoAP+BV4o
yIPh488l8x74HvlMtaMJRkwtg6N4IXNdT0Aygg3PJns/QjhzWjajKrx1Vy9L
Y1U1UaBkU0W8mwPZ4D/VxGXxKWNPc/oQuSJHNaNz+PggRSzdhhAzChojus/6
/W0tp+4rQJU7UZTkTr5ckUu805FVJDqSZGudTMnvlUzmMtkZ1M0uHn2SeBp8
Yp3wH1sCDAXb2Cc3OEatD3F1NTJsgcLjZtoYA+BE4Sd6fYqeTgIHkNBKfxm8
7xhCjQjxYQabgPTWFJ9uTi8PEbjuPnCQc1Nd7q2KZNbGDK06EiFOxvmMGNL4
nao7MF6eeaJEouVeuESiRyu3T3XqeghpJQG2aU15HwJdM+9Hs+maQzUEK3dA
X/Y1vq4hcbvK7k28gHEVF/AqEsZ+U2bpLN0gYz21jxxbHA3XnGjyqohW3uXY
4xVZqFFwpnEZbPmvROgM0SY/yYFpio2hphJcZgRBKUIgjPrJkk4QhFA7ZIpK
ptSJe2QqH2Xtsx1j3pLLpkQwsejq9dAjqroVbznzeSIvj9tdqDEKunHAd04f
e2fuYJtB4XXiWIHAkeTt70y3pjZ7Pv8y5m29DSuBjediD3GSgNjtSHB4xktD
YyucbfUV/XVJ5DBwfRjyxqXWzoSpAnlVtIGpGUYEz2JarGiAJme4ayvhlyd7
m1ulbpZXOgrOlGzzH12voa91DINt7YAiN6SBhTZAaAzMArHkO2jyiTq0LHCO
rUKZ5edJlg+SBjyFHJOfNlumZ5rsWxLNtwFyqItNnM6WgoAHyw1e/UZbQPQH
KzQLqr+goZCrwcBQhmpUeTAqh9eyMlWJjedabS3d9QOLw5MOBSo6ElKmhRM/
xI014BR9tHYsphuy9P+9l+xGQoEuDoLJFU7UkTKZlotJqVGPmeMS4XOPGBv9
iT9z09NDOrm2r2jNgz2YctQkP5PIe59R+8sxgIQwum+2aT9EVXHAux+4hqKE
E1vL66CmnZln2yGt0sD2FUPwW+5OzIAFTiNOe0BDXV8TdNeUpnbiZlFi+7IO
1BQjVNFMJnDJT2cHUFFzr8FVFDmnP3rlT0iMgeeexLBhzaaq6urHQeD3A2km
ykencDd9XhLQdqtKlcBLyYfaKWvnB/N3OC7Qtt54oUdqOxMIZgVEINK+fFcG
UIJPOeML53+eDhrVB9oqdRiAi5CdwwhfAGDHjwdNSbh2FoUEisRnY5rd5Zu7
aLbZXRDhGOkOChmnkBDTI/YekXcgh8PAXcNEJcpdmIfHMdegaY24wbhGle0H
Gm79DPe0aGDGryz0lg94OM5RGRJukDBw4lJvJ3BVi25TIlIEW1CeOsnX8xxD
3KxvIp2R0rDlUYsFPbdhu6VBBfAHPzkf5+GqvWNZ44okUKADV5s7spIXPjjS
1u9qQG77CRvwkjVnfU1W/9izNOn976/5kkOmrd0euJcoU+xxCvL4j/nA4dK/
kSBTqJwesaIhG8vUImBoRB7h2eABan3fWPx97qm9HWYmdfaKmfeiGd0gQ1st
46qRP9lZRxenF+uHTz/SPNOkKrD4GI/2kJ3jufUWDPArgC4UxVTTlIJ4Nebf
A9N4CheZOmX0a5QQgK9Y2EaCJDgJYyBAFwEu+mbBawHbje50YV7FrhLxhSVG
eD9SodSh7DucIeuFgixtyDKOGVkJbi+/Qe++p+KIB6ktsSzCDDAhF+ioF9iC
W/0svmxRZDnM++iQVHdfm1X2WpGL5H+IQSbxPEGL/0zdHJ/y5gkzifgeBW2d
dbqD1DMCpAzIGAli9IKbSmC75wcc/b3yOrhs7Pc7JVCWmPrm50Rl6R3kKYbF
tvin3YZiQyJrYv3srqPIGAU7aOGLBrVtoahQgyFTFfPPbecW4rmdazylt+VP
mBeHaPjwl4KWYTKK2VRwHUT8WQhdLgvEpNiBPrqKW2ke5BcNDzy2l/1OMVgU
QABeL96HuJ+yGHK2ivnRPCAS0BYvtIZJ1aSZRP9ZdHfNx3uh1r1SPRuObnJI
5csdMSzdVY2vMAdLChieWDz1Y74CSi6t3nwTOJt3MMHY3pWqkE7LvZ/YGV/t
qE1YDU4E3LIk7vsmuH6b+Syvsl/lBOjaqMCAo7mJbTpGGmLYxAkMTkjUrDtQ
9wUmcWKUOlfJbJifNGXW2vI0BO+Okl9LqAMhkaOwMIF98XgKdAbshtoIJjn3
bd26pwoNk5mwv3VAo8+bbJ/L7luspbetCJQEmZIDqkHlwvG9DTuYkVr5OgxB
KZN8OSKr6U4PrS7RDd+sS2OKprdA+TNqGQQx6WLv+Hwy3ftyyiZ/7VFus4Hc
fI8LMP/IIKlebel8uDix6uuCzgDrljT+YiuQDrMv4I4vYU55ibVwP+8kJfAM
DS1C+AVnetbgkAuHK//da06Rv6OWQtK+DTMUX89sDd0DqDx4AnebJPE7AZEc
mx+UuSar8RC16eLrAL8SLVxntZt1ESJFOnM3YVbOx+LmV0Zv01AJzIw3ykVC
Cnh8npgnYBux8ElrePegXUJ3ceF2K+Gc92y598V1ruRfF0ceH2pIxJAsZRFo
wFpFMKcerfJ6lnjkj9b7/OL4DLXuJyaRZ6f8URKCWVziXegwzBW8pOn+82y0
hJGqRSqQVMg4rxgfDVA4r7pOO99aH2lNMtX4Z4EsREKhISDb+PnkIYK0g8DX
yeyx5h4CT82JhGcXHTdUE4b1t6HR8p4yhCNdJ1xppLmrUTBn4KYn0ZI0bd9m
sdRL6YW9g+KIPJDJC3EAHQPz+x/5VjHPQ8PtdnM6N5IGEGqDe4TFAC1u8EPx
+TzfobEodMoPg2Po0+IOUTeYraw9Ns7J7RtUS3HAPG2FOLS0Dc8v03EQyQw8
yxPdMqSGxHy0UT/6SI3iYnHM5KPcacWvjNkGFmQW7z7jzBEj9HGxxhuPQ0lp
yBt1T4YTrJ4gv4xsr6ogb1xceI8IIeejUjuetorhRMLLwq9NZ4BYWBKOW9f3
cuAbaeCy9Kv00f6WXFoCZjGOT5UZps5sgi1EtBDqG5GWPp9II0eVZfvImQ/f
d7GITwDRm++uiukjHsi2I8AJqGiVsfNEuHDUyieea2KVK7/8g2srl3NFoAeM
EYmQQDBGqpNJrMAOtqfjHMVvb3Wx/2PX47MCEcSlCczWNmMtoBhvbdDYxuO7
/Y7M50Un+nX/1Ytz7tw6ledZfPCjcJKqLl8BLKzm4TL01Y56Bc+/o4JcByy5
b/jquMhKailT5CvIfwdYUlh8RjRVoH/5BQtC/0m82d35tfEPh29DwqIvNw6P
NZhDWeDr+3tdFpTE60gpkEfAc8ZVNP57qGZFXpOUaLPPusYQIWfFXbS5SPA1
VauqJhzwYLl0TnpJfv/9H62N0XFcgmgNWDiwbkX4H2en1UZQxfEbFejxI9iD
Nt0fL/PDNZ4PPBGzHzDCtenVhYTDT0igl+v2S+5Bf8wWmn5sNXH1kdEEW70t
eKNcaptnJfE2sUJM70HkUXJbe7xSlYsPsnrBmUlGtNpECx0b+ShgTinRJe1u
5C88RgoYyKUvw7Rvm0s3Oa6BN7X1xyvQK0woP4EjmonemBf+5gXEL8u5lE3F
eUkZ7Hk3xC0tbejNFEjA3TltP2gLOLeSwg83ilG0VhrqfrisLwOhSB7QKvDo
NMb44nYWDnSI5F+GmTwYwt69RNq1TPweexJJ5WBvkRPYb8nlmLIw8NsRy03M
NT0Rj5Y+KQF8TCXiiljcORa2nzxhG0k2oEt3Yu4SMW4s6zJLux2rX0/AIXP2
QTQq03l9YzzObnNKlNXiDNn/nNJhUfe6f2aZQ2DmQd4ttuwh3OAviVTm6wYb
Eb5gROGChYfsOPLETEWOqWu430I5XwOd+DvG69QY3Uyq/56skf3L0elRuKl8
gfzjBWybkCnjsXCTSe7SJPuBHbYp72KUQdkIQsITgbj3SGzSQmGuvNgkKKJW
KlPYDZoLaLZWGhm3mnKXr1FE3D6VF8Lv1OuEq/rN7+jZNAsHwiqAFepG9BaC
f/DvA4JvX2eRnJU4ivsq2O+uMJnsnbkm0+GxnnVM+qYkuUf8aCKHMdkcYm/U
y8at9YkIplW7YFQ+uRcivCIonMCs5E4D7bz19artHcOvrxvYyYyQvVxBsM7z
3GgATRo60Yo/2ZhcfLP5aN5lV30j8q6UH7lt08jO+/vSClSwix0Q4fnz3sWz
ZHtnAGIrwaGOgVI9gc/9ljvKgvPWtt3U+Roowco0UGNLu16+nqOFLytychZe
gwtTR+51sP4YT0Rh2y+zlllEUpa6UDgX/h2APbvYboRxZGzRDwsjTJVMHOJi
3ZWGY1XoDy9H5P7cGGUhp26tKIKZKt7w3tsSBFSOi7jaa7V8nKH19aAoDaPn
NwleMNvIQkjrtCCUHHAr9xoiA9P+WyxnNrgmYZ39+Z/Xdt+ADr7qDSi/C9vM
ZLeq2pp5EBUHPgb2IalOydyymR0thEetYWxUBV0u/crE8yMXSzuON7uJ2ZUo
Haq1gCLRTzngIUleEhMGwNkU4yvgSKXKKZs7E/SF5RmIffgQ5pbAewhPYd31
poFhRL/MADKrCJJ7e1lkiRGsBSnJ3L+G/jxWP/Z9gTHbWX43DKFGyuwWJ9xE
D0Na+DCY9Z1WYPEqExMzpgVRQZPtxWMPhbHEZul+CG3rxjstm9g7GJZTHw1S
PmdLyKo85IzNhAomW3tfouOzprs6HX1On8yGSrhQe0TYT0vNgfdOZfAh/MWU
P8nltE9hXk02V2DUsa7SDoqunfcGp3Q/wVXdc6gWFy6XMEv8yd64SwCIqoMY
Ozt6OH9KjKYBgPQBeAQuPSeIqbvcysDTmHGTzIrh10+9On204OnNQUadBiJJ
COIzByFkqZWa1WNhWHm+BAPntMDa2mvIYP8v9EaH+UqLmd5pdJtpJSQlMDY1
HQhJrw00ODsIFymBNSJk1x2IAVdDUD8cpGi/Y632YJ132hWq3CNCYXwms0Pt
FovuZie0BDQgpFN84EPazmnasl2LkXCSE0eeTyx90idv6yXIWY4eeajgUsQ1
YwVcMLBCnUOlzniVida5OrhHwORlsm6YhlFDo/fiS4iskWVk3hwJfGkYANkd
uSztiSXdkfcodGgfPHkrsHJxK7ZJfr3nor4wr0czwBt9+K789KFe1o4JjUNH
KgF1mM0D/eGPi9DWEbmK0HJTi8I+bExRNEr4qkDfH5MGO5iYs6MWkbbdTllg
842UIFHrKYzF1cwEw1fXGy6FuDu64G8/bhgq/68fcoxDu7ln8AjMoU8G4Pxn
R+OiKzQNUbCDCLxQeGoDuYRTKl7KT2NpWqEuCAN85MuYtVCwj4hJNPfmt6yR
KMa4Mf7tLIbduPvXFQavvlQhxVs50gFJ1JT+w1XJktRhkwSbTtDBQVoOeoKX
6pzP/pAmbAFj8X26rH2gWsqMaPs1rCc/OAFptjLC+0sIBPJGE5yZU5hh6Qta
pzvI1EQEBsUEbsKdYy4CfQGNnXwvGjF7Xkb2IcMRdCk/IqCJYc4qxBwIdvHM
MT6zF78snMDM6ytrrFz1fpfuwoKPbFmwEDxKnFl1SId+NQyTPl5aHKvGKu3e
s4xfcKIPR14FCNz5hkFfLY2iYSJL2c+HQMA8RD0aVggXD9/38nfzqGywV5FS
JTM+qAzKMhbO+V1EKihWSvzODAwaX39yLJn+3N+UiGl0ByU1E3J4NbasJSDW
jpFc5GPaxgDPF7+wuUK2ENXWeR8Oq0uV126k63a5z08WIZr0fMwo5brVpVU7
/RTc5msS+t5lQDNzdcUrbZMFl/fLkZs0H4YdFEVZaKPrexFPRZ4ADQSFY1nk
mD4GtZmbPCVYv2gLgJ2iFAtVqya/8TeYgxQmG4xkMoN4o/5X8lcIP7U1OJip
FwiCjaHgHJhLilIWUEmFZ053f3S/Nrdb0uYeEfv+9Dzgo8XQLMt9tRSlL+Z5
/pbQJMaPtwbWdZmaDG/ERu/hqGVaodubfJftJk8DDuQ+7xLJg7w9fFVPeb8d
YEnSUicvexMnQ5L2IQnpKIjTcNrOniYouKO9dUMcH9+Sj5VgQ3uymRn8f8Sx
r8qt8kTozXD4p4GqRK50OSkFAtplS1MW5/WhD1OVPGX+cI7Jc/8L3BIxaUXs
kPzb5rkNOTsFsx5LVa+oU5lEtI0915g9LYNbGfR8sxE5gtofij9vJLQq1SD2
62shemjgS9DaiKPcydduG5wCAVqNWEaw8+01Ls0D6UW7Pn1l2n8w1afxXFWP
pYnuFSehIMIC181yv6ANaP9oXbXtbnAgfcRygIl7UEReWh4M4a4EQaOQTvu/
Qxp20KUKyaQe/QU+PQ5rrpwfgfVhfGrJCK1qMfdKrpFcP6bZbiDde/7LaZdH
SYOz98fPCx6ULWafGSdap2FLen5yO9JYil1wnQIFUaeMfVM3vtIbT8bCUN4N
rte82mouLVZYqMQj0MyVYEC8TqO1qXk0P4YnopM9AcqkBFyR/y5Ejr2oWBRP
kqljJwaOxy6aIj2XarKdVEiFGaIdMA8TDdY1vzwSqUMKaFQbo3n91ASk9fKU
VxIe33nctQLWuN4twz/9fypk+BEKs6H0MT955lUNmch5e6a/0CLuigGm1YRu
U0kc+CrQNHAqHPGIY4oNUyXyhvyQQJdwmADzus+r6TzJG+wMJoe3xjdano5r
76/TEREVTWZAOk1ZlBJIjpTsLcX1O5evC0ggtXQf7wxU07XcTAzaOttEAO+e
8o2OUQ2L9b48MIV7jzzCJ+vg9DoZmpZ4qOFVecZsmKBHJTL7DOtYnSvLuzmV
qVghgKgFQwr+so4qhyllXRnIiQWESfGw2tCLlenS4bryv1Q7WB1XhoxsPyOs
O4mlLt7pSzUSIke2WsOwsAJekpF5xA/XjL8o2AkgYc5pY2MYENEkxjkix+7u
1OhZTR0SPUwS7TzmaKZrKypI0Pexc70Plb086lP+0+ccm70fDctwpXF5LjUr
lhQVN4vQrGNllY57j/+8tBznxR7jvz+VL+ZHN5lPgC8rky2zX78b5s2bctWE
wjjYodo1s6N2IYn+L2Nw/OzJSv31U+o1a1DK8wod8sp6GR5mbyH+XjYq7rh7
tdy+VOFBH40qjPKDSmB7YXjms5fLaJygXXm5Gy+2Bg741rbxkyz4QeOu8PyK
9WVhgxUPPIzAUTMKDtRiL2y0x+U2Mlq9UTh5FKSkB18evcNBbMTls5Hv7FQ6
bPCrApsuyntGNC/j2Q+LJojEFBBNO8n0QLQCMnQZXYKdVWje2cfh15mO9/mT
EpS5hixOjWnq+f8bn1Yzcm1MNnsrqovSTgmeVvov2KcNXvwYjIKR/rNlFO4q
KCwF+i8zXZmtBgTU/lkgxM04i/3p3AtY6EF6wSHTe5llQyPut6/PuFgb+Dix
jwFxwAI2UrVJC3vcBtjbVlH4vgpXn4kQoNPZbH6pds9S4CVR6Nki+aqq5e10
srQPbWSXHSQuxgZndaBWYwIdpIhfcFgTqYZsbXW5mQX2DsUud8/pvRGamOBc
bHgrbL6Dr9iZhxh5IpNG1Lz/detOYhJhlb7qeDevmW82c4ADSurCF5nZpmW3
AoU62x58oeVT5WgSRf9e8kerXqWnGa7XcnSjc/J/CKPox0PMtNMsHEfzb/4G
15pm0HZi0x2msKOgoIVgjiRom10ofD2FMQqpy7Ra3fG5f02LhQH2H7s3qxVS
Zd8+xBfx378ZoeWC1rf4m5npH/0l/17Lnz+mmA+itznDWrtxnJDuOYhlBu+3
qGcKKpF+0KNjfPTaimBLLYQFnYP0qwIRuzwbxyTNOwksShqUP6yctYG7Q7uC
mmxDEGj/MHwU8NW2lc7kR8/S7f0FoIlQCx6eYFQpdAtomw0p5fJRhMtkKRvA
KP5M3XaC5HiM+2+Nj7HANsiITKYu1L++u4GIb5nyZcindvxW8mjjfEkagj3I
6OAYdbVLOCwSgEC8yuBEDd9EaGz7gWGQjNNSgaBICfk+qj1WNOi7aApPsp8k
4DrzY1tEtrnp767cghFO/6EW8+F9h6dT1FqOa5undx/qpW+4DY+YZSkB6C3S
ggx/+tWPwmOZ65jn55a/zfJ1OzTCjacXDneYDmiLl7s7kkXqWG9BFAXZqQ8W
79m4duaM2Wb8GWTdJBKus3OND2yROKd2KD3LWa10eQ255iZBJUSB+Ut9a5MG
cOd/9Fa+j+/I54Z2JQyUjO+sHtkJnGEs+YuJ3LmSRYaLAve8fjSRpTc441cm
2psP110K0jqkmu0Ae4QSuKQzlAuHN7p+byu0fnwVqSVqkH4cgHZJtNN9E2bX
Z/HBvJti6wXSiV9jqXXyMyy+dS8BO/fySPjYv4kvLL2u5VNqQrbEL+AGOmMR
ueOwyvnzlGOhtFVHXYt/HPRUagyk26EQNzDomObbpYC+KirXq5RhuK6b29no
XpVy/HXtGXyvU26/abKtW/SIJij/CJAnnF6KvR6ax9/dPOxdvoJStWPpUNot
LhVvAi0KMgte/w6Y8Z0fqjXjFUN5p/+ZeYMHkPA/ginTA6ZhaO5NGx8EKGyw
SGuitRcWP2EK8zHokHFSCm8YCXveC995OCL925WD2lvO3k75J/lZqyLMmT/3
5Ln9whdq2rhbtcMnKMEmtF8WZoWocxzaz+FOZF9/4iYks6uGxpqSPi6CdjFh
cgIeD4hFObpRIvNbzte/vvfdGWWGVaMUiwDk2EUb6SqPs8mJ+kUbwNThpDPt
UvzrKGv8pnsdCCVYUX8APksDSiPeGD+fU3P5FOiv1KPOc4cAA5cjztI9WRB1
TsGBnyrewg02IIfZUcg3S+ep0bq0ul1ffilGap1qTd6cPcI0uYOXIH5zVjJ7
fP2TJ6iZHEqpTGZgabhvjEqxQvJ8javYN83QGj95TBPyhHmZnSSIxYwP26op
1Xp8bmCWE+X9oifTKpXNhnCOPD/PaB0btaV3piOsfBp58hKP6TWelSVwY/Ic
eOBl97Sd+sVgrJPU/vOJOH4qSMgwfDuSKjp+RK63pZwf/dwH4hkP9YXbDWuQ
3FAAUWvY/1emLrMU2UjJNcroIiWYDnIDTYbA5hNFTsH9KDzidZlqj0zqu9Oq
2pJbuA7jQOgj57nzvV93CHkc5KJD63EMjowTvJXXgTT1JhepOXVBtD8VNTwH
pac9V5a5Rv0e1LYv8FNFnFcx5E9V/T+GY8lqWggVAlouu/M4xRATsfw/MXa9
pCfS6MJ3ZmB5OU1ot95WrdNsYuLb0h4tVuzgbRGFLI5g1trBYQ1FO/+hF96b
DDvfPOpj+0SpSjLnVFJVMXwjiCPWpzgZiOlIi0KN1X/+RLEPJOJ2aDqC3MQm
l53GuNfNvHFAkxwZOPTF4EskstV22J0o/SrQcPnvfm0L+cDLcqMtkuruxr3r
k/OAv3bt0EKjVmtCxa0EotYZiS0KUGxZmiA8Kqt5Nbv9mhHkoahT8WwKwiku
rUWOYE7C+HtZNMRaayKZw5La5L5ljI3ys5gna1SEAb5lo2MkfoqwGuqsJCEC
aM/0ogiGgF0q0m5wJMFpzT3WsaX2umAG1MeMFfOBSY4wdme17lfuwGvsFHKP
6AHhQgRnKREUuYX7fAZ4geq/OfKNaNqhYty9jlTMl8zVhHul6I4qRggSQAN+
/1xrEgc11wgIMiNQCEipxPfi1eIxCKn2MAP0hB/4UmNqp+B3F2vH9H1+Djxe
xFzvhrAVlPee0wGBrTAH5AIdhpLknoxirE3mCHr1d/B9RMtMhrvhWvZOTA7M
Rve8o+9hgbJ3vjj5lzQz4eE2w5A2I6CnmBzX1QIZaXThBBdo6K+shAM+YEn5
q1Ci0glrj7R2pOtDO9WLG0rjEbeZFjydtLDlC0eHWB4h0Giz6wOLoHM8ZoxN
SQYVQGbOrCqISo4+ZHzQinrhW5r6xiHE/mMxL/kmTCO4g0s5Ks6N6CxXnnR4
038/tYE3BnhbOELg0EgJAeqo3SbFAa45PJqgRp6hhoNf8qEdmR1ZaPUa/Riy
nAMUZNodbkZ8MEHqm+PCsm//QdF0fp2WHQd6Z87gm70xO222vlCmJ5vkekz7
ZkvEwLCWkNngXsutrhJf8Tnyub2NF05/ROh/axECqhzJApUTbXfA36XM9bJk
hc0680Uh1qVRCKd60bGJ9aD7Zgd5m50SbmxqrhVpeB6rIdlkJTSlt5UEUCW/
7LVDJHYZSN994n3JuUJmhOfIzfSpgm7Nks3Kvee4i/dGdiGwm7bD5eUfJObo
wQDv48OFHLg2o1HQvGb0ykk/mbwUdaa1cEX0s+odVkb/ixnfaGtn4icsnl7E
CzErozO1Bvbpsq8WxZ1cE/B6EC2kv0Jinb+PC254X/kMRX+RCadSRrU3AEdh
++HZ4K/VqDBHQ9pQQUoZbotCYIqP2xJWJP19uOJr32IRfAo2cTWeoI1/W8L6
9ZMIrgfo6yw8HuO+rE3JBOKqGDQy95TdQyLNH3G3kHQGo+V1HrK6tPX7jvWR
v4hUyAAim8mR+dBHjOQJKje/YD2Za74wAffQM3v18qmp1WXnBp9JTF0Xb5WV
ax/JKZ87YnVLfSHUktWeO9oaLWZUumbKyuGbA7R9UzitAReQuUYMHFLdD4WM
B+WfnF1I5mIFSw1ALia9ZrokltCXmDis8VMk43UUMGcDMvBgLL/acpoRVKji
aUZWZwj0JXjdX5s/Z1IEpMKPYrMslLgKHJbOm2EEYUikfX0I/HulNiMpe8ou
y8JoqTrsJIaTbYUnTcWyy630URytCvEPD3rQQXm3alkJa1e36ijbdb9/dNcT
KFIc1b/qZwtOMWEvsS5bCCzeg0b6HEH9Ufc5GdR3fA0FWw+fg5azazpll1z+
Gvc+ww6BJT91VTlh8KNnLSCouSW6WAel350vwASw/EX7kokBz1EqHf/PUgtw
rmn3UDsBz2q7XXd1Havrm/6Xl69OFj5NZFraqYlGQFgxiLoTurtPvUZIopT8
mgMyYUJik5heVIOiSBwyn3CwFryxH34KF1oSipdr+wyHtaBE13zDgPu3YXjs
KMAL6Vy76A+Yn7V6ZpjnewjSy6TN2nVw6f2tQSNapogN7F8h8z4dE793B02H
9dVwk2Wk2Uij5UeXsU114aoJn6EIIWhqO55AIz4Ib4+22xp54XJAvBPLdDcj
sK0hP1gV9jedfnUIYTGV+DoXZg6P4csNJGLk+UBcaUJkAjOJSh0D+1X1g44U
iwqf/7H/LIibZLalCGWYVzfIwLtM7z9Fi8lAI7cNfSAvcPxoeb6NvUcwGutD
GkqCgJz/JZrSHhnsF3XTqj6Dk/HvqNizHdpY/xfNkHDR+DpQs9k4XPHBXhqe
Pg01RKOS7AP4As+aUvRkX1eM6ExnjWFjuXHmvblHudevvF9dzhbdZaCf7f7r
HHdAFkt5eAl0JnI7GOhzhvn9bCTXy5OmyXwRIm18jCBE6PX9/cmxAihZvhcu
MuHLCn6iB5g+M70ARo2+rATHHI/fYTwl4s39E40CyDCiQRzaFfQNMHJkR+Ji
DZMqTQWyIEBFUKOsaKi4GsMajnucoUxpQsMrbNZseMVZ2i0R58srhcVBQZO0
1TSkT6KSJ8bqv+luj8+3mvtDXP8N4MpGmOXr51iVb5xKFKo0s25481w0Rfec
1m7zL0mjZthNqgtLM6bUz7nsyPpsoo/C18OKBpYc223iNgQ5e4TqRSoj2aZK
/WJYCL3XUn4dqsq2B+ZwW6GVtFZor0UcGFm9SJ1mApuJ1uRs5rWVp5OsDPeD
+jPNbCUOI57e2i0QyHofnmEZu/HFJquHZKtWFI82qxCslzL5pCXZ6Mtn3T4a
nMFupsbeYZeFevThfookd4gOLqutZjm7dn+97O41Nhug5Xog9x60+iqGVq7M
hjGj5O0QGPsL3kmdqmhYk98mZMUsn5NtZE5cG2yQ1oGO7AMJAqC9DAKaf/kr
RIjZvZdEh4EQDd37i7HpXYotNOJFdpUlr1l4OiO3+RdHujYsDDlO965OttLw
4FR0VJJBCl+eBwxC2I3331Nl2/2LkxbPV284DW4lTh/j40eo7ydNP6fCv3H2
PGQeaDJCu1x5AHAbCuDGuRAvv8KxMyq5ERn49priONmnfpDaeXv7Z8/xVHai
yxAyjanfzAAX1Qki1XjeMRxwPQ5d3FOn9IQAFTtkbJnPtUq2P7yLcOA/SA/i
5iTAz9pJW7HYfx5/Lc+69cYbgbRy+tqkyaiqvVuPhCRvySB/pKRha7Z/jRK8
7AuFx0J1Yl4X2L+dS6llE2dmEMTQ1gazA1Vo4xb2YLw0PDl5j6A169rxUm6n
l/zJa6NZ76VrECBbpTKpGcboYxECelexllNkCSwS5rm9OS37oxylPKd+V4T9
CLS6RezpEFjLPCJtcSNIup+/znHkWtjMw6LralWvCFVXngT8UQ==

`pragma protect end_protected
