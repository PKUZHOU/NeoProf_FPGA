// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
yCn+fcT9cMACczN8BMvh4X0+7vKRSMwYLIrulefXcGsAi/b/7Nqa3nSIEhgobv1MyAj8rVxbAI8q
bDXW8ILPtukONdeER6WZXRLigLWGbZU4wKf0d1AzL2RioRLPrPlN21p3BjchFOJCoxRouvJ3v7IM
A8Oawqt+pxEdb/BPwoSQ1NASaMDbBJeGnWtYEXCvk9/ZBH+10ouKeqGdLAUREZz9AebIlxGP9+lf
1IKuw9haUZyx1HYBRs2wfVYgyCj7O/vSVp3zFZtCa2Vj7848HIRhdPUMQDDED43kHvxpJy+J+msk
FLyPZaEAdIl/EDArHHK35yV+xr9JyFIMoSB+cg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 29360)
ylLDVardinssIZaZxWwwo4ToLidG9aw5mED/MQ5OCDCir3elao6ohNknd0QE+/iuYtw3oULw6tWn
AbtPMhr0m27Jpz0sh1Rtntoo0MZdmsJuv/fqRXcTrvKtBFV1kz700dWyl8YKNp39VryGlhJ57OBI
DpE30ckae9UnXQfHpbJvNsSg7Q63peg/UwROhlNW8NFyX4UBqK6Bj1TGv8ISF3MWv0+dOZdQx+Qf
Z8FMBvQc0FVvgiptlH7w9QOeCEZeZrNYqV6wg/ql8anQNffYoVS+lN9X1gBFawq75iDNoKKdGywG
8o/tYj5rbE6pld0WdPCej37qGXxhUytwwlDQT5eDkaYut7GiaTBgDoC0TsZfV+RidAsmssDbPJlS
bnvPN6VUqhhAaN9SzZ0wxZCf2R/APOdTngHh2c5kwmnlGCt4Bfr0SD283bZpvFOjE36H0nI1bxka
/2UpWNPSk0ty79yv78L79QR0XXgOAGrMx+xI5TV2TXWVKjdJSuO5ePHYrA/TsImFJEUsKeZvGK3j
0Rginovm4RbI+y06avY7vOE9pNU6Xy9zeduzJQom4pUSPWhwpOTfHxbmsaugavODmUFSAonEAXug
7PMdm3IROipSrGV2E1eQVfFDpB1txDcs5bAhCIsb6iIK6sCNKkegzhw43y5SXvKaS+eVJj0fiMYV
0efr64Z3arXchIS9os6hGPLOmx3DSID2Oggrvk/QSSq9L/ynpv1ggziNaQdhaKDCTv+FKNAulU0D
JloFCiETB1fMIxuHGw0I006yLb9TB4uhY7C+IDnyXFYH+z4Ggo4GPUVddqg8KdkxqJB+aXSUzvym
b3BT2WJTYO9Igy6GU7yRBN4gXBMyxnov5EE5XNmskXbiSAcr67zJ8CXxCTZOUk8RPUcizs7iZLcJ
DndUPQFjjqDTc5sBwk+2F1Dqrd8cIuT5eJTBb5ugzDDBVpAFjusndlSAHjFEuxJlXFFu07Tucv5N
5va0J1R231mZc7hiDVOKnjFmLKguD85EyakqUURwXBjw3cvf6ylAh/mPWQbd1NodYoikKq9a9jvQ
q8Qc6k2hXIadX8wmyuRQBVkrE4vbwPPda8Be+kTCoeSP1DthjZJA0mpUwyXskLugojaiKdt18eT7
NgZBIO4ZYdbPoAFNV9KxnmdlNWLzBQhEP0gJnBDP7Cr5fRXvjZTF8bjcG3oW+SwQMxMd86QccQKW
m/9Hnfdvyrh4snKyZj0vDZBoyJ2HoCMPLxYAIyW2M/y3Elo5Md5jrtdt6UuVC1D1gIeozyIMQ9Io
vkhoFh3cdHLMyGpdYqec9E2wAxGO67HmIGkmbKbrfokIZmkHoTzo2sKXyqAI/wsK4tZE/lliv3Yh
oQwLdYX8Y37aTAcUV5Y0xVvpWRfzlWVjcXw1lBrW21lqFy9k+m7KQFFROiNKwwTxwlsU3DYHuMUj
8DP/18UT7R9E1ddoENtqcxi9Bj8AsfvNQSsZCHZBUx7Pk1eI4/mWh0t94GYHAdUoDa1rankAqU4d
FT2vMqY0JPCg96whIHFs5J3Vh5ya/ZZUiaTF/Bg2T3RrDQyn38as39GAYMgNX5WOxe4gsXHnPJ55
1/BFosgMCJkrbhV6ZtDAqh/1bouK7TeQDnAvooJWbGzgRzM/AYxbFXURN8MJp/iiqykywGciFdiZ
wv6DfmoLkFZHdtxP4ucvtPeXxqYt4K8OZESmR+051ZV/Jl/BoJrIP7eXxlZCjnVKwzbVpalwP5e7
/ubrwMXQQ4Qhulwbxo3y3TQFEvXeEpsPymhgwt10JnS/IdTnxFBii9LfKqwc2m/XERowODhTQYRS
/w4yYT5pJJPfA62HL4l1rPAMnjSRSnrFOyndJwgmE2WY69RjuiIaG0FC1oBttXauLi1EGSpGT7R9
isKBZxNqZqJpBZfnkVUdAuumtGyq46nagHzleEtsIPwVtqIh++QQiiMNChQVkala5Prb56bV21Vw
KDNgum2EXVroB35/4KVFnMWX1WiGs5xO7b/Famg4UFmIEQB+Oq8mRDINXm9wTGNNJwBinw1nfE4d
5Rzcs/tgL4st7Ytcwxhr52pGpOOjHw4g6pA3N0QDL57ysU1eJgQ5PgWncdnq83K1QH8KyqMw1+GA
QxCOvYJvXBV4N/HK5rsfI84hcY+yO+th0RzS2Q5ojcghNWUU2y4UMnnJA4V/oPEcgsfqMg1FOS/K
6twq9X/loYCAioFVH1k+3JljkNVNrXv73XunjERoxrmBXcx1Ph5DGHIRyRnCZlPIh/4MgDbRSDI9
0nI/xCuisXzhAtwWPrCkda9F6iPdEu1bpjMJi3sIybGWmSx53NoVyQOSppE4U/PDT18v7SLxjVfo
i86yjy43TUOwu3b6NJSuMab8Pqx//44VTS/ATizVDmytW/40zEUx9bMZVUPsf9fzhLCdcN0DWc1n
XPRWL7iGSUVwYBTczB+wKEffrHpMjm+S8qO8Wk1QKvQvtC0fmy1rE4y7dVSuRAuCVSuZJed7tERa
rcM+fvoq6HXHvfYXUHQbptVvU1WE8e4CCU59OeF+eR1YI4rEUnZrz7UPB2fc7lUfRAnuBzeG6Jfx
A0kfPo/ntlYXDOppd/EQb+ak76SwvkqpYhtjMPLOd2GeWF7Q5mRfc3Xn4rMIMr5XY15Wbh4ITfhz
5FAKlkVvvbm8sc6dF9842C30Z9W26P7bPd2xs8dyEj1QI7HuVo1WaGZwP0KL5ch4V7iJF074ME87
bz/q/EiMP63YhyVzdlF34MtL5RGyy01cDAdQmxQqU/BkK4x6wEl6hHyc3f/HtOw5+UZhbJggp3/h
dPVuvxFvhyYAuxOWp97/UWPFrtTlRtq7Z6ygh4awA/w7M/SA3viauSFIjLDK3+lSJy5bXtM4QUUV
R/BWfp+y3Kv779lnAK8PaPMpeHZ+UM1NQtFjraF40yFJ0xQt5nPHIgh6UQcPu396J2chi3+nE6Gc
4Afd4skQ/C76gnyU8vqq34fJ7WFlWc297NXx9eeNvz1e9xcWeAtK4gB3Mh3ihO0GqLBi7yCWs8Jl
qZBvB/DH8PnbOIyzUX9mPqqDTBLezaA05z7ngN46pcNgW3e9vuVpK8+JhP2VaN1xdfi/+DR+mvb+
9sg+s7M1PKg4LOMqYn4/6bRatOAbHPaYx/wBkb9UQfks5xXUxhI9yh6ZzRaD8ZJJdrmPtGhySTw4
8Jsc9FKCMIMd5P44+oWI5jBieB8CVEOFK8ST8F7f3DLwSC+A86wDPR5CzJ3NG/yslli647hs+5Xi
0Qz77uuS5UHNEC1mcN07m8fDWeqribQwVS8f17RC32Kd8Nvogm6iPAmmggijLDfk7qWnY8X/slzk
ABepCma6tQ7x1Pn427pTF/GvTmXidLgdUjehHHXxjDXL0r+7ok+zP4s3TX5rhBd0Hr5hUThmB+5E
mgjejb0kQ75WhXHDpeKPdnGDIdcjbs7ZVwP8iMDrmUqtM8aosdxkBiCq6UD9NduTVcORPs+1N9Sz
VAiRUFrqeVbKfQlGzjDtvXrYjhyqLKz2aS6DOWkyK2Up1J9kJy4bV8FxX/ybIIkY19JjoYWK+p41
bObQlYt1/j7ANVhMp99wznkay0fPuC+H65XAVv14jK7TBJ8bNDttU63PSIeBExkvoBn/p1lCI1Yf
IFtm5mkRtBz2I86ep7tl0T70OBIuqssA+GDN2EUPegGqgAJtGH1Y8Frb+AFbgUM5eXHLXmhAsh4I
febmd/rlkpaYWM0BrsGkPTrOMbyAdaOaOaVVUDJWv97bujqkyS47bDuODVqFPTQxWqxwp0A0yKSd
0UXoTPiQD0l75VS6GkYvxyjkk94pPCinHj1yc4G4PstSEA88A1o4eTcvjw2ytv8HeDt5nCJ2snoP
vFLmssD5wZ9bDqYsZ8QHiwtMMLMlaH5BUp8dJXF9W/6ZadkVXAxdh9p7oUcFgoBnbc9Yf2sppqAU
6Nx8+BbKp38ik1+Xg+iFGOOF2TstWBe2NuVEzHbgHKLvpHetcpAQqQZ2bXrC3UUWjEamRiekyHAm
9Z1wKF6tcL7iZ5eQFKKFSNo9+N/XBzM2J/nRKR6h2voY2nwMpGXZNUXJZccl8glAioAxg21R5wwt
+fZvbj9xRna1YqwfQ6oDkVQidLpc0wfURTPPTzrg+ABhEjcuuLBuPOBguWqagQ5SGDzHX/trH6g3
g1Lmo5HqH6SUsmf8DriYTyWWzzdqwG3Xgkyb/YY+FJS4oGiohzkP9z5BJA4Cp5TqZFLyq/goFCnv
diEBf1cljccSlGbjpxd0d9Tcy/ao/+oTPK3tIRGxrXYy6TAlkzUg+jTU4Ipt1eisBKKE0qeNGOo3
PQRor/fXWAmiNswzTnBp+2XrgRImEH7Fat3+3b343Xo23HCt2AarfYVHPlrTxTNpiIChw7ZyONHf
AjceVATIuTOkCMg6mZgpzNDIaN4vvXqIJ9Ylnt9roglki4Dt4UJYzc6gdLapduaRJPdYUQGbLRn4
39EtotuTfoHuVfBV7/0DZekt8ydJL52n+kair/FmuCC5aUT2dQv50pk4UKLWmYzCbkbeh2VZOSJ8
T2RDrfF7t3i0nEQVGpwzYEnm+1l7GbfrWIJwF/p0dImlpJkunHapv3t/othDtgg719utTsQaRRC9
8/XCWzo7/Yy98KFHr7goXGi9mgsNR81k1crG+X0CGn3Rs9Bs/zQ221DAjx19ptDO6Bk+HsXAGZi+
eBRCuwfglHieres2YCmA6BoBsDxyd6vPi1LS5+rP67kiihYjpqBlwSeg8s8xISj/Q7waLlGvl4dN
F9+Jdj2fyB5LylYIBXEJdw6zqBMDIrohRr9O73F4Q4fA4eF/xpwrV6StSBjcsltYfMUX5CVgsaA6
NRjIAeNuoiT//74OJQDJEYIOnyRonBgm2j87CMcOhhYMOXNUDEX0h64ZQY0+avpKBQ+Gl7QUGrMt
sdkthseXPV9hVt4xr/5SqVxfnD5qFSKjZVMK0Dc0eYKd36/xuwFeOg5daQMtYXlQKfwA4z5kspp0
TjnxhA5VQoEPYL1vNG2T1SSfZ+zkCyxh9QJ1Fr/+5uJd+m/noJ3/C7FiSbOSnTtqK322iv1BDkB1
6B4zJZ9p9yKUFzMG0VkryaMjr8qyGQoQP2sps/FGIr2TnYj9dElq0iIri29AQ72PabFIQXz+EReX
7KbyQ3N2hCFpk+RzCCmEI6tzqxuCuXQhShQ53hABZB86ZYjf3+ZgWRGjdj3B/92FU0IlGRlcm2lp
mYduUNUX2V0CYjmvAM7ips/k7g1eyzQXumxAgzf5OH+WfC7qMBgx3d8hKqR2UIXtTp1O8ChsIgZN
nr/IZTE18HuhCP6DiSVEw+QO3HZXxYFpqvEz9QlRvCh9YMBRZBNSUojjP5izEoFtiXPEY/MHl7ZQ
/y9J4iDo5XPbtuSJxLeIsckfLIgTlUNZXW+eqn2BXn+SXBMdtd+Urt0/q5EH4gxCZQOS1K3Xn5f3
JvXLlhJ5IZwEOPqCNPplxmf33tBKWPkzkvE6Nk+JibJXoRT06lUxUkCjsXIdF9gCQCID3amN3MV6
0yxxHBeEQvZQ0ua8Zv36Nl7e0UCowqZ0z7Msgwmkclf98UaoyYLp+LgiDr2bWFSQGpNNha5I6ahL
pb874JlMSZhc5MniQzOizTVOgdaDJlmG3rFXtyU4UHNfW5HRVczLLma605yy+vci8h2Z+KpHvhKB
gcQ3/XUWMMKZEKFFATywdBRrw6x5g2Uz9jdoF1ie0CsEXKjOxtO5vjgriSvN2hfyUzZT/Jggx5dz
IfZ9H1lo+f35hcTyGxoKxWRlb8UUVy2yga1TGPHGFyi4Kj8fyFIKjHhbuUm5EVnxzmii63NXEYet
Ioj0vOMLruwghjSiWf8FB+RHnur+OpDTgME1Rs+3yQxus6MCwNONViYicyb66FYghWEq/H8Lhw5t
hv5qy9gdJXfsWV+KqNcLpvnPI8TdFI7EZZkk1zqv3t2FnMveh7zOVgrTkNvcViTCsaZmmtyqTE02
WREgoaGY+ncMSUPFkXCIOlotMi8/BO1mEFkPqL1KDgaeMbR3AYw16L1H2IkSON59SiG8NDUzehAy
GlXtir4MDaxKf9pEdKFPN/vVhfqit0J4lZbQb4FA+d6o/GrNHNt5a6QmpBaJBPTz/1rv0d1JT1ex
/a75t4Yd0IHQr0KXFD8u8IAMc7VUJ2A15e1BN737eKh0VDGji1hVMx/wsKhJcTycr1KOEzBIvzlO
1b6xWdpfNDcxODNLZ//OMzXMdeq0Nxp2v4gZmYPIpzZ6sGjgd9v0ZOwHm+YIVgloBNu180jcOQ1k
R+UARxPFWWoKeiodAiiPdNr6kp9XHrTb7Q4J0d4qsdB950svPf0QqbBfXm+EB/Ix+thmTJuWbIOu
M5G4eQ5WZqbdpBza73C/D5PL/G2mNISpLJL4HU/0A8u2H9TU+5gHqEoehhm+dl+YTOEFKERX1eiI
I5LncihX6ii459E9c0GDRLk5vfXN+Oj0t50nBH8qS222Xj5O4KexRq8J5rHW5/unYw3bpwZtFXM3
sCR5oqNOIeDF08YkIBn+SuVDlg6VRv9laZwMe/RP1/40kbLlt8zxd3Q3NSEj2HGNo3r6vtRjwVsd
xHDZwq3h7oof08NsZpXGSsUUZa8FYdBXbd8CyUgW7kf20/zLNLNxrF7mNp3BDzDa487QurNlcz6e
f5dSGr/+zAghqFrmqg2a0pHAenZ3wgmPcd+21bYqF4p4g3SoolmnL02tIxdQ/NrPHkL0T1On2PvQ
i9zJBukMvase4Y/R1cVDrPmZaqrd4vyjxX7PPZEaDmTS0sutW9ENRfYzBvKmjq2TghsBmz0ALPdE
yzq8JMUqY3XJjyt+FvNUadttfFLpKjaCSDhxOD3poLc42/MQP7jr3uYHXpPZpgr86q1Qi9Z+Hg/l
oWomLdCjJDmp9CPbQcd6RyAv+zoSt3Rt7D5luNomh/oen3qpAk332iFPOsDLJqh4w07rIBOOrmFO
bzfDuSHLIsB8jLPmf4Iu+1wYUdktLQJWUHz0KE+07RTkuVgefnXCnRXguiyLp+vg1qpt6a/BGSE7
98Cr5rzq0BNwqQnTohZ1yodHvQHWvwEnutm+IpCLow1n2/GGyeeA1mrPZrH3Aru3hBr1eQluko3g
HZQsLRg70CpI49e3Ea3TwNMuEU0r6RbnfuRQFijaMaco58plEXaSyc0OYFgANaDVU3FRTTQ95xFG
9ApIjfN5yD0kMf/aM6sEKc441a6UJWtnpkzWbMssvlcCCzYulNsV8mpFwqHXB6ti/2ZAABeMTMk1
GeoT6vxW2f0HAwDlGIFeX8Xno4yD7ZRgvgq1wvRcJXTW9SLaD5Syi+/uTl+3KY8YyOyqUAUZyf79
LtEk/WPHY4jPuO4ijQjbWOl3JjUV3Sbl3dV9Po4+IhEWwBzLNDtoOek/8TL1CM5aUZqDmTELSL17
oEfbjVXX/+aBRLVbZ+OIkdcBJlTfyFDKgD0zn3YeuQdkIYIzfRYrmgZAt+YO2lFpgTIp/dGu0OYK
ms9f0iiRuVzsHbgsF2rrMh3cuX/uzoMzkfv4LkQNVMiaifRX7JwuruAgXeCWp9y6LvknhxGo3o6L
Og7/YaiR1lXoiFdipM3KQxUhmFgNpFark4Rr60C0549iVpSHzW/QtoS7qrw0tUFEG6+LwGh3J0w9
cX3c1bYJSjHrt+ccupUdgaOFZRd+Dda+KYKtD0Ql62/PABn7B9573UaORGeIRrq3CzKQYxiSMbFs
r3fBByXN5M5VDIHZbnoRWcf/lgOVpSNuJe8C1DUbNXsi8TGSnhMC8ErX5yLi5PJo4KG4fsdHuiUh
4i1Up4co79+FMs+EXNE1UE9/ZW3zTAgAoSeMxNmzY5U0T0CuPF6dH3GZ1SlqZeV/mFhF9aqQ/8Bc
6hVrTH3GAMvrWYLyqfRaepScFspOcKI19L00TRKjUhvoQM/LFdWWUSXfDCifiijWharMQxAmcYFj
usvJFqPn3KBB8WXG60BsCVK8jPvT6A3eLMdXelvSYvR+L5Hjbgf347/22B++HWyMAgWf41ZnydC2
pfuKK47MW6WEQLWUWAmipX19CdHcA9jFair/tXUx9oFL4odDPHZW9f/WNvB8LZ0NBVI6v8CTb6iY
d00dDPPBm2SYH7uOnkMqvOagV/+C3vY8G9nAglPxsvdF0ddLgw73UgCISBijeG3s5dWcGf2z1H7t
U7dgU+MV9izYvEQXw06kM7/YR7Sfhk9JJ+7R45D/b4ifcQehvJhKGoQXehTDZyi3Kq2ozxGTYpmf
UJPJjzikeNwBHfkvkcJu9zV8RjfVnDPIFxmXLiqciRi/GEAlrxyYllMF2zTRkLJGohXxBbPrEdek
5jgvYgV2MfwL0qcUk6gyM/RUPKqmLBSlb2ncuKl7PQf8DXGR2Q70FC0dbHYx4dycUaYI9eGcx8oW
QbnbGQ/STzaGNc79hAdKGfQL/dv9U/h7AUqulA1DUcpOXh1RhkL7peXdkJ3pLC51Qp0daLaR0cml
YDrSSZ4JYT/ckSCZBXSoHFJ6LTu37k85CHFbZyA0leRVN9ChTEZCLCUCR8g2NOO+N3MtorGok7QA
FL+AklQgg+RumCVXRN98q9mtAWXXapXk3Y6yt2xo7zNJnPnTvlQcDuXxgbTKgwEabFPABJMjUd51
mJKDVgQ5CVNeylZogY60zJ5Ju7GR+znByfh88Yj3z0KaH3wnYuem3qDcZn0r9V6cf1UQkEKKBnRN
FLQkNp2828QQFo/HP5UVSbXF5NajBW78lDkgMT+CL6kX0dOu3Nyo6JBjrsIKcJ5Lf8/At8pUC+b2
CJCJwVmlzbZJu/1Sfz4mmmsZTVC2m0yOKb/crTY9jwMNWtChQRaRoYGl+0ndxGMchuwDY6sHA+tp
Xcdv6F9gLz8dyoMs0nA7vU/4TjHAeNAc7MvlHkkL9ZJ26XgDTCQsLqs4CMn/w7h9wOAmQzHWR59W
mX4Y18fGTUJwejug7h/b6D+qjQQnn+XJueSHv54whYEwHzWmKUlqXscVWlC3HgKO006pHCxpwR4l
2lP8mjoxAwVuLdlK/D+8C3xqTrRY0Fe3mK0Cv29eetXbTarnKwqsRVkpB/xysAvqauAgLO1zRqry
xubjz1r0fDf4nmTsY4c/DrkQqCZQ6mugXmiEltGTkEuLqfmlUvrOlzFxHwvLteo91Q4TPIIiEYir
ak4oCxGnh2BkK7vbJ0yxHugfUMQYhIAfcwWI/iBU7fZo/2cYkMlLREfmY5tM7ar68AzCAU5GFRFA
ybq+X7ncnXgfeYZQlgi4LX8UqX2gfgRFPEf/+v+uQmywHvok9beQm8XFx/G4R3EregP3uiNYI3yp
NsPOkBmcnENSUy5wj7ji3wMgSHOTBnKZvL5NBzKv7/0Kd1Vh/gAjhc/gpmOpOjG9dZtfNJjo22DG
2LbQNRbeDnj0gs4tL+l8lwznLyr+HAHNaYjxrmaiqgb2BQCMILBAbnxt3s8yZU1O8YJPlpZSFfKn
x63SMc5B6PGLWesuDiLat6TFfFM+Lhc0hlv+jWKMwYinOVAtLe/x4Pt8OiQp9K5Ff/6KJwdnkmdu
BUDjaux3twjmVPRlfVB8xMKEVVs8NjDNIEDgfE8UvULLG4JXSAj1nK0yjNzANd+jdSHnI1bftnBP
6qpfOESwdWPYCCa5ZaZ3tukSj9IeqL5YdMkp335TNHjIFsPXtOIr2908hwWZF8dSIBgiN/uyvd9O
h4CmaCJ4zSCF6MuLJUaeGuFlzshhNEnU4N6q0AJvot6fqNodREGyAUr5wAB7t8nCru+SrGiLZwLL
QKnoeOwxvNv+QlKFfPBV4rJeCcnWMn7+qADDcScxqODpHseKPHrL6RsRqzrw6o620cWuLhFze35h
COpjI/ru+uZ6eISjDC67KhsmcBy0I4V7B+/t0qf87qSqL5/x8wWdO1V6H3Nkd3rLCE1MK7J72hPk
nGyhRpGyVf2EGC9tX5/1NskA/16yJnWuVLLynWFREJG1l30ps01liesoKJ1RKYznISw9tRubGnAc
Sk4VX87f/NnlLjGlqq+IsPKzV9HcIm+9VaX9eyFHimGoxnyG/v+wnJRiPqc4W+LX2RuabiUfHiR0
W1VVOIw0rVRaLcQaoSbYDyIpvhUfB4HLSh6PTHyesX0ECZwsQ1vmjsPamA5PIRTCjueMDXzU7s0U
ImbU5Q+8TCRx2AnIPNGT8398IdQ2OpaXffK7HidDXdmYMtI+OtE+5VRZOUgoyOdEp3ZR5pVjGxEh
j9R/mg5IvgSQ5QbtrnAlPDIb11jJra7JN4yqtiaNN/h74HBPqLMJ6UdZqZ0dkioMfjUV5kvkHeNa
Uhpb80i1DmkRLZcY3LcqH4D64HrXVinTIBtfr0+5vwEAwmMnRyJtdVizdRMxuK1ltPSYIrGTbgjE
EePCGLwBKL64VUTr2r+R8qk30o9bc1GW468KoHIuYbbvpd87PCWP9zuaZzN3APyMFwWNAgyntggf
JZlhpKLN2cCgZ5g7d1ulckRH8jZlMIO0/Dsvx6mYkCmMOs+PKn9when8mnnXgzGxZQeB/bjqHSVW
NEJGKrr/L2oCS93Kvt6sMWlqH+jsaKmBHiCmi/HMflQt3luDWAGq/HDlW/Eb9pE1lEuq8Wx/lDsF
Ur5WtZ0sb2nweLot6GBL+MMa6cA2NFxNfP7YmxGbTUltFVpK/0p4VJLVij0EWDmazIOwPxSBEfpj
V/xcAUsuXFUhir0xGakPQ81sFvmw+Vk/3B6z4YBGTc9jUYHg4qgNlWcWRt8MnsXJnqWQ/3mgpUAY
OkB7HNUYeIksZI9hml0xOzYKQ9jeX++1cVQP+pH5cwdBy3y5Vj3RbICO/NU8xOIX0f+hrdw7/vGX
JnKij7Q/VqZ1lNUsytMTNxoD48XK+MU3sh735I+rBsFU3mmh+g3u5G0HZxfYS2jF5/i9sgZHrz5q
aMrt8+5mQD+g/fZd9QnqI28YhZadJyItUBnAGXs+j3gKSTEe5ZxQWH3ZIot7X/5ZGw8hHY5MkmIS
/KY+m/pFL82mssjdt00wn/PLGAojZ83D945MW/2gI33qx0Gi5tj/mw7ZLiXD/ln4yAOaEFrGP5B2
3F+UkI2inPAsfgwb6yfed+bWGo1LQF5llC9RbzWunhmsPvTKPhCIgYtg7mhWzk9GuoSDXgm77sHe
MJr/fQ5XXkNVBVJgGdDAsYIg9qfucUMM3uw3cjnWjuZpbOHBZpX0XDeJyjHugqfeORxApRRiWQ4v
0TG764ZNWT+nq2cdolKYnrpDMnXoLUFoD9SevOyOsKXyW0s55LSdNIQ9cPgF5HdDiovX6T90GrCM
jXnz4lVYb1qi1K10gHIfl8CGDhKLIahHJaKhgGGed67XZ6mTky9JO06csFLOet5Lp5e72zi9tN8R
lQ6wD2emijNaW3J5inJekfjtWs03nI4OxQOZ1T6AM8lGZ/O1Wsa3/l5tAxS9HCOyRxZaTyhLfJHe
ftXrozAzbbmgbazkTjfXiZEAiVSYqQCknPBvBO2neNedlOZdDC63YOByro/+/Jdflb+/2p/GAohY
g98qmByfF4+SlIrjZgsfgoN6VjOp8fMDs7dbRFuLMUFJvBO3iwBMTdhdHGFlIjmIi8yvMcpHxmaV
npq52x85ym+GvyEJGgZJwofsYR2ZzWGYtuQAMgxSog0lpNlnEA7ybmsTYJL+7+bpbco/EvaafHl2
606fkcHkRc5kkkyjYz6JB44SUh7rG9SrUrLpt9O3jLOFAB1zcAH/iY17sI5IjIg6Xvq4B9mCv1iL
LjVwdHz+GhwiJ9AWQ5PREnhRqlNUEnMR7VzDNLhnXT3ibK4qQYECfex67U/z5cbzB1Wq2DTpBkB+
cWRAHVKudQ3GcfyN+MwOG//IzlRHAoyn8qVK65tS13MDrCwUFW+E99yZ/VouTYIj0wKNs81SAZrS
0bds2OFS252PHILiy4MT+Tv6F+6KStp0zbQmrM4g+dVT/WWWKZQGNWC98BJWkcXvgAlCH/Ll034M
tKnnvq8VQ/RR2asinYRFrKQiJRiLlNMFgzWbWkAd8DI9ZrENNjaSFQT1AzdeZp60XWjoRL2NfnlN
skhSTIOXRx22aexSuHTT8RsfPkwcxIMpM0YhtLuDAKefF/8iMepYzfRDKVW0mMxpwlAIz291JLDZ
HIW4ESb1v9akcmo1WHpeCtOBWTm2AYC0kMrc8lSh7773uLRIH+gYD/LivkMKxmZTox281ig1w10l
prkc4s30yHjhrau987GFMDYSWr7X0OxKW12wsElhiH9uwmkPuX3ubXQyTacCAj4iTAzxnSPA9uFj
gQbduBzlupc94ANIffByhCKunSHLXJrRM16Q55S0QLpsCUI1hBks8M30v5KaQ/vtxlVkMyyH+7/e
FIE6pCSe5NzhLIAkaPTFRqjiNmfq05i4Bu3f9AAE+Y8K7zysJ023eCyXbS11bePhMjtCYf3mHaRE
xpqrYhbm5ig7xuIQpNGx8ul1UwjiwIEzU1aOUIRXoFog22kgtPIL6MDlbRSYZEFg/CO7vYHHKsWs
xsmlMxHLDT/rnJEQUQ9RTUKaUcLFabChdWJutRKdHLeTDuLYjprXV6s1ytzd8ItJRnzNzMH9Se/b
5wAMR6wvQWHl9GuoMiXCCWzhIi4YG29K04XGZ04rYog6KRGCr0vYI4zBpm70pUViwPIFs2cH0tnc
p6pg59xGVeBKxB0sna3cNG2+1rVB5CPj6+hIDEw+BI2nYNNDj5oxwxMA3OC9B8FGbryy7udIk5Oh
3Jyln+6mjWPBng5yaxUV7Rg3dRMkUO1+r5qpVzq7e0eT9pMgcmZsvhrarmMHgUXeFt1VpG3gKle9
o5F6mGa0yNRP8ZV+bZ6RYteM1yXvDitTOoTFTKNcyNG3OMPzVdM7Tnte7RJRUvZEw7XvxMLsOa06
Dn9WxkUUpj1ulIDRUgQOeaPN4jZv/X6ixxoFX0kqszxb5wWb2Sw8s+651HAmlx1+abGxhkpleome
GHn9ZZPMbIbsn+BkZMJX13M3r8dVdC+UOK6Zb7tn2kBOT6V63bSxHom1WQoWDMT3kmHYdm0HN3v8
iy/39V53vWn0bZXfu95MKvOFXMjbVJa2zzjrs9m6j/Mjg4VyZMFSMW2lGNsNYV0cP1bQVg02T210
ITtHLwP0h1TaVXb548ZQqqS9Ytl6D9luxQX2Gog2KmM01vSQcCEZWg0XWympf8z8OztoosKkkKRL
qvGyB8PrXPCVPyZXxkJqkSpfWaiiVwyvvs8pi8Ep5bai7V0BOd5Z0GbZhIxSEvwmIODzk+On200v
1SgeB1zWjodIIXAB5JtN3AMUa7sp0xr5OGNeMJRh/yacp3BLbVa57W6ILeRhBKYm3dJohodSPTpk
ci4CWuQtc9libKw+C2/ajQzAArBX64LMi+PP8OMlFuKCv07fHGz4erW5RjGVuyLL07rb8hZw6FBO
JWuB2cspOgS0SlkKgmXERO9A5kyfO4ObuB6cVJeWsAhl+t/WJNOWGefXnYLyLi78z5IhPohIVmQp
MUhvtzlwGpP8hYKcludMHpOTIp4Pk1xPxmntAfRZqg2sgHqq5LlySG2WA/cVdjYA/CMz11CQTPU3
MLlPkDQnNdmnU7K5XXfddMop1xRptu3/+3q6HWov1hzGEFPKqaL54D1OCtLReGmrm3p4OYUYm9cD
WU3Nhhn6bfP4zeQLkr4GmRrweD0ATBSBfog2Yqc8IRuVjOUQChWipMpdj577DxC6RHIvTFkbNcxP
qyOLWTJbcWc/4j8pj6nnBAimPkLdjb20riIz2PM7mmGZ7PcGbemxyIV+IiiVqoc2JF90IkHNvkKT
OgiCCB+EprBNAOPJd4jSNOumiTDeTU/V/aBNKNgGCyYpISmYsf1C9/IsOfuSPekO1CoIRcm9mIjU
QYfTbBc2ISbN4CZcIkU68CNJQPi9b3u58csFROiivQ0BZM9Rvt3vSCqWhvdWtJ8l+kXvkTNNrpEB
pJFCUar2aGJxf6CJ07RjU7KaW67Q5pJyVeaBWmcyOw71wMYGoqV8+5Kknr8IERlzP2wxsVEENYWj
oUof+jtiqNPffepa7/FLVr2GhhaH3FipC7hVDV7ElKG94OHw6GoK9anaTatIR79uKUfcUl1+0CTO
YMio7RHpijcge/RCwGH1UGBELCjx649XiIXJ4u+bA7oCRe3zMExdMSbvpYlP/l4rDcfqqo5l5vm2
FQ9MnnlSpSN4nMYBQLVj7TBkOH7wGhK9ZfQAt5ETrjx7tZwdwIBz323jTx+x1Iz70S1QyIR0mDFK
8FtJT+isZyXLM9Q490LbSxakhvuTeCbaMSlxQHTLI+1UV1QK3lIq8M5Dk9FcCdxr1rrurtUx1nC+
f0cwlq0PQdl3EvDbx7WanaKg4WBwFg7tyyF0YPjpudrj39v3UvscArMHririDLWrnR1GyIMyO2SS
Fy7tqN0FrDp6GHR0gEjDSxgYbCjPgDoZWGNVngthMHpFrcPrQMpoP+axSOL/eTtH1b+wcvPmJnzw
hWlQXJfyXN0iWs1+yZaw2jcebAjV7XlcraPR695UO5vYPhvtm7zK0G/oYaiRrDbLynj/Cy/GWnwu
bi6ooVuqKwmXSpEazq9Y2EnFOokM0zSakZ7cvjB3ZA4OBz14oseBeswOoXe9kBLAdHNQ5BfPDHkT
0mHJNrx3BFebDLPLOsuRZ28kgHZTaDnASFuh1XWTJRc6S0b1xhZFWfNrjtSJlPfYWGgEZCCVeR+H
NwiB9vR2lWBrVI33GPpVgaqKydZjqY/O7cUmVUsWtRetVmRVLPponaygqdbT9Bx8HOPmyyZFtr3W
eS0K5LapfPTLAu2Wop/RjEUfAzI/5rlBfpxtpoRC3U2C7MR2U1EFqTnpb0T37bpIDCJa4lp18s/j
lLa9xcrDVwLb3ZGtZtqT2LERBE6ooA0f2rRwFIhwNcfiSze92WqUwjIU9y/FoFXPNbpR61FFgddX
i3eHLfRJrjESMyVHxpinUyd/aOB9L0JokqPJGU4zrbwbuGPm5DWdtQSkgJsWmQ641NE2jhVngNxW
VjKCKAUu88FsrVGJEKmR77++x/2aI04pifTzQPkXA1NOrLMelpTdfNqk13ff3ZJJd7QGQWroFYJH
Y3Tphpqrdr46/OgbhhjiU857ZkMuSXVFZgp1IpfI9nf/uru68SeP8VcfYLPr2IrFhOfoKbLOd1uW
RoudLwPeS7YpOXmhykhXkYlwVAYU4mHBF6mhvHZfCqcTLYUW3PdSxbX9z1C5Ebp31pjF17PRSUPr
RWDkhLeGVdnOvN520kcvKNqkosF4kFmSdugBvIGFRDjMWOzfc/edrCfvOPIU8+TePDGh+xrVl2J1
AXO8vk3nAz+dBqbMp0dF14FnJcbOtofOY/VUEhreUQX6hHitkh7wU3zyA1bzsNjSPhDpC1EfPX0r
1Q8O+qshe4uY4zZ/W7k9s3OsZ0/9KE5twksPTzR4epYjYugQNljxZtba03DtqUcsi3UqmjAYbDSz
CEjPrSTerXSQ5CPZ9aAzkFcrm+Z5PxV6GmDPaY+gXY5HGhaw4EGF/0fR3zejWgEsdfHUjl90MQHC
4XuvdfDI6c3wl1wmMfI8qhrp1bdhI7AgyrSTLB5hgj3/MSvRzbTUcg3REHpjTMh0pEf02vxmxkz8
u/sGZul/Z37HjrrA6bsAclVPyBOWmS3LnWbF1nc3bwK25Bxiw84z/cxSY0IGvEjHCA8XsKk9oNFB
I3t6Q+VlQngf55P0Y7cJwRckRraQHDZB0W9DVcwgFuZapJZ4GywWdYSOu9nNBu66XCemvTjYIkp8
ETBkE7c1ynlcu06Od4f+XjlP7InsN/OFaDTvpdta9uOy9MU+GAbr5V1pP+2NdmaytWXKPsO1pWdX
KV8MPG1ESUWQ3OMgA733qHQX/TaFp20DyKLjYE7v+k3Ivpm/LVpwSIJaFlqiLg7ThlBL/+yTo7kE
8xdtm/m1OUPqcZKKE7kTpyVJEvI1NwBFNs9eQps4OJ0eO1JOxNT8/ifTNQunuJZmBb7bqNBSjcBG
uLvxPPiTOQhYFh3tmzq7xOLw1i+lr1dYiVaTsrxK+hJLLCvA9/VGTBBMWQS7aAriiCwB5+Kaiyvs
/5laIxpW4qdoVXQzv1do/0SnSvMIo0kNFJkh14PUnb/1zZAZLprLE9xl6d9pfzX/NozdXrSQOEKG
8arGGXxWHBLznm6dc0GigZYdZ2nnT9QjYVXYLUkkBeiFaIb6OR7In9P6uKWm3RKQmnOpEOiuNy6s
CmoXuZ4MUDsCq4oAAb8M8l+nYmE13drfM2xcljp0HGFFy5MEgcD8txxIVHB3syK3xAIo8NIvx7eU
Ssons92DnS7K/oRqyVrMRF77SIlXMo2bTwZqgBLeJeZMt34O8CM8Oq4N1iaLyd0j6toNRpLpbJT8
l59bJhF6K4YB55FXRFs6+ilbxgmJT/LuPjgVNdBg/Zteg3NQDC6miqaL3xlLk4SS6nn0VsWdMh7C
3ZnFpqBZxV7X6tTVvXywd9RwC2m7qMxgc19JtWRW8xR2xQqepZWReGsagNrMSixnwUZ+TK6JhZ5W
IIMHl875eXnocFpIFU7HsR8iaOijU6zkwYbEyF+51Ae7QgaOJ5FxIQxkCbSxV6CKvHmirVouaMbQ
BPem+HhzAW/H2X+RsM9tcVRkQSWpwRW/lYIjm+Hs38q4bSzergEe62FK1IJxF5R+O7JPg+xBJ3vV
tk4zwuBV5Dw3d/2zdoWsg09lSXHi25k5YGxXYka6BY5nBzJmzxixag4YroYA30OCA4gyQV0vDW7W
C2RN26+4mMDSaMCTw7UyKQQuk5XbsL1H4ZP8WGr7fdmxci0TxPODJFPtmvSaIfJgziyvcYA29erW
3yCXfQmhVYF6xfjTqGEn/gss7uEoVqCQsMYZlfSzdsg76v6jzpVW1/zDJZrg+vNdGdGVlko2xw3N
aU4uon+JV8dWdT10FmTNTkGgcODCsW2IKCpf87AFi6/Adk4qleFNFLAYE/DJbahiJYewnxzcUKVe
pf1OV0ZZEaPCcblnmYSj4Xeul94Dp8iZKrf8l1xnDA0nSQfY1JS6+/Idht3sB/5kW6vH699HEVzp
Pe9l3pmawvXPKn8FUfJrXwZvwxzMEKBk1evyJ0Kpdedh/2m5oG/JJGFlaoT3QgtBXzNFiwE3lgqV
lG8CWKdVOUI/HcZ4lpN+PPjlEp5I5QvMKzuhjm0yY5jZP7TpFbcLLXM3fV9IVqJtB6E6rVzIrlB5
IOpvNKXqGHSKvr/vBiJEfSzmullZH+U3NALx4Yc6Bpoft3GSZ2DKTuBhBuxj0Er/yLm7fhFebvqW
IZVT4rApzNTRIdMQI5UfJvjMCqFoSajS62A4vBYu8BuUua/L+Wx03l+G0Ce3VZfoWP3L6zm8/4PC
Y1OvDH9+5a8L5Y1u/KaisLD0FvDEQyHRcrAhWHUSMVXPSYDgoblb0BzGTpAePFFVUnyVlrawnT1h
LAUmMUzYVhpbE3gSofmjUuZX3PV+Bb0CIy0SlwDPKnSx3bgKn1ZZdqYG+msC6BfRWD1DVCveNhVA
9Q+LA994WCDSJUScurOnsEot6F2w4pmj4SMwx+KuGx6HTguckJgmB9r/Xm0lv7N0cCQI6l7eF9Uc
5KE1H6ZCQg0zrRsdE+sOuwr5vhsWVQwL6Icgi/ITAPSj88KCIM4M6uq7xEmuH6py4xt68Q2itv5j
39O2iQXziWS929ML9LEgZ4PyShNzXQW8TAdS5kExvYY0CAQ5vqat9sZq20e97XL2USKG9AE9Pp8S
4F0IILS+46WIHKvYb3WgqMNteDAPcDBFFbjWoUqwHP9ZPkDm4vTSXkorpPUY4/9Ssg4xF6IRKUL8
1SPcZA09/ZARqJIn6nQAK/ss5apNL8jNx5/Y5EWhKUJ6icSpHG1U3HfFWuMuvDVpgnTN5TrNJDeZ
pBxs4buQvoQR7j3Ei8G24QDkMnX/B5YDexIrWrzdBtd2HTlRVTAJgJDc6cZSfRfE4ovp8yZH2dop
tX/HmDDnjd6BPpC+cwpu5OembXHTgboBDGvBBIDjHFn36qMlahYH/btaaii5kpKwjYOykQYs2Eh+
UJCkQhk8ot2tm9197C1o1+mVMe/KE900gu08yyOk6y4YYHYOwYYKOJHmEenAejsfGvCsfpogLvV+
j7YDo4/gjb+J0CD63HypT7voLbwL3z6c+RIVUmrhDn+ltGze7DOK4yXxAtPXgzTguhJUmkzcpkXx
qfChfCTgK36+ENoPLyqr55xhkjDHunDDbb/TgHoREZ5OXaAx91Y4v7mLT4lR2FZqwYyAJGw1pYiT
j0TZTbKJpGMNzhaTgkh0q8kSljHriORLJM9Y53t71giLwBfdru/pcafIe0uRPHHLB7U7I+bTTkPV
J842EDwO9wmMhp3tpvMOZms/98m/RCjyvOXZ8Rloe0/Ts46XpS/Wmo96v878cNK08KI5Ljsm4t6b
nkwDEjTgXaYqtwup3NW2DgHVQYItaNeOtFQYEF/I/RoxK5x0sQi/QiMOE2sffNM8nOizvPhe+NWK
S/7tZmGoKx2KAqWBYICo9AK+prXFauN1/OLMBUGI8QschWkSNPvaIetbPBJIYeaB5rjrNaOmOx2U
yGGUzst4TLf4okbgjF89jLqHwqGlPfdt+luBbHAdMawVMoIAw6qwgg9+1rQWyXejolXO14FhqaVA
O7xIu+v4Ucn3jK9N71e02HZ084H1PrfwnKD+HLmLqiHXAY05wRGwZucCuq9itjWAtHbo5PABj/nn
/TVvikE5QamxrdJdu0rquCJCMv1tO+GgTcA26/7NoL+cLYIv66SpBQlQ9JIS4kPnKDbXjxUlOC4G
bYdQw7tvi6ZWDzOFcJ/Mozfwm5mJmyTbwL+jTYte/7v3n7kUqvhcP1QKYPkVtbbeyq/icdhusyE8
VchMtVZfcGVQKxPxZoXtqNm3oHLZ6ejb3fSY2uIXzwNs2Ucm6tt3VYIWjQd2vLnArBUKKMF4+0k8
sxLDQfsThbKn9ZDvpa1GiqMqg3qq+toqB8CKtOFe6crJYeNsA3qN1IQ1xTv/oWc2FuW2Gqx9Exfj
NPQooInAcycn8zCKKuJnIpYisf4N38nifzknoDnv+6kN50uqyjg6fTOl3u1cmybcZKp91cpVDEiA
Tls6wDFiyWHgcOptbtPVvOvqEwiLXwgus877oXyQvk6d4de3Z65hSavu+jLUbBZAK/zVVQYgMfcC
vMmK9X/FixhQe02uFy11Nvzd56Ugl00qLUW+dz1ZfOIjO7HUAmcSVVTfsIbMi9rrABhgLD77ewop
7n0L9WIWt61I80sACP4KTJ9e0YwfjLhTkLqBgMkBdKZXT7BA0Sfpi8pdqAGfPQuAi+RJocbWpfLO
/rBilxqaMQAtmAAjwowDmOeIh1b203ZsNiEUySeP5U3Ugmh/I3A5u/dGgezpAbR0v99fz0FA4dkq
sExdZB0yt9iKM0FzgkEwFBDGK55g0HULZFj19mG6RzkgZcu3EiA5B66z7d3QyS5JBUhEbMO75q+z
/+78h8oKGFBL80U+c3CNEeEd0b0vnud8IO0kLbe00floK+Z1CqxZfgUCXfSesxUMufCSifgFMSid
qOAiwVzSTfsDyn4/PsMawv8KxnsPAbhIry6yh0UPjT+sUPVfDKCuB/iVAx3zXrDdCFeGIGruGmW7
sTwGsaUlTEn32/JUEeTT6G4rVvQtCSR055SzPfRKWXjlVSR1CLQPuEZR708r3ysUUIGP+Vn4qnIQ
nEvadM0TATKb8/Ikz6/yN+GzWkhCA9jnQGRok0P5oAxMojDGSXLvg5VaMaEjzmhGWWNCD+ygfC1r
0TbVWGyQw+zU0ulWvcV0KhlzicRgg5VJ6sk+IFSu5xa9ait9o7RlwurOlCYZHgUgZSX9hdZtz7hh
JTUEfiII9SoteBknndwJc5GBTlP17uXmBqvNA9hhHax5nxbufYYYqfD+qIDITId5RJlSFeQbQcfk
XxANday6kH3ZGyef1pD9ZzjZ2GmsRy1ZTpZAhoSurWUs76sJGM7Gafd1k6Apdtymvs4Rgah3nD+d
WSp8z9TkuZ3shxYXHX+VafN+/rO6h+rhBBjV+XB1wWsA92ibLqNPrPh6B4r87sQrdxUB3WWiuTOa
EwiWLar8ShZjLGkISGqRog7zFStpIxFfNYz71fvrWwtR0V8ktMs+e8DGV7+Kj5Gyr5WplLmeOMZm
xoUAheB+NC2hI/BjpUfwUB4cMw8H6Z/VyffJP/P3SusZac9Wb6dBS0ZbeU54IrPxhSdxZ634l0mF
930OnRKPer0ShOcZGbzeAUdHo9N/RTyALZ116zs2bIp15tBsEUY27wfvtODalue4L1hzMtEjDyHW
XD/hPgaUKkrq0wplISl678X/gNe4RW37ZS6YgPT+NMbUXta5epvqwkxPNiM3jVp2ycmB98dRuYhL
j71v+MasAby7Vx5ltRMT4sL63Q+8wxCz5okmDusDJpBH1ePNnExhxcdsWxXgUI+VUCemP5cYVlyr
GKhsAPU04dEO2Yr5mhCI+/znEmlpywHVEs+Vq32l6fukS2LnQK4GOM8Rg4BC+IPbs/4OYSur4Qnq
eVLN4dxGjjH6b+NxBnjM9hwmKSEdC+EW6UJMQ03oq6xS5cCQbPgcNzrE20PFQhmcMSfcnvUf7Mkw
vCWZNTz/9E8wqBFSOmSkxmZC7cDhMG6seCiucSpmeQna+7FAazZJDahCu/NSHItIxS+lQWPDpB39
DsxyQhv2OMoohSG/ZmpD5bYLxa4tvS44R/Xb2T4GBgazEOxBMa6UAE9uel4eYpZZ+/fRFXC2gfsZ
ykpISJteojjuAt7KQgLOnL99K5jSzYsuG+7+bIitcl1SgWZhvugzqPndUQLtBjOhnEbX9Icql2r7
Lki3QatbZ5QAC+3Nh1x1HrY+Ehrl8uOCKu531s/64nAlzYALfatqzbZF7t2mMDvdzTDTT2aC8PUX
Kxj+jtgHQXw5a/m83wbM4wNQWNONaISD9jo0O0Bpm2YporzJXwSaZ3BKkNCDMhyBxKLzsUUvkejY
AtCc+drkpaOjr4Q7YxxuwktV7Ze3vEmK5Zp/mzwXUWk50EK3WDUZGOxIkHEoF8mt7qE62Lfr/l8x
m8d+ZaBK7N5ffi9ijgv6/xS6ZMQ78XBnOQUahXf+HGbDYUL7p3dwnq/4QIkHNc60i15oEzclfdVM
AHsekuifr/2a6wRJTZbjHL2Iet9haX4Yglio1EMiOevGx6du/XY9nhyYSLbrJ0WWl1QIJtM0sqct
pe0Qsatv/cy5hJE9LLEcpoAdlq4Av6XxsdPD+ju9AHDgJc4wWxPunAODFh88sO+5hWXPPL7OwznZ
pocmmenpzlL6QsWR6Nx1rbfk26P9cdEo1yvhJ6P28yQYqrgJffyJf12dz8Cbp7LmaCir6ygrpZkF
HBUxKj/X8bys440qPmOokg//aB0Z/sJNahX35Zfkf9xCzlSiovYh/ofEs4VxyIn9crCXWUdX32Ls
QTVYiVu8MXvpERrsewAyqAt8d2S7rj62pRHfQw/s6oOJCwpsDEWUwbrHe8klJwNDIIfgpXaWjfeN
yI6dhMRIIHyQn9g/DeN8tTeSXDlxFV9dlAQiQgi0ebBPMk/tOLlAt3/MYGFpmifW6CTDc0fBL+fM
iH55kVuVDnSsY61PKWG24gGHPLnoHOrKDQF/zAMV08Pd6JpzO0LQlxd1ot5ZiGhZBZJjIgZWYiS1
1i+4KHeX5JZO/7DsbZdaQt9qLcrMkZByLzRu+2gyFLEFMEV4wQXIB0iSRsCChmpbhzqUCOIlH+DA
UheQhcOc/HniDu2DFzgyDK0QDUTi1J0PdVgJCGbwexJYI4BkSyFLpuPHzNjlGJBGxbeNpJSk+0Ab
DNpRtauCsSGKHDQ6+KozTZoW/sPLLUZcaDuve+ODP8dbu5oUjebrkiuBwd4o5j8E8RtbOxB51Qn0
putLUrAZjpfq+ag/QyRUmGC4y4jVs9cAhaKPOiuoXI7Db43xtZDZbYPfCeoqHDOsNmw5zjJW98Qp
kjqdVbIW0ZMNCPcm2+truzcYgPMhKO6CH5y0djOTQNtt1oTBqVOXy0l8dAsfZS4BYEQbXnPtQC5C
NHP+TmA3S9MbXBJ8GdHOiYOiJWSSAny92ioL2c7S2ynPep7BPK5uvFxB6+NQ6MAEoJK06MthfTw0
XnplOxUVMoyEyM0Y9BqItV7uIpOg91cvXIr7O7YezWbAHpwjKFlmWzKY97CWMeXCu8qgkcvj+POg
YJqpzDCVPbG/nNiedj4pFv9q7fYkS4IVhBnMjWPbfeFK4jT+b8Q9lCHtE/osXrkWZYK32Op7rN+N
5X8W/jzvOnrNMfyrTEN+FE77zT1TYPr+/JXlc3aaVKUaeC6wVoHif1EXEF21D0gUHYMMCPm+z/zq
akMY9EITdpiUNCvgOxbpJAd0NNfVIGs4EDSiSErpEiO8IH+9e/wtR+jbmuNXnfoUMQIpSopXB/7f
1U1BRpo1yrKOZ0xGmQR3w/JYNm5impmhYnGIA5ouccMN5GiIIFgCKcU+J268t/fQ3gVtKgN4zKN2
G1jvZWgitwGCH8B12JCsqzN87gdbVLM2F9POHB775tryPgchIvYjahn0E1my9+2WrgmKL94oq/fi
amTiMu1heeyx/wwLpiC3hFA57FUwQpPRfMYKfVMRVBBuY0701n6ulqdtbhfwCpmMbJKTT4TWqJ0h
cnonXwMiLG60qTrO06jdhDRAS9a12AStP3qFylt88QMr39oT9kNacZ4nZsXHoBjFQcrb9piFoDd5
3lz/WZ6xLPIyJnEKwtcZBSCugGxvwqpnLSfDDObRfwyIMBjv9ZAYLZnNhlNLCjIptOW05S/K2muy
dyHLhW+rg/GpJ6XRE3ipw38vq4wD6jtIvR6d7XPHBWrjRXvu4KLbWiwAOxSh4rJDoJHSQjLbqwdX
3HuAg/k81HQtJoVYHg2h4KYkIlgK4rc7s7hfoyzcOsDk0ejaYVea7mn7f/rXAxDcRTeLi1UCbOix
P4L7iYDnIx4kcS3it/wGEMVDLxWLmnlrPYy1HgDzqoEpxI4vbs+6W1vQmJ8X25gqiTRGubhn6pPD
bNLlLfvd46NfzifKZJrFXxu+bxXHs+v2McVEu4UhQ/fpJA7GcW7e1+ExCjbxgJnZ63kYtR6a8meg
haY0ro6PUw1fT5cQBbovPvMvvj74pzHeby09JEvPvbyLn53zZqs0zDzAkILEgMzSfdRcWukecBgw
0o5CF5oGKQ207AQm77wKHgB3iq9JK25/OzbExBkFJdahwY37WSH984nQl8T69jYAfxR7L7ZkOLP6
FPPl7/EjmnzEAJYNNgkNSjZt8XB45lTn55qmbwZR4gE50E/2tWTsuRQ2sJkNn4pf3uYyr9xbGe/X
QS6r8TtdFGueNCZnAn16o/qMRGClUO8F2U+a3DT+N1BTM+VCjOCYNLdHiMa8NnPXganjMJHwcXLR
exERVwEs2Qzko1LitC85H207fkRKbyi92Bd8REnSIuW8nxbHtDvxOyrLSPf9Fy6SK9f4UKkWMybr
CtzZR/A0kDNKijRzEHahZykeCUcr6UxSqw12/PDxaNKX2gGqK4kDVqcT/RPYpCuvKeP25WkIqQAH
d4+GHdTCLbDVkd/H+tSg6yVhXezuPcMGlar4CMgl40fmwhfDUFl8vRR8w+qU2RS9LpUVY3L51az6
z+ZfjqAhwCgCqEpJ1YyUPxXlnFmeK1pS+k9n55Jx3vz+63asCmXpQ797l/MDcYUyEYOC0drmhaF5
/QRW6Z5kHfQAAzS+ytTPJVs9wxTjLYUsEG4FkxVG4ZijFXS+bOguKR6mdTn7hvECbrUOw5Y72AGk
WqovodE4H614W76RYEbRdnHzf7uRVueOGW0rVfPhaf40UKyUSEXCAp440p3TIowvqVtIEf9hAZUu
4+T5YgwI4tFeCFmfTbbX7VCeank0zG7WsLhseTN+PqIRwik20UBJ0rDl8102NkMXujjwkzED09xI
3Ban8/IEHdzvYhkBn5fC2+aMQPgTf8ZQ2BFXoy0ivAghhRz5QDYQGr8Ts8H9fI2yHQqfnVjFA/HS
yf25T4Ts5VysYIIiAceWjP9kwC3Mnz1JN45jPky8Yu46qa75RlpLadQdzu2TPq8Io2vh33a/WoPg
OIs4vO7GgMcAwLqdhZ2EalzNU+8KSX1Ip0Iv6GhanxKKp9BrcoA6xiTAZrOnzB/2d5rN847TxFf4
Tm0Y9sGUVNZMGfYEICSvF6sZyuQMTtaeTcerTfBS363GfTSjHl5K+OayE1SeBNBbNXhxYPNFAk3O
dKOFqnenOcmpw/m+etZFl/a8RROV06LLBzkCP1svH3owWrMZz2oVD+kdMSA6CL9Cg9DaYBUDpPCE
rxpIuIodGygMLTon3Wc/skAEU8OCOPGChze1/1Vo1hZAPqBM/a/rtfiyEc2oUSit/aIe+gMIht0x
GT4R/EloA/fNDJ5+7htecdr9y8CrhThYSlRWjaMLqDciMfSMRpzk9wzxXOavFhEnH3yJQL26nh1M
Nc7eEMFyCB1pjRfgyPLLsyalFunkH3LtK0qSJB/PpNg577Z8XnRVK6K2HFI53xCUjzMb2UAvcOey
l7x389TOYC4J00TAiHQ63A4RBnMg1HJSwIY6IEDU45qLRySQZ42xWg/IEhErZxf4Rf8JXj3cddT5
whhtGohgrZnYfmqGky+DECMu5h3Q9qWZxsxrfDiDQhISVyUKmx3CYquiSljFOI3HR08FI3oEjMYA
jnFyKVp9WPotwcOV9q8WJzlf6q81lxdq/3ZZxxbdw2VPzJBIaxde7Dxuyz09pivoEy27NUHlDe4O
/CfzI6rbINFyE4eXqT+SQYm5bo/HqX+QcTCEK7nagFnQJ6d6AM6dcFfkqO42ogyrllfXHR7DI8J/
zkHMQDBYYRuIK3LFqy4chy/TrUS4H6QxmXXMHi9Z9LrL0C0MbkjngzPL5YT2LCyA14hXH4LiU8rL
eKV/DP6XFXvi4pd/el8UC7x0kZovLer1Tf3FQ6tqIZyWS4Ve28GFvVBqlal2qAGzFnSXm8LszFya
lFYo19kunINYJboy2Grr/OWyR9TuDk+7f8wZY4sx0/nEzA5k1EIWJrqa1v2WOl4a3OMT25mvwNzF
7KzdlvIXvqnFB5DDTe80muxsHkPto6JBiWbsjtSw5KoKY2XkLE1Uz5OF3yix64ukgnGxmmgAYP8J
JLbQ/gDvgVfYjKOvLwTp08OcR2eVHX3lu7eXp2H1XUzT1k9Fo+RVFcNCJdTTPIzmDcWdzDochprJ
32bA1VIEwSv942kbEvRvnf/EiH+PjNbUNLwXz42gQUCwcdr+g71YN65L8fKdRAoFG0NdMbo811Ef
ByScKEWMnQzagNcQn2nXj5nM/R2nDDcH90ltc0LtTdt/KC1F/VKQIYIPSsjsPW3sqPkVyDnXH2lV
oj+Lim8zGQE11XeWrZ7L18daDBizDs/thcMaNVuBV99VgQw65z+gUpcPpd+ssuhsGGRc0mESvzlt
iEVcfJ1WOOsfV2aLkIq7kWni0Y8uNL9vVo+7F17ZsJptDkX0uo6I8Uii+mAY9ojIaC5xnyDUXlEq
HNENlV0us6jO939veCDMSdUQ5N+sRhAAagSXUQol2xK5yPyhAeQNXT+w0avvyx5FSJzIYkdpViiI
czg9kDNtg2P4uAZgf4evXcRdtJxCYa43/BcK+riXTHo5pQXMB8gQIbfNrlbTrO3aTvkYq+e4dlCv
htRuvwyCfuJ3teEStdeR0TVP2NO7KGpzXR4Ww3uQpumATYd73hG+9RgxayQfplznNeNmDgvLbrd3
+tYC/FdGVrvq+l0ZjmXyi9vTJX9JXKYA6O9XP3PqjNRUG1LSd0MOVs4/Uca1EM7FaFsseXzQLOXM
fFqiizRisHlqMTOOSYWVAk/weeb1MwH+gdiOfb1rA02sv/gRDV7JmTOa/ROVZ2dppCt6STGIu7vf
TybkAHHYrfp/0IGIFq2faDlQ7rPAhG4JouRUsxVLFCIwzU9McmteN/9zJ9gFMJnl8gaJ/lQLCXcR
MXxDfGclwEcgkMwe8g/hFMa1bDHZ5Leuojo5Ez+ILAGjLfLzWVyfRYXd1olgJ4nMwSw+IAfoaTht
+gSaXqSxQTk12eTWs6GoBmkesOUyVyVnTRPpeJJJ8nm2uzigeHa6NvEkj/LmLUyDM36QZwGb1qdk
XKpZBGXTy3UXaS9wH7K8Q7nuV2hwzKU7MhbCk6NbNGzyZ8pd953jwpn95ZxJDV9bpDX1JJTPLETm
RS+jvBOBJzjyaDyXxmMevQFH09M238CwB6nznkJzmRToCcPUGJl3UXrsA1XEQbHGLIkUtr5WtQ1S
7Xg48TT5zcgdcwCsawTSoZj3Ahom/pXhwHqjx4PK9VjJoxW2f4DrQYx4oFNtVcUGdfS73tRGNm2V
ReubGSJZ35NQiMIsAELMp8U5iO6ZJyrsGmUiT5Zp9QfBhl/GAfGaZnGYvyuA/B5bAtx8iE18uSW8
Thvrp5HRhE1pQOw90tDBhaix+uitsQpwEmsxG4OlOXND1U15R8SoPFS4lk+vpkoxZPdVb7pyjHYF
G6HKNsdBk3pfqPOk/mxeld0fr5mR7d0AXlgkE2T6ppYiLu2coZhGw37i7SkmC9QIHkgLwBMnogFI
6d3E+g3Jiuciq1TmqLtR5YmMZkB0UeC0w2h4JN3XqhuZP/+jKsFlTupNRQdzPRU/c9E4+QY1hktx
op4Jdjrz/QkAk3b7LW/uX0t9+peHTLUGDPjcdmNBMn729ZD++zQ2cbfAsfeV5Pka2aAvVgMy3xmn
aWibvhiSEwx/clkTKqt1V9qnKApgv0htSl25CqqJa7LzeGPla8FGW+30Iy+B330wjEeJgL0aCaV8
ipgO3E3anK7yJW7l45TJNSvcDW8lKm/6GbzaNanrfiXTKGztx5pf6tZXGap7U+xebgMcY8VU3bmt
GcH9YkhiGlxFuhAqhGLibN4kolFbEUMTLS5lr+yZf4hdi3d+hBHVUot3sny18YekQcKQwBRttOBI
HKcq2suVQBlKBrH4YNan+0jF9qf8Qe1W73dP3ubAJYHVcPfd5P91bM48vKWTY4RtuwdApdzBjB69
8mhjBpYcaaVe8FTEB10aenM387OdOU6liercGJ9V5MvoAgP0jHvLIjAXM1jHhfdRk6Iy9T6YF/66
j7mOnOK+k6p28ggpMNOeRQAZiygDSTojZY9ZMz3ZXDSm5OoiK6dql8cbEVHa1uWHHESz2l1CVjsb
zM1UxbPZ5OFYPXJBem3xB/pWQf/enOeflPlU79DZGz3GAT9up9sA5SJU71niSNbTh8keAXmgMafM
pVPUyuSlUH2vSbDo2hA/ILLItQsNtKJlM/5O3Tw0aE4rdJNmYgZnIHQnjDqUyo9l+izd44W+eESU
A+hCcIYium/Rycitzh1Ul6zOaI0rn0Rbc5/6uCumhJspBBLQlW0B9CylV8NjNMhUx33Fhm936C+A
FPcZMEEvCy/2DXCWtnMaUGuLngNMJR3y/VFjFexabzS5D5DeKkN8Cj002UpvswqMetTG41KEgJbp
cdMwJiW4TJ2YpAsN4veQqkxLTdPafAIPEk0pvRfpwuVgEprd/mQvKxl/KxzaI3oGVcv+1ft6J4YB
6EN2QC3Z9++ktp72mQVfKMS7UBFR5LMQcl/YjyVyMXxHC9qlWkVqtxxfTkprmaX6Sma85fnpNh4p
H8r29Ei892Q9cwfqAHI58KAzbTdShJRpqEF+FNfey0pc9HK/XRBlNB/9KDK8Aj84YKd+cWjz54/3
SwgjF+AdUhAjqg5tRBVOMuNAxTSc99cnTkDCiFVoomAaiMRchYbN/DTieq/+MiD++KMIsF5MUkzc
fGi6LAWcuB4MqQBR8SnAKCIP6RM4vS6x59+KW4PGJFwQJ7H5HtQiH9hahsfTxkp+bqCAYGBSU5wF
LhzhpbRzVhBO/J4E2BPTKoCJFEpKTovQtwKmMwvW5124kXKmGGy7kQpi7k7FtkQ7eTg//gnYoTdc
W4fjroy5cYmGBiQ2mSNXqBb5ZO6lbiMK/DBv24ycofVJkaKWKogGwofILrSSMFBjvxhsBStdm4Rr
NUTQGeBdYz3kinPA0IfYZ9xrHK0tl6KzXOwOorj9dMiK8unisifkZgy0pMJAvw3VYNdfhfesZWaD
Hp8tECbEvBiytWoE+zIO44v/yvlVt005nXSqeO1QtRZsKQckr5Nt7EDtg8crVKbUfJw03p9aw78C
rkMObEJXONplm74Qrii8xbNIjka3EbtcGv45ETSvSzjOgohOQBvNIDrrr/DpHx50cynXB5Y6gMpG
H76zNwXJcjXoqM5B07twXFZjPHA2MRhx9GOw/PivAaVndkNRW/Eo4XL4xPL1S50hp1DCZOv6x6U0
avNkSS0GSlrej1v8bgKkBiRlFDD8uWnKiAAINZ6Bvv+OlgJigjuuRcbGBkWnyVc1kd1Mwqf5brcM
fJxyseQbdn/T1Wc92IOL6smjHE2/yakaVAfU/TBrsF/Z5rNhvJX47puHWuTTc2ZBxLj3gNwLKXw/
RmaHU6V0ROK5nbqpCwsG+GSH8H1YufNppkags9RWt2eB2Aalaqi7RdrXsEh7n+L79cj4/nkdYTeB
SFaTMJ9ozJ+BgkZ9M/mvR3ZUuEPOgaGtqWeOlQCdv0KQOAjXs1pa3qILIw4SoJDph7Xfocz7p0Oh
j8+0fX410DQ9QPj4e6pp6/p94nd+L1N3VRzXW8fzcMtONm0Ywop6t3tELvVRgovhl8wLUaku106I
4Hk2wPRoxkt/5YmCW8CAG9z0BweOI42sKZ4r5anVbqCmKDcAkPz/ZqLiTaGJhhMKkFzQKj3X4ezC
UjsrX7YEDlSrWbX8EjshTF8rGngTrfW+I7SCo/fKeDBao/TFZal0IUBqDSRyCeXP4StNNAajLOn7
/p98tEqqZ6+MoNoyEL4G65OKnOX5HPgn9CBU+hyZEwAlo7N/DhufIE2Rzw5z62KEbSXYkBbz1Puv
l6px5nrxIUXeF7/gF/tGchVI7u19m4WPmOwvyc+fQs2QsW5XS0iQHai+JvvnB9InLsFvrIXMGBIj
7RlDmn0dH3AL8ot8CUAo2Ua6I+tTzyjmsG10M3WCriKXj2NHy3PSbDunXtT5kS0n983kj+4NQxEZ
7I51UwdajYF4PBXayEYSvtZLGyrM1A9fMF3Vk6yLVCh6FB+skSDQy8NxuB9h5OmEfWCV8AG/4fc4
LWu/QlQqVHlyIniPsoA9YyYJRwSpyZODSeiWQag13XXGdghRLgXdoVaonEKZfH8P6mdd69nQA1br
kI/pd5deLyjsrRSsHFRDNM/+z9rCIi6GK7oVdFWpnWvddHzO5PZXhvTs9oaDMgcDRCI4cJR8m9VC
I834yOE6hamkabgrCRoEsPaqtYHeFpbD2/GbeLktbMQOAYh0dUaEWStMODR0Ckh/Ii+GwG0qwhER
UUlKOE4bNd2S0BjEQDRZFN+KdOmoXtj4dByPqCm8ZBkxWAf0uDZBY+uZZhO1NMcazLhzUNcHWNu7
rfPVYniMWMG4a0kxucRrABp0D2vUnsUuuJwy7USlDCevm1wEBL4Z/N3TDoN1Upee3x1eFgPf3x33
yd6EyjzazAjWKf/r9fDcZpVmVlLIKd6D/PB57cGV/wg8m/5/0sE833o/NDM/yAwAf4BhYnf0DPVM
B6CWYZttKud7gD31yuSGrNEn6hlTifcodELep8/6sOTlIrfdS4nsVWwT8SRyDX1vnXr/oDCwb3/x
hTpWDGz85Nol8QVExI4YlbfUq3WhL2/IuQ2ToumiblJC5XgadqyxBEoDWMEvH+cobH8b7OGlz1rF
eM4zhpoDTwUXcCT2mAbaq5Y3NStMkywTLEt53NjLpRKm6dsANSL2KVDR6DGTxVXxZycSHxMIG/tg
Ez1EgQzKWlkVywyTVyr6c9fiSjV5RBVQ3Ew3eR70unQNTu9njaDif9ksSbhVVXiXKoA+XW/VAKAU
hVBrfNv2hQj1AbqELIvnfYnOvuBCMxSFSC8AMKTvIe0IUivwZtLRAZGt4voPozB6Vh8TYc8L4ENB
6LrKXO2neH9lV8RKANv5/xn0hrED4cSk0FDYdLEHSN+Bbj4Pj5ZICc0uFQOKug5cVljPDU49HERv
fc68TU1oi/B98TGQ++OsE6Y+G9sW6jQ9p6FdN3z4AONxLcEhFmdnEabHNBTDmkGLrmYItX9LVldS
V3gim1pWoY2ke7M9hmcSP2sPUG2NTHIFyP8SLwfbwwc8rjMFJaIB1+HLpswE7MofvzGPMBbmg3gH
19H6rLy3pZt3lestq25s9iGzVq5H/o8Y09ItKjCP4jt/l4e7qcXkVjcMZa1jkea0Z+jnIkkiFN4W
0sliTVrKUQ//K9Vxdk/BNBRZsGAWh4qE14Qke8/hDFdF2vm5wWb620K/4Q/WwZvn8nzDeEwCP8vY
50Y9qGLyZDiuOP/QuVzU2UKmUDpjoUZnMnOtzc8BhgyIoAjvShoEaEjE4rc0vdQZ7DW0CqWj86df
TwSNuNPfQlsrk7y6QrrpCn4lDm4BBuUI9imen+c8hf7k7O13cSirt9FL/c0q1sB98Q9og1liTmM7
F25c3RGbgHGjTdHqlhqPKr9ZgCRCl+Dd5UFAQPuMhw+6jnymXEX8Gl7a3rgLUzDb2mAgkJYM/7MI
H8BaNL+o6HMyvaH4W+7HfAsAafCg6u1l8zZ2aL9V5v9SQeps0M6qjm/4UN2HrEq345a4bX5HnNZx
xMmqQurLvlTJBIMcaBECbnqUhnwjjM7eDVDN5s26E8Q18TkgkrP8UfjaoiVzmc2rmpxuHGG9mx/d
ESLnC0Y/3x249+AUiUlLUDWlaIcnf2G9xFSvekl2SCxkYu/NDrPLVSr0UxIUfrDCs85JM7haQCzp
6ubk/4N4u82iiz7JMAbsPMiRHrdnme8T9ac6euHhhKJU062ZDEDW9FWZPC+O9YVdEbIm/cB0Foiu
jPZR61DCNhmV+axrOvYrRly2VFKmpMwjuHh8qLEw0XGTcw0JZ2RXHlBSjIbYnjB9hb5tYX7ebhmL
J7iLaZKpWl3zU3bvKI75Ie1FLD4DO/Ozbu00IQGD7VK8NxbPefBGvtlbGFKpfHGBQc7rXBUbXpXq
ducJLNkre3o/X34qDgU0d+sc/PQACaKjzlvYlWThkRmzMU1mWEI4orj9L+W132E+mACFWIprBTKl
XC98pTXxQ2G7g77Z7Y4Z0EJidTglTHX5qtMXZhrk0M4WEK9VMa3oTeb7CBn4U2BppmsJeTa/8Ujw
M0gxaojddB6D1hlI6uViRHidaQEOg10Qo5zqAtKg+hAwPVwzjKSATtEGrJNm9BNAC2PD9BSzM9Bz
9dwU5BdWuWnadtohNzo/bDw9WQqkO6wlFXONaGt4fehr4ZHnUitc7gCQCgUVn3ETf378eqCEr2d8
iHtTqJfChrehT2P0kPBhXQAW62Nt0yxxS90hesQ64BySbeE6sFrPKrrPuZRq3qb7Yzq3KAip/vKH
+7iTyKq4upkpofxfUffeA3NDpT3KnqpTEWjjpt2zrZYb+koi84cq30iA49abpFnLLBUK8xrQBIFB
ZgrIOohlFoKNM/+3FLSkf9fXPB0nvyDk7avX/nx9q/q2af0i9CBxIfQjBh+MMe/RkPICwpQwACZj
lqgdb23MLfCnlEOwOOQyITAy5ilPrWiUXLN6aUBF6k6cylDWmTCoA1gQecDxztg/k5XIbYncIDtB
vU8n7Q7fY/IWsIZOgw6kZ1D6G5UYCzkXmdbSA30Y6RM5aFeB3h6liH2YJuNGRXUHYipf8vZYUfTG
hcjlacDgNUYMpUBvc7aKUemSQlOPd1MwaPr6wegwFFROV9G/tlBbDPiNwCpOeu0X30C++rEcOddE
o76lPz5mRcYi7ukygeik2wqB5yvt3I1wibYEDsT9sepUlK3KoA6hGJm/zIJqD+C6EueuiGX+VCig
dEATDVut920DNG4JLGwDyUbxdCyWcwsFSv3OoGnDsKNMjr3//7LqwUcRBQx60XW8lcP9b8+Bj9OC
dnxqzbLsjG/fQgZTwetz8YQJoCVbwTnvVREocy/z4SVxIVLoUCpzJgS9sBNwoTO1EKdDw714zF9d
f2F3gemZJH7xB3BkniSxUHH2T0kVPBQ/AQ9aWzahMx//2JAbupmWtTNSK40ki1F1JHapOkpphWFE
ZNIdAI3lTQwbstOUO4B++48jyAh9Cqvon9EMgS6rK33nxJn0zZ1oqxD8TvZWDZ9mXNAFkHXK67d5
1l2+SDMtwc8v4YkPidMXETjM5YiTCkH4ZgzMsFAmRIhRcwH9dmW9oMqNJz8g958+X/vfC0UQpdGr
mSaXOD9sFT0+4BtFjlyPmVhQE6I3kLOUpL6t6QHt92Vqfn/ZbkJJvyQNdRFAdp9lq5I6ko/TYtLK
HIM3PO6iC61xcP3IPv576qGSeRclaaB0tT2a3gzOBQYvNk2riATSHh2/OvKlPKF42EuxmNaXk0ie
oIBkvxiTEB1XdKaO7sS3cBQcmQ8BmYZ8KoyJNJA/s8IlXm0Ni1EMcj1R27Q1TsH++hiUny4giPkF
q1AFfApY1lanyrQBjHNxAtD2bvWK1ETc43sD0vown+LXobRNIRtHnc8tbymVJlhO0t6sYeXxo7fv
OMSMEV4Sqp58t8OgzszLpgfo+hTXoCAjiJV07GXEtie0/anRwQJuGrg0eJkdl29J9tKEFozheDMH
qCXfZlHXnpmM0SWgDbIbdoCCzhk/VtO7447LKiEfpbJCwWD8zFuEYzsGfFIwowxgcwIiSBAVznBj
VJ6CUSq4qPO8+Nn9W3gCzpaorZrYK6cbc7rifDzE1sKo9Hns1YF2K/nbAxabUVzc1i7tJn5wWPHQ
NYnBsMppUaSJWh08eWy+LJfVBAKY45xuCh9vgaTlQ/ucTftBWu6mOIRM9dqs/b/6aWe7QSVKQigj
HEiBm+plaTfUhua75rgYdxQ3EPuaqEF/k/MWHaTPxl4mIZpLHLfCNjQ88zBmxWsn5qg99UlTZcy6
TfX89nxVtYBRMoZQBopZYweza2yCaWGTCSelZqlGC41f4TwOzH031BcTWsyLGJAyo2L2DXIvIkPZ
7beY/Cm/ljMC6BVI7kiCwVmw4eDK64dk+nLnkHZOSPdWXsZ/FhNfd3317LIrHAgQnQuQ6T+4Hxy8
MtCBoT2uxoRKqunma1GufIzLnx0F/0v3gjyyLECYp0R4NsV1By2dFN3JlQ8bJOjZVjXzsHEr9BPl
w/XT1J+dlQFYIaGVkXiKNSzvhxxD87qUzRtuiYy4/XkJ6shY6Bmi7uUGacwRytsXxNoX3Qa3rlci
EXHkI4h7EBY/TODAyC5q1SzOyKT3qdtKARFDr4fLZk1I5kKoBiKS5LD9fxlqF4sMExWMCqv+BbTU
32MOlEBgz69LXuhVQoD+hur0wODGWbIpxVUZQV+HzmHUjVTWzi6BAQsRsj4ffC0mnYezv/apgPQa
vpd+ZU5swBRi5pPQt6Qf7j4k5YMh1k9KpmWcVjHqCggwj4ImaD7YgQWCrZj1fKMYnf60L45qDtjF
JmNJFCfOna8x80zQoBuWz7pp89Lk71jO0Sf+Il8SWONhL1M2uIpOS8u7eQK1/1/+hFCSwvgiH400
l6nf4OEk/IwYd2SDlDwqyzWrYfVHGqjTTJO3Ba2LBQyMsTrhfsVQXGm9lE5iI+37s1xOTuyOXK1J
hiakBoMt+KW1i42pwVp+inGyRA+Vn4Nr0NgYCMtcqMc1TyTjhupLTh8SjVO6jysnI3rTLLsc2Nrz
yHEnlhp9M2kpg5zKd7k8LGnGeV9JRrksUTCkLK8zQ2/QU8rqh5VpEtUHXoxm3m0/yqKT2IoF778e
JnOYPa3Z+6u8eF5dGEVzrReqCM+zHfumS/VPMWJuwdiul4ipiRSWCuN52Qa00qU/zixyFOoV9Oq0
rgXs0k+e1KSGy/Zn1cIC5MheT5qAJvb5q6d8QekEOIuSERnS6C8mqinbkCcnHkb2L5suZAkf3QIb
JL1Ij1e6ieysIsPVFS0p45agOtBde2Kohi6RfVUI1aF6g1CpLpByLtIgXQat23PEjh7ikB7c8Hup
Q5mtEM4YT1V2T41UHgW3kDmUZ60Jwgj14YHnjyvZvcQz8RqzRYnGz6+jCkobblSwJftuk67IKUX0
kVj+OGPEHbrTuk6revXifVJYci1Oj6XRzOtNCxKk1EiyTFE+h5onGKrO+bKm/IUcZmkfjGPbOour
zh0ZlL3IknvbtfxfCDqGf1n1ItDIIlpId/uCAR8uKewf7GqeoGNU11rjjUq099+HsZAYRFifqBta
pewh1B4i2bBxIDw1Jyhor+URhNpBipz8wz5h66D8YRWTOJnhmoyYL2+KLlkRpVDP2vnOphD9fnMh
9o0qM93AAxuLnB1tut5pQDKLmOjMfTWsxA5GTZ1ns4YjijEJ8HWqk9E2eCLTgXvbrtGTeIry0xIN
j9KyVYRGhTfFWTifz+LFuPeMBZ7hKc+Q05UYGFcAuoO5ttGFGMlaNj8Xf/7axX5PyqYmvDDXae4v
ahUzGYcra+KEsvhpxbKrXGxSYksfMjKq1D9M6rAAz8gJpYPxsoalbI3k5+jeYxx29DeJ9TPUsITJ
dzHqwPQJt/njuy3I7PekCDjcUxrU3JaAm8v7K8n6k65yA3voVW6njsD8wo5+9G2V2kcEE4sKTGiI
cXAVgebRbTOSixHTCB0XB+jpywJM4xKysWXx4/TCfhO7qFeA34qKYP9kv4FLnwlnwJBa9xOivRGu
Pa5FLp40sPWAMrfLqqGLk1a8eEMOLU6wlcJooAinHY0hoakzNrx3ND0RrmVPmDBiCR4SfysxfOAN
wZsGAcfDQ+BEZps6p5CqlwliSh9sxCeBXVKYWu9Itu21xa0a20tyxn/pj8taBsZoShEnMF13/JRJ
0KFJ0nP6JvcmU2wppi7S1rHfYb22Jw1kkJAefK8XyK3Kr079ErdZzqA5eqwwy5T2PCp1vYPMI8mL
ALn6MbU2NSkhCARc5IwM0aHdeIoJPMUZGlo7wIc3bhK8/nLtwHOJ2gXbD+UHEq/ljMUeUHFmq5w7
ScmAA5uh7ZRpPIXaYsJlrzzm3gqmqjgVh3reK9I/h3xlXluo77fOuCcLAksHJI9YTbzniEqVl1Gh
zAyR2dh0HZowuyMWuh0Ek7hTwHHpJxuUSoTuhPbjhNCue3DlRTfzUziPtHqdDN4jMnbDK4Kbekcp
vcawmPd2SSa/a5g0m65Z3AqEU5NYa2DwzNBSbHEx7edMcWhGIRjgSQHsDd2sL+EZmZWvAUac8MEy
wwtDsSlMDCTUBGcmtfhLo68zZ9K16p02AZ4JqF3LpmgsyLuRJPcye6989qhGVARtnvh73fR5ATdb
UadMBBPWFHXtV+qc82ZG5Ci2SucNb1l9hSqqBlzz2gYU18ElJMPgI8bk5w8X2FM2MafUuLRAG6fd
VV88JyOLGAnYiJbyMsJnxv003tRv+vKJQPDGgkdnmcwntonjDqXlMYyBEynte22cxMC58N4IiVIv
69jUaiWa5GcWLwvOXOWW+HNkoTLePWUW6QFBFU2Si3W1P28okOLwOc9aoR7kT6GeWTI0RikRmZLq
YRHx87NdZEqlmBAReZaY1F80Z6V/aepRCo7qLOFTJu1oBg3xt89NfujORDYIVr0kfG58wnL4Xdrt
ZXdubo2mM53ZFuAergZCgg+gE9ICNHqRNFTCCf0Ntvu/C8lMqKT3HxpVZMsBX5J/q3XHSymf4wIi
EySrrQiUf9Gwq15KzvNHEKW6nG+2/H0UXgHKZIV+IN847YcnM+jjRY3ffQBrAsf2bcP5haJQTFj7
qprCfBZ4Ys8UA2iOOu6VAQGkUjIWD2cZ91L8iHwLP79uY9B7Q0IIohfE2cOFzDQyrYdGiu/PeyeY
XesPUvxa9aYutmkAyBhs0SGTjXZwCzs0g5GG5QuTVQGygEPKbwExy/k+2IeTUrdBoyuAi9khT0fu
YblqF1+EyT9x3btPeuQKeWNa7p426jx/43qG2SQr7LuQv2UTB/UAcjlWIYeaaM918RCdvoaRVmo4
i09IufstEUDiX/4psAs+nlH5esPAxPuVv9ckgyXNYDSXSecMlrxIZQJIHIgF0iof09wISKpUvO6w
1hjSGbpuOd4HM9VssCJ2/YSl4XE4cdV9RZwW82jtNVpSIFKhI+C7NJHvjhjeVV+yhj08qH3uWhuo
MzUerjoer8VDeo2XKSUXssPKDZ9nw5cSR2hT3xRDK/ytlHBmX2Pp9ysxKqxe6eqDfNISBvURSb47
TGAtxmSnOgmpchIEpmhDqmAnzAn+xsG18CdnV+mgr/nmGJxgauyv/9+C6jOul8/b6+rBH3NjiMwj
rNfAPBGCbk8rLX97/atVHI7tMeQ66xDXM31hX74UcezUuSqFtfvEfR/DYaN49BBjYPxSloJzZ5sQ
TO7bSGDzjxSjlIRZZHTlRNoigOOoruwbzuy9blLRAQge4M6Wy16ncpC7DZwf0w8Qc4951GN2weCN
7xgdXhfFYb/uuPxE3Co/1RgwPt9OPp3h5FhEJ2DdUaICGkVdkkRy6X8OgB6Jo+igxRu2mPJaLcqR
8Sb0o/4bYp+DE6ehHZhef6DIwfTMvLUMda5cCU4jgSBE7WnAZJrGrnNSlw3w3Fnj+tx56djk2Pa8
hL424LZkie/Q9D1usAX5b+5UCctWSR0X7ikA24ACnW5w2l5wlAxBdP0ywJDXJcgqTHppUefGwqLF
1JhVbB38NnQQoOfFElV0T5Nfi4v+LPCAYkawbSd1BVJkFFcL+Tag7MGjPDUL8ZYn00kU6rvrQilL
EXeUhnH1QnF1dAWXrvaWaiXLKWfCahAeEb+hBLLSaTNkVbOdooFeVPoPRI24CIK/xHz4L5mDeg4b
9b9cAPH51ahO28LJ1mRMeESbHeBVaj+EIwy8Kud/LWwCXG/NVrCTRaMmAdQuzvJt7gkQYyFCeCmK
yKtZKso/ZNLNUjAZZaeW8UqicZG/J+DcXmc5RPQu/MdeWu0ycSyKOlWUGFIgisR2BLz+f5uKtlu5
TqwMZH6+5wGcCnPTB4TvFqoNAQ9bKxTVvI13DPp4A/uVHM5e3hY2jQlNv5dXc8N4I+29K1Nqisa1
vYjMYPnyPXSj/6aNAiqmmEWdm64hpyRv5DnULRrvJ7kmXQ3fQlpkr8U/BVqqQUwDcq64C00klJth
0bSVX74fzLwnWfHbxesEdMw7S9Ui0O9opNH3AoOu+yOxcgE5AWRfheqcCei8qVkzGgcg9JmMbc4J
wQ1OJ6AMR8abybKImCDL9Llbxbno5hMoSqXHQGNxxv7R2coz8aICpn+ziAMXmEOmPgkTG19zcgDf
3NNC/LRmjGWTBKOvBWe3bjlfgb2xIEbFc0Bj/8reiqQfyLpJj6cXEam0wEQU8snBg2GGX+EJjQsC
dwsFPNPgnDYbAOlAKd82llIqje6So+iAO73JCJTSKGeUSf0qnxajCiLUphmsuyaHpFGI/PgldneG
izeRESYU1NGqkWfrIHT2yyQJWsZ3VLlzpcb0HzDh4xquLv70WDfbOkg8G1XvpzTZhZTe6+DI7Q7O
WVNNTOWfyvd/NzaEB3IqoKAP1nWKS3+sCb8jk3AwSyW4Pm+WrlpIb7HZpuBEQ30/xx42mNCfz2sJ
5aZE112KNBmMTsaOM36WBmUVAGl4cTYi0C+kafz55STPC70EBPnl2kOS0qDy65ix+aYQYfDovZYM
ZIGlpQx+uSr8hWsUFQ5jRV5q+l4gpcDrQM4Qwca32zcH+NqsMmfZf3xHDJCpVm+kCsIiI8Cj4Eb8
gmC/TCgd0hZGXgo0PFrsHY5Llr+svcfywtb31OoY0iCszu0CoG1jTAQ4/Z8y15ImC/Dk0mdx7MSo
Ah68BaSs6dKxvJIxTD1+AavRN5hw1n+eNpVWiSm8d8+FK/evkhIUKk3cO2yh8sy1mM19heZqDqHX
oF3dDYO/ZW25R7sitoOsS6SYbWMPH7WK/PrTPmDHlyccftL0YLPhK5GdJdrnwJt5BLuYejG4urhr
MWvAGiu+8zBDX0RgB5cPyLSgWmjl3x+V6DZfRPXBJ0eH3GIA/9t8TRhr+EYlF0SjVfM+rem0e0/t
R7J4slAnnd0HeOVo2ANsIqOS8uBktLKkntErjyUsZSdofVtQ06Et4cgArjQWhiUlZDeVzo2JbukQ
GvX6AwQDiIhScUIjOTvUvgtOsVw+bui65TpT4RX3k7ouLPGNEycZXoixKRsRBjYYpWgZO7tc2Sg3
WTP/2ck6x9w8snFAcal7mAjJDgQGkD8AoLK60Nghedf11zR2zJu0EsN7Iz+yAG5cNQPqahaMMX0Q
0/rGgKLjmUEDMOkTKZt7V8lreXD/CzxZSvGIGxEmyRsyAPZaDFHVEybRrddZSLBqmr3Qwn+doWpy
sK7MOqcXiMrjjTXo/rtzS3RdsRRYF1EunlJSpYER5pRi0J2gqRDJN1RzTkeGDYb77pSPhgguu4Wi
yVO0Dh/0fEJG9rd8KnW1FNXU6Lm1qgfNuVvNIlHxkkTOqz6aXxfWP9fnfY2Y+4KOdN4KiIg0Xrcj
u5vq2ixpcI4RgPoFIYbMO3a6Xrn5G94wQehh2Lb9JANBOvULSnHhCdo8mUoCBIH1wZb75np5yJXj
lSSkHXkBi1ajcrraZ20f4qQ48zae7cRWFzo9j7SS8Pua/4aiCeacByA6xx1s929x2x+riICW1qXD
R8obdkjHUE+NaNUN2AS1mK75dcOF/lfBvMGNap5o271+GKVIiIx5z+csun9tEYoVeoWiOt0AlbKD
CMNWkuZ36Lh6hZk4GrER9PMOQxOc21p5CeMiQzAzdJoZFav8uy5RY0fOHtIiUBxGmU6jrgr3AIKx
jwzjVHhrTzw9j3NhnjWCJXOhw33eGIwS9wTfG1my9j2vH8N28PZkubYUJnTiJ0S5XD2urr/zsS4q
5/TmApvh5fx/W7jXO0mZzegViNQGx4W4eqgtjD855O/WI/2WtS36lz2qIlM+JYv1cOLs27q140g8
6JQLJLq0RbHMJikbp2fROIqcKL+I5rbS9kZ0aPU6bE0em3cid6LqC0jSNRmgR87rz7N5KegLIGFN
MqZqOLI=
`pragma protect end_protected
