// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
RLwrboUyQUB/Ph3DGT4MJvoii/Tr1H0vt/k+9iIahYcd4W4EQJvg/S+vOVnV
IgWVcNqRnrFwpbx3FiHrz+rHzO4/zKsGWyMs9Kr76+e/HnvT/rmGhqsXHByb
iSJuvPFF8hgbROW42v0WS/J9ez3qY8TVoKCbFUkRrcCA3wbMhUi+pOWwShxx
n/JzlAOEGSD4kUzjpudhNdiPu3NWjzy8s7Xoy66Alc5m2iSqt0k+rXMT9/AL
3mAQyDR2LEgCc7689sdjtBGTIABrHSIv2ZC7XjZ5IP09jsYHcNGvD6DS416h
1g7Hwjp01bGNX/NDQ2EnlwGJKXhv7fjxPCvVW6tL5w==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
I9A2M4TkaywdRqoNL9GxbiYMR+2TEZygstk0uO2x0rXGc3VfSESFyI1uG/ss
TN+6QdsIsO0NOiM1mMYjvPX8Lgqq3Od66VYKVH73fA2gKbAH5DXxc/GMlBjn
tJjGJGAVzcE2Zxq786dPMGoqOhQ8hQKCeK0hOQKHltw0yXgH+pxGLN55QtUk
/WTbbhy+I5VGPnHN4TrnRRqdmwfvPm94Lc/luHmPrzDy7ek3OdxuSK2jxDCV
2dv4KpSXoKVn3Exkm252FuwW3N6zKs6T7TxzNsRiJ8i0Luxl4KOSFw5TB+5H
TZn6rTYOdnY3coe+2DSnW+SuqNjhDdd6sLu5npoWBQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
R7i85tYBQ2bzsjwLiLz302DnrKlsoIdY1iQhfvy6FwtVSwSCdNcnf2O7FPN8
a7LkBNJPK/RVMuF1AeM74pt68NEu2sZIhgBrWiGVNpPynCj+mOWFaA3Libj7
EzCbl9OE0ogIeY+fsELDIW/QnyINslWRYqNGhr//KNmr+D7Gfzt3k/HaaKXT
KB1YgngdcMR1JUQGmI+2cWSxVxYFTMQme4THCozonTHW8riMZlHAwaJtlEo8
F31RgTEpEE4BUwRNdUSGtwjI4KY4vvYdpfMBzjAb1mXKIJXOWt1Q0tRjvlf+
RRPSy0h0qy/dlWuXhCiKNPzMGH5KzXSiR0QdXL2Edw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
cJpP4uRBuEfUfV0YwLwZX6c8sT2zKmUbg5zsRo1Cb7g3a2QNjQ7/RsSgbC0H
sQ/+PqEdVTTcGQddwQARFknD4Zw9W95ELEF6jNzj/czZgYng/t0Hvpk6EHAb
OJw0vgLo+CJtPaVvHXijStEljInp3WNDflDWrcpmletnY597YXY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Yn0nCcz4KEa93Wh1Pqttu6kyauHKJ9x014wJopT7wUr3xpWEoIMUJVsjfoLC
rJVa4zBLKkp1u2UCM8TkxeEmaKRjPbr+FPaorQi/yP8HbG7OsvBMV2DikI7m
Rd8fTBoc12lZzrrbADCeYLjyRoiYSAqt9pu4zbLpKZ5Wcl9G5ByS4TkBBO3R
b1kVY9LiT9bLOszQul0PWaVPEfV0yZF1gvavevYmd0ud9Wed9ne4sBLOFcZJ
m/IDYKTr1h6CkPakCciJT6MV4EB9IHLHeBBY3QsA35y9VAPyA1UcZgW77xqB
sxrUt0akUZLhq701ppTn38ianaQA5x9lMsAXdKVThgn5QwlTuPGkC72jkg3U
uQBNmHlSY3RdJX2oInNsIcbW0qGubUuqvMjsGpvKLO5HJvE/SkHCbisO0e6M
nDHT8/jR7+356dnk+zwWWimHwg2vSTYbVqfUU25yp7034rVRYBS2fzwsn34t
yshNMyIWU9S2muYvWhMCmxXay5EPcadv


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Edz10Yy219tVs4K4Na/0S/9QL2xHpY0DEffrwjFxBrNPmvFBmJ7SIzhnWNJc
jKp8Vk3jsMxZVGtgNHhVkUlhkfuR2/OfSRD48DB3G1dOo2okYxSO5/haXeDC
ZtCukihfKVlHMOHhTQFG3sieEZ4yPTTdnslQUj7i/K6uO4K+2Wk=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
rzlmtpL5a0ahrxGH+umGPkjzD3Bw/ybfJl724tMRQR2ip+Kx2L5TSSbVm0CW
1ffXKCUIKxkjEnPSdAzFvZVppONfH15g6rFnZnDweEbwGqdkdlYNTejQlbfk
xbhObQGub4VBUNIS53HAEXCwn6vkYcmqAkTZDEhtLJHUWoXBgQw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 3232)
`pragma protect data_block
h3AWRnzov5aHN+d8/wOT9I8eO7PsfVOGW498nu9jISdbjNE5FaIDMoWLXrnP
9tEezTQkMZOkm6x8lAHaCGfTJroSlAulymklUJirHJhmx8p5lzun0uKF+K+l
uAlWEcRmfpmZP6TNg21lP8VO51nNYZ0lkclv083hYFTIyidDcjTVLBYHO+A4
1J69Gt6CqGegeWCTq09nErkfF/eAOYwLh4XKGJUrW7/CffGNMR23lp9X5FrH
Z7QKXOFPPbM4Vzx9RqnDI6OGSFL1iMtfVpNdCoc6NsMqlFNozWk1RDKh+l4h
FjuQPNyb6hNwN0g93FAf3PY34bJEp2zcuAb12ITqF0O41GG9NButbZu7V1ee
XTK94PXO+jYfZwsRMCY02CJl1O9qfi+MKGBGovyLhp6mD97V0WWldi+kkMbk
yq0OlupxQIdI0ffyPx1oU2Goxqo02CCoVm3j8zTA9C0hxDF4A5K8HxHfM2oD
xzj2wRe3ysRbEI/dpa8KjAVcj+0I/Xg7fWCCOz9iYH7V2832RK0q4EO8uaS0
+f8nCgIPk1a+Ci+AgdR+LCZ+HAHAR36jf1YKwZTYn4C+zzNNUvg4iVgnx22q
dec1giHSQs1xEReCChRtmBygmJgahzjaKLEiohhf50+lYI49VoKdx+mXftMq
TOeoXbWM7mw2Wa3VhHSyG6NNUwDQGlPjtsErORFe5/TVQPkrYhESGYtpzXJ3
YLL4BFVTI6c94BXep4HZDGD1GFlKQc0Ofn7+xkGZOYSGH0E63/PljIidoHT1
FQVP2SUc4QgzLEnNGszHZTWhRZ6nd1FVspOq5wlGtNvOhS+jx4Dtjyxco1uE
Ou1z2+ttYhqFpgaNTZK8v+5WipgdbGxiHlbrFDV27Z1E1DigdhkVp6kyG+uF
2LCXgXTPYdVYEj/F63RTLQ9MbfDFIUq+USBWaFHkNqXUQQjZdmCKUUrYxErR
EX3MUZIyZkWuuA+go/uj3C/qS+9iS3oetrDR5e3aOC4JSt7nVckSI64lWsGa
mRj5eu5mPM0xR9EMdh3cY2+Cg0lMkj/WSwTkpmKlvz0J2M5F5RQOndDQppN7
eGDlttJI8yzrLeOSFMeKSEFXPN7ZLQf++lv3Gesq81KrCXkGt65jCfLbL8fe
OmUH0vDernwCbJ2ULWIWV8yYJ2BAjLFCHiMAUATxmZX7ltFb2tCtNBzkUWdc
s64f30rpdPoQ0LxNaFv8Vfn+FEDwk4gdbTv2Hutc33ywCGssn2+A/kdHx8dS
iW1hukUu7JAxTRPbCKYU2ml09wUVdRcJNOBqI4YpDtUQW4AGcPnlnZna9JB1
lq4KvD12xM9A8qXAexsQlKINtPvD29xnV12em+0rpjV25i0vrQRUewXnCEEp
WGESkl04zTlaCqtxJrq7Yj6+dQiABw9FABx9kSdxtVR22HW2AM6yWhBFdW8n
eOX4+cyX0Nii3etO8UHkCROlGPT7IuFCeF3L7oMqjBqnHkaWjr74KNjf9wFY
FpYvOUzq4yIukYHd6FXnJzkBNhXUhb38cvbsNeP/ijM/SJz6iFfb9ds9OIjO
QR4BWCn6K1LyYHGcSDNN9bMoEmY1rhGOSk8ncdpz+KK6+PYbnBDr2KaVNLf7
5QUBtgmbG1FW+YHu/+3MNbXCE4YP3AQCBj29GxOtpcwsc9Hkyum6DdwsjEJx
BfYuWz7M2l+WW3W7bzjVIRbSgtyo6jb38dXdKWq1nhXW+wgE9oJ8Y+w5ueT9
8PCmjowQqk8hPR9l4vn94vYyMqQxdE/o5Hp7dY6S1yhT+GttZ9i85TiYeWBe
4PyjV5T4tThjRUFdzzOl/617g9WJrHPu3KPjrOOvMq4IvxxPfo0kknWDGm2+
rzA4y+T1EHTB601s2/wzAPKRTYrpSKHD/xABnc6Z/U5bTwSvlLvYh0krwPbr
NYw29FnQSYb1NlaSm9IgdkpAhS9c1ZxXbHIu6A3MJWDHNbKM9x6C8Xuh3aU0
Rh8hK8o/pmXYlL3vVvAUIq9j2UfBItLJ5dk+e9jtjo8p/f7oT1y9IoN4bIIb
hBaoDK8vtgoVFiocxSO8lUHFV4HHI5lE01TaUQ+EvV+xFFNbNHkRk48kP+Rm
lQRfO9QYPo1FforskoevEUUpCa5U6vgbMSFjLdViFy6IXwTU3wnZNg1GQ/LU
D1JxLVP3urnyU+cassNEmW8TVaC/Rydvw/dNd4Du65gCqC1uhkS042jcO2ph
S6Qw3gt/3XfAqrhb9Q2zpwihOF3qRyrIl8brAUA2hnYc2i47v0sBGNhaquCY
5ZOXL85VT3ptsZPGBtNf9O6pL169IUgmffTx0s4UJ7FHPk6DmDiBSsyZBWW/
AVR2RbB1bBGXuoZB+YJe2EW2ypV3d5s62lzerZIRqJ/Qb6GKrvEsp8y2fxp4
LJnGOkrvalpFT5aqzbyf2DNeJPgMdCYG0kuvRy0wIrrOyDEDjSMEHJ54hNpg
zvomTtiBY6dxGbs214qlRJsQzGByg1mUqUvrwqEBlx1o/aTbYixmDHIjXP/e
4xUDp+O20/3nD0o/fVQ3CRTULN7ljnn8Lsw5U1SAPUEygXt7DbVCnVAId+LL
wQdCR8Po1iewcM7cXVbJOnW4JlpSGSLaFjJVF6rvrb7r/NMBZhGXojPj4yel
hRU+//BTWxuRC2YxcETq1nbfzWHtP4zXZIeV82tt7h68LYNv870s1wNpuT/c
FudWefYJKrKo+j/jQ1+nIDrLbCxpZc9OEMktEocrCNIx8Sjy0P3FSalucWPY
KtZZpS2MSO+oV+9m7NkRhKETSjbWH7n+tlKj1Xv77XnU8nZwhmYWHPuhwx5N
6TLcXPjctgB1JkW5axXYr3srfj+sxg45xRzRlwnYwcU/FJls22ty7qWjOXCB
uZ6oZcYTYLTe4KLQU5MvwooQXRZLEyTRITRC78ezhTvfK/upt9N18cM1ZrtL
/c+urnAEb1i5wGFwn+wo1uxV2lal2BY1Rf/uDZ0CbDj25fqjfFWYFhHaSgQH
MJZ8sO+ZsWqPOe0GLRO/o3qMFSapX3T9d11YcIFHksEOXQryxiLDXvZG5jSA
qkOvlzt0NVZYHOhPi/Pe4jMXsDnEIF7DhpxegS41IfDtIhrRm9aFp8ssccna
kN4a+w5F5wSC8gXS0yYeSj1UY1oJ4N4Kp18lZgNqSyOxH9gXzagEvUX1rlF2
fQqEsu1GB4Gv4miZfvXCXA9QIp111JJHCiD0tUJwv8UmCp4zOA6D1GFC6It5
cW5dMqlNL/1+XOrLBbyf1NFdSLuLk4hPVV+DDZmAWT+l07XX1DQmS5AQdgGN
kJ5ZUeVh4KBbxqrvhGaNWitHlTEVyiIgcLsDwRt7FZUllHWTrn9U9T4maNq+
zg47BE/Hm8PVeahkVTvupkS5rKgJMukZZYMksGdd7vdVAF7azeoqsABbaAFL
3eO1Yg3JnsOd5O7gG065Mgk3qJGihlgtn+qOGI0SxRtQMgLMgpxUoTkqF+p8
KHszibamI89icMAbooB2tHiO88hBD2cSkp7IpUJNoAnFoRKxdX7CI6/ZOhtE
dd4U1d8uKuDG2m8M47+GqUH9Q50YSpCAP9Mv9dsvZXzAONXKBgtIvmz3jiIg
JlQ1jxe+8lCKATqgj5GBuD9H2snMvJiIQWFap8L/ywkahmqnruLA1+Gk16Yo
3atAVeC9WSzJXmx1jngLQBZBR3Z+Ft0tWmqAtq4+Ul0nSjPFxjPT8Fh8SYqB
JnfzshY6wD7JWbRJVRmfSfzfqDb3YM/5Hj9EEpy9VsRl8Jk5dnMn0ilJZkEZ
bdfM+dHvW2kjDSdLURrPW0YIyKEpbi+cMVdhV+LSCYzNe39JnRYPfzVtWSPC
EzUWRF5YmEoVEnWHRA+AMxsd8a7zBb40G5SWO1EcbdddoGN+avt3NiRw6OlN
Do87XRTtKcPehfi6S+c2O2tOzLqIKkvtEzeqUQS936/13PYJcbmX3inoon4l
7JSafF7m+q610rEL25RogQmcEgDIOCpWEvYS8pYlWuUzI6CeoUJjOvHS0JJr
WJsygwcYnoFxdjwN3myfIGqK2Xi5isE7f4k7uRCHGZw900N/RzqUttOqcx9g
Ggab/WzqMRJvAHqPikbbECsa02WVkB2FWgoUHPp0KMkpf8nUy2S2ax4nAP92
C/Tl2fZwiDMgoRZL8iABx2ZB9YXPZjNxUx2B/YW+49JZpFbW1mneL3qI5eyM
Tbm1ZC+9EW2iBm2kBC1MMnesM8DsBBkwtTHeVDvGsCAjjtQXtEeAPR+wtO8n
QzzF4U+jch0+hyF8m7lwXVJC5OMvFO99kvsQ28aNK8C3LgZLOg==

`pragma protect end_protected
