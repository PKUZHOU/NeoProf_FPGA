// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kC28w9jhHimC9E6AuhRLlMu9Q5rE2Y4N4zwQEGqoGJfVyGE7X4t2nboQzyzR
rBzTGzQ1I5jBnlYpUVb+kppYhk9ptE333Glanog9qP4owUym+biboI7EsCdT
WeE4vfJNXf7qWSjwRdUxZh+hKa96W6ldeYWUTb026IZKDoT7swZ9j8f/uit8
yCLCtOKz8QGGo+QByEe80mqtD1VXwmGWADB6lAVumUHXiBkxL6Qjfi1b1JP6
xwnrdXzu6XqhWts3Sq+27fLmiQ7dGs36bTe4VwLOaQlYlA1jdv8HD2CQobnS
MTHs4ZPXJEXuakakHDoBwXV+bG3qdvWRZ6Py750qtw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KZtvaHDvuW8qHa4Hp95blA5tphMCZejOEE+lYZwZRQxL1929ICfyc5TVlUnO
I9kGFxqyVh7wKIeuJJvY91tEsk7wyHSr33Xr903Hge9NtqIQ+Aj8srK1zdlt
4aHc/CdM4gY1qa7mRVQFxCT7AZnGzOj0Esj025zIFdK+UQDn///z/0lHgNRB
qpk5QnveX68+/nBLUxXtq2PXEv0Q0O02P2MOftDGuKPZR/HsSPxjDvTeRD6y
oZ7WPOlDOhHLc/0/JkcI+KZbE06rs14qeXeCFqDwznTYU4zs8POj0Q7MblAr
z8AGBCq50+nNWe1N2m8+XH8UGhywkn54dMszYiEmKw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
SsY52hpuzAyoVzCifPKYYnqXjYEiLkVT2f8u4jbBN/drOgoUQQS1Bzdk+a9z
5VBsdXIt6uhXx6KvpUXlGM5QbnRDTeiHmgGfECtkNJc+U/NkoS3bGm2OR7rS
MPLUS/kF7N0IPHsbNiuNY/xvIaQhGdl1rO3qMITOx3nW8G6CJe8GcTlE5XRn
6/4xKwUUYM4+UOU5tqTr2LITyDBB2E3mdu0YUj3H0bnmuSqVv4UVhZwfvtEx
fRGOVYYYDUgmPQ/P+YhXHRwEvNg3JVdHB6NRXd41XVRW+C7HIcdheljobpxa
4jqOmVeKo6CRbqac7KUywOyoOQti38XdybVGWX1irA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
aZnzRNN5Z0TVIWD7Rd6AA3fCf5MIFNYWdIlRnlmLr4o87pcowzho4So2pRQY
3/ljHMeJNURH0Qj7NYuPexK3s6v/SaSdOI0qmCvEi1J2go4i6kBXviNkpk8D
2gEXOOC9A4N0x9G1wSC5WD9woz/le2IQIaS8Uh1xlZ82tzZzSSM=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
IDQPCl8qnCmBv+sYwATOtYnvMUfpRJblGrL1RqZsn4mbsEep4Q5K12v2VQod
wZZhnbfSkx/p7KaRDkPBEVtXcGYz1jdia+UcdmriUpoOs1619b+A7TH5x42E
dDRpq4RmeiWr9IhvdRihKDAHwThdHuGt+9bqc+1wCKwCufUtghtVQ+epN55z
0uGncAd6CB3X0ICFKHRoq7wGelsBz8GCYinFplCpWtPSxf9/YSHDOpPcirYe
34oc1L2gRhE97RHyXcfG/Mns/W7I+/AeXnyCAwG1CQqkh6vDIH8bLIr6rFdC
8x2MmtcoSZlo0VVHVHRzY0lGpk2CdCDSfBeC8/4r00Zapv9n/dNTpjYQ7Ydg
qwgZ40LYOi5f1318wGMFe90eFZg/ScXtXgyyz1joYLGnCG3XuOJx+hdP64Dq
2Ecomy8aTm8H0NrAClKGIwPFhnhd+ta6oBLBcFRT5SX9EbNPG9X+vOGW8Hh+
wWA6PiIi49+/df4ccfuW9FNo5nhRRDsU


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
GvRkwV6W6h7oVchhfryv3L6CL5Ffw87dfyEQIOqIuHnfWzNSBeEFZjRm/TgG
ljndnZFhumTVbSKAwJOE+CKWP+a5N9FyIEwSa0Pq+RlJpb4FHpCAQBJ2lb6Y
wFGqsCAnwxNT1xg+W4H2WNT+80AeNxylC4teGGDFvTw/3IgYvy4=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
GCxsQE9NytkSctDj4vJpisuJjJ5KWmC6sDl95M3NTaEKW98iDwGGhQbjgm3X
FEbAtZuI7u77eRocUjaQge/3pFMkt7PXC8vAja6cGrpGo2ZG8TEweFUF6ZVS
DndfpLGTXzovupPhXkhru8QnNOrotMdWVJ2/7zVfKC0wYHMOi+U=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 14240)
`pragma protect data_block
yqB8hXm19ZNhzcuMAuGq98kszksRNg3W3p4vg3Lv1SdiyNuBX0qNuqrhHvqL
9uvnYTCfRFZGlwEqonPlWO7FJQwJH6K5b1umQuMjG7BKcTdtrwaucoRUPwJW
3CVqwfS3FsJGQhz0JOvM+MJw3424nF9H3jJE/SxbUEnwCoyFGjzJEL6zNy+2
YWUNSm5fQieOAIvcXr5T1ucxiE0/Br77kqVNM4Rc1b2ue4eflPZJ3RTLVzHi
7tgRmj+ZwSMP7sUKa6T58x46dW9eIbtR46PXnZBde+lRLroYVMjuz+OtjcCu
J8pJgh/CaaExiAgPmElQOzbBvrLU8iargdVFRMQAg6rF95QnbHuuAITdzgvS
FJdPSND4EwPobFiEX3958ukXdz7xZ09l8Q2BnedW3Q+yMFTzDb7yBHIWlvhX
GKqEY+8Usc0ajpAeJSiTfvry0v/jmDh4OpRaN1RRN5vWoDqZqun9L1SU7FTk
l2VR1zVMUFqvpPpNvNTIRGjJHnBMinlSiqO5NpINvLKY/wauRFeHzA0pusyk
KcFqF1mtOP9olRK1t5TFVg09Yvuk+NDZWIWNCVBGsyMNvHlehvVBDm1NqP9w
enqFzN3RxkiwnPWKLgBkSmI/DvBL/t1E4KmD88mVhzS3iRrRvjAyRsBGVPaG
8dup+QGW78uXoxxN77LF3VBZk2/1ZrqMtr4Zff2+X9dN46EIiNa5clj9aKGY
jWNAfM/BbSufCjLvWowzejDVlVz9ZViWdVimCNIaeypd8ukncS/mWFAvsyQZ
mNr3qqNOVA9YD1A9UehMKIQfdBCjMh2UP40sWvBj9PRZ2q+d0Quono86LrSK
L6x7dVm2SHu/WH9azqdbamYQiqtj4ZTOBJT+FWvMJbhhKi+vIFXTGGJ0ULi5
ZwhKcf6gQc04/uL6a00vecfz8/Ews7w7AU5HVZrFsmcnQJd3tNqP9Ki6TMOe
WYB0AXe3End3TkpGKYjaGrdCRxbVeDCHQdVMbnrV6HjunomYQOLKWc3KsVhG
EAEvWJWXOPulzjN8Tj6c+9gk3723O/OL8x8l/qwXUa0J17kgbhj4m0Py3YPL
c48zqXcbVLfytH8hX95xjCno3nJi/PsxvbIVyf7xudrT3RXIMt/oFKfXxz97
3gbSGQ0tzVrW+8R4okue9mdAOn6fP83JO0l/Tfomu1BAxHWvQPXULzm9ZHdH
H1YM0Don9fkaEFF/dAxvkJQxYWr0yENsYJ0vb13wvS7gQHcbbXDyDWF4ZrPA
Ypl7dPe5NWsyRqIdQHKvZ+W5iaKbDo7iXDhrGZ7y6WzMsGV3B7JExVJyjlpb
GGlONMxPuYxGkqzeIIw5x8NqHeJUWkfaReI5iipBVS6yNZvWKmp59y36dih9
0oCFC0Wf3ysGC/ZIKLNwPRMm9dJUsvxs31h2HPjf/wd6Ev1J3VNPsHGLTopv
hwVXqm4Qx7yIc40sgZZPjK5vbHvg+qUNnr3Zb3EPk9Ar+SsvThCPOBMpr8yh
v1HhzDhZphjR8MdPrUMJHHOqJKsV+kjP9GASrjJrHiDZG9TA0r6D4R+AE15q
3Oy9IbMvq86b87+s6xZll9iLQ3/Z22zL4TQxWJoGnnXM3sndvUHvLNotb2is
X7QMyA8cu6wBhgnxUFeFl51e8MlMyKUapKuKbFSofDKLCbNXoFuXyf0Mu8oT
Uwn9NwGoLNcYcJ4X0vpXBTP23V/tpkZHS2uiyAPknIUZpHjHaSMDcq6ZIKFs
JAR5i3qpzuMEhU08+0NFFxlx+N4BP3l1RYHQ9W5NI+L8FoiCj05Y5TEEPJWH
MbvFKQkPzglZIYC9FodnraIGV+HDarEU7tWDSLLpkMcrFwHuVzd/qjXpivln
fC7QHRtSKsyBG9shvzVbYGIw+S54UXxoTTo82MeCj+WscST0whVwJPVf6Xwl
3XQEWmwciOFy/s7n+GEuHtQMeVHZcJYpfgm0yx1tVkcVA/iBc2UAsNhtm92Q
/l2NnNDpcJ3zjsYOppeytThRI51UtwZM6HdMyRC7uwEXx8pcyyv7DTYFIXTK
cCo4tojLW4z/lQbdHZVqgHhOC8thncI2mlvh1XP0Q5OkpNHUP2uQkwci7erI
ighrw0qEQJ27ZhQRjQ1pb5wD161x+KbI4kTc9Co5CSpcz7ZatUnH5hvHl+7I
mY152aauN5e+lX5F0FqYG02jtpg9TrzF16+t4JfBbF7+EQnGODE64ZlhNiJW
ysmCSjW+uWwarhkiIV8awhecJc+JZpO5vnMN/UAla/CYV6wcADygjqBbOxiq
J+vWxS+IMzyGdLFc29+N2oXEvh0bGEnrdwrT7nLriZ3TijGQhbG/WX06pOj+
zNCJvqHGKEi0Dx9+ihn0ww3Ig6KTMaki5eiV8z1Gu+Bfmu4O/AouOfFmr2jo
tiw2sfyaH/VCx6pqIeYz8pGjEVDz20C5u19VW9nR0F4rdzOYa4eAPNLXcW5M
8Rf/XgD6o2ZBYqGF8twQP3VMYzMrp1cqmEs8XkaX7YLe4l1LaUcv5GnP4pDf
X67tTGokjzXewRDhEQhMLMpriIJj8+fKuTXP/q2DyxV+bUcB0X0C6SXMafxR
VjnTWjczdaoqzC0f4WtGn9C2I2eXnTEnm3yPWnhj6cRWE1cGc1Org2b+AmUc
EHsmN2pTXAH1ICxswgrLU/bCmUqZ7Bw4RIeXW96X+zS38HyiA5kLidR3bwdw
jmVlB9hpkaEvgnAXOmyjdyeCzEOpCfyN/9/SVP5Xg/0mBBKtPkivXNbJVPu6
Hzx072obZQr0RowufQ6YLa7SIKFnAcFNx8DIJ25/dHHbVvee/UUi7FIQdeq1
xosMwDD+mZczYfJks4wG6Q7r5pSBPpmrE0pSjHfT5NVuwfrmYZBUoYkQHQZK
mKyoZJBu41tWgDJhOQiuaopcJjq88a02NgbhvYgP58QSxetb1LirlrkeH8G5
rWDC0xe+Qy78wUQC9NmntVWLPTfGttyiu/cCJgsb+mwJFybj+2FYEKCf50wg
tukw4yT5L6DBeKf+QOH20HQ/JXkbfd0/Edqbum8X7UNJwBt48bm4ZZR/bS1C
Sx/nkx6HvQ2LfTISidPbNdMiJrcbqrspR0VcYE6N9aPxnrmCYNWQ6ru/IOg8
bHyuvMhqgCKhgXNZTaEbZnGxCOcZ3uBHhiHN8KDYnzPNdXkfPdjrMB8iA4up
gNN4sUPoEM5/rvWPP1tNCqvFdVJUICTUWiHtlFJQ5erG+7ayAEm/dIB8tWXH
iXcTkyHTaoliG3qEtUsZRVtxvYBNghs9XfXkUIE7WS1h5n3J+scMbxBRnPbN
OMjYpmS/yEB6lWOJ5p8YVf67uAqf6+Eqs7L9a0d/2snobb06O+oKue/SV0Zz
EosQQyCSfp5LJhhSmYd2tAtvduT+A7IUQ6DshSMqJRnUAWM5juUxO/7k9SJv
Mk/IlsCfv5MyDAAYia1z7j7fvRIhywwMKutNkUhIf2Auzw2QFZEyxSZ5BmBz
LJrfQiuR/Vc79BOZBhOzhCYBkIyR1V/IpZPAVurnAj7aEgRwLTT1Gf/JtdAb
B5VhPeFVEG/8/t2yJM9+ZHvODfIY2NHZKrmf+cJfJrURP1/TkRmabjJC8s49
NyTf5buKKfNb+vHcJBl1pz2I2BFVuSa3D50L3IOb5Onat/Pj9dCn3nZM8893
ALQqKvCfdyN/RSHzZ3Onr0JVd74H/rZ7ry78mbUy/gVJbEw3rQ4jXrW0fgls
zEXQDmB2i/Foh2BndyO1aY2/36RvZaSN9ljEY09ddcLGT4TzxaPpnigqHjOP
YuXAG2IFfyQU0CllRdKDf+p91E5VPjy1loTcEQ40TDfB7ceYPtB22e9VppR4
O5pQ4pwQyp2YvtM1FWSSD9xiMecgpo7l+kQHZwd1sesuVWSoPPVoE/pIT6p7
/uyU1jnSR9wCKUHavImga4CYOhjylDTxxOmTdbp2Q73JnFvJK/L+7j14JsSL
dvsSmXpYsHwws8EQMswjdmr+EiTix0xDSqTsuytkG3D4GF1Tidzcb3khGyOE
sMbNqBus4PuUMvUdcgl3PxDtg1bw9ey8nlxDJYuCbG6Wvv9rm98tYDzGXwJF
35NZ1Jg/Pgje+giX3nxfODvyLFvZs38FlLNvQ0a+0eG5kNe1mAsVymhc5vwa
iENYBT/qPTgDBJBvCFGSdC4DBiYRF+6DoFFWpy5yPE7hb7Vm3R9Y+1RLWQVh
AWqh/1hiS2CtLzA8Z6jG5M7t18lTqMK0teA17VBSPhTTPo3MmBG7dLQkDsxW
DHYzrxQ2nSniK2ye+7Xc+Af4lpcZMeQVw/SuAqRNwDt8mmw9scOBExb/FoIy
xnhsaskomQrwVkciufDGO41AlnxCt8GFovqjC+gp8YEB1+Wl/APGvYhYvjSx
vYLZachiz/v6pdd78L5d3bdRGFxLKmfS247fnxm606O/2ebUEsrRKnuPzZwW
B/TAWy78IT4U7Nl+W1z0c6h3cF4HMNQ/qfsMqnzuRvfxSdxvogwKoiyytoMt
CDwOdPBKmO1VhUJb+pinnTkAFjZQSBbURxXWOwiAGbhlTZIFSZgulZ57NNLg
hGgrr8ykSUJTTzFgy/gDt4+M5tcHfI0gSddB2f52+vvDacjDYqGnKxxW8/ta
ZQGs24pyxwODaoJRhGv7fsnH00PDzKJ8W2rejWb0/YZ+9cKiHlIxrcDuX36f
dMt/+oHQzp1JCujkUC6uvrmMfcY8x5FWhYNf+z6kqk8c9weTflC8kUxbYOmG
uXERK4oVnPiodP04AIy0cTzxh7mwiXNk760xZMJ7dN7W6hX89xPIo/04krH2
XQuta+uyp0Xh8yvbCT73p51DVIrb4JJFSeelPQLDKziO7lmOqgz1LZNJE2d0
bnZsV9+yl8r5OlE36eZR1bn+WeAHQRZzWBgcD+oUKNyzPCspvKxncSr5xQhx
n+IbYbGTkyiR9cm4asRu1sghNtd9XW//bedSzPNtdNTe4DBnqXcGGgCd7wYC
93TSgrIytLPGibvWg0jVsYhc2QwJdo7NTnGknzqrD68dLxqu01A61H0pYv4H
rqwxX+K1KdcWrPopr1jVRt6RyQ0wIq5rTlXhSwUQnhr85r2Lstx1CMlwp7rF
H/6zkm29IN8LDqMG6iPFW/Q9+AZB4NKQOEX2mdP89cVdAKT9PZfzD4S3lHFl
447eW0QN63xc27g822yxAjUDeiDxkcV+Aye7aqRj4qZZtBUhwkB4wY8PG/lN
L3m7NfiwehQxWH3FrEZbQd3oV4xp+2lNMzVA3X6AK+2047fejD7pIKukg/9u
NEpFUCfHo2l10v1acZSt8mLU1+Ms3hZeMd3LO9j5xHDZ/n/NXjXbv6wLOt/R
D/+J0K64MgEe3UO1Idlv8jcvUduzJEJzvAJNH4nH28xsdStvWZyGyu2bSw0j
EG9UAPaaXhuR0lmDO/f4+diTWUDmAdyg7FNFUhKYtPJMo4d52PQh8Mu8NwgE
BHrApJZOubqlfIynOl9pr1SSiNO3C7nK2AnPfMhdkBUSZ1XpyNAda2scnhgG
Rh5rFqNf9QUUKQy9ik3ui7wDN3AeSXHU8hK9ZbksvgVt2VAv9xjXdrPvsQB5
pVHePIN42oy0iTX2lzp3CJ9zz8jcBUbsjaJ6WxUyC6LI/nSvQsX3zaaqL/J2
RPGmXlqfevqEJHJ5eu/TK7MJly7N2AtdziO/tcIRPQ9v7wTGn9yTCnAafVmV
cY19RPRNwHbKHQNRzzHkG9/OM6oPe03Dr/wEnOf3lPfde4NI9Cl7YvC5wE5X
PNIS3vKVxi6cLbqwRnPAxpb5v3+S9FzZOeSlTRuRmj13a/SsauE+xjWetweN
yH0XJ3VsahCw+YMWfiJcVMnZRAQ7LiEVD5ysTeAxTCBQxiHBtfjGIH0F8Wq1
P7Mk1jO7KOaMYK/dXg3fPX/nZQBjaKwG2qwHV6HV7yOd6rSUdOyu1YMdT754
Sfe4khf/jnijzs6cf6X7DDRu5XuhMCmJOb9W1aJmkU/zYby21SUZrOJ34bND
YcVPBzvdmUAGpOQlE/6aVUfDrfnKRHy9DPxb0OotDhdRKh3UCQD69BuZMiUL
m7P+UXfQrRLxBmkhnT9xYrjRjPVbcCTumU/6Z/4BO/dHzmuabYjL75pndOSR
tuApRaJOFK6P/ICHPLdcYfW4tT2m/0KPaVCorLEiqqK06+yP7UHUEY+IrK8r
mcmuUctCsDY9BSC9nj0YyUrhLimIkpEfySCt3r5l3CqMc34KXbOz4TwsADsz
Cw+eVbvBmzrrXanHdIaDoxX6axidrvfX7Ml+jrEuk0e6qbLNvcdurjENTm4h
vHTKcuwiHWpZGzdrglRO7C/cBIv2u92p+CAnYxlilfpX0mHC2pXow4eBs46n
alSKv5awEPvP5xMGI4uxcUpYngs4tVZUPpyp5J8cyb728A3EOiwwRLS1Rqzn
zFQCOz1ihCFpFNQyd4KtYhAMLIsmLK3KGDkHzLMFJxw0f6+wNDXxZQFGHjfa
CURe/o4lc8IdOZslSbU2VNEnS+9Jc2WTDWSFPex0t8xGHzFf9/slmnxjyQFM
/oaquJLJMyvdhL/N4yc2iAh84GncxtfqAiRvpmGaIDdw48QTOaN246oFbp5P
gN3AzadVJ18lSX5f0X9VmHVXlmbdyGmsoVAaCHH2S9jqCMKx00HDuHWvFKK+
2cPU0IO1R0Wgvj15AjyvyIx7VJn8DYpUpJqk2tisTJufW3IaM2k8QIvS4Lii
xid4KBwS6LKn8uHGDn41cWV9HtgYSpjigW+HyQtLrVT6d20zcUPx+xK40Awp
72FXDbD/U9iK5DlpB6DgkuGajrs851WJT8kN7I+A19JigcoJ/o25j4L7emwu
cPKSzlw1NK6X+x2PeV81Fb7AVwwBv/fmn/eoba8ymhe4BoOJsXymWq/lzr4+
u3MQwCqBBzg6CbAB9snuEEWFPnDjargBeEkg+tOAfYNrK9ssVMwXLCDchQSB
Hs1KBS99DIENZ0D4JORbyYlqBO2edP5mmyWFxcbZVzIByQEznO6Ttgd8lnx1
9tJ1oHs1SqjApoTsScPwEKkfdhwNN6xkOlQa6N3EnDRkmRDkAFQ0xq70kVEF
S8pD77FB5DkCqSbIkkU3JnE8n0+kg1sRx/dJDuuswH/uVV/Z0q3+5/AT1XK7
diktyEuLlwW1FJrPMwgCaSkzAWiVRcuKTh8TPyLAo/Cbr/nqNgdauWmOCzGv
trCgTzfCWjfYl+yM96RMWQL8BIVYnGxyPj4kvrlCAQJ2lYdZNyhewTXJwFp0
mHuKM0HzwsnbgfBlyrgurGzufoMEuS1ajB2fkG2bpOqa+QljkhDeDs4ULCvA
Z2TzZ4Pk7HRVsIl31G4yOUcZ3kuoYcoPQl2SjbN12OYUeHPAgW6T46BK5MKw
9V86+s+celt0eotR0Yaz874ofxHKKH7TK+LPzyb+Z31rlIoA7rkAtyejkZoi
iXWdPUE4mqZtjjlVdL7SvLnEW6TSkAe9iw9f0lDwzcB3j/ZUfFWXLvaPMEro
YK5NGIMWxuu8fcnwtnkOTzmsJilXcUCU4lqVAQB0Ym/mOu6pS6QwK0De/Z50
WbGdVYoJUzB/Xyywg2EnJprQ4ayEFoJglefaCzazvl0TLEDrBSPoZ8fYOhEh
aSVnim19l2BDPqvo/KALTm/XtSWTmhUnQ0fDU8ayaErbNlw0zzs08lsVaju8
usiLHb/fRai9TdmAu2G4s6NlmGrHXZ4Qe3SbbD+ifEhgkg5nPXlEADz3obX7
ciNIoPPXHlB40LyKvrpmeHrW0b3MhJ2TGZTPsfoV4/hJYDxDwpqxeGjTWLqY
YYdvKJtXf7ijFwE1ebtR/MeGvHDnqj0UFsWsoQ1y7KV3sigQyjr3ZzrIuJTg
OYw59UBPWBB/JqUZDiHlqsqFoBSPRlHSbU39+1oByO34bvTlWcteiWHmgHOi
oWrl+Q2JmHlYgRXmuFQNRXSQkCyxBbKqO9MUXr1zwPB17OJinyjmmtS4wv8g
jDqQDPVNVvqaPui94xNKfgGSM5OPKU1Wf2U0BKH/+nJq1YjezzvKc8wmOckD
IEISYagH3oYb2RXqO29Gwz01X6/FN3OhOSxfIUnr+igp3Bk37PYyqJkGSfAQ
kYbiWa0ZBpqZqMOKC7DsFUCjjdTuxtzPmBdnvlI6B2XVgDX068yfZbXPdI5j
oXw0BhqoXPdRisv6t32vklUzPDhNWxxzqOThM8ZI4y6fXsxEaDAf6/U3bK6D
DP7Tk7nYtYA4qsMruiNKbUzvM9jVWhGg7pNoPC0xf/x239eEpwMj6mVtuLy3
4IAOafOnhO6ipheU2//PuLMtIW91fsSxhoGEUJ7/OJssSkOjzTrfq7BpD61J
4EXx8wEunKb9pOt0m+r1ZAIXzLTGQ8/9mXJ7tZulLpgsamijtvYVj9+MlMfJ
2wKlByqwcXX9C+j7QIH3Am+xnD6SQRSLgHzNeYpbeXFVoz4EOjnL4xlu8jmi
yGxsZ1isSodapdGeO/bFTpFqALOydcKj+s++zk3DYFqjnSL4IzYW7aloayyH
10pFmL8wR6VN3T5s4XybvKDoYmddYtGIJ/Hz0d9EpRkxnpMSq/Ak8JnxlqvE
yE2XnrbMXc26y1ea/q4iMFmifdzpBZH2J6KaP/hlsMfHjmQ8+PITBlRpu/iZ
897c6cM+SBQ8WEh+H7npd570/bbR3bShX41oAprTf6/9sBniYc3S3BBpNK53
x9J8YH217ZPORHZ8oUZ/lGKfxeTDuiz2aVRkLLklHdWeKEU3STcSNHFRVDwi
t4pVukAP/OYYrMD7saxl3j4oNP0uhSE1Gknjytooo49zSTIB2ymcpYvLKQIi
vauvamuJ+RMg4c2P1BinnIs6Zql4+BNQGAs8aBGF/vZ+cEYL7bw5Vfdc0Hrp
xmWkMyBjYO1W792KzjWWfPjYRmpzn2VndPB2B4tXNfnMV8YVUZGrkUWLrvaH
hAZuhRRTL9U6V/03JOXMiWw/xhaQZvLND08td3mpez3LDgTVCd4JDNKnc90b
CfTut6YgRk0HSG31mkjwm9m6lpaDkpN3IDigTjGDzxRGZNYgjmPTnb5KuhGM
6/mYTRbbRbaVsjZy8O4r5GrqWFqv4zwzvN12rhgqTXNlAEAJMSLyvTT07ODQ
+/iISxJDpeJlj6uITLMSA4sDGYr/gL7bW3ATzk/YP4BBWDh5+9W5I9sRcSVo
/yISnjKOFDT7Sk9q1wCco7QTLtzAY4KbbWHb1t7fb7HvR1gv12fumHVUSkHi
NTQ95H61YDIJ/u9HOUzKu5aES4kUhf4CatNFSZDNxN+4B7u/RMZSSpTlIxja
34kQe0fX0atrI5BNDeemBI9GFknFLMxAqqhQ81s3CVgOuCcUHX9Jel65j0C9
33PV17oFGg+k+C0TQieCmMYvrQMnzJDOsj38b4Mx31LuNnRboRLiAS+8i89C
hDH7EQMSU/TtuPKqimvsFHEbhoAfKUjk40giC1yTKUc6P+zAL7ZYNSX8af+r
pDOg1r/fcHJbDvdexgfoT0oPevItYMbKKkW2Gqk2m1xOUTN6YZnDfobj0CZ/
I3rvqlfkRXRxSNL8lKi5I+ExT2gRqpbhN6m1q8tNiF7p3R3vRtENagYKtIJZ
zOq/Wv3Xw4dkZCzizUBGNQD6PGVaLnovhJG3VGYWkSNnKuhnQHaVlYzKCgxr
t3WP+vbahKV6tN20upLhUAioFU6jmx5vB/uuYYuDwONhfVmgJz/Wd8Q5OycB
h4Yuek/ULE73zbkqqqscGDG1yxOVABA7dV2+fItXlzRZLmvLbo8gO6K2xunQ
M8QTJan21rj+k6uQzNhtk0fL7k3oY+zUvcV8vIqNZWvbqfmyang+avK9Rixp
LS9LmKQr9mHCzQ5oTrIXV/UhRvzV5zyHs8o3rV4kMaZgY21rXDcvF27rlRe3
TlcUalChtUcVHPxDGUabJkRS7mWopYFYZG0BsflZHGlMPqod10x4tjNo+Z9v
aJrfd/or24LH6Re+yN2/jU6F4yKVm7YcgK9JpTKhqb3mZLFmy6Rya4xlwdlQ
6xySYxUT09nCGtyu7oQJGm+s6ObcEk0NHxIilY5gR11XczcPtvWgp9f3dON0
S+OaaChadkvYiD5Y+fqtt84ssnN9uqIO0XiWNbARySOyxMjj7ig6UgczJjtg
rrn492bgkaUMPxUWOggOnQM82ntN2WI+6NTzb0hVhGf+8XSBIGlQUmwdKAp7
rSsE8rTPe3zB17RVD7xqyUbFF3YHxegO4QyHLoRw27Bbf2KEwUOxXq4x0Cvm
2vCju+RHOWNFLkh/kNLTUBZOrVE/6nEo/YPwiq4TrkajuKVeuRmHxwTSzSbF
6+APc3JithmXoaDxx6Ohz2etT0X219iUlirlATgAUc+Zgs20LHzz65zUJdRA
MUIHhWm1WpmFB4eXtSDskoWmTL0tHlBRrmvQ0Zbhm0fdYGQkU+s5+URgL1LG
krEZ/QVAbDW625MaGET1riJdEaPUx68XPJRmwtLZZ0QFUUKCbYypzeKdWMBl
U1hoBqahVUgFs5mFzOD+rHBmJMLq5S4SM+Tjgv5k2yEsymmnMdN48JJM1wyB
5bOyAo/lciFG16gTicLTcNQ6oTWAa+RggU5i9tvDsAq3oCl8y7MfmD9AGRU4
eG/+rMdHs0rkJf7//+bLW7n5K0lB9+RI+iwNfZ5EJO7786k3phckr0pxLxbJ
O8p2k8aFM8R8gMJEpxGzJI2HQnNBW4QJC/Dl9r5KrsUHSvsXsi/ofs0oiC5+
DmgnUdMJ/1jA1FqcdP+xHKY2wFGetY4XCJgpcarC7qBz5J9CjA1Ue0w3o/ZQ
AjdL9xLtwqFviZUxqUXrx76J76rnbPJsOJKCnHTZvKFhOH5E9y1+H4VRnkIY
EEY06hYGoqgs7f7W+HAC9LI7WYeXXRVwoZgP9qkX2VSPXdaeURRnuFzD1Ra2
QmNXa7PTh15obdUct/qEaHIMt4T1zwBAdsjbplMSBCY9u8ylJsL7YIKub0xa
12USCMzZhz6KBACc9rAuZbHUcRtCU8eCqGFs5VeOFWbU2hQSWCDJ5C9lpy3L
+NDgvPiYQwCKKo6Lhgf5M0wP2b/BVi6akxcWKgrkTSNO484NdtQgH+WlRtHo
DTreB1BYYVd8pvL8eBg/NtVWfMOa9oXPqoqdAp9jUME8ckqohQgC5UprV4AR
nJuozYf1vQjJTeIxdhu8deTLaxt9RxaYfkzcz+uzMSxzLRe983lGH0H9DpkS
g/OJu97+kKdAd7Ep4mQKeLUnNgRx6QpwEP+7ff1Az4jwxOWyxg1/iD67H0Fy
6fQSqhaXUZ83rJSOFdyTCb5NYlwRfWPTnKa+6H4QyhXj5tW0kDALE/a67V8/
7luRCz61ZFCoe2lpy1FePuySPNpb9AXDsO+w13x8sutBoMSDRtH/3qNfCOhi
FWGo2wvF8HKU+Gv+UKSydszo4UdgbknwQ1hACj192X1UPsKMwKrt9/7k0IPE
0wFmd1xdEjULlmvLy7dXceF+VMg5Xp5AUFqkZ+5BW7gKKY3r8SSwU6JSi75A
3fVrAXdblrTOG9ubg3xPNGwYtUBpunaakmpygN511gFfjNIK9iOXIN2CeoCI
XaHqrWmWfmthKg9I99SmTKP2pPzSM5hDxkP34XcVUNqmSkCfrfSVpoF5o2bp
bP7JEiF5x+S3pCdWbhz12lOOFubqvMKb2IpfsbAQ/34YkeqHlJhbMFBAHYdt
3siLuaV/my3btE4jedwlnfmcNKoLQRiX8zY2zvU1JHbO4HFjr0J0zIv7B+4s
RAXMxeTzH4XKbZ4xQR9NogwVojiPfY2Nv/aKDJlSACDB/Jq8fZQtGYf0eB9G
iLTMMH24JHWEvoQd7Q2ho7PS8r597W8qQ4amdaKa1N5sU/SHkn5esOs/yewD
yz9JI3hJoF0MJWMWax5BHe4T2g4Cj3okLnImpYnCnjGidm4aC1zwdkclWQOG
Ci52vVrF3aTIFuzZyKIWEjOQy0UEq7F53IIkqnI/Zr/47IkKFBh/Psz5ipZO
Pim+j0HCcNOCMmi83K2hpZ8RE5r1SR3wTlOChyoOcDFFoel6KS3Boy+yfNvB
Q3PULwHFKkkZt6bCiIMfgwJmNkIngNk5zJlfsc2oO1e542JqUg6tIqmlp01G
AM6X0YaHnLfDEWI+bXG4GOeXYHi/5M2naSPpYSOCkCFVVLMJpMpYPB/hj+m/
mzy8w61VEd/3SYZpwPlc2qbPuY4lKH9U0pzz9xu5PYC+ijF5i+DSimJKZ6qH
DYkj0pYc1GjKWl9ymVYPOU5zRAOOzO9P/a2iot7Dm+9Y0nf29tm3i3gp/nGn
CyAh88aAy94ogHoDX/+HAWsaKdSE3emCze1bJtGILUpFKi+8ogWiD3lvpno9
1jqNI3RPxYZxLv2WFGjnXeK45Bink2LnI0aFsGWxm1Dr5DNYrPNf6PnruISq
O9CrQD3krOvyePmkcJ+/nWfkkoRz3mm9sBL7Tp53T8Jt9COYFstNIA4AB/7s
Oi5Ap3+scdWq2q/7ljcD7lMRa8Ji7wfJVmd1TWq1Jy+OrgWEYoaOQGUNIFhR
ND32opfAwFbsWraHuHOmXfqpcH6VXNdOhcv3yGhxkEwyOini1ny4eYYxigX9
4SBfYAzc2w0RSWZHJuZshkPer3d+enHBAiUszvgrvs/0eu9KTn3HOUZQjQGT
1WMMMqLPAZBDFfqPhlWTXZzscyWLMej64EuGud6iCHYdd0cjeDOA9wi4TJio
q0iN+xkaFUXzzTeMREajLojsG8P+gDvO9asRStcuPNkP9gLKvQ0MWtSFfVMe
yuVqzC3f3u4z4fVt2xvML3r/bZrHRI+09YZNorVoIBseMXXnJnShyVVoLsfm
n4ByugVb1WDcqkRW3875f6RCugUWIesTEuCUGyRWzZHxBOr9aacUvP7QDScx
2kVhUzlmxYcFMxZg1m0yoQG4satGNwuUpO9aFNqUgD3urUXsRhPTU8h58Brk
oPGpCv28Rs9EacMPmDck9sm7pYX8GOphYQVkYu21o8nOB1LvGFoua7zu5MFF
/GMjS9bWXlNFoF9JDcujIt7UQ8reQcdC9W0f6XZ4saPVqy6iZ9pCts1QkRPx
utUhArPwLBTY2VhV6zlE2MyCKMjmJVMJmxBcPw8AAOHGqcHFsVv0P2Hm/5yl
j6BwFok0fxkZkXyCx4DDsOcNBK9eO2tdFVfa5/nMhiFesrOgez8Cbb9Ir9Ir
NLK4jhbb7d9A+kicBN8rkQJGkkHCGegJudYFB6IwNabdogJlZZHLVF9PRCJv
PN3aGHJ7RYpe6h9dSQYckJ560K8BxeOtXVp49gmyq7+E9dmAYiF6/SgSAIkt
yHtWpJteCwg7276hIZIrmSskh6sdlPodi6QqgFf0h44GFbUo8aGayqGDGMzK
wPeRizh42Ghi75A8HPdEFa2RJbFyc8Zcvph1i9ywguy9vsD4o2SP/R4ELDLK
rQUFYOVOfdPKlAhJSBTYnRDc8Y4NWau/sBCqA3Mh0i/jP0JEE54K6bXf4eSI
DlZ6rjBC60EP48d7GJtH7IVf1myuGUAvQIEtXDX1dalYN1C3+TVk/ERJ822R
Q4+zJVSs1G44ezMoFHtZuOqYn0KSLG3MVcTY3NP80o058RaTV0/rElwAGTMs
mr0TdVxgjE9Ypa7IbAX8PqeeA0mkHDISHrIxq7lLaXUQA/mioLTeDx2vcVHE
W9Y2Ojms9DfTzj6Pc1zohUlhqUeUy/iwZ5lu7SSuU+z4l+rb4S26skSH5XYp
zD2qZw6lHgL0ADzDpMKXd2rdtrh5/hDYZWt/REuFyRugq/ej8zf2CVzjeWuU
K7j4tBtUdvTPDtek/wlm3YLOhiXTTwyUw5kVYhUV4kH9BVzAMguLO79bixKW
jK12J781zpHfk9sNfYusQzp3KCCC5yhT7Nc68Kc3V7v341Hiq+p9hqCtco8w
Uh1Cek0flwK0BQZ68rMLOhvC0RZbv1WHTUv1iGykVsLHf2z/61lBnFfrEBeF
ln2tHUxZlvRdYg0PeHJry4v5oLPwaFC2LffZTKjNIY0bWqtAlc4OV6/DmYx2
Z9csQwrzv55tGIwuMKUrFfXPj54nJm74UooR0ehYTGaPkrLpMswCgE3UN7JK
daRPzlqO+PNS2QZ11lWLpPTmZnrBgmJ2BN7fOtPP5Pn0A8C+k4L8FpRo/cd9
NLpeHCJ1N943i4p9jWRAknkwkR8Y3VU57tVYD6qmsEnLQt4oWxsvHTm8ND0z
A4QP9BBPAK0oHDnqb9IOyHV2V3pHsOtn+mlN25IJtIOgPCdqmmRlD92XJzGd
7ImZ9d8DR9jR/SRKrbFkr0g5jG8lgdqD7RNF3Oxbew73SHOnaz50aaFZLQ5G
3Rqpp4bcsu4uKoSn74coczzLtt2je6NkfMfJP3l5UGanepxyV8dhHzb1BxJf
YpI5q7p5NEc36dgQGefLa4dUynQJQgC3obgYj5WwKtd5vE7cF0NPZjYYOZHc
JfL6Ucdbjdj4whrcbR5D0oQ+0MObd1frHK1zW9XeYbHsKVIRsTMkwl1B8dUk
itCvkEhsJSiRbKK43vIFRtAW7EvTo7tRv/FbisizwuSFhIKoI+ec8YSHa9ay
YX247vkqtUIKhBUvGFhD1KvNs9i3PaYpInniEHH/4EZnaoKY4kopZk4bQiOK
rNiKvk8RyBn58iS0MRqMQAVJIl+P67Mo6npICLMjLGHh6a2RuySgmKjleEBT
6pAwBHmc531K32z+CEvpsKp08yR5JF4nrUKLFAxj8wz9YAzQGQOIzTDsrJG+
0bPYfmcujOQ8bUIhunZJeXaz2H+RwkVQuGCl696JALuNJ/YjnVI0yUcIEgNr
GpYBonImJIO/orUgwaKKVryAAwPJjFOEV9gQIWliSg1iGtV1GqNY07RVz9b3
LORQTWOQ7sp1xxGPUbPHcj2sAeFBA27FIekECVbcy99gfEEZWc4FZyUC4uAz
Tac1UMRae3ewvTHCzo/TpJBVvuCu40YGmVO7v9wVePd/cX5dEwgCxGZIeoYs
srMAIColrPoJ4t3Ac+s2EhqWPxpwa5fUvedDLCK2eEyTGaXbAOuN1TBzVL3A
AMmzez4CQ2wf/boULquplzh8h6ywBEtflnmiYtjZhROxQk9FYHcp0PAzbUPc
AsLhtjE1Kn8+up33zzADLnYgRb8yP6JUqs7kAakuC/ExnnDfoT+CrK00wxeq
xBDostkNiQVxzMWWgYrfMzPe+wJPTAg+bmWEnbeB6kCnfk+YK2TVuFIy2o2z
z5QbXtZ6IQk3zMTSGiuaPzVLkT2qIWA7S5dHFO9Sob0BAgaTLsPyeZA21k89
AIE9+1RETN+0E7DEi3JfYtZayrcAqLaQtrFzUhRFpvQEWIDQj5aExZs+1mRL
Ziy7v9IrNCmRQWSJBeYA0Fi128S+rdbmhsbcLo0DcCGmgOROBbFXH68lKc3g
73+zCXAKAHhXb1s5sUSX5odXv5z3jUyBLEqhAEZL/39DAYMxkCoBNnGiY/Kl
RN4q0C5wv0+VpFBJN9iKim+9EucR/QnVztmZqUv1F0zjmohD2xx6t9XXNCdC
9macIr7sc4o0hr6R2j9rQnOUk+MyCR8xegPtKc4yFO2nT4MlYweA8KnGqw2t
RDGBu8xE5FY+IoAHcTqWl6hYvox05sh7Gy/988AkIsh9RkOfcKr71kjNgZR9
6h+OA7iC9XfiIFfhBDDJRZshjBRsD4qm4ml3kevCpZSJKjE8e6MHE6apmfr9
x9wwGw1FvNlIRrB3RXVCK/esFa0+EjCwNDjfN9wl40OJ6a7OfBz+V0SOc/Oq
e3y1QYdfHitW17uJ0VemmEKMXf2JZWOLaIr9i8rUA3OFB5NgPzFBfQm6UQf+
5zD/b2YiEyZKiL6yubPTqS5+k4X0BTUaFTDHG1qNPnPJbXMh0/bQTARaMemA
w9q0CEgyS/1nSsK9F9YPBMajxho9c7k/M6JwHFKqdjems7eQugJc3K9yLuGG
uRs9clRr3LBD9ehZ5Be9OXulDdpdYYsXf63kX3AOKk0AZtE5ZOqxSSHzcBaz
yZ9N9VgUF2sLOLGrzdmS3SyHGgK+uE3ZUDwvqsqB9lPvFRRzY+JBEv56vpZl
9bM/nuC+YfFSLe+9SYTo0WjWH2EIoYhCctqf6jjkxzybRHNbgihDsPv4X5Rf
dtt9bcjw/YWldl62lqoaE+iusiP4Q/MqW6rhGQETkQbVXfgVtcR4yCE7w9M4
Sla4GPanQIPAIZh8pR35lG9y7DH+yg3rHuAF4fS+7/e6rXG8F7NrBvBUdevZ
LAJMkZ+GFx/BLTdxdeoDcrljEQZF/Vic/OFWdgt7qrHt9y3crB6fCx5pPHrA
EpBqijW9KRebpXbTxHxRfHyMURGLX1KfPIjI/AJt+B4f7Enudv+jF1xViGW2
oDYNYdxF7QONak+GCQG1tM5XlOnAtk1MW/+0Sjrd6MvxwUaxdfLxFa1IMTEK
6JJBb9jGvCwqxyRBFiV/92zdSBoEOGjq1x2pL6Z6x6MgtXlzvePfAH7GxAjV
1JgkmAIUg9Fk8HTBXoDAzLbqsQlmVxqIkLjTf6FuywGH398PVuCB4Uei/2tL
NgQL9QFw0ZLOwvqyjThvqCmPTMmj3Wp6iGPHQOUPuj1Oy80CvkcoKhmObh6y
L0G2TiL6oscHjyMPQhlVpvnhOZyJ6/fmeZJAKRC9I82aJ+5cRKFMsd8iZUbn
czgY7V+Lwoi56eAKh29Qad2Dxy6B7AuTat68jenn13AkSwClJuqLeuj3IRDO
0t3cbFMN5tIsLtgy60Ovklv8ien5iZsK1Qyr2nM9xZoCkirxjf4aCYS+rwJy
CTvoekWiZwunI29pBSW7ad1RJHbCsZa63BvSrsWb9KiSwwOzVoeHd4i54kNK
OK7RfTySulIRuVZvVdxmywAvIYVG4EZdZggGl/IhAfV+KVTxxvoD1xUfLUIv
JNs689owNkd6D1SmEu25pbkSsxxJg7wTvBqz+tOzPbm5NxPP4oNceBLvOHEo
mP7H3eg4Z6JT7TwRDjk+94cqeN/C6ZuS3pLjMFgJLVBc6NblyV0voYKIJHHY
WmZUtpfHCz70L7RnHo/36tGodXkutA7vl8hYjCGiFvhfA6ytlWxq0+pcNUu1
1me2O/JUBWeBy1tHb2sxpIaKtchNzWvj1bolyUqXLRpV8gdQf7OWmIUeKCKq
L5H6jSjTOnPMwwNZO0tobKjfv7OBK1mk1TleBoKmj6PB8IUdan4ErbxeWzZk
kTfC1JER3NdoHvFRkBtHR0Hw7XWKbCPIOUXVzLU5fKwQN9CnG7MnP2XLzZGA
YHGCZPtfWw21wBDIsamtznZIk7bKujnbs+zYT39NvrwFLFnzijdA5ngyhqZm
Ut2yn8DUyLKXkdkwR8JoyS7voBy0BPmfDRPVEPOKC5QklDc/zslWUf+77/4Y
hRFGrmtN/wUD/quH+AMj4+RDu5ZYzUQNd9DJry+bC/9ZvZOMMONVp4WqrZEw
kcuEol6CX2fHUdVrSQ9JwmYEhTnQFrecqMNSkZUbxn5IrbvrQA5S6dDLyj6k
f0iUfuDXiiusGnSY3BsRC4zHR89ziTMnYEqW1MZkIclAdDbjQjDYsgwFi5Nn
qsioLxupXxW1chbdw7AIPDhmrU9ggarKFvm2FZvM0jvcU1WJPleX8jiN3/9a
fhIZ0+ClKLZQSoMZehXzg/A7GYxFqH2xhy/pDa9jHKqdmbE02WyJZ5RWZ43h
E+DTvW9cZsoRsL1wJWAlEOYANneP/w9Th5mjDUzem943qADb65JIkA6ZX1Tv
2u1LFdysM7OGmOv+hbkcggUcwTsmAEgGzwFfTv7q1pqpNtAkeD52CGR+m8Tj
Qoyauhw+9UvgRoQlYIdFjdBMngCuKmeRQr5N1xl34G4rj4afjL9VLn76Zlob
F8jbX46y/qbFVwgNWANbmPn5xUz4ZNGDvAUgb9xmcDg6QqF+ZLOCBH3zFTcs
5gJF6FoaEo6B0pYDFPNTx6NsIgSzVfLsL9VzGOydZ5sKJtNdqJs6RqqYGWOT
PwK9wTB5vaTPSWA/OAuhB6dzBC9oNwqnB6DopUNqNlNnzkCKcnJZ1KWhzDsR
QktSYNYnObaFzmDI2JqIPWOikFVWqyWOway6vFoP/ohKDT7ZUmxlBzXjIjnG
wxpc02sJL9391uTU9aODuPwkzrzCBNdb1hvYW0+Q43SU+NAV2UmDK9wnFXCB
xciIK8pM25L8DR+vRtujzXpba0qoDwHzUzb//MMYgNw/D5OQ5o0ZEhDaSy/B
XKqw6pyy4EsawoIcx1oKq4ov5UlVSPCttraLbjysmUSDe33RgW1YQKc6I/Fr
ksEeLljDzzS2cXxfmyJ2IrM3LMJWwrpYcepAq4V9fWlwFI83KJkt/BfUkFwX
xTxhdG0JWN6Ytp8UdjzAnsPCs7hi0HSgMIEBp4l7shoiSN0UAitko5W24vzq
tN3pbViGz1NzapsYrUyMgw5BShNt38ceFPNrEbcl5kTMt688XnClcbTOgwDt
3IC2BfbzSc3usjpuZXnF4y76pIKfSD9Td+7Bztr4dQr3ck8pUfrNOKHJr8zn
9zxMbbm3CXclQedy+VsQgtMJgYc5B2fko/LgWhdXhdq69Rtx8SfhyXRDABOI
/0XEOanSAawMWHgIzFplGF123Q7Q+Fvg1WxsbdahurgeYGVrpT3CuO1L4IVV
HgtUXv5w8E9C/lvKpTC9kJn4xioViXQ/1gNJ3jOI50yN6Xbad7FmB6Q1ydEw
udqMwPqvxpBwb3GaD4bDQL5lmh1HTUGKY3dhPncLNltSVMj9/XhTdaFDXUk9
rJyv3kkdb/dAsM8L0vJ1yXMURLy6sZKJ5XhdI8ZKSe/ovQS6Y+45iTWLGGvu
x7P/mc62tC3arv5OiOBsbfEbbHBp5aT7AnuNoDdyzvR3U72mK9knfYctrpo1
4npcfUGmZAM2sg4cjNyQ0Y6Jkpul0i+TKtbQUUiIIfLq3gk5DwiSvY+s7Q8M
2u2Le+Cr9y/s23hTEZN1RfVDDXE=

`pragma protect end_protected
