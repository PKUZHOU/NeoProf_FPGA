// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
5iaf5wHzn8WrzC2YFwbrzFM7/jXN7NlK2A8AVsfSXaYgqYbLOryRclj1yHm9dDrq
ch3JxJ5QnnMysojXlbENU1s9Uo+4ipUqmbjfhnNggdwTlullYlpCpp6CnNu9xERS
TKS0GHzcY/b1bIZlYhCEo5hGiYPKu2k95iGsR+A8loxBeyZA8KX1rw==
//pragma protect end_key_block
//pragma protect digest_block
TVW2CstXi6x1++uROKXNFHfbNAE=
//pragma protect end_digest_block
//pragma protect data_block
FOzL61Cu+wXtzIcgBAm75TQ2WfwJrXNH7pMCjLzclseQqOazL2qMY0bp8dHtdocC
g0Oa91nrQ5U7RW95w2rNK93AV4ecdRz9R+rJChe7A39ltQ1qhXcnk34NWU71HMfQ
0ELEQiREHQ0eRvq1Q0i+i7Vm+DPgLuaithwirL5w2kBy3dg14KZvxifPgNdGfKme
sExPjbfLC+BJaFW1q0WRGGsTLoJIPLnElbeeG/UawibUcZthmtTpFoTcKr0gHGrw
FufSNIDIYDz/O3Q5cnF2y+KaLByBrJwjVA5KSck8sSXnGMD/WD0CxeJMPVRo1Yf0
xTqdXuuQpR4DoD2G2OjgHFovKwAKeAump4dh1GvIonXcnCUezB8igEWHqCYTUOt8
mRhw+R2ermhFvPrdkFr6XOgaZwQXZk65curIz7A2fjuORwUDqkqLM8F6SpfrJhoA
1ry/QUlriVJ4xo5f7ZXN0dXSAQ35BwnDkzh+Pe4nDoR/p6lRcJRYmWlD2hbTyeNC
ZE1mhGIxcXrXj8z4xgnF7SyYKmQ+1aJBQ3OPyNVE0HRORxUKXXauLugHaL2x68Mh
djiD19cRT5J36jYoYfOwDoOmEy14nyEGleua9cmz3lLvLErq/L6WVGeot26yoqAM
y4p5C9NnFyEhKUjqIaN/xTWFWHLwutsiIBdPrCQsRhoiw0FKfxRXnFrJaqFtOK9I
x6vYd+k+iw0D6Vz7DyTYqq9RB8LTrUU6QaIqga5bAU9539X/zcS12A4b6ceVM/nY
qvmpWnmBcZEwI4Zof/mmccK8u4eQ+Cv9NmUTlGyho4BHuuZ19o0+BI04Pk9PIA05
mSp7ThWPT3r5sDK2GilzCN8vXK7Bi02G6ItuoBjA2m+9Mgom6ASYg8kxec8MNamw
3NWWtOj/f626HZvPM9bDOvt/aydA4hDUHOCFNMhuVRhARKu+vXA7SLLTAn+eJXM/
fzz6b8d7Hh8KiGDWa9frQoqNc+Qk0sPWPlCXQdRECyoJt2TCwNyRB7tcZFzGUvk5
woVR70f0ESrtyoMO/pBtAyTO+mJveZDBoRv5coozTJ8OUNEN/V2gFKV9o5IFx89I
5LlO6xNxUKaRWMUFZCCBW5hsUvcr8ChzWS+37N7XjEvbmRgRmSc2PBKCUYxl0Poe
vKZK5A1wyFUhcQbgAIQxo1H4u+HzGxP0XUaG/3Ng5XylD6kGYveGYZ21l3grTJH9
/jsoMRE2aR9R1mlyM7kHvK5wpA+0kOpaulm/GMcLDXU7LaLQavBBxSIgOEd2M3Gq
ZF/OVKwgwKgKCMQABOiBIwdn6AKnwYvGLKjLH2RscJ471m1BcDa1HlrUxkwkfw9L
hG1I11PuaYX6Rg8BSOgoe0SPzLM9tZMDuSjC7yZsPl2IgxgkVhfzKPZxmouPh0j4
t8p8OtfQy612+9t5AknLn4QxnbaNFILTRb+stO0WFFUtN0tRGTuoDYiDxi3vplGY
NvKrm10d3whaIAtNfw7wvG/q5JQT5K1MYHiVR/U66KKXxDNg5IvH13BIVi0m6Ho4
2DYflAYopD1lIY1Jy4WTpqgdx09b41GSNic76drGVh6v9R3YC8aolvEgCJszN6Ct
fmBvRB2SBos99LYmdyaZBeEgHRUJX22BCg/TUTLKg/9qWpS2eQY32zmwtv8BlibU
tENRZbecJAxwDtIlzabtbptsh/bTEc8n+HbGlHcTcgWdH23IyIYN+Gzogo9A9tdR
1nm6WDJclXiApepEITBDmuC/SD/85Ig5Uh2IL4xM3C6RT/kTn7BHmAmH6NKHh7YJ
IqJ+yRuOvh/15uPEA2gPtysSpjiwggJwdTfVweGup/u7LzH983tiquhHEG3WqXOb
AxgYZwyZm3C/dNgF/szgIZn8PofLcArefX83JUtVTEMt5PKOsH858bgMquhlfPYW
223AsT7saS6swyKuFndpm4YxwLdW1aKYIV3h8KHrdbly1sgE11ZZr9FWwZZGXtv7
oV4yGnBOv8R+C7RK2G0mMTOtCjIwgLnnbEAJtrUVeKsi1d5llFgaq9dNQekKaDFY
Erljz07anmzEe6EbmJhtqvV6BaNHK8DMz61l8zs8gnv0gpjTMHzcFf8mERozkRax
XKSxSbdqOSX3RLF3dT1eHuStUoXvi7pODDP6UlowPK6DEjKGYVVfFIdOChdChJmq
MCuysioq1CbJ+fYnz4MQv76sgu33Q3UugaNCFkyzjnGU4ualcnFf6qYjKsk6QVFt
1ZVxtYqO/kWnpAyv3wAZEWoqqUVmZ3MmFSHQpJ1oVZqL6wbCDRC/w4Hrf/IKbonG
Sc9B7YV/Pwi+lhnfcKdQ/Nzzb8sbm/Dz4+V9FTEju94vzeBof+fu8qrCiawe4hMc
/UMPBJg4x6PdIfmTH4Hg29YShIYBlQly9RUWaGdN8CpB/nZwJQ6aLnKJBU9IErUO
CEgkoqdnPWEOb2G606qdwAxtjXWLNypL7JWuKIhFHbnbySzhWeYvaei5zpiTLr68
QYD0AC7wqlqRp/udy3llMyW3fwvJYyayr39mJKwCnvaGb75x9czooxaoiWIzyXI0
aXsSCXWg8jXZF3UwOi4svFZ2gP1lSb731M4eGLAYpkTK50DWlR8bs4DH1/8c+5wZ
NRaJfg5sqmhwTL/3XMRUtzeAfTmsUmuP+ehk571EKeLp+/w7oRulEk4s8JvE8PSM
R1HQBuH4YjOy296Yr18MNgR+pKA/qNcXGPgydCq1fQUozpHFVrcJ99XC2q7pPcRo
IhMcCSXvXBp4YVNPuB8YypSm5NQqxZ6Qbl8QfHpZl74eVefrNvXg/4Rnt3SXfcR0
b1gtJeIfH/8Zp5vtwDeXEfdFMSyESVSzPpIfACcsseGWA5gGM3AEb76iTcyhQqOI
dqGWcb+/PkfqeZGdQs4oIPPVyJ/CnynqFsdtNEc2fLDtr79KkubV4ieAC8KQJ9/n
CYOucqX/Y6+hyF6qwY6n11vPLAUn8aqPsQLGNPgv5PJfJp9R6pG8symtr3HZP5Oq
K+OSfxLDRAv5EWWVSixOXXhYm8DqsPd1HfL5LbYgq1mUhsk1wlXh/2z0p9BRNXxH
Iwl4gsQ/9VVmwjDRy8nlELGxuGALjrJQykOIPVCICAqRWNfxN5HWNNJDV0KnSvZC
dd5t6hCDZkjhNEHdTXmRtXv1/XAbPS7/wkS1RFsCFPr/u9sQXYI6sW37Y7dlBfRT
/knTbdwMBa6RMd02FfUEOWcxzapZuZ+2rgXG/BFaYMNWoZzsd8IjsuVuZ/3GYN3k
UTxiZAQpDsZeYUnyhsh7N/NQeu7m4bv2A3C6x/yTr6xuXQcGAFO5QTpalicILMzh
zomHAMdvp5EnBVioN3fRFQZZ/Ytr2a2WWP/aEHnJcwjf8RokOjncppjTt6FQOowr
09lJTAd0k0t9H4KhRxKdixeLBF0Hxj/SfztGLmsz3R3DaFriSPHjWKVNrM5SMuoS
vthvjCqL1+JO+d2NxCUSGx9TCHR1QpD9gGirpnNfrnjawIidX457ZeJqk1Ti9cNQ
Av+2BOpIqznTRjg139V6aF5SnxMfxxvFHOyZakMPFW/zFUG5kaf+h14Z4eIuNntF
SnAcrIa0ie8RztmbQ2z18UrisMIoLbDsF3YWnXtiTbpjH/ZrpY32SbbO6AvRBN9z
CBwAUEkpDPw0DXedqfLQTTAIaSVzw98mBZaWLUc28OqnnJSIqaFxvmgObCpLSrI2
LfbWwVDJpPffgPiWzU3wHSLbPZX0AessG5J1VqrZFYEWv5E8/4KJ78RJwopIO1Tw
V4NrWK+F4Qk9nArdhPZg0l0TfQ9WCZeoSlCDoXioEhpWr6dcpcRCYT0/AUw50mB3
L4LTw8qNitGewNFziyp+ErXyDXPsR5KeNd3OkuT6Ht5sR7CWm9epnCKpOScpcgzu
xCDuTppoDF36bWqSaUZtGHTSXa4qz71iIxZPpR3OB1himvzxL8vq5fqHVd8m4K1l
0CuKmGTNSucVEvubbVtgX6mc79DVY1NvBOrf+MgUqXMIMdjn49TPvgU41FMIN/Cf
dUXwBrpi8AtUKKE6SzP0KOapQ+NmdcBwLhQdTjfWSUhAaQP6Gz0FyDeA7UYIOtJz
T2bpw1xQBfUQByehL3O3Y5/qPaF/MTGrbowxG1LLJneY1rpXwf7Yg/F92jRjLBTh
pXpBqFgQdw++iwam5eGS2saVqSl9jDOwkYhYDRQthrE2mdJctO0RFp4ZdMdQE31H
LOteOKLCQf+xweGVLggz3IJoQh501Y3VmIaWEEMG31eIgn0H7VRQGqAiS4Eq8TEC
05e/3hU3zI0IiSH+9PMVBF7m31oglLZ8VcnKYU7XniHmL3GznMjJa1Z1CcLs+Naj
gkYIBf1H64G0CLa2ceEoMa4wpXb4wQewxc1Gbuk2xowK52xLH5/1+KjBCIXHqTym
ZrbIn8SQ8wiyRA9UQN5WW8Lu+JT0xEv+2Lna03kUtEiVNDDA8op33P0M1QdhLrnU
0gKZZDyYcea//V73T9ZvVapHWW4KOfJwcpcaJVvglykKGnFpO19PwQtwrs6rw+2U
C842Lskmqo18y/7b8xXImFe65rWL5rd7ZqNTtGhqlL/S37RFd+UfLLUfi7kT/RXz
BM9qxszQlXEkYVHY3Q2W1G8nNRl4QaNP0eofJ90DDAyk5ruAT9Rx9MXrrn/Khq4R
+WGxqEP4mk4Qj+NOl9sNGNxGRoJ7zA/LdrvbT+kwUoAKd7a/PEnE30qZJxN7jXN2
wYRuEYALTawLSqliVfHrxL2jgIGl+a+scqYYfMCnC7km0sKTjH/+Xu0G1bjDQh+i
b+V/W1yKkUSVfqr+qTp2flNXwHyfabcXxoS1rsaKpXJ7v75YzvRyWPv8BJE2YKVU
uHVx9lD7neypwdLfwYVQOxIoub8pn5d5K0SSC4O9VcY+zt/be1uCSsN531hAn15G
OnY4k93jjtFTHAsGlMRyw0FikVaKdb9Azs+Ig5tXPpLDo+jDQ8Qw2Jdr4zEQSarz
F7zJZxRRyzFJao0o5RkiNAu6Kp+HYZYNxy445sMiM6ZVwfRiIC4+Ul4cOhCkHz4q
fQ+qC7EL73bybRKFVVOInsqiyssT5/WQaX4u/L/vnRh4Z2MlhjhOscroAdZKkdOz
BresCQ1Su1oiNx6XQ7TyXLjGN+8/2E2KS9zDnSBBcCgpLMedcZre2A4mY76g9NiI
5fU8ENpLM5tgvjQ0u1kTqYVVJMFBzeF3yTwlEeZBy6DR2BMkZyF4UXI6zdy47ecw
iZ6b4a2dV7AhC7DQShc2tjFSKYPHnbIKE4x86mA0lgGzUzL38sDvXmoWU7HOCUlD
R5uNJ2nCEFZ9dM6VY1iKh6v9Jm9veIhkrsW8BiLF1N79kmqVR0kb3R/l/X53gjP5
Ve8wyeUJLitBPbN8RNXjyE4iDN76Nej/OXEbjlgdVsHYAFWXxRz+P0wuTFlYRFqM
RJof/BpSDYxY4ouot3K79nreM1dh1M4uSZjxR22zg34257U8akLJfidpaX5uJhK0
gh+ruJDoVkUlYopD1hY+a2kYb5oBZz8AUbGvSppgES6HdMjOm6RJwQj24Ja2vvri
Wj95iagOzW/fofBSamvkiBiQrmx9dsAze5Uu3m+a+hhvwnyoZ6qCKZIBmUqK1CSX
AMNtRSOMzmOWjMi1R86Qp3To1ZOrYxYkaO7eQdl9qzKe2PIq7btnzfWbsyGx7sY3
pQhFeckvJGCDGSgyYlsuMo+AY4r6dOtHlxLgg2MNZKatpYoCBxepgE5FbPpQQPH9
LGqlgW8CoY6lyHpUlji2zbyr7in6mmk8pJEMsqHtbnYg7QsY3KKpOlPmcQ27pbpx
EgA+8+hTUXwwv7wphEBmswDvOC2y4BKEURHhzpDiflp3u7WgCT6kf4TzZgizBg2X
Q+eBuHasLi1vdstPCGjAM5/XECVAkyN9o0YlVLfftgR+3eeljEl6D83+RzUgx0vh
i780B9yzE8CBG529r0HX7nPY+7M8oWM+PAWkIuLyS07xNrAMMgfMBF0O+rzKaKqr
nCl+oFMQuPSPRKeYw2l35u5Ao8e1qKGIYzVxAM6w4uyv8zTKYXdn6yGHIO5TRVM3
nawLVuGu8qGmp9p2XWZlhQzEp6N6HmLHoRKlfgZjEg4CzciFP1CPuve6pJWxQ+l4
9t83YB8IJQgsB/FeuIW/p6Jbj1Tm66qf1olvykk7BwPu26Y3UuE/hHHhmpWXIFBE
leGnf0xDhyDqinD6FF7leztUbk/t3vD6Mdacrx1eiKtuKDf7i/I6l9H7GHhCipd1
+85IJWenBfqAZlOeT/HXJHxrH8Ckr6U1XvG8+uHnGnt4wRoaqKIiurrVPtM5KJ+b
8DGjk+0GAi7C8qMuespqovIaL94ZzTx/cm/Qq3KJjZ1bXufBnKeGxm1kXIodlvjV
fjEN1Wybjc3RaiRHmBmQpRz7V/gqHrF+BiIM7XPXyYUW23nzyWfqhNVr1IKztnbz
g5vrmZq+xnYpGW9U/xFApfR2vv/8BSuvY/Omhf44Iskn5qex8L4ybFJExTM53fIH
+3E4yl9v8eFfPxBjeqKGJWyOfNiL7J0OOjNXeIxlriA4zXWlyRiCQgIyF+ur8lfA
JVvNbqKSU3RYI6D71V9X6NABjsFYbx2uTyWMyFA2Nl7UICD2a8PQOWk8rasjEWEy
0yCjQ6DthSQS1mY5pNkZOEJuEAobZ0W5IyTLdoXsrIfm7T7RX8MlQESgaGMWLC0J
AzKQ5UUpQoPk/iinKSGDyHnEz2P8W0ouWg43LY9yGIcL93HcfFkdxLD4duL6rzWm
0fU4w03roJZ45aBkWXO/3DWcK5Y3oimQ+fV2/i3q83u8LQQeea9HF8tuzvzrlmqK
ZkV1Iu5D/NgNi2XLc2ili7J0WH5pS/Qjgy7ocgv+gFHOiGYaFsvWRgvOV91F6gM3
Sz73ch2XXJu9rhu9glsRxysS3Y3Gt96Fkbbafg/OuLn4Jyhq0tVsVUzn+xnzaVz4
XlVcZOd3zaKNohfBstOiVTUjvojwkDvFLxxGwJ6SXl9FpFxiinMnkUYzSM18It67
bUv+0iUW3RSuzUOKEe2VfVNq+FGALgk8zJdPyZcYhzOg8x2hUowMtf+RvPMB78E/
sRWtQlM0EsENUTIrvLJ0WwuP53J7uYFq8goS31IrX9P5nIg8a1sPqXq5NaBeV41P
Dx4iOVOpuN48CWItukXgAUngaImiR1XhQUgN2MNvwYUMCRbXWoSL6xfXGkPYNHnX
vkJYz3++V0l7kgRYXTMFt3sC8XFkj7nvkiou/vQ8x8hznhkFOZjEdXmwp1sjRZ5J
J5MDKkoaeh5LItu0keru9SSn5r4eRqTAb6y36Sh/chTAggw2ccphyxZkSfiOhNXS
tSCd6rzd7JRdMlTy+dCIoZKeURbNK2vfHGv9SVy6/NAhWx7Yb/bgVAoaayOKOryk
g3NL7FsQ5vik7cWRpKMU/cvV7Z/8OanNmMbGTsAXYEcfxkr7EfAF0zLbKo+zAwT3
NBfpTh70c3zkENm5qrprH0oL8tlvi6ocCcMhGba/Oi9OLLvfgUFy3Gvqml/gdXcR
EgALcGt8jLau4LfSQ6RaFBiyNHSkfU+IxPToaWwjiXQkfx0DGt1EFBVCCTrRSJDF
S7UqxFoH78cazcCa+Y+7M69ZJQRh8IVazoEbmjmh8WNrp+AyySwhk9empVK2U5AV
vnpzww+UzweT7TduNEUqNQqBVEggqujs8eED1rnnutqA0EF2a5UUfYhz3jtkdVCi
tMnml/KsGxwnDE/NcKaqBOsw7hj2Oe3jgBBsCcOubcOElUR/7NYqIgR3YrOGhfIQ
c9TLmcdbgNfJmJaxGewUh1HkhJzSSGVgE4dhUHURvlEv+flOjVXYLDaq+97nufeO
242wVXHp6weKyOzzqdg/KwD/Xc2LSnaEzWCv8lZ8DRKTUePkSGG0uix9dvqVe5N1
x9FzBsA5F+TUvpk+jwM5KVGPDdYxB0njqQuGQYHnH55uYadBFxUigQxQKjXiYywd
NB5ysQtYqx98l/vQoP6Y/7FuZJNwx4FJLN+YLzdbCLTCEvg0xpvPmE4SJay+uiQZ
tgYMYrC0DGGYDzwW+YL9MOOhpZDdUDjPb1L3XWS0H8Aqsvrd/Y7G5DWnIxi3aTLC
4SmpPVttx9WSSE7HE8OEW6VbibrEBQZQnXlYSIkEODoRZ7iquyk5rVYlF1+tRYYj
rZwGzbmnMhAiDuBvRsrqUhJJ/hcjhZbrgbwL0f+qOxb41m+vrEwICU3jFRmyzuz0
ZltVK05X56tYNYn6jo8hEyrjwto9a97S00ylrL7+aTy7vocVVnxtiFd39MrRavIg
VWYvOsH9jcJuqUHlBdUboQdC8i8nvPjloZ+2/sSQfNSpSC0mh9s4nQLcX/V31T4V
YngqS7vCEiWtF7f0P887PDEFh+/CQwY7qUictvhPMquoocKCjXCjQyQmuXyWbKcQ
CZYFTCmC/d9bkPe+7Ls6QGnOY7oIicr7mTVp/RFFohYBbgn1ZxaAvoLe8pcK9SPy
T0XOFXw9/b2otivh6NdQChHa7/DhESXQgHOTMYbirG2rIqarf3onFw1KRCitlidV
WxRRWF3u4Fa088ItCL7rtfE6TzB16O23wKmh495uLMrDYyimYsu4EBTUbj3W3IS9
riJtAc34Z0v2Q5QngT202snT5yTpQ0ajpw8zJurTnIMOV14FBm/LinPO0FL1SvSN
xH7AjG62eBtclx27Z3qpKGYx+D3UjFwiYZVFJT74WbZhdTAnmybnN6gp9owzKYVG
7JSOtQNis5iDDia7FICC4de+EQrF6ZCBJyPfC2CpjXYFDF/SU0TeMelT/9TdQs4m
MaeCbed8ZrrSB96LMtd70BGRuQ5pKZaCROFHq/rrNuluUn30943jTVBX+13wumNM
wI1jJyQj7Q9qk+nSvpjsphztQj2iwFO8DT2c9b95UGf3zd9IP4oGhc2TGhkSN/z2
CdFdaIBD940k+4pQTTnwEGufpvug5Kj052yESLJcIdsdSu7+t9kMKtcLmEX8iIjh
K7hHCcI0mJ28ZCZmuGRFkEaX+TGjx/uUdiHzAXDrsVwIl/5kWYaIy9UTDTjgH8k5
X8jVkYZ1RZnM/bWeN56InfD6565Xli6Kc2epzmZuc5EMfalZz0+oanMlTOsqJfwQ
mzM7pzsvH0dI36fFOA4T4uY3ekOpBo3R4AmVfckpm6cM+qkP+D3bS+uhRLMrvW84
cOBn97BtgLkXCRL/8BNdt58Mhgous1YW38iQU55r/kDKMW6GpljMRALtI2ofPOBu
t5BWgWSpY/fl49EOapqWtZycdogeYKzYRai80qEJAHHC6BdDsAzwrud22xD74Yf1
HTMFCzeZ5K7mZ2kg9yb6If7LhoiMmFlw1iiCdmOTOfewu4q//2mrgMYYpW8+iwzb
AYpMIUyx1PsBEOMXFE4X7YDVSQvJ2A/WImYQwy7oSshFdaYRhw5rscJwwgFYGf78
uDXj3M38GqHiCD3nm+ppiIHJ6L4pJnnmfE8WeLvurp+2wNVGADpz3wh0pNboUWLu
0bZwUqwU/I88Gwb41Nvk0nLTnycM/DKvZ/1urYTytjadqb7XM4CwIv5L8RyB+78G
pwLyMWAW1VIRbXBtdrXIeafjvy7QpfvlhJsVA+8F3MzLFtvRK00v8akTCGEA+MwW
DgzzSGb8L3ByAanvHr0PdKgSJEuo7BsS9yPOs0vX8BhKk48Us2Oa8HK63ZqeiqRc
m8Nz/OWGcpYbvM06JdwYMBZgGUu9YBOEU85jstVUJUnb8u380qHPvUo8nC7hNCru
GFaoHK+LAoViBNd1AzhrJUYUIYV72VxmEQzk9MXau46wc37EgFywhg2ALCJIQZ6E
VSuFDQCbQgV9BznxyCo095zjz9SYOqD0/b6MXlaYdkHTErQe3H7UlLfMRR/kper7
q4nl/wgW/20nVa+CG0gylWTugkAHYaWO5aEgSaZ8mz4dqpEYFELty7y+YmJwH9S8
QTy384FHYaoCSUxhrN2TK4PR0IpX4nlBdvoSeSwXIvBjTXdxmIpKH8ZTA05c79ST
nCckds819P42Fr65FyiiG45i6WHC0iRLHb5xWrFIxGCFOdTHhX47EmKwBgFO5g/G
7D+gTdXsZ6kwzC/QnEeVr6Xu3CnSJTR/UlgQTWHtXvxL6hZGxPkzxelDTTmCM8kS
EdV7f+tgUbVXKYr4TFQY4QpLHXzPiYznvVpUak7pVB3IDDUrJuGc7ucagpYiL1pn
fgk/e7I7fZ6dbuQ7qNSDmGk4izq0/rb0xcKKSygEtVbiUNv2otB6wrKLf1RTJMG9
9YbFwDKvaD1YB+7cvv6kGztDCB8eK5PD0PF8Uf1Uhi8rxV7UONARlZHjoocT7Z3D
b59jmRssB6UgnfF7anGKRQDL+W+cdLMbDgsxKMWsmrl4K6uNqYNJN4K4QGIB1OoG
44LiuGZbkiBxfdN3eVSCTBjcnnYUckfCUQYFS4WaJ0eNWqI3asDpCgBvbooBiyNy
aTmALyTq/gd/o5eXBEiTjvCeCwrP34Rm2wvQpqk8qlv0b/3ON+r9/NKJn9tLJN37
vJ0vwh4SU47MwDfWsxG7BN8G9hUyMiP3qIopnO82sqtB7sNw1txvRFXTYAAdtE2Y
oZ7+lTxL8WNzXHMmCdfkZN5s2qyrPG9VuH1fgJQ8vaVYKUvRTwuHmCoZ9eSe9wGa
X0bX+iw8DSN7xwT4EQKncC/zIzrG7lATF14vuKitXr8Lp9cZy4BacTHXV/HnxGzS
vDLhmzjDPeBEjIQxETJxcE5IErv3mguWZ6v27NLL3EfgaW9T5XXcC/PJBDKZyKbK
K3uv4T8QEwB8AzIzXkyzgpwzQZ0fOziEL/x7P50cKENC61R8YDAs//NNI77RMBKP
UL/g2XUVtlrde3u7vtJRlDlYO3/UThFiQ+As2sj19vgUd18LinikU+gkcIqfiSdG
q+d77/p7Svj8qmpvrLX8ICJ7QwqnHhRXBbIwn2XoPk9JzBlSC+Gmi04+W7r4IZD+
HDSEk69BbHUtpgyfOoJcxWG3AsDTvf560UXD6f5PrUiNQmw7tLI1+zY8BFqN0RYt
sGWpyxoelKHod44VHbY2jmHvhLx1Z5/CzsDmhBWggez0XT3NRhgYZ3JhUOJgTgP4
cPDDF37WCLkcYSiP5eS32qrEhAxHncBdKu5vTJ9bCWmMv9Dg26S3VK2/abgWiszl
qgE7R/S/Ck2z0AUdX2YGOWL1JFHTToB0BFl4u9hyxA8/S3SO1oU37XJXMK8nHTfD
xgaZO8ryeI2TsUhR/QMdXHuTGaHkbUI5pX6WVQKdjOQ1PQ82Pfw2iK+ZV9GOypC+
cMppkO4OQd2prF7c4k7ihif8+GMSpqubTbuBdlg+LxwB414HOHxtNYaPD2Qk1Bl7
KomM/anS4yxuergGgCoMUF5qm2fNpI4wqYRWKWn18G+MBkXsFpF51dxqNxEbKYxu
MlmkGx/AGvCPShBK+BMVGxFwdoHBBced65FocPsJO/P5KmMMxYicH5wq13vFjDvH
TGFxQRsSBUT57ni4s+7gfjtBYg7XNNxnF4vwiJLUt2TrB88Nsth5qlvuDs2nC8kD
6oS7WNCHQvj9H2tqx+DK0zl9gINJLqXDY4gxBS+whNbKKvPVUyM9AzLQv8BB+wuS
QLXqLMJdVqYzshDqn/r7f9FX1MLorUu2DM13+BPZqR1ZPZ3uH6VngDTuiRI0S/A4
mVgM8BXCdad16+uimb754nWDk5zHez+09PguksiCz6Ee+BAn18JScD1260nsdrdR
CyAsHpGH7PAanL29vFvFzsMtB/YdW+M3b92Y8WY189BEjJLObAuUqEwIUJLUU3Bc
LJpeQp2dDLwdetxpxyqHKdoYVGGrArTsk4JFZKJ3L/hRaPWadQhlvWS6dYxoQ8Kh
3Si1HPxpQPZM0h+Irm/7YMX6eXQy2vnxnQtzJNBitJBnQnzaR7pajXUsBXVJPi6W
lvBMGJgoQmwiib2UWcz65VX9SuxInfXqqFtOAV9LBn3ndrwxv+X+CADR9m+ec3il
eHnjyTR6jXaA8Yx2w5Txa+r8qR7szLmEbxboVfk6Kf8AA27WRFmZwTH3qZkKVUqR
cpv99b6dqpQ2VaDLGEaxJbRl89aXHtmVD1SIb/iHOAViKxFZw4Two8YKZZ+SX08Q
SgsrvrnsLC9AuyPxliLPRuEvsZJeS1BbzUFaxmO9aI4BkGZQQG5fqmcCfSzz16Ow
GRv1QTxrsIp5xrzGXdtewelH9f7nqN+Mc189Fny31pInWd8llrmBpR3YbPGYTG42
qnS+EJRZ3egmvHJOvQSS1Nhg/XLYLPZdJBODAYuxFuhmcUccJRdi+zS8cEzfn0w7
ZmD8n1bYay0XD86UZ6992Hl2/EWyo9DtDwihwUm8qksO+b/nJW6XeXUtenZoDDTg
XrkDz9KRLZROYFnwtBK5iHWsj6RiRBE0ioPyzXLibmgO+ek7ShwdACqhjslzZk0o
B1eUSwUluB7a6GO+apYhyZ/XghbOaqtNKk8UYik3ksiKMPd3omy6vPr9If0LEruj
v4EKG9ld4uCKqJFshJI/BfKs4r1JIKYgdzKyTeNra8w3sKeU+/2NzHcBWbAfYsw8
QbemwFM/swXEaHJ+CfKGImGP/qT/qHQpme5IMD8Frm+uJvRGexuHk9n7aN3r5X9E
jtfYVmQSI583bpXixJBK1wJj7WdiSkG7mNBp1yeQmzKxt09FO2nL/oPGqBH1ol1G
NFbtKEHxY8G53mJX8h4ydGCeODKifSAuJYWaCMzzrdGWcWbIg3RgGvHSS5vzfR4V
ZIXfLngRFJaTyAYpcUhWbdXz8A+iamIowHuCvSnBlCMNcJv44dgKeNvepVr4IKkR
/dYMrvbj4dkvXlFcMOPfnFED5lzVWKiPl0f3MA3b37CojR4dPcN3MzXnP6CMFN+O
YzHLM6YpUjn+SlKSqOtlncMnbICyn+FN1wZ9mog9mypI7KWPkqt7bLO1JW4wMlXi
/ikTltWVXlPV1E8BQpCH3KeI7bB2AKvT/FkC6BDEK486xo0cmDRxEMne1hvmUh+Z
5q34pppYJACSgBLvv3kBe2NeP2aLDGAcZS8JjW7jLYnG5NqxaJvZ47ideCKRLnk+
9ZV6uPoU/eUCo+H1SAdXuM+1LW1GpXEXqNp2kSE1aa2qKts8CXEHByqXOsum2hxO
jQPciuJpClPkLuYTG4dUhp7Q4L5O1b61r7huTthZkbA4KRu53ErnQS8V8CvKt0q3
43o9aYvHfz+KWyF+DZehxXN8JQ3rdFY3tNjBtg/pkl4Aqq3slvlwQezJMo3VeTwp
bvWSc86Al8aR3jbLqqv4x7tUIIXaTfLm8VXlazh4lrMumOsxreV7FOOOF90Wp7OA
nZCEDx8ozCsZonc2DraAzvjtExA+IWD9JfeFtPJghDoR+OTEHIEyCRC4sMibz73o
YtJWaG2jc8NwoFKXxnWKjr5+DZ4Y1DnTUcEpUMwQw/fWzOo/pmMDLEzVf1fT62e4
+pnjmKzPddbFotcStHnTCXScPPnM758FydqDIYUk3N2LgG24ONjWbDbgew9/Kqog
lBKr7ZInilEZPERB9z/TZKt6UZa2hmD8Jr+MXla/OW4zG8w2kUM3GNHWxr1tRP7R
3E0jBnMbk3sDGwNy9GrBE51RmekE7hrUhTz+2gQ0FXxPfH//g36F58JxzfPjqot0
g5iHPMOcIOXFdVqj805GZVwuhaLy6JJmQXOTxtVsQhsvCkqj0iKKeFHWNYZcaxs5
fsrwE650201Qb6Z+Hh4Qf/eOb1WIJigWPa9PLdpU1dbnR84M1ymCopc0eV0ozAHw
DJ98GRG7pGwrW9cJX3R55KDdLm32C2za3bqQQV3r+XD7xvIcHoByADDjad0hJ01w
sWPSAC5f5sQLLzY8vzVPOJk29/jOKO4E+wZXx1fKYz25Ig8t6ZAEaGuR+CQlXGqM
dtYZkoBTF90ux+6bnsFNfrAHpWjY1MiK6/aYpZ6+4DmbpnKxYyl3jbHr7kAmzmQV
B1vVssVPgYYPfJF1FEDUsk1u5w+anmPFF+A8SVvmyPb2Ckh/N7ZV312y6AAhjzpc
uy+MeAreNeSVyHnfWY9jm0YQTrag+y2w9OimsTTdDvd88t+rLFIk+iJDg2oF/7Q0
Eu8Fm5y5BWV8xY/Lx1A4a237BpdK/0iy6+RdDbHY4M2fvnOH59cDqU6TlKwrbxb1
f3BmRZ4ADD/o7VD5odYqJXodDxgJHb7aTrpYgxgeOYZZW168I4IrB8r4theA62rJ
9BfjuGRuo7JfPxSaOyNWnhhm8t2mGfi++rdw8aJyDs/3WYO7pDwcf5roNythEHcH
SBGF58gQCAoPh78gPHH1P1mCJ+iMFcrW2dyM9UFsBfbCoP28TjuLa1txE51cnM0z
NMCbZNR0HOPkE0rAeNOTAX/qLu98FJRC0vIBRoW/Bh90Zj329CFlF9i1rRqlrgEF
7BK6KEKw6cT+VHHLxGKdXNCwLfubO4YfYVnZwFBuhA+Y8aJqT5yGAiMTfyv8PKrX
zXVkFxfkCC/F+T0zE+tG3RTZls+P0pDDn/t5/Q5AnJLglhHZRI/D08xSyzI0LeQp
kEr2KbyVE8VjHmOIKkGj226Fkw/ljCkb6OFhdqe21FPs1383L8p8Wp5aLSiv+Gq7
9AvW7Y1ZXAIaEOQRgg/sVMqYVXsIDeRQfT8dbFiSZhBRXDN7pUVHxGm9B9Qfveii
BWXxyOrQyHVzTX9QUlAsdRc2sxzBWHQe255ccrCeCVC/3ZZDXpjHHSpUGWT2Bcvh
3gTeP5PhTkruQlrdz7Kb04yM39ySf6j0KEmNxzvGfOs47xvXlYNUiIbXsdiQq+pm
VURb/PXZk2YNulPxPS5J0n2TX1QcjXbE5q/4LfCXEnn4A+vCUD/LalxvlqfeaPG2
wgdq5cmClgQgqbMODUqD3Guz/6KcgEGSyLTkZI8/FlhdsAHHT7n8Tz6+z6kWGefd
BSGRPAfS83K2IOhBV0ELykYNw5MIRUleMQleC8n9KkLsCaz2qipqkAa3o9Zmza8g
hoafNSS416/0jM8uyfUfyLMtS4wu9KTtH87XQnSvi2+on+979pnOcAkqwtLk1ImO
1uTHFcR9J8za7+b31GXRNFaLQP1734LVenzq6Z+MtnQ=
//pragma protect end_data_block
//pragma protect digest_block
QbiKn8lG9GaRUK7PnkbsjvSZ8sc=
//pragma protect end_digest_block
//pragma protect end_protected
