// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
CsMfPGCsWHcTfeNppLhIXcB6OkewoZXB3fRAXPPSnUQ3Q/6MVoh17WguDsP74HfqXgixSvJ5oSc0
8Nukc85eL/1LGIdO5sSYdgGB85Wr7cyY/H6lhldEBg0lUl/spEyAPKCldrLjNuAHOO4ju8//PWwe
iBS2VerA9eoklAvksD8CXzcdQF/GI+DnlOmxZNC85yLBIsxyEVVh+hjCcYeQMKnLNQrNT10Bu7bf
4KeRWEHMFkowsMBHuKtcygCyzvQW79O/KPwoJtxE+xPO4O/I+WkxGDg/f4G4Cwnah6O8oKh5RC/X
O8lt3jXvuCasd7sxkXp8i9+1hbXVpUDtagTrWg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 8464)
sqAABYmrxDZfySMaAu/4Yt9i2uk1ZALIwzIdcQbRG3BBY8GMTa3hlYLZUqSJEDr9ihSjMA6r1JWs
Z+hVQln/qvYDLDi7Ksfbg7CAQLULqs3BXnTnxW/OdCjV8Tdev/L6PC7dkHH9ASa3GaN3CMp/pCY4
XYsQm41rjszcbscPH6oHLedr1ru3OQ7S8min35iUyAJr7m3z98mfEV8/79NzuUTLUplEsdA/9u05
u1PIZbWNozxgOzftFhBErFFhEjZ9+TL6/WqRJsiq1CJqK/4sywbhJ0ri60iugEV2Is5cWH1RcOzn
S+m2NY5uwevWpu9Ce9cm4xtZPfh+GIbufGVK+fSme2D65bUCSAKZQIMo6tDh4TfDu2h212SOoLLj
hXJfKh8wnufi08dyezY1vbZ+8WjxUIegzwTMm1Xlp6Ul41e59b/akhtWWpDnMqdU2Y5gaIWFhkcD
WVR45quxCR9o766fp+QCpgtfhrb53q18XeB0Rx57r5AT6+9lEW9yKQ8F/3KHE4wBW8hHjmL+Gn21
Avurri25iyVto0qZflgtLkzsgxnZvlEDPtt55HFOS4M/Xd0WSELV9JxmAONgZARqXab9YQ5uYGmT
C8iInfAYtsvBgvaiLnlwUR5+XKBtdJ+/IIs+oVK8vd4e4B+AUzsdLW5tYyqq3hQxSQPrl5KpTEpj
gN59SsovX9RgysDwcEjOJiiGq12tj68q4w2ZMb7GNTUt9NHz0QwrPyqYWuaQMYqcv3dKuTF7tiY/
Aj4i816eGnCci6Iap5XfKnNw96noPKwANAO7gTidOx79C31/HCu+f3ziclcnTMMvHWk9W+PiUeD0
dHuMWRk10HS42wta2fONTGTM4yR7D7rOU0rleFPw+WYfKejH1i76G/KNIwopu/NVmoH8D30bNmcq
g5kUaNo7aXi1cmjXoWXyu5RVDahAAGFUdQhY2d7EPtUnf0cHKX0Hv7Ni55XlOpFLfvD5GeOz9QG1
vBZeHmac5qklsBfFL9Rh87fn52bW0kPOugXZ8xvglP7yfCZ1UHiVyQ+U3mmnKllg1I7A27VX0LUi
Ory5FX6NpWSuGplrDEu/S0MUYnsDb8cxTeob79JteUp6fzF5yjYUAisaMXftmvuDU7ufUYphdYwH
EjUQ4+Jy487OKVQlYPB67WvsWEz3pDzayY3VmHeji3YoK/7TOrRvbopq9NBNAfKadIgghrw09iVc
SS+vk3qdwwXZCslxpxZnjdEySlLmlTn5FzhOmyrQ5Da5tHDbRsHneC8r36FjHpnCczD/7+j41ULI
G4fbwbgs23AO2j1L6XwaIkyLTcKNiULzME3HfdtAOedSuiwI1rBblwiF4T6844N7PihOZlaHcbti
6+MQNvKhDMHXdUHK5zYkO8zPEJJxnxqkd5R2mRPjNuDgo2d1jidP3BDVPr7qdSp2z3VztABEN9ug
y/y7TccqRPqMg+4R5ddsrPTo0aKM39mfhlRW+ZUZgfyuDnC4TVsoliVUCCsrP9OkpOfoJipE5Q5j
m2WoBeXQDQ/afe2ybyujzbfmDXEk68rK8Hci8qaofjQaH/jcmQXAL1pskTidoixn6TaDMBdXhPzE
4kaaxPB3X56k0euy7s0M/zej0Aqi/bWBJncX6tCqSs2Vot/SgbFZPSEF5nYij3g9DcbXOgUBiNdH
U0zF7RUtxlk8yc4qIxzvFIxloy2yYtkDtHLop3HdFlAgvrqFIaGPGBxWun9pme8RN/RxeF9pPCt9
kYEan6ve7JZWiOcE0bdfYPWTiuaf6efM8fullRb188hdzNIpQUS6cFWPjVTqRj3XVqvEo1yHGNCf
Nagatt9mAWZQApfBZDX3OKIqgENCrebPeDNm8XFoJ11v/wnsw560tEI3oyQJf6c7B2yxwW2r2Sok
bOUqk6UdIqnm3XGi+uuPSIZG+0nNRi8mYVgTgDPNlxtu/m09pME+xEql3ovXh8fFTi8F0wcUhEJV
Y/zlkpkfRNsKpMB8VUSIU2UqewjV9euU4DGCvAvpELs3etCgx4ea+eJ1Yb69TbHu6hSl7P5+0cea
mEIj3E3NrjUGgEbjKSn+D/cs94HqPVSJoB+d1XrGOKHwfD2VZAnr2G1U413ncqkTMqJtOGXjx21U
uvxgFY/nEQkVVJPD/kO884ZDTvAl1PMoAanWXMrHXB5A8oalE25gqCleYQ6+gzY0DWJOh0JFGXiO
Dc316W4mn2XTiCgs/AhmX7PldArd3/Kj2fbSyPI/R35kMg23z7SYk9/jL4vIl9Ta/i5ZklCTtUt1
woANOer5V5lW9wG2CP+4hgmQRzHeOjoAtyStdpRGr18SopkTquAfgBYLwmJrycCNAK7kwcnrZWbh
/GmiEc11VRDbh5mq96Gjm0oRxL/BIhwCWP3psPkfFDV7xK4p/L2MeX7WPVlqUnprEu+v8dW8nkfO
uR7mTiHMAQ7RUVAGZLvMKZNNPIPhJG3zD6ZXv9+lIOB+VhszsWdnPbc9OzvkxKhz8Mo2xzjNcqHP
GrPkFnDb9MbA2SBbGVBEWsZIXa4fDu2RIBShHjRduThoIgW2avP5nUrsHIoSl4RXuoGvWMjGBMp4
RurJaHcQbauZm0hrJs3VwAjvMgxPXUOOXMbatU1WFPI890a5hWPsYQcztHxfyJFn6sw9UNhFWsf8
MrD3PL6fiBOTCyjuXj41GRs3xt5wzKk0CRZ3ELujMmnjEPbid0vUg/gM4/Ue2yC8MFKwyrUGXAre
nfFdOflyYIRuWIoHRv6WWX5RMKEI+vz8cZBpDAWDd0bUvVAMiAQqLRbLdSu8MkyaHFAJhPA21Ekb
qluWWdJ/mElh3cZE15U50H6+EDgexU0yb2kpd1BA2UcU46o++Glyv3vQhLWnINXIwgGLYeCvxPFq
2MgplNO7Cm1neByZPnioZ2TqKtcm5qQ1gp6YllYZQJGK/nX2OF0BBq+kuldJkfg2Hku7uYkCLnE7
5KoaQX6ai9ZoVA9phKtK5G8RlhbXG8hePLsI8O3fGBVQqhQkTOam/DbMG5s/Vm/CTCEVPpr6rQ5a
4ogBGuheQT29FJdO/j45qTknUCH70ShX8R0KRKqQIYwH2FQqo0pWi2znkWpv1qcYuPVwjLt4ebwa
vOHOVUeg22MTZNtMEE8CeRLSkAONRewohwK3yC8UZy+nbOEc68moFHfxSIvfZhlaMIpJxF23SZTx
WVCUeb6v0kDog7B1r4ylXaj84ZyR8L3YImsbH9VIs6jC6dxO5cFF2AEfWztrhd+/c/Oq0dGUggyP
1SuZ3xj5B3W0/ryYbR7DPG2H8L/O1HcMhdgXm56x7AIWu1DK4Sfa9M0TAhgKKorkiPytJ4usvW7/
XI1oYIFhZ/WDSFMoukHPAM1PLW2AlL35zz9wEx8uHW1oaRBo4lGfOQai1s+0wz9TmKGFKQSD42G0
h9S5uCTkQgERlZeib7FNNVDeII7o0lFfvIkRQICSwo0elN2+a0RZSVi8RAmvWmX1BmY8fE2N0Xp3
Fc/TXGSbHCTTHaxHLHP6Hpm6O7sQoDUC/DoC/Xne9hXLAdxQOxSItp9SC6OUcXcLoR3JUF1qI4gV
2RBqrlgKn5mXXJW+tKYPHxOavh+QhIr3RYZnq7ob335DUYSVYiaedmB22PY8MhxsbpQMz56KN2Ev
pQhs2sVJPInTqVs40icUDUbDhpGSZdcHp9PtJxV2OoOXDIAAcpWVCeeRxdWJRo6ZlNGFN4UyAIhP
6cT/dWhAHPLE3QsZ+lpx+iK9v4ZgvdM+1+gm5YuHXlpaC5Kn8c+SPayHHJKZgOYNFKmEj4un8V8Q
blWkuRWQr4hJd94WaW8fykU9yyOb6F7LQU8Ji0YrsE8GhF38EtR+NzHUHHq3OBMZhxyvPPX7fQF3
jl8Z375M8KDpIcAcR5eIWBl8kTFzF03fDfkSeIadN1/XA6J2YpeKheCS6G4xX2qJMx8fW4Ppm/g4
D/Wnk2rtvkge5V3bx9w6x8Ju6sqIptgF5Uw9V3a23pJg2o5PGHnMvG28JsMEEcdctJ16tc7vJw5D
VuJ4hHvaHxsiOU/1PZAd0ZuSxEm2aPHyfmeYiojghoFydDrw7h4Rre+oJySzFzd0tVfase66VN5J
2zN6lePZCbseMQTuad7JI8QRbb9hM8pFL2juq4pXawyDbSgqZ6r77udArVdSOfChAmlhhPSxxChr
z1RlwdsyhOWBhe+bDDU1Rk/MOWgc+CU1SzZLx+XFFUn3JchQ1Wl/7i+CIf1LPu7DxxUyo3MfplIh
TUmGSoijWufNikX6XXW4/LF+AQARgtSehbbZjAsNIaHysWJFoGN+PYKdUsllXmJsIu4nOh2IycuX
LcfZQry2Csw+uKgQgC5ks7a7H5AIKlYHX5q9jTwWZnhmWNLJEXLXdmo2ScRI45WgifKrw+CTRHUb
tlYZYfgBRJr63Jl7UtgmqlL4b0jCarPqnoRuOx3o4fgPhte+R6TLWDaMfmvhT31o2hVLLfqmu9Lw
m66xBwMnoJMF5O8VdQjOleQuDDKeF1s87EhUNk01jiArtMIn+e3C1IwEfmyBPYnxq3RXebZVzbn0
6E2K7bnFfrnMB3S8BSTTDH3n4MygVq0YFp14XW+hzWxnSuiO09rdqBR4cHOmxus9RGgh84cNHf4f
U/amGXK2u1bplXFtwJc0hIgM6O7iTeUvD999hGlPtgrahCzRLgv91QBiYAyI+4FkOjx1aD0vtBCE
0cbRm+jrcO8kP/2ZyuKLtDCtJ3SYKZvASS9nCkxhMs0UH7RHzujlGFl9yh7Nvo7dJ8tlkNyFPn5r
zHDHELoVlGBiUbjUcJtPKPu91cAUbUwqnadIdWsr66Ybqogul7hAamU/nhK8tUp7bJeYBrTjr43x
vho6gtG44g5cFe+4pN0wluTuSYIC0c99JuGhQEzCNxbW8i7B8lNLGtScj6S+H1VhBjLqUCKHx3wC
YPRrbrt5l+B2fZQJfs5mY0CFNldkGlJQjIJxm9FFfY8UMoqF6nv3Q7LOCVzWehr4OYo2oZVDLaST
whu+EteT9Q9jHJPoQRXXopaTf433oh5kTWl+b66rqHxKofQyHbwE1MelL06XG1GwuGmYdcpN59fJ
mQalw+BY5UoMD/fxzUF+GrB/y/Lh+2qpJuaRd34oFU7YD0ZRmb3/061rQIjffaWWzFcLpNda4XBu
sCDBh8v+xydV9jqazB38a8p0kL/peyqLfKE3QouWM6q4dxklT1cIqHaCINQ+IluD3fJQ3wGDPqQa
6fyFm7cRqdXc2jItQHqzoxTilB8FSSgN5xH8uikm8fvfrAPQzukvxyzTH4K9WIUY0aNZEe5a5lql
niT4ZAVm3B8trSoD/W+jccJgsAMOPlV058oT9AzYJaYV4wOlDLWBDFdoA8Y2FvpRG/zqn+snDQc2
dCmhMvjo/ODGtLEerONvnYgfBgkn5D+jFfhyf47S10H/cI38/Xe0y7BFIHODpIRXFlb/hq3r7v5j
65C//gsPP8415aHBmvG1p2fxFpBqDfC4cP8IiJ+zGEQucFFcEyI/UuEB3gQu458XIctp6BYBBw34
jdlfDJ9Bsx/ZgOuM/dIpOKfvheckXinj5WE3F8wxWpFe3ZSZoKsCLkNB7GhQHivh27IOMFwGU0Z8
ZluvvpXcd3phTsfQNW3GBI/7OYrVwaOvJlxahOn2YozscksALIQo/X7KWkUlQzxQUwy+Z4c0UzHs
flX0qNC3z0mk+rZ6lz1ytjaWLyLhyaE9yPQffDgkSDE7KY7iFTjq+kCpotmixKJyautfYBjrUCqG
OWrwQVP+PknBtNDwM3BDnZp5C8e8MbHU9J3YP+mh5Di8x6e9sVz/fz5aLRx3c3bgF0ge9YD9+vpv
YqgJagxlXx56FAWEfJShqkRgBCDUjzSzgm7NqOQBgUty5RF2R6hHaXX6QGnMgi6Yuj7/xBtoIwCi
pNue51U7yRg3khAIoEbi0ILVu4c7u58hrN7v/uYC4dTlkHpBnZozeJY/47/dDt4ye4CApkwLBhSG
0qdfIBEEFfjomwiUN5q1SY2Hj4TvdWuvtlmQPt4LYVdFghU344CYntJUvvy/zWs4gdJvvn38hvUT
EcV6tUaAfteF+p1nssC5NmKXudv77WC3JyoVBUnHf9b95rrakp9Nc6JbrLMJ56muGMOqqsmOl9ih
BmHV96UNyu3H/WgtyljQ8/7tC6hIdLKrpHxy8BlrmwPssHe/5yDtved95u/YUUyCChN1G5G4QL6Z
plfrKr3RTlj0WlueOE2N4pEK/KHvVRGb0PucfFBFRj0WjQVLlvHyAbhs7vJ/MZEX7JPc27VkHLU4
3lvcUEiNzuGbILZzCkVYNTU5vTa/X3Rt8UA4zcMsZqOHmZZzRoKlPMS9ei+a24Tp/c6j379tyutn
qKBED1iWy8RAbDTWcCPoSPO3IGHS55+blWGM69A9fODwUaZU76YSR0vTZvBYUUwkz9FCKd4kxSR9
vbkQ/GQ5kpgffrOnGxq/jmdKcpfT63TrkUA/LTnTF95V24V6sPfSR/Qkk9H2aSttjgMPme37ibOX
tfomoBJz2q4hLaYKPf0EpyewdEkk1Vgqq/VZoQ1jQfxG4lmjh9lK9ANeV9bygpyZMmcHOWzBuoey
0bJGXLcmLqBJM25lsw9P/FREd4VUCmvN6wiRNRH9hTQtEOq44dZgIPX2KxYXC5a3IjCezY/D5v5K
hiK86DMdTwPChaE+VmcguVT5T+jwqVSRowfhsxeasJZzAMwnT22SSQsAACWvdCvN9IJ/LtDPEO04
NQgA0LsPKiaMkuonxUVBl+wL++baNC0IkLQko5yoCS3XwYpOheWJiK9xZWS1lwvyecnJydchcbpi
NVicNJFIODbXMNpvXllPEoq5aW1dij43UROZ77YpiCRpFSEZonYSANwnZjthafT/14MDE3dAnKrN
Y+EB3+P8ZPfJ0mcjNWJND1u8KJHQbpSUfnujsFZ/+xEjvlCqnT/tlOThGiQeZ4mHyRPB+//SEJgV
eet3qUaRZs0oqHV9QyH/qF4Q177mZuiccJjePxq0gLSyEF/HwBQ457eMhJ0bCdizCvHNcSqf96Hk
7lQnxUYMRIlMt+9IHWEx0lAEHRm3GenfWptOpynpTmHb7H5JBtbFcs+vDrNrHhbFnYTDO0HfX+6e
afZ6xKnZL8+SsaoIW81cGkPF8z+/Xq+tZ/MZhOcLgz9vNL+za1P8l+w/EQJLUthJ6lnSPS4sokwd
OqzS+LDx7wpMVwd3ExVgy3X7bZCtix/80noQVdmNl/txxyYBjujVMt9aQ8TBskpzjPadYoekLhlb
B78sVjGiH5FuR9iYzFoSzkNnqJ/9vDPwA/6vKFl/uHgXqAD/G90qhDhb9XttXkXI6Sj8ihFgukpi
cM8WaY+LIVLqFxedIFIzeUOad3oDjDaBQpbmS1IeyKdPxfc45a3CRcAUl5cA26iADbvkpva8pFPf
rKkFlStbwlP0+RYapsU9P9a+BR0p2xDuK+/ZbrEg6xXB2drwBmB6USlNN3iEbYW4XqYlckv/XoEK
Htuq95JIVlObr/5W+32FSDKbL919jMGqPXli2wwIRqKlcUVRzebSPli3t2fQEY5g5LnQSg3fi8kw
O3oReI7HgmGIF5MRLoeWcyDkJ+HAU1W2dH8mPg+qnzMiAg9VN6ij2U50Bhwl/6+zJVCPeYj66qwa
ZbSwieFL8eXHxEwYxdqhYsZtPxbkDHZsv6bBC01ahtnLcKBTEll00L32JEPqutNhWdyiCQh7PMl6
u9YDvtVMKNI4TPEr+B9E7hq3ZTV7xSq4d+YLD0z8raOnpDRejQI9KDBj8GSYkoIiukWv1dVBUCFN
Vdy9zTgyw238MWlOaz0afcj2McoEKqJJVfikAkaN2kCmFAGgXWli6xLRwXuoyGneL9XusPEg3fo1
KIRapHXy+aXHlAHnxYCQWHXc6hI4GCzZys9CJOajW+G7Q3YwQWENKjoCi0zU0WVSS8+tkws2nMyb
Q1nQ/A2NPzQC5Rpu3CxqOq5jrkFsypnQG7N+eJ3fqGv8V4Jm42nU9nuMyVlr0oVM2ZgnI3cMwg+w
R19yrg3CuNbSnWpjVZ2exx2W+TL1MZQDZVR8xY0/nHHCSAi8L2k6TW7l2QZzWGF6FrCfXNxvL+a0
QOA6wqhrTmcAD2CleFL1QJC2yKAnsPHwqo5rxHCIFihG9VBl6N0Y8/GwmhQ6Mbpw0ghe8kPKgjvo
BB65Nc38rmue0HgHg9riURo6J8awm4g4uq5YQoN/hxmzRY5Ws0IbEgm21nF/eRq1uy2xOJjRLPA9
wToZvR8MP9eaZIySRBnl2Lmdu8rd2RHIRemnXpet4OP58lMFbGMRwn01PmxTEuVH8W1FBbcswD4r
CVozGERKlPFdG4e6MXwR1812MIUNX6aDpcccobZMN9Ys5F+4cMDE8HPKoSurkfFAtko/BaGdhEDX
Bw212hoQ7DETOj+jeG2SUy7Q9h+phdj6znBo+BhafZ1DricOSf8ZO/+kIBSg805HoqOIJYG3K3cc
XVB8aZDUhb5trVRbjV9Ug1QMZkJWhcCo+e0kVaN15qiTFFyH1VdJoWfsIthwyA/falWE0tXGBnOF
ugnD0DTc0MALcg6EYv42pp6y2Fgmng4qmbu2JopIhShzkSwNj9x0cJv3X3N4BNmSDGM2LQfRu2b6
tTuYpAaMG5WNPOKZ2ckQT/SH28Xz7YA+CvXtJF1tmZ8PkAyXOgVKljF37+6BPz8vxwf+lnirYk48
B87OvIk9f65lsh1Gisj7vcHVoxh0C9/nSnzzhV6KtIkcPzg9/UxOlmMpKKHtIhkfui1hIdejceDm
MB/0miUn7B+oe/n9ODhUOaBoIEsSGvXTFRa3+oO15q7ugG1YnKEswq7EFlMroM2yoWglnBCtgSYp
yHZvmGNtnVEbu7Z+j3zc2elqpdFRqdvJP2YTBG1dAnUcA3TfeM6ZY4J2Q2G4F59ltjpEMvHu5sb0
rX5kU+lJ7bEhwGVGy+ysdOJa1snzRLHLM1WlpLZtTpcyTaBs5+jrjhVU6DsnzYZSW0je+p3wtt/b
aEmbsmPXsUIoUy6raMq85qgFn1X+BlG1K5hWEzDsw9UZJKBBN1WFC5Haz5tt0ykpaceM0PZjh3Ie
s4RHonV7dITsS1229tu7Ar/y7VHuWt08N7z65yfiJ2drD7xqEkLVieXmIegmPCy+spZrQKDObuW1
CPG74RIogatbJWrhA9QCliaRvZzMWscUdeLQHB64evj1C3755UjGRtJNNUy8N012TRW2qun43vdR
MlhSxoBR4QAhWCT/rrHvuWZC/D1kQFoMIsmJcijoa2DGpQN18uR9Yeb5RJ6da0Q8d+OY/Ad0tnDg
HkY12nb/6WnUaz+jaHzAl477jPByBXdwqFOdi6S95d+EdN7rWJPHv421KE1Ml64eQYBfhsySZ1Xq
Ssqa0dIfbd6U3jC2T0v7AEmr8kJtDZ3Bwy1P9mmQ7T7CnUICdB8Y2W2yUMWcMaqQii+jIeVVqjRC
WiHJHoaZO2BbLdiU14peCkJWWNyy9Do3c1pbD8QelLoYQgxymkzFSQjb4mS++0Huqja2CmvH/HgF
VqnvkpMzy8QrL/hikDewOCzDv69WiWHmJi17T7oOFMCFjf/LoT776f7qZtAOAU/cECoZTMFz6I3k
83ryEt2jn0VCqStPNjlv9htULKwgvpADlB8ZbBUk+30IyuWWLUw3OjF/anvtJVqtlOShgQCeJ5n0
s/vEh6ZgDsTisJEOgDJopNhEav38CFqlTSqye5sjzGwmJqsOV3mvjFUzZFgbNmv2E0FXbe1CR96h
7iUMN4+diYo9YMcmNMRe0nQt4+JYCvw8NULW3r6iaKBk3u2fej0fyYDrxpZMtFFwSQrN/DodDGUN
SLPOumUtchjw87R/4Ax0a7S63fixASyzcPDAx1zFdq/YuxB8dw5I5GRSRzmKx4DJFEMB4ZOYMTwV
vnQTLcTbo0osmyoJs+V4yjPnqj8oOcxtQo4UBbjPa7UV5eqzrS5oS5glCZCX66Y7hhB8x4LpThit
8vUL2KTRj+h6/kAJ1mHFkOpjh7YoXaVYK1ou1+1dNOzhYol3wXCYg1mHHf8nZif5yzqmMbWuYMVf
gz/L76ZGFTK2vOJJxTmPFk5UfnUQ/0epNQfZlN/1L6seX29melHKV5BVeuYWAKKQcAlqSGtDEufG
POk0MDRoV4Ampz/q24d9H9Eb350GxwtBBHRbwSGGdfAq6340JPj+FS/qsM07Z6N/AcJcKUWhuVL2
xGXrcToTutOzRNyI8R8qzdrJEdlc9kXKLUzi5sIRhKYpfaLPvnCuvDjO3KbxmOr1emw7qg1VNQBt
HJo/2+p1+LxvvrwqTthOanEgzW/nl5C0IoEhPa6uvBmPDTL+6Lx85gxw2oj37xgRYMXBIVIJEXA8
OjRBw/PVcTIaeevJM3uxLltdCyaejRLnnxCAtwyHmDMrKITFtDj8+Aetik2/2VhHCc7qZqleQZVH
7iVfP4y82AP6cupkX23+Fym4xyDaX/TfkTaKTczUgVevGJykSqlz9GQT9frC/9JmVojEqcbThwQo
6fwmymON5+6vQSMiY+dBJqKamcfmhHUtqXGw43byeFu4XmP7OJfX6M/0E71xlSrjGrUByzxB+1Nf
kv7YQGQ9DXMSBthFBVhy3k6otfmduuZJu9OJ6qMcynm3kg6n+81BjymisMSFP0RR4W8D3Frj+MYC
38f3R9asVxR58M61sqoHY6/JhSKnHu9IxaIgjrF8WqsL0s4df9SBYpvEpZlHlB8j6w7Pc//m6CX8
kSLokF0n5JTucT0kYKIACUp8TqR26khCju42N32lYMOqXnkteC4FiQSC/AdipDIMF7nL1BliL+H7
9cOIsQ5hsN/7cMFSN9J8wgdJwL9mQnhgpm4mZ4iq+0RPVFoB4+xxWNycwYfrRLMR0hvr4mDDBM1E
uLWjkkZD0fCGiWmG5lOwr7drf11XnvxhK8KPdCQYPP5FVrM/cD1ILXEE+jGljXcHRFUym1XVPrkN
eLGNn7pKgefyyziA1c2sRP8on1mk5/WFw1Tig15h716DmhuVfX0oSADrFEi+O8Wo/MJRyAFcqUAv
c06WnMUukbCoTzXzzzAIKtOLQAUENfp6tikwZ8D84iIEh4bxBtUstxW4RwBj3QWwdGD1pPmHHt66
KKmYcEPdEcRWN+yjwjvjjPGCeWiJgIMw/9WAYznI7rFL/K2iHBPIBn9ZyO5pHbNSAHp3rpjAF3UF
fBYvRD9eYUrJSOBLgroFuG0VBFRS/YgZQ5JB3A==
`pragma protect end_protected
