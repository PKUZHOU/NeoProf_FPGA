// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
uAf3tnLy61mLBAZo/91En1Pt3jbcPhPfn8hoY/eIVy5X6yqVAp2TzGVbPJeF
OrYLK3DErzYtt+bA0ELDZEp0Z9/yRzUrhKg5l0XkSfuOxcDDvzAlk5R7wR32
BL7lnAI/rYVqNi8nnr6UXTUHzfribSRNeaBXxLYvL0NIQhvjSFdik+IxxyTO
u5VouXThxrxijwvWAFdaIw/FaUWTUeH82wbFR0eGqnoIk2sjFIe8taKNYMUt
h/CzI0FOPJtLJMXIAcsdb/kVSRKbIT0/Bl3vdTPdbh5O0+awms2/lJQqxvct
1YAysu7AjzAuv0pCGjHm98MOkhupL1N8JZ2/EE857A==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
lDfRg56bmhQFp/F083rQ3PiTNIGqlW13xu2F1u4Cntt0Lbj90i30+IfYZ+LT
hOJvTRvCjtJgW6tEEBwlRasyv1Wa6ByxXk202bPER0KkWrXTJLxCsJ3pBxKb
hkwrCRRyM4cYSopa5IewRrV0PYyeLX29+tctGu92nawCBmJwBYbVGDxPfe0Y
jmednJm+v/s6dbNHPpXE2462IVAZtXHh8uOvW52A5hw+KymLEBTopbneQdo7
b4bfg8xgmaSNOFqJ0yFdzCVChRwQlIVnlR6CNsnhherkRCofH+x4s0qNJso/
T5L1H8QB2RFObYOwq9TnK0G+IJvgGjj3eeU1RWD+pA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
g8LKIcMhfn7fzngdzAjGCmczq3uDtFfhqVxi0oxvWib8PBOOIDa0kX87fIS8
guvlIEPe52DCiYIDhv31KOuzwYaaAsSWsS44ADzp1zegXskIaxjiyBjssOkb
vA0dSOgQxgaXFdcZu1z3PlD2cvoDliYQS58da1B478/13OcRMZ9pQBB0zHrw
lRn61e74KlP6VNd0PbK6eIA4ulHGhs+AdJFXqPUuBa67Vl/xxO7o76yweHeZ
Dox7PX3DSTPRTUni+em5gLGz/pXcNYLa+5RQ8IwrrCBGWfNhir0NYZ0h5a3c
lfPfUlDxBluPyYZL5FJHAz8FibN0hpwG0SSQxgWPqQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FRdq065vqv5mRW32VQ5ODMK5y5EYzG0EREBP/Fgy1w9CaNgEMORZYZhostDv
NbUwp2qpH+NxnatKHlwalEmTXOjLP14eZVD1n8djkB08oJS4IXgJubtpA404
WXceZ3YosJmJugjgHf3gdY2fOa3CUVaIwCLDavWmIcO8OtlSeqY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Q0lw397HzdsexTdqfPj731n9eJ0dlZsgshU07U5rEzpMxWw0cXCX3ViKtPpw
KE2IBglhjtW4vAjTotD4INjFbaZ7kw4MrtXtwWyOOcjsg83qp+dZwBOSodFd
cFygCqaq1dI4HD62roF5ajx+fpfQNTLSpJ9d1Mew8y4BetMcWSoXt5BofFPH
EnZwcgls4zTPsDXkY6eF5r/oRBEoZ6F8FObnrY1ryilw8/sKbUNBDAO7bltK
s4Y1iS2lff9dtik64tI+GpK/siAg83ha4sy+jaaDct9um1W2fa4U+tkZUA73
yVMvAG8Q1hAw6f/EkP8spwcZH+xabHC9+GWfGGVA5Wzhal7BFQ5keh+N1pAX
IdAh0DFNrVko5J3tzIkkrW8KOA0woKb/PE2Du1wPWdWdNoFnkuXLfF3MTFvt
edjy4wBxiT7Y4owlJxHfdyb0w6KVuv9Qz+uEr9XV0BdXwZpWOMmTqJ2BTwU8
a4fnLsEwwslqcdsBCkM+YjYfydISJy2E


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FoiRur/Bc4Frqh1qJHh0oTGux3Vlmu7oAIiCJhCil+PwbyC1CtybFxC+1dyV
0HS8IOwaHIp39SjMAMtiUQIClFKqfVa03ela64DY/Sa75RRTiHUrbrKQJ2h+
sFn8sPIfHVrg6k8xmnSzLQX0ilIVd+3SSfSEIh+VsJbMVk/xfcY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
DEtggobUc0BINGy+JAiP5iTZ4Y79x5LcZcJDUWl545jjzYTLJq1MPKHvUnDD
Cr7oOY0JapqdegoMKV2adnigioCA0Mc2lHfPPJaaqoTEh4r3kvIsEYkNuLJl
Liv3Z81/29CmZhyEhqQo0TPS948f0awdIxopzsx8FOmXLgdotGg=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 10816)
`pragma protect data_block
n+VRwx8PwzzUWAgknU+D5/oNdxx/GqNI89sXgvNgt6wwSNT5ZKiFmIJs95Oa
fo8DHlJYZpz1ckG5M29Okz0LakaO1BxvMcx46dyAfAKzxRgLg4I3BDoNu2FU
tpzzlO1QF2hT5alpqPmnr66G0h8Fgz8huP4j7m6KIkBKzTxksqGGFDZcgwva
UDTbNMrv2gQhPaJddczWyAUxE215Wtyzc2EGQMkFPie4D6qKCiNfUy3K2eqo
E9pG1Ug4Pb7O6CyGCwYrF3waLyMsTGz0PZEHgq6EI88IpMdsiYPWAgp62k52
xSqI2hU4zARKT65lPf35fgcMX/QqLeJMBRN8/XHUuGsvweNpygAvlFW7vAtO
AhB40mNqkmKDq2jF08d0KXoqF3DQOYcCj9Zk0NpSJ7pj4PJdOCZ91yE6URTY
tzOIIgy607plFBssABVQSJV+OC/uDzj2O98PwmWv7xRCkvCcoF8kQujVA08B
zGQwgSxbOR9Ke/lvpIPiyXRSCY23yjDjhvBVuelfkuVvTZOgIfYNLLfcsIKO
942WgAWh72iR1igPBTbV140QNuqqloeP4wIFh1fDPpCOaSqWTnTGDj4jDFzr
c87mV6Daqz13F++5R7Dr4HaNNySKSrYCSJj0pid8/8RGOKaL+7sI2hnRGFfo
uuQXSEUinJ7fScb9mvJLzMlAQakmrxn9rVVXJ20gX+E4VvGOhIubQBNBvI5j
GMpHSF72frVAENn7xzjdhHBF0GUo/E1Eodb8T9huXTOAjdkFdT2WFJeAVgQq
1kuwdMmcSmqiggFO92e3ppep8rw2NvyAtJOMdpcn1l5I+DAUqed6CGbrzrjk
mV5wLXwqC3WYsKJF1cBpT+TI2GUvhxYI4Qf8kqTFREVmsyeSKKDyBBFsMqrz
Dt8c0D732fJeJuRzVUz12dAmaEQDksVorHIS5HeQ/pc5L9HVJhZQZNw7aG0V
JXukNEVuaTIj9AQKTjzHrYS3QOBKwRLOptPeclZ8uWkJpZrEuLnt95/hxnXY
39jpmw0MUiHrgps4y5SkXJnVVr7mF0SlVtQ8BDMOzp0PtUjyx9l7aXy+AKd3
h5SPSP72LFHSoaf3et8m9JO1AXrepPM4KJdr+sGVMiBnbioQd1sJ07kuquNq
6IP37c9lgi3J76N7ZavWivPoEiyuQ6jbliqO1TfQAIps2SXE9Je2hYkUsQ01
v6vAyT/bJpDaFzCwTM21Vj3nZDgm3qFW5KJaHKwgyihazLevFGbomC/FaGGO
BG17ezvitRAJfVqPWIfXBLAWeWbeu4ac7VavQXFR4ZZQipzQ3nOLKx31X5re
TXuU2hBcJeeFCrTJ/cFaTYxON6yk/VLTFYY3KRv7AKqpb7Ik8r0BI6Rcrxzw
jJwjmBsrSJiJjZ6IDGL4BZfa+T4TK/2ovSxAL2KCMgxR3Q5W4LXF5iLI3wzp
/Qq1gzHxyhlg2TuIzpB5lCoJYGvoEgCFZ18MnogG23v6d/F9upN+FM/qSkCh
E4//1ONO00hKmlXZqGk0XxmnGIprxLETtqj9Aqh2lPnkWJ3DUuNhtAJV71Cg
hh3hZwM9ajb6E7xFYyrnF4YRMBFnsvlXYQqPCKPfGrsYVNhwsQdCJnr9ets5
pS9RprZg6a7rRtjEaCRtd3E2XqbLfSnijWMS2cPLX9/AUHdOSGbc1UcYK5+6
17UtDO8t+Ver2TV/Sm/ELraXL0IzbPyQs1d0pycCrskIoFYgpztTQpHhVtoj
9S8Td8n2hh36XLFaxDhaNiQXJE4faJ1+tDe+yDQ5eNtEs9De1K30AnBxT2JB
AE/6IfR08W9kuuSW41+0D3WIRidUWXACZocJOLGAPm4sgti+Bn0F3jqPxRyZ
1rOHUuLQXNjmGluCDhEuJhdsLfz98GhTMuykopUk/NbdvlKGxrjN1IAQrfYy
zAqnkG/yC5YfCyKcQid0zqkimUd3onz8PkiYq/DjyJ7B+Dk+KxInSr062Tgl
Q2M9/743uirJcsqEFf5SsyntBxMLLpygY+u+mw7hmDUAuOv5wI6fGsRKVwFP
xRP67fueF/qS5QcRFIwKfT+LvcUbdIPhf8qfSWKgZeIvEvHaveB1guXUrq9P
G5yLzjEGbGNKGDHvB6jqh4iisabwxn+hPaNwStGa229+7GERvj8kv32SxxrB
2m2jCFOclmP0KRjFy7a8im+2tctFj2TKxNnWFwL9NCTwngTmHfxCc5Xezg9H
fPdvuxRvQzNT03Ze2BNW5WtZW/Qm2vzwODn15y0SfMbkJnXrCEixht4OLgm3
fKx66c079OuZfo1DNDlvq6JGZOQ1rnij7RrLbZsgEcQWow4S7wKAgcnpMz1d
xHFo5XMPEephlMQYf7EiH6wGmgvKc1T4BI5KDWNB6k2nNqZE7iK3DNDBq0F+
aWjJnJ6+YIrxKyC1VAo2JpAKNO+MUu4GsC783tfv4Ffj6PgAx6nzxO9awZbe
JZjcUqxJp5ch5Uh+56splvqbXLi/k7uF5XOYGVpUGM3/VteKJGTkSPKkzOKx
WqcWc0/ak0HGsZokobRS8PpG/P8t5aayN1yMQByFKeARQ1MZXgGmC2tdYL/s
F/ZzeH89V3+EnXjG76SNlwkZSEKOojd3aU4StArgsMd+s2hjwsR4kpW0u+J9
+nU1jCPJnohoH9863qzGUMN64VuPaS4zck2cRMAVZscz/rPVabvW3OtjSiLq
eG4gp2rK2c22LZDfyPrw9Palx1d9HOzryMBxJjq8Zvy2rJRA6OWk3uOZ5/bN
WgnqMlD6EkkQhp6LmXA+0ZbbT00Pnv+DwzWLiyff7ppLCZD8g8LBBZQLjCDN
aADRG9Xf7yQRPE37D4cJ6nbJh1l3b31V9L0RFIRJsb2Uq8P69qKVk9yFFkXP
HelP7SkQ2rjGqgZ4N9dGvtH27iaS+sJIpEAj2JR/VW/FQzlWia0zq5YGjbub
8lL5e45efecNi4XgowPR1BNRpznjo4qtFOGLCweTeGU72O6U9ErTHzSPPw6J
4wQEVofLkSNWadNALVL445FC3dK5HipHa7dCm6TjbCOOBeu3CMmuR39WreLP
DHcS4tn3uPyUhV/teCCfMe0fhkTWma3sCtfhBbf2KCKToH7/Hsf3krtKX06z
ET0omUJHqARf4XxA/9cqFnja892ORvNmiQRoHO6qe2RhJtxhF4sqtPnIPiH1
kFYHjr2ydBRkuTQOcKFXtktpQElrCOMEysxPP0GIyYiCb7HKklQhlXAmnAL1
bIFt3Zs7Svl41/SLQU5T+kAIWFOouOARf5hHeOL0z3H+GDkdo15VF1u5Q9PC
ffC7vwasLMNxPMCF5egXJB6N6y8d7QUDZU1RJmVR5078eF/4edkLfFpxXb3r
plfeZLMpP2Z23SQVGJF+tDhz/zl1Js/457qyw5vi9x7m7flLJdbf685CkfIj
2LXJ5XuAONAsSv1aol1t3XwZLqsUZetDRGPjvoH06BgUjDpyMzw+OkWMDEN1
0CIbzG73FmSo1nkxoRcJTJLiQqojt1G5fDLifMXwZ2+90z783uqUyqIFJPY2
JkmkCd6Ab4lSvTSMfABMs++d6akv4P5oNw/6R/QIGDuSdyrEgjXFXlnonzdE
LynXrCv65hQuDTDOsxV8SQ96zaKkJSb/keVSnz0FXAXIWgvBdV/8Q4lRwGx5
6it58+k6IksmaQoscAlC2ricVBLCo1YTzEHXNgxFwoB+xUoRQfn0otMmKWEX
/rM74Z580Om1KXOYHwR2j0zZUpgXl0bniiwbK1suRDq3SeZ/HPiBN/62xctO
keo0nR850k3oaloi4t1nDGTJdig2y6gTPPSX5T3MsheyceJHnJ3ZgxAQx1Lc
omozs4rN9jJe7TWf29x7KxC953lkdhVwJGcXARBqT/n31tEGKG8W42ll49Ob
v8MZyqEDVof1q9KG1gONpuInduDrZbxywZADc5FM2rJ9/wnpPAqP0a1D3NV6
cTZfA06P1vdTSWSFpGT5Hy33BigHnErOOtKHdlCc7lna2I7wrz2A0JE0ihgM
vqrb1Lh4SbL9PJrcfrjxe9J0Ax24g7VEm8ytBXa4rGwAI1U6SFTRr3YKXHMF
pyk+Kgx4WUYHMEmUZekKuHlmt7PW3TjXJZ1iwasVmQnnlxsHV6GRdWU8JOj+
nw2Uqj8NblrDbMewRDl0XGZzwqHfuovDEaPFltK84gckMCGQEZIFUx3fLLxr
TzClXhF1ki0WrukCz6fiFnB4/FYfgTeY3ncxTMpuo3UA9O31QNlan/gFr6ay
a3AAPpvnovhcZ/Thpi4qhCb0e2eAK96NG6Nr4FmlVTw6uMnRuzD9LCa4inyr
daWc/fXQ/QSH3jz4lzK4q6aNSpB+R8cFXk6zjdXS3HKxDcUKkcH8qSp1WQXS
s3ufz7LnesWyRGZGBvE01MUbCCAtDOI2LbgXinRi8LqgNp2L1R3wDKSJmvQe
1H8BbMW6VPlxMUSRhI19+dNt+7TvXpIH1IlF77cUZ1QqpRbQaLmw0KDon8/b
tl7YiUBpIy2MHo4/Zq7A7GMUhFNUL1Ml6MxuIRcDfeMxQp+C1PE3Ldn5UQAS
ZComnNxNjHkPz3VSRSLE2+47jUeLLxpxVleg8DKM7+JqPbemKr7U3MaIZiSZ
g9vrnm7OsFVQUVG4yBRXdsPeQRCQCQU7yjmSEVTrAzlXe+3Xa1kR89wKhOZe
4HUAI6irL0iZBQhPUB46A6JVz6KS+JrvvcR8YngncTDX5lcfMaMEBBMbSia/
upIfOCSyEaly9D0WX3gKZYPnUiWPP4Bg+OEnSL5ZDYd0bNx6RqvNzCVlf949
TJN6+Z1ZdSrucII2HqcNKRe0+H033NmcFUJtRKc0mtpDECV7HCOosibXjUri
QkxVQUoaGlmWPK7s9eiIJ5ucBtRuI1rhPrtdOzoktgg7lqkYt6vHbbrpfSTg
1qcy4F+picYnPjK9zTEyTIRDxZY5CVSkmsjA1BHX3IikbkgU6RjAhcBSNpVq
Ho/5LLwNgE6Vfv8JN0pxo7sWuu27ByOGQ5ashIqGlSEm5zAKE9StXojtWd4m
NuqzvvP+4KvMtA7EYKHmP2oT8YhkyyvC19NB7Q4wi0TdB15SHz4lpnGqWqQx
u+nNm8Xku9YjugP1O9l5TvLJlFTLG9qwuuVsFNlgLFTZVN9CbjNyNzzUzP4g
xd+3qfJtSuoHkkX+JUDIPYoQvUjwwSP9ZIruDmIXhREvIlfcjiKvHCHzOuRN
NpNbT06oYv7/dtyaqXxCBJ3LLq1A5hWTUlMG6SpN9f7/tTpa3zac5WV0YtTA
/iEDeFt38Qe9ADyAAJlzMJNJdZSbRdOyBQevH+k5hjszGn68aEEQUrUUJRoQ
P2haleu+pEfv2fvyfouRXigpnZ6BRPnAwHH8BVHfQH/nMu8GJBwcqhLo/Ern
R/emvZ8jY/hDinGg/kIhzyZevhRKp9EO6yT6Hlqs6dNUPC91nTCvnljye7Kh
yld0ZEcyRb3ktLLSNQiSk1r9dtlI/8mZixaJEfFcw82eCb8ftkCopmKXO6fJ
bn8qrWAzsBU99hWGHi+pyjI4uEwjal7ma4TdZvYSvU60ul+vzSVRyuYVMTPv
0OhfBzRMmRjBOL4YxdmqIe2moset8HwgDOXioS1o8DfdWL4JgmabxVfJdQYj
8Dkmhq5Hsu+4B1/0bts3MnnxpAMkSh+tqFdwNyA8lXmPYWgwo75secjc+OfO
q0IHhuaPpoVtV0MV0B6xmghY6Z1marsm/9jCX/YK2kbAa6ivLZEZyGKRqFRa
RAaHOifxSdW9n54ivXOYstN6TUw9p/fkCgUklfsmWWAAWElX4hdT3aUobzkb
Ls9Qe329xOtH8SMnELfWWJ6YY6yzbv2zXGwEQToG0AydeVDabtG1Hhx24p2y
STlVm8sw2l/90EjHjOeinUrfuU4PAoIyVyyMia9iEnzJsJsuUp+n3qDc8OmI
ZjjoNephV4NnFWvd+gkElEC6hqRYmO7+AJ3FQ9XEkE2D3yfcLpapldRX+hXS
C9VGksi1Hjco5xYp1/vAt+REzDZOxsn64AgL9dpuedzI24/7KEIgsg0kx238
DYzZcMFU3oQNYbSQqP55A2Edd5trmUQa6U3vONkFe4FQJPI7cmjzSuLf/S9/
TLEJu7/6cf1ZOLeygibs39SY7gO0X4SDXBkFNCXHTUC5Hrp0H0xzPHYzsQ0b
FFygKKih5ll4GAydNBYHW15Lnyjbnz8vcRHsunZfWrvz7dN223VPFiR63XEz
+29FSSP+TuIdQ3NkSK1RUJnqyddlJa1T21QRyd5hCkzpSs65evliKYNhrdZH
8ZOGe5pV5WlTJnPfeKnURZfwy0gPVJ5NiB0ARih/XJhSQcYCoMh6FYl//il9
el7lr3KIkTDEfLOgTi4PVmLVSRcpFVkkYUdRvUPcjRB9M17wRh6HscUS7x1g
QrICWoEoAeEbipa3jW8UJbVDXuMbELmlalWj/so92zLmKkhbUKhfMSGH+tCN
943SJ+ENDiQRpbi9fMHdhvq09gxHuXNvLNtCoyOhUO+vo/fcp2oeDqHiEvZG
rbBPjbZq2VFCAq+tCcyyZfMk5VK3tibFwz1iOoFgwf/5A/GU7V1Qrw8HuAEk
AtZiESGhLENtWXp/MX3/sxnCOs29Mk1TFttMQ9V4AeICmeklBH/n68iZmhU1
BVBdic35f86+YOp52JmtVrW+AxizVVGIswCJJn14/8GbaiC1K9v0l6pYTS/X
bMwK+YLnoeFhGE3b1IzTtmwmgA77eQ5ZamgUPrnRxMEA5s+QrgESgFx2ouxU
NS/BoAIUG1zHOvTVJ9m/Sv7OPAtANiPTNFPBQaJ5hxBWafcf73/pPi3UhAp8
sBI5WioDJ7VSHZ1OUUanxQwBLRfbEikgoN4HxErGcV8vWtZjH5cwr321udqM
4uQm2xl4IUZYVoANTiKcCzRo46mQQI5UPW4rTUfAXIekAosfL6Vzl+utwTld
iUZe5d9vUYoApYOs7eVv2Mjwly+4VUaSF2IYFHX5m9PUPGu3f1WhG6ZYFKx7
MI+gXvia6Ng2HunDfoPRAufGyv8+a4ARicJxRQKY70iWxy+GCq9/FAnEhsEe
1BOZFetbgVUoKGkp2fYtJOY2/0k1q/9UvWiG1mEltOnzYtRv1WlIK5zr20n/
1jYbaJDyLGzGi1LVzHCWwXHoEOEmU1fpHMdN0pBxW71w9UHqVqpwS9J6fev7
J0XW9JBXBAAcrNP2ZGM7YDHqZVTpMiubjGMgibG6luasuacyz2sDFaMM5wmI
N5/+XPYBHIOMsV6dcPX0LJ2r7knanHuA17l1R3jdAyE8vR4oGcD66fQDm89E
bjvrMtNR5mxrGzhZP0j+8qTQpt66a22JMlyK7sH5NYYdyySJUhluxrYTIdgB
ubxVIXh7yCeTWOPLBSKdJxZjq9UHmeap2pMmdoJGtiu6c+lDbVyRrvVup6d7
Lyw+oNKWGtsnKZBnvi7Yy/ZPBVdspCj0lzk+wyEDDiyi9woCidDf+DowV/dd
UXf5S3QhHJmIeub+lYmNFmaYhLWUqoSuXyYsFC+j/JX3IHeCpdVQ6EoiaKvC
zL+HCzqbA+dO/eyIfFgnU5Ke+m+3JxuV2q8Uxrs2sZvgDFLm0nSZZ3nT4DzN
HjdbLnvDIFUGYInX05iuhke8MFPhUkT0PwopUdoqI3Iyt7hr5rldwk9hP2xa
ZFSpsxEJut5Rj90ocQ6sZ9DyF+WoGC89TYmKnK7EVP+T1VDfm4iABHtEWJOO
svjG7OE1PHo2RGoAF/gusuxdFVIW9qP6y/TsSS0r9Uknn1o3GKJVhsXjVcTq
+aTH3cf6LKJ46TnhDmHkemRq7ZqXwCSLXX2DjR3Ex1hJJnbhLJd2NQomJnc8
YoMlBQpveuoVwpH+sf2UxkjpZx+GQo1C/kH3ZnE8+8mD9pky1S0FqBuwdC5l
mL20pX6RCF+YgDKn5FNNzibcL9SH6s/LPtsQnKgDa1RM33EgQFwFKVfLJbSo
cuK7ejLeiy0qzFYRjO/kL2a8UubijxDN0DfmzcckY2Q7eU8P7RRw7Xtrpqsx
TzRvDA2tq8mJUNQT/+CuEbUQ6yO2+1gcG+3qXqM5prmuS7upp7P0rKlrGeLT
ukFf5YXZX2QYX72XFO/EXq9s94+AqkSEDLKsVsU++ohqR96Zz8e7ROrnvCh5
Xqy8DYEzyCZbkmIUiG5K7hzTO8F6TjoXQLU32De7g0JreOSd3lBvQ2o/g6Et
0MlJi7p6zMSnelucYEgim2NeagV4GGFWVM9zNOKveqqOUae+UmeQFcNXQXRI
u70/sznO8tTfI0VJexcFUpIa6WOWmQeoEtlts+Lm2ily+uRBYkbSjJV4+SiZ
tBmvAZWE9ieuzxBmOfpXoj8SkGk1ilnwNUREPaaYyFz6FYRtvrm03/py/k4K
M8EWA0PoJ38ZnpNW+58nuZCyTWzYul7McGjTD4F8Iz9C1x5Drte7hMa9K0xD
pg+NFnWwms/aTvUl3jyW0FFqkAGd5deaxqmjmQOe5griEG5QGqp10Bksxh8T
2oPJuP0gAsXQX9gqnu9PrSlb2aCg0d5uucyEMRYA9db9KNfCgM5n6ARifdCH
cL2LfV5GXuybVEEDmFouvR0mHfjUy1iNnGDvBtGef+LUJbFIIj/2G3aPEj+Q
xitiOj0cM9snHYi8vYk86G39Mjxo8wcUeyn8NPS/moood9ccZ6owUflTYfuW
gP1MO6mj4ZU9vqjE2tzg7CG/kzDQUUTPWRJq27erc8U/n3yFdEvHMt0wJXdT
tDISrjZtOUYTLqmBDLu57tObdKjzfipcClt+BCvaHDwr1gHDdEHI8l2D2fVS
qj/7c+IeihIQdM34hkWKzMnrP5mb6vDKzELkc//UHjTPA8tSRG6txBVg2vO+
ghOW6NJWEgIqn5FiSmsYxONQg2d6SvVqP9IUaDSyzj5NUKVFwB4DXNgjiuTc
KkIjD8WgtmEvdx73i0VPlnADWiluSrY4UhDu5BY2DnoAeqC47m/e+NgRnuPF
T1Pwh8MvQabmD3tyCy5odFe9I01mPZ8JRlxCYtKCg4z4TjO9hjl1SrDmMnnV
gnhVrO/46hbxCOmQ7kuoOnZQGr7VtArKUwvsgB752jPy71p9q4X2IX3YGCOw
FH+qQCji6n8ppEiJ2NSDSYv20ORb6FvZqdu6rvMJpbjRef372OPq+Yg4tfKs
6SroVJ1wjMm2I1DS5Kz9A4/lhxs+bKggjZ3YglxIK3k2c6qkXCFOp1mVcsjD
vlUEABo0x4CUKUtzn/H4P3GWcnFXQiRtrtbykS/Psg2FVy8mQop6RH3a+RJp
4shd3wtQpA/s6a14BSRPfnigF5HD2qbHYsqRiTbcvFbfOyfD6JjyPAY7XXnz
9cwe55jjROSkec8ia+GIvA/t7xzFExjBHu70cWeX/rPJvZE9cJRsMaTKT5kh
cWBq9c8QPqdMxx+xoOFSmZA8kpuxndnDOCDcCR55INDRkjyVtnPa2fcw3aBy
Rc7Bc2hZACEZtHcxd3VsaPexa2NkNR8nR9ZJheMB7I/Qeuq9Ezimo5Rc7dpN
CHuIKGxF5JSyRzN3SpsOTjaEq+Pdn2gMsau22yTlUWf3PZc5uE6FPeZHwMUt
A3YkhXqYZxnVctIqNLYykbHCA96XMzyKGh6i5j+jU1tRznxgj+HXbwrPh6v1
twQPeOnTmtlOmHORvjKoyfukccIqHV2N7JjhLN4L7g0cKGpPs0niQGDwdoHF
zLezh8Vvqtp24C+nLhthTuyRQbqxwZldu2ImGG73Nb68GSyhqHeGXoHgbXsV
hDX8eFn3Rba/nA+PIqZrUa620KXhz31hHKzmJT9vbZuPOD9swltwJgdF+Oxo
Fmtb8NwGKH6m7haQX7VvtsYMXBEzb5Cx3FllcBvjkJE+8UIF1sWVjQNbkhHo
PeDMA/q1zSXqeYetJCl42pS1NhblSfu65QX6wgpMiRvwf6Jt2Di2Z2MaQjc1
DEMrIvVLKcisMTp3q32lelO/w9l1ZfHb8p784CE4R57/obIgCIeeXH5nTPRF
W6dInmWEzeZZntVhSG43Tt5wYledb8DuLuKDK3MIXeQElWCGDNDUEq8nhBV7
b0fZy4cQFc3hhdCRoVM+0E3GTpe9oO+oSZmka5GiAZ4Qtm1zNkeZ4GLTha26
gCsjwf7WXUWgwTc/q/Y7JbCStYzS0iQkhwL3x491sCXHehu/FNw5ItuBMhLj
4rBuR3OP5pJlhBMVfnKOVHhM6UuN3zOtygaIMtqvz7TNDPFUXrU6mLpqfTO7
QkB9LNWNIZVDAwYkpsxHlIGYQcf2cPWFG9h4kMXPgwW6kywAodwPZoWC8Bgh
k+yoxzzr3IUjvX6/6MbCsd/cghMHBvVa3Y2gPtv1jRUzy0bcndtnR8MjKtBI
sUM6DHi5L+gBNo0bjyxCHetit9YltThvadzBmdOzQFG2JRspZlCdVgSeopDE
xLmFc/KSoqsYLxFv4cGTbVpEOx3zoJh97ZUD38RU1HmoV8hiJOLgcFffSyzr
OyGpSgPOQQcYKCXEDRyBKMr1YRc8estYH5DFd0igFu8MBdTfh96xOajxKtBV
a+ZA1HRRjWIgA5sqPCYBTDjlvD5lut9Qp22bliIF938VGI8DycJysA+wzFz/
fGBPCGbEh4Uud4DL8t1g+0OK+EKoaHfjUZ1vvQR1L8Ty6SCFHP+TRjlXn7CG
Y11aoZ7CYgxlSeR2P9F87c9QqPurzFa0CdO64ESxMV5QDzj7WAIYPZiEG9BU
X1JJIqN51XEsu+wgfgOXuqO3gKugVVq8I023JLTQAg/0u/JGoQmnrsA+s3OA
4hoARKVBqGnAzv5oYyck+AepujOsSL4Tk/YuWMsu+HCqiwL9kFCk0tANWCkU
VUfW9LQkiZE5T3hE0dwQF5V33cBL8EdbOsdULWIBbv+Mind1wWcQSiLj55IN
o+QiMk6qIAxG3ZzmqQTFVmjupUHfcvTG1ZG1OOyHW21xISMw7qYYE27lFr40
ntUoeWs0WGhSXSUsNpY36wXtopgBHLmg0VOATqPJ29Bi/UUC9vlb75q/P8NU
0n1kW+BbpnpfqP0u+HrgCAFwhcCUmVbqnGnFyLnoQzQDJrF9a0AcmleNEyHq
OHWE4+J/k3z8/hcF7WKF87NWHgSZ/tYrRcsiJ0ZricIwTRg3iysc0xpa/S8u
1u8h/oNkksEASP1FvK5vqPrlvrNLXcZIt0YL8yuU3/1arbQr/IkBa10QXzlb
gJiZ0JnfLKDVxf+wgNvH1Mq50Iy/0Rph8FjZkeaJFzLd/kf4BiZNuyjyhH1A
wykLsb+aMl3wD8YsuiPDFdF75Obe0KRFr1Bxg3sVdUfa0yUvmqNclz1bbRhj
wmwql9UrXxPh6p+gp1VZNcJgAniKx/c+e1SUNdBus6Wz7omezFEhXmjrWy0S
Te6BqG2sCDJ+3Due48BiycYEWdObZ1+YW7MeUzxFnbRXvBO1X9qAaT3FTjNL
jLE3qQ/56z/Yc+Ux+izLdVk7yp6tEwpJqP9jTeQuxDqKdXza8BZq0YWX48o8
sd9v2w6m2l7kWKx9cc9f6jUtGWDVWdSa9+N58tz9eCnbIMWhTwluvjT+bFD9
3uCLFgw3ces0hQIMuQvhe5n26TOlXHwoQJ+94Do2QqmwtLTQVPdwa6s8M9P2
2OC5GGTna0uepuKVuEGhS7IRIKAJ4d++jefxDVwkBLbiTs3QVM7+OzvI3EaJ
ave9ucdy6IozCZJx6OLExOlwQ065ML6VarpJn8Tvn8HJ777bcYb8NuKO52Tz
87McnRD4gsqD/4HcieB33CJI2CG8y0BTqGa1wXl8sJmqDRahPFjlFLoT4Bia
svu/ZCRuTaRuvkmWlgnkDvLUEdrufUPi2fYCZjPsfmCNyf0ft3qZ8ne7DIeO
FpPzEcb9Og2P9z7H1QpuKsxjdUM2hl3OFdtMFjZ+TOqNAaZCNu1jIsAwnYGN
TxWx8Y/5kR5asvHL0G7q95wSo596khgmPjoA/aegHBS/h+h313hHFVPpEeb7
XK8ln9yIQohzyyVnQxzCqmN+5bbo7dVyXTEcIZpZPdolC+lyiTlyvUDbXtXQ
MDUF85wD2ipW+OYAhBittdgfx6Rs+JxI6B3yjJUH+gHLIoMtbjKPFycCrv23
x5zUSPb4HcrKe4NCdVEciGvUaipA130xG1xelD6IOXCcd3TJQxVeOB4LQ8ef
5aJWsRvwK9WDk/q1VQ+5aVKXKzAPXzrOI4BfZ9qkDcl1Y20Ri5b++ZUZZumz
AKpJaRK7uwzfrzPW+jSQho5GJDMfDNzAZLGNyIJK8R93YmskxudtNe7IZHSB
R6nBcPgqENx47y+Nj3meWYIyzsuxuYIu2Myq7xMG7pAU4jZ9Xs26ghdAOQ8v
25qONBYNoxT3bEHe7rHQIJNYbNy7J4EaKyl07s2mQ5hTqUCxRCFGfog1VEHC
q4VhqpKXiEcp9gq3gMQCF3hxQoE+2gulTC5VYC4kvR8UOJ7ThSnraqRr4jLO
5R1glZHKt+LxKPvMYhPIR4p7V4IMJylqJQ+0BEUBzSPKPhKAwW2K6GVmsyoS
R/fyenrWcrLgGO681C7Gy9o/J7BjtnmYEiPpNqhZXn/4o/hcbbpWNItvGDJZ
P2PLV9zqCVePd0P3w2B2nhClSxlbDH778CSmU5ofeY06BlYWNQxmRC2yMnW9
F0Bd/EhEyhjvINufqWeO+OiHF9JmLeiO7AMtjQpewcxNbdbU0LMWLJnbAjlJ
BdJltEX0x2b1Q84fXOMFC4+WJ7zRu8yMEbjROctzDV17c0bb2Z0ALmtDSBo8
R0TmItb8Fp0M3VYZrXLhmsPOVplqKFoJ6yn9CrlpePoo5m+iUZtui1RNTPpx
N0S7Q78Pdiir0nVEIPK+bzo/8p46WXADBvxREfj/AohEnrcBuWV8ZWE3gJvF
GtymWkXZicRZ8mek9DC2suUVh/8orBRlbYM1FWAUYqPOUbVTketJlG0DmWEi
0bcKR3vb1b4ylmewjcAPN9OZF6hhOzEgavRXcTXy8ZP2marqKBiV+k8zvqqY
kKPDdrslCfcbadwp8wCx4nKkEOmwU6DLMX0zARzfCFNcgYFXIQ/zPuzLSxqB
bkhP8m1+iGj7W2KW7Xg4joVg8RalYURdKHLjC46AjbiEwi59mTQXzMH4F2dW
BTIHkkDDMneODZjBy+ucZ72pAq3pS7ThNc/WAlWGczytyWHg4ssCgXLUW99m
Im8uBHP78E2GNgtWKpv2aaPnzurezb5GDENUMMYd5dKUBMgyLFGuN2zNngKn
TZ9XSusGfnNDPQkSxE8PSlERLflsGRSC2ENh/ePn5ij5w4Mf5xxtxieaJ7xg
oIHsk7ayE09wA2oZnPBXbqG0d/mTCtXpDsx3EKdp+rchG5csew23lixlxoF3
g/kn7OuqOFygqdVrHk+Sdkv+YKV/OFWMP1tKeX1kT5eABAuM+LGZzLy2Lnga
G8ha9Bac9t/4R4Gof9cf8Rb142AsfhwGOuBwmkYgv3lSSJjk9fbBfbsCa8PY
5hjr9Lm8o5uUpL0O0bzJ90h0dPkKGPT6N0oiypNHWe+bucQI1fklcORktOms
U3+4dovw4DB8dFMY9xRAHIzYoT0JJw8m/p7YG1+VdKPDtg+Fv+RxpBQO/Z4X
fUmEU3Kx+k5njkl2W5Lld86iIauUSF6SLwf+wNvOBRyFKLEncxYCP5U+4KI0
YOQDKmyGeaKG09on2bM6FGTKFolZgfvcoJV+fbhQsAO4doRUsJpFhWiMvqsw
QPHDgU8RJB3rh5gPJ+amad0Pu/ROZR6jKFASICQIbMf6sAAnS3X9Dc9g1kE9
5dDcU1dWDlq8MTNwpd9vY/7LW1h0Ajc1JnJNDu2JAjZ93126ToH1HwF7F8/e
fZRurrLPv2cc93VH/MtfAh9YHqi2KV4QNJWUMt55YcSMrsjKsCZv3HF5T7+3
rDU+ZcN9JuTelTXdk1ub5E7+E86MLngzBhgnAWjgHVWQoep3kNLXpiTBfznG
OKK2XROZyFyd0hZHT1qZEUr4Gb5TEr/xYZ3NF+BbgjXK/xU/hdtXnCArb4oE
tEF5ZzGrBFIK4ImJtPYDA4vqg/liAQ7Lx3RY5CLRlCSoz3lzbaEBG7Kw+HEy
IwwTdodOiil4lyylxGPDt6HDyG99VzIWcmH0+YALUePL1amoyrF8f2JpH8Qf
y9OrV21fpjAVKZfgpdBue7oCAWnWVBKzVCI+TcOim7mTZ2okdBSgiBWnYLDm
8FFE1SFucQotitEmxVEOWWGqWWHMvTIIchdEKqDgyZvl5OQ4EfYwAUZd9qVF
IxJCVA0XHNguIbb1mFBdTzgyjYomJmTNNAOM07lsW/3tZG1yhZ2w5h831zHE
XOjRPQnn0Yn8vHeROPa+0TeThLepFb6qFHYenzPKs2tZW8o2HYnFQ2iudaFA
Ca34m41yrOJJrm7maSKGDw==

`pragma protect end_protected
