// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Ww1cpQLDese77WkzKK40Hf77vmgcy3rJARY+ib4fDZVf7ZIWOGJs7noEQhao
YunaiOc1L39g9SFsUuWFs7+suGYv1hGyub75RiRZ6lCWlIy8MIPbNURBCV3y
YumCf3D218QqTaCWG1cqo/OWp3J/wMS7Gl0EJ77FheCJmqaMsTy3X58FU+3n
V1YRmT3ocqboiCM71PBi+sxE2NtdJpqEjwCUTIKV0Z+heEGqe5hwyLTTfexK
1wxBq+LhBiaL4avE45AFCDOcDQd7QNq3+Kza6NSyzFY/qkMWvqXEnz0cqzWG
dgj4RCxDsfEGQLqoBqPj4M2gY3HPkBZfMuS2RzOT8w==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
A8EfHsPsYgqzYuL9k0ai18UV1Zfw0w/Ri1s60LY93yThfmpI+DtImPjNBrdN
gKsBGvRfCwEXr9IQGUU66R+P76BCH4EmuDj1lYNUrWUDElVuHDXYFTzZTBlq
sxVMAhdwf2RYwxXRk6xNbObPxEZaR2ikp13IYQzlVafn1wD4W8Ei/bv11UE1
lwJiBrX/AV4uXerLvw2ymo7j4xySuHI2SKkn9sovUIk3ufvuR7Ldc5/sHGFq
NoCvl5NqyL5qmYkI2V858cUiHP2weEz4It+7QG6Vdsmz+B0XMkr/X9qQ/9yR
C1YIQY2sVpPshXk/PY4fUt1eyYlWjYXLpQOgDaVG8g==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pTcZNx6nWZvsODhXRUakingpd3+BVTyd0UqxXFQn+STD+/Gr3rGO7uCR5s7i
1NApv0RHixsmEr8tg6Rk1Ti2EVK8aPDKCXNQZIrqvbn6FBvnDbfotkqy5T2m
T8qr5YiIYh4clEtlxcweqkLajjWtR934VLfVsHwH+dYIvixHIuNj2pWDPNdG
8/r0vsyBeFoEyrpPsY5b4XIa3NjHSZGSlNIssFE7S7d+XQD+JbdIEwssRUQq
cju0k1WQTijAuGbHZIfMHqRKwmUJx+vHBhVzrDAeoJfLIjLcAOKqvseOVdtY
3u8xYs/bHZ/0hBy9WeVBPAVebu9vN2LqZONOspjwxg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
M9+AYCiEG2lrKAHhm/SWVABfUc/bmS503uRCicijuFTJ6u7vnHPp9aietHSe
jEz9F13qMXkPI4RPT4w/GDTyPg5MmHebef2dJvPjgg6Iy6fuA89OhHYhjytS
xPgJySTPskF/WYi3fY03E7XAuVqpd1kGRqZ1uGUc5IjyFSUT2IY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
EbD5j0dUFwyjb/lPejc9yJa7c7rjEYHa+Be/eVt1L3F7hdUnhoVSc61Ulqgh
Z6Msmy/AD+2RMaz5wT3HmYcLTh+BKpvqGQjQLCVoYZQY2zBdxAuSlkRkMr/p
dq+ys2FY0Ia3d1vjthkuFZfD9eIPNNym4yHTUXXrDyul66tL+AKkr80twi3X
JNcwBmMJaxEQOODerI97cqkqByeNBffhgmIiEm7NY4uUJ4p7KJV19A9299M2
m83gkpxuRrZgDN7EpbBYQXSGCjbX+jxnnX1wx2biomQhqDVBDCS2mN/GbSjD
fXbJeFmzkla5yJFvs8HPJm9q1Zql2hkl8IGt3VJdZRsSNJq17epy8S3NqV26
JCYlVRgwLZ96gBFFvCEL0JVoBnjvIOrLHuFtwt8Ttyts3Ippupq+9rQxGLNi
mpqa3sVrKGjHr0p3/dppP9BRQjViBPxhwZqucdJ0UXkIpLmBQI+hff7C90Qn
smQkXq/B2BWrJ+OBGPWgQXszWw4tfXqH


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
EHvOwhMLak92AYOjLnm9pu2k7DkTwrBVummFKX76TCkT0Zr/23ChuVM14Tw/
0b6+LRIngluM1lWfJ5A6XFqct/uzNYjSonXyXcs5+ZoQfq5KGUUNpaQ7TJ12
7k1gUROAlHOrTfH6i5kahCD2kU3bQT7bYBE9kDqpDq0Hax66ReM=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Jmq86gYJxu1t2yQQsLsrJVTHkQxwbEi/SIFKavP0+sx978Yjb97VfjUaixVD
wPpFo69e+YKkAFcqtWzjfgdTGQ0U5vwdOPipSv2qg8WpoXz/FCj7DvalSt5n
WRcn3jeu7lO+hiKlhDsKaorTeW+at4CkeH3FRxe4g6xY0/0ZlfE=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 2064)
`pragma protect data_block
T38SxlKFC8xlVNMdOCwW2ffqu6w6VVEMQwKlNujycLmlwqUFP0/+YvlSWwT9
2gfsXNerdZIFLIE4bIaO2jSdVs2+bENYZkSscjqJIeD9+tq0oqBEuVBrNucu
mGhI1qyHj/clydLRvCA1tl+s1yqQrjyLdv51wOAplzEG0LWPs9/pVWFJ8cw7
7lsz57wQyxqnI84ms3D/B1vAxqqKyDYcyUy0I97Ou/k5OtuCLPY4+KSkCIdD
zQJy1Z01kysvYKBqQg9y7GxGX4hFjCqbsJfT8L68EM67M+ozRSIxsZLZDvfu
G8mMCfIPh+8Aohe3Tmtgz0U8nLZy2iculJQg1Ck9IqcQBQIEmVHvvuzVhXOQ
+VQQ+W0ZDmQzVgstkR5YzjVPto2OPEuDHbAX5Vz1Ud7yZLxSH8oDITWmRl1E
69Hpnh1WotXocsapupD+oIAvSC2GkAlNfAISNt3Rlzkie+R6i47ddBcxPPez
HKGJObqo3yroFbxhFXm1bwZMpQcj8oHZRhL/FTXiuLsry3ILFn19S0dROmUk
2DOUM+K5mSfb6mT+zDnoYXS9aBqzByxH/LMkDH9wFuJCl/mGF8m7FZBeOQKT
/LLfnvq3h9n6B/+7L6RPKGGPt0u8B7bz7zMU6+9A2LU5ERAV3lZ784cSNqhP
v0ufikdpFqFt+BhuOdtN7o/wVwdopIBa3EH4tF3Y+kbxd9ncukkNzxUNhB4u
an9VSvAYSMBhNKsuqul7laDGkSXUYZYtoURElGv4OvQXckkRoFDS50kZxyaJ
k0g2fsRrXMmzSlI7W1jrII+FMsnwWm6k8StT7DR4wBiK16l8yEZrn1WRw0nZ
weKq3sbq6KasdpLJ2z6nsBE8tsCReCDJ+Nre7GIVeVZSjt/EeLpPvXYYdQXd
t/iUV9Q/rfaPxjnkDTSy9gKdGdQGVwdw/dOuVReJhaSV3+JQ4jHkL5LujB/e
kxzGPDL98XSxSTTqibMNgaYzXItJIKujASPvOISUgKIEQ+GU1iMHVU8XaTH6
+X40b47KR4kAh1prtwSuJPdNKLrNBZnMfqLqcvII7ODgRJzfvYmaj8M+OwZH
iefUoT9OLNmgol4WeyxbIs8NVJV5gvDgYSAS55z2ALagNDNbmAA94BdeSHVj
EYS/Xd8gNjE6Mrte8rvqTHUpAV2bhLWoNCxB7CTUtCt/QMrx2ywLz7WMK0a0
0eOirhAGugWzIzZqnaYWholKTzBLH2qyumRDPNLijvRgNmDuyX3GSuhmQWvE
Lohg4svradqEen7k8IJsSbz77TfronTKCDePhRNVcAZpEabUiX+jIDvXN0kS
fPdlToNK2nfVtYN7jBKzLPulhPz6DDBwtpeWQE5jUuR7eysXSwUL02c7DnL8
FEjD0lzwvPX+JLggOjGOQE7u8SZC6mZqWc4oQ6aRtBA3Sa30QLMXBtRwYB6f
f/sW7S7P37ycoSMyYy5gMKHyFowlhm4VPAvV1gZkXmsyI8b2+7jsId8fGhBy
9W4ySi+7/N6mNTa5tbHa9D42mh5I9V5bpLg+4DNYQGGxT5VYRx9Zx9XZ+C4C
u9/n89i43k5iwfYRAvAJks1X8fxq93UWLXTHpAN7uoR70U8qXhUZBdHljWQ5
SCMySWx4MW6pVWmgQVtOPxc/DHJ0AZuC9bB0kuyPnXm4tIoNdiVdBuWvCg0p
t3uxFSfyuldjfYCBDa5JznQfP/GI850c/dAgJvWODrAk30b6Vpvu+zHFu2YB
r74o8RdN0kdRQ50lBw/J//6m26g+A6/S7h/VT1xLxNdZl+jbA1r1HSdPqGew
n/1xMBeewC7r2hmf0NUfTM1uimIg4TtB0TptjnBJQP1DqPHkVZosk/dDEWah
SKvRwHGvrbV43uXTWuSG/w9aKWGhC1M5N/NpJF00ByZC9EhTwpncvKYrISwO
XwHiGrxKczvGwmIXk4NjoqoNRFFqAuFQGFc9rV9xu3SltpSyCTpu8XvefFg3
vNgCf6PQMw2TxYbT9IufG9XCg3IOcKFib2bJ2Ch0xI2C3xxJKNOZ95jcH2Y4
MSHDbDWRPkq9KMus7NHpqMmxtj4DY4ndjzpE/P9j9FOL6AsQjIH8XTYJOoPm
Qv0BXrrgVO6A4G0plZijsQfVV2PVhgb9nqVzL5xPcCDiRIJsr0Q+9lgw479P
gaoQb+2KeV/nINyJSoW6PPs6Gbo+SFtdAAtOGwDBL+DNkVROtFwaIRHXaC7y
1JgGww930kIqFUxMk5aFlTQz/IBWHzWwT5PeBnnj7kjNKY2Fku7e6AkbVJzw
lclB5LZSujZkuhY2ZX8FTZlc/EsleTznoIpstS/oQECku7rekOoaqz+uB22O
rGJfTJxPi7wDhtb20CNp8BdCfp/F2GEUFaHb/9ik1bOOeDsM9GfJ0s2kcxyv
E+YqPwxjO/hEHMYrNYuKwxslUO3xGMr2s/BONjWD1Gadc9GiXhG+ohM+q58X
l7NJAfAZFM6qwuKa2J5xiNfamd5N0wqfluCpjzDmsslibS+rHdkaZBuIorDu
P2ePXMDsTpWPZHRjd0OVx200LqhnyLt1gunT6A9YsnrOWlDKueq4nWRzmWyn
Ni6U7EuEc7G3NZm+gcgnvD7HgxkT420f2W/B5CRv8o9/5H3XyD+bDZI5BQvJ
jLVADC/gv0a7ajUtouYrL2OvDscRkXNVDJzgb0Mo988alz7YtCoD6DxziYVU
WQZopafqPgcDmIFeaI4kdWj+rOtdIyfmIQcnjQLczSgU/WYoIAWs

`pragma protect end_protected
