// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
qLIqLwDQQ6l1FGnz27xgjU3WxWU9oXQVLuxLPCbXl0TQR+PA63H6IbVzcmzTitFt
Pl2XIQH892b76bimrW+IcoWGDnsaVOCj0V6xO4pK3O/VIduuoGov6WkGMqPlzJ1q
4R/6bmZefmr+KkeZVjTCAsAnBhOVD6A7BzCNdsnmC5I=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 21936 )
`pragma protect data_block
6whu27jUuuiFYwvP5m6wdRHpznJKCmg0PkiJexVz0UZKMsnRq2qr09HMbp29Ka9y
n8bjtRe4E7viQsHvdfjGlZYqBrgLw1PRTizGrtobRe9FuZz19UCNkUKKvqLNh7Qt
89qRbN+Cdv5FGJualI6cAUtwg0RSs/p/+aHphH79+Yzc62X1WrekxkxlnChupUiB
fHRLaaZPUsnZINlLWOKpj62AyTplvYDH4khNPQ0DBcqF7mWzTamR8VMtxJkRW1+q
hL+dXPjZzZNhYsGGhL0I6hGD+LmtDjADcyRFH8NN0LrwJkocb9PJOxukv9A+jiTV
0M5Qvkp9JXzCUqk11mBo+NQCTiCF/OmFVw/FgZhq0VyeGq8jse3saLDgCCRd+RVh
hofhEXyZxH5KD5Dr2m8zQJ+BiQU7KWakv93Mptd9+cGT6UabvlXvAzwqs8LKE0EW
qNMPjuxq+dDi682ajXKb+oKd1IDMai/7bRGZQoN3KYCT0ivLQxZe/S3DfOkuiRI0
bDutLVxby21MekE3nJB/dJ6pc/5+G1TusgXkD+NyjjFf0rSAsntdEPkuSDz9RuSL
fPeVcU6qVeL5SHjSc9HCT09gWR3fHR9wkSfBVUtMzigGk9wr+JI5nxPRFNRJEWnY
smkPMdfzb5SqAz+VGjQc+ro/H2Y4h0pHtAQKkVGa0RThQOXYY94AfY4B6kdyMZ8b
9Jbj5ZFK+xlxAx/75rRVCOkDVLQr23iq10+xrTEYsoA2XaRzAr8FJpzjdAUZClhQ
GTesvHzJjHzW1vPb7Qgh0fsU9/CIRXUuxLqq5NdSSG+dl72D1zv4aYjuauEEvos8
9ZcoEDdS3HhbksDfnH4iBu9Yw42JBpcmGguPfp+CoNPuTExdKU37ZXDhaJmgWJnE
nPz0535ERopI9P3wDJo5Vr8jdhIBT0S4Ixd7HDhm/EbFDtvWP8+bInvljsyijbXG
wb3VKDiy2HyBrjccr0bALQ4gS1cwFwsdC/SNqZZqoGKUw4TDKX0OIkUt1K8aDeqE
15V+VSD9JREJhFE9CRbYa2VunED3kGzd96nvlJf9qNPQLCoaaNycUnCH36Z2sM3D
HoVlHGvBj8lpIHx1I/oQzdE3FGdDidoyEyXz28JqyEfmtNEC3wELnPPCiunDjZ6B
Cj2OKwxIDkfA2vS66mhezAM7o0xRq/lCaTBjKkiriPqrTlR1nvuZWJJ04DJxsK26
7EeSOQK2F0XTGdMKOeS7AUJ1qxwb8dGzF7yjLJf/XHqWhl6Z+sPg0dQp8YNEmwBZ
20fiOhTFXu8vZR06smRqpOChhrvmbrFZMMYPv8hJogs/FmXK3IQu2nkRmFOA1jW6
TmDgQTBGO21hEJRo9m+5kKACZ7de9PXTGaGMkGjNnuGFSDiNpJBmOU4fBqYcpHyB
14SeApuu+nORH1WH4ja/1pX2f6EynmJzZOdTAjoR77EsjCdXqyMZNpxeHLrLkuhA
Y7NeTLco77xs61gFFuITm8WI2uuxn8z5vyZdy65bPdDJzAs0nDVHzQAiCyv0Adn/
I0rYuCqOoqd/iMK3yqQpbFXTCYevpx1Mu0iOLU32SImiGr1oAcIqFRcz1W2DD2VQ
auIwCjKSccwP5nPW4XNJgSARHbuuvLvSmbBO9OZ2Pfg0LFfQJtZPwOrZB88eEZVC
jJK4LqOF+lCUrVLdm3NnHAOngyzUqrOR1d/XL0n6GWqsA+HHgFHLptAYMPLUTYO9
NlG3KfhYUJb6hzVwg2RKAb8g4hb9dxeDuHWBgz7L/zMSIvT0gDFvIcIs4CBtfBP+
imhlm3G96ZfKyP3zF1BU3E0HqWanCZja78qIUS3fIgt8I2MoiYyFrPNTlMEwqd0U
TF+2jQKMxwGlNbJOcelMWG41BFnH+WwMEc9FYHSB5cRD9BPEL6WQT+H0l03PnuZC
5MHOXMsDjm40RnZHYM/6QYVK2Pgbmt0qVtuQlnyuiu7Ai7lWq4vrhe+5+J7BxDLK
Y3ElD3w4gVXTUAT28pBlxMongiJE2vo4VaW3M6wLSbUbM2YxLa0QIXtiMcLXBxWv
I2oTtS9pPgkhbpMK6t1CT2Q6jySSU7MDhkS2mGs7So52F3VCs5j5v/ory/nfoMmS
E3F0cZompDjO1SUrOiGm+aiUiQ0mMucfglbQ+/SqYEuD8ZEn9WM/r9htNo+nr8Oi
6oZYZ3Y3mnfzWAxDDlh0lSs6tmF+4cGLDrpwEg+Iy/vV9qjPOQ1t0ctzlOvbcMy7
IrHlI7vD65b2OSwy1h2cOD5s4Y+T0nveYdx2J6mG+6NuyFEpCTNp/kvxb2oMaoVF
vPFjKBFb+GbYybHmFQymC7oxRy86bQ0Z4lE4pDz7Eh+AXToay8NwCY0tUnUGW2Jz
gSy2pMUHqR7Tr8oMZTCpFyHUxF6okzRJiI7UAXjmooGObIsG5If46e0IDsrZchUp
QTZ0jigK5qNwDTK70zzh20XTvV0L3HlnSTly8juxF02CZUCHLBeOzj+9cJdcIKK7
Cn86WMyr/8iXgB1GU9ajI06KtOwQCzSPwiYEeSPNlULs5NhgBMyD3QLvJM2PMicT
a0wAK0L68JEJK6v+lMZvHtY4L8ZJrBs8k66oq5/m4seVOCGJoXcyw14zxy+unRqA
0S43EaX9kSgvSsWr904UkWRrHQu8VMUN4PR9wi2QEl4yI9i47Mo6bh/5352wfEXZ
TRHRot+pp5vwTe+ZBa/2icBJ9OWh8rVeqy0mCvoCi15IDyf9ij0vBiBA75kgA2aV
vbVZMK0Op0MbLdAQrsQ8YIxdZxbUPxd6TROEjA+KBsCu1Bvzfle0YXiQv6nlgQKy
AecfgAu5mQgJK4950ubfhJpdopHQjZqkOnR5P8dpDPOr9waeOY7iTrDZ3X4Cg4+s
YOY31UYyt7Je6oxDpFpLoHBPg6GaXi6EI84uY7zjTgxpqzSHfDMufr18/ZcwZ38Q
V7BeEItHty6q09cmvLDcIZaAeng8zUxM6GlttMAd0wGi60jCm0RHgRg/FnfpSemX
TwD233PpCnPrUFHmsUkhGBdXxC3iNqPVqOu8n8zkpLgjk0xXqnlUk5YLhaR2EPK5
H67UM2odI8fvrWlED8UKdtMc1Q2Wm8Cauvj13QP1eovJAFnHwuo6lNrpsj5RokKI
9qt4l+eW6y/O8ISQF57A57hzgRNmuvN5AR/uy2JZRuRFt1i3Gf/R6HGtDBKzJjZA
Fx+HNcLdmgIP9rHqltQ2BiW8s1e+oKsaZCp8fBgA1wa34YEM+lMbe6x3btkLaXag
aBs7Q+OGsURyp422Km4SyAaqwqf1K9Ewk75tE+R7fvce83/weNBDXtUowZI8U58Y
xpqXQTKgKkax4zK4QJ2Qx32uxvvDrJ02I5SFcflazTOd7l4SdFwPH8wzd2QmBz8Z
nxH+/0fLR1VTOFIEpgTVjzQ2/IJXcqT7CWycBv+2jipRFA/wE4FKQYj+EED5Cda2
vGMmbyLgc0vZyrkp61e8Or6qVbHpLbX8Rd/5/gn/CMWAHk8rOMJsq6zjXcip1SH/
azm7HCOIBsA1Ty3VI/NBPjckF1aUIKhWR/CVfx/5+nBY4lwldzQq123yzYtUMTlZ
/yzhVdDZSR2QNRHytkkTWLSNovFxdizqTfAcAmUMB6HVZ5YWn/cDBH4j2E8rNPca
ronwgPoZOPzKWK3zsQz3X/s/bd7EaO9TG6x0NHqqixD1gbeQnK0kjiLitXl5V1zR
/6Ijt0EUrLBtipMWgpczWMBortqvvEMbDSeDfk7U8d1rzgGgVXV/FfI5CEh2kqA+
GpKUucSohiz+WDk4cDGEc/LQGjU8iDm6g4lhW2qjydulSYcHwXnbq5i/e4cBz/7C
9CszHufFEhSU8+MmvUfYQKK2Yx5BCe7lM380pgk0NBFY1jxWpdMJVC2NaziTM1ow
KVC+6Oq4dr5ewvqc1blTxRRU8YxtklRAge2qZp5JqgA71tH6Mlysckc+hf2Avx6T
LZQeTZ10+fF2f3ZL6LfHcJKwNe/fFuX8YiJZVhz8rMNs/LX8LzxiGsYMocLrUwHc
EZTKlDuLn4ANoWa5oDdRWjPgRxUcgj+6+LSijBD2Pc4Y09mRwh1XxMtLJZhi7QkA
bhjbY6cxjQC4K+7t7CrmKzv+lwUiX98+UcRsuB4gHWiB0qGjr8ukFminb06OQ4X/
0Fu/opJWu+5UOWrT5xmsZZm/D1qTRgHi3ksy6VgJg3HE5Nast70Ok5zJUOVl1LCJ
3MVx5RAyJGVosl836NpB3Sfe/DU2g+0X6uPZ2RqDNql+YUHbK2lRvEyxqHhmlusx
7NmdnbwHHdohItmOsPFgQKrZv0u5jIL7kRT+ofFX4NhRd3L0AS1M7/hmRVqggncz
AzphLvo/y2RzNaeGYIHTv9uW/uI2P2YFEDpAqIgFvMbq+dEz8iomGwUUFFb6thUg
GaBCKlCEX1lbKGuCMc2hy90fBE7BpPctPtyxrzPHTY4nRCiNomD/gWkh2S8fMXRR
UBiQauftl9tR+9d4+v67+4SnhjizTZ8KKjDM7UvRTBynFIbrh/OOrioSeWONuOAj
Xrzi9YGvV49HB2HBmlYCj8Ox5ATM3pIulPQcpBsePmKvAfyxdfpFEuhj8rlxda+o
ekGux5D2M7zNtkkmqUxDQVzDHZAMqhlWus2roymUDP1QbAtcdaIYTGjqKF1PB3lj
NZXfwbsWWvJ2xxB3/Ot76fmjB/u9g4goAP96eD6MuKRRfFLiUUWASmyiwZEJDZFZ
k2TGVm5+P1h0TbBbTOBwXItBNOFdQDXS3HF7PxEHkhE48beUmHeb795Iy3X0+Xyk
d8AtpuOwBGOkM6b3jHyuGN8ofZwlvQLBKbf2jeniTh2yiM6FvW8wjv2KeJ+kEANM
XDgSeLSg5okxJRQSpTvQnj0R4Q+Uer+8lvxQ1eMXQU1JQ68UHXYrhU2EY0MBw0ih
TzQFs4AIyS52sSNkql8rRrpOBdiYBWJ5gH+6neEM+ZPn6r+xNVO31yEa8QFT+Aj7
Mu04iEwtq6D2bzVFzoq8CmZIGn59riHhov7FO1Tqwz1HwRXYAqamungwU766oEbU
VANHZRH/HF+2EvczaQlGUgbZ+Appwl5i5h53/b2izUpW05BoWmXeSBeOAXlWTqG9
vcXWVrMoLTLTaPuQbZVuQFH0JySLbLRv3A73dPQmjqwv0MqCWzMh3bbvuqs4ZRS8
yFIKxGXX1soRzFi8iKbVAsqkC6wN6G/YzKLuR+LM0ktfGGYzkwzlFcu0Bme4rAuE
V3umNAdt4XMm6bmTlhMBqiXHIvSB/61RAOzHz/qb/yzejnPRbDG1a8G0zGIMW1uL
yCf0BMg9S9cJ9ikO+YMPf5illoeW4Ttbbd0grHjTY+ZcmXQL/OJht1qxFPzgF77y
xu1CPnjoQBN3P2/aQT92JBOk9I2S4x5YoxtOESaEOK66fvqrEev2qcsHBW6Rfcrf
VdcSkYrrl+UF9knQOKjOuDR2aV74u3B6NdXfkHT0h7wocUTf7qbCkZQQQMHPyVxZ
4ENsjNG1P4mDOxsnDK5hZQyorhMlZETiZw496ASu50CZZ5ZuuOHcbyWAyvw1AbqG
ftJjUuqHV1SyMQT3OAHVNcqCEtqI5rScts3MDKcqo0BV4WoJzKnbU2UHll329fLL
3aiR1rc2etfc1f1IMGGlxsxzwuZ+ZPBHFPL12MfZPPVnfv2Vx5YVt/wXW1iV5/zu
Xmndu42oFIbc66GDRjvGmR/4vyAJqCkX40q0ync/1VHXNzsKBAIAf06xaT15sp1K
vpWCZ0WG4yZ0/jUMg1g8u9cIFPLQlvvddgvimyKVkLVeAPtv2IX/WN5GPuiYXVVv
I69YfmyYTWO+MLGXjHQ6ewwqqwqQU/0lxRcAbofTEBrc1B64mNywefivQHgJlO/z
iNLqeO62anQ1Rs9/aiVKktPFNrU7g59zra7El35sgtNZAUL/38nJjr59YUqODcbr
y3vEG9p0myJ5XJk/7zNSwcVoLH8amR/Wnt0vLPtt3I3YTEYYXIQajFJTj3Pm+H2d
jSX5qIdszM3TNSDIdNiMuAKbzZ6J763tAq7mMHmLzriWW6IMo0ANBa9E8jGhlurh
RMNy4YNYZNeStscXdikFTenTCcEzokJlqUiJX503n7muRQwV7wGVHdtlV6hQeGYQ
72L4gNkW/csI2bNgwDLulLAeF5fGjNrxIcxuRzbJmc1Z9st12ey2zvdMbXiyATZv
M0DqhumrGOHzpDo2Zz8UrDihcXMDcOiEYr4ejzmBFQDd2EFbeL+i+IGmmmP+fG6i
i/OjgVFaD62DU7jrURB9Gno9wMWyMRPO1R13xBkgDrie4r7vzFRjkFkWaNxEgZhZ
JKnpb00yOx0JwUBmg4vTyx+u1+Zz/MMEPbHef5TaOV9L2zl19S+pgO1MP4dfgUR3
1CufZpSVm3BdSvH01Rqdmxnru90ys+fdC4rG21RsWjGAw0dH+vXjDwfWx59rhP0B
RJj68OGYNeqLksfuc0dBtfE8oeiGVQJN5R4+79cGVr0NmWW9h9wQLaUpJQCU+Dx2
Pf6irHgLuopkyrUIOAiXuQllzYVsoiCdKizdyw2ZmzyPIjiOb9zOiE5AQzJ4UOqg
qFquFVz3CX0xq/Kk0ad4Zup6FJGAkxvchgEYRshZB/xpltVEYrSH92FL2mwzrkOG
2rxRaOXlJ395rEELh8y0OG6K1KLpSOVLQwiNVCkAsSxhSSZcW7q/5wlVYmsCs1lx
uz4RyMiG29UU/Gl6X8mwLGXLKUK1Oig/oRuLs0qpEy48Gs0Erlqh/YbStuDFdnUr
f/iVDW1oCrr/RuHlnXPWbCj2IKUPHVX4a776TArLvVVnrRmC4pkopWhw18TXIj99
WJd2cn+UVMbTPolutq4eWy5dPfIMnTNeogP3LDvG2HBD/sqNFVbIumqlFNF9eSa5
Dg2JVCNGEoxUzeu6pzY8U06sHOKTNHOqL83obHOdiuPwfBVtVGFvq1rZ5E/348K3
7PJJqZeqPENdsMq5gNU/aYoJuASibsRQXT41YKZzafDBvH3rOHpVOwmsNXN61gJ3
SjFnBws0MAgeLttm1ID4cGowRKBYtxSAcX9iIE8HhnyuLRwPkLjYG02TWwnh3apF
5uqTRe1SnfEV8embtRWYTFKqorw/TWcAYpSM/OBJywIBBReU6EfdkzXEUM6dFA3d
NMmUtOa/IcgoJRIAuACqXSI2ODQIf2lLeTMtA1AztLnZPSGRHUOClNkKEHML9lCS
OfTiFoVHFf+ERv6uQDwhEFHeDRzSO4eF0zdu6f/QJOS9FJ47owuLKu+82mSx/Z55
OkqZjyK+8kDW/RtrOqd8jcWr4EVf9scyyjHhUHBRYjy9R3Fv0x8vJ+hSdPicKUGg
hJwiLDSLD5h/6tCXg9xRIhaNmeaE60ZIVT9OWcqtIhIXLhZgFRF5ubLDjImnCJuj
avi8WTnLukOCCv2twdiefXgmcFuwflSpxZ9y1tji/A90LRIrxjLYloRtEqn6+/6K
dqB6FY2OFTii5ebW3/d8h1qog5e66fBccRj9L0PrXmAkTZkOHMG9j2dHUByx5gRl
XCcWAPTzLywiVaNCYxp+KMF9eHbXj/VCUSAEYjbREnbcTC1ff5T56wPfyOzep65G
wGkoBRn6x4TXV3jCA+S9wTyLx8TtRvQJuquUncFvdjwmGpFYOrZgBzJQbpMA3tCh
s1BgA/P3cYNBR5aqSWWRGFWoqQRrDR5PXcDM7JKND9FUCCXWpXDqDEUtyWYxbgaA
0sdUf9xRpA3ez9dxgjbohW7Gi9sM7MWYAXnBtTGNBp4viX3F9U+uiuH+QSxZYXBo
8FibCRbvFHwVmaXxrQHGT+pdhBmmSP+MqtoxD8SRxlYqMInaVYePIqNhrbZRg2Lo
i4KlCyvlmuaUjKu0ZeHuqZ9a8uwkGZt2N4viLuNlCtDGx3s3UR2xeW8dy7Ewt3EA
p3Dhs2PnPFbjBtQlEmEbKanxn5aQzC0C3M8bnQ2FbDwCJcXaDPqjUAOvyf01GFxd
LlQGP5LGG/vBWs+PcEw7pFutRBjGLLikmtWVAs88UkczO5zVTpzFMRWrZhNYIoAl
YEfV56tRmDFQu3kP8orY52QK6E7IRlySe1Dise2zCAA6uxEaXgvzC0uT3thlNqNB
4C4N1PuiuXgrLtekjYr5vLGYox+6TiF/++RAkHut0KvX1ttlsyqSOw5zkDbFb1oe
Z8kfokzgSqWpduQGcVjFy8I92MjBx+nkdrdEy+nxJ5bUJlXGSIX/XJaD9WVOuMzt
ylkPPpvxLefipvmVIvwEktJ7WSNzHpXANZAh2HqjoAZws4xO8TZeqKS6IQcZ0rj7
8qyqL25sRH8kOmaeK47v9DuYdj7+nO7sFs1QARGmWL9zjJVDdcOGPWBMoIGWoO8v
tcBDBZeZzhFNp82v1UyjdVUZkaTRzg2RKCkT1p2hm7G4Er6W/OQC4lVACYt5f1F0
tu4n12u1Sf+J46ZWl47K4u+AOhwHHxAQhpSe5dC772eSsm9faxa7WxFL+pg1+RN8
bJmbnpCFvXFF13NF8/SNysX6sv+tq5I+V8u5pZEsh2eL2oCJThTtIoPMXmvJ7k74
mwmwdylh82b7sW75cNOrnfLQLXTixH6x+LG9UwMQd1aIKW5UWe8a4OhAEAS4G46Q
00oYj12cGwwYrfI6rapNNo+2ig+Z2b+gjvTQ1u/1qnMOCTABUipyEb4qRoRcNdrd
Gz70MgnE/ALZ9phhoS6F5ynS6IOdwWuoBqDWOKNe4q1QPz09V+ZJa2g7mMLARera
wDmWsjwtO4TnCbg4EJGuaAIQpmimAypXc/Z6s/pfFykA1YqC8i0ugUs2EusqpK1x
W+2nobMMvwNFXtba3faJ93ogjf3yhfB+2wg/8FpDi05JhE2SFpO8Ulqh1vZv7G+g
gGEWLJOwZRdJRg91DYEutmj2bpwDCfB0hjLd9jnq8RZq1bDpII4Xl5b4FYSd+08C
5Yy0bz/bLM7IXRWWx9YYB9lNGtBr3VzIGjtEGvG7NNm0t34N6D580rd5lYaMtqq/
tXjDl/YJC2TOWUbQTdMF5kvJzVsc3Ts/vgB3eHcAz9aVATK02XH+u7SfDTXQE+kM
JoXjGV06ZVd1qO/pYzD9BW5NS7mBfiWCsxzkLFbREmOrcoP2gk6E7wo92OLKrZ8x
waMnmZ+oQ8y+47KbDo7SmYEfnPamLb278Oea/1Zthk87tYu1JB8yOjjgG07d2K8M
k5UyTPZWq1n1QD5Wu9Z7z2cQmMLq2JU6hNmMkT+pOtREoAfBlw6k0tKIXkCMW1e7
gOxUZSKxXCLl3VzxAmuBfFOUsLZNVDVNYLjnXKs+fv+/p9b8YvfZ5qI/Q0DGixWk
lEoGl7pmDbTA3iNke3X5JeTyi7oBYrwbTMjamPtgoM5agybidzDl04sQLm6lpvan
GYnKKoDO+BLNCLIafqX23QNII3TZeUXdwgG4yu/NvkVIMXFJGu4N0SKjA1vgE+u9
E5ipgqpUYBLD/GT9IpL238kp5rIxbkZDIv/qPBfcWj8tMDpJ5ndjISZTGwdalg/r
DGGacXpyMyu0awfvciDwDsL1zIdIe4KOkTTSWXlzg0SZYYievYn4UxbZ0rhZ2IMz
2OkSe7y7M27scdieWEelS7GuK+16JVMBjXBmD85SB7ccc9q+u2c/MGlhZYqLiEuz
4wg76aR03kJs/81Gk6nnUlPjSEXafPVS/d/deyjbQlFzwBTgcHSDelLRCyuj5Bft
AVMmhbCZxnzqBhC4nUn5B+Qqb+NDPVFaWIFBxtb7J6fRbGx94Hz2iwbj5U6IPl+C
alpxV+yMGS5Gm8CDKxuLjTghdjE5MDKkaGr00pPw7UP/QuiQo3cfa+mTKIvX48ip
9aozadBXLf0BS7Ar84iHFKWoj9VgjGxy2soR2D5wPByNFCKFREdqcLIOeJWJRADY
CPMlTPZKSbtdaHUVNcXmC+KcL0gliyc/bfQnvgTR40L7OtdTsWT7mq5IJBmNQQU8
O41Gl7+W2i1CIbn062gu3Wj1YaPFF9BV+sAeie3dVoX37ePAtl3bWKkYWclr7oLk
ilvEneIaW5djGQ96OD6lFGTEP0yQzm3IA5D1H6k6ZWMNcI/f6vfRYzzOKcyjdz0c
xTXiCW+8OUHqmKNuQm5pFwS2+8tYa4L/HGkXrw2qUHK29GyF8SekIZzZ0c06yBo9
6xLOSFc/5QWVAkudcMwOTZeDFqnqlW1cP4KuLzQAPCdkzT676Ap+bpNxZ7Sy+I15
GH9Xh4fW0V+b54enkr4v66PAc0e37DQUB/lpPzzuaYbKhYjm09pHxUHJOZSYc6lg
qoqzvzuIqqM5sGMUnzq4voraEO6v9ppgp3b0L67Q0lswkCG5ep+QQeWJP21as9SW
wlCgXG1UnWFO3mBJ27uObvaUehhStBY6Wl+YqUAozVNlX3oJmXtx/mR+f3Jrm4HD
2wyiUKn7cYTc9QWmulWNA60yIYKSHDL6uTrf/WG4fLNt8wqdyOYuZd8IlEvNe1Dx
Js8SpbRr+6uA17NSZaBCnCE/qBI6TG3htwpoG/TYu4gsecePJWaMG1SHBp+FhIoA
5f4aib1glLOEwycnWMWn73fGqC44s2f3hBQTSLGlF1yKx6raJ2c7Ca9ZrvHAzDh0
Sx0fl+RBzgJbuKWlV/BUeohtWnDv5JOIjoGt2LbQtRYXIh+lAHk2u2b7irlp1rG1
Wl7xQIwiG/Ry5Ta441nf+HzaG/U1cQpQ71Ebv8UDXDJrXFk1pABSIUns0tGrtjCh
d7xYo8lNcwwn2up0vVb7Xuveu+fUH2liWVATnbANsZ9f2lYjIkuhsEAO73NIAPgr
ydd8M5IhIVqFoifLux/jl+fMX7mgn7D2xMY5FonMBLfTOp0BOnJlJDi6AXFUiE6O
Pi5V0YMhMvSC9pXRV4QynmeALHDFvN0vq8FWn+4JrsutPHL1eXJy2ZvTjcpOM/u0
u+vEaySN6J7/ze9H9AvtXMzizDmRNsmVtl+MMJOLKHErzhK44iEBzmVS267dvm1y
PczQVi0uFx0CvzMdxx/Po8bGHtXlAyvtRKzWyEUipt1HqVaT/mPO5z996hHpVS5d
MKout0rG8XS60PfQHHOWGvtF7dw7nGYrPMw7KaDKbR5DwmoHqHzhToe+A5BKd2+8
SptAjGuaBJLCD/hJcVWQ3EIEedGwaSXEYbMLhYhFR5VtV/DUHR7xVXjLZeAI/Lrz
AWY/WIV9bN0PqMlbL4n96IxsNZWMZeRLm0lU9DbpijwAgiFMpUQ/179bM6TNbEyp
9pScBo24Q+fEb943dXH7QjFkB8ld6MQOHPF9aRlesZMnkDHYdGl36OUkxKSqNFIB
dglJUaUxUfaE/kVT2AIUA9NuN9Noay6gygivoQ4j+C0jHM44HcrDrDlZwaYdQlNU
34akQMIWtRE7iC/IpgQj97ZKC6z2TDxs0WqmE7xLgoIVJknK0w2YG5Y4rhHI050v
ngy5eYCxoF/8n/Xk+fzWol+lJfRT0R4K69hSPw99h5vESlnzXOYp+9/o6ErHnmJs
PBOcqlR+qnlEnoGo/FLYc1x+ElBJlNVC4867r0bKHkSfAMlFNCDrD/YSBad9cooU
JDHrqXhwgN+3wQL/AmrITp/m0GB8lARLRAAzCRzIHpf2+Bc9SD5XA2YVEXlW5JTl
M5FgKJ0ikdT9p4e8vXBKhO9rrcnvueDfst/eXlBWxzWoocWqVrlamRCHrHTG4rig
o0RM0EyjN1WxsynGT925p6LQBwbcJKWo2iCDNd1/AaFZsWyci3O8IotCYSxhWeEe
8zTIq9NT3AV7xBwgGfGIzpWL/huDmGiCh75GbmhzC+G4QCyOvcar7pqZUUta3zuQ
1YvOdgJJnfnEm02e1YOxwtdKkYJc0FZwrz6KLuSz33AjfGFULI9D3TVpEQTgjtD8
cYXN90n25h6Y8HzdE4NdIdEzQMoRm8tLvRqP7AbOK/ydLwaVUigGD6K0gZxtMJi7
fF0/YY2MxV1rhYymCnvw6MCaBej74zYSq5Lc7HI9nzBg9EjUm27vPilSAC5Rs29V
xtjz0QWdHpRQdTdz3edodEG5bN/GYjJmB97/PWvp0soDquYQ9fejQ/oXio4dWCWW
LxseyoqazHlybo0CN6roIIuPxhZFfjxgOhPnKM3NZmmk7e4lcLZt6YSS2kYt1ibD
IBCRhOj3OyncJv6WNj4gIJVMC99nbz3PLOvS3dAKeHUdDTzcLKNue99Dp6rhWGTD
Dligu2dTx65QwNxugPsEJVXExcwDIDRpR9I+0Yohk8tMnlGJnqMPy1JfSGcNewRj
NprGPbIdvvyHD2m2WUUYXJYDrVKkBx4lnnfpAizB//qP2QhOB3JR92RCp0SbvRMn
iH/+sp6RBxGmv/46Qf6rpZlMPOkk9WZTUEeWz23gLruIYApEhoPfpC+yPGms8T8n
H0GjxdLkLagNKhYIhRw4hhf0Bjh4d6X1a5Z39UgaLkaAuTh2a+W7YrfVKma/Yiqm
5/1sDa+M2uOqe92W2ZMZJOr0tPsdCvQlC+A+izRXoG9vDDTLzw1YIBBGpK6+fxmK
fUdFx79DHB4qHJiqYRBpPh8Mxso2hgXJUOnaYpxFAsyysTAGWJ51WjbRnZsBG559
ntzjX7cmMii1Aave4pAnYD82cdSDU2hDo+xdbRNMemvlFhNH+UNdymrCXNgS1tyo
nevxWdCDq803i4PxFt4/PmaJ4GFcuBNVteNAC0eFbUh0HntupqMqFQjhw4seCfx8
WxvjahSf/Ow1uoNrhfPobEYZydB3920WvNo0kNkImHMKyAKsp8g1mpnZtmR2LgG0
ZdEYISdMVQ0y8aDdg0KaXb6IktzzGQBVBwtzEWQPC688C59q0ZzZcceB7TUSSYLW
+rvmZ0ZGuzx9/TD9FdHMwR97F16rx6ryYG7/JFTG6maQXVmnz34/A4z6zwBYLk10
UoC3HXvfePxetdZEClKEuvZrrvO9HaLl11zRP+lSNShzGYyaSmhf1Ut3qfpKsduO
qt3Az28iy+lTymDprw7rVihUGRtgFPCLz3/Pvdsv4Ak3/dU40V7QYdiiZEcbsIsE
BcLhqreWMmpomDdTJEf/KxwrRuk8VHnbzVrt4OJDxmc6O0Wfj+3q7S091iJQwTuc
gnjZnj3XYi+rxuUry37SvF2KbTiBwdDE16XtMAPLZCwNyK3ynRFEMu6bLlaKfyY+
gB3yqoyhcTwqwUE0iQjNu47s3DOAN52Z+Moj6lQD8sR1fXDGchZ1XxQrBsEqI/vM
cJpj4ddf4mt6eeKrzrxud+aDAgnWP3VRBQU/vXutnqXmZSKnAV9tznaNDEfpCgQr
HpjqENehkdDG3u7orNavuaNhtoH6JWjRfi3pj+Jd6zyhqgSDG3BTYG/xTvJ/oUSY
IX5C5TT4PVUnjAcRBfup8Mx3y2PB8tp1dln16cVoMerWRktFQ7iTh6Gi8I8yULw4
VBOjirEI/AeqdGKxNEepZCUBF+Nb2URRhXkHQxbvJ39YiL0HlHHLPHFQYR5o3EjI
fj+pgsWFrWYY6u9yu2nkGy7Jqx2MYWwxwY4i3ww0HQgK4owJ0a9vCOSeieyS4lqP
/W/0jDPVsFOMeOmJ6651vIImfnsbHFKT5Bkz1NrOVXxRuRix2IiiBP0qbwTALzZj
nQLZrR3TIuyhveAKYXW+NvSAlpUIbNDSp6fmgV0ZF4ilEo/PUtgPpagRKut296RO
3HgiFbD2ZEJpVr+WI/sh6qmgJHxD/jEFGA9EE913nYoVTVbNQghp35AAD6+gkOcy
+1POD9PDX6gUpSsKJO0T13/fS7NKxv0hJx3mHHwQnuI5hqvPUfU35DLZ+MqPZeG0
G3kHXh+RHYN5k8MUAFH9DlmWgjWD7dE3iQQLBUTMxQqbPakF3xbnh6kBDD8yz83W
cduk3nYj4+k+9WHHi6q5oi8LuKUCc7/sSNCphrZ0sv6waM1H4rIU/8aTOmsUS2Yx
NI11j5kIy5apRJmznteHnjRgOvPrMHOvnU5XwNhOzJB4WGVs7l9AxwDXYHiNrPPw
NeOI+bsEY33df1h8PSvDebmPXN4ruZoa0aLFmWjRQ2aQg5DGgs3T3jWOSzEY/XJN
nxf1UOARiIg5bzRi8XbhhR89w0ONEMpSo3TTN/wPIwSEdFF8orEOiNh9zJ4DAUTZ
VgD/N/hDusTH4PCyXeb1CET7d6SHiMXG5Bf1vdJtFIIASv2HvVeESoHOG6hAPlMK
vnwzua49Boz4/HcXFG+/30APr2EzD9pFXW6SnZx0Bma/pTL1RZnAOlKXk6F67mf0
s1+0Faw8XDcVSRFC00gvavI5R96Zxi66kuf8eQ6asU8SR3CYf+ZMyurZofVxVzyM
NZMkjE8pVEc75QwhQc9oAWpKCRckPYxRK/rK7sbCFhV4G3qHk/C6lUuPfKH3/9hw
vQnt2f9Kmz5GIfH0JvV4XE894ZNZjrg5exRWqf9vZt4xzC4AvCfPplF7Vp0oxySv
/L+izssMNdgXRNMe9NcxztDBoWph8JqU3+rgkVy3zXVAl92bxCETW+4rLiQs4PYC
++n9gsNc3+u1WvUb5ifYXyDMobgBnf42tvgYzUt7LgWJ/ZX9vmlnL/A+6EwKzItR
4ctWo+AHFxjTxiDQYys/Dl/5K39nbKyqS4Uu+cpTjn3Yqv6CE6ONhzJwRkY9d9Va
HaEY3/uD9Z98QbpfrLmuKY/qmu9X8fb1nPTRgkltMJOfLWZJgMlPFB6PrjPTJoU7
nhbmXNi01nbsRq9M0X33OStUEDPinSHq2G5X1IulrY8TqE0W3EuAdwgy2TvNyxk3
RNu4GcafQ/V/98Mqj0hOkHAxjPZbSbNQcAXldwtd9wBc8X1vzemaApUV/pvpK+qi
cuVdmcNnSdPKZEsDDIHw13c3KeMDwnQmF2w00uGDAvAqSNqSHUWAm+cd3uxlNo27
pFTGGA6PBsr5BOOYpCr5IopBpOxANij0rWWdxQRJoTE0UJLU2Evj6KpbYQyxrVl0
vZEcer6/kXV73nJsKUrmSScyvE4AVLKEGhzgUYUgfR23mZapmrolJTeRI9RSZZ9Z
Wyg/PQJpqbe0wK1d399EiMwM9hV84HYR7UJaVIPU0UQkx4XlCSBRlfa4W+VvqloW
Ux0ACCzt6B0fieiKN2W4QcjOjvsHYngcd3AViaDCNS3qDaQaO5zCELCW2jUo7ix0
LQ1D1wEdbRszWoRRItXFHlYkrr1iT0KfC+mgob5bvZMaTme+0ZhvrrO1kbsNBW7Y
PRyyGdBELPQyM7AfOjfNNIIJ3nan1xrX9ogJMYXdVbNfmo4VSbdC7g14lOQU7qEm
kByaYsR4ghvidLSERiB1Em2GyzNJhCbkCUgBjP3mivzpSgUDh23OQ6lsiyvSM/Yj
0L9V2GbJ+4Yv09uSjzfHIS5ad165FGVYWwd1MYOl3vJKfBKhLjhj5d7aJnXDJ+Xq
F0IS1rZ2tnSNo1GhNL657XQ9sTc2s68BkiSmX8H8yT36FlkYKCXCRWsA4t7rHvqi
Y/738WBIo6rleDY24Rvn9ZSTOcaCCH95a1sQTHmDDshxxgbFOzqLcspNk5pqQtA1
jthO6qWhcE7RoIrh8lrX3O7IbWyrr8tDqLzjAL7h2Jg+bmEBNLAdOjQNkj2kZV5l
KyYWQ49Ru0Dwda7ESfyZHlHYnzrAWuyQyD5rQPKh2CispRHk4jD7steRKJzHAFTX
/DXkaV2OYamn+PlHBCcNbgy+QeSjOnd6fxhDMSkmcsXybQA+X4ThAmup65Bbqz2r
A+LmGoA/4wu7J01/lbSClzD23h80vqLOYIn73hVmKx4BrW9okPaXFPCHlGfujcKs
xCrC31OYRuToB/RRdJ2ag2ERmr08eGTUvrlpZZs96fPwJlwRrAmJEceoWj04Ow4x
r3vZ++pCw/atk8WProYURL+P1Znb4afsdfdecvZMd3OZCyklustGRBxt+EG/HFiZ
jUIyNWvxiXysTy35uK9XJS9/jF9toaipLXF8iRzwMWJm4UsgwTi4yACAi1k/+Cak
uoN+WDr5wn8OwfprwkUFjD+bTm2yXdtXyro7VYZ2wc3lJlJxm6ReIUz80EwwYyhS
CnNtQhnBjmWf90/ZoUuiI094VlgF88oyi/cK2LD7uhnHpv9cWfyNX3aw77MVk02v
6NfI5KXJnnlgW62jssMrA97X9JnVphEBS6iJlPghhW9d7d+NCGKFqCFrB4VlVmH5
dFRrm7gVv/0gSiJ+Ky2wQhoHtNRQtSM4+0CYjPJeL27D4jQ5vXjm330Bean2/pVr
FzB9tfl2mmC6oYjdFEqScH7HeDYcU2QZ0TgftJwXZ/W1olXVoKh232ivYSVn7XDQ
LQmamsUfYBrpe7b9OSksusg8ALK/Lz31AtkcWPH0uqyYIssJ8kAwAJ3yR5CBvs7s
/5aqjtvVJ18BXRbciOxPmdrUEiF2vw37pffEthN2YmfJb8/o7iEBeuuFG82m529U
Wpj7BYOFU0Dy9NjHA4ntewn/E0y82GIxUB7vLuX/Rsb9GbhHkuEFMOTFqkE1WIGO
xoqO3DYG99JqRimPc2XJjAeyM3/bFP7Jk7Dg5SIFThKEPbbVeMvolISyb5Xtr4Gi
6Ode8MbFfsRFYktLSbc5J6KD/Zker4S/hmQLk/zBtkDaSlSUWsUmtckJmZ6tCvuS
fbfb/TU6LThLr/mHD43yc7cq15dbNrxjma4IZbTriz+DqOJegj6nwD4d/QU7c2ZA
5Bpltk1F5SW0/XSNvPRptIzeCajjZJZwqYQCVhtQkskl8q9o40fZyejLwaqcXWrQ
Lg5FSQWQ0FAAvv2crHotWNvhggSfumhAXcC2JtS+98TMsXbZx4Of5PMxuP16kgll
loAobZKe3kXdb05zBDKBDYsa8HlWrYfLBsb/dXomqTbfIatm+yCcmBiWMnpqMjdz
svWox7ER8Ad72Y4nUeekq8kcTicUAEUVLD64FduxSC15sMw4nbJe+SgVhpiHJMat
uH6FJEZy957SZ/aoGfQIom1/ZyHFldwQqQX9SJYrHdq84BDXqYKQCHnQqttLXWgL
rdd+9M2wTHmnFk6Pnjljd5XgVseEg4j0lf+lkxtkYcHHmPaU57ZC5BK4ST3t5UnE
SiEXqaR0n2cFFnCm34v+cIG/Uk8tcOGg1xfqQldM98s4Z5fFdjZjWB9IG3+ErUFW
iXo5Qfw0XhCk357cWQ5XbRRJy7caaeB2A5dnkaKKx1c7i2cgfum74Sq8bIjBtLil
qqsqlJcdZC/btWyQL9UQAJ9ko+eg/ZzdjBhb2oTItYFuUMvnk4Lx43uDq0OnGisU
li66R9hW8QWTYp8nUTRDtMUGtYL6klRMDQX8ywGs7uqxJ3RG5t9zkZWMTmrH2jVI
sVD1cDpgr2tDyk70OkbSZqd/VN3xKrh8AdKcY3fR91NRjvTs/A+iiRuI93ijB7QP
QT7tDJUQfLy7KNnoAJcAm+G2P81/B7i9Ysylk3AAgntgzV+hsGW67hTAbDWjs5i+
hRDseCc5995oJV6SPB/zSzas5qGMQT17o4S0gBFWLBO9tA5l1zmj9P41xSSQ/OJP
HzwYx5PHcr5GV4DavESjuxei5F9s3JSZrRVi28jufNzlh0fwHX8tqiyvHtD/xMwg
dcG6AZBSXET2undNEuzEu2aimGkhafp1+315ud1NWuuUvI2cl5rdteKElgHKCrTO
0rVrcKMk3bORYISWwxBDblH+Vtyf0ypMpCqkHvvshOSLWJr2X7Ucdp2myvFv3WSc
D7cUuwdgviJ3G+Ple1Ddoz/rx4uGx+Er4mZWnfzHan7nfIhafVaTEBMWIytqoVH0
rTRUvk2bHbUDl4Rrob9a/Vo+ao7ANjiOTO+jwwTb2UKUvbW4rJohtbsujfeDZeX9
Tt0y0ximlfZgsFWfK9bcD+0FEvGN3WSfHXOTh7E9KHwrRz7pmR8wyk2T2D+DrRb2
O5bEuEKLrSibqycMU2JStGxbhR1aG0WpL27ZFc7HxfUHD77Xe/mHKBX5cRi4IO9R
9GKc8QOA0BGuTv4LWBJboUKHq9OhoXsMjX2zd9J33o48RuOArjHWK1GBDnwZF5IF
8RyxDsGR+x7+USUBIW95tUus7P3nfqhlwdKVfnxvNT+gDWDJ1W+OIb1H6qitRnJg
DUH9hfIGLTslzD0qEkFLlN40ASFdMK5yZCcyXKZ5JZ5WvOPigQJM0NKFnYolpW0a
D6sE0j+XnCPvv/FtTOYZjE5aJD36iUpvzC+6clXJSqAp2XBE0vPidVt4FKnbAn1M
We0/JpZStl9IGy0QVLI8+6UruftKOhE2ybA8SjxIcPFLppasF4rG4kl+TxK+n7/r
UrETlVR3FRqT157hoNQcccsXRMqTaqDgZdQnucCagBqksjHHTXuW4QFBKncHH1Vp
33VxJdXIYDB2MXJeDBW8vLC9kT0j/TPJjc794cPpuKIvm6QJHMOxB78sXlNH5zBH
lnrZy9+12jv980ruqR3b05f8xceSIOBUAe+Qb5Oz690sTMuMGbX+A4TaKpj+A0Li
I7RVdMKflbPLProYMc9NnC/qoRcQ4qfsOF1jYYO9eF0jir/6X1IJ7lA4ELebxvbU
X0n+HoZEf5JMTfZIf/og6Qvq76FYy9PnmxB0OXSogDDU520wSNiX15kV/aMacUq8
k6Z847AjjXKsWUZmDtRk7/kNHaj8WtvCOkXlb6OTJs351EjmMAb6te6VBolH0FwJ
Jb4uJqWFCZWYMZgly1UZwF+ko6hKBbYT84FRjOMhIYBa9BPeFmCj58RnWrlFkydU
7D2/lxPyVk9XaMAJjBS7XK6gxZDuIcFuzCbJMRzpREDDZp2W3xGSOga/1WkNqEw1
rZPRfbU7qO/7wCq5hJLIQYj1Xk4WMV0QuxAKvFx1GdNsx22jkOKuBtaWhKj56/Tj
oDbIAO738hZYvtpnrItNFrr+XzwxhuKFgvUdOkF2A5Snq6e+WpQfzrNAuCEDxpWa
J3G3ofNe/8hBRLfw5tDhOKQtNkPrlpsqnqdEc2Mj37gSluRx9Oc92OBTY0fgtLib
Wf4uxvJb9nDctITNCSopceYWI1/rqJUU4MeQ3JAGDbYIqswxSAnY0EQRCF7YjRIi
1l8a2OcwzFLbPpOkf5HwycH3Mk+EhdebnTZCDFRJibCQYbvmAoRYy1GBSnhbyBH2
OlMQoRxTcxEcBrHBbs4Rj6IxvWYdkhCIrorCbJ7jQKVmFu/pk3qsOWw28uVhC4F6
GxT4tjxwNcSaqM3+NJnOklHWKjlp6PB+MxMUYy4luG5NMG2Gefsfwclyh4BE4z5E
uaqcZEHsR7TITjOHpnLYsshLbZKUoDRfKE3vuVsMamNKKTl/eNAFZKhvyABeGJvU
q6hMjmJyyoiGdkNL/3AE8BMjb+XI3J1SFmPRKS1kMOvkrY318RJ5u1Qc7PL6VLp4
YWzozG8sMduivrq4CxuypBYRf5SaScCEyCgGh1HBVpHVO6QFq92oCDWhtDixa5nX
NXS7GBuzrHIyQwpZe1EaleUH2E2nlDdpy+MMMEIshSb3wgBLU+bloD0NDe0TrS+u
iqVJapTrIDlEYAak93hKWS74flAMa17Z+5en+45EBdp6aTiHtxQbKyzgyHSr9Xlu
mo3kNTD5EfRU9FDs/4lWonz0b+B/zYYp27QAQ3/8KdbdK+JvMlgVomy3EWB0WrXR
gb5QUXfipk70ZPJHOZdsco4sGqggBdjuiuYBLKoz2gRzQg3XQ5OnWpc8bwrP6oFb
o89w11Cx1j/jaJodvMwgZv028eGJPkxB/Nn4UCzU2pjADqSBif/KKHEXkcH+uvfB
Lht8e1OEN59f5G4Is5DHlx3PEQ7YqPRxTbzKvCt+IyJxXcHGBViMUa9gPch9umyF
Sho42HMSELFeY27C1lLEWV2d3FT+zpmfAMnGxlvl5yi5O2TZW+MpvwSR55tE1LzV
Z+svsewXk7nieX2GnECH/QAX2T8esA71qaF/27vDjfiC/01cZ+ucEUWL5clinXnH
DuB9/qMrT+48fSjYlfKlZHCHRe9zGuE87Rkt2M6bmDNbNgcy+DV5roW/vkrmYF1B
LxTSIuLR8XBEVK3XNTSKagaBhZzC8hf/2H6SP9aa0mYxqdiVnUpOG0Uy8d+MgE9P
QIK/a0JoTlw91pDGkD7uO9CzidpLYipT43LCHiLBfNKcU/lDoGHgeaNlfcB7VRVk
wdUO6M5QPm5OhJ7d2/NtK+RaOMnrFba2TDVXFZtBGpN0eZzzo5R5UOxOOpZ/+ryt
Wqp6cSkitNnWWmoPp1eGovVXEUiRxHSUTt/e7dFC2fZG1JSUlYEchpRvYDQsuUOb
u7CSd85cmcHcIE9Ob7AhAv/DD5WP7geouwSQQkHTs9CStxZI8UwaEnAmYYgl2a4h
Pv6XNjSqALYtFVR5DZyb+h3SekX8u6qWqJ6llq8xT3+GieRyVO/zPQXx8Oa48PTu
UutQVTuiGmcqbAg4pVmM1BWg2Vrx9Tdm0yBveFKquJJ4hwXhmgHJmkOFdKGTK9F7
jMS3+QULnQAUxemXHP+yZmaMEey+RDqyngAcd0sPD5JHqaTBhkKk315GxIOVgkhh
XGx7gjdsxN9rx+A4RJnIezr5UkAY5xifWxq0NncTZKlBYro14JSs3vu12XxIKa6b
6roInXSuItPOvfB2i6Mi+rruvSbTRDLVAxrt/Xsmum9L0QHauhRIme3DSmVyBByK
g0DOM0mr2bcaQcgtn6g6+qWCPDTol2dkFl7qv6DoPC0rlQInSr72cwST/NN2qVRz
L9SzAp9WABF5jQEENw6bdRqtDBtUAEk6ZZ7qdJpgyTJPfGFYskZl1PZF17cRFylw
4cvfNbcY1WFwyA6RP05MrvbinJ09uT+381jjISYQb0xYRzu4Zbp3i+gerI94U5q6
weAzLswy3V2SH80i/dkEe6GfzTVdCnvPyPZR5v9w4vRUON/9ZEnlWoSHUeClWx3C
oWsWwgLpYltXM1BjQexK4aNqLVb8Tp6HHMR1B6/SKZfFdpIvSnLOShDjfxD6j5Ro
iFT+ETLfke+MXnWS7kn5vxlUKdjwHHTf+DulMT5Uj8BqpPuIHx8R4jqJgiIZixjo
ox98g6rrvdJlNyfje8goBG9MLiwkMN/wIULEi9qlXUGekGEJGERuvdsVBLGFcwx6
24g2ZOiRgyb/eEHrQOV8DbgD1oTmbFjb7XwR6hraDpqRB29md49xfDMpzlV/GFG6
CSiU5fbmcHWeH+Fsn/7U5rJRXS+ef/3lNmR5WFJ01cOJI+vh9sAsck3Sa6ashBTz
Q+fTZ7B5+XhEuWMg7ozmDBFFlcXpdFrTruvYpSXC8BtjgQXjV5kr2+Rxu/hAADCP
Duc7cJ+3vSFCrlkQ99ZYxsySPIbH0XYEKf5gOZcYLJ4fgF7MnXA4OYwJHx9XHh5n
QvXkYyrRw4+Hvvj6gIGhLjmNJLZCpz/f/wqNx3gVH//SBdXtAGcLYBxcjcprQ+8y
pfLztWkQ+btXXsGLyKsbxnjcCz2qpIoW2nhaIKX65TT6nasXzy+ydB7GK3W95JiY
9Om8OzrVzGskhWM5FZ6GGm/wQ7numZiv/z+IyGjTuVk9lY2u+IGfCrvyBc1UyJjR
AUF8mt1UeVQ6cILXNoj32Z0blVCbJVUJ3ZeJmLDKzw78t4LsOSDUdES5w6qY97f2
vBub6agB1d7d+TBuD6G3YrEv7UpG8lyw5BV7wp0NULLxRK24hqhfjRkh4K4Px8m+
CuPuHccBNje/Sgpoqf/B+6/8CyOw+RYyZuKoaCevGC1oh2CEYYgeWsKp0Yg+2xGM
jvUNPiAwgNeJZw7mbHH1OOj2RF34EVCe/bOZtXZ9E48oXE5pEdSzunfB4ccmIFj9
Er+fcNBDqaJmTME8x+RV53DLLz0BDY4J5eCWaVREOXvnUtkx7Odxgc7QpYNWh3/t
lfdu+cnTp0w7blTl6Er6tsdJvG4y4tsTVt67QDHo0WLxkJ417Nrq18wLJ1i64Shd
qe560mMdamamqDwWf4+lYpDYlqZwMqFEids2JoKuxxGhplLLP5jIE9QW7tfHPLA0
gsTQIuXHaS8cwkCeytE1H025crJ0NNWrKYT59Ha7KsVce8H7KGo3Z1Eyq5KvYvn9
O+L19/4xn66s3zFq6X+26DC8dLIIn4BNnRyaln/DwhnHGtE9n7W+jX2exrayQPHX
Um6xtde7VKUMcHFB1IY/0JCeXkDJEVy+IiyJL3PhrFBeFTY4pYAS4vn7yT6UAwTY
xYj9zD1apS4NJLvk4TpmfGnuo8kHNnXHyFbnfk5+eyW5WQhspmm57lOr8KK99WFX
QQ4qKf5Iye8lnCEshM92OdKPa24F71DZcdrrv9XR3JLv2pgJZQVAAr1Dhpip1xV3
WZFl7dmSP7MsTH3o6AAxTaNSpciK1278962UwsfzTgtpgSUocumtXg69xpvjPTmy
qQXx74aE4z+Bn2AuvzKDe7dxVGVjlbtcIyRRK+ciyD/UINw6Hm1aJi+S/er+L2sV
GRuVpZKVbufiV7egyi4/1yZDo8s1a8dzk5aZuJ6iHR7q6fpsUfvemD4LHa2/4Ave
ZSNzRRY/igfdTtBu4hCcoUWa19I0VKk/HB/JtUBB5GaNyyCAPe2ovVXnIa8J73zT
1/eckfw1t/iIaSVEiWReZSWjWtOrILFMQFjDFkX7OHOFbXDQ7Dg1pVCCLz6ODxGr
e2zDOKPz739ymeQ4NkLrr0b+r8bQjnoUvFHoKwksVZuj4AMMYh1OO2lSoT9ikYnZ
hxUcavJUJu/afuitevN+yMGMBXbowc7PBxyJbdzZ05pthv5EMlj2Sl4V+sc34Eop
wNQj0bid3qpCE/IdinUDXkzdJxImebkdhEpDeaAWCZA9ONxRZoyPAbe6EUAsd00p
hoayqpea+uQOn4tDcF9g+S4pjY12J0KTxz/D4wx7+wfM7vRCEpmZouWu9MSp3P7W
C/CFE5Bkv99K/oGvDEpqihyYMU7IJqn2u+4VWo7/a6y0Nnp1TRnUwVXFmnOzdF8j
Aqh0Dr43A/ObS61D0OSjP8k+upvdgca4aifynaUGsmkohzoz5ab91CEASPU//wOw
YcSf4X219dYtjEQz8PGXzMqMeWQ3uRniMwPwqsmsawZCiYLafzpBIw0yO3O9u4Ia
2mJS76bdwnOECt0tY10dD3h+og5yyNo2iACTJwkulyQI2B4JSG3XB5Ui+eVaaKEa
1uFYRIqhXg73j2RxhKD92HeA02X80/01VVXC9BqW+9Qo6LfvqerDUSEYWiuT7QnV
Gp+MvhiQRKDSCQAXV16yqlJcQParGIw0hFg3qATQ8InJNQ/lto+KWPc/ZFnwO7Xv
ccOwMzKLgf6bV1rcl7hVSIMfaAx7ZeHOtr3Na88wdpBsVjk1rh1rlfqlZMr2vhW8
sYpScguWMHonm4XU5likUxN3GTrKI9go5QsWmIALFLmbcKTEpUDgUHnx2cnpnjLa
4nWvo7LH/uGHaqZwzwz5dooLtEBeUbeLL3VxpylmQYbGNUPXLlLZStUKUjk8ld6q
fodS6LxWncTK8UI7eydRAdVGTBlMUTv3E01g47KjEUjVufysAtkZw4VwJefs84K0
Vuzf8mrNlekISc2hwWpxYuJcsMUKUuiPrKDiXVySpCHCIamBv1I+xdBYkKKXuWrr
KwFHR4lHOKfjBd6wJ1GytDGwVORD5ZFPJ+/x4AoJnvwwy2rpu12414cP/h/SiX8z
rxKsyauKdjBWtE09llY2ycTR3dIDuE5E8cMYlY7dFbk02SsUl/VnxKe6qQFWPT+e
j9QrcnlfOUxKhtwDxI5v1IZX7qRJJFxvzh+11RuTKbFsEwP3fR7jPfopUi7eIOtM
fFIQYtWGs7DxE58RYl8E1rbOzBXFRd8kFebvL0/Td9E4bAgdrGKieG2rXAqMAf5A
YKSbXipKvxQ9DcckN/jZaMZdO7kW1w1LlhvGB1prkUJUZoghQryzWIlOgLIN1N5j
yFCFhUKmdA8Mw10ZGtsGODUExU7Hhkndfl9Qa5rFWk4EVh/GjH0fltgp8QztmO2/
jlXW8AFWsVIYexyY6FLqxnxwfIsDpQyp/qyJlWBQ1fVQTkyWgBR8vxvwIhRBbG6x
8/OG/FkYPzYJuSs6cGPqgxCiY6WDqhBkqHIgm0ZM0iLnp0FTxeyb3E/mUMiBJ07O
3hy1qtTgjxapQtmxt1R8flEwwtcg7BHk1RXGDBM95eJuIKn0+gTzDZWd9QBRWkTP
nAj/F1n3mAizd4wyFlpT1oDONvbZDb+KaQE0iSI92+DHCfl9tiG8iTr8UGBPjD+O
bmTZvckQ0v/f9JTUfaa0h54SworKBraPBMIwkPjHMUzaclIXmpUkxtGzZGvOAPcm
Jqg2JGdvCQqPGaligyATWIuT8PhSxPeFI2MckKPY5Z5IKXK4KIveFKvjxfGTPNFe
ke37caG6dPhKJCTPWH/Sd6E7R/w80hWxNun6qdSDlbvzBzQktXeQwoBZjL96ipsf
zjPTHK1EMcfD75Tno71ILvP2MY8XiWA+GSEdHk9kdtVfLHq3HLgcyrD68uKt31Ny
CqSaj/mWtv2uG8iPF8pSO1ACOWqqId5d7mPI56xXV0c+qNS/2xOeYJIWWDIVFOcO
wf0ljnXxCfvMAnHZpHAJesIdeY9PmvbxJJjhMuyMvZ/a3cI+phix5xof68muv1XC
+xZeuLflQN5NccByFKfrw8R1lccSpH43rZ2NC7LVabVOzR6WgwpFeJELT9ACCluV
F/WUqcAqKXMseexxtpAU5osFfSldB+ui3Q8/SSCqejzLLlMdIu+zCQbS1+dsVIr3
2Cot1FAyG9FhHMxcAi+18AlQAf2SCuNvGc4KgdiKVGbdvl3H+/EdjlHlXW6MOWHk
rVUqF2GaayRGu/5jfukRaV6e65wge1x6FibImNRN118eb6NLWgYxzIv/8u4655OL
zSBSlO05/rhW2ZgrfzywoVHZO0oO3K3rc/rAuS577fjfEounWv2SmTdjtycWdfDC
EdtLPFK6jFar7BpmBBeU3XAf/KXsnBJ8m0Xkvctc7wZehnFdruf9xwrObf0gZibG
FmSwEbyclmOM9fR41X8Jbt9Nz2xqoPl+qoaw0xm9zGaNdRnF+dMHyJgHFDK1x5Lw
9pS3FsM1qvKWAZJbnr4/NISzcdNufBYuiAPNr7CnNV6mOlmG9fbmsWHjU+O13i2e
9jS8QkTBNtdKvMnOEhS7KFROsxnCujPFlLL5E7K2aiCebV+0ZAH17AT21w6tOTBm
nLPfuDMm2e9Dyb0hIXfOnB+mj5UuaJqsOPpikYSNoxtwSqKW79CGRiFtGI1f5rkP
4UP4BPBUyVJSBRmojdAoc0I7et4h8SIGXBpjaIcEgUcAppAJbYQdEf5o/pWWdXZa
yLkdo9bD3l1D1mpv1859vh3AK+Pt/1jW+WDwslm8Auyw8r/F/NO/kVbGnT9tjbFq
BzUb4E+byiZ7hTPNYFE9BsKXIDvH0FxrAI50qC+EV8qDbBwBQsQB0xKarhfoxD6R
DlKmn4a9yrtAe0aQggUknyZIHgAWhwPz1P2oZFmXdMShK69Zr/MXR3SAjUDHkunf
uhGC7yipJrlI0uYdWMH8A92ym7+b9X1mCpl7H7J2nOc0Nltic3XWI2Hq+5WuUcdc
ZAkWFttK2UrY1PKqiplcD2+DsUK61lvxROWP9oi7OrzxIxVpLFGJ4WqiKDZ8HAg3
RGmvVxCfCmKOr3z6FtGS1AplslISR1s9HXWeqMJb1KfuPX9EWSGWvTuXJSGMDx9Q
qe05YSj5NRg9cdaDOX2mtYyay5IrWvzIUpui7gR4jUtebFEpUxJ1zXthiHnhjUn0
ArKaevJYmbRnqxmlZ1ncL410BhKL+LxxMHD5mG2+ApHj7DTZ1rzZZJ7pvDVSxDdW
XZDbxURxjsbzW6P1C9kjjuo9J9acF6xejjgme6nZ4ugY/XqMRaCIf/uEDMdcQs6I
kAZ8EqDpVq7jERoDmthVJvUAR12CZ77ZFSkST5GsQ3kOvir9scQHuBReCwPaPDBm
sQLWN+Ovc+MLGtA7CNtfteNYnp7gEQOvThY48EPD0CLRBmJsEeF9gLlNAY+V28TZ
tu9FdaF9gXVxQ7iNKPSS8bnQFjr1AmAZfUc4xODujKz6epK3aLHlc4hScYeE2X5X
OEGqiVGN12P3jaiVBjoJ52vu1/fvQ8McLhVeNBhyMCS8iUXuutSwCBn/bskLM+E0
JqzE7Kn+9oH3hNytsesKKk9bM1iuH2fRzT5flQN98L7T3aFX9qnh/9mDsBnhgEQj
YezyFwhbDbi6vU2OyIAWIikfJqG/FwDTioms1ZG6aTHJTTOZjikJwO2/OQTn0B4R
8BXGTb1txNcosSQUN5rHNrF5TkrQqAghKiIXWABfbugnrwEmCMzH5FWw5Nydw9+5
lHyftpOkPIWz7nTxpm9MMDUeVWkAqi/8IoaC3xmwEm/C4rahNrYgmO5t9VVWK9mP
c31KEL1Qx1LRp2runKTQi5MCEntUr+dJ0DrN7Bml4odan572uvC/JZ8DfxhWGcDy
rfewd1EVhCEjtjXpJwgwNOmZ50JEMz9h0GA10gPbeXpOF/joU5tc83e4oiCdx4lb
ONXofecg+f3rDMsKp4eSJeWe1O2ilgOazmYeZXQaPbV+yhkBDjUBdZSvYu4U/sRx
NQ+GIGcMrLdO+Zdrib/iad4adZGNTRuwbWEEU/Wmroyal40PXlC26xt5Yu/qOABc
lu1onj5M/rjN0mPUSwDohoQ17v5vcrLd4tYQPfCGmJJJLbAYRWkSjsRRudjRnCuY
ExZlhxkk4egXGUGYrY6kJjGrnAW06Sxeffg/ZiArSeYjeO++CqJ7kyU+hRkLTKAD
q5F4yBaP+JZDuTc+eSrnI7Avsv31zwcIX7HhD8lvduf/4ARIITIN2HIHUvnm7VZq
hogdDnCa3sYF9GmqhlvVg7wKjj9IdBMykZkbzyXgy/iRQkFPKomOYB1YrNgAiZaU
J018TmumIjoJGOWEbnws/EjAf8ZakbabQbuQ9T0RcGfDIPMi2nsb+Q8PfSSqJdYm
z+Vdk+Hopb45vyCZ0lgi3D+z/d8+GCaiPtGZ0vfPjN74+CbMM9f5XlRUw4vViDXT
2YidKoxPutUsaPvFVjOVaMCuT4+O0a/b1nfL7HoCEACgws7IzQ8s77h2ssYdNPiR
KQxiCRMfzD88aSZ0bU7K2GHm5Og+Zwg2/yrHuRZd+lq6+CfviPg5DczKzB4kXnPc
eEgWzzEyktwhJFwZ2dFCtD7Zx9xWJOUU6kBvBLGdYVhl0RBpmfEtRep00A6TJ4bJ
IhI5aZqrORETWX0mqioLm7sbVEcZ2t0/bCHYxOBts9q4aLV2vma+RhPwVt0vPHGI
QPKoJxgC91r7VT0QRd/N9VS8vYMil3VYnt0HEqhvKwSqc5JJzQpxEtykaCUTYwIn
QV3djGi+qFm5lWU7rwDfPw63lXGX24OzZFLBsyMBJTA3HkAqNToAWWEq8Qn1fc6N
MZWa8hPM0HXXHu1ka90xAGduQw72IjFu/M/P1wObT84yXkno3abTypAef0r0PjLW
kiXx8uDAwEoJtvBlXHSwD0AiWdcwSbVqVK/MpwjLGxERgGF+qiX3QIcWsVmOZT8a
p8FTILXV0gSPlWFDJwP+XJg1zuMQy31w1qZgZnPOUPfSQMl8K2RXgx9+PkTy3Iap
aPJ7yudHNN6kCTMGbrQI1crA4LRypxjp3QlzzBsfjSESR0tqgkUX7BhjmK8qShzl
rNdwrwWKVkcNxg8MMDMJcnk21Socl9riciwB9umxNMLfaGO7VZIWM3tg7Bx4NgVL
CxDhLyMV/vURkC6sPIiaD8Wi9Xkd81ZpFMrjtqmMSNx8j8efamq7Nnwy/VRsO64B
d2jP/xrMksggwcJjyqD2Z2mZlVgSyBM3bbsROzxE4mdJQ2eH6G61hY0HTm62iW7H
L8qN3fNXITB7W+ZOhOoxzSwH/zpIvmhTdoUhEepCUr+tmD1s2Vcb4jrMQcgIBX36
rduu4vMR93KE8B0peGjwRozHX57JwT0P5Xi4zzI0J5Hl8DvByMKPwLYnBv/VDdL9
SH+LQl6wwYry7VQxJcSb0hk0j9xdugnV5uy+D0VC/n6ClJ4I78TCliQLrHrG2okJ
fzwCnqBElYzRxWqE74mdbKVGazp/T4d4ffXYEl6G1/FpZl49Rm56NfOfvoksEL03
N4pVdBcb0iwn6AswHzp3Ao4pyzxlUKJTDsQ3u88WjXiXkBfydACCnq2gaUQJWN0R
IFtJzT0Qrpk3tBvWV4XR1P/9fA6p5XNNDYXbD16jICi3djcDty/egEzg364i90ss
OTX0+lX0xtsvlANlKbqAV43kmb1uFef0rjYR26knFNG9XUbMNDoZgrdOMp3ARXRL
L4IZYUzJM+94i15/6RExWhUyvlUb1r23hjFgkXJBHY7x+TW6HAIoKAytQi4cshua
OLc6Spc8SNdk5UPs8JCm0Ap3RMjm+0gZ7KvDVaYe3rrfYK6hi6eV4hJmgKJxK6fw
aPWFQWqGR0D+GG31VlwbIBY/xEppOvS87lY+IvbVZcCmwvGFblxGvYfswLX/Nx+r
az+CiX1qPFHw05KAlJx6jt9bsSSklnDYYsj9/sUAxeyPUiMDEy9B3pJG18klGl4A
bQiQUipSEhZP+IUm7dPZ/wsfRe9cmYTbTj718RbaFRyoy39TQKieTJpmSYiA+sJk
7TBM1hBTVPwoB8jV4J7ZKDh6Fp7rMfkW+x5I+3asEtGIZxeBnSzTArOEYQMpzN8A
jNsgRwo67mAL372bnW0WXiFfwQf130eO53FSi50qsGcl3C/xK1SubRv73Nar/vz1
PfcL0kCaJkhuPM1rmZJ16gDiP3H4Eug6Bau82mjH4a12frnOoj1AUpdUeIAZPP7u
VqstXYy4tbhjI39e0SFcqZq0LmJLREFhF2q0gW1eex9r7o3ez8/1Z7DAqoDUr/is
mNwvyTxidhAnL8GjU62if0jJuMiSFb0zaqEJ7Wq0ltLjr39oPgrcBixnAmNP8LaI
mH/aISPZa9GmtkccDe6cHXUElLu6O3mCmFWfAUaZIrhoexJdz0sPHy4Wzfu27KjB
MAjBEJfD1HeNNDZfgTXnnE4PXnrJE7r1OikRBV2y7uJNTgc/xe8u+1GmbzQYspP1
5/sZslyWJ4ex7n1zBW9JhoJzdq83m/o7QCecOLTukWK0fBg271//72sCVGnoJN4V
VyLB0VAvThOGcIvY19JnVjioQ+pY3K4gfOEYdqz5oXMPSlUaBdG4kr7Xe/FjeUkI

`pragma protect end_protected
