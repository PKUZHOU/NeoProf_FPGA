// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
AKSVxdV16V4zcDvDntXg8Zk27zY/ITKhZT/S+JM+Knxk5x7aFzBw+A6BEHvC
HQvGIWTNeQYs/G9dW/bj8UoYfR0jmLH79NYMSuTb17cDrV7zhG+MPstk3gSo
L8F40c09loNT7hT+zcDF5VwQxCy/+a+4y69f4Hn0H2LPjBnkIaqay1XhnAfX
a8EXcmMwNoF2mEvU0nikzaRvkbxBCVohSGSRAmLqI4mGLaAmUq6JbHdtRhJ1
Q0UV8oSkqGib+jf2cQc5OQdEeKLL8wx1YseJ6Ic+bYJ3eSR7IZ506/Hnj/UQ
2MHO1gEXQpYpCptpZakIo8Duy2BySaeQKF39sjEY/A==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
E5qfj1rQWTM4K4Z9o6z1GqFBVGkW7VwMqjmf+SUGbyAlbQL2B+XsEtaXG7QH
/rxyZvy6l1CJQPtpFdKoIPrMf/Lt4tHXGmTcW/DPmTPQjnI/Envr13VuGl7Q
ppF1ueWhTEpzNIitNyArjJoDYpvw2eDPXuJR97eSkb0yjCjDUl4Cl8NyF4pj
Q2+glVJP+bOegISif7sNGLMqHDwpAlcfGQR8YRnpjkPn1CEa6+OgfQ1qadot
T4pFK5XUCB2j9kTKK/dsY32Kjur03B0tjaGdUK2c2Ule52Ko8h7+TM7/nVzf
A2uRN/QkmAcawu/yOM2xcRIUAvlYuqszokrLhpzOQA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
N9oYMivDd8KppC0ZX7/yibRHPOdvFLCaxXNphdZdWVOCgguM/6lPhzb3tZOd
qiI1kmwn3qyxK5IAd2G+qKRR4k7eXtAE+YrSFU5oIqRw1rBi/7QTg0SUl3MO
nb69qLY20EitRv474grxiwpMCbLLDAq9oowX7gYxV4l+rI7tQAAJATnV+ZwY
fjTJsOKg1NIkblMRqassHGwsQWfFj+AKvG2e4HdjfOff39RYlpt6Oou2odFk
LxONA9RhZGCbZzJtPGcsu7uJktQHFESk39Qgl/mUO4Wd600QUhF+4WWTrDhz
qvNOrmaNRHOkjluaOCKNwJVDoaJu3KVBzoh2j+lUVg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
fr+cAp1YFjK04jHFPlOYplLYT9pYjKQ/uTYuMHlyxPU2sfT3qE6DPDFyj/gj
kPQ/DZdt38hPpIaAiTpzkAks5dMSwyupGsPl+X++HemSWfwMZsYxV29RrIwI
Fiv8lMjgpnorpCEAn/uJAK4y/Rg0YEH21Wmop9THXFSB7uoQuSI=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
derw7QzIL8PlQzW4I6QKGhazN5VS4LFEYa1RiXsFtORZiqG8SvqcFYyeuReb
GOf9VQ73+h7S9hRFH3keg7OeaK/aLvUwXKbk+N/VwAbBJFxgDaScRtzUzbZO
W8jnMmmkXcfuZ2XdxOoKMJqcknE8XAPXs5yfMlLorcypzWU72404uVm0za3m
0JnXqVSFfVaEMrUITashx3uP3qRyPxxmT88arVUfnG0ts2VpqhJY521BfZhw
pUXR0Ehd9CH+TSUCYThkevDmhwv9c9GIu0arDF6GM6xQnHpZIJlwuDSSLAYi
heOVnCQCkmHQ0yF+osFjyL9gcaDmvoVTLCTYrpIcpAdxUUmbLfca2aqgpaos
FiCkUjf/aiTP8TVJLdzRr9G7LhyYXo+It/L9ao+pHOHAPWS7sgOGGOOjotDL
9k0CrfJ4VLlCWn2KO0iuC2ibPR4YhqUQVWqvLfBvHEq/YqNrPbEA0048xprZ
2EosyHETRWspX051Vzf0+Lu5bn7Go4uv


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
YZw+3xWT/RA4Jh4fph3Vaw8UC4YheBMj2CazOlUYyjxEYuKw/6sTJ0u3WBGg
mD4CellQLr1Fgyr31ymdgUbHal0rvxeISMi+VJ1hie4xInadpqyl72Etylu4
8mJLv+uQi0GIaQBk6HFa4etXY25IyMRnBXUkLQ+98oax/OsHlQY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
VF9igUasDlMo5DMs+5sRY4TYe9IFQ21XDkT6gyeHKSefgiHw//tiLFXsjmx4
LkQQl4qeuAWvdW9g1a8CdKc47bVWpzVMj9QNjwYylht9KKocac4TBQ0CM1cM
fgloMTWoAwxqN5jHpbydRlGXUaxg1SfJ+nY9XLGFZE5xfrbSg7o=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 16832)
`pragma protect data_block
F0HGteJFgLmDesI30sQCbQiwhlOWnBoknUoEEh4ggzA7li9pelX/HVLrrat7
DQ6iS5stmSnMJVHvwqIm/pBnZlop5FRKSRq7m7BEbMOTwU/CDZHf1D4PokrH
xLt90+zSEbzRo86JuC6ckXXdheBDeVZE0fnOBAsyC3Bwt838UiOfwyIOFDZo
SUdlHB5OZk3WFF9vVxRfnI/LQIyyRJNmr2QCihko0MJnziD9obVlKnvYbzB0
pdVDuPgeLpiA3OZT7yCh38zVnfCz+DdMjjEf3cYj/QJysnkvg46UKN6a6jwU
DXrpo3qFFj/EJvK7XYHMAm+eCd0ukHEXizurz7vwx7BXmg/rr8QoMn7Q68pT
YOwSbx/WdRrDgYSaI/3rvMn8F58x5KpeodzhmF4o7Lu+/8Ui3IBQEX2Wl/A6
FZgl8bagoKT59wkakhdDxEiB9qNbZuDu3S688efm6AtZ0Y6zhHg9uYCA2Ujb
RFT3Rm4VZrVC4e+rd8LDuo/UNyyanr8e+yHxQVnNDqrC+uKgk8ZpJC1SkJot
0TQNhm7oF+jD+eJUyUt8POSd+L+c5a+xRaY0lQ/6SxTYW+KgHnvgcWveEkS7
ZkXrqcY4c+qKVS6lN9aIxbCIejBzuv6DxVkljAKmwccYz7y+AFFmo1sAgsCJ
kPbPutd5DWDqW6EWEjMxC80nxZrTXC8xlV8KBLCEcx2K22Mouc60EYxyaFTL
QEP+r2icUf2LG/QBRJM3D2zpdDR8/kcuHZY3AaMoQfM71ClLZx3x8J4BDXan
VXcktC6w1AyurlgwO3UCAbVvfjyIlHVdFEHV4Cp35CcDMLvVX0vNfLKsVxUx
X2WE59NfrL9zh0obg/47ql0LxitsL8NAd3KVNr+XIygV8YyZqvSU/0Awo2j9
CgDLfZ4mrEFV9lob1lkx2RDQZPONzTPfNYg8MLV/TfYbUgceBOsLpyfuI99C
W+o96UtpYqrcy5Ok4ekVcswnl6n1GlPau08W7B4pMB8+JrdUxt6MLISQKWqj
L7wtgebgLsOmcvSiiHMZb6EjsIgMlZIVG58m84gEPMq9wcunWTJO3GykGY8V
qb8U+PkbJ2dAG6gnbEl+YJQd65egNKWlwtlQcp7lOAJaujS5GWsbJG5Q9gzZ
miEjGqW03Y5g14+4uF7N7wGO8OQFZNkh5abNQfJZ8kdW6jh5s43QPNos8yw5
w5qROfsGUuoVGhuT9OppM0a/cBvsw+ieRbQ/VGMSYSHNa7cPnn3Z4EgjlMiU
bs6KdSG7QvyuFzMAxEJqVoBJoPNqSqpnBBE0iqs73jsRrd3JGwxxy1NY2T+s
WV/62akqbuEEudMAW3nXTXsGWdofp30O4yGbEWJc4wJpu5K2TnM6mV1U+dJ5
+7bZnm1JfbGQ7+wF5vLc2TrXh/sYnQVXvux99SMbEiVMUX0whLNaENv6Ww2q
wSHvZj/rjYD3xG8Y9GhVIPbTXw2u3OFbOBwbdDlCoey1Y64FJeyMKEDtIE69
UTpSxH0tbpUQ0LqQ76vK+URYBdKIJzsR9hpuxKng63m/KKi8wKu6hxCbMf+V
rA/TbVk/ZhRL3q+ltUE+nTOczSI9ewD9ow3oxiBF68vC1+w0pdaEEG5yuUuB
IllKf/kBlDBy2EpqeS6B4MZ0XmDUFXLBs/AQlGzE0oEjDohIGlpbq8Ob4OOw
eF+2j7apimtHMV0YHeA/ykU5w3DBt10Ilhf+4Qb76rPLRsLUFI6FvC/PflDC
5vgKhpwRMhqWDSzbRJLPHLwh/HpmcP4Japow8xStYvGzhlG9coajC/xknkdZ
5K9L63hkQ7uWpZxf9hSLb4uFg54aPEqgH9EPVwHU8QqjHKweUz9FW+pQZrKD
40pcetvKnMLUcbHfaEc/yOp0qHMLi2p9XLzOpgMCmcygJjWZzWsqcw2DMcaj
DuVzsOeOXP93JVI/2+AGctuQqManGwhmh9G/GY3c2eySukaUyEj85KoJNnch
h2qjdfzoXHeIIIljQdba26oFYSwOh8WcWOyJcC4hifNoBbI0RvgtvjRkOEBk
JMeAXdjSVT0OoH7VEh/jCMXlK1PH3jdaBjj0g8mpasYOstIfAl72BZ5yWiog
sbJYSfGrZLzKScSVQRo96zm9jKi/I2Bz12bjotW3XP7/M6gaVJphnqwSICk4
yIuZrSAYfUxSQKrz3vaZsbEdiWwAabkieTj/4JdJRQUe1p2LLxUf1cBqtawE
18fDD1omqOJQF/R/guL5DHJuCVSUDSUoR0mPEJgefqV8FuJ13XiryJGlcC4F
CjFFOyy0s7GyyU1yOrC2l68HHzk21KJgFKUJ+iSVocrwaq7mi5T6zv8Nr0CA
vND7divvIG/tNYv5tKTjlzrI+vIqqU7h+p4O3z019IEk/DEOOvfZF9A9LZJk
ZFTzvywVO/tpEnIPSn5LMlR6G8u4eiGRPW4IipENVaofC44kmhuQV3buRvkz
IYhJOxpCw+3M7OySKBt7G7bCbSjaN6bUCMwInqCo1U3vv3Hsrb42Hp0KaoNm
0Zva8VhN4yumUoZxYjfqYXZcsZtqHFJNCvaLpWtJwNwa12KDxBBEZEPG9xj8
pptaeAD610Nfo/6ZFjnJ9qMPagFiYUZCocIJN4zxlryV8siuACly90gKPAPF
GgOuNQywW86ojHmnKhWp9Y/IcPk3Oz2i58cRqzKI20992Wr5WiD6Puya0xpf
KuLubyFQO7yeQzhyNrAR7ndxvQv+uenm/tTmVzJEVrcf+9wlzQdL8D17u/7x
sRr1z4l2d0aSjTgqpNoDNmBBtRv9hobyAk4PfAIk6ig/SCCaH9CGY4T6R9fH
9b4uO4QITg/wf9iueimCzz5weFLBXowVYe/rAT8M9rkym2plzAVA9tpWjY62
9oLe1TnkKXZ6U3/u+rMJjd8+vx6W742zmQxkTHb1RHKsQags8xqTiQDlw19c
i8sC5bmhYlodzgG0FPnVsxGL79P+nl4x5JQeKflveKyd2wAdD57zkCsOCRAi
wJ2J8LdsrVcpOxkIzYOgYbr/WGyafrRvan/8pmUwI7iv/SJgSD6DTp1TLD8Y
yjpWQc1b8MqvLkxaM3P1YceNUXZENElQ73pLuw9QzRe/8ugVvu55Wv0dW5FJ
BuVUVsP5LUQEGFWh7SSClgXsi5CVUkv8dz0E3gTREifZV8YHtZHRZ7gp2iPR
vctAVtOiDY5+hPaDYX2aNeOEubGq1esig+13Yt1M7S1eVlfJPAwXNr43kK+i
RWWxN/QAEdjezfSHXpnIjBsh4YpP50EqiG/6vJNZM7N+GFcztjBC6Talah/Y
1yaAcgJS0WnGH2H/5m8x9+wTfCVe20jxAHCsaDCqKPDgoFWOS80yHplOikdy
r4PMMM15wl2NeWfCapOKh3rpjob3nMjJKb/jitC1LH1guOVqbFXTF8lbbERy
XoSRgmsXhEWSRMQ8vjyEe0OaF21rLd7ysRjjTtJ8zJ0gUtMZmwyh1/bgoNgR
1+Oub7sXxFnLn+sox5zaG6SNFHuY0QSWKrLA7wFbbc5Hj2XYBkj4IQqyk1ZD
4OM9jvaDSq6NqgSW1YuwOv9XVlGJhhC0mk5F/XWCV5jfB1CiF5XzA2cGlDtq
IEdBpzgLfMQnHpwmbBp10N/h4sntVSNcsR3Eokl/7dkb7F1ucvs5UFiGVsBw
ONCI9/bx4c2jSJyXJslkSO2q3HDLTj3UHs+zXRBK91lAcYd8fQCbBpMNgjgA
ap5nF3HmxJ/YmELBAWsyev4J5g+UdLHWgl4amg7PnOaVHaOZVAfXmsLllKQR
pK+2+q3bpuU3qAYvnJe45jzuN1mDKiWYVcMpRrPLxEL6fwr8SWWGz3We11vJ
4apA43iuvST8uQ7ltae7RlxXBaM6EjAAtqbftdiZuipg9pBlC7VZySESlI6T
TUoCTsaMx+mvHdkou44Y/W3A2viGDS4oe11h5eyAcgInxjVljT9XCriq8sQ8
1ERb33HrYbyXP3bPnX4tYsQ7DWutWVvSpi/BaxDndjnIgw0hbcSoSxupa19+
fRKH6Rfysg8n6tRyhVzP2mxawXuRD787sczICmkWVZRT3SnNH3pZSHjv1FKX
k7UYaXMHRd8OS/zaF5kAvtiPoUNiDnuwpoKPwsH7B1Vzp/AZye+cOYcFkPgg
LZ509bO09IbcajPCvNUorVQZ+DBEvCvFTl5cssLdF8ad/f/w7ymIUBP8EtYu
MjXynX1CLhJPmfmRdCOBZbwbyh1rQEYoBfH1h9Znq9+TR+oEQZTnvjiZDz99
5FBoctqeDNwmEcO1ldInCMBpbasd4XtsnbxM+4EO8cp2tZmNgh91gKMAGAE3
vvxgsY9SqQd9Cp7mrw0CpOA+0syNVkJcqGQsCUZhcerrepviBEfPuMsODyGY
etbqPOPxyNSa8BPg/hU6jfbWYM2RjyWvCyItIQo2ZmuhHu9wshj04PJN1MTn
ypjSvDRFE4vjxN7u4Ch7p/IGsnX4HGiVsP32oJTLLF6uu9nZO+VGmbeVmjAd
vxtrtu24Wye/puwl9vUWTKgLuF9a1fdaRGRxmg6b1sghBg7CaICNZ6XxoNH7
0HmK/NpAwZevDUuF1Y72B1Z1GvLupOqNMaIhsUM9FgoVJ3UUWwt2TaybLD+N
hPGkjxycuXDZBOG/LqG6FPzyR/Fj98EYqz6qzybrtZwZRmfB23bFr66n+dAx
X7giCIMklSHc516N0d5Sz5WR7nayrF8la41evBW+SXL6H+26Y22jy7VQqvBq
gJEb9Vjw07UywhADj+OVB3Sj75vETD37WqwJo98MRMNDet8dLA9XYB3I5hsz
kGebOiGb4uMZkXi8IQsaEDUFlqA9QUjzCOJIwZzK76/nqZ3IRoKQ4SuQBPk9
FuphSIL7OsK0CTCvD3zRArRmNgX+r8l+IL6C0fzFLQm1rukhAwe99WAtTwAI
la0RG7FABu9sqIAUnMbhanvJGVjFbLs1MVm/I52TKjlS5d45GoAzINCDC4aw
4Kfy6iQ99zXbxYaZn6Ts+VgK800yb+lV31PgAohbIp4GksbyVxHMzgRa1eoB
jHjhRZO1XWBW3qpOKtt2q6HRA6AYH7WtJRmVdpnZKGIGlhSHyzwlP0TmOeJu
1L7d9ERDZBw2vhWGWek+AKmLDvPTkPKF3YmC1/uyBRRN+PUCa46hNDYq4JXh
L4gRE+VKCR3GsSzdEXbtjClJCzA2hzJ5r7+c9GQ/rZp0CSAlb2VX7rA1U97V
r78xgwHpQEx422PgowRgFT35WZUH0dmtobOAC5MZeab9BJDD1g9WKUAY1Q2B
vx38JDgB92uRGKvLz1bLjfxoz0X02FZgQ5tcAJJrQnnwru/InYvcNBr+ha5I
4iifmIQXwkFE2VP7YUtOxfLEdqEVZCQpmUxd0XuW/heFsdKM30Wa//OX4YX8
IW73TJj1Vd0HS3P1oKXzKFYD6uvsOpof/+3IGUy0hmM4lTpyjK0klnphqWpI
NX9/n+IdKrfJ+EymqakKqFy/vxgYbRJ4m/BBudvS6CNq3OsLsrCVD1rHlttk
FJH66QfCsjWskRu9PpJu2gm7J8q6su91S6B2vZpCxTC6LG4srumjNYSr6knG
JxurHBiWC+/k835d7IiIv3glMo+h6SCkmkNhcibiWEtyhkPkWPcomVDONz7e
zHSTnD89KKTCDjJA5rWvxw8aJmv0WsaDS18ldNe+WtcpA/N5yL3lfx/uBsbr
GY/B/Kt/gHIMPGQObThKA6NSK+ZxIVVNdKAJnlkxxEIOSR2zG3C2iqPI12Xj
+7BX/cH42Fr29tPDTGmygO/5dfXsT9b+tzqGWEVVaufQuSZqYdnm7lWUm2aZ
kZ+n2A6sJGXiw8K6TIPG0qXHKi+k/wZ+lr0WIhtbqc462AdQznDwPaTpFfL/
r8Qvo4nNiO0M3iC0OP6aMW4g9JfuBQlxNyfIfX2jIqh6LkawcaD8Ac1WWkWv
vHBG3CXzpzy03KuoGv2suSWBxvqSgekE9+s4RQtyiHeEbQyx6dJhjDbO9j8e
gYkBh2fMEDWKQdQJU4sIW15pf25afJ3sQUCpnN+rY/9cCi2cdpLyBlHovl+X
tpZtdgwR0I5CjHx4v/nXQI8/F77LiATm90ZgFDocuRwQRzDAhxdtOsdizVY7
NUd0tg+lNYPJVPtdwGMWaKUJPYe2OyxeKPdus5rPm+FEg31tdkopXqX9kfk2
PYWXJbyDlTIXzSp4Oyx6ZqMhe59HRK6/XwfD75BS81P2FjfEuAu+KrC3Dz3O
WvvBcZd99eO8FiQPOVdIIqyzhT8lSp3TCiFDLHZ7BW0N4nn8aiS7KyKlP1dH
82+qj5W8Hrc1dVGiHAaJxPHNCndfjY3sZWU2x/2oZLxuKrScm9i1G/DEJMRM
uM7fjdFtAsdEjw89Nj/CKEk4AH3d12hR/7bUM6qtTMWa2wgi3cZ1bv9n5wMr
5lkMR3o0EAq+mtUHTL5Od/vAIWHWUM+SB8f2MwzGgcXvUchTv8580/PM+0ZO
wA9h2ux70yqIPC+Jedc6oORGmOYpzWsQyOqE/6fYnvJTCELJFSzkWJzzeVG3
VyTF5evcTGawYjrel24+JuB7d097+7dIR1mGqiv7JZsJguQCZxglBcOdliuo
gXJkc0zRLIVAtEbAgmOsYm4BaC3fGQRd7euqnIVgYjLVI5/yKKXPuIUSm6D3
Kzq0GnJ4V/wztHUmz08+fcp5kCgc6uvOcSPYCtQzFBdMeNnoN4yv2z05j+m+
MQyPN5+HK8eF3d98nd5wLf5VTv/zKZUCEGhO9QTOXRIRYXV1r1LdSeqZAczi
hT2jM9Ce0Ixn+nFJEIysSTDhC4LPQBHdgUNbMlr0TLTRxpMhbx4ZhubgzE6N
3V0xdyIQ4OE+XVsjvuaRrTbiyjo9hMPPjPxWp0hAdrHwyeCsYO2z9hOMAf4J
XLIvVehcJ+9P/jKQLac5cDaznAAkvJvLwLQmyxnIMb/KrK37tFLnvgVdmc0i
WAtmyQobNai6f1izCCJoAkb4uqcgiIn01IYwNwKmwQTS9h4hck5zYNnDkDq5
T1rME9UTIVlPq8Vijm3qss1MbCcrs6mHhMPtvsyr1phg0t9ZRqXnMtZZP9Py
ptnZObD+j4eQ5jyG/ots2qEdXSv1oJx2JCQnT6rQVTfhHXffc2uCgSMf0Uab
oo2v5CI68o8HdXieeMJfuTJ8bYi/xtyvZryAP8+gqXLdPnvmzfMXJz1TGsf0
ASd3d9YUwQ9tgvY4wIeoBrXgp2box7BSepQ2qdTyv2TcyMRSfWgxzHONagwE
7xMxD3v0UQSONQl2ojcXtn4vU3t6LptzPSin2sz34NoPfuWhAQcnWmYy7x/K
va4t6FyGNBRgFOIeZzyD+E9jzFI6/yRQjt6LRxICStUGCtC93NPc/xmT1gL3
A2LmCmv82nmA1S9is+9X9SjqFeg/OGJ7JLgiL1AJreDFTmpRGt+6KqyJDtiL
EDDS4+NbcqCU0tFUUJ41n1KCXSafFT4VQccjBWoZUit6aPITxv6INMKc9Yij
tan5YMjBWkaBHqJOG3AE1lp3jV5kol1x0RqtUUnF82zbEI8tZaBGFvmZvwVS
kW1GAYrwz7wjvM61vnBK7ZQd1iyzGnj4+I1vGkOt6ReztXh6k1lUnfs9U4Vl
xsbzJOqP7kPEVRed+HhYNcFhBqSPybOsMxjAyxPm0Sy/oaQnIq+YOj9UtSMw
JmMseI/fKSxgHgVBKVHXZ5Wmr8ORYYLlRTgkSqNSkJTpsL8mclNM249bXU1A
iTwxJocCbqdGYpcIRQAgK47dK+12FFVpLUxjaaLFXBG6P8QMNWWDWEUstatM
yuCCGMHlzAwcUn0NGyXJQ+VN0DSK41wN14l+I1uXGyD9wl4Fs7MhiFnVb5eY
Awa8spaTo8tdLFe4fbZxAie9+nyZCAECplewvH4RXYWCu1+Yri1+9B2A0JkD
TP/ULiSjtp8WgBcn0bl5aaHCtMxUtEiPlpq3X5cw2IHH3+ar8+Q8kULFiP2e
HIFRIJanm4L4aEyn7BolHz0wGd6bEsbXt1c36y0kuPNWYfk/HFFT+hYTOvCu
4/adKcpFFudWlQJOxhF23JlhI+YBFaTb3SRp/cHmy4IzXJl8RFyTyR7g8Lp3
n50oHhm5FK3oMT6VS8CqDv1DqVeJH1T5BPtCwsCnj0tuOFy3wPbatvIWgs2X
w4Ci4LYEVUFbycMNW4k+kF6N+XTMSiSomnr9HYUA1YhmmtFJ/yvaxSoh1lGW
rf5+B1Tuet3pFy3gwAQzwwwYtf6wxViiEzboeNKyvostOSFKGxOMbnOuWs14
ZqOYPe3L2qtdlkcMGdfKsQGyWsZbpyac2+Ie6pt2cgyJ+1R51E5rSgpi0Sax
+M23J/Tn3fUnxGwpOwa+0YvDHT0hfzHB1HZ0Yv8hJPAC7QpvK8p9GiffvDOV
mZkp+sH7znYV5Q39VPO46oEDm6z3ZYbMK1ht4WN5wSk9UsyRoYjXr2kVZ+LC
pWG1IW276zoDFYlk2kbWnWOtGeJdsIKB/c1lNPtVZDRKyeC/L0j99O+tQ9kj
4FgkGk47obAxDmtckqn/qAED4g3cMDcdtze6NoUYph68jwq5nlCnPSHPn5vx
VLuPryMB4PTgkhc/Y5IqzD0gXEi1V5c5Sp9rYjxlul1QvXkbM9WJMhOS3HKr
Li/6bcNsi+gxCUfqeMJrJVBmIcuo6R/ZLMjcSJn64BnTNO3MPNduIPQnsBvL
T5D8DvM3r4m0JlGsBMRNGcIGPUauM1aLKITugJcyxpkVcz9fgtGfMXjirOdn
HFJweJ9ZtxSRs76kDIK+tkNOOfdmmf6EX5GjhcLu41jQA6rYNQjlwYUoMWT6
A+aGYqfMkB+6xjMS0woQyOlkJWhQ1d4i05QSOns0DdJkRtcX/0Kn6/pXPFq1
XyFJQm2VUnIUELjY3l3W/ONR++l+j2h7GRn7D3FNqQGDKeIqZiHt76+iXJth
24U63FfURMVkHNmd84dp2cgjW77MlX+YkyZf74REdOc0coIQxg/J49CDQyA8
xovo5qBBmSi6KhxszsfuAzVcrjkW2NUPuO3OiWR67RQN1Qt5gbenxQ/lM4gS
yLpqo8z3nj+42t8M9KC3ap10hG8cJok1zyvlHLNZH+DLV0RSzYrphHiifKxf
Wy74zoiIRHXrq08wCcYdWixflbi3Ky9/FK8qXRSgmTClCi6LnCuKs5vmww9r
Z52QD5wxBt9yNr71BwmgrZzlaZECVdCB+FH5Nimk95QD1CzWAh1WnLjCm1LG
NYq2LpeHkp4AvPNtD+y+w19EG2NCUe7xs9PnAQFFKMsreZy4WJXBm03rqDRy
Tri55I4/Ufe2tStFI/DorAHaWJYQfmw14aD6sKQvuCfRlb2kimEV7k8upsxr
PYpT0+dn/KF6+yQEdP0K+voPVElBMVV20X51ToSXFkKSFoMZ7FFswyVgZRbe
S2qqLhaGXezFq/Iuod+/gmNIrHPEIZrlkfPmxu2N/zSHGp0PXMvyiOl/WKFf
WZnoqEJJIKoNXMNeTplByKYm/zixLz4NHWOSvlW+VbGxebdzr1aUha40yZMl
UjyzU2tr26InXnPo7BPfhyyzL4T86cJoa3oUDfEAEnSfSJfUlaPALsgSyMY+
bNOmm4Hy2SKtM3UmgLPKyT5muJCsqmJwI09pXIm9Nk7D5xXqt0tVhCDGeZ31
6uRMq2pA7bZRxjNyvPWdTdvIR1IL9Vz5A9Mvis63w8LkrzXrypm93VMppJiA
SW2134fuKK4C4NYJOqlT7x/pICtLYCKK/2AuI6WATYFHder2GZzVXyGJsRi4
svr57shTmJzP7g2iSjDj9O/vm5hZgPT28w35ydbEfz8Py8mpEdOtG8l+g24f
vtPGHZjKuYIBdN0S0E5VhFptHQAV8k91KT5emAmBY1GuEBZP36kAjX0kVJsX
0hMq2iP9/f7qBFadj17PoCC4ST5/YPa0xKqJ79CImXZKmC8DNjSuxpgAWbfe
h4VKyWqR5GnVk4qHRBHf3e9s1QmLFZUiwbitCu9hjfJ7/DJKcKUzu9mpnacE
7mcb4bNCZzEQEioIpCIotVhI9j7X5muka+Bt3TXDFpR0pOpLBJrgPw8Gb9ZN
O+CmCx0aZOOQ0z7Dp0anjD9DUAka0afbhID8jhzOqe8gSqP88Iy8+nkSdkwS
YlUiNJoWctX828FpoUP2RvnqJjj/c/74dY6UzzZt5NU8h/oOhlkx2E6WBa9h
O+dqrBD75yj6ViE4KdA0hYowokSbmR3c3r5ir++Ad3+jrKxidyw1P9CJNDHZ
YJb5GSkVUmBvjAR6cSnp25q5mwgFPp8RdVyxMtsVu57ZTyduxelN1HzH+zy8
9c2/SelnO22F709GlgA5U0VFaGS29aTfTG89ACsTQg5mc9bx54WOeOaTjtEd
WMEO+0VJzFOeq5fi3vajMoUZNKn8LxlOzsGGSmBxVnLKexRRZ6+H6Od5Yh2p
xa/97GO+w8wqM/BgsXBWWLXvg0J2svSi+zGTJsSEveNP0wWKugdtgOO8gFQP
WrI5pO8jNsDcCr7WWZ1t5g4O6UxoReT6DQw/gHx0EbrUdDWQ+kfj+Rq/FTJx
uEu3MCJajwz9RJDLyGfCy2WVtS5KO1G036srveCJDQTxJ0/GizzacumuPXzI
AwTv7N/wSCmAEW5HlJJU0ss8NdTWRd3An3BCwxI5W1PUWUIw6UrX4Z/CE910
87h+cleWvaGFQYqXQNlC2sVmA8V/OkcKm85fIzole8ZjVVR2aggH7ONYVtjk
NqmIpDsfpDN2OcYJfSW/2uD70P1i23XW1uTeUlPWBD3HmSl1xHsm4ZLBIHPT
XjR55JvDuy3HW0/pYkA6e/EFDd1u+uOOVl0wE8vviC5qE1ynOdNyOh1/5p4C
nOn5cSSgbLrwq+D19pCZZOTutkahUez8T2PSdwkEMz5u1UNA0tRvg/MmzWWn
iKid8b9NfBTlPUWUJ83tS+QDfZ1o/FwlFGv7HUqu7uF77ABE5Lvxg3dK6U7n
P7OBz1e8mecXFVD+mvH+e1Cpgjjs2F/XTjh5QDOzB9+8p/KEWBMQbzAoz6CT
fLND6HRnp2XveRpMAk9uABBkakt2xtWZisZgF6BwP7PAnzcRCrHcV0ZJVIrZ
rLRM3FNRAHXDDu3/UHRhAbqwZ5UW18uqKptIu03eHcgxC0I1YUEoVV63zi2U
iYqV6UmnccIfZDratVVLaUPi6zegnf+V3bJ+WHrdd4UNY0lcAaWKcqEG27To
rSbUBW03MgBAtUD9UKmJ01kPCO1xrUKi/O4n9QUuDhbsIvoj9SES5qHdWrXJ
vEgFC225IgBpuaRz79fEr+rVvMrNGbhAgrjTcrKSYxYa30Q2v8RgvY20E4HS
Y7abHD/vnpTb7WH+eoBHUF+s6MSey19nLuaqkklubgqSE5O8CLbqv5+Pu+ul
wnE0Pk0Y3Hkcbeiw+MGnR+HeSV3rvdYcOYchFkNZSXkJwGbEbnek4pLqByfH
fvkCWnMjGEyK+PHx2Vv7QIS/5TUSqbiHHxAt+MwaSDeacX2dZydLkluALCZG
hWBgdGHHzKXghPgW7psLbaGyDRnbEDOAvUvFvIAialzchR0Yc9noe/1IszGn
fllaj1IXPgFefgABgsy4avCDJFfxw+O4H6obF51Qy8BpxO70/zTWzkhz9qEj
80ECiA+qWsw0NKoq4K+BC8BQX9GMLLeujYzki9KlRTx7Dw+Xc068LptRcV/f
uSyVy2oR6FbeJZC0AFURUc8aJcl5K8QrA7R8HI7NiVOPSfAokdP9Ynzwld58
Iq1njmUtpfnD5iPE+ouqo+OOsgq/wW3d9bvU94AnpMQOEV7jTPhrqS2VoEHz
y4rNaUWBNlLjGT5wlWd5DBzFtzFfGnSuhGvstUVHRgRVTHCsstssX10jGPBI
6qcQ/BXLnUbx4/uskFksrwUJbF9T1TVCOQk69L74v7IrNSpk/1ADsYpIjLpC
vRz30I4sjNe0wNzyG5NxP2kgHk//9jwnvm6H/d8HlOIkAnM4DMGchCkn12jg
v3hc7qMtzj2/9tIRLPqxyKh8fmkpsw8y3kEUREtGWgYlq3nOXoOr4ImTt1y6
g6dsn6SjXL8cJieyVxq9q82VQY1kibbjab62TF9Jk7ObdIi72D4Mp1uYnmMK
yohXxP3DQSUASIaxsg6cuSbPCR5jh89M6035EaaL6b3iSbAezmTng/AQER7B
Tyv2ge904qEv6AyyZ9lJht5wAYowUw03RV1LhGxONAk+YTWl2NCuEytBKyqK
1UF+L5ruuz4njONlm77AdrvWnt/EevWwBjWftdSUQOOpcc+fNYGFOFH24xB1
CnPYYeFkY+VOvWqylnei3KjW7S4ZenmxOThjrPEtnVt8NpmSc9nnCyRuOfRa
w8Uhc0uexfHgZ/6D1zAQ83u6qglF3bYthzIkr0GBm+W70sj88oS1JdwjI4Ev
3794USjEkcR57bM7rX/9vl6xgNPBsOs3kI2I/2NzNw885mol3ul7TDEDot6a
xFzEe8Mxcyuo/1R1SSdet9UQEifauf/lXvGrb2uO9q54m8210aCRtEWycfwt
JblVIFBYN7PGX0pGg0QdRkzF2/MgxAjdaSKUXR63SiGF+s73xvaSvGOOn4GX
w6YLptW5ce3mScHJ3/95+XcRuEY3XhTaDNh1sKecrSDsrKiG0znxIjqcBMLl
CxnEiKDR782ZeTvr4cA6swBfUhMX+3TaXFcSqxGMMpTbbNZ1MXOjmk9oCX0b
3Ky96Uw4t0iZkU8uWVwhUrIiOBg2rGaW8NpH6qSpi5bMhM715E69RJdf8o6T
ezRVoZrw8wP2OMhMYMDnaiY61xRf3A9BU4yVPuNJ0B2e2jw8t+CDHxl0Wfkg
2HlnWUAlon1iepmN7eIC8UPIy6H3oyNBk0aBcOcoctx5/ArWyNKWK5D+RJLD
eRVVoBMvRYKPa16tAbTCOjEUssMiYuwsQizUSh+EyqR3OyvJTy79LoxepmYP
ar1bMDHarFSJRsMqOwoUAYgPhl5xOUk9D38aHGvYgbsafw51cbShN+CpT5p5
ieLCOGdyydxO7JcYhq8OMW8/mESvc3o1Zti0hxclcfW742nvf+jJEY+hw7pR
/HkRJGsnyKE8O/unHC6fxilO9UzcZxBPQ5mJfFEbqp9dJAN9hkUjNTodWrgn
YvwVo5F1xIHUOzm/buuUH2ULhRehD/PPG9h4XpOxggMcm5mr74oVunpemSmc
lonsa/+wV0xVyKnncJJDdAInLQyJjuqXJUy6iDpi3ax6TJu27DJNu7Ag7ib3
6+D1qfRicV7cToSqBSx48DZ2dH2bQc8EahcIeOj5OtpN59Y0dvusLxjG4c9h
Z9PMmDkH4FgO5a+3Pi5x28wYNr0tiQjeJpuR1wV7228/ouimd3pAtwlmr8+4
JOLtekPEthc9lykFQby+nazzJGTbpZcZbDTcGCT5plfGU5ZlFtX++Zk2gMc2
XRTyR952wTUOcGTZvMy/FZYI/pSuBNBXzNDXT/ahSYM8y5yqGPhaWcR4TKyh
dIy7/x6iuFnxAZW6JSjsciosSDyzl+AovqG6GC/MsccMJ2ZSeBkCD7aQAuLs
1j3eaJh8Y6mfIOpZdqwBpHJ4n3oggUobYHTaEuDFZ1vvt+n551zwPBcwM4TR
ds3yWjW6+z66agtx+hphRbZj2jZ+R2J6QZbJv4rjeuudOTAKcSwyYFrywau4
q9QDaI+GA4j6VBMiVGRUmEzfKRN8inwFNb/ZSX0RFD4NpmzmFo/IRtRokbAH
HkQG2JGUXNV0kVSziQsuljJ2C3EgpXNd5p8zyLUXnzytDHCMMD2CVZyTXLnH
G4zqQau50AjoOFbfhxMoNkcwQuws4fLolM+M0nWkPE42Xk7Kfj3G7IQiF7hk
zu/86D8fVDo4x70xiVXZLqUb7A+JBluRK2Zo2YF43SqsW4YflImZlpriJ5A4
RV2bhER+XMuVeDHNZzl6SLi+u1n+/NgOSuguVtqCzfh2vLma4hSUF5aoaT6Q
bsctmzTMdly45ZsiHOOTUtC9gxWjiHhNOpWOrUs5iznuVrQ3/as68pdA+LCW
P8kGkx4pZ4folff+Fobwof7Z9w3zOqnShgYdu/g3ItXtZV0Nzu5HhoRrUayc
118q7vkoP2zIErN7cBqCO9oX9wLSDXpEVCux39drgK63jrYyPzhWDIHiRXo1
CsXTenLFuA6lcw8c4xpWFb7sbleFqCIF5vXI+srUJwba526sS1PsCumUHdLM
k1KqQLTAuJHXyoYYZNGll5q+i2T6cq1PIuPlyP1y2seR39s3bLsG8UeXOc1Q
UOjo6QdRJVqK3Uq6q22hyDr+tDsWly7P1Gt5GD6PVNaCmghByLVa90GS8i7f
87oPBWUT3Mco/E2XwAen8Jx6UYxp6IJISjGnt+wtTvt2xyHpMJgfPSwacbrg
x0HBG0dRGoI3uLOFAjIPMZEYTu7cLbNrNRcVq2yAKgHJLb2wUP970F3SEsZu
SqhJRrSOF45GYtycnUuGKU/KTI9YK+Q8y+2xhHA3sXBF8K16he91yN1v4glu
sS69v8n+n1c0xbbmMQ60f2A6BSnT+sVfon7ood+mMQNdXirSpPFXGCDK0n2e
Qwrb5Q9HySEYxJjkQVAlbXbjKEdSePWlXt+Ag12Cj9BJAIpOEH8NmT7s2nqZ
N+HN9K4R9Om3/sAZQZ/p2D5ZoeGRLeJDWFcLmKp2jjtTgyva3pYHP7RycWyv
svNbE1dsFZzrH81EfblWSSJIJbLk712O4nKmRc9U/oujiG9/7K0/jd267JC9
jsYbwP/P12vQbWJAr7GUQPrtD+BYpr8AKY3FahuMGcYzPdoXxJpb4ROc2eM3
IfD9pOQpuLd8XIYevuD3a7hkI+eM5K9QFbjMfC8aC5rwAAKITsdmDA/hWsD3
ywFtREmChZGOsUjm+JImQ4MrcrsLyXc4AXj3VGLzAsMmtr2oJwukJ4BZponk
CGVq9dYlNRNYkNofOZiIDVb/AG5grzCbD0bWQ9HAoYBT2KBAA40kP0Dy188+
QZu++ZGtJwMo+lFM3QfqC7yXqoyqnpVBKMs6VTJd4OwE2P9Ct2oH3PzIVSJ2
UzZw+tCSKLprnp+5QQ9CFLzOHJ4czbDH6awb3GiWR88Mc4z5KJDphJEWxPll
WtDA0IngTkUgueh2ZFsHNkjT8ECqwGphaB5FqvSMRtP4C002J2l45Ow2rdpG
CZkSmLdxf/me2eGsyT4HOB0NF/Dzi3dcXjqf6pCFmggEqihiWPN2E3UeLxSw
klEZEIrv31RXhApU+nY/gsRlcJMA0xwHdoRzd2d5L2J7V/Bo7lk/LjQw8zYq
lhW6pI2BC50v15UdUo2vjLBrdzMYOrc9PglIYxULKCuL+AZiM15uNf1tPuYx
lwVaXnEIhCoTKIe+ZkI9eqMq+IxqJQDsGVkweXh4UxuvW3Hr+hb1D7Ua/sF0
60Zs8TKqiWkeay0lYNGguSZdxIQVVWV1KB1WnVVru3DMb6WF9iNTL9nU0eay
5nwO2dG9PI0kYXN3x6fLd0w1Sz7/Lfa/AR1wRg1at2mWOBAQFK5sAOBM8stu
7aST3nr1+0iAACjEeeQJ9H88eESRWvHMy/EZmadf9S5VKa6V2iHe7OqqYun9
AyCGp4hTONWOqjxMVXyqbyoRAThNcy5ekY5j9ZtrDNx8YFo3ABGQPSHXuQk+
Dcs+At9nmrdeW9PIqKWP/W0bdfkUNoG0fEljSsLch/IO9OLiYQ/v1JXQwlme
AqfMvzZRq3m0PRxb5lJN+MNlIaWqVjTi4FkjHe576O9XcA4316wfHVG1BNme
ZKmvw4xjjArOCYuHkY5x2HwRZn71zZ9I0Cygz/bm9Xn8rPJiVuVa/+V28iwU
AenyUWIG7yoU67fq0BM8CFOr88avTIoJNrSNaQPcwiMYoUQiEiUG79HIByGf
iinQiBniFRaTWbnZVilH4GcjvUtKsOjYFzzIEpNRjHmlHi1uJpvvWYDBEF1/
bX4s+Ks1wWW4ffTLik6TY4pI8QoPtVUgTWvdnU7S2ht9tnm4AQkE2J1Eq0AB
WlpNNrTGenUsRpFqto3GIfYcZ516bqNcKKfvptJHT6e1fImS/pLHU3IdCt6z
X/kJcFKvBLKiQdlwkpelH7esW6+sv0UaObil+U440uWvpfSMUO8gjtFBK4DL
dd2CPk+M+u1nlgEm2y/u/9WwP2zqE/m1oKkuJ1t/dkLbVoNjt4D8m/3NDol+
agM3LvUYhbH08yVXmyeoRZF7xjd1Rvx0DLevvhaA0eWruOXV7OuSacA+Q3Vf
2Q3/TinW3KA9BJhdz30cPQFkFlTufVXqE0SgiCrJ7KcQGSN33n+xelul5nT/
TeVj8eO71RjeD6s2yegVFyGZONI2RSH82oINCVp1ANeNhftSe+jbv6BlhNd2
/cltTk16m2JXVZA/25wIYx51oHrxF8Ug+RnP0IvTsOfl/Pb1mHdcJobn/9JI
zFVEqdyknU2qm/gBdYtSLs5AvhuZXAV+Baih+G3KrsObp9h2ayiAAjH9HGrZ
LWoxEu6NwjL2UMV2QibEURqVLmM+U/+DgrLEO//gvFLmAXcpkvrnfXzmFo+D
oHVekTjLPWGF3hDaYnTNAf6VIYO7H6DPCAYS+XinxURIW+lrfCNDb0gasL8B
vjDkpvIPFICJVLBcoMrJz/ZuqJrBpb74SfgseznIQ++XM/HBB1NxjJGDK6PX
jxOcsw/FBYZE2vXF62MOq/2ThH2qgjV08tZA/6pjh0PJPLzVNPVTtqvi4iG0
yQnQOVPyzzWm6ToOCRcrH2jAEh47gJQxw3WFqWCyNZgXjOKCcAi3AH48DWFG
eNycqJ4MX350n3cfJhP71qFT4UMdsNugUBc0nM1U8TOtyzwMHFOVl4m6tjfC
3BcG16XiOT9BKbSRCCYp4HPK7ph+12kZ3Hz4GnwbVrmSy4ZUvlMUzZsQWwe0
6ZuVdx1g6kXTOuJfvhJdGDwRBkSl9GdNxIXVCyEhmPvWMwTZ/jl+kzsXoSRv
8fHh5jCWHN2zJwTJTeCTKZBrgg3MpE30xEDH1RdEAto838hA6ScL4eQZt0W3
ibkFBiJ4PMS+HFLNSlRhmNMGHaarJhhIrFNXfsEVIBFGh2L7x+EpRJBdFbXp
hbXHd2AGGCykavM5QVSBqUzexwZk1+HChb3RHz5oeSgwV0vto3AQ3VcJHBvF
lJLw1lXvGNQ2cdDDY02Idy8T5rfMINI3NeaJv5eoeQ0TRG+Bd5rIJ4Wf8LeK
9sRy82mJjIFsqRGZxfhUljSAD5wH5Yb8BQ+ihwvBBLz+mJDVH/Ol8Irs8hO/
luB5dECyrVcZn8HqiuJhBWU0U32xuKBczlyMRgQOPSOaNAGaWfONJhwtSLHl
x2OTcTrdUJ3zilUjJ5naY8tnxghPWlRnVH37cGuSRsklfFGfEfDqadehH8+E
Vrp3PedNxDY+M8zdB7UjDWHphhm1sPyHxDFRj4vSzjQJy823hM1uhSdczO8N
+KuTSjYF6F0F5+H9mAqN2NxRc1rUaImLypDoI8IfHKo8/aFOpWMX6H3bhcp/
VgUhquAhawAVDABpo9RZ9cvXi/AB6W/79ufya2MtwmeI3pEbT2x9y/m6BQUP
BV+2KTcA36mUzqyj/EixFdj8SZsnye4vtWNrGDvsmrkiikcwZYcMQN+oQIOc
BzX69hq6DWyDa35EaqGisH6jlLbx7ji+cAQPuvqXy61uT74e3Ip+m/dSLpTf
nMGhiidOWzF9jDe8bExYo3aBoLwiCt28WSlGNC79TnqOlZmV9gfpRZF9qhJw
mNawux8FNROhNHCtqbGopKn9A+rcngrqStLufVl3x2Ur+qVlpvknoJ3fTs6W
DneJITUMh/S65aBMlDTAqmlJCT2ujsgS2NJhcSpYYYk4aJPI72UwPPfYIOYf
SK2pafz89Yhd+LJ5lEKRI7ox2vH5PbaJB7zt/7Ua+59fWbNMVy27qLPKVtRP
OHw1Ew5gtt6xhwMz4MZKBdQeqgQNtHdOFwO5DcgFaFNCTvBjf3Zj0hiiOvMA
g97hFeaLPbwTuE2ODkHEjEphJzIHXEBYQPAG+ASL/0WRPt5XUA5N8dhS9lQ5
hfkhCVnkQoSOX6QKnAUME68NIxR+yuB8xGDUTEHYMOj1z9tfa3c9+/01lN5p
A/rPl9DdJDdgLiHnAF9/MpmMVfpb9jxL6KRRa62yxD/D5U/uvX/Wn1B920zW
Lb6MFEqjQEsoiC12sVazi3BBYAstZMjNyyWDO55obpIA/Z+94Wh1LcslE1XA
/YpioWWNPpe2ypWbtlEGdxe22Io+6VkyZ0hpu5HV9AbNvannEmjeQJ+EtmFl
IUAJatPiVLRA8ZBjHxZ62dYS9+o56T3FagsNExFxcOvh55Lg7haR9xKdFy7I
x25A37E+sSCYmpmvn3ofUvVG50+ZdngljKu17Oso7g6XyVVzk4XTIO2c27NE
thhIEM5H1GS2323wCawMfi1YATMsTTX11Uuvdwmqs5XBxSHLtD9GppX5Sx1O
vB184VVfandE5BThgjEY5bWkSWDTZJxLWh7S+IE/7QB3b1GrhVBGHJ+Haf6z
mUBEKB+7K2xlawYmmdn5egfkzJjo0U1B9j1udJRj6DtK/ViesQ5EzGU5L1zG
79PjYs81Z24QegJDgcxcqhX4M3M6Cbec3wM63W0dbOkHhD3JNragowo4sDTL
zt3NvEz8MhpELTANpaliqTW2Kt6j4aDjC0sj+jG9fG1KJkLT1kisFWftaHon
HWckkalXyvHu2ikK7aKvbiJusbC6bsyKEIMEJVD4smvWo18b4OCk87I2L+6U
V9xqCOMpsQGLpr6b1sWk2KAH+S7GvS7UOb1FaN+pgV/kdz0SCzguZn3NUxE8
hrhPAtrQyujNGAkvDSyXNqICdxAaI7xLck41UGYNhP6lbVXnE8DdyZENjNuq
+uZLx7MocE2n9gCjjvLJQDNgwSWz5G1lhK11BRT3RYnJr8nJSBAaiKHV2DJ6
tPTB/pFYIdZOHj1RfUm5XlEspipDUKwnQUp5Inm6b+FiQnjWyx12jEgIkXB1
VSCmFhniCaCdGssOmLh79dbob6ZQt+BxcjxnSXxw5Z2fMjVFfjFwusRQduWe
o8xoovX/pz1hSK9vSPdtKx+kVzmgrionaGleHtZwF+OjkoC1+AiT2KxUgu6O
0iu/sS9rb2qm71H8MnVEeL8ZhwMoP056Dnb/zqpaKVo3to6T5C6yR24rr2vh
hjgBIuVM7MVfgPPHRwW1IHbhKg+ijsmqTlW99I8KF2svqO4C//KnVQCNP8aI
0jyY4QUoY1LN6x4D8LKZflJgxuyR7/GigNkjiFtRCfqlts4n2YkTbPNBU5RZ
BtLt7Mr9hwdoom+KbpBSCOjkyB9rh1NRaEZaufGmWYsMTI2VoI0orFEZg5TB
qAT89s4AuDqaGelWgy+Lp6eMobfryUevAXuFQpe295stfm7W41Hj/GSdRG8F
irEp3GcsvbPVVikjwGnWCA9AkF8qBFiBmtbxFHgZTC0bHzp0+NsA3aaxpRYH
nh7WH/SdmQ5v12Hk/eUR1kK0FfZPCoB7bWVo1psRt4bpjHxm3TMKLwTNHrWc
CzFynAPN+IWBdOAPd56V2eDG+It8WVZMdulnEAW+aZcNiEl/s2NKATCHU0qr
kWwUaLLgRQI4n5je1sW9xaFbmDpynrijAspkk4JckPoOVZmZMswSPatke1k6
MJcOyELjYZcW7x+ucP8hvKJ5wD9228hjtoB1aq6Fr4dYCwW75mQypo5ro5Zu
BDXhaxMPKT7vpYezeHzkszuxnxkTHq3RMKceWH6m/NIktZok/DKEosG7Jp/v
q1To/qpI+qpZ6vwDlPl5lyG9ew5XO1sBD8nZ+VW3sBl1+GiuQk3YkgRKq+XE
lcUPouJ2j+l7SqlR+UaJLxqnfc83shhS0GNxboxlKieLAm4Xvop+cnRgSpPP
m7kitT8pWKbBuVVkeoc2eAgRppmra+8i8iMlcJt+qnOYovJO1ga1itYS4WkS
eqcDQ8PN3779LAC25KdNeKjJvbHX09JVqn9vNZLyi1oLKLe3k1mjC35FFSZl
KbW8fKHpmSB83KQZRUHdW4n8sdnEypNsy0S6cKW1QZoFdtCf+ryPiD1LPxts
uQOBo/ozLce8RDQxvnVsO1BdDHeXTPyICWkw+M0DhnACOiOTdCaAuXq4Mb32
hOeRo/BOHxUfngEIvXM02+5+z1YHlHAakis82kYm1pRpRWcbcS7Qst4nj9IG
Urd3hkkCy0IcZbelXPxLxpkDwW/GXCFb5ikHdvXS84Hmvql35nxzdFKk/PDR
FiiNyx01VXAeWe+Ko8UCrJzJVocBJpSZ5Y0sGKxHXdTcgwpNW9Si66Ga4vjS
kM2gR0QxemBvYI62OyVtVU6OjdGWAUY99vjdY0ggXYwoK2NpqkVoo3xkxKB+
z0QrdytMphuqN+MuiNbf5Y9NOIUvmv2oebsnfCcSkRnq+B1vBY3/8a6iQgnR
mfZ0pCtLm9CnmDmRHnDixEs7aOnqu4iTxWmMcvhY7yHnXmnMaw/NhUHUMnlK
HvTiaiL+qLUXg1NvxiupUdKzu9c+Y6Dl3n7bj0gfEd9vKgiqC7lPM2k/TtZy
QzfDQUIq4WUVrx50ONFV9RDfepPxbk+5y7WLFIZyAsEdHokk1T3lO0EbmnC5
cvk8HO0+CaVrqVvLUTNq9O+9YZgMk3zx2kXiWeOqJnBlquEx3R0XYW/q0opn
7AoZ6kyPHxWyjjXfxmzx/6uWVfYSjRm5gy4X4e42d2etI3imQdg4ZH9cl50j
+SB9XRtGk0UHxrT1Ud+DTlJ2NePj5eCcIa6FjwzR7jrn3hja5jtyO1o21+Gi
rYlnVw7uEeONYiIVVQURJ04PsWc1CwcaulJlfBLPP18fKJieHjVk6OrpEO9Y
bKnRvNnIsbtUv1R2MQZl0KGJ9VR/HaSI0OU9kTw15aY68yyrzclWYV15krK7
bCATXUPPNXRmmQ3ulwZRsOwvYc8+s1Azul7UE8NPMy6Xk+CElPBRhxS4Pm3j
NwX2s77IiqqN9klwV1aw4fUdty9Vw5VDMgyQwU4VNu5RtySSlyFfXKdVrO27
GUiYSfix7ZIAIqTNyKewzUGl48s7JNQaz9yq2GZLSmTAS9uoXfTjtIf7EZgf
Qh0B5nC7W/tkG8qoFSvylHJkiCUxu5Dpcswk5A1yd6lhD1mh5HtZeoxB4lYk
qKxHO3tY9iFnL8J6AqXl/+zNqY8GODR1BkExFfyjbFE3dDV5xZ+yZjmGFiQm
saKLoexyoV4c9Vys51Allie1KVk8nkn07CThTQTCshxOK7xRQuWlL9o7EaEp
P5zHBtDxtRIlD7ExcTO3eJePfyK3Mopv/xoVWX5uKg03Ju/P/M+Oct10qnpH
kb6MeYg5s8x5k/wZgQhuNIfWbRFkunjDLVaWnABH886VA+Y18wOgxdxeS0RL
s5BCCiSUHquWJlZ4kElaup8CY28XzHilpPf421Gjf9kOOaX6gWuNRTGJOevk
PNFN4KtbgYQJ2RtRq6ty38Dxr9Gkp2sGEKmWvFCF0Rh9JpEEfwv3R65nZIn1
+xNR4MX25Du0KyM16ap4r2JjlP8TMm5sy9Z5xkUxyXvaxKVq2dt3BsfsaMjq
YfDuwWoqnJzx4mHmCAoucSx551Sf1MXthvgIEDr9dzbdA4TTariErQ2uEyFy
oVSKpugC4I5+eq/z04o+EYGM/QySjAlKIdPWrXaG+XN2cGKSOonsxZkd35jE
PK+pxsO5BkZTyehecrdv7p+JUzYWUdCneFVmyMzcJyosD/rhOQfRKPcfLRbE
9fPmdvSKCCw85fCf1lwSJINY9HsyMVUibY88qlOOWgxFnWNLa8BXcrYFd49/
GFaNFbeYQXg392x87/XMX/vMsWV/MXnnobLz4rgobR1gqPPjUGuCfeEAsbGq
DAb3/qDiZXzli4y8aNHQUfjAquuFbo40lVJdzFRnNCmvxuWW+60YOTrhbr7G
vgTMK0vHdfvoTbHsnJvOBthcDR5F52y+oycrqX7Z9EnH/cB3oorudKQ1nG+G
DISQEqpn/c8CJ1NbvFF+NhAR9QiFz7bvOzUqn1+s37XycjAKVhxCmunRKFzH
x6gc6fOwcMhGa6b+/DbhDCj94rgkoGAsHPRviBlqSif68S7dAFK5d5shd6Lu
1FTyNjAcVu7gKNu4U33qtIYgyL3RkXcBTGzjWx6lPEiJ0QtCImGCfNozuEwk
kQiEDk7ZxjPDCO0ndPGv+d1/JjvN0f1EOACQTDolO5H4Esq0ReZF0kQUWiM2
bINTs8W2/iWr2JBeY9HJ7nIOFC4Y3KpFIYspkppipkvTlD3pU1w4ig1L+wj1
h7uBGlm7SG/hYMZT7diwXPmCFune9aGgstFtzCDsOloKXyEKK3ULGfm5uNK+
0Off/NwT5VbdqaG2dxTc7qWemDnAcSgKRsPlSex+kaQEL9N5U8Trf9iTZvn3
hFQ=

`pragma protect end_protected
