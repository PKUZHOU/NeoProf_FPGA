// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
AsXMJyfmtnVHALWKdUKaoO1GcvyLJomZMQONj+HtyHO2bGeBsxSXyh4yQDV+0uZz
WofWAuiZqGWw9wD0eRX5cyfx1FdPrJvSz0ztdeQlbgCp/v+K9R8o2qlxjc/XtRcE
hmBc8TzY68HiH559gMjoRAyIgANWLMY7AxjJ51bLh8M=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 1012928 )
`pragma protect data_block
Z15lZmDTyWZKvbFxD5rfMLHeKxSFhM/KevLz0oDNvUFrUm3BCK6gjUu0h1JOYmOs
x/i8P9MYlP8zy+tOUVL+K5YrXRpxRAyIAVtkXZPVVOm4ajbMPFqBY80mF5uKziXB
hzvFctmgobzD4YyqcIkgAGaMPjhJ0GiXI7m18gfs/Do7SIJEry+EDQL6RJCGE1S1
Pmrupa3RqA4ifZ9KmqAcwisGJzicHlqddgxFR0Oqna7KXJxVYGHHBv3l7NPVu+IT
M4Ga6givcHuSmGiG/i3U4yBY2P/VD/cnTDxKd0jwxobMncs8kQKDeu0Olo7F+UPP
GD5ffifaQOO8IcdPg+bSNWyj6Jjq/mL5EXwmkCiEyRWfrNoxGa7g6wnEML+Vxyxq
JXUgmSlkgt+v/mlCRBZQdefzBseAzPDryx+MkQwsj6YtcQNqa+5eRpoZVLVa1FOt
yrXmmPaWYdBYZMgA1yUNo2RElmR+l5SMQmqIGMOBijxhaYf64CqA7Hm+AWjGD+ur
JN7xGVFifv1tqpYhbs4p+yEeD5X/2CXgI33kGz4Xhomc0eDJfl3FFETyCB9rp4Td
Q3Ct9fGHK8+bvvcmCm3V3/hoq+2NHFZXsSdh90aqWyq+VAjsr78AzHDHuEx8mA1a
8xpRDjb/RXCn1mqJVAo0Bx6iIA3a5GSrH42DRSizBIpbzhzq+jmt+E9ljt3O13fd
T82V9eX4xbJ3cMOxXzrZ+mgX5LGLlpq7m+koEcXFow2bnlOTPo4jOnyjhdHdR3IO
Bd/ZEJHTfrNX0ZM5ClleBIzTmnDd7seFm+1OnYBCHBw59/PxaNNRTCGUQ8LURH5m
VzFfiJlzbNc9oEHLmeCJFqmMvJkNCiY3ILvQOhNSAUCRDQ6IJAafkAo0c6UW6574
mWS9dyBcRTajeFlOiRyzuEnIk2/4d9Z6SASx0jphQTtaReRPxFk5WdRn6o9thZzp
5U/dPoICqn/RDsXg5vm87+6gQ5UUwMPIve8S8U1zrNpC97qZFzJsFy57ROMxemAD
wZ2kmk0kOYShwa3HsBnWcVGa/0AjfP/FYjIS8LQARxCJSKn6G0ZPmLOHnNJSt9Sc
ya9DtV4ZohPUepUzbY32l0AGtS5OjBovQM3umZ215t+4xixpgnUlXQ1KcqJGkxZ+
Pah72jbavglOS1XqtC5C9RRKdPzl+9ARGtwF0MDfWRFfvH+NaKhHuQjZJH5WzYKs
5qSHeUVO67/m3JwFlZwsaX2xNSfpi7+5dk01GEov3YOFamDyvC8zGDpa/7R6E9yE
9GXOEjlbY0ZRqNnXjWvEdEDdqJNfPflnlf/bPZsPaQy3wAhflLLLy/W7h3ZcgZDm
zvn+jBETkEB7d2OXVGPcAbF+yLXRzFjtBJdabh8zPNNcKSUDwjlaG2QT367V48WC
HTJOik+Z7luIhm24zNsQ86VGVACCU7aFa40PMLvq4ymJqcHmiHmhoTetDkCX3YN7
Lx2lCP1G8RuXhw0XqTK3X4LgklTVMtLz5T0flb+AgxlLCSaku9uFLBFS4ShRkQ78
JoDO0EBmkEG/W4hfWqdCNyKHqRSpDliMXhVJh6fMhXTh7I2CEmhZsPUecUBPlLBD
Um8G1LrNVN9P32Iov79xwep+gMqcsXUOiAsBXE2odaK3j0bdOGlwT7RjFh16bD6G
goED10l/mE7TRFQzY+wAzmcqvCv2U8MX9SZIBAvDw6miY/VW3muBZplMT252WFWF
ODv+85qfGbiICNX86noCq4HLZaQX20gPHh7gdA+IijcxZArRQSj42OwaFjmSwZ3M
H8S7pYcjJqC5k+TIdDmYggVHf0fpqKaKNNE7f0EB+YJPQow2sVdxpKKCHgLQu+XC
K/WrNT5e3p4nK2a8vnkitxpDyzZckxAgnP5e9mzbW21UwqPHix590n6VYDBhvnio
uxpQrmp0raWBQ64gFurrxs91xbyUEW2/KKQK5SKjUor3U4pEZpiIlzzg3ImyvvE+
TjlmfCCTxqs+kpxkoCUA9P4+EOu0yuPjNRbpQfbRp/bXgjYC+n30+fNcw9UACyNL
feNM3/mUmWvVmPyYbdgUT16T6fWc1rrnSsqcsRx8Od1H3gjSANWWnJJfIIY3kBPx
33ZRQS8WIci1+vjQREEB6MIAw5oFsDbENDWbcITUzK3RX2gbwvjcf7apS0kUuacj
wAyxBI5ZL9Am7vSrjSXeps0KU5pPQlnpZLa2XN2TalAvEBuqaGMWlJqRx1+owF9V
FubU3Td4ddLrU/GCvYk/4523VPn0JqecL2yY18aZCugss4Fa9/3c2udPNx7mxJcm
ub0xhyWEo5XJ4WxiBD/fpdi5ROefsDPI4S4QidSdiJGdeJXYWfw2pSp/Lhm9BJ7w
dHG4SKoEHB/QmfQk7t8GUqHQNX1/Uxu8c0B0Ud9IRRboj3JGd/RhfXg6aqg+gos2
Vn57fVWFYIF+EbdHYZbWSU/qhJ+KYPKCVyDHQX2VjkiOau9ztSdvSrESNNqPluVU
mdExg8I2GmWc2OdhszfE4v8LgHeNDr7Zp2FXx6ILUw1moUEp2NIG/lvjG8DCHH9P
yqeOlKoEccNYXUKWE06KaDS65mef3Veqj2+VP8LF8uBvVhdxvxw1H1aBc7Tr92wc
h5Rkfb+u1PWfBVxFDuhKHK+JOgH06AdOZ3+vIPhJpbl69P1yXe3DtoWCE+eOYsqt
iwr5888rJ1AblnycsBopIQ9Gti9T/foYT+E1DBAaBr1Rtv1b3OUiBzVTjtw51xPj
QMD438Ht7vrC63poxU8syPgyobqXAMThc1i14rp5eOnh+jKELa7H6QXyHmr8cd5g
ebiVw0SGfowUsQ81VTREhHgeuZUXXdrUhELkRj3UT3eZQS+XT9TPFS/ssf4JPP2v
eZ9tJZ/Va/KsktcjqbJX+TFZFfD5hhrtMrmF5hUgawqMgma7Xu2+VRx+T29egr9N
Hbco7yPhPzVULG6Apl4Q9HrAR4nBGwSLIEevNTQl2Rg8aYrl4gzp7C7YJ9m3CwR6
TFgINS1vu8D3ssHUpPwU5abUYcaObdQ+x+SsvuBRH0Cn6JiDR2c6XqstApHNbJVN
1AYU9JbIyrM00KEP+g6gBNuNd363LGgqIXT9HKHaBHq5GINZNMgVSITbcWBxoPPm
5mzILmfMaLvRBtBYh5zkI3cTORc9yyrOO+kkNPP7dJYBtOtFNDOxElrX+yIdt2TC
ZTI6rHEoQ6/qPn/Q5F7UrDBnti5RLA8PPBD6xYsGE3FBQX4cpc/yUqjLpM3HO11y
T8ijKbEZhRBcvkmYv410SmPdFtqDj54ILt9kvkvDbVR8MxKwcdP/hKWltYtQCt9t
hnUb0gYDpn5KyDphiVkOStivVfAxousZtC67W1baXXl9XBhCfhKbk7JzMxeLpHor
CxZ/QTcs26fwrOfotA5Y6bJ8xFLcU7Cfww91jXurHboNDW7g7JDd7Sv/sn0jTwa3
kidb3hC1stD7A+sOzJnR9GK/00q8lo5EYOyVBYMU6/jt8Q25kX14M2kkdLbjt3Qq
BtSoFBwTFezAzf5M7oj7aOR1bLK/kcUR/aqT2sbq3G91bLbi9Io89FUtEvMa45bR
FuYuISEirJs2C1S+pWyzgxYxF5/8V6iVSyuBaT/Ie/HdUhdykSpvmL4s5byqBwj5
JH/7VqnBFElNUi2ZPILtylIoM3NRQ347kCLv4MvCNg+eOr+9NNVF1xhU3+7m7rf+
qL715XPwqGUloMyJF/Cv249CIAYQogVZeXh+g83jBm06OMatSP+1Zyxyz7tZkBlf
Y2UfLTlP78Yv+OSLc3Tsqczwd+4oIJm3iPOKgR7x24wglSg5BD43x+pdjbjodTfO
BXUAaVp+S/IJSx7lspngW7SqrNnkAF8COw5nwMiSaYWQ/IS9TG805JCnDmroK8X+
KJhoTy2hj1lwleKKjH8Pf512KDmd/o7dck2kuVjvc8a1s1jhTl+bCkAcgF6aQilg
7R0i4QyhAbfzNOpFBBL7mkPJ4o5X49zIGPRdyVlipHIUHf/RGu6bm0vqvnXzVzxv
VX9tsgH8A2E+bjLomz2wYlzHg5pgfFtLke7ROfiKkxH8ag36n4tV5Bjt/LmwTC+/
DZ9e/6O9TVb2UWKUq6g0vwzFTpYvDPYAnH8pUpmeoyZEshX9miZgMy9QaAtwOI8D
GcKw0fEpliVlwaMoMIgEv8wni2aYpbfsy0ehVp0uNZnXeUO7t3PJDPjkQnjomzJf
LgejfGTZZX/803r6uECICSzwKywkVrKQAlExYmZpmd0+3jc/Ih2IqAlnoXmWnCfA
+i/6C8HZhsWq3ECHZmvRy31/HcsOV8mJtPMnjygstXyfIaaB195yToSLC86wBKPo
fIpYPQ0fgIb42vsNwGJVDa2wgP9ygS+8mPg8Sq6zd+V5TIRKZzWr8OGmOsQtSL5O
OP4AChGNn+F5LmBwfku4DXui6/eLm4+PqP72Tf+cl5XAQMJG1i3vcbMKunKH7izh
4/sCzZ12kA5BNgOLvOHwtuojYfaX3R9PYuRFPhECW8zAnw1nxiiKFlhlfaQnwY5z
275qYl7etWrGnwIlloEPZnWSbzvgLgLMuGtdUvswgikD7ORS9L6Q2PkpqdXscY7i
O2mC8vk0Nfy7k56QFErgYIhPdZ3h/98s5SmB7dr0Kapr9QoNe38/7gWVRMK+KzQ9
tWam9fPyWBrFDPPBjuo7TDJSCHohG5oInGbVcvfPyLS6kfUGljl/BJMlwrgdqNek
uEFPQ0RxahHw/sf7zdn/F7zkcwgVlQ3YyHleknm1Pezcoau+QSBlG9BvC7MDCay2
r8+BavNBZldFGM5vt4WBEkYB9l+71Odx2h+DHxxCRtYT8qYkuGcSLEWMJ3qYBCJs
Db0Nz995k1ZUWGkmVweu2Ef+CKZEnFLnd//GVmKfpDeCMvnBrdGOdNRr1ay3PEly
hpaOnexhAwxDa6r5FY9TQB3EjQK34h25is4Jy69C3aNIU4dSHMNoJoEuTx9jMuKM
XsBQMdgKbtlGyaww3FkS8lY2nyTQ78onGX6xxkPfAmW5fLrznO0UzUkVLRn+e43E
fj8Ja6ujh/ipNZfhFJ597+wJCvuax/thjmO9ZifbqN8A/P/vyLiZ8fZicVcIF4sZ
1g28PgeJFZ6iEYBIhGcJnnGd0qpEoE6bssc0uV3lopfSy03eh6/W4OEo7eq14RfF
xd9FG2LEmS0UvQVx9guC1Juav1qLAPDpRdsEdOBiglJcq14rKpvbKWEcRsDt//nw
+DJ+PhVH/H3k0b/kAdsjF3x1uTKUYVWfiIfgS7iYd1L0sJy7v21k6Q+aW3/mJ+34
lFNvcly1o5t35q/UailthPpD5UKzO2K51v6LQnIXijjX0YUMSKotEvupCQ23E15J
1I/O5f7lgQmLoqbYVLOHpk8Bn1UNDoHd4hqTTtuGPQvPIVN4h65zLZ8O76L8U45b
eiqQsDAd8zoyyZJ5GAeJ09jlJRqOukcP9oAw/PlDBWZ/z7fPAYnrDHTwnwrFtQqO
aDklwKZCGCVbHvkEz+nkfR/LeGsjZL7f+9pc99BBXcJPtlJ5+vYRbfdcat7tWmQH
+0Htzxl+I8LJEX8Ttp6ZYISKJpKKUaCsfeYWTlq2GgMLjVazBMbjZWP6tvvwzrgj
RAgRmuabau5Ak792CuW++3L+/XX+370GJvhG+SlsGBf4QZLfJbN33jUJEJxRsWIp
vW5YSp8LSIO8qq4LT7gkxUyzU0kugoxRZR58lV6iIxDuvUloej0hccxwRrpUDBoV
Mf173OPgq1gDoPXWSBdeVq5EF+qkQHKXpcxxLHvS2vOVcpH5KgkqUGuW/pk0frCA
CceoXcHjwJOFT1JDWNgyDAxxB2UGsgciVcCKV6SMYpNVLVJMya1KOkypMwinfdov
1CRnSRkPOovnPhvhRZFvBCewcN0WxZ8UIwMRkEbfJBDbEwSdANjsPPhwXUJFcKvq
pQEV2CUXJhYch1uc/UTNWqQqjCc3eYtp5D1KTat7cx1rxSgljJu8wNGHvH+RvAJY
8XFVNxSv/vt3gir0hxvC51PZAyNCclgGlBnd0X29wkpXjd0fnGFtQogtnS7O7STe
D3coKnkP3bNYRM3nZI9pP1FxMCH1YY11VU1IMKILoq07rfJxtNytzCeaM+ldXpZj
cuDdJ2zj4Myh4B1+DH6eHLSUc6u+mkA/dN9CiYaRmkw3pMcnx6QzvIkJlVYdqzgX
aGLxDFmb4I3gqUaF+atKOGoKJTASNdSpgmU9d7DO4f5HJyiweoSFdMbum+RlAEaB
e8ZlKLSaUeb734Nxp0wOBAie9yf6PLN/qZp5Q6bZlKTMR1X81eY6Me1lkTncgxWA
+c2G70oRHoP3buS5+6rP61uSeiTtCULvZG4agxgbk2a+2RerTLMqCBuuha3d8c1O
3mb+v5me3VTOlDB4fSWPSEfI3mrWt0H16MITNOc8BaWI1VjtowVm8jTm1va/qiCc
W5my7rmyZlaQRVc3hWWdnHXRQe9Q2pQWrRlPXxDxdn4Ra/nulQ0otWikBwCnUgi+
ZWr24fFplOvbVFhcjVIvvnCjJ+fdkvGNuL+p9Rsw/PdPT5DkuBdf6MovXh8Tx1aa
lEq41xL4JGyAqglsR2i/pXyEPm9pYpGpQM+ua8B9uX2Simp/598g0gY30oGH/4bH
6bj0a0sXOJoTvrucKtGaROc6uZjAg9ZpP7YtR/ijY7vH7MooLWFpbG4jdfU7CNKI
kkfBwTbkaQeT128SQM76JNpxBsAmh0LwiT5Cs/4Zh09rJIs8ebaxyHqkXd/bkjKT
xIpc/QNcPOmfleXJbP5iOdyayjKh8zQOfZk9evTgUFFSv+LmFU9DRGwdtxsImKvT
Po5aIIRlnlYBrFUaqFWTOu6Aq4VEdr0v+lk4LO1Lq4Q4e9sELTvZaOgomoPwKiQm
KTG6YR9L5u3gv6n0NBFyLFaS6i6RK8CQnvPwFGJmI2RJ7pvjD2Y8fHTlox+gKmwG
lfUvnhzDOd/iFDuN0+fyIAPmjqF+xDQvUTRBTe65vKV7B4FgpDirLnECBX3Rp4Wv
DHV5Qmky7gNtij/Acn+WdvxT0NL8ND6FS1ybaGVzXn3lGQpR8GhON2ZfYv4gVPiR
XKpFp6tcIdOSZ4/yGMdopyUsjNroJpMVRWZuc9YeoeR+7LG1ynKVqBa9eF2bmyHz
chN+XfFgCPI9eIaTQ6/jq1jHs/kC3cgoJk0S7OIWYoxhiSZ+Uk6o2cXHwGpldXko
5J4pAdGqpQmdoqrDrTfQRzsaH5fV/3RVjus6lpPWO0eQfCCTFBE/mLSrSC3J4sf9
kLYyYxNDfvLvUbq5EDcNOlu6a1wl6eEGBEKcaIT+Sj/lsalgrVl/eH0bzQM1Tstk
zTuosYnE61TIZcjR7b2BCkAOcuVtmRyzA2pT113NXy2TPQseEQLhRSJQL8cMizMn
54Yps8zwOYE9zgqUvL5ObhyBC5bKCDOftDiyvTTnKXOLo4glmMNt3XCZAoSGvk+y
919/s7RKTRMyYsdAg4OxuS59fJTUdRENokpSPXM9AsWONZg4zrvED8WeBo+aDRyV
0xD3oEucNHwdz8Cmamb3T9Qe7SLvoHdKnaGyk7QC7KDm3ewSYH/w+iIAX7Bz1Ot8
cparseO00iKtpD8LFwLM4pb5r/tLlQLJUpuvShbbQ4C0CwPUau38+9QWsJoblcro
tULhYQ1KpIWlZ02gg8uRf5/q2sG9SuX/Kg95uH1JB5ykvhNmB+AZ2w0NMEbZJaCE
Asza6KzLoasSd4FdrmZ2wViQEZHTet7ZucFoRUxv3G0FlEAyh2CbZ0Ff0iBFYxNG
z8TDzVtoad63c5H7UN8oRNjmo/bvrOWUs28/9q0iU3HkueWkBuvWpFwa6/tvQqwR
fg9uPFPZOUMYfCVWgrI5Ue4LHXmsvjf9Ggkljz9EQSrIqhA3Z1TWpeYwtm6ijBwS
q2B7yu9E93vAj64Q1U8Z1htb432NGrTyvtwbacd0Q3MH2Rg1UTtAkBvJzw7OYLTA
HgSdieuecHPxhni1X2ttzAuWCks7h1QzYYZVu43pGl1hUiY3Cch/ATC74VCzicQy
SuGwt6rrnGPSXLH8A9f+xDRQmeXdWYseDRcUYiV1QKfgOuiMh3aKZ4IpIKtoQ4/0
93CXT21e5znYgJjTBU6ZXpRSHaX0JMRiN7QBP0hdkcx+WMHlmQzriOG9Ontnw4/J
eqypsIeT0826h9meH3CQqY/aDdP3Xuqw6sEgoIacnYWT/QWHVIOyJdKtDhek9t0R
uh7Ey2g/9Esr+PV4n1w0m5S0f+1PF/bsBvi/di7smNbd0RcVCDkuabvqaEXS2/oY
sXIImaE1ipXfTcdCI9RpkxlreG45oyZ4LLl3xsskdj+UgERLo9epdCzbl5tA/AGj
qW0IQNohioFN7cjVu0n1/2b+Yg7N4QVJTnYFlEpw7VTjQvx/qn3TiU4UeTwADfTB
r09r418+X8nohsVXQiGdnKY9Y+nmziF2XS5T11hugq7V4/qpqUoCpqes5kwQhPTW
klZrBloKhVR9NISgQJObn7wOqC8ydTOl4I3KM8ZPNxu/IKjQHK1MOyjNIyJaUHkY
px+Z2gjvY/YPAVpgebdJqv8YcG/DoC6ALKpvHykPtHXoDV6WMMPKVTEbR+5KxSO9
dwQIYzkaSvACaL/oPJ8ERiJB7MS1LXl0bLEu0gcCQdA8eFpw+WhCYf0GJFaUz38F
kVLWIT8SvsonGCfMS+cZRyICvHsprDwC4ixQ2cEqN/SNtd+xwzhYoRbCqze7SymE
3vpY36Oyb28wykLFbuAEcZwllcbGCpDtDcjnmtAWjLOpe18FkjptoiPm1IbKIQnw
d0HZ98Bj4kRtNOypx03GH/X91faxdGeddSwwTHIa3ctqjxvbKs2l4Xzp93KVWb8a
D0lPSr2eZVK6Aok9qhdmXx8UUyD7WQ5hKt3ONM5O5hYQvMMmGIwtKMx00pujGLKE
goasqL8VlvFpcOEHfSHdHxHPxuvam0/EoUHdHZcnku3VCcyMvd/2LyTz6ZR+yCfq
xeoS9M3WgJ3SXNVaIyO2tF+3H9sFRAtNuYMx+GsGQPdhHRBtjlbm64TdOXKZANX4
4tdkKRvFuVI6Gpn338jvzvsDVcUcJqdl9EZOXuyXZ3SQj2ZDjdCGXAviRrZLmcoM
kJEC6VpQWrmIufGj/+UkE+bGHcoPOqNAyhPkvU0QEdoQhfFKCR1JuSflKZwQKRAF
tQI9W7GPUZ0uc0MpHj5st0lu7g07SfYP9L7xPJ+0VsjmIP5zuwNSV3HpSVtmaviU
XmlGEEH2X6u9I81J/aNl6ps++4OB0gOKHkgfrXQmCMMvUKWkUn7yatbigxIxXWSc
BqdUYHIt8wk9AgJwfunHBfw2zvFtTbEujXbBgOCOsRQrI85jUnO/vY9fYbmRmGfH
LvyovV/CYzdhnp4R5tq3kq4ZIanCzXMeK9vctF67I48lf0cMYwtieuhENvNUmehM
ZszzKH2M07qmyqnrwNYMtdC/NL9gwbG+fGa1uYCTQTBVxVEfXU6trSa0BRScO72w
B3x+JEMHaDidz0SjDYUki25+/rNnWqb96It5n3QGTTttnpDSfVzQirvs76RCVkh5
zxvoWk+1BTQgBjcxjRdtsPnm8IFGxrolBogFQAkKF2cYeulP/SCvuWD6qIRPp603
gy9V3YW57nSIFdCUkeFoOC+cdAYS6tHzTlGP6olm5OWWSEknz/IvoaouBQd72eiq
DlOwhkyvmKzlSr7olpz3Xf40gpATYBnhI2qhNJqXzUHNs8WxnGBVgM9GmdfqYjLn
6BTypt0KhcU2OIoPnf5v5vkN48XYrpSeer3C4EpdNiog7WUf7jRobgmI8ntdFtxG
D+hEFBaUt+JQtFmO1cMDLefIaqmtP5IJlUlxlMaKj7AOkQiwt8dnmIpWuMnKBybk
y+AGyuBMshKO04g2wwFXIlSZXjOoevITweSSoFN489RmE5+alvPz2D8PKz6U5uLa
F3e/iqvvI/vVq+bw/Kg6lny098VCTX6of5/mA4GGIp3EEy1EhJOzMwyYl6w6DwpE
yQ7c5KFz7wVCehExv4TgQLX3HuDeU9W+753LTRlS/tROAPCInLqaTsfzb2as2L31
hC+DcrF6sfbDfcbPKjw6uQde7EdGv1RT6eoa1q0LB4+GjYXpV/2Hy89lx9LCedp5
COWySimHKDtkOqAIBfbHLudEvNwAghJMK4kDDW4rqwlOVIeriWwCXVUsaI48Os9Y
mSwTcGCJSJKVhmQwu/Tz7zDzATI7wsFH4fuYN9esIqXNqj6bgVLqwvUUp6lFK1qo
8IogzdRGfh9y9rO7MY3S7eqKmvCuyzoIWfcS3gWKwddTIi9tckC61ZtNk7J2HzG4
P1WRF2u2KbEhT3fzvUd9esrE1NVd8xh8O+izloFUOzliloJAVudheiBoMi4PFe1d
Htr1gG7hcRnYRaSNq4zo80Xv3RFgBE/8FCsbacCRFnQV0VI9zLIXGY9UIf0dPo8T
PQiNA5tmgLTcxqs7G0O3RQA55Y6SHSqp3iMYg8+15KIMvaOciFfjA2mKaYi+8N1B
5zB+0jshjO8tB8laQByZicvStEnxJ2zqOC9UbdSNIZgfzGZzvQe03CkzQH/TZUXe
MqRLeucGLPRb8B1IonX0zEHmxKCmlS+LQpQwNIt2OdUrwv9FFGE2caAjd/KDRoFj
OujNKpOiuQSD3k6t3yOiyDkrtcTtMHa0OpcyCKmZfqyB/nnCrpgfS48PiH+apHyZ
jGHkZV4koUBMrpk3LtCGsLgwqZbqA8410PSUI7T8ABOAGv31X88XJuTSYo3FDpqf
HcnpMbP5/F9SGsvi32aZ6rhJrCe160e4EKU1l6ybuww9vO5/VAIyO7GSKD+ZY0s7
HKx3mai20AqLHKRaG/st/6aiju00A8pS/KlH1l89nCYtOCccePYz34soEeJ7tuOW
HK6xupoXPvdL8DiCD4wSyRpSuKD40bBkii7Yykr2I7XPxiV42RIguLFYSLqR3Qzp
JhWqW4DPEqYFNWWCD3WRlAbMsw/+mBTozgY9IV7SUwlL3V3T1Qb68jj4ao+USwmU
q5cSX1ne+XTr+02pE5bz2mm8XAYUnQLg1lWY3a+gphBvvEGt2PwxXroRtwZh56RQ
J+ZYMtIirwOJhLyoO/dWdCJMyu6dmsuDn8ZfqW/5Y9ZDEU9qrO/w2I9uIqcMUEvX
SdACRiZiPUJNxYQEPf48scrOhE8DpqGZjAakPf3x5VkKKK/67OWKE8yBirOz2bOW
20zK73n3PO1fhaF0DLGn8JQTuqCDVDMBrkteSuf5qORyww86QJjHa5VLn3lzvAzZ
Qn7Xc6qr1lLDSrCUHRp7j1ypni3deUxRlcQ65kGIAQwQFxcUe7Th+5sD/sVJkxpn
4cyxR6drv6SxdUX+ECKzuuc2Vkp9Oo1goge1dRnaNATI+BOwaQzm5e08mlO6KJP4
PBWsmOmJVfOkl/4XV7+ZecQbLnb+cVyZSJ7U56dD4/V/DTsvmEmKQqG+rN0DHhnW
iFSHI+EEPXOFrAOg6VZbYS2+D4JiDd6ssL0oAW2eexEqx2cOiCQ9dp5JZVR+ZGzZ
BLaXl80muEo/to2VpvbHAlFCbr99bY/fPVNK5kJ/37v92HFLcJNLzbrBxZ8T39mw
6RXQk5PIvK7WC6LSq6VCeXbX0xSVGR2tduQ+aPjWE9iJbJMxEfzTfYun2qvSDc2C
leGsPU4X9T55lspcGpYCAmVH0LyOyYFZYaV3ptRXsKFF1MAicF4AZ0ny6yNtp4la
TK0MfKxthtNPdGggD9CdV/ZB9YEmrvmVQjgY7qm7wXBANm5cFKKRb6zK57zJego1
+1ZDC6UzTJXBtJJ7BuICVkwkPAv3ELuAh1emvc9YHNOgU+TQ6Ym05UjZPx17LzeI
P7ZkLw03sPAUaXRy3udPmVQ6XfYykVWLwit/+7bb8VOSuwnwdSrHgI5FjIsItJ/P
oJRi+RJfsTW654qIokyuhBLPzdIalcUlMFb8++tBz/UJDGS3uf/RYURY9j5p6fab
T6XCQp153vH6PHg1ak5isc8qhzWXcrMFRIPbner8E/zeUkBv1MlvQ2p9/JCZW7G8
Rj2lbM+W2/X0U5NxzEKD1EN7DLqCKHaGQKedHwdHPgtPUYRUjsIV3InTW49H0JWY
yjGFERDsHIBhgkq/cxix/PX4JJ3KktDiXPnnRWfua+5098kY2z4zGdI7tp844Uu0
vu1N5FmrW0ic4y5K5vzozGRFjl2olFDG9n/mRonIuXYf5IdOqnLW7ki6KWDvoYVo
31FVjlNJsgSNJALXRzg7AbROpa68tPovTvTZ/otsnJ660sxgOP93QM7nZ81UXUiq
7bp+WhYtr4e36sLAkySYomB5d2cgdpkHFXlTWKj2DTIxcbnA5xRXFjMs72avcvVO
ahsgTjbqBZD5BWtA7TZ/xTckSE5rVtF5JN99NzOZB66EKb5SVYSn1RpKm+ZeNgJh
6dJDlFcEMTlrXc2yNbQDWryDOmY2g/d0CYB3Jx30fvjZ7K0B1ospYLj6kbQcUed8
0rkUSAQdTdhdMuhGbPBOm8tVcx0XOu0jge0vOgXZgTON7P57pUr5bVSB3HNsf7rB
xCZz4UxBniFc1w1dFcsq/xAgyCjaA57QuiNubX3oH/LnXz4EYOsmrUxblDRk8Dnu
JriiIRN7DbciXGMyzjQc88qEkBQVx9ccSavC8+FC3yD5gLIhHU5UjVgbso3o08nq
KK0MnC7kLM48DamkZqF4akgUTMgXw6F6Wa0bwtO5HUe5u7xRLEahXkxamrF0zLby
m7YRIZlWb8rtOyegkLNoSU5SisCIBpTNmqFftPFA8TxLyx4MTBN4ZSsuk5kWbImB
na7N/cN7E7AOauqRk78gOb9xnIThPnkoXy2IAcLaRhv3E/RKVZmBo7sM+8+VLesz
HjpgVeVZXvZ/5pEBGeKWtmA9ePdMmxrJ/kgKJtp0YBfvBSTjrv3PlbgiyCLEba+x
eU/sgtRtTxcnU4jLlyrvU8hfVxuVb/G2N92DewJVam4KMpG7q/SEFaD1/72eTaH9
9SU2RQtIbn/QUJCQZuac9ywhhEFtEsqXAYWkRrvMOrAw4R5R6GC7v3vdCCzF8UGy
jSRTYnUlti7tOxMj13FJ+AgWquE4t8Xl8RQNliMNpYFWxFrneLzRCSvJhqs9Dxoq
SQG91eSLzhj2g9/owZGUZna2HiMd22AciIoxyJBy9c/ItJKcA6WfpBxn9FTt0C+0
m+VDsUhpOWNNNpcxcGrOJipo0worqEGRjl0iJteAk2K9nUCFtr6GmMZMXDvSd8Zt
vOkQsaeANPBBtS2Ea5JKf2GAwtngtckScigPduMEZjMBx3l1NOkC5NbmVpwFUOg4
v/r46V3dp1R/XjWabJE1HtM+wZrUfie6mupcrhFF1nIJX67ZaOLzWXjEkhhZo1gv
ckniF7GyOCMbnmFhl6lDKspkOogUkW1PYj0K3h6TYiJaCyDntkGFBzyTDEDNzyBX
xR5BBMc7sNYwa95l2rtE1VutMLxebYkn8Cj07Q5sQOQRGhJt8UsJ7oUdDYVfBZ6I
nRP56pNoYDv8c5XF/cUjzUe7q3aM0c2kB6NaGj4CpEgc7flvkn6bGYW0KnxI82Q+
KtjnNUsmbwPqeJOUVfA3D0sx3gWfJJ3JfCojNjbEfP0AEISD6mNOkRofTCveu208
/p7aINoVXGy72HOn9Nqnt1kI75vZpfTXSoy9BL9FV2KeJY8B7sz7MUs2lLZqTgcs
VCe6bluyDYG5MYWqnH5i912Ap72Ek2ie4SLJmGvtzz+EmraW0fKTe1z5Kht01/1u
eK+9MfXpA2NVf3QvxV5FFc7wNb8JFvTX18hcisyGARH/gbUubsZDvFgcb3nbkDJv
CKEqUzozkN5H/2Rqnm7kKAppVq0yhktDNj0yU6Pi9PvpJpFf/3yWf/Wg/s8n5iO5
dJ0EHQyjIVuk0ae/JH/pOIF02RqYG6b7aj2G05x4ERX3Jqru9At/21xrktQcDBLj
ykpSfQTwto1WhY8JjSOv0PKTaGtwxCzPNvqpQPqtLUYA9JU0H5UpzqJnMkwiXNGW
u1IupqnBQ8eLee2kkUzuqaW9BQSPa5Du0/VoC3lU9YVF5NVD9x7OIMH9WUFGfPzc
evIi/tDuHncTxetQUbxgupyx4qlyL0757hBCjVloMhkbD4BGwCKjYypSxASGZGsZ
oN3/N9FdMaVpfmkUMtCOfo4mNFpyo4sB2dtK31fAdgvd8q+zOLlpuWqAQ78RlewT
/+UwI0ShRRK+8YhGAj4UTeFe/ZEMDsXHgRsLU9bogLwJqnsgoslCW7gZfh1gjhKA
iN+A+uNu6+bpQfWln00t18T+/KkKqPlFgsF33XtEubIGqqaE54ppEpsi8CvteT6F
sZ5D6COTUCA0R0EkauxIueSKt7oz70HE5rbCIYZWBah7hIGUlup0DLSoMbjxm0Qx
M/9BRIr9//FyQNEJMu2bknhyuMC1bXz4/EXwgXdB3WxuIbJErRHgY9uiFA77gecS
TAanmeb8/+0u014mjwnGyCbjkd+x69hdZgjf3gLNg1ucKafpWImSIgqq0InfHpCw
LSXJ52g0lQAAAg52V6AeLienLigx9wqMfR1gYf0U9WgCJ5Ng4EzQY05C6B4aBF1s
w19pkZ9m9G9lB2bdMf9L6n+Q5dW4PFKh8fJeHVK9ABwLOOMaSGW4zYq4BEFN0+HW
RaeJUV/8C5epkN2wnggdwk39ntFzI4+BvSw41D8GAYLAbPdR+R1judaw+Z7sCUPA
9OwwhAEeQEDUikWokRbVJZ/H8YJkq2QmaMvdfygqC/DDFHMu5VPe2dWTF7B3hWOy
4svoDhL6oIJVtbi9QhJCSiPm5tTH0x4DUK5tXqFCZcHBddioiXisAVBMsT6Wl51/
qHMvT4RZENqpERkqz6RIJNusj8I6cLxLPEWfEGY2hiSRgVUcV5YK7q4l0LnQzSWK
sKdYDqk77vkMB9vzJPKXJrzo6eiTshugbVvFufdmSgFA+p4YoHRu8Wyr45p/jf1d
0jUWhJl2Hmkx2l4ggtz5wDkHXOCRpCBS/TdcQiOyHWQ/XS+7d7BYVdyXWds0Kjgj
W0IkdXWv7VKr+PWRioU0HIY+uVQfyDTRpKHM9X+NeEPIdNUrR84fXaXQUr+XU69N
p4NHJ8MmD2MYNBMzMG+54scABFbD91PYMUwg25WvrSn3hc7KFowIhl/Huv1n2LeB
OJF6/Qa0L4Lz88UIqoRmk76TCGmAvmSFBycwMV5HLDEhJLteWk5KunjUYblpbcEJ
D8RYNjh96VtdT3J7qq2Fzq4ylg1qm+V14HfqU8imF8+uq4QAvXflcSqnTbZVmTwz
oXuDdn5ODMzQLD26e40UMJRPoChEbQfRe6hxrgTkSUI2M/S33wWuuUZXXJ1oE3Sr
5eItGGJpNtDgDb0yi3VTGNPhwUELiy3e6hAiqmXARfpLZVPG8F3JleLLJqf9Dq8c
Lq19RLt0vEpJzUfIZAohJltwFCXYF4RbHvAMhTQa+wRP1eJkH64qgX3S4chGGzdp
GP5BKPGjQYsQEqEndPee9x3W1Vrfznm0lA3+g+93LJRE+sIfCVAQufSqf9/+bONi
BtcqspcCCPaysHHe+OyTX1p2vl/B5gl6lY3vb6HlY6Mdt4DsHi6GzLLC292wRFqd
bwk5Ulwgbz1XkjEv6KxY2Fa/lJGaNz7JJLX5/AOTaTy9Z3pMWUYLigRDTpqA4Ye6
r6brO6sjeIuEG/gbFz+QWYued54xM/ElJm7hvq23EesN+DXJjhqcfBMTEJXZW4Uv
579JMcsgjTcc0HU5bdzNR0j4jspS3QT+/jVnW+IabU446j9Xbdk/MXsO7ID4qPdk
6GATM8nKuScqkgcrXifeo/9LmNFKt+2JvopFpWUVDbKxOCoSJ3o4AxHgtFwlg0ji
9KzixqbjAcsg16xnCdn3oGG2nuhffU1sqqRZsjYkEoaCje4g3x/wTNrdExbKeEY1
EdVcNHdA3ivk/0SbQJX9PWyGzqKvqhetugH4a7NGLqsCpoUggvyB9fn1ESd5e4Yd
DXlA/mlVU7D90So2rmnXlX9W7L/ZvniTLt5toN7d86Zts7c7n++cp+eRnoCD5Tph
iXm9Zg0+uMCRko2EmqGEq8NGNBNuSBhfiMJHL3udowT7t3TGJ+CNyy5+C0wOl7+P
C3ORwZuYhNvnpcI8a//cJ1Mat0MdBznE9yL8eL1G54JatYas9yXgpMfphfzhPZkL
drMdA1ofn5BLKyORstgqFoLN3Ve1p4a8NcEu3BeBKygj4yrNmcPc6uwiy5fM+rXO
Ag4qg++yol3Az1OtzPCxPMW0hIKshhmJGMx62ioGAnyIjMlCAQYAZrfTDbT97V6m
NqjHq21iYvKg3wjXXq9KCoElVLwMmSqFRZKHxu4NdLtCLAZKqmr60vgakm2AIF41
4+NFM4N8IPXVxzOc2Zi0SBhRcFCAaE2xJecJieLCM/GCi2Zc4xdtbFreGhNEEBhx
hFYZKevjNsdWYXeedvNI9keG67NNnMdpz5U94Fxl3REvSBdt9HQH5fpsKPLa9SRG
hNnwSAPMlCgQlzS8SsNYBVkZGoVv0OZjfNXeLBOgoeEmj820sU4bqqEVsuhBPFSy
+3S9rGycdjaeHAK1n3s2vygjXncBXZLoGSipV+Xx+DgynA7eLvB9mufLoQugYMBn
QYhPEzDVKnCLih1cSZRSjwLyJdennjL6MGo220KqKZPobLl/yQSsA1PTshDV8eLU
lFgS0u+NtzoQ82uhi/7hu3r7YgvE4VuhB+vwcdHhySho3AVM/soK/7Q27U2b+0WE
PREGX+NP9hWSaMt8jPz6r+VoxG+JJFm8mvA7OxKsWmZr1SzRR7/4wR5I4oRq1I2E
1Io29wLubMW7/II+77Ed4fHL5Tq/iXrs8ODRXvo1P3gTOtq5c6LfbjyhhKRzq1VJ
D0JBOebOxFolnHWhHbpZIMvhqTBYKswJ2C90oBARc53grankZw4jEs0CHHsegzRb
u8pFQCqVl5NlwJ8CF27lnldbOyv71lzoFWVS5zOTHX9hAIk54Z6yFm992SO3H/Af
9kWdij337lpWmPZo1fW9Zt4mNDRgL9CMRfyC0SB1JU5oG0peLcEX6QdjbKTb/8dd
CPuxDnqpLIvHleyN9zziAm8Xtoa75Xq4B7W3CZ0hd9TPJFXewy04NagqKGHGUhpb
zQlvnTWJqBjt6oKyeXLcqZxwcRfWzOAGTrJTaSPlIp1/TFNQcNscXJCrJ5T1otm9
HwHqx/xeSa/f4cxX8aKvOBRzVXm/pw6QBnDOD3yohNPX9NlqNffj++epuddYks51
J9Vsfykkwq2PK1a8oz9j8r0LtUyV+b5u1TBBSe1cA2pWcrgArNNdAjgnpIyiGhA1
M3/NRlJ4Jt9zZreQG9EkGYJHeyqkGNnQO29ZQPgLE+AgWawlMBFTo+f9+nparav0
o8ftNeEqs6MNAHZXztRz5f4OTTRXXKIm1pZa7pyOmEocD/kpi4meHbAL7yWCkfj7
c7H5vr6L2SSrQEKx5imuwnFuk2/y4VaYaSBnobPLykFcNlUMUy2HWDk7E42ozebm
xUM3NxBWAv8GGw5H8w70rMh96nNkwf1onmm+pu+z2d7GG7c53D4PnPovBUEEIYDE
1/BMeEoSssvDrO3mDiIw9J6xOh5uGfnSy1b6qOnSCfqglIVziM2rlYd89r9A6eEF
Zmmokd+S3HZgZRwDFfdDD/84zbcYCa9fxxLxAPqgF9udLFJB745f/g3t2VuWWKm7
v56i559cFqt4+NGBcuE8DIvft3oCUPt41oullHkJtg8pTWyjAjFQVpJjjyFxyMVd
Af18trSQXIlA4AkDA9kCdD23cMpCaLTnjdIiLb7qDu55L8BPN6OpLrkY7/ZmR/Sb
0QjVWdAZPEIYBilpG7+xZlxBI1ZFEk+fSronA6wDmQ/zpg1cGyqbrGxJBVu3Zb3M
MOhIQxg+FLgcvml9ykTwHP6yfqFtOki8xGPhj4iE1p88VMRj5JRBwRBrfyEsxmS1
BvDWRb+K4U2DpyYQO2jMfI5GrQuRm9tywfT1ZzE86JeRhnc0n1MDXa5UIvSKA13d
ZtB/TWHyG6MMajpptjQ8gyxCZg7xsBGago7SS1MDI6wODbipV2WggivLBoeA3FUS
noJ3Efbbb0h5wuzWX9yFi1+iy0391lxGgC1jAUgdTG2POf0K8CBp65Ez+AGgYEVo
3JTidO8rLdaRLeA/O1jqiuRi0xZPIumdaDZUkUJ5OpBXSHVpbmiceCa9TK7jz/Mb
7rGHPBePUAY8HUlYshl/4QuUHMs/BPYtTHWaPqCuyO4hQLJFku4UOsIp0zmWac1Z
njBEbJmDPHIsxX5HiewLlk/KzxzvuApQGGwuhTUoPAYDu2l20jrRu4wSRXSIdNoz
g87AFLdalW40rZbbJ4QhUDgZPdESTcv3dkJBzFDRhYnLk2vFaGhJjNr9wq1pEiKU
8NGaFIRqbGz0jlAnQCTfyH0XbxtQtRY73H5WUnZbp2MM5Wgmu9UOCmfcY/X1BQVy
Hhq5YDe75m200rTKQliVSc5Ka47rOy3pl7IpxccNBFhZ8+lQkcNDv566eLv22hFZ
ZzVkNRfTojw7SeYflpOJP9E7U0lny1QE+zUcg2cWoE9r9ZZn/bvCfue1Y3trmbi0
48EOd5vT1qub3n2MQjfkGAgMdHSLFM2ORonVfGwrpPjTTmC1hWzkQzvi4Gh2Qt7Z
FdbAKViX/jyT3rP/qJ/U5ytdSe2cSxSQaaW8L4w6O8TbHbJblmIwFzc8uB/jNifC
r6RzJjLq8e76JshfKTA2UeinXOd1h5gZOgBh2geZeOUwAImXbo3oOPW5dGUk34Bz
K+WOLRYijdim1uKH7gvuTRPBIVXpfK99oKmKq83uVQNZ6tvihtgOcRfhEezGmccb
iVqKFJDOHRZKXs1ZDygS8s5u/PbryTQwiRC6FZYasgfadBKgX/qAsHViQc8YE4h1
QUg1U1YvrzIeilqQfJBBPezw3xM40diin+LrUcuAY37VYLtlDRQcOS8bcGsg8kVM
9k5kFbfHOfzKHU1uzqOcL7h03zudc6IX5SjeLNI/CZp+f3UiUBxcARSOGA0uYmN8
3cyEg6J6EFMg5B4Gq+VcDmOeGWVpZPnek22IFbodUqhObXWhZe05hf/Y8P+KPPaZ
bnsboxwyEESsNUSKEPUXEKcX+W7z8X8d26bnkKpOrkwrIKBtDyoUw0LIbLOjdjZ7
M+knVgv/HoRRh/h4fjTqkxGioJLk9bNeu0atIcjTue4pXrA/EAotiMVjdjGLcLOV
u1ae5jq0ByRSio8l4u5PsD4Pm3YGoaCgNL4qgmHEPmPs5De8M/izZqVMufiMWv0u
zxvwwVEXRlMLtFCJAx+pPXFZEt0FChPXRfgzjrvCnIBOiaVZ7WrVFz+ZooxnVpEz
hfPTYGNswUfqKLsQ+9o/VIejM1NLYH6rxomM6DwBNakaxthXXxC4vw1BFFougbz0
ZAZLYUNNRjuaRwi6sVFp8ykvztEImPvU8P33EcS+bQU3xcMDhE5+Iknw0OcrIgc6
E0v2OYESdTNFbR5T915AwseScNBJaDjwD8dcNmfvCO9pe8tFv1CzX7JWfQ+rhxUX
bvZRldZtOmIzTsDXNYBth5gVjBqK0HQ1qk4N0KCUfScYe6uR8/SIPbZJSOQLz1dg
iZGcNytKOq5tUYt/yMtyOpinQVdtfdskq078h8BdGf93wziZObAAxFkkd6WuPEgV
qZL0EVVKQfs4H15qEBR0HM+R8xllbuIUYE9SSfP3NPDXGEMVs2qiZiubDjQzfJL5
7Un1Wk4dh/FP5MocnWxNVIE18vgXzASYhIsBqFM4oFqA3/a+ngNhHJiqSzsdNNQQ
IlNp25bi0WIccuDZApA94dYVbNqfWCi5b3HZB6/CN+pP1ctObSFTg9nwh/AnfMS+
zecv3MKEq8wHZgr4e7suTl5b8raXW+Oc01eJ8YyWODEW2EJWokIbTtrPh9Pr79Vc
vNX117rMLVOnyFQSVDUve3EBsUMl5HfTfme7EecV+AIQzNLbGYlDpVH7LS/RfAbf
YnDha5LjzcVilFCpkr/9fgXNHgq8GGGwV40J7GXFVyptIlVpNRfn92N1k/TajWFy
HX+oXiBBTNIG2q62iPiCeDPwf65ZdV0t02XifJH+6fbE6yFEc4MBHqG1KDxwbpzt
yEgAMw70FYn3lwCx8CG+vWVZSmxvv0icGNcGo216l7ai/BybzffxcemTrYfhyMlT
sVKEoeF6Hn3o5m6j1gzWSsaBE+8VKsIZFlkoek7OiEh0JTdIkxSNllAkYK7pO5vG
95A7qoCfTjLKftxNHVePCFjjwlzG3zqn0/2FNiOUCIwmF6nYiNUEJdcZN7/Slt7d
v5mKgMjd3weAqywX7vaAFJVyiZCxSVXCNcI1AkFJL2qGmdbByrsqXx6gwnOznJHX
XjiV4xi7pEpEObuGfnPPXfeSMAx2fQbX0YNmYfIIXRlTdCUGIDRx3PQxo3eExrd2
U2byV5v0KCJxKHTq67VQIfqE64jaEpv2WGwW+yYkZGSUl1RHLCc9PbYEdZeCdx/D
/GDwBNdwtv4l8vGiK/vRoEiqK5posEQtITuoKSVVEEmvSgBp50m+KPgTvH4lbmfm
jxC5XQ9EJzKDpkD8GQfOeF9dLZwn4P+jCSuw8tKVfxAhmUUutFjrrwuArcBR41hC
qHm+z0VQibRB+lAelyyRI8ODZHB4N9nmh13pZf2aAPGbmByGOdbMIiWt5W1IVVQ7
/FHEw8yV+VvYLx6D9lLePfdPW7nWRWr/hUSAp5fFPJrdQbRc65X0l6cYVyUvS6jG
jYEtklBBuxDw+9KT4ATCBUCUAEC5A5qnETmlbNrnJltSNZF47O6zil2fZ4Y4mRla
sWdNX8MWvHjQ+AF8cCfILl+KUats015AqPx8lEXPmZmZVCWhqvR6nzuXk3ar5k4c
FDSHbOrRrfq7XQKN4mUzjV3CHVfrQSwWelV2CBQbI2rOmudhk1dAq8wwVwxnq1gx
W8fQvPCmbFEqBPa5pP+dOKb2kZthuxqNGgJV37P8yX9xuBz5rAbTvrSagzDF+r+Z
F2XbYPnT844AcA2gF186Kra5Xu6taqtvgzxSVmSa9FYgA6/ye/t/QLa0YTn0crnH
a7FS9ZRwP4DZIQjlhzdllW+VQlvIlWxxJ+bgfY1rrLJF5kv/XgQbyPrQtPYDmBqi
JPsd2FUE1uvkKwdF+p/UOkc6w3cwWeyaGOKMytnPckFU3HrH136mpd249DL2p36Y
odzcglaRw7E75wg6fxZ5/VyvDSrwTU8PXXjR+qViPnP+Qus4nNKv9ivd/QxCtO13
p5eNWmWgNJmgIh4adcafIK9bKTwauzL+QyobZ5o83cRbTuWnaXw0EFzYmYDHc6ee
6j0IzBkAd1WwHZXByTHqpHjesPp2lXIcS4L0AAda57eM54YMeRiHkH7wYujdaqaf
/7T2VtgPg/ro2BFg/xKsqDgPjqyVbb+lnkaag4T1/U6+5EYyxzJWanoFnJsCBMKh
gJMhWw7AOwojg0G9hAUziFgNEOreVvYgzYS+JLsTBP9mDvBit89AiagNG2RtBWaM
kHVex0eGB0Rms/vhti0rvui11yQ/BSDK65mkT5rt/1U6oPO6biZzIsuSitG4RF00
Mdxbx3mMxwCKCCYS5E8EMt6wgWzXCgwSBWO+Q4Q782ABwAwh9Uy57GHFYAnu0ACp
/v3NqlBfTHefqWT7gTrH/C3FzeNNEpjmZfW9bON4/LBe51mHNPkBtcpM9iB/2ZLG
wiIvrhCqqSKLrBjJZhIgvnpdK0Bozh80Tznjewqaeighny2MnDcjN0L/TES/8fY5
QrEr2OEQul137mIIpHsUJ28PmS4+gl1e6VFxRDtYk1nGNmUQhB137FjZwpRbW5Rt
qk6I87TcT4yz5DK27uo1Dqgw7wBVZQRox1q4SQuIHgdCFU94EQiGsBFsty88xs6E
q1ejC5vzTonV1G/uIusXOJuFMrmT2RMZp/GO95nykd63npAjHqAtmENxehndyhLn
CEqxPJt+sG/nE9e3d6z8P4pCUZhmMTxZma3l1cDdgMf5FG47rjbhD1y1l/HrVCDV
zA8HaDdlpSr2p0CMD9lJCb+vy4bOWSSSJOt6Bjc8qFfw1MHVAQSdsfIYCxJputHb
cG0bNDuLmFySwk2sNu7DrMLcwvVh5QRyCrkQ1MXqgf1anhba5+kUHgJzxiEEbfN6
odha0fWywZDqadDke/WoW/N2zAr/EqdlNeCk2e0LsAwoRSYxr0HO8BPm19f+Z1tC
uxHLMFhO3TxZT6rMvspzECW0k86T/EmjRQPXdJpXGkZL/8DcECV7nA2IQx073e7x
1OYXkt6W0/rf2EA/AMaASdGKorlEYsM7Gv+mt3lHQIzF89KjME+2nNRhjKKpEbEH
jnj9SH8xE5KvAaQnwrGW6MVV+4A8Wr4t6uTk72dpjHu3FKAjMK2bcZc+G9T8YH9Z
mC0plQR0LSsiKZCkIC6b++RXMxWoULthnDO6vhPjqwL/ORkB2ADRlo5yYvJT9W5i
Cm0ACIiU0H2JtP7iETwfO9+u+RhfR//xutWG8tCL2iCYM80DbvUe69p5G36mdSM2
t6JwwXdfjurR+dQGqYquPtvgf3Qg6af9qp3FGw8BA/CRywfuBUiM8/OfjkYSsVCu
fu29txVJvgVh3Z4PZwAq4vGFDDfF/h60w/hqrX1eqyc1AvMMA3aLxIDIv5ktjprq
7zRHCcsqXOKX7Koy6tIF64InolzX6u0b6t/tDsPvKGEGoIaQwnD0YpsQLf0zh7qU
XC4qrfYBaz2k4h6F0bEoZFN5Oj1H1DrdyzkUJgzavCzyOE0HGa88N4m6b3r0bXYC
dNre5wpFi+7gMCVHouBf02IzNkZI7pfFnScyDM75V07mg2OHuqYaYTl7SS6ItcuY
Iy6DunC6yPLoO3NI4xDdb+TDHf1msz/nfy01mpasNTcN0+XHQnzdPrJh6q2S6q8S
6NBHhS666UYoeV/nw1uyN1rYrT9Td+d2hFXvEZJWuYIx27qdwlU45CnCZLMevuah
Wn5+jK9eIF5Ves3FCfkCHdu3qY4EO66tBID3FP6BKMa5/8N1WVmSvMMTUvk7AZJb
5PhcDYi88jV3u6+vsUxjjF5y4R3XfBY1CSjxQegwkmoQ8ltpdzHN9Zv8BhIpcqv2
mX2r1kKEQg19gnhvQeAi6vk3ctZsB7SJyObcqkbU9SORo1eimTN45lU2jNQYMZSy
agjaGmrBKx58WyTSqS5PmIjVl6WjKD3e2Jx3NnD7/znPaGonLX4nE3f2YrTbkHJ+
9GRl1W/Vl4sCdTGnS7FqLOXbnfYrpRph+d2kAaZbxrJwk4AP98bNXIal87b8B8P8
333Cy41lsoXko5V9ODfiiAdlxMBSrp9UUiVPnblXoigMeeky2RySkksdDigCjaeJ
8A3m2GP3NNg7+FrygntITCE/++cu7Ieotm8yZEUfdWbCDWov6AUhIbWz4BbJdlNL
gsS5ANSPaIArGttE9QVXJDAYI7FcXgdxyVpDaZJQEOsWOWe28YMYkMIBYnw+ePf2
Vssy21JYH0fTuU6CNOF1Uaw+EgT0pj+sFWA0A+KrFOwpDYPSydWNmayKDCbCrZiZ
P9gWcQMbqqxjS3/EPVR1K56BQA6Ga5e6bfmtJbkACn626HrJxPu4aMKnPB4MvQs6
CJbzpKrcWfnuPGFJIHw422jxPCOXoTvdzPjTDHx5P/snxo5aFdBApUFo7Rrhr5bf
9rzIf93+7wN/w7gBE5Iy96rHUiOGLHuiq9OKVvxzY4oXokbo28TkWf0s9R8OoaDB
IDhOrcQX9VqrOKo7ewA1fuTb/0UcSy25hgr8lnXztsGZ+8ohcv3PmCx2YLS3+ptH
pqzAhlbpzgJg6QE0RIA0t0iRiYLiniCdJPxGWRDPJapukOa+AXROtp4c4uJsR86W
0CLQzlRsJHQAF6uScAWTOXrcEUl1H9f0UzsaQwt2tj5U7B/cp85sLuSrJ8Y7SLi+
PrxHEFaCyMFJgz644GbaFp0eg24rcMCEAEyjXspCTDifWsydCRoU7Hb1aTKO8SKE
SbCIe9HSYo+pdnQ3QEK2Ulb9ycimZqc/agpmcEyVTl3lb8KgJYRZWz+ygOgd498Y
czVJ73sBsdrNFYzpHCYdmH9f6gSk5m9mNedv2GuIqzwKFG1Nx4Lv/5kvr3eR4dap
TVNkfgCmivbkShK8WroPBEvLNNIg3i3ZAXG8mT6K2ANJy0KeAQ7WqnAaUqUb5DSV
eiXKXNo8tM0awHOCuUOGBn2MfK2+ozdm2QfoHnARirjsEqxQXyGXxkPkLZAJepqK
eJl01L2oqBUcEbifS+E4uppZxNJUA+mGoezaoAuRPUeUGCXcSQ+QOIq8n0lqn74h
lJi4JpoULAntPdQalCherGY3SAJm5L+RIhYpKvrqvMspHI9pPHDLnVFo/qpZdjZN
HFfLgsx/kYkHulGdLDkRy60RhORkZ41hHWDEEt3DmavTtftgqDwU9bcpG2Wc2Rle
IRjdR+22189RDVmAvPFjiZx15/dM2WdIjFhrLcaLmfgeRi7dXR3h4ptLIG0GKUJx
kPZRVkwL1zCb1jriexZxJDfuvyvJWyvz8xp3XtY99qtQAW86Oi0WGRR23BMXCMtx
9kqLXXtjYwyHCymW4/SkOaQyW9L+rkejBqp/fBdacpr7YxJnQQ7xzkiynpIOCHXR
SsRzBKrexKy3o1aEVhHaG0J5H+oTRYwQ1PWKLGC1z5j9BXtcAYIxdejlfXsHU9gs
nxih0jT3dHXjHWC492wSXw9KZJeebxTGoY3m5N/T5L/lpLk5AHmGoD/OaKlBpWlB
5rkOho6/+Fe15kPVzZchigOQnrr93218BMGhvInFvW3PoKaR59BzBCzQFWboWb/C
82UO4KduS5O4IpyRhjNdowTvzF5d06YEKPIdoXntLQ9iK/c6snsHhulg8UsqcoIe
NkN+p5bPW3P4Xr3ivAQU/H3EH0VXBjwwVInd0myRdHiNV1FDElbRLCDW1CH6swkr
zZDI5M3btOUcM3+6UPk/bE0n9RS73gvIZFrRYu9RXQYiEgt9YyYsW7qf2Hf0pdsE
VTe4FmtcL3xT0Ep9NkviTLq+fcqiEIP/V6LU8Pk3AWaMD2lMdaNnJ4H1wGBI66BV
Px/bVYrX+Ig9Zg/d4XMEcFfv+xITzvZs+WY5CQ7WzaEBgEp6BJ4dIwg5FSI8mJSB
kf8sClh3cG3Fu49bC9n/T5JGJ0RrfyK0YF9NOZuirVtaQq5+2qR6tH00QavR7W1W
FHcSUo6PtgKhyaaMteUxgwerDfF3eG5WwoMTOdy/dByG0BxC8pdXqNmh/DiLlQiw
VQROkLw5YhciGXPbR/fbHyGMZwQkekPuPgDC9zdjq3ABa+EyHcn2jEC2Eb2/TWwO
QkPmynyIqcn8GKVVgejYln9+7+NAQwBn7LD0qxy2FrcXLZ2VOUQu3AUbFK4TqqA/
E1J76awc+YokEeKUfCu/alVIrshsqy6+8jQubLp4cgM16U4Djqag1J0nkwnbtF2r
6Ei9ysVdB+3KN9CulzIvFc5krl3bp84sbelHsuu/2yG4ihhexbAZT2gqnYOGtAlO
a+wWW1jO36fhoUKKizLPP1I0Q/Q2MySxfpNCwc1I3+YA27BgGDiodnfShRa2VUPE
tz2hqSpc9KPQ7p558cKtYPCsOn4Z6lrUz4fVuEmImtvFo+AckltRBfZhJ0r5jjwV
vHzvQ2KvGh8wvSKDACvbrAJi6vlefEbZNtjpPv0rlUgeBxfaHd4FOBXndPEGPkvE
wh8zO2FmsbO2Tb4YBrO6n075kB6sNFjM4TgEGY8guhsQbiMSPnpVC1R/6IKLYiFW
HTAxr/quQaek1FHJm77mrhYecKvuoQKe/E8bpeyvA0kD/7aq/vo3DkbdpJESDK2K
q5fnabquJ6BFCuzVVd+jnpJ1kpVdmy/v7+gXzIxE2qVUaUgqcmqajspub6zuVbKd
2Bhgq+NvHwZIQtQYJBslwsHem9GrQ3h1LnRjJU9uc6DZ+IeVjV87KGDYoMryoIKk
mh4mh2oGC/4PhxtlCxaFWz1CKvZJSPFeDAYoU74R8qTJHjV2ojvxvGTIs/lW+NmT
o3J5BqBHaE+ahXk65GQHpUMcfWFXUWaTf9QFMG/8gnN7Q0naSBHLg669yQTPbM95
NhnpE+VsECHNRvxwCkoas7jOBmvPlJ/gP3c6MVY4pKEHaD++YW8Va/7Rk9lyEqpT
wPpiQpMW+4IfyKsAO6Wkd+1tIz+K01uVqq3EzHKe6y9grCVtOXwzOf0BrtLAXT3L
mdVGWCSajM8qL+N1KB46eL5PDyT91xLlrlApd49BTEIdwdyLlviaq66Gk3IxR2q7
RoVYadcKefOmerav2HtBY4W1mNFRP10TsBxUC7BlFnYcDhSxEwZmV48RxeOzMIJG
9CNZhC/q1G1SGvncZZ+YCfsG6zBQsSOFbf34NLJD8fwKY5pz/PqDTa5Nr/bFBCwo
ERNwu/5c6P9M/N/vn0BvpY1TrsRnV+oR+E1Q8HSFq4V7F1bHgx+GVYwbu21PkF9b
ylf0mrrfrcqNfRjozRrgchZHzpLr2yJfZ2iY3X1H0x0mOww/NJ0Bvza26hwJc9dG
7xkpMxLNQpG74PwkNE7eqUkI0mIhMMK+jvtIm6fkLTSmbLaHEBxrREmfTx2nf+7m
uYUnReg5bbvb3PmJ3QUZq9ejGnmk478tBzS1/VvIvFltLP0CvEgIzcrmVK73dKhj
GrRC7NIDqkCLh/eZ2fSUDg8eVzf3+bSYFAXWE75jD/w4uB560uRsz6y8eljppCZI
4Yy/ZnvV/0Cg6vF1lm9gTZTGtL3JtwFcs4LRlTRVOUKCEsXUL1cdTF+CyYOM5fxI
BfQSAj8Jt6rMSfE3ubNpd8TY2qLVgi4Pk5Orv1HZ6NnHa92kheBFQ6ycpq5+uAsn
1gh/e57nLUUxenKlau5E+FYVVf4eoW4KpkMUHuGiYvVUiSMdVZZkHZor8Fg2eYgk
VAPlRqh+rbcf4Tovk0DuXFcKenV/nrPQ648FBB5C3Xvt8gHRIeZu8yLCyHk4XTFU
ekX8FoeXghxlnfr+x2M2gmMtFC2QUZQm/Oc+womD5a0DXakgJTKZt6DUiVGR0w7/
zdtbmISpqnfsjfu0mpjB6gvUB+FGq2+kQxanIy4UHX8Rb4zSqjRC3paOdqUwTntY
meOLzdzbDhCtTs0YDREbXyq6qGuCcsDV0RdbGRYOY72hBXjvv5fH1GrO0/gefpJG
McAjbdiL+fCEobNRFKoOi/IcIgDHa/C13UBak72avz+TE3TMja+9XyX8KWLE1D02
jFdXESUapZb2M1ApFviCdVLDokfrohlK+7laYYyMAzyYJulNybcyWkVKhctHf5kJ
OduPv2wtPlZYI8Z3VE1bxvqt+NVMZk3vVkjFR4Ad4jnCJV3WYYUwDqtZXvx0LROs
ceSaQs8/2CqT+bGwQATijhROgEhRR/rLie+D21X/Rufx7ErprC/ebO+tiIE2rRlW
kSwLmEQDq50AuHqAYcTjarpAQpa6mknrargk2suFfTwen1tjffn5AW14VgEvPU9H
3Smipizq9ZD0/7+D3NDuiEgiWBnGeCqysFjGH/6FN+3OLJo8v6Wx2OICD4OY7Bak
073ZAoN4pbNBMFqFvU1/7+fweDR+thQ2bRYb9D7yvJTub6pblZPG9Vh0gX39J0DF
6Bd5YllQWVDv1UT1qGR0UzvFyEJdCrp1P9kpVT5YDw2Adht10T73MA6VLmwF2ueu
fwt8NJMrxuljpcJ67COErCCqAWHtEDCYNhu8pkraWnmDYe2kgos3wt8A500FeINd
IFIHW2OYKWBPNbsM1tyr6VnR7Gt2IPE++e/KZDWTcOZdtciTxZio4MEQojsIPzlY
qBpu/e0zqFIlvOmKQ7bwoUTlKEImTpsR1Yp5s/IY2EpFkox+GnZqnDKikj5VjVKl
X1GVJtGGoMUFkSmG+rBCcl5k95dXO8ND8HCqLMyUFSPIwTe2cuQLJSdDnjo2dgpq
elYww8E1nIEcoIHhW2TQZ7ol3B/b3Tl8sfaiVBmg+zZJ9dME3MeaDu6jmD0YJ9oE
EbTB+LJWeYGtMx9NhJV5OZGsdCHqaA3g6TCV8HAKu/EewOhJ3vqHEqYz82uOiicF
XMYfqxcNbEm9lV4BJVs94+z0av+VRsjON0zi5e/j3LT7oKEZGGo5qz4ypShi4+gw
xgwjuurJRO4lQRlzaJNJsGxBvKK0/ibKYWm3Lj83qbeSjAvgUJKuMkDJ27j9dS1S
QSxC4Pkpk9mR1MFMOtijbve2QaBXS0sVSvvIbMJjjq6k0zyBIU6DXp61/b9VyAkL
kT5rFp2XhBQ+R0oooUZ0P6C4TOfPRZAr0H73GgJAtfzJX+Tby05ZBw+SRSB4If4U
JErc+bEACTwdvWzDufbkgL7ZaKwOD9ld2pnXiK1S6ZD22MOo9bPeaNxQOX4UZ+G4
aU/csUvy13PnSJy2dA+Ob/7t9VrbSVf1d2Msg05LXVvY2dK5e+rEUCf8h9/V8z4C
VVRpOTmPvFeBHxa0AgH/BFuzvfw/Fud3UUKHQwid0r74Cf8tGkM8NVC82oc3Y1eP
b5ImB+2ljzQmbEYo1TgREnkcu5632+zs+WDapHZ1wZ6znUA2JAKIa6t8kmU++4B6
7QRZcYyqriWSOdbI+hNGXn6VUpyUo0KL0JT4gQFuf/YZ3QAnb0FE/cSNIXXoqgYD
cS23MFJbROJjCDKWtr4KJxEwTh54pBvXyEPRBLRCGejmad4MXwSE+ytsKXqCZ8dX
o62zE/8L6gf7D+ozJX+W5qFJPhIEezEZZnbveHhV4NTEoimlOfuq2w7NCDgi1TdR
Hjaplmz4yF1V3SIwEAun+1jqakJJyUtPZi1nZOpzDPikfT5lxb9e3OzIeCrx04YJ
uVYLtsP54QwoTBv5GeBVbKMyPGcmM7LFmjg2QiuU40/UJX6o0pSBkcWyi77+Gq/E
5f30JgqJHqo4P6+bIoIBZe+5gIukF279IFNnlqOpb28eATMnf2vfLp6LA6rlE4Yr
O5fecm6WQV+0SNeV18jkZ5avQRwO9v1SO3L5ELRkdvifNCGIgqiVcXhD+7TVuqUt
Gvcg/A3Y1mkbdGSBH/vMHvuU+sZKjMtHBxQy4FxHPfYoPzjHgKgCdwG3P6+H7MBd
s69xmJJxAqF12JPLmkQ6ddR/2CxCwiG7S6/HOi204miR+xQweR2ptOgKZADgSYk5
HkGRwe0PM2XAzQFUn1OmgPx4sssv+LGijg+9oYjXUgGsgcpB/xWbyqwgmg25Jptu
M9JX/yNZiYhHb/3e7KoPpZuhL2/JXU4idWcIB4JI8ZXdqsWJ+ATISdGtD+rkW52I
GS82VCApRN2oDnLFoCfJcM9fvesrwEE+pFQqtWdbb0h2Hu5QllKEaDOnVkGaKEOA
NPLmkPRKLZR4W9Ru5dm6ARaCHUDt8uod7ZaBv1hx3yHXfI975v7gnlF8KakhnbMx
WLPWwEy90gcD1A7jnVc09iomjCYtdtE6BytEWeFYD1UeoT4OOei61XMqCX1aujph
Ki73T+nq0l7JerSucD9+ukEJ8JRQdC7ryvFwmap5h6XnxHqqXB7Lo7d0Z9AMBr1n
NgZ8cGMELKiXuSRLop/Y/z/GI+w1nqUQOquwLz+8REcLmivgEjlrVmsgJRU0X/Ns
8iwrrui2FmuYlBLKjS/kl38YXQqtr0A2gSvM/K01joA9eNv68zfAs52+QaaedKog
y9c8AXQRhewlDP73ubA8vIIIeNynb34/YOwpewTX4Y9IKATZEA/xxMj0lGwCBrCA
wgXM/J8Tekgto/XLlZ2+dV3QgypD1FCMOzeBmiVRJjN1fq2L24i4Rrb/yQU87Mex
hluIcutpArPK9VBMeJcE8E0yCyfpGEOKuoo+MXjdtl8W6lUlAtdR9hIQsmQjWjnG
MptF2uaFzJOn2pt8wYxWsXA5Dl3Jx6L1YbzaL4n+t4JuG6YTuBY897+JEafz9M25
Kb8wMhd9Bq6/L3nMf0UKDt0US6uC271MGSbUaZT7ISewL5q77ebSYNtNW1vl9BXe
mPDNbYK9rQmHAZgcuVdNMxUAzPceifwBCELTKljQy3N5ykyKzeeqsrdr2HYmhBYW
7MwFrhFmASujs6MccQID6Tu3HvwX9zQRTCUGozV/5mUJD0u/+koR9uMNKzEUkpj8
tm5AT8/9L2QVaR15hedbfXjnHUV0UQJI/Lc7U1AdmHtVq/Itp9vgu+6y8M803nO2
URwumN9BaGjSYc6IEaUCwQWeTsMJ/lvwnd7SxqJBAJyIsBzIym9pCrfStZKfD+RC
3xd3vTg51kHXnkIfN6rECxUMUL5s+/JQ0sXqLtAT2j1sKFHed1fwliKKTLMikO1d
D8aTGPorbJDwZiQ3YmBxPKIZepZW8BuIzJv9V/tP/aRYlLf/8kR4/sdu2CHd1BjV
/h6J6wyuj92Lea6ar9bsX46GV3CfstZELUij+LeXVfr0vKoSxPuVW9xrSMwJG0rH
EwMI4deVnh4CHv1Vxi21e8dfYJMEzJXrjrxNz/0iNk2T4OhkVjoRm6jUNBWvNUyA
tROVAzyO0wZEFjNKIyDETxYHVzRI0OQnhbLgInopWbPom/tCCXkTpfIIo5ZG8l+f
v0C1BLFrUQlNzsvW64KUxSHy0Tf9RpNwUn0Ix4Lbd2eLRHTEM3FumI/LYhtjuTvk
/cXQpQQIHdZZzCJ0dc99Lo69IvHdi4mr0aEfej8NrtgWl84muCY54J+YmmhgJL4L
qSIYiGxLPFsVNcUzuT6J80fQInKMOE3Ce1ZjB62knMSHc988rCzgriBxOmCGhKlP
lyllqd3RcIiooiUTieCUsqAcMxQXW7qpvm7uE9sdqS8ptyreVYSgoBRMvYSHceb8
FB2DDEYTDyCIIuRoD8/gJ01p3fvnbiny/V7FcbFgYunFxqwcoOxtrAZKtSYjmcb8
lV41Aw2KMWFfsGDFIy4uwFaPOmj8XGxoNQ9E41aVJ5LhXp+Lk7qdZAhxPOQLkSoI
sBIBxchEW+/LqPNXuQIyuaW6oxsltCvYulcVuYP5WHHt31BkXCxCsExA3L4fI2Lc
aMZ4Us2kXSHOL45c9rQfB7yIAvbb15ux81F79+AuyPaNqAAwKs4n9gDc+qn/WGem
m59j8woKRBq8NNWarUYX1Q/ZdLJQerfUUpHezJ/8VxrINrQBzkFAezXO8lVF9txM
8w4vYpjjSMb8ZK9o664RbY8226OVPioDExmDAecIwiBURq66P0RfjNSxvNojM+sQ
CqMnfZvipoICogysBwnyj38uZ6VgE7GMsEKPg4XXp7ZWFXS4HeSgb0iYc6X5Y3Lc
3Mz/2dTKgSVq3CWkH+TfOwa6JkYwIRDC2VmSBFg3y8+uLIfduHrEXrFCRMLRgRER
04zzog7/9Alrh2zWwa+XifQlcQG+SR1NE6DcZNuxTp2lVyLrUYNGUhqE/+iHo0QO
9OTh0RjGhYKxUzrh6UeBdbKJhLH/5SYpiD3wdRo+xbcDmH4Oy2aTI5oN72JiBeiV
KAByNy2IIeJMCKh19y+dkwyjRy4WwqrpbEZCnTwhr+ckqV+ZJI1XaFncMKtntx1t
IXAgyHNtCTqO2kVSrQ91bxArvEa1YAiA+wZsTdab6B24v3fch182Hx/52sjTJ+Q8
Eplof2WAZW4EUx+3IvQpQiB0teY56Oz/U0aREgGDm3Zx4oiGh0dz8iKDbtKw8ZZs
s3/SjV5lGun4toazciy924rbyGX7jLT6Clp4pBgUvv8NS1jGDfkAiVWqKG58dWdA
KHY13r5IwZw1BrZeL1mwoY+7eHTqFcZ/NOJoBzIvWqgibeaIMeRUqd9pscyo45Bs
8H7pJnTBsBfg+H3B9FqICNgtQle+GoBKf++5n4n8gDY0QyTkrRnosoDWM5/YTf/V
S0GhuLbWNKcPdzTnIRT0W8pPQ4J/6shKQGF/htfE0i1Xyi3b2jfHN8dqWtlTyZ0H
DNOB4WZimoLG4o2HZo3BFLUJHS9ti/kjGOqlH3zr/VP0gRInr3MQw9cO7ZMN9Y57
h1YyQ+ZaIvCGnISefSls0gxYPkn4HHciG1zq1t7gcItbtzsRgxoVLbf98WJ9QFZn
H68J0Nfslz75y5Gzn7C+43hbNe4q6c4aJj87FUbYtCAYjG01FeeT4CVBuE6YMMBK
Dfc7CiyaBYCfLg103opwgejlIgQVKeTveECV+PtqQxfM/qIy2GdvNGI62Bif1XFp
s9rRzBtL9C6Y7SmWJ3ZJPHWIq68FtP7gbnBltjK7jaHgLn3hK0l1ZLTmo/y5z7dT
Lj3/7otYDXNojLRGVfOIz8thY8LA2JqbmCY3Q7lvHnB16oygDYyxi8V/DG4nUUgn
EW3PTuWhk5XBWRpiwlUe34la78rA5QyVpTWFwe82Vq6VG7HpE38quWpPiTmDf0AM
AcBzglDjhM3UP1UvHPpwLIDF2ld+lE2YEcKauf1jqas9c8Z08VOF7FtqpZMOYJUC
Wrr7WetroA7q/kChPOweQ8xLWJsn3tFjZDONY9ChXWXyEzaTf6OF4WLqkITizjew
OXsFUb2EbHBBjTFXEv53zvTReD7oNveW1dFVlWhOXhogKx4o7mQ63YbuojAmKIIW
x8KHI/LulBVmlBk4rWXkkD9AHyHb9TLxy8V2ICu3zjyjXzGfAGKcgmEa98Su+i3K
ZkllTFWTuqR7RoQbNBIvBwErJ9zjSJdm41LHPKv4zzCWXWKTPdieQRENbcTEerll
tDSZkb8SeG2pv7fi8tHnRMv/PznZMZQwu/sRuBftwx3iGXHy/tazNbt1UlY1x2jK
80abphnXPfx01TOmht6SUKmKQfSXgbZW6EsqInI90trLNe2sV51KnAeMDWWeC7QO
QvXEPqknz73GDNCnsF2eummy49mp6tPlLyhHrnHqm0ysYvimwhyPXgiZeXQCUOYf
vyFQTyug0LWzMfgL0Ymx8dU58bhSQ+j+HRNEoS5RBPl5ws5ZMGOh4P9WzaA7WS8y
d9ZOarkHHD30Exv1VPqwU0Fmf8ZShBzQZpjRsKuRNNi78UEOuSRWatHN4jc/NbHM
tqF9EKBJXvJJSu/YPBCY35T6Qwz8oPXj3qRzVNuLhJ0YsA9+6lee31oszcrzTt6W
KHvrL0vETZbSgkzvCB2yRIHpe7zliaBtT2TvU2h5Pb7ZkoSbJo2afh9YjZwszi3K
3WY0pNTj8FJmC4BvsKUwRT/yCP8GX7QhD/KNiPElSpkazBIjMsGTN06caqAG7UEa
WmnVFkQaByg+Wlo4rZD2Yd5/vApf9dTMBa/nB/I/XDIvHaHtoRTSMqP7SC9CDX+E
Hr5MfunHu6nj01P0AaaOW0lxhNkm5uiq37yKg417SY1p/R3rtqPQp7IJTYydzaT0
hpNpsALvhzNz8ADRZeuEsE5+4GAxL2ln7TVPRsa5rqamnn8ZsNxd8VAp5W6VY04h
TmPxD4Z+3fVrht3E19d/Sni2o/Aze+ndIhL60dD0NEnSLaVrA878mc5ywbqerJij
KUj3P69TME+Q+AUPhmpouefdnKTav466Pnr5V8iCuS0jJq7HPgvkqE74mKtzt8mF
FGOG47GHCIgr6ozST1GJ/DVGOqzRweQ6iR9YXdCd9pef+13q/7LbJoD1kgh0PGXt
2iaWQWS6Ip3JN5ECXBytDyorUajtEtog2ikKuwcm5pX72yh2tY3YtVCsDQOEf+Dq
CX7t6PTZDqj9mpfxoRw8JGG5ECGZAoMrQN1AzI96ai0drj8kmzNtpUDnAf4YBLvL
WKtYW1/9NgmQ17DU4iVXGmmZK2tKGeD/qYL5ji1lkbfXkWt4tqZfGYfwn9XTUnwx
N1lAkm0jlbfcJacxO8sH/cQcObe25ijofo0gBu8h8lSlsDkpX2b6fFHpUAharRWn
fuzRjdtyOUFy2zWbqs4Cf9nbfna7DgxsX5+dAMCqXaEaIF3GgUVnSoNGz3m8UpIP
BX8fXVbS2stznqmKQguhzLdGmJkP7haMDkTaJ/PHyQKREPpOCvyUWvbGZ/nyMOzY
UOyUut3jaZa83PCKLQgWMmx7ovchlQpAr46N900bX2beHo4TMIcllVZE83lp6gKL
zc3VrHyi1YGT7w8XGaL+7oU+Y6HWc3Jt3TsS9Xll+P/K9KXmwk5hp81oe/cikJTc
v3XGmmYlDkYmnBK67IOYhYzO597I//YO37lb8g5SEzYyc+fBDTuve7gEXXd+yf4O
rT0tYknav0BObfPUKlWl6h1eGUifVkbC6VOjnoesCCp5ZcOxXNM4daqbOVB2Z69K
fknMCbFU/qt5CH7bQASbpxddRwHj0W5EE6kujIpWbE2OS3bxSEKqTBjnuePUyO9d
QPfc9FDbXX7U054UxWvxCD/yOHPd9QLo2Wvy9x1EubXtMcPy+xpWnR+nN8rIqjvm
5FV82Rj/2K8wJf97QRbWNM0b63lgVUUqDZB/Bdrz0b7hQhNyh6weV/8C0dWMZKHs
pcEjXLPl03pCxcwZt0JZxsWgI7nePf5AtkKCVkyM4RZVxf9wWQpz7AMIl6NyLuKJ
1XD4598iwutPiRCgVBgUr37TtiNinRv4hQ7muJPGxmI6/uHAVY7/hiUzx1hfKoZO
Zb96YyXlmI4KyKzo6maLl9v+X6FlDSgsqmPhvOyQDgYaH8rKrLabEIRebwLJB0Os
diJRNKxqgNZpJmNz8T3vk40cnsHDDqej5pfuNw34Md9lefQHkOJZHJyNd7Wjzb0W
z/sc4Czkp+FpHApNfgZnEbd0BCNu71s84iPi2EQr0DuhM0+T7kCUIJknMBYZRj+h
gVLtvPr51OxHNxdRkdAfLHEy3WyH9J0T9EJiQuMPnxPWJCv4B5G0kvLpZNAqQvmu
6usCrcSmDoSHHSQkcwHn+VpxZv+PFGlL+ZoxtacpHcwuzyHkOgmfDTvpezGo1DC/
yGTX1uZePlAdqS0VS7dM+nfMj4r3QVHPB0KAGwiDYgrmlaPAPTK1vXx2iZbOMLsA
jvFPPqBLNfzZiIBqjTXm8idQzD2jJcxhlgv2ADVIntQEFRs0tnGUDZcKjvRRfyo0
+ebsqoz75bAgbIuPM451VHZkvyRE/qnxRRByNjMNK3ETG9ET02bfdBPedus4qgfh
7eC6ej7uD0moY2CfAeVKhudK9iGJ1PLYpSK/i/ydzKlKMip+9A1lqM637EeX1y+D
wPVLL2xZ1FL/py3Uwj0oK2zJJtw6vwjFmF8yG9wBb8pEgG1aAkz0UdgXgY9RCsIy
acHZ5C6DjWOLIzc6qHPGIFRrZTJ/6pL0wj97/sMbHq3nA2VB8r+KkEA99bj3DBvH
dDaC/PY3bhCMCm/mvTNMQ937jVIk6gKN7238Y1ewTHCqJQTtjOUBFFB+QGN8Px74
+yYT/k8OWrVxY1E/xAVB4MxsSMMxsr4VF7jhL22LXFb6+qnvszmhMYSz36cICwyj
acFjxDlL3zQ4JrAUIGQ6eu/p/mdwUzpcwqSd6q+BzxQrL8yY9rlQtjnpfw1HjR0N
I1hId1mAgdCW8pXpOOU1yoNnoh8Vh5CaBfl+IuT39uEPBCvwbEiw5DL6UuXQzJAM
eIJGGSmLnX5cwpwmp9SS2KRJm/DAnoXW9GhkunGRFrwYPpi2C9Zppd0BLQplqi3/
vlCIwVE20FcCmvUZN4gY08tSPqaAwrdDspw3YvNE9KgflWXf732PMhPtfHRGq68H
Ns9BjwVY0Q/5Tk4k2DB39ysfitx+tJpZ5IRAkFG6/tyiF5gqqPForgT7wKkbJaQE
hrkLMXSXhQIfPuXVSUfs85546e7irP8ephQWG3uTjLqI6EbeaL0bjupSn/3XmE5o
npTqUKXeh9EMYcR8RMH2uDzUiGRve+QTdHuEYPGHKY1BwIbhTqjCSR8QzyAZiwW/
DoJUNmjOa0IhaOHMJVm5lWfMNhnGPm0mxIe+jgMfa7ZWjAlZ9KMz28gC1SxO6sps
tCv2kJgn0izeW9nECnO8N8AbQi8saldbtKJmqeY4Cu/NMPfZ09RU+EdhmzIUGbmX
9odCEOH39BRP8h/NRwOqGG6f5NAYHcGuz7DRVbcG4KGjFqqwCBA0uL7U0q7wCkeo
NmKh7TDomf0QazUHSGwfYnDYPck6m6LBtYTLxLOrlkW25+8hkt5j6Hik0wMOC57S
IBV3EvGxMoCm8oSmIutp2WJz5k9yzh7l/ucW2ed+chTDY9QJB1PjngwBFc9Ww3yP
Yf2RJO4T8E+k1MkTwL6yW13gEm3chle5E0CMEZh0iJfDYFEPeq5tdexNeu38VN/x
7vSpmD0oLunfT8bfRuzibegFNyJ2WZG2SoiLr/8xP51ihuGCoesNHAmZlx10Ax81
H7e2lywQabs9gaUTPBjpVj+yNmqXWoveuJoh2VvLtl94bLvPaGWssvdeKvIx/NEP
qsnF+UqaUvSv2fLNZ1etfouf/6Wtv4EwqXqWj69s6RjduWGndsLIQOATJ9N1cSbp
wpBpM3BFzhH0Ouaq2Xj+8AIV1SRl34qSeddkvOG/BN2c2Gnc7Xe6Edzjh9NoGzs9
IcKlOCBoA9SjHdVLuRg0Y6vLC6ydW/E/KBNZgzLImnH7Vh9uHY2TzQxJAhAbcZTd
eril7E7xEsW/9Qtrq+6DmgkBhAZUZH+AGSagA6PY4/U2idKejq+OmIqANxpHCNOf
W9mTyR7h8dUuX4Jwnguf1Z9BJiDf4oWYM+7UJUETd4tQ3DU9aFUUDZ6vuj8yhLBW
Y3NWnQvmCO5eptGqYjoD8GVzDzkDP+RRdUcFqpqcyMgJ20u2+KZ/GmEp4D6a3wJZ
6e6Db3zu/l0DAjxattZcX+jsukn4FZczRv7icpWNbmclJov8FnpWLp+jezt1yn6k
TGhU+FMBQC4toyFdB6SUQIZ+F71WV9TIpRywUorKtpuXiJLeeN354kMsoJdMq/nf
Z1zMqJbG5YTZFfflPXX4u6z1j3gNq9f3KtQ5oTIJ7elpbgUyUCh2bXx0VhIUJH1S
dmwLFzIAp4f+8Y+vi8QdjRkg1hY8yKotu0h1IekxjIAVc5fog2MZr6vSon6cvX6/
sd6/CzhH9r/TqI3b5GsXajGXhb6jmciufCBlBULgRbGuKIqh9C+ZQjIkpAA2YPix
whhvA2Jkg+8xU6XyjH9JAnipJimXAF76Mcs5ouuio7WhT61ieOQSs2VAbaluRhIn
Mt/hiZIzaNUSS2kn8sGAt2xkAhU9ckBvPN7aiOa/e3w0sfy+E3tKsrQi7FZOsxOO
hG7V9v13f+6AW8aHszgtL7mhLVOwsmS6s0duxF7moH2TemnEtWv9gcLNDMCCS0xt
imCQqLW9+IW0B2Df4NunhpNmzzKSSbe0kHHaA+jN4z4TdYT3O/F1EZniw35iQIE7
cYDkpXn91h9JldlzGkdnS9bLtC+uVlFlwAhNGbxCpt1ipE/TdzkmrB94giB1od2i
QjEufbb4Ar093JU1K41dHEtE7BTPuySq0dx2ZMw4Rj0X3XVTNlPNlQ8979NYPPGD
oXeIkXF4KVuLaepEvjCJaIYsPmhXJ/v1NIh+Gy3VVycl3jfHGcsuOnRpSV1eyr/s
k073uM2OUeuZ/bFhsRYDv/0F79v1GGtwym1G/5RdExj0kil3uRKiCpC7vWGzdux4
irQbqs/nLpPbfItq9KrsOciKQZ/EB+wTJpvLOzWzIUNoqFCDzMm7PE54mEWeDvU8
lqxbJnnL6q3wVWdtrRImqW6OtSIvVMyNr0RSjxWQ3WolLPxHqQSVS7BWUZjwfYI2
a190TLvtiGZfMpRT0vCrQcJoweV69MEoRH+8uV3X2k5uOpKntVYSy280eC8Sxb2m
KbeLnrmnojRISRaJ99BZkdQyEpZfJfxmKv1nhxsd9VWpg6sx/XGupB/vmV0vvkvs
lF445yHdg+kI93vaoNj9baqe7RUKhqD4q+5AbeNzwyJDBPg/MWsJr5yzcNaQmsLL
HOs3L40tiv2XKx5D7Y+y4Rj+sFB/9Ljq29wFA1t71Dj2zEf2yPlFIMwxIy25JIS8
VhS17vbI2Gr//59OLCMSwtAGc188TeQkSuoSCKEntb+HVqtFpV5T8zDSXLTLjZHo
fvaIo4wU75dM7pb3yVBb7azAF4rji4+sh8TmaJDrLDK6S7DE37PUrchzlQSWXN2U
LZCKkeYYLf31V964Qv58RV7nT7CFf1THq0AUD0qSJoXQyrFOjMjPR+H4RGCwDnKj
2C6WRub5s9fb8TYIG+o1XvGacou+cPQYjwjAgd9TXzXkdB9ueiXBIbMwCMWotosM
0uBCr2/Shvi1nc5ld4hrsTMlhKNk41sHEi+gbImfd7IRh2K10radl1sDyitgZyiC
BzE2tZZKC4c+fBN8Jttr4b2u6qVc6c1S3g8L0KdV960ixLK8hYcX+GZwTJ94DEoE
6egGWF1+qOVQV2z6DqilOcG4QsYyCpUchjestj1CV1dfBX8ejcfvhXcRz9GwU696
0W0Pnkxwhhpv5I0E4u78KZWa2lUFg16Seft32gOFXtAQAmL0T+nqYqXrGCT8vOdp
rGGvr3LroxLMLq7egwp3Xu9fgbZeQhGgtsulgBARtWaDn9TWzOI1cVS11CxTrJI7
avFevBjMYkkwzlTg6frRn8KoywbFoSGAYq0Dkdy2sVp54Y8qLpNDD2+KwV9LPJMW
82WMI5E2gQqAB9Cnp7cai0xwwDYmgIHnrIo9f5ehIFVi7AHbN26VQzQaMpvIBH3L
E3iID2hjCyQpAGMI9Ra/FhXTo7WFCIObnuio55LeWEIFanxneny/dvR88pe/e8n9
GXEBC0obJGJUuX2o/JKpMJq88OKrDxX6BfOmn5paet9MEcH/C21nTw/aacNEzlCM
vDJwYy/gOi8HvSBVXJaAwmlWcO1RxA1MuHG0x6RecKOLZghLDdcDay3pa22KXYGS
qWGELuBI2cX0e5IKYpcrn3CC2dv5n/Qkml+qCYAJAmEk9DlHwUUvaVOHzipGLsfI
zNAWKg2itssKyQ1EYA8o7E2JgAE3kpOeJdW7eh4I1i59WKKVD+YkNe38flYherOG
xAPlMrW9053YgX2jJX5yeWU38TqlHCPnldk34oDX6jC0RW0UiDLLL8b7SiC6Jg9l
bbp8K6m8BPha+WUboF4ihl34ci6c6stix4l0ZV8AN+xtySZb+qtKdHBFqhTgiOce
o/Upb+WqK8YLgXDaZ6XADo5d04RIlNCN3QC2DD8dPADYQRdWwSZFuhlvIk+hdB8L
0SLQ4sP7cyREFKI4Gj53W7XrTb7GcfuIZh9agrN8KJ3Brhur2GfLHRRxwJZcFzJ6
k5T8u4zQXpjDyivYop7nIOSiADTakRotiIXlSMftph7MPfcgsVXmwRB9hIpXy5PT
028Y5Og7z3utzTRs0zpksBoR0INRQHnpXAGNLOnJp4NaElY/LhGLvV6pJQcXZ4Sr
3BLT/Eu8IM5V61atWmfwUcyrxOSl6Q+3Yuxf30ntTvrZSzRaZCmc3VtKElcxjHqg
rYvLSvjtfnd34Q03j0Sj5hyQYkxh0iMips17qSiUlFnBejcehKdJn11KwSH7xIfi
zNClpErMQ60yCLP4pCTqQ66Y6hm1SLg8ZB3jXfKZL6FgIIxRvOh2N3reoWtSASiw
/1wc55qQ24N697chB7wM/r6D64vzGiCwhj/KHQmXWnH0Kub5ZllIwTM+Z7nYjRv+
+vgrgpIka5MNe0GxkLX6A/19EuxpZ6BDxD52BiqxfRhDk/XxlFlVyrkProqh2mn1
xRTqy2gPOOx2iPsoiJgdQnU0AliXmzj4rYrWw8PZ3Bhtq8HEqQ3WBbkxp8Obhv/Z
2YM8Lctf9/4bdwe6wqFuQ1TFu4mrsnQIgr6188U7mThbyVAAgn68itqUyBcl0Faf
tEus056Pzy9din19eMHrAgxWLUa5riwwCIgAeDslIAnEU9nZXGyuTRrof5XuHIyJ
AHpxDfC+gsUEY3S8P+VWUkHVcvZFr88Qhql6B23d1QMi4nM6raZq1QnpQl4kDH4m
Velqs2/RhijW+DbMRcnvAv3cOmUAxNB7akz0PovX6YzhCRZPCgQjCcdTK6KdM/Ul
ooRPZbKxgT/s6WrukCWZvkKDlC3hMUXGVRA/j+IU79e56+oHhTBIL3SZxJxK7pQ7
zYdt41ivk2+IX7UORk4fLqyvqCRG7Qxh4nSVl5WmwoBHagoAufYZ3gxNPe89jU2i
hkhb6jv7YIjoNUlozk+buq40eFjf3VrlGAPLxriFKyRAibbMbQlfcy6Su9ovW8F8
Hb/TeebDCn7Kzvl8hgMbk4hbgrU2RyFVkb2vdFYekB6QrmV04lUhaLSAPhZf68kt
05u56CZ31PvxisAhdPvHwq1QZtR/XaP0fPp4ne64Wl2yoc97dbnqwN2TC0qA5Kph
hckvYdb55cyPQ3+z1mG3NnPZptuhyKcpVhbVATzRvRRT6ym1wAQM99PpimQuOIur
vHJJsmfOrqr0OBhLbK+VW1Yq5jnfZHdvfPEKaY+Ch0ec/ZkvWYWVy9gbp5ABINie
2NDQUEYmTn3PC3FzzlzkSKix0zZnDGmS+Sa3MTt+TC0xTQW1m65jIP8lmfE3IP6u
ar4EDQkVE122LuyuMAtzn5Mbdfnn++VRzLuKiL4X1WGnB5B0zqPQdY8LEbqnjJiM
AoW8GtgO/8yFkKQPxDuMm+w3pEg9Qbb5KZlt4745BRQL+jFvfD2GNFo0NlIIOdAn
Mi6LqrwV2NxWNyx9XBdfHLRAEConSvyFkIBx+LD6Y3YjoBIm6mpVbJ1WhCAIb2XJ
6BXz4a2YDooE6sbXpeEQEYWhT6fhHxh2/AOGuhruv3MDP0NAgz1/dDaJeD37fw2O
dBkoYKQeOnz01Ruh/gNnAJ7iwcSKMir3sDvZWo5gC6o8hYK5KypkeFZYsw6SeeJ/
v6q8FrFgPJBrgHBiRqcXGrWjTBp2M+O91IDOYXRU8rUFJak0svme6gvM6b26yNme
6j5oWUQ1snGvSVuJeJoVTdRws/U+SXkTZtF/GbogkB30zJ8TNn4B8KCEiOOrkwvo
zf/IpXJoKIMP+kU4MYfv9uFVF1TO/vxoaO6pAbW7EcbE+fylwa8ZfOGL2UzXVbZw
0mmu4K4WpZfbutoms2qQi1EDs1PSKXkWaD2UAOeKqbPvkiwN0KwtWRopnXlj5BZI
ZXJ3BiQuq2XR6SAyQwHJ92akZ9doruaX+GHQ17vuPsWxW73W6B4wPI7UGEU7jQzm
dPi+71WbnmnrJVbUtCeOcWwtnptNxhyEERRWjgVrbJ2PMHRp8J+FnXjxOamqam06
37GKVIOQeoJwrdRslO6eH7EODDDMwFzon8pvWlN02au1vm2vLXQm0oE9CEvFypdn
jNXLl/5kaJJtuewvvkkd0ovUHaUgAW4d4Zmc0VdgPkRls/rFKMag+62kDTgnrMOr
9auTfYidCd7l30lq+9lsRxoGJ9nJPG+IAU44jx/WrfsO+DaYEZ9oCix/Y8r3ZOpA
SmX5ycULBNvDg9WLkPwQzYglOioyBckzrtFnv4Zf3YEEpUetV3wYgFBu6L9IUKO/
49WXpa7+R9NvBdTvSCut8P4bBUY+9CPCh8va/rX22olOemH8gChY43TcEmvenKqW
+LrhjyYwuaHrvWVAEo8apuauaLLX/DZymJAmGfwDW9P66XMViRZPN/pY3gptYhf7
OfaemZpdNTkMiUEgSojtMMz1juOE9jQWnEO+CIBDCsn98Q4USG8LuHIq5Jmqnp+v
1hG7EM9C7TF65uS0swDEiVzWgbpM844T3Nto60WRdZUPqoaqfHna5TZz0bxSqF5M
QzVsDcYFJaNXBN9R+tUA0BBX/WoN1ugzgORakf62JjxzSQqPAzUAMMQtBliy2MKj
zx8HBZv9/la4+8WyHydd99bEjX9QizY4gkh8n8zgpGnSMzj0OOelO7IK0BXVnlo5
Yh48wfLi3nW6VBlZtieKw7hm/ehKGRSMij96zTdX7CX2jhrLN12oASk5KOiXMDEW
++e3F0y2JlpmKUwf8q1Ne52BODupqmKzjdwfGB8OUCVbUA7hq/P0ZLI/brBCqbq2
WMaBBh1d5yoMR9ey+FxY+cjv4cUduJpcr4BErpXSh/G488M5s10ApuwfaTm/5EYJ
s8rcf57aRRuIFl7id/49mr03464iv8q8aLvFGfBbyCHZ8Yfjmf5pSvi5pKKNn+Sb
AakZPpZV9vm3SwuAWZMhxMIzQYpoJYllOb1alqsqc+XgmwPJHFIu/gw99vrFLuhd
ENt/dOkuEQcdOvpHNnQf9twRGsKLlYGptSW9YDjVE3qW7BBhhBqyYw1L8zxEe3uf
vR73yNLnNtasXSOcu1+SliCWRr/KuSer5sCpuxOduCctLZWHk3hQYNmJtPCEkt3S
XKOpQo1pvFWZsdqNPA5sGnn0rnCinAxUfD1FVUW5objp4bic5KwVtGAuhU/Soh5F
PbJ/HDAISMdAWLMDWNL0WzgN76NZKgzGQovOgOYyUeqs8RaStzB2IPaWxy5bSD4u
GlLhJqTxcP355jxZchXAYIMWFv+pSMQ3CmtPv54TvFBKY5o832gImqkeAidUR0sT
yGAjvD5GLGycTKonmOFCgnno4UwErgRD8l9efBFygjqpsV/LhHKisd4kfHPrL9T6
J9Rkv9At1Zpfuy8iL1OgYR5G+718QaVjP2awrxQTAisM3kiiUtTz38OrtAU0JAgP
HcQOn+ULt0WYFFL33tYQ/P1sWdBXJJm0YThvrS74qRpkqiEnX9mVsRisLLnToVQv
oFW+wvm43GBRVd0JqyqME4tuA6hRpKTVGDy+6DI4vnn6kJZLhGaxMqn2kt8nOvCm
DVf90M4w2riQ3KfWLdhEQjbJDzuyx3GQUO1+JT3347BIG9pcWYPO7FZa1hVxUPa4
QS87n7YkYWWc7zn6rip9hYpcDYLbhQCtZGr1cXOID9queyG9mO85qwb79k9gdsLT
L1YspsVuQFJEq9qJPs0MXEtpcchPX/IOSAAVjnamBUreCRvftwNJfLIu5EVmxDJN
GVq+Chn8m44FHpalgYTpMB3oLMPT7IMmJSiWyKIlv8vV4ZTh0/GwbVVNuYa4eq41
Gqxgz7c1YKBPVB3hCK1uFfNuTivi/nmCv3eyDGNZ2CQfbWQj2XrlC3F4XT32Dqvr
B/pE116XqILXKdIa7rXH4mWt6gfobmbteIhYQDeb9TP6GXCehwxEM/h+p/GBgIs3
H9TMubdKngre6NdCCCzhRjOEAkugXf8/2DQvaLooSoxbaBs/zYuoF+LO5T0g38YO
hh6Lf88vkMF2mRUME6JbVF3y8SQ9l3efiu68llUKz6YtcYPU9XLNDos1Qeei3Pcu
w/oJiCY4AVJF6IHICODL/JPmmQArk3K8vj7iCaC6YWJKRXoPJbaCVDUVv6Y5EXYS
hC4NV90Pe7YBgvzbD3JRZ+51rHIabbVBlPs8GfAdTAGDetuxEvr9/xUofF1m9USf
EYyKtG+cDhTIfI5JSz1Wo+Y5407FWstU3SBA+hOYvFptyE7kRmmY0YBVNnpPzkub
pFA82hIbbHZsKtcw5ncoB95JXWEUGnOXiESptY5jWuqJ/+8+fmLa4Ivdwl6lYDHd
uhfEaPfmpRPcBkBCTUgmA1zhydM9yhwGVXkKHyZJFmBya6KcK7/GRZLc9cQe1zUE
k3+lsHiEA9ihj1nbVc+xrpcx0ejkPa86+EcaZqjXqepTL9cgod9zkavOZIZ+mCEz
fAZYuPoxtiCbXo4AE+5e2Qq+5Cp3mzVln7gizEg/oYfACWfF6W1/wwBumRDU78R3
EIRfNeA502AgDsFUAQeyZvNn2CqlqynJhsdnyAg5UPvc+eaywYIs/39nRhzDQRBP
/ZYkVneMeVysdR88DgPeOACVpUofV2FSqTgy92QQ6CWmBmlXzP17tdmxzgMlXuaL
fiNMzL7wVqzgl7PvuOttbM40cXi3BaTliPZpEL63nYzEU+OvqqTMfioaYpjqfw/m
JLnYLeZGZ+1+StkIVLehZ7fZrw223sHeBcPm0j068Oc+50KUWhj611Q4GebzHCP+
w3+Id8YNfKP6FqgBEdgA40cr37vQSC4zbfflXFSG0v1zyxgd32RbUky+ZJCWs2ut
JloAqDB5dBTYQxIiTogrQYcQFqYcSdqT7juTgBTx9MBIB/G4IoVEKyndaebnnlty
VVRMAzWyZ1ZB4OvKA7bPPtIsu8X8WslT0O19P/QnqUdU2S4tDVSIJVLab2vGlGQ6
m10Q9Zf8+hUfrP8LzzkTPN+RHvRj5UIeCAN5RcFM0PEjF4cQaPFUKrUVutn7LIXe
aEpcgoZfdPl5KQKnldUixRF0kfAqZ8EJvoDGCERduWYWd+nqFN7YdXgxLKmYwUD0
gjjDqcpo7RpRlWqmsX7ocxwG4zHuZ97D43+l9JqmbnnQrteDyDPlOp/Lbg9N6O5w
CJOc/2RP3CHvlcwSd3BqJa4X1Ms58hZbpAyZm4PvJ+9Lo98Mk8l8sWNXQpZs8aPH
YR1fnE8X5hqRynnapSKlEi6Ev/RQKF05O2rbS5QRncQqRI16y/KU6hnZ/0NHIYLB
4F+aLTJWgsjcj6dFt6ToWHEY1nIT0ZKtFJsFParSihx4xn52IKsXZybu7sEwbeJX
aVWRG/dq0rBKWWK9i+8XOg1FMJzzy5h+RY8LYj07cFjd9Ze8fF8nPtacZR0vNaTX
B33uznK+LzOQZ5gdlPWkxgbduUDQT5FrpOYMIYry1EcofG85UE01eWFBgJZsKnCQ
kEr833B4vACGULim1S9hnLaVspZwqGeOXNo74GAcSddP5VUMZxhOGWRxWhldjQ4K
OL5PTWhDMJg9svqpy+oGMC/kCaWHm3r0+0co/X38PtU8UL+AAImgv0W6lO2flczW
n4WpDRIsHJbbGOk33HjJeRlyd4dU8wBQbmnwtCGUUIOMI3+gAFu46gRrorqoQjMg
7iyBxtmQUlAxaajPA76KM1TkbXzW3wnJ+mcTzHJ1ao8Aw1yFuJQlAmfGf3QQi/iV
vaC9x8BD5GePwmHPe3ZtdUxg/UMjApOj2NzkS85iFhk/lW1I4BOezVSMra0iBhJ2
BR44SiAuQrbqbou4YvAhYzqK1hcCp987+2WFTnUhR3qDS6dPg8R6NdWFzZgnN4l5
S4briGknIq97X3xUFNCJONncNe8KTL2cWN5aVyeJwwsFXW+plFXcAof/2x/q7t1u
Pydl5bTqiT9PUd0Islj7zXELTLeJ1FNdt0P9DvT0xIA3AHhaayScdsC8Pj1+si4s
q6nFYc/0VpVoM309wv2PkOpxSwyrtycU4/gsmCOjLM5KEJZGSCWa5IY9CpbFEjdz
DF2xVndAaiC90SLrIW4/xOFw8cwufXeN2RBn29PtgZjXggqWKVGezQI7PH8ti10H
2XK+rKc0Vq+fS/3UUFyo65rwJbqjx61QGprAPJ6PdjUBvEjc581YlAhoiCBTVxHc
IqYReghVNsQ8mgMggRLtpbJuG634eAdPbRyYHVUNhIz97OBM3EKoWWpvQt5RlAeA
95nsgKtCzeLjbITvPWZAwP5ktZv496gzviABkgBeMsRYms5WxaPbY+mNZ+n4rEaF
ANmIyfvWlYqS04QwiaqNSfK6yz2ypUafToXuWoGHnobs8qo/hc6KO25eKIqcpdCM
QGOgBvqd45odm0GYNeXg88HjLYkZtDMIM8zc6M29Lc6EWZzSdN1/xckAcKoxvBCC
IqXurjhQc5QvhzaJPBKweRoF4r6Y+fmYrUA9yjESKJU8DpEDT+1G98LbR48RnWn4
rlgbTceZOzTCpXpPHqB2xaYQ8twthEA/P/jZgdgC3XLCJIu8uBWp4WfzIKQtEYF/
ZEm0M1gBnaUIb/T79FjWbREvErBkHv/IWglDy6RUw4WzmU4GNl0nA43ORaJr1sIb
Hltlg3tV+T1rrcu4/jevnxqFaz7fx7mYdrr6FT+XU/yWvZltRbQiZ0LMMIToEnhD
As19ZA6vBx3UdAMFRCJE4fNKyw/Tu96/Z7uEBgZVwJvxp4dY/fwwgZY+3sMOHSvR
Jn2NFwSCuISI+HKmJGdVdPZUapRCmkRF2C9RKoHmcIf+6+d7gfbvgdNOCpaWNlmE
pu1dHN41D519P6QmbTio07svWPVcqbfKA4juab3hcbzfwGZyCTu/DOE+yPIHS4Gi
aIcxDsUpx6icMqdNEKiFDGqwcFt2YsgTGZiNX4te1i0x5LrAAQC5NjOXmmZ7f1tu
a9cZs5S4kqL1sSbJOFHd4aIofl0D07yKUSLdQaD2q8AJgDp1E/5G5DHdvyipHmBq
YfNM58DZD3OzBfHiaVfpFG03+PHOsalYHuJRo+i975B/flxqhWuLaBe26khSu/YO
aQB7qtmEP8ECJ4pbchht8uZ8ozBYpnDrHBlmN2x9AlYI4NuwoV9bCP26MzNwahdK
EE/LdDNsQ8rY40PV8Ai1O1CBmtA2V0O2H6DSMAMTG28ETFTjJkyNU7MYQ2pYOoeK
h+fWQtls6wcvbMM5FXOwrAFSFLlsXZ/XaeLoGYn5O2L17qNjde8p4LDtwDnQJ7vH
jtBSbVGNeiKtLNVrWygIHGfE0CIr4R0QIwgnJu5Banb5S4XsCaV2eC7BztrB2xIN
3x3o/pgeqDNFM+l+jmodtIHBaZV3M/Luch6BBZlSwSyl8Uw5EwHmwAWk0mkyPIUs
s1lL3bGGsWu4LQjHKPOH6FPpBCvv9KqkBxHCD4k79KAFfLSWEPYiOLJz1xIoliXY
V5fcqXEzkXZnKcXi5FQDCTT3/0mJMguFPD5ovQjz3EyPoB7s9GvLlAx+zigsSY6z
62vL+SIEiNnF9hnugx0Qd+qDoiemROjcjgN2wcvMXXA8kcfk/WYSXv5ytYT+wZbk
Ilx8/zy1whaxmFbRqw3mPouEVh9JNnrD5JGLZCBdq4MEokfom1Ayd6uPEGow+2o1
rkh4h/Bt6ytduX2XrlxLJgSgVvAyshtJPSere/u2jj4+VdpPUOzTMBZ4sTIKcOzc
rcMR7Czwo6kyj4S+JOkJYBw52K5RFvz0ULKdqxjBqSIkyttigeTEz0Y3F9kzq0Qg
CpJM8PGcjHf0xl7ii/3v6+FjOy4RFPNQu5NE6avOL3v5rzw2bX/fMWD9THLIGj81
WcGLFQjj6VCZKOqtxCuQk1B0R+PXMe4SSoJwAYoQrbhfiUALrqryuql1CNNyBNPJ
PsVN9WUVTDqGNkxpNHVMCDE2YOHFZ/82Fd3p9zYMdx3vEEZQGVTgGHSGZN0I1ja5
GU1vPY6YNXKb31lzVU2oKk5q6XFubBOEJ4Om+H6ZIYpO+wxgVdbbppu1WxlzRWDc
PHUR/aXNnDXYBTFmyPxW9hmt0pAUqAFskU/i2YY/CyeGuWcPQtUE6EO1p+2SIegW
6W8PqxxK8hV2sdAnCoQfaQnlazQE1/R/PFB2J3rnquSN+E0C9vDsvZmh7P15Bxt+
xQdLWCByGPkXEN/sFhBBeDPrQBXrucb4xtczvCXr/V2RZBImwgERKXoAKq8HLNtG
w2uTeZU/jW5zouhrWCF6Etq2juPMPyTnMu7sZLAMOHYyvKxXr9xh4JALj57PypIp
tC8JH8WXy0x+tbEJeT3NoZ4znNLzVTovrBJ8WDe3gPlHsC6F5hj7iizxExIXYRvf
s3Zgp+5lkkD9UEffawhhclgIbw68HYf9ipXdc2pNumrRCoJHlH47uifIq+TfZdKU
Fl8yv+jZKRkYFStLJLWj/MxUu7e7+IOcKnZhjmIrvn8APc6fSw3avTPeeFA+J7AG
hopFggoWu7i7qHsNwzd3Wu1xKijInDo8rN61vGRrCytJTQMlD2/ISnp3Lq23lS3y
oUaGDcTHh5Z/3XCmYwRmieKN013X6XwqxKMkd2crPUi2Pxnw5Zv41jZK9V4w5IDE
XdQog2yHtTLAnk2N7nVQU6B2FK9+JeINI8hoosJ546aS1qHVKx8JFqOwbyvSOd9G
C807O9YKAn+ddWq1Fz8bLJw3BbCIdR19z6eSGiSULVRGXoyas1jg0g9RE/ELQAL2
sVdJbnyqsn6NbWHPWUpsK3tEHnNrqbvqHXi2KuEoYgkmoyduR+KeZEvsjpASEDwE
XZbf9AtzpJcJ/C8k98le+ZTv7nOEGrq12UC9i2vve6UOMZJX3cVpFMOmrcPbr0qn
OcFEhgbzDjDNuY1cQhd/TE3EWL4G9dV4F90WZsu1d5YraoBYynIc5Oqia8znqHSA
LMzXLZdBgIMqf8KhSc7JoRNUBMnJYEjbeT7NW1qjy7V93bsnAVi8CrdSfS5kVy7z
cow56DjFmdniv8EnAqYPwVxgpNps1/CzvsOSBH2JBDDnVpQDLgAi4wrmEZWelTAG
fe+6Tm2izqLbpGIsPWO1drt0jkjzk8dPdBLhVh1f/Ac1syU0RS2PzD/lQBwMqMv3
q1aNa7dwAfMoDk00B8DOQtE9HO/h0eTocXr7+THUsqYE6khAyLD98s1ogLqssGEH
hGx95OMUsMCBHZqHfHoXIUCa/0NEQpD0/UUNc692K9JWkkPWyKlX+1gF0DR9F+DY
uGIB7mvoMB20h0SnWrfkWw6C1u1UFEbPdmV52Pm8aWTaPcoo7TnHrT2FjAH7tWZp
XJmHMGzCeO99BANb19j+a9YSq9+V6qYoVbBwJbhWrMRcvIaveYOh3C5gMV2GaFmY
n/9WUD9h/XV+42h0HmJPfyge/W9bsGckMx9Zj3F+/kZXxaWLXHzlmNuu8Sk3ZqgM
nAxMX9mm5TAit5jnkR8dzFSIfwglgmly28DaoSU+Gvs7d12Y422w+L7wyqGgS4ME
fkYbbnyKegQwtn5NcraC+R5CCCQah7uP6Qgb5+RZ0Mkbo+Sz9QecA+vHAhkVquWX
NikHiFbJU38yB+7paTO31MLk1T2YJHWJqHwx9VCnoK+VIatXIkdjdAzGa5d7rRD+
I1thhe91ddtZVY8N/J+8zF3lz4cdkFzhVOSJ6VMYdatBF1gK4YgUIz0kJSsRdYyQ
NOw9Jc529ZC0hQ4B1fZPL8Fmmh0KO6luRKmu3BDFKi64DvQRUQVDChsVuRfYUfL6
JW+ULf8PrMKB4QFC2sFszLAR5J6AiqF6p7WyWN1PsYu9P6S753Tvq2A+rojmm39N
LpkHeduNfjFGhjXq/B1pW73LWMhKm0sZNcwuH6CNa/XsrI0zc7itjXpTc6QBGJMr
QHbAHOEUBKtsGbpU1nynPFXSNlT/y/VS81M+a5X6dRlopkkp9KRpRWma+eA9Gc42
q3ErKSUG+QE+RR5mMWQTd2ycCkUKC4G5K2ghcRlFCXdZkS3rlSQ237P5wX9md8O+
pHgmUZONdfjMhD8msC6jMlD7s3HDEBcVAUe0cN0sI+m+9Q29WeWzfZ60nCechGSo
KeJ85LUvxlz6/mOdMAoP/EEE7q8f4Ng7okj7U3yNBLHB+6mMlkGSdReugWqJ9Jtj
VFAi95EP/WwmzHGoCpVjynjky0WiVYKuM6EvDgImAkgIhxajZfzv240NaeF2b75J
WVZn9n6MS+GKopVf2dF7XuIWN0FbMs/1m9N7LGSA0FoKP8lxKpiDxewfnPLmHRIV
XBKKpOYhgE5mrYIXAVpccoFA6wHFfzga5r7kLMfiYqzkqjdetflFYwgpAkWuDWBF
78kqUKmGE3UOYRP5zENJH13tcNa8i44bZKvU7Ap2B1Twcow9SKztJOYxuUZ/DERc
cVAXll0uPm0AP9W9iV/f2uzFebgyjPbl2Id0pirEmkNz7+AQfdWkYFbZINhnF8+K
npWNJbetiTiabkBJifqs/R+jPJ/3qMoO85Bq36WSjF5jxpiIybTlXa7o7V6ZYy2U
xabbWA4Ju9o8NijF6i96U9b041tA5SMXytvWFDIVzAcXK0v1AHKUHCdpFZ4EHHj7
D75izylfFSgWkz1e9ZobKD2ekLsr21Vu2CzHnAwKHc3QWUBBoDtzxSUf3tVqGbmR
hpAZ3iF0wHiWhwi0TSwsb/IAvLDCcySxjKHNFvDNZyCBPZzv11+R34CwgCu2rrB2
NOjU2X9gFog9dsuTUkyVU/IfvRlDrtxsivIj0hHCxZVwPTyJ1fvs+RTOFMrFRgA7
0pfou/OwsZVY0BjPdbh8DpJyDc/ICMzeX3X/3tRODKcI4snNVZ+bV3ihoKIen6JM
sWCP0tk0xx+rw/go21IxQgpOTpby8jpQK2uS7Iu4ypIyOtOw2zoqNI0Tm6AmZjAy
0wGG+m2HUfNPgAKrx61n53PyrAX4hi1f6NI3DDHXSbZUX5YPH/HxITRNpfkb8mbh
7Zp8o6ATPyHbw+me/u34wXzANFVR6FCFt/Hpd1k2nsg+G8MZmaCoTr6VQ1ZMCPjb
z568qoE64czgFDTH1RahIWe3uQs9AqZDDwXba7QOxiq27kRV7jrsg2F511FYfQWw
CawYDY3RXX+DuOFnUdsI6scwE3HwriucMSNfsT0ZMbwoqsSaKkQFWye+YH0jCkAZ
CN5AJNdRqEcFkM6bArUkz87DKEO9zp2xYUa0fJbcvXWUjiLXioY6PFjsIplP+/SA
ueCagF+DLFAEOufrUPrpC36kkk+8GhU+PRz6TPh6h5KTmet/gF5jPdKbHZie6InW
iLKivl2d/MUN30uSVX3Dtzm91LYliE9yUEJtAq6Q2Rq54FZNvAiGfREhhFEVzUMn
fWT6PiFLMirruUYGEUKfzA3HPmMIFppEG5jbLnHisOnrVO72jqi2pTBqJH4oeW+Z
8lm9kHwSQOnvVtyami7H1sX53porEQmvBU1FpJ2rHd5BHZCXzeCbeUEDkR+qa0lh
PwIU1kW1YOm2jqwkQ3GXvSqQCXPKZmMRHgk/3fKAf082+4N5QPSr4xCuUqlW3Kq9
Be86/ecTOGMtXRyq5QACYR3Y1fplgPn9ilmw7hJLOr77yx7Gq4F/DmwtHI6NsEK6
cBDvx2GpMcdMors/HBWno/CY6pLeU8ELX3Hjg1e0pl2qmfoI0Dqf+hkYbHpdHLER
m8katNPMJOjLn1TBkGyam8zlDvm2oKCTM7tU5y6pXEqoJ5mqYHDkkC78E8tfM2DH
ViNow0E762OklIhqDZzvS+KlElYt+mKd/Q9o+BavtKz9w1GHZKr/OfZOhgyvf2pn
Uv6K20u7ubwhRPd82IbCA1jFB7C1nRO5XU5da7XP2pe81x6ffCpv2Ww6wZUSc4Fh
h56Cf3rb3XmzZRKG5y+8JkeEFBkSwGIpsZqcN3WLes1fzO2rqetZ4OF0UFdHYe1l
rhHnAebFoiku2Sn7j6EfHIHXDnLvgPmOs/Qs7HX7fsnKOs+ZiW1QuWYtf/fNztdW
E3Hkt2dbB1Mcs3roPoosag0e0JdF5t21+/BRscWBjt51NPRURBkGykzxyDOuq2Su
r1wQywykYI/VeauYIPyKM0VEwamiqVmPb1hZmoH81bdWbrd9SGBNZNyCkyONdSPV
0FrRuMuJUzcLutVjsV36mxuGF/hFx/Rth573gBaCxLJbTfukY8kQqQuBiLyTCEW8
VaYbIqJ8SrzMd+O6zZXC/U7NoflM5LmOeol3ZcCJwCj+j3IjDjVBrh3Y/UiCgIey
anKTwZYS4ogZv59PYaCOPM/dyK4D/qqEu/7ONu3xNB/GAORJhbgFwOnXPq/OFsgd
iEd0LukED14kIT7x3wHGm+smMwko8ubKmW12S69RJiupZ3kXnTrYOI6pCHSOm8Xt
POW/yE4k/E7JiNLlnulq3wGHc/uFES2qn+TNo+OXGjDGGPp/HwStfcvs8PP8ecO8
rR8Q1Jju6TGOjXETDeScKahHirm9lHpLOnmzw0ukf8UIE4DoB9iOocBv5ap5WbIi
Gn9j3rI4MjOJAfogrI/xvs4oK8z7xn3ywoLoKw5Srvwl5Zw4Ynk5s2p8oafl6N2i
cKR6HbAv36j5ea+YUq3+tZSSdF/WjM4FegAwCTBiSDjQ5/QsZhBaBxLXzRmmw/xO
Wqpn1jjbdUkFsYUl2f4HVKwnu8YhWVcaY6p5tjbdfGhMHLtIK7EqYetA3Dmi/Dpr
+hNdPqVpeyvFD+Ed7mprzTbd0uDh61jZIqA+Lcks/gBtHeuKRY820kbPpfzSoCeB
iFF13NgB69UyHr0Jds0e/0be2EPKLC8n/4rBQgrIpycQYk1vGn0JufZA6y1IIITa
bZ6O1rImBBbiMCFYiGM4j0aIqPSQZRRMG2ckLIDXGBhyZOg6S16NjiLJyBvXFVQ3
yIf11kOvPu6wYk4a9ek3PN0Y/7uXGY5wv1iLWZhYUaBq9sKssHTfHdKNrBiFy0aK
nXvflUXiQrcvYFolP1AuGKaGVW4nBOjlWIGAv0H9Wj3GpstLu2hyJIQ8nNfBRMTI
7fJ721miKJPLyHoQ15QX6lK1r9rInT/l86ifmFe1u/DNU2xKiJscsW4PMEWLtHwf
h3pf1H9gLtUePnn3Lbbvz0YaELdkzI5ErBcLKc/cTpHM45tZ5XV3jslgD3KcWzHu
JqhlLzwgW9n73BWuLB4Li/oBoRYYuNfMpTe8lyzTuH4v+BXy/oY2S10XAvoGpKjW
qFOasGrZCVeEp1A0W/JFi30YB2Ru+nlCqKSsgCiClBl6yeWVzxihEtIDVaHUNev/
M/fSgHBRZ4A4qwFSDRJKezg/H8hmMwRC2z/o2r4Uv+rMTvp8VMq+1KHLcNYbY2TF
+ExcKqhULth3OCKhvpaO11RtQ6MfbiG/kmOTKL3f22dqTerCucDCBFCkRjosUnhF
oCBuTMG6LQqvuQITJfYvU4kylT11SLIbgKyE31ta6I9HYGmrtqQcOB8SZvvT/BfX
XKTTqo1e6tRCUCr1dIv4oROXVIYEFofy5zk06GaI1bbY/isvcH3g1zBcP1kvdNcT
n6HKqk2hC4L6mExMj6xBk9i8OCvhN4pK0cQHLATDiaVquCvH5zPascVwLaIk7+kf
azIniMnGGK9rrRs6sQg1gEX99QHf6ueSe+pBOG3CmdOk2qahnfBgR6iAuFHjivhZ
PmiutbRWnnXC2WVcLacUbZ2G7aeXrtcx4FRMnqZs4aa3QZXYuAkKgxGYhONKReDN
RkJl1RqvMGimmlKAaZn5PEOTJsRmTIBxC3W9CgPrekjwdKUa9zrDy0VmA0i2EKn6
ingxlQHZNlApSDaLwVeMLyA5rhlvrwJvxakVv46uFPq48MGHc2vnlGK6PCHA9jn9
bU3267uctawQ7IqrlUDykmP2w22JJ9jrKmlt/hCCNRoWd+outu5PcfFV4Y22C8+R
XmmDsQwd84IOYP4PAxcPOaIuVBhaQHr/j79pgLuhD1stc8EuzUCLuJJi0cVc41AN
/H0ezuok/4qvgtqW4YCN6cSok8qUeCKoU9F0QzXzlWSdkXzbtcvmzF28JdImbI9r
6/2KC4sWZ0GwZYwa7TUZZw8WCTehi9dsLVfrxooZpnw3unQPIxlm3jsOot4QM06t
T6vD1Rnn4LMAFsK8TmFY5Q8Qmf3Z2DvqONALQ/h08HFGggyJ5dIDayTAPk/N4KtK
QtDlN42JxMZn8PnXVRAaqqcrCupnLAqb3Q9Enr2doyGCoTddVgL4AipxK17/ZpOy
da6Au88vQJvrRzHlia5AjhDrj7HDGTkDItDc1VBQLCTO9JYdHf33Kj7J/620A6TB
iYHX9DkMw/GHjmU6n0ZNW6BT38iwuMdD39jigwNyNdtxRvje25RCWOSA1cPmxgV/
DxgDHDRmF1s1wL9ERtiXYnlfH3Je9oj+r6TWVD/QumlGST4xUeGsxbeB+xY9FMyT
hi7/ocCWlv3tPiB0P4tO+OVWAqjDUAxMpmBCxtVivKxf/85NX71t9juoRpq6NSZX
SnfcATI/5lvnx2nAlu1LW+lt+nYH3mO4fcBg14I0qiHKhJSN8G8twaRYeGTEhpCF
Dj/tUAioyu+vxN749t7rja5qo+WqehUm6ZLwPKYBw1oEA5phjFYxYuoDnVmtRHnd
uMYxRCE2ysx2IQD9H9xUTj7dGk7liEvAYLVYfjmYBcP3zlHij3JbO9M8E8QloLv/
U3ejldPauJjtUBC1Q7MKnP/lY6rOKF2fiJJoX98TWpGd88Eo/StujdsAox5h6fO9
wTF9Ij42ApDv8qqYZMucqHvm1OtCK7oXOGYvHiiBReV01//ZrbBqnhN5IQKkb9Um
ro6JJGIsf99nrXBr+Wn/6aXyw0ksqmTUt94DVqiWhJCwmD7h2myeH7Vm2Z0s/rbz
F2Ej1AlKcgJjSkm1jkTzkAHBHLyRwKkBviXGaQ5bbTtiGvvb157BsoKl9VrvthL0
nL31x0Hb7uWpdcNOQn0fOVOj4IEWO1PnvpHub4/AbkdPA4X8hbG63BRUgWpVSrlZ
WnxO7/RVSRppBc+hywVluWcM7Q+Ah1Q7LYPWtSiRScAF+ZtubErI2zOgmpmbSkOC
f8WbvM3E9ClLxfFGfHb4Fv6Ohvia4Uo9qzX9JsuUhJFoCvFuL2XFWXNoa1yusKqg
86JbACA0uZHABDw9j/d4bSs+LhCgUgT9YD++x1Z6RipZNUUP6lAmdU+V6OPJpKT+
RFM1omkZID8OVTHgrPqFViv5rqg9C6sBC3vHFn4df9dYxcfc3c74KJVBcw7xtS/f
hqHkkoUIz3vbHxOxCjCYOWL/oUm9xsTN1LuDpJyj54HxGTT5teL31oX3a6Q8H7A4
LgqPcX/RsKER6KqOSDk1x2saPOlJIHoBwGrmMvTYUY45zTrnyEEAYag66TEj2GL5
hnT+fSgMslXvDZuemhN7dE8fvxiWQQppHRAoP66vOefiOow+9W/vQ3jykyWizCdJ
vjlf4iL4PMM0oqN9/NsO/tZXWQus4+6NZL7X4B6InJ99Jf8xp30ZV7qBwshndCsT
xfZOwvNGOsCC31Aa0u/tmwR2hmwwcTVOCpSDYR1gOXl5ex/Nh1Z3wrJYOQTDENe4
EioOka9uK34lVZxj5wddNNpYU7v08FPszvN9zxSAs2z01F1d/UWoJQB4IqgeyFf6
prnrHCSyAn3UC8cbHI1GLUbfw9ia9sebpygPRUBK591LoXnu67mOecPVNuEjd354
qW+Id/XSTq9vefAO5Kq86rgnXP1rxSLjboo+IfCHoyoaEaW/dIoR9GdEbNxX7597
6CZsF4FeJHcw4PBsydMuKVER+rwBgrPPhlQSTzSi/hBvFpw+WbXqDKNF76RcNT/T
QyHt8HFZN6ngY0EZzveMEynCwFPeJJvTFRWpWCsl2sCCJ83zS21z7hv1q+d4BdqP
2CWtgY4EwX9HFlN5iFDSHb3HaTnSkT65qcnkB3N5MZlL22z3QRfZmidBFeq1ynRU
SPInFGEqebw6LNrfEz2SrrvpNeNmatEoMv5Zo9WEVLuWjZCW2YYc3ETNgSiEZKlD
/0Q9arHeCFNHAxk5ADNUeW4laD1LLX6/RSksgxGNJs7v1IuDquIavcG2D3SVgVdL
2I/dvp1c4qIoDdEC049kINyK4NN27ffYqg3EhyEUy4P1AYt2EYiqPjUDyPGp641S
U5cIyYk99vG7HN3lRFh+EWDHHPgkhXuz/udrGEwn3RSaOuUGoe1tIJxGchlV56Q0
cP89DEIk3nOfGzgeFPAJj+RWDGRXwTt+Oootml3CvQElpSw546bbe2/00g0jt5gp
g5IhLX/mhEi6X2f9f/UkCL7ku1m5SuSxDj3vHvQI2FTrs4r04lz0Pg7lhflbyIim
s4SW9RrkoxjQFvSIPB51n68xK+Qu52U9N1UAQkcsl4oFPyijIMjSZOr/orvX/V2C
2OiSVB3CHw7eeXNyr08SzPm73IQjyi7uO+dx2oQPOWtLGTtKhgsjvBEe74pg64m4
Cb0TGknLpVX5B++qamprkuFPsKdprGxmsuLFGLaSwcwnXyqy5aMJF8jK+LnlDYSY
CZ2M+q2VahqbCspRwcQPifruYMc5CkcsUCfNaRguUnTyPpfrbgVByfwldgAza5XO
4gCW415Tz70W+JuZwDBIetyz8cbPpnLepa+Ra/aYrHenj7L9oXabpASR+lwbIH+U
uRR8AUFe40Oy4swLrT1FrWyDfAZjwl8xVd7vkInQNtNjEI4J/Z0rX+6VG8KPq7Dx
K4gPV7XOoH1nAIqyNbFvn0Jxl216d8boKzQSVxMtdwNGTjLabZX0xAQmAPMbrLVX
CXi94hYT1H9GtYJGnQjNpCLwFY8SvsKfDAJDcZg+Gk2NXyqTHRGF11oZKqij00ld
CAs+w4dyT8+QNjn5vbds4QnnFFHqwX9ex0PaiBjwSRF2oCGPTt86w7SBs1AixiqT
OLW9h6wBH2ixdufJUKTBCYEGBklgPVPc0fOIRLqp7JVkhIEiNW88Qrxt7r34AIFf
fsv6UVi4uMhdhVshwbrzzvyA5xPnsrHJxLee4AStHAeYMDvOMMFhpeBUyak6PN5s
wnxcxbTxEdJ5+zHtZHe6ZCqcQATkAIFn2ktEMMQs1y9+wV7P9Ufu9qptgmggErXY
rqS4J6r0zD4l5woLX6zsXocHieSX0IWnijbGqsMh47vb6MfWBubIl2hgLiwkAMrC
YE46fpkejZXDoNLG1Cl32lAZocP1HVAThek+A7zmseKiPpWdk82pqkR2QEg3YEr6
s2K6au0jMkvg9jIHwRTiNZBpm/WcFvUmw+M/3M00HeuDxr6wZvlfjIsAh4XQs5K7
5j0tZAR8xp+NJcXmAqw9ydThmSJBPO7qhtlBJpqvjZTBMGhcjM+vQvw3SFKyeRtf
GV0H07gxlRlTfiwGMi3+bZLQh4JXddp5QL+dReSq8Bd721J7+6kKp6DiJ+xabbkU
8zqS6SwosgWC+0LLo/j0leCEhTAxQXTuFtDUYNPoGdpOYz6YV4IxDlNTC96virVi
jNHH8Xe5wFojs/i4MMWsS3RsyyJEQmohEYVVGHlV8IHrsOpD8zjjqsZn1fkj7Qj5
i97Wwa43N0tq6q/7WqYIQQTtldYUQjWSkYjV2KiQzToz7y5UvOV0r/sx3dI8MzQF
aUKVUkB38GVp0qeAnxWeavHlHovTv6txnbXtCGC46760UBMwffaIGuE84721hObk
1/NMTL4KR1UaWgy3/cbVeI6N8N4dD7qhYcWAk4WXaFnfeqEzekTWFHAaLYp1S7qB
Y4ZcMQA2lxpBAjkOxlyH/+gHDDIl8FsdX7brDty0a411xv5qTE5fhDRFET9FbVBD
mex15jnY8nvXSSGy3Q7+O2NtV7kl0fDqMFoQ1lhRn6bsqOy9wvgmVZ+c+7q99phg
L7DiW0ABp6fR7jlJ5+NMkGYnTIyEWvIotc061MYf5sjdIbqMXHfMRUtebhAjNjDd
68DYcpe69gzU4LaSuA3NRZW6D3+Rxn5xP8GvakKI5LS42d+wwMSYWBVxiFczRk7J
PI3z72JOP40zOjo7A1p0xwug9At3pMlupS1anzmUFT+m0fRNr+DblaG+kfbv7kdC
360obj13GjadtIzFE6Zj4oA5F7N7xw1gp/1TBSWQ2ZlqhNkrEbLYAsjINduKFHaV
lFDvnjfGKb90c0aX57gJ5+Quz+9cNpJuW7KLZ4C/89n1T5VnR5SXJ2oIefhjxbZO
pYhGImg89mhqXvreBjEFzqLnsOm9TCsHo6t63rWCIalyHbLBbOPG6LKLadmXS59w
hkA2BaJ/T/RbY2+fI0gbHjbrjsaJh4xIwyutEqXDJFKYRVXP/vuduSJ+urYpYOnS
xYTHlD2Tzx9KkeoMuUJzyLerRUDi9UUKdvOuHqgJFxOYLTA45nhPYrCRLhL4JnaQ
UlOMrxiKXTVPeyaz5JczIAKFGFeG2XBaz7r9ru0G43ecQSZu1F4PDrvWPpCqceE9
z1TIz+s8FFU5Bzojer52x7sogoiLcXgEU/zID1wMPz+n9xwmwzliudtQYx7goXL5
tTBj88qU+fnXCZ3qfX7l+Ih760XfBmyxOdQp7EIFftV+RoIlf4Bd891g0SbvmMNw
qhdLbWDfa6p4cck2My1givigrI56Y/AP1UGxUMNhue0AbLAb5vQr4Qof0m2V/5HU
U+HX4VjOTPbaEpFAJ/MbZtH/3tlqOv8o8RO5V9q8J5HxWD5CsGX9+zCZBSs1L2s8
HC+/dCYufi2xFTwuWTczYJyp2h6FDe9bGLjkrBeDCOOwDqRVANjrTi4iNNTtwMfb
v0Va9RUd1zbXui+aDUa6z7wCunMsromrmMMxvbvBb6aFFk7ohyca9UaO4wjSgQPO
0+bhDvBaSk6+QiUnGrpCejtUJVtCYcv2XmL1gMD9Nqb8LEb5ggGLmYFwVMsn8cKG
R0YcaP31drvqbpI85pz75BnWy3RL2kx1R1NzRWvxtOdKOIdpaN0G8/icCoQjmmmH
ptcRBNSX8oY6T2NEBt3ATxgvck34Xv9OftjZWkptA5Qp5Fdf5oARrYEvwoBzQZTv
UyHjqEBZ33+YNkcoagvgkFLYl5vQCrr31Uv+heNuKZ2T1EdzbJSH7aU/B+QKDWQh
yc+GIy/uQTxBo/BZ+K0u8OjL9x1mDHaqSplAILFzx96HUhBHCNTAi8tAtVzN/Ftz
p7Obap5NZ+uqjCO6bpxBKbFk0ZagXKQ2WxcloYMsUtpzSjHvPCMOfFgcHcjKG5Dk
jXMjUKtrZMvngAme2/rDW01AKr+t29l1oOWj6plWhWLz7FMBmsc4jYGvEzurlpQh
ZwL3IcThvTWEqjgDHqrj10JxMjsJK1F/ySXnOyB2lCsWRZmih2bDJvLeSJ+CFuJ6
Ac3EpT/qG9zrFzTlHT7io4ifm6mrJ8xODrtWEfMaxfWq8QZw6HCtUNdRK4L2fC2X
FskT635w0WomngpKTMbTYLds2Mqlr7s/JljVZwWcRemYFIDqWFSQm62m+1Th3F2Y
1CblGBiUL/SYTxraPs26AZ/rslXSwgRXFWBm1QKLrPDku64y/ovV1zd+/9ZPhCY3
2OrGnE+/paElA2XXltKR29gy5qGCnlDILIwkXl5RbljLqFesf6DGVWWK5gbxJeQ2
mOMKXdQCkSoobbj+UB0KrrlkjkZmltBh6swVYKq/1htkjjuadfnSMijg3qb0FA/f
JSN7/7zU+nMMGOT6sBdoO+AZITv4Ma8Xph683dUlHyezdht88eLC/l571mk9b7hL
eJkpB9CVrEnrpgFohHvVF7lP65a2pZvjK5bFTV6eaumHYidK/dVs7k/cYBeVkib/
zxhBSzfFu2Vo9JlJsDGPTymuKdeNsfje8IiqMiKyuxJfI1lAdxf/D4ymUAMKmuiO
3E78a2WBUYnfH+73PJERLuI7qgLY/swtA8xBHpjTdSoLcP6oEC3o54AyASgOIuJM
a8BAwHVknZuHJSVA7k8idvGl3DnX+HiL4dCE/xCEEvOzEpFbziCZkur8+nrk5NAB
/v6wCv5Fl01P0JNZ1YaxG+oDC8qRaAPGVkqscRVXV04cF6FFVoXoRYAX63PkfY0L
W9C7OlDx4EFyixroCbN25GE1gqC56OMqGucKIdRVl7nUZg4W0KSCM2uhOcPTGtTm
xLPXGNMVXhX1IxDyZ53r3x87XF8AckzvVK5ISGatwJF9/PXDWHBuAeV5KJSVgCuk
iPVCM+WH2vjN1TlUxg4dYWljoaE/g8+4wV8alydieyU0i2y4STm4+z2inX55bGln
09ySLlry+wE3Ef1sIWFi7KbN4a6w5opuNmZkwlpYcp8fEKnLQAs9Ktoj6HOJhVhr
tuNxHQJjI6Ib2T7ZvxNLQ9m5a05lFGl4Xy86PdhZaxun0JVQ46S+kFJ0Lu3koRUn
+B2ivVG0adqf/PvPKmeZs2rcJMIepe3dVvVSIgDxf66fuzPw41kL0BsvcGRljSnl
XM+XSb+gQ60k9Fxf2eN2ewrWLQEQvidCsoQBQ6z1ybqxhIh7ZLD27VxTyZwo75Iw
0PIf8RNAqmvlo0mY5SSDRULiFckDUJlIsVpGmDyU3QPRXrDsgdojEVC4hW6lPjoJ
/OHw64k0LcZ8XN/E9sW255qo6lHDIIXx8FUBgDzDEJoHFVjzLf7nC8BfivUHZ+OU
GOFE6EeCOMj4B3JvefcHNlCegEMoWlxefTkJJVUwFDvSh47gPK2fAWKfZX8Dg5D7
GxjlL0wK+6UTvZZF1QcwhQdq7ldBpGD92PFzcW2oDmakxgPFp7qR4EWn/mz3eZjn
hRMNnEDttI+bkv20fjB6gUrKNFS/b2aqMq7EhVo7NLu25bJSUSnoB01U7rzI1z60
Rh0GpYD6IwA1YgnZKOJnXy6qzCkgFwbRM4fAh9pqcNdP9ZNhQSqJMLeu2T0CkKnU
kDSSgTT/rgC5npQbweQQ7KlB3i0Rp+1b93eoRBiRyVRCB6ZqxHIorvAb6jnL7D4R
R3lMR6/2hWrius7TpKqBGm4J9BAdU0O+pW3H7sNpHp3i687PTUKAWNc7W/+oRrG8
DNYgV2odMpwacVN+iH5OuXb/BTIfNsTKmwyIMMkAgsl8u8Z9zdkcynW9rKPuY0oA
pH5Ir1eeRYEqwq+zIJa9nBX89kk5ixiGWAOlFJM6IaAURmRBqfQuR5pPjq6g0R2d
7LpM8TAWuPLlkdLWAb21OmbFoVFpHTDk3rM5L1jhx/dWfvPXRfHe7Ti9EbM1CB7g
RBLmjhQPu8CQMdfK2b7aIZqf2qGlED7aVLRilCj02d/9MqKRHIT1GjAYHvDmV7w7
SqjTc+WXp6IS3MOzcckUVk72xOArVCgFMYD9G+5TuSBoOpPT1QhlS+zFxYzLRUAW
dAodi+vgNVKcLCshNQ26lp7eQiVtQORMA7h9Ys6NoIcc16UfE/utnLR2McwIIpFW
9RFMp6ZhbWfVDkDLGI9OKm29c4/DX/nV1s29hGXgbEOyp/msYM003qJ0OtIeSnIn
jgW9ScSlWXAhPSUf6fWt+4M3QywJHficWTJWCBtGDTV4HAXKM4tJCQajbuav54Uy
aLrQOm2o3D2qk6nUvFd2oOVfywsYS/PImU8U6kZmFkHig/JDaoj6+POng2kIkYX5
hFE3HK1gLSvf9JnXGljjIeqlz/ZKp5HbrkkQ/L4N64sriuAbsLT21bUlNzAL9oRZ
EvuoDBDO5HpvpOPAL482zgBeqYIo2v6Sc5kV0QCsGQrCLAJBNYRXlNk97hQd77u0
wzQHkWuPbwt5SRe1UrGp21rOAPSZtly+VGt1C7EqXRsJaTgub8qmXdhuZ+dCEyVy
OM47Qcwq0C6Szbl+O6r63GTo+slHxmXnrVk1aV2Iwyu4sMe+i/IiIwWa9DKtEfCT
mw0fu9B8yrMK9uR82JsW319/RAup1PUnsTWtP480Ukegdy7XdvecStyVCzE3LBpQ
vjzKY35q3a/+8rZqX+ZAlJTRoS5jMv3Fc3bSY7SRkZDOgjW9YK9hXWZJCtzbXsQM
AKHdk3iMtHRlp0wARSIf1+zOc5lRWwPJeSuhcpe0R80RFMk1e+D1fBbJufH0UINn
mteYmhvi9YFgYmV1Bn6aon00TIyzuBd1ziom0lrqoetCGXQtgLYNeCWgag0MJSLb
Nx6tT6n/QeDnkqdawgi1DZ6s8eBJi3a45n6srNy4MoqEipD/CfRTt0KqBcr/Vi6m
q8Q5Yy7e6g9F7zYpobV6wrmQL9yVm7MqlP8BU+/+wgjewKmvxuS22c8FbiotbL2x
zJ1f9YePxFJMnuzp91JAXfYSgOxuqsGSb0prC6Jxk5X58f6TYeBh77bBG1HXvkDz
r7TeNYQZbG4jToHqEcsyOOViLjbuGtXQpMm/nKdi/nBsxlbPArsI5bMQungLetdi
Ic9An2ZMX/9u4PI5hnbbYmp3ZbRNklFRvYSfJzfpMD7AdJe1AE4Y4DFe4aa54tj3
prNHFAhjqNxeznFtLDzmaRQc3PgYvS+uz7nvdQ0xnFZ9LqyTgexzq2mDLM9kFWY6
04icRZvXVvZ1VSBROlnj6l0/Cn52xTJof+Acf0zVMn5F4x6AQUzaCqLifxtURXPT
n3ho/T0+KF5J/GigTPdqV1Fy5kbP0gSjfJf6XCa636nwIkgOH7muRCGY0xeBRobk
LwQuFK/5y4U3HRwCau5ge7iSrGRKJDTsODS9U4oFrn8Q6l/pigDVqfBDhZsHlMrr
70C+HU2FSQboCAvM2hlbQkeRI09Q3ntituUvi8i+65lEvaVSroLGISFaG6mbxnur
k3L6vqOso1oHjLDbwmt4DhHVnVYzn9CdB5lCX3V+XjTXLfihIGrpUkIG1fEF6v7t
lXBql6m+UbuxkvN1RcK6twFxfdjDkDGo5fXzD2UMp0XHqcxHLknWYcSNSdsPIgR4
fItS0jRu4wk+TWIsiXBTGkeAXDIMsSFIBCyf1ZsUssxcuVvZz9cAWdBq55LcfGnF
+GLouFihPehpjIJu080/+0ayQvWKGBQKBma8mKPnBdxuNO4pXVZLS4DLmE3eVJ32
JUxlRVcZmTjjaAdXIgeqZR23F665Y4foUatHZYoI9m6khA99OuYt+N2Nb0QJQrfi
fvbSnbnjv0Ul5reOCBeAw1npZCAgmT6Cx9qcL2uJQ9dX6n+4oxnQn8Qs4pS7ghHo
MVpzci5HXXK+Gl+zeI6idYEB6oxL1ZX7oKm8dsCjz33nxc9hFk/xf3CTc0bZAFiE
0vRGSpjvUgMmN4XusFMYSoxdIwPUUtnU3z1wIzE3wevQtVsoTMHlno4NiNKKmoxP
L4mbfi3cOl5+raznRARypbCO1dVC8Dozw74hDiRG99y6QHtt5w0GMaN8CHLJ9Nbv
totQiY/ZzI9i8Xz7Cam1u85sFtKeSKoMLwZK0WxE/UUtlEvzjR0cjKoJr+qm8kGm
3fzoDDGcOPksV12RdqwhRSMkHFpeKXAMuVJMj91CGrCJovv9c3ZEetyiiE1dUaIc
uFehWrP2b8OZ2j0BqoWSkTWUibGmrPi7BskBIj+oo04K1VAugM8zO9TxqSAZIOve
i5FGqoy2Sqj+j7aUgdV/5V7ypN2NmRnLHmTjdtEwf4OlulpcItv0uRMI+Q+a6Mir
OWcOJ/GloCWyMVcscgnW7WpurfL6IvSa1iE/Hqoikx0ptXofMvPH8YbIKEga1DWA
a04xIUduJZuHtY0T7wpteo2VB0pXuk6YltxKv8QwmMSRbWqo9w9+G4NXultPAj/R
0RWMoAV9CdlSXH7qC5vSyLIM5XMJyoik/vgzOyfZkP0fQPFfyW+tb+A/GEwKWnYT
tCYUK3PMtwR4qvMm4WTaupup3w2yRTFsSvG7B+U8dp8ZFFjSCAVrU1pXmrCPgBos
YCSZ3N+rN3Yn71Rdk8y8wNy5VNvOBaMoE7WyqkOYqdXXlsyeR9l/9yE3kMd1D+oU
5gjXnsMTNddkzStn6CLz+dkbqV2KzWKL7bSgqf+oduLru15LC01HjRiZElzwWXNz
xDNUT8uzvIiNFLubbKEsOsxlh4UwV/YQqJsDlU70ABTFe6RYgyZLoZoX6o3sAR8W
VLOBuoC4cNLCOKip3J91xk3m0R/JrKspppEbo5deLHiDwGqQJAn4D5MRGAD4J8z7
4VwiSE4EE41pIgIr3lkZHRy2v3FsjScYJBnlYk/f4wq6W/LELtS4rudjXxzg/6J7
kl5h1gmwbixeFtnh09tFQDWomoelLXEVqRtTq6vLpT8A2EVG+QiiDnL0AI3gyTX8
p/gXtHq/POG8CElN8ydhjLBkgZlI6ZAqpZuxL+VwjcYDZWrY9Mys7n6nVpbJYXEF
q4x83Facxl5Pir1Is94POILlvh/aQh/zi5tGNxmBtPfT5QMCs6fEE33ham05M7xC
BqUb9rmn7bhP/y31V63ABZu6sZW4CVEtOLdE10j3uG1pViTq6rtZI4E9WSSuzBN1
Z7tMSDj3rGUZml695S37DL9tJv49okaIMtMW/VkPNpPogKdtFpWc6qTsRexdeHK0
dSSC9GbCntzfRft9f2sZR7fPPkcxhn9VW/C8Nru2ebn6DXxfxsa5ySO1TiantRzU
CL8CEFXFSUOxzL2lm16dwbUoQqKv2jkmiRzC3hBDZqKKdCSt1jfrmX5Tuh/j716a
5BzdeAxepwA2isTkxiuxlD/MwBp+qpN3EfaDZdHJ78ZOWdodi6RaHO9Y54AitycV
nm0iigRdg8HkBEm3mLQNdQEa07ccm7UgXzqWT3r4gOudSDoTYqHOEgVmP8BJ+mQP
MnFrKxncWlSTnbzI7jTDXEP7eD+hPmSrXbE7wGbiWYWX6Rm42/eaSmBf0x3DtBLd
by8c2NAywvcxwCvjWn4C2dZdEG9BowhPfmqXrgm1N1xQwZMQsDFo+XMqTuaX5gzh
zyE0W8Gu9AbykJcVUQwSlFKSXeIlj+8Ib6zyV/1L7AOvMpHmK39Pg41W+/hl9SMf
0tbNbJER+50iHXHWjCQlG5Wtz2lW+/RmN41nGY3HqvEru2eikIIBIz3HP6RgGnzN
bq3TzeELg7tSFrnSN6BKE2wRXsBhEU0I5qzZF8wnFoL3GlsTZpDIhxZiikdg75ZJ
Mwzga5/kGLwJa7fd1GHcU/wTjRuDvZVSb3T/4m04zhBaDSQeso4dKhkdRtn/OySa
MPO8UzYSsHqsctajvfuNnRYx8kbufsetOsGTcJhjN/jI0YsaTPw0C1vXXVUxUFRq
FTaAta1ISGQ4XJnmcJxXSaHC8/YPyNwzLplYoKMdRe0Ja8R9/pYUh5/LFoMija55
6j7C8V7z9fBLid/lOQoFLJlC3GJrRlUMa82V6JMBbY15axFTQWWqQeG+D6uk0NbB
wscxB7tn0r5Fbvd3tK6yghUUoTJe3KQItjOFXPo/CK+jPOeKW/V9Qy8iDfXy2ZDu
oPKo8D9Zld2OMVWcP/kxw1C3Q18UoONrXBIVWM1WEhncBOoPtlLoLv3LS2fV7Su/
vqcR6THnzx8T1F9oqBdvXwTDP++X51ZkAfnTlQDXZRPWr7/BhFLSItb4Qo2wpL8y
LN3Hg9ERjshxszMrubDJ3q7gAVzaF8bZbR43m1Njq9Xqa8m7N6uVFL9SbggUSyOl
X88DZtUf2SyOYp1hdXn8JZdNOSf+FiAaCBUMyTfTcL7ueLrZ8Y3T67mbXvXfKlka
iv02KvBE3hGio1GdruT9UbMQCmFNB/7KJN2ENSG2AHh63qIEcapzEZXp+ALCOjEk
u5lxHYnybhbac6Vz0cCxQuM6oA3kANt18bbSbmN9hKIvTZxLk2+UonxxqmzyS6yA
aSek/CYjSXlcwlXhXveiKR6iEQbQOX4j+po8acrtJIUTDVg4gGokyAd58hiu0l7B
Fe7qCTCEeWKULxKB3tBfjd1y56nG9So72fFsgzTX+8Mcy91FFNNTWHBYbnBSUgMu
UXZIA1Yq+wN9xjt0ydzfqcmGP+N1fP/FOEkyTxeNO0D7lv9XR1S60lor7iiK40wR
eNMkidZ+O4Hxs4USMXv3Lg6/bEXBgrXm/MPqal5b86HCxVLa4RYYTSRClm54jw0u
JUmRRvkutAT89tappD+2dpnNTUQ9lRNDDCFUtsx0msXGTrBTPh/XmJ/6DTo2bCxf
yvfvy46iIng7Zu8Q1GUTNni107MnqV2Wl5OUvVfVlF7lNXNdaffD1QXhtsR6gArJ
rzXLEKN75Y7929+wavHtlsNFyHpobxGk3kWzuGrXvk7c0uqI+fYNgV180j2ERGuJ
fdg3qm7sRrgULF1eV/jFIdfGj5Gfz6MLF/4B2kbsV0R9VoGFIPY5GBtYsjzml2G5
po3CSyjLZiwmG8llGX6Zefzc/ti6s/t267NCtgyBwbArcKvFaTcdGRmGvKsoagH/
1pb8UwMUtILQyCFh/HDu+80Vn8OgN8gk4ddEc/Gek8thmZTWUSoMTWARBPXt1leb
+DbAr7BfcV0os2Hj5MpTzHV7s6k8ShqVWs/2IS6iHb9fZ6yIJcCKPvcNmuMIdwN8
wutH6SbBKpqtQWIzSONJ129n8mVUyfeOyXAUCbC2tgbO/HRiUWyxqAeBWwUR310k
ZGEFF8ENOD/DSh8Hq4zvTCqRfLVjIN+CnkMnwOoi0EcpxQhbM237g3I+LgaPInkW
lPjLDd2TYOGzLc9ThKwZiVXzODB4G0YNJHT61ASDkmI5QphPTzFo4cN8dJUVfPBr
XFZyOaydXsdXzLSAPl0mTqQdsQy5VWSgT6lUjAH4+Cld+XjkCzUZ3KaZWTZbWTXO
PkcP4jfMrPjM3fcKYdXNIDPBM81rcDF9tD6jhIY8w1KCNJ1OIQW/O/ZdDdIC1G9w
neddl0CSDJkVjGOrn6aqrUEAYvv6sTIC1cPiEj/skMLbtVOPY+ttqyZyaJV2//6K
Mkuxu3viWoFhV9C0RKyzwgfIQ7Eo+tG9PdAzD+YJt0AiMOn9X5WXmKdTXsbAiqFL
w3wrJO2c8LhE4kmNL21JdW54NrsYe9sRgZ7eZvjPIfDZzK5sm8itFClPyGoUTwtx
5z/8wAbzUov1nkbh3YYBYXH40VkNfqylxEGRnStkUR7qW9flWZNlwR9sC/0k+/Bu
jv0CKfIAZTeXGqaboWaQ62QrwE7kJQ3g2oZ5yY/jgkrabW0F7PLVlMyPJjcGiyP0
h71XK8Oak3c2ivb7hrm5GjnEZkgEM3yviJwtDXWR7WQh2K5G64TIYieg9PKu1Uq0
tyeMzzi07Z3bRnarZweO8xd3IB3POnx3s+21vUMfA/BtO1mnXUQlWXOesAu6f7my
5aAI75XPQtlGXUfDMjo992LfTPtACE0rp36g4vC1cW6k1dMuPlmyukJcjgH8Y0+F
NAs3tthpmE20njC/WL7BK+IW/BJwzpa0/dHk9bytCJy53EwVZ0+vOwIgrQpHTUhz
cw0PrVn9PwMAFvklO9dAN/xGfWvviNCQCh927tEL2k7DuMatI3jd2GBgmmxFVvL2
ePTdSVG+i+OEV+tlkj6sPiAUIEDn3r1G2VRqmcqzu1SqNJWcAA5Vaur8IkoAmhjI
ehiPG4II9PqRiv91ZhKgHR3ufUVsCSqR9hDtUlBnHFsh//bSh2cKpvsepHMFRscb
IWvkiH6x+lI7AKwRl3hZtDEXubWETK6n5Fb55MnWqOc5CqBvv9PKz8YdSPd90+Ku
H1pRCFSonCptjXdh+7gMAaLLSU+uy/ugtnNPNTZZh1zhedLtlFdqYe0LewNnWJSN
HZgcQUzoHjGPK5kE+OxTb5uCKYjTU5imF+ldAvFkBqedZuhkw6L7g7lbly3ipd7t
vgP3ZDTesPLIj1ImByVgRNbg+t5/68GGWZtF7r9yF8tx2XueB5ZiuBReD9qRShOu
/cfEG2X1s9hnZL5D4W5jdd1ht7A+a2xzcVXu02SUac5Lq3bW0wxylfrgXVjtyx9R
0wTvgNUofuyTdkgw2rcaXOHXgaBPpHSYMfgmtInRUnDf3wh8ssSh1e8QRxVfo92y
+WsAj5Ft8WEsLdHohRv1FiyjzjqN1oX85pjzSQFtkJnha6p4nANMCqTYr6djngcq
KeN2fShPQS/iZvvq1US3E+VXBgFWLpPCOHihC71q2ijwn42E7Y01CSGYDDaiGmYZ
cKKzl0xgI7vedO9LkRAj58twjbqIaGEIEFY+FpSwwUBQJVMX2S5N2q35J9FpCpxB
m7GfzFJohGw/OT9PUXiTV32JFJMZHKL9hopV8mEkABJTsaA5AkOtIfRy4zB7oqNz
O9ZzWXfmah/xj3Z54m5I2F6KjBsmhmGdRf15QYeHVTXalVGV4kGKVh/72pryP1ug
iONC6j8VThP+CDlbgQ2dkWohxgew26P8RyiEvMrHlk4H1++OozgvSC6t5koLi6xN
SJ86jkfIeFBZlIXdasud3pEpEhXKh1MgKYACptpIvCHl1eYDygszWz9MVtNbn7Q5
GTMUZBUaFrrkAjLX18bG2+54C+/Z9plTk7fs7rJIJtSeiMm2IhXgWGMf3b6tXzGG
vKEEU8twfb94Nni/dG+ceWcG+hHB31n8rXFbhe8iLEObvffPuBaIhnkG5tDjDRMU
G4dIIhqf4GayaxGLznUsy0TpccA49YtAyXPM75ZZKqpJJPyc5EQs7FXFSCMR1DQ6
WuK3YnJIhTyNgMOsNMB/h2bGa/ED669KiOXEQmYbNhEqCle6eAcaoxJGHT9yNY1/
FME1OshF6B6wi6JCcsLlvWAtw0/i6NN0yNIkze7ra7xqMJzsBaZu726pV1a3G6XB
9Srzu8o5cgSoFQuwFdE0sKgtPqotdCLpH61X+Z7R3BGoje8TUcdhtkieiIIVU/gn
WHLnWjOQQISRIYwTV/4MJWBZWkqBBn3vCdoe9i9PbJOvPevMlYTrgZb8P6KKGjrf
JXPQImB4FnuXMw9WIJGVCj6XwPUYqQ09MsRmHO7Nzoq0RdCthX41EJF6ihRZGyyh
nvKHEM+tuTArwxc1dL5+UGpOGOKvEIG3gGUDiSrqD7wnSsi4DDrhPPmuWkRZX+cA
s1WQXbEjKGR15psXMYQL1OHofk4DuiFWo+Ws4WG1UTX0/xf6vZM4CfBFoh7NhFHX
j1Gbf+cyGCORL1Oy+3/sdg8ZyWvrajbw1M2rKl6uma1mUHzfs3sVVdMnosxvr6qP
HRCYrLT5PRMAFCFVdqPr8DIJ8aB93a6vuAPPi93da+n0l+3JzNuB4XOSs2Juj/Qw
+0yQsvDMwkCapjbAAFXkwBjSz9a1Js0kPWpW3NrsHeYzSx+a7AjEydE1xYasWCW3
y0kE2Et+iFQ3nSKjubsiHar19b4tcCvjcNl35UaKEz7eNPJPFPr4uxF3bm4mD25U
ggqqmkpNwMuXqnODQXLQYp/TKO7nSctbiq4vfPm8/ukkvTWIK2cflfV4glWXureC
/VYM94FbS6cY7hriyGkSBcE6WPzgbMLJnMGQ2G0RStzlZpp+GZg6CzjYjyNEvEbu
mOAKjJQSlSAZCeASYrjaogUfqGIy2PkiRW6ArS8stC+SkuPEj2NSCtTkdlF9LUO8
nmBeU8ujopMP+tlYQrRXjSv3C/P6w5f5ejRMaeJpzecRIpWuvsRYaVCI+2O7OscW
rfLxss6KZWNtIwOyDvrkZzrIAMihuKMHUuvyaJDIvBnczPE++DkOaBsSac416uD1
NJGgEWoI8Dc9IJIIRGt7Xl5TEkJE2F2BRFfZAhQzZrztoRApovUVsZ24ozIM5jID
qGSuETilsut+xCxBt8upH3U818kzYN8NWqMt3K0H03HEERb+rb2Mla7BVGtNZ07P
gD2CZAuGjE9mHzTvSFQ58/DBZ3T9WftKzBQjfFhfq+I9fIxHYjMm812vSDCHBpO4
SYq9L2WD56hq/xqaimtPoCna+ML0xIztR186jaVVIXujzkFZ8UwM1/dmFQYnfCWE
aBPAow9CKLRNqp8PybjMrwfk7XZnu0Qs8EewkuZhfUY6vznML/bV7pDra2Tkh2dx
6D1nEEt+KQ/CghNffzQ1AbhbkTeqDRGP3EI6WvswM6ORaDBgEwOI3jFpXV3jn4A8
lI5D/l6fbkDoVwtix5FMXVc7BZdm6RMY9yOtx8rtToOtOOaUoxUA7Erwh8GUE4j3
I8pJ9DKTHP8KuPxxoBHg2vSshFKkelmMj683ZY8nJmE8FUoEMQxDTIV+iX5kuyuB
6UFFgUodTnqbQxDpvSmDxFyd4Sw6H/Gcbn4b3ed8ti6pWd0tqsg/gpGHDOpPqExC
mKvxFf9a7FfYMvCqMqqDU1fLt3Y/qMDWR0wOCRrT4sAbcPKogXSRmnJAFimzmDY3
bgtFeuzsOlre+RIPNhBh7Alz5y1iDJDpQI9t8celSWVp+ibSMODKvK4H9Uf1opE+
wlUOlfiZ5cTfnfzItAkIejzqT7JZhb1cRNV3fqh2bu4Of43DDnqYKZx6ANjvYuB7
lY0LkIhIvQ5zf3rKQ5M4Tq/xmuph7F1ExaXqcqi1R7c6gSBNLar1iwYCGAJAGLnp
QrqBKrDoKTugPCbpxDbZJTFUTpeuIFg1kNls4jwOPjpvCN06w43UyxVVhvjqxjw9
UI6cNpYoCABs/KgXBdORFzs4STDBYmp8oUtCSegVmxtVQBJXFxy3x0cwqNvBfp63
u2vlKuCfL5+Rh88PJewim9PbsqdMgxOmLWp/mp0l0ZEP3ZinFWs3wpwVEtmNF0zE
vQdkNbmMWgtuU+HXSqBwbRgI+EcGc+NeQcStMO1HjFW2ZlAb8FXGVNHGA6E+cpCM
FKXnA4/f2+8G2iRtRqmbgt3S94rmTwzkjblMP3JlsrETuNECU5TPwmj1RcRtUJWa
9i56k8igMVFrmhmmeSnESlFbWbUoo8LmMAjb9wxRZhCBQhhuIZ9JCsOdP8YW1NNU
9gu/5F0inkcO8C8cWTA3+XPtUsDn3NdcaFCUUJG288OLhQ70XtVZ6opIkI+VrKP7
zu0JmnpSE/reeSFXZRAYThhinE9sOJpH5rb/c115LpbVXpw1U701zX+IdSzti+F+
++BAe4SyrnWznCnSZQ+FjDJcv68sH0XEQMd8tiNhXV+GI3X9SxQ6ZnvPSQqtuMhM
12V7ct/B11JFsxkVeoaC4j0ZyS3C9OwFfflXVJAvqlIgN0H8wUsPsgp3S0nbiniV
5L0Sfb80igM2SRjp4jXE9FNGWLdNGQhdlALpSE3M7LhNxQkaIyvj5G98QXlU6GbP
BPuF1KFVAxmOKGvnP8DYi9mIVlx8ZspF0x4nPDjDrZEs0nw+3fVslUDky3VJujAH
9IbbjBCnloCrv3i+bfkIcBMNjwHwPuUnFX8M4RRM4ZDprrMmZE/EfR8L7junLHJK
taEypNNk/H744VS2KuezkIFtXVc3QcQajaY6dZXuymvKT5/1mZJjN/kt4Ngmd6uf
+b0rrEzj/AWML9MIYRqCKWdtwTjwfQz17MJIqMErmN0nYWWfVyKZvQDE/DZCOJlS
4sOmyWUDlHgeui467TzrEaEGzLPSR/xE+rDmpZ/QK521Aj7JBk5VR8/WVYPiUhMb
hN2XVGjmcy9Uhj5LLcdymrvAmAfczrQrW8p/T+XqfONQ/amuYLiJYJRH3gVd/G9I
BoVlB2YN2M9o++1TcolXMzcaGEmruOUPNLr53PMaqeXvKsI3HtdPjpT6fkVepA1g
FQN8zxa34GCOwrXLTQBc8zDIzUqEvbueB/UFQKkR0YfIRQ1ZD4GS21sLg9Be49j5
KV7g6m40Zqa0+NHNnDD/FgQPNE17cTJ+xmeLqD2zQ6lFuUWcsJCsmdhOkKKuqozc
v+hTLB/kAB66tkTe4NjHpLQU0tYdxZv2WKiNoovqA18vMj5juvt1v3Hn9zGZKXvy
5P+nXIGmLu4rSDVE91ZJfg8m/ui4JRdhXKzFy0nTFXItdJT4EKyrpQjQczodevgK
oXv3ZnUpkv34G7cbpJlsEZZNDKdRj2ZDSab4pXVszdklQK40T6Nn8Lb8tOqaB6nE
5ZJ1KErftbCJXYQBsGkeFMBsoBNXAYtqp91rFd7nQAIgI3T7YBPkSQQbqqesWjUq
VV9nXv8MBQfv1+uyOATv9nO3tEstr9a8yD/qlmMVNapZaovtfH5PEqsLltXKmdDg
m81mFsx7V+Z80K1FSmgbC5bkoyYn83OpRLtoJ0wawy+zGS8KuFVuQte2Z8hlcF8+
Fa+gre/9QRPMz+hveXsHgCnPQqX+YgRgBZ2mmOcgKnpAkiBaEsFOxmJItzTih2E1
lKzGoJjVSYrvBy0cT5C2he72jJN/agVwobn3HQSKaYZ1yFI4/10ygysLg7YkqQmV
GCH3rIwHzMYWTWAa+t2Yj+/AveoZb7G4ZXkXRnzC3Ujb+GZCbZ9a8bUSRWCDvayQ
K5bWDrToYwfz7Kf8f3GqbRJPAGEez4+TtL9rQRE4eOMu0T8lNk74te2hKGOv4a+M
vqyKQExCVsL/fg2SYaIMl72NNGrMNRFnYiRr2iPf0ukXDL6P3+tht8BPE0eLLjeO
2fuMtceCk9J54LSMFD6lPHjnh4unUzVthLv8Jld/Ffb/WXA4bq0v1hduwA5L8hEW
oSYvkSh36nrpzmJOJ6AGE8qssjFPqUBASlMVMKrMEC94QXjue+Uen4SX+NkFI/gX
4K2hKmyyqCs0hRgFCbUbQK76JCeDaiLj3VIUQQYTnHpca2+CiEcQwgoI4xD8nqwO
q2CmlFoZRv/lR3vNECankjMqIutSAtFxNdtzRTNjhJf0XOxFg5YPn+wtGpcczE0v
ANGPvv2xKx3qdvYlvwc9a1JnyFE24WqJupRM/Kagp60/Wpf7K0Lfp4d00jk4JOR2
ftoRhYinJQs8AFktV5fnLMzi5qLzROjGwxvBvkGS0ztGWTJ/RaOaN2yw2W71amys
18ACwuGhyGuca/QajRA+WHSeBz2nh4rrvZR5li8ZT0K3TH66aoUrym3Li9Inm1Tw
746fUc7khGtbHp7xBM0EVk2y+Dli5AVx+iB5BOX77zTDn/wLiKRORPGUsbyRiqVi
s40x/AYYjC704PJeGPQhsmb1DpIu1Y58feNy4xdeNrFkK1KuZd4/j+Wfcl6uxQG1
k7iK68Z/36lDxmtP/1mD+9hnxpKSsxoZTigrbW/4yNCBwQDdwfHokstsZlX3bDyq
OD4JZy1paLTFvVMIp+/regcq7zhEtm8bP5vnoRwdHGjWFyujgoJ9ZJK6CtcbP0f8
NchN5Ai2KCEWg/WPnTXHyKLohaqp0VY+Qzh8y/w2AaQOHxaLmfkDl3grckUEXB9/
FvHGRw2EscbHVDtT6h7lWXX+KWMAqxXO70IoMD0HC6pbcjhk1ui78CwTmbWi7dy5
MH/47e4b6IPdn7L8ZP14XCTSb4nIiOyWx5hVKx+cVQ6yTzZP40vIhQF053b5yUbV
axXbAvpANgYNXE/4cVcR6cyP5qdAkfRHYwJ2RjmW97YoGmpUOfWNH0v5ScFD4Lil
R/A+moXnrLywPFcNKNd02UDTfAYs5gj5yqRCaG4S2Z1D7GXcn9xioKGY0wOS29cU
qPJrS+O/JMYAxxBkMF3hOxdJsiC9GQWRqFWSoW1WaNIWV3Q0j8HXmTGHWXxhyKcl
mFhWo6wMSRhstT61inWHtFq2nQeYs2rODOTvQ1870icS9w2ZWjkKDuIHmMnjD1+d
3owOhhcMF2OdVZErtpAcNoESwnpH1ceh5iIVQHfiEeOXlfVtvbXmeckdu5zAA2s2
d4fTa4hBlCZKS8OXEFAa8vsKyVvBsDuVBwN0+vfY9BdP2G6lYpW99LQZRZa6os1h
xWBZ+Gi9ajnaHhz5XOtD1YInDzoKQ0GRBO5pwaYmsfkyAr/WyU6WmAXRcQCTof7I
+0cPFfeoWLNfcvJL6U2GDmdfaBjW8NKU93ZmPtJBHMXEe6y57nwFZ8882PIpR20g
82o+u2T8S3eAru2itWy3cBj/ujDSuWrbfCk0Es5ERZUpimCTO+m98LXUoWWt8Pxu
6wU/ERQU/G2KRFWBxTUUaLpx06K+zfMYJxzRjc5fw9jhw2taBH85fH3VbzJqBBhu
bH/xYSYkv1S/AmQn+r8h6nIuE/ObS9tM9C0Rx17akteksajPzglEqtCDhmlQV5YX
VffZaGvZOd1NIo/VJXQfP27D84OvJlha6WF2YMs2QAPxTBdSKB6T8e0Xshvd5r6l
XfyBVRpn0xfXJKvlBY9bdzT+HR3s16BuAX7jAaSicghCi/3DKNWSdeHRXypIPUhA
JyRblpek5yYYdmM4rMb22nXLjAGlG27SeQRmZ4yh5DlwuYsxFLeGRmhudzDrV+Di
UhRnhjwfZTvjKTXFlGhAOkdEFUp+KNbinRQdexTT/C75xZhPFV4yzlzyebj/lzXY
w25wfc/hKeGi4nRb57v46OrCOjR8FzTrrNf0556WgcGFZoUzT2NvyWweyZDoLxc9
eXkpe/q+k5TIJR6ORAz8jUf0z2F/KRjIT7YizFytLSmDLPvoymAwKjPIUym9Iuue
l9XQooUyG+9AFZMBnFISzlU1+k9L1gMQMNX3pe+WggWRyib2hdxaBsLw1U29PDHt
0NnZ8jZEyoUQ3MtArrF0B/2qJRDm2AmF1q/ALE01XFTJ1looAuqU5H7LyAxyG+fm
a2y44BwZFrF+iOcoVIsJUragD3DTIWjh1R0+FoSUpyIRxkv063hozboeTLDNVYf5
56I4CQ8ACoucytGI/LP06O0fYkWU1frHS9qz1Mk39LHa24RxG4EhWs48B8gCdAGQ
aX3/fQ0wJndMeOfOau8UDKE8BdHGSnQ6th6XnAPYo8jlOzftfMqPauZspG2vjA31
BzXYYPO+8bpWeiU7HYTLAXyfj91eHgJK9cpXMpobSI/yzPkr3sAB8gTLpo/MGXH0
z43B7MYCCO1pZVOV3AXt/+3AnhgLM/FY2CZLJTYwxGz/DTUQZYvuqHZLQKVks8h1
x3ScCPdIRzU6Cf/4t7bxU9wHKRVOZAp5ovbIe0D+HlCyKNYXf++dgPqwtkLMO5s8
ipZhFdeQLAAazgjADPRxi9q+ONIgB64pLKpBeo1Gmj/oGPme0xj07+xcFpSqGb+h
rPQxejqg5tmCk3JAtnSLG/qbvM9RBAc+Ihycr76i7uktJ1ejowhsgpRQA8zSk980
TXryTOyva1n7pgg3frL65nyPcaqtZLgG0aHvD5tK4PDCw5kz+uKWTApwK212kdt/
UnQTsM/sA8aBav4hwYz5qG34BbMQLFKrkox8Nc3bIoAd1leHBYLfwti7QL2STsqG
vfPIddpokVn4/radRu0tS5/3q2+bPkkGtRNCEpliZBRUVadJkWG4ehvrxC9ElTYl
8BDdbohotFBCtKhEMD4oT3XvSl0JDGymhWhKApEtvnVzHeiyelEvOwotB1dLTJ4f
zBm2j/5z5cOpX6rfIFlO9lRDN4/MV/JaqOXaFPWmIEC+4C50LeZiTYK4bGpAZ8pB
qltnvkyjrwqdeLFGK+YVGMbg5iGv/goULu0yeVmr9HvDfjGs/HW6jhd7ZZw0zen5
OQhenjNW/x3TTxCn7dXiDwUafjj/1fIrZwSApJGaCdFZV4+F48Cczz9BNuk9VXfN
J1dfwHZqYCY4nQDOrhZa3+lACg51Z2aVLyx6vvgXGz4CgyE5uoG+4Ryq8GRZtVDk
JHaPcTIk5ljbVm6NAEo08/EdmxLCUPg+zGA76M1su22qQEcqXIr9rVj4/7mLGBfW
R4rGRHYQSEM0OmJT8x2VuWMGU9MXBqA1MvvEaXkpbbQmrQeJRTIftJQF8q6A6DdI
vIX4BCnAuxNrpnrF9PvmMiQSpPc4PBXYcgFkJvxse9W4h9mz/oBHDNxQOtopNSzb
qQAf9+TnedLfhtDQlEE95W4KN8t0YZS4c1pXFt6LQjmNd1DUOPiue00YKtxJUcTt
ZoFKvCXTDTEfPuxPdF4V1P2KuyHSu4peAT0mMK3ucf/HV693o9dCMVhiL1MXxe9p
d7mx/vxSSf9bP3Dwbl0nc5nSLXEiK2mUjuPqLsYchHhkcLh4fZQqFKEhQP+uHExZ
hq9nDpswzkiiDB7XcUulWwI+PDHVacrMnEdWVYcNkKYb0wbJhxzlZQF0mASKOE9X
avEXXHHUn0Gu3YH2eKgmVxxqGMi0o0Fc4Uq4Gm9qWKECbYIrKWNzzJZen6zEBUIn
vmyKzQbHMEq87shzWBGbhiKWPASHvW2676jhGuK9pH/pybvKmo0AVjeZ+9RaY5/C
CvcEqYGVKTS8bhSsJ7Zh5Ubn0LgD0y/Efh2mmOJE/0xd6LMcFHWqN08/MVbYoU+z
qDApxM5a+iMFepEdC/P/F+KdjDpZ7Hd0YARlYcYmLRrs2RwNnIMKD5SLpP8nfX47
8Y0uPEyEcJ9CLBvlJ+NKIWvxJAJuR8WHEAQFofMv4szUAmlGYylTFJH2Nb6RI7Et
x2UG9bQOizDTpOvyeYiqPROmZJOVXQwFEKK3t7c9e35WZKkLSIIWryRXH/ykztPD
MDHsaRuWcdizmQvEpqh9A/tO/KBh0C45vTm1R+wPzhCiJETsT3CmZLiWGvso4R7H
/VtahZNaRjYubHSD14UVnxJ3FDfgbL5RcWaES4RftEyQqZx9lP4/KZxQ2Ezvc5bJ
Ae5UklPcLvzlEZ0aJv5IwmBEzTyl0oH8nKkOmGO8+kG/SwwtK2HRc68lshN64U9m
vm9cFzjcLlEFlc7Y6Sp+giD/K1r/xxgqsEhMrg+ImzwDUla8ylKFd1AlEvnDTipD
Kn3X2a6LnLnlACkYwcQ8RbwV5X5A7iSZgfbdQyoVjGz0Zaoh92yglLlLwG4OI0VW
dr9KV1tJEkb1liUey03ee68ITmaJVAoIj2rdTyyshYnKx6Hc3C7Mg70U08VVyQNZ
srBfvLkHCcTpfXd9ZSiuSLk8b1JozZwDIZfwj2oNFbDcE+Hp/EQjEa/qfdZBiD/n
7KNLYGTER1zhrf0mbDwwkgneAM53hfoPDLXdLd3XglF7zR4ydLbpdEsE4wjYVIQv
QJvYhG65DMXKDafPe0+aUPHR6O/n2jE58kTB8UxqSMBvWrwc/DcMwh3ci0Fgimq1
yx8QuJToL/LFN5E3hWwUdOXy03wjg5X3XIj7AIoqi28MYdKp7fXxBmJvw0gAG4Wg
BeBczcobTDOndRjjqroMJKOKLKpy1GOwNC7CNpfYqTKXIOX4bpXoo+rEKke7Zw+r
BhIVubSETcKz93RjYHKzOsGy9c+sIsKi0tkqOs+z0t0VQ+1p+wxISMpCGnPORMPR
FExi28npEWBsHlvTqw6V9MaknD6BqFdG2cLQEOnHxLtt85NMR1cC+E2Vj/9rGL7g
JhLc/cyNEwTBzhDh9pxbIin/nzD8OgIKhc9xv3Jg45fTdfqWCrtvD9ChoGWEuRoh
ZPN7E9Hhmqjrys/qJxum+fNWIUjAhxQQRL8BL/r12fzHjDhhRAi9a1WlQ598cz5s
2M/wQJwwi3fZzogDn6XfXMt9eZpmIHKcy6nHbov0vs1BohPILjeqfWv8D24KYTlk
AnHimptTznha/joFU5LrI9d4dt9JwMFpAQDWqctWkA5GPClJgqD03YE2vMIVppEK
WLgUXN26oZK0peQDNYQiSXLTwnos6OUaswb9h+lHlxkVIVnKygPSzKydSp94UC/C
eIKPkLCuiBeTruOY6I0393s8qVjZ68iSk7sDaM4He15DRtLn/dcqHqK7zQBA3vqO
IOewWY4SHZpJT8wwCA0Wdy6kBPBf0zw2VK4Iq1Xtr5jb9+0cY6tjVUiU1nqCxO/9
WzOdGt+AzG2AI1fmFapVBgCadG05imZ2nRoJ7pB57PNIS0MAYpDZauEfh30jcqsS
nYIQkruOABKTbTnhY54U7X54Vdbyix705loNDBhbXDDUt6KpC7OSCQLUrsSI2QTY
6h/qSrIBAmh5xO4tVdH4MLUi2sk2q/i2UVKM2TSqoacaSPLTJCIvidQV+uEh2Agt
eab5I0QjUjYVRn6U6oeYRunjXq1iIV7Gt6er9aFXOx99vJ+d53KmLabV8z6ilIc+
Q3IpmRtU2MOZnLy6AiMyIfxkTMbDhJXAa8qvgdO74F4t+5fJ9rNf94uJlJLudEdk
KQNl+UGoU3nxn5sa344p/i7bkz7rOzMjlHHlHsss/MOCXNLjljLUG58mwTpw9vFz
Xis6PIscGy+756SBa2ASU29NPZVHYLHoiOftaeQJHAMlEOgdBhAfaSzYfrrBy4vk
uLyejaK4Jjc4i4nnu38cGijSVQoKR0HA/4fA8dvgGb+GxQ+WL0lkz9437fsblShH
C+FiJvfH64+eWGrtBIIxh1Zv7S/Mdmdau0+9BetZv/evU/X7QV6Z3RBsIBQoEjiG
M6f4rX4UuVljIB+sTco3eiohdOoTfpr9Y2lTN7j77bTNZvtWQqQeieIOXqQvr4e8
y1oh8GXG0pBzD1zMPRrvs6TS+tlZ+pAr/fpsLl4SyDr/Yjs7mYQS0CmseANvoctR
WZNPuC3jXOc+Dd+jx1MUO5DoKOvrcOZdidPOHY8pj/EYcCtopcMUKMtUzq+Se117
RusHmiLk1/TcH2vktmrMdY5sovl8qLg0TiDF09qsa46UX4Sj1d62jytn/ez4jQTW
fHHjqY3Obrz07MLTEUN3olxn5hUYMwo+yqEzt4a6nEGpC/lmPFaFo2FVbfc/Dq1v
LvOewpw8U3vqHmzIxD5mbVTFW04yYeuVUedPtkkR/L+gKx03nfCmrWSXhDrsS093
c7Qf465ksnRe/H5A546kTIxQAoexvZ7CwE4dmh1X0gEXAyoB9yeQkJHRabLr6lgu
K5wBdFC58KtzmIPFOtKmIXBQViBSX9Molf9oDCpFEMYweeYcKHyFNZRj/k2x/Hin
OQGPMuR1f0tr7AA5vMg5tHfd0BvRwsm3eK7eSZNAeyNIc4cb3pl1g3N+UVqS8wSY
RVQ1jHGFWiSGgNa0n1Ml4Aq9QukmEG/2LAm8nDSjuFxAVgODZ1mbu7oIeKsD2l8Y
ZGSmutqJbPwNxOincPH9C3y4EJezAGzURYT5/GPW17ppwnpk60285LQqHH685KnM
OfASvAoY/9thE2dc9z2BxVmD5Fpzsg1m+9792z4Hq5RfkExKguRKr3MtzYtyVeoW
iFPVGTQzSilcHuIZh4oUw3MCcmeGV2vEQ/kGvvcRMb1y7TiGBwne3ivKLH5+S+O6
2tIzYtSFec0fqm9QJVhvxOyKrkfIQEX/zVBedg0geXJlVJpSNs+bEK9U1RNOc0Db
Rreo+9+oIoYmJZWR78Ql4xhHooPLm7uI0urHU1ljkoW48gAdc1H4qPjE/6uzoear
mb9jX/Sqzcwl4o1EPfR6hPRUjm3/QuLJ1Hvs1XjgHrY1hhmNGBF/lBYoSj3kzRc/
0d/khn3X1cMuj5p+67E/MHT+PLAJg8kUjahJwKZHNHQmQooIYOOq3wc2/fl2I4UO
uYe4V5p3mBvobPpLyFHpsFpTNmyuSQohAyCXalm3JGJYsQgjbk+o10kIF4V7rUfA
7lB2zfdfanoWnOdK5WX7artB8GaGhExuMVlnyLf4uwUoADmSqINTn7uzKOsbVZ2M
YoydQkI1frUzVzyicNCQLcnyNXfyz4UUmZwUGllo0N7Vpw6Hwe9W+GbWObYoT/va
oxhg7uRMVTpk6tJILiI5RTvfGcZig0ZAA6eL8tnuGwVbzC15ETfvW+HH4WvWAyUH
+v7SDWWCxEQT95ss6hoAU0epxTWuNOk629LXsqOmnskyqb058hTkHt/RvNaoRgop
MzsvKhUg0WpByZAP3ynoqGTcrqDHtBIuZfanqxdsvlOlmLYyObpyfI/8JTcKxDax
+JwgHVcg38fLpBdfaKhc5rxEdmgRMRRvH5koIF9bDGyJyWGLDrEJJh0PUN6qQqad
PknbAqVxPUbIOtB4pfL/8hJfoOkB9kOtR1D4f5UqgWFrO8KF7AnyZoQeMwUpndgu
RmuytTfKeuwS4Cjj0YfZ2h1PxwAQxU9ZHJ00wKnXVseaDgortqOo75HssLv58zfX
6xJTNQ7ws2CP8mpuBp8+Mv+RsvIp78BL80dP4U4OmpDQl5uYKskpt/gWPfHAKW3l
q+eloeHjfClJLEHKw51uUsGVa8Y+5EVuJMxesXSzDKR+t/i7yC7kNuf7s/0c3EU1
GICQlNfZ6zkGomKexM6MP4EgpAICNSVtqTmO2xdXLEKUtrTCtGkzHKv2ql6Xf1oF
C6loolYD5Wn5bG55XXkUmUJqf+jKvpyn0HEdLm/vx6OTAenBl5RTr7Y6VC5INgop
QEuZ6unFTDYLfa9L48rwKmK8thQWTVFh1Cg1YHO9n2unsdpHKYU25sVxLOsYcX0l
Mr04pzIogWK8fz61lWv6DSAC06Rv2gkiTUMZyKFGWJXYoBs+Cm2JhS4MrI+T3vid
LN4Pr4H72UNxlK7Pga3r5I48sqjQZk+CAKpmDhfCnR0wx8ZXKpLHCQjfrXnDPM39
rUxEkFgmIHvEJLR7mPlDs71NSbaO3Fk5+jY0b/moJWBN17ADUT7iz+FEeY/+ZDla
IcDA0Nqg+zTCvxDZ7uAGrSt8lhYQ+PzhOURyXkoVPx5U79hBAREta2iQf0tQuuge
AIPS6M9+mGqaqKtJI+ong8iuGJcZGcONnLWyc0tB3qaZm7PBXMBP/+LpEnbZ/nA6
Qeu9ekhcEuGy/LhVBgdE/zIc9OvXXZpSmM0t0VVyRo9TcQpZf2y0bNv0t+Al2CtS
eb3gvmIfekPrcC7EcaoUr3uuPsMvHepLdjpo67Ct5TYqxN0+Yzb/gFuWRgwbKtb9
Gr5sSoiVoS10Fa/X4vwGTDpK/n/eWTjH6+F+/dkdsmfTeApdtrk1pJBTCnqrNqWY
jxYXbhMpRVPKmz/QZXu5TQjLbpX7sYVDq1btjOMOVu25RwzrpoZdObcxeeagD814
zlz/41CaskxdBQhOoQwAK323SCWAMqt2UiiKcSngWVWa1cZ9oIEMvqVDB6FTu5D4
+8SCzCzAqWZAlhs/p8kw7CKISP6sivXbpqRzm3wxqx6NjH+ktigoyO09NoYMAEaZ
7SnaX2+14EcDAvovMf4WlNogWuZUDzhuAIYJVxppA/9+u1zvqswN0iumo+O59t0v
szvC27PwABhzP3uel/B6XrSptW2u3HiS9rGLoOgC6T7XEQ/ZpHISqGYCBgwgqAGd
QpnuNOYAwKdgzdu8KGP3rGMSvcIB2fXBGngLHpvVVtzE3ySEWEOOHUSWs4UAesW9
RrANLziE8knhHHItUYCh7Jw4LJQp2iKsM6kMMrIuZk9EXpvZIIl4zaCnREUp7cwd
WLgjslHf4PduAjUuaL4CZBm5ZCJnZd/AAMfp26/KVanyCspJiEjQa29akTMUTEsI
d3L6Z+2wjx18oySeuSMIiuVmxOQISv3LJ/NOzJUXBt9/OHNAnUJpaRiJCTSBAdWg
gox/T9PnP6lAqDDUVclCAZB8kdAGqoUsBH5Z2JxzioIJXKVp51A9u3XWdrTQEZX+
LeO3ST71YGtbBy0f3rL+dBa0D25sdb3CXaGFwKBg7i/9youz+p23hI3UgKSqZdcB
ajQihEfnqITWj1rEwpGtS1qoqFBgfRS2s0tYfdONta16rVxZzILTdPo9adOTtL2v
q/aIN7jHmyu5BxioZkwgWdxyXKE+oqfcnSjjj1Rjp1vWykKXHzJEz9DJLIOq4Kw/
VMIxAGeYWEQ+RZt0QEXLlxN4Luv+8p0P3LuUM8tED6eJbNZWFHyW7qf94cnC/2RF
tBmuK3L6nPzSJdeowhFIJY3bI3hDbZIwYzGR+6cCsVbYfKRzZGTsAmsVyculGo+D
y42qA59wEdaRJw0yjVdZnL6ng9WEt21zToZao8eaN+TIQdhIeUBj8xOTCMThdztQ
47J6fzwEpsqa0GmuustqcXpTfjIl2hTqSxwzz/oj6MHvMb1Doa0jHLPpaOcQsjvQ
veUjpVBIl7QKa/ru8wWlTXzN/m1xT115TXjnU5cA8w7EoPG0KZZP5hVwagOsBQse
0bsjI+TOpXmAZ1ZcaJvNiHHS+lX9Ns0GGmHB+eobVRFkG7eaj1BaIyxrx3OKhVLc
693c/hc3Q8JRhMBWRBVVnW3mX4x3eQxW1yPMNJ33fqFX3PlHeqaZD/Nkvly5Fd6o
YOR7owovWgqCQZlM3Wt3lHnrKoeFmbGzZPht55JRgHF+2doNlXS5zSs5/RCcqI5U
UiW7PANLLGMahfTtSr8XFfAE/YOQp7YwMm9rq1JWSWCSiWSw0vTdiAL9QclNJrv8
pk6LcLMxQDPaLNR9dGmbeHf9TzVVy9rvvlDP0wPrsI5E84VHSUOeJgYVReWb4iha
DL+1LrYzhaTOQLWS5kRpA4oKeFNe1JZE9+DbaOJX+ItIZRmeCCZ5vcESb17mXF6V
kdLco5T/M5JwkNCzh0oMPpxla2oXGlZ8VoPpeXpMBTyEIARCWVKfMBkm6YxZi1jO
wAujhX4L1CzRlB/rSQvkwFn2gS3MsszbEouyeagK5s3FtUK9LzQhOC4Q0+7FU98w
stvELgxqRiWm8fuc/i1aw3P2+gtZurTAtxztNRntGQoIqtashAW12xUPuYpEmubc
OaT78r//gMIoz36ubgTMzu78GDnU/w8V2AdPeywAQxbTozkUhO3QpufgtxB+eEDw
z8a2dpzrIImgYFMBcebleV8w39csDS3Gu1Ul9ZImx/wxL5cYrFtrTv2lG9F1Cift
2SEIiJSarVwO1pi7D/932m0/QeKmeslGu1p+xXnwHt/UfN0JfzX85LTj7k+HM3HH
FjvxqVofvgbQCf1JJpwFzGsMrwttsuNIZiDIfhSmgnKYxrvo0Jn/8bOvjqnKA6og
ZO5cRC6QhvCyLv7omOHRPgYhbW51713tA7xHML9WR+4JaBKbutgM/hiv8WF7xyvD
37B+bUg98sp/b3Q3UBhn2a4y34EQgHoAfmHzTsHi4K0zhw2HBX432bOVt1ERqyZS
GCzvywIeiYYBpUnT+nvUtEmpTYJdG60pJpE4oX7XIcA3UmWnPnYVX/qwrcEE/FXn
vzR8HrRwUf6k/Opk9P8QfQKONE4nkQhlJdoloo+Txv9YqBSXawW5s3zzhXZ3fH6c
TuvUQrjZIcP/jrZSgSg/bS0Zh/TuBEyDXdzOn1d+dCggEsteGnm+x/DXLQ0kfDnn
fjFOCwSZ//ymEGv5UTAWznzlMK09+TyqStklE2M7BwYfD84CI4IVOK+j0hjkj7ay
jdJVtNzhOZek06EY4NUBJx4lqQoDVCTEXBvX0qgkbD3aAfMEtzQZvH/XqOEdWbdO
0WR881gQOMVAfqCQRaPBW6uFXVFjs8vH1h7tsGfdYFBIGGfb1IRLfEKBfQjoOgaK
6d3IwsCBPof5sdS5CaxVSX6cm7K0SEiOhdI0if8DVViEyhIuAg9rbyQEWo/lF9w1
aF8QC+6fmYSwtDKldx63QNxSPET1faaNuMV6lrFFuNulcoYg6SUUEqOjyEdGsRix
33nWzimJUtq5U6cfMZRwONgaFBeO/0ewDo5npVmRYYHxZjesnx8c1JMb1Sv/P18o
RRbRTlkQSMAjVglIRuhj/en3gF/VKddJ39BSSeiF/MXFrvpFIpKeYbiXg1/gmws8
eXCR+alzMmPvHMdl/SSwZAJjhKq+ImWgfozntAhBowa9NhEnjj0rz3IPvQ9WHCza
CzSCVqrvy6tYSBeLjMM98UrNMQn+1KhgWmbUlroRH0VMXBmZmaE9O1a3wN9kYS6T
uXKl6zKZtuiV8ofN+ktM+mQqinN/ATbzHsRLg4oHRHbY7yAjUaYj8u19QzjKu/BI
YBP6GO9IUHjuoJau3wSAPZFZcFtvULqrlCs0anJb16sQ7locUVIBTAstuxbbTJwW
6vnJyfKQ5ls3opBNlqPdcjfqmQwyvmPGRPsxMTNiM7kxU6fmRVqY1Hc5AKqnf1JX
aa9rRh8rk0Pgn2+ax90ojdzW9QXlpnta91L+GVZPMqjCzZPgIGLHuW58/cYT5Jup
N04rDvrYUr2mfom2/AZoX/hPVH9kTiVDJuJxBwDuNk1BvAt3i+73YXTQl3pCeWUf
iDWQPCqY+jptAaq8nD7tyd5BAVQz/uRbMp6IGAU2okoy8lgBnyGHIYNsMTVW35LR
tagKL52DBYZfcuU+Cnu+zx232pJSJ33q/3I5hPKsSgIPeLMt8zQCnZ8vnghmA6am
jUPzqvbYfprfNw7Oi74CaV5opR2+7O9go4cduvYWlPSpitVBPhwKTcJJv++cPmtj
zNRAyTiFzIN7vAP5d7yX5A+64aijKW1UsutmfWEfqeZlpAeUU3kI+/lg1Ar6PLVu
/Mi3ksRgsUjDbEZKxCJZwd2wAq3/1cwGNkG10+RVyVZY+LVdLI+i0nFNJHnsYGq8
rLJ7uxWsfcUbR4APFvhjvk/QoZG7AYvMLhdt917y2Cg0HYYsag5ZjMG0zjIa79N8
N39aYTe0op9M3rURTCOBUOUsTE542sAwrrKSAbYGGuuFKsWH9n4kbIz7KzIKAHvG
7KyoaYosLVCYAAH9bkF7qjDuFmbCMvRqDn2GsZEzP661DyjHn3uHVKlVYuK33IdC
QAL6fftXMVFIdqNtQfozArvkEVB/xzVR2mc/EBsTtHI9Cb2EeHU1Ri9ZDOrGV5xD
whUS3OmEUnNF6/qt3F7MlPmGRdwKRAsWKdUAoV+xZBsbKg00hf/f4mJpyqE8R8XV
N1Fm/DhZsaeFJwsaGSAB83m74eUsTGyr6HbgUhWDoqe6FAXHx2DZ90Y+2vIOFfJ3
hlB/FWWkyBNiFYoBsaSq1h/3WLCvm5d1HykPWY9FsXC2kMuqh7vYphWZRG5Va46n
SbpETTNVVlOOJefLBkHw+ChVfY0GETzLHacCJ/YED7dJnUILRQmDwuRO5ZyFl7U9
29wgv+RtF+Lx+ndDLqTyKz1Q3vfouOasmAQb82/Iwws/8XQK3aXZDwW0iDXcfbOp
lShtNZR9/HENOXJbi4tDsDrIfAKTSxlMLj0q0UDDgPzjBrmuChgF1wxHWuAIHKz2
tSBP837us3d6dbpWhRaPORCLY0pcnjwfgeOpmMmrZcp0JSDHA+FG1jeA9N1OSq+F
akRnyWPrzxdI0Yy/9jzLhU668uUlRLqVBwK+ifvuxCSd0cr57s3abpgJcFQj02B4
b/0YNNju/You3u1POV2IqCnZIuEyFTn7wQVeiojmEOmAoISlN9C3ZfKSsQwbP/z1
xRU7Ap0gY6BddlExRFLJRYrkEoVFmewbhyPWfVYf6BRGVtcVgvDY0Wttp9gX+8Ni
B2p6FWQUEHMMl9qdAsh7UKiwSnk4Gu9AbkFs1iMW3pqiaE8BWnCq8eExfVNX9MQZ
BP2zjSzzf+iTei7rswRFxU8ImyWyYIg/3j08IR9KgBD7pj8g42GUKrLFsxf9Q6AG
PScHCxI1IRmqUVC9u9wdbqkMtSyDLlhkjClI6t5c0kBTgrp/shdPBFfKScY01G1b
yvhLCyM9ALxNchBs6ArGXsXMfyoAcRyunqo3SksKjEIk+r5wpT9vTuhe9h911uoM
/BvMxyg51wFix+0OgfQqAmKTVM+sx+tRVTJO9KgfMCJ84J/6W9W2dEhplzqSjMWk
yQ9GKxQ7oxUKGlHeNwG317IPbIx/VxMvt55qKOmuN27NK/SENGnDtxEfnEfGudk5
mG6Dc3ffZRdXYWEcXwxn6PEVksOok7t2W05p27jVw6jU3qcim3jh38uc5Ii+MGCQ
rjnXfauJFQ7TXfhFlX2A8PxGbZZuWCDMRBbUi1RL//Y2FDI1xvFrdv3KmCJfAZmC
tIxu/0lR4xW6NbV81PrCT9aeyqbupqhhQJajx+fvVWB8MVUf9xquPifAAWGQOJFn
PcwcLrQWca3hOlzFb/+FbCki9zrni9ay0uvnJ4MQ/WJaY1kaAIonLHidvwi9GFUj
S9iP9He30qMEJu96/IS+mJ20thyQoK0eSHFl3Tb1sct2BTXqi8oT+7BzhM0R4Rxa
ignxGK61qCUn2QceXH+JjS+FJEBtG4rd+9mM6g2KRLZiENLNryYalEVnxWvlbvVJ
0LCwwQKSbWELf6O1CGKwLWgVKA3yJlI9OpdjyNXZ65HDnbOOH8+G1SRgCmrG0kYg
47dV253Z9v6kB2lztwsS4bsIiQOTqpGA6ooOURU/vSiY8Xqc5azQ9SCpPs+FIWbH
VVwaqxNc557HMBOetmIwKyewrq210hqx+CsyiNCzgtEnwQjFxxsS/S++R2HQil23
AeHqLBiWxqwPLM4i/P/rsm7+CUrs4BhY2nweFIbNxQqYsp345JCqyUaRlhCPY6nr
7z9VQvmCLLFDXghy2EWc+8Rgb6YD7qil1AVgR1LZwL+mrwgthCB0ezUUJx7esMCc
XZwlyfUCK39zSJe/gMJuxRF7X+dtKBlDAVRp4AxbsDLkCrGA2ZID1cIzDWguoVxz
oZv0mHWA6BkZctUmlt6v3R00AOlwHVvSIMDpoYLLCsXYtYPHcO6GR18QsNivhZxi
zJLBXFSxox0FrtXse4FfSWJ8k/ClLblRAaLuUXgQ7e0RY3UTjle2W1rRAm37tC/U
t1tlFSpvTbn9h5UiVZYx+2WpCOxHbZrJ13GeTF80BGHW87fiPb//+RtrOzatWAks
rtRnbqzxya1uJc4J7X9gnpxVvgE/pzrnZHMjqHXLrWz9IpKsFuYnGxDxbKNMN7Qw
V1dNwMHAjGfSvj2foc26JlHJ2EWudesidx6DUJu/U2WX3amUal0o9aLQXLFXu6Su
P7ZV14d0JYJOGO7xIkIJLggfHyZT5/O5AaP2DpxAA5hnbtmRbSY5Q38YSw1RP5od
GrHTgBqPPvGA4t//i8xV6HiBw1Q2HZX0b5VY71KATekVB/TD2vP1RetdyveGnuM7
HFohQiIaeb0RluLeWcLxM7byK9QC18TkZ17JDmN2Db1daVHkzgnDwzmvnToPdtCL
W6RXghc6KfcT0CHtVjhcifJLONBjQSkbTxH0C3xf4vxNpvUcoEy4NKq01h2he3xM
1X2IJzKIwQoNMKUDnIoIwr3WywrGu5EbR8IQ6daDVFmEG9PWLkn4PyJ7opMU9SRV
2IZNVw8xc7qtu2ysXTJcvlSWfYjf8mvGbzFPM42MZFK+jV8O+gHTqzLWMsuuwPPh
b8DVPHcc01/GgJ8cMYjl0Xfc5Yc7bWC2k/R6ZWMzF/Bk2N0kpfU4LHNzDz5zjk/n
oU6Odi+EUmrc+w5CTlxBO3L4b1mUPICzLPo76jPmJc2TLCYDfMQQxVwdEjpQ4egA
cTo4SqaBbf0KUtFkyK3BSrXVgOad8gXT4c5mXJPwpWLL3XhmSnvC1nypCb4BaDcN
pHX0ysdAf16LD81zWFQ8epXE8+lsIAFc2sF6+UtZov6E+46aEoqu1U8EzmqsCf+g
Xdyd/75zp47D0nkwnYjxXUNE54nSn+HKoaEVAfPAq/uFXgXzYytPZFO7g516GG4U
nZhAgbFivMsvtJ0wpT0ehZdef3CEUJBEf7qNeIbdKsGz5hLDtR/XiRbPVQqZHJXs
ASi+bmslqtglP31G/btWqmWWYLV0y41VyMi2qP0/hjJqRod0+Q3ZitFKnqx12Qjx
ICPD4GeW9DDfHzGRPOnefZ+tTnT8eMlm+XMnbrfwdsTSVgsOmEEXygskmZv2uasG
ICalPYxV3UI+Ak7hJG6xR6/5m6gNKkHnEx9s/tNsblT0scVDBOHt8h+5y0dImI6U
ndTBg2ghH5rwFAK/RL7m8oCzaz0w05ALYZQjbHiZjRU4XA5KBQo0/V7ar9G7DFOb
BYieYa5Lrim2e+8KA9JgiGVpenkMb7j8Iva4ih9IAaH4cuT/SdL0Bcsi5D6VfZFW
65WQQ9iUJQRQlN5W1hkND2W6a7fU7YyiSQl7o/5GuV7X8SZ5uHV4EnUjuvCcnIvd
CaN7Pe7j+i3wDfgVyW6dw5TpI+NHeJc7w86+x7r3uvx1ooKXIz/a27cLdlJt9b2u
gxC8KCjCk/j4+gn17osKidaFT/C9xIAwvW5ZIFg0+eWqYRI2S+eQrNAr90ynYBii
Wh8HS3n3NEL1lUzsL4+iw5NEivjQjZ83O1vkf1ZeFkE4+dxT1tG9T+dUxRESBrXU
OYy9KdClMFILDrrJNU2VvR7+T61lAYBGDMgQDekHM0+7u3ZL+WDWvrtXlTXhyOel
AXQLUuEZB6zbOZgTMqqwbTg+6Rry6o+1S6ogDkdlH3idExIGSMuhKpYM9M1MkMZj
cqK5nAdpgA5IreCIbjTiMt7HCoyvwapqdsmzm4KuMYuydDot9OOEPWfdlkkNRK8u
LIZCmPMfH9v9Q/ii7f9ZzL0psYWLFSZISq8mWqnSb8H2tNXm1Da8Ig6ogme4xBy6
PmEyxB1JlgpG0aVyQ7fCulfXgb/dltCeMsnGmd3QwcRNZD9ZnmuIWKZ/oEG3sEou
Krqyi7taYBAW9vt+LSfySGyHXJIEq4g0L0siYPo7nxroTgg0emAeSaDedl53kyb3
ozIgpNVTHjT3HF/6iwU6W8Ctj1MSKv/bdINmL0izLFTc5bxwgC68FbniopGsvCKJ
zJ4IWjrw7wDOyXe7uqkQrAlP9ywTKKT+FUEIejP1Fof7dkTZh7SHrSQYwV9sLtvi
04krgInhqPbxjeT7KTl5p/yt4AXYmQQNmdaj1qgS4rdM0phsh+esawCmNcCMSgX1
gcARyKT5vQtOWCTHGG7CYFw/Zy6zE1QOH75yYfccnrTLGeb/TH/LSBhXfsqtnO4q
xNO/vYNeOxgwrnFawssNktR/hOGi35fB3L0e4aHgZIjDfzulgzp6ZM+t7JvsPCIY
tq6Oh+UOPJg++pAURdf+i9Q+Z2ilWJAk/JGJw4E+MqoZcm452ysFuJnV7NrcCeej
rIfcAyNe65iCn7rbi2sMdrfn/wFntG8omJsPqUjRo/LebbYfzEILUDEBUEkZ0xxz
AfZ1LXzspqxuIugXRnYTa5ZZLs1e113v2lB+PTgc4dDgtgAtBkp9q0d54dWTRGcn
GFTxTEEI34cHJ82Ff0mnnOIp/HnQhJLtHHpmULR+1UuOB6Y7OZrcZEb58lmVoVHx
xO+feUHswR5+AESOPd8gA+yLsbZdpQ7IRmru0UwbKqf5ZOPNnTG7L/zE00kNIw5V
jswMV5zXLvEWKhAwRXMGJ/ijy9iZC5OuCZLNZShxSm/oqzWda+L7FL6T+dN/biwc
S1wfVwFy9h9gPmPzNSJez+1i62dl0tAJ9OwcLKwH+MTzTb1u7qCgCAgqhxSyJ63J
zVEUZf1OQ9p5vEFMJz5gHW/OifhGUU8TxX/qOTVG9mnitXZOw+4h3lq4KQLYAT0Z
gumxDyuhTrhiLJhc58hamhGvEbUH8l+BY+gMGUPYQIhkUPG0mXZ5nf3to5SPbgZd
R5UZcVaBsFXRmQBM/GT60yng4jEnUrZhj9gRSs+eyVAl4pjZ2jsH3LtYp6lgSm2Y
pt88hYHUnD7iXGCnKtQtDr/hUfJHdonXL01h+Tz01x94KbHWbxb1GB0Qbf1f6Eks
0hvXb8IVFkDyBGE+PJr19wT2k79sRaMbOOqvxbolY4uWa/nLgJvhCKGrEtjRUxnO
mOg0q0u6gzfnzn5NWHWfNgeFxTMvcQH5C6rq+Uq+Y7q9kTSZaWby0X8Z7criSwyj
cVpBefEpSFXKHXcLYTzB8NpCYNqkSXbVdYRddkVCr6Lgf46Ksxd6xlsbe4g1wIjC
fa46RTMGSyoVHZXZB+Rta735waZ/ecJv6iAV22eBzq5nb7woqcypnnmNPxW67O7Y
z890v7U7NhxPbOvCnEoYt2N4TpxUZikJtYtO3cL8YU/g4wBArwqe0mr9NMupyOBm
vHXMEG5fcaVhEeOyvIDoMUWrzFZJL5de3BU440qNqkJWP/s6xTdSNPbKHJcPxGYu
huKQ18PQoWDqL2PchJNO7Qh4N3GhMh7GGaWN9Yj57fzmJ+rYfMxW8IED3vVgkjYH
VEZh0utRtnDBvEFVO4A0LOuxB0ThtIW33K2meUnwNq/Jr5Ee7kAKD31Uk+ROf/o9
PEsr1N+5HNvlw4QTfs4JHD1zwp5pwCklxK/73eMdRV2he2Y9MJctGPPN45ucwRjY
lfjHNRxA75KyLqaqyyP+KqySMYEIRwyqnCedNEC85f0scXgPuuyuYWH5kXKJphzf
FgJXWBmjMCWxqbY1MZm9p/4+9Rhlxx5VH9JK9oYvgq8N7yyRMbU/x90H9SA2QKwW
tuhQefTr2O0u4nlC2sfTe2IvSnIhQTleNOZezRTCt6XDIN9xhfGPRFffBBtyGFPS
BJhBKPINMi+RUFduETGpqJzFPnvdWVTwOAcfxsE0PLYp7ce8/SG8Z1d8VdTZD8c0
xH+cC+7xNkL+zkWqclMe6sUonlumCaWFUYhLT1CD5ut9MXv060tkwa1OQHomt9vq
KAmFE3pcfXc2AqQSnZEniS2Bdmqwf52hW0SyHZmCMmWSYNvHPdIUg3g+NeuAFxxz
0xr4nbi2qQmVtOLG6RW1qwuZQgcSbI9nDUawVPz7p3NF9HQyzl48AlrGBHTRdUKR
wLABQNsaLVCiFDrDH0yY2T64lDSdByANupCDU2N5si3Xec/q9oDOCeyq7XutzOkq
xKP6gDEYSC1nDCg4Rchpl8PylnQ+9jJQv98TmfRbwCy0BDcyyKypdu/xHcmLDHOe
SVYB+etNKKSdrV879hdhBMS7RyuqFv8pZdoPISYhryDl6BvDEXkLmrECn7/WxYMe
w3uOHDXvy1DSpvP4NjIlNNLAN7C5uX0Wup+TWnE6ybPNkRx/WANNhdzKy3vAvBxB
6pIcl9k3zfRNy2CRFuzdvF6iZaZypcW3l1GHlPH6lgjmpWdc36XALiU6YbrFAx38
0GzF4vvwb8wpKagHzDyXAdx5hWBK9dj2Kq1AnGJxB+LOu1ziZgR/RA5nM6qER3Rd
ZSH99Uk3jsafFy6va2GIUt7jUWVwm8NO+2medM6/3uojPXuZ5kzykfd7RMouXBsN
JTIlTY55Ies8BazWkgFEZYcJ6EvG4ATvTYAiB8OvblOp5KN9Nc5upOu1l4xByNgy
RA/59isxpmd3z9WjCMiAZQBPmRF8+0iZ3z2++4q0U/Ef1M0Krqlra3WSkHHoA37k
qcTw9WV+V054/L5p/QvmrqsxCpRcNwYvqsz0wjcs99ux7ijVuuMrXW0Q8g0ISWlu
caQ/bOQ0DKT63/VnUTOQXB+EEPANsBX+SQEO46QIwm3o2SRNkV5wRy2hMakxoMFR
oPoDqz4D1qilvoMCD3rHM6fZWVNuJUzAz/hZh8Khd7TGrtTPR+YQJoFtgQ/aYrJ3
DZlWbYl3iQ+BSHQFyiga8yD9RoUWGfwDacPtleX01Diq2nhjfYq6YRulU5hf88DN
w2lmRcQsjQt41a6In0hlwBavhaLLDa3bFzpk4DuRM3YWF5BZrnSKvJH6HpLmFDCj
GQqD1AT88UQpLkUmM8uPpReGtiZ+zcpZdyq3xVjS+oaNgVKhUAIPmkkDBcsNSSTM
9ZnC5CAD0Vqgh+/zpriAAahAYw2EAsD17g3jnUvXSDbLwODg+tVQDQ+IzgRm1Nrc
DKaldw9h+PNzzQen0Dk75Jcap0+UyZ5xgngRszrh9zssqYi/3k/tE8QMbQKp3i4L
XRNjBh/VMJYhYhOQpzfVr+yoFWR+iB5vwnPKyqiV4rrFScF+dWpbLguDKd1yWp14
a8ogjGSDBawbYa4ntm1+CL1Xb1tVU7xpPGg4KblidU9LE29uPO6flDXLgMDt5llA
8CkXfivemsd5+Gn+/8V/vtCwdVamH42okHn21N7lRoiIkA1mbdl9tfqRIsT6dsI3
jBKSNUFOwA6DXgKpAVt173pFAPW67sNppBfprQ6zmL+Hx/q4X5aPKjLF62IBw1QS
ua9k013OjsXjfqEqATmsBiLon0ZNKaMFBICVtKbgho5NoX69RVVSXWowc96u4KBo
wNAJKksnLV4DV0oI0Lfyt+qJywwnDUssXnOWbCtbUL8MV6puZ9sH+6RuuMloF2T3
42u6I6S86R8YPrU8Kh46mZYICiiKzoi9l4VhIJ/QQEygDookCdMtMpdXlfvkmK3f
NpohHCet/pHS6IwV2QILWxW3AGAoQvTi6tYX4Hi35LXjhgeLU14Rlzb511XWBq+A
6w6R6QFdPlS/gqroZeSuSI9yBdGcQlg/iJdShqvhjgepb+baTqvFFP80XEFIGbds
4ap2Eew2DRVEeOpNXTmxhd25k2iVqX+QsTFscs9M7xSpEmsgPM9syI9YF1ACL/BJ
OcGIkl3S52T1ielDqibEOq0BSObjun0UCISBL+4v9l0/cyWy2IQfD/yUAIRiMxHL
yzHMepK/CS67job1aQWr01zJ1dDKXR7Pmud8YcPpRzbUjudICmagnvK9CefQ1PRh
obnHp9v4lhmVIV8cJ3SMkWGoHZFCN+fTS6VLdL7gjs4yZzp706sBV7AAsJdm/ZEe
vfCw4Y/nCCeJ+VbNtp1MBV83Cycd2TlpNx8kumb5qOcxdi3Wj5UrAS2PgT7rEhKj
gF/8Ei1Tg6bvWadIZmSjkf8wFg9Hry9Gpj6Os9zXulX9m88EmE+4MvScX1MwDzJ4
4g1EF8jmDlnqkKEcRWtryfh3cmK1m+opz9lbNK+FOTdwapY8QWYKRjOVpH+2MLxm
36wgzuEFdGau2COWn4IDBaBAhK8bmVJQzdsNGedsXCRQoSes2EwjLUw81wJDFOKB
7cW/kft+hVJxDLPMBMQCoAeEjkbULaG0EvSK9t69Budp3C/+XWjqG0E2vMK9XOdG
3vsdhpf914B226itkCCTDJvpY4JrsXtmBdXkDIBGpdr7hTWcpS+ewveG3yEsaIL1
KQw94w3E35UwqNCKHjUVLmAEYCxoDjfd7xrX4WSpnLyHq/iKVskWsWf1Hlwd4211
zFkF4oSOvfoKr2WtmhQsUn951JN74d5Bbp1BYtg8VkSMa1I6LrIYt0SdQwnGI4bT
hbgcgenEslMTOmW5AG/WSmCi6gF8U7qBjpPRR0EG9u03oQVMP8z2S8OZoQG3IT0L
gN5wGp9Z4FuML/h/YQ0c0kE5OtRX95+b9uAWteSFRlhK3EDb5QSauYiYfx018tUx
1c9YlAizuHcBYF503ROiTMl9eIxwXkdGd8XnAFT1b0Zddfmt5it8dB1UM2rXMWgt
9k4nmR76izZ7+bwSw4OO4SMTQh8JN7ACtnYfo0CcZvSBj26QfLgYH0j3j6E9eb9z
0jLw3M9aNV3XGNfLaZL9hie0Cns0zxRPlfBUe9YmSUcnMwnyYZqF8ElWduILLFzc
AZFlC5xuEGw6LlQpwf8F7bviFiuI155JXxfgS1WsuN62R0zUcNv/k7cnHWFgWLiY
hgC3Aldikg4/WZkmJKSoCP7shNBcRyUTj/D9O9qHQz3P3Zd8RWrRNEh4PfuJOvWC
oJxBm0oPhsuSN8MOCkhQ2GtCowAjK9BRIP8e3ZlssrxBUBPrqx30VA9SwEwQEsAY
dUdgRPT6oY8fR7dzNxLdG4MHvgt3Ps4x3dG3t5RDnJ8kAldUxTK7JhJPDg1vBGah
r3sknBLuUU/m3Z+TCfRe0sfkyNgAq5j7iNzMsKwHi7meYpvXSxGAuybL6Ar9VE8v
rImzGSPc6zx1ScI+JIvG7eBo4puDxemKyykhyRBPBYTCqw84oC8UNqtWOO4OOXTV
I064naH7ALIHJusKlEnda4taS9W9D3ZrAnmfAIHoJ0Koe7yWBXkmGelb9OoDPTtN
THDEDFYpM03jQIX6e8yLr8A8Wb15++x9Up9rOXgauNllOLAdi18adtXiUalEkZWD
VkfgGaUQXtA9MhKknN6taPZxkgAZR6hDndZ0oxeK/3H9v39fntDf4Txg+WUahI3b
fAM7rkeSGJpT114wbo4e7C1Fw/ZoaR/+NzoyPRau9vxh0k3MCkuq9ysJEEOvmanI
5np7+jtHnwuB/vobt3n1UiDyON8oHYyYC2QYf11GYoD0Mj+ACerL4Lg0W9taXNsp
0XyC56FMkjin40IDLagude9qmlD6bLudwuO8wuUxmD9HK+MCb15elPbJnEOqbFxr
lU7tU+E63fL2VGJLi8PoyRkBqA6I/WNALM8TFPS24HlkCMMOqVs2xjpXDnRGmcQX
ODI9hF+m7ooo+9MEv9IRJa4QZ+QWEDe5+2rQiILj8LXYTwcatsi8+Ie5qN3JNkSV
6Gn98JyMHxwvILp1yIMM3rGT0I/Tmyj10bb3FKRbnPFayIAq6cmQ2ZOApkQSJT40
21E62c1GK9Jgmc+GvlF+pjuKQxd3Scwr0rx6WXmx64PrMNZ4NXyaf5ptNIg8rcBN
gWgsPCtH+bW2XnpIxjkdvEU6EAyEs8ODmP/NXcvon6P81QTZycgIdkf5ekKLakpR
EtNMlk7TTOrqZ2QwpKGB8rrlD3c0izhHLgOk+mBwUIHMDdC54c7yjwokr37+pE8N
eMobPQkpZg6gyukdRyp2w3uXYQdL5u6Ks89aFr/fICsgeC1c8dc77f856zSvf+CW
6qCXJlWy9P4J435+avgrWKJ+5RMOb9QWp096eU9v5dBKxplzK9es3UHv9RdyVQP5
Gu0FmfZ6Xv0L7iviAgJxjPxKKMKc7s6Dhrf4NaRwpUJtfVo+q6kgpZa7fAo5Vwpu
yk+/b2f6DPXO8o6cqwrmY7vobpFwhDBgejh5jiyS6d406FusoiAsaBpIphDCAzvO
kyDQ+S/WiAGiLqRoNeNCN2zf81uhMTfdF7sGVpkT8RcBdp8k9FhK0zJKdXEdh8Lh
033sqJGsW1XL408WRTQejkGIJngg+g4920GglfRZgzIgKbLg220M74fEcCFhiCdS
m0YzfBFh07WkVkZIG4aN+7+zJyaqjycGA1z/tbk1ZD7Ao+XgvKkvsMeJnDfzuTKJ
nleTZ8dE2mH11OYeR4Z85ALb0e/LwCm8/rGw7AyvF1PRHusT0VgG/Z3BrxbJQ7pm
LtK4BPZP8/3PsZ0mSp2DJULLLFtRfOq7f1Qj0yT0Z9JxT3ordGHg2SkuYZklsg+a
nZSt6RA1bxsuDQRr7sqsi9X9UfKEnzxomfEeSm0C7TRExnIeO87WWYlL9iybbMhq
Q6vOlqpfjRSm270wv9r7nLQpa4KtvD2qnG8CoygIN1/w6CgzuByMLKOgoCGCdLAO
wEp3mdJezGJAApK/51keh4T8rwYdcOcr28n+gTbNtuOG4arK9KHnS78o4p597JAx
NWMBOEgdSJT+5wo8mEO26/hBXjW4sc7MCB3VvS/hKwO0nuzNNWGWsW6PMvK6S1KE
uqLhFaEtdTWp990uudQwbs6EO+SppxZqcztwNy0tgYFoz1ydXv2JtVro4XFjKA1m
N2ze/dNdr1se6/I7/kJ6pdyu3NlMQEYmHS4jY0TpG8LF7qCfYv3rscd54xNEk2zm
CkQBvd2nIlJxES/RqWAyGhvnQ4Awzf+qzwY8sXuEUGcyGUGHzSEYXQlOwDFCKr/3
yANl3wIX+pXn+W+hevnQMZpIR9mG0E1Hc5IeCCEY3WiYACgjoHImDWp6tL5NjAgR
9GFYAch/R6j5G/zQbb9dQzxMtdRTfaMHmvxg2uVIbLUSyEcO+eZ+yRfMaW7DKLVg
h0abAU//3M/qbo7e/Hi52mLPUV2G+SxIit0mA6rZr00OdK/CAGIgJoSEVpNZerFK
bnTM5WmehkkQI52xBK801FiojOaKm+HtwQBReR6+LD64VE4ZNrDx7ZmvwoBgfevc
qqvyEDAn+VEoo0FxJlt+ZWjjflG1RqFnCRi4rHSgVOzvVqjPdw1i5aSFVWwd0MXZ
gEXj/TzWLVoSghFqp0CneS/JukslkUioWqOUPWnn4jgO4cbJaQ04rvS8fla+kOhB
i6VtDN15lgUjXTZRTSF4LTKEI+CEcWrz5nWdvS/ki2PL6WRfQfvqX00T4nU7qoQH
6m/urEZfgLFoZixt8Bz0UWNKn0jIe4je70n5N+W8sOmILnnUjG4PdX/+AkPeauDS
fu0EH87eXecu/rYYBXT1YF2adWoJor26I55fNBaGnLpvOVucHd5tXMJzEnsu8jce
D0dcc7o1FX+clakkUgoFuHqQxDefeQHLFHEbnFoPar9l3ucIgYeN4he/BkuT/B+G
E6e8l2PTmedY1KPuQtDaFy/KRwhAfLTt8Lk+fowX3MS1fSnVLFBnkEYGwqE/FIQv
X7XCMlMh3JbJIEXzGw08auwtrcoqP1Whz9yhNTykc+raVOjDEcqbH+jCYPaX+53F
rJCWKC0qsMEBNSWbkacu83OYjRZppik45yACIvcmYmKT0vGhgp2n1H9BGno6wYJE
pY6JF/2wvbgMxSiyzyYrrHZvyAFq/MXxTbdIKHgZ2pXclyssZ41R4jaPnlmBXDDY
Dzdi0krK+RPZdR1ih6TgGJIUKRq0c/MMoJ79yRCSW+BoXkTbctL7SezxGaXPtPn0
mZjDt2Cr9pYn4W81/OLyX/qJG8ahJkRZo5U+YqRcOnCywHqShRWF6kDxN3I4cUbc
ZET1u9xUYCBKZrPHvuQ4brzhBS5Gsck9TPEFTTuMb+0+IkoQPP0ormIBSJsZ8J1U
b+EJJuygcGLjudMHGurr2yIfhMHk6KhgGYDtH6Rm3a17qw3cxOfPH7hSRh7XJZUR
90sMqxaPKKOR1nT/YEuUuR3nzR32sTMtEHLA4ixKchzR5/cHo5Lpo6nKlQg2Re6T
x/MWBSZq9R4b1RUjV4d6G0n52pTgocQyFDuJ2WfUEBp6dyDwDjRc5KMdC7cAUgLU
tcm/KiUUlaJmbvlarQJX+UEthrePH8V8p+hvdjAAmh+s9tinu3PLQzKhNy+S4ng+
PU9OMNrDIZz3KIQgBiLwsD3gMCcNsB/6YNsi6T1wYyL9+aiR8g1iYCX60xYVOaAy
MMuj/4tnexwBJx1jg8vOD9IUI16KrqhN1ojAweQGw/IbhfOuiwS0jyruYBiHkPQr
vhBRtblTCf8Fs+GWK7m+1CrX90KoFC5tUIACg0rsiPpeBbF5pZITB9V36Kl5uAK7
6YfVgnqjtgSHsSNdHYXVvV0jBlX9iiYCC+cEU8WbyxYrEwytPnGCQWVNpve7Ic47
WIPdHzImKLIClzaix15tR7TSemqSvV8fTiQL/GcA+3ACKIs0LeUpWiHa3akzxyj9
1t6sNHpEOhgjOIMEKEfJqYLoAkXa0tHo7i2H8VQ9l6ZIAczjbc3Tqf22rTmBi5XJ
zJrURvjTGLKLM1/RLAGyeHfSVWe6Rjpjeqr4UMMJFtnbi2/sbfByHzNeRR/HSHWS
1cNyyn7vseFY03D2san8cowueCYqy7vlVxdUu1RJivfbMWIKp4njeMwqVKcEOiIa
ac0aevWK9zw+KI6GEtqT/Ho6upAilUuSwe6uI6RdyjNJ2S+I0uTM7Li4clRPFbIw
UI/9HBIaKwR39E4MaSdtT0s9YGHKwbMv9aR4xMSggw7LhUQ+2KwistNztktd4zJV
gVfECakTvmvyqMzAXToMHz1Dp+1lAT5m06sQwLEs6l1ahGDTE9ajWarz8HJXVcpT
7SsBIdq6nOo3GnMGQpTcSrpJlOV16R5rd9fgBzEaN4LzNEFZ3K2eJAYqB9ISVoUw
6R6G/L55rZVOjQH1TDnO3TVvFFOURs+WB70Qzh/qwGwSUtO7bY7VwXwgI6Hx90Dl
XM2/BeVgWz9w2LLMMXtQSP5vOCEGKD8H8/4xy50Bxh6haa/T0iesTAbOhUMtVtX2
Hmjwgf0ca94lNadUldEbm1+1zO1ONOfoIAPhmgCNMd+8BPY/jJRLHo3JMspt8yLI
aXnYSPExTNHsep30T6CyrpZSo/IdDG8uzxljeuYsi5qpphVmoQ7Xhu9gR8HTr6Vv
/lKY5BCQKfuf7grAq3PoDsvD4F3efUNUOysv4WDKOmMzCO/yBqz4m6MWBeGb4ab0
cScj+VG3phn1nVx7eDfI0ekkekU5I1qx4WOeWN8fCQu6H32ma91af25wXSFvTD6U
AyMGXInXjWQ1SQb+tMvd+SXMrlJjJnb9g68a8wG0335pV2K8Wv6qgWCNEG9OIX/3
GfR5d2GPpJrk0u/IBj+YkEJe5O2TPFIewBYhYK3uBjsttXxMXDu4JwxkcKpKaYR9
nbAP9q62I8ku6V34Svcz6GsPx0ClwXwayUxLlIe5xYABBazefXKhrqy5wEM5fjNL
Td9/kr35pG8pUL59Uz11K6l6sHp6SWsiAi8rNNmFq52d1C6kpLHNqe/sE8kpbcN0
JburUCaVjSgYCvL9y57ZdIydzXBGtcAtJpeqZF+1TcZ8rrOIWOQ96ItCPZYDHne+
xaRUC3SSD7/Bp0Usg4yT4hm+9VL49v5UrPW2RvL+S8kuBSg/v+46h0YLfO4kaJep
AZpG6uAPC3/IHF31gNDMDga9pQEI/3XRFJGwcDlwLaLs9gK6EHqOO90BGXhN3IV4
xrj2DBhjRxZzu4akk/nq7WNGw/+yVTB24w0sVEf7xcBPu+VNplB+8q1cqhnkI0KS
W3NKitxFqlLVWFJ6v5jjbpUrNvf99fX3B72mC1R297TMplOHRiyxeMDPq467btRj
t3CYl2Lj52hfBp7N/R26jzqbB6FCCK3rg8JCPTYg8Uev3uNIYH9gRr4GnJ+uEVq2
dWAG+BhIVoRiqBb0FdCfvPmVSNDEUkcpzViC00vfuTCI8udCfuTCY80KgCUAbeaP
GBa5PtWFsiXz+HtZWauEsg2iwt5HozjoOVHWn8twTs6MshF9SMHcpoppGkWyELna
xiBcrxTtinFLV2TmC6MFT5N5T38dN3Am1RJph7eftCZQJRQmiScwGEd0EHj27MbX
pqwseyZmyXPuJ/zJGShEBKp8JGGlUbbuznCWUVkqAee6WaCr/EIzx1gm3TmcT/xI
4mQ4GeE07hcWEBvcQ6XW6j3R6JhbAXcAWmFDHZhmNCG1nika6zqJWq7JUIU/tgTm
Sri3KmLWyW0IPYWzkNt7OcWFYjjE28p5lY4pE3icCFMWUplyxjnLlb6rQTq0BQkE
sfAq24D5W9NANVJsM5fJhJPp2eFDgqRN/WCEfm+fih+nkmTErnM4xFb1K2Kl86Z3
TTrBnm5Y8NhDQFZJOPUf8FZrpyFCTgeZ1medHpAjMLdw+wbMPnW8nDjp9DgdDbGn
lm32HC7yILymk6Uh8y3YGi1yS/mwJaui1EqzWWZtZt4xF/nmDS77w29eBIgDRuBe
NrqRA0dbmZHjgWWbLRrOfIQRCfAqfKNJd08USjrdd5Qj/wSl7I4a6b7OzU3EB6kZ
GtBEAJrNrJwFRi/oEvtl+mYh8ev6NfZH47QBqXjUpitvYp/9kC1bJ7UyVGk4ahAM
FfyzinTvKDkRxSWpLR+OmYQHTnPcGatCt8bPrhkZSuK2iFNO1oEnIRbgIGeSqQR1
P6AsgWvcZB5j6QrXSvK/wYyoeqcxc2TP6EOoxAYC90W7bch5s7kl0vWwJhvd9Poz
7JiF7o3l5oncJOGmznKtAIhcGvLHzjfIsEws8NmJHeeg8d6PAxd6meZ6bqD/375f
gN594raRST4qQVBPvN+a6dqup/+sYWl4ej8jPDyLPaSdNMppGMuRtwBjO3vzbHMs
zoAPSfIneC116PNtLdNxxArVDHk/36n8bjj/gMFpXYR2WmpIOtunMSTPWz+uIAfx
+9SHObgB7pLjQehQGVi18N5ce0/MLvU7AKwplH6npAqPYbGiBQ96vZQ4SsyDCV+h
D2GxfVJtlLYFmkYPd/UJVBPNgD+1hTuLWc/sHh50S8xWhtV5wLNvSie0Q3UHXfFV
jgzEgErPR1LdidDPhaSJ8+iYxm5fSAxK/Hxxq1mq1JCFhiy8z+CKzXBwirvYoFoA
4EL0gK6XrwPQOSjoMJ1exuYCu2eTOV3kH1yTkN2rdv6Ox9jYcs+eN8pmHud415gs
TNMoVOqEoUBmFfkhkh1MNsHUddU5zFdkvhqSJhhCImoWFiFXQro/XURw2avNuu0Q
LSMhJVE8Gms2Np4Ng1KTDkOK23wfFhwmL3au6u4M7mDCaRa+HWEtlbdnTDD16aEx
R3Ycj8KXqLI0nM+hjQYqez/lpS6YTehKgXbL07GOTrAEVoXyT7C6b63SkaLJqjvH
tjZzHhYThOQjn7D5Bvj38YsAefPIMTAz56awCVd2C8huOwxncZfBAZ26ht0d8jA6
YhLxWW3xWXHOid0NsFx5jOPl3ewFgakD42Npf5yjReGJQKH9N58LqBeDcKX03VJU
HqzlhJ6Vq7jP/oo46pUbnoZAf4q+3TXqqpz0w/RzaB/liRNeHHzquraZACJEa2pi
p2p1J6exLfUB1gpWmaYUxnxCSnsjCcyTGqHtbgTfdseifncj4ypk7B3OPMe37ad/
YMOsZcZ/ykdd27izUcISiNfqtqK5TJH2ltN9+TZHIkETmeg+2tlY1lsU+UsNVXwR
36Jvz1F+AA/T4Msr1wX2mIsjYnRcB+K+/8W/HZARo07Q991mhDhwkHh0FHuYhD9Y
ubLp+bfwMItDbdQNPA4gzsnxxaid/a3tsOmdjD0gDyprccBFQNHovqTVPkYJBHq7
fOJm7v3ty7sBl9cY6yT7KPYrCRBQZ/dIcs6MGHvIQgA8ROcn7iojRvnROQ+ReBga
YOF7+Drz1vZFaOiEPeNebKeKr3hpcDCM3y/NiFmPSCEz4YyLKo4tYwcj2OiyvpLa
1BvhSblqd28K4Y4sQXERHcKRoxgSc1766nmbLhfzV+uutwxN6lLzV5HN0DnBiBLz
B4ifi//AsrsWBZ7nSy12PnDYfMHivMGsrl5Va0XkVkOhHmwJgxoCvXLUGqj6O/w8
xDcA6WbIr6HZeBsgxsRfPdymv0pCPJnjZJQH0zXMb0qKWplQLeETo+oFcKnkhI9N
Fec4OtyXe4Z/bUnG50Umvp80hGJ7AL+Obot3k4gEq3tf/khDySLeZPd5b0AQYK+n
FJgx32006IA1L0APfeK74rV2ZAEcjafU2qwN3eUM7IvfZblbxdbiQ5epvx9F4F5F
tPxj5ehoXuYdID/qgv2RFpLBUEk4QovsTzgdIrDJwRMA5MzyTv4o1DzWcnpiiD58
AdexANAv903M7C3D354xDN4tVODJS5w9OXGh+cV45yB56R5sBOlOg4D/pG8RIdev
udX4iMpJu65D85tZ8bkIqicYBgweWJshH73JQ4OVHk3MRMay8RYSErc8L/hoqdw9
lX8HB92KVRlfunXzd+KaU/FNlfBi+AeTF7Tshw+4izZ5gOH322RVxgFFQmMmhIsR
SlNSMVDYhiIJ6LFQyZf7czSjC8yczJOfND8nM09G4obTEgehQx6Apj8lrjp67oQ+
oDMeMFeJjfU1Am+WjWgKH/rGOrG16urK1N8A1JdIlMxK1pDFdlG1uR9LNRyzm1mo
xG27VlzC57kWSUaWV4H39NbtnURoxz7PjfSNq3utO0q4JdjrxaiPhFx0YAWw6IPc
Acf+OylPGQLvNGUopPe4TWtADb5tK+iAdiFmN6ALvuCYnUDCEDwmW2D1mxphPxJw
NzGPbD45yxeFkdlQNq0jBJEVbvRQSjguJvkLQTWZ4k1+uLpW5ByCbfahX4UcRsNO
kOw4dBATrpUitUp18qsNU84o9Df3pqqqZ2WAqX7zMNp98UrLwKmQYLKntKo9wOZa
tIn+59eviK3hg7M4PrbrHehsSOoNC7+Lwn9bW/Zvhn+My38CwfYwaTFGw9+pOcfs
Fl153/W0b1j4Kz2aiOoNFeS7LaToakTAtTy4wvvLoja0OfYzQf9D78aSyne4HF6m
fNeRFS0Yevd0DMTHbRwS0NrZmGLrmEb87Iho3XRgBOK3pK3IYs/LuP5f+wDTVVrQ
Kzk+nJL24gu0VB9gdwRo2C8ScJX8Roc9GiqsKGa/bWJDa38Yaj1rZvFH1gSD5Vhw
DLgBLUIqgcPTARtD6EU516x1m1B6T1mzvdkersWHmVeDYyjxCry2FACGCba9eEWS
kSy1y8vdr4EBrMc6p7c4H6DCO8muxIH/yb8smDDqLtqwXKppRJUPYxMCsbjQr63v
3TigWW3XYdzhJh5hX8HmSw+lQblo72TacTqjsTczk03plmoa4wTUKULgjMhn7MM3
Zc2/PkzA8SRSsloGeAu5K9xbSqetZtObHZ5azcoUiBsx3X10A5/rkdDaG94ygonM
VgYuHZxAOI4waMNRwd2oecyJ2lpX8suWxC5ccth3IV6NhzwynOpmhSSJ9R9aIIDS
MEQNiEkY/tA6sOFTEoA4P5bdsdnEA6yS15UoPMFqngbGVC76RDIcrnT1fEy0RkCR
HQDbSOcWG+5WEB2cs3dkdGzxDMIiGDvloHlLMs4SgMAFo7SMaAH/+CzKRN33wGVF
wXUVFAKocDmlCVciPOm3h9cQUSkfz2yHKfcR5MviGaSRzd7V7fkU9/NdMDNJ+n1E
YUBXoLFIeuUWZ1/wxuYtJnGkH3kdXGTHKOc9ExBdS4cQFC56w6c0Mgjz5MvcENBk
G8cEct0hVWxx9EZKrMudmZxiOBI65zh9cc8e/6aLwBWViJ65t49srdNAyzWL3cBN
w5XEA60u8F6RYN30ADYOq8InjEYVphZ+ifzZymt35Mn+WCGckzBuvVkcE8Fc2I+P
n6KF7cglOIGXjzt6wFTJ6nDHlyQLUqO9kfibDH5n5UgQ1GnzaIkc5k3yVXU2QEEC
OEYkYZV7FusWz/O2TrQ0NDePt7elPoYRztVXS432wEKYoWJThJqwBgmCKaTghtgd
JInboFyOFQwpCY8zEdF/ipHdlBYI/JGGg1tBObk+tIXuicfuoY7DU+W4reP68FP8
rZnHsqtz4WlVG1PogYcnZROY2YBjYE7mY+rM1+oM1MYTdsIDilDITLGg2ChiJDPO
/6ph1MhVZxqCbPjxfgue3fvVkm4plb8Nt7xmNV6ZLpK83yQpdH0xdlHzTazBYY71
1QJP5t79YvP1fI22n42gmPgK0I7K41JhABNtQMeaa3OwjV3cdZm7WO1kSQSWIMVZ
jls6fSDwlXDquzJxjdG1s+D6c33mmgU0tpTiNkapBifRUX5E9IjJpv348fE83BtT
0MRTTXOyP3pDa96IrEdqZfoTBvn4oJNrl7XsuV+LOQWeSNaO/NnAbHtacm/YjiQI
zkwmbgU5Vd8gTyv84r9jvyaKoYX8UL1oF6vnmLnuVIe0MjuvE8lF/910icxaOnXy
SoqiIbj9gp2kXksOq62mB1Vf+TszmNWy3gzC+KLgm8c0rq5ojOhxFZ7RcdLKrhNh
98w93ZBC/sn9ltPQUXP5zLMHPqy88GLStDEXkPnrwczipKsiMqRPz1zJ6Xli1Na7
ZGg0ZAwG9o9UN87tqWd/UFfPxyBnRRuMi2BDA/5GPocCyTGnGH1GvNp1Xm/7qqlU
odbtveDJLkvR2vAICqoom16rWAibTxQRiMjHxL2Hm+GXkPqwJ/bAVcI3kcjWoTFt
2VQWXsD8YV3zpviRIyu5eI4kCGzRZNOhGXpjm6cNOM15vdN8Yk5ClBc/NvGlKU/G
QvUHJ1N4N6R808zyMeA7/R9ur9ZjF0lO/8pl5fLhEQOCY4MdtQzFGfC93gVCUDgo
OkKsYv3btjCLXtQpvow9J2JB5QHZuyIviVSNSu5YuY5m/S1NFjLgVnVBnRRQOi6+
R6usnL6IMp6I2yLPFHBALIJXU2O2AJ3Q0D0ZKbRPg+2VJBwr4cjinKEQ454WMPWI
ZpQWwqDGWAprmxPXYXYRpHc5qdiJR+fvnGrRkwMprxXi9d2u3MsOauAe0Oi9jocK
Fbqk+brSnAs8qFB73bwkN+k+3S9cVNCNWkF8chrTnn3fwSrgkbBxQBytoXO3JhOI
8yPJmhiGxrnPZB3ZPpM+6ZuvDu6ZU8aVU3XPR3UmhjE4h6vx3moozHTfmeXie2WD
j+h4hStWWP0vCpYUL3zOx44BR1U3RnSPefJJuqwZmeZY4Ly8GNluZEDQJDW8sUdf
qjEFKMKVX9TmAhj7SSe+66Eo3Vaut6EFkW1ZVANNYXqx4+V6b+qPXj1tC1/nJo8i
HBJE2ZMm3Ny0qD57MneykcJpgYycqwruLHht/urYOlJx5X+/hmSVVVeCBSukjGTH
vu0CW6+xg/N0EdI8QLs2QiSbfmy34jmTHB186A0PzhTONvc2Vm9d7Sv3gzgZtzJK
5gXxEM/qq5Ro+vN72pM47/m5UfKMun/eTASIPwoGhr2WIfztv7VLtmOW03TadW/S
HqKl4HojmwsfjMqSWE1flDnCjCuETTfGEpKqa9Ab1AcSNJ6n1sr4Xriv8gPyhuWf
AYV+XmdrQtGoAKJjuAGyAjL17wiuj/7lwFEK5Ed8hw5Y3vVMNe1SkPJnPKXRNizy
pSdSvn5QN66AHwchwG41fRRzUu1/WYDBJZVDzRNFnZQjSHVEb0j4BgMDVo33wPVw
wwAbVziCyDiQoEbdC4FBv9+9CiMiCautkZ5uZ8gsT9jfuqkEltR9zwAZWMtfKixK
ba6BtCa7LfFLoqH+jWpBDogmdAb2FGB/v85Zb8pRBOgZE+ZkEr1ptC5I9O4Ttk3u
heSkwRSFpsqJHflnObHPC4gLSg4fBqiWMlYR4wu6YNOakJzFFWdV5+aag2POf8/t
Xm7AadEPCgHzhzp1w3qr2LJmG0+hiDrbPNPEbjRFLk4NM/nONk5KzAlfRJo6eOeX
FXcc+8PJhBRjx9ApEC3Kx0ztmE6iuTCvLa6HDKyeajDTRz6s6UAkoUKixHKw/pRm
AbKdFB9FvLAkgi74Ylh0paF1H7oPE2DISApt92pPjMpq7cLIb3z+1NFyxZZ+f56+
t9yxNOWFjc831jmI1XWWf03lHcQsf5LE02MHMLqSrANNxAvbsG9SkaJvPf6qHcjX
6/P3pXlJ0L07068sooy1OotgwslYjevgHW2zRZReKcF6SYtZD3PohLHbhtge5Ddl
4PLQzyQqCED/qWr+TuSKeV3tUmP5efgGaQZTXU3pjR6dhTpkgDfYf76tQop4wKBC
5jKcRjlov3Pu3ii4ZVSdGkTyTnxY9aTWoFKmYcFu4TwcH3g0daYfg4Cd8aDb2y/x
ZqPRPL6RwrOLtP7iT2LS6EwMsJFKmzkTQ/ehHL/3JWpgrOnA1PAOt9oC6aBqYCk2
/rY1L/j1w4SyWHhjnGnE6v2IcXWK+b7HLsBqUHw01PIsIsF80zpiMuL85O7C5SWe
4WwMGShANw7m8ENkyvE35983rwo6F3lY47PumlNQfZw1Tg9bOmeKbtseUejuzql+
cbZD0mNNMGlUN+UV09jjx/SAtflbSjSxt11vrRTExL5vySP6ir5GYeDZjJlMfz9B
HJDIBeUN7We/R1znw8o+6NR96lxhxfur0t6jhHYBQuQjpCGdiyOj/AhzQJiZ1SIZ
I67x6OauLCYRBsBUhio8S7hyrNjIRBy2F/nYNjTL5pIgLn3bHBCHQL6BbI6phJW7
FrWZuFwntETu/N9toCTwh9XBgvFcGTUW+4hepL6XVlno28ikv4pJMiOr9hcHIYVo
HQ6HfRSr/DA2S4IJUC8sL1L+W9Qxp4IBsMGejot1OBp2w+EOK+xKWzcD95yOoSal
NibLpXyUxnhOWFOYYBLAziMo4JiD2TDh+HJOL477E2AXAKwWhmurUZHy4hp8V5ol
npqZsiKsYtSlcFnaOQ0d1zd85cAyjrQSvFelpl548SdxXSF3NJlL9Xf47FEQZ4sM
BasVvLMV9lcKRxRtg+gl2v6pL8tWN5orA2D3n61ul1gjWXjsn1g/xtU7/1t+mPUz
RNBS3nM9LtSb16lrSn1xB0D6vO4Xz5/SBumygYq90V/e1LSXmL+VtJt3REytaC84
Yk6p+4Mgj4M2AMiDvFVobBqP+gcGuDrWxRBkFeeM4I46ZQNkmwqbrx1WaBBWBjLf
ZXsblCobfMNMk4WitJI8EK4gEwQ5x4h27r6Ttd+yRRTqsxsIb5ACbJtRFWe1h61n
OgdDQIqPlE83+d5szICsBhnxbdsR9w911o1WUH+FBjrMtXxfBk0qFvlR7yNRsRTi
ANrJyCLXUmJ1ZbTqgYAg71fH4mYcNvCTTWrYPsmJsHXEEEpxbhbVbfwgkkmUCOw3
9xqSRtHOYLzzKF7VFldFi4+6jO2fLbM67PuBc34TxDrH2zAqiQr2Sc5zIxqtYF6t
lhm9SYs8x2BvmB51JHohgHMbiSKskGUmkAwFajFic2eLXpf8MmQOHgvzB+DquO2N
J92yOqP8nbymNdxpK6dJERL4eJmcCYkWilc0J0FSJWd6kddfSxmRagTcdPB91zow
Ime0aq+zXurLV/T/YUsu7ncmwwHO5J/0K45IpWV2nUdK61OOJaTkYj5FE/SNEAPS
nxIRhPbnaRKaCcIkyhjfVqmWSr8VTCvjiu7E61vO2YG51n+v8XJ45fEDOrI9TzTg
Z/NmjZ0I6OQGRt5NjOIGl4GKSXH4xLgbI15wZA2ioL/oZ2sYe5SfTAqguJLUTzY6
yrYiRBTMXtkPI0W/DTcP2cSZQJlmeM0+75xD5TD8o4Bb6IVL1HrWBqlJ+HYmr0CP
IidbyJfPkk4UwtgMVgZO6p9yZeVaS7Iqv8MyqcKx8mhq1QstHWYOTHg2sJGJrBSv
Isz2fhYEmZYo0oG7DMC8Czn4L+EuK/iWIpqMPiqjyeZKaTaJjQ/PYOo6s3ZWSB31
wm90/ODDcvYqAi9G1mP2uTkhXAhMJZZQ5sdAq6ALHFdV1EE2Pu6WxOCoI2abs2Ku
1VJMvNclkt2tlTioWLGuYSyMY7b8AajPvqjbeolAInlL854OQ3hnK0/ovDFAKztl
YszsJYOvWX1XYNmmWg5WSCN4rNxzygL+J64rViOBfwkw4DQ4Y4vS1ZfDxu1WBaFm
5KbziTOYohoCsjgG1otJhOqHZXoQngXgHkLkXNSlcJBqWQqanGYb7whRD9Lxlz9O
23FMgA3QusZxozIsszc5gzDrVsr9A+8hQDWloiTkJFXSaQogwD0x1YmKYtCMscid
EIKVGXDvaD1yb9O03xHtgsRAYMH/bcjQ+TsRxveTebnvNTgAgNMH2FCl4iCJNBBP
Trev2sefZN6IIAS9LeOfg2fWLMBcfGEZQN2Hriyh0fla9eAzXnA5ohamkDWjbx/Y
OLkbfehlZBACBOYd81Or4Dqr7ppVYLzN368TGyZcrw4OELCpO6TXYN7imNW6YJz8
1CiF8yboMjcQ1uA2R2GOG12BvO12ZFaHehjssyN3mRUGmtTGZYHoK6C4VDgs98b4
uhCAfFxG2OVkc6emrgNRdpItyf6LT6kPrO5tgn5KyYL0uMbTkoDzYz1qjY2SGwTc
6rBVzrHHcxpKA3mGj28U20xP+StnbhenjRph1k8IkhD5HF5kFvMAeaoz3ptTzsAO
rT2eo3ZJE2lu48FuZgBibLZwLICK3bgRGipWl3xt0dzMOYM+k3urV/we8qK5alYT
opgbnWUpBa6VTmb8QguR1rwNr4sJ/SJvdjrAG0BYYXbAiqymDMhkWJC7INga/vYI
xQ19x4ezLBqRiFeucfSVhiHreXM4AIIOQh3FaVj4z0JxLS5BimKABnJXHJKDoEmh
nd9kHXGxy4Fc4vbqDYYW1cD2o+PBogcSqCGJCedlgCeybM8AmQn33LkWA7gaCm8i
ZYjIxnjg3p3ZiBx9LIw/uhdhSGhmnhfdgxADb/FEAU82lp5rSkpxEQc68Hy7/+3f
ahpFEXIxm5LOSlSK7Zxfp+xAUHg3GDxZQLy2VeCxU8UMrnbiEnzS0nJ4GECM/eK7
5GjH8tSG9HOLq6c2xnXR6j2kfMGWXzP1PYkbuJnx2FEPanRZ4uUIkqdpqlH4A2o7
IpGXN4J5q0lwqqw8Qfk2Qk3FMU6mysnUApngdD2OuyA77d9LAF6fkkQRDfE6NInL
1M/RUnqJ+AvI5SdgfMEOzQuANANJFM4p4c8DD+muB8oyMimEbg65LT8xTxDpe1+/
NfXOaf5MnoeiKs1A18TGO9R1VWV/VHbhaFzMR3v4vy6DDAgWnp5KKgJ84DxA5Fpj
KJitehDyfsAPH5TO50RQKfl1bYIBBCsrf/YaHFS3rP3LdDEA+ezCYBIw4202cmzt
VXJyeabBNO43AqITX2eP1yz16e5GbwKkughvGDTAtnZ+wJIMeC70mUx8I3bvK8Hl
KQlBij0rP+50hLFJmHD+GmVAPKlxf6zttm0GUeEs5OZN1Gr2pAOLagTFLtuWMpF/
JbooYsU4zaeEb1kJ1DkgHRCoBnhKTRjeqSKocEt/OxaTZuAiCgQ0CbeeKhkKuS2Z
Y2Z3JUXrM9DtgEVLhMjMoVlk5wQTPmUgsq4CF0aQkJ5cp5J2O2lSYzxt0KIMq01V
qbDoCecxbTOqeFT549MV0OZWuqAKzLdR5Vxho/xQEkeBe6s4WzS2/ncl+JZOy1xm
a2ovNdGvLIoNql7QpQuIqRrD8hEMqS8Xv0pEdB64pdYc2qvV47ilYcNsEp9TGTHL
QdgN4+QkJdCKV2CjT82qiden84Tg0U2tfgyZGX24qYXxeBw3DH3Z2iC2N19jaDlg
faInevo+72dKw4szaZImqeJ4bHVqOES8hk4/b1OxEyxwYOZE8EA0ucej+VpVY1fQ
NCWecWD71HQ+bZpVqo0dphdrilZinbUEl5/j7/Do26CCrvlVurUdF9s/mJHYCrLa
/zr4YYG6WRxew2JDziUH9vXNXPKtksk7gykjvzywEDERQk69yHg4MdBX+Z5B6bGJ
CKhHX6D48eF50egHph+hQ5zRjsrTzGwZr8/wCoitl6GpUSbwprsILkqPW5bntJmb
2aZBhgfM36mu9FeWRa9uV1sZhsoS697fAPK3oiJnfEOCS3e1lRt75+L61JHE+547
3fhJUCjB7WXGzo0OsCSI9MDu8XS54a4ngZ2b9/hd1LbFyF+JNL2cUed494/4a6v4
9asE/qv8uegj2mvvYodFZ5V3bUoCGxf2Kh1EcvxtUpM/zb5Mn8l/Dk9XKylKgr0v
o4e5a42z9iyZs+fDFMvyyiUTj77kzsME+Ad2LXMUDNm96ze8maVaMN45K/5b8InQ
5jwRWPUCQs9NS676hmP9ZKWHtwAPGC057yxhBtokNLwZCsLP9F5jcDu7NkdoeY9E
krx9SVsBPGnI6Cod/Db4L4MuQGMC2NC0RYqN6t3bNX6YFMFjWKxVrvTZAcl85sXY
UUzEyzUnsTOIGBjzUYnHvF208sig/f5ThbQsDqqIgdmq1hl5LvSMCjDu6CtWYUkc
2yUKNd01nPrQPVQ6tPHEfDi0PVg1DjGPnNas+JHzUW/YPTfqoudD4UtVJWF+mWsf
ae8gTvPtgb3v/o2c6QJ0kAL4q7TZlarO/w/1mTUX6nTAmQL7PMj7pRVyqoEZAhAs
O2CVZ6nCZCJzWBM+nJ417vvamM+EhGQkk2J5l6fgUnsD7aMLWkfCwBFebITZ8Iup
XdlXXKPGIa6/p84s4Y0voYG7lIhMw7prjTrM3xcwmUaSyBfPGLz7LSYEhhYCkVUy
y1L/xQOlU6J+Yc2dTAJwvJjI/d7ZEFpBZMegHQl1H6Zjcq0Ldv2RXNj6IkjE27J1
p4LSdO3ye/0jDTeJlXl4QouXf+nrUv3m8un+dxsB6k4sRwkpT8rX3hjt4D/2OJT8
OxZZ0U7nCQRRVd1CFjgQxLQorBV/W7A38Maw7c3LjDm3JRQr9f8JmQH9IJuU4hvq
Lgpdyq3APvxIAmhXy+SkIDpxxUL0SzJFA+KzAQgzM3TRBsRlLsLGZhve/QydRThO
xZLFA/W7kqwc82BxIRMQrthd2Xw3grKf27KB78HqeQwcrLzQpEfdRaxIHaGOHD3b
s/e7Voqo+PfsTj3QKjXM5ch51PI52RyrZD5n2cIn/7Zh8KRO3ex40JdABeHPiBB+
JE9pk79+1kMFtsRo0WoYH5HusgcvH3kv+QAnOn0xmZDoSK1/atTN2anhCbpSFurj
OyjHAgN6r8zQUEk1eXq1RhBrPpSn0guJdk5bZkUHAUwsI4TUGdD+TfAhn48GT04i
+ViyHGWfFrksORo0LgN5gm3f6c/cML2i3wRWnaD8lN9YbEi0tb5JUM8B0oKtEWhC
31jDCP8E0J+tS+zQiYAHuQI+2Uk1996EhgCP6VSVDtN0lXRmItKIk7BO74wynraD
EU+CVoHXbOXM9HscpWJjmQSgYGfJO6aqqTvExOCWjMkzbxeegXOY7bs1k0Y5fti0
NEdLy5Jdv6Fd019XQ50MOcIF2jvThikjc1rqHf+qxJhbMeXfJTGpImyk1ZfvYdrI
6Ae2kFEH9Crhz1wQi/W0ndUJAxDaRPur1o1mCKVk6vOi0Z/GakiXAyXC/7Fkyqu4
5uMLKzE1+H1FF4axsUrdnFOcuTNZYbkmATkvonq1grudmQB8ocLV5xhUhQefbPeS
8BNha7wAdNFOFo40D6Q7d2vO1wJXlAVVHe/qkNNgjCPYkbN/xUgqz0SUjKHaHbGU
ewIDCJ3cAolYkOxfgGoW5L/0s5o0yQK/Tjkv9N+P9LqwFH01K/eFRnP6CVZ5Q0sU
RnlNxDP0GJoW8rV2BY5uaM5MjVGmfsYIoGzAHMHCObpavNWCfZN3VWk/bE86L5vQ
4gGiBcpRQXfe/JEPuvgyBYwmmccEv3YaD2X+j/oXV+sst7S90PteBzRSWswBHISc
sose+WW9o8L+jx87tHEOFIo9AXC6Ad4r/Q7riu456UZAljodDUiTMAja/8F4W0XB
tZzH9aZmLtck8IA1rIeRGgcfBxmTSdpD5LzF+sgEgHAWDdr5vXybl+GRJB/5U/QF
IZULP8/h/jQYNMwIIankgZ6LP/krHQyqr/HvtmO4jTR2pCM7eNIjyKF+0XmGO1Go
Tl5F6XerC8o8u/Y1D3+ttcJMPswc71ZEWRNeVQ+34QYahRoQmDIRetvyHjcOn4UT
lss4jfaTpLm7RGOcyGU/BzR0tTQ3Q5bT0v8dCQLYADkyY73oXc4rR+7teg7udkWi
+3FeI0D3Y2iux4quFvoHj518OJJwOaB3N1EH8r/mQUySoEfR2yXTSwbqfVUUGhvQ
U+WrpTxvgAkl3ngZHTjGe7nbAlCep0NJlc0j1azxMENrbcfv/1YpDQ+guc2TQIHg
jbU5aLppB4fw5C1eNTKF+3gjgd0kOMMCE/SLd+fZhSsbk08dPvTv5ZFFOqFBoQnJ
EjgQQKTGDD1nlIc06hKzARalk6OTqJin4hBMJtzggefpBZOWjZ30cY0HE8P3R31K
/ptqACYiTdcfSwkRap0p3vcfJ4ePxzUTKGIEs9UJDFkiFa4IzVmq85I9ftKGVLQX
Zzz4oX19usYDG3xfQxiUufXowxafHc5vfwcaCtk5OAo/wlVjuv7bxj+eLh1E/7t9
sltRmw5hoiV8YdwTnDWaClf3eSlnhOV9A+1/2R6SF66EF6fN34ld7cgBnJK1vtnM
zzQudgThnrAJYLWEC7mBY5EK975aKjTjznL/ewR8JHTBdZO+des6XYhydGZfA77e
3ltt/wGOKyVbM3anvS5mpZAmajoVopZCIQkrG9RL+6MLdq+3NL2mqnShdHdCC+EF
fMLfY8o7WHLm7Mmm3i14itYuZsGZ34NCqGISvuDQJUH8D2SF1oTF6jsq5DMefuDy
JRv4GNsZ/k817AFj9Xdy5txGwR0fb0QKX8xT5pAMoyijg5G2ogmuWUIiEuO/rxjl
aZ8g6l09ijovkvFTKDlF2PKagwDNQ3iEy22Wi9ycAxRaV3s6Ms6HdGjpsWb5078D
7ds8fNtZNzM3xTdHrOK05rO9fLrLo9vQXFbveTSxLFA6zfJnfrddg7yV9oR0grh8
YKXAnOagV2U1y+iC4cYaxoAIkaMbdbiOBHomBvrLaTj8Ga3X8hiJb0BjAmno2Db/
J/mkACl0AHDa2ZIAwsfA1mxXcZTBm3u6+zKhzA6eBZN6G6+haAVh6DJDYLFaLfG2
WYw/R5/8OtdN76UfYr8iUzTUu+I/qfc0pv4ps8fhwgRTNN1SC3uYD8FGPdozxoeZ
A3w6EVdfRK8xuC6c0L0Hy1YPWWbAhgzqRy0iPxxQBlntTlTzt/jE2kMYSCbx3Ity
P7j0iHlaUOSRXMQMBSPNhxtA7vBURxrY0lrNKNhOtQatlRkkuglQMAXfZ0ABMADH
B2RxKNEfh17XADWmwZGdTbTRFlK+Q/2awYfOB5iM79b7C6jOYn6MEuRVj/DkJGg7
oynF2esPu8DhD2qgY+M8DwR48jZhopVVq7sS/cX5DXqnKS9s8df7euTJYqDtWiJQ
WmZIC/NSeiisvfdtnQckIRgZdf/zf3GWFya/NQeCVtRJkcPTQsUlodXF1Onmhus8
wqWrumy2lgR2lvta0c0nqKJ0F/4fSHgk8PWfcUhQzHMvzkmCzqMS+Tipvuu8xa4h
fUILU7HLSOra1YtmKZi1F9kOHHO+ofKAR7199FwA4oysMkYE9AQsFsAXO0DKBOuL
zMTv1wJwwE0jSBq6/gU2BqIs6oWkNpfPCEwIs6sm79Vjtik2KI9CMHNSjtlsuwW8
kVytHMCIvR+nOK/Ghm+wkZ9CWH7G10Z6XfncAyO50lKI4GqXETRfrC18GegFkLRe
kElRojnwoNOf+73wThWJsZFWOWWuemkIU/HHAxlVQlfI7J2V1Bna0+tjLy1WCfxl
Xgkbr6bT0NDIeEHlSSFiuisDZtxbNmsnR6EML1lfI5uT7HfNyFxC/4P3pHsQWrUi
1RGDHaIyKIaOpvuzLRAki6zf1ZShn9pIsDwH71hwBg+DpHfUirvsttFNEm4OXOpd
GeqBIiSO/YTwXaiKZD2LJZYydlM9sBl6/Re7DcpvOvQW+qzhqkRXFU899dXS3BA/
iMF0oHvJx/KqLUhC2qxgtkpte9SQ2zhQxviiKSucsD8VrkPFDBg5eDjIk58uc5p+
VwWRTr+KCfI6rlMmD3tzUtCcilfA46WTtDJLn3chUww3scjied7FHaeauQ7fBxf6
2rw0sYhYMRoPzErP3+5y2cvUVE0kos1kauPkjvHbHNbjcuq8V3N++PxdfvkWUNtU
MeaJvpghRBpV4rzP0FwuquE0PvRkTGV7G0u98BQbEp5148pXdVrGUVIVHkEoSOtt
tNVG5h+LPw4CUL7D4WGmSpCq246yuvvkPX76SYGmpy1f3aWXvCaJ7cefDsgF9vAj
nRe6t2F+3mll7ctpAOTmONuRgFfOT/C4hOq3I5wuph7Ct8seJL+CTyIHxilAyNkc
CuZAV2+Um7pK3XbpuEXlMjBMLw6hhLKjPhdTh2nYJN0vUdwSe56jaHh47PPw4Hfw
cFFDUbATy2SU6CnxEYQqHDo8y2BLpeTf9Ff6fZMlCSBZMAU6fG7dvu2ukp8lvlOR
WEHWB6/7mS4koTW7wtmE78emx1efupRX8IAlZF26zzzoAPmUmPsMHPo0+HYMo6On
uj8MEe8yeuZeUM7AeUH31ccHMffFv1/jcstvT5vVqozuNWfB6YDzWpf6S9BcgiOi
bb0gclHrcogLGQA9KFrKV0RHQ6M9Ms69fyF37XL+gJnzwdYV8rdzgdPhmOeSW46z
6eWXdOdjHEmUsIW+d1b4pDJd046FRVc7NS677yD9mYA4h/mkFa1LZSyEw+PnkBXp
J34I7fAZO3hueC418zEXlFROi4lydfM5JPasgb7Gyvk4AKT2qjFrQRJJ9T0BXNEs
uJ4BS1ih7Igvw5lBg07l1uN7/sK6WmvS726JndfEyNFFfOi0vlTXnCtX/MR+qI5+
E7+ffttlVhjESfDm7IjyX4treqkwv/xVp5DgQDhBJzXBxMl7vCc+BbhzZ8fVaGWk
DW2q7VtIDGiHDcaZ74a7iby54kN2N3GED2gBBjSE7YtkteTWrpZ/yOjgDEVEdwd/
A3RILabF80pjGhyLjF9zXu+3Ev0XS0DnBkdpoOI4sqvRdVzUlN6GH8IK64L+Ar99
VQ21hSVxq+ya/qcnPO4ALaXmC6luqiGxjRy/wRj4nzvhLqoW3PDgGSXbpMxqhZWn
0/sRcXMXzlOds6rmpITjmfaHV51AA/pDJPn7ltq1qIVZbuSZ9nH/VKyUsIrqjEvr
GHZhCrbL2ii3UO0vBluNGgyk6P8pi8Qg7D6F+WKswsRv1OoFcQRLkfV5y95T3oUp
WfHTpWjHsHmNQH6SolkzjbjVmIo3Z7Z+pgWmw8ct/IC4JYX/G1e4eoq0neme1oCp
h7LIRBORwrN4vrQUDl2UwO+xrrqZmLT4OwHyHgPXSXKVFtQMMaC1plOC824VD4/l
1darYF7rHZKiJThi/mE8zFRI4c1XprGNDa7HM7P/ggXA37qZ31S4MdJxpMKUtBza
zUNzbHf1UZ9DS0VXQjnOBJmzyYozTjKK42xNx51fxYEjnjD1gJ2ycJaRxa7b7G4Z
rft/8XweuZWCAlX7rLtBlp4ELS6OwiXTRXmn0ZaqZfQcuyrE8ACLd9aUc2ynvTBo
WNKB0uNl5SN+frkrPDhoMW2UW3CrVnBSqmPCIlDaLf/i54SUpbMWkc7UAXaXdgQ2
tj0gnTyz5PUi1ciiZ+2OQZecZ7nb5X32MJEC4CQIjzu79k0N+nxFFZS/c/8Z5Ph5
3DkBOxMQRhdV+zK3F4ZqxaK5po6BTnNbWtIgziyu1QtPKAUTosw3kJOZ9MSFdkVG
8yMLGc0BlNurnunWCryiPpend7FsXLC5Uy7D3blLFhHsh9UZmQKG7dr6WW8DvhbM
OjAEfk4DjkxBYiZ2fdwOGRaPYhU9Vo847cw3jCTAO3YyUKnMvxcqLhyEwiB0iCw9
da/5FTFGptIWQf4lcs2stosvpCm7SmbKsbF9FUXgFbZJaR0JD9pNDGenqdPeBqF1
Jn2GmwftkGilnVl6seOgsgXdlvYmO8LZwBjog2AYy/rUwXL+czV5OUBiDVcLyzcp
4H5eUSwV07MY3yGN/AYqJBJ6LB8D6kh+0j+HucGQLx14CwVS/pJXlzcOhLvWRCX8
Wu1Fqsw0WZHAkJQl13rlPJ22aaIt4pNZ65bc0ld0m6bxSjY186G3zhn3QBgFUcaT
VIcZBaGDlhi8kPXInKkqqxw4h/Jco7s9GOMVc+gLfh92ewG+ty3o5JzcC9UEMjWO
1VAXibO1VGOEagr3OWd7WSGqigYaYbYuh7qm4zgSK13utMQlKhJoVCAWPSodr92v
D/VSa4vq2jU3+ouw/l4VmouPWjFxQpApRxtsiBc23omrTCo7/N7VPyPpyV9lxGMJ
A7KJiU8+XBj85CEwPbyiZOQUvJaLW3fcalh4YJ76mdodoUGGKrwklajlOUnkpGW4
3RyoRUcWxRHOgl83ph0Z1KiwYIg3OS1Z2oncQripYrQIg+0CABNAiKNnRnNYlIQT
vUTEw8aAyeuYkfLi+HRJiO7IYzGVIqRNzNvG8OIfnpbmPwX7Tj+kUpoBrID2xypx
ZLwY/kStNT2Q+Ndx6PCaL/FQu6wmBC11pGahi64m80O+RPYKo2+aI0HLAkK5uY99
XzGg+72ELoFp3WqWJnOUEVDyaKXByivz6zsWVtCuUAdwYm12fpe4XRvMF7UIzB5r
1evtKuKYMzpQok4gWCut2VuturpYCvxAVtHIjbXC/FVc7yPNsDgbONjSum1LbcDF
ZlIJvMJ+IkweF8lRCsmocjbeo5cHmHviWIDqILB2D0Bo4lNN1Bg85+ykQ/V96lRQ
Wdmvalo5E6Crr59hTvLkUQt2JQEnBofeYCRYEJTCaOf1vB7eJKMaWwRfGv8LQxKG
C/DV8KPdtlIeQhVC99CJ3F0JnyvtM7fge1Lm94wTlA4L+Qgg/az3kVBTK2ywpwzI
ka0N+6xE8fke2hi+9aXHPvjilSvSgasuZUC6y4w5bP5pkQzN+xQnwa3Gya0i9DN0
Y+KS8RJe7gpdXcoHdj4O8U1bhr1Ct6XnZbV1pfzIQua6MRE/aaa1ToEOg4OVoaaH
1/fwf964J8hwZJJNmNr6Pvkzs13bfLcc7S32z1OlRmLR0dbRuS7zVcv0VHvFeDCR
Is2MnUmDhpYW3lzkKiTYluOP98yQ+EknNrVJgljThvTQ9ggpWYcOoT3Lc/MJnZTO
sGMrY9MBtags8fmy3aEqen4S8eYc1OCNbSs/0zcVlSNE7W5/0Ps7etz9yvqrOFUq
kWFaLAr8BDDxYhYjh/aVd3Z6FRdALZBv22A7wwmDhHH+bOq+5SdfxVHHz59J42JS
0VRbmkNYhEGPkgT6cL412QDMXimtxBknwiNuO45yH0h41yqJOBW+2SIdrfDtT65A
N0jKdndkZfUaefnoSAea2lx+Lc2xDn7iNXJtUBZ2IPmBj+hspos1odoCVnWa/HaP
53wJ3bdMmBA9qO0z3A4PgVRPDzmvFa8VcSfSzz9kQYgftPR4HMLmd4/KU0r4jYe5
GKmR583pvcjUdjctsJSmFFQzzGwp45NSa4MRSEHfguzf+XDulgDRsemDuo5ApS4j
Bd62IpKPqYPVGg4QsMDmaQDHS/67Oab9yHh5pF2kZSoOiwEdLzFoLap7m81gIX7c
CpEOvgO/dJb5Bi2UuXC6G/kY7eHFfaN2BR1w0+c5QrH+ARo6BBJ5CjrsNU5Hsce7
1r3Nuf0mTf9BLeRT2vzhM+wA2dpiMFTskmpifYuLjt1TN33WWQA2oyI32kMdACLr
/IOzFx0MmdqjMbDW5w46TlSaV5woEBehE6GcMwbHtlNFF90jFoylaGilB5c0DMB8
rO/VC61UB+wgjNSNZ1rgjibxT7VAT6dyl5xKPPV85s8T4rODjMQnyzTNJ9vEXIeS
y8ScuW68NLr8gt261QbtbdnfAXN0iYXve2JVO1YyPQmTRHTH2enJXYYBFnzID9l+
l8QGB1jfTyqrPq4HjLOp1UE0uTEokqv88JWDnxdU8LKqnh6yAzScfYSxCy0d3az4
FW3ucU14Vb0EuaCDLTKwzzxXuBMn59JDj5RuvtPi7q0y3pLG2fFWiXtdRo/66BKB
9PBePYGbRjIkW1Y/X63iA8ypGiWqoCuTlUazmWGjDAuhzN9ki8/llZuk3dtLRD0M
cauBNncHV+LyVS2G91MRVfYjqBDcWfZf2sAd+3VOrcMw+v+cpSF7t5NQrUtDMtLH
AgLFmcDN23BVnvM6noChEbO89v+kWbIc63jUGqed/r45cpMRP0qfvXv2Td7GeXHx
U/DTcSNVaGIPWcDd2eiUCAboHMVjcmhlLD3ZiDapUbG+j/oFLMUMIAsU+E7TfbLC
d6eaQSiE6VUGVFl5jD5I+huOeFKA2KOwLRu6MHkjzmuvdU5r3G51XHIOjtP93dH2
macHVJv8H6neIu8XSyyQTnPH9S5zki0bSHDqIX613rgGEwDi0vGPCYN+5RJ/EnNK
i3Qkv9JFQYooMEI0nN7gM+MGGxc1Atr6QlsIURlSPLgkrc9hrWlzDohXepCoW5O2
uiujp/er8s8RF62LiWHhooJQ8zsjmgsL2RutnAxZfLriIdo6zuWu9thivsVNqmui
vkQ2v7G2/jn6YwY9wfqO5duayhq81gBpXcsXo3sMWpLBaRdESkzIs5hZ0aMZsQXT
UBYBty66PQQ/Sjej/rgitPuJWeFH8MSBhjyq1hu2MNXVzo4UXcvAEmo3BoxTH+sl
2qWXF7hZCdAGFpg3Ps8rBDtvOAUMQEkKmm+3kXZwyq09ftkoSeEJgccKiz9Oz6oa
zIQs+BgoiepeyixUf1yBYS5FTaToy4APla6O1W4qMg/wWCpMKeGtilKm85chvJkE
DFutnUIl0Hs2cvuFd0L0Bto9p2zwFn9e0bZq826Wep9SudCkRfHFl9CSMJ1qgnKQ
BFqjZwxb8VCmoc6GUQZqQ/gEf+4Jf2OZwU/BY3lKGJi5aLLPRfcnPIQ2Z1qfS+dN
wmzJjsg3rLUVp2scBqm+efyNkYsNbzxQ12fWfPZMDec5kb18sHhvSQzz4ry4qLXe
VxCkjcS8v6PIAAgsXEOblrs7F3iR6EGRL9lcdPqCdTOu2z/oKfhoXN4I0QR6Vf3L
gmo694fMoXM/dQ24nV263FzTT99z/N9qQSo+pF8Ixx2MY1KPAkAVYleGzRdLUd3f
hPM7mo2WULQTKy1NnJgjx+WaAJNH2ZvTP3xZYFbC06dGsDs9VA0Z1BTpFYCdWkWk
bt7meFm0cb6LQZ3aDHsgkFa34WthpMiXkK9Sny4OcAtrZ+cw7OqvGcebD/yzKlI6
1Och12qZwrbYJ9An0NfnKinFeefBIYFPKB+SbXovM5fDiTBOC8LCeztuLiai3XKf
l1NGpbK3XGAyNvse1CTj4xpfyEihfwo2KY5z8AV+ykPqX2suDW/D8OTy1g0UNE9r
l8W0aV+rVrecaX6MPldUP/oYEu8O1mJoA11DxiLhOmnhDpvRCeUBbj5/EcyJYCXJ
jQPH5lxvfZKzj1TIz/GH+2uLbaSxAb9+fqA2h4miqn+RRamw7K5KdsqOAJV9PnX+
Wk18t8ox+uHLiViwaei//yBCASUJGiXn0aRNjqql8CaMWyqZpwT2B9FSwNI+ozfZ
kvJoooFsDGvNue25hgJN0tccYssXZomQ1xCYMNTRI26cH5MsyVJaT/NpeTETuK5c
P4iyMyg+IV/Arw6fm2agdUt53oYSLtLouznLnkQYZk6dp7gNC18zlIsoOu0KQKVM
dbJqvVML2zpvsnr8LfItHdKTmdSdFIPk4pdPNqqcg8siGpQfc9z1e6A7BziB0UYC
aotRg7MXncTI+DIwsd+KAv6uKl+kI8kKPVV07i92V7mpxXlcN4jeCKw3O4Clb2vK
uG+kOvpfytCA9+n2mV/HTS+cg0FhPyZqRwEueckdLQaN9tkJPLVJZ4vryVW2e8j1
AhsM59GcwmWcjIkJ4oSVcgTOwhhzyXbnHsUM3YtAw/fXd/HgLUlXW5qREhc4c1Kf
j4ECgfy0+Vw2Ly2Wjdi77shC+UhG+1GW56xNV18Oc9BPujjCrPERD37C8no5qRVN
oPOLQdF1BgpCPfrvdPbESjjrV5S4R49cbiyMblD50Pu5DtIu0oQ9gFws4wyly9LH
oUcS2eqQwCyVolYTabp+bKcV6keDp3pZngwL2dnKd8KKaF90UoOKsgODwmG91wOA
vfIkiW3ScSKdbqzWMkJrnLE4eqSlYt9MvAqvQRhntwVOwTUtcLn2izpEu7J/PWtJ
bCA/DzeHwiOUUypnKcai4Ph8nxWWlxdvE92g/ouAlYpboVdlUE1QNGVZl7St4D/e
dfD2AKSv+OYN1fS7cffR6Fb5lFHXokT9LOc/Gp82oy4YY+Sv9MAe8VY0YFZfloLg
IHnAehOkSw5oPYpYxA4wNED1oN02nQgKMg59jXw7SMHxOZabDe7azs8TGj4WL8uw
BrW0Ig2QC5vIoUI6I1j002FJuCXH+4ttRCyKolK2HRvBFP5k3nGMb6nhou/vlwPq
rKosbjhbDpTljx0og0QmQaQSZ+Bsd0W+BXbg1kxUpaftKtffV8Nbgb0H6eh6Rdp9
DZblkRl7ahk4w/3FjvIYMUam3d+DlMjrIQ+ka5iPMAVuNEj64GA5lxnedPfopFES
b3+YTZaypFwIkMePQeDccKVfvLqn+d0VGoKvGYppRb36k8X4fkInrDQ6tYMJjp3G
C1PaAmU+z32L+myTWp02WtzvBV9jTSBdJoaikwFqWjJzN/AJ6DhayLysUDN1W8aw
zjbkuyfIlgES8IFXDVynMAbAbwR8jOlxydWQtex2Z0+9MhUhPwkKmaYJKLZgQHoj
yyfo9WM4gwFk3ZYo/QvX0zH+sEqkNojhe8pgp5+hvS+0msifGhERUaCTGw9Q9m9x
u3nUNvWtQpvGyvlJruq2w31xZBYdSEdgN0q+PRWaatKzcjznkrGIdIsJis91jpwY
pBu4dGJtIa5DpQYYKLXeW780tBAUCZncly3xWiGmASUO+ZQWeuFnNnBpkbO+3T48
mDo8sV3yvR1+ZxUSlJq4bjrrrQfqN1ztabB8UOHprg/SCNSVA4ah1AdQaMURTohk
fZGMiKZlZ4q1/W2EQy4dvNWqVHEuQyQqpLEKtsl5brERa7OEJW5MB4+wUVrQnWJ0
iNz2vfSZ3hISg5z31J6Ehi5G2NkiFwz6kpVZV32Bi8jtSR/PkHc6oNQRVfGcko8M
RM1xamjWPdMC3SYaGg0vnAprdJmyPD1NpVteSSXed5KLnwODC4aP1/nKTGDrQru4
aC6Bh/3ixloEBtKNJE4u+djFT0m9X3Jo4P3sIKddAG+d3EZYUVzDJeb2TINuK/Tx
lCu5cDoBUBeZJ8sUFdfanQfBQ3pkfNCiJibcicwQ0dJYlpIN3ubKgpq0vuESyfJH
9ffYu7x+oE8K0Ubevr8GSRPkMM48B9QVjx+u+sltaupPIKXLKFp4RMeQP8xNDN+N
miLFA25x5e5Q8R9K26ixePvFRuPLenzeRYaiv5bO5yaF7YYwdLQ0P5u51fhZiZGJ
ASHkdsD7QqYPaGqT5LzF0Kfiz+VPxepSDYX4qC6cJ3dk+NZuJ0hyKV1Gzm1wzoe9
ztZG84EMbwLZg9wO4TjefOuwh7TKo3kW5v8yce/tk9BuWmiyB31ZbkyNtQBPsAQo
+ptxcoqcDawoqRh/OZwzjSqc2IiWqCs32YClYcZAaR8BQwaeiccvQkV2SMtJE1KV
RlLFzkel9zB/Q7BMkWU96mLH2ZGv2EcO48RaJ4wbJuKGfNY1Ccj6D7yHwqKIAPU/
x9PbA78vnja07W3tMsIJPv6L6XitQwz9j10GfDSfnOUGTxB1LAFd0Jvou6qmIiop
LyexIh+lXiQP75f8Zxm7K6BYlvP+WsqMyALuH2Y8hF8WgQJFG+gUmef+9A6QUEnB
mFmUE3FzVAV4y9DgMvzUja84DpRDVElvkmZuniyoxP/0nGMOMR8njkXLSs5TQ3PK
3j4H1TMmEYwCgSJihqxOsKuPueUOMIyLUgFDuBXYPoLIBfI1vs6i0rTQk8Zj0rIg
MA7ZKI9MBiQYhFmOiM0CeC4R4j9vooBo8tMY6mquiBupXFdIuZSc9VmiE4kRj/qJ
JKcWt8jBGw5TWGh2HRN/i9N9a1dFTvQ0cSS1N+P2BcWjKz8sZI0Z2eHoOZZmlSDD
ChnPtqyGhw08uBBx0g/Rv4jmrappHgUarYHhj/FGDtiaEmQ82tG701yEZmhN3bfW
RVCtoHR2VdN4G32+ntWHueH99AVKPUGkSqKMj+2/lRwtKO+vF1ppH/2Ydcu2KIgS
dJPlnQ3r868TZMnDAB/aKtA7HkDlgpJt/JX18DXJ4B8seQv37ecjiMyvvlDefi/k
lbR9Dx62liaC7Zer+s457vc1bODP3tgduoUoQ3aj33LwEucVRNK+g6uKcu4KFDrN
6rY0qJ0zIByXiiWv3IM6NOWUsOjRYbcA1R0ep1ospW3RL2NyJTYKL62nfItVlNuM
lyZbW8ixCY9jR9gMsdp2ZZEsDBvs7N+jqweTsAXQ5SsjLMqOXXy7CPeesSptFX1D
QbPkh4UZ6rXPS5yjtWrTTuMxqjpbdEwqgIsgVjYnu7EGaLPAr4aSywKE/WRYANO0
lQRdTNlVkvInUyfb9rO8JhS6bdKOoUBhv4Hh21GcbWjV2dwRj9kGKsCKJZOH3bgr
PMf+gXtP/+tNG3JS2GRwZt6nUbebWbU70pwtHtZERlsUqey4iWogisB+KYbctrak
dIjLjdcgatmAZKbkwc4k+snLxg5FlsqZGvm+zVVRSxAi0EjhQ74rScCFn3qnpEcr
ScIZMvSX1tKWh+PaKM03XIhXLfNHtdCOcjKB6FkkcWoxshsu++7HCg64k+KgcbHJ
6x60a2fqGvU09aL6r//StSKJaZr4pKu3zA3l8kUjZKmcDSOpgfex5bBQESQHU4nl
xVbEsTRWEVynGsnEsTWuq8ShNtX5gwJpE3IhMC4dXt4egWSY45ZjViE/tbEaC3B4
kc6MM1NloEexbIJZjKbZMP/HmcnMMaVCdydt7H81lLLiNm6RubUuZ3YLZSh6n3rH
cOEHpG+21koy8nLjtYg/Juzdc8+x6DhmeQ4hZLqlReEqvRpP5F1+uCY5KTs/teIg
/rUHXRJc5D6NsyKoy9BMoOHP0/8tTWvKFNBJIIjDkaK9kG2u28rpjREsG/osEE64
VROM0EICtjDCd0vl3o7FEt1zjsj2Palg2TXxnvECa9kacEAxAObgF7MuzvSvFDSD
T50+L1MS3Zn+au5S6jR6l/RppxnKL7BUxERuMaqU3vgWhvEwFkuMEyKB5AW8G3dv
G58Zi5gs3HUHWKkP2fnygqa0pf88BW51oo53vBmQojzJsm99I5LhirtEb28x1g68
aCAbcqtM/ducK0xj7mvmHwf4HYSh9HNsSOGwGqzt+CsN//zMyAVRtBgwDS5vU4OY
gl6M4+sqdo7JaQ4pNCdv5wr7NGBIpZ93W9BY7FN7q2zE+dDtUmpXiuvd+8lCGu01
e7fwlu0F37SoyRTeEpRYtX5oh4TN4qDwKJuzZHZRDa4W3uqYwZOvnRG2D472q3ll
KQnk7qzd+zeggkgmSBbZgsSVYbyzql+Lv/74QFiTW6GZpvXXPGYMJwmIFF4aTJsw
6MBFR9VISg5ojlATrSOK1YRgnciR3RnwyiXmHIRHXOmx9XZ+VP4G3m3T6oQaAUkr
5K2t5hiZzLRFHjN5B3bsOidaEKpGc3RzQJbfuoad4um1SippEc1+XZspIxevB9Sl
x1vaJS1ndu24hMHTun9mgY3JXx3XnfHjLqAiGVTHk3abbJCPcmbHdbfLEqQeoGRD
e9zKBp89ivXFNdgtC2pZNNrOMX0ThTKH02PsWeiiglVRjRajuBUJJDqbKAE7dx/F
oe69XnPguY4DRQcbm+nLxecXZRWqBOzVlw4BjFJeUcLZ9ne2xlAUKFWFCqdjYPd1
0zwtrARd4MpK5s6s1eoVdc2YPTAuXPnFmpZNkRdRKkcVV0PdK7OJKDxeayX5s/1+
R12xrXCO64l6v6G5/y0oAtXvq1fKPyzvH5wvlIyPLBtcwlk83fQl5wjwl7YfGXty
aT4cCaiVuqNpunijdTVPqbiLfdfkVfp+UxcELHacDHi8xTTb+fZoWHh9AwFjQnky
HlUQ2RyH/CQ6OxIKyDRUh+RoSbjBWf6TCqojlYhEFY+OqlAOJtC2y2+cOdKxdMYH
EKpV75ALv8eUR17pCoG3WJigZZxfB7Hpavi6va4q7DK5+f2rIAX3Bae3SFkoJXwd
AEEN1mhALYUFd46rrSnn/01jYccq+ycZfIimz6Bi37YFDBVRznEdyRXkI2sx4Y6d
i83u0DIX0JUdfjoLKcwobMLIphUrBO3LlALE7r0l+YzoWGC45lcqi1Jw5e10lilI
xLfWNZ6BTfKrHt6/U564+/AvTIIqnY2iXjQs1rEtp2r7M/zWLY3y60FwkDWoIw8u
XUgnnjph9c9hE5N4JxxJEfXtKpcl/ePyZM9Ndis6KYGHTJ8VxH6DUQz4+wgluKdn
TcsLBrrdv988FgLOMS8pZ5Mub4OKbmUF+HxUHt9cYXCBQC+SkwGSjRixhZoqhMCM
9Ck5yd7kLmtRgS0wIzMCvg6mVwqI026Gkex6Tyk48lGkM0ygKTGdB0ZkqDnIsn6Q
GONNJNySQiEgr+M8J1c/CtTFrI/KbDFGOXjhvz6DGS9Bur0qC+vMk5llsJnXPw7Y
rvxDkyuf7vNLU/lUi4Wbf6JjqKPVvmCOvgCJ0dmGPaCenVDN7EtgNfmw0Qwq7V3F
BuUirbsLWaLtGI2G1hbmV5eNRKmdbHVE1nk1YVZLKIzeueeFbGSQFApZDhPuyG/s
J0eVYlNPTpCcCfgcnHLiCmPHSmwciXwmXTUdYSfKTTl+f6kAt8YUdWF9jsX9DpNx
eZ3fSM8+gw5e7axWHJV4r49bNd/62/+RFfG2C2wwXsTksKXRz/IIFhUdexFEiQIK
cpQQ7ZQt/b/mJPVF25J6AqZ2SS3QcoVKbZ76XmYqYQW4HbxzkLjY5o6l+gh9M7+H
145soQXANDDsoFm+xJGA7ZZ0DroeyjU7e32Fy2v7ApM1K+u7m30gnTMOh/MOU63I
PX4Ofbbkyv5dVcJVDtZOBlyKcmZfC2FIsKuTGzyJAMADkld6C/PhWrCLis3NQhnN
WUfEzRPAF2JKxeh3tSyoJ+kBW4k0W/jQe3HDkF9lazv1eV2sft7uO/IoPG/eE0tY
qhxXlKiyw2Z5oW/mswlsd7ghpoSFAe0WQz5tUxie95zCJ1lUQZqAkbDIhTmg1etK
RO62QgfkEygs3E1yQ36+L9yZ9W8B2iGft5PCAZ21cIfluh4zzbSq/jcmY32IYOMk
ZBx/JVSUQRtDRJ7vp7I9g0RYfl7Y4ledvKtSDdVorDb1WH/eJ8/V1/WURVo68L21
93Ldb2ZqXzEKGCqwXv0+KJmmJs1twsl8o1ZPDvEM0R4hghJmSZhqEwVk4BmGXCtl
GQVZFbjBCob0JCO03DNejZYEp029MuNXa5sxzoBH9h+pG1JrdxRdz+ppxX3A/ha/
Am8qFNoc3BrNy4lq0bND1i4TZ15/cAEhmfbCkPeDGSRCYn5lI6EVxW4CE/W/LRkB
LklIlFr2JuzvbRQWgUSm8RIV6+2d5smHn0EvoRvCbOo9UyHwsCdIv5uDV11R/VKW
1DwOdpZQ8ENX0LuJMOWKOYgEtu18yWqGneToL02Sq9Pt29iJL54btuVABdZAeMYL
EI0ekTxfTAIVUFSo51eNuIU2WQOOqYFYT9vvR70OkhPREwESqB9Ex2LQDxX0TSUW
Hz2G+hBC5HFS13kL+pHgvKFr+99JCKdpPPcaQ4+82HbU/i89IOpwjsEVjS+WynLB
S28lkobhKDS48qjw+u7a1atCwY648oWmyLUG9sFguPqNWtBwMEI6O/E1iuYKot9/
k8eJRWvCCjinbP/m7u/11eSnd2l9OnQ5iQHglyANtAE/ERhX1TYp9oOKgzyvMohW
CafElyuv81N7u2pcmab3OKPB2wLZydvB/ILu3y54C0MQd6eLcoQ7Yh4PtIOcRC6C
CMWgl5eaf/eiCtwFF/nKBiGUE2S+ot6+dUrGFTReo7bIhPmoGZeyUAah/7tVE5fD
w4WVsMkl37lkSedFAZTZ0vtyko/CYRmo3+rkaOGjy0YCEomlAUvpIwb2YKC8At3u
hnWr17KC/jPw/RloI1dK56LpJuKa3dLgT7ElbDnQIV3XgyS+C/Rkg7Knl5glrVLz
/XV1yNLbCWZ346DETwh1u6REpF0sxF9X+zKCTUjlhF7ANFTFlRq7jGZqmCrLeIp5
DASW/Tijje5c22irNpkfS07L9ppbvdqM+tYBAX9PvfJq9qPa5WrY61Qz45C6Etoo
6he7xBjMyc7oQ9cOHWl051IlrsSDCf3IGB8OuEaPEwWSUwtwxSXV/khix1odNtoF
ZS3XRRjaWC6Gm9zqCxsEN0MU663jT2ORZuLD87MZ4JOwQudGHurm+8YE2BixNP9Q
WnGvJsddnJHKhFZRfOqgoqzEPdsfh+CI9uMkmLyK9+95zqP/Ucxp9zzsM1F029LA
z/7CVN6CRc7ZzRlY8GwZY/o1cLv4WboI8zJzlAWmyTCMu8e+zQXybqoEfk/oq8XJ
UEckzgXr+fty5ODPlcdVfLk+wwrIDppQj9cSn48Q3VUThYdsV0hTnjek1aSfI+eL
R9WoVZvUIQ+ClYyl9fjUL+PXUPOqyCz1euyWv6AMFpRmEV1NRMxaQRAM1aPEnLAy
rwLG0dpavDYCFN5bnVWMjLjJFDWobJbnZVViZnqkeOknXrLqyILR7L6I4USi3WsX
9yLS+OgSceMAM/729aP2f1X7RCGOZ2VBdbf+Q4WQ2kJyxSQ0Pz8niAzKwWoNk2NE
SvCfc4Loio10jN9TPX9KUnfZUFAKOUH7nLn9hCV8gwvxrj3XHpskKM22Ux1Ag7v8
h+U/cACa/0XrCV1lHU3MgvsbB9asgg43U0CBxTnS5qZvNcVAycPXKk7UXH0FVA3X
CamOPeYq81qrEpYr6hFKUhIhpUkpXvvwuFbjmPjlsTHRA83mO4eJQj/TkoQuH/uO
nX03N8O7Egaz8QsncxYg+ouwvLTQJInn4yMSeUSJhz43RvLCv1xA1lueU6A3WcVJ
53caYZHbj2sq3yzKVAnQAWKUcYUFX6tMSm8nsqvO/ALpHcPbXnvOlknBCMq4RngO
3tWfcmp5+FR9TJujDRQsPcu2X4eIEdeIzLiJx3w0yFH69R2fr5k3indhnZT7Fk3q
EY8QbX+PWOXh4m1BpJ2yvBtDsitcYAuifR9Jgyjk4L/SQV9TCut7RRpwbH40uUto
VrbiRy3BCuP9Z6G+xlxQ0dI31dDmpUw6kCWIcil3QZI5gxbIl1GzCrS+aOzdSkhn
RyS5Tp8GrpUA8taUL/qIVfsmvfPs6zJHKqESCcDb8otELFlyn02Sjml4f6IBxSn9
RPCujkr/0NHyVxFKmnLt5NDTMpI1IRiLpQvtIvEndVB2WgIk52J75VCxYJAQ5Gsb
c3+7DuX3m0SmrGbwzRXZHWNsMOuoeyr4MgkOSJcrrpmxd6PYx8I3y5qAEpzrUbtW
IdffDGXM78DvJIG74qc/OTwslmOlSgP35RpSSeKcr2aGuSqCdB3MOBiBryA5OQO1
e1KDOKH5SBz4tWD8MKNLZ44IKnLKrfnVbC3ymfRjccDlqnBq3Zd8m4FOabqT8tbL
Y0Co+yANChJzzgnVXIMoP49Ye5ft5rVSGu6hG2RkjACBo0xA9eAETMndWdIIReg3
0pwYyHyOr8/xg305dUcjpOAu/4gcX4xD20T9RSismlNLiDvcI3r5d0P8GndlO2Ny
Du+4Mk7pUp1Tk5XBnAIBiOhCx2821j2kLLbVrUGeTDRtyiTNL6rZyjHN2H+gP4TU
Wuh6v9ccZ6tehch+MEfN1WYV8DVTl3f4AvF/1t1kWXoVMOX+///vPkplPfWChTv8
cyLKEWHc8egQSKJsRHZSOR1s5CbKD1Qp+xugp0PF1aq6b0Xaxp8rucLdn+IyCu1/
Clse2V17QaeCdVFb/rSkttl9bQmnm1p59DoJfh5aRtqX7PUERxgyYFrx0GC6xA+0
X9jrkiszjMSy2ZYx7XLDDPFLEBH0OfIN2RDTaT7WUzRFhmc3O7C+55voExLUWSUH
0ydvDKrxg+e4Qx6eFFWnZrASdoLxyt8VyggITbsRFXcFEukGvv9gfOhHjfWJ8vh9
T/eK5cucSFs7cuwbOs0Saz/xfz0xhtSCJMSiH5qOACLY3inIhAifav78RRVuJM48
efWr+8MZGa9ke0pSxyi5w1Ct4G4tQEEGFEHyq0rybDY4l6h2/9R6IXB00pBK60/C
o7HNL7VN3bFsN0pz8mnI+YH+2D8mCedDWQNZyw3Gonae1Edg0kAhzN20WMgX2tyB
MkhPlR6M5lD2Sbfprd2v4MX0A9xcli/VQ8ir/UT7YrJ6e9wrPc7Mk8bdALGVpk3L
ULFYeoCpicr+lsg0YheJR3py42dPjIs8ORiTMCoLVvp0pXpm8oXVAx2+aUbPfdCy
2YUW3rAgo3NuJ/aBsoMlg8Qz4OCfU7YgnZvi8fO+GwLYQcx5ijXpaLK8CvLcntaj
Yukng9rvsWgZkld3ciLx3MqwDNHsVZmQpvb6k3AEBWv6ZMSaQr4R9z85FemQQp7v
pgp5G/eiAbVkL3DX7G5x57IAGqVYK/gDhdLCfmRnYGBu0yyKcrReslE+rLt1WUqN
v9L7G0n2uRRhW4NagdR0fWjE6CSjEycQp7GJIh3Vjqr54AwaZhAIDb7nG5DioojY
9dbM5ceK6+qUrPQUmRNT0nRgnB5tBMm3i9fSwjVmIkjZ0W9zXvb4J6AQ2hcBkZzD
NJMNFUvlGi/1NEwom7tKeC0sifLZBdtQZVy5K1ZziBjr5KGCOsUHde25Uc8I6+5F
QHQHL9L8M4TF/4gbFm0YfhL2I6JdNnTrceFg6Nz9AExdBB7/veK8el9hG55upHng
PIAmZdpnFfIchbTM5Fuz3DYWaIJt0pp/OBYsDA0eFiYT92iR5rEHvl90tV9QY+00
zJCSQJpME7eh+MdYA3XInS+8q0YSG9+EE0CFTLBpmLdoLWQRhYe+umiEFg4AgPKP
JA+lalLJjw/y7KgnULSLY5a7QVTn5LlKJMbeLmCklu1lyn0u/q/AT2Ox1Z5+hQTf
MbnkDik/srzNq91X4mGT04heKgmEAPz/AwF1zBCOzgZZVhm8JYDtvquKZH2P6wbK
+B/r0RMBlfH9/2hQqWlXsL5w8y8TydKh0kAp/wcfmRQZ/N2tUxescHp12BXJJRDr
qSQR76FtiCWIpebp8h0K9bOdrFb4OourQYkVDB2fPPJRlzyWo4ls0NdQhjZnaL/K
qsD5fKuOgGAqmMytpQl5pqiEGBuS8LDbZL47I4FhKO5BuVke07HaM+J8BfPiWneP
CQcM0nrUgSg/a3jhYPXKoDYKQgqxEHnrx2ewy+wiMAKEKcEG5I0gKhenc/KAukpH
y5bGCpKmW4LMd7G2asTyuDE/nzEuiPSzpT4n/I2bVtNv+ycuXHjehGVYqPQo8+Jl
kl6sxXHcRqiHvTLzMCdhEYBaLoxmBka+Kei7Z3/yA90iiKm57WwePYse/sl+upcg
1T2dQuK7bfZnWO8d1WxNRGP618qJ+ldprNn3MK9/ERg8MAFzJLk6ni5PG24Bt1nq
Or/tJwZ+PBpkNxY/KGSTWesFdnOOMurP+eMxliT5zTKR66g+tRLebkWOvq9DfzWJ
kW5lLm4qL0dnPBaDKTTw0m+Zd+ZEgW1XxojWplwNaU0s3VAhZ7OCq1N7DKn2c8xe
ossD0lbFCpHRirG1StpCzifs4wQsmnwUkaXqE0pounfGOfgMjOBqDBgWA9hJm5MU
5uD3G3OZMPe7N3hiaWHoTUn7W+YATpUkLhO6PsKWReLMP8mFmBg/zopHU5MRYXL1
3PPo5DCs/bUkHnqv/tNPo1TCjUbtdnySkrGHRZKx8bY/q4KSSOAaK+Hh/7yVNQKL
1uN+YiHRJhRDOYUSUqeLZ3FTkartQk2o48s7qIs9kIqipmw3kv79XSXW8+FY98KL
9n0MYl1otrqluJeRWUGvcLCQvkZSfqHr2X4uf4QsH237i6cYfupS92LF+amGoLL7
BFxKwho90tw7sZ3ljXAKWHSEqpkz/8CynxVhHmz8q3vnuYSDug/SQE2BpOdk1Va6
dlti6zqgGOI9CBAT7cDnHYFh/J/oRdr9SNbTdUdCDPbiU9N0/rf2vqkTSwbU9zDR
9/ZNWXXLDkx/8qo6DlXxVgeQCrj0UJ/7nF+JADPppTSRDCdkFKtq8gW9nvxOgVWW
vgjjA8SjLyHi5g70PC2AZM8SC7QldcEVTYaAnRHIGA2rDgbUgjf2Mw4mgdS4YJ4S
M+KDpXA+bolyzRBl9NmN49sHSETgmmFvou6vXQTh9DKs6hQfN3hgQIGs2e/pK6+w
xxV/2Gt1IC61QEhI8PW1xJBqht+WpnPIi8NP2lFCM0O/SGj0X/KxS8mDkHjVQkou
NXTrqdatla6Y11g+xs9ymxQnAu3U7jD+A9D4zjVaeYFEUl6pgPBKUv034S+6wXT5
9IIK8k4Dims+6EI+CrPG55jv0MzCZGPFTjQd+AMBBC7AUcUhEoXzVmnfQSgT4/Fj
VD2OK7QCraKP78DR7vCOuHD6L70hbAhMiXSQdYgFXaQfGt2WG+bf2pf6A+VEfOAl
uHrXJe+/Il6hqbBtvJkswsTD5AW9e1zNaiXSMpJP3BJw4rFwuIv9oG9YSVgMvhMY
W77BGwo3h1RNBA5ZwAUX2MgokrD/1AtzKOkXpOtxyaBu3OU1jHXuT56qGENBDruj
CrcKq0g6Pi45pZA4j5jc5ht9t3ck0beMjrcqHFOq4o1unc5KlQM2tKa1S7bLC9OR
B+8l026yCtxNtJPzlHzzSPdfhnnto5QLiQm1KiRiFM04naIQAeV3Pv6PTztkzOl+
BqMkxtvA68ln9pAz36hihiOp2kt1+fkpZcdBgn1rEbnTgxAGa2Ejl50m2hiLY4Dt
mwXh6EvSJ5lP1xKOWwEKJZ/mEhUP24aq5CwzgN8X7wodvVpyU8HJP4eh27yJf3zX
kSq2Y7S4baQFJuKRJjd3thEjHCkseZhOQbrs6RiPOb4cwjFAeBSJ61B6oi6If4FO
SrolOP/6oI15Wn2E7Vcf36+4QYpSQHuyXmfCYAT0x7MtFIRg7KZz7DmbcEGekiWO
8FmS3wwegTzD7ktCyf5XUlgdU6nArW0xQgIMxEnY2K0mbr+g3B4nSXlQi8YdBGXI
bp4glK7pmJxl+yDS0Ncakbhb/Za0eE1fjA4JriOCXOhB6pzxYdUchMjej+Y/Ne7i
i7AfCUpl82Mu+MqhRVsQXsyerCj+6gjBWypJU5WOmF3pHuQmlrCciUdO3EmjFcd/
neoiP0sW9Ds5VNvQnsj7WcSCqFYijMT89NKZnv/3QDScGphN196TmlElmVXQx4un
VeC1yP+N0iR9fueVtJuphM7Hj8KHZUOGYq4HaSbtRBc8kc5HEFnNiNoZvELKT7sU
rVpjj3g/wVq+BsrVu4ZB9DN9swspleQB5kUMGfEgaaW/9q8UwYGgvVI9+Ca14Nm5
UrlF+hs1cDEkQRV/q3NQARnslS11FLDGxwuIzmumH57u0oKGpBCxqDZa6kJJoTns
GWVVZAOYuyFcV7htwpfnlt3hfUd3QVGyTRuPtU5GbkeuTeqsmpX3NZT4EstYZu2l
sXq3GUtxpm5/bNTb/vEzdJXG4+hCPWcmsvPOK6M4z0VwqZ8sMqAXkUW2FrByWkcI
o3ANIOJScD6X3kKI2U9GlLicMbna/rmmsEKW1wYSkxQhiub12RHdf9oEro1B90KI
uKM4SCo4LfHfGCNBnmPsWvpvMkvFrAWysSkitLH11mE4daPy6wazdugRc+iqvYi3
0mBcHLw2OCFe3Lg8yw/bVGveX5sBO7Ggt8AMkF2R+aPzEY6Ez2KMawNyizpZN/Lt
xNNkzVTy3DXlcz7RfkepOsdqwTEJyvTyeqmV10HMStYA05DO/w4F8DSNNA8v0E9e
PAheA78pP3lSkoinGwJctZ2BjOeJxbiGI0fpzR8BZ3J/RrAMfy+8L2dnxjU/8F7n
usCQJ2gmBwr1EYbNa+SFV/yybTeEpp7+TGvp3yA7drVlAqRiBGPldB0MttlRop0D
CEIkapihZub3npSDa9vb8UhiZrWUMyhK71zm/miw1/P+dhpprT6W/cfd1ktkJ8u3
7C1X+s7VE8NQT7jMhtywZ/UdFY06NWE6R46qWuC5dFcJOS9Hko5j3FaYMTmQ1/6Z
dxZ0r9o/2S6EmHMU6T8/9UZCU01SCcI0XbTfAOqY7Ws3nHfMEzTaQIaHOrE98VAa
sKBl5UjuSRwgsGc0/bI42fZ0gfdg6yHzfr+jS51r2kYfvPPDdNOHE7svH6xERYjM
mURQhjJDOsevV9VsAvnaE9vT4Z7Us+YkxvVb+69CAIekLtq0u5PTIDjdaxDf+xlO
TkYsbdInMoKOed5aqg2BU9uqWxwj7OXR4TAte5YhuUVc0DqTvB5KYPoJ4VMeUaxJ
O2OTn309TiNu7cnItZjKR+Vb/SWXOBwyyqFfFIF6SH+2FpqaNpGEnoT8+gH7S/+9
4fWM0vsz2/koeDi3HSM5vtq7CyiSToY86GWRn/Df2lZo06H04fjqoGoBBZ3mDBmb
DNQ3SrkT8Qn3oQ5vKXtfDAbhRMpPumypl0jDb21mKgEPaHcXBGCo+ndv7nJpy9fu
6Lm5/pd7y7Glc8rL0pFDSufnlqL8Ar4fN8CLvPbGAXoWTaUirISz8U9eNMsOmk5Z
62HUVW5KixjmBHsYqYYOiLVhy0YkVbUEjY1fJ/YhG/kyomW+IM/PAbMey7EnJEqz
jgPz5nCgVnWLRN2/vvYdfePj+FIa7ENTk4zE+TdjVI1wviaJOj6MGGBrH53vA/EL
naTJMMxVlLPQ3GhOg23JySqhy3PGbcXD6EJpuKwIFzRjY/qfqRgf110tNLY5nX6h
jc/yF5BdC9fgoSbxyGwgg8a2lygxuQK3vyyY7YldqkrWiLXEvL44b8Z0bw/0knzt
vZI+0Nq41UziicJvsDDij45X4Wt6YtW6mVpT0Ps0+67pyokXTsp3dHUOFd5t7r9b
AtmEqnS8QaDTzdA5kXfHYSmWydAad3BYass1cksxNAfhvmN9EI4vexzBZ9vbssmv
djtPJ+diz9dPViNQ/tDKB/H9NOuhcQ3WhR8x+ufM1JuRmEmmOX3FJZxknmUPgDXj
triDFqTONSe8bhIKTc81nx2xUEQTQtFgVfFxvJcEjRL4Dgi0nzhEGbmSnwXMPaza
4tqfP3iRpu8HgB68ltbnoLqbLxTKGuz07vO+8XBehgybT63n9uzaT1lmXMeLfY3Z
GPYybtYWpe+pctoHqLpj9+76oXvYaaQls/SgO2lRC/+gHeIAvW4J8PaYp9zA2T/S
IcdF72R1L93eZ2oOrCieve2g7owIKP+X2NigypGxJ3/3T9YSjTL3t1fpq5IpJr+z
sr4jE2dA7D0Cz1Dr0g2E4VDExZn68QtodLRNEj6j2Bk7IPTaxakf6hUG6f/kcILs
YkL6YfH7zSStq/LGqTN0c/IDJ478GU+nJd6OTDV1SEU5Qy141YA35tXpY9n437Rq
gXMAJLrmdKNC/AtMXBfTDeQJLSTUV2hlVqyNtqorPUB8VFLncQPjRzsLzxchAcnV
BiRsznI4Xm+FG9DMlqibNbcFnC1hW/a4X76tZffw0X18/2sgh0iGFYP7uH99mwFr
O1SEyH+4eYMoCijkPzVHmZST5JIRReP9xKQrwSYQbtekcazXcTceGnG9LW8SJWdy
FyaZ7a+BqN69JhHVw4bobA5Yn6ErmmuP2nB9gvJrpXCGYASaVdJBP785FgFaCfcO
KoEwSz5EI50z5Iu33cUhCubOmoQWW548kHaUwbaEuWdCzZR0dEn94RRwl9vUM8zu
wGCTa/3TUB0UDpjx4eLoYYCLPUfb56po29e8B3BL/SFqoDvkGfOSLtBKptDbCoMq
xuswVxyTS79N36NyLrxjgeo47Tsbpib+g3OlcCOK6DAj4kKVAexrPwiaE8E77VGZ
Df9HUuK0l+FC5xkSkXtiitLhKPYbgscSOdcWGbZ22dEk3nDCjVhnxe/+vOlBMrRt
d9UlGq+C90Ju/Xw9HZeoK+HkeubS3jAAwQ+M0lTD4cakCz26aLl1vYM0NgFzxHSX
wg5rUNF/KrShh6VuwDc+tOVxYJxW/Fp11Qj+dNil8RLstMGZNtc/p+WBRQzdmkJA
j1T41xAgexbmsZP/hrVlyK9eLXC1jNHTmUfGxZRZC8FbN13F9tbwDpvySk0PY0wX
EahV8S30ufFXVow0JQqeIrRfet0hem8xOwMJ4DRTq34fgjpCBWBxmbjXQBgXH0nM
o1plQnM28XyJYA3NF3uIPOS4iOllpkl5NxqdRCtZRls9gQVG3AQaCOgDRJk+BLiQ
ymFWObm5ibb0hBk3Pn/6ApUIALFgMGN78bhlb8kun96UQlky81IbMw9EKhlDG/ss
3yZeo0uu+M7aH+whH2lF9Yqq1tBjMGxf5mNatAVfNgylfLyLUsNf7gPWiK+8H5/g
uFAV1y+W5Ilme4hCUOsaHQFT7Dz/7p+CdxnHCzQ8DE7oFZNj/XIUz93+X480oLZc
peKkJ8nS+tNjJ/MFoKOh+fQQAxhZmMsTwELWfdV5mp3/PlwOQnJc2SH7p2exzYfm
FiBxsNBi/dfll1UqoZv7QZGIkjORXmjWgZfpRIPEvRKAaJEec4u9DFec2ku5SEAe
27pcOAqS+dC9cE+opVv5ny4qJop3QWdsU6gaiwdioFeJbR74zXMYOtY8oOM1Qkn5
VxJqOLsd8rGXAMQ1GleOXDfl3lpvGbDhluk69+K/3PZRbG4rnLCtvjf3i/jitGbz
cLM9Xsjpz9wBAqalxuHVtnP7AzQu1B5Ly8fpcvAGLPQyPSEqCNS+1h2SwHpgZS+6
yO4dlgfhqwYxv025yxSyoSWvSztM3jgN0KNm0c+QB5p79piOaQU1MnFR12mQKEwc
MtyKzipPt6hKb1WuzmbyfNZTXBa9BPkTO25iKAC2o1aD8KM/yqGmErylmhy4GX6e
9RbHV33nFqs51fRZrTo3QU76mAChnSOPAG12LNQbT8DqybQ/XDt8P5mK/afrjVje
jC6g/1wWD47noP5cjWUut6K2B8ML795HfvFfoeNsLLT6mqYHv/mmvbax+wxlQzPA
6esDMZYOB338FEERL+ZUSC54ucccgbjmgm9xXn1ZhqpdgHPWGB/NBONq0qV7IKAL
Xla/pj9F/lrUjbBw0zwETjLLsHaHA0xstflGwVbX/V7ofs7d/Dr/9dnFE6z5NAZ3
hcdPynzfR0mC+yFRLnkIYx3lMkZqg09MSFcZaXuQvGzik5c7INsIXH21wX2ihC9P
HMxyfsvn6+ba3/04dhoZVYnBISw56uDouJ4edbqpWaSq2WPrhRxGqTLajOMn7MxL
fBocH6n3xChN+YUQnMqqV+p4tLQkL4HVP5eoymz9PoOmwdOCf6KLds3tDqHRmW0n
5bl/3Q8KQZi+dqys8dmxJsS2JAwSVA4Cz0VflQfAvPJ6YT+8VcuHbSE3QsmPmphj
9mSkCxK/TJjE4jVf+zWS+0xx18IfC4g9qXDHkL0zDX78Yp44gqD1veMSyamKSLdt
oLhW4UY71ftqrMtD7989xQUMCUbgl4xIQJCh737rKpziefI0Lj5rY4Sb8UZN06lr
ij6gJUR/GFckds2bCzBgnY7Fv7vJ/RluOGockbUkZaB8gAeoJQPIXBDHkAZBpnat
7qUonppD0dMR6hOsSZeX86zWiaXTz+bgRLXgBhxplmfPIW+QA62JyZNWeQyh5vIY
Sbxk6a4iJVEIAl1tQMS0B+Daz4ZxH99fGHEbQsvh2sB4H6RFbyQiiPCUUJDnDXII
dYPBc7Pf2QO89C3BW4PZe+rWaswo2kPpT+M53i4txzCnZij/Zo/Vr8Qbr6Mws1tq
tlROKIW1JbcldEZkHP8w+Xi7YG+ljsvVy6+wN59EuyrCuYn7n4iDqpsPA2KtYfHI
ko18m03TWvDfN6zZ7eK21m+h3RWPsgr4zYIHQVMVyDmh/GHstpBQicW/Rmv8jCB8
/LmmguFtTb0iyIxJVGymXeKLF6dnz2dJaGUl80cd7f0XJVfbUr5+s87GSE/BsH7I
T5FElOfRYYV68HHRsdmxGbBmPLPCO8lZMKAfVA19JYhoVwx6SxTPNVO6rWLmhsHZ
ZAuRR/3naxDgLT1b9vdoXz/pclk9C443ThXVweyeSTDqHcX3QS/GJ79LBzNBTMc/
HqNWNZOBPnxUopBbjaKOho8ehYUBsgDm7CKIC02fzb6a6kBL3tYw156KY5JmuGm5
9f4hUruitVXxfniJO92v/15NQMxip9aKWumhvm3iSx0XhZROJYdEXXHvtW2r7Pol
2FGiXSPPdHVURT7jpZHA1Hqd5ZEhbX3YO3uL/MqYqwV/Cka7dawIHY//fMHl3vBL
b5/FKYRwStCgOtE5E0zKCdtmw3HqbuL/HQBqv5Qz6Nu2blb4iAmzMqomE9ev9pM2
GkONF4FoKs4x0tCCPCbJtsMG65gSL5ugulbBbMJgikIYM7iWjAlQXen66rRJNF12
YagIOnqwhTi5lHNjO0WEKwTqm+Z7tFWIZKFkD6FAq1mox47tHFtEZUcpEqhZiXjc
9CGnReMGm7tX+qhZnkmadPnJsodxcOGzWIZFEM9S2AJzjVHJgHKClJZCeHYH9wKH
D+UX8sfJng4qrKA3hrKqAQfZUA6FKr1LmFb9JymDtEUiQErOO4uRoVxU+wVPVa2o
aoyE3tV2KSdWi1VpPWj/ZlI9mqZnd96Vs670nR5aGamsQ/g0hVnv+WdLu0sBwEFZ
euuUDTJTPO76UYI2h45mLaauDKQqFqsZApb6jO9MfS4eyctkgg5xRu4tDvMH1WDE
2WcF2V/UsTj76/h/YexAoTTRR/f19jA1yPhupL7nAjAvfbxIMbmTTX5YVq0yOJNc
EzI2PoO5/RR7rsr3+8oX078HPYLxzgVClvTmoGNmq+XBZutv7CQIxehafYpaQ+S9
1dmAV/Wb/XJ8SgK97gPd5vFA9p0vS5gsLwtQDdJg7gSbyM2JEiGPaH3qFfsqGane
BDXH1us3LJKdD0hVdQs31Ts/2PSO/73rBJuOc84HQNTXf9uTsPbbDmjzB41mQQVe
XDhUIqAF3e62DPFcel3o6zeEDOdvNRYk5HwhxN3u0SVfI/DYQcSVpmJpahJLGD2j
k5C9ZdXQQB3q3ZI6YijpUqoQP10xQSoWaqyOWdL2XzYBaWWGW9TS6ybLG0DgLyJ4
f/9xUlHlb0boFKttBl/7LFD8ENx2WmDaJQea4iQp+M7Db0PLeUxJ5k2PoudUg9dp
TuGYtaRB77qJckKnbkOA1CDYi6S0spfnDf8Sw39zXce+H1OsLSkBU8ZNMP+vHAfY
8D7TBIAk6rz9r1nUW4wsfseSzjaJrj/TM/wLHuKS4ng28XC/5g7EHUSKZFet/+1Y
L4e/AaklTaNGvTD8VH3uTLL+FH9EIMg4bXwwPnGK7QZ8UV7AUkxkztf+LMbeUCFl
1sm/88osVbN0dboTQaqXyOLp+JliHHfreuvdqNXNNFVuesGxG7iWmHwnG8VQcbWC
xFJcv7Cy4eVP/n5S+FSbchlAZWsQV2sF1xnTuPNVtQvcYAU+RVF88FDnjGAJWafR
QhpEdnIwI4KS9aZth2kLdiRghQlSXqlwEMH2dbFCUoQhf2bWJZs+r2SGeiKpKIHW
76o4L/1IZ7Sakxiv3IKr7qoN5sjpz+OPXMiRK7tlC7ebOPIwX5e4GEcLWTO8vRYJ
aZYFAkbn0Ole5RjT4ue8fK/Fc7AyJjKFgvtBCjvu8vwyMeSqpqybMkH39IHkYIWE
c7N7QCsy+/5nVZ06Ox/NBnj+wxewzS7Au/nFKcrHJ+CZkLWWbBi4YSbI6MmozohD
uKi5ot84y3ReDjwn8ek/sbeN7Cl8Nv23HDXIdEulBMXVnZw342u9H4TYrNU3pHlj
fjimYijWTCl6kbcRMcFsIavThOWDgXoXzQejgtwIag64eg6cqfHXKFd75OceKAUk
uSI+H+Ap6i/T/1FAwTfnzQcRa3eEcHF3ait29QmhI0rAkGrrWprvCzTWP8vndohu
NGs0YzSDeGq/s6ItscQdKHDqWoymkN+EBO+2AI75Iwei39Yf+8iQ6LZNTMz++9A2
zBwxcjJOOu6LdXG6fvtEDj0z7FU2ZKBObSP1MnuVhH11BylbZ9cSpOhdOcskazPc
ceS05AsHIF3uKiesvCdDcQxbaPZU/gCx6OpAjFg6BAtL9HE1aUD9Za2xlZ9dOSO1
XTQBw009tToMKayA9QbU2LfL3NNIevJn72RBP2CVsLNd1SJtGPXvll9IRDVLFgX8
ylT2ot2lHTBXEBwHIuxGDcaY69+n1h6JR5rgUyN6kb27O9PJMrdFDt/4zLjDm1zR
J+RQW+SO8zpgHylr4uucooEZpKZpLBosAdvGMExH6y1caX3eijODZPDM/0xrMWL1
jYXcbEGlxfFtim0C13BAxbX+aP9GtiI3t1BTOqFPQgaIdwMHg/zA3xGs73Ka53ve
D98+gq17sshAxYJ2pjJ4nDH0posgevx2eq0yWXzXLt7JYZCjiiKdXvn8qykJg3Cq
4cgtZbrkjt0K4m649KwsQiKhewZvaNn7FDzyeik3QRtgzb699rj5PCjMBFva9jgs
31YdtnGPjDih0+thukcS9xLPR+zmulzcC78oaR3H+0wU2DnfEQGldZ0X1fVWbNQ3
eqVPxtT/4bH9df6z7PiTKHi+t2357Dic7rs5jMLzCtlB0b5K8QilbtMRy3Q2Bked
q6Teb3jc1jO5V5hQnf9cy9kzBnFVpOtFBQ0vJKiqp2vA0XfZ/054ibgV1ngBdwEP
LARY8sQ3olEsWf4yHCLKMlFIY/7P2lm7y2JECdsxc+USDLrwiVafofbQgenv38z1
Ss7GCZh/FLH7eC+vOALWFxQViccvP0drMqZ3heMq0COkmYKq84DJ0tgk2FvBopEy
BKyhSp+MQ+2r4wM/+m0uES3m35yZcPAstSV/uRVJYcgqYQoLEk00Xr8hDL3BQphO
RZ9E2DKShqGkL/3pjijpNufajZx7NUHORocFkYUDYQtOKm0JgitSJ5PEpZU4rBwk
eU4BFU6/dv3TtxyyzpzYy/2AgyBpJ7LpOfipkk3FvcDcavrm8jbtSzdY+MrHwA0h
EzijRJ/s5isUSwK7GTFeJRANUhzvXsMs1vMrvIn63Kbyifai4Tml6MZ5DtUOK4zb
ts5u0H6lUmGGxgodC0xL83TrVk7YJn2gHfl1IkAxb6iEjK/R2CnMFnS2MqdfSByq
1cj54W/Q2MI+qa4jBfEhwrESqOGVHIRLyaaFGklOVl7zJ4Nt8n1WD095LYaeGm5y
vB/UFcZtOumBslGWKorMpyHPNRk/hlNPYZrovcBtyB1Sr3HG7VdKXGAzMboGCXjH
XR4v27kIojvlXty6i9+GkGmCFC2bfpGayQ7TQic4U7kSxLMcKC1d0qV0bcxT6XqH
9uNYkef6yRfg7m/m7YtZGxz3veTGNDCvzp8cYAGnIHRVHlJJtQi1vf5vJRD23MDj
FJt+Iacg7IVdamP1RGBk0Q1B/2IMPL3j4yCopuM2wp6yPhGkDFCqUjoGrFjuttJC
EsawSPR/Kn5gIODj0Q9ThUJuiVRQA2wbxVh4BlfaYJPDqa11gACuk9gDkhFrOw8Z
49YQ0qa6O4QXW5VUlsHCqc9mnbgUIxS5IbDYpf+pTshiKmrzcuCpCd/xsigU1fgf
9WqmjRUjXBxX3QP5srRAQKXzkWRmQRS+6NsLu1iW9qZLFiYAc87CLDfgUd5hfSxZ
l+4db8/3MvYQK7n5UDHn0tiOB7gQDGtIotIP/6j3UAlr6O9uwx8Q1Nnkplpd8C73
ky/9nIFptNfw23bYDzJYSRIXJgIlVh+25T0qZqeT18Eul0+CF83Wm7g5+PEBfkqA
9edcBv24u8lBv7cc9Ctqa3gInVtR1cyDHc2R8fWsBbsAK4clspdt105ZZ+P1dY8x
dYhbGd8uPeOpffyM6IUO8sm0Lw5+ooUU/nfFrLzawc4W2q7DEsdBgym8KW3JPZLO
5mZ2Gx1/wKbgAR7XSo6MQgWOEwN+oQcThKbUznFfLg458ceHX87WJpg6dDdXtlM7
4mpyB4Zg4YiON4LSpbvWYGT03+UtXzaO0FgHhzu/zu7YDY5BUPL3pUiWh6W3G89s
GDf/X0l5cwCI2xFlq15WxK0T8oin7HJ/2AJcJYafn4u231bgXVr99ZKm6meELAXZ
SYtK/AL7TUsexGc7duut2TH+Pphea6G77csr/ps9MhWQfUorwauRyvTxyJvmu2B1
uE/XGOoRcyhwTTrvxqQVm3dYycLMnWiCdd8RB1MXZYYw5GQFPkq09OHesJ3d/YJ5
KFPIY0Vs0ON9hzanmxYGlQen5CNqKDX1qsSRiuOA4/WIG0SptZ9Y+dja4bgrO7OZ
KY/+91LPR9gwjsaFhy48+8D7SI+wB0zPzs7fOXI63g3g+Tld2Sk4tzvwJRvr03PD
BT+g8Kj84sKhAwNEmnrxsHuieYORx2lRx3pbSYeX+IPFxjul8bCpOOXsTwAdx4w1
tIUHnM+aJ1qFsQdS2jUIgO4XoppenDVXYGERD55otkcq2EgLxLGzu78XuHOW6OvT
41hoCJmTTvl/ATcnhcJ1hJ+bO30CsYHQT4h8+Q441qhiZLceL03gItizj2gpEWsJ
1AIJ8lm+iLEdE+oEQzAy1sAWGZ4P5gGnzR25QDUlv100pCaFo/97RU6E8AU9zXsP
em9Wd5u6AzGmiYxaFWGF0cRFP4QBr+tWgFyW3j9cSZqvDwSJW3dR9YRXMJ2i96BX
aZZ5GcoQw0N4ScLfBmwt7lSGEAU9lUWESkzS6rY14tBP0X4gsFnYo6oVgxnnCwJi
q/33a6nrKltZcl7/kWYMWSL53BdziEBGiCOasFRG7kIjN8/ierTVWmTy7kZBnYPL
hh4ofw5k8Kctnect4yDUjVTUy3c/HBPGveU359Mce3tnyZAGH9ZqHQ6Eji0GyyKg
0jOC27BXLpBm4LUo8RtJ4YD7A85/h+mXKh5ju9VgPnNXiGwRqknfLr1uP50HsxBM
dvMnLfgJkolfn/6tvpUvFfBC2DYRXQKVDmVrt+QnYklmmft0iJbvaOygVmC1QmNM
5EdIleMoZDlfvTwox2yhINh0sNS5fQktbuc/TxF5RvWtmMAEFM3rPhMCRJWpfSWr
qg+6IR05MqkMDjrv57ABwe06l7MsBtBydSXwPlBH7b3QKuUHjNyE1X3aGBan6rMz
cIOMC92BW9D82c0RiQVJFTWltb71vPVGf59Pyf7YsSCs+zzmsfIRkBVOalhlAetd
Pn4yuUNC5I7YbqrAM1IlSjYAOvcZIk0rfs8q00oxvOJ33y0OQ/OzecIFy0iwZUJ2
IU6jl5xB0UcwIQWR39CxqTgvxq3UBPgJJAoQrIU8ehrRCw2/T8BSfJWA8udjPKOZ
qSNdxSqScSnwmuBGxFtrFhXekHSQ9ZdrCCn4V39JGTfAaygxidXpG2GISNqK3C4j
R0X5g3V5qIoeYVVupJvZxuFsHMK2hwk2K6zbgYnvQJgM4W+Ls/rYXw21C8tOAHRl
waR8d5PB9qFYxDjszD3oq9etsjIgmfUPoD2TqSSWPq/GZwXLqlJlZya84ST00H9q
yyMCcITcY1OL2T5irx3k1OG6acACi4oxTEpGqK/EJORuhFLaWiLsS3PIhm+8kpr5
LbygR7waD9c48FnMC1tY4HBVvXt5gDOmXDl6Nblnmm3ZQQpgB229R5DS9CptNraa
eM32EBWf3c7WPyJHn9Tr1ok6Rn4nE22zL2w2d63PkJu8I1qRNf3n/8zdlLJycd9a
nHgXMdAg5IZIebSoHMLmHaRGqsTTbK8Wgq3y1kBKqz6ixx9b1mFao0Nz6i1w17xG
9eDuZyK8QK4zPUA7WBtxtlXfk6HnLyb1aShKDgMj5hXfByqZmlfTU7Yolfel5L8B
3GT+qopd/oKKFxrXFPfcStrVBMKYAcKA7jnJkUKsPk2QE1FocuqX0cvYcDk7fblm
nKahPH4Rkidm7g/jX2pOgy8+nfHj1BOzJox3dkwn1dK9CJRfaYWOMuvXIP6dovjx
6aSUeOgJ2D0gTzef07L72fqBXa/1PX45zL8VrgJ0kuakftpqzjPnzUiHDJT1QSwM
OP9/nWrW296e6jZHNcKpOm7V/fRIKkdBSiMitBOkykiUbb2m0NKOiwTnip2QxNQI
CPxJMIel5LDB5ZePotx3uIeniSLJTWSPhEs2Xh2GLlsWglchKj4iz4/3Q8OhV2of
5tCrG70yxrOBs+Z32L5xrobD+KrMxtottAanU+E7qLfcvSiPrwJVp3J9s3wRnFem
pIBRyiUbKQe73LzhlsBZsiybUBY/dd++QFTzHSWIp3rqo6vhjEj5KM1NotCzsXJ1
yS6L19w71G9TEPq/3LbLWUSSX8Ozz++UAhwPXrEU81WOYdl34z2MmiHlfBnzm8vl
9weCVCXyxoRQzs8pls+IoVWIHXE9T7EDJL/NCbeAXwnx0TgW1igAeu4mm6X9b0RZ
/tOkDUy13bRVlsDk5j8kwCUHzz91q/6Nq+trgVT0SL4EzLlBdwiyMNzlDvyUs1hz
J0S3mSWvqlQ7pH3E30E7uA3AqgHRZWkojwptm9XFk9f3fmboCEuRab3N1e1MEWuS
iZlVh1Eqa6KXU3Z1uGhQKzG+P3sfQDbIiVaXRb/aOKO5lcXqd8CVRJPHnoUNSZBo
QFkYS4wC/SLjOdezQvUqdRVO6eG68tV/1c/dn8jWbYDLf5Y+gc2Nu8kvA4BLz17U
OGnEC6kcgXGvr1S5Qnw3qWjWrd3F7+slW6U2dqW1NdS/XYrvxwkrGsK8WG/3wAxH
1fQ0zhiBMXQoh5x2twElYcql9bZVqt2ndHvSh6Xhsk2tFjQLVFLXBShx8hs4TkaB
4toKS39trVr68qPTvEVVx7byYIaKOWeQQOX5PDkLGYV4kpGdOyFbOpE8dgvwP+AB
GNMgIuzgtwunOvg1femqrKq62lHd0XA+cmMA82mlwCpfmTfJ1nOh9XYzggBMhYoH
Ji2hBn3L3jdHTG68yEUzWYu7P6fciJiPazEnf9XUpN8c/AzbFT2p3RykXIUkdQgY
/pW7O52xdxkuGohX/n4h++X8304jurB+ibDgJWT1E+lC7ABuwngHTKHYr096eVBP
fHzc4iGyT3GnXpH65MlsHk8tbPbvRXLWZBq/71uGDFF6K1GbUrFI9DU5364wdxWi
/3OE0Rh6muPmvJdonteKXZhb6zT7/2pAaRSxfk8CBnfoHvMlcfBc9ceu+AtSqpCs
Lw6lhIjltfKqVSUDNiSvO4r/kh3Bip5IqbFW7f6tdFWxygn7v6AklHdy+PyPNva1
J4wfmzj8k9y6lzS83dOD+IzECgr23p0NaHRBNUIk8Uwdtmyizujk3EBpjlWJ6lpD
trn69pWFract6liui7DJdUZZRGJhcbgfTp9/5jmTsLZ65p42V/yE4OMRBlusBMON
VFU2AV7gfUmXlDgI6NjfdYcF1OivWJMhdkVd7FMIxLIZ8zges4oe4BE1hiIOqH9v
LDt1w5EqeSyYIByW+uij0WKKDp+bnekcMTmWPzmvLzHoZ57IPyBiMlGZzG/IRcs2
BYZrIA9OIvgQBbqEtFRL4o9uV09A5FFzsDjcoxqtLaBTzRHfjDiSdL0HkFBSzXMr
s5KZyWO5oqqryLApL85PslcmFsH1zHy00OXq6pd206DW2E6H1pq3DBr5f1dG2TUC
E/rfbhDxpLQ/lDKW3UIEV2D3MTQYxT/7WH8vNrME2L9wz+GXTaQLywqccnAF3O8e
+1GqHhsZKLUBgbJUI3bfD1faFHsU7i3tTR6KAh+V/BViLrpo/dJtaX681wla7M3M
YRpM0ZEshYtewFENl/A2gGrKJpEndzDHjIoO2jCCXcph4NdLRX5/y0jcAnsOal+a
YG1O/NcJZZRP/jiLz+wsnHDQ9W39iOnl6Q/3sm9IgYIsc2SSdk84AjYosIA1AFyA
xy6H0dNp6hl/yjo/6tt7/xc9X/q8aqt64r8Z0/Sp7eQ32wIvEEQyzIFePwh2HgX4
olrNOlPpWWRROAt8fmK36qn1bB9F1DnT9uT/lWAxOi9p8Ytb2ejjf2XdnZqdBQpK
Ei0ykXiHffHrqON2I7mmQKkCts2iUy7V4LDULPnWXTLLSEgdGIvo/B907Bpm4GrU
5FAUA4dh/rMnz0p411tvGBtsIWctoez1IcB/qz5OiPKPjqG60rtAzYA3AKMwgpbz
sDY1EaoRDAU7reKr+wUIDRHnpzFLHT9JF0YDIzJOxK/ow5fRQRA2ZN07Vp7dV0yN
Ki4ITo8WzZnLri+RqIfLvzHKUo20pXCB4TLcygZGpkxQhTopwhQQT5wXoQ3l2APT
Uq4gaU0Z7YUMrkB9qedO+B6ZjOahBkFk6xnBk53UQp8A/jyi7uZuRI6aFgv3xhGV
zQzkQcZULm44+ZbLIMuphjWDQG/TsmkrMJ2NTG1x2ID70Wp2BcWJjQdgTqHcKjY1
xs/wk+N6Yux/YuDyk9uahaJwdcqms8YieJMYQwocZjvVeQHP6X28e65R+CvQyo7x
uqu0CWtrYKbbtgGGtzTvsEnUFxv7XDRQc84T+P9T56xBkDQMvDXfnXB5SrPlhXqc
jOFdvPbiR+yWVYQqmFdO129I6L1zf6D5aGVQ4sry/Lm4AZ3N0pKTVYnISvLS2zN8
zx/ZYCiWP5Onm047soZeht6QY/79VmxcQDvnJ0z+W2enOOyV6G3gl3ViglWIF0+x
Gw0IMtX0Y2l5vW+LVekloA8mVisR64CiXfzNuJcVwK8snva7l/8Cn0PaHcKpTUD4
RqkeR9xGvmqxDubnLxvnI6z1ZFmSwi15wPySsgL2M4qxAc5r5EGCxs4fI/vBPzqZ
W2jp+gQhyMntJSbeHgXPNkQgggVoYnFj2w9IfKWtcU1VHjZcSXtyStBbjnrjliTO
z0SoUrARzxuoMsvGOXkMi81pGGe7PGZkoNOhHVWcFkJuFmkgtx22B38ZDwOylHur
qnAyCsgNAd3EHrvWEgvuqYwVArCkC5e9WLYl5+ZztmQPX0JDA4pGpZl6zvOOn6e+
bH0eUnryKe5rwZMqhhFa8+phqyEKjdPOT3wc55Nrjw/4R/1//5Nt4z1+ejcZX+rO
zqbkrrSEjoMTOenvwDoEFDUH+SP9S1hKO7yXAKmvUEkt/5cHCvSGtYdnuWN7aKvr
lA+N8STl67hP7w51T+jykJN61SE9l1R/a78Z0JtkXmfa21LZtAYbVOy89S2IAv7p
SC8HmlOltPFzPgCwSmFyy5HeHuvlZwdm8Ehqo2VF15p5JCm4YhzcpGeGA9niuVSq
NB/cQDSzzVahOEo4dEdzurpo9WJg1B0Lr16UeLwN5ALqxUVFXJQmwxIhckySkCv/
WdA25j6HUKebb+aw4qAt8kPkBsvvgtpOiKVsoWmwRTPjrob439w5yEslxMoS4vyD
xymTEHvr1si+TpmghsnFRO2mls6tmSHz5hqUhTxwehek3Ky1N+W5iaDkScoR4+1N
VdRFtUVQIj5KMVxfpeGEbnzOzLwlqhq+JdTm/p3GnuCXwEEzt/+4JXksVmho2hLE
JE2zdTkxJU/BNaPcvCL2fFtHsxVaB0FV8QOH7MFOBadnuFgP1Ct5W8eUxzJbXpNW
00+ZzTf90MytiYlFjA8pq4AC38aHUEnsIQnodbHCCGMaECXyKkx+Ie1m+JPE3E+Y
QbvW0Za6211A+5dpFrDjzP159JeBAoJPkx4L4bVf5ZKgv1exomIti99hdqlmGUOr
UamU4DCt/fkJRUI6uklaPfI5eudtpLQAk5W/w6A9FR/oQzm1X7EkhG+wMUD+Xkdi
pXh4QMWl7QfeL+UEForLsq2En/7cXcKbsinCJIXgOdROvmKYDC5Ij3aaNZlPP08S
PhWnqeyQe1yeMusjvoHsGlOhNbuOkoaBBM6T9PKRvmv5fen7tHEG6gdgH65NS6XJ
vNM/Nr4ykxqI5nmeE3beAa3p4AiN+UiQao7htgFmLXYDR7aCpzw/KOQY72hPPSMO
i79VCDbzwxfyiCYCl0SlfcikGkPP4h78XERSoFLMdMz0zlDRNj+q5VbZ4j0+CB/Q
osIx3GJJp4/M1K99gxjzQqTzMamp0zU8yUrPtrN+T9z7rMD3QftWjBTwK0JJ4J0p
FgztYHM8TVUWmZYHMbum/I8L73dI2uPy3YzsyPqjD1jvCMoadhcX0yjxZ3feq7y4
iN7SWc5JY+qk/7mKyYOPk2vYqIJz37zAWOtoRVW6hRwhJcCNpPQyFHrREcUt6uEc
nQMXZBaMDqT8xoSeqTaRWZIV2zv+zJ8Tvzxc+56urNjbp9KWeeNpjEK+H3lXCbYj
+NOZBehvROb1dBeI+yA6A0WWJEPRfm03zyLtzCjt0VQiLcGXW0ZXoGxX/TJab+ag
V2zZl+ZO+g/HgBdV+lOfpxS/PlnV5thqqB+mZSLc7CWkmxbP+X/TVtURvnA2AAYk
FLwKi8MXs9qIA71zOunBP6jyPeBqUWkdCnstk3QaETc86SITZbM0pONtIyeXMoT8
U/KfEBISDABzJKXDjcCN8KknZAnssDmB1b8gb1qXTBgyXZFm22nHx6LPDv5ordrE
HYNSdfQlzEzJc/xsqd3d2qrATebLMvM+K2lbrP5jI0e9aGfKGn4kzSHItTB54nqH
QyA1g3SNov3otbse9/OhmwGKNIFrKnoLGSdV1MYEitq0q7JUQqMyJjoWMfm9M2KD
DX0WgWqpqlhO8pMRhUe/eABllbYnOmoCG5vPc8B+XLNnenZTOZIUOzY9oMwtiiJO
/mqHPVTVn3x/18jDS3Gta86CCMSKlXMcBxixGoLuj0fVoXMvZK5PFk9CVEoHPDqO
sXcy+1qwD5fCTmg1p0PbUS9JlYA6PMHcm68u45X9+SXEqOPyFD7U5hg+MO2CXjEh
3S2ZNVb0z3kfaTKQIEKb4GhXVcst4ZACAD27o7oSz7MEB6igSNVTm3vY8/T5+3pN
hWMXderlk/FbWefv0UJz/OFd/bRGYse4R8YFEqGk23f+Jg8wZJOhPjAO8QbsOmvf
heonimdbALg7OqjoBOEB7EWRr6usy47L9/bZpOCDmYP6jigQvhqllpiNrG3A8NCF
QEfRp3TzWH5YKmWH/tsHopocYTtzbOF7fgOG8F3SRpES+wQ/5ThcR78nzGb+zhQj
dR+CmJax3LTSlnK6Ni71toqDw0PpsDWCVT0NehGQALQO/IzqD018HQPOYfeTR1Jp
ANHb7GLT+3jThYnxIlyKvv9CqhyycsfLZTk/v/2JOOoL4en9iOW30mIZ30l4STNW
RFv04YktwRK5uZIxgVyDAGlaIfJrPecY89eRCZQhEH24Yth02DVGk16Vax2NKp75
ySRF3v9vHIvdHbuHrSwv7RU4GlvMiwcIK2M0Ue8OvWLXO71/itcbRnL7qAsCT5C8
3m/5kTjZhsUywSr8OC+/nIAaHVH8pB7UVq/HEARsLBYuNDTBkoU00fuYzIg7UTk3
fFc0fk3IN9Wi5b5dew64VMnINM/o8dl+kh9J2LL/T1g9abpLSllHCawG11Nx9hKH
FpoW15GmaCuvQBcmO618l+7GJQXESPv+68xE9dTCmnznGo2w9jyPooCSXzdwE8u+
L7/EM9n+ywl5q7QFiTeS77MjphnW2EDrPpYoPGBV7JyBAcvyEAu/1tqhP3Q/ac2T
i+FYWeB0lWiRNa7K75U4E99ItScJaUzmNizev8drGWsz6b1eHq2FL2XjDuoxLiTo
vk3I0bfhv4Q6D/5/pMyfquX0ef3gii/jMx2Gz7nWDZmJ5CapzJ4i2odJRCeeE6OY
wOPhrPE0hpen578FiUnloSEXJqAGTqZ6dwetkVbMdo/tILj2eDmW2/+yw/wcWCSz
hJolVRElHBXFIyGKmXdlPXQMpuWU54t40CU7s6SSbccUe07MVgH4jO5T0pbIlVM/
PYOa6+nivpHcpZULWwQReJ/nrGGIaJyYBgE2SK/gOrjDVIgkB6PR8V+Y1VommJ8U
eH53bC9STPnyRVtSZ0tfjzZz9kBmhSguxxV1HpUnYlcOObi+re4YCmSKZ88HU5sG
SIOpwpcpEATFdqMSFTAGXnHjxPNwCcZx6e97jRNR90xHdznyTcZ24pOyJTMf8/k/
9hsxbLCqZF3iLwoESfXFTK76to2eaVxEEhi7uTxsGaaixcaiogwfYmFbmCRtb5Xq
miGcGHC4NUXfMA/pMtuU+5eOfL4Dc9+dAJJB+iT6o8WEu+0c+95Bz8vxtG72JFaO
DAm8ZpjaOXPSQpFmNcKKan9GWrK7tLHcaZ7NsHR3zC0USAgK1IOGcvhi/TlaAnFc
HDxo2btj49W4mkzamO0GcqSkkUVcV2oRe5wG+ou09Qtah4zs9POk2TgbGW8E07i5
JlLczQkbkYehA/lB+SVwGzTZ2mFNcUyNjqeWEWfZXSru2VLzJtW1G9hq18b7Xz35
reqEwQE5R6LSSer9zpblwpwJWlOnkoveadLZEOkiUvKwP36d5eYvI1jWhFbqEDqO
z9s/Q/k0V8ianloOSNVNFp9xQnMZWZm/cix/NxLrLw2r6xlHT+QDVXfV/XfOpXDK
XTZqO+yA2SujZIeCag4EhHIVxiXbvleMtMYN++ixvqeuYtcS+R5Qr1N7lZMqGMzC
XxDmxtM+XKT+RQLI+bXz5LC2/qrxZOv9fsJ1EyYoHinC9fSIOxpr5V5IoWc6vIiY
p6pm8S0pq4LTp8sE358HE+jnxnuKQmAxawh/3qCmm7512QAomX5wODzRSg9DtvL9
og5fdjvqZi37TuXKr0y+R80doAZvWoIteaMMTMK7sD88Ou6GOvavz+vrKTainWYw
v5LcqprYWUFDZi6nmLbOsSLIc8nrhoT6Qx4wYhW1aLWQNmUPG73FylQUuQyGK53v
LvcWf5556S7zSlJGivd18Qcb+SO6VC3F4GxCxrUiXDmnBXNdml9IescnsT7VUKto
da49S8Hv7x8Z8s7wap4VbpgWZx+3LO19YR+zXrDwMXSItHlsG8dtAiKCTe5uZM7N
gZOD7XJSiXhTPVFkWlNMlATa3SLjL2ydLaYHcU/SVMezs9bMJMBW2nxQM7QpwGjU
xnh+BGMu0B3BP0BFz8g7aG/5Q0IXsI+5EcQrSLIH4i3O1rKxmcLaObajmsgC+VcQ
LZHYIopLo+L3YYWUI5jK49/M/bCJfwVMa5W894WHKr4vU97W0ZvglAgFwzO5fSsL
XYWWFLvd7nnPnDlfBNlMOaTK70yDsXf48CqkLF+IgtzUEJEdcmY2r+tlt/4RYCuj
EUqYVpEoVfJBYolA13jgkd/1L8nZUjSxz10UjsajjlplGOpctJkzyfEdQjaleQMe
8JSacJtjFubrcG5AKCFt2Bh3qK5rKr4j1XNbJBCfR8pIea7in/s9nYj4gPtG9I/c
6Dot3WbePHt9idZElDrn3Vkdjm6fO7OI3pYl2edgoObTTqfyI6pQ5VJb/S+P5evZ
ZUPer9e9nl44SFzG1wPuCUHzn9w6mp9KIKsifCwUh9TYpE9u7s315usZJDqP4aZl
0HOd9miylW33Wv0qWxFElqdF0b7VgeE7PuSqxRN5Uz56S8x2P6GvZvVvOaqPXmhs
pTRt/ef0qTUFaTMuqY/FJ3hNnSLyoGtd+/KME5Zaa32LZyogcwm3BpEpEQ6Vjc8L
dBnmS0w7sVxzQZvK+cKHJftiaHOIs4y1qUyJrlEcyeo6UyLMMgmIfp5xzzMNLv9D
i3kM0vmnpoQdiOUJXyMHr3c2kVE29iCsv+nKGpoezBOsi7M9XdVsVkQCiUBpgJAT
oRmXSSkBWKeELb4zg4JKSZ8800ojnvWjsQOPnQMpTcQbR8k4+JSEvC5DS7ZWM5vt
j5gL5zd8egY6WbA2cvzXNm4wYc41paLhsMXc1qZVy7TUMxzVCoj+i54aIubBwUsU
PmoXNCu0dY8/prn3c+yuObIU0ybB1DaUhd0jXKksMXCqgIYC3TKyS85RITCExOQf
tlg2CiLH4JH/6kRJK9eI0MvgMAqduEVZ9mt9P87m6j/FcFGsQcK8A6in8nNYZGYj
Enut+OUpapxYh/bx/6AZ8B8mzcqCE6LT1ccmXB79zyHRzwqyfTIfbn++LyoHpCuK
RTYiwtamJeeRmbYiJ88HUZb6F05Q0O0GZ4PHlmZ85Q++OnOhl8wCQ1dHcm/fmzQS
V6WCSfpkv0ybimfssk85QDHgZK0aIw8kooQi3bUmeNcVKEXoteqPt0fQELy/qTf8
+JoK80Etr22/Ejp4BuPUSjsL/cTA5BtRh1fV03TjgEWbLkgqG+NQmG8JWYAVNZes
m+m/11jpJNK/yHYBK7/khelTpCIVZFgZJHbCK/FEOHJXHa3AaOWoUVdbbNxaHQMv
EXW9aQ9bPDVCxHgdJcV6DjnDdMHFSJnGWQiXoaGQKnNg3xnGFKBNpHmGzUcRuG3p
V1qIENg0jXmyZMapfFjFQdtVgp6JN1HjDtcHwF6NozDyWRkbs70ITuoFhk75RdFn
3Ndvy3JGNngoSJwnwv1uyWCcVGhAizoiJcwVV6HVGwlz/QiW4BJiQ6egZG9mXmoV
3DaVVVzfs7+m5U65FwycfkAox7DBfx0cwbm5PrsYUMtxo/cBC3iljBvEw3XLoN6u
p6khqOrTb9w0erw1Ck+L2/k6W7vOVK4lqkiTZUNC/x4FBJQY82j0eqpYRBTzINhs
pk4wlUbxWXROjCtFd9p3+GsltK8++An1sc+KDgqXF5ld6WqP9kgTeAVvNFtAguLj
viD1NMp/Ixz0GEeG30/EFkXHIaNYxmfkpcbn7gWvX46bXX28bhztMg2XrB2oxipz
TWP5+17aZqAaMP4iyV6LWOJgH+aoz5DPhMFcVqMN79tdtQlVRmJ8OeGtJCLd5eEJ
l4pNhpgpfoBntKog5KNE2L7E3caZoKxKxnkDlN83RNCKPvNt8O+7GurBN8aRVkg4
HLhFcFnUp2Z8lGmkhCtFFSllMMZ5W2vf5aXROuuLfRyt8og3hDBsrpOCsg1Qns2H
GUuXHgF+RncOQ5vt88PHu9QfkSkjyaa952U70AXu9naKNHRSBJtSEsWHhKI2HnDt
Hn5fYqk24g0q7/Ho8JOoM68WcfCZjBPaW64w3ZnvfMlELvwg/sMx+3rbFPVftUuU
+WYMziDXGXFBE/Hg7wq5Bu1KDFymLxjkTD0Tejc6zKQZfVaTLGZ8act7cDNFAwJ9
paJV/HT2fuBa7mZZZFbZN5I0zcdxlKQP+3i2aV9i5qWS7KYjgWmC4LsXZRTZRkN6
dTc+lEc4D3Ku3+4Tx8q3ab7zEuubDOnVrgVjt42IyEsircAq9vZ/9ermfsXYWBI6
wG0+dwiw8U0hfewV2HYRKhzMGIFNPNjukDWwVkDHFs0g/aUTOSqGCsIMWmqbvcim
WDjSFzu0TxQtaEmKtJqLfisPGu2W4wBIkxI+FiSpMj7yhOS8wLGpMGwaNPIdjPIy
a6gqP8hiYvvFwZKyUk3vMud8jGAeSdeBeZ7IlXr9Yho/bA03oImbDd9O8ooepZEV
VI2coyuu9OTfONRUrb1VfIPvLs5laMaKy2vS0XFKtoYp4hBAfqbPkKz9dNlNysFZ
yWCPYpE5HRY3KlNKGa34tMRCxNP3HXZLFJao9+dMrauQzrO9IXqC7Amd+UPB1FdF
Z8715wPk5SaX3YZYun2uM8b+VguKn+bo9a2zFUNH1yyTMTwa12AgvOTJX7/aC4xf
10QxsxocnIKicPhW1ojsOxUdpkSn6L0YRSOvKs1ZZLfZbi1MJisRhvgx9WNExENr
570rPEzEF5eYf1weCjDfXkf2CFhdjplVoX0kgnBD2VT4y4szWQWZz2qwsk9N6RNi
tt4TZG4SbtN2dhArCUSH83E8QFP0eU3caCHbo9IHUpXD7ZeIfDKB7FMldRmpNyH9
Y+0pBk/12tUQV9e+h5mCQtc9V14/0aRSz41LNJsrBKWZRvJ4WgoXU2hvHfHtfk87
glzUukhlwQfbD1Ob3BsCw9cpmSZcDQVwTYlcVVdxukFUkX7s/8ORA1AIzzjdlu+S
z9Q+UW1NhqofY5XX5EHdDG9xG9iUgUE56sMQpwOU0rgGHPON/9w0JicvHHwAKKOQ
0TgTF9sYofWCHMrr3DzSGWjr2gE4Lxss6C18lSsProxsFqX0KQBlS8JmdYCA2+vg
Sv0ofjlyjtAIvhFrrUJCA2fZnN2mwoirfkOhF4GXZfv8+VSKYkEhrvTgjx7vagr9
hEwenPd2qPdkLZVtvpAkGNdilI8KAAoTZzETNeiqwlXoRwt1x4KjbNeWmDLDAaHx
l2LHO2AwGUNRad+k5ZqkuaZWQGsnPrGgvoKyABby2X37vECnuM+6JtGlRzWoa3W9
UvBuZmC9S0XDl8FVqNYY4fCV01SwKil3JwY2u96mY57d40CUATw0VhuZrPHLtHHz
P8xV3bo9nYz9d/rmTHZv+RAMYmmvi48BXWRsX5IISmtwozjHnoVGl3qfbJxc8CfX
pGx7AT+qwstXHrhOus8lMlIzVMkM79VoV4Clu/X4Kei3bjrQR7oqcB3bfjb+DPaZ
HhK2Tjks6pje6xDGzzSBGM/LElGLdT+6jWRb+BByibfL3Hh6CxjG6j5+UrNhXakx
9m79+lqJo9WEmJ393frJxnA40M9b1WaLodR+q3hZXtT7jkb3T4AmiTXUHzsYb1zI
LtLUq+B0o+6sisRW+eOLm5PJT4oVWE7TDP7BsopZEPgJwCLd8abk4bFpHEATbC5M
a61z4ZzjOMX/QpwEeThuZbeRD1/WNURwvmq2KjsxCdlhBi93fIqPB+aE7NHRRBAs
HtEKU7zG5n0iwLLxc3SOCfYoerE9UUqoejJL4/V+2RZ10Av6IsKq1bmkV0jU6CmL
xVkf5IVglUxNjaav+EmNf+xPTgOj26WTvOF0rdL4eCuKOTvpk+QoB+61H39TmSH8
9YMripdDwf1iwXQGBqOglSU8wKIhrXlc9UqOOfAjBorpIAZTxW9mocOl1Yyg8kB8
SSVM7DHl7NPfNrU29fkoFmZTjOIjD4j2Kf1SHENApv8LAzLUd66Xpe4JpDWuYn4a
qWRxg87z3MXwUikkBA/d9bKk2PrSLg+gPLFCiZer9c3h8LoU5859ciMWYeIN0Xao
c3tYmFll0hNvi+P4ouQzvky6SU48QklNRv2aprFiOZXTa9FcZ8VXBmnJKht9X/Ud
s6GWbA2BVZp7MG8uwrpz0ov9Qa5sJF8fJWoo0eYsqdcazK59FfessM19m25J+GqN
2Ag0q5pBVDJ89KHWmTj6uMe1hxubQUdBmiUiaTQQi0CHQcGcCcCxqhPpg1SPLVk8
Wvw/pRLlL78tf1dSjoIhvblyx7bjHnayuGoiE9/A7e7eFv9GXOZaQZJ9gHJaOO7O
NK3/lQGfvNSEyq+n8MCkSWO25Fk2dtZ0+tKHNgxuGztfcnf1vVehQ/63mMLIA8oD
TzekE6csiWqk5ntsI1avqPv8KkRsEXFTkC8EWyvAdrhy58Ya8PQJI8XtXWeS8Y0j
fpbuvBCL7j1zR/cgkSnJZnmne2yfnMShJgr7vNo0heB8HmdfzbxrYiMWRwOp9Toa
iAgWXBwOvSqdL7CmcAyuMxdeJPpkyMpt36snEUNir6JHhZkqfEdoVKfwOFdweWnR
n+SRsd5q/fnxu6utiQFL4JL3oAMp1f9r0HD3NU4ZcVseoLYfymqUDX/D4dfw+zGO
TIOui4mqWGi3JOcZuVDbi+m6VaSwAMunczW0L8bPgipkjyDoHpXtQQRb/SBILuUU
kBWC6dF5BoZ0YeBGFg6gfUT97F3PwHi1jdoDHFQMtbhRbvuutDOZLyiC9trVgClS
VEMDdhEOSbLFF4561P+EijVXaEgNbWcd9aWEHf486w1MziQQBjDvm3/owgxDETvO
hm28SDTykI1LH1gTqMvuVM003fzyuGVVdHJaB9zVfjQf6dlRVWUxZrisy9ysfnhb
FRNJqIjuHG/cfU7gHOOj2m7LZV6wvYnXaeMs53nBHeU51u43Ivw1+kjvqlEVtVml
NFxkXuPPoCNbPvWTNEjzaRb5rXG77SyjXzQ9vr/qFuGHD3YpOa7kGpML6AAn0d9I
wMQjlRd2ImmqxE8VJKBi8BP0NM9Erlke+8lptTdt48EHVvFcsITNbwejEzt8LTHE
+uOIOgBh7rWQFTeK6nHlRN3d2bJJMANYExnst+voyBXmUmN0ea7zoTePwL/chClL
7YvaAef5JfSRGyq0Tg+oQC9ZrxcTJXvGyj4juYUXh8g6nIxTbfQNHtuDspPJ6Fpg
xd3bckCQ+gxxtky3IFUc8Ju/MPFq+PBWOdaQIZfXwJ6G6w62iTjMZapOeRUqxAQw
BTYfSqd/pDE7i1PMdp8hOsKckqAanV87iZf8m1bjUKynve3DWmYOaaBDuQLjp/s8
avZeEcprRWXL/VSiIHMSmoMTr5HTudaMG47fiL0gBg0xW2PhtRI3ZKdxSaX2gb8Q
zkO0avM+4QIOd9vEnZOgne3lwhQqECCkI3V4dml/s1uqtauyklmmH24TDDQ29UQp
jdn91JPaatkuZo0QRyfAqLl+agYkHrI1W6jjgQIKmoG4CX90kwRH0ZxnHapyZAoB
09EUH+EF1DruUXEOxfvsMTDuhPjUUqaF6HH9wfX49Ksq3UzVsS4AwjSWv9miBOnx
iYw8EEwWjiqWM9RbOTTfmGZ5Z8xZBJ8JmobCAS95cA2CcpPsOQKKBjXZabKa5IYF
Reos7nSyVY6TDbtyy9k4/xP/4l2neHw97fRghAYP7TjzS+5J5jAU7E9jafgP/T/S
3YauP+PP3S64R/Owt6cv0SKKfWSS5gkB7oGZEpkRrKYCNB5mDApO7/q4dthIiYP/
UZM1Gs2nRPaUvCLpk0Xi1EAdz2G21EKfR3IY57uUGeJXqpmp7rRVPyVq92+Ab2rb
ZkmEir+6yCPKRLdBPuBZ2l2nK5fRXtAXZppdLCWPLwQpVYSmYKPYVgxECKOZRVqO
KBiPIW5AB7DJ4dAQJUDtFFeN1iAIE4Acj3AVSGIqzzeZ/h/gS8U57fmKjxKmYQdv
US/5PzX1P4Swd85AVtq8Lbf/D0cZMxl3v7JtzBAHcRe/zLGSdYi7XnKp1iX+Y273
0/Q3lecCeI/xmypV56ZfBcShQ5kZtuddK1iIHlONtbotQk4cDl+pMAWN0/pgQn9T
FvWBHFs1jp0pvPrnFW+EKVU8lygq9ktivBbkXddke/tij5aeYAaT3zcyVDH4M7Lp
yGQECtVuNF5vbJdarcWHHKXqC9vIa+d0nbEmAZBj/n/lI/UNc3Nr8slbnylbQh2o
1sL0XJEZhYRevZ8dWBgkxZcU2gOUbqfy1snCtKFdA6I9DD/QL2ntNVEeXYkPC6j/
+49PGbuz5hdk83Z7PG/VqePJHnUxYta4eOctheKn7N0eAtVcHuHE5OPrCqlijNZa
8BrsZsPRDPUhc+NsdXTnJp1CwqG8nqScwfwG4aM0XT9bDMJK5cMuYQXZzhtQ4OE8
5N13TH/Klr8x29FgW+ujI7//d4u9iMHOooyKZONxed+HBo6LmIoNzzECDctf9fzK
ss2NZNqh8fC2qUwCUbeplYXDnlKc2pmzQ+8ztGkku5g+WE6oWLnxZOPxX/9/0rBV
nfmVW2NCa9wiJPysHbtI7Cz0iiQw5XI8qdraPrWzAGUuCQN4J92kJSLk700T5YWA
mIFv07fnI7kp2Jk149qRAMGjSE7yCaHZcpTyRSKF/HAGnDzQuEqi6a43Qn3ACH1q
qQOwlTdzPnxkMips+yBbUXSRwk5xOY0hOqwZp3S4eGdExAWpK/zv4Y3/k/19ZIBc
4EwE2VUpn82mFcZ+j7hM/PLhiUPVkHJxAuNVucAS3VY13B+I33GLDiD9TtFSZkEb
UKq8FDXBMbFIa5C2D4q2P8K2oT4IauGeLXme11yapUTHJ2lhSSVYPVTDAiEZMCOu
+TUaNbO7wO4TKL3TN+ffFwq9l+fyp3amJ8Vj6HbeZ8068ADOEAPx12BXD6jjJBkW
KClXNWK8jkhn2oMqcgE32rMoPMuMWtqQB4XbaZimXJXgYYOsGS13n0p4yCls1WcJ
tRFdLp++1DFPYd3+i9PSI0lz6FSajC3k2CfnEt6R1BD3EwMF7O8jDU8Zy9O0wpRA
YD1DlywLI8+r/fhmQ+M4R4YjrDBzotNkxAV/VSuA1QI5IYGhZaFWwCu4nCfl/t0F
HZXmXx5IYDw6+JPnJJy4hbYz3FY7KMQhDkTLhwTM7Y7lBRACXgnczzp8C/YfT+NX
Dc4jCfT/RZ4wW+LwSJvmKh0ZsYLH7XSk3sdErSxDOqsdsxuAlY0+1auIpAuvqo20
ffDS6Bl9KsQJCx24vNKhFPAMMQ9OVG/aWfFhEv01oIfDMix1MALOL775AVjy489P
8MZPbqwn+cimKJ7lD5ouJGxzPQ6ewTGXy8ap69MGUoZZRvUS8qpsPzPSFsXAy/dm
rmoJg0oeePfyHDupnSbm/6uJr3A+k1N4hOJ2Ldg+7mXShxnDuI1HlNx46mG2nh5V
IJitbwCaha4mNvyHfVNbzZm8PlztUb+r+cnSBp8YvEwiqxn8YpA2g6Pi+bJBTICS
S0jhJ1irrZJIew5/vBblsDbLty1QT1XWFgDfrbwtqSO13oeiww2oJnzjtrvPBrGi
//bBwXWJlSDMHl3UZH73jwtAlaGInqIrSo1hUjDRWL/GnI1F5oAX7tKzDoUEpOB3
wwPIr3LyfcGf66HeN3j/hiif3lsuXh9lfOPFm0aisRBpxcb7yZXRdSibYzaiq+eU
eI2aPWVqnMEnfjuUz4Prd0ltY2WqSV7ol46mN3nT1rLJQdlktXva2tnh3LkIndgr
kmjudNQGi8O5OUMVeBQRSxdsf5SzunnJ+36lpaedqBOTa1wvfALgFcAnLV9/BTlX
HiOuDeIgaOltUY9kaecdbGjJyeVSKw9n1GIJuYOfpXS5fXpSeeZsy+QhKw+f06oN
Ui8VF6QHHnmmjvGapb9uQHsmfp5RSRmCee/Q8ibqFP/AM8V3mPsv5nAj74qfqdjy
qNR1lub5Iu97FcxKsqouOuuUurBeyauHVpvgM3RCcc7QV54rJpouBj1w/lw8FPm2
Ok7tZuyFMPVctxte0TEi5YAPVsxWg8Ktfjp87NHR7DWWNqZVQhoYd0U6+6UPv7n3
h3YFGwrnclmkq57oFgd3PJPKSFo8VpQU+ba3HhX3lg5iHammkin9MisZO6A7fDYk
vAhNhMW9N4vOU6fqCmQvYCRp7BL589nVVDEk9a5mb2byWTFKMi2Q05ftTpUwn2hp
IvG5DX4peElyYLp7iLZt3H0+0YTktsaDVTxJ3Bw33RlDSdOAs2FaljvvtSINSyME
yvDQ9BeqdfWf8Yaa3W+JJnjuayMZKr/7QZVdmlfzFA2HkGY9IaPzlBmAxH8/UQCU
fGiSdVqPLRaKVA+0tL4SnqvIs3MD9hTm7rqeM1NqZW7dAQjkQB/d3ASrMqBBhYrh
85qthi8nl7NNupkP37tkjA6GIQ8i6AvsiaTRpHbOQ6zb1bqgEc+WMu12bQMx6Dtw
l7KRNj3MwYuaMUwt6Tal8SfnKMeFM8yAQ4Nmlx210eawepcf2XednL0aVDba/c+5
nZspab9/p1TKgJo9VRxVN30gn80IiZipkcaxfIw8RizAiMS5H9rMtPvVIkZUEuE8
fEptydPJakhN3iBZRW/GElgLAW5HhiJHADr6phnHm1XOo4Oxbk+d07HcutHEY69s
bkqaEIGqQqVnObV/L1ko3OtF+tSc1Chj7UN8+kgbC4HfpXAjRqlih5g6UBnGEbZ1
kdwFn4BD7biFQWh4w9ntmBuCDbO9OpxmKUfc7XwTSP3ALFrZ0m0J5fu6P/2l00Be
YaKizM6pGCY30FYmBkiMlc1gUY7YiRFy7EOjqEcz8ZS2AzZS3R01OijIuFLyiTIe
QC72p5QGUbSFSX7uQjOjjgwdXTOFaZ3PYUbV7WrK19q3m6KBUzvC0P+EFY3GaFEa
NeG4BJabqKFfoce+CqlfDRaC4DxBDsnU8dFjcDevrQsPFQsqi0WcJ2aDOMuKM1Yq
bfEJe0MWBWbATYFGqz6Dx+5BJA8Ling6Z8kY2BuVwlY3C8UeBziR68/jt5prSB64
nde9LeUl2j56kMgbYsSsdxzGYLgw5fKN99Ezo2DNsTZmkXC4mLpyR9cSLUWAXt7X
zKgD1WynAHIiVWWEaI+VTz1d8dMPqCi5urPwM6VhaPIsq39GCiP+uWYMPklRIbNV
DAaD5DgjcL6IZLVKYsN92tCcFD8BJPNSNAFOqvMqQ3AffU3yXNmTWWBOy+2hxD+g
9I9ydelVU5YMxLkUETD1owKnMIFzHMPrBfBOK3WP8ARLM1wTKivNuothrwHGIG/p
5EWkeKZAw67KXjgRIk65IMPO2R6JvzIiLBuQSDSwJQV7Ny01uMCtMFKcfDdkktJs
NOmIJ1UPzUsHvyqXDusbUdnbXow3AR95uQyim6Kai/tuSHGk+b9/PCLsUSs/21JU
mdX2FYpOB/rtZ2LIoBujmh7mXcvFvt5oytkz/4sQUYSV9IYDDu0CM+zi47R7bfNj
/Zf9KNX2E5hp1vNYnNv5bcq/oBZJw/HzcX208NKKpTLXrTaYGqAl0xgqxCLtk6cw
O106xaEM/fOLhT1o1MbL8HXsE0YSvunm3JRazNKg8hEGPIPfC/H0nOJMR1CLN1Pt
hIM+fWkcLyBrvefM0WPAnbHxxAOynnuHiVRODIZBM2aMJQempXvwomsE+kJnRY+4
/CVMkZMSXxyqHRf9YnT9UrpRgt5mNPl254F5R2FT0jwB4L2u5QyfVFj86txWO1nA
G1IGvevgBgpy4HnzYtFtDuWsb9Sd+IbnYW0PEHfgTTyf37qGZet/XmlHfUydFe2C
Q7ySgf6gZGrG75BZsIPOqzDz7BHhlDIHsDF60GEvA7JVgzOibysiIZ+G4hVMaJHe
dsHVWQhZYSJQ6kn15yUn7mcw3wCFTPWWlJuvvg7pHyKygni4qN80kOHHRu7UM5ke
Uye/5Hu7ry8wwLKKk4bTBFj+SXCjCfneXBxV0tFheE/Os5cPLxNbrTA0P57aX3SM
LUwuJKJLqTlOuNkr7HeaF7uM/ZtDdV7x+HvSG7wR77vWrXJAwfqvMEci/lerBZ6P
IHqj+NAxWgxmKCWgqnjkt1U0Y9lm4s6Mq0bd1QzOBGWt1M5ZpH9fO3uyOxisd1W8
VRYKtjCJFsRSi7FOeeZNtntgiredxwGiuWvZBZk8sg/7pAXXIi8wxo4Kzu6EZI3R
YHw014PY2uNoUkZ3YGIT0/aSZqXR6k5Fb4mvMvCy6cnVaFc5LZVGiOd7KDOzOGJx
ArMlrI1K93x1+WNN7iX94jERk4A+T+yeIz9Uv9hUrKPUsjL3wgel3AdfvYZTDrxo
JYm9MwFzk3YUFoOMTJzWbXiMn6zqMbyihFU7ZAbwLPcaZBHB7GwkED8lVEFUXZOA
HGTp9OrW/SRshoi67S/bdxXltp1/vzz7xZA5RW8xIolLiiW2zkw5/m31Ew8aAXj9
DrrcRN7GPM0wELc/Dry7J96ypSwnexxAH7UG0ckBuWkLLeuZEFkBDDtH2F1fhRaG
LWV8BMLbMqMcGUoVFcUUwawJqxnYPS6NxmyBB91aywH8R77GN3ajydyNp+OkBa+U
9NuSaB7jWzVu6hLyt76A2jVmMYN8UJIlpAhEfgJ9mqdnUy8oCG6EQPsKXyzAZ/cf
spedCa1KSCm5jrsTfjC2/TIzI6ey7UM/Een3u4uaQmZzbyXhR7qT/o81mmD5QztT
aaQTdf+2IwfuHZTS/l1Fz8ZOzQz3rtdqNk28iVOfd/BSueAFKyvSWKDpGCa91BoT
vjRJ8xs7H9qxjJKVaxHNm18MnaIAULGAbrOj13sO+4O8/72+vd3P9TXJHxySOIr0
JCFADUZybetJeox2oYqMT2qrr78/GZsSnFuFEjyKmSpVTSCKunSgRcjUmNfoedMq
/UOrJb+ayl98wxjWDU444Dqr9eHBS05snTya43MduRqhUC+8f/oelqEPcPEU4EM/
knyikLZrrOhDdEUpO8HY7Z/i5yG9yKwKUluUshUjXviTFoDvGhJ44ClucCXgwBcA
oPKXKOVp6E3RX4eBJCpgH4yK8cmSUoxrmbbZzj/ZJHO2SoDvlGSZarZ+n3znNDjb
nhmfHIU33dc/uRvEYT2WIc7/kEZe43pXUqVnFW8yKPjDdo5ezdBlfOr4g8154jYi
BOLu9NYNyalJ5jRcoyLOQzMRmITakAZMI/7KHWyhVahSTXA+aRnvuO5gVLSz4lQ0
aYGzPHVDCZVReoKNzOCcd1p2pROtmCZ1cc05zTpzvmaHREDz573IPZyRAKFnBYgh
ex3YJIq/ZkPYWWKxIVH0WuidljPPtzoWYYw13O4NJ949gbSXIsdmKVLTLIafLr9/
thAoKijngxbz+CUKgAanLCUN59DM1vW0EVn4xGRWAXI7o3lG7hk3QcPwfi53WfCG
dvSofqoBYdEJwlHN17806iBWIPxbAaKXoTdHKQVrSyYzxclyr0kQpi6beOMv/dQB
N9XZB5nsnfTAfkITkiDsQnLwg87BgyuQqyY8m/DE6vKiupYa6UcvEEUSLR2CcLJ5
mFiiPHA9U0cdADEO0AGuk7777ATuJb2bbb6nfAFUK76Usysz/eEhZo2y5rkl4BRK
hZSXDhwhdzfJoz6Z+pw43dRcVRf4bItMZFYO2xcyyEkHR0V6PaWvHAXixZip68Zo
btznfN4ldLCCqttcK7rUumz0DAlkBMsYIFy+z4hoqoTH728/eJ0/UGKjOscr+ULa
I/WlYgyAvFbZJIcQFd2iRb3ITcvG6mdaZlqJoxW7nBr4RVEglhfydyA9kG43kinw
euaLNKOiP36q2ENEbR0dandLk+CIfMpANAlo2Rq3icKcur5TJguSHSwnfDFXXsuG
kUTzsWnQuYWmMBsz+b3etZ+8+TC4dLfWumpnCxvfmbuk9K1R696k1fqHd6zU4ZOH
wHeYgkURhy1whG1Jzz+bS9DmZOs8jknT0/lmk6U8AWxps1Xy3L1vl4K+gIoSF4QA
BQEoimd7iNg6oZeaIhoaqxGA7o1z0VW8lB2Ie5t0Ry7oNdL9qT4UKxjda0trvACo
Cyeszv8uVJejDYwJK4lHyw3kdIz+p2mzRbGInaUiMmDHelwPRMYPGWODYH+LDIca
cTZt7lVZPfecKGH6+LZa0WBwHeajYDR6+yCD1rs6abmw1AXyhkuHKa6FWu+3SHwM
YdWTSYtSYHekZDLE09UZmFN0UR2LJeji1AJgQcdsZdWOrBska/SCYkzICgvvZLem
HxEB888L1Te7MsV9f87CqFyyy+BBPYmE3+htk8UGe+r9hME4roM6nrTQak4751h6
iYKddNhiCkGdEuw1L7FX3B5oCorgM8qEbGfoDlCfMhQbnexUrLQ63Dg98Jr+ZaF0
YFTuyp+55n2xM4VTvoyhS/+J5ZNSPtpaWTd6fBs08w4NpdvCgdrS3s5CkyP2dIGJ
xhAE5vqSlI/C0qLAh9dyeS76JIlSXFjBn3STHMpERvSoPCpm0db+CQtAzJSxR4U0
wq5IOlTpkxPyUjl/NIiNltxcBI4L+Sz7V6hsCs30p2RTd/p24rNyCUSj94GtfIWZ
20jrC6PuNmiaVotuy7RTsGpYC3XAkg0vlA85miW9Skx+bjzOOLXx8K+9YMy8Cpo6
m2shzaD52+ffQR6abIpF+1a/Tw/74v1EzLjftKtQnlxMFdu9DHJY5p3MJK4GWf8P
xZxN/HaqfKH7tQSNpRco+WNGVmRlpu2mpvt0SmivMHNy9dOs58Z9YMW7ML+IYmqe
/scUxNE3A2Okrcz70k2SzetNPczQfdA2+dwyAMwlLu8icym+7zYwfu2xeJAnF+Wv
KKwwwgkPVrxsnCXUflLelWSolNmUDN3K+4nNMllw4wr0kKi4UVDWKR3EudeJrRcT
28VnSyaDIspH00+WbuIW2s+Xw8piKdu/iEbHCK3uztKSm8Lobh/oWf5detJVT0xy
IkIhtKJGh2N31b6PEPhCke3OKuocROXfl7IL9Fk3vgiIvxSvWUs02vD+58VVU09e
snid1y8emcndL7q2GsHf6LOtX9S6vyBrd6xtyz3HExGWsTIp7FECzNOOPKA9y5nj
yczHdv38ezF1kPiIPm0Io6gyesSzjakFNHZcLX7MvgCImQgnSNUE48GiYLH7WG/w
8nWlXt9gJ0SoCiqybSqzXMzqHNzMwU1G0swpx11OjbGxC9+FSGJF6JGVuhoROs0W
eLLJBBkCUi+0FLYvgCCv8ubwwKaLIQ7KOksGAeisnMRX3b9cK0R1D7ctIPdERn1/
rQL/QVEbi9tL6jl6TKHngqB+eAVjRtyDuIKyXt0iGfMVhcUOzTfNROxsAeU1bFRP
2KRgTBRRKN5aVM7cvofRWJIgvuUHZvQh39uORVpMhf9ZgxWhaqO8Yto4bGt+zyEX
aPS6do3onD50Ksn8UkFCVuWBrr9lM6NwSwKGfkevY5Qn/fWuZ/zJwAyQ+4r9+b3R
ID2OUc9Qy9PsoGKxtW+vmEH1BI2F7MwUq9xcnDrkWnZkv02cYXfS49jxEyt3qVjV
/Nu145fym6X3mdrW/95ECyISkGLSE8JKA7UbOZjZdxlnnNXf+tHUj/mg0AnaeG9V
IEWSxNAxeEqhMJ+LmLhc91jrzIs4vxr33lYVEy90Ev95CfIJvWM1ejTUfetXAe2A
h2MdJ3Fn0147eBaEFowRsxMSi6+hPk1K0M2GUOvXWlTBF4On+nZau4KIsWtpi9gC
Scb830p9ZcEJ4tHEawzB04UAbtA9dpFmUInyFlO91X48IQ1UlAAT1bboJY4HoD6b
ATd+hMO6NBvtFDMUATL5k3DHWwFU9ufZB+MTohq/YIHHss2L0Drz3qD1UEtSoMGj
k/wgb+tTqT7NyM2BRoSA74GcRTqWOB0U3NmcmxrGsPy+CCset2ABPjk8806VT0Dv
Vu5z2PsXuklir/0EQuRENrbq2h4xAZJdySa+nBF/nLJbu8Ud83NTIz9ZZFGEaDj0
/slDo9EQUIl1VUtMg5iihoo+ifr8alq2c2FCDH7tF7RqOXnrqMLarxcqzTDP5OeF
lLse67ApRg8MxBYqpbtX4F5aMNbKVUohEO3lCVlFxB8BJhQhGwlfLcxBQEheaQ9L
NQYPajEWlbauLVs0QXRmpomADB3cccUe7KSV473IYDCsKtXwCIi00ShXaaXW40XL
90qMlua9Gchzd92pe5rslPWc/LaYNTZIWOt09TGwrfIQKfooylyAGJMs0c/VPexT
J86PNJQ527jblTvMQRc3k3/uavLasohpMOQABrLGRbCXbbhKH8ukOr/+oJZm0h7w
iJz/Vt/Fjvk5wi97iMcEDU5p1z4kSLeTtMn1mmOrZfaBdoRin9RKQ4MyfAoI7uXX
oxz7nbBch+XB+90Vpygj+sDzloY3RX/c6DvixddXvD5RnxFwLU7e/vgMssh8hk76
EBpSWT2az4nzx6Nj67EtD0aV8nb0u9o9CKKPDwn1CfAxCQBeE6P3qK66i3YMZ1zI
tIDmgf0DSx9MGYTYNWLhSc5OVCRaJL1XNIaQqJsjLVZbri9TB45m12vzo63H+uL8
dWySMILSzE+dcVn3+1NmBjg4DARxYF5DH/lzD2uVaHTO46ypC++Z174AavnFnJAV
xbodaZc9Elcf6otLrOyfpx7r9t2tsBnDKWJS7SjraQWIBu6bgWE0n7OGxdN06Mb2
2uDpi/yM+nTL8uF8Shdfzk8lROpQfdpe/IS6Yr4Le+tfOkFqPfw2fYHBmyMTNeb5
E9F2fj/H5q9Q2edLWQ7yP74MjSz2Y5WVhLi1ojIKHiHMpwpSU/kTxDErcFPhhizn
AnEawJq5ItI9/HX476fnT/3VgnWktR95goLgaSunpRyBOchOFsYZ75lpRIKf/ZV8
TwH8Ow/s5vLdYutTQbahAGR6bF9slQCNYtRL5ZWCkbrjWq+gNHaGNJ5Dlp7j4/bH
FPV6Gij1spw/ITXzqSL/tUErWqqVVgqetT82W5dwwT22QYw6fpvEF/PHcnw2OuV0
jCiElD5B4IMM0tv2OI7dOYWDrW5AQawW15TliReunY92BFfbxyLTlEwoSjP6fr0J
9Mr/w++b/pi+xH+tlrW7phwiYXYlLpoRmQZSXyl+DgaDzummrLU6H1i6lYxKKf//
jYYGX5wsP2AIpHbS7OishvporE7LEsAMlfXljhTl646Rsuovn96Jph+vY9hb4bET
XiKZHtITuypFk9ADZnZ3odN61LXwI1j/5TMzc9THzJa34qoL8juuk+jL5Q9zjSIC
EWKQIXF0FKRLJfxyj+8Dzls5xAY+WbqBxIf9PVaupUra2d9iUruGiLGSE4W1JQlU
/v3885MC2/8sd9cYKBe2Ye3tvYdhsU0tagYlEJ/ghRQwB5Xru3PqILUwKNKKqwS5
Yb1bgkzDLJuEn4F7B3dW2PcrFVAuWYrTpIzk6sJFcmcZgrrtHfDJRR+kQw+mzYsV
G6zvyze1HUbS+ZNeAJJgzLys6rB+kaXLrTv+kSTQabCQJ0g+XVDeid8virU3zdjg
UeqS8KzFpdFApcVU/s30zMbQj+HX4WlnUAAi5cou0gm1Hw6OA4LRSmO6HMzHEl0r
85GAglecQk0CVRDorwfZ7O4oMG4b8WNWedRFdA+tzpo97YEY4dCrHbnC6jbLcXVb
VaCt5Lew//NYZNiCovI73+tcqNN1eamE+DcjEhOOft3WKvX8aUzeHA+G0E1NgTH6
Ht7DErW5niHLSOSmZjP/ivYoUc2r0HSVySzKtX7fF9lfv4eQKqkSUdiuv5N2zxq6
L8aJ16KLF0Qzw+vsujPAFqOMR7oQuds8rVBVikeGJ56E9jsrnZWpWkWbJOwqEClM
zmO+jtGhKcp4ze+OLEcyJpEVwYN3j4HKYG0rR8/ZCrsJd2UhK5UjwooCQCUNDZfv
RtyM9kWqehNrx6jCe+HEbPLYzm4PgQzedzvmlOYpCauNVewt1zT/UFe9SABYVnGE
pkNiIkHARTNjcs7svQHq8cEAClL6xAdowdV6zc5eeQKcFEzucak1sTlsOGqxRaOC
eQWzvdmWhhPmDUKFeA9rZiU/z2izHp49V4CuGG8+gmRz+llczZoebHFhWYfRUpqy
WvwnIfPU6O6AVZDeBW4Pp2ohBZq7Cq5aiJFnrKuJmc5BXVUDNup56Gab8JPMKqr2
CUZiixm51F+oxqC8tz6fF5MWcERY0G6uBCu7Ciov8D1SBdaNfFnJDUVWkj9aoXqk
eu+xPNgoM000hvDHmY0ude1aCqppJ0Q+Bzsmns8bRlFYU6ppz+3fTbX9WLMFMEBK
bF8JPJQvzHVp2Kws+OBwXTOKSMPnZZOWp86+lkdT3QuiyNqREhSEMMSZK4bJHmPk
38zrC3EtgYO+Kvj03Qgz+m+wgBavgD3R40FXOD+gkLSNVZET9lVRnOlUOYUqOIfr
fsXJHlH8swZyknr4E5bFYmX+ZONpr78g3ozPXz4SUE7gOS/EyNX+/AISnsXFGZ9E
yoaYtgEHOs55kR5ZiVERkUmBzvTsFlOMjH+kv6IeOtJGlh98IQPPnQJuk0EizXya
x1Bu+EOGYp2kM7TCZ88VPfbCfDHjWX2FbRh8nMOJriqJQK0gJRKnyBAf+5PjU77P
lLzMljW/JBFt/tK1ITAobKQInGOo4hWVj9M54TqHi1O75FJ6vIict2KUs1Vc7Hsz
hPH6etI3goSRs4a27AAqmgXKCRzAsmMdtJ1kKTMgFGKhKe7ywEUHQe4MgALWh5ho
Cmm+6p2S9IDQTQhUJ88O9LTr1QaTyuD+L7PvJ6LG+LqZZ8VFYno6uvgE7DTH4RSR
HKOuRxdt1wmyi5CznF2DjI2Qx+SkuHqDBVdMQjSTMXCqbvgaJ0iO575EcxVfIzwq
6ylF+ebuxVggAkv/vQMKdRNS/V96Fa0tx0q20KgnhrQZFEJlKtMDVdUmQLVIMRqH
wqHPpsNtcUMqDiF4pgeLmd4d1URuH9OB/e+xTjNvD2hWfsRLybyGQIHxSnm9ryYm
Eq6565vtEp6TXqik2hbiqm1bE02gByqmYIdqaGE+vaUExzbLfUsy1CzGHOaFbpXu
F9pRH4MGZbBD9Mc5/IaHbuhFKbMGZk6S+oqgXTxKGs8nXDXzn+bLo6nyFLnt252W
ls6IamPsPrp7ZmqV1A1ZwK9QTs9eDq/JxB9p70uaVTGjSTbH0d6MRXXwt5bXmKQD
EPCJagTT/j+XtvFG7T3TN5+hvCG5LMdyZwD2x9DS2EdAthN93155ddscd1rhvoOW
nvgc/RgrsGRBZ92NW29mD5gV4eev2hrgnTxh38IeuqjHVC3ow+1y+Wc/0vyaeMXl
qpEoOm+6GAIACMHY9dCyMYF/Ox8zRm0HuSsqTbIw4XVePaJ9V0+wiYms1q94wnCF
myeCok8ULns5IO4zc0qdN9PxUeH814aQT40GIHuZHUik/JeMpm7n+NKPbuzVHQPE
PMsVC3DibK/Qsq92d9ixOZ8hsjq/ym725gG+SVUho9NzXWbaL1O1MtWEYilVFVtP
ZRzn9iSlQXvcj74CYaFxhmYGC5R7YSFrQkzp93SVYqRStL7zS68aKDaRHPVIsiLL
ZvmvycNC0nSOJ4wtWxpTX0Oqx8jqhazCcYmbcFxvdeWit7MDTYQzjEvnNqrlscpi
Yl8JWaeCrbGD5C9JsYH7GT32tBpJQmwlpvJHWCid84cukbKeQ+Wtxt88xahb1lyv
pOee4QlAKyjaVihqee5HTQTjgauc5l3ABpl4bkaTV2bHNkdsKV3LHFR/0b0qtffr
OQtUuFnGCPKhQ3YLGoRlUO+er8xXkmHk1ukcKYzSagCO4ZJeb3Ag0YiNjeJ4qFou
YdmByIKnPE3HzX635pxM/AafiQj/XQkLoFGCgDdILURdYD8IADe6kRP8Ce27koSf
5OqPhiHFkyTrgFGIOG+jg8p5F/vxQe5cCwY1KPXhKFCnuwZ8ecbKxyUjrfMmXend
SUfAuFInK8ip43lzg3oSF5+wAO8OezU8oiGHX7pCzPZBO5dQq8qI/wkjhnkQB5wM
wNrZr4JfJvLvZ6CIkZeQCYG98OzSBqrTwle1Q0nBytzyZMoL7hiCvJcTgrLcl66Z
/gXPgXic4hg8PIBwdjGe3BBHNzAgYfGAogFW/ZQb45YdsZOrAEwVa/jfIbiITEoO
WQiHfdbQEeQ0OWm1MZOPzg6mDKF0PyEBeUZOSMGh5K89VlKEMnMjPEpGAT2X4cSJ
rQC3a1lBPplHovVuYinmZt89OcAK6jBlqABDvx0VCwa9rJYbU/2myJJxWhBJ5AQJ
TZ22a1QxGJn7xJGXDO+gQNbIuhm9iYU5HLhz+2PDGQy/G13VhgU+/1wL/o2uABbx
jNPw0qRbTuJiPVN1+a8Ux/A7/Cv6FWA+mzT1NQxcyjPX4QUJPwdAfjby5ZvNi1gg
ATPbxfsIWnO5+R9SzO3xIlX5d92pJlbmMm+nkvRunD/cI+1A+fF7Y5EosOME36fU
o2L3I9DS5CPIQt8Hq2LOKIGh+UV+aNvYt6PTsAaqzIIgkO20ERxznQ8VCqWEZ3hT
cletO4TqhdB5CXF4yjptUHltg07rtWrzMvXUsT27jSOkw8ymV1lv80g80ZA7hKen
4NMwe+5v6MCdEqwTyDM8/nvhiokt5KVJWldkhE2MF8L9tkwcMKT7SAol/OKPIfEw
4AZAOzLhZ0JpMb8KnDM9j2Oh3epMOKgEpKuJdV0VoYDlf4jgKsqNZ6+7EJSDcqxc
csEldFfEZ+SKVpW79q0+GB+b0+AO1pn4tihPTrWZKmMEefCyrgS2QYcC95v28R9I
wXAC10anBN416WeBk8OmmFQq5odQVadjhgCLRoWBfToHqwuH9K6J98EXLgiA/Ax0
CcDNQWAK1kkG15bX5VZKMlM8DUGYUKEs6FGjrpGkyn3zFwW/6e2LZE4hv8yPkSLl
D3kbQ4lAnzF+iT03xMC1iDz4GFHjxJzNx6G3dulwgRScehlpTNOCTK5XwnHqx9Bl
JSjlaXdZn5D15T/gmYSUpTUplFf6bbge4NzvF3gT3hyYI+vTIgsnRFkv7v5zJXG9
lOAjqnV5C2irrRMv2w/vJ32RoICDmslwQX/Q7Nqqtya+6mTk1Hbhs7X6FFeZ8pJb
PJW7T5m/alGay7LDpu/Vd1FmWayrOglUtZhU1/asO4XxlKVc3xJLiazyg73XfRkK
k6tXnYlZtoVtyUWfLs+Vc1BpipWnp2i+qZcY1AIHg53AaMmERLFRzXHHf/XkSOl8
7CXB7iZ0x2Kuw7tmgLACjYhWwgHMYsqHtxNSgvFK4ytfDwuUpx/XKJ6TgikhZCkF
BD9ORWOzyuo48YrNq4y8/2dvl8G+TqK5Je6iDRAvdGC8c6CiRXutV1MMi/xicNfC
t9g4fo3El/J6mnLGgtT5rd6MtaW0xqSdSEhCCM/rNpV3y2xINCWDO9KBJQP9OKsP
Y/T9Q7q8m5vNs9Qs4f1cBY4txUMEyYP4V9XlTvMRtjY4rOIA98hlCN+HNR6cpCiU
CKr4afTMOHapfwIYYiHeY2ovivOUJpYDynHj025NJCRbkS8YkMEQTSd0uwy4yPN2
o3uucKm1S2Bt9QamHVd9q1dGsQonEL+Q0I1TPErF1fbfmHONPxtC36wCYW7dao8L
G1EtH3NDO/BrB2HHh0XIlWW0KhdfTDcJGm7q1CGfFqBrbLNihKlZC2L8ja4UqJm5
XetOsEjJ+H6waE4hq8oBGNG0Mk5IMkUbF4Bn9yNZKbmcSx5IsttHN3cBbTumzXCA
NXyBChAXvWu7x8EV31X6fFPEQdGtIgY7zcJQ0P7nHJXM9xYAjl7M0tf221PKtpJV
8tuST+VAvTe2ij6uus1RHzDWLRUS76yTZAeBpdiRJMSy8bMlnLVevPeYTUcMoApy
Bo/z2/ORIpxpNaVoN7tmKErNfCjYxT2vimvE6WYc6GUx4cMms/JUmO0dYNfmYdPh
As71Yh3ctrZ9nn2cHVntaXhd+XlFNTwlnyTw2ue0PC15IMnpQa0YCSAdNwEUbTKu
2RF037df98C/BmUwF4opsETRwSN37uItd02cYhTWxcY2kItpLpMbtSMbH3dS/9IN
uY0kYMT1eJ5cu+vpG04svBgDVgXxum7yYVw/R4V5USKjpTj+ajptNhhXyRpHa/3I
E/ir30JQqn5SAQiCsbU8m7KjowECbYqPq3tjGI+kii50emhmrWX/BPRLPZE/ys9U
DQNwgmw9k1aXCDIf+ALbbEpTlSUlZ4NiCWfot9ovZko4aitpZqtf0gBJvzlxDKGh
uXcWfpfEdaVCDDb9D7WFAlvIarb65sIIyYkUB1vKiddlMaEgeat1riLHmWofEVQS
KZDoC/eMvj4gpthQClnUzH8H4WSOdmivSBls1FQcbnAY/o9fkbyNl1WlE4Ch0sSY
qqImgisNj+5FlIXC5wc2hZ0IUUb0nmneOTPJ4SZwMP9TaKWHrq0ALZK3lvv7tDMf
Xi4XWMKis0IBClWOgLyLCcTKlHJcMlmfH+ONXMC5al20sBdqBTMpmVpOSKRfGcDD
jgfJukpIqIWqolYDwonEW4M8xssMrfo12FrOFFHq+mfpHXkQECHCgaYpZq4TQWXy
MF08vjY5gdSvVJX7w/GE6JBZDmVeV6L7EHEGErc21REljAFAGP4ru9+eMkAUGPsN
qHY17rRJDvv0zjBn8qb3K4mn+tWkbdg7mPUdiuBIYZqPIWMNs2JIZ1vNEFYT938L
RlFZ1WOleSq7mKCVURMBIstw/9bRaWI5ujxkRxkW5JQUCa9fJtuAcHEUNBdKDGTX
7TkMon4qa5LtBgmLw3OCWi+iSIsowuJc5lMPYMT76a3LDaw+WGXm1yxY634MAqEL
ljLY12lNVwYRc7OapIv5MtolgtInJK3U029eN+6hJKrtDg3Dke5XExfQpJ7JdnYR
3pbYeLnnQ2dn30/mkZ9ATwNdxjsRVtjNNCV6ZD0sWZqDUzFVHn2YG3pxiUOf+wTQ
1IJp0V/wV0YRzD/iB9GCqr9BvB8aP0v4q6nWjfBMSgiwJ0+j2KpH8cCJHEbwYrAv
lqmWhfVM87PRHLDDaxP0eQR3wssoK5nW+pwHyRWvLo6162vEj/iPMxlJ/DQAj1xF
5n3OIGVw2yPeMeHXWIFEwT06QPvZja+tGdw6Hd8lyz8DYCSlss4VvJAIMBJNGjom
kwgT+a+0qjmJwlzOpeHaMJaCi0fT7OLb1thromWIZJfvHh39u12X8PoqV9tlr8v3
79epXgV8mQj0CNnmvL75jge/ExFwQaN/Mz+4n4475HXjO4ALCpn2Xpyj/M3kdHka
ohnW+LWH5FWukyoB6i8N4SlMa4fI/CdA687fE+KrvM0EwQhVGIwWs7LYVJ3IW8eK
wTvvw2orewqEa45zyXqaUvFzZ3B1sbGdUBSuhBmNDoV4fMEJ+86uHEPWqkBGSJEy
dT5bFMOQ9deL5gC1dg7oEHKApoBo3188lqLClEuGqrdoBYR+yi1s0sWKwvkLwLmI
//FZhPktAbdKTRD0DM1WLYys72ML6dwgaZmKSXwVW987ZtnelV1YDSiYO6Xxcc04
50rMF6dLz5Dc63qn8vmwzs2ce3xhwTIb6qQN5jUxYUzwFhGLAlLGIw3dm01zzFfS
Bm9tLa+nhlrzy6NlHYW1KnzY5gFkrbp67IHWdryOf4pN6YXO/nKeLUaBpew1s0F+
c+SDAyj8zBKIt1t9knZtyKFFga58YBMMVcYGEZ+puBI8X5DnXxzGf2j5l1Pbxw4T
QzSjqlVHutG4fmFmHwp+ZwfdHLarggYwGAJjYIIIfdScCsBymih825jvdoXG4PjG
/rgajEJv5fofRJ5q4VqaXEOHhaSfYU70NhaVUfAFDGhv13hgiTqxBKR039AUNuKn
9sQSIs9D8jLWwE+hDnyyodNHwqMGzUQ/jktnCZA1oHZ0zSS5ggoG33yB82OWF/xg
v2FRel3mKIYgWg9PvFNxYWQHpe4DIa/+h/n5uzgSYfk1+HpO1LDvf1lvpu0m2GNn
O/XHjsXHZNzVFOKWMNwdEPatQL/KlwfQwSVeecQ5MsZAQlEg7LI0pSElIR9aQcOI
hPO7lcNGPaiyIJ2ZAE7zlWz7o5gE6NtnXFbDMxYcZ3vRk/H/r9kZU6f0wz9jY6JI
3NTR7D5fXjuJxohyzZ96CG6LszPurGFStXE/8M/8ABhgH1fi0cAon0WGKLA9rQsh
+fHj0rxbA1/GlIbtvqycsncPRUTh/svIr+NaiqR/DX2jrNajHDEsvz9pFfixb/V5
IBD7443XlHvITRh08/a1e8gicSxSYcT/cKA5nvUYNiY5cje/W7GP0UmGr6nfr1EK
Sas556q0oM5omWxsN8VetX/p5STsLpwjf5UjH8vZ+XhM25ZjZsCc5GLqYj9JjYGP
WIMsK0QaJ2+gjAAqTajYpfalKfTkzCpdN5K/G8R614IrrE8SHB562vfHGB0zDqrR
uPY2dK9PN1M93pV/bqLb1WLtl59gYLAUgee5Vi/jRNimgMq45z/g5fDbuK6sbNpO
GJ8TXoEwRG9EeS0ZCzBKMHkfUcJ2TeNy96ug12RUbpIm40sQs5bx7XgudGxogD/e
zV8sPoPzQ2nm6XUZSXc8ldwRj32SjZQ3OM2aIMkRWiYp7SZb6+DwsqhwuDn+0Tp5
JyGdwsZyljWYWHUDgAmAkIsLr5qzYnPNS2qEZ7AyrkOR0H3Xxp2IEA12ukafxS4Y
cpBn2G3G8tXEJkZ8MBQ3kkLLbcNtqR8nu0gHfImxZEuCDoyRn+WE0BCwx1iYsBIf
nPcr3gXVBwwDk15eFyPB0OvFqFCTJEgh2X52KEne8PFtSbY61UnLkvzyqJ2rcL/n
bJYgqNA9IupQ2+S6FKGiQ96VvZIwlfL0C8pOqF3hTv0Qqssm7kPP8wQaH4Gydi9P
2uUn8nXrrWFuZ/iI6pB6MSuj+2uWkFvEWp4j2HPBm15EhXPCFqtpajvZypqXfy0J
IxujSp4xO35+qs6PK73oXKhTEH+nuuNl38HyqYI4kfQ8vA+312aH54Au6RZtGO0/
nwFRUROL7H7lpBVxZ1piwAeI2sN1bpEYUkxfP44JU8h3iKsWJfN+AvIcmGuwHkz4
iTsImn0eo8jSeGZqVZe1pr8QGpPDn+2PJX8zm0hp8D7fUZ9gfNRuPkq/NOSmLqJz
76a05vUJw1mmWCoh7Ld9sJPQHCeJn+dgeUfXDjLn2fimrZAAhfn26yRoFLnHV/zQ
HWA41SzA7PiqFUkzuAeSa2I2pUcUqKkP1kD8kU06gfZShjBJXloyh7z7r/+r/aMt
GPGxWn3/ewzQjZ/J6iASyynf6A3vRRl+j6hyghMkS/L7hJmtZ6/9CMn6yP1loNRQ
Fn+sByqkBiXALkaa2/nTofddCKjNTqmVckYOgfz4Q9y+ZckMo+qe4w/IGxwnNHC9
WqHXInrht2AYh4DsJWshh1Y4xs2kw/GEliLAS9C/WQ0zZEH9fI4z2GA90vXNG059
UKxU50jnRdqqzVPtuFnobR/2Nv4iotItvHnuXoVEyhAWBJIuHMX4W6Bw85eXMU8y
tuWKM8OXwlfp7lFii1je6IsLsWiEpzo+y9bMpko7XcZCgdQZQhSgAFDnJIj8ici5
U31vvmF+Hsw+IXSzTuhb50tbeV8SFo72/UnW+faDRyMd77rsi4ogN3sqAhCPJZ3z
YLWzlOoDiNFwTEIsZoSRgNhYnJ0096Hx9comrLsC0ujH80Ae2M3nBRRTovbL5e2F
vJavR2NEAcmqARtbAJX1RciRuEWSAZnp7Axv/iHwCxaU5vfol2EraCwvPgXxLfuN
yKCkfXj2sux6sWZCs4x46k2GfklEh0sLfm4bX5c5cUnKTyAhkneJmY64qrT0tPDr
QS/uPV5r1fmVhgv5/cXEDMI/j9XWBLTMnrPkVF01QmDmbCjVg1PbsrewDDwdygIb
4nTvDZfMGriZUyncEANitfkIFMTcTx1CklQS7dksSLnMCEaZlvbywNGIZ2yyY6o8
LcOv3sJCfQkMN0veTo+4wQakU0PTEPRBWf6MBI4zqBKo914CgBee/nFJlvlQeTE3
HX8gWlfxjuIjKWOMglyH+cKFh1875L3UZLlnXD6Qe+MsW/bdk2Eil0TR/8MrkTZE
4w3f+oHnutRD+qFsCPw7xBa9ubp59Lfv0Bj+pzO5aiM2bjjao0CDI3w2OqDBLxfb
kTLt47L2lgoWUxd3Z+aWivY3uHCZhE6CnYhU+1QHhd7YXQJrqUiyLp3Gy70qjnZ3
wKojvSbQjOzQFKt8NBfHk9jVGKHlU4NyKitw4oRNeWFo7jAhWvNREFmZgIb8R9IF
JjpPu2MEzWvB2Ay3FMImJ1zW6R6/Cq06QnSyG3zL2n5C25WF4aDKYPodTcPif++q
RlKpO6ur+Vn4sq+kTY27y/R4CZe6TKEsDknjYSFc8MCzBvn6Cbtz4/q4pNU4j0Jh
7f0a60TorU9T5u1io7efeeppxBb2HZH6XoJ3CVtlZR1BPfH1/FkDPiKbVV0uT9pU
d6CUomvEchY62Yv8dmLHoWwSQrgyxD8jckXZZR3xjmcDoc0B5+25a8KfnETe0tGK
1nZdr5EvIJ9USpK/CPDn2U0pChXwv9Z0Pmy31q00Gmf5jnw9Obn+bZX9bgMOvkKR
pEPswyR1MF7IrXPIYjgTzJzpFm1I82oLORoThNZyVltiW7IsqIDb2D5h5cag/eJU
KPDjgypzlTx5q2en81grM2FMRUR3cKz91WdIrJ+Y4zBnrXwVkeG1knz6f2GRfB+Z
n0w+URLufP1YNkHCzshKZWUegyTYN+Q5/dgo3LcpydwLI5qamnHzuUl4rWOjNW92
QujCsjI0u629vEkN/EuXehvQekDazf/BSqVvKF43OsyQx331ClSx+hwCWFd7ahBu
QNsahAnIOtj7jVvuh5wSO5Ar9ardj4fA5hJoFbsBuEH3tPUPpwqafvFtjG+yPFOM
qn5OLYLAAnSFfjw4naILuvqkPUKxPd/+g1NOcO3ekdPwuSPP3kpooP28NSTkZyTl
M8HGaSBDomZLbZfLFlrU3UY+VkDDRdg0XgHHQAsPjdoREClFPVH1kuJBoggLcnOr
gHDWyju9dhDKUXoZb6PI/5Kri0OtE62u4L46Lmiupg3ah316kTO/l0QUbCeatgc7
2+MXp1eLgHbd+tmTPmPjb45XTLRFQgPQZaNc56fo4huoCyGoKPQZVJs6El/KMHZY
vinrQDSXnvL+j21eMp0O8eJCBbl/YXsnbdLqN6ioQjeFwTArE4WMjT76nBAGJVQm
NvWmGWfJ2s1lQ3AHE+JuvKxQ00stnhZerxL9PAR4JWkDKKihBpQqfFKwvv0uk3eD
bKOKLiYYHklnnZbbDn/JE0KF/BacGVzztPGKVueTApq669JGcbes11/uYMB02C/s
eyYjXvHpqGiCOPpr7HfVsdkx9uNGj7K9Mv2R6XWpfZbW2Bc25rbwW1lIVt8vznyX
WvuWCsqwVI5ANmi2SY7gk+hjBmk3ThjsPQHrl3CHpTqzHWzyGYiV9EIqyGqbtosC
hWK9J9l9w7h7C0XEVDYo7Jiiail4LkgtVdkR+WsZIQOa01RJO24e2ro+nWULGlyX
nPXZCwzNNoH6w+y39SkphBOvAQjxS1N3k1lLZZAwBPZWU+V2rA27etYeMkrTBGqM
HZg26Moq9kyOG/hyKGjsc3/OVqKgYd/T2C+1e8B2wCeiHtlrMauLsn2XfggZBzkQ
HpddjsuNNCdLtSqP8VCc5yp4N0oHlrCHwHm10v3ohYsNR3ur1Owdv3hex1t5eAdd
8C0Ru4NM5ccDMMwkW/zKpukYTM8vgu3Dob2SCVSRg4z8lG578D5sAOSPa8pCpnVE
U341Ec6XlyYCHTn7QPF4rumGhgH+iDe5LP/jDRj+qwKs63bISpH1vZaIw7f9i+nG
aj/puDDdAHdH1x0rRKcgBr9n6538Z2XIqUYiioVuttZgappOfTWpYT8U9MTIhZjg
IuJkpGBl0t+cTzoCz0z7XqDiu/AGn85VhCz0bUqlu5iK2pj1+yuyF9GI/GyT0k0H
+zClaThrQpTFAT6RH4UioS469hO/HtaT1c4vBHk3yuEhZdFaIvmINZ0xuFmyfwde
EUfENqzQmqQArFLz15l9S17ipYVsk62aiD39Cw15XPAeRKTwRlV63FNwfXDzoCtN
wzP8C/0ffRx0nzk/aEHLJJNbxFVxn2ZoTLP5b9uwnmzYohjuYk8UkdtEAsh96ynJ
GhA96cfULF1vh86zJNtrwOAL9z8EHNorq1kCWByktxhipBOC0bM1kui5B60vIvkE
eijhgkDfnEo7luxmfw+U6PeJzTJ9yMCjxNgjx+jYUbQeAzl4WfVQeugsgYzTFEVv
+ImdmLeegb/xXJAi3x37JTg/j68OaT3W2imysIINjaPwpefB5KK2nURNElVksHGo
Io3h+XIvQLTLCMpJYDghGHmn0KTAc9+8C8KG9ilRZx1zoObA7mpuZe8+8SBlLWCs
5VJ65WJWj2C1QZNz9v1JnwRFix0sOjFNHDu4zf8l2W2Y+2n3cJAd8BV0RHPgpGWe
f4D2K8gnGInGr0EWdv+VaFJC+equYGqP3uyrNK6RzpfEhPPoqZFf5LAvLN7n89Yv
+Cr9W+NJ0S8djvpunsFmLiT7QdZXmDAcRTK0ytdraymEArvOc1qM/1TbdyxF+4ZD
z0nNdK7YNhzjkNExIEnCDJbDiGZ8RHifenQopI9JTWpV8CiFeD6OOkPo8LWgodxV
nVzWwZij0WnE9ibHDHRUb5dNludg/kHYRaE0B4aEO/7eN4sVzg/QKoV6hY34iCK5
lxegnsth0JoKnOL7mz95pDVjFXvj2UzYY3Gm3+YfMY4IhzZ2Zac1b64wXed2I8/2
r70AYCwtyF4ALWftZnXDbmqVnMpUav8evGL6FdWVklrHqI/wIk9hhzTI3BGjRDc7
HISsli74UPqD3Djht2sqLTkIuUFYSVHwQoWPtpdpHM1KlxQR/DcjGwAmVpkIibxv
MHy+3nVZJbr7v6V+nATTesLAzI/QgzhRb2RTSc4U3YFe8vI2BGBQsE8BGX21ihHq
MIdDNy2eZwoqEl9wd1gNK2Rry9LDLvbJRp6uABJrgh9Ng/22gYHRRckAuC//smdR
fjbXj+C4IaDTCNy+kXkU4dvn9ov8H05KfbZylg1p31zkNmhhHppHqdX+ldkQaWSb
ilD/EC9Ji9zW34z8MSTOx68M545U/zYGf/MRfT9k7OteBJsIJPXh9osMjB3+hS0A
RQQmAdDCj68b/DGkF1eeYWVzlNxxHBQG5xgeRppZcWGiqYXJQlZ9tRs9WJQVlOOV
HAnUwt/RSMPzj8DWsKj7alraR95CJIyNakWPNqLGnlwBbilCqtH10v8WJzkMkBHd
Sdfx7bjW4Y/mjKMR7cKuhhQuoObVS1ECoymq20Vvs6PltMphr6wP2Bt+HHWtfnFa
ZOTTkQ3dliLUOUoI4rFt3hCUOKzrK+gc2pXWFcaBMQAok0HS1/8K/IiMeiPNWWQd
dy2lAvLwobM3cSj/PXRFo+Tes798fyBxJh0dPklbweShIq2DwLBh1Z6Bf3k3wk7N
Gw7r4RwSt+S4X9HDezp2bVsxma6GQrKdwDhO7JbRBgvPeaXIn5pkSf+p7umg7JTR
1flRygNPLsKzR2VVrfwi6qC5mAa1EgM2ufDFNMzYc/wRJwdwQV75oQ0iMF+zXSEQ
xlsXsdkihPq91tbjkBTVrKCYFWAvxr6K6hVIsB30njaJWeWHoVlLXPk/wX0DwPtm
QLOnE+wpu3Je0xC0JiUjkZIX8t1MFZSBABUIGczkfT/PXDEAVPfKDXjyk5JjGZMY
Po3V5cyTJ5JI4K7sJtGE05dy79orzL5lEvTgx3BFUbF8zP7mQeWE/y+vhdgy4hQP
qUdZHyNqTMGTBgYoDQ2WEOatAHMhUjO9iN8/0Q3yKPa1ZwCxv9fvuHs7iH1aHbXf
pN7Q850qw+FFNJC2Vakw9Y25R8+IFTxKsiZ/O4SL061jbOGPm8vORdfvU7xwqcd7
u0rWbUjwGIWtADvEh0VZi4PlFNn/1WptkgaejM+U2XuC2GUfUdiFHlfwn739hZcJ
AbvLNEw2VG4WOSA1+ojRVGM22589Sl6zoXU9ez9t3sheZqpPOqkxpUqhMFTIcjDG
7iqX8TAIOilqQyc31/Tc5QxQ4GzgdRwI1nUe5LFaX1rtkDLZz53TrcZpH6qKfmmO
RNX+9jZhy5VnNzevCybx21S7KgNk7Z+wDizRFEHGfDUvLiRuan62AulkuR9pS/iP
j0d9C2AzMqsJdia21/D+AbQBDVwonyib0m95RZ9dCavQ9BREBXmhWVW0dReHaD64
UQnExAEOy12vhp9p7YdZ+ed/CMbEqtCso9d/XpFdYJppNA/Ikmmpk9Vs5zXwYKIL
XFHySWKrkBTcClTEk62byp9kw42KrzTAszYIDWrKNBoUAaUKM+kjYSbnFaTwjeZF
+ARwXzUOBo9+KQV+RsUkWHSb+eoroX5kidDAk29GQjBf/INH649/KFAzSGINQ6gU
buj065aog1i1+Ggrps8kWtfdYzwFowozt8HhM5/P1rVNgBhipE/G8068rklDYmFB
ffEXlGhqNozmqJ8RCzU6M3i7xi/wau7KbVRSRoNLajzazDMoQ8p0VHvaR+S/xmov
jHbezPQbJnf28qVlHYs548GzB7wfEbklN7drXLRFVirSYafs5mYuYuIJ7g2W+aQH
XuRdWfJy2kiOzlbdUT1wGTYHXXTKp0GmSsazETY89kzPM3DDLpnHr+U445799WEE
75TmNe+oThD9o4MyuI5c2k2ZH3AduM0osY0PnOwSGUyUE+qLMhV52Skpc8gkm+ey
daGzMsVeRBk3f4pRTRtDZhO+1pexgtbdEj/0uZnyoz9WspCI+74aqguVk3joFZN4
bzkAOaRkM7lc5LV/ucGwGffJubnrX4xLzNrLCn+5Sjdjpis5DmiFU0jcdb70pyZV
1gFyYjdVLGIhZzYTgFOr7i/+V5N/EORp7ihHoz3WbN9PPIG6/5mR2yGwhPUKh9xj
3kMmvGPPJHTIgrsD9O/Irhq5vY2Cgjji/wRvFm6nz7kS0Vo06WLBdZHkoIWiZwWH
25UwYnP1YDvGzsOJ4O3di0EdQ+jsA84IrBkGm08xUsn0oz1BDvPH+7HGPap23TGw
cWbecCOO8VDYaDYdobYDneuiwoZNARJYbkEVDAvBaDbmn2KoEUDeQ+Wep8YNmRig
It15Ytr88+iyTRS77w0Z6NRDc2zCZGXDupfkW+TZHiJZn01YEaYh4QfdjqyB+VOe
J9dWklhqwoljysae2TynqkI5T+EwcyVcEWy2zFJNJrK+dpq4dWdWkumXxnF7UvhO
WpPd8HDaop0VEBlKklP16GL55NCBmTVbw1vaww+AP3viFplVriZn4kSwcZiD6GTq
CAKdlxdTnZ5E/CkARM2h74Afm6Sh07rYth0S4ePm0qcx2yn4DiaADd79XYFG82h3
RJLkzx7lOFdC6+dAB3977bisWu01zEg/w4wrhpumvEM1nYbHUY4yZPMXUt/pX5ZS
NFVRCZvrdNH+CBfaV8stp2UFSpqMu0jOOcX8fMaFayK4rNA/n+VqifKm5H5WnPEe
ka4CFp4QxhR6x/lYMdNn9/AX7PScAZhEAJTAe7H5NBe0XPtvBNucJYKptgvdviIq
HY9u631qv6+SvHIkXzFoJ81n1tA333R88IcZbFpr3LWAaxfqSVYAQJ84hh9vSrEG
tVrIdXe5XjUbpXwudPPYyXdmrbLWydu1RBkTto6VTLWYmEqhsMf1YZ+dP4lHcv6f
QV3kHmfHbHI8wJMn6bR597sAeTY+67cZzLgN7l/BwUK8ZBWrorDZdR3oL8jPsXaa
vZlOMXtfzxgQDJbCl66qwHU0Z5rweSeFLLV3vTzrYLb2C+XqnYSWBVqwbFwKpmmv
6RaB2YULZVBuUoUVjk8OdWHIfkSO4KwqMjbIiqtUTxOA2x/K80vbVOA9SX3qpGGj
abQVnNbYCHGvQ3bfFxde3say3SdCxDavPPNu/xA5sE+bmkyIYt5CHruC3whEaFdN
KW6uZwWXi7OZO8+7XGtighImmdAh70f/pfkjpHVWcJPmcDZyAxxWRW9I5orVQOhX
1l7w9nEKdHB9DGdlYSYaPfx+M5dbLAIaKH6bCwK+maQt2FYMQUf1Mo941p44lmxn
MYWaL/MdKKhcrbNeDuPCxQIcme8+JTiRPWgo5abG9GoNAIxbyNmQ7ETaiCEWFoI0
cdSzHAmQP/hvz+JU7hvhxdexeqdCaqQLcml6HCUNg+XOpW/+zAOUCRxwAvjmaCCZ
ZZsfbu9KPHQ496Cz4ehUGZmbp+3J8LVEwmaAu0RNus8Ws0g13zXte3cqTOBL0YdT
YbdhvbTyYs7CVgU2IUg66dnHNDkjnSu7i26dd5qRiV6wgw83CuvZnKlyPWru/GFi
zrFXdv12rnVgGDMlefUH77yP1JAnHSgwJVhPMUUyrLTh6jiM5fqjK8yDsea2yaI3
UqRUv/0TFENk9qVKHtUAff5hFIX8u/7K/xDwP/Jkq9ZbiQQWa4mruNS2OpdrbLLS
VY1fNFoBt1xe5K3/WVwPZ5iLznYIXxnxr72VlflkIEghcwk0hPBpjMf2z8MlXSFD
SfMK2uT41iMMWLp5NwNZg1z51L0gqcp7myZWWvMQz4eUWsFKjThLjc3MoN+iHebW
XYQ+AbITLP9Xop++0gvds9BnMEubrtFjMzziuuJEM717Vn83bYdqXZiggww4FjFv
7TiCtuRXIc/Oc/6A3eJynEM+c6UkrR3k9f3taBpDcZg4fST8ZrYgymzf3yHRPiCp
bhjqeVHHE+/PchPaxDCKAGx+C+BZH5Vcdev0yiVzE/mj0sxnC90wEfrBbkkLhAkp
PSNACYVrruHltjUsYZyE5TiG3gY4ajOCoqnGlKXir1p8uVd3Ab3qlCOTQDJLpW3Q
IKs/KrvSwiP3ltSyOQKa4LX2KKwegYcAqGWNrUQDrmGGSywApZDcFm4GtkctzdzN
Pc3WvHJ8H0iXqEzZnMbH0pqjQ5nVJEzQ/M3f5Wjs1m1qaH8QuXf8yFJooXW8Kd+a
aBCrTlBpFPRim2Ro3eyFcRzX3VR3g20/XpKunInDU/9kExrudMaRd3X2IeNWu3Zt
4WicFIT1elyowpgxP4V+p7A5nC7fiInK4MsWdQ1UXa7Ekj+up8siDsncWRy57SJs
ZPehFzm/XzEQWUMrEHScn9EeK59fAWLk95zj7SdhNx4p8bsdLPOhis47JwDymcga
lkYoxUY8WHLbFEeBmwS0d3Qgay7Nc973r55VJ8CyhsyEVo6XsRYMXIGeZgbd2dVK
qOJ8GKhbMmxuZCU5VxutEUTuO5cUKqiLfsNsx1FfDqD0mBACEoC4UkAWCwSFxkPe
iKQeJ9H8LElYcmUbAlTBjNTrFLLREgLMdQQDSdVrSzGFKLnWcXDdz9pUtdbvl6mf
03YyybaJtbJ4tU7Jiri97VX77Fhxcr6miqUFopTXf+qbrHhA1WKV87fFTBzsA3sK
9x98p6nFa0mnLadnKSMNod96fq1BqOniPoQHqHVnn+qP4WR2PBnZ9e0K1OVXcLah
VmVRH/zgsxg6keUW4qlPJlMh7C6WzGIDVc4d30kiN+lD6d2xnlgSjGZFTh4MjM+L
Z6stiL1XImeHDLRzmgfB84UP5lsGYbr3siEe+yp+Hdmgl2Rmy4LHG8Z7Gv6AhqwD
Eyz+mAJJU7yFEkL5B61CAqsWneJqwra39eksC2Krb2RA6/vuErItE0SqBQj3HN2n
GZ3BeT57u9jZN3Mm/Dk86I3bBBf0cOJ33EojdTqER9SvSXQ/ogXM71NPNyFGX7fL
tWLjpak2E4uoFv9GeNJTE3AgKeocgh2zRY0m5eUl/SVc73yP3VXutyKtg8a6X1H9
eYUzfO8BPTzqTPuuMQOIrkXLsbjVsXxL8YRJqVbnYQUTWK+/c0byVw0bJ4HWJjCw
wXXC88qwIHanpT9olL8GnvhAivzfuIEdfXHC/PGVvl+iFbCparN/L8XHniQLo2lK
ZEsqma9usTaUhFlrfk+rTWV/1ttb9lROTbUcAWCHM/OtG2cS2ttqnrwK/GlUlud6
KPcZObEvTvQq2LXjjQKnW9Fg7eza5pzKlVOgsXhYoNl9NIB+VPDMvpwewWY+2OFl
T5B0gqmxd6oJQGKcW8cuKA0q9RPNzFDsQsPI41k41c/FPrQljmZWI1folWu+PLPl
R1DJ7hIHqduCY84lAQ7ZTE6hCxMZvGlKBdJPpSJLsnCzMZKkLM/kOE9QjwSzuT7a
nhecSEiOY+nDwVNGwX0BA8Wpxys7ZBpmFZyNZ8hf1j2fz0m38SdgbmIMGuHoPXpN
61q4fwMWCpFQnatnopkOCXnEQFDz55olw2ymdBrsnoxa6Q/CbueHiPdas6ugCbBO
Ixrhpp8Zg541haI7BLfDMugGCHdZ5Q0V0USFA9Qc4XgZ12eKuLVc3KXfGrgAGvUA
YCNj2KJ/bFBo5ccgPfEo3khS5lDssEPH2LN/8gfNGzsn0ytg5OnLC10MpzTt5c44
WEp3rZvlNvwxlf1E4fSiYkTAQeRC1/4UTD2FDOZXCB+p3lt/EBVOExb/Znrj0s/r
KIoss9AImN/qaJNtqw1mbnMHAGRZi5/LxRGYggI2wmNKHH5bh64ORaj8IQDi/NVE
OdiW0wMIiepW2Fpbmf5pnd9+dgg9aHHObTtX5kO7Uo8ffLEngksE974PIDxs7mNj
RwiljnemURJDLyFI+Oc7Xs8IbkNZKGPi/pXRMaxmffrByIKLq2kMRVr7DSgVz7Rx
QXi3teB+ppmLMSrdUJQWe9/KP5XjAV/wwK4IfpaAKX2Q0rQFTRraU7luxGsSe/A7
w+7At8u69Wy6lAswrvtXvPkhwXzRj/jFhtv7ee+1SxvyAU9jg+ZRasNNHAhRl2RG
rvW44Pp/23DyVVDh2TaoZ4ZabkFOYzYyeacuWDV9xsL0ohnYv86HaPQQsGifYNkP
hm4SYg+bFJOQ0V3NX/RmsL6Xi7Vx3tgSkHL92xn/JF+bwPSwP2fa5DUUJDcnKW4c
UOqDHU257rY2wGodZw8SkV90QUtkWkaK9mx7ikuWXOeeFPsoQ6lQCtryyN0NEPEK
AIzsVGwEsJEqXiCc9rjNvBlZg0bhj7SxYGmtuHD3v8HPwPSO2TN/phgucLLqlkJ/
ZDROtU0yiZuIpL+MotB/aYe7lCJtq6I9I6LYMjwvAV0a2ltQIO57J7N+6taUgCbi
UdLwBCE5z7cHje+9ppMg+oNG1X+cAWwyvN153ss/5U9+Daq0L0SuvZv0boBIjK2h
0ZAqaAhCARHpFIMrPs6he1ch5n2jdENY3/CQTPwS0qHkZ1F6eXMoYAWytJaMIti5
d6dy01qdHK6bKL9wt5ZF2OL1YMXlVvrBGcylU2sjLXZ3G2O1dGpPWSQHDXTKB+S5
Ms9SiMcShslsxdezz7Hb5JkZZRICk7QDWcKWtoWTviWSKO+8au4xy40NjBkjZ5SI
jLaqOQbV/fnFzqTbYbe4LtUeQN9qjWnOHkFqfeaaFHzJPDR6pqMiqYAt5DH3G+wK
6e4m9n/oGSkkKbYJujQkkkqDPFnWffGJXI5QlEGrgAjXN9FSRfV8HQmlG3T7v9gh
DvOd/ukvqDmDwiipkfUX1qA3M/UBImRkMtuWvXb31tEvWHLqpeKznBUhS9PV7bbH
Kb+wrN4llVkzFmM4kAa0hSolkfv9WYv7ONrleqDTaKK4fTNAyPyERN52yHNOCVZd
iQEfF9gCh5gFWK2kEKWD5Y2cIu7vgzNsf8EMpN9/V3LuVMMzJOdcaW/yOh3nON78
hSoUB0KGhNlRcncybq7ZtEgVaO459480mr+1JHQgiu6XZ74uJUGLp25V4E0mstxT
uxh5flvewQZUPYjnkK2g+dxToYYVbZwWUoCFCesVuge0pc24XUyeM3X+X8oEuf6N
W15/Yl1M+9iC4LQzGzBPFbyaTqX3YYZxq6cHz4ZWHTTs5dK5htzWR1+zwqchvQMz
wjCpkO08vA1mHbuxcE2QGGCFBmdnUeeJOrvhwTstQdpzwXRASWKx5ckB0cTTdfKR
Rby4EDAKcxhCeuzAJMGOvp2lY56tLzxHj6Hiq2jwqM/3iDf82fYN9KqIxT3Mv8a+
9fU+lqUBQp+a6+vx8u1/0tj/8SahuI7j6d2edkqg7IXSa2uwwtuOHjUMemM+TyGM
1ydTk4yShQBxWMl/1MIirENWQ/4UhoWuQmmUO6J5xz097w+D4/zyvX+wmfc+0Mp+
BFKCsoantduds9WEdgFGtWfY9znPOs1u9MRx7OP9qszA7tNrtljheMhILq4HZeZw
tjaH1UwKvaa8FHokX/BvSQNCKrp2oWFzwZw8olfEdDZAMzq1x2ZUKfRq7N+ZmhGY
4CWQulmVTC01gCrlpm8dLUt+a9zAlOdESaEUrjq1FJ9/V6Pfl9G8fGYYMGLFDv6U
2Xhyg7o3bWsiqUj3hBO71Vlz3H/HOMIeddL7jAreBHAWErG1jeUEs+9RTN5gCD0Q
xzBt4W5t3zl35kGmAUnh1AQ9BO+8tiV2xRvQ/q/OXf3do4DinhZ+srPm6j1K0QyF
G6sNeJIDawfHuFNZTpox6yxbV4aW+6iEFkVHA+XKEhock6cJBS4C6U4iaRwiLN34
9K6kFULluT32Qpr4k4iWl/gLz7nUFVJGuGZIR7uTHYQrbn5uHO/5OU4n+I+YeEUG
NiRhsjGk/BgVrhf+ipLMO8tg/Fh63pGDAJL44KTQZZj+9xq3ZBMmLQRZMzMMLMbo
M5AF8Q1w25NOibfuxBW12asnV0xC0KMhvH2vZHiRaxGxx7Ao8j5/m+WrYc8Dd8Rd
DUTUCd7DampTgOz7AHapUvLWMXHzhaqx6Pc9Um2WFeeL2lubBz5PuTNAsIb5x7f3
N6pkwqlRkSoNWCAUWR06CUuMB1EtF62lc87/28dg9kBFLI1ZobUeG7cRtapqZ3G4
M0PXa4yaJRGRgGbaHF4YzESM7+h5qktr/I5VZdDbIz+d5U02yRDNpDdpJjCbrgcG
Dwtsi1JQPsFZif/2Ir9MitWDZQLoI3OHSfQLDVQBxBfhM7gxUwctXdOg8bVWUkWh
DabESTPY44JbEhOPxcwFtIpBtTrB9QDgUfoHOeIv0gGI6YHCok56oBLuw1OThV1A
WlSP6jFNXE7su/bN0UjA/MCJ7vuU06dtyFC0yGBb8ifrfuHvVlgzSVlqa4CzgIf4
fXmVBvh4uUySXXgEfpCQG2h8GXuJa0MQR8BSv9nXOVxYe6ftkcSuormG6/Ptv7qB
sNFTfFWWm+3NIEy6ax4QVcGpwlbiZUwL/NTNQCglIzyYzFd6PlTETb0/R7g3AC3X
cp2QrIFqWn4U1OSKlB1alz1klAuXs3Z8c6Mgg8jwOamFRGiZNJO7BFnzPZJ6Dcpt
vw3iLEf19tbOuHfy1fL/TbvzIJrKTn25zfCqczeDpUJZLoi937qj5Nr1SqeEhPKA
QHDxwNqzh1/Aq2BfTf8mtGEuFebSr4NwY1sIToJ9xju8BT7JZrILIdjEFi2US43P
9wrWof0vuFEP8YqvYjteTMLls+fsncKZNWRTsJDDFhF+N9lj4vYmXh3PAjBuyqFs
gXd/HfnLEqfQVaYS7mXFCb0BOCu/TPhpjodjCAQzSkoO0tp/Wvjg3V/bMNpIoqaw
vJY0HNblgkA9PvjygLyPmv5/da+JHBcAt9GNOpFeU3Mjy4nJVIbHcmqNA8fy+Wgf
aaw39gKcbGJD5/y0IaeSstRzktb/IBhje5OStoqykYQFjfGC+y++3IPTxzkCpZxZ
7Wc3TVuLLMQLvRgPhkBDOPaCVSz/4qn9B75UMzYoGNLbLFeb5sbBeh8x3NYNT1Ci
frwSEvKNJSYn33BPgvvwQ+zDFoHG/5Ai3Ja9AOop7xz+ITlxQt0lXPJV3HsAZacZ
ati9BS66fnoI2FA8w8xauK6NVh0vj0zkNyX9L6EG5ZHrtFzMjwoq6Q5hspuNv0PW
PO32Twlj2boxEKvOSVCaKRpWFfLgmytcRH/GSDYYMdPN0vvfZRmzvrWLqbRUiDBB
dfVDN8o7aNpsq4Cy2KRKBgjDsVMYxI6GF3WBqaUAwTG2Xg8OebPOEYNSGxz69Kw/
ng72d5rNcv91jyNZ/SnVoM+zprVVpRiRUxkl5RyKi1lcHF853smqozwRcuRjVomb
/clDZpcSmJzVZQg9lBIjDLlhxKur3n4bQ4C/ZdsXMIYibbEiEiwoZEWwIQE8zT6Z
Bg1ExGZNiEZJEFlve4ubU+n6TJOtkRXW9FELK/+gliG0s0LiVcehlM3LnKuHv0BR
6r3B5YziTbWXgoZBP0spwZ7d/TRdjchgbQnsPPPcHE+02Se3BNh0FfB/EiVKjAko
dR9+I5yAGSpeYfiXdyH1Ul16vp+9A3C2OTLPTP/o9Pnl71xHeieBbyOQPpIkRANE
hw+Dt4VDKkHtROlSC1f4jP9Ivz/kj4icjApFDI7VZjvAhvXg0Ppz7iNbZs+sjN1U
djavyU0oKRH02dzDqrVamG5DwbWNpYLGzBdJCCNdJ3RitXJP+1XW2DpH6LbnsfJa
MLzrWyZa+iwksrN4HeX1kc0tdWmiOm+EBHXK2Js32axGIWjlDHf3PVuHloJlB9bh
NEBDGTlrwxNhqwtZ0TyEsb5hRh4HNCK3Ty5Jj60jAxtE9ZEnaF/fc/VasISWjV+U
S8sH5AgvMuS/YjtpTyz6+z831ICCEELl7zOKhNTVmIFOp82Gt0l11ehrbSlEgPKb
PWamVJLUQwowr9dgjh5nsWDsJjUAW5m9FabyOjN3Gymwm3BnXh2lMlPJgSearKd5
pAtdIs9OKBC1c3ZWtMpU27pcydOCB4m01aiIhPKrj+LNWXPgu7P/2++JqKov83j+
oAFdVUdu6fzuqKKtiV0TU29n6B2YOOyb7n8lWY94yg7tv6nQwPbMY3BxFp3FocL5
m/pkcazsHGZXF6BNPAfs76Qd8F5snxtzIW7+IJ+PtPxHEJn6w5QiIqKhxbod1A9P
gXpeYcaoaWEhPlYKXq1q1To3ndPdeayt+NtvpCAb0Q7kf12lZ0bk3hJudepPMvEA
9baioxU/9pIeBYtSer3p0+f8rVGjF3f/JJRUSTaCSGfFwTPIxWQG+qnAIngUzZiJ
cKwkJH/0E3UpazkZOIuD9q5TTZW26bJ/wZhOLJlzYnAV3q4A4ClhEgxp81QDE8b0
jQMz3FWejPPvgZAl3I2T91Ph33pNoLwQG6y5vjOoR4PhlTqZkF3l0aR6bXl/XpUh
sMaZxSmu1Pb5bVIWf8PNMw+4UCWVwSck2A0+w9UYJBPFwaQtM8x/enYHPSlBCo4k
IR81eDOjDKaEspO9JajC+Lz6GIoQpO+2PifkbbMkHRbrPbyL8jE3lCDt7ux4KSz8
CXEPNsU5H6wQ9uKToLs017bnOp9ElgHRm+iYhgIC380Z0Nv2/HnxUti9cA0S/rLT
3AeYlbs/fXZawSlMoLm1U0iKLQCacJBP5z1R7t+8TONR5HkrNuDNUt7rmb2Do/CG
K5/WPCE1BcEOXufi8Ddt+kBNawXdO4byKGrLQkjQCQl96xdqJwU4ihOqXcgC2lNz
Ocrl0ay3vRvT9B1MpON3Y2ElfbC80IDv7XWBl3xX89rK92f6m86tgUW+b/ZToP7L
JXZXtgCQKusebj4/u7H8XeChFtc7PN+T8XwYj0A/9MBeW8nGkmjHUUf20bja5ViG
r0W62NHtOhglrB9awg/hTy4WAMnNaFZ9ah2UQkFS89pCaXE4vwG8zm8vW/tjIOJm
JXeCXEmrOnr4LFG/0Iw/vDcemvnDAhHDm8ZyA7wK8pvjh3okLrpPykR3HBD4WdKM
bTFVA6y1rb6SxL6pc7i3jOR+VyzEnhg62hMwaJ6AcladBYrmuw0KiVEQRgWf1jxG
p0Fb+D4CUy+Ep4/2JfRxe6r/m2JRW8AXDiSqJPv5tC5mqvSN8sQTY8Er58oZZtb7
3ObokdTvuKoIID8A4dyyGHmQ+bFKXBW10huC7Z2treBJTprBlKqRXMGDPR7BoeG/
h/6ciRk7+LRixBUpopo9LtiVQGsaSYZ8sVABeJ9+ZdAbicLzSlP6EcT0awM832SS
xiNC+MqGnh/f5H9BvsP1a7H0MGy2e2kjikoUp6Yo6DXFQk63UNH/VK6iXPFZWUQm
/XBoaF6QOtu10PZt+WrzfkHkXmbjY98lmK5w4LYQyrfZEqeXfWY718XQ2ocADoQd
VM+2cAy7lzooyeCRD/xSDzY2bn7/2ZNrqaZOwiciqLcIRrEnwVq9kf/WlfbUGdJD
FHEyxQBFwAMeoESZx6H4XcgrjQvSYYsEvmBdOrTbSOdErapHeU+CRNYvxptewg3D
onza6TDKNc26sfyQfNeE90vjqTMJx5VmiUAe402JCBIvNrF/LdZ5pV04W8L4sybS
8LOlgDE4JrYZ0b+jh87B57hTHvsE3wVWJQwku8QlwTTycD3IsQiqqBYbrdFjOKzN
/vOQHUClfwfC7VC3GSQtxcg5mSlQVxnUpc+hizAKWR18/5HILh+mQIxD7Gj3Tbq6
WgYtFtul8KCdXuLLlkMXadBUL8TTNxsN1LlpYqpCT8tzsp3UeVwxCdf+XMwHvprH
ppwCYKZnIwOsIoRfbb3DmZZoYHSGX3QYtSlNhBhW93orsSUAVSEBp6doCeoSZmQz
F1UdKTBCihFx59G1zJIISj7Jz98yzlno0VT8N/zG9oJCcA4xFKdzazyU5TMrkiQ+
GaPa2KHHVftZqRt1Lf/aWGFlHpq2J/sUpi00Sc/He7j6CtRec/jQYcYC+KrWg/Vt
pzEL4uRneWA2dcrtyO16iAQPYcKUrtKKVM+Gpj+4xhPjFGh2heSuc/MqgMkISrCM
9yFKbOEvGaiTh6FiIJ6u4bdgHNU3fTjCIJ7Tbl9fr0mypFXPTFXY4OlgXvbK5Ys3
wZgJVhdZtP8iXwUyXwIDlAskUv1fO/vlLzhjcbvnErrq2QqH4idOaoJaaPYJXf8g
qp7uQpI/C8yFDOiiQGjyRSB1lhK1s8K7RbwqNSrbEOZ8LxOuezbFDoZ8Cu8tGOYp
Cdpk0YVZarHKdNQ7wZTSOUShzjHW5OF4j/uP+AqjD9aLLBrhgOpJv5KLP6LaURWL
7s3NI5fzn03/V6di5NeSYtE8o8+bzlh0z6jRVNK5sKLwn0hHS8q7eGvRpeuLnrY0
260X0Sprw9NHZNYj4+eIX6omuTU8Vb5bvvnAtqSq19D/z/4m234FNRjW7qxUz6CL
n9urITYe7orzznvR833DTDcttvL7Ke6caAWxKBYdFNcDNXncz2bVsuCe/xRlFLBH
9Pw5mzQEbQEBy7gy/Cfw+Ig1KfF9JDEt8a+XW6pTswVxkNqZzaqzE4uecDfz9Qbq
uSu8rRQ0sNzO7snbqnuQGxkfGyqPNXosgghcafagvSnYpfIOoMeQ3IFdV+WnhJ+0
HPDLC//Ls2lgDKHpIjB70glrHw8YRh8bfCB7NaMXg3xnQEp3/LO1b4cdafzZJY5q
SWFzND2twwcmwP4afVjcSSW/D7gT26DPI+8iQqHM2KofJV6EJv9NvcxnQiaSomG6
MpMwOeCEZMbqp0tUzpov6cJTcOM2TS80f+5z4v/YXF4lpwWrHae9zm8iH7FIFp0R
yo2p0Opb7KJtgPiBdMZn+PvXkWcQxborj/XzmY/dF9sq1BX4SQR7sRGZ+jV8l3fX
Q2h/AeOMxTfr1RkCewCJunGqUNi5GMvTRPU1VyfpxGCAMD+YAb1OxmtFHEhJe0qk
Hqh0XefuEOzL7NYwqiHbMaAKWusDWZFSx7iSSUBzU4uPW4a/vKldZeNItw5h3eGJ
6uVcJRLKayYY49aENq+kk9No/7fngyZzx+Rd4SXFBOsAbIVAExVxmyOmdIXFhHLC
Br+38O8zfANrnjZRkLtzyilTC/fdFyw1TWn6ujW3MWMT+8CTKhVtMJooycWcfTHY
1gToa2H6TJVQKggFuDSCvu7mgeOfWkRm5d614SzXLBkNN+vP9uyugAWpVV4RyDtr
l9Y7/0l91Bv117CB3k08RJjubx/qnqpN32lATW6YFSHCc+KHkpa1rgTFepM9R+kZ
AplY8AFKRQiu5LRktzOVKM024hv42EA/jGXrY/kNsTJ3yq0Bt1eq+W679tkatVuY
/5RFKInVQDnwO5JNPjo6TVpfRTY8ZxAKcT3YMyL/ijkxxitNNX33W3y3NWuE4Wr6
LDpp7ym40wdMpr3tyVzh4+Tc1v7+OSS2SkkYq35wlAZN2AqQCD+FGiOLmQq9ZZIe
5qgVgl3VDy9uXFsVQhIWhadqTKBmucT6wzJJljhTpE/0yhpLQqUtcvSkoUfz3ymB
UdX8Lfh2ka87ewvvbR/uVbF/TUriflRlsfDrercpBFB9To/6AXMaZNZgmHGWwoj3
d0lxpsgMAVEVAWyjJjKxlpLejgrozkrLT52B2CMAtrun81HXvoQHPo+hFTBPaXnt
G2IOGWdRt59YT0KnvMppiJbFMkM9Wroffco9a70Xw/2ljrwf79iRcb4JSyAvfb3H
FCcBpd2ZgbCAxw6GXpBDfWXtnfHLhusyluQhvHW8NoJvBt1XOAd69KzxtbUyRi2n
qg8kqZjZscEMTDEEod7SctGmg+xJc/EhYX/mlfuONHKIoyTsXkVvXUfJiQNpp32J
ig06Y+TxE5P0uT6gmqEH8xh8SaqfxgUte5UXNz9mM8Z0KbU20n6yoLmQsHMBqolp
vdkqb3NJKDSP8UBaQr3izWGkbjR7MVu3yXEZLeZW2Gjhf3vQj/8fLo7jMZqVCzug
AE8swT55jv2rEJr06a9KRrJiCQioKrJutUpCVz0pnZ7QIcbXp93NU+mfKzJpKDnq
N1uY5noEQHtgren8bAP/d+k50ZxlrR0QyEKKjNJ6dtFgvv18Ul39CEM+huXX30BL
/ZypuZyS7mvKneaXw05hwtDelHgXM/N3bwC4kx4BhpqdBD5s+xxYovSXDlP3pRIg
QpMKguRibhT7QKdZUWUJYzBiyfvuXG0wArLgeXT5ONZ+icfTWJoQmqkGRGRJRlti
jE+ect+7sw3d+gSeXQPNFOJbn2q3VBSV2zC3LMh7367YjbDTzdNoy/bh4i0jgvcK
RsHuyAaJqWFUuCXkNrnrzl8PnD/K5nxVH+9HDZ6giNJxPn890NBdoawSEo1ctnVX
WhK1f0kXnJy1m+Y4ZqO21+vOI5UdFnqTTA5AdpKCihqv8ohzbVHaZNAkEi2ZqXOv
V82A/DUhDpYoR+P9SD699Tzl4QirbXe78bwtthI478AqLWk9EualMMIxxeaay3Al
egvhwoUVV9/lIlgi9vxlgwb7+45pLAnvXU7E4lnhMeZ1UKcMMiLzNGWYcrnNIpUl
gkgGXy78qmh5CqPPZh50H4JV2+zt0riJg11cgU59Fgum+jntgjPCfuaIgGDKmUcM
Od4fJ4FVSY3WiUcbhBb8i3N077Au6JRk3WnG/rhVoXSFGHhhYEvppJHc7oBexqxO
svcrcRfd25T90sxGWIe3DsDB++7VjoaYNEjgQ9X3Z/ks84Uw7/zNZ5auE8U6Il+G
VsXIpTbsBaPVPM3bIo/1GcRX0OQGkxZ2srX4IARI87BXBk4Q+ZdLmqANH98e8p88
fslRWCvrgFlubyb/N13064/rMhIcPxdwiAk0B9lSG8NAioUOQwaJ/au+pXp+blv4
RMlRjSbnbqnkBUe55obj6OBQqKbu6zBBmgMqOOziJXhl7eNqWUj1Almrfapd4uBL
enJsSWu/deFdZ8Wl61kxS/l5URc91bpk8IbV/DslO25cVLst4B0vhSAUcXo2AcDL
7K3i6dTWaKZlhO8B/x7+XovJxdvL9Kwf7m3NwNlB7JB2JaEI0r6f/J7p2ogMYJoH
BA2Ywu88fpKBdVbh2tie+rdzSn3lcjzv+wudm0iVE3TwkuAubONNK40FCXBHZnED
naK5O7r+nsfh2+MltJZjlP0vTm1MpEwy9EBZzLkdN7MxVrMsI4zsBsCb+qV0ISZh
721BqdHv3lJcnp1O93u5rUzOM0RHZTbmmiKb2dQgvas3W1wdxQImh60rQmg8RWum
Q+zka0ycDgWE9kEekLWXtf+4e1AzsxMMJ0JzD7wf7n+WHbc4wggJZe4x9rH8nt5o
PwyLsnSbo1hwEM8gio/THqWc5kPRbVtA8UE3xSA2iy3ueBQ4DCsz8jTYWu1y0aNi
r7OvsrufsODwTdql3eKd0urzfVXqQej+VU+aZWafCirSBR9vK2xO7Bw6/0fVtnYn
tutxAKPDwtMZ6q32t4PeQ7KALlnYUWs7LwTyLjr3Kes91cBqpiiZacrsz9VXlJWO
idKmyMp6Pgbdn7tCrexrUxzSJ6ZZvuLJ18qS55IGsWtJUfWJ8R3Nqr48vZ9PzT3l
WofUSlACwxld0XFs+TV8uzclK5VbSwr5moJ4YADmibvgOXulESikBQqUknHhWh88
gGXAOs24kdeRVCrKglyNoqMbh/HK6oIjUaXHgeUnDdWji6Ndry1XrsOJin+G356I
8b+X06mPA2eUoXLm+Mk7DY4+Z5KBjg9HExGjU8PgDeiGznfooTDihLE79CQoUWYr
kNVHrPa1pNvk/YKXk2UJ/LS7jG5jDiUN/x/ikLJ9+/nyi8US3OK9mKBNQsaPUAs8
GayGnrzavr8t7YtzSvKyN2eNL/8hNyix24zISwTv1Bb9Z4j9LCJHbXfkodf5GnHs
XNm5kjKLSAiJ4cWZewFCN2EsS1FMsDOv2zwJOAFxCXIjqHc9oFacnFVs+zkZkiWA
alisKObQcih4DElfPe3qbc1kBpbX73cbXnMMTBZw+zKtpZeJKEV5wn9kkxpOIuyP
DK5UHKHvGzpQA1rpukH1gGii2j6XJzmkHBJ2PF+6H1JJteC2Ke9L3CcywvjYk8vh
UQas/52NxjQW2rr6vqz9ZFd27LOgWulRIM3Vjof4X73rzvwX7P0CVXdwdtlDZ5r6
BFsxM7bvsZKUBkX8t/aK+n7F1Pz4LZTD7YFM1Z0fTbzfEX8Xkdk+O5m+wB8B8p3l
LF3tYQ/5dyvHVmBG92iylUtQ/IXYi93WLDHm2E1zvm3Xanr/nhiF/QgbJqIPMOvv
6pHPp+HVRX3nxVYg7wOL24Jcpu0rcR5/gH6927lx1T7jnxrV+5haKQ0MR9V/sbzZ
LoxoBoUGTjmA2iXC/iZAn1qPIqerzMcOHFHv3/88GG9CDbdr0CeDO7cdYm2hiSb9
DUYPu/guSXTr5Y76Gi3vXOtdv0E+Jmr7+u2a86D5FYlNFySnWAPhzsgom21j7YW+
5BYMl+W6BTLN6CPOuzA8FM4QpzmMSH1j50B3jbLs9wPKq/BAiqVuVWs73Oksbnxk
DoaPYFN1hH2wkeLZG5rtmgNlLiyqiPB81h/K5yCMBwwVH+kgHyCvgkpc1h8B+PJi
DJVWB3ssnl1hQvwkwEpaNcSZVyVvIotWImWA59yJb1XKZkX91gF1IXhWj9/YBJMt
vYtIecRwRtWvJlq8YcaQ4USBhtjt/GJFDKKxmqpzumxySckkP3Hd1AE/gwl7kIfc
EPaxoTeXNC3C7Ut4547vsMOcrF1uiQFqXw66w6kQE49gC7aRZ9Fe1Bjo505cMCyu
QdQ6Izx0krxHXbQM8xUhumgO+/LZfN1dVdDVljH+pEl0c8AQJJsgSVQBkT946Zzf
hpImj+B+5OynJqyImK6QuwLD8Jzj3z+JuWndNAcV+p/wgrkXk5v8Me47aios1MvM
DrqRJTJ+ndqrsRa4V/f0WIypA7dND7ev+6DHcKeSYUccarj6dOygfaZ0jgyflWWB
9bUmkdhnfxzJFhhMkt1IMI6QdF0g/pkdqWsHruDxTbvKhWTRS/GJt5f34cZ92lQy
CspSdmd6bBUFBYIyhgV8qpM6Yr2J+RxzJc97LGouoh60w2rpmjG7KgfJuG6f6uf2
Ki1f0p8uU1ZiGpUIXyXKja0vF0avTRTv3Qrb11xnOl9VYYa4MDPtCiFauohpGleS
vS5iK5KcKDC05n2lwTI0kjiPRysc1xxnoL1Vdsyz4eYqpvZQDkvHOrKoZPOMc1ih
hk9l+gRtqykkH3wJMI5RxMkDApAvISPONBMwfEiLkJLUUF7Wq6YLIUnTdquLgWwr
elR6To4cmQX2azEfyUXPzOi8vizJkiJTmwnY4CRoW4NnXr7K5ygUc8Qi68k+/pPI
pNb7USvgMQhqKGo3QGurPOjUtfQT78ora5r3BDMoVOIEpRWxwslUs8zStWSxvyH5
jt3g7R1aat2arFQNIewW5XbV5haxLOOe4xbqRbfiMw3VsIVnnMPTk4jQVaFbBd/W
45hp4npfgnVFnwO6R4feENC2c26tTp+mWHTo5yjYTG6iXyqiQTDV4U3RvEdDlmwk
9jhG/gr8H8Zy6BQKTsNlHCpxL/0FfQ8UYDnRa+9jyMxuAj+4X8h2P4weC8KYMQzZ
nHuOm1nKGIS7OGKvg+W9zHcf6i/OrTlN/rMMHe4Thk5ttEBNsG4vjUCpLpx/+rs5
y8BYCzBpNk7GbLLsCUyrTFGgdG3rjWW5Nq4GcIua9Zz+6D19ov0SMdN0GCHy34VI
GKwwjwxS9aOwI+kkBMhSF9vVLl9TtM9jELkKC/32V/OwXyE1M8vp8J5Jh3KcuXRM
eH1hVSXSmNaeyw8kY0fVA4CPWTJcdttD4tQ5/11vGzJRyJ4P6hxFtNUBeXLuo0lR
Fhzfyow/zq8RKSza9xq0QfAj2L/6RwlZKvrFJx42iDKSZKhu+dXKzMjo7mZ4PSdE
Jv7vl2H6UDftS+hhsdnqE6fYfktvBMZowgm2U2hmJNN8mZX1R+lwEGBMU/SF4Shw
m3ow7gF4dFszv1HEd7TU+XU4Y7cWOvE1Lk1IzvpweU+U5bfAtqrBBc1kWLwXC/7T
c0fL5QTL7iNZjhxsUF09gNQtSXGcSJf6ImL2UPIaN+V5+yQZLMoZfpYoViszmvMu
Qkv3El4EvhKljLYQoWu0aJ4B0nn0sTOTFH5gv9Ie92S+wNW6WDmWtq5P784uwPnj
M5fFULiKJabtmu/kIbmt8swoQYXi+bs3ZygmBBWVcwGXN9R9c1iF6eihdcMXhnHZ
roG07usRVXdWiJKYuWucqc1U1OVgUKTku3vlDIKoGDxl4vCrt2Tn/iadqNea8uCP
BTDXV9ZkIb/cJRBRjU91oz1FqqM07nf7ZvwstWjI6wTl8RDVxyStFoM3MvNg92xX
V3xIw3mHRfDsaSoNTrw3fyPPU2FtTs47r8nlUKUw+60FnPrCmyIadVRP1yVF+abd
Qu8ziQGl7ffTPaVLPLyerxG7sKF1PgBzojFqPCFRMq4qBuQKejv4HotzmrZLMa1H
yT+7+fFcF3Gm/ACx/eH3UEMYtlv0PcdV0Hf3icnJla+unSAtPfYdM15Oj1j7R3R2
/o6sHoqzVqdRSGYxQ12lBr8V4brJrqZTsJ7uzkh0Plel4IikB0HRFAkIcTWGniCX
v862GlsQ42GeNkOz8XDEG7rl2RZzj1lVuJD4UEKxl69I0GwD9LiyfKe5l7KM+r+y
vvvHNwVgoWNFz9Tlq/B/AwUHTFtJ8ecw4mIR47lSj1t8FWydKvrUv9HAI9JjWF5+
+vcH0eXdbHpgBHxjw2/llFEA75OuuHQ3eBNQoSeVMMkJcF+upcFMOaVQMjDV186e
9bmD0doEFZRWOWNUyYb7M2QIL8KHAATL7KF323d6L5bEF84YwO0uKVPlMG0dn9li
y/GIq7Ire0K8NXYO5vwcYYLRjoCI/qbfk3uHNCDDqnZKGniGExdnVlPCyhQGUql9
mYIy/yswHzS5/mJgQa94S+lhdekV2ZV2XPb3SkIFI+ejMcT0fk/aw7TNq7/wNRmN
Lq9zZWgG5WQsDz7ZUnLV8HenbsSjKXYrofKtQOLFe3DWMCEf33g+acUWVpvez1WV
vfDTWSPmtqcY6sQXzs7DAvdWxmUkYx46q/BNEIssNxuC/P+Jb8uVdzs8HN65vWGM
kS3brcdIrnRHxWc3sHoAj2HAfl2r76ByF+rQ1xJ6pe3QNXkzmN1cKPjh/4CmFpYb
7ke/3IIUblKXzx13xdFffbCOm/1GUSDIBJ/PwkPsE8Wh+MBrXHKK4ouNhWzR8s5w
Rt1E5ZOX3NEfy9WDWW6WY4239EU5MyRvqVUQ2cKJUiGFKTe97HQMusgK+BVl7L2s
GVkfmYzxKsk78Kg5XHjb88KnnQ4HSw8x5EuS1FNn9vbO3Vq4j3RjuRC+340MXvhe
2lAS4hX6sn+v8Lnt4L3O1bkx6gf/r9wO23Kqd7gLjY2Rnc4GyUniv7gXAxkBWqBl
0g9xRL+zaADLWdqs1ybznTPSxM4WJNMLkI++aZ4Wc3fvwFMP+bQQPQWnm+VsusnL
lEXekwhN8Ut1D+twkqPlPgBE7SLr1JPOkA2S1nr0p0sdmgiUrj/OjJdj7QrJHsNO
0mB1gfwFP7ieG5I5eAufxxHhIJMamHi3fEGBL/vV5PAliQe8FvkWcE/lwzmdosHk
cgRW09yrSNcGYH+vULDnllsaFpGWSAbT6ftX15Pn7zvy3u63Ybszk+cc31Jo71UY
d3cyaQcUXwWkM3prjVHRJjoUsSeElS0eNSwzfMFk1G6qBd8ln8rkMemcUhKFSW3N
ysF30+fLxXDfATPZjBAnCkTjxNPFpUOG8NL6ez1sZoSp3Te0TOS6c3tjMEZEmKYC
RiV6aw3KsIr4YwFqOxeBByRJKBwkLiISt92HArq2rsr2erfp7YPK9KEPOdFxIWBT
t2A3IzCmSLmwn+ADWelf0QVrHof5602wDIJ+tePEeWKHFb+PdsNL1wU7VZzMPGxG
hoTFD3MYEEfFaCgK1Uq0af23uAKghqoYaWJfj90SFyQt8Wg1MPAm4cbddKrJlV7b
EzBehrPOki4sjqxwzPvvqHA84x6AxWKFDuyTf8F3coo51edQrJghzhqWluozKpTo
iI68kXiwYSTHRMzG9IM4+fkDnOOJkVbiq1lC/zlW+yPK6MLPOYQKi/3Z1QmnNqVu
O+aQYi/X8fp797dff5A3Pt3asRrmQBblPp7T2I8rAPAYZrcGh01hjBfkFw9JKKRs
tE35xDBarQ4cwLaS6BqrOKH25kQkfDHJ0/dFY8p9g2hIs/wGQ5UyyoK+B5X8mPSa
LQfCgLYezNyIZaPD8zto4TbFPJx+JKocnXmeThLUlk4MoZvOF7rpG8Ux0RngaDCR
EdNNfAD769+PZVGWrkGi51UzkncubqMxhSNUV+PL3TYwRMTXChl1N2sR/tweLSOF
kJkRWsqtN5RhmOhB0HlQoS5h5hf/dyIkUzi/hZU75q3WkCu+XgsdluXEAUb6JNOg
O4qctDhlfobzgCXBpPjaWqfpYjgH1JZMMtlQEuLGBnvA/pd6CA0RWlpgOMJ0gMHS
8l5ov3JRCLIyboWwJE9odcgGrdVikgHA2CSQO+7ShcGCtLubzj8S01FOXYM6TIoj
r8KjhihuGOrTWlX+6IWKHg0JNx/dZixZN+3uQXlRQXLXszwq18ttCqt1dcPlROmq
mjpZa54A1j9a7rFr5MKoZG+idZ9LDQcHb6GTBVbFdxgFj/oqf+KOVQmCDyI1+GGC
J7YDveUm5iFaq8uFSTqbTQOrej2RsQcxoHa8ANgRvrn4GtlmEVkTSFaLXqzzoHvV
D65t8aIr9o/pAxU/yQt0shnnSu5M4GhajN4ucAijUXwGqmsrNHbjOmKi4AD06IZz
r8cUdp6wp/Fyp0BfsKXzlnblqCtrWCXbThQ/v+27XiCSjCatLC2YPYCzdxnQsk5p
PaS0c/zpo0vZ31NL2cRNnBUho71l2ZFBtalnH+okZaq2otJkR3d/Oy8V9e7+fzL/
AZ2PproAfrP/F8L9zeAFi0w/yuyTA18S42+XG2523h7XTaceM+1fqZQ8JYxqO33D
+kWy5J9EEwI/Fg5EpwieB/cKgcfcqGhF2GqdW2AsIVphoQ6IOrSP9Z3C/85qvPQb
jat3RLn26pIqeYxgU/a6ZQ/8chSf2XrXtTQt120zq73oWm7WWQ1fhqWTVZwWZHMN
OoqSDKa8igk1AXeAQ6RrPxeL8dEsmPQak6Ah7vhnbDvoK68OdUaX0lH5FAv6gafb
xEmOn5044SIPMuypoppj8KO4gx44PMhj2JfkybC0YGki2r1RhuwBT2F9G7Gmp0KG
MNuQhdmBtGutPfZ7fuZdHyTQ+oUi8Z2ctr6CU9SeEsbVHTXzfu4BlfSkmfCCSXFT
9jp+syH4IhPNlkRRR9macipc5IQWaI/Hd0Vsr3gvKx+fhcIqUIzIwTMFOOI9GcWv
WXtYW/MVfo+ihSWmTul87BZiZxr5w06vQMiJMjXa1HZzDL8LGnJuxzudcu8Idk3R
6jKUdmLUdAVZ5ch7rdwk6tBztVvxuXleOpcoNf7oAE8A2jA6OmROTOeY0B/sg6ZC
SjcrFljvlij6rxf1mK59DaNwIrNZgvqaQ44F6XWrFfcC143LNPAJxshxP1J3Vp08
1gj40oHoEwMtw/gpbWWqI1cuNsrrqeisZtRvUoftkRJSscqsJzv8575qvwPbo0Ye
47RrMgyDJ5xAuU5kSkyWT9Um2nvSFJ6y2IcoSZ0xDONO8ypDrToTsKMoSwU1BaG0
hLI7vMyhrybSiYVuZqgWlDo0wBxcrq8mEt0grq/E01cVatw9z88pZB+UrfvM2Oe5
h+gGGgH56eOmS3KviLjOIrWcrw6zX/UmxTxkJLG2sNy4YaL6UY9uMTuhJuZNuYLb
WisFsf1eM+wBx2iIal6NHhmNjkmGqfv+jl0sfMMAB1X/qWaaiJ6/S2Rx0MxSrUrv
zL7dMu5MvL+9m+mhKg8GiUTpagmNWk00LvMaWI0AB8J6o69cuhM93TUwiU9xd2kr
YXKCdqjEBiclZ8GNGuIfKlBlIJPzhbumuI3S3kbuxr61KeCI+g2dOOh3/AD6W5kR
0ucmPXucHiVHMnMH80/WtxDUkhX8xGCpKJCP8nCzYJS5X5f57SgMMPfTMbLYhyCb
BI+cv8U+ueItyGdhq/KYdN4NaWcjW8gTry04f1dsuJStRl3NsbC291i7wz3DcEVO
wRp2fxxvDNb5kPbFGUy+HvfqfpDw5Rxi8r7swI+KTjHj+/4ntVWV82i2wsBcVuMB
onD+Q9veb2Uj+GhzEvy9mFYCUT6ziIjV+x+5MRYXB3zcf7Djfc3PmDeb0JwCJedc
wsawRSB+wFn3H3odcElJwTcOeCKOPdfDu0mpxlXCjN592KOAGBPjdDZAi1TgaBRl
/da3jP8qcACRpt8oOD1V0cLUZ+4S1jBBYvusSlM+LFtFtIoG8ja1UVTQK+6ZZAug
yconSm3v4efTaIsPF5cdOvHQhTS0jjowagJWQY5NJawDuDWelnV/BHZuGjzgGv+X
JogqDbqrWVmHhYZ4H2gu6Gh8IfW9mciJEVf6GZtaEGg6W38SJkTlFl4d8cOAWW+h
Fa4uEpBrjH86qhEzx327Pk7VRCRQ494/GZm87VmE3NuvOA9FuOUnqXK/nfxwb21i
OY2VlKenjphInX+rT+8J3mbxngB06JbD+RipXMCjDQiizTOMkDdQlJcPMxiqmh3G
OEqbS2jVvMsTI6mcLeXehFWSlyrBs1f62QkyF+HFs+RgJVJA8E9uUUsY+apx0nXr
e7yNJE1hWZyihwvRn5R1XScQVW4S67cxgUhh9NS37MZ16tzfkRhlQgp0nmvUcp4w
q/ZoST26/Reo4ZGR+ikX0U/CkWEZZ65sSD6bs1nrerORyDMdO+xwSt9/FRqjsJXf
MxxyhaNHIRaiwlEuWKURDV/UplcruNTTzJk2eU/a74TtuMsBM27VHsKTKK0kUluX
X0vu7q5labNMxmxXLOFYS0aNtjUhBvZXfyIxZ7jzd1GQcfLdZQwscvcw/dXaSRNI
Z818p9zYEPEwjPFho7PIE7UfQgkz+syyUIxIosi6aqX6KzkKSHGKQIYH7QfBttCA
5k7eo6KI2m8KF10pTEMVUYQPVj0O1aIB97z6HOozNqv+qeZcLWmjDvJx6w+g7lyq
3qEYP/q/WGwVVQG6qMo8KJLOf/VRZToI5jaim4ir8uCqcukrZGGLjs7n+DWceYVj
dNXQV9QNW+z9knBulAstIgH/XOvzO51QpwnX4ygfch7ze2e+mNjvJHG/p3BYPKBU
b/6tvy82KKpClq/C3eQdpIRwrJpAp0vST7WDA1gfg0cj+NM1n8fcTOYY0bmi2eUJ
d6Va6p+4NMVVT3Eiy8CbdZRVIXRqZPc1KsNAQjVjRRzbbG4fE1woKTRatsFptkZM
svnTWIt2fKh/pZ+dkOTAL/0RJH1b+ZghjTXXc2Aq7sBWazyJHTUuljhXnf8WXFNc
8v0hYzs6+7JaaLSuS4URSAk5RcCK2m7tA/OOyUGJyXBhl5WmWtGjjwAZAzFxxt/J
4K8Nn6HL0g9w+pIjKRZybvrnPNG9w9pN5TROK4p2grh1B8hZkrvkjgBHnmxTjr/D
JpuXuyAuM8TOBd93jsbGfAtM77ELb8mdZuUF+lrF1H7r0Qe5e13aU7b9Eg8CcuOi
vFYSrKP/Fz4psgRe3KpUTPsobTZbHzqk4aujO44eUTZ1sBmrhGSFWBekqR+Ms+nf
CE2SFJ9Eo+TO6nEA8KQtdTRS2v31wV3AZlUukJWMzGYUw4hk9k8vArqTPbndIToD
mFU6SASPPR8NY9335H7MKWo/2NtOJNVhPHyTLBFOfBtxMut327eW5eFlS2H7Qw+K
B0MK6n50qEfvUC9I3RLqG/W8Iqb0NHPKvdb+eWm0Z6O+WSImctFugL8Q56r4I+W9
GKspJExtxjvU/m6+LdHIYbeE5dMTmyJnNy18E7+CQsptha7Zno6Fu2gTp7uzDZU4
PHvQZg4UwWMbcahepxgGYf5GOEha8nxM7P+Jzi3LQ8KRHO0XF7tTVDSgSohd8eN/
+hTBIGq/V+GflpuLQH1p8VNK0c8Fb8MCIrmwyLs+Pg5yEvdXm9uvQ8d2+Kky2RHO
qrTDCGQrAJm8uxK8hXNORcqu8A3nAqxgOUjefCRsvZWK9lAg7Lv7jGMSa1GY/iKA
2MmiZbyuvXiXLVZJP+HXLGn73mDMj1iEX3L9mAfRnMbygg8fST0m8TNCKhZGIVWD
Udz2RnWUsTcv6RWhuSBpbuSkAYvwjB8teSQfuiNi24QRkZR5BgL7wl2hpvXybklA
9ZbavtghpjiB0f4AAcq3uH3gv5+glFYrEqrQloj4hgKEkTElg1EylRZUapPcRqCR
YFxgBY1JtqWdOEuMFMfKz3NcVNDvD3/3AbwCB++k/GKWRyDdy3+mgEBGSpfe6k9A
Czu9cZ7D6CQmmiENGSnpvr0IgpERO1VflLQZhMhMS6YJhjTKkVd3MgI3wGDA0zrO
0+ehSaA6ri4Q2UAelc1ldQ6Z9PS5d90jdBviQ6u/9rglFhJuLLAsUjBm2Lk8Boum
ALydCzlQhfOmvA7A3VT654mejIHAE0QpwHIv1Lf5hmLgUkoF3fCMQo1GSk6XHpau
m5HTbk/+PfG6FZKTL1c89/PwRyTfl5OtAasM4GaSuhe/9/jWg8swCuWN3fSuvgpH
Jv/fpW8WugJTj2NG3Je06FSkB2SHSC/u5h5wu89UG08I0r/c2YwM41WnSLSlRycB
/FA8CAJUzhTlUd8iK86w2t9Hw1evK6JSkuJr78+TFf/XP/k+vn4cbzgmT6QXIIQq
XvF9Q1h3AKGAd1bCrz/FM0aiETuTHA8qigfj0xkfG+MK3w8grrjc6tLZQzxipbtC
ykLaO1NhTkIjeVdLUKAEtqjEFq9YOtiWgurP+So2G2MJK4sylDR1xqcyvQ5WGz3k
l24ny+oClgxg7wjXCi3kULLS2w8hzYce0bRvO01FxfIiZ2hboD+ATXFDaa6G0pab
2I7SfA/nTKgqQjP/5ZlZGT4PxJiB/I3C5+Q4eBDowe7ukXUUsdLx0DmwbziXpZiv
z1VMydv/O1OYegbRIxWH4daMPqlUVWYXujG+n96Fdvhkn80dbQ/SoDkS5ATEeaEu
tKz1kFDXVNC7Dl8HxnzLGXQRz16TpK6cFKxo5tWJ+wu93Y6LCsoCS+i29Y/Fhxpq
mqvEDJmEC+7V5ElMXAnraW679aLolk3IFNZmHSpEB4CC3RH5c+k8k7sJVe1xc7l3
f0FVj9j7tog5Re40rRkXhkvROgOHi1VhmceX51OyWA1JfK8n1JGkEWL5UBx0k8RL
xEhD7+oK3t1fYTjy738r2AuB6b2ZtWBtouC96/+wWEZeqGeFnYoZdporIh4Jyib4
Tjtjiw8kaWtti/htafHx6udXmEJwUZ2c4kKyB+6Dg92ay63qz+5hiYcw3n6PQcdz
0n+rl1ipr+dJAF7oti+c2bQg9XsG2CoRSJ4nGXUa9K0BsFz4cTXB+g8vdGN3ZHN3
VnCUTjYRmTNJuNvbO+1vuuHPv4YjW5AkYCNP6JrVeX7PkMtBVpYNl56tRv/20OIm
c+bsTd/3GliGPCt29lLEU94EUMuhNhRGH8S6eLzDsmfxb9w3/JwmRZlAWC0jLkya
sXTWF8UT0ISDY+BKgznhQEHHwAd/0QYox3MdAT6x7T5p1Qc65L0Uchz20LhS4CUl
68KUZaG3xtwRC3qZt+UlTtfoNfG6TH+HundbFFjdgbnk/cnvTaZ6PN+n3508ewJp
rcBt4UF7T45BpmQ3noXNe+E964P1zhKL+BbwQXpAIJa5fB1oEHxXl4SNt1jpm8QO
pcbWx+SRvJpFih8hdwxWD3fRdCQMJsBx0pxcudWvJ9d97PC1pBybk/J0fbi26+Ug
pQtSUdf470lmBX9hCv5nCrj5k3dGHk6NuuEe9Su/p/qnfixJZP6ocSK33OIWZnBK
6sd/UnLkHSc4bqRkP3+3b4nGn4PwBMw+inCuQvky/hngFAHnsgAVvcsBzqQ7cAUq
T3GMpACtqvvbXguZ22q2+tjs8Uq6YkAUk9QhGbREyA1xZaQs3/jytU6Xo/rdVXBB
w80NzHH62QDRaP2446NKjq/ubqjQ2NKJR3P/yNEfCr5SVa5wZXRtVBk9nzJ93mxK
56pPVOomyQNvDeFewpJwBCQw+ntKjB9fsjKF14MFn3RKeqOweDUazGOFygka/iJl
TpEN855xi27mx7SLAz+0wBcw56C2Rwxzc+q0ienclB9KYqioyqMV+1jV2iQq5EiD
qxqgPuKnXKYSXj/DJH8pB5wtIPtdKNWLg4Y/ujfPQ4/TsBq/00rpfAK75UHxRvVY
MWMAIpKygl1kcTMHnk+KjTh0c8Ar0i0gP9onRgsiQAxxjnYD/hc9us16wt5CrrSt
KcsBxe+izOUfjdiJjk1yhrdLxwqmc1K86ec7H4L9xG0KLdMJAM9zwpkFN1rzTsZf
MxKz6YJlNHIKXgmswovv8/2IgPoq4V1e1M8aW3JC3X7++J8P5zXagqOp8A78jNY6
2S0OIWYPBUMuUTojFJT3Y4lIaeEWrNBBjE4jyPx2TGEeiup0aRLKPa5Zu8uItgB7
F3E/IUcIalSRA96OgTc8BFvORpFD1NsEdI6qjGVqPLjycga7ss/q7ODxpcb4aYoJ
se8hjWoHygg7TPnekzG+uCNDEZuWZ+02wnjO8MidN8nY6tT/0AtHW6d/g8QuhkKS
bgSGTXv1ZU0y5Sm27f/DUgagtdM0exHqffsEw7ES+o6ElXmtJilKJ9clX4FJO2UR
ki5umAkXW9wYO3v1ie6CHbHH6qV2D7ODGLjAB+fSSQX+xH2TdYez7GMZ87vQ1+t8
fWQwbcn64qrtNptKyE5IMeN4J5AJv9KJu0B6G7uBoUkyYQQOcigsBnGBbJm1sgdQ
MIHSM0b09zMbHcRCOFfsXtDjCGmqsE3Oyk/68wZXerZqowrDStQYONUw1/08oVfY
z//fN69w48EmfqxecSyHRBaSoiG4x1BvdgX4ELOZgcGxnSriRDdW5yzeQ+/Kok7e
EjrgqFp79YXTHMHxcdTJ9jwkVEoeocYp4usitNSEzC8drEG4BmkMtaeZpr0b6aNQ
a2mXS1HkKHFTWJWRw+TnFNejcUfzsfwrK1Al1X70Ufp9tggLP0G8/tFhvB3b9zrF
6co3/QSFaAJlJbJ1LGA3y8pfifH1zKsmynh6cBCCz4AT056LKT1Oz3W9TCVYr+3F
t82YmaXe3TYdlv6Cy3hYgEn3yQhg8CUpWPGNIyhwXFnC2kO+btoW9ApMpZPfGDEG
E7REwyh9OXHBegvhneJk761GHctBwROBjhm8EgdxIzmBZq1goHRKqV3ddHtEzBNj
qY7vSKZZ9YM+EVhyGve8+l7RtPP/m3jtX988dKwIy0kiTu5SjigShtamwY8/uJ+n
ZWYiT85XvraaAGxMJ/jz/dUevoJNkCxmPkr+c3WOuqm9YLs39geKrMWBckhIneF2
LOuLRI0oIRg/Xwrk3l0sz9uJA99ue38k6xgVtYBEJ7DJQFmbNJSohr+UnulWv86B
w3gIimZeoJhZZT8YoEFwT4Hzc+VreFLKuc2GHnCeZC2P+cJFs8QRucHjLW2INxUS
UPkFEbl2X/toOGhKunaQa8gLnu5nGLIY+3uj0Sec4qqnTijJK7Tq/lwZ/BXGKWPh
8+ndEoWMp8H93O3vVyZndPA7UmEEQBrpETGGlP2hf6lKqD2AYS2YamyhAralkWmF
+swAqNNqgAspCOcEDK8Mg9hOvpRh+5OaKnIkW12EIgXZG6LTxfo1MG4N25jrLSHj
usNqv5MguxHx51D4hKY9ax6z/aNIWfp8GkJif1l3mZNvbTp/CQXRBevWIHO88LNf
szH/d2dLA3fvS5akiNPVxOdEgZcX98xXVHFOjBujHh8BCiSbz1z8cHg/z1Hy+K7V
ljmmqLPiAbCC/tf4SqXUqhVLt85VnKgqLYcW4Y1iYF8/BLmA2I26hNO2m5BCuT+S
YwWzBPjzmL2j7xuDLfLvlvs5IjviC3d0m3oysXfr5W052hvxd8N/yiyHgZzgrxQV
Pr5fY5iBg5sXr914WglrEIVdleQO2cTnCr23MDqTt0A7ekwqKkbNfPtUAdcBgBcw
ojJqJlht8JoPRlYluZOM8Lgj6M2V2bs94dR00ufq/fzl3AAInbXEDFB1es9YBcqW
5BGv6WOj6fDyduTmrhPgUUZzNrdh2+705jv22J+YLimsYywILhHburOTNrbWHl5Z
sl9uaMm8mV9Okl7Rknsl9o4KGmu4N1ogDVZmsbLAT+7iMVtWfBlvRKjpsqjWML+w
N6hOicnAYNcPoP58iL++zXK0+3VUb2S8/NwfmXexlGNsqpn87fhANuhvdGc39M0+
28c0ASYv7DGHTZ60CnoN4S4LpeyCo/PKeoFZo9ncOiPLsHZehx3/pO8gJg2Uy6sr
OKI0w523x6x4O6SqTmHClnif8lPLYnNon0Z4YswVe8a698IEh0bM9N57dmpJ4nKd
Y3G7m6eYqD3lvf3LyC9wFg7pB3a58cuf1RG2VJQiqU8geLuDynoWxwNZvoq3zDAX
7qVWpbZR2NUvArkZ0bEtDgymq/FK8BERSSUYYRk0Azg/TOcin2F7W8tcIhADVr7z
NsPNpRfZ0tTCynuc6cvT9SQRXkAFMv8DDO0jtZEYQ+ypPkJAjvLbqTb/fj6apPD+
BxTPj9Jq5gGqwhaSpDeL18jc3m36qCZwWikBEZ1CuGSe+mdOSB7+XT/kUzBRZRxL
qMkj8+UtfMnQD8DiHt47tlEwOA2GzVvfJpNPeL04RcbhYsLKMzuMMmYKA8CB6JYA
zJoziKhVcfUYDD0gmI/m/ogK4Y4rWJ2JoB7CxFlOYu9hmaqDJcyXu1bXNKCL3ENW
nG3L84xulMPK3DkGNzywebrW6aTF62nqT06JrhBHyWTXCKVBxCrJh8SWwQRW7KWz
hgoaJS1uGrykcDScAAUZg7jbtYdAo8sB17Dn7T5GdaL8l6YBFosLvkNM8ijePDiY
3dQsJvQB7hYxvu5fDfnI9EBReazcpcgMDoYEXW9MMcVdi0JML6GJ5oQAe9ZEE/vc
NtxwR5yRzNYs3P9VlNLbJeQGx2rWwI0nklFPUBc7QzLDWvLysDcA4Q5BBvD41ACX
RYTxyW8eDTo1IFp9xlGqWmfTXIeUoP7p9m3oqtRHdIKIonfIBjUT+Z+RwWCQYe4f
NJQKBMYIaIwReIl8HGrwNANXscNXeqoGYott4ajtpkwWB5sUweVDBm2viez4B0PX
mlIJuNdqE9/t2UXJdijzem8WOY7dfT2THq7IoemyLYm/ByQflI93t4yIA2s+1lzQ
CZHpyo4wssA1cWWzu8lKnGYsBdReoDTs3Q5wm26h35ayQ5Qu//YSfUQbFVpPNe8k
ybYosS24oY+/Iajd1kOe3A7gstVx/gWRg+WCdNVCvJ0TGVr4Yb80Wj2er9nb+CSK
zvsCCHWw0vK8BFhfZJvdYnnn9Yt5S2JBdl9kp4iIgIPIfMnxKSL+NVA6+bAKak7m
mqcKqGohyc/2GJ5yJdsPL5DC1AWr5BSE1k8HH5NZGag9iSGpK6zmxYtAs+iXXmx5
vSuSI0GNZ3P1fVO+ULFctsS+irs/ulFXW8/janglze5pl9JGPHyi8H/QQ46Ta3KP
SzvsCkiOEaQHteoSngvvgQX0yyLXRwjm+xaVLdbbKUVzQ+f/gC95wMIPZRRajZjp
dWej7Oz8nbwTK25Ng329s+ooyajytwQ3YSkuBRWaJf8Ms9uIvfbkcQ/1XuxqtljO
Fl/qszXq0MdNlheXJCprZov/ekKskueacTn5VqFAAc9WctT8kGbPsGlUhuP/k8+X
z0NQOnllrRoh18RZmn1tLiFo5qrKWOVaTyb9jZH5Ki0SbqIKPPd5QkG4QoSo4mO5
cagoOFwWrWw/fEk1/fPWKkyc+GANHPnAhPRcXwkn2lFt2p9YrnpnhlcNw4S7QZrT
EA3oD3HDZKDhrXTLA+cZp9YHXJNhe/N+KHXcZkEFRAd5b4+i53kEszniXo9Ff6QM
oouf2hLvJjsczaDtFi4yF8EJuRcwgD/7UEbbPwxjYwSQwczecPLEA2joBql5YfmM
PaNtc7BH24KZJuZkFmwmlk3qwDjPik7id0SLSshMkDqaLtUj/hml6nIaoFH9O7jG
VP1PGP/IogoknM/CO8bLXoHVqRbxSR8V1vbtMqqfmk2EPWqqayodc1tYtSksc2G7
qXGZJL4D4TfpiCgMo+Zi5YAPj8aI6+Dxu7cUpJ0DUxtoORVHbIyW+rneIPWmORGA
JMvJgrScntbOwip4EzkZ2zVMNcvE/beZtDqao9QfGIBOH5JYfl95XbkNwo733fD2
Tulmn96CaCrmqg9+0GF/BTfjyGmbxiThcHImcDNrNG6JNroIYtMu1a4VB/clBsP8
V+gRk/TVsMLt2BxusrlCYc+mghCqKBf0qH9SfVkTLceDOlYrX0mEcYrJLddZK/z/
kPTU56gO1sMlCoSOG2CEl3RpGfjYAS8CSKOCEPq89ll7VeD/yZP0EPEP9a0uTDVp
QlCjzk+HbQeL2a3+jVfxhKS+HxxhmHwsX62zmfnIvtrA91p9r3M6gEEM8cuyrE6r
U8Xs4Y2CAypxcWpxdGPEHjLaplU7RmGfdDe71Os7ChgU3aaQjx5BbqVnePxhyGgx
5oLQwMhVTQt35XzWBi2ZCEyGk47dae1lPMyURmUvml7tRCQHt5RgSmKXJ6qiyvyb
KM6tqtqADHXzVG2eNR8ZAoe3XWwwsS53UuRi2lz5672EFr/ypbpY+EkTaTpTJYDH
KKKyPbZFAXZ9Cxa/09Cxl86MkcUpj848LgdhW6WqArQ+vBKZnnPVHNOjXv0crltV
7IK0xwMYA5qGwrz5bKIw+EXIZA7Mt27mtPpfeKtt+DvkguzCybvFxpdyECOAx2Cx
2u0Zz8W/EiA9oo4Ml24LYzckzQ9yTlMek2rGNq8IZvj3JtzOO1EkTokdQ/3NT6lb
QEQqM5ONIcXAWyXEFzE/juKhSeZuY4w4GReouCO0vVmP5jhmoarFBADAzWFqRrJB
sMSz07hvCT8KXZ7/upS+WCaJi0Zd3eamIWEIzj9jB7eDTqirMSvd9J06XIrOvAOl
bVoGCJBpt+NIG3eyQe35QzqeqXiCl+CvEuEOKISfiSofROtLqVv08bXd2JFZlnGq
KQEN6EUZVN20rEGkHOWAdyN+l14xTbrrvwurCE+4FolXsPQ3mumeITS0Be8WmELf
c5xPQ0iZAHbg9RXIhIzU/l8XxsNyfNp+COi6gj8lYzWt1SzJkDEmkuuip7RWk6zH
wVsKDT+izrFBY3mwJikKVRLlTGh0EAhhThkTXfiFi4hsrmJszqBTZ4IW+gJw0oQG
0YvNXOMNvJ2nLQI9Z+nNdajxRcgtZPR8M2hdg6T3M5GqT3hedKNKh9EbtfUpT6jS
tIsnEy6i2BHdo3x2MjgMBMLJskFoqzMSS76LdYxKXAqBh8N2RGQf/mfTaaM6+eSG
7ldBtXwaQ+fB4QGzhiD3bMqfqd8R42y1nddAbJzY8nSRC9/3wDEw0Q3MHdIOVeJF
HL9csPIfQhGi54KCGcTunPW4O74PUZRXh2/UX/XiTppX5rnZfnUiPxbZvjKyjhkD
W17hlNqc0MAtySch4RxAoqeLAJ2wBfVQhRTuIoZKl5oEpJs/KDZB5F6uQi41gJNV
qjY4ynqYQQamXftyn9LCq/tMrkqJ8X4EUiJnsdll5uZsIOymSqHxCmyV7Agn9vIu
i8NIanxU457SUHIhTPFqWC5UrpAXRFAtfT7RHGoSwoVXIXbo5csCBfVMtlcfsINb
VMQhcJXC74sQxBzuLn1ymU8Mjok42e+OlliUOFxeewPQwIeziCU482OW1nFGSggl
R+gvba0pGWb69Zq+EFz2hLvjjDTLKquN7A8ADqjwAf20dZC1wpW4clKL65R1dc9c
32QX144FgbuahoyziyWvvprUz9mX2sV8OqFQXeSMV9x9ImeQuhjqftUvCyBh2ER6
PQy1h0CcV7ax67xMojQHx2MxzGvWkPWyr02yDMVIZ2KzwQPQylvAuAnV8u9/sfms
aTz5+SQb9lCs216lwfWMZtBDmd7gyiYEPUiyCqWB7LTd1ME/5ZWDshIBDL10ED9l
fzSNsf91Slo1nymCi1rjFEOjspwdKLgOe3vHWUf2Bih7tB+GExnR4CSdHKUabLWR
z5CmRy1ajNzDyeBBwGTmQAeBKGh2FU/AJBrOV/hoXVbBs5qLD9iOhsyFaolXuBjp
0lQjjxT6uP+BeOjBXvx+219okx8ODlT8vZrf6cXyjfXaRhTp6NDorkeo2hJfWYez
cnWX7xrIHMD8f/YGlAIl1+D3tTZsHQLDmTC+DQUBaDjYK0e+g+e/WNRuft2JUa3h
/y+YwrV1U52K9SQAaNmNz9qB05tIMvtXdpvya37xiI9hB0ruP0eluzRSu9j1vRuV
8fch4g80eGcM3iILPNxo+W0GZOGHriDxavF6TsqeUU0GtoPM+Vpp5xEqMeovDCq2
z87C36RtBoh3Q/l5XLr8Xr2a1XqzzqTjRnnOsUAEcZJUe+SksLnGIEj03azjX6N3
EyMPQGhoNwDHIOQc/xklPxBCJCw7Iw6sKZt85RDq6+IzDqC5opffNGglSRWkwmWy
y2Ldt5eDhS8LvykVbU36GSpeUDNCcrPyy82NyD6hPF1XE/2O9HbPt4jiCqXe7/WA
oi5zUy3MIjqz4rpXwAr1VxdH6HCmg+gCpphU5k5dT1B6XoeEdzNVJLfkOSkPI64m
nqglJaxmJJLQMAX+9jBaOwSO85AE4ai7S7bTJ1e8pvD2AQEgRCWRxbih9vk349qs
gvcFIoLzdTCO7kMihCgzoyg1TKs0s4oeMMWZZz70uPfVyXkF9WZQK0hNFcxcT7Wh
sAHoObk54jOa1t4fr4qXAkOUXo0enH7WV6qv8dOU7FzizOu+RM7G2HSD8RUrWTLn
a8DGwVsS7s3ksyq+xYT1Be+Qby4fnwTVU0UMLZfJr+eDQrQ5MyibbKmXk/7XyoLb
lmz8GASN8rip+HoGXceFdGFqbiJD90JK/eYswVPHz+/pzs7euqoVdpLLO+jeuSOP
aQsaiFmE1guepq4FA57paZ5JVtqaFvMdJdDzGiF7ukNfIadm0lVeyGYxMWiryeWr
SSbVClFNpX/GChGClr+1N1ummnH1oHycdk695y4lPUXgN1CzD2dKdJzBKs3iJLXU
VdQDW9LXTtpkPwW3GfzmKnUkXcTBYGtTn3yAJdqsInREWTm0yvsj6gp5L9hd/wnx
ub3BDqvnMIEuSekmBkYWBLoh1dQEB7iEZ80jy2CMQT6nIg909sr772E/NP6GR2IQ
qM72EtuQRYV0ECihLBUVt6HlkH2DSZTLRU9T6Bn5odVLLYlG6GAdJnlOO4y4oji4
d5sUw99OwdwLvyWSFFysfPMlquh8vcymDpfAzDJWDSBJB8JkHmgf6D6Yl5pHg0B8
EYjskUeiw7CipJJ8fWSt+6+70tAQhu9lYBEQ1Gb4bm3iP3kuopk4f19+xGQtfBJi
fY4R6J3YwaqHGXWBz+8wNCCuL/Ak83qTcB9c0NBdjxCj3gC462V/Dt293lkpR25W
DqiEJRkDuhjjz/DvH2xFGJPBgdsX++61L9KwF1Xm5TAN8wWslRXCqg/TufszIhT1
PUG8HVmkRt/1CRNf3oxQEtyvgskKCUKmMJsyg84M5idTpJAX3zYSfZKer1dzaW92
HQbQ7gNhGeVVRWeQw5ZsGQdd728mmT8LT8KXO8TvytLYpxbcj91kK70WlxihyNk/
n8fPL8R8fw0NjANv+ZKX6k44M1LAU29mtFcCkRYEZvAl7Wz3o92YIooih9D692cd
gv9miZQGCoPShyNicLp0+FoG4wtGYebwXygEfundKTbyq2aOVKwOUNk9cTwSPutc
QEvB9yccD4abC8Bn23qCL2jZARhLd44+FRh+iN94vzs4f+6vqcCHvZquHxMCQOaJ
w4BeK7keQO8P1Hehi6oL+0ilQ+vGEsZSxKSDrq1F+oqjR22Xoy3LPHlxIYM6EhZt
gNenL03NSuVKGgLquChl6C34GoFLtLg16Srmiac1iiZyNlvQMnoLTDh27i9AH+e4
vTReESfR/DvfIiC2e1TJDdakgpB3TK9TwAKtRVFRPbXpNycg8Ydcx5bpLUe3tqCy
UjaM/PYmx4LmiHNzap16sNDezhPWY40kTuSyc1UNo7HNIJpaSQatMLAAeEuPYlgl
xVUCWi3AQdf+bSGn7bbTmrtHrguSzn5W2hcaW6n1JmTpu9Pllg5mf/VC/0iqyyjD
7bK5+PS1AN0frQvggyH3jvZIuweZZM40uYbK9rUyHlyYAmaBvbqKeLRn0coXNTKT
zVXJyDk6Bjf3eU9vKhWcOFyVdtx+onr0lD1KlcYHilGc+icFHuD3LrpU/XzwwSrC
kcIAn3VLROLxndysPtPVREI98f/IfjBisjGzFJMyx7LeIQfPFMUB2BB6SmpQpRae
oi966Qe+y1GLFeHgIo+WSbjSsaWPmO2b9ym1vI0XErrqFS6NocAgZWksdtGvfgtr
tXXa72rfELvzP7EJdD3J96dv936rXHJFaPo0jOCVH+F4qXUKCj0ZbmjZa81j4Tce
oKm3uyfpnOVsHGYFgY+W9MsP5iyRZVtnBH8rJyKVk5P0dT7c3vBt4voXS8Fb+02U
dQOvH+6DhAYdJjiAF3JdK86u6Gh2RTYIICNpcR85XjXWVSF/eysBZT2XW61S75Sy
wCGHO3RH9a63jp2cvjmeSZaQT7oN8/uQr+CpE7EBN3P+hi2nngrFt+pfexyXeFT8
CZ1QjLSZZddnHRbPhBsAbhaYlv6gfTHvvKjxaSeuhHPmUs0qBwzUasMgOn2IL8V9
0FfBF+gcOm82S1rBPKrNODHrPXUSnKoXvidc7i6AwbBq7LtC5CBC9XvsI8vEn5Fz
OTmrkZ+s8+VO5Jt+B9CIvKrzn3bf20f2+rZxSAAjBGXTpM8pPS1YAkTPGg1qoJ3Z
zt0waDLzFtC5dh+jfHyDO48x7X8BhvcljcZO6grrbQiKyfweOJOvoZutE4bK+6CN
wcUJTvNqoz//klSSIJBHyJoM+9cwyii5zSuGt50q7PTFlib86TFzhhL9nsJP4XKz
a6+LCBSwSIzmPjHEjv1DL/kZyUrR9OD1M0BUONzxZZPBB1jMf/b95Gu7JsqhK/49
kS7StfjS0U8h71rN8aKDzV0wGhwTRbYI2fUQcgX8Hv5L87VMfN2y1WoPUI4P4VLn
bIlTjjEQtjs3UotiF5Akf4PZONM37Vd4RHEvt4YVqN6I6vcGInUxQpAGziC/uHcS
yxHauy4VsHXwQb5rFvLvmX2CA5MVCDxsNJ4LMkSbhhJw54a1W37EGlcZxAHsHBBB
0lJkwyjrzynRgMI6qAPlNd6YWQxED0uv6ucyQJFPn/StrdoQr+STVY6mWOQGOzUC
LU0VAMc2KkWzXnF8vQ5KUq/DP0rxgyprBekv4shQS03gtTr+kQ4lll8jMiGzKd3c
DPwxeZJbLN1YXqLW6KTYhNs6JjoDDzfbj7BtLh0m1Q6Jhy/Ljfi3BHKfq1+NxPrj
vM8SYdVvl/Qm3naN3R8+cV1p7Hw4wnMtmvZmU0aRQn3gvGLGMP+zGzrsP4pY1KzX
/TyxyDN9dVyDs7KIN7gKsKmI2BnH7TtfH1KjhZzqG2hi4IQjC+E+gc4BNECcnLXt
7LLpkh2LKZ5taBY2PeWh9UpyWqwFRr3uPIWcD102f3tNgq0IBUzvwT3tx0bR9+7Q
6duULPCiI9/7RiJ3NWUDGAl7rHhnhJDOUUTq8ELNkR59WEv9O/IuIxPFslheTeNL
UvcjJ5jr0UUtrFFWacJ1mQaPF7AaZBTC3OoTfLXWkGhvr/ChIT4WTH4aAGdF9cwU
c5EzkyxzshfiICjIt4+l431YWKZnOgAFcr+vdAjzkBk9V5c8ILUegZeMMlccNq37
aVNEAyr7t0uSx9XYo9sqwwnuNRKCliWF5+szjQAQKdCCD7Jucl9dK6ElvXIzHCUY
vkkCjleSdSV4PoAuPGQAzLqlPFB1fIqQq514px9kVnUQDEAf5f9ZYYguRuw+Sut/
F1dJDwVDFKN7bbjyXFYu8iqr7nME27LuBPpr5tRu1EUoLxSVG8N7Gaqkf1rl43IJ
q3QoowCx6TeOp0Zhu74CuFFnecIRwpLfaFOufaGXK8/5Hvq9oSB0+WKEhPkCowND
PeA/Z/C9SUb8UnjsLH/PEbv8bAnlmiigYkUfY0nb7RLCd+0LA7KJNRJmwzQtnS9d
UwOTpth7b5Aent4zwAqqkEQxwXgFUcNw1ndUPYglWVvE4+Kz6KJJ7QCTmyC5LPyR
eEoQSaF0/aDnE7Fb7aeg0fuCkGPS4xdOqKMP9lN+Zl3aZuY+KN+KXSPtPlXcbpPf
6DzmIRNj96SVTDQ7s8NMEvGJ27HvDMapmN+NtIayfckp2g7ciiCq7g437CC/P/Mk
in/NdVkgtRAgqkx4hGon5IfmUX+C7yfdNRh8OeIi7o/ZUQLOpcQxUAnB1/aGwZeA
3DovOYLx+19TDdXfwluedqHxkNDc2zmF0cTZNBdGTpKU2r1QFlqeG2flO00XxMq4
1gH4wmD81HSD4FQ/jHJDTAk49pgej2o/Op0Dzto7X3GioE8iW+zL/xrI3ofXD/WC
F/pr3iJUPsEniiJL8iJaVTiebCoNwbEN8wMFPM8VhjXQU23z/lOcSrZXoYTe7Cn/
jgfybZgPqq+T16AEGtLcyvm5TkAZDYYWaL6MngbdRxpVPFws1A7lscjuMOMqHc+/
LkF/Ejtq27l0iH132TPNTRfvsOwPdmc399YBnQddMl6fwG18hTMATVbqkXe4tYPq
qfX64zOA3Ttt3tT9N6lez2n1tY+rjloxgrIcmuZO1YqV00aIoJmz/yE+irYKRQ7/
6p8joKHvjCjZ6+JtGGmKTVTsg9w/D7wpy8vVoB4+jEcsZCi2xH+ARBVkmVZIrvSP
VtmLzdJQAVusDcvlFzsy5vn2IMNZ2uLCw1yB2M4AcHHth+t3VU0pZ9TNfZWP44FP
j78wCYpZpyYM66AJOC53RFOQ79JHDhPOIQVloevz4d+k59cvYS6xEL0JAH6pkAYK
vfa9vPZxtbTfhvYoLRcQX3u9sOcrfqn0lDa78PJsgvTWkNpxnoVcqrzvm2xhBVBk
Cr57c7wd+UfxBCpJ5tnC13Ne9ZdTkhxQ1A/a0phsvKIQDOCSlCeteVQuU26B92yD
MuXUsywY2zaXxhpqnSCht8soE7CCv/o1wU4SDy7LkUT9XqhdQkM+wh1ZcfBM4e1J
LuueNXAsu/nmStYPVL8IDr1yLle7NTnnkpsR0wJoms45vZVbsB/2MSHkQydMxexy
RVDor6lCjkrqeZm2cpzBfFa6EWATd3fszX193XosOn2tjIkebsRszfZqO4eyucMd
ZDCA3LOQs0YCdk8epl2CaRBU6BceTpTfqevcg0STyhPtL/jK7GEY6Sykn0Yyxvlf
cuoOnozrVSPy0wfSubDW5JIb8gYl+jHFwz0MmHJxaNCNyx3hwOQeoV3Y8r5lj9bQ
iP4S91fbrju7OzBn3HbHDqkzZPXx8pKvWHVzSOhuF/WRldPPTphj+GGyFUcIr1Fs
xieXIRUr+GIQCxtFagwDMCN5WBOA6go7sWcjYKIBG4I0trlTuoccWkDXn2m9N7AY
C+jD8I3X6RPEV/IyFJ5NstGHDswyInGrkQayeKi2T958vgka8c8baEYIQP5XLP2f
lp89ONPtaflw6MQ+lKbGiAlNrZ1g63yrfVGyGe+uXSY/G4EFSh9Son2FwqeBTKJA
A5Y4fhXb6BOj2+P5cb42jqB2dL9KbCpyORedDYwtQMa9Ui0I8LZlcgXi0Fl1LfNq
tBA9Eg0DKAsCQ1cqKBFpVQMMRDwrq9NZRgsMvJvFJgjxubUAGdx9MQ8rkC/dUDDI
QsZ0PbSE7SHxVDn+SoZSMJkqafI3VKWagCCRGuqhpEYDbjihhWm/zaoC6zHCp7P+
nU6RA1CmFm77C8GqShzuL2pVy34O0GqrdbldvcX6BJ821y6YBelifnaiibpVYvTG
aMqTbINMXTJn1OPDw+OTctLsOy+KadxaAvdqtMmw3oBL5ZC2XS10JviXjLfjdIk8
9OXQUWc1QWjuYUhKIRf/8qdbGVlJplf77DVMU4L0yBcLYZVEtkaZNif9DbCrmWSD
by8XSI1/oEU7heWcYXcgH1L/TByMu2+GQNO00KRaABuTqZf1WxdsS0BFhtsAAdFo
Lo3pBzfAPw/863k7pI3M9B438wWdqSq42O9SLzZ6NEGYNY+bE4C3B1KbUQvieeam
JujCgfYeGrK6lC7KYduMVFF2PVKVFzZUcBZM5NeMN4AjjtAiezUsCnk83TCMZft6
8H7MiysVYQcKkHV1AoEg7lD6Z4O+OoKxDJQeiu8H4+A7Ojl5D13rEMFFwMxw5MwP
cDg+PtIB20V4+ay9rIUcsoS1Oqcf2FgeQghLaD6PPqI1ZGE6a8L/cBSC5AuhN/BZ
dBFpnftFdll8GPtSP9Ca0mlxYXMevwDv8dvuOoI21aeU8JmfBe4/luzvPo5mfLIp
0+f3FdqfF0K2zoL13lUaYMbTgz6wAdC5h+uller/z6V5egsq0+wG2lQK2NnEvwAR
mBkAhHIBHot0eDefdkZFi/2/ALbkEBL6hZkTwi0DfT66/5KAUShicslrXEqOgg1E
rkx+14AnEoBGr/FG/JUlI9wUftBRDW1R2cQv9qw0eZzhD+5aITAGrwfUlq4dJDWS
4cWpN8iPB79L09p2sEUfKoDX5xKiE37d4pl6iKirdNTlQsYKiy6M7O3TykQUY+YH
Vjcm7yvEkPFLZrZPr0/Xfer52rbBwFbRxEJpVfn9b29jO36l2l4+0VNSzwfhwn+I
WFDSMeaXQPLDgBGpLi0ltaItKYo/TpjV5EuGtsMiBfAyGXkUzSGlXGP/9Z/x9SMN
E7X0mT7OwUy+aiwTD3qD9sY50nlhLR4/7FDwncy14qiunRXFv1V3XPlqZ3b1SpQb
j3/TFp5VR8LdtYCDTTBQVVyQVPeGGGg3LsCtCxczwNZoF5f3r6Fv+1tcANplXZtJ
CcKh5ykAv+tLXovhKNUgZqPFIRLsxuKyeAYzGGRNbMpEFTxAev18QTUw+EUSEZb9
7EjQtLjEnbVm1gZGYohvuY3Aq7anfWsYodEtA4y66NU6xNT8r8kaf/hcIeDyJ1PV
dmDOk1F4S6NtOH0bE7o4wmeXpWWp9IgMp1OVhv/bz/k0N7DldAgDqtgFWAMfb8F3
oZr5U2csbIZgp7zlDXtelcj4RGkCsHWVLNBZTjLudwtyj77jlkpg1R74X1Azi0T9
vufm4mduPP/IjQjaQK0pWh12Tg2C3Vf/DWD3Xf2jxU+OTZ9HmgM/mEhCmtkNMRel
bbnnb5Ux3aqvQVsBnJsJG/XnE2268NULxwvpcaYBeZXAPpiBdp2hNX1etl6mDaAC
9Xr1rhpFWn+8cBrgbHRepponUhi5Tqrpw2ABMP7H54ylg9gucT2uBLyE9Uu4EeTA
NH91/gcD5hVAsHekbp1Q/483zZUYL+3leqnn0F9F3auPNPpQKlCKN0kxN9fqpEuh
BfzhT4e/kClYgAh8oHhNhRt2F8/ZJNa0H8sCZOHNMQABrNDx6/jtIKyZ7a0CpmwI
sraatCd3ifjQOi5ZuW18oR+6ZUCk456i85GpKJBfM6E107XNznYW+wEqv5WWmeoK
fgyEcJxe6lgTIy2yLwGz/HRMPonvl45wYRxI29Siq4mtf19EJXx2fjl99E1CBRqx
x6pILTxxQeiC3hQ76FMv7tlH+m6C3XWeegqX2B50Kyqt5CgAaFRP7qraROoAYFgS
EJpAvNlewwxIeOk5MflaNWHZRGF2ANKNXSSmNaElLYoYNi52TTr4EKROjBmH0+Ds
sstpTMhiuWR6KIi3vhADrk5HgYI4lls+NgMh15wM87kVoaNxIeviITI1BQgDyosK
wjQxLwKrtng8qYqd2Or70ZF4tGgtAgqDkYqcK9RJ91ThcZoK9/Xfu//nfkWOeDB6
Efv5XNwo3AaJyEzD7z65PycApUH4s0Z0/jFrqLifgKlTEXE7K4k6Pb9+/N3dIj1T
ynj7ho23Jh0yBMVNrokfV9mh+w4bovFRsIVWzHJbl3ROrDYXG6fJ+oS2Lv0mJTdg
8n+2C5wMy0tBKqYuh2JC9jYZ0C1Llgr1kxOcGNU3vKY01rc15PEYod32zy1d7N9R
I2Wm49RfcAJiA9i/bzoJ41uraqWB6R7sn/7Dc8y1z9Pf8JYkGJ/cPykV2P0YLqao
VOo6QYVB7aNyQPXSsJVfsViNuwMhSzYgDG6w/ZtQrYCmbuJIgtTXsI35SjAWYN0D
hg3jmV0DrodGrzo0rPVEJP3moJKVuajoBVEoXhhWJj/71hAdtU2XGwYhzJMEYUCD
dYvlozfKLp+oP4REYhh9WntHKcLJRICdhc15slGNkLSK/sfwpVA/LiX7ZLfMYWrp
CrpP0XutIjHIdmNHsrcQLmcj0EaxvU5QN+ba+Q1Vw0PCvKW6msNX+o675qd+N4Eg
rqHpSnp8ZgmM5SHZNvCoY1ca91nwE4ER22ZguTyb0WLxBQdVbkSyD6iXZx/+V4hB
wJpid6myYYDPK/NjcIgWAFDzMiv7YBF/ydXzCNVThwTUbXV4iDBH6oZKG6SdGc09
oNZ06aeb0LiL75HwDZxhs6aagsomjSUteeq1CFUx1eP7a4+PKz8+bH0XpeG/UiqV
PFgtD/mO2KefZWBOLvdNC/U9UEr9xQrHMs4PoH4QJdR30mRyYRLsLsXXd+paj/EK
nzfxNRTsjU2QaI7Eo/esjImKSgeGmx8PKPi6iHhbSAmcSHYrlnHkag5EiN9imoiG
Xy/qeGq+KqvNPunS+NazvYtQnG2w3TdiOFmynpzZ/gesMjVn4CfSWfrArVQuA1Z3
MppB19uQSe1LQCudkeXc0sxBM0Ogz2ssMhT+j75YILq8sx4OSblbttVeP46fLEzh
IlqUTlZSqPNn8xGmap+AaB5ZeoZjse7/ObniKr0AkR8uEKeNUfPObGcyGd028rTc
8Dn37GACoZTMa9Y1FVAE45kSNRR5sUO2hxBc1abLfhX++fndQGZB5Is5PvSMp4wB
2EwlhbhFi+8HgYWRB2xdv/xwtoCErc58DjcDblZQI5bj7NCenDdSr/Npl/6cUC2t
IABf4Ia50iMWnKROzFfHp+pa9urZNRLVxMRTQU+6wMhSE6223cY+BIUtSaNR5XP4
SpqvBGEn0VBCvPcdxx2rsgGMYl7nmscYgVlF2/FZHJnDs1fJH/bR1BSe9A6Br8wa
qqASZOd4EeABjjmvY9tR2KJKGsHfzEl8CTbPVrq2stsih+LtOxBt91FUPyCY6A9m
SodYjpQ8HZse0dzpwNEwYrV4oUWycXS1N1yArJ0MjaK85UFRvcMQ9HvuPE3C26oE
RV+oj+uw3VRak3EWyc1G2M6+tPPFoIt4QuY6RG13hBN+ZsA2r4cP9YUsqY+++e0i
uA1KIigJ/LMkUp2+Zs5U1dB6IUeEktTIBwXLBLitwX9aLKykrRADYGYAKpn7hzZw
xiTXGiTX055UVJ4e4w/pMKrrHsgMts7/5VjPwxW0JMxl1AHb8jbUhhHYDfVfF/r4
6jRIAxdS6e33srzNJ+s8J1M1mfN2ui9X4hnbiuwn6dd6Mo2R+1/VG3vG5TLSDblA
Tk31LUe7tGE1jIzsa6hiFsKkuG2MJieYFFH3akBTcfhM/EpLoQmnv8Aq8RYTYLps
OWT+lnOnJ/zI/3gDMGyR6sB6Mluw/M7mExCf/VB9o1YzyqeQ8MWd9GfjK7KD//4s
OOo/NU2qn4iw3G8SmlGavylTfWZUcrkgVTqcJArfCqB4TRgYc3VywJfJR5BIne5f
DBcTAj5sZKASVa49aBFb9n1ZetHFIq2dquDqCnu6E20976DvHVfmDcmJHzOCf+SM
g695QNmFaj4NQVIFNdG6rCi/RYUmalKj6Er3FiJbulsFVDEMo+9blBHxTXfGTlEd
PM/8Ixi0Xx/u08wj7m0o+JdvQ4a3ROGGGzioHbR1qj7VeLf4eo9+KVydSWdRvylJ
jlJ4Z9qldheT7xdW/6MVunqXQpXq06kllgNvvSyZaFh8rPdzQa0lMARvbD1SNj4k
96vYurObjoVY+d4GK5vHajF0NuJ4xVqQL20CIrRQolnghRgiB48pK14/kV8dhVGQ
jgB00qboAOh5grjW/7oabIqdOfu6zDvahFm+MnzAYebyyQ6T6zxibCZoJ36smuEa
FkSA1rHIEIn7ugjFtE8vtZuvJ9TTcnscGwzBCgx4/b62ZBOAQKg2Vp7vZatT1N9r
kCp8tSu7dSNkzhqVdCqF7t0l5l4KQV5hc6kT33G4KgSTS9fx4XTr4Jw2gJL41wbz
uhb4A79wc2fYc+abosism5brt1pZIaSBw1XfWu+VqO8WpLkLAvOP4w08/on3h95I
rIGcVj2Y2azwXnfzzC4PftTjubcB5bGE47EMmWKuPK8nVx4PwdrNas4oI5uxzP2+
qk7hoHLvkJhN9OoF3gLcPKd+vyoxB+TaFkHDGkP1pCBDCcGPv5lY40p9bbCVsBNX
asM6RYSoREaukpPquhlV+h70wxaI6Kp5BKy7jh71FdfJIGKd7/1f6luC1dAGBpuC
j0ECg1jW8funjdb2ZT0D602DOUovCdLGIkYJOwQkySjIkKM4JsSp6BQHLcAdgAaL
kDUkA9ZZ8cMjXPlEm1yYLb3Gy0Njc7fmwK+6o3+vY8rX/xI2npxALI4r126k5ulb
fiygLLX7soegvWsPHUKUyt8Oo6Jxo3fJhaHbjQZ/lZqvO6dlJ4FXG3fMKj8ZMQsI
Ccpcorl9jrn5rIVB1awGW8p0XoftG/LFiBQEvejtnFRKORsUxWOAEmeC0SdW673v
5epMTfSx61MQTTpDzXSXXgmJrzczOkF2BRZCq35IHFS+rMuzpYE6bmwS4hYoVZda
NszC1N+h4Gth8lZAecFYwQJAVel0IDL9WBzlELHCmDZER5P5+6z1r9DFLAwFdJyH
rq7n1l8AhWphSwkl0R8KnUUgz0FTzQE3SMCTZ6hYMb/+ndkWXvVblD90ZHxu50zs
RHj2Psk95xpedUyWD4NeU5eWEb3QGl6wlNMn+a+fZgeJRnN1ORhKQqfXRE4s0dJe
/5Mf3158yFCjW1Fp8KHk3fT668YWLCCfGZkaogOXGgRLSgG8i2CfoeId7rI1SnM7
uYOpCndGkh9ICQ82nrG8NgkHvTZwzju+YyVlBaTYm/V/bKttNfQpYXwnJg02BIna
8JYC5PXw/K4nuzb/qE021kRtBt2yGGueG/raol19vFIrL7MykJiPRUd+nk4k7nzH
RXRm3EE6bqOIXw0yO0nGBNy9gPwKIF4N6ZZ4u9UqslrmDG8Gx5ib+0UgSHjNVjsB
bB75yqsw833QjnyuphLX6ReHBa1idNAQnmrrK/jLTaA9cJdNXym80zvEYYZqWGHe
lDZOEpbqstzrYNBkDAWDZkrtk1tnhnS74IDVZhyrbKLfnbK/oNJl02BY8Ky0vwwL
67ril0MiZRhC1sUz7nBh7EpZMrXQ/tQZG3MbkbS/JGOsJD20apzO4CxvhKHJYAbO
qpJ0zTdlGckZIHbdhXRDzno5+mCxAw2LZHnhrnGWxfa7roKZpXnhmSRBXx2a3U8A
DoblW/+Z3AID/t7X/KtuQwd/WT12j/7BJQQwnbcUJSx+BQKCXOimhBHA3B7IoPI9
IrQdF/QarUghNLToWuYk3nhn2w9JuJldHTvZFqUPGICjJ02RfjE4P127Tma34HO/
7cdg2D809hN0+KSey4xWAQ/H/tl+RwKZ30wr+7XXoKM2KIMvCOPABh8IkTOIqbhD
PqqU2wInKIkIehEMc+iOHLY161KqlxPXnFB2EROb/wDN9odIziUrw1zFPuazQHjZ
Cr9/yg1+G23T/LHc7DxbfyYD4L0oEmM3mEknpvaEbb2MqhQKNo3ww82n+YOkV9Ne
2DmhR6VAdBPZKHPPcQVs8eMVL7ohVGTZaLUlM/Z24ZoGFBlZY3cAwwa983U6CXcJ
iBSAqZa9UcZvimcALGUM0kD9NKhUdRepSo1pLcMTcNjvjJ3LQvognfQGEiKdz5Cu
/zqpN6+21FxZW2hQmfMgpEN26DiwF8OO7u/8jTukq0hVdyxKAxhrlunroMRWK09O
Jzimhby79YBvpKvDJ/9hrp8MeHf/UQMTqcP22ipmoZce3LViJxkOg5rE83b1Z7n7
q0P2wnd1bLMnccOv89g9ifMSpv4GVBAHNvNX6REOYILwhkWC3D2STxENOyMhL47k
Anvr2SLLc5rIBFo7Kk8wYsyrwbq68+ENcS4op6bAIGq2HOGwzrpy0zn7DTImyT7T
kQ9CYd/7Oe8a9bii0zgUObcAJW+gBmr/862Pmnhg47PxRpuormbpiaR9rpjzscU/
VgR0ByThRgs/DbSGWicMHmtGaSvxcWg9Xu56D+dLUNpvQb/Gyd2dgmAO+vubiHkK
6tUIraFuSNX2Eq5bWtzPhvufUB8X3ZDz9LSjBLRRCOL6TZKddidZGH3qiYarnteA
bPiRmg85YcJswvzzMtpR2b3GrTyvnRh/c4+lTZHgPZBXsEKJ3Ilrc8WmZ+hM8Ffb
PmQSs8l9MrstGWfn4T2Pd1aJBi8R28ItzQbOdkO/X7AqRnD7frHKzhtPELE4O6uH
qixcd3Q97fM5SEuqlkppvJZZCnpw9uxOTlmOu9t6FVk7DRLeHWpVp6FxryOEWw0x
BHBWyeMOJOYcmImjVYZFJI8CKqxOuol9LPlUzze7XzumkShm4PENlUrbXoGkEu1S
U1gAA/H+RZu6r/kshcRhIKzfM0uGmSVdLmRwWMC/auQtPEnNVCKWzSmpCRb+R/M/
iVn8HdtMIDq1/QT+BTAJX2mq3jq2FCEqyBQHQ0Tw6TuNZPTRSuFsN3nQ5HHrRAO9
5N9sHvV/nuuBpoLVtroVmp/1Fa+aLu1SC3giXZdn+fL+RpL2isMaSrBRwB7IulNP
v/JENmtjVIVcus5qB337t+WbiKmIb9ncqJy39nkV8u/w3V2Gdl8vn5mXAfo2pbSj
wip6H7o8VCgLyRFVAiBx+/8Fw4hh2gGFc6VzdDuyFgxU4I3Tz7rpuH3kZNa6SH7v
Ogqra6/foLF12NMVc7poTDRFcEVOTdtGq92vFjWHVt0lMtRrUdewMB2ElzqE3/hC
bT1WlBes42/gH2DP77Rk1uGB19Txj/NKFcs3pZT66xW57xu4XBuhuzdZVY2ywvqY
VdTgNPMUpuIGh1k4vD6GsyhPOrCWKRhazEweWaSVUvY+9lPG+2PYfxBHQX1x0A78
hxwK5lr3R7fSvj+0VAtNWOFkRleWabimPHI9ko29raJ3ngqPeaMUp8DzoSZBVloH
LoWAmayMCgJ4QM2EJXmJHuWOlOuElFd/HvRp90yyguKKKVOnwULREofT1ug+Al8j
5y7tzsjoMWTKz4VCvRX+TOBa7HrzAsL3YADWy+ZgUX2SirKlJ93ZSqndMi5pi9vG
/FuGNCK3ndQdZOGBrM6qE+l0bSbKP1Uu5qIMVo4uWuniWDmkUI2FvNCY4vo4KxNM
6WwsCJVL000WOJt3hgJc91Hta544iHqpZE8Lq6PtTQ10x+d/4Wh1DY/98dK3CpEH
glsO468UBt0yD+AItzfUBjfhwommLOF4pcuiKU5ieeUsl79rewMxltV+d9IZo6BA
3nTZKhX4rCIYL3+3GpDuxdkq+1ORIdOVYwFKr/rTKOBEZqikoGy9wHpIVJZSkJch
k5QqqkxnyX9N+yro6A83nQ545TeyQ9pnT1a4rMNNwCm9/H1I4ESxrHzKmf6lZTgl
Lk+tsQk/WLiU/BAVDYNOVgWsAt5yB2Ul2TzwwOfE7a8IuYITJs45yjHLCClQMyl/
O2+sIcCvBFpgmXxOJptu8UhzR5WWldNAQxZsCwY5fmawAXlqkPdgLEZcj8xTiHcB
HZZaMOuhsOpJ8wl1DXSvdA6rbz9vKaVL+YPAUNNiqg108OsG5AYC82na8Mekqvnl
kmYrKNZmPVdSVP2toc9PgEAp24yvdSm2b2BRC0mhAjpyx8ogmrnfFMaiv/RqnliP
ryo2+/udjPhN/LiLdC5eB61ZUtmqZwp+FSEmf2xu7QL+W8Oe1hPA54wzS9O/ziSb
rGkY2+KVNA1rpYm6vva1KG78pN9eyjBXLAkUQxDbnu/i3GwVcNWUriEvPFSTDaA5
DbWvToBUA2AR2rRn/aQ8HRw9dCcmMlCw7Ndv0MxtGDKvucfY/Gy1CSC+YNlNyu33
pjkBiT3dBAeNw9XhyjTACa/SNXZDrWjwlwpwaH87F1fXncbsdjY/2xXxUmngGMxK
CISa6ijuJo+NT7FRM4R9mvSPKjW0Q92i9d0I4BojkNypgAMwJaoRz8K/T+zkeEXP
BgVoKxF+EnB6dJ5tFr8y/zg0DccFeNuh14yuAHMKwliFZjY01RGFiuWEjaDn25JE
5IoJXmaCeSMf3gvYp6c9ZmBVxmmwvzXpr5MHlBDIGaxsvOLgPVcZG+ngiCFKA2wK
h5CabOnsl/OMnblkMR7VFbfKT0TcVJnYZjxgdP4mRVvNYOLZi+8I56X+vmuVsM47
sLQ5jDU0W1jKPU2fFQQl5B9fyoIa3dVJLH1IzgtHJ1CFl8ENLIggfEo132BwprqK
JQb4g2rHFtVPUCBc6qfLINCSecIJuI9t3AICLr/Hk0OFZJK3Df9wkvHQV17qGH/l
Qa75UIqtgGxa7ACIulbuVkHzVNN+8zjBGoGSa1CIC7CD3i/d9r7pTfO47fZ6oDD7
rP0+vmMnPwD2AMvJE/m3cuwpDwexr6fogjr9LJq15MdUbiOWlpEDodhspn7vkmEL
j4/FR+l2befzf/rfzPeizMsSTFJN60yOxvzdbsebr1+QwZxrqQSO4uKJYVkWWEHh
Gh68mu1UhbgIWqkKRx3c37nB57UsGcMeo7Q03edh4BMKZdy/oT7o26YrMsu5sgi/
oFfe3Fx5BLcccy0NNVMsd7Q9Ls9nOLHrbZPJIA4tTTGEBeQz5/Sr97uJms4j7t8s
XGhsgCfzuc7Ia5IFva7Unjpo+xU0dN1iaNfx4vCTLrVqNDCkwA5vip6MRQnXu8hZ
1v8olp9LlKgfuQkZNhksNY4mRI4y8Y3AxSDM73ESpTTWSO/UFEJIQIPUJRltD9gL
HEHVLToBaUd9PN5Yvfzrgn1Sf7RjecBHO8YmxVVWji8I6y60JgGg7Xiz2IzmKS76
7/H5XcO1VjtHuW24yq0XJaMHnESWRsbELeUtDXQ2ZCJ07Hp1HITF0vbxxypgFkLf
0fNmV/L9Rnm6d3zC3OFMQmJr8cUWgZwmrqg7fOx9eYJDHA0nUpnFsZMkt0rhvLTH
bOHCIG+ihkV4ze5smfO2bikbOug+M8ZAlZLIOjbXQ8f/O2N//SBSI3artHPMH3vw
xJ+TznKkD2NaC7R5dOeLnCerCxGZ7j2uOMmhEje1AHYxFBQAeq3TSpzR9A334xAb
g8j8qRd0kMYQTFFUejYNWTP8xQ0QitdwkAp15ChUoZvYSAB98CnCABPc60qqrF2s
+7fky8StseuuY3a1xL+LVCSDvWRbsx/FByyiNlCgrP7AhzSeCcrW2We+Fe2V6tpJ
TkfApNO1Y73XwEzXcDMQsJw8jD6BM1yiAkq5wiJVMuwq+WM3IYZMHrAwI0P6oSjc
Ni9+nCVUS39EyUe6itvZFKo8/JuXM4iDdlsnBvyPSfeiDhDzObfSzMYdHTZ6xg4H
L9XltkBKpOYCxaY2TlbmeFwehJ/aXpzXZXAOLg81C08DjFMiZUiolg03ka1+c5Qv
ytfleSW6jvin5VxHE3QpLbXQ3MzeDyfU4Ftbd3EFUc30KwCdo1pKTWa7dZv3/qeg
GYVYyQ7K9eyuff4KRoeThiSSFg1xSzKrj2oyC/yhO0FP3K9JyNsU6K336BPwt1Nq
UNX+SHypA14SfYMNOvloKUbyugtwIMJ/UlpdN9ZEyeOgdJnqH+fSmCodcWwn8o+a
2bRSSBzivoJd1EA8ZlbgcANmWNLd9LnU5da9sQIqgSzo6RS0/L+BRl/5urSP8Qx1
SP2KVooknjKGvNmCj8scbifNxhLKpqd6a9eQ57D6ZsBkY1CjwQGLn5R05HITkgQ4
3sufXizuvc+YSMrRnjjUTnKoDsa3irW0WexG96PjYfIKvUhjj75fj+6y0tcthpQq
Y4/O+n1SvZFwb2Fe0sptY3Wao6xogZBQKfVjyaus5/Ry/jcMcqMvI5UcxvAuCLFK
alBzAV40iihFWADxF5sv3WRWOHl81XkbKTmHWcnqbl1fZeE6bqSNhkHDk/MgcceD
ezlOg3V2qvS1JvnkbCDGWFbW2T/pSKFn+3E2y8vqNUZr6oCNHMucwtVf3sWag5xe
0KEC9SiaK2ttG+E0fHDXidJQZTBKJDbR1H9tHxe3s+3sjM+B2xMEa2rY3tk5Y033
TnPSIfskUsBZ6/gMNHOKHbfh+mNM+0ZFsXtyDcyouUSFjkhf8ql7i2Mu6QQNE9DE
gAOefnuqrlmX2g+SKXWtqxGY9ZMyfP0YvS/iOGuO8GFiFhZhzXtCA6aeEX7naoWX
9kDHyioIIIelgpzNSVxoYWUCBP5BJwTfAfdcUezyeP5l/CJ4/oLijhQgFq+3Lx5v
EWmdS+4usUC162Rk4s0odpi/3KvQgcD3dtgR+DetOV923mV0v6V/ZhziauaeTryq
0BXC1jfpzHIxoi0dN5LYdVcMu5J2g9fMKRvdmF9124hMOXWvXi458Rq84iFqE8LW
3QGcCSinSxs/KPZ0l0elFWhjjAttveexJ42Nj6ITkq0E6BC1kYYrG+bk9BBZ3jdl
KSihvL+O3cEhyAM1e07TAmx961eTJ58pTjZteEHxqTsGh+gAav0wZQ8UaTPtfXHw
BtEfrV9UfjuIGrSPgaTEuyhaFdo1IpVWkCfuqVTGZfO1glGE2oYooMxeu2m6unVR
TdUd9uSkIhQpr/GVhEFfc99/cP5jIlEBrPUCmG6AAOoH8i9ikO5reo1QJQmHz3vu
1S0mhxG1JCjsXIPYZ5b+BSOzxt4IcHrcIbsByLqvuPW3928XRgvqyR1nFSabl8T6
45MKNnfml/i0mTfY8Dji3fj70Ss0Zt2A6V46d5XTsYYuNr13rjkDgmdFoGJr4njy
89SgaOmU7qn/o2KuPWYyUtsQneQgFoTxLVztB21kiJnGfYvkTeR2hv2gNr9FMAch
MvmzHcUFgg4RD8OSmKk2hOrTnwzFDNM/LBgmzHvkMng2rBpX1iQNO3W8K9BmkN03
NsqXSkvHNinuK6We0ycSKxrnf06qJlHFoqE08zRNuz/LuSZ9RqaXS1Eblsk0FAzD
KmKcWNKaB8YK6wc5/0kbVPC51taSlS2vCC+oIpgWQwU/EtlG2Tmuocsi6kHJKxjs
mdDSV1wTaWkF6Zts49zSEMfSUPDuPAhYxJXj++nrddAaevIOeR7yy5xYC2oo+WuD
7R9aFzySJlw3f3uRjyy3DYNl07je0NpZkAfW2/OIFkMOooGlCC5csznTxgSvw8Fc
cqJV/QKo8+o5a8qTynECUcnRay/kLvsRPgk7d/Mf+chV9lyUfA3Mh+wiYlefJwyA
YUdBDQPbyU65JLfnb8ctZmAvVQ/CUgkp9bP0SpmrlRS4+Ae2C5y07mAczoYpNXBM
+/kP0wUboIliPJhSbzJQ5JUVkh8FL/WGz9FWZoccNxD2QnUJCGhwcob6j0V7a5V2
wILjynP712mevcUy5+Tq0Wzn7KCd4mVsD2lpUNrYh+YX+eQ93MhewMmUSwVotEVL
DvdetbahA8wzUBaN4BGJRlTFgXOmxdgw7ZKWdaO2XK6z82MPBb0W5QRh9/wnERNZ
nF8oReGraAHh/dF9L/48ZvgHWTteTT6aoeZayNjTBG/PVQFPPd723YYX6BNfXb6l
610+KOiGL49TPvgKmCIdeo7JzXLVyzpXKC+GNmhYh/hfoqtqt15AR25QQdOJLUtV
7TyvQKGtGkKTlW6G1Tmfg1nssmMJyfc1SL4QFk6DKyZLF4ZTCzweCRUUrelMPADf
MrdquRkAAykphDE/rajRnGKpJ8zYAQ74/cDfvbZV/AnUgSnPu0+htTer1yAleCH0
jKCTy4Xbk8kTJMeUvuL9GG8v3A9FP3TFJfHZYxSEAFRi920RDrXcanteQ31AufcC
ERsHnkSonw2/gZve9EesJXJpKu37ATvhx3CV+Ci3RFGnCEVPeWaioH5FL+3lb8n9
+s1D/L9LCjF8F5zG+SXstNjAkia//zqOU+069pGk/bboc3dMRKGdNV88rsXo5luM
1Z23/2kCi6GI2kJDCJB+B1aarRmp0jRygVQwqSgqU7BVYBtqWuypaJY36rqij66h
7mbwvJ5IJy55J6It5BFUQ7KUR7+IJ6GS5rF+sG9Rzn7Rud+NktOuyEIt70NvCkrN
bHsUN7hQ3bY/QYMVSmMwecistZ9u8rtm0iK5RKBqfTQjfoWNoyVcPd/kFMNsheLG
Br4n5bj/0MVlsZbgSGDUBOSYDmFt/XvYZQwHcvuojKN7wtAC55ZNSANRpXZkRDIB
eYeaalqKdDt0EWHGcSGbzyXbmMcyL0tgRWLZ7WhZLFW2fTZHC0byTSgW74RnbpSN
z8r61HZpYwoQ8ElLTGV9Dnh3e5wan8EyKgyE97j5gI/eUtnGdfIp1sVlONsbJmL9
GhxO/z9SvF7PKoZ0SizgsGdhn62hsxL7w3MzrgBlgWblFUrQURX6KKKvlCcLkWNx
i3zNQp5IUDreFS982CH9HFQ9gy326DwDILF0dtGHrC8hMHl/DMMholBUI/dGTYC1
f3kJUPiVjoEPrqhrLRgImLwhUdFHXOrxfnemAAus+WPrAy5t8OsOEgHrj9UFlqRW
ImjCellBIXNILX249qqS6u3hufIT9lJ19oAiSPsOFeOf/wHu6yuL3s3Gfpt+f5V0
yXp2sIvsA+m3rfKgUvZR1TFRdgL+66dmRhdHq06uYdfQYPv/hqx01z/8qA94t/Db
8za9AMjqk7o30kwUZP/vSVauyiy3yt6KclWERtZLz1iBWlS2dorvZWzQGVXTpB7l
MurKvn4wBgXYlBF3CzlHs/UsDO8k0DX3CZ9fWVU8mIZ2ZCxXZoRfuVN8jCL/3XWG
jYdpywFT3EvwxgaBBHlZlMnpecKMHGYrCRSPGrOVDQjEBEcrH1LbP4xxVru64WCS
K0qfE8/So9iQzqUcmN3enHufA5Xp4cOgXBDp5BH6eGejL7p+iPjN2h+slXEMvykD
Cqla80zHchvm05rYxhswPiZW6VZP6/hHZ6AnamPayAkpZm2mWptZ6baidzWjxEik
zSxZnEVcZowQXzXK+YRSNgUW1fXVxGkjxsVWa3yU1ySpv7B4ydUYRP1StgU2Atjx
HKcAmOxyVT5LeADgw9EMi+rZFgx2DShMHfnH13vciu7FqRM1SToGuZO03aAyTeEn
Y29bXbu/hj42FZvxMBnydQ6jB4MPz8KKEKtXThKMsM1UG71cN9P9v6AEz/uXIDaO
WjYt9tYT8ROkq+/JJtQjA132WrAQMRNK0pUhZUyzvvWIskb2RwRzmLgkQjq5MdAz
R+Mv8rE5OY8tJDOEcy4drstpaISdzxrdVQ8CSd0sSS23sChZEE5xTISu14lheoIe
OS139uOzeUVFQUYhDmQZljDqE+WeImGTtq8Kj5K7WB3RY/2XJbMnwaTB25RdW641
7DWX1SeCZYJ0TbhiMWL77nqkfqYNShiqgCjVjjgmoe1DFHbPPrSTnp5e1sVaIZfn
K6yrC4xI3c83GuMd+ohR4rp1HUbgC1tSIM1oizrTYQKaTFC8PcU2Ah8tJ1ks0Ubz
VZSG5JY5z7kydJD1DpcKMuMcCx9rC0TF5TOS3xHAoG1kZx3WKqvksAcbf+RBAd01
vPVp1QxkEMhmqZ8zLfH8eNoJ2BtJHcQwnjnIY+UZNzBEnqIoDGeNaiwA/V1nHqHF
EmiGWUJMWFE8Ky9x/5qz4XG7/h8ZVTyOGxY0pGcOo1CP5fxj8tOohzE6hg/F3gWp
7fPG6AXpR7mEPWfYjJ2yWKvo4p2hG5Ni8kDopawv6atX8sREeBT/GT5X1x0DtGG3
Dg6ZQer3vY0udV/mA/IMUwlYSZ377smoYTvwfLTt+PD+siZ31s/+oyURPPbVAnoT
PsKuP8FAFV8P8QOQghatCokTUMV5gpcjLsGqvrvswS0vkDd7Pn7t3RldnPVdQMEj
+FNZCKS8o7bZ7ZW7QJDFT6j7iA4GsZr84t314juzN5T6HDK+5JawNPgjUOPBBOk2
k5ryRH0vqe1DqGR2K+PvucMmpu0d+9/9b0e3fMKrdpT0QrbBfniWbSw6BtIZ+37e
TV0kNq8kfEsSO5yS/1Z/TVoTfsQGzAQEEIhSUhQrFJOZRnQ1iSWRKUzKk6EQ22cE
lxUhukH82d3d08aiBKsL+w7grX8LPdDONarpg7A9r2iiI1IvoN5VRhlW0SjJY5o2
c1TPhxxnrdAe3gWctoDUZgCT0HO6PfT6mLVXAyXC+2MPxxEjmjm2fkzb1qTXIFCJ
+nmmyDkMeX1QnbENaOH9l9ujlfg4DPMAnZiJS8Oblv/q8BnxtIZqmF1dXkhMcekW
oPN73gfrXzHy9uKLLjuB+FZ11O7FzGr/53QsVO3ELiKcUupE9G4t0S2+Oz6D8uET
IEG88s9qf6vCVc0G+lV1+Q1WP1a8k3VYMx/Eg/caPYUxKl67EoAkqMYLSVWLSyVw
8P0TNZ8D0+ZFX9UfF5Qa4Qe4avx64JfBGETRaRWWl/9I9vh6DjFXgl/gGCKnt9wd
XR9EuSNkko4eLm8jPZKGrfZNbS8N1C+uz72DCawGncbChOxrKGyoiwi55r4VV0MO
t70r9NvwYM4mHCmQo8yMee3wMyidMKSVciXRMtJQoZ4en29DNdLIVGTLo1Y0ipxg
sd/c++z2r1TbMcjd772ljf4EXLIwCFTe4WBph5xT2sVKoBEG5Z26Y3+XlXBACLTc
W8kknpZ+Kvbh8I/+Z01dJEhEsI8Hv1bQ3Xv9LflSf0znYimcbAZAeOSF1GIImNyL
qEXYZ0eILk0p2wIlMccl/j7r99tT0VK/iuRy51zQEUm1eZGbvt7yRY44kOlGJPla
WuSXwLjt34KKRQuhrqkCWWqmiSry6C3qhGGFFP9QAYZsI5mKqCUfx1CY+KSr10pm
LLEPzVlWdE5n/qL6qqpYWck8ZoZb6u+LFAINtXjTm6Ah2tiswCtxQROxy51RgLUY
STnkpdyO6UTQsBulb/uqIMIAk+oElij5/rUxf7JVhyNomp/QCInDWIwiuyt0tvGt
u8pktitG2m21m/6WZQDqPTT21MrsngLvovoi15p1qsHx9BIrCDu8kZTURhC/rO+a
WvdmUR2qdASDdsVdpmMtYRTYgsfND7q5dOuzXZkTi8QnrGjYoVM9D1Zsg/YKjWH0
o4y1j8etwcVb7H9Id2b6RYkwcaX906Rp8tf3/T1UCx22IIYg22uY96bpV+zhfAcn
sV1yEroM4vrXskaHXEfa7+Om4a8JpcfeUIREFf+Hp4fkibiLE1lYkWiMRMO6EgDB
jqTTZmFSn4XxEyqYxzAQ0oTtal49aQp5L1rs9k3Akl6/IjWBsj+iYNOdyUB3QgUF
QmM41CmZoUZYM1czeg8sFFhiOY6Lpg5Gg+KnfIhAHXEGlMINwaH7gO4Iujyx4LXC
SVuVX8yn5WsFwVixxiUvVXhrwWEn5EFu7CQfVzrUg+qpDyYii7OiKQFsx4pIpzhY
JHq9p8LPuFT/R6ODSDwH2xp7C0KQaB80C/eWGpWqOZm3dUsKdraSUmdf8ts8LGsK
mix/Peu1A31Da1QOiqkSak9BKyGfpiJiR/eQQFlV8USMHNsJ9YqkEN5PqF6Qg/aN
4ZHEmeAZcQB7fD5809if1TyNkDl4lr6/YkqH+zlNy9OM3LpDTFGot94MD9UETxQO
TO5JYTasqqmTLOqPg13cYYBCmW30OPcMX0k305Uz/APVroH70vt/EPz/PTXf0Gcc
uzRgjrGY8j2+D7DN22J2LUl9VQ6CAOsJ1omO/5m01ic16zbHDsSKvXr48z0M70X/
ShQ9P/EcCSTztK83Hak5HKbgfpuAe4OXKCNqumE3+lmv4kFeRDTeU9uR4BFjKR5c
CmT0fUOZMFLRpZEToZMMoIopHsbc03H/qKvVH6d/JQBtOfB8CeLNEANLnh4CxsEy
Pp4u8D7+LLmDF7wc0apNRkD3Z31U/XtfbCuUX5jk16c6uoZGgav9TJF0Vj4qpI6x
Og5Z7afnm6YFGWR6LfqeGkoiZuowZpAhS/Qb1Hb/G9DCJMZ5hulGF2h6O+K+rwqW
FH1q5+UmB88RRYjeYoXQWvO9mdvwviAiw7znwrflsjr8/rfjZg8QoJjv/9J112fH
oNrVj2hXWM1LZHH1DrwIK18F/+nRNU2m4rlprjd12q1G0/+TYQV16W0jjQ7Vkbg4
64JuCHSpkUQ/ICzQHDaxlbY+YwuKRSYyBP0rtOrY04U2uhkxQEt0SdKYvbSuFnrS
OuBybrBmCowgfXHu7XZ19BcPeIG+J+SFGZsFM3aX6Mg0PEv4U4J6yCPyTNAsd1tS
u8nFC62cLqKiqJLnbs+jpHEcvC92qOpQM+mL0y+Z/xqXXIFTvHC61oqGwR3EQycR
ClmXDIKtTDGqVIeoOJklH4for/Q5BRb3oUY1wdAeiX2ZDXFTRZybxVOCTh2sRtf/
pPeONAWfDuOO79XJeE2m7O5y2biHqxvQxejn7qSxFF5pLgtd7zTBaMexKspjlVIF
bH9WkAa7LPLKbq/DrMCUzZNiN9KnZGQtvJyxEXpVifo/HvFvzXBngE79rYniKtiL
Y+YUhxJVDlp6zO4eiNPr1D6O0GOcK8Na7GCZK1Waw2h/nYMwksoCisyPlGdGh6Aa
G3sFOd48Fm/3QzNL4D29pcK77YNoLu/gGpiO+jeM+rPCmTLhEh0/nZBr+K/FDMD9
8dZUAy1oUGWdZcBEwwdoPyTwsYcPTXdrObmheZK1g6ccN+LxDBL+sEDHhHYSvLWZ
0Yxwyd25rvNz6B1chOBBjRXLUbWD/FvuMc5n00LxEFBxKxev0aigGRc4FBEqzLKy
yccteycJrNtEiF1XCmpzNmBUydYYoeigz+p2J2Zebhgm3EZPGiTbjhcOyZnt/qB6
ocGds4MZ866Qb3KHOBa1zhHEyUrCRgfY6l76el9Nk2+KgQwKaAqj3bxA6JuxEgGp
5o13V9n8yZk2belqHbQi8LtBRUkQhw6mhXtBtPc23xbK5qG+oy4DrXYK16l1x7k8
366aMGw17Ec5L34pjT4q3opjfCmNJ240AwwN3vFJbQSJL5MU2gy+0iMvtAV/5pmJ
PYhE8IShRBXoC6DOHB8SwcgnOvD0VeB1egNxGje/eGOSS2A0/hIrwqt6Gro7R7hH
j90FWYBDvp1hPPi9lZdPHiI9C3om0MIrHBepGtnTjRvgzovLbm5aRw50noxab9RU
jnMEjAOWmFDGMPAoZ0dYJfUBslj2wgGKKWhuq6dmNydBT+n4nzZxL6IojlAgB+3t
gGn+zjkZOPyiqUnvJH603siREXhREfKBXI5O+MqXRVQuHJ9x/BxbBj7bweRKq1MU
YllwTyFVuvW/HitvRwEzqrB5qQi8h9eL8UHF9HzddCb/r3rsSe2JF4iGKn4VLSIe
grc5LrGvTDhpCy0lqtw1ipxDbyZOV5J5l8fRmrv+syV0+jYpqy9UFC2GgyZ7L63J
BmltviWc4bPTuI6k+aCIYLO1kl103kMidCMgE7Qy9YKhnyptZ+fWVonQHgQz0+M8
Mf6IDqGLq4U4uNUKMYUhk6Xl+5EjQN/0HPgESU75Or0rPy4T4F2MWK5eJBGarcnv
zvmH7lkAcFrRe8jN6Hfb4oL7sNLO5P5GvyIH/VujPGr1HjXiKWUVPF+ilT9rvBf6
VPokrZGN9dp9KKduLdTgHbZP8iUZYIokhvadDyp9JRy4Wlbs63GOOq0FyTYYbEe7
b5u69XpwGue+nVBfJ17S4oeO2EHeqbrE8iH3wLFERI1XIyUht6SjZyMnwUABd6KM
AJFsuW7aGx3Vs7/wGuhCHBiTjoAtnDmIW9dIYBEKdXwyosq25UOQ2CobSo8744/N
D3jb4e6Glt02ABAKWlLU6UwjZcVb+BtSsoE6hBXqnh3qPQqFA8oNb1U3SGzIux9M
GaJBmMrpAALUve8dki+vMjDbNtNzmqpKWu80AkIYZhdeftap3Uf+26LKSnzjw+mi
z04ggzVc8OqQcre5Ju6lAIN8VXqUsufNOfnpYXIPM585j+GP0i8wUCiAvQEV0OeA
iNRJ2DkHcHwGg08HjZdWi2l2fbJuYZDPUvvDw2CBk4tAD7LQBIQTtE45Y7wUaKv0
GOXXTb0rkeuJyx5P/DaVePHclDy5dvH2OcQG/Z5xxXx1c8si2US++4IhvDZ/EYPb
hiSBRFdB9MszfUZuDrmFMKaeg2AJCAK41LUuZMqcHgjAiCGqV3P2N/iAnBD020FW
/cIn2sdhIFhH7Mjaj1Gcy3kgFGBoSekLQy5EcI+LJ3mbSOJWluzj4UAVGGUIdxac
GPKoDdmiPl+GyTUtbHpn7zWMSbNtcKLvpvHAjFcnpSJ8j2mDptALk9ZyN6WZduOE
XtcZCnvoO+eGvMm0dOB5HnYt1s55Wmko7wQ/dyr5YNZTOtoNtgMia+hsTdKKINC/
rRHa0aOA2AoLHN5j0kIsxh1ca98Yn6Atyu5GFBB10qBa8p/YbwkOco4YW1UjH6OM
7W5FcZkVBScTCWA3vYHfMYmjO5yyVYWU82E5V9jbemSIAGFvgmtqnvVSaoErnVDI
24xuEhJhElaIGOmAKIqKQcbYxk0x1U7PFop0PVErM2yQ78iCrYb2FHz8WZgG9xIO
1TqZJcATEd9GCk+i/NabWe1Yi6NGbXdPAYAaQra24CtUupfFBnnD4yM8YU8wp5EK
vHRfW8pNSo3BA+9V2ndhAib+S9Nxgtm9L2P5AQOG+Sfo5P43r0bEd9Nxqq2y1S+z
ejzQhSxg0a2zRMo6dYofEFSoq4J0wZgqvqGZNU+1+UtfurtXEwUXzO4zzgjHf71V
RW9dlKc5OrDQtwX0VXO8P+xfeUl0s6ZtAB6xt/ktlNOVocfPPVP/J+n3xTZWiPcl
LxcslN1Gbi0bwiuSqZjUzt4uHCyIXcTiTVLI13HFkBu+dBd+I4NvLfmhxgg/gT+0
IeRocBRg2S9Xy3Qjbbf9UAlWTGLnFcDog5hqYxWDrkBifneGOgkuM0QLWxQIDlAl
aWMuwvG0zJJ5c5clIB7gTZUrxPLwwrKzBGUp5/IiMyVDYqRTBEAS+HvxAr8+idUW
RalWVH+a8t1+pZ2CqrR0fVOeo3nt4ciVvC0Ri2XpcZhgkxBwpZN4ckTaQud2XmPl
1prrEHTHGwZtxt8JatpK9zYVn2UemYJb8Ay2WIIjtXHjsrgfKCMmUnRscBkORVDb
wdSv5RBwPJJ3fEDTUHsBcuO72lj2xmp9chvul1TYqo8nRrkv+imGQdFHzoSvh6lW
UweU9T/Tf1OD3xmP9ch16l8lxlH9EK7Ym+6gMuC0i1Qe8l4KU7WIx2f4uydYo96G
wRWQQipAQbK3Db+clbet+Kx34FqeBxrpZuwAc4WhcVyY+rRclrZGVpM6JaknVHWp
Oa+hsSZUQhhKdXeX3cy4Lr5IdUigVeCOCC/tqocQrq/p89P4ROfkvm5K/ne7DxbR
To8y2E8TNfEqp5ZJKmTRBBE8g9d6C7cC7k9BFIwZE1KRK4q/D9Si2BAf5Vp00RHJ
zgC310cX+hVBPfNjn2j6QC15u/TXCl5NwkM0UmDR0X8saTK5Bk8vY6nRodLY9dlP
d5dMDYW1DWnEoXjZs8QEYIrt5/D9mrEPlWS+5Tzz5FzDZGm9Y6+te8LtPCn5yqjj
+FW7nLM6rVdiEYsWVroXRdgAOposNVnGTgsEIu2SFKHXOmNAa4mMwXPD9DhIxvZZ
dFhTrHR9Nvzxz01O+QmfO7gMgNGhN5OzHdb5iOThIRzXMi1DlyXwI8IQ8kXnp8et
RVCzuJ2qPinAVU7VDQ3/Kq+tpkfejpUOs45/mnzDTzCL/lTKSyxpimPhR397Om7l
1Jenr5vZwrWbWgzA5vVXsCUloIZB+mMUVuWvrxYa6RFf9tMx4q0fN91cECoAKnmq
dCuL5E/kMENBEqvmG+SJVUDV3D2DxtZ/owjpA9IE0Tu9Dl1O/3parVN4IGrYDBa3
bGCaYxx6+oqxu5ev330i92U8wJN9MhL2w5l/grGOmNgAucQXCanOnnojzQUlX/Dl
pW3H5fiCJ4EarcaIPT3PFOYunhR/jvvFcA70NAgroperYPaUCoYwLTueZU4NEVa6
gSgO1fHFRNCZTINzHdjzv/69Y+VSh+vPZtycj3v3X0lbvRMTr6PoOCegx1IwU5Bt
YBkDfSingxqDxaO5U1Hc+nnI/WDcWOddj3i3C5OAr0freXOjfjuM6sTuOaOQSk4t
9bvU0GBS86FWRgDVXCxez6DAmc/jo/0zEYHzLXJQFRn9Mzwodcg/sLuWS6D8gABd
XWVpTKure1e7f+PmsYTqQS23R5uQCYIGAHo3eb6cpdjuYmjjGLt6pqSLoL2rC4Wp
jiCJfysnwQsZTZ4kCh04p3WXmsmN3x0v0bieiJulCrrC+U8SAImqE/mscKzPW+5M
DsK2eWExurbLEo5eQauK7sWi4CiOoce152l4tB+W+pkrEbl+Pt12TNVzgui6itZR
wSJPh3E5254FNhgBGAXjUa2Veyhm+uNZemd6z7SCVOKuMBbP52o3B7KViw0tbJhW
09RF4dJJhoxYHPmx2Qmw2O/THTKpqumMcv3cJ/UTqh6G/8TzOBGcmUzEnHs812N1
sicX5SXIwIPKfyTHeGEw9BJyuASxko53gsX9cVpgz6609Qm7DZg8DcIpCJrjqz84
2bbb2m3ehx+42RC42Hbw6ukMls009EJ5vmnoYWfNwBCWXpdEYsCjgnPtswAleIQ0
5+F4V6ejlLf6Z5X0FSMFASbv0N2XhVu7B4UwKVriTLwmhxcpAjqsTBipYTSYciUQ
uXf2x013IBmypLll6yKiaMAQ7YumamiBy32NTNfMHgJp+6JRzMkvXTrF8W/nvjA9
P8DiPEFmrSWRhMOSvGeyo9B22CB74Ze234pnIdvHya6JlZx9xsCRPnO8fMmdajS2
4QfoZ7YVClqldK224jWAXdiHHmpIKecE2oMFvDTCH5qFqy6Rcgh+ouklNOJtLbI6
HJLJ1yvyAaUDwEc/8bf//CdWdiQlRmaYu0UTDpIESNmZdNoUCNH59HvHFzL+UcC6
PsdpgItz8hd9lUB0FZoZ2socOA7gX+Dtnl6ckw/deA4dKpdW8aJ0LwmzJQ7xvPPG
9d6YqUVIRgw3N1vtB7JGfRiB3zEgZazcTQKWR+Woqdcnt02MKzwgJKzEUHdhQ5Ui
d6u8RZOcGOrIY3xP4T2y5ZCQoaljWuPRji3Ixv4t9j9HLJWtnEh74PVEtrCeKq1h
oP9WpCdabL8XIDKtICQ8bcL6GTXkLtsloQVmF1NYi4gl69GS4i0BLQb3q7kXQPfN
3Vqq9H1d3lr8BQBJHgR/2hwGHRW+CMP0dC+EG9DuY2+REZkctpmpI+QOj5gYh7WJ
AISe5VPH2ZpybG/N2m/lX79ckbwQNab2LbGN+X9SpdKmp/619VubVkUS19A985Z5
nS7u99GGflbPvDcUyCXdMJ/0m2ogOvcpm8UWO8S+TAPFPQOt8+/cvuIuuqyHgaYK
WuQGQEK0mAK19n/4T8vusOyAz8KU+tYhGZYD78RrBt7at1gh1/F0Aoh8Y2thkuwl
qjNdWnAYk6RhZZSMicS37+AOOtEiXvCwGjEgU+PW64SygFUtl+M7XiERv2WYQo6B
OP+GnZ5mQS39lIXXRKOSgx7vD+MnwX3R6Jiy6DXaIkECUg3U2PqeDAWrj6dWCk/H
Dtig2GBAXvhEHGaCu4Wpc32VRnmHsJifcdbeweGNvmvaq4Q5950slSqNnICXM617
t5JfiHbIEzOCO5tPzyT8J6dSjejG2eCWz4AclWSdQcwPG4zgh3dbKG6xl0l0M0RB
/27wFtAh1zP3ksO6RfauneX2ap/TSxRx41htLqk6m00fodNqouNzBKgjjIlgcQMp
spYmshIFrIFttNCH1usyrW4LgG26h5BwR8/DYntL5nZaiikbLUHW4C3P5zmKPSz7
OqgyR7wWoHWRxtvGf/nbNL6kt+zO9u7kfKXWbPvLckr9+8VmXuaevLY0HP9P/dzE
qZdZ7HKK6kZ1bA3IYtwMn+yCHw7QRQmDz4S1ZN4Um0BDn5KAg0s2jj2kT+WpFDdN
6lYcOU7c/3YCtG11q70/t6dzudbsC5bpfqMR6ym8Soi+l7tgOekMkXLvWaqSHEOv
Ozjfy+4fVkzWM/QCbb5yVQhONm1b89wbxvHkJPNV9aEZt4/qUfhPk+DinFLlT2p4
aBUvcZjAh7+pg6hLpOYLGl/3WEIsFOFBLHsrS1k3xw2VmpOQXgNaA5gQayz2ZMMW
wvdFud7nMBq5Gsgxs8jbMY04x1hjlQPah3DYWOWBJHy8ZbWoMLJmopnPz+Bmj3tX
cn5ILruDVG5fWvQ5C6V9yfehhBBn4IKQabMRohrMK/szLw+Bn3L9W8/O8T/yTT0E
V7zd4QF4y8E5AqzEfif4viC6zXjNwYFHbtYh8zbOGSikiR58Lm66SsspbmFOdMv+
ePRw7lK0/yPU1xbnPlQCGeYLKauCq80KGPBI0v1PWxD7UlY6IEi2PHQOvOEJ6oJD
PTPavsC80bOoacxOlpjLeC5e6FFvQvWXCi+ZjPqfTOQlLlwRzDIZgen26L4Wm7vj
TIujDda4Z1wmKDMMoxdyr4dSsFss76cQoKvHUQYnPZUifkeJPkmK3g3X+XYMqQyj
YkI03K8Fqr1nN1sLc8KGwjLwCJXUzHA3E9RqsW2tXpGiRpPlpoUxkhkcjkkzIs+8
nhnUaNPFckFW530wZeY5CgkD4qvoYjEwzhN1hTQQt72F6WPSyDjTZQF8Nu603Ldt
2Ib98O7hMfPlldwkcUskVe1UtFpa/LwuG0a+JE2LHx+XbdehwThz1DknHMyzjJah
FTtd+4GZmcZjCVYNCwA5CukOB1+ew+enEJlUnW/q6T0prz8A7Nv7wfePK9YSE3MM
/LAr5AB7+AgOnDmtFp/bj97AJH8VQDRDR6O1cnm/R/VPldeyTiQIyMrP6SZD53Gd
vHI4OIMSg3fJmD5z7fajXJvk+Ozs86tih62IPpqbT2c4RD4aGTE8If2muqLI8gND
BdIxlz8uvpuaVELscQ8K/ikqhB962uNJyJwn9qaoBx2HoRhMe0bDRPuAGvhXzyXp
GWDrNxBEakBgvtbVY7rZaq5EXo8r3P7aaOLZrMj1enDjYxP9ALNt2ZYJ5P2tA2eZ
8+hsAsWhGJ6HOtTywDt4zWuUuY70B4dvs3e31ORNHCnz6gzeMfr135xxj04JY8yt
SCQhjVNwyFFkbzwg5SkuYwBgqU/6wZjPPqG81w9nWhsNREaJUWvBnHmlJk/MmHVk
YBlfopJH0hU0ShImnSnwVh5EDJ2YAKWfuw5eI12imcOKVXcgzgrgAno097H5zb8+
bhbyONOAjZHghPzvTJD0RXWZ8UtFyRKKKyI/5DD/kDcKKZYfSQ8qSPvKCnWiS1yo
K7PArniEHTwe/1xTy7Hzg83ZZZKgiHmaedDgbbIAniskNa/AfvNBAm+p4wjCHDPa
nTujt8dgmWF/4HzXvyiR1tD6Z3rwv4QebIA2TsHeiQ6Umt9HqDBY9xHP/ird5TYN
Xq/tmsdA9dSDraGzQr0Jx4xvhbCG1JFeMO/eZ+kWOLZQGxJQ9QUI8mXnBhx02H/b
UyDyppeg/jyPRvll3vglwek5MvqCoxz87GmAMEx+rECGd5z6CJHYzc9S/r3hEhat
1W7ULuToE0dKaJ3q5JAVUQIMpMQ1hlrfHawEQKEpQVt1+xb9j6uJsihy0KQJzEAS
NImciMMLoO2IHnK3uPC3TJZeLOfeEjrCO8AXWMfOj3R2n+D1CNSeeIKzwDO/0i47
vimox/Y9IeyJAb6toOkbcfsTAX7FZwzwynzooatlRH+gFoiFrj1yyjJgOYxnAVkH
TEXdUCSBzRvvPGZMNhdo7qb9IJYKyh0PbgyALMnkTnutz29emklWBNQRlRHp+CaQ
R2bPUOyyuqud9D7FzSEWo3XnKgscB/37mJC8/jn/wctDypOonLdaQ6DZJRvF4aXu
kY1dVlhUo18puDba8J/xKenQW9VwG/DD/zWGzUo/MdVaw9dqbD6SYZG6iX47E52R
n4+c/WzYficYEg3n7FYUkYDH2ZyeCnAstrxPb/rv+Zucq4m/ZletweZLH5nNpuf+
EYv1DnLYgSpJjOLWFtSWxGI5ndTpCxW9MUfGlVr99kWDpDd3aRA8RnmbS5kXC5ly
W8FPhYerAWzh3qeYUOamFgORUzeJNNZXQtNjdjd7yGOdb0oRKNLFJlX5k/tTIPkN
MYCL++P0/xRWXVnm5LbNEOzYgTOk72uQ80boarzRr+CxGYfux+onrktj2X3H/FS6
BY+3kD02GSSBhlJNFDl26450FEfYcn/ug15ZXD0yVgVdPxbSx1yH6OAkZaf8gbvg
1AnNvQKVYj8jvgnbZytEeIsU+AY/y86HB4Xng+UhNoCHloZSJyPbQNSmXbGx7sSI
1t757u0WKWTKJQNiVzeS2h+uI5HYT0PuZWU+5vV0FgpGMWwdVRrkP36wv6JSOwo4
3KyIGVwOCcIVjM/yVYv4NyZK51Gyhr+vOVhcFC4xOwOl3FrB/7a1hYwkF2S0gdbw
vRIN+liG97SI+4POPCGqnsdPUnGcmge5NAx9d4sVd3on7H9FWnDFiaDzkAMqSmZ0
YEHeZ04qJ2KiE3skqZhTsSDSo/x0HJ/K7QqCvs4hCyzuFq2J9W13vJgqkcYQfpeV
Gzvd7B668kI6i7q1Ss3cv12BVPwSHLqxJgnJsumlhnhsxjl1LDff2gth5dYeDJb2
pmW2oildVXxEuHSMkpnIlxninWh0JdXuvv9ti1gyTI5AMVP1m/jXQ//6ObzrFGKc
zS7/w4m+XS7p+mqjdPV7Ubjc2AW5OCvhfNPcW4v9UJUBHMKHzbiovP6PMdEIK2Ih
BkGErijgNziyXZyG9eYwQ0MFUy1NJHV2WzDGdoDwN1bbw8GyzqT8C/JsuEHEILvu
4c5ovacJyK4JVqpjPThmWfw0dtkgOY03rfc8pj2kokr7SKJj4VKX6flC9Qea4KYl
sTmU8TbOlsbuOf3ufYwKIZIYDknuhui9LTRP/OjmnYNGM3E/aiMDae9SkAsbaeqK
AKaGVuCtl8fCyOY28kCMfzsJS2UnrKtg68BqnB8MsD5JoKFk8FhW8CMfBMsQldUL
HtIQclH22pxIWMjI65jQok+Dy3J3eJ9TCcBBEnqPgf6SI+S/aUL2ZpnqQrI7SeS6
7RtmFguBopbhWCx2E8aQ2vFxr7rhPUiPk+8PWnDn/TmlLqEWNsWsGVUCAMAN/fF/
qvX/055aYOTndWf3AP5w7AraJ9jBlw0dyNUUx1XL/AyR/MQumYRBOaVOseiO+R4v
eHutE8tJWLLRIfTm05AROjJX6LtYV3Xw9ccjU8KAyTZbYoWylYbzH0QYw8FTr7BY
PEmoC4HhtrizIjsaKNms62Qm5DujQHlJALa0WXtNIS6oW1I3/lUxXOllTexsbzSo
7sL09g9e+8jm8wMsNVDXv7WnU1yxsumtUQFnP4TJ7pXdWRpjxKfmSD2vff27wZOa
dHTyBdr8uuZjVYWH+FHBTJ46kBiNe+zU84hPHje5O3gVigr6hjfcgihYj2Z3qlDR
Od3zkyQOZjjHAPvQ2kCQV+ONb1l+Iuc4Vam/qFc/ba+Px3haQykeYgXjHXKQaSOz
sG1SDZWx59ZdoldyGEPHjIdTgvBxBV/UobIIAnmv1Oo8dC44TLC2llHYyBpt29lr
Wp+miilU+u/I9chGU12BEDWhaVjyCPbR7AA+gUqZv8FDosNAj80vNUs+54q9LZ9H
343B73EG7Nz0hQFeL6e3rjzRHad7tl8pT7hhnjPXlTMIU3sCQLXcHR1k8ofuyfTq
Y5oH1T5XiT8ygatyGhgJKBG7WAi+HWu0KQbiQkJhFrh6dXUfPKBo2KmAPtw+WrXJ
ZNsD6Ta+l0rPwrW6LI1cqEv1xkue34W6oHIAmiKuTkX57tTo3qtXBiwJYCd5ReZr
IO5j9kzNDdyqyATKlTOq1OgCsoLOiPyzStKU+rpFCHJPEWrjxV/dOQ/nZzmWOs0Y
QQLW3uAl24GrgiNZJDYQB9c6cvgLypkWf00hk1NJIzbmNIOYstQ2szjbZKfvfNb+
ez8+xZ26oIAtwSsap6QdRuQ9oN1877IpFS//FjHO/93qx0/u7TSxvpP//DFHrCke
OHz0OdZUda+ov23wg2mNJVq8R30+kN63yk7IDrr93jSlzQfTxPGj+fI6iiC/r/Pw
ZmUPv/AF9bQgc6DLZYLqMJx71eFiX336AwSW6BTt8E8Gc/c+CkPBDDZWDggYHYAV
G3lZV/mfDezExXwNKzVkinBrgsGvTz1FS0/v6KOozD0QfeKfn8gA1uJcv6sJmu+y
3QQ5KWyiQMyOHluCP53o8bXc7FswmXtXefnfsKGDFVbZDZK1yWTSanx8+4hMbERQ
KF50j0N6r6VPdiYjghcxrUbyJzFx9pruHgdcEfvsvYFYu28t2U+31Qa5xUOfaaKk
ZicbbWfEjs17dkmx7F52frfIgnAtx+dlnsefY2WH16Xu05c+L45FjtGbhnmsnxue
M/roiRoNemMDdY5OmKDAkZq9ueepVqD/FHpxojFs1aFIkuXgo72nUD587vesj6jP
YMwGoMd71xaNP51Fotx/vXzoSp51I79WI3SyTU8m9WLnE988R5PDbLqDHJ9wpYem
f54VAxdcw4fG9j18wCXRYDNuXJ8UQs9u51mnqdXhs4X1CNm3it3kvwYjhfIPzYY+
i+EDnPf7QR5UiovVodksxXVoGGwSOesjSChGsZq+IMxobHKqZIQhG/8/fbPGTWIK
diqvPWcUwJR8bEtOfZKkS/0ZJLwdHA2WjtMf+PiM8YRb//sAmQt+VUEFyUxw1KD1
XKkx8UaP2fyH2jxFKOMSj2Do5hv07VKjuXdJ7zHRPe4q2leDbCgZZUKKUKAIuIkQ
WbzdeYm2H9Fz9/i8EDmcqjZrpKSF8JesvAJeFLdvRR89G8dvc8/gGohyps3n4UJy
EEr/ywcKEYeHCKBVr+bRp472rj+zkiWyA/Z0FnU7ogYf7nVQ6RvAP42ZMqe4N0v6
rx+AF33MIkqfapwBmuizvLRoTVGF16AHOTBMfb6ingevEi/ywunz58i3HxOH7Cjv
YzNCxQGWqAJrS5ycxjQ7cUvPwlffXfYAwMqAfKlQnrvh24lJ/B2Yzve/Y7Lb+nST
iVbMAveOTP3l/BDHqKsJwL60Cz94wP4lz35VlYiCDKCl2TZs/xF8VqcyG6RMPY0C
X6HTtuacWlxq+wxVfXdfqVm9fcmDOo9LbhOZFvJTwELBbFvuiDfGCLIsU2JMWv8S
ZK7/mP3xuofpo9ANmUg3PJ4hDkSdF/tINQiPGSMHDKoqfB8PxgJFne8DHqwb1qGG
RjkT6HGjgfFXo5QNhQvOlBjAsxQA9bhjxrCOp1G7IT4AhWVb0rQGqeWDQBMr8iId
UFQWz/3Wr218DVvt1/xZOk7u3Bm2Ff4HPszd5ikea+hi0dtbK9ORBqLsQos2TD8F
zX/0Rf730Va1HDzsCAm/F2Y7kcTUYG9anDAN7tGZfL+goJEStPr6MUQZxcCHAeP3
kfFiwlK42gsCKoka6HfrlHnwquyB6kdQzNAtnGbqnm+dI15UTfljlGLvxMJXgaVV
q1RbpQqs7RtsSjczd49Ri0wcX3nVdMZAc3ZAUnTsUjRddUqj/YyyuwKFlAqkJ5Xe
Jo2dgm7tt2OpGi5pIduPgOpX4ErSj14byXanx6hymNer1FvGMs3X8lENAdabzJhC
A9G+XZCLhupbKWCMNM3bEEO2bbaQh8FFCknHRsVlW8gnaXJ+sB0dl7mCKXfZScwC
iqrow7Q7pX3xdfns5zrGYyH37L9CbmxrRwqLNpO5lTJDHBy4Fjm8ZTJSxp8r9S3n
pD4GA05hl3G3bh+OwZ1xhz1+GKDzsIHCYVrPsfKlTc73R0rN08g+ZfvXR2uIeKKw
hiXt01fGXEjWFE8ssMhlB7mYeoPcvFsm19pnKPHLvkX+jXu3T2ShfzxwQ/iQrozJ
Nj5BFVBmqROr95mF7wjeiUPCC3j2HOF+u16APPgTQZiATQcoRpEQUaniWj0yySi+
rfQqeHSNRg6JBMmD+x7Df9ZOI+Za0hO6UF2QLaiOvpup2BWN1MiNZ/WN1LiyKAlE
iouYTm9MMhPiGqVTC3YG9HwejlcvpHijts3ZGfkdLvjQe/KC2KAF5Qj5FtTbwH+y
CbkRGxKOOAt3DpdL+fj+ZG48Ak9OwE8xZVG0xsoHGkr9JEOcXTIQ5tpAfM04wcst
GB85pTUNXbEjDjKQ0dE0jJg9W6CxXzI9X28w6GeyZTaRtNqMMrI9ucO7wJP/S9u8
lXV+w/r/lGCM7Y3xIVus1/HPM4kXBdQA7Quvfy3FV/ExC8pydePDy9nwWGRAiN3o
bxFskbEcpCuKOFcWTWtfGwlpI0YbguBJ7Q8VR5UegoeRIL/gr78sGXmwkRkQYbzc
p1JICynSnAVegX85odpTP4hdtpgxtPzj4bHjvM4trSeu564FnLGqbpzrfLcC+wwr
KZbTcs+wIRRdLJZF2jbCgUBZz/gcse9VZE1iqJdtFMkJjtcHdFQImg8/Ffqzlur2
HVbCICtodLh7zN1eZKT6aaALuFeX030h8zr1t1S64z1jUhQ3+ea05RmrpbjuW/1b
EKfJ3SVZHZmrtJnhTJngm+nKXKacT0MEJWHeYHWE0tc+Y1xexK151W4eoye9gZwD
wtGi2iHbJiBkrCwmhOSFh5OBnQYw9nT2zYTBKsTxJ6pbZEK0gOKYA5V4/llpD8z2
w4lwqcQsHOrWwq2ZZF2PnO/2hzomQh7BzZ9Jhepi2KlBUetD+HkKPVHMfDN2PqzF
cQmSeWN/m3+4/q+JJsbtNHYYuA9xRU1c9aIi+pVb7PeAgIbJMvsQwnShh1zP8Mxz
m0VICOShRvCcOMj+sGb4dHx1EQKhPwktHQzEqyq8Wzt8g5TI/qxcttvyRy+GZerY
20a4aPa9hG10Y6q0z40TxdF48GVgpgVf/+lwLP6uwmMMm8Ysh45HsnK2b+8quIJc
P6NqojU76MtaDiyT3g5UCzvpNCLW8gvlaeIfvyaQP6ok0Lm1oRYEOimc5diEQpZB
M5WycujE7TSUAarN0yWcGSQStvLrRp9sNg/aEQsKZDAUiaJji/8HDB1UFzuEmr1a
QLwxO7rc+ZCy3exHQU/0kgujwZvay/hLSqM+DdlFznYmArDazTDG45TxWQo/yjqX
PDqbUZlFf0rYBcdcagvIbClEc5IB30ZKJXD6U4pt9VvlHASqXj8rKSmeJLpGU795
r7sRIer1sWe5sIn5ZZuVcZDEewFxl1uBOyFu46p6MTNUXIokLDeC02u2bpX0loK/
igr5OsCadRScD98DEBiA+ALtYqU5OviZfRaHkNkX7HUeJVRJEr2XuuqzPqz/9w7m
gmQdlMF8KXYVj+YVK3RiGb+DcDk0zgKIOMfIUI8qSUAUoeIxPLb3/QmzoilMJ44c
tYAxmKEGWyUmuvaNJR1IwIAYywrY6aR5hnk9AMVg1XMl6K1PkIQTBIl+vDGNjIxd
wXvrJk/wydBglZ35N2YWqh5OOxD7lPN3imcQqYMcMfTcSCnL4dmQ/NcB+y8FsT7Z
bIbMS18MmkX3hI7kAjrsTfE/j8ObeYnyGSfZ4BqKKiqEUltTp6JPquuMJguw5qdk
bTyi9bzHXxxbX+fivVSsKqkyRzyRIdmKMAuNFc4wynEOK6c/TzzNHDAeyv3LyVPS
zGlcQiqyztNjciDcKCfKvSTf9bDMYGRh8WKESA0EqrwNhNMSE3A0FrP1WNVNMArO
un6ZLbwysGpbOUfSMgzfLOtg6G7EQh7EYO2I1m8FfV0tHuaSG5OFPllkqkAOavng
yVo+GrgrKKZ2OxEWQJ8jUmO3QH52bcMuXDCEf6I8jn5nSRBs8UokY/IrdOIC4C5p
v2LSj8GZtb4fpnpkn5Ei4V85wbPiE7p8YK4FHCEulKdBLseOtb3VbViqQMKxWIfy
ExwYlj7ns8DRrkix/fJJ+US+65P/1ohbbkEmzdbhXZci3X7lGjqGXmxaXxE3Hqah
jf7ayttc8m5/LFFZCwtgb1adAYU6tydA3f3DecYUqUp4VwXYdAR+/UtrPI9mb8su
JR3nEUAcj8cG9t1yfE/L0wod3wUGlN6nG8IBVY34nErsEqauOxIXrgkEL9EJHeMs
TrDw0yAVLfz9FNZKc/Z+PSh3I7BNb/pwPVRq8ukZQp8DF5mytbl4N0lMTdQZCqRX
RlVnTVsxkfqYUQXOdJMa3j1PySm9Erl2lJU6vFMbWAFK+0rkYOqo+L9H/WplC9/I
y+pUHtOOtDCneuGr7HbkALUBxwwDMSYxSbIbDm/0gPLcwkbKEt3LAX6mXQtBFivA
aHtMKAlHxuFZy+Y5G7Y+a7yJq/dFnsBpKQIcKeDjRBqiFPdusXAJkm264O0yNoN/
Hzacm0h3QXqWyp3paSYvb6POvKYHPrJZ/tkOPiWVtyRhXsr5aRPCAiGEuryeNr37
UbFbsOsFUVoE0SDmHZYchXS0pi9q3s1QULrvhrBcp3cKj2pBhYRVt2dTX5wRghwb
WHpSiNb8MbNPbLS7TEg+mf5bHqtNWLN2oIsmGkj/LK3gg54cxhrD6f1XConq9jl9
hSskDRx6/kOAfTfyGim27vDvSRwzNBjPODcHNXs3k4UaFVNb70Cx6Bm/AY1SUhl3
657BErGFQrL3Lw6iqXqMxBNXsTsyCoLnWkNDgdngaMiZLaBbxxai93VGW5MYAJwO
v2qI1Vo6mro0IbwWfoengQlU35aMXABQlTkZyaOFhEhAam7e0dQgyjnL20dEI2P+
13K9jWLO/ZxB5uSy0NMMgEVN6wgNuVdG41BmM3OMLblG1EXIBqPMShDpOxM9Y0Uc
lq+8HUmZh2IrZZLDHLIxbxX87DjAXwiKLbvVTxo5LYhIcCeXbcFhO5lAbkrMqnLf
7+HlQo7kefEGNoUBO1M/8nsgcCHWZo/Z6drVAee1VoqBtn1zwyr/CrUuYp+zjqa+
TrfwiouLOlPnvX3aK94JWfS+uaNfHcqKVBtY8Q1r9vikuFdXRskDRSj7ElvXJ7xw
DQx97f6OzDir37TGb6KW+MH17QFLJRxcq2u16LTJAxtDLi8Vu27I1Z3GdALMUymy
ibUuNeWKmfw/fhiug0PrrWhWiU/xLvYyyHEqPtjluiZF7olyUpAYedqR99XuIDXk
hjo59J0D0ozMp4X8TZbudK+Ium/BEj609DYlIJZqf8anTrWVzc09TshWgft73apF
pT360UgP/8oI2Mf0ZqGt663jcuy3YgwBmQkAjqAGzHZyYdlREOU+aZok3pDdmUfJ
Rbt/D1JtN/HFZCSSkyNbTiewcr6QHY5Win1n7kLBmW7mRtRLMYyc9PjKtzfXXv3L
XA8zgwkE8vtxVLkosdxMkkP1bTuQj4zyAAlK+N3HIJn0IwV5p2XNu5t5a9w+86Lb
v1bNLs1iUSrqedPwQKIxb2Ckd6j6VtmZGvwbImIftfP9AUUTB27THhGVhhm0aE91
H1Hi5xuOY1OkBStxPYZGBgcXb3kHDUEmhLPyfCO4PUtzhz69VWNw0F0rQOpMWru7
0hq9d1UeVr/9uCFINnHZIpMWnlp9LFCWL3T/YfdC5duFFaMs4WFN6X0H+oFNnjqF
f7RJWx/rWd3ydZ7ywUfU6p1pvwXNHBDN3rocJWC1KYa3WaYCYQLzfXj/aqGCr6lk
E8hq4foRri21xd7dyCPmuTuo+Aey7zAdcaFQHzyp/skAsDwGm25clU6m2YftBr5F
19OXduleMaU2fJGaa16ufOYqKfc9wAgwGNj1bH5eWUTPqd4Hvd8SJdbpDnPD0YZa
qDsBIJJBKLi2r2X/ytCzICtPSrB/sbvz3Ho3NASdvCRuhysg0P0624lE9jzXfwQu
CmRwU97qH/e2sBLapdnp3K8dr7l8iyeEg2XWcwauY9oB3aHt2h6OFrBVlF+QqW2X
3esLjzAK/x4sWQepHjo+O3l4cIdSpZo1OR45i5YPo3sgMoCvvkqQ/Z8LJ84bHUWv
YRph6FLiyMZylZn+Ltm7Z3zIRdOPxktdj1jtEw/86Cv4Nbp8pXbeWG+XOQx14gpZ
h9KlnarXGeYCkomPXdxdbfMEACLafMhAarM7/5b0D0kZaaRm52BzxGxwsyJplyBG
zibZn692KmfbfS17SkhHxgMXVXf2QgYlMhbpSAHLkx5TyQqF9gGdQZ6aLUjKoAqp
L3ttW6DcyUExtRjydCGn96UQuI5acOgQmKeju+w9SNo0ynbRzSiYuuhVKbXGjahn
pXGpLcrCTSGe39IerI4qi3s7HlqTtmfz0+Dyy/rlEppy50u0/Oa7a0sbCaMdrgpU
Q1kMYWDtTHK0Y7qj1+uPenN79snquLx6qBhj0I/7n8OGQMD0Uuobb9csJ9NISRLX
CDAVhQw30NqdlFZqXTu7ZABr04rOz8G6fZQb5FdK46WQEepQSaIo5DlCGsv4Rm5b
cTqIOmY9CtJOKxZorcvsVW51KZ6bSt/rh/TpQflUt9hR0CEQOxAQREN0WO0Vp34E
IQW6JKdAJc5gehicFUNbTMgyfu825dTXLvadqbvONBljk/evx17/PRD2WJoRWLCS
K0ydCaP0Q14DT7PJkdZ11EtZXyzvb22JJyyLG4VVA25MDAm923W3v4o6SCYUH09m
J1jIWYNhvVwdDfVPk+2QjtSTZHWnPaY9JTubQGL/0ldKwWaviXRLDwalke22nwGH
Ob2cBfx99mKG5OQZaLw7xIVgAJKueqiNOikU/USlIuAoGd5VKJ9CzilkYJmdc0Qc
pqtwfgT0w0Pp7Bc3lyqiuXZalM5wQ6a6naYrIQjHSUoAewomQQVhvg3UMQLINABX
xpLCyvCJa5l1T9ICcfWv0EROL0WP/RVkCX/m75zX9eMeFJZffGd6v5zAG07L2IQl
oC32Hl/jJzrT26sGDPRGzRSBqJcoq3/QdUY/Xpmixyjn2rGkZMxKIJFpOhIyZoLE
92CwQJHBK7Zov8jvyhqKmDM/yYXP5dLeF2yQVZz1BSBoA3bxVYyT/KAftJTaA/0J
8rD+W3nkAFknRhEdysvNEjRdkgUoNW79gUXVThbLo092quERm5A3FIFz0XtelpeQ
dlLOzOEveLErOk0enY2fQTTwo2VDSajVA02D2NaF0mtXxB9f+baIvEYK2zetgwE0
0OQVOJswjNtB/Aw/DjWU6flUSQd8xvZRgw2OZOhbOyFQFmMgPczhZZaq/g26Xn/O
rPIPoqZCg7YVL9P2+n90xe3Nb1r26BRYn1rDY1lMK0Ie7w/LTuC/lFoJSWKotZEi
ZhtlBUTKxGYpGgXiImcAtdkFft5MfWSXoFN3Y3sq2d5L0cLlwN4SMfjuEVY2bkfi
DgkADnGbkp+LxlPF42cK6xBfrZiRYia0f5YRJ+dsT37+3KJIkBOQvo+7G2eeRrw/
DMnpfjdkkosVVpp+2t1FCuOUOhKqok62yhau1xKA1IrmYANCCZ+9mzlZe4vDuYC6
S24NoQ6AkOH1jnWjnO48UhzQBbB94fXozs81hNyDlNAmZunZD3l5IaGIgk5FS7j5
6ynmfdgjDqfvw0zkx2hcpo4ZzzBCO0uFlw3MQha/WtSQIcpR4uKDkc56vpEcjdmI
hOOB7LDKNl9sRdc2WauzKVv9XZZ+g7S4LaMeY7UhCRZg+l8FlpRKwmn+xYDf8Vma
V370kQrgxTICzuJtAqILrAaMFYGeHRvP+ZvwCHlkOf35jcpuUy/UYk50sMQGeBSg
vYjICp7niBTt4cOo41oOctuhzZZ6HGsARH4cpl9pn+gTBuPZ82Si/gNuzGs0OXr1
hIA26gcnQG4hOAYBvL6PaI1lEMYh4hL2DPP/stWi44cOJrO6O0bKr99HbastZzx1
CoixH9XwbDZG4Gy6SL2faAyEcs7H/bLLIn/TqjRxXUni+ctIj7QvyVYsV1NckITh
QmMJy0DrEzj7qjuFt34qMM9NRZuHGoNtt4Qx7ndq30bHtIDU/bTShUwoF4rkUlZS
htrR945vC9IvPfJrsGQDLyPN24n5pw748qHzMcs2dkru98kWnKwZtkKGdlG1sMg0
s6ZTLSMkz9T23nGFMIv1mnQ/64PhEalI5nGRbZ54Btc6ZLkvS1epUxRGAsdHyl79
ZbK1bUyoQDOM9+8iRVAiMWStb6rFJjpk/6Z6CGYraaJtC/oOIt6IdgMRVQV/FFmM
3i5R6h7qt9z72Jjq9wbPFTV7JDKgwGbQrlaN7vWGClksmh+NkbobJX/fB3Y8BkoT
x4aBZhKrVZCJOH4UmcgacLLOl3a8Nj8SZTZowIe0uMKFPhAk6VHlIqxxln1PB5GQ
Oig9J8APUIt0/x6Nmn841YI2WOCeO5DU5S1PEjcDWzgOatdjWhQdIj32WysLmkf/
IJO2dJKZBWkoTl8vcnTFn7oSLM+iEf2+2L77FXQiTkCeR4mxjd8rqGpFe/rhW8s2
qszSmtoTbPREA0a9iAT84jkfJnAfCvTs6hSh80qZeU/8Q0fT/lry6EY3C1jtgVsw
rTfofi/JVa0BL1JMAYxlHDvoF6RSRQOLOMFu5zjBFw2U1wjv3pHLYVMb52A0pGNf
2/zLg66HXhHX5VVUMifk6u+d8m9cN+ZVXJFTRB17M7zn0TO0HLRMOcRhkUFSud7k
1ymMWL21eUi6A/LophXxhvO8cqYmkApSH0HPkQ7cv7JDpe1+Psy2KH+cPsocY9dr
ZKWCwOD228Hh54FdQ5V4qXqv4zHiQY0AyLvZpmeEpX3yP7GwFCLnNJMyOyM6GKPO
04OWUpzoZiULohIskZA+8LoBDdsTWLMsccAv8qhtUIFUfIG45VTIfmJRMyK0mBSg
HhRdEP62nI1Gof8IypOToLBvbdck0PG0YGssrBabmk3raE1m0q4UBqBXgWvYJotd
f7GNGTGYE5KnHck9VoVxLtzZjOqOQvuEmdt7DdMGx46j97eRdCG3bIwuIdlnHXFN
JQEG6UvD10ErP50vQSmGV8RIQKOlfgXaw2GXLuhji4G03iAsTDEsNiu7stgWQb4l
cCA2x98w8gNJtSB9CIwV+UR4v1T4iHF8TS69cMCzqIVTNJBwwdNDluoP9wQSgFdZ
/5zr1wf1eAsAXb/xRuy/7VPoVqoXdHRoL7dISKN6yAQkX2wFgr+7iKoxWheiAw3Q
9jyWkZPKsfRZoPnGGd5lYR1TeNpDf6VNFcpB4nS79IVCHjHvmcrKPHu1PJ9qwTdN
QwhZl8RXZcIaktMNx0mBuqfbZEE4AjM9MEO2JSeQ/R7hUjo0ardLA4zclwLlhzIz
u/EmTLAagvnezLKaQVVHh0KeNeHB/v9pkhMx1ZbIVs+CIsK2/AnSWPO5FqdOHQRA
ujJ4045LQVYNtVM0wqYmevsmJBD5syXJ4q05C2vZhW26kx3IanLEUwxThKvaBCLc
56w/RYuq8B+nmbiXGKTbcNgG43YqXwSCOsFhfKWZYJCAm309kyv5T3IzRoFKWXte
uYrhIZs1O66sdYoj6BVX31bIbEzorqhvC2YrO+iDROg4e5Mw4nayHopilYwCPirs
RQwfXiGH5c8fgZPG05OlMTYgG30VLrTgaEQnkoRJBi5zEoiF49GOuMJ+aay0L87R
5QQO+30Qq0KAQQEVtlMI5sPxwf4ywi78TyW4VfH8b7Izr+4Y2a3kJWHPgHwkW1Rk
4FPtKsYDR7HTjoc77FNvujtvZqH3/SX6I5qytdQJjdyjnhXahHTITonMB2drF/Kt
hssHFmCtlMEcH1vyQQFGbCvrqf9hz+bdHGajtsvO9GZ7QUVukC8nhiVcs/HVsAhe
ydlVm5qB9mxG3e+E+9s6aH1p9PNmXB2o9MJA0DsbQV+UD0oab9fv2tn2qWKNMld/
tYbqHpxEaPohBXmUnoRPdjgAHvy8/vNELKy051uaMQRtsOkr/IlCuSzwZCd3pubV
9mOgi+GFDVunrATEfFVsEuOvb8KXcnDM+5F56hVpyUj/bZklNHY2rZiZlAxLc98l
F3b8lSKno1680hqNp4Cl2DjYvyU5n64ma8pPYrCZ62Zqyfe98N5/ID94e4WYPCFQ
0l+fNO2s78naywtS94BJ27OghCn4G9wXk/KITp8D/gYFlPJNGABNdrCdgiyLzOrs
AvufaIOHebNy3vaP+8Cbiev7Hzk8NMt/gplhusaqA0O67DtmyVbfN6Qm+MchdTQk
urw7iLVrq5sVTPF/Wgqa5Kl9bvYQPJHyjuw+DoZM0NT8HQW3PVINfmNdgVSC3/dJ
Jk9u3OknVidozK0DEAqaVIML84K16gBtaAlH7t2GAYGNTi+9bHNTvAm6AHzpJiAz
PxcbtMFOWERj7EyeZ59EpYmTiEotKniKn910OH636BSw5RebTAevYHBceSBsE5u3
IRm0Ww7hKt/RY+oWKmkirxKfroytiARO+rq2cUC+UTaicsmB/m332SSO7Y26mCwO
wJOfen9SVKKKL2WAVj5LESm5BP4Z+z4CAkl4iEDSnEHdvO1Q6Sr6Cq/vs20K68Yb
QgsB4uYOK8DKKjjBkg/HKzgHs3dQLlwOsfa4FgiqfhQKaKrUNSgXPPr+hTynmzVx
on/4DfCmN39oXDQQj1UqxKFzLkvNXgUNIKWB2T9RA0+X5CldqUXcZOXeQS7k9qH/
w28fwyXADU2nbeEOjCwls71FNMuenp1kqx0nytyoI2NoRtgGiM0SKPlj4LIRgrax
Ms1ffy1UvuZ6toXsj4tYn1mXDrcqpnJbjZQ9uuyx+WzVGTqR3pCYPiyq2+wwgQuv
DFCd2/i6XfIty6DMoRpNJ3UgfesQnJxkQDnHrifR67A9w66MIcx+gY6aH6z2IcpC
RIdUTwc/i992MFa1CwsMqc/JgUBfDNOELtoQMXnJOPsQQsBbUEAVsyqHOiZXP5ev
l4QGYmQMKsL81MdIdJ0iMirqnXiyw/1FfPAFMJbiuV3LPkrEb5Sp0ihAILA2a335
MSJHkHJrelbnE3UFHQxUs4nlK1EuwoNK+qhlD+qHZlxSihjEtQfWr9LVB9tbzp6J
P5GUz85QJO181S0Z/xbUzTLcHjryICRvZQVI1w9bmcTLtu/AeziCW6Guq2eE8VOP
DV/rXiAjx2BsHjrxgxiwQ0vcIlbINapBAT87r2PU+hVT7bFb/hiM2FHEITa8Do3U
9osMjhn3WpWpmQ07XTmUtXMYZQ7X4mNJgTMed0vFokELa/TqJHVBGSfyK9H+m6bj
dtQMFF77YoQT40lMhi8YDRucjscaVUiCPMQqzuy+QNboRWbuECCGa1EN7u46LcOw
dBg7eBiknqeJEQ0eOdoG6P9YvQ6Hy6b2y9q8WX0WdPGR/iFbEcQk67nhq+rAQP/K
awiyYJuy+LxR3GLbB+6y45tEWVjEukqjjsQrOVgFHwkTwi0r2iNmBvcu0nUyUsJY
Cpg4Ao8MRq6cUJxAvaYxQl9tfhkdPxEoja1j9bf46cchM/FZo/TTjeGYkkPRgS1S
BvNScf2EacNDhL1P1T5Hfbn0TrylLVozyk4uSneNSEBMF8axjIKiwLI0FKjI6ile
qCZx75Oad5Sjpyv+hBMwbxO20eRH9xc1xeauyzyL/FJz8wIAn01QO4umM1lWEprE
lS1Fd7n4L1QyrcFSKIYeD4rcVPZcrK0slW7m83SW0027xmCe5Ut//6J54A/c5FYN
0jba6cSnNi5j305x251QyuVl0wUj7MoXf5yz/wuujqPU0hdae7Kd8xtXBvr8zxIt
7FomTFsv8ilCQCPRGlzFTfYqclRJZx3eyvhAiaqUuQjL8Cey0qgMg2UXMBFuasTy
WgoLNP9CLxWhD6/1BdvlnUX8YL3+FCqv8hCi0WiwmKSS/S94ymeplrqqoIFsTT+D
wXYqg8pgjZBKbMO5ckZhq9lCuQmzVFD4ujF+jRHkhKR2NcQY7SbIVzT7W5ofFbiz
AOS6rTOAM1wfrPkek1e7dDJfy1ORhsYKjmW6A5+VeMT0u3hSAR/gS4jkGZRflJG2
zCZv9s0NqtLjSFwmKXNE4d8jvt12XmLdnqlWIL26Ycr7KFFjPjYdeN+rUUvaQbIB
JPZD3omm9txfsshaJGhqHc+j/WhPdTy83sJpS5vHcdX8SDlDmkIWoUJCWTkzjyKI
hXTrhAogHEqvaiNuVH3Ggnop/WsdsTXmNxVc/CnZTW64fEOzf+KTSkrynzeXF7/8
o+Whi89sDGjwB6JymQBziVUCoskTOE/siP883DrLdWtYwDEGG4p9JchAZxhUpljk
JsucskGnrQA9fzpt8gQHAprrIXgP5Fgjv5KM5IZWtgaWLk06s7Clks+JcYouGHc9
g/43Ry6ruLq+xu/sfC8iIr7EwlJ7NKsSUnmZVXW8jeCJU1qoHeNBGxGHaDNlB6rZ
Zrp0NmEP8AJSRQ5oasRoCytf/iITAj+xIXHHReBNoFdpRGqVnHtN9lmNciZVxiKd
Ys7je1Dt2eUgUdPO55Mdpceo/y27OdjQvm1j2zNcjCZpG3G3ImPIcMHkLWU5NVsg
V1xD2SnuetcZSG2M/FqQK7kK6+hi33lC524vRjAJBrlrqCPNUL76AXfwoNoyt+52
TPjaM7u3EtDUJOVE2C/tqnamVGOd13JUMIGrbhR8qRxHwlxlsW8ZoBGP0RCGtYHF
pOn3QFJ9nFS0DB/NycONwSW9ZG4s2bGpPf1KFtOPvLQlS4vriuGmN9bGdlz6i+CE
O/6+ZwIZZDX9JhPPLNAKLjuy2B+VkltsCPBeKNkKiYihtEvUI31SBr62Oumrz02I
NBajuqvDcjRMMxTGxY1y/4NFC5Dhc8U/suFaDfzgE5g4psE3LUc3mNdpvD0b91Rj
iLmrUHN2Y2N1U6ODinOgu7n0xx7bZCS9TY5lCtLXrlMhJbI1NHvHy1D2vAWLql5e
cfx7std5CEXehtgXARWxydWM7evp1a7J0LaK2UjADXHzPzKUIoHmAz1W0NsfLiIO
vd0DwymO7ykOMDKGVRPTVrCG2Aw4i5gvObF6hFyG1MEJCGT1OW26RrlKGuZyDkCf
xC78lrvY0HZrfwxQ3coh/uuRKsPcJFNQli6pa64zb3j1fdKXqV+tTj0MdprHXwOJ
lNLE7CivriECbPBMIF4EeL8QhhmYsJN8XQ0QFJVGDFduBChYqGOYzG2yvaAR70cJ
lh2wQQ+GIf13SFXkHqzc/Udwtsq4YPcVcvetCAjVngp7u95plJZJmwsUUDSZkymg
oEABLD8DAbZ7uGkpUt9gSP73VmRwsRgZ+ZjRDel56bu6dAFZTJy/cXybIfwUtJb2
B40YhoYYISYfoyixJwPwZNa7sX5j6c+7Ic7umpz61p6qo3nP8592xhEmIt7eYMPU
jx3FT+2P767pxUWk0l3rsnidxNjp/QSYszeRP4UFlteXDxDkwnoRxklOwTEc+S2E
TJLu1NcuAaCf5R2nrzTdYY2Wuepvlib/V1lxLnOk4xHGHMZjS/ZP5Ncs4088rESA
CLoWbVqXf5TPOdYStZKkjvWV3+7xAIJGB3+XP638fSJ6sa+aCjf+shafYLI9PhE8
sdr3L5elZB+OthU8tQPKcuya5Gm5+lcTGgLdfjuhTAteeK33/QCTv1ZLbeWnu2NZ
w6x4rjVxFJdQQN802eNZaacbMt4TkyAN872dWheXnYqp9HF4FivQZ6lNxDHtyKQN
LrOIEpVWLv8e6LZEcDbbcyZj5+j29U+9pkppWl6WGUAWZmbeNmPvmHGP8P1iIOlf
g1dxYv3JM4jSbovCYx0AMc9qQX9hoKbYVaQAJG3Wt9JJdY5jpXCDuTBbHt0/wVNi
F8bkwHpk8bfRV7Ierd1riNAEuBBEbhQFaubEY+rcywwmqT98JiH76idkW3q3TSjm
00y8TUsGneWQRBKjXetNQbi7+NqCzEiLAtQNJ4EEPJWlEMytmX4583dfl7D5UxKe
QpobnsakIxjePUUfY4aGRICqhqx9laKDtf0pZZCuTdQcSM21rTu2SlaVKHwpSZhZ
nsw+idBtWP7OEJMKvjHTA4y31LcKCzbJttqIARhsws9Pc+f4TWttsSdyQOHFT80a
RNhvc/ReJeaY8ydMLe92Me3f9gcYN8sbPg0/VJ+j4ddHgAWF09NmrWTNFDNSJI1h
hHIRExa8sw761Hm6CzWNBTs8pNJDaB1lzRmhUeE6nWfKLlxGD/Mn0rJf0HoMK/Np
x+/ba+8k8aEH24cIhbYH8Jw0bCLiKGjVrWnCJtcfrl9bITHwuvX23eZnR4QmJK35
KcBg3GT9XMN9xJ6Lzh9hDExqTyJcGQTT8SgGQhwQgyZGcSowe3GlCIVLHtMixDmr
QA1wnX01+3geVf1E5/BFkxRX2/jQs8SYndKWTnL1ebh15s0We/H9F1RTxkdoWlcb
/rLS510eX2R7UxK2IUqUv+tzy2WfYhaKbG7dkLXKIauzcwz73W4eCrixhQVv08l1
AtKcZzAHCxfoK5GNenxtXQzi1YSXivURvk4mkyihWfYXvoqhwNbUy0F6BBSkTJye
LPFWAMiyHfBC3argzjkE8JWaBojaco/cNJ4VqrQlJSYmXOEWUCguTtN5VBAj93gh
8tkYHk3cBjuv/5bi2TvSWK7T6XQyjZLtJVcXm2pZgThKugvKuaFf46fOf1E0fJM3
0f3TxnfM5KRoY6dHMjEryqdgDMgwgkKbZXlJfdMdXWP+BnEzwF+IpU2iK2CepGFv
IVcRrvUlHyi4C3+ZzjO3a4DZHwDJpFtpSs8m0areOSwiml+bbGLwNylkOva+3P8w
tDQxMPISL5M6i14uLPdXnRsXI5s2buI/4OvB1mXVbsSDEhvu6APZqIXApSGGeZfj
DOl+TiyKNy7W2Z2IsS0BggvmQEoDxiEde3Z+OslmaFFrVA21w7vqtuwX6H9niR+d
dyCFzl9VSkr4MbACBwLNcg2oem1huZoqruWpbF1WhT1KuzaAQCa1yeoA9wtfFxwk
r4y5/JOXxVdr5w8z+Uobps6NZEArWrjbKnFH/CzJmFtlPIbnY976RtqkamlSlkJu
xl4AEmRtOELwNFmzk6e7Bd8z5sO1gSlzsB3o2qaRVCxa8ZriFNRK5099JA/13Qhs
tpm6KQY7T1xV15IcbGYdJOeDtIvZ7lwmF1iTGQzr8KidSvpcniXLqR1dtR1uAgi6
95SEEc3unMgJqlGrDK4yJ60ZmEMk9iR3InivdCgjj5XlMo3pLznsi5+QgF/YsmkM
fiWkb2TOKGvb8LwyiduN+kZjXi1vLOdufgObEfpKQqcA6CTROwpqBzp0tfV/Pp9/
1aM+gymE9ocwD14ZXgKX5GibFKOSgcXZ9R+NXU+se1RANeU6IlUt1YdBJA/yZ2dY
EiLKAHeiZTW9Zuyiw0NenWBzTPC9bQh4dT8/etTl9UhYxjxPFupIYJeyXhUQzoj9
uJqPrDvFq59XqdmkLDc2nbCTi606y71SAxlPs0WQUox7QAoe9Hp1BKDvPlsG22Cl
DopSsdX3fbUavUj57//frtY2yu63RFTrRwaZF07SvR4gy8LF3ymoCVxvjB6Nf3Am
6xDXJhDkE11b9Mesx0sammHu0pgDPGEYzFJuuJ06j/umNSMk38kybS3pGldskG4o
wf91cI0EYlCDBNlKFlTES+7zAQSDJKAn+RIkhdPkEhJjEPlEnlrrmWP5I7JXoITs
+OSVRKdiwXu8iM4lTKmAxeLu3kbOKESJroh32vcL+68Zf/+ZPfpDCDqrVnCEU5P5
mwyfEbtR0OotnTn4zuD1BeGzMg66cdcZ/2lC72pT2iR7ebu2Mz2S6uCEKOXGMGO5
l+/xICt9kEJWfxKlo4vfLqO7YY0r1qz3IT8MJAPjwO9O/24GqyShARxue4ORoZSB
dXeAC/CWab0dSwymkbE8lXNX0JtlhLMPdTG9PCTS+O6QwBplAPWHY+NQfw8MOGHU
YYu0smAYN2UIYEVkj1xPhn5TOJeVILkwmF2+OV6Py5jvUjBNEYddX92I8wqsCAN2
wAX8SyGkz24r2KEVYosWj3AwTFcOjHOawOKPMAQ4I6tIhbDU5SgoIGT6S2b5QvN2
fsSm/GlkE3lDeNpEqlU12iaMmEYimyp5nh3eH37AyTutkk2bnSvQ5MSzT4IAjAXk
BSIHtWLADmO67jso0WVGIAaOWvJ5DO4RuNUhcanPoTpQkQUMDAj2p1bUVeq47LJR
ctH+kL3VDyT8XDpSHofz/78j7FY3dEDwuT+c669n5pYBhCoI7kf9pfl2iSH69DRx
y6HC6GZIX+QFtWO0NMbyU7Hag2yCTN0RknNsEV+ci0giNQlVvi+1QJ7SGg533Xs3
6Z5y8I8euc74NgD73tNWu43/towVGf/8kIqvzbRgGvLZ2kAkY7JD1PsZRFObNcLY
OWN1irB0NQrjoEODeNSELY1VEvrrPdlBL3Vs1Zeytf0T0Vl/OQ3YymUfJ3qagTYG
yjkdo7kOmwdSO8Re+Eq4aCjIw9P6pY74Wdpes1Bn0oaglLQQsbp1GfUSlh5evG9b
tlXWNxLuKRYA64qxlCPMVKilks69Ddh3ZP/M22wPpmePNLc8Frejj96WckfP7SVJ
yLKC+5O/jnJVQK+GPo4o7ulagf/uAzA3qgb/xq7rlZjjo1/2Q7GxbxZGnK41naiu
qQBbBdSlijCFChUQGmzjj1kM1ma/hVjFMCCHwIeJkddfh2ImmJm0c0Fo9Zmtk5MP
6jmoi2gta4y7TQa+5sYslYBVB5KaDrp0BMl36O19cf0D5Phf1esidEFv2vYgSxSC
PT6ZnmRLQAbw7h35dMZ5q/oyj4s+9csHQgc4m9jAHbi4LkEFGY20efg0MBVocz8/
UknJiiMLpqJJRHKvGsnz5cLZrvvki3bBpogIyp3XEEMm8oLtItYInZdJnk0NcXD1
MdgK8gGVGT+dx8qStlRQGTBsGJ79hKVoLtYJy09C0A/KQnZn2osny/Kkz+47fn0/
nhWeSYJdHJGLrVTNtf/yQx0cBEc7LS5Jd6ZtiiVrb5ElKw3DU9AqXK6ADd4NSiTk
i7wjK6YD8RDKTvJq3gHrxlRoQ8tGyUumiJLGMJOteENt8yQxhapBa82QI/MafG5p
MtMH5Dq1bICvD42YilliOAQMsCDkZoIb5z8zRiV3pheGKe4DhFRIuHXABA4QLRHT
al8eCtXQE73RComNV3/u7nY409O468KxUL9muNQ9DhAeN0xmJnfv9BGHcKZSgwXe
Bvol8iTH6MohKpBzWSx0Vc1aNVUIs/ZvJSlZhzSsMpws5iyA+dtmzR1sBMbfFyJY
12r9QyfwTnkjEqN5xgvvhNtgciO1S7h6GOXCwAyIMD9LObUmMyoGRd+kofNGRmi3
g/nQsPsPIzjHQK00wj/Pa40w2MCL+g1oilf49LzMOok2nrDA6Bgv5FoBmR+ZSolH
Gpgvjr7G6jpEwL+SIB2hySaIdxjWNOegU+dz1FfnaofVOC5Yrp2vgdDzsIIiCQCy
KDKX07yw9fC0z+MC3xF0/MLCpgaA+rXaO/8gOku4p1hxXjY17k+OAV3WEqZK02EB
BCO720RjJHdgJ3hOnQIew6rR7mf/sRR98GHLgWXOvChAKRaD83c4T73KizfT0SSV
j+WSJuR+IZKDe31YVfCFdylOt+LqLyOP33Ek/Jhnm6rSnvjb/DBW0HK7C9gxAACj
h2WdCW67Sk+S9xkPR4ZB5N3QL8Jx8yDS+lp8/M1PHN7dmoMb4Oj36INjDm2xnhiU
pmiegULfUpUehteKL6zFWKsi5HosahQr6t23uqviaKSjPY/c51q5BHIMGclMibyo
5DOIL3ONh/Nn0q5Rijxj38+wJnMQzmcbVBPPMbs0sjeuprMOvU0QaWTrBLJVXYYC
x8HJnOCJOcgRVDEU1ghgL0zw18R0Gf2FfLM3/lGcNZb5vC4S3xMtZqrjB+YqzZvW
zE+JAO4qZP+D8Al+km0yhj477ryLFKFZcqM4eZXwrdM6i9XDQJRFC6j1u+D0RpKw
1bGA4q9+ffrSqKJJK/nuiADNOl/IoVHRy8g5gctq/Ah6qtUGH4W/DOAunDK7dT5e
aBqpCdD0W3eXOOa0ZlGx+a5eCtxebK8nL/o3twbBlxasxyeBHlzF3GqnjMPwtIhP
UgfzYTrbOQCatdrfGC+6wgLUf/yRWp3wN/9PpkQThSVHAhn5ZtUZL8Jo1xhTdtC+
+SIOTMb4kYWoj5EghkE5AVnyu/ABbUvNlmjkVIqRPkUltYw1WniNQN/aWfttwpoS
1PcksFJwMGXZ+ndE/wyPE1DwCz+IkzlvfnFGcCkZ/6jv01+2Ic/WTN7mmWrtiUEq
LumnfnWBdnS/gqENBuisHI+RQ9bUCnTleQ/xLLxIK7tueSvv3dFD0tt5wuufqdzx
/jIf9Mixl4h0IOjP4vqcqC813zfSZLn7S/EAiWza1g1rRa0dq9/yyOefJ1tjQg7F
UH1tLTAjM2/u/nVQl+HcC9u1PcgT0LTBEnBuzYtHQsalW3Nwwjc8j43Yatb7W15E
2wGPheunbQfXNTavLh/1r/3GDmAjixzqzstGUVv/II6N5basISW5v/bkfnk/d74V
LslH1waqQVv7YsfizBDSdMyWaCuruyGZrHOrxrW/5maUneYtfC1oxUFuYpsfg+hd
ucWHXfON47C9b+qYMcRR6/rnub70vvT5wM0B0rKj2K91/JOCeGq/tiK9kfviHy4j
rrrKx+riErVFde8Yv0QwYjeTqHnUFdZGk6OolH2wdJiE0R5/t9bnRrwtiJvYIxhW
E88um4T7w/yo5MOhGnEP3NAHzcoMDjZvJdjCWkYp0zpiRIgIPI4jKtVT47w4KYcH
yjU0OugpuO4yvmcVtfcrWjHPxHh/JMbdy1SWC5fHjrM+c/eImNOmdL1FCxupo+Gj
ptiQ2+kS/LZVxs7ZIkmR7NtbAZ2jFHoXaQTeGwAEQy8YZ5HFiTnPVY5GEgwwTEHC
Q9q4WlvggOa6vHftrRJt5aIZsDWCwuEMr/iz2xByn605BIfJOETl5Vo6rH/O/mIK
NnmJpBRP+4C/sUsSQf9tqF8XpTcGuYHckzU29Jnf0H4wJmwUJfVBIsHQcucOYY0V
VSNCqmVNfkQTkJcpxnpEj2vIrn61jvksBZN9tBIUFUz/UmV+/TojWKYNz6/IZEhP
lrgzL4uW2CvLJLcbSDns+vfaFNn0iY9x8dGS0VNNYgRO+uwIZ5vakh/bF2idAb7f
YPQDKgxJTpXoEB51RwsMuIPsJnTy9wcqu3EDpYdkrar27dfGnVgcSqLYQMywzrR4
Sv29HlzTAFyoOZqUMa6hHvlj6G6rt0m4ZCVR2tCyIqfUBBqZBv+91l1T0OjVokdi
vfQsduWcRg3vJG26GymqmF9ZRSnRfIzZSp/IvMz/5syoad6dXKuVxMcMa3DhHonu
25j0GCHGMsXUFv5nOEdfEDpMFsapG68PmLDYeVzmFTanKjZxE6yqyJtkvcHbNU+I
3PhW/Drh3AzUZO1V5Df8yZO45WWveR0rZIqm64bFVL1JF5tokQ7eAhG+S0E69ftc
4YxUf+9ByG5UIECx1BIzbYQJGMHHpytpY6+M3dxhNwm/GjoOFc3V8hc/ST5ajKgQ
zWocz1/pzBecXO/trBftytBtloH4XVFw9ruO5XsEW7nhXZ1n+qtfuvSO5DG5IPB0
9hcH96YoINmqZWD9vk18nblQlAmGB7cHs61aZ1g++aBJtsoTni6BI+nVXhDE6S2b
RrZcn1h45ACAhLzACO70ixGDbWVLONQTnrnbOIgeV7ub08Y+agYaWhxns5prrug+
BP6+DLsOaHvpbacc6NG37A8lGzwBEtrOLuC0Op+ZWq82JDaO1TK5bVL/2evhFxCD
cbvbgo6xqrCyjZLjr5ZAWiJV/9o6yebyYbRQx1GbEhUxrhNpUR2Aulbd0us+CB5A
QISLciXWI16Q6vPyXGKhFqaTcDzMBYMAxlH/3VnPwIj0Fmln0b+NQW/eX7o4eBMC
KIN6yjXlGBxA1H0g1tfGqlEziPultZHdHmuB2C1OvBKwPl2GMwCfyJNCdgLnDs21
aZr+b63bAApBwxEqUkt5ybPQ4wmlqgUK2mtFxXl/c3NuKevU38FsHbCZvtTnov77
Oi20fvsXZabdsTiu5/gITxrbKKeRD570w14Epuc/yXR3YmWwfeGZu5eCA2yp4yUD
EjfxdgRFJSjt+wgK8GSu8oLTh8cKPhWYmhAKvAMJoMs9bIYnOVxpkQaQhS8KJtOR
/BRIjdl4pD/dNSF4NFHDnUtkoXHA62P6PcK6IvQDFDH0aratMKiiAsl/8rYjPgxC
I53AkqQGUuX0Ww0AGAsKam6TOcZ70UHet7DG6i5S1a2/O4VZJcM2hpVv7n+SygrT
lq5mQ9TZwMrgMNwJxMPO5pGb2JOsvvunqtOhp17dAVm+kIcq1RJCHDhy12kzah5/
bsvq6uVgOi2fZVtna2tcXmBdqmt2ZXJKi9okAmTtM3Tmfz8yNnYklFG0D5opfM7F
+ccvy6NIMBNfBP1GNwTEpwlrA7SM29FpmAj84NBrWjEqJRalj3A9p/rMmRyjFu+h
dQ+R5PL4hryZRr/LayCMnNvTWfIuQnd1ckEu5N8qmVsBnl40bCDvpI3G2OumT58P
MIeW+ato/PGlhvoOYH45UZF94vYY8gGj+G80mLzebdDqaVeB/ZUihTHv+CpTx+yy
6waFotNcjQ03A28gX+x+1gfu1A0sxiqQbJ86oZtmYJCMcx6YHqDbWZIkS812EZZs
URraIeayv4w5YFQxAwJ0IXLaDFXRO7thW1MLN2LCCxl7XOH0INb1kOjRfpPQh5pQ
tEhxzVehgGPyhENRXG2ZgHq5FZ8feOhqr6ePnI+d7MqnHjsTN62GdJRoquOp9n4y
AEfUw9H3AxZN+lEnaOGZOoGhwAjFV9B5NsEZX8LzKAr0eJqbUHMcJHniCJWL1/KA
jl8liGC5uSNN+rPkbmOndDT19wg/jVuRw/X+6po+jq5nyXO4DdV5jxPEpfTO3FnZ
UZDlWrnfiYVnpwo8dIaluU+1FIQbCaJOKFpDT7/CM86CcdtJTH/B/PPmBqCMFQo7
+DyPgHMxDwfgecEmIoc6ZkprzQpgs9oMN+XxrYPj6iCZEzrB9RGVKeIfQQit+GIl
w0ZmuwTB12GKlSE2ndZz4kxdzNGE4N+dv6f4aXCIfxWw0uATpAhV2GEJAtDUvjkI
8yZam445AhPWMQ9Mug+sH+TrvzbLUBSrtD9gfcJNhYVKC79BLQSA1kHq8oCL6hbn
rwJaU+7VleRCl02PXoJFnKlSxUQLEoMqWy7FjGO3a53jql11q5U79/vPrbvxWefE
ivOff2bRjiB6Ny6YALejuRwlRzedLNuPeeX7ykEOqMqdQMUn8vQwyScH5Gbzoymf
UtDvDDKYSvOluk+Vu48XeXrV7wx6bMJXHsNXDfLCS8a210Hn/pV9ngQW8qaebi+W
ug2ms+OiEqOr8UP601NVypGTqBLzeItqWsu32YA1jO4XZERuxmZQvGLfTMqKESWn
Gu+l51ZaFf2WtPl2q1bA2AD42bTi7So+yhaPoynFopGZ2RSx62vGMUu1o8tUUsO9
XwF2uk/tMlpjhdDwDaTbPMVKF2TRfuQC3Xs6WblKL0XFVFTVen+ZOjNEMYm83kRH
bEieLM+YY6LGtKLuZaPURd/W2cuV6jRdofDichbMZ+y3TnlS9YumVb6EiqSmuqW0
hP67ehnTnHPwL0OSvRem9do7V46x5/YtLUmhQFs6I9pTuuE3b3r+co7pbaWP/sya
S28nVM/wLWC0WJWHf7xNW4jOF9b4qn3z3+GqWDLEML3rQahpap+D/mwXVBWsTzG6
VPm0R52Q/QQqa0ELvM4EP0wC9fYHasPVr0hOMhWgLUdaRRAMRPRfrpdgi2AWXtmy
JMwIgzmBHahpxT1xIhkzLm41oqVL79hVsxoARHjqi8uN4mgvI8uhxrHNC7gYwnkg
7c4HTRlkzLnp8AD4ezujM6uW/u4sOK3hQI3XGP66lH2RL8Acut88UUNb4gMbcJnj
Z/RUBa7zSx4zrY/Low9RYXqc1Omgx4t9pu5inyoiEh0g/YH28wtTxeMnJ2sx2Miv
HCumpEDIIUDCKYPQVd9MINqdzjst/yWG2mkWnWCPKKIBSQqLiyEG1feQti9rZkrg
/9jtRFp0KV5rLPz3t6rqqpVn3yGiIXHIWdw6hnkHuz+TS9Ww/CzP42rufrWrWH0v
OEm/oIGVnd5t9dq4wDhM/KP2pPKGUMtE09SdeTxRSkCvvtAP5TFixhx//19FJKyL
85OhntDlVEfJYqYMwm/mAoIR5ls9NgV5qf9pEbGCN94AGQafVHvexCuY+3iqQeJ7
4H4ZuDhIHRwkN4lBzM2n0/gJWzkvj0maYDuhYR/VM0B8ViCdL2FqFTgzzj81ty1w
MWhzCA/OZPoT/NAQs+ggnSdLniQ/9wGLFE/Rn2Y/TimAQz23dD1pboHMS3Er7UIY
25nkXQSorzq//Mgp61bmOrWbMc6hOae5dqDkBy9BIjD002fJhWKgnewD2yZi0ukq
KyWll6AfdOc1e0KIA0Z17NEYLPZ/5ANJ/ox4jV02O2h3/Kv4OzOgazbb7ViIlyPF
6Ik6MYmsmt4aOKW95MK+gFUaJwuHog+zWPDBB+KAM4C6gayN8GJbRLsvc9os6GWT
wDhpPEiqy0rkKOl9Ejx/XWldCVaECKwKFspGtL/rNvWfrlFU0d42H7ufmkrnuaGJ
zCmrhVMpWvt9ES0nbtF05f2cn+fiUuJj2pwnvawyHW/z8wMIORJVvA6/Umgn9XL3
P9cpN/iAzEviqEY/H04m46tz6l2oOIPmKeWhpP74a0G/nGEaB79Gi3xV7tvGd/0e
c22lI4y1MKiMUvyGLuKKeiKER2paSmWOT7t+vxJMgS/elacmWWyb1H2Yv7Tc+bVi
6MT899hiATAxArCkJUA1Iqn9tSm46+HA6LER3s41RVsWTqsLxNloT4OKjp/e2Xkn
r3PH2uFAAiY9sDhgHnYHNGeHSyTL0xXe8xNYdHMubj0edU75nBB2hWX+J14c+3gZ
DQA4rsumZ0VZYefCG31BF/NZhZppbqAUxK8ycGF8rGk7L0jO4Z7y04AfCTIVsLKj
ONkw4yz3YCmitAW6fEMJ9YxirEle1FJqVK12uEyEiNHGUtmyk7ueo+Cxg8EDLyN7
KOiNjpP92bIocDVQaoKCWxpaItfGcMHxG21MSUPIiobpvkmaJceqLQoOLGahZodX
TfIGSFzBm7wyj7gjz9D3hB6QuFt1PIHgS2/aMlpv5oOgaLqmsn9quaJj0Jyn42gX
W7Od194JUViQcUbSWBqx3ArpJveURqZT3+boTuqCfRgTnoWMKTF1Qtx+VIJKspZY
tdrs1IHdAsz9g+/dlFHgkZ38kcQ1z3+22Jm98hgNFHZJwFa8QVRQC7FzMANlt3FD
a7jW8A1d0fwTsvi+vNKsZ++4wvk0UIJkJ524nNLatMpq4ctU70KRSksKOiPzu6jU
Cbi5OlSYjRkMRSb2dQ4DNM4Sp0AhV6fjFtA/9v2umRw/mRRHWkqEfChpT+xjm5sD
/A0xBCNrgl2bb+lJZTxP8EbwL2K5TZSfE2wDGhn48evwKtZH+uZWKZnqzbDZ5qAe
6ThQz05uQrMVTThJbQMLbWHQeFctANjSQ8OD7ATs0aqnSMvZROOveEbRdPEBL+zy
sU5SX9bUEYUb4V3N4tv1hrz9doKtsCynN/tLEn7slFxSikZiVgKoTnadC/UQ/+Bu
GvT47WbkzXnZzR0KgRWYrxEnt/NFi7sKsN90/+zKP6OGlBp0raxkVzM5SfmZfq1D
/9YMiFB3t6KfeDwtKfJjlDB/EOtHjvt291RbefeJ/O1iame7df0mvg4fy/YeMs79
viv2aYeJbEY0Q6RsIPx5iBnyriJhoseZBO1OPiSTr34jWEUJ8/2TmK7t053RlKsI
4LXqvxpaQg2l16+/Y1QBmgGGVOYEZeHmdtTjujCgcRqzzRDwHcG1qlE21bIBTFxO
hT1N66Sam3uNaH2Gvl0Uxapg/c/7I3b7dwZh75gTqWvQtwcMUFeu+x5/kpzrzBsu
0NJK3TmTiHM9DouU7l5+ozoYeBgIvuZBKrkMezaB13N9dWZarp5qRZHqVTuDIAhA
bpJWlz3KipONlsFaME3fTBB0jx0zupROK6EUtEM/KXitw+B9zz9VnrllC9gEw3DL
6Pv5gXg494muHujd9S/1YD0NOe/AYS2/3opykmD6uB/PpN1smNx2b/1J4rLN2zWP
Z5I7fukYgZNCs+3PkJfyqdXlwqgSsVW+kHTS9PguHZQ7WURQhnkrSFb1ntjagaTt
3G78g6NifmP+A6QKiFd7Hyf80FKzPMedxxgWRvTTvt7D/BYok1yMvfi7KAhu1xYU
Ww14XlGLH5lFpJBlM2PQRcgtRymYhTO0p+ppMOjQzHKn5/nwFtHdmYmbUKm8t4vE
hhBIE01bc1xOQVKUSJkgqduelHUP2ytekbTONX+LR325Fuy4xWpgNyB7rmc0rj82
faAJly7YdhvQ/0auPkWoEN4NRH+il7tLSeTyJL46OwSeKH1/YAnri9kej/st20Vs
3IjiXOrnsyxMop3Frl7dbfWI1hglSx2LgzYTFjI6hkVEFvZ6RvbPvaN/Mj2gYhDO
0pAF0iBYeT2Ug2C4GQnZTV69IWpdEvmzGLvJ617YKYzFLksTNoEQ9zTg6zfT0i+V
dDu9bc2XiHTWy4euuAgn5ZvGpRMTEdbqnlMELMigR+xiQ4iEb+MHY5DTAUUDOgZE
XsyA9sOuKLa48woDFahQiPMvO8ErkXY2quiUdask6ZIiQm5uQAONJNYxMGOdFdas
9uQ5fAyom82eC/Ro4qScMBcp3kiR7h+MMGrOM2L2f/MG6pBPPaq61I2wubPUTdws
gammZzKPIc7wvel023y543gRwvjxdR+favIPvWohAgF6aFJctW52Msza2YQ/Usc/
TU3XUCtOpwlyQRvIRMB60dRXS2uJvKwgTZKAp/aGV07GaeyAhMvjL2YT++KPGv+b
Lnf507gNwYRCCBCTSpGhcXReqEP1IdlcgZ9T/p8b1Du0nSyZXLFAr6yGDb4mRdl6
j1g0M80pi0BaSW620KX4VcqxLTaGN4L1m85nUNJnOpZUyF3eb/tEtftQNU/Y8R4i
+2cLmGX5PuXNxZU91ZTg7GyFoGtlsf57hHeVXLAi6stPnedI+ZpKJtADzGQvD44s
MVj8HB1g/kCG8ANOzIgtxv5Tw1Y+JZ3+cCrMIo4kMKAshKSV8nVUIjNy6mbpx9sN
nfoHuFU/NRFqOYlC4uyPRrsUiS4eWnOmUx6h+Gkc0yIwQPQOxbyY7rEHKE+FSxLX
Xs8lYvKQsWOSNLM3fshLO5wkZp2lWIE6QQ88ktt11bwEPyBoCx2wnrXX15yKXx4S
eIOPeFDFK3annL0s1HNXjaktRW+7rMF241lieGVpwZohEvb6IU+vl4ygYpPC5tHX
C3/2uiBjTanPzxgIHAegYk2ZXu+0wINaviFthiFan0eX6iOV5TLpYCkZ9l880MT6
WtNv1j1RDSbi48iO9NmkA9rXaUYox/QfN8cwKJF7fdqP6J31UgPrgFXbucMCJulj
JTKbwl3BKEQGCEPrUJv0lcFyhABp8C3srvCzxut1AZ1EK5WMLZJ0GIvbsYMip+9B
p7lnkJobWKdLDKRf+yPk5cfc+3iQfBZntBjyKnP4mRukA85KjloZpC5ckL8zmV2P
SE53myfJV4YWoF+/Za/DgaDRZgJDNTAFiJxJThJ9O6gSx+LxicTL/HEEZHj/xg5M
rQRR6xmJ/qjlh+ERIb3efaUx66bYIdxgSuHzoSPK2tKbB+jcvJyYCOL5dxeaAS9W
TqgRLb+yWJFIIppunkCOXZwydBbRoLV3UPWoVEC+oBbLT7TY7IXO8ruHX2E13Q9q
ze9AZOHpkfSHpQUuItCgZLSNdv+UVrt/Ug8tZPXLhJAC4M94pWu1i44ShGeB9pqc
rjMh1V7p5S6JffTnHGEf+9c9WLSGfVRgyAVXiy5mK+JvAHAhdUqvhiTbkyYn76md
ZWKCqD9T6ZkPQFWaiQzfdOHRTkyAynm7HqB8Ppcfjn7H+Jo6NC+9KqedVgqS0s8y
Cl+eipr2B9m+o5H3iWxCGGvVK8bKwa1sx1llCxYMcili21rEl9SDry3Gj1xo5CF7
+rlkfh8i4hl04IWt1tNOfQk8Q7lTqhwo9JusZMLOFm4TdVcEfhnzK6XrLatfEkNu
uu/9zHk6xxiHQ98JMqcAhuRAPUwBUtWVN++MG4H3ELKOUT6u8W0r4SkcFD/GSFEP
VpVPHxyCi2OW0BPEbanDltSEDqrbUCj+xR7YWMfAF82D5cBZhXS9qW9ZAmk3Q2dG
cBPZ4ftXdQxImN5fOyb3h6Vl05XLh/eAjT3db5WIzZguNDJzwvY5dmCmuJ14EN9p
AlQNmgbjl+bDDuXPlyj5dDA6CechkexwzYE4a5WntbqWz/+nO2JYfy+P0gxu1F6z
8RVi9OX2kjb42zzZLiBBGugQIKcdt5s4dUFC7OawZdWCm6LlyMF1mKF29dhHE/Ew
4dOnEBYluXqyCn3NKq2cqTys+g5ZXsmQtTJHTai4eCjB37qBOSymqC+ekEp0wJIT
u/RRAO94JtFSNY8ciopumIzseOPALfLKdGf3baXnMRtfouxLIOYEC0qD4tWyK3WK
o/GZ5IYUjnqdpBKkJnAGvyivJJ7N7a2cH/hP/7I6ezuJUJDs4/jE9JOYavbWWZbc
goVhakuPTmG7237QWj6hVr4zaAceU/U/I2iZE1TuLOB4nZP5D1dSfwimC5tJdQM4
Qr8qsI5GVNr2t9+gb4q/AF5YBm1xqJztc6hL2GEG2wa2OzoasIU1KmjoSG/Rg52X
/QA4u8Uw9ta/ABtxrXbme0qGha2mAFyOrjo4LviWQdinYACefAghyIIrJ3kxlCXf
xE/jI+JQWDhC2AxICHQQWrBYa7VMGusEI8u3oC0+6nxSPEZWOSMBDl/ZpiCfgpKL
pPwTiMbgWW4ujFKfdFhuKKCVucY2ZlYrnY2xFRsNFq1wN/YPc9tmt6l/NGRBXDXo
TA1O7v+EPMYyOwW+hSqGNe0XlRplXVXHylrJO4kFeB+x489nUP+yGv2uzBEXnyCH
Op2mPfNkImP241PKRcfbCxOQjW+85aMmd+/Mhhb6556utnncE2THzevvhroG7bGv
8MGgbw3DFvoOKzmSuuSG47xruqoE8+AoTO6N99FEm29Vfc2OtW4zj43s4or1l1Pm
8daasSqoQXE/AY1j1wXJJYsl+qlK0MfdtMtfAUZOFl8Ny+BulrpwQggIsRfxQ+cZ
Yat3vhbvPLG/X+tPLaheyie2lMRr5VRpqQBkWZ9ixukQuTQO1zcIhK1Bj4LHOMt/
Y+gRRq3KWZUETkaf/wCgd8YJqk9CYR40sMBuZxRJXJeTaxfrfVfK/IM4LAz3hpr/
7HnD55ZPuJ1LtyWLZqhxvqMr+rcC3wvqHRMDE97CXSLDOi6ogWmBatdcxB7FtfuH
Hy4vJkmO+rx0RwwKKxV9v3qseSIhjoCw/59HFJ3WHHwDQ60AzC3IZuPIgoT0j3rh
vIKpvnzob5D++jaCoVeGh1V62ceMnqD22qFzJV+GsrBb50K3+Y13uSyVm49z4BOA
jN0V2OMR6WQZOPJyYbFEKDpTpQvut9BjiN5ToRVup5jTRi8lUp5Pjad3NjDMTXDJ
N3l6O1s7BAOcBLthaCkageuxJ00CRgqCGE8R1IkdRhM0xuLum4Jdpy89E2Tx7nOX
2k1bhN7Mg9ELxFdobzN0CnD48DNNDfJUqQlRiIfH6Odqk/XZzgGj0i9qjcCxE7QO
krIuz2V7q8ONYU9J/HNDkgNlrD7BEY1ATDZjqD41iQWFGcKgcoMVJkt3kd5CtxDK
nydXSI15nqfpPOsDKzmpPTwa5aZvWpGvZIJYi2vTZpbGLtCrU4YaD9BqLQVwOK54
oBytJUv4Nj7PtMRR0lVrshenHkNtMG2z/NGxM1MDu9S+HYcdl7eIKKuJcUfvA6w/
jSVphBkX3zlSsDJIHIeW0IuwMhU111TEfKbskCcVqrRZWDzH0Z3bLaUyu9bbLHVt
9pvcKqfKluXPnyEFcobHo3B7xw+FWR+3H2su0yBdkobDwXk8gSy2RMW5mhZBJH7H
CmSx5B7ZU9ekKPmxpepFAWIEhx4nSPI/pElfeOgEzxZH5PLPB7jizqk9zCvSPmSM
ciUecWPlCAVEQ0ltC78y4eoZmPZcyGetoHya3qFw77/N6g2hwiaLQR0BCMP5jYn+
yywWQzEVWWQgpGhz6kUv71QEiwobEtBfdpWs0VC6oX4seuQVU38U5layeHKOIVje
a8Ib3kPp5O1mnkbaGoq3g9BM7+mG8sMHcCYANPlJFGhEHHfUaCwguMv3HhCy4yML
XoIZca/4oQf14OIGL9Q3rHc95VhDLyOrES6uB1bftnSNDr+/wDT+X2oilfZW+nOv
L5a/JH+1uhZ5co5M4eNT1tOHl1VBZxTL2bXSGHC520QhkYV089aafu1RD3B7Ltw8
YO5RL/lsZdxbKRws+LULDL1AEfJI3cFC0dc7zKeOYSJ8V3XSavTJ0kKfCzXK+4b3
0GHaDsWfZHzsQQdYusA131bJzimUaE6svxVvBX6AQD9QPi+9mMZr5NgoCo1nDjK0
p2rvRQQBspQjmL18AextdXI8qJS4H1nH01/FRUJa6ZAXMM6FNEXR+heusaiDPZW+
OzOHDg0DQHUzTGUosgnVaaE5cm7UFgr3AtNHjwGF8zYDM5kV8bjbtguMURmbe8ff
wVlbgiVCxOiUiqQs5lIjF9wuEWqTSN9gtiEn5cUmDRtsdQkKJxhufXEBGlt1WmzI
4YOBiCrgw/qg6pt4zqjVAPNraYBLBDiBwGG2NQblKf3+xa0Fc4NLvAlNSrFvHhbd
5N0yGkOZMyapUMa/qLuRnNbZ7SPPF+uyDwIpEkb8BXpgyafcRiryW6x47R/66v1T
J0VgQ/CCjokTb3Hj3jd6trHgqX1anxa9s2TsLUTu9ZemyyWohYKGbuxbZXceeFCa
lm1SqD+zNUcPQZOfLhC/iOZOga6dp6f7WEqNYltUTG+KVNvkhboKZ/3fE+BZxiZO
AMTQir3XSLMgyJjfU6oMcSVJ+s0v+AIMt0JnsCwm9O8DC4JDxqrRQwzP9HrJ1ms7
W81CNOaIOS3kwzOTfrNevGhrZDMuxqlaGGETYsM1FjQL4vktMU1nDrQipJlGG6lN
moq/dAmRB9nXyZM48tknj/9zyREvJN13JcbkvD/lq64XvXzCZXjDzNjZylWfV/8C
Ybx1THa6QVKohwVCTDH43ePTfkyE0x8kzSNQ/hg4QGaaPH2XK76t4Og0KJIowt4N
SXjgtaeRj0vb6j5AeAQIjbnDgqgvxzqtUB35+no+pLgOgJhislyxtCNz42vw3BG/
+fW3IfbYlabYCA+mRUakUb2lPE3i9C+93/jmmRypkXeExrt+eTnm6YM5nGILLRON
Bo5aMH1js3BjUov3/sFwpa1oGa9xx5rsw5zuF2bi/ChHC+f0Pj4n8W77FPdQFnMh
NGt/QbsJ6h6W739eqb/JQVbO+Ft/weCF6qWbwAJZlsu9FySjyyWeiljG+07NE9Ke
RKWoHlWuTGZEymXhg6xhKesV+YsnDDA3PzGalzAc1Y9wTEu8fUOKV8Gyg8CbS0c7
PniomIweeAy9YlyxgXMKm7ylx4mCxwhGyVLAGS9dAiOH2jPvNR7VbOrhHAxIuDGy
/LqBwh+bWlgcIjyuvKkLzwBUNUrC42syujv/IlcklyqHY4C2iUsyy3dF9aTfQDyL
bMcxwG15hhPf0UQPYKyrBgyUlzTN6lpQMx1oGt9V5dwdohV/VUPSyK5Ih4KDn7vV
gvXF56TGP26mwOFGBWxufAb8HUCm2xwV+1t73krBhdKuWEzzVrKsvA3OPN+VSw5y
uSZizxnB/yuE8Vu2RdMQREOb/pFjkpqGSLBxU9BUfNDKfrKzXjZyHZb4a1XpsznE
ibP7kWrbea1+DTkPfkdBELyI9dhQ3zYjtKVUcQJuodi421+ErtdZYfjt420rtk15
00TD/NKN/9Eo0Mv/Cdvu4CGJVCinJ1TC3aEsceQnRtrttXFw8Z77SF8s7l32QAPw
oSdrc0hnCGiOqZjHsNTDZqLSqfOFLMgus9hhK9c/5/bmRXxgYWeDxqLfksyqxI73
kD5oA/DBiRFUGsEiE3Io2iPo1ZCFYLRkFgmyrztqZckQ4Asq4l/CAjWI6MBOME7R
kyTWzbvCYTqgTSo5W322rMvhQePGAGjjg3Lo87b4VaI+H9kFpoagQI6+Y3wC216d
p5/BuFwUulgJOGuhTwNVqRrZCcfphyyDRiUJllSQQw1cTwdDt7/AAeO4sKsTAgDL
06Pgx0WvFCRgbgnAQ/To26eXcv4DXAHieiut83SzjTfWRwzipfrlvlBO1fXTrXAc
kUzjUDk0TyTustDRZ2XQRdlRQDGDj/16wCdqrNBO+42lLn+VCqGa50tb2PJP2PxQ
n/ShUN3IUkDAKbuasyVc7bMa30B0fjEgx1SIf7L52D1QtYj6JXRRoyn454nOEW6T
dqJ3z0jhpkR9KSZfrYnloU5MZ0eg9LELns7yipTxVPRUXswPL3NJ3znCb+QPO+Us
dfguM+Q98BJwVY1jS+dBySHqW85yEiG0AjtMZe9tdZRXDyNmVirIyd7NZOCPf7dG
DFpuZ5o5A4P/aj2VpFjVThx5jsI1y8vgzod9mcsJGrH55FT1ef6W3R2BDuUz+4eY
z9AWJJbYjDlVtHClEqezy6WiYb/DT2ldn1xqf5Cbs7WNBwOM8DvDn5IuPNZ0eTfZ
cqzJZdZN5OsIGs909j8N8PCUjbIvww76iUj1dQ4yAzBEb98I9s4Fnf4cpasjJprm
IHq48IIyoIprGVJY/xA/hU3YWpgNFOcdFMHChtKNjMTEb/eBjri0nQCZkxEdwZrL
qSJBNs9WafiN+merStdHFOTUIDjQ3beiR/Ur5kfZAbc/73W1xVRhYeLSk2XmY4Z0
r27U3xGnVuBb/yKvlgefc7Gmiruj4tWDgJQp7wU1aYuAysJDqh3pggDyvXW1H3b9
8dygLecwnJt7YokbCgc2padglwUi0pNSlnkjLCzI5qVl0I66qjWPCUx3Wo5vqMjY
y7WcE8vn2DUaTq4XBJYPQZOgsACLBj7n9zh64lmQd340d6ZwYrLWkltpuG7dlmYW
uviLGlp3krFcvQz1Q9ISIAWPNgvCTo6FMlOc+4aGWN499wU/ftAIw6Y61vbRbDhl
WADAYk4XZa7CwrSypjfT5mBesX+HJabTwUQn3/7ndbA5Fg8cww1M7DsO1bSB/0aP
n1fr0PeqVFsUg+05PydfvDZllJqAwYrWGECo4Xx1UNu8XLmwKyjYiecPRH3cs1Ub
I//db0Ev5p2GnS0HaD7Du3HAn5uWu+3yLx5Zs+0SFWpMFJv65O7wuJjgdlrqTU81
h8tPjmaqfsTykvfDAc952usEY2nmZUueC9ghhBh+WMSkTCErRVJhx97oyF0KSmgm
D4MXLFp5tNUIeHDS4nB14Iy7ogf2f9CtToFFeJeaRkGkdjvhP63q+1kk0Lq9ikpD
egKf514DnwT01F3nOjgNnE/D4V8cGv4nrjeoPU6x4d8TqI8OJPGN7NWpjk4dFy4T
6bIixRjO5wJv8ABFDO8H4FoaHCR0VMMWSUJcbe+ujJRX5WKvMbPP1bs/q2koTqmb
YqQHLJwOXNCvJCUrjhX5G9LxsOU4VBjLdptIS3n6pfU9X0DWR7JrRjOKCTO4CPOE
FXRsV7LzAE/5cFJHPsvtHvhKTARQUNSxMhx/torCP08GXwEGPA2GlXNrusEv3b2o
GNKFWHV+2miQs9QLcL9pxu6OdwJpLt+N+OE2ukDLuyYZvye678AV3f1g7RyHlPXW
DHYRNtdwGFNS11TmXfNj2sn502+wcQO6gaxKd5HokJimJnB4xKt2R/gyFFJvVPY2
m4Jsoh/R2ja+6Hil8zw9skAce6QQlMjx5mthfYMdVWqGV2HCun+5H1IzGWpm/AHT
O32SRE4sKafbjP0JdXGg0+uCRWveBgY0uVkKBfQ2jgvjxANRSGpUZZkfV5zFnqa0
IwL97DBwZMfcjE67PRDyYhXQQooHhq3V6ZtOGwDJu7l9QP+TatomP9jfT/zPx2hO
iDqlDflHGSimHYBiTzPlBCwHtmqunfpqPzdcYNqBE0u5oricQ6m5a56E7sijOIWx
EFD64nI4F8cs6J6BeIltBbQvKzzA/3Qj5B9IxaeY/KZlFcpjBAqaK1EBSQ6rqjhA
VK+lnAShMPPnM93DjnsfasNxS4GKGcN3p8akHQGxVuCyICuFg+I1dA35BEr5SsLK
3lSOsm8YPdH/XFeAH6Hnhh/yzS/bcoBsjGyC/PsglTAF/a52e8J6pOkxvxxSOqig
hYGh5aWt4oVqlNnvuGUgq7j2xTNNDvJ4kjfVslYgDiKh6/wa0YqbqBSOo8iEAW/h
q+RtlL9LySwKoiIOubrTYidLcezhWMqlX6ACuuBbkUFQNWTABm9aqo8MRU4snOGs
TbwzdHsQYRm1cXDxKTPgzIGbo+XQJBPLn/5N6FRfyfrUWom0zlla0l9+Ozqzf7xa
nj6ll/DyjlaX7rR9Mm0p3tjdaGMmjdMt2wZYY1jS/ByVV3+RSGVt4/JuCsMb2PJF
pRRbHZaf2hNZD0nTt6e8hXzjefscCrdNDr8LBekYMiIC8I685Z4AU2PMoLKLFH1+
mLz+VrURtPxvY77Lq3h8ajnNnNJ+lxrnjY7o9FTUVUWaVjzxxsX5GCYFGK4DZ24q
SaWZObjqENkMHIFL2g5smsW4pdiUYUSCRqZvVrPEWY1nR8UkQZCOu5mAHeazkCVq
oBCa1RxfSbjhZl2MAgwTbRRyrX7MBuFf3eXtLMkKGMmptDP75u8QyDm7lN5dFzF8
oRkpI8Tj8acmGt6trd/hsnVloilm/XxuX7gfCTGe7kC8uFloEYDKX3U1hPkFvKSi
S7TjAT8CAp+oSKu4p89EW6Ev+H65tvXg8T4mmLzkg0J20VTMpjqUjHTyWCU+kQ4W
D4XIgGnSOEvt3k9q1IUvcpLtAqGUr7lZFCbT4VcjuNc/bon9iHtKnYXgSiZXQcJn
RHJ/0etN1tuwD7MP4exeZYMwnnn8vs5+xo0YnSeoHACoLsaXFctBgE9Mvww3Cwzy
Qa+td687ixOxHKU8fANMgFhgRATlj7RkeGGN5peLOushzciEIrKrdRmTwZxTPHnS
2UuSJ/4tuRwvjuaG7vaJgND8zq81O7Jf0cBHJrpisgfLuJL0fbIV6Lxe5CdBXU/c
DxO51yklvTVjW67Ryicsh/eJIBQHLRsfRXqChZNaXdAg0lcZAVijB1cniLnKoi8R
es03z+qwyXoeUn8NmP45s+32h/4Q+EEmA0WU+aOrKcl81MqkH1UqKehrtfhrEbfb
jbHu7AuwUQj47ia8jeEER73ZyF2f9Zjz0V4aT/F5LpqdXLyalPo6cIcnAzaKbelr
WakZy+lIYsiYVUf05h1qCyuKunxIQ1/E/wy96aHlc5xtUqC7eb3lbxqVxD9JV1b6
KHojwXTT7789VDlvn5srY26p18dDrRRrSIlSsxC5S0dZxQJOk8jSCfTOklTmBmLB
iWUv06eg52b8DgKBsq6Y7DfanONf4KeFbkjUJHv7rpOFBPrGiB/0kSq/SYrtWqG5
5OhknMcx/2Y2cWi06SLkh/88Fgb3HxYQT0unQKSdLiOC0zucC4ggM3fGYWxYsgjg
0eIL6pQjyxH+w1Wg/mxMRW+O91/+m9d60P+F1zH/DNTjjFAKSTwJ7F3mr5KxvoxW
rOq5+1KUg2m21tNxrMDNQr4zY7MeQ3n84RUejoAX9LAtLE8PvtH5N1AlPSzYPQrg
KUZylqioG3zm1h1ZamdtZGg6D+Ta3QCvyrq2bfiFtNLzMzFig2l6NfyNECqO8Sxd
lhNFaNNNsZD+0BG6pyCa/L91C0N8E7M9JhyAL2zgF59ojS52EaQXXk+Riv+beKl2
e/KRMEkSd60FWihpdiUuZ/+cIywFV9yqmIxz4vg4ovKZEWPpJYhGQTiM+PFz/gQ0
XTf25x9wsfDtVXdFhgJjv3TqntU6CmcwtoFkOdjhvkCTJUhmSJXnAADImO7zeaXA
NRol2gbW3PS4LDLMCihybvG3k+gwPleK4oszTIhCU86jft0jVpabRrzwLWtu2vLd
XyU+r0LBfHZOQsPRPeJqyuRHDfUK+W/LLWrk0ebp3V+lMpPWoqCIAX35sWI58E/4
TuBvKHysMLhHYty71J7w8AO4d3rcvaHmbrTUxgSGehqRQsx2Kc/yD4zL1ASZ8Ew0
/zzUdA9HftiLWsKzoy1d7MK6gSbhs/NVOexwM25ydnEPFAAS3VNqltEDp+rMmpKP
i4al8HWalYvUPXpw/t4AtqWqDId1K0rQnM14qA8pK8RPNJeBB7hLuzUcueeb5pRY
vVYFMsSNNWRrWyDZpEioxgX/vqjafL+auKeuPClhA2A5EPchN3Cj680b+M3LSxg3
4a7mN+cUq082Bc11bgFYK31Tb+8fmmPcX1MmIz7QwjtD/iMefkrCtaZ/RxfEqrry
URQmN86+Dv6uEpWWadenu4ZGXj/wGgoFesrxeAyopg5jYnfFq9oHNpCETrTsgtt1
hNkLC9Zl21CkcUhlt3bCFTEPmJnXWiwVHbrzUKuqqXOTdQ4QCs3k9/Bxfsotk+eM
Hdfc9AXREqHDONxnrjjjwxdUoHASm41IgKpHtbdbEHtrJNl7Px5cqRMeq6jx0Vsz
kWe1TmX61Yi3EuVFvBIqlxv+6W0muTD+XFDiuns/WzJA2Z136hMa/wRrOnQ9E34a
yj4gagyL1heOXVmDwHxMB3SmGO6F4f5q8rwzhYN4rV40m4bOOsqjaUjYeL5jDumm
7OKhlc3Vy9h46CeRwqXQUwelT4hPZhoTIi4r8vOkNNR0RQ7/saHjmkBpNpEAFC/W
9m0cWi1v+nOWGnd5SWGCLziFE8r1TXYtcq9UkOFRyFPeiofxWuSQxlI3SL+SksXq
ZtJArrgvtYbAzXB8n4EjXwPoM7JMniCxwgZGfnSsqjuiyUFxRMSN712Jyrc5Mt3Y
31JXtljxvnvSgOx0VqjxduGU27NAFveARJuOL5nTpOns/z2AmxWe0rMh+zUf2f0Q
2BCWtIP4oYj0Q5DiIrSDGKTEJGBjFLcb5KVYZUTYQ7gOOucBOvKhFYROY8xzgyrt
/GdYxHhI3AiysT4IrutvOk02ePv6oR41yln7lctw/aS4qJDm1bFt0v+DM/eCl0D3
mleD1fR3nScZZrxhvYZwule1v9c+MU4VjVM4Q20jT93OGbWAinaSrSCQrUdTBGbC
CUJrKWJDf2iRPAD/gedSIRkFb+xeolnidz2NngAlQrXZy0dT/vR3izaTEma9lmpP
NzOoWhAPg+hZ5s0ivMXfnhhe5NP7sBYzgN4Cy97pEfXuTNL9FM7QPzwA1GdPgvmQ
HymSGs5Q3gs+j4JRcmczlzAQy1xapx7Npr2gqLIu1S4WjKcUvZ7btLzWeoZxdu/X
2Vr3TSrM8uThh3CXRD2NYLXcy25AlaGaAMC5qiEDBp4OnvADfrACU54Eu1iqyss6
Uedfx3WFq/e6tuu5GiQ/culPkI+LNaRZJVkf54m+RVKtUvn+xul4jP1fIzEaS6pX
J9oVvJq5khFaz6Ht65sUQ4g6BizEx85ffz10+vuM5eVCEk5+W8rm7egSR2iIbf8N
Ke4Ogau3wAkd0O1FghLk3NjXd5FaETs8Kz8gK9oBTDq2EF0qtT0XT3eO6KHQ+SmK
u9tgkhGvttMMyTxdla9SpYrt1ncI9LxQx1trv1ETwQN22mxzWENNwZzBhilQWoB3
UNaYntEEM6JSyDoiXkf2d0uT6lcv2gPXNTD51NpokKechX96+n12xS2WhZOL/Rf2
2SYaxMLd59hbZ1iDA/TsCxFBSRo/oJp64+gkeFhTCcmC7/eescA5/C2D09mJzc/d
nlou6Y3LaHxjV/9Se9Jc/bDn26PM4CDhnBGx014VJbvKrdonift+DMJMrz8n4IEU
kmB9E8LotDA/vKXMSDXhRJzrlssM3CxsMDAXTMCkbIQKqP1C9Hw6ps7qrsLYehqr
m4E7dO/6LGUlNlIFX/yzDKdIuIgDOJELZZSLXi8vYvm08jUOSlRosA4Dqm8UcG2H
MehB6Y7vjaSaqX+1kxoE2EpmrZmkw5/qjuR0Z4O0mYNtxj8xhAO7z1K0RJSC8nXB
t5NfN2KeP83H2sFVwURZiYsBOtizrjd+V40LBp3eJlJJmsIPQi3KddqCfpuinlmt
e3DsOlv4u+EeoGoO53fcz8AsTNeIIEo1oJTM15GR/Jc3Uz6C3zhBl5zc57XH34aU
h0778lQc5Oj/Hh+wCJPY4XU3/4sWK84/zuAdplR4ibabXLTqxeTurixru3bgztRp
gbqM8ufK2I+TkFtH+Yq9ISysms3eV6AF5B4NAuc3A4pMLHdOiuTLiJh5nqNEVpyP
ZY3qzz5eq1mq/kVe1cdh/5Kac180wh0632qP8ZRhTlp1uVkN8CRZyWnL8BXX8UwQ
nwHsdVXk25YTS6J+gr0/mDKbIxnNuiW3sOgOmwE537f814MhM6Q1vZc+NHkaTBI3
Wh/APfTAUSWvmLD2FyP8CHeBHXFcHjX8G7jcYxUfGzPvZpjVg3P+tZVRdfMcnyiV
4AiTwUZEiC036asgT8Mdza+B85HrSkMR6t+cjXVnxj6axm+GDPSpW/kPuIwCY+Rg
nIGE6vCilklzhaAWl3Qr3U+6RD+3hsaA4HN7aZy9GKKIvjuXvejrLmKQhueygs3T
XMm53XoNZ4a6h1XDk1K0MEA2DGFtBmQYFmsgfxCrQNxdPPZRbhjuu0uM329TA74p
fonBX+yJ6beYC1rsa73hBB3LtJkKN6sp5qA60k5q9VNTsk9Z/5dEsMP68lQ16P9w
hrYKLzVbv4c36q5hKTz+0oFZ3yTNo+/eKp+MxmbIOTEO/4DlOhS1yxaWd3e/1bzU
bk1HTVin7Y8cUI81CQ6kt8umH+dOOGzhczqMPiKcvk+5UcsqSHS96R0q43O334Pp
TToRBHqMY4BQMP0RqaRN7bc35k2/NU/FuTr7+ZdHsMcUUMZ2tTifmbgbysG3kqw0
1OzWvi8224TWz6zyQjipwtzHJfSzDZiUwLjRAjmV9wPgezkTIQJm95wrYixjThUb
oHwhGeZROkD19ZfmjhuonFOzbkllfn8PAuGtu60EJ4JFHPMrriu5HkOIZMenPoyR
AdbzRwdO/9nxAXrafC41XkKXOYDSSpYuP0/E52kFiOjbu2YzeIxJ2RP5mjOrPAby
MQPxid9CmnNvpBeCoEgQArg3L1yzKSgORn43/w24kJhMGOeMhzpvPceb69HNz/TG
IW1Boa+1qyB1PTJ/Dg5AHZmaxlhqcHra2vaWKZTDykq27xgJ8VcETDs6g3f2LypT
+P0ujcUj9dr15ROvL2PKs1lCYAvdoKzfBpjz71diStzu5hfWu0e402mXRaumn10W
ke5slod73FqYeXF7GsUerqqm5yyRqbj5qwGuDEHqF9zyOayRH6RbNfm3CCwc8h51
KMnUKaUUdf04xn/B7xUFoCPdWQmpB+JgSVAvKpWNNqTTovcOgL4k6HCcnshis7jz
u28zLvkLhSTcKwnwM3r1tIarVR+TJWY88pqmnQz1OxtRdL6rE5UHg2fXPZ9ukNOK
loj8DBAfZvTx65wIcMFTGb5dnqG9XUbp5XE7GMMQvsjhMRFcjxgCHnMunldH8fKQ
MkLI/AhvywHYMnnCGf/qsNW/eARRyH1zUOtpKvhSAAWbxloix+gv7Qrww+mZAc6x
LiQ38w0szLNsWYCEsoIl4IRLg25qsskK9gvKRqdPcJc7A9tAuymcnrMFBs6+4WvA
TMg45JPjJlz7P1bk7CrYTYjEqdQbLMQEKxtge8ikL85tgmzBNh/cGm2svxT5JfAJ
0ZFe4KHwybNn+jTqubopFqrTi9AmB4Jh903Oko8x9CVPoqUcFLi05c2bPd1QRJth
75H8b70NAADg5BVFxBUZrTiHMg5rfdZwLM9WHUUuYEctSxtakkrXaXN86fArEAj/
d6CDpb1EZtzato6rIZkQe0i+/eMRcfijrcmachsiok4wbha178Iyl1rjYILlQUa8
yM9Be1snw+66Dwyo9Q5dWyBMIbt4dUtcoV+5NQdriI4WJHdWGh5MjbkS8TKyzh0s
zqF1ifiJKVc45pVOSL9pKZtjxTLpIbOp+kE6yi1Wp+t6MAo54tkOO/B4viFc1JnK
rcrIgXZFccPnzFbe4lcljNymP2nNryIdRBiXbKpBxGB7vgZvomZpG1bgDrtWAn/r
tJGdVV3EnV5uumNqrRYv6IAl1ZlRd3eam6ok8qbiKFbzb50Qop8U6uwV7raCEvvW
g++hhlv1L/vOshuMJXef+Ox3isHEGukJPPhnj5BPE6mWWhgjy0drRarNhJ7r6DlA
3tQcOo53AkcJ3ZCDgJPJfLvsIMO1BNwH8MymM2PF8vlJqbAGR8cWRani5/SlfGWU
KFUyRykmr3CH/ROqkSrL5guyANXDslYA/QLtzcOKGUFlzPYX+gwNmJZErAKdGNSQ
WeK77WilvixenxuzQOLruQDNXHoFLYe9aoygF7YP2hsaKDqtPqdo0D4rT9mBkJyh
6ezpYqG0ND9bpA8SSbZYdA3aGPC29Hfz+/cWcwQDevjkYpemZ0oj9z8sg6ZShKQb
gN0XpwX5C99k22sdooGOBjEbB9QIiMVb5DKylWNWooQVssarQuQ7lRv4vhQpWACB
aeswRghkOqqMYiqCystwbMjoDGdZNY6BvWdiHioAOVL+qqihVDK7y75g8xSrEs3n
PjC3gam1HtbivO5lHBHgj/SipMVRQ1MPJrMV06uYgMjv9JXfdxrjxmPFxrI4vkiT
AETKbTNFYOAE2R3ViaM40QjfVW1NEKe5s26N0S0sDzS1vlwbLzaXhJFyejmQm77y
whnF4UZ6YsY2nbfQVDFq6/rAy37JWuDQHMSHLr0BiQKPeiR3qRe/hAVk/M36eDy5
NoNyuZN9eSwiPJiyJbQy5fLGYyaOw/2P+F8g98G+YgFpbdwI8kRy6wm5hOZYe0hq
yxjr3wQPgwHatztuWETyy0IrDNxkjbLeucGdTP18RmDvmXDF5ZorOiCIlz870U+H
Aji+sgz0t4nbmK8Aq/NViZqiX43FceVTAorzeQdm9y9Sx1dbER+jkTNxKaFdxhk+
dqtVF4wIYT0P5a8XX+5CsRH3TnV4mQ+twpDZlxgp7QRjKKhs6ROnEHZva992Btwe
3+F/m5P65nV9JjdaMXu41UuoNtiU8MJqzWUEIxQ0SxUIrzVmZUen2Z5GlkG3eg14
FC/Vcs/Te4ff5JcMysp9H0LAU4sUvbwH74zltSFM+xVYZARSF5ZNkQbKaX9xj9ct
9/HiYx88xQA3TOCwxBtx747btltHLwoqHl22mgTTiCuFzCWwbDJ7A8QPOZEjZmop
+pU6p1t8naoOwgVFY1dI8riGM7FFlA1JzAHjeR7n48hDxp2AtjKEcNlNaVOWwqXs
pwZKA80N569ncLOYVI5BEAIcq/4qTgXiZm32n9jBE+bWp83YbtjRreNaQ9vxp9Z0
mxjrugU4oaQUsO6KWysSA/opn5HIJEhWfTetSO12doYxo9aqOq1PELDW3Sj8jRpN
kpjfKG6zVPXxMOrEreMMoO67tgNSP0Sq89BMmkfsWCG3WjYuQJhexWECbBUsTinG
oERcLBubo4teLSA8w4SAjnmjkX3NLEkVim+rsHjY+e0LQWQVu3kt+nZWlYsVpGy4
YqWTEicC5QqPpXSXLW+HcSGk3pbMbBwBB8STcfGat25LvrWHvcTI3IlME1O0ap8p
PmqlO3AZyLvQrwBLlMhanrd/8azsr0Z1AdFPncE6U/fAt19x2k8BuqmSEfrp5xdh
JMuejpqlAFsmNyA2l1/Zf5kxpFzYJsax5msXYOjsWhx5DneXOZLKG5qymIhkYbmA
A0yRLVWKgBpIERzAs4NandwSIS02vJAJgviV59xkOHMpUcdbupCz5r5CbasGytIO
ezCPlpEfTkzKI6wRppbcbFd0zw87Y9lwWswbpt20Q/19LZ2lXcs/RvIiooLCIF0V
n59ZgxqC3Mf0IamKR5xkt+9Uib1wx583GQyCTxTEondh/hqyU28hWqL+klUE3Xp+
G56gQwXmw7/8CIWa8q0Yep5ooj2kVXme1QYcdglg84YQSTly90Iel9fvNSPcKcQW
3JAkVAuWwVQQWl5GMSWGC/N6y61MTDf9b8wcSd8dQwfY+R9SgaX//BRTeGM/0rfA
syw8hKBBbipgXIzBEh+J+lX5wk0P5voJUUdPFaRCfh/oB5gydqZwNwD+Uvm2GqcP
N6m5iUNSNyb8eUJhmEONMFU/sQpdWDyVn6PW7RxRPAMDzxXWws6kukD3u1XdesoB
mr+OlMfJb2yO1Ee8KDM2OvNIPDbkI2ugj8K47i1dJDK70RI5nKhHwDyaX0mQZN3q
s2kkf7cEQkI7AeWNvsGschq6C4mYqII+uA66heOdqDmU7N8zANo3hX52/EgUcR61
m7ezG4zdWy3X+inp4WVwDaRWhGXlB7vy5KPVfouV6Wisz0dUAL+hpiwtLqCQglwV
cZWMlVO4cpi6h0bSMQWMaWH+Myc0svqnSqkq7fAmpIRwIgSHQMSV1YCunT8nTLnq
i0enIc7j7YMN+40FVPX2KU7hOqC1eBCPzqQQATcj4+PM/MiZ13sRZn/zUtKjH9OO
gLkfQpYU54fThwMTzaEnSkxBmIDkE/jt7j2I5S1alb4JXIMdgSAVy/vl4bx+dosm
mOosjef1tklR4jr2/5FoiuMqiyhwPLTAIn1PC5YIigTW+lbdOWagC+9Y7lgkOzCj
OOVajxha9ANua45HUrXyBBDRPk98KunphEuMn0GZ/gSP5kntG+pOgKJG+HUhsAbx
33p2K5A0+E5tgZjj03Tv42usWCkfCuMqhkBH0jV6q3hfkS1Q47QfPg2xI3OzSJJT
0xLC3q+HIehokrlISmUEp/rLHxRLEjoVlfR2RUT2MlJ66TaTCbKXayWv6e4oaUcV
+AOmfuETsTwIzeKpqkVubDLnuPrMi1GUMGNBlJU482lgF4lvtXa2W81lsp6fW8Wx
fMpDcCVYzKsaIfejC8c21jdDQBPXlVWn2kVRS7rOBcxhLEQDogPk6UI5vZefWUhp
ar+l33Q5hcXbUW3rR8MAW2KZNq1P5GN7xaZiX8kEW0LBcNCHZQUU+0sg7PMEzOUC
EIFM1fg5xuGtzy1AF6d0Fr8AuSi6IcirVL4zlAkIWTFv/WsABizkIrxtl+SHSpKx
SuD7zCKjiIfqoUVwNIE+ShzbcQl+GN9BIQhsLu7ZgFxpr+4n3L33C62Yi/UxHGjw
OyZo87+8czFb+6T87jD6thl/dziI7OiKJMXwiQukZufURtNjncj8nxg2ItSpIvJD
Udu4Eu6f4V8n4NLHeSul/qSeYSPvulsCmGj+mt98B6G6OM0AU3+kGR2ObgFeDxvC
FuM7ewt4SAGmPu8mvMHlYz5jaSgMpWx4OJl8Hca8gYtAQH8eu7TCIO1G+kEPg6n9
OujRiVA0cXThzaaH86hhpJniObXE4jCgyCx/mj4Rqca6C2AnRNuFa+NMdwxmOcji
kzvexFcnNClxIn4jbCEaH3ZEEd29wJdoeeVAaUI7KZfx2Q4WCowGoy71z10TYZn1
36xxU5QWgZyjd3naPMHlSLRpKYjD7p4++usAb/MfXEAFatI/59iDKR74W7I9lbu7
nKe3dbKHJBh4oPKcEbJJAkvujNC6I99mT8/dRE7/mH7yKiizfmDcuSI9Llta6Wy1
XIpZIQVB8ogj3lARS80wX484UkCpeLbJrYJY7LFVFpadU0e5rbTQW56PMs1aawPO
BP4x8YRIi1FwRCjdW7sZDrKyYudjcfe6RwahAFqiuK3MFeHNPpQZGVEdCpwSvQe2
WO8aE/HufSRocPHmp8t4N75bswt/R+4LGl/O31YNqotKLCxkJJMDcMVs/Nk9oymS
6eW3h7+ZZrMsxmbWKDQEoJ3o+WuOVA00zq2roOJRydoIswnZJONiOk8BfZ5MA4kb
USmwM1/GwaZgnpRWVW+Qh+E/hLcZwYSJIp1YjNb2OkkrWnY4/Mq8eXjwkQkaEQOH
EF5ba5Hsf1IbVIo3YKt5yrQpg1Fgq+VdAQdzx63lRe4M8dV+WDUvpo2i+YdjBYgO
QHxFB6KybvW/719Pyc/DbN4JQyzGpU1r0y+818J4N5tQ+Q8SLMHeYHM+EcfrkivF
Q0CCxWOZSeVJZzeTa1vYKkvKi0iabxVUwfw39iX8Gi+5odrDMMHY73dVVg4GgUVK
OonzVlC722mBlnWk4Ooa+TisWy+X2h1Qq615mG8Mw39hYrsafKYxWwmmwsWyW6Tv
xYw2qsYqd5ET4ol2ny0red4L/GkvpCOl6gKmnPIx3eVC3lQiOWScdBL4cMo06ZRo
HL53cEXS/iG6QFgyTdF96W3IojvkT4DH4dNVM28nqQAyewdZCvsgFB4zONYWj3XQ
TlhBq+blSlU6WWbXsd+EhFtVBER0SXsCA+DrRaff08DmY/ET9yto+I1Uvg51Plb8
vyelhj3YNZstSJupbDm3zr+EwrSvVQ+aUXaDaaQ1nUT0Z85+PWaq4TEu88/g3XYA
KeDjHAtH6pYHe15Yf5rV/+v0eGBvOu+B5Qt7zi4ZuHrCozteS1gD6Qe+ckKTILzz
QLvrtno6tDxuhBpnqIfsv2WXFGRRIOR3VK6TThhu1mv94BiGmeyAzy1YcxgOksb+
XRhnex+PDTDBjetheGG/5TAFYjEOKFhjTPRtIcNAbZ8aPbstk1eEhCKeFxPclBIy
0Al+i2rDJlx2TdH9528+rv0I8Mxjl4giqZVBnDQ4LTrAg4XNgIWUuQ90XRP2rgaV
uUrksJQDOiEX/rXf57N1Jbl3+jTr7hNWzexsBW5WXJ4d6wFETGvQyB8bEeDifGkW
mRNHrFVDzQpkwWEQcCA0mI1MPT3oUQSr367opF+2pwQuFwNgfs4LAbqhn+lF5p4e
GwPXT0K4jzwZW8xO3dVGhu/TwrHR+477E/+S8JkMrsTepnU3xgbUQn2IoYVQ77jF
4BkXXlcDKSupSRQGXHkDmLk3MBBNwUsWN1nd0Av4bRw0xFNgaR2sS7v5sBaFCEBb
AF/GgTr8Ux3PYWTzp8AqudbzY+UwDX5usn+WjjrhOyHfQj0nnu2edudl8oGxxipD
NcuyP7LyRMkBB/ekg8uKI0seYxZBIsQRTflz/D0JdkSpy1ryFE9rglD2xogza/xa
S3qteXyJ4VhO8/fYjIxkL8/aFYJBzg4ec6H0X/TLKYQqmalnPrhPPAlboQFox+SS
wMtPQWj2OkZIxe2oKBPL0bLC/RdqcSCzA0jDIKvFPUTXKRrMmzCFTMK9X5cNMxcF
9rHgkAK7mmwUjVqGB9AR2j74TmO8kUrS7f38ItOmu/FgGtOf+aDpo4mn5ps5HZwt
Lahen66bvxgO9kq8ZjdH7ExYXAGr4EpmZfaSQGhSK2P340MQMRPWavZn7h1FtILI
Xr/QZ837aG0FPceIgshIp4HuoeaCWVV2CNu2shUD8269TqGrQcrCezMdl3Pl2P/I
aXgAavtbkgYC3DQiS8xdtfPcUWSAgfDwU2GcUHjxxr4ziyvbzxqS/nGsoH9vNtXo
PKaTcy66e+azf8EDE1i/gMxY7yflTgXFFaj3S6JSsIilQSVJVFlTlh9/rKj9nTvu
ovZpnrKP9kevO/HkERECNLNP+v8hZ9cx9qkc3a16W4F88yAvpCPBknekkQ/DuycV
lUAFms+wfhobr9g8edcne4TCL1R41L3J9LgxIApcr2uFuxdLsUvi+PxeZHAJyuKc
PVmP92OLf3/LBHbC+HQN/UvW5XSfD+hPz2QC3wafq+ouvtGfXHp5ssvk52OLV5Kd
J5n5Enlh93P6+H0QfTApIpN4ff7y/3OqBHOalzoAa8oYQNpo8Me9M8fodClzHeAg
7/vhD3MM6dNlQoZAr7hw9VMmwVHnayhb4N33pw6NpsEFIykQ+ZkriDSzvHgGk32O
Aubh3DUq+VmQ9mbwFeeuAb8+vL700Jk3Hd4XH11EHQRFEq4HdsIZavI//p8myGiQ
jOHJCGaQp83RV/Kw4TO8XXBLX/0Jmpuy4+RQygVWdD7jrIUs2V5LM4pcA9o7ThmS
0/UMOd1qzxZ1kZYmzWVm88Wmaqf8Mei74RPd9JQprNoTyHEss5edTpdohuiug0W0
O83kU2fDAeHt35/4T4lEOY/dBCDLRqj4ySnrs/KKaftj/J42O6Ralgy2mR7jmNps
474njy/pyUiHBADne+MaAWa8xJgRmH4NLIiHq+A0NxMop0pAhpgopin9isy4KiMu
NjyfEu7WjsTiecFUFHlkuIpTPUSzfl2buSOOj2nT2iai9yFe3yv6lB465pP0xQP2
5go2VKB/Blu3U/WJPnj1W18jEfo3SrlOVpjU+USRtHurITJHlLncGrR4TomtbrWn
QarP+rhsqVQL1OIH3BsIgaH7KgexeYjs5aiGUMqwpi2/Wjs5PyWaPxXtUZ68vHuB
ypcxzv4Ef8OpdIDuG1EBtP4ZneThSegMKb+UOTAfxe4SI+H1oUrXEDAKAFwqRpcI
SEVq+DcMBLlUTVL8udkOakQ3btGcWeXtqX1hsHV+Zfi+nGAdVj4Gdysd6a2fZi3J
YRh7eBb1kBqkGMXgefwo5osk5nmaGXyVJ2Srjd+QbLEmrfRX2pKRBCwBYlz51x4V
ouPRjnPdN3TXqYMUc8Ep7jzqvEIhBnGcB7et4jEhWru8aabW7loinzHF8fCBL4//
WkvwIoShn7GkPqySHpbU2esLK7lmcnU4Jz9b3H9/IF7OJKSHMH/FHxx//CcCIsAs
QuuJQnHZelUqsXukLUlVmZGknuJFKbbdYP70z3pUWqd5x686iz3uz3e5GUVXmJJC
vpIzDvPf8PuqazUJ9bl0GTl5YiwfSOSiaoRf+LFqkQY9qqUhOclu/6lxC/PtTfko
2FKxjKj814gFLi0MX2KeVTUe+y56jCOYiHpc0Cg25VT/C2+wM8+9v3x+Uxs5I9CV
5+ywzOMR2dumDF0WgKv86zdi7ZPJgLZCEunCiMjLXhRgeBzZSFpBHwdfDhQOVoJA
sX4IbwyrBfR5HcfFBiaVULf5+z0teu04hUdLYICTYCa6P1XVd7wjaw9FFIs2E3PN
jdNpmtpFHwU9A82ItFXFjQ4GzFU9crSePIY7H3dWpPLkvk11TGbqPUd/TPbkz8+M
GVoSc/vNzNRL3qPIwwWH4Lc8hp5NyTB53wlPVMsLS+Zl9UzQVjNvAtSK9Rs3nx09
L8AAGpLqaTaMI50BuK/tbEMPlxLVg5oP3ZrfiOM3WAdvuWvQndABcrMYMq1B2Ckg
grnC+aSExt/pTv+E66qc8N21lJetjzr4Xxm6wWZnCZ41yRwuTpIm3Ltcr28ywC/F
bkDNS51lm+Zxj51XdInRDbQSR/d5l9L9vZNlsYt3Q98X0CWmFA9Ra3f7xgqKF6gB
9eXvaYelGqxVi94EqGNkbId1l0kExxBVVuBqu3BgJk/3iNUkhusL6hMc5daEDi2A
kG+0QqeioUWOdWRDveBSrjbZUma9NZqbLWCQ3EeRHnB6WYguANcg7DukG1QaDCFA
CX8r2ZRbTOkWwrluKa6nIXikJ2ZsX9W3peWxBDJ3pAmOK5/MDvoQHt7rei84Mgjn
Sxj2xeJlhpRQ2D8VM18zCJOFXy8hUcyNY0N9i/0lx6Gt21s91nw6XBS6axJn16i6
l9rpaJjDLbHeXGCspudgT6/EmjE2+osr/dVini/UHFt2M0GJMfNh5XioplgnlaqG
bCtpqKPeRvMaHtWWsUMprYic/ISzvA6jHHPQ1HhrjPYyC3827GGYpdfuysQqj/Pl
2L95sxsjqLEszJ/EXbaHt+DFi9QZote3SSWMSwBJ5369KLNZYU5iOtGoPhTQFPDs
AONncRZQUUQiYUMytOBE5cjOXen+SFqWtRpq+DcfLaa+VzEtwyXJ+xdNpu6RDySf
Nm4dJeEP+eo9sXlJrBX2V+xmIPrVUwaflF4DRmsPBOpO1Wt5Hx88lHJZzsx6rKQm
wTzsDUdHqaLTys+KyB5PGYDrZoTC+MyWgE4ViRGNHll0fupW0XB9vtstmfk7jcq6
tvhR/w1TdqZdGs1OMyha791NiSOM4fZqQ4gqZOskSMFvJJ/VvG5UpIx6R9uCmNT3
mvAnQxaLtq+l8dT20FOPHApQCicEK5era6ddzSjQ5KpklAENS6fYL4iR/HE5xRgt
2vvCpBKQdLjzeIP3Tjin4kf90oBsPefHD41/m95bn6Uj+yt//kchuiyFoQm3uPeA
AXnOcUaKVmWE/MuUFcArsD4TuVJ8fazaErmqqR+H43RcvGCwvJEf4lx2TwfEiow6
TNGoKQIYL6MFBq1Geh1+nDh0wrUlB1DXZULaAisvOHKZ4jJliVs010BBL08cevnp
Cfi/T/FRQbi7NjLRwzfIIPF+HUVdKkXj6amZ/4NYor7gTr9IKLOpbj4eRmeu/rdO
eq3+1w7DvYClUcntaRIbhwsLSwKfjQAiEEFh5wCTKxuiqYIGQW3KCx9yDFP76p4A
6LMbSJlx4h5taicPxMb9r+iGe1hqWAHTNLvGFCT7N8W0Hy1/tVUFIlai7LeZq96G
I9geZWjuamJN8UTrxiNaFAMk7ZXoWVSlkVFJxZbOiUzqnJ4Bn1ut3yrLknuwnJ7S
1z6jIBbsj4IG18ZPSkJrc85zup/YM5KIQYYqcyBoAMA45a1KEq4tUHbM8d5XZW/y
Icy2nDKlN2VEeX28wHeNudR2wn8fm3RWUrY4x7TrxT8t0VIDrDDLo6KS8mGjfm9a
3f4lkN1WCGT+XLHyRK2iyUxAtVKLZTRDmLHnwpZh5wuPZYd5Mr8/HbcoEqTOihsN
kp94O+30f4MAz4KhWjLxlBOidP0RyF1/77AiGceq63BFCRjBL6yocbjRr4kfWtXA
hPloqV8rJvVW4T70BV+EG2Zps3+Dr0eBQHgLFRnd6FJdLYe/DJZL7fBeBAihnQnZ
3Bq0KtPJltmFp+xhiCxFAUo5ynsBTT9oZQ3BZAxlSY/YNoJIEaEaGlgQFZz67Eke
WXWh9GGOl6aJ6ewaSWXfsiFM2N/LiK0mXs6P1TDHcFeqsajjrlBs5ZiWQuis1Bef
xOubo2+QGSGlcOP7jEfhMiyw0aOZ8OHs5YVnYw5+mxGQxVJ6wRVttQfch7H3hTRl
dPw7mnZhSvmluYxe5hSBJze9jF90+BVeHASb/Hk2LPOrRHGS+A0IiWfrqJpXKve0
GwRLqLRXHb3whASIVqd8XUqydwL3Uz9UlgXBJKiMVyxDnpbs6t3sMcFAtH27TS/g
IXcgweEaY8IsEnA+accxkuq/Hr9zJyC2ZMUbaJ+kPFY5O8r8mZwdqCVcZrj2izm9
885R08zyCNH58+RNnsMU8hq8b3cu8PjTEnlsEowqu7rNIGtH8usVD5TvkZBbcbLe
u6KYTGHJgzVh2AHTAKmCeNdjo/hb3rNmU8OAf0a1ZLRMO6VxZ/OdKE+YmJCPY9cB
dNdwW5RurJM64gccnR3L7atHjFdYMbSOBtsfBwEqvWdrqeQ/jjrdJUL+qUZwietv
JkWXZ5g3RAW9AN6SUt1rpNLhZKjw+pVBIAd2OMXlGgznCnnF3O1UDih+o2uEh4B0
qDvOJr0+BZ+zv6oAes0p0PPCm3qAA+doegbhCzfxLzyj3iMHXODT4/DOt1fp1fqc
ojKzgMspyY7xH6AM0gM3amRfBO0f5HaBE4A2tuAGbJKDbNYIM3pO8WjWQmMr8+qD
XgBDjBi2frF0UFEgfUKOyGgVJ7GVHZhwBk5Ymy3TgMeEfKQ8oQ4CHs2DbpAO9QB9
bKZpgJWLyuIbZp6m+J62VYk3PSWUW3Fxb15hIO6xzzh3gZHZci19O9IAK/FfYJBl
fWio1eNeJ7uoeShMMwc4daqtmJLTLJBIWYX3C746h/NaIOPn3ihO1kBJEm45s66j
iYpFyzcW5pyWXSiCaCEC+ufGsid52jIfpcfW+XBKgtWPxfOlm5GoFQsq6ns4uANz
pEn9wIVIyY3yY4vRQwXAQJv1LBPYBzwTsX75/Dsw1S9avNoMg73i0MM8a6RuoTPC
lZIDZwn3jxi39VCszfqplMPxSUM7y9vHT0IF6wbRq+Y/1DFJhHHoI8FtC8CTQpIF
YOVsbLjNxU+yq+Nvl02sJeoiidPbYxN/53n5RLmWSnYhvn8+rYuA6wqew9X4sWXZ
ISmW0rboQKXffPcIiIB5NV1UYQsVWb+8cGOcZqIJ6OpnuL8E+3++dRSk3STHZxBn
+NdgPV8XgUcmPi55cZUuX7Rbo0lWw9E0P3vnKo9Q5orVc7jdEAQOnsG1UQO+TN+B
qLtAB6eGYKISUoC7ljXZgQoWKDE6nTPvAQV6mVh1q3YwMseu3TW15Qm59XhG0J6n
wR1dWoM7GEdz4+9s0pJq2VcqImIV9ZK3bkn+Fn/tuZGobfYgBQBH19M/Owkp7D4+
OlKLUCvSN4+p5VGkkpuIlJ+f8AIJZGa089ysC0tBwZc9MA79u/QvxUGd1UKdXLLL
jPxBhWdGY/yXUeRK1nIAGWCMGnb4emuTZLlFVqZISMIx+8aS9Spg5jhS276ibYzj
B6DdKprVcPIo1+vd9CA6566X1UnL8Lql8XEiAvxGVH4xcOlE5CRd71rtgtN7efBr
OUborPSdbjwBjpJJqED7c0b6d+RtX/gP24TIGpxZop7QdZexWg9YW4cbLw0cyY+u
d6jbEatlJFcS8Oz7OkGO0Vlkkyal3CNII5bXxF/yaysEYIexRle42ahfD9aCIEuA
vqvDBu6fpvdVTr04oL+oVMG9uiEH8xXOjXibwanCZurZGiKx2gB8fV1+XUiDajUz
/iSMRVS1cOJPWeuUwuW126Zk+L7eguV/cOQ3GUPbqINoiCpIhWglR3alBTC0nYhz
f4O2kujOxjLTmyJljIM6oU6ZuC6NjDoRPfSg4h18yNzIII7AgLHvwKw4XNDrLvGu
ZntYYYpmlFymz7mheOr5YJOyqQe1QNzwLI1RJ3/9Q7pbZwDcbPuUiAXRyzNsAhBX
981amFEIkPahzlbJboUGgbco3C/IR41L4PUqNkESwZTh/gOHKLf/BLra8+4S1brr
xey2CouKVx/EgljpoBcz/kQJwpwQvbVfhZ1Ck6By4NT9FHbfkR5voVcL2UoWhGY4
k58pfcoqpH0FBRG7m+xFXwE9c2w/HvnA+5cxk5VrFjel8jDLbmTVK22TwghQ0Isn
9BYWjzbTBq9JI4FmGdc7HoXDUjV25nHU83Jc3hIoej5mTDwK5V5h0x5ghfyOhE/9
ReunmSTIC41tuXqgLrF1BWgaJfQi9fGsq+0f/GL6z+17yhrBQogHPJaZfGy8T5Kb
GjJxIUFetDkBnCPYhubznKAJKV0UhmXA7iIY5we4v6VQoaZ7/K2Illb1mDfRM4Bm
TMDvKhEXR2Sg+LreYwSX5Tg3wRe2ttNuUg1bMtZi9ZWp2XHQOxz4SQ1lIfAJvHd3
niJyNOBYfZxejKkFqOMLMNfnBy7PEGbuIn284bnZJ4Hvba5YZZ3mCWtP40KBsw1H
wKM9dsGIKXcv7DTk2o6nYXkSYfxImNApUTut3u5jNMdbnaKGR8xUtlxQYcp6Z5VB
SDtmPAB1SvosrF6XGR7fYFBDULEXZ5n/ujuPsXqbKwEO0Mjfaq0UDn9+OtHA+2vr
vIk9BUCQ8rakCguO/wkNadxnPKqjUq6brkIBdTb43LHmJUbEFisJxM4kiV0ZhRrH
WM9/h0RMhC558YAgQwaGYlhXccgDMxcFOny8bms5Zmp2sTXGEqQ46R4SHH/E2ima
lTFHK8hf1mX0fL6mHU54lrTJfpS+Mmq5zWO189v3KU1hNwdr04VRSS0h6+RXoY/Z
vO3NTlP+KHsqNPzLYYxZdtIeciQFH4aZSpWy1Ezm/HW0rvFkTup4/UTs+/bUGRfG
w6pJ963Sj1YxAAcsxfY4TOF+4oqEiCf904iUWkiAhTQunvqrW/lQEQ6ApQR02lMV
1vFlZgLRiFSlZ/4qZkbX1FWcFt8ReMH4SmA63pFmCY6rNhvT6Nefr/+l+pdRkvEk
DnZMDxfeon8QQzrhAC5InwS2TL1yd0vQh9rNfnjTbsc6LwkAXdy4z3mXNyYLWhTC
IPCLW0OZcSLz39o2/Js+mDGbgcXrbvS1p2VWxJrI8gl0EXLFtWNtwMVg5/03QzPj
lxuHMkSPRQBnWD1eUDSeYL1FqU3UKq3i4+9w2QGE5F34BOdrRECXrds70ZinAy7C
+88/RqCwSrb0KQGXpAIFUpUcuz0g7xYWpixdl7SY8iJNRJIZ/Zt/uoJttmrZsHoh
hrnAoJl8KHw+dkDm7m/4or/o/iFD/DYTnhYqSMUFry0b8IM3ImTj1FjDIm3ifcEc
meF+Pfzu4GHRUBDS11lnX9CoCTgoapLr8DvYfh08fB71sxzX4YB0cRUs6wFdbfcx
lSknrOdEJCGZiWp2VyZwjXN12orCcsP5YAjY7uEkBctog/DBL5nRUqePLChXflJu
PthFM/ckt3ltv6Ih5Qw+KhOrT0Hun4kuG6lFVO3zgQVa+eSF1qVAK9MV/0NQ2/hN
jiAyYKVxEkoSJlW3ePwNNowPcCKnapkTWGPlmFTQmHbfadt7N9M/iTEqKGhBrCou
qqmElDNlITVOI8k9GfcgxN7P3OT6CdFLKADDsjGUkn9T6jU8N6MnEqQUGHoZ0CWq
KzZE9T3nz3gp05NCI2ZkwGBCM4BBlbfUbKLBnadWEUlwt4UhX7jIsqbAzBh5HBMz
81VfNvJZX0Mal/FHLoRPm71p6YO+XnXaUgC9MGgy9UxN/vU2xRoy9+RHwo2Glg9T
k0G6ZvXgPpX9EGmNRoSiVNyUbS+DSHuVAOkKAaod7jF/12jhB+qbSUgHlq/k2w+i
rtNNbSYJbJO0kGHGnRx5VPRoQV68/fARm6jlgLto66nJwOn8D3gs7yYkeOWDMngT
UOlf3j05TXV0x8aCgrIHUZINBxFV2kNDESF4qKC6etZzUSEbMbsif9aFwoFXKf1j
60JLUhcfumrtfFHsJI2RJlojTRs+eis15Tcotk8b3ULGd+XdhQy9ceI8305OZw+h
CGaZSk7oYHTyuRxy+rCoUUf49mM/l42u64TkZJpxa7qD33EQbWjD4Tf3dDNmZqHM
bTQXodkiWbQS0SMdArnealrU/0ZW1qZo2cTqOCheWrfx3kWjKUi0/xrOdugYEAoe
O6tbprCa7K/A5bov3tVqAJCwfTlpazDj56Ru4/snizOoixScQEH/zx7ujPXx5/UD
ODL7an1MZFB0B0HvTUIeNEdXNHC848/Kz7V44vAAUe3KGHtr62wALDzk9mJwdgK1
YXkGHa9uIbkyCMvSBi/6b4YwhrjAEX2HKoaJaO2SdHIdyz70341KgHK1R3EdLm1q
kUCkeXLVRk8FLuImT/DbX8VyTeffsV5k8dRxJi6UGlMUhdb71RPDJKjgaHsvs1s5
nrbq3sA/5otCfyBTTuFbCmaC674qA5QIfCKFGs8XUDEV63kRMpiQKqx5PhVGs23g
2730TomrxRoCgSk+ltr2E606u305gS8TDeWSbQSPNV+7wEI8x4F179A3duVGTFPz
/3ZrWlA2co82pFpWsD3KEuAQwNelEN4BxR22Kqm9e6TwmZ40dQWX88Xz3p4K0k3P
j7Vo1bZVoH2jmN0oVRk5PC6Eu9GYw7OE0YpE1KPdIqZcAqpednbVaSOEoQYtLbco
Z5wVicCG5E2b1vWWzuIhb+7IuxHqNL4yQf/5Y7gaR7HWL3A3rEOvNXZtFrUzFsUO
9p5HHA/FUxm2VSBSJs9o1rUoIYVwxKToYDnFYXAT+zxoNtHb0BURX9i3OkYfaYEJ
iqQIxYW9J510s9ZU9VMiJ8DbwMwMzPKFgPJHDtJat3rVC67tQJJ+xiFvYmHmu2kQ
MW0vlyyQAe826T+Y9GA+w+hF2T9OOk6/k+haEbjpX803r7eOE5R53NWRsRWgl44/
KnMHU3kBoTXNvLE+sqazDXrWEcvX2rV/jvGvc4kk8yZasvuvrxsP2lRMupgcB+Hc
NY+9fft0VI2U3+uXg2fVQBWvb/HatGHx1Q2zjJDXKGpd1d4SJtL0hyxKnn2XZhmv
GiJT98BnIfnCIgZ02vOAklIasF1UGB0tznMzJdvLSovnr15ROJ7RS4Ij4XQO+X/I
J20hW0zRPql38ca4934uz3IqZuV9vgv6aFZXAAI27ZWgw4x9Bk8pOgcAfjN0JRkZ
trUBc3J9P+wnfVRnrJWDiyg3T/6syHDd2PD0TJSRVjxRkgGaB5R2/R0lJG+RolbS
yluN3S0K0ppxJ4QRYtkoDVsA3tiIrJsIy6X5t83l61+dn62rQ3izgvFBCcXnQ1ob
MjxVQ+8tLQHykC/qOJI0LyCaiKpzV0nfIw0Qq53o2HGKeqBI2TBFAbj1+KTA0dEv
StpGXtRTy8KmNZ16WPA/knZCpX1h5kfDzLAjb6e0AynH2PNXnsPosI/hOdn23S+h
59XzWdcKdqY06abpMTxFDsafexnMubnCr5avWWaY8IotMLCXeFA+GsvTStBWpxWl
4NM5z7BQaZiuFLsP5BrEqQHoEWGh1PconajNqnr7drgSvRk1Dr2D8M7raQ0nPJZI
0jnGaH/EubaG48d3f7NP3BEjaUcqQz7cP3ToVjGmtYZGuurYP3YbeXokCVjZZUnh
M3V1vr5Mw+7BVTRLoas5X2uHe8l9p7cCEMqVTgEAvZazmF2uYCefenkgOPErfQzM
ifHNp0RdMyEwqlPJVllEpjHpCnBnnAdpHUMb//Y/9f+xRtI+7PN+LEf5WHzk+L/U
2XhOOsBqs/dz3QLX2X+7y6eBOvx/coWuVA77eYLUOPDto2/AmGncT7UQnyXNo200
2uaKamYxnPaF3hy4vdMQdRcBK/yFzBkXl3o36gWyP+tRea0HqxUSnK6AJZQU1eNh
RQPOwRwUux2v5z5NlxiT/vAtLQsQBrWed5Dhc3vXbWvUbwNs8g8hssiNKnZDvr/S
lgRifouebBwVPscuShiikPbE2Nbg5fxG/v8U7qDI0FPpB7NJQt9tlhSLUnRDhpf7
Vsv0O9UPaiskGyYjyTVvjiyABhn5dLQNIqZKrDlyQWbTSKuWsnmHFjj1O0dg4Cj/
r5wVkRSqdRY4PI5urgb4FwjThENXaZF0jmjmmoRYmVN2A9uHkc12ptM60dCZ24Vt
g0SL8angEpaY04paZyRVkjVVYetWtBeCwOfR17MpMdvngOJzkar6FYEG5IEWcNa8
FyNXswy+vVBk7Ko3hTqcchwmmmNGC4oYGZXnrE1Bxrv2wfCzffJ0s0wbWJi7AGNj
fUOuBvH5v8Ir8lZnV1Ig0wh+rdrMfWqzSMfDM3EGqWL5Fs2ukwoCTfYfycJrYJP4
FrcH1SOeDs3okDehck0d3bHhWnuLJXZdwFunbRW2bxT51nIS0+AJNZEagD2KgdbE
ATFM9HgoMJP8zuSLRfTWZ+VCKs8En9D2qQP7hkVD0NPpPkgF1CCWQ17lhP7stU5V
vl9xLQ+4OoKEJM8IPPyDDnS9i1tkzzYmJ/eacs+Q+oArG8A/48F4WGi/gmRa0t2q
mFfVHpZg98aNCiPoVUAXBE1TY+xyHButgnQWiWTeZtS6v7AGgCzhiFn4eeDc1cPc
acyk5XVdvduLaEvPa68DVxu7PKq7eyJpc5squ+arqWZlrrICtx5ZiXUO/uuIrbU0
GSy+ZGhJViWLdOhv1pJD/1Cg4mXNjxIzxUrSxv7Kt7MduRQdxaFqhUQH0R5vWFjq
EoHFAwMeP3p1u6csz7tt6owlu6qXhsIPRqCxOIYt1c6N1my480J6otzhvs3HbB3F
ZTH4uOjkfuJELO+EKCEpqagimjeXY7gnnn0hl4l06GTdRv4Zd416ohE9JUiBIWSw
M+2crNRQCfw7tv6RRkb3eatId+RGERNxudl4p2cwRh2z7VKhm57RW9MVmNxlD1ls
2IicfAOKB8+CJ5uNfSg8orldmItewweZKqCU+d/Q81z64wMDNxU5Q4G0VPxpuP+r
YNYFGNFOkJtbvUnQhdObaiUUkuq3jprFKxeonJU/ZrAYQyvlhuMV9GxzN4gKBvbs
OxijvQDT4XULsKIF10aYarA590LWLlmHWgjw00G332w8JPDe85kSiIbrt7FFH/8p
47nMjmZds2325VYE2yMEsz3D1v8nRrrNFBQBbj18Wa8ns1U1kViS3iIeeXRjLN9z
4I9wGzTlwNAUyayN53Rq8O3rmitfgSaadr6XcstEo9mgwgKbodwHVjtpsddSEl4l
DFDfnttR/Jv1aiHwevkpln+InjTycZXTqaHfoG5KxrKjB7I4gO+bZu9EbEswoc0q
XGHwc8ePio3GBMShiEOIguu345uiIllJjHWTXr5LH8q8O4368amvryqulyNYWiOY
OeeellRGpShp9O6D7IV8wLvv42yTuMtz1LwAE78pdQ9MqnPPn3fICAYh11vpPXEa
aTVTzpx/ZzAHQpLjDefYg53ST53M+BCqfqsE2u+SrugVBW7ksA1xuBrVBcduhob/
Q9va6M6xsvjfBixPEge1w0WNUloBOILIUsfFtZTJNzYWU8TZTdYdnf90jn2fvo0/
VzFhi0kcVbijZvjC7rRyTH+moRJ7vZTlwVOKrDJiEfGdbUcP7A6oz53F1y5q67Nb
VhG4dnF5jK+4foDGGNQ0nmA58KBCCWO2D117yt23F59lz59/MjXyhbLlm0oMF9bG
JRtOAwHcFD/c7bl4+Kyu17huYSyEslcQMthAYfgaAWfhrMvDe8PLng9HWnHYYPch
ubBozud2H/11kEuble5A60eJ3yTRMNx5QS19i0/pyaYoHvbNecD7Wtj8g2Sxmcgz
U2h33xjeNvVvLS4PTfWSWal9OzIeHBNUmqZDQSgKLHIFYSXnALwksmoLhaAaSKyU
BsXC8Cdk4+k/Gu/fQFSdH7Gx3Q1WsHDPlV9Azin+9ZH6gnjNPKTV9aJvkLmy3v/H
zUycPvKtk2uMMz35CM7S9IAMmmNS+I5SDXj13AyL2+APdEScGmIkHSJ6FuAK4FGJ
luh4dPt7VVfvcxhONgxrmbgfWDJ9NflJLLt5vtXQexax85YGPJ0Mgm+NBJ57Kphj
7SflPbSQy2LURxuJc2VMLf3uFnm/Wfc1XPu8JUjhWNTidQ008BtoIPuS4olhR4Pl
IP5hAug4USGDH0d0Ik9P/oNrL0T5qJYtxtSpJs2eiYPzKpo3ZTp0qyGt4fSXX5EV
J3DvzjA6eqkp/50A1UAqdgA5DhxkXfvfzuLHgSfEgQRl0qsfXxULC4hLV0b/RvJw
ouVfko42WMTMkRbKKVa4bD27sy1PZRXqANmzQVbsmSfl2Gjgp9V2UYZkbtnMPK9m
QtuWy/e/goRZCXsnkRDrUosONx/cm7prA3nYGvAOISGHwKVPQOWHcSDCAnKexU8j
gOC/wN6TB6AkXcDsqBPUwsdOv9z1vrys7uC0urgPu099GZ+j5j3U7/1/tEb2W4FN
/aM1uVMOtRPdjENqZMhuwxh/Ij3uB14JEhfd/E+4XoOyT2Xp+7+DtHq4zF13Faj/
u9GtjDKDxpbVy1YY/S4gjI2pPSGrxhgX7mnCajRehgjaKVRm2QFaRnoA5LSbctO/
nBLefwS+Ig+RVr8PcXPh4NFx0BwL0oBMz/LEKbPE3EdAptLivtg0CnzzFK/hwUhR
N53+yOL5zDzhGnCxXU4OTLfUL866nbcblXnBo9bB4Id3qW42aFUugtN27su/+uvB
T4ypdtX7siavlwpGT3yK/9npSeV5S5VawaYtdfhviicUOsUC2zj09l89DSuAg4JE
regZbnBdxAOE/5WAkIoG+mNxfYllUvog45sZMRTgB+YyFwOYkkl3y5eOtLeL2UN/
PPqy925LbHM/9i38tqjnwtd6LT8m4jNsO5S429fdOuZyfeN3my6SRyOzKYRbRX4W
iY5O0NMZezzZdTc4O80p7hNIQt0ZDNguR8NUz+zlda4TOLHTO4R/wxobbeTyIibA
Uaf2xvYw7/ruxeayVU9KqOaEjJkdiDGLs4wrjqobsE6F2PUNQgakSj5HP0o/JUYE
9q0nZTwYK5iWRHdS6NUfY6B2MRl8W+Ko4yr+l+56LH4kAAHItEnd8YSRt5bL9uj6
FbfptEx93NxsDRar118moKgJ0ClJQiK9zT+IDAD9Evl8prLQnogfpmElz6kSjK9F
SYCWDtCBbykOQ0LbhKOb4JqeOTswuSuooj42pqY/zBmeM09MVumuVA2iEFhYBbpA
3oByYszmCArp0EWTJ993kNYpTzxU6meyoUPZOqNJpv+WHqh2qz7GdK/7cw/dN4ed
XNUw/HrPisB98LKrbI4L7uHH94sgqseSby9G/Y9brCeErlDnQpQN2w9XXWSlu8+I
83UuiJqXrcH7mVmMkbHsG6SiX9NyahvYST/L4pcmtGU0/58MA5b19gvcT8MNPQSE
lMHT/Wkgfi9jQ4jUC9RNc3DTyfL+Z7JTeRFpC25KgFNHCYd6Mg70GGVIHBNf6/Ks
FRqlM9AwgoFxneDDE/hfytOVF14Nfpr766B8oR/+2no8zp1mqXXpBekI17sDtSAu
5Un/dgAEMi+MKD+LTAajteH3WuXHrfw6xT5Gn5flnHVU0u/8W06FMl7qvIY3tDEP
uv9vSUEOBK7uhp0lls18ByAt4ktPnb/owO/3AzHYxe0V7Q2BcCmxzpHQtdOZTAy3
/lW/1E87gQ2Ujqseg98nSu5PJ7KR4APrETp/bptrUi9beGx66aOXPOYdoIqSKwVG
L9Ic5r/gxDZfpOZirOmf1CexLDNPuDv1inKBzQKY8UDHknFd7R6KIzDH+bM5/zZp
3/NX9WAri6CgXDxvEdS+U+jThWNY0vilbz+54aU1EVPj4fZlZaHs1l+TdTaG2Nbe
dSIvPVcu8DsZNTJbchXroGr22KykQ5yTezBzoYQvYFdqygeWt2nzzOq8Pa2R+03t
oNYmvPjfmQ3srNveO0pKzXWitrAJJXS78KHmQrqL1Dnb/zOZ+pjx3xU6B7JhuN03
1drUN2R5bTDtSVjGeCakjnnPBLCr3IJfNbwRpr5J/7TN1rpbgOvbjQrXuu06jBxv
R7iE8rvVjZF2ykaP4+iiKlXbn871z3wtOa+V24N5nhokSsbHm7QMraSHl/HgItjd
QTBaZ5wVjkXS1rIG30N0syKKzAt0h+jB4DYo8mCsMiNk/F6aavdUU4Lm8MYNBi+4
Icu3F0iV3Lq5ZauVSQ9ZsHIv8JNbwRltgwTTQRr3o0RTvZH4Pxv8PlYUmLxGX5/h
Cu5fDmVh8agOIJYb5C5ovdOmjPPIGn0jjqL/jawnXjgeU97loRV65jLMwr78gT/x
uiA4EKJ0aU2EqrQpAZa4cXCBoHKKmUTv28oJkCMAQLEy2tSGo4QGGKGVACSwu/De
6d2RkGe2n2UYnppk4XQ8v2ipu1nFUkd5tOriszQnXeudf/pNjstZidnYXKIhy0xo
HldiL1EjuYbm0U/IouuzdIvAPhgOWDtEl7JswZuGs53LArcuhwiipqxr66eof0Vs
MmZ+g2yxzj+bd+YWw9ThWMpuX3N28rhwzLCz8fU+v5sAxF2TDOqH1zOHbF+2ln3I
JTGsC1xgComlD6JMvNYlaENDmt3feIBFoSlHHcdOFU6S47rVL4y+B1bmqCHx/JZD
I7PnTwnHWztSx0vkWX++qYqtHkMwC/T3I+fBLkiBGxCmIsTIAX5NlpDf+woD/JQ3
bYkFzxJSMUbb5pvxij9DkqLmLqmcwVIrxq3HcaR+WgD+7y58so6ylSZ/YZrFlkN7
cNwi1Wrze+n6CFOmR0EZ/CgJK+EYeVAeXnzyw7ZK6PbttfkG8HaqO/zGuXzY0yWi
mTTyV2NWYj93/xE2RUJmq85h6pGJHUZAKVhNnWY9S5rF7wKsLz54F/iKriR0/Md4
v48jOfHgOQpqSR/fCezVOaB44x4S1Wdbd3QZ494bV302lKP7d0+ntjZN6KDN/+L9
r7PE9GYLx/aessO1mBCSQmODid9wY66yFkrwgZnGy0Bs0Et3k8aKkhyg4znu0E7e
AkpXMQjwlOvUejfpSKXJ0eEBVPheOvmRvU/3NsCJo0krjFYLR1MD9QUSHWgu0pV6
J1qkfaYb1UPKLgpbS7IJJbbh6JqLDVifRPboCBerjw+QUPTM1vagcyzbl3KQa9tb
zl5Drek0cqm1mnLHCJ8pnnsN3flb0JLhAoGa8GeOiMC56qdF6wmXAerhsSa5pjw/
JnhN+l0hbkyg7/1/hoRfeJZUME4yyOe5kVqxlUOYqdIHPRdMutqh3yzzM49HZvmG
8ZhrUZA5onJywcmrzsP6xPERStAN1UgFni9NTxz5Fn118U8VuggY0xbJx0LtIlh3
livY+bpcFA/L1DXlWVAlzRmquZz8LmBVi6nie6RtjMrt+hpbpGLAxtTlHbaoEimf
IWvef7lPSN3zRkneDquGFIVPe7cJIUU0JK9s0a3aU45xxigkHc5yyBP+l0rOFxzp
0BBLCSLU4DN0ulo4DH1Gsj/d11pl4wKRvu0NOthJt2PNqJjMjKHMP7ZE1wgbQY1f
2tuVFhNCzqs7cqNwiqg0CA3PHMmJ5XXehUGPs/eZ79SHnxzuDNsoTLP/yBT5rLE5
BE6ojiDmZX38wNndZpgchk4HGUtUxO2r5SXHluR2GApFClsAryQQFg35hWzW5b84
agUqZY6E6zTQaL2/QU2SohUv6LZqLWgJqZSz6+X1F0chfmvDIuIu9UbI4a+FBs9m
G4EvxLAWo/JQyDtc1TCQgfvfiCHk0SbhxRqygHv4JwDt7NnNxVVXcC3lSzhGo1M8
MXTG6dn/xYfRfQNkngYUJKM2+P1NqtgF1Q7ZpiJ34n1viwEWtnJ7uWV88LSVebrL
ZQuvXC8SLqgjThf/O59MM/Qe6PBqrTnPVuaH8ph0h3yInQw52SuDK+C1dySD44N3
NNPmH1gaWwVHDEuE6f7oFBmjfsXC6f4AdiDD1qC71JvkzG9BQVN1wOakkHb9IdyI
uLe7sEc6Tph3Nw1PkiTIPZ9rVK8+avri4PHXHyI1nMUs4DwfYdEps/TaRXMkeEwk
9Lt9/TPUa1aXChpjj+kdGkumGAk+OWbnPZcVGxiJ5zHVwG31WgsirwjU2Q8ao0G3
OXBvwbv7rm8qaJC4ihLyZROUczZhGrcv3CU9eJ0UZJcKPzXLRy2PotxhNtBsArr2
3Mp02AUXKWcprkLRice0HTkIcIHpE/lmrrYrSS2ifh67vOoj6mqxf9XbuAWz03aT
6x7u2VAxm2Bm9XF5gMs5tjidYaRotwPo42tpmW2zPlggSxSCyb9uvmcErF4Eb8Bt
PHxNW4nEmrKIjlWco4GuTpAaMWMO4/cClz27tmbriVo8Ka+xSJ3KhB0tl0sXhB88
uZ6ysVa3BMvmjwbkCARlM3Ou/EdovpSqXf70rDcDhS7p22wot+htdJs/tefTEzmX
V41fQGvMK2PIfWxIV9vXq3WE69danPw1OIFJRP6mi8xewnNQqHWdaAgxBTw+Ks6N
InbVHZ7qStndzytzGowFCxlp0W7WUW/ZELMpTlbKb3QXIBnLqGTsm8y62NQ3eCpO
9v2QgT2qGg6UHeFOGYvqaeKfDbtJXr3rFJPIweK8W7aphVuCKiuvzAWSHlqBxWI9
QKZfQLlaefFzK2pwhPKs1t0u8NvnqWBUcGxQ9g4TuNcy+KFVcCtRI5xeo9+qAJW6
XQkOg9gtRMq8mINYSEKtewAltBaP8CCZDm7dpsnRGzjoTsZa/K2uvy4pwU3gI6wy
l3Sdk+bgeMGhhz7qZb30RJKJm0NSXy1x90fMH5hcBhg4nzrNNJUeBNknnXlezsXu
GWR6RQeoxC3guF0ZNOzDGikm8hIB60DoAQWnOePz8PuL4SoeV8LTPXtM5VHjvCDf
F55g/SVEL54T+BibsbS+9Qr8iF0Xq3792OFXdi99W9HhDf/r3zQiAc1q3HxSEZkf
Y7UCoLNjQGlfqlSKUoFh24mYOwKXhAzb2hPJJqOhZwmkCUic2k5w4UO3Z2EUBWNZ
L+uIMkuNw/ZmCDa4oVyWmu9hLE+4m+lVkvtUGYFilaCrVFm2sPU7q4DPiY5K6oJw
qv5Lp37m7B2yTHVz5v9If7j296XTT83EDjI3Ugg4aFENjjTkdKTnppDM74I+F1FF
p0C+CH0vj39gh7lOStqnmUKtWwDsTOYnImGhSighDVRjzeTb8bsKOl9e0q8pIYg+
y2k3ab12IEfQ0HiHvXy8XQYIBrjgvYh8Ygq7ZFlawwKMuPR+8IXfUxqum1G7kfxT
wZpySLLi5ApgjIq58sAfEfLvvzdUupY43jQhcxws+xvEwSHto2Oa5P+DfuTJwUVJ
4FNXVf0Gzx3KlWpp0hzz1vPCnMmDckzH/C2DwHzyFP1JpPAQKaXuD1lMD1nCrVHg
hoQvnw+A/X+HDBLMgIkKpVObo8IiiyTmVskvSwebj65oKf9T5N+GjZ85ogxEXvrg
O5QyASkNIx+qlkQSVWv8bJWftgHK9RGrOgAtFjBGleFcDHIe0UqctuCQP5MmOsgS
XnKB7KtR8vmcL6vTXEmbOzuXNwoc2frAQ/90AUw1pKN5GxtjTNwlyPLK9+c2j8Ia
6YAxB3EkzvkSaaeECEiV5pCIHPDWxtW7nCsXB/MMCKlw/g1JceV3qKLWRp5inAs1
lwG7U9WtGtipj2MtTGqsL3hWzx8HIzoXDVRxgMJxi5VTllcudRcitKCr1eGfPygE
KO2MSfJouMr9tjM/YWV1wKY+GHuxES+oOMgPyj5Tfz+OrapKrOvT6eCc63JKMNIW
t1+opmr2fDoVWTgVqSWDMtIbzEv4+DMactcvJ8FrfQoFw30P/FXZHj8XsmgVLWts
0cBaSy4JjDEqVp1xKRlse3XDATt/Vsf5RZu7sW2niostmM2cd0h8OqH8CYYNmoV/
8d2HSHeSKJPDv7ag538mQIGmvvk0xobx9gc80TS4JZRiI/G6iZAP/OQIYrKqx8i7
Iqgm8sF95/hNc0VDjY4zkc2fQ3XDJfbGEzpShKaeDrb8+Qq3uF0lNmpHSJ4iQHAy
LLHaWvYZeYqzB19r5hq2lIH0DyrW/U2KtCfns4k9VR0MjhgdtnaAZYaZGwvLOWUk
CrWo97DLkbyxSzv4Dsy/10DcrWOKuiVUGQuAnXaEZWP+meIeV8rWBXqrxCT95Bc8
qbdTfWaqqr9JQXOdeqtYc0ULExl28XXF/MroUDCqcpXm5z8mR1bJnExRe0SRIbzw
9M/l5dOKont87yI+rdIxgrLf+j75cY+7f3dkQvcCpLaPpcjELoZd2Y+jUjPsD/a0
3fv+3pSHd7+N3E3+1+g4yGCN1hYruW3STQbn6XCjtQT4Lt3v0N7gqo/sq6JiKmbb
l3leIXPG3br6vuTvL94V6UNd9gbYM4/FpSBc5CoMIrj7mukGLQmrBO+STf3zXJ1n
GnQHsTx9A++moBjiltPqh9bieuHiKzXpECDOkVHprpg+n3x55Frh/ZVPTjYMi1y4
Rz4yaUYy+Jslxko4iV1gkfS/piXB4rteYT2pSAahtipJlnL6gQjfLOek5CoGm+VW
mP/Wb5+MoNux9bbLs1RcpL5hXru55D0/i73dgwQ5KYOBUkSTDIQjtRhPn7Y5ZM40
8ldpfuMYoAwV8vgaKVEjhxJmIAMXOCD+HGhzMBf8VTpE3SHoXLhHYTJLUsZyxJ6l
JSbbhZYAJtRpllbVlQfRtvYfJ0MTGrGnpTKz/pLkkIi3EkjboFBXY3WvrdOwJwmq
tl7H3nAiNcIIJ18+HH4A9CAbn1tNk6bzzofZF/BbDwbtIV7e8c3QjmgpreY0BqXq
/EwSNc+fOZDmfxEGQWmW+oVQMVMu9NqLFL3VEVR2uslxmXJnUX7q+3jZkVhxyMXt
BsdQF85e52whgOKfvu7ll4TRSzsDccWh9U8fdiMOTrng+40GvLVwFp/RH1WWrlQO
I0dIJDpKwwk5DE6VQhXER/HUwOYtQFTBvPqypRFmbfnMItWyeaqrctnD8mckxo+o
zTFk8gu5QccqbaZJp72lpIT8tTcmkYq7DmkJt2aYq8C0bz0x/46U5j6PJ5BZaYkA
SmrOEH3DsWsVlEoNJ+GpOAei9gyR6OS47ePpQHOETIoKp092dxi8up96ITa/6SHj
K7MPj8Oy1ZlAhaw1btnQGndnKntYg9ESbGsZTDKHStp6lcUh0bwgLt0CCtGX/bj2
mQWf1KiqSOom7l+/Kx8h/ZVbcAy9OymPO5riTxuQympHVCKB6WaMxVQAoKppzrUy
4lMbyWgGQCg/inqGEFU6hXNozeVqoFLFbn3mTmZD1PVa39HCSOqdCN9tHcK8CVO4
XeJ/1c+zmKKe0BXGtZhS7YCjTGBkfNgqb093H241vQLovl79co9U5FUbSQ6KBoGd
v+n9HpvNcRxP4cMo4o6G23lg6MuACxXX/T9IGBFZe6eH2TBew349R5KB9glB1n2k
URW4rd2Fzt+CrBkut2a0p4fyRWlg17FlFcDjw7CoNzbkUbSNZ460lblZvGofOm8q
Y44IhI9ECEkjMQZmkeH/Vd1noA53CItEoj0N9w8SzJssvE7X2MH07TovOKPKO3Cv
hSKs81s9+LOE6Budgm6WT1fGZ6wKxVjAHjXQy0EKBU2XgHqR91dlmhIT4KPCZZA/
NrrrDhH/bVS9alQ6OI6U3qeu83ptdBNMF/EaHIC1s99hNOVKvSxBiDYYv1ZDRqBK
ULo9HyyTyxxMDaBafK4/9UV3ZIDhHKnx7B9asG9SZMBpxa54uSKk9oYX0WUw19PX
D0jRZu8p9TQd+O4l8EB/HEZ8VJuZkMDsVLQ1OI+xqEkQmqkAJHWuLiu4JJnyAaKp
Wki/qfM4Ke+TqMUvcwpB7UnYlbPn1eNyHmle6N9+3zzrZkCNT8ZEl7KaZZiJQC52
PTwIPYyOZScJRBACivWbhlvxwZgGvr7zhIj05X3NxAFWzzVZ8jjK8va7LpY1sAxu
w7Ci4r0RRJLTkxRYRpm70L7iKxeoCsBNONJtxS2Wbhw5kQ/oDINHd6m7aM3dIKop
C2Trv5erZZWhSFvAF5g3qJBH0+rOO6YoALibqESdsagTfRDjoeki9Pk/nUmwh0zF
RKmw9oZkxkd+AS7NfjeMW4xZO1ZCdHicjkBeFJ7nVdiNrbD0OdzrW+ouCztZG9HO
obpiLQcewctj3y7Aeee81h6gaiQ1x8AVIE/rFh8Q66Of0p3CR1/XoUnnGivwBo/s
p45cg+WnFEHI0M3uuIlXeuwuk2ieoJrGSrF67F3+8mlq0Zjxblsb7ntawPwQw/H5
eph5m1OZTlRXMPecfgrVv5Sl4tu7DYRspdKrk929ngF8d52rgQIXk7aAsbz3u3Ho
ktOP/btJgoNzdt1x6IXgVdHOPcf/cz1O/VhX3yok8O4IksrogWStsX0SFZfNMKo3
CD/Ih42cBUeoFTDLAmAEJq2W8Mk7ZzlUkLLg2G3awggeCEmyolsIFvkRqhmNUSu7
75FJ2qlY5i28arXHELltQMEV36QOrb9STIAON0xy4AJJwowSYQiQKvrBsxj7fjtm
gHkBV9aVdO2bq2WyO2/rZ90VCzdPU7TSyjMFxT4aYqkSgb0rigoF2icQK9m22UwX
JQjONWPL7aaH88i3r8Z5ED7hfxNXJd7SrH2xCSYGL9xtECnLdyyOWwvxIumYqLrc
R2ww3d65qQIsPxeigctq3xmXF/p/zvxY1Ht3D4ZwE2B11UIL+kiFTb6VgkJiJ50z
N+kexigBoInczWBGzIdBv/yQOQ0GD+z+p8PftQgXGHZTExRjmYyU/po5X/Iry1X0
2vg+kY4EO+qbAeWNioZnmKVB2rcOzaiubGn86EA9lxrXe3xVeaOEFuHxsNFzPoCV
y0SZw+f94wuwMjfhWG4WrC9OAdkEMrHe7EjQSnFHHUNTswwfx8Tl8SQPbHWHh6b6
/FBaJN40cUIpXGZHBX7280Su4Xt0Q3BBO4qvAu6/njHItRxdnWpeGHLlF86JEUUS
4ISDDIrQ48MSCRg5raZBQlyFJVZV/pu4Y+9yCeDWBqdVyj7HxvaRELEyzdwoPw7O
tu4p6B0RFf4wVb9ZPbac0bz9nKLcNX5caMdgWeYh5NCqAuWY2tnckwPeVga7cOLa
91SgTehI0mqKva8PcFJkIsLnwvA+ccbC9/wVGX58fETq4iHsH/VvteFssEnoQJuw
SaSPtrdCKWlZGGQ2HSEbTZAuQMmXEzBOCksmUcDLrsXP0Y/bpKuI2iuTsBjloHn3
mqAG+XcoiMsi/S22SeCUIic/Egm5na0NgglBKqhQcqzM74LtwyFLqNcHFBxA1Yt9
2k4KQMCpOZEfTRZnsFtlD5GT11rV+J2FJ3BNAc1KuC7UCsHRPVP9YQLYZnZ4URY4
j5ljC+FXVAC+tvD/M7Yf39lkzPMDGTyYvNGZCLjtS94PPcqsRxcr/XJ1Yqwic6av
cDhMhg+Ficv7czkokgAMwRX77tgmEOhrJHEbhzWE8hiXD3hL9XpCazsMAH2qniYZ
cv8dis9IkLg687xAdT2fpLdc2QTQrUlscS/DPcIWBxqf57sTBXa5PEMtVcO9W5Xx
dgEfjv3r66DcqJ5X1UY/gj0pxpiYTczhMjSVeU2S1+o+x7U1JMGoKW2zagBCNCbx
Z5lGybmDo+WJalx3VeqJxckLEKywiSsWbW3HjIFIP9Bl6M6/ruVp5fFrdHaJyIrl
NicpuAGBDYroQt8TgSke5GvEQNps9x5WPDnqcJ4F9vSJSyAYIWAedL05GZz6HkwX
cRInLx99aFGH78v5zjBU+Tvd1SNLqciUbfFbyJftx/1kf+9XKYiY76xlzowoCoLt
0Hxgj6d1n1Gwa8iz1AYBpB75+Y4Ru2XQHPw/vrrr5qElAwDq9r9UPQpTkex+Ua58
qR1p1m/00sJRZ7xK9pDGRgufNd2t8fQIcRNemqdRRWEnjbL62jVTFBrsirJk4B2V
pM0iXU1ii9VcwEXz8kGY1wtoNuLjqMege1AvLZIUb8RUN25V7lJTEbsa/i9GJO3J
kXKAJyByBreSJjuBN1aPML0ezfd3IPnltIWrGaFXhgnuluiE/XlMSIXuJybYnWX6
5CTkUp38eUSUaOMOL3zBhtbQ45fSxEZ2jqkoWD1ysuJK9bkpFw+S4vI8tZRiLcb1
k4mpvh5McebZRvovYNA3iFPoZF6kZeE6rQV/bmRvb7WGDHmspRrIre7s55kwLngw
UHP/JQPCtK5iS5+FHXkNjZZg7PVGnYbtDogQmEIQpUmph6Qof+39rKeJKuZbY1PH
JrnYankD7P8aLQxSpr9E9sejTaUMGexsAgRJea82mmFVUu8vaKbCicoLNmY3ZAbQ
tgmDyhnxypLZ8IMTYvGihMVD9Mgxi3uG532zbZgsGJWQUSPL2pZqUWSCU5nZGpLU
mTQfVASw2FJbMqbzMuoweDVZHeud0+0vMpM7hH3wDCcG6ALne9Ck7xiCV7Lr3Le7
5mXTX9sWCuiyludj1pGLmoUMdxJeXEOI499Xq/9nf1Eym/asAEahuZVtVN1r0tyq
t7hiVG2XkeEHRWmPe/lx4q0QepbLKTKReolh2DBGmfL3OHP8oBt5uIP+hVCyXZu+
mTOPb1vr6gJdp9aqhxSIui1TknGbGD49EB27GnOpH6Vt/UHXSwOYXWv7RmwdxMIU
K5XeVSChYIXYYWQcaAceXXjSR3vlPo43eAhmyRN/5/EDizcyCYb+k65GsOEpEaWw
nUgLYa0rOBZuYAFlJqHP5nJ9SPXKYs6e6dcdQ+eD8NgBzAl+w/XLSaAOxEvQqrTI
KemWG6cgg4UaGYw71c31X/17dNOGhD5VvKJE+9gWRnYByq4kMB2UN+yoIhYVUpa3
p3CVS/40YNgpANMD2AiNcugDLAlo2NlGwOw29CcqH0NKIe/8SDwtQRjJ9oaQ61Qb
Xq5RO/GNw8wV5+hpIKvZH7WNixg3ofzAtDtCH1OS0iWLw67YoyukxcOTpL4N9TlM
8Y1oinfvU7spDCp6UFwcUTW2P32PWZSCqHHAt0K41FHzy6cSfRQ4rhWpjToUqn6t
DyJ52+o1GYleyGNZbi65q3iqT9b90vnh2vCrrv3QewaJcccK2w/xV1OIScp8J6Po
+aOlUSvSdb/jMrmH/bYIO44HoLjmg8Qe9zaGdc2P8ksa/dwVkn7t9ApIJtLs6ct3
aKIBcsaIIh1jatYW1C9mk+Ar5be3pA0oDFBEXKPOMlnKualaCcZmjMesPfmzmBKc
thvWc5yp1U5IeLmXQmPKgAn5bMm5VUnLUTn82BKhSw1TJ7NS18ZUjR1GcKGii7BQ
wJggDGmmgRH/pSUn+vl/P3oPO56OD79CGCTA+6yJNqHVjPojYcorO7ZG7zBinzFz
w3RuALjX38Nh5nZh5V2l+HU7pgNFAeDIY3lBloeq2YtD5lM7tBXAPke0PNYzGov5
aeUlWrLwMfMKVpHQZIuB2NO3qAG4p4PfSI8vHCrQDEgmtnU3bO6oN+q1FQkGSz5H
Z/Q7FWSlMVEUdtW1ffn1VAkb18h4R34owx04h0L+7vhhKP9PeIVzyPFWVF5LKQI2
av3tk1GKn3Jx18PEXa+p4cJK6h1zTL7wmNEiUyfWryz8zy5WZEmbfaSQIWQbE/1K
K9xIwOj+Jqxu7+kGZ5eLeUh4PXLQleNY6LQnlOUsRr1shNDboDWue7nHvQAKdlyp
liXhCvqqH/epYD4p+vYT1eWzOdlJS4iqQjzYnAD3T08+OaXGXEUd92G07G0LNJbR
T9FFhhyGXvghmRsgrTEytpsw6zB/RMucaVaflABg+Y7R4TxPYLuHWdnJAMBUVcg2
5jdNj2LJRJNbkzmb9GqY83rbpRff0VFvCVUIyqU0EZBDPyGkChHlGsymge3HrQ6V
SYI1evt3h5I5fdhWzCIvk6N+lg0ZRdK6yfnwLe3XhEIZftOjE+Vyv8Sj+zc+OmuJ
hy9I7AqeYUC5VGrwjNfj6VIqAMmIbriJgF3Xuv13QTSyLn6hH9m/bz9tgefT+N+D
m1C0ijkUmtsZBGvxuIJTi6wrcD8dPPlyJYjWTgT57HI8qy4XWWqRDxIYiBTHE2gv
OqOE9ekhh8xiH9DhwN2QPN8yZvStJRShhVlzd9j/8qAIcCC6o4WnRPWvQNQ3/vNy
Wgl42h8VSUWEZt6lZBwa4FPiJQ+P/gxxHU6vWFRHtmd4+ZWTAPPn5pXbvzizFGwq
RPzYMzMgZkPBk8OPNtqfSXFr33EwezifoYxq9E0J5qzxF0TZSiqvwmHQGv6X1QLD
TafSSo4ZD7OFlFHX0esMeKyt68MVCxYNebMK8cAfj9AH2yVGCfOg0861LKxjNEGa
4Hsq++yNRu2Cohw2cYYpVyaonUqKs1wUZ2Zz0loJgD6MWwm73Yl8QCuRSbkkvSej
BzS70TOBVTSJh3fDtBt5vQU1XhC+jy1+jOrp+VcHglnd1Uf09GydhWeOINL94Y0h
9o7fl+dKC6tSUvadoQuHjNbrso+gOI+Lys/LgUlfj3HM+XojC92lNH4rns/lcICo
QYzHHHt+5KA5mpR87sVZOjvWuZNId6CQSXpIYQBh5jqiNxiegt9So2KzP/csMT/X
jdaEPyS2T4hF2sWQLXrhTo9ZRxPkfbLHu3wM24za+WWSleUicUHKOHfO9ekuNcMv
lHAtQQ731kQXQE+CDWF0pGupaxV73rXg+q8eD70C3yZLs20naERc1YgL5Hh/N8NI
ewongj25HJVduldHyJDNeobF2oIQ53/Dc4YUKXVaEgyfdjE6ZPxDNYM73BSB8clh
j7ZAshLpORdM1ncJoqzsiKVR3DGkyXbb73ZgeCPk8xX/Cjb3xocberSviw2Uv5LT
WrhuWc3JCYIafqb6p04p+hTm8qWY57T0aBWOeolkrBAgrqhtbD/OEuLBTyFIJ4kg
ODxJNX/o4LGUvO2OfIKnlxu4tA/u3e97AwktDoU0r9FpyXQPOuaDTvAE1aInK4D+
vzdzNaOFboQ0jxKVgCs8fKbCJKfsdcdvsrmJS67WpLPrgRbaqAJrE5c90A6tjR6m
Kpl/p7CMAP6C2Ww93/kmYz29MM12y6tuPXW2m/6H/T40aNG4LMFrEgCL0AKedEX5
p7IO20zyW6qb0MYlNiht0tQJYapBzo1G9dSpiwZsW+t0VrmQzAUbC1/j/pump43l
W2pYBp37U1c0Obm5WjWZ0T6MVeyRGVnnL6joHB4mC6s+1YtSDNFxPQ4AwU9Tevwp
FOD547VFSEHRC9WrdSSNHGCgVQqQLugV5eFFLa9TYfS7mzpcgVVukUdAy/FG+5EX
YSbsB0vVNQB0D+69KpPXIfg2AcR4DWywD3ZvgBDL67v/ujPV4JFs44S6ZgExOorf
sCjEBeHhYTJGqiz5eeVqR1k5yhv67OTLiBAutXtKziLnqc966jxoDzEBv969L7JA
6kVXjFSzpAtPuNXz5zOid1iIw11w56/SnNxiM/xre/+kztj7AzEKnmyqWOQPMm0Q
Jl+X1wnA64iSirdgppKnKHI46K3D/gqH5d0Le02tSvOcP4c14rrxr9vqId3LDG27
8tDOMmRH1dYqV3LQg1L3Xae7T8gB1peCEtSA+uP8AiYOk58b22xMzkJ/fNJPZTqW
zAqKWTbv9PlDgHJT14ubXnCS0mQDViISd9RQnF+c3HujccKO0xuuYUbk9JoJPU1J
LxcD9plxLZK6AKE3R13L6L7T4aFqE8hCyXvQxgt0Gp7j2xpKFarGpk/HCQRGk6eZ
+IWuyVPcj4i70JFLOxC2Pd4rvEuXvoqUwx9R3guPMluEyfi6YjwXojDDCmD8qUdU
niZveFI4QwmYCTIQvCcYUIg+ImonQoAUkidHotJc46T+mDcdPMfk1v3+nibHuTTi
WvN38aUgflHNp5K3aiztHBi8bLTyMp1QU0fesu8VZrZBFC9ocmiQMwuzHTkaFIEb
A5BHgTO/dJDSeg2OfpjHJ94mYKxG6vBRaV1ufDsQaFljYcEFH4a6jVbkq462TLCJ
Hvw/6HRy5yFkKgiATUBQOsXw4I87yjoNaf/BOqS4s54pUtt6pSxp4o5DRHm04KkG
ixi0eHAKJtfMtoQR2rDoYe89iyoKOX3ExBiNlK834qMFZXvNunP9dklvlEUyyGnj
EsWyWhh9Xbj6ZVxGQPndi3r5hhNbBkOexepHTaqNJ06ZSo2rusRqcKALoUFyBucr
tuKQM761kdRohaeS8vvADtRcfNuSeCXvuGYVLBgf3C+NRhhi5ZpapXjHe3YZgS4A
OHlwmK0q38JW6NR6AnkbIeyWb11/v8McFdaE7EEiV308Mp5rDn2zR5ypFeqn6QwS
1BvELi8zkau8wn7ZhkW0DaHawVbKBvwd2oxTjl9n0nVRdvfAFGPQJakUD1x5qmr8
jiDDCaTv9Mb7Z9HOxIgAYIjSZua4RPG+HNFXp1zARfsfTktWWXFSCDJRtXyAxah9
QOlNCX6b7y5Zb4AJ8xdy9IYhrCJ1tbLC/stchWuBfCoEle+duaIJIw3pBzKuZS4l
mDfZAizniRrzF3QoekAA4GVPz2UZpI4sXLzloDKXUnZnUDpHvXcCLKV9BV3bi8qc
Ae2Y0p77czqZOHWCFRlsx1kEr6EqtJcByxFZ0CVPW1JP2T4GztNZVJ0WHroMQDF3
xJ5mZ/K9/RWFwXZQ/f5YuxXgXDCs0v6QSpU74oYpBuPh6tkIdKDGc0MnGY1G/YZo
PFPGFP83u4yfzVNZL4LxuVYp9rY6npJdpT+qkw26RTNcVKYbQTEiJuV5hRaUVOHn
Ab8dKNa+N1NpeDTa2AwobxLg9dDtJ/Rw2ArWgy3miPvv3K1dXJrjrPltTjNdHNkk
10x3nGbkffW1zS7PzPpT9g0eqBRyhWiNKMMc3fvjl64ZHLoD7ZnMgITDCU6o/nNj
CCIp4ylmBfS4bL6aEY7Nyi6ey1O3chmiBUM5ddzKkulzxn39PbKMn61RQQmBz6mL
CPJeJeMtDaKSlMhnm+UfyWtpM2+nRS/zjO6GEosYfJzIVikwoJ7zW39998danlOe
Khym7EkSy9QNIBfxvhF3gciKmoHvAzLf8n6Z9LuZoNpp/GmVrq7ZE8ZLOYIJUDhl
uvzPy6P1WmV4gSLLsdBjuxDIis08Q7q1u36ibZp8ZiwCYGh9VUU73x8Opdz473vB
E8pTIIRUhrxsT/DkheWILZCd+NwrofcjaEuNvUkcp5o7hszK3m6YWXDnBY04Nrzv
54gqcd+NhEZrg1A2yLW6nOEHofejqR+CVp+1wvADwyu1S1WbOJhF+yhIt5JX4ZEH
x4PWOnNvixOqVRbOL3d2HEoUqwYJX9j8vWwv4LyVo5QQnHbLys25kkDlmnX6cbh6
9Tgwed2ZzZ5d3KPDuX7i1e8b7smYmn1z8uo9UnA9vEE0z/ulPG1ZuaIK0/J0QrGM
2MHYQ0UXH3jkMeCl7S+PSn3vBwnjl61OsQSDaYTfFTalMdNGPV31rP0K5ffAddKD
foLyebiASVjkxsIkD19Qtd559GIC1tzp5DNPqfgV/Xrou+Rj4jqS6f22F0wziKDh
HLGfDEBwAXp1k7tee7tnKBFUf+tefHhMT9tEMpPZ+EEH4bOfzrFWTagGdRNPcQKu
d1s/3fTsLZ6O+4rVBZVkg51U8Ofi6Eey9GKrIL/uukF+LmiWbQAalVr9pRMGPMqy
gh01DeBOQgqIEb+ocn++nsXnFrPhyfDnHJIUEaysXy2SqjhZF5EkoB0XqBvRJxB4
L6AhuerffHHqMGQUPabzrXW+WX8MhUhRPdfznlChyNIQ2HyKBXPHHhHsXxTwpN7d
cTrUe76YsdnEKM21kpj94mPEeP+fmzKbprgBogh3p0n1yLTUWhAK2P85m+86JyY4
zaDbLcZyinZ7YsNa1xhmFbAggp9MX89xH0SeWyyDi4ZzOLxvwT64ZbwxiZfeqQGF
0ez8+3o7PzjUWFraFVQjQq0VxxT3Q5JTvrsyruAR84u7298z+rhHhlnpdaZqy9K0
Zm9Ej7u1mgYr6f0D5qbQB8S7R2K2VaIsaEmgGYgVLMyzK9LZ/JMAW3MUqQbVcRo0
DG6OzQng4GlyogA+Ouk19kdx0UvCINFV7xEvwNwp8xUFBl+u3ykp/rTjkhlDzbJ6
tJckc5KwFp80N/BurPQDOLk5t1pXGgWf3vZ17+v9s/WaAywKZGr1Hl72bTb/GYMT
j2OLIp7i3MxgWp5yGrV2EAzhLVeyLVffiZKu7Qo5HDuLL0071UNA3NYpPEXGmoLV
vh/RpwgWXkkF0jB1L+rlY4s4dvsSKCSA5TI5VkIZeMFX0irL4IMpXkFT8R6jxMWS
F//IdmN3jr3c+GLCYaYuIrjDXL22ksiBIAjv07DfrMR5qPUBWZC71tlX1WfFZm4U
DlVXkqy2iJbOcqsPKjL2TKVngjWB246AJ90VCB7FCG69vRwYhZ7fnqw3gi1UHWRl
XpYNegTkcBjN14G1OAyOcvTrD2dh2Okinu37DZDXr6uX3uSIm8JPUQhD/gThwpZD
ZDbAiT9ih250hBC623DUrtdr2uJSGgTm917iAqAbXTfyozuKto3qzCkmd9N0tx5X
xsc8T648YrDTzQEEQY2Pt7i+QX0k+QVCPrdlBnGToIrmDUg2Iyx9sMZX95gM/eHg
lzuWGQfNiw3wagUmN2UaAB3WXLPBJR1Sua83/ZDo9qi0WPDi89+k///6IpFPuMeW
TZEJhXHjMBGqosgMn2vOJt9OurBU5P4AwlmdRCM2lkAkTs1yHyZF4DRkAsLp8wOp
OjHz6g2K+a/Lvviqpj7RjLqwcy7Vf+qaG0ZaVAp+OF0M8Uxf4zg29wzf8e8lDZeR
qxk4K151w7JUH0g3/hyWWgL4CzHUKE7KkDISktM1A+vjgbk8C9PBTK9PgnOEYl4o
jhyP4OO1MY9JWyr4dlu2QF66wp2waJPa9VCQrq1SuRj8QA6gL3IIB7+Fpy6vu7JP
SJxWshNJuaWvj1246W5B+0VQKYdaN4s2Fj47tYXd547Qhxhgx4yKJVcDrvO1u2hi
Es8vCaGZ7sZWpgZ1KtOzm6QtAgqP+/0iSvCy/UJKqQxzvqfLsMlTweJboLs1keJG
AU4hx8iwNYy6KLVHtrg3D+EVmOlLeU1fpXpxkObMtJx5XOduuWhg7BSfUSxoqrJH
5q3bn3Sv1LC8BuFVqNfpPOw4ruTk7s96P2s8trpInk/hxL7FjzMz8cldX0pb8VgC
2wMDpQEkBAhfKVwGkW5CGlzzClgL25Ex0kN50hqF6ecSsPBYa63SRpSqLIvF9AMk
gVC20sD9AWLxMJ5NXE67cvr26VB3lGnJfIzOCtBlM2MAOnAa9OtSyxk3tX6db098
Q1yBNS341q9nQ4XypqeehI3q/Y3ex8xPnCwsJUI76+wCcl6siTdEY8sV9IMU3oio
1XJmVv8F6dT64jADflar6gDeSyoW0DTCcSHg4Vv3eZcd8IjaawOrvkZjOvDwNOaZ
QVTVXRDRN0QKWezYhoCwg0WLOHXeDEsr5JqQOF5bQlZhoYSdUv8hIBrkpqjwrPQQ
feWlRaMt21By/VUovsmTObvJkPJpgxp/AXLKFCf+KYGl1/u+/JDWIGt4xhbaU83e
sXUhOpaJLPkid5EL0HstD01FEhLIFnNCtSA18KKkw7AIsO18kDVzxYTQv6krkze4
Y3+cEs0fbvnPuHFxLs2pUPvffLzBXP6JprWuDiy70z9MI/clLc3KAHMVzCIgB9Jg
sqc7f6coY6ZZF3F3iuUypyZ/2mRqwYCDBcZQPQCm2NEOTmwYI7oYe+3+ebbDbY/V
9qPe87eZEjEYaubiyAxaauQvqmVlRvbJQT9HLBm79JC5AAqekFGZY4iphjQCzUv1
Fo6AZteNo0NNG0vKOJRscGKPxW8oM56rwag66ZpEQe/t1vEHeUfHW94qhoylu9In
ZUXcTYX3pA8mTudZF12SxJbH19LS7E0d6fJxF0o+jvdzD8H9eJPZU1h9kqGvKCPc
a3ZxS7t2RXOYQ2S4VIa6QxtKvssAJqEWFK12pQtSRq/hdHTTCom0CYoDa9t2nLRO
ql3JOk382EahTP2X86mpcL9KqH4NQGp7vI+Wu3PDmxB23j5lsGg7b7oMnaInUJ2B
sD/cZ5Ot9B+RgG4EEM4Ubfm5rRilDzuBgNQlhuTaQ6IIDT1nDwvz2mP0o65Cerkr
HX/irPzo4Ug8DzOspY5QATqo1Q9fP7gFV39zS0PZbAxkGGK3x2rJf4EnKsrnItz2
aarg9tQRSLbb+Mmwx5sXkUoJB+HINHCZ0rSwof8l46kU/t8luNM21t3Lqb8gzox5
Mw9Z7V7OQ9XAGCRmDKcWfPm7t8vzhKpVT9OZddGUz+1NF+KvTBLdtftancfacRU+
sYwbs+Xq60Om61AY1jst9nKTKPYU0WGg3tXG/4NqtlAaTUvF/5YbRGjzEOub+kCh
k3ztnWF0kcI6hWUcZgI6DoklzR+n6+lG9DUss3gaWWGgQmKOa/MHlbRF03cSjEKW
BGdzO+R99PNRku7RzZaWBMITRzN1xG6ING0UgLvZoVAeXZj9uhDIW3mMW79TB6Ax
voaETWE8FG3leptMY7DfdJ+ZSuPYuFFzUmehvlfhMP1imAtqphUvEkQhbl1IrN02
Z/2p9jF3gpGFdxGQVFHboJeyG9YcefzTzLMPYJNBsKSnSatHjjMp23biDcvR71F4
qqyyH8b36s7+0610hPK4g5Q8r5wC4Ioc8jBUxePLZUVEUVhVar7f5VnesFpv7gCF
FOkjFG/Hir4DajDqZgYAqVUXzO6482w3M+kBtKk7FvBDWWDekP3lWfCSAE6di4Bb
zMQHdCZhrmvmXNHPXpYZk0MxZhaSTMeVkbJ59znaXlUaNsxPChi7zkuQbrNAIxlp
Mz5M0+odz8BznIfjZ40LOyIxOdaX2X0/J/gIrS5jEv8z01CjCAvHNP1Z6VhQtFEB
ybSWevXkuLKFbMQMEbaJPPCEMqzpzbX61xuCEeqrdD28ZZfb/kVmQGQgIwhhhKI0
i8O3Ml3qkiPLIONy0STogm9PngCjznLKzykFRcJ9NvKH1bFy3pqbUTepqn10yIy2
I3l+2HYJV4cyQ7C75qfiYF2KORx4fLBWLJHy5jt6aO7lDFFY55qz6PMAFQ7UBO26
8viomS03ZzQEtSexrj/FFJGMggIrfY40GwLQ7YfsIM5gT1KVgeZpV0A5tWFS7JKB
pdPzPXmRehBTx5gqSSilgFzcf0e0I05mI6iRKRdMT4BGTu3iGaVq0MAfnbVLPc+m
CkpEcCr03LyL2YgozSnL5Il0+KL/ZUKOF7UJzbQD9iGDGuBdmEWl66gAzFUk3zch
xv07jsnu2OxmQs2tqHyan9z4seCW0/hyfuC3qFAHo+hQFgsT7Iq7xLhIDC7+vylf
z49Z++K05qHLglZY/ivppwYyft62Yk027cJIQESJpQCbL+aMWxw21YQsY9/8sLm4
2da8F1ylm3qKkQVeQ3Fm6UgoxVNbHw0E51JOE/AY4RvOTXaQYeUxy8LsiRp21Pvt
4qjgvZPzetoO8/fJ2AfsaxMq12qF6mA3iSybyWGl9JSlN0tQ7EwLHUrNhH3UO7hz
wc9ryCjmdKhvREGcakEm6BpCFh+Y+9Mv03KNebWRWMt4QpLDjewTkPHyyJdpOFKv
wlZaZlXgHvRaTbiosYMwO/zT3Zi7mEp6O/LF69JvZnllNPzCDblgqjnShOWRjdz4
vnw1fUHWVVmiisBda7Lrx7CRNGuXNOgfOvezFJN8j6d0+3XbIDgBEUxT2a/gW/tk
h+KSb2dPB5Y4a9Y7Qntio0DmPOsPJnmyX4ZD61nQ7El4FtIbsQw6xs3Yyk2Kc/iy
Nn7HnmsgUxal0jRONyy7gbOVhQaCTCQ0s01QDOasZJZ5qpAB0R8o/WKwcWhz3IuM
eONyBDEm/uCDwlLAvbLXwUy8BWS6grpU2nIhegfBbj6atfFLKIccNZCT/QczJLbt
lBziMq79Qwj21uEOqP2NwG8tkZc6iPuhmruDQRe5qhFwLwydwoyLqU8R9eJ0lPL2
GDqo6CiuHr0C3X15OACew3mIBb2R1XeEFR0myc23cgFyZm8ZL1k5R0M3GVvegwg1
SFRKH7Svp19Fysmxc7fcXSff3vCLTaAGBbJ6C2/MJsiaPCKt6ex7SBC8kUAeRRYi
QjLnsOc82MXJImVQxk9JJNF/Q/tbKsvm7HDlRCfomDHXFBdtRG4g9wQKA0nxI5qD
9X05bVn2gCMcwfbPoF8l9dLIx57G6QdOz9U0QHAEVwhof3tgKjGIwB2+SSWgHF6z
cqynFVKeXyJYP2PSrvyZGVyIQ6GPFeH0WeU1as+VyPEyTLyGTmw3XMBeFoJB1CDh
5U72k9oKvGAxxZBuMgjUE3MEcQbDQSdCnJoUe3iuVaH+9Dhh1BNWE1Szr3M0187B
4O7Ty//NXWgCqhiAPnNImkahzcalietYfyrmLFDs9fRPp0XVOEM0XqC3du+NjLxb
mTmoNbJN37RmSLf0EfaboHpyNObIQbhyr2RhkVLnE3pyK8Hy8J4TQ0SY51xQksr5
SgPt9Vg1JZxDn1mOHL/dRVcrqgx+X2/1Yp7JeWMdIiFhd2OJkgdUyQynyFVSh119
ahJkcvNj8L9jbSgF21XYIXyGXd7ZgEpt1eUHWtb0+Y68EtgoHYNIukMnngJZ8EjI
hqIqMPPV2O66XR68DP/zBGx89TZwRl7jQvo0pwwVopf7bc6gFRxuxqq9p7zxiyj3
x192y4kYY9Mw1RNWxD6leXMthzCelR4GFHoja/oyc68i/zTWOOa2CywB+Z5rUeQ3
nNtaxb0LqJSpqyGoOg0IMw4Bm+CakXpGhq7TIrAQHD5VZfXo2PLo8LTb1taKCDom
BY62KS2HNvlhk4d/mQ3/o/0FvAJftKXrBjIW0iCCcJwfQ2eCU2rua6y9Vc6qdia0
yjim9iMcYhEdO2v7/+ARquinm5DCUR7W3Z9qKuRbXmZyiH4HzkdPTHRS+TxNtqIP
i6ZThQIu7sr2KmUl3+nEg40GHPuNM2C/AN8pdW+CcviCHRsD1JBSOu0bdGNIF4l/
MQ8QZWrVsN+9J4/KhcmmPK9kaHfpcAF8vR7LKVp12L0sncrdP3cX7rZCva0ApK1m
bWBNw1GEsHGOVt9lzAhP8XeLBjCjws2vwCasnFpdVhUYhRLZY0kbz7x4ZDgYTuzS
gTMQUnlCsZP/tKgTeEeFm++PEympFz9OGJMx3mCaObLVtiDcZXNCyLOND5z0D27n
y6GoqiGaHaT8W9Cw2sZzfG6e/Oxrbnl7xCgokzXOb4PuH6ve1Sn0v/mvRtzTH7LO
IluYC22JbPhLGX3MRVdGVlg3cnFMy9QGlSl04S7tOu2d8yfBVkSYWXsHVeQk2jyV
lTEG3lV3dEqoWGOAUpkQdvVY/RLhbTWLZ1IYF6c4DDAxKaXeQRv3FLhM46uTxnM6
+B4flwDqUm/P10mzfpdvMq8T0tTHOu4iZScdthu9rQrflU7yfmVrpwaYXHOXtdrb
KhTB89UtqqNCHb7s66X6GHaXCneFcBm1W90VAwLKQTFzaRyhjE09kAintg9aRcDn
GTEO+swL3oJkENH9rm6ePRWICAY2y1FqrbCsaKezUMRWhXqxRYeqRGU/lPU9Cr14
NEN6jo40R0k22Gp/gJidgqTtACtYHRx5YR0tU0R+WY+qbvgJmFp3w0tqL6X/EZ4Y
axK6uYekZUeRes+SEfwy8vKNSPxHy/RC1nu2JHHQzKYbQ7r7e+i6Jl8TBvXvUPlg
2yzPsoPvTJ7oSsyWlNPW/ssj5GXdeEv/pRMTlIEruRcIfjc9qpcQD8ApH436JWqs
/nPbiGQF/Btj36G01qi+zTAVETnz9dm1gbEG9NojvlYci0RFSmI0uCrriNAwheBa
egwUlNbfWLAo49BBRoRoMFWxH1aCjqGokshxoufUMTHONZn+L0iy3JOcbzNavtAe
Y8FWmpuZr1BDAGljiBFntczTrhxawATtQcy/YWBHPELmj4qKN1S7H9omoBlINGcj
xNJRYmd+8mM/Jw2fxrH1ki75J1Xx4/rz1AIgWH/y8bgFiVYLLLeApKynMEREWtct
q6SWV3eTWbrNGH55xGe5UQGax+deffw9cG2Dp9/juHqBSYbWrpQ2XX7UvtXJa/mX
/41CmAPXW1twjVOzTVdZbYAVhOQaYetlfLfU/ipNxxkzCItznxif6YOJA17yP/Hy
n4Wo0kBtY7h6rrDZMxmv/xE2ZXNpYn5UoV2eQ0aulIRevvfAW+j+hX6KW/bhbXlF
Fw9R6Tg5dEcnwyRq6utKn4QteKnBGqeGutR9d53fk9vQOQAC6rliYNTXgJNZYVEr
CV02cfVMIY0dnTI92sEdiKLbFMvNt7z2E4LWI3z8D4kCid5igxs9bdtz09FGCRU+
GNrmxXK6LrSsXJsOpJ+59/tg9QkS7yTy4CzCN6vKmqejLfWy1P3j/JgzfI35ct+1
NLGeWz28FbvoZANnukKgUqlApJmhsxm44LjIPp6kRwSkG2duqvVC1VySBAVwxYvz
hcBrPNYNx7gS2/M1g62NF9OcTIQDmJ/wxW6FT2yV5McYpPR1rNONGaLxHe/Ef0I8
Yqm5ktOTFWCxISmUQkvpM9mrfi4oioY+jYqxbqP03dt11ANfkm4yntXULCOQZZRA
SBuFHMgaLmLy9KfyzRDIqWR0zkrJUj0+gW52butl47qaWS9Ml1IQydLZw4VfBJdE
eWbUzmwh4mXfg58LJd28EL9UgU4wyAf6H5sy+slwYJiDnVdsAz/tHK5lN+yWROXN
XogroIzlQUuyEmyIKAgQntcmQ09jKV+CbuqRNLv67qqWTELuG7UFN9F6mYJkB0S0
uXxhK2aF5CJ031Sf9IU9JM6Eng+mN2ladlPdGyLDQrnfSealVEEV6CCSlcUIklwp
Nfp2tTHAG46iCoj4gTMM1md96iuULCSlGmxUJCdaEVB2l1hBYgVflUKV+XzG03Zh
TQw6ZhvaO0SqxWltgid493+PcaL2HVnj2Hom8o/kaQIc8/9Cgujx0DbP7S/Iudbc
z/SlX0FXXRR8hayGjTJhUqxTTyWQt25FkslL9P/iTEJEZJ/nrqlvb1MqsTR0gqp5
/zSiE0aQ+02+H5FVJXoeYQzirZyzxAC3yZyhiLAr+mBpQXi1a0D3rCG4xbBbaPMs
TqNEWc1kL3/QsuD6IssbkkgVnq5298Ygr9kCoUMYZp9/x5UvPJw62jsNAPisP9bF
sK4G369hcIRPMsYdIYtWoybYYgC/lOoVAWcn5qc6Xdz5UzWJCOMHjg3RIoypFJCR
A8EPFrp2YGlj2t+XLNsbUq+Kj65B9BjKEroLmDwJLyQdw6hVlwNZZ1UNmVcq80oz
VB68dyDZGpj6RZjy7dujMF43HPj/XdX5Y0kVWGMDSfTYVIUs0OjnsSdCcL51fkTh
B0eNZDRFtGuJEG7kUqP9GAPtfDq7yeFUBzarWCoBn+5tLqq34baGQbpu4QEVX5iN
MAMleoY4oR7AHYssKt2/GvGUdlkYU6keeDp+5EhqeLIsuKia0Gl0hX9bIAr1knI1
2a/E3LZp9EiB4FMqv58CcmYEkQvicg3rkn+zaoANo0ARG26HwkO1T85D4zsPBAYU
mRHIypRDtpfVq1e/vk5lAkKaCU1nKjWQ0dsKBsBSLjpuADP3fLbbAItKxi25J8UD
M6RqSsXwEeu57UePiQ5paISczZ46znrH6M0CtUiD0V9KxDrrKO8htaTRZiEwy0gg
CZiGSAkZ6qTt+eeoE+6xlrDCKw+Csnl4A4qegR2UWCs6hoce7YWe3Pzjk3FZo0yW
KUN/ETnecE/xUOXrG79+HpTr0JUIVxMdn/VBCBsqZd3MaA7XapcRbyoYa0NqLyAe
8RxJSZ3jzce9EeL183E0HpwvY31LukPD+468+ELL/nYid3a4vr1hBhhYW7E91Buv
+JpjDPJ+ZbwOJZCbxbn7ZYHhJ1pLBJmcLqSkfKv+h1ljSsb06TrLooLvwbS1Mww/
Ym6KADgYIq21wJzvcC9cudCecv0v7Qs3Js4ltdxaE9/aZAcYfZe0mEGt/rTrKpkJ
6ig7tUuZrcg7CFVcE8cOZJFFE+MsL0u62Uv/yQRrcX39mjkKBe56TlT/SGSPsGjY
J9AEUknf9YydVidsTKMV54q4rn/blAyVdF+Ep831OJGiECoOeaaM7Lb1nq6CFXpK
urd2MVg+RPnDh5UO+u8Y+gAGMMIsHecwmWru3y7JVPEWw2NeX/1deotg6v66ZuxW
MgOKDn8SLVZn8LgIn7nm3S11GuCndD+Hve7RNGzov+pDVlrFPr+zrlw5O/Ej4++g
YTB7Z8VG6daPbxgR+3yQOL+klejj95UxW0Vh4gPJ+SnzJhcpZw6aCJbZofsMM7K+
ZJSgmN+86+6gCpV0gf53IjzAMLHzlCis+lMecTzlBQs/3AHsFt9+xBt59Sw/j6H5
pWqt8hY4PeL7DVhNrZKs0LjATj4if1fNNb3Kz1iYDJPfzQkwDZ2Qq0gOL6W0gpJ9
+X6ZrfOMMNdTzfhlIsmm4uQOEK9hyDOAgLMOTc9esXxWmbh7MMYeHduKdo2Ov0n3
gozRuyxyfsY2JQqATQqQOAzCWAG2m9NpFFqa21YPX3G4h3yQNzc/13xZKemExfdc
4GfD5gAAhwvJV/w/ss2EumVJPtAz91TMQ54Sc1vejcGLhRBCjK1VNI2OOYjIHRxK
ITTK2dKtAn11VIA5i/IVEYT+zZvKF6umZRK2zQRNX1XaaRP4+dZNL7GFXZYplBUX
O/90SWWU08BKovdYz++cSeaItis8n90B/L7uDf45HruawXt+ZBk9CyqEfU2IvHuy
bDTv8YvM2Wa/vsTMtXwfhYLUsPuv2AyPMXdsrzLPoMKZBMrScSGKAXQuOCmof7gZ
xof/BEzmF3KyYkvLnNLbsokzOGbArObl9DaO6NyQlObZvtM/bDn8XYFQdvyH/IHH
tTajWsCLaoSK9ULVSTsSHH2seDRGn4EfwLLIgisdLlvs0tgXHZtggTjev8d59QQ+
kRR6siQ+OhEt22eIJ1+Q/2bp0xoNW2UOPq8r49X8RPIUj783k/RtA3WP0e5LHb67
NW1RBGcrUBSE5uX4grtVzKA00dL6KoposM8FniQJ53n8Zy9JaOVA8zcmMO2OmQkO
mrC8T6t7XrmdvDCm2K82w0KOTEMkInMrhb2r+luKImgZ0SwwvFqWpo8j8SorR9vL
e7hABJGgAiXOkVbTpTng+f0swBcHK4JVc6S/XeD+lOwlN70AiT9RLw119X4X+geQ
3A2QA8g9Tyz7M3lj0pWXzPsI+0p/mpvcQ+nK3Q4Y7cWes4ZUNMfiJsL+ilXvRkya
5kfQBaL4ZPiHifUdSltcg3bw3e+E9CkLNYv1vlRlA6hd/Ead5cUR14h2SzEk4c3M
BsZstnMBrz3aGOJtaBBeQuP2e9cImxeY4YB5GiTrX+rJA/ZsxX/RZZS0lZuMcYuM
WP4NXBQNHlb7fnCEB/G+tqIsTZy2PnLDRFr989pbSffmbP0ZQ/hvddgQMv7XcQUW
i8ncqMq314Jovghwgw00PgNJLrDMCiizg7/GGxjtq6GgSp8vrPZUrKDpXK75b51I
wKLnoXB/5peH0eJdG+o69d9bIfAkZVSeooL9MD9Plm4Jg4CqRG9rbTuFo8sZkg3U
p9JaQ6kLb04gbX+gvtTQ0UOBaw/AXxMUpj0FaArFyzxM5+uQyR+oENUUG9mdCfD8
IOV2H55baAfLrwCmUc2b9AZNSGtiVLR9YCiLsV7VgEdcJTIaWGqkqnbkLe2BvydX
dFmuVeAqB07hDf5VPMDN7zVlEgsq3uhVVgCx0ivQuALtKbsjCCmKRNGGs9lmetQ2
OjI6CunOWUVcWANTgK5/M3pQfuzrT+yABV/XZvkUm+pRrPOcNd/EPj3M8wUAXWtS
uiPcFFRd5WaXvZO3xYc0h9ES++ZwAoUkG+I6GhDGfhTWk85rTEgJ2Hx8j+N7QHCn
f0Kg1aChuPp8FmFclVKijfHLlss4iXyQpCAR7sIGiBPQULle11nattVuMVKstdC0
mYNBexG5nGVFXUSbAndDWfOpliZqwoxWZO/vKyy1mXGXbHqRy/whtu7tr4MvRA6U
VLB/q20h3ip+VXHYMky6DbgBdfpRxgLg4L65RTsEf98oj3y1Ne2/HjqbXPxQVQuw
xVBevSuFRtFNHy4d9Zn65kxT7+6NrxwIgaRqcmvb2+gYHqK35Zu0Hu/zqmTwWNnV
GW3Ps4kyOn7yo7VSlfotBdmZqC0k01vHItycL/6GA1hMCHCWGmI8eMHadXUHpa5W
gcLKNcxH9LAYJZ5hei97ZTiSQ5heDbHWA6u2pOpTeqHKNXBVuO+nuRKMcHkMDKvH
WYwACSZhkBo2ohf5ztGyRsSbdCZ9Up6MpjVjAeSdWp/kkXb9T6eMSyPqzeXBLSrx
kpj4t5g39MqZuhELwLmwWcuOn2SWw/J7dfVV/MF7v98kzF4dU8D50ohITxoQ+1VH
5dX1guvy+GtlS45P0ZdHDd3M4WKHz9dWc+4N2zPRwhvL5PLwWjxgBwd9pd5fcUu3
6mT5I5dpKPfWW0dolCTUN3EuA/qVrEImWdCGpJB/lhU956OuzjtYUO8b6wgvzFUk
MpS80bX0SdG0zB+oYzBLrcu08nUD19+UijZ0xdqlbgQ7viIs23jMbhhHXhXssYCh
2cwvl7qBYN22QjEJStAddOryzei1Mbiv1UJaWsCijQuWnwnDrDbY2ORLOyB0rB5v
YqIpaI+VqADef1N8oftk50+xa/+3zZZGLjKjSWbzhgzzpNQkObIrXfarQiIDdhsy
4CdvHVOkr+UHxuVOKWRrFOauSPPhdQ8Z3AoOuHyTPFM7ws3TSbslizZyELxyseMG
BZRfeaBJ0P0ONDqOVVCpcrocd80KJgb0x+4W+38+fcldB5S5Qh4E8n6Lv4yp1MHE
el9PdAK4TRnF6NSgL1ETbwIBDjdm9dPWa5vqKzAyS0swwyafOliPNk6/t5XGr72R
wNiEKjx9O+OGu8NzO5M2N9zM4N/NGXbMkb+FntS9rUrwqQiN4loB9Ux2oMiYiibN
cklzN45i0i4UrXRiU8vjZ10xOGoeP/HaaMWUYsyBwDdsqBrYwSgH5dUadEElp4ha
STtZ6+9Pwf9SwpPi+wXUqhPru7ZfLxokrPxCC+r7BppI+GegaQ6Hi/3DMqVpMLkz
1nLDmzw4AqDAYy/OPF1+DsFYuTKJspF/O8bArVsbZDswkBXf5c7kXrTgLbCdm8JP
+F+kSddOB262uEhwuPuCeKd5FqFhSLpjLgqfo4NgGnDHpFroLZjZuNSUY2n4cimc
FjdMibgH9Yoa+ao9Cy1gVsWwA8QjTgWWyamFTFGp/XDf4v5Txguigs+2bbcF7tCI
uquh+69Zq9srXq+7Q+d3Hi6q2fCoPvv9A0pZ5wpLjIxp0ZntXX5iBLgO2YFbSwLb
9dchBCqASN3Pf1R3NjJ+P7jQQdJubPvbI9fYX8NuR0WLX2L4Zd3Hwj7HK3s0h6zI
6NweV577P5LCdL5MvOCRXEaMoxqLVkiHyJ9CxJsiNsJlykI2sG0+jwRD5Fs8CXKE
soKbIaJCu1vUIC5rA1LITEMiUN9L5n3VB86Qvp8CAjd5LPcKPgWfh+AGMtP4/9KE
y8aRtADDdIxMWWwzjb98+aEVI2mnDcWwryyKfBG08N9HsccdM5Jz8BqjeAkqKlcP
gm0YmVvk4Uz+gzjTRH3RAZMJcbr5HuLuf5n14kggnSWcq/xP/eGI4awTKzIE+t7N
YcSPEO+C8yGVE4+XXCDpMalqo7i5uoW0unywCRA6qwZ8zfXY7LhSIOlayvIojsGA
ufWqTqdKlLdYyzmWLTnE8Dn2MXDPSK4Pfa3v7D2g1MhIZwIM1N/rEOiE2erO/O8d
4tMQy/inNk7/cPvZ60MJ1AahvpO5l4qHkBQPkYBlHb3ROaxMMOY5Ex7iYOpR3f8V
1LJCCC9CdQNMtkFBYWEboywHTxny7g/HsCaqxUhjNrqCkKWFn+XYw8GpT9SddtRa
m753fAe8aWZsN2WVexSBdlOM4f6cILpRpcTjVTWWsYqXIMw7UfpS8PgdG/s+pyB4
7NU/BywBwEpVvnycEzazVddI6Vtz0zGuCRP6lYefs7+Q5MOKhUvtZJHTCwLN/cZ1
FQw/ekDPfzD1h4TC+NjINuGTzRqpOuGsrtQwWeboHSqN4X8r8vYudS8CRGB/THtG
jRyO92nsmUgtnHYNW0o1b69FSZPaMwSm8rVHr3lsts2t4FHbzxkY29Lkuiwh81nK
siGyG1aEx5otq70+vqRxWoD2ybhWMeo3suYT/v0eOT/qA+0jLd2SInc3VX0CUmi+
+baC55aaBwh8UaO3zkFHu1wTOFV5/RqdcEG7xCxCk+/umK2HvKExAQKzc2d4lkQA
2TJ2oxFTmpFmUoNWD0mqBGpJF+GmwlALUoN3coy40Wfc8IlnStq8L752jaH5dfQT
sKC+5AUGMkjQMXiZDZUB6rCXDpquPyFJ4StLes81Pp/Qtd/N0pHUul7Y8+z6RWDA
r8+v9GbaqFROb6Sl32yQRXVk+bRco4qQTAp9rZzLXwanALc6KzWSmQ/Ciu5MqBp0
Bj68MlGCwx4GfbFtqFp1KuQOSrMUCI1mj/1KppU9ufMo7EvUpd3USoAu4i5BOKUp
8rre4erMs0dYmJ37+NfmOAXAXY8DXq+Cu+7KMUDjolqoc/4/jHgLy0UpJwh3eBTi
lY7e7Z3jH25hhxWinCI9uX79CkkeDfM0oj5waXbAzBnXg1w62D9vjse0SeRviTvK
j9LHJq0Q0qxgGWVY/bpEk+eeT5xgjh8JW6of/l1VBo8DBtGR6q7P+9ilZSsIpOSu
eKsQLpvfHztFebl/DWlclkmTTh2ctbaaDyQOwdtNJp4QwHhsNcn1TdTqfB4fk+5I
QzkYxNBwQPZrj8T8CMjvTko4NCp3kIzrnX0469B6xUwenWUj1T7FUnS60nBPEvzl
Mm8Yg3klcIQZZUIAa7aK8f4HMIHPBVYtROE++k2BP7UwDgOHxPuj0TBaV/ttkShN
r63y0QJaE8rBrHL/0CMNBUi7onaR2pqiD2hwbxFnYE1K/k+BS61xhU2FyirYdIUZ
FfFS6aPWsukwEPDQLEI62bIL4gIcQONoeHM4Jm4nr8mvYskqoGOVznnE4dD/lQ+Q
/7RgC8YStX0fuQ/+nch5wMOnxqUdzrZmlkCMcb/pdfmxY7SUlEehT6wYsQAgokxy
W2QXgMxgD9YMkcK9pwU2gW6miuxjOZcn98xmSEiFAI/xaULrCIKqPf/WLQHtbO5N
c0KG2ama8NOtC2pV1KhuHkbqI2W/oDVqZt6CmCby+LV/5Y1Yx2p0LbMfiwEQFLsj
zT9o8msuwIUAHfMBVo83MH7b5JRvzcquLy4f+LDVzrb/qddB2o+In9qLcllTOzLa
i08tVb630o7ZQpRVWah5Txt3IW5bA6p6EmbsuO1HxPGRPGeXsf5WaoZco27Cn4mi
05Hi2jwBtFEvSQKsOaS9l8/bO+keqYsEP+0PHM7+e6uIAwiDNY4xUX7yDL/fxRLf
Yh39J86asFE8OO4ffvhwTybBRkPja+TQYMw4v4UGtwWowPKcM7rI9qfmryTGFnKj
e0FLR8MTY+NHIH1+d0h5/s/4SJQxlpPGQzl6s+hWT7Cecjg0ud/ZSN9adExoTmIf
UHh2FR7o2yAqWacX8Ql8vsyQiA81z/+1DccIaLoLJXFf3oReZrqC/iMta5aOZ3Qx
mZ0Og3FwhM+ptM+UUHs78wNIDfS+ZzsgsNawnmhyA1LwIxI4dU4wjjsWPa1IrMSp
1IVPHtSIi7g+XHgGJWjXSLSCa7Wck5Y1AyvYjgUkjq+CuOeGLz70aJ2PVvFcsB8S
zfMLPo5nQEJRJiSsH9rjVr8LKS0hfoSbQ2Vy9gfjNkWMTj8QDwA1GKPWmvBWIEta
WNYSXhyxOaSGBZF7Tme9loSKk6GhQQq/GTpsztJraXecLYezn1Jsezx5uiXlzGCK
KPctpxaEQGdNrfOwtmmH1pUUp7B9ZvuTqFyrygr/pJTnvxcY4j1S9h9mQoO8o3+D
lVkpatJjxEnkLTb8OdBaU/kge+qBKzm2NQygxtdEvJOAXECqU3VsGCtygZNvb+Zn
gAv6JXSK07AulwUhe5AaHDtbtt4JuQoT0bzptzZz19T+QQnfpcmBBMFRSYiHuFvi
o4xWXqQ/e4hNCh9VQkKeN/CzElkE2j9Najc8lq/m1C9uO10s0HVTsgVn60WPd+rb
XTf3tdvxinynd6dcxDsuF/aN8VnhT1p9OOAG9Q1okOeyc3XVZOzlx4KSl6f/TD6S
ixHSRph+1q86BhaJgz0zd2TRMkrN2T6kCN7l3j5zg1gzl6jHXf7C6P3yTf1SzerT
yhFZwC67QOc7kzMLTomNoj2eFRNS+k54HxmfyfBzMW/XtI+iXu85S4lNdn36F0fe
li5bq5ktvH0UAOw7YFvSqSWQeIgU+ORe3eTQdl2ACHuDpPzgGYhLwgCjVQTyDc7B
F8lNpvkIyGu9ey6Ky61mq9YH4Ezam3RIT9era6FLQ4d3KALcQAf4xjHd5KRIOSuv
1IaZebLKraWclZu/Ja2jnaCtTBN7lsfgqXStcxf913T7JgDQdsgLuow+P9X21stX
XK3LDHkaf0+LBA8QrtMR0j3ljYZclVEKCHW/ztvTY94et1KluZE5YQCD8Xp48oD+
K6ZbgGQcvB/mNImSNFwZZAQUFn5lVk2ufzZFdOzHI0UB6wu2tt1kk0IVoKJBZdLH
mWLQ440bM4KhB24st9j1LGNZfAVRteQL/Q40t9fge++0wcS3QG3pCrA6D+7ti7Ov
4Romo1SevJVeOCsbfpV+eZMbkXjxvynqX1u4QIpX6bEpgjFP8VcYpj/912faDqIJ
ucnzPr/AY8Xic+mNZKpico00X1dYtJ8DEaN9YX9J0oB+4eay8a5yIglqtbDiShCK
rKfiMg04OLCGRMdsIioDo31o6YUgLsX5zx62wa3ld9g7iBDNFcabD4LFC4da+YQj
3gZXAuIpmgljN57+zAr/KIe3s8BNSb1+5FYbyCAQWcknq+zgwLUDX4mXnkxl+FzZ
E0TZePWblJNjBnbrDiA+2p5uRI5VcDUelLIzf0UTctF6zCNIBU56eLXv2h9aLVJm
cl9bgJ7VLwyDXNtIxWc4ht2A7ad3V15HS6qlz9uIo6KgAFd5p7eRx0PAwyQGA3kD
X84lqDyH3GmqIOola3MfYDXDkqb5oAy59w1cDWUsI4k4UjY3TEB8Lj5BKWBHjFvL
3vY8uUqMlLCCtET5BLrIF+dQbzlz6ZIslFLjkjdLNJPjiqZUVfWy7KYgPUlturae
ns91gEx4mSzDeSDCSttbJGEmNgh7xskz+kLTRQJqHDlNGPrjt7MwtzT/CoEoV5D0
UOm5HcHM+uuEG7Fs1lt25C73dQxioyOpf7wfybK3/p0mrsGNIb1BlcXBxonDPk9k
IV32M3A/mJRYfYQAogSFVylcilOemaxAQtwB/epZRE+q7bOlp7li2tYWI+tXYV2q
Cy7hrzocqvcnMzPTGrrdf2r0Zjz8BKMAYeHQBb2EQd6PusxBKu+nY3eRqP/SXsgY
AJFI0uZeW8lMxRHq8bormBZLnx1aaif8KWg54qo7YAj7fEyG9NNRtVH1BhAE4PJ1
cfQ6qLBsYOlpVnyrSOuCdzSq+4Wv4hRbskGRvyuvC2ahQWHLP2L8pRGxIiL1GYTb
+nUEnoET7gTAOhhJ3g7GZ7MgjupDqK0fvYpQ5zIlxArYLkWmD0bwUVeF1YKuKEtX
MjIIu0jMqiyFJKUn7jX4kQJzlJJGhKlZmhD6o1BItkoCLgR5XrXkbzlyMKDjwyuJ
DtCdUGyp6/noGXBAodv7nKVcSBcujOW7w6BBP/fELaPr2FjyW9N70MxG98k2xWqG
/P5dXCSWJ9R25p9j+gc/70OYueiOyMrXmR1C2dU5jCOSrmu3AqRjj8o1b64pPMB7
zoKsFCFiUkxUthRuXwVlt6ETV7xNl+DvXlakRdMUN7lke9ibJKUMMi5Ks6CqD0hL
zjAUyhluGp1ynWTgS0Yh5xamv7yMD7UKMmT4uOOVg351Y4WI5TYs8mMMSEHA2MKt
mQmn3ha/uztsqskUdEbuIj56KNPqJDJX4w1Qjvz0xaXujJ0XoPzg0mIMXqFV2Pk3
x1HoPcOPJ0FfX3EzmQaE/wi6oE59E2osKREtvg9x8ZgdJZz/6d0qXM2DxulOCFlt
fyPS9PJLJPeMvATCH6MlW7xPEL3hY4G5VwE4HBCVE3yECePG9jSgVoAGKJ8P1yvE
FBaGY+6sE3XBWCWLwizi3lAg+Ku4xv2yJtLObGVzLuvH9BKUR5qLarPJAra0nMkp
BusiSL4/IOUrjes1oDOxL53vrkLWj95EGIcCWuB6A1HAdiePfsV458HrpSTe0fr7
dSx1PGq5+C1OPIRJHJcNAw1gve+GlaUusPaOuZAmVSPudBmzNgZGGd5niuYkwxpX
8a4e+raf12A/g96eZ6Iv+7DMOXZOMbIcNNzvuWbIzDFpfhIc0Wddd+JTfMbxuE24
nzQasrwF0vFoPP6BFP+7cevM5EjFNDFsOt9CB9lrygA0U59Ijm3AgFDmqny8Nl5Z
yvk40sZgWRaazhT0GUhZTaDuYzUgn/XR3yPkcexFEj5lTxq7LaFR3/0jUmGiwSAv
BeQRw/pGF+k9u9F/jv1sdZfLAs6aoNHZBHwvh3193OfPGeG7qa9d7h4aQZuO8G+f
fk2qHE9/YHgcnqTTzTwZvazqXRinLD+T+XIY9xFBU+XL/ECfocMOOqxq3N1067dS
YRUHTffYzOkZbX/7V/tY+CjRXcuKfl+ZC1MAWoMB/PGSfhmQ2vCPd807I/fTlZVP
7tjs8xG4wm+EsMgUsbBIAWeroul+7vW9uFML9n+LLqAyyddeUpMrC4ZLWVcHWCKo
iS5q4Nmtc8RQngKtz/9ItBXZkuOIxtW/mMzkRBZhwgv/nsJkWaBXGz0wFe5KSgil
H3gwrY0YqZAttu8uWlPNCwSsVVKv7IYhEDXgomtHKvX2oiW+J0GNJeUypBN8RqbN
IfQBqqVLCPaeI9fEXJNz9Z4XkrlQ3z5lTNRRLx12MvHTHZsgjv2tubpc7IjJojDa
w9CHLqSibQ0jMnuz4XEPWKS66yrq384QAgSBtv8P5zxunJTEecqnTPB7a+5NHP1F
a/upli8SVsBcNdTI9WagipqZUzuTncJmO+QNQOyAxLkimp129RITlkDelilIegwd
UC22eWElHhzCq2gOlSpU3mL0RvOnrpVACf3s/0o+f3mTR0skigEiBnR6UYX6I5VS
SkKrJkZl18aEOQSFYRHQACDIB8Sfu+4TlK46lO/AkSY8zcGsBQSXBXR3C+2A9I3M
CgVwKjKf8sxd5WNbUqAYQZDmGRohedm0tlrXdaTJXNBbOax0MsYIfR4ffMqGwNa4
mWq+yfYH/0EPu//eusRja781ImS8PaYoJwMCA77aie5FY+QjflDkihAj4sE+8iFi
IS5oGHs5WD51c4LhnO9T8QFACWi1jTLOer5laslZLzTPjg4E+hfRuUf7S5wR/n81
FlN06oVrMd8Ap1yNhSceX++hm4FUS+y67rk8AWlppNI5xjGJM97nEkDPxdEH0Gxp
KtO8Nr1hywacO6bG2MGpdtaDkcjZDb0/5NZUPyb6QIl5fHar1LfRiq50EBm60MIx
QuebEKrJz4xVyYZG75DjNkXLiN1rcAR2qIT4vAFpXXOXqHDlrw13/USP3vZ5dtfI
xo/jLZpMDqW6hA47Jw4u/Jpq/Tx1Gttz66YOGKhEA3xoUYqnjkRA0PU98VC/7d+T
oTPsQE53jY/AWlR9ZkhrKNwRCgzmtym0mS0Z/3Xg4Jg/0UZBn8eBHbVE5lgGxd9F
yhR6RW2+cTyNpLnHBkBjQIx8m0ayUuwFnc5kV43sJBFJjjgtKIGcrslhnjJ1jxWu
FaPZy8V5mzjg1LdzwLJ5qerSj0sOpAd7bRKzWI4Lgrgm+3TygtM9aMbtbz323Bkb
JeydLgDv8YDsj8BFcaVJzqcrSmjJ3VsdFJIXNV2yK7HeNXZKPtm4NW+zt5jX8oiv
6HpcRpsYGNBpXz0U0+Xm2iGztD7JTwBhZHlaMWnxANdRQ4TNFItAsxuzZCgcBhVj
l2H1N6L42wGLLuhEvEiUOU4KJ3KIEpTR1VoGSAaJE8ewDu8fH6bvnKZkYG+Qq1sO
RBEAF1EBr567IWS8EyyJMfX7YZnf4/5knQCNdhuAUSiZFP4pfdvRUaLoPAzggKkt
YEXhFsSpnBH3/1FkBPwV1l0lAbTTGVt3uwh0ClwB9DS5unUWdoKZPnfIWztmxs2t
c9DhRLUxKcmZTPHNwSM8ia3BpDKj/CV1Vmc4j7JzwoP7wqiBIlLtmFDFt/oEn2wZ
jx6QlZk7xfxLkXswPhLfKSsxl2JVnwR6goK/ufWOFZNVp3bLFMTlG6rcmWq01iMv
YJMmO/olU4Q+yLZ4CeUiFKRVky7wWCSNPMS5M3CMGIWSQXVcyikCBJb/fX3iA3Rd
EvlpUyL3Vh6QxGBBvFz7PzH/O+1rR682wAnKzh1FK+0WGVb7MzTYrSPCb2eqxO84
1DNvjWk1G3FYWbaDYGLu8E0gJQBGWQyj2KOSVF6y3m9Ocz/1mA4ZmANxAACwNzPC
ql0bSHin7WRdGdbp3sa7QR16UKMtY3wt+UGmo3P0a5aYoTqOGC1CxvgAF9TLuUXZ
cMtV0IvoZfn+4ybyipBq4zKa8X6TyfovgIC7GnhQR5koe3UcFSx5+mUr3P3aeWS9
ULYIFvSTzlOV8irMcZa1YdBaB3sLQwIQw6NOnelql4cQYUBUStYNGu0KvlT4pSWW
C9MbCGnT2pYfW4SSyMsPrUlew/FyHame7bRun1SGeE6P7XJkSo4qukjwFDx+lkSy
D5JKqI0/aWqLPXWZolhkqhfYshV89Hl7su0G7w3vYMRINUYFh4DH83ex7Z/P08Bz
zsixLQ2uxqIcRGW4q+jDf6axxcbzObU9X9qt9l9yLKxJA0Fw9XcohAv6pAwRnwjJ
RgVQ1yilxuIBtSh4lUZC4gmDzn6BvoTkgUzOp3kuHhzn8pnOJoBZQgqVZMKi22KY
mS9Q06ujR/EPGNlTySnHiZrZ7JL8FXr6rm4Wt7LfJkczpKbjWb8qwjDAjBLl5Gfh
p6ujIFTVSjoYbnyzq2dkBht3z4NGLo35G2zoCzU2NqYwi1WNFMUkUjmPilaVAizR
RaIwhubMCZlxmPV0AE6fNx0LrhsM1bEGgV7NyV1RImNUkJ4STQQ+KXY5YuZEG8A+
KJvh+WyF5mOgLD6BXM0PbdKXuR9DMz1NWD5xOxkq08269pLfz5MtnZvYQP6VQdcl
//yMyYHoYhQquIYTfLRycGmue8ScCDMfcmnuwiVpSzuXIaKj3/o3zAKEEQej3DAG
Ka5NTJt05NtucZ40JEgnMtNo+4ulLRYSu3REJxAmRsN2TNbvRfR8/52ENXuCnG5r
Z//HPuy61Yx6VJNqPaYJIEwme/2Ob6X2KxoFXnEv7KHgj3p/rXKsTLl/1msIYRXS
AaMZdBzIRhBtT4yzSw8YnClg3IhqzAuDzB46Y3OX9guj9iPVBMWVczdKRSwLWYC0
7dJSY0TbfpBuypEMZ6baqf63GRmeP+LSAgOTCr39cfC8eLvjfmxBgJRJya8bQmcB
ccPoedMh+bjWAJpIER40iNRsoVKL6fbg+ECywg5Dh6s92Whhi+1NUOtmdFiI8gPh
BX/GbkXrP/tA6BbtHf3HpPgERRKCMxXCXsSY2H7bl5rs34N0rRsVPnOtU3Llfi+J
CcSiyrBUbl9Wz5hEiwVoJ0xyLjEjBI2IgFIbnXmqwCovjBDe75cSYBuJCJc7CxIA
reJCC1BDAMjEjByzRNE686eIacgJhC8faCXPGvEh7w8WUVVlGzSz35pOPE3hFfLV
YXZ6j7lSdTVgFj5kRD+VZCLkslt6E1Q5NG/P7vUDjri7n+fKjzJYruJCcDfTudv9
focxdO0Mja26hUacbquvM8UgwZC1FuV9e/Nxlc68iZKdScBLEMV9niOSk3S79XYD
ho4SMmOcg2seAWUGr/wwnEkSv03tDZybZS5R2tPVyeg1LOnEbiyC+fkrlKrbFMn9
8t7ZlKcG5rmFaX07gjGfhcL2c2hHJfpzoP/r+9fgcUThyqgQHfHeYPMfT6AOJSuf
0xr/Sp0FOqd/onPmhcewXADbvgEJrR+Dky5jaKIuB/Cx6YwLp/Poj3wH3QThIvYY
G6xdZxzo4mQo+rgWVW5lTjKnnGq0+ec2bnvFi54bZjuQvFeD5d6hLeNkkb8MFmwJ
VbyjGo+AJrjlakhFcMBqLSHrRLDzsS3JR/9aRsylZAalqkl8Flcq5SHCbr2vuppc
RdnnHBSx9OnDelShXdarO2NUc98mvA2WuvxfdztBTmSH5ZfxU9f4t3WaxPSN66y+
cokE0ym40HmEAjCbNMUT3F0mWS4BwEr+9NPvJEjOB8dtCfqreW3OaWRwmbAXNkt+
RC7mriWXiG0Djzrfabrt9FygIX9jxh5cul+/fNr3Nage53unpW+bTlnYQG073UUY
xWkDOtFwynwVvQq2grVDunule23wB3jaurVg0Fy/NGK7sXCTFhmg7EP3XIqVBMEY
dHfpDY9o3picl0Po3R+2HZVY+nSfb1eSfTk/I8/3zmSZkXuZTqg7Cjmi1fXPNoPX
KljPE6Pwifqvz1RFUA8hHRDT3y9PhDC4qeBovvfwsIm/+X01jpOFSqdZimpCPbeX
StTX/ClhhYssrnC/GjPwkAhrfTWDQ0XrBE4jNzUC/MUv9hZIG1ZPz3ZbKFdf4gW8
49JLBfvnFVygeLq5bv9k50bYYqufKeLP+ejw8Q9Q0JTCewp3LXl/Wn658MdCd7UE
X/P1LfDfs1sNoqIo9r0J4BG6yQvbR24+pbl4I9jmfOjD9J/e/qz7hL0UrG5Vn9fs
SrSqsfb7UtxsvjNpvB8ihD2TIEmdhe9ZUBH7fpePoOa34ExQpMBR/HN96FKdDze/
j73KTFK8Kdi4S/bf7cVaxyWK1iJ6ACcnJNEXB4C2ZLQw6zSf70JwiBaFkiTwLvAQ
wb9N4+yvoJUCU2+ZOJ5asg6Y80jWFCvGGwL2Qx5zdbKd+gttKPgcIid6ir/czkut
ufy9TzSD1ugPgd/SBaYpMGZjOw1q/MMzgh6KzVXLK8FtDDmKgKPFBwBXiNSTV0g2
6b9g9SCtc1r2tKFSNgqsilxSG/Xln4O0i3vuhsRtZ11SM+Xx3eRixwHGgE/Fhsfc
TWxK3ne3njYqfYM33+lZeDyPWAfDxxksK5j3on2DbD4FhIjrJGpUZXsLmdPKGh+4
LYoN15AnnPnHCUOHufOqG1b2+IhALwVErbf9aCvUxswtO5Izq6VH8j6p5l1mmRbf
1t44y71l7Z4+vUn6zJc+lDw5kHIggWbKOocGTnf95bHBYTX3/gcGVQDxF/LTCkgo
V7K7BFFtKsgabFZTpkngysx1x4H4w+5ShJ9bUG8uvyTlzGm3YD312KxnJZyijpH6
1DS3SPbDIKQRm4SYqB01jBgwPy2MVY74cCq4MiBz7DC09Hh97sgYwX6filkNiEQf
jmPuKR2ImGFgdlnABHuVTSZzUGKnUGwNx9HDPwqn8qInLUWCaL41t0vafKFUNBTw
ANXvXpF3Q/QzaMWO8ibmhXOV8hA86HVXrNt7YqOS8o+Iq2B5jQILGSwHH7A7tcgg
WxFc04+R5FhqJcAbJ6EFrr60q9+k0bzNrKABz2XjV6ZAJIm+VfPUztu7buJYFMjn
hfT/9qcrKgvvSAN9DUy67up6vHD5BOVKy63Qkpd++3mbbQ1s/dUHPjWQp1wK9HfL
HpuH/xwZGdeMcQKxiLgrKqWkge3DYspcpQximIshsGCbTIxzoaOphjIdc4p0ivH5
d7yABXcLuxoMCWh1uR90LUFPrvCQC8V38THSoafKGo/5Mol5a825MyrKIx/a/Jgx
xnnwm412EcJbgSKn89yHwBxg7eVmqMBEDZqqB0KgL5WiSUjg2lr7AAoIO28QlOj7
PaAjvms7qpoucT1Jj70PpD678yUSzhaZRdag1dWADeA7BsfF/0yJji0dxQ5oC80O
WfPPROkENvZ809xScS03waLiZWMYSJCwfk98GxYlEUCUK4V2aQ9SjqFHo/StTPt+
1NvLIkOsi5I1uXNhAeGnsjVsAfhl2WvtHcaC1JXcgWcAaL/3KDMf44/eWBs0gHMg
cv0x0uxfo9nAsb8/NZmKv1oLoihkDK69wiqL2cX01ved8ESryKiwLdw52LJzqn3e
a8Am7vcYLk9yjMxpI/tnDjt4w4zAw3hQto/Jw0JmvEgc4QDe3tQGtbMKprXnogHD
OqrOUoozHuWc7cahmdsOMaLMWS9UrnBb3DOtzdGDzYKgEXwieh1zT/qJR/70sqev
WnmWWpp5GaNmpgbGA7DNzYdfTAAIh2B8s4h/P1BuAltqUgprlaAnP27xpZ9DzS/h
fzt5DOJt8gDTD9MzbSq7aIc4EIpy5aI09xYT1eiBDXX6Gm+eyA+8SOK1jfMZWWbJ
CxO7q3RgGe2YeDr/opZ+uF+6Js+mk7yAHDLATV8ojPWg9Yp8ZF+Xn5PQietM4/u6
3nK/15M596O4dneB6VfusJMb9Ew2gSsmURMZupYM4dW68TCCuu3uZEKFQiO6jVXg
ZIEEC1XjBVW714t9gGsWH9uGMyi68TSCNqBOPRHAcQcRdFXnJKvmXCaGumik1EoB
4WcoJkO1OVv/FkSXMvKig+e5TV2gmgA1X9qR+noD7BppRiBj5bxz7IN1EcdAopSM
VKcwQ2oLc8Cm9zWtaA3MKUyRDQrI8Ir/Y2RfUZYrA8hUoap/Qz3WfJcWE9oo5Pnh
h8UUrJjFdKj1yE4rffCxu25YX2eP1qV0cHHoZ6wcu1LQcIoLpld5WgqTxvixFyTN
NnjN4C6a7JhjotmtLADVFYcYUGHUgT7ABkXSl7gDaWk4Uep4S+AOdNSjcslzzMuD
fTdP6Z/UMBP5pu/+UnwE86QGUI4jhbinz6RCrq1mPNF4M/6tjTWAHSIuPng5F8t4
JsjXJAVTpfn/0aEqDCAjYtT9scxEEYvN5G1c03Z+ahk6P3dlkFdFZ0kzTyQNYG/X
3OJyGzpx/aolpEh6vztCPkb9aZKa6zK59e3Us6zQE0bCVNgKAEEsGu+0RHTAJIbZ
Z9KKUTw1Lp5jwwiIMvNrfXUypZ55AHfyeDaOztBHy+KAVJ06sy6ooI6JMSZ8p48a
+RrQR6Cv2Hau1CkXwvNTGL/V2nzKcxvb9Eoyg1wZPmdVlGSPoRh4swmlhGevjwAE
UOJPmeopNIJKNMcylIgbXh/9k8ye3IWkrzjiO1K2o0/HKHMCtPNcExrNsdMS6u/y
C1TyMCGsEA6+TRakhjI7cjvrHp9cGdXtW1irI+kkd2GPsC89RKZPKaujIZ32KI+t
3NkjWcp3yRxtPnA5jehJnHMhbWKNXhIsa7OcQilnj3wmXwWCFJiUH05kH1TQL4BE
6sD2X/tRgAOA934XfEESDqaiRFkckMYd2CHEEQ5un9PtZkAy+7pyN4GtFz33c/ZI
q95sIqtFQQptwHFYN7qYvfuYPFRXKWVIAh5c7uNTRlhd0aXxqt2YHzqKbZwmAIsx
RviaoZExXYY56o07Mxtk+pImjxvNvCoW3TUVygYqwTRTLHUWrjtKP6t2ByLu8jWt
3mdB39GS6VUJH77P7LGkSIz6zx2HImve9jOR1gqHCV0xpS9X7LhM1dJ3UevvgjfP
HKmvTNVLBJCV3XosBmK64paz+V+xqCi7PzlzSFgQ+zXHi4cy6r862s8N84rjf6Ks
InQHaf7sDVuLQOc5oNmVUKIqax8XseHMPbI33M/gw004CkM3up8UbptFaLuFiz1g
tAtgvSBtZz/gs1NJxRcIyDR1Ie4DCe/MDAjR0hQrnVhRz/whZRpEqcrQuSSw45Lt
62AphRljbD/Fjg9ZQ7GXq16TZwHTUo/o06u5l+h32BK9GWVBvDjoP7+lNIshP74k
6PKDyDtrU8JXOpg7CyjoMBxUK2i6iv4FYZyGZFR2ejaoz8OA+J6zmU1Wsk5EUj9f
1bubum57nsaKrFBrM1CjdCL7kaCcc1kQW8x1E+/WEnOZPabvOaRA+XzjdudtmgNU
h+3TBrfosRS0MgIU/yQRVF71BTV0eQHNo179sGx0nK2M43M+7S0RUEEwbhscMBGF
q0Gii/j8+PYlzZD92i/Evqpk6svbjAVKKRx/ri7r5sav0S1O6aD2dGcoELGLwyRv
TpilYrTTNoNz+sxT4uwgxrPAnw1y6yOR7QtiGZCB1Fi2EFE0/ucQCjm7Z3xNNnWx
7g3CZsctplFmePlsIDOX1YaxeUfwOB1H7sjCRC7kdUlhTcMcguF8HcCNBEvls/U8
Ckqb3V5qOB6+SZajMRsVaZqcyjCgQAegCVbCnPA+Wk+3zntPrBRmhNryVYaH8J1H
5m3MSAcDoXm9TNDYX1BG0b+Paem/P0A7l3PkIPZQaOo/IF4UYKKKH4P7xZYTsDf3
sdzExjmVp/uIEiqTkNTDKGsu57oUCLyiqquFPqkYEtm/CIElxmC1VSYjb3sqOYks
3IN6IQrYRUi0MElz2ROJRtD0jPKM4O5UG3EqT8qX69TVJFhcAbpGj96eArr+H0RE
9GzyF04YWZaN4+2i0DBbf9RUvokslexLN8NaWxsVyPHsiLIVyTAfoNyfT2SyY5zx
8EcbaSTEWBw2ziRhk+7XLGGy9clRhIKZ/X2p4B2jSZ82pNPxpp2Mz2XbMe29Jxoh
R24PfahDvXEvwmNJzqI1b0TzA2I1rWFqFXFx8sIvXbYV7Rb6bjnenzLa+PIIcfWJ
qKlHJaAhDtpleH3jNhAxBStRCZnVa6XZh5BNW0HWadGji8EZHdAbW6yaNa5or2Yi
EDtFHWw9S76fiNZZGQ2j+aHKHRcUOn15TKzoYBHPkx7Wl6Jgn4XH2e19P+ok35Bd
u5QDEMdGrYgBoWt5mZYYFSWhR0R1Lr8679rWwgO/bV6ZMaeMkyhXGkBybLxBeEuT
YpZkSDAAievwN+PNEGtRL+8aTlLxwFOsNlrlC6/lAL1yHlBxqoocEQjXBb0ege+j
P1zJ65vtzIm0tJTkGHD/TpNedI47erRGoMlf8wQQJArbmXTCamx4i8O7pDNt/LfL
/JhHUeaUcowTex7YJwuJOri9se8fMHb6Zega3WdMMFbcsd1skWWm3Wxki/msSBP3
MKYSPAS/RSNxV7mMo1HwUd13EFI77aNkgZd03rS8CMf5QM0sxk8wo0SZ5e0UuG0e
aFPrT2IKiTVigMB7sln8bePmgeYLdmzRxfDb2r3hykM6nvSdQVgmdrO6J8uzuJd6
R2/M4DWrZHJ3JnqWu/UFPizN0hVlmDsg9xrs5stvD+d1cf40UjTkwiGTaOuOAUll
waSCxwARbXwY5WXeR/AH6qm3o8f6V0EfoBMDDZeDpa6Dbbuuv/nRFiiYF317YDOt
DbaMrPrZgmCk6Cl9ZqSRzmeH/bDWM5l3xu0M6gCxyOeYlKtOSKDO/AkfDOgBeZyy
ymCFXjlrxL9+ZMpMQYwkQL1gI787w/MK4VLB2eZNcihHVgJF0NMTrFmxo7bFAVLW
mLb4iYNvwkNb+FE7fAHAQpRoJE3gwEqn94/BWYd8sWVvFBoMUplJp+oC7vahqVl1
9VfVxymlVqsB3gFITG6yrSAJ9iTNJbxsl0inPAa7ikX9axlyTATOHIyodJ+etckK
TvJ7bMOetMZwB3CdrvABoGTmKVQq/NNcOA4K4KpH40KyT7rFITIY+VUXDtOCiOSw
0p0XnQWxan33fR1l3dgE3MJhfSs0h8Poa6bBKd04lwI3U0bbDhc9i0C4xGl5tfEl
H5gwnMQUycTMFhviUsyanXPojO0X5MRlhnJ87ba9D8IIVl8P6w+Y/m5syByaDvQe
XD0iV+2oE487YdOMKTMEylTiP1vFZOyaWt+M+o0bEsy7msMM73qqMb+PMEHm6xjR
Ribo+7/QH69JZM2p3tBOhgP7ifS6SFJ5KYN2+gQns9GlczHMjNCXYVVbTmL7Fpku
cHwllsMyp5EeajEYv6KYQcpEaGdZzFLuAGn0wJn65sAbBfsSxNsSa7FavuYrPGmE
IB/ioLLA+D5udu6QL5v042d8IpaCgOMXfwTqCEWBnq6mOWljByho+pTO1T7a1PuJ
eOpWSIklZ/Dpf3VlvVgIlYJ+vEno8mVl/DfG5vACf3VAy5s0p3+bXRwJZzLo/e0j
+5hQnt5tflrAsr+deiL1S54/018KvTyIOH4WCF25DgSRixdmEd6TTXYasxEt19Zu
Cn7OnBvULwx2uQ58zMz4uPWCv6uu6UgYei5iNzBxMi6nI8Y+VoV6IFIeTD6zr8NY
HVjcBmh/At3BrtrizXpS9YFyaah3tJBqym362doPop6lNGnWbVxl/4tDZOjeH3wA
vnW/HaW0SlZSCYGEjfNQH0PGq9MsegjjMp/3Sj11wDvJLvHPZzAiTJmAIvol42W/
RwtPempj8E9r88y+QugJ+u14LNLv9xXOgTO+fwNOH4Iw4I/yQcbvVpKmpyLku+RC
j0UgjQqKaXnyG7QW6Vi2YxHuH+eGmcgWXGX+nbnNvlh3u1ZdgaxU6Y0LRsvx+YPP
oZlKldP2lVd5Ioa/o2OQ72ZbS1Yde0h6JiSbjPI+PKS7vPElRsSLR548j4g9rGON
PsYoyA0HXEjiXt/Y20V9Nljxw+Xgd5ZnYreXmLpNUCvBLYs8iFSi7n9F0FEPHtNv
0xmwKoK73fUuDvHSxKntWHnOdToRqHKRJp/gRg95Ce4PdBPW+dFdWx9QxpgKeHTJ
Z8OxO7XVbZ0uwlnnoF1ya6Xv9bd9dmIRu0EdqmbEc57Ho22LL7lz0NFITBr/gMfl
U1bFSfhVYIWpSXARDJmW+g9dtnJR9GupKoS6E+iwyHR005tXYhUgEhhsCuuKQAoi
oPd+4bwjXa0M5m7FpIRRj1IwfwFjmrhG1o0M0ViJSYiTTBaZjudUJgdfFn5mspg5
IQZ25KTm94WoewBmLTbVcCYRUimF1Z7qxzEiF0e3KZEea6SVx2vrX1J1J2GxdCvv
DbnqLOXRJCaihOXnZmg08YUEPmYKmZh96eUQZGCQKP3LRX4QXsBKeQv4udV+ujXr
FWTTI8G0AHT60EWIrB71qNKP+LTDbzhsi6W0gcUITqeI+0z956gwtioxH7L+cg9w
+ycPuncFwoVVAPx6OiwOQMTmBRd8FZqnlz3ycT2iS4HixwNjWrw6mszy/cQcVTR0
VCPOsHr5ECwa03IqPJZduKyghbG1DD9cIgEdT9NXsJSFlhfSaWxowx121a4Lj3yW
C3EaF0iM9UO5oI/ws4vyj1BmOkIzbmLQ0RcuSIdu8JBhN8QWvFSxc0jNJvRoq0Ay
5CPpDJt1JOYhFe+RIVDqwZZ5ea56pjPT/aJvPyP3dPit15aI28WIvZL+tpJ1TV3e
li2APtRhLVLOErzva+49sa+CFNWPGp+J01pcwPXScmr5iZQC8d1+bGVD6jAkFgfk
6A20pVoB4098hHepA+Qb7/wrqRWjnl66YX1cEP+u7uo8FyGL+JUR5p1szAlatrjS
2T+M1QRehyI0E5j8nJfOCNAL05XD/dq7i5RNfOx+06zETKChwNvtFMwnVdDgZv1Q
knqReXRlaKbttM+sKOa1nAVYGpaSUqxzd6v8fFyP5fCuQsV0PR6PB5pM9J7nQEs/
M7kZaNenNEDo7re8OyB2YL2krMuxb9bEoIOMIdHs/sUT7bgW/Gx0ZeA9wXe2sAGg
D/vHPnKsQiXX0Mrqg2weVkM2SwXXzzBDt0uIupz/2Tg92adwexvgp2OPy3oefnPk
wc4Iugfezuw3+66l0fMkdJuPSeQti5IqCigxAUEKoHXRwUH8dZLK9yHLnelpr+9V
BhWbrtUqSl6jyW6MYT/U5JuFdiUv6Gof9tlmIQdkGcNqOuD5pRka0nyGolNkpxXh
OQYI6LDhwg7Ss6l4h2nlA3n1ZzkDRnqHKYFuGHBW8XNDtsgyj3RnepHqngRt0MBD
dcSxEdZA/MJIV6/u16PX7d7+dH0Gf0znPHyz5KauXQAO0gag53wQSCguXtIxw4GS
93wJOiiUxQkHZP0A9jNDYxbsWD6wCHRmm8ApECfKkqpd/ZhJruF9hi6Vzurs2lOM
/2Xa9DRg7BxByVzkpmqMt/rc0F5o6TF51e3rva+LpaHlJegO6Z2zRGxKZ9kRmVq1
3VQQ9+t1cY4xnIREtqF+4PegK7s/XyMQ9Yp/mkIad9dYa1yIp/hrFFpmLUBpknSj
TfL+7TwTveMTxY4gH/s62XiCzN/Lcu98XnBSzmEcP7noy1WRSKD7UUz2R0+/d2t2
vN9oSUltCvALeLjdF7iK2XmqFhzJStOaU8MlMUuk3RxliBoGoJhct9jivJ5vIt+9
NZGKFhHUFJ2hRta6Uou4vwn6R5Zo4mEYqYmjYjj2+JXdZytm0lT/NDay5DWIRzUs
zg+IYeNeF4AZ08d9QhT6O/erI/9KQlXupTyoKvupVmjWY5Ism0Z5WPHOxggt8u7K
uxzgfviEBAWTjn8q0A4CYbYS/Ss3qIdUGd1uNW75J5p0RxJsDOcD+d87cIDt7DAH
3yGbWc/u1DxL9Rm/boP3855fZKFUvlxUe0wWoZhwPsdqKlWYqaj8YL8Mz+W8tf3m
rN2T5wJNy7p5fJsa5+8j+90gsz9N/IZddWa/0yp3k1+oLinck2bE4acbLD06oIzN
V14fBmDUabvVQFsf+A9rk5WirlA43ecur6VKra/WMjUTkPgwtrLUFms+CgVDozFX
OSG2VGBgJXgaHgulSuZ88dwADU1CYCwaC79cpoALNoabo8Quw2vdcPAqpR5P+z9t
hfmMHj/4z2H6GRbQjJm2Nk6XlZVQIrWr819tjlkDjCIjZEQG01qaEN3G/GcAPaSk
zXVfKSZJSBE/SrMt82ncN7bNgLQ6RbCsf9keirqjUnxo6WKm8bzMcUZe4v3Bt491
g19mgegSCxaE2t3VwyFhLfxgx5NpCzHGb5ftbtrWJ9i513LrKrkIZ93/iui+uTVD
tSW+FjWTIc0mieT0ctKL16DGi/WP4jLe/JXeDUnWQQYzLDzaDq8KhE455jO6zIYO
RqSsioVOEm6ppgJcQjSt4SGu1DEx3YPGCKhbhOf1zgljQ8XWbJbO0C7TDjbBgvcy
l/Yp4AlCjCURtNn7XVDn8rI5ufofzINHOsYl+Ij9Wm5zWPNhk6wexg4K8AtoVYle
fP+Mh+wujdmIrxQwzYhgpY3NLNLOR93wd2Wc7dy27NOMQn0ylLklHBerLYbj+paY
BAKYEKLYVrLoMcJqX5HY9vxIyJMt1KRC/VfgjLqrEec5b/AoEyYAo1brovY9bv7a
Ws1P7g/tn6J7USuKLBiqYcKiTBaWEOIJPffaeMphnQK+ijotPtwrQpyQEcot1Lxj
KUb5orh5bvpunXPPvGGP3yRRZYKNBa1JFdR78I3a31m3++OIzW6bM/qt2Rs0uCLI
Xg0eRsxE1De9Qd4LjNiTmrludfCMZCZMH0Z4BnbD7CjVzavKJkqChRlcCIN4cmCN
B6PwNqoeZFmYRFE8ZihkYFA7TWdj/kaDws3oi7o7cWScxdsAWLl5tupbhRWyAVzG
8Zapi03URHO8bTohRj3GyVJOWuOhaPs+iV7Buq3O9JEC0grNMZO5N2zNzWPyW1fU
dUjPyeFtFPtsQwiCPolLBuaFrDexiFmWIObP5sDTaVbnjpwcuLxvT0fGqVrpKsh0
XNEHEhx5XEsKmYWw34GS7unxAvF4G/aRTZW2MSY/t58o3Rs7Bv/1EenBzInLyLDZ
Ofj6Ztv4YKaWAZxvOUE+uDgD8MVZzCjzXpC1zC27v07D6eQ7UYwE0iCSGm7ovu6D
+CpiQKA/ePlQ4GTTe8sLOpyos45V6jBX3El/0fcEuc1ywbM1AfBV/FvkQY6LlgWb
6uwO5n1Ccd/AtqTOe19RHCWgancGE2DR/c4Tw0pvOObTCFS+oogJIVcKM1anz/j1
6j1FSbUwFeof6ZDoibAv85DmjhUZG1gZRICOz3x4Zul4fV4DiFCCYImFuc3FK4EO
zMM8SBvi++Sn/0mduYpdDMi3GVr57zkmF2Se6G0UTic9K4UXYibyiQF1X08kt38N
4bq5mikOseQ3STGClzoWxA8/6TqSg0pGAa5OkGnxlkH821SGuip1z9gBkwu9+lCF
uO5a2k+Cl7UNLI3kh0p2PfM2wrJf7fpBF9BESPJ7kSsNdzg3AUq9lpsQBi70Vnfl
gtj6zX/W2pZ1cT47w+8z5sbH4xz5BFJ9X67TtejUt2dF38Yc63qC0ThT3NJPvEjJ
s16b7kmRkPsV+wK5Vz+qn4r8Ncy7YhBcLez+9C8e6LNHKAcNRIHv4D2HpHJ2jwgJ
xplbrxsqHMndfEk1+in+M+TGoz6BdjzipupWB9jMBVq+iDboJPpEybGZBrfoWbf3
/K55o3cVC3INZTZvxLhqIdYTe/Rss81XBrs88HqgH2irv6kfewlLCIAqSuDbAK29
pNtSKLdxBeEmejUfrpnv48MlHYwZ4vpGIyl/I2+tm5g5x7eZ6Dda9vwJAX7uyGQb
IAL/F3/SOdPTU/usPIXyK6hJCb6ptyFzrCrtqCkgtxGm71dv/TsVxVfQGMREvFzC
UkSWCXP0UC5s+EnRT8/7s5XQTkz12jszKh6h7cwUXTQ8CBOalEOdG39UcKJuzdEK
2Jtk0W8oT0D10pcvsbZcRrE+ifDfHa8QVDxfGOaaYtrZWbrhKJ/acN2RA/fD+jzq
dHlkmCDNiXhVVRj189noGbvc3coD9QtPtSmwM5azNTEjov703F/W2CmbmZI6F8nB
hnRAHpL/QGj7TzRkasmHJhSxk5jdb6NlUHUqSFEFXPKGQurl66vdsF56AOHLWvM1
s/bh8tOrLkTkX/Wa04J5youh11mR5gR5VeI2ZypK2SPTzDKyw9luATcELX5rbMk7
VCzOZbFH3Qmq9w+8BErtESPsGKbkJ6UFfsqX0KYtPZ0VTe5FaJw/ITuhZ16jc/1O
LSJu2eEfpT5KNZ0LSzj2cYve5JA18BeFRrpFGr1d/52ASutbrtC/wQgMbwyowhlc
eeMm6n2wUnx3haR2rvziXe9kMGcbxVPKICtVIb4AEjRxetGP8Bd3BhyfoZaYlZI6
yPH7gr8I9huNasIq77q7uCpBVM8xy/xOx1zgMFjnVoMq9pWujWjr/TcaFgAyB5f3
Jlzma6hsQyi+PWiKCodxRtBkj0CW7m+JyzXl5CFU2qG/YWHvyiJBjnZCbBvf2u0N
JDHQEpq4JnjmWuauGim8B4nB0xo9H3cFHjiwEqVTsQhMHaTsVGXYkG43HR3Pff9w
QLlVimUov6T7x3KcQzF1MKxpkyzx9f0KfT4oK20CMeu/p2aWTlHOPF9uzwrb5G+t
tW+PyXLca4mCw7s2HmwPXUckq752DT19w7S7mIaYBV/cVCIcC1scvK/BtWW9KPtC
fYiDeBJECP0yTEHoKC2m1EcvsLC78OVJn+f5msFKOBbr0C8jfQ6CqTx3W6tnSSVJ
tKLJECP61H77onREHVnze5toL+W6+DHZ4uAcMlcQKMUJjMH7LwXTa1ZtphsBowDs
POu5MYo2fHftfiuJVnIxckJzDIJcV5ew8oRdDpeTCrE60ZZUZaRQgx3bLp7Q2Fga
5QUqXxAi79SecQ0SgiA9SzbzR84kPXVCLolQvepHcofbq63WTLO+NkY8lFa4HF8G
ClwveXTDUslTBaxaJPdnY/ciZwVosANRiE3q3z5/+1ycOlwbtHVOF3+a2I1RWpDe
HVqCOoBveZhf6VQFb3mgbdIfK+fvqmEhgk1rbUxhYEsb8EDXBkL4l3eUY5irxXrO
9cmr8Weflu8xphATTVl6N/DLovftfg6ywFqgG15FJHOEhuKwbzmsJgPGD5S7LQrc
UssW6PHLJ0MPrO0EZ+FMBIZm07AY0WcW0LRhyOfkpE8oP1MamTasdyOqQf74eETT
hzeXgCbdt6HuWdSXkIkLah5G1skT2OrEa/uws2s3eNMR0XGgQgWsVTkNCZMSheqF
boAFZsA+p8PvQgp9iGS3YLXdhipgS6QzuZnfeGEV1j4H9jA+iud77gTcuaOCEa5i
3nr1DnR8VTHnlTK8tFG9EMVRVR5yvuZU36IGglMPREqW/eZc3Di/eMPqB+bFTSYC
tvtouxA7LfxJXccETNaSTuSAN6zHe3X8bJG3VWsA06hELGilAdnjE7uvJ1nn3fOy
iyUpNVQUXYejhqb4TuL/9ghYT+IRFkg9JVlDO4OYrErnF/vFH0dR9YA2Ols1GMBB
FO8JTkiYB7WlcnqGeO6CCk5zZjdybV70wSSb1P8fD/or/xkJAWmgr/Ph9ayDnwJg
y2qJOi0Tl2tv73LGu8FRlj8YspZQA9hB43Q5uVvCNr6GEGJLirDw6eMOOWsO2kWl
m8OBECXkZOhbPo4YdDA87Qjbz78TNl57EVqbAJd9gDruElZ2Rdd0/YsYIWkeuq5P
xB0wwOjtyh8qaXnjRz0DNhytvW8PqCJ2xmFjdFQlRmO4W8kqkuQCEZTETFYTWTZ1
orqES1jIzr3tG66WQbTsdlYiyoedh6/VM2in3nMECsgkPhrN7SYFwuEobquj0I80
3Q6cR6q0QIkPDOdjTerPS38luHi47658chlhjL1BlD15bkwF8mmoIyCROL8LQm69
QAfIMpWDvJrSUdbFMiUU0+VWHL59qsmQhR4sj1P2zo1IRnou3LdKupGrJESovuey
fjRGt7flCH8zBvSYg2qZl3QmGYAsbv5Ysnum9dsneDo3hX1td4lVJSEFWBSRkIZk
cuNNRlTm4hhCQtl3A3diPV5ArZP6iBLWZhOr6uC2m/rv7GlqGmWp+QjDPAWi/sEp
NETRVOYc2Tg4phkJ+y8UjoJKW6epnjpGcyiEkve35Uo34z7QDgSTgqybePK2Dzk0
EsxgCtVQQEjFbrdFq+Z2k+3VdtyWJ8IqCbLGqn3LNCXjJ4Z72kK1i/TMocDAMXIR
EtP9g1tV9t9adTqUo3pp36046AibA9PwasCFhdKvXYaVJjvbezA/ulNOJ5EgGEZ/
g43Ed4t9/acUfeuEdRj13LbSqWE4QJmDz/f6upaaD0H1BRXrjryInHVAPXPLVEGG
ZEzjIVsdehbP1cKmCdlefnHh+s0OQ46k2PaRm9KRUyfrZtvGfaZu1JkEntzJ0/de
kchTosTHtPCoyiFa0R7J1UAJPE5Stm6RacOq8H1BusxkRQ4iWCGfTs6/oEEdP+8l
syAIhJ9OLUuHViGvdl5XzH1EGTVnahsy/ZmE0JAgbBeXtYDH2rZAIcUbo38sABYL
Vgq0nHPp/0uh35rArYZGrZDlixOeqONi08GYFBNDxLm0HjKvSf3536f243PqJtX1
7qgP+XvhV0i4HJr0REU5WD0ehKP5PiVBWNM5/QjXj/GMMdKE+rrX2MSrFJ4l5JSa
FLxGtZrzf6EKs4b+ofV8F0yRJvD9854Ac+mr+ByVrsdObw+WYN3CyKzANGEM/ibO
3LDnlgxhi1FCfr5Y5tnKByKPmt7hMoTsgCXfbJ+Ib+ufK6oznA4WqztlnVzZOYbl
2upuh/t1qiB4KgLHJVkhMuljz8WEpKLZENuYKw/OU1QeNNe9NwIFy8yLYmpWAggK
Pyk41NWaX6Mg4tb/G0IKbicD7n/uR6jCqzN49qn4hWP/hT/IXjfgFwnQimbKBbXa
1B6LyxBpTr6cqsGQr0x/9FE6Ua8rZRJiQDHBm5azRNIi2F2YdMlZkiv0E+DDiWHx
XqrBJPEz5nOQb4N5w+7lhivBDej6aTUxlOXPLVolo8crIIwLhjqJdTBcONxP5IKT
VIqbRrcsN/b8FIyCHICjCyjtbEpIcgenpUdZaUmYNbJWmY02H13n8/AxJyUga6WU
2HSHLMRsu/fYlXhkBi3anqoaBA9O0h0HiCzO3SVPF9ljqND0dpNTPcwbmbcstLUd
GUDkw5GR2QLUeKHIxO3nAQgtOeTZ1d/rB04Xu5nJ4+RsLMN5YGUM43lZJIUoSkVq
qpIWObp/rs9srjwdJX7k7b3F1BnHB/tK8+RkBl9n3nQQBy7ZwyejkPQKBZkMzDN8
QSOOlj5ipCpmXZ1cO6jd+m+iqIvBL/3U4wEG6VqjB+jXAo86HXjSSwHdAfFPTBzl
99udlpcxG+QA1D4XRWKmPMtY2g0/xj0+TfkVkINeK9gUkHe/HtKGIb0DwMboKzmE
vd6APFsSYBVTGxUOl977AKl0FD3oYrxDPPdqEOVNfObl3kd70DfPouJdK5Z/ujWs
L0yWuWmk/fbJxWq2CELN5cKL7BqXbzlmJW1crefq1wol9Hc9SBBuQ4YX6gmUgDeN
qScWD4r3wcNCkkO7DoDbOFl2rZPqEFcCRogPTXeKfe+PYEIKDYf63jLJT9NzSjXZ
JgJfOy+vH1OBYv2xinzCLfVnir2gSByLZKNXc6idPxpVdNonX5Zmo5gGjP3Mmrb/
Q2dIyrOCA3ACdGFusgTUAvt8WojWFivEvHzqRi42ZwUpsy0SDzWz1wh64KDiSvyC
cHJ2w+I4MC6WOlk38HBSqiKBFNrohXP4oD2OhHTlbNBNziXUlibqC+iroeUSXaVP
n0pYFCqMizL81McUvWPMI8WA81OcTW4H1/dXajqUdNSagGt8m1gZSDI51SHSuw3m
H94VUxBfHQvM0NYhgC4g9+QpQbeHRreM+M+oEKDofLl/11j3umosGcuoZG1rwv0i
I+TSq/kaCT8nWf3USZ82Ncy/WaBDlmHsRLr7GHxHmWATAkpVX6hQd8mJi2MGCN4D
HpKfcDTduF7IC+LzTxHRLMBsfWEUOLc0JCi3P3ErfnDOHj/yZ0ljpGMB+Jpjtj1r
G5vWNOUY23u0UXLqUpgjeUz7HmdUQEps0pP2y7ZaX5triYXea1+W/1NZ9v8cX+Dc
1GfD3k0aQPTCQGm6yxAMVnstjTSNJvv2iX2TUIxF4XkZLLFTvKuY8yqb2EM+XOTd
yo8F5+Fj28yIq+YbsjEqs6qUk8dFRc6DEiSOs7YPCyjpE3Z+8Vdd09P0IochPyXy
rnayiTR4LGIpaHKuXfxZAm3E1Co7eR4AtvEET2XWgwXlPj98c2UJVjhIXEEbHsBe
fzAF+0Wrz+tDyq/FRU05oDbQZoKSJPCHXa8P2fnuzr96wTEGA/WXSfJBpHbckzoU
dPNWvw77+ELUqEkIwSmEPZzP6xPQEL4eyH/rJb1ZaPjToYHXrPcfTRWf50XuVbu9
6GpJX9VNS+e7uDUPK6PNn4nY9FycvJEeFIZRCGczkck+KiV0yVYVKTCDH9jsd5/W
dnXkQDUEv/dkfSrGCCwS6Kis/mm6+Xw6lOt+YVbKqxFaUvwCXFHVdWXLw5POCFEC
N9zTlJ6xvvMod3Q2sRkICte25Edkb/2JelQ59fA3UAcWJAkzzPYagBIRvy2n2Shl
D4RnX0K/doKXxnaYKuKNJiZghb8xHhHIIyHwbTTP5wSKCr0YJ8ZuD5JGP0h4R9YP
kFHSpryjPZ2ZGnEUINYrQDeBaTg2PdmneSUgDe0H6AAetCtrnQqSfxyrT5FReRBT
nCtGG/6TzuRBR3dvEpx8vVjtx7RwET347TUAeu3JvoVxrzzSK+CdZTWHyKVL5aC7
9qpZOBNtG1YX/b9skQziO3AqECdfo7gkDZVcdVxWubRmiPvy41JLj7rEaGjxnfpi
KYEXXHZryjcUUBGa6WNH8aqUZGe7vgGGrWKidIKrt4sTm/Ses9MU6yv3HQ3MlSP6
fHPruFxsRECD0LlNNPkKX1aSb8bhhZStfwdPE0Y1CuLoo8s1t20pB1+xGESevAZ2
hrRix3cbvGvyw21G9KV1m+1qbeMWUMTfba3K89AHVqGgv23QG6OsMlw0mdWWO0os
Sigu6+9uHzQonPJjae4eyraWY41SIofZGD9rVojgTPpFacuHRLOKjd+fXvwn5yBi
UejOlEGDDNyhueS5ww6gzFbGsc01kdptjx8lAhR5TVDOQmLn5MEIr31Mg5Aw7mIe
cQNg9dhjJK+0sdr4bKPw29B9+jPh5Sy/hGCXqpETK2ea5BCSQPnRy/ndOYXMJ+pI
nJGT7qZ+NPjNpy6G0a2qoN340D5nI1HYObaC4gEZdxb+BJvFU00VDEluxJNxUleX
IQAeBs2ocC72ehXwDUNvaIis9LTDPS3UoNdtgIQZG3B6vWqOiZwy9bDQSekgdNSQ
07RwbfHdlBFeD7E0TI9RcpyqpAbJ08vIDdYz3Uz84Xi6g1c2SUM6WmZhtCbgodl6
CgNGUU1t+VQjXO5hZgkjgsDWvFJiWHFk1WsxoXqnHj907nklfqFOC+dAMI17tVIT
fn+22g0ut9gLqNVDlh0v4N+Ea5BVOb7KnSq2xzJKSLg10P27LlS/qCTec2VA/SUF
foQtLxcCn2q9scov/jYUaTFCe3rGt2bbbksh+uidpLbaff6YiU3MSIMair/I6/vI
wE/oAB33PgBg4lJSiKeIH9FzRLLUrpiBRCB1r5C/SotJj1Frl+WwJSPuBEUtzv5U
DUioP5NZ0DrA4o0nW0r+c+8ytM3qrCsDzZcUAv2F3EB9H3kcwdP5fWGssDAmf1z/
tS0Gf8/18NA3Umnm7OKWI8lnE/cQ3cM5HJcgTebBHh1zrN0hvoDznmXZQG/eXToc
Fy2pkxbQuO4mTlxN/DGjWzJBaP0dLBpSU7Itza3GQRVXu9JfeTbD0aR1zXkzvJuW
2LQMrcWoCkBwLaYVcG1/OtlqavOR2Jjlg7ecsl7EX4zO9DWQGKRsuUBAf5C7Bitm
apAVvu7Zj/abv4K1PxAhZnthuwt1OkDVex8XlQcoJJCHmDCkFjy3Th07RjYpkeOZ
VZcD7E0pWn+VFUE8aVLasGrbwjA9ndeUzbsFhUwmalOv30CzwnqE2RltSTwWdsVq
CmG74uJmkE32j03aLUMJS7l6NdPtV60qm0GU7XtXmCWTOH7qEfVA9f7tuSPh5vMq
ImbgAsAoUjvayQO3DhGOEt0HjgXxPBEIqdy/DEKogEgsBeq8Ct3uC4oAZsO7Aqt8
RAvi2K0spEvsIPm+zc+bVUQ386BE3PQ0EnvS47lpDH1DFKnROw7Gr822WXqqQtsv
lpd7oaFJQSS6Tjz/FiAAmnpra+lGSQ5II7Ho1BU35PVlB7G9QZiCc0dnPHatKWJ3
S8zeBKJjCMcOFi+CTG7M+659vPT2iC91Nj6iWhGWAd0G+r8LQsUC2IRaFSI9uHBq
9TAdsI/zb4hUVzdXe3ZkmsHycs0QavNqacDTenHfRu0K9bT8S2k1ssB5MCZ72dkJ
8fuIGjuRvv2edtHKGCWVMXZtEHpqNMNNtmVJnFjnsbGeswD99OGgIJ8Tq9RDPTjz
3jaDsWrnEkWEfBUSVgYs4A0xBd/h2wRQLiMSgA9uPrbAaWApENZ1d2HRb5TXroVi
ANRnKxbgot9Xqc9WYJxTM7adf9PcVzO1CDeezu6+9V+Tr68gCB9VZYF2o72Uq8sg
/2gQ9KV6gmHi/vYTDIUNeOZjT5ZeIgkLhilVmf2JlAYFQPcmZAlE64LvO+udCiZL
nUgPqaNsUj6+H42FTNZl/Tp5LcC6WLh6YeriZYFkCcHNgEWUgpjPD+WspvL6IxOU
es7IWuh3j3m8dTZNYo4VGAmnk/Sra7xpitIFIVJg1NS9Zt6AV2d7HVaT30AOlH5e
mUqZmDsFQnlgqruWeNOR6/7JNASZblIjtiJqEH+/GaptGTT+apJDpNOj9vcLiuJ2
i3HcWViIG5GxE9PQuY3QzZyDS+jJwVMfmZPyL+MD1qhtwxUGYlPPiNHWb2AAaE7x
HdDkSabx9HdqjM4umpaEyMlYxpDZwypJ5p7iZTjswb3FqvQaF0+B9bBHjLON22n1
SwMO2K1Qo98dNq+ZSi+7mm8uLqR2kfBH/pkxGpYvNLjne2EC5PCBdpIvwxcjzAvg
EM7UOvFq2EIQRzzrgy93zJzdjXxM8xq6EbCiJXuZ8/CuTyH+L9yVIeIb3q202mJr
x2fSK3liTC7FsTpQoXZdBIsACxi3DjCqR5otJ4BOl5rYzBx7/lo5+oQ+AZ4Ky7iF
xq8NSRmMFMLujVgJtmwkJiCOq0mf90X/+/EHDp85lrtJDarwVWfQ1KJBEkxpZAnt
STQQ+tPDxf99zlExAAczMB0b2/8TmNZgQo+UVdSHsiCXNhFfdNlH/66Agnlvxnst
OCR5bwLlURavSHey7IUmytOCOBMvjoMBnCg11UbMlmXLS9utBOW0U4FN0AWjwp5w
qqE4vavazxMT6tXe5rol+URet5eReRVjSi6T6SVz19iDGDh/kQekytsYeMlLeUbp
gzWifkw27c1md0N6R7VSLz4GNIfiUL9h0JcwWLr1N+0eQWl8m3edNVzoZMyl/i1Y
m5fuzxUgOuKgnsOjaORx8BZ9vhoKLVXxOGa4TTS1CcNWqlCNKYOmbL/+grvOCt9k
ATf2V0C/W6mdmlad1rdtP1vkOCJW8g/E4Msg9VeWOrc5ud0UP37PtR1LbttSE9Mv
blBYuIWAQ7hgSGVcQOWBIiA1n5A5zxandZhTpiZxeLq7wgsCT8/Uo25YITTbUkhR
N42xt96dRaNOizyV00ZvA72Y17vDFiccvGqmL7woIdWxeZXVfwViOMVyrWovBRsL
rONJjrQhOGIYEibFXwqzy+iEh3H2fqkqZbdxkCANe6KhUW/1tZ9ncliJDdNF15/e
WYE/4jxFeohInwA1yDx33kt1pV0CoTkAuMeRi8CHjDZH0q6bn1zGLwGiert2e3yN
kA7TJpwSxLyg5mwhByIW2zHPMfjC48qdJgK5gAxPF3BeBcKDV16dCCEpArLKyOMH
DZD6GZirzqP7bGZjfSDg3vjBoQGAdrigO8EGc0E+a+exaWxUZQ+emD4+zOQsVxeL
R01bp3rC/9TJsn7sLQEd7N9lhfL8wsBhcaQDT0nIngFBFsZ/rdgLKkQPsnyS1rZS
yzlUnmXGGnmSVzNKeTy9GEa5+bPM1EtN4AcYCl4nRQmWG8NWh1EzjZNMdP1wm2sl
AcOHkZnHCUDW87GuhI8nKXfgW/ul+O+nharT6mw8oGvaFfBpGzKuxWjwN4MWagxm
9Nt4N5VTokJVcUXPB1g1mgilXs5oDP+LXX1/50CnPQ/KyPsSfTjz+Se8/f2aI2xr
2mG2R6A8rUJq+vxcPvZ7+3eifLWfIONRSwTK/wHgoyP15ZZOCHaiYkQHAU252uI8
n1wYNUTEhvHs3ERmwOJKxt5HpB2De/zpwBIzXczIrUba0Pli8PUfhpb1w8xSAFrB
CNL3/zm/3w9DyJJ3ue4+UsMAciZcHEMDlpZd9MBVHP7ORdqAwnGf3DIrPSI411WY
Cmvc7JNT1LzZqRgBUczOOlkTMOedzpoejMfBn7AB0IpbOVsmuzsB+Fl6rfdgWmfB
UuizE0d3TthmXxtszywGZDNCecfLXoK67vpg1DDFR8b4Mxj4bFPXW0ejMKZJAeSb
ysQ0uFkTUL1hSnuH0PVdFdEUHkQAaz0YE/UCw3NQtOuICchFxczDOkwktYHHg0Uu
j+yuCHYeUAL/MahtOfmdVS7Ke+46r+JS/gOvnpnZS5cwYLxoh0C1XhVnNyt5K5dn
MThAOBI4IoNIlCUv2ZQ9eibz3Ia4nn5NW5ln7OSNQ8vrBnaUMME16v8L4gGy5ZvR
lGL2JIiZYtk+DMFFkzOfu+e+wY7F3BwoRC3+OQ46+NVJVrB4YfDmSzMqauM/j6so
kRDzlIrUpJUVlaxs3jSIslbuTVhS9qn/j1c94kpsGRIwYO0plzp++kPfdIykB+gB
kou7ymSZ2DBoshbfhkT1lf9g5dNvSTQvm+qGLDo329saIrHEa964E1R/HJo+ykjv
mDi5JDWrq6xRyNnlfI5XcwLLOdkD9QAdI2csaPbM8YKYBetGIjKqlht+VG4XSmbT
bhHajGLmpxq1WN3ne0qhTAigsx6bZlo6W/8tCW7Y953L2UfvUbTpGKuZGKe9dWAi
yAFQJQXZB9aw2P+aPaLH5TXX2/LRYmbpJszZiwivsAirW73XCvsnPXERibQFHNzX
LztGouTAywFhUOzyKHJQdnY4IPhOuwV2j6JL/NjzMobh7nHhQdyTxyAS+gByCemQ
EyDZcSld8mJvY/bDtIUGHUzkq9SsUVjUrApj10MLUVUjUJH/A0FbsMBQ3Pu7ONuk
LBh8jSKmwuC92FGE6kZ9bYWZNwBkuSVmWRY2w5Im955UYiVcDVviSd3wCDn1UqwY
JwLFGdmHbIR1ZqSHOE5oOXOcmxcp43VP1VW4Rt5gSg+HJPLhHDWP8/D/3tGyBOD+
WptdoT+NzWctCGxK86RLDbOIiyp4c17KUOOkdhpFwbuKhBQP7qj8Kv3JneCGF51F
J61yotyn64vA7vsUt0jFivPWeRlbZDEqIwWsxjRId/y1BWpb0Nyft1wjWeLD7DcD
/tXjByQOIDpPgmxUCCZoRSyF2yGP1ZuUV5uL1614ggGJPUxPJMNuKIkgdyfoARzw
Dk5cHlG0k7f8Mr/GbY5jEZCz5ts+KAZymqyo2eE7ByKZ9QAEIO7gKiVCObeMjaaK
lshLP/x1HZDxjoKXf7e+KhAbeunlz5rQIPIQrGuRxViAHEEB0ubMbTQuSmFbIKVu
TGWtg3UISR3e8P0N50C88znhb0xjuX47k/0nNfgzvdjeb7IShx7IGTCZ3Mqas8Mx
lbOew92mzsP94LjUihN+UETEEH0R0hO+QOnBeTKuxcPy1bkDQnpcuuGTsWOAKSHb
bjhpXNy8gPxGqKKv50WIq7X0Yc9T9fThlK1Sug+zp59DR3JvIfq5xJfMIJ3DpRuy
9jtHebQUyFAD7uqbvP4J2EX3ovZYzEbHlDDG9Yw8an+fmoKVrlvGz1BNMhpZwHPP
fQ86CqdaoMP69jQf7hO48jRkR0ZiY0ghgJTVJI4a9En90VjfJKPUz9ScRay2Zpsf
euGXIxCDwNuGOb9Kvre1YrSImnT+jhcbDHW98zQQ4lL9eCZXzIB5lJknqFUakgK4
MNrajxMZSx2zn2vR3xm2fHd7ifBP90C+ornxIHtOhWIfaEJeBgDyxRX5V4nZFG6g
cVFNJIUJQfGfNhJubWGrzYBumpfWsbsyARPOOa1Pl0XKSYDXTZ7l6Cv7DcwUNJyh
kjbQ0rdAfWzfEJXv8JOGSjo6toxN4ee0T3ah4azezcyVltYHxS9gl0y1pAAXmAZK
CfJaLVF1165MQdtnONIufo4lemzHzVj+0dchBktI70E+HQyNKSKv/CBIT7WHjjop
Hv36StX8dTIFuMvrN20Zh5RAj74I8OR39/1CiKis5b7VxIUYQvYMDmunnCs5ZyZU
DxhfjB6qafQgK8Difcq7f6qysVKs2gD23Z1VQD10g1L2UnjvG7H/YbrHRUFkXmXu
3Sjdb/6RyjmbfzimgcXGfEIDbQ7LdRPNkkq3d4/niFqRuPMqv0uxHbSx6Ywa/ef/
f6uFuiKPHG18bFL0vrinKbe565xXCerGEncjNTP1LjNQp5q1HHmsmStzDK1McVRj
05FodwwsDvvKAw742lk3dhEGAcnwHyOgK8JNP+3vH9Aonul/tRVCFt25LGa9E3sb
zLu37hWZ+ksjhD028PRbD49Cpe2Y+wNdUjDow/QTjtjt+00Hc0HFur7m2cByTRDj
Ee/8Y7YESOchGoM36rhaExT7zFi+OSMXCsUekbNIh/Wp968cs89HwRkkUREAYqBz
7AOC6yltBE2UgYsq5Pc6m1QTaPJjPOPTKvKnwEBps7Vq+Sttp9w552inRAnV9hXw
0gz47UckVNNc6nhKw1Q0Ue7ZTCNR462kvWQPbPE7OEUq48uWro7xEX7ggSacelfW
qi0dQj8DtDrI3bo8PGH43gf0BW2jVDj13QeM4+Kyd87A+/9H7MoOi0SMtJVRBogW
ZehRlMLLnqrBM9lqTquCY4gRxhOcPeia4UpstK5G4bZez8LAWUgOIX89NaBsR3No
mE5opyJ6giPOyDcLWZUOYndEuVrCNajUXwDTpUMcB5HdMS1xULQ5yPudvmxBES6j
SlqdSaNBMPKzoz0AYqP/hKTqOVQaBrsCW1siRpfdbfzFSAznJ4Jakt9L+PEOhFjX
+HQXdpVY9rjXZSlgFEwL7nTJu/JKMY6mP4DXEwwuDH4/kokI5PQljsIVQsR2UPYr
JVGrmqHfN2ACm03UhLJuAQoiQJd8fN54npNi41BYvfjf0FmnvAtunPps7WVEFfrS
pfpsVMn5wtTOoV/i3F4cOEcoy3GBQpbQ3vMujN9iTEvf7b648K55JVWJXJUZBsC0
yhDaSIJVauUyVF2qYhfvYguDJKgMcZ9jVGrLygT69edoYwPc9U7mcKgevde5qx2W
IA+/O3eKpu5vY65okR8Nm82z11Wd4nWmjiaEjBXMAFeds+iGwfc2ckaS8ZV3996s
msuPv6QJ7SG/O2f58EV200YHYrpjzRMi07pnZmnDdalERwoWl1qI/kYfjwArHGVH
GYDe7UuAlmG1lPRtAFZyfDtNmr2CloTPOhbryk570dSwuhRIDPgYqyh7uff+iPNE
QE0K2vH+tNGEsjGDm+L3dAtlOJ0EYairLaPMxJ3wBSabzpq08m1opB6RTJSCruM6
24siGF8UmLumeLIV35qL66GpIIUS1CXBaDRdN+d18PMsFEWW/F0XqSbg8ijG/SjV
f101zNlhr3ud/wkgLNi3CRJNto/6tnBHMLjPE78iIWwmM0Rt2mOtPXuAr8i4H36B
TXnr8xK0jh6u0okvMyaGRah67f6MQ+uKl84GGq0ppUuATtvdiDfK/c7U2ioMcqSM
jOpQoRR8tw4T6JeZwYNBWsfayW5HdpYNm00Q5JcJm4Y9G1NatZ6FJQIuDTicgflC
eFQS7ikrfxWpMQuoF0uA4RUn3ENV6I0SxDGuVzib/TYE7ad2KeJAprTS0LuEeFVf
FzIHpKLX7FPphEydFwhxMHIC41oYPi0B5EPnv6qtRBU+fNSeD+UbhNPOwxM+yle4
yXpBosBtbU/wIUU23jtU8b4orpqtLuh9Lu59uIY2ddV1tiEfmXI9dm//Iuo9PmRR
BHdtvS9YlG9WeQe8plXU2Z/zDoPZT7uC4JX7J+kK9WzFhzp8PaEuNUDc4T6D/L1Y
bEJFWJBul9/6aUg+IcNsjwfi7iDkY01WDD4IIlVe+ZesL6yIx+RbnZ1Y/GQVtaAM
cGBCJHwgN0wlbQLRDkrWK/XwNIRLtEz1ZauvuyhttNyGaKmSuIo3N+9lL/aqIVhH
m/KJ6/SZWlFm6fNHatOi+80l8J2Y6dsMG7Napyha2W5DAQ4Xcli2yNxJoj1vIbEI
byLXB4nW0STnqGGMaRmjRqogO1BFuUzvtWFhBopbGMW5OeXzF+Flv/wHJQYExMjf
mg/jnhgL5WAkOuFTJOwte46Izjyb+JiJnaitfZT+OnwdwiBR6AA9NqssfJkxHroJ
GuPQJfHsrR9vTCS76KBruRQ4m9Qq3PGcrX3vHEKXMFjsJeCiJXpZTAqtyBYeFpRy
WroEbw2RwTU7sN1c7IFsH4OV+LF08+A3ZNjbUpD2FI/NkRsa85BXrkgrn8sWqKE5
/+bzy468RP9y9Lqy75wXoBKiOvRiafGCL+ke8L3W40VsyaHzRhREMxN/9EiV+PIp
Sh5i5LP5de4tMx0WvNg5WNa40p1zgY0gSispBDKA4w3u1M6jp12buKjPq4P6Uaf/
mXR1pi/fexD9wGyjQo4wvESNCt1YPlfMqEcmKtOOnk06c5uMZhjdvtNVo9Zri312
nd5jkkd2lTOvDgpZJFVlm7hx8eBnO8c5gxU3av8lkvOaA+gOJzet4TThWbgL8pAc
wt5taCM8RG2BrHPgmyx4VCVFMhczR9WTzE5y88T7nXVuoFJZtrwXBlaRrNQPXc/q
d+PPuxrmeVLkK9OVVlWG21aXNfZvSFdxGpk4mxEEDvrEh++99IdwxW7DRva4j7DM
nRuM5RIT47+RM2G2pSRApb1gLmLyPXJDRZ2GgmMtoJBAOqVQOxLRKhEJ/XwDANdx
uH50UKLbFXkqGou8L4TaIxdHCE2ReKLoPS6yLrmTHEAN3Wz4MnHtCPvQ232EGxGE
4BkvpNumG3ZqG4E/zm05N0f9yqi4xx+qPTY5pTt3/MeEOxvKRqbGI6qnA5e0Oh5T
RT3qKYm3B0iz9y1iw2xdVPpiawWx3wNoIgVniANXIntUd31QoVTc5QNdy7tzAfGN
DNkvj5HLzTJ9cE7sAEKhv7ePOF0FIv0S4TU3OPmRG+k3Ue8vIZMWskw2w0AqOFpG
0vtaWD4ynAMouSqTqB+rTBWFH/jtP/JKQ2F4mBFGqsJa+NTJiEwSxtqYbrAfh32C
dry8QMoZih4autLzc9Le1/bgBiuqE8vGI1Ek110/TMAtUK9I1F3NRF9gZ71pDTE9
HwIDcRSnUBJOsy12HcYxofBjYivb1MuGT/PfP8/brqFtxR4dQGh0m+CGdvEne2ca
vaJm2GdziDW2iC6JrMGNvJsACf3QyyOqNuEh5XLkmrk6nRKV2FQiRhKz5uq0jIqS
QUqZUCSsHUn/7+XyGH6PGB5Iay5bjgNzkTufS+XdrgelZ90ovTfiALp+4sSWoTY9
ZikGu7e/m4oAqeVF/FJK3d7lZutR96edmVVZ0jcikGQMXSwat82Y3jLGcKY99Pze
nBvtOwL730DqLimLtxwbVGYlGVRb4RiDS4ga7JvWakt7ehQV2y4HYVfniJprZOKz
n7AV/sydsVulLp07cgwCB7fTAc3DMlJpOkGjZRdsl4+eaYoTgLeGZK6/1oCJVZ3/
b9Jv039BoVy+R0aG3HIW+I+PrC6JtqCgwp1qJnuqbKo3eu6cciNHJluI9JuFE3GF
zEtdvxCsXxzYt5OIyaOsgDis9Iw4DuzD60UqCzepRyEk181XVReYSzyTJgaWg2mn
jW0+ZjfA7O27oQEbmKEO3Qt8nbgoiYCKW7Z0WHmc0Av2wcKLWEifn068j+lRu9vF
V0FILaO/8+8b7uf/SRAhT8Vk2K/JGV1XS3qhO7FEfpwJFKXzPYgyPQTZP7ixYsg1
G2HlfFIXLNNPc0LPByJWg8/y5mw/O0gA7cY2S0hZPH+1gz4880k4BzKTpJ6hxKn3
rPTwRHIYa8WvNEz7J3Scp9OnapXUgnRtTAUGT7bsN43VhgUiM49l/i08c6hUbxmE
zdt2h2EBIEjHoVNGCxzyO5u+y/o9+AXQaHvQtAJ8Cqowbd6Z/eTn9g4UfC/UI+iw
TmxeDbAb2pR3QaVlc6GcBS/NiVzkNlWDtVSgL4/dOsom05w49ssWXdr7jFx1nMYH
JJ2UnFneYgRxpqUvwqDqJZmxO9i3aK2a9YOGYkwN9vWwfvScIsKd//m2cDPp9gqP
WSwl180ezMzUstAXVpJYHFO4m7h3tgB+CVIgR+NYYoPBMNyPX0d/HQ5RXzQyJ+vX
x0hb8G/jZyE1kq4cmLXZLRsa1Es1DbfeMuak36uOnCz8gzRMo5c4S3Ub+e39kdmE
mIzN4IQEbXQ7atJjdI63NCPwytMQsUhk3R+t935LG7qg6iUExgZCPtNXiafA7K7P
cBLS0PSyBwR4FmPqRLi5YGBK1ErXASCMYN5g366vVBaJkLeN4+C5NOuQsPlyltjc
dA0I0q3G6x+j1+xIVw4j9TfnTLPaXW3OLFXVD5EcrfjkNXvsWf2sjP9Ewv1F1GzE
Y6HJEP6Ss9IROgexvsWppKquyaDVPvliVwH+32d/SvNnJSIy2aXcgklYf0GEJZC5
ggjO3jyTUv38qACBJbcHK4wQtZYIJ5uQno1AjsOeU4lbqKh/Ko6UwhsI9Nqb15Yz
0D6gIX6Mp0yI+T6pk3pSjb3ozUQ9mZ00isZMWAZ3OOvJXlSOh/qsoudgRDR/HIqp
UQp3NCLMGGKdmigNRw4X7u+QrHtOW5LuRgfmbqm/W3AsSKLoDFzhaFPvVGSpAuLn
IRcPExU5iCNehe4eEfJYmaBBnfFaYl4hZEdmk2w6yC5thjv8FdGqaA2lyRJ7VIh6
9QFvr5A9ckHxV8habOQt5jAlWAy9Kd2pml91mkQCXai0cv3HzI/SBjV6GyK02RHL
Rk1IQchEGwCMWQ7Ga//RG0uy2legirp85UPM72vcuV/ebcAW3CtEqkg8Y2SDZoLF
XRwwjFOScnzGbomxsX539zIydk/MQ3fVju6W2VxZiPAo6L8KIcqXNiaIU67Mt8x7
u6rN8dDMCVnIEFhcwA3LDd41ifnBP+rT35BwubBdoYWJSR+7hTNIhYACFGKcozQ+
flGuc2Rw3oFhv7Pt1ZUQV+LchkZqSPoYYdWyc1xM9TItSKPaH0jPtI63vQ/q5nYP
GCvAISH3EUxcWK5muOZfeiOs4COh+5j8/BQeh881uWeZayI08yDAi3CihZB2Og99
pEGB9zTZydfPSi0cuPtUHcHrh4Q3si06trx6iT3K2VKh493aqG25IvK+3fQxekvL
mgtvJOGl1GhT4EOK4niLJbKjQXaTXJJxJBuUlMb+BZsdm1BqSh2/oWv6/TKECmDd
BOy2L0RU7NSsdTzU50aYGHCL3d1Y5DQwlBJ7oed5tvTp/yabYoMgEmxBLElZPR3i
tUZBbY7LCbLBtCR0zN0m6LqbRVnLOWTPlK4C2xq/XVl3cDN559dqSRRvpfmVUYKY
nWM3lCHgrPz0BVynt3fqfdDH0AfS8n1o075owfoSqEV+X5qfmHBOfZBGXqy6Y0Ht
AktR65fBrU5dr/JP1a8HT4p7YNzxilhV73SWscU3Ye4VkMrlrry3vmiYsoqruzqI
Pn9QuvCf+d59hGef9WFSJKb7dDP7sWok0K+tOt408srGWJG6EQLQgDpgx5SvZXmT
BECVNuPhMehZtwKDy+IC7kgKptkxeeoLijCbTVWgUD7XBju8/gMcU8Ez3/rMosch
kZ6a9x5bmzphHieYeZdhSYU0pnXokERdX5DlLJwK0q9RxK+t1xlxgoOMkRi/RayY
ZFKEvEOimrhrmZGWuUg60mieY08oOFdk2se8S9uFzFjH7iEH6m/pnUxd2RlJR/qF
GrU87q5MdhXZnS5IBw3Dy+cUmJmSDR5enFlxK+OixyhsGMoBeo9veuvvv19vTdpc
5zhrfFR66MQGZA3dRqrQK5hR4IrxBkSytid9krplop5/2eN17TiqFvXg/rd/6Twn
nC6obwe8b6TWGLILgUl3YzRLk3IYI0Up+2avI64MjQJjXWr9GCKeMkTsZVS3eTFd
1OB96SWZHSsmPhcy+XW6+yotxHgBIlr6hRtH0eR/Iw/ezfk1QuqCwIrh8YuoqOiX
hSbYq/KN3ktz1pilYyA8YAkyoXbpCjLAXLSVJrCyvxEWCdsrZJrxtcNUPr6NR3sp
S/wC/DFKmcA9UP8RrQ+8I/RGcXVod5+H94P5zXcMUUuKwojG/FIoz37V8DwFxjC5
gdpzXt5LgEI9Hu43oWsGXP0nWwoFek+YjjL4qbbE0HoYgDjGlf04eJ6RNFBIkySN
J4ydDLUwA0CL0ZOgNlFIuEAkuizX0JLc9DkPjKnYvAdvejuNdAbfFN1CimTKOY+B
q23vKb0/4ArGVhH6Njzv4E8bxj3340iYKkoyY7dZISJuG0Kx7VbdxV03rw3aXlEA
JxnpIEWU27+S9RE2Ahf6EswUn5VxX0hGwXQ5Yy6HCbty/xGVe6EXZhAFzB64oR7z
ZTXi5BiP3q3T8zZsDl0PWIG+t8P4PKYfSzb8DLPj8f9S21KVPVeA0fH7C0BbUkGq
qzUfbLPI5hshEGKhtDgCrXlWtNM194Luyoqi9p9nBZAh+yhhSFn6tDHwGpoGrP7K
rrMKMXfBu/rZXJ+YbP6aocVnTvEldVkERrtS6rOGHx85BGT1iv08sRUuwn8jKH9h
5cAP9BCToDTMZyF5NCtMUtz9hHYTKfcbdTcLG/CrbPEwXjUPp8wx8UfYrw+z9QcW
Tqr62hsTjch7SUZcREdB3xIXxVOAlqdfAZC5SDwrN7Tn6HeG2FbEqrq2hsReo16m
YqGKQccCKxdblrrSYii6Xhyh4dcSRXAB3Px8Z8q4vK/OZzEVywhRUaaCHHyvVsGn
xWlHahM05sekuu27wDssY4QfXszlWwoyRT4cVsVFKReL6GLWUU6ouOcJ7B2Z8Non
lWf878VOvja1vw8YqQ5Eh6qzHLB89AHXdgCNqpuvd8ZHGh+mX21Xwk9mL+/qNMtR
bVpuvgZMwVQZ5wQaQ14xO5DHheA8CH9gBWwiB/NZLStbxJfVYZARQOaVPEv+LjA0
VqN9A3wzcRNIGQUJziuUraSfHYKB0h/mYquV3mLCr4zsKxORhHDVJWvywCrE120/
gcwG3pTg7uRRtrOELnnCefv4pBSNl9nFjhUYW5N3+ea8Ax9N+tQYtlkuC7HK12Jc
0dsypZsh1040DZwzqiHxg5w959PPEUoSF5qIdYUc884NYasH418KrWp3ETv+dzF+
zzwDyU9qJHxnV5R1V4FlPaMA6E5JkqrngBl2kPLmXMO6HzHItEs/zWfwmOVGH386
BLp8pCWgUcLVYnF/1jc1PTmc8oU/yTdoYw+tYIEz5YjlE98X0wD1nZ9idHNBwKKx
RMsquRcwFGTf6BcF/w13RNvbF/gOP1+aZKm7Nsi6ORPXP6PMz+XsmDXlgXvexmNJ
wZyPdQIvGTZ6mFpD4otvdfZCfs+UB2mSIVG4nTkSzrIcepppeu5q6COc7ct3ud7Y
dWasgWGYWjCfqDzH6o0XRCF5EAiGCFps8GyQ6SS5cuNISr3TcV/2ABeYrkLK5agX
F5EbDY0ij/TosDW/2YeWV0HNzFCZkI30qzdOU4MMp9iBAeX3D+sEaSbxjLVrCaae
J605SmGQIWvP0zLua9bWSQgAA/buNfm/wwUEGaoabwRBwvyrOix32NsvelRBY7Rm
MyKWKPFRisizcWj+wM8TsbrYZxW6opHLu/UTUUVIDURKBhQcOy6GshNTvkqo0kBO
4eRUWaQWpUJgKgJCWJ/wpueSKzTmmfNNRy8miy0ytMc+S+WvXJONtibkRnAItLbP
KSE6wDx1LkJh2LW/t8VMOIrCz/+bfPBuMdTF3xxTDFfmlBtGUs0g9jkW0nD0OAdb
LXrPzO9sIAGLnhiuPkH9x3q3/+ZqSltdTgnhnQLGkiqop6KLhrTqgxC7cKIUsNEB
X6AuZEjgApB2okNtKvDB/ywHqVdFYeMC8j98qnRRyMXkun3YbkuJIoki+jXCl+mV
VkIOvEhsNQVAcGzUv7J83gbn/MIBrVHWaC2FZl8+T8f8tONJPha5X6Xebd1+ORs8
r1BStZBDBPmEMnLYkd9YABh74ovUyrRtD7B7tjOgbNX3+h4e4w6G8ssan0XRGi/3
b1pvUw1645AeYZdNmxQRtNiMnwYeehgr3Vf8Dl86JSah313RNxgQG/EOsf+DsKPW
mA2dfwpxvW5ZWBvp3pSsX/Evi2RBJjQeuI+55ap9p1JwBg4YwYOmfrVhn1r4DLa5
eOQN2pPjrtsCDA4vnQnIJVNDpLjWQjk27wSgk1nY5Okcs5WJeLEJQgVaIYC4cmlX
I6NEXrN68ycVrAEl3QtvYz4Qtf0sW4y20eKu2x+Cd1x5EVMoZgZyqaedsM4BhhmD
xqWcWn3FBFaVKnrGRzOFMlx2tVuxxuJd/Nl88/nQkTMLN8QqwIDSIASf2kuz2OhO
rJM5Z4eFd4hv/c0skz/l3v2tPtEdUl8HmnasitgdiaPQHeWSIbknopSiOc9He81u
6U74MZuLy27nDUwoUIin9Ezu56zebYX0MOz60SoaSsaKCMyUuKv0zKPFWSOqznyF
WkxBUTGPgSR6tUZgz9YyfeHBGF5UQ6JcTuPlr9ArltKEg7VaUV+vaMrEZKsrowzb
cIkdpjm9oaYuG/F8JaBPPQvwkUPUt5O+MYg5QltImA1pguBhAZ64vvetJXalDvwg
HqBce51+gHnl8ckPvCygyTYlqWr3XjI7yKwRUh6bYjdy/K6jHmSbH1ma4JBzNU16
+cwpy+NI5xQ+pgzWOVzK3yhydGQYbr3/sB3GDcdk0bvOm5+n5hX7Notf9dB5dghW
lQZ8veltvSe05Oee/e/6GiGOEJyT51bdNV9YFSZDt/rdH9tBJ48USiCaMIT7Riyq
lZgi8Y4DmGL/Vdb6/NbuEb+UH8Zv5um5YkjsTB3gaSBHPqPvEvpS9ROL0fNSy6aM
/bm4jmrWemv4Yw+bhKczIIAQBnVJUJwbTLAWZkYW9BsuvI2ICYtpiArIXWxaM2pE
d7TZzTpR9uW+CY7xeKHAbng9XbN832tInZLTAqEEInFXQZp3/krHM8ew4EdLX0Qu
C84aa/P5eI7OWQQNMwtZFoj4KXOgVULLisbKM0vbMYHAFAPFp+I5HnY6cp89xEHV
IbLU9gWsJRPktiJ5Kj8bB5WepWlI7bnTkHmI6RrxaIxtnXU6BBoyGOOVkf/wA9Id
aAN7HiufXJ9cV6Dwn1RMyInJbcqPXZULBXwyq5TZWBZOM5esQzXN4zp1TjgZRlCe
/dL/Gp3iBy7WrP306u2R3UPFDCx0Uth3bU0crIa6AI7GbBmHrArxy1RylFeGI0DE
iDRYE8gNoboriOrmJ6H0HU13XsNqRdSZJbs9IeqVjH5XusWogtTsDZabc4WSYGTa
W5Y+cjlRZK7fJwf9vp3C1hDwi12wsTEo3cwndmrf1cMdjcXZ5oTEjb28D58/I+Vi
BZC0sUOOSsHSGgZuNewXqbD21F7ifAnXB0CydldHy3ADuiis01n5u04D+KY5dUMh
/6r0l3bn07Oll3YlQi8da89BL9YaI7d/zcHP26U2MhmMaifV/i5kCIXafII+vu+4
N76d/ZWp1rKs5FVyrW2i6In6G1AIaB3uDkinydqy0yHk70vN/eXtaOfKxu29QWRr
muaV0U8wiTdlH14Ou7ppMYnI1SHIve3OxEuwYSLXDMbJh7cN1f9+mWAFBxHQoFPD
QwT1MDom+mJV2wz4yk8CiInEegB7RDw9UtIto56Y6eYa5kn3lUA/P/zIVGAc7hQN
RuPHGVmYnFcnplQn+S7SS401SBHd257HIi708gmSWUUraCTVnlGLxgiCTNzDzMh9
TFhAeJHqwLoK/b5dWdMg5ez9K9K1yAMcbOT0oLGSsyBrP6ouvw9hyWEjV5n8uwKl
y1t9GLoiGOud2VutYmZEdKrEnPmQiR6drlAVINP+DnFb2oovgB4dXYOUkvpdWH99
qksJIbdJbmZvUkNcHL6l0zrtcAupblgo2NJ7PVrGv5pIv5+03itCE73CmGiLuQMv
BTpBX5rG4cvHdw+CQrboxOCtpfD7K5MOlE3p8Qw8qMKhoROrUZ/ETwEf1gO7MLRw
Q7OtIiZSgShQEixv8/sk/ZvnDl/ntkyCVRYPxcM1n3+LVLwUM3ne4txxuJ0OOELJ
gnxGaLsT3vEhOUy+jkAUKtVEIS5vFBdGuiYq4m3DZfWAb1fTzWPvbnLIrPCPqeE2
sk+o4CXi47fsj4Ep83J0j6encRgE4tIbxtGKSN3mYeXxaFRz4tdTG1ox0FphH41f
NTXLFLT4O7kgD5zblXnVCPiY3b8cYDT5xh2frxyTRov2G0N5L+/JePLhdi1jB8ae
N6SSqHRUIoeNVKlqHx2tZJGSUTvmPi5XLSIg8ZNJvzOTsBpwOW8Onqpy+4v6MVaD
02dpSPN2D8VCSIQPqM7uTBM+k6oXWIWjX8TbGnMJSWFm+41eENDXLtNnNmja64Oi
fl7cSjko+oYmswUcKqszgXPSM6eq96rHp0qPJsq7VbWLodxgkvmZoLY02Y1t5duk
Zn5sLCsZbWuy6LsXffzsT46gbthFQ6vjEKgfCYXlnZuQ9c8FMMYcKIQ8FsyKImml
j2uZVSc4goGsUA5IGkhA3y8cHOu9l05FRdt9DXk8L/cQQkFXBFPXwggtkEer06UV
j08/givPOH3fhjssrhPnmle6EDEZrS0BYxf4bwWNTefcJQ81LlqJRVthQMnXu6Yf
NjVvZxIeBjRvMQPHpicrmg5Yrsrr1UiyTH9PQpLKVyQwkgu/oKjS2m4/lspDG+Ou
UvXpoUfjKiRiWnBOon3DPwyPa8fzW47hLPRt5WLbN4SL91aZP2W5FKhFkIQqXFbX
khkF0+pz1VP0dghe6RE0cPja3Y+fKXBwT6pUvbSM/TVfkwiwovcGXrlnTwuzo4QQ
FZyQ1oyhmj9vqSdkT91Z/l7JzDUE8MJZlSFGAT5czHkjl63AgTM1u7AlEJ6ryssj
EgZIZSZQq4tk66++rDRw0f6AI5ZxNjMRmxdyYYsbdmkIuduqxKwTW/Y6TsmMvZbZ
wBuEXBKGyIuWVWgVJmz15iAl0bClFZ6PIG2G+0qU/JuAFaEvJkDgKfkVTaTJ2Xom
I3M/GmZe4JOk+Ukf0s9+eOIMSHALC44DAg6JCOg0/lcRY3uZxFj7pR8NuCUn1prR
iz7PEq3eJk9C7UPCk51iI1EpLVWehGlTiR3J+7L/H1vRatOYzPe7qZMB1VsRIxvN
elZEWYZOFotCG5D5w1spJ0MEcG+sTpDPeSnapNgUKfEx9/LQvUbO6rG7ATddwoTA
Dyruwim29AbGa4Y4DR5ou0d9BDACv8wf//qVbhjY7PFcuBw/kvOr4wBAAZ9vCxIo
sVThC270oJoufvLEmTEJyyJg0OaLM/1HE5zh2oSPdXlgvqKQYCo76KneL7l15L9P
LwZkGW8d/Y5oyT8TAKUQf/MKS0V+Lrh1xez2p3+3564ZF0GIti+hc33zch96cEhk
gYWZ1VPPIm+P0LzH8m83IvTmu2USKExO2Z878iQZIius9P1A69zsPGNAv45zS47G
Bf/KXICwuQotiU3l5Ye66u0WMXKtUWq4HFaYbJz0/d5wCqM9jNJVBiJf17etvaLg
3f0VWUOI1ZrFhLF+nxEQw2Br0GHDeBjwm/PuYR4pYIQaxSZ+hkZrhPlXrOvOvDTI
MYJsrvxppTlIF8m7XhY+nqZG9HcqdBqFM+0zwARoDxE6yMN2pmZXqQZE7L59qUAt
pfzI7PRMp2I7oSQbCvUKOucsUQ82M+L9IwaPgQNu+JWD1RUqqizB6lsctvz/TQl0
NSZnX4BLfZdorqw//B2dcb2TvMJF1a5VFr/crVklx9dJWEJHlVyh+EG/7ZGCAKRY
WSMU7wqtQVpcRdWfVt/lD/AW7VLF7W2ZCNE5P3KqiXjrRtUD+A9ZJT2fxHIN3YWC
GzSZN4OY9GlEkMNVopoV1HqzfRWJ5AZWs4uWmSmwv3FumVfXHW+DnXiFBDHgCNfy
OVhwGKLWvEVFx3M7AMIdRoConbaGDPtk9nt867VUp5qigoAW+tzN+p4tjHVhIF1v
BWjTuHdA/2cj6Tqf3oReLxXBK2GoTGlKuolyeNzuF1hHZghyC8OsT7TNJmjK4dGi
hc6vaeWODRz9sxVYjVbPheISfNfuAfB8erVH6zOAF46CbdXk9iiosMvPmjgvzhMk
K1fnDJNq6Yx/HqVz+j4uKOpSgyNITv+gRs1nsIsCV+9K7ifu8Md+0WefjFMNJm8w
9WcmyWI0DSCTS2b5loMNq6Qkyjd8nfSXWKaX9tcAK7vZHE1z1k+mG10G+IoltGcK
IAGw2AnCxX5nRHaYnV6iab0IgnzkRz/lvRiAlDV0BPpLax09jpJ86+k7a7jaxdgt
97a+MBplyoz6p314VAzxxUQ1psNhOVutE39poV3Q1UJvEwji7O6WKmDZudDcgNnj
DzsN88uir7GO3V+yQs2Pa/Vqlnd3+NnmEGfUvXWICliRKliGZX4JYeNbBMED6n4g
iakfCVw6u+cbHXZR7Y8BlWysMmbYsp6t+9qosR1N7AhF3x92j9JaZppbs/EzMQ/6
VbiwxdLc5g6WrtbmSWDx8zjGAO4wW2uWAu+kx2m/BpMTI8y9HvEZx1GKnXDBuam/
Ai4oP/zL872hVnRevJQYA1KeeraRuzZRajbn+0nuXgX6/Lafs9iy3l1h71R5hqsv
XrH9/45gY1XziurlejIV0qWy4YEZDqAv97qu/yMZln+1FVlJhzdXc3ckOBox7r2M
L6veZTJ1DwjTGjO6AnNiAeitNpEYFFL472TWcKp8Tid8/uB7h0jOEQaYtHXWT6qG
dcHLVYrlPAyQUz3zh+TvO45RFgnbwhaUNYeVBK1aX1KoPQeuhcatvyXSwC4cFr+X
l/pWQiwUXqxeLzaTCK6TVq9KEVmhh/a0CxZzJEGNtdoWSJPnrmQJNKOAar6vSCYm
EkLsloYBTE91Dw4pPD5Qz7HvqTJ1mt4l7Vc1vI/OKLJNOcU3mp9k9kTeExPpnoay
Ct/qwMGaRyD4bbjERY3Q5KtMvfe7H7ddHQ0m11S8pPMdEIDfJ9fKk5NvaMnIkCQh
5B+BLponhVIGnJ8vjdOO5AER5cp21tI39g6+KF1B7Ym0V1FvWLVgfVf0YBwI/jR1
HB5RATCLfBJ7QvKmbx3h7/X5NczgMG0gKD7jteJCD+HhITZVoyxgPdPlYcUJlmgQ
Kn29MTtKz3J4T8nS+I1ds/BElkG1nYYpmcdxCpnEWrl2n8QRKF4D2DUV4pjuEDpd
772dQYvhWEBp+fYWj5pM189WbZBNllFLDQT5h+C7NYSjqOJNhLXnUyDqAjiz+Jml
N+4ZYpxKwrrdY7L4MmaBpDUnDSdJ99kJsZcYfgafv7AmK965dBNuTeWouPPXhSMz
o429+HkDtfe3BUEyWs4cjBgbNjPokBjqoouacaZA+WKrrrXk8xNAQ8xUldtV8fon
Z0yI2i4W151sX3l2rYfhP8dttU1qrjzUrBo1O3VUlc8lDipfAanRExy7n+GaU8XX
m3uR1gZZj7kmyCb5AZek5fwO2z2i4ZnIdTsJL0C/hN2VFh+BbSUmKJc4PNrr8vtJ
ECXUYpy2PxLsorXB/IE/25uV9UIWZ+7U1T05t0KywUs3RaWw/eRGVnH+dmN7DqnX
lkD/H0HGoLjtUsW+XTpy+LdgaMRDfKHu4ZdB4RLCUlXOMBEIvo6VilN/VN8XaQVB
Rtl750CnAtT105k4FeGBf3RaEtKMCaRLqS6muXEbaJEdbQtuVFize+GFuR14wrqL
tG10Mq6ktBXZ1KZmXKedLMp92aMyLR1qnfN8N5LIqSYTD0uibhLzyfatJfZTfV9u
k6lspx639ZWeh6wmNYFNSCAGEgPeFKAYeUFyl+/RS+FEkSai0VyVVwch0o2azn/u
spRA7ZH16liWSIeKR423WC4KFUMPTWh7pXBm+PoaZgUVipsFXHBCYyvtOhPyrHM0
7nEXKIzC+zdlkDEs0ZeYQnZvkPcek+w7f80PZzOHTeZvaujmvlNd8EddP5XdNqvp
HH+ErNWYTLj4Mkxhs/4i8WjGa8/UM9DypH/KjYSNyZ5J5xHVcfsBiNKQce/0GiJh
5wld8XeJ6PbQDdOT8htfDrTJUSoGYCvyixUj/xsLDsH530+0mjhbRLjhSvSrdYlt
xwABPQiEMIQurXTNBi83U0K3jQLO9BlteZ+tDWPkJ9Y8xV51WU2IFiz2pzdJDcLz
8noWGlvRCgRRSxiLVoMdVgH2Ra6V9ohPm7SBU1mqbK1IRLa81A4kPaJ34H+tLEt9
Bzu3MUgAqUPElAl2kcLtup2q3N+ZIru1idJkVJz3CmpiXspR9Lcn+CsrDL5fmPwU
yfqMYfWppYyY7T1moq8LVLGzf6m+fy9bhO+ppMlI5BTvfZfeFcmlYHfPa3Xlr7FP
s1NafPXh+r+aedl8pCSn3TDBbXwoy0Jdmzk0d9CrwH0eSwhUiTDjmn2XS5kmFHUJ
L4/eWz+ZwILdWST+X79/n6R9FwMSo8qk8HkGuIFRBA9aVGB3ZYDdHLHYcbjD3Zw3
nXsYBKEGuhTxdOiC1Ki66JG7NmJfL9utxg+DALY1QbLtB39Sv7EB/xp++kxHWuI5
HqiplLlEtAVo/SOu0BnMasIPnT251Jxe9LXYOCebV2pKkH7GI6kb+D6R2Fpam5uH
izzPNNtelBrLbSQhSDVdj4vuQO1ed938MWU2fJSb7wlpJNE0EWteLkTsvfGOgZec
YyYczxl6XRzEeSX5pxk6BPG3urmR9ZOAuKW2haOzasxclgWeXq4Ja/QbMRLnVTh6
aSyLr1LcFPSFR9Zjqy0TvLoanhhbAeFX6yaJ3AcXypAGDs5+cWytvHKiPBXqP0W+
LkT7wWEGbW6j1oSbO5YestmPOVwCagjWLe4d8bXqRXtoO6ojJOPMI4IZnd56opIo
F3/ASNifpEQqraIiIoIptSHhh3ORMpGF8e6mqLZ1imXi4TvIKwVkU09gdfyVM9BF
TCwiyfND9SqlfJrdOhdgSWeWUw9UIjC3aJZYHKFFjlmFi1Z852VJSHh+TDbMGMTR
+r1lms5V/SXNuw8qi14TsfCeLfSHfkDkhLI0t6C5YqnzA0yjU1G+irRbIaSFsLxU
JEIeH9IRvdU5inPnMSzACHsjWGKfNlBx8OMN9Ha+4hqCntcLfVybOBZG733jrUt4
QrlaJkfW2xB4qZhy7WqrEmEfMXA0lbOG0qj4yWvS0u/6Mpb4Aq0kRvjzT9ytVFpH
M2Aidwh14OkdZwc0QhZ78HGRKMUkTDbgGy9xoQiG9XYFJoMi1EL+dS0LTnJ4wD3i
QDn2nAFpKVJla15wrscvKVdelLhQMUQPyP3Aoo7x3KwOpfgCy7F2rFPA2IJeRujz
izcbusM5EWPKDOrurQpGJi3KADTwSzOzCJGzK7hF6zCrqTW6AqLIEgsl0FpXNOf8
KwzZU0m9gdvu0VgZc/3L+ACbmOUQ8vUPV17JCedCDuVVO7sUeLD9ztwyglv4uPkN
oyZiBIMRGCGl0K3hqUrIboI77q4F1eXNPaoBgxB6PBQtYVx/3GeuWqFbxEn44gIz
Z4dRZyBEIjFdIVYEen4xqCjj3u+pfl1OkFAy235FoWUaBloSmvkzAicnfDNCenM1
731rTuCa7ZuWzQFedZPHpM9+d0n7JOdnDGGEatF4ufASb4rHHbhc22C+LG4mbyRl
yRfLo8J4kaj2PLh1YIN0BZ6tsCh6472Z9INv7QsXsjjgBlWCLW8UXixLVHDnsg4g
2ezBLIouQFNDqcCrJys1cv0EIPUwbJ3ux55TOoKKIzwgMhilFWGpk92xuIH5t3HT
vUl7jMxh0fsaERuiUFkxJ9+JFUdakftozDO9/6xhSajBX8gAVPRaY16aYR5CKb90
f5dK17voowRAzoeY4axsWXEjEd4vGraI229oMzRv5y0BRlZ1dVCnyYEKokWvkLK9
PGN71plJvXuSeU/BVZ7LLkk0a8b2H7tunXNVPF1c9LitNmf4TqVUxTGZ9eAr3dN9
DHDheQATQQ+vrT2kB5ld5JslTZw94LELLifhSEeVROO2KfTh5DxeZqr7qawn0jHs
Oul1lILMy1VwYG6y3pQ/FokI5xO06CqFubVtsIVsZeU0SCFe3spP/6jykEnyhGJQ
sHt69PTDN/5+U1YhuEKayJTjGCsBmKZfZErtO7xGXsNalEo46+wdxksNMFg5rR/o
BMyy/z2/+gSO8hoLzN8+Gm4o1fDBxiBsuxB3pR59XDz7gCndrRa2YTGONoRRRSs+
pDuJudy6X9M1nCtQfyjpUZZqSmYQJsmf/wBHvglNASIxDzDHHmbKhoz5V8sWZI6O
tzc/y+PoJV1OOpRX+36ZxW5Je1eRd+q06pQf77RDyS2v8t2Ya6BjhHIl5oLHj70O
7DNpLX68QE1yiYKcQ1yYQgXSVqmdnZouDPu2Y5kqSS+zPFVP1YtIIK3xmLuogyoZ
RJlyqn0LFQ0mK45YWBHtIFWxwgzlrI3C4xXUhq3HAk//bhybTpHASlkR3jJkki+N
NtE97tmXUyTKUUARB20PgcDCOT88GHFIvdaD3rO5R49EPyowXFbtmo9is+9O9JvL
Ros2DeFSoK/6nP+/gZIfWkMkitab5UpDm0E9kTTxW2o9yGcTfc92/tbLEvQ4M25J
2/ls6Rdx4coBIXjKMIXGmGQZBHSfnidXH0fiUS0KvrDjiXKmXikqo3BnxQ0T+6lG
aZB+kB0t4L0HCA/y4pDp07/50kNcqEBU7SD5dAX3YJ1dJcG18/UwEce9G1JvaNEi
hk/uX8TkNtavilFbtsmI7PQDkmxQcrwUX3oHDUdnxi2aRSONsLVYNab3GBNRy0s3
7nCEiv23FdNjG+n1xV6Y+zV8Mz7EkoRZF75+agcV2QtjhSKJIyZZptfGdbQBtYq/
opidu0JE6TyqbsJvEyE/LT2HhJH0b+dPD3jPPcXzgLmLPFnzO6R4ZZy2K7OHM5Dx
vMCQC3TjfMjLrvLDIOVg0im3lXhSIXsH/l6Ame97IOrrk+2ccc7pSN2mw868sOqG
SMKvXKyZSYTwh+Yz7A05EihQyYd+3YSjJ46aDX2ZpY3p9MC5UG2slG5Z3vkvRT92
/Q6/BgwXVvI7MujtCl7axIr3q5q+ink0RYUixIkWZTbNeysYYKb7hST7nNHx6wuB
amtYj5Ba6LK74yUXGinK301MLTu1Ybme77Qm7IMrWpXC7NX3b7X+vOY8fZUZxgmc
PNQIb52Vj814DYASQR7561oFGUah3K6/9kwPn5/o0fL+5oqusb0vs/SQSzZasRkC
8MXC5newv1ypvDyYfWjcki9jQGpaWBO1DG6VYV5eQcR2DB+X/aLScC84Zo/mF5kW
pYMjkuIC7U96Sl8iyWJ7fn6M8dWx0w2FvFBCD9VOcJ5hbWyF522RuBgDxxYbxJkW
YPpoy2mjGZrFstuMHvhmRHqVWKZOqN5HBCSAslNd1ULCwH7Qgdgab1OxBAsoegmN
cG2xldMm5/tEDTBL2LZpte7N7zI17oedcRPARKRuWMQQ+knQxoTGHDQzoVGk6w4j
JO38Wbf3wayT8M2VBMzLQ4uaPkKLWeRSusBs8iY86PfYm2J86NRmwZNsb8iljOrw
2lzQNNiHYQhAomOrgEbNmt/ZbuoT4olaVmQ3X7xMeE8LVn1iASRNGWFzyS3kN4CA
fIVtjdWlglQw9jZH8z8NEQivHhjfe32DV0xkvphDuXW4jwcrAdJBoXMPVcEHTphF
uKeeFZHbkFYP19V6OlXkc4o0EOg2eTOsW3ttOF9YRQPTB2z3SVNIAadgNTx6sXaI
10qiWhMeZDweW8kciduBHmObUsr5jveoz4XxXgVYJnJUsp6xTL2VJVUKQVah4QSV
g7NISgQeBl61tOYxHqYdpQxXXOg8BICMgarYHQ3IfnTCz2yscrqyA9eO+kFiaejT
15OTNdF76jZ3HcIo4wWXtEdqIdyAWIfmDuZixDftB5FOTgkImigdpXMZiRQwGlf6
0hrSclPSY1372rJSavD8+x67S0cvc4aEqNgbfQ8/v2h3ciIstrHMuOiH6AO89l/I
V8inS5jJUk9KRGuOb81PCiGhwrlc6lqC9GjXxMB8SBYYh0clht3DgyEhnBzPYUFD
7ydJj13m7pWOHLlIpFmGXXp9zGYKtiA+u9N+37N3DqCldSw6+8sBhXYnqWgQwBuP
tiQ3OImTDQMEj3TrImkkutncOnkoC+CcrM4Qzk4DV8X7U++BSZ0Btx4Bdj9wH0y7
wNwPxrriL8nKffhFohnu9JzpqQXgFtlMGNU+yq282ETz3xZh7FZBSbahNZODrnmf
iqQhfLYfCS8s8Au3rA6l4defb/gAGAEoviW8iOhpj4GcL41EHmtQYN7WjSy0EZmo
6vDfmvIwRN8te/NODbfRCSL54oUxLQXOHsCTcTd9hK5tLcULewjJ5Wzj/jiQFdZt
W3dnIOIGfytriIAMTie23ZimdUtJgEptgOmShxueinBn2//6T2H1fwsd43e63kho
zrj6z26W8zY91kP9oUN3Y1hMKw8WM2ulTv38ER4g465mMuPOvVjIquGWnZnjXMsE
vPJm3AhTCNeUfMa9pZE5gPyZSbIJ5q+10MrEe6BR9TqMUd3fx2Mj6b3DL51RLyGQ
TPw4+C6nB43rU1pwVa3+k5yuOpoX5+2oBEKlr+SEjYhxIgyaU6Fn4OsIv0bUqMQr
29v7WxnE/Nnh/5FCL0BX+e2OuZ2Ys+J9NibSG8NxZb8MyIEeSldZsSx2z2mtuiMN
gci0VBRqhh3yYU70IDFaTauyPUquI0Osy5dQsEoMbnpu+G63SRYqLgFwtO57VSwe
SZcBWiSRo2A3BD5Qj18GfPAbV315IgaIIFMrkKnYmTuKzBr5Ig2d9696E6nqQXH7
chTy1hClA1j3jnzhXUXezsXpYp4dlQ0Y17WB0XFDj10p61WEdFRCp9g6t58Lmq8W
NaD2rkIvOXkzxicN/IhEKW1dPmpf36me/zJwbOOrCZXZ65H7IElGFZL49F4ufVFv
1Yi3x3Ux1MAZgsorU5Wfe8qcanXqhUb7UjjYMcK0tDgkkOlvM6E/DhZCyf6epKjG
MouQcl+EMNn/rPAgldEK+5szJNRcYJjw5zPFj6X4bfw2EzL2XjKOMTyaAfI6Pqb5
mvWPW7KVQPigIqyv57mR55lDMuNXWbG9J1sTl/Da1wdo912xmNjYD66lNCJiYw5F
6UVIvcRu/T3VTCjtgr7O8uFEXiZpEHIGKVWSU1vI3jxHGfoZOoIAH0EJ4MWfQpPn
5vM1+P6CpVxWYef71Yte/WBdxdhaVnbMO0kduJHwxJ6luBjhsdTuuuA2qC6GQK26
ZGXElkARRMygXi11Z/CB2fTDo3Z369ny+wRQHtGz/FDQk1AVUw9y+VSz8dJGew9d
7z6h+Pz60cjbMI/Ccdx9a4z/9jPNWxF3YSKg8O9mGR2WuylCGRiPv+RKtt2cs+sx
wNIPn3mdR1M7BBE4Q/nCmgeBQa/WLHddMIC6kaOPllgPRn60PUyO2U5hQrYv2tPz
hrrx20zqTRI2jTKaKtw9Du2gbEeDbpxk5ecu9Ko3gFbmKzx/Z2l4qoKY7z0nQqSF
0+1yCaLp2Dt7/1NegPkrPc+E7pq3UMTyBVWSB6RIYngMcmFG3xoAtkNO87mE6zmb
8n7pZpfW5qV4vohZkXn+3k9+5qa1ZVcGjDck6eVHIN0yMIkANQQQK4YWd8Z8aFDb
TvqsgiEApkyxqKqKKTbuvLc25YKzeg2wHIQdHmltoXStwDx6CpaBtZKMFVLpSDb6
xVdpn9k4ySsr0BFOIes4bAy5WF3VyP6YNyVqG0opyVNM8z5HjhGhig3WEQHXiJ6W
VPfPUs5kYIDH11FH/IidNqZ1coYwcc0uEdXsTm/nYjYw4UWANcfbeiebE1T4k3PD
SmkJfZuAnNu+fTmWio3lL12HoFIPSmn3MGSn73iLboCW/SWqLgd/Q50R8UDHWSmX
7UxAq5kDvVjc828LWvcggPeE4V641xfRPqObmYPyoipnCmmwzrpVja7z9OZ+bRfo
8w7QVplYN9NLS45i1mEBVthzLuNYHMtSmNxBMrE7HH5ALDOVBoa4ejnYk1coUTI7
/vK/9mSKmGFvzaKdxEr/BVUWUDJhYcZ/vqA01Bh776yQgdCD4IfnkYD+aLRHfBLf
KFwzEkeIlVCpYGgLfiaemDA8+VBfZ0jAb0QFpdYzrwv8mQOIGMh7tq/Imv7dFElu
Tb6lh6keGdLRyjjJrusac5sjCne/8QvS+GgZsJrYcC41HD3ePO5fysOMUztm6c5n
w2aQeA5I6r9tLhHUTjryRiNH3IxbM7iqDxzz/H1SWlQr9Xwukk58v/Z+EC+zHHHx
DpcM05301x55qso4XJ4wynkot+INJG3VSp8N62EI8V7OH8LW6+h1QbzSTFC3AsiA
B0n5nyskUdl2niCl+38MacigHSvMtggtpa6d+M9G6246Cv+6W6sUT8ru9oRtmjtY
9ntxGuQjTwTTVqRYyD1XJXfgTGsKFJRUjSEUa36wqbrlqmaI6M3nJVN+/z2h83f5
amV2eAT/DTlUN2GwRpo3bFi+qMs68HjkEwAq56zc1KOBykplIlk9vbg2UBobSYwo
hGu76QAwivqnYGAOaoY6VvSKKAx92itvpeVXzAFFm3gOkewNFOh35Om208W+Tv0F
VlD53HrhIJ31K55NBE9qimqVPZw43j06W/JZHj4zoi7Qj4UBgx990HwDy626xs/s
xTwfojG8EgXCK5kKYDTGMiGOlclZD53fyUBRB1rnIKdhxbnJMDOwlUMY5/PbSOM8
eL0/4MKUf23kfXaYSU3/dA97RqXbFqS0CfFTPaj9+W0T3Rt7DbxjI6OiCk7Firyi
9bZkRpM7VKedyyoNO65/NtUwBLNYRHzRfLoLKeXAErrx+/v/WlZuOTxdgAg5243l
I3RVVZyrtARyxyrUQF+u4z1WYm9r1HpxCpC1cc2u0xhMa4TtKg3ijx/Gq6n3uj1t
GcSHQBFmSTIZvT+pZpyHE8Y7wqlCdONX1T+ZD6LezCJU250CxthWA0pD4CYfkSnn
Bgvd/FDN8p24vxqJsex8gPnQTO07zDf7N4ZQERi3aObWRSpijB/j+6QCB3heOBls
eXC1layx1rh5PcBWZjpYAJcFy3sCxeMCq9qt3e7KkwHUsEUCJKXiseKqM2aUcuxs
9Mc7tHyIl857vYWjh63MCQ3GZbrkluq9FVCqKFXuWut3Li88zA2atw7LxVdkfoL3
2DsiOWWb6ngAm5GOReV2JVJa1JGxfll9Lm4AUk5FJJY0fv+x4SMY+ydjN3Eghmpb
LdYAXPhj4HizvBGpo41w2qACg/PgwOXSbR5GppMptvkPVbwvIoVJHDKyhrUuTZ6S
XJGLgexr0snhKJB2Iutpn5ePxEMXa7+TVnuCQhNwqaJ+QMPsYwFJ+Mb5wlhsaHl4
9A8rIZv7ZSzQzePITeyyL6moYowiY/1mRVYjFx9j1c1l5vL/YJMlSSBZx3yX6RYg
Y7yzEFusnsZ6W1PzHTWoct70RUYLpsD6xCxEYF7ErM27gY/DbyOmbLQJ6DMHFY2I
mh/PIycW/cnhnZXQyhvUu5Sc68/eFbKYSS+Hj8dS2ijAGsobXhc/slOlO8LgXDho
Q01Abkz8swdsQXnQf0dB+EJmK9WJzV9EiI0lV/5K/2nPKWPUKcKBuzdG0DXcCN4y
DZiA1lIuBm3JzTEgikhESdYrjeiLTYvG3o47PxIeMW6WnSe72C1WBrgjtPggEvQH
lkxCtFlmCuahcJeQ0QdUA3EknCRHQYtjcM3kGdUt2vHWf6G2b9i2vUD6rc9ukTAo
FyigpFl3APBWm5kjCP8riYS3usNla3OM+jQdP3bkhnhRv2XdnGt1aNbmhpux8N7+
fQiPgAo555+6EPkhi7EdFAKQYZymu4Dw/quUKXgIKRBw0Q8kKyUqpZ0Zm5iQMrM/
HcVgAqWkUphy1CFnSZNIX7eWgV6pRoKFzo3qgCAJUYVwSDxqlQbWv0yJxgjOWJnK
W5sAUNWIyIH0+807PG4oA3ugFXG18NsmcHxPFiVf5XzPBV7jbbkNZ3dJj0zKfYl+
DlateCb/tVuUwnE3IgFafSyHBbukol9tQQGrq7ctoRXdOmsR8Bo60VFTVKs7135N
Z3nfP/ggTpcIVitowk9l4N7ZJAzUC6TGqGeIbzVGSQ7CJEvx1qA3+Uq+/MaCwUV7
CV8NBVo/1oAVz7C7ZKYy6En3J+wqwnEmmuyWslGjQjasqq7nwE/vbFDw8pUNrt18
A4YcdLYps8I8jWkwAuBULK1/q6TT+SPZRwYCnTkwex1VW0z6BZxK/M48kcqtZ1g5
NvZTQTA2/4slS5ManxF7tArTzCHq/1FKKQtBibpLCh5Nk0IWAVXk9gB1mlfRkdDy
6THY4o5TOnckC+lMii97jHRE1Xn5kw9ODRfXHQHGDKrJKWDCGuLXZOzwTG673n9k
ZQmkG3gx0+UheToOZKa8WxYhTifA+pmRkbuG23glMPQSCg5QEaHvgPpyEP8gIbuc
srSyopyzkXAdOZjpQJL1Cf6svQmaUFYauFYwRzQpSjmESz+sJhOdONKdSH/Hl1GA
s6buou7SHo8VYKlEYjJ15ZFxbZf3eP7eL0PP5bI/bH4XIUZibXPDZXJLKuUnfGcE
Lx7WOlsXF0qMvSPYu7UR2Su6oTeZSTEm7bd8mxx2FYjl68oh6Mc+sgtbwUXkeaiV
+dfeLrzKnkjvBSlL4WJcMazYsBRzGb9hSpE4Vz/THErT9MvdSoPrK8tVXxyOWf4H
ByE6SzbIQQ3okR830z62ZOxd133QGuEfLQr7jaPL7AN/b4NniEa1lwUSkzCWM8I7
64U1IEquHravBelCf41GAqRZXLyK/krWcR31NbEPIa8FFT4mXam/q7QlsIVj8CDS
sXNLCkgtbptPI12OoHvsJOdOrV5HqcQhfk+HRI1P2aFvSo9N71Zyqu6ov7CF2zdk
g5w4fOFnSDBiDab6Eh+Tk5x8g8btEf5JDHdF1GU4jvJu0lu15Ely69nPEA9c9PqU
ffV4yxYbfQsh091dAZng8agsQF8j4QlsNIPUikrl2EBnvVtWh8YY3vYFoyzJY9Sg
dY2Q5tN22a4GRuPnHSLBga7yqhsob8qJqYF8V9DZOBGN8a6GIYszoDyLINc9Rbd6
Lky74xjVieBnvZ3SOiFZMZ9pksUN6ZlzAMBwmFHxLo5oYMIxn5ig59+MXXPzrgtu
JNSHrkE7QCc9Zuj8o12e0RcXTOhnyXI+I0QNjXluRONWZXSezoR7KWk/xVp8ix+Z
zAZ4F02iNAOZYh6hbvtc0tK4TSnq+PbtmTQttmFqYr8RTFb3V1spLrEMc9sm6pwo
lTAKOhfvXrBY9/diruh89h5YJp5/AEMxN3w1uGiITEeIeO7J5yL/Kwlh2CKTIEa8
uOY8ovkpp+X+8/rM+CzNRXCpPjAlNS40QZ6U8HbCgWK2XMlWRmvVhQLpHRdoNJJe
Y8G7dD5Ek5Q7gLfKi0/vMoKegU5DVDAZTvyB8WT8hNepMtPaO1rTSFCeZ6VG6oZ1
3iBD+VNlXc394bTyhq07JX6W7NMfgRzAV8ivmfU6QZ6FEs2nPG92OHFcdlWavdlH
zl2dimsAnI611gggmdxNorqg/8S8hNXnKCiu3O9GhFdWgxEoJcaH39vT35L/M0ZQ
Rv1p28qi4V/UFa6iR1mDCd38eclN4YloH/4ilojuJQUGxri71amhhd4JRzJw3vHA
frMPCwWFcrMGQHf2N/0kfM2dmE/roKjkZrq6kB8BGcgJExPA3iTq847l5VbMPasy
fKXjr8BAoy57vqgZ6k/OeObxGjYvx5iMe/Sf8i2JwtXZq6kBudDKonlgsIj52u+I
kqmTgi1nNHKtCRbK3qvPuZxRaB2+nNqVOz0asccPB955onSdIxTUZQyWsF3pWvZ7
WJmk0cua0stcLP8vYvLGLa/B21+u0Ufhw2RmeTiKoZ7mDzyTb6YxWoGCSLAdMsAD
WL7HoEvx+GlU3sCnDZ1FzEN8iyYAZaq0w05I14BjHDsvNq8ImG7q5zGdOSLrC/xR
owW5S4ILdOtONQIqLt3YpGALynH1Nd7XlohsBLV8bo9tKFcbpihnWJRzYHeLYeLr
t8gCxblk+UVDU/1LJi5I0r+lAV5hZar6TW10GSQFaaI8PujSVQGCxUO7Fhx9vM4T
ANqQp4jdk+016H87RHtkv3UwRwubwhgxUHeOwPCzX32mHHSbFBmxFy5PaPRtVm3V
0/6l7LhgdKtpZL3AIKtwXW99i+z/8hSmOsKWpUN5Wtf04+KrRKN52yenUv0fFtXm
jbqe2MqWIhYUBkD4FZY8oY9outp5trnWEwWRZ+EZ4jhIqSlbujQe19+eVLDLRdJ3
GT/o5jsvhQ1U8hVMzWE7XK36CeCfojoNg/OfJ0wPsGFIeJR8FZm++JCfKYsbyuTE
JC6Wb79uLaV4NIFiBAGhrLhG5TWQGK2xpd8DRWpRmUpT10aAW3Xd1XcJe26qwHhR
NQ/gY/NxOgOYGK/iH1cfG16INv9cQSA4FvJWBEtlmw/djAG2jtDeFsmC6S5xSK3x
rqs6Pdrknbb1ZyfwO2dFeGv5+I4+lleL6eaEpzrVp2P4aCk+HizhpwnSJCRSj+2T
mpX/cmEMDJCmsPtcVUfVCR4bk87Iq3u/5v28GNReJtP+pDhY7fr5UNWvA6Pwr3+m
nZKmjodX92IlfsKMNJf3JmBlePi7Y5PRDD54+svOnehF3M5TclUZIchxXDabCiEb
V1hbem6aWjGCOAi7/6mQA2zcFZxLpHTrGIfN0Tfjpk3Wybk1Um5M1NNdR8QHiu4q
t5Wmf07nHN7JcnjT6byg3ePvhn195uJIaSnriV1YE4oJuu6maETQf9sfSf33PiyO
P+F2FKOKbhx9XuyS7vjdRHdmhzRuEepeaKceUIFPZkpVfx5UODvQCgHGD4IueVuL
wl2jIWi2oUJoNC4MgZZ2qRuCV8mlidIk+ejw/yu1wO1Nk2/BUHl2WUQnkq8UOroF
g2GS4p+v7Jm7R26YaaJMiKJTWC6xH5XFcHxwnq6ZgD3/hIOYPksJpTfxWN+S7EKq
fOAy7rLcjXisBFxv6FKgXOKhWoKVdHQOxOrILN3dj8S1sScbPropXYIilnmuSvxr
TxpuqWahpsCldeHEKkW0kX3L0tNdrYWdS7LF5fNmIbmJOnhNAwEPyfuzWhird9mo
NSq34016gTwDkHEJZ6dNseCGipv2F5MlD7gTAmozPOI+Wrvfj3GHzJ1O7Y5WLh8G
+D+cyfjOjj+JJpb7VmB6uGeu1Bt8LYoTtiFqw6Kh/xWvY9sEZAOxKiBLdlZquWdc
6gCVpmr0UjMTWbO/m/4EgK3gbJATTv2jHNE4gg2RQKnP1e6C7kkcqlOf3+NeeA1p
e23cG7jyFxiIQkgmLYNRYCg+5+obW66CGB5ArV5lk974qyb3hnRKWcs9n27eMi6a
W+vvnJek5/5HasEci98bDfCjjMVXu3p0k4lcP3SVDsglkrr5N/R+hpQD3lRzIEiB
O5BzokTQKGoMEEJpxA7GJOujk2kFMh+amyPJ01fDN5p3DgFoWn+WP4/jPqEjLOHD
MjPlqGCboywrhgFpC8z6Lqp1RYLFWnx4/UwNztSVg5mmX83kMCnEcymPYKaw8eJ4
Pwv7774h8q0tCeY1XTc+Mm172K1BVg6sNwez94o2cXmMpVBRJYDmyFjmfEtaO6Gu
161ihBXAiDLH4tEqwhvP27DoA3rjKRAHmDqguB0H8hI4oun/m9v25DuHmEas7ABf
4lYS+yooblpAv0m24K0sGB3Ua0RZNMb4+zviwb+AWClEN6iIx1zowfLP7eeIXGrj
L3F+/zditwsZFohAauz+CpKuFSyazk7adk1604B8dsBkiyGuWr4RVD/EZp/5U5Nf
Zq4ePhJwjJ1rFO+scz3/QuiGiEW5KiD3s4ZRX66bwi/tzJkkX/6HaT5V+LKvxUi3
i5KhgaElYPZ5LXQ6EiZ6o3fSEMFV+ytBsnsCt4+DucG9fMeUQa5lgpf0KFwS/FPL
I1kVyRf9PtL7F+O2vvolrkeKd+0cu9xvt7Mzyh3bGF+Hu6Sn73uiIAcDn2O+3FOL
w2o1o8p0EDDE13my64el74y5cirEv3pF4wNY6d8rwe3FcIAsFu9bk30K2S7RMQcu
HGxj8e7i5daNJqBHjyj6+YHF2Oe0pDq/Jd8TbJiqKHaBHQTu6QLzOYXdxPM2ABMq
yAnTd3I0MI0oz25mlKFnuiLeK/2fLkVDFAs3wZ+ZEOEwj03ARz9Lb6UoOjO8DWCJ
6Lw/9Lr3EhP5UVNnNtjoBrRgWjh3fl9FTp3SJjXoivOX67OzEwcUoywJVqHoAnU+
Wuhc0JMmun+TUwcKCXas8QHEVajM3kUmRVspv7xon71dDNE8sEd7tJEIBCHjMgJe
KfPdQPGTdDGtFcBMdyrrZKTSv6OkhSONgtTNY7gK08mRsd+KhnidihAEwo5ot9bP
fUQnmmPsXaJwI1lZ9k09PqROBX/aLC2OfY8QnT1Yrd8m/PKUtC5lJ5E+uRVcPld1
qFY0IOoUbEPL6aLh4G5iYF16Q6948z7HYIPk+4uG/kzksa7HzVMsPLzfstGKDai/
ukHGehQ6b72qbsP1fDNlfrF0NdggGMPxuf/kwzHBka0n4lhCJGPfRBJgwkoEjb6c
51s4aAz3HK6HfnfjjxJRI2gOxlgIoGr8j0lzxvAeavZIgGs7cFkIGGvBAlQRVgRs
HVLTVMBWM3/RqOTLcWFQIlhAWv/I/TCVim3bL9DqAwVpnNgMOAwi5A1Ijib3Cr/A
VFbgQKrrL+ifKCV80C7dt1RQD+khlV6yxVqdU2Lzsmm9KYPIf9ALf66v8Uo2jGVH
4dSjqq5UsZFMj8As2o4botpcvaVkOwAv7bQl/FLOZfhHu3hqGlPHvLRHA9Syl2+i
ZYrrXA2yqCpxbF+fCa5nLF/WthOZFOopwBXpgx6PnRHdscjmondTNUMA+ewwaFnJ
Uit8sj4UC+fiiO3ML90e9Tg9GjeoNLuKlFpSYzZF0/NKKdOx/CtozFilYNaRW0pI
YMxzVipFMLm5n813dGDorCfnv49Mv1UifnU7zH8s9KGTlCmWx2pT+wxeMKOBtNF6
Y9TMiV/4bxrnON11/Ogf7/ojj/hFgcNkZFTOuCle7BMLJzJohXL9MKaY5eVokQYA
kURPkezgzYygQEFbsW15lt+vQhScJ2e3xa8g9E3C9Hn8D0ciycx9lAQKuGR/E4ir
cyRhkOihThmV+qoQKhwtr8t9O1P2POCTE0hS7rL1am0MqRX/XexqJrssK+Qr6xCo
oy4EUah9/JAl0NW3CRRTMQi65OsMtFs/QLV4C/JOSGoqQ84KJz1wevbdpEJ1aTEf
5OX+RJ7CH+k+F8YlkD61cHg26hg2PjsvB4/QbZvJ4ehUYSfZgRtAub9TsD6cusNy
iEmFJDXyhcEF32DVluXhOhRYKD4GzqWxaQ7gZqfhdHKZvNVMSOD/hP3tJwkDAhwH
hprCPy4JxvozyKNNUEWK5z72nLECKwgVPjZ9mzZ5LdoEEfu0fViz6l1uhJNajyhB
0LFFR0Mz+lD4Wv19gGH66XGQ/ZDLDrpRhXhafm2xUgVKqHUvOnuqJ/bBS9rseIeK
FxUPmcdkAxevbdlou3x2VmHMSuyBzeV6uGMyxg1NQcS5x8h/U6IYTU9YRWZhwvq0
GewFnb8DzhYXqe7r0re9WyEjxKsw08va1qR20cPGncZGCbvSjhEEMNZHSVd3ESIV
MP7FE0vbFTsqEJlwJBoVQOylYy8FHACiM/EBU977yPxpsueqAohMqEiXlVJkbXqf
INBQak/cDHGlF6Xx1KIherJ20oo6kdbfM2ZUafZG0HRtYqDGnHAfB3RWpYKrjlmy
SUgYFAJG7hJUwnNdpBAj+ZITAZMyB7lhwaxJbzSBpYbnGMLLtqJC5ztnu3FZ45Mh
Z1yUKW5WoTC03PAiRDQo2FIsSpuViaXCMqecvP03J5wz3fRvxAyJ0DVOKiePj9yK
JHMieLWHfQ5EBWMhoj9cdNThHeogaonxtJLDhoCDJWkT/NESUi2JvHKWl5iRElQU
bG9ALhrH6e0ncjoaQOL0YGnG7a8Z4+HXDzkqhugm9fz4vAAc7RpkEcdGvEfb/Wbo
C3ptb4M45VHPL81HJSUKNJ624nCm3PMGEH3kDN4R+QexqeJ/8IWxxrWTkZQXttCr
PgN5CPKmVhmmFm8zpHokdwNpiJ/GeaxeKeV7l25IBA9KtAQI+ZCYm4poH7Ba1HY2
S9aTCnNPuxaIJRsNjyZ6h64Bws2yy/XS0L/US0CXW58QoZ+hLhrOYBzzY1/FCAnu
LCoeN7Jo/zGzmScnypw77pinvO+s7UDGUfFXxj/tKLBEDLbk6v4evusGAcIbO3Px
QSE6JJFsKdfTCM3gvCs+g+/YhG16sBzn3FwEYF2s00ZUdL+vC/FL61o6LBKz2TCS
CR26i7YbXt4H1GrXouihAZQN3q/3gslbP0Z2xRqra/5rYyZZsc5IIDvzQcn6dTzJ
kPCNfKLK9eTJXqUNiuiWWnm5VTW47CF/GYZwvDq5pZM/W8ei2cr9iQt4fbB01OFp
IhV/gFz2AGqy7zLJ8/KIh9b9sU6Li6koiNxg/7v3WJ83VqhESkrmum2AAcMpKbkq
sGJXcQ36y70jnhjk+rY9GT9FDNemI3We74aEilo4Xonn/l+AEnPsvwbRtdPgROli
vYcGwbUUi0nO3TyesHqnZ7HPc3y9yWdhPmN2wOrlxi4aVKsHZBvaK2b5F3Gv/GhW
npYCmU0epoKzDAhZMACXw3DCZF+S+cj3yvm2wJZQWVD3RXdreB08u1XgMnV32DxG
7HfOCTFJcbYBb813EZ/Or6EapWVdhrtSwqBpUtvCh9x8vqIi0WWas4l7pcRZ4mD+
4qEjWh5aeC+obs18lyhtbcgRO+ja7MBpKKo6t4IqfF/rH6hskiPE3b6YlrdvNZS9
GYbgmkun+vqvwifd9k2r08vQHmkIJx8m5xVefAoePM8r68lvaw9XaVnhoeepQ33Y
11uS8WWuAGCqf6cRBKQD+KrdHDXNIJmlI2TG9d5PbH1VnsLLnxR4DHoA/KIv+DTH
M5v/lGLFEoFnqJFWdzOyKBv1jdu4H5FyvsLUwcYvq93CS7qC5vzL7HyFvcdyJV31
CtkSC4GByHcSyDJ+sgnNYDwFxb4knKNXY3A6IBeSfEmXsdXpFY8TT6sXDi6IiD26
49GTp00x+b2hjs1v1l3IS8FabqT8iBt10EZK0Q56ukVz0VYJ2TzG2Ntct512zycQ
KIf8djtQ1i3pO3AzV8XE0vscpZUYuBT+DVCaOidrUCx9avu9a5e9cUc+y9QNJXnl
bhquHd+ltpQVo3O/iM5T2+v8rOPb49Bu2mPjqhLjsK3pZeE9gqY2yU0rvebJv2KS
tG3oROGsndepTj0Sb1kDsV2NcWMB2m+3TGexcqlT/A8W4gWcuf1M0GVBAarTzXP8
jVNfQCa+xAqz26L0yMtP6YK2j5mr+lkFobLxRUuF1kUOGgd0efx7e4PGz7Whwkd6
FsKnJ4SkC4pfnaTlQlhHTEY7lzvtuzILdDSjGueWB1RFFZnBSDy2+b8e9E+rceJB
vjCXZalW9Lr0saiyMhzp7uIakxvqUlvmVhsVFGhZFUYFdtod+rJQ71e8VWmTFt/S
KDs9EBniFke/uh6qDOR6EMsFB1a1VHfg48kVOnLsPGr8EWSikPV1/WrKWARAizNa
Got49oZd5PA+wR+MpsK5Pb7LwZqYslHZbxGeC5zmtAgSkUGwvu53PKPAPMeb5T05
Z1XCBsqlfuV+0E6SYwfDTc/kghUBYTgPeBfVN73r1E0tLtvZ1dye0Jlc2dO2j9zC
HNgYfmh7ArZOn9bxpx/rRp7pf2Zoy4NzWzDjBUhucn95a7HiRVAQzrQhKontb9IU
5Q81cAzWv30/kuFMF13DIX8CvVq5kRbrVWrV6yxil/pIyjRGpmueSAfCHVAmbIl8
ZtcK426QBC/3BG3TRaBW6CiACliawh/NTv9/lRyKUDz/+z4BUaEEkqsi9GyTzG2w
iNE69K204imDyNxdUOPuWv3JCvFtCBc8XkyU3LSYOYs3gyLs5bR+kiGocbEVkg0x
LN0kakePIWFgz7czGpT1VulPMleHA/ZIeE2yq5infmiBetT0q3Q0PDs1b/3BTiox
kucghkX8To6NnPkU2Om8w27JDe1nwvq7TL2Tt69kWXgBcWfdGrXlYejMrcPRzV/d
KS+1jrhZlelYbCKEt8m3flTFcrTvpWKytGF1860+eIMVInHEEPdcqihfqDHHH8KT
8b9Wwt2LIkBrXhYbRrDRpaWBTwuAwCY+tfEwZ4MFnz3NsVWCSDfPqBSDPZ4taKl2
fRH0Gu9Hi0Ve+NyMLNsUHLrqKHGby/sR/g+HMqk4V2GUEAyjex5kpRZTLLcZGRaL
gJo3c5W0/Tnz79HOvjdbZnm59CGuIMfPolVvy33XcRa9YmeYWiBs5VlnZ4IypFDz
w3Dk9ma+BCoqi8JFSH7V6bvxsIVl/xZRcs97JcfPqfBxiZRLnyYm3zimFxRnX++t
JPTTLfQoZWBmonjDHsyYmqjpyi4YcZVZfM5sYdvKNdwt8UqhC73TO+sBr20rG+2l
lvP5YtDamJw1STbY5RZ/osTUg4m8UehkOSB2HtbQBnQtyeupnd9RJvn9xrFqJOYT
ECALvgud/yG2qi05Xtf2xlL80T4mnELN0CszSqyEn3jkZAY3V07hZrc+rtzY6LAh
y4nyqPFNVABq/UBoGcCd7b05onMhxdm+JDnsYzaivsUbG5OVwkAUsoIIVLZx6FBc
hfIK4410B+JSMqOKMf9uQNKG0/rq3qyPHM5rW+eObINoVh0AXKvDDujnj4x5jyh2
iGi5yO/PC0EgyVTme84Wb9OoHYGkPyJXSPhyFgsjnRumfwljfzmJuJobojR+mv/s
mwVEob4uIiGfCLiMCxhAWlOZW0xdMSnreD0ff6PzYpwGeb43y+DTzhE5qVFgA2mj
d0115kk3GHHVLuuWD+jO5HYdPi+ZewwtGmu9crIz+5XfcEkxW+kvGmjJ5HUNLvYa
150bMzXquxdlY7PRBVHbRh8zj0R8Rd3zvdGq4ptT/cCLY6wpfwUnXUwf+3UwUyI4
xuOrvCQDYGXywkmIjQycg38xRLomjmISVxULhaNw1aJGw+X3fufd9jDbR2SUSvVe
BTMavkJ/rEXTag5OkOv+mnVv2DHEmUwCwCK2o34bevqsm7R0pviu8MPikcR+naFy
KxtkfE/K5Av2JPjNK511ugTdeUCT3zjX4it+PvDiFeXTubVziegLGZ0mUYCw3IMS
/2YgUHwgRyOTlqudty+TN2nv803U4IHCK7z4eHzFUc5yH++Ret222zZRnAFRQDrY
HvMhJ3T7Rdnhb9U9gz8zuThoHc5Sm3t9T59OavqFIogUZoP1M7FbjxuYmvsgYAxA
IWUynSXVtUx5HNsvoJ3jgdTOdiT0LBbjpdSVK4nvgmRXqLLvD0WaZz1VnNReCzVC
wm37w+oaqp9KIyvM6QJMnEBkJvxpWqjqkdOGXPVmStFu8LgT6KuHOytwduo9Zwli
39n+2yjmaA343Zbmiv5ojHOb/2usIDpEH5iQ8G8+jG5jcpeUG0D5aE7hNuq7abL2
5b2z37N5I0c7ogWUv2AHs8hx2jr1Y0LA/bB5cSgCeiH6QcOA1VTTGoSQmOCjQwgr
vZqR59Gt3gZ6ITkMRxcUkpdCiEonH9U17fVElcls1rXHfTueh4s/ZLLegjE8Azor
ir1szeF94WkE5QsD7kHmisqdN4Shkz5XKLNK4z5pYYRz8HDrP7uyQJ/kNj7r4McX
BL7rMbu8/emUNKzIOiDISDyUNU9kwdN5KbsdujwjzGn/1M9tUHTcAtlmCFVrCGHl
YhhRK59vDOfAtPVbRUM3+c9I2TvzBAZL3kXmw5VlXJePZqVnjgTBpI7tbmDbtonz
VaTQJhENu5hVSZVzDHKj1fF2GftccDINSRVwE6h1pUrjM5lcKLuZL/SBZlkCd8mn
lW2/ByVfHUjyS9CmVZMm4/PaRf6DJg1BajtZLOome88fFGnwtzATKz6IMWed/ZEa
6sseyeUszqwEI1T9ELMBmr0OQphXFyFPHkVjkga30dexaqdereS1/mSQLotID54x
awfSCgtlQSayDf5aCBmv5v96f87zKuHd4EWoirWMWdyhniQOw2OsUyuHTCByyC3I
y6tAfFyr2UTPWYnvqLIdofxM4gqgVHWuOVqrujiyTS3reBnTY/rPSLwePwtM2P0k
kzF18URVBpVkN0g6oLSocG9ruUWiAmviPFIIrsVPEcHPzBg6jebTHGn5KZJbsyZP
PapTWjYRr9mgAi5CQxSfRG1420uJB6E8o+DywcB24YdzR5TRd9yHVbgA70LHlhu4
pd5vuHfsjRkpmtXVOuW9JcUP1vSOhLMR+G8ihuiTHrtvx7PkIPn05yFYScs9jKxg
dRKyQK0trWZLsIIeOM00UyJqvAdvp3V0pf6b82QOkFfBtFYhldrH6EkccftFQXVz
gNG2DwbQm0dkeHhq7RWmXFC7B18FNbAmghnSPHuw4HNFSCH9MlhmndyIixZsNMER
C4yYOQU1xZACGLNFy98ath0ESMmA3SLEmyAGaaDic45px96s1WorBRIhhW+d3lvt
D7ZS06BV2ElEiSHs5R2QboAYVQgSMQhIdAB9x1VILJ+9jZzQUjtEQ5kUoZ+8HTrP
7bxwM9YBXGsTndTwfTZoa+o/r3UqCHTQXr5Jr0i0WdKFbU/C/LZydG0NaiXmlKLA
FPT2LRWrYTTKJIWec0hELazQsqalOPWokrK4dtZVcl0ZovTmTngrrPpChVuOjLxV
G8rHV7evM7BiQ0vQEy9SC+eR8bDfpeMuzmii4dvZ6qzmCgMCSdLqMiH4u9n9uC2q
kfm8g8RI8ChLIfEjFnKLPezbALgSvhcZB1B+601TD1HvatQ9p7Mhjlv8Fuy+wm7H
3wNVUm8WWzeVUf0JeSyXb7T479DnquU4NQOwvTzxGgbXud+VF3ROFwHyrO+TPNFV
+G76OIZrt+RE4yUx/Oczu0wQ5brHVzruRCohy9EDSYFqx9j8W8agkjdbxAC05fDS
pUN57hpOvRvsH7jVl51LaCVwknNObQMoQFRB9qCakOKg81T8d9FsCkkpvieCGbZF
P8SVeb7IrurRSmaBuq1JLj8weFltT36veNKWB9RYQomjXMaTZD1x7gbMvHc3xnSK
LrInmh9u7trK8S5XEi3CbK0YkcxPal7gJo5DumTmAZ8cIJjSnG0kkEGKPNaWG847
lXWOxa2n6THPLLyo+4rcCYZsCtl9BOx3YIC22Yao2o488i5t3wHK799SpD6L3O9K
nBJUIioRsiNYYCZ/JfMAWSED0dBkLUyS15fG5YKhcV8vDocu2q3sTTuCgWL5pbWm
RPN8Q/Vnv5PVbzUgVXoLNsUzjzftoPWsuT6vNU6W8RX4NrlUzIV8ZRUlyzenRqlW
+mb5jNtT7yMjjaVB7l1biRw/8LOkOxPeNNg68BqAtTxk4UTllclpFiQTwg5iYBU4
RMEdm+8ukryNoQhvy0i31EjmWxTYVzeXadWzzqZBzTgpNXjLduZiQN5vkVJE4bYN
lNLAHhMuu/C2y99xE3slEteK01/XAmBuC/36ZY3wgtjmV9zqeB0YIWDVJ7JP2Ea1
LJ4yS7St2OC1Lji0t9xkjuHs3PpgqmcO9cb+0HR0A6I5uUIKeXcmve6vRuA7Vql4
gMNjBnOkY3sAEAa3L/ddguzz8UGgn+hzdpEgNRl8bgf9lv8cv4kIvL/Kj9VWy7hu
1g6HHdsDw9jG3Szv7tIhGsgM52SKDw5KN7bAFnQP3ncbGMmoSx1mkv2saBxs/EHP
ovSG/2VDQpyQJgr5VQgJvtDd/aNKKyC7ySu5zH3yOPCYlP8oeMDuP3JxdkiWBVWo
AqwY5k+L2NKuczyM2Omec8gPFvbPbifWkWCWiyhGbP7mbAF4gnsbWm2vc+8ZEyf4
DCBvAhTplmnFwtTxc5NidqPYbScoSwwTUncKxAprsPzf3+28n+p/72zWQCSmXvI4
DOMX2+QWore86JpWM06t9fzCYP1yDI0LVuep4S9o51q7eLYV1hZqXAlPZe00TRHJ
Z5+9lXm+6VNvk60qDQ+vA7t428hz2IWLmJnaq0OwAkZtkkqsqhqxEQp3YsTvVtN7
8TUonya4/0YNbHuiYlt5E4MydLaZVE/3DhXX3MnZXWOGKYO0j1n7Z5V2KFCge85R
GH6MQJFs4lH8RgOkpWxvzVL+6UGsimu60I6XVCkQaLsoGTBUad2RPkaUw+lKonF/
r90HYaw9jWvgeBSXAPFYO22Kgu701Wpu5TohRqLBJa+0ybzl5zt78HyMGRebpCGu
rjh2aHj5dT6UnS5iT2il//meCP4sqiEBWgv52LJ70ifvIpvKNOKj5xT1otroX3PM
CKPpSU1rpqAKG3ri0STJMCDOlxtR7gvOgyE9fWJYZZR1p/iMJKHoEDhMgzkXoVzO
yF7KfJHr4Mip/BzfsLhhrp+JAIIvP70sSssbRxxD2zBv0O9s/5RkYQ0Fc+jDv2I5
bcDhk/7J+ttetLvSeKF6HSaGlX9rcA3ykDeJVKq9PuIYRz1j/eQuM8mawevaJfJM
M/WoobVtIjqdHm6q4iYn0s0pTktDHJLyjPCju6G+Y9uJ7t84VpM+HVXVbkS4o79q
eYRTsWhu5w32Hf/BTLvLhO6hlyLqcvZAqh4TPTOJphg8a6OaiO6hlrTd0WrjObNo
Q8WkwNyHsRf3Hx8TQMeWnSqhf+UPQOS+NJFfHlDuYe6fIhbZZHuvSvm5wUXk/Px3
65k3BgbifBlJLvf/6EiqgzTtgVsoduhTpqJnbsHE0foI4ly4RrVle3LRmwSjYB5b
FJ9e+ZJJyU3Ii65nlrXyGbAqJbFK5JVtZqfdjTqukhHMefsMPAl1VDCr4YL0+N5i
9/iD3W08quOr709o8C4C3V8oOWpPEtqOpW6OLUwj3+HIRPewu/5bijPoFVs6vA2S
2VdbvtSPQhuVrg8lsc9QPxoRSSavS5vzn4C4OnP6TXGg9g/GG6Xaso1RHQEMRnFO
10r2SUhekdy8MCZu0TCzaLU+Z2QAwQvdFcdox18qNBxC3U3Zhz8bHYXgz4O8BWwu
l7VQNa5IBftW4vmredqZMfLwd5hG5O40/0GmGMqrjNmuTfr0DOOxrizbjTApiVrc
YFNlbam5vCDkxod5cwL1S4lCHgQvlk3AQGUOXCa9/ZnKLOYiT5xcM27Oo/d9948s
ghOgiXjX1tkMuzxKzVSCws6KhpyL4k2HFbBpPTQr3R4xhlxS0qq5nCosxoU8z7Yy
BQyhmV7J7rOFWchGYYTtzwBt6ANj3qq2kmEJaeK9ef54I7ho8tgnxQ39mRNWBOBA
RXZHsYbdx9PuuGVtK7iVsz7PZNWa9d/Ye7qjo3rl7WEg5VOJP8bPBODdflRxr02+
yfJPCKNOXN9jz7944nucuvl3m5btYiOCMUkMF1wRgGuDXUtd1+6262JyNyKmZQg/
9Bhnks/Y7iE3we8PdlvSYncTHKCCGwVOsBE5yvBG3SzI4gmBmbcF3BU02cfEN/2S
B2satwKA6KSn79ZHgMd8EqQG7TuFyF0eOQGKzsng+TWnS0ZmpHoBfZ+WOzSHD0UQ
wtgoh3AcT2QQXe1y853DehqGp1DMBWBqtu744oHR7chVH70fdMUVTqfQ7PiSTUMM
AKDMDhc5Hlb+nELdYpdblypJvBMV/Jok6au05mQXAlYKjLaPgRLht0HCB45h7Oee
XqH3+hN+un/jyK6O8MvTfuVF0K387tB1Cidl9hrVdc+o4Hm6RY3G1fjSQetAwlwk
nwAxDszSblQDMaSkIRgYytPxcSWGMNlvp1EsE32BcZAfsi/LCCvSb3b6YGQuAA1d
I1iunlRsLhHDmrgcWQzNDcJF/fWF5TaEwtsskkEmeO6lZ5tQk9O8kXaAf4vz1Ra9
T4V1wSj/jA/k4FYi4YJ4CU3D5XFoWnr2QUa6gb6s51vlQkKHKLSzod6fcuVXtnH9
IpNkFV0oICoiUGd/xgmv5PdFNjv9Q2dSb2wZhEF2PXWRHL/GYvp2k7o1bFYoojYY
i8WZi/iuh9PjCXAgqSpfi3iYbCPmVMbcaN3BO8ASGPtfVwkV2OLv5Ch7gR/AESLL
KpTSvl7LhJYyoB5JVo7m0RpwxAHwacbc3Pc149KC0+xX6hlbMvgf6y8IxevYqg20
uzjjfNcNVhgRjzZlXeKEGQUUUI7JovTwmpXzbr2w6L1aOTyu0XESltHXtjoq3Whp
C3wapvgNbIYD7Oiay3FBo/d09idqV0F3RS0BovfdZ5osNdGnVT2h8NOMGUBQLF9c
OK4Fw+yOoSG06iwCCI4/849vpIPOZ4tDZ03wm5pELLwJnkm4br639ANZy5br7w3U
7gKmIOTYrz4J58Im6if7+jTc2qFbha+BQ7y7PEs29+oqBAcnWwpH76v8+4gPzwH3
gex0PQLpRD1zsAHYicyFw9GFCl9ddh8Pvy4vg0pb86awrTfT5Nj9IWM+H0Q1ocoC
YA6pQ2FSGwWnpyrwCB2ZR8/qJ0NAmocDvdWMrm+2O8nahvnlfHgo8WOE4fiMRIQZ
tvYPB2539TA9U50qpCUhBIlNn6KnSG53/sA12a/GBbeqQetMu1WZ1T43AgToUQm/
/WheWhKOhxAPy9sz2SnEKVM/+f4kIzOex9cdQkmu6onRj05eMNdJG5Q92ZbQ983z
lwu/DCGnu5tKWqSP+UUOwT1S6Bs+N+4Dx1zpZFZZrtJIuM6dPfEcQIHJ6lOpWSVw
q0Que0UJuJ1aJsyWIsIYzluNr/Fn1kJTnMcW4tcDpzwyi1sKc6YPhfYnSd6Mq98I
FIFS8U4aMpTEzUt8prratbQnxpZERTkh1xYDqP2CmCuPKmuPgpEbbRomhr+9s6LI
2GQ+PfgLSjf2X/KRKlqoi/lfCHxmXT5ZFnymPa6JM92TLGpA9nSF98QJMOOjNHGU
LQyuNj57YyvATOgMBRL1dIqL52nakW6y6L34XSxShqDdP2yDrVHgkTm7PLhJ5bf1
go8bBTyHHklDgC6q4YgYHuMhqLv47xxIFeNB6qxUrBbd3qx130PeiHeysA8o494Z
TgSfhYPiZDxX3hlnSJokCOWxwPzwIoY9u0DWZxbg/iSjBqUQxtOJqEDglb/mR43T
5MvgqNm1WMBbxHRnIDH2dGE3c6DYu+IG+P+rWF+SvTW3HA6h9JRjD2vY1e/LMXEs
07v2dtSkY+af2kkBYRCvNaScpgFLvbj8Q9Q9pxkJZIAclCG9W3Rnj63H9fwgvGWY
cFADAUfqsRVeq7t16bltY8b5CPDEK/I1QoODlMmvlMraSTVoABItnfXTjiHaYalI
vIzvHLrrbqtUMxwHv8Tsxk6G7zRTuEJ9E2nFDWwFGx10foElur/XcKzkgAJ5Svl9
iAZfelZvVbcYz9SEi69nePN4ClofstCa/GBDTEcnWJM4KKWYqc0COQoGxoISxFiw
QphsEY4y3Bm4gDf//M7JRYqQjyvUIgbowCIiLEOtx2m0dBSy9DwV4iNvBUr53QA5
IGibM8V9nIHUlpEloDKGPvnf0FYOzUzGlQsWoqFgQE/BggE/9vUrWK2Dt6AKAeO5
afZqOyEoFppOedJU2YY97FZhtMo30VacQJd/U5sKTYLOLbRMk90jjzt0woQhpbuq
p+p5EtkD0/L91+7VzmPXAJO7+o8AoCf05YdisFSeAQ0A5Gzm4aZ+hEfb/HX+YCtt
565sAld3vXBF83gNw+xVlPjsrFyeRgQE5OfrBQFL+lDR38Jto7dH045YOYTu4Zun
ZGONsASuwEdH8JVZ8/CLHe9TQV0/J2wL47c5Wcwut76CqjYuj67lW37+xhgAwlh3
j2lu67byf2Ov/PSa+CCN8NTvL3khWSn9pRrNOXOjFS0xrOgT5SbM51fwfg/1KE4G
9ybpKaSV2ayubuAOEpCwEZcULnKjAiRH6/z3r9YMBi1RkrKDWoW/XZMV0ZyWj5zL
3W3A4iqYsfcBpLLpKumW7BANH/15rHmIpNndBYHkk0YSJUjp2h/b3fEe93uIOf7q
p4FsNQRjojekAYoZ35Jkwm0vZqFbdsyi9hVFikoFLDYFKCtSYdgyp28r/cWsj8na
784CAvY2ts7DF4jYKA7BHtVL8EEZjkYXLweq9pQDYYxyzVaZ8HmCxjnUL68B1r/0
0GZnzBGtQs2JCTwdBpcBPRDVvY15WpOEM/oOAjRymvo1GeiVprBGaJw30lyHNLk1
0OWt8E+NNjsKObx7LqJ9p3RWy7po8Kf9Zmba4AIsbhnttOovBku/lVxUnee4o2BZ
Rid5mAyiDa7IyCwcXTDkm+4owuYqm1CyoIp47xl6nMplL0M6rq2eo6sFjNqz8Klh
Z+TRdKeFP1hEC/4uFGti2JaPxTSfh/T1VQfjBdU6qk7UN8uFcVTrL3snp0Oto/Op
G+cRfwdFHdFKAAi6NMgVmrGG7q4nv2h8iBTldaseJqUA4pk1BwvP+7fZzCXjT1Hk
NBcjTu5C42571zgvb/SlgeHAkXRR+58WXsI+1M9zL48UIAjTit/bnWOYVhAgFQC8
2XU+SZgvKPG9pQSHHWleKxk6PFJm5DMfX2nvlHuqfevFB2odFIsm95DzY8bT3G5v
e5/xIQK5aYrlY9q5agyUBM2mZHp9RBPGVXHZLhWqi/v+n3FnCtR4RsVy/lZNIJqh
AEIvkqsleAjyKukV/FHtcIr5xrUZ2thEmxcIHtldr+VnEf2gB8qouwSdKiLpu/vy
/aLamtHpLtvZ9NX1WP55YLRDKZK7fDmM/EnaJAaQ8McoP7PiOHqTmw4f1tAsLcXh
14R2/Q8I9OPLHVw08HeR5RtqBKqqNpvAk6jH6Ql9ABPu07LcewFF950+i5cBtpn3
RTg3/rR6/OxZm9w2fU/sXDyFcnSXTt6l8B76SzSNzMBT5yD7e8gitWJa+PY6fDSJ
hCq+zCzyD/Cm7Ix+NfkIUvIZj2Pnupes/cSxeapJXJeqgCFNCK612vGYqGSRweRt
pNh7kU9+vYpw6oYGwODNvzJHJWQg8TmPUaZEX8FRuXD7EEM+80TE/gaVQ7I3pWk4
3Dgho69SgQigW3Kap001FFvEW6EeAOdmeAZyy/VA1oGMZfzIaWa/BAw8UthE+0k+
9fr3dyT49JJgNfP+knLjIfCAAEf/93fgYMIQo88ERg5W429dEcqR4iFDjlaIBY6J
flN906baYdjrtMyvB2vZ5JYy7CSx4KU22oTb1qdGDvp6yvy4lRxZPpPiBfH0toX1
PlrLhjaQXW/2x0EIhAd5a7YI9OqlDQMwpBKsgv0Fsg0ksAEF4h5aHScmFWSPP1FX
IjXrR4hGJs099gV53OkTwOK5KcEJ4ANVUG28QOQVIIU8hQ0LS+4fo4LD3aXf5OCq
XwW9gMom1FpOkrXKMCjo7tfGIEOpaQ1potZu5rIrXgvM91TSTLLAIlxPFYWZgTME
PxrnbD/9jSh8+DsyHd0Deyw9t7vF5UvKWMeiqG+WakRqbFVsC0xRhxWC6K/Zx7/Z
S8yJpHjtoFl6nta22eEG9mbkJeFg3PUSMANr7ovwMjbsdVJemFbquT80uL1EAerU
sZIzhofAOY5xErVCyytWLpadiWAbKVwSaAsHxTw6uiKzkgUWRjaUiQEIDRrQNKfR
qCj0qbvhiY1xJwbHshcs9TUMEPQ1VdORWLoSKBabvo4yoABXRg7s3EwH5EmJKUtc
PJIrf47UWqmwsIRQNQJIVP1laVID6HR36Org2Ova6l42YmnCRL1vE6wqfjrEnjDz
nHqkFynAdOuEDqsQ5YhdfuWgGuTE90fJFSM3dZL5tHmdI0POwVj2wSZTV7i9uAOa
uLtDb0CI+79C88rCaytNMoyKIsJ9X99FhIrTxlw7e8dpTw2DBgMectVol9VLM5mY
Axctk/RiXyASEdGT+Wh+KIyXACVG/4XwfSzLdmRhkHuTM8NGluqNfBcO5MgbLHzU
o1+MpnkUvQb0/UhlHOOxUBRQH5CDoLp5znUjIbq4cIRwKnyFVyKve5iS0dA7On/h
gb0HWHwAoqeD31wm6fzZ0IWkEKanXIwQnmJrVhMJUP/CONGzJ62TFsHV2B+VCZzm
ENgkqZaFuC0rgtBKksyRYX4/pqUlr09uB7zr05DQuVMGrz383hLMOZNdd1R7dcjZ
/k+n/42/WWilk3CSeDcIKqsGk5azruTEN9f7fPZPgIKvE0OvRVvQwJSwnO7p/Oyi
Uj+9RDaO/uJlJlCLV9qH/J5r1RLQT1iTpeZy5vPNqri4TiKblhwyxSe9jTFIzA7b
vsnA/9wkhqwQyN+zOdBq5UZmD56lEa8FjEVp0A9nurBnsuRQ1CIhLQNFDC7gEdUp
ABoSjfcGfwSSlpV+Zc1KnBRfYSE7iPH/Mur2vcbTKlKWGcP8ByLIaDMpMx+QxTzu
MOtkhEFoSnj0q9OhAi5yEjY8lQsBx6CUkAGByv/H3G7DZ2aMSuAZpuLWi/O2ZVTH
lGnbBaOBZHDFUdtT3I24emDDwm+mHmopB57GlGTRNLpR1aOE26b0gs/bX+jzjOC+
kUBVxPXnC0hB9sC2y9uEp0BD5zU5j8HHerP+9BXbeEeVkSZPxDGV23vyU9Y5258I
uJuMp0Y0XeBvG53pHO6t1ceyZ2JtfM4J2nil8BnMjzq5svlzEK49c5nKd3Xw11o9
WgDue4k3Iu9uLVL4LROgCy0koohf8SQtzaILRKJ+syJabJXn7go3qIvnWy/bQhO2
gdBrTLUdXHc1tPyzrNRuwmzB39qZLV3tWQZMCi0sTdGCQSP1kCFvz1MEL/cCYloL
lVC4SnykCg+QiWCfahP3CCcJBpEednXTXJKZVvIbEruPhfTF33flea/2OfaBufK7
Vo6ame5zsA5TM5liDoq/ARaqI91nZY/gbBV9TM1tWLf9rsU5l/0bICJVC0Swcm6X
LE4b6R7+Dt+HF41Rq8BIPoyXx6gM2anfn/f4zyLW6XgEEz3w6EftlxPsE7o6lQe8
Zw+hvCxXkKwsGTCqSmqse6B6OtMpZ9cDRgVGXqbV0AN+15UuCPb3fUrB55g/JhmX
8vVaJP6ejKxjNwXk4pWwdorfQr9ffyz/n7ecWrgzm2LW4rP9sNRBc89GTGObtpnU
5Nog1DqxmJz62nvG7f78geXCYMwDEabdM8cIcau9zdFGbloMkIREsKLm3Rd29Sj5
h95e3FlvBc6+K1lYBaUJN4a/7FK2ZY6Avid9daJmK0VCjoob3RyhJB5QTSpI24Vi
5kShoZk0kx/pTtuEHYKiluxdlGwXIc6RZAI2M5gTb0R704+cY48miJ5vmvBVl1OY
xS3pDe6EMsNJUB6kMo3HSmIbFKU6hMJ4vHoQdaFbt/EBlfX+gg7rdmjDDxlVwu/K
UGvnQl20846aKEAM8TXH4Fqxn/vrI98RKNL7JjCCyUJ2JQ+oTHysZY9WyLxVyNT5
uSO+OXYtLRh2nHlPLXOknraoieYe5DOEii8OoJhDxMfa+IjO2AzLqkht1oIIGT6I
7Ql9YbfoOdCDGQkWRdQl+yT/S+OvwwhVx979drFYSia1O8beXUqF1sDquMe9Ykze
9fX5le+O8woBHUPNTRZUnbb8JjkeiYLjNciRRW00mM2GhY2+cBM+VSS0pixGKsGQ
gDkadHeMJuuOk/xGrVfYCUEMa1Yw6JBkgpMKC9hdyrxNl7PKoPh7evTvane9FDfX
Mn+L3wVGImvdGNtJdZ3yH8JH7wWA/NUvd7G934vNijJjfK0/+a+GHEkbpYrQMipq
1J9NYj9JB7YNjKU/VrTn2t52bdxCj8spZtQnersEuxbqupCpFKDBjlDrkyo8udwT
tIlQLvG3C1RN4m7cBPabtHzNH5aNNC6N2YMGfkXmsrzpqAPebFTMaCfJPxW2lCuV
LD8xvuaEbK0syCA2gDdohTMRGHqwMn/GYA0i7zx1cDyffWTcBZ6Cb1whv9C3NbLj
bZPWkvWWTFVWL6fvVa1XGnbPiDC4ZExIc6iUopgHQFZGasAk/Wf1amzqscqrxpHu
HhDlqBGQ5vYsQZGzE45FfD72gXgC25OPFIGdVySA5rhGbp/1N9wNSLJTMG9d/GTr
9W//LslVBAWHdA/nsSmlFp2JO39qL7ejYY5W3cr8uH9GDWrwyBveywB4Z7IsCry/
B/P32ZFUtYtYmXdOM1FjO0U+4HI8VlfQq+dfOFNM0o9hols1Zx8x03NY4GW9jz9y
Ufb9+LjN+PWlt+GnL5OXNqVsDiLwfLV8qMDOnU4eTZjeTjazTElXw3ms91fWBE/G
cOxgbrrGpuquYw3yFe9OhHhuvzrilBVUZbwe85NUN3+8/vTYYktAFjOZJ1SdHL9O
PrgFyOw7/EMCohar1w346ZICPXZsrxlckarKYbkK0ufKNyNMyspIZKhhaDD1EZyO
yfVyTPCr2x6RdyU40e1TMcCOsv0XjQ+x4SVI9PBIHLnGdfgY8FLgAM2idH4m1dTL
daQXOpOKOYv+AZopJzaSShqsCFATO0eiXGBbs4c7RtXnyTmUgeK4hkDhTjBSx73L
D+OLotGb9ll42jDxLaoB0lWOoW+3KYuS/WMC8yyq9QTg4pyXZTA77562H3fdToHU
glu4E6KbJX+rkhIZSeP1gFM2BHOCwDyFJnNJ4DN4E+yfE6luYkDlDB9RqfX1ZLVv
V6gep0KKpQKcDIYi3MtCmzHkUkV7Odna3ZkB1KGks73rEZYbfk5QCLKF/pUQKZYR
gviTlp4S9h8Lok/WKcCdcKQLHJXgxWDPVSR5YLMn2Ti0r/mIjlANW8+0BrH22IFc
dWhpB9Vn29dvTTmsdzf+lTW5p2Vfoo+g5kRT/q2+JCoAmSqQZm2KjwAc48VHV6VP
ljUnuWwfthTbggRg/MyXVf+I2esHsXGlihHG9+8OCPElaBb81gVEzfikPzQh+Y/K
gTQn0cpYtX+Zvmxj5bw7r1kWXL0i/yc2Y2WwKxprruDRaBfMEn1FJkf9DzkZASoG
eV51rDFnT9u6Ps3gI7xmQQbiA3EK5bumpetvqti+r7xcxoZuIDGlAAxjVH5AyhDI
dBlv+2xY6dprtgICTXYxe0NQp94XkpUcC2rKaD2dRsvqpgjLfoClldqVHm8sdvTo
CD/J9qNIwAYzNx1Mreedggg1ICGiLE/VBGBG7c1br8Jrs6xboEOJmM8xWpRe0Uiq
eLn+N7C+Sc2et9UMDa6WD/s1Qfsn+Qo0dZ098sGTDlUbC4al5PJuakIVO1HBvuCU
I0LckX0Uc3gcdUgI4zwqO02LlmbZ91Hj5uoTdDT35JrgJVYTQFcXbVVBVkiXeCoJ
W7C5Ra4ajW4Exx9Ie9z/zTWlUILQ6maWmKUzIaNAeBog1nym/+6/TFu3ar24PFZV
SzC2zapW6EGQiQfVbAyHEbulsE9p9h14XWdLH8dze8DY7wWy3V+uxOWNxZIUZRhb
9e9MoLDjlOgc/cI/v3Ve4ukzGczUXctjvbopnzNl2CTGY53RmdcL8PGgOdmOjS+p
ZVpiKSjbj7/LHB6K/sox6XznRPwCHAbGKJlDDgGXmD8ND1FbMDFxox9Hd4Z5yqo0
LW4CQoBQmcFl0YRTBi29G+mCbgZNFWJOMoDvwRnemdA1QsI1tsa+n2L0xeSmEBb5
hZ82YkLot3FKYUnFVfyAk+1UhLJgsbRU2Ot8a7IlP5biIdIzTtR9w3nrIjMRwUE1
YYuOdEyroAfJi0qkky0D4gLjOGGTLQNVgGD40i3GAElMkvEskVe6CP4QyIy1CQ6E
Ml1NbA3jhC9mSZMFi7BLJNUummfZZb6NCgm2XNlWsVznwnOyJGcvFJVXvwj8btG1
eTXMcYzvLb/PgXp9mpxO8ebykib9/dxIvEnirTTEIUYDRPm6IO/Bd9ltEbEEeYhT
pUDHtYOpLw2GZFMxsDwL27LGq6JFvIDDNujc+7C3oSE37fakWf9ACL9lW8sab2MQ
kMTpFnfVvMutc94NXqSOH0uS0+x2QqoKiJ+HTOCh2AEhZ7rQP4TZNcVZVs+U+1v8
VUlMzNU6wPbMgXBfhIQdI6qbC7vjrzjeU4bLzFP5bjhHe8zaePQpY0pjs8QzjsE1
I/MsN7UPCBNwOjn1qJiq3Qf2yc5lb7nnSnmGJKnCmQJ7YqzSpGF0/YwIVZQU+fZh
6M/LjLvYfVAvzFYTHGNQqJFHinVQIATBDeuJLrYoROiG+zvKKoSzAlWb29smHNRx
TBVVDl1q/I0utfnoQb8+HkXonf06fHUqC3UrA4UXqKycLqn14YRXIueQeGzsyrfE
TtK9chAxyHAAX86B/wXbqREKx7y+7ns8B9CGYTkY+GFi5ncm8cEqlr78IRA6zyQq
z1JRdLC3oB/C3dqyW3vv+ncK6fwDUYL9l4H2Cf/ICsW1W3ef/CbeeiQDsICU81Cj
L3fTwauZmmk7dBSzdv18aYERgcWIlXqO1zIIeIDfPeaNNOpuINv6aR/TkzlePr84
Si8SIrlc4jsrW7yxpFlAtKlNnoUfCLCUvp/GZUZ2KeXROSyZA4EUJUVFW1p+AWeD
AmUiSGvFmtNhKfIkg9qANeeYHtVbfVfmlniEJLo2xsgE7ULPqfHB/XKoHev/4uHL
rc/4P3rhrx1my9ZhK+fff4kYUuc+OmeGB407fqUCxZNXIGvxZaB5vGxLUVHatJeo
DI0tBrbCE3wymiPiqiETBj0ZtCYu4p6Ompw50VTmGV6N+klsHaxmUkNpjOXtpxW4
7CRWu7g0/uc8AOHW8eW6IDoJqy2be5PkcnMkmcW2vAt/tq3Zd6AY6xKeCj+Z1eQZ
HwNE7gWmxK+LOsEpqrjfJlOIEYQoLdMR3AZHu+al3qbcR9SkDfyYQpZtZj1zZdoT
nu52r4+HfbnF49+WQTD7p7N7Kk6VIrFQLNo3mgL6wPJVCeU+VQfWe1jRJFO5EfDw
r841RBgjBDW4oxSqICTLpY6OIxBjEdaeqPIfr9z246PdymzHF8yldgofGePRuqmA
IpYljxYWPCZfINwJLzWhqeUqckhoucTggwl5lP7/NBaooJwD6CbJeX/hrTQXfh2J
dcnLt4FmnNaQy9ygN2V7D6vXctmBj30gk6S3WmAByEHqPLpXpefwA6jPqiT95dl8
/LFDk67l2ikJPh4YRyEJQGjWUPEmokIIBfyEVZf3Kn6NZi9uzsw2iarz1dqpsBkc
Kb2tvnrHOht8nbnnaEFG8e0wzMaUyFszO9alq25cvw7zQYwl8JyBC3c5inUnb19k
Ma3VRUnfdvjpIXskNbvSanXth7ycztrTOsMRykYMHozkppHUbpSFlzIlPQwNNFaf
ynPo9oLBYInX8adcX1+RDf30/Cb3a04YjB079Ow0mebYzL9OVUJX2lQsM34D1z1d
ynmD5bb+aI1Q8bVWY2AtXOPdZ4HHtbtpGe0Hj1WW2DqcP/rdhqZBZ0/3lcVUOMbi
N5O+hCqERaiwV0GWE9l5FNz8Dn9eWlsKBy0vzC1lFTdvqgl5ai1t1oNTclHAyIGm
SyQsiAB7X08Y6JOguBedthmtPUEXJfljJeP9liIPP0HyBRjpmXfJWJjS1unn8bMP
txYiJHPjhVKncHddp7/E65Tn7B2bFO6PZ/Yg1BVY3YVHyLfjSecLhzfp7CyMHo0N
8GaDb2tLQany3EmFzzHQqfTd7S179FmJXnqP31aBX31mjdQhO+ATMyYM2KbywBvw
qv+57HwW8l4htKwVwGuamk0q1KgdSZ9d3M9Liu9glFS+5TOHv7sCXRTHIvGI+5lE
CFcT6woISN4kHcdQLUxInkBGjyNOa2dUYJUpYnbt2Vv6nzqf96zZc3740t7NJh+O
XuHtidduWNrNcp26fqXm1E8nrON7f/3e9q1dHJ6lVshVh9RLxD2DlCjK0eWWXBiz
VMJiT1vSldHiuugc9HCmAiaN4mUkOnoU7s242riX8VDbYiKYQhujxi+CU6ds1cDv
FZevx5wjlBEHaV1kJg6Wr0l6gFlzRbHMij72Tjf2WPrmH1xfMoSRe3TKeNAca81n
4pq/xe7WGYfK22stgkakakoT5rp9NwJe4vASpsTAX3ooWM6zrNwY304AeGAjIJcC
12kDU/GiZDWLOLB+TI/Z6jJ7LxKRmP1MnF9QdvY1StxR537d/TdBmX2ONVS8KWJC
4AaHBjh1uKFXwwRSnujqMkw1Z2Zjml/JfJ62EaQfYjnOkLO5lidvyLw4IqLh7k9M
sCl380+ZKIoyfyI/pIzF8hxJl1XysoMhPUOl4n7aBksiRpvd5DdS6rocAnGPcuG3
8nxcXc0PljbCxq/edKZsh6tCXLXeiGDohUaL2fiIWiIICET2urXqrJMBMZAm9RX/
zQGMkF9AOSvmFQ70SHnHxc9VFo9K4ZAD0jbtvdpvDQSGQt8eSDLPFsQYPHEp0S72
M95zy5lrkkpgYJfiX6ASv1APEvb7soR7nfdl+CXeYF6Do/itvbmWA1EpRVAOYVAy
u6qiUhhAhrKn3dSM6s6t2r+Ofq6AGDOWVXXi4fV4FnWPObGCvEa6J3caJrWikRVm
Sr5Yny0V8rtQB83XS9gwXNgSIcmspFAY7Ma7jXqOxRrtSvH3NxvRvQecbYLII9CC
jCdxcIq5iPaH7ckrFsSSkgmXNOulcoKBr5O7l/u0vBShmYyyxWUtYLCDkGvf+Jbb
d/1zu5+zQgfTrcmMho79Xw8QuqyeUN49WowN+ztT+zm7v0Mi0qzE9G2qS/CTXQvS
PgQGMtZqIeRkS5OdfKivKU1px2X1BjfRVBttXRXJY2yGrALmWSlFcGq/Evty5lky
ziQ5e6wcWBTOH4sDFPyv2eV9ZbMCM9c7ghIZb3qh0jME6gjooH2PuIzxLi05Vfh5
/RQMrOHsqnbJg1aEM9lpYcY9VcBtaVbUuyTShiucbWB0ViWDAbcdLBXjo89Go9Vc
rC3ZcnbyqQtYMRc176zvWqTgWn8/nop3VbBUtEt7NjGaDbizLjEKZ5+/InsMTDCP
mSTOWYSAI9Q/+kDlxlI1So6j6b3P3gHcw8PNqNihOH07lSxGJBCr3twcK+7zmtqz
D0ab8CRoK6Fcnj2/VGdLvtaZYWYG6f4vtfzVrRPQslYeeUrn8FEmV5SJN2UHItiH
zLyYAASbfORpDOA0hE7vt2/QBV7HTFJvwCRBjEvh6asqajZkQZIETFU75604AThw
Ak8BwxeLIwoBOq7Mo+DVs0D1w99VJqey0awTQFMxwXEtMZsgdQ4b6BABsVoExvLw
CcdUtTTIEKLeJjrWkCaRuVFn5NKbSmnTvhabB58tjn+/EAw2ZAJ75OBGRwm+6aQA
iVzXSsRxCqFtTrHZJLxiqxOleB9mscWsdtuIFpZ6zQxvkRNBdO8sWDnkfDbbndp3
Kw0JMz8ksmB7PrGb5+jgwT2Tba7TJwRey98tZ9lfrNunVnab8hC3BpPTuNbccMJa
kbw+3H0V88WtJz8Th5MRy3EMFvsZkO7i04SHsftnyaMPCNVzv9KQFuOKp5x/NscW
oHykpyloZIAWCmUbpIVHASg7V2ecg5ETvSalIQfOp/jGql4aXAs0Lt+tHbseve0K
bOtLAxClO4+jfoL+GES0j0lGX+jmaNGzOV71c/JeKET0vOa4RiM94c5D+Z2zFjNj
G2lMuSaMQnMBIrPZOtYy9OSyoXRv1oAsb1z5d6bXP3sX3oG7mhs6AHTTZF8RPhrw
vvQ1bOYaqDOYPPThZtmGdakKrOsYrswrZdr6CN4dkOqWjKTis1JWjktSQNHV/w1z
Gjyo7LNA5cq4dJDHKYdl6+yzpK3F0xdU+tw/zWZ6ctlkEWMzMAF9TEWyRTntxUnc
dvJSW7Jh8a4yAfhc9AvMAiAby2NuQ/8sRIzJOG2KIs2OjWEtTfvQoUAEG0CO+/18
wMKh9cr9uLya4tWsEEiaFY7dHIifpB0KMHpXM9BuWD+SK9/xP2/FUsSjbT88+dVH
9uMmLdvyOCIE6yJ4S8KO3l8L24NgwGF1AjTYRMdyuXtBySoFYO8RLx2EEKjS8GmW
61RTVx4Rp21nzeiTJvMrFLa+SSbyxGIyDRgK5J+8XKxKanaNbArIFDwci29fKPNg
/x+1slBSjGi+Zv7THu5CTy3yamHUBo+ShrSMK5tdHbvl+6XDtzAxIuniKe0eNhTk
3qdFtXmFe601wmTLgxm2TSmwUF1hiFuPnlPOs8x/9T+1f9jk0Z9OH2GwX484JxB9
qpeeNFYknGQ8BeexMAutgZ8+rJhX0JKxdhZ8dxUG8LiqncHFzOZ0vxfoAL4YlDFA
A+1B6Nu+Xst+/VQMSiCPuXpNMBOzms1UPFLqEhfLpmwpJCb2YUmWkBVAd4H35uNx
j8GDOfQDrH0ri4l4yD0nVTQdV6rbBmLoOmYmEU9d4aIdRUr0WGWruysf9+X9Xtqt
3M4nwVJ/Q58PJKvjPoXKWR6XQr4Bg9BuLJ9ZDNALu5UFQX2O5lBHdmUjpwfDzilY
8GDoBW0KU63fFGOlreoQiiju4QtfKw5r/lGRdg9m8fnfedEZ7M0yy4bT4WoGUz3p
/dYWYl7eaxywHrHCIQLbvpFVvlAvIpOl9z97Encl4RdENTyIKdx14FGfFdP7c1a7
SqdnHowzD4Yp9ffrHxg1WiaE8hyTQAoZoDu7s+mWY+OqHor1o4OQKnC//Sfv+Rxy
0O2U2fjU4i6IpulWuUlEZqdzhdVk2qMbOuUDW+ubYYwffr6QsT42/7nPYLY9VPMU
VeN9VhZPM0AICyLGWXKRCFV8J1gWJJxSTY2Vh4IkWgz0CeZONd+X0pbBOy68WA2/
oiSUyEBWDjZdbp66KUjZn1dDP89zs5XtBRUCzlCo7dT47LKJUed2f3Rt4SsBflmc
g9uHinmtwGq/uF+nUaB8GBCbJbGnzXF/tuA+R8jM7gxwH6kDGH0JyZ5OKsYNrfh2
EvLKR7lPeI+pbQ1wDSjhTtmYX6cgNfNeQLJrBmWqRVwne39VVuuweJOcCnDYMEP1
5VbWC6eKSIhg2XCWjAwL1qjWYKRhshC4YIVffUnqN8TvZWCQEok+M1FJlb3YNYTP
CZLYGZG2eoN0XoYJYu+8ik+M8pe6y6xnm3BH8SC+eOCRM3qVFXIpFvU88kFyteD0
2jdED+pOuxF8odtjI5wRQeNkxIH5ZUiPD27PQ0TIamqLsaB7giOeQXBa9tTA+cY6
U9mDaITJDDiK+qDK3nNh1eilHAfDoWRjTQG0j49zv5eB2YAdZfr07dcmKWJWI5S4
G7hS7z/5JyK0k9ESMd4l/owzBAjRHt7ZcQ1A4oIfoq8XToRVNl685RwqykXuiPWY
dBRXuPh8o6wmDaNOfx+LQE2MwWiHYkhYY/YwHNQSUYr/Uo+Hv0txCGp4LBDbsTny
qKE5zmKuCtnyzUJH6iVaX+4TKSqVsUZSpN4hy38idkCJDxihUn1eiNQWc7hKtoFm
9hhgpAOvzVrhqgWwG8qyqeCdLL9UocFxcD0o3de40S8kQUR/svt+jZ+YNz9fOJI2
uIsJx1IaJDTlGK8ZERFIzyub9C0Wgm28Qc648VBuRNtRLCw/jEcSkBb/ydjnL+uy
pO8zPgnlL0JaED4m25vqI5Hvq1NysP+aid61lWoqIz6uvySgHlul9+RXU19Q22y5
3xHi/xqFWwZKG2QEFsprSp2mjs6bWGM2v8UrGCrgJ3RHjP/GX2FlDe4+GywCqkqg
+ymBIXc1G836EdbQlXHrmALKTQUDp1DSReGwEOWdDdMYRlUkGE2XSM++kxvhWtKj
io4C3ju5KEj+ThxMLhhf9PxNG/s/sq+eWFs2acyCcFhxLQN0ZOh0Yy77EJgnncML
KKiSxDp5JmnffpH7Jn1+Ui6j/3nciCxmCRN9z7YycyftS650N4UqyIF00x2lvN2c
UVblZR5meC8rS6h9d3EvmU1/v0rvwEUPC13EQ+69c0G00pRepy4HYDJ+SdSDBiNL
yD9NEqadaDkpmJMEWTS9HN9kviaSGvX3Fd8kmZ6FMd75tHRBYDeiVX2AOFfvxck9
P+P3fgiw1PXcUaD/hheMTcjCXSdHAnA0ZKRCYfRbQ+C0Bdjieqvjw01JrJcL98Su
f17vjdnGzTTssg4g/YmvqVQVqKJ/YiO4o7f820JpmNDb3FKK8ghB3DmBbKrgEKHi
EuHJY5JxVQ93eOR+pU4ox5O47iq9jcEhNnTybLQyWu6g90FD5vlBP598kTUXstxD
dAmbCVkJ/CM0nE/RDyae5qnqlmUmBB/5DpvyoMGmKqOPx5kTR1PucEyZis4Idmum
LFA/6GsF9pYXAmmsgj0zbc1pq0ZCoCKy+6C2gnQJSCX4qm/0JctIfJ0d78vbyrWY
ni4A1Pphu/6bpt9WOg69TqbRRzUWx233mgsxS87U0+TvWPUVYICPCAE3kmvkLygw
zXx3TpHfspuhU66suWl3a9wBLdQSBST9RYjKOpOBo/H8+QDBCcWUBCbHIEG+v2Kc
iP4Rb+ZQHraVGXbNG86vE3ztV3Ifvr9EVVqUh6j/FDfhN3VaTHf0TA1aiYkKfIWX
vMOVt61HKUHiM/oEEtBcwsh0Mqm9j+svyxbuCxLL4uymLISoWDZ7KJU/PoK3yyBu
LIK8btU9UMOTFjbB9soErIVhN+M96lQpvbh4da86Yy3ySCGHtYthlPUYKZprk2hz
w8JOtTWSKOjo7Si3djVKWysaxjPfvP7CzeNoIIyrVD3+ww35nspiV6Gqa6oEdGe9
t4fX7EsiuDk7xFyFHV5yalJVOf7O4jBq/eD2iw3QKD1dvmkqRsV/DUOLWHhS9eMy
AOQtiSmEWgKRvRmBzaZmYQk+42yiyAegZJpPkK+r2WZGJNYHIRBAw/ffSOPQVfN8
A9dfDpGaymsVbA8huRzmpB/mo1MrHouaRC4Vcdenfgh17aDtLfdrtELaJveW5CjB
YLXTCmTMkFGwcbg5qc03zsc1iTab4y2FdyWouheJF8WHDIJTHOaoF95zD4UgV/Vs
q+RfoucVK2qbE3AwuEL8WhA3VrNgqYyiHwRe9GHlMSdXZ+RWqw2/ezJ/M6l4Yryj
2MQukIIsj9OpY8EGW6Kq5tl5o5HH/3YSBBuGFLvobUz2GGzxA1dio0jCqLW12UHD
t90q4mGem6+rFqfoDHgFq+FhKT1k6vui8bPEqBjOx0vSY06LMON96mTQmpzIPMZT
3cPQLHytibZoIzQjl/FXnXsPCwYQz1bWc4fceZBNsuJ5Yy8YLPsdLqYQDZK4ve/P
ZaH3o48AWfH6Ayaz/WqU3LedgcVCZ2BfRKLmJ+7i1ms79AO2XQww7WN/RRgFuXP6
6SFm3svgQPEBmtSbhQsykOl/nejC1gEMO1qDjJ8LJZcR94vGng6fXdG+ya5K+G+K
bibbV97iDw8kkUkSnfDwagaorumgeutEOesmiOv5eWVpyyIrRhsNO+rYlmQeRVLY
zXWWPplmAotaE8EIYbmmeBfWMUdAm6loyAz9dpKn33P59KefuTWhsYp+fpGbGJoS
zBgwj+NI9eMYTpgYPeYWxecuJf8nCuriWjK3Inc3Vujk7tIQe2qTVFgwt1T6I1ho
gDb2+C7bTYi/hhi3jRr4MNp5BvZFvFE0hkBkdKlTi3lWo7GN0IIxbWyOpMGskc5V
/368rDtIERkFhpsVVcaCe85hg84xIUtRXBYCFrnVj31JTTxCH7YaMJc3F9V7wWaA
G0jH/UD8FEFz/SNvoyT1V27by+7lAwU/Uh7U35zR3vcUhS3qsvQ8umudMTtFp3T3
OPNOntUC9tOjBRyEjjpODbPYPJm2aZqytAdajiFcPNVbXwdSlrTYTkqv9fQ8Ndqa
2eBxUmh22QOi8oGO7T/CccQB0fE55hEaODY5RFcRIrp/KFjkRbZtwh8fDKdPaE0u
CAaKKRbvM//CT6eKftRb0/+YN35k3tQCWoSgpmrdXPLa+pqYLfDQ6+t/3SXBFNyi
PHGj4Wgj+CVWn03T7MLeJ1l8lIDUTzHOxZAkU7o6khCOD/pEXUpYP2+aHOdZgs2w
E9H17Ma/6X0hog+f4kD1IGxnltoMiJDKDZdxsbxTUUc0cXO/DgMZ6T/xp1C+VAXR
+M7IoQB7WhNqzkym+hoEME+VX0bx+K3kauQRhSO3fYDlmFzfqgo0tkVysQcM6FMC
0iHn3umeDlTditSVnSk40+4dYXwoHT+TCf0q4tVtN2lsgdZRcgLAlu0rb66Y13jB
/LUUTACSGzv5pK/JEuek3NUhCfOWKEqg0o/ciZAUqsahuxxiDLqnJGD614AySMhs
cF3QNdqIenGgSmCyRJjrp9hGSFyEFI+nLJFbwMADekSk+b0z+1JneAURIAKi70VR
M/E11hL8MyL+Ypz9GFG9yVW8Z38vkPiA2CdzR0KU5CTuarxwsQIO+qWA064OdAPn
OndDusInYLJulTxGxutd+IlEmzkymk55OPDIx1tKixVoBWjUz4SBzv1KrMeJRZCY
RJgmLFh8POWgjhsDW+PVlt3DyP18Avbj6LxxaeRrIEJ+xJLGZJZXeWCan6XBTntM
NvPceaeUrBoBXFBVTgW94yBRxy9Q2Y8jpeE8h13E/jEYJCvYAxzhGKDcl7KJO3ey
Iie1ceVJPC2mr8OeqON4frsLTwgF0RciNx7qzOqyU/TZfrb+9IlD+miJ4TFteYr0
ndloEnazWwGkV0VHqrt/gdwOK30QLOL+2rFjP2f0yN8VVNkQGtW0yH9nJHQnyHee
EeuuwNO6Hl0Qj6VsmrxNwTirvLH9l3e5E2DNNbj+N/fpRTj6J06n4TWbIcsc8S50
gx7gUe0fIov5v5chJ2cq/pwZ9sFsDywHSUh6nWl4gGi5qWm1FFLHfoc/YO1xU1Lw
G8X+KuJYtVNKB3T6nC41eIKlygDJVYd6NzZO54qitJeAVCObfLhfn8QS5ESnLXMr
fY55LQofGpKZVvUS6xOlmB0JCtNvIDfVTkEK9itLI0KMTCUwZhwiUqCnl9oUc2Bo
pGYyjyhhKQfdGBOROYx1Xl6HI2RyRcUpWSArHNwHdT8Lt1q5FZozKmLPvWYq/e0J
gx4E/WWVXWXIgbsASZ4hYakFCrWfq5hGQs6T5Oa2zwQh3pu7yCkhhkFX+07OBvWV
XNyzk9+1KbGhopR4czwDOpzX0f9Dd0jVqssesbSkY4A7Jejw8fSc5ay07748jBtA
hnkgM5skbCm46Eho8XSkAaaqUr1wE0WF0QCYzDDtlVGqqdb49YKmh6zjf+fIoHyV
qsmC66z+QRi9WBr4AqQ4i5jow5ftQ67XMbf7yk7X7llVHB1BLk2rGMHUNA+G4DH0
qZLzm8K9YGBVY3oGI1P0P8imp2B1ga6x5/9SZgbhQB1ndQowc/m7asKkTJbKo7T8
UE+oLKC3eQ0IcXiYGJuFWI/3pdVvBsA0MuqSXAkvwKXVO4777qIHevxWx5WLQEuL
YLKFEKWSkgWaTCZiPTpVmKazzf2Gi8ZoPEeXRN026NxiGB9Hl26CelwT65zkMFxh
htxhBKpOWgPrct60pSVyYxdR92h6HmBrbbvsXjmcrEWPF2e1t6RxwkZI0Co4/M5/
12+K0eDFp0d80bGP69GyaENrefacYESlCzu8jmvWceTI6q2dHqrFaWLQoc0qWJ0B
I1P2vHSm1aqtVJ1Eef5gvy0+Od963FHHSKjHNCAtjhm8p8oM2LGkZmygjBMvPGyo
WfghgrNBokepNpiiXXHJT7PoHTreqfqVZlJdg1xXgEin1hpnYZNwU75sKPnHhHyY
wGEh/ILH9ZTEb0PytBs+meMKwYEWacVX6ch1+afiMlakJ6mVXZjUvc4tFFZA021o
LK+GWMKSxZLXxU3Mh9MfRav0GwuogUutu6ISdk/LTBzLAgNnQ0VZN3O/WOBiPUjh
5h/ImYr610BpB06DSuZBFHla/ax0maj5bnselQhXHUYyMQtjfbRDP6zT5+l4yQmH
OxeoM7Ls6fGZq6fBMJjZ05fpZ4PVnFhnbH326jaSvJ5s2VxqRTb04Eqc1wz9autr
k8Idc8MfKsmzlxOhl6dTfWJHDb/Ag9DU7pnFNVLT/4Bz1QAy1kKTSXoODexNHSNZ
dwQ68V/fRzMZB0D6Lsx2GqpkMjanAkinfGo+YeARZsBf/R1AQYG2+5bgAz2PIbul
Eej3qEBxX6audeRHuQlimgj2HU6f+42pt9rzXYL3CpajD3dNyu3sRhU4vdFv6t9/
DJpeuAFshgqYbPc6AUl0XeoEpWxnH6phM7s/qtL6ue1fqj1kiXQeHEu2JNvJeuB5
gHmpaQ/10m1FgRyXkMB+kn8bcJb0NtNztQLnLavD2y23VRdcUlNtaEQ9LTKKcOJQ
aLLtbKzF9gJUKGnoSigM1fSsBMRWB6D9p9FRGe7C5oSILIFrDAKOXW2WQCc2RbOH
eIzxBgK/V04EjM91wfzZY6b2RYCpnJIg9f+XS3a7g4hKGQEcut2fFNNEZXT0qMN6
XcF7TXzvFszEdHIwcPP0LLJg7z7DXvVuH9NaM3yCcVpEkgoekKGjc/JWFPrEjo/j
7wUXYPiE+OS6QDmrDpi9Q1pt02eoywmWVJQfv6uxdMlJctTF3c50WaG/HSQDUXGP
wvxOxvjpbTZjklyjOQfPWiSThPlVNWJOuOHcvOfh61gS2ssBqYnVEhnzkFUZS/e3
LMS0CTwhF9ChCYlFGBY6Mj/MtMFF20tOLiR3SuuuHatcA31JLX5smysW+gA5t15Q
cvFzHyzJ+3SPGN5ipTbmTaDNBgXRcbJKpIW7ZxDzwcOklld/snMzoGSgisppVEZr
CT8nLxsApUtyGrpwIFicngU6McTd7epu3G7N9vKgWNELN4qly//DUsXl5dVdfii+
Tnh94Aid3fDhN5Aof4/vJoFzS4KNN4uRj30t3d4jOV+OXEzwZ3vpp5BdfAt+ynAb
9MPHzidFZ9FCYWtBsFRCVpG+gvR8rpSqScGzfsRxoslMg7kamwta8CzKCrCwNPV3
9g7ML7II5xH0/iosOvhf/kqYmB1Hd/8SuR5oAjmDLrc5G00Vxgpk21kiyU+pVySd
g33hOAAkxeakHg+w3j3IYK7eS2WvOWmkKlHBR5MbFzNYL6TkgIzRIu95XbLyvxd7
somT9h6bJ9RXngZCLtmUnPUlvjIqklhtw8UJeVf7HjF540vvsw/ztunDH3vfQb9s
fCqa5Mb7E5zTx/A9c2nuR97NUFXTnBeEflHPR/SBK2Jl2NOG3B1xBKbqeq+Mz9St
Jim97y8tbMqQcNgf1rkNTIRXIMSed/rDj3xNq1iU5uhtcXB35j0P+EwlAbaIVnxA
Io9FIyj+bC6lSIfY4mIZMRTY+ZZEDixk7tJrBK4OW9ruvsl0pTKZBfOltUL4bczs
YJw1JSt+6EzH+39DXD0k9UM3trt8crXNc7nEl+/dQtw5tt92o3uy4YoPxT0oAFCj
pZ9Pwm5lLpqda/acRbyHbBXYpyyNqdGXSdVv/wEIeHBZEbMgA2Ca7Xqny1cASx5c
fjPOL2mzjV1FthzodvOcmqpzjGQxhid0hXIzKI8k3+/TqcrzW3y3CzGZwdO8mkn/
kxcfS8ubQO6e1eFpQMU7aenO8e4ztwkXMaBgzxyUSvkAydcnOJYDHqRm1eyCH75B
1Enj3qT+R3H02jbq+Pt16EjXVCf+AkPwABrrALH9drSVpsSQp8aLcgY6FGA/WR9v
CBDmUzVYakKiVo3eyVFWrdGtzOHVA0+FV2fn8OZOuye29gwbPhuSj767bvf6wU6t
w942TzkETdKeFZOG0+y9g5xVWJJGmjWBe/DkCRFAQIyafWKS8UtWw/x73RUmWa3d
cF3OYnesWXlDahjRNdg95IzSVvWWXwCe9EGvxIiD5ZdDlLVdhsbm+6Sz7FubGk9g
vqkXeM7f6p68NztzdtxDqJheSUdZEMA82F7NoD+GgEWaUzqqEzVLCHX2DIlNYD4n
AQbbxIYxSUoNS16rrJnLjGxMPbq1sG28coKilYoipC6Z7Q/WAIoOGlwtyOo/Ndg6
atT4ZwBG09xBF8EGO3+kZPpcThIQNzO9JqbkiygDYIhKusMphcqhGBDWyNS9dEML
SfXMyYCB8uHxBNtDf7aqLXrZK5XKF7jK1MwGbYIkduGDYxID/HOk24aRiURhX4zd
Hm+/e4CqmdRmYtCRCuPbXB2Y3jv592Tf9Go22OXXKjZw0aH4RDdMFUZRlNjBMZgP
wYM6FIYvx8Nk8X34+iKDw3QnTkbYPfK78LJM4x+V3wwcwqiZroRPZq3t+em5lQIS
6Jrby1lH91nWPey27wKIRuDQuSMMgMj88cXQ0Lp7G4pGe3iilvpAgLZsblpgJblA
EBxFov4EwmIoKJ+/Zo37sfXwT7PrAW4OZXPd/cKbefueATzUrj5/p28aORcPjjZl
kfxkZ2elhzcLqgt8sEBbT2F/TZWB6T2FhXgsjYENV2vbnl/5zilm7zpErFC2iSua
XBSnvfbpmTYtS5rc6ywUWoXYw0HUTTW2GZML8U1O5AB6r46GjgO6p3j0gBiA//f/
bvJ4XHQOoZd1ZDuIngpNSWqq+H9F7OuL8EbnNFeM8gBJcie2GcNUohx2SiyzlCc5
AQ4Ams+GD1nXowkgn5zyZFHMR7PLLplJFmHIzacjIPN1korkjpTqfhCIgWvbi5Ok
Spn8/4cYaemDq1qPr1EIKM8mU4Qrhmeuu+RndBtP73m81urYUpIAKC9TnL47B8y2
RiiklHoMk6ognyJ8hC3X6Lqhvq3nILJPPmLPfPCRegpxg/EM9F1vK3B+gBddX3wv
9gdxF5i/7WqngrYf7drxPmiKzk3WOblh2wKTBR5PnOShoyDD7mrgyQUfY16idf+3
wmDaJmAU95PYl2oqN20c672FZKVnHiWOpSLDpoVivcGIeAJKOhAlupf1aZBT+tFq
ctwiMvOhjk1J2bTHXT2k+AlcUFbUKg98K0cMkA+bPDHJS0pki+arP32QXhZxHyV9
LGlGOgKrB67uArI8/F72MR/JSb1bmBj2LdDA1Q9DEOJ45HzFkFjBs6PZUn4uI5N6
sEXejZ5D0/MOaQiib6E+hMPDO4YThpFGfxAg8JwSwKi6++09bdBOch4wZItD4J9G
by4Ql0ItMaINmj+E+E9omOciKG18VSaPy3kSlWwVASMrbKZCBuy9tkTRMCWIIKLP
w9ZVsqI7FoOSeDksA7FgIVRl9g/LO2gw/OIGDqb7wHkr9ZF9FQ9OYFY7w3UMqfCs
Ssgc08axMpim8eoSfNB2Z/d8QVWNkzaLJYOjpdiiC4WvI3fSGiAqQNsHs1LBMrBB
SJ8wsVvL4OcEbCAMtv2/W6kpEPh7PNAaeZteEBqhrLzmLJQty+mcn1f3dtq/tqJ5
DETDV5ZecyTjIuwgCHIRHe4hcwRS48ylpDVMJvMXw0ydc67IHssjxj4z1NjdnryY
IR4Bgyt3DIrneK07zZqoFSn8hYNzQcc6gM8v4PGLsC0g9/ajiS6PkGdXWPfVYcRd
Tk5RNtt9w0BMkBeFafxunXcbp1Frn0hqOcBEbAe/lZzHYkzGnvwRIcCLK0mu3NbH
VaQidT5nQDk4n+zQNeRlIE0Su2Ai+WXy/z+Vgpjyij971hT0FrwKWPV6QhZR8f5M
MIonfHBJxC8TYUKb/SmVEQhHQmdHM/iYxPEAXQ7TRKrH/R36rAt0nZHeVaCyVcVa
02aKKSoCEOJ29AAp/Pl4vjQfbssHeBmKOFE+Gj2T6vim2oEeGLUssfmAGDvchvP6
NejnuGC91QpDfj1h2J2wObC0OQNUjq9+yQ1pBoOYC+/3CPhOqUc/rELsH966iPGo
Us9e6xohg+yLjTM8KRnc/e5zGetqLYBwCxkEy+ZlYxzeHWwyaoSAhPkjR3ZrDapU
hxUN0ycGNn4pXAmFQAmQ5hVuICEJ8Vv09TXwIdErbdRAMrJbepUpQxi+BVpewnpd
+WJkux7x3SWYzpCdKx1GI4Ncq853WzIyU4hmx68xoTMNvlxZ9GQHITRXAlTP7XZz
ZBZ/efE9K7Umx2ICWO9iKMPW6Qu/7FE0IcGUM2MVjaxiLp2NgjhaKtrCxuXn/mte
sjZzJ1ZDFJzyet0e4eE0Sz11+2Lm4Nb+3VXDA/2sKvoFWbgw1DFggL7jX8L6yvr0
Z2C+MULyF/a3+irgft4EWWU0tBh9pbbQtZV60gIrIrV3b3JaE7NNK+ajlXxDSINc
YtvtQvo7jCd5NKMfj0THJRD3m00ev8AhUq4E2NneyV8PdH06HEP1SXdg6POWcVlg
PqLFqBrIWlOI+Y+eMN5Vdlk6LsRBBobt9KJnXoTYRuw53nSCrt8iMcwPBN1VZifi
M/FQSo5/x5vgECcfIU/CSjLvLc6BusqfLRL+++m6n3zwl+qgsXPJy5LYFJwQIB3o
TE0mSZGYP+kS2OKzUGiW3yZtbvrwg6dI7SFRcMK2CixmO9npaL+R1ClXttudNaP6
4NPnbVwoO1G7+OZcPFEkPdiOKXmw1ddMBGzv6/YnRiXgzDNohNtHe2BwGrSxwKgM
H+TZY785BvHEhbHZQcdv/HiPiBomo2UCmO6NdEfJ5b9Ya9ex3pRbwpaKo5ODdXRd
CYty3Z1UfYAkogF+AJ9hdkPb5t5tzMJgAgfk3j+jcemriXP5j6ua/4ZFF5R0PCWA
/EXHjvZXeQqmI4+1YeMqnWQUF1RSWqUYFQEbC7oAKrFZjGrwWBrvmVN9xvoK2fYo
qSFev+e8W3ffRIKRJx34dnTfMXZSUngR7rL6T2J1upxQSnXUUInRCF6e5M6mc8YL
1Zn2SCk8QFwnHf2bFzBdiO9jZU7Izc7KU5SstT7C5WPY7OzN7rl+25UozDQq0SbV
9JUdYMMwv/pDs2pcLYfkQutgK9jA+QeM8LKSx5zwOQevjob/74K26bX/qRG1MDP4
lUIKSOIzt3g8ICbxJV9pF0Ea+kpeS6NS1W4myupdxJpNK48mU2wO6ARCnJeHOBv7
vY/S6uLIKvGGRdVe6zA52F/ninyo8Y3LtNbcFhizQumiv8KbOeoik/Ej2jjfPt9h
4lw3SwIBI+7E5IAc06WIXXhjoY37YBFstNsC/409J8fWMMi68+GNg2lXiB2OZHxM
fgj8npuIDCoi46zRkewJf+HcmETIWqcwa99hYiP0FlMrRisoVMrysGyXrSsHzPg0
0/e+6eJPSl+ynLF+hURwe41aKWjKbFdDadjvgcop6TYPLPzHOzi98n0AFPSYWtc9
Cv04e0DxFE+QA2Siw/nHImPObI8917qJwlW9InC5cM2slY1VsSPQctSPbr/yabIF
eJ2NFvYqV1JHqs9zCw7po/ByTmWOi7CVem9R591KzleaHK1LPHIOAcZjDHznLu0R
lDFU95a5S1L75gIt4oZWLWjVu/X4EG5aptV+DUHSnsb1cLdU3dtNrts47l+UkmST
YK2WQbsX9gC8dYq2o+2ws2VcYy5e3CaeJVkdx/vyIY7jhhNQVYCe90raNWwrv30w
sKoXafywCENShi2jW/QLdjbaJttmiPqKMHTJLYVTLgCiC3ObCnJ5noPaSMDl2xr5
gLRyTPWYXWk5Z4W+RgTyr6VKO+dF8f1XuT93B2kkDmoDZxQsCYB8mCVx1W1FXhaD
lGdRWsbWO585LvKskxn0p82NguIGzA9XhWe/iLDVn8a4DQ3weUCJ+UDLi/PDRm3f
iokbaCswdmNmhAGikC28H7SIjA3aFTg4zQJxB/DCT83PYynDDaLo1cKQrAuNYSZ5
Nltw+BzO6DZoqGvavF7/vVx68EtrX496Cb45Gcd9L1FVTmpl/zkUOV/rGOksJ2fZ
xxtfEP6o2cpGChjUF7ZASy2HK12vOcE59/NoLOnqawBHnYb7Ussn/Da3dsj5Ad77
3ta69i6h2aJEkPV99GZYvE3MvMBRv2gLEVfiShdLOPSnSM8EqAZTq7YDHoFrtgrB
e/WItFWWkRzB8Qdbhui1qGwBS84SZCsfaGrL7pTQy9x3HIU5WTdM0b71hHZY/1zP
kFgPrCblkxgoWlp8nEOpFt7cwRfBQXK4JnOHj926RMvJoiLt72rQeIt9m0q6Zr3A
fGyR0BJzYM3RpwKIQ4m5GR2aIr1DyOmrRW5X4KaLMquKM6onTTpclY3xOVxTCfZN
KXBreOwLGwdhCOkyTPBHp69LstJvgM06ipgvVWpFUSaeLjeM+Q0s7TsLtFSRhMxQ
Hm3mmcA7RoVq1ncuMfYEVs32q6ipGrbURMk8hn+Qe9F6dezyqZgGtplOxWp2ht9E
Y8EWwFV0X1/NWhYn0iKZmJvARtGCIxPMAnJe6gBLAAzB7Kc+KNK1FzZvt1YzgGPZ
Da0xYqs7ttsJ6DM+4fCS1X5gfUEuo53XX0IOGYWUYAa1rHWfqyo6kQ5OcfDBTBE2
TQNP5NmjF9sfFIdKhnoYzFGPfJBDRJga92Ay3GSK2eTHk0zdaQBgUIaIP0WhQVqK
eCsuI/jb02mu9zazADtF7wSj3JnbMk1HTITPazN5Igormux7nfnBcfX2YtTjB4ii
ADaN8Ot+xqPeO0VHpYLhJd+nWoethIilEybceOtar543y/KiDkX7jedobR7mDHpo
OqzcAu21tXrNGmStaaM5v00ajg0Y2FnuTe9Qdwz2mE8Ek1+vFN4GDjy/LgX3Fsgv
FogMVHhIA1qDSWJwMNlV1JO+9y4MH6PvP9/PjIVz03JrU6gScwh5uWB0zFshztBv
FluU0wo0m2854cIi2litMqk+5t4Qcz8736RY1fvP47NKvoTQL2C0z16tZd3e1lmY
bZVjJhblpRcfeAL/auMacdhrWKl+FMINKalAspsKGRyUjdInL4Yen/QEy9C0fSEa
d5XNPauhP76LDLdDohX/zWeSqJ1KkC5Tlntxhmt5Xz+JduDLDGD7E5RmNIbJSpTF
XQ1/rpNTiuITrJKtmmhW8sh1m8jj6ZI4nLTaqkX64mh25uHD+t4B1T8vJHCkJJo0
alNEnhMt1MvaWfnyik0RJ+1g2lhbn5hVzhxsRDv8BL+c49buQnoZy2XEADoWLZ2h
J0FVKf04DOQ3h+i46L5WY62hb9djLcpOl8tjz8XVtaSkZJKpyIM4OlfRGggbBhYU
UIuLBa81la1ImknLoRWyUjOqxGNRfvJS1sRPhTfzKzIsMI8XY/3nkZPCALba4dNE
ZQnJKxGbO18RfandhiCgMXRFEurZbTsSZEkppavd/bQyRyIr8yPT6tOd4tJJNsLS
2dyQgf9f7Z5o6hSOKwtvwKPpBDcDfB5c/GMDdSj+aMGb+SgB97PWBE+iIR8bmMs/
8wmAKDM8UiOqNy3HqnUJ0j2bRqyaZJumaG8uH067Mmrr1I1tb9ShtCTwSpsgtNYA
NuDaB8TOPGvIpF3+g3V9I1astWzpgi89xAQbHflwmXBlJiycARqSRrT2VST+gqre
qYQjyqWPFNw1Rc6Dd7bc/AR1wlEEp3lXyRSmUrMV+fFzo6Yn67Ul3KQfQsRAdv6M
tK/D0Y+8dukJrN9uZ0eLOXCJQZ3n8GtavUOH4DkIU6gS7wBgN+BXcknFlpdUi4k0
6Rp2lTJ64mV8X0kIUNCzxpUl9yU/oFSHA7F3Cv7PxuiqEt3HD5LdL+WsAD8I5o/i
rsALpvcf9+Uvx9JCtwoIFXjuVNH9KrycaWTLW+PvjouF5cOdMAlAKnwNCLV3dNCc
yaS4FuXwS/wnzz1eZXPexfpPDEUjl56dNtintFsDQp9q7EQLYufs1xiT+2HsQwy5
kg3qxYDD6t5RY90ZZSk85PxM9s2ed9+XLF084YwUlv/S4zRm9MsJycyzI2wZKUTv
GBiKbo5HIIH2+tHJ7SFK5UyIWEZuafKV7BIAuBo8HJwhVWDklgRfVGwqI2YoXm8M
Kk+tqhnoDrS3Wh0B0gG3TTnautElfT61bawnoIWqs+6yINjCvDIQgDwNNL3aWtG1
go9qAwd+aX0j4u5ob5lSyHIaIaFtaYW7Ek8hfa2v3qgStc2da5G+LC/msOzzaUwf
PQrDZbx37BGrnn9hrQRIEpqPxE/kku/qAlKvPjy09pU0J8Bi5Jy7s5abmRaIaR/l
cqiE7myFVJvXrHxisE52h5HewgpIj5PtDSVRYWl4NS5MNeaHEOB4QnSDkO0942Tc
s7ri0yjHPjNpUH1Hey7zy2qrQSQFpn2rDSGptv0xKi9j16Ht2Im+N5M0TVGqjvSx
lyZ64iLyTCr/JZbsoz9eQ7igd4ZiJ8JkQRwUK2H5baW2d0PCTyvCQbvcD7PBoZan
rpcIC5NwQuhbJ9CTYnENjnLWkLyMg3WvCwFsUPRRYJFI7EM8g3koClpNCeDUvdm7
S/7dgnYh7o0ZJgb1zyALHnQzX+tEsLusqfNCHXVb4tW63qCjqmxCv9JZOn7CFL0g
m2hp6VTV9fcV/6o5Vo/PbiCjAJOVUmDA914Y8CsJdaW2xjX2KWSxhJ/DLmv9bZ5T
CCiuqU54FfMyjOTvt1oKLiooLuZO8xjLt6qmrXLBlE0SpMF81mifWWYTZigLSajV
O/7wxo++hKgzx6yMdISBYy6zY1lVzw4VajYzpUBovhRWUu3r8xaBUOIAh7lMptPE
VXOlKwgRmkLdB9BLb+f4CYwb4aH0MAGf4h4f4iLM9/7XgiPMKsFa5O9Sex1V5FmK
IqaKfabEg9ClKImNbGkK7cihtrsFeUlOQfg6/ooXw4TvMgGJs0PAozZzsaZ0LYLu
2q7NSi/84svl4OVTrZHC8NUIicw938Jt3onvsq4h32OAp+URtNbvMw7KrVoXz8Tk
g38oRSWIQ9/i8n4+1D9VcwZfmjfYO6d4Ymkl7GPwGjLPxG3/wiUlGo283wO7fZsl
u9+MLo3XEIwD7SUEa4MhrtABCNp35ef8byOf6HooZufo0RxUlRkHZH6Bsb3RHzWG
HG4ukUOZBL0YcPX1FE52i+F7bEPjgk7ccjOIldnZ2gEAbr3caF/krqu/OCedf0I+
RvX4TusbQcuVrUyAgdVc27O0cdMfKenblLW8Zkc6qosYmLnF9Sca1fm245OhQeM+
E+WymBNjOMSK3ouRggaZq1+nVAxbdNwcxuqLPJevTepWL25jWt4AuwYCVOk4iIcB
/Zz73TBXiDi4sqVG7bsJ2CYrvrKJ/jmjvj90zOz6oGWmHbt7+xLv3U2cwbCa4+yD
mvWy9OJxEeRjfeCvuM1SYyo8TUwbZ1AxM4pR8ZOXSL8CiDvzrXGqZ4x/bXetx64d
gdu0xasJm49/20BTP2I+EcjX/I+zPxrP5AbIrxR6rpnPquCy2CLI4zRAcVKhMQn1
UjglNpHW8ZgPEFRl7uina3uFC5arfHXa36Ak1gnk2xJBUINdaD5KzPUbLjkQDjEu
ksuwJ7B6HhQ/7YOGpH9VgGqVzdT364vRjHUYfg4BTA4boK+yF5nQA5PCuR02UnmE
1Pqsxioexh94Ryvl++JMK8XGosuQqfaeBMgt2LyLU82bfZpHEO0tKrKI8pRViQ81
x2ROHAd9B4xsAdnaDvtFCli0eAS6KtNzCzKCAw2S4umc11KwWlMiLOEQTeQEuHG3
IfgXYK8T97MFCiC8JbbleaaHJGJdth0EhXgNh0IpYxtVrwurK1QMpEtCBxZrzfmI
ZVWTl9Tu1/lFntq5AuNDoQyffqCmdmAcaDnqM1ITJY7s3KZyd8Vpla3eASxobTSt
AnUcz2YokRbNXtxq3NK+lYhrKVLnXfzuXFUO3L79xUJqePOJ0lek83jx9KyeTblU
QFYbtHyPTNnfxpz03uX2ZZbIkYlhulo+4UAoMF/RV1oKKK9wYh68aW2/3rZnoB6K
+gVmDOnnI2us30T+UjcmWdHDZ2C3Al6q4VONbNGArLv+iKXecUXD/qQYawaEtY65
oLG3dzLBF+7YN1N79wQZM/ucrXV75aSgRpM0DLUyEZRFLGK3yGv0QZ4OrMUl2Vak
0N4nVquTBGq9MzjKX6LbneuJvww6zN8ShjOQzZPxUPoVAXGvGVjTUcu/kXwI6BmS
6//2tcc0fzSJPjfg8wjJNLtCxz1ktwuKtgzJJhSnw0MwVSaZAloVAIacV59hwmqN
eN3eQDChjLCKVrNcFXJR7815WLu1ofIAdlXtyNqDm4JAdhnFsrActiC3wX/Qmhba
ALFYVsrftKRvvJA6QWXihXMrsyPQ+GFdlX7hp97KGLj9cH6hCJRPyVXeUwC5q0uU
CjFiV7sSPyfYbf4d7yIpiKhoyAMxf6Wxn8UupD6+w/90B4MQ49c63y3oO92jteeG
wZAvzn5bHPMT0lb0vFwg5c0Kb/n/UFKRWGS1dSBkO16bFS6mwsxAGngBPcNKnDkb
kdoEf3tZAp4LRCRhx0x1IJQuagGlIVmoDfYKE//cVWoxrapCFsnZkBgHhSTFe2Jq
q8Hha2Vcb+J+bjuMrNf3yPqX0LxAgoOXRpGh43OWLmo4b5DORA39l0vN4ZqCjJUv
ljIps1NxXfmdcVkSXNJka6C9kIhLpY6k4Cn8L8Jrk9ycE4XkNPpzbNj9gT9c0qiv
wW9TPnD47oQp0o+C8LiL80EgvvIC5bA7lb4Z1w4As6A9lOLllZG0TzNSYAaqojFk
iull48tDzEl9oJFJYptwiDXTLB4cH83nnqYhkGMh6/PDorle1YL2SdvRRoN7vobG
QkskObrc+Wa9X2JOnaVKAYqtyMoO8lXNOv6s7fFMXGY6sY/zw2Kguybt8TnJrqns
ePjjmUNxaxhklUfa3BQsE5lJVsfnm2R6P3aNp2qkYlOzQjHZZs18rHJv0NsOEK1o
w8BLKn2qCjPsBjnt3gpYsTMR5aMfESJCFLg/lhW8TTGJi+aLSevvUPW7CLLyyo/7
9RWf3GS9XVarWJyiuu8qgArrtrVFEzcRG9CC2I89lvf1OulHWu6aL5GlDhgy3QfO
tXkfoWjRbQ45c25dxwMb+uAzR3UoMA7WUEfaMPJAbA+QIlOlHFH/RiKLgMhNW21h
f7QOGq3/IGSb5sgO79j7JzxUIbMGbP5poSp1+VJZ4jXnQk989XplQbGcOQAo5lFv
UIWZmqQc4Qp9GrXVnoSscxtdipPewmKTl3jF0RPTAhFWXQIU2i7+VWGycr9Hhy2Z
4Aa97jRBRNj8r1Amu/e1ajacOWyeihWzEdAoZbOvpj4GbUk8HC69zrZtUlpK0PEd
YefXTS3K0LHu06Pf9O+0/GW3ocT/TEmrk7Kl4R/W9IEYxmmKtLJRpVSFuyxfbk9H
ZoFytlgHMp6GDXc902qLzOkTibJ2+4E0+vlGOlNh+2VMBZiJJ/IZXDaMwFt7HBKq
BFkU68VPjJG90oXgNf7/OYEWKut8ecHtNNTpoVIBjL2v2v6ndIBBf9wmraY6Bj9v
ZDJbXEi97i+WyBTFSacmiG5k4R1xkqxG6UZl3g59F2YGqRZcu9fItNJV/kwNQ9tk
CRFg6gAl3cDKnsfrxEieOZWQmyc7WGJz1+urK3D6Qj86cbzF9ICsjNNd095+Ti6f
53vpusLSc3TryJe8+5pKhSuvaGGW/2ZUG+eUmthwTP086xH/zJ+JDOvf69Ilox8t
AMItDod7AchaaCPxzN+3e9unEEL/3gFHVoqIPOvQzblwGDbIissVv75KW6QuWQc0
XKSa1reXc6bCwwYD081btsUZ22zz07GyvT+8OnscL/TjRrs6BMSF9nmVjunt1j9M
uPmwHRCh2RIS8+5VS8+0E/92pl3YM9JRc3oqYugIQW1+WniRCmhSGITm4dLOV3L0
BV9qhDODYiFIDBFOrHKBSatXr2APW5CiyToc1nqO3+kaX8Qgr9xNKy64TvOggrJV
Q2H+H58u8c2OfdZGZrbBrRjbSoQEBPxTi3XaVZs5ROi1uqKP6ozqp/4i2X9x/iVk
V3a6Faz5NA94zVNfDNAvYzoNrlH42ihBugk70Rux2M+QOwDot3pAKAAPWG6r19rW
nuxEOmhJzjIdwT86Ms9c8+Akal4xmGmt8U0AdYsvoOsxIHD39tnQwzi8Pd+lmloP
kgc/O4G0ji+deKNqvnM3JID4TW4MNYy81JUPzBIPAe8c1HihmugBKs72caL3Qo8E
v2UfINjmZofONM6riqjaJc4V9HwINz+nJy1UlHMnN/KriyXcFeD245BJILtHxnFo
mXePCR5i2W66WdHUS6t7A/an7DlfQ/yLlrp95dwWKqfCRueIejlICrwmZzqmyUAW
S9xsSgApy4dMSWb2QOs+hDiJK1lqONebUoHQX4FkerwVoQqrXX4aVmSSjCzDGgUn
fF8dHdwTZg1YxKCd45vCSOM+MVAlaOdZ3Z99AnsXp/iBeh2U8zaVShnaIr4Gv/k8
cPEBpPQ60MIVcg6R1Dlquh3JGIIBAmKRxNuKTgBZA4w2GNt3BOx/hs4E9ybMKQZ5
pFnaK/53sAffKzBnw2q8YOiACXx55OYEvRV5/ukzfgrq94uupN81/1GxBwDIEPDj
hiox0ZOL1Ic6/nGaEs+pj6DP7zgLmKgOreA04cQKtifJyfOwb9bZ7mDFHHP64uvR
aamSkCfPLGTBUgGl5ZtTzdpuw4LKZWNlHD6oiZORO3bhyMXxcC3g2l49y3f1ukmG
LrJIjVARF6kMYb58+EoYTtoM2hq1QIOPgLL5X83iwSD7KYmHM2DoYlguwHui6OpM
i3VxRyaTDHsmz9XS81q2m9+8cX5V0KeF83qrvvAz+c9YukZJiaTbSwxJpV8irfLT
/GT8qDQ9Fx5G3Bgp/Epk8WmwVmyYlJfvaD7lBUNEGW2Rzacj02TH8ExOEi6f0m8F
Xypx2SJAJ3WtMzKX8lvbFaAe3rYl/jjiHLc9NXthouNZbRF5yObqwM0W0qhxZYAa
GINRRuHj8wR5TFAHm27Tx1aAOpf35qs9zPKg1MdZD4ZzLZG/HKDsI/5ezHSLAxfy
UIjQrYTcHYwu5pDSNvN1xvWT3+Z4sVmYzrIb+7sdbgckdx3YqznA7xuTT2+EhBR2
EVwr5a9+8NrWjPIrBj/+eZR46cmXgWYqbwAyfvRVIRDFeTeJ0vHudVbFXf+s2Sio
vxfDsflhX2pcz+DROU9h4rIrz+jsvGZydf5V5wQH6vEgztukyXIWh+jmrP5vXf6W
ynzn37bpskfvOE782M5AD8eQCFQAvRcFVmSb+HuLuBxLqz9e8XzgTjge2O4udR6+
NpdYnezeuYHwPbnt2vVFM7WDq55ZcQkZYjj/SaYH3IMu6oYqmnmggb1QnFuSBNnB
mYn5ju1VonluPwdyf3ns0e7cs/UKxfhBV8pD9QYHRU9EJUwdf5htKT3QOv/hZ0OW
28BSXXR4Ri+ILFy9WUeAC2ui7V40UJ+ylHib6D4HIPrxWh3nTEQ04aOiVjQ5pqVH
umIeViFbvak/qM0RmaCOiJprBSG+3jcBMmp4DuNuclzG48qkUUwPkJOjX+eFxayV
zkW9WcjTg3BchD3DqcuPNRNR0+PvJNNy8SRg6bqYlOCk7zS73SckepZhQStnu8Ab
xhncSV4MroRGAvfjN/TfEbxM1DT5okQmQZ7bVpwnCu17A+HKMPCA8Q0fMbBT7AhJ
N6uxKEX1x1Ha3v2u1atATyENHRkZxwM9ThGHKvTMow2zEqaAws/J/UKcbluoOeDY
TTkeEuqXt2SCQbj803MtlaAYxGVZAPsKzk/YpDQpIk4lKBHgTDR3Qc7xARZf6eLs
vCi41FSob2RCRBZOdikkJt+KwbfbrZ3g9RWSQ8rLJwmRlOf5waiLE+/NSXPARE9S
y63ocX9ehHtJX7rMDAK7h4CGzY5Ud+KIsUuRk9iqT3IEaI2HbRbxKWg5/9ASTw59
mjldblQEmeNpThlGOYPPlOjMNdwD0efVXdrL9CeQpknDDZi20Ug2iWCrK881X2IJ
jbmH3dsJC/BtQ5FZqY+hwJ3MkM0iz/8qTEpv4fX4ikaxSrC/vIvTJkUo1Gz/Tsnd
GD2EdHCHaSp/WToxSkh3l7N9Xis/HyaCPlmYzIRZgq1VsUiF5uLNALbS3k8o3gfN
keGXJWfyr0TK6O4zaRx9/aY9Guh49CcoyRwMAMLpQvXwv3zfVrVjsQ2BVrC5gUr6
eSHeJdJNYIWBLZp4sw42aupKenJ3GHGizmoZLXUFr1GLKRWMaL12v6wAU13Jgk/t
T571HP+Kq3CeR9U3QYSrjl917z4zNPcXaluvDQ1q0uXSkZJn7HARVDZQNb23+sbj
6YkgZvIz2tx9X0iLEz98hke6Is4GGQeArQPNeq7FMs4UUjTg5rE7I3wt032E4RS2
TyxpovYxTm84ecaPEvjo71HQN+XxOE0FZT7mugZ3kq/Ip4asrnFf5VR+sl3xAogD
Ua9R8nb0MmSNgqLjsEo14+ClYu7PLvujuTwtHrY1+R0+JMEypFy9disaN+B6aWhU
Ic44wkH6Qfk6HoPmvbjxv0R8DLAKqTIdck1QFtx5bf8hqjabfGPPQiFqedDHPh2Q
7ilLMAgHKYupmop3d13S5gJyy47k2Os3hal0UaqKbRXUohi1iFSNoavjk1ODSPs1
ZZfd3LPQQ+jVypwrse2dVNGtURWZSOwvsvRrD1r1AcwGh9sCPa1u/hVU9Gt4RrIn
i5IgoVreK/1PYdz6fe0tGc0ITg1v4qTAXRMDVb0CR6lnz9xrCa2NHGP12/hsPXiH
NakqcnRkYEubHpncDKetHXwhVGPmaO9IUoIDHC7T98rHtLeyy6vUK2wZIJB/ym/2
DVezNv41oatZcJ7FcssnIKq9rs90oNH5rM5XhnDj2QF1eH/lphVyNut0kfjxZNEE
2t5yUPzhH6ksu9YhCWDAUZXt38ptZAAADRCYQ66liUiiA16xtOlLjrzzNVZTwlNI
WF0gCxX37uwSRJkBJqI3C+mXjkP58yy88YCws7u5XOUxA3v4uDF8xOV1vrwdCL49
X2yKO6rRXBK9H++q2v2bF3WZ/0r4mvm3GQczqwsXRlakTJDsS/3/geAWvrnkGrQc
4JKWFqLo26ZaJsgDqrY3cR9jxGbP9Vn9/SbUrHlZ/PGziR7uws30BB5qNL6oq24x
pe/Ys583Xa6Mzw2ZxPkCO7fCQT4bFgsuxpAMq94N3hwSWpWDNghLTKmmxWgvitlk
UpI6uUQUdjPi/2L8NOEn4Y3/M0bXwfuiE4rwQOmr9MUDfMe11oCz8sRsl2zmuGnJ
A+GITXwJIiUj2Y2Zf+HoNGABrZwOxWXwvwpW/bC/S9gKBYcLpS0pEhFljbPQRnu5
5XqpWjbpb5V2pcxIv2w2fyR2aootuNS6jAoaQ8CW6fwbiGgsPuRrErEy8nmLt6uo
EkPBEK0Fq0ZP3ANx2ObTA3FYSXH9L130lYWRiXDFD2hiY5K4dctPvXme35Hz8ElB
S1Z2WopSfCHWh9iT6M0MVLwoLD4PjoN2TZL91sXPWcLbkE5wmI0mH6AnDNczLf5/
1U+9QsYJCU4UgAE5Drm3EuyXUyMX5qsI3G01+AhTNwNVtJETnkxBfrwYx0U/Y8nj
7fxmUIlsH/5M78+XNzE0meWyx4sBRMj0lCQtAS4KkkKt6ZuF637p4mDrbjmdBIzO
5gNVfD8B2qI/fqlfTfZ117cvgvxSG2+x+H2XBhLDceNByOFssE0eMSr5UC72H9sT
QokQnbdLfXhY+RhpmvfRUnOq3yL9oQ7VKdw6215Dse2JmzHcg9c3v7xVRCQ88i9K
F0bKLV+k5wKB9ernP320pjEKoBjdrQRPeSF7reertf20yigwpMU0pASAY1y1Pvne
JaoTH86p6Y8lmZXJ90++xrtUxX1FoQU5mhFE7Y+rhhunPbVOlHcIj/ahPUq9QsAK
Dt/l6c8gh5Uvp8Da94wyFWRb73jcROoixIO0sDD1WDfu0TP41+x0YWz+k9xQZIFO
NM+sDbM1CY76+Llus9LfcWFDRNLC04IHK7LtDVXJx6XPCt6oUttp832rd/2XC589
JWmJo+BNd8C/6hpyjj1Sa526iOSeUL2+cQBLsyZkp7wNv2yVByOPdij+UH/JsiRm
44sJzByUyIRT/bZXbicXMl/pIwnJRP6s10wKo8X6lfiISN/xwxVoVrNzzLqTJ9gw
KVkghRVKlZ0WtH8qbTU2a/++V2Ku9YB8UbIygaAzOCBox4G83EtuMCWOqQ9Su99s
OCMK/dvaXWNj0iaY82KuzNoTyXvWg/qmHgs0rAYi29ot9ZK9MJK+3AUfXr6k97kB
x9VyGG/0f2fmQ4tyQmgCPzuRXjkNsJK9FU04wgWq5zqtyrCM1wcJoPlv9319jdBA
5r1ZSNLxdmGAcrM8zVMiYfvI4idH6Qs/Y0fOV0Bo33MO82oqzkA/6A3WLZV4lUpU
yhY8NheO/TtnDgNfhT4bk7kPxiALgzNQ9jUKoANlDeo2OycLxGGaBVyNTGOoE4fP
zI5seBPkUYXWJoSwa8gx0POXccMYGMfqbksOXcu2gixO3yd0NudW4wJlFtTJVTst
+IIXNr+urWiWUXDAzvUf01N71j2VpUh72isC9og4U9sN1oh6U/zQBScJfDbqXWoG
Mx/1CppilOA5WNqJEF07Y89waAkMlYSjGfMEyCVpxNRZZ2hO1tS1PC4UzCu7KHHH
SUw11AdqVSi/1fCtPLrxSgl6wl1ndliphkF6OwmkNTCTQX/Z6oYLzgMDg/S7EKF6
P6bfpHbj1jsVf2HsGm7MGiy5srK9dY0FHBmNXdnIW/5QbUUIxRXnJ3HBttFnNTcO
VLdwRSXVv71DL26i4gySSpyzDQxbBtvyEKnQE7jPA7DAH1EyY+pEPpfpfygIUjj9
gtf6BHFehDWdywGgsuN1TOcRG0pLX4GH1mASvaQ+e6DtuMzwkMwVMsKhK4y1ZBMu
W6eX5WmKCiFtQfDS3Vm9wi5I92AhVGkJA1z+8ew91VaRGg8HCIaWZXAcV4Tk5l9N
VdJgLUnqJaQt0OxiKbqq9ll7CD6vkJR1t47mWyielD60q3YwfydvEg0MSGNI3WDL
G4s90zpzyrEUG1RRope6HcZtT79kdt7+gHJcortwDG+4UMKExjuMYSxTb0sbD9vM
L5ue3TbTUUBnbLi4Z8sfl4eQ+TzNicsV0G2ZxHTE1N6G0c3+Kx8AJYl2UpdcAXiR
WInosA1URrDgaJ1HPo7UeiO99u26T5N3b+L18UU+SnQcxJxV8kgag7sVA+jCr5E4
pyKjhGitR8TRaSFHVuy3XgJlT+JsBhv2DQ9RUIPGsmRbpO1Vyl7TfH9FLIpb/03Z
RrAwL1zcwWSre7IVEjxJfQJbWh71rp0k1QoGJgktlT3ww/A7D2mYzIKvKYmSfIxF
V3/CW2CXj00czZ7czH2cMkbh8EUxUI8E76zUIwWSq3wslwvZX08sKwzOXShn6Wdw
hBdY2w8RXKfjPy1F8d/02nK99GmwbOo6k/Fgk5b903fXO+2lP48/UXyjlxA+FKZ1
JXBdS2VPCwHcQznd8dIt4KWgWz4VJyWdVyDpohh6aepHLZdod8xVQiauFHnqZKLC
Y0VaRu74G1q8nNOjX+namGeLfvBX6KRYxm5GNElV7Ky7HNbgIdbqaVoj+AOIBv5w
R65u5n/dQKN9DVR1MgTWJwjPMdr+U/RKKdHD9ptHyHzv00J3NtdIv6lkwGsK1QWX
SvHqgbQURv+R/UHWrh4fTsHmLb0P106ZFJw+2WJeVKDuizF/vJkOPdohMFNqQsxt
wGPR7miUxLfVZMoXVntF7vzvrpdcc6DrpCQhD2Q7bonv82+sWhb0H1zuTeK7H9z8
DsNIsJcVhcWCOnmUh5UfAa6+AUiTlVC3k3MvcGFIWOlqEwSA9s594Ko8IA2nv2Ew
LnS1ef8TS5UT3C7EdM01j53gusX/vfw0qHu/3IggUeOVk2lSagqpsD18bQhaKfii
8E3mR7b0wySFdywLznaIJtdY+aVKofPZZ9FkR9i+hDBIj9cF1F2OdCsMMxx4mruZ
Tu214WruWfDKWFzZq1NJCmVlxw7OAjuFcK8CaQzihN2KDnnqhOELdOy4EKlJ/FcV
/LTH/aajlH8A2vCtFRWnY+ezNlXT/XvPlkcT1GK77Vp4UMZyVx+U+1e4S7OtU+mY
AOAAdknbvGq/6ktgbdbY73cnTpXOLjKKkOQFWGhrlYLoJ4iEdDcll7T0tgNTC14j
IZfXPmx+osEcb7R+V4U7IKV/q3HOEaU7e013/mWWtQm3FU4DHbEu/WNlNQKWO192
Z4BULFksFVnq/hDezHmxVHQvYqs9eSl2CI0UBeVLMlImRvVHofU+5Cq+BttRkRSn
0LWNtDzws+lolCcYGPlHXMjqbCpEFC81VVCAJxWUM0mDXi0gwRGPhEwRCi7GCSeW
V/ujWLpgXkg6MWU5Bmv3zZ7gfvhYpDrPd9vPlTXCF+1XRMOhhgdWg/5cyWpQfSoP
bIfu9MEi8uFLh7D2a13yceUBin93ZCj4WT7LPccyrbEFltdS5WWZXTH9P7v9zL/H
L380WgFd7LO/iRNU1irtr97rNMwLX5qmhzGTKO+92UxNbaxHKgNOqwsCN4S/nmra
SIdMYvPaHciCAGK9/n1TEWYW3fkld/GQDzPsKCt2363FByivk1kg8LNxDPokTb2O
9+ZAX8FdzBzb06/SZYAqiZLCjddi3853PKEeudsgTucpdTU+6BT7MqfgZ3bRhWbA
ECZ5v2gpnV9sn8jqleMk6KGnGvQVUkSzfmFx831zBhu74WrewRSb+ywoiGhiVlJs
TOHqBqlizChrc1nh2KlC4b+KJNkcBEuMeRCEwZXWNlDpddQPhP1WmpB1Qz2ZVwqW
HRHn3s3CEK38H0YjCFvpu4F9Pvs5bqSPWt8bnAZLK6qy1VkwJIprUQcrWn40fZsI
qEsjMM6xvhuSe75zDFT4xOHITWbjiLWBR/xUn5v6Mj3Lu5Uuef/vy/Yq5Hcafq3M
5hPrTMIWYqpK50mi3KkNaW5lSIskb2opusZcKX/V7cIMPdz0JDLHErIoCBi12tuH
tLnHZRihU9EKPzNT4Na+/Hdtrr+7Lvz0f1ZRfCHM1++DRajnzrEXWwexmvz+Lxsz
DoF4vGZoDk2tTGStNUbE5F9cRsFYTCEuZYNn7ctqwvLYWQwOmgZ11Q77+rl43qOp
+OuvBRdCegucE2eMGxU/P++zXCR9pbyj2G4lnvnkQOnhfSb1tUTQEDRXTMn+vfIz
Aom1jaUc96jGP1Uk8vN9+WCTnW+6pXir3oiXVs4eevVql7vg81jzcTrZyp6hl2su
zVbjMmuzthCHEcW+crLdoMT5TKctkyl/ae/wpJOJ9mQRnZeEoo8F+6NeoL/A1R5l
38K09dvi8bxddEytszGW3QEBZNVrVv2b+i7w6OzIT9aA50Csv1xxjt8oKg32/U9+
MMvK5Dq9dfgQyxBBtmKJvKtqhUeir1PAUW/dp5bWC1guQ2qg/4JL9t0HCU3ly2JK
cgjcR6l9SmkqG7Wqem8XWHh/a6mtUYArzsjSReepilpwtleeAbC82k3koJ+aAC15
C8c5p71fzIIifuWLXgYOAsW5a1KQBjPhPyJjDb/dHrMMExeW5LBRWu19YXZYxbfH
rXVadw76Hasx/Lfsc1/EmkqS4Pt2jRr7xQ+MZybOBg7Ga6+Hvvwfg5SIDWT6abVo
6veh8n3on/wUen+QmqYjU0RNikIlSnNDwfNo59NtkYqjLd6kTcPk054ceEj0mS+H
9UIyOmi6wogXGD3GPjHlQtD/nTNbqEl4/mY6+6kUEP8zIMQCPBol8LY2S+YNqKhX
1YqUIPCdocqDMTpWiypP84JZb5TKNe9odpMF/yLlyjaZrcJbEShGNXeUHA9qEBt7
Qqh66Qy8x2RqlfrlTirD/0s/y5omgNsTng3of971WfUpIzS96cRoRLlFBNDpBTia
e5RanJRtnXPbHGAWBjfsdXSZDEb21HF+ftNPzUSzWLVCziXD6ivSM9SCUzs0qSYP
ugmCXpes/4ponFdGzJT984hB4t3dOirkKqfI0BerpT2T6AJV5S3woOQcr77o/vdc
nu3Pc2ahyxnkOuBTmWv9BPNzl2flzgCYaxzFZwAooSM8xD2UpzmBZSLFPHPx8sAB
uCT78F5RIMXpuuMHs5nEj+1JE5vGTJZqGxhvJ1sAwaDrQpWZkHM1VpKKm+vuqJUj
IcrMyKtrp8lS4dOlIbHlIQhwVNk7S3X0wJwVauC0JI3SjYBPGVH6BRYN0gL6aq3w
HejqRAy5piyHROPf7nvNuaJAafBYJcaifEwk/ZE/80vX6A17gFH/8Yi0+NnMfQ+m
PLl3qZbcs7xiq9tfG1v52zI4mELGjsiWa4zVXKcJ/XzUUfzDGenHOR0S+DB33fKB
WF4CH8f2+O5aWzXOJn7/8SXlJz3LAQ0t+TyKQgoSfjN2f7XRwKHiWDd2FHvVJYWx
15wNLbgAEo0Ba1mPnBvYhbxXNbWGOiVR5EOKNqA1rVEWgfaoqRsTiAKgBfBFNp5K
0I6zY9jsCLsPipGriiiu6+FQHHH4uWFF4DjEasS1RxMB/5I0Oe21Pq6k9OvO81DO
dVqUCgv7vNSwygzSkGqzfLg+6X1VPadDGBvZ07VtIbtOGmM44f9QhvtUZgw2P6Iu
geVwynL8hLSugVA/K70EBIBiJastXtsUOzl21/W+ZY/gbDNhyC6HJfVNuUL3hGSM
8LQxTbCAABhBmxFYHERYZy1e7/e+AZxPZg57VJ5JJCHloP91DfGwqHy4BJOB5wwA
t8iIK61wGAg/Esma7ft8wO+z0Eesv46TX4SCHpNrZPpGZlXB/3G25yWueMwRsU9l
GTeYnY+iYmXGCHPPitZDbguEjKWxygwG6Sf+SPriEYthMNoqRqNhGqWdHHHCCZ8S
6Z6Y0PJkL1tQW1nYLl9WdzMuuioZ8Sh30pyEidyAWIb6tvB6YA26GIyqFBM7OwuP
m2pCOQ9wbrS0BZJG6FCPY++KcxLmm3Hhmll5vJ8xne6MJPP+mVtgIIdD3X4ikh+J
E128etJDtmJrrT4DCHwmTuAZmlrSbOxSzRGu3iJ1HzZ7I9jrAJHZ81Pd+a4yxQ/t
OX4dibydjsh5ZgRoEMygdnqgA2ZmO2Sk6jkHtXUvSZzCJ6uzOmH7HCydeggvDjGx
6tGHyTWzgoGEYDgXVi7XLZaDQBgpJINEYmMPMcXr8CBAN0PXUd+XdLRk4ZzKd7pB
XqJhUKGCxv6su/ohUDuaQVVL+n/6QWOyn27dJtRbblpy4tVP0Id/L93U+kZ4q5qH
d1cQPlM8t4pdxoFYEiw5N5CSXJt+MBMYqr2tYhLetQZYD0KRbRrK9EEsEaAL5jLh
rqFrMxEZwM7jpDSb9s37U9cOvSZbl9zsmCeaRpI2Lh0hyIJHmHHf7aLhK2Xvv+3C
higPXDPcARlguVOwd+loXSmdmlsDPRhfN0nnldpZNRw0lZK8rbf+DUFjFPZ4vCm6
MKd03kaoOMpPMRkMbkAOjT0rECVntCx8Vi6YXszNLB1nKGoseS2HlBwoEcAfpFE8
E/mKzbiVbPAjzh69Ph1lFW2zmnokVt40PD12DLX3WEPMP8IU9ZntztngrSu0m6VL
u05OY2ghWLBovRkGh6X1Fn2+sPYyVjnrkldutc5o2gFDEBjIiNAemTUcrv7iq6bS
wBjpRtaK0X/OtonYIMLdR5ZC/ofECVio6QRhWLry6voUjPGvTuW9IgJPg4P5eZML
MIZVuQ7AyHhf94DKwMLzTiZjX0lbFUw8Qcf94K1Ti9iv86qlfGD6/iq2J9DfrGyz
DreD5/HP18DsdqFwkPZjYgARDof3Am8mlBfR8yGwxdbd2poFkOTBHNOigyJ7Fr53
NR8xEkR+KI7Jx9ntTr+fjiAkOWPygGMk5rUKDkBIpHJKcCOqiyvr5nMGEf+DBpNI
7X8iNWkg8UacfO3vq8V3P1ag4f2z+W54sTUUyDaGlhVncG5jZ/hGy4r6w5H8FvME
W86Xdc/ir20sdW7zjb2FzEaBvA88f87vATmQXoULHFJOoDCmGFXmX9gG2Wt9z1bG
vE/sOEgnU7MsQAb2mr8vBudn3Mat8rzr0kQJfllbLqbardaFFx/C0XWSkdSbahp+
BHlMfuqoyX1GJUBbY9VUdRVIiydVyVoo93lHe7fmr379oNlH4MsmdFrdfOLR8b3X
mVmlVMZxJc58UuyPUqBySpzoEa8oyJ3eqYdBLBMSkNYzy9y9EejgTBuKbvY4vfKm
Z16L8axyGuaGlinshgsrCAYS/MMX9G2PoQl/ne0CsA6mb8JJBbfFCStVOE3ckPb7
pp0cokqpey6aao0Zw1o1GhBqvc7rkXZ6pMXUEA1XlBuzKw9GRned+7VOqI2hFrUa
fP+ha3SkZ5T9JyfF0UMZUrBQpee7zyzmxyU/Ti3MnMUobP/lLVreMN5ZQ5lDmM83
qGe6Z6so76eOPMOlgv/XlMFBsTj9QiM7tP6e830qQyE0LDIBoQub4IpFsuC9sgdi
d5eNmVgnAsvkWNOMPvRe+xkfvo5LMGMD2P2g0x+kEhPUqc1GOQ+ejH4hXgZzk+zw
UdTUGai+CX574n39N1R5uTYYScNJawKBoxX0jWzgb3iXURt0BfxXkv5+KdIJHt0w
99I7ya8fBSIrEpMWpMyOMJIteaGhf5q94OVcaDlQT3xWihwYqzNNoF6VYiSA9Fy+
Ea2vHBf12czZRoUqAcxu1Q6dhN8TC+LnRwk24EKHrKIUm6FBKF1BMIg/Abv2ExDK
ThnMnZOMfydZw3xpNTDYoef2U8wmLR3lzfq7UgKLM7FssS2y1b3tUAFvECLK1lIH
amdozU75I4LVcZgDjy5Ct6B7jHJB9ZlLbEF1+SDcmfL8pMaPrg6mweii84cidm94
5IizxqPkemEhGkhY1joNliVPi38j0kraqWrUx+DjPHiw9nTwOSI6MV7ph6rq133j
l+MCT0GMMfzS1/jiqdSaPqLY0TIR3MGAg1qREWv/z1CYgUVuIRuTiJ07LGCSBCvr
nB/qnkhSLE1AGfXrW9JwsrTuwrCOuHRgmJ3CBfdLYgCdg7ODa+f7bo/l20XAHj2N
7XoBlP4HNvRfkW2qqa2J+xU60qqmDKPkx64xZQu5n2NZxrQ2Kf7WJJFnoXVS2b+G
3fGbgqMcPnKarkA8MgOosMpbGn3rp6uiBXLzMR9kVewjuqb4XpkI0Niu5+6Z7bXP
n1RWj7Vl91O5ubYAp4p2s3HQr2vhRji3Iw9Cfa7rIb7iLvlcQc8xv84e0EvrvuQc
X9etyDAsuKGPow+gHq9yHeJ8BOQbyNrDCWibDSFDZwtCkqCFh2+8/lurbFIPbFuq
ra16Z/WiDYy+VBEnCm49LEeeVZ0DH46jdoWRpKfpFb/9ogYzcUISaPTn1tkXcy6B
UVdWhgkv8gesIHMLes+rtv2ToKuTNSIVIGqSSN+TqeYLvfJMxT7bTky36zywcEvF
xWJKVuUL1N8ckeFI54jYxPs1osYGKqNXxI7iyEmtmMa0ORXNDdT9jQ0lGklD8sja
/XnH9fBzKJdPDc90/6j1PNcTg0Qq88XG8sRljImpOt7bxMaWaV33HGCxVhS03i6q
95IJxFkE1xdvuTdHe9PTRdv5S8Tt5mb5E55Y0W+QlTSMZEGX/+ahxQCIrtHY7Sn/
Ea3h3uYlDxCEzxwhzaU16ncsJiSSedvdzhDfVRt+OAMTyFXE4BfvWyixdorFyPRE
uMddFjFh/rmqRtdcsdn4hRkfhZ5K0StQzxUft1hMICyA7UEE4zgqGFDfzicRDPwe
5DGRfGCAfEe09QzGy6DfOqMbE8ia/3Fsim0bPd/X696e+b3rATrtS537TmnMi8lg
H6gqzndpCIqrxi1wcxuGmBpbMYXjHwXIOygnbYOx9W20uudZ4We2sQKxGMbBqh+G
ZW+b6S76efy1uchJtlL7RBv2Ko3vu4iRmoK6xuzHU2CS70JS1luzB5W7lsNr+KOU
EaF+px7Us8d0+NQYDDFM3ShQC8Xq5IYR31oLbxcCIvSxRY8ZFu8fSBar4ZdaFI+T
3RX4E91Kon1gJn73g3rozf+350r4B8bLuAMDY+arTg8QjfCf7FNTAmg/H5m9nHQh
trEEViypYS+6WWYs9HHLMc0iZClaf8I1VPWS7yUoFYu21LJfRKclrD+FUGiPyiG7
VgpAuhmLIVHEvBG5kmlrjUmflpHFjlq91zU9pgOHXBrz5R+3KUxNO1XE/XKltWNO
fGqLq+6dgxjQU/3sp+7VXokW63sq+Qtg0RTd3m+XwyzoFGPQ1xSPyIBnUgei+Bd6
ykhTApshoYuigQp/meyV2REHLeyVVeihvO5aIg8vwLyDgFR02H69MNgLVK3ZMPEb
Cq+qoEZGNKs9CGqrPD/ouy85ayA52tnqUVsEyNpjRfHIczwPOW5uzU4/SCS00lIc
hEsHcOeb+yHHlYTyK6BBoisoWelck5RFpfVp2c2Pw+CvufkMGcTJuK1u8YPUFvFh
6vmJsvCNhAkWVdB94+ZpfiGIam4DWt2lB5tHq/9YEKG0WP9/ei2ObqSqYE4hovmR
tVpxRmQAc0/05qcCl5y47YafObRu1MzLq15o6M9twJloSBJPKsx/lkpLfWvVXUyX
IqiA1BM/RtL9WaF4zF03pVGfvqD32Orv7VQ8sWwoCkWFuDDKdT/Q1UiudbJmQgEQ
8RDjxrposP4UBBXy2I4zdRURwzxMNCK7BD0udYdYXO/GlFNQkfcQoAs1rVCgfOnP
TfN/5M/b3ej9KcihPIwxX8D9g73Vby8hAo+Uj8jnDaUESFDawHkTmYBu2VO0bNDZ
YP0ipycdhnBOpHyAh02SIvvGtKHk658YWwoIeCC2uDaS/OGVpgNA/mG3XMDRc+k5
S72/xniP/BShLNz55L3DIQCucviESMD+lOUirWoEpJqXOYILl2GCPFk54MhqhV6a
u5M9EVyF0peZnYDKQm2aXu9eVU2cpjPttn2XACP8i3GfWtyOLF/ISPT2HF2UQBbL
U6jxWqQRUxLjZ8RCpcYqdKHIgWZycnODxjbJqI/98U38DssmUsLEfAyp/mTlzYwd
MQifg5S15NKNLjqbMxHqeHnlBQzX5bC0bV2umqML7SythRmj1EDokrad6qU2NE9Z
b7E8yVH2zdQnphFyrlraOnZ+c8zi0wN4LD+yx0iwM0JsoZhCc3fQWmJN1XRmaNUQ
KjWNoPY4DvXa6T0y1lN3ryS3gdBv4rZXkUzjBae8gs/PZFkyIlk5CoPuMY9qMnZq
fgCJwn0OYlAX7tffn1ckhnvEpvmKiXCEoYfWDqvYD9vWeycsMJ3wMfot5pEnOP8F
lM8JRfoFFnXpgr7eN2XKDe1aPhJut635tF/OVO++zY6LmZZUBned9t9fMXaYP2RP
qJ5IYrpL3j7jS22ag3ro+gy2HlF60W+VKSfHT5cGx3UkWTfg+vtnbL78eLvyQHX8
eZ2dcaC1bisiPESkJlp0BGi7UlIo/UFC66rtCDH6KqNnqYUYlzyxtlEeYAyRwiVY
c5jifsNStP/1zPuipRi8viz+BpwDCnSpUcagOfVIYnzA0znphsKLyJ02FxAnvwWc
Dsf8hT0SEQHKrjrjkGBMG5Be/ElAZlT61m/bPmUFSJlNliz7wbmRFohCtsdOAloB
jhJ5LxdLnHAyCyV11TRIBwEvJXkxK+7duepI91NuB9jG1QF5hwRlMZxuuEnIRM7K
n5RJPRElNoEeX66th96rcp7/bcEu8VT8aAy4yxxQ0+HbIvHG/Ysx2UYt5LBusPiu
Pnz1hdakxI5SnNguqkgkQ8zhtPjLWK+gqPqv3Pxc3zXYMaBzmRgLi4XlZufi7Hxq
CNy+ycyuI5SKj4oTGCeO89vAB91QiIRGN72IJE2+WmX+8Z5HPsMXnKpUh0PUKCwL
M42XLMTIpm+cpGAtHVEXLksk5mavoSd1fzKrRhGfKS0aCiQEaMhI8gpCI+xRLbIO
abZ3If8DAHzprUphuJSODs1yk2HFT7FzpmXZNGz5nlcLRG4bbeBd47Znj+TXRQ2/
E7PusLKIRkh/NwpeZLShYRlTyhqF6bOvCD2/dZ9TzdZErjqQprp0A90xfTdWYcLl
oqOz5+1sD4X8/C5nlFY4D07Fvuhz7y7+F99qnrHHJCm4+cdj683sFXVIW34J92yX
6qq3iGNNNw2xxu9yB0OBWofHc6F+45WV6drA93zbhNRdHxHSPhmZkqw1u98GTdWH
o1kFSkizLDa7ExcWRj4Ckw5o8VtCLQj8nOSCont01AZyUuW5VPAcD2wNMUM3x/So
tJvxeq/GfFW0wmds6u4whQ3wJKVZjvFMywj30+4ek7U8/N+2wyUQHGMpgtAmJMig
8Ebahp4BkiCbN9EJpo2DYXK1LBWUUjKbxREJMbqqkNdodrA71IwoMYMlAzawkPLu
tQTkCccBIypQjFz56XyH+K2Mg6rxvLI3X9z4IJAwsmV83oiBFYRYYENHtnsSiwU6
Sb6Kljrulw4aYl94ZkVtnvFrtBGmbY5HhP7gMmAb0Yyuv6L/WgP1F2veUqB4njxb
Eg7FaGRS3wTK77qRDTJiLAwQ9VXB2PtKsgvt6Aa1fSIIGulhf6sdjcG27BlP/MQT
LRSRLDWqtZPaTPxxE16nDyJ5we29kpftvosRGQhoyNs8deGboo5J0E+wC94yacjt
1oZCJh8XXycN9pqKUjMHR+Z1SAy6r8D6i4jjcBsudJQjhYfk2w9KMSSD2fcuvh24
GGkBJz3J/h0/z1Q9EmI6tLplupZNJftG14eT6v1yLoxPZErP3kqBU6bxKGXYNA93
bVoPRzu2UyqK6hLHjgiH5I9HPj7kFPgQNfZqj6Lf1ihxFbR6ocs/xDWGJWDm6HZ1
2Fy7ODxzi5CZdCTYW/WmWclTpHrE175C/ezMdPT5gHjUIyn1ejVFMkLAVZIF4ry6
Qf1VqpIUDytpNVrOXLe3N3Id5Bs8HWyD59CkeeDFI7GEEcnQx4F1rbpMM/OWP/tp
ULZgFnJTvqZquPdRJW+bjzM+l95iuIJILNXn+ldRHCI6MqS7b6kk5fPICUCE0Zb0
9J09PEuBaqzHYnDE3lL0QIOJ15HjSdLlWl269PdzBFepnvme2ReIp8zeRBTcjECz
YA9vlQ7ejJDLDSe0nUjV6qN6Kq8phtnGa1Ekw5pLTakTHQzbpAF/mhAu5NGx1B5J
jzKbS8TZC18aFrYG83SYL+pcumySfT1SyWClkEOk2Qfga0fLKxN7WoqxPl2Tlfew
f+zGGHkBb/2KA1jgSZW8tYM6TwUpn5pD9YeCjjFzgiVDVglVE7U+m8xWaUHUS6lC
28MwhizfNSS29XexXHCiXwiXw2wxrfwTyDMtmOx+LosGULo/tZfbOJ1S6ixw4xpX
QQy5LpVKN+rc6BBqzj7iPQDlB7iBIjSsqwDIfw+nGCQO030giC5adt5r2nNHfIzh
SHFt2phNyBqYZZ/ukUACUiJKexn32OC1M36+ePcFPl2/YHzjsRb+R+rPqJuCJ33v
ENetiJVJII5klXMbirmHWWuERBnQnEUj0CUWbfS2cwIL6r/8UuTKGrCx77LcrOEc
u5HUuD7y1M7hon/6U34Fy8lO29B2QBANRvuquC3AGi+2i1Au8wyPStDz8gxFJuiP
z2pF+24vyVyGIS8Zbbr/gi2Z7ybiR54WA1zzT6/i7Cr5+/e9RE86UW2czPONnAn3
PJuoUxWMLr+9IZN8Vm9Um6noOsnHWSaMFtzGFjjn81zltw6y4KozH+gKSbefM3mC
SsHhTFsoWT9m3mM7Kdkw824X+TG6qzTIan16zcwlnObaEgrOQ68a2gwCdV5g0aYg
rC1QqKXWgWlwhX4sa2fBiygu/u43jtaS6/QyOupx15pFxG7OcLZa0vGA+vayxdcF
qENFZlm4Ouw+PBT3AvkyCsWR2M0QyFsUyXBBidl96i5q+xOzQ9at+0Shcv0lVb0S
miMcFeOtCTqsDrwV3P+eyDs7izC6wwbBa7yopUcilzK8VjaKUnAJ4IlwdXjVjzMA
kf7qB5Lp1AEmhaDnE2oi/5uSb+e47XUkrYsnBnGbSIlqx4qMCWvNR0AfsSUkMHRz
xPGWox7IsBSuaYo+q5r+WR71hwAc9vn1o4veJ4LQQ3BOauBkkzXMdyMLnqABPUbo
QTMiYXCaH0T39wpY3ySxYUT2ZS25XRuMeh90JLXT0faX+/zLMtRBxx83h5nl5V61
4/oo1OuAH5/jzFEdGqKnMpfVrqZ8kgVzT89jbstYmpzIkhKPldq9DwOhpcGJetiK
5wJoq0q4LQdffl7EYRh159BDBOjOhv76cj2jyPI76nOzXpQr+kSzS8bH/umIg/Bw
G7Fht8MU+mpGJBD+2zsIeTt0ngUpCWbzkhKKepAeV7kMstzHLtfV5sYwdnX49yIX
6e45ElgnKy0oGjsJgFwxkAAZnObjHQoRqu0RWQpYgBC/AezxI1BuHIa41rs0sf0Z
vbGBo4S0m9T6WGm1hfAltePFjJiQPuuRsglWwkA3ApE1IwGSGAEBcBYHXKoQYj2M
Eq68ViZGI9BAr86Tfk4e2U2wYVjml8i4lXXOuvDQG8/Zf4vN81pYrfHLZz5ZwuN5
My7NXmY6iX4v/9pJ39X0gpENYyipKbCnUftO7BPhrCTi0bUQz4k7FnIP18C343CV
FO+eqdrG1u6NTG5ZB85IwJbcZO62nf+dlNl7bYMp+pIoMTMPwlQVzd5Ih+UILdx0
LU7FRlgjKBakIJ3D/HZ/gcZWdY46WLc2mjk606QvIbtDAFuKtXRr5DkRPn9JvfOy
Tc+56z8lupbDGczKjeKcHwhOxHyUEratQFmCK/ZOLQfKEoA6C+JabztvyfiTppZD
+VOSrFn+qSSaM3OOXNTZ21v47O/pJn7+rXNXMG3VUuwjPrtCFNFvzlH6MEc1AlgC
CswMWoRmU/d/WYnT3FtJl/HykHi/dn6E2Vij++pdgavfb9M6gvCtHQnZGkU3Chcf
4yrnhg+OGQzV+jZFYcXxZIQJmrbPjHYpljVDod8phwxV+P/1hJSwPdpT+t2bbdx+
gBYxJ7rNbGnuS73Hw0qQLMLTe9DdlYEpwuByrrLRYPc8/n+/9S9t7/NfqG+Z5GHT
zvC/Yv566MP9bXSepJMOqQswtpXnPNxO4dlpDnh59mRifuDKP+M3r59qWT9OilQ7
O9Vj/UKL5Qt2IJ2wV7B9djZRAHGrNWtSgRF7Df4yaMfJa9WOMYQN2UhJ8g7RzGGn
VXX4oXxUa2Do4jCIZo5eJPHyjMTopE0PWHTpYiDx1lYPCHDAZfZBHDSnB8WIMwYb
26NpUbZMGd+ahzjV+MVm/CtaHBd6mTi2txxKk+nUFejAaexYAy9NfC3U8yjHc3Aj
omVyf2kYBvLXoLVcOLvrtGQKCpMC9GYyDnNpsPbb36t4RZbGnOfUrxQfZb1sEUXV
X5PkN4ZHWnug67vHIH1S3gHnvNhDcZjmxeyivfjxm4lA76w6DcmWjI9tCCH7/aWs
46EQGp+qHcyvH4+PCSuK0GkFpkm3GuHyXlFsSTPIzFp984B8Wy/90/3Xx+w31371
W75ghDB/8UPMA1tJnnXFVcbZzbw8hd3RTgRYlgipLCSj5QgVnwBs9KQSVF/t102M
GjJBKZWsDP/upKZW6AmFjRyfS0w64kSR02oTxB/JlRisjUBuuTZ61B6UJXrIaqVo
vfC+Yqft8oOzD5AfclaAWY6a38CD6/CVcQ6PvNK/nfCvCyraMqen1L62oa3Wb3Ou
IQhISu71Z/P+5zQYSF10D99a9abYpjBw63uuNvNFK1qmQxQgIYyR/9uT4LbHtK96
d0Ycqlr32j3iBGBou2kji/RIVzsKgg0qg9dngqaJ+Ho9QB8aHjUez6dy4ebUC6ql
DyjJIzCd5GEDEu2i6/2QawHOVVZl21lU8YCs4tFcAwuKL/6ABwC2lTYqFFfHnfZI
R3Mzkfyl6bQFeJxNwHXXsyQffY25O/Wfn+Y5Cov5xavT5yBfoFx9nd4+ugf69ftf
iScin27jnhNk9jok/XjnsqZCk1/TpO3xbqaP0Ft/220QCVBt4uqSesbpC1Hslt6W
VKVO9kcQ5wiRFgdsoCjF54GMNw2v2n5t8BuCsg8Vs2mX7DzwfOFEzOmyBl/KIDg0
soxyiyVu48p1gUqSgXUbo1qZMcb/yztjeYvJmiXA11q1OzW8L32zcjwsQxZ4tFkp
jlF5edwlrSC5ddy6PdfJ8cUcu3YGCI2kwE/7KryMYQocz8It0USqQNRv/eHm1GQ+
XrifemDxujIn1D/ytN28kIVHdbGoAmTc6FjQOKv8n4ahWvGugKCgvHFPj/H3a+Bm
iYvf3IhT9+cO0uy2GLG/8ZfaCgf773tJlEsruZvhYZwbC8DLnQXjVAvMKUYwUIbg
c5RhQLUCcXc6y7IcV0yqCxrbLh5sbsY9MgaaBooCbf5s/jarnAMQy7GTRIdkd9fu
fBvNVqkQj9EY81Azsm72O7HS2S5PItqyFBae5PmvFgg2yftxu9OaXZTKNeHl4G71
LFMelPe+U5WAFP3IWk+kIJ78g/B6G3z9OetN2TzWR3TtrhjZHPi4FHFWNWx0qKAz
tb3KkYCLhHmJ9sxrdi24n2TN+47uEYqhTfETSJlXWqer83HKBnLmzDGUHG2vcn47
65A34JioGNvZgOUJAmPo4sBksgb33KJyJ/kg7dy2m4sNQIBkVyfkTqN3MoJW7lY1
Mz86sypCOWKK7vmkHdTB0dbsb/2KEM8dEg/oAZuAIF3AjKLLYJ9Apn6SMJV7fHR5
eymHf/l7BdlRFCPlfsFXgm0N10FSInx5e2uU7MqhtM3rkC3ytSoNQghcncmCgoT6
ADUKZFi06iiLbe1AX4baEoY2dlXHelDLIc2qx3KPKpRSEQR/unpmdLpSW4IRIiF+
d1ZpfMxGkZNtXObklzismnogXVmutZ9nS/PPgEa6bMbuPuDjM2zBteZy/zfzXja5
LCMTbtcHGgVo7BRQRZMwovZdVYRxJPDjCV6YkHGTpGils1mZu7fee886u/u3w5pu
pyOVAgFJGQU4pjJ+CEff7HaxFfjwNU/ZZNGM2/VsXg1V7lQuGPSln1DnLcaSbs6L
loM3QW15QrUx6lDdeUTlZQefOBwLqEI1EMTd15LDMcdMI5sR434duW1dX7QgEe4y
6LG3CDDstWM+Wf2L+3QfwYFu8zQfyAQLKiR7iBOG0eVPf/hOCEMadtEMKYb8qU5E
U5qDh7nNJK5IuwLG/E7NyW9J26GMARKVMt7j323YQ+vxfrMp4x/8QoBqYHf6ELtD
Hounn4oVBVwsMRrHXd+kNxUmpM2nVuL88PmYHaUndOhIfCcGYrVyaXV9v7xI+L3C
ib1l56Yjq8hUY1NfR9sIizQxwY/6pbz1gTV7CLkRwIhHjxKD+yEhvEj2RjimpjW2
lopIwKhILELJduM8MXDoam6g1k97XlPTEr+wfxtzDcYdl1afMaDgo2isAwlEYidc
VHGyfrdxmz8jFwM7ekDsN25Tnnu6+8uzgSWrumf0UE+m8vOVtzGdde7/NFIpD0L/
YUKnd7G+c/V0omRZIO05QjwVrky1dmcd1IS8violyfFEkFcc1MFKKiayoCveCm5I
SWiDIfQjrl9iv64uvZpa8As5GlAaDSEd+TE+UsiXJ+s8MrBkfqq5QrwkIytjtIEJ
tWl0uM9cw6GRvLqulx93dKTywmHbhP/FmK9wS6ilJXAWCD0TK7hP1jnRxtWcH2tO
vTkXOkCFYoEqEQXQIQ6kNWMI/SN5b6knDvRWOl/TkKXY60eSogCTpa4jR8au58tZ
MnYD7NuYUqTRsHaiLzWFJXsHBawP63+gk5lsvXxm/hXJfm67EXxn3MbL/FeWZa6M
hlnOWHQi0Mng24NSp16rswds5lw8RkTo+mafpe6Omaz86trcZQR9DveRAytQTq00
0ZnrV4sl5zIgisDZyD2W/1WVtvxmAfWHQxbkXFlcCwdsiwVr+STZon/hN3ctjofA
/HWRxl9T7bnUpieFQhQ4IuljDZTqUoLUnmntCUWksPlvgEy2ej5ggRqktKF8Ro+p
u2nZTQjxPRmj/do3VTG5RLhXefHPTKumX3cRi0RuYlk2cpuBLGeLHP1pbWHjb3PY
FMPYfRVpeSgDXk/k6Mu2d3Wo1itP8o4EWaquZQoOBgbEewz3Yun038kK3q1AeWWX
wDutrSqOw7qGS+fthYSHYJSEsnE+8Uy8oajCfZXHNSnUNTkF+RASFMxoIkZAHdi6
rhzE18wNwN/831cs7kjAu0bl1s1uROYE/mSVB4+dgJZogIInncmTb3AZo8gaS9gZ
b0tUEvU2BtRy9dU1cY1xgUM9NN+XZknQBYKItRHXWasbs/yROIebEjUpiNVWmAjO
1Jn8v9hK/0/DbB5A5S0Ls+0iZa3SPSkUBXojYJ0ZHThLpVnyCjI4dPc/uOQJR2f+
xl/OIwNeEI8wC+3hYdEL+5w1OOWn9uSSqHqyhNgEU2zs4NudC3AXtC8lNpiA3mca
p1BMWi4uvwVejfmgeXWvCDNqFWa2DMdER+v6hQSKuIIjE66D2vplVcoHH1vfhAmW
tT/3hcdQnAGMnH9EXxlUllLvuLgeszai9r6XB5ka2/aVS7dPiGC+QGdvUOaSSN+8
exNCImMTHDrrgwnAvf2/FNbQESMfz+/7EP9qxDuNaNMYHp+EJ+d3n8JSJBOGpDsM
hf6O5H0IPm5Z2IVMn+C4a9662llxptQZ3/rJ/RjFGnxccNyj1ToejgPQiuQTr2nd
WnbVj7FbzofTmagGxjgQcuyL6jwH5S66fS8gpGAXwFqx7DU2+BMXk0d9G7KTZgFb
Ubhz7rAD7fDMEm5dsr8PzEkHjracMdOEv8CII7MRSDloTSKkGuo0hH3fna93gpi0
SDZqrcJ5fyh/3mfJ7dGQaXy5dnij5soszdXkC1el31IdZmuH72t3pljBMO55JTqE
HGJCdXE4RzgRkpByyZ4fh29JQK+KFghjYhIFdGzDW/bH7UWGPWBiXUBSKBBzNpKv
Na4RKPBBbKnR7rfKAJLDQkhJSiNzQZbGhpiKKDeXdd97cN2/CiSpn88HlMhqSjmb
XlQFgxqhPlvq/ModUDzNChTB4UNnYjNauwmsP6qRx06DBSsjwVrNrqRaATdiQw4m
fl5GefW6/I9PXMRRvXejWDheTUXcqofLGNntu25hOM7JoFd7ARtKHWd/vOF9c+1b
0esHVosCfC1YPmW4Z6Anqag9hPkWgh8i8LhWqhJ4cbEun5y88H7U/zTLpCC7ryVM
ItzoQTqw41BgsfzcAA+ITbzkKmjvat+a67/Ep19a8l9625/vx0ncKzvDey8ZXuow
pGmfOdhLugZ+WMYCzvZQSbJmUKcAvqewZHZjFQNF0eQPYBSG3yG8G0d0RfpNzE0H
NkqCFTWgFCikLHhajraBOJBOHcoma7SuA3lKIjZH4Y8Ae3MR48Vn4tpnTahcjgqT
+IDLRITfvj24Z4DMQx5/apb3JBg9OB1GCEQEi+S++zcqUoxC2ruoCtjneR+ng2LV
tKu4r+dqv/CHLg5idYxESSaY0Skl9qXTXCSQQt2iPSWA/Mfs1gdaW40OFLJapCAl
t+1GgXkV8+P/DVq+EDW/LVurcb1wxrOb8bwxDenZTLMA+CPIglfHIfuEngdS3J2/
40YQ6EQxxY+mnsbuA2vPZjIFtQCHTxQrxPV8wtOdjWRWinNv+wQjRQcGI1m88Igo
1XMg45VpoAsUftmJuNcRr7dy2UfCcZaGCeRH2t7VOHMtYjvPLPLcRSWRuewCS8m3
vJdcCX0n+NQNSNff3anZD2MWQmdh2RlzeaUcWK+u/VYD+OQJav+khgvAj9e67GTW
squbnbxkQSogtH9FB3KudDvcFDYpxO9MwLRUZr21KTXoghApvLoOakjUyFbtewol
x/UuuuDOxQu6ZTtruPvgA0r0T3FBOYV+2f1xdYqeHUxAYL5n0NMPyUKGZjc8hzSA
T1ln+5pjXQBGTfnbeoCFu/XtEuLzBznUER8NcijwXYKNZGl783/zoOVsMHRqGRnl
8pqfDl/KDBIFjQSYBYn/eEL87sn4edPsmdZUMuQJDRaCHNmycVAyEh2yJOhQYm7I
uj+vMeqveVHNBDYYXi8Li/6LeSIbS0OT7EgzLnO9FiX6ru+PV8oLNYwMPLbQCcVN
agzLvGXxNu22EykuFKbetID47OnYF3k8/i9JWIG0CR+SASExgXbhppdetXrErnCC
bjcNvwthmhflFCcWqNmc1pv3SQBkO/gK90P5GUrHNKEYVGW+GUzl8qG9Ai9aroz8
hgodIQoJjrhiw/0fDy2GorqNZHCB272yOE80nj0kiFr0JjYTgAGei+W1tIM1q1ld
hFg571S04aw9W0o07JQ6AyVpg2+rH6S9pnm9RbaOXY0DRq2v+hipLXTDNdB2FnTn
Sh5lOx8pIMrFLzcqmkfqzyvvQnWtse9rP4GKuGaDVQKm2UM1q9Mhud8OKfBcMFtM
ph+bpA/x0gch0lhKN8b/aKWtL8a6DwfO65NmTmT5R1FOcqlwmFOY9Zibg323axXc
y7wEXQzYfbOXgKOz81Dw16siP7FY62eVJXgqXcrFnqR6yafZRTUD2z5eyGvLxXlt
iTyf4Siw2MnYQyVj05rOU4FnPw9Vc2vm4XbcYl9QXvPYs7VBIBM6GaJzvychjjgz
TrtKmNnKYQoyZExyfo+2kuwh5/D4uVAbf5MX9K1uO5Oz4Y6YVzwffsQxRUJcMEkR
DgPiRxijgGOY7gDY/nTbXIta8tF/gLSJgIuZ1rmlJxzXItB2whOH3wLYyXz5Fd7X
VEFmWbS5FWuq8XMgDXdK3UcE6KMgoiJTtY7VyAqxcinCCfHIn2hw6peTCmfnJnQD
PN7rRH8/0I5Z4jDkmomyZl5QO0+iTovLDQ7GV4WRP1DT3YOqNP6JRISZRQjrORBD
sMFpml7do9Gz7EZ9uiNObZeaZ4neSgLh8z6LLI/MzJ6frkGwVt5Rs/3RvuJ+ypv1
hezFaMdyaydjQPj+45YIsTxV2AHzRK+L6T2S0SW9idAtSSvNy0F//Oz8f5a60+6e
+Q8gOCc2sK9OUH5+Yx3AKawlwslT3okuo6MNtEN56ajyQ42wQrVexgNk1Vo1cLUn
A3lkmSX+HpI80pkoxPIW/hM5jrb3W6uKw1Sb60eSct3m4q1Zqxl9EAQeF+D/QVCG
BNbWixpn5bOwil1HTeNq7PU80MkOGTx8zrzemzmdQ5krZHh5J67fzUcJsLAfCT71
HoHTC8z1LUwb3FLZfGhj2ISaOAYztnG9PgzRgQJy27Mq4ig7oHbNKaZIhNkd9DD9
6oowuAFftNf/tD07hlGY5DDll0IEbF5sxCBaVMUalZeVzKrl0iUSdA8kCvObuMxJ
3d98LEKExedUyxXSRAZK0uEhVyQLIqs75kDXq0/gPC2S8NH/NXgTRvrOwBOirlLN
CdWfyAOzWaXBGGnNe7z6Rv2qvFSe/uLcMruJN/aj1trd2Aozg684yU9JsfqjPnR7
gW+tB0SS/AndlreSNtlxVuKJHzR+LjvI4d9yq35VkgeWSDd9awmL38CiYd+n11F9
aFJ4NKa2Cen8GqgtlBc1aO/NhVAW8co7rNKWmnojxpU8a43iRxsv69DTOcCwS8jb
U94F2sGHu83bcdzFlGND1yBACQsaLufqFfmI9ZQkOqSR9LdAE2/sqvxsIsxcw2f8
T+r31JekJ+EcmOPOHhebT5XZUi7ymAlS6pm3EOHisEf22jTOKVks02x5fcT3ZSZg
Tb829p9hoXPm6Nzm+p7kG05y4VjT0rcj1JiwskPZpZn7mTN34LXTZnP2uCGtOyyK
N54JzcUY2YMnYlgobj++6zIwG7THW6LrmK/UXY0sjQ3XHVAOwc07kPHuEdgyRBzN
4WuBVpbfJckh38oxCQlp3kbjs+O2f0J7QTKyyavTS8SH1Ny5m1pUBepKxGidG9Hu
hmWt6QrVveRj8Cf4uXTUujdDLW1kWmrvyd92oeGc92UZM2gwbRg8AnisSdnXmhqt
4TVN/KVGWirxKhVKfDMvEIlhlQ+7QZB/AkW02LLE7GlSSOZ57oChRh2LRwwAYcNQ
HOKO+dJEw+3UPJmlk23hzAN3KNJUQwDSuMT2GbfqqBmxZA46kZiKEgtWVWIrcagj
5EBzo/oOL+HQLZbQXKDg634XbFT6B5HnVIXLjZHdvFYLYh2JM3P6duBmxsi/V+I1
BRPnYDrZ3+F6p+znTJ5dZP1VLBE1nBr9ZjqKxv/SCxfPywqaGvpJ7UPAtBwTC1Op
ba50+LQWEQHgI1e6pop+BfUhYSsEcXiQMMsWCUVCjx108cJXMfj/fcaHO347R30I
lddGk6wbjVASMcvs5Jw/LY0ygvuYnO5rEwzcHTqrfPIY8CR35q0fkrb7cT+8YnIH
W5m2UFl+TVAczGUOEthS6UodZXnS6a7Pcw5ivrTfdzU4zdctUzucrsak4tjmmk/4
UliGtQrgAeB4ySeR42uK1B+xmAc8csNfd/lQ+vsy1oi2L6IOuauk2UFXTd0+wZ0Q
MM2aR1ztEY7ZaepHdeDvPU8uiHWlrCM4gJGHK8HF373mm+7AaHm5ZCH3+q4PGOCw
evT9201KaMkta01pI0zID30wBmlTw6nacxZ5Oee6wvq/lt8d2VCwLyk7Shxyes6e
cJJZgcWrkze+WKgp5wjwFPrQsD+lPVQrnR8xbFbl74I4SEaSdV795Wqg9jm/efO/
XTDjntCN29prfqnte+wizP8BZrUFmU+LQQZ/tM06GM1IBRfQCGlj1DT7w5G0BW33
hynNVVJHIQ9r9RtK9wOn50cRRNXBwyEHQm6r15GfLeo49pno6dBD6Vu8YXBPjRov
5D1lK7OblzrJudwXzruWvkIBOzpNuQD1gEbUd6zdnuJeCJcHacZxZVqxoiu/8DeR
zSmGsDRti5jCJaUqzNmVUApfQgelE6neMwOyoDxtvnDzA8sa68HO7ef0oXB3r/y5
HN67/i5Jc5vu0Ws3NE9bM3mnuCezSIj3WlvWOMOHzIBJgnBiMvhFknGSc+A4aMZ7
PXODO8gv0WxKf0VTPSWolwjHfGVXPL9v1dJ4+u2YTISwtJI8twI46s1IqkDa60pJ
jCD9FhopibsfLpzWCLRJIANtClk19/h9cSfmFuQHO+Uoq7ee6D3z0HKazc7AKTUc
j9rYxQx6uD/2sDaDxwz5yX+Mxlubrjpes69nDAO9M7OwCalQhD+Bk8LvzIg3gtsL
JeZVVz1gjvQSWd3nulKh3ub9xyzre9sC/HJWw8cIaHRl8DhFLqycFPBvLFbjY3nl
BeLYRJ5Yyl6aNhWHxmi5L6pyHKR76FaH0ezzFHgU2YfIBlCbcBF85Fk8GJeTGwa5
ymxNacTIyP8xhDNwG4qO33kNoZLB7VPqeBfqxEJiLov3UDIRfnwp0CqJFQeVdgxh
cYV/wYWSIbuP6SgPTlDQPauJPRvIh3KtTEkVZQdjtWZJekJIMKhOydVnpDoK2Cll
16NaZfzBu4Xbe0YC8A7ovYLzI8iB0Nq5G9J4VR5mWtFezGJa77ngdDZ4ZjDFOWaF
1tELruoK/PNIBwYkzISe6Or8/9+oRShCTE+oheVky8a/GJWoOCLzpIpk1YrKA7MK
zX6/5qnYsKM0/Ftf+K7pbFgsnxJHeI1Ydt/n3FkIshS6S3PpBHUQeIfTdHzh6M02
1drnE+6qGffE4HUzW6OrVUyI7FQP1KOTxhPt1m3SVKc+xfeJ45VdRs2bfjD0Q7SR
zfbH3I70dxDJivf1txhxaxa3NwRljiSyvxTu3sd4MWsskv+/wJ1zrcveGth/j419
NZ4i7B0oG2huJ47RWhq/6YNgrdIBvbhh8kgwlxs+f6KK/fK9sNX+w+LvRZc42Qih
TadVpdsuDvlVJPOoBYNk6SgSvp3tbSmAFgj+iUtGsD4YBhA1BhzYV1qjnqWsstSc
0wIq7hzdn9hnwXkrviU5ZHnS/V8mJNOwtLV1DhhDeNNye6kbQT9geTHq3QwMma0x
VpK1uLus6eNEXPwCLvVHodyTvhrMNl3jbJ2HppeUErXcwisfpSOe5fVMr6Kp2Zi+
bHYA6BUSRm9YO9TTcIDqiq9/7g3QLHiZTpfIm03qAL7b/cMopjQwtYFZy1JJ9mXG
9xqoHkSsAnsa23BiOW/tPbcZTJYXP3KFMUJvbgq4R5gk2VkEKi7AiiuE/fBfhT6E
BwzA6XTkQDZXdGhvq2dDI46L0Go4DJCCnRHHs5Xi5WzVF5oN2ptuqU1YOap9fmi5
UnZZ+CM3wv/ua1O/2fA2xMN6EQyWeYvKGCD1yCdWK1DjOA0N8pnHWWOcjrsEJwwl
9RYKeCr+nZAu+WvEx/A+3skhg9Qzz12o2TgZwvrAIxiDGa8/zW5OhklMQH9LuD9O
SVXrzeIYkXt3NwuCuskcuatcm+STLkpQhY7TnKxezrVxEmseD5vudAg/XsmFwLBf
kUhhIglTXvhAto7aamY5ITyY0EgueI2cC2traaWqw4QoU7Y09hdn9VI+PqLBYpdy
k5czAH6MiFWXMh7RtUjzDDR8ubfkeoAxulOD6vpBjePyMVg84lxmGEnTHRE2TSAN
+zvgEC07JAYseca5XIF8wBMZbz+octSDltST0XiiZ9P/FKSrYTp4AS/mZNtrzURU
r6eiI+tQr/HWHuOzc3JITmG/DAHyAD4IjpnwaoSyEVQoJDRBEAIMa/BxlGbq8Ll2
obgnrPJGf1fJuhc8MvYRFNumQmPnoaSrcWJnw9fBglsYLUSzxrZrcTKhoSLDffHc
bXGUiTCOP8/nFQ7OTbQ/Btj4dgF4rZFXU/JZAsrie3unwFWpGv6H+huQSgbRGRuT
1SXQudQGCQKLiDkerG7XIRQ6G5C2z7IJh7GXEsgHYQ8iQFN0sujVHIrzWqzljd4m
S8tpcsOPO77pl4gRA+td4wKhxgSkN9MYqH00LC5XB1LngvkzHMjrsMNl138oxn6a
O2NAWSZcPhHoCOTlsQTEJ28bUHBJCS8TYyqPwA5cTZcI6Kt41c0IH54d3lRj1xGt
rwVdgEyha++G080+HBhZTY4V0B0GWZ4Vjk6Gkkck2MCAfRaRgBe6f2SS01oYZ6wY
1OeCr3qTmucWMBtfXBRGbxtQXNzdxUa9jidKK+3g0dROJtcHjSSaAnVhdWGGewDs
mV6pKUohJujsFSTpjVgK/rkP0SPYmizzjRoYC7JwyzYVgS9EdMyBNSK8vPQIuBCb
I4GYQrRVhH87/ThEEGzWsYooxJCB7ay0n77msqMzHV+AuXpK2SOvASowZRq8cTHM
zRhGQaaIgZE5T4wmvijKP2tbQ1mnC2QKaznKXQB0HMWuzQ69flE5wXOHNjCSu/7n
6qUqGDNrAciwtU9c8INFV/njrfmuKg1Dr0Sm58IW4ZybJ3OK7XLnH/5+stLjiS+7
rRj6dU29zVe0z7CppyX0lINVb3RICP3+yfbS8vDAayttehfoQwyH346/c0NIHGWp
j+SpoWQWOvX2HZ9BfFGynDVPd79XmzlZv7luUdKkbKJ9dZn4Pp0BLYARBIGgVbjY
NxWhUj5kCplQoNsjAzrxmA+sJGPJKS4A9n/9m8vOmcyveYXjyq5CD0xi4x9d015H
tI6rPlQ+A9Y1369z4mWvYUI31DDmnhUgAqGZLLoz4u/tNVWZJ1EwNfZDin+GxM5s
v9WCdv3aOZdnuid3ARU3UgcY2HakYeIoxmCWlvo7eo/jYQhlF3ZbVZmpwwWa9Uwy
xViQL8rF2A2PWaymEp9+vUZM/sX8ytubc/2t+Tv9oYS6g3sGY/w6vcYj8HQpoNeN
tRSG3hyndZcalz+c+Nb0/VJJWFCJbn8L8XeVufiQyg03eFimBDQ6RDtwfq1oDKoi
EaBUXMRG4kLFrADxfvso8NDELy7iuAhQbxXxRjRwAQ6WevDbYkkBw4VC/alwn5Wp
gC0pNX40KrZc/VcccIEBKNJBef909/x/CCqWyT/YwH3fHeSTyPZKIITnsa6ZkFyP
feEJuEsBN2ZiwWPgsJqWxG+5IhZ2qQv6Pt18i6+LoRzsqiy3wO4HfX187+F435NS
FiRr6harhdtfuJGMoY0CATPkEY/s0YWEYWVJ0HoRv7WhpnH4OxjAv4ybgy28KyBu
uaB3uOVQy+mFdrhb5CLv0pGKC1Rc0rCzAiUrUOh+NuTTQl9tbsz629FIckglRQVW
e1N2jNzUOw2tG38yeDXX4FM948yabx6I6tH3yzXgdyjEcmOvsxAx3l1JtDOZSkgZ
Y59MvCbR6aXLVTAaunVqnrNi87eyjmA7OIzDBtRtQbLCEuJNa26ad55+ijSLlH5K
p0I4f/A20iDpjkonbEQu2WJJ3g5lHZSeViWnpjlKLqbCh8yI8E+uun6JK8O/PWMa
8EATQtxuh84PACSKqYyDPN9V029KAEitm6TqlrrvZZ3t64V0/qZDu2KDeUxnoyf2
5EE06nJDvDig0iNu3jcorvPmmUH5vCvTatpCxSwvlLPkwHVCgs8SYlVoVtbbwHxu
eglG79mTelUZ2mCvyv6YGXzi/JaFwAsxpQ0VzuvdpfIqCDtDkq+/7dxkBxMvXjmY
X3vGwEd2AA1xSjf3fCYYklBN1raomEdiZxolIhhuZjH2EiVlmdNijNwpRlYpd/Ag
8FZESaMirXnErtHR3ZCq5G6E0xfDq8C+pR8TU1IIWygBZ0uFam2yg3GNQIHZcDz+
KWgv6aCvY+qDZ+FPQTiassneUDXx/t/21VdHDeezC9q7EOBvRHcQ0nNqGNd7Cwps
EYi23SNQAihe24raWCDlRM6IaaAAgJoB1pxaq678islXK7lxH6CXmWoEf0GDaLVl
NVwJcdI9TAhhiB8qvYfDL9TF4Yo1eJ3hBTH6I/6g9BQlqzi48+L6JRHr3mGJkyQ4
SnFmcB/jkM7IJ962/hBITHSaSARZpY4sQFzK6howxfd9RGSdsX75oJ5LZCY2d7U1
IVCF3qjX5BVxf17o1amLv2SNE7Ya4yiuEl7aL5KU1PkwFdzoIJFMHdVHEzaBAeZu
UPM93jxmUIfW2UHYKROusc5Zf7KPUlnFc55N1YqcLqMfVBSe8b475ZCzqcS4q4Bq
5AqkIWqr28IJX4N8REw3k3C3f1Jm9mO04ZoBSI34uBrLqZfI/iC2qr1hYFcy7eze
NK+ef+7Tp6Hu20Ig3eG8nhTkJ2439XqJfiPKaWdVxo4UHJ7BvLQHo5N7P9Lt1SvO
F4KTtZ+ny2FiEddMf7fdlTUVsrwlZJaGYBWU5/0EibEom05XU6P4LHR0OeoAO2FW
kKb8P3VKjSHm6mQtGQOvcEKEVavKab604tEqb2Y4MuV6YDR8voDiUkXMOmo0Mab9
H9AsYlLzS7urZN5STreUUxHCVYPE+VCmHHZZ8Y27rgXCtzgIIFIY/mTicdpBLoLe
HEkb5bgOb15ZbMAzTnzOd5zFMJGSy8hBlRxTECaHn7x/0hCnluImL5zJfMj4TIfr
RxzP611UOpMuf0WG8JgIj0sv9FRgX6x0KwCKnQ805/vozTC6D9Ewr2XNlrRJKVII
vqKETw5uUblwR1xG9mwJpwjuUPyoIASh4yjle+Z81SOZ/J9brmMNyU/CmzC70v05
tJq2SE76/A3ROtgGsUfWtwP9iKc+AtT9xsU2AmzfjrZdNCBGDWQd+Br+7HV3SnEB
Cu3poqFo/VD4kUERx9MZzmY7vJ3op30RvfRzUHeuF0lrnBffEcaVXvdicnVYMTIh
zbsHHcLApowECNYNbwdNTqfF0r4a6IRB2TGBeYdQjwCHJiwTRkBfZuWTfGL9worb
iesKfWVpMA1Q2YGB7v1vUd4phJyGfPy7lU0Tx5cwX2sHXNpF4MYcaAYlUBQeekPr
jEQ4abxHLzfP2KXEu74DBO9y3jCn19bw5JFPcKwagkMpDQtVD81TukJE+zlP4tJC
oVQeukBrtuChV/bna8+vz/ijUCzxsdRi4jTAhJRFXjNjeZC97bMVFxDuDNLDNbzF
kCrt46x9eSAFps6oy0ldwx4ja1M1hgAgUPuJKZqetHbTWez5jtDrHrmFHAZ8TQiS
47nFRGCDlhi0ZfudJhxH69Lx9SSqIUXz6g+o4PtQeUe5ediHxKIAwF/qevHeUyiz
FlDy8gebwHXXwWVukCPhUsMrFZir3DsqmkvjQEYWE8/JMBghwAfLwXGMWfgC2++4
3eJx1X7YGtwC3AuYRzMMFkAuBV+oXM4eKD5PnKZagVW5nR7CkTybIDT0Ahy1Wr93
Rn/tEwiRpc6XNiNQsGhB+tCHtlOBpxvYcDWkqiMKugk9NTic2iyrwrP+lfgLZ82C
pEwfbmag5RXi7lS7FEQ5dzO5GJdpjcTf0IUD1YtlFpkAajYpPWTwXT77basWEHNr
jmObGf1HHf/4FlyczOm9YJ4pFbXHaeODjKh4PgQxMDWOdi7U5qLrMY/8qYDsptg0
RPnGqLxdwqqbWOEGGFDzW2pC05TuIXQgFKOQ6Wo//I3vDp+TIeVs4PUTz4Ut8mct
1m8T8Kijgs1aBe60/iynAah16v1pNdxg0l038MycEZ4h+qwR8RQxYfxfeAV5GNnN
fUeZ4BdhdJaUBpF3jdapikI6Zc6I2gGnAhcNRncCsPKxlr30EeU+it4LP1oMdin1
zChwfjh6/bbl1FXDa0Bt39U/TJE6IYoyN24iXsGUwOVJcxi1N2nNUg4vYqPzmFOy
P/Sx7dXLkTnHY353Sxw7QBVmk0thyswpG8p94dWmbcGcGhIKKgPrw6GunO8HmN8F
YbrHpPYGO/rafjytT+oQFJZK+GS83nO4kg3cx3hc/hMMdtO6wIqQAYLEbkLrqkcC
Flmna2mE+LyvWgpmQ+Qbpvw2Y0EeAVcjW+K1y/Evu5a2QS73GDvuiRX28FbCivPD
snyKxikERu/ogkXZe6QjGcd0AeRR9KeVVR8kudqEr4M/87yfMgVE8K1ByfcY9+C/
s8ImdikxTZVDMWhze4b/FFhUg3aKPU8l34xxeUHPUrOUscEu5Z83T0asjjqQ5pO0
AczqXBRQEAfceWiDBQc/r9HxmZyKU+jZJmm6YXtJ5LglOsx6CYhKxMKtnr89ra+S
LJM4w6qjwm4uc0RRUXOwZaGy8AVuXB3w9JY+6gBdErt7jlxxJ82XkI5P2Oq8qmpM
ZBnna974jdnoRIQ5qcb4KgHjq+vfRNvGs9y/olHJz8Y0eYIe+OqxYDXGuy8u5C8M
LIRTz8fzqfe7g5+cnjmDfaU5zA+5eGsGjqXp5+lj4dJFK0JgY3BFjF8oUZi1LY96
3F5c9ll3qCM3VhzMOzxYu9m73nsZswSnayllQoXNot4tjEXD34PY1GHZbPKpnri9
ES1Tia62MZReZM5ZuE8uszeUOlJxl+y9eqTOpo3z3DdT8tqjVHUXXwXcgoJaqPZD
QEO9JBYpt9bybVHbi82VTCkyIcv7PRUFaTM/hZIarzGY3Hn74J5LjN4WayNRa9XS
v8rbIlFTZi4thMnFt+NaXX+EyAK934Y/zB5b+AVjrdc1HjX6HeDKKOkV4xEJ4+qU
wVypsG9rBEQRH2iItbinNtz4wmHZ/sYrH4xPyQCZczi32OdHmdR1Ka0cWNBCNQT3
pwGXmXYdPRQxxy/xZoGn2GViEoKeQ8LE+l76+OcHyly+MA3MZTfhbPTtrYMgDIx9
IRXrcXy3Nh4hdB1/htd/cSkDbL0iBWHgU6EkYn2OEwmccDBmP/qXNv2SytjjcZ4T
yc/PSuXGetbRUA9pVJcOU1Tw2ijwdjUtpIljg0MJ+bfg3DMwMDvL8T1LlOieDeLm
LSvcZijNV/arZQSw0Se8W/2Gq10pHuck17KjOifFbn64OJgi2GNQL5iNzvebaqPt
QVePpjKlS1Fm7c9P55fhHSJmpBGJ5fKtVVJZCz7I13C4MYN0Z87LCtlRwFHhCrX6
CZzrjN3auolSJoYYzT7eaudU9OTf4dMIhFmMtzoGt3dralOZp7aGGTjv7CeE77iC
+NJ5vMTftvTYHMzfoYrCfcnpDM5tH23FJBVvdxTD3OXJCIVFfUB5h7T31hJg3zdV
6tKfGvDtRhLS/ngmCrqoOLV8HIRmQ2ZJ45FtX5QVm34pacAE6vSfMmwYAmE5b3fv
jxp13v9RD/x0C71Qqz+dhTbAG+3ujkCtb8KdoKhAb7PJc5yBFoP4jp/YjmtBW9k3
pRDoYOIWzHDsA8AykQuKe4GhCfB1dGi59G4d+uYNbp+5UCYM4o9ndvBM4QDU7bpm
JmCFuyPLW+mDISTakB5fWjj2RdoUEJ0uxBlDlITQFTgfyjy3b/yoz3a9QFEQUmA0
bPLDqIi2hYIPoO+ebUnUKeJKFWluvIapJSO7/GoJD57QYZDAtFhlbotmEWEYPwK+
cfuINmpu9e0612KHF6vyBGuiIPm4MGck1x/IEmvE5ih0q+WmZlRLLzMoUvuFSXqN
T78FP+/s9WU7FtjGuX4iX3f3Pu9HFmo5M1z5nu8PsOHoo41WGNO4AxLHT/w18bJk
xJBVOEh/djs0fcmBK7Ad7+4dmCryU/VW4Wlj6FHKHrMCLULxlEF82O0rnZcotD/K
41xyXiDOiqj0yeRj+KdjeTEzEdDrb1uhUStSZSREx63CM+9tr/o9DNBzT+aR8ngS
sg+3iUvOz8QZtYdQBP8KbK+zqJXvhze84d8Jn2jfM+YHv9gWrWDVrOQLCKHtNlJA
V5zezZgrPOAui54aus2yvzQIBTqGI/dXqHf4FaOCp6yg1dk2ZMWYM+7s4s5hlPME
HzTIIxXTMeo9ibDwDxC4T2t+hiHSrahp926rlGuOXfcq57q/oFWjnc1b+Vu1/b5c
qWbnrCmkxjX2wBL6pq3hsWfFY15qq57GOm6DtsSez0VYRA9mU27S2KrLj6c5JfA2
55ZzME1bx6ivVFbVdVWE96hjbMSEp0P3QjLzVIFNBSfEwtL9oZiFU2Qjue98pnE+
DnsTiBNajkKb+DKLWNrwj+cHjnSrvdgSiu9NPMrxaetvqZaqgz4mAKGfGevSSkcf
9rkdqSkoWONGtlZOlGAyuhpDkHakV1IteuDVTd1oABoLYtQwLo9i+uFzvmi3rGX5
2KpHR8CHfzxFpvGnoUJDzlY6aIYRVOduBY/Ruso9Nu/sD25KerniERAlLIlmOS/U
ff4f4g+fwmIizIdNdzpeYOPguZUEf5hGCxxL/xiaW9qwutKnNhMJTtZ5s3ovCvGS
IyfWcLErD+dfTT8sVmrxbo9zLqTm+ZmTNeDU4Ms0exyOLySa1cVtAwI3UNTzbDY+
i+cWwYHegZMMrNIVkrs1+sYZ9KrIbY1/GOmHNOfumLHpERpZSTSrP/rjD5RWzClD
50x8t1IhxQomhuDTbSBKdRnBIXnnSwGeNVTH9hWhGjFtKC+mqaM5JRBkM+4TVowZ
yGCuQOc1IYHVVRGdNJcmwyQosYBLj4s9NqKX74UUiLfDfQkXFKUhol9Jv7rxypVF
n1Zl1+/atHKAhyihd5yLcqAZPefrhYTsAP5kLBHlZf8VwEno10AdFMNvXnPgjxQp
DGWkJOdTinZ3dLe9s0CKxwftt+RW4qS+xrE7sQT4d4+lE9B6zkyOlerDj21cWeB0
2rJV/afvq2XMLg07OeklFqJpwixU1vRevCj/5uoIURjNbxRVrIc8HDVbjqroW4eL
Qa9sveqvAbG826Eji20qCwkAsGIh5l9yZAl2eFYtdp9o2wxibY6YyTfsDpsm6xeF
FUE5n9FHzJwNYoevrlxH1ZiI9TtOw1a4/xVoKIhMKAghzk6zIRM25zXdKUoAKiBq
LRugibuIZf7V2NyPvyA7CcfEjCohTy2gySsDWL56OZwoPnddBRcmiCw5q49ZSAa3
HOpO1YATxj4tTzwbv6lDbRqELU4n63k3DFl6+w8EJH448vrgJnCUxtF61tAjPkEI
N/f+ba4MHVlPtCn8E3O9mcJ0GEkkw6S2ZUKU9rKHH+ri0OblhkQMm3U+3NE4u0ZM
U338G8lUUY8/S1GcS+XLM1I8U0j1GeIDmC0/v2jRGVEDlvhutweQhskHhnY9n9sl
QEi8VUP93N6+J9xNnYUBTqJ9dC/QKwDESlZqbu0VwCwd1zeySxtMv8/34nSVa6Ic
T2B5RCMMrQh0/y64J4EK3QL4Id5nbe7fAGfnyZKTPxg1fDCODWyRTTov5t9JBIJp
7t5vjpQ8iDTNP7FRJux69vte9kcs5m6rpD3VCxsoCIyetRZ/0cnhesdc6dz8SBWy
S5nGdx2i2jMggxB88D2Rwg3BB4xoXwqmTctSPnCQ7m/vzVEgg7AK95O2xd2hfuZM
WlAdXjtmSL+fUhVYvAFlFjUrX56tAdg3SVjnWESV9jO21w+3BU5ebvN1mpku6+Fe
pLd9j6qGeUVimbpIW0FQY/DEZA1Q9cRXJEd3SLXlWose/U2T6R2MQdTH93cZJ6sY
E5uYsZeRWmN4p8TlNOrRGMcN2L6Aw3sRlahT8NW2qslWCkNNekBdlR89uK+b5JUJ
9jJqKCTntht31fVcnTnWc9AbOxR+2Yb5wM8520fwFoEvBMbDxVHeIhnRBI0ZF/9O
fxIv36a31CRHKxnnYQl4ahqarMIYZlrs0e8DinMZNjOLaiWdJMl2yKO27gHzbQYY
iiQB9JYTVF2ysNqX0z9ROZjs/9lFdDFqoOBxtmrvhAxQCw+dtJHJS0Ak1kGHw75L
o49qPVsgCswccr9ZcDjEOgr6uc23Fy+Guv7coWTrX5/4Y+uNcBrecXMp+bRxyGah
QOymRlB8yqDR15Dd+l/uK4p8KC/mIaz80nw3WRabpjGAUL9sxsGcAgfmREXxsar0
d0iUCoDM8s8juXUkARJROftsfrg2SBCsTRUXaDNZCsnVoaMm331LUum2k7l10NYt
2fp/VUQnymZS9fvoA2KQlSYNPRwsLfaVchRb96DVzYrBmN+UiehNA+F7yRwQIjuv
qPrgTwzw71Mf5Ne52uy/ttka+3XQs9hLNKhM04REo959q+BhXrWmwGVEL31oovis
t2VGPejNloWAUXADkhNoA8aiQIL8Kar65o6mG4i9dy/3q1kQzLAjJBGQrxD6nhBa
CY+IzslEpQCUaDII8gwlb0XJRbR4qwmIq3O+KlT4TOVgqsIZeSz9/2WX93zkOzj4
e5Ujs4Hnu6d5YAkaq9/WQsw3DHT7Dr/iWqSbb2uw/L2hSNKXquG3Exw0AetOivpc
B9B74wTKCtAn8hwr8sP4sLdRlXbfkoX3Ya9W2AN3WRPprVBsUC/tOZ7HmiZeZos5
I9yNVkqUeSK/k+N7AUwKHMkVW46l5+lb+Y8SuTe+/P28CC2hItrxSQ5gCeka3sOs
J6MQhH+HeuMWLNnPT9ZpnwgCQJSf6jLoj3idyWewJoTpEsEzq6CUz4dtJbvAi1pG
2YrYujn27fiSvuPsWOgKNwbQ6n6Q0Bou/WCp5hEiRBxpdduY2D5Waf7O+Ks32glF
TIqsMiL2WRQ5nKF7QnM3/fKAFJ1HemT/iAoULZoqAz92c0MuIJWvzuZLNWJ7hbn0
oOviw52lcAnDTs2yB6/oCZDQalVE3P/DI7GM2UbzKvx95sR2BuFLf1pJmBdCoalt
rvCQnJMd0FUty/zk9d/oMaWUJzxi2iGwHbWBxO+7BelXEGVFgwfaDOBIQqHfa1FV
ya1gH35ePq15N/GZsG2ENlwYWiUY8jsKnCa2Csj3+VZibbvMrOHjp+eA3Z/ib+Xt
mSs1loUhq2vcWfPv67WRxh4Sg2U9Yl8NIoR5MRn3Qp0arhJ2si+VR7hA9EpDGg66
Znz2na6iKCtOSyr9PvXhlcp9XO4O8zcU024FTg52ptcB50ZdKS+N5xqdJmdajSB0
y09ifjCk3ldW/zrD0TOXfpzxJqKBi/cCvxc5HZfx0W2mAFXmfYmzJRpAFzUKFPws
UIhRyGPmZEsWelGO99haBb//50ym5GKFtNtktDcU/95aAi8qRgz2a2sHfgukUFts
BftbiEBRmLp9mUk4pL1tgETXT+l3FIPh5Gn3pgsPFbzDWNaRRMEemVkFbj/fIn+C
Ael42Wo+MGGqqESXQilhlFK0JnQaQmELn3ObHvxmUZuyKnS0QkdplGFuqGpk9ogf
FbWz2MucpKY0UAaXDZTk66iDc/KP1lIlHMM+pkhKfNmIBzI04Y/Vjh8ivic5iMXv
99Nxun1La25vb/Q53m7jRFgyBKYwfj9tfxvdGnKCzzkcV9dnXTlnPjpiQzTqAYq6
5VhlefyZXo/91E9aAzw6E5VxusxdPX5TKQpHTD6tfGe5IuLZ27S/ZcL6L4GeZivW
ulQJCPZdNmPDAZaGQoObPDIqofwaVo4c7spVd2rJP54+ixRyFMiZR2T4YqTrhj0d
ZXQXzaXE/rYHNAwmnhfHdROcI4mKJtNDSzZCDzi0LXzJY7A5Ou1YTJNA2Pg5llEt
JDbWZo7zNJTtE3y4EUgsbv1fPjDhCZfvvXAK6fp6ENxQljGLDg3Ri8hig7av7eUL
4tW4dJ5Sf/VGR/R5fhSijZR1ZBiQTNkgPVazsbX1MsZdCkmDhsuQ4+Ncd1D14t98
pzboap84IMmxCpETu4CcSCoU72Jr94XcxZZ8tTt8/y+BUhe9EjydPwJbOcGUnC0i
Vi6WIv8Ef9kLt9spqHJbpIIlTAuV/DNuyD9D1Em1k5Q4dy0SB/7BHVOMF287SHfE
Ui0y60bR+V4QQ4lhdEdnwnw89MAqcp2s1w08LKHO7sroKc2ujaH3nkum+EtaK/V/
lzfSvcbvWEaNAgno+diIvp5ggJWO9TBDUyCDVJPq0OCua2DhYNj96hYBxKYsp0db
9s40y672U+Q/sR6FCs8QnswA2mr5loDr5az09QmxpbT9UB3/9NkOiixOuA3fv7I5
CrFCAoeR+g23JiH+BGHbHyFbePXSCy++jASNW0Oj3hlRxs6Bo1iWiXP1wSq6CsFN
mvmz2xM6aM5KN/PBv9oW2EV9lwszDSmL/wMeFTZSGeSRaHL6sKPnNKVKrkGZeF1q
H7E9N/DwUEZ3qWp8f4XwvFwX8rpxuPguY/yuc6/GuSyMzzvG4nt/2MWXnMcHnvLr
obCI/XjIsDtCR0OAI6nIBqVrnk+1QSPGLoPD6CnxV+QZVAEFqbM1SnWp3reGdp8n
IBa5WDSXldkkzbuV7zTy1eMvxc9e5OfbX82P0K0xJqFjFQ8AiveKXemFZbikpyxY
aguLoJBwbgc/Emz11dVe6gde5RFUjtrC64/9xH0yXf3yDpstRyhYaoG5XiuyehkW
t65mfX94rDSguV97m2njUKCQqmt79Ak/ndX+el8QPRY0hElHqjt8YjqtT2YQj5v8
/YwYeaBCa7qkEsIWgrb7yxxr0Zq4aHNCnkJG0QPMhmWtAPDfIPXINPhlqQMRQl8c
HtgvrZvEKb4qmO8mQJiRwpN5VsH/gvgEcQY8STIAsHGcUXhtCZXl7evgrh5gBS9f
OJa3gchgYDltmWkwdbrqy/KabSRkyZQZFxJJymRznwt2xjNUJ6Fbdf7ZhciOg8Mf
3AB9fKTupaurMOfpcOrVBdGddLCgqgr9WD7FGNJ5FHBfS7E5xr49dQPoFQRxXbss
lBPKlX4bIajr8RX+EPkzYsRKuJp2KRoTNo5i6XoLjwlbzSdDxvaVPjsXax9M72Jk
2cP3yq+PYHiQuX4GS8Oz56qkr/tRRFQQgpNFoW8fw8t5rTokrAwgKDMG09nIV6pY
yCa4eBhapfRIZdkj0YEWIFsLCEM7WvpvkRBvrMGetMJdDEqxH23YUBQ/oS2BEqMg
Kg+hMYfLcEBjpOAIOPq7TZX9YJsKg4AIG3H53Xtzb3tKrTbJ1NhIcQzBuDOy6yyf
QnJX40a1Bp+L9BVlmi0FIghzITV9EuiNOm9WKErS/eGSnmuIZ2qvthtZka309sc7
r6ayZZ/+Jkgnp0280sqnEihRj+dJ6pE815xYS+nIiDHdIHotbQQyTxqze5paOKJP
U3LLcxh0pKD+uPLz6CjGDoIij5r/OvDToXEYxelkZEikyqzvmNe89NN9/bFdojYb
TDnXk4LkeN1mF9OYFnhdLyQP0p7MfVD6/T49R6iSSOKE+RC/SRvdCOhUy2t/UX87
YpvoIrdkdNvPjOWENq0d3ZAZA15JTZvGv1uq90LOlpbcEpNY11T4nwBu+kF1G3uL
HRA4sN+UOt8vg5YPopacjr8ejKK4M36FQhiebCZ5qbOPHySExQgPXBvnJ+wh2urq
cjrSkSM4sWsdzSSObDOcNZt5KvbDitpduY1EHi1nCvMli7KFilbcahbOdK5gV/lb
XLINFlKXKqPcVjnEvTY2f2tuwsU7i+ce2LkG/IvpeHiNTv53dRSb7xHJEacQhjlQ
mmdhbuwBJVDUzLQp1qebPLTeCDgxGxVIPFs96m180kYDxLMwP+DdLVFM5N0K/cGR
DYAGHBVFJpLvRwSo5B2cDfSIVzkPSLFiDxQffGzXntoCPrbEXzJHVh0ONg6NiK79
Upex+SnYFnwmOfci5D3O35wELmDYrmWdJvaQFxKa2v0Wu/YNPZTVWeG4qjjfdhuJ
qCpcLPVfVYgxfg2XSZmZw5B4rZYRQ2gTRDvvPg+GmJ00xsmoroZAHJu9LgHqeT2v
D07ISupx/wfZe5bzkc6M2HNrZk0sPJYolrcZhtcBC8K0lZLSMf/rhgl8DKS+LNpV
qB5PJKe1fXbcpnyS1oUIoM67JUm6TdX29trnAwLpt0dhqdHaRTack350LENZuT8X
yB/bsV6Fl/qepRkTybpcZgv8tc0WAdCE8ixjC6K81C2z+5ph/p2ephkz9bYiFPGg
clnEB0WsL6PpgIMBCYXpMO/I+tUSLAnOHcB6sdARF79QLUrIRWT8dz7KJhzkCCJz
3HYLGLTiBsyLFKNDugMB/kEMAWncCyGKZOliozbXW51iJKmkeYUtlQ20a22TrWl7
I/8ZIPHqoTDeAwHgLz/8nDzWwQZp4cE/r7zqMIXebMpc6yrcmdLU9R9V46G+DE3g
Eer3V0H7TJO9E7stMnHpP0oJKcRfUOr9LtIZjCNd2mxGXZoaPh2Lh15aZ9pWg3Tb
vL3qMM2HEE2jAGjbJib5cM6YVAOXj/q4/KjjUHOTyTtNP+cvBWBnuxonf47dME0+
eBnQAzBSBYDojb9dCtQOboc5YdYKD07ag5dLP4/M/lU2/kav/WZgZpCLuv0ipGsx
4ssLAwISIsk5rLy2fTiESm53sNXfDBgh1/5LMJEteUPBX5X1KXCIqbuNTXDGNuxs
F44DqcsUrE3Vhn1yVbhOelJvmjeABD8dMjXdNDj/mi2ouFIV/b7OwNKGsTmEl50Z
VutKHMhkWXe9Vp2JOIkLVTxOMyoRK6ABhIPj7VFCLlPLJ0CG2NmQkYMTSSlT0Elc
V4zuuwCSy6PWK42NHzuAAUb1UulN3TdhqI088aTFNdS9nkBCwBXJ7YFtQjOg6Kwl
9Pxoc2nGK4gpr2+SjprBFJMlJRd5LM501QVLCLvlg7KLycCYwcTqyzGxnfGioCWP
ZNP3UdJOCMvziCidGhA+QTorAZK/o4a/fOTBj5qn5B0ctYF+Ix+s0NaXw9nKsHuh
if0bM8pRJQPlgimNPGm0ePpWJjnbjWSwzbAZySkEXPTX/1aZt9/cMvbNzkYXNQAT
s8j+OVlq06/k1YGuam2jX6qXOsHwA8RiQBDYS4UAXfNYd8LMumirQAVlekGLWTyc
Gj0EhmyAkGbW/4xh7wZBq+OrfhSt8wBWDo/UNPasrKHX8xYj5PttWL0frOvRzVzu
U6Tkj1dgpZHH4qY4jeaQKRr6umGFvdT/WgT48o4t98DZSrwpe5kWlbSaLV7NpqtB
HVO2hmv/JvRsmka3+z+IYE4TJxQ0K+D3NqPvJMsaXYSnoJ7jLmdIGoFXM6gsWAJz
didjrPJv1a7V8O27m82HWW3n0okUhJ674dX9kjn3BnCUngVfIM8Mzh2YYChExxK5
/yWu0NKaPwP+PY+idNTmgCVtvO8ZmgxMp7hDTz4dNTi4OkhnqfgoUk+Ut8+2GPAl
R9dtiQPlnH+j4kKWL8bBYMKHLXCLCrA66roiSuaCYo+X4kns+l7grPCLYhWwEb3/
wAdwDFT+qF7PEAyK8ON5eAPAQ3MOz7J2C3aa0Ir0yREvDEDu4P/aT8E1nGfTNQty
9CW+IQvwntvUWzvEtrcbYV9n+PdGEyR5Kmc2MihdzYhvKrqSz+ZSQVDWvKklB8Jg
7lm7xwfF96AnVKj+zZbuCWvVv0/Utc94XG6pZzf5ZgmWyVpsrfIbi19C8nvL6M11
tBQnPpYeetZw1HHplg5mRAtNRyCqFB2AADRl5ZzWabsAXjMsnBWk8KpGHtM/K2/e
7H3eFne8OPGzUBkhJN8LXr8C/vKnhnJSHFb/stOiEwDP1VOKbdX844MifQU+B5M7
hWPcLN8llKvMD5Yc8wtptuLfKa0qrYOUgsi3L1g29H8heItpV8YPwhJwWBPEQVGA
4snmH1qAAh2OZo1x3CNwdpHrUwTdWG9oD2a+RDe5a1WnG8C/mBdkdtmsbZiRW81a
rrUHz1a/cW07UlgGRRif0vTtdLz22wmeYR5mxBx6wCxYTcsJOiR3yO1pve1/eNgX
xEmwdX7qvYeYQxCxmABXPXFY+Gz0KZvmnCBs6nGNE12HUHHjCTJM/c+w0eRIl+Ac
JduPNl/81MDVSW7/TAFKZYoLfNivZXGXZfWQfydx5z1RrPkkA/DAygjkWzgZWZF4
VC/3yHd7ebrEUwrsPFF4Zl3AGpNAKqJSOnidygrqcnuOoTQ64xkyh7VJym3jzqW/
LWyuht4GXSt06ZwVuD2xIHEcVbmSSKWTB2aZo98w7ZZ5Ktt7nSWO0sFwLeCSGpZ7
ia/XQs8BsehWFPaFyXmEWQMWhOXu/QUTE8p5HFfY6c1DCRg8NBSrtUoNVJhDrzcb
fDl5GCoxPDQb/DTm1Bz9zzdU69CoECZIy9m9eB00RO9dDf0ptuAoau6hIplvLk9S
xkPqWXBcsG7v/JkdIw6/VGdBwIgWydKlEtSo3wsN3hsju2uEyYWjISY0o+qaEEwm
sf+pZ0646pnxRhhAVUxTq7EiK8aJvDEsfD5sVOi5KREc19lkgGGcRRxRWKLC5rsH
nsCPuDoyDESJzsPC3MYR/sCe1yzRg94STE0I/E1abuKwXZT4PnfCi4iuSpv4MrQO
g7tvdyuf19CBBIFA5D1U4x3Xd4hTOVsPg2wmXqbl9QqObLgpgta8aQEGRulfxESs
RyguVjC5biVRbOYcPy0jUmfbrxg2MpnfoOh1iXTuNvmPiNR4xlmF6gAvzv5zQZYA
/dLJJHtFNIRLde2vDcfUScWjf/5LVb37GUgoH4RunDIFiMe32MeeJ9WUXHD8ONy+
REW09mDz3PzRKWDOBY3cj2GPeVWvPSiME5f3DscD70luqIiPcSrpSbAkEJfa2wI1
e6MoxwCWIkWDUWfLtCdKgssRpTjAwt6NXkxuro0Z20B5llWFepJPXCfBjlZPgXgH
dNjATTrfpFrZ96bqvCBG5Uwqr0iyzBs0SBCZXKaiKgdhxs1aJv/t+4vrbxHrgXYH
x3IjJ2H0/DRDGUGhkXxsWCS/4YxLcHfJcoAgvC1ng3oINreFCmepIoPxERTtSWVV
XqqWoUoyy2lzhB75bMpjm22r8v7ZMC+e7KwSjKb5sEUezlc77zOuL1jcujmj99O7
dg/cY+/ibvaJBpnABCy+kLC6yOGP8FGpybhJGYgWmhUmoP787UjDQeZV0c3qtAfo
euTAz00swWmhdYJi5uZ0wycPR9TqOZsZYzET89dMrBe0uoJXq+YgJ6iT3vD4gHqL
9FWq8s82cCZ1lnC73naMg7h/FUBaeyKswhWs+hJEF8POsQa1KR8v6zGs9n5grENv
Jd2zt2rso50ODAANXELkbp6oAOixrcBjJw2Oe4o5LOkxRTKz9ctoqBsRoUT+mAye
lz562wh8sFIY8wg2Qt+1KmtAhtSWnSTbeMiHn4zZFOfABxmJZWRNMk0R4Do8ZZs+
r/HT0jFC2LcPQSE6ayAMfatnHh3UR71bqxkOA2w/Fm3KY7J7AevaYo4qVuZ+xv8N
nSxRWuvfXbjCyM9eMbzxfdI7ibdVaJBZqP2kFmvN8Joc8XPVmPuaWSCuiWT4Ieic
mujoWhCwslYySMewMFo7eNNbH0WiGySt5V0SIL+JQqyfshMGmvD+fGcgCExPerDB
WXZ7nc3xMPaEhum26tKjdxkVplqslfAeNdgqfLMdM0AizoPeSyhy3KXk5P3XJtU0
s0cdBWXc/RYA1NSLlBn8t47TXfTSJjPWfRkvNdQfICLyNGAWpsHk3O16jUtm43lI
DGPK8gZ0mI1r46A/xBbTT80oTDN7VHQEHoeIeun8UVcBR8HCdvDOJmPUP4zidEbr
DH7dvmcciM7iaJvUAFhSYFoEAFXY8evfeTqJrcRaIAFVIxCZmqWpMoqhq4iDNf+Y
Kuee8dJ+yRqj1HQcRgDFL9vl7MNaXGHNbQ4z0QwmBqh/JiLQbU9Uk5sQdg4Cj0fK
3lF4YS2WuPr2xk5AS0wNcyXa+DdgGL44tprwQb3MRGPYBhZdj2UfmM6OQsuDYbgB
q4/DavY65cG8i9HlhKyJQ40Nm7JLD4CKWInV0XWUc4qMZPcDm6Dq2erFUMHz9K2g
F/s00oihkgSwJYKOCH48blQotTIG3TpIv6PG+r09FpfRruX+HuBXKmeAe/bFfv5d
Vm65u/IDN18Sb/lhPGc0McrPiJNzmHgEb9rOYHAS/f1+H7QPOZIMCwz86dR8HkDz
eATlI7DBurlPjIsRqfYgk6cZzAhokrmD5U8xne2ZWZKvXFkBPBr4JA4tzV3XDc/+
M9mOeYgM/TwF4Kfa9u6Av8bCU9okLLDkR8im54YG1KAlECInoN0HLUP/MFhAw7jW
ej4iwQ29rRwgqoCiOI+pWM/ZgwHEsbvwefm+tINKlD1LFEwL5GJJMyHmfnrtzw9Z
1dVE56bQ9X688BDtXWVjjuSBxhflq8QKeg9S2uWcRlGqfgqyJPispXmcRsouPDAk
CxC40HkNWxGHyKk62MzTTwpSXBiWeptdP5gjSH9XciRtFC3gadhWimZoPhntMgce
dNggZhGC6eaTUnqVQxkEyVDS2gP9CBvLcrcM9MdHj5+u0xo7LdaQJqOyWRYgA3v7
HEWSyKdvrBMKsEDlGKkEtVeJ+mMSBo39pxQccRfldq4wbDgStVmxYhBTwum6wzBH
BuTeao6NlyD/hMwNVcbfWapbkCjI6tEmVJH4qs05uuRN3rVhtUgeorJCbQ1RT3Ex
UTWMB9AhyaH09ErRrSRebGO178DNE1L0BLWB6sDsZmwdpfGWRYSAbPUtKMJXA58/
gM28fryxZJ5zS7Uhase3RircNVhF39htg49AUTkNuIKGz9EgWXkIfqpBNWJu+TO0
+uP2zSq0wVE54S2HR/Pqxw8x1/wxZ46a0zgRJdpDRWpsSswhTNgsopvJ6cKglK9J
5biZX0K+k7pmn3N+1JV1IeY6Gd34KV4bP1ICHflvDEDO1f3p+9sZv80+UkJUEViD
/wJVkP4GD5JCHGw9GPYXMxkmkemM3qOzHKaeHmUTFIBR5bu3DZEiGB1gAJvxgPkS
2DMfQKantQItiBOF+52TeZC1v3dwKaR/p4IDcUpSlgL2J4EO+SlRuEzv+qlmo2EH
+BqwAOrwgp7Lqw07aso2XOFjyZGmiavNFvROHhvzbDwOrmq6lGRPYK2h8KgkJJbB
oxlFD+JVN83LehxFqMdjENfFLkpfYyfIVrydSVMUpQ28PH/LmhVR/plQ7KYIk6bF
ofPuQdFsIXURjOwGJgkg/O/nPgKa8QDRWecIcJQNdQ8FxpZL9HluN0zR4gtKrXvj
xcY5VEymr7Uq/NXdV9jz3N1ntXcwZzYW9C6HUBcpQQYnOUspMvw3xN+0Uufs0/G5
i9BReveC4GjZR1PZ0fP6w0svBGRa/69Sr45Y/Xy5ihscnfF/Wn/5qXvO5uZ09p76
ScAfybrJGRb73zQ6qrnAjjsfV5Kz0Tv8hYgJcvislmslnn6BtxPAcA1Ar+4Bogoq
JSQGa4/N8rUjzG+STYIg7828AQ/91uNdHL61V3nmQ+B+SXD0mYxusCGBXdZizILc
pIYOO/oY/wb9c0tpEsqzNPmaSMqW2+67XH8xf6Eqv0zDyy+kVAd+NZ9UUorSnUeV
qQj9o9jJW4PDz2HOVeuCzOEGF7OHLMRZk0OjcYGm8Ei0kna4PN064GabQp9loCbk
AAYAyJvyxoKh+69DKFAghzj+Ofr2ujeshrQoqTFqQ5C983FZA/99R/2WoOw5DF3H
/+FibiHnYxwzrjfpqVtHa7AymWzRMXEh5K7gZmZa17uCFha2oYNzms3mXLmRdFGE
424fppAfHJVBfYPp/bxSKaRf75X8qoM0YigwBM3k4SXmuCFzXAbSN5EXJO9C1zWw
6tWxpZNJXpKp3lPXowYw3wLWgaJ+Uy72ik2Fed2DTSprVB2r/dHn8TCClFUijsK4
DWNWq4VP25n+rx79S4ZnMGmaDy2nQVYTJaZSJ7Gjg4mEQ0MAsQU3HOW0b0evsWCM
mL/Ig8Of7JYqIJ37NcCEldsrjVf6MGBAA0Fwc+Vul07alROduENy1NnhBF+K9NXd
wOf8wZEszng0iUZOylWzqw/+P0+gKmhKsi1B6I4qgTRRpzMzqyUQooBCI+enxyD/
G0tIHaxdvN0kY1naPlWauILRK99rLSl2cPbfPYSkgVYIhIiv0bg+agZFNvCC+TX8
Rc2X3+x/y8OUcbZSrG/mOUc75AyN2M538hOpFMHmIP60ZVIofiSLbodC9nSliOBa
xcQnIVrAzO+zsAi5RmdZDMjQj8lTRQjIe20nuKSufyuM2TUzNtvD+PztVJGv3q81
zOS/aradYynkMkRKBXvu0fske9sW0a5ChYrg5vD2BlnFAa/9RaEhHBY2TbUEtoIQ
fph2EsyxnTkVjhjbK+OkmPUCcOepIwcat1zAz3UF9kAtOHGeeDZcqQiTshuWRbkq
tcjzRbx8t3/LLwWQSipxrjzhRx0Z3EEkmAz6UeCdnVi9U8JdDaLT3fnJAsPA4MLy
O48I/cpuNWu1fe7aDtcEdRgQ5s6g3Za5imzfjXrp2bUdXckHxqDZIgMigs5LdXBo
lUGmvUwVEnDKrLMJm2kc76PtvWRQaDOhGGzxAkqF8/43eHdrGhe6DYL6Ms5OAu+M
LU8CJMJglCGIUs7c6wCsA8ocUsd7tweIylBRnI4t+jpl+AaBNGvzppbiRMkiwBLG
ZwWAH34zMiVntm4DARnNKDW8ER3LEtr6SiSoRbsWOOt7x1Ru2jueotGD+gSCkYDL
w3stEA72rvHrfH86CdFmjYjCPVQvjdYr4kfXP51cOgmA1GJCafN2QyKiebksfNuK
LWtXrZDuPlglo77E0gxZmsicMZjqF7w2NB+oanNPHFhmktqzWp3tn4j+O7G75Cu3
OOOEtDyX4spo76wQjSAdSWYjS1AkTpuPto8Js79hbK/1cmXgekvMBff779Zl8zjb
2NvMLEpg2Uo/gj5UCH8hGA5dOr0I4OFO2jNF5u3gj1u4BK/MMbjvwHIT5Oy61L6l
R4245adw1F/SetXwatIaasKddl/UcWqnLS5fAXnfrRBE3goVmgE4nns2UPuA6h6e
ciM6SgG4//7AX8D9xdHOESjZ8ksdMxogrGeiwTxxES0IVSPQnhB8URK2yFIgAmvv
acayZD7gaxh7g5Bby6HAd4/MEfq1BZWRIBcjPWYvh8HTXli/ysxucdZ0Th1Gt7gn
d9YqKdZ5hWmaXvUuX2Gnb+ANsCWH2gT4vzsv5CCjmpH89Zwg0w1vz7+C1lQCNNNB
Z/vvq98kn5KRQ9g2ysfsfhS06JjEQ8RlaX2qGP26u+7oXwMiGL2CaXgcqGbHHkEW
OQv0NrvhI3E+Xwgo/tV9t7c/hWBS8087WbnVakRPKbpxEi8cwXZd9aA4tgj+os9s
zi8oNpsrB5MYeLwnU9LECdYQ+dwQz01whGtu8PTXuy/ybhcU6qPtLnL76WrHVzSn
1dXD2SSJDjGnmrUKYWyyP8Ds/1EoV15sBcQoJiQddxDW+UgoXffWP/BEcFCuzJqL
IKNR9sjlGqUppLyhjdvG3od1XMvgaEkZzwv7GWh0HY0WrIJe4HqmuqkrT/9/ECRE
Es2pl3M2AcXn8EZfmYBA5ob/YJjIwBxQFL9XkRdII5RV50C+MZPZ2FRxrWAl5KIM
A7DZIDh8CILhoYrrshIG1LFhjTWZ7XX/oVWKHiNxDGCka5kfZvj+/FJObyNH9+yE
G1hukx/m+3mIDALjzVj/tV0ZSc690UIuWDeuObzPEnBQUWd3OwdWGfK0o3Bx3l2r
Tu5VlkCdkrWWKf7xVvIUS6aaRbFrrR62vtLyZUfjVWvrJtGKbwOqwN6KEOijWb6L
Mvucg3dVC6E+Q1eCtPlSD6z9H7DMsYOqLfRnvHRBfEtA+/lrGaGA6cgH/FLgQNSz
T6dQ/rUWkJ/0c4Oh7VqiCQuViLbd+XaZQCdckKiNWXIey3sxEhW9gKc7eueukxVV
+bwjCkDITzzBN8seGKNU6BJh3eYrzh8IBjplharfdxOUvRQGUaDYzzVJtKNClnnE
+ANQ5pFbjMET0X37jrQ7RcW2wYp0i8XbuVQ8/LANSvas18rKMgbrkBSFd1xWRpUb
weIHfUX9L9hiPCslXDf6wyK+JBh9YVBbNPzr0B+U7zQtrk5ucRUePas59dmkC7kX
8CvNppEK3udSyx2GiXbud7lMx88cpJ5wJXhbWfsaxw57o5vR7ZSYfGPRyBZArP7h
kQVFXgZ7p14JX6Uv5Fj9hUDmLBrcteyjA0r3BmXuMjKekOjZLA0+lwjpOTyduKgU
C3WNLc/h+XlToTdfUjWtIo51bUGMS5g3698QwqN8k83sbs/LBV7yT7v4K4MWaPxT
wjoTBGIyxO5X6vW+MXRz+09n9irlOz0zdW9kWjMdRgyvtoej1JOHnmD7DGHeNOhK
v4KfmDbw6Owe9Ek+A2ZEHnRwPMDlhUmRAcCk6u3JvK0S4vSBKBJlH5cvd/eO8LYA
jAXgL0KCfF+7V7Cd0dlbREQSMOrnWXHYY1+Qi/C61GrNfwEhW0nlitCMyaQ6NLtG
jZz4S24JjURN27tE11lFukFoJD+s+rro+VatHiceHGiwMOUB3uCYrQ8x02rUDllf
WYLW5b/iA05m/jMSM9avBfxmAVP+vxvK9cVQwtFo6jHqZlDPza6Ylnd4zndd4g9B
lDiLOkssF74k83agU5BTlmV/MlmCKcOasYqIwwlr7FvrL6lYgxb03DAN+btRnznX
0YNOyg/jikDm2P0Tcwuw3RxpfAl9CqP7qBS5SAc6OEju81IBlErIee1eE8KHYjD1
cr5vPyNCf+vNw7oR7ccKDyzAlgmpi2nCpsmxf4TCffUgAnSk2FWV8BAJQ6XYL4Nz
1vTP8n+cSYBMuQS1hf83hhw3rPEY7sLNm62vUp5AVBAnxjBpC0QDSoEpdM2WmwsF
DCRYem7dj7hrmblTrmwOVfADrzQUb34G9O2uq5R+dbk8Mb0uS7608DXAc+LJp7V3
g146olYd1WhDmdBAu5XumCtF/LibLb8V1F2kTb600C9uT/8Q+KJthPpVMYPLV/7J
o0e4a2I0psJL+uqFUjTh0Kd4v04SwiwDeRk3yYdT4OhTT0PxTbF/qkVCM7DHSoAC
3eReVH2hH490sSeX1YEUvDXB8gpcLtpNchrQDnOQOS4wE2y46zheq+ZlBjtxu3By
4jvgW0GVaH8YK6aGOTg2KfDf+FLOI2pAXr0XmfY/d/15yxAPuYMCQoky1z64LfJe
KZBakozT3XMlxjgG2CnG/c4rVkfosz7sMtXjk9GQeayHFCFMVR1poZEPX4w9Ofph
4nX7yUkEslH7BwRqVBpIrfsOvH2i6hMIPl0hnxChIJY8rHHTN2Q+1DrZmByiwlpi
dGQt+zXOzekhtuMpEHlV2nlwQETccSKTJZ1/npRpQ+6fmNYWBTSbb/Mne3DOPEig
7RlAWwtVvAlvhvCaI0UdPGG+lNseomnEeM5sFPy1jSWhhVSRMmtilV6EP/iLQ/YM
rvikI81pI1Gk3mC+ioQaquKoblgXSuJTroxEONBhnwrKsK3L9A8k5IDZkB+G+w+K
Eyk3CqROIhuWz9tRQvTL8P5Ap55IQxXT6885keHkZbRS0h3dQVkIvj08+D/ayquy
My0A3HfbHBPObaE9aLbhAsTfOuMFn6y0O/SNT8biGjcaXciucu2HKYyEtWRjP/BW
hD+6ZhM0AWjAuBllHmCotX+e4fGufXaXiA7FiIIPg7qrRkDXytPd24HXyPH/xs+Z
rjJnXk7fy8tFCM7ioU3LBYDP8816EaRkVkbyaL0h9NlhbhW/p4oGrnmn8q4cyZI1
WE45uwyip0GHz8ST7Opbr7qhjYVhzzUkD7uUdyA/lufyEFFNggdYmvw9Aq9djPEm
VaboxZ2WsvjjdXSDV/zKCwHxHVpcyQbRchYU5SlpxrYXz2G6lFAKq73zLWapU053
m3xonRxDM5JR25bzBpkd1H49iuoacffWBmH5WIIUDlvXg7JdOF+UEsP2jIgq5sqY
E8IJXKDE5V40kuofgzs2ZtP7BTF6hO8oWnrn8n/6HmTcA3It86L3qcVyLzw6Dunx
YeKqXpEvGC+chKEldeOxRS3LtWNMl9BgkUsiNYjpLjz4LF6KWE6UwMYCANn7mKMm
3++DvS3UHO+NVPJ9/hW9LD//fQrKEq4lH+t7FCNQLvadpwu91iJ7eA+ds3T53are
12vj0sc4/YRyM/cc6Pt9QEKvMDDXzHiK9voIXAiioox5xjowbk27SOVaiML1kg5z
llYZhY0Q8NjYnm+Gp4l6kBnavAAHAKLG00NR+lGVfGfWDDO5TbOS0oKlYvqE8GjI
cwgOBDn3xGtabKswXbE/5qX8vWSJQzRFXh7THiZB+/+MqFKSD+Zv7Wa80LpfCv5E
VQAL9WakLNFNYTOreqW5YltYQJw5DLHWYHzVOg0XTXxM5eEKUEBgqq5dQqr6tmcH
LZZPD+Al5wcMZQ/WFZvkR7ndbgOiPx+OcaKlYMtuihkPOFh2Lf2AviIhN65Lt5Rk
EhcLBDd8iqcpRPvP/UTKkCfbEeO6lnMkD6cFvlS+CmGEKRiNQoZYXM++mcli+Qxm
29PwaRHavpZHbUQ8orYWBcHGCbVkcCh3Olgkj1afyyjZviTASTyWE3fLaElynFPy
wOlbPUhhcuoVuZwpPCHGN20GFEsWadFufqkGMHqueIkynhq9Nj8Q6o0fghUigmqB
7nuw+355zxfbdmtG3yKHw+mZygI/LD3LabiLKavI75S2EvqjIrmU9cj+H/05iCPZ
A5W+NSZUSRcjSORSSdxHjkLKUm+J7Z2kUdEvRYqqMh4qQFVwrngEihPutvzKQuHR
0TXEOn4a7P3+IipsHKP5kzArPg0zIMtSrAKbpXy4iQzFxbVgb7yeMBpnRqKG3WFg
cjCgpSx1+iBoDHuETkZCVZmekOiAJgIpUYgYtA/MrNHijPt5tRF2kcLRgyn4zqfm
bbVPYsGOa0mcl2os+N3E7LXcNEHVG/L6zlemwoZLD7to3wNpXer+VJtnEmVVVRbW
W6S1jUYKxdSX+VYQhHLls8RV0bhVTVc57fA0ZqsddMkZQBQ5asaDoYF0I30mot0H
ItcTuDn7uPy6a2IPVr0Fz8eaByLaz7Zs43/qrwzQrV7erj5TQY6GvKq413ehUBbW
77/ET1RsI2hH69tSu3+UewvdzrPBCACatBvBl3mxWtL0MkZD+gKkVhxRa705Z6Ur
NObVFJJfrFHELxPJjSdJyCyc9Z+1O1JdMj0Z72+tAxJpYGqkmcjmvFQHA7pYdMrQ
x6nOw8z4Pm2ZveJOYqWPGAtaqQbsZeHA8wr0253TIhdLsGbxYWIELny7Zcq+jwiH
X4LOcWr+nubSeRw8P5lW2omGSXA1XN6gHB7xHzdraI+j8+gEkdSUgY6QmnKMlz5l
4UdYzJ/GtKuq+oBbMDotefcXLrSTf5yKx20A5QvIc0ynKSeC1KHbsIRwCVUxs7yu
GxjncU5NHOb3cPXkXXWKb3tqiNLohGdG6k7bhC0EQPGTfSX7FpG5yYYlQxZQ+Ehh
T1kO2AfVP21KEki+sgF6XddolyRuLaxfDMCTtuuL3BjA0DGLlwjnoyusGBqvgkSG
XldKnnkrMULgUiR+snQnqE5vd03/0pEYwrwOx+yWkkucZI+iXLBcMZnQAg88u1Bv
1Rzoo97+oczoc/0q7EO1YeC8VRMFL9ohKgqSvN8ADRqKnDqmhBn7mVCr+D1sAq+t
FaDKT6sVds178Tc/TiPdkMOZKb3qI6GW7qQ8id2u8fhpZqbe4KYLJiY6gt0HuD43
dUbPJANi1vZV5JrvgYLBGc2UdnifaZLIfnfuAnVnzVoYGBYSVprTF/9Piy0VG7Lg
ToOiK/GLx0PtEThpAJ4x89qJBHWBJwJbES+dOf/HFtZnOKf+VhRy1yMGelrQ2fJB
BIEu5XYr/wcNeNkMAUUdjrvxrt3mZlqUgd18UTJFe4O77BhqAg4LreSXaUHDw8Y8
3pcNCWD7bYq3MlLBWrYTAxiB/gvUv4JtY3qkTsoZoHjhs5jnj+p3EFNbkLprcpiP
jjhBAsSL53xQeDO8M9Nxity8pFc0jJVltx3dDzzguHMvJs3uuEByiKU7EQxLNIIk
mTpasBWCfsImXdQrflx2bFOGV2T3sRYEQVGUTBF7+pnxcy2BcKJZqbirLGksEYmW
5+sX9h2Ko8G2+J5shaaPpgLbEmQQ83qEZ5WE40bE29rNiG9Kwq9erN3gtHmNLCAv
/BV9BcxhNeUss29XczietC4rvfMSGqVwDnx/3VFLJBO5bnczZkAMto1RRlI+I6AT
1oyqnwwHZtCxSBBeZxRSbZg0vau9sG4hVw8emW+ZHVEAonMMQTCDMoNXccXPE0Nl
E6eSuuTL0P50E9fcQXNdqTVSCZMqR4MdWEO3FwI4CA7hJ8u3P4fklbUfU+pmxDZP
Wjlxyh6Ovtes4VtuayOdAitPK/QBK8Hi26SzqLTWB8fR0gdYYQJcntCPTHlNUwSi
vmqf1esD2wE9qnEa0uZ6zP9JVZWqkxvnEc8I/3CXrAER7/OXXUrW8iP3cG3c4F4g
NVi02NaMFl03CAmKV++cc7OtUZc81dvYOsAAhYkJlEM8l87w81I0OWsbgSZ9puD8
ro0MzRLffgcwP6GVmx6PnsKrjQG4TLp4nRP86XXCmxKqX6npu4VcstTAdczv//aN
UxxNPjufF/xMCiCylhLMxyaSzXwEhSGhMlppM1VTdHuJ4/6MvNZV6eP0os/1SMya
Q/LCBWk5MpU84uwou+jL9duv0DY6QImlLCtb4FMMnTqlIeYVtjVkUuAkPCuoUCT7
cYUnQxAIHknEScpL0cRH3gb8/xRiDMrv+ORVkEGbDvb54zYxXGGRm7qZwX7d6wHQ
VQuYjk1L95zpwR0+tJ5n0perjA1/U2SGqI5VeZkiHO7DtkqtaNomIBhC/Y4Ne8yG
g5DDH6QE4MxgtzhMwnPXWLNrS/iOpUOWZaboFarN3UxQkylVXOHzGld2GNtxkGrG
/N33Qj1N47PzXlaTpMU46uOSprnvY7WfOL0AhX3XtdDdUTvYMRbaK/llX2KArS7n
xfXcWp4d2tFKqohK6biXgjbOvdKCr9DmtTL3fPVN9sP/CZ7zT9JmHQlAEy1e9j1H
77BhI0hmDMyxHoY4uSm+utwtoL8XHT6+itMoJa7jYPOire0uJPVJiCd6S/sMvOne
2vMfMbTzqZhF5YrUDxYCzTxxhkFYahWUvICqNF5Iikdj1Q8IPwioOT4v/VAh2LJi
XC5hPiF1ZWsQikXiVfT7Yz5mklDQR8j5dglhw5vPeGoH3qIWmoaLR184QuHFRKSN
UfKcDgqGNfXM/oCQZZ3ZQfu4g9VaKbWnSyYjzzm/6qkgHAwU4wkIs2pDvpAcUrir
pqHihNE/kcKRkV9uIc44D6N+LVrMqZlL3jkH+BjHmTj+smcuKqGKFXgsNsOglqQ7
qrW9CqT9SOrVlk88gwbpNzdw6/9LJl9NiKdDrIapnC/QWXpdf3p+qupYCZFnKpWy
AQKB5Nsl8nuVBuNIt7h+Fg961sym2YKKGo+69TyFn3l9xh1TnaJ9j6b2sllm8b79
T+Us22MkLLvwqxL4JSDBN7/MFH27kRF3ZbNrSQUBsdWuXF2qxN7xALucotHuBHte
zK9xQSGT1NW8G+3JeM0cBut27WmCtwH3CahPg9qcxBSQgErf/aQu/hxRJWHTDrjr
pa0aic/UJKVTpd4B/zgmImFqRRZfBq7N3iKRtfdcvLJ9aVDTHE3/K3YUcWPxF9rr
guCgNtZTou78Bx1gAIz403/ytL6kVuUdWGLKQsImt2+SY2XP80Lbx90xlJ/zt/Q3
2rl0zObz84ZoufIM/lBcn8l/UuQHBNqCLDxQ9oHjaz02whTbENGzBCjmEaJsuH56
f1ox1lJ35aJTQLK+J9XVxxUGan7+JPLcKzMzVTx5/Pqk/uitEd/3cy/UAnE7/3w9
e0+YLOaF3I5fEKwlxbLMAuCPFVSN4SwIJ4kDCYomqrmSliLRVbH3EbdkAKxvIqG0
EI+Xjy2BYrD2eT7BtwwNhZ64PefhhZnqvY5Iwt504hUquBHAKWl/Nq11UgdDNnUC
s1ygc8Y+r6S5F0dIZDLIKlfG8aITZTroFXUgteiaVzqxeg2ICX2nF6s7ASQigYC7
Rdycuv/AKzGwfnGPMTHurl+ID7NYEG25rXW/JKBKF0Upm6GCFBNKYP4zNyWRAH+v
opcHznLR/RteA6I/9jIoNDQZ9IJYV2F8Qlr2qk/1K3cbz2A2nPPQxZu6uVwN0Kx5
VPfXY2KKuyrWlD+SmxqWaBVoS+MJmx5mUbfed7eQpcew7qpBBGmPc3GgoNxVPh8Z
9RAA+9pfxEGs4iMKw45wQTPe5cJm7a8cXIE+LIfskim7gDroAUcbQKXFV4ku1rax
+x1xH0lxJoEvWxhbw6guj8ytfiRvE9RgifbDTniD2LpYVNbG/SEqyGA4qJHbf83P
YUYClgsEtfYzCoOCBSwiu369f3oSuIAZgF/BKZLHXS8tW8zPfoZ+ROglbqkApHMB
gpp3XBTIoRK6+tPZToCfaFsvK3AjrBCQ8WGqGYw4F/x+94BHpIYd/T5Ut4aqTkax
JrtI6wiJx+PlC/AJwuuM9QNBSeguhUghlYs9UWY2bPiDysjfBAQTjWByEldn8Kkt
Py15du4dl11XLYuUW2Twdkq7Z+94LtJ8fsoPTy9epwsNTDcgUKZZybmOLC4CT4Pb
VsCuERODczvMeMLrvcZzp9w5lDbpoUzg8KUBcQB2krYexKbZhkyfTaDA/mbhKkMM
dCmDaRftW+Js1LUEGNLL0c80XIm08KNPgY3eVR3/6LJv+Ca1Ho7NfPhz3DLdSvLS
41kDrsya3BP1PwDbcnCxJr9uPDiiFhcxrD4rLXqxoSpARmWP5pQKOtYURAsnow3u
4nSDi+kF8bSA8MXKTqoSKxAM/qykc9WlFRPmyKiMXGMuuAMO+YJTRQX0ANB2dCGX
otsf4vS2gsEHepYCOCvutFoeYiPda42ziCZKnrtDwr03shnmNAkQ/JL9JTQRN9j5
+bjmTjWk1HIhI57v2JRcAs+V5epTpr83w1/HnhL+EBeVUP0DfNB7HQ18hrkgxLKR
gjER5WdPMnGfe9U8r/tWxYQD7ev+nmlLD8nNEaZXXVbEpJqinc2+bS2EU07l0Nyz
idcY8EVsgR/k62UaU9NHcgK+nDkGtxYhMyUud/jglRCdllkxApEf8EBI3X6MvZiu
dTuuWnraBUf18+hgE45tOMa36Fa0n2HPCLJB0ygVoYQDBqdxbncN1tCcC3v0Q79L
ck0bjJ/puIvEFMaWvrojw+zgYVsYNS8zaieiOBLpHLJNFOi1P9R3NQERYURXwu7d
R9CTxzlRC9x5928ZFCfK0apVIa/TVDXWzr0GGtjavUXkcCxJzdBb6FXUoJWlO1s8
/1Z9vF0Wp7ap0E+QEmxG4J4Ux1kkkktPA7P83nGY7ivfu7AzhndqkPxlrmzKcydq
DE2I4TJ8NisjhfxwPpWZ7PHIjeDvav9LZb0D/EOf4ZCcroqArY7lwIdyaJcH7VDU
ZvD+K3Oy7/3PuI1aF4H3oXRJ/9G8N96WK/90l1ZZt33NB5blW9qI+8uH/9Lx5hV2
f+5RUFs/flOzoqQok2ReDenZlCu1HL9Tf0EVlNjszX45JL1KL1MrnELlRJLR/5zD
qRypdZyqJyKP10S7cwLje727kEVUZ6qmQ477Te382GwIuxufYhB+pkgBg+aTbQHU
WjTMQMhRkQTJLGfZ6dNX0ZGmIJ5tOenTDUrJEHr8PPqF7kfuutx9RatE5jifnUwu
o/UTVJ70QAF1zEKVoq6MmwiR/PEqaNAOZhtZkqqNjmEvapHgUfu9emiL61V0FMEr
sr7UK4tgpwIsW3f6uDoA1qE7n5EoU3g5uAoLq+SEhSLzMo+NgpEniYgeBXvt/ewM
CIC8j4ofBwitHf/jFTtENp0yemC5uiiVCVDVfYdbiN5ybLbfE7bstzkh1Niwk4GH
nuNhnpy0pWxCCC/NgddtWHwJwyX5RsT0m5EB0UbJXOcJsFRF8eA4oaWMLDdEECNU
OC0qpdbRDHE6loRg8yeZn8DER+kfKUyy+4QieV/+J7mbOO9kITOClAYR5njnWoSb
FwCsqpfQd2EgwelnQ7zyBGUe7XhCBo2KnU6OIBkbVwgOOC+BTP70FJBwluIJIiAi
c4T9O8Wz8gCuWbBhlgA78Ox/V9WS9Vmfr9Qot6dU6YErmW4ykF+dHNL7SdYYRJ8u
UmtXCSPIoFGcu8hFgX0VapwY3y24OAcpZWb8IvWC029Y2Sid4IippK0k6jPJ66Ut
ZlzPeotR67qaaeb6e8nCE4DZdE1a9ZlPS7cneZyEkxZdNbGjxgbFMKEXAjDiFJ7L
sQ5qkP9NneWmTuZ36oaLasbs9QDbzgUqEAUg/HcCxzVIo86nWFs8WYYkTEwUp/VQ
cqJYQwvdh4MSOxB4HvHYV6xD8VMfDQgj/FlVKNrnu2Cg8ljfiQ4VH3hKKC/4av6V
rYWGXN2dEun71WasHF6lZLzBnzflocu6QZk9XpvpDjOXclzmIy/yXZLyNzc9XB4o
PcBNFnZpcOdLLp+7mFmXfJ7SFNAP+P54F/KWD6GtFWCm0X5ecs9miwfZ9ScJuFN0
nCXBxSTH7cKtrj+eOtXhC/75EwE0lALsEYsfU3YvBwD1sF8UzYn8l2mLiVWhpJp2
3lk3APca0f8+wlvQmGChR/UiqYTY/4rapNrb1+XHAEG2f9OIazT98zOXN+7ZSJC1
UlZ5OG4sOkgwBS1UXQRsShYaWYewzad0/b1LBFXvarBKRtVrAy5B2Z3l+0Ytpmgy
Ui8DJse2cu681jhj8a0Gjn0Ep0+2SmBdYJI5bMrU7cD8DEz2B94Q/Tsqxi5RSVvz
dzvWmyUnfKlley0m/V1HPnxdHBK04+6l64Ha4yBUKZpJ0/mmVwjDvggSXMJOvE6S
qyPyvNr4ZhfT8Q4anWgsZJ87wgdoqiIgYhXf2dwd6ws315H+WtONLg2G4nLG89h5
bhQ6eOksq9lqNJxu659DciXTW4Ixmr729lfT/tglpZjI+xAkx3eO3a7JzCRqjmeP
AQzhsUknJ3CD7/x8rq+wH957FdzL4/rIBeumQRciSPeGlswdUknRWp4SCC0ZpYie
na8GTyRLaShw4sy50nJJzPvgbj3bW8OxFsSQoO5sGTVttt4lSLp0RihRpRnCFyZ7
va7/be1Gs4hMJq3P/ipmy4Q0TR5Elwf/tTuCkGTUxka1y6qrbO2Kp+JoN4ty3w/o
7gVZAYHXaIKIspKS5KaQUFJG4JnJYyQ3eMKdH9+H8G/D3XIZoQ+2yokB8286Awsy
n/UZMe3uwSTyvlUuR8LMjkSLhHUgXEg4hCNGXuArPCSFAzNKWVxr2WI/c79Qymvj
tw9XL/2gI7zRRtDOljhxQXCbiN4+/eJvkctszG0Yz54y/9l4s6LxF30co2BDJrJI
ywZvr7anRI4koxIJohhMkB6IICm8jFSbUJ5dIWJUEB39KlFgeEPwQMp4k6DrfM+W
6OJG/ZvAa4s35cEbf03yAazBnM4u6GZHI64ZC1G9zvV6PDp3FEGmuqj111OKadrf
tDmwGIgjOr8HIz/X++dmlQd92818+IRGoEdFQEBeCN4ZEF1lQKKCo5gfMSiRsyoQ
Ery8YjtiXA3Z0DR9Jv6nqhexrESUE0sgAZgC3LGuOtiFEb4Y+fpWpX/BtlkMxT1L
WI2CYW90uFCMX4IZcr03N0vr7eg09xBC/34HH9nvNRWhaa4/pQ/hO7nZtpQR5vl1
WJsIzwqM1KMN87ej+bInqEp/ZHILl7tnNdPwvpQWPVs3q1Qd86kbuC4CHxN1EJ09
0qxsB2NKlT4UlgWATcqng66puT1/5/5t/ehWC6ZNopcf3bo8RHPIqbWNRsX4xgsP
J6hgTOwLbzSpzy/NYEcKOd2eMp1Xh0h9MlL5toF1wX0aKCk+zuYXMwPxnPFKXBPM
t6cbwVeJ8DM1vLEBkxTzZRjb6k9qQ6jDfWQgY5+APQE0su0PVq4kwImy2aLRK0rm
oTjBhcYfQ5QUwE879SRAVQlOZctrgcXSsHGLOOHR15PodVEkyhKP7ROsWathb85T
gbXUyV0bV/hfy9/JZXu62TWyOfEfkpbZSQriLscQKmjNudnEi1mxSY5+s8VYjT/H
tPqVENY7gMkQYohfAT+Gd43eqkpg4mH1LwEr81BmD3mgc6APLp+cIq4aMfyxQ02j
WK7ca6kfT+1ulqk8nbROTaiqDiW3RTHae9o095Ffyx793ubLk9JXGgaMncK6e6Gf
Zg6vAKs7olMrL0w0zsaxSBv34Hpz8ej5frOtfPYdDSUz3EMeEBKJxTDO+NtcRsrg
J0hr84TO1ftM9vD5o22qcMUAoz6STtMwhgBVmuUxyBKZt6TpZwJayPmg7SFlzRCf
32HnfDgLqE8rs4nAfhdoat3zvtt4blGpQtNWaFOEHvo4RGj9FGySxIPNgyg+TI67
o2ZaXmqXHXDWD6bRfvutw3Y+MBTy+1gB3ImaKsmXdL8suIrhWuN+dcuxp+ixQFSI
YJDl0a+g79+U9rmZdVUJX49HGBrSGbIs+FUHG21WKiMWGJudZv9wZ2PVWqqEnpU3
o8TJo+CNu6XZtkCfBCf5cLNJcabttqY/L3m3nxfm2XPcoXuuDuXBCa615SXg5NVp
atN079/FqwEf5abkvVTpRzh/Jcdm/905hjG3ZeS9MaxjRnrZEyO5M+CwPNJWIVE/
itE7EPAuSMW8Ct3ierx9WO3E5woVYsRwG98hzYS9Kms+CTek7Xjzrm92R0IO3upu
WnPK21KEAm9SNyycKSOKithM7QQSrh/x8mr1uAy/LZiVSfGPBCfekOBUReXycyHI
BgoHeyfYbAg4XRmTRIDehBeFjkJum4efgNAgcWCsjymnBm6pmhXPAM80sq8os60m
muYacby1CrVA+uxePDLPlNGaCdmsFjnBDHVQSWwgrvNjssNMKVsn6iX0/vPYX6FS
NpazD25Gptiryci+JKVhVhMuISop8KOiF/klVZ73/g04Yyxy6Cd9Qyy8EF72Ih0V
OyMxZUetrASidVqJdeutpKmIoG91uef9q5IWxtyfO+PKH1+Z+VPPEKd7a3LPa/JE
WL8JKpymvgJhsk97ezy7UgblNXZzZQqS0RUnAucMqCakvb4XXzOV3WRgZQt+V5a7
JXa0SjHJTTegjk0qv6Sl7OJ5HM5itKpmN+gi0APJYr9AYP9tCc53wZr6sStiC7Nw
zJRYhJfy+Mu8eDjpKQjWDUW4XN9PPnDIx90T4kWH2IX9l7VlOiFMsnKcVmJM3bNj
apf3bbuLbgg0wmlpTGQaQ64rVjhoVWqn7OLJTPtkWFUaIA6P61mkXjJdGyDb9tiZ
UC9dbutpUnGOU1xCZY+uFujA9iJJ3w704vOfCYJQzmfJ5W1fjdSiQIukVwKi886l
Pr/Ovbot6cOxdGpVvOkIeK8FIihDb+phzg89ZTlSXlC2jGyFX+B1Kv5QM5O53ibi
fmHu+/6EojngbTk12CJSk5BgxHkZemhgz/Lh3MaEq583WsyGhc+S+62YhXIQuTvW
XKWHaVRjxXXrQhphH4ABh4jRNy1lLfNXY/qMtkZX3suPuA/5lP7fY4EMb5X5IYvc
pd1jHH67yYcn2QebtkoYTjbawF0XZ5eA/VqckxFyLiH1w4lNd8JSGE+4nPvazqx/
OoGqWDb8lsokoIwXehPCBE0gFsu0LRUd+NWHn5Ej5bWyRyh5kKbuKZHu2k4n1HAf
84MVKkQzMqdi5Z6BRFK12lc/oWAcmO+aWPjWNgTEzH/83lNOehRVlJnMeCaK3Rwb
IN9T6dHuECHKdjbiB89l6V+32nGTWVC65EPoWEPhH8fMf4LetXBU3ZNPF6rGvpVn
pTjvj7DAX56u23zhb4/20XGyG1QOqAd0Qtct62k1grH8Hb67R05GY7X8SAXIPFov
fUTT58c5DO7TdPo8OfdPkAhdBOYq4wjpFGHFepIaPRaUwk3CINm35yQlCq0I3rFd
5dshyymqvMb1ZCwT/ragoS5siKyUIDD63t2AN5BNd9MzODjqUSYLqkwjo9e+urEe
qrH4r2//eQlinn4tlYBng1f5HC4CRSF+5f9CCkru+h4oqv680noCmuS86nOdpVA3
zi9CimLvzlQLKlJ4DeD0bT0vDyn/MRE+z8uvICCq0NlJF4WEO7g/E4oiEQ8GM7jP
pDgz1zRJEnD85cMTXwfFAhrbqqGe6NiCR5pq4MUlgBrRE+oeDih6H6L5P1tuR5r4
oQeXit2S9yzsn2zjfk/8w5cjLFf50A03KCobEgiWUI4nkZZolJCM3B1l7CvIGf1i
LCfvxwKga6xQo0cNNoIzFmWDc8ZylA2PAKSUw9+O+23oCwcQ415KUTXKj0KNHq7f
eFXRDuiLsdBmkxFrhMV8/xbuaj5ROHJrDTOWrCVn/Ramw6d2Zow1Zis2c8RaeEgt
WyPypz5KhCk9H7RA+4TqRVSnUmEatzwypls3oAXBk0MfLNn+3cdXii7BPENZhKf3
+g1Je2Kl5kg+UBDnPjilYy/JKgVhSuTuNOQPNCnkjMYt39t2gkP/7KSHRsqFNk98
3gVVXARUfrFxRBLnYmO9XptM24aydufUasD/TGvOWXs7PSj7bcADXwtfM1DrITin
u02a5K+NtmDs5RkR9PUZtkQQfxWfAh/lYaaC4orLPKdKuTNBWVofKDlaRPAkAX4Y
AopJ2KKZJlezVZE1dHJG+y3GXTaV1KBzoGep4o7aylJ4YujXbNmTdK62toEtP80j
rRFtbJjiWirXVg6sWdQhzPUVZaDYQcm+lRVDaa3+6RYe+0G4X9BZj8s4RgTqcC0z
p67GBpK6i9AWGylmPfDwSjFyqx1wtmXA8PsHi+78Qq3Z7VgIFQiHhuff2O2Sa/Aj
+6ZWMcM5kK1Jhkw9WUe74uDhoXNF9oRH3257VJVbVre20l1IU5a6NMW1WWr975Kv
1anMJhNMQuMDrdYne7bhv0VLvMeaI50YcNDyCykEBakZupOVsPnrxQw2lhiIVrRi
9x7AoCbf3SPgq7czuslZCJMvD+hCqy8oIuTtE2RDucJ6bo3CVS9af0ZyAJvXAP3P
NZ3U9weJC8Et6DBlQHd/qHf1BRj12k77o2TUcDoq2oSfu5JOYUE8vBMYg5lem463
UqtXE34oPvxt8S8a0supT2OhBtVc5LZGPHwvfLIgkvGrWhrmod51sCPcmZp1s9b1
b00YOU+sZQdmGl33lGb9R0OCtzn9vTWd0ngmEP0PoJowBt11zsDAeF1l5jFTjPba
QDnw7d7LehoRX8h9TP0T8c+F9LirxTznUhsvH0ZqrSFGj49RKeUvNQ9J2zpVmn4P
Y6rAzpWxgUh7Ot9Xb2IxrHxIww91wiLl2KM/c7s1MZ6Wix8/nhtHXhgGh2Sek3lB
8mCriojoR097j+dRzWp4udm+w6ImR4jBWdpFAwDf6+s3Ft5M7tc9QG9roUK42gfn
X01GzkUD44rJanbS60NtzdUUjTmDl0Jvcke1KikRRJPewQsE4d3QWc7tEUuGKw/0
AsESO5+xZlvQsY60M5w7dg0td3DQczkZsKJDxAxdMX92HQ6ovMHqNL1fMR1T5qhG
NC8mmbs1346NpypgCBZlTEmrD1scC+EOKpvK+5PWydS4iJsni/ZH3WSLZ7e9lQc4
6bGpue1FNhbvllvRZienXG4pvVTsC2ePegAyq6xKNaKMP9oNC3x4X28u4F6GGAo5
Lz9PGtKmuredY7hlysdeeGe1w7aJVGeFj6ItDBrIVOI/+hlKu5KMSJrReK5OCv3z
5JViCnYoP2DfuVJb73LQ0BtN6KZitTYas+0QmW/1YxWAhole83nc2VciID4JYHHK
piUKyVrgo6je6wPCCbAOtV4tYdwGpVEnPBciMrNk+g/kMnVm7p8lbnyIoNLDSeg3
dEdaRoXOICdRpQ7r0fSLWa/P71MPgYPUAO9o+XPxru7angpt035KXVKhITZgvHcL
vXF1NAvBCgQJpm2Z8oKgP1jRiJsnuLfNDtnZTZGNYjyDSe3+4PgnVWAzWKBxUHI3
tixGajr8u38MQiWnCbNmAbCzQ9MrM9ZiV3H4L5ZNwMy0pOfvGkE0HBYmMuvtZhLI
1+fe5C4RH5dnv33t/OFfYeOgoU2gnxy22JXhosNUuNnmvTPI8J9D5kTZOsIZ5E6X
OjsrStYi3uqt7O3dPOw/r8c9ospWSpguhEHLg6BIbTWM7+8KJioOEooPFX+60NxG
kUmJsYOZHbu46jq/8UJOJton5Q3LYUnk3fY5hkUCQkOseCLHx3uSBWMXPCdPzHOL
vWkuHQlwl47EVW2+5oetcEvf8hRUF76kkMC+uVJ97r/1Qkps5HuNy8CBHqbsT8Qg
dj2FFdYepfYnP3ar/Yj7Cb74qZckCMCjMTacREa4JJ2HgAfnP+2eC6jAuDsB6V/l
MR8DytYKaxMTpX2YHWCKU85+oB1lp0u16KvSWdQslrWf1Mplnxv94Co3yg5kWX7O
CDbteaIV8ij+8IXNjog/gVE8i8TLggVLwN2X+1OLTG7QmR0bthjAx6dQpOFbl1I5
77GIsNcQcmox+9VEloxQw6k6ZPZMrwDRNSu1UeSJZM5tZPGuXNBG6FiEcAs4Rnc1
QwwHE4QAuxoUdPBvaemWL8WJ/iJukQxQfNNUpB9zrSqO8Wt9c7qee86AwooCPvxg
Y4mDY/gbYRoEP9BeHVmcoxNdkedoPCCkbkQ4Y76qg9oBazJ7DEL9v5Be2ZsqRshb
XuiPwY39icIQl3bCm4ciqw9ASwyEYclqRG9tJ7MLl/ODoVqJGBvpjnbPePBSlB+Q
GEXHMylrCOToxPLuOgxx3KKFdGZfjba3txiyCSkaj8giAZgJjjU8W9mV1xGVU5Eb
0CXS44h7SyyjpKVa5RPv/t8oKqK/o+2VTZ5d6ZaNEYOAm8x5uphqEbnOHMJCSgye
KyKlER1VPwQXYeWo/ssMMTew7utz5OP2e/KAj4WZknEt8ktj7++NTeaWJGtqJXlI
Kz1ub1jzTiXN6cjj1j5vaWj8npknua4DOpc1l7xold4oZn63n1LyYWXY+9ySQAgn
LE/GDZFFqCp81IXz8QV8cL3an98qhiRWpsXyYOrTPKPeOUuoVlhwiA44XHYVrZHe
u6bosCkUl6CIQuF8B3HM5u3GEdv9DiTxM9DrWpC2/ekDtOa+XI/VgNFT7gSkqLqe
goxWIvOnV/V7OU9SI/TbIxX5TzP3D5rCaxv9OGgqR7NdXRaaY2txGZI13i4Eo/G6
lGSdFiNdzfR93AE1vwr/dpv5iJnIL1Hj/TmCA/qzzF7GadjMj62Fm9KP+BID9lbt
tpbFos262xlllh5bUGwycksxWrpDbHyyFkFmjMw3+YEAYhyZsPRqAtY8hIzI5cpm
ADnzDyipoAbtigU5tfO1XqHgm01+lH2/EmCKFsyzkeIPZtpr7x9E3oEZrzCi1sTm
+fjaChSxtFd2eh4cmtXjLV88FH4hBbGHiZM3jXV3/yj/NKfsR9iAD5Y2d8ExdDXc
YXE3F19hHGAMRrW2SpekF6QYz99W4DRucWiJLD55Jg9Y9grZgAULMwGtlYowHTxm
eyB0EdxjxBFVAv5JS78SOE0dAIuledM753kU3SgpxpOPnl8Kg7XtABV3mJMdeFXr
maoC4v6I37/7FUIGvDMDnZ+blyolpQFFV42X35wlpMO/vZyT5gGr9EplkaFucGVU
55DTnHk44KaHODTQJCtx7A+EjZQle9rlcGVc30HyQ9lsX3gVmYyl2hBooMBoftwn
Ckfw6E3O1JeuFizIK0u8Vy/W3RGyrRjPMKVWRMhQUjqrpLry30kjrOMsuHcVUXCy
M9OXJYm0Hgt9xDxjGPWWnRhVaGukbvnzp4CnaBY0S3Hl6jO/H/QRtqpGoQdj7QPo
2nBB5lFLoVbaT6EHDiE3PdD29grS2aJBCChHeTSvrP+qYoU60K0DB5dK2a5gbmO/
b8Spi1eC1ip0lD824905npFBFfAy1OaxQ/XmTIOKTBVKDbvyS5+ovA2F7rUxRHU8
KUgAPX6h9ryv6VAGv+VWx8VWmBP0lzp5GLjskvozF3yAXgdgrvsIgvZsdoFjlgUv
mkNADxzaa1X8UDVUPipw/A6XlegZPZJ1Ny1Ca+lmZS5SJSTyKlwFLr+y91dBe2wc
chdyhKxS397Gvvhjc+HpJyRhRqqtC8+RMdPqRNQTj3QYO9vyffg91G8InZsot/1D
tAKU4Urue7CCDHXTGXFXjzvHDQtNXErsf/7JAHCHHyHk/5vPxPb/vDXi/0MzhJhP
5CgzAaLZxEDEYiuaUD3jTW2+1zJ6PjZ5v4E5ZxQB6gDwdrFXER7CN5x83jDhvcbc
JL920aaEMnEYrM//rveiKuqHiHP1bo+BDM4GSFAOKrpCYd8zUozgJUT4hzFNiZ/V
ISWeM07Rr/G5mztPhq8mw/2R2+xX0GaHUJhpOwiHFwYJ/YfxewymCrBmUWPq9Ij3
JSzD37kvGOmVmBBZdI/NyVN4dTlPhjpyawMiyp55chFIeIxPh+2XIJtPAFVILXYf
uyS7MWZogzHgAyEA9HDMfDyr8Vf3lUCUY0V16sPhYMWNtqfdS7FmSzdA+NbETnn3
w6qfZOHWtC7rcLvHp8nVfGDFAk9XIl4JdQlDCKfSphljqy64E688iFcOxyexMtFa
8/SI+4wludQ6h8cDj7X60gXAbV7ZtfL5QJ17w0AxvKDj0nHeD8T/o+6nF8esWfBK
N5yq4ObrsaV2IP0VNGmTzS+6TU0I07oFSsBYQEhoQi4Ujtqcxzziz4HxVoRiVAt6
7mAQR88hOmreImm+ZyJpZLemBHPtCjq8L+93Cws4haucz/rXvA1CFp9ziaae8KF1
iqlCgGZzZ7xIPNcryOPgIdvF37pfqPl9gnjkovZT8rBccs2gkglUQwfJolzOvULL
aeUxo/Bb+S1OrUlzxE8pZ7JewmvCcc3wBl5wMNOtIFyIDhHVRSzK6uyHPIUnSBIk
936HZAAWw9IfDXy0XgaYKTZobpq1Uy2+8p99+iXXN3p2N2FVFVd+zOWJaEDZ4UH/
IluGItTT+jbCGLPfDVdm6VckR7Rbgc/XEFz7jTFIvJ+qpOYyrVAEEfVI56pr+CPF
7+Xvvt1+S4z9ip1sghS8cTh32CsnZircQjXN1WlzvENdrxhqSllkXr51haDx+/td
ZQPiNpEudIUJL5jL2X8QnGOzlWjFU+URfKLotPl/QgHns6lfXk8MJLAHiD4O+fw4
fTsShEkdB4Y5bkpyXqj08V3TDJ9+B2Dd/y+ydHhWo0qSsfuy0+zY+I1ioKYp6tGP
9381fGCC81BYf2/gUh5vaHrGtJ4zUTecqLtvUy/OEjLkf0WfX3hTQrC01DgG6BBE
EqdbNg0dT0nFYucMCTbsjcfw3vS7JczVryZBad8czwcyfgLR4brOZiX3BY+etlD5
/iafvRxmCXfWDbISV47UzXmgoV8rZxE3rSrgIEPUMsqDxR+3hIqVCzjZkaJoyYSm
scheSpVnC0dTR8+NkjvyPiEeABurK2Ar77plMN22bTFBVwtzTny6DgYNUgYJ88hi
mGE2lwjLe7w7XsBcVPMFO5ZvcBZvY1+U69zrwothmXnIzQsIEnPuV+XAYo6j8Fkx
ehLxnwkJZkX3hrGrT7wZCRrsjWpzQFXdkyWBiS26+ws3rQCB4Xmc5UXMk39dE5XX
BEqAqEa9snIyC/8t3pvjiu1f1mAfg6NtlY9VYzfzQS33JLJIZfxjrlunJtBWcDYb
N5KkYU4eYM/b3EXz3h8tw914swezR1PC/KYsjqxmSNjyICqQA3g95iH0Hpb0JrSy
ECmMXIOBG7N3T7LG+6FCN6YgXzeyRQPIUdw97xG+0ezRV39A7n741AXGvZjkBUQe
fZBRQKG3FAyQL0p4a3+BFcshM8p976CWsi3ttymLoZ1e4QmTqLn/bSduB4LVGmnV
iub7HDFltGdtdWn8VSePGQWLQGvJZhCCmn2niDkDi2VfRCzU/Uz/LI0NO+2+12la
d4IABht3hTx248TXRKl8T1J9xBPsACeRw/2QjQUc0Vyg94QZfLECw86r+Z7Z7uE2
JJ3pakzD6FZqCAzTHmcUEKxThK9pUJM4xdAGc8xJjZsjRQpON0EOA5ICBpfLNJ7X
syXhnetLtLbS08uRp7mi5Ehr8vh2Zj2/J2U8T21Szj/IBjocdVb2BHAhd4ZaMj2h
0JA/FWrTbsKNwTqIGrX0Bp8ScXHriyYVNe1VS4kOAJCrh3yH3eNUQF50UDqHMVKi
ZfUq1AX7g80qLa/dHQppPnhhL4WD7vw3bIPPpnIt1o2bHk29VtJ/5jsmD49wfvaN
Z4GzFmKZ1y92kI3Kj6rRhHkRkvBcHFrHfAEwzSMKnZ8rXmvSS4OCw9O6ab+RUP7U
ntKfUX3rH6x4TSaC8yRy9mY4891UXoigxPeZXNuvtAQuV8u5JA6xrzUhRmmE+nRL
0HDW1qDrOaKS/+k9y4ZStt3FT+aBEc/DyuQZeZMYC9hPp1JZPmAdWRhhi9rWR6qG
pLFSFBud+jJoEfnzPY7hps4Mh5XM9aDvBelCg7LLeoy23qQGdq/IuIB8wil0Nq90
7r4ZgqMogiWhHpX6xZv+HlY9iiISKx994UOymwK3ZIjJSwe+/Q8a1h0mSRNZpBqK
0LRCAVagzqPLotQ5h1ML67nus7QmqfyGCAzW3iTP64MCJMC9PQGlQnJruX+Tiu8F
4LlbqDfOgwyB4Du/2kzV9D0jsSEMheg7MZnobcTtI7fkSSSAyGUgizXSZP69RuNI
8LBTFxmLuKrogbMTN+vNHaEsrn1ZjKh2aAFlJzj/8v3tdqPRmOL6Vf5Hhg7zr1wD
qakzcuTCITsXFbsfn48c5B96xKyYe3QPN65x7B0ofCCyzpyyh2LHsb3erYALaevB
3zNdqq5eqWc3HkH91KMVLWszHMhgeKeoD/E2fCDubJ6h0InryHRskPH57aUfMYKP
1KBvyJFidMqy8u2RrKqDB6I/ML1raeX7JXoPnvm9U+uTFOVWwf5ZjNYdjbWIbZ2c
UjeMy6awxqPV5/seaW6kN4pv4byCDA6hAx2HrEN7J3C3Z0rQgbAJUVZ8SU1uXZf/
SkCUlpPG6LkgOnDxsYOamck8BI7QaYAe+SSlmEwEJTkJy7Xu1Mo+SzYT3Dj6CRry
5OmZjfmgXQjvs+7j3byI5PxLSTMB5Yj3B1a/wWSylfc6lDNahSF+tDOsOaip29lk
qJA0Ka3Z79rM4JpB2ssWq0Txhvl6dUiGFciz5RdnETm3NEhGr5M3XvZOCAPxMGhY
OJbD2Uh04h1LLP1FlWTolAam9yUiuCKNTmNOExmz4M2rErYq+1GsCmd8Ab/Yp958
BP5Ig4p4UFdbjM6eZxYVNMXhQ1+2u0afhPcE0WpqgCm9yUlG4uF1O8x5Bq3CG/ko
lrqQEJwySMxj2V0FbDeueliA/yGZB3yFpyrAb/epevlm1+sklaqBiIO921WdRtCt
6k9Gm/ReWRMUSFLKIKZCeSNHL8Fyu44S5wDU7iNKk+Ub0Fns5/1d2Cn4lmup0xB7
FaS6D57iagfNriEMFw4hgHK6ak98tdwu9e7c6mZS1EouxsoCKtz7OK87Cy799hbd
5IU98IeIngrbl8a0447kzcg+KqVQI5f7jZi7g9aDA4zsPqHUc1HwfkYy4WlasURP
CUSDPJ22OjSLOy/Pv7yZwPV8kh3O5OTaC7C7C4P0ADsODDCqPhxoteHGvf0qZWMx
E79ta10Gf8eTm1vuKRGNAS8QdWhuOzEpG1ESoUCMtJw+C2xFCJSQsitLbjnAsOgb
4zQ0pMC7223gkt3BgXoVCfDM6gwOGQNAGr/qO+6D6IGn6EGwc8dhUgRc/uQX9ZrY
YfgsYJ28xBAn6eEU6GF/yXOpKaqDYVZznUgiPHn2vgE/lTdq9oHR+ITYRj57aK3i
ucZkrb7Osg2zkTfg4do9EwEzfQ0FkLC9ar6YVhTk2RtxHrKgvH+xwyPQ6HDuGgv6
mw6jIhnjImsUAlr50POHWiBljVGZOaHyJ26xqODR8VfzfP14MuQvPS1Hpa1EMD3j
7e3LYb3UJNFSQKKR2+bOFWRq4snBtaZW2Sykalz+sczBubVijyjX92ysNvlSzSDx
XWO48lCBKBQq2lBNx65GQAbT77yZvX1GVr0mZU+y4wHFruQY6Lt82HvMjd4tebgw
3tS5KG0YJJUVGW+EAKUJ6wHFkDjfQe3198txV2D1uukoAa2kbfxENRIqBRV2PWS7
PyKpHYzuSrp6acW6xzstS1qGVVc62u02IhB+1luIY7YQPkDAGy8uJYopiwX3KQjf
0mx/WbORjrNlc/1EDYgSepQJ2ecR/Ldo7eIMOuHn5RF9ngSLIKoAkPQS82Z0eOl1
QtlSdQMLepi9yd4fv9i5pip3Qk+wEWv0ZqjwNlIWixjvMCC5Rzo7A80opYu4msyC
qmXInlFgHx3UyRQ1xI0p/oHQPbPfE++rgpkvD+87ix75bsF77Ri5LuHnm9QYIj/i
cuNtRgDryYuyWFU4XkwEFCqeGFcOttK9+RnnT01vIPFXu1ZxS8GefFTz6X2gD2E3
vmujWP1ldTmgdfW7jGniiOZ8NrqZqEK/P0bIhdUhkThbf7zgJGVwzfQqEj2OSJ2R
5mhrTUTphi/PMeteHZi+60zdQAZULE382pCd69oJlS3ldI2KJbcGnanVmrMzmaUs
mGXkMGtlrL0sdIwQhapxEqz5RY9OtZ7qL8fbvfzVsX2/0yCZ+eHBDuemNXvPia7c
lUjGBUWW1tmc3Gw8LfTt9iJg9YiFlyaC1nZXtYUMOU2Z42Oq50qxXysnejs3Fn63
v5Qzp9TbQg5TUOVQdHx2JGjsGY0GDARAU3jc6+vVQcUVes78XGxw/kvFqrp4uYoK
c5HSLM1G9v4LNKADrLjgoMuBX4lcyumsiGbPOCTuHqy8T3VHDDpilgaCuKIdF677
1funK7QZVVKrsn2aI0aKreUIiLYEv/GlzsDQDrT7GGpBj0G6hBNW6BWw+DR8Y3HL
mS+/+S++CD4Jhk1L5nU3LfnXIVp/bMHX6SA1bFQqp47krvY42I8LPqnOpk3Nybk4
1E4+kMvqm+aDgx9BYDuRv3n8TJE+sX4Pvr1CSa1U4c3Q15p5H6WBBVqOCKL0Mu/f
rOzKOkN5EDbqXKf3lyww9CMA2p0vxwitY/y8FPtVxbY9tzEsQ2pPU0vzjTAXAYAa
5GQ2V0B1b8Ii+3LPJstt63osKCceMsjfAx4/XIJrtVEE/RfTlQ8VPC5TCPXWymv4
jzOis5ooQMgsEss2R4oaT7JZoiOQdbCulCkln0rtg1l9GA3H6NfkPiFAcTUFH+Z6
paTGR7MINCyoZA9MQNX0uZnuiaGzjI5XcMhjInsDYrg9y1CPvERqbku4xoScbwMD
rOGcdDjt3W/8jLY5i5I5LVjsjxJAGQpLWwhgpx9oWFupKTkgqYz3OzYiaIa2heL3
h6SVEOYPwf01fQ+hKTvb0M//yI/5DYXdmTp2GJFb+IE1RyfvFXfb1bhBFaFepmHR
MD4ZlPaGv9iOIeQO7qit8I7+nI7HbGTw9wALS9nayVUYPEbzogEN1HsCCGgvrhRo
ZbcB4zm59jn+sLqzKNvvHEf9j0dUnj3+rny6c9TQOuJh1Tdb0rPLWhhn0NiFzA5s
V5mUG5GTph0GPEDnMffbxHeXB6+f8qagsn5+ecENPtPMlkTPV/INOVo9IptkCE+o
I2xKCanwOSr6oC079sanbSjj/Pb4hkHqYmqn2+WfGnSzmguqci2OwWOCfHFbUHW6
1RT/Xv2jOYtYaL47FsHUlm0RyVW4S2TwRc53YVwJv+2GniTG45ND/mPir8GLzfMw
AmKSWrsBdraMta6rMzXU7NF7dXiXlQ8CrMaYzWdiFtZARWp4UN578OBI0NbFA7td
OiXZ25eDXvPj/BCUJyauRI3FfrDXnwrCPjuQHDjRVUDtwizlEFnvs1K9XQO+8J7r
qlZz/QfUIWD4FtB9OVu2t34oe2dtBp/j+4He5FqKJ2CedCoM9iTxGIvqUUc8YLW+
YEZtpa18V/Ch9oxWRTRBPshHDt16Iu9MDNe+IvamG21Xp/gx2h+PbNb27r1JHSaD
i2Ld9Tzf84PmNm9JAXzvyjebIXRp5lAohgXd/UCCuJiH5G1vrkmwldJ01GHH8bwF
kd9EgEeGXAn2HREevmAtXTAuJGissCmP3QCFh60Ss6kHboTjLptlwrWOiaTy9hEU
sUYlzhqavKGGb32DZ+fTcc0heyw1ingz6F3c7ZDOeYypKsWHLPiNfL1vSspXPSiQ
c3UPk40Q+avQLpy5AFdyg28vBXWjrcTtuxsn2lepNsSdSpHS2rDkabZrdQIQZjZJ
IVhAwMG3Kztz3jX0tF9pVqGFtYPKYgp8oQOPEjq83TFXa0Em1peFjUYLmwLeKoB6
nEpiWXd7YTMsDUf3EUA1lQF+ibx4kMpehjcqXMXiIJNMa4E8DpucnHgWxzWmvHBh
OTcfCFXjHwE/eCZwotoO5az1V/CW1+Nj5Ze6njjP1RFCmk6rFn0tHqwp1Igg79su
psfQLhyvXAQ6A/xMqx60B7JSiJ53Ce3V8CklAgg4FWgGV1Kf7op99K1Wru8MLVgt
dzUwMqXIFBmwgWFeamMI6CpZgJHN6XHT5XWwaTFwVfTIrunZrt0V+Ou+Q0gtWuMh
jqU3wPGC5Pl3jKZkIiSVi6HPpm1kcMaAOJO10OKODme/aMmXYj0l6QysmGmmVcAp
TmP1XTVcDss+CeHKeckd8mZxcd2DaIoENwBMoCo/U+5/Y397/et5/ez2QoO4BDXG
lSy4rr+yI2Q6g4Vwv9bInDqj97+FQAC4XgThWYdFeKeDn1N3qccnZ+63gXbqpXXJ
wZuaN1LV/kEhNSVDuuhAPhrGRdX3k+haQ4402OR6qyycfotCkOD9cCerKb2gWElP
W8ahMqIDd+hRGH8JS9I44T2bbiyyeTCXk++Fk1mDpzQ6mQhlxfUR3yHT3Ts7tcoM
nNFwsHYsEX1oVphSAmatKv0eSbkxZquhk4EluE9nsFINylfM8k1TLkdBtjTeR451
q/0oToNlosh0s4sDE22t4oVv2GKnpJBPQc58xCNMNZuyWDDwhMAGbDr4GdsX6kAP
niXD87N8UUhTH4igbAHEDLO4kLFiX63+546UH67Fjvbgw/vcfnKHONIXzEXTDxp5
iQC5Ue8wLV3N1DXyofiOtB6EotPXNy1lv1iHvd9W4V0ILgMsRaDjlDQYnZY5rr+W
Bq+t7r/iylEoyDwrKPbFKPmprnwBS0nBEOvfymqpp1DsWkDcrEatpiohtkPu7EfJ
jjHxH+hlzKTMUOZeYtySNMdVKziB/wePjLmGGKciAk+ME7sOuFbtv+SulX0YdJaw
b81jqhvjN6CxwauXI9s5FluTgWTFS64y3Oh+1LtMGXQERWq3oa180+4OAHOdD90E
DQ8ImhGU0KmJdds5+TcuMbFYqBwsEXK5k6aITgZ/Aj9BLK+w3+VeAUVre3xtDVn1
h7WxOsac3TyJi9h+uYdvr/CchvnRbUo0YJlnN3rNhlhBzSxs9PUl+aYoxeLbzwmG
3oGxYENsWbr3/rYHRckip+1G/hqZTlZ2PQX5YK5KBsxgGYG2cMjzsnZrjXdpVBVS
/cqGw3a+GAyKxlA5J59/8aLP+JbJ0OFrXsj5nAfg0G3hmYvEdDQTTPnVfss4YKJc
jQSgyMIKrW1Ma4C6XU9bN4bd44m/H8V/OLWdiFK151siXUH0zUSjUVtKbQjLtWW8
Nipfy1xJyjmqFIYzxgII+xeUZ44+Sll2uOBFS8H3OYD2DDX/oDKuIDSJ4MDGgXc8
TtbFBblOZ2unre+tMXl6v3gcxFN5L8sbkwYs2PMQqOZ5KTXKfCqYTp1yJwR7Ycl7
Mo633dLFzP32+ivhHooG8KYSggYobX3uH2RYHG7QBM1RqQc1eEErK4f1Y55epTOm
G6cxBXa625TAUt8W5sKei3z/Zjt4zcDBQTbN7GrceQ/Odo6KkMCeKWkmeOjN9Dds
e+NbiQCU+TuexlV5Gb68RJRYAgBzqsLATiw5rmneot1rPWEBhwSMh06VQv+I1wDU
OFA6N2E5j/OfEz1tNUtYceMX4Y0pd8dfmV4Vw/d6LQOtQD/M2kDAanJ9jmE74FKH
ez5S8ZUQKcDOFEadpCdMyi3DEVw2wY09pBV3yu5ZNf6DXPx2tSZ2Af3pDyOROkQa
lPyi16x0gRR6O/2fKrd9bPnC8ALZO/9USdOlIM2nh6NaoIl8+42LSwEJnG5K7dL4
nyFO1qtL64iH4DgmXrdc0u30PxyJrOdyLT+t1aVbaPUfWYP1pjqGk7DHQkr3x8m0
5mvMlE4eZjpAzWRt652afgyKbq8fEtl8DmfMpW+htATNAAMNoXEEzhDtMAxkhhQ9
qo7oHdA6KXitEXZLn1ef5NN2jFMmmmij7rkE/DH84EnvtShN8GgSAXSTJX//dGqf
gTw6nwwg0rPnJUy726q3HvEEONtaKyTKADqESjL7Xfk6WtLzI1XyBUrpGW3Q5mX8
9zxZZiaNvfCp7n0wsj3zUmbEuLRSy+kfVUKSlOwrHXVkR/s/rxx9tUXZIWLdEIrl
SqSSvXFEPGs/h9oOAXHhJYD+K84YUeT95+RpKHlJFdYlcEVIA28OJDkyYtOnCq1w
nE9FGs1iNaB57nRj5MIaHgMb82F/3z8YVj3K0k0CQIDi5NCVJE6OOatt994h/NIK
Q6Q51vxiwHQHk1Wq7SlDseqVDw8yA+c+M1/chx7Tzh+wFK0SWGbQno/D7kjdYMcT
FCpu80WErDJHpz+CSVZPo9NiWLXtaD8LAhNiSbPPffSqjWuItBcoMxdNFj9iJEwT
OsTv/Mus/HpuQEhXpW65tuD7pZHg8VnuHUBkaxur5TzgdM+UCexhIDUDuL4BHxIT
wsYQ+W13BxbjHG9svvK5bEHvXxV3rvoCC53livlJK4XyYWcu5HDSXpwzpKVRQ7yS
7RTFO1+L6NdiRbNB3nDVUBqIBYsE1r7iZcL4kajHWnFGSWmgbxXrVDa8pgpCiCQS
nx9xt9A9GH+7LY6q7PigjEm7XNngukJL0Y8VoG+eEJCaGPM4meDQS9nR8l8XPzmv
m4zNjUI1bGjcJyt+1FmnHHtIE8eniAJcxKqY2M2BqyuomWhJrjLzEoyIDwA7nyzL
z8hvgCyx07KEHy2MMUf8Gs3pqs04pIW5vmisYxaXNcz5XOOCFWhZSIGT/zSkN5kl
X+K+GruGPTzM7QF98rFpbz1LB4c9lU196P8lRVRV4Lm/H85StDij1TwMEntN3+zo
RXT5BFLDTK3U6GJLqeUhLp84aPARcaAT3ntZ5OMUnWiQV4ZoScDly+LcqvZarH5Y
LvT5pASQBPJPkTSyE4rDBsRO/2Fzc9kC2ujw/d6mNmo5Hiyob3M+Zz1VmVpRGErr
0O+rl2qqWpVA3QdXizdSM+ns0Nms/Z+iHoRVsSe3oKARuIG09OaJFprGYjRDZCF8
0UkV91HiQp/6TiVlMYoTx/Yuet/EeaOZF6hvcG5kK9ExdIaB4yBbkljrKhFFzFnv
5GykELOJfVa4Uh4TE3b3FXcdlAXN/4KGFwmYtPxhStaQIwCADD+LSd4THvQ/Arus
oxMSblbI4VG8CtK1MF0raA8DvsCKnJRGFQhYdFNXl903fma6Zx7K96USDu1BgjLj
S2VMQz5XPoiA1sR4A6mlRun5MfEjHWg5ndF1ZsUMw1YKvCXVcJBquuKHGUYzf/O9
JUE68HLpje6fiThYCBhgc4jd8CwEssPDlp+SAGNoXiVcP4CQcPCn0FspNidViBWe
Fd9UvhFRWDKCwaI6gp7HWYL27yk/BH2GOGtPBAeqF9QKEBUId5lyZ26iOupNWBGJ
kqHZSJS76kmHy6WTIqPZVD4XOAuQut3z+qvwbrHQFdQ/1e+ippZjfdaL83Po84wt
eZ8qLiWLdoeybpSlm5aqCNSAsc0MbCpWuBDH44dNBwvbLxoZKw9TnPNhGBpJFYJq
tyGzJcLo5QpNQIdsp65TzvB69HhRbWpqEglB7hUfK4aQSxIb3fZD/Vog7SyARS/7
NKWQ3DSWuuVua1M9irT1AafQE+sT/ujDcwjXN0FQ2EaHyFvxJws1MIUOAC6/VWJc
Pf9uVqa1EYFPwuROjcayOGM7SV3c0d9coOZKnsLw0I6nslRrTGKZ+vCjL4Fq+8MS
2f8D0Jvdv7t2WjcPXKjsq1S1XzoreB9oh5/p9crbD30fghiNUY0qgMcJMx/NbQMO
fEI+b+vYhlEfnyEkHISBpbS9pKA6yhAd7IpZQ20HhqtFYsZeJT55f2C1VQELCmHU
Qse0r94tbMHgCYe+y6isX5yRtbIAeUD3luMmxGHkz9u9Ty857lxb3pZXttk5cwwi
ZMjXInKv6lROctRXKYO+mmT2t14UnBnXtyauMcMlA1u+iXLOoir4Xuy5XSf4Q3Kn
RTPXX4q8VIsE7/V9zc4PwAnYi0iTlisDJmnmRYF36RjeUS+uyXpXq5HeHIbUFgYU
NL3zKXe8pSB79+w1dwt7ECfmgyZDGAyIYtZDlB8csYyuLi/JrIJbDbvd8sknoboW
nv/Quv/qPtRxPLuut/4H5GEqpEfC9KwD2jorPkf6dnwV76sBM1Djx3ZZ3iEf4Zn+
0NcRx15yiGB21p+BLSrRJs1JVYME/XvqzsEA6wlZ5GDp+8J32sTMLQs34/qKIQBg
ABc9fdwQ3F6RPgUK/vPUz7zo0Z9zXDJZBtlapCt8srxOmQSuaF28JtoCfjVvkbay
8SHvRQWfMajDE0gluNrgmWPa7T3PSBZRssE3UUZZ7BruPFtaUeFywB6pMQnzBQsj
VCeiKGR82V+hB8pSFvsF/8xY/x8SsjgeSw04VnemiNYUSnajtkD6fqTsTs4dr0jo
29lx8xhOUtsEjKMuCYefLnsRb3vgAlSpKolwl8uoOMaSlZQhS8nrzMNON9RjZTu2
XhiAKw5OZtzFhT1qnrtrZEpDbCykHALhGqZCas3MV4l8WVU1K5WAFICYoj2gvSpO
dV2limrD0yuiBzFLJK0Sbtds+oHqgsnEXIqtyEQhYf0rX9R1EJBSQbRxUGnVI0Ed
pPcfH9ej921hmztdleQ9WF4jn0c0tVfoJEMNyT0Qt0REAtqiHbXpTvE2MD4mOG2h
+O11Wj0IkznuRxjblqlkcGLEilqR9sbEbrkRVrCtyL73eiwqHtTdGgcF2WkZkp56
nIjwQkLpOVYoDZreUf1ktd97d68pUo8RLW0vhpGYZHh4vRwQCAF5PnvhBgaF6Maj
R6AUFLqchKRmdK6f4uuMWAD3l7AnaoRbFOoJ5k6OPofo3greSUBwvajauKn+O1Wc
yL3SLJQpcQeA5vXBFmi9Ij7pc8XZvDe2b6jnWj0bq0/iZbBnoCtHDryekuF1fuoK
fj7K1UqhDbDqNMMwtNgoomJwsaFZCo1coDSB1/n/aUJXofFk1mEMuKIzGROtGAjn
ggKTZxczH7hxCXGAZiI6T/yeWJwECXXQmIitRLdUpq/saXiQiJEhHbwtLcDl2f7x
FjYOv9+Cgyx5O3Jt1fpwyCSkc4hU4ZPSGad6ryhNf2+mEAR9ituIsAolmRDyF63Z
M3smjVSMSkmugKouYUkcmsROtYYKiSEvNfOdAik7ff/FAMNPB/ilxFsMPLxoM9R2
efyqrySZuJHUtFmfokMrleje/hWIrJoOsLd15iUzYAAdk6/bAvAXppnsOi4+at4E
T7pU2CTh3EqamAtRUkC72rrH87RGV7Ib6TzVGqjEHyxBpQGtJwySLRHiO9hCNjjo
HsZykiX3cs4MfDB9LdgDpiY8GWSL2OAuJ4cFhzmPBVs1Shr6EXUHa2zX5c5XjZi6
Wz8VXNA2Ku5p404Ep0VkoQih2esXRIC8SbOshetO5ajA3W3Oyngfm5r2lo0+mSb8
RrPrs+GUSVlAOmW5HKRSHJg+ZfRCIvFy1rbXdRUm2G/tj226t8y73xnhDsPx4Mpf
TRiU2b62HavZt+ceG+jpH+HIpxba60jA4K22SA1+i1PV/L8Ce9NafK1ztsA6xg3p
weCgrju0hPOA8fPGjepubYdLsO3IkDtCRRzlsFL8FZhhKZ669x6sIZdrDi3er/gz
yMVS3fMdFahWCusZblam4WxLl4Xw45KrEvE+Uxy/DXE4+eg3dPV+/7coN2+Rm8QY
nnE9eC8hdo1pNci5QPq41IcKZBSkw+6OeuvSLrTOVUr9rVFZsIu8DVwj7fObx2Wv
5erZMdsLwNQOJ95vUjArU6lBg4S/q2SsnKIxLk/ddVDfuDj8U5IgN1lQ9qgfMt/y
E73BLQYwv1gdpP98eWZMu6OXL7MTIqkC4kHihc29fIJrrkasq7hpie0MURYFYw8e
yXRpTPJdgz34qDsk22drUzVKwNtD6mOYmAizV4AU9N68djtZ7gLCJ5q/k8DMPlix
J48Sp/NK6y2eGT+Rn/Vb4futNb4DJh6wbAb3uxE+4t2rxsnoMzSu3CRc5PoGiQo4
PGkQgPErCd6Gu+22WBjV/xlSH+pppPwfO/5XNxzFwZoju81E7CbCJKsWywA2GwQV
eq5p9Cmbx1iwOuojCIDZIBpzh9j0aVvFfvs4nk0tM33ZAj50gGGtKUpkSLFqUbWw
djwF+TYR3CC699hrtN1m3ituelpFTaCgoSbWkcxNLEKdjy4hXNy+wsIex/0iuN1t
Md7VWKLdTUtfSsl37ivdoR5Xwu4Gs3+ArfFNMgekqDjmIbtyZ54iFilmLVXKIx28
QTVLefQo9+4aSVxWIM2tLZ4/W/NDXAZFvG48H0FjS1E7XwRBY/WLd4Moln9HaGaO
FREsbcdVYrltPNMz07LrQgekR8wR30bf8XY78pPNMmKE27Pj6tJ6gWuy+7YwIVSJ
ax/lYmAIgqAWdkbPtTuAci84ZZ5iJ1y4VnbODllbde+zvYRAIg85i77MPHRir8bl
2SFytOSZYqA6pAf9ad4TFQjxMZYsWIfyT9sfPngMOYDUlyyHWo4d9uaHTOMewVjG
hC7iympILp5g2IEqtpa4gFbpBrmmUQFMQkHWF0E40Ul2zlZFsFeRNOVXLcx3CFdm
KTASALPC3HfG0iqlalfa9JNj8QpL5xlXNPtJM6xBGu51r1mtTlOpuW9aC6fnaCCC
u8StjUh6zp8FU6anBP4SaS7vTzQlDfxumxk5IGhc6o8gyFm9YoMyq+4gODiE+WEy
UGAHbn8N/TQ4WnzF6L5PPMfjnG/iUaLpfwRlPtgs3JpLKf1I6fhVaxdVjukp+EFB
HM9AbZjXIu8SqlyFUk6BCSoJy1dTQH/ZI+6C0J7ngxzCLdPe0R+TpHtmOBTogxDk
gk0EbM0iYvh4RCmeouzv57/8bOVOHz3MjqqX6a2ThUp3eYKBZPgm36zKllGrO41z
2YoE0ygrHRURPna38t3NlJY5X8QaVI8Z9sInndV1FobMntKtuOhps7Ezlj3Rvw1e
Wd3jK94MPQhLAZVahX8W3S2RH01rqSEgLQu23MLDmJaTeI1Rxf354eYnQ7R1KJw1
F9xLebioJlTFXQoETlicssSSOg1PYzBz63YjPhsdSQi5vWx6aT8UT0aFnm8eiY+n
mt0VhZtU/S8UJrBUpbVwEdMbOwxOOU75FwgnmpkE+PaXtMfGwkCc9S4u1oLapM4N
of3gO0wXytdKwzpQo1oKibtWSGNW9MFygS0CEWpkSjg0kGxm0cTZY4+Kkbae2zb7
nVtgjY704TxPbOESWxizAJ8GtfJWGAYj7AnYR8Lj1mLwQ6jN3S86jDUZJSzVFoGg
o6ntYdYlnln51iRE/X1i93M6cLNuJxl2eXSFdVzNO6Id9rBxBVWe35t7bKiLsPjy
K1UtWd3A7boyDW8sjfWkYIgUCkcl7AJafpWM/yhtNE3mHmEtH/xP2GOLne+r6Ylr
jU2eaLA0897+BhZ2hJnd55+HoiUDoGQ6L+GGxFJhhYhxnjeCXHG6LY/qwRRXnCNp
kptcc6OkPX9N6qY5AMAK3T6zmt0g9inz8B9FqenTbgINIjjMyOjmqX8hQmDzeNvg
jMEf8wQ91DCBXaIpdsmYHcoIXhLGgV8tzsEH+PZtacW+qXKDJv/3/sgLVmvxGPPX
TrGwcChX2ston0kW3P7luW0pKWusP57n5xb6ydAqvrrdcLdkpXADSngrj1QZ5Hq1
B7l1QxyDQzeKk7JiP7FkJpcQw8RbK78hFFz8GHqISQEsHLlZw1BLVManjAtVogrn
UavYgkGX8Ek+GB8epk+tV3CtSJH/aUnTroiFzdAA9VbnHln2fBuMdyxokF3OcrMj
dohLoZRtUxMIrzsmIvpVYDAFX3m3r9z3WXmBWRkW9qsh/78Zjf4RgUXl9n8t62ET
5z/5eJP2nZrScwAOxt0QbLf69azczf8ro8YeVHkzpONC9jDjrPcn/t2ZM6ZGuVl9
WXXLMDLGX2vnxmGQpAzLBPWC1S0a/rChVRGTLmgE8Zi9FXVkw9NcdWMus8foAyAR
ar4pzDvLKomURFZHfslosAR7hIHDY6apz+Fjy2OTg22WdlnMvGi+mFjo2Y+b5/D2
EDf/9itz5A4koGJvSxY/JdD8jN63g0qu4imVil/u5ZeK4/0pFEWJeztGZ58WWC+5
h204VxuajR7XR3otMvmNysvsVFzVHec1X/0Xz6575L74mZR46ZUl/1i0sDLdQc05
pdfUltShy+nPf+EKo2yFx5FZzordMUgDXOKBkzl3Ihv/7nH/sIVaf8enS1uRZjze
04Plh6Rzjht6iqaJMoTfl+05gI5Q59kMePNLGtcnEqebop+3tOBO8BLWUSEgGeMX
kAFY1BAFfktMNAhYOxgBvau8/nIxRtJ1bx6XYnEyZDZjbYDSVz6vi7GxkAZL+dQx
rE8961lZHfreIzQZ6E9N2PTNpJi5HDKHvhz1fsMRDRUfKru65wGhLHtWXLln/FcL
sHVtzgoyiUaWHqs6311PKpuTdb8EgUAVIstiC04+15dQoI7TlSRDffTgru5BB9SJ
Hzc9p7tc60/Yihe79tqDocxLew11/tO8gmGM+BIPAj/N0Ck6ppO66UnOj3IT5xSL
8Hj9jM+sQkJn72ch5q2G5oCMrh5aVCh+GBKvNtJgB2GMGUyecABIQ7UKJyHoJVNZ
SLKDLth2OJo1WnLBHgoHMKELPOSsq1VQwn/sY3gUQzOBp/P+nJoXEUCbPtNKfi+p
sqglanzTs0qYkxWtoFcLVivKlSnz6ORVIYgS9KP+rXF8VVbNQFBTnHwCVhC/krXI
QFiu6JrBzPxNkVbaUYZdjmm9DVEDpTHCr3QRmrVyG/BpRjVA0/oso7ltPdPRKOaJ
VByxplBipHHHRnSfVjne8apaDu3wYoV96RQPxrrlprPhmqY2WDz83r46OHFWi4nN
BlCR5Xn+o/KsctzVosMAmM/P328wNp21JUZP4e0WYvJwhEc9h+eQLyJPeBex5bBT
Dm34cw57yEiYgkqPqhqVwhabYf02EG+neV/FsEW0YBmtrhN5B+4ta4tmPJS155FU
JwKA3E9lHGMzefM4ut2BE4Vyv/JwSEssYuvvk3eA9F1RoYPXyNqLIwLB0VS9TibZ
HDoVr7VPxJM+JHVEPWIcK9pA/io/H/nAsaYFu+19nenqIILcBdbYGC5a4RJGmCN6
KGtE+HKDDiTfgEUMbvPJR0Uz2H204SRf4q40WFM+ndF0jFQWZM3Lh8EeOr1Fw5Xq
KnzfWQnlhKHXya5f3yXFZ9oB9QH8Fv1HmPSb0LrNpl/129qClH7CEGjJLGU2tnOV
0a0DpCorbe01G3Q72tzlONbNqFpybyaNBmvM4+yqnKpuFXIyvgF4X6RUX6wP6R8C
TTst2Qd7OChdmgNT4yVzCXD6ZqTk4SaOpJmwFsJoaFncFy8PxISytigNyxD4eDW+
Rz7yi4rF/P05cj5BXSWoPHQMnRg9JO+4T5LsNaMBE7XzTD39TcyutYSiav9MJ51J
6Se90U011diXaQQYLbi89BDAejjiDVWK37cNE8UVvJECcfS/e+MHHK4442zrxBP8
J5id43eaVjBAX+QFNnI7mwdlnyh1rzsu9iktF1bv2BQnRxuh77QYkM8X8cU14yuK
Nv6Y9B1IRpGPNSQn+6lqo1r4hYtapR44WVpei7yd4PpD/rirRHzp3VDY6J8Qk0Se
QCDyUFvyxdpkwip3R9cFAXEIF41e6NiCFtCXbELkTOE/Ze5U9kQ15Nf8kTPYm0kf
9nWBWVlilEIpFtCTIp8zjPig+Ehr9WxgnIYVkTjQcxS/ZNxJWMRzn06zHJvMjLx+
rCJcj367K2GO2pbJ/tb/n9DBbVZm4M4udwJSnu2o/T++ATEDzkcwArsz0Fuxx+p9
kCZvRKA0vACdILzGBND20Da+G0UWrQP1uNf2mnNej5G3frGoC5nYndNva3dwGevN
ZLC0M1f9o8Yq8M6xXPMKWUAHdsONUlnRG9IgLArKdM2r0SOp6NVcP5F9b9Q1/huO
pVzW3LtgpNOGyVU7Rg2sRSuRolmBTdZuUNn6xYoDfcXAB0AvVgFWLfgRXs8V0XHO
s/78wTGWPhQE3hDwewtrwMPo+KAmLHtYJy7w/Vc46FxogSE+bUPn/2f0RroqBCzx
bH58MfJi8wOhoMlAx0WZo1cR1rbSzDifUsnOiANiyPOYGpY3z0Ae8fOkAZQA3w3K
jGHuPOMFsUMvsTE4Jl99Ah/o8msf5UImx/DrjpFx2HK/xMxHpuwV3X1/fy6hYjTQ
vz8RTMiaEnyd0eLJTRHtvNgFjjyqKhp0604qRrf3Hh7fSbnw1YI2TNZMa8NRYeLO
9X4erzUycoqCc03Pn+OHiLDT9EWJ3JZxZKWbNyVDm/b/j3K/56I/gYrVVDUpRb/2
eJLw06PMS/4kxKQWmF5B064MyrBr05uV0FrcWx/jgtrmUpedF/eSk4l6/gj7OZBA
qtXYGk+b0k/UXIaL4pFgj8huYpqfQ8I0PcTU37irM7rxko2wvTbvHFLi5hIR8dFw
afXJyb+XwnRLvqSxdrPk86/AxtQ8rOE/eMRwVTzpHIIy2GiFX4WiyVuN0U9kYZHO
sb5fvb6gLes8bCLR6PI8z/mR4h+gR7vrGrwP1JJg2OXc8Px8UX9JXeALGH6w+6S4
YQ9BJsVXqL4/z6fgNfrSptX3L3h15/6RBCe5G14MET/aAgX+wTUt8mwpYj8prS7K
EKstICCTfEX7CCBGqoWKAJ3/8BChsAIS5y32YYYLCgvzTftNEkyBXUDJ//+boJLW
Zagt6Ur1RzNOaGG59rLMYj/yVPQUnbss9wc9ixRQl5faXWPSMUUBZdimOOFr4p72
ejWPaFL9nnzDx0ae3I6OATBAfR5CfU1PjccYMXJvPOr1cFXKywQuj4OwOKBWA16H
UQBBJjSRY3JapMINqObe2W8aeXJYnipnfZtqYS43iNlGFMXcykZ53gYKlE65H3G1
AVCzbNmZ4DHNZf5ackbEYyMxRxzQz7uSND+QXG4zqf5bLuc906c4a3XA43H+RHGG
u//KomECKCM77J3Qweu/Mfpzbbcmmw49pPT01+m4KxceKuDNn/XV/Q7WWKPpb0lE
xrs+OFn41/SiNP0HcK+TKniWfTDdrxBo8WVxhU4vgsd/KuhXId9K8gFV3tu5IIDR
0h6b4eKoXyDdjvXwoZa580yVNKg7EAm1JDkfi+U3rxpwBx0+mnbH678d6M+JnAI3
/o/FyRzNUVUEc9DD4uoKyilznnPcYyT/qkLhi8y+0FV2ypzfmHLwO4heAAGDfiW3
jdN57lhO5XNLEMWm8JaZd1L3D4/GLWF2aeF3YHbsLkaa5EHGuBFq2XHKeftOcuVJ
nYQO5dcTUfx3ymx5apjDSVkuoguoeV2X6fUTKP4uVNKk4RK12gOLjRIV+tZzODv0
3PNCPAFaFb6jKj8Sr13il+20b0MdPDf5tPrnNZn2ijjkxVuLpIV40hvXoJ6nNKWb
WgVnvGra/dkUzuszOzF0axf2HDeyHZjpNd9CIamKsr2EQHHfAfPnRkuemlPCd9pc
KOAHqg+PW+oi4BM+IEf/x7OeV16WiANqiqBgICwNAl54qsvVCxdItCoksj+OZiTe
rlFz2VL9Ap3BDQXjBgfNoSTn9Tl/bP7ylqxAR/IgiSFrXz+1x+NCnjciSSEiZhho
i2T8/nbn3+MN9BoVUKoPTbWH5itmogKUopoAfRqlUZsP/viWBhCor9QpEVgtBqUb
yq8IoSSPhszH0sXiCy5KYZPCL4i4QjW76mkZudEwzTl538SDtPL2kiP29yoTVId5
tbVEVSGkaKq4Hnnng0r5ylV58YjfsWkd/7k9T50Kb+iGZWn6Q+6wG1Gb4SNWWMCs
9QtFjPwTW6WKRXP/EbxhwBnYw8TBMqbdYboTKrcwDijcf0qXIbfNeiCNPpQJ9dLA
xQL3kiH0Rlf7gU8YOqmer2oetmhFmbvQmcaondxzbJPd1ixOC2FgZsxKGOdet03H
XffgElP+gudZwH33IxPbjnbpU3e7Q84dpHXK0jdhsXiTBUpJ0nq5xKdN1CWsWHCo
LWNnj5pxMm6/rnEN/VfXL2hO5XzEcdPaRymWIjX77CvrWDcvasWI2F8oilCrNS3e
b/nnCEnhb5zpUC3BngpmLoDh0t64O0OpEmnWwyH3etBq0kP24a7m5i8l0IPPQnsx
xbZJ3zUoVWYxaNyRqVVtfeSaWXLNtgd6oXlTpCuGMWG6fc2C819s8b3E7zBbWUWo
AqEPF9IBc0acdFmXGdDipf03LD1f21V+YHFOJ83yt/S+V0nHaSQkSEDYrHlZI71u
ix07OpTrOvnsCwjXVLAAWMfW53ew2wXljG8rzgeazOjm6jd4jbLLOTbt/3qpcYwE
qzan6X3gss62WjZXWtEeSjUy6UdJ+2ZtwaykGC91D0Is4ktE88IVBPmKjES+ELYm
yunXRcETn3XwVZ1b+4ieZzBr5Se75xfUE0Dav+5Uo0TRyVlFKBT69WHpgwBgJZB0
zbyriuWn56WrAo6A5jNxyWoBcBhC12lkylnS+1YdXNT1kuM992UYUgQdpKHL2YU6
OAVH5Zo+Tl9PFbHVN3C8x843UPYgys9maK//IFI9k76QgZRkxNCpPaA9GhxvjuF9
MPWWL1+a1uxOhaE2qR+4J+zIBx4cRTWaDMpoRBRpl84BHSGCoJbmlzpJI/YQyX7u
nW1Fc3NnyX83ap82EOkcdk9k2Hr20tOno/HobUyWj/Yyn6Of/eg+0vhb4OHIrFJj
mckRGmb76wweCy9ed02+9Er9gUWgYmY4h+YvkrP7mTlOwFc0v9q++FUJ6CHpCPKq
+3WOB3MqmSigk9Bkxc5ebjj+7sBSolqkPCV9kczRtpLnPGj0mGmlPPNaNaB4bRTm
O0azvacGjLEdbZM91k3UFIH27hw9kTyS5I8QtFRSE+8JbWl3Qbp52hSEobom+rNF
I5wrNQh4PNNkT9BRhS7jgpRS9MuUgnEUNdjVL74vcZRLj/ug9ON4SzTiTDM4uL6O
vAxnSpbwcdXztUMmKx9iEVRYlol9BHJzwXVdQdDcs3w0o00W3uTCxlot2ARg9phD
fHeInLFqbzSaDadXNln+QYVoIlGbKo8IjNpF4ybikjlzdnPrMx6Me1ha9oeMvlga
lJcchb/G64jncfGqxORwU40d6Lp6WFOqpudoXkrvadjEJ8SiVCiYPzbSHS92TFZV
G3OdeOeinp7yGvautgBm9qtTb3l4h+nkQMXqmAVRtwlQdVbwNeIEBEPyYWmLO6j/
Iq3c+gsOcIoDpfBs16NvGTdi3BwgB/OK9FO2iZKqfHpFKdC2mUq19VD3cwaxh2iH
VKHioDosZyokHdmtwHXFjie8qORiiaH9AYvH0pCEvBCgatv8Z1yLKjKHdNhTszhb
Zj6gKVm5DTZR0q0NPSW4wZrHSxdw78up0v3MOQLuBIYs2T12hPVXF5nnhMh+eqYx
/JXjDqBOakk8cCLfd511tc6WYK4kFFWXlfpzuIiHwe7cuk9MX9MLzT60S8EIqXTb
fppZYSDdM+4g/C8zCfZsaVKYpqVqfo+g0p3ydrViWUeKPOMvsvhvYDGGl9n3bZcf
QG/N3h9NwVFnmHMEVrPVKJTuWQNO8Lsk6CuaO6orTwuhWyOjJqUaLo60KEs9ksJA
s/O5iXcUSP8BLIW258qRcfexbzCqPVxN2iwPxTKmw8m35KRF0H5JX0/4Y+vQBDps
lwKkzh7bTOOF/Ir/x3N7d8cQWrg1d3skLHJPcgbRsNMjfJVuyiyK8xAmU4F4SFoH
JGzwU7HcJL0d5MrgRLGrG9c2mRnBO5MDxOmRnOnICHC5FyRdPasyQeeN8lywByzq
oEzIq1czsPUrF2YqpCNpaImhZPAmWuS4UWdIu2Rh6yyFslJ6SovSue0kiw2fr0ay
n8YO0YSKv1SIphWAjMijw5lZ2CmRmJ81KwMNg+VOXsEKD0I0OGx6egP9Lz/OnXgB
9FsyWwpPfTCnvCdIexGCmkQSVkrUXYF0pCwQ+4XYHh9WEsDdhrJruoLmTuTDHVZX
SIV8Zx2/EXTUzGcTY4z93tukCphk09VaTkc+nH+sYZukdwDSqyoJkaW0wVGQqbX3
Grn1qfZ2/J7ZdiOp+pbd4pMOc23Gl22/aAX7bumH6huTgbTooohu0xQP+2e3FyHM
RRxL4ajTV0CPoL+AcdqIzMhz0NMWQl6DSMT9w2u4V9jTQsPa7giOT7UEPN4PU7Dj
R7UHu/d8F97xnlod0uuBa4m95nxNaq4d1kaPdMLuOw1O01u5BNDVST6f+l+RvS2w
MNPTziwHtvnl92VSKdQxWqqedc6YDuB14/IJApiOeid/PB+LW9sWkpSI2DpkxlXZ
CtR2qHvscaCeVqPJR3F+NcI2eZTFjjIoYE7gM4I5KNODOWtcjIsM1hF2ZKLckGwi
1kpI5YnTpOm6WENbUnhzU4ljvcrq/wztLjbMHs1kjvJ9QBIAQPhhumeJHI0hYxnf
VELFM1H2AE0x5ln2ayGhHt4+4Gkk/5reNOCDPOd5bsEq4pwB0QLZE1wFK3j5eCMH
cQDVkaeHF4wOPawEmosN8v+pFYenftYmVJuOkt48sNO6nUjhyC/Wynp/KGPXv7+N
fdUgJPrEhRDRvgm9/srUEPjiHbFA8d629s3sksM4KHyByVQJLmgpVASHlD0bcGIT
QFBBa1NOtWG/w12HfY4ttoY78jx8F2gXZmNVRRUP1QuXzdrxd6WGFq87GtFPTZOJ
dHzmCcJxupEIPvVZcj8LKf+lAG8LYMI0Cl/VgS62JLwaKgVra4QU03mDcmokHwcq
1dw9B4WUbW4EcmJaxvGgac03eTFgHyTqD0QW3TMHEJe01OrEQ7Rz9pm+1P+CLudm
lZzqYLnEvS6pODyv2/2lpTwojEllG5SPp6ds+ukqR7BE1ECvUWSIwAdF2FjxEM5I
NhZxo/FbFIjHprIXTzkIv3JrywnYDws/mHEwcDuYBmVxb8VUe3qf7m531W4t9pFE
oyFdiXWQyajFPuCHpYoQd0i84NzjPNfzwRQUQP3WDhYXqSwd5TUwRAvbpr2EAjmf
qGqzmse33KZ1tKlGx6B1OKCU9tatxeOhqJ181CORou0BhinCSxC4nimktCBHl2gr
uTYatcVH90g0pOy6Pb2jbFBdI8tHFOlFfFwcDAh2vUGqKS/lrWGGdvpV9HY5D263
/VhhXR1FV9AIa5jgX6jbzzyJ43F05RvE8HXBu8hkOGo9mQByJlSgdNfQtJIPd9lL
NQgxfHtQ6ZOjVrHRyvDBe56EDN99+vTuWMAKzXN2cz5BZfGvHlI2VgDJdO1yGgY/
2N40qGz6Wor6CVDMwPRWLCnCJONnA+m8x2EgbgDU+uCP+xSG0nzzCAJgUJZ5Up9d
Qd2JN1cPQwki0sc2b9V8FFkSW0vhfSRfSGcqC/RM97/RwQn9xiEdSJu+ITp0xZQX
aSAVsRSmkQpUSHGv3IbAgKIzbisabR8S9tMPy3Pgh1ULAK+1huEus+np2U3F2pcI
zRYyHA1MaR0i5IJZqRkYPzjHr6yeU3nFlnZgyHA2jR2imaLDS3sv8zM3YzBycrEq
ZBJ3nvS/eSwRTDQNquG8Z+Uafo1HCGNoVS8Gx1Y41H6rOl8TdGfOFSZvEW+Iy1S7
Dec6BgJxGKpw5xp1+wgk3vdXYOXR+lggIz92ACM/t9WKfmEunjbxNKbi5u013DdK
L4z0NVtesklLaADJaucVgiGCLv5O+YE+dCFrz9O3QwGGnGD5yAQN3y+jcwUisLpV
yWAZ9RPnt09R+PI2XUr+5yilgW9ngl0aEwriVpRXefK9pzOORQcrblrsKuj94X3y
lOukWyYurjW4KfHAd8Pe32raisxeL5i3jQeapx7ANw0zGZcBE/C3eLgm+7t4lAJG
MhdUUo/UF/gSCxfvzZphVjd6y86VhAi3dXOWaYqL0R057XyHDRn9yoczGMf2SgJw
UwkQZrvVukLmUqGA7opMot9i2mVJqHaZPnlM8mDu3WIzi/GbObRkOWVhRnlz0jpK
0ubUnlfOIlfeDs/1g9/I8qyZiyHJ8LmLX1u6AG2oqTeX8HQ0nWpTyqQulWP2dMGa
yEWynnKzsPQcWorzj//q2ZS6KJzksQ78puQyfqqgYtGe5U3/1kEGAoPukXaxB4Jd
xR52ogpAWKKmb0XI26jwo22qow4t25yz0ehN5xNzdoQVFL8JF75Rfim8dpogX05j
bHLNn2TzngQ+HF/lqBbReQRLZNwwJNhf6d2g8gpUcfZbNoOxOEkOcbbR5QZEvoUK
Ns2YedqRP1KhTRGeAZor7TFz/txRqPPotGvS4wNtsQdO526iHvjpBjx2kNovObOp
KdUxsQ6m+9gmNte4Mo6nx1z3TkaHwGH8XBYrkPDuyU0taAkTAFDeaMIFUSppmi8l
RYhRhEYF6cCwWsIYU2vOtX7PN2aaAOHYgArInQcZunAwpKTBezAu1oG5149eVw+F
HTe3I3+0AmUB5iOZvmczyRaM2cwHJOO/FZOi76Ee2pogGTKoNda4cS2CyjiwAvdO
VWqhOQLvgYzZk0o+Ctdju0fzlwaxDCTAUrzS8/s0RqEhZwUOj+roloCKhVj74l3S
IAlOyZcyHOAYogPvVBxZG289ZVvWZcANuPKv9FL4gmW8Uf8XUPB9xC6TY3eQrjFN
US4ngYXBEfJRlgi4LS8hlmDbx3WVNVebr4F3+04c+3rQ11wXplX7JzXQaG5Z4O2N
u9G7XDMRk856mYWQRIqzRRphwG2F2Z/Vb3X9Q41O32XUlkwtFz/hFmYI48UoiiqK
KeJemk0u3iEt4kcvpOaAdecnpIgDNtvDhpOilt4mbtFMV7XYnt9mg0L4UCTS6HCb
5rgGGLUOOX88anUnkFSg2wnEWnrP3oWpUpbJrHnme3i9KNWEwEbDtqeT7zzl8lpW
iDGiXNuNXfqATzKDM8oKGz9p3Fu2VQ5n5Pew7PBTqnjBqkuUD3aMYf2OVv7lPgrd
235K9EfmZYw55ajOLyNMDG/P84yrsoemzWmcK31sMVVSmWrc/pmkPlpWuCnjUtit
9msNMZiCci99cxVEJV+zU9xCdtFVJapALxjWJmk5FuH3m2jZyPM6B9yCN/fXoMZu
aTdW+PebyjOHsNU2X2/FFaeeaZfxZKM89N4vkEbDr699Mi1ihunZLXG5JDrLwSii
rI/6mD5TpdVbaDOisokPh+rcNbiXky92pBgW4wzagjPBQUNSrqFSCrqZ5QxL+Gxp
5MC2O0KWWKxCg1Wf7rLar8/oqwsyMsXZXm5h1G5FBIWigsVgStJC268gux8pp52/
8NfgPZnlsUVVTr0z7AHb5oCAQ0vkC1Fd8H9eX8saECJtt9ruiz5oObdURvwBETKA
7NfGcERYoqA2hc+tma8QdECKpxQ8pkentDdSJDjvAHXZj4SSOnTe6dxx8fq796tY
VLZbx5fd1zdP+5qLiLTsFrEV7AIIDDRqJFuCONPL0CLg9ySv1yOEWmqCuWO6iLQU
n6bhKOSHhkZOr4jKPAea0UFeZeRKbQQm37MYTnEnlCpXwqz5BNde3id+wy3eFGKX
T8ItRKghs2fg195uPtAh4eq4oJb4gJHSbsjIhV0iAF1l0DLD8DEFqymUiHvz+afi
z1cuN6P4ZyidroQHOP0Yi7U3gKDYRW86apKr3sJcuc8ZtYrWSj7roCMXVOHfYFkK
VS/KkgpwS8UfpDkVA939hEUvdcnQSyP6hbZht4m2YxcdbTC6xQHQ/euCiLzk0QP6
JSMWp6yQ9vxCPtKY/UPDHTVIDpryTHrJysnmH1wyUeIlW4tFxXxM2dbTdWF/kenh
bKy5JyJfke2BsATYDWzPSYe0CflbdnJV6OBuhxKmEmJRvaKVQRtmm1gpELtnorO/
DAySE6BCVHakFEopU/4vapPyD3Q2L9h2N19Fix7BbaseQGoQjCdjZCm5vfBy4Gsx
iLEv1n2f2CjnLnBZzPWCY4O/W21noUMlUA30/lVE57tYhNx/QUcIBO6tLSMsp0mN
8CoG8aGp0eplUUuqRgnZmuVBvRO+vzy6yn2oNtoxRIFWTgteULwZwE/Ro8XKADKp
jHXBKKlJ9jxsjRkzDRc9OKhUqcsVOM2YUyAIiVwpT+3cdGsSI2ITth9r2gLswM3j
Au/ZVkPbUEM2Od4+xblEdCZ6xDBd+B+lc8RIU/7wQkcA8ksaRX/Vx8GYNx6QTUK8
k2dZQEoI6/OU19on8xOK3M/TURWARhJlmq00xVY8F9Vc44h+WWqd8A9TXxZgL0OE
bciW6RfK2xmL49KsthUIaA8kPxdS41PYKjeJZ8XyL2Q3bUNa8ARO0czGw7Nyc6AX
xV/EfXl2U+x8vWE9C3mndMdnk3WAWiWrviFy9PMm3YdoG1ujukEJBqjsb+Yd6aTR
R81zdg97NIKnEkec6P+DyKpSOJkNthaey530jhQCfoSXzpEtQXlcYtu8PPx31O77
2LOdv4YFFhKT93zif2yuZqsvahJch5gTVWL0lhWUVhvvaKzkgAEBIb4VkPtyDaEA
3bvRuefUEQhwoyJiJ3JJlsaE+j4MsYcgNJD0WPOm/HNhY7yVZL1LOxic8vu5JUA4
wryD6z2u4l3PsKcOl8lKZo7FDkjOYk+prVVHH/2Pd1PsWC0neGPkvj2eAryP9Ata
7bK3RUpjNR8TL3LWnWQc867YQwmpYrPOFG1SqZT7vZBtzJcd/g/FCKHzMStRT3NR
od383lB1m6zzapRmgWu7KWpd7DfFB18G3KBSTEseLslJ4F1wX3aPke3Sv+LEPnl+
A7f/s6Eiq74YvvkFCkeu8In0C/luzElvs8URmBQILkQDu88dH6pKOQk2z8/aTQre
KsDTjq6KVyURGDSR+ffvGIq74QacmbSun3nPYF43Cx/u/XhdvVqJ3sx9CHWoezC6
P6fweLoEr0XqVLM9mI0x2C4ZYLFE6U84ALdMD+t/pmyoAfTtHx+pfzZAYZo+X048
fkqAvcOEtERbyixIX8YmechC2MBG/eBEq5OGI1L+14hndPh+c53cLBZFWTuD9pxw
AZsWw0NIgKZ9bxFhtms5Wnh5Vjzi77yTE5t9QIhmg939gmIB7Ap9qGy/xKVcxMHm
+8P27/BUl/QAIMNQxd3Ltpl7YTkkC2zqe23iD5kOesMoHTMzck2awTyNIw/i4RHG
Ir8LVPiCNnyQMRMhL7Q0UyvW+Vssu77yOoJ9TUMKDc3FYZHFb01+00VUEx11wII+
JJQyzPD8d8LIhXsYDb/ujopP7UpN9sb9mXjwrsyMdNeNj/19QN33ea/f6JPbTNgS
nNVUvq7v+ecco1bT6Phc5zLxStH6mCHGrj0vcQ9XUkT07uXosAYsbwxOEprUX6TB
95JmU3npx2JxPu5yUZPpCPFgICkngbex6WFrlL2EkX54c3d/X/JjArKjRPmdGEHJ
kPgh/UupgfUJoshkVAUM61Sxpa0Lr7EAHPgUar/ZmETLX6JdPTriwoLW/Or0LMPT
4b9WIpjAmCPVlxbAc7B7aFg8DjyTZQzFZnKek3uYGyLL361MriFwaXrfjEq6zW4n
NdU2ATwSkZMilTPyK5/YRnL0DyMboMbBlvwqvqyucAq9n25foqdmHY+Yb+lDIYoL
RI9atZ83UCKBafPOLMQSCdyCIxTjBRtiAdLjyomW6nZxauuFXTYXsUg8KxYOkqfH
hvwk3wQ32j8WkR9euK5+L8sj9W3xYzk5TCHzueNQheeeb/sFHe5H7/c6qB0MtySg
4kM1Nyz7ReoUpMG5ZRVOjyQITdnqd/LeRyMEdPawNiQISzYZsolsZev0faJ1CB8G
zQ6xQrPoAc/QX78gI+W9h681iDVeuyQFmX4iwgv4dj1DIgUGeLp9ssBn0mqhSLOp
w3NjdW+UFKH5ZdoN5/UvCmGuijCp1uYGGZjzWghXhxmmGqLq3HU3u67FcoY8jtZ5
QPIHjKFnIpId6dgfZq2BGQUSobI8vg1xTe59LQPB9x3/YgRsnOUWDG71TZnWe/ye
9WhTxwtcWl/iUD5++XGUJwPPxl392eqpGp5l7sYHwq6xvunZi7ar/IQhYqIK61fx
lFwzJN31SWK32+epTpEXYsVmDtj/HrRi1zeJXqYqgWH2fMU2gX8zBz2hc6NJg1LK
OJ2cdxeLB61SqcPPxojd8wCGyzafiPMBUXej4e9s2c1mTRoCM77QAh8EokhfUiUW
O0dvWSgHrkbrXYwQ+2FY40xnTzqCkWhcxSTRSFcQODySGmpOR0BKPzEQ1w5sX4aG
O/V13l0N9Jr8oPhEkgAUDw5p5PM7jsVc14cw1he+A+dW8PAyNErkkm+krXHMvD8z
dBwUWho39txTm2OtSZBxABWcYZlsIDy7oBZzTDmAeBf209Ltb8fsCfu69tNuqnZ3
udIkcGR7GaxNCQOytm6RATIuxVvPUnWZzjn5/1QEzAyd9M4UH3AECNuytqMCrMnt
cvf8fSJLsKJYU9j7KwFz2sq2EQRYwTvo2u+IDzBJcQgC3meHf/MORczMOAWYB9Vy
PUrVOXbB9j6cHaAifwAFBagkyTKWiiXTXtDmozTMuODcA7vicE+z7ughsFswEeDz
fQYbfxXLY41ZogmSkdtXbbKKuJ8ZkjIGtjpkZ1w2Wh8U8QfbSbvp9lkJ0/LVd6Vm
W/P3SBDAw0gKSfZwCEJo3zZgb4cw3PK3qkbDqwEkKpjW7lat7R5AX0Gcgcw7Qa/8
WTFG8yh3PbOm9mhCzspYCU1fP7D8iURnMIjpHrA1v1RXeJSD+p4tHUv1kI9xo6jj
LJkPRITRejy8NTj38jmjVKEHZ6mHqCeaLyecuNJO4K3BCg2lMZ1Cv8KTIIEn1bV8
Nd276Hl/HGkSZZly86PDLHlJnqApc0kfXPIA9IPs45auchXJf5ywP7jAj5AQaXXR
GPUIQClWg9TkX7SEN1z/yeL92txssXg/NP5QNLmRMOmckEyY0FvLXE6eyD/QEIzU
M9B3EtBjDTPjspE3yyALW02AsStgN0Fdkj8tezdhi4Ol2qGP/MkFwpKlzh93qOvP
IL5sRoqTr+bS/NoPI7bo730nX1NjEkutBaOweYUhTUE8TbtavVO+27Bhg/H31meJ
LvUpLEeeaKkftTb88bb/nfSd1Q7SIb1Thy7tQcmCiTtrVIgsv7zDv7HTZOdkFtTI
N7uQgxW2/6raXk5vjTPtzdNJNYjO4idRmeO3asiKnCrQaPGpSBjIuyClVFwfYUqe
a1zDnrKBB5ElKqNTnv+u/bNCWEwgN1wrzI4yDfa3n9IwcqeyPulPhUq9TGnT493H
6kPyKku+JGBDSvqRYHSRbXe/qYloKalDGb2BY0VzQPeRwCMJ+l+dODpBt5Ou2Gge
hpAPHArZVuT5uqlgvOfDhcx5aNPXpKUb0Y3bfPC5Ikdydw8ZodNn+srZ+jaCiK/s
Co9N5y1um8xq1UwLjiikT71aI417u2wNRjmO+XiTbnerlYV/3nJBHFoYQbED3pPy
yeFU0f1s+524xyRiBBWp5hduvNEL90Zpo9eVQ44qwJ0A0jB20sJ5/SBuUn1gkSHw
sIuV7QZcV0GmzIDSC5EhYpc4O8igkugGLeUc9ss9dDX7KnG2JxuHzpngi8AtjLWC
iRtBYN4nV5IS0Pdu6NC4ya3+Kk1VdAjv1epqOfmFK0NTiIrQNrMh0wAgT5f+JEOb
75DaR411JnvLwDHW9uPDrrwSTPxGMKem5DaAtWY0wUonzwP7LwAhB5Hqxg6bHrH0
KBYi96c08g1i00cp5kZurEXgt46bDIlE86T3SVgsJCbxBHgSZ7fzenwWMmX8VrST
vvbajTYxvMNTBoLMX61wpSarNj8oyAJwlD/WZHH2QJQ5DVVDcas+L+ysiewU63Sm
4m7bt2mMLTIhbT3qhT4NhhrZ0U/if8zQEJtylJxb2vxyg41G1Ad3RK0DPVDw1fWs
2yciceuvFJ4wIDbZiDziq2u8mWJ/iAI5bF5Fn/fXJ3A3aCr0cpiQgVfRK9xgAHln
EMgQDPY0rP2Gm9hI0F1Ol448zSuIpHvGwctvIgAh335Apo9StvIPt/sUkbI1Hk8X
i0KLVe9GonLQ/iwX8Ir7Noc1FhHdOCav7SminU9VdX1ok6GDeiwsTA/mSFjkFcPn
du9kZHH2HtqQCB/uNL5+Y9C7CY2nK942p84zdoV6jAP/dZcH4GaY+INh2bhOu0BY
xChrVHh4BM93JfsptCvOfW2SAG8jUrbNGUJKE/GcqOhDHsbOH7tszdsN9Flbfx4g
DEbFKJWkGmkxLpSWUIvr29QzWfp+sf9Pb13dXTRSFebpsRVVNaSACf0ME37h6Pwu
lGjKYZuQ8f9S0kbUMHZz5K/3E9tFfvs0eLl5yTbw/PXrO1uXKI5UcN3LpN4LMw9+
VTOhndmi3XTIWQbsUFXitqdxJon2PO8Bmsq5ei+60/A/4o0OTJPn/alZHxCjuMW0
/fEJOzYzD6IYqcRg2SMP76vFzzFZLCqsjIjj0N67oFuQ+7D0aGJ2FCfTtK9G/PCm
9RKBOVcHFc2TG6DDZ2PIhP+O8dgFJqqe0Lt9WcTfRnmyDpBBXnDoD4bA2RUg8+dr
+PKlrfWogUI70hxZEM5l/YnzHO+SrFKeN9G7LBSe5swsn5eUaG+/HS2/KylTK0kj
7Wzfi3Jw/gT4A8/FPw557K3IzI6eKoztR4CYygoEDc24ueDLONWGLp6EdSoLXfpc
pas80fTruQm7PzjFwuTGIbB+lN+ES49BDWYX8cbznMX5JkUkuuhQIcwtz6FtCzfV
pABIyJobpdq5ZrxALMk3p2Qh8ACwirXDc/kB+HEC3KMaUCCzZNS4vvLROE6p2+1W
ovrNa7qbCJE24JVnpvl5JdkaUkbNcv3B9v5E0iGXPMJ4zQC4GwNMsOFvwAmMgfdQ
s10AbInotsPrPFmlpMhxEPrXiHKObq4yQcO5tVTk+ParklFz3YC1nywFZQEhVstY
3wcHbPXuDiA5SyY2YcmmFQzPPVN5KPmP6Az2vrHTxO9lvfInlnXu4QYMzEych4Rd
CrQUCR0p8CEFRQ4Mdv9Dvl7HjT9iDBgFGveb4OX+fQYDXmtz0mYqK4cxfE/TpXbH
Wj4nTMCOEO+ZTFL8HoimHRZImig0QylcP6EG+42E7pkVbzpiyuMDHBGXaBcrw/l2
wQSSbyxuGQNDxedPUqCBQanBEH3JsVPlwSyOk/3NQm68bMfdR6rmZ00e7DszWaec
5ZwW9F3x1f9/4AXXGxqlM3pXWcZUuiXeSpfOpG4yytr0PjcM67gDCyBsX/YaBq8M
iOpsxfrL40jZRSh3e5ZwhMjM12sqBi6umqQshrymWtrRc/am+TmJjJh7qnVYjDtJ
YRCziiRiyaSzBBrK2TC7jjcwTYEVUYm31nFbLT66yB50b5IoCClY9S2vafocDD2V
xmpxIzaZfKGaPD1kJTWdubkFk6PJi0IdfuqgeWNDRiErGuRmND3xpOX8oUJrF6yF
JVd4JE+0sVhdh/gcZM0J3UXJYdqbrCjzYHEwDcNndY4vPBKS3/sYK61TbSIjDdQ4
aKROo3zH1qvQjvwYHYqNUtCa7JZZRCWXo8FNAJPcRoTdPyq775ORb3iYFoh5GxQI
rCtFrk9iLwxV586D4dkE0lEgWztBtw5xINaiO0kfH32wcZyU7lQx8VcUG//x2MNS
gToMvg3M228TIroufUQPQxVnBHpUD8qwRfaLKK6cRrOwjsWxh2sNDkjEaX0OOGuM
a5bImU2RSKIbNA/ZpHCw2jmZy+tGZN/GCU0fgLEF4DpluXp/AENJAvShtlwGj+3R
5n0QdBET5QJEL1cS7QQKe52Jd4YO2egYt8AzbgixnldBiGalnQkTaa3wsZK51gJ4
H9YiU5XTpcAA4FzTQ7aoR6/gUVwKu6cpKAjqVFTBGW/HWybFqORmeg+f9V8VXg5P
bfyZR/xfIBCwuWCk+qicXgMKZ5tyz0Tgruprl6DodO61+MDwpVzNzN+03d/fRm74
v6IrAR/igFBm0KSX8J39lokavp0FZiqvAfZlQ+oV4OzNy3rMt8ywykE4Vdt0HI/l
gKs1Q1MAtyh+3DRsQ8MHcXWB7R4Nqt2L0TY6bQ3FGUZ3EqDaG3xLgL1dCAinypxp
Fk7fFaD8b4mRSaj6pPAzvMuj94aGts1KxHtBggimj8w7jbVB84Ckq5S1VP+cTWjh
jnN6FLEu+RGjp17wMI2xV1v8Na/LBoaJBu9iOW89Cc5tYzyXpyIN41XGr+lvOj4x
tH9ny3aJld3HuH/GJqVqLxbBcTZ91RLh5mlmRAb5aEFiLeVNd0bm6HDXxMQzYFM9
8A2S1qhcAU7vLFwkz8GoK1Q0zH+AzgnZK15TCqs2V5jwAp3PuxJNquGdR4qlVbVR
vz7ktF6LxH0Rv7Sy2xx9f2iymWgFs3S6njd9eOPziDd+y95wddBkXL0R7S5CWdhd
O3O+0B1hqLqCDFs72bLmfHBeByf9m87AtkNc3fh6jO1WAliafUgoaOy19lIpJqHU
tM0pvLS988Dmn+U/w8QlQoo2RbGkQxGtIaXWcCPU7JMTezLLE1HSnUp3pk0P/jrd
TOToeylwvBLFQCD+seZ9VNLLA7xxFNRDSrQaWCzwb6pj9hWUPPakopiUIygsTYjf
IsS3N+QA/2zb6nho64ktTywXyMdqQZ0yMCiJLOdaeY0QWnXvbLJNPZq4eZz4KTeq
mSxEH7ajM0iWZjNgU07LPWXMfvlRI8wwxJ2XJUtSFqWfl4SMZgBspwrpphCkGge0
Gi8Ps3ZBZGIjSVSQMUjMu68c47rJRWQX5lHLHdvssclil2VrGQZHBC2f/TWUAYrD
deF5gWN5zzyGBNvR6baIfwb7oJnNJ4d0+SfI5iJLaNnvr7sOf8EWCEMQlb6xylbO
adfvak2UxRw6XUOOShOciShZJRSKm04RWJ4+pkBoElfeR1z1XQ+Zds5UOVkKJ2rG
MdnSsLi3zQss6qGRfrmYHv4UMqnY+btQBgU4exMEo2YSisE8GAf7j7gGS/C1V8Ia
KvKn/JKHkc1CgPLxkPjd2sxneQ6Q+P78Yj/pXnCy4P5YJJZ+AvVOzvseHMApkMcW
+hkZ19yFLtnMH3ezshgSljymdBguhnuzrsg5iM1QiR4FWTVhKGnmOJeNBjWZodpu
Mj4RGBjar7Y82tkl7nt7yZLCbfBmeWYiHsbp4gCSNoaLodO9CEQsf9BIGSwTX0NS
jXQ6Vhaj02gTjXuxKIUB9PV41Yv1JRZ1Wz5/7x/w2nVbWZIdZvdBpaPhM3Xo6VOK
AemDicZ714xOTDBeGoPYhMdtQgpQD4rc+R1jpdGAqiuE4829CNPDRdweoFwsYLn4
1zMnlTm8B7WaOyqo6ZWmAfnduxNuVKI9pz0rcDhWpbOGljRPFWl8rlyriPJGQmSA
SaK3aPKy23Up/zXd/S7cTiV3wdhuqV+0OY13uAv2RdcIgjohcTLjgboIdb3WMq/Z
hS9AEWPiy0qcMvPzPKMUAee5I15W4Z0otzFE7kelGKXUV1idTBRDXTPLNQZxs4Nm
z8WjK5xSCPYWaLltiC/JQzsCukKyr3+nfa1XMx7KgDVg9U49cK/Zkx9j9UhrHFPV
+Z2mz7Y+ts8ZKySZoPYO2hjXmVQeJQeBoSVCjjyRhIddDWsMK7sQ1kacO0fLuNEB
ENyz7eieeUSuHWH5vU2pS8AgnVP6nvVp2ab2qpTSGnEEvNoD+iq3cYeUeNOcr7+q
YbGxppI2sMHQJMzXXwOOOC2VhqGzdSJNR+BXhpBk6Twx+7be5M4opNg1DvlSkfk4
wMZxdsLVf2IYkLY19/bs+IChqoV9AsfunD8sWgqpzLr4r3WptybRJ/6/yjLA+WAs
8kulN7yxSmA522iX9WUgjc6mQZ/19rqkTk0dlCEvfprT4ZhrTcm3Sdfp1gcT9nAy
rF5SS2ubif5q2IeVpB9lbW7d1KaBmQb5NciBYJ9tDiayIfA74MOxifoG5BaeZ5nn
fDev/Q9uBh2YlKUnJmSt2sjgoSGFJcxkljPu9IPtx3xXu3QqPdpt1aZYPhjRJlhe
jL7W57nP6E+noXpKFYy9UJpXz6GSMX8d6NR47lAmdmWaLfcY48W+dGVfzciDGGyS
XGPNmls0G45/wOiJiX7sfyqoPFzM/fx6BpatQYSzYmmm7ifWUEiQF6pdwy3wT0Ka
uampQb308QsMYUMXimX32D9qeJWIdDg/FE/3INOe+kWvR5WLTKMN8eRrosb1117Y
W1eb7vd/iCxJYBIrfeCsOKAZI1OLWQE103Uc7x5DZRCirw9uOIUhO9RygsaTkESJ
hRyq/Ll84BOmECznYyRK/KjQyzPBb2n0unnDXFUzZ/bztOiK9npJWLEwRo2++o88
PdVj//jYUFsTHepa6smHlD7tfW+m9ue/4WKENJlm6IBOZUNxXST0U2zxXu5S4EXJ
jn59KU+HrYp/vO0abAfJaFgQUO2RLsd4LtcCbtfFe+d2RyYaZz3Fd/99ffWLwbKa
E5y9FfgVmu1CtLRsbsf7XMi7HazwOQw8VnhgtgobkQluUyaxFThKjZJoyst3M0Zm
X+ce/DrOmXHRGJte+rckOR32ZyD9CihgojUBfIHfMbcuv5qJfSQKkQpUlL8jZEzA
wiAdUNPH0bY2S31sIwh+sUQ9F/DYNbZs2/gNEc+m7MHHGS5IgDns+X9c0ZAFDfzy
REO+1C8Hze+MT+pCajHRvUn2PtxG0QcJhOFedyfVUWLx4dyzDuq3AB0pBSReyt5/
8f8mLQJNPG1qc+0upYZd03bqGy/VDuAQ9FBXBM6JEjbOZsjI7iLMXo4dDCmRyVrO
huH6pK3Pcq/tl9r9rn0ZJtcS7ihDL2S3KCDdnmUkIIY+R0SX5skeji+OLW1Iu/7T
NQ3iBJkY5V9P59XAOwLSVCg92i4BNBJUf5op7x1192WHsxigGsnGXSVSSbXIjEC4
hK1QCIzi+yiI+aDVs4se0uvALkbDGeUZky2KTo9S1TURfEMtiX3Hyf5IMukSKumc
RDEk7cGSkFeExFwDbJmc2ywVSvHhjF4wpNf4EkAgzuk68ftdq3kGiM43ynF/vXuP
vCfvD2tm7yAJSl4GdB4+KndSL7U+sBryUDjGI/96d+W80OsT34v+gWiBADIDE/I/
c3/6RyVFO313OlRIZIwwOYiqSLxSHb621V3HVXD/fBB7aeRJNYLmA6Dyg4rYJwVq
N91atAD+p2DGyt/rnNAAjJafMOlM07zXZHQUVIspouBZMAe/VMjjErDJSXXSbMfi
601e4KDWp81VtzWEHAJtqr/RgiIZ/AANbL4G+xoitAqB8BgNjrnOOt6vJvEkkAgW
6WtAmYPPOJKahgVAj7qnbvm3FysWfRb/BNlMIqD05KO6+lcHfW1Px2OiAKUJ7Qm5
p0iJL7F++qQy9OCBzdz7riQ0vjyTYp5ZTBwPjhUNqpW3RKQouxMbO4L400jqUtNw
CMqIFOY1QSvkOr/4nU6ODO2/UdX8tHcnc4fzUooGvU7j5J0rrWb52PUxg8hW9Bkg
42vuB7HL8wbsVhGmP09qAfEJ1wqHlGRPiQkEQjePD9JRiK3x9so35o8dswAsFs1L
UVxO7vUfQVb07FxyUftAHdC6gf/Z1NIJKF2RzdmawlT7u5kk7gzybM1fOt060Bp8
8QiCDaOlS/JsiY3uGmkL2JRARexWtvfAqov4UE9c5RMFyn3cx6QeAJN/MDqxvi6e
QiIz7/2/ieMfbFJs/ZujaTkCSfi8M6AI3DfODZPQsoFPuO2PhESYhKBaEHKlD2nj
hvz+88HdIs6FFgwuHTu3XKRpZCr9c81UY1RdROsAhuYfX07gQShQt+Y2FBi3GTkp
P1iDtZ/x5i99qU4/iUxMZ8pXPl8JkaOQINrpiFTBEzGrgRTqBZggnoOwJ6Um07uZ
fIOTTlTXV1Rp+LDajewAY1H4hM8gGU8So5lcmNrFwSOa6x//Tsi+8nhvKD4SVMR4
UlpKDmSKZJE5/vXWgeAVEOmgVMzzt5Aj7XerWOuPbbRxCwBZe7NmEAY4nxWdzBAj
R66nMcZplX9SO8U4Lhio6xL4pWPVGYIMYKOpMGEZB4vkIehxRlyqm3LscJ2lPBL+
3hAWE+DNCBM9tKEOJso6V7uVb5F/jV+yfhBLozj46nnEzzkAyvFm9a8l/6wuKYqz
HGqJ8a0OkXuy1tOm9/6e6ILuKSsACqcDj0mtPysBDPx75W5VNBIIVVA6F3+4V6wT
eTOrru67pgEFVaSg5QijabYPmhA7jH1Xrr4CAAIhO8nzl9l9injZynDCkOKiczcc
hUvbcDxkDQzdpTeykiOiOvvCIGTlnJX5tm/8k2QWNi2kVgRFpzXkU0ZaX5nkQvbx
y4AS31S0TYceg/qZatCw0A4MOUIllJCVH0gXObQLZ9FAK2LZ8mpDW0jJdOBVUzSn
DO5Mc+D4tThVrqHEAkBka/Jekf+VVmG/AxZkv2fVDbYQl+O4W22eXMOBAPWXE0ht
F9+7r0MSybQs91zmz7C1XaJDkVOjdJJ30xVJHZzmlhfTkZcE6ymXW1Y2ccVuqe6k
OWGgRbd7eSb8kahyrovN03YR8gxSV8Dy99vtOHGxaHRAG/HEXWvJAI+hQ9WGmsCM
tCyXIXG5wLZQX16xFHt4Tc6iCGfBFBAv1Gr0IcuvhfLl2wGN1AbpwIcxBqnsoqpC
eEN+14Qb3y/9Z6RfkzmJKDKXJzlzKnBlx4WTVln4K/WuamWHHA6Y2tGHv9Ewvanc
FAE24UGr47GlxVcpkPDK2SPDQu5+vPyXlKpnK4x+GcycS6FzSgfSgujPGZzGVgok
EeKxaDaqrt3UurAaujdCtDGCmxIzsoFSUFIZUI+Jm00eSL0P7x01Z7c9pK3fryte
BH8XMlK8ItTPiCEGABlYb7p46d1f1YjYiOosssYqM51ASqioTCjy/Fu/MBduUxYv
zdUKQPwWICBicLvR8tqrt/Ch0x42ZbM0nOh8jkRnrQrOZOuZgyFcG8/XlU954pEc
tzoEkMQ7c//G4L7kLx/KYbpdadfhI2eXrBhkXJ1rRasanUnjjQzzaP+8TXoE+wPo
dbUdrf/lHFnr4zci737V0eLVbQRDniWBkGbDnCciK0gyVLGkQe5cqBGOSn/kjMqI
8uyUFg79UueIhSgr+0A+K7MI973218ZA8i1ehlwauppg5U0ku4jIbVRUE0ijl8oW
MF5c45bGVJBAvTS2JJcLiHIkyELqKBM/tqJ8dINELSyXNjZ/JnL6UeqmSjuPJDFH
2pPdBGyk0xt1tgfgzvro/vRxc0vg9FDbvcHk2oIHYkU7g1ASF8SC9sRe82akaM/Y
TDZe8c2gqsptFk/hRly8g8HHR2EPE49cfF/Gf+lyRGJiqGNMsOmiUWz6Yk0730Bu
fAOssfixmlwxE8j62oePokAdxalB0N2KAQBk4pLcHyqlYtVzJvUlEyJz/xi7w9Z8
dW/29NUr3icORh1ka1NxFB05CFyzNJ0DvdCsE/ZLEJePsWsjG6d3EqLKl9E1c9YI
1dQ++Z/mzAMJhXyNUikjq+QTl1ye8domKPKCrAukg0bei4ARxW1xJgH+WV9LyUrd
Jxef6bUZqmmda2ix/Q9Ev7CPBj4/NWLTCOteSCf3adshkfEBXh7liijUtaC11Y2x
Iw/Gl4348tfnHJ0vyWMokdgxAYivTP2dEZPmsNYQEzfiEbnDiugwEwxFESOuW2SW
clA1YXQvgv5m4SSwDsLmmErn/L5p60rQcqS/9iB09BzsR3GYGpPzsar2ozpVuehd
1X8Ky0M2ylbeQjXu2stMTadgGRVOh4e1HTjkD/hYWyx4YdY0E8GXQjjN7GVMlHI9
uweNq/VQZcBtIHPwuofoCvtpKmnkb8XqDkcZWO9stLHAwtgx84yXxpSnE18UOWe4
DC7/7iPM8vyj/+/+sJx05tHW7Pefo9quse2se/WqLPEZtrHC34lRDbH8JBYveFTg
GC4+mvAIaXTbBJk1MnwdHI+tjFTSXQKReSLoti+zKlT3I0q1tPjWsdoIBxeNFRvI
MqMZk2XfXkaJgjoj9DKXb4kToEn3WqYlHEMoF4IqqIEnE0973w1AqtU2dzeeaBFi
C9mhhI9Vlsg7Wc9tDJV+Amj+40tCsaeX1k2Tn2ORS/fAiVmZI0MBso7kot5t0lPA
GLTMlvSwlcJo4Q0H8+A5+hx7yTaEHRfMum87Cn7ODJCHOHfdGc5N+yJz/9FUbhA4
td6WgnODE1/LPYdN4mAbv0CRF8+kkBZ8XRyThrZ+0pIqyv0EO95mgInKdfEZah/v
mZy7KjMgmr2rUaqDGpFoAcAId0Xijw8xcMtYb6J6KKPp+Zxk81ETop7sEV2z+r8H
1PleQdCoJM8+R+Jt6wO9CquFrhzkbVH6LXp8AigGepjv1B/Yh/PKv+T9klPQFm4y
8/sHpTy5uBl5BJl5nw1//Yv5vztrI43d8r9lB1cB0pqU7C1AyuLSGAOghPA97cZ7
8DeyQhjs4N+n69TVa2+1av9hPDdEIlAXXdfDOY2ZmMK8mjk4YkrvTkLhf9XiZY5X
vZ6tApMyVeQZw3ZVsr/+lk9YqLU1Ryek4kEGa2vd5dsEEXnLMMn4B/jYFZhNqf8i
QSCk0uWqgX89dxDbXZWeugvVRBxsl7fD9ZlfVMcbjS/6GnmHp4MKzi7ikQ23yfZ9
4aaQBcHWWEnYFWizdx0zxG7dJ+XDwEpdxic3JvM7XI+K0sEs01KGJmWrJCD4pQjC
i7WXhkVHnVIV+Y6GIohVQW7iWpN/gap0m0bTg/8994F3u9oxltK6txytmUyw7vbJ
yzLPGWldQFlPnoLlqb9GYtzW6/lhVLLE7QDeoKuG/TJE+pPi5lDIReAlgQUMplpG
QaSuaRlXSVnNOqpBg82R7brXQ1Jr9rAT8mckG0Ain7/kXLNE4kACLD+8tJt8SMz+
IqVV/KrHxlRPVjutOSLox4SehgBre78X2iiL+K9q2OuNPKO+n9LZ0TDMN6XiSoiN
TUHYMH3sbCJg8NCHeqIrLVmnUXp9iUJW/8Yt+i4SlVkdoaPBcFNojL1sS5nu7g0t
t1n+jOzCkg1Z5ICDkAg+dTMsIqnWp8cE/g75D65+B4CyjoA1mN4JDBH2u9jMKbjC
39NAFSznu43US3dfRFIho0ojoDt0oZw5R8BKhITX1sGZXt72qr/Q/9nQPXN5RE8R
6ufnbaw6lHAtG3VCVbftfunKVUJa8blNMYxTGkvw5P5zIUP/cCvfWHgjOvRUEXnM
FmyXp14o8wClXEjVzBUknQ0IGsW5Cu0SwxgzTp3W/2yONFHMQRlKG10fY2qsR8ak
l5tkCk8agJAKqUivA4CuxI4i+uVIUQ28E+a7nHXQ4wWSiV6zugJwiQC+SXaQUFwF
njs9nu/C60xULXDNqix118lUh42iXbDskElwAVA1csFBx+vM30EDID5C1aRaDCK6
MqOaAyrxjZfYkU335RXUYBV4L4XkAqw1OpfV02jdIEup7NinLd8kyfVdt6kWM+mb
YxJ9NL9qZ5QHU776pn73oD4mUknyl/wveslEK7+7itzfclVyiEtony8K1huh6nHP
zb01Yp1AE//2UlQ82SoayH++I2BOcEuxZnPk1MKapQoYHS2N0NpNKJAXrT1thLoZ
qLTCVftrzaUUy9xI0O6xtqKkaXCmkC72yFb/AnoqXeCTYcbirW3chvsK83pLw9O9
9E+3GmV6QIbFS/EckDkVD3vvGgdAj/NnSSRCSZXMh0obyRaCPPF1veQb5LUJ9td7
uV/V4LN2Cj9kHAjb6lvdx6mIHNytyLS0YuEywewHPE39ZjFqMLQVtpeP1cZGBTOg
4tamytXiHg6vgKXtjQJez+nVTw9r5Fcns1NpEoyFghntezRmS/mQH9MFsDm+e8CV
oq7fBCQzqWsGi1FBkZ0GDry3r2TjCMgBVGmoujmKOEKuVEpsED3p7pMu6nHOnwRH
N4X/SM2mcsK9w3oVqP7C+JFm4ty3eC2WMZ0/RVJgVBMDVggKeWYTTkp6AsR271jT
Fw3EMsPXjVtO48zRB7EkfW9LlIomrTgm2CKxcqCp0w5w8IZ7awmPnemDzlDwigIu
bZfz2O1mTGh7Qe1zbOgdiF1GQC7gf5bTbK0d6+x7W6QdLYag6BhOowP/1p8kq6pn
oeWEWwy8FI1kVvaEwhqG616jSB8yBpASAp/Z2Sp+wH7exXe4vDcE0zb5JqKLf3jt
pGWOxYR8/1Dz9HCjj27SA6avduc8qP0DWGlCZrKdTuvJacCbDjCc3hUkkda8+uah
8KxPLDogtUXJ8JFl0INitkYxolpVdnJR9CX+cAy4rLkxNaAc/OBw5GIKnJE/F2dE
ipHucQB2nko9WsLpNBNP65/Ps3Foo7EBgwg7mwKVTLJiO0zI6PsTWSOrOK5EXF2+
8+PXxEldLrvPl5VvrM5cW9ES8lBFIzqxPN2vAUpZ/N07TSN9OMiec5bqYB3LVi8o
qY4GKOZtqGhivP52Kk9tiMVI2EgxHxnCNFFj2uV8+sBUHAmLCv0/KFNfekIH7gBP
ZXqW4cqgVCvHB1XHwPFc7NpKS3mKKg2ZLZacurTbczb8Awf8lyMpKGsHhAUlNEcd
a7leaZOlf3RFScr1qhZCn++oYKoVCrEMx7GA/naXdVf4dfmql89GmbUwtNXrsjQu
KDCOycl1VvS7TymY6C5bJh2P7Xv/gATh4RemYVQ6jGJXlh0UadCEXO6M9jFLP2mJ
hIcdAO3n1ZoLemAWCORiShScYv5kTr8WwXnanFC9Xc/Smg8rrQ3aOMsn2qUYKKKc
1/Tq5JrIwOc1tgfMtYYZPXmICYNCI9xbinaP/qH1HS37C5O2kzpELispXmzxBQ/F
wmyka9apqR7ez5L6H7UAEz/GLXwyx0mNrZA/rCZSqmtYWgm0PCHON5v14htg/qN8
3RU014VowOhPn7cYTTMQJN8tx8+rua9Kh5k0iaAQ3uhO1JXAhcfcc74Dnc/5gCSG
+fJyXWXxD6hGeqL+23PHfchnN1vxDezwcXY7rxKrmI5arxsBqazmgW6/0v63///B
+gL2ho+/WhWrcXP/khu1WdJ+vXbMlKgYoIrQM63RzKVgG6QwryoD/lXQrzGWkPQO
o32ZMVMtTXZU8dXTGr6UvDEfTGetRTwl70GPJGdF17gZvdW8rJPHtLlcEYC0ounk
4QqRL3v2r4SIdZ06/iRPKKnIMAWmg2Tmz/yAb18BprGmtSuzF4TTyA6P2njI2/i4
bG3xJ/xJt4chhCPd6dFdu7fmNmeql2cxd/e5utjq9AKDpFgLl1xi0l5iGM+gm8Qx
M42CjOQmSgJMo1M7IfDSX4wADKixHXsw6fmppE0JNvn9EDJxjzms2/ldM4xaMgd0
VUTLUAcD4OXSj1ikzbI4a8uWyUK4JXyO0hJnU/9ee6NX+LaxKn3s/L+1iLwTpM/W
v1Jo6HuiCxbaf0F3uKJIbQc9NWEPo3iiVIITkISNz/896eqbSKuAZ2RUo3eT+NKR
FLskuGRvlXMKRJKsKc8uY9XQuO5qr/rC2JR2olidhdZiwg9hyuacKoMS9bIqy/jG
IeYDZNPubEbfBcUi/idC1DckCw+XRCW67IxvKJ/rQgHYwn097fkV/Wvq+mDTsB22
FaOgu9uGZy/JRaBE7Xu9ooNGLCNuR5O1V9lCs7XB/SdxA9M1JEoQPcGmppvE4ZF3
P1o0auBXGgSbLojJjaJmiLT82yEQseOiCsslONfgx8epqMC1NeQyyMz1kveV6FJz
3bjLVthYWjCMoj6GwHXO8U+alNHk6Go7b1AdOO8E77lSxisJ50jY8DwydOoiKZFw
wfbJZTPE0hsr6zzLTUER9rF5Aux7KLsOGfiKOKrQ0Hq7QFymyoqH8kMRWBIPHi25
c+8pgPO/D8MRuP/Y48E+t74U/Yq2TGyEfRk37/Mzc8ejTf3Pprj/ignKBQl2D7Y0
LvQt53HNcBwExK0sbzZxiiGijt8rwsqfDs6BZE7XW4XH9VafOXdgLLymgtxINGfb
9RR2uiD/N+XshFdU67Gb9NhETr5A6YL24MPTsU/Iv/gEpONfEtdQ25MUNoOWlR9j
c7oc+Jt6/kXugIfp5fbEjO/LD3m3vZR5k36BGFEcu/58CiGIr+3gwXclPN07jdKR
ZclC4uHBAUDgQYbuUstJL9UdkRhEFEbTNhk34oGIHEjywWJNC2bD7W+SAsdNsUUb
noZ0sw6AUeLe+iMrRL6MxwPwhhtde+qjUXR4+M8uLPmnxVtDnFomnAPpTsF7k80q
7wlcYLv4izxHXJRvj/1fePiE4XNujxxvicTmDtVVRVP2t/TjAbLN7B1XvATcdx1N
a00yGcLf9qSS+lwBJBBUh4h4sQPGWHMP+Rz6oQQjY1qc/frjBGGof9re47iVQaQp
UHXfhMmOMbW38ec6pNFenunFXXY7JKTT7hNneft+SgvH3NlxTodapQK4GXZtp5DL
DLNdxRzjbldimZtbUYhAy/DWEeDnZII13OWRUU8cfr90EZlxaPJd/J3XZI7HO3dj
aTnETyteorw0Hr0vuP1B0krOYq30o6kHJEYS7ISoHR/x/Kx6gtdTSxwVqy+qwRXB
/x3egu+Yty8LqYIzC79lqjmzwzC13C4fQ6zSuxMCHvvK2C6l/FDc1UrI3jwOXzaV
bRd3wanAnzyPdt9rGWT9Eh27p91Bth8R22IKwMm99Pv9ykEkBRVMw01TuHBAZoup
V3WFimhmAcu6ItLZRD+khJqRLG9NL4jQJe4oYeH91wBTgrKAY/8PTQvoQcszM9mG
EFB04GHiWRlFBEKlX306+JOE6m5l54ADc46eLE16dS+AiYeIQsyvcvkkDmzmcq39
sh7hOnM9mnxPqw+6RsDuPy0VuwJEnby04TdHeZLdz7jWSKUrtX+XssmDSacfVJzb
GRBxsc4t3YCND0rVL3d5roFHdunpbS/7RaHjhpkUCgfE8O+/qyiergc6untK17Jh
dN51GJvejGcOKLMD/01Q8NTs+Bf50HhRk3Wq7BH40Aei/9Dx/Wp6p3RAfrV4AFj9
47YU9oE3QRvHaLbN2AGTWp9yq+SifssYQWjVJJ5bEZlpNim7j7ATDJirgUBTHTl4
fvVpOuTEjOSrgNM00WSpGv9lA0Go2rKTOJLrBR8TEWiolM15vFdhDSOzFQE1HS6r
eR4zuCpF5bUhNSE/F7fdnjywMr+SJFNCJUbDxO0ZIXRkq90CX+3F9xLCKKhnHkFn
tpTbK3HThE0yXQpi8K3MZ6AyG9JfeB+gAEmSKsm79y8dtHAVN7FHlsMyATlnu7jM
VnG+FvsPoEoJaZsfQGWDiwmrUYj+3C8s1CC2KoEoYDsG1jGCBj0ZPas1SdJFFaUJ
qk5jxOodpCJ+r2ctqiywln4s12Kd8S3L4zPWw3S8SCIEphRu4ATpSI+O98Q31tpU
fA4lK09RX7NlHktAb2XGpOwrFZZiHW/Q89RJRB8nWj05xFwr6QqCrlrsp0+tOhQB
aCdWgBejWoCFP8Gc2PqNzbtfS1AIrt52OcS1z8he6MLJCp3lO23IVNQiyOyA/iD2
piGSDGTYbIaTt8NzWuFDkPd2zPA8MHzFhET4KSFNVIONiqHfshEqfGvQKqG5pZm9
H2s+JX5sPL7u90RaInR0iZU2xpAsUraXbhOE6G8vheX5VzbaIj18SWL8ahv2Vg3n
V2OPyGRkmk8mXkRjJVlduiFK8hVrfKQobjROkWHYNsLN1SyYR67ZIDc3r7mH63MW
0Q7WynUlcdHoQaRWjifEB5kOA+A21PseyxVhnfjLItX2FgTmUmFP0WYBwM359t54
5j1A40paL6+BruU3Em+2vMnx7Ze/Ag8C5neVcgXJohrO11I/LhIU91mVZYlBmESR
WbC1CqpxuwE4AQpRZy9MJoYqoD/5YQ5cFrFmtqZ1+KN84WeDpQ2I0RNdGyhHulk6
PqqmjwV6+otyQkSyIk+gOKN5/qteEgj+91GzHdFKe0cH/uIhZQWIIH3SkEI77O6J
rfYKEtEupVA4bBxyMTnZRc9+TDJ9oXY2sUkV3KvUWC6U/lt3nP30eQMSSZ82MBF0
4heTUsX03rrCUCv+7QnX+yliaRGXG9LrVTdFtdHcE6Q72ikYlbzh+UQKEHXvHna3
sKfliQtanNTA+mjvIZ0stGJknh1TR2Waz77nN2nYEXGGFZvIjjcFHhruu+4XYIBj
sh3oM4VgwPnTwVk9TJT0Hi0M7XzA3OgfSOGtW8R52YBo+KG0VzW7t2oDhtrjB4r7
ocqplyhqru27bIC7XgyDBHVXMJZUDPJ5SvJQFHbyBz/CoubgU2cTecl1umZtSkrl
12VzlsC7hgMWpX/cndQRljPZ+sSUxtFS4wIj/P0Lpct33BL3ZbpkVWE6MSjQJpn5
3Af5185FFAsIr/hOJQFPXOg/WTDH/JdPPVtVyWVn/2PFveMyOiLhm94RaBbDLQA7
iqoJf5N7s7BIiTTz3C03vTzIxE8M+6Ei73p7RGPBOTojdmdIbfnJZMaGa9CvMhiQ
cdNQXD6C1EPcb5AnmcefU5DASQYyvnA5PryId267sLwh+E2X+zCeDeLzoTYaqcYM
QgjYFrKbUIOGXOfmYLhfj/jO4WV8u56+lycTR9wgEWD+kZ9EmsBYjC6VL/10JGQl
lgHGQlOSu5JsgBk7RiMGZ7i4LazyT8QOVGuz6udRCdZ+rUZoN8UNI90NFZxeZzZq
52UfWO8qGYUwjDqMCU0fbhY3F9RZ6e4Yb7gjGOMU2sLvqRMX2Gdk9G2Ea3hGqoHv
88Ttqa0gUb1aFBOhE/atB/1VWMv4WoLyLVSOQPEUcbym9h/DgXlrQGt7tZWTNwWc
U40nAUBYhe7rjLELjA5Y3FrwRf4ltnp3LZGYvwi+6M/ZlBeYck307QafoPRuTF1z
KSMOW6WJ69J825ytvofDsx4YObHzBydgWJg1yjNEnIleH+5vV/4N3ltUfI0Rst2e
GOPfrB5QOd+Y35IgNQCxVwgfKnnrNNNzPOFMNql7lA6uNA05FksQGOoH2eqtFm7f
bwHOh05YIPX7jjNEdcwAhlDGD4u76m8X0mhSnTF/Dji9lu5iw617ghzmT94o8/aj
mKj6srHHP+dDAf6bfBKTTeWcoF1467krAAQcBJa5VVg5XiWBCYp9fxPoJKprexjc
HbtF6FKiTbLfAX8iccg/LoeskG/QbUyYfmWXVXCVzMXKXVUqLZiSM3MzlUcK+MCO
Ln6XoeItJBfvLOPkI21fQ6sg5TDRYqu+xFettmPZ4KfqNPS43n6B5BQhGhZVfNEd
AdHF19gzMvqBTbICxQcSKWCf9W3y9n22U4CpmNQRdw2dy/SZvK69cfRVg0BKByOQ
2qByPvBGQR+5c43NFkvtztdbfhaUFjPOyDbRa5wP06KjT9NAGAMbVj15N4HR4VP0
M440lUHcah1jeDi1V6HgBJtkGy6mIhAYYzDh79XRWunCoSwiZRtl4rOVQd2b2JZ8
6jwsYkM4bL8V1CHKbUwVLTH9jEBrDAFSST1kK29x4EkhqmoLZfN4xW7wa1CSXGsy
sSD3yu+hg6x0JR3sdEXs5RFq0nslgHFSSerKGQqnMbDuyZC9tBFrenshgBcrHC5z
IpMsVMqcCNDh+pmGPLO6rwqMTNYbKceAiXvZeQFPcljwIkjX/IRPMKs4jYJDy+tw
0s1jSXhX0THESwG7GJ3xGngNIZivb6VNJ7os9DBZJiWQ9kih67CgOSm+INe2UVZc
1W3dsUUgj+M06qDud22B19f2owVa0RXjScRszQxhQLFJ6FhCvaN5hGdK3Pv81eKd
C2D7wRYdDQdO4ConR+HjZywZkz0YTX1ucXRWBbc0kHG4P32FXStsl/jIRsP8GytX
iyDElefJxNprIglaFgfmInpqQ7WIFgfHpapjqqC3z5myVDCk5NEmSUL07nhJk/wQ
z875R1OCVepjm8OISvYhUOwtvYii41GYG8YdkiwQVSbsMUBiyBgl/Sjmf59dds6Y
gj91OxEvlufPgD+9jd66VtFjsVQt1BkVKqdAfnsuVXue7+UgdZIHX3Yyvi4KYkdN
XwsIeXS/XMz/jIvQwQIv8IQSv7YP2HijtXdDHfoG7QJ5YYnEZhzy3iraUlKAng9e
Yf4fJ5hicRDOEi07BGCjk1JS8MX6XVXnKG1988QS777UtrxDeBuAFYXLGlAUYNtq
bBFD0xFh3Vl1ejmkuAiHxJPTf7X2T9l41nZyzDTfgzZajJCvHhn5BOlbJTfMgd66
i9MpPw/sAkQ7O2nwWGFbwtKK/HBHBzIhOeywyxlbkXmlLNUsU7wr4LKuz0UssbUr
o4bYLY6EEIs1NBXA8M15vMFt9mwA4MK2zseuyCyAoB5EPRnWWIkH/jtP2LQH4hhw
B9JQF1l3li1FJ6olGDCRBKZZBB8Y6t48XfSpcsmUffmuq+5VwVCUa/1YAf451ibN
EHZDPbztzXxXyv1vu9xOr1Lc5KoUPl6IkdMCEGvauVXD2Yg82wU5CSqP7IPjvBNy
+W+CtzGh25ItjRh/qP+qifak+/lQAk6DpSLCmq7kuPaH1uMa4eVYB9Th4rQP40wA
/0UJBWaqk/xYARzdLT05SM0Y6vYx1VHPb6n0RdmRPbLzvjqh2RCUNrKnefqSYzC1
3MIWRtE67/+Y8ALUT58N5/mlDDN8LGg8XndkXd6BHKKSUghdhXkLM2Jde7Hb5V4k
nH44y9ZhfcVJOQnPHNQYx44Zo6kB0+6O3lcxcNJs7N2eBwgSi4MsqcNxOgEyLnTi
v6KA81E2b2yL5yvzDSXeB7UPTs+79Z4M+D9JkONikPyRxyj6kKB4kFB7/lp4yxjr
19xWFl1uQbFYu53IoWzHbvIbmr+XY0Gb0gfzDnw3SQupnUFTDBZitq7dhAh5IykI
YfDBnUcWlajY7dJ7nfY8euCeJeeCaltoc+tl3Y+x18olj24jll2nGPwD5yJI+SVL
nufwKSQA2a2xnxywXx8bVeUBhWLx+/yucckbyA8RgLJI1ih9fcjKtvqDvgELNsbw
xX0aS5z10M5M4s8/PKy7mNDjOvE4K7AIF8MRqX7yiFRaqA6G9gzuEbQq+on+J1mL
B1VP2er/gYGjxH4e2QByXvgA8myZ6D0XIxQIR1rIRNBUB00dhETHMwtecGF5cgBN
onDutcQ3UWVVl5wMX2D6sYbU1+RkOCU/fh8sm8POvQLRb8PwTXyB7vSwsrfMh4s/
nL0aKVfCNgMz4dzWE9Xe+lsAyBlwrqnYpj5+SRu1WSfReqJUldKoQMbI+YSn/NiD
48XoQC9GSTNdM0qOng7WNgImfnhDGuhcPYUKUw5jGeByAPX7hHQWnaG2wv1cZVVp
asOs2bmQ8wB7XuWXdk8tw+aS5K+V1FzPbbbCNRlC/d07Q2vtD48QpUoXqwznJErL
xmcdYI4KBG6HlyLpP7XN3glGdzEkzlHY6+9x5BaUW1lA9wLQ4EXXfWp+Ua9JqrNj
ydTLZ5hzm1vNf58efyxzCvSrbFMdlIHgUikOEm5kZNEKT5zO2rKAzKRkunGFfdpy
Gr3a//b5wT2fNFa3rPKMQGvc8pNOEhCVOMENMsZ/dRonCBB84SA4vM+YRvIkIiec
PfgA3EDYW2YS9GTlk/ObFC3jHOP/Xa9Essjpmk3aYzbT0SMUeXnER5YfeMYK+v0O
0YT56iPqo8o3cox+wM+COJ374EAF8abVR8mhHSJy55L3tPTx4U6DKv0EClgyUtVk
FB6YvsuXB9PM+L0/cLjhCDYtAKW+xk899pVl5BVPGxxWaPn8PisUSMkbTeI3omor
ufTJAnOhc2XdKnLQVOh3+MIOwGOuAI7nPppni1XSIE7QPSaX7fR3FTJVxxEJOvMX
dKcn9S/zpOHDSeb5ko84EZ2xd8L0k5WX5XFIm72icOm/NAYQN/HDpf+TnCQV4awy
rM1aRW4SPu75BY/fji06u/DEuHG8ct8uB2vUgAma0eHebIDe8YxuxVc7AbEfdQ7S
qLS4Qid+BDzSuhyFAg1rJ3NU7x8LYbz67H3IPGzZ8Eu9/bhn7ntsjEx3o1Hq7CGn
JtCiCSQqkahSejw9ODIDOajDgfWhZ31HCf7ttVffimQrF7PVLLj9bZdu1/hJ8j3W
VuxF37/bQLBEwNKMEg7Io9n7OBMyZh4yXMmyj97oWRw7rMyEDJ8dAkg+JUmHydkZ
6/fY2CIL6C8vj4zd3r2RQjLw5MMo2B9Oyfczs9tuDiTvkEXyzA1JmDZfmU70X3o5
LBMVFRiayLIqLvz57ntcwe46ZqyROccE4zVjvbN9Ng2m7NIuRffVNIjSQLqY4Rzp
HvlHFwqEcoi8WXRUr5UPDwnq1sOkbBD4ghyNRIQA3oQiLldTGJLalFr9IkfNlKns
DxuPU9XFZ7yiGV0zEd2lrdTW8steIAWO8zUQ5ZEBZ+ipwgGb4pH1ll+9B5OxaHHl
6Lsu0fL/olN66FdrqVBd6PqEEC5AT9caR8khDMG1GOvCTmWANBhwb1MME3i8vI2G
kusZwgm7dnsgcuCWlJIw+TndKxPkI1coVSK4LFN7fI9veq3MizLeKCRpZBF6To3+
X+lpl/M8fEDy9Akw7NGXlw3pssGwJMBjexAgkpwmtCC4L1lnKtXxuFQIJpY9AIzz
a2hxR8a0DpNTvwtgxk42a8CcGU6yhv958es4f5l9Gl2ivNp6X1gZaGMLs0ADuBmM
m2PtbX+SOCdNfEsrNs6uZlgxwE6biAchX13PxwiIrpV15JRy54IvqLVJ+Gw049l4
g1HInXB1/ytpWub6a49WiQo+504O0Ky1pDI6I75ggxexwj52L8p3VhzD9/pWftHE
SAx2a5ygqKiaiiKsrHhFBUfVHbiBcGexz6lCZ/tLNrOdeRBgraKHjoN9GV8dODi3
ph63Inu1hZJhyfCYlWOyec42ETTXkMK964xUnBXUkcC7dVGKlElFdCDyV70o9GRi
l37wV/bO4PFsKXM8d0uKnWbd97DjIGbhzOg4g9dEwQl9HRwMms/O4XUYdjnp6lVR
9WEkNOkIqU4JyqVorfDcNrj54GbdrxhYp8XVWw+d1tAwIFpPVQq8Z003ivKUDCPk
28rY9AmDpIKjreupcomIVwyt5AbGUWHo+uMvBX2UMwRsMdl4snhm6Gg1xDB2UEWn
zRLJejqWfWQnk6ok5YO1VyMS3NvIxPsv1oEt5zcvvnjvr7JWq/yvRvzVpJDRkoJ6
5UNO6vOZhK8AbHe1QwNxZi57aaiMd3C6mSVmb/wxWpjttedCbPJmFdjzlWQzmzL8
7V1nYflZ4UIy/kQZllEwrHANxzey1uJAaebZutb7Gow5bQKvppGbf7Owd4P99HeA
c/Ecfepqwb7eH826N+t+YBrTaMtHxG+pGSbpB3G78ur8Yc2Os+Zww3fG3h0FxHaW
aGJkCXWIjtQtzpMojxmfP3ogMXaLweYeMrn5rkxNlwZx3qw0zjK5mKlRlHN57Z49
AgKYyPr3bLEKolTwaO9wjGA6qZfHAk1Be92ov00SDLJqwxhS13PdJwRS36Gs6DVX
WWXaxmxfszuHxrl9oUzf1XgbiF8Nneg5GcjQCLg+yaXGhsS+77xQmYrtjU0IiptI
7q3PPMmBdvBtzW1XIZTy4d0VCv+1+lqhcERUcD+aYv0vSR0CDEg2B+Qtgalpx6QV
pFPlHTSzmzlYssJYTWqXEmLxtmLuzZgXZaYh5+XTXeKdvnvynqNWCtvNSVkbTm4B
iRLRRczIRLParrYxmfRyU3tfY9dAHnLPAzFPL852twA3a1jgu9IWXyUsfjY8H7bD
KO5vKjc6Kzf/o1qAnkrVTnMYdtPBwQRKWvfGQHWIfnIqqOSm4xcuMqKOiGha5R1R
KNvowDbi/YiNr9i3yzK5mTQyxvNT+IVg+30QwdlJ6e4sL1nfKfMb/titCO6Q3o9l
PvRod9PU4XpTdIMX5irrO13DozsJkfdMTvURtPMWtvRvIMa0p7i9W68MfictHx9j
CrdyajQPtCAX9JB0bhIL1pFPblPTTECjFm266HHbd3vKwVa38VZfxSnF5W6xDG99
utYBaGeBvGcW/17idKYaZksCd5hDFHDJcFe9r6aZkTBOmOPffjUIpL6oxqf+OpXi
5MPuUvR87+ku7nE+CBp9mAODQYluxIYB9o3CXHYschgIDHnns9oM+QbKjHbnG5o0
R6fIzsMYoz6uyCJ0mxNZwDYt57qpoa/G+F+EelG6Fa9PYMOu7bOndQQx0v9Syidl
35KarwLeT3dQ2Fh3GqVg5Eo7By/ZX9hQ/+qIuLZmoKm8sGE6yw0XP4uvjLbOoGZs
zr45gj2klvwFXy873uLPgAmBdi/h4YZsOTPnOjK6X++n2LYx9L+78jLBFHopcjet
J46YxHErk50HEPeh1yWwrvqa/vrpSFbzeHaaCcWpn68LZuum24AEEGRlhnTj2App
8BKz1wOHg0iHDFa9pMqiYjluTmlTHF3OweoS1atpVR1sq2vzTbJU47dN2doIx080
pYIt/NR66l6wB3O4AdQ8hAmirZX44Gy6u0xXCL7PS21p/dD0WUKi5ZpadGcDcAMP
NPH9tQ4iVAXztD3MeigmRAhBhjYjxcDc8hnAsuQsoVx6avWgzMbDFf/k5RM7YvRS
qlTmB72AG39aGTHLv5K5fUBKKm4kW+W1dBDUSf3jMeHjnmpMh/rsHssSf/UL7APZ
I6YAzsS5tTnRGE+zhk4nByx2NtVKeluy7s2/Ko+yDPf8dkvkYcgZaIVw/xEZjSUw
B/VM15hgRN+tR6QlASka2jezL0bTehHMjd4eJFggMVMwHO60VIzgW/6Pv+nfTLaV
FX65owvf/+u9tQ18mNlwI7FjVVpQaSn7MO5A89J5EE3zYCp94Iq1nc+mZkzrLTPW
djr43dDzPmcc4YHH+E5P3cWwHlVWtbGKyw8PivCpKqW9e+dPrhYVl/9+ooWiOuFF
/U8E8ft1VhCuzDIbkEo0Wt9F6MmaCJo4hcR58S/cS089l3McTbox8y8eRC+GKhXK
80ImoB03Wpxx7JlnDWhor30V80VjqHzXv07/+thK2IA7X5b6eFGDHI1mUJahWf0i
vBuJrX6iMGv04xwY9ZVwh3TNoLhxr6ly/yY4iAMziUPgHiMQG7DW4cvRE7tKcupL
DHV6fQYwoExR7LtFwVUb/LFQ0eeUfoZHTRC9gOB+NQD03lnEWPJfbXm/IM2kIUI3
lMk86e/Ixspgk6k6AlMDjpIPfmHqEgGy2yB0Bp94tR7jChOWvCm7V9/CAkpNX1Dy
IvG7Fu6yH80Sexy1ZxMzQpSkgVr2OWwSvKARaba9WrwIuPLklZ7jMci9vB0ZLL/j
tGsG5oZaX1Yw2XMyrsVVLE6Aa6mByyZGFUMtQeiL+M2+UPW1dcUX8v5kb46B62C7
gfYAMttk5fYA+gpbZD3ugQ5QY5dfM+G249C6kxLEPbQ1DncRx7XXdqlIaALN9XmS
rdTcsCEk1X2OVj0+Is5McNm9mjBa96JWXSNmZf9s3iLeaXt5D0CMqGhKfy+XpxWL
gLU+W7mVfhrDi0NIYNwF02D9O9HKloJwGF0kY+u/o8OUf2GkHfUR9opYlF2+lDvt
ifNvRXt1Lsezj1JXu+EJFGb30mhYE9NlAh11CgoPS4tLXi1/iGUJvF2YlNczgu9B
rAqZkVPjg+4/AeCGxMJvwpES/fhA3kMm4Pfj7x3ATQ4GW8vic+17eUx6XuE5h928
S3TxhWHQx3t/Yf5mQqSR59taDamssdI/CaROG/m5Geart3VSWOnRv4X8zzEnPTw7
X4ijmmdjZaYQpT3uWmOjWZ8E23D9rOqzlQedLnuAk99vQG2oTKZNv9MuMOl8sbN/
xHKwNCfp5KDr0udGQK/sXKFYfE4RLWY24dbXSWBkhxYEwP6cWepCeu2+K6I1uACh
zcQscSFltixiWzg5nk+JELfwUlgtWbZD841aNg8aK3a1NXgT2JdgNHAg/AMswMm+
HerWvJ6kFiye5eP3Y5bRoCoVqsgTd5uS4Lf4WM8PD8jyrXCDs07iEf9cbE0T/sWk
zbiWJivUTH+F28zr6VqfqlZJts0Gl0YOO4PqswBXrSRD57IkFDxe1dwyeHAFk3Od
jbfs5FaajUh5oLZl/bL5MxEAxPmtIZRbZSrlKdHq96H9LZ3gOBAONhlcaf1xc+zI
fyWGjK+gKdQOpHxek/HSweP25Rdx67xhgGgewy1hc5MFDr+URtnzXNLmGx3H09PI
8AsjMtMVZg1RNnxNDnbpJoLTW7eBILyj8SFYON+KQ03J+bYOkNm0Br8K2FyQKO4F
8RFM4kvnrke/HJTMQawBHBJv0Q8+FdFBfJtu7/+aqdKA2c1fBiQ9Ql2QMT68evUs
G2LomnEF4pZ5+JwoFLBkF7HsnYBw4KV42wBWBLvyRRGhtmNJUy9JY2DARMUxNUVQ
pcM/Ft0Yj4Yshe48NAH4vlr0LbA812P6uNI7uo38VlhfVMWmJ2iWz+LXVKyMrsJB
nBB799rlt3T24R08Ml9Ni9t1TfiadPeAHaCm1kedcTsddso5IMBk5Tt6mJTq9pjt
rliF+VZVjapWqtUr/2d27TSyDyqVhnl5XmeyrMsjNvSpLCCKwDe1jA0q1JIoD5q9
nepdZmMdESJflY/v+hKBN1jvs3G8m3zNiBUcTCPvrlCB2q/oj80XBEL1vhzynqqF
DzVGboZz3Eg4DK4bsWFIpxPZLp8fCRm7vCrjl3DlRKR3R8JGOSb7Mc33x3vdt3pL
Iz5wtoeTD5nQhFkaM/9Ci8gem4OYVmykRQR/fYHSKA8iVsS3J22St+O9czDDXHCy
pz7uCwvkmlv/s5pjhFybtjPdDXMkC2w17659kg+F6Xa+OyCMsjN2CQ6s5YME+fec
zmLpoElI4D1E3DcKqPRAW/8yxqEEu31Fmm4pbv9p4fF8F030d7ObSyiSQqSF0Yx+
3qpJfECw3YodfHm4SZSIdqmwgfG6pTZTpBOTs+XZKkb9shFC+LEG5JjgvQRivvgZ
YAfqEdSZ+rXn7CjdAEohaqQFEeeQ7x7DKOkBLH+Z83DJZssweYseiPU9MRF/V1TP
3bCtdjpbomqpP7IIPlgjrshwMve2V0/KaVLqtu9U/oUi5YCsiunP8LP5sNBq6UEh
+Q4RaFnStbIjnQ/An1BSlqGh3GtsWJUlrYF3wFc7T+LiJqMXT1+ppax4gSsN0Xsq
X2es7cNk8Cr88dWzKSzfATAehi53GISqyWRbzpfZ59Pl8RUjYtinLaMH/u2IzTNc
c4HRruSO2B9jeLe1MicD6oce7impHx9Y3SdiHc42khmN9rdLFHEh7SGHDxHM68Ak
W0FpV3IXCNzGvvHU74wg7EKUNwZYUpbCor0vKQnrGIypapl1wh9JXzZtDQnmb8Mg
5o0fCzU/nD/pKbf11mO9LA1Wstm2hz6naP3ZhtoJj26Qoh0XVjRZqLu3a+s/HU7w
Crd7QmV1TgGqjE+ZaNPJbVrFCNA5OD1A5rn6PKScKOUK1Pj9gImr21hqcZoJyG8V
FNqcvvaq+hpswDuos0ZWgI58GVYoc3UBlU3Gd2ddc5J+YGTHSRl91aOqk3FHOBTz
dlYm9uOiIGnqjqurdvGO3MogyWxepxEyBEQAge+doMTfavd1bD5pS2Wgd1tCNz1H
cZ0Ry95V+cNF0pvJGqeZ22EcJVRcfJ2NTJcMSU1a/NnxBXtMYcnnuMAU+2WM6qSZ
24K7nHwgDUPqiouzpitTiHoV+xMAVeK/OKaAtt2mqBFLvfhpDNofzs+yJql0gCEw
RGmcLNtb0UeJB6gRmmulBQaxOCtxfmTJXW1oURDfGy/hMGKBxXA1W0PJaLHq5df2
kcb4nwHVdwrjc9YnBPMjCc1PP1SG1g2/IACQ13uRd5ZakigK7EkDvNQA79NPMhoC
OmRYwAmCMfebpGYlxKul6oqbmdRbu4f5erqD6lsIQ2/DZDowaFJ8tij3XvLCwmlt
BZwiHlKnJJFlgtDhPPQfyuH/nZriZZ5PZ8PaqNlGILjmETucYvphtiM1ly+y2eIl
Q7HaE2P0Bl0qZtAJlLdONKSf4dt1yeDkhlQMpsAD2b6MssxfrHsI7yPIx5H8q705
AiJWXnS7TGdyKccmMLwOqd6MAvKzQB4RVhIfYMOLQohXWpQp1ddjZGEsx+FgQP/h
GRoB+ol0JGp4Bq4BTlDk0G5NtGQRVOPWe1ETo6XXXma9G+dRgxy9G+GUljQLVjsc
r9fg8AU/oU383elYHj1TNpm2oHR4vBjSII+rzdIWzvgUk/2vUxLJdc3Qty1PDVe+
KYTHaswO2xv+hw11s4muN2C7qF1NrJbUcMYob/xMOLNj6Yoe6ZKa2Z6epFCu8tod
2kCd2xwpW9m5j+yUW6QPDvHxXkSxzLXWjk8uClzwndiO31/WU3W7KeRU6wEmWwHR
ZiGyQs68h0C/sb4k8RKBPtzb91vn/Vn7+XSS0Z1lsDPKT9ii+5mRAN+MNwfD9pEy
gihNVJ5aPydoHk9S29eO722JDLVexikeqDoV7nddlI7+VCGghtX9u144Z+1S04T9
JUVWusubl4EfMW0LWl1bPwfQ+liAUkBGE+kX4XEqlf2vFP+jROokKLvBBv8yYfc3
b2DxHmT31TVRC4sx7BXmFsDkVF8s4xcU6iqr3/mmKMR6A9sDaNWn/V7DS7bmBONp
QI4162nnp3ZKomefgIN1oJP+FdCGL/5x6d6WDe/Ee/ALfcD7BMP9laZAgwF4pX0O
Z1ltm+7/YBZ3fbwxEZ+6R5e3vk7/PyqK049tPTrtHh1B1eG6zvin1FYUIB9MVyWK
8NWq1wq7jHRavs3qMJmTGF+oKjugGG3tskKrupDI24u1Gz8Csz6dHIUBR9+5ghmG
fx4XG0sf9naQmlJfjanZtxt7+9eCA3RVQD7BgOV3ddiXE/DzF+HKsrJ7Ua4MtxVU
DvLQMBOGj3el4k8X9MQGxoYA7iGGiLT3CPI8vgSEkh4Ag9tXblw6sfghE+/HMOqX
hTV09NaVOIjmPJ7eW4JKiwwckI2jtUDiJEIET5E1Rg6mZKOH8h9DEdVm6o1+YLTv
1Nv2+meX+r5VnbcA91fSrZqZYemc9y9ADdUIDuOfCOZybcgoYSPC1522Y55y7iNB
PlD+aoLE4Aj2l4ktpBRPolX2zrRdZxvTffx0wFsYLogym1rQxpsQr0Rb3xulPrdo
cS6x+p7ZC6wmyBFpBY5DiKdPgTmknHicunbAzMuZkuVbcIgvQq987CtURg5OFHwN
YHZ6Ya5l4q2hCKEUBQ/+zexfOfM7heTmlF74/Yii/+DEOlSQqa+vt38r4LW76duI
8CWxTfCMfqcQelxJEgHLtq63TtsILn0yBF4nmJR+h4xXojCL8cxfNKoMSl/53ave
3V8L33g0oraYGfKBBn68uBE0nHlFUF+ainOw1rdJX55VSzjzHitCQ6tMo2pY1Zqm
qXiH4tzLWJWBjJ44JZTg8R4n64h1FN7owA0LpGf+CiNr+NrDJnEX5Ssx9SX6vOs4
nZybP2VuiPJPW6P9bxIfbAXlgMCLAxWgexIrKnjNrv+RiCyCCFxYjaWUWdLCtA6w
/j+hNuNfmFxTfUh1rrKXlwJq2tpjK+p8lLf3ZCr5dma86iNkuH8RBWVMbjTvIcOe
jAqd+X0RmZOJNm/zJWD7Tin1izYCDYAVA3P8rSfpmy1q8bF4TF+0oEsn7XZugRzS
gQmXihkPqbbVVROwANbsK/tle/sxx3pkLarc+vfxDA1Dhp9+cX/vZgv+G0Z+rmSv
vMPymnh/KMCT8lFFCfGBZuzAq3dOSPiKayIdIY1paTOuhKkrbqhMm5UyDFqmkzTe
V5HqfF+nfFD+u2W1E1pvd5d1VHzQHfkX8IgJ60ZE6Y2/JH5DYGxttLfGiqaR7NjB
jlADYWuNaaK5S/GvhUFG48igvu+O3cl4oWcHpjk2+Fu93m5RDP4v+uWUII2JJOu4
Fp+PiuYxijEsIsRfNZHXquI52vv48KI9dKTKiSUubiT+aw/jecOyKsEvd39vGMWi
xxLF2WVkh5KxUnOAWRxBTDgRu+ibx+HvSOHtsu/fcK6zhVGGaFseXz9GmQPxCmyM
n4d83jqdu5mrQS1Uue/DsLtZRoJJKbtJ1VVcPLkTUQ/RqCCuA98L6L7QxyB64goJ
hodaIgoMkfmAqADMF7ItejoRONLmXWywFkjyTxIV6zdLgWs+wDWI8T6rZOAm2j2e
syrvDAoYoMrW18t8uQk61soaj4lxwu+s3P/aThuyvfry+NjjSO1/HW0eyGMtDmSI
RrLyO7ZhkIG+S4Mw4PCuKxXxiy4mPrri7CuYOsRkhaOPyeQ+WfcsdaluFFFWcpMD
c9Sd2RtbV/CHslMrQB3GmVXAeUCdc1DdzeXqoUuUe+5+B67Dv5JQpq/v/kSOubFJ
4I/AOYUjsYDSr4o5V55oy4i9dTfEZkJv23oNQlXnnNBp8W0s+sLmn9VXDATKPkLA
EE1VXd9klFVTg1z31RjwO/mCHjmbgHguqqDj2woAxQPM3/MdHbxrnXZiDGynxj3+
05UBA6hHnyTXmal1NJrMHPnjw8X028qhLlfkHVbYZL3thNxhrrD8CyQXdTjAmh1o
CDMyCbTcVwzn7U7ErKRuyjzjWwXKgdzbeS2nbJt1K5WaFkTLfquvJh+Tq9G7mL+B
PlXcR0jUFjM8ublirOFzILxHGKTUr1NKVqsqsnA0gwLRD1xnlXRtGEbiBzOZxMLc
ubf6VKBfyx/G2o//CY1im6Jq4JrtLyjru1Fu+MVMlYuvVxM2j2oADYCNXXZue75p
6yyjzB3leXqm0vkKnf6Wr922c/EtyIwkdHJ6duJ7RL1pwM9sFT+Bc83ys7FPnm/c
eVn4XO6edtYeWk+xqsHZ/bAONG8XW7KB+/YUmaFM/JvFAOTyCK3QJA4HWpokOFmE
mNHlIfgielUfAtTjRoAsQ7eu0DcCjE71W653aCIsM/bDYoQseUn1f4uKcc1mhmBF
2Rm396ooeR7ygnOMq2S2zT2rnew70iUU5i3C/St3q44iPuMDQm/7J+HpteodXpI5
unFOaueCHPjKdC3htbqk+f6s8V6i5NabhzSbF3SFYeeOT3e3qPBgFpMQ0aU9dCyh
dGKqDWTrO0bO+xGb+XZePXgY/f519G74PnPXtE20WFg4S475YL977EOI2omrfFI3
9/aWKAq9cgG3KkdXvfo4GkLKb726/eecdv4PCoidU+LH5Q+az9CrAw8psvOkIi/a
vxTUU6WAOL11NIdPBmn9Xbj2Gqm/SYe3EQ8ieWLOTVF/MoJW2UxFurFr1lrFbsgz
C99qTU2FrpKKFIo1dcv6fD8BSSRyfk7ndHTZV/J4n6c8Ogw1+8fNc0d7gNgoyvkZ
ADU3MEhlH1/oMJAwqQkCJJq6SmC20UgcpO3vxdgyhnaLPxJDIqDyVTZtn8ZbD0p9
BRGVp2mssAAkiwI3BXTRSjBpdCtDGiZ58VTnpLD7LR3Z08xvdaVdhWi77s+v70oo
/XxC4LEgk3cwZg7YuGcJdCUKx6H2L4yX6ByFVmpXgFceGs5ESLGaI43SIHB4/Tr3
YhEnEDHIpLVC28PVJAmfRMoq2b29jJV9g/8AXqk6KJHyTskRBpx2+K5IqPoRCMKp
TT5ccl/TQVLIO6ysHpQkxSR5PQpE27XA0HMLlNJ5V/Yci9U5xHfhDIRamAtz9Ite
+9jCVVxg4T6zgVZMzQmbSqybBYhGOQaZKik80fttr+impH1OKMTIGival+FIkX4w
MxNNMQx9bxj5j5tBY1kLbl4dNWA+pGnbitSESUfOCgJkj2mH2hv1djG7UL7DTO1S
L/zTCWOgEv37WUD1UJICg323ofBO64kWiyts4DjK6V4a3ISDGMUR3UUAzo+OBuTl
Ufmhpz76id5/GD7seUshV7NyRsGjdUJFDWzS0W1lPQgvNrcNUpiIICZ/4/TQapwf
VvNnFMQ2peu2zK/WfG0j8lJedxhAbTE1yuhoi97VlEJv58h7okyCScF/YFFG85zz
hMMnC7bMpAk3U6Q11HeD3JUsChpJHS1JzpbUCXhUDYQn+3jMtajvHFVFsMrOkUkv
wNrN76vIVfXxmyrhyVY2EU9G9FVcnYae+NvNUJhFl9dLVvXx6yoH8rCYTfxN0jfg
WYwO1egT9e+hoY6js1fWWt1Z9QImFk2HK8PPnGkEDkEzB1L69CQHdNzLM4iN+z+s
n0MOMNZxQm+1WCQPrzISwV/yzDkL5lMRFdVOycIRByEaR4FY0Kh4ay7ebIJdhkDs
nGT2bJTFi3MJmSG7SEGJ2D6UQ15EzZs3xSFcVPS6JU6hOhHJIc2+8HB2ymwX028G
ttVELY8k8ORY8G1j0HWl/XMxuRLAgj95+OFEXWC7gi5lFj1VdejpBAhGkFRQx8wo
5ee8Y1IKYUUPP86CyqGWXHH0CiDqTEDsGkXT5tKcZmAsXl5gYGmRwbih0FS3BkfE
zMLFo8ui+/gunPgMfYxHhOQ7mIMwfcmAUY3apEmJLXgdPHfoi9ISsBKtiNUl2hO1
3PNlO2BOKz4zsh/K58NYLhI3JSwlS+5hEmp0DElKIjhQferINRl9+9ABhh+roTLY
E5uCDLOw8q8J/wloNZwiqEtij7Pq6x5MozkOmbV/KPUriOcNBLggJwqGeYS/F1W9
MTnSfCgGRal4zIVljSwGnWjhdRMiMX+94eNN+xqNQA/zPBOyc+eZyJ/aRSBUFMvT
xFS3ZREehyEqJ9RB4OBa7YLlOL1ZK1vAXYfV1Ky1gfv4ir+C5muShecF+zYqXpvE
EWuXcTSg9rev+IWu8zYA0mIAFpOTJLOOEEmgRzIBNdXEVo2+E8gEaU4ydwOzpWvr
ONTNfuLg2BczSC+ed4Bp+JaqUaQJxBQE+ZK562oX80M0Y+uxW5yFR/K2JeBio+f9
K50OfoRDRFo3F0CUW8NC46B6TeYrD+VMo8C/4eKIlaRa7FLx55PSbR+OUYWoCZnR
fmUCOe/V+Oeq5EgUd/WsKVWbaoMUDWxbD256mAc44fporTtPzbZtIaHmxiKr89F7
GP1dtlZ5+yB6eTm03l7LYbgYjUM9xpa4tolxIEu6WfqWH1Gl2pEmZB0NISCWqZ5b
E/579+BSv3sZrlZ5lVa04NUOZeE9S3aLGbceOULtPLXFfJ71TBRk1ULWhZEWo1CP
qWp60Ulm7O+FXpskJc2pcuiZWsuWTfCcCxenOUov2pEdB7i67plMi8GPjqkFGBnh
GUdwCC2YbmdC6AOlrOBEvUBS+lh95jJCONeQMbbhVvzvZz4rSgwd4DVahAY3cotM
tf5vstWvWFnHK0j/SiwaiYp6fpXHFLZqAlUNwIOFE+FTPRsSvo0VSs+lLnR6MRUH
M5gct28D2RJFz0IMtCNkMuQ5iY70p7vAA47s0LiCeA0XJnETNUGd0IJ6MxTtYeGF
gAZ2QQqYk6BRLgJRT8+6YTijRp1E18/Fi2k5lmLEbJijvkbPRyLjSIKc10nJ6Jbz
+PRNOnb0ZBGd/4lEp/w3WrMQw+UREBneK0b1hJ+SEXHwG6iE56OA7+NUJnKcuV/U
G4Evu5NtDyGvOga9dPUrs6Z9xlMuezdurlNgEh2X5ujR9de4dQc4WJvXil9fE4bN
/+SjsO5ZqySJ9IyiSsSJfd3x+x39dWob5UwH0NIUFN8hkBIHjzZtK+KOztApNj8t
+6sx6xEkOVODERm2vacHEg0y/tsDX993SxGtumKLkmtKGRk0WhXGVImQ4nd2A8WO
1X7iAD7g1u272bD/NxX1YAZwSGdstNHdblRFCvlicX7pnXTR+ZZ0qD0RhE8iPDWH
XKMQI3duhNxUP+w4LqAdiBaJKkIr17RXnwqioR3Pg0STZ3NLs21S02irQ1CSFqiS
IIHrnI9REjGxtFnMxYK9kc5W8QPiAoWCW0X+pLE+Fvemx+MxSDiDNFAjyX3f5yJv
kJANVrN4l6q65NVY1WQyJqe4AEixql5tjpvd6M0cNBQL1IPLxmgb84Qeaa6pLMVd
yNwjmLXViHXYT86s93on3GlbRTQ4Y3Igfxh9UKcQutTDwhcdw6MlmRy684EYus+c
HejibrRpZj2JVCBRCzChZPtw/KcoTVx3KT1SY8KTVhHFolzfacf/FknSurrALefx
si9QPzNAcMLpQZFkQsjofg3xgmlfsFS/ECPCvY9bUROHfGYXj3yAFG//E5X+CxgO
2xf/m99JeQkrYEZfOfRuSgJ4O4k6LFIxLDKVF4msrWbZFhefLHwLByLP0MMD3iCd
Bu52GGxrsaRPwuXOCC2ysbLYeWM/DQqXgltE4JEi8augFKzjcXbcSXNS83P5FmxA
ckkRjlBfdswBF5J+MejBINIe0z0oFarr6MqD+itOFVOmbsGgnYVIBq0YHbDQiljE
wBZIUdQDOPgz+hl9ov454sJBip6BU7pmfkenq1A1t66iVa6wiYkbHdrQOW2Bzy+A
JAP1O8LqXVo04wGk7sYA0qt1/EE142A+D8HjeHU4m1TLCV3cKTNTFAzf+hGADVZi
AygP9YZOzeVkLYexr6qLSolZB6BIMoJ18pHe5CL18Ia9Gzvxu8WVaz7XeF/l4Ycp
mxS1/IApg9hr4DmvJNqELgFpJ0lr3xQe6VZB/1ie2YCg93XllDz7q7Rm7ZaAFGA9
hpJkQgtSTAswO8rLY5QxAaH9CeFWuBDuJ0r/C6a6O4B8Dsh3nPZBoerku+LQWMzP
RZ43ozLhMcS2xY0FbvAxL+rFdCMJ4Xwb715X6AnBtqHlRPqEba+KKloM7Ya4w2BO
J3uWV/tzqkhzDgByuNk49RNkThBumjyiSGYCiihlM3JuZsmW9uX3MSAbdiRo3N8F
2+pQpxVBnnK80GPzZk/eouLOJ/LrqihatXBrCXJMwyNIdDCq9Nd3B1iZhkzywJ3e
rh2CzmQCF5aLIoRhcf6K6aH53cO2oeTjHhaDBzNzg74W/4vAHAXopZZ44jBT9Wqe
7QiZCNinZy+FuQQn67s2FKOZr6VepzF+n3xRWTVhhQ6SQpKvrofomW4PLSYPQFoi
iS8uOT9H9XadXjQn9yt/pKU1Bfk4n3IGkmug5FffVN4V8/jXt1Fdq9ANCY+oBJJ/
Bq89Xh5LD5gGf7zFwEw+6WwR+v09tOAnxzgLVPIdOnpxcloEzQkaF7tAO/Xh2nJn
x+Yj0mv0syf5s2o9q4iko3zMZwVj5b4VEOeb6SiNqc8P9rIqE866ItF0VLbtilD6
FHk5RNKQo4Pq1qx6KTqTueVzdO5Z+dxKAvVlgMOWpdqe+KgG8NpkWq3PmKUrr/zP
jS+irij0KiqknPiqcrOhubPTc+Wq3Mf5+iwJVKX9u6BA2txG+oWJLKFDlmmsVuar
2dj3/EXqPbxZPfR8jMjBmO5mmefKfxj4xylckfmIX9uw4HqPRMSnE8qhPm2LEDvo
b8nlBn0wmrKv0/U1cTutbMJRwYpYyTxoyXLgbpA5eMjYr/eSln5shViFFiYjTEXJ
92LPbRaAStFrAFwMEcglCrSuIwt44zeQ26K7Lmlw39NFHNwCRKilDlJ2FOlGKv28
9ilSF0/LqKxGG5HDacZJRQYyCUrUX4rTaNrQ8bxQn624Fct67eQ6Q46w8wS3VoPJ
OfIZxufonu/smA5le2Zmpq6y/GE3X3L305AwvXgmhb0YDQG/dq9OkPu2pd0psas+
3Bj5bYf07VWL9FmguQR87r85N7uvwcypnqZbABgcwXaslQpGZFJI7zTh3Ub9Pxha
IkypQEjlKwGHfXMM5hw3aHWCG/uyn1VeKw4GfvjmcNEfvfz8ndOgKDmipOllA9oa
/I++Aat7FA8Q0EYp+Flm0hDAiqVck3joTY6PBy4L94ebQbRZL9ucaCdlR8ZJ4CID
NTYOnWnrqqLYbHZ4UVK498ycwKW9hhFV842TlyX3L8wuWUa5Ymo+IQzyLDrj9280
wxVdf0aVEOu7y5VZQUUJT9mfMWg2AUUmkljJlotFme/L1nnO0fLV3/j8VFhi8DA5
Ae9OWPfNiBLk/F6xrpaVV2ax1Is2aw7QAQ8D44VOQk/03Ng1xeyOK0IJ8jHWRAXv
WFCI2AV99ZrSiWOxorMUEZaPNIuGsGFRcSqdcjZTHdOnaGdDgOGFp5+hjKUPKk6n
M28NV/fkpytXJqjkA9UCt6lJtoxaSH5T5xtr3TkACpwP80+liYdj4zok24LFvmGb
JZvxHIjZ/62qdILOARpdUZVLpihpq+T0SCecP5vCk+msiO0rUSnq59LcyHa6SpGN
ErkgQhb7wfqz2IcVszWdO/492x/1rKBUw0L5soER1INUr4cWxKbxOjpNAKV5Oy62
BH/8FJAXyQY9zry/ahZPa7QAzW3nOmBD0ZbO1kRQuvDXsd9G7po0s3FyGu1Y+oZK
1VWMQkAUQtirwR8R++6ByjkXjiFL9YcxTvTmFEOn3h54O2wJCDT1eFhvW3k0qE7w
GQG+pn1QVtqqxp2gCBRw7d6pOrIWYpfua1F0xVZo+gCkW7qUJ6eFob0xAASW20rX
eE3648JO823Uj9A5zaH9acXd4bOmmx3T0dAaFicdz1O11n2soycmtVZMUjs68Slq
fcVVTIgV68mcIWa94pkeuwAvYK3ZYReBfTUvbdl/AP5RsCUwPP2jWlwF6RpHovin
CD7xNbqKIqH7LrdpshbWddmFTPNeVUOz7cPqbq/K1XUWLc5y1pdi7Hy/gD5Hil64
8qYaQpiwAyWLGflyImjTglLoCELs/GihhVr0NC68CHyigcPe4ut2cUpvWZoJtpaA
4kfFyOXouL9BpCRChAQ99x4LO1nRFaVpEsSUW+L5D3bkQ00PrquX6VBjbcHyQPIC
YctXbYvSKajcFw2SOw9J5GLAaBSnzz6vFHnpqKsCcUHgevIjAUrSHlqyLErBD2JX
CVXaMyset3PMGH9VyROmj0WiigfHOsmZxn62GFTp2gQ8sfQNDN8AotlFVm9mxa33
oksTrcxYHzMbLEcJSIR/54c4EBDdnu9EeEKoU/ovJg0nxUgv7ajW8aYQ1gqP6YnA
LyRud6VzkNyaprM90ZqNHi4IaHJgk/P+3oBA7cD3RE5LtdRlDhQUmnUtq5AkuXrl
pFUwr0nYXZNiylolJJ0M6U4d7+2eZMHdXtDOOHVvvucOr6KUU3LpQ1xdsMG1/cDD
OF5Gk8hLrGMSYYODaVNgEZQ0PPVZp9Dlba/xzRivXUYixw50z00STWZ2AjWaiDKN
PfEMtXVqyaYuBVa/dufsCHX37fhYORLx0pXorD83iEq7+wy0++CNz61/zYdFncqx
Du/WoRUehradC0asdGjTiEWmEEpE5RdXphZKGlBvNvwkMUDCo3dTV8t5QWUrl3T5
bXgxYM9JBK3Hes69xiM1mz8kT6QYoS1nJ30eJqGQymSNEn70hKiSjt0y7X2K6Kzu
Wp8EcO9i6ZlioLYLLemsqQ+8cQZTQTL+111LsrLk2YlQHr+1APfrozB7Nhql17zx
QRGdQ05qu8gKZQAdsAvgdPk37REpcWWBdton07uISP/uojCf1a34kaiMINO7wY9Y
8SqQHz56Hm7K5Ex1mZoz60Ct/AjulrOF1uNrwelFuhvgMG9aJwrq7Xz00hRYmp26
clGhfeAFtc0Axuk08ySYDMwwmEv+53JsHcsA78VNKHPNMM7txNLjcu6qvUtWS2e1
B82NuPYQecJ+jwtsiRX34ERoP5MsRcIOs42vrNLj/egdkPBG7zehL5nohLy0U6y8
lyM1mGAS4n2iOFAiAvhTgEbvS9swYrPzAM5FbPz4BJ31po7VwQhltbJ/aA00MAi+
OaIMXECBH6hIPEf8imRw5T2Yw0NhO5NtkuOWF7xC6qjXIZborJSs1d6o+GVkPKqw
NpnE98FEL1dkg18NK6etKd0iZM1IP8bDYnDoJL6poddEhr9GMGCZY6uh6XKRXhSb
w1JdScdHqSQEyMcHm57n3ubawi1wqOD5C68REH5ZAbYotMgfkqd69iItUFE1dhpO
4dePJihjP/jMyqBtJDxoIsMANvy+JNroswV4emsd7oly/SC2xv+0tDyfPVpMy7ft
SvlVvuCusz4pj0YkQPQVteJgLZeEO4nO2DIep1w7o78vStXTqxbd6QPOfjHXR0WG
1BwMuKVJuW9pQKO3Xns6v5gHr6/K5beT1opbT6IPw65G70ZMJyQYB2QanTr1QbvZ
7h/5YLGNPI2e5sYPfUx+0C0FXW44TreZRrdbGBiilyGpwEvXXhR8eEkNwov8vLOF
AXe33kA2GBM/maRdw4XQpN6VJT8vaPBN7jdRROsB3QwdbIV1/voCqzwa2I2a8Gqe
ncNVq2mxQzVuIYAdQVojivNWSXZN5JcePrTUC/KGuzhhmZJqd25x33X5/YsAMi/q
KbYW4XZELuwwuMJI7oVFxvbhs3ZiNo4IK1rsc/0Z3ftFOJu1FXMniM8LJExEe9ka
h56OlfulvejBym0m700vKt/AY7qlLOwGPvSIMtcS/xJIL/uIFERgvWyX+PUrTckm
V4vRunBEW79CblmEipAFWA7NZAiM6pJeiRWlxza4pJl/b0tTtKVMB+eMzbAysL9c
sjodaj0dmNL0xsjhpW5IuT/vT7AFjWadQLel4GQduK+7Kg+QS73L7VZY4k0t+aoi
Vm2rM2FS9JZ5ENf1SHk/R3ieutyzRksk4bkRJXT/Mdmy+CbISbJrdMg8FYVrLoIh
kcWXjn36NkUkzenOxM+bCdoPrESBJedaKmF9qOKBJG2tcyQ7bR7Tpuz81wOlT06R
vHahbhwSsPEycce4u3XEVxKGysxkZSBDoiADB1jHQTslgx7LWQJ3eUHqlVVs1TsG
+WnO1TBtH438CxbHU5+qyr0+T1U2cxi80gycOSb+zBinu7LhTriKGsesEsz4tKwb
1oCWIcQbxUL9b8wme16zOYxxMHFv/ATep3/Q6Pb5XrRyQ6NtBSNOYAVsbh4Gs19i
thO+KCf5iGJswDmZSV0qPggODUiXx1/a1+Z2ArPaWVH8Vi1aFzZYBpsbtUkeq7Qn
3F2GFSk63dQnHpAlN8ToaIuLEmyKSZtu9coNPh9QsIwkVaYdZ6JXf3JJv5uKvu0f
GfqoOUsJwyWNdUQykxr6RGH8UbROntbdIzlZiHg22gEniTpihZ1s5XxWmcUNfQFZ
euVzVrEVr731ATysdbAngtfEVHCLVjOGNzbqjz8l0pRBL59UjG2S9BqW67plFoNn
E00s8u4jjGiLmT9TFoRfsawArzmPWW4vEnDHzAy+NaKOmidTsNhPZ01KocFwpQfG
U2dF7QsaQm4Ni80C9jqvkjHeVIB1887xX2tYLwtiDijueMYUaI4HT7sXTwb12B1w
LZmlkvpTBxT5DwRh6kH/XjUtgPH1wiBhxUcXi12ADwAJWsbVZGL/vfdMe7e0WoaJ
+zCtqhGbRoys51v6cFjJnaGyqQft4IgSPUJNK9ropsJYImotjpIvDaXPI+I821wb
Qqfx+4b1E6jRYWAsKxMYMWl1p2SFNAgnYONR6OqTeU27im2y5lZOd558t38D2zVD
PVOU+xpNBzaiP2JaIUGWnvhoOQmJWQxOM0xpYfZvl17jytkHSoZPO3Ogs9zRNpAb
c+7jqjuUmnjDIR5INYct3q18D94VmoJMsVB8gbb5Ad57aTGIMHD2Z+IobK2xWxE0
cS9G9C8KUbGj1NYpa0Iy1kKygginNUSdO7W6pXi8WSKRd9w08yg7/XSP7P4hH6lb
tUlMeqxRb7OefLNsj8opUIweZQnVWW5kpIABsFLpZJ02Ae0/0biTa1XmP35R6t4a
iflthvyrNJoOh0whDr+1ugMbWJTwsDQcYFoSoQ7HaKs0HE6zJFTvf+TaUUb1p2i6
arZYscLcDRBWVpAV6FK25denYr7x7hL65L+J1w9h/AHzBTouXK3yDTgwaMKqib2s
DtNxBtlx/tbXpiyNo/G+UEBf6H56rQzHVovhD65BxeKMKay9pUUSmaH6ZgecfP5W
gZ7qxO8YTqXEN4UTVscPr+y1Ik1rwGk1Yq0t43R4p67U7y+VcSIfO07Zryog8Dke
RWIbOR2Xp9718Lg8MOEMvRR/EcFlMQ6kcWlHHX++1aoZUYIdG6WQldgPvLH4VcMW
CSex2XIktAQDo0qGq6igyJ5xcJ72+PzaShPZqVgSYsOnWkHuKCwiyO2AmjtHAxeg
DTSf7eO51U44Af7jCUGFT7O2c0+NnWqHUa/wfK4RSHws2+3x0LXy7vLmzFtGITuj
wP3k9fhWAffu0ewHVj6Hmbqbij5TrXlCxokmpfpHRAFEV+hxI/95r7N8Kblr8LaI
yPW1jUX39wGz8rFNr+qCyY/xQuqtE+lRQ2CxsWH1v3iTF4lohkqpBWt0HsKYO4Rz
h/Kp/wHEGWnwDNp2LJ5aHmoEDSg/Y4BHGzOeARrcigAs74hYaUlUgn9hsDfaCi0g
2SzwqGGzinV3DFrmu8CVEBIhoymFk7taY9FW57yqLhJ0B70yh8IHM6vJ9+BdhynP
nkSrtcizmtUoGh38683kLSz2WsRvQZcvEhaf3J0zNQ6sCQU86xREajaJ3zrpcYw1
NBkRA6fSktFapZn20RmVw8bheKgsl1oFZzDFSxlClnzx+sog0lwcRSDzl7ckkRJK
VRnlsEAJNm+R08T96w/rMofPnC1s4OVn487clrvtVvBgEhJq0CK25S5ZuypgHEVg
sbdHVSf7gu5Iv7x8LFkh3sdjX1t/rXGTlaAYleYWP+KEc7aFs0HWo6gae0o7R/Ko
mL7aNKqgkcMEoWq92TZt97y3JuYjZyti+EaV5aFQa+gfdobHTOlwi8St1kFiJEtY
5hx9FaXRLMh2qiErytpkPSeHHddH3O7VkfHXa7VhM4cbxEeReO+4sL493fquNBVf
H8Z+5C0fd4PlA00WOG2jGYXzun0JoU0EPlQoaIDiutvp/NChi0jI4wLLIXz4opsb
4sS71Be4jt1ii6mxi0OVlPb8lkt1exwKR8Xh6WKpH0pjZKaM07v5sO0bbckDDhj/
ij+9omTw9AGD3EW2bt4bEDsrlDb/gLwMw8RunmZnyHFXqpEkNpicDNRBJjQ1hZ8U
7W2M+bp1Zjrv9Lz2FzqaUpUh+R9p85uViKNW7Y1LNlVxWGKehOWT9Js0DOn9609I
ztmYGIkupNnGWvMaDLGJ+eabJq1vrJuxr9CBd2W7tmpx9PoP0Kzm+CeMUViecNLB
5MEpvQOuMrF0pOtYO8J0uIUhZeoVdXBo9aFPXL/Alq8e28PL8ZQt4j/A6/XqOrwt
Mg+0F2BsZyyclfLYdbF6tpEVKNa85KsnAXgkmYhsUXxXLyWRfV/TU5TCSj87E2F/
wrCdMmcCFUBEoW0WQG2Ncq/glxO+pzZdsiVoGWqdroDRFf+e2RM6HqJtknoCznSD
NSqBmINUMORas5lVf0MDVlNYmz4zvurCM+VI2OY83WCfJtXW09kG85fyICSAcZ3c
o2TxjTSyzSpDNrkbyhGgh6NbLj7/8z3anusNWjsRuNVBvda/Jd+pDCZBJ9UTgtwf
F3kOWUh0V1v/Q6hCk8iifx/M3RtO4FBWEcAGs8qrAIQKVnkIKb22/TY7a26yy8zm
rX6csKXS6GGmIkwknzo/dPrXpSTKg0lJYeLBLMr8I6HABZ7XlJfbIof3E7QPhsXd
p432wzqCKDO9EY4iOe8BPO56noGUVU8S+P80CRNVSo/FajMTukk96hH8Igx3e1iN
pVypVuOJqmfUA7WXpk3ebhDYHbr7pKnh9L4tosYUfHw9uu/c019QZaFXBkiqt+1U
fPnQz38Zzhp0GLhcIquRRNFFMhA7RkK2VZ6aWhFqhnqWWmisT/FqZZQWxfkbBfk/
D4JYHFp4y91MMlcmDib1ZFcFrtUlhLyntku+Xx4z6cM5ZI3arPxAsBfxn2VzX85x
iEzXmj/jKDx1EBd0VRcPf7QZbktxMDRk2nKh3war1i/TDj3zNgALaA75hc5ylmkr
7aTutWnveNpUwJDst+iX+C/kljTS/hNFnDY9WObpDwf7gTUE86nwnv2uug2Qvoh7
3Db4FLLyBYXJaSLW31wn1ow5jLyC057YDjH6XVuk56j2612skQwwEwya+bGMbON8
YST6Hh6v+2fV7SyiHpiRxCjO4O662W9AsHFD09KXbPdIYskEzUW6TPqJLGoaivRW
QLnRodptSTkNdfbVEuVX4sUz1pg3En3aUDriTYja5GGelVKSbjfCXmdmP6IuSGE3
TwykJq5vjGQZfyC7jTUi2zsbHPmvwpBMbv7N3zqaaWSCU915TIay3D4XeLSAfGYc
RdDdOHGg2SMhe1RbkCL6Pmu7Q3IJjbdKriTFZeuaOhl8XZPwIHDvV23T6Dgvbrt6
nVA1ZOywgZAfELvelVpxDxSuoMcBeEzxZN2sP2GrzyrkFMP2jJ6mrVwueeVBnlkH
vLMvay+EXERSmvyr0jaRPRpD5MEWB+SzUXkHIN+OBGOUDd2HrsIgCfJTAmZU5ivp
GOPsCRCK7dnKoCtpWLrqAgfPnfzySMRGrvUX3KF5j/D8DmdpCw6EqYXxRnGcGngf
VKqS2ov5SMRj9TozMxuDvCBdNSuiLagtiG/+zm9sh0tCEOHD2nKbqU4pcX1QwuUk
lPN4IZCZB3DCfhL2QlJG/LNM0irWz9bNWVmC72RMspjLWHarOvNd3rhEqPY9RceK
CYwWEBS5xIm3zUx5MmIItlL2doDqgtkgiKPAQCjz3GnLUlp4QASmg/HCeyLHT46c
Ju/SxnuXqBnOguy5pT7/c/il92qIiPgdAvkDzZsVgIUTdG2k6c3QK78cWbun51qO
nMJMb6TlZdbQczdc9STOdEX6jnzcv/4RWIoJlZZba0xRBZVT7vRxQSInmhe2i51O
/vRUtRSvczeXbSYIS5NpVj5CLGqpB9Aka3U3OC+3aQeLxMFlNWabykk4VbYKvG/R
al3ssvZMxSpeY8gxX0Uap6khBPcpTfw7l/xpemQACPX6m/I7TPfBQ1+0C0BC7Q9k
WLpkgdBmGoP1ffM+XT0IhRWsahFw5KRzNeEmC2FwROlxDlcq8ko1zWqY7o7oQBwj
oVVpH6mWqj4X17R8wAHb579eg4aucUDikHf7mYSlU5dibj/8wAhAUtI+3zbiJdh7
iwyUUdc5N/MHfEuABKm8L6CxsOs9Kw9UEqMfz7d5wMO+ohdwYEpkwSHhPzf+OTGE
ZRA0PoCufstr7glK9qGs46EKwodDQz+5w2KU24Hlb6K6khCG8O8G53dWDqPxVhko
CV3X6dRj+f7OqwCGexJ3/hkTEej5k22hxXXKl8eK3o0YG0FeTwdxhuXt4e3ZS9MU
GeENwkyKYhcE5ml96zAwB7WKRMTmXwUSx9EUwK6czACcB2nHfYfp9d/oTLMT2zEB
t6gXXjJMTRrADlNLw3XyAYFckPtWBIdCHKX27uGC43am0DqTTtBQQJ9/MFwJPnRw
Ol9X/Q4QEULoToE1Z69250i7WWR0Pj2oJYSpnNsS5WjhTx7DYIst+nxLtFPfWMNX
4fhnsyuJSIl/dcVZOgk/75wOglvpkmc/vtaP46jbFafg9yp/yGLXBccdiXnkr95r
M6aoN8PhsRRr+ymNpnBFN1uhto6BU/BhXwXcDbJJt6OG/Sm+xVJkIo8j5BG6y4a8
/cvzlV5CfiDrsIuZFs2i5fryvi7QirRwlcQUfFTW/tZwOK/vzWuR9TgsL0dVcy4G
n5FZg1cfUU4MGV6qd38WDBiQF0bNNExbRwgQX20J+6MTfAwPBbZC1EvPnlqiKWkk
THETnJ9LX60LBkL9QeNWnXZoj5wfrvUxuIFWfUh3O+xA7oEgc0cP2oLl0e2Bnx2r
2ioKpcCLiWWTxx+trWpmAFqhZ6BHHELeYuCsoqvafQveCqF9ueneejbJb5AGRDjd
vfxfGMEkJVqTZ23ZKVHZ9r3wOiBcJI8hBdP4D4CmL0GSY6gWx8YKv4MuifGCHUjE
ZckUxIYFfRxkUy8BRjAql856ZB5YJZO+CihYGbayVoDerWyZOcL/yvatPXg5aQJO
ZsnJncoD0VllffOKz7J6e3zmPqoD++ZdYD38bfMf+AV/vGu8sqrt5Iqdr/lFP1ZS
pUmvejdco7GillfwPN9uz56zmZq/ryCMw0qJ2CM6ZI+InIIhdABbZZBgVEbtXojt
9923TsPd7Sm95pPE8PXx5IK8UK9taYZi2I/O6ojUpHZ1lkElI0R8ojFRr4orzwyl
ZvK3gKE0pOoO2OKCY4VxiybkHdl085ZoTDzb5h6D7TXiyRGmYmffWY32p7TCPmDs
837AUaXtsW/Tod8S/m6/7EEyi9sI3ZN7DQ5Kp4b63xB8fIjj0ZQqFeH/zE9eA+6l
td1/NcCzwK8r6eHdf2IAtMyDXQpz3z0V/woo5i8zcs/od3H6s25WWU/Qqywgaihe
CIYRwGUJkspy3Mnqbws+iOGPwtPAKm5nRoBfjvvWzDuIwIu3RSx6eYhLEvB1Bfqm
1EIuYSvk9Uk9zQAWtw3jlWhK5OcjLIIbobO5lJpStqRNcbigVhTzCneIrASOqdTr
K18MNRA9yWsMipA9iKCyYh/idavQ3JLFKGnXVl3MFH/zhlMvzKgAVUH8jeXHfTn2
ZGG6Xt9Im7JrJMeAvsBdditNG+gE5HuJKtDIrvSPQzZR2nCXWl745HtB3DFsXdW1
/R8yHssMq7U2JGTYcMfqDZyLlXS3fEWzmSWdZNw2xZ1XFIAtTvileviEUZd36znu
Addt/0X449uQYvaiD+XZ8z5hPru/oyJk+cDzmJnWyxLpKXWZ34p2h4BjjiNDxsDx
Ky5hR0sv6DbwOMGc91V/f+kCbjDArEkWwVmrHGrSIE98DNmHZdeK3CP3K/gZjh1O
2x/rFkdc51JxYs9vlcBJPLR6YmhV56U3Cy6Bw0XukYk/jZzkG1qVPJaFBUlUbmB3
50Vt+JqCJK5b+fArA/j02X4c+n1ceJBEs6BElew38fZrz8FDzjam9MPbGls5nv1C
DuzQh0mzel1QsgKm0YjekCLdDMYYMJkVBLOwch590Bd9wSdw0tCaOt/PPKNKV6fM
JKyGVrDRJfVWfk4nLLZ8gvcHcFSY9Zs1z9EyaBPgSpMXeJnvVgSDMIgBHpwaU2MN
K4D062xOEAim1EB7CulBkLxrXwvESszyccPnPOyYGVPNcA35Pz6p6Ed/2BD5Fd8d
M3Y2hMFxefYFNZ+UR5Ar1skRbTikCgKgnXLdT3D1h2bIFq6eShxtuxNsDDVhHhld
yn8bGxuxRoa6pOwGO4yczGdh8QXjC9ChcG7sT7CujElYKRT4ngomXL7knXNJcjkx
2zvJ7pCPPlVtwreOqxtGDUGIYsHoACJdA7MniXfqcNFMKRs98u1LRAu4ajWIPDCP
WYYkvTQ64EhvdoWLgOdS8QL8oXzxvpd3jCQ5H84dzq2khLw14tsUHJFXexeGB065
WEsWdfRiTudGiLNBWvttbeliZabGRhQ5sioh9LHFlKa44LsTbwMuFNfJHl08XTOm
lUEUjR8VbVdbYUKEVHM7qmSOvdn6r+fiTMQUE8Rox+jMWuPz2/1hntNUyNRi0CW5
eyrDSHBo3rfaFD/JRKwPW59bois0GI1PMTvZH7uFI/Wk7nQsLowOSBRc5CoYtHN+
aoWcwFUpeui+LoHqeZaC9wrRd5cgBk2gATzTkfhQP9anG2smsiA3d81M58RlXl7e
6O32t/atu2/8FzO527WEDny/zcVSrvrszsVVAdfMSdnCqnOCAPcIBelVTdauw5nT
08wwcxMJb3/GY3agxShYo3qXWIloW/j48s/R0BpO5SYjPgxDTykF5WP55BTcNge+
KOJ27Lf7JvLS5OpWeNII3tPvpF5hZm18LC/OLQvfyCe2Z6K65OddjAtWZW4OvN82
shdvWpXDKCNjwQY7s9eL5bFUHVfEl9ZhqArVQ7avgQk3rkcbNVRPN2eTM03CCrhU
D0632xB6szX2zoowNU6nznwSrDhaAW+FTz3SXz0/7pTtRj5YgudWCa0bz0PzHCvx
8azdikvndXUhuwsJQ8/NvojP7+5c/5WJTdv735L9elv4M+YU0NibNW+sXGH9bakT
7a3LtIeXbxThwjhvf3HbEMg+BQJ0L80VhnQnSiPNbDXcgphrvmIpf/zciEwVe2wX
WygvpgsqSATohXyjBkwELu0BXHufZ7abLt08c0XhR0blJiud2+CWadw8mxZnrw0N
kgbfvp+SsUiiNuXwO0IgK398KfzPXs0nPe+KO6GHRhmANR2QAnyU9U0mFjFlkAnG
xPY0dmsUk/9nVyUeVed2JdJ1BQTlsxCg6YRgohk62WjEAB7+wP7jAyzxEvGvtneN
U+OmLP662wrB55uZC/7lSkWSm3ZOCOp6HUISFzVeTkGy9gKuJ1yM+9gytQx8ldz/
yiSPaLa5k8U0wV+gWnInlnb1Pvrg0fMAOi/fWLs+oXT2r0dogt9/pqRRkqVbAq8q
JaohnXMNqZwfsD5g825jNb1CPYKwfYVEmuQjmTenti8bcAtpZxe2wK/ERNCxjPIK
z7nA6X2OzuCrDeU/p5WD4/0miLQW8nEdy060NGayE6ASgVHfr3aDk+IzinQUK6lT
jpvypajdpaYB8a1HkrINJzR+ndKcP32GOuVXlEOP7qNWjwKdnm9APL5w042rp4EW
VxyFS6T4x4vloMCrtGNWMo2iRIEfqIYdwU7ewiNWGPa0hU9WCoGI5X4E6ovk0Ocq
bNiwgTZEkbG6pXLHzzVPUJtv8ITLVP7gy15NwicL27StWtXASYm79JwAh7xI2Tkq
ZRD8iVNsi4ny7hONHPeb+8K5gAXS6k0brM6wB9DAwc0i8F3RkiSVXHKqkUlx06Vk
Vjkk4Zzr3hdMaRKQcKVjLXBBGnRyawDnjpiOvISJhJ+JMWuUm7+e0luEHzdp3RYt
FeGX1CXTlq4TJE46FNOG+ZW8huovJ+aW20O9kDDsU3HLVjzqOLqpfIzJB5gy5pIy
UfkJUs4Pub0oIkq3HLOQxw7gLnSPukMKJZWfPMypp+rZg6Fa/9r/vEh9VGwVfXIt
OO0o/bMgWTZ8YTuiYIcJnRf995xflrxyZecRJxd7IbR+vL8/wep7m2wTmjhpS4VH
6l5vB/FoWRfsIFDpjY6xM/ziVdw0jWAEWwu9mYm3LVNkVXY71nst2K6rh5Hc3JZT
pLjhX8D0ImZ3D/0qnPJ1t3EZcX/aVNG/L4AB+adGbA/Ivn7Zb9PZRU8wac/MWaHj
sC1s6OglPqkcWjFf5B747ChlxJaLHqZ2pF9ddrjCFX+jMpJ3Y7NhbS50dgfnfmSU
zrqW+Bin2kfaOI0eA5YnjCNYZqcBP9eEeRHJlml4NG/Z+DfXCBqJsmc/oJO6wwXX
RiEx/GWI3LyrGKqMfdq8zaCM5B5VocNJ6KWJu7+23B0Foyc6eNxQ9sjsWw5NUkcv
9Q+9Ncp7vMdZvV5dpXgpSpSqZWfKwOupg000zFZBNPK58OVVmzxiQp1KxuPNNAEY
6FIkBiLwWRJlZw22XoaoyY+MJOiCpUHfJrOoDTfmzV0UyxqbtGlP/ba6sX6a4g5x
CW2BPx/f61GCTovcjSHZOKkTP6pb7+mMNwaas5GIJq5FDWAs5wkeL2jAmbCYCYsC
gxfxPQIYDm9/oA73eN+6/QtQwzod2jYFu/B8hOv+LhVipKzqDrxGoPZMQniVYXpb
mciQtGO2oEDbcw5m/LJlnJgRVK7uRjnWrYrsmOnU3ZrZqANwtyRygYhIo9j1UtAS
vTtgjC6xovE+Rle4pEs9S1QXBr8EUyUpFi5pnjy8BCdSKWsDm5VTmCoa1c3q1wUk
YjtteEu696Y7xdWfReqClTW/BZt6s3EIV/F36S2waBrzLFTGnVyn4fYdVAIP4qzi
KZgoPm6jIwQz9/qWESGFQoDj851nnQ0IZzCDA/rcqBekyUu2OJc1JB4VmuxGmFrP
mTTD2Mh5NqmPgJA6AtiIQDh/CmRcXQKfEOlWbzk6LqcxculID/h2m5B7we8g55aT
PWMWjnjyTk9rTL7rwlQ2CnprLcp14dbv3ura06tPa2dIn6JMZtyJ7ULwDKx4k9lD
1Uws30/U85/mMaPpM2Rw7tTYniZmtQf4fI6odfa4w1w6DraS+c3MK6ed//o88heY
vv/NTMLtSi17Lwe7CubI+4j/BEcTTpWNwJrQ/E0u2st3kfn5ZieNET+79cNXDFa6
BTMCUeLhN4wwLrlvVQAeFj4VLgUV4Dj6QQ/Xuz09kzwTCA0Bn0sm67IvcdYR1nn3
PDNSwb2jpci0RsI+szhL2gtoFlMKRJdliK2mCgN60ReZh7tDvHmRCPHuTg2H0dxx
p4nIpBZj/gRTghHaOEh0lLttXPzOrCpHbeX50Dv/ya/yWc3NsHnaJjUMjyo0B5Ib
fQzhlti4p3YYDHl7W85Rn3HWr6zcmmTZrnc2tmx7ROd8XD58647PwT9lEfsr1vUE
8iZv7N35Pyun1PD/BSPWiD1ePoXWVJePUUU21OEdKsmznDcxPfyck30z2zRISAT0
PptBuuxps9LiQGWhSTGFfk9bbLVsvG8G+MVITB5eygpQyGjB4H+EekWWQjXyKGds
Ib7qPt0TF55ttaQaHiQwK/qQHvQpeE6/NzrijAbZxVmMwe1NRfEmSiRym4YXGZPk
Gba0Ey5e+PPXHbhRcofmm0SZA0v1pULYWLR4R3lcn5vzahKPWzp2tw9hjWxwJucX
cwjed1Ez1p33S2ClF4qZTZ044J7WTcW1I6P6tRs1xUVZ0Mac+ONCQQsnt9OXqECS
BPGu0/u8z1oYxbu9eTn7kdtKYqgsCcOLFrS6uGD/rotr2PEjb+R71bzYjOyE0Rk2
SHKfqCCiWcoKJ+ImhOG2mbWz6mjcpkH1y07rf56hqeeua4weKIzyQZEJMYxoatjr
u3ccVtYmOUnnQfIp/1334XEAB69v2RjQTIP0Qw6ykilXnZJlj8Lhdkb63FAsOide
GDGN7dFW9uaOPhluzq00H7iZHhm9YG5lM+hB9sL1v1e1pcNK4+vyX92oLpWhF2fI
DtJyg8Pmzyq7yY1tZ6MlWWqhbJEs2sRuYnvyYW1Z4MAEgTUn9uu5+M5lildhl21x
Obxz6ikO+TztN49BP+E65I7qfyVSL43yPGs7WPEx99VUt9cNgqhEB7WQbpuoOg71
TVfmdcCl9oc1kg8HW59i+LKGdDFjiq0ryOt6Bc2remPQstRrP8WWgrpq/rOjMp1H
v+0Xhra9PEIl01QuvRElsBpzNE/mPbdzkj4reBONwkiFHt9lyfMsSOw+9MJ3PMOx
ttAp6hzwFTDKrcM0rTMoCmyr3eR7HFzQtsj2fAvJ+nc1bGOXdOP63yNi42oyJUfc
EUg0JFaYaelQ/TRH20stCPBEHkdr6BISsErK/qQB/ShOm+XTd5kZ4G7QY735RJsA
uY4OUm8x1w7SbCpoGqqDrXDEHMZieJqqqTgosRCUWNZJwv2UtudMRupFip+6vLKo
8uLIYf9GTXqSdPfelcJczJRYj66P6a4jeStLmW3U9nUXfu79tpua5OW3gZeqfph9
5L2zDbVC6wTec9qphh7WvDitZxVtjTRJCe6An0XTckyrvKWWPWh+G7ji3GcxDmOM
m6fLvOSKkSJLVwx4+J5t3Lw6yD4qpDEflQDy/hnN71rg52gF0oeieP/qaoM1NQ1Q
Sj6u+rrmAzrXy3sKGF7NXaG9r7cemOHsl0r9LVUf4wO6JH8tvvTf5rbKXzaUM8a6
OAJ1uixxg2yT58LYXGS2HFBMHc3QEKWmHaYGqrmrT22WVXn+/RLHYGFFoha3UFvY
SqnL2LUkZsW7Fc1D2halDsx0GpaIR6VAhsRYflzgYVFFLRrlAEUm+BllCvgisFTP
WAJ+nghyKT3QDFQM5uUunHvww2FaNKX+AS/ZQT6opa1IvKFY/1fi6CDQV4eRrbJ1
i6SXEGXtGDHph/gvjPxYwAWJYEQxfTW86KTBEXuQHPqUV5ilu8Fgb13mlCflp6Oc
SwNPljd3M1vi6zUXnBXVnBt3PdMYRlXjuHyIBQsiGzxt6Knafn4+uDJWuJ0dVnrX
sDhDtasx4JZZYoRdsvpNCVYoTgfi/7AdbViV0fqtCzkiLX7Jd27oKhvaNEcISNKR
EEDVW+J+vAKyosOFIrT5Tfh/k2OCSLco0gMc+nC9yZwR05X8wtDhHzW5STdDBqjt
tqkVYA0/2KF0M/73vSrCUcFBHOYpH+FvQaqzNEDirntyguQNIQAPftq1ZidhPJ7w
JRazDWZ8nJbqFUkXiOKrAOgOMpdkPZj03d0qgsbNUEwFVmsVrVm8DIDYf8z2xvyk
CwVIc3OZNKyrn7hVLBVKdwG4MUJaK59rQ+QCYUFKFBdsem0/Fz+qJzDWlyiu13K6
kRctsCrwfY6VHkVd/dv3FNQiaStMPgjbUd4K68amQT2ZZEkwBF5Dv0rxpVOysXks
ffkGVO8qxWLWWjG6VtkK1PBpLaMH4jSEeC02N8jlskogJp6Zdn6dyB6GXbboVa4p
3YzIuwE/IkuiNy2nA2Cm1X3syUGBS06S5hyh7Cyh9hr0MZHXSqCSMqYdQSx09+dk
iQkUpLJVHOsfPVxm8KMSkWHHG3G00DJq7CwjrXzDCQIC6/FbCLGmlSUwE5OZ6kU/
7U6wdhDurY+Ltq97ssTPVeBr89xRVki+7b6y6FgDhvvcUqceyBIP+sBlX69e1Uwx
hnQzfPKqcwe68vS+kzd5he7bYZ/Zwsl95mYVUz3oLQwjOxKXgLUxO8DHLMVNL+HJ
PB6IlT52k38Aafv/JNEwORnHWb2Dz6MckCRxQpuQ8p9/2Mr/E9mG6wb455AvI0bB
T68TYlU2jajD9lShFrLl9hXG9KZulKyfN3bRhl1dUbV4rI9V7ptb99yJjOY4IUOu
Fcff5eumlDwO1H5awo7DdOuQFpCnZEUrCTzUYqMFoSeBYPf9CQSu/Zp3MnSZQ2v8
kRekAblCttqMlHbxIFj4a4Vp7Yes6Etu8NjOhBrzZDhC9eV3bVTBjFZi4LlthJzH
qoHRvswygDDCQKUeeP1Wi+X0MBzUXIHPos7+qD2Q/tGTZHBFy57VGHy698iRj+o9
IGqUm6nffzobqYGlhFpRIbtGE0F2n2tIrthW5UnoISvA+ku0rRPTjA46pTqv+BoD
7ATkEMDM99JHyOGedcm7KeGqkhZbqSW3yqzP8QoQxWf7mJ3dlfMKGxZhijQLbSnq
cEsQb69POoTm+zCZkChKCP1NjMcbjBTPyPLWkHpsHR76/1YJqop0DLZ2PfSZDcMw
BkyTfh+MtGY6U2S0a41F/9THzwa2OqirhVySmhuJ41cdLXNA6iygfYi4FNzk8a4b
Hqq6yEp7flkAJ2HjrMv7+0jjSUjH3Nl7igFfncLq9rAEeiI+D1BrCaVLV5Tpq01s
Y69RAPzYPPYsH34G5BRSrS2dxl//i8SB7MSgjx6lQoxdqkNoKgW+u12OSlGJStjt
HY/8JtKhu63+eVFfSEaXFAnAztuKVQIHowziYMk4lFNsd4BxKcxZsnjRZ4G3lD3P
tnLlPgJHs0ibdcqtAdRCv6uAIzISP8/xF2sfopjSkaG1gl96Qwf7wdso80OZgoNM
mDXmbxVEC/VZthj0+RHI9Z20/PeloF7xUcBrKgoGHuvlSbOKVbQnQ73GtwuZnymV
kpfKQfVGlLukd+VcmDd1t8DaCseOJ/JJjyyXctYjxwaYa1yUwvl7ku7LYH+rcvhZ
WtL2RB2pEVeTqYK5rRt/G9ln9+FqPTsaGTRMzzqcKx3kUf78ua6tYIqGsqf4eeMS
TapZ7daW2kB7lmzCIMlqhCkk2x7Tftn/YzlHDiC92X9pPIesCiD9nrn3RbCiWxI5
dM4JbWP4IQr9/TmHLuCfyha6Mf/EPPabEZhWBopYRvK/0Om2YweDZj6kJDeIBTsv
KDm+ODjLl7ZebzVJYcdSmWoLWgTfbBtWevnxL8eHNGA0/ONP5PWgw0BaHtjS/ODy
OwgrrfCEXc/6GhmtVTqcrjPkq33V5l5hvX6Qk2BgFXFkt4ChGwx3CqA3E+dqAMCF
4p8Xa9zsB9nF+KU1OOMj4DlOJyqEsfezcYqejTYgjf3kjWbRHLUgB0RNxxv/AKVt
iP0ZMGL/5diBF5uZfj5ns7mt9nd+MjCPfQ/6M9Chdhys6AqvgNdJC3+8BlKfQise
+hGILsndk27/8GEPtlyKZw2bJSRmHeeudf32XhqhdNe/EkDyPJmHt0yfHd3PLmGo
fIeRayUTJv9voued7fqoXnZKC2aPOqyW0bgw8vb4zMOI4nVlnvNNJnhb9QUc9DG9
c8FtCezGwmgiwQSdy4BZaqQnPaxRfZxFMgX8PhXD2E8Yr0PSGiU34+d2jZeaU5BP
tjq0QYhGI5QL/OPgNuORprjj9Wh1CqZkIEXhrbqTNarIM+8vNS44mhVJTuPRE3AN
I6j6cCRBTWgkwegBDNK1QE9T7LaFc9Wrzwag5LDlKKjYFER0ZyB+yBNVUODjFN8H
XZ3OJMubev8AozF2kgTSD2jX/e2hiGZSLS4GvkcVRQy6ZtCAt2HwbE4DO0fQuFtg
r6KivHut5B0I30wcujpdO6VbrQsuBb9Fyib/P42IqQcyp5ejL1j/jbShpP48uMPa
T55qlwKczBSSY+Mb95HTEjH7HO1G4guw2UV4o57vX581yqNYRJjnh/0qlzuycGnw
uG9PdnUIrtMBwZr9o1YQlCnMeRSUao7RnoLpPaFbDxTH6dxVi5fww1sKninaexbU
Suhcv3xFnLloMsmnsBwawtnZcyL8wWsGwy8naK76Fwa6kXyWl4Tz/R+bi4h9lZDE
gJh3yeSV7uBr5hiV/mVjqCk0VuA9xp9ooQpEUUg+6F9bJhL6cz9roYmPyt+3rVBu
n/BAcoflbMyZ9AtpG1u8IaXk5b0FGDhtfW0zEypMN1gQYR612BZyTLwOpV/sHEdO
hbCsWn0je+cXebOXH7NzWxfh8i0tRo7tH8uuxf73peA5pSGBAXBF7RhKazFk4tED
Yji6JBynP5ox6T9mtQhZ6x6e6rfW8Ku3PzenLQ5tJaxnHvx8XBGPhMsOkE06iuM4
lTJnPTJNWE/cTLvuDBEXT9a60am4ktkt5ZybJFbTYcmmAXSZZ9boEJifOYrJxfop
ZYLO95HBL5KMn3FFUFrMDxFK22YewanInkPH/tPosocDcP2HOgJZzMjHOacNKAhY
jPPnlkcO+/gYaOOrIw2T8aPyVw6C4k+PC88HSRKiXjkjosdaoZy8NikwXXoPUCB9
rE/4CAkTokvrvV/q4VXwu8NC2xZCBGrMdNLDBYHKKRXhKOkXDSfqkd1eR3KKMDHH
oLnukZrsF3/BfmPVYqN2WMnDbjziPK6JFqQHshumFRqGZAzYO5hlmP345qQ/kTyS
2i+3I/KTo1ObyHUZ9sx9DX/LRh9m7thkfqlbmM1VC/jUtfAnxwH1T2mguCEgfxNk
JknJnvM2NxQ5jSQzNjFjlXxgQ8lFkxh3T+d+2mXNj4pP4hybr+WEu8cgdXt2Lz/7
HDweyqkHonqxY7vZXlc21A7lpSA9PAcLxDe2ARQhfNM/WAZISPYINVU2MW28NTZk
kQAxdHiN3vWoj59lDPdb+vNANm0VN/1ACAlt3wjAkqGNdV84hcxi0Laaf9EeN1MN
QfYmYv+I9b3mIMr4l/xDHgj4OLtxYirER0Nr9KpXFAPopfTx6yaI/BlcVQN8P103
gTAGZaPtH9dPrxt9o0PehUfJ1HGROFWNKUnbt2c27d7VuqnkqIykxoT8XuXed7Vp
BO+t1BIaiF3NjrUCw7AB1wEByvJWBnRfT73sjId7zqu5HLtjGT1Rpn0VsDtlhflN
xCXGQa3Q3MuAPJ+Aupeu7UxyJ9Pp7M14F4GYmXy0zB5XV2FASid6vZTGxgiZPrvG
hy+xN4CWGNC764FdtZRzbhB1RQRLVHRKc4AfRh40KJHxNAtJU8TKv3nPgzB2Kp1x
Xc3yFCrJQkSZQrGvFUc0nh+tveenA/jOtT7YZ4e9xUTzcoo/nSZ/fktyQxoISs9h
gzx/mSsBn2df9coDr9dNRpbPJE6LLZtQMcl/2NvsYGd/K1uesdbf3tNN2FBuUneS
pJFuZ31Nl4MBwPa1oy3cUkDJ8pBN5AdMVyIA2Cxg52tzYJM/o17yXCOEMJfmHP0d
wwjRgAzT+IO8kX+iJ3pZCA9iLbztEd+N6Fh1dxT1XmCs7QILaQEVXN88p35XdmOk
0e9QRIIJFuOCDSulknDodplujf5PBnh7IXfH8MpMGZajSJoanB40EGyy2kEMv9ft
qX2kbVLQ59Ga7vfX09nvyLzaYuci9dG37FAGo9AxK9UPVewOiQmz+59j7sMIcJgM
Ay4RZXDyY97+cUbTNe7A1Z6T7BIQJLGmxW7nW1FrR+aweNxzD0YcO/l/VBiF174c
b7fqpO8zwL/SJpUxtqs2FcSGRjyNtO6aMqv8NcjryJl6xkMlxx+HonOdXCcM1e1o
kFos8L3YbuVHXTFymNIRDbXbli/HRP3Qmdn7bzv2zEGTNcBi+lKRssz6KtnOxYDQ
Hsf2+skZfLso71+BZyu3nAqJfAh3QHzEnTWmy8eA1WKWJ0FvQBDw3YpWHhNDIu2L
rAbSnMlth8J2j2rzAGIFQAOcxRF9EmNfub09ii41/gIOyO7+fqUkPB4JQDQy3IlI
49/7og+MZW7cArZy3kjZ2A9GeqDiVTTu/J9Z9ODHwOsBT/5Z2SK+xevjy9BA4bXu
Mo3V/71+Y4SMOiyWxHQbUheeJ7ymCtez1kuWuuEM6yPNdILjaWxqZSTp0NIOXQWr
iOlaptpxNbNWuePAVrkPom/eHlEEopTj2IyiLttVy3ffoYt3Paju4kFFXEv8xJnL
biuUel7KkZx6HzQfaPLsyg5PUVGtlktuw/VVqLXViYekPBIDed4hv6YuSID/MJI9
2fQo1PudmuQs1PtdSe26LwBKa0MtDicC5J4NBiTnAprKAnegJp2Rmq2y9+xicmWy
uEww0ZnH11bMV6zH0XhZ29pKW9gdAWJmQmwTRkVkJkDbmprRfakBp1RzOJtyOrbP
KDXC5rGvRVMZB/f985w6UvqrfQU4Kgi+39Ki8F1NdTkeWMTNiPAmdZ+N5AL5ur5K
f6jVjxSV5Lj0ZvF3hOMatK5dp6EvygrqiBQ5t5qQzMNktFDDrt87mBT3c/YLL90D
4AgS0iGfZVFaXQPqU6JW5M9OTuED5JQk279xIMBf8uB1FBw0R/S2TdHzz3QTmfuM
IsksX/niYAIDni4B8S+BrqecOonq0BcqCjavxBa2duyhMBTPPfR6eOYkdBrV4uoi
HVPWXEcyuHxYNeI3MmpEdVuXp4vXCfcFEZmMd7zAvEKrZ+jlVtiEEQ/xUxZdXjeV
N5I7h+fVG+U7auknRh84+ojZaE8YITGtFWqZzrSxRrTopYcZsDcZKlgc1fL1MA5V
JPw+X6WVu388BnIA0trI5tlIJXu8CxusJF5G2cOdPXAK1JvS6Mokg0tN1P8VgTpq
OvTLioz12tXVt1heg0gSSGTowi2+OJOAnhrOHfXB9nA7gqta0khMx3b+Xz8x3L48
tmClh9eCD9fUHiqmtEfhWqPDBBNuJe0t/ku7tjDVtLe0FZp8iKkY5Dg/9xHWX/PP
f0aGhM9/bnLPPV2Cl7KggQ2dTxlquKQk8DpX8gxIkhNOukev4hRKoEUqEpuI1ZmG
EvJD4486CNG6evCHelQY0BljCfx7lNBLAaGwvxF7CGVzrLYZBCkLTKAJfDj2/ILp
U/tXrgcItYPYKBV8l0FvJHcgBsZpQY9hfBMyNPKp8RYumQJAOnllOF5wRYXlli4j
opSCnFIOt4i/1sJSTMhLsjuJg70aGjRj9p/t5x/hu7OxnpT680b/mWxbzu6+WfHm
JQJS2jIkEGets5uXu0WG1oxgv+4/MI8ccVCsUp2R0WYCCb7KWG1TNep8neE5uAvr
UHR+1g0t7XbHTT6Hhl0yYc+Fk/YTSFE0JxzKFaXDP7UL8RjeWpF+QgEuR80Qja5I
KW1QsU6mj5EKZwolF59b+CgbH0lsN14scWO8seDb6U8MtnK7f4RK7ZYZxoDu6vsY
2fjfEGiFH0Vmd3hKZ75x/JdgN0UYFqzKqwHZmRunF8vfc98X9KRfiA9VsP5S1X6u
eMCuXCKiH08Wm19l4RPeIzRYgMtHlxjhHhy6qMIygjrfVXUfhI4zUHX+ln8mbfYa
50XYWy51eFAibTAfJUMT9tLrlfoeWQtzHORYr+wNeL7sFYa61GvuMqo5S7P5e9Mk
aTVdwKc6eO6s31YS0eGqUp07HyOJAhzfoB74GqbMzCHvQxrJgYyNthpND/F/dFgX
3CN9tCOFrRaJLfk9uWXtth4EgejIik7/DtYTvxRQvtMefmW0J5fuDHBnyVa185AQ
qlBMhunZ9/BtVL9J9UgZE9gV6M83iXRFpEekuO3l6OeM5za4Qr+dHHhbWPAGDKUG
vtk7DiF5L3CBXxbkcE985s+h+pmht/IkeV2gXfrqmwkOPPy2E26BAcJu6B1mx2a8
pkwZECx//2eCA1RG52AtXQLkIn9FxjTIbtzaOMp6bre9nxTgV5h21imvq5cJFBrq
D+3icXRq4Gb0QAg2bM9frGixOiIyHo09SsthuSq0Oj0PuXYP4nreIdCEgeBRO9yV
IKmZc8DZ9Kn2/BpfrfCfl7lXYZtS3j3350ei42Ko+YOGWt3wyajkx2XVtEk4ExQJ
oiFUnIg/AiJo1NvHUh+PhoIcMUtdv2/PDL76v7NrlMkRVyNcUxrsQ2k/eg5IwB+y
imC6/+y7ZoBi9mOY9FZYQQJp8tAZMGgdjb/aBSK6bOg59YBFofcsNhnebVQFurll
krfNRkuKzWSLCNTQoSQ5WG09vAYRRJ3R/EZkhF6yN80QyXefi23DxZPvDzQgs+sL
YdwrCloB9YhQJDwt8Iw+G+5bqbeOigWLxCbH+I6ZR/eUHMXlH5hR460PdOzyJ9nO
qph9J4B5jrP2J9vW2r+XNxexnwT97cQ9Io5u3/xIsGpJ1wW5/J8luXXrWcab+x6Y
MxzcOxNEeASGFd83TrQ8rGpWXq7Pe+LSX0N8BpWXdiACZfxUooQnPUZY8DG+X5il
xdQ6Fl/OrqfHgKOXLGDAut9os/PWxCQcCRjDBwohj6mS/HrwHjmDGBY8HQbx9WgF
SXMPclJEsS/BeS0zJ7GqTOnauHu+5ihQck7nw64nEvoSwmLsiVYYnKWFJ0Etdk5V
c4fDQxtOY1SgRtqqDVAHu+Nw1T62mpjc2T+78YmOexaRu322+OunYQUqzddhYc36
xAsGqcEZhmi+qg7iUUDbWuoSfjWKHS3/1l55qiTvmkgKexQHbZbhq2+FY57Ou5dH
ngY9+zJMiNYhkDH5EENPlGNO7p19p8oDHMOTlzXMV/xS0+QLx8pr2xkvENIWbxVq
GQ6b9lG1kOUdob99lHKwZN9IlwUK2GKraFQakgdb4EanOtCBCTsTDMHwrD/rN6Ir
7SEmZBJrt0HbpoVQ4sYIjC8nTEtf4Z1d/zwwMALhmn8cSsMbha+tOGJ++UAwmdu6
dr4TqyAFo6Cg8oPdr9oOuad8wADXI9ls3agYPXi1Ygj2UuUb3kmLTLYbu5Tp2zPI
nDaOVdbfMjyMXs3XsRfoo9eEsZ69oudf/R7/RLlUb7V/Nvgs9nyI5H3M+4Occn73
Ay8jCD+3BLYM4HestTI28Vg66Qz+Vqsa1ltxj57362fSZvmfOiLUYwvGwmSuTS+v
vd+aveppO+BkJoFPbF3BY/MBM686cjLmZhvDy2svbGuOcOiizAB1JJXm6i3vTcL5
+J+/7rSelvxTUCjtdZCAgqV4N8PsM5R6109RAXuQi5VM+WF2B+O8b0KFoBExJb+v
ygCZ75RXlyyryx8wcLEoEesfTyag6fizLavyRZo0G6xuimS4VLT8onAqkMO8bUp+
90IH0HteJ8J/b8OWkMReJbMP8S7frHl60F4yDLydqAk4GEzmANXcbYtSJPEXt08e
ojeQb1UDZu5jeJObV4dLraic3+YY3JbvkwJG4XSWgcds65KmxfJoXIh+Uol0art1
aeG9tYh7bIYIwbfKY2IfPbxo8hSfNuc6qkkYj7qbOfanOYG93nJLVzxfXe5fVDYc
CrgvD8iBShQleEv689jGLQW4jyltsS5CvIx8OEOve5vsiGiOl3ZtpE6JI8jZRt1o
vBCyCbakCKDOPk4S10c6gHNvxMCztVNZcRwR4u1rly8IqAQgbtRBV5yQFjQe58Ok
etNEIcwyq21USah4UOb7K6sGC9GI9tR9h4iQmUgXK86iuHVqN2IzENRFoGA4meoF
VraG1yQUFWHj13xifHo0dk6kKox1JVKQa0TZOJydpfg1PfowLz80Hf6SD5lXroDp
88gNQqbd7MSXLQ0gTOjztqVNVu2s7uaphopUOuRL6lvKVvTqOqXAb8PvlWP1rsCL
2E3KouMDiQnKTGDcg/M8EuqWltQWq0fgLyZH8re4qCH7hdfb4GpEQEFporuQCy8B
dvaaEnKPW8/4mVQx+v8b1y9jmS2aFOudnl+bA4lt7b0RcfscUIMl6r99tIMAmckX
Ik2Ki0RQ0e5E5hORFu+b7iiCEIaXB8dmnu2lFD9wKQwBj9NybdtaIDqzvDCK4qRP
Ds08e/mADnBqC6H/55iCvEk3iO/e98DG00EYSKCG39vxn5bZMLNB0No6IvHet3Lu
7WWlZbSXMHokTAVEbsg+1sIwwqwaBzkN/j/oQubR2b9IiimAYT4umHGiA2ze4gVr
QoGe4Luupo4mZl/54y/NG3IvajaBkdBk6CJ4QApZR1STNrvBrJzaFisUOQDc8fm7
AgyMHSfEaDmoEwluOmPbOKOHkZs61Fg6JrBjvqOzn0K5319W+rpKyQUDI3nd7lfM
Sl4/seKttsid22GCmXpzPogJHHbv6c+QoKIZlKtR/vLfM2eXPmdIbJQEzhC7rTzJ
SZW08b/HC8PDxzQgejPSG2j2zXJM21M8pUFj/lEUZSqXHJxHOE4VZ+ECs8UxRvSD
AsYr7oGXpvOzSWYkB/uw2kJcF5/bCDg9n0VLKpPETJIZ6iCNy0aY5jsv9SrZ2AKv
lpOT/mdbrqJZeNXdBBGbRrwtj3hks9/jT8LWKuZ89WUipMQZ8MlQfkySrQDetnez
7kMmGfcNigvLZyRY6noZUt/FE9pBUEsqX97OghMBGQ5QL3Ic281Unv98O1HNTtze
IjCLpVfAW6+idz3CrMzV/gTaaqR/OXUuOdxC2QC0SILh1g+EPFNfickZLmzWW1gu
XomAZeS4L1L+PcMPnpX0uabFBZoi5QefMbj4cBZiVYh/PbJaCJEFuCpEHNkpdRDH
zSq9eT943qP+QczSY246fG3Jt0ZCyY7mFBxQuzozFzhh7ShQu0fW2KJ+DTNazuVm
Hm4dDEVAdVlThqd+yXsmDKC9/9Jo+t165n1oGwX76Rehpnmgt1WhgSjOLEo4J5rI
cZMumg+Qe6PiHacF3W8d9NtU620kQdcpdbmWSmiZTrc31jVrsJZaAPBVnlpo43y1
m0MKuLphmA6cJ6ja/jm49wxPRxPgiocpBdTIGp0shFoesud555rBUkObxFjEVGbN
tHc67lV5O6iZYZQNRx3yccpalGfrIM89ANuN5IWc5Dw0f9Eo8jsLS2Ss63PgtMfk
pK3Rs00eqk3pZ+SG2/DWQG8EcOxfq/pJim5eyl21dNLWVmI2LKS9Ql2FoK6yv94b
C8spBZNF3a73eKZFPt+zkBzRTN/OR9tswrgXeBhKjK6UaODsjjzPM56QdJl/ZwlM
gSOuw3BNqrniSfZwt/4KKoGnhUFhhKD2+f7MC7FX2HR2Pty2eRDfzeegZ5sNLBma
RzGw7H7iOZFVAFJ/z8pzdT3OOf+j4reVsKBEFfCnn4i1NmdKp6cPsz2JfJ9ZHLAR
v82zWHpfa/lG2xU7EdBr74bQaj+LsP4SjV0ltAX50RQoduk9gVTHfFb4G48bVkwh
qWhj6L80CSUvpkZjPbggtKMevujfanb6AWptIndcV7+0eN3pW1VkmBSUsHGG0PFl
FKvL/Z6jRnleX2ceD/3zwSjJ7owZzeDxrpDAr68pNG+2sgb808c2H+p6cXBgmwZ5
GJLiSjRoRPoH6QX4/mNkk6aAMkfIsdK363fT1R7f4TstLeoMjx2GNbOXLK05hn4L
TUzHtiI6sXtkjcNacqo1uCWlOqfVruPbGmRVmQNyRqeWB8OvzeEJ36oAG5/ohmec
JOcaTJmmDxaf8ykzf5qKcrFsyum6rcd8VAthv+Ba3RQjSqDUw3AmuFAkHdiHQpye
cAUH0H7XKCpy2m4kAV323OU1BSrw7zIJsJxsKgBL1haaiTm1S1osRNKyU6dNkLH+
DlaljRfz+hhMhNFZZp6TwX9GD+3kt0Pv6ffGP9DzE4na/UZflQtPntivT5ivmXh7
dC15vC3YvCHAqCG9qHRzmRfKaAUoViAaccTgkezympRN9PYCq0q7pWi2bc/M3wVU
j97Vow98spIld7WJLfRD5I4VSpBSAAnH4jXwVaRXpVKiE/cwx5KfnmqFcluXzSc/
QHPCVeVmuhaKMLazKPkqY/H5VmIrh/ybuFilFHnrSkjfbNMZ6boNysHX00H6NSpi
SMD28XSBDQGAPXAdbb6e+5/hIbUwJwL8yABm4Yvomj9vjgE9R3YFEpTIGusdLNqk
rMnkzaGWhRR3prPgTC/4D9ydgMTmw3Ke0k37JcG7EVW/mIOaxlzF/Ou2/YVgbjWU
8FtSVZ2LWpegfWvVp6hELf/Z1mfGDn7GIRo1cwrb8BDikrUO2JfpLVgMXhYPEffB
Vo7OZJ5k77w83CXp7jpN/gryspVSVOW/RIt3E9jPtq6HGfZH7rg9xl9X6iBLdzHL
ffrbQRyrdRIbqivizjeaeOjbiSr/SGqdm0p4Z/ycCmTMwYEUWbCPOXyACGh4dD6v
3SSevfTK1BbVEfP6GRYCemEx8et4quNe3/KqeZoZhf3wYpB8v6T8Ur5MiWbTlmSC
KJHrOd9iDXa1taDbZdX+8sevcpYYbXQDYU/Edbbpz0ciN24lZHtHbQZ0wNWzCx+c
Jscr6XLWmAWPw3H9/c+452TBMXx9n0XhG2GW97kdIvUaFyJRIE6qmNXYxjtx2r70
pGwibTs3qGHv9okQ0hNMnRG1sJSOkmec+tXxnsT3+eG0YXh5/fKE12e+V11j1L6t
F4y0fHhvNHVj2ibfNCz4cHZ0ukSv/iJUbeAwFKQAZts6d0uziXst87akZXH4Jr7G
MRGAjIc1NbpQDGb70zdS2hZ2usma8R5F/pdE/cOvc23lhHdVRJH3EAHtiODIwtES
WNbjA29Po/ASJ0IAN0GwLHSYXGDAifSxmExuTr+/Q/I5LmXVp6tFinKHf4cgy9B2
uGB2VEw6SMyr9qWpgfjjWLxqK/xxPUAQbGfGWFjh+nwz/q77SdxxlzAWNG04Pb+A
jnGui8QgheIBi33G0HZe1KmYOSQasN+z2fwOnOkygA9e1tJhoqVcRsDLohtb5M0k
CMOI6uuwCkSqSI9rGLA2ohEbTMHpzaRMvniTJlOYOZ/d6jQ/D4n8J0XJ5lGpAtHC
LOJtZkcMltfYxJEETNHvWj/BCvq6c8F9CQpeC7SI4ttPkLxKPgYqoad7Ju5bT6m0
UQ0/YlHcZUr+6K5vbhcLVAS9vvDJHKUZvPuP6FyUAcRyE6Rhhnw+y2SwhYKbofc/
HhY+aCq3mzImbV4sDw7GyMxhLN/o5ZfMToy5FHZw1kbQaSATZiGJu44BbQAEZd2L
qgF+4DsnKlGCB2f8h839JN5J3Zf228+KCJdcohHDhLYtVHL+SuamuN9Dr9oc1sZ3
Y4WhyiU/TUYwKGh7whVeLPlU+mnlBse08MbFDrAQHouIJEXZ/ZxVjDd6KrfIS7w6
fL9CD0yaAGnTHNLWlkfFsvM3/9JVeoy4PXTTHmojshwBGJaNI6/JJo/NqpCGwsGo
IgMIhZ/kBctCqqT3NFaISVBxvXlG4m76aPC9ggylHKbUfto4ucazYG0WUmXJG4WE
fhk8zZkiKt2H53yYNUcMUuHSMzOSkvRWBXMIJ4sTdS05ueDkQZggw8hHpKWImSvF
UZRk8lj8lr9Bul+MGJytRirlzEeSafnnvDsDx70P15euqOedLOAr8UmDSc/rnA/e
3b/RwnAAyywW45LtVdvY9GFksqSDUncLkZ9LhtfvNmGVvIlWiP7v2qrgreFq27H0
eVTLHCjEuOS0uHhD+oWS3yVpFJpMaNUsMT/egxbPcQY4j8OubKYDP6aQlAo37mrK
nwNr+BRRINlykxJRRE1wIw9qPdWUNMQIPk7xljbHfImAXsYkRCPEuY97i3H01EY7
ISbg5feqqDq2x0gwkEogIGHJHcH6jVj++v6sRnyNfN2IjU48q8kC1NeGri5oDUg4
Q1To7iUgqO5gaFXeRUVGzpfkWDK9T0fUQThO0vccnrtDdN1wr5kcxNbqbVTCX50M
Eqkjyfq+f+zwiYpy7KQGaWRHzeTn+Rp1Rq+49TqH2lXaHmkKpXDsGAHN0l/fOOCS
sWHTNpGXjWi+1Jybcw1fb7azPnJRpSIkziuJhpubTRVLxRxXHy81JNXMnUoghv11
0c3inFy6cTpNt/L+bZfEYL6peOcCSeLEw7q163K9tjncluqPcCts+LYIJc6IyFb7
Cg+NBb0SJtmCSSC00uj7ukt8qV+NE2UyjyOnfScFea3LDOYf6CZr0bd0CVLRys8l
sNt2KSYP/XJRoiaowgZGUnSLhiK3jlxAijmRcQq0DjEQKu8k46BS7RtDuLr4IgfM
8Hh7NNgzVSebg9oMoleSgfpT5RCmyIJmITehBEM4vxQlvYOPz2mXSuQ98XE2+6Ns
fmybrmNwED+yaXBa2Pvupu3lauoDxykYXKiGWwH8uh3428YeofwlKpv2uXthn1XX
eLFNuG1RFgWBhNyXiPN5/7KP8Yy5FqY7VAk2xyL9A0yeVAJ8cQ9day/QgxP+aHUB
J5i0YcX80OGurvXW8g68TJrqIz1NVNiVgmPWDKkSddpi29fWLUWYD6kVzcaAfdbl
Z1j57l2M2U6KY/DBueB19KyUCsPV0cA0+0esFcK44c8CWBFZXmKjKhrZu5MhCELo
/l0kOtNaokqTgocEOZwHrT9pqCsLRnsgvYTmz8OIFqq7SMkMu0rx2eKnklPP6PkO
0f/0dUeD117yy6rJqhR6GJF+8JYwrocHaQUXhEv8hLiQywbKoJRTxMksgCYtBrp6
TCLDUrg4sQS+bx1G1wn9unEWIRQC8XX16ewkh1Xn4BYN66MfVlk8tI+W3lhuA2FC
T6vZ1sHr3tmEvzBD0RqWD/wXJWJH+32/s0o74EIeO5qw9zXV1IzJfBeQ4bxyE8qC
2BFK4hTI/j26FxEptMgUlT598Ne9Pt16L+TjAL8ym6vQ+Zj2wSG/Z5W/CSaaO37J
ZVxbSOdzKSqo1bcYShoiq4/HOQzkfDt2RqEr9czyziycU8lKLMnUAXYI3DMS9Poz
pQy/pBYQSHqubuROotf3eVox1JnCZy44VtihyrQ7Dfrh2CsnEuvYwuf/BEjUvOCf
OL64V7uDhRdUlGi7ACf5t+Gp3ZMuFJ/h9II8vA9zUKlICXhgU+lR4Yqa7QoUPUHr
V3nnfFsHEhLZ/1hDBxoSTbDw+wRRyDFQO0+4VGALKBy0MEY+1vX/ZLVgqSZowJlx
VfnoY+R/H33HAsVBigPp2FlYlK1PHtgcqmfbr2Ynt47+WQlSL4skACA+0HIdw5x2
XjelTTrEkIHXDKGDF8btAldLt/IhCMHhvdJMCjDD8CtmNBSnx5nnFq17FX7OXHas
ufK5oSM6kqBsDp5HD6O3i+stvrT3RLQMr4049YKdxsZdME2hH6zW5TpWMD0hz8B/
y8GPpkF8GRzE9NecxyXjeChlYca6+/z6TG1EEEOKTUTn34RXZVAvi3vWaJibm6/a
oRFTysFQpfZSCbVF533WUupaQaoHA0w/DUR7j3sd2qybChiOOLoRL9pUZlUPt+He
INlP2cwjP/G8iwt295yyE+juUKDi+q60ajdgcujNw+V3ZbEWenQdu00JdyvbBMuz
TtQT5olNITR5CN1R9jK/biiEOCxGCXpIpimessWuI1WqeYyb47Bq8p32NiziRrCY
CbBKl22KopAsEyKpT1XfLhfgPqk4XMxDXa5cAssBsrxO5N8hgxsNYuc0HCzGnf3a
EnVuXgQS6+uKqcdtGLoPO2uJqQ9nKWPe3VtiFhA5RBjNW8fNWw4hieA8/aVxjD8w
dEYUuv0GR7xiu5szE3dlxEg62AxgI5nHzuWX9sfT2OKcJ9v6wMxHe8wTqS+g+8+G
iINRmHiJxbUMEZI6v6eWfIX++aT0+5zbgIdl5ewGaAozaMAiHapCi8+rfm/RRT60
mp9yoVlNwv1dg0PCFS3NLj3PYFDyY0imb06/T28iI2Eqdz2siSRw4d9yjRTuZeS2
4E4cnggkYOCTEkZIfR1prKkPe+OaXQjUyuhCXWsNX/UwrPALeJlFUjpre+Cg4NlJ
V0z0sOuA7n/DRrEqPCY5ina6dAwpONviaX4zqKD1i0bozw7PlOofr6TnfSRP3lYk
FfGrmmvd+od7wFRQGPEtIN9X9syODgRcYa3U+McsK3rPLZNRXsqB/GD4mb42Uvww
UL99fj+P+aje7yyROmhRnGu3H4RlGl6CvXo7XpvzJqtAyhj+hJfuA4dk1lIbaz/T
7s54wE6eOZTMh8QK3ilNT1o5ut/iYueGCg5NLaqMmyiajmzIOOOMzyim9nrIzTS4
Lmlsd339UvsEHM4u/E1mY6lF6bXltJDgGwKDibe1P4PAEbCKhcvSKUapawAviqF6
0W4tlf4aFNsEGOrzMxxaQsgSqBHBEe/5Tv45I6mzBMNS0seij/12jCJ01MhUG0Lk
Z9uCB1TGKHoy/CQkJKxX73SURHZI0JWUr9vBr4qysYYLFm5rbuQI2J1vfWbEwaNO
OmUBr/dB831GTejoIk2YL6RZkYaXwUdb+3PyhHBHGsIZwrXPIYwESBmRDRgmY0+X
QfCdiULAbGy8Tk3hDj8a0RaM0MUmwMnLjRr0xAUvPhO0kV5rwWq3mDhYLvF4xgTK
5N9d1uTwvfdlCgBCZkq0+gUFf17e4/kQ+qd3KoBTP9/WfkSAHvGlDaj1dWjli7P6
fShwef7VJHgKlnR6xoDA21XLWsQAT/k3gtwkYdRi9jtmgKdXLMaHK/5vX1pHC7DR
0JvNC+s7eRpRbVtCvnjVDysCgNSr0+4BKW44xMbXbDBAFgc0GWEnR3lBPJZBfxsv
uZWm2TwnesAl2Yq1GHacNmc59jyK/e59cU+xeb4+aGIinJZGm0CsBxkaBr5tOfw0
ZjHvgpn9VdBXpVfK40Hpr2FvqL/kziBFFRCMzkmmA8d5otzaB5w9V++GZLXeooDa
MAGP5Zz8M7/Lb75KUX6lc30avlQBbkp97q4e8XNS09t+5Xd8TFl6nQIKJZnQujwb
wFELAEmPihoQ8vEf1OH1Uq5SaHxV2GFT9HCwDMcb3fLBV79E3QdOVxxClRGvgbtG
nw2cqoV5NdmIh0ln/hmpWHNCYsFfrmX9Q5iQ+i931CsHDOZjtga+r8nokEPZu81d
P4O+GsC+zOaHjjYBCcUqGKtGx4UIGTUf2qiZGsbUPR71myu2HrtllCGBJgodplMF
fqvLZkCejHQyfiETzcxbFOsNNqDe457IkQsCe5i8PjU7rAUklORA+zA66LcYb1PA
0PfvjfKWFBxtoNEv0w93UMVSr+jThaJEwbVuOT61c54rxjcbu0KrCbxfxT0qzU4T
Tuhz0tra64j0ToXCIft/VU+V2QMSWd9CzRQkvVcNV28OWRebYFcFDe/j7Nmer1+k
djVyuZbIj91VOptfGN6gV4qOa9cOYYHt1IPljL1CQMmQsSl6eMBZYs/lBefq7Z+R
EvVpzLpkBNgad47vZzJHX0Qt7rWDlpAvCg+tU0K/l3weTy8EDv41wvqPR3+Ipusm
E6Z871IZ+9/aBrLuVc+E+W7+FhUbDxW9jk0BKOdrd2nkvF1sv68fL7lWa1fycWjO
yzOSj5cVfir1ni/4OndwiZR5b40a6s7dG16jt9nXjGvGAwR9g3/vvtD9gM95lVyo
Vnx4W/kVK4uICHKQauNZT9yW+ivBMBg6EJh027Bija49WTC7rFBDBQzZn2gC6p0v
/nmi/Jd3RPJmdM1S6wuotfZc2TTRCkKnNmiO6svDvYGGYEbjISRPwJldVo7vASVV
EKIiy9n/TeP5j5Hx6Nl2oiEvb2mhpctJLK6PMTqJ+qf80sbVJnJomgiJxCfHjhHS
AjyY+qkcE/gFSIly8MGHjacyXFt8bO7XxYKufnpKOL6qc+l5DikPEJQCGuwuf+8o
K1/NgZ81X3IJxJ2xnvFV8c0Q0DypPOHI5jw60Vh/NROwJOSxDfL78U4cekUBaihb
S2WVMJz+4eTV89O70NAiwckV6ryFJgv99hpM8CXulFvJmg2yWgEHqQNa75EeYp0c
+2DZ5CKBDZinSeD2X72QS4fEmOQ5VAt0/R6JN8d+QUTrBFcmhUE+3BA+nTZM1AgP
h+VwnJaLGTXa5bd6rkGDOQFnk3GGtVwyQjPX5Hirqq3d2tAAWV73NfO0UXcBZdIX
y1WE+7Z3oZbhv55yjniNnSDZ3HBwBax68WV2J/n+ezbkwXP2TKh4QqLuJ8in/d9e
d/ZKjwKkOXX8svUh8XVznfULNYG/BabU/nFjayjwh1Fw7+2uvHSSj0Gcwb7ej9vk
KOcRKHTkkFyIWJZjROc8AU/KPDz9wRlgrWLG2NR7BPrThCv5VV9d5OfT7mR/cyv/
2QESfTez+rF6LxKqtt+WgDRf0isxhNybccnJZXN2BOCiUWwKzh/5nYM/wxJCuRC+
GIJ/r0iaueFMfSgFH/AkMn5N1Zo0Mzxts59cwRxhWnLLLaXxSDdsG2Jl7e0Och7u
20TBKGc1nULp6+tG8R/olExLAk7jm1VdOH70VJPOYshu3sdUU8RmXw3eDCa+lpBL
V+wGjm9TbZQL6cknpX2BwraCq1o05QatUR2RfbgcxuHIowaC5eptSjlJpdky7gNy
8zyVq/csR95ZQUKtrW5hKly9LDspnmAyAXmC9VzKUfJSdHK0ng88eRUjm0IJVtcM
Qw4k4jXi4Cxio0ZWwquN2kNR2FFM6VTTcXo6QS+kATJunnZFJaSiNiL2G4dh1eBb
ZEI9+6WWe+0vchpBp7sz5jJBVBHXPpFncgWP6tN0BWSAGAio/n/LI+CdjleaCoNI
hrLeBW+sDG/CNqM92jQbyOZKrZO8Jqrqbl1nWRpbUkjTc6SgqAXw0KOmiJGMpqQN
iPjavf2oLRDDtTa9cE7L2u0HrjhlAOOZOzKm9aiF99sBbuVwIVOIQUoIkTM2KYXH
9oivHcRffzGKai8dw8JLhYzWXM1iD49JtUt+f6+i7DhXFPrp+SxkRGTHhafRWTrQ
lTFv8gzMnf2eL5AYo1XpPgxR+q6LyEW+unD2tCAkGc+N9rruQZ0B8Jj5AtetXJTv
nW1HISzIe2zEvYE/be5nIwVQC0/S9j3F5/PsYcLAT4G5Tfnje7rKK7bWdm20hz7U
2T3BNCxijoL5LdNmMWTWrEj5QT+w0yyKv/OMGneGeLe4809IMBDetVMxmjYtUC/M
d85FTJoHk/lkJ23gYBki2F0+5JhsUaXwzO38mDxYo19rDMIHIh/V+uS2DHhWZPGa
0ZwqsrkUnHpzKoohTXY9JeFBG0qtNS1OyTsmEc+B2VUgIvPQ1kv8qs3vSrCJgmlT
F0J1B5QBC+9K9lbDP/CKmr0zSla/B5d0Py9Y1Ok4OnDBOFpqIvGJ6gzLNgpetQC0
askzGpKq24AhfbUOWlFSrzA1EaV//5XF2SO1ug9ja+VhF8i8dAML0FHfzb6swiYg
il2xlDpfLNTwRLwlSrfV801CJhyYIGd+7sMdZoh1fgdFp+yGQVt65U4kdTALiQJ4
+dVRN0pBAPvdGMkH+aRC0fD4/YinP6mzUL2By+fqfteeY5P0HPYaZ8Z/m9IkkJit
otz9sJsSHsfJHR8GH3sMnt+IK8gTbA/RqyjdH+etzMHJfWKKoYT5zkbVSaZFHbNf
TQ3u2HKY37oUFiAwFhFp/lYlS6oXJg0QwHLXKWn1tqgTfg0TSh6gAPgBZn6hDYLJ
ugyzne/HWAGFpU7o8rQAKdk3Sv/5MGq5eJ4RiUfBMyp2HkqKZawL3RzZvbSA7QwW
k1n56V0gtcWK8QjtHLxlKoxWWWvyrb8/fL09MWjhHyo4jR5toAO73O/yC3KqIpXg
iubVScODjzJ0I4bF3tgWRGhHGkLBZWeowS3b12caNYf/2etHXxHCXXjVMOEHfdEV
9AQvg/wdGVjW9lG0bD2U07zFquqsTokV4S15AllX6EOaCGwZ5ILUPHD9tbwT6xlU
B0Y8Cv9GLVx4fOQsy7CnnlNXYAkeVsp3fvrS+Dp7q8UxamEegDAZ7E4Hjnm/m4FV
a5Jc0j/lbRTAL6uAwfSRpTVuFAjo4S/mtmRCCU8BZbxT6HuyPjcG5ACCnLiXsdQ7
vNCB9KIVTLhBnzkNrbzYYXUa9tVPWsu0hzblYqJItfCItWV3T5inxu8gZAuOzX0x
KVPuONE9KDaj0l+qdp+s/QnTlwUFE3G2jvlEx2AzX1YbifW8IkNVMiADZzaoMDVH
+w9DDW4qw4jNm+ohpB2uX016QkijubudbR9KGedTeeqV9UxShTHXOR1ykZVySWf8
DA1YmdhkhYTnTQaNUT5TPGQDO1Aq3KJpVrDVHIh4HK5S1ukR82dEljVn5aws8rv6
dG05ji+suPEd997IGH4CfO1UfucSBnOEOjOEF+zOevhJMuvGpO6qf+eAifD1i/Xt
4HKme0NDwkjmwaNzW2fORAMG1q/wENzFYO+zzwOuizLVqucIu+rmvCeRbrGGM7Bb
z+IWfCqAS4hCu6vdz8CGHpgDeiV6dvfbRpCGsJ5zLS9ap0pQMwsEBSMt/zSveR1w
LpJFbbpJ1g135LbNmLoe1WYi8AS7GNWkYJSRTk35BmIOVkECci1ZClep4OgCHGSa
lcyJIavN5hcy4N0Dos0wWu8TFwbv8/f7p9jSnWLM9ujsIwKXC173ZJ8R936xl+OH
ywySAlx9wctRIEBJ1xf9NKUagKfGf+RPe7z2YEzYlUULgCyrLBNyHcBosUQTAyiZ
Dkv7ckXGX+7OrjJ2GpPM/w44WGbi4kKjPLzgCN/t6t6mU1sCcY9HtYW6PJIF4k+T
o527SVHqldA1BKL4foa+neRroZJFLe9cIAxCjWkXtyUXFpvNqfhh/hzumtVa5NQH
Leq9YI7T6bqVxlhwqKMWPIJyx7Kr8vcuSYRgoawGzvhAwESGQPyMoUoIBn7oGQoW
osQ8HKOOqd9vfMyVjlQaD57CAiAroQXY372MC0n9aOd4rDl2XHZrJTPCqIwM62pj
OZ4aFZ0iHA4vFt+dpLW3h1HwRclnCIx9yy47/or+Qd9kCphuwd+9LacxBq/0q18h
Wbo7HFYwLS+KHrYplcLYx/JTMAXz4LcGv9uUwS8RxtuCgj9sPrcNBLoTSB5/WqUE
bqsrZ45H+9mOyIH17ppe+E4XAnw03N0KxZOnw0xJqzN5H2vyuABYJgdJUJHbi4xt
tqd7kUfxHaz9vF4sAb0RS00Mf4F8FNAgLIgrYsZzipVmG6m9WPA6XWlRC7jZThJK
yd8/me7OaUgvAnkUrDlEUjtVNAeCg/KQZzgpWBBOMwwLsVjOEnk5GwzNxgn0jHpP
k5IgwqbPyq0rvo/aTO9/aVIVjJG/A4of5l+Yh9I9GP6IxQKnyOC/QX7E1Ud4b+l9
zg5m9iTDilObLjv9fiSkCDGTi8F8pgXrnPf6Ud4v8gHd/OnGMsOWcZzvbmGrWL+I
VQnpci4f/JXYp5ALi63guCgn9Gxh70BzdGrlC572FYOqTxEeb5Y/4ALqGUQWpyHm
mHmFE+bKi/orGnDMMpagP6c+IRuE6hm6bU2ucZw1BMGU+mz/sjsi2eHao8AcSDbN
8Ul2xz1o4q9AT5U5iR3deFfBgrgcHecMwFTp2XL5mll0uTfCqMXX8I5lhoOaPrPb
AIolSyXfZa0lHNb4WvC/twSGBWtOJmQiY/FR0o/zRhXCMjpcqZ2CE/4aEv4Igi3W
NFIrHt53lmP1BE+SvnPDYTo254Wz2DEl1oaCEBzkDqBY3U1CJF7p4wrGkP0kZWMT
ndOEsSH2HlPi2nnID9kqfYaKA5OWWxvUA5faq7BSiDRai59/Gotqbk2eAk4ZIXO9
/hULrA94LAasjeyLLaqXk4jVjHuYbIyDrs2p5kccey9K0zWcBAohTbEUkIQzKZxQ
hgyq7FYcuXFTmOxbk3QwdAYjo6znk5n7gkdG3BDR3Q2WpdOCaD10NuapGf7B+DMg
GZRADazpqvgmwbbUVT4Xv66ZXABRC1diGjxeUUZXfLiZgum1xqjjwc+YkboORLdm
ECBSDWfieK5+uW8yZHpBwQNfUSovdxdMMJCMQQDB54JMUiu0BEfCzyWvoyTsVybk
w6ujBOKyqHUj8B4BQiaSyFpxIcouJBDntLGSZ8/U4CtLsDPs4anLPiE+WbWs5lJD
qYzKAsoyHH7sgY4Ddhx73Chcd4/Ya6rWkTFMJs684++Ed1M+coB3nXiBf8P6IXa/
4xUUAp+hcHTZ2N4DRt1f0iozJ9RBeoIy8W38x/7OjR1rQO0mh+/8gDxu52eIwHAt
HalFon3ZCZScxTD+0sNXUCtRl3YM7eYzhH9HdoAz40PHfDI4UehSBJ5wa2uvbLFU
EysTPYVZBjxUNk7DUqSS/6z7/htzugwHdkvWtIAM1O2ktQa2QjfMy3sPNh7VDqme
WEXrwJPMMp0oTRlRF+71WoAFRL3oYcGhoFuwVP9hm0vpV/Hfs+MLWMUf/xrr29Yq
fspqXjzrlfj9VMTEC4u/8JkfP9ANavRl4ss3DQtW/uAl6gvc8LUodZ2pAEujxmHm
72pFh2scPalYfYGKD/9rIXJYTihDVasCAP9gyWwnh6aU+Dh6i+simyVauwHR8MR6
ItuYfSM7VeJg2xNjONVUHFnxyQ1BZalrpuF4KQeLescxDrNl2w1j5yckmGW61GIg
Mk18KInqW9JhWunFgznfzwJENOyFuLeJ2U8rh6JUbBK6EuRLqftcCtVszQdPw3Yb
HXNXtzOMy/QVDaldD1eFbAcRUiLxQDsGFXK5ZTe8u4Tv0hsKXSA7r5X7for+Vlav
RotouJzDNzJfMX7U95r/dwEX3kiFO716sjis2LWFyTCxW5fWPjLd1vQIer+py3e0
7P1/QDEFg9Wolpz0IAiL0Qe5n28OWXAo3nKs8L9J2IF/B7pycZ3gFLBnx63Alqyr
EMdg+TwPbwDhUrCJowWh9IAWYLDYSKsmNIvz+tY9YYdpOdqcO1MbybmD5P8z0X5p
BGkiQDIbytBhmfFsn5wSIZJWM7Q8L5AkUULxcvg+zeKLig+xK73xqO0PsgeCBxwg
1fzVjKjva+YON/SYpGkti4iox6W8tWGBsmoNzoX3bUFkL6GZd1XNxq2CkYuE6wxN
GmzaVdjf/K7KNNHb6rrY6/vh+V/FmShllNh780phbvd0Tgr1MOHwAXTa4TsxfWl1
LMSP4KODqPeQEYcZIl+j6scxyHA5Lay1dOag2uifzbY57ENGBfwfNSbQgtSCNCas
/UD1bCUuBN95eg4XWeB3XmeM+rMT91OX3jJQZFjtPyu0zzsBwRSndL34jzOLYwVJ
BH1BfBUNuqecTj993bU9Z4w4tjqmJtGIA/x0L7hEqKBpmVph5VOC2pNHdgT/QP4W
KwWtkI8JYu6It171MQI1vnOHrvH6psPQK2yHSNcpBaIyUlaUagiKlGwg2RHEscTN
S6yzlwD63EQhGpAfZMh5gR69VypG/3VHQFmiN3cAbth0BofZran/zWzAV6qULKsg
UTmMD90btPtJJxgZhWwLkF3XQ9hDHJuJV30Ng6qZNcZquNGESVHdeQ34BpOQXVEM
KJ7X8ZINFbrrhwvnztbtv8LwgJ8MornkudDSQ8XYxuju4g8LCDnDEHdy4awM+xqw
sOqA8TDc5tlYIRASLutdEtpUxECiTfgSWh2OzdUQzFOswCgtXTb7C9EUdkAJW85h
PpcE2fwN9uBberby9RhohSHtt9CNJtKkSHbURu+mite3BsQDKgmKMy9iRdqA1eax
MCNpxUB9kGIOZEo9qEoNgZHmuYCuG4Df0VVHSeG+D7X0UPAReUh5AbzaVeWd2E6m
x/2RJA7JI/iZ2o2rnHDiGZl4qTnv9/eORsENFOWnkKfrF7wUlk0MMqrVrUD/F+nj
fXS2iSMvwLOwoLVQCeBnQ4pjPgI9rMHNOKlnlXo8qFIaHrrXQ/hsBDwEil6AtIIr
LHvhPUWY/QkhjHm/cuzk/naMrlZDb1EmtD94nVoYCRurHk05HLvi/PhqrTbr1JMB
FrY5AM83VXINSTAJBoYGVF1DUi8mU8xNzryd6Ef/ZCckLPg7FiebOngljjlghCUD
SgJSOJ0lokfbpiyF/bG56S6APE1lAmAOsceYvFDVeVu61IHDPeU3G7lqFIbmhRW4
bPdMtK2ee8uczvQACpkJqLD+r6O53wqkqHOnZmvjMJfaacMDhLf78cpM70zya4LP
uOnaKC+wVJs8ME/FRa0UCZnY9KIMxJRcNJukeRjOts8JkIVXyuuYMiWb9519G7D5
HynWv46Q9Z1yYbvw6yj62eAo03kmkRzPLXZr4nIWeHqt36V9r+ow4Cm4c+GtldTe
l4Wm9pex758IAJjf0Mf2laY4jm+LQtqateUt59dzCUzXueykCt4v11Uvz+QQaZ4z
/mf7PCAZrLhhV0WMI0A13bftdOY2xRw6WXSDJpVxZ7/+W2p3+B3ebUb58j9gDvij
s2LH73lRBQjgbNGoCF72F6Qoa3Pv96+fYaTDWlhb8twmuP4h7KDpqz6R5iTL/lWx
QndtqQajF1tTKO0iRpQEf8JaXYJcmhB9FcYO873SV0pDJ+NvppQraDziKHf3qnSp
/A9EsCvwI7XguyP4oul15Ifyj45m5n1hhEYtsqjWaZXa7z5IUjW0+0iNVKAQr1MA
szAmCi6m1jhqT5oskNMMax8ws2piTjzeg39yzfzmeJEuhqL17yevUBFAFgnwrrDj
j5U04jSdao6hQVLWxBRKmL8bv5PdFFgKlBOTCnIDacIg2Ld0dpgtZeZP5mfKLygU
jjNfKiB9R2zF4nNtB1JTY0hA6YJmBW3cKa6LsAOZGHARUMY+vJVHf5xSKzBj1FUP
KkSyt/Elva8nDfaaUvUKhl7H3DhRyiU0EskQtZrzpf4HaX+1En4RkYQTjYPxugE/
ueorj5V2nY+DFQT1bzzN9ito4f3oH731IxD9boorGVZa9nRGFuFK2hVFEEZbmBzw
sp0KWXsO7XdmuD5MH7+hqHzOwQ+J6QTANDQOnDflv1aSCXS21kXJ22fci6HbwtFy
k21D0FC1dxkdFxZ/swh9UG5aPAp2pfKepSdCfbI781m6MmUYkLPovB0cIQSizEZG
nBy+B8pgk7FAPm87MLtExKYogCGh2IQsPReWDetfDHfdrB0GBIgY/QDMbs/8dwor
YRggwNb6F4oMKA//agNfrW2RywJdUtdTrCy2YoWeg439uf01973cSisqeAEdLNu5
NZJHGogYuxy0epGmrwtUz/cAW4BFtGdrDpCp7AlBT/TY8f6pgIVSw9VrZl1arIM7
e6bO2x/JipPlqYjESDicYmX/Bv1hopu8G4lWyZoPzwuDnBQz2LgplQJ4J2jjqWNi
U3VFJdFu0uIpy82t4BwDSjJ9WvymhFQMfSULaZlA7njJXrSjatBZ7zSjS2R0SXIc
at4xAD/wYmEUgTOMO5ZYsehw9ufStQ3Sl7cJt/T9ga8OeUXkjNnwS5ulj5YFGJG4
ND+vWgg3eWon6y3AyWrIbNcWkriqt+1KL5jydQLHGpxJ1vMlXxOTvlSi19cIcVuy
TwIPvqC8oXC4nOOi7Oal01kQNoihdsaHK1u+grqI68GCJ8oRipQiGeHVnMFNCb9C
eGt/pv/H5grl1KcDvw4pAYxM8nMFc3Pmag7+O72+MtCUntsrTLy1Z5BeAJqh7ppv
m0wgUGqdEGQzePI4eTZzIwZ8cgc30ipY5r/i6WvcB83azEM1nn7e+O9hH/6MNxbJ
xm2TEJNzGGmaRLk7V7s3Qu0aS8ZLgS8OBsEiQCGNETJyiMiRih+72Yc4l1m6Ot7t
fGA9SODmZC8vOmGdwiCp3Y6t23+Hb+dYWYdLof0uZ4+SSaCCcRvT0EeEcarqthcG
KZDUCrBcdAwnH9oh8s5iONjghf8PDViXk73w2KJbQ+4u6gmlfkVocb4IdjLuNz/w
oQ/7//g9leE0/8CkIi6NRYcTxEvpXP/+rPtlkC2r9h8P1iftyx+RzsA2BQtmdgaE
ZJvXThoy+yhqsCM5t10NvDr6xoTEaVPUP0lLtNP/Kxl0feQDHgpSJZyItYq5mBGA
HU7nnr1TnKIWYRgWvkyvNENYtb47RBozCX10QXcSABg5oBqm2szgR4fyVhb27lFv
ZNQOsuuYh65hpi5RkkX27j5eP57vPoK6SCaiYthT5cKmvLIS8CE6+5QoOjwvKfMa
BoHb+uS3UekvPiAw+Kl63qQn9RsmNg+Hmu2cTNjTY12KRsRUIlRghRkQC6+H0awe
670Lunb908TP6byp7iZTI8u5ad85DuvXVYNLegIEBUnyC3PKPmYAgkUxgX0VtDbT
ok8BmYuIlRujumUvLdx3Aj/MHQvFmeMuqL7t8PCN2ciQGOVmONx56FLlOAhKa+LT
sG1IHmZSIqeNvqY7JSKqHryLiUNTWrnYWdU6yJHBkO2OKbQ5nUloZqYnfIFRgvwf
xQ9PYrbRMJAuM4Obn26dABsVfW20dmPO0IS8XcY7e+md9wnsMmm9LOze4V49GWdF
qSXciEkTbJV3zSDSbVckp4m2xAYtdRrXQNyIaxZ5llkqYlMGxRTLkGudvXTCm7pg
xluZ2g8mBPfz+th1KeLpEdYhmejiX6DE/rxzBu0EC/dh7GW3y8Gjd8u9s33E9zY4
qnafbARNaHBu+4FbEnCSWs5plY70THRZHCf8iGQgN8SA40AIKy+nUIQ5VsbCGOMv
4PkJD4q+ve7nC3SrWYfFL/Q1RcT85cdQjBsSqjD+NxcueFn3P3u7E13qV2uusFUU
c9AMGfO9u1oZHWuQGom2/P/sCIP5mZFu2LFRLtFb5+rnEGO2nHdDpsS5XeRGKZzj
tv4Zu+cZfnlE+KFj7/6LkTAa19aW/0jtzDv8U3P3PWsMgU9Jsh4uI/ikAZkQ4Ng3
GJ0jfSKGnc+Xz4CFFiJFX4lyRHvI13j1U0W6a2RoXIlg+7W6JzCVZAmRVcZ5GpN5
cRxm6Lu2BrBC06wF7/kWwuWVRRlefCaRTgxYDxWVr1lhvUhMnUIZER2cYmpeFuC+
R8xfzLYF09hKAvL7SsaUannBqy9ki127/OAslCajscO9W7YqrCszi9XS/9fTREgW
OHYWM/XfEWkXEtLMDv3ZBnvanU3cUR4LcPdweeyM74KzjXB/FS+Rpk4wSVkAD7aW
1UejkThaKzRjL8FftwSNeXOxVSBk8FZh8/QkRpQ+yhGFzDthzXASRTrkmH7CfrIH
hpeBn4xqfdPPUhvdQYqNK7+RAh9M3Tjkc5tjy6O2KYf46tkuFJ++sMwzSsvP5Aky
OOGOL9/6Kt1m1Ueopt8VJ35czjL2BxJplEUhpwtgniCcMrcqg6rVPm5wZIKcuqGH
DuDoh1HzU8tqOJO8uV4DOkVZa8oLjD9cF/Qvor3dfpGx1tWBhVIPBhJCNr6KfaRS
gybNSwUcziH5es4BM1gFH9NBuVgEjyTmUOhQsME3LZQuvSb1D9z6nm84gelU0kwu
WcZ+BTZM60CYdAksn6dRufLI3fQRmpFhyeX8rtCXnxb2dzMEwDCuQcJnXoBArucH
o9BxwwTl2H/r+LjxGCHhB2xJFaD+dAdnDXMMoaMN43NWMG+n9N3Q5aXH3jGE/lAc
XXAtnW7APr/VDK1Am+o5RbPsVa2BpiDmJpi3cg297CIMhOI6UuE7j+eO1tHQrAFx
XGRUj1vFSIfHdymKvXPd32TbVsBd/RvpCxu/u0XRlnJo7eDMsR2Mtnf9lMxshLXK
St3IGX0HljWSNMNL6pj7p+yUUEeDcrqorP4w07DoewJkiAZpustTcyjFMuBqOmeI
7tgDPEtdbDkrMpM3Pjqw0KvO4i5LA0vYBWpwomm4usGMrgSQMUrJxLzEKb+AIJyp
YzdjefppcyeDhiGZyDSHt/Tpth41QGr1/qKeu1PGfiYdjebUOGraUUCt45FiKEaz
XnATURw7lxsFQ9z6UsM8aPP+qCvKMnAUMU4krMo/21O2lZSJVbEj4TZdawDYo3qR
JzZvDXkM41BOJDZI9JQvwZXEHJaBH14hEFd2z5CRwb7POuf5gq432K026kYT+Qd3
SJgw/lZbb2D7OzFMzB8IkY6/KLXOavDH6S6IClFF1g45yqgZU4r8uQAZN5nipTG6
AghOkPiFo9kePPzUaAyZpOggKJX05A8Wvvk7gMTI+f5GNOThBojc5yH//sWHY4+T
O19uHy859gyLN60n2Knu5YGwuY5D3VejRI8GBxdP3M2AwiCHvOvzqInH9ZaiAWBW
anx1wXGWSl3FfbP71QVhbEEBqT7CiRiUyQfVwqhCRwK3ej3CzinIWgLhRUC++m0q
+wBjxyg6yJ/klMe5FZyhjj5GlrjAgX3rTMXY7WJCujatL1B6jDckHe6gdVTgkXxx
oQViYbbUwt8bTqt6OShjmDWbB4L2Wwr073ehmuzMW8QWLVHchFXX3AuJSAEDadWd
s/AMRuTX2/mpn9ZntGDQTfFqeYlSV+E8JKCWnxk0o+HMSfF7gnostLP6LpTh66dE
F5Xwxw+IfzYj15Olpsv/IfcyA+L9RBDjNgcmDS3dNF6gpv08vZ5TtDt4qdMdRoZA
1Qgi9vSxZcrRAezgvHs1nCiAaqrqgmgwuNquC0Or5Ybzt/dQ75KYYuee2m/WZZwm
1BNPzqzW+Z7oIp6hH4gDoT1FJosF5bh3Q+jwS9Q/Je1puokiS88HtBwrOvVSsD4v
7SyPsMxO+WPNy94Xn5dSaDrq2yHL4CYnf2uZcrJCZ8gLhD/XShsU0CDo+rC4Wq4w
jDoJYR5JHHeuOKO2MCXKjaqBMwHq1LITwKivGWkEi1Ui2nLLJQK0I5p8Pm/3QIb+
xS2v+HpR0LyEnJmUlbT1wI8wZNB9mEiDBTOJyFuNC0Hz2GA/l0VB0BZt2vWaRh2L
1dJyQ1kulj39TuGxi2tMdfMZ90D0rdb6vLDuY3OYLAy5s5sOPjDmOkw6ODwS8nY3
JubXDWbpQ77WNO5w64sc/Ukgm4RROLaLB5JNFOF88IZZwA5JZrkUlvtwaULcjAQ9
tNBiftpM+Tp6Z3asYj6q06VidUoy5jwrkP+7TFQQFUMvPaLBkXJcJdvpuAKp2iBz
mODROg4WWJZm7t1PorEefAflmWo9tFWp6HghAjXL647gi+TubGhLzf4Ko5xLpV9P
VyUziJa/YXYaibmkhP4aTrTi3slWDZKz9FmdTjl86AapIytcgNm3OlyN0grtNS8h
Xjhu3bNJ8drLNgJYPbrbbC7cR4loXj23xZd66ItZcrMe3gMIbR+G/BSDVcIFx+cc
rcUbun8ZBNE6vbL3z9xJbSflur0PlIuIp6kCI+Evc0t3IYdKORK+UBkgsyTc6KON
+f4uicU2u6XdQXgnydm9+Ot/fZtvKTSV6VBBqN2Cw5gO0ow0AJEB7J9SZ8h4xndn
UT4F/xFTq9Ffy5uDCvREs0790h3uMg2GmLEmEfqCpf+gscYYR6jrz+ENjuTPb1ug
kAUAu68HclnAbenpmcjXMcwsvgKeuj7U9bvo14qfVONpcx+55eCorbRSiPUmDQLU
PswUhjvfWeOC0l2epER8JZ5eGMtXMyNZ4ZuO0e7k18qsQtfrUWlFMsEoqEAjEF10
+79UFiFxSkOHN1b51pNQrU0aEQ52rxnlPuooySvWYBKWyu6NJWJlK0rJaveQubdo
pzEu1evUH5LYJ/xzPVHZUYWUrRy+MKAPYb7SZolqTDoNr1puqNSQP3oCNEaS3+h1
FjtZ2SG/HvgdUw+u9Zt3kVNCq83BsJjKt8rLq6sK0r6fAiTnCv4ICQdZx7wQxfxI
n7DWJhfts/jXQ2JXaR213SLk3Hz0Xl66bdo3dt7fYfFUdV24PUkm+/DyWu5sCMZc
rn5noDxjB1FIqPC4d80TRzwLDdx7DtQa0j9eCrixFUZVMhMidKJHQbfSi5WEO0G+
6Y4KzC4V0qjrC9TAPz+Ssk6wbhz2MJL+JRxcejqC5u02vwGx60SecrQUOij0taex
U9I5oxacj/hTID3yeUeatdqex9kDtxYgB48ngx4xHTRLx9Zns+mo1Ygrw4EkKpYG
dxEfcaEW2iBzTlH9CSs5wBnRp+ZBUPGOEZCzkIxK8ewZSRIjt+LL1MnjYmR+gDAx
YC0mRkZaAN0LYbD1insVVo1fsTRzUlNesgjdc8Qtyc4pNanFLAbbFPY7xgAyG1p5
0FJJZzdh5Zt6Z8rjJ5EfxUf+RpPzGn1zn/4cOv69+yPnECxMpvYs1MCLcXRDRxkE
34kpJnd32FeoUe4bAFKe/yzIKGudKfK5kfUFQ0B6XCxRl77XWaM8wOD7UsMcnpnD
m+tgM2p6SVY7cD2O+6y2Df0vraLwPc4FBzE84ZBbRvmcxT8p8X7gEnBWxRDVNy/x
L88Jzow9Mjm+uLJTtYTQZ7dQoi/HB/osFWK9JTaNuxEjoWXxAsC0Oez2upbR0cFT
wjL+C5eYHfwM9QEpXkYCgSCxJ5aJsqwEOPGnTzb6+UJ1QBsGa9bIdKHXlLkbptVb
iMEQEa57NsCbJN4BMuIYOky0Qr0/BQKp2p9hHb23CnwZjxgSsN22qtYCkHgWVQmh
67eXzVeogOYrgMjx0r5DzQOb7O02WCO77IkujqPtmGBMIrm64PMi9Q0apfZgsAoJ
BehT37CjTmGUDcTZIOzmJcXGeqXUW7uXnX2vGRtbkYmCHy1X1geRM+lifCxK8AbS
r6n+KvJS+ZSA3kH/RI2XUs3sk9E0KXOtRZRX+ZHR/P9QDfGg7fadiqLfQAKtIDxP
ZI33i/xB2TYRj7ZjCesm1ecN/1BErl80bG+atSRDTAF7hEmPpJRVmKLa4tffRV7d
bd6CyYrKivwE4Iv+L6DZYSz3FPB3MxCUfttnmm/BNQbeTgbA7yG80eNHynzB8Gln
XKXBoidYl51jv5YN2d4yMH6b9zOe7UfQVELnmWUzVvzXfFygXLbjEH6LMmgvGQMF
JKNmT9ZwREYdya4DAIDEuzuI9lm+4IDNTGasDob/QyvrEvQXxr1et3R7hKeRrXXW
zaQ4GdFUN6mmKTOptXC7AGKmhUfdrqpHqYn66VbkugdvuUEdBlr9ZnQODxksRdm8
jwBY2EvWUKh1I5DRcDfQrIL/KhP0g1nFh+uuYDi6zllY9p9GTRjhmN6s96qnuIlJ
bmJFTldM/vcaYxq8IEvjty9rp5ZOBXfRw87OMnaqbPAACJlpDhLqpvKc6gPzYBuL
81GwNLOMC6vyvhJSRVHi4uqn8Tor+B2rTrdyxcajvthjLvzk4+RiUHln6dXaSF3r
lrWtyHXpuNdcQstwQ7F2j8O/qe28aa2vR7PtYVAXKeOyxQuPBbaj+bb03eHRaGgh
NmKIK8IflC6PWAu/MovrlHavhtAbB4Hw3OZcQB/cCmR3tT2wiujItxpLmfcicIGA
o2YSQgghavluBaEaT82kFfFoIaZpBVrFx7iDFrtlzZRcJb9N0oF2gW7xjsbn+MMq
0gvO1MkMLKo/yejyGWzfwkx3olBQhG5XZ5h8OPLwnBpNf9oSy/LnyclTPpWfp6N8
vv/AbOyszlDB1/sbDlKpMXg6lqoA82B1nVJ/DYIeBOhiGUuRCQrq6WA8Yxce4oOd
CFBlpDTZk+kvFmwciRZhe2fKDReFsOKGHfqSZYkiJVzurCbdNzSRBwGHjogY6IUP
7HjTixm90YY5RQhhwKHAKMefGhqOYWs7/xLm5gtRcw+X5zEqpKFJHEBUyCQyMZKi
17T/18bfRsByIjiLJQjNGToh5NzP7u8QRHiCalt8oMb6n2WENCCTunK1ZU/UWtx6
yotW/JKjstbXuG6F1cYux6/xshtfzyoSfv8ACce9k4sGpDxEehHIS8X1cAZRkVLU
LOISEvrwS129JMEr4xqacBuqx+FI6V6y9EMV7Kx2Qo/98mtNklsyvNmCUTAVAbXK
+hjBC87/Hytkjq/9hF8oBaT27u13weedFjh7GA43NiIq6lfEVAkrotE5febSYb5E
8uOzNP8x7RFh+0c2oh9dByRtPWLhfr54zPV1k712R1o4vqM3mbtQwAmUXVM/wzxu
Uv0U6V3FWK0TrlFBSlzWIQK1l2EWCJwu2k0t7RddRB0f4AfO/GPUkBs/ex/qGeo6
+oLklAdmnphww2rP86qsrSQCWdGpZyo7zCA8/etnD6/qcN26/dHHRxN1bnRiObRX
F4OuRdKXRmSHYr4oSCkdLOVSf9PruyyR/lvSbCLPcCdTn6fn6q+FFhlN0Hw8YWXL
Y9iS+eB0OXvTFnHS4lmaV3NsTqv3CeSYij6IFnlpIrol5LCEHUaSQEY4n4ywaZs5
UJ1RcfZdpdDaTfQPCaJcqCLG9FVbityezEmwZaSfUZdMkVHm6Tce2/CVVFogLCa2
OjH+NldqWfXffjEB3ob/UpavZNG2BS/0vKWeVOdoGg35ZVot9azVHIFUlXyFCTBm
fdjQjpdfsN0IsbYMCGlyqCe9uCwzv3+KAOXhSOMHPbZm6/E3JILjvkc9UlWErvFu
OBRGIrAFYhVnYCIUmKuS537Os5cUbKTlnpSsdZMWXJgxcDxQLWLPsJbDXADIDAnE
Dud1B8obxJ+Nwt3WWrRvrSdvMLzhk2fxCGasTPbxhLMfYe7fQctALgDNylVi7Pvx
LFIj/+67UfhaE7JrYS4F48g99qopE06oTb3tR5N1+4FmJl1AuZZ1IxjVm3UmLi8q
D3LQqtwr7P2l5Y5wZtlsRRQr3BddRNfez/BtsIfjQ4PjiO2mIznEvc6aZi2Jk6k9
7tlcmBIYRB81IaLJhP398gt0rnAf7gxaltMMyCjQtnUNpU6Hw/dLnpiyRUgwT8J9
7YTGESssEJ6G+0euBe7cn/lQoA3x5l16wQpg5ghZ+fRZveYT87c+mBMgFVVHtIjZ
sBGMpLkndWB4vtrYVyPG6EDjqIJSpsqGvevi+kgjEtY2sWRBJ2dyZPZ5KH0loZbJ
VnOQbyczZvpZknufOr+pKOOsCepkb+H9K7B3BLtnlD84xjNy64agbe1lfwfM36cA
rUv154O8mfpoizUzs89Fjgaj8g7adNLw5bO53YTP/LZSp0VNAJQ2iU9BDfC6cIy3
ifJAqe0MXfzdTXq543Qbty5L0B0MoECloxZpkDkcCBSaF2ShvPIicFPkL426TDpN
ccSY9jUnGVysCiszxI+0dLX6yV1rLAdnWXXKzi1cHViV5Lo3O0NGL5OIHPy8yl7g
peWPWo1i8DN4pjc9rm0DRmzQAM4HUsSm9fo8a1dtVOzMt5SzejInGNHx3wfcSG6A
4b4lklwWItUn9nb6CMaTkhc0wpOw3g0KrPqKtDyFUeugemOmfxVqSDZoGugP0ez/
anpgvEKYwBr75AQ6K0ccM4XNQuGuyrvrCFORNowISaLHT2HhErxzKEhohKxNIx+E
BN8/F22KmuLlAj/Qc2ztQul9zdsTf23tz6/pu7pZT4BoBRmC96XFV9ELDY0oPx7o
0tIuktAwX4VP26iQ5HTRpl71o1tVr9vKZzbWGK1lUbshNDpcOz09PDl5L5dKtNVf
+6Ev+Y/QBvQXCr/6HotJl6YChUqmZnPpzb1CXyUK40AVQOjHhPsGNBL2Z0IdQXH3
sjswoFNBcACAo7Z2jtVrTcMJFGUIz/bhQA/Hjh2eAUWAbzJEh6ZN7IWyaY1D0U4K
iaB7h2/bDhpVBerG6trGYzQHhR6J4M9IM0iO50AKeegJC0PGB+gMSXb7lqD5at/A
XPOHuPU07bkeH46xNzzuw0pIBPbw8HjPrBQC7JoeIZYnIWrQLvzEsTyb63JO65C0
GeDibxburQCylvJD7jJOzEo9SgUi7aYuoftDreDWj2R77uoPCW2D1dvqACIdzKE7
OMqdHmGlOwK//fatZqo3yOZbbXBa6I0A5G3tcUzlReHNvW/3YR3/JkHgHf36r+0w
/KkamWtk7QEKD9IwqFeX5xPH/w069C3+tx+SXXUm1k1Y1FmyYbztBSvoLcayWmV6
q4E0ohrQwjGhjZs7683DUz2irAA8MBl4h/qJyXI9nwQKxeOYET8l+HvAlNJjSgsY
WXmMgv8YWHAY5lAA2Oxpp/ukBm7xrg7HuUTQZeeXxSAfigCd6C773ju3N+CetgwS
hkPwIua7Mpz/GvW/U9+o6WLGp7TC5mY8+34pirHFvGmPJJ+2sVnhLD9qA9PCeFoQ
6bBVenrgmCbFnpncusDU44pwuRi8v93vOaVofnZDKUOqFdjMTKzh03ji5VG/xIlq
g+5e6+atjLkD6/PL1zZaPU/x/BPb64sDm2rnVq4wEy+FYEszPLkSpqALY3LTP184
RmeHAvALuKzZGx1nWjm+djG52X4DrhbnKG1vPbnb4vH2K137azjtnJfdVEO+CoZw
jOUU24U4wkAGhIqqWhGsLwP1pMzIco8nao6OeFNElvOQXd8dOSd5e+Mgg5UoUBvc
Zkyqq272W+OAzHFghmzqdABpp/DBIPkYgSJzxawRsDlcquYQcaIRh22pIwQlAF79
Ip26Hu5904iRiAR82oYC8fI1vOf4Eu1eCgE0pgxw7oF7Tq6Qk9KOJZjt2C1qWOrn
saXWKg8/qPhDZrRAxd0qu09IAWbjCujKHVVS4Z3iWwoHSt9ChPuvr5FMHtnRIYYN
WJgVGG5YrBdHYLyHOYHtxsUo969CYG1pgmti3fYqtlB1/h/5Q0IGLu7C9oCnJ7LP
lTKn1Z30UX2xnWTVAaP67EmVVrLrnHsa7lrmMA9KHz00FxwSbXVzv8w8pWOCRrID
JZhMUm5sUCcqZJCAgq7YhDZHMw3yMHiQ4SuHYVmR15Y8uNrcbceOG/iIPXSntiAT
usJdHD4fAbfcflf3ud7EN4F3EfEliNCMlgghFTNWqZPzI2PctAEwZbboOg5Elx8s
mDtRCH3V8oQDVhPO6YKdgAELjSQM7mMZl96DWIjYsZgj1zMtW/wq2SEjQ3UpbyFn
nAOQOWhhnyASOyqtIvF+Sgn2ZYbxedRBoHj+66yczP1aXeG+Eqp3PVSrltvPLZ9L
MStuD/X1aKADhGIWqhty5Xj6QY/QVUeSLuwcHeZXqHsXeDPp59l3z33Kfs6qq2i9
Tt91fHZxH7hwYQiuTv0QLnwOExmJULzy2cNsGMvq/01zeMydHYWCWTtYsq6oKFJM
ob2VufCRBPFSOrvavrhzE00At+cisxwwkVqolBex4vlpV24QIxLVoYtvdeyq97my
VIWb0TuvSs6UVyEJwn9OveWuOwWADlkNFov/Q3XV80cMLdbfbvgaqxUPSk9xlq3W
LtQQHgYeY7IOXaTkvPWxT+lMj8o2UeyFnWMhIwLLO57NhKEAmQRGvqGnYsuVQTiy
zC2yVGW6dNfA4CSKBxgQ2OYo82+FobnN+18K98tRhHZSdqHZkQ9aOJvPGTRek1kQ
etEVpBUkE7w24ZUKfi+87tW3x0KXYr7lQst2yaZxYIUHUny7qCUqS37IIj5znMsW
IQURWs0BfFjgJ3+yvnf/l5bNdKHFWmqOXV6W626I7x8Mg8Gl5njT54NCUzv3gS7y
KJzdjnUb+lF74/p5C2ofXxhhaUZ7mlFKuTw184L0oPfoZCCHVmnUm0jaGB2Mtysq
W4AN6sBoI2+eJi1RhzBDp3MDxKHZZmquErOUjn9gbIqpbLcGlop3GF5n9SZFVarV
MQtkMK8qlbNH3UDNqGZiYKrVtiwZav0a1qSqPikmgygfRJGpC4NtTLzUdDXw78A8
o38cso247xFG5XOA8DxdBNEICjINY6MRFSyoAaqfoKmKfB1ZvAsWLwRHBeuvHF33
Y66JEISvVwgXs/9rR1gItYtbRkEmulm68PrYSfVDIYM8TQmYpxnlRjZQTXRPaJXn
0+O1cY7BMw9kED2S0lpTIzUHiMBsSnMWtGmKauFghBQ6T3uNQpBJrA+9BS2OYDpT
EaNJepcJIywMO7osnE4aVZDNv5VAkwGVHPBkA6J9NW8fKY/p5G0Icz4P4Uh1MyWI
BN/LNKym5SR0qivij358YuXBRIIFaDGcRGKeYECQHNS4O1upezloIvrI7Ka0X/v9
WFySFxcGtmrHwQahRDFdIuZ1Khloakgyuo07STRpt/Iqy2GB/rzCIWWHQu9VF0nF
CgAwUG/NQ8/n8W9Vwslo00AJiSXo+9uzjIB5JRKojGThwOgjq4+YLs6JIFfLCEak
gRJVeUUcpHZWp0gm3oTQCy4PQN10GGpvAV8fuz2kYGdSHTcLpyaNlryKEEWPMJxZ
j0yGwVw0M+Fm2K1FOsyDcnFBzxIjeQvGtcxOF+Y5cUb3MGoUuODBGQGIef9aw6Ds
cvXVRgpEdUl0/J5KvQhqNpOXsKKtoFeJ+tL7aSybnOAWPVmjHmuBP61TE8HdJVN6
H9bMDbyXFDFIJF4dJSz2kXpf7uI669wUi+N59jGfU1cj/vci90L62K7foQyC6ewB
2wHh6PQgo/FeKfJWxHiNvmbJvYwKp5FPv4g0JZGtAhKyh9zpHhqXNOEx45zhxokb
dKr4C/OBgKP8DdG+oAlzAfodD5F8FZZKr2sgqzqIGRMTs4qVlBOOoWhDu0ovgyuo
iKk7B6FrRICW9/s/QJM/UABXJ5ezXXEWPk+DW8KXktrSjHVl40i52M6RF5kOA0UO
R9GqKCq67kghH5mXWk/Y7y4ATb4ljE4vgsf7mWIcTHVKVDdb+tBVUVyHSWvxwCO3
1ezcIrWT7Ktq9Fir6GEHWY4Cu9HDmDR34io7X61lbGCktfTGAbD2DjXySpxREVSd
K0gX9eWKDOM3feLw2mJNkth6tGPm8xbpDuxxN4d/wovj695Tz5LniXyoyBS5JvQD
kZkULqohzdRXN4OGQFZFYBr/GbBYuoT3oCSlEjs5JteEcdbgncRHkqZU6P+HbnlE
OTK9hVLL6KZnR9f7u2jjaBct7EPWu4cJUuaHUt/s5360AYymxxGICOQfgl6/edpa
mhO10ijtYh5WU2VayPZbdEj5E90QMgj5ijnAWv72EMF07XH2cUhg8Mc/z1MEHKhe
AmH0Y3mWyZ6gOhQKXcV4gz9nz5eq9eviw4icvNH7urdn53Wm9EHzlGG8WRmsFJEZ
izt5FbfutNOHbEm3NWkM9sQHttSZeQEw3obfwrL4K2cM9c/5xaKF67N63aivqJU3
aea4Du5pnw6P57xVZmttaOij7NNagyBkDuTnCMsbIK1BgrNB86XWW9Jw5einRQzB
JrvPajGaxlHxUNdCbfUyILVbQFsJ3Np7xfyEl1h38thKmYCjBlT5/9ltHphlA1gk
PbyH7+u1T0shX4xg2+mpauDzgxVD/QRqgO1JMbLH11GJF1zG0SNfzb4f5hfuZMze
n7TERryzhtOC5r/srgVfx94G/DchdHnw+B1RX+8Y441gDy8gH6uIpix3gCzG1qb3
bJeXpXnSop8Ld95usD+yd/DCSPDFhJods9rOGatMDkyiWL9sS9eE+SSDDWsZFGoi
hdpCTB4UyogO0KXMbY2BOW8289v6yiKjiG4F13FzMgnqKhV87/aQfgCBw+7W3abr
EQTek+DUr7Hxo1is74bAPsIjQSXjV9DgZHbC4dGxw/Y1cFu3K7IC48wJVBu2UnUJ
4yoSJjcCFU/rgl3Ilx3K6AocvKUuxXGbhux/ZPK6RONNAu1CqlciGbpnmVRUf6EW
EX1KkPzDqmgQ300dm2vjA3EmKe/21IiwgvzDrmohMTMrQslgIGAfHEgP5QP9MNDv
C6n73xGO9FRPDo69NJslGEYKZok2xHQv/GJ6xlDGNKL4BGJRJgSTjqN4Ohjs1/GM
EJIbxcHw3H+dGbDPz6Ty+vvzpUBooBKk52Hv0bSEm3KHEI3GDSbKg5zV/eC1Kdnq
1OZmopbQn+s+PTtFN6lbdhhnasU1f9tk08tpRTQRK7Hg4ER+T01cqY9fixQdHCtN
lsMm4yPnqdSRm4s65HiUsBzKex+FW4vLWQqdT+zBZy5cptHaq0t1qaEoY78O2PpC
lbc/h8+SRF0WnhqooS+88QcBRAEe+0Uumpkp1Ji3yOcrmeSMC14/mcij54ZfCBzC
GZCSrdn8Lh5EgV+j1UkNhn6wSWkYeTneOVWYtlYoDog2wlhZgVctXnoEsqSrLNPW
LTBfgQRP6/VLaNwXGcuSZjhs2o5nteaCB5qhNMUXlxQd0TS9PLpJ3YWX+f3pVWKC
R5vgo0C5GTL7atxyF36qG1lZ3D1Tol6bW7XTqDS93ziOmQiXMHOdFsn1j8Ggg+fd
1l0K7ZsC6O1DGx4upSiYsS+ob/t5pqPEboVwM5Bl1p40KNAABxwDHfVcyUaPTwAx
2qUD17lli+E3iqJTJ4q+B9G+BSHOoUDTGr3aDsL4lVd7ugbK5sz/IAoYpNTTPR6f
aVxUVyQyeVyNEJs8PrshQn/4sst/tzPXys5DwjqsyjCiwTvhP8M3HTmZncAQL0ei
mSV1QzMEjVQ1eufVsnSNAGi9SaoLXyRPm7sB2MOFy6XVL5ZXnfjGemN5Y6g2LtBQ
Rzqjpqq4zVUiuRv41shnR5+Gr+liaDrtFB4ac4sdhkoT+1JcPFdg7++pCktoKOiF
aQZTSCFbQhNXyhWchzKFj+s74T7q2DzBqm8ocSr+qp19BsQw3OLuIsAmUzVR64hg
eKJHG4LSUME8lN2nEmZJCWNLBgvRnUO2ZunSdyJdnapzwAzTC6QawAecXTyp7WJb
x8szu8UHrwmKPQKDFOLGKG+o5B47TC3T44w1WDwYtXzFTtSI5t0LwIyfWS1zmzHL
2nDWbwNsn3yi0UJvaMu2PRf1vOHN60gj6GkMeXGBDy+N7ORH0njFKri3ZSTHQ03p
W5T0R0jcGgWTtnPRAR8RbppqrE96KqbpunFibGkFM6x6c8qrHdFRmcMM2ugQlqV9
5Ow/ej0zHUwhXmtvBw4yYeKeoPIs0FdWU6T8NuTAOHpS8LdU6t1KBQjB1bvuDUzv
y2xfSI/huiidE1MfQUXqlpbG9B7KAuL37Hlr1jxaXnh0+0FO8lmQZz+28NuFTfP8
tSI7MbogVdajkV0uO3s38rcBJhv1mOPmhwcG2Zdgq9KU2tORecyNFR4/h/lnzS7X
LT+kwf0jlpR/hr8KjVJDyDIEL5YaZYZPsWGai7xt0fP7WuWE9dYh0HnbnjhUskK4
e4ler+WWrsd54H4dkrPV4RStPmjBKIKPowxIlhdOz1GuouRp0VXHlMNeiSWNCqSN
HNbvnoTZwyQePF4De6rUv63VFnEDy+X1AiuuMM+e7DSSeCEBVo6Qh40eFzzkF3NE
296C2vIOxg7RZr48aPptHfp4/R/mcUELogdzEYSWTED3ZXbByS0yEIp1T9IfjfxO
NpptuKpwpFGXoRYF+C9UbnUUkR/o+0hmsZY0upqQvy7H1L3tkpCqRnGPfNo52jxI
03vyfMvvL9SUBxcp8e8t8N25vFNbzbdYqnDZUm1moCB3tpDEuS8rHHYlB/S9JXpE
Rgy1fZV8+7R5epn/5JJF8EWxtfx2+j1b8RJ2dvOtPmMQnFHZS2jravBNef560oXH
M2ZIVlLC29WVkwJ+hE7B3XPYpUrF2qR/3B1cFn3Ma6wQFZe322bTLZ6O/pZObEvF
kv3on7+hIu6PFOTmSjy2LgF+7+veQWG3+Qr8eKL9aMXZhAUpxc7gWjmbDO0nF5Va
uWyJYnX+MG96e/lt081EoORdx7p5WGMr06w/Hlv04tv1wweRhwll2zw2to2XgNxa
oPFvTRr+2og/VwCJK9OvDyQcwccm7Y+up/LygHvNh9PAz69oWO2XArds1fIrEarZ
9MGSvI8IQhDdz7sXqehAzhETR/NUfd7aysvoNWxav+F2qufJC2nGJTqI4moEbtsq
eGP9FBYOmSQZgD4a6iqqmcf4m7OkgusU6UZKYZiNGHgwc9bJTuzT3UQL+z/rs54D
5MkKOReIj/lxbLVfWdbKQUfGauz1xz4XrBlfTLRyhVaiWjkE9CqesIhgUMniAdBo
xTKyqvrHNU7/4SGDfm8+OCU+CC8PhBc9MFZLYKHr0M+dIz0K8wHNGiI2BwZuKtLx
ydrtbkHgAA7+otyh0+znT76NNDI2ftc6wMIWRU64Epmj04xomGEzCGnPzESwFjgK
stQNfBrEmUNxhppN91P5WOmZ841Tn6Fy8rJn/tkhf+tVqE09QtRTPoG/E1NSMR+N
dBYtjCu0srCSdu+egpaMuF4zupw/ClOjS5GrxeSk8PGTU6n1GjJj8rET86tVsvEu
LHYaJcrnpVtvy3WzDFXBe37zOLiCfDlf/zMnrfnruZYc+OMvZxGOE5OvHrsHDUxV
dPNSUDXHtFuetah8s2YjfQk2s7/oJ/b6VGKxrUtRaz5CLBqzHb84VLap+ewhyuOb
zOYYdBwY3O3COFqe4/288Z1PzAF3Zxn33MVIs8jy6HFZMpMJLM/CRnK/cXWLUGDJ
kZbnKrXIOL3HE3389P4EMo+GUXI4pYQA23D23BbEhJ1TBGsEVAl/u3arwSA0K00K
FasIOovcmELAWzoFVDUu+vX1QVZbfSw54OdybLKwV03nSlYSGWrJD54VTfibG8Dx
+6fj+TG8JS34UxyNHmKRnMNd1uVzFBTwdbEcxyIFr2M4LQ++77cPwQBjxRUFgm2C
2aG9LmdQDacvhA9CurbTeiKHN9mslIXNuRiNqVTJzHrL0zoPTYHEKdxGq5uKQSmk
cwzd4gTsXqpYw1XFxa7LxZN13xR42ee74MYCzGW2N92EAnNVz/TLukkzM1F5hgZC
JhjFZBtZwCz/MwBEx9rLeJXLaoN1O+kWhPLabWGRas1QbL/KLlcw1Bg9SU2/qoGG
+5+qrjwijBo6fFs9QPR/ldy5wOlSaWltd9WkqTUVP02LByOFf4XDlKh0Nu9Y6riz
nhjmrT+sgLBFmrb+P1Pi1hdpbZrwgkRvUs2TwhQvRy0HBEUELujqS0VttcTbvqSx
chZkxWkGgM2kCECEGbgDyCTKAHAkOhLsdZr2gZkrym+yYB8N8uDM5eL2S4lDT8fA
RxtRnoIOkimkqmahQLzaiPm1F5G1JZi6vmSvvLzPtqRCOAkmGVOGVdOo4L1hk4jo
GZQGms2IQZfrIw0kP/9B3AhwFzrWNQbFNf46McesT1J4fJOCREggEhYxpWJ3CBlc
oA/QNpzDgBQZiaRFzO50zPucFNrBYIyLSDwFe+wjKcNbdzOQ0SXsvqIPrS7PZ5W3
ZpQhz2Id1AJKJHwkYoYrV0kQudqhzkMRWDSXMt8xEbTjFV65buHo3fHa15AspSex
gxTcK4bvQiegANG0193r0+3qR9bL/D/n269x06he4HNAbAk+XEA//NhbKwshGkmb
P0Z4nEQbyarUXGWrjvowwSfRa7DRnXTcetRqgehYg8X3YYc+HzL77horcZhmX7DM
80aJL3EFBoD8r7A8fvmOfIXhr/gN5Ykuipfi/bdD3/SXLWXY4BLJgt3HhMFl/9tQ
6LhfnwIWBNsrTcMrCVeOpXuM33rhipZGQRQZmb+CPBu/6/43FCkM0tR56/J1c0JO
R+ONJwKMc8ofnis2KhsRueelqLlw3kwZrEvXN1fv1DJ8yAey5jI3r9VzlAmOAxgf
BLR1uWKwCnotuhThrRJe3ftqOxh+pANyMzpr5AnOmj98up2sdIDWuaCAqZ77rHWk
N0HKd139ndEKxwCxvoBHCVbd2YFuP+4nuprbo4QfC/RSRgQGLYyPd+06KSgunurV
zUwiRF8yRA4Ak3WNN1+k55vUrZ2RWlHPb1L0rykigDYGrbWS11MOH8+NmvXMVFA8
vdmUFYvgpLqiCcEcAw5OMIJVcE+wUvUq3+NFNpL3iHMaVUG1vjNBie3WoqMDy5tp
bFdmZYP9CeBQg2vhYXcj+pPSh4KqcUc8VUU7xKBujPdZgtNFUzXSD6VVrqvKRR9g
W4QEpj6YwiBOiBNWFt6tidTYgI2qzZrwOLDUQMG6l6UyJnuj0H0+VpyCPv/spReq
BMUCLOAncGWUi6qNNxevMwgottKIWBjl1yyyc5mTKe1jTdxVww2wt8g+GDiZvjVx
tQIzfOrxcoY5/gnS2gDJGjevHl4i8lSZshgleCfD1usjmoB8/AJf7rLRO7zquXBU
AgYgrtOkath0hx6WiEHcpjTKypbf85OmUKnhpCKGH+Q3009SvK1C6VovoKFFLeMe
skUPp+26vZ2rzbncguBg7ERvTiYUIg30XQmbP6NpFBjMHNO2eVkulHuE70V0T41p
GXkO6gniw/ZFh+VVpPIVgQ5jnQC1nitcDF5a/blXoqLc+kuLtRujRaXkZPvfMLpC
eZ6/mbeoEvcJZo45psaYp4WpzXUoaFH/8z7TssVhJqdWi/RG1INGRYA13dCgf41Q
1QIx61uhV02AsKx48IVHELkq/+P9N6I0ct9A/CrlmAf0UGn1OZmMk0u2CmbBVco5
OVvhjblYlJWtJ96IGM72hjuiIY9dhTUoMGEzWpLvtTq6/XAUTL99tn/DhrYqN2Nv
6pAHw0PHSTUuR1lYHUF6ezVGpB/P3R6n8ujXHJeFN6vjTmEVu/xifFFYs0N5g0tr
ZTmiV4pZd6C4yVGU+VGU6sZrrDZqA3bUrFBSI3bTXh5kxCWXLTYiN+hm1dcSsmhR
NahGihoPGVpkc3DMIyC8CNwnTUDwW1uQy9CfNqMfVz4Lj7XCwx1qYIOfyVawidaR
PIC9kyf+F+wD68tFE61DZXEjoBo9E2Jo9R5gOrZFoulty5uC2jAp/gejmxlvVZrY
EVmSHSBdK/91E6Il5/E5/uI/t6d9uAugJA4anyFZJ2ow1xafU2enjEMxJX26j8Hj
EYqEebdHzLFwwxPDpbtSYxgIWW0pU2tTmfhxwVQ2b4Iq3XUHK+lH1PkSGP0pbIvT
PDutxmhaF4dk43a9eL224atXC7nh1dRQad1d6Jxqx1Ks0gE6+2/a++kUuZqjaX92
9QP7WCkQtQMQyfoNDtrqBewtuDJ8YEkFxrnrnGyV4K4I5LW2LWPSZBtmHRoM1K4O
ttGAW5Xq+6xtyAczaUM309y0HSie+Dx31ned+cSswbSvl0XBuEaEY5gEGkHrGCsU
xkOArLWqXCdJpretGEwQGHLOOdxDMr6JbuhxCNY5rNPwvmOcT2a0O+mmzHmaIatM
VdHhMAB/Ch3ADFRtfBZp7yHdlIxVTvob9z4IXBFnopeVJVemNyhldd89fraog7uz
7NeOJHL7eX+PI/LCXsWsxaz0TfgXzBn5A9k4so3AMQ6PZb4D1uELkSBHh0xCQ8LE
9XwKZhXEtkc1WxyLJIDwyjStpCdfnCr9YqqKFhUrCeJKrH6HuAx2NGHJVvYkFxJj
6qkExHvsr3bS5VwYtwnX9NNOhJhAQBoFtlF5XoKEOycHD/DUNBtL4wgkTUgQOrAK
BXrNfBllGpAhjA2NGbCae1r2AiVR75ZifcqrAP7h5VOfe7lE2IUwbGmr9CF7fzzL
UkmmWk1/dsQX1XkTfmZB9zL7TQ3j8EOL5W3P/8EWixIdnsacZg1v5nxSY98m0mT8
JsyNko+u3rmbREWoKVGBAoq5J/ZbpQPjCf1Apd6YB0keefXGd5czWPQXMvwdVHpW
X9fzZQqF/4PJJ9G6SYAw59RIRqmw+fLGACpL9gaBHFfNeQc9o5SBZmkLI2wrnhYh
WB0LpX3E2S35n5cfJ00NMtD2c0lDB2UpIXhGnKKVEp9GpFrXBm/OGfp6IxJTsSUA
crwvv9w9JU0mP9la9wxI6+xJiVbFdzwEOw0SP94gY+ub4JE3edd8RJ96omgyc04Q
1TJ8TpRhM/7LqoaVuit00n5is9SMlvuLX/nCjOk3HaIgGwPmHKrULbu5WKDSK8yz
Ya01g8T0IYwszHvJqq0WItbOpu9T6/EN4YkWM/NURxrHbrH1vv0XqLFnHjIVUvNL
QWC2OZfTZL4z+zLy6+ZKoBhoRFzfnCVarVdGE8JBIi4X83svehpOneVzX+FnnOja
Dd4iSs4SG963tE5RRVdAp4RNaokKh53Tnw8pILAXdUEi06/FMrqmX0zGBhs93BaT
RP7C4b46B2tOYud0rDzhbO4ugxKuxsMGX6O3VUNu/jVx93b3vSLB2j0MHNKTineN
aEDh3QhZxW2t9e58UPyAi5hsvJ8mxcRJHhoN/+ZE/yqKbPO4N21rn1wSN1cRFljA
GEeGyNgrnZGBAUpfpNskijQ2hOmh0DzKL/J0au2Mn0MCeNG/hc1S4JvveyBTEwQc
fVzUVh8/Gn5yx8l2XrIFHZ9YG0+3sj9yZCl5d4blBYYHK34dalCORj8w0NTKLfva
ozlFq0rqeUU4414H0RPngVwBE5KKAqwEKhOohPh9gvegygouD6yyrERXN4XoYNGS
LspEtN1C/Rzb5oHhZw5RU9ezODqNaNHaYEbgevFlUrplwh4AsRBlI7HoQAEnYbqb
Qpj5XzbqzCj7OOQSgZGQE8KwyDWENwdrr2GPyd1LuPz/ewEWLyI/FlP+xhq75wC7
oCcgoZqx6MYWmwDQD9+c+VddgtDoJKa98VsqNEBqzrCelTWeuBsVJdNyVZh14yBm
4z9Rpx0ZyglE4pCY2WVUq7rxW07EuJ0OsbDzHIENhrKyWG0t0fOiUkbRwBfhYHaL
UD8FnCSQSZdD4GMkQmXAfXU3DucxJ1rCuspNfX2VLsn3K4Baxi8QOhQCcfzZkJyI
ftEe7appT6FrKS180wqytUT3vQ8rEHTM3aSvCWHswU3us5Pg/s8/+ceGTSlauiVK
RasG1hH5EykIY/qNbzTJbAO3+/TtlfeASlczh/blmv7xjW+KihkugHsEA1pRo20z
YdKvNqRCaocypQIPIYKG7aImK2oVoFnnVZehpgym2lSKewNQUv56IUWBIjb61q2V
YNVl8vpKIn0TXMHQuq991Xnwx6UQOtuWjY5Nvn2ekh16ERahiOdBsoGpzMY4d9O3
n7kF1F2yRDo/cBY+SkXd16srhKZcqOW2Gimm6otD5dgul1kDXa8/P5cwQ5Z2mJiU
pPp1/DY/OC0+EK9kcTmNP0Kgt1bqJ/oadjVxRNWe84X2GwTwh2c5Pc1+BMrpLoNK
UQ3d3+YcZf7v0C2jcqSCFeiWRdcXNJgwg0Aof8IOX/M7zWNqsrxd66LYc30qJe4+
tjwDKje9mqMEj3u191giDGUI20fr2M/D1rGKTnAOa0+fgei7XZ6/sDpOiieasDR6
0qT/xQkZnjsEqYeXZEJjjwwCIy0Bgk411FIaEp6cmYPKu69tb3X8nSv3FpBZCVr1
JP4ZZZ0rDk4gyhzuESFDVpqQScXfJY/95o9GzmnAgFujp1SnAONyZ4JCI4CYEzXF
Gx8+5hJ7CqqxNRJUGMrj/gOxQTmgs41AVgbNTJDGvj/M5s845aeRWrzzb3YmAPLa
oOcHTn5vFtC9qIyfbEorGy06BWpklavTGxF56qSITM5uWuKUiMLy3yDdcOTGiYWy
DHk3oEwhpB6tkj9I7VxicTWck4Dc1Vplytv79gzldZ11Xu65Xzk3f/ou/cVQ5BB8
TbaJAPmziKun+WIhbvswoVlnaSqFYcc/UKaJKMcgov+kZgKNG26GzsxFLBz56s7P
cL5lFfwDEuVzlEy08vPbUL7jFj78r8ecC69482x1W840olBmKRhAtjNNzQ+BL2TT
XZcEFYmfcu4CzKvIqwCN4YqAzIGkLMCePa3GSpiol4UOXgI0q+isCe3mgAX32539
T4HmlwlvPffIXeoVF4THqNTnUDQJHNpewhFeJt+PhRYIpmaAjTu2XpfAyrhx2Vvk
sETowAtj6WaFtKKntEMDToQT9rJA6HVwtltQENnGGWEPDHAJ7IuhfnxDdP19pm9E
jsM7UrjYJyTVmwqQyFrgjnbO50r/x7K6jAbqptDjOIR07PN6GbyksFL6+N0tCuxk
csqWu4dg9Q6x5fDqIYCM8L7H2jk/qBCZ57X8brqgdjclh2QDDbgQQD9q8IlPITeM
lbtLfcYBJlR1hAXDdpavRouZPmRZI7KlxDjSflCU1xdGL3In7Hv1BuNJK79cF34p
RtZLYJK7uS+6eo5Dfoz/wSusj69QQ9lSpRCqvElw1M3qNLhwD2uEilMCH6EVIUiP
x+E+194wgBRdJsMWLOhWQqwS7diOz+iK6KXN7mxc2BI/Tyor+XcDlwxzpUGfvyg9
m5/zgGi227zd28oVK48XolRCtvNAslq2iTQADGaiJp4bgHzHzbmcM2F3Kuqo3Kxf
CdEWWogqhV7dvZ7rBXRiJdb5FyUoF8s4RELzmI2Psqbgdud81sLqA1hdWYRXVrgV
WvLpjNPTU6OUAngXVlfkQc+b1DLCkV30y8sbMgfSdKLL3KD2DDRP4HmjNilaI7RN
16kBhZJPADdgEWy357nkk5nH204xWdjFRCB3or4SYdydC7KFFGIhUvCbxpxl3wDN
SzPvrwfwMd82wGaTvhyci8ghFghcXDOIeFOSUkr9uXt794zFM0mOE8Q5i+xpE4f4
CCp75f1zAl1Txn2qk5bE1RkIrpg1XPWrKZc4cct7Kor/Ti6owWpabWq9rVFo8seP
rAFsQHGKP5VF3UYtq8C5uOFTXZBHMCd28KTJ8kPSKCniJw+4hhTgSGQ6H4ID2vjK
FmX5sihGwO3THfIkgeAu9GJlOYSdrNogK2RODDNJtHZuz+LbycX/ZDYIKfTzibvS
vNlvD46MZzm4GqxVqXBAVwFT0Gw8XYFvkO77DMNtxVvnoIwWJ9j/6kjlK9Pd2aun
bxQ8p1yItX7KvXS8fRoTqaBQgXJ7IoUHt5HQUOPt1HUCe2CMxc5YUfL7ECQCoM7T
+kNM0G8Twj8ua03BuYEfRTq+Jfkkvpn9GckHNoqepdVxHzrUXRuUWL4gldkwM6Ca
n0dIJKoxcZ9RF1fy/QPp3kCt1KVV7VPYKkoBleitSgvkC3nLOdGgL5+ghd7K8mr6
TihM5pxjCYJ32LWLh/eDhjJs+d0Wnm9MxWpSS87wLCQvUdMZSyyP5STmuaq/wt2w
Bxqr5jNJ/euWiLMLVNmxa/s8TrkOijpOOQaWZ4de2NnE2tHZrL+yroHm2QEIEfzk
I43rQIfjz4wbyGTHsXzrogR+IyPRSTyHE4OA2haUrQPxYjD1SqDXkY/YbzkX4MbV
dWsVXVbT2ZJJz0S76WOKkYWUj9cN0vPYuTA7HyKQa+xzWBBgi76D4Dw8eYNnc/Bn
wWmysCLtmO4mEplDtSNaUSLvP2ZTpICXTZvYCdmVgUW+i65ZxBN0aYdpFsVhFxYM
1hY7bnASJSWnVkrOgSuHU8uQ7LFdHFFaiT0hHKaIPY9a2e+d+cnm977tWLryyBbC
kRMEOtMrxHDyVmvTEjX+t7rLK56wYm31Nmf4jF7GbBcPuyTLbFsvzt/u+2NFPY+s
mfob5iJsZ2BPYBGq1lSZE9OwS3dSNSYd5gUDlvzJ7e61bwGxWHG+TZm8wQ0+GWQ/
5ukkYIP0FEQ0+S825QahSzhhpFkA/vobzruCCriSMp4hQAlJmQ4D0QbfiRTQh4Ti
H0rPGrx7PUgZrU3tQnHikv5vofrxLbZsgV+KYVBoyVfeYd184Kspd94Wm3Ugv4Qg
d9TV4N95Ne660UL+t9SlwqyF7aywEgRKEiKHQvx1E5iRJz3qEd3FCuUkhnCzXzZ1
h6wvFI3mSFxxkqtXFPDX9yj66GiGHcSHLY/JnxXUC7tEnZ2hie4Wa+M+ioNgUWVm
heN2hhDZBa8BJ6/76RyGzQLyJ9QWRgRuahmF/OvTHHQv6vY2VA8AKXEdH8SiEFEP
PnvCjMGQAwxZeK/tQ9sHPeFJZ0FtSNsseQ0f53b9LSvrdxpf5MoLTf13HpVKKJ83
jzygHnR2V5m+gbuH+qnera8fgq1oYJASRL+fJ2g733MvcnXPkkqdoeD2PSPg5VRJ
wLA7sH6mBEC15ikW5PJkTP21Kjla+scrVhFQS7ug3DwIH+bqdRDETHxgFcDtTGoz
wT7VA9zDwCtn5iFN6XSkCJGfstOXimHgOiZBRRoBwlN7UgIWRtXTksoFOH1vBW+r
jVhXsYWGskENn/lf8FbGOv3UZPUCv1nFGcPNpdH4hgI+pnWAxEKyymz1Rm8Eq9Lk
uzSxqzO31eaBeokHzkTiAwgnkvpYrtqsKuSdlYvYfvZX51amxYAqy/MTI3f6KO9S
rrcIMBw+2Zj38JfeynFHEG5pyM+ouS+PcTOSJip2Az8m9WHdgbXTHDFgPIwImuh2
Tu+yaGNqNl1rfF2GqHCPZl+L9F6bgRCSZHKJShSP3YliydbMeVNPx1R3Vm0i3B3Z
VXJkAbD/2/VqMyCalZeNqrVAeCjPrXWLLXqaOr2Y9bZ9g+kH+KjDCo/8eDu6N2nC
aH1Tmgun7k8G/keAWFcwQhb9TXiUgxawh0VxE7X7U6/pbRvai3Q/W1A/dmTBl5HT
gpIc5ewOaIFP7/lXJKpvcH5EUc5FyPqM5gBJMmr4/piafdS31X0WhGtofe8No+RC
Ww2AB1Ui03HEFiefeGpmsqKw1qwtKmXrKfvSdHileOMWs4dAOWxGNZ71OVBeUvn/
aJOfTZCQoKD0/hMc7dxkN4jnh2mbjtoEKmpBi3Uv4TK6vjT1V+fwYPCdv51a5Jy0
x7FQ6vG35o6sLqSd0JJ3QJxbELxsjyZ8R32W6zgAexOEbuvLP72ox3nYq8q8L4T1
619zieW/wRy9UMI24HYhKlzos6WLUvl56xPTPSSFZYlru3rTl1F0lGPoYzh7dMlu
TpiCRf1Ibag524FGQfDizDWhkdPU6xVGUPFyK9itGHfldWqHzModgwlb2vMYbh0j
UmQZITrU0naZA+723cmf1jSJChfzkqCEhXz3t9FFoNU8gZ0KLDIdA5Fb8Xmaj/mJ
1KQipdeVyUid8VQ7LkflNZqknKMnAEHBtNJcFhrBeI/zQL/VRye5JlJX5iPaTSkd
79UpSzHWRJicNFqCeY2ofrrh+3T+bWBQaVLJ7bvytweanD+LBfK8rw8FiDDGFNPH
e7cmNl2SZPg1D9LjpsJqlVXQhC0xX9y7RkdxaU+st4cyaAlzVSfzq6kKBSqaKTCy
hzd6uoZO0rnWBJb78No5PM1OKf5KQ516QMKd7xUthDIuhinvVF6ZRvRtlXgNrQmW
puPpnFrFOJBuerojUU8zlumcok/9C964jokzgHXpaQCwXOJG8Yat/Ew/6UN50n05
6dC+KjO8fqqfVZVI4tj1AaxN+l+h6Lf4aDLm+d2BrkxTqaDL/RHmrhjJHimeBWbs
41xq3wioUbJKDPH7t6FIJGhX3H14rm074+zaWjpAFbJetgKj0/54TkbpiN2JQqWd
9lYPXB7hPbjzdEf1pRGMH40MgMG1OxDSAt5laW8PPKGSnzNNs3LxclsIugtUWhBD
ZNf4X0p4+Gymx92zVfhJOS05Ya6o0jS/naARPyH+rD3uhglBa+CivJmSlDwR4rk6
/UT7nGxYcO8tyxWRq/trKUDsjrPEDJsx8IzDHuzlKgDEgx2CQ8liVB+Q9eBFdsNg
kL8FJ6ID5YeD5Q6QPj7pveZtRxpYi+w6wXLnV5y1MjAACG18cqquS7yYAln1A2Kz
iwPz1A0xyxefx7Do6PMhdTR/TA28EZOHbBg6XQKAI99b47RrKIWzVmcBuS4wdlqf
pDUVleIeb9Qz8zTm5oG+ooLkM5M/yVpjI60OovTEWPS9iI+jTYgHBtWSlaFq0V2D
f4Ul/9ckXo/KY0UFsLP6m/UUzbS92qAcfrONPZxtLzXMR0v2jYMWfwg8dVG6hS1L
vTaejI8kD59Og+bwRiLjIN8vn2jBcjBD4CFBMLXjVVrKdG318hk6bxR5o4YGl2RU
9cFfWnMbsvIrA0SdBaZqNhL+t3gn5szyeMXHXkE7AYtvje9O3VdtfGnT0IaxG5Nz
Z3BrwZamb+ozWfHA1TlDWQFbTRdlhlwzx04ZsjKACc9iszzdgzweA3OlfLe5OXBd
HlSvMgK4/T572EGRLoQCwNwpCjydE1KzZUN6r9FmzOQttR6meZXU41aL0kGjYyoc
05bXSvyAm4n6EksF2T0/VMZU/Z6TQQ0By5z18ZGvfoj6c+mNGelXC6idQZH596P7
QQNYKIC7IS1x6zdsP5aatkepDc3S1PZ5cIPQplXyNUpBNeMY+ubHH8UexkWtubFF
DFV4SBIO7xnwwrA1qoVeDbi8Oj1nQRhE++rcqOI6teaZpXeMtTThfwFFbSI5yO+d
MBf2uY4Q6gRDL9dS6VjgGuMsh8GhsdkJY4k3VXOC8w5DGM/SYeG7/2A2bsSTGbza
cMYK4RTE3dsWzitoKRdk1xeNxWN+k1BBMrMFYSHlBq3ZJA8Yn/UOPELQbm+cgS1e
uX404UgmwoT3p4EPJwg3+W8M405UqCtyqud9cdI28gGYZuMOK5LUhMTZdHWyYZCJ
5cnyd28WAJx1Ds/ADkhPGpeasy5kqqXs8hFHMDW1HUSwxrddN6BNCOXoPgXm4P05
fdnqVKH2eSEZF4wgtoCbGppkbpU6s1/ExY2Y9o8hBcF3oIpobkgq2nXBeXbV+BGU
WBdLpW/YXLniugAJarWmW+2GsJBeXyStqHXuxwG0IYgHNZMRvPgNHUkW5DXLP6JU
8PUgSyiChFWxc6aPsbyybxK7wuRY+siXjB+bt5Vpg7Pgqti2oGjm3E+56rAv9HTq
g9h4jamtq35cta6hz0oL6ALu/BGKqFYz/KwHbuiklTw7k38NXYG/1ZJNfFD/CYxw
cjCFOebHTXXz1GXkYfMp3iO7VkaZMSKuQRClRsOOG6b/589OSKOVCV58GqYnPLWH
J71mTo74EnD7ZkLn/byo5gwflbvEnop9TqrNm3dL1hExggcdz8LSEMx4bnnzrhZi
9ylapQ/f6GK0EYjMP6ePDLeM+TN5pvjH6Kpf7CDLfCPj450tv4rf6JrENzi5BBYU
xUkxXT0/s8A2xReqwVGZFeNpuqC+xoyXwN1G38W59Bd+xdY2WFKXyN9MFn1AcLeJ
3bWdEUGPQD8D5REeJsZ6xlDX0jB/EKZISNlkEVAm5lSRmmKK4S29dtrBm9+hkuI+
RoMse3VFRgVB8pNvVVwF3zmYTY5qTJ0o5qRDul8IVtP1GZKtOOX+Ixql2jOB09Iy
IixKs7EEUmz7FjjOKE8CivWIxvezJ+cwtOuXMdWI8VaBoiNBJFuwcld0lsGsyjlp
A4oL+Gka/k6LgPR91AgEwyNTfIS2FQLnj1ZX4XP+5BgSEzPrdqxutpu8q4Oowyrt
dX72rL+6SCVrExU4dHdAGbtmWiFwmd2UKH6DbQjJPrQcFnjcWprCNazPh/QGX6oj
TwMmbtfoKmis/95mMl4JJPkRSefCL51IxhWTegthWCQDZC+s+zimXl4g/y1orTIm
Lg5WIHUddePA2lGp3VDvIZNCP4Ohw2Otu+xjjrc7KkPSVXy98EELiAJ749u/uqNG
UXLTyKOUX/XBwhSsTSrjzcK4h73Qhbg+ZanaH/gqBBKtLwRv8XjOx5l8g7XlqapV
q/VhyFkMTJPorAgVMBNUTqNHh1afvGMlmpUBdLE/XdSBKmEKNkr+N1V6YsIH/NU/
cfvDnQzVWVV5CCFaH5xZTSVTRns+VOTjrvhafw3RpFo63f/F9m4YEfg9bmE8cKzy
UMqf+/lxovI1gcv9liQVNcQ+HvEoMuxMWopycF+s9fRqPlRssYAvSE5PWinry9tN
mniAR+8yJaW8MQB86I+7NBMLCe5kfJ3c9iFD4epWKvElSyI5E9/AZdT0xwgeV/gl
2A18vJFFuy+LM8uGDMsuTNAM03+zua8LQ1F7sAhOxIiJwBKqPjZA6BNGtN9+bNmC
f6bX/PrdBJjR+DFniHHed2erg5gKtmPkAUw8uxsBA/8b9ejxBOEYtv+OgHF6tz3m
RxqBEp54KxOxo1ZKIVp76FnKb50C2FsdSFFMjD1bEiQQJFs4uLFWb7A/4uBMZ/JZ
KGeYaiEaWK2PxaiJrIExZU4Ypxz+mSFzoofk3E7pSJ8zyJ5f6MIFWT6vcl1fJpV4
96xwPa1tmkdWl27Agx+hVxxVSKzSSN1p1yrIO6YcdRFoIjN4FV5eA72LdnkuTwl7
Ma563d6tB/u+WG/8z56ZuUO4t4EonJi8ZTaFUMb2ZwZsD09HXVjl9ufpcXgIiH2U
l5DEQhN3Wk1EAdiZdcC9J5zmzK5aazaGd5EbSsrrycypWGaR8aEWj+Gjq2p9aucz
LMDX8g8CJF7gUNeoMCEbn1BJPgS4VSLdTGqXnhIq5hF2ls6Tm2sIdJUIGugLhjsI
9RIh8bGmOej3N53GXEcNfpjcUJ2AmrjMyxg0qTPRepQzF0FrYonh+XGA0m3RECFg
DYw2FjuZPlQa+UrmOWhl9lTY5rG5x+9XLAyN2doVtCZSuXA5L8qiUHBitgY/BpBF
JZxnPemgBKvrn8rSNfAUQmNv3oivoGrWlm+MNf0p7dqFsXNVbW99PrAsJyrIFxcX
66RQm4zhlDLfmlut3LUVbSg84TERlIp+MIi8cY3wHzw0q+KjEMiLAxKhCPw3rFuR
9DzuWYle4qMCfd2aPTELUFk+AnzLpibYv1ubXQbtmL3b78uo5IX33XmWfFEX6cHO
jBRDEZJveri6d7D4iS48gc7la5gLiSs7hOPtx1suTVlzXvDnYuWufIaMrXWW4JJ0
ruSnAEjFQpnTa6EcoTNptwf9oc9GJHw1LbqZLLjtGjMBIbi1t1EGTBFrZDDQ730L
K/iCVWBpE8vcr2hIGXUQoEGGJoa/QzDqWQT8M9quQMe6iLvOsIPnrh4MlZx2yaiH
DRiJcmhNaN0lnYak28qFSgXSPE6QzzpuCHbkSnLbQW6SW6QPMa0mNPS94JCeDVS4
G0/UtM/g/G8ZOKwE7g3DISEjejLeqH8KGRIsNelf7rlXWNp1/UWzTkUh+u8ZOPUO
XlLTrgqY4ZRWQQZ+XiYlersvNhHRUjHKAtRv0oG/eUZ5VE27/vvsgyfUZxuvNncQ
TKW04lQeuGFPmY9gZszFkuST5tHIm70DiBY2tFudGM3WeRsRuYfbTybceuaGUbPx
+9waVan/NprrHupCElWRTMUknLEu0bLGwTqaYnQCiBaQVuwGlyg7aDFbhHqIj8rd
5iJV+PYEJYNVBu++R01NKLufJJ8brhle7GG7ZtqSRsJzSGPrt5Jzt6FAjSRx7ewH
g/3o/MEXE4HUAUYC30k6cYXP782JdCdkp32GqUIkIXoeRKBEFb3IUTe2vecSVnU4
PZGYpnxdEFYchOfzJGf/uP6g1iX2ZFwyco7ipolaBlYAD+prJpX7MEfh7sh5xEMo
LrIthhFsjIsV0QrIsius1yHrAFijHkvn0D2aoATHNd/8N/glBfXM1DW+QlWTUJmD
cKYtBnfFJGInlYP8hzZkQ7vPuJxIrtwdAPHqjtra2m/Du29tDboTkgrJX0O/HjRJ
SAoGgKNUYAS4qUdvUUI8LvSsPd9jh5oAfjJcx5IFd/YHsfFrLjyhe2ndkuGF+aiM
5HVbP9VIt1iFo+Uec4U4V6XJcMd/kahonWN/f9Y/uy5qFrw49EaevTZ2DVPaMLud
faHbXI4g2o8VKj6FzufJaEdrIgI9RsbhXkF/v9yIatdXH7NDvgLTOcKRN4sxhKW4
tx8X2oNLfAR1mQBEPcJGQuD3KKDFxQLqZeNZ1JV9tgtDSfCqYAaPO3EBrumvXrxd
yFHLQubczZS3/SdTjx8RL3KZtZzbA6adhFbv5p5/nIr5Qz3sObcIo2ROa7WCHqTn
rQw2NgXXlAh5Pk3bFoNihHm/opLm0jPKvnGMnlIBbRHSGKPi8/94YgGtv9N8g1eE
FUaf7ci4wEPMbz6gdjsD8/TFk58IJaaNvBF7s6lrU0mWJknrs+I5qZPumyWfMpFH
26ji1KvuenHhE9rLR3EYRST6FxuZHLN/2MljB2gq6y3Ai5SbhsOjZ2+bwkHsVROv
ZmGo19VOz2+6GvzlzrAye63CQWp5Qrp1gdAJGw1T7UqA3PltMvrw2OkE8TjNxQYf
dGWjTjwxdWvFqi5aRJYHilJEzAUqLZEY6Gat7LyYJtI5VIKNua47jOsC7gT6ofNc
iDtsyryjM4uOhs0MjaYKhAaJOOGAfy7WKhqtQEmWUVsxM9MvUJEY81avXWB9T30T
T7CaI4v/bzxhR88qxAN63uk3OL3IX+Em/HVzE17I9S5Tz9JyClWtMPfwNcRUIqco
HikNT377Nminc7u5rT27a+pIQXBYpP32IsiAq6owqUdIp+FPTQu9JD8NjJiWJx3T
mHmY4ZNDZ6aKKwlzB2U7F4DlnBqAadzDGvl28Nxp/Q8J+kOvkfWr01Upn1C6GulX
oxGALjd1U5Ms4bzcLlMyzgpdSwEMQ73lmSIwAq2rr16uphIbDmOT59+8vMZMSgwJ
byQZADmsEUk9tg1FOs1Q6a6GceBrZEEspLR1GAhxH3X++uV47aIYb9OZSGmuVU7d
P3GPxaLOGRgCgeAn/YXpBaat9J6cj7rh/iAq1BD3HGEmo0/WQ1eOxt8PV5mfEwTa
nGyf506z1+c5zOlVFoliId2TyYmlSOfpfZXc8+uXrNh5vo/zqTduT5xnf1eyjD2b
5N3gUwFq87BBlv6wWZNMYo7hV6ttp9mQ6emiCw9mdYeK3dmCeGyrPUqzP/0tkW+0
+HvKH2I+1zUbhsxZqA38E/GNhFU35nhVx6Gvq4z9whGofL7Tvpjgx9cVcXudXIko
ZcJUnZ4xCz9yP9nbl6O4ZP5He6urZhB0S4yJPQuzzRo+53JPP/8oiRJciBPpL4Aj
ooiljiBlhUZT3mqnw3a4M+sHQ+4h2o4nDhS/BvwL6fHaycS1lDWzkXMJksRyn628
QgJRO75Jg5VMPy+EaNz5TJZVJJSWEdnk765byuLasB/JeCr+RILa5lwLHIe6LMGM
abxQBcwzP/3Z3+chCk4ouKnIvUizJ/2UwdQZ+GW57YA4ZWSBDHBig2H41s1xGv/E
Sk8sgEfgfbDtlBmEFKyK10RjwijJUu9EztKFcZBEjXQzl7lfmhFBrtaLyd+JcfGJ
SxKb7JXXqOZm6rduGQgdCAfsd1kTaHYLNgLAIfOzRYl0LO78xUsxg7JFMh5OsTM3
wSJmGIvsOrDAOz/HqxBOMEc6SbW/VRAKJ08mLPOxFsOmEa0H/Ee1l+zYICYSbqPs
HdXbyzeyFr5jtNO1Rg67KbFuFfkfuZeCfyLloitB3KUeTxprUe6or4bE8GhjGFj3
omArxyoA4PmD8Kx1XOChKq355MaT0/bsxw4aPr62FTIifmNrHuHV68nSzHENe3k4
O851ExerdcDAOHPdb0CwQXy/pmh2S79c1ttKzFxSiTxGe4dcBTCiorqHtkrfTA8c
O5iv16DEIwnzlHHidZcMl1kj634xLoU2hd+YwUXPgt0ICXMBRF2Xz8LF7+M3tSzS
2MJVjuz0evDj+x5gfKIFQ81hNxJtyMIDSR6UomMVFt9CILybwIqgkx2W8x2s5DBj
1qNCiK6wTKgHIAjBzGj/iVZIlO5hImbwVEosUCg1QidCGNuY44+1NjswFvOdBLRc
hMrHkon4WwQ1VMSm4bu4DDqceMdlR0WTREIz6ywp1XhjaSkdgZRmEsoyz8ydGcnS
7omGMrQVVz2r8hgHIKQL+y8zo6f/FvpxtSy53O5s5jiAuXEVN/s0wgJP5wX86B9R
giZwbMV0vJ7OvuKHDyEYbSYV5fJKPd813RY4Pns5nFhxEg0aQS/oPPphim2N+6s6
hMkhUqNaffVw5KZ2ZoUPV7ynLY4zH2sjpZr4jCST9EUfMxUMkXnQJLGr6Dlu62V8
bOsJAeiaVuf+TTzOidOQQGgRlNuZedpf7jvVzJkOClHlHoBNhR2L/P9LlkT4DoJx
kClObjY+sm1hyUqJzWhwjO5+OXwS0PmM7JuscmC7sD2Z9Whd7AfQw+khYvnPXKCk
kv2jJget4nvCmMiu56u3Gjxcv2rBxRgJkh1Ql+hAKGWLnRh6o+0EfuPV91UnyhgF
QhoCH1O35RYgEb2ihf52UDhexsh1b61mQ8ciyLcU4Bibg6qX8cf7s0M6xk17fjZD
4UJpJfb06vKRVGpzJ5XFSs2BRZaK1fWEG6uVXrLNh4KFhQymhQ0f2R4TEcy/oz7c
ZeqJjGleHweOT/zLFippVyEbCKQvhyC0JAy2FxqYyoHCN8A/fRcqgTnkKjydJkfA
5Ld7bkDP+E6UI+AQ4IPhZhYk6L6X/AV4szwORAzbTUT+ZCdahSLtOcx32dyerHN1
NvA2dsBe93rXxFkQoDZO4kYfeeIcphoR2QalCYqEj3ocoY2dF11zCKHsfmOu9dBh
V4Tzsay/KmoYrDHPlrFgd7CcR5B6bHGZTmhp7YwXeQ8G7sSUGfOaZLk4u2Pt2Hha
L9btEQQZuOEfZ3QyxVnYIogizLf/etkMCUFEZg9h8+gBfAM0EgfHNhbF3MwO85eY
UQWtf7g6vrqQxojEUO53ZdV0v9+Sl3wisUj9AJ1DLKJRZ1kn+mZfQMxBF3oM4WST
ltUYBVMRJZdjMb10vdwYycFvaginKqxJhPMXmCeGSNmD56SwKa2b8MQibOUirt1F
OfQpVeO5gq9G3k2SGFz91g8GUVZLfRH8A/QoTxavcVGfcnveMumAL2k/eICG5KUQ
90sHDZ4AOoarMmE7LYC8iV9NAALIivg2s/Xi2scOCMyBR5dL3mwskQIGYp4EAQIe
icE8u56h5sVhjt9sWH+A3u22u7jc9xKql6RqSqxmdfnz6XUoa+oKoikpABueOYzA
jxY5oI0J6llZrS60MIQr1lzJXIcr87AwLxKqA9SSY942W0VtRJiOkhgQ8RYm6e8w
z/N4iG7OvrbK4vCuBSliC0M1DTYUGpC0js5zjZr3qKI9rpvBFC+yoDGM/xPdIAXX
zoKmaBg77ot80oUkEusyOnvWsyn8U/exXnfmEP8DslDAz37P2aPiXAg+H0BHvUsP
dJuZs9Ctf5ATuehINQCfRLM+hTj1ZgTriBPz6BTwFGIefbeJkI82aFIW0+vtJGhU
Ks36X5RcaTc4K/3hNkKwf2sBjc2m/WZ+I029vT0gmbRdgW/tIVnG+tQ/J+xqII0X
m5/PpvTHsG2WAydjYRepiUk3wt4Dh/Go7425MjAo1elfzT7CHymHstaoiR4V3xRh
M2aViYWtOHKmOO1pO4CoZSmQrR4dkI15+vxTy4G1fMp19mYgXyAaL11QqbBYQHDJ
LbAVDvGbSJVLjBWtMd1fzk7NPqibXBL3bDCWx7bbaaAig3Q1uEh1uK7zh3SuvoD6
pXcEMmU8Ydj5dvGpV/56LBkWBO7WkBfoBplEJysx2eZ78cG76Qwx+LrjPAP3xCxW
Tcxog+lu8bY5jTojqRHbvAkoUivrESi6fVnkU6witRS2ZulNFynlqD4RADG34mrM
ImBWsumM9fwFV6xNQBl2TKKjQy3sJyum8kM58bxArZo7dJSs7/fEvNuxG8+e4TMd
4R/5qpPsjDjDSM1yNrSO3vPco7B90578UUOqrEqMCaE+9he1b/uxnA41P4z3mot6
118rCCu+pkVTeNLpymvGAyYokPqt25NRi5gNTQF/bbpcj9Fx+jkaDbL3KltJW2dF
RTACKlCnOEaEfrr2KvyRSZuzwoeGi0CaxL/+eMjfYW2BZOvZTvEJaCnoLaUdgYyC
j8r0beZcCcK3ez30l76mRKH3DNYuAyP1DamK1WFeZ/5v+pklBksbZPj07HLDaDjd
04IG+poL5Qn9WXSUIKzImZgg+ahrwjpTchqs283B2O2HIlEjyp2+mEtd2Abx9/oJ
3/LmxZijfBtrJbSAMQzuTaYEBrtvaMhLsfe3J0t7/t5nt2NmREdo+g0f2QQ0wYDL
AsoBNlTK3mFK+tlUgBVbcUe15Ol5RHLhZy+ZEP9CdeAja1SntnW3khJFxfWHHEtq
EA/iEXpxuL3+sRzJ59MjKUDJ4DrCsmxx+/EMAziTrLS8qQpHFdKfcEu0B2h+Gd5m
FVn47bI7LgtBCITgBEaL1dj87bjXA6D89QMr/66whpmYtnnsXh2L5Scwghgk8OSH
iHazkbDpAATZcTwE8cFgb68FJl/zFVBdDJZBq6XlLGarSG5czkJVWDXnHTI7yajX
00g8xxetbT4CV/KU/v0LA2SgEr7HZwX4Af3BCiZhDuBBaIZR4V5oBBXAALVdYJx1
o1m0H3Bdi/LdfQ+Ruw7iWd5Z4e3PS1n6XatFr/K5NkTLJgeuc6ubjxnmFVDt6On4
kyW6EPV2Mxj9eBJc9l54HpWfPg1VGN+8/TxJFqF6mL4XzFqidPCBvWerzqhvkv9V
GcbLGsWG7OLKymgQdsHK6U7h66NbCF2d6s+6CXxdDl0VS1VJYtrPGT/K4PCU2Xtx
KZDLr8dMoqcRyWhQelGGP9GXZufGC8Vlv8naVaDZoE9bSVws8/WqQb4FDqOCQqjN
mNrmOfTVAMlbiU0uScyQa0wQ6B/NGGSqoKl4whn7W6olniaxHuwIgpPE86EfBs+T
/hA8byVbulvob0a7WqACSaSaCXicGglAie3aasSRgblI8j32Sh53lWie9BHlTFgT
gBEck8/I3Fg7m8e1rHV7HgqKn3EMIyuF2kbzlit6EQB5TdVdKwOpXSyvP71796jV
utMLWAAgw7N+5Gxq6Mca4rlcUYo9/k+v3ee4Q5Z5Uv6Dcn6si1BpBHl8ps8CcyMV
anKopdEguARoGUP+RNgvKKrGnSvGmHiNxDwznaia7FcooTY6iTPRe5AzhbQEttb4
eeCrkwxR68GsDN0K6vKieXP5viYkXo7fDnFKNbzjdzPhRCE3zJ+UdWHTf+fC+xks
4RTUvmk1z7SPLVR6M63FZgE2vZQm12G0OHwJbeWzhZXnkSjNSNTxPH0ie6BdPCEM
XZBge0tK7/Flq4pSU2h4zFzrKbKEr0vMUofRPxfEIwo90lbvepREzPnYOxbB9Bf8
z3BREa+uA+v1LCoesX3hNB3dcvRgfoRhXB+Z6Xf1A6fxeTVVOKDfjSxGWGeQB7Fn
Fz2+W1WELLTO96hC+QMk+M8/GHQxQT7H7BlLQXSdaolKqmaGZFHTelIOcHXZ6lW5
PQrHpsbATw5kDYr+/2sHmkYIsmIwY7lUDNTCO1VOLTIvl/80Pc9snWOa4qJ+y/s8
mr7g/kb9iczTDOaQgN01uGNtLBPd2p2Rwyku53vpQg0OTg6SlhdnHlgGn6nI2EC/
KxcoyUJsFtT4IYhmeg93BEGUiT85Pg/dNboMtIxo3n9Ly/kvupKSFzjQOmJfbWc+
VkcJZFjaspiFDL4WW9HEVMAAOPicbVc0opI66+LjjPrhP/E/TzZcpkFv3LDDQgkb
7yzttesHzyJiLKInQhEAEziQaoStNPiJ925cuE2sfyWyvFHV6Z2l+e10SnSqdk85
TJWMBysarM3VSO8fb+eyDuyeo+MxU5t+a8i+iF7uDeoMGpDWNjfLc9Wexit4gE39
CG9lF2pP2yfp14hgCSnpu3hhV/PqHfWsaRkyzru2MYALpqvs3RnTAZmPUJ7AMv20
1FhGhIbD8m47AcPWRuxCt5+k0r0gmwJdYrAk+J7/OmWjESRz/Q8Q+8hfN8dVDKKm
iasvI42NS9thI8g8Zkp5bGFFwXtlXayIxyOvoHlYKY2YUvW0vJruxmMr2QASNrG8
9G8F3ej4igpi3DR7eZDFABkwCxS0IouqbyMVWSBQ85xGFMLPYq2Oef6EzpSs8KIR
+Nz3B6fkZMNp2oPoQp/5OB0uAp156t3kbqd/Rp8gWj9FrNTW8/RqlOvaCKAulOka
jds4xhzHWgJlmAL2sstlYPV78tLxmtwt7Y1KwfRhIMGhrpu9+56D0U57GAVFkphD
4Zo0ymsVvwZezEZY1+snvDeHlW1bWD4PVqXGgfcXM928f1OVL14GqjZWzkCU8U6p
slbby/psHJ223kUuLP78VSMUq11fx7NUw+1z6ORrsozhmO5R06Ulsz6BwOJBwK3Q
ItzNWXvP9emJ2WxHOglmNAvX/agGtb8ppQT12FPj0LbU6sBZy3Dr/eMiIW63LYA3
dyZHll7zz5JjxYq/uRNHuYoGwyj10suFomdjHyfxxLC29oOR1CqZsltKGXErYKbh
OaC9k5FY6P2dSSChkq3JjvTRGJ3cLFf+iDttrbNqua3WL6D/yeMxJ2sObMuVnUdT
mAjJScpkPZlncP85YBs6Dh8vcRsYtnbhDWDP0iVqbR9svhwaFRVj8nUOpJ3a/Fg6
TeMO3tfgiXnZnicGfLgQ07YxkG9MWRkgxtAsHLPlr9XUPQrIQz/D2TmHNxYUPt5+
FQ+oNqaGfF/N+TeiCDo6zGyIA0lYwPPn/bL+QLefe1/MFvmag3NXw3tiMBXuvw0V
ZL0nrT86KnUqrUhcJT8x/xU0QnoOhPJmSL8fzP7P0+QIUp2EpPPc31h2gY31vY1w
LnEUbazuT9fM5CYcpwNgQ30DZxmYhQkew+MbCWB3MK0AhKtK+Z8kUZPtaiEtcTTR
IKpJKzPjipdZYuk0otRegXgk3s35Z99th5EH4Zxti68OunLwR78LaNcSp9Hr4Oq/
BZNQSRFQT00zoumBnccvUvrUVOgfhcez1NcDshJsdkmQ8Z2tAVSXLwlvJ35nazBg
RUyprTJ0Fsos8VRfzHBRLcIvw4Azg0qHWrPZRXKbzd8VyYHbJuy4ddCrON1E+rt4
/Hm9lOCa0+Xpd/PysXG3MKm8l06TUbVQg5kFWY8+fhLtF/0VAkPKTYuLozH4odmX
dzyINz/j0k/9042BnB3nM2j6Dfvl9e6H/lG/hQCvVTvhVUZDd1Kk777GJKiE1PD5
HTfCpamdIxLbT3kZTNk6ce+XnIL7XDO99n3Y+ovteep6eR9oFQ0bxYiEC1TLPDLj
Ff87Idz84fXLWnghqG7gqc4lVBh+EBrlY43TsuzhbkqdRtHBKjufIFtzGy6AKjt0
+Ohyyx+Mb80fVMp3RiH7MUmRC9qHy9ZxQwDy1iUnlgVeUselwBEPItxV+AqnuJ5S
PTE7lvfNTcnSk8rQ8kg7CJH4+/ZZADcmEKI90iidGfyqF2kvgCAZGCdawWdLTr4E
VouupmxCUrdIZcV7O0N94FX6vw0wxvcQLlKCOSBzlQfO13hAdnZnEHNyE2pzqvbZ
1wON3tHE8c7TNtrU8jOtYag1/0ZG0hbDvunouqNGWD8K7PWji9rwuNSCPYKO9wgI
JuqI309HhHpGubxWp5pZvZ/DppmVICxeBFSJeKd7xVevWtWBkzGhyLmAHr1bymeU
d9o1bAsNCnVyR96urcm2C0+Q2+onYwMKA05z9f0l2RnHb0qcjtlzAIWv8wHySG8g
eHVSh9fwX793243G5Gn4x887GVVZosZ93OsOAXypzKhEtXoh5b8vGSZvJtT8Nzt8
2gsz4ISnjCleqtlM68qMr8mK7aP500LBAq14BkS/wVRKRDHg5iGAN2PLsI22P0XA
vAfDrP+AgnmwqOITbsc6kTSpMG8rIkne5vjg9WtKADS+f4AzC+KBhJaRvpeo9cDm
pr2BstxQ2th0Tk0uVCDb4T8NA2C04TcMRU1esoUeR50b8ClUFA3eozHHXMGzeHAW
O8qZG9UNfyiHuHbxmbQ9BZlkbdL++RmvWKHfV1YwpGrwe8Sl6rh9Clj0LoGXL8Ea
wm4WpxrSPP2T8yo/VFfIM4PBUjai2rzD+lqN5xqXUCOCqME8OCY3qpEl2BqsFoOL
ZX6x7hfU7m2BWaCkhyzNHDPP2QU+tsy3tYv4fMjHRgmNKRI//TBFTVBChKz6bLdn
1fYuLMG1GC6vNoIfS8Q84zdGNmJQzrIU2f8Je2upi5xLPVYtBD3ZxlReo+m+LP7p
KMXHh733WdCC79T0ndBU6IAiBW+i6pgxUW14KQp9AmPTetJD/R4s0gD6ecNpvyob
BDslVsmVrCWqWVvIY3GBpDUTu8gS2O8axfVGGsgNit6hhT9PKqViI4umwKP0YiPU
+qc/OLOdn4oewN9ruKZ0u2JHlFeUt76zvOjpfcVFlc9NC5uZuG1EhVGGOqTkxt1X
l9aO4AMv7zWLAE3Ck7gzvTpc0NgjRvAVpxc07rnVgfC3In2fxPRKcWEBy3G1lvGx
E6zi/JkkEoPl7BpV995r7tEBLJrKITZqINgUwWYJC2elF+d3YOo4OviW203M+8qw
/Sz72co4TlFCf/9KX7qXoXkzvSACZH7e4Rm/eT042Mw3nmeXIgVPErYt/8ztwxH7
dJijFu7EKdvvgytpYBrovmNRXpZHxNn+SXP5dHWk2Z7EP/Cee1Ue3J1k1IFy1bR3
g2Qwwr0qoSFzosXiLWu35nYS9ht525/Dz2JEZaAsfK4uTr8hXDkU1W5c/XxaJD9t
VsHwAUuYLf1W++A+/NwHcpWpKysTum3AEvTunLcqE+lOljG8qlXyzxvi/ZI9bQnY
LObXVyDxkSNEtoFPVNcDwdQUg0cm/dExqcDdFHgzHLehqrZRJmwDtnnNOirXiI57
1ItDScgNow6NCAgtHyRIrUg+524oHV6roATIp5ab9qEGlfymr95V5Giaih6F73FC
kwNZY2mS/OMpaOld2yznCIf0aaVoYGydkgM/GOKZka1PLX6tfQNsO1uj4I76OscH
KroCXiahig11vTST15tg+k9AqKQWTY9hHSfcKSZx6ljTVC2+fCbOE800v6I9PzB2
WQ2fJ5u4ODLlZyRhzCjBx6QKu2Go/CRANQGb/GpjHPLEJfX6WLJivWu6GqdDKuG4
9qnPkNYtxGku5Ds7t7vlWKVSbAPzUkzRmiqftaXOiZ5tJTe8imGA5Ly7wA4VFy3H
e7eWlR0WCuXJp5+swXv5/ON3JjEOZOIuhg+p0g4INIttUUMtAWjfnNcOD+jdHjm0
bqPFN6htljoZ1Rz/EPHESaSegxEAkz0/M7nwlibi0Fd2TCLnk8A9bZMLL3bgVcVD
TYkIUULfA1UXipFbx2D3pguqZpQr+vivQcxdhQ7bqJpJJSQSVZmUmFgIjIsarLAg
Z+tJJXBL1eTIYOsqaxzkCOmuy61ut5ih3j8eevGPAk38xmtkjJOnVz+7k09VMtt8
sSRwdc5rE6qBh319CnIFIcCRNgjQAOoemr8wEDIPbjXyPlI2UipCDcbLiyjgj/XY
AETGf0K/uMxUMM+Y4snUMe38OWjSYAlBkhfLpVlS20zZ2vclko6bHSifkLJaWzIO
Ep97wYtCKCIJ0OG7VODcrtZLF21wDZMPlXMPLVVWPjlpwmAgmmA5s4D2QIcAPLy8
A6+U7YT/QCORLv4tXIvfS3v1gN320a/9Ic4YunEZcPQWQ8wAZcmSZH36yOQA9vgq
VRNkJZuF6M7swG03s2rxFjG7Elz0UQd14YW41l2b6bxAVS4Brwo49/0XI/oE9rwH
rCzJwwwCzQVocQ7nSJEelGcXV2dqqak5yLKz6/bUTI2eOurMO1L/IL9htP/PLYc/
dN0MNeZvQOgiD0MGDCO/ozB6GEc54383/6DuGb3YKhzJRo8Ng4bnDyiurRA1yBDt
Kl7oUiS1HvGvRvVFRmogAyBj4O0imH3LvlFyIt3OmDNyy9G3EkUDmkiG3paXpVny
QXAf5KDUpcX61lrhi4lZCMAYFCj5JxzPV2zb6Z56feULWwPRQqjBgB7m2lY/vRRx
whg7Mpu/F2uRTn9cu6WnOks49Q21qABOyP+V3BHpgNTJVGydFelkIfpwlGo5KL2v
aOslfMy5k7ZVd4Yq8odslueY6Dps7RSkO4ClmzEGhzMGHRfNlofUhSSKJQljJG/T
KUDydnEExnHyZ+s7Ys6zB5zFeb7fWWGJ4j3rgzBjE2huHB4FQDH3oJvxToTaP0vK
aGXMw+M9EqpeFHEzOJjCjW1eJ9CzqPfoOfVv8yyJeIL/hd0JptksKw30lDOSgvz2
l0QOn+uKcIVb+nQKxZOfir+bTASfBJmz5dC9CoBtWMw5WWqfXS5Jal8dOWB54Vm+
3Twbaj+dxRlTINhK8flWFALzxGIPDcAzungI6WLbRTRmvdgkhdzAVcGSSWjSZR4T
CnDE9wRORWCUkVYqsO7TKJoMxY3em+JfuovPyUZdU+1U4Rrz6XfYtnXKj09vKv6E
FbFLcgsXv3vMsRv9+8V2DJCb2FSI/GDhpRofaou+7CLhB8W18G3ZEA4yCHvIW7I6
BWWavfYj8qV3OmhvYXKcFPzPtJ/+ayipNqL7VdYlPXjKz/QueQJ9+6OW1A1mKI9J
LPskdob7elPqyhC7ROa6QOJG0wwTTNLg1iqhdQAe+1VYJP5PgqF0oi6XnuW1wL/R
rGzpqjSZ17AdaehQ5aT0eU6xdrPzkP6w+i421e94OvXaHDZjxgPvU2mxHKXha1iy
4pf6DU/Tv9DDRk4Woe3djz8TDdnaJ535w+t1e71TksQl441ETssPgjU21dvUDITS
FWSElZ0DT7lylmu3ZgSHNL6iNmzWK8FgVPEkBk1ABy3spq2Otd00+zGTDjH/inRG
DCHeQssUBBXNWEbuIPsXd/3ukzn3ps1Dw/K7TyH0Bxa2D9HXqbmjQ3W30MEUjptQ
pI9J8XuYvq/Blx5mKLvZaHXTzaXUe37qOaOz9bNB/HKa60TbgWtD1u5FJWYRQ6g+
2Hd58Vzm/SOWApi3XHpGsup2ZZEq6Jpfv/If5i2tIi0iq+jQRqwsk6MZ0dIfGHhc
dY5HkGTTxbk+UuTqX9CDRvzi2G0pObBatbxx8kkugSDd4h+0I4CLqyp0QExHnDbu
q1gBa1iIOgHnTXRF+HZdGKR5+L+E7NtGZiwnFbuV5fziZ3kvkGUWMqL8ua6wkfmT
4Aqt21p3W3zpoQhGfcBkcvqvCKaOJlGiPV3dUt5gJVc8+6fwZqvS+7jJ3z2atNEB
rE6Z5qJ8mS0rENrh7jbtmR4ZRpirTTXeaPnNjE9sfw6X4VH0NfXXyPgzAuF3R3SH
lvaHRqrDuH8zCdSQZZH/YO8VPC+L5CyCgcXiqtVpzWP/0PsjaG6jKuMWY/G9QjQX
GOViOjyc5fBnxdvjWNoYPu4pt+fOyhKlGXlNJtxc00mn4TRqNwDdpCELJuwKLajE
anf+bDd5v1hSjYh5lzur7v3NJRXSfwn8dKckNqeioA+fxj0WiyPgHC/gkd93g4Un
XCEpTM2NKav6M7lpqiLxJ4EdJ8ZVamj+d3rRy33bYvRSzWqF9tfIjIZ3nsiIK0Q3
3xyrY/EHSX4kqS5ErblkgUozJxt9f5mNOX9BB3BMMK7SR3z6wJqsSP7lIZ/juyxc
te8zl0pUgpbHai9U0ZZIqx+rNLG1wuQU4ZHYS6sWRMmm6//CVM1fjoS7zDmzQxH0
9h5w0xoO3Ywnh431mnPQagx/SVycthb+LQGB12a8wvxF4z2P+Aq4D45hrY9uj2gF
RJgEE7zJfpLSyiz4eKIvvxTvrwfqqA3Q69/alMfbFvMcXAP7ky5D0ZNWCpHwIdCJ
tg8gbNTxquDZJYdTtAAV8TPFnxdoY7Sc0s1RxSK7aidJEg7eXqJhGG6T0leTBjMd
R0M+ao+54fCTLkDxKH7Fq00L3y9kWgG9q67XYnUOnQm78dGRkh+9hSKQX+Jo2YsY
q6/wRi6RZIlB/A3+LnQ3VZXl9s3WAcifI3Fs8mAixMiOgSrs/4Q2IrrfMza8xgvj
1CrM/pRdT3T4/IYWHozIo9xRfMkqCRfxJMVeV63Qis+CWjWNhVybpzYOP1w9EQ6Z
kO8SymCkrUFbxDhcpxdxaEvestKeqULQR5qJnUSg4R+r742spJU0kqDCC6gkTwDd
volr+uec/wpHvRO/Ygd9/CLnOzFnglWN1vtLTGZbnpJik6HF+QKZxaTOvdACVCTm
m7SxWcmEN22am2dSIK0K3572srpydNCcBW/AgZN2Fjl2FH/hBz5MIebnMcAqn4gF
pR4NRWhSbaAjYaKNXEI4oonkc6R/ZT4PvkhsUi1wcM33OjJyGCnQfsojQkEyoWRx
meTes8HVXNWAEo90eT1yhsm36rgloCSPuLybEDPAtNq4ixE87cqeMyt8xLMIrfv3
ic2qFjKBmbpNjsQeZFbGAU6XTyGs2Ppy/GN8Kjjn8gLA411IIeFsNswH333FPbIu
b70QWVDLF0ELWOMCLbhxJPXWiSsqFJPnzi/1iCgdF7XoR3R0MgQEdZu/SgoEyjw6
oqLkJHn8qSsBU3+Sk2OYWj5K0p8/RF1JTFd9VDy7mDrw/8AjVk5z1ie5u8Vds52C
LplPiVPvXQBLqmfiXl8YqMy3M3TdnYMv8gDqLzVzrIsYD+H02O7CrvrcdmscaFN3
UdPHuDIZyQceKIbEUua7B6jVh2wwk9EUT3qTFVqdRSA41M1gr7N8m9DPbnDe89wB
KDX93h+AfQfDQeUqFAzD5dGxYxVZTTQgXaCSPSE7r+8PVYmkQdsEu+F4deLZzURl
U4HETAgL3770iqXu/5yY/0/xuE7EgoxQYAN6/i7/XEB/nj0ua4Mv6huPqZ1JHRES
44rOz/b51iXE+UHAp2A0AoOcT401lJCtHineY0kpgpCIb5vYW+eIPgY++jr3+kQ0
9Rla6JW5frYRR2dbBAW157lAF2KxJwVEgTpXI+c3yQnES90HFc8BW7APe7fP6Rdt
Cshc0nND7Cq2l0gJfEP13iNnkDSOuWY3cja/cbtSnSTxD5ojGJFWRMF/q3LnHDjO
7wM4LCGksWasnIO6Dg7R+Y0MS2wuk8vSvJul0f0cT3y2tt8SjOZl5OqReE1xQrvj
JnxtrTdGMC5pHiwhVz83skCAv3cXaDelFmgSuh/XjxHw+3eqUL2wYJu9TKnzc+Op
wbivDrMB8Y762WzsrJ+n41PWtMmLVsjEax7edd7Y5ctvy4NZFyV1iNSWR2Zvw38P
AKXiwO2gukL6fd4NTnbL6ms37WcZwgTR+PIEvfPYjLayHNd7j2UHl2AhtTU+HaJl
im/rOQJxmmZwykWET2z8ju+bd9sKtdjfoQr7uJXqSRSCbgdfApsEHiMz0w7ZqmSY
bVu5aStNrwqNNAkK2n1QEogTjrrYszxgoACXHdODDFZzWvRVyJ3ysqzKJWgcLEDy
nq83cGd9dTsVEnLOhL/6Z7fKsa6XCAu/XPnzjSANWvyDsTif+Dj5xnCS5Jm2qblS
+dJ0lm5erlHnrG95HKTXFqZHfPgFQTJHR/TX4G5TdqlqcQn6Hh5BOVPJRcsk67bi
FAs98+Ob3bJFTOgpPcHWFzaSY55M+pCVQes+9o5GWIoC7KZ7cWEhI1nabjyj7kIG
+bsMBMTo2byq0dcupIo9+ZuVqziH7EUnfO1Viko/UYNJvtSnuMHj0kprQGVFxNBS
vG+MaAFvwnWPz5XgXFy3t7ogVRxwdCiMCX4Ocu0JYCCscmx6QmAZDFkWSt+K8O8Q
tl/GutSKxTGbvniASFeEMja63G6N8d7/X+AjLlqnOcbF/JQ59z+BMHvnYOfaSoZD
QK7m2kAbswM996WZZCD8RFEiCwrUlZb2gNLBeJyjZ22iROJWYkK1bTWt0CfF9fzo
BVtOLT2ltOelDYnDnUJQWIBguRzVxruwRhDY2tE8UubK93+2OMCl/001l9veY4CB
2dmA9Lk3peAosIxAMfNJSUnZuKivshPKciAUWCJgeIRTKG8EzrcijQMhPs6odhXL
pJuEv5zzPnyrsV/IbTvX4/nPQCWRt9qYngwpZvusYMZVwMEzO+jRDa7gB//+UjlR
BpqJzcwPi6iB1RIx66wGFxBkzaQRoL5pGWiI9TD3PIIXjcK4hPfajU295i9NnlDj
sSBbCa4ed1s9iMYWVEJtyxMngAPVANzIrK+AzVAKCxaoW7AJyWHZYoVTmca9aHVs
EiR+h49oTmxVCD84UV+OHHcJp37JW3X38V/ncTDM91Z7ZStD8IOVCjsKnO7UTGWL
0et+GwPwri6hN3wscR7jgInWmS6/2ImllQnvCPffVxCrnN2t7reX2D1SVk7LZIRF
SfjXjsYaq06HgRfA5PbYVU5lUu6QFdoI+r+0qG6y8NPeqw1V6LhLWrnp6XyqunSX
tS3wMnEqsmWFZSobxVXT1G3K98GhKICWuBYaeYaSvXzNoU8cluWMQEWZKTl5EtAj
fOAzc/xGAz2xuUdJ005kH304GQDx6SLF4QpnEUh6WnJn8UZR1GS75A90RsM1laGU
saQu7FUfk0NTiPwxkizxD54DhyNCSx8N7s2fitk6v47yAFK46sSMYnj7lOfNmWPp
VpLGDVfbXPV1z/XGN4jmwcEC7R6bVeRGVXnIIRRrfiX6MpaPVjY4Gr7gytVoZnzA
cl7pGVctjauet7mnW/SxT2ZaJ3Jf7EG+O7ZD5uYBHs84OZVwIkq2QzPjIoRgIYKa
Qh2zpSBXi/DekHDvgw4SXnX+lWqHNmqupwkZj+r4IIRbZWp8THb1UDSmTXSnaiFu
3GCJhwO0jX8JpHpgv7EGUc3gPOV3+J7H/iSf2HZDaLVK5sZRH9EIx6LHoVYRJHuw
9Lz2Ks49nYnT52aMGfFRc3mbjJaYpTIafG/d6LdnxnM8sPPcALKnjMPfBtHgAq2q
3J1eyzkONEK0w/8TuV4MEwo7uTYFx0ZFeLww0r4ZWXhCz49XS/CKq7Q2aac1Iryh
fWbhmjxYuj6TeX/dpvwSICEEpMLmKNVQQ6S/hvtZQ1IgQJ16lO/kTy5hXv9LQKyS
S90n4XJoig5/XU5t5xA9ffRrRkaqxHv0X/nr7yioWINOyisCp6OlWZkBe8Q8758V
3ZFhA2++/oNgtEuM+5xlMlrlau6Y1rji7hpt0IAy107n1/jmu+ktPdN3ySmeVp5D
v5xJWhVYnoPucjF93KxbO9vrWz9XbM6yxm/j6HDxEFDVyzE1GITzLErBqJqyc5ie
r3CPJbNgrmRY7gtUs0cWoyRJQh4Az0G0b4il5tMPJSTmG1/44Iojo/ZgDGVm9aKQ
umArvDUSi2bcfk5CB8PDT9rxSN/+4+hj74C89UteXKQxstUT42Zyf8PJZmm9uXSz
Nyg2omu2g5qlNA/mdMmmdymWwwMgrvifAhqUKaKaozp9olSztzJOULP1gdgBjUB2
NjZcenUlSQceQo5eL6KaMtjdxAwqOGbrmZvk1T0dqYK5BKJfl2pmVUXQN/M7Pm06
qgRu7LV6ojcET8ntWK/YlJ2P0OaNNgoeK9pvdgY63tNL2hBF6Qz1us9smCxetnOM
6p6rrm/guBwjP1RioUo+JI66BRHFCn36oq0UvEuzhsEaMEJeKaY4Fky8HVID2ebY
+ltVHKEFuEqaGn7qCkmbEAiEUWWAE5MRFN+dIaRYnWYaXBYNxdYB6FiH3It9iPgK
FKMub/muk3bI9wDAbkB8kDmulFFmSlIPDq21v9MUGNRZJD4+cWJFB7STO4+Z2Iyf
DWIkIZ4Chq57KneEr43i9Sou+1Y3cAG01qqqSZN0uziTUwWW7D0uzgBSH80zavCj
0ChicDwzSPLCfdL8K8uLz39r2nyCGIewTvd0jHJoTHiosLw7mLl3G4lCcTnQLK/N
+4rT+Y7coHGw/QDl9GGewPRZWeugFq2dkkeMT+Gvg+PB+6aq6pnsM/N2373JDo6A
SC1r2Z3+nP1MT3LCAr/3b7A6yGRCt8PXAN+gioDWyIx9LsPhfB6ptlm3ugHZXDzX
Q0bxuypRgdiUuP2PrJDa6wDyfmwvXBE0MmKw4nx2XysZrbUK72a9ipBXU0pxe7DJ
eFvH/kpHznAuzvhkD3Zlbt/PETSJkimy8flSeCW8pH2+eBqFHEnTVQKUD+TDMYAS
9FFnkvUlGJdK9jZcrou0VOWfNt5Snt/68dbkQy7nvhDO/F5t/wwmHVfNMpb0D0No
WSK6o84VOa6RGlvauaGfQbTWUmUIhAdkImlVAglfFPVBheFhpkSXDAucLlXmO7A6
zbiomhP4vJ77j/1DGmSDTm0987SG1/Y6lE/Nk5TuSMer1LkqB7OOit39rMX8OnDa
NUL26KZjh/6q7cP4W4W5B6E+TBZx6GfymVyT6c3XkX02dc/SSjmQO4Y47F9bzwEn
5aFo3QY4bAt1ucNt6TSLhayD0nX8F+Ak5zjxkdadcT4BwpKdmGVoyeFs2vMQCtMx
KbQd6rrHakbX5ihYjtVzGAwrrPnd0nPm1XJyQH525Efs5vjizZdTGa7MiCZ00rIj
Bm08irrRjMIx2L50pM494SuC04/LJ1QigLK5+0JtAHarr8v8aEyEjBL6EKl+yUxd
aZ7jXEy9SI93X7zg2HdRh171dhl4ltS21eAIfD++xC9TccQECAnDhSwOwC+IUbce
5NMy57nc8Y6y76FXreU3e5NMHXttsLyCT7nwvphSzV3h3IFM6PprfauZ9+t9mwF2
Rdd2AyZ0zQdocB/uog+DTRyOxZDyLody6Zqv/dh/x/fDssn+3Gbew+WJknbi9Bth
DnjFji7FNcaKgpzeeeldpgejzQIbTRlyYwe2/ZLvlO+65JRM4GTuwh0nmDfpLEMZ
oJKcSrn0ehwGzyTBoVKzTd9frApEgfYqEgQACaY5Yf87Cgdhliro78yXDOCMtGeA
uB6fS49WPxZSCVK/DeWCYBzz3gkwQuBSssHcBLCq0T7wYGl0CgQnDkDKI6KipWRw
4zYGRUzk3SJ019zYKg0wdYmxBEbHbaVN/d5Ncq+H/F/QmfIBnykua/B+BYR7D6Su
1CXVmEooFHPQg6cY7VrwFeAPAYxXzLL9yW1yvVoWl6r+f0ymJa1BrhZ9luqyWjEz
QBpNIcQWX8hvuVNZejPMEvV1GM95GAmiPuKO3tNW4J92TYkAWwx5hRGK4ffH4vom
HPxeI946d0f5CnpPMJ2Y/T1K48wL2k1bBoQhEblUzn1qh+SJeHndXTu7lXuDFZSC
ILdVVz1BE6Saav5YXo0EeSsrBpMeTqSdITNwbPA2+4TMchpPRgQ1/VzdsAtzzzDe
arLJlxBHJiNsLH6PNvkBrdq0sv8iIlPHv0yUlZHlD9+72IupnXq0/m9WjyoURvg/
8qxdCJqxeZVH/ZMyWuIshXJNSfkqOxxZuQOMQSBkTPsK3PaUALdQn/F5muqOMQIi
1IGzJih0qK1hs2HEM2IqCCg15wnp9SMhCcvtbPyfLuOkUW0hioND5h3jCuiseRIs
Rlo5fD/ylv3ZORHs5B4cOoo1iEMxgoIFXTPGU/y2z9mJA4Zz6u50kIC2GnMucc9Y
vp2chsHT5D2N8EkrVe50WhBq0VNa8xLqYLylV5RVMiJgRFZU139z3TEJhltI+thW
Gu2iYixejXKxOceqLvZBzgngDlk0YEUM5K4Ndtde5GwJ5lIgQe3E14NdwUcrcvg0
pfCasREJhcp5+FKd2Fv/cPX/BVCE6XGObCfh0fDRq6+HO/Q0SGNe9PoDXtRYP/yH
V7MIIUbuIpV2XmV8E8sztAIDAArCg7aTBRjwiP4lOopcr1vMD4Lf1HrVMz6bD7Bt
bmjpLKKtoglM++z5DPsgg1ieBhDqvi8OKZDdCVM47gtmwqrDuADsXWjIuTEi9eax
oT9rXRiwFFrV30I76O2gZaxVh1VNB3uymcubO4PO+nGXlF+nQlF+SevrxK4grMDk
EDOZWByzWq53m3JDmKJYVpce2lh3v42Jpdj5+AvN5aD1yye+YNspFxVxhoNlLn6C
Vc9VLunT/4tSbHU/UBLsMQnH2BV7/1vvc1GwDNZwNzuSv0gn1k5liiS8OysGzaxJ
9YEySbM0tsqatA2K1SdXHIReVW94UQfwyxmHDZY8BcW3UWE7BGwEQa0gfoGzHFS5
eRcLxun72whk7WmwQ2Ktzmmf+sc1YUIXbxSlcJruuUXKDLIWjYTTlCGHyZyRX3TN
nmCBz8xI7NpjRDXAIBe5uX32EaPUWzJ9gImK5f9zL9UzoHdhQm2tfKw+QbMzZGtx
mbMoy+u8kuMlHaPh2ZIwSky75UN5XYghXRhlkdw/H7eT17AtofGppYzCd/PgRcku
k2xPbdkuG23az0wKV0lUDJxawRTMvR7uBWhXiHfTyVwDcWCBdKsdOZbtIudNALnd
FziBf0O5TLcKWSBgbNATdTyarUJbGNj/47img8bF7ssWAX1vRGv/bWSrKtjrng11
5B6bBOCMLgwnnMG2cY9UdYkHAZ5PsoW8T5OkfeyfZVKig2/NXo9lnlYK3Wg+4yWn
6PmQ/+bIDMqN1uvdBITA9+OY27GA1Rmy/eFldfiMKOUL4VoeQOZK4eKwJe6Iwo1m
CkXBzUJhFB9ya+IUhcQxi5NLTcy8NZMrnm6Gl0eXTe1XPg1M+NeIPlgBLU6Ywtea
+YDpKdgPes6asAW5NNrVe1gWbRhgHU5p7L55qJkQUeyd5WAXN5TWhJtyeIaKD6hd
frN385ywGR1cGoDOx8/oLEU0pz3GgbypI0JRrYtqky0q9RwBcAN9MeDpfT3gjc1h
gNFrdawG1EjmDPJL06QUJGH2Vns+ahZ5J8TXCnGa/ZNLkHszaypWyjaX3KLXBEmH
HaL1RqJal9XgoyQHgbs76eUIYqEwbMTSwYgu1s5DWkK2SKq1dYCOz4quHn6lTL0e
wZNygjKF0qp4AlWU0WRvwaLb6RtvWV8vOPuKzRO+8T8aWrn3jxXIPa7tHfG9Kpqy
BeCVwO7CNWbrt1K2l+GcNItZfbRhBXrSedNY/gQvIt74VhT7LvcoukqmBVrXCWEy
GdgY7tSjOeyvKaV5sYoNJQXaG4qjA6H36d+niV9iyIGHoCWXFo4kQfJN+a1oNo+I
kXfek2TuD8nMJIAEAIurF71oNvelD8AMUuCKI2Sm1NdRMv0Z/OOxfxaz5dtrmdli
sbTOf6iICd2aou3T2W9LEmaAcOi7IKVU1SZMmbdrvIbKPNvZp9qv+9Q8t+t6ctVE
P/SugEtucROXeYta6MJWWQE+7coaxHF8XjUKI6qDgbeg5JKmfE2vpim0lScwC0Qw
Mdo6e1JP06dJYHwDp1ScYEQvTpndcRhVqktJkiBWE1KvvaXNyPXexU+QrPe2hcwn
FF+XjNky63EjP2xw+cw6lrEZoIaH141wjUtCDzb8XYmP+rrSAfwMVwsT2g6lhuFm
IDibNGWRF596G5Z/0Xers4VXPRKfJdJtKdn7xKlcdZjjs6kb3yaYwdTomDj7Vplq
er1dkL93G7p+0LVVEr6dOQeaEtVAGnzUpIXWjTpKS0i77YOfAdGxAqPuOa2G2dZb
V+yvu5rO+Sfos6qWA0mHUFUjsl2njkK1n9E4LV7hvpfYjHcVTG5OjApokiMyg3Pg
fdc+sWIhHmNVCQZgu+nYnrzvKFQGe3wBe9ySLKCUmnvNERBmpJBKnIheKJBTbxwM
Sh4zOX56EKGQwxjNw36Taa0U/o/qQQuFgqhM/KFMOXBXAViDeKJGQeqqVqrTnICO
EuW5ip0kgK5jvNOdXrK0WPmKe6m3wW8wQFyfhwizRU2WDoKQhagLSuCkK+JkRcok
XUORfGR6g8INu1mzqvJNPYBGMqN5lmu/Jyxhqal0/bX8yjn2hKLneJeubbTnyxQt
5Dxd6WgbEpLJxxm7HhCw0zNtnQ6Z3SQPccbgXUElM319QFtdUdITS8zrnMvx4Wry
0ToeEguuYaoHriWqn6uSe7JyYSProGW9NgGz7pJE/phg+C7JDprg+/7GQ3GrYDWp
ppNlFYoBEKXSzaDzuR5FeK6vOxxPyDvHBF88L9Z6T9momg6OBUeF8LQG3EbAroVb
zIhjpcb7LXzopXsEitE8zFAUXLaAmTOwHsia/gx5psnNANeYMLUgBY4pXKoq9XWc
H1Cb3QLth2KRxVm/+ZSBSroSShPgZzs2a/CeHyqlOGTh/p9JC1pXLSF1FCd2m+Kq
R5Ftwx3FereQW7wKkdtkNdStLAaczm0aOFPNOslyLQmp+2kRiPWsOagjIJMeIp6E
F67e4F3OdBueGsk2C1upRkhBngSxfc/H8+a8GX+U28PuFL3txtcH8tILAx7VXYTz
yuHtXgbfeWkqfgGttKWG/gvzP+oAtiil7XfZLjKoj7+yBTzJ+z9J0aoYslkI2r1J
K+pHefZkKWzYb5qAlKaroNwq+Xvx6XJHqigIk3pgFlUcJrDkvASk7q1jR5wssjUl
t+mohqKJL9VJekyeyXrJhbb2oTuM4PV+EOxLA3Jlbk2CDKBbxi3WNKuNWA4wiaFE
qaJuIKjFIbmGd96cxpNUm6iBgoBr+6Kk/3jFIx8zVoi48B9zqDmbKeUCOht06HXe
RBl+aUAMekgFCygctRYWvyVBBQIKxjjwpUC1UjElSzmHia8h0yue5jS0Cd4+HpKH
H0oCkH/jN039k6jgL7gmSXykF7TJbdHPYVGVdD3NjiMLq/u0+tOxeMXvRjFP1De4
iKdyqcv0zM8JmZAnfb7Pbe7RxZCMOIwLlAN5BrlIE5FpMgQKCDRNZem9cYhXtd3C
D7UQLUvp5xIckTjtMvEPd0JH1ss+JEodpS8BIhOMn0AbpyZoaxdgeQdjmMSjCQjP
FKiky2+3FS/+q7yzdB0vdK5e3Aqj2Km70z/ckBBStDbwEVd56ZEZ4Un+zpMoSi1f
70LeLIGhgIHPQb3m0ECzd0hq/O7uEHwX0W4suoXAHZvuscQtLYW4cBVy9K1bLG2r
dw/ePpNitiXD8ZsxVPrt7HfUqV3JsJHMgVw2sFAffD/6Su+E8PBdG9SVkxk2DB/W
ZtJnhN931njkNxtWQlFt7ZcGS0fpD5DdfrSLSCQC0iwmHD77mfYO8q0wXFydYBJN
AbThFGFCOeelhLjQZcLKaD0Mi4CWFxwGfFbZIDb/5tMZrUokacp2VHUwuS04ZR/2
75+VHOR4S3UAg1bLw4wD+xtyVocTq3VhMPb8unaQt4gxfWxLppdJtUG9tMMAWNP6
0GMofikWEK4NlsUsP0xE+5i+4tyx5YvkElh7weGr9lUTdUQ8czo6Uz4uaZ9yeUeb
kMIWOEuQr58yv/OKdOcNgYoxEqVGzSg755JGjPOPgVlZoXrPh2NYqgkvUBqC+xlf
BVUU985YLw5zWeRUNoUpdFkhYTNvvJrnpyDg+lvyPcLwBMtjZWkOWkoucfbca1Ws
89mUZpuGOZbwUxCIvgcTtoLRXuTCSwZsClW9BSFGlGfHz7lk1LpRHsD37FPXZ4SJ
djrMvzdCzWx4gtraniJ5f8Y1Bz80liMt7QSlmeeHLLYt1WEAYnRSz/6V8kq5r02t
yVbDA44eJMyWofNTK4lcqIzm4t+dwiS8zuHEi7Rd4Ep+o0+H6LMvhJeUftPIii42
3lSGW3CREonTyTkXgFE7o+6dS71R0t7p0OGJwxGjVTTssIKZNaAcDyuWpy1mbIxn
ASWG/3IBjkYpSonctnia4c3IBlt55vNSulcdJvtBMK7HlP9+xXCnsC9hm81dQXL5
qRnSRbXDXW11W8VrcTZVbGjtnkxbwpz3Yr6vxKbiFYqntE4JCki7sg+qpudgpSXn
z7dlXAj6bnUSs7k4k7PuC+mvJkOS26ttfDRhBL0Qt6giVKEyPfVoE6d2jWS2krpx
yzVDsDAmSavbzmJqSKDLtfuQSyxkvzTQZMaeeVxxborJPl/2rMDGeWmqLnn1InsG
U8hAjEw0A0ASvHv84VtFjJcKTGn00UDknYg3uun1Qo7baLByIDD1w/902nXaXxFl
ICPRLX26meTKLbY/6GO/DbFSGsrzG2rcf+sQ1A46Lse+cSZi31tbOBrGA7eKSOjj
C6pl7zGYJ/gpx4h9ENH9PBemuRtNJ14ybCk2ad9mM1X40XSi8q0n4Cbb/ZYxvDzm
bVGxex7AzvJ+9qDt/K6QZAugt1yAjLBd7nAEqjUbbVJFlB/3E2gaL864ywS3IzRO
hk9G6Tw9E1jQXG0FG/X6Ewl0yMP9njNXpD8jFpuMsbnzInVqvchRByrRBijgw9Nk
ix6yj4Oj911WXBapXxI7k9iW94EjXgRKknYLN+7HsGPh3DdBdfaBeNDjbF3WIggC
i7tb+UiVs9njWBgWQap7NIDPiA7atn2JxPElLXwU4xP7cvPY6aHWjvGeVH3W1HLV
D3Skd5/BatbFb1Pvg9GBdNnRPP4qhiviQOdRd25k5oRNzlVPiDpbngK89w1wCBFG
1vGYTEqW57kHbS6+GKnOp/Hgzc3pjkuBsJUSVhg4Rl2Iw54Xl3KuVdoyBEP9Xn8B
+nVvdy7xGsKCh5vYZtgIoKR0+U3lK2YM87o3fl2UwJH+QHfRbV3whR4Wz9M4ubU3
/mEdQOodZNh/euq0gYXs6P9xRjkf7AE9yMo3PaKbt3s5gtPNh0AXrHYiEaEvJL53
UUwVbEa1XSA3BLi8vQ1IlR7Dj5qGxdLn6RdKSI5v/A6W3GxH2gHm1Tusv9qT3WLz
nGI7PZRO1xmU/Qxh2CdoncuheM1gy3AO0KbKATy7EZLC/ZkaVzR1DO7msd+0ZexV
2QHhH4X2QAU4Fj9KlQe/rltbmj16XLvfchI/TkezvQch7+9+MdtP5ympmjW+YN09
pPvQyWg9dbI8Jc5KJl+ez4NzavrDhRzwDc3tQHafIuhqXCp7hpuBrbzC3tLQ1ubX
KnrtCXgRbzByzYBkOX5hZ8CymhNtvQ6tooQ9EYGSIas0dz/qG/OhdjwQHX1c2qa3
S0vq/QVNsNb5+5+WC3PpHiCKUNCM1eVHHP+RSPI33D+dIMIfoKC+ambu2nOBoBGl
2ngEMtbqlMxhLpax5ShGCaunPn+QKLn2yFnJivkn3136qL0DDQlS2OJ36iJ5DnZG
Qv2e/mkW8ljiWp8eirFoJXUas1Diyd79BxEvGH/Ja+htgnqUn3mTHROo0NJ7KAEh
Tr8A+dqanJ4+dg+XpsKQGVXnownJ+8lpS+Nb9UyskR5eTDMECcLG0w3CFO6or2+7
Yvx1S8fzFBpzt9Y0losa4L4AjpTGKEWNTZl0/tpkBI/JyeNv/yV6EXBP/qb4l+JX
gzEG3qkisuC2TBjS0mY1eZv5EOrc8noYShEw+P5B+dsvR86Zm7//1mK7fCWxDx6+
/DAMDLypDMM2EMdk42pxbJJn5B8mzg5+WfUsq0/kwTeCEMbFdeYFRgQGtmmEYazM
H7Qt+vPGeGOHaKOjsPyVy79UmKG/zkasr4/yLFWXjhYmKvexxgi2mJlurqxDvM4r
nn+5fF7rRDDcoJ5a60QK5AoquZ8aDFRLoN4sev+ExFvF/bOZBRcpbrN2jR5zDUJI
n4y0UUNZTRj3tq7PGbboTwoamEORaFTun60PzUY6nHlHZr/pupKd/LdnWeuGbO1r
L3ppAVppHEchRbwVaC1Q+UFr6NXNyb6KKfb/wg8rhNk5PBc2nMtEq4QfA5eI223a
rTYguqAQn7nDjusvb2J353U4IOHYThOn3RrnlyyVbR17Wh3l2tUlz4DGaiDSu0NP
1pq6GMLg4LsW1ggm40N7KorO+CN3KCzO3Qz2WuPz94+tZelD63Jlg85cBYtB9EQ8
RRBbjOMzE+qaaogk6lH83J3DON59Ra3XeHC8hFi0T9OESNtMIrMjKV8w7BqLG5QG
WGhOMHv8D/t2VsiIbBF+84zBgQuOTXzeLT8pzIu/Y+oZgUaHSuCsLm7274y1MDmF
hbFiOcgacRlD9OWPwDpB0vDkmOpzN6giPjekLYfXKueSoLGfwteAY6KQXukNFoKs
YHaSYkQY43OHCbrfEovZf/uwLIw2IOMVh45nAsilbNEXKDa0HiHOo+1mZiRqHTk4
asbJRrw5ynveXsh4K/XgwRWvVvctFTVYKbunuAI7oDym6fLURmPN40BgWvWSzDWS
3yUvO6T/4sXAaZHy8UScH54MIQnHfAY0oJC7mJgTK+HR44/7P7ck1xkEhOz3ZPFd
oSPzvobrOQabJCgPiIgBZX+eXKyoZXJjvpqHSLBKiIR2rHPUdhulT91agTTkZalt
UuTotk4em1NDX2rSb3TPAbItGbbDqAJQgbE1vroGIV4nQrvAxelJjZEbkJ2EV49e
ac+hO93bRnJCjqJvSK6TyA4h4N2ELAy83WQA4sTCGWG534opwqjLyL496WHPp8t1
+avsKK0tRPZalHCUm1QL83wTRjZqqvEEXUiI2ycNicJxQRV8QEw7siLn3cvyCKIp
z51YV+tHwzxLd2m2bsceepEQsi9OnJs8phrq3qZRxnAMtwbFE+hpTPAij8yCHEWY
sR4YVvJJtMGlowTGTDnbIGn8w2c5hH02Hvmd/uj7T1gHWtR2R36YyY2bJgr47HZr
9Ginaxp4WIb+oQnp1Sfk3mavhF3VLu2sMsX6xTRGTMSGCy05gY405GKx4B1KVF2x
3aAxDLmK2GZt4/2KwYqDMQCQq+zo6hl7JLBlFqDlshGbjpnNKLtA4+RDynj15jD6
AL+TuZXk+sjwH062wwZZdoxbDVIdepisjfzSbJXLuVMInyk6ctwvU2ZRPxUY6Jk4
IJxdIgCiuNDSnQSdgHMZGCLRZdUtKWouDcXGbd1Q/LNnFNA6rzPRV8UgWhJG3Upx
fpx4VxNOfaPJHkEgDQR/F5sxO2PRN7pDyPLYk9fY5FiiGD7vdOVIT1y8Is+jHIHq
6dnCjoCjLPHl27yyWmV8gComKdCpXpT1Ca4NEisB2MaZdXi7LV60fcQWR9s1Kz4T
cRXB1L78ycZPt5xJKJI+VXpjCPv3izh/ocJE1/wZtVPWo1OKd8W3qK+gGmJ3Qvsr
g5KOXvxbr22daA5KMhHjOW8e+2zZfLm4pG8IG7FpIMmsvn5j0VsvyoF1EZQLvj6S
lnJMdlwYJ0ynkhOmNnOAtdjk/TcXzoWF8LNz6gjPG6S6besn5tGkzK1w0UYUmonh
TgP8lky2qSQAcsPXutsJFFvIo/3d0OAdv3kkbjZgnVFt+1UKU8+e0qy9uV6M8OBd
Ohl7jwVaOPhKT/caVYb52Kx7TqZ18RyYYQI+lTxTMOUBMML9BF2WppxJrwcmCCOL
fFhhFeYx3nMNKdpdUp02BWL25Uc+gC6eL/0k/0snOHdeuEDlR8qZDl30RSETdi6q
bdeBu76HuRFKQ+1lUgn6UKadir+kJO1N8Np97lzIjx7ZVh+4OTql8IN+RhqooA3j
XngT/3uigvmQsOIDnUIhMQU3R0x3bDXLJrUnLh4dz2BzVqCdKaCpw77pTKLQsG8d
3dI41iF5iUzdkzznGgzlpl8BX+m0vqkSirdLLDlylkWp4gmR9KSNuBjI2Ddna23j
f1RL27DmndKzvxLG48QkD0rFxHDShFYjyeto20IpL4D5xdcQlwdDPg7nuduYKMLJ
Vh2/72X52Rx9BEZP8jngKqitvObBEtApdcxj67KLS6TSuhxSNs2oCsmqcmiilfiq
IWrruoriWEj8gTtNqhrRks+nw/9Sdr0FQc7eg+brwAUzR+yL/Q/ZE7v5bRMTrV8T
Hurx8SxbnGIoAkSAwAFM50P6oWaE9a2stCYu0HewXsJ29ONlR3uhslEarJN2cZzq
4icwzlcBHcgM/9Y0ZlgkskTfBxfktW2PsbIwAm6ns9DtjfLyRq8PNXJKuYwo4aZh
aJudQvIWQ3AnNgf11ofwMJDE72VsEv5R7mpcjDbQ/82DoNJrrVvHP3vOX9VH1qAg
b71nU2SmeDXWdd0FVqBTaNE36gdhLlnrnpTWZuQFURBu3uk3f3HdTqd3F8eQyF99
F+yHdWaJW6D6W8MpS0tQSbSBGMNUeuvJBx1+U1KUxdDVJtgswlT4FQpl9a8pIhpq
ehPyjxidMD6iMc9w4gjNgk7TrnJwNaONpx5qYXOSvp7mZgmVH9ltmGtTffzwtBue
5b5t4ujkfe77GfF7dwuqSq/eUrPiVN5xIZi2JA2pYyVu6MCeYv1DSG7PVIIO7tn3
5q/Bn5h5fE5mPB33dRP8Fls/y2Q2NhQExS6BMuUJxDbBhpv2josfnxwMCn92w1V7
46XbjEbFtsKxqHR12lWSSvRi6S8nrdlW+uxnKSORGE+pVmV1bY95qHlSjGOfYz9u
oM1ojqiXbyM5BWY04LwNd3iw23InK47wPDmOnMotQbfI55J4v9ATtMcFtw7wvDEH
Nk5q/9aqZMCqL3SiHK3o88LAk4XJv7GLET/4/QMNMcaeuczO2MVi7uxGPwEYTerW
pWvCzr+NjdeyI4pTNNholDkb4Vu5D7GvScCF69lRt4jqY6P93OmVI/1RyXHbrsAt
/IKOeJ4J49gDuR3wqgjmdFfOPjGEiQzT7+1aJdkwANLh4NUShM+V0kF+OzK+/kBo
q56CrQ1S4956C46EEIHZldDAh4dvI6oweRPsTFYKAslMJOxKUhuxaNN5zmHUSu6/
oc9+RFJ3msmcxKDcwzIp9DQgFzI2ZjulGtjMCF4eEawDvDukU4aBRUpYsoV8vQxb
8ddy9i7Wo0NlE4nvYyRT3x5q00ECxMeixgQ+XlxRsyPpkzrtQfe229b3hI5VuvCL
zF7uEO7XfMZMFTXfihlDYXWqa0p2O7W/mUbxPR/txHcV5MAC6YbkEhI7OFIb/HDy
tF3X8AUW0JVg2s2etlkFUPVdrLVumGdiez/rqZ36s7pFmNYzgUddTvmVPtLgYKHC
AhAwTvj0k4aDc6edqGnShVm0g6O+b3me/odb3pZ/7S732jeHhb+U/FiTcPfW9Gvc
tJjo8fbxnWsfu9k8W9vRjPSfzVWrEEI/i83ANtVoOVz3TikVxfuFjeDLWLQNih9t
qadbUTwn9gUed1+hh2arC3fNoCl9vJQBspCaN0zm7LOzeBxPn0NWeqZaJGIwJGCo
khhBrlVy4quoWby0Ya/Ei2GtSm3J65h+8FSoVBdqNXnMvqBCu/nLkkkLC6VHlbek
F93QDq1BPVTOjx3V5glmyqMb33D98m0AN98nXPgENhv6XBc89FT/QzI8OMjNt6NK
EDOkX1tw+zNBst4csn8yD0nQATFCJNPxMgIxaX+g0ynoBfgBbLd+rqi/QDMbQiCo
4NxJDHy1TO4WEHdRvTSGcwr5oXxqMKj7XT+XCrNm8CeaKQw3ya0xepRYzqPQM+rj
5ZqkBjrRDtKUqMW9NSYH8uKkpm3sNE3IXI6l5cV9t4UvOZuRmrx5gOpBbg9zFAVC
B/3mVD99Q5x1RPxNkXnmhE0JeAKB1ZYUYvySMSlmsqyitZtvDleRDaa+KG3E5xkv
ytblf2D7jmasS6pjUE/jLKGKNo//QXlYnwR5Zh63l4ZDjI6Xt9xbZBmGQEWXW/Ps
2rke/LyzxDj4I8ehyKRMIUJocgIRjwlEsBg5etxd6QNUByf8JjC2EdZYn7b45wJk
uuQ7PA7Sh3/BKkYRK9Ya88jOP50A6jUFpue+uO1HG7BdvPkt9O26zJzublMLwMoQ
dNHE8TImlh9VMTZXNvOjm3F8q0mqJJ/uvDed2+X9Bqnl4s6OrpfcLM8Vk7TOhwHF
9QFSOLDctr3otWsKwn8PnfmhzuehvG+/HD5zgNvqLABZM9QBo46H0ucGrgLs6Hgx
ifHmb002vbDB3102V+XZVpXqytdl2hckfE9a5hbrfTGXJ4aiswTW3OgvoOqRY0uF
pRwmC1DBH0cAWhEb1KXlQfQd3fPmhTDuHNY62SMp694TyFmQeBD5ZpVFSW43KU8+
8aby4Wye7ILjSpaA2Zz7wEOizpPAMKVyMgrVcL2j0vOmfCS9vYPLaCW9qdb/48yW
Jn6eh+XqffHFiJJF+9MH4qqmVmwTzNjyjbZXyb7EclAHyUSfvmGSstjbZjiTXyDk
XqYnrteoC8OmOpqsF3p9OoU+bw0K4ulVlWXmoCh4iEvFu2WtV/aGgk+49VbJGw2b
v8/HZr21RMWlXpi8s8AsXtt5NKgFSFUfqeFb1P+1g8pjZ2btaPjEFQHSQKbAYgCw
3Ommk2qIBw16727bhHdIK/PFMOhY5T7bp8nOa00XGeiTo0eE42AjUUKO5mpSLVvh
XItHBBNJgw4sdidzPi1SI/c2GADGKzzfCa3EmfD0ysmbFPvMex+/ie4hFaJY23ny
AOBW5PzxgY8TVGf8hQMl2qzFYcSWgRd2foZW6rgrhZiuxOqY8Y9d2pJfMf2QVgmq
nPoLA5zuvBh8ybBzMN1czizgtwVI4cw4S+lDF6OV+i04JNUiVvbl/RuvEFJvF2O+
2E2ZxT8SVA43AJnrsrnBPe0fjoGbiAdWz5yBuwXS/Sun3RbTQ8MoHDm7gWKFEue1
GREy93LeO8DLcPE7YTg8ER5j+m8O2w4/YQwKr7zCnrIgspDTEkFu7rt2kmksjl4d
x7sjaCmswvKovkzvqtHRNfBHbCLQPB1rjGu4jqxKuyxtk39j6+BK35HVDe5aQykC
qTHnhnzlxPfmPwBwVwW9yXnGnDqHkUykKqakJ1akts0maGeo/40ilnltVTvAJP8F
w/bp99jsfQEf8tscZpVc0Idr6O5NkBwFtjQp8rW/N0Krtwb9LxPYC3Op8R2OmEK3
RC37NjxT8YD68fkmdAcPjYjPrfjsN+RTkSClukg5XxcvAVz1gjqeBdonwFAL0S9i
rP1/kKEfFLVIXtGFchKCbcq8ODzmv2i3GdYXghT22lMycR7iMdKaBdQkLGBV4Kyx
YUs6yZ0NjazVkT/q8huOEGcrNqUflaNZzdfVZPCId0+ZJ60lc6IPLVNX/iS5NT+V
ur7BtGIXuIY4lcoNXwbRI4E8+F2XG+onhkoAwF8boCX2koVdJlz930DvVOhLmlVz
ve0UZkOxx/gLbaDIhgD8xEwza3b9ZUPH0jW04cgTVQYNPkEGh/SZGEaKVKOnSc0F
TAUw9yFKFtqaq5FmjcXXe+VEsEldHqnjzs3p0o2YmSDbwiH+gMRryVaOlIcjguwL
GyVetAGTM9gDj78NZsg3UJofnW9vzlzdFURaSvK5+cKs34YKQpMSMIpA8duM+xN/
x5iuIc7EdOVhmkVh+dAAPAL2csyTlP4rVh7rNmLKJ8n5dxAQpERX5+y95vmqZvpK
VpuMjouYNwevvO6AXeXoqCsIyBJq7XGztNLE6u29SNDXddL4Eybmbh9/72oRJuWF
rZONrgJyytBBwo6GUAHRGsgtoVjE7laQbPmZYjqlm54tut1tPUTNT89q6dzValN/
flAbLm5jXpqJwzZ8TSPgjb5ZsOm9eUACWzku8NWLQ+6G1M4oiwldPuyJGNp5m0u3
HmvK33T/VIIwPuroX0alsQtGdY1znn2iaXnn895WRkkBwUUguo5s6u+/Kcx6rAtl
p0ZWoxoQLC7TGI7so4l9d9/eWGQdY8SHxLmEebtEVGSYqk3Qp+izEgnI2SqOjWX8
jaLxWwrtI7iF/ypRicBTkXs8ZP5v6uxmXI2+tCCa3FK1cIAv1cUZh9aoZuYbnM3z
NEByd8MhUYHWnpcrYZe8WpwlWm/XvNa7iMOOiBgTrXaU7XpeY4Kq/I0Rmp5Atkli
0y1nzbLWS3ie1l4bqnYV10d0ckz9sEYEjmerRWtCzaR9R8Mw4/Z1TSOm9ZnPTkcO
E44L/QfO2DcNiAPW41FxllZsEDt5A12L20D06t54vOeTOiL3S9klfNZHmo+d9PVS
+0IpOFLtg9M+aJCYyV2EpkikyMW8k+WADPxxCUtqVst8V/VF1Igz8kOW8gEkxWWn
XzqYh+B8LseQLEzJ+t/GPCM1Fz4smTvKaBlzvMpAeyl0M79wHudYC/pzeD8GPOXZ
UeBt/Gda/xwPJfm2A9QnENbYiZRcAJap6JxmSX45fBtUMB+fRR1/zdkP3Y4RlxLD
1AvlBb5NA3IeJ8Slo5AzkspgeCc/Lrp6bDVxl2vk8PRTMvnK6b5Y+FJDVv9kLCRp
UzttX2LZ1iThgpC1tu01Ucn+gDSNYzvWeSIk3s+cW3w9hW+UwHBLr1onDRndpmLU
lTl+tnjSxGBdaNV6iWljGuRZATovbpTL9DT0wOaMzKK+HgxGrwsD8w2+Op8mtdIl
6sGYcRlrYXnVg4h81OL9aU7EJdKtnkUlmo7wMSywen2VDArbRn0kdbPiMdX+2KFF
npWMdlfJk3usx2DP8zVIOAZyxp83N5BW0B+DeKh4Krkyl3O77EE6J/Bd6CsRyQqh
288sC65UGhQzXk79mJGReyBl7XykkSgWtaQSaiD70MswWJryFD6V5rqT7L9v0ifz
laD0XHFKB7pWIJ046LOkHoLVeUS653Vk/Ksti/GqSEEdIFlbi3XbGPE+Nvvajex4
wi7nKOSEB2oBQ0gRH61VTJdZwDFZnaFyWab/2t5EWo4QzAD2gN+UOyxAvNo+mX0g
HX0llojxNOTBsXaRP2jgCq1/QqKGrjoYr3+vXk9z1inPg+7QnOg967Vhaj2v+0ta
m4/8/NAbJUD1EZVclS7hnt0bjcwlS+W3G+ZMHm5VmW9gkv6sAOF9gVHdsQXeVUBP
qnhJQAXvCkoSq6EUpfQrEthc6eGj+YeAgfGsFYmzkM2yxbLzEhuDksIJRNKPvT2A
nmvrxZo5qDbbvIURev5dm3eowyAtpYneGx1SkHu0smflm1cbHedRI9VBXtXqFMjJ
RTca0wyc7E0UvUIfgWQ9M1OmhvI+gg9x5b5Jl8VZ9yU0Kqzkd7SPSbSxhhO63bhk
CKl9L9RtgjkTNFHy+CoqFj9DFE339V60bYbqiJ9Z5RMreQH7kRZSvyMpM1HHMgrh
V+gTkuHaVQbHK5FxKn86ngAF4DCuEREHkEjzx0KD38R2+LIrUeN3xqpSwkttU74k
V77YGngIGOjkzDm6rSRxB1Xpd5qQymCKyIkiia3K6zCITWSxUKANkKj/iwEvTUVK
O+7OPizEfVDXjuqlgZbE3C7ByuW/sBWzEqP6LHI9Dxf13WnDR82OW9qNIjAiggFQ
vrpOscjKhzJIXFbJsshRd+mwfyNXGFum+KwCUF/1LNa3yXv/dauUoebMy1zV7CT3
etV7+pBonYV/l/usJqghBCXQtAQsXxXSBr2l8sVMkNMz4HxX/K+W5aws5CwvhJC+
RtnZR6SSyiffupWOSC25lgynpB5HiTP8VYD+LwZP/oIIE/7W/chMvD+KGfXpUsym
H0mJmgBlDv4egzSv8mhgnMS5mN0/HUp/WNmFke1+XED8W87kIUd0zIFrm2IP22ug
5b2LIyKCtIfYY7A6Ohx21lfmRQqjqRslBDGBiOc8akQnRE6AUejzBn/nvmUN1Kzh
8DPxKxJg1FCXFcuKxQpL0Ggaxr/ggMOXysM+tZ/XulCyEEpUxMdrtxxOb+Z76IJj
c7nKvwGBWIjX5s3EoNiCMohMIkCfCfxyTV3E3lpsVBAmjmM20ketIPndCrZbY7WS
6exSR0yfRpqzKM5stLE8ALjzEhABUKNwIN/O0h/3YI7VxWxuED3VqooeyPZrWQXb
l3mtwfumITJJk7s/e++oUkF6jb5iRhOJw6tRv+PA++g6zDoxh40yHyhpiJh8uvuD
182wMcCXCJiYdpGgANc3LiMJ2kHDzD013Mi34xbjhdahxDolpZy6ToseP0YVYXeV
7qUKhdbdosqaOtfREmZJu4WZaumVSsOjxsFFplz4W66unmGivxYxjCFTTO+PzYue
615TkTgnS3ZHGTVdcQ7My7UPxeTy56Sx4FPPQL2dtSeC0Rj5lZIaeH61tEJkB92k
q13D0dM7CMSZeOBcuynRQtWjrXZXEsc+RFzKwCL7MzigfVmjY2+/+J6VX6OgUuT4
xhzCG3Ls11Ga8/yMC5FfBSJVJI8MD7ZurMl7Hxky2HZoqW8s2+MZ6dzDlYBGUter
MlHjpcrtQ/RJhhm3siu893Rzo/LHXmI9kThgB7p42bo6O8J0swufXPBw1MDh9Uv6
eGPeyjeBaUHZ6eAcSwf0yKQbsnLcOMxGV1IUe7X8ODnCt76Ju+QBHrWKYDab5rYa
X67rn/iQCFQhIsjHtAm2qi64Xd+Ay88ewihlvxxG8KAL6w5x7ockPEiKBOfPW0iS
d3OAzrRXDKRI14+0KBvJPa65R5Q94WGm9s26ovRgelvaCBY1T/GDYbYSnSsyEeir
rGJ46+vJfxF6svHkL/cwdujheyN10l6ux6CQl3+MWIw1O9KmsbQ5TWj3PW0yAdyP
lOu0FrBkZ3iPnBZAAmxi4AP6C3KMGhZ29/sYe1Dh/XtaSPWhYH2alK9XHYuwgsb7
8vs4gjb1kuUHL+XwKr3Z7iX9B+Wco3v7Xrt/cvqqNPTXJECOHYZewU50zPZOEtYW
pW4c3BGblLpN3dGkUZ3ScDFkCzBKInR+6PY6zVp0cAQa8QbVVmAVMzOJQ/1J7QQB
ziAaeVBo9byedDqSMtIRf1ZG9eHVJhNqY1ocYPxBKt8Ac0AIj1s1/8KaNkG4q/Mu
qv0HAfCwqJyHFHqh/Q+COvXHGoedvJydK7HMQ5+E7pCdoOLN1zjMfH6FzmeMT3uX
rrkqzpnWE9fmFosA1zUGwPPjXE+A0MINeEOusH8/FFcA+0PjZT/066/RJCI1+L3p
QM2kw+833KOGEEK+H7wXWmdXfE6CnBqT5H1SW/zlXDYJAGEigS42TPZ1yMg/pEc7
k+HMb8u6W4c5NBeAJYHytMCyiCTio/A02PFIga2r2MuIJ/ZhNQ+Y0irozJi7f4zp
z/IZ0oRz+7TmkY31UJqG2bIyQd6qY4c67efsgLMg4+p0lxir+ETSSyr+5nHf9rsa
gK8/KycxK2vWcGr+8nf4Prb4u+hsLHhFKn3zzVziKwc5ZEFKWFSy4l1lfNZtb55n
X9v2IF267fH0B7lw2xMpOayrsIx7hsHd0P1UBvyJVOix1iEWs2s9bfOwga1kLj2j
Y+nhXi1xBR/+8PSBVCJPX+JGt50Xu+Qa+/ZOVq6xJSclVQjdqmW54v0cRiT2IAbF
dg3XdtlbUyhTbxAZz8l6eZJRFg5en7WzzQpzzylEz8BfYA9hu256lac2fADl9GUs
3K57H9qs1kSgLnp9vyBRzIG/Wyo+dkTTTAusW6T5vk3akoow49Kf1AdWmHfcurfJ
8SnsQcLsyr3MqFuN2wy7NS2ZTKgEPo9zi4jute2K1QDf3Jd/H+qUWgoPjsEesaWf
Ql8nx5k3winRGVXnGc6M9hO7dS3uozVjGhdCIddJ+FLf05R9mkrZW3P9HIYn8y1g
IhUvd1Q5GgoqWPXsbn+s4OXr2aP21qaWnbQ8eZl79W0XATNwpgV1Oi7DPPMhVX1w
IXby6UlK5NuPRwpigIvXC0rX23SQcAR+nz9S7zMIce6oD5avu1cdGrcVzH3Qasbn
SGnovwbw/c6zIaiZIIqpgva9u0oGTPnBaA3+WGsKeDJESAl8lGPcKKCVTbCk3u/a
pvf6fEKmCgD3HqRnXMW+Mu1msRB8oX7Y6coeGCj/qFF5iToNdGWmHaoehALwVOGj
UP5BnRGnhXftu0EzZK5p92480eEuHlIff4AdNaHdGmrp3P/BVc4zEfZd4yEJgvDR
EEq3QFyxDjr9Ap3gZ0dEGVz4jeWJQqWT/Xy72+sBa4tsXM8OuK8ESXAry5OVgg+v
8eDcPpuGRYCP6X2qKeCcHAEW74Rfa/Eu4JHP+UOp5DXiIZ0mg6TbLjwWQAlb/zEj
u2Wm+FEdwojZvv0mtZRFfa/tlJbNlw9/hrOi2c+sUkgLLlKH988QPDhjrTL1fZgi
Hg1YxPIM+d0HudeFKJvOG1F8y7/gu7DxjbIE/GRsQZfOmPhQQ1CT/xohz4kQvDQZ
85s39GiZHF1dvEayFjosKQJnt6KRV3ItYm1zGgZ6o1buYxW9LkK4kkj6qvAgxtSk
+M4LwZ+uQMv24ki5RGGemGgje5wVb7F0HemuhQOR07UGVc58k9WuvKnX8xFWOtyh
w21iFuRnqRFWPkMgr9WW3A5xdWxLp9ICtnEC7DBYdfB4NCstlPsDIcAt21gzqjHx
8IPVTFmc6m6KFxnvXPzATaymAW3/5lKpcNcMO/DmK2nXXUp4LQWPduTgTk51erzF
MlPDwmkwEvgUCoZCsl/ShGbHQFumyD/OVQBBzzcPqwy0BWrfQUXlSqxDG+AaVAhH
Xq3A9N6Un4KWX1bHoPtC6EvvtgI/jYXd2QGZwOg7gq/l4V/QtpMfTzJgvhsBV9gg
bzCPg/OSlhcA/pSnHdB4pC0dqQgKoI6cwi1WYCjIMY40V8YkZU39pNN/sUMMoyx6
EMjEuxNX5yLS8EMzNhBP3SAOmOEm68KVluy53GYC0krL8dc2FRgKuNwgYtdzcOdZ
GvZ8uIvNVXfszfqIcfmeAbaNkTNTHidxJ8M/UV62Vj67HSNXfD6ihSBSRF6LehWr
NmMaZUA2c6bs36b9hyGHeeBR8SF2f48wT9q4CaYn4wD56TINhCh2a3wcIuHXrTfj
SqxXklCx3j9hj3gdgDiJng2RtfSmpugp+/zaJepbmPMWBHndBBbtEkKZnV55yzYm
7PRictQ3vaB/K19m436vXX7OdT2/VgnZvoV2k1eN2s3pGnGC9YYOg8sgEvMsvnXY
4SMnU8IzLg16s1sMv+EFAy8FZ9P7eIlYV9fPRdzUV+6M+isFj3jqRfWQaRCDogYe
KD6hR5CQ+MNtDzVFxMMWciFMemRA23I4WQRLWikydZFdMMUIVDaYmC0QYZVOHnoL
3VgtNDR/SQ/tfr9+5phvPp/v0whXuCbo6GLhBoXRmvOQ6GYqgT8fJOkCPygjPNQc
JEDDGDjcPbZ5yf8uvT1E6wg9sWJkz7fKKbBK3nPgOerDkiXwfU+ymUDLvrItP4Z8
n198G7/ymHraD0IE5IUmmVei8qisLm3R5KGxhK+8d9lAanQ4j2xnDijnreQDqrLR
BLTBjlKNYr7eIVZxVvrgV5V4FO0wYtScH/6jtNZdfXOcBtQn4uH39sfG1oYlKezi
vRTWs/vIv2VCTG8VZmc/gR7BuCDafIH/AaWIywnR2lOrS/Wn9jfx7sQ18B/4ZZ0f
AjF2Lm0TlJM8+bWLK62p3Gz23uzwJepAc1eVOdO6vftDnwATObiHzNOztnIBG90J
fEYg/XniI9vJ0KvzlAV/1bTmZgkxTfdSEYroI/bFhEBb7p66irXyb85jqKjsruVe
KFK2omt6MPax0xeXVYJbYYS9kr7muI5rbg5JqG0nbn1360VZ9gzNWKCSf6w/6ahj
G/8u48iq1dZxfRTRi+uSK1kqfYuXxba03soE4+3VkVN4pwvg/L317e3EzKlKNPCu
LQYLQn3Di0O7FUYmu+msjwPhLMRlv5omsLZI0OFp9i6nubRNAvgTxuZamJUct12y
UiMtEp2LwTrbNFjZNqQit4XudBcjmTvddrhXGkimnqaWv/7z5YS5CTqZRKTICTUo
jBjUC/hWHF/2wB4aqwBsK7AE9HuA3D2XgSgTlUYxcUm/5wMEFEO98pFOTCn/CmIf
0o9FXUqhJbVuCjWqSn+rI6P8fdtkWQTu8W657Jn9OWY8TvwfpssYan8FUt98y27V
lZSxpJqa3g6CKjSId4cU+mPAJpWDgtk4RGVzyMxbCWMYb6d6DjliwFxkwL7yOBiw
CbmjoIy+l8Y5fBQwL8F9yEGFM3U09rrFYuw1DgTiwoH3Yq6jXobe9eTBW4OczcIm
nnEWLVZCs3GbtnTJzTZ6BmHYiip2brA5pmZY43SJ3uJP/1ThdHLCVgwdAie4kAA1
oOkMR6jEe+vTJM8v6SWHLhV4O6prtKXOrHRXwj7wyInl9EDaMJ8StpDd2TVXtwPK
zZlayW7/R4UaodLQabfZDR1lT2uEHPP67nIL7mAs3zA2yi6bkxcV8+ZZ/094GK4V
nL4FzH+fkcnLoPgG8fYMB5bmoDlMkU9VzUwfG/+fznz+SeOpI47cY3W7bh2d22ME
x6M/c59M91/yZr5DKlVRW5TjeDqa01NVRWjKXH9iGYEmHQKCpTZQGTEDrkHBD1cd
ukXEwkprVPfyxXkYzAXTNyyrM9JpfuwEwDSHFBTNC4kf7YZwQ4Hmxgq+svrRN4l5
sdOCp55HDHgAKcLkSu/TIFNvQ5P1aKSuK0iZU3bIQV0zcEeZDd9xNFk1b65vROID
gCQdzEwlEG9ciS5RVxeBOxLG6VjRChZSMd3X8EbAtKvqHCMyDXm5hP7rpnk6Aajq
qxJ5EWvgEN8o6v9sC/5qwBk9TUrDu/zjqRvzh608Xx6qiguOeWmRurwAZzSHn/GF
ZsZRWNhbT9NIzkO+jjla1XZ8As81Q9Pl5CHpUGGtusLwtFG0HTbVa5wkraQgDGbs
SOR4kUfzekIqbrwUh4GdTki5CdrxH6ePFqAGcIfP58pQhC/MF0LaPgcR1SajlBIY
YZqdNETQXUcHV82IMEuyalSemW/YsJdLHceYFtAyzjIS6W/OLYPs5707Dr0I7LEU
m8L/8jY2IFCblFUeSHLQxuBb6XklVL0pB1iANa233e2x+z1U8BgsTtgiyAm2EwN8
14pRiUCIsvHIxacYhqH68jwNQEbtEvfjaMvyND0AkDndPJsJfeM1MWcx77GA15Cx
Lg35K180DGf/OqSAEtWZDRgfoPFWWk70n+PT766ZCv/EWtS9LqbreDJEVAnkHjC1
yxkXPVFfQ495W9dIBQBxTbx4FzcT0RmOLq44rH18O7HHTexCAL3LuIFGAElNtHLV
qOxX4y7sO6HQ+sAHd3T10y3/aY6UUN/0o/8i4V1euY0uingxGVhia/Q0kMY37TDa
bHPZ1KjHnG7g9aMUfwUrdL8eVnJ9BH0dWDK91n3Nc07TMZkYVm1pGR0wdGS/h5tL
MMyY3F0CLU1aglVl4tm3f9YiZdWN0BXcFyQttBMqC47kKA9i/etv9SurSxWNguAq
bSDqt2FHgjPrW6x5tkUbUQxwEyoHuG1DqOpM8358tlb71M8b3q9gpCuMS6CZGgLa
CJwxWs0n8DYv41SbttwO9fmqsJQTlPKOqzOq3lN+zmHIw6OKKb/5NVSdMzCAC9XZ
Tnc5AZr+cGN2RzhsACIewdgiNqy+TM8+MyBbPI8CFWcFIgx0UHuXPZWOXHyBK0qK
aD8GwmdmjqB8YSomj+X/OtuPAkLaj4mEjw+G+QiGk2vtwllikowlY5YCArpdYljD
Ht9esXp1+9Xl9GJbnaflhduTcgXBo8JUuVrKyLJUMb3yCPv/aGHqNhW6vF60flEG
TOU2NfIdxBOFrfyxR7ljB3nu35JSVaolYNcKb0rqDwax+AQ3dgU+bDG8Fhb0Vhr3
6pr5f+cSNls4qZqa5IYI0hhkA66rxK74kKknDV5ReTGSxHGkEfobQIL03Gp5dTMN
4iXaD78eoHDCMqXQXRBW8BEmwql3YCrwfBbNIPiZ4dRSV78Mru5nmPQyvTsBp11u
DA3LD1rQGQoeKhTX2lDzos7/UO4C+yt2BPnTa/KuMzW6/qcI+IGcoUD8qT6rE+Kg
LaIDBHpURSUjD6lqqbxa94WpR41EzLvJHwd06+31JnGRragvF7exQ/f9twsLauV4
zjmgCJRyD88YyButV5v6v97NMYc9zVJkdeJWt7iO9UTlajdcyfFBes+VI/NQy5HD
8vqREgPIcRfh0H+v3UY+ZqY1+TCLcLrzTioNnTs+ID7DX0olX5bmIyN37f88gnBm
SYGtm7VVi+yrC2S3H7Zwwe9Gntf3wUB1/O27RkzQEMVURP39eK+FUUzd7Ni4MKmd
lwKcn1wO1rfAQrWQFADbGY6f+jVmqhBwQEP71Cu5ZjxEOkm4IquAEH1OXVtIHjgX
qk2UMFr6SDJs5Q26g54KqWcx4xVLa1xPzJNO0eSbw+ymM64Q/3xZrU25MFFYZxLQ
BXtnVnFD9j1Gd5TvB8w8MlPbd37sHsfVFibrrcKH9oTkW/mOjVBukSEj/eUvs7uy
Vu47vc8bFLUB897RAe2Mf/ggY9LUJq84MCvj3hZlheYLNM9PKq24EM72ODr5gMNf
0pSiJTdGbHHgZEvXx1DollyyUPccZTbzgWlAgqiK3USSjV6r639pdHGyh+sGoXFX
sdH9eAKl9ml7Vo9amB2Dohx+yQBcPojYXpvChRT8owCVqkolAFgtCqkVAdFhSRr/
nMV8xbJpLb4Rifcibi6NGgbthxi4+Cb803q0+naPr+kvxIGHsd3edMtlX6PfcDCV
EA51MWkXjw5EjFdGTYnjYo42W2UOe07Z9wcRxQui1btd1YG9nvs5ThzlXcTimm+S
fQ/+SVEmoseKzHnzHNck8Z8G5hAQisarGfcWAoAIMb/jv23nFfdpkYokA9M/ZeY1
vK/16sjScAY2UKZNKAkF5Twl4SIAZ3+GSFDQUzbHlSmD7SW/OkHldu4Yisxn/8Qk
kKJClju9os4iwOAEmm61kjWAcmlsJ3GFfcwhp32rOb/3BpvlQ+FTqEQtvy3wvr3w
HHtsNtmSGCAozxJHuzDDveHonrdGuFgY/aH8q1Lm5RAaiEJxp44J03kg9j0dYRc4
MantHOG5HJnWtaHfpmhdnb56YrmHSLBAP8FVMxBXQUzgPHvDbuQTdyFhRh331bhy
c2PtzMn6qlFe37MAthUOYCpUvLfCevEGCY+fyvc5ZWOPpfe+MgB+1SpuRmMkYmZF
3M0R6YvLAqNHSw15FeGyeCbgAjdZ0nt2REiqABCBVFisGeqHbkTL67efqwpYx1Ch
oOD0pojboTMxcTLbiZylx9xnF+2l6CdSJEwKd+zOm8lMurTBrcpk08tWltUxwIuQ
qujANMIMgSbZs+gzV23wv88Ir3aeX7FoQGDIaebEatUNWFpbfEMbufPfMzd9O+1P
vdDu6qVV+vr5aEdx3/DtZf7kCdeWJXYaz2eWl678cftaaSYMxL0wBgnQZtZXZiSY
KW7F6MKqdEd/E6NdRVhMCJtBR6aqyVC+MFK/eRj6OBQq8/zvuOUHKnNPDWtpi5It
Zlwlkn2ZsDuQ1I3ewerX1mipIMceRGtlOi0eAgeBIjDlmrkBG6BkayFzzASoXB56
Zek4fcku3EnZ71ltNrVxMJ/bDM5evreAtzJJ9wx/V8Z1MupeDcf/OqK+DeXtaK+M
n2fVxefmJIyuvJQn81k5q2351xXs03RoYCO5SBvxpgldMgCjpG96RaTx2yVrKAVQ
QXwBXBmTHV+i0UXOrQb0lPhzZSnsQRFv5BYHhVacFC4tvN53ZR3ydqdnG3DwUUvO
VwFWLKI3lph3XvCqi25iLCkiVkCSxwjBX/y2AUQn5IS+cxpDtNh7N2j/aCJ6bP3r
KOaLIwaaPP5ZwnFKSMd6zv4xpbXc7zqW6HbAVGEK0vTlq8XqfLK3/E9XeGZO5Tgx
5Ddnq7J2gMZWM5n7pVOTLjJwLndhJB0cuk8IYuDHth6bob0MD6IL+uvPizU857+1
2Gy9rwv3AMfTNXHW0MTlsUOPyCBGRiicgx292PD3pX56aNIhJxh8aVje9sGxDwVi
U+IyEyJSXHpSIYnjmbxlTNTGYJCqh4yzNoiLNP4jNEvNvlcQhGIJBv8I6NSX28ui
dHWITjjHzj6MQmfAc4x0HCFcYlYH88QErhXAPHn0kc6TqWXY2HSHWWt/JuqWVIlx
st3YnsHIwwo2cYvOsQ3wffWtR1cmpi/NmrGZs1bzuU1PPcon6dOs6B++NWqeW5Ou
XdBM4ZwIq+1tASvOMOzTV8hS6Zu/TTtcCS2kLE+ghhkSUCsZqQAEwZWr1Hy8LLk/
rPWRHklsKX5khY/lr4CwDgUdpVj0FYHViBKu2BMvg3GD9Zz/xvarQwMockSz1GN/
gU7v6w3DcmHqqnIdemVzL6ctNGao+/neAr4DzhgZCQ7U+G83/I5HgJIcxNw2OMQ4
0PS6PSOXWqZb8q7LPfqxi7NY1gx6rGZyHhNKKE5jnT4b6pXc5RdXRYi0H7E7+/nq
cK+PiwHCCphJLovuJbyHmUjvCQ1P/yReV2dC8QQNjgKpO1KKPUbYV0o18fqh904E
unSqQLxS6R+j6iiZ6TgCCH+mBMix5s5ycIXj5UpsuE8GPyvacJPhiUbD3clv4kaX
SXT8kKCEc1thFlqiseVVOkphcHMlkLl8LXIJv5+iJcfWFx95/oVgdz+vi7Lf+8ca
3ompDz3t09/h1Vjc5iPQQxJEV6u7/9njY0j8mOW4dYYB7qVdprBLG0Dsqnm1afRt
VWs9Tvb0KMb8qqozQ2U5WT2dLYzIHwrFZWwtT5jAkV6dxjfdFpj3dOjGjSnw/Mbl
/G7er+wn9L8YdNSNDvCLs3Tp0OZ3ZBBWdlNLmtd7VFOFuc6DPHxYi9P9uGEWCw5+
SVnwO1LHlgxPNvakoFWNIVuwA1XK7a/5L9aYM6quKP11KRM3nxtW1N7pXjCEEImS
4IpZwLT3wDIRxGhCjuksEKqCCj9QHkZ4khmWacxuioQ0pvn05H5fR2JAdV+J7eoe
zy/RByExhvNLELGJSSCE7f2gUdX6iYLTLJCVAO95n+34luY2rompVfFJl62LoxM1
vSWZNEW79YwBUTeOsnklpuR5b5W8hFb4YcmzCVC/UHoF7yfFbVJvCf+wzEua3mGR
PcGEtz3w7KtqvNTt1/7hcl8Yt0uG0ia7FTz+IEeo1OORJdKOPmNjcgKDNmEaCEbv
qGzfkOfSGW2P50alvWOxPTc8Ow0XsDhk3o0b7KER1/3kHgNjAK+IxoTrDlVhSy2k
BDHsOCs3ddyC54uqUzMX+hvn38WctxOt0KyLV7Ej19FR1SYgIVpLy4qjcRS//apG
hM0Kb0ZqN1CStunwNzRD1rqifD6qS7wXjeSb4Ks5hJz4ABkKbePLK6ZMugEvlr4B
L0S7yfqE7szm4z0UM/+a87tMgU1iG36k6fu3AJw6aRdbbeYAHlarJdmKglU1DRju
eirhmkr1BMY2igWUs7C7sBuNqMYVe4EaxF36HxshiGJoOTJFjT8xOANnCCPEMk5d
2qgtzQV29WpQ21d+HvZCqLFa9esokmJwauJ68lvuNOtEBLra2tR5JeDLOX/9WHKY
r0flnVtjPZdwmimfhoRR5ab1Uy7DKRUmbvLuDv9attTuXH0VaXMRTowaN77RqtCm
PrpWpzm0VxukdvQf8oXF6qiBs8j48TBseBQXGtn9ozYz6lTrAq9Y+grcxITo23u0
MZXlijvTAa4rV6104NCXbhP9V+mW0MLF+PdmWHuytPGv3uUTERWXseQfMOqTrCOR
h7sCpnTDu/hR8Z6SaD/QZ5XixxyEfxNE7kzeXKA1O9tOt1wqTHaynbR/3RCWgaj3
eWj8JZs8/QTb/hPKn1w9hUj4XXmzVII9Rky+gQBWZRsb5O7rYq5dJpStdC4OuElO
vRF4+gu8O+fSje41gxSyr7HiPuh36DHBVY7edm37NMNUQRVXWAf/SgQNOez+89EU
k0LzsqKTdR1qCeN6iCeG26A1s/PRHkz6FstbNRQoQZNRC6LFDiSUhJo8U1ujm7PZ
eQ//HYoz4qX/nM3tbEMj3k+ToLcxmWM6vALOW8ccU4mWoAg8tVseYItQffQyvz9C
0ozKmsl/0PjPx3ew/KPaFQfK5RzBaEU8oLk4QpW6jW3U3bm3ORI+BovWhiNOP5tj
sDJ5oyBPma0uOR7ZyivGgMZIRFduPHDHIrHjtzGIe1cXvvkF499pgj6k0hjaz6/c
pfIRRaOCOqMdrWNpV9fTVo3umcNzvIoPYveT3ohYAHqGsB4wyrEwSSeVILVW00sJ
bO1nLk2MDDNZIbjPeXM0dftXLlJc6FGs6ydcGTI4yDleo6bj6ByTmw0/o//K9N9V
K1BOvASmSx4RlzWzpgB6OuiD50SUr1ElEYAdxD4MRob75emX9W+J1JF6IBrA4y3b
ZonLYNP/NSOVc6h6ff+UQAMGpZ/6+osUv1OnTXnbaUj7lGfD6xIupdZ2HS48nEkG
MBMND4RLt4wMqy3l7FeJ1mTJ/w4nCeEhsSnaWp3EMJDsim6QzUSTfc9dKl2djWjv
9H3EGYxDfRQ+GVkxKoRxAdpHypixt1waaVhknjQsBvQY8XAlQAO4BtG1OByqU1mA
N58lkvWMWmoxbx6yM43JL1sCl+emehBvmBYpn7Y3MQAsSfvSmijjZ0nXIqLYZUWb
HP72asEbAB2wYtb7VNkRAEDOdBvMVKwfj8aQeGRU7LITQNlmx1EshY5EIqVLL6Nd
CC6VJAc3UkIpfd3JTSXfWM+SbA66ddPZTnd6D+kO2EZ+mmzxn+WPQwopzFCDox8c
a1vsAAtgH9Win5uW1c/9Bg6xUa8ea9/h7hK4Li61YbVv5I6KwgsBfz7qhngXhWnM
vgQ4ubhCsSOpnx+Q7+fzi+dXpj/MQMeEp5aE7xADU2lkrcXkR5Z+fylWMYrcvoiu
gl2UDAKtT4hC/D8yOcLw/8lAjV/14AFD2f34CBGmpjTiSDlH5JT9ip1yEykDRSWj
SDhDU6pzYDmBxbZCzeAaV7STJ4YTDvlOe/dk2rY5383BYZLzA2r5WuIvPZr6yYls
9aGagGsRhzeokKvLyjy6hPR3gUEOFDy4oqT9IbuhPLRTw8iib8HkUy3bA7zrbWRk
uXhX7i5HWlm+5nEkdIHaLPo2jTsfd7yH/6Ar19wKKS9OjGOyEQWmgvQ9B1GQQzAy
JeVEzwpRD1o8kb96570Hwqgo7siXgg4OVnC01AW7/3XdZZpe0vsAWWwzoH3LUZgr
y7DLcNNJNF4oOLNx3hVkaJEWYsAB/PbFtL2gd0bOfGjbJtGXa35hDyRH2eOqBN7j
6TWr8oMbp6pgHOG2IfFsUQysMPbtD1LTCYtDg6lzbfISWuFLZEgB1RKl4HtFZMrb
ZhSL1LY6YRExMoN5GHqoOC8bxaG82wqixQ56PM6jDVvt2qpyeijdsQG/xqim8C0D
ROi7KGNoCSb/lIpQYU35UyFvcpXdj2kaUYV9yOw2r3spqLLsNvz/lWm35j13Wp91
SUwIutiTkK5OqpHHdwZd1TorV/MEjm6xw0oWBfV4QCcTiDP4L0LtdAYQQjiJw+T0
KUlz9hhYL6FRFAbZeX2gqpmPq1+QVfUdTjkFGw3AtJbGWZHSmCToaYs447VqPGsf
tMqeG55ul6IyglKzLxhlx0bKd1lbPIA9FCX3alHuRZUpnzWijLp2jR9vxe3ApCZ+
tiIKAuV0DZS7XPO3s0pGn3iouT1K4zIAR0OAETfYG2ge0ngpyAek/eC999H1hwcW
PUevzvIaucQyI+HOBYjpccv/HnjEPyCuCyCLFhgZydpKTDR6XByUCbZRoEvxLqkW
H4bd6+tPBGTMcUXiqmP0w55ey5hzyESto0/TO4a213btOw4mySD4KTuRxU3s9BuE
xXlBqfU1NCXkM/FPYF07n6EITU7WYqAGUNabZO/PzBlfBfN/gYqazhr3BsIuXsNu
tXGGwWhkfZ7IhpHV1OcSqnRwdymnESkGgH4oySNI28b890eRkTKeQ6HzYV8MtzuY
yTnna0sEXN+ZKb4zUtHAqcos6UzXOOlK8LM2gyhob1I8yg0VoMC3fXABla0zqObn
Z/au6Vk09JbSSf2uDl3iiYKdgwJ6VU33vqUsyNVdDFf6QCxirE5VSZiYA1wH1Mqc
/ZVzah22TlWpbmUDdyMgFXhuKpJHOXUB4wlo1FNxTjx6kHI9S03h/Qd/fKfkZIEd
n2lc1KLt3zlQ35at3MjBkF4lE64zyUubyBuY6hGEYWJpLzJnA+Dt35I6ovOe1G7F
pNa9w/0pi1SJZVY7/n52zh6TN62peTfaMZyKAxQzVkefH3Xs+tegsg+LOTbGu7Es
1kkhIoofMg03zL6ygMFxeBZIwuqaIKa+vE26Wg7DS/4B44U81YJ6nKmjDwAMWd0E
tXpLWd/Vk9UfddUIUFEYOPnWXYOU1M1co8W1dDYEMCdmefmevsx/9B1DLA/ZexOj
4WUiGMOvVSWY7vKq+sRljkhH8z7ZPq8A1GThNea1jxern0g4X1tHb3goGqnd6s8G
Qxow4xpkwiREAfGsSWCleW4oGTO1iliyshnkOXTQjJShqyhFoXgi9qh8LgY656YV
SFFEGE7RrZDAxOETSG5fmFeocEUOIqQCXbHPrptedGZpCg3ekXDRGRnEFgn5c+SG
IW0h/4M9HcTqiqOqC0ORxWG94UUTPF5AJUAaft5pq7sbsAi7fRNuy5BKCtJa0WTb
aROn+9qZ2/QENUsqwaS3V+JY3UrPpXsqg0XSrzmP2scE/XmqlW+OBOBAi4gtNU9z
S4YnfM10YzWnTRdqpidOND8PkGZPiecNfhcU8TMnu9xkFhqp6PeQK0HBQnYti2DD
/JRRmrBzSdDybdAvVbr1AtDr9E9bN7GQxQqfU6zq+IkfU2PufkFGcNm7X2DHcT+o
UcrCOxWAgt01LVAl0/SP+TFbySJnMFtDW4szuiDKXxxIThmfmWAyLvFUWUrYkdXI
Vi7RpOsQ0IGjucEVTPE1AJ0II4Fsrg5mECTgjb1TSgxTH0JFPfbqoq68JjC54O3X
Vr306+T4CVw9sina1l1hc3Hadn8CQ+xx0nAuoBrZ8tBJO+EVdyoRgQdkpBxrOD9m
km5Eunh6whFGeim4AImfGAwgZ/zGdxPN1fZwrGymm3tynvbaXxKTFIVSbTA0qp0U
biKdQAErv4xNj52G10XDoktXxk4p/0lWFr4YTPF1tot799Do2c/Bi/6zhEZles+e
hp5VYUFx3BJlKI9PewRe0RDrNzRtTuJ/Zc99GZ1uSUlgYMB09vDna52xU03h4HHB
emtgrUmXKL76mg9TIYNUvKdW3b+a0QulHw8eXIciqCCINKnnATZpnfxbDvv//siC
Vy/IO5Y91oCgCIFx0K1GHwT9yEk8zR9Bjc/67ckvbTflmcJOgmRadhNVTLe5WkQW
0E3hKWBgdEACNmSdXkjFQXiG6/OJjGmERe/u3DqhFwKDsDwUkfyJzP3oxV6537Yv
3HoSrStBR/cEpjVHR6DbyyRxvpuPgDOpI3okyB/PHQpr4MisJiT2O8DdeBSqJH3b
tGFHARoIg/85HmYFtwNmsXkBbZUKQQiyz8+VQfQ8uOOO0YAF11fyUAQV9rRDD8VO
zwvgDGh97DQ4khBxz5o0cJBsMqmPLoNZMH9qciCBTow1b8o85Z+RDjJdmFydqJ3N
ILEHHESIFWedUXJCfkAbEYetxiLkmP8E6vnefLeqz0JoAmiKE5C8LNHHgyyxpj7e
SHAorcnhylQB6E6n8m7V5s+3BowbxqxitQa7ycCRrQcgJ9mIIcQIHXcf8EJNPBgq
iyOTEFmjvUTnW1zvTQ2whv5BnCeUkusr+uJZaf0SevPKyGUdI1By/W5rvfKg9xFg
JwBp5v1lJYb/qmLj7vB4LO/FCsuq3F2ygTgFDLQ2PG8kvq4eMSEkDg23Xxg9P1ws
/Xi3zG6QIH7Z3EV31c6iwD2uGbwVY7LQFOP5cUVhOQ7BT5Qsxq4uq8v0APZwtoSQ
jk5QDiTIvGIAUytdrh4WOw6c666Fh8AowByJK7cdt9n1zUocKUuPXMTcH5/SAgIc
IvXXfwDMBF35FH7F8T8QndrlOrQF7Qy4UrxYExSFEBu3zxznYh6lpZj934U8Gz4+
9rXHMnhJdNnBcC8YXM5C0nySEJsjHj1TGEk14WwXO3xmCrxKaQMyVheDDJq6kczF
J4HIkS8Jmll2WqLDaKdy6Ihu+fZ0kjehJeqs9kDgCNxXKDJcoJpWKwW09gFSxtrV
g5OjfEHKCqr0EQGSHr9PPGrFk7+2tSLbR/a1//Gaid5vFrR9lnLmjHxQyLlyb6D5
3nUuT78G8aSfdWGZSMhL9lOnRConYDZFl9cJdZ/8YSchIK+vh2/MFZk7PAzcVl7m
dxpW68rKGmYgqYhoGd8dJU75fgQdgnw4+/xvTqOpCFBWpQSWqiFj2ObGhumH/u22
1f8pikkfyiL8Lc3oFbKKV74CzyPvgPAj8e2Fo8gi3cZe3FRAZ0GflL1wGBGINM8Y
YYCHKnme1UDX+1ahVwsw/MSx9Lzpv8PjIAb51I8FXm5lC5ZraRY+VdAGlp5BDyfH
6p0/4WwQ5E4UzaSL7WTDAF8SfQ9PqMYf1Rlf5KZld44u+ClBAvlOi66urh/UGFSl
JOoNoHEv0aHeuqJfyaxfSW3DBh5NDqRUxh+bankWwYTUvlH+JQbp63q1JkWTV07c
GWQjkr0kuvS2mqR0hnCHcWE7h1sVhRtOdDB1Rle8J0h7OWqJKi6i693CSnnqRbSW
bdIU2WeLQRbZAFpgXRxGz925WgcETTQjbLT1rheedrZeLC+5H0em6K7Ucte3cXUa
3um5QDv9HSRW985d8oyTt71riWjVniiQtIn0SII0wD4mmS4og0G+fzkEc/wOFm2x
gmDqu8bu4sXtB0QHdfXB2HQk/YgV2RKY8uAb1ViARHkz/yMizdVCaXPbm3ztDFv7
SCJibaQXqSShpusNT/UHYNye3fdfPHWzKty9/8SgdU02UbjUFgmB4C/ApQOuJJ7g
YA0XovXFbCUeZvGQid1ymyVpoxAbwOfMgjxIn4w0nzViQqJNF48idD1ZwFPvoTmN
1A/dGPzFdQJzQss7vMKwH6qvBg/6eI3pDKSSzcKuLiXguZF0lK0j1D0ef/GwhToy
Flb1CE73B5Jy8IVjnQtRK2CKJ/vluaiIMUIbBIyS8U3uZ+VKmMMGkgeRPSznWztf
smVGk+FLfjUIP5EgwZBhiZ2zqbcyxQA3ZaICnmqJtnQsaf04zv+V5VM+kMiT+mqo
RsT0Hf4uegj/3ceeuFMREOVZdHHBLhW/fGkocHpg7qvDGpZ518HS389Ji6CaBqpA
B3UCv4Q/tyB7whm1lpOAy929fUEVP3bDjaTeJaDZvu1Kjb9CDIvjx+cbi9LGc2cH
mHaqROB4v+tuHySzPPYflS7hgscy5Jqe6t5CddM4Hn6mHe0qQcADXblNigzEsr2P
Rh5UolxrutYc6ME6l1iFWGOCRn2HXecoP6q63dpfcywCl/ma0C5fV0EsCHGHb03b
KF4lS7Jn4jkrRrZTOZwCNH0EbLeYWoJam4imXKn3ilRBbgvD8/DF0gmL05oFgKhk
7KMMoLSwH8PGSA+/0LVZ6yjfcESlOFgRtiFm0KHvG8cMTPRSsI2CjWwS0TzJ86cR
2i+0T758ixPLYcugxK4SRVCcKe7+Rn/H5r7PpQcaLv2HdbC7Co/XKQ+BC6Vm7G6d
1Z1p8+kn0G24apDor7M2ikgQtvStDW00Cd+CH5RfESz8Hoix8OmU5Ny/2Dnyzl0k
kh+FK7GAzedwPM0WsbpcVN8Dmpi6sL8rCm5jOBRyDnQqcyWIJhyIo3lyF9BO5Tgu
zrn7/y2LiF91PcVzqw0PKcNpQNNsA1X0Fyr1jHtgRdAn7QbI86GQ6oLNfSV9Ge2E
fN6B9yEH7qwJTBtg1fZvDiPRPlfXGxIJrm4mNN35DywwdecPKeEKh2gKGAyZpbER
hWjV/yFk/SvzXJcOvUTp+cr2+Oe/uy/ytsbJtAJLcrHzUxBy2/KfotXFGcm4jrDd
+zCqXlzdvwbCuCNM/xqspwOcR+CaofATLwy5PX+xeBmQD44zakC5nVQ9KfvYjB4m
26xh2RGN8tnSD2NkOXOC8b8hScUGqDcrImMHD6jzRtLoVEH+BuE+rfB4gR+8o/M3
u2Wtcmhq9JoONG0AXN/D1mVjtRL+TR1g71BNYzw3Ky6a+EV2cyM9jvY0vCHT45Gv
58PK8nksQHRX4Vzeur61ubq2AJbDS5JffEREumLOV1333xsTrocZuf5egU1vkv/R
jhdP0fPHZ8tBYTUqKUKuWoIMyFPjllAvWWQ4oqLii9ryuxsbT2l/qCI1vCVJXc3B
QgFmPDRa3WHCW37zIKQpyx7Htsjsb5xsqA0cHmAWhgPS6Y6qDK2VIsND31DeA7MD
5xbUSEvapIZ8ePm1IoTzYx8DDqJNejltgLWCeU1VGbpg0n441Y8CkFPkbSV3Mvjn
IJLffC+ZQgFA+sMCWgSncrOpeU8F3d0axUXO3Zlt1xG1OSLHhevkDa2q3pLJK6d5
+OIxvia811yHXzvoZ1jWWvVj6wibXGhkWxlZgcRAPeUdwgyVMshdUd3Ag+Bh9ERa
4mYlaxfJopIzzfuFVGvWMFeIWB02q6Sl0lfJ8tjpd1GoecfYZyYQiEQXATOG9hYc
wJew7wMx+0KBbV1H2/XLajRKnG6rbyw48zJyIP1/y5DnHdU5YABOaBs2AY7nid6C
nhZTpmpGX2w++T7eX9yOlXN2pl6sUgXL2SLWMc1rqBBkjRv0Ux6aEX93Kgmc/wuc
yxvOP7SLMcMkN8Rwd8DkxKzMCTusXaC6jp0HxAz+JpLPUI44Zvf57aweAv76TJxO
727aJXnKy51DOaNOAaBv+yOo+eca6Y8mSeApDCVqCR9VuiNsaF4SpRtu20K2W3cs
h1zLc7A3R3pQ3U56wmu5pyNwhrU8ljlymFn5ox7InFae1HqZA79nNdzihMxgpg2Z
EdCxs/upU1ikctsnjTuyZdjDGJJXoTLJFForjiEcfSYreOCAZK9kHXPNs1ESA90h
5QaSNzhGX+o5q6S5Up2ZGeq+XPV2HyGrWCm58gMvHC5dSHaTMxcazeCM1jsHVuvW
8phMHSa2plwO4F6W3G3cJe4aXfNoPhcNq4vBrTkczkaxSJfgYsw8xqe943ineGUJ
0wt589DmJ7nJDdJrNrfgws99vbbae6NiJ9NooKIIcQvcnNTsCza9fuwcIjz2x8BI
W2Q6cFSErymaN+zwq+Z3A2sdie93cYS48nZwZWo+74EWZB+5xPbtdq1W+/i44j5n
x9aPsEx7D7682jsxMVwynrZgRSJe5V32ekjeYO9LmnpOzlkMfLSmRAJo67vcrXOf
5Zzqq/P5j1Y/VWLDauTCKi4idKRSZ8DLqIFYPu8yS98D0pk3CAM56OvLm4Kv094d
RJU1yS8rBgBlywI7iRgHy59Pfjm9gEkBGdpu/Wsezw3ld6nQgUin/CmpdvT0yinS
7g7icwwqlnr0pcGjPrsWqfOat8ViXV6tzfSJUZW2BFuyC52yVMxVd0GLUx05EU2v
IZvGGndcZq/xI95STjxFeaNpnJ3Gub8c9tVXBzvOw0upN6TlYVbfDqvootEiKvGA
Z8ZUyHmGCnFJEcwWDqRtNYupYLvMpLJTKHSSla3B8Vjk/Gw54RZ5fbYPVjzkt+fB
QgzXmg5rmeZFxuUnSgznoIu2qKWrA0kWbbF3q5RSsk7luPG06r614+1z3Oi7bsHp
kXWFLHkc6GEunTMWMC4ALdKyQJnmGxuQ3k7HVHrNUOyoiNfJm1XywYIPLkcbHfOZ
h/Tw9+TB2R4ClmyNtVQjeiOnW+h1NQWiuPK3EfSYfZ8HeA/c5g2iEX56YkIfGcDN
IGZydSDQf0J/pg8jttdydeM+HyNwGO+JG6d4nj60v2PKP3nByDj//YcFWLhvQhap
dkqb9G6tUShwsCosCoxb5wpOGJSOMaPKW3pv+sLxIyuX/mhx5mJc8y4C0RBL3RfK
xKMR5ffTu9qIFdVKYlpEBPi1dgNsZKCNhs0OEXPxaCubAycSAj7GK01HfKPQ6okc
peHguVJNy0pm0RJGYN+jWOcywFOV3FxD5e3OYW4Zo//8T+Bh6AaueXJMU2/D8rEp
lpqiiLaMaBffBfblPirx8cWR+N4yTdC+kXvdiKpiTeHpxfsrtEXaUYX8XYVYR+aD
yRHeWUHV/qzwVr1PTD5nbCLeU3Kh92WEGg06hJKXOUS4F9sIDYKYlpNJPpf+4A/Y
ovvbhkEkGM5OXt/MugYbH8kIyDCUytA+RkO59IHRfoso9iAltF4F3uXlo+zO8Mui
UdufNuw84D9xRAwknLt7sMIowLYJroXcUgLrVEDWIetKSE7TVJi1dqPL9R9k+Vz6
rqiaLaxwtjuYhNd8G5qYgeZzOeJPUK/398g00tJixBDG7bEHbH7KXOEtJlTT2yOS
t6COU1sur2SubyhRfHhlOQoduME3ZdZTKsyp5GDU2BoyvAGZ5rLO4NTzPzg0SNTV
X1SlloSmr2jJCNQMiGaQfeTKQJ07WFmS2MqWwgndQReLC1kJt0+WjczzckqeUYhE
OS9AMwgdrKv/GNtuhRldnJObRd/qRzLsCK7Sr2KqKjlFQVjgLA9LVGssiW3PXuuK
9zwR7JSapkNMXRvkwhfAzRcj+roNlsRkIohsXc7Ib59nw5dFU9Y9VOQG7udWOwKf
qV8UV0GXmtmjMbT//D4wb07ujRTFOr1lwnrSxblyBLGd/A/SDGAG2epbRDMju77n
zujI6VyPrJOzIrfCCfTHwl8hghzioemm3Kl7uqpG76EsVyKjKB0FCblNIq9AB1EJ
dbEvg6Ev9cQBo+50480r/LQBQ2f/4d5wgdD1QwZnBQ0A8kh77lLW2bSyRmcuxP0i
g9nEuJ0GuvoWlwhdGQPP3C5gTZXMBIBqhSp7HLbTAbtUrQyu4q/gY/FAoaA+I6Qb
NdAGszYnfgYtRgzoinbFpwE6i6YKLL8sZegHp9Mg5Tza6oCtc57Bjo+axNTxeQdL
xM5cetLnmbQuXLQaBbwH5EmU+qX4GQlxrOwWMyG71fTTezrOHDAUG0AqLTScdK3y
M6d++WJP/sOPJus+zkgz7IrerVBYbwt+6F1icfbKSfe+5w5RBFkGIWA3OQrUfK1/
i31mzan3pl4mJVuvtFUR+ElSpDNOtw2YXD3R/jeyOvk3Yy+ZN9frDT/FrB6TsCPF
up4WUPhgzNte+XbQuiRum3Uw/fsdpFUKumCuPGrSa+jwf9/9Cx4H+tLF2FUx4PR3
2tBfWQzyTg1VU8Twsc31zKblm4vmWviavtRWGgKIkh0P4p8WbKsjGoCL3mPHKG/l
uPRnolYKJ6HFPnmhxuFO5rkP3eTx5bJDzRS7tjzlTGdh/kpZQPzH/R7PgQT3dxZZ
swgj/4Gu4Ua3SGAnRX+N7NAA+cgqEHd5M6Yeuk48UajO8ks/7+AB8KSZxG3jswMV
h4wf1i5Y+qaHoC9xqKH/2diCEY2/9RgwaCM82PbZr79nfx+IFrDYkvb5jR1Ns5mf
TNCDvG7wOvuF7K2kleEqPHAlOxy05C+ZUvDa4hD7P7o/RV6QHIK0SOJeKFe8RiEM
+mMsotk4+aPOK3Aesy9WpZrcnhvQg75GuG/q+GS4pOlZa4v9DLMd90TFpcefcBAT
AUhFmWLWXg7CfKPie8v+ZqLU1QHgXZOMBiAqMMhCjs/8qxTS3XadVlpUm6P5WEXO
bO51J6Vy/nZ5+1BnCZAIX6kv7Eyh2256ZxUFLXox1H9mGAxHFZMgi8tjok/yj+e/
38v5yFaNkjVsHYgkNEwFcHzJaJUH1Jr4cN8DDaQ6a30WALQHq4DMBBJRnoM9qaTU
vIbBa4u4Zu14qz1SLAOj5hLMD+NlfJKmPSccIKqDH3reiN2p07XjUBoXSU5sLEsg
zkRBJbqfhQHUU6qPesmsW2K2UT9iBiyCkciveCmmXAQWLnvZ3gjQHnr+di9NmS2m
6pC36aBjMjrp2Yi7RurfW8mRsiSsFsSoHHXZF1vPiJZ5WTn9H7Pvgke1bBK5LzAH
tCyhQYSKmpPzy2THg7iSOPqfYPfNox4TbGcDsRL8BYMFOev6hmvEOyuVQfG/6eur
zQfeKjsRdHyNBE+fahmPWX3DNTHA+7p7CeI2xdatii50DbfCgZcqctgDfSXYLkQC
R2b9L8Lnl/Ht7lnkfu4g9OiNCNbtbN/0DEdc0isfy6BKrGrzkP6QVDsfkuZqw7wl
u4t17n1f8+JSSBNTlv7iJ5FS3rBPxNumctfbjrgtG07F31BMmQMVMxAzmjr3ALgB
KudwzqBtKR3+W6ZUNFMjz/UNyGIwGnISYzIBkumMZZtS/s6HeaFJNyj6ZrttskHq
v00FcPaEgTDNV7U1JMCzeIu1PwGfZGO/jyDXtf57rG30hGo9qqzsuEon1Jm/CZ5N
tEir7j27BgBl+7T1fshcXi0AwPK07+vObRGUXto4iJqesphIh7DFWSJ3ozxLp76T
dSbXCuL3eG46IE8lL5qnwFQQrVrOEiwADlTptTcxtAWM5W/MeGwt9Y2Q3ZUFj4Y4
FpkENIGID8i7Z9bLYfwhzcg30n6LaY+Ljf9TIf0vudU1xXr6cd60wI1e+D5eoZn0
by7ijE0iVS4nQD60kUC9m1mdTaWixZXvU5nrCdbo+WXJ3IpbLXcbl6MdNg0vYQ6M
86s2MXKy7v0cRdI5GrH7hyZVvN+cMpBir+YE9M6Wu2noWG6y41438x8ebmsXNwkj
9970vezUmUF8yJ4fFYWMWfZX/99c5lym12OWd8TsL/ZuGzd91H7q/UCLNqFAQLBe
Q/YDS/XygReKj2qyCsH52nBvuZr2zUH6qZzh7Q8Gxik2toYzhsBducW3/zdZRolK
3xQjT0rAYAeFFO8MnEOXAf6uhOjtRWA7RdhT/0VkdyIa0+nvzkXGJMySFXxA8YWz
3dpys2l+qxNqnNvozRXWJUC+OZvY6GbSpDq6CaXcJBlWECPBprEDB/A9tbnbv32j
rAmimE7ZiOqYGRl6KwQYShkPK3TTHwDHxn5P3Yw0E2BEzYe7yWcFFwK1QDXQgFCa
GUzFPo6het3dmBVzkAohD/dCwLLS7Abio3tPWw/MF8ug1Fvs83G0WuYMzqyqnbcq
xrU31K+ss4AMS4R7oYLvcWzBTx0vKu7lSO3Bn+Rc5a6K+2B2140JaEU8hKCdqYtK
FBOy4ThFMIf4yZzaRbEZILHo7zP0KVFIcWw5FG4JNpl1ZtSbKAW49PEhg/yo4L7R
HkoM+feYXlEUZm4/bFseOBxcQ6wk53D3p8z3DYIBndKL2T2cKKJ7xWDFVQmf5Z4R
JtSobjdlj1KIk8RMsds2if35KBOiMGs2RFf5xqEI6mQywVvMiwh80JiaKIv8d5h2
De4Ro6QEpKm2mlGzHy2vfw1Vl4EU/z1T/wK8OBrvz2pxd+jvZ4x6I+GLDRgNHhW3
cK8s1Luq7vSgTmFc8Zhf6Scv0HShLuXj495nSPNtmH6nBUy/MkAPTdtvVJnyB/Cs
o55GdqH02OAA6T5EUZCjv/1s7rvugCT+jT+5x65YWZCdGN/xammmHjQ0wZZyJQZm
Qv9Dne67LzuERSVoT1AEklMx7751TxhDeWFIaE8n5b1e5w3/ZriV3AByC0lIrubg
Jh0F/fLCh2gKYBdDwhthzw1PZgKBMZyj2qfVGas15gI3PTawsOEVOaZoSaoD5hZ4
IkKbnt2cdxANSO4nNrvvixnDy3JSm8Xv2TGB4+lSpk3HWRQNR8hPPYIYc5QBXQus
FgO7oJsyoHIsYjvQLYMkG7S4/0NZ1TenzoC4H9BPgAfxAjvqgYK8HYA22TiirlN9
M/g3DwKoQx5PKmVJExOdy4Hz4nPl7UQqFXruPgMAU1+UEMHBA1jdyZsIR+x7F8A5
YRCVwtUsek8DWBLqSe6wp4GMmMNTznqgAdsveNnd6P69To5BSfJdAk7j/9shsbt/
SoUve/eHLC0kQdl+WiR8JCrATqfneB/Wyf81VgIuM+1uruzF6E31yV39PtCG32+D
NdSxJ9pfZ2qXTBIv1xT7Fgthn276uPrOm7LC2EdXGdYoV6sVczSxc5qhCRKLsINh
0bt1vVEGtaqNyjlPbG4aeCCE02zbVZcpaeN2gircHQW7Dotwzux+NOOddjsCJvbN
Hw9JPOvntH4fjo0M4HbjeNbr9GeVZjLsd1g2jilq4fkv9Tgdm1SdefvlHplkebn2
SWZn0vDkdAA17wLN+Twq5o4MFCFKa0omcVkbNX1lPkkOYwdfMXKncmBn3WVaIMSX
EZcmq2OtcQpiFUmtAjdAx1gyrxn6wA/cwg5VGYB6EZwJ38W0ku9nph69vR9rrHIc
yCiZut6jKZvEZjO6+ZjKrylMFBCWZP1A7Y6le5O53y5of7YJ/h6tvOfBcyS7139a
fxGNnPYdj1n8zEL+TRDvZieYdx0M5eFZPqQkpV/Xz8s3nAK0NpK9UJvw4vCkvL0r
nMJ0R+J06AHtIapptGvRnLL3+FX2V9Sucjhcr7dOOF4kRT1LzIJJZcPUfeEI//Yk
KeM9sj39Zpc3hqt370y6CPM8qmJsOx6Nz8SYA8a078nzWd+OlqUEv+KOpboGsJEH
T84kVb1z2KVmw8nqIRjsPQdY0nK4ufV/FnSvLit1uT/pjG2cQ+UtJkN0ZzI/pzeA
vDz+sduxDlsozOYqR+Jpb0PZ2T1XVOJwMmRilgFjhsuPmkP8tk9yZJtGqNG3rOJe
+B8e/UY0jIkrXPubdqOQRr/GiAe2k2qxwwANQtuema3/ISbe8w3cOpt/6DU/cUbo
wLvCOxQi0tBkFKNeO431jK3KBG8OjhH31tQUfwOjAaZXywnq1m0rF/CcUF78FIcC
j2aAqXHjI98f370cxquXirsLm7eHn0JsyANUOGoXCWo5926PJ3Tnp30bKvzrpdn7
Tc03w3GiKmFTf3OmulTg1kdO4KDhrE6iU5EGGBzCcZbMrlRQGCjHs763wliWOY5K
cfd1y0G+2D9Mds9CbvzizcQkiyVH59m6ravNqrEQhs6U3xUNHQsRJ7BXMablmjTC
DcGasvOi0B3nKGrrWQye6Di4I0s6eG7ZdHjzBshi6/H9+Q/8vDDefXlOvrX6ep3V
tD11ch9zyKIvOlgCvkTjnXDeqKqKftQMDN0Lh8kjpeI35ApOcMqJDXfP9uAW/k3Q
siQgIEVOXi2IDN2bVDKj56DitI+DSkA6ZoWUJxFohTKeM56COlcrVFiaCkFS345w
lyEYaurkFOAKJkhf3NW/+34QNN3YXL8iTkfbVClD1omD6hFFKp3osHGvRMmo9NQb
HEYKy+13hPiNtH4nGSpM6EGHDRL0jRqYA7OHvINWnO4F5w0Lpzaafybpi7QVeLNo
MaLm/oh46wTplWg4Krib/T0bJMFawjQ7iDYTKbBLfl4AqFNbM3h0WaXEEGgDpsKO
7b5mG2YaqBCD3z4LTWmvLNBNF3y0nneTsDypCDPMvyFqa/tKYziFCXcSpcMqh+/w
Krub3Atn7YJeH7T+ewg/UGgbHRvqeVU2/vj+UmQVCShSVkAZyMlKoBs0qRrZ1B5e
Fqg1k1UZN2r6dbMCGs5EYOVxAm3Q+UkSyAZgCzNJZvKYGd6tueV3RdElydalbivK
G5P8zeVmCChmAFZLBB8WfCXpX41RLqqTR9HX0jZHv9cRvQQ2BDVR4NFJdofT4D0g
0xQBlpl3asBBaZLjAW67h5jXaVyUVoKCc5cw7fqrbV+MeoGcuwcyA80oz/NnqrXm
WbVOShn3riMxirbDMSaOTIJ3dS0wuU/DNbd8gMrz6oFluE/+X+lqEAB0z/zmzvQM
TETkAmOz987i70fRA2cybzJhxmvAa36Q60T5cIDFTNTLS9VS0QG6ngQmDC3zg6MV
Nw6da8mnTzGdbUrOVm1pM9GI38/L/Gzn2G8ZDyLar04f36QSMvFJBObhYs3JttLl
Q4a7kklbbToZpxXiHmdjgNc6LRZqFhTv0VqsKoiVLqpW9E2NUK/nI36Ne28Vur0S
0+oWVl/k7FTAS3uKdy1k5uK/uTMxkxKkJUgkFFelV6e8ubQCTP+SA3BlzAqXUR0n
yvo8x3nOfkJb1U7ZtAnuyFEFRn3z42SmrMS305xVAfCUXBAeAtud50gvZo3UreOj
0clzLUM/d4zAKCJ1gmH3rmoiBLinSD4NoqpYoAZ3WGArT/TWk56EBw1uyTpurix5
Pui+pWQN1nKsGejku/KBYIj/0RT/WrLIkSkKlso21dAiOYDgTVIancwsvBSoLKOs
qLzaFNRuZfFWOMqO02DIE6e1vz8vZRUykdF2U0rJ0nghZ4QC3+nMp9A4PQxhXS7q
SaUuX+/lPIIoZQKdnrZq31JyDiYM1H+dYBBJPvPAm+AniOcfLNogln0QslnJ1/aG
qhF69IOc4xUqA/AtTlHpml280DkoMQGZpcsPeDH/MGySK/7ief9rYnXrlG8CU6Kh
XaOSZ3b/wLzlwyPtpUD//GtGJSRSaX5BnLO8oowQkCue2cA90HHfwfj7Ve1ivkZS
jfn1xQ/psmNd2mFZgef0ImEBVUdnqSkmCrkJ5obp0A8Mpj0Z3yfgmk+B87PQFtRA
xaj1jsqkBGG4Cnm155N5R+rN6kwvP041FbXL9mkUml0OLGvn3rzaX5R6iyZ0Cx8V
+JfOsKZ278IChdZyu53RJPqXJMvD1826sD4gJr5X8rfplP2u7iMNwNGWhhgAyfgK
pi+ipV0jVHCNw7ia+aEyhLMPvL20hh7N4Laz9HUZqmR1kDYg+2hASp/Vvm76QtVb
xpaplE/+hMIueRqh31bwmLFzunKHQ5xuJ8Qxs9vbyqfGTa5nhdGRn7e/PN8bwZQw
ZSOZVRd2NxGrs/intyR58L8UX6oNepPxuTaZBie7Xx/14OkYat+7F7Sq6pQ+D4u8
qLQ7tmYIPi6jBiYiiIq4pWvtR2MM4LpHVRDendZw0zsGC8GHffLib0IjRKwovcQ6
ivpPcP6CKylR6poYuIFGc7aIDcsc8Xgd2yhe6jeNqzlEX5iT6qO5jJclTn02rsra
+TysvA79szffwtwu0ZXgDBleeGXLiheLeKIMM9IU+Jw1d0fKkbELhjnsfnGN0gpj
bGoAJvtg70ujzoDqlTacBfcnVA2aPYq4soXAmXyN2JVD872ExKfmy7AgRoLu2gFS
SBjiPdqPbeY7U4MM9rHGVxbona7xlMN0a1zOyVSIbrr9itiENk2NQ84h8gQcNYxy
NHP5X/AqH0Vxm4u9OoEx3Sv1SncAwN7AlquHjuxU9JiUGVxgl9tpHtit/6S/3eFY
du5lV7PE99XkoxMRdLJhIm11VDFoqRnWHtvkTuLtR2VBjFQe8vHeRlY12+IZX9WE
HCx9wAK2toKdNWc0lR3eZZBYvhtLigI3MazoQvPCIpbcmxRTJ+3cCBj2bFgDjC68
zCwreXq01YUw1NVhUPAuDoIGre2o9paF1UIkPYNOwOhNN13U3mg7S4OulN6PY81n
8PMqgVF+oDSo/dp2+gx/zIujqqmMfkCCwHBBfUfXti0nLRnnzZo/IjlFomsfy3tx
8PsU3cn7SJIgJ8ema8emlVEWh98lzPObneK+Gx0jjusU8CjE/tBrIafYIEOYvBis
R9CyqeF39zYCgnUS9wQH8VfmkqcqUl8areSDuZV73HFaslPkKV3RYzcpVmqSeGrd
PgHXKA0Q4OCcuyGQ4FOEACA6kJHKHQmiN/GEcpIvO9KKUr3ahyMaiOPCT3ovc4Ud
PBqzoaVyqCfmcR4ulTGLz2PFtn4ZOQ7MM2SQCAvpJ07ruBvX6TsRz6UQqpCqn+Go
RpIJmxmby4xSQTyetONRm1/QnOxKx6yZKYvcG6alReDihzMmW7oPJfJx+J6e1/Ya
vzuhZxJFuGkqWr26FybhkxmOyJdOnbdLNbqXr4mWeB/Ns1oBms+bb4aaaz1vJ3P2
tNBg6HI5K+oFEo/2Oa0+ZIiLOhz+71er4DDmchxWpwtU+TGCeijtNuAWXLKx+yOf
NpaTvgoDEhUnME56xpvVKw0D61pC9mPRR+Eqd7QzQ+Ko1iSUe9RjtzR4wrdkcv3+
l+gZJnY0nOo9dV4CJanOCUYQTyjekpmei64ZuE2weMUdhfAwNKNEpKqc/xVihUO2
5RjNIuYho81DvIm3Mfa5zXjvR76JhuXHvnROTWraGJTLI3DeVhQbcJQ9glK3rJQR
pRx30F0ESU9CrV5L5ZhPiV8QMTZ48J5HylwEMjtaOZHB13nyNl0yehHBQfmmypcN
VDnhuFGkNwd99RJ119cXo3ta0pUMQTLW6bhHhTMD4bOZg9lXF7Yz7Nm0OdjqXwBS
/KPkeMZQeKLTJ3DqYNRiwgXTrejLD2KDZHyipUGOHgkCxqwpPb/eWlPXvdw5nXBV
Nak/E8/fuYPFKVW7IbvO2VbR6BcqL6fMb+oA26Qf19+ZH7njYUyGi+XWpq+IlqLg
v/g73qDPJvELbAf7utSU8TsP483QO/5zhLjoOr4FZ2eTgy28kF5jImY97dZgktSt
hklMdnWkiiBf9nxP7RZznxF7YvjPiu2TsZ6WrJEXo6Ea4u2XixvFtEUjLJTPlHeg
DkKuxLRBtaeJLQxs25lvnjxgSt8YWKsgebtx2lyirknEdQDiZixLA7FKsC/o/jIg
/MXEW6iFLSoF87V71b64g97p2tiapIT29b84ufN16/Gc53eUGY+sN1OuIboiY8NM
lLpdF86RbsFi9DO/L//z4ZyKmk/HrfW0DcttgJA/CfbUmAaXAv1d9lKpz1hZ/xRv
Fev6Q7PYSn0fqdx0nsVPgcDO2xtxz1CBfEP2XKS3Ts0xoBQk5WNp8YsIwrB5cam2
Y6E4rDx6pvW2HL9Y6lc1a1AA76txRQBAzmHvlf6bl0GxO8N/Y3rpuUSUiZXBGFOE
6T8j8GKPucyelbp39Q8m8fTKj53btCAXJKfmzBWX4IFPQOdCBj2UKulxYlhCmXhJ
APzV5sPdhb57q1TFkNqIfrOuNpkKIhrCJpjiuTu9+B5hOINHxIiwx+NL52eCEu06
lJGfc6fSnye5NeOv1/zJkrkmhk/ihYt8X+vzAYpJtd8WyGJig19IgiTdgk+UAs3Y
NMn0jlbcsJaOAgvwjiin7FHZCcaebX7wZaWd5NKuv0TlWBP9KC5zYyDuvLNQb73u
9mA4RpUhgJwUpnbC6GiOjkmCi+gDWg3C1vKfGUdFCT9OnoFgN7xqZLQd4xjDIRnX
2w6niiFlIghB/4FkJMTP1BnMyLSlekHtGgJ1jwssOz2fdkBfeHD49vvsgDaiaCgd
Yn59JhFW4yPd51adYKZ/Gjw2OhSgOY7udACk7oCiexjxC41YiiC71HoNoS+AaWOs
NavNZ65+h5ilnKgG9JqHO7NI0XBLJ4E84wn32c6nMoqV9rwU3arZ2fQYk52r0h55
hBgpOofZKQwnmGJqFTOJIy0uDZlFV45iHYQRgQlchZbONvKuz7CZSKgFnp7VoeJo
lHoZ6LhhsC3wlCGUhVKZ+ZUYDsZUaPXx/d0VA8DuUFfwEq1EiIJ5bEhm1+PZHTJI
9AylZ2oE9n2LALSlOTssFPadhlBSTP607eUANPFXKw3tVQFUnIMJ9IfWrIfzX79Y
njbOZ2TD7oP0sItOGr3rbYF32WoUnVOB7/m3ElyaHHVi48VXlSb1PwevKlaiJKKC
t5sRCPa0krXI27CtkKP9L2ARZYrzSYXLyBnc3auNXCaZZEatNiJN11LCs/O7E+Kc
W9z9e6FiX+L4CkxmAoSKXaaHpDsafuDc1ajb/flmwuFstvRW4vUs0zE7LWB/ZvUt
ENn0jWUHQTW7s7OpmAvyW4HKyAs1spd/NAr3OGFw+F18yMg+1gjyCew1ihLu1vPN
BpooqZgvSEeqkNzVY2J9k+tmgAney+duLyNpGT/tXN7C+s0wTPF6Wwj9k2bd0lpr
9Y/vHcyudGt3lwdj2M6XC0D4KFOqVSb8COAaHRDSxA5NPhHO8xjiUpbC+V1OfyMT
cMvkzTZX4gO1Fc2JckFtSVhFcYoPLJ7O4xHiYwHKyx2xFSn18sSWNe9sQzOd4XRC
AfdA9fLEIdy9/ATAEj5/D8Sv8ecEAjIx5N+sB9J1SDYUW3PlZbnHLPQaFI54xBLx
6eQBwIdFzkzDKS4bijnszJYKAjjvudA50HodBE77sA0DxmWB3Go7m7mwEmN7KI/M
AR2uX3auWWXBOzm4h/j9wBlVhR8LKiIKxl9eqqhQ72BQolpvTNcYRdfkhO5QYF64
p1/yUNuYdPc/yKlgfp6WOxPgrQgK2HCqUl1pF+TIyFutkn+FRPWvjZVebE/hLBlH
9VW3DX1NbNfFc8ZS7JO5QCsIqyNlEX28w66u67tliZlTEgsI6uT4RUnnxPckHpip
/axVq2E407VO0aXDz/bvRVGLx61aMZGJv93u/2EHrPWGswmOOW8hDlzNZtF7Ods4
fIiMIhh4KqMcrlHVey8Tq7CRRmohbziRTF56hw+19jsVDo86Nj1tDSJOtSLQNNXZ
roUW9KbzyoPu0+HMD0Ch3itoqARI32Tszg1xT3OtC2fhMRBT5s8dbU1N9iytVXBD
4qJg5LWDaXs6PLB5Eh4mh4vphNRiUjU0zJZMRXO+eVm75c7rtNHAev5bFrE0x3YC
lluCKAWByfKMtG9lBV3dIvq5x3jAt9AW62eYGNvNeom/y56kjWJRBKcIuwZGtVFv
1CvuTVA9DI8MbwHYChJM0tVAj+ra96oVc4v5f/eVbmT77YlBYcmhms5VKtB73sMW
29igcwjxivUo8yHg2/DR9vmlRh0CpHpOP6d+35jjFG7QphPtK+42wBbV/62Rjhid
rZJdgyvF5e/+snhdTgZ53BiVTkPSyfK3qbzpT6cBrcB2LqGAEdaHD3a70sHOVXo3
YJM93xcICl5Huv6xPPzJ302dh1IgjweM29NRcG7zYXAPZKrnIfyu77DCJEhKznxW
qDOmA1uAQTR0zGAxNORyJBA5JMeiOcW7Rqy5qzI69/3zlJMAlvGw/gsOlZs3CI3t
dbkSBQ2KWz2uEOAhbTx1y/FVOapH3zEIvsNJXrzCMZ+HcyHPZSz4ytG6JwEAvHMN
OmAmYJlwhXZrqgd5QqZM0QqNRwb0g35SbnEAXgXJAlYW+y0Zk5ldHacauTpUEc0T
Uk5EcrMBULM++LMyldHIx0MaMaOYOdFw1yTKGG+mjB35kgyRibnQwvdurmitexVv
rzPZQ+7WaE6jo5sn+HCiYzppJqrFZVQhAjxlp3z8WeuGIl/4vMr4WznbwD111XLj
7JttS/CmV95AN+au6TeS0EYsf59MRPPUZSLytIMuwISDUfBhj9r0PjwmyjOGjhhX
IHOo/70i/5dKYC4pezNF7zx6G2G6zi704fKbQdqNAebSE4WtS5XFgv0UlQ718cvi
DtajlH5Is4pQ8b5ieaIh2PqehzGoC96+yRR05J2xikSEDanaM461WalmJ1prPYku
lOneOyC3usRGZA+aO/M+kHear4RQYmBOOkqUAjI1e7hazm9Vor6vAZpQxkRRbgr3
UL5uVO5DcQUq6yadv12OUhxMfVO6ZjD0ai4NXrURXk4MShv/QApNXKzFV++TUsS0
F9Dmy0fCYBQaypLWi8oYyyBtd4w6h2OnyZrv9S4HvHb4QIlzkqmqcofRrXq55dtG
PCLaJnR+Ek22+WvyB9f+Z53/WaGQq63lNJUIQuqXH+nMbmOtoDYxHST1ZAJuHtPH
hQth52X6GugbQBbWSiUYG7wHvrybB3p79f4j8zoKD7llA7dLRvTfu4nncY+7ABzQ
Smyy7fDjanJA4jVHgnP8F8ZN1vxeci4O+iWbX3YkhKnTdLOjp9AVbFHFORJ8qGmc
z1wnzeaVzFlPO74tI1d07aZySYTWVrOg4NZt1E98sbE+mqkh7p9u6J3dg0dASbYe
0ksLoGwje97Ft+0NPck6lZgcCG9oQ2tDMnsMRpDp3XavAjeykAuHV933R/0WfV6f
bh0a+ZzYgkWd8HmpzXiEIV4DoUCyqtwsoaAOTLYwjbemos6VFOfKX8XBuMlEG4oJ
iuXGd0uD1Ep3YEVrQzXdQ15gAWXDNYy3G+3AVWFIEASIBDELUUiu2gT2FHSk+08v
0DaHWIv4ljsQ+L5BGGwKkKr4XZAUSA38mT0+hnSoJn9bpMuPyMO8EPHybahnUFBC
pZBdYm0jPQ32QI6gF5lu8fB+QGr3Sns/OUcglXFScA5Nh0VTmY7lmVHYshK3JY7q
ZCNnlrIuYhVxkft5DrI+5MxSQnRkwgbqmbLomyxI0D0Ny1Gzs/EmUasy9Vo7YYkf
7tAoEusD3gMrqObbiSHKaO+D5HajLaH9nUjsJ6T+6p8g0/Mj7QxJVhmH8fttgaWd
ymnm0X+o3ygZ5AiuEvul+7hSN9kYMOL2rH/2+7JujUF4/Sn99osZc503Zym3bi53
26mUnY5qqEXG9G3lq6C35E9wbP3gM3xl6ZvBS6hmfzkunMsF6m7RZ0/1iwpLxG2W
zm8Sn+xyrkKcKnyqbdSNpHklBPZMvGs8awJDQ72SbNCFQX5KAxPJfzEnLG6Kj4Td
NM7+sDLxZZ7MW6Rwq8CdFDNRIKNHISzZkUugIs7kD++N+Q9aWasWObkG52wJCA9E
qbZ5sDbFCzcxH6PYqAHH3vgNd/39FrK6X15PGIK2RJPnyqrOaW5b1w3o7/o5nSea
5VRWLkUR3He68hHAsx3qOBhgWD3tfmoLZJlMUFVGSWDxQCsTouYtIOZkP8mgfiqm
MXhhy5PhTHwhp+qWh0ypeGPNtv73+bSAD1AxYkHA8MdCtseJNYog9Y387WhzC/up
Pj3RLg731fKvOsAnZIGiru3PWylHWNIT9igJ31IwZei+K+IKDpYhTxhcrh0suwDy
jw87XWZhPOtH/OhwI9rkABNefdcLK+fL+clbIcqs1lDUalq9tZ4FQL7IlEslh/0k
Pz3VS78fnrdFetUFtBUcLQkX0xbBs1D3QKaV3fiME8tGwub9bEv3B5jbTxwVIymp
Kwfc4+Kmi8SghCt8wXEuxKoP9Wg5WN8d/d09zVPFQwuuh6lJv84BRISmeKXP6i+B
zSUjYoaRFTGo5unJURHL2ONXXHjVmK7/p18aIEOD8bDliR+K/JOr2y+tgeSH7PHV
Vj3Clh7ADeAp1O9clghEcLRJ1S/siXFDh7Zf8peknhu0IAyf6RtLNHirgCp8O/en
lnPOB0JE74F5MIGi8YUO7cTsX+JvDF/4k+qEmp8Uheny9AMjlapQ8cMKaMVdJYdH
aV4miE4jXnwLIn5lObUG3jUCxOgysjitB4O5YisnjGlDm5DgqYUyh7S8VEt2m1Au
hxBJv1HoaVvu/INk40vHlW6AvHCSz4UOk/cYLkmuL/fH8ImQHRlrwAe2eDMNKGrI
UYgjkJp2jJbW14GuZrevpCruJjy6RHy3yrY+LLP/LfJHUI4L7Ps28AI8i11MPoJ8
UvrQBf/Rs9G2LC7QRyqnBytgsZRPcuc4+DHUoGuUCjb54HfB98Gu7QeQq6SO8h0Z
UY7ojmNDgZKQyePsBox5Ff78RcEgeWyvQE1Bw8b5oK1Xg9T9zFadfjNggTLGTBxy
iFwtwHgHcXkk96kL+Aty5w2a/TSmmZ0c2szh4/KoyZV0giEtlxtLqiVZnYj4K37c
I0iMLgpovD0G7m9/gUvPSUusZMQjueu9KrC8LhIA3gMik0wN5izcN4bhSIeJqlON
qwTqLXAICBtZV1N2+dARUABC9jDkMmuz+EIw07hDK3uSxwbNMgt4ZTuyET2RnLJN
jAfZj0Tti51EcBE+9YVbyHMXrBsyPSgQQnS5hoybqBspcscLv3F74wwtL2/uycDi
CYSXD9zoja0nw7BiWLqu9yOFeiskcWnErD9J7/riISqQFhnmtYOcXCa8FSw0i4fB
tsCaRr8tvpNzj6h0viQUW343E4sm6Xq0eN5GlBkAaFPruZLQHVmdT6/GcsGYsnEJ
4w204z3l+8whw1ym5DAL8ac9FWOSEZjWtMagRN9jrRZzbxub5Dk5/QiuD0Zk+BPk
kL7/z2tFYO56uulGle5AeZrALE4WILuAYeuXvuLx3y3yiJ/Xnz5MWhVXEPBM7cEy
vjbXqqFt43qmB3H7QxAiL+igE8rJcAy9no4oKPogcaaHwOhgF0ucSDSzpxDSu1Cp
s//s5zRt+81C0YY5cCiUYLX4SXITdkLLwfSB0iaarhS1Zh2/Oz9prZD/0ghH+JM6
IxLz3o55gbpbDlltCT8u1/pOhfBpZY1iONi5hkYrub/YDZ0zjzccoBOZXhqEKKW+
h3puoKrsxcnUiY8u9no+r91JO9PsYpM1EPzIv/Qe5FEnRw2tkgP1mvUPuNc+JUiv
PU6LLYJvA/rMasjfEd1WpG2RzVIBq9O4A+St/Z3WpT4Fhi2RT4JvCsXSRE7SUyoz
OBo965973jH1g6AUZfx9FEp7bqz1q9t9F4cM2ziVXEERKaATVXNOytyKTyNhvgbu
wAwCC5PcRWrXxHrPdNMfkFtkn2yQUdPfO6EuzLMIKK+YcECR70bWKWuFJeNTacpW
SM4xZUL5jNNiF8RoBTDE/WAvHVY604BmX/t1kA8J+KIdcp1r1gcYhRAlPwsPrYJa
VRbgYoSCUhANdIFBdy07HdDsBcWh0yWBXEl8DhsqAXvO3gWdSWJdUi/iEDh8i+Kd
5KTnkN8vYHM6SmwZ57mPkl3akMj41vnNK6urBVmj99i2FjB/3m8CJFUqLXqM3q2C
kZoCfAB0uDi8aNDAkCaiztbkHA+VFcShWSV2jY7UL7v4rdlr9Nn0mtt6u8Z3Uuqf
eb/g7Pv6f/7sQoF486/kJuk7E6SlSoWJZaxD+HpHThxLv4j1tAt3/PODLyaMnG3/
wZvynb+vlakegczKLUkyflSI8Wx/DmW/tILVInXp6laOroVxN9A0ja4VxsYu+6tn
bKSJJ8ZzXzLLFC9ZdMmOmIqUbQjQR9nyY2pOFMcYZVeqK58Zecc3w6hTcSUxbOtu
IPbKRMaPQ3o0qiyU5SEGwSEE7acrczcLz74JLirvcHW61dncenxk8dtadM+YVkuS
+Bis4forfqmO5Rgxv9LRkBsxnQXx0Diq+dvWHhs3txALUqRnGx5XJeA85UNSGost
Y5TwYUdxKnBdThxHvmU89nUX9qoYOlmXDm+qrjHzVUmQ3DTNvJHHKFMfU/OB7W1M
mPHrFSn//agXJRpfxqbKXIVX8u3Rn7idfH1/51K3KI2ErjdmN+z1T4KWqfsOu7VE
Jmrgrh7dbcW9ZXUiQo82sSXaghIr5cFSWLyK/VoQFINd4SEkz1NfJBYYPBYPbuda
JjXaS26qsk0H6ogAczpMZRIrL11R8D/58UYBmBvzpniDbhHTBfZb7xMCUL5o4f07
XiHf3pCJBXrlg6HxW/mr+4TxIAXl19Ju/27QGBt1lg5bvlpMKZ3Ta2g0aF4ilgIH
YH1BnoG+Kupex+khp8ffIY9IduYVcR1YGkdrOebcpxd2US+X2VS0aIGWG/wbBSF1
P2EpBygNolh6BpORWUQPDAvbrs9lBzJP1uvHs3mpIacLLB3ku/0lhGUrph87laqj
CBwZEEh8IKOkJCJtQje0S5fSdSEo/fHPxnLTE3HT/B17YXw1XpxJbU5gwxn90XfR
h1NAH2jl/GPLwjNgWbirO9/9iJw1zIC8f+18pnZbXVOmvYqyP5AYkpsKguqYOyUm
Jnw5bsluqtUVT1agTMSCDpEqPonRn10gYoRnN72F0tHALT93ClljjvXRz+zwA+nj
0aMhs4yJlHuVEZlIA/qn1LqwIabRgxeChBhb3UJWT0/x3V9wVAwMOYdRHTwboLdl
2i5+r7smgxl7tbFWGcb3npHxpXlrn0U/m08Gj8dS973YxwiIXVk5gWoFED/PzClf
IITWqeb9yCyZPJifK+Ux2m8aPKEhOEZ/IRH1yyeZl/+z0xszNI83yDHSltxoz9O1
cDQ08937BQ3uP232n/p6TjJA/1G7F8zTC9pMv48U0BtuV4G/N61hH8G20L+Ubl+m
mUlIbj1EmFCdmozL1mcOse8QVD35CLYf18tthtLtZQqMnO+u3zAZ1x0nQ/YbQX+t
TNLL8K/+sAG5ICcBMDC1YV5A1F/El8Kxcn0EjiBZqRDFSPhz30dxFlr4YqfZorpU
8IMxEpVtgrgnJUsFQOoL3rPuyp2NpphzjkMvGU5do0i0Yfy18t6rsxa+QfQdMgZC
wvRaBQ2GvB1bvw67j+wmFtCOxF1cQ2heG/+JNkMhHoYEI1vEtzV/FQUGIK5zjHvO
GeNMcUhavwtcM9Xn5lp4iXhCmOKnC/Kp9+KxafIT68Su05iINOsTN+1fg0wVcgns
h8NoS98pQvQn4WqlvunQE/w+OBUUx1vQlFsd28YLyRYhtpRPcFdBzf6dv1vWITD3
zashh/UJDJgORPqiPSbjZRfAzJ8Q8AhjcVVMHQDB8icNENxERIYJph/BToYd/y1x
P9ykJb0z3H5kRTmaf0MBRxk8c4GMe6MK+pH7Va/Lmd1FCSGTwKJRhRmiLYGdv6ZM
vSU+Khr74lxSEA5FfepX1ep1XMRdCBxaeq1qHzHyeBO2Rqjrt0EPKmbZBQVGn62Z
ci0UMP+cyn3HsdO6tSINokF5zm3/BEgJ34tVoFeUg2VYBU8XnJUZPCGEdAUsbwbA
5M+l6jKzyOkBWpegQpcMfGOg8d+QQLArEiFyFVaeUido/AXV6vHpWKTnmlXDQd1/
nFdXletRKXo0jpcQldLIp9fIvhgR/UXH9Nr8Jn1E3ye7Hw3O9J5+HIF89OjK4wX6
a/V3XDcbX6cPQ46oiIZL6bKO/5mLI+v2l++rbN2ZRDLcUlswb3W2kiJfCs2aEeo6
XT55dJHfwzby2lxFeLVHBEClZrkWFO4rPp70YfOXIavgJfx0gga48+Mla61Njdw8
AX0OIcm2Z4ZKuiaM5slReh8wBKWVBaB5p/Ynuow60g6mFyewu+NeHHB55nNMBriw
8CoonR5MkfKO5nD4ZiY1fX4K0EbIYmxEkqQgGuYs+L8GMPtaRw+0WPwe29kO6+R6
+9PhT4NYq8DaUOWJNoGs01m9PuylRnz2r24uIaxdqaUFrfMUSd4RaNtRHYRv3uwy
bndzvxfgLAYWTifcs025oV9x6rsyfcrG20VcgWROX9RSFfpn1LpqVrsT77aJ2zU+
4Vd225uq2R9p1DZ+DE2SJSyEBmfw0kbnDgvMX/LBk/QCmxdAkzrBYpL/fUja43I5
6+R8ddNRwxagxsvy58dyPTTZuUWVzfe+xrNpPu8sPaRw89ZQNc3fCgpNVXETf12l
jpCkwfaiD71of8xcAnloN9KOfxvezgeGMkaFc5YcN/R7J8Tf0lIYAPNOJSz4BEEj
yvFPK/rEmIwc5A+OZF14jJOu+oeI/OlYx6b74ZUDUur7lvAsXoGLK9BW1Lp4Fdcj
bLccngWnmeGDO33Brv6ECgfKXS5OGtP1EA6NEQvmjcNM3w8IZk65jBSkAWoU39HH
em0b1by6366S7on48hV0O1u+Y1V4KWgqmHwq0EMup+gSTeWJU+QZPEhxJTtwF9zh
QYXS/gzzPBUCnkY02Kk/txwKxQB7Y5UgQkfZq2LkeX1xoP1dIByfl4wyvEgXeb0N
2/AdzgMUH9jz8ixhusIMircruL3GAneud7oa5FPSzcK00mUKiVNwDS0ofwvWa5sW
/Gx1FH2+zavAjHZPbncNfGAyLFw5CQiU1WYiSLNJDJW7PZc5HjKivwsANJJPuO1x
Ni3c3J359Y9hO5vqA4vHU3VHnkgHIThHov6uwEvHZi6oPVMXJzZm+B+NPJhzx55C
L35QulmQ90npsGY8wMfz7pVB57Zp+gPAjOH4skAl/w6v/vteyGasWzTYK65EZAvE
9vQMLUQb0oS3tITlxzfd3A2ZOEV1Blfg/CTkQAPKPu2+EqeRmw3+Y5ci0qCSmWxJ
KiqsxYY9up58Fub1sWIYRDIlxu/9PgHBbT56XviH04y7/mtkSazxkXXDLgR6qiJl
H37YOZwxdjr4g26zWD0X8POBEgwsZ9gN7qBIwNv2vh/4Atk7OPj9km1wKzmBurSm
I1jzcQIlBuAAMTWf4m1on9mwhLwCh+CN+9X6kDz6T+weQwnJkxeroeCpMowIayCf
Xd8jEam7tDDBsiNHDPaXzl7TOg2kyFBzCBsP+Q6BbvjLuX3lQIyp0ihIMFFJn/mm
+RGPxaXQUcAJyHCg//zxIHMLxtEsOoQsX0vnEyFi1UNZRlCHkGvyoNTotPvH84g6
2/zoLNT5aII/sKfMyjvwXoubKWYjRAc4WrnLgIMhsRrU0QtIk4mA2EuCDWYqzLXb
Y9uyBvKzHfPnNOitXouqRIDIQ962zR6YEwyFZ2IoSuVeiGuVdVEsFemO6jt+5EcG
H5rBdctuSUwINd8DiIKMz+i6j5BSdCY2Vw59Gxj+1i4wsckqPfX2leNKxUlgJieL
3H0cdiq5hOBkFbgN04a2uT23SLOIkJohT3YNo2wrywc6gfjvFurIRXA10hkVnsmA
GdKIatmpu6pUnbO2tJJZP4/KCcnbNv74+6x3OUs7n3DxfUCQ+vPpovBUxrKl6+CB
jNkEqWJa1pjm9gDZ11145kgt77bxTOV9gy1uQaJNxqlgScCZym/j+AtzrGy9QM/K
yz7wuXjM2GKCnTedquiCLomMVohD7G/piIsEH4DVhqgIbn8a5S5W2/STdSqavJ1i
KDlWii0erbUvtOCd25sT6d7I3RRHLe8gzYmLEG/qvIV+dvjj33sEuPzY3/MKccko
OEkso5Vh/GeOhZYw000FJtdMNXcnqvUDGdwZvdsrq/8Mm53KYmt07v76YIRRPSYS
xQc2VBcU5BQuT3BITOoSMRvxLzMWesUMnwTaCKVIT7PLU5Zb0XoV27WM6KGQBMW0
sq92o3vo298nB/dOMhgCbqb1PyZVLnr2uo5gr5Kc4CeaCY6YYZRsaZWFm8BhrUsm
s8CutGXUSrOj/XdeHBEdXy7m9EJ5iAT4NCAIWbwz3yBRgT9AY1x6ivdqjBNb/1Wl
e0s0ljWLjHf30ikXsroDn70DT6SPMcJ2Ihw7JOJ/yOLT0f4cJK/4AjEqrp7VP3bt
UwiIavvuEhn7af2AXve7H3V6iB7AvbpNo1K49Xz1Grg48xkkD6rgxZUqLAojsxNP
hb8H+Jor0qHSC8h1HODnySsxgmwz0Epcbec/EiLfrHKWANKiEHgB+sCkGRBcqWqL
8Jm+nEKSpo+oGWTWcH/ppoFw+LoKgSGb0rMCAn8MAj8ec4td4ytJJzX6swdKCQxl
OPTB55qY/xCVR7nSlSGV4AR1O7ReTxZQa4urgKCLLnzdu1WeEEPOVxu2xRgG1fz6
e3fBTbmbfpS5+cSj/rttfcr0CTmrjGLmON4Qb3RBM9l4SmH4+hsE/GGY8iNz+HGx
VsvsRG+y5Wom60/FnoMVZImQ6asuDfw18cTnmwt9Ei+q280sHG6MrrEEQ3/ek8Bt
KgB3Dt9rSn62I3FoBeLMBO3NoMeGbwaUhxj8XiM9fr6Gs7h51H9hAGL7TWMhJQ5k
SbNRmELJiDgf+l6eoQfy2VkIG2ynp9OwL8dXDZ0AYNv/82guDw1RNry2Hev3Ue4H
F3nGUgE3OtMYpnV4nMWCYRH+gv5bY/yBAVhCZUgyfmlubfog0ko+nLrVNg1ZArj1
KsU0+ohYY5v1wMBdEqZQ35R4Yr/cgQvcANBaX8wXyBlqf/bpERADyeJ77cB1koOP
hpdzAGj1L/bwt6kqyjlOtxcb89k2xXdeSsCJC18q0f7KXl+hEm8Z6ql6ggQ7eEeu
ppoUzkfflSElxt6KqIK84yvSF7t2wiUIUJAFVQ7pbb4DXzU6WHUUoRYAafrpgsq6
59E4YvI6hCtRiWJNQRQrlfkq/qPrZHelJVKhdoJ6EqKRg5tNooqeR0Sl67acRzpY
3WtplQ0XhJJbzNqXgB0wI8/AUd/XBMJaJl2ADutUKwj6aRY2eJmrFBbeV2JnIzaN
mlnEIPWKR97zkH+Ko3cwp/BN/cH0YDcy0lhUdPbK0rSaNpGTTDXZYHSYbTm+1sdr
yVBB7lcLTwbNVMkZ+tdIjYKKffLUs41wKMTzrMgsXfOM1n9DgihyoTwRz4f/qcjq
kjucmD83Afq8q65vQrdBPFYYETy80fN2fOokym+PEuZ1eBpx872C/Oq5qUQBH1gr
8t2MaWBR05rRrmdhW5c+5DSrwjQ18e4WHuzQWY2uvR2Z9kPnX3ShOInseZCS0NnP
kb7UwOD9U6Tq7ZR8PH8rLZQ312h9I96ziIurvLhzcLmqgzMCOHyCT8nRgbKRbELC
RNnXgX5xB/BNYwGG/hdC7KWikRQuo3FDhCTV+PERCNUOc/Ukmd84mnA6FCKXsY02
gDSyMMWi00fhc76u30TiXbe8GX2LFG/RXL9FfSFwSfhwFqLWxOyDa4guPd+Nh4l+
BO5o/WoK2OJ8QAYm2ZDFBq67ZmMVQPKowwPQzA/myPidw1a9OU5U4rv4miuUQbRD
AdoPFyq3gslCfAEtK6sihckY9w56D2UmcQAUUp252LmefrwWna7udEGEg/W9IKto
FbREDmmva4r0EQAfrVa6EmgviGwWfoybP3f/OAeSCTeZcHUXI/65wgl3GAsAbRMH
cCUjUfKE3DsOxVRR9+5Xta38tbpwqWWWvNKoqCXdjEC/yRCdx8q221pchFR4HiBs
WdvDUeDM8HquFt7u6MVSh1MqtaBj2ek/1EwDbgfnIsprVeGt9tdtsaeUohP8eF+f
vwMFZxoOHABbCnXsavvis+RiiYb3LkJ3SqdAgo2FhFmfNGo0U5KDUE3rshwMpu/Y
2GaynQzPkYt8Rxa34HlEswnLnddDbcNTpV6xdJ2zoJGZXHaTbJA7v8tCG+SxEDHz
YXTNhwcoGu2NGD6GdrECkAVtTxGWT+3oxTDFoNdgpeVV9H7QSaXZmDmM3BL2ZZJT
XA9IyO6acZU0nDRI6qe4po1lijqjF4JWWTwRsPiaG7dAMBFUvWDV6k/BGT1K1ySo
zsuf7IO7RFTlmsznSztiXMjfuiEGuQvu3GxLfapPYWMH8K66Qc3evvUkmtWTOPjZ
WBYvknoc+/pwUlAuRvZ1Bxn6i2jcxcWXRdXD3iujj9pkGYhCDIFbQZlXAtuEynTs
7AC6rZW0+h11I1GEJMMYCBnZ7GXFao+2pOuhRMwJsTwdG0OFN3uRIXTWqoNMEwFS
rV7X5K+UOBu+YTauqeiiyRMRwj+ALPRo/5xV0KWfR+vNe0uRFEwWQJlWnInMJ6AF
3dh3Y8qqUu8iXhzMRv6O1u/Gos2AqvBs4sQ+WZHakT1LdXnyGPAz+v0AZpYxt3XS
+iRtLPeA4/eILOrDpCMgLiBxw6a9i2xW4VhxJLdEpeu7zYnblNAfGF6OiE9DIvqj
dwU+8UzMLToK7rhjDtbzNG0e0tnFEwCERZewiLMmpnA2mc53pm5XkHHUmTvNZoU8
YvFNCHcwSNDFMwsXe4K/etXBOUS6y0GcCtQUvIyRkRPg5CC5ZWd6j/FlJwG3pR/C
ljVPVthqNbHciyA9fDorB4CiHRfXQxa8xmCPhuc3E/F44S0kOMsTVhYT3nNURRnD
rEqoZ7g2buPD/Oz8wEK50ixE/nEVDyIs9IVqP+4pS5rX+oViS6DIg9rO0aZcnA+r
J83x6RIYy8/mltS6NxRqOpucMG3RzChgRTUUGCYLNqKXnlkfzzVPApuOp40C0BvS
9k+yXkbL0VOZ32VIo5srU/00PTYrhOIuSmL41b+pbGtLk56UrHH/4NPbR2PQ2lx8
KjfJ8eTK6DQEcExV6VstNgDdbD4jJ36eugOInfXXbZKN+ZnS6BJeY+jtoXwUcj+r
TtMDWamSRKYaJWyrHxWAOPavlhUsDZ362GmLl/K55zecRlyVGeJQOebVnuKoJRaY
AKecFjo86BSaBxy3IBFsVfmJX06SIps2sU6Aij0uHMagUYOQn7KMFv6v/jXuhTG3
2C35q2H9ueOkl7R5Jzd5uawcMmLrqNO3XbAk41VY4UZy6IOY/53f5EEb/Yjsfg/J
6B2gQ2BUEjhTsSLvzUGIhwvHFPz3jWudtP8wY0Ect0PZypinlb/7BybaTV0jKmyR
xGQ6R9dmIJeBx0CqMQocwLeEJOZ7gD0srOCr1TmzMPheiuEzIs/p00SU8OgTCpQX
/U7bYKhDfwh621b5p9So1B8mwmLz1qVLdqgOVV8u4WEO0mLIXBeUR+PHON3i0Ylp
NiQxiZMPghsvQpQVz0VtXesD6cNh2S5mSQzcOm4m4+YPfFaa6zcf9h2EGTjlWIvE
L1uxJgIq8eSRGTKx6sQMwODIvMIYfjiBAq+c4DfWrIozr7HFs8D7lZ+Wl+Q0kEjP
NMJrzdJ9Nw1EKNv/NhBR1IcLkIM6gT7SJn3PmJCXlPBx8Lqvk+9/bi1QofrQ4Pu6
1DMwd/QwtcIZ3yD0I/P27mKzfporPdyHv4Dfo4bF5w0uip2L/KvCGnfiLgpo4w60
59xhFsx9J7eagOXYNAvadRFTNcRC9b43EFoC94WYk51Y8XU0axCf4en5J7E2Fd1O
bFwVOPnVkXVpi5z/qjlyXtR8G3Ec8vYhRZOqalzM0nfFexulrXOc5Lr30S9cHsb3
h/a7DwofVNxzk9l9UU2HXMAa8V8gf9u8cFc8L4qU/khYDv4R3NWiTosE5didoDoK
0OiIbRKmCl0EsS4QCzwSw2TIizmNkE7OEAlku/uIntnXH9tK07IcBcUw5g0+cSBO
kbONb9wCDNKjCOs9i6oKlEjFuvTJDi0N2lz+FTkagRhFkT2V671jzHC85Fi/36em
QHxxVSEGB+w4/yEsVFkKTewwy6ubavOV5K4hwWhVJyIPDMpBsAFf9t4LF1JTaVqU
0reDraHQGadDgeHrj52iKhDgcSB1zhq70il8WdjHVEDCCXawBu9AkH4tI0JSgVkY
oU/TOKm7xs9BiB9lHZ0pwQ1Clhsjf87hP62rt5MbZsqNiJrx/w1w4ZORviOMzvIq
9iNUszz7JBLZC7Wk97iJyL96BZJJaHA8wbQxn5DLJE1uONR2VZq+fUUlC25Smtez
y8QalZbXSMO1gfZTvxHyHqUBaVpJXZr8MRzXe0J5/wbHisa+1Fc/4Mj0w+hFQEgf
q5vEJpb34tBfYS0BrsgPt0N1DSEcGYjC1gF1Mk4hByF2PWZghIld2mdY1t53rIfP
n8oEGJt7pc04UHptPsGMpDOMnwPq1SKp5JQfGD4Tc/nsPq97Js3bGE+sR76neFL8
Vn75uqHSPuq6/nERB59Z3whNYQq8gg7y/CIE5OT4+yp1s2tidn2OlFSpSfOEDEpD
wWgtsXpyRwVqN1BgGMg1IDj496zMysddtYV3lZsqfinA/HrXMRmlvVMLBE0hc9QT
+wZBCzjKDM5c/2fMWst9nTsMMOKmKHlgIx4w4oL9cfkgeMi1l3XgT4vfTaDyIUCH
M8Pdc9/+i5bbcd5fBjiE49fmmiyDjxUZBnfkOLlQretiz5eNvCe4ofCfLlbDT/Rb
Bmlq92dSjrpdWbBtMk10ssKSHzP0jqWl8xkNVe9c0wix92p7sdOYhkJwwWC/8a4b
atBpmNReZxbMp+dT6LKptkHuqiiERltD9mcN9CeC47AZCSeSP2J/vPYav+H3GjY5
2G6iIzOV5mFJWnjtVyVWCzDAZMg1eXSIQXuoXerXVKQOgIO+6mPwhmjuTeW7VSL2
CFaJs3ck0M61uIqaf+wg5yqqjiY9qlQ3P8RgPnwrA/BQWrj3R/078mfYZMjCngCm
2SwgAxTPnaH+KV1Ikv/yPpDdBjl+qKthBfuddxC748iyv1Ru+e3tNEpPhfXWwpDU
tsFvxsoqe2I5sr64ya5FPgqCpSDzv6gPRbIUVeVUC0yNFOJ9mIJDbdcIW5HrNBWh
fxycl3TCdJUeDhErkhTe8FObuMrr5z30W++Y4ikrebd+7bCHFbtTQfUSbcNnUDd8
CUnZM6kdzOu1wmHGHhGWliECIx74Q3AlZENv/i5K/+uLisSv+/5GL0oX7y558DV0
j5DnyUJT+45hsYaS0CB1Vz+2E4GzL7m5aRrn642VDYXjfvFTk3rQRVuAX9Y5cX7e
qnFJZ4YKhZH6hHeytRcdnJKS3yiCGeTW3z+yO/hLFS+IGZK8eisdzAYRufC3s/EH
Jb8qrcpIogiIntPITEfzZ51r+V6HbiRYZu+zKclV6gySsi4/p9kDAOJvKJFSNm2m
NkMKwklc8n8nwmB3VgdfZimrzrXytqqt2aCdTTcTEkr7U7vA9kNc2cCzIA3fO34R
1R1ei2pzfBpZ4I31Sa2kHYETS6A50RlIf7q0KQ7x5VoqbWgsyPAL69DyxUE+fhxb
8Q2NVVRR0hDH3TcJb058qTRhWlPZR8pf3h3IcqevSUDCRlAEj82KR3PE4IFqt2Cy
4UB4eSz/X4noTEoua5OC9qOlZY46Nj5SOySeDMDGVnIZKtL0ADLsMe6xt0ADp3Rh
7fXzqLnLun8bjEzEooHZRvcbXAsxydOx8Mq++J4+2vUSaoBj68J1H2ZJ51uolTpk
sn2zzc4C5Ml9nbDVjPAbeCzBHTEoKK6d099ehHHwUbabqh6O/HZ22b30h51ROT5Z
ow64SBzJXddP9/xXYXHr/8Vu9X/0fu8Zitr3/Pe0hfY8XW6QEVvC2YYpBXZSLq73
OXGpJ6c9qdcQ8zMDtmjr3nBMD+HEnJVfvKQ2PqeHhZ1gpTppw6A+eEEcFXOTbspF
rdjS7VdxQLfHOHVDKQ2eMXk0IKzQrkGAxILOH/hylS0mnFvklo9QGZXjbU6LEkUd
82Nyzn+jmcPLbFw/xo+gSGfOc0AZPdHxoref6IMWiRC1C0hPe6Ng93wEY6icRIiW
cv11UjdSsFR4BlVevV0AryetE1/mcCxjc5ahw4KG33+83dN84HyWZEZMZY9v/Xi8
sgY1WOCWmaQbJ4efX4z5tdat3bn6rS5p4Ddy+KsUYOdCb8QgyFOUmgG3YHX6neKJ
SM51xCehA+SBulZpd3CJfhVFBgl4BHhZ7zibpjSr5XIS4+Vk2CZawjqLu27D6B/P
rV8o9JxBwyqYXBhZm0tJK9qBrFghnrGIMAn0RTOUwtHwEwMHQYMPfpcCmXJ8rMOR
7xn+771sazZsXi6xNpLvr9piA7jmB1LCCd/jUnEquyBRnjtfIMq7em/h5BOGSt1+
1oIbtj9KOjvOYr5w4wTGss887GKABgjUT614D8siOZWMUmtXpBiW5Xe2wtkKWe1n
6quvfKuzAP8Uzp0iakqR9A9gsxbnNEe5QXnsI4NjfAcmiWWMcPqYMLnVgGTreJD5
UxzKHeoHN6hX5jy2K2VoL7rtbE++1yNsPxHeiWu1ZdBVtRCOiPw4+NIDAxDdqelV
5jgePv4lBYU7V7jwB2eIowCDxzQGX1C6rO7q+6WI+K20E/ltBMSk/9SAeWwc6ajA
AC6HrGPKnuKLZWxmOClmrj4KRIq/3am5eDYEfc7Z3169aJTSohOOsg6N0+utrgH1
Lzvi5+vviksqVbu7gJbTzOFHfBLvtmp7Zggs9gU7eN/4mnu+2HCPPW0ff988XXG2
ZOVprVhbvUC4DDayzjEZ/DRCoOw+hrUE/mOoa6JtWzi81mXDUO8Zpbf8w4JdG26X
tsYLVJRsMrUXRhfkFZomTY13SH+sunHwze6vuyxb/hLCAkHb+4+W5ukq3L2PtP6k
YyEPaUvTUKnG/ZstQP0njXfO+tpBQtkv1t0XwCv9/uRTO96GkcFypgap5h+Cr0sd
cvU8TbW8868S33Y3I8dKTMWoBe9i4+eOGCpx2lRrI9UdyH9SnGBmipxMce9UggII
MaOBX5IrGBISzFg4TZYWSGWIuY9od4lhdbW3O6zPYQHblF9vcIpWbrvjylYr9fcN
uBNvT+RdzJKujYGhlSEpcJIEp8Ua8j7esES0J9qlOPO6wQHH+GsxiDoM1wxdVZlW
3btitYZywGhAGw9Ueu3Tq2i/alDqqID4UPN1GIcRyTcHWowmvBjPvJ9PbKGGCg0b
GZl3QFD02cmOgW2Iv0PqPwg2tg/7r0Uvz44QG/mzDUXT6lCFZDP2zOxHxj0b5Pyw
TgeCnqds9PknSh35um24iQ7knxVYdLLbCvmWlJzbl0Je662RdCP86OY64tX5pTyu
rZA5zZEeb0QDTDoad1iFZiDh7Dir6LHdpU3+Pb4EIFDmOVher2u9Jk7HS3UhSK0A
9vDfqY2QxEKWcNr/oPm2VhxReCHEUSQat6e4iVm+n34zEtbNgIME57vN8y5RFEd4
nsvSuSc30Leghr6LglHLBaWsOUZPfmvdXx2s8FJ6hr1cGstjgaeK3F5E2YPIxVzs
4x+ctgnuoe+D4s84MVCpYIRdfA9j+HxzGEIGNxAk4a0BKh0iCJt0/0FfAeixyXmI
tWef2ZDIMt91uAD5vtwGUN0XleFKyAmrQaobyO3Jpa1NXBwh3RGLd6iIIaoU8LKw
twVDB87mb+wz29wQlezMQH2cnzaqBk3+9nNfVlkEPZAisoduUOYOWtgL5wHRDtwj
5UdV+o/RqFjb1wKkNWVdhewq2ct4jdYtVX8BamO9iGv5AYMzbmHeothjfCfRBIPF
GId2NfHazcQ2dBsh1dbIz8HG6cnBk5yCDPBfkbMcPgfQuuNEyAMmFSwZM9HfHzLw
NnB0uMDImzO72det65ZEnJOfeoM6K3OHjeh7C4LIJbbng+l9PL6fIgxEq7FQasmO
tHiJ8nLr+4rBhUEBkvt0n/xv9wIinlvSfaVbU3k/miyqahy1WlYD7iX9l70YV1gU
tWmj7+s+yFs2JGD6zcxU53/06s+25Wi86HSqqIQEauYsutrPawUP3F+x+o4zWRqo
VP1KyScnhPuex0vjnIQqs8Sjr4EqoBaLeqwpm1Hw4rFua6h4nRoWQfGK0nAtz0tu
eOytkRtGt2qnf/FwjuJLrrhdsftXv9T2Uz+mm2sAsQuMH0rta7N2n001pNrQmefm
3A8w5grE+f/7yeAZUKYx1BMa6zXjwVp+X6znVjGeTHneDwwqY7tgvrNGC/DZV6jc
/+7v7SiBSWVve/cOpDsDOLlOoy8QeQsZTS+U6Y8yCV4qeVqkT/iY7Neb5Ft8S6K3
8mwfRrrOnhE0FijAq8hjU7XJqNjTaS8HAooOa05XuYVo9tRFbVp41k6p2/so5hCM
iMcBxSLc6u4bPdS+u9hYOAu9i9smXZaa0WJ9iZA/E5wp5O6VBM34VntMPMfb/ZGi
n6WuiOktbG98A9/w+/FBbc6EuvYgXZZcfVPSq5Kh/eZUJ8rqp71iEsocw3D/cN5O
PaY88FCJRGMFMkYuQvhgLdJCauvOsm9R28iSxvDrdr0o0y/XclXkp1Xx/nDsg7xo
98YndYnHzBI/3RIFZrJVdovOkBYVMV40Sua0yTTkZ8bTMy8qYQGe087FhCDGxqOh
/RZ5HDnLgSceSHlvT9AjB4YFMgXNYaCxxxZtLBanrBNm55QAt7J86MwpcGbNO+PM
do9JAQJE8xCIFcOKNNQeWgWdu8Q50c9RrMPK7Ih0KDj+AoL0P/Ja0uz0y5wj5wDn
+rmq7JASl9sPyjJgyin3uMX+FC1W57V5Y1v7BDdfJ6YvILUYquOywClMO4tN+54d
eExf/RzLq5jzw7f9aktiTNl7yDy7su/ma1UpX0ONVy0RON8E+K5ykMq3jt6/tvrP
SI0rb0N/VrPq0HW4l/F8uQ7yf1l07KyIVzLgNAfkb+rEXKFi0mwny/95Vzs4hXc2
6xmlhJVyuvyJTEtSgQ1mIMQMjnQoUaGu7ljSCZqURlUt2Zq6w1wfNIfx2kkr6X3J
avRFYL4P6aYwULPW2LZyLpsd6KUHzqyUC2J+ccaU0gHGQlWK582ztsk2lsXSLK8f
Ik+7hmbDZ/mhB8zcOD2UPvZ33I/mx/rrEqTXY5gmMPmOLJFqFqxrxrv4giLCSKWI
IFf1mVrAILD4JFC634xcWwbjekehxTc2/aZRpMo2xkRAYadG3AadH+GibL/K7oJ/
jrBRuKKsa6BWzKIHLGt2PWlNAJwLRsDZeTaFq/3gAIGpjxe++qW5tlD4Joip3vqX
rb2G7Dxl9WIjyyF+JZtaTWvXApp4LJJgQxZhS4lbRJ3IGaaTrUmWm9f86/2oNkCb
gsCbRekrXlQVHNPt5UvrVW87jayxSaLl9LK+h6LGX/KHU7fXuqjChVWgDJzUE0UX
MgXhEXuxNNh1yjQlqkR7pjgE57A3q0oIADeXGYH8y64fipUHt3zSgHRgVcrJ7XIw
gMk1S5XimpHg1p86mqouiiS4k/cJetkyyRjWWzOGZYV4imNf8WHY33p61FyjQ+qM
wJdABGZRfBGMSuuFQBPWtxU3msKhpFKonqGOK58bepRUuAeGrXADJqDha1ow4ANi
ixup6LSZY3tq8uA9006p/k+29LDVVtyl98xcdFEg10X4J/QLFnNkRFBL8Cq9ICe0
+GHwN/2V+tJbIvk3gR635CD0KJPTe/tfa2349rRmgyb5xLP786e5/GnbhvwOEi+C
TFq/KecHh6wN/1QVaJIwHYvtmYHZbyXBfqlx3ITPo5iZn7V3+ekvU45xYK0KV9gy
Sk5pNK+F+NJPD7ii56pGxiokTYEks08UShLxQmvxgp0K50a8TCYLsM20rs3VqPdJ
fGIdvJ7G51s5ooPTqkgP1dOJ6Pv28oPa1D4zqyH4TB5g5IU4pUIdbpdaaOiYChYd
ifTcHSP3hQxuy7k4XkYRxkAu2GZew9fK5hefXaWuRAC9uxMghaGODoBBugPOSkFW
7LtXqiusqqF7JXg0pXSsYarj32DQ0e4962F8BmzyuYF+hvkAT8nCeSs7rttmiq29
pV4sTjwvIwiDLQeClxTeXcKMEFkRhrmddTHyPpGhhlB3Mf3Z79TZ5PoWFvMS6dLe
309aCm036Mop5oDgpIlPdSzFQdbaz6X48IAz9aMnbpkqLPkrRwMQS/J/o8eMdNfw
jUxl1WJ1vuu2pykLMi/ZfKoMip/KQrlH+X778RAWnY5LXDUZ0vV50/y+G3801fEl
gMF4eKI3f3Q/0w6t8qM/+WP8nPF8Uo+jaM9Lnn44Wml7tmLtNmnL5HxJBk3cgEJ0
yj6/2lcK4RoaCjnIaEW+pU/RDdv1ls4hkC66DBf3kWmdJrMR/y8QaRT977fQCF9l
1/ONI/3xqJbzeeE25SLITM23MHsA8LzjXq7wRnfYuvq6cBATs9FuhWfsDj5nRW5b
ZEr0+BkkyW7GGTvtqFIK/excRXtXIPk1Pgfl1McRvt0uScBLXg+U2ghITelUN7Os
krI9Vkqu0IFe387uJCVABJuYBYR07za/n0v3JFXlDNhWkxX3xryYbbfSg4z20CoF
H3LGeUMNUazWWYVZdje7NJpsFr8WiBLNngzKwAh8q/fWfXAZNBQ1eB8JXpT54P8t
PZ2axNOkndFtKrZnpkSQCEM/29TCHHXOlTrf9jdlaQheJsytx47Q8PCgI/3Z8JLJ
vXPQoLqdLjGtfkKbQAYknEIlBg9H5a8wY7ObragR6aP5SBI7XhRakfMIKYv2F6Cf
9Hk0/JUFcxioBOmGaOZPK0LYQdtNL13zQPAl+1R+t0Oq203vDOsT2dnbGp0ikjc6
BEPXyWKpF420M4gNK9OCpBkn0kEpnWOVAPQB4ISaTlOXr+aSIJnOfcHR5fOGpNnL
l0eQur8ZXTrXp9WUosaqAPGyGjot3410lwY7V4DerwPJuwoEZ6mSXSBtLwdo/qEm
gRWsgidaK59DLRSbpcuinw8926eRqLsvo7zlyYQfDJJ9lksj6KdLj4fGgHzW1AUa
reKeJciytRQLITwk7SK9rMW453rfxeUNinmx22OZytOdLdtxwCClBjy5w1jDpECG
CPjPI4e9wHuoBK+sCjzN8dx3hkEMZsOeFQBW9YKGj7IKZMyzmlo5t2wi7kt8Ayvo
sJxpJZ2wlQ7QHnNQgLeGCJXDj0rPlK5iWor128j1qSjb2xAWB3oy96OV5IEtNvHt
PEl6YWfqfv5gsjY9ioChPyNjuyYssaM4m00HTouDK5QUCdcCCbtnKysq0i/Mhysi
ROu1wJHukkxSgReptTi/Df9WC9dwyFPpVORvz+FyiskC3SKdn2jYY4FxB7RQ9vcy
Z2mZJzmBgtWYFPL5rrfcws35lWS9m1Oy6bok83loQWbs58iS/2J6vwt0/Tw/P2E3
UYlXhNH/1dJ/OC1WpdFShTAflbd1vnzsgG2ZPmQ+3XCBud4+VBBZTfyE+iwL/pci
8jambWYxEj7PzO8xhsv8vZltTqJMpdZ2W35y2Pm2ReCXVdbuPHhKKlgoPISdQNai
1DcqsBUY61rcBkzflk7eVf37RQKqd/ymYIIAzuWyCb6bC2PV063PXKHySD8q8fbL
FlCk3MgS1zVN3iPjXOs9w99efMiBXbXSahac1Ir/eZTSyXvRQPOT2R9jBB5yE/v6
8E40mZUAvePHxmJQq4cONCrYF3EvPsexFGmhGoib9BmFDCwKvAGBDz0qasF7alK1
PCs+z85Ve2MqCE1wkjvf89gJ37rjcHZtO8SYdFDsD/bc2cmh9i42R8kVj1ui8NJ4
pf7BgCg3MgH+0ItvNmW2Nsk+TIG+e+9f+eZky6pbBVzJ7evSGnaki5XpukcEHEuC
zIFmpOq0iw+7pv8p+uxcX0k0aR9RqKtUfLzat8TmTX4o7FZvFy6m8CxyCMLotk4O
cRWfktlIigjWbJPW/DBU5oTMPAWqKiPcJvlP84WYgfMwvq2/UZx/DeeHOJA07Ao4
TdQtl45qNyP6aGi8yTdaEQ9TSHs4GiBOO123RLg7pjo3uODxMo8wEf8ztJdxAntw
irXPeaDr+ikiTmvdWdGTFN5CxgGwz42GGk/mpuYMcUU2FyPVWYylQz9Q6Tgh7eX3
VeZdYAR+CxRYSwlDB1aFDZYtbn4OQcS/yOb58vC3KyOY/qgcIWl74L2Re4D+pRm4
6MxIpc2Tttd2RoyQgQBL7P8VdHdmHUfs893tApqvQKgD6aVMr9ZEvhxPhvxKPU1u
LlEYcp3ydToALgJIXYfy0Mqu5qhmcUInmjG24KgrNLEx4w7xQ2SzLTh4WqMECqfN
L557b7e3O5BRJr0XS6hJtJVZnGI6TrRCKJWOcscWlx8QXoKF0qEUREGKrVhygIm9
ukzCobaYUrXqlRuugHfA4Wk4XIIjiFrgWm2zz+bkz3ZHgC1ZERtrcgejKWvi2WKp
Ub8t9J6a5pJfRMmbZn+GphFrrk9xB0JRstEg1ztFp0rsonJuQzxWB5MAlm9fI8wM
UClBO4u6BtJVnhfiKz/tJGx9UilvclSesk2ASiwQlEMzNTA1MXsthSa1pB7VXOvX
9Az1kyuBFYja3UgSj/1EliS50953RWYw8NYsKbamX7UUVuZXsUCfTFqJhdUZdZgb
eQl0V9sDMMb9nc8fM3CEDcggRYRdfDuKu7vLjHd40SImjoOjSu/stS9FBYO0mOQY
hr7LEKQg1f9YboaAmjCPufTKb/GpuR+7dRNwZNhCLpyo2Fq/1xh155Exoqd9juoR
ov+oUn5ri6YoAK7ab7vGBVqKA86VnVi0Jn7/wH4lEcE6l3wBWwWrAij5GI7dpbIL
xlwEiKgGC447vatRhXgpLaljhua+0ccg17ftnGJAV97JxzTSbHz3Uf1F+rk+HxGL
7i+gO1UsxwKR5A/1jdsWhm8d3MGRwzygJvAvOwX2DSj2TPx6/Y6YczFXMCYNca4b
EqAgf0TBhAV8WmwoQPER35YPvvyGWk4OkzSzKlrxD7X4gQdjwLR4xLo8TIRzzRQT
A0/lZ85O0M4/CqgXZIOU0w2dCIvJpELY+UPpOiqyrWvN4dVBOOO5u8XSKHAZTgJu
cwH1zSt1V7qH7WkqF9D6o4zom36wmMtgRIdTXJjPOf3itIM5b6pTYwQZf8DNNUUq
7ZWGAB+A/ImxjRiGuC7YGgbWxyxfyhv6b/6DprW6YENLYW+AQjRp48VbS49XepuW
KHvr7lKcxit8IoLJstA2w1VY4jfduANcVcPUpoGzzcGmG/Sjrk5JYJoQeSP9Zgdw
21Zr2IvR6r3YVWLXU/tbCbZMrO9dj2zMl1U4va6e/YjR05Rw0hPEbSuah8J6v77e
utxnK5jQ/LTFLzNuYyJrHFyQJkMa342u53/vjzDc2lUf3k9w2OgDkUUZcjU8bqyh
Em/Z28M181kD0ZR/SqwVTvInz7DewreLcs6wYz1cgKV7OTruj+J07D1JaSKze7H4
uO0tcfTTwl1JE0mJ3X2aiZEMEwz3es8lnNRvysRKpjkEhHJ0xOxTHL9h6jA5YV+W
j1xC/3p0LbV5Lp5Iegn8JwUYRHXzAxB//sGWO1Yn144da6rGJWQmlxZABhFdJWPo
jONWYqWipJIji0dRs6ulNSOFFnK12+WNl9DVlh5OoIQuMthm8p2QeWBwn335uXgo
EHUsCxG3x7wZMzOYMiNBayMsK4pWQtVdMa/ylLX5QIraqd8Q3RjpMbI7Y555OpT3
7GxqM8LZKYijf/aJyCNJLEUedOe8WBFCZ4wz7ulZ4K4SXf0ltLXXDVnTiILssAr+
6OlvRltQSWsgvhdPqv40hLJwnirH5EKDE2m91Z0WjBMPGOPkTj+jv6xESMxtC6rz
SeisT8OIn0gsw+DwaWZ/20eZeQS0zEPftV4YAMBTEWtBbE0KR9ZfkQyaWnkxToqL
8BHTrGyHOt9uSwJwCzUA0eQi2UI80zFVbEWLllXqovGLxje/40ZrSqdmC4fEst6H
h66Vk5TYvd1QCTnvcMvOAjvcJfR7myR+qeDqxGxnJBoDoDyj5GweU04i5u1qu/oy
w2xg3H4fNRepQlanYGmDRo9Duq0ehjUCMyDRr/xD3Ans5FGeh67FzlGFnNu1cbqT
YXWKs4I9UvjLNlenGbyQvcAlfL3xKUKuz7iome2UNlxNr6VAvAODs68Q+b87olm4
NvnHiDk55Tu65FhEL4ALpI4BiVDBvs+y31QKRhC1dAz3h8JiHoE9Aa1upDtaGII9
Q2D0SutWcI6SEtqV61BIi/8DrQkDj/e9HAE5OBAsEqXpAq1RHKwmgZEWMdRZH3Oe
VWf510SnOaiyzqmNSXW4GntaBRDgGhCSPqyQ8dgqAXLuTL4631FHj7ooOSHESecn
bgS8k1+n+SuXe4MBXN258iqQoTLGhgcwX7vNwDqUEZ8KrpJKahNdB93tLdC9UD8+
lhOULd14h2sxmJtM0koe7LEDekdPu+2VVPSeKfj089XkY4OF2Z5LwlNYEmfxNyb9
b9BXdxIf59R9VrSF5s8Jc4L83INkHzl/JiSQl7QdhDDqZwLwQuhlZGce2sF3MWha
WrRSQwIkufuVIGIrhvopXpiRYa6iwlLMpweon9BuR6+kx9K8axHPIV087p1vNbvL
/8Wszwwxt36AjxBfu7lLZ7PqoG1K2PGxQ3rVNBuZU1b86XXa2afroea1OcGzehuN
2+ckpCPZWCIC2uCx6hz+xWfahURFfpdE1eyHE9bJMVT0qIK2akzu3WkKpCO8uHl1
7c9j1OvEJxVonbr8SP7zs+mrhSazc3Uks5GgcVgY9UlbP7xeUjUfZYBwRCM0M5vd
AgoZoZenJfAgV9gPuh/yNXS5yt+J9sdqzpdvdUIIE/VbcXsMJrGuskDrYSwHOSIz
dkwFja7KRS5iO6v1d/Jd5luWKlwot8XI6XDHbq6IQzQQJyZ5mO+Rwu2gaY0Pxy+5
VVf1lhjGiZ/kjPI5TBvahALTIR8JjZ04UCVX+gz0GX6GPyX40D4/gqmkmZVNTIS4
p+sMbCPwsHBSyerG1QuxptBSQl4NHKdHOzaTne2n9E1MuYFBfD0+ntkEFEA9+m1T
h4kg2jZ2huG6ytjtAYluYIY1hqXXqGgQCFZkTI34u9wuG7oTo5zY9yz3hy1FXgJS
/Zu2YgN7uG0T39fW+VY7SmlcS/dt5S6gRNXB+f4cSymUXayZEFRAnbLPLiOp1zOM
mPTeDWywC6QNP1YUWRB9SVINcLh5gQ7cE4N0vYiV+2cR7EFbKHqzTNIYRSEZQEym
4qvucF7yob/HCpoZux7ygyixH+wqnFjDYEAUwOgNHBgos+N0yTjjYd2ypdobseSK
kgXDAa7ypL/Q4aw+QqIi96GGkPfm3iTZ8wGdSJzvJOOnb5rPw+wNyyCx03+KNXwk
xyINKi1izLbFeUJPHCBU5WbFcF+sy1v4c94N/EkzQAgArNy341bzf5RPfQzgug5I
r57QATslHgefByZDECBvvsR7KBKLHugaW6FwPoO6xrRjczZKgtWX22hgLx0+QsSd
O6XB7rPKlZB8Yezy1Vrk/iLi8as+APQ1zhgR6A2GuT3r72mKVTwoE5MArTOIEV7/
+4txdvByzoR0+TFlydqYJqA5bYJqbCJThjipMPg5/wqqgJxUV8j/cwLqUDT+hOIi
9FFRnmoBkHbrf+32w9j4e6vGe6dU54AQg38/T0n+xo3NK5sI0Zyt3ZxBEWZ8vvfS
QxQyxRptq6kg26LfSow9PmFlE83jILROC/cIf7B0A3cVp6n21WGCI11BFgTHULWw
V7NYOylvKP7zouI936n+bmhOqpXdoJjPB47deZcFhEf3xqjr9inGx0dcRLbPPYzv
rMXzURGaeupFStlPVNXrliF56VTrcXULxfbNnFDP8INM7SMogjmS2Di9r3+JXlPR
5opX21ij1EUCgDl7xbteB9f04sWTbM5Ph9nOfxPzcGsIhLU1XAYUtQHUjUMGEEln
7BVAlb1EVg5StXbmOLzzXS7KEIuWHD+313KQxi6GSslVZYzNq6+/c80n/1Zcps5J
+Ru/DulEnfzYVrLz4dLo3uHwFfTO+3icL6MRBAoq/Ls+qTvCYZEvaserSqhXbNFs
Sz7ux/TXPhYgZL8LEoTfudKZpQpmPjAKe+QSp9eKGwKmZZkZmITj5uDnrCyNUUAt
aAVHmSjn8dbMWTEfaCIYmpZBWNJvsu7ZQMqxEnImxkdKHnV53HG0MnC8HJk47KPV
cOXB03re86D6Zy8+vsqHcjjxESectIRDDusWRBTVDA9mtUxxmRAKrxZ3J3O6lD9D
j3+QCKHha6GlIHa8hb0QfrJmYZWOu79zaseVqI4X4ziCYxaiQOB47vR7wuWidZnl
Z3EtrA+4G7+zEGE434ao4y97q1YwOjaDjs/1cmHRyVfi8yeH9LGk1YgpLHXjd66W
TXnUH670zsT51pwiOZjN1SQgB4iaNJZP6MYay5gLAWF5u/dJQuSHo0tvK0D0feEE
u3IJRJo7TmwrGZWN2zwa4ZNJNOSVLZ7MbH1hrQeJ+IeuVtqzgI0t9PGScvUk4LSL
l5qi3bdqrorGqNxvWSGBG+FiOHRGz2reti7e+RzDOW6dhh6IAEAdFuf8v/zYSHI3
fInwcLTNqXNd6tshPI0cKnU3o46saNbXlQ+WA0nMKDrp+7KBcYC8nbi1n1hpwPv2
gt0hzsx4Rju1Hyh/+5BDm2hCh4xgJBmIYJ016dIwUJ7l3UcWIjI7rPqfVCGjsEbJ
JoNFVqRPQ6EEx0HWjZJKUFW2QlJUcGw7G37sC1+hXoBvapwy0mpUxQ9WNlJTS4Jx
Ej/E/ICHH2MC2a4lMuOZPynjjHdkdmIF6gmfP252eRLu/fXFB50/hB+sEekNm3Ad
dJ+lTm0swmLpSzH/Owv/Rx1eAQGvTMAG4ilWW0AuFWyLbfTbd5zsP5clBU+IUeJO
4jlSsbFzA/2K3Q57s3I8LQqeJwmIBM4aVmvqbKUwOZhJwjtFCaJnSBnz0k02ACbh
C7C+uHxpjp+4hALHKwgl2hZaQBqHzv8N4PeqSa5Qj/8DtW64dbevLXEz7DXIEs2/
K6oG3dz6l2KRBT72aL7JGUR/ERTOJZcRsD32MFXrXveh4obLAKSSM3H2sDLTCaYz
sf38yhtJodh/2/AKPMPsdddO3WCFoAWmmmSqe2Hx7ath5XDWm+8/fR7IH90Zx8hm
LuplM/2i8XnAv7R5OdmMQ/vbVRoIMftuPZEkDfY7FOPrwnBrh4tEV9epCj+efcGU
QMpJKTFNJ04EAScMPkjC5RB6LYF3nDkQylsLzyZHUf8KgJWrzk2PiHNgvek92maN
ExcuMDtOILGMU6hMUPeFZuJGLGMQcNfWVOtvH3CtQSztXbM/jkKOxLDoyN6CovEn
LEc1jiALRE6VxKn138Xxzv5wA3nNWHZ5f1u6RCo0byOOdyj9+8r0dlTr7DrJ30+r
g1TsKs0EvLT6UXlCHMAARnub7n5SMkZ2uz/+eBBgIwFsa4ANsPiDGdOGdsm0bk6G
pQBpRDNPSSzmhzeMDF3zHRtLs41IvCwXz1H3d/GI1PaCQIWEPgvH3QAO6mfSAbtc
UtV15DRX0GmcxmbX2qNZgN0xMCDaDwgpk9IQxyD6wY3zQqJS9gQJd+XrOyeb9yCZ
FCIhPnqzeUKNnDNNtAPaOA0tYBWMq+aWE9A9jIDN5o921fX98f9V0ECOQlgojiNJ
sD5flH/RfXZbZ9RG52YTRGK6bBWXjgbGeA4ALaW8Ec3gY3oKozUfgrMuUxh47Ch+
kK4FdFbw4aQMwENvgXMiMACSWTsr9MMk/C58hTcxVHQiT4lXtFHO/XXiKiBRLpEN
AiHQ2YlOL2ZOUxJ5AU/8WX/OZDXyvNbH93Rzc+gyvhsGwtrs8dw3Y7jFUQoGp0TX
AYpwRJj5+xDvf2GPNmQJzp+ee2Sc9r/r4N0J1uhs1UneYQb8IpXrpVsoeWw5DcUL
+GqWa9vT6PAjMD3vl8IxNarQROj2vdkPzu6LiBsDXxSnmAsLB1wm0kgVV1BJLznF
qaeMKgPKpHNKl1vbIP2PihFmeW2AKwTCjPmF1DM6JsCP3Gp+MveBHwSaUG+IZaj3
c8I2vZS3lyRBe13YUqIoHo19lJlquu3iNIQZUBvDXgkQ8X7g0HqD7ThCdxK1dE4c
Mp3KZ55UmraHtOKQZhdtP8SBbfCdShNF+odneDzEEIHVpbwFqzp00gz13WdYOX3d
jpnEAYNnIuZIDaI3GAJGKklnNWTf9nj9Ab7OAL0IAew7ykO3u1hA+3SGDZHrnF/l
RfNkKW/zYEpuMC2uDyeYNsk+zHj+cVvsh8AUXSPTpnx3DR2AmiE5DG1B/l5EqAmm
BaUU+dh3sBcz1I38fLFyxEg0gMmFaBR96a7MjDaPo4KDn/Xa3pSfAocGjy7CE1Ko
nJj/iQNCmfHyS22shryMdClJrEOBUulLBzPGcUPZzVzGGSZZfATB2y8SCXF2MLrE
NLncGaR+cpg8GNQSVfNbLkTXj2JWnt0VEGn6zSTY6qCC8Oc/Q/z67SiD/HcuKvA7
+JFOaMqWMxJA5qWmsTmKiLN7B9t4ZaISZXdAGvAHQOQC2FtQK+8oRtmx7Dsn+Bmm
FIW5rJNMJ6XZQQVqzF8jd74GgjtpIYhz9dsuFbNUnDHfHEE9aTZp6Apjr8UKcI7X
KUfiKLYD5JpG8Q8WETPNu9I/aHq+2r3g9l89awfsz/sASMYIaNywWFUIADcM3w4w
aHY7Wc6IzHLtcLWV8Xspm4wTt9Q0ZdL/gDYnLsRnxDeZ4fints7eG0tGx7jXK/rF
+oukoYvqVwoV/JxsgrLxVk6lyy23O5QfX4/gvTWbdGBe6o/SPAq8jpy/zJAb6ZTV
kakmh5OQu4ucj6ZGPAY10yLVS3fXAPlu38LBPQdqlaifhZ5MIIwuUWB79+VTs9+q
8c0QjdLBCsH84tFAn55A5YzxOdqmtvtILO2nnHeiquijl2KlN1LPVfomZF3P+Zal
E+rzTj48xTi1Veof56zKQtCVgnxRW6IU0Ja9Rugtd0ywU9uk9WioIhK6XvrBue83
Qskgg5TkAhpXrw7sjgLpU0hipegJeAYG9IS2Mc4KQAOQzdYtPZSybS0Cu8JkGt+D
KV5bHH4U/TOaX1q6L8MmBFjAITOD/wonIONyj0Z5PYZ/NtMHO+U7mRYSJiJzfrfE
MXUPR5i4LIvBAJgTg+wi6YwWfXXqAwCgU5+HqM8aYBgkaYe0BCI8lzMpXLBpGFe9
fTNyntirAw94BNRrCCGqISA9x8zORhD5imqeu7uL1HwoPH1D7VKHZFCoU3eQgYZ/
oap56CD0yW0OZN1D91NgwfOrIW+myMbMM5FTFn4hYiyibTM6joeBGI+BcZq7SLBE
k8CBqd6Y2sN8dIPzR48IMltIy/SD6v75WV+ZXNv9K51YoPwsGm3WbPwliU4zjDSR
UkEWvPtIVWsM7oFQH0TIyG4RV06dflAH0lR0eDs55/9dinVk+4K7JFHosej1G2x8
z2hGNeI5isYIvWkOh6lbWBWpeBOnETXbBdGLFwbSAksEUkz5eTPX176j9ouUcyKI
yGhxmL6OiG/C+w9aHErb95NqRmTxo8k9XOkcGEs3AdjSnutso31+VM/fNsy2Msuv
3lTPHHzdo0QHqfIIBMOjkWemoeWIxIxkDW7HU+jwXuGyNABPy6KYyOJg/oRS/OjC
smdYKE2iWJOYkvFMV5i2UcX7v8OJN3tN9ez/LoXtngCa/RuCbLETqgZhlEnvjKvV
fZu7XGraHnhV3CjNbGUsmq0w4UJlOg44JJEU70zXp6+ok0d/A4R9P6jWXsWMWemk
CbbHmQztvpCtn/yYiuanHsjxvZx8njfimwrRrkpqFfcOAnbZy/fmU6T1xlnUV64a
heIr9l0LiuSmnm1lGs0PKw+QS08AEsIj5ykcI16EI10uma9odTyvOFHptdMRq8Mu
SG0ewqPBQ5/NnLuOjfkiXdf7FV+aT6yAAY5aaMDrO3AjDIqx8P+tnhmA5DgGy+Ka
qm1OKdmIfx7eglvxgIuPiR8W/Uw+L8OEYlus5EcefAhtCjlf7U6IzNiGD6VHhDrW
ob2NEyn32KDJ9Bdpe/tXZZKamuT/pXU4Slizl2iCNMzdJsaZWlFbm3P7wUNT536I
ikO8JFclu44d6Q5vWG6HhcOY998iTQ8vApPaBGhAoN4+bLjBHWUPrZOi6IX/R9TQ
uWZE1MlPevVLuTq+GhiLnZdRyHiTzZvXUjsBpuO3vgZ19hFOeEL8862KdygC8Iib
hxFXshmojqYdNNjDKufDV1oCpXDDwCaCU7HWbUnI6JZo7iEZY1FFzW7wIr39UatW
CqI5oZ+JZAE8gUJF2VYvg71qMVD3ObgUaU+q81SffDmirrmC7S6NNeJK5QVJF/FY
oq+BsZ4E3GLpaydke/j8sTzoG+uElI5vu8prLl4iwru7IXu1BSaJ6JzfnN6HUW1V
kr8QLF14lkIcBeJQnHIhM0AgR1rXVkyLdRYQlLGJIDgiW/AQ05T5RU52FjV5rVAM
x4AE+RWgvZdvjMd88xDeYZbAOBkCilf3ZowwPErl2eWzTFsY+OA4Vn558qKXtyb+
0xasPTFCroXNdOs4fIr0Ur7REtNfoqNrFgh/lqR0rSeA+RuGrduuFfdrw/iFW3np
UUvw3vlsfpQYCVDW/XLtF8O/UsrmCi9oImCBwJjho/STd5lKacotYlp+qoYQAzTP
Vz++4i3wQI1bzwm85tWGdlY4USreSVBpo36bpMdUGCQ8fouxY3kbkOwWe/dsxxc0
bcH7PLqcF8Ve9AJBe/oLiIoFToRagT/AOXkEvarLf2W4EwWqjYL70M+FgyijhV6y
+AgkKUgoNL9RfyvCp5JDy7Uhsr746kQ1iHMEyFVpIApXtlQxJs68tRtkCCJuf62O
Pmvu5DWxVKaE4Ud8B5ABSIzTsCx5zzIyEyEQfbL0GESKRetQQfj5n5ZaA+F0wIXL
QHBLQIXpkp0D0L6e8qYazStpjOTlOLg6qBbHim9HWViQCHrIhAH6OfiXpxyAQ+f7
tl4x38olWX5CrUuc9WXuIFNFq7O9z7tjICZG2RFaCRFdNN/Z8EixfN999vX8nyx5
0HHJlAMdv7VOsqux6RIvw1J320PY22LqkLa6Kdd9oy2daSNc9wvdKlkTR7JZI6O0
GB0K68BXLsXPASSHr337Um847tqW7SGKb8Al20vM2N8xpFl1TFpY2wg8ZsYxTzpa
voMp2oPYM7A5JX2cNRNlmBVDATV7V7N8zHMB6Phio4P9UxanqVFo8an3zsOcrEyM
wSZJvgvt/uCiZJFxcSqCNaYaX2fjZOoFjZg0yWtDGzNgnyPERKKFxztmhF5dlDbu
UuqEF1ureMUqWBT/fTmLM5dzNwNcP6v2548clsD098qi6ow+SUaeWyhFRDSFd5ku
JjYtO0rr1LqEiyf4D3hBdETKfF2SgfHU/hsC8iSDXU1FjoZA1k4CoMaRLi01n1k9
xe7BsYWgmoDJG0cKsdy58R9m3SD1LoXG33Grb3vB2+chkZRjWR2Y64/gM8wYdWcd
5tktcSjR9kK2mzLbECsRA4KFlv7MgYvX4dKvYlN1wj1sTwma9lV0HLWPFYiiCezS
8cm+HiNFMo3j/pHqCd7x1spohXxvKPkLVWNHKBaR7MmsQb94/1tQcb6yAw1kTKKg
jZCfrQEBTEV2gF18hHe5/yZaWL5M2BQ2xSa+K3igczr/VmdJ7ISGvguB4YXX9VNH
wC6woiY/zbLsxk62waNa1TdxT9qfAVf8PriBRWBryyJuq81gj0TMSJm0CINAmNdC
cIeQcWdjYSLl5DTScHaDTLjOJ0g+DUY/x6yuKsU1jMy8tAnLsJgX+tRZShWzJk31
XSabvdq4eG8XeevK9DzF8w/HUQYBaodagSuUZkVNGbi/sBNEW8b8XltmvJU3iWIa
+7TcJE3eBZHrI4Zr/0yzaohrw7rhOiMAnxn6Kd8Wslar9kLXnUmn644hBZIk22id
CwP1NybJcwJf0wCnxzvtNUvt2HIBgrwRA3J7FANosyYjqIubWUiooH0/8DB2KX4C
vUt7Y9qjB20gGuzZXyYbtbfHpzJ+w7RqBqTn5cTmOyE2oeYs4mYPO487QI9iZ6PY
rHsDZ4BB8HW0GDdkSuk44FNh34fHTJC33gXaIbkm3Qwn6ryFnBolUCSlNTqmWhtx
Ogkgn9UGsBNEqBqyW+DG3pnXk4QQKz26lIRcBYUc7fwSR1ZCCCiY2zEarXut2IMw
7FUGcLJs84ihxZ8ebwjVv/XmfuVJpyepWSYWmD4GuWSr5G4baL7+G8ApczdttHsD
ZRyi2lSrMrzGZwO86ebEu1Ecl6uH9SpvofTaab6UJJcis8IfpOscNH3f1S30GSh/
APsz2zyyjQEuO+MBazrD0foXldJr7eaVEmxSUxdOK3+1c8M/ZeYYfYjJ17MI813g
CgyUyHpQBTMDtopa5aDn7GTEHKoMqt/MUO+Q6J0Qno5vjRC5C4npi+RsmH/WLXD6
1MDAxFFKfeArpB23YZVR0DE3TG4zX0TRImwOAFfL9I3rI+taYayHPEnpMQ65/2qw
1LpXXPKLvg0uba5wplNDTg1X/vSdr00s+THS8rBsw6rYO3LFGw5Iv3d6k2FKm6A0
+zUz4pCJL0qn1K4w6hPMHt8T/FZ4HVBDM8q85z5OZhMLgiwtV0sDEhevEhm7VKd7
pmSNQlk3WSpmw6vr518yjQChHU64vROvvLhEPVQiOlymUTIXXVZTMtpc3NDPk3qI
/N81aNt8ONAIiK5qz41iITibwIYWTZCBOgiDD4EBAa1z/pXf0TVaLAEq0IaS2JFG
i/QNRyh8oPY4Q30p2n4HSsLLOoe/H1rvE9JBDFLeXkWHWGHaAIh8WwNV+3k3n0s2
Xnv49CHjf/qJIVVoTxlgbAxjTBVcWBVgIR7kYjnGWptJUxmAxoC6bAZdISLtaM0F
NtmyV3qhcIg7sHXQq9S3Ljr83Kw/4hWjqCe7l94uMX+i8uvCIOAnMk/aPuil5aOB
qjbCbuojPNMw9cetfBVG292RrXshfjL0M0+d4qXQPdz5lQ/e+D+3UaZzNZoEQTyT
bx79/OoMMtglWvOIna9vzONNniLQmECi8oPC4jdlZM8C7nTOoEE11xEtFsuhNRfo
iAzNfveDHTmJFQXK/2NBsjXVwpmzzJ0sxb19cquLgS/UCEzt7l5NiNQb1DLpO57q
JHTvfvYLP93QX1zISj68nP5+UfHR9z68DrJrasqTsV1VugyP1tGbiEH8PLsvnS6c
jo2qtRK7s2DNKchYcFcRvbiHS6JKU1nWsfUdZjE7tT9HXUMzBVikkRrJnabj/h3F
qewqUu7BWlax3lUWj+2bnFKS3D1szW75Ykj3eOtzUjndErquuIvsVz1+LcPgPtTk
Dl/J6qUvqylcwTVNmho43c2sFgO4281Xq1y0RYg7oNtpxfy7+5pNwtBNxvo6juMV
xEp/GO3fL/SrOhXWbT4umY50FCfPQcaSjGXHEs4FYqIYIlpbv4KLsmK8Tl2zEHhh
q7L8AicfREGUphQrLZy1ddwMj/oXYXXr9laoVNvMosPcfAQpjAqDldYnGQ/ssrSD
3YXDSCS+Ini2/i+zOYcq3cOl0GU8clGUCsJutXJDzymteaA8Mx0/2+Upwqdz4Lz+
PQfKfjUMitOUi3iQindqq9fMP5RtYTZS+OwuPao+CpCswvsgUlZcceJKCemgU+Y/
HO8rDwN9t3a3z3b0sosErOXC4X3lQxqXJfWZigXC3WyAhKbR55XtYmKKeNQGgK2s
PaQSm3CEVmreChiDXzb9BqsuRjpBDI3auxSgbde6tEZguuKB2rCK20oxi/ZCXP1c
Miw/cjNKEdaabcJFrN0b2imBSK8/ivLplbVPJa6MnXzNIh9xbVuB9pzur4UC72FX
XC3vG/48rmHcRvU6hgSvl+AKTcy7mbcXmQfed2DtmvT2+uEl+PQuJ8autbbc652R
OmWDKgrGsGszBUQpn8hm4WbvrYSK7yKqiNRKVXRxJgq0PTYc4GQCXsEoCz4bikdV
je7GUGPpqWw7VjGo8YThH191OrKHS1tsKg5IUdNnqsTdAwiErg+6BKvv9NSU5lNR
CUbe1vlBuzkJn8PuS0iPyL/coNxMXwjz5UT1roigyQDaHeOGDl0jRpE8f3oY5Wn8
CefyZYXG2aiu5+b5/EV5LUbyO6BD328AdVGEha1UmoR4pa+Wes1VibDFaByFb1e3
6TbOSx2AqaZTA1zlhaWu0blaT2ppo5lQUvco62+fgAcB16bQwFmxtwgLxX7a5NsO
V55qJNXrDvWjCplMyNCblyEk8PF8MQP95ZVK0IjnNca16zo861X1sydKmx2HlEYy
eqPJSiUM9EIX7E4EhfddfR3Cca4NyqUa0bWLOSNHBwH7FgVo5B9W3XDqrlbr0YjE
M9S1p/8Se44pt4oALfM4uvk896LMaeixCNmEbAC9Gtsbt5U3r4LqrxxtCMq4Zuob
XBYFIpXy2iiaGvhAeHfpi8y5vMybx5HMCVB/pGF0npz0p+IA0Z70JmyuscXxevKr
6Z7ryYdVceSjCgKjLfCeN+mIoR3A+HQXaOPZjcCXji3/S3yePyqJN31uqoPTi5AC
6uqjGHXeoItoqTq3lPss4JMsg05uvSmBnYyLoZPkLSpHDfjr9wO63e5mwixRmzIE
BoqeWf4mj0iDuqjioli4ANibLevynxtEir0jWX+GI9bqfC5nv1FJJsdF0PjF1IHM
ssQnJMVlvtz52YlAEKR6GA5ws5pGjEh0KcZ7ET6spDPGcT1Pu2L0IauglS/C3/bN
TQ6q/2ftrDhQtcUkeK97fkt3gR5KlU7t3bdKo4sl3/P/I/8T1rv1RpgibP95Ibgf
TOCDb/MVYFO2+awe4F05+LNkQaPa4n/SLwKPpLksjw762/BYdM5/1kWWMic9f7Qr
VyOCmL6IyhkotFqHEIEhL6WAsemJcBMXSmGxFmPbBygRsnNxYUkx9oQdQuwjjZhc
bMqDwnwStgWa1Gw6SZ22AuF8M8QvR7voYNhpH/Xro3VEmxo6xqzwO47y+nnV6kwR
vL5YgzN5QFqs2j4f5bEaGmNLNayPT2EszqcGhNRZJyzZM9ljhqIVS+DgqgGUGgmu
/u2y/E1Gj2uNWqiN1H11owqm15++WM3NyH0ekOva0sEUExdi7LYtjltElaKWvs+W
U6z2e1MfA5jtRocR12ok+Ni92S7SC04MoFe6hIE00q0eDRbWNj9xBVGCL7MBG+qv
b+UWKOU20i5u1HpBCxnHQk9QOFBOxyRpgGOYF5uhzxc9tlImeAuZK/gHZvQIL3Ye
9AZhP5X8JNWYakNm7cB+l3fjzbF8nz2krL+C7PFRdogfRTjRtnUYpxtnl5wLBYXF
wCtza5fLBB1RHfF/iVXQKaT4X2oqQeBYJUOTy7ZfId9YboAr8ml7gRIqc2BXgdz1
Wyic3FUn5Wp2T3fSP1mn/sGZbbrTLF2poJiAijxJigBxvpkjiYTuOjI5JD3wGxcV
6VAuDOBN/uvpodUjl0deN90XdiozdCtEkcYLf3uWUWUt/fySZEPDNyQJpAmQ0FL1
wpMBNT6YSdJoWXR1fzo7zzyYGizikBn/eVbPX65DS9TokaFcoYk16W4r3Q/SnCjW
NTnezyg3ECbT584q+is9Qe3MACrUsg+uVXSRFxe0rUioG75cETx4n6iqQH3wh2R/
bC1Rqtw1CgWDkRQpwR4Kf2FB0/0orvj5bfdIZHL6qYgTwyt7jF87VevatJ9vnFsS
XUqHsqouR1HG+ED2Gc6GIkW6fPdbz2evzoNVvvfpnVFe7uxca9gJJDK/Qqwm5vPM
v/qvTAKw+CaTE+uvtYq69hCKwYDGuJrD2w7mUWUE+jY7UKKgr904whRnazsQPv4V
WQJf08nKBZwTbp4vmKoPUY/dgx6Q3cNpYvMZZSxNVssEwd1bq/P5I+tB2mR8d/76
VrUrfV91X6JnyMTDCBudWXO+pKH365mfB5NDVv7uBlqczNZcTvZzPdt/d45PtHch
23ugrUeXsBE9dQGHFEPZ/wGP43qcy3q4/lPnlREwl8xSsxR1xfQjU9sDfRoituTk
5dY25yoDX2r7qM8BFuMG+9zrmkMkqs/Y5YyPFbsyp33WKcCrgD+ZDp9+xQpWnkWD
2vxYaD+WciIf2cb6inp+pEJ4BIDvh7IMTPrlwX+Pb9vifU8xhwdobgGm3Kpfd+qA
s17cX/Hj2TfokSj3Nt9jaQ1JmzOo4sbV1siYwnrAAJU8LFPDoGEbMHSf2NKWatHb
8WhyGUbTPagb9SQVTMAGfdSWW3IDfY/NnzwM2einFCjRMIeVwzO6Cbd7ouhw2JeN
jI6asQ7FK2+LFe80ijNO/GWPTVNLxcjc5lRWr/GemTv4oFPU3YmcLEFqFE98iGJO
fGaYIUnw5vd8Sz7UQSz9514FeVxlbmDhW+YVbZSNiCCsZIRgYfVoyFnyGQSs97g/
qGHLPmUVbRUhVnS+grVlEdmR+6vUx/BmJbXkMLuNxSL9nJhTPy7ARQyxz2O9WOQP
zF/r2j31IRhTKtks1nKTlmBi2lZbpEcCqEuXKDyIIEgxaZc2eB2mTVptLKl789XQ
NRExeV8y6PF0VHpR159kBOYHRhJcLxY/QiE7T1vcTUB6rDXm89XEYbTvcvmZAvk4
qN4Ri9sBKbkqx/CofaCgR0ukV+888UC6zIgCd+X/7j1CLWtHZDpCoODNy+urBolx
A4PP7Z7RIxZkY49Uzho72vj6gh7ipfrpfU+d+qviDx9CyVo8tfzWJZqAkLD5JbWF
PTpYcs/GGl8MecIz24tcW6WZZ45OsIKWkwdezGyq3hURShrh3jR3zNPoH8mKCRBh
jVPjHSYEWCaB3AhMy2OKy+bpuzFBu9iebPFHeQ9GUXN25G2KNgOAM9tKJ7AHW9dP
lOJKSMP/aeUqtCs7rjtNrHnlJF/83fDk5vkuewOs2jJ4S5yYfGNjzbAFfIUpD+Gz
ST/Oe9TVzDel/ZAg8t+kWFWu+7iSei+N/NGP5TxXPtxavS7Zu3T9DzFX+3PKqyko
1c5bw0dqsyl7AIaYgUX0rdnMetqZAhXt3b4246PUI2m5RunJbJUoioeI/F+UNg7w
FOqDX/PLqIb9MxFLjBz8ZuyaOs1C5qjPxRrT8bTwFDm4vaf0vBce4+Smwvce9cta
EwcJp2eiS7NbXrXayQkwfGyAIAFbKOu1oFzmovnD98Qb3EZXe1DotOURqiIc/1Kx
aM8mwUXjLrwnI9e2YX8ZFy1iQEMUb2Uo0syXeQhebb2aOsDO67P33thHwMM6nY3Q
OiGpqegRuwrLTB77D6WXRta1TZ4Pk7XQsgdOTc8tORLROJiFNmlHwlTiGbaAqCJH
Di/yg+bC0f6hp4Lz+eJX1wBEXpE78BLX5yrpqjYzUlEl7yflkcJl6dH4D78Vubor
ZdayybbXavsKPd8ifDptiSaS8uj3oCwptupjtMJsQkAYC2L3r5dtlrealmgugODb
nSWsMIgaxCyl55E+q9brdfMWYY5QYJM8ldSb5tHNJyN+Y/Nqr2nN9PRqZdm+oRTF
JFXD/yn0MrwN+MLwQbphZUSHQQDy7Omie4PKO5uS6r01s9Bf11UNVjEh9Qoig2Rm
n8o0X9lWdyYewNcul4RjHTxZwCD/2lb07igxHtGu3bEDiHLaHIJBzoxwVM3KYnuu
ej8kAjHzIj9kRJVtdaUTalKJq036XXbRTAnIL0EbSyfs+fRJsYhnYPuCw/uRNpYm
USVv1tXkCTPykFqnOODtaK3xS4Br9dLj7rq56+dPOaL06O+HwDxImvNFxHR2ef6j
fbnbtA2D4xstiTVl0MEyPRulfe51A/PWS3/QGLP8iusBz0pxSad7KtXRDbdr+2Q7
K2HeRQXXgtZrCnakf/Lv1AwHrqqu1B0DOLOLzwD9I3vEssFV5ADtEhyHBzbzQKTJ
eRIWf1qC2NQMAkCXGPq/0PrVBTPSgu9JLpOdAZ4NbITRL870CZY4BUld0w04DM4z
DS9fqvpgsGoKuV+LnFi/t1PhqwIL3yyUZnFUlfO2QKW842oXBLjErlnhvLMue9j8
g92Xv3lKWIbGuV5psM62g7z5EkDlFd9tPElRBI4IsyWv7RR5m/CiwSOwfUxsO6gO
2/r0/p1hBLxJ52FnPdlFM4sL7BALVlQkyVDHfdNXULN9Ci6OLjKSSHx/Z/3UO3uH
8QrqO3a3RDVYhFrj2eQeeW1Y26Mmrjqt5QgtSBYpChbT3QRNs2cmFpuEklYFlV+b
GNZxbzZCQkYgUzViFwEwVEnUkQ+ObdfudgFt1bUeE+ATBifJH26HLpNoMix6QzMV
lMSJ77i7yH1H6AxCeoDmZ4Kl175U6/huyjOm4XEogAL3pPDdvsvSSaiRuJX00uPv
Qr7B1NgpNtX8lpHBJxXrA1uMqsOnfO7DlNvtPr4gI938dLcGBX8GL581CXZmJMLZ
TqSzgAZc4umXk48LvMU43NicwVIhQ9R3WuKh1r4+Vv0bm72dC8AdE9kGD6+awwVV
u9QSu35zozuqKQHawn233B58H87zo+N2+YIrMlYATH9ye/MPPe3MQZWSv5yxeeG2
51X5avvhOLY+NFBNQspdut4AzPET4WECK6AdYUWmusy3qqpoPZliW8A0wqr8+AQL
xHffV7ynayHpGVXv9VR/B/beqNQznbRD+TpdlP96kLAtGENsVpqkMjHSOSrRYWqC
7CfqsHenWeW8dT3/4zCDkO8ughQ93M4pdOGxVYQTmX3B2EBVvLONKVWP4s6ywQTw
T1/bivD8XZ0gTupDqZwWLRpS1VwG54g1QG9+UzRTmg+PI6vxYeOHC9I7rG71aMcv
5FQOTHVCm7yiYkLNpfj3ou8jaGITPO3nwLrdLV3aIT7IZ4ccjR3liBAKa6IZvAv8
e6p4dvtpbb/AxcNQvKHluBGvdgf/Vyznoab0GBRPjdoF75YbdcAPyw2aNrGUZ8HF
tTXPNVNfVXeRCRgYQlK6JHPUq33Xldl485kXYbuaTm86EZK1IEDv0yu3ZrtHy7ZZ
A7E+PsECb5uBmPvKhuBFPYlCq3oesUBom702Dlradi/1qisrMvdaf3+6tkZPCEWu
rM9btdRO4FLJvmOcBUmkukusje5IejzB9Vk6J0G9fWW86YnSQ9oDEwTVpCEWvO52
uigcSjmQV0jHsAJ4KXS4DTiXoocl4RGq0A+plDLX8adC8B2g2jPIn4D0h3mxmGkw
ybQ3F3Q1rhg4PGYTTXqkUQyc/KBtg5Hm/CiNQEyKY6lZvbkRQV0fwMvtfCbLtcXw
jXETFsSg67/pbeg2JCMvDX/Yn1L+6B0rVbE38CIBMWuK8exZdRZZiMKunjQcMwWP
9jXy4qDbstefVlfH0HlDL2eADUHghtLGBGYmEAyQNd0FVydOoNr6LTaF2v2Kd0By
QVQwRhQShfL1xgJwOSxFOIDVn2RgobPcp5Dz1T10qcfC9jz85M/veFvespt/Kk9f
+X4rfYIC/BiuUFmFKc4v8WIhpHFSj+42UGqQtStD2OAsxR2EufJbgWwf2JbAtpCD
UZITF9vND3qaGHBtmwV+DWbI+sbpSyfWc3YrPyEXFJWBxSYSSW4iuR2WePkdOaeB
FH8Gx5455ZYtpGdEDZfap1XabiA2s9sN1BTmdXvgllvcHZtyAu/NSzTj3/zTgYac
I8iFQNsDaPgiEhzGNV2oGQh4P/6DTybujG+jUiEo5GaTP17XRGKiJDuwPZJwN4Bg
l1niYwk2Q0V2cmAgDQf4YJH5b5yoc/znYJIQxawiXb5BwDE2AzITThyrZ7XKG7pt
TBKX0G2IHJJ8uIPgddKIPVV2hnFMNmsXJQcdxjr1kDZ3kjHyF3PC9kBrlGL49V8v
wCP/gyPHNhm5MyUNuWjICAL4/jktRtDZ29V6CYiqZX39/lDSm9kDhF25fNf5RWzo
aTiuUuKgI48qkP7qHrjzyIlJS8QECMFisZZZH+zVj5AwecuDGDEYJgCVVhN4KzRv
aXOzdr/jlStx8pauuJyPKmecIhByUjbpm4dCrdDrgaZuoBtG4zv5mGeYVCGTZuif
i/INFxhCfAotup1k8l3F+f1T26YaTEQL0/6cv8Ed/b0MEJwx0IbjkeDZPSa8+9+p
1vwTJCwKtq/cDArEPT0O3QV/miG2+L+TnMuD5PbluBx+DCEw1ungMmnG6noBCGFL
VnhdmlGw8NcUweRVcIsVRE+twTFStcL44ESAU1P3rthdJBqOOApBgAxICEz8dEIc
FVBIOM46YprdYCXbXW/09beHa1ij3WGC0W9YJJR13eluCAXAHzPezOsmox6FFgzA
vt+dgil+slQTMjzkKofEwvAWVqnIcRZQOHyVOs5tKmsCheUd2W2b0USwZk5MHF7p
42H8Dw8B087AhosqWOe3bF3wH70DbvWBlh2YFYABJ4isLlI10skOvSLsEDGDvuQz
MdcabFGTY/Lr9YkMIAw0Z6lvYGBggroU4gTQTfm8HJ7Ggy0s4UkTNeI6Btr2EEmb
fBo0Pd3Py4cdL3n91NuGVuTafCmI1CnIBrmJGuuhIpoxTvLtU6wCIt6+Vo4vjx4z
Mrrmywci4dZlrkMjvNtPiDcQIp3D9qtzSg9KZhNzVALM3OGL6PjmXZzfiQMQkXZU
HBCkWxRiLjg1WueghCaZK5kNXkUepRoRPS32qYXtY7geedlmP86tlfAWaj34hszg
0BH6b9s9VwGmzvyICqPYWJjQQYkchI5td3ricCKOxUHFZKuo/cvXPdO17DtM2Zed
9xMAb+0bAq/IDT78gou54mkOfWEU9TRh/+69MSvTPoOgzV8bJfB3uXoSQsmp/bw1
/7NY/N2VULESuFCeiHvxsHp2HsKJUd+MXLqOzBoNMIGrj2faLSh7bPTr6dQ+O7wG
F0VYeOGq4QSoliM1XU+1kWkUi+xPm76B9j9MAB7d2kuHmRtMifSKaEJBoT7wa564
jHe0wZ5grU/w5erXWO+BpNKm/+m/w9nHBbR7cV/Ncs5nC5l3MVV2Rhs6ffMSvaE0
0SjjZusMBYOTUzusCE5OybgejFgg3u3ZZErZ0XwHO7HTgw3HC2dHNY9mq6q2P2E5
ZBT5+eiVOtfAXjdcJg/74aTOxMkH3j9slFKTvayQNnEmZETKF0vAFGPzDiBKPRrv
k60Kpw8j7W/lCA8/bHyWDgw0TJjokr++juWB+m+Ih3cf6tzKcQ8tM8aNdZJ88Vlm
gbd8ONiJYLK6Vh4HWtfHYcJI00YWHKUF5oCZIggJ2whF+ZOXoa+oEu4N/bMUvIgD
IudkU+QaIFMNWvZ+4ICB3mLy8MfN0D7nCia78bNYsFaWi3pDKl7RUxMHq8J7gv1U
BGS4uYmtrWCQqy3i9tAfBHRMxtNbfZKwu3/UkdMJJ1yPEwFnMjLSFpPHVwBBUohk
oyp/GFR53j5zTBLeBDYDaLrU7kqhDsDnheisYLn/l1MWK+pwBlXeoNqgT2rRcA9i
qbbr1ypbIOZLQrX8ht71a6jmfTFGGNCnyc7EMSVCE3mgI1uSApPn6qAEmOA3zWcA
KJKYQIcws8H2vz/ouq7aMLS90SaC7qvSoWMZqcpKTNiXE82Tm7C9crjwDNB5DHC3
o32G0g8szYkaQLe0WXgqm3IG/QKhmT6KpwpxLtMEFLGUHw1TNZ336by/sBOOJsR9
Fk/4C6xbQgG6cPBf1imAKuSe46Kcjlihrob+imfsQ9wzmV50AlBTdcpQ2onLW3Zl
dqIMqKkT871N9S2pGZajkBm6ZC/hZptAmXMBo7GIziizA3ILRpo/oRoXOALDvLUg
eGR65T4FRSxc1UmkFQ91CaMMWBvDPvDmTeO5dfxPl9P65cI1FrFqGJS0OPqKf3Up
dgWcODoAT0c0tHchqIqwlOAHEm3WXEaS4TsVkfUoNqtQFfJ5rSIIGU9GpaH1brgJ
/sNaDb+UJ3HThBMiKtywz5t8Gk6gjg1eu9VKoxv4VnyYfXuyJAOFJfSg1DiN3/cc
z9ZtSZTdQtCeC1JlncV4Rys9gOYe9/v3YxJ0PYlGdNmSiQnSHtTkUFEtIgW6O9il
E1QZJn1evgnpzItANfjYeH2ciTjTlnzv0dkWpKP5fQxsVqgYslrnXJfgZMqfXc8M
sGE9ipNOvsrl1V1InvKml1NB0w18EiWIjfEfJr59nFlj7XJYQUe1yh5XE/aGvptj
mnSvlNrZ6A1rCM0rdWJkE3zO37dpslojmaMD/A03gAqkrwtAWnGv+9nhl6/f5OyS
jaP2oNcseKAPcRYxuxLx1iIFHmI4mzBsHlYJe9C2Xk+79A2fK1aIjszSGkSJRFJC
w3kyXAT76Pgip/y5fCXUeSge3MIrpSjhhtKjfTSCIB99jA5IUx7mvQb/F5Ebr5rQ
bDKugGfFFgGtxovjuTIE3R6gHBESH2SFnEqk9OwHY9Z1goFcVvrTqoTxDw0AElJT
0oZA+gRGR9ZkVmskqZF69K/c3QMDTzNi8dah6qVrr4YfdpdtkTglrh44wUWFJtAx
slmjNB5+sCzsZV72/7fP0XElueiMBcQtHeBboZ8G1ziyCdMTnsjznPtVVpuffcW4
HtWBNMdwJTO5c4LQBgUdty2gcGyr7TGrI9yg3DsdiInhp72CsSIoN07r0oYqydaj
A347Nki9pgXBhzHW1/wnGQ1jbBBb9INMg/REp4mxKCU9PRIYnTgzksSWVkxMa6UC
VoVwDbANoJhMc/KC734qp8sU53T4oDJAjGj/MGdc86BK6wfZCsQYHTDL/7zDH5y6
ZyJK0mONsztW5hUZap/iwdlhYv8j0SSJnCqW3Gqs3pzsDDPDh7MfhoJ6OFzgbcbW
iEnn/5uQ8+S9DdaKxK1Vb1a88CaRsbaynAv1IUHbzgA6/zlJsiGWuU8OqGfn7rYa
wuxKp8A0UexaASJTG73FoRrBVorfkYYPLeh3iQwwhfdxLZ08bnoEhOuYjMc7UgX7
FdZHLauPs+kYKsXrhGcOP9dXTQnV7xwE6359CxlBppgIUlay2jJpI1N7Y1tc59p1
ikTRe8fv0aOJy6rdBY6zggcWkF7Meu4JotPMKpxdMya5DCam6kzWUpLxVWQdOojK
zdySg6jx1yM5V1SnXV+ZbxNXoVryhGlpUwEcvSBvEFq94h29AI/nFW5GUprNO9vz
MuTrpwk1U9FMfZniVc2JIGY0yIWsuFf9fAyVoYOGi78Zf8UUIxm39l2gzc6iYT4k
mry+FZ6E3TpDjkSCrKGYx+IMPwdX8DvXkDYR+BLdc5YwUUvYYdJ1sukR6/rYFcVj
49xNUA4QAEYBFAZBYYQVJ5FBna5SLETLjzZwNIP9KjtNuN2uI5Oc4u53IbrCrInc
qjIF+U0zVZj7KHbWLqDRe0zOuK+WXn53Z3SC3tYu5RbBiITyxyR/+ddWaNWPFKL2
mu66iGzbiORgwgDBE2U8Ge9rNzgnWBOI//o7Vzrj29dbvHJR6covgTmCfLQ5qktf
P3ERcEAOwhJ/bMo0mkg7WHqR3TbThm10s1o2/FiAqq87Qczz6cMURZoNplteNtgb
x7GgRgsEbe05NeABOUI+Bv3l/p0ss5KNQpiTwxWqSPg+7TQIIvZ3DIoBBByX2vZC
SMrWj3gKH7PkTt2qXDu6c92Y/rfsEqqxHDOC7N0dODQiREP4evK7F8TVgta8yTEa
O1Y2z8dlmVeB5w8PIZq3qQ0utelGeE+tUAxFO+CKCra47epeY+MycWQSBwyPIqvr
FOrx7l3iNIBGv+EUp8dc0JFh5KprAnT7MgvwEExmnyKoYp8P0P6Mpk39W4/4mbZt
TWT/cSre93UU6DkAUegn3awCZ+MTjS7BM5v27T1Xqw7ASE4a7PxlaQ5XYhYHhWh2
3odxF9f0a8MOy3okZ9nK+CQgn6sBypyUWtg+MeJUy1jA/wP43vFIaV6Jljj5+wtx
mpj1YpPzMr+dG06dVKaoVx7oTf5+ynW6E13Aw9V07wSKByEdrL/3Qb4aITwkYJsD
Q0Bewq9kYPmJ+mJcSHC92Ux2f45fi8TbKmDQms32BzWDgRiMjo6ti06O4ESpi/r0
2nLfkdw8d9iLswXgzdb5h+XsjRbCtG9YTSDxKjDE2eXomDDf9rb7PZdwD5y6Mmh6
+SE3iRiT1bkUVxNxYzTxZfCzPDnFDZm1kwYoRB0UX6w+4mwjruC1Biz6WRDyjfwK
k1NrrCfT8JNSdvCZ5AezSJTw71IDcw7Vn+V1dOnFeNrZeJ+bgG9NWBAUZDPSV2Ou
19hRUkyj21bna4n1xxoZ0iv2h9Ivkhi48VZ5MSgmFDhzMdSGRiJE3Ye1pqU5EKWD
9hM2Rm9uEk49I+Q10pEZvs7t5keZzlTiKmrbBCTG7ojuI33gm3cV9EEPlFo9wAR5
g1DLMJYBiguVXf6eN4FZuWH65cww209KoLdIVOhohhznQ0nE2HBWRNInzA2p/MdH
hdtujWwqJ+PmNlR8XMeX7GMuGgCbja4bUjMdiv1p+/+sXbhW/fw35end1K+hKuFF
MwLZ4qXEwJOoMJgtR5O036rFHZSY592XQ1hZNmRvkndiwX90+VD8eybuS8zH0t0n
7gz0xE75w3gQbw6Enhjf7aXnQfO03rZC6dgX+NL2wR83PMHQk8Eizs8qjgy8JpXi
kNwnYFgIEebcM8dbFAMmNFVjCMAJxFGN71puUOvlT10PhhjIisWdLwrn1slDtKgi
vaM3+u9lnsgknWjA9Yl4LZwzOvSRLgpPKG0HPrUOA7hZNUwJpHMVRjWtTm0RgkzK
Av03R9DksDVmyrxoLePOmHno2N+r8Y+MRNQVk0EdajAVBMPbMhBqSSsYbsXfEQfb
N5J2JfTL+wgoz12Tqx7yNGhwaRZwGrdIqJekf+4eE8U3g6/vhxXupg8wz1kpQH7z
fEG1zoa5LMwKcgeDzEoryyRtyS0kf+VrMMr5biRp2HAHXQlFV0Vbj2t5tQfKPKvW
q83A7Mi3So0cMCMvnl+mSxDyASNJAIyESm+TS9bPPaSgwlBLjlPK/4XT1mhT/IR4
vM5BWr2nokgmnPqQ/xMQAIwPvjTWlI3iVgqdH/cyfwg/Hndu+l2WtVkmNoZrO0iQ
+aK06KeBvy6eB3yxRlbVWHNMG0KDCq0RsMEMMH6O9MzHJIcRnnHu6iXHp4aOfcvc
AuPql99QP7tDwxIVeS2aGNlb6qFRjGXbIiFNwb+yXnVVWh6IfRiJ9T2f9QN5bk1X
X8bME9uOrga6af40El6y0SltzN74MhtYROVGtysmUMjAIwGcLXDLCTYsDvyKZfEf
cMOmrpAyFVHX/MhX2s5YMWeW5e4h2O3KKvTMivFzCulzhGXGSh/xOusUZgPDBJrC
kL8oEwVA41fuKK19rNUso/OQL/RxKHieEH/QyML89QczT50uWE2e9McTWHpWYB7T
pFDW61r3Dw7G8/+xcr/YDuYZmL4t8s6br9ipSv//czwAf1uM/dgrgtEDdya9PhSI
8mPvSO6J+h2aXO3JgyVevP4vW4DEGuop0GzcAsLK6gT4Q9m6pNMMmbpWT9Jah05p
oLewgx0jfkUDPVCAhCaFk1SSXTdRalYu0VqA4ERDNpmUfltK5WO2IY7tomrahlm1
PFMkR4SCpJG4H4Eu3Kzwi+SvkBlAfh0EmgtpIEJzhn9meNaOB49MQZZ5AOTgCkXx
ovIeNQAXF3TawvT8J01KA++7kG5QE2MsmVORETqgukzRgOhXK0aU0ujWUuHobXZM
/fXGhzhIjnDfd0UbeZfl9iEseOnZLFovzxRrovWWJROSrHan4stC7V75bKBlS5gB
+fRNF0hg+LAGD7RvZS850cmBci9+ScLYPYF140b19vzQC/jBFw64B0usyL0uRH75
WbyJJqWSfA+zAt7C11+pCqoSKKCAcn4xmeC5Giryu1dcfhcS/5PJVVr1F9+IA4AB
R+WWDzeJJBUdy36B2wEChOndHPlcMPVIzcqHPvoij2u0f4iLe6IpBzGpobRP1r1J
UnuSguJEIxfnJIT+wd5dTasYPnWAdpQ9hrtk+chLOWASOhC4rWEmqZ0QU4kKBcXD
JjXB5zlD9IMp7UzNLPmnM0PbPZrDHDR01hurGrA+07//rJ/PnUlortrAmCb2/+ks
qJBOsfy3fZjLemdCRXgSoq4bL++TtpiDXbe8exk82NxZNkszNSJFQWIkrLVtCsbp
YA3Vl/OAwhhMqoBMr5wAaByZwj4Rv06OmrWqKKuWyK6v9e6MCHPjmtcgIriZGRMt
fQ51NZwA8HWEnsygo2mqruxAe/4SxtrC2K90YerehTJIesWOHqnj86zjITG4f18o
vy0JDYczs/14+fiLUcu42/pN5CweXb7VpIPenBrlLywvyF/GF1TGkPgTPPk5is3D
vJ6Mytt2FwU2jQ2EWFgVRQ5yK6FEAonqXD+YC+qJhERxXoUwc6e87WIaEYFSgBh0
WdsYIaVzyrNULnXCULepd9AMQ7O8LYi/5xd80WRLPB0JVGR8PDYX8v/nRjnDx5iN
unO7Hk1+yOxdnNjRvUJns52QRzRvmT0Tm5XofcMrSP7X5LMlboADA48cwr2LgllU
mRtuU6v2h/thHtyVvcd8W0w4Og2aZpzEaGHwTCAgpvsDtSjxLswRV7Ti7DilTk13
eji7t9fIEB6cvDuigOGs4ZzT7tR0ISwj8WmSVMf9aXtyfHUoCdyWafdL3xHMUoXK
N84RkSCPDIvTVMu5m1nzwHyy/gDK5X7Ic0i39KvWJYgQKoCstQadB4wX/uC7KU+1
iEzCpL3H1+LnJ7RiYtwy4tqE82TIx9H+b06DCAU0b7jNyfRjuU0wQKef+5h6Uxxm
Auvsbx2HlKrZS0YDC4gz3sg1oo0hBAEoEwI5740KveQD1/b09cnCBfaYe7oD6oKQ
KNMIYbnM8F9SY4PgE3MLbdkIhdQ7eDH7pUuWZlVAhV1QqRL0aXfT6Vqf1MieTSgD
jquTGxyUMUr1PBpNdAdGZSZZekr75Gk0/JlISffDbYEBPKIfeoUSjqcfTCR7DLFT
BGs3NQe60Gg02Bf6VULufrQ6qmdEx+DZRx+TtwHNlWOYjPDB6Ro1aNUVK72eezzh
xqE5qrrj452ppYMh1LUc16zA2pA+7r3cKtWW4Mo+InsdHYwIyFn4UKOe49bnii+r
Ym8NRRmsmZGRZFN2IpoE6916Aj4nauEbICs8oMP0swRI/o77/drnNUS+Wm8PxmwE
ZeCfxdH3ATCM+s2y/jVQbfxyYWngZEYKTeEkPn+yt5gWgsFVNRL8Up4jQu52tiDH
xYzEHTPIckIFfB8KK5NZejODnJZHKy4qpQpm/Cpw3PsWj+qBEVjOkeZP3H4Tv6Vk
qvml1QmExBTf7bK1/RPRrQoLYC43Om+u4paYyAUShs8mCb8pX10i6ExriM/WGm3N
avLz4spxy5mkO1+OEkNgoU9bsARBzvCF5qRR71f3r2qYW7FULLi0Rviu1kp2yS2T
BfQfSv8YaXShdYrTG2m69c87O2RSi/g+c2G3pwdHKemCPB9leIMigkkEUVl+JJKY
bxQfk8BS1pmCz34boWvx8FakU+hUOqzyGTIYq8nEfiik1Hh/Oo0S0w/WtvuLvc+b
1BWiqffTYZla6XhySRQBc8MKy3oR1DTWvJqVRhKFzjz1nAHFyJZ/b6KUBd5Qx1aB
IQ3U7/Yv27w/2CAoYGuE3XpsWDB+TEGLR2u9XoVoYj6gOaIsVQZjZSMVhjtg8hb7
2635wvU6P+oSkvJoelGsu9XcR/al0a25hzNIrjt+lTebmEe4qi+SPUfoVDCBniSB
bdrEuP5zcIbaZT0cxR3PVR3wMP9xcq/aApn6UndSHjjtuyeXyfwVjYhKksMISvMu
EZimX0gwR3EEjdAuLu36AXOKE/MVfD/ZRsA0Dy57UQgBNjjFINFoZ8DU9hA1mFtD
LqorTgddoLQjzy+hFY+mgR13WsvQd63/Jp3WVI5kBG6dH+z+TVe3ErS1sDFdsVUi
xh88i5YdpS/9w+9PlsFNNHMuzd60uTV5VucDePy3I2/aBy0KGHcCntEFyQPYofmP
8hUjQ/LSWDCCLWKdETIEL16Frxc2iWMtHCh79B66dgdWmPacuxU3yGprNDuie6GY
24YW5+x6mgYValOUhn4wrPLUWKejVueop7+y6TW03soeBWEzNuocG/2qEiyx6W1W
36XsUMkxkveHYl1610/ZM9u0jFxZo3GzNObBIcxNtB+v++Nunxahlgy7nxYMohmY
4MjRF+2PROBtj+9YbX1UXxPD+ju+T4u+6eciwHo+jq0cZwQ6JW+NO4a3wIhiIEZu
I/BVXI5KRn9Y6P9239eWnpDnM2PrwmYtLPFAca+U9jEufZV7YT/wpvAXjCV6TolV
K953h+7XB0RPlFVTs0IfpY/FHm1VSAUFblTP/Q6usM8B7+UMbVqIjNIEmj+IcCRx
2ZJ8Z3wuahL0PKrnUqzcnpPFCbFluq9Zr4Wvk+GyeDCAhGYRJpU9kMm5bs4Dq7LK
FXt3URbsjHk1C3P1b6VcHPkh4INbf0D5twp7EY7GUycQmw5Y+xkX9qfZ+MKSC04V
2UPUkyxTQ9b2Lvcgs5sXClDKaU+3sCgs4Svn3zSEe0ZzcVnIfeCK2/P/oS0TPBqe
BOCWpF83k4J9YIGuMoQQoGpCX/Nc3S3zd7xd/F1UROQKJSQzQKDc9Vwas+TeC3qY
7RjFvigUvnJRtlVCVvp54KiGt8KJKQ/rwwZUvgxYgA6dQ+fOTiH3YO2zoffi5O8P
/61/pJ3oAp+3iGtrXbh1NEM1rZ/+6KKxdb1txY+VPUw3+QPklQI4Z0jRumI9txNo
mh9KZV+lq4NZIQWL44mNG2O936hg656thgU6ldLhQRalEYhpnnLzaQyFP/W9t4AU
ygE6a/ZhKIMOTwx46327eTLB/AQEuPIxOgaUA+NL2mndwqVBo1ClJEAiKYiJ8oX1
OQaHrYrwk/pe9ce9HuFOBjGUP59yzDGUQ5oaoejhFD0lFeeBMkpegEdPtHYBBNyC
OBDU998sYJ0/ORPPyEs1TWcXg6y3VMZ2moWQZxvA8AwLshnPAXTEUNXLwkB+z9ww
tVMQdYAAOnnFQRN8AJ2rIa0MTwjLL1mvtg9BPsv4HceloXSl+iCpZe2jjF1SNPFE
kI1EiPyPDGZEpIr9jgehktcejZ7mXkDjOZWmt5kBmsIdCLmD+WitaCZEVBi6YMYV
4nl1L0FslW+IBBqg3hN8ItTTcs33jVzus9iUidXmJ4jaQCDyMYbHc7xZunCtZr0w
eVJQUT5+qHGRxhRjfmO8oV0kAQKeqRYRaVNANzd4y3lR2j1gl55DWlItdj+VSVqN
iTKmN8+QaxfyJV95jVPs/dEZ46AmeXQFaWoJHyOx8elVMRmQdKJ7z149O5weUNFs
zYezXU8cyaHTAex/JT+sdzYW2BscmgHc+y20v9hFQHODhEc65wwHN/0wDTk1NrOI
s5rfrcyhR7k7EPJnJ9x0x4PLiVglBoX07PWuUZsr1pEifUlD+Xi2+vWI6lbT+TcL
TSvft4TNXQxi+IZcejNg4/aswhpZZwAHDh6k6P3S6W25DhH3XHG5YjWVvgDk0P4m
syn81ncxa1J8gEDM8fY9ej4hL0LDmMS2Iq8FIb4dvW7hLus4LqVk2Bas2yOdfiPi
CG2up0dHrQkCrOM3ITFFSOfSlSSYXMC1Nj0noUZKlmush6ZxFWmUTgEUuSfS5kPl
7t707BZZ7onxtkGaR27J/wqwRZ8JL0naq/7d3BJLATHk4ovQiOjpK0sf0+NQxwF4
6gklNHqaXMPXjEFRh1+TLwqrajeqocwGfXHVZJnIf6emMNpaqMjN9W6Dg+di2cqZ
YfBYnTrwDiHifTxSwiHsSPuFMOM51Su4B74uWLfkwdkK6l8JoOOELs2Wqa7lbG7W
lsKxF5Zin/XuN/8/3pWWusTuKil9lNPBhK3t/f6LOK4FdJ1rh7obUwT1mXiiVOPa
B7s3znLPd6Z5nVo6OHnxHl0lXiCKKP5b3ZZRNfchofYtYv0sremX8i1N46sZ+zeL
hzS1Rt/YHABe5E8QyJIPvvgh7/3bRMNyX7cVUPoXG1NH5dlYt5y0me1iL285xBk5
aMVtC92iNyyzZAOWlSzymOoV4M1QggP3RMyGQszeUudkQy2Zaf9SBL2FBMpr7hAv
ArK6QGXkhwwFIP3VV/GW9Zmj0GDk8zljVYeL5RyEAdC4QaAIhMi/wiwT/Rx4WZBm
OeTsadqdpBQ21QGrD2ezQfpQHFvAzg2n13RYsNIqKEuWc1pE6hf074Lsjn2T8WTQ
RkJP/LASf500OyktzW+NJpUgqXoDAryJJEIgAqr75JSbBDsJYj++Tiur+Vl0r2Rj
2UTkk9qK/JBsaKQguM+ZQxieBM2brjAgfX7xzjkNAVNEfWzLqXqLyK6sxmlKWsWk
fr77EtTZk1bnxVi4IvHkeUfVIYkUXFHrheXk1k75Gz1x4aEQyOmmEKR5KQNKYQUk
B09GUj3ZjDhDah9NiZtMjABQ/AR8DnGYviFq+f613gQpFzuWdJj4K4O59l9JgRzz
QVIdokUDucs2QxzEd1F0qaqIWBpEMtNdJyJ7SrkJXag0InLOmzqm4EX2ljpRK2S9
iKSwp1DcBtYVbh5eyZ1i22xROaKbNlRjbcQXRTH3vlYSmZir7EKf4VdO+aovAvme
enmcH3C9f49R9AOe/ikzQdyxC3ZNHNP5pV1FIgVM0KCz5sqJeXjrYaeYiWHHm2QO
42lKtUdPCA0sztwxNKPv8M6ZEzp7Dj2S4o2EZoRV0jPaZUKnCxBwWMY7A9r3ilKI
hfdM8dAjVsQTxTi/BEipjtv06h1HwA1WkjkqktEeBSIf5aGuTR1Zj/BkMMX7qzYD
l6TqxiFJfw881xPq7i+hjg6p9FVH2XjEXZzYvwqtojgLyqUgmRsiEm/HXbNp/rcb
u04nvhB9I9541CPyX0RoWaapXblU7bnS3p4GibWz9qhV0Sn2yIeZ1+YJEEOhfDxN
Uy6Qxh9ZtHryiho78f8uD5yCakPxJrpxgzcauROTEmAkSipE6CFtnfuXFgGQRgNm
PvUxleVB+NUF+2VOFAV6FiKLmio/9C3obN+XoHoWKmUeVtHP7jnpDMmycbfimyHf
/VsnTB5UYwhqU8kMttqPLkWutcKw82wdjsSUAJweyDdanShiiEtbfqtCWejQtwjH
ByW3OrL/Pqwdt0/V7+FHIp5/x0cn3Rz+5kM+QevxKOOD8erei3BvUJDOPFpRlf64
hW5TyjZkJ0ywOYqTFzN3ajzDWp3RsT2biS+/Hv1NAmk2DQa28EnOB4ZvHWqzOlke
LVhlOfFnP98Wr02d6XvlWlVQmAXwNB0kQYaG+j0LXrRG4zF1ojVBnR9focekZYDv
RbHnS/gh/pJtp6EWinIWq9VATvpiKhCIS+HI9MLBkN5FH/lO3V6YM9iMyAFtgR7h
UFjylt3m0YepjK7+Q5RBXWsljjASvnRygsER3ZRzxuW21NXg6EvSdnL4DVq8DPZ7
VY/FTtIjgiN6RXw43h5oxj2+pTDgn1WZOTXUZtZJ+uORDutoJlnS8NJGb+VYEMr5
s1TUfZahHcDFV0Z2b+iyCra8MrM2HVHma8ZoCI9eiC6+RDzBkzKLFfSipDMw3HuJ
HtWab4Czgi8KM7NN5nXB0Yc9JnDeV9TcC/mSqQoTyVdc23UQENiU0vtH9dnrTKBb
FnaI/IYJ1TpicfFNsvt6txMSdZMB6+BHMLO1/HTJUwsDV2xTS6R4sMzc7jtFPLbL
RzWsrqJswF7auyJvdQIpO5V4sVqJ9TXrmSzdi7MonY12fGgy0unXo/GbI8AiXNiI
c8p+kocPwU8dTO7Jd7EjACAfHpAG/Ag+Iv51pXi2ZjvJo3n71XXYlfc9tC/9EMd2
m6XDqqXcymZ1jECW448mNZlHJKNIwS9KJcls+gE95oNym+cdgukdXgwYIdFEB/Kh
BQE2Evz/uoR8MmKMXIDv99Vfe+B2WPmbH8wv4qWbWm3LBfT0RYtF9HsE++4iexIl
NMFKoHSpHW+ojfrNUOOaYWnxd1zRojq831JXi8O2An0uObKM1d8C7iQCgP3IzR0M
QFVNgzi7/o2a+88B30ZL8wvQgKx/x9kJM8a9dmXyZOBCk5scFspTVjV6I2PNIvxU
mfHv4Jj4OSAnsjnR+Q0D1A/zXW+R3ws7tsx30fduKTjhAsrG7aj44YdOKfGCTDFH
SgHPurIBjLu854nlV89cWm24t2kjCNXpsDxuvP1diFVRKH+571ob5SN0nk7vp7Uw
PoxJiuyJhp+Wy+e9mhYebcD58EfeiubXQetW1uU9Yr1P9ZkIpC5CmoAKJaZ1BqKT
b0bT32bIW0pVbAjYK39GzulDo6KO7JtxBnfoRm0nwogNHAcr/tkSi23SdcbN6mTy
JIyH55vFur9AZBMNG3pjzI386hiWYhHGb5pc4izOrsZtPS0I7uVKhWGlI3G01UrW
Puyx/aNvkGTCQ56bnDrHcdGIQ4AGULlua8GWPZfD29TC06ny81WdDJNGX0G33ARj
Q6fu83ISbIe9Vsel4YHb93JoplzD3jmr3OyaiZCc6HSfnZaibuu+OlFimrVFw8nY
XwRpk1Ckd4AjDWTtRsDDRWT1zZ5ih0UhPzdi4HDyUXpA3DEbvHQRr+cUSbAaQHcV
IeZumkvygv2RxktmbL5YTfssLKWxiHwtaAJH6Ps6mBs/mWBRmjBTau0TIEv7kRz5
LGAp86NZS8ulbiat0s5JAb1pi/f/CTf9uFLf/Y5epAtG0oC6tqdgkXcUwgzhTTit
c9YXnClJ12j6nPjPZ0mjGlUPM2fmFCtOyAE008GIHlojF5NmtFNpx1PQEarkHpnE
Ha+C9HXJLABxBDtQSH1au6MzUQ16eLjmgYqAJc8+W/SMbnUNvjJucC1iT42YavV/
XIm72lyzXR+2/fJRYc5yMVVZV/Koybn2K++8EN9LVwiXUIRgDo8rmB6mz/6fRjd8
WbMzbb0Dw3IlQxCJmiiPf2/a2nW/tm2w1DQJIjAK7mErg9jeH5+ebasYE+pR6cpn
91LrnEUO+iFXmQ89C+bhRFJthOfKldUN9WgIhUaLu8NBoB+TRH75YpKYmkj2qQAX
zFbPMmdpqoNfjFGRw36XhVxXvwwpxyfEl5LG+QZsJyjgIV/c0sfQlIvC0iLtB9VU
OcLIeb1F08hD3+7uyPJCD4enRSWtgFrb0PmNhjTYcMnIZH8faap/j5c1dwe7jjca
pARcRi9HHs6Cbo5dxzZtBBHdFFDN8oK578vBCAx3A374pGhO9RlXpvlPVsNpVP6w
3TehLuC1pZHhlzWgYJIib5lxHJ5F6ysGR+BlZp2V/UepXyE4uycBVtaNfcb151MP
o7xbrdIfhzGset+dE5wwMN+edtIxhxuoYWeW4Og8iFqDvbbMmTy/dy2hQWBGSyrH
BTJAPtjS+owWc6VKuWVgjKaSqIPf5FhLi6bFIV+z5FM+i9ewDP/7h8Ll1U3LNBnK
DEfEaaTsIq3WUpkDhfXc06wINvOxAj8LKIlTji4YTvvztI7CEIIaeh1gLFDL+US7
CZF3Y/huBEeaH11FqYwl9jLGgr+BZRF4uElDXOIo7PRcMrObhsGGdWqhQ0wYYRnO
LLjM8Vml1TvOTd63mBSPz+BNEZZ6jMoAZqgbVNksC9UncQGJX2f7R0QwT+uT4O82
cBfU+hpunop3/15QHLg8v/6Wi5K0jQU5o70uF9VBfjBcu/KQaAnSePZ5h4ev2cSS
ikHnNjD7Nz22KtDE64djWaQLlsEc9c20KzRa1AB0qXo40NcDWiKr9UzOi7lhtbrM
g6sdPpCp1woks9kW7SR0QftmTBFvb91ME9UwdsHyLzCTNsBpdw0G0MAYtH2X/PWX
yI6eiijZBgiTkQEMCicQ2+xVcoxNChBfQLywOfEQDUl6pHweRWYdVMuShrTpYgY0
V6Yi7ldZn0EglDaYD5L9hGsKJsLht9yYmSXsuktYYh2WXN88R/1wxzShtwsGycOb
9S3Z90yja202FIgtf3RQjgpEMV77zYHsfGsgykzWMgk8BP0SD4bFzw7zE7dXjb9M
52CJhb+3Bn5mgPWLTkpZH43EIId6Ul8KeIWrKBF5+X0+/MsFL4yyNGBtCnu23EAa
dl8o7dNiLu+nVPURfRZwvaAKfNB61+i1MaoTCPswKLLlk13SwfxET353tP1PMhPs
5rYCi2Kb1r7ZCF0cH9lXlf3TD24GHzE8qmCDNGf9sWC6iztD3g3+7+rZZB+Bzwab
nmrJ1BjQO2Fd9urNf8dS9nfpxP/xFhrJrMOJZ29HXUyz/njd+hdmRzfcOIaiOmyn
E2QeAupZNlDy1umJbLrBfiij304lFwCa59gvT/AXdDclSy3ZCDH3szsH/LrijD1m
163yBHPMkDNwaxISVjP+IS7The9HuoSC218jQypq+B4xjfzJIMimJHYAYPJOQL/r
vMYMai7E+PA6k+zWJoI7MEl56Ys1rFCmmac9glO24LFcpXfbNUkPuzUR7sp35zAV
ein3V9eVOU1l5zSAFbeH/Nbod4WHET3PpaAJ+a0/DwGmVZhRahenOptCH+v8nWL4
8fqjOk7mx/TtjkHEMKqgNIgG55F4V2UHSXrBIyAIOoFbrt/7GfLhqS4EqxW6yRRs
2sZO5DHJb76titLY09C5IpD/qfV7g20PLmnstH9nA9X+6zYv8wZkJd9g3yffUn1T
FeDndPkpCNvenntOiHXwqwZ/uaaP6IPxerPmCBEtXL/M91OpCjTIRXYAffk4Uv6M
Xf1vP3eqFLAX3GBUHUO0ohlxI/ds0JqFRl4a7MaJK8Tyog9BENViLQv930tAh312
79//94GYu4ffWMWtJkjkhaP+rGdHJ5xT6AMP9RvnwznDNXp3YIQTZPTAosCp4DdW
xwcHY/eapvdj9Ot7vrvW+PXc/0Mg7wjrZDTk3r5wlMv+GFA1a3kygWIVRj9Jl9q6
c1Of8LQM4DIfMWkxigVr5M753u+rqR2kYvd74R3L2X6d59PHIV+KmaA5zA3vvO7u
2nEFsVW3O05HfdKPnxBdumr8LJkrEviqONYwtLMM92jlOxnYsHd18ggzjTJDLgaM
tJu1jhRFYQqPhqspaamm8JmouGP7rFaCylydjOeJCak3D61OFc+qObszl7cTwnTw
N0/gAn1LxOj4QcZ1aAw5EtLEdLMrtk4GaDpxVMt/ODtID7QcR3u+MzvZORgAcoro
lBHFh1LM0gy9bOhnS2huBGaoBK2Pmiu0IyXE6Ao0N6Lj3z0h6GGklXdA8n6ejBTg
YOYqZI82SWPoJEf5VEfazYctVg4KhJTc7D8M/XImmtiutGeEODMFphzWaA6iY6VW
9zhCewTIPdLUVv0lUv9+LRSfGNpiu9pRWINM8EYplEjZCv3c4lOGgpuqp6sNIO4A
LPmmlrjqA7mjxrpH2kE2ELZc3upvkQLQuURusbtVQNm/nPkzr5TRlZqfnYWaamC7
SsK/zhSyzOyeL0LM0LpjmQ50fTT8WHfKOMSHOr7aWMIs1/Hkw4VYAXonIEVV5lO6
4nweC8gb7/z6lvgWr60s1Rxkm/3v4/5PdbK0DV3uvBncZh/03dKyKZeNhnLbcNwC
HvqXRVAReSD9Cvtom2yyap6FmDyG6VI6eBsFz3W7OEkBL2XWfA6MB6ITvZ+I0sEa
153Ue24oTKxZMdtKl29OFsjWc6N3FkZTE1Lrf+kxQcHhGplrfWlNEmmNkL94+epu
xSaeN78EXB0F6jK4v6GkuJlUdIsF3pIhOmbM07yrWGqrwfi695rILAkcMrMu9gOy
2GEqIF+rw/NuTf0OrCPzl/d6JdQbrGT4lz0yqRqr4RvDFvROkwCyytHkc4PQP229
9Dgha4uTAyDPqMUPF09s7avJNI3ZaysESOp4Y3PJKoYl4o6JmhABAlaXePsYzXur
YHEWPBpHseqT6wdCDbIyiklsbf6BZCveB1DbG3u/CaHzzi6PnVfRgQina1uUEDY8
7wB6yT+dWGeSIfmIZgeCkvk+kHtnCRhmxZljQgnC7RQdo3bow7xp+2Q2BajZsqK+
vpK/9MX77zsz7k53lcakdraVLH/QDblHsn7gOo6cVuxVnXxMJ770A/bTTQSky+3i
qW8J/lUXTBbFHJETK2aiuraAON26NvRz6yC5gwm8wTcO6RT7V36oHCr0vwMN3IvU
HNsx160Nypn2I3mvVDBRmv3pwv1WSUFpVGQZ9N470qv7kVv7dFaLyRZhYkbdemVY
+ZcUwsvQ6wIb+4D45z0SAAgNiCch9Miew3VS/y7isEoO4/w6QnNuRvvyb382A7qR
8W7pZSwKdADH7nreB/3mLV4yLMH2i7/YkfptQbjX86u7ZkAcmks8vdqoIuzKYmG3
DqbMlf0uoTCpaDgybEaRu2AYwgDK8fXQbFRplMhVTwnRA/dBlVCw/NynxyPiBKQ3
uox2l7y6jkEBx+82KwTvBXB8+Ci6PieuxN0iRxeYMsJ3Vd75/SHbnT9j8SkZbKqn
vSaW6iWBpLU6SDkq7WqolK6VkOY5nTGmECDNPDRxjZWVQhXHhe+rVeeNJomfoHwH
5yq1ltCcmZ9bbJOlUoyqIRDb/JyHmGGGfGEevp542o8PsEXIkcZq2lSWiDX7L2bE
VJtar0Xhn1mP2o2FNPzYmuLcvETEA5JHxg9d8mTubIDkDrg0tJsPASkXpTDyF8lD
QaSWjpopIls/rKS+3qSlG1ge0r5zlgg1hovgEb0SoQm0+O0PuuPwIsbMewXvlZyH
k/vivwK17UiUHsu4tJgB+D1F0pgwyB0I5sJhoJh83994Sd5AnREfIbYIuujR2zbc
rWp9mLQEcdo8xKOCXXbLqD+ZoVWOlmKCPvfC8rnIUPecAyFYGdCux0TTMb8QN1QZ
enIEGQ8alU2/i6Xf6YHwMDM0q4zb+PjqLhqQ6CeEr2w6VLmraSvtZ5N/pGgeeZWT
k1sWfHacBGotr/MTd6N8xhaWWoRzbbDslsXaAZcZJzJ+cs2Q2YBi7p+7e+LmY9D+
lffRQsS0PuoWPCzlKoOTdN6UuEoXP3cI5hIzJdPrApfmRq5VnWkhkYXk7JQwI8EE
peGXGFIDzEzcs8IPsnap3zPD3oHdlJ7fVlMXiWwr3FPPfYY91dCFG3Rznrc85Zqj
GkE3QDcBy7qxFQO7uCxKd1YY9SvVYnH2bgvDLPYJWVPDrrVk9sO9ZZzCkPHuuc2J
AWSTYXvojrhL7AUA0MqAzn1sCAaumky6w+VvDZfIwnpAiT0Xke92W5RUTbv//qCN
Wve35PEsq43jbi1nV5V0cOvyD5eKWKqY4tbUBGQd5NBUIjHb20788Go1M3yyEl+W
9T+rjxSv+Db67mt+3fs/GolKDCuA1KxFY2SWD2JR/nTltnVxb9w8y9Amj/Wui+5z
k2sCOfR45Jnyci+T1OffnSgFt23R+hhf+OyzGaO+G+8J+lF2Mqqhy5hy+c3o3Pum
Vh3KWvoeUNlXg4pxIKHPHeNAIhXTRfzIjW5d7eug5/Ak/4YqA0R9II+ZsWhFeCSE
F9Nxio5JBr5D0dClKBgoYvoMo4jaQtVr2QlCLbyYH2vS2tUNJ0Imz5TEHs/1UL4k
zD4RzzUKgrYWXQLK6gNDOSLpSe3Ylt2EA+6ecL5b7KsRG2avBYKoTS+hMALXphCG
YWCy1DXkWItYlQLh5kyrXtmI9ktphtN4jjgg131nI0NADr2UdgPEBgNWgOuLt8yQ
P1HBhDXtDrP3tiBbgGsI0GE5PlGP7evF2Ab529GwnEtE+pqAs/Ou8BNvDtO9nBSg
wMmeRPRQ3ahSeW5vgc0djoML6TOpYJdmOKqrtHZL5IYtYyeJ6USwa3orzb1oU5/1
ocHLtbaQr7dBx8DASIFre1stlqtV90IwOKc7fHFQr5DhRGrnF91+w5nThncLDvMS
Pn3BMBU9FKM+1wEgNJ1zU4RkqIMiHnrzdpV7in78n38Khcu9/Oc4sXf9+chKF3kp
rFd2VjV7AygB/8IFfPVjzLkkKleEd4CT7PeiRusHoosbqOsrDE/wCRcX4SMm1TAk
C6BHgnfUT9rBs72LLvCYOCYl8a0ldoJdfMbEigKj2IGAWRxP+4utO0W2yJP9jkP8
z84+Ux7oO8wN2nLj2x7xkgNYo0LeP7nHYzj0JgEcHawBVRf+mcrGUiHVeNQAMWml
xF6EzrUT0dMNj4mFjUNppxdcz1IG3Uyc14o9NTkV0Pm8G1AftOIcCeBln+1FMpDn
YukFz4my+SauHHgk3m5AymDrOTIEAaV5qgbiUvHeXwJlioV1hejSS8SNASWZ4+Us
WztWSf4PvNbopTPqx7cvDpYyupHm6peI5Y9HlMqM/NkiCeOM6gZv7yQlbnEl6QWh
tqx/8+I0LGfRHQseEi2EeDlUQ2FtVF+5cRpUz5v8AZnkkX+kxPCvj0cGZ7TbDNmj
IPFHFTbs3AB4q2eJc0adDnkJAo6FdmdEx2Hiw6XKGgLOSQLNRBLwFxAiQu9/fOxd
dWq7Xx8406QDLuQONkh7lK11Oebvo8eZynL0JGJnA7S2m7zI48ixYJLXGcZcWjMW
RZhBT+zwrRc7NgXp4VjTahD8KJ2mV6z77Yhl4Q0GY+AjXAwBY85NYUzOEsuocz7H
997eeyKajWrlU0ZAPJsvd4SBtdl0HEL+b/7HxrtXTY2AygPdhUD6w0mV0TGAyGMM
ynFZqaGTNkDUKvtWq0bAjnLFWxHmjyVK8a5bZcyHZkhvJwpKt4mwlJx9OKG7+Tnu
9e5Piet0a8OixruBJhXDMQosByZHYiceTENSHDWeEBvjfL+jtrnS9QlcDhsYuRdx
/c4+mgBjTN7L6swvsty7NH3yW1FOOBOMhcdQGkHqRsIV8jBvjqNWi1+aNqJHqQ+Z
OLiwBbnkInrkmuMHTSDUvJ/9JAWu0Aca0/BrG8aw9utzZnDL7KCgoajHZ12gefQ9
h6pCE81R9sPqSaLNAUVUyogpEf6ydQvBU/6dAQJlZ1RtOWQfwGQo4KDDo2SVTRxt
4B8/W6KpDImlw8ikuVtzsWuiWyyekSV6gO8nfyRaC5kRDdIY7tzcbQOq2W1F+3ok
HmhSFYL3YqUWmCdxgy3UFijzziwzdaDMGZBSvYAtU089hNtbVXR16Xqu0cb2u+7V
EnxX3qKSU7YWbD+MfieXjHro8WqI+YL/X8z1jyEryjzBTKHwdDPhFX0hrjYyjvVp
Wmpuo4nc5JMf/u2MqS+LZUs/D4zxtc/jtFlam/5QGyHAupNBZ7DohCI5ezlG9C9a
mbmCF1c3q1XM/91Rvmim+q1MjaCR+dDuCD5TjETwj09HnQg1FVoXJ2FeV8tPkBYj
ZtzdcwkoLQIDqkddqgKQA0Bc2ECcdVg6F9iDLd1X6x7rSQ3HS4eGPMkwKBFk0U7u
beBbGh/7HS9Q34fmuAGPdaAOf9MvY69zBWZMtzT2M5a5ZGi2pHLgOE5asZEf/NN9
EXbMSiNV20F5xaDAoRAKJ6sAQ2+csF29px6ko0AsWGTwbof6Uq2gDCcrC+CxAUbJ
nHq4lj5+WrieWqTM1bePXlSKOWb9EQIZ1NFVOc1hC73JhnXKYsIwyxMZXhiO/CmL
hAm1jFhhajf4506pay38oJpNa/F/U2Dz0J0f1dQ99Vn7xJ7HlKwUVrVbFebJyuoX
by15hNS+CQP9CtjjoPae4RCNgIXiRJc7KOphaJqBFeyU6ToDw3STXAM5NATB38NS
x6TdM5V6Wpywbim8Vj02hNLSdwVYu3jHx2i5TaWrKv/uKISZUTsloN1J9muSpqdO
Ih5c11OOaw1tyLGYb+HBdOduSsshZPNzo7L7V9WbfJUzJMMpmnU0+BeE4zc30/m5
UNZiIJ14z41IKGYf4Ws2hGlZaZSuwAaJPkOCZyC28rbOStPKVTx31GO8MgzucJrf
LNoga75FW1A5hSGKgi7CHKGxUO0EYTx9XEC1vfQfzMKHkbcc7RgPGVV7DTW4p0XD
XR2TP6fj7O12ngoUFSSml2asHxGhIqy2xWXayI8wtk1xRSyEzPtQ1ISCEyXuMchX
lJECOuwpAxOFhwKyrK9iZx6iftUT4eQOoW3fMnxi/hoqR2rQKsLnt3qWHmoR4UT2
E4X8JXUdLd6kopH4YUUO8QKHjN882vuWYkWJu4+8s6hCaaikpOD477q7YhCiW7dD
LFaWSBfRS1XRElmMpf2sQscd8JG24N/dRhwKuzYU4MGSja1Aqaby1mWB2NmY/GUE
jzJA4GIL2z5nmdgu/CM+CVagkEbvFElbNKK40SA89Z95Zi2TD/+ZLx/mcSNlkB4e
CmHw8ekQ/BNIQSbjcGptvGiCZ9w8Wpe6HwAYNaaF/2dq7GMP/QPM+M9MC89vGBSC
Gd43EK3TdHZJwQ+oUYvV5YhRxTMaRAlnbyc3bgmwjj9VK0OnZ+OSVfDWw+5LAjsp
Cw+asvnaVSDs5n1t0jU+6T/jGfZcZba396Y6hiMt3p7LJZQPD8yVuNVtlpB8bVSY
Ie1gMxm3kmrVknhRnBMlJ9KWOGmS7Ex57Iw5q5GNdviXr8b2AvGI9SX4sZbF/O0D
PB0OAaHdeZ/NU3DmTin+BzHdHu9+qjqnOVrijnEK9aIO/CIIzHGnLnkXmqZN2rpD
TP3JGHw7ZeilcHebaDZ6qzwcS6aFwbXSIqiqSuIeWHg4IyptYe0DE8ry17MnZ4hx
NCN7X5ah2xQJOKbQar36NKPfNtCgqdjKTlcZYfKVGvR5DABTbyaIbqx5cQFxCz8p
6f89bvUc/NkLCYWERgUnKvSKk18S0WjlH5ePg8VroFdHMLU4EbI95rYQoDeHiw0D
THYrTGjnatjUtlRWXChc1MieMY5TddEAD5/srRlm2Pks//OPPz7GyOUEiZlNhRCg
teRM1OVbjSdfGxg89eSJf6OHVd1n3m+7hJ3sGxvoUQuBndxdWAFJ3e6kUdtC7C23
NQ2dHUgOMu38TORngLmBSep9P3okh8cL0TbWeb2MWuidPF1UDffi0QXklyPgjLBO
uAoDgpkd/GJ5hAD9EB86WK4A6L5ZUGjMfxJHYqCkaBAHk2w5IeRuZOoZplXCV45y
D96npwNG95SCRDfKrioiScauOY/0md32DN0h3UPhtVRbr6sVoQlrEixSVxI33LiC
a9jLG0mNK8pkFdhnZ6ZK9xozzO9B/3mjQdrz2i4Rc/doSBfqChZnixNuO2LveKGK
QrUawRzlWtuBvJ1CIcbdPuNXYLx0OQOvSrv0BzJjHNMxuTt92PHqCEKp9Rbbpzcx
r5UHwDNgTuXNFsgVYdnp0eH7SAxzItHFBCJzyBjtX4fvjXQ7V/eQt8F+Uwk2yjeC
F/XZt6KOC66LwUkByLJqBIWCxs/bspTP3IfQCJPhtwcLrVhuLik8L0yO4WUTeA+a
5y5Om7fRHc+utsw8Kj7on67URD1QUspU9w6eqvvcMOL0l0cW3Y3tfFzeuAnPC1bc
LYlcTSr3lnQXGXFd3MPK3ROYdsMAzUTQVL5wDZzrxgRbODFgvbFaZG8IQn06Xrwj
LCPkfuklA+8eFJPhsB+wmq/tpBZVhxcDXwp1n7NO6CIJ6iePuFlvRaddngJBm4+8
E9yAgkM3guFboGSj+chpRIAJ4LDnC0w2BeIZD019udy0pCOLcgZUZiyXLLFXWaeo
V1DQ8SKljSCIjWhrUqWz0aNGG5hRtdvvYUXu42h5UKfn2BEW1hNg7ZUu/3myAq41
JLmptZZ0z/eta1Z1jjVxoXXUc7SpfeLDACDkwMDKeejYD9N3KbLGbv1JjAPzcHrb
7/u3WDxmLUQqWkwk+7ffecwpPne0L0X7KUQRV5RGLRd0ooZsw4iFCeBSZlcf0Q39
zG8fcQX8WnF1jkln5eUS0PnIgf5RDhTG7IMHz6S+oRcAeHE9MkYsXv+AD5opJR3t
w8oQaz5CabxMsLwN3ndFyBLIycMjAd6n4my2t6e6jUMOp3oG2Tqq/9Ync6+lRnqy
j4tjlo1IaX3LpnwPXKlEiOrjN4ep+FwVOXhaQc4zCzpQd10oW5EyXsLtvvpz1I4T
JiOuodaOvP3E/X9xSn0q3GruErQ/cO13bq++Bd0Ye/tnb6Pnc/pYFFmeXoqSgIPM
Xrec03trTrvT2AVnwYNeqmwsUCaUU7d+uf1IMWlaEnYD5hmCpmzhhsfeL+CXetQf
mTMvbBwjfjiyTXRYISxw/xCb8F+gRm8+7IqFbKSzXCdeT+uiqbWOcbv8gKp12jI/
pqKlAgmAP0EMFU5pOGzAxrk+vj+h/6nifBqKxYNVNEt0JDB7H0NOb5aNzYfyXkBB
LJ5XugmEjaDjdEnwqG/38qkDbgEMPeINcbzQeXtgS6MNuuuiIoPrMJFZ27hJlqJy
k9HC/nzn1O4Mj8py30SB/wK5FYGeTsujXotniw9up8ZYFNmghN+Su3DY83+ea970
siu+KPS4PJExcGMWAPqX7tPQHIWtUOLg7QthJYu1MnB5QSra0j5otbvX8FBpPSD5
9R2ihKm7dmOWG5OP9MkhNRaUWA2m4St+3HAi9iXT2JiqMHOVgKr5vCgeHEqgKl5R
DwB50tRlvnUlGsh0vh61YokCC4LhN6MnlIgT01LIpCbOfrvu62mDRDd21GDvJpGa
ep/suaqELAKT6YCnjn47xyOpGL3ld2IcqJlb3/R9KfPaCuDdBWiFkscVgmbIgF6B
yumXOxDeWHhZ+TyAdggrDoO6d/erFt/aBHKXDjy01NME8y4DDInjpmJpdp9BDayw
Bp+rXP6vKnU4QibwZqlW4ZO+8exZG6riLKuhB1t0KL4+agfpDw38tyICJFqnAMQX
9HDy/MIVI1sS8pZTioBbogPMgp0tnCEhUvTH2To3/GqxBuqond/NcCysVqMeWKFT
d1wgQURXwqaF5SeZjllWjz8MyLdhJQZ+4guNjeg6+t43jiMfHb3exzVtp8lGKxIg
C+OuUDUqC1lE5ia22TZoMdSx9+iaNYdikLTAcD2kuGAoZhEloXNAnYpdUFEm2tfB
ZZZZjLFINzoO+tHyf2j5RYYrgFAzcPZRdjQOWYTICqdtTo0SO7XbEfinkcgg1Rat
p5+e93JCp0++rT8pkX985OtTc3tyAazGaK6pBGfPkBhESvg19tJEDrhVch3/pFMQ
o6XFnEa4KoX3G5ODmVz+Mctr+OOeq0rLNDFv/nJNr1DJMspQrKgajuvTfm55pKr+
fmmOY57vaI3/koMb/8MDmnM3m7rQLwciHbg7qvXqnajhCiI22cKJgft+a2UmdiqO
qN8b42Xv+E9m3jZS+Slm0DLq05JxptQy7J1VqkmYB7f+xuBwVNJoz7/ncnOVNxNH
Y7WJSEUWUOjzoYRBmw/K2LHBuTwUAoZR2DjnMrmYhwsOZyKh7USp/lJEtiCZTcKf
xJvQxC1Tyh/i6WlGxF7PjU7sQyGqgx36aQi87njmFOzooRYPlXVIBYjbQjskGj3B
/gQbZae2H2yAKjfPDM91tWoGa7DMGaYZcgaIngnsvhmfqtthnPddXvUWTvDKcqEV
93MLqBM++7mA6PvwwFFpGpCKkOre/JQN/1YKKfVO4I31JT9bI8HDoMKaG4L5ByLr
rTVohhUox73/C+8Op6MiViRFbutGz0GGzTCreOzpTDucIxMCBxqeNmSeczDDs/SZ
I4wIGbwpoO9PmzHM/2gK8dcW8/Spv38s6PmzoGS0+qysemL8AIjZaaezyO//6Gok
aunzXfuO4T33mduE2Ougc6b2SE68oSxE9ZlzSYp7LupIZNpdRBfvk0cnBni+ZyoG
grCY6Rt927d7J6NasKlz9DPyRN+hTcFzZF2rGti0wNOJ1GtbZCVapw9/e4E/IMLZ
K8Ur/Qgm+UZiPCBaD60mf3TC98IFKtAF1F0oau0z3kKrj3wvfL9uZr6cKPLExhjJ
oVKNEDqK96vU8oS/6DRUVX06LC7qOAclQMscj9MmVNJ8cduZCDb9Mp/A98RjB9mn
UY58JbKml9Q2oIOAj7sG8W65gZoQ602k3cnvbtafyJM0iAfJNg1LWGCrbY+MYVYh
ypjrhGpHAmG32+/+i6azffqfa5VpmmIdLesyfickFbAcwshns6bBDA8nZHvJyIOf
uy/dSctd77NgvdrrjqTgzwWQcKzQJXJ7XG2wp8uRwEYmBW2BG3tl55YbjVFl3xMr
aP+njsnobqkYtOR5XWFFwWbhXYGlHn1zJvfsTKoSbfxJinfgjuhUFyYxNDut/YR+
EW7El0y5wxWnwAUmHFU2vTnOJNjoZY4YnzM+dxNdY6iukRharFaXgRr2O/ncYmci
uqxLN8YPh4iuYHJc7vYd8ufrV183iaGqMqQRh6a0b8YotmGuJ0ntGptyPh0dLCpL
WAOFkXCBhKUUi61hKDH5YJyyIaVZT6z+9ePciCEIBm92Rl0uccEKK25ynKwIhNrL
+XoW/Lvur0wRJ+QEDp694DbMaCEHo4RvznY5jqc3Qt9SxE1eudmnpTs5ho80TuMC
H2CUzhDGF5RCWcEf5LjtoEKB7p7VGt5RRrMTWrs1YuuQ8Hl7GDVF90bueAU7NwYZ
RlJJzXG6poM4+KiG6fLNw25rz9GnLacr9KS2x0O2wrzZLMm+LcbpyzMYugqknkHV
ShlDIXARl22pS7Iaj0PD3OmpQgHBbWK5V2QwotipLw6JIAaSc7Lm4ooxfyoRn/WN
BREeSSWEDFJs31L64aNIHJK/b4C8JG1O4wVaP95CEDx84IQkm9xiR22fduo0KmCs
ZMi0IdLso8WUU9/8xM6S59TsXtR750g0r+fRRz5Jy+GWq12o5uzOQvZTv2BttiFd
gMzCcsoaVIkHnMZjKnJ2Rj9sslz70PuDTtFVholJNS5qk9VM7dgPcQBkJ/c9fUgu
k8DK09rABNz2IXoNy/x3WIhGv35fPSZSiGrTTfWb34RsPoS6zhiPKZkyb5wRUafF
OA+WCUrnmNwEVY6pDcoX4EY98KzbqGnOPrHqcEw8nq+vDKe93mee8s8HaTdprisI
R0qg6iXPBWBE5LQp3wb6Hw1lW3IB+/El9tD9c4t11ncmvgX5Flpa6PyeMlup6hW3
q3arxxTNUJBoEqh22GRijbYlYPP27YC6rE3l88PWVr+HaPz+maD9Ehe5goijVs+D
WK7KTvaLUQWSWgq36qReSY5wt+c61VppcSradmwxQ+jC+KdVsb61OYDyMJT1G1fU
qygo3hIY11HuavX4iCX/Pqfk/dGiIteMvqvJBXTOP82q1CU6gJrGON3Vs2r9mSw8
8d994OzjXDjtVOxuYnsE/B+TFPualBOZy+xwb+JL66onf0tCGzEb7P7UnNA/fnK9
FxhpSwNngCAyi5bmEa5mreCw2X+Z+RxegH9mQ392qRMOvedTYtnMMBd7c4z0ZARg
36F5qrih9rHtLJDwpasQzKIkDljnM6+cduD2436gPDV8vesbL6/erj+eerk1o+K0
kqI+xabiGiPpIwSj5Akkr+4Btgn17e1zJMMAI/GzH0LlIY6zKwuCcBH1HHFJ3I3w
4LozI4uFV5Be//nwMuTQ4IdHOUtGuPmKCYcLku9Lgvf3OH1OKPI5N0kSc3O2RKtH
tMLZULODNpnsxmjRzfAxJnqWRr7ckWUefihURDoIyZRXJmt+SkuHuhLjgc49dFCn
mK0O3jlMM9T7a18aVzvreywsQ6jCrSI4+hrnrGRStePc+q/A48wbi8c4CLboCDgm
lmKr2zJvUP5DS1a7lfTZqYOCggWmdjJstn+bx5p0KQz+2Gvvne2qjQSDnN+pQsQb
ZuTqv5hrhQwWfmjWXFHgbgU4lD3G6jzbz+cTk65grleq5lC0AXbkOigiu/i+xsSi
o6yHStBpLOmrCrq/V6kmLYsXdM0y0ncVu1IWkLM6Qqj5rHZEzBRsoK5mA4hLNXXK
yNCYP/6w7OLvaFA8QGeLVQOUnuYesgSuM3keVRVKZl54BjkOm7elV3MmuodRN+KY
aKa3Ll0QGv25wcbpxarXdsyOCEZnDRbRxfYXEOsTLHdkpJZMZp3lkEGU2Il9pZck
VNW161dhbVMM80MTAJOMN+7HHTOqOgVHwF6g933AEZQuMpf+NwWTumQJqyh+vEcn
6BwEO805GbnhrEG43hhoMmpZWnXcBMkv38r5sfHczYoE7XHMqtEG+9ksPvodcj4Y
EF/KzF7sxwn//ZwlrEzzsuw6xdHPFCnqv8h4okBO8Ky4ntchjI/bO3GF7YZK9k4e
7NQfa3+gTAfVSgMcNOMHUedyVtwuWkAC7jIO5epXaAfm95RGrfvVN0i9yKcBFedC
uCvvG/BLQpghb9mPghGt3wZ8zpX9zhW0MN/kWoxWQ9YsrKIb8HOdaWSBRS3kOz/V
hDRGfCh7PJXj4pUUTvUpIYT82YfCiJiWtRWeslaFBVAhPLNEECk2RQe+QnzuNa+s
lUaYdgzRpvsKFEw8r9cLvmJH/3jrlBzDR5hZC0OvQI2yzg6KBkb47v712PnE89Tf
iIYf2kVxknBFSKBTP0Ld7j0QkCqsf+KqIrFcOPY+76WGQ1osektjRri0stlrh/Pd
u4RBhnV6L+zRNGZucRbkbm4YRFMz1p8zX24In7HrAEWxf/PSKs6tr68O+5qgsRat
DzBHjrhV6W3qg4umzTXD+XJLinR6SlDE9S9o1f+/Yq+5cT+0FvwO46jaIpc2rbGA
aKR1NVzN+PS4brttZOsNd7cEOXGwlJV8OqaA5B5R4E+Jy1t90ZdtngzhZOg7M0mX
AFNTdDlmmWOQ4n+BewLkd1Cx9/3j6fO+GkqybpKFOcoHPfHyg5TcQ9udbkgVT/Bq
PZhPFRr5Tgl/oP8ZsodqiWud4D0EfNV4IjC8iMkxo6AHCjqqMiz/sGqvCEeH8QVB
ah/Dt9YnrGZWpH2QI4qOTEtnEx8riJSgJKpbo/Kwhl6siZIE0BLxRhr1AwGn0wEv
k8WXOEGk5nmRg/iMTNKf8RVo6axYokz2gVeabDjx9K2YE/FqKOD9VkvkdyZefp+9
585bXu4Yfu70YzOURgl4sH/o/V6tk7hTRVUHFPlJwQl028wwD3yek2JwhitCfMLp
MzRKyx7OWz+rGXEI6wRm4v5D2pxRbiRcegNPVptucoHFsSQ9kqGIqITWO5vcuwb6
OUkO/LcwaE8se7Ii1+3IEVRsgVkMckaWhz7PBYzEZ+cf91CMVXDBFQ8+as7v6moz
oXq/+w5jpxlq7Zi98FEo/zV9Z08YG29IGyFBjeiqjQk5XrcnVzct51I9HCh6HTZN
QfIvpANJx/HC1lNBszFFFIu5LaIk/iIM8o19blgiTUWLvRrRCuJWWY4cvy3BtDba
8x1yJIByoGO9HUWnmbaFkvwt3aA7yBs46zSeaedt43ACWSZmGBfwMAmWBopBKweW
av+9L1UXn3ss3dLL/LflvMXk8NEranyHvVzgapgGeypzy7WoMZHi5MTRsVe1TSMQ
Avt2K8B5iBjqWOc5oNCNAoH5u7xcAZOel/aCvIY6xdtdcyGWzFpn3kUQG0UNSQQ5
mnaZ9H8riwTc7p0TkSqYzbC2U5Ct52jF7YKdgAK0+UZch4Muba0YfLLwrA5i0HPu
5o1kVMxrYPNv7bwXOnQ8QsaIGubZ1n40arl2APfbNhfteYdnRrRUh9WlH9BghUDR
r6S3fENp6X7poMjsXMHREN01W0iE2QqLPJnYBZY1wGrZoHJT+g5sWQ6wYUemxG72
Miw/Xd8dK/x793nS1TwDF7/rQv+zuX7LspgGY+mJktDRXP7oFz4c0Z2VT+BIT58t
BTtbHNpGEqNONmVDkJiCLCmK4g9kmfS9UgB/cpAVCeRfskSnOdlA5/Uuy1yRXwIo
uyQZL2JS2BqoNyuzQUpoMpeCQQ9rI4THnNXCVlC1IEb4gfCrnSfln3v2gSSWGx6/
TllYd5ZTe1sz8DXXxYW0qS3wwlUUCvVBVwUTIECiPuZicXaIwIxnQkuc+CGg8Vg+
d87xWqAGOtUYZ2U4PWrCO4nCId3hWOdSgucbOtOylz6JiwQiMjunK9+5LWcRqwh2
9KamOgQ99g1gejvjE4uKb16E4rDSEj8SeDox/93evS+/7WypSAN2Grf5L21GbofG
qzHAJzFgLnEJwuLvAVpv+9IHT51fZ4EX43LQH0zxACXwgjm7xASm0Ac4wm2abE6m
FFboOVhoslKucmgcEW8jeqFyOeqpmPgLlsKTHkFgs7lzI6RNbmXpQ1NaFLEzw/kW
ojx9wgIPtyh+1aFfOri8johOZw6U2Yx41iLq3nFUBQCb/G8l2Ed3AqnkFaW2waW1
QLNTgMnrkAG8StNPHFY0NzpURGXgQYwaPmUUlQiDcdehWR/9pRu0ufQX1lUfYr2Y
jLOzeyNUD+72HvgojAELixmwXF3KCLW3PuZqHJJjVvT3tc2RG06pvSOnn9PFYZJU
jLLm7K/VoS/u/cHZMVC3+1iJuE4qBolMJ0hV8vjRGvkLLT/0/Ki4OsZO/6PPxVOb
Vb2EZvEZ2jsTkutxCDB+zqhXB3MfqRo6LV7jgEeCXIp9sJfVg1uukSvgd0c80via
TWuDVwA8N6IvEy5UPTdfYTZrrWZZKqhshhXA2ECH3yubc7BACjYsXtQGJfIk0boP
L6b3RDrQ00OEv+py7h/oOuxOCvKgeJTefiDgkRWMWzRpLKkXhqRt6BXeuJUnHp5b
KtpUEVdvuZl+nF3SUEDjJu41NOtTYsy5Gy5yGP1h6pI10wYsxyjaNMoFE1BCKZTi
2nKTPtGQOpfthKoLlrDRNgVtQpiwplIeEUMBX8Qpo0j5/obDn3lrJmnJGBiO1gRN
qPO+3lLEAcbQ/zD1GVZ4CDe6uV21TZCu6xMvzxwIhFyZvUuTbbhbKK7fMP2HlXU9
Ke3keZYcN2ytZOXm2Y7samMN7abVZ4LoVzRcjvULkuhB/7Yr54lhhrQSbKQaRFDg
STuOVPesPCf3gzbHBD+BaYIcU+xxdGuz1KX6rlDryXexaa3IL7HZOf8qt5UImi0c
e+LaxVA77KtJ7KYfAd1NFd7kkVkatJbAYzeJkmVWJdcoxQBlbezrFaiqI8Wu0vvA
WTIW7jPVDFrO2aEttfA12DNNKx8u32IuieEqjpEF/Levjc9tgEOG7MQoA+DqO2Ks
lX7RvOJM873GDftuQgum5hnIQ2EZVR//bkPYhpJz2SiIzVO5pNNvfLvsdLqKZDj1
iPXyquSvt2BH1C6g69VlnnNL44qOrKcRBycWRuKy66m2nDmOEPrkEFN4n1qLjxws
NEpdYIPaPX+aoA2SUksnP5BhP9zklOCFW+ffSSbZdimxWtCD/X8E8f+TSwJKsrTl
Qi1+pSgBd21piC5gzMzvRCMcy5RcMz41+NvKu6Ye+JMAJmXXGF5zpu9iAKr115KY
oNDwFOVsHW8w1hm5GdT3og38ae/TxG1e6GqrEApVOgZXfXaaTTuFiqUutPxwHgeJ
InRJW0Fr2AJAhlL3JEugbn+VRdURUrz7qiwhC7ByzLQMJB/JGL/MbQR84X0c0dj2
Qt30gcJBEj5TiL7ICDfJ1Ilim7rSxhCPmwlWxHGw5ZouiS62Pjod6OC6XFPGmZkb
u3c0TBxyZhJvmxUS4NQuW0fPU02Qbj/fT3Pi1K+9Mt6YG4J6MRI17808xyLLYqiE
im4znsO+f6SkS/wBHTSY1BOkjfq0o4Yvwd1ruibQPIc4byPVjAfhtHACysk2e6zX
XvQ+912VlowcPO1yiYgEm9JiOqxz+k2e9e3lMhdsdbUZN9mRwwNsrRK8x/zs6ggo
SUXwdhmyLC0BbkG9KEPhbHgcu7OqcQDtDZygMAIKxoBZWQvqCliDjkKEdsFS5w4r
VKx1vWvdA2mRWPYRiiPNlO/cjTsQdM0i/c1fPj3ikY2sa61EXl9zGOorfB6nCG0G
KNaEgaKPpxt+4DBq5zcpZykNGs/Rv0v6PYQ3by0JN0yKF+RWBgnFqUtE064hfxf0
1julGHeyVuGHER5nVjO6NaN0NDdXyc3uIO/rZBgKzoFEkq6Wio7Rn5HVTDPSe/90
VFnI5OxWYcq66tfHvQxw+dQLUjzJtEjtbVo2Tg7WUcw0wsTuTjT094RryOVzPyVh
eKk9HWP3ErgSZCi87nMAhDHJfFvyRcHE1aKocutprQ604+zyLYGg0mNES36yR6om
O6yw2VZmOJKbiluLNykbKuzI9hiENEWEP8Uvkoos9WgS5BddztRwlCOcrh4cO1Rv
QmRGwawjf1gPr7MWg4I9pAyIn10BMDzCTaqcxnWFFkU+0mxX8yJvqZ11SZLlrtCV
OL9rJjSARXsGzSd+X8JUT3vOaXwzbZA9rKXE09thDotWlNL31G6icFK38qnahiMy
KaZKbpI8JU0EYaarlryvmLLWueMrwicaj0fu82sC4svx6bwxVaa9XOzgQbbG3L9o
Ki8anTyS3WruCcfNBL0SvGLn9ByJuJvjg9CQSwpM7mEY1XffIbVdP9v9t8RY4LUe
1hUz2wyzFvgQRwpgOYjSezR/vzirc15j1naHTu38ZdCcDB0t3J2HBMWmeKnizxSn
grzaJ0pFkLtrX01aFoucMiSRDqYam7WPngayBWt85H+1gDFXYd0y2VTpD3QBP+Np
LV1+b0ZCdf5yMs9F8lzT7GfjTIcV70n35BN3whfwt2MbrK08fMWnL+4GQ4Ve3aQ9
G9BVbxnOR3uSaSQXk4hvr7u7bRxGtyHtDkt5fRkj3h4pnaw/ool2woCFzRsFlQ+3
2s/DzylWsAmF/sseDtk075ZJcb6cVFlNrb47DIaz6D14jdoMz0bmmzjw/dPsKsx5
AfhXmknJrWgvgK9Elp+TjkJKZPxEn0mLzDIxDn8q/8VG5sfJHUUVTiPlYkDyVbSZ
7smtrzm8Dondany3YIjoTBPdVp/7u0gsRv21siQMyo9tGIDhTL3uCa/dHilvFCry
upqwaVmsBRwyYenW107P3gfELFhjWTUl+lEB46qIG0J+enx4q7VInTy9ww5zec87
Ev8iT+3f1y28seSIe/2oiy6akjjVhgtbv+IapVflV4ESpgrgVYHn0hvLK41usVCH
CYTWG/jBo5n34t69yWFUT7nPvpeJg9Nor1txulSAm134X517mcRvCd96Z2+Vt3+N
0nG9oFznkEWEjF+rhaNe5pO3DbsQCmv4AtSODxthawY+K8eZoCi4+Yw1cMlLSCru
VfzQSp2Nb3pJ4PXNOnoba/1df/j8C3T5rcZEKNPKdXxfPnkdUi+sCvvgQT4XdUtv
LVigBEQlll/V3r6E6oHLGF/JEB54eRV7LTZEDw2TREJ/dx6VBtkaDPRwAuM7Ggir
69LmYExQ6eipc6bzU1xnvvaL1iszWcPSAmicUuMoi+WjfvNpIwz9SkZXBkCMOOCZ
uJVAt6aOq16fM1KN2EtskRPi0A3l6hPfaVky+vJrbQZeiS7euZj0o82PYWJYHIgs
ZHdQYlowIjrzsc8Mg2Er7YLAskfQmVLOXl9bQ5CE7cMuOYVeuWij9QGpISd5DfT0
Me35td5pypTNgvtcWJQ8gzfR2r/z0lqFM91zW7Pah+4srzVqYtG7iSyVK+E4vsGX
cMmbF/zjBWJEOwu+AtutNTgwX0BNhrOLm5STAYQ3Kjyz/JzwyaebgmTYyvwrb3rS
H6NODgz69oIw0RpqFryogTY/DFyomp32k/sJHCAJSCOSrQzXSasjIoeiqpd9nQcU
avqs46lQFtfgH5ulT+oC/4Fj2GPXfQEm9eO93tCZDu8hJM6xcOd/EXwdrt2SDcWa
/XNApH779KPe2YBa710rEOaP4gFILm85DWunUMl4ymCSOdgguYSh7ja+H2NHYfIZ
kqC/xbIRBHh1GMa5Q/ekmKLJIqxOH7kVVzYD+G5C+pTEppfCc7iAPVoLPaggjGjr
zSHlnkIJQ4dXl+X6S5nZOSJ16YKc9VtFkZsCaXhz/zclwKNnWtod26E5Qh0aprVV
y27rIfCbPFIp+W2paLOvHMavoXmwzL8LsZq/OQR50LR4W0UAfyXsoDoqVbex6Ged
6FpPHQDqWS59dnXw8g2bk9bqZkLxS71PwckCdBKGfDzpzfTmN39X8agd1cIDf18C
lw1tP+GKE8LtvrRQk9MEC8hprSn8oTfEpunMTaW5gatEemf7rg/wNyh1x8vPSyV3
0tFVFSOngGBQSCkZ3WkoOwlxbI9QmMv0DtXeZUE8B5EA9pmgrgMlYAjoQMfh3A4p
BFNPPufDtol8HqDmQHJHHNRQZ+x1f4xmjguneYHws7cC/kiRu6ubiS0/ix3YlKFf
yworGqwUJk4D6EyBd9iVotQhAbGicIgdaoNNjxZ9TV8iZJLCEcbIeDV3yZZEuob+
Y4gf6RiTgF+vKn3FIzMpkYLjdmZnY83gKWEXhGMEX+uQLncUqaB9xcmqAsFUxT+2
gAqbhjoL6/Cgy5a4psdl2TCnq7EbHkxIZhsYkamTHGbEkVszT8RJHwh4TnAXimOP
g0PukhJ7b/el6JUOgiONEmiyPvZ66iE6CjSw2S0NNdoLcfpdMigdgD8D45px8Tpg
qLqW5P+wKS+XfLJt83padCpJRQ9/Tn/rCVQMDgclJPrpJ780DF2kCE8N2m611M8J
hzrY0BaYOW7Qty/6MuW6pYWUKqAxybr8QXke/Td3IwvR4gCqSQ7nXAdrmWL2ZhRt
qizN4sbg3OqW5sZr/z5qlP4/WBtw5tUV22dKqB3ezTqYPVyDyC5Vntz0S+xnKULJ
zEqq673JUueENrx3sM07FUX7+HRizIIui4gpQyHBLFuQHFmLyuBKURiJWaH3tNaf
FTsCA16w2smY9uRwrvrJRJuGxInu1NddcnCpcJK5enNFBqHnnInroIUg8VpNRaAa
wPLsK74uB3RBociEpPFumN61UerO98jPn9UutfIBEbmbezNby2Gz/VPGBD2xKZAx
lS/suxrsyzGtvRb6huNHZLP1oh2C9pgrZMoxOJsykeYFqg3v7ZnGzZY1Lwhgzedx
1eLpjf8gcp3CTsmk5MtJHR7G8MP0zYIRwNB3L4LHV7Dve9B3HJD9mqULiairPexc
Ve2B/QEdxh6cpAeAT6CIthh4ByM9WMHfqdpJNL9OqUtSIf3JX0mS2GejEEbrg1m8
yX69oo9QVgomTj0n62HZNHXqkYwYR1SaFtxPbdfq8ccPuG4zGUbqX9HBiAaUeepV
saOj12quFpa6nyBQyzAi2ozHg4y5syfEsoLlguk7Jvqj9O3iQx4plGHT9p2P9Vvz
iUCeGVwZR8oxWKDoscWUUkwoIff/GIEh8y52iu07O27AUtHq4Q3Q3fMEU94DxEVO
cIpLI6V28z/gU6ZykVWjJos/8V7uyugiGhr8DrRBwAPFGwkD0iOR1s6bqK1g9gjO
KjXkjZ0o6MtKjf0XOkZ6EkvPPvqM3X8ewx9WAvxZSCpi7bZEkj07oypXuWrrQAPC
umLb0hbOuQjii3405HpuTzaCtAFWkxvmACJD82kG3PVvEEiB1/C1ey83k5n1NCDA
HPe5N0dKesL1fxCA+HOklcEPBGqFM1CZbSxtHmIe7tomZe2XCCTW8AaOgfrMo9y6
+IQyrZvyqXm7O6Irz//hphg6YkjAw5YBh5+DPWsa/W6zlJ2GhjmOH3sxlKAAxFqh
lKQKQzKBnh6yONQ/khWLUK22pSEi4S5y2yDX66WY0YrCVIDIBeQvQGtzRvQXenpI
wYiKLOaglM4fzfG0qTqsFosnNdJ8H8FFPzGqlKXJP9bno0KpBoQ4uNKUSjZ2F6b0
dw4Nj+DApfgNq1/mTs5tPKLPjISX3H/hG4628U7BqN8nd4+v30okXBku65Brj8Lq
wGM6BPYg1kO7KtSXwMe5tmyHzbivgSV/waRgY0XVdKWRUXmn+2YeXSqHcuU3eguD
qyJigLFwY5a3PmCEdHe8e94MZiV2onw0d5BGAbU+zSet98szVzJYLkc3nr84oNUL
DqlBakGkFGZv8yqfyzxeADT22eWeSXSzhBY2JFYxfql+N5Tf5Ei3pw0Vl84CzU71
DNcM0+bmMsuDugaKOuksHEh3izaJGlsZawxMWPsiawcmPJF+He9CsnTlE259+5oq
w1fKG5T9gKuuoVk8jje6ZpOilo3rp77m99IVBHLcGkwXzlgz4V2efn9FiLcB+Kqn
QzSL31iPfDt/q2Chx7xOlAyV11hjHN3S69L/firuZ/gHy8mDa2v8kLiQhBxzC1ag
OQtrtbreZReEeXJQKY8FD/9oHQQdUDi7aGXx3Gd1o9G8+t+8tCIQWsc9OEXO78G1
8UJ3IdVdZbLMwjba9Jc2vYTzFFImLa4EVSxEMrfWw0wRRD0Y/+rf8QVCeztgpz7t
lhxczvLzxrxwo248Ml33HrKBcpLisiEiNWZNxLEEF6BfYXNQAoUd0Q75TGB55CYu
YiiBKvZYY1IIahlZx9Q3nsp5jisEvvxXSZ3bpazajJ04PV1c25UiTV1sYAiyXIQT
Pdbt5EE23JOKbO5CDlbP+C9Qz6nAcDgYsdBatandhpFCKf9GdLSytze36pIvNtwe
vldvWtfrDPJg/vm+Fy6mFuZ2GWBzQYesocs3tK4pNcB/h7BLhZYcQs+HL62xyne2
bQCCxYwggtl/a43upVMNyW7Q8HPymGsbKcz4JnuyV7xBMnTekc9nSTR/I7PzIaeC
3alBeKOa0LGn3esayimXwsmEZHylQVj2rVZelbsybs0UcQbCKaPIVpK+MX15uwHZ
fh+1aBrqTMEiP5ZtwIoog2p2TBOeK/Sx/WvUJw5wf4XFwLCx87KGT8ezpY7pOtsA
T6kLjqQ3pmxvhi0UIMJx4RCPHmPJrH9VzRcCtZ+nGfLt4JvXAIVdQcr7D0ck+X+E
uieUJVL9yo1iBv5tg5VsYjWUndgKmzJxa155A+sJ0aiTMReor5nuMqzl9q5N07P1
3lkI6Lc16eClT+vuXgW+u7hfm0Ud6RhkuWj3F4GzOmHdWqXkfeNCJv1ur2+hhU3C
0WHMr4UJPFJioIXKQdXL7xGP75uxVo7k5XFLPAM0djb03OKhbCTFwT4zEu1z6tAp
euGkOC4hz751Dj9jN12XtfZmD9137+7ANvvQS5B0xOcvbhd4HD7qe1i1sgmYzh08
yZzGxglgWggvqVo4GdDivkv7BKPCKSlAKCu65lyeaJzH8oFfkzLgZqLkO20PPd5p
dhPqy75WIqIv7O7BHlJ4UXemWE4uv+fGwOB2ljjAiSaGIG2eW3IHgrqwg3bxbwT3
BbjAb+vSU/RD2oyrvlhqrVE27K26a1DMSQOxO8ZWbh4TsD8pQPPQgWNPF645vZMT
ygDxIKiwHGD0gYy2KkSR8yHW7YLYef/MFNGcaYcjp+UQK0uoHxvSg8UIUOtVsM3m
jJhbBCFxuC83ojBwmm1vTeLJq/99d+jy9v2WPanDR1UuQALqu1QRlrcQo74rhdYv
TMTrQS19MRimFEOtS33fI6zpPASwt/yua4HTIwX3aCnuhDcjaPMaJ+zRqwb5/RSE
jIBmNH1ccvdsVOIqoG1TpZQ26eSszqXbcD4wriMJZEwBIzz00hpWyTZ5LvxygyOO
RvGNbBqJvw5G6PuGa5mI3JnDXJ5FI43DtD5j2idwt1ahSv573no6p1CWMyR7zDKy
GqUL3oz6cZK6h7SMmRxSrTsZ1dfKKeJd7JMglJrc+x/zYVLgfpKklYrMbUNYSJPs
yiHV+QvTIATG9G69iBvw7vdwk3x56c24cv0o2fNDpumyrIqhT4wbj2qWTQ2XvwBK
opp82vZuwIViU+DvLAO0xDhhAR1CECVu9oeonLh1RLc2mso3+8fCulHV26z+xbtU
KSzkiuqcQKoGniU214Hd3N1KCpOWjDS25woThplOsq7F0UJU8rHnZIhX0UlVtsiV
hJR49cBE4dh7IqZnERA/ajT46NrSBkO+VAKLr4iSkZZIdrgzwWFRBC9L1SeeeG6m
gy5x1S3kl2x/UryU2tE3GqCws9HXXB2ItM8eqEzjTSPxoFb5CKeJA9Kl96sR0UbI
q/7N2rpIr5kxqwI5N/gjymNWoKiIh9pCYkZ9ddVgmf9yB6pKfN3mbUM31f/HzpJl
s3dXMsd4AeP7Vo0yGo31ez49o9pzwTebHQ2PqT3lqsq6Fxw8z/pC6nV5fOi235Wn
VcQXWE4Hmm4FXibHcvRaNRxW4YBu6CeGyvEx3r+L/d4drYhbBTfDoy6vRluhuht7
tE+sN+NuYMshJdq8XefFQQ7MYAasBcnXjFtJj22vdk05sMUBtAXm27cwzR0KmGQK
robujnefCKEyl+jWQ5HOVNmNnMmwSDEsDBtdMB2fKV6kAkNvw+yDrIz+1BcEYtRh
fR//IVGYlbzaekgqkNsuAjJvgfpJoQc1+LSHLIieP0OLCn9fHikc+1M5heVbp2VI
bGFAtHnBeiiJs13MLX4C0GweSspXWmA4dsl95JcOfTjvdBZWEdhFOkUFhXIWAax4
eUZYnxKeiaIGYJry53ktUUs8dIWP8A90X4uC7WNbUmrfRPc6aorgGilyvjOBxxf4
B3V8TMwBQJU1cqEBW9AitkavFnhuh7mVbv3/QBUNeJfI3tLH8qi/dOaEWTkNKc7S
uLb7zEd32Fg97wcB+P+0vSeFKgXezAVomn8oeM7p2zvzVuFZpZzKOvvE0fD+CqIB
V6J0Mr4xmCNaf7/vLfAGVZ/5DBjRNN7WFYCJAGT1/3L+E8G8EQXldr04nZi0hV55
o+xmGppv5oA1H0bN8nixvBx8rP2rONITZjJXs5rsTD6k3Rh+I7CVuiW8zA980gOE
KruUxFUCtopS/2qwAkLdo75pPMRorvr7qhOQLQien7ytvA0j03GHKdKLDxDysK6p
YcjKEEkrxY/y8VbA6CEYZex2NGYL+gWSO+KtjZNFy9WMnv1agsCTGO65WdbBdBRg
AgxxRsMWK019eE4KVvGD+n1ixjdtifQU7G7wHxn91/OoudTtjtM2q/+RmG1vsWZT
y73KIWISlNWJ4rDiBfoAeGF2z9a91nvp1PNQ35afwHANseCc7HXz0TlI9bCY9eeI
ulJvrPOLlN61ehDndDmp8irIagDK5eeeZDvC5v+CGK1Sf5QU8BTdbadVHXqrUkJC
xPhIwvCZn/aejx4hv3nBtnuBUuppxaUzTll46jJPUpYHYUsS6swy+h0KWRiKYnlh
n3g1xQGVFXiF5jrbJu1X6huZy4/TrrIuCdbPA1QZltIT41uHh4kmq2HDze4aFTsw
JFWQoS9Ij8oXO04Ks2Wyx8GkdGDHYhtUAtdw70q3K5JODffeoa7L06I3Zm3EW2/t
tJyjuxD2cF6ZdWdhFQHeiTfQ7y1+1i7Dkyqa7+INZTPuDW8ZTI58HPwENrkEyoLF
k326INyZhzq9VW19gHNT3MVpdXaibbc0zzxlo6OkGZkrxk11xVV0MQ5X4PBm6Vyz
VpmBeZXiODA/1C9we9yy3VALF/3u3JqztStqEME++DIXXHQPCHjHTJrbzA3uRm9N
wzA04UTVyhOTSFIsYDII2BnQgJ3oYs5D7/7ihUxXLj0hwoJt8gvuAtz+1z1W4wLS
1j/l8e6OewR4wV5AZhgU3ePT9611jcLKhcpSrCkf2NWkNfEnQioext+1pwdOZ2oA
in6ygD/HAFUyjUv1Q6SwLdsTErks3uaO22OdKOR0pzwlM8jCuZtWRaYMt69hRQYW
0HFpQLgDGuOvjuW+ANIy77aexpwhcRSQuq05aBLnbcOijemdWRuc6pvYVjsQyaFi
vY3n3J6yuLUhGBdojhsx49Jw7DieWKORzLv+5pDnTJ2VGOxPwMq2fTw7XmEUPoAX
efTw3RdPZH3lrz2rsitvEpdt97FcfJttI31ACba9PJRIZVsByFhx4uvWgKICmNPI
ryf980+jrIthIJSMtDLeR9GOSPFUcITGRGd22cWbdGkseP0OdgCkSgAwxOqAS16Y
6gW+weWtIl2Ka62Y7QYiWKHAcxTVcH7myCuNklBDyuhBVaykSNu3hUOO62h8ypZR
HbP4uNAem4Ru9fKHdRwOfXaQXZZycs8bPyeHNyvSZUtSOId4fYydxzDsrEcnLo1a
YCSC8SOGez923qCMwszRD28UQleQiDuVRBE32Coro3gDMqzWongJnuqzCu6fVreN
VjJ4ftn9j0qBxyKmnkSpKfV3ejFqrh6K5xTF1E/nY5Y0KEs2l3LMFFv0U3o2G6DS
1s3tYDGUCz8201Rr5EqaK4WC895jNY26tF0DKw+hZKQQ05ZxXAN9etc/n/A82f4i
DJ5gxO41m/wZNZt1CajUkTUOACp6w1XUL8gfRSjsFKYPoREVwWf9Qze1IrGYqYSB
Se49ycCWyAazhbZ02y6rRgZeO2gK8nM66j9gSQFPrPUuh0mmmT/pIPyPW2rLjbgx
MtcKMQt/gCFZdcav8V8Sh/aek4R8P1iUm8pK+nIumKK1zn/eWTrXUlX8ehrQcHen
zeesrx1S1/rnP6nkwj1+frk/EPoCY/mQzavDe0LF++6tbmk+1VJAxvw+5slI+tyC
t97u6rnP5MzvE6Y/wlINqtIpeYVNm+3Yf81bPoIjDz1n8nPoCX7xnbuJ2B9cvafY
cIVvj/Ac6HBnIjJ3bu2R7Z3cG9ng6N4X20nwDYQlZJb09+dN0n7uLcxrePE56nbY
g5fFVHXU2KHgmnAwPN9w1YNbnYX61EuTmtwjHMM0skWxlzP6wDbNSws9FqEZxmI6
BuoEYlq4aa41VCTa6a9PtdPbbnS5myaX7/yjzvqQUcdQXeE1NCTbx5vinOLZKGad
X1/abRIyVBWPoF3mgdvUijsjKv3DOJcbXQQTOWQPRAYec6uBZvTAPMxoCOzCvxSC
WFx3e/b3uQW3UcZgujRyqBjOkmcTP2m3yPM2xVendN764h4Fwtjr5eQgs26w16Un
qVfq4UXu33YqUAFYU9KIcfAqsPOauHd1wPk+PGrxgyLuY59tRTKzp86ZGVEITQOx
/UoH0JdxWEyti87GXssSdQe2qGYjdQ2YggastrlXRetGJEhl7DKNiZwTY/Cq5ZXF
uNJN3FqZ31gGbIiu80KjwY7TzB+AHDQ4V8BbZa6wlRycVEYca6pVZmD6ZnqV8DYr
3j/KJgW4kw3XbOp3YoMnIgWYRkVoyZ9xrrX7qD15xys66t396RFauxTDW8nUaP4k
VT2R/0pgq7rtU8iGVf7Uw0A9CV/HrhgQ9BgNR/CLtBdzsaCd1aeYAUnWt+SPFKpR
6HnYhja2BW1wzTDTJ4FK2UyHe1EN/ZpZFAJeXDvmMgP48YVVooEi/yereHHUZhLG
QH0k3XUdoTiWhlcYqeaixhoMpL8F8LsVFV2puVHRfGAm8hRiU8GnHbr0YdSooSLS
aZPvq+vs/rTQWxDQ2N5mgXBtiQCTiztItdqWE98S4+wUsUri/UytKpR30PJlyWt9
svNCqlCxK7V426LFzrHIacUkAQt8QzmbR4VKz+66LOpWHtmZJQAImV4x1+qycz61
da10gqQVhwG2jB6Bz8s35d+rA4u2Fo3kHpFAr7ZZHUrIUBMVm0E2XIMcFxeuK+Mi
znqhJ52VtJDcYv4bt56+0AYKeeQttPAYOL9e/lx+IhkzIadtzJt7W+VrxlXHX+EQ
944HlNxbKSJ/lDi/ugFGFk378wUYkPu7r4UqZhi+KMNkpmY2yaHLnAkzzfs5ZQkA
JRTa470xc8N7aMXODYWNrnhLbyu73dHgHMxAw6WuOda2QL08ioT13zjIT3V0rwb6
nowSjaBblrEQ2ootfur7gDxe2zRwnarmRpz8IDK13kkPuSKFKggDKYadD3f0WYyT
xsAvxrwxv7ZyyStoJpj6vTwG/vdhkjYFDmYXwXbarBv3GAi/eSIoNZKYWfeKWRR3
UfI/QXsMcEVbFmDA35yRUWZ0337m34lbXMAtwt0hGNPhTHgUIaL0h75XuNJCaFAu
AayZa+nu2m9kZf1eJRdx0ZhTOqPVNsM6oV82JGd8PrPRT5NzATdGHj8KOsdWKuqB
HhbOkmOfMRaBNBYUvhTldWFM7beJzzaysIbCXAvZh0IaSopSpdLAC+h3F2mmNQg6
DdJGzMwMiYoHsB9UQ/sCSLKFE8CTVSAa1FeCjQDysLU7CDXRC0pYKh7JMM5hy+/7
q32lUSxp0hhNwxgOMHDKrfpX6GnBQNtmsJfJLyYwJUQ5+K8SH4423EJbxnzJ5XcL
cHf9WL9/FS+ukfTPjimDMIRcPIXDVcTnBv+DG68NIbhxB/ueBqlkAYFQchlytzXg
eiqZ3T/96WDTHm3md2bySMWI7g2q9pyQ/y6SGVG6JIVcfhV1/00uNa1/zyfK450h
GmDIjCshkPFHKJ5Lp5d4NX1WJLl/xrjUJTFi5fN0H2Iu7P60E594VtjIBfmm7HXx
U9mel2zaMNy7Wk6t2+Rmv9FrDsuG1vwHx205Czk++1uy6ASjP7zgKI9SS8cCx0eK
y8+P2JjwYClpz4xNhxb7y08GpD4i6ARS+4b6HEWQOu6wVKuiP6GuwvgL7Grut81Y
0B30EPFatGwL0Hg3zsrVZiyGM2sN9nwvaYmBViJoLE1yL0K4h8HhqHiJYU+qK15r
b5RIbgJL6yTodx4KsnVYWKvlcRHmaLmRK1C0JNs8uFECRjn81T6wX+4cxqcbDIwf
h9Oe/Bf38JyFI3LZGciF4xSxLf3MNe4JC75Rjo0z4L1td2RZdmXKhhE2+9OzUFWl
Zj65SAItcYTUQzfppy42p7GCx67+pjVmS0eH2KQmP/X2gsVZoH2HgXSUAKryUnwU
rHGh+ivf10nCiny8bbQAETw8eqB53NBj9VN+ZbRWL7qsQFkZAIwGz7qAMXZ95qhs
aWAhZkP5XZCP75HmsHcaSlasbkP4327nBRZRNm29ww/Cy5ZXEwaB4G9YCgXC+tKU
HMEAhafp5T3jkloFdTpEdXp72pjsOpSPw3QsyqqP8iXu82kyxOTmowdNW1BccKpM
vVZBQat+tsuDmZkdZxa2YCcrc7z5Abr38KxievHq52ixCXqcUTTOAXPe0Cb5iZhN
eIvDngP+QmvXh2TaxKerbXfFGt8Og0RuSKTWfHSyWXDQp5ZC78dDtVjxdJ9w/DI/
MWFDJ8ez5nNawulljtr+xGH70A4KkRVdMk2MM5OYL935SVmpMyHzzxlnkShMl+Gs
Z+kJ9w148OtuyERDzXXL1BAGf33NeuT/vmVyPYZqbcq8NYeTP8BCokhoC+fn7a8z
QhCaWaryw+p1zkx2mJB1Sptbu0pp2tzAypj+Grl/+KJpw3vdgK1mgwJdhdBFqZQ4
fHPWhcNTD5/Ok8RFVkpTqTOqCh3T1zVEjOldRtfBh5Sh/cQXrBzIQnjA9SttRo9S
ZdO1gy0D1Fot2twoZ2DnaLobMAHxJE49KmtGSwCO7QV+MD4MJ1XeDRHVW6s9Et4y
N0kGe9v7EG/7TOjnnzrUaSlP/Bp4qHgQH9GGno2jJ7u1jfFfLzjDoSZIG/gRtQBq
ZNqsoRinBgWjfNkspW39iAl/Bs9lCOADWaulcFicpJMCDXpIeBLJvME1M/S/U2Pj
FdCp71ABMNR6dbNPkgg9d6j704Ct+HmJ3H4T0xRjrA2t1qTuEG2SHe1x34b0nKqv
0EzeRhneOiyeb3m0q7rIjxGxQkPYMsE5Vx/6N5gdb+KD8Fl0txzmYZltjfRXuH1V
PcAPpWd4yCOEMPNzYkEvxXGZgGe2crZqqOIlHo0gwlbg2tYOAhdV7KOngC+PYHSB
m6zoZtlmxATz1d/PG44tuSJ+CuCH25PKr2khw1CUxPN0JCl5rkQFPOLLyx5E87oJ
fEo2KW9TBL+lAnSD+EL/sfXCNi6HPCnkY3etfRqr9XX7cIdQXl3ezxMz9d63ek+b
oNSCClr/qHiM7PY428ptjOmEJNMU7tyevH+jnRUQeX0b70EYMsTKaxaPWvSZb8GS
c1Kj7spzmwMNrUbcvREgib0Oc5MsmTZqUpBX7iQUG9ARN76nZ6OWE9h+/6pemQGL
hwEyzxwJWPftfTvsEg5LiGhU4N1uRz869dzt3adluM2ZcVYEGZ4snb3Z3NFbBiip
Z0fPXxy2DK5y3H8twtwTd3hlXWrsaWUlcTC8uHmabE7RPk/RSS/YuErX3cpNIKEP
0nQOHRnAdTRugow854YjstBm0zvGn8XFPHgAswXxnoj4G+J5AvoyETx3WXM5CFK7
95e5XeA+oZsSy1G4vItBZtL51mXqc8MJCRL+qYZw1OyJwjqNQeuFdaxZYsSY02sa
VQJZ8UgPQWyPG28wAjGN7YkU1sRCuni6ZTouRqjfhpRHJYm8aCuszEG0XrUzklfH
TcXuXPdov6obGnZ1eqDcQN94izfBkKcYOYI5RYtQGst4LXyjGvdWDI4zZ1I+8D3z
KVwsNgDbavTo0ESWuA41oiWAIDBzxJBoE5FHb/hhJJxCaxJJvI1qWLOCyR+RYGct
+Gozd3YNVjAts6gFN3CgK1dWp/d/jn5AJZ2I9lAouaJJosAKymDhdb+9Djmmt1gO
epvkBbFdbroAdhnVVzBAIhXHG/O6xNOfWdEdkgh1w7pzcOyUSZURIxyRnJbXthAC
1Bwbue1V9VIKSKkGfrqOWKjGhHemByBEi6mnjf3MzmwwrXedCDxBtJM5C+8oLEDk
Q3FvBuj/ZtVrbubob+xYwNxRfy44hNB+7IUCTmtgtkBgbDIp7FzFuulIcQyM6Olb
RIxe5A3CYHI26yr0B3KriiXIyIqF6IOBUFyrz0Laq5pxW7aXFInp6bFnZiqTz//W
aNd1bOcRu7AzsrUq5Dn3OKsIm1gNOKf8ZQ7Nz04I0nmEaoonm1gQE1DQsOkbYkIb
8vSgq73a/5AtuZ/mr+aBn31gEivbuiZmjoqD++4O4KppGazUZdPbziXhFL52+4mr
TwpmUV6FA8CLhpQkVmnpHPscrPigr+RLto5A7bWLuEDsG2/0okRwQMNOR1afZgto
NfZuSpueF3UMdZ3GyCtuMbk3CXhqjfMlmThjIGzNKr5/yAEdCF125zjCJcmSYoYM
b7H+oBgR9Z/6sWDrlLy4OGyf9BKIUWe42q8p8mvvqb3vcfwrHmLUYIS4QvHgSPlq
YjsRdpGlBWw+E9e/FQBg7R5FrAGcmSm1QlQFMMB/ddDZxjtT1ccW3THkHWuJFU0T
dUaGea4s61LBm5JuBMS2YCrRoSfN+QrVghFVeArDDv4T7h/2UNVRBxehmK/iJkYx
rSm0GdsRX22WuHVBrFXeQh7Oke+xYm4GcK4XukWP5Oy+6PWWVssU7PdApxCXijfZ
ubg+b9MmItbZXh2RGZjFHzkDhNKM8rM2bWr4OKo6F36biJPbnqx46RWA+tEagygu
veGWgbgi3UNIju3wv1tcXbpqPbn39eUHJbez8Sh9dHvR+U+GX3xOCdOFRrZNcmkq
9z/wzZ3em93vsEyue+/XcTkd01nuqyt0Aw6AU7v+RtXhKUuCGkHdkqWZ29mQJ3uH
WwV/l+gXCU5OCwOozrkSSn4gP3jLqgGaMrDVTEWVLS0mLERIoNeG/tYs8SMUXq37
t5DPAH6FKMJS1iVPWkISHzmybU0ZMSCx5aKpCfFM3sTbA7c6sqDX0pIoRrK8VBEY
tTHCyz6VOdLGIIZ8igt8x020Pdfn4aYPgj23Ws2ibrgvqCyGyXdtfcTQnlDH5Pa1
v9AhZSer4m0gZcNPCNXSCxT4RvLppPvAFwzslN78UihCy01TNj+8ydRzIlbaOXmU
uGy6PsMhzzYj8qZmaPLi5c+5S14S2PmVseHhfAQaU4Ud3zb+Y6DS4vUaPB34aaV/
UTChWEwYeVJohI/T7t/N2S9qHOMo/0EQG60J1Co0UD/7Mc02ibYx8X/FaGjDOB2G
+PbSDqwRlvvU4NwmNCdD6Qf7MgZEJSWwM961hNTPiYvtbd4HzTjl1d6XHDFvkuEJ
hVXuNKWjoB+vM/LImXnj4kjl6svU59u4bV5fcnyoaGooC1410h9QgEfx7BHvoTWn
QXI0KEEGl+y7Uu5YqEuG/v339Y/mWCjzYTnGh48kUdYr/4hiSyeJVx8Fnv/3xqP5
7LqlJqAdrU+vvox91cxPD3J32tPpIGPtqKzfewnAI9BK4gWxiUkxSBzZFV5WbT+H
aDqVPp4RNMnw3I+Qad7A61GACf/nuCRE+FuXr25++JAK9GW50UMKVNZ1rcVbhKk6
PkCkqu/6oOYRuMAKHNzK4gF6Nb9E9BY7w+lBIp9epsJRQEOkrspfesoxrDdieWkg
v6aHBGFLmCQ32RZEARVYtbn5BfFOJaonOZra/KDUVDrv5Iy3Do6OwRk7gijCVzMe
BONqgjvfOU7lFevBoNc4MLLbNXJ5oJEOct4JrbssJZUnsX7SEmSiBXPPg01Owlkm
FgwKvyc6GJA1KaPSlrLrEOhiG2SCJ4QQNvSmQaGH1jsPLupip0RBMB86TLizaz5V
/k661Z6+LGj/ur1MMDPOjU/BfkTI1ObCSeDj+S+V6HB94eYZkBh+OBMWM4YixXtw
+SUaAyzh+ynzIbAfVzGnA6riHGY41Uxs/xPFW2NDD1xXT8TFEEyymMsF6kVzGDsN
kpT+EM1J2xsnRjYcsqG9rwOmJ9gF0nZ3PodD9dMUG6TyypfYD89yOZTuSrpCbx2o
893v8ito1M7EhPZJAxfhGSpjGd75D+gh8XXdDts6kq3899qxPz75JQ478dFRvvRa
dtb47B/l4NicVxlv3X6GeojttEe04APkmsE57vYfQSZmH2tqg4N6W++Ugttda4iK
W5hrLCs9nRFzezUqO/QgMuRFFzO3GBjujPeop+oo9RyHIsPTyMbDpDnCJE2Ck2Er
jzwd3l24oDxQs3lKOyBv4+9XhSnoUjusinRsez31TRcb7vvWjGfEMpQ3WVFEYewf
OB/pKFm/zbK5Yezkwonjt/IXdQB4hsvMintkxOJc19c9JbvoEvD3rZqsSjLbfCkT
tGueDHlfEW6F4Iupr1y8+qx0/OHxfP8KrfaSl0PqBeyJk7DiA1jQRDq8GIR156J5
yS9rGjVWbztPJxxO9tvyh0UI2Uv9UL8B04dPw/2lYzQECBjKnIfDKm9gJhuots8+
if+EIJUcuD+eUBxseLDfccInHO3IkwlTsXq/pYnCTfbc0pwU51jCOuym0m6KTAkZ
kgYRjEzLOCFHZYL9nKLgZeBzQO+iZUuJtlk+x2ULZSB02Xf18c/rYUZAFi7+owZV
DOW6LMllAMEJaXUYt0HX4dZXI8y4ahccgvIEyR0O/RT5H2IWaf9P/05rH63jNs+R
pQqI/LTjv0SDppiKrEisyW3y5lKhtee9GsVmchtFuD8UvKDPpaP7jPUYKQbs5Bk5
sRnsnz4sKqU6gl49YwltOLNLx9HIkrAupavxZx8BJgewPH3svJmj2PCgt9JRPzOn
2oZlA7sdp7ltgrdBslriGtbQXXwf3Fci4HsBH3gmSR9fh/RJRqmPX46cQ+jEh11I
KfuT9zm7YhFPCdzQiW/rmJFAds2Nh+RrhD2G2bEO+OG2U+mBw6JZkf2mpeCTrxqW
+q9CKxW1CNvQOWJpswBUVAggCtfiX4qKAsWzla9rXNDCQiGKJSoD+h5PXCd27xoj
9ijteOK6tNgOKhb6W9ejbWmhBXc9AZUH2Z+wEoEeqvGiT7x5sjGDQ+GlkEJC3VUM
1u1nBBqP7h7tvjKRXm+Rl0nSHBgCQcS6sv0K/ADrQ+Mga5JDm5dqGNGKRNH7sp/X
CfIGz40fyEsuk/HH6XQKPhfCRoDpBaJQqVi38QBEVUtaDcw776FyDIljtiPBhT/b
nvEKxrjmQ6IcuoUoOdKNAfJKk+5EKxVKx0TJVU/iMGNL0scSz653NLzlMJhwHTMg
8Q1iLOcPvNnkjp4JKC4Vd6m330zM9eYrYNuQoTck0TInG8wIRR91sSjsDhzwpZiP
xlYNUrs0Gb5YHoWPqDlYRo2ESGqODrngkmiBMeoVMuqzVh3lIOaVhwIhM+FbTmju
zcOEKZrdL7d+kALIRwpH1QL8XBWZsiMZjQhq+CHbLeI4ueIvOa0c6ZVX4HQulSK6
1g6Xzrwwt14JdXoo3lRI0vQS2EinenrqAA8CNmSWwU6eutFrtvOeheXRGcTaCJyk
lr7UZnW3n2uhlPGh9Ir+ktrr8YGvcstb2yr8KG+QWYKIcqWR0jSiEPPXtqjSICDR
J+7NztspsmwaeN+o4dBKUvWkNqNM5MpaSNonRA6EJCmWz6ZEVFaaH0poRGxZszWm
e2q4gsNGn4HfMRHMgEeEoSkJaVGU1mroVW8JzvL5cmOI7rxy35Yd38LcuahyY6Bm
qCaN15K3abLJIc6uBvAnYP+l1QbvyJQ82tXr4Nov7atxslJNdMtwNqRzjJ2cBay5
K5/znXn1ybeXm+2q13NmGR82heCGNnVZdd1jgEZrE3NPvRttSb9g4DyI/J/F5KPT
aaNdBs3J23yrgbVhcynzH+i9QnDVP5yc3FXer0tli9tiTE5V3ynIdoqsKGi7iULv
JRyKnaxHBIJ2lnKcL2BB4mflny6JUoSqzR549tIXOZoICc0AQfsyK8n98o2G5ozH
rrnbTLIajoogXc+0xiM6nloELDmkadjLYliXC752qtoKw/U/0+v6jreRdWQCeanT
+2pvYqAN5gGER5n+Hhgs22ELgmKlIKkOyrh1ljGsU5W14qeeti2wEMhzeQBNr1Vl
Yhwsm9F4C7++KZtbCoSi4qxJYNLukmJrNT22h98bPA7FqG28j+8vJKDRmyFjd8hS
+n9gp1lz+6G9ki5jLf2xDGit2QIWbGGq8DqJYk7KbhGYilxT663iTCUriWnhWv/V
CUL09pGZWexEd2FV4uBslVqo6o4zc0tgFvIR1WsdEDyhLDpv6keiPK/APTVh3umA
CAWsj7RtlV8TTcm45FEbsmHmxAJtJqm6nvn/BjP1GhUjgAVQZcX02O+cIOGCvyc5
3ri936+B2knas6+7ig9sTpTDqDbY8KsiZVrGQBB5YBe701QEOLjeoChwIY/H32ei
qo6pxY8e5uAp+lm44MjHadCo6G8Be4VZ0Pn3mhmqu54yRccFHNeaXQNyEwU4V3VZ
j6YXq3nBgQGu6lCUAXHYwlBYgSJBhJ3DNCkH+yMd1PMNjHSMpq8x/pawrfMroM2w
R+CFYcqUrfd7OYFMdSK4LaKVw8TFH0lGL76HU6mZCxZkP8V4nZjcPSPh3NJQ0V9Z
bPFLLklfDalNTizeOGFoHdD/kB8dGJWP2Sby4ME1dOggvNNglqdPqFdTDJdWpnRs
2Dx4g6hVELwjDxn0+iT5riewGL1eHm7JI+z2NnxxEu706tDLy+L1ZnkzsUkqHiNh
pu3yWlfLfD+1mlpGvqj5MRm/OZFiIre49H47jJ4fpawHs4yKLmxvtbzW11d2jBPH
kfYPA8qR5bPq9eVLmJecj17J2q6fy4/GX7k7FTIE0YlighaatobNcC61037/Pmce
cEcogW1QQJbunBRsSXDobxbN4WvEGqJFXUM+pFLNg0RjIfQnAR4lme0P+F/7iFh7
Pk2p+7vUVE/wsyupeYlx7+KNooPn6HAObDRMHIhCEtuHidPeZHGsAQAgVy7XPxWx
5EsljNON4ARYZtwFIG2ao18Aru1JvfENuYPwuXTUODgIn2Lcda+TQ3RWLIDIEmgi
BZCBNvydbGhaDwDCCZmDl4DDL+PTfkuU1StPhJZOLfO/YHj94Wt8dKAxc9oigANJ
3+NI4eEhOX8GRHFmz5enw7QMkSKSX0V18+hQosZL2+poMw/Uwy2OG4+J/0qRYHo0
YBafrbFCgoa8dkusngcehgE63KasmYJozZ39AHjwn6N2j9LdAjji6LHoDWq+5usQ
aRo4efeZLCmwxll1z9o3AGnX1HHgZbRt6Kuyw05ehpQLW/x2phAeeAgLeB3Jyiuo
FUbeqNBxbXKEAJYraa+h6JKsT3p6Ugs2AGnWoMAY6qnmDvpnaWNu6SQ90l0woG8x
J7FHks37qf9nLj/keyfkZp57MyYmP77WqLFTCU4HVTv1LxUpNmj9c7aPw/0A3i4a
asgpcmcUXg+AgjBoXEXv6pJcJfPjLP409T2nUYTrlQnhGbV6RTw5OqgcOd0+4qT9
9IIcS6Eb5hsgOpWVsqK6bVM3M2CbgSdRpiKM0aH9CXsXq8qB+LemEaxT4UQajDjs
vfhwt8J+ZWB1xU2fpASBDyKgcStQ9tvyTxh0PG1+557STRFSlvyh+BDXb71rPj2M
sDxAFMSEX6TVx5P50XdnU55TbK/5Hto8WBGZc/8O+HTWd6dfMBa8xmg8pFFfI4k/
Ar9fUpK2vJyYnlKmAlzCSxqaNAe6/Tkj8Jerr/lhnVyTVg/cKwkJMgjuCJ6MKcuW
L/m8+/1mnW416CZHcXVqeqNTIOQ1TZsj/a0ebQIxMwLfFdspUHeVDr6F2WBReMEj
pecEF94U7DPygkS9HBsYSR+qJIKa/TiYwXMxuzatG97nhOMe1wsy/UNutg9+Y9y5
cGZk/GOTIfrmM0/NhMgTqHo/dhAnHDZffgdfImcsBX1di4H9BQD/QHVV1LZDXyn4
PxkwjJqebh+giPE1mXIxl2EncCYDimYuE2eE6XkneJrjv1fibgy5FW1uu1uyfQ/w
5xOkzhJVlspM1kUVuDI/dPy8yX3HqP2i697VAZYi4pgIF711Ho+QNC5UawDbTDBU
J8g+HCHZT3YCnEJB9um2jWoj8CKrUpXcXP4a8iizS52iZOATWvEaRxPth2Tqsrmc
PwLlY3WtW9USf+bGXsz0AoZZjolE6wH0UlLUFjIIft7BceJvNMNbfc0aRN1KdKZm
4ephWt/RZzCI7BUSWgaNd2/XqVrySNGjRTNrFbdiXGqgLJTbI7IcZk7ATJZxnzIi
KoY6DXkAhdaWwWJ/A//NN/Pkw5LCsgI7qcUvV1p5b44MYqfjZayQiKdhC9nABsDr
gWZ2oVbkUrWLoVm4XmM/71hGgf4E7bMh6tWDBjSYD6ReUhZtrrPgAAO9T6XVeA6u
eggvMZxOHpvlgNlDnH+oCa9ir94b+dcMmJK92eQicptGWz/Uqa7TsXS4NAXG9v8E
AU5Nq6b1YmHrzJyA5Nd8cJiSfLlnYiJXdbAOFH6fGpwDMm6huWPjG4lKQlCDHh9U
kEGmMGQDxE5HNwA+pOImOUQWFG0KWwa69e9kYkcLVCbNgLpmqgpmI6joh5g02cvo
cXgJ2VJCCyeES/eIQlhMkoAR3f4KA2V/Qbm9RgS0AGDWw3GEnps+2NYyQrT9kbJY
acYO55ECKOohLNK0lTjSL+ukBWP18XkNI+go0wJyBMsHIhr4lvNmXiUKbE1fZzCx
32h6IPp0SgVn1frZ1JZfe+n0bTIxDquoITCo6NfIZ69UdMi6kyF+CvFG7FrQRYRV
C0HmidNO3jWVOuOUBLKXpwPIQNy3OuE3Rsi0H7QuJeRhgNPSa03/KhgjG8iFGioP
lws1T4VwJ+crOSksChif550aNnfYHn5R98gObTyXJvyw/+jeY4r3rhfHZ0ji/quA
QbAoiv6+Ny6ZA/FhCVulnW7VL610tIp03MOChym05i/MxzT8CF47KUSF+4GhwTIH
/k7xqzVleeZKIuHajWdpFlBuF79meXwbcI/zEdMspXlFKF57o7lEuFn9ETpVq52J
wWm2KZdTSl6Lgcadsb2jxJUv6bv159T0lUPCRbKmD3KhnJLxWr90rwI+qUh4kJH4
uBW/BFq5vvRWCx5oQg/MhKGQ8Z0VkMmV/BDID/3Lck9fHLzlhA2FUcM+YscWVWpy
hu5QE/JNeLlMlspaGC35OQnXYtjxwIHDJqeRAnxdwBrUI+YnaxgJcxmZvTzPj/5T
Kc5n45hZCTeFNp0zIt3zXUByyKIQqFrP/DDwJciDfOknfSWeNkm3vKpedk8ZFMKN
VRymPj9GF2sG5J7sjRIZb8Ah02KtD9QjyPN0wirtAhmxol+77NGs4NvrWqQqE+RD
90EOu+GQF1LfAfnu4pwced/j+zdglma8AFEHFKCOrRCtQ3aQML8enhpWXz7tQbOM
SumZWyWLuP9ovbaUtd2CBDcZpmqCr6LYR0yoFu8oPp64uBytqCjYvNIZ89rUhkU/
kBQxelOZwg6qGkXo2ytCvcYvlJ2nrBgdim4cMX4OF1/O+BIpddhm50RnAn7Cub/p
SQ9TMRTOlTDk6ce+Kg4US3bJoqSulvfiKpo4xSheVqGiNmMhVQIDVQwbzFuyyyex
Lad0ceqRmrZmOaku96Qxcv5TCHM59boXH+2Bd2VRvPkRHiKYgKH35tOO7yILalkn
Ea0FVm2LiGqt2mjl82BpPI8ANg/bNGOwmfRqwP+eiarM8BX6tJ3fLWCB30sTSOyz
wB93DXMPYDMkyzspZrooBNMVKLhHVszmMS6GRjOFKcwhNgV7fi7kYDVWSFsLutW+
qlP0soptIjqRx+9sD+QT1v+nxQ9T5qZbLy6rfU2K/bt/+c9+SUCc0NKDZKIho41B
l1L+8xxgGxbx5nKpEv3bqdCop6tQuwd3VZsd3Mzs8HeLLGu+0Lc0d+pYRKKkSLWw
QN5pTU56ubRAVlmbW16w1QSaBzq612UaZrjJf5y+Jo/YayWBMzgpP2ef2qkX01J/
6j6hhZqb7RqEJSRW6+rG1y3xttTRch5Yq3FF+HvstDgP5pK83eV1iEb+29v3wRt3
F4mR336eabeupt6FbDrAXVV3HDJGkToecmnRvL76hE2HK2BDsn1/5qRuWcnWLopG
H2J5gqLHAJysnbeSWxQvc3QpHH0nxhwtkAOHnBymc70YMpQdTCbpXbGwS7GU6iaj
iLF9MEfcXPaTGon6zZeNEtPkQCZ5+xIFxHWzkK5uP0U64h3VgPE/KDHhdLlZHLgu
dZQpX8nAvzDuWudYCXHMQC3+oG9YKi8V1nUYtLRQg+O3ugMHRFTyMaNJ6l7RmTmC
0TVnrrgVvz9qH5AC3RyQrdiDPJbHvS7IRkPVCQHXhJm9ietySDqyGlK+v++SIYWE
CT71lOqRuaEyV3TIJYM7r2hghBMwjqM+ZVH8K9oyfvlwhCw7WTIhLDFg2BgUgc2l
OEKPKd8LPmjI7JE8fdrufE2zwiz8QFMi5vBPyr5BuKDp73rtjQXf2qbBRQr+6/Ju
i8hMNjp2OYCRzbZxBIC5nkRLRrWASsotCs8/aKXYzZT+tR3t5JAT962xYi0hkMun
SwDD6W1c9WG0oT2HXm0sV330K/QlKWVwVkizKDJJGKZv75RZC8fBOjlYK2JbcBX1
lLjVKJYYw08KC6mTc0CsAMzLvMdCOQNM64BSO0tRoPegX69iqWKcAbFHYeXxwNnk
BbCTgWUA2Z0imU8y7GRA7C1FDcHtX3jDRC4B7qEFObflumvc2S39K0px81WX+Aue
y1Hk3S542X25PDLSoHKvddGX7/y5wPW2VydBp+ytHMUqNXbYMrwNVn2t42P0mmTW
rJvahrW/pRvV7D8MjXCDu2WKRpg8XX2cZbNhAwlLrBTBAW/Z3jZ1+WobM9KlvA7A
ozpQB6s4SRA93JB3BT3C7bXtCrgrN7ayw5qld+7RPxZiFlbSEEACU/XFvooVdv+/
XqqYc5YnTvQgczmKWl4bKiXvmLTZzHzYwEFY/0QQM8Ba/XtqmYZK/PtMhM4zIg30
I4n6ZEPj4Nvkpqw5i/iG6i/kizE7ay/A5AcLAfbM4hdOwpIs9stPNqSdcnvHDp1u
mJH9c9ESUE4JN+m33dL7qIuEhhmS/MM+2mE9fyClO9LV6EKaKzgink/iuf9PReTl
DI4ytO/rJwLjxuI72od5i6o2i601q1UDeX7okIphWb0NQfghFiwzBkNJrqf1UdaN
JBa+heH2MmQq1/A0ZTdd4p+6PKDHIQs5UQE0cFQk5EL2+gczipcBBv7vWztMm+TX
nAAqGOMTJASLdkb0luqnNRYIYAXfVSjketkRGTexv06EHejs7G5Iyvhm9ElOfpTs
Dj8YdlXDz4obHq2ApN5t6ZVH1o9om5P2yQoPb9OjMboNji90jc6MyqSrxOndlfrE
+B2WAvoFGg4KZIzPQLSg67f2ISmw4FKfBElaQj7AI+Dmxi4lLXo6xg7PRGiNvv2I
VzC/1iJAa0Je4Oa3JTJWhph+mINm5kv/gIV5UJkcqCJwCjOyii429MO44h+QbrTq
44mOqcU9548O8mcymdyeLzpafSyoeFIjFHorfaUzUd/yQtcqOJSi+2naqL/TFiP8
eK9bSkJ5aNesnKCisJfbYXcGhA2lGIv9N1Fy9ZGg0E1ND11h2ZrZJi03Nl/utv1o
Ymlo1MFF50dTuJRHimVT+3GFGBp1y7TP3FzWJcd9J1FqPbY2u7hK6Dno1NQP4gjZ
x8eWQNcReglIlmtKEUp5OHmatQ1TdO81h8CIDdlkcKovZsQ26nT23pMoYlm5N9lq
UXEpzU/ijgNWdf2vK/OHue8UnncZrK+31D8b7IZv/Uz1BMKT2hUXQTJXwyakstDE
LQE3Oj4oz9g8NL7Qk6XcJaD0UbOJ5F/iv5cI21LW83WwmQmgNA+WH+ZwgNfo26wf
u9TROig+jufahau6/e4gz3nRa7TA2FwSB87lLBFdv5XKE5mVHZMJjlLWiyZKljIT
YtjpP/1KsRm/SgjmAaiyVnOgRNURgcNznPqFrxNIlXyRBNWhNzz8C0b001POrrmC
diJRAj2QsOLz/sJ+NtsXw8qb+X8+51lVe+n9ZsWXOOMrNA1mLPMbhsZYYbYD5Mbv
DHjmpLPqzPPk49aVaJtUhpPkXpFUks0gwhTDYHPvZa6VOEJ+CogA8u/gjO5JtLMc
lpBzQjx3JLvsMAE98muREZTwrHE2bL2EBrj+URFse/QcXgCSAMxCmqsfsUxzs75S
b0aUxaDM/k4xr/Ag17pVYv9zHHmWUKaABMTl0P7niatt3mptAxYV9U4YT/w5hk/X
5Vn3J9aXcVKAZYp1fmds/5R3iwBB8dpc5LfrrgBqcefYXTyUae9T3ucA3rmgMKvZ
OmCzJnq4kKB/TpgmgUJdTpS9KUb89QMdAuhrbeJXebIg26LAjuHV2KaculWivtJJ
yIRF03+9L7fRXaUYxQ48Xx3dOop7xdoExtdn3l+ptyFDVPURVIuFSWzAP8Ta1sCS
Urg0+od1zuZCHL0M4TXdXJ+8zXFRyuNqbd3dIVyDoUYxekOsww7FWgoJN9+MNaAY
/SBdMCjej6v2PidAp4f2pzCIBbNhUMNxTNhXHj9r3vBXXR+93o6NteYb/Oh68bU9
q4fhl9uI1q/CEjr5erHEYvyvKPrmqsFMIghquIUvPVNQOy+TWVTuErFw+xxWqdxe
ljEgSfyc2nNIvZcuUt+kKIZE0D48xuh4WoLiQ71VqphCibqtF5L47l7T4DFYMMAH
NHZPhDylbbH8lMzfmF28c2jkl8d5Yrlp5jN+8AiR9Ik20kXYD5gYNDZ+1+jI3A9A
KjWWTwCPNvh2IvoJ948tS0V2m1D0Sws1ZAq3CcY5Saq8WJv6RfX+U8S5TFQYLK3S
nJHjOqBjUy5J8bSkIob2wJ5mfGQNvXRwcW0Z2eecoE/l8d1ayB/slTTx9eLCs9YA
H779P/2VUHJ0bLdKDs/2vkhgFUo4ISSuVEaBDJUgJioXL3AhKVU7xCL9mPO3k0sN
n7+JkQAQ1jjRuRWrfyuK4bTwvw1T0unWwepzo3WR2FZvee+cLpZw3hZ/ZdJ0mzIv
Xbfj7pqGscq/h/GsFl5FMPZLatX5y9MoYwVR/8jtEVIlylxNln63/x6Bnt4leRig
1ZkWeNsmvu0yZNPXQLDJzSyi2aA2iKXrCY04AalKcyEAypFRd2/RqvNt0vkdFjME
teqB1CYCE0Z4YpTPkXApwXRKRgb7raFpek85DW3dJKuWrxdWE37rUQYKflaYClrB
BAe4qf+2R07G7rTvKJN2pc3uFkEn05WTDQjx8v/MrjXsv02Dqc6DT5p92EyNz6aq
FuTyYpTI3+ZQca33yA/KVPA7Qn6qKzprJEQ2djwrOEhKx3a8omEGBL9BwaM3xVgq
Ydf3b6XG8PQrJJkW5h1/+NjV3tLDyLVSXgV/SztffHTFk6yQSc2B9FJHl4kO7NqG
0ILiZMguuif1C1PC4RyAkxppdyt2wRZWbGIwXoT75ADUKwcnXagDQ2N4Qw8M7czb
cm4FFQImIUev9LzFIFiT3Tre4FMey1uxMj3MTTIMgNjaOkAmCwW5q1Z9VPdihErG
cGqBZ+EkKkLt0cox8ousPikYvuBm2t2OaUuRl/O/CTgqEfeZeZQUveSRPjy+gJoZ
X8MmjZ8GPMDzg3Lj7W3O3t1qazv0eso5ZJNDst7yfaz7J5kL9ZJO42egrzuWtMdC
3X7nNXNQppLD875DVkwlwAT7vnV87w3xvfh8CuvwtQlHmwxaavYxXcWfwdNLKS3m
5NImzUnbsk0YgHNIcJW8gjA3881YIKstXTSBHH2NG+U/Zgzifj3KWRTgcME3JCZI
kZoGMSurvnLtJGSeeS55oZOx9JI4XD43W6kWlHabkjFjezT8NL0sNXJWC3x2dI5d
emzmQ/oBScxEuIZo32qba/7eeSb08DD8a5EtxETOYws/luo7E+cSq+wtAAyieUcu
fPE5lW0gTd8TmmeWNm7s9Z6u+k3mIyWanv4YTKA32uK87iW+I9iI3LyHm1D5Hh4E
vP2j0fXvDUb4SCkn5/ELdEQO2mBwcQya4dg+5X0QtrDwYma4ssaAqZrAYLa8v+7V
6ELclR/SbQlCUad+ce30CvUPIpS4SO8V+TLx9ncb25aexomo+xr2LIck9IIfPkCG
LukkXYc2Sngo0NfCsdMhp+oZrJKOGd8uxrY7P6eI0UvVH0NBTKMNU+e8Dhd7g8dI
JVsrKBcLpulpt3J1RlD8Ah2nYRKFV0Yiyw3S4+9CURUxAREE/s2IQT6ujLcrjyMn
oyBprlAU3jJ6T2DLLj7eLKq+DdZmHZ0xjqvxWKM//j99yMIohwzlqK6T4kUpJQMX
TT7BlNPmjzP/HPw4Nl6pmhUlSUR2slRrmH2Dhsxt72Ajq1fbSXcPKtQAsVPW94Jc
j51/na3Uwwv0eo/s6/+Vem6WlMJP6m+dvNw4pnaAkcP7/6IGdkmviSP/tW1fIU3i
g4wOUSn6ghIkIkIpBfccq2QGtc+tGh5hP/joZoxBDj+YgyvfGD8zaa6weVH13k+2
zLbIyZse/WTQ6Chg6nT34pfZUUWUi3iVmSKgu3igkmbUOe+NcT+4yz0JDTDj5muq
hLZypz21DVNODWolUPea9wzeO53G0ayc+lGg3cVGT+eQsBxgdvmero7f3gfNcEnn
bVzWIY8YdOCo1dXXx4REYwRWgQQs0WX8MIrwmaL5o1RhCzMeY+FFD66pXP47Fc/M
stYfcAU8rl6oc50YXqaicZ7OcmkCTJnqHRQheP0mxUTMpdsQ9pA6/Y0o2QjWTPLo
uvt00rbw+dNYhX6xWbHGb2l4JwbYgvt5dqdbLLIu3T2+4xqwy/DXXl9icd9+KSFh
1ttyIvibYKPF4cRmZkkcUl3PcgwAVQyrO5pAf8NGOG9XUvtottLz/2ukV7gf3rzQ
xPYfW7ACA/3NH9BJGLne+picoZBZRLC8sXJrAZ08zPVVu+rLqylc4ku3ORPPWWjY
fpJVwFzHFMH6kywYQyK8up2pmtBIYEAWJaawkHVNml1ALXY7nvKFuOnW2NySFQjl
I0WN1SZhlHCT9GwtK4vXp7ATXhPHSJ8msLZmoDZN6WQSu3a5rms5+n5fZK6Ahe7v
SkMGrafJNZbsgUOcwmISGBbScq8kKZBq+IUW6PB4x7m8EkDIdOGy3t7xuwgPk7aI
Edhctfv9k3GJljx1UYvd/SF6l75OBuaCQkFToUf8gjaB3/IkK1bRhbeaSQOvp3XF
AgYeV9EsRsELzKx5+3bFZhfZHa99+6OAYw6azu91kk+YECj1PabbWoaDLi9RAhfD
utp9cK+dpCT93LY9rD2yDfTgvoKeMjLrxN1XgU1hosger0fFxq3Y98SqhZ1Ha8ew
OEKR3sXHpDT1G3NIykw4axVBiS5Nsd1Mk5BP+cXhOStYslVl/Hk5hfrjjefLsNBf
HTwjx/EUucCIQy2qM4qo+eYZmh5sEsrtJWvXB8i9GBGNUf0TrWmVNMxdgNTJRBjH
8ZSytWW7M50BBkGN2BrsoXu3HRUiisHBgg+N3Bu9VeYXH3z3V158qgNiQEAggXic
riVuDJ2oChdLe0pRodyjGFo7cI8OFDMQJLUzxWkj/UahybQBHEk7HlSjqUsaFQYX
xCP//dVxkxmpF06v1jMd/3OtRzsPs2BgR6qKm4bQspY01k1C1OJ8b9JcszYk0BfJ
bwAPhkq0BDZ5NnvnqqwpKdI8xNTgE0/BUuZM0Pp4AXWVCa1uuLxLv14EndAbN/wn
lYrid83aMr7mF6J1c+E1knuRVAdKb29m6+8h9dSLCCGbSv0bi20LCKNd2JKGlxxK
RxJDliaYZpBOdYaCs33vB/aBNV4jTE2cneyz9nJ/7KHVKbBfikNQnjmM3doPaMP6
gUscD8aiNI7eXePcnrzGqHVLsNoYMeCD5e5FgyTlJ179bd7b8p0CH15eOgTs414n
uoFEFThewZrT/COVaR5D+eh41ypKVsQ6vt11PoS03Ow+KBVkV7PHD+9liT2XmbhI
q9RZIVu23YoB4+yriuKMuZ9idQ13qXMW7fAkr6YrBHMwUlnOMv4Z5dbiHzeeybrc
LBqS5BLRjCvWkD+8ZL1BFBjm5socy8qPNwaml6BYs6qeRU4hu2NudIM3jcJerP4R
XY4QUznZoZLF+bg4PwLwCzfj+7ECJ6cB3B7VHv4RnQYvfIaokLOo8J+43+voc4w3
Jc6ysKP+RvJlD2xBqcsrkjJYKZb/0jtpL3NLc5uONcxrLopmBegraiBS0xeHUxua
35GLedYX1vyZVpu1UxovndcLdG4Q9vghzjUmGv53uKQr7dmzXcQcnd/73qSjxTQD
bn9ZX49QFg41d5dvFvM4KD+PeQWiHwKn/F07kKkTlo551UZSOd2EgHZ5Ce3QiBOo
6T/XHMaYKOc+ct3+ZyfctLScON6LC8jU0RnSZj6XnjC3+Kjhwcs/Bu5YUO7CanYH
VSrvdGTuZz4VhquErTSlwmPA6fFJ3x/eEh/to57nzdvCvLY37SbC9A3vFZkrLVfh
9xc9bdAZUQ3wPQ/dwhjgXA9m0M5Id4r81HiFHBFK/Q+nrjfkuZcOJXxxrp5CJuZ1
H4lJemaJVoZZiLr8fKRzEL7dBcnYB+rEMgk07cCNdgiKI5q11mLaVTpHvrMOnVYK
Uoz5nmo4HaROA+X+z9ImQFedy0/eRGKW8uIQSYq0mevrRPC0UHkV+DIBUMzicB0s
6C/vgxVMgloeSOJJwV87C7jdcuxNLmGD00dEPOxopayLJc0J4OPg5kAIKUOwu3as
g3y7W2jkHzr1sm3+tQQQvsYkm7kdsAswbuOVzwmzWMtt6Xxtwd++xwHuHAUIodxd
o0Gdf95tBzN+B1eqkbMEH7tRoQ8x4u1PE+0kQ+fDzqqIxRFpIe1/qn6pD5J9XaZB
qboHmbJueU84/jYSoHHMYavw3BZhdX5DFb2PV+GPK9sfmxH4m2PuoB6HPhS3ikfx
XEGf5VA4cBfozERaIj0carw1xGgUqxjvwxSLclsY3yZTo/uHGFzE16t5knH2YRzl
Lgdu3rGdgPguoVbxcXmyTXuvVLJxapbuJPPKqiQ0LsxgSg9/EZxExutG7Zm7bbqb
IZqopd7v3yqauOBrXxeogASqKBtMHGnaChS3eoNB2Ub6xvkT1vs9TsPmthrhhcG4
hymoii7JfT0xgwOlAi9Ox8Vik0LWxNh+KHGA5L1arr2WEMuUe4Yk5iVKGsqmTnfu
8TtRzFfBjocrWrpfVjzaARHOWog0thRTb9WMEzIG/v0+i00N8avfmEQg8qwx8zyB
lW0aVJWINseciwYen2/1CoaUF7WBebI7RoveqpQxI4n+vDI4A572jKdlmQ/bCZRD
D8P8T9QVDIHBK1xITnln8I6vpEHDsg7lxzqBO8RgJY+aaKYC/V0QgwqxRR59NytR
9mbwQrFG65eLs3jPmR7tsHDmRFlu3LCib8PlYTk31Eob35umyJpDEqOe1pzg8z68
FEYXMNMbM4dk2wbnnCfuxQIDA3CcaXot20Y6RJ2wTUmklEB64kHHr9AZNLHada7P
sqoSNsAuXqmPlhoMyQD09PkVXlnBfLdp7SVulizi+th+/C6s3GoGqqlZs9Vr/n8h
B+J+noU4FaYe5sklZxuUIh0QqTtwgjh6REYAfe9gG7y+fHFVd5nNPrem3qYBs23d
1oazKCA9u5q8XPG//0o1J72TabYq2ZDUJZfAnO7WXtpqau/U4Z1LlJpPMOQeXRkM
7vFt4D2U5y0v7tpn42x4f5ym10HUGwiz+edOm6bfcftLewbLCIhaL4nIw3IM51r9
+OpFUSp8DYh9YXJ8DybWcfAL/Z6Td5LA8d1qNv77W8DFndItm1Dv6oi5ZgHB4UaT
3gOL23saYA++TGa0VgegqROeQM0skOG0G0xvNksQHyFNSj8TyANpsjXIKy2VsGP4
SNuHsZ2lFSmLXOEDzu629WoTzg2AY3LMKfnaaww2J3WW4tkvZDsfCQbXY5u47nfO
9RfNjKpKPTtIKcpjjMMv6OIJbBkiB3wradzBLnyrkdtNAYRmmvntOoMakI8NULUl
L4RfaTe+DITWIM2itfsDrwMq37iHdjvncSj0rcj1lVBVqEWwhWp8UUgSVB0H0cSY
7V5NnXgT8Vu8sw+hRTDhQEcr1USu8HFZjaQwsxppb9wxZyhQarxrUDD/C0ycYPqs
OVUxLqpa3rv5nhA3hJTrT0N5sjX7xABfyqEtCuh6wr/duXIWN0s/P8CWJLVQRwxT
b+cz62zgg6soNN/kV6X5t31WOhUxwhYAtgpwmmlJGlYNteC1Vjjj0dvfx9xoocqI
j+gv5xiDj68hAO4/+LuRvnSHESTQ66NSXQOv3f9IyrQgjoPZWzgEZz979tTkRl+r
JAD+v1uwbwr30qxEGz3tj75wKznShhBogOizemLBYnXzyidKnV+E27VREzuiZBrC
yuuR0iVTf2fcezDvMdmzgHQm0eTkhffJ0mGHnovBZ+CF+3dGWXkAxeb21Clj0ZeP
ZpwD+YHuDgPk+m6ZM0B+Vg2Ab+9PTE9THS3mQFsGE/XAFHCKC+Xvzflhn9XdoE2D
HHhiTIcOJC7TzDi+NzgBkR2H7iVdkoMaKnYzh8rnEkvft8ZZX4JeR1QyNvif9y+c
LZUigJoImLzPcyx7Bk4erGBbBQ/U0P1cEf9LAGFBXB3jYT2WrAUg+r8exfd2EUsU
9jbvG1C5LdmhnriZLvF3E3yA6aOzyBMPd2pVK/NtC6vH8r0klsnbgd6vssU7jZ2K
ivoxUjyukMalTZeLuAadNnFevoPoa8OHiF4UlAbFlCkeGy7Oz/cAZXS/jDuxoItd
4EMsXYpPDH8PaDuhh/Apxjro1kC1LJ0Re3ISGh8gxLoKCB51UxzzCF0ZO0zS3GRW
LopfrM0b2MwCuyywhPRzYtwHgSp+aMyrSGqFUpcjUOkGQMOzvjbQW0AlxRBay/vM
t/e023Wmxe1F8tuhHf1bRHhNAODk+Y92XhkBwcjITWQwFCUKmecGui9mLbpSOc4Q
8yqP7X2UcFtPz/v43kZCBqx2iIXH8WVdpx5kgT4D9m9K4IiALOH3YlqccX1Pr1jA
1SZVr25+bolocdBP+VLP2EvgUZs7K07Z5zOCEKa6c//oEZEYCc5qMmHppkt4ZPuW
Wmur01hqWE4LqZX6uU05dQrKVzlBtU5tQSQ/PblagVmWU6fY+UVOfidGX+jTLQtV
2ptnvkpJ6oSoPj5WH2oZDzn3RvMPwqFJZ8585RBZCM5xRBVTJqaeByDpwRMKOGpl
pI10nArZTp2VQU+JCdqFIrSMASd+IpCDJWb/TxaXgDNE/daYMmcVflDSnU0o8zFL
8ht+Y663ss2UrnJTY5+2s6++GAc1LDXby+GqYgiEUhiF5sr2IGa/TNqVlLNYSg3m
38CgmMYxRCDSKYU9DT5HsDwZYEeIHFdk1gDRhAlyeIQH2zLxeORG8dwNqm96fm2G
h7toLMKwRPy5aA2NU7S4zQKeduccaTdgNYRhrEfI4igpu/xBRpF5fvDvEmXsjERK
uxRE7E0kk+7J//8/+8Zrk42IW2We02uz3liMakXqcmqF01f/yvxWroN4OehVFu5E
Bc/Fjv5QKHH6Ma7iNkaYX12hqpRYqDWtCifuOY2ErRDX2V7cyj9tlzwY7oeFxBqV
vsE72579cYmYo/a0HIP3phnCz1daFZtieTru788gZaYAWT+njxcBzIuVT72fddih
y0GHIYewL9ms4NvNey+BEQEVfQwDp30tSB9ekK/UVhruK/0WQvZYU+b3btLihWCa
BS0CXFWQq+dPonyIaq26X17YXic3I9Q2Lw9qOmNl3q/1UKIC+0e7TimiHJZ/zZP7
jMGyUWTqP0kP5YXZHguEnBEXtFbWwDHv3ZwZbOsgzqhbwKrLmflmlAd+cWxtXcHU
E9HNA/pMFm622D3n7M+SQtsoaYci7Oqm7GyNIuYs+MYA1TrYOdKGSUzo8HC7tFyf
4tO5o8LSpkzIzNTUWrvYgCDz36+KfAtLOnQ0+1KGJgoMB4jzD70iYNfz8PtBOrMR
kSp66cZMeBDMuWJM+JKH+WxETK9AZjA54bk+V+NNUj5jTCHZODfwObQlHk4rDVkl
kytQ7oLAmd1oy9mtnCDjdlxyFScFDJskQ8p+f2DT0inB8QybZicy38knDC5CfgLN
9I7T5a2pzdCxuKNoqJyh1zCKXgwYsDzefjDwwUZwzv3IkJv0IeSe33PHDpP+rVNR
lI1AeO8epl0CaxfSlmFQZF0wkTo1cp6ZRUJJXsWIXSShRTHNoOQFg8f8TVgUOOb9
o2lFtSP32JNbTF6Zln/u5ryi/fdMRbcuUOsO4kiCY+GSvr2FvTzvLnxlqVJICrFb
bLjixrC2hB9hDkweuB92DdzLhyc76wMV4yYhlvNjUy3us9GWSJADLYlOa0AO6vtz
fBXpBCvKal50SrPi63eJ1cr11REyd5XdrQ9vNH17YeTsu0S++gdIdTzK0QgmpX0j
Tg1qRAfWqXj7mihvC0QGOHr3LycllPvTGE62x95fBIrbKc1nyYRWWDh1aWm3uSmA
vxmXohVd76om5U2gKLYmICT9SzOqOhke6wrtfe6ZxPPRhUshgGjtoeOFPCMBISjv
d+Z0/ryZ0s4eXhF2A66blHyaUKPvXCnYFUxztSABKyU48sNtAHDYKb/Ut628VkwT
wSLRvjv8FPi9gHWbhGmCFeTlk+6f/yrjB1lPUv5QwkMOq35WhkEycQYBag3qLfAn
c9oaPDNKHbE1prSVKxkllAe2sAhEKdvJhVSdFLieZnNoeyPh9q+Z1DffA5OmvLxe
oLidS9qh6B767PMRgpFcVIrdXksNQAfOC7GrauRsUhEt1qIfqmgKdmCAigLJIWTD
3nViyWOxub0JL8hE9oouwRdZAPjp1o2mHNzBYdYVAbRu+SM14JN3qN/l2zv/plpv
3sp5+LugMXT3l96/Zi1wviNkF9c6G6DxLU/GPR1iQD09DksXnhJuEqAm5fKoy+NN
tcJc5Y9jLc6TYaqrtIWur1v+JLkC5U5uK0U2lmjT0I6mHkn4cEXJdDfKekwObQZz
VEzsAUH/OmfvGknG9Iw/ycLq8/NWXKMO2kOVNA5uocCBA8izwhp21Fza92pKtAp3
l+1s3yBwAQH2ZDte3oSEaN4Dk/qxZnW9VQNlDOl2RVS3/pBcVHCfMPgV5JaD8FRu
nFqJsNYJQDV6+Zs9RbFlDcwkJlS4LptwRrWdsYpZvW20SQIZQkFJ3b0fHfnOS+FP
mb9MP4B7SQedrgNMaVmIJYgvEbn0HTza22Hr5wHF/KNhN3x6Te4ky4pc8aaBByT1
C5uqd9CFC1+A65xCzCuqbGXUfD+fcOWEuXBirOXa/POqiQCG0UZCHOnlmnbqkbHI
6MJpX0Fepg3JjMl8m7Bv/tsaj/ljm64s5bKY479x5pfKrDI0shHp7nN1/Ep6jqtt
HcM6NT+DoCxPKCiPFSnyU7S6quewwzH2amXdhUtLV/muBao0QyxRxtCp8zmvrw7B
C4Hi59KUk6VdmEdM5mZ0qlNuo4Qc/9C9vAsQNKEdukxqmUQnKFctpWZzvG5t7Zj2
LhByTFOf4VRkfPhrppyCf0Unz7iQeSQB9n/Zv1aUkxjSGnfafkxkwAumtSgHrYXB
Hm5X11JmjtcBvHFLr81JMjUxOxc4Ey879sLwLu3jEE/QBNEnfXfuj1EvbZpSHw+F
PviSMsRveQxtQgqAALq8Nln6I8VIu9TyZYo28lZv15Ne6Qwn6E8+UBuAoctwMqaw
DWLTYaLnu8Ee4Ary0pn8W3SFGP7E5QW1WsEupoWXZGIz4bmv/71Ux3KMSaexfI39
hq4w9TR8wTmvNYxPQehvsV+pEMnoNLNSH0Ie5HSBBAoVBrW6hsbn/wcwKerOBNhs
8isWiNL1CNOm6+EHgHXpGTs3R8g1FM78J4uHLE/Em9Q6pztyJo9U9PtTIHfc86Kw
TF5wba/FbtFU3vmGGFXnDySBEmEoia1RZQCZAYhbDUDgxjgGoT5hV+G+Avs+cGpn
FjpasCx1YlPpJXtT1e50TT/lYO1+MXKTDfhdq2D5NWsQsfKAAKFM/vJfqiYpfeMD
xItkIIUWJqcXXblB2p9lx6Zd/G3Ok0kI1bkTX1Nkdsle+BExCtvSnDZDnnjP71hJ
2OH9/FMwgWhsRk5WW8tv+QTyEJbwFQ8ho4Dxk5fmVmjJiz+yVXWUGNUrkRf9RBuo
I0sx2X+Uy1c3Ip6EVp5X0N7hMFBZndM9XARp+ey+HW5ILszPeFPjOkdSwIgG8Yt3
BosQyi24c+E5DRYjUSjCJtjMBLA58T5rBbfZh3uPvM3DLUtetiU21njX8/0zqLAT
49EdMjB7flcjnb+sQOf/v6jkz/OeI7dRshvDRtYFptRFMF8OkVkWe+cyysg+jvOx
a/ClqnavHZRfeRcGNBEjvnY4ooYf0V2kj+isMVCqs2IcJ6uaEBngW/AykYyMHwS1
2aqfQc++7nv4eKEbqhzWLgWHzDch46e7P9dNFqKNs9HSYUrJ3grcxjiS+hNiL3tG
1aTYGfTRnY1ZjFzwMKxJKS56MrnwazPfqIpdj0veTY4bXBWpEiEPxxYkT/rg76h8
NsHDs8LZPVj62lAxqreWTT6HW7votx2G4pMQLWnNvX7hgYeXJZyekxUz1PAWsES8
gslYMfnOEbGppEUaDU+sfIdL4dhNA5kI/3XI9tTAE2yR2Ggcy+ADqN6RrpDUkc3P
4jm6xj3o7ASFqb+0LlcLyLB468jAELQoGgRWwxwwMef3l5R/HVqTFQIab8+B8X+v
ACNI9feeObU1ryl82hlUsLBAvzGj01cNLTxD+IjWylJUyxXARV49Jy7nBwouuFQ2
s9v1PvRFHjmjeaIYk3HiX6XIR4Tspp8Gs3leKkV46JUlm3BlEAs4RVN027Shtnue
NvrOrYVgx6H7mdISJKEfQFVjf2TEUPUPDu3009loD9Ay2jMKUOKm2MrYglkR2H0W
3rZVA43ci/zltUFDAsjzjaIAlyYtEtHMeBVDNktShb8q07U1rsn24Kq6v+9lK+xq
P/JqzntVpRMKHNvUCJ46Rf28qawaKYBrhjV7qoulRNy+hnGt4YtWHmMMhjhF9xns
RZwAagiso+GJJH+8LFWKcGavgIwAtCZxuoUiHAT2LYkSacWAi2KGRN7PaZlPr553
9Pn2EgNC+X/gvDfcKK/+GmjfOQwdQFhUdBkoYn2GjnYgT2J6PLW4kW1Dk0swAsXt
+wIwmTwPmrJHO5UcmZDKVIzxy7Ia3mApUHur6BetvTV8MPs7W0Y4i1zlQ5sFbKev
IriHLmwKsoHgIdMzH9ki8BAPcRjM3YVoUfKN8ENKQOhHJRpXM6EcM4GKkp2svZbU
V6pkFRrff7jpjxFLB4aYivi5kkll7Fc1ap3RrsfgddGd8T6fI8T4yiFeVcJVQtMu
WRF51J1p8/JsgQjd2+HufsexHtr/QttSCqG0a6UYTqcYZlxI+B0o6eAFipaa57zE
+7sP5d5yMv0nPbkUmKlMK/At1d/ZnvRfaJxCKzeleUvzvcPTmja8XHf9a74n2gyA
oHZJoXp1kdxZFDmBXgCsU7enyJX93K0XM1yrfjMSrKnS8uhh7KQvgmRRWV4CWgLG
rEUgqSyHTPqgaJKgUfx76nBz8OvOzJ5oFeUPwBYn64KKl47YmPr9OEYztNUlJ/7p
OPtBqtUl5A9hH0i0bkSbL3su5ydHeq7ue6vcTNkij+xmlUOEI3ExmHN72zdeIHtf
oaq/uijgrhFzy+oHPJ7PYYL99Z7CBvLI+TSXnHh0SvS1jl5mL5MYvJt5Wd75uRs7
356g2eeO7cJK5ySM4DO8OP6VLTn1CdzKL2wx8OIhXklJvZMq9qkC3Jb1FDYTa57m
jsnanQQnnBw+t2cvYRiOYk5NA2ezuV032G5z5v30CAKaOxjpRHF+8iojKWI9ErQS
7zTUEoVm3qyz9ZhJzbSEI9XwqUD4bnx3g5Ozka7wJN2tURKoE9aQtXWRv31QWfJM
jsyullt6LCh91QlEgTvirxoiT/8TKSab3JVSS5k1nDqEAtDvoDgooLBcvIV/AivN
kFMCHhY464qGz69PjewTa0C4QkNAn70MARraY/azJ5Hemr7c80144kDPL58Wwg4G
TD83i2OyHLBDrSbxc2xfoOze/Y7FqLslMnAneIsPtGVjGHALs7+r4ZrbEB9OUjcS
83fCnb6G7UhWjmVUG9ygJ/nYhnHD7igcGsj7irEt2WVHcUzJDVctDf7mwRhbAvsV
5/kiKOHYKNNlxDeHaE4ODQ7dP+araT9Wml/1/57vaRYSw3bkx6v2HifLv9HLK5L3
y3eVHK5MII0oqSicz3s2b9qbL6VPaO8hYtj8tWDKGdVw/oT+RqFzdtZwIgi/Hd3N
uk6SYbyPYZlMuHYRKsraNGv3Ts7605M6vOKkFAlkPZZp40E6FV7900o3x4L22jIx
92nr2jO5xtbH5QTSlfGDoF0jDTT5sS+EXy9xM2sV2elopGl2eU1+JGLoZPrAIF1C
su/XGULQFGfsTvGbPMCN1LQbEFIenKHTG/kDJkeSW998iXB/8zISVoG/GjK5ZV3i
x5tJ5Z9P/bs8N4Tji4X3gcY4im0F2tBP6V3uvECVuVoOCvgf6YV1MMTy5ZFNYtgR
xRWMhX8xsW/lNbTbTsXH4w+3gUdtKOY8zR4iTCxp0GqoaX1xU7Jvp4NsWD4pZMr3
ugsZ6Wc7hOBRfEZAQ6fIBcjKZAYVFJ5+qWZ2ehys2ynCxaGaNRy8k0GAI7DOOGPt
wcw2c6JRrjkYLCvwY+pWn78FhifIMycTrhtmrBRDwE+ECdFjjG/XE6GeEME4U/I1
hWjIuyb/D9UAddNM7C/x05anuQk+iMyHgZzLUw5WLbtGcCBHIiqd0K4KVXGtVICS
Tg75qkbbShWmEAPBSRPHllqg0JwZzEH/p2Xe1wbI32WL4ggYK3hIAho/iV2SB9S+
e+ZNcwOuI2O8ATn10K1RnXOkbhf+PRO6iPrC6+7YIdSjRdARN8gpXASllFuCt5I9
2zcgYK2coaDBnk3t/jmsv28XKz0MatH9BrXEQ5fud7UzHzNyXNvhxXM/8U1Hse/T
TCfLA5tL4Z8T3ODicQK+9XHCIW/IbWbyIRXUcWpzGuhmd2MozJ3DJFplwSuc8IN4
C11B6D3m/tVkBJae9aZFwl0YqErBGFo+ECvtiTP4JffOwl3mNgy5y3L4tlf/7Egr
5Om3tjKKophCla5Zxal9W83o6GaYSIC22bkO2AMwM7nesz+hJoDZVoBK1JktFNDV
xGiByOiPkjZRhbyu384P4Mr0inzvy7JhRyTJK1sZvM2W174IDMY0OFGJpvAVgyUl
v47kAekZgrM1GUz8EJP+CXfWl3h1BWeY0urnoYt7tFB3Yfupk77XijW8RxNVwkum
AzdwXjGMlUq+4N3ZksuAlvd1qzkAB+uaCehxR3+CBy89Yr9ZVcKT1eZpKHWiXDgG
IXHG5XoRCPxlUg4Pgf1g26LA2wXadE/xBxDa/qVdp3X1CPmr97X+aC4frfn47I5M
eJqvhtNnNdR/ocztQNPaibX+oco9At1NS5YxGjXkCNOH/88M1XBUDlRLaSVPt5IB
Yn4GTn2oLaYRt981lYfYqsL5V02zBF0173nb6K5+t8qWS3lH+QdqMhGuWCajtrPK
pfjLjW88X7kORRv0s93vVwBQncrzcaOo7kjs6rsYrsiQW+zFDgdjOC8pqWvYwg5R
KVfEmKSKNxHoTQiUbyHtCS+1OVQaJ1X1K/tS3iuBtQE2RH0OAAQxfjogv0PFVGnz
YxH5nGyxa3yO23pPzXfq7cd7taTuTXUENoWEIblqw3if4eLbAsKH5/eZbusRMpc2
N6kWPIm7d3i3GbI/0XgHLvYCuFaYYAfJnsRG8RrgdUhdpRw90yQOcHKx487TTfat
PW0N/fq5+nCqcuziq2B9BukQDNhb9ki/OP0DiMR/t4+kaHWQ0o1ZKcuePH0C9gk1
MxKjH9VxAR9gyIzHMspGzUz0VyPtyXUjwEG3lUyVUcN0t6N4PygSynJrAuXu6PiM
ecWG5UZr92EGCZQyX7DkBKcK01Xp2onaJUVIBz01tmJBkj85aPgWj2nDm8Fx+cuf
haySimUJczOm5oI8MY2sQpB8TAey4Xs1jY2LNgTMoCXLsraH+cYacgYQZ4L/t9jY
5Y+STFzUQa5iN8QLEyAEOOr6fVsrxcoRdUpFdLaoJBjPILGxg7ppmuz7loj7FgPk
V6J11WFXgcCRcfdkQiitT771yoiY5JK/5TW3RvbUv9s9ZzRu8Rsp4gn9qoIGaFCg
k25zfjCocFHNGS919RF1kay03zUVWczoPpEesNJoN4M+u1SxRYoLfwo+MAygk4Hv
zwGv0LLViZx6SI4cTSNgR3WmfCBILQgFCmODnn+fjoBVX2XO0G2CpwFjLEmC58o4
qUQYsmRlKvyWE/4KhnQNOxaI07LK3K+MiiY1z0BSfnNSf69JmPsq+X8XaflmBSI3
HrFR9QMUWIw9dEFq3o4y4s+TA0gasxJCL5U3qQZQ3iidqWkoYxRB5e1Q4y+Wqh41
uSSf3YFByDFBbTQu3P0OCfKBnmqqQty8njyaRB0NEUSg6ggc7oH8J+T1NDWhO0Ev
fFFNTPYQ8HaAERw/JR+LjTJqtzVP+p7BHgcJ4gcLMSy17Iyt8t8Sm0BJJlZq14Zk
PjiR7ZfL8U9ecBmB4D3A83ZqUsZHEL1kr/FV7AG60i1e4kOthOj1jdpXpFf1DIjm
OBN2TdPK/6QzXrOKlSGTwdEb0KJ2LjgFI7CHs+Rft4wTJ1BAz1GgBFXtfidygpXV
SgGb/HONFoVrlBRY2RXfiz4tMl2Ws81M7E9XWqZu9KztQ8De4wnPd0R5J/rh5s1y
csiJcm5nkEnxFqciS8qVGg7Aag4xRG5xr6fi3uPtCp/U6gJFLxwwes4YrBPxypKF
KoX0x8T/wwVngniSFryHX/QQ8ikFatEsGuj99SvfMhTyPwyf+u3mFn3XFUmKzJm6
R0L091YDcLaDW40uUa/v/hjCeo9tSSQ2HtDbQ8cLerOxNlopxJ4zxCi0X+XNzI0E
OVSl2nmb4q8OSHjv+8vP+KtNlRD7m9mwzu3c5+WfQZj9W2QV37JsIT3J9QcFR/Mm
hfadXyq3YNeudspw94AaYvXg270dEovrzExHKfHakfIoSWXt/qEuFTAryxnvBEiu
Z/ClGbdmx1isSzDtY07qFmbSyf0IlisiCHnBhTj/XFfAJbeG3SorCU0Wet7v0TG4
D4FtYdO7DtIgvXzDGEHRweuTylAyXfmdD3w27Df8n1Y6JV4zKBjtxovp2dyWYM+E
kB56R12KjK6vT9q7jlYZ9gS7RjVI14F4vgZvEYtnts2IicVkFmXhoye96B9zOLLm
4Bb5p6Jp+SemN1YRbN8aMCVSWKpmIbxUopkY6W/tW+kE3YL7eQEgZDU9iSxaVF4j
AxIaVcx54P02aOk1x4KubLcBHHyytVL0Mr0Rg/d2Uxs/DC4ce1DYW/KZONO4gZw5
6A0d3Kz5HleBsdKWp0QEvDkecBQXDegg59bJUHO1lxsbQ0CR8OlfgLp0GuRJpoKI
3B8DkIRdBUpBnPBAChIZEqGKgPnuwlCVr3Ocm7EYm3adH5TkKrj0M75DzlIdTfh+
+tw/bO1ljKSGBfH4o76SrfKKjEdrDFXkC3wvuXNHVnqUFeYW10IvXTw/WjJF87Yt
fKI9xgp2P+TNkYLmuLX/7wjkAk0GEButDx2vemMdwcg7jheGV1HCB8M9Qd9kKSWl
v7FpgWsN2n+DRa4BXtjt3uQFxhFGgu8XYRccebqj/wOhDDf/uT+3wAr+oECIV7w5
mxCuXsad0rjY+6F2GRZNk28RRqIR1OUF7nbW53z/wRNPfokV9MBwZsQU8cO8ZBnp
0HYVdT43Iw2iWvwYNey8+DNdcF0IoL4q5l5FoDNPbPzMzSGcSgfxkKA7Ux4D66Es
xbxQ2tgKYFYPN74fiRSXAFPVUPXblGHKzFlTwbfmbLTVkzJ2r4/hSFCh/vzFcEnX
+xQO3W46YI9nZU2P2+mreUk2Y5BKK4R3qS+I0HqdzdBnb76N6t+SsC72gbpFch/A
IePYvn5BQH/AdccIrOXRR6zg9SCCZXRQYrm6tJevQBZ4O8Ps9XkONNJSBFcvl18d
eAmv28SjC6LrHxtKWDbnqN7wsz82PNuNrIcU42r1w7VwdV2tA/CCr9nE5/8zHoUt
sAKt1y6j70Um9KlTCXyKNFP3gVWdWjwv6fS8a//7oz+WxaYhDJ0+kOlDnumNKvDv
JbD2cWHOGIDRczlI3yJnH+j5v7xh3t8+RoBfQbSFi2iffIE1kLjsDQlPfULDbcx1
JekUs9dMOeQ1crmIxvhQsSH0v5YEPyvemJyjrwAWxaWZEAJtr2+7fYteuD9DiT4R
IKydR+pT69ZtIOPKlm0Gn+94S0wSw8MmvmjdJVPW78dcMzuI9p2ub5K3n7A7zFfi
HZ2aXhtZ+dcW+tvJDaQXbR4Rby5SOdHyrPS/5xa0yDoZWdIOrZ7IFZ6MEj4f5mDg
vJLSU80ZXBbXDst56zc4ykLoWiUfJ/3REyOYseEbjV3KtH1cjdXvjwW7lBlFIswy
1AwlY+Fz1RJkKhJLoMvtZFRcQ4uIyPO7zDkvugdTqXo34HKJGKoqweP4yVL5AzJc
a512dZk2T3AI6jY9BKSUlH98xxcWJIPnYsw9Ey5S3ZahgkkiFomfOyjXxQikMih6
PZqWEg8kmh/sjgSoQZ8AHKGhyNtS2BPseHPzxJHRdX5G0riYboUiH8yMdpy2CGFg
MD2opnSCFnTzVMxQACxUs+U1Er5G2ZbhoJyAIgaxSiRqae2AuYZyKvil9o2u1b03
Z6M6zp3bUsIFh6QuuO7YOHLHMBuU8A1AnnOYfbeHD3arM0KebVrVNLC/f8Vn2m7i
BShoxYYa1GSw5o3ZmX7tTZ5iedaHCh2hteR2RmDqzix14sMFh3WBBBUDNmTwDOyh
RFxrlaAhjofI5DsstcV5JHTAZvlGD6HlDuR9oFx0VREoTbkNET3weEocCwNAJM5I
hwtxKn2u3nZx0TPUemWJFxeLZdmiIeFgZWGP4Zpp8U8RhQ6y4Cx8K/vsOka4bvDk
Ba5zj2S6r7VyfXkwiJVy6w/rrJYr5CqFKAbPtJLmtGu717aaLSebWVoDXKu5gyaR
CEdsPTCN4zmvs7ax+tPouaKEHOK0GUBQ7pEEWSmt3M1zCY2QUz4YYxKnDmpWn3fr
AlAL0ABuCHn/PY/rDukqfwKxEh5Uh3RPlfYbVDinAq5fSQHLao8/C+5CMo6yyqFs
SYcAmoZbcji9jnyjW3i+iH5sZgwJPMBW8YUFpqDfbSeXhJgluM4zZGHMwWBTnTkZ
eNuGHdFJ89G9aIudT+eq35BOQf8Kkkwo3HjJiNLIm+/QNOBjUAkeH/MtfYjZBql+
Vysc4F4WIHBihLEkzifLFKnfLUNuK4WhxYrbSe78blVKBWPuoWQvdyvPHYXzqaE+
FEP6ia4U8ONxT7ScrOAfc1IFc+hXD+Iw/9EK1R5/cX/+lsJyIhnFok99g6JvcBFi
gp7MonmZJDrbDkc2RTrpWSWmzKsjOQ6iAlz4vcGh2f1dju7ozUzHvvwSslds1DYU
RK+q/Vg8ovURkvtqKqL+KEKN37Su7dBiXgfzrEY9kNGzZVtGvqdt6pKjzug3hvm4
5QHoEUH+O2hP175ONocFVLURNE+tNFBe2FYiscJo77rfYTXFNeXIJUj+VIuT1KIw
jmQqaHRErxH/nT0NAak2X1Vyp+EzH0HX7kFmAr614BbLl0VnaBWn6ZIdWIcMUfFr
ZiFOcIcycfMhC3IO9juvPyFj7Sfto2f8V/DTBZNKmcY6XSq9AMV0sei8nPuMnCfe
mhmPj9aokoe8vsjqs/PnLN4Isbke0H9Cn2VK3KnZPHZ0mx7baSVpNIxj7s0BS5Tg
I0URa4P5+FBDcbwmSkS1S5/+CNxXR1JJD4JLI3rxM3kGxhybtGMx5b4UCsBaormZ
t7fYPk9Y6mzC6+cvCZ9YANX8UUomAxwTo72uU2aFYtuLEvf4HiQo3mgWr4mrEKdT
VgLGpoOE7pjmXCA6FuCqPfbdUovR5RW0ugZGOfL4/zOdG2ef1OhGNGUtyZP1iQXs
F9tH1nCDLgjW9hs/ebYPjxGhrgU2WAATZ4FiZuJ0GyhDHJbXkCqRkGwNuLCkD+q5
KER+Q3aL9ZhJfBlTPlI7WceTy96XJTMNJ8qTKwezQ4z0xD35gxRJK9OxVpcpjmmC
nugB3kBpB33dW4TBLRc+OJ4zlx+yEsXcHNdCmcYHJdDnFfmix2w8THq6BM6CEWSG
riybTUFh4w2VA7C1mWM+/AmKDMFu+qc3eOZxXczywjW8p6+m7otzhSqtMyVdOPNP
oUsbHIe1DhxzRpcf7P8eMOJkqrb0xsmhT9og8dFggAr3nLK5VKOSkS3a5NWcXmi/
xL/5Ijki0g9Wddij4XdGUCIgFdJvpewDA8Aag3/MGElb0AmgK6JX1TlgAurN0Tzw
BjNb57NchFxCSO8nEu7EQH0yPNoGQTyFBwRGzgJiShcoylTS5rBeOGnu9O97nxZQ
9Vkh0DkiO8Ftnc96xOncNLZRXKCcEBkzbVV2c6RIl/f0lkHYBXkmNomgwwLW2jOQ
kwOsHzADg898QHpviVDym+U/Eoy7z4qNZ++LoJ1i3Vm7v+VKNubK+y/Ldo2MHNRO
HG5+JiGEm7B/Uxxva18xHeyzmH6zMAGudka6EVzgWeZQwd0t7/d1tL6xP8Ctx2fy
k4FMXU3UtzYHBYSa/Kl6bSCQRF+yTam7GHpm9nSbgjSjDD/M4eT6UjDvU8hJdQve
TFD2aZmddI2TayjJZn1AjEpanRKM3I35WRkTGw/F4NYxPKdK9YZzcYp9kDSriwZZ
TJmClnY2/lcRq6AEYsmBPxdThnv+w28sNqjBtq4DrtaCtS9t4KovwLOAsGSaKCuL
pcr0tiKHLCFlm6+K4CX//Hz5jYGA8aACO0YbbbDc2K5ygIfVjU8xfdCBN3MS+Mtx
+uzjixPHc89etAxBHlg+VqxuGSYh06BtYBoKQ6AAS9b8UfCqTKL4gGky3csWEB3l
ulwsSidxxsbEA2DXTIfAKZSVfxOgqI//GCHrzst2KGZkCEUhklSgipw5ViBv2u+2
cuUWndQbMDPQb8pLERKIlf9aYK3N06Zxzqcv9N0xvOVpshZI/FLDW21YqwwMGGFo
f7H8cN25PDWk3wsM3MrjM7+5MD+fsiSbK5XbuKugSM3iZvzYCC4Q308ASx8w/LaV
MjJy9YUq3Trp8fK+YxrPyNFnolM/lb2eofr++pgzRT9fNhJtY55R7s6woL9Q58bS
PPcnMDlPqeVgtk5Rsogkp56YPdfDRz/1k2goryv11/wXbc3r+YF+JqtD37kskKIg
a85iEs6WfnJISunQmR/Rq4IBvX1iCc1/zhr4NsyV7FlqZ3YAqEvgO4D/gPgV2k2/
ilPPj+30nVfoMVRrrXDBzJ4DQsQGYN0oP6bXXnxFZM8foID8+LyFL6+OrXhzFxX3
EQJRqYGe6YQ482bqfC9ZsdOufEGuU4CF+Jvgl6G8VjnBWlmw/2WkaCs3WVS1qaRU
1Xki9fEzAnom62fMTJgV7nPQdv6ilxEFr/skXMkxWeogeubrMe+CgR6+Cac46H/d
Uc+xIbaU/gHaixVijIu666fFhy5bbiMMjddOUaEFE4ore58UqWfIaDnyTjaxkzVW
XiKd8sx8EcBFdWdKP/VP5eX4GOwTVr7K03z+ADTnvDwLs0gvb/jbMMxV/czSyhvn
8D2ZsuK8cHFzex3SfHC/D311icG2olWPSv2lQ+mebmFVjZVJQGQrLd71i3qRoDp/
rLS0hKTy4e96qi4zrx6xDWAhztTzSkPbnvmKP7EJHDmAnvu804tEPDRLYLUTgCgf
vHHkdzM7iZzk67tqaCbbblFwPsFiIxSogIbBOcpdwbo9N+54Zs3Wq001TWNYhuns
sxmaEcZ81Z0zdHXuWmeUTzWd/baLrLbWFDu6XGK8dDCLjWQXkiFuUhgStXHKlq4S
zo9XbB9Swqgm9VqYRNZRbE4sj2TdPbWGLxB5yzMgmb7XWL0ZS3/Gh0+T2+49+hy8
5G4c3csvry1b4g5efBV8vP1QxhwSnRUOOY/CNEujy97cJyU877E4RwFAF+lcSzyp
XZ2FyU/n1S6Lhpl9uO532/nj5pnq8/vo2QoVjosLRf26Gqgq/EB3CTYHHj7zOQk1
HgD32eeQPxI/Ye6inOVYV6HHEELrD9MJxWRSt/bejCnJQqc1GgTaU2AGYPv63fBe
92wdBt6+/25sc6Dydy/P0Bfx6xouPaUoOrbG+8nUI55KNtE0fiw3y2zdH3EGKlVl
tGPPT0xTwlycHs6Sh2gZ04LtKG194UdPeIj42PlaieoYJrbRXRMuAwXeJRsGd1MU
8M/V6orktj+IK/MLF9Z0ohroqj+XpKaOkrx1LY+eeweYUnM7mPKiJQUB/Oftum8J
wJ5UatBN1XV7N8oglUraJjLxArfKxtAvrifoiPxTiGK//GvAOddAfOjPV8OB1daZ
ZR0GD9uuARE8ga1MtIzJv0dPVSxhVYqK35U8HHIqT9XfLFlJmadPz9Xy+i426ZVO
cFNe3G9l5bJZJLLEUIsYvtmVS0pIPqQqE/otspHd/gfg6aBqaArHpHBUQOTwwvCR
6OVPN8td7AyQQuTPZK5cIEy1am0yzpaQU+oKwCue85S7Nd5C1uxQrQpmuj0t4K84
J3EsO6GELVScvA/1nnCBnld8D9pLW3b2REqaduHpb3gNl7PWzxh6a28zebbqN6nQ
idYFSYeeYoSxv44nzwsy1afoJxSOrpyxfF8eGkxxi7z16bTvbtMYsxbwshoaE/Nd
P3gaHr8xZPHhGJyDTuJopHZMpc3fSW3XaJ3F1SA8nMfWFLCyMTEcHu2y0tArP68V
RCQ0bpJnx3WgWBD9ysPINuMOPWDlkfO4iq76Nq7QrcGFs/bT06NP+ObGQBzywgXG
N/AjObthqLvYqGR9h4udDGU8Hah272y0J2Pm3GybkfkJ4HsWOk/B2bX/GDjwoyaR
JEJNRXxWABkzqOhqyIJMKVbmOhYK2Cjq4hIVM1VL47Y9hDcDnHq2mJYLN5FAvuu1
zHr4oKrme87ZG62LeeOSRwTscmOYnTWiIPQoSeUL9XPa8pW4AZFU2GxMMWqPb0es
YLCPKvb3lLj4vG2iOtcBlAa+g0qeRJhbJ9AA6vsKFhN0063pIDqsl1rfofFYUr+O
LI+0AH1JG8fOdvqyeeBmYNjKbnPjQlFlSDbqfHzN5wPfB70EBe6VfEnvocYhftAU
tY0uMrJlJDwGMSSWzVSmNXZpBPUudpvOWwCGYJAK24MGRqey/LJa1SvbTmiwrjkw
4gt8N8gSnGASfM4rJ85UmGIDB3PpRiGeuDQHAkFooDSDtDiwITNihACm2hcCPpXr
0yJByCXDRSjGR/5q0lv1kpPKYFOjMBsSYXAK8N2uufla7DBNYN+kobklGLARGQJd
FJqcnaj4W2UKpuNk4JswHJ9F6EH0toV3ayHWz9Wn7ess0wkDDO5vsSjjW0w712t5
k2L5YRJbqtnsCOVbkI6nx/vRMg+XCUTK15VYX1CphaJxEmkPxEXgD/31PYYNKTE9
tT8yRdz65JsyqhiJkGvxqL0QP9dksregzANGubs+jhHygkBKnH8vf2yl7r9gc6jk
TyXzb4chJVTKY/WxDGuoutZEJsN0T1v0VPjwj5yPVvKkKHywhtE57uwr5WL0Axgf
ofx8E6gD8AJWu56J8FkkLQ07gxI9TFG3iM+7KDobNCmAz6fnjauRVzDBbMyHvzF7
WTIP7Y+blQnCLjPYy96wT3hAM1HguX9m/FMiYh26ISkH84aW4MSA+9g092eFFt8o
mLIc5QZz8P07+EojQ64BNp4NCUzAlrZ+mC3ZPoCjr3jJB8huCZ9dxxYSbaYOa/q7
C+7+aCiswSlAvPpgxcVCSOOdru1BtTuq7hlZz5r41YrQRXT96V/TTktUmKGHXY+I
xJFlvxxZLnddoAejUQEuFtti424+B49WPkGM63+yvjrDl80ZQfR3sqMPpAnszts+
U0k0M4Ds23BUC5fIO/GrHLOcJ/skul0BMqvUF3IDe32c5yjVndq3TniZq8Ezyrnp
/u9j5HsDqAXN9u+rTQAHCpPz0j8t+ARUqQUTmIs0DNjeP7Msig0Hl/HIrIWHm6aa
7/TGAG7uXvy6u1h79KDm/wGulU45tB0P47iyq39HMPEjO8a0mgIlz4nDhtHmSwfa
oP3yLqkYu9p9qwY7RnfoMjx+ygL3J+dUMEjziurAbyS/wRKpyP9fav7ZXZb7JT2T
OGLj+UkY9jUxt0zF1r9eOCWshXleFR3VYaLU9pJpyaYa9SjP+1ZXRc8UrHKGeOBf
qt8Omc47FXbe926se7z+Vroc6DkX+T7SBehB2GHfoDgqiszRduJvc6bTWfUWfpo5
I45543uGHW0ooMyHsqMuQ0Yr/GgRAoIJ6yOTCbu/TCGq8bUJ2LMd4D/B9ubCEBmF
YpDG4CXbkA6d24kxZwlXD1A5Vz43MCyYzLYuFMFI88ya/RCmgS78xASn0Zrx1HUS
OcBdCZnFWJ+Sue8hbflYTPxSC/VwB6/TxIv37GQAxUu/SPDc6baSJIwcaxZJi0ut
N0A0XvoD4LQtw1TGaiVUH9ae3SHHhOdfh2kRdlZMHzNVI+WcxHxY2rK5o6XIA+w2
jcOQzMOO2EBM9mbBII9694GJV5B0+/ky2f5NSq5OJkTL4xtn3xYQggvvneBw6/Oq
3wbOTEMqf0wN7fd1H/HQ+nnpr+wtw9U3fDp8O35w9+Wa8fOytpNSdNAhSN/8n6om
9DPP4ejQBrMNR0cvv7izz3gGdwgvkucIdBSZQFW/sN++p+tp3QaQ7S9Ul7RdQYSl
Atpn1wOqVLJ5QvrFCH4yLOM4K8mlrd8EoDxLBhXPfjlrR32+mw4ewqBQbkT4bGVc
FuWLHmrh46+HCwwxHT7SE89S5tbv/9wQZFzS5G3zl8eXsa1aP1cZLy0ThMtYBLok
3kYCXvfSBfF+mTApYlGOud7+5Ue6bNQPZ15AC+IQYUx1mh8AlXcJTOZrKNRseNU8
cbgT1khQEdI3gdTq+MYX+XfAh/+56ke6AeZ8gZBKPunroxugkQCEKD4EeDayAd0y
GH/rSTxqyF/dNozMm5Ra4uPMkpXVCPszOq+FblVXBAzrVqyfQOLnCuX8Sfo6Kl/e
AjIO+c0mZcnlw4nt/o4bj/PRA3Lbpd9STF2ebF5kXKqreF73oKQi0hmO/Cu0kEFe
YioMU6BqVSgb0An7Iy0YZp5gbuNpkqq8DxwbzAmmlmWBRqHzb6MbLo/38qcgZSxO
VH5EsT+l+e0AzExSxaTExRZtFNXzDaT4em4sITF6/+SE5F4oxMcDn2AU+wvjd3EU
N3TFjb7/vwxpLGKB+RfDhr+ZG7QfOZRCYlSvy0Hj1W9Lx7NGKaxsLEZZVU4e5ycK
BEPnklmN33asIpSo+aJYoB7RaK3CQulS5zo0HhxwdeaDNm3JVb4zA925xiOUMPPJ
RI9iq1qIJshpJ6jk36fLBt5A7RxoQBD/gUoGAzgRq1u+7PQcG0QLvQg3d3Y/i6EQ
ZvcvxLG+1EXpuQmYG9TlA4ohUx5Z7s8rdjbJNnd+zVCFD1ufGpZSfB2QrZwZWrQT
DpvpAiuNDqg7+tEfPUiST008W+ckmi5dU0YOHPsx89MdNMc1URY9m7l86zrtwlrT
8MHlLO3cJ8ckQMjRCxdEEpWzZwnea+n3WYHyQUqcnDx34RVrJPVmdu7dfEJR6u/c
QS+SpkOOkzTrnwH26+KYNRSNJWbkfZs0wOAuOormXncs/9c5nY/zuoDi6eDXZgUi
50q7Qn+IV5ciBkQY+2NnbMZd4puUf4heoPqHoEfUnAj7VzY921lFvAeh/LtND2Zl
DB5x9L6e78FWQ2B73dJFbbU+0rXKNMZFY8dQwQc9WHrmPOVA5xxiT30wjKbfCG2/
xCcVGYA0MRGXODUlNKoiYTdkhaHJGO/8FyyX4h6LPJe0OOP5ixHIKv30XOWk1pL2
An6b5K44osP1tnTcIDYSv6FX0GPnwOipOEzw6Ky3ag4xwuqGcThdXJ7hjKRprUHd
QBLQ67TX6AnRhAsGTgyDRLvfZ8ZdxObF1f1KGlXRasnewuMJDqWWYpOetNvAwH1T
n9Oc/y3gzzP49eYqFAjl8mo+wAwO+V/RdHVrWuMG33PTupVAXQe5JJbxuL6ulV+V
uJPdVY8hxMLsHCORV8fnFUriQOOaN3ZZghkJg9Ftstd6VLBKShROOIHSvYCx3Ze8
QV3FRx5itxRgmhWB61w6tm7ZUzJqkKvCqwgMzhowHXMFs6X58TfKEH5wVXvmFLq8
+VUuux6JukD5GhfP3ZDYXx97/GPk0SbHjaZeCOsJIrcgKnZq+/EM5kh+3cRDhies
KnBMZHF4WUYUKtAZZVQHuEW3uuAAmonKgJmNt1QDsIDq2lSxdhqxba2tYwqSsKOj
SiwXweH9WiSi0nsLvCto/oki/gN0VT0TxzJNRWZs/iTyJD+ZrlghRKQgVlDV7RHO
7d9hjnlXqjGH7SCd0OaRr8UjMRHgLteSwdhpXj6pYmsJA/ziR/rOyAgd5JdvR7bL
zwCcbhqCAPWqHipkFuRwHVgRohBskmKZYyTKQB0R5B18rxPCjzfQTetOm18oAJe5
fmrB0IF3NRrFZ98lAj2H9Uqr1GAQnUXpOKeegzsKvEcb6tka3Qkm60AdVxLVZXxI
O5yXihSIkcNs3NhN3uav1YfUgu5J9N6tgeU+SBiPL1pFBy1UxUVH0FhRrdGxzjk6
1wcqhi8JoGCkrBQk5fqy06qooEZaAGc+/KbYrbN5J+9diJLzgDs4sSrfNxNXpiF4
q5gpT/hbHpdgNWcAal0QHIEWfZC1xK+PVHM60ONGNhReg6ILvAeMzC9nijVBML3c
y8x24MT+vO7tPLaYVmXd0ywiGjHofjCZ3wWGB2NF6ePjeMzHl1PsM/BqWT7mcjKj
dti56jfKrhgljWVfA8e4aP/V6Xw+qj+6ArHxp2na9ahfFqO1/5bNT9gAse7HKHr7
BurNhHNwRH08kIXkFo48yseJgffImxMO8cOqGSWfPYzC7bdJBMEl7Kxyj9At0zb+
JZLuZN9LYwlQrHqPMwDD7NNp5nx350hlZq28jC61uabIwvJCmYU04Q91Klv118mZ
wJ93TOMsYRz4y9tbzo2285LfvGK1wdj3J/KkykF5MiPadIeM78KyirC6EbDf0eZS
ZGruUN7XNc6PJokmrFdgIlg5Tad8xvj7/0MMadyOZAGMBqCz9GqmhNuxPrcsXsVp
qiHHFnUCOYQGcRfQ8JUl15OPZvAtjy5bb8dviBpqFQknbFxPnSQxJWg0HVhZ+SH1
Eju5aB7fOGRbAdgq89mINRXqlY4qv+/T4ydtTFgYmD8i8UQ1GkGvyj/MkUTtL7U1
+BfV1XpkQxeu/PU7UWXHNVpYDU7iRESs/YTLqV59VFAb3JyT79BYdaeBymRwvNys
YeG7L/BiNSHRNSj4z/LmbcknhQUviHViFNgG515eRiHj32oL8K++2Gm4WvGqsEhT
N9rZ8rwPXuzjqkw5yvBk+hQfH5ZcaapsP/mQrmEZYXVa/wH5H6pbWt+AP2H4mmoc
q/b5lxkAxha0CtCVsx5UZCWGC3dQMSIDN0Ibe0ovHaqgk14Is2QTGLekVkLIqMHn
4J4kCS9mSIpAxdzfgK7IhiYhIglUwbx5liFt4SpkfUG7OPobzyR6sI8E1GRehI/z
MGWvHXyxRJXyDsn935/dIe7sobubcaoXCdhuEuvSEiP2O9F6Qjnk1OR0omOcwN8t
+mSFlTKewXOL8lT4tyud+Uupfcu+vvH7CylAAA89XIyDT4VDlwZUIWsBPxhVz46s
Pro5dfrHhwBai6rqNA1/5Osr5slV/bZ9057uci/Axi/Zpk8aOfuYEX28O6YBoZeG
MAorBEw8L3F1estDlRXwMBWGH9ZvFe0jtRy09BPFRqR2GAWNBE43ZcBlVILUg2fi
Y4SVwH5GVzX6i03FFdnt6q8yTMFjTO0KpLqHK6belRmC0sR7jsUP2NcHG96xGE1i
lxGLX835GfPFtHfBqKPLPdjORLmAKuEHV9qw31uwxzWbX3sKIF7nnb61Ay0fohP2
N7btS8xkG3s7yz9WqBSlZo/beVk2hmiwiQ1KZ7wbEUNpLslabNs0yESXlh6E5I+c
iTk4PNOtRikcCYO755YMlWV+MsHJHiTsLI4i0sxKqn7QRcMb19cYq56ZPD71OsU2
UAEjGm8HRqDuFLk0SVt7haFJSdqXLDbIo/YfmI1DdPoTFb5u2m9CHnCXM1Izm4QW
BM33kf2q5fA/X/491meIQS2IMV+2Vz9xz50N0lzrb1qdnkWsa/K9hS+dSdqT+UND
94BgZ5x6yU1Y322F5nqjrzBNY1PbxLxrnMt3U5a8bfpEjFjjdeaSbWeODZZzEVJw
uD4TJ3uk4M+Tf3LcB9CbBITUWe+7/XlVI3elm4XuV9l4sFr5Df3jePentglSAr0W
kRf6CFTBQaGBDwJmXTXl0xO+EVKm3gaxrzJ/8bBbamU2gpX/+ptEntj92vAVzSIl
fHCuzr33sp3BqhNIUTvtuSzTFtJuPO9nZxxImdfS4iFeHvfrM7BhNzt2Px49OiBe
koRRqz27BVMSLO0rFXisDPnb6rBLDeEc6SiWwDlo7SN/Wd2/O0rtjS2hAvUN1xLu
Odegw3MnVJWDCcdEm22ApraSljUeVPqXIRTjQGPS/hr71awDvFbHP2OE7GPFaiYa
7+KC7cUhM1Uepr8TOZ6rzrDbqa2uXKr1Pi3RICPZ2nbl0ymbSKVPL8MN3zzP5NUM
LSraVVG6gxgtMGD7WwOi0x21BzlVgbQH0CURdbY3r0QB9aW6sd1jgzVDIXYrOUaU
ET9CazGEfWWG2+lJ5QOQWF+RAM/SzxYYiobENY4w85jM3It7RA36e/INcPzfW4UV
1XAc9pcjHPOpnx3nJnKYsEilyS2RFXy4xSDJA533+cJru8aIuhPuJFPeHWnPlOIr
LQzr7627XnB3THKFigCC65wTxGQomJ9IBUstb6Vp4oqt88TH1o6d2Y/rWKsJ44vV
jmMMGya20BbuyFzHnjmBEGVdd/EV+3wCDOtneVpsPMElMCaelurxcADKimSlDuvV
RMQZRBogTLalickaymB/Wr2aGUKmclcDm6thDJmEnywfIoVH9/OWkt++tOPGispC
6Uy1uEbiO47aHKL0EeYaxmnFeVxd8BR6V/rdoBJfr98uzjAaw6FOtyKbs173LJNw
gpCyjUtijpx7WHNsxszaKkQ12NhQjCU8mRyTj4CRx28IkYgi+Haikz/UuvzJ4CnZ
kY8pqF7fN65NnfeyfndCL7RC5lh3PUGpHG9i4ukuo9+edWoTe2zRHmaq4v92uFFU
NbSXHB92j1DpQIOOrhlEUnP39+cN4Bcj9pqEklFdoHLYPyBTGI25LqLBuSbzQ6eE
cZ1rTOIoRoyPYtfqpI2IJgsupmjjWwLBYXpV/yxD9tC8n2b0DfHbYceOUCouvuwN
J4cPKVDeie6wG9CqdiRifewa+wtCQVhm36mH1Lrz0jdbGYDKx2s0uHzprYRSImS4
wHsqlTKL0w2tHxEDs1V4MdMnG/PuID6m1Jw/dDoIDqoqTlhV/qX90qc/l1ybR133
oaFrrvujwCuEmZ12HbSj/PTHhosMB3fkX9li1JMZSAG9xq5CUWt5zttP07QN4IBg
+f18dBCGUI4j0w9Tnpiql3sDtT/45n95QWuSMuWqo4S3XHua49pFlD4AtDnT7urV
prmYw2nPqOAuiD7aluLztS/tPAfycpK5vgO61hrk6C90/jdT6rZXsUihrvbQPJjL
Z0q5MylDZ2E54206T6QOUO0rDgUQy26WRE6indyuN5d+d9JYPWMQPj5zuDYunyNR
MsdnkqwyTYdZfoV8CdBDdvhZRbfXnw4W8P0funS83BE+3r96GYxXOpB62PYmaUjI
d64RZoHZvLhkkSKA6XKFVMzvByud+wy8YBU/X4fEr9wzGF5w84kL/HNKqDg6CEVa
Hf+Bh7MJWgi7TeyTmiRjob0UzvOrTCbYhL2SmKPqODBYVEn13hE/xmNDCnZ16KMe
SRQa7PK8f2A6YQzgxhqSjarnrcZpMpmoKhy0B9dU2uIo38lSaFxkXxvKn4tTBJ2z
Vofv5ojNx9SL8XtTNiX8T5sBfJ9KedjzgYWmiJiZ9ule2lOjBS2jxtI52sS09MUP
fynazWYuGQBT69VwZcL3muyofNfp0lVU74+Bwx0ukhFZCaehmgCw5Zii2dGhHi3v
pqFVluQk06Gf0WSmHZz6Qgjp3IHJnVKn4BQPl5v9wFejytkfqHTelIU86KrqrCKM
a9fRymWhkbCLcypv3nS8LB9pmMNqhvgj6QAUGYwnb/uCtBupiweFneni3LJSt+47
xNNOFYf7F/X5lGG0gUAKKU9WsEjYRooWFb32CMDhpb7cM4uQRczKp1aHzG6g/+oh
uDjX7ccE2FIsuuZeK+AGPqJ5NO6lSWnyscCAsQ6xkA+w26sh96utNT1zQ7EcY38m
lPor2JLV1IKVCCaJ5q4t8ywYgFfrSm6Mz1CcDzoGCLqegcpNFZwpVDznlqDBXGIp
pxHHxkH1NQQWlAcfH+SqJ+h6tjFtuZ8VL/ndK5HcjKubeWCrcji5NEgxSwRxZShq
9+L1DcmUY5ihR2kiJqqarIrMYZiWNzjA+kWCTMUvjqGY5pFQmf2I3xChSzfe5WCC
avNtXkQmY+H4VFsspnMQ9xBTFQcg5XyjIh8HamVvL7JdjGOVQ2vV9k8WHWQjZKmt
77PXTCU8wPbjoEvOckKvlgd73s7Xd7mG7iy3lU7IvMn9e6ba0EeFN8QI19oAhv4j
iTfxw8ngG2XE5SQ18zs9+ViF7ov/G3e1RZWKMXIxHKEHqDchcaOngENnhp3KDH0u
DZNLnN/8DNXzgX/n/883XNV3X9cfhzZD3OLiV0/6zWaxV+QrQhs6lDWTu3ipz7MZ
Dhd01MpUhrY30847ZkQWC5t0nlmJEmZKAvuXdfU4x60na1z9iY5D5BkZOxWm9y6y
smy3XkOYb9bVVHzegFKDMJPjqrXP+lcgbSepW6WM2cDr7zXfyuxxmv9KNs868MUh
qB1fboPV5GWglszjr7sepgHuJX/p8p4260nsmAuIMwUpuv+pwl1X/YGvPv2xBfwv
HyMvDkCG2TOe494Rugq1zJ5TT7I0jAL9W23Vml/cHJzJ35vbxO7jPMf8lI4AzwyX
nTg0xrl61FPnMI7wSrPmwa/1sW1Dh5Qgd1LVplgth4T6Cf9tj7rsLiy7MfoXkKoy
bZ8T9nx0OJXV1Il+lcU/KishspxfmqBZG+KVS4c6OxEz1cNbmk3I83+5/yeHCpDN
+OvPoNX6qQBKwUVUTDFF9I90zF8jF0fVbt4anvXJzA6BfiQhfM6ilie4/K0qDpVd
rQszJSv+BH42Hhm2tBrtr+CmoqiIGA3uGltkpni1j+Yt3FoeZHUplL44qJkND0lq
ayWPfkMrF83OOnSHo9cpKXLTXWZh49wPVVy1ginKMcfUbbrf//Yp2sazcSe/Y+sY
nNL31LMVYaz815lqCNh3/JsqBa64/I1IU2KlyRY8UtqP2DmkBrUm3pEPq495lwvC
O+KdMUll+zkkaEAeSSKoy4UfBAZ/ENVYc4UPKw7vR4V8AUUQ40LDYeJLz8q8sgjl
1hTWGE0zAW2TsWLG+uGcELxbiZH9rResMwmFU+3zP9pAqCMn3A2uIfi9UD3tcQkc
q6Yr81bKL5bWA/t1Nmu95RAhb9PsXprJosMeS32vEbJR5+I9OxcvAVApXnqPOxQA
2yQ1TIfDOay9h8J8OsmHbq98sOPJc/Yb1ipR3hOTuxumyvedsDwVPxGytlkqVvP1
LpaULxT99PLMO5nbmx7VhLr7miAr/OJU3OpAO1G/1HI/bbZyr/hJecy067PquIPi
FQG4e2LtbQCAB+EJROg/7K1wkNt9oX1Ov+3LzJKvHqKk3EeRB6T0AuX6O9Z+1PlW
j++JES36MvXRxvPxM4gB8vKJ/G2MwgAhOtg46eyfGtjJg0ClW1uUlok2eTUo0BoL
xGZP8rqNQyUUzwIw2ksg2lakMnPW05wVLwlJ463VESY/GMZBoYoHl5b8J+JPlBQ5
4PnE/iwqms4ISsCuIEU30+2i7cwQ5EEqgvamdb0TUJ6ck9XhZxMtWSaC3zebafAt
flmqNrmBY4Q9kL3hA4owaUlOt+ilmW7wl5mPm+LEVVR+UHRxVQsopVwRVIkebHrw
cMw0n+ZLbbTtA7Habn+KicEZViC7SNHEvaH7TOpiKbkAot9/OH6av5hGZ5w79eT5
22+R80qEr0hnR2JPbFJaeElHxuGluBI7ELJC4INKcbUoojdiaV56NN2egMpat6jm
oWNOUpN8MQwgVFijI6GMP6DkLBKlJlPIDcKCGjULFnvhgjf9zraqtqFi3bq6HCRB
ZNlp8yLRPCyCwNXIuuizDhbIKDWRCCIFYCU3upHvL03t8tF5ndlfBwhb304x8gvR
uEa6xTTfenxKG7lAaqRPkHcdUFxNiZ80z6ZuO7C4z4zW1s/1YWBKuYye9Of5DooJ
OINQBMbMTUYhKJAs/jh/JKMZGs/EMT0HZrqLG6L41MnCIHMaNRpG8+fPe+D1+oGr
4ol1X9NVbca6avWms6gZO3nkZBY10raULZBjsKP3RA6IwFSZQbbXHxDcaqDwPHCs
cp1f/uM3+Ijxuxz1yzY630Nm2FozX83qcogyG3xh481oLDH6USCZnWjaIMX65KdT
F4Ye70TK0oP2jLbFBUB5LgOd/MFFXkdWYQ8LVe3J6hKR7xSRX3AnQZE7xTQR9F1z
O4UkiDxtBCJ/d/qXs3Y3Pj/fVqv30CgaJZ8Bq0syoH1scEjPW3MGJLigtbD9fZxt
mknVNtiQEGc88VwGbk2aDXAzZ6vlbDvtlP3SjorydowAun+cpL2PnHQAg4wzfbbo
dXGVaZuSJB97FMup3z2UzenNYpgkPH2JtobzmzK0RtJrZoCdqDYuoXbtvHorZtym
b+0iSGYkTs8UpLGwjckzDmJpyijpGxNMge868d79xDDz64n4huERtB2EsUNJVRis
q4zELs34eyHh/oEcLzCiRf0fneN2hI5MYJGcs8O11dkG7rvuYh/mfLDxn2TUuH6x
KDF7kF/ZmdENiIyAgyZusMHgolr9wEdYQV8iCs35IdO9sa88J9X/aGQdR3hC4c40
ILo69didcL6VMqBN93XkxSUWugVYZ+MIE9InQjcKHxDKm/GEjQWV0aeg/nHwQD4S
RdZyzKrxLOx1sRKR7XbJQZp8ncVqrYjCokMKOvU1+Nn2DnO/k5TOSmjsoQxUKI9S
EE/zTs9K7VwMOd+5BpfKDmL/xU2SF1w4xdStvRLziWm/Sdv1GP+SbBG/LdAxbMmc
YjvN9qzbKk76YvbIDSjlQXAcBD1ytwYVdvClQHRL+EYeuguQpst8ZMXNj4ihBbDn
diDfdiKIJBhjvTIEVsQikSOyUzz685Io8CpC47+ausF5ILkLRjAVmfX/HoDSACAq
fM/TblvYiJN7qakkuA8Tg9AOK+OiPBAzFP5EJzP6d8w6YDsTHrSLrZOfiMDvkHIO
RddcEXMFylmVRPf7GjTUJ1D64rLVOfScQ1g6zpzGj5dT3KvIzE405q8zNbm0aOzp
AzzOWJI6GQoZaQBbFihxwKDIw7LrKYmK0ghj0d2hVwBKprxQSlQ8r2WeBX3oRW92
wR1QuPsUGSJwyxtqoMGLadRONTIxGhHlEkTb0D80oGpEs0lHPE6MPrxVXflHaUQ/
xYLayWJouLecfScFPS9wMINA6DG5Rb1QlqKctMIXa+iyyuXfcrBfWCiBpqDiWWMO
OdqfiGHbwidro/2d+8Er9TJnt5ZD/x387+JnpCZXMjPjz1S7hn2QUTe/dbwpd8nM
3qzoXhgCsbEWipBebjPuwt0BMZvSsUoJqgIGlBCfVqh1Qu2TBChXicTRWX4qfYFn
KOZPzce8fSE2wLi4NafnZYq/NbJ6yX88Rpz7fZoPpMoxiZQmZxo+qmPgU/c4/8YJ
Ylfu0UWkSVwdOxMdg+ENCNPWdf74HD5Ztp7hVjWAfaf6lalAzd76o+KuBaHDZUwF
1tCK9k/Jxvv3yHHgA6aSHFqX016TcvJp+ggg3CGISXtu9xptVu8ASgl6WgozJOoE
z9jobX3GdHa9xSPm8nqY44tomL8ey+tPAi+szUiJ5/tyJaXvXi2ndsMAMHhU9fEB
Ap1UzgyHuMege6bL/IDUcQW1BA37hhkhWdRpq1EcETKRcImWxppVwPJNNqFrYiQn
oipnyhwwfPgT6PO9vr5Go1a9ZYAUnbMEnYe2hTd0mwwQ86hsfEAqIsd8pEmYUhTn
E40WGTbsSskOIM9LCnHPovs0cNTFXK+Kaqsxk4ft8dV4682sSIpAfBHPyLrGJV3a
lACE1BspUms7Bl7WQOwM+753bmEKIw7+LbIgnqindidT3yj1YXqTv2IFK9fdhEDf
aUMwVZe544LLtnXMUEOjVbx0kUsFfr/ZNkixmDwVj2G7LqmAeTS30UiHMqXki6T5
e5NyWxfPLnsfTx2uWUNFDh9T+IkvqLdHn8pfRs7gM1XfDTFNHQm88YMFXTnmKuWP
6V/ApJHZ6O+XiyflJc1HYCZLJ65aGoLTAKM7uymz1qx3BZGI8OxkGmiQE1eEeMh3
4rVhMq1Oz9HzxdVLeIbjge3R5Y/ORuGgeyed6+aolOvUTlxQmOqTl3EAvJ50fDa5
a/TO6gWQuzlFg2sLrxxN6LYhAiMDiy//UVhERjxc5RxG5ipkoYcW/gVKmWu0W9pO
2ZmaWnaaI93Ea4TUrM0T3pV/g85u5RsbnYrn143gMdhkWzwY8WGUY+cN3WFYAeWY
Jr2pO8n4rllQWTxG5qsgnUQioVjo+xayskDLLsXg7iy0SBDLzX3RdzWVLYG3Z5O2
uEXsI8xM9+rqycJSAU96QqH7nyomdL8U2yPeHrtlTZgZKMt4Oz3wuwU/7BwGUGvr
6zmRaftCNdWk4ie7OY6So+5cXVUinMFPFPS9vX/tOA/KNevwphyu+QSaJnyVi2Ak
4fJ1cewMzCQlay8e47SqF/PGIHaY1YDHw5EPOrlW3F9+yooAsI9RGG1R9HnlSdjq
8Gz1TSYjgF/PZvzBUunSHBm7ZHHB0zE0o8yHwvAAyWfkaF2bM8n19suxjZnLWNYK
FlPnloYED6y9oMZQYylzfH1GET6VteRuIS0M598XcMR7xclKr7WM1ztz3Ju/5bUi
LS56ZaCOPqw5O0m95vgv1jeHJqr0XBxZ9SKvICPkXTWmhVhStOHIrXBQnWasVRQ+
iuFjpOYoWJ4J0N4j1mRG5T3YqFzXfd/T8UiOugAlT4cjHqSgfjyqIfBi/aBah0c2
JKh/Jto2kXZ1zJ4bRFWTJEIovoWdaRuV+/rYfi10GXR+Hxw5EmhW48mi20XvR7XK
/dx9t0Kk/yh5h5QkgaJLpo/k10tyKNj1QzR2pYbMZKCCS7V0aAgpoTQxKvBbNFeL
VUOKDRmGjU/e62t2OIPlXRPU4MHuKEYugfB703HRKTQHmHyG7Qdo9RtoK0cZ5vV1
5fq5n1YsCgfFB1WCrB8jdFKTYLPQJNFN0Gr6gYXPCP8wG+w7fvxA7gdJE30PRiB7
aGExi8zY7VrTX1n0fmBR97nlgsY25i/6UVBJrIYk7N1TeFNvbWTYaBhtue4itfPn
ehhxdf6BvQixamKZaOvhLQ+uV0rynwuUP+stGKDjbUWXCB4aKxHtZCbBu36TOqE7
bwQdzAx9zRhJJ2p4wqobqmo+mAmCfleb4iC5B8TC6BnxeyeWn794KdC25PUh5Uus
CNCpqDa3s9G614NZelQ3TNA2FrAfH1lS4il9usXsi7tk6ScF5kaEmgmnvrogtSkY
gKzvgWfeHtGT6w/LfS6eO0T8mYUGY/ob0T7vvsu+HqSYYlSeI5OSlTE20ZRmA877
+AEPTmYY4Xk0qgl0Mv7hr8Zn4Wc3+Ug0sL29oVSmYOIhXn1K+ZiFVQsGKJdUie0q
VrgeLWICW7xpQG7QJGi1bOUrA9nwHOGu29kwb3X6MLjoFHi4BlaWmjM0xSEZtIad
NXRlKR+kh31j38c+2RYsEfGDWQR/QTWCjh6UE1DQLvY9FrJzwNP9OVUiZHOezxKB
0nAzQJ19OWPYXBHsE1JDOdGCq38OlMFPi3EW3m/Y1j9/5lA5xuPLmIi1ZwXZSPZZ
gJ0HM21Kx/dynxrgHktDjVL/NGZ51lnTPe5pLa1zYH/h0P580a6nqvOg9gEFwKYr
FIefP37QlKo7tMqHqscAPfGwrVaHHaJt1FXN2iYzpBqgSDS/6btFCYi6o6c273xn
3h667Kcft9CyVwFCBWzsni6r7jatbLhyNkHnk9e6WpBG3UWHDU5mZf6fUdml/BrW
fe80iYfh0t1UeQgt4TLOKXuSEyVaVwgkK864d9nxpJMj0pDLMrQHKrwXKCvj2NDa
EiJU9AxMeMLSXaK+kjywujcZ+/t99Nus4PB4UAF1ORhj+9FrNjH3uUWTTjU1PxDh
VuWsX1ku7ML8UNNnO7bkEQzBi8aXPhJbWjzyqp9nggfs6ALVvfe53SBP7xbHqJIa
wbUofg5JNGpGnToLq8LuWFOnwF0xb/nwpE7y1QIw2p0nbSYrEzMP8qEPE6DydBoK
oc0pBdZ2reXC+yTAQIm50Ic7qLwXcxCkFJIrUD+T7Ad0FYSmtgauV5YLBzOEwno8
eD7oWTa5HF3sXKu+dGMGqbIB3p52lOpwVD2ige0wB3TzcEmLMfaKhZtUu0eZyzOm
oCRkY6F60Sc8DRG3kUblppIRaxHsxtow5cvmde68RywiQDyoWcMOBrBu+KpS2CeG
To2QKKFpqJ0OzNIRs+LxvtiU5PbFo3ChoYis3aTsn4+KapdKm2RB0iNxMqBtugoB
zAyeO8y9UhToB+Q3PDVuO6gPqnP4ru5Ao61BsAM/BaGnY8jC6f4Qm6I5IzDSxNZv
/va/PDsqJpOIcEc6fCZydf/D+yHCeuhIIGXnEtnzvnerFt037M8KXKu4y500P7Ms
6KwsYpXqHI4bVcd+x6YuSrb+PkQQDM+AhOMQAPuInVheeh66dtNsjaTYhZiV3y8t
1mCzn2kvoSpj/B8oy5ejuXDWEYyiqg63WpVsWnK1dEs8MOTT28GrmwYhpYmBUcAT
y9cHTZ5vA12DdZXaP6KZVG88vlWhJI+c0bu82fKF9DXgtPgk/F6VSnTFH2Z68cD5
zCEFh7LTlz2NY1dR8iOKgY7UTDjlrvvkmZLYxlHi1/Iq4my7xswRU+EaWM/s03+V
o+kB0C3kc7qcd/mHo+nw9hwatiytFv1jfac+ObrZx72G9ldQ4SEooQvBN4O13tkc
bAsAAsk7yUJea4ivZn0BazkDpybSoyGL811ltZE4bF/uXE7Z4LRTDhD7eMsNqs53
58kY1P8ijbzlpeyxvr3Gbv3J1Jbu+FiQLzR3eINC58gURFl0yrA4NandcOYHelGh
rA0lZu+vNAHzRWbdxbA+YcGE1laJ7TWYg6+oNu8TNM8Uj4Cbnye6ZuyZV6DKqN/0
zp44vtzqYeWp92z1hKmyMxCSRVc/5DeZde5kZvgr1RIVnwqsAY0TgOji56ODBhWp
KKiSB61FAan9IN5kseuS8Hbp+ZUYI6ZfXW8Ztl3TEO6fNg56N2RigEJghrXYMXjo
1y59L0obsQtc4u2JlQnkg7vQAekrTPumE7j2f7ZT9ggB5jSgB0o9V9WK9DAnnnOm
RrCykZjnFM3P8hIVpM3Zl2zTZSmY1EWYxO/SDePF1QQvMKi5wRCftde/GeGLjbbx
I1ik07DxK/Du9PNqyW19Uz+mtZbhI/Qu98Z0AY1qlSAANhsGmktSeQFWiK+gBjn6
usROa3H35Pv2DX85Q7z1Ud2IfzhA+Pzwy8Yog8JR7zMtvLBOzwJeWwd9n/D75xhm
92Eq9wTMtM9RyfOR3z/BdYETWepdRaQGhlAcskRAXu+echzeFUvEKU7GJa98H5uK
7DET0wz/bPOu4pq3jpCHpLb7GCqC9eMa+Ddk8BVUEMae8wPdKfrw2SWxP24pVxx7
Ft8e0Bp3+xy5xjpaD7cCxMLh+HgwjU2ec47DH43o3Psiz7+re4CeKaeWbty9zxQ8
l07h1TbwSgLvwSrWLV51WFq/DIp7SIMh7wV++MvMaV5TVnV1ki+NpR1qd7GEQRUO
c+/H+NMwOgJXR1jub2VuzWTsdzTzi8jxAgk6qTA0qg+ceD4N+krz8nSH57b8SPwi
R0wSh6D0Xfu+vtr1RNnk4Be5RjYAiBBrzUxjQ22C9rZUtVLvo8Na4Pj72SbftqHn
7wAiM3DORm2Oz1MLQMHMfETowQbdaYceLr8ab+VnEb0Xv0jUaEptAyDksy8Heq75
JsWC9hEHcwZpy2E4f2zaWpqId0OOGtKUk2cKD/vu98/92wP3SahHCqLYTQjbLqZ8
RNl3tfLWKcd5jzOynsYGeLcqb4VTAPhR0czbIp8z+StSqY5sF1cAIHU95pgI1svI
3PBdIHCOghiVDdE9KbZSUtzpiWzMhtS6ULPev/NJQKUfbgbEPuhUtYlKAODWEcZi
T71WtZQCA/i6RkczS5NivH+7Ax76yW6ZtHgoeN4jCFUfTZ2cvcFjws/QNFLyPQqn
JLGu7Abv3Dj+WNnX84kRlZx/QLArsCt/83etnAvgz/K5c2jhDyrzh61rqXdmdQsb
7xvdXRVN9gNsivZaE7LTlB4hSzHz4BzF3o38FEYzFd5BETWGzicK71VPb04Thzn9
xTquA9T27NeZvwIscm+ypyniZPnQzaIqM3KKRzX3CmexoUI9ciGC7Se3ohgysy/N
W+ThgJ9cxZPvGYtHd1BWlRfjf/LSg3gSY2vi1OUK8kE7ihqjLpYviTKDt3KnQ/6g
7vXk794nbuZzgGU5+tuoPd3hknJ6InTyufAq1lCHHmf742oNPVte4Si+UIMetUpO
JyPA6I7B0ZuwmidCi8dKz0lOST+z0jeUKaZJ/6o63aHzXr6EzeIQv2zzvlaVyK99
fH8zBDtYPT1LIRAIQ47d4XXxH89R6TLY3TqRg8nK4Cr/zTrz275cpf4933sdReJF
p49n5b0KOpYWWzE9WLpiAN8iv+oEOYWn42L6ZMInkjm3SF3IzkHOmkhgDe4p42EN
LRPmEkdQllO5h2UOcHeRsZF6bclwqqb0t4p+F3OrkGEq2aEPLsSYS77v79AT7fV+
S2GGaRKPIBR4heUfhCDX41sxZ+hWqXsAZd5pvG3llfK/pcR3SuQNS/nnsJuiAPZm
eOyhQmAkxpoEBKOfHn61PcEQ6I4mP6BHV2Nog4PdMEK/7I+heJ+ApOh8GAsZd7RF
zk5kcEfoUyuXyEZ34DAa1fvNyyQ4cIIKbWegLfWNki0SkEfTwmes5YbFB7oxOsHG
JzP8jxyHpNd7M0u1cXYZ/TuFLoAs56Ilhjg/7fDm8axoMQ1mnEftH/jS1lAqSEVF
dQs+J3aQSe5J0BOhAlWq1SBdLtkT0sOkGSD8cW85jUcqy8N84f+MWJ/yMjTFagwy
Ncio4Ko+NWCzk/BSCh0Q4TT2h9jerhlJEtNGnUcRPV4MlEBH56FfqOruo25jOyno
lZ+FE0H/nlF0pddXBh4g8emZ55rGRjDhRh4xwhO/ilmJ0q4Dpa9Z2io2dcdvFPG0
h8YMx0NwHiHmWpou27U5W8aJj2eWV2P/DLGYTaB3SN6DfcxRiokc+Xxmzi2wAzv5
PZ20yV3h2y/4oQG8dnGsLkj12g2075Jh9ITyBuvBNwpaSYR3fnh9EQZceywIy6FV
R7ffmOE4dlJPNY0jZOvK5kHWxEsC0Wcn95fpTSu9aSr/aVY9Hy1deRg2TDAs5BP4
7/qX63Z6BnVPhIGTYqrtDaDZwE+1E0IUT5+iB8J1eOorv1on80JFlDVuuQSHgU4h
T/3ZJ8nC95iau7MGrKDvh0Rq/vVUfgu6xoLEWWf2G9DtfGbH6PzwSceDMVQsrt1V
4Rw732rrJz6ZOcIo04VeP0pR2i0foJIekE35rrx+OSl3hFSleHn5wj8enADyI+iy
0pyI0nAGVtE6G3rrioKS6eqweMUd4SDqFiJyzhPiWmrfAvJTRHGWrXYxliFV4jPJ
rnvVwjvHsLVIH8PShxM1OfW2GFEDpzaQeAnGuPMZsgvtkPDIgbnbfLa4Ib9dhuJK
dItlpUniTCk0Ju/35XmeBQEYOWN0PCn/fy59uHHqMsdmneWpi9dwbbo2uJb7WPl1
iw3DB2OK7ffgsVQ329WUxxo9J74lpCUTjeqMi6dPwb2S2EMJs2igAhKYRM/Q0bkt
8SgMUerI6fS1fRxKol47MSMIMAL5iLcYsnxcrHrtsWuyJ0NETbHn5zS8Qu/sKywe
5JIzxlNygug8J/zEYiAO7uGt/o5+Iy97OXbwwITZJiCmqY8jG4nh/BhKXPCBwfER
nkwXLY9A4h6t/nuSRZCQXHVy00ssXPGSbpC19qUa27dqEzL+cjWZ/F/1V1gM4Ox/
Qbf71443WReFlmhoQY+JWtoXyMOW9AxnOmyLe3Idv/2C5aKvUv8LLwQbaq7EsCuM
A0D5whdYDdv15UILc0OPRPPGrLv9rpQIiDUpREMxM2xVYGsTmxcWBhmaGDF+VRAO
NAAEHli9X/zXIWAz4opkvT3F5r37H/3oUX4H6qPPcyiE6x2g7Dwjc8xn7lD6uMJk
i+Z4RtRg/pwLG0OJTQ8hi3xuzWLAMhzjCU4zYJQl+41vQ4UXKcwZRY3IBDUxQ+2Y
dqlD631vdL198faOXFbk5g458QSqK9O77dJHhp+vQj7G6UTuYwYzM8A7D9KgJdgf
HqXf2BxK02wXCdVKUDS7jecrs+qtxaxgFh45wphJRYkxuBu8DX6YC5fMpmMpLB2g
CE2Igdnm/LeoqRrRGu5Wbq0pc83IWXl6mkFJDSJ4oDZ6c7jt6KRkvYdhZGU5K0CT
WjhHuUCaKpATPv6tUOoyREaYFckcrMxmCdWZxLe7sej+X2ZKoxc5/4H5h+4IFnqs
iaLUHLWu8PIHgRrPVvdS78xdXuU9QfIZcCclwTmUIMHxnfqswdO1JOI8767aa6JD
0JSiUN1FSWcM8hAIYL5XvSiUtpTcphfmJmleKp9Z9EF/ZSj4mbgUlAmPnH0BtYR3
NbtyGwL7jhfUNgFshN6UJRHkQCW6ND07k1x5cMWGe07TY2q2tOQ9cGGvhevg8zHz
YWpecQKw8fKedbTDTqhF+ClFv4W2I3p3t5XXX4A3Q2rvrFsMi03DCWK1oX3iM641
dVpkgBYK99TLumGF6mQGRPMMXg8N+hdX5/k4FBwqLk2d/i+YJoi/q+A+RiRruMMK
oVB/TUNlQOs2kPb913mE2vhTBGqfXKi9ssXGzI1r/oo/nSp24zrDmpDEK+PIPk9v
9gbj6lRHbKFnRuj9pP9dbLsgnE33KKaJt2iix55ItJQ+kAbC0Lh3xXym21h3rkJk
yE09fqA2bIOls2rvke7ct0oVQgf89aGiZN1+YVhVh6m4AUeYxeNnJc5iw5KkSEmz
v9mJt7LI0SYzhFnt4M2dHFbDF2QqkTGfP2qvhm6kc+HieCrbeAGQWg1B57kZv3z2
+jc85Zx+N9nUc5YXTl8pbdqg28P1B5uXtcPSxBR/7MTq6jXD3iQzfovTgDFRHkT0
UE8+Kh8mod6BaQWjwu3W31qJVhQkAGo16N6rGvYCYIFDZ2dO6W65H2qRx/XZGzCJ
Sodu3Rs05ClNBeaWpCyVtTrtSfUXyS+vezCYxYPmLcxzXRvDTmkZeNQf8GDd55VL
zEGypJZDD5uy/lunSk8R5M8YnvvKLpGHX4KTf2zZu16LesDW9z7N19ikMIB1nP0X
DIM/9b6tuZ0wpJNxREc16W57YwVB/7hdUW6zkyYzWae4wVIBbEU6i2FXjuAFo622
eTYkOu5eaaCQrWS87CA48umNS8yW/3yJ/U9L656fiGl56/XVbzxbv+TQkjfjz5ka
FD2ceekGyBykNM6OQ8RexF1AzX1VCIzOvPUppHyX/yw3zyM20YBXOxRkPceJqiuM
v3M0kfcgCbI6Awwvc+um5mCCO32E93tBFfzTIx3rwqTmLvTXD8PlNKLnl1FVTAna
A4J4WeDAic758Z1yTEAFMUO/RDI89MWFsB/qab+3pZQsYZqw2xWCX3RarqH7jIHj
n+ELbqVLoQNt6cJoFdnt+4Ej/hRd9F/Q5ZUMh7TtLumQQRGJP/l0G1hv035q00Fo
bN20qZWJYY9aPkxOyzZlbY6YKjLkkQRj9Kmsr1HOdezwo6jdVol7DIxqoJT5Mrby
v5i8Biz0HL7eLHa1PfX/GT2AeZhJJsTm4Vv3NtsiFzBeHto0koK1Xh9sWKy062xH
Y0jxdmrTFSkfoXpppnf/iqRGsHeWBZMvPVar58SYREouHwN4r/IoJkGd639fY5zp
BX9f7sIpwE8WFMtaMDxfQ/MgLMoYQTM1Wk5YnBC1MUr5nTcYyozprtCjxxSgFGlg
ANPZgoiCqBkGmwgw9jRa2hCNe9feeIPQvNqtLHFMh8oPjUZy7FMwcTRvt+9BkB1A
dkAA5riTBGOgj2UdXGmCrwfux9Xev3JWF9c8OlUsebEVPaQAdG+osRK1+gxlWGgP
/usnXxtdadVFA6bwXA7PpeqOa0dXeoQ5zpbk9MlBiMk1xo/ekOeEe95F03kKg64K
3rCCnWaZo0cWX6wS2alPo9i2sTMoLP/I8HZfSPjllpsLdJVsGn2OFn/CNBcOkYhK
FY4czCIvg6Kz5MS47jTLHtR0nG85mbA8BcoCnE0q1BLvGr8zf6HtEeqXyRjMyacA
E7YGK3rKnQYYzVlIbfCN8Vjuk0i+h5zdRIXC2VpJOq0cMDQAvzMLPuh1n7bLHrIu
/6/jGLxq6QhrXXR81C6FVFuMq1UiaTKiOXAgSVVVl0a1dlXh2UW3X7qSVxFSFcrg
ATLMHxPOdAURmIh/dI4DWoXHVbNGI/3if3+c16WzMQdaCadVvWTyqABEFplpTWCt
fWF8V8r9J4ChKG0TXkPd4KAC1lKQ9muUFiMcS8KCFvFvlOAt3+uWGTZAAVsYgIAq
c1s4vKvNTpE8YYohyPvWe+57A3T/bVqHSNrE3+1MlmyxovuU9pmGb79iEEbZ9lzC
Nkh/c4oJxCHzyGcY7bO1tA51rMsX55YX9k/vOrDtcIcIociArGxZE3s8XqkU4KVE
edFa4KlwpjInOurMKPCfTLYs/N1fhUOQCevWrrAVmqL3gJfc8hdk7hgsf6+R02cx
AKiw9tGJy/P7APfLl+FksbmoSPsGWI9OAKUFdP0QdDVDMwb+Sohcvz4iekfU0MqH
ih01PKwQpWdd+mpCQERuuv7Tf7Wx+ofX8C9ba9ZdAqJ0KQuZoA+Cuog3dOo8iicK
QGZNL1Bne+f5S9lbeSCkjs42jxb02VvFrfvWP2uETe2Ws98APiSCHRix/T6cSCC5
3HgmP3+Bc4YSh0xdDVh5meM8Mfopkv+CtYUhB5LaWpFhrBuZgJijAhIqHpwgM1q1
JRQKAm0QDp2iYiD+l2KXIf8g60PYW5b9jjBvfJIO8I6oa39wNAHPqk1HohNUh2Dz
7FyGkVwjvqAXEmpASJuimXS8TStzd9SvsvpOLEuDL/0d3eVRmAZleBjWhviVnieF
G8hXCru2+qhzmWyZDoJ7OWyEqcMsu3Ftpz5xf48g1xns2RSlDNMRAMOHvCNn3Kjm
Mdp2GR/xZlMtkiEZpcRVwxLNUGbemQ1auAXruX9HoKshhgqj2EtXYP0oLAtSLgTj
VAtLdCWPfACSxOE7ej9MKN64cqbTpQ62bz7QmIUzUFSmwQC3cOaYYAr2FT+DsZkf
xIlIgEBicl5EpuML6k+VHJV0ppW5NybG4dSzOHsYCOhJ354bka3P/RCSXUFfd6Do
EXVGvTw3hEsZMo0hDWAIGUL+0CTk/aOnUd3JQjYD5QJl02Ye1c0FuUm4JenxhLbZ
B4EHETDfSg8Rm52lXqhju4vjOcUdPg3PCEBni8YiaD0Q4g3Bpx1tSi5yhQn80cBp
6q3+4YE9pmCBxHO4FNGF0CvSEh/Pyaj7Hu9CO3GOWpynCmAHWwvYvzvBaYH3Jbum
S8pQN6aDJ2/AY3UplyTBCRtbVBiDWWCbOWYGLSPnLJDZ03j8m6Uno7HcgOA5Hjhm
I6Gyc9sRrWztjKBBxsf/p9dnbMLW3q37ldNf120m66IlERYaIPavddIOjVXdp1El
KDQYlf0YCRxY0vHFKk4o5ndlMh+GrUY7DH8na/Ympxdki8PWgdUgApVNy0NvZX8V
t9F80bTxy9hpf2Hn+rg7BwPCrOm4wgi5qVi6YTjCefCHMH43nBeL+V7v833rnjNJ
u+Q0NlW2p0rz92XWuM2H4Ei32ayXHitAff1Kk24w88aueN62ah0NFrHNO1D46KIF
tlAOcHA1r2tbFLK3CrpSHTN/56Il/AvdS963jAkz3AV9qITfqslODvdGPEAZK0vs
IGil4NcUfEqzGwr6b2bNTxbc7guUaBZgDSbzFqoSh8ZKkRrogkWfXSKJEHDw19zj
pDSWyMW097iaurWdJkudEQkfVZLLrw8L8En9beEOd1l+PboVYTGM3K5ezAnwQuJL
eoNnoDpUXrJ8Y+r2ui+dsCL/YGsZYBNbYkdnMl5Zx6tF4jVZTarFEopeJYZpT6gp
Zo/1xLkgQC9wC6E2J1xervLkeY9sZFiK126Iogs0gQIQEba607wT9piqB8svywtc
QHnJiyV6NAKge5K0rpz5Qjx0EHT7HTS/b1Yi46jYaz8abCDNPCMuVMTjvIHDJd9d
ffYr1aJrJZtozI1Rp8cn4na4wPqld7OuGhtf+GO13b6FhmEhg16gozsQXOJ+1d4A
0h7Tn0O8Ao9GO8bkwRLKEY6X3IqqmCwfjOs4RiS4kBvbIUu1P94mzOYH0ryEEzHe
FYIpZVd/uOrWYeyAHA5hi6U98oQ1HbZLqaQi7O+y6nnTgPiJ0RWuAHwvZzsQzn1X
fKppVrWdEbpy557HrgNgZKGAxd3sPgtgPSuKdS2QFl/ouTbaVoqAWGybotyu1qY7
t5pBZ5VOBIS9ui2kq6UAJ/f39sv2kMP+TgLwbPzlnx+OJ/KGvKKxPESCfV/kiw2c
u27cX9TD0Bc9qkS8DYD8z8BZ1NymLQiSXy2KyhO1RlI82sRXom6+KDwiOF6m0nw/
TK07zcXGrlqLCdWhZ4WuJxCzuhC8OyZsOu+d8cokxF3joEuofkGlqo+z2jZmEZ+M
b7u9sJg6mr2IKSj4jI6o6nUAhygPeC7/3jECqRQ09h24OTqU10bK34O+esvWvk7A
ET0owJy9snubAZEh7MREJjwLL/7YkudToYp/uPp/BfWfP4/jaYmYvZyO1ok7OPFf
IHXx9fFXxded2iE0uhO1vHZS/wMWcgAaBUnHEvSTY7AAuvtLMKuDsQCTM7ol6YQZ
QFiXwgqOOKkfuKU5jSZM8ezkDKOmjXbQCo4c8XADWevRo7Z65ezZEulTxAQPK1W2
b09JL4LanP0/qHmkQn4Zva/oXnqqEDRibaZu9OfxRwrn/9auuGsW4MiCl4Byfgp7
yNBoA7CnTcwMMZ3dvz9t/fw6Ig5YmtNwe2QUonv3co7MWHepTh9KBqPTJSK9xKnX
uV/0PukQdhrf3gNtlOmZt1I94eLQZD8t1IkrGQMeaDFy+gpXIxx3aBMlsqyTQ1IH
7nrLwNUtFmxY1Pd/pfVbLYmBqXRtChAJuXqVVbvxPCrtpKw6KKIRcw/O2QjhPT/M
oE3H9gaFuy6hnPozHR3OuLLb65H0nQMIHfLhyFdWqVpktk6YY2rqfUDQu1l8g3Zn
zFYm6XW+UA6MGtgcK+nd6+BfqcyF7Ic3S3Mn+fJ548CeJzcACXaSELo9GiFQuatG
V0DDg+4v3wZTvaa1+CvfnmbBB2MdV7KdAOly/thRSVN4y708RkXU8OzdzPLmm9/6
/eYwIyA2XUS2MnvleHn2kanyZCeTL+cHi3s9olUP4ECD90JLhjg6XqYIU5uVzh02
kNfmdavqNdnaLhiKqm9oaDEjAckDTvTLPv3YYXNxtX8vrUw1npnLRv/1K5Bb2td5
P4g74mf8fIuheGhrtIyQfv+jBzAEWGXbrx85H40H3FdDXf+r9PlRp9UB6+okkgTv
VeB3xV2+TBdVIQgImdVvFh+8mg0+3aGpClm6DPfz1Z7XZ+oN7BGd5K2x4q4ukfjL
7DRuGv22vCrxqv7frEL4RDkGNpP2oCfS6OmpSdMgzH3K2BF64F9dG60OdsK8IDhG
DCHDZ9+PSquBk8cER2JcoPndEMkZqXqXQ/q/nXOolld2cRVrblJSG/Kkn6ONEUp0
gZvdwyr4709QEVWGSk1m5d8VcL1Gro60lcTVXiOmWS5Z5AknIXB9+tsUyKItNW/K
sTR2klVWcxlJUqoXwVMABdhHfv0q4MWnH/9/gY7zSKk/73auKB7dKtO3ffLwTXFp
ioTb4nPOvmH8TuiS8wAA5jtnlKRTtGc04xi4kT9/TM71xkrzJBbH1zNBlfYdYb3e
TVsMTLu8vkG0dFBqD6hekd8HT9CKBhwqcX7MIOtieoZsskgo9ZZpvKKeCg+zmRD7
lovnBAUpxkDof//wkCeXYfhxXScKSa4ScF31LbKbWYhvXg+HU0zFeVEBT6/TYPLo
jzbz92lZlKGTt5qGy3wsw71lySPKlV1CTbjfMgcO7GHTKn/EP0y5Fq6EUmDsNgLa
0Cjp21g4oGcf6HZor97cIeJRJy8BlRdtMEf4sJhktqbURy0mILXljV7eNhiYteSi
aRqn0B9DAAkPZuPq6kLWLoB2uvUL99KvTjCd88GSHbir5i242qsK9hrH3i3y1+Mx
wmDCpfujIBZnJ0ZZIR/BmiT8cUh5+4kotaMaA2bn2u9IKV6JMNGxi9aWYapKoc6M
tblU50+TcadUIZ4LWzKvaE7MMNY+gDoiH+0PuiqdMyKnEvwhNPKXcqj6mjU7jgTW
R7ILHtQpTVD5R5fMCNDJqRkW7H1X4hW6KZFIkMrS1dWX+Yi0fHS9uEJH580QQVUr
X9uJ/gzw4KLhPZD7xxFrzEd0E3Vf4FzrC1AYfyvvGRjdE6fWxx9Md0MM7Hfujl/V
4qYGf8hSxWrKFlb6i3dn3XTZM2Fph6g4Mazxr1OY+sXhJET3XdW0EUQZ/BnmJBAh
eU7C0Jyz1h7Jvy6eGX55sA2TFsDPzZcJHQ0ViPYU5ljDJQgsw4Fe5IPT1oGS8s3W
GGkRAo0owHJmJNoqCAPByigIkp7dMeIxkbCZQUXSM14tqidB+lcOBcnmXnz895Wi
qwcCkG6HXX5wUObU8N+87tuH9CtYuiEQ6NRzURjCVVjOobHLDmhXCkPPkf1EJbEB
hSxTrL5hAm7DpOCDVcZEyLQWfUEjuwDALLCPGTJ2mQeih6nlTXN2Bi4pyxGkHRI6
Gycr81NuxVnoG5B8MVFxUfYfBr+9zp82XGMPyAGjceknrWOb8veKwuXkyqnnFjE8
nMZASX4VsxEQ8e/ncbviQnl0vLa5JS53+TcaMV5KOfquGwbU6TcX1+mme2oQ0l19
F/fVAzQsQRVmSyb4y4QtGZ8OtgF7XFwloSNBLm1Y2zpaezo+4hnm9WX1fEJRnj5x
nFe9dXfT9Dl44kITTRFr03IieNSV74h5V7yVJ4UKxSpN/JNDpr+QllJaALGfMncS
6E9kLRggCvxRSaDjzdAtzkPTZ25LwP4HEAu8SUQfuEf/g2ZMCXGGm0NgxS3hKpbd
nf7j/9Bs6GBzva0Mdl35FwhLdaCsmwElw5jcw1XLSA/p/LlPupqAkz3NPMPqDqIB
QDLk0ygO4u1qx8TpKcdOej4XZL6e8SWczub4569PJOL79/nNLAN8Xymg6KmggnBx
a9zegMBghdlRca1dK9PBPnJascdgfsMO4P4ATFHqmKNqTEn4ajSDGfwRZfb+jmoo
mnDDxZxYfS5CUIN+XQUpUDsUdVX0kRU2t0E2Bqyrv5OW6zgqL+efFDgdj0BSQCYV
5UpSnzh4NRCilHf6EZ+nn2lHlH0JYOFPqjtO2Yki9TvvKh/YyYaVjOwdy44GWFdz
vMXMNlVRIPhabt37xiZJgDaJnKIOv5zEU0kLvGrTXXmUyE9tE68E3fWS37J4hw/6
5RoSNCA0fKbVVhC4d0gfCDaukwohIDDGa0z2jgoQh2ozywDXkF2bBDHdcYMdytHH
b36VRn2xoDR6IL4li/BSJoo3pByi29wLWW1+afMus9QME1qcjYn5krAdtCj2D3at
c5AiYOGOSFNNEkeMDPxEkxOXy7FfY73L83b1Ms2PkxQ0kvTgpna+duE+oDdC7EvG
JobUZd/iOUPbSEgk290d+pYrDPMpKXsFgusXG3Ss56o1BE74ZNZ8Hfsr33u5674I
F53lmgc0giziEMmp8wFTF5D1r+6/frXsDYzHauAej4pcoLgOCgqos+XW3jubpDcL
s1l5UctYC4g80EtDGzHiV2pNKDsDg2Spr8CmJxSAZq/7jaU1M/ZedrGnUmMhIazA
fis4d1zuCvTQZozBEbw6Fol4jcDqGPSp7yU6xgH+iJ8CTeiQUsyCzaGk2JYpD+kU
Ws3YHOda14anblNUleVBSHOk7rUSYlQj4wOq7tVs97bHvIU+du6MuJBHYJljFKBu
HvBq2YMZfXzA2ti9eDUQO3pVTemzTt1ybKnSDvIUXDZZK960PTn5XGcT5dnlFrsV
s2CjJw0Us/CUsRB/xLsH8P/4S2CCxyelx98nD6FcxAXWuybQpx570xycQiNcVaoI
K5jW/ciw2Cm8JtMg0Q4z4Nu9b4zc1bs1IgFb9KRcqL1nnshZVtH9Uh9N08/uVMtJ
8XzgPHXMVPUBfC7TEcULv+wrWw9GtcnNMOz3C71Llt08mOr1lvVSrs7Zyvxhuk5g
A4p0qIW1v/HxF5wyCXKtnE4AjOmK8POnhb6vzYUyqJjBdjZeoZlTv7TmRXQq/2EZ
4oqLcgzvxxXTdnFmdBXLDSr1LxIFGWIn0YBvalciyRIpUsfgk8Hvv41sbs6LOGvQ
rKFNqiK27AXGkBbItBbqbDofWperTaIE695tpiFW2oNK0lR5MN3Nx4a1v79KDMFV
f1X3yNVadPYswxIgoOH3EDQcsRcJbjkRl/4FpQGtSThersC4dbeNYXHwfGnJ7cAD
PsSTF4WeRFEJGB5n0Ac4kgAD6nlbQvBYyI7MP0/vNKOmtw1Ivo2tJvKkjNE9EXMb
2Zu13XyTOZlvsCkbNwx3Mug38kV878acb6W+2ODqS+suoU25ScwBXv8tScB32h4x
jWChVng9o14Fr30rcP8GACf5HFTedjKzxM95O5U19JXJYIeJAMkKcVhr5kuprZDM
xXKRpnuYywLjbj7EffSw2tx2X7ecRtJXSA6uuBY/gK+rGOkzr/YqpeJoLk7/vz96
Ai/22z0pnZ6rZLVknmOS57dmwLrHfC+aG21LDNeD9J14vrspR4Fb0nasKaYGZkta
Vc3KayH3hOB+JBJxMJVhK/x6eO02VrNQjtesWYHmHFknqGVKRwlnAjLXu9FUazUj
oxd5d597lpjGHh3/q2UZANdfkBJkMTc6gf1FfHm1FgtS7Aalq5Elx0sX+AA5Cdv2
eJfJaLsc154TwegpqiN6FSakopFzqji3jWrNJoDyhwtTNiNbbruw2bQ2BoUD9Igc
sax62osQzSq2V3AVw1ENGcicxDosHERbNxcEH4PtjM3vSeE63k9dfZnW0qxQy3mv
bWgNeLwysnSPgQo2NPdGVqDheVHGzTt7JGpiLgeJt2IIh8En0bU/zZ/XIDMDWBgK
ALvRpBdH+JbdflT9ERTDL/F/N1shayE/925jnthLkeCgLKaAicd5NWfJkS8m/Cl2
OBJMBjckV0hzebC4VdX3LUw2zjhogluYah8qec7+RbhmdX3hheOV4PdAyq8DwlTv
B4g7ufFwD4jsm60B6ha8paFowlsbgNu+VqEmha/y7c7hXcjBpLUcvqrtR69Rkceq
59RYr+Wp3HpaYbxR2eaeEuvbXQUkWhTaHvJqkLHbPjdKcgVPqREHSiahhJ35DCLW
0bLO1y8DOb4HFp5PUddiWtvl8GNryp3S5RbeiSjTnD1CFqKmQeOkPQ8EuEzDTWd2
/KN4iZXCpBFhfOZck03WcDC+3JJYpoo135GJbjn+QHFTCYUxj7/P63sVGcHNj7hS
+TqoxOukc0FW4epMfnIgyOkGb0y62/OPr03w+Nh0E7dPN+XBVWMx52egna8jsiBy
UOg5XlIjqLJpX4lw6I8dRtWNQaklLxVHA5tpKdb41/Fqm9kND/uRguY1LdeOw/v1
NVIBy/g2htdkPUK7SpSIKDLKyeAKB9piHieMwok7COc6cWP8Q+JRUJ2DKZyQ6k9R
iDUuwN7yBc+NxuxUWUyI8WVhrOc6Mfgps/ADGUsgWNLWYc64SKpNabpZA9ej78eT
QuCk0l9Sn2y2KZuTzhuRWE4dxqm6Ao9S7JNA46yGtX8PlGpU9c6fViTbONqwqnZf
xjzkmhyfvsoq9yaemo+OFdHZ6pkBadaPpkcCV64j+R40mU0Ojir/yWj+//MwDnKn
b9LaVHDfEnAxOcq3t91E81V0Ko84D9mCjZc7UsimavCOVN65WQGkctPeteIp3qOJ
Exqt0JUls/PPSbHGKyg4I/nlXKy7iRrMiLdVF7aygFa5FWMmyCDzxGadkFVYzt8B
4dzTlYRGliQ/JsYeU9D70VrEG1hhbW6BTnMjWhLGRdMcmwnjGFCy5WOFGCKzt95o
lFiPubjOw4euS7SKvJ6Ouu+QFKL7eE0coOg+vNdmkEZc1hF43UdmFLD+zc3EMSaH
J9xaZd6+sPnb+cTa3gh5Cl2K2H4qRsv6z3Co42eVQ4vG+SNIiqeM94Qxzxr0Zzow
SbvejdmiSPiGONU9gugsiRqqI8uYOmmlN4k2bPvzbbOMMCEYlZygbeUyXu+CP+wl
kW/zxN4OGyXEfeniPYIlYsOivJVLtiPB4yP+sJtifaIlvKf9TAEfPQjVFWtUe3Jb
MaTxSgdspk/vxFDw0cE1rFKgo+B4YD0ji/GRHHXiafQfyoWxtSsxazMUMJj10fac
5k0ctmgdftN2nnAOIzUWXkkRYXykGnc807J+3UUouD/qlumrx5hBEA8he5F5c1xX
9EI0NTM19IC3Tokz0BifkfwCN4t7ZdkiRT2lQqFWUqCK7gue8v53vj0KAMIJOE2L
0GaI59HUGDF4g67CStHEFKFx9wwfzCiKZTgnzpul6msSCLmWKGAT0Uktkc+q5dPS
IdARC0pshVluqIlpXOWFZ7qIVfx6XNu3c25UnYrCVNITqStgyIHwcZ+6FskiYhH+
oFfXaYa8ub3019bF5ROviEcEPxDsE+7BQZ0Q9BhkqrCnCiP14Dsf+l9CP3w2PkCz
jBWo+qNwG2oWG+iBxpqt/NDXjNqzfWpsVIuAXqRVA5nhMKJLJyhvf3KLhNtQrlqX
XcVh96IsDFdEfUpX39XDutOA1RTG2FiIcTrrZfAy7VeZOrbWTMpndsPcHVs8bkCJ
0Inczd4xBh8Xr2VLdVB9e1QnSwE6XPOcPIQ8YVV9y1Tp6kmu1dfBhPp+ghEZnl3N
i4Uu7BPn/hzYfnXYdadSi+Zchw5oMUZ2anNePC931udmHAqvXFUhJvxbCFgwUfQk
jOwFbVS3hqYak7UZ5uHOcs8pNF94dRUBwZqkPXsJeCggauumiXyKctc8s8U8IFbf
oNCU58lTIXMHHMQUdJiCNrjp75WieR1r20cJCOTu5WADq0sk5+BkAYLZANI6j0SU
DqDwTJjtInXHxbol99ijVxzRCdokEEq28gURc4dCbF+TZFFfwjt7jpj3geL3Z0kI
SmGe96sDIjLpU7fSjxn8ZYfe5xCTMCl/pzjCjogtsv6Op/9Rs5uX3dox6tB+cNT4
PoODsiFfRohhF1eHYvu5BNELWgp0CngK8hqoGep1w4Az/fhGe+Vg7Ahv5INKSvCn
sPxOw7VJ7c/B/jiBMun3awGN6UIPDr7Xe+Ik2c9Pc1CnviJK3LvK9MMf6xzDegUA
frMpZ8hxybsvMC6zDsBuujvYzgJrVtwTz7aiPKOQTVHXodjBZLRqGMsrYUC6d9re
Dfz8VIOXUlIjSMqAlYE9HGmHa7DpshpAzpHoXBUcmc/FrXzNdt0COlOCXeCM6RiD
lm49ou0ekEclaksLLUvydL5tQ4gVQ+YSsLB7OnSJHtJISmSYoj1xp3gTfcy41WqA
CjiXkh+VxchblyyoT7Jou6jUgkQK1WPUUUyC7r00u/eiRyZNW04ZHGPXaE7RQDYT
Ghm3VsiRmN5/3IyekZ78BwLgr6/AUsaGwXRE2dmYan4Vmm/iZP2iYNXGgk6I9Jqd
vVekoFZk+y6ztMf9UyrdMVtBezxrQubOw73MdoUu3sJJ9VOACwPwdIICkGyGEtAI
FbeukmzWEGnw0BPI6GnT6Yv1X15TqI1mPRLtbfFyZvcPLdWARpuiBZwH8OiXB0UU
t4fh+sRA/abouaWFtvMa48S9ieQWNYwmQvC+bV7KK2QrmxiXKmHtyT0mL6i/HFgD
z1N7KveVshKjKQHGc5U7c4LI3aOllymePSKASFk+1K/rClfwEvCHF0ehahh1vpfl
TkcrWEmqeBQw3ZM1C5dBlIfPYlVhBM6KlXye0fV7uNDVOTCZ5jpjt6KnBFFUAXzh
7wwYObgEIK36VdfmzOhhx5pYP7mS6IbjvJmCcQo9f6xCCswJ4SQWeUi0bhkgTfo3
MozJlKxu9lk3ST4FDu/c3xyFwHx/SD/Aq5VlyqDs4C+inUvR/1DBgq7M7ggaY8ek
ydl63+0PHa0bHlDp/HvQMzYO+UMFLcQuunCTRpKwkmv+viFCmy0Heiv0XEIe7R3v
SfQJvmOZzQwuXE3lbJn1htYJNeopKcjiX18EFkVYFvFUNanAkUqSI3juZ1flTJym
4MOEm+vCHH4cSPBHb6LTYGFDPjCcYczLWlMH6znLio5YiVxXbf8qoQ92uhwVKK29
jeFtvzhFRjIDwokwfSMqK+XzTU3zVzN5X5FGiSHsw76oeuTjX44O0iuk5rOiN1Ax
uNpqsBWS7CNRrUin2NVfpm0jK9GaCv/TIs/5q+cnKZdUvkkTM8p3DACvuUPPa6T8
VwXGxk7gE122RISS4gYlPXg7pxwAK3XExR2NuapjkvlirCBC9KF1ohYr8q8IAAIP
W+YslBLnhZn1gcT9lwObdFq19VU3pUkUGC7qrsDMFbf3V5/mBIyGVsy9GWnToGiM
eRTVbooJuifsmvM8mzZn1Bh6fSIX4ARABQbkHkr+O0FbdJLF5xgEtbtEAyHNBEqF
ChqfY79QYCnN5hAL9NqO0kg7i+ddW16yJGxIcdXER195yItUcYMGtlCzBNNdHf1t
Uz8Jf63E8B0lMh4/C6JEQSHKDcgPg6FYyG2ItRMlekuy8jRkaJP3I3TVHdHAlMgm
5kz2/RyA/o41kvk3CCQBFzAgBaMsB1YcvlVsnR0XJeRBrWH8eO2tWnNve1xS5gb1
3BFPCS+LdEL6gNxAyyz9FGHcqMhFv9N8z2UZtfBlt5XrDuuaEOzagB8nrOdgC0Cr
R27b/PDYwM8MzHNaKO3tbSaiPPMixuB7FSnieHmuEIFTrndPj/xuCpTUOscd0xXD
NcqjNc1vpNdrlPZHjkudEs5VqBi9nQLTyuEU8j0gYdEmc25ScCiw1f72rcvrMyWb
82j/2J1GgOA4o8iq8bUJrIeMe+nu7EJZKV5q48W81E5hsjWdn34pvEpj3/3t7sRN
HaDdje3bOGPQ7GsLoGeuiADinwHi0fTD7fuCsOvCbDlopgnGodOrQad2GcDoczKR
wRcj6cCzrQgFQmk5LusScn2rXesblDMiT68sRhdyxKZI62uxQa6s7h65xpuxHbAJ
XJR+zMJY9HOF08jvF0RXXNEhNWOJmmNAE7s8Nwnow0IQ/3ftEknkYKXU/swBexN2
IxQgfQS9Vkup2UBJwMXddizErrz4JMA2z2wF9xbLTO/vy2SbdOdUMOFp7CE3GX7x
pYsqfB7lQFiOIEoA163i38wbP4kjeWGHx1jjm/9VLEYNGTIPeGB5xrAWxTe58kr5
ciE7CvC3OzMrxZwEIkLNPyv39b0gvi+TH9CaV1cS0Q3ZTwPVbhD8Y4FdAmL4FXBT
ro8VPUlVy+MzxWgvVESU4Lcrktasm+KRDB0+zdyuHON3ud2GuKF20odo0rAcVIp/
mRTn4ReL1IBsRMGtzIjOxm0oqr2lTdgUgqi/hD8cyOI7NEoBB3I6AoHgvbS7exuM
dWNlLUHE6KwdsIPRCwhsoW7eyR4aYevLXY683SgVrME9dtuQciLQCD9nc8ei2tWD
oF2/jmGAsSWfx9wIVWrfsCZwfjHYojPaOesT3DOt+DTpMB91Rn2HYMteJzeZLXxs
2V0iTOrNhsAG+kTZ+Pkwx4PX1KpoInP1H+TmUi5Tnno+CUFj98CQHo4mHmbcN8aN
IQPRku1WjTcaOoCULGbRBq77ODOMdbg7Nyw9NwxpjwHva11F1y2v1oK1RtJiqrWi
HU90bbg3NWt1UbZV3JE3buy3iTSWa2pGxWUJhjdOS0g+uW8lAmU96g1f+FddQUXB
MOyt1bFat6gtQ/+dVpjVequ9PniURHuOxQYZgcG00XB+CaEeUJUeERRcBjnQ5HHu
pnaHFFZwbAFe373WrW8tUCIDFbXBNQETRtgJAN8prVJ71GxJPSIv3NRg8v1l5KJ6
z939SOnD1T5cjx+lwNg8kpI+GHcW6AC4g1r3x+nACyjBTRJYC+GrLBFjKy7Xsw1H
JnpIoyfg3eDEetvMkbeLXSRZdUzbQti3pL7W9rvqeGM+/hO/saNNunrrMfZtJ5wv
ewRCcE6m/mfVZpQHJBgvxk0xJWBI4gAQwRueWqm+tHcE39dwIU1WsuNsdI6DWaz9
wysqTdkv4jEeo47n8dYXBbBLJTgk/gHijTeVvTsZAnCw8F4dccTYagSfmOoWi0f7
yMGosjgGwd63RfIwgo/fNikZ0PlRHW7icLeFh3dwTfgheSHM18Mmk9LCfidSQDpa
1QnBXmlazT0G1ChmfeHcJ5hQG/m5Msxv3QbhzR+FeVSB+wk49Jz6vVJooUsJcmIb
QlJw6fiIg57YArm1fBOux2SK9AHMUJQNd+MbQ65Tjjefj+7kkvcquwCTnDjupEpj
f+gOszd0YuvlMu/AQ9oIrmYgkwJ/3YM/fhKrWTYxLRs4t1+C+u1XSRqtrMv3lFKZ
MySiMpFvOiaPjUccQS0UET/GJ9rUzLz6Zb8beqz4yZOIemaPGvPyvavLKa/+Z0vq
uQKZwmJ9GChDEmdfIrxPKbHoNm/XvlXMCIYYC21ACUQA+cxzDEQpT8DCzp7dm0ui
xB14Oxq5Qrd9bAkvtKLwN2uGGjytCfnto/r+tgd2nDD8BMEkOcqYc8A3/53cywnw
ntkk1mMm39FankRy87wONkG1VHyoE1FYt+mLFmm+lb+U/uiruu1vHGqUQLX+H5Vw
9w2jGcQSDUcbQrdS/kTBoA+gyZZuBo6vBuy3JZ1dVQVYZarDrAymura4UPMR5BqV
XHCR7JeiTEmZbuXu9Ya4LhCceJ8LTif+JBvXotCMZnvtpcWqfeqU7ydCitjVpomm
CQEjhIRXCHpAf44QvfuiNuOs6tBHfX/CbOiI8NZk7mTTZdNWrG4sX7yXpGpqJ7Mg
NgYcdI5Nx8/MprQBIRG7tfcCU2nauaWGeLZ7a+zLmVM0VfYOABkYqJZj7sgJiC6d
n5cKoPn6KPyElWPVVuyuyn+NM1kyF5qCGn1TgcKn5ySOkC/PBfN0zx+/7TvLCwgP
EFAvAGA/u/6DrIH30lgvwXCVOE9VC9eUc7/8hDKj0VPF7EGa/2C6tAw94Yg6rHJu
Q8bvTd50Vf1zpdVdv33BJLxF679O0EJG9NKXV8Nt8oCipWdchDUyHEPP5jJxXDf1
ADV7rPjLdoDkWuCs6r7c6iy6BtVBr3a5t7PVAHhqKBXqGq8n4fsydtiCI++biqcD
5Em8saDNoeziyBpuFZnR2Fvyj01ifL7BsFVbDJpDIO1VvoTi7sVPjgA+3DpzkfMd
eH5jYZkxqjmlhm90y1IxAdgXOwWJmDa+Hjo2Uqvb37dm1tYGMtA0JiQo/ctvdpmu
JzTG2C6h2x6CzPdsBCHBbAQTvjMewoby7QjLP+ja512Ahusfe7XJfX0VWIUQFNO+
3KBXrQ6VeCaqt6JTtTeBHdHPzaJJ7Yl6XVpYpbA6w0cFvRP4n18fxep/fw4YE0XG
+BPP1+GtQJx5Tl72aiLl5JSlCpm00O8CGr1k9SJ+vPxtQAvvBQkbJiBuh4BS3NEC
nlDKh2didjYE7lwKdwZ70gkQZXGzdS6WzzEL6c50ctO5ccU+oDZ9rUCILS23ZVwQ
QDmofDXJTH+nQ4vR0Uge9IUo3iHx7HXD/NxTjl8cXNzI5XWEooyY8KLI6v97KDCM
q/d3G/hDdaEOwifMZm4xWnbz/s1xANonJG2/ED1gFa1wNfkhL4cU4ObgneJCH1lD
dHbIt5ZNvNP+L/ukNgxWovnBsJFTZRkvVaFHVrhNfnBVOdU0LX8NHcGH1pkkwlPr
XNUkkux8WFsk5N+k1CZoRxb0dANplPfF6ILeOwoRl/zZkUNpWt9GIqkqPu8xcJsB
TOKuKYV6jzc/4EjyFiSgIsckygi4c18gatAOwRN0uIoUBO3z//uGC6QJvSe7xguw
cGcZeF5EFRjLUFZNJOGiHLZ5a08EoVrevPRPDT551VXBG96hLy6gZNItpoy5wNCz
Izr8WI5KGSoMPjgD1vvMRlnkSxXK882PZeIz4VwsbXOD/1xYiHYpADwKdR3JlWld
O5OcbcJsd38Zn+w3wDQqYqubnYpvo7lRq7sMF75NYItja0i79mC3c3OuxIUFe6CQ
JtOHnvG2Nn44/ek7rY0hLQ3KZcLjpVCTccGgNhDoE9KEyGgd7ObLqPENtqrSCFIZ
25sCr0XcXR2MeAf8fTO/7dgSyw3ILg9YIxJpeZsKqfZwdhTcgH1KGvJT7bGHcEBK
o6y/H4oC68TwNienxe+lbDI/9AoxBI0hGYjfZICQoHNsJiKP7hSkf32617qx4NV/
fKMec+N5gPJkZChxRQU7Q2UHWanMyLtQBWCVGs67wZTVVHFMfcNddhEjncIjbRqe
zCoXdT1rijmlGl2z1XDRuLot4E3+uftLb5I/P9o7dXLX543YkwSlSnPOFtmL5D8f
Hd8DVFCHg7YxuL3rxoaVobulHnISnLo9sYoUTmhXMsw29oQ8msDIAV+yvDQh5HIR
WSAeCsa++uTCejQYJnP9lxiyizK960pSVjA8eXtRt5rSd6gmH4lInnBWq+RDAMt2
QnjxMF1x8yTnpTj56rd0LTLrbQCQdzM/j0KnHP0hN4fNe5I/q2whZ5SDwyRRJHUo
CY9aBD2FxKQAPKrB5AIk2KiV97i8X2mt8VlhEoMpWmNut49NQTjZOhGF5WU0nuev
kvNeKH9gKB+WmsytjSLi7Hru7SoGkchn/6vIOgQw831GhgGMDYI0mGSm2MzWbsYp
mPixGlLTSbqM5Tu02h4rA62TriT/tmibWC2OxgVSeakw1sEb5i9rk04i+rajJmgG
LKDu4QH8osZ+j5GUCVh7veMVHYOgVIn3xmkx9fjEP3EHcWC0uS8dosd03JDMxLqe
uraXFN3sccTHwYcwMWEyWHhbNNVOU96+kPHpNV5J/SkOfYnDLDwDP0lupWSKqoCW
UixD5lyjXa8u8d+wHKjxodGcXARCNS8NyQ9X5J6URvZeX9Sb0+JSK32wuJACQZ0H
SI/BfLu4TqS3YaYiLXX9W3BcAUdCVvr3484Hur/681ggJzfUc7X0Ad2w9rO6wqB3
DDBOHGu5LnETyYDLK9x66TWJR6VgZkKhI2FkiRJzZOGd2y71B7vhUPgbteDL8FM7
LhTF2BxnuZ5QfMCng9Ad+k4HVnbqu4y0JRVtjULZumld+bT0EMX8z36DL6Pn46Xo
RhGrgs9zpnaRSPGTZlUwQxHt+HHi4m4HA5lqHxLjg8cblYjr1EXy2m+baMybQlEs
wxeVDu5Pv1ADQzs+hCcPun5uGL9+76AXx5kiqgDhN9+F3Pg/g9zJ4da2rennjFYp
085XAQfQQ235wMLfmPqp1w3W/4voGl30zGc3lUQ/GKoX8lZrKyE/pUUrvyS0T16t
0B+aXECTtYkS5M6TWDbsoHEd0DfJam/Q0p2ZaEMQgPjScypGuonBZVoH8JnpJfMs
hG3xjZb2pKakoyn6S6uCyf6leiFONy2+hK4ygtonmDJPc2nrWMoiaDeTGi/71w0i
jzcCn49p5XsQBwTAvGYX3jDGYWFDpl25cNRGvb5Lm4NxKA1e+2x7uuw+Er97uiKZ
4zNzqFbyHL7iYRJJZ+G7utI3jR6HmxY7aKjTgvsI1vca5C1Ff96cu3RyO/Bov0XZ
HcqImUX29uDxk9VAM/ZuW3HEJ8zgiikGYQeOmWpyr1aibTG0fkl0Nzl2Aq4Nu/OT
eFyfHyOECLHtDOdC4loLD00Wo6dLLVmge5tM6r7CObz32aj63LGaBneW2mTim3e7
4XoY9ecn1Z/EX/LLImeq5nD3ktuZQuSXBeLhAGSpcz3ydfH1hySLym50ceTKf1g1
fUCbzVNAZGW8t73n5Cl8XPLU2csNtLSrMaPx4we3AULKBrNQ7eBVdJ7pg8sH6W9D
hP44C7uNTfAQdh9Vj5+2mJjKbrnFxt/KeyGXsIbfXyPnr6KecM7NCqGT7VM/wRaa
HTY12sR7AFdNbWjf1y20zuKvUrN6hoJeBVBbruOblQh6ZaNKTQPgxuGMlnXqB1hv
KSznGMWz1xzeQqoAS0FJY1X8u6Ir49Z2hwWSQcC6jDeQnacvaIAioTe8NQmeeJgN
pxZWv74pJAXfC1+fIr+EjbG8wpg2j1zJC9eRxvuJ0OAXVSBOZmPA7Pcl3SLkv695
sDmQP9lAYdiMceBXUr1IKRYp9vxH8oHUqieC18TakK1jaYrGMIgWpUTZtvOq2wnj
5sfFV41GCgdYWovNPwuajWHJL1E/SDe7NDSMARZiZhBMznIykuhAA8m6nlOd1uo6
RKypXOgTw7cdJvWaLQFw1FPxoNuliagUYtIMSUYN+yPdwLZ/IU61GHLU30NhA6mo
w+/IwLe+IqQjYJKtoF1t6VMOIeF6TSfJS/qIJUyoCzLtdR5I3q2M2qlrE10XU2jW
/UkXxBdUkLhB+mSKhEGLczM4yya+/vJvi4qEX4TNtjiApABwhoVWrizD/Eh2WOBc
sVxZFXwppmKDQEhNfTKpsGiFLo2O0bwNd5Hs/D+JK6XoawkxNCylGU9T2UKGadcF
4X75GChVR0969jUsMu7Se7qECSdb+Xa/0DAdPm3VQ3tbbiLSKvkLAP6MzWScGsdV
U5u98vLxxHWByNCgNQdjL1UhyRZp2ot9yQukR4s19RlUJ1qvpGQkkDnkeuqfeiEo
R86ZQZ7Q2cokSHizQI2UzEUjY5KaNLFRtM9KDvu1b10WTC7CV8uRgDnlUy3jNzos
MDqxxR34cqSIi7I18mVV2FHxH16QQWavnBtnU6Acj4OEJP7KXMs8ZaHLjQzl0yis
WEbvua4l9j03vvGkfojxGzMvIO0wlgnjwm7CaAB+RhnJu9jPZw+JS5XRcRzQox1t
zysLixw+lY8Nxpsg6DXXlLCsSpKe+3qb6RQ4HtXiL9cEF7uK4DlAryPIUQrp2S+6
4Ennfv1MR8SZ5rfv8f3aNbxqJFwulKileg0kLvVD1wsKwKoQAhuPw3yo2IJnFqvK
VHq0wGPgT5Qa38XDXANzLUuVrOyq6LO0qmw+Eluqn/0AsqtIL5Mko3LENFeAtj7Y
skfx92rbkFSuDFmCKnk/WQ7/Ro7bU+k2VWZ8WbDdS53KvNsJfoDd1OfG/S8o5NIB
fX60fpn6QJ2h3IzVBwN8bAFycAPNjBEHN/i4XyKX9YVcwEhTLG8n7mJY23dfdpU8
LrDXtyF5bBwhYaqG477MDtAH2Zm8dRbeqwSCR12BsJP1KCV711dffSf2Fm+gbPFX
uZ87AgqfhsggtFcL13Bj58UjXt6t9/H4H21Q7/fc13xrY+WU8op2VRwE6FljPbiN
WrjQ7at1X5L5Pe2otofZeDIZzWwxyeaN1oWB/fWF0UpX/KA3H7HSyS+H5Q+jiArC
4cv3tSpPjN7DFTn0F1joSUDcSPm9Pafs6+qwjMUeneOxYtbydg4Do8hSHyObDUQA
w2JPPxUVl72n8Jsmb3bxH2VrWWxWADb0UPPd1NPSOgg9S6cjQXhswS4gPgQpJ1iS
ZRnhQga+WH5uYJzhnMX2Djc6xYOxeCTINRUUaxFBg37C20WhJv76MjJxPnzcOl3J
4cmbkQBE/eAMpulpJv3SecYdoVakhJ9iy7wLEhU6MVA31h0+eX6xf/Ktd1gZ62eD
DT1bqdsUK5pDQZOwhnm/U2hAHfSCOHoIPLEXuxtQBnRHyKiVDlHz+Eki70NLmlbI
k6VawrhTYQkyu1RjzF/vaDa+V3O+Yf7nZrFWBH7h1roFn9wEUzXyujLt9n/S+9dF
PwhxUMBHioacS24qfmimCA/3RMXv33gTUNp/Im4BaJs30DebahrLoQaGsLIUIU92
JgVoHthFZ6DKHGhQLy1sZWyF5hhy/0FD857FpnIUuobgcDdVtx8lptuai3StECc3
yXN9NP5NR5Bk21qE4pESvXA9H0xK15eeOrenjHv9A3SmGnfJ9RBn67ITJccGTOwr
fwHoDXdnWMyrOgr+B7t4r32iDjt1XNKncN3YvcY1ej1qM+lGh1UBRT8qS2KIfa/b
GizrjJqfDnn548I6NWLq5BdGT4epQOXsPkEUrYnGq8e3RBEw2COWJdD5y//4phF3
JABBVMKeY9Mi9iJzs1vcBiu2Ngo8q1oeUKJLdMMY51S6VrSqU2LUZ7sIEnvfhyvS
cPqTQ4gNk0oxJHBz+kBMKgacbDdfX7suutFvwFuUK0yg26AUy1nNnNa59RQhYlyN
toc+aH/1r0GL9mTTyZfSEmmSt2Qb/124Pp2qBUvJjWPo1aFFLLVY2r+IpqCTxdeS
WHBdvygGCHoGclH8WlB2yqFYOM3NKeL2+6qPzU9e3KARePJi7/oYmk+Cfdd29yua
/huCM+Ti+nxansfrKhhqqYYs63hFnepVo2oLRb3z79fWr21ys96EKnpMs9oV2+QN
vV0Hk0zWkEl14GXwk+7wWGQcXjVg+OXnpaxv8ZHIRiYcoqeySU+lsjJ+2aXAZzFu
6XQpwpdXCz1bRlnogpVGoOZAWckqrGF78vNUYsUkIdVSBPJcDe5gs/lSh0iy+jQy
PoCFFKy0QwyvKxZtrUOacnzIb8QU8Rw1JnQrpQEG8dq9Dg6DPP8kFUx9MB+UdF3K
a8OyyKdT16gyqQsvheTQjyLm9a6LPfR89Gc6ZyELP/YdT1QBEm59awFdM/JVAwOl
CzPpivIZwT+RNx6+eyVBMy5VHFzg0699d4QoCt+3C8HrJDnx2A+/4/Vo029d+1rp
MKtH/sz3/SUqJ64oE/josWSd2jlv5zoygnakGfAyxlB8+61KvEIiJjcMqiQBR2zb
ZI7l5GY4IzT4zbhgSH8daWergF85PZ3o57fOFv5NMmYoBmiqCuZUbASy/kaydyqL
hxj5V61Vh5MXEPS16CEndVBZLUTLWbaZXiJ+PG2wkwEwXnqE87ITMqg40vDY8sUa
j9bY9dr8eClYpDDybciyR+ldclFRF+LJT9m5svv8kV5suPgdISXvDAPqBb/EnrlI
JvFqbyFG5nZ0MBbOcvzWA+M37cNa1+4Get4SljsmhYf1kTmlPsqRZeGOwqXbOeAK
IHxueje4YlhJnoM03TxtJTbcsvYBGXtbT0YKuUxofqL9+gIeXC70qwwWN/AwaKS4
9tIG/hxk8HmWLKPJCWEkP5+k0ULB5Ikwf9hKR4QAja79HFCXOqG5sJIkJFeisZIy
zmdfKz7WBp14n/qKFkS8ei9x2xo9dP83oouoobC0bli/lHGpJ9Lhix4QqKhnM2wi
kff5LjbWmC9ehVzoQRFLeaq9XzYvh5mAGsiID+4zgxGxjN7MZxeIUXUUYHXE6NFh
WVKarN3yAvlEJRfvytNiZ4QG2KtpfPi78+Xc2JShaxNG1prh1Q7MOw2j6iNBLgbM
sRiffLosLv0jtmeKGRGwHI4gTP240gAqABS0XUzBHebf1+v0cPKDpy79XtX5VM7d
aVQZfnLtgcFBdB4r/rk0VgYBdGzg3T5YxrUTTNawK2jtt9MMK9lmUVpTFnNR+5bZ
HV5INeG22VOxCtqwNwl6PDuTNN/yAYXofun6P7yhnKy8Wfn0qmB/dn3WQMg29cAs
AbUhxraDpDYTUwCyiHM2bDLqupVLDY6WBXiXmZ8bW5LaajJlAUYwJ9vi5b9BcpLR
yQobKRbDkGYqOoEpY0WqJOXIMTFLzp9zncWVKUY3cVvhXxIURb9iOqPOnD9rKjc8
FFidrIt9vhCbjHWuvRPXdBJXEIzOiXrAnewwASmgCgnlcp2rClwU9+foTgZuSXeZ
yXn80mr7V53QwR3ONbBSarnbiK9x+tE3Lsu+bMdFDpAeQWNMsP16I6guAdKIC6Hv
2OW2b4M3uk0fs2vrz4Rph4OAhrERB5Q/VcByBQX6Gf3miFDrgZJQloELmqH9vFTV
8/eon85X4ITJv/l/5RBY51vp49vN1oLfRZK3j/Tqt2IwCSIvyqa/wx13Un4xyZAM
T+bTDna8aQw6PAATKHMiYAj16vKS7jXyoDs1xuTvz57Kj943h/vjoq9tq68O/RW4
5gDwrIEO1HXdiQs0gG6rdtgNNO4Cmp5qCpgu2/JyrkRyAypBnF+6qb5VeOG2guoI
/aV0ixdOIHmKHFQShYejgGDUOOhVuXHv9pjpZnzIHBCQSh9ERmsoqzm/SbMFMk+W
xvx+mSqEdQcLn/s7hUsV7exg5Hp8PxDmFUvcl8t2o69tHN4DlOcdESRhcBp+TRqr
mCI/kzIMGt7aZHjFzu+vtpLOGjc3TheDHWSzlZTmHrH+NT3VR0f9UX8abqNELB27
K5ysmsfmqCaCr2wrY0qRV7pCI041sSQUmGEYxBdMEKAQSvy5biEzv6kR/r5bxAAE
Vq1jSURpDn+b/w0A1sEBQSZsr5N+Cd9Ae3wXvnRM1x0DpDJs49Tr77ucwkOJz6rr
86B7qrv8IUtHdy4MqBAwdbc6a5rtWmUU6PWow2owHXO4tipU2iQy9JePlcGFBXcl
P4561r7J2vJjRzapdced1FLwpvSTIaLccEwTlO3ye6FbtV67WsagJ7Zpy0d2N1my
mDjIfaNQp92NDL39ATCGZ09lpUeVO74z0Sh8dCczFQaZBOZ+SXKu1Exz84wfuEI7
Cj+Vh3X5Hxef8m0s4AWviVLKg5JOEIRqRqvEfd0vNVlmSzUdRWEh+L/c9/lkdL5b
tPioBFWEut+71fzrXKKqeLGN5fOUDd2QJwR0TDeZ99b9oRGsikNH2GZbs95QIUc7
ZTFWjXiMVsVW38xAuxzm0fHzn+rxY8OLjzEttLTSiEmAuS9zbDlAl+lJwY2Ldpyu
1P5iBwF+6gXZi/Wzzw6hASlkQLd41QMERPoeLS7YcQg8RGNC2xAohS8N9ZCM7rxB
sB/9t+xANWv8X5ETZ8M68c10lULlkCPSPjNko2I7xxwt2048C8KHAJnjz3UGxO4J
9LGsaJvd4Kx41aLI0GQyU91wkvGsq0biqV5N87PnB9CFiB0K93PtGlY7+AOibfJ5
5Pr66KGgq0QAscPEX5U6/NTLYQRvaIfbpfBISlIndmkoywaGeOaCoyXQJLSRjP18
mXjsvsB7zi9Vp4fd3L+dVHza+f1kTd4Fte5XDjQpSQshvfVqVO9tgKWP7KDfn8gr
r7a4xMtjEK+YDsLER6/BvCzmnPzPScvYPMTAIr0QTWfjeLQC7K159OWXHbwkgKIv
Ku0Rte/rTd2+nc6sRr+//kkbTZja2wu3axr1aqY0+otnzbtRFuuHKLo2X0IVtsJ7
IriXnO9U8zRHyeu8luT8TOhtd2mtqBJQCrUH6GohJ+170wTz+O9HWaEPGcZYX0KR
wVgrE9edoxvB2SJa1poCeqw67k2PN2xFdpJkspSXtpT1BRLxiUcyM30n+APMCCyT
ib9AfHG0ztfs/AiLlEe2GH5WxraMo82Xy2mPdRl3g/bcFIRqPlNaMwNmqYTSbjrk
TXw06G4jzYE1vC5w9KLsioFIHKDwmQROFu2klMYeyfrsLWtgTE0Cyh0MaKGctaOu
Wwrcd8+wu+VNMFXq2nS3yh1wEfUyWp/vPU5DhOJRKk9b0FXLTtIkcoyOsvNjlMjc
8C1cdSm4xTViyerCaZMxUhINpaDwvUe3zzusa0y3KFldpAbnDOo5YgpztGm0HQw3
2UWaX6yLAA2xwh0PtVOKFILabrzOJvUwB0OQQiOQ8Pbui/44rT+LKL7mgtb2s3Iw
eYj273gCMNpPerO+SPnj1PUi/M2AByC1NInuf6CMBa644X3DaM9JeYuq5Cye8YUp
BWDtFsTTQ920S6VZJwUVjNB6D/AzOAZfOS8X/D16DWs0giSYQHn8qaWHoHcQz0SK
un7HudOsn0PfLMbrmnap2x7LUBDll7VMgQ2IvNIjz6LQgegcB17oDYywqKSNhypz
A30PM7P2I/uuH0WHa/mtjXgR6Xd8TTt1OcomyO/EEmFbvsF6CLQmDSvx/juJSw2H
OCzXaCgB+pRz0f86TK3+oBDl8WNZeYxoDF7SZbUQ446PKxN8dAQ+VKjDRrbGIBye
WWqL/NvAO5EKXnIAFgnKuPx9WQ9tFbDPgOkFNUyTx1gQnt891WYvuYb5iw7//fEM
Kps/OEYeMYzs7sZZdnBROC7ASJp3I+95Wf0aAIVdFy9AC+wEuydBqqkHOn3Eyu8i
YAXr9mtej10JhfdgbcS9tdQE3XbjHghNIdIGhfvoiXGU4BVzFd9wZ1mCm+FgKBEE
IW+hTMSkLKW8HI7j2jcXeuNtrKpyPyVIe/eJXGqlWGr7lj+TZRZByPLToHj5ArE/
7R39qBXQ4KKcGB8yVdsCIKw95U/dyZhivL53KarAYs7jpNiAi6t2vvrLj0RFTTT0
b9xtLwM3Qui+dnB6V43goaK3qF3QI5ggQvVPRbfLnx1p01eF0huP+gD1G+9Umkks
Ax88FMW4tNHn8EOzv4GLxyjyk892EzbqpEGEcIHUs3Ij286d4jAxMjRBo5p0yCTm
6hqXLv1qOUbsNUG5+OnH+j5gUS3suimhk0e54P/oUfPXNiF8VDD7WsUGWQ92oBo3
w1g4ZVtJSAZngqeZKPM6bGNz/naCvfk2L99YpzaS531uBHZb/uo99JTexjrHJxP3
yIdsUwvFN5fwsDMyzTpzUHicpaoCtTJxlIUXAqWNPTCNAMQmxCNTt0S7nSoJhmp7
LCIn4rFcovnhR6DC5Cj1+eflcoajbkX2ZrsLagZSeABjFtezb55ouPLm86JdvHLl
qL/3Szb8AzPPsX73MBTHb8Zug4ozQmjHFrGuv+fJ8WL5er5Is//SmG/G+0tRByDv
8td6z8wl0vrpkwRKXPDbT2rGoJL5vzEM0z3E2k1oXvjQg0FWpnIj0Evcir0qnQyy
7H8Lh5olwZTOsXeAfoDSuX60pMD503q8HVuPggnPlt8+vlImSbvxJtLTiAcPndA2
TyTE77lFjTGPAVpgtj/eBE+PWvaDuVszuRga/Cht95thL2P5764ltbXFN4htGUqd
iQN/szgc/K1JLkTfnk1A+S26JnG2FWEAON+FVzcZ2AqG2vj9yXuL1kY8DiON6M/x
YML7Dtuy/S366+ufkcI2jl25G7UaDCC4sEeGbM3tbsZssEQtD8ZAy86bEIkcGnTN
Fw8OfGdPOAoXIWXOGgBdwyBJP0kv4VtRIoVhU2/ySLcYg25vxqREMt+MgZqXvSa0
ObJtB+m1zUm2KQW5HTxLELI9sw62Rn3ayQWsLeJHeJIo3iVSW3suq5FZI3yKioXv
9fDQWeRbz/KDVEfPfRY6zr5KgVFgKIU2xx7WNfDd4GFDSG/9PdJUaD0ZrcqaLLVE
opVquS8HKCiqjSCN+ARahSvqYj2xtYDrm8MluQqJoUXFu+QtmYP7s1l8i2JWKBgY
+TeoUxJEFZ8e5hWfGk/pLL1Yzv1/0pbZlpMXPY5SJB+YOWRDmUwsbpfKLVDYpcyi
FS2Gs8yPuFik5waQiTIM5Psg/o1Cn4XY5m0Uzf+nj+ihp3zOR3zi9ZhyBgthcyQT
cB8uXWti6HI8K0nsuwFxB13rH1qxFV8+XllJ5V6JoFDXwMvvikbL71KnXRnVv08e
w+SNcvgwuzli6zOdqOkHKxtN1pLE5UcQDxeHu5zZ0yrOw+GPfh8JNoe9P4R8Dvzg
26sFsAf31kRopzGjiuzknnYUDFJTlR2tr4xSNMCIPskPp5lEz8d4E1Bej/SHJrbA
Uet+C45ao023z9dPjcJY9miYXL4g5k0tgcj1oRujQ5rklEPUBEYFpxuDA4a3MuTm
xNeKBDImRgciNEVXjqF2FnVqY4/ITzA7qkiMQAYpShfFAbP40gFis0d/i3qb4W87
W/RCk4FFBKOHteFRmmQe28p7LSN0avu8zMgPuAWDoCRgnXP6FCoAgDBGcr4gdM6L
8W3m6CpiyrTeJRVYgvw0CcXziYDAFGIKsBVpy6cRrZGtpwWgZKtgn0w4irF+rAxj
wchowAJJfa+PgTK4hrkZLXmhMahj6BtpKiMwD0Zer5xmYekdl8wkONMCLHFQrtTp
J9eSkGszbD0k8EX6uu0rd6kaOYmOCa6BHb4AZpfFo9JcOaJQkgLJK4cGnUVURQwo
1tede6mt2CrMgEXQJseJRmCCFecIROxNlhRNgrSFI7FfleMhO59rUcT79qctwoov
CNC30oK7SnwFKyewExUVJsmhvWD+Mj6+uyR4weVfn7RH1mvwY9cd83/wrAm1KHHE
zaKfuPlGRskldWcSU9qf8qJTmOolrwohG2WjLYPLGQw3c3jPaR4Xi+REfeNj42dd
Fsbjx4YYpWGYmRIGtF02fJjxuLvTgoSV+4CCxmkbLS3hgQenrhvpJPI7x6xXgjaA
R726fifNTrVTL1HFnEBw9Ertmc22louyqvBp5sg+nKpAGIWVYkq2Y9CrCJmEOZJa
uUHmL2MCf9UE45cIecKHu7Gf41HuhgWFc1Mqpwykc07Oc92zOUEm/WbUmRbH/0o7
HHI4ymq1qImanDf3KM928HYytr3oxWSIxIaqOqgDSldFLYZQ8QCEFxh4m4ubQHqF
5eKAFA1xXt80RmAiUMW7Xk6w1odnC7D8Ree09HXvphPYs8XgckykdDnt0aCcFebU
/XuT3GKRdzLM3n0TTBw5jjMr7QLjE3NVAE34adzGVinVdSH9fJHNlQxfh4aHaxlr
uCr0ZnwDokCmv6J3cjt7R/rDEbQgdU6TK4ExdCABLrwurVNp6tHZkkPOzaECxn14
07979qk+j9M1TeU0vLg/ymDtsmhhuQKH0MkywHlQ8FYVK8WC+qMwMTdleeXehHjs
1g/p0s7xPDgoRU1MqOHXtiihcqF/m8CJpBtg2qSE/96js2HFADMopEgQgmCZ2P7A
Ic7iL31DjYq+j3M/GgSl9GhBvmB471dKom23lGhYV6p4ls2qeOuHPObHTiPEOMc0
1VzBw67ZKaFHVcclf0e1CEw1AJtaMHQVT2HiY/7dBEFBUIGMc8WE96ZWvCc21TbF
zdaxv5X0RDLJMFeqGgqH4EoavR1+KRwzgVcNo3QTOtnlvbZ9r9aGV+comW4RIh6k
WYm3tkvMsuCoyudW1/Urg42/wwkCT1mRLG6Gy2/Nc00Sf7wPtWkksyEZuOG9XPUn
yQNJoMjzvd9tRDQ5jUKs5UABpmCh5xsdk2vrEge1N9wsQCsjq9ufEfpjDJG2lqEi
CpV/iz/fcMIkQffG6vXnRNGihEw3qqi20KzWxK4RPpeJfiZloKaKUZnXVqnw1+mE
YzDZVj2kpVQVolbEQzHHzTjczLB5TEltdE0Qg8Z9tlikgQNxm7vtg96vcMIzoy06
EdyV/zht/yTLPzNBzrIUcYzLJhO13neRxpLzyu4trfwZ98gVdEmWKhQgY87hNJ1E
2G+dLczZBhR1r3YC9eGAfUEVMumrn/hM4VH48a3YvXhL7UgD7LdFA5yE55NCqz8+
mhAm8PrST+cJeJCNwSyNtbKH1npWsUKo6JM7NSgEB65VMHaNg0TiE5+qV56VwJc/
67tZ4L8wNfo9UWQ4Qt8/CJP65pMiQDcW2iFsYn/vcWeKgcKjawo5SEiryQpybmal
iOqHgQ9oTi6ufjIRLAKe4zsP4gIq3tIUvD7zBxVye6LCUyMqxSTDw+Fx3GBEWYKd
Wz1VuzE1Ym3szJj08QbGm9S5455ZQ6MHClG0d2zBTsVTpAi24qiwJR1aBm9+6pi7
vY0+XLO3oi5sTQJ0KdtDK3A2hl1m2NJFsOTJ8T8Ypzla0BkQzBrkJ9CebdNHFA05
3FYIrHcRzQikR/LDBQup4sHRMTe4yq1CTuDS2GdDOcWSt+Fe39jv1voEyP+zUdeZ
0jzNvVS5vR965AK9uHTPiBudOM0RbUZB74OZwzyX1bHyLrMm/fsFcVvCYLJpMV3b
ofUH8RPHXAbVBENU+svd2ArIO8jNZxyWxhuP13+dYpHaKiRAepMbwT3F96+aPvm1
YN1gstpadre/+V8JTAYatbo/lrOEJLVDiXpD+F2wNAIcjaqg8ekjckP2kRa3jdRq
JNn1Adkt2lcjTWkEM6hOCAzABsbD2sQ4wy/u2TnUar63qF+JMC6Pb3siGzHK4T+j
ZCsh0wgYYW/dEqVULWcauxytwn+hs+UVQNbSEwKSSXjwSnH8KAqC+c+ol384X03r
rPWNpZ0IrqtNqUEkvfqskTi0wofDo435rHTLkpo0ezf/AcEsCJArKSydQrYCxmAI
3m7862s7Yag/7tx5dyxo5lwf8JT0GNxh4jIJ+605dBZgtmvlD6fBloqyN1AQYb3p
79mmXT17K58ADLsXDAztdi1tGppVmJdP1dN9SLWbQqcFJJqNGK1Qb6qx3l2BfkYW
biv5Hrxy65ZmySQjvDuI7D8bQbPNnBMbDCWUYB2BIz9b/v8gNFyS/Or1qXZgmC7K
KZmM470k7+dk3orEYHfxOOKbgDxNenhuoUhc5qI3vNsNP7TKL+n1Ogd5YGSgiQUF
i/hPiL4cHqkLpt+jiQhnnsFOnNRt2wazkn7jh7krB0cp/60XbZBOFsQ6tahgj+Ia
cROHJvM6es8jVVWCclMkPE/QM8XRVljIK0AYQkhurRt9nFLyRIOm8ZzfPN7u7rIr
e0oWMP3rfP/YkNTVobqqm0q5Io5dNDYGAmgI55D+BCO9Ajf6UeElwCN2QddpWx4v
qB0SrU8WJCxoc8Tq5r4X58SJ/hlIcGHGjYGXwW77f1pVGECiLmkyOxMzMJwXOq3C
ZHqhmUAhj5Mto0nsdbJtqU3Sagvfr1coZkbMc68GTeH1PdprM2aGFUEN/O4psDhH
zQVCELDT99trGE4tH9s6kcc2dHhzwcgr/g64QT8ND9CBThmHAvFMgk3MX3eoKVy8
zxsBzzd5hSOuv3CRYbhZlfYqAVXKtdqG2TIZ0Jo/UBFuUoJH2nuyaHrkkGQlsDQd
NS2zEy+mnfjB8JeJ/FKng7g/9N/rgQdbElWkrGh1eWdThsUaw2eR+f+TIJ1KCMAl
dlDKk+g2s3mH4Dh5ur/5Q9y9o81HaxjUb+0pbPl4gudr3ADpN/6GJlo0qT0l2RCw
UPQ9Lu+mdvlmXxTjT76ODcMdJHSF+6rHLshFTfdRjq2Ie84oFCVXE74tH9nQkCF1
GQMY+n0VFxpWujJlEE821v7ETEF6fHieZAlPEaZMVK+rgxX5U20SVTwzZZJy3gm9
KjVOYXd6q+9LUXjG5WDTioMKjG/QdLI5qtYHqAKT5fpxNxTyYRv5vDjTUj2JBh03
um4nyTyImtnmdopn3Z3AFmvPo/CnZSVuTBb4vTOZDqs4ZoH7oxIqCMeoK3FZ0i/r
ViVC3uo0N+lKjSg6/rtWZn5Gd3mddSZvYwU1j9PG5x7g3xILL0sCv4nLaEzcJpkX
JE58Hw2rMZlfBVFOgnOHfPoggmEkF2N/DYCnQMVYSikBRzz3cQeoRx7l1+1ZtmVI
l6F80r1qS6xpLIhk0IJ6H6Wx83PpmBTWyXQ2+BBIqmKO1BIaSJcuhU74qNFFix2U
6ogqYSBTuhvIdQAEVuB366441VXd6gj4UXaLb5bwH64rSkfIbhI3MYDsEtdD98p5
eRhIqmNrA+dX1BIXbr1M9PHZvM2cl1aNvnfManOpV4bbdGmmrqKtTHoIfnu36FkY
rnZECKEBufoktMhwmmNhuPypu9zy2Ako/49KARR7827TC/J2Tz4QPgUmriYBVWlj
FX1cz4CnOeW7lYOaPMawDhL60e/OlgM/H1WQaLupdOIBCd/LbGbcONy4KjNtiYn5
muXgNBi6qF74EOW1hNy9BO+ItNq8PJsdX2E55K66umEK7crbBYAq6Vez1YmjPlqu
2iudSzz3yUl6SNuYQ4Lo+gvTY2xvsfSlpgK634RZl3+0+2rfajy6aR4fp1IzgSW4
YnXc/nB6BoRbLmyy3JNN0hLmXnhkw0O9zwxllLxnAUDO9xcv2E751KAjVVpI0Zw7
eCv7Y8/OPIw6cBCK5+p3WkYNPVHSEpHoitf33CMkgFIZq65uUu6o+0/btKJAjtHC
ynKdLujXvT464vRVFLMK/xEuI1EeFqtOTiwSdoumspaPpzm7EHof/7Kb9q2Vmv/0
oOhBR14efPxxBYpgBdPKmVGpusD/BTarv8gKGO+4Hvk5yyhoanLobCJhpX4FG6Kp
bFcYbyyStdtQi+HWxkXASL1N9YvY+Rr2XOsJqeAzZdrYHV2FsUt1xpR+E8Zk9bxw
TGa1suNtfavDaMPYzsaZBivRnMr8oZJyZmFS500+SzBxwZqmmaPfTKo9CPCP0FM1
sbsVgkKrRQJ9cjmFKvmI3Sh9kQp3aOEOOL1y02togjMVy9+k550JqTfL2XmNfUh1
DjxWFjlWdwHrXSGs5xiGHno31XIzrnPng0zf9Jk/ArWEBTBSgohj6Xv4FEYzzDHz
pe7QAWAoeAMXvpknIFXYwPScWjraKOBRdNfmBOjJ942hfmv12ntvAJ5riqoHrrQj
kGV1833/tOg+K28nxq2wT5eWLOahVB3AzkMbSeTA8HMNT+pfIXmsJaWVTncJ8vmt
vUms5fRSOlVsvIL/7mO3oojSoj5ksypuF7B2nSo83aoIZrHCFtB+sMKyE4AE8b6e
6/5Wu3TFfZpwskKDsokOhxBAgjY5BTMvWtI7lzWauW0I3MtwQHy+hdQfslpas9s+
Q/dKxx5caM/5fRRxGpx/GGC+aS4XBg/sPVDiW+hNrwmcKqEb5FQ7rw8atsu2r4Qb
mvOOUKjez5aF1t4RH9S/moho9ZEeZ/5ZLEhfZuAWVF+MpYac94+xjWHBQvJL8/94
Aqv1ueDLHaBb/f856DjPCqwqPA4LThL5cenngw9Ht+CjAx59DoVIvlYiN6H/9IQL
mezk6RSZW5OUCdnPfQUslDwtkkcmkBTSn9hfFB+cKH40Ti/g5/04PeDqDTK7rXIL
9NeHxQw519v6/AnOZ+VdAkwydGRsYXfiqB5WxoMmUVlGu0369Ss5oVe2tm4//pdj
jf1ovQJ58yzfLr7Lzg5H139Af1y2PICAkIEnG5RDnF85+36KQsqpKxCNzSBZcg1+
Mu2q9frgeiqnJGcLK2uknEXzl7V/CNS4aOfrvlG1vx8viILL5JbVbjQQvGHeTR8S
/NHPsChNKIDXFLajm9r578wD5ZaopkGeJG/xIFWgMj5JDUyAjrgqqyeap/CMP/Ob
ca4Ov3jn9kIuBTAEMNa+Sy4T8CH+qsWTPOPJAHB6ulb1Lu0tQAGyZW+Ejh0JRbz+
tvu2hSgwUL64AOiwHAXAMS+NT+82MtTKM+YeEjg8ienLRNCJ0TxEkf9fI948PPrb
OT03Id+yrHDmtIHoQUXAb2YtP7K33QPs7vU6qZb4Q+frrzbGaNhOAicoZw1NkQ2Z
iWJw1LrYBSpTKnNPwRi4/oLESoLuD4A7cPHPaPONKRBOxAtQ9gnrWG5u6Efn4DPl
q9O7ddrss4vt6/9VdzXmO45ULaruXMelhxKiJugccZLeF4RWgngkc2Dfp2NiCdUQ
/BK1rawSjer+DzCKYSpMDSDsMeaiAIf0cPoTEMx/LVvyE8w+T6bLmBBb/WTBinR6
JOlsUAfxFvNUS+D/haRhuI3GR2OfoAV4PAPdumj/lfBpOb9wHwcsfYsNnKk8dz16
RkkeajNTG8euJTVSsQkTHTutdSsbYdeCREpxmZCER6feVsCE7TYgzvYw79hqbWx4
Xslo7j8muMQx4j+sEu022x5/FMcyMHAn3K6eQdNoy6lUqCxJFn/Gvj65plcm3Pqm
KsMh525+VWZTGjXWYY5Hsymp5Sq46JqmAOdkajf0imYHJGjuCT64w9CsJEYpUsGt
rgpN+0zpSdK0RCCuCa0/bMCG5qMkIXxPGV/WhKG9ZJpGyp+KINZ1VMyBPTSvtg7q
rKNzSn3YaA2appKJmzd8v3pHB5hckpM3mhcN4KE40Eu8jnmUn9V+DgRvD16F8rUP
+rVfezCo/YIiTF36udrQDeHVXdy8O9t1MaCDAUvzMT7dFmIaiK8oPjTiF8mXgen3
woETEMoS7Thd8PtsV6aALZ/8RuuVceEN69I1xpGc2veovg8yDKtpacqtjR35Ih7X
GcEuqP3ZSTGmXdyP3rmAjjV3wu9LCs0jJncGXYllNu4kcma/zZenDLJCXcVIjmFy
mwKuG881OLGPLuUIQsU0N9kJumbJTiOpTZtUP+Se7xforrUWBdZPXqjDkJoh3uKX
apnwKk+S6uhyRkXzPJnn1m/UIbtPLk1gulHR4y7iZPjrtZQjSV96RmPGe+Po91qm
pjbQE5hmCHiwr+ZatvDb4ANDcDHe7aOd3cYHELuS4jIKVG6adnIgQgIsaQgdbwTV
iKfpFnFUax54d0YyhXJWw/aoWbYu7DYvkD8MkfAD1B64EO2xHFlkj3F3L00z3IkQ
M737w9dwQgYMCXXpqlX5+RZR0h75ZEv+25fxyJzJaGpY6YnYdaQFfktetHNc9jd+
6LdxGxgUSLqOC5UkusEUWoJWOb7HcSb7Q2Rx46fGotv6EFOsxhVkmY+zqJp2CxGS
7BdJbgUocqKKoPxrt6hznR36NLU+DYfY1ny8dNdV3tI4q+r+JNoB6JXQdBcxQZZZ
NlC/y49tFAPYEQog3e1uAzBln7L10Gg59jCt9C/XLFLHSJVi76e+Np4PAcLZcCpL
IcW/OARZkMyB3IxqsRNepYbm9+Ekuql0eCENDh9vgIF2sQefHJ+xIg5h5aYuiWxP
hVZkt+MKTXUz46q6VNPoUR8PNsquZw7UY9QULx8KEDzTFhEVjEluGIu6Fofifn7A
39Ju5TZ9cAaFm3pwniqNMJo39YHW91q0ucWEkNixRXEjQMOKhsp4+MJgyA0ZgZ4r
7db4kGaLq6c8wUqN6FhzBBCcNH9/LY9LtMvA4ZapkFajuWKLQyn+61o+qTcMHMgY
w6uqMX08bRH8KvFelThPI6heInDfOtf19IfsfkoGc/ayhK7UNfu+r3ScHAi+OfeG
xvbJfm3oFM3GHEZ8JGlU8aeZFSSgXvm0RdO6Kf9S74Sj0XSIUm8Ez3hh+TuSO9+Z
RvMNyZHMwfjPk2KDdZrWXguO/P9YgkPu2LcSJofKtGKBfNfa6gyZQmOMVG4Vv713
GyAir7bVPtD4sNJXHm4vbDXCNwbPwaMnvF/TIbWppS7VgB+CnLR0LyvWIn0hQDzK
bqXAW4zCT2TmORhBhg7nG38KD88/tn2VRR7WbJvKIGWJRL9xbjVxa+EIGSbyeH6G
vTLCqxDRaUtFS8OeyIsw8tYY8WFfq2bBhIUiDV50h2d2jooJuUg37VjV8ynMPYOC
3ADeUnUZx2fxshKpu3uZmPmzvEua9F1N/HsffAh/xadPo3QhYT/EVZdsuWsFU9dc
irao575/kZLgQlBwKZU8YTUMvQF+ijdKq3UlLxRUMCmZ6/KxIbnJ2uVc0O8bR0+d
ZXrUAhHxxx6ojrzUxd0tF3BZM0SOK36mffu/PD1EvAMhcP7YRZ0MNLImYd+m1Hho
ve1ZYx8LCTminZQk3XjBjyhdA8vuBWzNd02tETS5ZG8RqZY0Vetvbp7CqeY0/2eB
yKuYQly5vvoJKTJEVTZzPZSMMvat0gwmfaARlUWhNYVmCk1qiSdIMcqrptF3h5UV
TykWmqcmF9kxcMYZguYFBpFsyh1/5w3itNn+icAICXuwY22zHkfny1tLRDz44A7A
rQAGPsu5uDTWUYLB7Kj0zKE3SGUfeOGwZ71heh+eqLF0h4eE4kSZG/4Qh2Qipnng
Ws2sHlQREnRnryG7YmGLCqoapie+RfG9Z0DxivmTykgsOIu4dojHTCAINPcsiJbC
u7E3qGVTNzPKLfg2NvHR3Nc2IaZ3bYL2DfYkIWAthDaDQNpXMdI1WORblXOURfbb
nSktUJ+zLxC4cQW9adainluwF1SiPnKC6sMkGKiARY5VK8eE1YOPxTRQPqrU/wOG
WHh5tmfqSbjSH/Sgip4/KuOuGirdEEURUFo/5RtWmd/Sna37RO/68Ip+Lpoihvvd
7kIRoiheQXedpHDy0Q+MvzRiMIIb/nfzLwjsjeUZYhw7ISaBImxT6VWkmfcws2OZ
95MnPeHiYvmNBKmwi1Ro+tLbsa8JXmqtoZ1OyEoIixwgEYEYB8uPrx0YSYdHIro3
00h9NiSmy8hucPOnWC2JslMzSC9nb3LO7wssln/spsUFC5fB1NnXGc+j8IZOK8AJ
Uz7E5N6tVvHhWa+tMMgasnczuDhUdcTTE0P6FdVOuXikDhZ5Xcf2Kj0CJCSSCYVS
zwhPiWK27wS+SXM0UT3NRBLnwL0WW6CxnFiVgomLG5spPWBHF5RjYxPEsGwZH6jH
gvCy57LLC7b4xYybkb28LsvxtpvVjYzxBfupTVldBLU45/ZKSGVyjVieX9Gjgp6B
IlllUOcqg3YeQ03XtmU2JxliRtntQMg8iK2cMAVXe2rtJu3h1p75wl2t7z7GfzK5
qo5Wv2O1YVBi8lZ85eFhe0ohQSMybaKIvPmV+bDcrdil9NbA8QNUjPTc7OemTaRQ
pMDTeML1qs0vfkKuRHQtMLy10fbN/Yvx174TwqQI815msq3hH58hEN9QoSBGl8Z/
j+MTWRZ3RQwWTZdbtZD57JjO5m8SNYSdchgDxZTzg6C7fh15wJqSIECZvk7BNsUe
gJUDK8hOOy5iIyem9bza8HkJrqOPMu4x5su5jFHsgSEl4slj74M8cdgkxjIc+xY/
3iut7Xacs7frWPM4YqTF0TeIlyFiQORDC4TLnTUvMW6dSfZFYBke0yr4zGLB2Iar
+ebzbh3I6Fls1sfjhcbvt3LHbUH8CbDHMWoTmqcXqbHzk21Yz7/Bq1LihUa6OWJO
vEcYyh8EKnOkNV4I8s+7xo41yGQAIwogjshaYmLsFE2lMUH5ZVlhuRusBB9V369K
jeTmPBAXCtp/uFV0qs5HMTDq4ITqzb4oiDTFJxDb/qmXaLmC6eLLgYD1jtPeW3/x
sz51hT8+pu07Q/zIdOniQ5IZxiwRVYBvTATXIQ1lzYxQRFsq71QVF1o5JydfNhO0
O1md/J7WFUsDLZ1t6zVZ4o//VplCGgoF17+EwskmkLB7E6Rq7mKd17lB+wBAIS6W
w6ng7gxOai27U6XiW/omvwyfNUQUV5oGxrdOuAydHMkkdEZ9Fp/TwP9HqtsR2PtI
emIfDqKr0CLgfH+VpdyXaZJ9w8oy2mFx43tyB/a/a51qeiPuvPuJ0jJY4rehNISU
Tecs8Z+jPVp4W03KUt7mDP3jiWruBcB6uhfA2zXrn6GUL7PB3Qex4AjDdJiWhf30
OGYng6T+/5WsnbxiaiikpXA3uA+YAH1+jj4On1KqD1SC0Kjy8qc5niBMvu9ZCZbO
bXj71YGgKz5OpsqHvph9hVloubeWzItA8vzt2y4MQHXWuoDtJLfvU7nNql8hSlnI
8xwdBUzjmkxQNJhDRKfittWjg4IXiGvB3s+KO0uo9pr+Sz1/AcdKHB25pB7oIkLp
TmvYZgydSrTCag6HqUR9cPSfkHW/IIN95oMxrzH25az/x1PsKQlOKv2DnOfBIVoq
DZ6wvSsAE0ZbdisC8nGQ+9ehzSP1anCJ48rb6dEIjnBNMg3N2wvQhpDYrxOacxS/
2ehnDuwLpcGqbiwf+fC6kp9G4ZM07DQ1fg7jyGrMLmTowxQLb95EZ+nH+mUszUX6
sMGYzZfavGS9pJ+//8e8zv73oVk9oi0/1cAuG8DYO8haD6Ze4NPfoN4MVdrmSUN7
Q8qBDlabtTTKkmW/ArnfxLYWbuVPcLxqws7QoajWUUafxwIm1y8X1jBudoMbPkxT
SrH+LwLRqvMNSRx3uMHp4rGaOESPKVbNnOZ55krqI30rDNx8DiamKOvATwDDFP11
zZ7oBfK5IecygB7a9WvTagcowhT0tsm8Qsvown6mCGz6RQ4QNlE+/MoPR0IDq34h
YFhI6ogj9bDr+eM4YEfpGsokjWf8Ne0wEd8yAhNeFMWz8S8GDOEI5VNUR/cUHOJ8
pmGDeFiOzS7KzrhmU9HGWAgnUvifNcAKZ6AGLHo6Yo5+ljZrsQ/oBotwW6gXPKWE
2HBzcSKpozoFlYhf3mv4A5AlTNtUns2EFEcjD01wnq3QVuSW/36XhDOvQhGqHlDb
nuvLWR8xAsrvfA2TalXo+cZzXu/4gz+uhhXNgPCgzRRIMH56e03ZuuaFIaxktvm1
xTEOO14YLLhhGncbFKVvJXW7RSUE3jeVEIf63yq+/1nargeDlZJF28zw5oAol9zj
ivJ1Lm0SvDwZWRUdxwHcDGhzpeL8Z/TWstI+yYMv4n/TQqikjknjxxaY3jdW9Qq3
Dml6dLAiPEH162sIQkUj0CPdc+yzjDv06429G0KSAL9j2E4AY59yNYsrtAHMDftm
F7JdBP/U/uM5cCYF0XD5ZhPprJrXF6vJRZaOe4BL3KjiBYz7xqfBDb4eTlCSMuQJ
E5DE+CHV/ATIWzngkI9l3DQyHGUYsYk5QdRETERP+XM3w89FhSAiY1fE5peAsWnP
Q4yP/NvZXvNLbZIHzUyMOUSKwZRWQNCLWKPzv8K4LZJnIAcokqOaydjXh4a+gi18
nCPLqq+X1E+LedEvow8deaICsbHRkYRuEfo+Ls7Wgyz7RBUc+A0b5J15fvkG/bnl
jW/ipAneGKf9gB3qbz9NAFSwZll9ZfYpwmYfwItqwArJopvCxniO/969tkNTGqKk
6klbWFoM/2GUDZoJbMhcS+oS+Y9DWaIVyq0a9uO+lMUTdbT7GQ33ekxjMPoFNead
yemf5llEc8t3RWkb3l6MuPbxzddBpLyhi5zp1SLFGVIDkEFSCONyoRxn/xMyrYdz
+TjFc2Xe0v8LsrZ66nGl53j8X2mlqUAbuuuKSy4Odkjn8E56xcVjjD2QieAUVDdM
t34vVzG7x8qVIoxmTzyjiSF4bZouAKnKsFvbvUu++rAWUXwScnP6icxy5RF8mDbl
ZhLqwCEMLR7mN6XnZ4g4FjIb9lAP+PimWkMARsW1TcUxRtb8pxJsy6KoCsHWv+mB
iDaO863A93BbDMYQHhsY6Md/gOZf5Fwl69MujQW4rfi9wYAbMgrajYLHw1IC91WI
G1bkm/kL+mwddNNYWmLv0GGNjJ76AMWDrGmyVlMeDYQkys5yJgXFNpPP7xv9D1LJ
lTH7XW+9DyXHvZMuyhIWBtxA/wM/3VIDJ/Ix6wzWGrOa28AhND00oNWph8VxDXd/
e4EfONAocv6ELU80IP+Ak27YTEbCZL8qsw97Wh6XzyieSfdLng4wJwMP7AZUtmGS
Y29j/H9Ne6n7GAHYsQf8m7y+BsNXW61WeqvqY3jjQSsKrdFqJD9JYzjdIqUjoWlE
qiQtn6Jem1rP7vb/hlb2T5dPLZoiQCTBy+8uYZldUzEQKCoi/oSLqxi+5fSEEwT3
2aJfp6189NWUOhYCYgbyraaV6PTT5XIQjL8JaVq5VU9BXXHYfhDLLpPSZ6VvkwSY
a7CJakIVzRPBoBOj5AoFn9aFRkw+TyQpoCQAS/vd4VRR5h3i6FQAhC6n1foqmUMa
UUFlVuCCSji8bJodFcHixbUL2SBKDF/9evdN0dxEs8898ZwWHrocaxUi13JLP9xh
7QnC/QlDQYi6Y81uwiMyQZtaQDmOa/CGGEzTBSu9zNbRys9kzJyVYwmYZIaJ3YQh
T5uaVThtHc6hj4TuXBb0jggvuSlGVq6lrrrODNsldm4P3+ku3OoEvb2ErBv5sM1P
trCUuoWJP5PiIZSj59hremz9ETFfBGbzO347gwysj1XKUrqG/r0NyKdLHLAWc6FT
6HOnbg/ueRbNBr0jcCy275FhfAFXYvm+O7To6ufT3cEHdEBOPinPj9pPHZEbltd/
u5NXYHi/lgNmceGKi9AX9N+YiUOTD+6TJis30fPH1rUR2Zmx4v6kj04tV+aapZE7
J76l2uk6d56sKcufNRyQ3cmkHH1Cv5CYyaw/7zOQJodys+05IkuGHFCRij5Fib92
hpclHqQvGDxNcNKAZe4CY9f1teKIfmsq9UF5w6RTZUoUtGUI3PowY3Kt+NO0/Fmm
CKc51jtAoNy4ocMopGboXydPFNX9aImt2v51xEAgc9In62GT9AqoWC18F5D5ldHt
HAFRwotKWWAOEo8I0U8POCL+Och9+29n8JktWoIsnfmvGdR18aE++NAR23XfH+aA
6tB+jxPd/nQloaSwjqSjPQD0Hif/qGmlLuADAA7RvkWAIqqR5n4duidq4i3ZypKt
qFWkPfMJ+jPVsBGrt6t9sr3aZJTUAXjrMfWr58Dv0pJvhaJGWtN7w2GmWg1IsSSi
hzqO7GEPLrZQ6H1c6zTCBmbJcmWZtOu8gAv83NvC1GlD78ota7Cwncti8T38b9Fc
3jAS+y1e0n1bNjzUcOOEIjci47cRddoQaGCEuUuy1DqrHBBHxR23xvbJKKd5aLY/
BlLSqwhUNPziL/IoVxVdR5Wsy7tu2gZWsD0s1fTU2yig5RFlTdCq6/IPiO89iWhd
OgM8VJ92CtAk5Vz/NtWuLYjFRc1m0RcV+JAmKsv+TGKg8RKPiqPCxJ0krj0TcYym
2gOl8KT6oSme+A/Vqt+wa2soXZT5hVm3/PAHP73JYE+rSQ+Pgw+ZTOgH6kXxRVAu
VLScOeiEKBPF2d1o4A30QXaSSvdbQvC/5nKvLBqaKfSCixWIMU+Vs21jeqe/JGl7
rjLkYt94fZW/VHkPTBtoZx6qW46I2vXoJuWUl0iVtbXM4tPz/wd7cc5MywlAI00T
CavqQvWkNNiceJ5BpecMNOZHatKSakdWcLMelyin7qN8SRNow7HfjtpLKwe/T0wx
+QV4Bvd+zO2j/wGrcoACfSDHmP6kJFtPmpMyWkgM26aIC2lOyeglG1XKWZlf5Y0x
/FwKr30PztGd/OkxPAoRtP2lKwieVtXcEOTYsljCy7qMaTg/3artIlkG/PQ5X4D7
yiHYodZM0nS7YF7SIBuXj++ak9KY/FQyzjtFKrSvukITlQ/aIKLznbO6dtOlmthc
l1tS2aF0LXeA25bRAQ/LXyz88t4yu3Oe9zyJ9v/S97t4Olc9ntf2V+/fUDcxObYN
lz/ZkiX5amUa893HA8oYLUt3prWlHJwZffq7st2/UujELzzuNDNdAcHnzMlpfVxi
4F0mG4q9ZqBy8Z5JqqzKFH6gRl2Rvlrhf1ULuvpKklpRaOww5ZE56zB3oecrlqgv
7WnYRVRzu3Wj33gzAy9tDB8AJu8wJ22rtaaMUniqa1837hZ5t0Gs0XSavq4SkpHt
Kz5rLS9bTadUNvf3K91p7+Ctq2zYryKZwlTPRsgimmvyEIYyiCe70b9rowx4sJ2n
KAEf1UU3w3Iyc0nJFfvvaWFB9SkLVitlis/0EzFFVEJ828dHlLAWO972M1yIScSL
9+Nvy/ERcuak6QlMQhfQQkFT0y9sfNvLtNMiqbOz/9QcdD1Q321A2jpWO7C5UYVn
4FaANGkixSpjYGKZRJsrFxmhuxnDyVKZ0E4wZnBXxOA9ZSY21NwwMPOlwEOWQsps
qrhw2TSs9/oTRuTyD3P1xS2mYJdPRBmSA9RSMS/xf440bVFObKL0yVz8bweSJBC5
cp/yGrj6844FtE6fH5RWqctb3K5gqN6OBe7nbqjixkbXuAXEH95rcghQefdUlYEX
IUBe95k0ubE7mGCS6T9WaD1HLl7ZpKt7tO37R5wbJG9IjZojGzMSmlGt35oRLIQ5
y6SKXBxOEDP1PSw1NDD24Uj2By9jjkhDtHGXxdvpJzwvZU6JQg7eGb+rwCm4/5Ub
a5nN+FJ5a8FJOIesEmg7VZX/P8vF3PYuwZrY7jnMjbnLOHcfYQvZ0EsUjnFej2aO
+AnSiIanEX6dh1pmfjRUnTndPDbwOPQH0by6w9NuFilnNu7yGaG5mEy8GUWLu0Rj
2rGE/F4zHYLFmWymLrMjvAMdaNF2ea5dsym5B+8RhKo5YKHvgi3myUUfQbQmmeV3
jLdh58yF13sUqHwX3My/P9VLL4hpPatw1u2HkcrHKj1ABjCKRpXjm1xY0434OfZo
LuSJWS1QIrapqvHJCxa/Le8WcGafhXe+ymfjXKBVatqNVnRbUpP9Sm5xfVpv2CbD
AkKJHQ8l9CuKg5N5Afc1vJSh9XhEpJUzVYRZaGdJand3mNu6iPY/EsFDHhUSUP8N
l+Ji5WMszwRg8vVAUj+yr1+S52WRqR3J+lTTPUNTOj01HIz+H88LwU6vTExDdKHk
vyjSJIIKG4HWKtg7II3sp9X/gDTWf2S+RsvxOgukj2DqVn0JndVCoVvU1rRE3FqQ
S4HfEalvedYFMnDysVZKwtp3PlXHNLUQoupBqqDndzhf/3rEsf3fB5PxLc45jBmj
RVwGH8Y+z6m+wCK3bztGxnfomkMgXL5ior8tC+M1jQnnlQwu+eTZUoRZO4ep6/YI
bY1Ls9SRgR5ZRfSjLtUD3LJhBxHq1pmP9CLw4RIrYAvSyv0t5gFSGjeTkEZE2pKX
HERwIhM+0GZU5VkO+6QQ5IpIWWcV41c11HrEdBWncR9793EC2LBfpILv3h6F/t3s
qEWCUjKOf7yMzU7GErkPVgoQbTTfBsmCcDppL3FDIZmO0nFAaicugy9e8PN3qha8
acMHzPQWLqL+bcd277Lq3e7BSR5cxB9o6yX4UX3Dq+DDCWOXwm75Dr/gJAyOx+0Z
6JybNMm80vfE84zlg0xTAypiajfVKTK6bMmBjEIBucv8ghS9ECDHKTSUsBFcejD9
7KEwtTb0nd0I+5HpONvguqwA0lFrX8vV0uEMD/CVD1zfbhhwgafUNDZCXBcQpZYz
RrUav1d2aybrF6ltdXBxZRBYIZcbG49BOe6vMSkgw28NMdLt+ZszVb4xCws+MEXe
fWUV4kZo4Yovkplh7+jrjuqXc+ktNDhbxN4qx/A0JAaO8vCVKeTlBccF0ioftnOA
7xnGElnVzCnC7ZxcnuWZpz1BWS34Q4X8w9YfAbMLpjDoTna5H4ibPAJABm4W9RWW
1X62GrmczSkDBTOaWSiG3x75bZs5oT9/z65OlHw93C0pCxyz8XRup2NOBXZ0/H6l
JQ6CqEj2gZI8l6QtyujxA5bnyh6BgxWcyex0A6b5YNxmaX5QTF/fOOa9Putrl/+M
cORYe+YPmZ/28RY3LI40aWMzUpVtSSBUNk+WYcD9AzEFVWnniJMCUF5s+pNLnhON
ZS/0l+wOsJtzP7+t1gxo+eGMWA3dI/dUMifVtBXhp/lySOWKGT7M5W6YMzlW/QtE
ygX0BAVoc6DlqGHJ4es+6ALlHc+AzmL/5RDCXkcv+1MC8Z4EXr6L01GZ6OHDlc39
CJw5e4bbUELJg+A8dfxM0SfssItcNy1IPDEKQsvcn69mMLJUjRFkhv5StfoAHh3R
BG1u6iOCnD8fT3Zy0K7so09Ye22zy74vGFRdjZ3gaxmkDtKvRG2sv+AAx1Dxyz06
d0/NeMR6ad74NQ5g/VGodAGNBSuUdrB4Jyb/z6bzqoLPPUfiEaGBrF+U31eA+C9O
Dol17oSr/+cFfqubHOTYd3miSUrskl8VqkDzHxvZJDf+rUpqtMUaagp/7oGU6NtM
tAYR/wb5SPUQFPoLDTcd0eLxNBK5uJBsqi7VT8k4qsT62O5VWS+h73QXhOZNAkQQ
xVIfu1tJITf7zCq5tZXMs1MAgBw56CDfNvRUOCxoJ92XCgMJLwmG/YzBdRlZrdZM
pU5zLZZ9+Qm590gKxGV82x/eZJFTefspF2vzxFde9yWa15VZrnoMIRd0Lh2Qa0Wo
uOu5fDeiuhXJvHH/lZoldxMSr9J832DKvgURLs8MOf4Mvf9AUceQW/PEc5uvNsTv
tTBFTH04ri6yd9wcUrNbPsj34BF6B83V4jM0w/pjNNRm5op4xc/fP6OkUbpvfRWP
rFXp4HF2quug9xm6hqJRcBt8tGR2El+gliwLIukkr+khnPpaPKyXNXqjxs5CVOux
7lFv38oAg8J6M5dQhriCOTJ+oW2f4wcUm9SLzXL2YBa4Ro6zgmMg5lY8XxnruI2/
jO/6CekhOBIaB+YkLifA1rcTNMOULbkXREG3AQuoRxBzchwp+0A69/mWXdgC891n
ihmMkxgNTZMiHNHFXomDyFUJ863ReLprGdSI/W6yxPRBsNeyCaKvy3nj0H/jolg1
xShQZpKfP4zKIlSMSB5snMc+EmiE653aTYsOD0KCZBHVJcu2I78qcYd+/TP9VXhu
mUIvONoOFTdO/KTvbVSzh0b5orc0YWoanDwUbPghjSpYh4TFyoC8l346zfbB9v2M
0AF10U+mrfHx8MFj3XbT94IIQf30/zMC3FsLOP168aRWLe671bOTPmVlwVR0ueAh
WBgzgTjDsiI4BSTLKOEmn7FNESNdER5eXr88lhzgANi7LvOqvAv+SGBmkMgTinI6
CLJQTkjgU9YM+75+OFh69a+b23qAJmpe41rztNUa5rnbuiIXT0APNxqMR0b31kaA
84J4Cx8SiTSuM5hGRGZK6eRGHn6Dj/PnfwjQJiVTKzsE4wYl+CEKMz9L7FqLQltH
gIgwQKkKF9WyrfpKZXNtX8fY4ZF8AldZ8nXtsvcq8iNiEHA6A8XwgTGFA1o9VAVL
gpmdy9N+BVofT9SgZ2Swd78b6YoWotAD1OxDmSkEtT5FSPTjkDZ5U35UstCNGmT9
FHp77qTAhdx2oPBxA1cGSUFwmXcBnl2M5SPIwbhNvdq9ENUYke5jLEo0sdTSNVFu
jYa+b3HPwO9pGFc83c91nnoXFl2MsBENZB+GZxHMKQrdCGuX09MMT5dAEDlppuKp
UOwd0wFkjjpmfHjyaD+dH5BjdPC07dfxUQ3xcNe38Jx5Xz2KboSdjOadDy6F/QdH
8Io890kNtinPeZrpP0vVMiykGql8QmvWzbKNC1q0G431z7fWt+abT6m9xUEUYqjk
32aWy/0Qc6mKxor4HF+Yckn9MeJJbcoco9SHtsh5eXzR8577WybsxmJO1bFQkCXw
2UdzFwGdnDXDgkMwtfO+GMqNSYAFGFLQ03xV8ZpIS1YY0If6RZqgFQJ1xcGvMLEJ
b8xQKs3T7OACXFN2njDKF+32h/k97Ma0KNqLD9OcwAU5SJgiszaTbn2/kOqi6umT
Cos6OoOY7MXjiPDgmOay8bIxY9u64AgFBeZ2T/Cssp2cj3RKegM5+edcvSafB6dU
q4dMRvZtxZXKrCK97bvgpDZioLMKb3CfN9kKRLBdHz4oMBgE1kUuJt1q8/MG1rYs
Atb0KHJwBoGmxtDbbImeqP5DgxsNGmNRcXl4Y4AKdf/2qUi9FknFNOzjUw89LYbw
e459Kmo3Qcp5XXhpW1kBnIjv8S3jYZ0EHRFRyIJIwvTftpC/vCFcii2dRXrUztuH
yCvJKjjiJ3l4DNHcZUglrrA3eVgf/OZWMkHTFLV1NJ8WV9MbX7xTgIDDvjaeusJp
hzoMuifNumYng6+lOomHb5IQcUa60WJmf9fy4zBp7VS/LVCdasmKWFPxPpO6luVB
1F89w7HUydRMo3gayBmkeaFORFPIOvRKFE9qmjg45Xz39Mooo795OlK5pjbL8KXh
GBKjuiNR66ZIbEZ+nGNLYHDvRZXdrNmRi73TSL3RUlrKyHBF5SxKUVdhASdB9HjN
1uqCoMEVBkkFNJBN9UhLTYAk+jLDk/m0OJaGUTbvMzBQ9S8XIPj05WSVJtjbJZWA
70yhQqezGRmN+stKWpbuiOFm/C34/9EuilWqZSilvcZtXrJlIi5l4dC12cAODGBg
S2m91mjVh+tbDKV0NZqBM8TFyb/pu9pTRkXR8U5Lznv9wZjS7H4+qDeRZSqd8khP
b2E3LJtXNWA9lP7um//foNsUH2EP2DnP/uNQrw1vigd9YDnwpA2mLXmVjxBHGWzA
Z55V57rnzD+3L4CQGYn/lJvdvpzxVFbW4CXzmGRapSX+eaM8ior83eD8Zi5ITTYB
bgRkU2pYLr/j1fo6msNxdXmpz9f1rwU9s4zduo4N8TRvdrxdMu5Moy2iPe2nNWd4
PdEydBywa5ZhwjiQ4pXHgxJrqHUU25E1yWJofiSMlHfWgoyUtWn9J5MqoMoyLbJS
VPHBXQEMip/+LIMcrkGgq0pNC/N03xciVfOhUFiJzUzvK1K81uPxuh1m3ediccKd
0W/+cKh8lkjGflc5Aza+IzKLvCYmxxcO+zNNFCEVQjZKC0tu4/84xDtd/guEI6V5
/YTSTB6nQ6cpXooqnPaHombxFkZPkGOQ2WnZa1rGjUSVIsLpTn/94pRNYUQVWU7y
vowRHkrtK6MGqMe5hou/b4ueSo4dQR7kk1OtmvuMCDwfZjXcnUskPlkmfSnGbVNg
sSnV27DgQp3TQtB18oauiKwPt6l7F7xKm4uB4WEGFs2IVPNx2LqomfDvfIuR3ts3
8lyZz089MZht7SvMaNmx0SFNrp3DtBMHYvokxRzrjBH8Ja1GjWf9VUVxDQ9JLELD
aHY8ciF1+DMmp1LmezIS4Fg12Hk1nDbf6szI/g96bBNjWYNVLO7dujWNWdR5ntEp
QvGkm0FRdMvYWgIgAx/S+RiDxFihKzqg8VWTXG8zIlFuaSjs1CkzH4MyTA+pRtue
wpdYK0s1X0OAHWiTCwNKh25PwLvEjI+Pq2v0d1MW1TYNSSH2Kuj0QMvAAUkAhCj4
d7Ea6Zva1LsJAGzOElCPxJEVocP/zOu/wHdlkYCeapf3ge/vtdltb0O8ih8PJxuB
h+erkMfmoK4gXVXulr/utrDBxb8ym1YndtdjOjwu4Ieh7Pg3LDjKJmQvlqwE2I66
I6gBLjEpugOEVgNb5602+hePNScnAD+cdphUUKZbKm4XEUYPlzUAFI0igi7Rfiw3
AOBkJpR9+p0ZkJKeFE+pwHH78PhZEqH+fc7phwJIQeZzPX1uUGqZjph0Eo7nby2J
DMG7R6NfXPyGk94UrWLWazegmBCgCUnTltmZ92nPSS5euUh6UlRDkgiNnJ2ri8NT
iv0H2KUvmbC/PzjmMC5y2ZDOJr/Wex0PaeoHKvaHx4QEr7HEQPTvqA14Kxwp9r9N
Qda/ExYmbNJK2zYiw8SJBt01lHRSAUitRdOxZJNftLJ/M4up6SLXSin4961cMCUu
eDBUwkZjoKG8F8HgzXmA0uquSGuSEQadrFGVVi04bhh7nkXIX0BR4UXFUhwRef07
v5ZJta4yupUXWHg4cUQhC3i89cwB5EznJmHGKsCdSvo53NYDxayZPghHvzrRoIt7
CC+zpgJCThSJBynM5Jif5KoHI5r53846pUDxLM57zs8ak7sQUrV1UcWvhAeMtO71
BZlKWmwL9Lr2HIpHvxeV3RgBwlyShgtGHi5O2Q+fMF1zazR0C69r9/CKMGZNI50C
3nmn62I5BWfadtn/pzK7cdQH+Ybpc3IOH0D1oC3UQbBFTT8AoqgazU94giwOL/Q4
JrSv7opiB4jNTH8QCxBsyvbk1nkLT9ZgdiGbI3f+ARbCV9JYy+LHrHbevzNtl/l+
usdX2kyXzukR0x7XOesi5Ai9M16tenqE34tCSJfgty+SZiaPa0y+BNvHpGTqveti
jqE8IlDaWYuXYJxKIyKFlSWziMUhk/xRi/xB5dQqLJCKSncMxpl3GwSqPVEPuthQ
IQVAxDnVysqDQDvR6BaxuYEju0gatV0oT3ZGZkSlVi2OOT6FvkstcfEVWKzwvlFI
nBO7StSJMLoh6/2dTjIiGeXt72QflTiS/RenefOKSReyLKjj+QUXpolwRdfKnP8y
5SSoy49ZuVY2BwSHkSJuDsix7sm4T6+wSX1+SgO0LJoQFCjeBXeDrRIKHmXBhItu
NFhcPFMPi7/URKftvFKqNyy/SEu4PpAjBU5oPeGc5HXnyEyxffEM7GjlJBSQNXzP
emDafya+YAaHyck+9xxnKccQWqph/inAkqSvLfC7XaTRpYIIh/Su6pegGaI4xx+h
m/MOTx81JLQuNGiROeESTO1IKvzL0zr8B7e9hzka+drKSeC8eQYH159nhm28/IJS
aq2cI1aXTrvtLYp3EgRMv1KXv83pYpXZp1Y2rPQnbad+JQQskp5CRVIIWlyq/T+T
N0zi6C2sV+rmSq7OI5qDsB5a7+X3ejRmkaHHX2OXJa6gAelKILJj3WrhAwKmaHPN
7GcZkb2rDMGxit3P3mWebveE3/E7HvS7M3q0PVYChyBQQLNk7Nihg3bDoyLDM8D8
oo/RXcnvOd4Qghta8AvLno4+Vpfi5T7Flnlf+69GwVSSIwdmORb9nV9pEQDcRl+6
DmhQjlGd3NuhmOuLgRoM4VHhlPd0/AXU4bLXoEielhOxFmwTGtqsXs95XoQHQJA/
LSnfvFMP6A8gcobXaDMorYhbeqNF1n5NXUL157Z7fGLbwfEWeiQM1bkcQJNA9FdB
DMUvssjNM3BPCdzhyCFokZIEIACHvQyXFCMEm8O3WrutAv36v9B8A6EToUzkQzJ9
WefvayRlS1TgTimYs4x8BCGpqS1iL53K8wD0to0IrAGjf+ozb/vxQ1BfMgHsr8aF
RCFzJPlmJTLOu75s5r8lwKouW2B5m4uWFEQB8RLg2j3PYEN1Vcq9VjWFaz2kvPtP
H1jVWnAQ6VuBJFbPMyaxgmRTb4SA0bWGkwWm/8PEdgBddB77WotCT0zwyGXxOJFW
e8kvKE8lVc7qf1zJgoaKTs2iTqZGgErt9d2kbS9yatwsl2OnRowNGi/GFYS0/J+T
7jN9x2QRNo8M3IqDjAhKNhOJWLXP2ue3jnZAjyegVf41Iy8qMtfgDXUq0QG0FyI6
umCDIW9Ox/esl8g/OF0azFtd2SSmcmahYsmKH4e9jEGws89+B5RR2ugD8cyamdyR
wZm5GVhsiffl2x3pONuQ7lIUtDSEC+RtMiDyJaikYrMBh6/7up1ztz84yJxK2q79
g002uche6YzFLmBY4bSOTkguYDs0Fm5UCOjeO/XspzrlReuapdKLu2CGaELenE2H
TpAbjqqCLQHC8FL3c6+7vdHAtmSnindyTKCW0z6NBUH2ZTbJbOlXyG1VqiHzZ6hW
CEbjbp/ycHFgaaKWdNBPuVQrVUvqLt9TAQKu4rQTEFopWK2durWlbAbOdlMCJYfH
YxeaqVICbe1BXl4unjIkBftNhZ7WZOOBbfs2nG7agXXB+A9J5FKUHV/5+UKcJrng
JzPXW9ZWtCK7k0/jJWAv0jZADDB77i3ddUYUjYy7OByYCx99eyLaHNeFWTv7Vvdh
olY/nKb14b14rud9g9Pbf40jL2Fc/HYJVeoXdOYIEiTzZUg557CfdUG6XYL2yAPW
0s6fiK7dh+qc0LNypb94QvVq+w99blRpTzWwZs+IuLfzOzUIal3ws+f9bfTO2Qjo
FhDcjw1jT5Omp40rsakveny6N+f0R1xu5Q2wpw/2jZ3XidNCaTUFQBkC9Z9o+F+v
UdQSq/ret294T62439W0Pworoiy7cvRjrYv8s/xLHEiLanf/LTdnT6xJOpBMhAg+
PwVy5k/AE5/tc33SCY1r5XFiPwTS7qgJVfGSLfwFqRO9FZGKvYEcI6bVC2egdArK
yqY2SWMytIXvlmlWkeTaiBi7A0DuU92+kbUXoqBr0tPehzZe1ukVpOaPO2VNbge7
zP0CwAqvBo92b4RaTaw+5uih/G309LIMEq4b6TVGl1kh2VmmPGo14YEVXkI+DGlG
VwfrsHDp9gc5UdRiW8fdvhHgG3D03OB8rb/SiLFk4KU2FvtjBCFlT3lFl1BXztk7
iVcSmqAR2T095ELUpCga9am9tEiJJ+DgDL1BnlcTJ4cFY7vnxxb2zhvrQftpMIl2
UHM+KcE7TP/LjNX6FIqAunazO15vT8opCh3Uq8GcOsp7fVpzWzSkgVsZnbnPir1N
XtUxh58kZrzEp0HsUwXGZW5bstkpztl3cZxEehcr/Kskr4G2oyttSYOtOmhpUD6L
3l5IkdwrjO9Qg/U+cffRRhMtI71x5+P6WjxjlqAw1h0vqZ7HydUzaj3w226aF4PE
OwOxE5G4Xm1FHfeeysJw20LjVVYKua4Cwn/4rwcq+GG6Rd7dm46kXfrOYWcx0uNg
tZZqtP+arXF0tn88v+VI15uDix1TsDmXtaPk9RKPjpqmtbV7OSAI+En0UOcBQ+lQ
ky3mb4vTep9nYF+oCnjrtlgxXioW0IHkv3Nj53zygzHGMVj0Y7naHogGJU48H3+l
j/uMk14w9ym8vW2Vu/aO6aWuH1OGYfjsB9cayX6U2E84IlGH//tSRRNG8wEx9u1q
qJjJsJdNZawwkU5NvwWIYGfJUDpJZigD6HgOXNR6fQIiVyDc/xOt/eNqKrtQSwKi
eB9qycblqZppsN8avmiULY2tJ790mfa7Df1uCViANydkxolQTmxkk6A9CkpOiS09
tssiQexu05c914cmjcZLJEUcCGi0MdzoRZxKSRdeesZfGkMS52bO6eb1D3bBaf21
BdvGdby2CyLA486L10U5yvLqFCQAA06WVwMtrpYFiaRjcT2o2fOpl+eYfn0bGtnw
wOBvUSWfzol4sgoiHlBv2kJ1QPx9NczUiDCp3gZuPw4zYPU0zWrksJOhTZo/WsKM
iEulZertvpq6+ADdLoI8JYVXOoGBnloVoiWtOlVmj6wMAFGsFpo0BecQL8aypeD9
JVrOZZBHPfPs5yDJeyB8kNnw7tOPUqi6R7H5I5MCNRJ1Us8JFYdhEdxXekoOlyEb
MtrC1xvFKdfCvt/UvO7wcSA5PD1qggxm23ICn/5eBkkSV11q9VgJnuVvp23ldBQ6
X6taQW5Yl2sU24tC0MUZ7CAJ6jx48Kz5YOAawD5Y5ySPMotoTzgpuRKe0wu8IhUu
jBq4o/2y/9hJr4H+gYSkvKsVJyGGkbn1MO/LD/5i9+jKSKeFoJNQGwmDlHQImqMp
thtL6AMjEBzT2qKdiHX8S9aW4rrZmoYM5COBPFb7tiTvoaVZK79kzvwzuCU0lWFt
w4scQxAJPDim0HxFuXV//HVdvKF2nCt5gM4OXimcNkwswJw68wqrWJP7BiNbmmaS
TnCxJIUM2etHRO3vDEQcMIZc3Y2oHlVtjzFrSSjeuA+Zx2QSMJyPMfI1xdgRMtx8
ryP9Zjmd3xD5aPkK75bAMvjDzYrRzG6prAqaQxr1Su6wVRiYKS1FMJJQLdTBQmaQ
94BN9B29JA/IJRNMcFWlTzPa9VRScGSWh8N8BndMLLnKujp0blzrWLAaNweiR/s1
C0qeuHEl0NH/BzaQcO3sv+QBQLsGb9ghbJcZcozCyaSWyNmu2i3zWHqjfCbG/7p2
Jgv4HIgzKPRbgttG0ORi0QiuyDKHw66ABl8aJTz7pkJQJFZrUzCGvPsx4sSMpVXw
6bRoxk34L77CcnWm7N9Cx8sapvMi4YBTVfHnV9u7ZOzPCPvQfEXW17BSzhTdJDdb
+ROXfyzA/XLF3tIgj1kz2sXsz1IxXdLIDcNknRanTrPiN3EArSMHAAiH4hzXAFJ7
KfVeFjJ5L6rmCETrJhMqAHwqI/Gbc24KE3uZPOVcnqcBmCdw975fyWmvijWI0YtV
sRUl1+q1XVLMJ4m1qrhHuX8Wnof5uGymyhSxWH45qpkeDeTnz1GWK5HYhaKh+hJy
IOrYGdYuJylYS8ovDM5qczRqOyrF8/8knBn76lgPHN8QL+kArPUJodG1ffJSYl8Z
VlDumc1dfWrvyWBneNGl+yk9Vxug6wWGmR5r9lWC6IGkNnP5x8a31Myf0RDE0aZb
BYjeqLFGWqgV7ycvHnyeumGfM+awk1fWYPV0VE6WNP6gkTnnPi0GJbES8thevObD
bHiSHnpMz68om0x8wAbTQd5ARkGPIScK1n8g2XQR2adX+kjStW6oexFezDyfqV/W
bRYIcMSy74Qmq57vhZiyHK2TuSPoj9RHNBfLUk5lWResvBCrUHkkvkDKsT3xp6ZL
Si6RpVvsFVh0v3dIY41lWvClelBQLM9tU1UXGj6WizFki0a+hgzir+TdcoJYPxuk
Q6j4JVR5YUt6xVxGEer/4Unw/JNhv5GjgXI/Cvr7ZK7EcBLIg6cHiQD2pO90HnQd
rKT7As2XtESyiqlEqO8/+O+kX/N8rWfhJGBDkta3xDEWJzGJLRnDpnQ+cB5phcx7
Q63khKq9uvUl09v1GOUvSUgYyxd4RnmXzI/ZsfWRfOLW4rpQQgO0pJUzMNe9QyuY
m8//tyl8f2Mv62uMSgJljFx9ESBlE4UOY8+rpwTBiNQ4Z6I1W1CjhQ55zhK+qFqR
7+N3+SYnAcuUP7p7buX7q5LZNGwY/E2fBvvjYUy4lsqTJv+Y4DiwpqdbpoDwGpr3
EVi5pAZzTQPp1l8vT4eOPMmnP+cRc2MGXGlvkeENbur7dRy935hINaoYFgOdmsa1
TPr60DnVm2OT5XZ/jPX8A6ii7DxITOHohbQXB0RuxqWlteYIauqLgrOClfXYPpYz
b7QB1BMdK4Q2UCrUcrMkk8d6QxJ4prng/rjcMihztVGk4S7vstMeX34yNCNYZLZM
7TcwbF7ECGNbFpXuuh9iWaz0n2PE1W/FroNZaG3CkKgMk+r5zmEAP0VMV0RqaVf+
nz6Zj65REw1crJgRhKuegmJMIM4k4iHa4jtWSyjbyO9wpYkNIodoWgslVhIKGv79
LCPw+qJCjIVo4/CqTj20Xpr7RP1CvCK0XVitEO4aXzmnbFuTJeAKa2ubwTwmLctW
TwnMG4uCblrfkBoSSxeV3YZWNcERMuPya23HJTsf2WOhv59xGHQSOQ/oXRwq112P
0SaeXsSOwHGLtfdu6VsyKPj1H/tRVHafYXbHmqXtFIn8tivHMXlG+fHH02cd+g7B
wW2Cqr6dz1X7dBFUpVvE1MnBG0IPBHSG+G9pTqS29B8DN8vQK8xUaMlKD0lQkV2Z
cdWLkKgYh5AFChGpa2gkPYvxsG5KrTd+0gjQuSMWukEK5hmG/valoRK0iulgkLZU
vWz3FmLMUllDEfYK3U0kDGM5YEvhVwSAXgq7XpvIoc5kljFNVD9gu0LA0+6TDqHF
DQKVaS3idf6ozVp9YbqVQKKhRTjdioHSpMd7Ur2SiGwX++u7bO0/2inv3MVC4iJe
nvbWtbG0vneWbISn+Cj2R0rW1Bw75Y03qvz2P2dcpmVJOvxfyG6OCw0V32pEz7Ks
+W31iA/f110kZ8aeVEed1JOfWSzp16dAJYJSTXckdTOo2AWNnIdHVWJIi6Zthe3a
7RIZkdEC8OVk9dZ4hgqKQX1n6dKEZGiugMDSnE8lT8DcgWt5byYUSn3XK3lU755/
D8+PBC7f8m30qz41lNjOlXS2mihn7sl5pdzK+1bSVYk9dKkJji+mSZ4iOlETroCq
U72S6Ik9fuUiGbXw2Gt1NoYvPl5XDbL6eDV6QwvTh7QYWloWyC3tZpWCN0N18SvB
Jfy0uv9l7K03KpU8TLKdKAFctzL90C/FP5EgxELmsCDpVBVeQ0NEwE+RZ00xEBOu
kCQ1J/+RaFzQZ+kQe+Z/l2EewQXFbiiprdhYnoGjcc3o+h86iu8T1rtbhdrJ3z5Z
nNt/qHYdw3j7Q2xM6TvYQESHo+3aUY9X8r5OzB0Uior7JpJetwoB1jG6v9WjQ/xl
7PFwiCx0mEQgsD+Pxse8McGbq0Os8Nm5UeSq+v/JB087PEO6wZjsP/2H2cgvoaOn
6CHXgi4QGMre4ZowOsZHVA/wdDXgk8yy2/vtX1PkmXKVuAA5wiLjlmYlHdmpEIx+
+uu9M6HDea0HS72FIqoqOHyLoVMoJAnQO/Yc7GYkQxOTyxDCa96q202xTXKzH10+
9Ekhj3iVT/mTEK4nHMDuFWDQY1ycs4fWi0bEMHJubhux6Z2NE3dgmjQ44duWBcOe
yr0I1vlzmqiL/5TmgqiUqAs4b6BXzFbVwiKLuXthltCFXDoOIqCE5cGBjhK82cdD
OmDGt0SaZBCHy1s4ebUTBr/HcoRkxRZURCrmR560B6Ly/31FydSlsHSddsx7/N7R
Nx5FAUrY9jmMwimorMz56m3z9S5W2OCVjtjTbetqYBbN4kMpy85AmPoLjv4YXAaC
vUF5kSi1x70KhcBDLrPWHo9R9fLevuWi8c/FXS0pSu0+B2N4hM/mBZzu2D6po04T
rQYCQE7AETNqOLnROP2wmc5uUYwkHcEIruldoPZ2ZLtyiWBvNMPz6wQ5UcfkcpFV
xR6LQgSyWEkUTJwytp8hDkbQOMs3GeJhg3SFTilVGUvAYBdCT7aAsyUz+6O9V2id
BfdLUmY3pWMR7WX9KtUghqrh+44rWsTkPqJFSDjFZAUyt7V28otWtV7UxIT+9xh7
G+ddi86kE1B0TR8P/Tibl6pE+OwQUUgvqufyewcSBMLmcubTnu372+e2DAcHIyk9
NNEuL/xCRFZf2PVDNPVRyLLU3GAuhEOBCGbLV/fDnHiBfRp2tynRUjSevSA9Kmyi
VR8KIKzmRmatO2jW6xWdEiXIXYif8Mvgwq9HJncM1YcqM+LOeyDCKe0297Bu8kbV
R/62Q1dzzEuXA4GeoHWAr0jjlK8tZcwknHIZHgaOiuP9g2BkAyRdqiZ84/2rKJNC
bJtsn6jprBajI9rbV7e7BtBdxqI3btZ6W1J+N6iZc1yJfM9+QS14fWRayJDY4Pfd
M1kGfpYDlOm35BrlIzkDSsQseYGyyCNyfvF52gVxUbPawwPsmM/0pTGJFMiPcsay
P9oTpHsX7kud1J/UoAAYcRhWPR8qiSbqdc0EepjKJv9rgiHPv/bvymuYH5NkJKQL
kFVyIbO4gcSwt0nmR+TUGsojhFXc4TpzDAHpoecQTGpI7CH+zWno20eBpVdxYox7
B2OQmsD5G6RJD2DZLy2HJdL8b1hGNgRnO1R4g7ueluPef7lq7hyVp5pSHO9/7uxj
V/yBjURhlL/iymO4/Z62qM+oI6UqBE9EPzJaXDySrBc6qBRQWf+ldPC4f5b16FvB
nPoVQ9Iy10f1qVaGcnszKS1M2wazykp74tRd9JCxmjEFmJPQ6mYPXMR26Tu381Ks
dlJo2vHPmSYCG3QhsI5A3t1+6e16/6QEWFBlkS4S/IvPpLpBtDIs2T1YEqyLO56h
53jJc/C8EZ44OphjlnOWMuTTkVzvMC73BrA+FyyoIdpUOheh3tMorW+NVrD2rxk1
ivfdOIp+A/y2gU21vrdUUhrBWKYWoKlo7G7hQZzI1XlK1Miqwclmkkp0AWqQAdk4
Vy2y0W07TN5wKlUZXNnsTcvDzAVn44Z8Ba8m6avMq/jEX59F8fUeTjMqrIz3jomU
PJq2gWjdstxeHddDnDm3++nDINOwwpCbkriU92axwTa6Pik+5VRNwkHHMht/pncE
kJCj0e8+Ltc4Y//av6+eiLh0VUP9pILARWewISMYZuWaiYuju8eU8AjmwfEYv81x
oig02hf/ZlTUsF9YNaBnoZcCK121sZVqqEcUB5d4+/iWlVifS7qEC8P7Exy9+17f
y32DRMw01HGBqcQWPhOR85rFfiD5T/sAmZsGX9XmEohNK5Tcz33B7JXwb7GqDxb2
Eh4x8VZrIOkhvrXdoqIGu8rR+3oTT3AAdYYcUTuB3DNU3Gv+dA+f1rlrr0UvSQH1
iJhkB1KrIrRSy2uk2wjnFc1z/4ekQWa+wcNZEvIxsk46fnFmsakyL3oRvQHiyL/z
dLU5cJ63xbpWhDD0Jc5RHrn1Vnkh1GgDm8u/MKvBRnsaysMfCLz0VR1DBX0GZpUA
/gx/IdIRJfPiDZZE0ZUohDmYes/QOMCTZbnrtWuieZqgs6FebMJym5AFAxaNGHQa
VH43mfmb6IDmgnO8QkOp6IjAqDwS/9F42//LAW5dgcHP+Ua7R6pBMwoPQySLE4wV
C3rorF3e4ItvypMrqh1u4FKeAIbNP3XWLvT1Cy3QYRO6ywKjWMzW+AQJkveLFF+G
Edvwet4kKfJawq0ixCcyaDS02u9KDlUwW+dtzRrQaHeOquang7Otm64t33Kfi5x3
YSHu39XB0LdvBzQyJ/BRSuY/ShZhZfk+Uxzn68FW6dMKoAKZGWxPwXfZYkcFQugX
3/hj1yK9n3wq4qqvzpQOkQ2cWTb4IqIbOAyZGhxdcj7Tj3Yk/Q161UgYJSib9eqB
rmm3Dsjv9lMSfHASnz3dyChKeDNb2OqRofp1MXLeEqLDg0yevI9DmieX8lCuX7fI
UeV2fuYRAbm+EQTNc1bVL5zcoR++ecAIzBav0LoXDdBXPte5Y7mesAOgNhyX0A/q
3OCJBhoEEnzHpjIPMkCRMsIDUMPVsYcg6qzF+W5Rmvx/A6jS0L6FPFI8EB2+SC3W
K/pvezDOE93akQhVzajtK20XNn7pXgxQP8yq8wVDKVyn2s9gYAgZeAQQHNnkf7l2
aTfb7SD1XWrHY/vcyzyEH3mcTvLMQ8oXFN80BnaScEsCiZmGnryC/VXhduWCdH2r
YD/PQgUC4wnwDAuNhvElqjkwib/AChZ7Ct0U0T2cc/19Wpyi5PTaLT7LnrqkcE66
dIe/39b0vCoppcg9ecwWC8IUbWAEn3ccvZpwmvpxEDpQSaWKA2/0i4AZ9urexJBl
kO6GfXzqo66wDHcjkEO9rFmnxwCHEJT53aPUGBm9SYN1x0sihDZtVeD/+KKRnExM
5Lws4YzLlxS8UPQtCfv2ovdKm8b+4YzlQn1z8z19IELcSJHPgARB4NbmrZDxYIJl
61esolePlzV2JXoe6/PS4c0bM3CLQIwzQohoHQJgavtHosE+aT0GsvfZqDeNIKmL
vpK+9QtfknW1YcutL579PyX8JvECKYVsoiCKt3BcoVl6Z38zp60nlYi3v4UVP2Js
4pyZAEXevZk3SGldiNoRSJw1L/mmx+tVW5YxTcy35cpJFYNm8dXYsQyln1opWTfy
ZUib4FGrIe/NXtR+AbIaTuMbDcdqwoTnsNsrslLKW4FBoIydsC7NRAeUvm65g87u
SdDq/sBnyV6oVfk16/101KDCMH3LNz0T+Jn7mDu2wevOmOwF07P6sR+sNPbIvKwN
OpxAC9QHdgjGzn8/5eEido8gqjLpm3N4eaqPPB1U6XWkt863LggeAaX9DXv1SgZX
RAUNg+vBQe2h0EatXVyuZWMtTUXY11vkjARsypY3a0blxIIjTAwbbDqamYdmcK3S
M9jf0zor4N8B5LYGbuuEBIINM85GHQLtJIz9rrwhSz3/Ic7ami2JQtHRCCXeyHQ4
XYtJZfQTdcCf74xI/QFSmrbUyrvc0AcYclK/TWE7Tpr+PhBy4CQw8Sl3c3Q8OHGu
nXgAvBMpEyujBdMC2X/LMBsC8zvHZlEhPyKJuGYLLpkvXRt+421Xyq4NwAt8NLYj
eIas6WnOhots5tHq/bX4rrd2zy7Qg41tW7saeXLzUmCAjZuQiBAFov285OcgO+1q
N3IwTjhnGa+2u4NW68Lz38tpZmARx5fghB7GwJMmYL6a+unsUNsdAZcIqSS+Erum
zqsEMk5iz3rvAX24FPTdQgScmMD+DI+hZK248EhvoF/Ml+ix+vUOAj0zrvrRQHb2
EwtnL16apqNYSs/PUBqrcxQZDlmk71YFGkaOK1ywNHk7Y6/49GH8SKIpPxOJLQRd
Tz8xdxqDvyAq0yVLJZO4KmtLCd81wbo55WxXw8Iy11jRKJMmyU1MywC7xz+gLG+y
RrVGexcCkZ7eRmgU3NgsHG5H8pV8rhyMYEvFh9CJaMvqEs+3jSf44EBaQ45O8Rob
m3F/MQaTf1sUVZson+kdVhffoKE+izj5LG2fNV0laeBTuM4ZjWwd0dQg+MBNkt+7
v6bxypSu59ocq3ZojaGu4ccIQDgzlY+mUXQBf2huPBRnbH6nspKb5aXTJ00eac36
KZTaqeafwMFuE9AMJufitVaOvUQVEXwc1iUNvDs8/kgEEBqankQsO1Pr4hK/Jbmc
AXyvmXpDndW3m8DskgPP625aCRmjlmWkraoBZQC2fNzwfofLU+djs3lU4rMXXn+I
JnqeE4CnMG5TPXeT53ZeMa8iODVzverAbxXFtvi1L+dtBpPbDuRZ081Eegx49Dpv
9GmGlmvCuvc9yPTfn6mn0VakXmb9LMtOiid66dr8zoPDvygbancn+TnOixgIsr0v
dCNPvZdpUglDhyktTDWcWoJx5AbIXJw4mrU8JGvnARl8B8wrS/YD6XljMqMScoFa
Yj3eYKvc+ZeMgZv4qmRGcLBOvwVpJo9A3cfVz6MqiZPFOYXiXq1zYhM6Up9JS/Fp
AZw0wL+MGqzuDyil8wyjh+ys57w4s8SkDz6KG5vD8CUGxUhajjakr8yxMjiPwc+n
2aBygEE64EXd1Cr7rY3QdiUgzkiV2cwGnFQisQWQy9G3alrdVPU3RQZBQjDh6Xbi
oef2WiVuff+c8TRqOyyRK1Vc9UTjQsbg4AeG9cNg+beCU0dXauNGg0jGQZ2tLcm4
mqsgSYDgGb6dzS+af3hyI2mEWMKkuMirLsNT3n8ZMr9XEtgLsjW7HHkYb1RH/Exh
6g8huET4nmyQftXdSlDQnc/NXSnDovZX5cmsZNTA9I8cf7Z9ykXdK43CuHTi0GsZ
Hl4Si1fvmO9Ml1p28tq8dy0SPv433SsUPDbwW32RG724cKNKk8OZ7nyfxJQo+Mcr
DiRlL6gX7LfTDwMTvL9KecWpZEitr9mqGntWEkd0W/3gZEm1XrjSYCljX9sBN/5B
uRIc9Dq7jwwLztDOo7zFIzMFk0q/yg2Eyc7O3xm4Af8EFhQZoa6+In+vG+bYgt8L
Tle4crwPlMFRPv5IxtzEjgH2hIyBgwU2Sb14jl1hrIkjm+Y43L6sBO9CmDQC4IGY
scl9K4VCY6eXIR0hDA0tYuNa/yz7B0xXxuDXRHja45XCy1++sO61r38Zfllm42w0
77AA22u0ZoMjJ6JtBRwZo7QKxvIZVMXRJsE2OEtvFSq6/Uzw+dggP1q+T8+XTd1Z
0Y6GS5dAjrBi7ehFP5qgMCateanImmC+9oyBKpd7jMSEb93nCf/t+uEk8ekfgEom
ji+uwmzV0sP3Nbu8Civd18Z+L6kWp5a+R7wPaLCyO7Cn5xcY/J8PM9p+vi1lcFNT
zs+rIDnxCmifBrJZZXoLGMkxhZI9WJHfgnB0QMEGTo5YfK+2HVi87gIAos/yFFyF
jgCT5xCHRhouQJNcQlyTpW4RVuToSiAhy2VnDu4h6FV+eVciPcEP7V/O8xyP6QQ4
/G82tqPo52i+1EFdX7zXUchEYXHgjFc6/lCtvHxQD9EJtr2t3xAulfManAJ0sSfX
1Q8n65DUWWcg5XIQiM5wc5wiia6GDGc6HdwSk95E4VbjdOha1+v9sM5/GXpdi42Z
HWBHXSOkkaWjvBLKwY2jscuWNMySUVXqSu/6c20p6FQ1P6WMT1tSjuE6GczNpSa7
V/0x/wJDc/xRtpTtCvifTMC9fyNJhBejqA60U1yPznut66KbLg5M8vNAIDdj6FZZ
G/xkV3+pkcSYoMJhISfdgifYuFSvo482wlmMGCiiNBi4tDLvLH9mAOWZ5LC2rhIZ
T+Qp/cejgGUYlCetP8RTdTORezJjKEdLPdbM2lO8LCoHnraUE4VIWxEHEPx0EdsX
n2EOVRoi/UuMvKYXN2MQx3MnXXh3MqRPq9tnJm4pZ3pBlGc4E+3XR6UizlEv8A0+
pCnWfVI/e9806YgSscKVT0v55rhMO1UKcZPXEyK+U5DpwpMS+oKLC3rXm9lMhO7C
RKrGqEn59i39hUNVbKykRRC7r0gfGgSn46frANL/Da9R810nZfzfycBfFvjBJ/vU
cIj9jxkk5rc3shhxCeBktmhxEE8j7ram5eDcqqAT+TX7WN66H0NWfOmmCa0xIm7j
FNIAZyHpJ6FcEaRtWXgFcdMVXlwWa589gei3P29CywJ7Wu8AOcnbzeSMv79fiToM
Q2+nMWq84tgrY+NqcWi1mydh0MgUEIRkvGX9u1u2r3Ra0J82so4ZbcVTw/vWniXv
S8khPqLm9M56SieipXomdCeBJsPTaB116tfiEgEt/FDmSYFiOPkrCGXOSXxBP9xi
v8x/qfsumXMRZtE4Mq5L0LKx968MaEpkegj0T7RjjfzOb4/DSYyMFvPaFGnQhXDH
3G51HGvswUqRsOIwlCRj77dFzHlDjWGCOck28urc/9Z4HXu9hsJ7hQYrf9soA+0g
eLWK11eTJ092qgpqnalukMGv59DIQN7uEaEg+rt+xVi5gLg0RjdJA85j9KePOXpO
4g+HQ3c3U8ICKQ96Xgbwa8aV+wxYp+0O4OhD0KL2tPIygBtGkLC8KMHu2BDmOYKr
hYRM/SE2KyqP6MihLQ6Zomx1765UZzfZSCtgBOoQKMU185MiFexWLPQIO1zqiF3V
J+muCA9A4ulamt0qNdznhwC3sK+ft7FvS7VeAJXr4+DcLAgwJQv5I410IMx123V4
oRo07eVPQSgsIcf4UXD15fyIXLZ04n9bW+QJ3Yaktzcr+r79FyxHf6O1qkNsiAxB
OYbKhMlu/GHxWsGNCbZ4NXRFiJJAjsgoIS/2dYqOajgFmBqS+2NHGUBdSvfuAeO4
OgIkJ6MzJ6NcfMzSmvruVJo1n74z96aE4h592iC7CnqfCYr0ToDHKPMw5qRvNc03
lOs27zCSwg8PUeN2ZWtlHpZSH6mf/EN44zHqjTwC0u4uP04+RZzbaqcUphY17W84
l8rqR5tCn+9TrETVd/6U+0EI3goqRCRXM/22d/WRXzepOK6qowfovG1j6mJ73O6G
7oXm+Kb7t9W4WNny8IeQ2PSYxCZx2RypS8gbtLdR2iqMcbR8yWN+Ztk1nNWQL9iz
k0HYbLPh76sn8oOFnCzIdeQEoftmeIP+9Q5Hrx3/91RGETfmal5G7SCdJbi9bpUn
iyQfQA6Cc6m+FTbwZauUmxqdA5Ued8uP2NzQ/itpI5lA0vBegLEnmyWIgEtu66Ia
Pxu/SsYOLiAYhaaF4nEeaPjb2ezzlcKkO7g0LLSbV1n8aqrMJQnsV1Zgf/3uIKVe
4u5Ze8M8MUOsW6RihA2PblcpB82mgFpV2hnhIvqc+O2DCQbmC4R5mZwzhhvcj1rI
Cu5lXWfD14gSY70vYgWqHAdHRpKmxu+JvJ/N5xsGPM3/ZyPIgD8fAJruMopvNA8e
/v9FW1mqE+vCOP+ZJU7eGXhJ5QhHDp6UlYwceelCnDlreKN6ZtY0ynJba3M1/LX7
lxdmZTV0DAw0mIcSg0VikB02KW7oR2RDCio81EFvQfM4gyDVHrp8t9O+78gPRp6t
IYfxJ13HTNvn3M9dJkC23ck74n9s+PNwWxdP5U0zk3Db8ohHrpMmGQwpCmHUKcqT
v41C6p1yDKk/oe1xPoUdL0HzUYwr+N9Czw0N30O9hrsUAY2nTvprB4XsCiSiQG9e
SUGXZ2+YJgU5UlGAaBUqwXrKE0RbGrw3RRbNpgAO2EvggR2X6r66XH5ThgO9wEyH
CeAzJ7ZJu9AaGTMPpBtNeEKpqUdtMVydhSPcnrzb91Ispo4FElMIBpAb2WnW/zcz
UQN1JGPWAwg+gTpdBxVBScv51L8BCkErsgjm9rLtAD49WVdvbxi8uguwbjHfmAY+
Gi0EHJJobjbiJvPtWyltyxDc9AV2aibCni0r9PGLc7B8CCCKB8SnFfiUWvrR24xR
MNqHOm/i3xLwQozMxojTf5GKTZlbvPskCGn98wiYSGe00EFzpwDK3ujjYhkSydUD
uoHEOHDE+NuuqHg1HR4HBUWHJ+/YAnmZIW8FBMsBVUG/IkLOTs3pWhHTre9pBgLU
q1/QK3lPlf3f1q0n5VA7IntCGV85xaFqcUbvnEpQPOJqu+sBa3cTrCUVcO/CiTAm
fMOnFAKBuAV1xsDM+eYFDfqNEb3IJZPC9CX0R4Ff0qKp5bXmEQQWvS4Kx0cMk1b2
eanT5v48H59O3ETIsgiETliLOrUj5YwPfEBZedluBSCxptG4aD2PkR2LPdzLMqgu
AfU7i092hkmPQIE6HME/EjqwiMm3c0u49MHJ4VAh25A6g4f9Xu0NdjavQryhLnAy
UCwEzRmsH/VnuJhtRUzaLdOXqLpO6w1hJxj83jFWJ9L4KYRZ4g5X6a4+6bwnizKo
LW0/SY0KA3mSumIhPMD3t7a/KDUhaP8GrSFAgutdJiSCLNy3GkmmNHmMhtiS+oTe
e6gUZ7yZE3e7IBEuy7zkITXKy4kR31kc2S4gPgXZ1GWATS8F+LxdyvfDnIXs8b6j
8+TyyjrG9CvXci3ttxtslnEVPl5LWxMxKCbvLq+mW7PjeqV4fzXIr/sXZk7iKJd6
dHOIcurML1Jd1TBXCpUrqCUPoBtB5q9Th58dviwheuS/CTYegmm/b83cgl80CBop
hiAW0Wk3GuBV7CG6LvKfU5Eb+59dQKjCDAq+OZLhLOKmCl41jHD5n4TSsTJ+pDb7
CpeMfluHqzRAZW5PyZ1xd4Xq7hPS4ajPEPZelM6dVutMF9ZSCI8hcjB4lelv8lIT
aFqEn2LS+EoIUu8FB8ZA/OG9sOxQ/3rbwZe9F+YL4ePlqSXVNnVosTrEPfQ83ogE
gyZBe1r6FnJPhYBXkuzFmMM6F0SNaf4W3B2agnX50Yh4Yz5TDWxW0Nwt7TGL2ICT
ghJR5P3kwGs5ndU67Vr1tQTJKrQktq/dB/qUtjcLwZllIdcZ701GxIb/6VBgDBMU
Nz85tWfaUbbvwtr7Ss7IbOml/AvDHzK/xMGqIvdcyCWIhrMwj90E2HEb+YJO2I7m
fbXKEUEQEtZbZmcLMOCaWKCbPdfI0fEWCMuKr0U6hsMgSdEAQzB6aewdITBemzUf
Dy5f3yihBj8C3c96tPVDMUfOIIswz44c+oOUlG0FGjGLYRgRN366SzzsOOBFd8u8
8LsapVSbL3SSIi+AiOX8mQsenQ/IxedXGc5kpeuoWMiSvgr11ervC+StlN6dtgqZ
y6ZJoQGR4nkeYyoAmINfmb8kZf1xbyKIo7sB1cVhVC8v7DvtCpuADY1JmMvG8H8y
5MUXkawM+b3UyonLmvDVcMZzRbrQy2DHViJFV8UtMd6rElutNtA/WeaV/DFoykZU
74tXejT9WY4no3WEpi7PJTNsIGsnaBq/3nRowObNZTIBRMC7bwFfrk67D7fMjnYP
IuLP1luHUvtD9S108SMUcFFnA6bpwtSw2G2Q1PUdZijfHrwLUqJQL9bmBWq9/wb0
iu6CaUpn8V6BirLRSWNlE2LrXbqlNIvad/brURgRrAh9E0eetW9eUgZh1QlVSN8A
Lwigk5mpO6hNw8KqAEpJnw/TiHqFOMP+8UBgXYzn13LVAh/kAap6ZKI2tOrM7YN/
x/KFUuFYD9o9pQthUvX89Y19Cf3yJPBTclEUOrAtrFzS3Hh2U5qsf5aoinSM4zc3
fIyFZsiNrAuB6grpZD9F5BHYi3PnvTRQ7/C19Pg+wGdkIEygOe7lSJxbKwNSKUxp
YDSfkvfkNOmAZ+7PouViAX1YZU7+CubPpXR4E/vjN75cWbzRa+H3WpKZMH8EPTfI
4bo0xiW6CpoNJrtCCApwERrZ/add8b/NxezrCNzN3EzUV1HFhrJrFe0OjV7Ctz+2
i8UDyaAxTzEw4JLWd/CdiU5Pya4sZtYkJD7Gz7t1CtpGYOikrHcQQP5Tvr0TBcSv
Iy5mtJDdG7uFRIYHk+2zNdj54ptxDKGpeBBUQ3TljhIlcEbyjNFjzBvX/vBrUE2v
LXIkPDYZmD709tKW8YoTV68xZ69RsncKgOPfkwUzUqw9qQsD6QFonQe2rMm3Lc9z
FOKT59WhZ7e84F8WHZF4ZrLVK6hgQ7qcqNguBUUQpqYPF5OgJ50NXEEtSGj9juS+
9qJSRBVHzLYQReZrR6KH5iqmaPyGox9iaS+QVk1RE+FiUgXEH11VwV3Mn1K8ICIK
R/W6KzPP3Z29SeRtZI4fTU5tqyBXVsDwAYC8PCPKTrofW2G0hXvKJwPXdwlGEPDa
2mq/1T7Av4m3l6HFIJiDADhuNrlka7+hC7djblm8UqnoxRKRuMl+Xw0o2la62t2i
Je45hdxyp5G1cX5unf4ZlsqhjL1Q+uwdLw7QJlrPN/tNo/sUskBZvX50llVdminM
cib2rCesn7nFTPshlyeB8vXDnk+SFJ8FcM9yJW/un4r3x+QVX1+wGYChW4oBi+1P
z1/tPYPgaOamSSpBMXAx09E5vO5TRPxdndnxrdJw3KukLwQAZ09WrwYNbCO/U09I
g1r9RB+0hwLnJf4tBhpvA/8Zhk+aOQhK50brS8RBTXoqj8FtOOJPw4hBsJI57kd/
lbZ6TJmf0AerqoESsHfyxb2JgDbUC5oiznKLV/dCtb1r0w+v7Ql3VYx71ThCSWcb
zNwu69ORE9yzu6t+ENREkFSz22w64MIFHaF2/hq00gF47r/2T3EMRsws0u0rfVOg
FdMfmxaDn6jFhdwzTrPFUxWZ32JCN8pLjapINx/ouP+sSLnewKLcVoJgydzFs1ox
sw20XsaoyxVAHfnuF7GGSs8iO/EKiaNhB0AiCnbEHH7cSzj3o35KJHvKrNwEvYRj
HyuNBGHUh5RGevvZdhccDUC1r4fE5BXzGCZrYk4ePG+hrKDaYgExzCG4PBhJ1y5S
/R/DtrynBUx3SLniymS7dKvzL2HKTZ+fMR6LRZJV4SQBqrvAhUHrT4NoJ1GEkld7
sHZZ6WgYJHUYBV1J8yNRi5AbIDOlUL3iae9U5H4Yuy8ygcYa/4PBKFuQBIRtMKCc
KPLcwQRqI9s046h6UVdCNi3gf2ye2Hu6vhifiWJ1QE7YLG1ooiVjCVUv3XsP4Ide
eBcPyGVh4Ye1zwqP8lOJUkq1CDSWUrlc2m5rQDd4GL0GhnuE+8iRAK5VvXK1ESrO
f2iIMM3VTUksESLdxMZYNI8eWav85ujwVox4aNDqfbp3gTZn6b9gtPpS0CzFl4+1
hkxXu3cK2hkdXOtZ2Xw4zQZZseEVSdUnawdfqsqqHNw+QJOYhItzH+pYS0r9Qj4A
2gajc1WhCOJlIyLXH+K+jnwLGqQM/ehjM0sgGHkn6zo/rDxIYoo4BWwa3Zucu29+
EAs6eCcPU7QN2Rutj29JFNjrFrAjB2Wp9FXuK/p42NUkyRqpFs0iPtvCbbXuqSOV
PdkUDFlTZoWJHyLk3WwIsYpqhuqkTJGdKh1uoBqv7nZGhkvVddw56auoiBbeqTFL
OTD20IbVIBAyX0tsJK+FNqBJLkzAZkt7si+XKhVadcOKC28hcXB6Vf5K/UPWbikL
D9Sgf6seGtQuapT313xTdY0m3Wz1xFjKBi0EIqZMsRUNkrP+OCV50RP4D+yxqCbA
0pK6CEoU4bcewpdjIbge9i4OwHEcOxtRlsfAkezKjp6wnmywms71ABQ9tgh+l7kK
y71jn2/v0gdhVDTt0kvh7dWTveWIgiLBoCGoQw/ftYIXZTdpla7mfCFQBDRD2J4i
/wdZM8Vqt0LjIhcK64FFq4sYMcUV/+isYpHbg9GWYy+Fneln/zm9Edar/56aQcDc
peSqY9E6legwzru7LhVNIeT1PfiKSssENXmhmi8U2pqdj4ouEfqrdYgueTBcJUf+
PLBrgcko5G9P9UEjvennK70FKnyennOainfz/6KPfwoEP8jgQbNvvBYrFB1TCL6P
+/OfU7kd3HBEofo8VUMP2crCKzoZY5Mu1ei82cbH74bzMREKYPICCpJa+sGga4Zg
woj16etIKLC8EynPW23rqdDyKJnJIYesyno2haHQ7yzo3MBYtv1eVESS2ugw5+Jz
dqe6+gwHD8r2dKShV37r/64KjeO9dPPp1VhaodL76mUnEV5Or5Y/nhwd1tScx54j
f1NKRGwP7P9kUZBgGcFmWIkXNmWUroJ/WPEnqcmKHJkDDUvdLivgaWuyqDopa1Sd
9GK1vLWbWJKdwACnPtiRDogCS8zen2ktN+b+kBYJDDUjy3T2iuqms+qrNIgqNZcD
Mn0jqe8J7Va09m+t7xvqCodiVDhnTvvHOEvbsYBxiB7nToW13H2N/pD/1WrPv9ab
sVxoppUhg3tf9dSr4hXu8truc1y5g7Lslant9vqEa4HJimNOCi75ypeAMaG0RpV0
mDTIZy9GrmdT+RKuPYH7xnZJ0wgfcjjmuNgaW4gnyV9wAiqt473a1w79xEHGefgl
xEWc3AJHUtR4P8eiJTq3s5qUdJu5+6zWu3U5b4f1NrFo0IwXt9Dslbo11onxlR+K
hoCEzID84pCfPGilVAqZTEBPze5VSlRy6XhiOOCvca7AXWoUdQuNXniWOe5quE0u
wQFpeElpEId+qw2f2SMI7s06hca//WVYTHlriBTdFfL+EMBTTd3ya5l6umAt0ZjJ
dGeNOjJ7URCYzE+b8zLvNHAAJYyChAsz8h4WpWnQU4FigpnXxIuM98R1ci78QKc2
6R34u/ck2FoAiCPqrz4n15g7fbbb3yVOS/1gUZQdjZBlYbn7+3AtAWviM59afask
hq5RMb4x0dIofY9gQcT7MB3+Ns3Pem9NEDrdCsLODGlnIK+6DNN00pQxFRs4Hyi4
6UKQpeGqqkYUHMKM8ZB4Z608RR5CqiAKs2g9wbZjEKoIn5i9P9XY95pAYXJmek5S
tWuIoaDMI8LRrqCF14/3aJ0z/t+pt5sphKL6snzCkNz1sTmyi/gD6jTRHqJpztsr
wEPOkq+ofMAwRMPQ2QYAupMa9QkS03prgPa7nQMYF2rR9av/w3xlGHmwi1Hxbgwd
F8XgMICbEQ2yKs35JDGKWZ7su9xHgbVtmhsQz+v0DYmIrasmpHcDYEzbrIFV3PAL
NNF+1VvUuIs8/OM9V+da2XjQPM+JCaT+xlTm4fCKq1KalKlclK4fHrlj/47qcQqO
z6hnmXWDK9/JhBqUZNBwUrSgODWTAz97DJilMknTNcxBG82vTO7YSgFeuJNTSI/A
gxWUeYJtRDF8HuBevsmkG/dqXn39B/QfX0/ALIemDzFtVTZ+xSIhQhl7WIksTC2m
qlBrE3VQzHzkYMaFSO5ZMTbgTJkd0jV/+CKMTNLv34bVj31z7TSt9SLQ9uK5l45P
rJqHnYJSt4fs+TwjX5PDg4f4QggHELBLo38uDOzqEFOFdQFEAz/4S0BDa3YVn++t
HBgJwHJRXgnaUzpFRR/SefIZVFaUjC/vkGj4Em7OhVk7hDbyh/YtOusZi0FTFMW3
NAxD3++blR+XZmuw7bUU/nWD5kfpnG3ewuKgbfhZ5LsXZ1X5IvVdFgjcWRVtmDv1
POXEN4zihmisd/zq3WAKtbh+OqlAyMZIXpIZJZHw9AbpJ9iAX6m+AJPM1A6eBhpl
SIhjXn9uytzX7S4Q8v6D6yLAX7w3Vq7frHbh6VbpVKUctpYLvIANgRQyqq9cWnY4
TrhQT8T+2EgrFgSqseKX934E3R64ZWG564aox1FOYASAfu/IAmUAv4HF+9gWLVwS
wSB7mBGRXDN6pfg0SEqgep1gXFyz/6w7yXoNLJSzFSgC2rNHgsDWKdnWcVl+rTBU
yTFK759Z1x+XBv0nE20MPPhWUGyj1ioL7zlMORXA2mPbshS+OiSjzk3Y2UjbzOhJ
2ASlnCzJvZEPXf//te3Z7P3bZhOVVDe27Yt9TXLqyWlMA4JfTjQPBsafIr/cKvyt
3DFLCqxS4YU8A4pQH9RKwzCVm+UDrQDN9r13o8RCIJaWN5AyvCkgaDJwsvdnwro0
ZThu+NIq2yKK9Z9mK0JdDpC922mEDrA1qP/7to+o4F1ttrpOsToRKbRIq0p2CQgQ
O5gzNSdPoVA1Kh/nbZMSnUXFr+ME+Fq7skFO5z1AVN8nPt/AZnec8es7VM4CzMfK
ZI7DoAxeLjoKVCVwv9arOL8eCbradTE9l4RacVmxDrl0ZoULISrUWz/thF3224u5
mh48F+2hdWvmtR7dmOquepKIrzeW8uS/jbcHA+hQZf8u4zqRIe1EabaQguyJu7fk
ZpIoyVL0nv15ZUJiwBdhy0LBdxzCso+5kNDfarhLSVZqVLwDQp0DZl1urDnNHMZW
BvKtlp9vndAxmg1zOYJg8aC4j7I1/wQV6tK+8pkixdXgZY552LcG3o09BdQ/AH5d
q2QvGDpp5EOP8aGxs8xlmksRZHv5Cxu876JLnUTT0WYlxJquhFqYPCwkcNxYRKwB
QPaJ4AORe16sutZrhEyAsh0e8FiDWUkkoza9UpBBstsoj1xZ6Su+U7q/dJKFBPp1
7lE7aeiJYhs16CU8cJ1tqZfWPxR0srB1xonKHbPL7sJeyb3jo8FImrRtOm9FE1Se
7rNitbvkaFTSE9G3DaqropIYvvnaQlfSa/MMF/k+3D7NMPeBuT6tbVMND303kQRv
YQKJTwwbOWFipVitXW2ZhGRSdECs7hS8RP8hfmsLxE9ll4ri/jYT7dcUwkPDYm9e
3f8ztaVju/Cc6627zz6dyQss5WVyiMo7kspxNpB/eZEiX3kQ8W/m+zCo7L0wmR01
YxIhJSsdMRL7MoPJGu3h7DVNHMAL5OtKc3JPqMD5uazSCJWyNB6Zr+b03gm+ih+V
WvekaYZLl/sipbhzX13kNfgkg6Zu+PFUFncpGP0ZujORJYc6nRo9OiU0X2/erCnz
A60la5q8TdPRWeDyDXBhstkEBo8TsNYGusL9UnA5jdzTULxAuQE958Ip6BqOmmqp
z89fWt+3gY1nfAMu2U1D0z36mxpwA3Pr206Ya/vb9UXlyTBvnLu146IxoFTTrpAs
3U73JtIXrGgxZ2Tm+gslPPaC1mib9vVvdRIylaksJgkIdKJwFZuvdRD7od8xysDH
i7hszc3IeEt9Hd3+1MoaZLJUf/s779Kr1vW4DkbOQAYfO5ocQfeT4pCDlOBMvmwX
1Ess7HxKvWIyRIIt7aKxQVbD+SAwydJLsyEB99Zmq+y41JmSKKuTy1eJW8M12Kbe
1phwBhMEMJVJi08TdmodGEMtWMMIU+Ude+n7J1A8SZl8KNSpvuHwpd4ZCO/4i9HW
I/eR+BzBawLQgV68fz2VKoVArW5IpxMM5Lf82BPcuE2V/QyLjvytoT6t6W2+2pue
U+nI4JhCEEfIKYFn6iHN2ayyvgyN60duz8ZF+tAZOQUzhiW2ycNPP3bjeNXN9wQJ
zcyK+tbAcqTcngM76W4kDBYNBvwooSbh4+2Jn5oWI7WqBJ9W4b5ycWw0gM/JXY6G
MfTNkqEXEn23c5rGTX62pWvFgql2CWK48RVVQMxVvhj0VddIRFYSgOM3HT/+B08m
UYB80o1XdzEgqJTL9+zhkNGdfsAgDEnQ+YJ+QaHsS+NaA6jEImYPqiHUWXiaQRgl
TgELYjjZngwDkW2kwATSVmYEdsQeLhFMHPoIE40no3q6J5bRFhPeHFuUGoiRU78X
lQ+KREyh651Sg5onACiDTOYdOmfYyOp51zsOhV1U4m0INfgoyNSVj2gaNslw6eLj
vObkj9TkRfJ+R71wisEzAlOjVWRnj+LOVFt7TCyY6OPcS6/JvA/wqMmuclcB4Hgd
5pTB0mykm6+73hyWtPISimpXJHroO/aFsu7H3MTKslPfcTXACPeUXFuC54zUVYxi
+D6nucWVjvEHBct605Xw7S6Z5tzNXGMORnTVAzIxSaAqpeyHMSwTFxj26yS1kFel
vy0XWskozExbDMnC8FvwuYCfzB7gw4y1jAKZc53nxPLcBazD39N4gCPp+9aIKOkA
AsFNQc7quGhQfbkFdyvM5WniAbkPHSiG3mwpNl95bVx/B/suJ9DgZNYcznCpb4r+
okwaUeeKQZIjEPF04iBXmJWGqXEeiKOzsRgID21ArBi9j3581WBEeRevB3NCqbHg
OUjb5eE6zmqDLv93qHUqqr+uyQ9bQAae3b37FjzOauMJsGkeSPrYeQEYdYmZhdbP
AGnl9iZ6CfySr71e2AF59JMk/ZVVBPRkXMY9H6j7lLXE80A+D7CF88BC/r1r8KvV
xu2QxNJ8AsAW0mXqWmR6lVWl63JStarAXDSMy9Xyran55YAcQUyTWe19i7TUd1DP
SF5Aq7pUX7V9qGxn9N8tCVEDOA3Tpv86Z19W63dtuR9nToLXCHyDmQFcMLhRwbBm
Cqndkg+fe3S3QbFUumgQaKkCfYrfTyom8VziQz5pfOY85EWyan3dSvw/KGsXmnAY
92rB3rnBZ9cNSzr/rBgP3DH6YE1Hd0xsFh+sDkW6EcrwtMNoSGW/MW+GtikBh1iZ
os3WYaZpU7tLAF8ZuRbPSNnrC1EI6CzvX8+EISunPqCr/NsXdnf/yFecV9b1k3/0
dmRmG7yhmrSvkcRM6MCWp745Y4WA9tqfOuPWuoHh4aDHLSVt927QNdZUxyk1nnXi
rqKmzInTx1mLGCDuFL6bMbD+7qaFVW7BGIYwsh+vYmcy7pAraWeWXslmr6/8dXKp
juYhD4PpTFiMmZrE7LSrpqNum1UzQr3ghqy+gJYHJFEOIi+SUvWOixrLyk3fdPcR
Ejx2vjtK9viOZrYLFS8DUfsxDaEPs824fVqJYcwThvy79qMCd2CawGTTZKbvTy0L
whskF/Vnc8ECEOjt6fMAoiKkuidCfmOUnQmmuSjfVLyeX6xrJWAi3QLgqOb0SqSr
o+/Br0iT3UfIT5MdAeye3G+3iqP0yVnuWGt5vQciBJr3/J1BH6l8bfTVEnP33FX1
vhwjhlba0zb8+IZz9scGKjIt9wrGB0Xgijgkjw0v9JaZoiLlH80+SHkGQZcNeu1W
S5yvPLMuB/F5LGlGNTuApj617CmAFGBbfPBbfOkiMeNDS7jMhU0lZzONAiaLgu3z
6pVDtOLkYWXAmo8JbMsY7Aqi0TDUMr9FGPPt7cQhq1pWhKmWtSW7LoyJsZ9yertI
/Yzq9n4p68JEYT1ZueUu2lcQqz4Y86lro4j80PgxkjtifgApxsj1zXjgi9lEGWQ0
M1p8Z+LWDYMde1gLrtU9YyhoZIuC7EX9k45pI4GBIyEtTV7auKBeGnqRfbvO3FZ4
NirwsO/Hm8WcT8pTKslPNmJj9TVWE9vdaslIZQCQA5R/X0eOvy2miKPNUBVkuPtK
tAGrB6kQd8BXAaeTo7PQ+s+CgPGOQjznVcHlSOKJJ5FChXCj2Jt8Cox6MtJv6jp6
uDXs8OKF18YQGaQIGwI4zV7ytVbUsNAheZyRkKaLMS2RPq/Pwx/Nd0XuhQYSTN6X
KoG3xr6Fk1nXKNk9gr3T23sQ5CgTNaok6C6xWOt0hsMOfBXWm9Uw3ODTR4MYWtIK
FxGE7rxE9H+nO0aYNWV1D78vxolsbOsMnH43UfcZwCCsTa2JNkBdw07+T8ssU22m
OJuI8A+hpRuW/KDMk4m4S5FAeI9hpqv0EcnOHl4uHPzPRe+Nd/FjiNy7AoYPf6Pu
Ix1VAstddGEOFk4f9xWA9uQT/L6cURw+4E1AQLo0BAJVQW84X+/tG6SpDfI3QZcl
TEsWn1vuTXvIYmlUSu2JGTc+dn4vsclxSPltSYky0FHk1kwarRecc/5t+dkYwG5w
PNdWkBHtvQ91uZzToplPSqjZV3dnpXlyZ+MKQK5jGiydfHBIm/8vaeuK0hCMetyY
0cAKeJrHWoD9qxkysrHWTUagpOoWm0Tv9dxyW+sZmGhYf4fyNKc1/MrEJuu4cgWs
iWBHiZ7fzOisKYm2SI+zin46euWYzohpxepYxEuyoSU7JkfHujxCq8wxnSHNfb8I
US5xtAk4iETwrqNKN9I+/8bJwyHIKDC8/Gy5UIBzZVcHnj+BEPw5CfVgH5qcLeu9
JwaOj4tH+Y4ta6rBKGoI+lE6nrvrhW//edbi6m4oW/7Iy1O16hjFlWwNUVR0/GD4
Vv4vDPxNHI2DyhSthxbEC4MDv6b5B+UGT0LPkZpKQL4hrHKk3EJpF3dTBxddJWxi
qjZ0HREfwzmeAnGJoA3eoQAY5kO7LquE6fBcYusDXFv3KCQy8C/0ScSAQrqzjXaf
7xPRAAoQK+SvzxoRrgVLk+2P9jf3EtVxnIZvr6eV3iVJ2kgzRFs5XjYdI3eiAnoV
h1ACsJYrLJ8EYJxSiFI80mZEvVX0m3W7fZXU3KsJxWdfJNafEp2PaR7LJKsaB6lc
4aezOQZILb5XnHb9/8iet036lv6KZDtCQq8dJSsA5S1MgJQ/mFsNkbjc0Z0uQmyl
KhTHqfH3aVlUCMovDoK0i9NKFVPdtQNoEICqokkainbZCNdkqHor8gRDQgUsXbj4
qU0RVfDoYXzZSYxNbqNi6H0bspuhKoi0EAkADf+xyU3MMImrk3ziO2ELGcQPv0ly
4KuNsCs8WgJNp5RrNizTsJyxAyoYm3sew0gJXsjMlnlrsAEdZh01zEvFr1euMj3C
PnHLbdMA1CWu46hPr1W94GHxeJsPX85bCH0ePbdf+hdSdakavt687yxMmC4zP9CU
r149vZbqXs5fxVHy4p4vtUhoGllSMxrwjwAj5lZko1LvuXgzGgL/5qBKRHKY0WZY
LUmAzfGvJZZUQ0cU4hzFoHbRyFN+otF5UTAcpkqBVaukkgNkBDC7i9YHs1hg0d2p
yBftrNYOwudit6gjJ8CkM/0mDur5UWKYeiDBC8hu63SvuEPu3hIJksWCXs4EXu73
jALgKB9LZvCovED6MPc0t0Z328AcVannZA+u8ehkFld9wOhd3H0TZg2wANQerjjm
8Ofa2ER3USBCfzPPlB5VA9V7kfK3Vlzqi6sGFEjMNhX28HgQyI/1XrzZunHgnb0H
K5yBypyGCwciA7mEakzDOG6Cg9/u1+YQiQt5KG9P3AXFF5SJtxTApFXZLSXrha48
us9GsiVBnzGorJn8lVER22Y3HuXFai0VPwTrtIqAEpAvMya94R190mAaerXuawui
KL65hR1M8p861X+yeiFlmvPtnT3Pd+40QxaqSComIAMZursnN48GU7zNRwlr16qK
46BTwFGsPPibmMBg+0sD6JZHP8RbuSWc9gRfoLA6bCvAH3Diu6fVDWcYFt7ja6Sb
mY73sHoMFn1C2BycgokHC2g6+hG9Pk835t4ZqHbLzYnaeULBwjU+lEb59N/q2nsf
RgY7g//IvSJpXVy1cuEZPdjHVpJeMfckDoy27JA0b1+xQBmdm9zICJSZJBrX2ee5
sv+xiLcgzKp8HnJ9mpDbxG+p0ASvDbSlbK6WWHmV3dHwE0QRDr7qTIFGzWUTucwN
OBR6RPMaSSN3I1kNPtV197wVGvby4wRK74CjM/nAVYHGrHJcbTiceHuHv+uULxLX
tHN9huLgt0cvOLlAkVsBMGzGPKHSLTFRP0znpcxvI556Vi2MchyCRBSAP7gKrTG5
eSEKwbQMwCrd8psCnEJkf1OFz9Xikyrgl9aPG1avqpbAezt7g7u4B4/0e+yMobPx
gSnNiyPM4Z3/e1de88kGoSogybzDypOZlIpk6BpCH2TnLpfZQ5tQkwZ8ijA1UwYj
zJ+nAqjNZAJC1SV/sIL+n6hG2eQ080txIwtDR0qePTh/vW8aydhu//qzBSCYruPJ
uhBzhKsfym3GKIGnhg0ZMJzA2gdFbwBhdfY8FhNXPiicACIjiC5vhod0MDQpzauf
aCKSPvmuqV3Sf78YhlAhFZ9qkWmRKoRKuZYXQjhnnjIif5zxOzPI1vLyGpLuJMun
QuK57brlF+7aiwEl/tZJZdqWW2lxUov6UYxTPeSVGLrOnQlTU68LUEyMK6X4HL+8
LwWu5BwndWZBtQ9TIn6MuO9WG4PPKynP+EQpL5cSZc6Qi1HMAhkC91PCRKUua8qn
Nr3wk03Ea8Ikba+69zT7Oi+80cfvUWahHUOCz3n+LFE1XBrr2eJLCVjYWnpVIuzH
7+V7OkjVAiiricU/r3+l6jZZxGbqshZBZwl8e7zmA4zy1Xy8Xj3CrJg1kA2EXI/d
XwbgEWd6E0Ttxne5Nyl7jbrMAtI5Tt0Ov3Jv2eNY8mMZx9QqSZ93s+ZonBMs8pIT
RxR1c1TFLemn0ObnWurgnNQzcvaLRE8z7Bvd99bJx5c3qEsQFwpY0bzQMSZ3Sn8K
tzfjpt7++oZD2sjmiFZ/tYTcLfgjd9PbJ7QVpPgp9m/XkG/E1yp97qq1LxFvLutS
ASj16LXrhKHqdR7xytNArhxrkFAdG3PX451ARk147VpA37rv0+yCd5NxUoZu/A5E
oYhWQ5WVDED0tQCtZWE50Wz8Zj1dznzzr7fkDn3/Hg33SJlv9XJ5o9cc8WpV8mUy
9KBS7HvwSev+vxS74q5j+fg3MK/h4a+LniisrLdPDW4BggDzYhUwpfRiCboxSOqg
EBAhZJPhc95T5FVkK8G/MZ7k4dCuP17RlzkSlNRqxzV0tUcLdDVqgHWLWlqvOPY4
2ODjbXPq+1mr5D9N7DAsvokIPQJOYhPTnaX56RouP5aOCHoGNmSpDjb6wz6dUl8W
mqZp/wwUd2u/mZ3GmmBSBlJ88OyFNCg8xDEd9t6YCWQEAw2iMsdLHGOpOga1CoTf
EStkO8JawK0a9c7ZMmWBDWjo9U+zbaP3/xF1Ha0jk341wWwN2osB/r/gU8ZUrX9X
ejLKGraRk45Bc1UkVbNEQMUeQU45QBEzG0jeVl82uaJ/gdsC8lhttH30Jd+w1ho+
9KuNLVNHmaxxTx73dI/svVBzXkor20bKhpGK8QSHrMustU5ZGbpi4Ereqh7fSzlV
qPjQhVsSWT8enuSuihidrXMa1FeER/rCPqKtak6OMXGXqCCO6+HdgsnoAfc56aEj
pcSZIS5sXABRFkuGG8IJwW6Z2rkGoZe7C0DkxHmkjgY2lhJnamRRW4dDBoag3nAf
u4/U0OBOrYYzb4X93Hzy/TfztUJwm4S8U0lprjFrjmFtk3Au0Vp/dyy/8I6Uwx6+
zBwKNaDKge9lUZoT5HAJs0t1zhzNE1JzMyHzFBcAURhvUb0GZIa+OT8POgm1ThZ0
xRkE4xTAa6T+MCz4Tgz4tV/TvzpbW3u8PzOecByJYjj2j6s42Tk2jGeLqp+rmDrt
4FT0B1C/C7x9Cg6WudgyHxa5QxCKiU3Za4hDqteICnLZrN0ZXnkVOXFYTM/CUUkY
3ZjsVKasfnRjbVXZH5TnD2R6o1j/CnilDRZfx68wFkP3ZrZQ0LWQaiFV3XPfjYTZ
eEG7O7o6p62XFTPOftyuBsc34HYzKWWMicYq9wlV+LEkfWcT0htjQ3uJajVlzG7M
2DepjdCyrHmws2uTilfsUahgv0Iop1dj0WnWqd1zr9AEmw47s44RxH/Y2zoZ/sUW
NZ5NbiGHKa+w8D/ABb6Ti3DfgNzg9DLH22ZN30tvH1QzRX0zU66/QZvL5JpVIcRy
xgY89iQWUkCdyOxrZ/CLH4YloguB5Y14dbXhudWNf6kM9FP+G4D5+2JquWV8HjAS
7pfs8IX6gDiew8dbYEu4nToE8G3qG+emT3gp6Uwl2ftWVyRHhvX4Z4aA1/fNsNac
NfrdCNJ3Qi+QhI2uf4J5kKtFPf4VOO+a/UZCuscZJLkUDhCbth/MzWKDpiHvCwkT
vnfDEUmrUeN/nfeYxiADw4TGir1OMJctrBXOUX72bzKx3gwein5i995+JHOUiKAb
JnyGsDj9fFMA+iKmRDsuoYxIiDPopcCSncUOXlirq4y2mp56Hd7tZANRdOcNPv9F
SOuIqF3yMUOnnqeYqlbNKP2NyQvtB4vZ34sGA/z4hCtZRhuB3xfy+sQNpmmzD2pr
gvO4cv2DpdlH0sdsG8e2yx6wUmHDrolybGYFHcFDGqZni1CTxz7i78GXRQCjzUn4
YMJlPds84AhTyDrqYxQQuBjsbsY1GaBi+dGpu1oQCYzzw/J/THWMhAAfx/aHWCnb
ZqAp7bnGXS7ichLL12YncJjR5+c7iAn/+ox69FGqw0mkA+1NsXmYlOY0Wku345XX
wJFA3MQiO8eyZCHuvBJ/swypXf70x7liUXwZswytC1qx3yLNkB6+zpMfthSiEeUy
IcTy8635k0Dg+nMWWsr9COSyLvSFyGkEX65L5xHurczPSjbCfWX9kZlpVKgcLjNq
XMGb8Y0YDvXK5pW8SbLDlIMShBtL5NSNaeLsK+0m25CLJEK+yJphsPU/gyIUg6lA
HdR4AwqYP7VFKuj16rAY8Jd0cyVHoB3LCUW3cbK6CGhMYXSHw02e8/XfQSt+iRvX
jvKvJ6lFZrUiSucUMalkvoIvtv2ogV020VtZVCwXLmtOIEds7lP83hv2vxIXgqjU
ZpfN8zeUnMX5c2lduw88nMqhjbujSHEFz4mPyxQJkubKpYY/z1vlL49IAT6nwqDp
Hh1SImc3ToVByuQLqGTSX8qGSUPHZA+7Qey5Z5Ta6MEBahSWl3v6J4U3nb8uuExV
LTxJYYDNHc4+j3Jeub2PaAnn4XUybXYKtR8BYiRQ28FGwhvtamtDU5ATygNSk4MZ
HGk4iOFYPeqOznEQY6HKUsmXuZZMjyqJYu/UjkDWo/VafOCAnsmMR3OzEau9hUG/
ROLSQiG+ko8myI2ERHiBEjFBfE/p96WMsaN83aBWBBq3VoRyf5fkPRKHTlspdd88
BN0rJIsc0HkS68lHdh5e20mfZHGi1WsvIsX6mG2d+/FyRvYA3Uba9bqLlXxrgDZw
kespmYcf9m9vAWjZ3pagDH5Rcckv4BSJApCpifMoV2/J4jovqhlVpNTIClQpYui2
sKTQ55W/8mYi0bmoOcU7ay1pVMrtE2UD1iIFnn9L8T9zB4VLfIn1nZcDgdf9qGAK
Yy8JK5aYkkAE0U5lnaBnXvrEXRNswVzlWA+Z9IUhekIp9MwHrY5onlOPY7iXdSNW
kQJxbCuKVnUo1b+ogd3Vuq6htfcP0UVAW+xDkgypXvojtXGyuxIBhidQFes4Po8N
xaeC+z9IaGYKEX7ZeuYI/wTsUmazZ0+/+F/PfZa6IYPiPc+Q6fPOinIAsDxIXr7j
yefwK9QAruMhCtmOxyj3oDCOH931avRHYj5xENJUmuiVK6z2YZmDz+WD8RMZHjRz
8M0Q1Moo3GTvELsmILbkubRa+j2w8je2FXCCfrI3Kyr7Q7Ajj8TzTSQuHRp/7dGz
LoZ1voNHBF23PZsHJAqpJiN5d6VC6Nqr4AUgTrKsyQmYVFZPcarc1iFOH8HY/rYm
jBgtxC4Xze1mBCUDtAhZ+/U2D7vFML2klSrtZn+SDlEF5oH1CHeRzVOB+MAMU1A5
JN5BeaL85qbS+OmRWTed8HJmKoKmlxNab+5JVptD2GUit3wrt4uRtkAd1uhpyLSH
EWBDih6DuO+UMnC+Gn6S4rrCA9hk32AxL4tEfWF69OUbuW32w0dvJ5r5fS8OeMOx
pJGwKaW2XwoOS5CtNWq6CmzYsXGyTj68exxQrBD6/8DWHYfIYmqNnTmxjj+x6vbF
qdflXOMehfXg/8txO5S7NSslE2WuTdu+PZ3SMi0mednordAx86KUqI6CQHkKR9W0
2Rwgl0zsXRha9X6TQPR9W/s4Xif11lM+Q0s5zsxnUdliIl3Otkzbc7AuA6aQcRCm
5cZCRE7o7c1+SDwI4lIQ9nGHPi2YwCTJCC183sZLtuHqwxfSRu2QiBHXV1qqTbFk
hSErS0QGupPzbn/+Y3lIP9Flx00eqAHtkZzW9xJzTjux1+XN+tr+oZY1FxPqDBev
x2lKZnKIXWpFmFqPTuCP6fei3gIIt1NV4Ujh2ej/53oWQV2pMS45vV16czrwEw6w
d8vYTPc9wr+18fVaAd12P6G97w71TfV118WEFEmDIT5tH//WGZZTXYvTAI7wy77E
WCnCgRHGmhmyOOMreJufWiqRBrXqBsvzrnFKAH8fmo/sUT60oAkcKHqxMTVNkL2A
XsGQFUavL3WonIf88Mn66LAF99SFTatAtPdepMOKA6cJ1nc22D+XpP/cEkgRezkL
DNv0W31CKsSkwDStc50Z+1jFX5y6V5djFV6Dt1HeJh6A1idsTcM2mexh9uW8FXk6
p7v7MU5aMzUnZuE7Sgjr8WAZA/xFQJnpKl8nOoMPpLpLfak41UFdAki7yCA22XjS
XixMKRBl0vcnPGv6zYRzg7KZp3sLndxNCdau66RTpp4AtGoYdUrRZkRDHGwilfLa
LogzMo3+VshsD1d/hKpVcWiFHLeh0LMTaYC09Gk2xcW9WZoTe6FLxxsyqnDhPmTp
8tBRmYpZEnUYyH9sCb3vnLT976aj8RbfyMUCCpqPNl2+OBCz4LZzN7+fR32jf1gR
dzFMTAQnFD9Ee+KhJGOfeVLzOH5cCdE0RASdq7EnTcmR3sBpJfxJOJR6hguq+6ER
AfVYmEWj92+OXXqg8rsFW+T+PKkvb9qx6GXzchnoIvs67yFfuHHvffmJbH+S0BiC
j3+ohGjghSSiY6hugT3/nIgIF1GBcMXcLdq7qEWGAVyYJhfRpCFLTD01meQ+kb+4
oqyWmStMJWXhHMYIspOHA9uYCDZmeG/Iu8R01Dly5wRAavyK4uDq43c05zBzTZte
Eo8RQ5dbddfZ+kjLnvgaLKhAF0QKwSlbvbCAr1Qt5r+WUPBL8HD1h2xCCcuvU45b
EqEwloENeiWpbqLSJUJmAUih/PsCo+gk1IuXNG76ZQJ9RwTcIsyZEs/KxRVhp1tl
JxUCifFL+FZIrDQWhdHxa7pf757tr2yGZqgtHUWtFVIwfZfXTh38ct1Zm1FtdO3l
DrnEC22V5sDFgWbKjDPn6fGMoaq2skXxPBdSgiIdRBRJzGPNCWspfOiEiVwjgla7
SwnY6FX7eToa9RKJOFwQqJH/d5rq2QHH8hGlbSmziNiv71PMlMvLzL3FbAdB3M7r
CX5XMCi7SvVP2JDlurbimu6B+5FmoZPbeSeQ3ghNja+IwzxBJ8gDRnnXiG/cuE6i
/fkrpFpcabDjuUyCPb4qj/xo+hULBc3y4BRP1GVR3NaTWKLJLIeBbLjMP7xVOgNh
ryAyvQSFPmerg9qDWnnZ/lZCje2lGseFg+IdrkUI95DLc5s6pyzRI/RY/CSCQA+2
hrtyx9PI6U3qIMOE6uwEIAuPXY0/+XFkm5EY5vxX8XR8SX9YSiE658mB+D7OAL9P
HlQ1KZClBRZTHNBP0UdxAHY4XQXG26bUqKfHlvO+VN0mzlY8bBs9u/foSmsUH4hZ
zMDpzi7nManX0TmqxGtMTlWEIlhOaNV3TgMLpz47SvS1nCKnNAUsjHsIlVyeaoXG
Gi+tiFLNdijSDzFzfnBfoWX19EaRMntTwHyKGQYCS3iKWmGnxsuzf21d262vCn8u
v1kPAYaxQU1HWOeVNh9Wy1hbYUHm9wXfn5kABZPmSCAIiIdv9WClLYEAlR4Uulm/
SIj7+CMD5tckVvSzymQkRpS15ui/qhsbbHaP6q9UxAmLCO40Ly5jEN6QxNXqnTAv
7tO7Z0oxt+dk6v17gTjhdEnQ6twh+PQYUg5GU2MvoTzjRtwyfnlTl99HqLvzl5FX
nz7pMyg4OE3FTiqKCGUxiAxIDjGPzkJHK5PYDn3jdZvqjFv6FyGGS84rZGddH7db
pfXU3l+9rCvZKetip6e9GVe9xWLmDN/7mgbMjbQKeC+0Td2MXGIicJJtfX/0s/A+
28tImF3LzslXfODfSZBTZePS0kV7c3VqO5ZpBqZ/eGP8Dy4Dg0jInY8Z/BhgkxlA
M5sA9wZamatnZJPNwUfrxp2jQLSEYRYW8rTBF9bx5oJSkiPvI9CpJpTlC2RE48JZ
gm2Oxzctv7jaw1aCKPec8EUqbSpElWyNAj9U8dxZ010DWqL7fV8DwDCwWYr+xa29
EDYPsVwm0/NP6vqQmcaiqCjM4O5UE88gjdPvhy31A985GanI7UpzJPmcgM8mk2DI
4rhj5moJUfvlyi9akSeCWdH8y4X5tFX2JetCdTGdiTQOQOBRQvIrFzgIcJjtwF4f
AVrqRZvTjja3ZVsHwMLjm2VXqD9eu9+GYs4yvpHlOoe98r7AAqXQsoiRzJVuGbKL
etpjnX08342owhRZUK5TNdzDz6oGDKhsuPYxprTckKeN4VYuq/9EHtAQJ1HVOMDj
oeoGjySdto+XERvKZcmyp+WNKk/HOzxpp+Cr6uMG3WHaU5tvaBnTKC/q0htD+EKg
lEcmQfMMJL9akH88h5YyE3i6dZwci5gHVRMsrakuVAc8FD4A9+FMLybcPvMYp7Fx
fFW0cf8gsrl9R6EK/T9BSON7itJgEQX5JCpLtJxYR+dCp2i3QbZvig9aEvhwGFoi
Lhg3FErtl0I8ViiX3WR8SA0OCedXmrtBpgu/1CdhpeVs0BWARABXER07hVpsfCcS
yBLnnXSOxlgm/Ms2FdeQQ0JeMc905zZhak3NLnNjlbz5Mu42edOpL8QiroVfqMER
xex/cKb3y2uu/sebHHAycQbm6hfLHucnIXRUXGQ1bOPWesMdtLNWifAm9qdP/2st
HoNcW+osC2sFcLGKqUSUeGryWqv3zI28rWdzmufn+vSqu2/2Go/wMlbZ0Nk530YT
IHm1nkxCFf2twU2oPu2q/1ZIhAm+u/NN8KeuKeWstSj4XMvOpPjBeNQB0ogA7niC
hYby7PFq8MaY/lql9L5e5PUs0bM4VPxqkzoEN40igeIfpHn2i5ABJjqx8OMGVSu+
lSWC6cAXQ2+GmB+t3QNYFLaTCrrwZXa+5QVWVoocW0ZdTy+lLblOZGTuNAkTXo3O
ORrywNBhqJL42Vto0PSPgWGS4kHbGOQw9FIIDiZlAh5ofPJs00oKyGae4ZW+uaQ1
j9JLUgAQ7dRvII4hSXgGydzEX/e1lkwFaiFaueTegCScywbpMz34yJB/YQqHmX4b
QgnD5muKoyCkBxUHnbGg1DQniN8pLiGOJoi5Z5NTUA+DSmddTsMtepuTDw3HFGjY
2BCjfP6jPGghS/wvwonIZo/mEUqnpY0Nc0vAeO5zPEHf7hy1hamWSeDCztLeyMR0
73A15D7AMyhMLPnruHxwr7jbqlgFBQWG7mRZSs7v8Jxef//raSYYIVVhydCIuAey
RM0+KeUalhOsELmcyxB/hB+xgAgzjNHTs+Pd1CCyiS8dc5P/CanxiLA+aX/q/lFL
GXVWwdok/osgMoqcYamGikJbSzKF2NmM865D8oTLdPTAUKR6H8lefs0+mVV2KNBB
fJcp2kfFycAmNU7dKKqX/+Rz26G0yX6VdM/6MTvb9t4FhVujvTY6BAvJhSVw5fb3
cwxcErRF55eVlDVStiTK26JxQEAS/od8ruPqM2oU4Ri5yAYo1wqOdsCApPAaP0zJ
HwxksiPUh1rgFEL7LCLZyBo7OHqosl1ODNGtM/+A17EVZJCgzjeA1Q0Z1k+HmrU0
vBV+IdrR9yoHZHU+Ry96SkGvIAcAo7V+mwuUNaQfEM3a785s5aaFIM3+IiSAcCII
9fymn0bcSEJpb74NudZwQhXpn1u5y9iu2EExcIDEJTT0Fjo95pmU6cbbFRPeVnHq
JrEqIdcgX9QE7tnBbhfH+gUiOd9/FzWuEJOf7et5B24iWScwh1Y+lWw76bA+sCVX
d+fjUSKiE2BFMeDOyaV6eWcVY1Q/rgTpaZG3qsEUCEGigpBfLnyztSUz1JhVBNaf
T2xXTOkqCOH7/fsvYDC9Gxce8B8m4UrmQ/ymFALwYFU7esCTDXHtu9bo6fiVRSy9
wgEl7eTXYINSAmeVs74WoeLzBrh8iaOEJL8BKX8XFTQ7eMCuuZSjmAC2VQIJX7cl
LnM3uuan455dAIyD5jd3sfCcAcUYwrSbFL7/+s4M3OPtdtNuK7bm/3ldW1VKeGSC
5y6pAb0iWiUSa4gfPXoXKotLoF6nMbLzEKuWuO8TmSqURwTIJTsPM6dLkdIcWsIV
C/K+evKWSlxfXVzupaaZKvC1nKaUBV8KxVwrVkUMqnvQnlNWPnTAdsZ0+KPw62It
tB/bNxBOfpRES8ONe1V2fUZvlGZVhxkv11uncHZWOn+aNei/8RaBlduoivBNPAFz
DzlBEud+17YXcQ7yyyOPb8urP9gyyizqHoAhz54b1fGVVjFMzHjb41BZKxzZfOrq
X6CH0e0aG4TceN4tVlx7aAiA+d8BIz+SUUB0nwjLtElidydtZNKUaVXLum6RNHtm
bVJAYPHG8y67pKpyvXehPYxz/K9nmlbUdhJOVuWZ8a/plAMMXsr/9e/IIWsfmIEB
D9muB1wMeHyrA42h5Pq3I5MfARdqr8w7DcRtUrwaLXFH5H+iSJ97+beYXN7GBqiL
RvtTwQQp4/IL8l7vTpw1w3RUzlCysgR55uUXzZkT55L0vfzN0vxd1g2FyrLbCvXA
ychWEfC6K8XPyhixZ5NUCd8tes6aQ1UqSi/293QE4wYETVXgXWW4F2KknDkXy1v/
pIBg0prZoN4QzzpkRy2fdZC/XX0qIuX/psTLu9r/mKXliDIgqoZqBweLyog4ZWZV
ED9kATedwXW/knPXi8W52zO3DrEc+cXT7D63RKDRnqd3kqc8GgnnK0Iwjorxn+Xx
vncaALS4bJK/pEylQ+LYyqZpuyzF9MRAQZfBi4i9INbwPIxkoXtJWs3fxTQi4vu/
QRPtAQKzWUcsUz7bApkkjSCkcALT+3Skzf+c9laVKEV1uI0zE3L6Ox0dAgj18eQw
vTLOFxy2AZ5OpV9CyJVgQ1+iUIWZi543jMNFT9aWtdfIYE6DIdDvitJOYlVP2jNa
3AlD9K4TJugpmgISF5T5WOpWdUOh4slHnp7CtQVOJHg9efwcSfOunNDE3UOGMSDy
GPiR7cz/RQAczZLlZu7eIA2Q1ZGNQWHVBABl3gJgA+mb3nMZDIFLe+/Pe1ckbvXH
9ZCBXqP83Z916BtBGbeOtBT2hgPFgf6q//O39Nto3JHIbGYbajkDL5Ayon2IycQT
Wbo0wwqiaWgkAbq32Fw4Uhkb+K9wHJahO944jf7RqtqdWP5ZsRN/qzNXOau007by
iM7VXRrcPARuAXRsgPSqYmkpvIBbrEh5EUShO5Tuv+fGZKLH+XxXx+8ZkfCWh9MK
Z2qaUu5YO7/7z//fELe/emFEM3JFxBGRYs7IX4tX/GY1/CkIWWFCqpj48QHl9Ma1
QqCgmmMztEYoYzArnBfZNBMWosHC/6kwggshm571EapiKThSkZV9KHPnvxbIzc35
ANibf+a8GZ9YWiFD1GD27sfoLY3WXGTvnaaAJO0Awrl4GxkreTEm+sE0XTe0PQU3
PQbY+kER4rqQi27fwV1NeIkWqDlOTbpyN0j4NddPC1hlo3ZAT62fCHVvPf7/WqrO
mfqGJ7vELKpErCuc1b/cGC6/8B8DlYSQkgTZbiQ8x/8cQQeKRi/ZnVG3ApU4Xasl
r1Lk+k2z3z4YGvkuOGzolp0cKB2D1h7u2lPK2ez6/+Y98haZidlPBYAY7llm2fBH
kA9+HbM8pZRqIKw6JBFba+tCjA+YqwjNlyaF56GL/yXh0j4/jpl8+E8Jx0tTcQYq
XrwJG03TMwvb0dGcLX57+VLodxqhteAw80m+D5M+Vf9kFd5KsvRYscwSw7yoncJR
rKwQp0qeqV3qSa4pTP/862NO6qkGH1VzW+CgHhJ4uY06WJwlfjN1m1qaXaA7mM41
yTx7dztvPO0+phy7STqLsdlAiljQFFl5qnmHZDyRiaygMppXuBkpR2M7kM6JpPWb
aPvcYVpzz/qvr8X4SjRKIv668tw1QZkuF8Eb4RqO6+22w61++7HAR+65cy8N4p3L
R9cPcH3xlg8Zor4vEQQi2ZtX39xQWyZJnAckTTQV377qw/ldAa2iutdVqEfUfALn
+tIbX6X01brcekGIMEzfAAaKwHIm8bUUVHQjxE/zU76m3C3NFBBzVrvsGqy10ort
s7c3kjKjqqET3ENaalm9z5jXoQMZt9XiC93Tde7kbCYDahzSSQCVfh1oX9yamzla
2FCGqK0qUZjNOYYV14864ljleHqYZygWbgQTWRpcLRJm/nKod0H0ntz4ZseDrS1m
uZnbOHewHFk5V/YQEsrWdYhttyLqjlRjvu0fCJoSMyMPjyvdhMks/uYwFdgV3dvV
9POKZd0xq3QxRxoDMF3fSKWlvfrCcvsK7jdycVq5Sjf4ZynsxMaqgARxFdGOGQWv
/qJLZbFGLUO7IzXbEJjxqePOMvLbqGHHYclDTpEILEuN8yc9hm10g8DMScoFwV7T
YEyI7ZN/CUFeTuaSk0YFdzq/zYk4lDPaPE79iXuhKRKu7X4Baka1aPuaKuhcw++F
p0gHoXF1aCfCaEhPZ6PjWHwEsqJVWoWpBH7IpWLyb6sTeaLsdattgQvbSevMs35G
z1KURiizzhsqfZ6rlSN5iuy+weKWehjNfH2TKBOpOpGwJZFzNzQiqe9pvbb47W62
4qT/CrObcYDdFqYE+u7oyzNROANWThL0CGR+ze/R/s54s9FGEA+L2vh7yta3mmfB
PnU1h/Gf25SNmT1Jk8mCl3KUPKUnZqWjSf+D85KDClNgRjaF/kmuFIBRDs06quYj
pTT2jia/t7ZjWYtH00dwL7lQuRWWe2BK+6GpgYQjPa3dNAqzcYglME3gBh3z8Zn0
ndNNk3r266pQ81P7KkdTe/MhnbBJAEHQR0pP7olIW6EHnS0TcJID+2yEPbAeMJyb
S3OT+mYsaUB7icGEXSjIq7M8vU8QIZKSfzKbxJj5R3EC7MNGPlv15SHnDZFSEzEM
wSv4sNPssESbV0Qc2+leke8ackmQBh0LnHIZNuU4SK8kweUqsm1UgbPmUbed++hf
AssjN7yydoRS99LEJq9bSDD8wLaIg5WPXJwasF8D8i91PmLi8uVFirkdmLDdKP6k
9nxyMZ+66tUfVyYwe26Xmsenc9YvYtrsSmyuCO6rskRdzVbl/sUZVkE1Do910Wdu
lL54HDc96aL/p7CiswXn0rQo58PGTysC1kgaIRXp6scPgrmNP9jfNRaDZ980ymCh
hWHIXsDlFglIFQufGmvJSn+ndBjZYIWOtzlV4sxVg9XgdUJtKnKchNUYU5oXf1hS
Ek9Ok2cqGqGfupL0/Lz9iiYkzL8tWGt2S9ph7imuY3X9Jh5WMlWkWO0vEM8EET6p
KFrEGhxgBk6vO//ScVrnuJIEatWmQ5+JIMIPqYj0sDEPFxULCpHBkjzfVD60DTnp
6YFOyjBxK5AqZm4KsubNt1148l+r2ywQ5G+tMP4bZDSpZwTBY0yqIKDkD9V62eQB
6KAMFvvxxrjnA5caBpaJ6CKns3vE6F1yGEyHohsXTzpINh31syfezXdE37R/1IIw
ap9Q37RX3Bb5Dxc1beCqZogqlR+BCqJYGFpa02dDwvUYiDWST5ng84jbJaEv8O/Q
O8khgEGFytEr0n0G3kjdFh7+BDpMN3QEy1MhTR7VbtFGHc35kd2BhIZI3u6uezuu
cCV26iXl8wncJmsxKdfE/1VWrg2ktvaihVKl8jeMk1c0N+U69YvQE1lrPVCAIkIq
0yKBif53ucSqj2ye3SIPNkv8ol1mv/kVsudv4RlmFks9fenLNLoTZixtFu7z7QME
+WTqRebbwPrhMzbV6bsTKoV1fmxkx0Y+bgUWwagjyz/R6u/tTp3vKqvnF7dvijAP
5ytxyKGm86B/Nil+FDRan/8tZzRFGNyQBNiM+xz9YVFcD2qb0XnnMda63b9dRr2U
+iJdrxEtNyu2N3R4S6aUwqmSVhG7QZyxXy+ru/8NN9XEIlfl3PAY0eDI4kBUEPll
+WHne/TS40O5eoigA9/fzECVIERZyHzVHkzB6F1Fp6LABErz70N0n97GhoSF0+hF
P95Rb6Q/DScK+pQPZHcHkCtrsBKTXdfvJiRc9TWpU2BO9fw6zquzoXiqy/ZcChbw
OuoC3IKj9YysJnZJm1CP9zlonAUzvRhqeSsr154lKQjQ8Zbek+AxMqE2FgCKEvZr
UxJnF0HyAVfnCo7XAFlaYwapoAAcdDvluphwelQIVObYaAbg6tLsmy9CeHqEfhiI
GCRwoNOb38bpK7dTRDRQEgICikbI+4S9X/p1+pnczHKH9mJMqekmI6mAoUdK5/My
IvGpGIFWmhupvXKoD4Q/0j4Ov1aL7Ft1vPNFT7aiYzDlFWDDxv+GfGgwDmO33zUl
rtUQ9XlXsio+NAczpnMjnvHhYgIo4FfqFL1aV9uBSkwo/CapODsstGQequrkpBmI
1W6rHAH8gPTEbxkBo+tGFZASMgmtkYMdY8OqEe9GuZsKG5s2nK66r3geofq7lcDG
v4Bjs39okJX+u4ktCYWh8nqjfoCrUOAJR8Q6cJHHcvkoxV/DUlanPlIL2VZDmpA6
v4jysu+GcMHiUimTJ/yv8fU/ruQKuY4oFNBVQwnBigIMbTo0ahiuMkq+EhYCWEAS
eH7evKlTZVVDJYVg/2wOPSOUpsGAy5a/TLKBagnajHKZeJDDpuvYbZOB7pZkd0W7
F4gLHIcz4jVtTK4KViA/03HzhnRYOSBaFsfWIHlbWTciA2F6mx1M+CFDouCxuoRf
FXyapPv5JVNF59tksNB4prPmiZKCMknxkjVtk+VALaLEtGSWRDrz6jwZ2FjdldCk
lwUprhuur3dzkChs5LAG15Qc6L/fwnvgY+Pw2Zmp2NEStcmldkJn1i+ZLtwz19gi
G99bc9A4wKDTUgFH/iMc0Fe4McGDbZ5Xmv4oW3VdVPMBSm3Eo16PxkrawUsj3TCK
nJLTQxejTq0bypFAWx8EE8+7CaFrfaHdGQh0HCG/n4H3e5dNqQfmC2TP3s2/agcT
7nco5pyGohw9C3hj284D9QF6orX67P3p1/mfkLqlZaegMdzlk8yfiyLkp/r3Yray
k2mtnpHAY4jKZx9x9p49nAP07LoRaU58ze675fXAAFuDMuUbv/sXxlJ3zql0A0wT
LgjFwoPQBki+ajEmKNG40Xf1jk8+DbT/dIhGNMMZeQ9lOlWY33nZG/XVpT89md9R
DbG0/bWkWSMiM51tLNTMOXOonVHOqzTx0KElRotosLRd6hkjkLHv7pB6ywUikreL
9KBLfMi0OO2Z11um9aAvPzFELHJk7km6CbmWYA824TOX+g62GAtdf96puZzEQ5C5
3clWzL1qHpfuf13Ue/v2oDCm7auRgAvtuaPJ5yQaIVIB5FAgjNambAZLOiVWoSd1
4dxddP+K1gY/XhwIFVz6lzBBCMlBdzH6I5/t2q6D+jdARDDoIGVuZFKu95sT4DFg
/UP599HXMcX/pnh6oKQNiX67dC3Os4kAlyjgL9WywZ9psomK3qqgFrCKElKtztLA
DTJYybxKM9ClwCD3szltAAYBFAlyVOkvwtws0/vNCxo6ocSYdFD5uKH8OrnKt/y0
yVOBkOs7Cp9yYhOOVYjAqhLDlZmxa4+lei+kSz0YFK67LzTM/7r0phePV30goFsb
Yr/GrzSg0L4wK1dE9f9iq6xDg1Qx/NsB/VnYwEfVQAnPqb33e+0iR0tIcJ+8F0L9
2IeUZa+Zvv1Qpk50cEIdZ9KBAIpTzesomkjlflOtT0uBaNGZUinPL2OnWeP89eY6
BurTDuWxAkq7luZwZmXomJXveUm0TbtI9zA+dyAnkud/Rx7J6R0divpK4uIh2X1t
TY7ArTqP5JX+owKzn6JExT1LqfioxZLLrcmqWLL8bTLs1VYZjjc3NxkCDnukHPnb
uR7zK4+ysg+kdtvTRcKKyHUmZqlLgb1hA23v090OaO4IZIWpU5vvNFEO7+QKo/gV
Xgu03NMfxk0pJPV4i133IBnoTJGY7hq5ym7DjbbvRL9h8DFicdRVo/nypTZsoEMl
GsB334VuKSeKNmRbxY6+jYegDxbrtdwDy1IyNce5N9XFfMitzYLBn861GIChSApP
UqJvUb4Bc6y0jZNj3EskKfbV35ZvD7sl4nx5o/8mTrtFXfKKlNQ2EqxE3qx6pGeX
cP+bPorRadMur4d95t3f9kEGgg/qk5hrNo1V1kBq8jtYM3DOr0nmLNxT/gyRUGxV
K7evLtLF3Vkgnf03rRA493Tx7gCKOto/CwrFceW0n72xONftzoIWRwNUp0ei7DpR
Te2+2EWFkHrZIfFbojq8JPiaFqYhDceaZW0Z1ylqu1KELWZDxnH4J0yGfzRqlMvR
VdKW6FCnp51QoSiBcZm9/8YfHvUTJyG1hEP581gYgisL2CJboGLpnlCK3vR/5h8x
u6PcGUgHTZ/jc43UEKSijo64szqpka11ypTkEB/zNEeJwcL781cvfydu2pabSOw9
DZ1CcEKi+rF8O0RcAmh4vDUGZtqzNufqEwy9/RT1N0h9nT9RfG6ZW+kxzTKGS2eD
dEx85AH/HZoYkWnxKULsXf/Dc3AWUNf1t+uuNq4V3b0goy31ghwfA+1LnfnV7Li+
mG2H2/o17d6AbC1imhrD93FsZ+HRTDFYYJtmL1jmJQyiY+eEOR6aaRXH8yb5O6k3
H/TIazXOD3mri3k/BXLgBIY/oohEp9rPnPX/UEE74OW+omTFztao8CdG/jB0nJP2
lR3eOPSg/i7CO9bjGuAAJmbYMgE7d7ouahtYvF/GXevzjxYstCGIc3ZUSxVIV4WX
H3lJyMxTF5XJXFZHOf2T17FSvmPwVKVwLb0KXN9NWT1bFqnjFBFZKPrj0hH+TfHt
DrVGetoPIgqM/IZ6vH2l7tXZZw2vLi0Ck4bc/w+RIdJC7/f1hZe2+Xd1bNVGggbu
OVTdHCmnwxCYe/5VSWThIDHEHByu9GcRlMtiJ4aaXc6UBsBAemjmSCyNvS61EhRG
5XaTEuRSoMm7i9cG8LPIi1eHE7DQjNYoDsrSWnXzBV7Pw/OOIxLQQ5oi+nRzU9KU
neRjeOns8VHO42EOqIqfGNFFIVHZK8wtLbQtT40WvEEmNBK7Z5R4gyq0V0RjbHoR
KiB7zkzhEysw8xxA2oq3DOaGSobKadpa+AIQsmkujVLcHP0mMh0q0hfxylFNP+P7
Dp0mBAg8UDYRexLNo0T0DHWXVXKw+p2/nPquuQxjAriF9JYurV9v7dSw6+IvRkSO
pG1zJRG6w5WbiT1YxfBF73HVTD1jpjLFAxvKU7qSU8BzZfqFUGLnIo0u62e7K5El
lNt8ykaAamynl0IhvbevYtNwu9aeNQRMFItRdwC+6OVcM9+l5tRCdC3dDP/v2UtJ
2BNZ4D5usJkKKW32TofnVIQ7EI9PIheYMgQtNVWlVpECJxe3ta4QsNPAkRYmACc+
bj7yOAu7eXzNHt0qfZBS3ulqIWq/cVur4wATZDc5HYaNG82uxj2w5nDQjXyNLyCd
gWvb8APPjSrP24aQHaujzNTCB6BCaBRkurZUBOBKG5aRDiSddn7NJIDIZyJUXiO4
FCBMj6BFVqUlQ3XMtHrx3rg4ZLMjZWxMuJJ42lKgGIeqr56VVwbA+xYOM9+JH7kJ
FWQmDC9dBE2Derrbpdo21mvi4IoSS0IC4uBKwVz6SVh0R4oXIIgX169asjr0lEc4
pdA/n5v+pDsWFIUBu5TQIS/40EDe8kcj3nL0iRrQIZmzQCD4GzUfVhktemRcf571
lBRKPBZZpFQrwZOxdCFX1EPN8yPoHAGqhIV4ksP6JYyUuvpBAYvAa4PfqTtcenYo
T6/UCX7R+V2yW+0RoiNw0TpqVeQl5kREJTMTrVipZlV4m/0zvrJqN3GfCut87Ksy
4kr42I/pFN/zp7XAHJaNln62NDdQEBPSfnBafC/IlFG036QNPjcHNGa3sR5DhaxF
9xvn5w5uAVioaa66ncHYFPfhAhysp3an6GQOhWPps1M++UmI9oeatDLeQyC3Lo4w
nJ/xVu6DuykzxvPUIKhtqpbmkI2biPagY4p4nuU9Sj/BijiyxfG6gEkwjTrTNgqH
A3/T/hYdRIilL6uytgbw6VJ+eYskB0qwBhtCXq6DHiT1CXGl12gV66aXSHRRscXu
IVmCyWNnbXFLWTaypgRVVJA4923yVKzphOmu/E7QIQtp3GCGsDn6tCvWDFGbTkRC
5UFoQ1RCdqHaQHc9pRrwpjRui/obolS/ZfShYSbDlCr8UG2K5pfZDxoic9MDnu0l
jQiBZ7evAT5H59LhIQMsMNN8tr3WVgLyqoX1DUQG7Em7oMrNVLkbrDWAdYc8MWJd
BYESeOo2RzjpODdzVV/u+szAn4aG9SSLgI0dPSJCJ3CuPSxpm8TLy7y277lMPtUn
PRH6P3m9BCTV17f+lzStTRSbJtL9kehNagoDGjqpGpR76xjKd8HGCtUJ7Tf9eV20
gDuZxfiZXQhS5M5LutQhXD3DqzD78lSqC9q5hq3+mCucmhr7z6QGeqsFLs8e/HmD
cL91KFEekHCsaZ54B47wQjRnrtPx1jtAyDi7AMBhfEldaZrpjtm2XdPHLwyXyRlj
aRs8VOxYjO1Eq+zs4kAjPxJOkpnbWyk5c1p4pl/PHcRQRfhnRZCIsw2jxy4FF8xj
UhFCGVGE0RutlveHYfxVtxs2uGY0TTmW7nYXhk0v30G6L52eoY9/8wKozshJGe8c
Qfv7TpiBcnUnTckdWKr9K4ASj3DgF+72ZwVF44FFVLtwH9PZqZWkroU5czAhn4ZT
v/Xbg1is2ip+6G98quC9jwp/EIEWwchcwrs9BwaktI3SsZDzS7bvr/wka7IWPDBC
e19stziyNU+0y8AJ9MeR75q5e6+tzcqoNrHCHDviQrXo1HUeDDg95DBtmKQ4g3ke
Hng8en6JqJaTDi24Cf5jkchs7h6qZgAvEQq7iFRdXjf+B2OCbzoQJKTEAA3dKzJW
4Pdtk01IWh8IhtrUDeNPkMeJ4gtpgIHaSHRAV6n3ASuwsJWHDkfahT8Vz6gvghBY
bRBUNJjuIiTS+XOOz+hOYOX4j61vkZfllw0oPqenFJqFBsMIvmmIiQWvHKwuB6Vi
zXVyMvQjOz9QcqRICYBzFoWAY53FbUhGdNlt6rUtbXHs/Ggyywe5umlbDFq/dEnm
+GtDosgjJUQUrCXA3I2ZoOOUQZN3AXlb9LVtIOrTzirkMCgsi6d84zF/j5+8p3kg
djD/P86tqA1qXmoZiICdLHk+0VS9GqZcWcqwZ7logN0w3VcTyc+Ofht2npBMPSXP
xO2e2q8o6nKfzHCnI8sfieC70/15xlQtYhe8PWwFbctGHnls+i6UXqnTNrBbzImR
yG29Nhex9TJR5HxHvH8Kn49HEsiCSOqC8wysk4XTVdHD5IE9SI7xa0vxyiKW5GVL
r4xpSNmGLhyImwOLDf3OBZJqDUB6d7L6rFAzHUnwtdRpt6AtlVQ1chINlVP6J4YA
HYVnfhOTkDvSW78rZvLVi3jMbmQqIASBtia7Glpk5qdqwGmg4Mamp/oweV38DKyH
CZoHd5ukcetTllkBFD3dknbArORN/zjeIv8jppGBbXQA5mkPWCLW+8Ft06W3oj1z
hiFOORpYr2E/vkWtqHH6puvjY0IB22yPMc/TPZmRjv4vyi3NN8PHIQ72prdc4ShA
EzefyQ3TMO9M/D4ETuafzfxJQr5JsL1VzlMuN7lmmGi7arjugkZsFH0fMxCFS9eH
/Pi77R9yj8DHfTQiIEDcfpCxt0+hEXSsm1bWhxo0iWmmbT9T+x3x10MbACGOMIFE
M6h0lTgEKzIrsPG3eglhhr5jz9laWNVLztRrpAiW5ArtqquTsMxWOgSQmqakobFr
Vx1s/oCaAqHs7KGzxGFqKBICmhomd1ksCv2P+XqVFIlTmSW7leb0VNEZApMN0YEW
EbGAd5kOUqROGMocCfuQ++sY6s82jUIShhiostgN6hhpT1ZhrThLcKcZOSSX70Bg
0rzodj+a9bveJ+BEK30nnS+TZxwP19B2xNt+cSWJJfDxh+oXT4wHP9A2AMXDBjLL
dGA1Prj6pme6H6x9o1Lp+2F+JLkTvJF+idd9+uUeu4V8LJ9YuIqzWAwbpf1Tdi8h
KBauKFWd/0oG/ptzGLQOyv2Q7otxLi6CMhLWtiAUIemubcevAP7iGmlVgh2nHmjy
eAKKPuQHJHj/WMoYgobD6Q/9NWLOUF0i2uKWIdbWQlCw+8GWzf1Serf+/d3dD7xX
0ti+fVKxa23zgK9jWoUHK9tNPkHjfTmJqaCX1JG7HB7yWtkeqy3SdfXwiVp+oISk
KofHhm3AdjLmsmPa5XKlBns1896ANXL7j5766ALlwf8C8xjpEcw8bzhFjGaO/2TR
r7F4uPRwQj7ZcePTGZ2zdjaDU82xtFoR8s8iZzybRiy+TvsPtTO/lFwKpoB8nvw8
5YnH0yEQoH7EfCB3Pyq4xI/kpakTc8ramscqYxjQ+Kbtq1ZHZVkb8dYamKuJkOte
724rj7fwAtKXvp5fs/tV+LnoXE0ly14wt3Wp32kZ5EaOIp46HcmRYxLLd4KUQNpG
u/g7EKPtQbpYBoDQt6KM3+E3++WSsOuU7rWvdRcsJkl/ztm7rfHFSYkfgzfD+iLg
W4TCAuEbV/6TUHLVmL8/T+uKs98sDdjsfvMMcUh7RSKCvKXF2L7S/rXURmNRX7nR
snLTg30Fz/ur1rERUkDsY9nxbsjttG23R56OnZ8MnE6oZ6qMP5O66dvEWxa/L1F1
N50shUesaNu94ent8DoeKe/p4L9z0VN5ii29hNHmBiRGjVYLCdMr7mEBxxhxpP8o
NJ49ZWh4eft/NGIfdXM35le/ijgVRBSKAS3Nkb22UU7YkAwlmjKZis9dgIr74uW2
icCPGtgBw0COT7AkpZKBPWnfQFpR99wE18cUbcNE1+umsGlEP0SOkx4peqzVZW3F
LPl2f928whX1m94IR/nGzgULE3J1/rwaWf0xykP33bsfOGhPKBrEL0WOqUmK3bYU
NKig9e9YkiNe4knKtWKogmZNrFVc81b9uKf60t1i7E590NxJtpQfJ6+uZKrmfDRa
wSiZao2M+ao6oxHGH+aSnFrpTOMuPBdJHeH0Ywa78OGgPJbevL4J6rplkBgZC65k
BHdjO/dE5bvG5nwpZl64O6iG7+JsyXlhw8jCBOgn3uXBkzSQ2QaMxf0uqv5VAISZ
Gq5M/kPPug1Bym9INKZrjTrEzcg8N0coOTn70HpwSe9iPJ7u9AJzHBm6A1mZA/Zq
+85/RzWB/yVhsoHejmN0lf9VytCvdn4L2GVZ2JlK2oiP+cRDIhQZD8xYTHy5SlCg
ph9lHlOrq8G9ZP1jKkKlMcG8Gx5FRm8oPt5jiVvKAQ44cMjcAI3LYoRhMCOZEpiQ
gtAtA7oqZsXHRivKIgXAnIiRRe4rj0WlhdQsM+KWlsQ4FHu8i8iOJodVEXGCHa70
CVJItesxaznToIc8wcZwblaStNPXD4HCFsk5QYFcMRdN2jVfZamw45wwyH4006tM
4sZAt2fUReU0i9ZVssZPMcxeEM/vhM1eOp4vt4OFraln1ir9DlPAByElXwoYRaUb
0mqOFRoSoopv1aNFW15r8nb+J9sJ3zyTrvYk/GjtucXNXHUggLmZkjbKrneQ0wRG
GqWMAEQfjlSUWL2qcblDZ0Oy3l3w4M2XCo/yl1dh4yPkWdXHX8oGRbWCdZcw6Gec
O5j1qjnqoonfpgsukxp2ZLyc22vo2H2ijAtekXGgV9JBi43OS/mGE17n0ijjbQL1
PnwdD4PIi5nXWqVSqHf1OwJV0SGUNiwmUH1wgkH+vwijK3Sw8pDOujQOLnrwn9WN
D/ijEUHLSjAeQbQvUI6OhngKmhUfA8UAn8RpCJ0zqIjD8cYznJ9Aw6Kvh6ZUnAwR
k0JeV5GRIAPUC9GEnFM+/Q/JD9l9HO+9JrbS8GaIxWT7X3+olAnZPXM1qClY4sp8
K/yKDKfE/BnElTex1AcueEv6UtwF+8Gdatqjnv3EzWAH/ijQJCFa/PDNxT9zXdKE
G9xRbPMKJMlLUk3L30aCL1eMUdVdxC5RhN3Md1kaas3wcG1rEk/eXKgnSoNu8l6z
H5haFqCdAQvXdBzz5xsKCibODy1BwpYV29yDRk0e/jFLoMcoBkW5eNL+1vNfxwzC
mrMMxAR9hFSW2jhD0qJButvmGbbBZm7bOY87xVHR1CyS+ifRLajeQP0N63sSNM/D
GvJugroxaTCJ62lUyHAebZh0AmpoX2pnavbdICU04ssJRgZQFX9nRQ2ZZcY4XpSG
HSOFCN3nQzlmWNUCun+g4m2Ia50KqKeEz8RYkpyh4OPc08GdNC61W8MRQnv/gg0y
edS3dsirzEHP7kVJu+2IKU8BMQF7yHHUy6Uws4FrWnYjgkxk+oSYn31edQoIoTRR
HtjqTji18NH4HSC1+qIXvNW2aHL8BO/0LMYatRb3NhDhiesYNjGM8um6oXdC0J6l
fTaSa989ZFpH3gBRXWw/+J0w0xlccjBuuAaZWgOPnncuGhOEKWBF8MjbL3b42Z5T
RqYx9WvCU9Sx5Tx2v9/7eS7wOUZMwaLlPx656X0ZA+QoYWynnKmCDiRZTC/yOR8L
P0uu6TKAwQlX7l96umaCDkCpPxAzkf7AQfq0EZ7ydlYQ+fjFTpcMZJHIePGtTpQH
Y16Oom+6fTuFp2BKO3lzX/W8PUf6Bo8pejs6krOtXD08eqwIRRuo9DjbCp9GkfbC
4wtuqXu/G8DzqYv+S8HSooc+oUWmAH/2j+syJTYHz/3XbefMCUExHD/PWsyGztk4
MPRFwtiPB8Nrzz1oo+9mvEncVRcNZxaYDcaNCTWiWvny1ctTmwqCxbWwMA+MQ3yE
bcNVAFL4/ZC34a+YYzH3GnCtZshUMM7RMgs6BtIQXxSIHgKa2qiQKy9g+e925NHB
dI/Di8ffeUurU5pJwZm1UczwFK5zdVOqhXFVa4iv/KMcLg79SdUjDEghi7EqXeVp
JMtnaeqrCge/eZNemRZv2eIN7UmhyEkwvnoF1tfU1/M+eMZfdg1WXY/fNlWq1gZE
3v6bXHLkUh6SnFRX7qaO1YBSip6urqdCC3gusG2haN15KrkJYFRiQO8DT7YFmKbI
sviLmvkF6AofQa61LIFT+WqRemMxxjM3Tvo22DQKCULeUuifpL6d0PIeeDZ4lckV
Ob2tNOlZ0LN3UzyEqhh9mH3nFXXFnhVyKs7uLP4+k/cUxb+pN8IiavjdfYnKIG7U
nO9MEDgXNcf8ldSFUBRKykoIwDHOeQuWZ6Zey4RcHDB7O3LinOAnB2Vv3md1IpnQ
tLL6zn8FfQLRx3biTtHYeDKOBnsNtJfyjPXTOploPpOHBk0RM8uTP2MbeRf7WFbf
120Bn3E60ixkc+kaySabHSVnQ+9urjsewuHCX8H3ndHrTs4feJRQ1AuSXOME9ZGa
OQgGbmgvmrbCzHKWgJWcKH+fggVUQrxEv/8H9HEtEO9Hai/TsCoKj8jSle6dyRis
IS14uyN75wGnxVntBH2en60AZljZ0FScOtBt+qe+sL9ctHRcxWqd6O4B4EKeZJbL
SoFRDJ4BCD/S1buJLH/iy7uDlZ7aPgyEunClgiGrqOfslt3tgiLzLeqD1+R5D6Yo
uY7vMjTVRyXpTLUQTYO3B/JbGjAZ/rYWRiffCuSYMt9h3L7AtBRFzRh9ypAaB8aH
g5jPdkeQg/mPB+g+c9jARbSnKEmEXahe9vDAJ7IIpEaY6xYyczjsIdS/NwyV7Vg+
asBzXWK7GxBNNDAkIrB5x7SJYogdU4S42uVL52HhfzuUaAdbBlU2oQk1nWAI0o4B
gGNzk4dG2i77elSYqTu55kj/IMeXuQVPv3KwKGfIsLuNpN5Hb2Y5ZM3CiJehI6vw
Iz4/z49uz8bOokRrSR1NJHeUzekZJWejFgHG/CkTsOi/LGXa49RTYipHFO+uMjUi
r1eKmM0nTq8ywXOeNsnpMqN4Le8Hwwz3O6CQ8G3jOJx8ojPTRvEtPFKKEhAEOLUg
+8AwTWYrxzGAE08uZWnVsgmMK2a4qLi6UftnXXbS0oCLaB1wcK+YsW+1RiuhOypM
JPMqAaKyzGtAnL4xo0mJ550CHV6Wjy9rw9eAYalqrzUZK1sl3zymUaI93JOToch3
vJ26v+TX/WjWAQs9WDe+tGejX79uQqRGaVDIww+A5a2SCEX9c990aBKhpGXwoUa1
/5QvDB4V4zreqmnWbuMUbl6VIdj9d2TwsZimuGZaGprLdjvCp+iU7K7ZbcKrQbYJ
SSuEniLAbhsVzx97cPkY3tM3SHqctI69jN/BO7GzgXLxwM4+i6LhSQGDrPJ6Acxh
vf34hDqfGrD2EehU3RHFKVrS9Yme2ufWRgiZJu9L4Y9o04OktCW7HtzLr1hgZwci
NXnLkexFQWk7w7jftL577LxPb7/MQngwffa+wZEMjZJEx0JBiMXqUbsqC4Q0wKn8
4QOvKwNdj0taTXv/r8ujH+M/NUruVQAdIogQW/y1AW29KzRI7entkt3AzixqPpjY
7E9C2EXLIHQ5+bQtfo0B8uDDKUOprpVtY8EJUX3dBMOG23SDICvrzSOw3tk4/EsQ
rDoccoqkoxgWkt7K9Owfi96NDwLKLqbLce3mgJKga/e2bmmg5GXpkT5DDyuKW4ad
0NXTn3GbCEZrm2FGJzD1yyQjCBYb6IGID94cd0M9lT22D9do5pv1it3MjPn2XOGU
xtGax+8O3gTO2plfjhgGAPshaR4JcmOtnd1KfTpAt9vqmm4MTDgKkDnBOhsa9E85
BT2LsuFCbgJimhCNxAfdnLHaf9GNHThZtCjNchApxpxZz2ERZ+u+x/8nANchwwIT
oLfm/lySaYtmIe7d7ZtBPtYOHiiuY80Djb/nGDnaQYwSTE9bT5+GhCs9zk7oqkxD
t39Dl9fe8Ap84fRjTcj3wb/tH2BVqfkJxYCVY/P5AkVpeonVzwq3RDIFiaeI+ZeZ
tOCZnry/5VZLfwpEvMLYVlaECMHwkvCElhp3BZsMzkf8qUTBcwCg+2UIxDAqQWj3
v5QaOGnsON1S1v14Z4KwwpkZU5hrFBFWYtlP5rLVkQsvsg1aBfYsNrYRwOf3Rcsd
U0/C9ip5nU185KRgvYFLZ4u7HziRq+o12eXvH5Uv4AlcSjBRE9DKVBlgxOCEIq44
3Eu/cfzvjmpswwakMB8uGNFfDxySJkxNodD4gp6n6jUSCOS2C3RSf/0cS5sIcsIp
UlkKA86SgpukmDIgqQhrL9H8sAcwLoK+XE2Iz15S8IZKYBnAIhkn6ieGRK+Vlb/N
LLTrIyWuogXO3iHSsZnv4zOgydoAoWDRnrbaE5swCny7rSNTKM1ScC/ilBiIhTlh
cnIgoF2T4rcoZX9pXKFi73rjndKPt2rcBgVtSUYMl0HszhF7nsiV7mhxD8fonxb3
o8LP1WTRKLGHZ1+4N+5rLQQmrWbr+eHd9zu6HclMpyuw8uH7H+guem3LqKrs9nOT
LENbLtMC+hT4OPjjRpl8FHjxhKcuaGAfU8b9zJf6xQ10fl90LGYcFQSZ2ixzIWMy
k8rzaGs67qntIX7/5Ecn5VZkpXHZf52J/oPAkFyhG5yqKOQwFiWfon6NtdgYzMGw
VcY+C5rVgeZcfgLmAUdFRwBCSdwCgCtgzGdFm+9OSl9Gbh0qV1/ORGJ5/pdMPqmT
1X/tgOjzPceW4hijne9oUKGrP0Q/kesxwF3Fmm98CeIj15AtSHRPhpZYHYXvjKRz
1XSFJ4l8PAGJMFBEDjh29PUnXbS7DZ5XKs5y97Nk3kNU2EypY96+/p2ZtPZQr0IV
5lBSRVekBLGethseeAngsHHxbOO7O2F2VkPyDzDLvyyeeHaDU1tRW/GBcFoY/Xxp
wL4hm628uNJjodklAbqpd+SOIk/QqbQYW+ymQadQHrVYcdvgU8N35yvH2i8ImpkG
YzeOOrzaMtK+6VuKANxYEWedfMKUtFgOnv8adPsxJcCEbrm8ZUOy8B21X2p9QUC4
X1B9G9+g0kcacGuySzZ7vU1j7aGlsgpUVtjLyUhE08Ia97H0+JdQ5zQ3nTIUQkRF
ruxPFkvFacDY3MXXGfgIpZds9u7eX5NmlozdpMikd2zXD69ck9sZcRw2uQuuEf2u
ajBKMASmUpveqI6GCEvHUhg1podOkKn7zK9Y4CToWO1u39s1B9/CTXARYLf1PpK2
aV++nIO5LE5/I86d+176daX5Lmr+SNithojGlTzg0yXChFRekjSobuyS4PNEJaI7
wgQ+mUFux5tPdvCK+Go0ubQw86SY/gonzgriNbHDl5v7iLAZ36UXi8bwNBdvmtad
XBym81einVE+KnqXDkgSifq6s+0nJ760IjFsWFWN3yTa58aeEjzlJrjx1eGO2DZX
GkXCXvKB+5Livn0TbqJNTY3A8X9nqxPAxEK9qmR5k6xfTKYHvZoLksRPUpIINfQH
2jG3pK/9cphTVpic90+d/8ZE89pOVoKihTeoqApYmDte51xpTuaeOEC39Ddai8sO
TM+HWPGDHBD3AyYAMdMSMZcl2j4gdH6ectFLCTQxBYZ3avRT+EIucFskXlgrELIx
JI2x1BEFgAmx7IRlao2KCnk+4cEx3eTQuHWQo3tdLWn9UDI6mq81XUKmx5n0c8bM
jnnTqCbL1PdDu85xqPCmbg/hnQEAu7MsLDmY8jIfQi8Fgmlxs5tqeEBgF7zgxVrb
h50kWFkcFrSyUA0wmSUgU9P0hJSgktQn9ZL1qrDpttc72XaULhBgKoX30DvaMmLK
b46JjpBSfqO/ceqQjop+A7KZ+gERKy7gs7W5i77ZGaVxBgDyUPjvID95dtRqPmN3
f0LIT4PtmkwJ56rDOJcIyzi6tudHzvx5G9Blk3WBr/vtnjvvAg1nDZQeKZuQ38DZ
q9f1/hEPnIMeUMJHtHFUaNpgx9ieH6DteAeO4gqlo/IsEaXnds+8DCPma4tVmkvo
JhU5sT0AqFPi6knu9QvWXJRUmo2J1YsEmmZH0vtWHQwkHO+xYV8LpYlEBZIfIsYl
wa1j7OsberBgj3E6xysCjQo8/VwfIPCsVXwFvqt74WIWcTvaImtuZ1arfPPdGKmc
+mfT3G4UfsKM0mcZX0Rpd1/Sh64pwCJ5ih3yb6gRaqVmJVeP+q6CgFKXTFwLlDYp
JbZfzbtS/O6B+8UcrXYjhjnO8wuGNP+bUo3+5YsTkAEftc8X7zJXUGuVyn0fP69D
nZHZOeUeDtApCqSzmllZ8yYWKLn2RH+bVxvDAmahEXt1QODQQO7Hts8uAKdxCcX4
I5lDvQmLG1GTvqTcSNeEfGF2pc/vSSSOCW2IfJjpuFHJTNS36YZ0lN2L6feIcdD/
odyEa0w64z1jPGyz9SCM/oTWq04s6cQItkr1ADC35n9AplH2p6PhBLNAXuaHGAM0
yhHV/LEIs8sQ2jbjWe0C3SLt4h6mwg0mpXapEsaLyrFtIgbJFkpH0FEhWtmqFSzt
wBFzPePfh/VeMqZrj9SKI9/y0VCitF1qqe4zQYHM1XcNRwNhHhKNLTNW9K2HSYEa
vwNr/VetTpqfe2OMKSUT/xCBikso+a0q44flgX2S0aOyrSQaNv+y9Eu4Fr6H19Kh
d3i4FSSt0X1BpUnqCyfPdUH9EYzNtNF4z8faaSlOMAsrKAaU6Cn197Is/I2vnkUH
iqQmexebDgjLGS1gXDH4JcCHUcZnqEN4dYPekVRoKXTCPwcdAbAmTCRP6ipx93LM
IYRhHK/XhM261CTIyxDM7AsqMUvlkZBvOc6oGieaI52eZ8l5+ncukO0FT16iGM7/
SwhWjjtu6/p9XOY3lgtEWdF+QnnqkPrCaukae4UXpXgbVWu8E3XBrE4UsuiMs+tv
q+b3pkPkvIVtyhaZdjoiLIupQF9M0o+QC7xWmogs8aPB3u5QDFd14TSMC1akBKNw
UsGaKMBFqKugnhW36xwZFkw++anL9CvY0ctdYKpXqt0eu4Gm40LkNtt5RaTtc2yr
VVb+41OpgJGEp7h0JkBm7SlwTU3d14TQpy/i6jOl1uOjJFHMmme6P5MqYvoggZSP
4z7gHMqco1o/5FVFfSeJw7KQ3LqdnBz+MLvu4OjqLjNfYlDP7g1pteiVrRV/StlQ
UkJ2VE9ZqQJEteFvgXnVszwWNueYzKr2FBYddi1urKU/6RhixYnsPmpviMW/g4s9
qhYo5CvEisuSdCNlG7OdoqWsSbMddW38oD8NuEP9omrjA7V/KIuljKsSq36ELMnx
KW/wX5QT7ktYIgNHKCekrigBEWFaPAcfbR9r0Z0Kf6iwt8QPKkLjMYOkVlSVmwR+
k7Gb4jUdgCB/EkGA2vFKQdpY7sdCg6xu6Huokm+mCPedDjCVP4CZdUkzMDPMdAVB
84rz8W0ESXqEfOr+V5sdtEIermbrwaoK2116EzhpNIFtsMLKjV8cUtifLLuEL/GY
5p2g6WFfS7QyknAOANA6MH3mVeC5936SiDpojmOXf5hrj4zEI+RF1L6t4lhQF2Dd
v60miK8pcEPgdOZiXAmlZXzWGLQ370oPHV7pk8jL/hwq1zRgZ9DLGG/YaO7nLlnT
VjBcYE8X7KNsJ0JiOyKd5doIDE399vM9HqmKKWwDAKChW08ZZwy5HSJ7bQEjRqqC
esx4/eG7bbttCcWJoIVokV8ZbkdQFCDdESgqvChzcPbI0Rg5FtVoYiO6TxWOFU/I
3xZgi2ThBHj6DDY4A//uXjv7Dn4KrjzraTEjF/2599WIbIMGctoA7I/LMHI8JRQr
62pTICf1V/gE4LKnSv5MWNeFD5zMkxN5WH4pO7vd2duot/IaexkDoJcvCQ2Nz9OL
C+rvNWNwibBFGA+aZqOpMqs1PY7oOw6iqoPLARtdTdvlBv0R3PQcsNYuaAvJaY2O
wVm5nppaDdrN/oxHTey4HiYlNbgvAvLbZyLZzXpPpRKqY0/G+oiXldh4fugjlRol
nfkNuNSLAXNmzTnj2YagIauNkRJ+PekbTMz9hGQVS+4WLf2AAAwhSfudgo99FX8A
qUZdUTc/sIEIzWtHjq65vj+b6tAK7MraXhgcG5iDTkVBp/5dyORNLVzJXW5yTIuK
tniiU6aihdYJX97bDb3ueeHGc7lcLQEkC/9LqQ+oQC0aiH6l6hPIegDqLSfboBcO
5LR+FySpi3l4LyIKcV4H/fvea58BThXsdZ5f3NJ/dIHRzHkFh6k+U9xEszRJJMhI
hMcv6g1ZQs2eKDRLTsjjn4MMtLbczzz/JznLPgk0bkaib+SLAEna+l6gor/ABxe9
vFSuRT+P8gFqIcxhmL6qWdSGSSJDEJa0EeI9poULi7nHUIKOsRkD9a+QH/FFuNDT
dT2+gdAcO6oj9e9I8khKfpp8ooPjz9bzp0ONQV9mAuhWANlj2doN/wEENqWXUR4y
6EgyecIJ8YQm/Uiw/goAhUUCAMEUCuvO8qmdSbLB1WDebdQNN0OGxGxNrHUHZzc1
95kO6Ys6Tz92jqeg08rwR+wOMru34TRkgZkeyhv/7kyW4/nb6vSuVivqDyV7zbza
6UMPvIb6kLAAF0ydVMOPJZI2solixnCz3qgjLt33GTPFSqvZf+6KvT3QBhnd6X8C
vTtw3JeydtKIeXBfofuUakEpNxUWPNe6UGLEYUqUyCNWym0guy3jx44nQOSmndwT
ezUdzbl+8bdK8ALyd+xlRAnvbaaOvtnIlCdvoGAkcR0EQD8lOdiW8kFXB5cbZ9j9
/ys2HrCvyDcmcZ62fQ24/c0+vO0Gdi6U+GnzKXLWQEq+ZG79BiVnIYJV3J5oK6Gs
jf72TPjQdKP4C0TBTJYhWCRJokkizvzT4tYBegtdXAcraKiP4n6fPkoSjt9bdGP+
wVg0FWFPizH5wkrKVBLApCUpOj93PZPIKiLhWpJEC/NgcHPYmGWNfnNqYWWfY3n2
pgfQHHoZ34QLEXp0uXK2/s7aYkCmCOQZdvRcTWYhpdwaGI913tPCZ1DD0L8QLCtC
mltbnVb6Z/w4jvXwJKfiMj2ZWITw6qf+hKs9K+U8wh3pyjFVHNkx5nR9UBxjHYBj
HV1rvyS24/FZgTWXumKOmqRYXhjTR67TWqa3U2f4Y6kYcd5/R0CZGNdyWbqfWF2x
cxdwZvpEujjRPDnEXbpdbi5ttTpGJpNLfMA9PzdnjIB5Xuddm5JOo5NDZrDk9pzX
eo0w0DqsbzuzwER/u5zG+li47wJv0SUx4InVuGdyJ0irVcWHbQQdMAkjthHMVYdp
T2L6BvWXCJDaOXV3OuR9GhcGm2FZUolPc/Pvlgz31C3n1ft1HeGvDMASk2W0G47Q
r6MKA92kOn8PdTMJt1l2QU0sWsy0JEkh/LTsTPQL4ajQ1wURANNqvHw79bzE53i/
0UXywFRbR+H0YDVaptgENtVR3pKuvr25TXeBRHI+0EzZbhV45JwHJn1YAFdwNpTm
X/1iYNeVdWhyF5/v/CbzYZ8/Bjjs4+yzdRijEieF+/altSY+LQyiXp7osCoj9L1z
zN7bHoLzZQOJ3Xjmi3c7luoAMFK11Xq45xHPKXl5Oa33Pgd6QKxYQgH8PyH5ahqv
QG7f7yjZo3Q8PX10IoeqLsizD3jwdOtznbv0GQq7jZq52UhbndAdt8XBG5A3Htnc
CL2sm4HVmSXKHnyU4tkduy/9eiUNZJ5Xr+wcmmBHc0+nOKoIzD1b4DhPPq0zkdpH
ps1yx9/31/D0DyQfr55IIfITYTldGLGJD52P9gEYjKIV3xJKwAObmG3YHSyPi/gS
qV/kGn/Q7U79HgR4Xg4hwI/ojGzmA1gGCtyWLhR2i2lISVafShYSSOvCKYOgnV6/
TCJWuWyI4H/JoIDNCtD8zY9LMv17mPxu+HcTVSwj3xRKZKKS7YuaE37XT/5ICDbJ
+BoLV9mCSWsnbxeJlbM1E1RWG6MxeQ/NJWrjiGeTWpgnTg3EG5glVbm6ZNdL9HrG
/W4er0yXwPQqz2Yv27mUDau1Rz13y0qxwrTpthRVUPf+gwqO+HmLxwNGauqm7hLU
MdQIKo9vMHFTBwq4kweJha0pDnCwMSQhd0+iP7wIOaI+D8QN0cyboVmptU2R34U5
mWPOs5OYqgiI03z+rdBUWzE5Q59dTnsB/UwZ+jhCd52uhoQ4HhuM2LDVbQwHp3fu
GomFsw9vBB1YD8Qmtqq7cwXvBTAlYrNsPdonfZ0pP6A/IQabXmVu87tH2TU+TRei
FYyCws7RBB65Spj8jv3JXuctTMakj/Xgi4cGDNwFHHpudt5Y83P5BTi8iGYtXgJn
swyo4RPz8pyFrBUX9If8BUzITAlrI8pP4+e8XCqIPSl7OWdIfl8Qod4zYad+eKHj
hFHJi2o3b1zpyrsP9HLeMLoo15UrWkaomSi7i0M2dTAqI4W4MWGv+ux+b9nndQGn
IEahWDso7qfBKrx+ULEL6mNEllhM2R9driUxBFdjwP+gsRDgAxmBIws0JFru70Ve
WRZpFIYup5b/KH63vrCFuR7Q2Yb/lj+x1XUmS+SqmI6g6FDEs8+W9vQdFaUZkyMv
fwaIYHivPY8XbWreYw5IHOMwfcd+eYO000PPiSfnRP267Ex0woOncRML9a6tMtcu
KPs0nKWfSzm8s3tH5VgY9t0OZTM3Dpu7/3CFBOa9rw6bHRJ5kr3JXGwOTzg245nX
1b1+lxMIdh5LiOwl18rFWifJeztFUiBSHp98nHtOkwR2+QR9Npkjz3TVOQkdIFxg
9UUB66zOQWzAy9UaSEOXBlKqjDA2ePVzWaabO7Pkc/FWTOlcVqKsm7GeA5EFdfmB
SZpef9Z5cAvnkD/Yne2Kc68OUxdoGZIJ6IxqEXU2ClsBribBpqItaCsDYnVdCTDr
Uu3RZbkadWnDOQprSciX6KkDmJ0Ly9N8Rh97hChrVpDbtEgcMNsnBAZgt8Y/wZCt
eAz8VGQRZbbvQO8t2uCAU9InYOOT8NYSOjlOiMLbDmPxRyVKxS5w21SGmE9F3VhG
7DlVDA/omXbAWn+JK4mfVSWKIGJ7QSFH3Hw+srXI6FTKkUKmaz61ENJ7n9bQDXhn
t8nemEtJAgIB65mcEZfBOoQ992Azkhxms2bTTpPsv6diu6mrglWy/SLK6D+ivZIr
7Q7DiPOug149r38A8BrWy41a6rLBCYDtoESPUSZC3NInDxPTz+wDmgqTDjw89RYM
iG4znK4trC+Ch0kLDg/L+IG2rbCaV/gFej+HHkFsjhaxp7L52mSVv7oWi2gYIvLL
GYojjjeyltF05mLXcoRHdFAAN0Ka6rMMacHd5a5yjijuDLV5LueBkjrSaj/HxA83
Zzpm1vrtnOpXlP1WqC7HUxrR8Vi11dobLZ7VmBUjQY4IKRUst4fQK039+7MKKq0R
xnmnoX6ZhvrJSUv5UF0N7gQevvZXuyEkFKaY/dn4+j0AxyqygrcV1wde5+Ffuwze
PxJbhnQ7RUXeQkMBJFWETGh1JSr00eM9oxTSQgXe1gsMd1Yw1OvqzuLz4R6uvrZm
bVJsAihU6rYKpNaQWNVdOYVWXCwm8XClqBUkEdMfoMPEd9HOlTP8qR36Wi2hrcML
VU7Mdt528RgadA95jlHnwDJNGSLXsUWLa7KSFgqbaXrRPRtDXFmWIvbr1wwUhq1M
sDpjOi9MH3KhBH+19tXXFyytPoeTf0SrMdlyliS+WTur6/oFc6Jv7jtyUlRAHEZu
GchQJzPlW5u1Rhf535sq8gnxV/yr1ecHdipdvNq9k3p2WWh2DBhWC4sfHxrCPccu
q+vxsEGsRC4/Sb3ykaHoWUHFRNlvgSobiBwxQL4Y8qdFloCH2rEVmBkclVTWwtQm
jVZ5/yRwJdPVXPwagIhVz51kp+de+i3C5ErhppoWGGrrOvwWvTxCYPFuD/OYX3Er
mV9U/ayMwzvcoZ+5D1PuTvKTXN/ak11pXverFfNTHR26869kix7qLjwmUp0HeYY7
lKB8K+LBRJMfmUTsNYjkdFB/XNrAGO1095GnwXrRZpeIJ6ywFvx9u+/u8SlBobWu
4DL6n4qIaEXNPlB82TToc4csPLOmf9eZKZAma8V+ydSxoG3zPWTGlFPuvxxpbQbM
LEVbwPpykFhYEkknhR8lCuJXx/pK197nTQ71ueg81Ap/d82pg8T/d2qyYk0BqX+P
9h8FL9oBx1n1vEA5X/pVbjUzCoPLF/w88RJJi8B9hoYnS3Okq6JJDVE3LMDrjWQa
i+9kFiuL55xi1mG8RKi5ixJwXqV6v42h35moT70uCpfq7vyl/4l0kqjcV4LzAL0q
QqZKvUFdMHkYMM16aCZIZYdSt2AUhYFWu/Jymk61VsTMZvre6ao9FneUOC0yogMU
aT1t1gwPSyrbfgr9dfJ8+Z2huFsgWRpslfr4JaXHCRiELPIaKeNjcrmRSF6lQxUQ
VZuAX7J/s9eyO46Ue/5WQz4lqavnExytSfuLnj83zrAMgAX0zjFx+FznncZnK4M5
ZPNfNk27ley8qTsGEmcNQPL4r5HbSwBhTPSP2KFLIiZsaZr/KlLRV25BmY8ddVcg
3bLsh6kJGZbJTqLDiTHSmRN8+UIvKzuYTEPky/atZzNne0YToTGycvlkqT9gwc4i
3xzzBPuDY1AjgEd2BN6nKspUEPiNYfMdbAmj0bF/oKDR+xlXyh8HZCGaorYtoKm+
oOVBS24s8iZ3HiE+J71+6OWDp3jjPU49er//yMsVBt5AomCU3sWtVWpDMjW4X1xd
Hc+52qA4nzIVWFcTVE67WmVmE7PoDQm3LDZIpv6oG4jfefE2rCYc/SXRLd2jyEtO
RlG5SI81z1GSLxA5QwXsGxjK2BOBLxB9p4f6EStkDmqfd7sOOh3CFsXtzPrQ1yxM
LLfyPRfbNcWtzG0YX/T+hfnR9WPdpVxPqgDmq6LMsYeIpGLDOUena1GbOEiYmQOc
1rZEycqEO24oSChLZ8FPzivEnDIzIYXbWbVAhBEpPK3YWf1hxbswZtEvNsiqTy6O
TPWI9nTqMA081JuFricOm5/oUceD+usIkWbb+ePXHhBUdUmPnf/784cZOQn/kDq7
Wjd2UsY1wVp8K5vex1Hy27DxACLY9zkoFRkucIIJmut61TLXDILX/LC+iqTEZ3Ru
cIYlYTsaJyjRDDUziOs/L2uYVpj3TdAKKBYBRp2XkYl7n8TcFSuPsy4j13hlYfhn
VOKbBYuGN43a4VQDFXIqnrTvMIqQt7WtjuHo/o4MY1fX9usYHWrk5Qbn00GDqryw
cvNNSF9g4uA4ogglICzCwdgrgnJfSiL3qpugRUDK5dvBIFJbQJS87W7gMxcGgxOg
0oGothTH3R/aZx10uynxx41RoVGc1TxvRyqkdPmFO0564CkFHixLNj8w9INPWSUQ
w1gPZl0RK1HDrW9Z9QecxhUlfIpyvI2jcfHQEMaKiUwLphTalkHDq31vZmkx9OrT
V2QnZ1kGSRutkYZsGsHrseBLRNSapjf+rITAm7zkz81YmzF1uhcnBwywTKRkVOEo
wz9QwVHu0qtJx0FU4CtDFsghPjaT7Mkig2hgxMWnKI1neC8WqHzUng82dxrK+QA6
XKTh72mVTJm322bhcyQQLXHlsOoh1jC7XWEzsYqeoIZE3hhiZKUOIKafOT31CmVM
VO7gsPaBRn1szm96lWNrNoglejzxoxyvJyyE8PwomPf0bqv0shbedcdJZCh3sY1h
VQdwFEYCb/jkEVFDO3H62L7k238IPYWNvlZfIK3SUUgHf3vNST8SDo+XXESCxk4v
6LKc/s3yhf0EoXvSdJcsEuFcr/P9R7lKp2PRkweckUT2GkrXNYA3Z5HWBWWMtl14
iI3GUAK9+Ipzk9KiaDZPkndtmE3damLYpqdyph6oDeNCIOaNMhCHepoi7ZlmcZKs
w+l+WM8XPHp93m7hcRWgRglVQ1s60hMOeOddbzaO/AMm7CgiC7SaWi4GlQMI3s9I
ieONSkF5UA1jFYSPmZUIhY0mIhZ+iR9Z83Yk6DdhTFw+aSKsupDj7dSkTFGnBlzo
6ysYzhMYitQsfqx+6Q1nqHhW87w76WvTqrddWfduVJIjJb6aJNWFrwNW6j55cVC2
UEy9zGj4CR4qcpngPf1Pjs/+M7iSbBvVSRJnWwB3yNoZ9uXnZAvyQYV179yNudt7
SmdMMo8VXWcxUB4dt4H435rVvxLX903WYuXG4i92EV1OISzH6SuBurlIRAV7FLhq
fk8qCsYtn7XWHUc47yNRSxJPgd9VOpHoB3FWW0RhY6W20RMcUwV9ksndiWQzyyYO
q8EY75cEI5atYPXAE7+2OCM17JJZY+knd5dC7rzsfFO7r+9QfZJK/SQ7RRoFyco/
QglH1NzgCRqzFr1x85/4Nx+ZJy14KNPQY2Lhj3beytEo5/3HyNH/+oMTqJBu+rUH
cBczZZBcOmZLWxBeSNPkcR4+J11+WlUmwXVBsj9kAe6iIh2ICoUycg9LvM6kPB+b
GYrAVPJDkdjDoMxWKn7JA66iGpQp/uOJWbhbFH6qvXWzVHlkBifjQNoG9/aGLf+9
nm/bmchem9mOph1uLRm43N1wybVG6RZkPzLN0BkxPO9p2qMdxVfC944OOwcmNgNL
Ga3xIzKsDsmgO7ZtYoePnNMaJ/ZxgS3sPMzEMqKiCf5ysJ8siZBZim+tBYZqFPPE
CFs2wvUReCNp4JiSeQWq+Y6QFYy3saD8a0MAwjwcFNYMSBjh9xSj5ghgBNrHacWE
rVXUI3Spf4OFC0tNkrkgRcvb1iiQYQMG7EpApuzy2H1yfBOKbLhvRssD60fFu4mE
GWJVMf6Lbj3TpTKUMuLmmsBJlsB8ojGintPeORIuSRylqNVakpXvKT+dcLoOAsNx
kPzgdIAhrdIrZeyy3aRfXN0iI+Dyx31opH4larr/3Xou//62tLatrJZOeWRAO2z8
k+TjLF5FyvqERnG992yCEqqgUpL99Nl7Eo4YHuC4s/yUq6q+Bd+xIfw+gBFMTvKk
CCHHp7vCjc7j6hH4LJpzhhpJTAF0cktGsNujl2JJrAnfmArfD06lu4v7DKObYCyT
WFtN7bxuJrT7PLTzGPDNAXW88Gyuc+3rOIMU7YBA65FqMVxCdjTxaC5Q471NeDRQ
hTuAS1gGL8yOP/PpnVKTRI6ekMAbGXrlHgFyUAfTgH/np0LeL7mV1njLxr2Zb+c6
5rw+EaNIwIVB0FA2W4UQ9E07XQn3OxAzvk7Ri42LtO5QJ7cR/bTYLtkYR+DiRm3h
oU3RhKpuYEhNwsSR0cAXRNyHuwsQeZvzKbCi7MLAKghohaSL3rLM0r54sT23Dxme
yZF/NCzUmi95CtfWryPmC23Fzi2HUlNaq1rtZY+T5XsJZ7xWGkWz5hcXLV5yhPNv
udpmX2RTpRmhweTnpMqHXVH+7RIx5Am4JcE644Qid+91X5/3R6rTNgfP9Jt89k6e
EO9sCQwb8b74H9eiyel0KuL9n17Di/evapzol7PT7qbqq/ScXc3OJ2BRtKfEgGhw
p8/Gq6sOWWgXCW808ukC1lMwkN9UJYgAgPjLKxvU0UHq96Xqy0EnjmUle5cD7tqV
LP+WkK4HpPre9E+VQzIRYlU07ggbEbWxP4cKkhChm0CZMJmjGIn7oMCC80yS0wWS
lvQiotndJuvZIyOTwAaRIhlvNHswFWznxo3e4o3R6fyBH8A0NKD82GUIHtGMsG6d
l+aqeLyLuNh81O4dVAi4GfGA/KW+ctR0DWIa5zImev4uVAqwDU7RWvN3ey/8ckBH
yeW3s5Qu9uMhhCftIKUJlrh856Rgo0ebHzNfWYLmHu2nFPDcTg+AaA9eCX382Wgl
txnnofIOvKSPEs80bhQbPLxnY8UDOpAUAxBQ8THqMXooWaeK48h/t0W4HhVDSPIZ
em7cB84ZkdO31v1kcF8P3jKPtjz4Gc6KhJPkRjr+2h5FeGzWonxsHeX66x3UfRJ9
tD8vAuXyetJGkaRjyIrhzEC4/dEd0mlCZYgdpLg8+Md2+1gkb82Znzb350Ttzbxh
C/6vXIynse4/37Hlu0eqIVHeF7WmAmBmxkhzk7191w/tPXpj0A06A8Zlc0GH0RXF
C0L6V+xjkwb3/uFdTSpmTZdRoz6rr4N6GIZWL8+zLwrian/jO6wSCCD2ve9+ix1l
Z/tiNhETBs2E3Y0AOtLeaRtN+BPIlhmXigLv8PH4vCPwKmVJcjKugIoAZ9zjtxwK
ENVlELf1eEQKn7yI3BfYXtBa6EvxNQZyTD6KP8KjYO/f6/eLdgOdIPRrZzczndtk
fVg+JU4uEHohZIUokv5rahqIRqA9aSOeK0Mx7Yh8f2RiaHil5jpBulrd8UfZRZ0U
PdQ/zXVIOImznOVpau0rgWCQr9V2O8y6Nr8JRCK3Uz/A/ys2x1Rlv2R/FSc1C4tk
LC7YePIoe8VS1P9hTzyHf+/pQbsGf0nA5NWVo7ZfZ9ORa7vSYfx6T2Lc4HY20RJt
waS8VDShTPufxrsHPN6thVjZD/PNxWLZz1CjjRiKWx/cf/SKi1H70GEUi9niRaui
5H49e2iuXImHsSmghOQ2qPjvIF7LLeL8eKlo2z2buSrYduyd7bN4OwGl54TiVVio
uu3rA9Em9RGaOQNZxgAc03n/+uJHMZyT6pZkGDsIjSPPe/6KyHbAUebhyhEJ4rWO
2HJavfQA1J3E9J78B4padQgW26amu/6OoTMFGigHU8Jx2nORHzCJAr00tgiiQNeR
ntD6104X50VCTlZ2MLaZRpdoVs9nMk1hp4RtWMtroCq42GZnyavo80c/pK8kA4Ei
BT3nw4NHG1vtJN+1iPJA5NPVkNxj/AGwP4ZsrJzsZWzj6/kQ5CwGI+f2SD4HXYvF
zhVnPs4dXX3bpJDhlFqR121M+Yk/MLFwx9DRjWfVhwmLolU15NcZ58A2ulSc4774
ZSQFJFEd11NhM+vOn+OV+9dQOukSiLP2s9Y1o0IEEMZ9fjO2BYur0dGbAjtQGO1Y
8Sfs86ysgkfkHvU6XYL/jpuISyj+9co2Gvl9hQtTXHfYveu7cPaa+VbckYNVGOfL
gBpJur70+HUNwe/5m+CEQuZNjGFrhQ5siutwkj1V0/FcMubJSXQsHd882hctbRgZ
jZfk9uRKxq2A1niOkPrbZxj2pp8+mXyOFx+6fl02JMylRCHS1PgT9UaQpioNrsia
IbFlSolZondvb2rsIV12Lt9kIw5FMNElur/KwebdCZ75SMOCPSFKHjrdBtw3z2/+
UTrXpu3eQvBu49TqgECzKYSIXugpxhzPgToECqWE4IC9BZTX9iyToNfuoHpbQ1h7
lukzp7xc9KOKhEkgLu5nMmkrQP+yer/4Dwt9+0bTnI4xE+zQMIZ8G8ouaAZFNubY
Q3cGEr9DoHC023KuEFZtVFL29c2EA7HLPM+XC+GPRHW0YG9uywYkkZ8shBuDQlFg
XDS9bItuRY5BxAVj2qjul5coR4lv8fQhZMHJgm6n+uS3WYyy79S2OuL0ZaOJpTVT
+BBNxZZh6p+vIUwC1wmqoGX9d0IK1Vo6L98OYj+r2P/0rPsh2DRVXm9mqxg5AXSm
EScosgACctfxMSVp3PkoTCxxPwLA97R+rzsx0NRxZQ6y4VwMZdsibZly3WglVMpI
zLOiuVihrJmP+wlWrrv9e671ogFa5JlCDS6/bz1lsAc3M65UYnBEX5z9HZAV9JtZ
086XIqmDRnq7bTCQJsJREah+XFd7ougV/QvdaNPkyfW3mjRJ6maA+CdXAjONnAO6
s9VXLhDGum55hPfat4WLYyM8H200uYGnadqY+pdyLY/3J/xvkQx2fVNoXOo3zV9Q
7xPmTTBMTdWl5QhP54NoAthX62O07WCOO0Cbn81UdeYWJMCPkal5j+SpVrT+CfAs
Dn1j/tHxoxODXpaly8KAk0foIWSKCOC2+KRgl6CL/KTNB/NVU3hIidzpatSFZBQR
OaTMh60eqvxgpN50Qp610XEvnyftPUOBAjdazoP0yPsjmpqRH/EMdCUUNILPFD1g
6/905y0Z8xn177bSzwFAxWzsB/F8pQhULNHP/VuWur0YNuzHk6KVkMk2v0T8YQNM
pmyMiRgO16o7f/ts2LmMQXXFyMhJ9uuWA3HaiFGfes/TmnnCnsqN9baK1BORpCAN
Ltskd+HS7kSbZrZH8X5YCNST8LuFsG7BWvcNzAQNwQtwO7pm4LgTfWRrRJiNwmW1
3GAlq4TgBgTnv9QjwGE+6a2iWuTbz3uZGKYcCaZIvXH+8R3mkBeAsy9GdYxl7qqx
TizmPhjPL5rHVdCvpCecfhvj3aRC6EBVhPNGo8PKZBHzQSOFv4iGogTW7dqlDupA
+Xmccy7jr5PwBAWS9j9bwVHvdkeDpr1TARraklNNZl21YRP/6R9kbrPhUaqywgqb
NygA4lRFKCVjWj/2aGDyloUoRDzubRPR5AEO+rZ08WjtqMVBT9A11C0t0rxTPd00
qFj7vgMJfLLIBAloraXkBJJ+4ofOucBd4VsBJio2KSa1/ztDhtpVFMMLeyL6+DiW
YaOKOLAqEk0QefaQBu7LdFnZay92x7wQKRrog2BDMgwFTZ4QAnWpPceAU4EXKrYe
EHHSyVAxGO5uz68kNzXf4VJLyy7/IibcgTLIQVHIN7fND4Xuxa2fJVT9htC7kLe3
LyqEvjCC6bJzbds1dr2Vceo4Z13LCqSt8Ms5lpEvmDjBrlFzcenwWyZjgNI9ecLa
3MJoYbEP/5K2FeGBkOX/kOZpfFn5cfW2jhV6VzDHbsoKwgTASKfjuFyl7Q0Vnklm
OORaSa6h4xv0FuXuyaYPIuCKuzsqByjBQOJK0l6alLKtIOh2oAiOHUUHrDEx8qlz
wTtyvT1sc0Ts55EM7lVRMs9PTHe2aOkhhGm1pSCCTn4tX5q/SdiPTzBB/YtHUWht
Tb5fdKlUVsb4DmKd9BpbD0YJVQcSPCggW6WnwNe8g1q54yUUwiOW/NAiXuI5X9PD
60Xpgf8MiylTwXZ2Q98D5tKQLbKm5cyPfGz5Nrq73CVo0zTAlTt084CoAYgMZxX0
C8rNQg0NRdV9aYMoJXxY79uwRhLLmJiWiVfKln0hiXkcmiQLcRy0u7ZcxtuMk97S
TeauG4sX0QcxQKDDjR8s4I4HOmhC03H8WwpjQ2HptCWqAfjuaZRlMRobWn3YiS5v
JFa4lJhCNvI7qbhBXpehfEMh57ebSQqVRSi14lZyKycx8FPeuP/xjKGgRczVGBQY
zulTiHXB8Dy6tWHFMqa9Y9u66f/E/pd+j7NDxR/w5K1ZcoNX2jdMHR0gp4LS01Dq
jgmbOizyD7fFNX1TguTq812BUe8gVBDzUHYfoIkShbEkNWcWafD8ideWEw4orhh4
G1WRVmTGwirK3htju7SzdY5V8f9x45QGGU//IjNfFlhdGYVX1/LokOYGGy8eC5hF
Ju7G0zTEfAyZ0VHm9vC5Az1vEsSNBs15A2egyvIiwh/utMe3187QQAtlU6/aEoyD
wG+qzbag+h+yv3KX5i8rjJHuhUeiQuFWGhztVJbAWfe04TqB2gNpkqOVOtSD2MYN
YAhAmXStW3R8SwNERfdEXyJdn1XFkJE3WZG/M+RRV0VfvCEKznp0wyQseb98misU
3gfmqG4bHnjeZgN/Z0BL81TWMMMVedGS26iKcvZpn4UAikQFKQ1jLBC6Ydorrk+j
F3WTFGSauQTikw4Vop6wlbTYgZN919BfdUU7f9sdIIRdmWJDc5ENobvmUQkUVGtR
deuAWLhqm/PC5k8bc+Mpv84NsPel6EEA5SVFUGDTmfjBBQCZJflR19RsRjtDJVlV
2EUscZFHoudPPcw+Qr8J6rQXrhu9tEmji0wlpugLz0MVU+3uPDuA1NOGoxCjDu0G
S3wGTWcNd9ibtPNV73qCtB88V/pTmqyGa82gxz7Uflj89ByQffImnSSqJy3VHz9S
4kr9uhkk2+UHvE2q6Ss9Bxl06QUFW8qtmVPMzt0HAslhtKEekf8tRmGd6UQYmCsd
HCqgC1Nvv8ta/qkaTNCxqSf8qwN1SkfH4+g+5dYMjkbvxuPV7ynz1OJaOT1WgoM+
xryG8kDPHmfcoPn1AGnBpdtlnVG/gU2T47CbKyaVecKP5aP2fyUwLEPW8F3Oc+eR
ikWrAqAZ+No5nRludxhoN+5jy975HhssW1KOu1M7epjG68bxkFNyjdAhxAWDHd2h
4jdds3Dy5AcpnuOUhpqFBku1oiroP+m8xNOkT1n8LW3KLqBuVM4ufMeE9DFp8333
oeBa8UQ7tswU3SC+LrxMpkRnmBqKVhWqz7slNp9OPpDMAl0WgeyLcBPEc12LXJgR
ltDhTlE90VIKMtBRpwMulkHQVqDjoksiXTSkqrDlJ1i55trAWg1YImIZrj5v414t
Dym7DZMjliHy/FDMMuHi37Zje5LrThfoRUj+VRA8J5a3V4NH78AK+k0U8I/OMcoy
KHKIKA2tbHaPSe89+dFttp0XwWZn2skHXYa048TFvsQ/lkapTLhRtZhZH4riNLt9
8uSqHGGGLWh6a7fFdohD/mqdBzIZPdrNCybQt7FxP5sNa5FJheWAEemKh3ulUkhr
7dxE/J+///aGKm8xRXbfKmutrLIW7mwl8xUaEorS/8FdLNU2JRl1nLTxqVPWTtuP
u23uZmLsrNa4kEmWmXo4Yxs7qSzxtzMMsMsxP7892zRT0iiM+uBtlfSR/M25vsxl
d27Aw6IztpwZeS3dgPAniz348i612pF5yhpa3bXGOVrwJ5gzRBdH91hut89ZLeSP
9dCL+sJ8c4HhesFIBC5A/Od8o7u34KQKxpzq1dS15H0tqzvy6y8jfOEQa61Uybmw
zSyd4tvVH2JDp2lxqlYAAwCt/FdWT6nwdyZrwgPxER+jvGhkxfiFOZNuD5JrgfDx
++CInyYYQJpOWxLEd6AMu3Mjd3FV8ZT43iBDrd+R3i75pV8tz3uumk7TsbH3eBLF
JScmymcxo9Um99w6MPhG0o8hIOezibHIGOxJjuUh4Q/VxANvaeh5X3XUQmgSrhlQ
uuCQEAJ4xRGGAmhga6KxNB9AGAqWx01f8kzk1o7gUjQfDwjhTUZhOaPVa3662hWe
Z7GhtsedM/9yoOufqtxvX3WSsf9Q3FFRdIci5mBseu3PwcdSFb0X9tA7GPgHLdCE
pLQ4hh8bb47P7/8RJR6p7VPO1TkEhOrjfFI1JZk0CBXNYm2iiKWgch8gs95Z+DaJ
y/gkx2Ggbu0gnP5z8Zujvnmuw8WJ3vtfqw94rpr2oJVJqj0Fn0Dxa7V5W0d0el87
41Axgci/L8u3it4pCMm2H0+yNJiwlZvQMyyyE1Dti+SV+QgJUV97XyDqdgfSqpwg
1UBBsBr8GOpX3arBaZqUom9csf6i6tSj5ecXSVYplbp1Y2bEtvTNfLkA+UL+cNIm
z9Dx3sJdtoiKAI5mJgde4d/nOn9fYHHSI/Br1WKbUWsJ5LOL/wjanNLXlWt7dldp
XPSyH1Wvc4s5dUmOg1XjC+cYLLbyVwiu8kkdBl4VMQakCf0KQ/JLjQjMxeuHfKrd
lJ5ojJ3+etqLxS9lBvfahdSMpIbM+uT9dv1OWGBv4utjKjP7fJNtLBAGrtdGwymp
qaUsnJeiq7rxrStlF/4dTuGNzRr9uJILgB4eNu8kKPqfZp6m3r5D/0yGkeq8nXyf
BbuoJoFgqTaQYET+1PHjjb/6EjTxXaGrIxPVkjpjxJZVoCh758ArxS4Z7pO0dDh4
X510uwlCGuD2BLhIyMYP3uOs3rMjR+Te4xjXby9zFcYHtx2NnozamSvoHyXFzZGP
zEmup8pu1XyFz4S+Adb//E22KIcInPfimXhDMKw7aS55btrz4g5QOzegWqaJY379
S57KJL85gXxPZyWwtmcQeiN+1LiHWkXPXXZKWAr27FIFtNgyMD7Yz+8W3rXgfUaO
/vVaRNWaQfTTo8A++/0eDom+4Qe0OOX/cNuoF69778M+LmovMxGKt29esfQBYKpy
tv+LAuzyJK3OTtWUHZwRqQYhj/WHP9x8VE0X9jBRESJR1eFdZ/cngxP2TEikPNC1
Ls7wWukzYl79ZpStfeaArSy8g6uPqGJcTrWOtJVH/Buvnrgw5OiovgM0ZtnzDNRb
xhvBbP0L8aWNKL67ejMJ7b7lMGnXL6jSHPfOHhHQY8LJ8EKhTuJdjgfkgJd6Anbk
aG1b0nDa67FKmmDXqs/AdS+bhaEBd3UIkHREq/DRLami2gy+IrShgAxg4UiwEQ40
VPTJ7eXZGHURmbdOXIoD3GIl7yWSZ79plY3x6z5bLpf8NO6CR1FW/UtLaoVgPa/n
D/3Gu3CrldZR/xKZlFRix2+0BCmEGT8BmMHoqgR70wqfjHE2HV/gA6/G/L9dZuYG
W6NzqcFQ94KwcnCUPJ2LAozfyCZVCZSZGokNoZWrtdBCstPcIR9N8IUncYRjO73j
oK83OUV/f8X7Co40MB7JJ8WQnrb/0HMNN5D+ggrC9H1CDshi4pYlfGrRj1w2BuG0
DzaIVQkFaAwc5n6VD5zb08uZrNy3IFZ27K+9ms8pr8869tVlE2LBEFlejqGEpqKn
0knlm9TtbyT4W7TyK3ztksnflkG3ft+pWQrts/nvBNZu7ZTwPcqF9yeIy6otc1/y
2qoEWhbUusSjcCuU5OjBQhwTHiJFi5PrnFIoDcAA7Y8ZDyQOKyb+ju9AAVcPG8jq
6DhCD6MCzo1Cn+RxB9q+jZc7I5u0CNc8qIf3zv/dCpEIhIXEi+buUejsPVMLS5bn
W2UTt/m0EaFnvyHAX1NEQic5Zp7GNM2vzNU/EQ4Dz43RLgcagBKT+dQzNBA3GBVU
WxYBKdCdqKdcjl0GjJLpwTrp0JlX4/3c6sLYzeFZm2KqeWXKxhCYSAx1tx8H2Q1m
nvvqR9vGwNaOjGtEOZG9gvXG5FS9RTMOmnrKpNjAnyAhFXwsYapwIR9m4xHB5jdJ
azN1kqrdgEMlM7WWdaa2AJVlG2cvpOgAVO36LXgkM+Q1oiPdoOnDZKEuCDhYU2Yl
pp5E5sAru0Y+rxm8j3WaJR1vMuwCTJfnNlGosCyw7e93NmJdlsZMYiY36wdpP4hw
GaH9bhhsSDEXW4ubSGux8IRB2Q3uQtUc2Tn1iCW4v34oCJ1XHFbXYMOiQW4FBQXQ
BR52juib7/dSM15YhhfbGSWBrHA8fFEIgoCaH1kF3ceLQVfDm9jgtE4EebRKNXa3
T4TjiSVDqnA07b7efa7h1EZGUPO8JGIWjfCg+t0oyOncNDR9ZAszhhm7VjlbEbLM
LOe5bOLyXVpVZAwoWhh2sQXah5/7FO9nWSvqq7fu4gs0eQGPD11jy+gfDLpKHsiL
OqxdkDTt+d4tmGQO+cy+W1mKSCVbC5apZ2jnI6LmmZ8IRRrGXnn2lgZtqmvIRTMQ
hKqzFVu6IUW2CeA7hFrGQ2k7MKK4bbKjBNweGJ+OxObyE/aCNMKzV39JoSjtc3Ep
L0cJ8ULOMFbeVpZEMmFkmOZLC3gl7BRZG8dT1IRbr1jBXdQchywL82BYVZDTgZpt
3JxpvTXl1fRm3wNjiv01dVWrpCecWvRFJRSCS2j9K9CDQfAikvpctKzHrCsTIyQX
+hjJLA1erWTsXO5zv2JPJ2X0QOV7F3ZrAZIoARoGr5TDM1Rs3QvxOhrh9ANyEUCS
mbevACtBInXS4n238mbQVf3uTvK52cPTK2iZQPeap0nqlkZhgvJIDsPz60J/Bung
wviLFk/uwCMyV6caN7VWA5KFRwojnjW60DnWCYFIR7CYe7BfXFrbf1Be6uvKKIou
O1ruxGVu7H3gQb+K1VHJ4Z0fL37wlGIfirNhpTD5u5gYFj7Gt+IZnwc3eXCfRbfR
+qenYMjwTNIWgPBu34s8ndb+Lgf6wACXgUR/yFwX0/y8VuZCW3pDG7NLLYLjpO/g
fe+BUWjX5H8L9spb3lv8A5vz9UnO8qKnZ03Q0a7HYv4AzCK13nj3lUS+1MDVRakd
3REY3uGOhRKfIiBJ0udmcNk/QfiY+DJrCt0d7CdUSyZteg2VcYjCQe3J5uemgzlG
tH7YqUWIUQ59pc3GPH0SFKdE5exffqnh9HwCxpo5+UzkfITPjeXILqzRTN16uq60
rrgDR4lAE6C5Kn4PsPuPCTsSthB8ZWYo9J17QCEN2Fe/uXIyPc1DY3sx+yG3S+O1
K5qOcqzpI3HNmVb88QA3Tm9dJ4PMu9fgWfaz4lmfvMMpRPUM4GwjwfmXhNJYLjBp
CVz4cPwL8N7NucNua17ZpuAeZUnaKuPres+mXnxOhxwCZg8beV7dS7lYhGAiWNZb
00WMelFmwKZkt1wBHs4y6V4q/MRjHz9eDJvwhnEGSNK9ynLjWAmwsxL6QGP12syU
ZyhOOxhKDpUcdzLySnkO/YingWWliK+5tlW+VQMotM4N+gwkKhtLqLPekr4heqN0
q4JnyoPNOgs3VcrxsCHFvrLjo9h6RXy0YttgQH27AzYdc2c9unXtD1PNarFKU+m2
gnVEN9SCFR6PTykPIwf4ZuNPLyEDrTUSx23wFRw4Buw3ztrrKVkG0EbiKpBwhUjm
kWy6lIinPwR4xPsKWf3mmoq2OUBjQl4y7/1MLvmC52ZM5hXuYnthzFLel3OLJS/N
14Ta6Dcn9v3W99HJpcaZs0x73/Enp0o5AGnHVVGscOcXFzN5psp0X4IBce6cTZpR
MCJ6FBpI43cYUZo7A95FZei8Es9LiRkMRC7dFDJIGGw6ByruiFEG7/oJebTEQOdu
JctW5Bj+6cFX7xpjnFSUZujUzwc1cwyjtFPVuLN4Cv1iwfaMq8lqs1wT27thX71L
68bVypdXiAPS6Ite4LpyBoFrM4zUyUm/BeQ7qImPPKAmdfy3qdqGnxqGxidvAbr2
+5uM+4YUJR84ptESWllZ3lNmKmZHsKoVnhh8IOytlAFDfK5cr/ARjUR/6/GXcPaA
gNCfUO3P4WhXoKyn0ETyL3o4EuHyEu6gdXZRvYGOgtfJ3vpNtd+PDQa10uhFRv13
f7CzXB9lZBbt+MFtkGqxlJCgxewUvrDtNeskLGHGl7rtG1P1+Ypr2DWq757Azue7
dUmMDeXrW7CYqay0OaDqO8TbvDdFsy6qo1HGkETqq4oS+5BxuUCGfjJ2gMwZ+Hfd
qGVXYJU1T6YY0x+0ZEb1cGZs1uv/Prx5OGclb/VCJLrGIOqlRYLIRRyvvQCeXA6q
9Jaf0oWUEqXKzrFXdLKdZkIofHaufxyVaDWoWukyw+sgdrfDJzzlWjLRvC9GDKmE
ZN4bs12i9kEFTGN5osKgRAiccHhISgBrVFnY4VD71tZEGUGKGMA84Lw4g9HVO6of
7OPyHyJ90APFfe4XhhKIsxMXoAg3GCBZyTWiBPoSM7wzb0V8Y3fmZ6KHUByeXH+G
aITqvmA/Pn+wGR3fTCVdn5A6nqPN7uqNGKGP4c5XHXtIQD/sT/oWEor9t2yBRB95
+GT6+BIOS3SGtMYFDhIgfBnGJpIaUY2ax0D3Svh8UprKh6Mu1T+NoHsznVH0hxNY
Yf2I9nUSfV3blLk6k1fLFq3n0Y2whukBvuMd16Tbq2jdPL5trr6W7yfc/5odkDUQ
E+QjWGEjA7c1B8+06Vy8UfGV5zNCreRmRNf6NhhsWa3HnxH6gLZJGxcvwPtSkiY3
gH7WMG8eh+MQsRD3b3jjCPUGBJAjlhBsyHutqaiDR77eCi9vUuJJ3miJHSOqwAX5
rl2DeTLIZi+jhTfGtf9kiEAx8geeWYo9YKhc2bBpkIe38enQSkcyu9O9NpR7UWEc
4voLqCwNAsZUsy9TFAu913Q/Vj+0kboXKqZv+Xl6jAukq8dRevD681Jx2e15A9Tb
h1TAtlIHh42lG+aI6BBW40idF/f/4oBE0PRjzDNBxlHYWUwo8FP3332WlsALGsHN
DpUmUbBu/lAXEoTUbkyKTCEg1KbwN9KVAYskkxIhCZ7v++AYpR6k0iqSifcmzOCO
zLkOBzQVII3QdzPr6cfHoNx06SFzY7nXggyIBdBw8Cf1tTVTh6HebhScr4WMYWz3
fzIVFXW5ZP1q33gl/0ORBwHi9ihW7gk2Qy7wIkUlK3eQh6feML/HSNrEMeHa+vgX
jNuhYYPpye6pFwhhCgcUBUoUlPeeljzqFMz+FgMhzvKVt6IlVMqKJ7HZQQgusZe2
QiNzqIQavPx/3LteUwvEQJX3aLiWjBTlutw8pgzd+ckRDKOykeQ+UVDUKJUTUyt+
ubvRlKmVsl/tGQid7Ql+YHkNmkNkTNR63zo4Hn6tjITvjYW/uVCiSSAs46Ysgnd/
ILXzQRm49ZGxSGm5CCq81IBwF1Q06PDVpbIl9jmsiIPovSIpHFDyfgDVzBMtmCsm
HERUND5lLgyHJta4vJtUrHaDtw8Y1mcKAF/tNV124fe9I+ChI/A+hqsViuPGGr2e
WqoETeeHJH3NRdrJOYVv+1CYY8sqbz4nVlk+UZgERKLnkPwGsoycWoTwIxTobV4z
L34Y+0O09+Bqf3rDIm+yNviPsxv7pHorc7VuM08lBfqzZT98l95bpcAfLiqb2gPU
3zZGBhoPsOpnAxI8Xs5n00/F7DGsYIr67OGmslcoBx4PYUiD0q/5R2rezAVN1p7t
SmjiSBR2eTv5Bxkx0rNHpO8R1onjk/SX3RmIwojBlqFXPXsfKzV1U8oEPLCe1Qpk
mNFLvNifOIdR3TpSSIhHImqk5AQq64CL1wU4PZdWHmCtr7wNqYJOUfi6GZvwrmMA
xzueEHZDV5i7Bm52clEzijAeBM+dxiPp/9m5o0nxSqApRJePUScxDox2cmPTHlQS
52Id4sjl/vYCV/TxpizE3IRTEPbJSAtNrrIVmeQLhcrRujRQYQ7KO6OmKn+8duiV
FgDgh4vlBBe28f46SmmpiUlF1PyKPPstFCn15+Hy6Iu77laYmKmuy110mMqzUltV
QwFlP6mdPuhoqhYBEdb6Dk95wr1E42dT/UJzRKcBpVIfBBM3TVgn+4tjiQmkJWeB
E+lUDgYxam9SQmfA7MERuBEYOTADLVlExcMBr8mHbox0yLDc0NoXcSEAMaf4otps
vvpl1pz0dNHZtdEVt9ZiT5r+o3/Onif6brjrHRtwS66q39f2nGsXGGIpFMJI5QAD
WhQO86MCWRkm/jXSruwtYvhG9OYBTooxkUOfMzId+9hMbACFtRI03TmWPgOfb43p
8uTb8k1aL0WcAsIaULVxP2mkppZjH0PZEXkuqUSVpuRc5MbBvGQlgcof7A/M3ECl
9wXfZldL7xdiT+kqIrT1d6G+w1hcGmDjZlvZq0RSRo9JSee+7/OjWaAkUlw2Lw/K
pMwwElQ4yFdVdhbr4VGsMDUfFbb23mfXpFRI2T+NzcrATxxa5DoDaAPNdjAICPij
Cp+7Lkqlaz9gN5s5gXWm5QwwklfGQWlz4A8MtEgeru6O2ITBm7U9tIYQNsAJxy9L
pjXeIqbn/Eli5L8/oUyyBUuGtb2EM4qulEJ4fthxH4xUr+8LbhhRZCRTyBVFcPct
v58IfRSGWDAKjW3rMkIIVJTGvoMRIe6qrpPvmFrzaP4C/PYFJKup5T4DJRDNb80W
vQggUeBdHBCDpGw00kYWiJrdPGlGfoid2TEdMBiC+hhvL/nbhe44T0bjf002Ont4
ZqGKSMHHrW5e38Sz8gQ7sVd08y0sCEv1a1+Ws2aSR1V9Lch+r4vH8wlH2PxFEgF9
M0N9sH0SWD4fLbRLjO8Id6VSoArvlbZtIfB5XshMlq2EqoRbhdj0o7N/d18l0feg
++Z0QEhJ0wEBbFqc6aRsv7g0Tai/WblKxfPTDTiwySALN4TzTb2cLrh+Fr/xadIq
t5v41ZH4UL11E9Qs1hNRMWd6tXFfgetDV+r3LxwLXvBMetJVrVrOSheFA/n4sT6m
RRw5ZPK13aS+gttkIgaJ2hRtDUNHdYaqYA9o1R1SrqduKcczItTGXtvcAo49mGUU
CPUUk95UnYjDe0KzTPrls7IlG0PDsCB/Tu77ed8vOYhzHSjltSfxYfMVwzZWfCHX
sePO5WUPCFSXGA5Ug0xAdKEfz4ZZE7/A8Ywf2IWGkldqZC/fhtiEPpNTkyXUoyyX
R6GQKQPIXgzIDgMLeRFG5LKUZtaxjEIGVoBhpnwuaIeOk6iOpYsAgdzQfPIoLyhN
4Xw+LyXnmsywRVLG6ahkFMf14HSKh6JRIYwgxT/IPtQ8gNNZt8/togQWZJ6BOXiH
Lc8OTTdRm7Jb2vYW4FIWvM14chR3WX3jsKcSko/axlYRqZVHwTWwFIZ8ZPrTPhda
n1EFkuU5YwYY17WQHSp0ezz7E3iVY7EEPahBF4PLJwbWuoRZ/tzxu4owJMIPvkco
c0PBajdfK13ULZiXMLSBSzvOgqEiittNXaJcVBoRIXiBgtX9C4LG/Eaq/RB35nQO
KGCPT6z3i9lvLXTbC0Z+r88uCkTg/UJgJuUq+lhFWxSKkiDPLZYqMu2sNv4AeX09
yQoBeYGbZ2hYEnptp3nlnlwcQsHX2PA/DKrJE/kVki0zDbJ2JGe2DhNetBaSkMIj
owm7ckp3wPUR3e3JLLacX23NezUhj3xLFWaueSPJhSknY3c9HN54Ug4yhFgQ3SK6
eg5OT3yLkVfhvhg9+kgQgljGLJYVMO7Mqi0P3O8ZxxWPXBx6XZWtQKQlfguR8n32
1hTZgPOCsJdE4rBFxU1ZC7a99vHWPdTgCeukqlQ8C/hMFQJoz2D2hlaX4V4ubG40
LWHxX5XT40oH88x0K4+G82Lsl0vi2iXDWR9pWz3/tPCGKZeWnWdYI8P5BVq0BUtG
o3twefB8ADAPQw0XjNG9ykFvg26qK4QquekiBl1Q1YRAeIab7IUXH28gVv9RSLRw
rQpXXQKQKX6BJiwZ8/V7W8DUkyU4R43Um8e7rZwm+HsH3GYwFEIilAQ1bYfPqsJ5
74y/TasdhhsT0e3c23TPRAnSJtAfcQT7gyt2gkUP1URpcNa5Kpp+ouJchH7xLCIU
VAHI5EfKvuPXE3UdcbIleObLGc35fpRjdt45fFy6Ylg/Uw15Z6WWZW6cy0IuLrvu
bUmoqbWoiMREBPIEWhxfkjW8PXtCpDkz6LC9HCIyrEzEHj9jGBh5wA1bD9veWVuI
+7BJ5hraReFbVnEC315LzsCJnNx5ERv0ksx9Pv6zUY40uftWl6XvA0mR+f/BntzG
cI2fn8fKfsa9znhedY4r6bTfoi3Tqv/mJGX8IakAXib6cy7L3BGdT8wrGhB2fecW
KPkDk26gwd4BaDGja2hBMM3bM+xyigqR+OiDezuViImbQUUrp9j1vHZCLhFMnomA
6uXh1EWHQBglWUmtcDHo3euCX+2wUt2mhpyATjgIu4GOYaCJmQeEdGCRqNjRw56J
NEchx7nTHalAl78O9SaIuPdnNzNa2+GVpdY/EZ4HmHsPbFPlQMAraLQ3ZTN93Pju
VOA3YZJNnRYFLVWlPpE7rU+UNUolkpIR0ygJVx1/+Q4c/vRLEWEE2RfgQvtc2xSi
+zPRW/DRkHM+svg9mkufspCkrBxol0X71g6NeJgsCkcBB17/f9dFEkmLb9hcD5rI
ppbrGNN+Y6zu5lSWecSHSaZECbHQkIxCiPhNBskA21vVkAfZ/vNzzxcTX11V/mPZ
xHqbQgkTy6XUkl4RdtePy4NH/SX01lVVGwTWSQfu2EqTjWZVuHcdeYuewzRMDrWA
6RLmyt0/FUbTzdiE8ozqV0+njSpa7N5e9/UNPT5iRE3GQP5nETzjahCuJm2Bq2JY
b0qNGT5/CIQUAGmH+F67Bi+K5D/yGmZ4pLSYBRe9s1pdS27DDulIx1VxtYxwToI7
i0D8PymYhVKAn4k7BNVpDcIs9RIqw4R22l3Po4d2gKsZeMWKmvhr3GOn7r+8nMkU
FJI0d1q1xTgueGb468T9E7CqALR+rf+q+krYBWDh/BUeqXizG3mslZtydv9zCFMm
GC1T1ILluzPd6JrN8trdEs6R44bmHWgFaoAJy1zmaDzC4HJdXmTMAfZ+S9bm1sww
LFRe4HcEoIAyDJKdx32JVJqqjdEx8UA9BiSSBR2u5troOr72WTJLGOQxcOctuJmE
na1THUwcu31HRHQTCDbBbFLH+aemoM2OYn009BoYxpEA70+v20/Eft+aSu44ItwE
+LPkO/AJBUNtL6JNFD0ep4VC0NdBLuTw/7r2ChPAigNykm14xqB3rXHqonsoYZxh
gQ+R+pz6E4odJtfP9kS+DntH5caxkB69o8ssu3mRJX8DlzakaNNCcTtaV8bj9uLq
xBTtIXaCQkZ7WHenR284MAWkVYCxzg70BLP/u35fOzHFeDwRSRIAz9Wt3pJS/tWP
AybCZG1V55eFK3t07V0Zu/eeJwy+VrDWIMl/Hts1tIG8V3B+f7YEJr+45+VkUdr0
qk7xcQcT/Mvd12mdPzqCZ1ULi764I75yZAmglQgJCwdtTEl6Hc3ULRBnJ/mRSqOZ
BpbgrWVc81QfcHVJKdIx8F8ZvB6UafyYEb2pMDYuHuOFV1uJiG0n5X1Pkth9316P
wbNKmeUrFw5nE0X3OXrm8JliYkEmZeNisIi01w8vsH61kqPgxhPqZrhYDc6JJHF2
Sso4FVLOwafvsIfDo2rSGU1zMUfKbkJcNfS+ArcNzxikbPK9YPuLMWnkA0iXo8Qk
4+cPNm2hzjMAM7coJzxoC5GT4kJgzNbBW7NkO1o7+iF5pwUw08ftURlIveGaxVFf
Glg7OL8xpLdEOb9kH22z9dfZFeoBltpjRhEkL1nzn4/sXg+oEDEyNtM1R9fc6z4j
zZwV/rW09+8yaJzapLcTiGmNYvg0gOLThcwLMj8iK97qYU+DYbRpHjWtb9HjaQIo
v1bk5CZuihmQkLUJmp2eSh/sjlTWS8CCWsCaSE+OzNmxjM96Tc1gqV9QlhT+aZFo
EuWByTLFSq0iFQ2WtI1CtViQ1nMsrL58YEarh7oLhp3UofH5GSmr0HQ/4tbjuHjl
TSO+tVGb+D6GQY5jCyEbgVe7wMFKaeGOav2VVqg7ZP77mh1zDlGmXS5IiG0cnE8I
uwvXZZY806AmJy5FCtGC6Kj97U/fHeJFhyKhoWJFZMWRv2fFr/e/vDz25ycjtd3y
UjP5X+D/zyzdlAZjvhli2HjkIHVQpOiFspsfGL4vm/bk7ljKSuE9V4bANJincUfx
x8YcLBxOQyLigKbEAqgiZWC2d7GU60OA2zdVTa0bLn03m6XA1EYA/yEpHxAHeZpM
5rJAn5wWSHFxkxk9S9Ylbh2bm7OZc4ovIT+y6tUHCRl/MyOs9FSejxOrfjIax9pG
R7Or2uGGmhovCTQZJEy722hu+4VCXZ7gARFQ+AhGZuy29SZ/BxdOAbq5MublakjN
eqNKYk7ENBmUV+JgZ3c+VBBCcdiz2pmp1fwl66CGrnE0plA/+dlZakE/5p17H9hw
pr1K8b5sa710MvwTDe1atS36I2GhDLYk+0vr76KnUZgUaPFRK58undKSjF+8yPrn
Z0q0qixtWvEwgEGjZEJbWrUx7rX44ZMwpb0GXhE7Pd6nzOT0pV+1AhWI7SLTLWVL
RuWDJbL17RP+XUmhOcNRfDjQ+Q/Lv7WIPgBdgw6l9O8KSVtvgonDTkghTt57S34F
0CmDV1VQcIEs6rTRZVpkreqrYI+r7Cbgvf58797Wk1Pv5/mBXGHtT++5jRyhtRWQ
gXgYRNW84+k2f3ojUFhbyk/fwBIqZYRuQEX8n9LETXzQjodyQnOF7TzuPkAuaaVW
8/LIoc458qNzchNB4pwFZ+frsb9rkrE9f+96WJDtRioV4ciH9KLGzFOWKLV++UoI
QSAXbJv8koPnLvwDbBlqv9ZMHl+dLLgOruRoYGX6f6PlPlj5os9WUxNsYpZjzym0
I9k+D2ZdCqWAjHcs849R101A2/Ez/me6ZXo7GeT6XQG3PpkwjfzmSSZB0lkoc5W+
JAd0JS/i8yRGG6g24al5Ix7Z+222zk4IxGk8setqrmJFPwJyi+UnoMgBB5Ez3qFD
tv3S+bVE9HgwTo5CPJ3xT7E/meaPUe0I6SAgU7Vdhhpz9mOKy59UGGlLc/xRX17I
gyiyW7kg0syRsJtFja/j+xW89HsvxtqVXjZxXiNbwpnYhGu1D+4VbkKBqlyK7Wlm
fECHb2l48hPFQfXV1jvKJw4LjcdMCZgz1u+2ZTi3JzeyrgGYOdrsv0WCT29VJzUD
NW4sLINDsOuKFExnYSM3UwRBbxZNqImxqbECrsLoxVOlwk0J34k0AzZ2Mm7xp5rP
d+EtudJCO5ERSdEstaTEAub1IrLfBfFZM3qy6wO8WTxIAM+9NXsKEvC2jChf45jh
AGv3mSsr73IEvXudMWRLXWczPMvdbOqsd1quhrew6068ybxVQ9MwNGQDHtRF1aVt
kPS1NL3RWhEDTgFdZuHkPioLR0U7dd9ZBBD3+4z4tB6CraNGUYibnJtipmroLxbN
HrhQ2MWtcSb01Q3g2+dvEqug3KdPTciv3Mslk+GMCL34dwOmtSsHHFHDkV+Oe05w
mMrVEL09iy8R/bQjv8ihG8CvCViZBO0/5gm6371xjYh6ZUPlBSpYvTx55Gu9E+Rt
T640Ji8qswz+PnOTWN57C38XR9GBrqlLJczkRdD4AdguwvYK2JPrtg2hifpk0Upg
wNFNSf70H6/cQufNQO1tvWeYskb6Zq/2eBXDtpkgZp0qINTrMvGMACzYA+KLfLYH
/C/DFIy96lxUFOGb+N3JDhz1FixtPxFePTxQFMgTH4QpyNt7MDQGjVEKsQyUAqZU
L9pNTHlTfHkfcYjUDwFDAIZLNrdLEMwcQJIU/95yQaYJAz1LMJwLroKxITS/VmqB
Qp76GjZEFDOby2p+244PZnCodL6cbm5UElz9E09URj0kh5qYV/UJHSolbstKSvtO
eKPurQyF3E/Mhhw3hR6jH/8cCNd5vz81eyZZ47sXbvXNPclVOLZmPBcap4UZm5+M
GWeiTgWQHpw7zj5/neckr9MHhVSTR40drhm4yYtb2G7OYy4ak3cRRyspW9cPFTUe
WfnmL1F45QaxgklXd94nr06IFeL68DaHhZ6n9WaFJonmBLyCOD2/S5uq7usWlIru
Exk7c/eKVSSfhq76Trtw7aShnBtdpoeanFekbAAePeuW0vUru/ImuXvewD0g2o2+
wokU4NOKhVKYBIkFAO6isvgDWEJf0ALFj1uqmfvuqCL7TPtvwHs3lam5/LIFce16
rxBZqY7BX4S/k4cYvSl4Mf+99a1HuCtjPItx8pcd8qsKdatWqj92FAENynXIt8V8
W80PV1N1Cz4MMFj+xBQvqT0EM/eLiRthudHlhE6SOt8K0rcjXNZRdnpb9/7qyYFc
2nvo6nI5sTy27dAEi9/a8IDA1al56HpjZUhCOZsQXXdCIWYCTU+Af5JAXdOlRoPD
XExEiaBzkLNnY1iuVRQzo3G/oq1TL2gU5HKMDXE0rtDVaF9jdo4CqdgAkeY7ur+B
laNwKLxDsUVcioyDDTPLOmtPL6gu0KHJ5iflL3Wbz+MeYcntNehl9EQ2EDD4XNSg
bdgae3MzF2/CdYYbrdO1IDAlQiPoPmW6gPEFe90WKsDtX0PDBIUhC9T0MNPFCh9E
UY4AkhM+aexwpuv2k4QBCBLEq60sJH3Pb8Cnhi40LtcrkybTtWSAqTMM84cGvX1f
UCYeAn47OwBXnPimI3b70idEpJcWYUII9vvnOSsQoTB9RbrX9B8uxM5u4OZ674nm
qPh8N4/jfP5ydbUyp1BXnmZCSAeVxwqsuJM+1VcC5ZwvJkmmZ6SsxXNBo93ofn/j
/Y5cw9xVGhKTmDOOIhKJBX+F7pvZuK+/QxOQGbnogUPdKKkIIj5LhVmHVUauSNXy
mKPuAuDR6nTFAtJaxlw/joRE7Ye7rnmclSW2zPUME6PS9oZxvvVEv09D/d7AB9kE
zmd1zj5/daUjrT71cdlhAoh+dA7jhPWDpCXdhUM/gVTjtL3UOupapfPG7WCo6sGe
I5Y3EMFW4A7hG3X66aRAK9Q2eS8yu/AaT00o/OQ+sCedoScbaGQ77a8RwpA1Uh5/
++pleJQXgUJtwELowg7Lg0Ptkl+fQbsuAP/PcNFvGx31XqRdfK+TKiasRFJjKX0w
rMxDweyAM9r/UcxXNRk2Yy7M0bHmzD9u/Qi0VmYYikWaI3D2iK9gPc2hsSYUwwBW
EEYhwuG9yfwzQUP7KNPCP0LygwrNwvsk0Q5FfmFH8VE6RjYqPC2mB2FpehNn72Lo
qzM5ojm8OfJVv7jjw78xgefPMaIbzDoy3+F9up4TiZt6xXyHBenAP4iJBKG84pdU
uFKJVYBXKjpbFvMIyoSQGQ7ysJ8G5HjUuRiYJ+cvwljxkaoszxSKBuYy9wsRDIV0
OVw4wlOzOE5+lG6FeW5dzhqmfNzJCufSfFCeGxJvLSpU/85PDg2nR+66P+PHv6lO
WE4fBoiUfnz+D9c+K7A5ILKuoG68V/5WPMfvgg/VY4jGzgVEVhsGO6NvtST8tYVz
kD1gAIsIIgLDpRC3eKjLvb4qsSrO0AIoJcQlFXCKatWyNqzOaerHYAE+Nw2OFPh/
rpRovtSARhATUyFYI5662pRrfBbbn3y03iA1WhAiX9Rp0cImgwvq1G6q8iZI460P
542VSoz6UDoAkHUHfNSPYRsGOsfJ2xD2eAx827jqMYtcomhnxAhTtHfIzyauGpEW
75/CZreH/g9v1KK3hZaW1YL4bMbrEljSbp5a8nK2+8KtAyvd9phzclTTRfnp3w7L
KhlNIDWkhvvRbEHpFuXi8XmtBogo3FghKkxkh3Pzj3tpokB36DQRQ7TTX6E6qJ7D
9yWyb7KIf7RWinMd2PEHinlOkFz0s5+9Nc6Hs1gpjv11hO9yjYEll7JsUcT/bvDu
KWMCTGh12IsjNdLBV0cttTL49O1sf+zIJlIsRlFfJ791F1hz+0wTIXL2QVZzlsFT
Xab8sdpczEVMaLocYi4BbP4nX+AF7dj8jDDVya7O7lm6kWSykMw7+mn99FIM6nOi
Z42VSkQCI1Ai4gvCqKFg4TIzJRzQ5ctojcPZOeBtSMPbokCqBo+y4tG4uoaxjC67
8DvtQm37wzvIfF/yW3iuiv5msNgmshekHFWQt2/C6wPJ5ovqlkaCrE9v85dvA8ms
hLJH4HCx/ICHOolr+uNUfv3yLVscoR4bQGitHcz+/X0IUygvkD3OaAD39J0Jz7H6
+M+wF4N5yKZl+CpAKK35x6IlrrDasw2f1v2IC8G+4zuHVz+6qLRyJ705WJN6hYO1
D69RtjcLv0grgqTBsNGNUW9Zgpu6TvGx4ShNL/ifqAyzhzP3KjDOWL+hZC4JQ3Lv
Fhi/VsD0JoPBPB6tKS5eJvvPDBZG9IphKLJvdpey1cJowcxk6WhKRv6kaBNGXRNC
bJ55dlALW9daJjrJ6PWGyK6IYM64sg+rGJPMsVmVhxzb5zpqPDl9f2c/SqfCPzTT
4I/BkznKey2fTUevovbmSKCBviI9UqJwdF50BMeSi4i9nqx9ilQNC9wBngJJwkFU
9EvK5ZoE7PI51+DrO7ZUEOK21ZJaigiRYwSZNcoeLrLZcpcYjDdxlQ62KZp9LyHa
pf+i7I/iLMclAf2ncZa3B02gALbV5wLiUVfP1jggoANGnC0U/+7yM3IA2U2oFHsV
idIVo0bsrzXgeR8bhS5+9e63c70Rj9C6icQxT4drNtXivhPzpVWxDZkaFNrKtWAN
rGBIbD/+P7dPnYBO5Eo/gpejuNolg7Z79MK/IsJcSaeEs7V2C1FjlbYO6Phuo3vz
1i3GoDK6zHIW1V7CW+oTrUMIfahavwvziIMb1ewQkaKPBTBUtWr1WzivgdTIdr9o
tpn93Qt3BgSEy6yti2UzjkGCLGp2iEgBZJ3G9vt46IoNd5OFrP2oGmcKVHDpUd0L
j1pOOyTaL1jmS97fro1jVe4CJec59azmCLiJIJFsTMPpnLNvYPqndpzgAMmRiKYT
1iPgVR95OyKyqCHgSmrChBDst7lXSTKXheG6kdwCYHHCeYqUrmzpETz+gUpD9TM8
hVuhjYdrrmyAkNf+P4Qv6SY+GnyaHfsVUOPCjz5hYun+79IxAecdm4d+CD1zt75E
cdlE555BfmTcJbP/K2L5eImrrE/oCEynsFCgjv/xiXbj8aEBO0M/yO2wWA4CQZAs
hURBNvVp+gou5RIBC2yk+UOd2NpGQZ3DObp259YCgKmFgST09uoLdmcjWYYZITQn
GA3u3C6B0AcbsL9eDjWv9kI5fS84G+Gzhc2I1KUu2bjaYpO/m9dvyxL1iCEUUp72
/wSa/REAPoLQ0LdfoM52uCQqY5AhbhxC4Hc2bFzIVqUDi4IfkrzZgFHIZspzUBcP
uGzZIgeuH9+tzVyofrb1wqrzZqXSWGKP2vPwn7oJQYkgGclZb65jUmztN1FQMHZE
gKemJvfX0e8bAqsj/9e4RA9YcK50uSXrkQhcDR6j8hUYSft20CNL0PWSNbdWnMQv
beN9z1y5qdEXuyL3y16ltqWz92Mw3/WsYrX8DEsBEW+szGoq/h3uiHfUnItQn6Up
L+foIgVV4P8NxlE15XMcPaaRzGY9p4SY7q4+U15gWQ+4hf774eCuzhvIlOCWSced
/dLCN9VGw+DZWuSHumJqU4Iia4OOtbAPiWUlGV2WE4uTK+n1nz6A4G9Ic6bM3QUj
CxNyqgHz5LR65EAlyjE/alYFaonq8v12XUGLW99TkDB3AlsCvqR5GZJ1Y+FPeI1A
vPmozvKvZTEetBOD8SOvdXhja5i0oqga+yLjar7IrqQucOShImaqD34T/47Q0NhT
9Jf8chh/U3GOVbPXDKVq1d8jFc+xgxxSoo8Ki3/9sKi8jcxhSkvbgRkagyiVRsa0
b3TiSRfRhNawMf9ioe13B0Od9vtbOxHe6VfFhtqbDbB1H6vUMbKLPEwGRqwiMtfl
HBO7Ulz2hgA/K5zYpFKWTaC1kJMm9ON23KOn1hMBrEKZFPffdO7wad2S+93Rab4k
aYNLXAwCcW8R5rJJYSYHGxHEqfwRMSgNIReDnWWMvbYYtdtzo/0EMBM3EhUUQXfj
xrxnNj0UiNtd1v2LkhDTynsbLi2RLeJqW2h2L/COAtEfWlUDsu1RTaTHOks5H0PJ
k3jHh6GJIxq8qni6rM2Om2fhEoiPy9XT3OG7qyCbFOup9bK6pPADAtCkohPQhHyi
cqIysNp4h7b2SoNRzqeaGu4fbdxCrjThtz825X4wrAgVFyG5Qcb/S2m1i79NzZnn
NLDVDd/pY2WDBs+0aK9s2DUdrZ35Gbi/1vu2856TKhxhnCJU3K5chr7e++9wBdco
qQsu0OwJX329zEES50dg5Jo8JF0gsp3uYAUDAURPJaRiVECVhdFT3Yz8/nPCmYuD
Oi3pIt9DGB//SNrUHy0m+izmaw6NLi32re9o460+r15WU8agTgUz0tdljPeV1WHS
1IJJAu3R30B70KIDPiPSiVw/zPAL07YdkKNnDQJZvpiI/p7hQHo+AlyAhpoDTHwd
NzqZvP2NCy2UMwFrCATWvY4U80PkRYzk/gEvengQgxnUK6ZafvHBdNITzx3Lxs6l
TQ1RpL5EFT7HPZm0daUhezAH5iGQIBcsGGGYMuGrYHtDJdcQL21/eUTLIeyrmDRQ
mqSFXi+urddZZWF26loMDhzvA6arj3sg8g6Y5JJ7oyDrNKfA8Xh8T9Cl2WBXv/fl
sLENgwR7Uyn+Q2RWfubt3mZAcfwLzi2AiEEBcpEJEGIF6MOHpPaXvGAZ/LfrwXsF
uQYNRuTkFUQw6LXhv5r7GW8rdk9jBrR7eFQ4apXgbzBkUocOLZP4xCXSFeSu3vdu
1/Fywd2W9GsOXhpxT1xlt+hD26pLVw/o+ZOJfw64vVZw3J5/EgesQpEZUnwgjbkj
DOCvkczGfgrgs+shcCxIUnHt7Zi1p+xHiBE7TY2cI4OUxUaqfap4qPqkzlSluGLx
GMlpYyGI7o3GPfEVX6o17Kd1DMtyOoWpxSljWghNi+y1AendDFlCA5+laxox/USB
JBXBzmfuoAH6VayH8kCsfnw2m1DyllF4QVqiDIiE/GrW9DFdBJz/BunZBv6T3RSW
7Wt5bYyazxTJa44yRYx8o9MxdhoRaPfzeCvccMxCLU4ENpfyb0vF4Op0ZWpWEQ8k
Mwk9woXgxjp2e2LZF3w6G/xuz3SMUK+8Vutza8j2YI9bXzpahzaTvp/OVE0e8W0Q
B18GaQ8CTIBoMKDxEVria2zCQT9sPXqrXCol43EFuvxAuS4ZJ1J4Thh9RCxHMZ/n
7G8iGy1hbIQnZjrnksvf00PtG2SgLpUU4l1llypO09VuYC6mTraGBUjXuAqpTAYu
dbjd83zy0GtwRgvmRmEbgxxQAuAmgI22wjcI34yvMGqWPc/FQXrWhJFgylVUjvb1
dUSRasxkkCe5vSCCunua8fG8Yvqy1GFX8Yj7KBjpfL5VSxr/7V2Z9vjgTqjAmSUF
FR6KBmQDnUkzk2c8IzbIDF35zLwK2K/t78bjqaLyPtutiqAvtG5aLa+YH7KH6YCx
Ts7D2d9EQHdCRx9WPY7q/8YghI7nx9bmJmEXPlbE1WEy5wnoggbyfPDdu571m6a0
rCzIAxX0IgpVK0RuJ7ZjTvSL/qb4bUku6syroWIDSZo2OjiA5fCYGKaiIbBGoqfx
55GGRn1E7hvmRaDnWsSixyImrAwwFPNNSNJjNtVaceYZ4J/ihk6o7vPpLGyz1fJp
ybaVCZOktqlfd2lF4uFatrpZp5BitRzuTU+WXkHAju6KKzKv64ei7jqPkq2EBypi
0IztzQCcqBmLQsG9KbNaXut5TJ4bLYxnc7dWanb/ohp99yzRvY23X2yW3S0b9kL9
xrCDkY+Ib2HYtlPM99YFTRlwpFr6ArpfjPR4dnXEQuqGsUjcaOsu5wcgmHKVHGKl
uZW3G8bBTJs/Gnxy1vSPAU9r8K3W/wThWYrQFOABKwTN8aZ9GRRuHEf7RuNNQGl6
rF1Gxu2YYIXtP0wN0doXvtVblgnXyveCeXi1Pb7O+PJl204O2onWHbmEh3lFu/UY
YBvm0GMWOWRBUFlxAxV2WB1AQKpvmO+/YvsTKzSoOqTLoKeXJ0Edjx9Mt+2ZVxno
5iWSmmFxYNB63uazS8fyAp53hqqSFafyY4zxTID6H5S4e8f5EG/hbrB/CyBRTA6C
zYUduHasY9Czlrt5ZzJpJVcVL4ovDHAnGLRPgRW+hADiIkGOSklNwv8YnuSlJ4Hl
5Xm6Jyj36Cp7LjdCELdpYJUaOCIfq8djK6A+CNoIjWzCj+N2ib69PwkI0TTvGspV
8NojJa5eB1QpRXhg0wPX0kWZoS9roXUEHpiDmNcB59iNTjAaz/ovSZIrw+nQZi34
npGyp3nbq0MpYBZAKfaq/6DElpUGobR/o1+jipbJE9DxueflW2sUN7mBVO+ceVPm
eaRKrfmYk0ALqZUe1PfcwktISBqXB37n0fZgwJBlE1Y3Wf9/54H//iQrdNZJ5o4U
DqsTIuYZiyLiei3fG0DOQcL7orhALwdM9XP8vSVEDtzF7o7Rf3i3gztrNA3qc0HY
tkE66zh5wJMkEGw0mVcr6LL0wBlGXUjQoxRPKMn1NkJIbuRwu8gLZWXa+AYgCz5d
nrjbIS+22lDHqJnJg3/s7jJeMKhbfuMYMVGkuBlr9BWNhvA62uyR+34C5a3zvyr3
WPWDap3ZZj6PTpx8cYYWjervNI+RY/lKbzwFeKvjWTXQwvkR/NTLXJvZ8tcpFWFG
eMh8kmYDCVLiAQZkg/Iy4gP+IiG79o3PUrpjkSLXPMzAE2VUqeVHh2EUJezQcIrp
i7Z0ibqO6i4ErQzKOY0pwRhSUPPcXZgf+/5fqM9L3ECzhSJh/bJ52qM74GS4vC+l
px0myzF+ibHkF7qRETm6D4Q/vhSu2PzNY7xF9/f1jTVsXnickmu8n/DsQJpQVBlI
RFidPEZLPJYBsnZpl+Q/OcnycqAvXiVOiRD1qsoAytBONZFxTV3UdGfRrRukOxvV
We1dOf8I5BwONYFsVFXJ+GOrKutPVnktoQww32pliCVVigDSj5KAjCsqeJKFXsXS
/wbQWjLLVISrJNW96sN17/7VX+FXWoi23ogcRwGADrJ+77CP+kH5XeizsiGm5HfZ
L8Hr19WLNCDC8GG+hU5giNqLJoa6ziKxjj18juIOHYSkcac+YjWkUY29zU9njdCz
VKi5Y/bIwv+g/0aztMVVEsy30BNkn78LsXqlwg/Xc90dk5F/a8QQkfSelnj9RB3i
qdkjwUtwSNltISAyTIcZna+ugYXI6M9isAfOyWIF4krinThPRO9KHtwcIbGL7X7e
XNCGoUQxpFDvU2a4lhSlPB1zZTZLO3SB2mGpqsUn4KptWgR4+L6zYcIXCiQqWn6U
3ogVg945u/31F83Ml0DsSBp+CUyxRFB22mlzyNi2svDXFWOn+EhGNbque5kraLV8
nDYOQE+bhC/TAaQgLP2DJBbFCaIA+5Z4De9ui5qo0xa6N9JRknmsAh7Pb7q7eWVg
tumX7AwwztS4kpPrPCmZ6+J9LsUkm3c+XxNpOhE8P+5Xre+ozkg63LkXhXek18Cu
2PMzSPLvI4Hi1CKrbmMY1V2dqI/6FupEiLJod2GPZxVXUKMSyYd2BKb7Z16NCpjK
ixRun/AGH57CgEcybPPsQyXmZtwo1q0GNEy0dc3/YE0y5Io7ch9uGwg4n900HNnQ
n+Kxo3wj3amcTQeQVcIQNJn9frsdeRvBDJEMvJ11m+b6ftlA1R/XAecAtkQOSChQ
lEWhDf9Bosnni9MdmLQ1xRWdWgNMlGF/4E7mfrGV71WNS6PNJP1D2VGAPyLsWZbw
tg2G12rr2HTVvnxSrT4/rmqg/vUsSvGTXPd36cAhVT7iUhPusDDXiKU2bQEckidU
EbbzYL4plgrQEExbALuLJFdiUUgP89ukagdAQ9IMsD823Y04vBSv3H94KyE+Q3c5
WSbSH5JElJFjU6pbwwaGocNoSuU5Ux0W/cyE1ObZXi6MMgp+/yBbsynhTCH/RU25
m8KZNUUVwxl1GvQ7Lf4EG97iURPZ/euKc8qNR43+3RKVmjQW2ZFYdyN8+GyV+fzM
Gi4Ta4yju3d+UUKAsZ+EIpnoCHBuJSdim+w5Ei4Hat7j2s4v20p1KyISpNw4PYn4
gLB+FjW5FlotCEgpVUDh8yG/b9IEdfSZnhXoUzCmGVDrjZuKxmlkbhHQBRvYm+C5
nsqQWkfYorWcmS+tmJ+ZaNghVyAx2U8h0TMPta92Nbf4dXzMfzt9lNUpFrawIRWD
VA7BV+zRiJTlgafVXoB5BgQe6PN1eQHoP5dPIBmryEUt4LrPeY8WHFIorxdjuPIN
MRBC0YbJsSBY0llxwqZ75YAkWvPEpZIZqVMoSS2OuTFDuQbOgSGjbuas5iz/ZrqK
XlvjXUAj2NFYPnUuSmKjzvMElP0F8K0KC+g5v4dEOOnqEfCuvvTmvSebn5jtwiEa
uHrfWwI0haTy0/ooBwXQK+6Plx21ulboq+zxo5Ku1r9wX7sjfBNaBYXmnKmLaM8T
7/SVbIvsIL/4g50127+rbq3c79m0Lg1TNdw28md4/3SPrBp3hZ+I9vvSVmleqC11
nhw29nBnMIUFK0yxBGkHJcTddEjtV2HmaWO79v4nlk899O/z5UARbheDpHNlSPzg
2giGSgU1kMDibybHD759giy+Z2BaaLbOs47HqluHOlV8YdyIryp5lYQV4+l7H/C5
+poT+Kyx50t5xzn3BtzCcCFGBRb7mRsJcvU6UdLuu/Lt56McuxyEKT3ccCMoiBW0
l4UBOCR739abU3mhBRh6IsRLmINStMpDVOwu7yCcRRU61VNT5x9YvWivl2KHq0ts
5OmRk7h0m9J90BqsHQeXcfWLuOMGSaMqvQoqrAmiLuNqCDSL0PaSIa5VjSngs13b
qClH7FilAa5UMcp7Rq0iMuR0vgOUHTttjitdakIfDPaorp6J4YnszX2mUfF4RIK3
l6I8Rmce+BDqLDzQWpooXT+ipjuONMy+gXpTD4GlaSh5EthgcEn0kfFwVbDZ+yrq
q0M6lIOpbv6VY8swxkh7trV53EAlYti8f6kbTOPqrFvjNBfQu2CFWSpu7MqiW1KB
xmcrNGIDiGkisq4iLbQ+Itp9JoseYYYR/n7QPszAbOqehBfViDNEpHJ9x07147rU
sVHWCHUjUO/NeCLssHCuqc5NmtPs/zC+GSlNLleMeT/faI2vTh0ns+Ktz1WEc2Ff
0rXOmPxv5RiI3N+Lz2o7npOe1pG74WApMQZQVSP0jE8QdOmrQ7uEzGjLvT6VSclx
vB7811/1FbbsrqNucWka1GTe0tu6SzbP6nrKYPqr0Asr77zr8qwcVIdeDfXjQrEs
gCbyOUKuenCdYwQrQDKaDFaOJUj7FaOzBRkkFQjxXBnBXBctMSUHyO1YRFXF0lU7
M3WPzSh2o7OV63B2KMdniOVXQFREyfuL1zJ6pumNlOkZAxYKrlkHwiFE0SOxnJFI
8yXZ8k6sMsGKoqCPKLR3hIDfDAdVxGZ+9DGTmRMpU++I5l0+XlDe07pveoeXE5Ob
wDPyXcm/HcljPtKvVGzwHwsvoXqGWsNc6l9xPRr/hJHnzzd8HcO86tzY37QC2eBa
KUdp6VBvGFfNFT3r2BgTLF38o9FUZnR0/IosuY5RIJ0Q36yK1bjjdFPYOEjoa7t8
wAYSm7uI0osOXtMm1tN61s9Qqp5W5LCoy5bElq7aUGNKDxtLFnALjwOEgSEvjUtj
BSgDzU3rqjlURdcyiccXWKNCQXZeO1gsV9aKPp22yr7ql9bwHouinqfR8GRALNYW
4WytS98vHdTUWI6TeesVAd7rqV+xch5IoJ57CuVDbN03m3G63raRE0B3wWfI6ow1
XWG+r+DYq5Iyx0tLHh10seKQcCKE6UfVnHDppGnsYjN9Wb7IXWFWftEqzXNfj8gK
9/yH3E37Ce9ZufQIQWSheu2qKKy67VkzvwjeB/qXbbXiGAo8qZiykDfQvduycRyk
xQb3pGa3uXVvSgZJ1n6ZEXCqdeA/O0Whnt9latc7LrgGsBhsQkyiOb63zLKpHpUI
w3oX5dvsSIr3afNY2+yOLxywnyNIm95nR/g/gPLKCjgI/zvYkUX1uP6TU9lSXInX
kvZU9QSQ4j0u/9QBQWJVnDlJS7QV0aHQ+BCsyqQYS2jOLLFHLtTnL7kpLXyHS3qf
jRMU+I3g9s32TzwkIBSogDAIAWJcPzvFbdUNe6p3EiU2FkUFLgqUxR8exARwdZFB
Mk3QNbtfbwdnlg4Xlar7UPgytHrSo3AJjOoNeTO7pECGuvY+YiaAVAH/bYWEFpUZ
3jctMzJUY6lWlwcf8SMbCORO9E253NmiwqGsUn2sLlJ3CPl0aIdO27klApeFYHhQ
0ysj0J60ZBKuvBtysy5P8MDmbXiX3fa2GnvxSfjkAA8uL4XVH5AqXTZ3xTmYoG/R
rSjtFP8oIdpeGJt8mcvvDv2AyRNPzJ8ERTgAkBrHaEbVaxX/bWpYKlH9jdQdV9fd
O4CtbCk0zVAl2olCPdHdvGQ2p2A3/x54JdA8fhMmmcTHRbgUHWP5O4L5a/LetJZg
VPi4T0dXtZNsZ7wjFP9Pl4cq5FDFxgmbVJ8DXayZC3+hIX+qOID18TUHfHhi2Ag9
gmgXBsxUx+VgFgwnqZ59wy1FBAVKUzFy5jBNnP6JTL4JU7xn2Qb4aBp3RWqw65i5
uEWS4HvAHKuxA27CYCnO4ADzLz7Ss0ADEJkRlcodVNAvS8nS+8HimXNI/6H1sG3U
Dim73fEHj9pczjuustGgfKJXmChAWoCuWKLDxWmk5LGR1u5YkYIA/8iXxIIW4rgn
+I4Oc5tUk5nIXoFhipwNoKvghfZU1vnun4jM5jzx2c/WeQ9uWzgn8pHoCmrjFqu+
gaDfJeB5Vp3D37RIVatI0EyjWuJxEgdkThmCs9NgAQTFBGDNV7d3pqIq/vKslm8H
Nm1jMC/BTkPAxj5+ZFL9E+SCpWihTLimgeCVE5G2U2h+R8oVTsdpianNhjPo2qM3
lwEkz/F/fVf9z5vam2GEgSveStxG7aPw1iBUV3jYKV2OqZ/TgcFTisvy5SOIqK82
wwWc8p99wi2QKIOIoqtSAmRcA7QSf6Np1snoRFLDYNw6jocATvrfG79CT2K9g6Pm
dgD/+q1zICzKHHQrBr453GL26e0a9jBdQb/6O3UGfaouszbUylmTzj44uM8glNvp
GoiiHM8ks6+AV1XM4njipexsKtOEnT0sQk4AoXB/i6ILD5Hv35dMVrIhXspYG+l3
uxQXxgSWILqPSRbTHUgE2yYi9xTnxnQSfGuQ4upBRk1q2pO/Q0WWmUa3H6so5Pqt
MtOLtk6hK57380l4kGOZXGZfm2f194uFwwvLgDxJAvFFDK9JQrhT4fa90pQ2W/AU
5Vl9/+4osQmNnXw0TxccWdmSxfYrxc0K5MlWsHARwkkBhABn3lZfUli9cgTxe9CH
tZK90EHWDpYBkq2g16H24umZNIlOpy6i5SuI4M9uowgdJJ+7T8TjV9670NjDKcUV
HC7WC1InI4JiFo7YRnHzlOoht2XnEhv+5mbjBIzE0/7ERMH2wy2utsOCuZQnoEXh
VwYdEYpKq2wXxZHdz7jIA5SmtbgxrqrLc+NtAbc1RCyvDO2/LgaR7+SVBc1auYlg
yQL7tT60MhwairhpMzbTI+pE+2uZEtCPbyuqErfYEwt2oVzezZBASHylLzSVzOE3
2nYmLhXJqj+qPvKuI3JcRrhTkOjAN+gr6OfIc/6SkAMGj2nsFT2pi0ChxGVn1ud4
kpFL06n617k5miGdWY1gCNHZKVWyjqvyeNOu/oes3yV952Ehe/g7wQMVJx4BY/EZ
bv4N6vkUMJunIQlbSSKWr5iIsnXVVgtlgkFH+FPB/cVkBseOL5J40vArG6lssv1v
R4jsSFlfOez8vrIdIUDIVW84ddShKNGd3jZSGlScyzDf4kV+5at1LdZfPKpJguzD
rmOOfT1jtBvYbpcD27ml4uzHRLHwEEXbatN4J3pDMVOifn/+pVJupVT+UOZ9yPde
KYQhBl4GGggF5WX+cGVRgpn5mmyp6KZL56qZx4ovq+tTX03alDxgxiDZ3RziMQp9
rQNe0gOifrtD6+gYG+43envtcOd6bdqVqu/S4PZyMnAEiaggs4jGqs+Rz7PT/9CG
FdbCloLqDc3bfninn3HIishoj3Kob9KHWFm/XJE17diLpAPkyteshd/jk+86XC1U
1zAoIG5SEv+VcZZ67F0TYpO+BgcT7t6XAm6+M0lqFm5DZS5EPLvsOqtxSV8pXEVD
FxwAld1vWXRdvGv5awEb8CO1RkgjHlf+gYqZjEF2AsZIXfYY8lpCJurh20Ldr7Gy
XBEouAjJTtuou5Ui2eo978zrJwbOpGsaNOwTBZUw94ulA9fjVTmoe1MqEBaTwCnl
U8om8yCeCD/AYO5jgNkrZt9nrbMDsIv+S2IW4sqqAN5PzCe2d6/oOJ3rpbUprudS
O9YePhMq2So5fSVc8Qk1UwppCye9UbqDQiAP3HK7BCT9nd1uPK60sms7ALtqkeV2
Xjw8YWAfoP4flPL0OWv/5kYra9j8+cjnY77ub2MEhVlKGnN60rTixV16n2epLvou
OPtp7TFNRHq6xfl9yNaB6fs59dBFAImyFYf4JkrJOk1XZ8emRcIv9d5wne7pB0Se
mAx7iR3+u9KGzygVhh3tovJrC9f2grJ61a4cot1sWY23P6tmswS+N2qrKs/2TARn
1bHQdu2X935PVr3T4EvT8748/ECe/JXI7BymzoPUKXuzgOQNbU8Mbn87SJ+L4tbC
fzDxAzDOUgTdrieJCud2psEbpjbucMxT3gZCfyAkqDsOPIAbSph8B/0U1jzrwIi6
w68mN1NpMHPWHJj/BN1fUrK9SPLFKJQQLIfJK3OaXeAoRe3cIK4nTi4bDsLv2lYV
ntS7TpjxT7xKqeW7NrKLMdOqfnMQ8JgpuWfveu20XSgQNqzaILKTMMdqhQ6f90WS
G/NVzwwI5hchq1xSrFhXIrRc1Bp/wtdbT9QTzxvNrh50eikcQpiq8M8ombfLJh6M
Cm9LWMGcYLKPyxhaW30c1Gfg646x+nIBteBxdsa7fe3O7pGfO/elQ8DkvSTH4OZ2
9VJcQFoMOVunECqUQJqxha6/WVN2OqY7J/+3V15CesZBpwndDB0IjHzA60DQG+5p
CsX8fLRxgj8pGiHKLgWdZXGdKwWl4Q0sKaTEuOCwTqBybpcZWXMuetDqEPet4h73
iCY5HCro025CEh16mCkqs7uV0k2KgGcIjOQDW+V3WOyS/qgQY9cvIvMHFAjIf2Ou
9mceOOgaeZqI797q6B/ViMTx9XrJof6A8ZGErSX3fypbKdY7YekcqXd+fe2tnCpV
tG5bdYMSdv2MKArqPIhKyUt9nqIKydpHO3jXqHv2oWoSfleqoREXF7zV2f+mk1ux
6eKCa6zfXD91ywxleMfoloR1/5BOEsUXQsoSBXKkzbxg8eOZ5H1garvHrkMKv0lP
t4t6AnmohHsheWiHP5n3DeIYOnTYcR+b0BRW8eMvEparIkFpxy17/tympXzJ/3m/
GV1Yoz8t4oMdOK7QV9qpAy6cBLR0QmzdZjjPrpTJiMLuON5hTADL/E76NCS/vBwh
LhoeRlGlkkrHUD5Rmp+5fN4Tu4hObK+INRFEX/LtWLH3RJbB+Vr9GGSVjcHMKvU1
yoHKffKHk46KobK/RefevXpH/Lzw9GLkmaIVTimS0JbdtUptM5PX80UaotuyXumG
YWdCaGtwBVau9eU6ykHtrEC5GD4n3K+jhBWmTYk6K8YTtqvPODezJJav1uPs3/Xh
IttZ+2dry2YIf+88bzpVITmjiWsglMtIDm32+LK4TD6dsN1lTKcecyK3IgqGv9fz
CeZPtgBdyvJxvWf3O3vR0/StJmcw0k1VxzbvzdULZxc8WbGTNj4gqK8Gdt6XXz4T
v1dn0P7P6dE9MxzlG/Bz8JFj/abDQW6G6xLi7eiTQejc/6uP2uqfEjVAbkgohy/o
LOxdR/gGBgXFhI9/s3H6m+Jh398EoGBYIhNHGmAYmZ9Dww50ylLa8P71/O6SNE12
ozIQzzWOXifIph3Rz+aF9VnqNxeV+cZC50NndcwaHOKs3tp39/Hw8KNAbfTLjHOG
TBhtBVgb8Aihv4A5Euxbh+lF8XrU6YlZdbNgI2rWiguXC5/KsL4yO0odDl6D+FB+
1ZHQ9lRrrGNQEz45/N5A+xODpnJlQnFyjmtNpVmzQK6MOpMsa++pErWKwNfROLeE
IqnDu37e5KYGihS+NWYvy70tS3joh2R1pBm/9rdkG39hgUuCDK/qIRViGCpuxA2z
Oe47TulDygkZA4mvMioEWikSfyMQTZ/mG4UTaGfR9oa4OLOC3gQwbN5YWU+OpplH
PGjK44IYqz2Eu5VyMHoR8NgYbsiI2n/CJ5N2UTFOeu7ff9O08NrUWUheFjTrKeTK
RU3MvY8y9J3OuAXBA2ygOKcYBDjBXmb6DMWd4CnrJwCuloaL0Sl8EFObCbcNsg45
/j6lhi1j823qOI8rWqg5UyRUi5VjlQtyLOQO+ndpOU3xGp0Qg+OiCROQ4LtwZaDU
K1dwWlyRjr2ITZ2sfLre+2p2nN3SLlQupM/Lg+iScbXyg0gQNAQA3Z62WpXOt0an
eo4I3h6bg6wxknBOv/8/BgVOg8sqjbcstuK4yIjz2mJ9HbGzgyceH49Xf9vdMScT
lQ1BWguHNgZ/ExO8b5CyZ5VegT7miBrf/3Edapm6CfEupQl3bY/ja6n47GLm1pYm
RHNcz3qwc3eatDZDiFC6J7lLBIQ8ofkCYOM3+Z/Rf9DywIJQnkjZ9H1am5idn43+
egQR6hpiZl97dflwlOFvSDJhs7zhPRVW8BfjTQHYi5G6KZAek8ADMzo1Hxo95EpA
Xz5N7/nPkoT9OnP9t/6OL3OblLzU2bK9MNey07yC13voFhI5Tqe7/3trxaftJyRV
Aj3gYT0VwhNqEn8s88Cf1eGiFg2emR6mo1TyuKviFzo3L5Os5SJ9TWf436x3Uip1
sB9V17EYw+63KvQzXuwEX+/vhTo+g/nXupQjVUIDpj18v2hC0hWVld+T4ArQWB74
13ccZxx5eleaeSj/0gVr3N1Bj91V79Op1IIbdfePgQyQyhZoTOnJd7vy5/3mb8QH
Cs7oQkfVTWdDea3CoYbHdnmzhxAQ5eMC5CI+lRloalft6om3ZByZpEnzemjwnI/y
bu4q9nQSsaJ9T41mHGAjKJt3KqEG1d77l4WSx0JSRNxaW7+xCzbDywU/r2YvexvI
GdsRf+/4t6mdukjK4HCFSOcea554dIAOL/hJLUPUjTU14Ml41yl/EzmI9lvS6m1/
JsNPvwrQgEmBdqc4CLb5esLjVz+SuJTzcH8SHlPhJmmYradtwJ9ahMdDx0pHuS17
xHe2NuhAGbCwA1QONwXP6qLRIFH8BrlKjCsp36WNYW8aXp8wZQ6tJhgGfSA3w9r8
o+gwE4bFtdpZsLy+42xQPiEGTmuE8Pc/S7e81JDhOTnOcMoXKNjQNlbuSTBX0Tkj
lTvCQE6/8B5cJyFxMuakcjUVFBKLz5LiKtt2bOTBDZzZr+WzlokEg6e+q4JG5Gfh
HmKPP27t9yV12afivlC1QWtNE2/5MTkZ7ORUoJal24pEk6CdLOc+YdQM8o+sRcqd
1GcLvmo0V8DAWqIwZ7wGA0YPVsF72GdeIIg4KZ2hHuh6/fidlnM/FLghRvDetZB1
WLABtuuTN/ff+rv6g9D29QWj+xIurbDvtQIR5rjQnLFZI7OZyw4Z2OzLas73Vpmx
KumL6aZNgvI3NArjRxxhk0s382UuAuIPtLThtzWzvWEdgEma2zDqSRAavjIXJ6rz
LO/jU38W6jldytUxYiccnTLaN/1OQVWlQcP8hJWer6xQPSRAJhCeAwr23Y+a6kw8
5uOxcCjXsBb41q7PPmuJUWOMzWQTWhfoY0+TAKRyo/g+1IFKbZS535ike9wEuSb4
xeVjlRh1OeyKwSxXG4umHZSWxzRit0o1e92n5uWyPyvx/KBKJhitxDf1VVkKWaue
wlq0vdW6DqpCfq9w7IaL2jJJodsQW9SRxZH18ZhjpRTHxlSD7e4hbrOunDnPXs/H
xcGZpZ8lNYHCMygocjINdZ7OzhIaY99wydUm2Add/MKRPUHlJxol4b3dndAaAe9k
A5CW3om+Zx5haHuDpWpYRvrYFEPuZsneDd2GbvV6U0dhAAuJjJ8Q0B+EHYKq7DRP
BedsoKu6Co1J9o7ge7oXCNgXlMLo3Z/73dUANPviBDr4+0/zthd627IKzKNid/IY
k1IZG8t9VonWBxw3vlUhX6BIpXoFbPLniPOGTLb+hsfEv7KklmVJKRRESfR1oTik
E9b3n+++6Ushyb21v1KucjbqPfB67YUfEVaX1DO9g9yrDv80MFsj+uwPmWO0fQV1
Er+RZqlxwFHj9o+LMCvQ3WxzsDgQdibB6g0DRVQpATuhTXP4qTgHVJYAemq1ZQWX
bejzs55WdcC7BwuGU94HWPG49cfCT4sRWn942WmF4iWXP+EOXQDxfffmh+17jXWo
ntblq9myWCMP9rxxWABR3AY8vbs+IgkV1Uz6Jya3ByUWyupt8gHAeqvutrY8Dl00
KoI/wSme14cmZ6nRYblNgrMYjVK9SQ8K9zcwMUME4arcZJkzfwObjHEuDe+kVekf
TNfkA5693BdjcjpQ8tS7jF5CESJC2mWgAk9czUwiMYoODkL7vS8rvlyPjZ3+DpSu
hKAOZEtqG1FuTjFyJQgQwH1I3OWMYi494E1MPlxMBvv8frhrf2K4yxSNWAOg9Myp
NMf4as8yzOxJvY7xmGJtazSdWIOfRZhKV+0rMNsuHOhd+5zwOhZf5CrVcAn7sPmW
RQSZ3UwHbnrrVtNOQ8CF90jXaYt7oWVw6zBYIpO9AJ3ilUBPxj5ai3Jws1xLBfN1
sJdIHBO+ZjLuFBj7ZZ5kEHpz7el30MusRiMYwYZeAzPIgFmJzOA5psoNW0dcqLsi
J2AtcRBiuTqFkLQTWzCIVMIzI6WWdVJekNEMMGdzyIaiYXTnZn2/kTEOAr1LQQFp
PtgsukYp29PlRMpqFoArc2tZ013i454C26oZNRRW169ptq+g66X++r1bETJfUwSr
zBSQ6MRY2nIGks/49ZTd4GCsc8ukROVQucTmqK6mSSvZuRrEO9nlTyTgCJd71OZk
q5k8q5WKGGU6ZbBBFPRGLawN0Um2jJzYQq3GHIEhlUgO9CMsWEiJSc8TlOC1wskU
JQzgedfGJhkk4/qjSb5AhjDSme4FjHncAvBttg5Uaa1xvXmT+Pkn6IlyrU1AIVcu
1eqy9mx7qxJHL4DnBZSJBGwx0MMdQ1uDg7V0StKzu7SKHEEEP2HpxyIXuaIZYURb
G6h635EBLsMPIRPRNXtfo3Q5LTYm0VA7/7TSxD0PfV9ftZKATwcuG36tiLggFew0
goY84d29GTIXwrrLmVlRp/Vtvl/oGBguFZJ/AV8mIhii9uR2iHf3lCosyQHNVMCK
9soJbLm4iw9qd4Zb49VXKWw6hpNtpLC2MHttJ3ageq4SJNcn7E+aTYfVQEBnsfv6
+1GzBLmgasqEcL8opzV2ltMzzxA4hehEj8DK0Rd7r/lhgNSw7fGdCNF4gBv9G945
OQNbQsLpz/TXLRtXLqh3hljmnpFDjrqs5NtJ24UHG+lcLrDy4AuWsfDlRaEwObfo
YIOxzu1bYPZlseOeA075tJ20MLiSRyhCGHTQfEmTmCC3syPuDD/Uk5XFJCTheVgm
zNkrevfcH0GavSNxOc09Xpqk2Q2w6CoHJkZu7eggPo1V14Td77H1k6hKbrLYd7Fp
tZo5kp1fXVx8kyhzgQmAUf0DhuXRoPm+u3sJ4yWJNVbm6sb172v9kJq3Uslt4nR3
kqFa/vOBTo3vRZMTA3iDZrc4eLHRYLwYsuuaDc4PPAY1A6BGnGnXIBXBwAcQUG3O
Mqhep7aVCDiT6hg5xxtxsvrO/8Lw6IEdk8G9NbPwWwV2sCPTmS2ONXyFhQqTMW+b
6lwauDHzgeySlwcMGdFatMZj+og5UDtoZ3rGd8bQ0D1e4+C8OYprwdwjhu96Sg41
BroCzhcROe/9LzH/+ABW/7ijx89GqwUHBBCUNrTLlR1dwm9jhYN/13gW7/C+R53N
NSoDjdOqyRpQj6ZnzDCzv/13VszeHhPILK9QuQYrRVtrvO3FLLF5+8zywh/tw5an
NSA3ICyeAoBqy1ExCHkb9KzAk4/AODOmvvD4r80cIpjzeH2PrjZ2cef3RQFacOZq
klRB+TJ2gYbGcdH5djN2Ty4tIJ30A8Gb330NsUFhOG2+k9lU4h2AgDsyCmu139O4
a79lY2RLCWDoL7+kKSNYvaPBI70ptsGW6Pc3L+xC1Vh2Rt09xagQcKi0exmjSG7Y
VqlNH8wSuqw52S3w74eW3GLi3kQ1YGoDIhBkNSCUeo8UNX1p6OtYvJaWwnCfhDvt
9OBBQJTg1p0CWTMAfHyyQ380YbRYA4eU5ruCT/O671f+dys3PtSQraBfxNtP+Dtt
wnhi+OTs5vlMHYUc7Hnznl9QYuwF+6uGoWusRDUQWgxu0LkccdickfySdUCoqp8+
GZiqt0W5zL6GWr62QloVen/museMOhAnWRIPDE/rpJq62JSVtVq5v1G+cq+5FUMX
qthKTthVZ73e01eEZgTUvOFRcMvn3M48IEsRMWc/BSE58zKjjKWHh5FawHz4sIs6
2CCNpThvilXRL3uqEhq0NOlx6DdUARRjs6j2JvVI7rXg5jdWDtlYRCUY7P24AGNO
wxJ4w9zcHCtc6gskqJzo1qz3woeuUo+Y4Lqtu3DBJlMx9bOKGvKOPRcL+eJNZq4F
5ptHGf4a8iH6VC0xDinw2cuM6k7JS6aDjezj104M/JURVsn7NWx6p9IOJexhmAwz
dydKihaRtuwQvBs62k5CSufyfB8mRF3m6QTyUXxAUlMumHj/0LMhsp5lVAGmH7rK
x2u4du13tA5vTAkJT/M+hPAVf6KT67F7XPMSmH0+pi4Zs1WlA94o8z0LeZ9lQKcv
Wd+aMF9XUOkOZhVz7NUK6NREIuBUOYsFwgKs2MH9G8wt+WZZ6mmuGmsuBphI08Tg
/rZZxEAn2p03u825AAWXXnS4iOp9+SSs3WDTNE3Qw3toWCzAFvmcVGNeNPicsXmT
Ykr1QIFA/PR+IGbiEiCpmObH5utKV2K4vpFqwz5fYvwTZzfP4LKNZL8Ni2kpmjCw
kFbELquFthvM8XPOFt2G2niB441Mzjo+4CicIB7oEUFR6DWoy82oV20fMidzHssM
WbP8oGuXHeAQH+e4jDjzM5Zo9nLJh4r4G7HPt/IqKe8PZz2tq0UTOg6zjGA6kRKw
GpaI5WRYkjCyz4a9teagRnLWzdVpPp3Lu2K5y6AGnr7BO8lrS8i2dv8bGM6pfuH3
0mtAszUQ3R7HcOL0pK9HAfyYsGoRHtrgkcToFDVAeye9/FmUkAZbXM3GSlIbI2+s
L8jd9qdVMAhuEJDeQ+YR6N4Me34ekryPmf8+5w5s5vkXVXKO9ge3NTuogGOx5Lmu
9v5EjT1Pw6n6muRR1YsxKPWpGi+FB6QVdXyqUFlPcwCYchZ8INXqahzDnfKTZUtD
c5EhUs763a2r89mkEMg6xV5P/PVAaDdjB07wYqS6USJCR3yNFNMMHGQRM99kK0HS
aPNCLb5t6HNF4H/vrCJ7sABZUGMI8TOCDLWMwlxpOgJu2Zz/T8Jlai7dJI/q/3Fx
dzkUQnbcJ2Hav0GGUxnzBmf5o2IzHGgK9xNT5W7zglPcfqex9ZV8hMnmbhKmXcMX
YXzjd316aS6wtVW7H5EWnuzDVLCIqJXPwnXhPyS+ZwxAziSRs9aUjh9IrMv7GB6v
20WaoNhfQGVeIoW5slzRDM6khbwN4bt9saoNnLWejl7eGGxfM6hRHBUjUxhrvWEb
41Z3S60ElO1g+xuDZdjKZnF1dTu5HkwDfd5aewz74Mkz5oivJzcwd9jivmDc/nXd
/H+z0jaXV1K1KwTWwfq4WpBI3+OTAva77n0/uBg3dDGZqucIpO1ZR4JoKU/Iu0JD
dh+engpqQBbab28yWEAAMOfhy8tWMGKdhO7oJuUX2JoKI8+N0SOcrDCVEVTGXR4Y
1Q9LwnT8OmAJb35gdvUO/DlRoGY8HDs2j7s2qYGO7zEew2yOK3hB5kIrnh2ga/Cf
nz9WEwR9U3XM1CE2RtwfttlrgXkjV1eNy55owKhnvLcDwUH66Ruht1dlOkE/4Qeq
3ADBgR7sbBEDJhyJceoQPWHP9bNeVzl22UGsM4+qpWqJeDQ/CC5D+x60x+EdbC7w
tqU3ynEhB7ME2cnulGt0yiisYAIdaAkBmuBmeV7+7aOVbE5l0QtQimiXx0Qd1CQM
Rtw2tDRJfVB6+HsP2aOmqPhngvodxswK2/dLDNljMVeELy8zFh1/OmmMV3TGoDow
Ht9DANMnguO/rN0kNJ8MEVHXjVJBNSnnHnxBlTRVxzn2JHw+NzNN3pqIs7RBef6Z
oahTtl7cnRuQdyPcNM87SMcGsdGbNc/aMi9j/c1ffRmovaOth89X6Xvp58N5MvkY
zf+vfqaFllFyDzfWCVSmfM9+j/URtvmVgT6mzb+YGCYigwCewywx/oKe6wEY97g1
KttYSPfA7m/RcH+bO/I7UT4b6bIaTQdXynYrur2qIxVBbz+58UMf712EOoqJkVVQ
/RiSk8TRyrkHVKfXOeVaJ1W2Dnys+WRGJ1SmmtZQfOrb/8TWC+eu7YjfL7aB0o7E
RTvRQCI9YLs7n2SlOIci+3//3aXxHykETibHrR7/eZZP5oMt80BqitH83QssCYGx
vkCYe2qeoVwt67szYuM4Qa0JTHh/0/nL6Fhr5UREubc9Zc3pTaVgS9onPjnzI17p
cmF32BUcefh39UqTadB+pqnDPJPbhfvNz6iPT9BRwcI4AfkiySJrlHVc+89Apgek
twmu0z/uIc9hNlN6PI75qU65osZHC5z3wpcAn2F/AIhxlMBkK1f2x0gshVuiP26p
Qic8cp0AqnabPStbH1sAFIMHjpx69X7Zh3euTDeORQMERI6icCMi264JmIbTL+qU
5r5oH1K2TOt7VW73YVWcrZhpLjsN4KKZNPn1AZLnfshHbdHlLwjh7Avgi0C06LYW
VQTt+Xc/eHOPgDnCVBvgNPYx1GFE1jn2ggHR5XIwypQ1OTKd4KJL2ATMs/o0vOdS
Sd+DQn6KeT71jUfKSLVlkUk32fsxL3ahuF/a87D3J7pXRAseEXm8O4nB/0CwE6q8
Y71C5xqRvWtRJ6LK3Vjn1RDG/NDnSl5F2UtTPUjH5r6erqooX1HE+9zXw783/dW9
rXyp8MiHBvbsMaAlEBlGnkO7rT3doWMqhadLxNcqaSYvdWR/Q2UHKEiydrkpgI4A
fWVJUlHQUh6r4H3DJ0T1VitU+ajEFp1nFcBb3E5XCKML3RqOPqsiOlrctCxdi9lx
y+MrhBmtzz7fWFZ5ml7HwSckX75ql1PTmajmMOfbrMBHjnKfkgHVyM02CzuzP1si
gYt8skeLCtyrteWU3cmOffRCCyZ5PLls4EzpkjeKO4XjUdwuAtRrDqpyXEBG0o0O
qwruG/y8Va/055SF2+vqSVdgEGKB+xhdunmIV+obzrgWtHFaXKHwgs/EyxRCHkHx
AhzzfNPbszgAHCI7mtFvMqFQGRsQ/TQI9roRzEOwNUhx3vdIjh1ewk/GP5Ddp2gW
n5Q4IIHh7l4JIBQK/Tv2/UhOSc0cPFv7B8Rx85I6AFRBAYK0Ha2W5kDZRAv6RkKr
OswPIhntjJMjC0XqqAvKCjPmE5l0XyNdMbKoltFmGg0F/a2CQm/vtHL394BoOkRK
SM897FfjXNKonCk2CpCheKyHvSySD+3bVAEfAzks6wvP+UAkw9Z3SmnvfU5xfSRs
mk6LVExti7QiOSeH6hk8HW6tVxt46kt5OFCnH/20o8SitajJ9WEwDkhgtUc0M2xe
n0YQucYlztNbC1kILwyr2KT9fsP2x5DgnoDKoMxb984Qiv+ToSZM9EaLnRT96jvB
EgF/JkqxfOhkCzAoMHLzpRnFu5m74ws5drHMDt+Y4ATPlZVysH8T+cB8d7SEqH85
Cd0vvW2eA7eltOxBdXTsI061/7Hqr9d+DPI9nmJbExJ1S3c4rYXclxOlNVSPKLtp
fkKQIH/tCUxt2bIt1qMV1QEK+IPN4+GcC3q56Xtb/Mbau17+jdrEwWq/qQDknT+m
YiFt9RWWePp+GtVCoL7fMaHZoP1FK9Bb1cz+gB1kOKW0Bi/r4PoKq33FdSOleUCN
veR2tkEUR1agUEh06fi7nafVKU0AtRMgMn0zgChhjoqzvvGcwtsKFjRoZnpekOoH
CQe9ZwZbzVzjLxpPamenYVGMye55SLqvDngSBMO6K93T1cQRFCD4le6fKUjIcOJm
iLgOntsoygNB0ZdMVZQOO4j4kXeZMbQvCysOgt0WoeCOiVo3gmEPkgyGjlEZVb57
+OY728O8xi6q1l4ljo3FzQKvCWnzKAJm0WmERhH6iknQc36tb8O/lwLsFIUkCZzZ
v23b0SH+XmwbGgcWwbpTDKgmFXCV/wa+bxXAiAyiHvn20KtjcGyO/rXxjh5GQo4X
FpPnQ8qFfsRWkF6i2PY7FDZ4Ga6B99NllSNDO910GIKgiOIDxlBqjjexY512lpGo
49k7ZEOBKO3jYkYXvhavJvDePVwCcU1v6MtCj8dXwHXQdAGG+d4NtICdKXqUYo47
sTtztce5wl20Lg72HtLIn7dcf0wJvACsF+ULX2UcdU+pBpn/9mrywyhRbhQ5Ba+W
z7fAW3oCkgaqVp0239LY9CAsGX2a9Gj4DmpKpKEK2ep3umtDa6NfxlAdttg7Tzb4
S6706QQhCN+WY5yThQaQJkfjyRlxgsIrVTPqutKr0o2M49ruPxPGB0ke3F8FMdQt
I5U2ZI0d9HoVhOn8sTc1tAdLYXd/HC60oiK2nxw4y+VERyojcZdE3pnZhKi+Pax3
eqUG+Mbw0lQzQFR362tivqiLuVQe9/lvkK6C4sE966vSR0TKraioTAsWo+ENuaRz
9juKEiPpwvuocDFSgevut+DySpLBoXeoLhEfPx1OGWia1H5faKGA7gD8X/B40Ecq
fknd7ACUoYOVcrLlXhX9Cv+dD7ljcmmAgWKwmMmZCspUmCHS49FcaC3YWOnHqf9l
F0WvMmvl/Vyw2Swqb1boRHcayR5H0Foflx3FT9MbpinzI/xW6vKfSC9IAdXUZ3Iz
pVYEqWh52ZXtp/A6tC4EzD+/AH9kE/ucbCv3CDi7+wwsFL/XxsP5l8gl9QoqPcLy
BYvooO00IX1JGeTejHHcxUct+o0nkKoFd+rswAtGs2PA7CdCPjhV/jrDNmgPVFgG
AxjI6H5Wzcvc6BcWZx/uYMc/XtqHsG5jqh0/V/HIMlSaZfBjZU6/TxHL0m1LOxj/
dSpDgbb7ZBNctg8agv2NdkV3loFYtT63azmAcPh8t8zkXuAZkLVRdFxI5zbcjGYW
9Qw+/pITfgIDGRCyF3nCHZwM74uY9VIqL4ZkijzqdAWA7er4BJrfFhH3J8ykCwbt
seyl8SdYamMX+0UMWIw+mcYXT1uFfWtfe8pWHpeO2JXQel0o4FWupw0DZXUZo+fs
Opc9OOx7MNRP25ueboxd9E7Looal9FQzBl0KIymrpSPxsMyeQMExKR5pkUiJq+fu
QZ5rCs2Mdx52UkLLMuzsi1hWXSvi2JDZ0UAU0UvKuVcUzopErPABulYm05MGOq9u
hJVwNX0QZL334lAUmglDpOU71eixMM+slra9MiGIxXMCw/9JGU8K4RcN1LRBpgJi
YxMFspKqS4ztrA+V65nd2A0FdVg+nwcAA6wBvToR9E5edbLVPQ5R2fQMHLk+3GLP
pv6Nt58SJLWkdmKNKBDeZY5k+oQ/v8WUi/WcYfmcAKbNYVWO0gEqh+zoE3jeCs+0
D5P+q7cnxCmUwZeGjPWqobrm4oT2CMCNIp5tMwU4Qf/g+Hl1NDhVRSPLYvlA0Roo
jAjKom9/ShM766827bvV7yF5o0O9ttcoe/WvuoNwy2z0FKsBnMZN1UFEqnKiS5Rp
WuT2OsdaJoIihDeCbnYgzT+ZhYx5+q6tB6nYLmc1o3D+957lWHv8E65Hztu3xaZ6
7DFi75kHFnHNxmwYs4tJmGUSYYoIjuItq0hxAOr1qccXX57nuwwhW4SrJvMQ0P4z
qxUhowS2IPf96kCg34oXNIzPPYA248DQH5tnR6UUrtPxpaRfy0jZBugckOSvkQgK
MSbGpmmkaJtXoDvLSlSvLWAy3Aq0UWr114CdmoVIWjIWZgaznsSKdV4mgNWHb+cp
Dm+8KlNEtD2B25bL8pOuiE1ouuf3YjKgtCkVo7aKSz7YQ8oXLWKn0NigpnMP+ZA2
yOMIj6O9+UcEz34Kx5rdleuwvnAxzJB50qF6VNOcqkZCm18VB8Xcr6kpJzJ+Vw7e
EcnGLHg7zsmM/xDv/DshGHDcv1NJ+VXbbtcDdyH0dJMaDQZGOY6xXBO+qxECHGXN
0SsYM5IH/Fw5cCL7qgi2a/i/AQSHNc2wOo7qew0opaT0Ti17LAdCZ8fRa52gwa50
BQWjQalfi29gCpegiyLECJlMxCbUCxjcfgg9BMm78IbjK+Xx2jrW/G/YyObNh5/+
c52wG4xdlZ6Tfa1UJDzVTmIvpUc1GmkqPsB+WRSwFfpwAD7M9LslkOSHR/MVjw8p
pQRlA1/QqsWJ9rKjICih7mRtkgJkZh3RRlwz4qhheJlrFjXFGGykNvl3zOqp5paX
vv2lIayCB3TYakQte0qlpmZn0iEn1r4S5FzO13PWG6/DuIkIjBq7wVmPS1saD7lV
QTWHcQB8Zve9nTX/uK5ls2xKl5vDV9+KriZ/EFpiWfrT2mGN4xSTM7lazGkBQ1k2
JS9MPiZoesw5WB4YzUnvw/UyNlJydT9bIyXdNyGQWZ3cizYsDbH2faweq3ZYgrsr
f3rlYAD3UXZrSDKJkqkt8+02egQ/IneRAoNgRsYzVnq/9T9zYlaJoEC2rLNeGGmf
t3U8FSqf1VNXgWfrMOJB/g+t4aXBWXPKYH2suODhQjgDtI0JH+xhJ5w2ioaQLBDw
uVo+xFWYXWBCCZ0iwFv7Rj/JoSCgnXFHi8g8oJ5UmCZEom3xckGrUWNUbWVCfkEx
2LNZizA+K16Y5EMotd4VzSb+x/DGIz1F/xgdftsziEhhCKULMpBVYh4503x4cp9T
e/xq6R/41Klgrjiqp4kqQDk3035POWQ1f96aH5Z4Wg1tcEsdqTwew3CV8x4aDcLE
69D+BVBb5j4LrHn61xfINdEJ09uSb6plBuYo6CjztjC9ph1pAaMIfdJeSvMAG0r3
pEV1F+cFEqVqKMrhPBBHk91LKZou4cF5QA9PY9xEnTGlY1JogYP59dMm7NTL0eum
ahdQFTx+MmYLmmkH6VSRMnQgG5AuV23yKBTae/AU/cizLrc73KH6U8cj5yimg/Bd
J6jkNbVKbKxT4yQ9yFu4G9ZlAoh7UuIJSAAdHNtYD4vLIGo0zQH7FV9hPp8e1oxv
ZnOhPMkY21CXCCEXk+X0A3dgCZWHvDatcwRJoqFte8flsvn5WY8jfwVu+6An2ZNp
QUwMeYHp4NTQLTxqld98masE4K4LI+PqibNrlJRaIianu77495tfG4RuKsmpRmUO
0uBG9bg1K2ZK9eVIql6zADYFm0B9s09erbruMk7114CUuIDKCgzSnLo8ILTlt1v+
O7tr1Ycqr8ECnJoIaj2EDIjL9SWDSPh2QtCbyM8n0optEgbTRNhq2jVbXPAj51XC
2d1M5O5hWVD3Fz/I9pAcIkwt4QGyfFHKoyWnjtqVBDEqwqUF2KiYCeiRrp56mCXg
y4lCxX93ctkSgQdfvFOkKh1PtTnhaRxmiWnnQ4ZCYv01zUB3UCx7lHJ7t2FKZQHZ
ueY3dGY2oF3Kd/0bpqFX/RldI8GsQl6gTNQnk65HqzszMznPF1hceCjkLsogMCSK
yK4HRpWxONh+c724wXgG25c96HNTnGPnskwbQv7uEZyAge5KQqU8CFpQghALUskC
TaKKR4Pws/OtNszkWMCj300jPllgG7kQYmF21rI7cWrUFxYkK9SxAXydA8JjO/eq
fADOcdUqG/4YTL/2GImbV4Iiil7RfKdE04EEaIHN5HDjtyqza5rprwEB14UnByz1
MQupY64JeuK318K3r2BfAj12Hsc3kvOJMuNOeWCRk57eKEW139CUwik+6Fknus0L
gakoMgfCoE2CqzfL6Bj58dkNsFo4jFer8dkw8Zz+S9RPnr8dpnFr2w6J6CgruE5C
5FPgu9rYTR2w6dR/BhqM5XvWjD/gqqQtIC+Cga2+dgYhgF2QTlWq0zTzw8rufhty
ED5cWC8D2IYRYL6pQd4XQFYjua4MpYEjdryzeJfvKig+L8NwSXSOdV6EAOMLf7A+
kB1Tre2T7Nyqe2plTQveayPxOB4K/M79fpx7smYWSbiSeYcg2jLX3IE/RZzZW70p
fNN61OPmFjZdx6iEyN+SczSy0GdO15uugcNXhX37ANdWzFeQCqBwy0Gmv0ay/oL6
EqtUfvbz4uqq0SePd8381lCgqyaC9lyRZLEQL/VjmtUVGxoW4E3BlElls5mK478f
+nNS95cIdXgGv6fuHyAL2W9uSHpLkFcFghhZYK7E5CAHoLr7r5aYy2uRF0rHlinj
kIJC5gPiKKCbdMCUjsAVttynWBwfWJtesJ7MWUcYnITI9cXKRTFJKeEya/xztZH3
UwiRFBy1mJV/hyPeT2aexsBntefjzqErIWUQ7tmsfIFkpwg3uu6arPCI5rvmx2U0
suauL4xXME7fbFcJYcO3DmM50kvUXISKS2Z8JkdkVcGtePAAQmR+KJzJ9cEPfgV+
axlcmXC7tYbXC81ppKaDxUcwmmcsBj4DFXZh5hQYygk4Wdnj1BlSNt3iOqarvhaQ
AUnqbNX2u+O6yShi+NGvEdoUheOXbTLs1VK93sXgp7e2E3j7a56zF3wp/kvhfmo9
jdvBQxXnkN1VLP2ziWNJhudIhwjhNk7lSc8ia8mqBcirAcrN87e0WUvxkE/uQdwP
4P7Un7gQLgHWSh6M0Qi8py59EwzTowqmjx8f1JyqhfGVtm3ybKuiLb/448JJIikI
E/xjGS77gz3cFtuAj13uDk1fioidANucc+RtbomcBX0t50shO3gpZ+GUTJ13gSFA
Dm+1mMBwdkuX1YPcXE5oNo+SeqEKNGPHBRadZGe1LKyVKGlXRmjIFpkEskVrdKoZ
AhUFOGpUKii5Bc750NbP/guw6y0T9sDav9ni3YkrdGQNu+jKvm31E/Ngrjuum5Ap
3PC5Se09v8iIkJoh+xt8QP511tS+RGn6/UzJ3cLXgWpI0lbxuLU4BHkI2lkH6YWI
L4eNcdDXrkxo62QgB/Bl5ZIqNsONFn+syVIxNKkH7DJxoWuXV7UnJHAzCkLiAKAh
8bs9cS5SnKEQY/Tv5wjt4RKBZ/vXhMWKr6Les6Ex4C8IznxO00L9BKdpKSJkzOxE
Za1trnUZWYmAzaoXvrBDDYQ574WpnjxYfCDF7M6Rp7jbd9CFU9JyYW6+RG1aWrgm
pDNjI8Me2JbAYkZtY/elbeYeVti/k4NvvELhgd17JM+ut24OT/KJ1iOG8TH6rZhP
nbuVjQaB3ak7Z0VTkAjUcHu6SO3pckah9M1n5JuCh2IU+PDlnz6Qjjxkpv+KEd9/
5AXv6bwcdYB3g1R0qXJvdg43F6CQmu0vbB1AA/uhmUgjnxsmxAKCJke2URpuLx51
d5DmBSZtDCzJ1NvRM37ogipKAXRH3VHsbZn6yL4Yp3XYuSA9to2dcYUehK6VIwWR
2mIk6PMj3sAMJ8cJV5nwkcW03PBovP7Zil/wOXeRs9LoMLjmmpezavRJpYFaHYg3
Mbnr6zSXN1zJEe1u7KISnjiS4/wy27iCPuRrO6+A0uLd7DukSg+FRBpNiwf01fTi
fgMFrHc/iAO67C2w5DINxZVlquYE6kDT5Uw7xi+sZADtVQLVlMUPAUWFw5XaYSAq
Ss/CnhJOCGWbWFXjphtxjpLgbqarj/c7g9PdP1r+mrBhZc+UIi9lA4PDip6gPDx2
rmngHDoJUOcAmN6MCrAKzv2UT08JBEMVj+u2rM3vMXrT0VfYtD9zjoT1ny1D6M5v
oAxpHNW1Gm54gdYpgq9ymLj6DIiH7HN+ee7EpaxDaB0GRSbqkDd5FMJmuiU8Th57
+jPXvao86j6WueTs9Q7fssyZQa2dA4JsBm2iUyp/WcYmesSco3PG8+kU/ChINJFg
gUJXUut8p9Beb7HumFJwYzcayBjns6eLzC+XB/d8HZbKo1l1N0Uqui9fDNhPNype
roIiT7IYkfWNWsMxKIEPPRG1SgZoD1YsXnGdPrTpSbFeHcF2sLHTUPAajU2Vdhnt
RNA3lHbEDVj1sKG3p6hNAIw8qz1/wIBDj1hOE9Y7bbTV/jaj2ycQuIsvo66QsJ4l
WZKlMAjk6pfra6KYk+Xqm0DQ2NlM6ageud7FqmQee0vcGY/oWJMGnYEqoD/x/oX1
997lbydn+QrIa0WAq5NYgt7e9xc6sozUCIXr2BnvGgEM0lrTU0sApw2mGbTg/OZ9
xjP6t9w5+jqq07cDXxBsEkAiWz2vUUMhgK8dP6JR3XFcpigqOaCatYO4hJUdn/9B
BXVl1ghZvHBz+X27u/vzHpADv4+JKgMZS49bHUWhEZtK3j2Eokkvz53GhYtVdzep
+toM2D6k5Ketn1U6UbZKri0B64mYIQ3CZVu9jEh6dmUyil90b6QGuf8ZmpxudKrK
Y+F0zEko0oYHl5s+B9ZovMmVLNLtRWNXLUmjshPuZ2ssjhrRV+Yd4RNmtj0Gyf/h
3an2fKb1Tr7Pl1Hz0ajWHy4tRMPbgmYf1K7xNga3vGipKiqe8CZJUJEhQxKOqSN8
FhjS8vLEqQ5o6QJKnX1HEcNcp//B1BCobI5FNTcy6diGQL4XKCKNRILWKj5CB+ta
DGD1f6XsRs40zslpeo2i5QsdlRQ4h5NV1M6i2Zbd2umoTvryvLy4Es0hksejgmx6
yX3Hh37hl3BeGhmOlepLfx3xhtmL5gZCt2MaJjNslDs1oQVa+YDdBYidyOUOw8f9
QTdsuXX7XopGrunefm5gyVBfnbnjYbVWBTM1xsGmQiGWQil+P6+D74uR8Qsk0W7f
df2SjcHUv6g8Osfa19RAgoh3liTeb6sBqOc0gHrACGmwmH+QbRI1ugUb8a220XlK
vu/n9r3tbUJnY6+8i4qRcpGKf0KKKdcU8K4Oqb2rWmJ2foUd8l4RmD8Sy08fDXIX
SWQG1ZyIrP3hFails3eY89OMRDQIJNbG/EyNcRkr5AUPoZcwyvvZIgLtmNa+MJLa
BfT9/kbx4DMfjkShLyXXWFJKm4f5ekFIHFNiQHO0LESt7VOMA8o2WM5Qy1IElZDQ
0pE1Wc+8SWLKRDhgl8iNRzWQLwsh+XIx8Z/PLNpHqTpu/DeYJpn+nIMpoYrx974o
Gk31H6HHmPTl6cyWb17dcS6qUa+wICFQjST5XPLdd4/aUcFIQfvHFcf9Tla26M1l
iy83XdZzRbEifj9o1499YoLDwnIv/p1DLy1N/QL+Rg8OHlssC0ChP/KnpItV/41z
JREhgCKNBRqJU8XgiyWC3tBVeBz+176PFn1yFRp1aQoAQj3x0uyeD6smF1Gu/ulR
FLGWG8+MVbMLClzrGMGtFOpBMxMb+Tk9nr1bk9Ethk3v4ZVWfgFTbzYyB8pc+jwn
43qfV4GWRH3TjYhS/Dhkao41sXnLAb1MV3vgjFxeXQ4vg4LQZKBlOZjsDh6MUDn6
oxupaLDoBCbQCMVQkZln+nUDUusAdHOulUlzSaP1QPyDMehT3cWQdZwINw5LSesP
Y+aR+63P9/uYcBQeuoUXsJGYcSMabyWBn04vrS69MDdksXXNj8rDSQaJTpoI3Gv0
zeJrpSpAG/TfK+NUYFhqAeYX5cQV6xvNIkVqN6eRhYWDVKIHNlooym6mcWroenYu
56cDpDuwNsqT2EwEQWtVFy08r40dVrki/2H13034JxQCHgaiiJlUBtRx+vVzVKDn
43bu+ydhwJ4rBH1QUDrXDA9rISlFxXjO8zA5fT9wA/gnLySaJfDNExMV7gPqZ+yi
MFUvkVdSLnpa8dddKcfLjAqcbbS1DghfBafGhDUKLNJcyQl4kxS1rAPk3eVj/0Vl
xJZFgPLD+aI+yJ4VpyLzVwu5WmKyhL3fO/qLDSu3u1NdcQWJThgt8qImir2Ge4AK
UhSaDjjdNTaiSWp5m+BKp/Hwey/v0b6NvpGfQxHyB5tRegy2josvc6T7nNoL8V+d
oYqkVtLxTuNtFUk/gUfMCsYuDdQbuwVxFnggYAL63JIB19SLlneDk9DLbBBPejCF
fYe3GtYbeSSdloBMO/MNQNwJg+IDTmh23H3+yz0Fk5kdaDzCLLsF4NguSKtkm5GM
4/6zFU6aiem67YzlSWv+ljuoAzlDay/go+CHzfXwTHW61NVmeqbIpPfAhN1w98Wn
F/ASj0xzFiwlnoCIWiZ/cX8eN8g8u8DTrG/WaArs+wgt3joek0qpg5IHNoS+Y19T
4UeFBxYkDyns7upB5MU1cR+JXxyZwXZnQAxPaLNWXcsKLISxlcqP6kQHSj6Z+THd
2QYp50eB+gN1ZcLos3/wWqKXgDuCrzFp7c3hPHgx8yWygZ2Yq0HKMiptbWXNaifZ
gXdBNxmIILD4ckmg6Mrkb4jO24XMeuO+xwy8XhAm7Gu5rk0vMw6CL9kZe9gMsLBS
cETLt8kPI1UNBRqWL3+0B3IqT74TmJGI4jbD0VPRZn2msCSs5CjyPLjYaGQq43KD
PtrJ2w3t9VfZ5a4rXs4o8EK/qGaArJLlCSZI1PrduAYkVWyKjqdrKSCTOJpDJwuE
cECeJniXTAUtQE2f63AQ9HJXvcFeQo7RvKVl7LoG0f7Dr84TKPvpG0UVRTuwVwcr
TSdqELlaaorHdrvkFZZkJxLrTPaAuZ+tNxBGuHTM4WyRiShSrMXFtpQzRXdoLibl
zOp10HCZ24UbmAwsQBCC2ago0cyUh2feakiAcjehQshrQKzaU8zNt7YDk4NsT95g
wMgB7on/MTPIKeGYbodedEviIVAXHi7nVM0ag8kWBPDdShsUZNPyzWTFyGluTXIP
vYPTMmVKAy/7fUFL57FbRdL2ajnu3W4ifB+myJCaVqfcUxB4hzzF/wOAek9dtjlv
X7/FTVcsFHa2TzAEyhkBbTMuNUGXwy8u7QJ8fy9CUZyPy3Z4nTI/j13KFa3D9yWN
ZdQbppV6dIwFSgCxub5M4fL573bfRglfRPcP7fXr94Bixn3G18QyXmIedVmAbGxr
DQZmt3AhdyTOZaG92/2KSfmslVDUu7z1EC/1JMjWSt6ovXSA7D1o2v/nK0Cidcq1
SDJnjYAoZLrjt2Fx4Yg56K6cHKs26JesUY2bhUTVUnisnUk/CSU023CkSnq2t5/T
2oUpjdzXdJjvyXKxDss5vZlC9z3Vf4xtC9DMVZnLy60fiK7WiqJDV+EbX7dWjzGz
OaPBmERrYrYgQQdPheyOZu+wV14C+r47yrZ31SD3OHhd5KHuKgDRi8oDzShYkXX7
VPM6FQAw+cAql8U/IP4bw36gtCsNAb801wJjC43ghQp4aMaZAj+q4qa6JG1H50Qb
doQTplCEGl5beX6T3CtWD7r6726U8I7EtiaE7XtAAgjYDgNAmxL4XsgXDCnXXZOO
S39kvcw7dUhmKftZ6VFegmcga4Edvd7J40w8skEMg9xzO5kD1zkiqx6toTmOKpDi
nrY8XitZBwS9lppOgKAAlCllTt7nxaaVstrE/gh0HPmQ+z6PDHt315Kp0lhtQxYx
n1H02TOnmGMwG4iXS3xFK5uc+UVT+UBZ2u3R852gQGMYsfUhAE3Ow/zEn25GLrNm
8CCka6dKEonbcwI1av55Z2AG2xcETV2tol//+Fy+uUyPZZGJJBv770KxdBSIgp9B
f6XkvV2gUf3QWLqGoSHQ5o+3DLftIc3fOmqE6SSlFDfZGO702OryhqLTw0ee2trw
tGYKO5TR9E1N7Au4dC89kBq+lU8x6gLQnb/LoqUgyw6GHr6EeEAiUOtyZzc+i6M7
Nrkm+olCWZ9TcomaIDs6pyxPjpkMjmv1/pXu3mcWvZGS8hhfDo1eBCUw7wlh+mfJ
cWe+13smTkXlKKn6hqerRbFbzIDvuph2MqVJmVAJCq1FCBFuQ5YWfChUwX5Kp8Qy
NdAlpuk86W/oJ/DfWluyeoyakhgodIPDVAU32Ctb16woS0HjP0tE6o2wykUjFlg8
NKEvxqZlD8q3wfQwNFiodSfJiirLHumOuMnHQIZtRA/CYSDwvlxqVl68HpIV8TBY
yZ3512hy6vKMFaxbUKzR4glaGcc2lgJlH+4XWtyRSiIYONlQ6UIgwIYIMNtmKRoJ
yWLJL0AUR7wiy7RbhCwFxRFNFmp+ZeqLncj3rl7pB03j4wUIfelcOspEXKWrohZ/
Qa7ZAwGEWzAd5c76YHjKbPSPlgjMmQpKLm1vy2SVJZOZ55xmVmWAIRGey2jzwNAF
kjtcqeMt90TPthXEPNdkqRSvthp9lNjfAFNu87UwOYC/KpKUM2XGjBUoctvtD3kv
QPrV8hHxbXHv+HmDLrYRjhtM7Dr1jNyrDlm2MCekCs5HYy0wELSFL5R7EYfARUgz
ZNHz4gvLMl0M0qcJo/yXC5zluQY/SCKK00PqRIc23U5QBGMc77RR4X0gPqTUq1fW
WYx64va56OL1IQzSVv6db0TlQiLwEJEVhQNljX/ywFQLOrdGuWS0gDNhzuRmq82Y
qWSzM1KBNAGnJn2Y8AjYMy+hlA3FR3tHka+crrjgHsrjZmSjgC+9vjvlX1f8J4rN
ZZVidOT4lcb9M51ish81vaPdgwCIc43sFcWsUsRNbF2drDSeJIq9jRCD2oB6Aois
oVvgcyuLcV7YExsVxL+DZL60UB51E72XVcwqqoRR3mgg4tDoYx0iidZHrzh4RK2L
Um+yL4+ath08C/DANxbNv2c0qYf3mTTY9gvSWu7eZzzwpXeKiwY+PcIeV+BWK7bo
ofOJHn5HBiTZLLfnhdHHPhrn9bksQrBF57MixpFlqVhX2+8ngP7mSlTl4sWb0E5P
K/uMaTlADDTMFqNHAkUsLyqnDH6z4RlWUPXDI4ylShun5D3BCLvoykzPb+eMYXYQ
Tckg7czAcTZIU8grBtIqxz1Nx5be1ufeR4R+6AETe5y9ZI2e1Q25LEew9Dmp50bz
xIE8mVKT5CB2xoC3WQDgGxBFqmZP+2JXNeEEOS1uV+bsq09JAwffuo9oU5rXjuZ/
9Gh5nS5ckqAyCX6zjUaD9kjq4ftR5Adab/I8fuhrJIehYpMb4TkvPWaO4/edsikk
MUq1W45ngOH9VNcwjel3cZjQt6oJeS3vc08+9My/ekDMCRJBUKNVJcwiRjInViWk
h/z8y4UXYI8R6TWeYocNDwXh5In2gs6xRVV4F/e65ZtPDvzyDIwe7tMF/UhjsRN1
b5yQ6lY6Wwp4Uh7it0a1uZUYiEKRXWuxrmqDMNimoxE6R/hDEFDfcq+XuhbwtXIg
TKMbXI7v7U0S+pAY45vI+cAPBW312giBzc5hS9D4bgzqu6YvCb1Ccs2uAflfXFpx
JGjQKtC9fsOX3b3w01rLC3uYn2WBr/aRnYpnUmSdQCYueM90+hac3xE0TPI5BJ6C
OEPs9Eg+hxqvV1QNWDmB0yRmg+fBoAtyaQxU5aWs/wjfrNuGa1jmFUrUgIQ/SkEo
hCvdppUUL4QxuPgq/3fDT5pzD393mW1tmn0Qp/ZaCu8n0LH5ZtHKEGLapHkeC2av
kzIOLtHV0pIK1UeVBhF0RKlh+K+NISUlPeXgv1puplWkeeFChnLaczc1jv2dM0CG
BRDkqx8N9coXVu/i5wIwryWcH/HXhjZHTQ3AxCul1MpjS4zxnOFWNrnqLYRjS5aA
S1iaBgb0xfJCjMhUQSF2yTqiUbaFis1RvzRPMSTqz//5QuW+ReJmr03wkbkL4gxA
7VHKNsC6YkeBhHf6ULqkR086AgVvKfd8HKKRNxnEd/tupCNwCEdCs3rLoUz5Mh92
+vgywM762Q6dRqmwMo+Oa9R/ocjb9YSvkyU+/hV0twqi5Vb8CbduB3ysAcio4s82
qqzP0RNSqA173bHIZYvePQVJkxz9iKg41WY0YtyLnOXq/JjfXoWDTSTnxYHQleNJ
XKzSzL13OXymU/uhynF/25t9lVJmcC+cSLOm6B8YcaIIyyUnviY9siKLDvgc+UzI
5KjAzYM3UIwx54jiPhUNQQlY94oxpRT82bqOGPxDmnayPgr0Il9vGCAPt+ESxbSC
7aHHeljrxUpqfH5Z11JxYffrlbWA/DR/q8zMHGFb6NUkXGOwoY4OS84ZEGVn1lmO
d7nttX7J7bqu/ZME5hZtvG3qN4hC3EISrD/HAERzlahywIGbaEf6RhtJYDfOkZzz
6bkjTSgOTI5NouQbvQsUh0rXTgASopxfrHXg7GYXQqzT1n957vWbocK5NZ9QAkXs
/CQqckPGxAa1kLfRLQRrZF7KMMXNvC6Cv2taxrGnRv4wGRv9eOhZksI6kIbgfVqA
of+yT8jsyLV2iBS9ct/ttTcQhtA1DsMUw/2rdeS0dd6ZxRvkB7AZbCMGLVNOuZEH
HVHaL47tz2NZ/Cl8T63IJdCY5umGgtqT3UuV+fZS1yKabcC3ypiOEV7TFOEhetiL
0ss272wumw4f0rvAOK6I7UOelGMMkzH3cXN92fkwB4K4V1PMPEOfKvOVFtbWrj8b
743O0P9sq8Glgd2OsFHvPp2CjIBxy80qoiMavb9jitjfrNn4koQVYEkV9CBeJIGB
htR5xRWjenOsZBn19c/HYPVhwRMyYRD5r20GsjZtHup2n87um4ZyCr5PNawVMxkk
bRb1K7hGI4kvGCC9y2Q4hQhOWmKcv9juQyFmpikI0ycG9eZ/OKH9XEOqktiNMLSW
/LvPmAH6gO9pjt3dAd9VqhealKgkJ57pG7hje7CVwZMm89kz3hbCRRLl5mnmbZdQ
TQqDA65y4sfUtz3Rlqs7VvF4NsEeIoAaKdm8F4vHWcl3IlnAMvzSBTz1AXqdG1jL
eLK9qMcRQfcZIodQDJuDyXmlC9TJDJzxsaiIHzADJgh7lHJIj2FMmy7lNhykiWPb
oM8/EdtluYmmVqtMjUrswLBOx59+t+DbpKpai6OrhGfIm8IqcHy2MZmAQhdVESZw
7CcnntN80z22mGLpCCvXG4C9l/jKvkccbr7OHo9hfdfnGq4IRQjwP/WfNmC3RXI9
QM8/ADdoHwkRJwiigGKXm8EMaHgnoQaZEHQLdraLmCfbQslArJhTlSAJI3XJnv9G
qeLANzk2PqyndhXRI0V0hDYaOQuIHsyO+GX4rgvNdvMlcgWuFZ85izuXP/xmYDyn
D7hUrHK8DCHc47/wr9IWiV02j1PFKbP30bM91R2NKnr2+G/lgu7f7LWNtI64gmVM
OTkimTSv5BBSB5XLKB9TwP1q4zJa9ID5A/JVms15hWH1wElvmiybO0Al1EASgmhV
1sNaAfu+h8dkYS1kOhX9Yz4UJgHgnwsaGk36srkn+lP1qbSoM/RjEPt7ldxKziJE
QB53o8wJ4TOM4yhPG8oJSij6lPqmtMSW8TSXKS8JjW0tJgaNrzISeto+ICkPlQ2J
vfo5Kt/mLa+N7/NmjhJm8JG9jyIXzxyyF7qgJr+pdQIf4xbi0yemIMu5xONaIAZb
J58j5MpdJ3X6i7q1gLGpZbrhF1Uvn0E9dUp0BJKhh1ejsFdD2qtXiCP6AcEInY2u
wDuxJzuaE6uOYrAWAueEnMnpUIps0HiY+csg81FCQmZ4ck2Xh9Tv58nF1NIntLDR
PpIwunXZJ6eBjwNrcT8OclCYA5FCqM/DSpp+sqo1jImuM0XGQZfli6e/5SW/xWwz
N/J/5BXntWcdoTV4hHJ3aWeJTVcIICG0/UUxt79/SxWkMrBigzVyPbP6I54SUT+j
4+jQA4gbtxAVL4TPaZDiyptqFpmvRj9I9LhYpkcARhePzULRQHEAOE6/7UB3ygRt
MeNZQ1Zh91rDysHAdMDnXZ4zl8pWbyup5+PP1Mz7zckGIk3wkNG8HHc0qRKZ9Ktq
W1XESjRzEs6ZlSAR+uAuPuo5COli02n7wafzKc+VB4n5H3jHD3y+UUf8LWAvMrg7
XvmZ8RYbiJcamYvtfnyULM87FPlPitaa7hfDYhocVat+Ck46KY5JNVfwn4YW13J3
uWSJ+I9Kqy63uEM/4cFLr9wbhcKSDVOudsDpinkfitFH+C6YTr7Z97U09AB4CzaC
VrRpHOWPmlfUni+J5Icj374TRhQansTDdgfEQwg+4en0s2HE49AMK3dGznHUrNwW
g0D9XwIdlMDSKHxasnfXszlN/Hm9qVi9t5Jofg+As/2MLAxMg1a2lTq1YlT1ErAc
c9Etn2Ek6g8+7T4y1lBkTrirTDgkKlQv4C3Wp2V253jIzfUTtB524Tun+bIMvFpI
5/aOufnUmQAg7X6kcQa8U1vTKGKKqohuaXUHECRRkPyKqqf7p72OMbboHYSbgSfl
w8qs2+V0mz9xmZcSoIAzHh5HE7Z2PTjF04U55jL/ucBl8Gc/mEi+ABAUmq6LcDl5
1vNMonYTA+8/Wo21BuLuUfMrSryo2P853Dza5DscTcseN19dUnGhlMyagAHdaRM6
SE4qxgzFjRV7qp3f1FUuuGezZmYiJjeP6nHxQGq7Iev4f745KTOXbO+v2GprJvSl
Hc3Je88dLiezJLPlVyJnkgkTTBE49TDUWTd2FZ1d9CtPoEiTPM3sunU18JFW8asp
Jk7dchbGrFTIJKY3C7AV/Fmxu3Q5Tbbf0THwQG4G69+sx3zhLOqTbOi+UC0Hnz89
NASMkfqfcyEKIN1O8rgUgh3RwRvu/ii7WnASioa7C3VjRhsdpnET2b3f3k8tZnXx
p4smisv9pPl4Kqb75Oa7JB8oL+ubG/TJv82khkqJBJFDrb3lsGOkvnvTF/kW0VOE
EnL/uJT1W/ILTvXYpRSfdmv16GMZFDkA36lAhVNIuM2wPm9AFP7aMM+ePfshKisK
28K1bJPlhWYLw/Np+zbs0usMBByfU93O2J1DtwQejwINTUVE+I5axplNvAOYWkEE
6WImw+C9hfAoZ+f7hypy6n5ulpcsflk4zJ2SwP+rQc/DI9Bpv7sM/4yZTCYY9ZdF
y9hlCDJQxg7sSEB9+ieeOPHgNjBFUiPoJPsOiQS1Nq49+AKPdq+vAQ57l9RXWtJ3
UHQHesMjVxSlHa+mKlWQ+jEym84KtHbF0JhI60LnfkAPzj9zMvYkNYjd7iOdxyo5
zOoC69mgUY/fI83wAi4t6ftRqYgmMGsQElnkMmkWFT3Mbls1JXGMKlfpg5HUMkJI
veE6/628o4Pli/oFEo6kbfA757FeR0YirHrNkUZFWo5s76wVoRZ9Ol8jjN4r0Xyh
zcKU70EvR910y93YKrFbu/lHrYHkDMT+Nl8yhWYp/ldvso3WqzKQPvyoKQRS7cIF
iev0h1hshEvUItNH47kqK05E8IcN1+Dwgp4Ti7vtWqqQ7rSfhR4OZ+g4WuRosyHP
WJ1ln7SLCu+jg3NHULTEWWrGQA7nloBC2Z8pHfHfXu220fBEEIBJ1PmZOJFflzXW
ZKaWXSgxermNSQjzUwo8334T+h3h4juL4rzhSBxbi2Wiv1YCiW3dAo1IrNbrmBTU
wKwSnFhR7xymto0JgcvkWho0Rv1OfJ2DUw2PNbyUzvfHfJpI9zG2lJ/21Wq6XD6k
DMrjqC1rbWdKnBw7wzv0M2Yzy8gujgZlByiHJae911H0P23oi89HHmSsCdtAAmHc
izZypfnIB07PpdkT3mSeqXLhHW6b4anB/Fz+ANsuEcACAlynnA1/a5QayyB5wdT8
+vLdIkE3eOCfQfksbfbEmJ9YWdmyoRhplGjighmXszl/ZdcH+PEICIG7zhP5O6nX
4NkDpv1Sjpw+UA8krQfGFBteM+l/DVjCEIgH0LWRRRsTGsvG1Y2wCb1pcRxYwH22
QghSW7vPu11JfypvXrxxVr/SLghMMZ/TTJ/q8ZjmU1n8ymUreXf1cuUdrGBMm3Ee
jnNZ8yO4sYgj8zjs75Ta9byBTkNFnDYGZWLeMU1Il431Mbw2DOcpFZdeJWnVX87H
B3Guk9Apb8hBgZljSVpY5Xciu+RZ4OwWEC5jSSyZoeFR1E7rKp+Pietp6zbpiuiK
LDkhuP9NCcJH5RF1uIl8DxeaiV3Hju5gt+sTWK00hu4RUBf6qIlR9EcHX/bt4odn
9iLdoBgAc5ktIqn6T6vGHdkKf5Lf6MLNKPJvsE4Sf7XmboSXa1qTHyId0wC3yO2+
kIKP/F9zn/Hioj+h8/foiCnJEMk+llQJNKxUW3rG+/PUKjBeGm4DHncvYlZP0+EB
qUtivb7JYm6RsuKU6LpYYIDN1ADER/kp9dsYHdo8klmiGn+C7QF86w9Con1BfPd9
SRyVxStHXPzOJ8JKIwXfxpWud5AEw0qnMlTikGT7oA45Ip22N8WcRY8OmmwN8XSp
5Vb8q+NB+Lnwl8fga4P2WYtRNCv9g+/VG54meeESQ8SqnrLF/lVHWAHKkT/lYjfN
F3O8dH4x3l/P864MXg2ZH1hkxLVKRvpyo+o7luXu0XBDVH/ArIdXF9dNjK0wGUzL
sD3O7QgZVbduKhuB3YAu9YX3koNChKuPi0oU1XaXtK/A1K0MRnzHxvASuNdrfI7S
WxwFx+vDCZcQiStaAtLI0QLSFze+MpAadvNTncma0+Pat8FfBbt5gIoT5bBXww/g
8XGsa5vaYNXIQ0E3c/+WvpuS4HJR6XHkkY/6pjJ+AzdWJb7vQa20wMnkIRusPrpv
gTlILMkIyL13jJTT0zMBJEBxDGY87qnT6VH4aK29E1IPpPt1op2fo/M6aLNXyVh5
eKp/DVpVVjggwiAYNDDzR9apPWavKvwrLm0y+7TFgYxgqcxX+ACr5bRBXrnCigQC
Wn4Ie0PvplV7zXrHIo7iUjkc4DO9esScdE84TO/10vxhse6HBYA1lOp2OKm/urzo
RRM8vTk3muN9oKs9WTZRqk+ONgrXLDrv99tw5ApRvj/Eq247THW8Sy800aFrmgbu
KlFCph5PhgJJidD2jbxbkJyJPilmyqINP61FedLCbxu5MI5EUqHXdkNRjrYlItT6
Kbksi+ypu9w2ELtd3nohjDHyyjJwbBFaTfm7NCyHI3fGDA+y7HJQk2M+gwA/8zyG
LYF2d3IpLh5Uvo+xbgUvI28tBiKf1MI1oPzKi91pxevFhb+OIKjBFqJM7nF4qDHL
G2r+pXita3mYLyT+cjAKeKp8S35xECxIiHrXgEo8y7lGUqQ6AGkgP/Fcq4PjBBrs
a9iK4PaDCI3RiLzMM6cz/4mDN4I8TIqOCRG9H4n2PSMkMusyQ/jjkXMkPppKj+u2
InFtIbIorS25KxFdo/3RHnEcciOsdh04VWcjH53vmDn6a41fRGaAr5/vWQUrSK4D
xFERcgvSuLV94VaSVdCsdlVbFBPWoOAVTAkkhpvMOUDudZ5yW+KbpOlMrUlMRkkX
Crf1aQYXoM9xjUkB70HTsY7618ebeXNXxijC6aTl2IUCgRpJZ1aaUYZHk0ZQNRjJ
bIHfjQbBGa53LjK+IedDa9EUG9d9uayGYm3jfS/QM4Dj3kbX1nkLuoOb9CoFu2Jv
wNtJCyJq4k6J8iR9JPdo77jwL1Fz1oqC0j7CqbSszHAFFQ+hhiNg728jDhazKi4U
Vl/i/GYP0NaPWCVDBk541YNpOJMefe0D6sktofWDaJNG1sXZD0eAc4JU59LOewFO
gA4M4Df4KzrIpq3O26Um161yWSsf4ZDd7fOlaQ7ZU+qYj2MBshpFoLtpX5oaJ78O
7Zq1UJxZa4c0k2fWJdZivoI7mwbIfob3oMY70O7UI+T1A7I2XJ+V20lhzAOFEJ69
ZagKf3xw14FDLPAdLp97Sp2WiPEvqIOr1WcrM2sX0oVBFBYhkbVfK/lWvEidBwbR
VQVl6s4w2VzJSN95ynVeRmenxBc0dAnbn7QuUSDl9wL35tuUc9bVPPKz4ZNko7yt
zXEck54hhfz5yjTlWx325ClqHgzQ/3p48ffpo2X+viG540Zkv8sTquTWTtlwTPDF
rEcAqqhpNn0D0To6PtSNkL+7abM//W8z89AqJPSalyV8jYzwsiAKLH9BONkkXviF
Q8/xoPLBIJNiHuty81IDDWnckrZeVKugiTDOJC/9+1fvHBWgFzsZnTOobvUVPQCz
9OlLMoVvO4qRcRk+4vCM3SzQIueSqUtoYlcUoVgc4jSS0vyW7TCq8T/nmqQENMNX
tkKlE1ophlHHqmjlOrBfIhjdWU47DI3czZZXcp3rScQn8ZHW/Putr9M9b8TqFpda
aClk/PoxhojlRZC/xeBkq8im9b4yhFOV3wItnz1VPfBp0CkFKcvVsuuDRRUUJ0c9
XUtriOoFuWNFU73VFtDn3rmkjxGRZfXB4PeK4pdfN5w1m0Z6IzI5aJMSpm7JLwZS
8ECAr9/xUc32+yTP8WNLT7JnEjvpQSWpQmLwxS1Mbln6Kc0bE4Xrxbhy0XwhrGE1
fX8feg0uBWR22zbowxnRfuoBaEKdb1OD41ZwOWKF976Hy5lHiI1kGWMB/mHsEhuS
/3XJh3N/aC9HsmFqFw0Swr3zqIaD6QCRqRUZkRYHp7Yl6jZNHwHOWL1m3Dg2pv2Q
OwvP6oeEPvAnMOM+JLcOguIGHto804uXmXCxBN2ntM5d10YymSRtVycR3DT5/VA9
GNQGcHNlMrzRBKgg84p4piriHoKmbdwBH+/sIDQUe6ViO0egJPygqq6mX+HHOqqf
Uru+z0WM8JHHUTmqqrNfoamtlP2qgSlHMqiwVGTPQh64bNWW1fg4TVXsnGPULm5K
E0cCVXoycedZFjp4gR7BDwI1p/FuYZO++dVDsXp/aNHawNGysBK8hO/GehNytO4C
W5/lry0XJV7bB8XagqqTe7igVE/jwIKIIWIUfgnl+BEuZj8bqw2a7LXZq06Wrx/k
d0heEt3ImiJy0IJoXD6LWvs93ONQu+BgIVapcjFtYKE2b3yqtfmXPjG6MdKOdBSy
eBGyzXYJYBlEqSycpLm1FOmcC31q2VqkVZhuVgq3kh5mOwlBA5TAujnoCmRybm0S
3PGimAGkYYkYVK5ga6liWJqzQi68yJ1jRMC7fwIb7W2FSlWIo176kAmphANw5vDD
BJet1p+D1+mVFzxqPJ3C73kzb+9RgG0yyJLnsNxDh/v5/RZbCOZwzvvzn8is2wbx
9VRg5YLQn2yTZR/U5B5Ky/cE5jHPQYS8GxqVY+T4YVRDM/vFk8oW8uI3m8PIWgbX
4KqdavbaJcwVdf5GLu2/es+SPXnA5xL4KRa5r7pVmhb5pND99WZVoY5JVIPxCXhO
h5FVvBgTAE8E9lV1nAI41ognv5x0zF6nlPEbZYzxfKUc3vN6qdpsvgAVjNgqaftX
CNNIkSLDJ8rbzz74zRAtCJtjg95YL31P37/tt5OCSfrc6+e9ClltZy/OGgYBrNg5
1oThFsw/zrnwxF4JiQiKSGJNcC5+Lxjvn3603Tz8/10S0/TXQfXdABVfYDXzavR/
JwDriQpQN8VrwtnDLKlUGFXeNmQyH0pHNRVGr2FCnaSar1O2QKY/H3xE68LnB96S
byxdH1SW24l1pJTndABsD9o+AD2yReyyOICPs0rg639ih6dlS0ECeCl8hg8bAxNQ
ATieR19Ay3Pl04wxT1CKmrhSZ4kW6YL3ZuFOjFpJVrsgHlIcBPMYv/yvlpNICRXY
tfBwf0hQ/GSSuw2kJG5TRyDnRThNAqn5CxeTMw/Di9snk9n+qsg1j959MHFal0g7
m2CX/UVnw59dpfnYPqhn1+aXyenQmEyF6OBnkomrZa4lvYjHEndGyGDNsLV6KwD5
scXvJ6P3/uXDYXeCTPcnmwTjL3Vypg5/Ym5NJ8KdrsMC77wFyX+yhlbPjKwUBP+F
9DbulAJ2g7m8rLKNGCb6iNweZX18Gj4n5qEbAdhk02+X7/8kZMTQPeDOVoXDRCb5
HOh2Mxf815fyeOYOPYfHlz7L/5xkYPMJiEMN0sWQF2mYuO4NOey3XwZdI4XILM4c
mMyJnIzJ10K6kqrfebcVaqcgPEMqa8tl0+diH0rDQqjLiLfRzdmMTkoa7CHunwu4
x2OO1EnFuurTW/VZsmF1t6w94YFu2GsVbw+sP48fIPAZxeuZbK45p/v6zsSUTYGB
enNGs79pN7od/qFAGqUbxF0leyTX2gJd4H/ayFpt530+Iwt/+0riRD7iX4AB0QNS
+6Vu0Wwemmieq0CjmkcEum6KYlZ1cwS01fSGggW0/6X5T05sKXvhD2ny4X2FJGWN
XLRraN10Hx1lvww6ao3pHysBbjJC6dFWX1DYQf1vi4pknAk4QH1XMHpglL27FZ5n
XR3KJq8rYqWh3zEQYDw5ICwH9rqUoL1QgRtqtOn3yUcVauGzt3y9qUXOWd7FF+Xd
EBU1WQ30JhXg3GGCF+hmZOkFebFuEp054AGIScpgCpPSmiYJueHTtWlsgLj9jSY2
n8zOenyb9AC7SyS/BLnyqW/Xt1I/XrAAtEZVY9hZ4x5kfCimu+oissHLcpeSw4V/
0I/FWpabBM6AFt12UXFj2cBTextvtd3sadVTTdzBhjqHBnVsg6WAVHab5UMtwQPy
38KhdG7xBhUuKdpFmk93H6JHFw2jvV+Uyxup6ErIpPwpd6BCC//4PZzHtoAF02f4
5f0Wt2sbOiRVuX5BBrYv16Ujvl5H8+YZYZjq47SnS/JOBRrwT147lQqpkoh1oJL9
BUIdRcL+dGbavwuRmI7Kf7RyavzuQotDU7QHrHa1S+b5A1Ppo7Q4SIXd67ien2v5
3H3n9C3dSfs00N02hiZz6vg4LSxM0HalPJ6vfvAFdFbVKWvEjpBDiomgoSLexjsj
YeQSP/FROrWU1pSrO5HuwknhgZ3d8h8dy492xgvQ+DsaeHoowyDgZMO6gmxw/c7F
BgikvlqnooFrVqPadygT/QxZvUNHNTnAnDhvUj5UfBiRgTX40F0Qt8CS8KW/hifd
7PQtsMdnIZPuYgCY0G9HxD8srL591DrNkASJybLwvGnJeh4Bh5xFVTP9LwhkQFJA
4xStLujBd09nZxUr55zmeoyOCR8IpHx0vdUUkuS02RdMhOJ0/tT7hQngGp1Pkq6T
JL2XwHgDr0Vc0/XVGxN7IlOXCxuHUbBs1lz7XaqadGuSWX2MB1/g90pD62bvNdOV
sG3PTHFJmxl/qtH0jaalGevpfDgFOkseFU9RDiNgoEuDUP96TfQae2n7jyRkeKYR
gd5f8xPXyRF8f7Bgt16qrFqhZothRxa+FJjNUcIhsS152MTbhjoLCdIOTsLmtSqv
oWuW/Evji8jEZfUUxuLE/D0lYAvNPXthOeyfzrfAc0YvJ11qzut8emdRlx5UeW4R
CZxeA5FvfVf1+FZ8RyGejrt+OQfeC8HTVfWS0IQsAhzS3eGLhC56AVEU6DEsdW+L
CCOuIix5QXsrZfsCAlgEgeEaE9sgcdZWXJhnnR2/XlflbzQH7OYu9BWZAHpTsyFw
2Pw20a9/6SCrhTO3OIxgpOahKBHVZVdJswl3PE5nEzEfvqlzxVJQDHp4J9g3q5Ry
5dHKRnWZcFUc0kMJ+84FH/bKYqyYKM8BJz55NGZXenL+2zqet9QF7icx5HJYHvhG
DjhgexMPnhtwZs5KokqYzElzmL5uk5DtgD0UNAVZ/FKST4mWSisbL4kWUS7E18PP
uUJKF7VHh+HUkrrjFqnMh+3HTtnj3WCLWg1TD8zAoTZILiDxBm8N8ijw6TpsayrX
0RpxiL0rahXsyGlYU1DJbFD2Shskkh3kVerLJicSb0LtqkluW4tJaA32tEOugm/t
tRQmLNaAu8K3Nm9JllfUqrLYCefQl3oG4vRxE3wuengGCI0hFbc7LjWrBuLWEbhd
U4DzfpgQuXAVYGhkWK0WWF60prfI69HzH9v16eIZQ/5L1Kd0tBOVr5W7bIYRWZte
lU/9uNbVKBWspJ39c01Gmk4e7TqzPM0P/EqFxAU0/XyIpnKC5KABx+Z/78pokUa8
hNlOPUvOlIH77/AMSQb8iP0PE8XX6F4H0//Df1WkaG3pIpTPGi9IcDzGP7dH259u
lroxTqCotzMbJ/82RONpHupCJYJSzy3OBiTndGKQnSRPBW17k5FQy5da8FqQAPJe
pfWUMko7bVmbPFdc+SFPhKQshTp/oP9Trbpdhfdt6J+AaxFI1bzz6VuQA1Z020gT
+TAdCNE8sVtV70IrsLh//Kk6o75S07n8S5/KeJZWMK19vCcUNV/nxeMyM7HlgRAy
f40yMidu8pGAwBaSOR9OpesuRZvfyG4WSnAxzELFub1ATny0zprUZGDnHSVRNg9B
fgOXqF24LnqQ5tdTPyEKK2YGeK5eAXFlnJv7giZcNmpzZGOAUQZuEJUt4iqcfrqu
alKgONnbuK1ecUJ4Rs+Re06Q0gvg355qAFno6OquuVp4PYxef4la2rPJ1GbOAJ1b
/zgQKmIkstiO5OWR9bcWh5s0kMtthYtGnhApxUP/kTTMqMCulF++47k3DMz3K5nb
dw7XX1nQz1k7PRkcVffSl3K6UCFy3qkBPgKPvtiQMf66Nd3syfRVmtz0oDyEeUzM
WYJDmqlwh+qU8GZSfkgPSJU6Iv7Ez1lHr2iWqkBWgeK5bnvy8Sdh2rOITkdk7XTX
fgFOpcy75suyaQXV44LrBusOrQJ93FtKRjm3v38WSmvkZGSbvHD5o+O8SfrjmbaR
lHe32HcApZN42gmXNBONSDZaEAZGfU5lz3QVjMEpr/GhkHvb+ze55Bna+VvaCli8
g9aqEW/hegzpUUjmOpr8aEFLbj29qSJU+doBYnxzHQVk7QBZ5P1eVZiniPqwgBqx
ErV/62CWBNYMbXleyxjlqc3qn5NAjWWVuhssmVqIV6rORe83lAd/zPwsW6br38I+
TJlSQKEU0KToxcFlwo2ir8QnS/kV8M2uczJjfnDnxDd3Wp/labEY1sV3xmfUrSEd
Yva8z5gjvOwCguxSssodM2aTNL8MoVXYVZGVjoz8m6GldiuJVeZ6Tfkg+IgcgErn
Ou90T/Y629HN08R4Nk7I9E98n2CK0K3b4y6fmD03E6pcAra2TUp7MqT8A6RCP0NN
OKO6Uv6rLyEANM0Qp/jHwq73nBg0L5KXMJEhFJL4bippGydPIiu/Lm0Y3FL45MlC
odHk3wakorHvw5F15axkKNaCSXpfR21fNuV4aJH1QaJHykgds0Q1YbLipyo6tI75
xwDStbsztJO4AK07XG3uLAetGfOPQJMwuTlP2UYZKqEeXvFqNcph+1R1BFKJsQKv
S/2Tc4VAeHWHuBhosuXQW+54sySv1mdIdH89HshJN8svmnI+JXSyoxlcW9/xitfR
pzFW3cBNxpsWbhN+x2n425y+jkxgBCyMT2WCmPJmV/tCQCt9t0H5NBY9M7FTue9n
n6n7jK1g4AhCWCGpmwn8vd8tLJzTsKmQniLCReXmXFYgtwD70yQXxLlw2JZzqP+w
xE7w3fB5AGQNdHMZUi0GVHfVkYEsyD6wHhuWjWnQhoR3yUvV4dXub3jVKrsur8aO
n4Z60e8K43INi6aIPXlJCD93pBlT6S6C1qHM1xpdcws+S5xI8KJaSLAn8FIPhg9I
WP/m5yY5QBz8qtuieBCBQYnGjOv8cxAKUweA8UKc4pq+60VCwCow+Kbs8yKtbSCM
7AyHQdRksjczn17G9R00F9tmNv10d3K35V9Xhvz+bkBmTsEDU5RfcaQuWlvLt5uC
Sr8Da1louD8SA8LXhrHiwYfvXPgMNL59eYYThJizObaw6QshqaWLRlub2Ydk474i
01soZvJ57gag8DTJ/kay46u8F1vPxodDvzUb83cXnKVCPUTyfY5RPh/aO9hoaeK6
4i3Tla/nZ3uKg8OdT11voAcEb+nlCgULH7z2jXh3JdJ6T9KzCS/H+zb/Qm8uvLXz
ERjhQ9RzL1ctOZPj4zMoPm14KGaZto/8lQVcBnpEmumyKbr+nqQpZK9cT/+y62XE
qPJViZiKLNJaqh0Nkex0sP1GU8SZ9xiIt3NbNUgERBTwSsEU28huBC6VwTccocEl
Ha0IVbkF83LVMZwpuI3CMu8NGyXi548rq48oH9bazHIKvoDR3ohjReSJGzasa+QN
P6/cZ/4IUdQj90fcqY3SyEGwfimCo3ylzsMNFCG0yHtK16JYwUJ49QawZ41dByt+
IukZqboGAXLdWyVGGrFcExNNTcv7CqxSLKX5n1ihv1V81NJjksWbeE+uBPR+1KL+
GiN5haYDAzCI5yFODGp0w3EtiWb5h3jdXCXDiBLWEZBUBT7thWTJxF0yd/Ol9y63
spNKpQ3xKwGKZ2c9jxl9xC276ADHVj9WX2Q5RF3vsm/khmV5H3Y5XloYc3hLgmcX
Imxdq4avNR3I5poklA3h47pbJZn+0y1Ge3Ha1JKve7Pp/1ooU7qAzUhw1whfsmUA
cHRAt2pvFaI1QUG4FZ2HAKuhK09AWMYXXU/7fzHqnS3LHmemcwKJU0FILt7GzXE9
zTu0E6Fw5xc0fTrs952KWTWaB1/uno3GHNtN2C/SpDtvEM1sRoH/ywwn/uOrB1VU
XBdN5+CLCjzJcC3UC/zrflNATH4EF870aYYW2PtASmaSV2joYN1caR/vLvXCgfZN
3ugt2o9mo4IPxasHvrzO+5aJNCVJc+/tgJCGjgBoKnYbpmWh5jIDxgBnI7bn9Zej
gXRlcOL9EHPn6W5dYrKvg7m6lUnSdsAMLpcoVzlA3Z1G3fAONmsM+tJH/RajCiBg
v0ARd7dmGPV90LOvEwe8JkSUy0lF0gksnfbGQKeH1EzPXTjbuzqmuYBGjvIiG1dq
ASbYX5MGY9G/lTKd77pSDzJwvNHGPudYvWBgRpamK8znsGKIDkX4BEaLU5EsYpLe
2tpErF4lalQF5NXTdL4uBupiVZ5j9H4M9ele4xOEe+g5gAj9GeZixKjRLc/jJjDm
4YDdMKFXkZgNUNyHFmP3WMufk5Ve6UXOI7+XVCZeN7GJbhvvyyGssj9Z0I6GbSid
sXYjlO+0x0sshDGrFrvb2iG3Z9HN1dcKVrVG6N1VcZNirz4SlmXVNQKDC0PKhHw3
N0uDQ10dZbdsYun4eLZ23FRap1DPDZwlk+yXfvPIx8yQkbIivOFT8wH2RWmidqOf
pF4WIhav7GsHz/xT4gfsNQ8XZougg/33XujH1ayuko6oNIQdMLPs6ZgfmD/JClFg
/ZN0HRCguZpIxJIdK4bpztrqSRcIs7JIld6POQrhmCv8YN0ojGD0F5I6qRM0zX/B
ofuxItnB4ib5MOwPMfG8QdcWN3Sg1OPh6UE2qOKTzuZtxomEFZcd4wU2pZK2ou8k
jLL9yt2UWr6CnlFJmaSQAiLai382jYYXputsX3XabYDv853ceLaFdeAuZIbuPZ80
9nkMKK1KvRycvr0GoGu485umAYhVHsSWEgKfyAaSUNSvet3oph2cKthHeyREA+Ue
9bqfGocOEBnpyb17dBaTAjqs/z4wzaRmH0VcCzqF/6spg1PiNEKcWp9y88WVtPdp
hY67a9Uc2UsavIAAPFdlQlkWTzCY4IjZ2R/8/1GkWcbia0jv9AwuXrMQLuc/g6Do
dNARLThv4eqaxRPqtf1vY6gnIqwazl0S5Aw63IWeMShGpx4nw2xxAJwrLjc2LcOd
mOZWO2K3isdsqJflwkDzGjSTD/2Oc1FK1/1Rb3nDGfxYAvHBFp6j/n4evlqApIV8
/1/PTdRB5+NmLgyF8dFmBskfgRBSW86C1XqzvHr2rsrWHBaZbuol/PV6PjDqro4T
Y0DBv9R6K2d1ztYPQl90lSUTo0XWk7M07eMIfa97PRODN99CwvUOO1no1ryqFAri
9/Y1VNSJYGJ3FXdZQbfxUywIi8gNwaM0m8VeLBqsTl1M9i2Ax19u5gFrFM2sQV4s
jrU70unIvIdVhuIpboeRKAu9Xpt28o5Msow2/u8Fyim1ipHyP9wJh9TgijqW2B2u
0eW99Nt2A8c4MH1muhgYFH13isYLhUNepQLUdLyLXLuMt7mcnvFw1bj8cYfcUd/V
YC3WhQU5rzYEpEbLiSk+/Yp2pSbIdQKnCQKKSsICJZyy7NoA2eiCxZ9KBRxTeRmP
sAJXVBFQFK2RfSp7sbBKW7FZuX3FeAFFdisEZJyIfwo28/RkIsM4ZJnwvV6f8dvu
S3IRwUnli4HA0T02NNx8gCo1CWJM/0kUTDPV6mzw+padvZ2T70CuirZRAOzEo2rd
TOA8hYb0j4x3SiVToYc2LnscOba2Az7+wAX2Nraf3OeX0cGomaColCWEwudhwgSg
PvySp+dh8wNT5auuhVKZyN0E7AZxbo0lhDUfB2wmyElhyHzJuEOFVSAo6pnm6QL9
b0PBturKAkMaIsNLilSUM3rgkxgfHUIItVby9df7lxUlSfAiHJzd/MGVasarYPj0
Ecc/Ad+GxTROUh1W/C1RwbPRr30aQrAfYeklWoMiBnviAxDnPgStoJLW4KkDvTxI
khRr/Hp6UAzTo78BIWBMpBfcmsuXxWoVgLZI5Lt9AJ1yNMS3PMJiHJOKDWgdxWrL
P0AeaADKHzxg4KVHJ9WNzv9xhaD1//wmwmGB85rH6jSxBB0Mq1veQ0B66G155RG7
lZc+6ymAxEjOEr0y7DZFlI1EB4K6iZC/QqgGG8oMYJw4QlTOpPn2ky3PcA3G+xTx
zBwh+RQheR+sDnGtDGUtpe9tzQM98wz38TCQYCknLs/+XXzLqvvk89SBRV9k2mlY
rLTONCugZEu7+Phnm6JGSPhijipxjjbJrxZt/S/TfRGrfQgdMUki4Wq2I0GVCjiY
B9gSio4WL7Gj7XQOFAevAmdLl4WfVU2kVsYGA5lMy08tLtylzktnwoMTYWUrFLgk
sFkxDUxQkkQIpSzKn+IVJpDBdeLA68lODC92YEUa3haLRb0xxVorOkQ0D/1FUUE4
gP/kPd+1ZBz6kthKvS+Vrmub69emsTmV7E6xORNL4r4ZzuyqpVAh8C7FFoA1vuiG
2EZvxls8ekR46zdARjhzyueBL7cjlLgf1Xufjz/w1lfqxjFLK42v7J60wOrHY1Bo
NZyrUdpELCrdSz9aji4hLfg+VuiuCHn7IGaN7O7GBhvHhgp6i9PaEb2UfJw1SWZ0
/xRU7ItrDifgMh6lsspJLpmWLLtwGWrq7FE+dQrvQTqKihNavp1+6U1lfMv2tcZf
sZr7T2a3vjtZz8DfHy+guEVGAgsME2yWRO/d5WwZT0eU2I4ASbHSDjLy+8Z+DNjB
Gh3KfJ0UpVfXzfa5aRENUyJwg+1E+MvocOWX5YOmWbQipqLyTp91/wovIbVXmHCV
ST2FjZ0WoMvlUcr2yVKybdK3vIHnDl41m2mimFhlSvj+9yh1vWHn+KqnecewQN/l
AbSO4IrhoFqft0GNVnlFj0T8+q1ww/h0S8C+uueYKq6cGNh3/V/pFDL8T/6inguB
s98pxUIFyDVWRoShVPZkPp3PMOuLeSu104/J3jR+M4M8VfxgSpRV4bldtLJo+sP1
Rc4jeqwwk+B5xaFKRIReyRi1awocn0x4MeI6iNiLj4PgsyZn0A7n/cwqr1gOaqvO
4piwpOx1uSWu6YakRGXDdZgma0iHbQxMVvPeIsUNHQ5bwDSNjvoR4FCVYdsSWtzN
vE1ZTnvnTzAkvkxDSt+YAjNJZ5Z+dc4BAKo7hTcVNjPCWXu0pE72UI0jipBHEoIA
9TzksDtxdMqJ5TDlUOQnykMFdVmHbbiW7yaZTM5EAEmMc8JPv20rWGpFMD44usli
wYF7fXtOXaxc2lnzO2CBs/2dwThJPnx01O85yHQZsOnvepWMAbqHnbf5o3/sMnZe
cuQHWMEprmmhsemv8BYHktPrcm9INTaGXzzIw1w/qNJE63HNcsaQ9Ts3wzQ0Ct2l
kxvEO993UXVnuNsKb2jHUvw8fZmD3UnFZF+sooca/EEW/J21gqJLkIeQ83MfYmPk
baSKBBIe9zTDu0JrP2tzDSMbN8Kssxa6icBAp0eZQXHQwCJlpDTApRJbyry9jmJK
BdBVRAvfBQc+eUNyUp0RTc6If8ZcO7OGwA0aMBHeoLr996Oaq8zQg/c+MITBmzxl
ysDt7NYrWlBZOUKFUqqtMJG14QHJlieo12YLJPvckxaQmAXKpc2QO81zqY6KwRVM
m4V1mm+AAAHa/IPPwpfYplNIzQB3y6KjRL1uxJcQEikagiOQw5MlF50FsEcU/UI/
glKOlIDyMjFASq2Y+TD5uFAizhKAZXWnGDXrKYv0166NjFiPJ04yXQjLxH9w/1Gg
8Nvcz4WQdRFmVgw7ZYpXXX+et0B1w2zYWx4HjY7H7aY6tFZtDnMDjY1QbGPtgXQI
bD5MQCqlfmZANZlPiXaHz5qglQ1cPRF78bynvPwkPTulr5g3ChBKqMjKsMR3uaqC
ncHm6A4stbVLamxh8cruuFPeWMwhS36UDXAselF4Y7kNZCdfnKfJQQZPJhtb7+HP
/DbzDBK84NTDwjFCokJneMQrgvldIhhOOHYSzKHr4yL6MIN6BL0qCzGsw0qIBD4U
V7WBjdtPjuEQObTzx2uOI55HmXxbSgfBaAiedOqHLjqQSbNbDWGYy8gUhcxm9+2R
W9O34tb8eRRqLKGfrqy/5b2dQDrnsFmzed/gQT1RdxLslCbrj9UmgpFYuMUcouBg
N0BVz5eHWqCXgM4rS/wfmqMbCf9IB/ei332+a6dnkZGm/FNanG4wXM9kV+wUXH4C
IBw6oijEtnFSys6cMzoCMjsae/slTQXwB5xptC3hQxLUmn/gois+MGocFXgVaz9F
7ZKc6zoXmGK3IMhA05m8WmFFhE1Vd87HvP7fGbvetaupDRxzLgV6DkD9p3rrq+pc
SbeM0Jwjmm28HHlpuIhsctwpZnRMnoc08XHMHAs14hj9revHSgy63qOmwrJ2jiyg
Cou0mqGbvEN3rv/E3rxTZw4u6+lNRiE4yUWXxWE+rvwvC+7rfnFGxidQfBHsmUqa
T1tqtEUmyZVFVNinaFwPmQlal1R5DwnRkbZjmbefozvSNUI/Lnlkt4AKpJ9OsRvt
DAmzuZLxu9kPeYekIf6O96N/uN4GiwscAWI/afr85a4ei2ir5eN4jWGV2/pkj2Mt
6sV909hWR04Am4uUsjxzO9qwg1kUqc6rLSxiSf9IjRkSvTnL1jJLX+LL6VEqct7f
phHS+WlKWyJZ1mEq+JqbMlxGgvfjfwDO3x+mbtZ0IZAfS6TtTbOfnpI+CJPrrT/C
5CJO9c8nv9Gb6jvQJ8NusRRuz3qUghR/odirgpaPml5qqg2vwh2vD+pSNCwHs7Mf
rzrqC3gUB6Dv9VB0SCx8cxCl1EuCQAqtlspjzP0bd8qxbda58i75ZsdgI3FhYg7G
j1Dreu1svQIme5t1dK5iF3VFNWV+AiVl4IyTVmEd03UZl0b89irPcWTN/IaHd9/l
GSoxMP6Sj72ODBno6tlUuPwShoDnAXBT1OxDcwyCr2QxzgssHBbCUG/6BlM+Uz8H
shiC2Z+bpvKqoVl60RypXktiC76lKFFFoj1B0wRJXtwuFBmLbOe2CLR90zQOtjxe
5dWXTOUtyTVB7KBthkqgZsxpS/enUr798caMJ4C4S5N6rYcbMIbmoXsH3dUYlF5w
b8srHTPwWIIxQDH6WexsQSFe0vk0ky71Wpb4p7F4nBqmuo1TgS7PFbXn53Lhbs8G
Fw6vifby5tnbwlC5r7Qc8Vy6yQeZIimsAymS7KcUOXlQplE4VhJla5RfDEG0EZ1j
u9JIWErZZQOAg5/cVc4EC9yO8nWUYHGXOIGeKTltKS8Xb4FOGmn7N+ECgpSPxJBI
WkrluJuEU2KwiizFfVS4lK4JLBn7+y2QeQFxBBFU2OjI5N5SG8MNVx4GcqaGEbq1
qlckEFwKfl/Og8h+HrtCufztyOpYScpsfdwrAiuEJEXwxesQ/+QzsDt7KFG+tiG4
qeg5vFAm/q51xkt1MWZ3r3bz93okYMcFQoSgNkUqMMkkhfGotIyTgK4lWMGwqpqh
fe6wskM88l4RvHxIAYI4TdoyX4X2RmUPYTWBS2ciRcQ3nC+JyQXHeHzovmNEAng/
ss6wdaVDm9eODS4+2bZEp2nNz7HNxaXhVD+sIotnpaDMH0uVhKcI9XLZJzbP3C3+
3fHCU0Sp59FIYoqadXt1izzLnk34Grk2Ve3GKykny+ebfhbXOj9ohmyYPK/vNDnN
nZZTrWt/RAciwVSJwBLJxBCFo2sFE6cZkHW5XbaNqCrYhmaQTQsll3VPdp6IALfq
MLSUZnKmspGg7TC2ZbGip4fSKayy3Oji2FIBhbMH1yu6dYO3+26vkWH4vAiMoUog
yiAqslWzAmMG07fo541nKu8ZDmiu4/51EoU9coQilWTc2bSlmhb8c6Euv4HjvCQP
uf38ie2txEPmGESK2uBP566rInpevNomOtdFouO9HMRiDNPsr4lZP+9lfUxHvwca
4kwGXkr0SOJODFBYwDuVnx2HdPtaBAWjJDOStThKWXb/6WnjudKCVT/ZCEGcNWkA
Ef7GKVlcu0rUeQVDNFPJe2suqhREarU7mfKXDgvArr99Xuf2xesFiJlZ/P5xfA+0
2GN5zaZnQMRhSNTQj7Jnohn4dIFckojSe+/OEuGIUdCbog+SVvvP+9g3KT1rXatM
eFpAQo4A3zdTdjVuk3a/qlvUWCxSqQ6UHqipLbrk193qAHCmb5ZYDbrSGXMYu8H7
kkkLyfuKwGXpNFPZeZyFV41Guy/OA0uuBDSxgpzNTAVbEfmlQUDEYoqJWKdr4bTI
Ft00EfQuAM58/BDMgiadbBmNw07zM/opJOedyKP/YiGdaS6vPxey38jiBh9GuXWY
sk2qUUs3SWiaSgbl4KF/x6e+o5Lh/4KNnuHEHNU/zg/T09LUFqJk6XSby0xF7s2y
Q/rmOtZ9ij4D0dHj2bRBvjCROSC+0YMOElvudVSdKEpL9sUR1smjbhJlxAr9fQ2C
Bzr/7tJtlfIW1mdfnkJTDaQykALIRAfRFeD+x35uv/pB8bkapG3XIc9Be3S0bFDq
u7UxwKB6qV5I15sQmj6WXelf6jK3zQagq5d5YLeM0ilHonBraLZ6cPCMPBVNyeDj
a32PWpY1DQAe1mcDwJHm6AMExYRGVFq2ft6S6RWsswxAR842676/idRa7HnCIbHh
aELd0+qMgjVSmrP1Xnk9m0Itl12sn8b+blzY2ZEGSPZBU8IjkU9z9Bn3uvnNmDdG
cihWH8pk9oqS1e/P+Z5EGH2QIeDY2IygdZkwyuUUOF9/ni/h48A44nA4YQWNW2Ta
v1flyNsC06Lpm49xIzgqXYPUaPO1nHgnimtQCidJRTLSmq9PXLynIEn1hgxar7tO
7E4cfVFu0grbKo5iuBdh7W2WSVDCVR4mYWiCdOTjnpa5ObdWteHkrd4OsmV0EnMf
dT6U9ILg21cec8x8Gk92gAJZu9rg3Tj8XRTzus+oAoqTy60NvVoAcvDj0R2SD3qx
zxYyPLbSNyeYU6GdyFMc2t9cGubg06kaauE92XHRoUdFDkjmnbM4zImx17rDIo4d
0E6I0CpzMD6FJ15iavqjAvi+DeCKNzbokI6h4myYmlIMYb8JONHzH94lOVs/4Ro2
gwzetIGwPwdjN281ZraaGVNHVhKBAGVS2H1a9Sf92MoQxb+Pf/URV7TemzolJi3D
P9YBR2tXKQNoahRngQ01E/hoEizNpanxv9vQcKEsoRN39az96Ti4RVG8iP3oS3t6
P926dj22CmlFYJZQwQkmf55mSkKmjzPlJThIZdJBawEU84H5CLZwUCMZmnZfi851
w1fXu5aFXAqZYzUdnVkRpK8rHo4jAhsy6FqGn++vogghoY8gZX8z1mPTkQ/YsPbl
E6fu6ANLt2x97R59RAYBVbCUYTs3Xt8dEM/Ogyv+wnbv24F2oL/l5NXcqy/HApLb
mxRf8jUwzEDRYZfjBCmT+IYGw1zEoXBUZAYui73OcqNOwaRpVaVMoFbH8mpvF0Rc
ySh6BTYQCCHKgsHykMlWHtPveLAZfugh2KcYnVwV8267tsxm4Vkf3LMPvcqycHnd
k0gqQa4W4dA9VilmIcDqi+yCH+yTbjjTM1gzso6qnwivIl7PTa7Jlju7zC4p9S8z
A4eDSw5WexhiiTXH5w9ZT7F379TaU7/PxH0BS7kyj1WWtCEdMG+Ruj8tUbLSGSTJ
1Xgh751ZYRskiTxedmZPYAnCddSMYOIOKWksSagFHdM5Efx48HoO4A5H8KMKrOFb
2Z84sY+iPER64um5eBQtAZSlmebF6CZPc/xMqG6jpV4+oEc6ZPd+nhZfVC7Xq7ir
uhun3S4AdwS+y8VFl8DYx4FhzfDh7dvk05jMzLlEfU3DVkmNQ78E7l6oq+hc/i0X
ESvaagczEsmxYeUsp3HI71mpaYoxxrGKLGj/+0asicrOct8ZUL+O2O0Kz01w4Co/
5KN10lelBNxkvnRuZvAAlikcCTopSWA9mHaFMuRIpped746byuoWM4Y1iqt3wLNV
jYbPVO8MkdKiW5/kWRYNOSVaQed00OF1ZdFn/8yj1FPlom29y1fV2zYOF+DkZui1
8eZnf/kApMhaWZLk8jpKgiJCzf8o+rn+vPXqXOOl1lmTgHFLXTxk2QpErVSKaV1R
3gKGceEVfu81M6x0+q1P4ZjJIDvezPvVEDq1nRHBex1iB/yuiIFIvU6UrKm+oPa3
7oCLNsn39koh/mX6eqw8BLe2iCzxLoivNefhFm+gy9rcEwG7yHqa6YjGNfBgv8v/
MfxGrpyYUDwBu0TFdeDl5cQEIgvnjmh5wuaHPCmKpDYBKWwtNSM2O0YzdwTYMfh6
Jd9PRLc7SuTFEZHBiIvPrXPRGL2EQb1GuOjB/3UDGfPsjUevHu6jUUs9UBcjfibU
PZzijV59qpENQm4quXnfsUFS5ewZF0qmJlXxgiONxp+S/cesdrBREkMEM9AySSwO
96AcMc0jIeXww8kw+BphJGoQyjPtQqK8HTt9n3/DMTeogHstV7o6WYyO/xcowCjD
cp2U9E/kKlqG5ky/ROh2Pks7+NCNLU+6q3EiNgtlMuiJGMz/27r3fv1MKZ/8WO4H
TJPXFPT9EBkzPhRPh1pMeIxnxA8uQhBEF/9GlEcwTKoWFVXOL2mFBuxWEj4OHwdX
VmTa2yYyqlGMczLecd9CEcz7ekUxVfK0HQkRW60NhDTBKe1EwphRju69q91UNwIZ
o4/Q+rpG1u77oP1BGtAJ/m63ZyEwUeqDKuVngLEq6ZFLj0QojDRxXbYXWWIS+TPA
tsTsJ1P13Z50an181p2jUwI9xsUtEdzzKvIHuUADf8ckV+iP0bjFXZq8daBHKe1S
pHX1Kqvo16GiR+IlGTKcUc6fGxF58TIfRvSIJDywm2bDs6Rf8cByq9ANHobav+KR
dsXTLFqrOfYQrJqlESsICxoN1s/HjUWQXKBj6Fn9p+DNzTl3D2g6ocRjhD68UUsX
MPZi3XxmcR2qpY2VkDCo6R780bdr410/SuFa6jECfl9qCf3BFAIHNFcGTNeapzdi
mY31hnyx0/s06vZWzWX3138gyZpID/nQZU83MGIIvQT/PES62DOxOKsP/mAtvdOQ
peJobJ0TwVmSHWBgNAWsd1x1/VeYp3X9rAOB1TWog3wUzLGISuh1b1CTopwcOazp
j1EHN9/p3lT3nvl8/5W87iQUUUl4u/skx2bNLdoIriHvfZeUu+teWj1+F2QgKxDQ
x/s7vvA6aS2cu9wH1eszaJqGk70rf3vFRHPvYudvVAyc4Xf2rU+xKjBJNYFLT0/E
+XBiNhIc3swqX9pEXxPkJmTYkbdLFNDJHpwDtvVMPz2ak0lBdxPZrtynmtT7C6H6
rWSncsdQ1UxKjXu7SUAUSdoroL8nhDHI+cxhlwwIkyqNLMmt5EOLkw6o7tySNOjA
BIUcqkhDfT58P7MAwFEArXEpvflZ41kGmsg0xS9VWV40jow7iumdpff104Ow4rJh
hamxxxLhaRz7ADwIaAVrQBDhq6brVSdpbX2ge7HZuz6C4izKyHrZRUrFaaCSNp5/
t7ZQPPMNehtXGTRWdSjIk3l1VMWMmdkXHvy1zh9Zp8HCnwMForc5udLS5it9BZD3
fS83t5ImmZl71g5DNcR1LRxKG+MV+8wZ1rfyt1wDXO2lORbzPTbcu6BvzZBsLEG1
Iw/G4eS9shIcu/rkcrHYDBYdbQHTNjBfiksU6F+8mtgEjEt2NuLIq4dhKxmGRHB4
9hGvqwDCHp6PSf44vQ9zDWmFsQqogGMyCaoeKKAYqpQlIe/AifotYdSmflDVUu3q
MlGIi7szsBPi1EUCSL6OSMIgWiwvYoRq9g96N7xXFhnJLhNF8C4E9m07HpcbQune
QWO1yd0lolHHVH/iVbW7nkB3dc8t3W4SKsBweOY3dHHNDciJo8U4vh2zwfmM6wep
XPEJe4loZYtk11P8HHYeyKNDFG9+xbVew8W5xW5hjxAnh1eOEYPabUurGCNf2ZoZ
KsF2hoqdzJUEutzRuprA65nPvKgONcXf3WjuP0WsOK6uNkz1jof/cjugWsDtYTPm
bylQNmIzH7rfR68vZhx4OjbgOkSQ0bD6zZ3zV8ZhPElzfhoG2c7JCC9/zTG8f4jc
wSxLPpVBjutjtpLaZV/RkmNyKiuVwZpS+Dg4pxy5FCzUDjEtOr3e5ijeiHXasXLG
iWpSnP964MYo8G+zdwaLhXiRuPX45Mzpx/bqbdjN6UiJUIwjWnphiWYYt5Ha8EUW
rLmgXf+XS7jC/jLah2H/5yGkakOxEeMNR5A+6Gkd1h8teIO/kU9gVrLo06QigBVM
vn80vFb0EPWJ5+T8SKxR2vylxKVsgAwGSV1q79XHPk7vm44xZ0QMRmSdyfVbRsI4
6ow9PBvT20jVXApW56LpIP01b1L8ygd7mwe8eEreoTsZy7ESzmyHwgJz2SCZPT01
1zMMG0xvkdwEBfjUU5BOcnu/FrUye+YVNOodjFmU8je6V3rBAScQ355esw7nfKWj
qsV+RQO+1dIf0PTVKyRjNA4CaJQ47nIlloOoDiltV2lWbM84KqXRxcAkG94MJpPe
Wzw430A/sBwDrjTfmqqXCC95x/LgDTXegTBl9EldMeubHApwo+8p7002IBVPaURz
6FaMgg+Ts/1GNurWHHVlDdDhXJq+6gBJiNerQTKlJdPdR6F1n+ue7TeJjPHnwnzl
dA8Su/qZKaHRGQSe4Z9XDnOwBV1O9C7rqCYT0CTtJVdDneEcNfzUU5fmNM3cfEex
cwQ9652QPHjsss0V4YS0kqoRKlaMshWd1X/bYnl31Ba+gtzkmpgQHJAsvVO+966H
M6eB5TVXHRDEkkwVnSjigRNkh+cYuRo/VDGf/6ZB25tRk66PlrBDc3vaeAE/fqon
nHvP2DJ6BvqyjipIdhDcv5hQZerGZ8zPnY6dFicEwhjXqVLdnDJmL7DKqyqGV78G
/NWynV2SwXCP93yKF+fH8v1Uz3Qz9gcgeZbpCcfhaOl8S3fphnG042bLPisbagxQ
RurNY7x1DDHlzPNlBXpJ8ks7A1raG5KOlc/siaYgVoTTQmDFiN4aedT+vFg6evAh
RFHqZ0wG3DGGcexTTAKjtdL7TZZxiyBqiwK39nogWrVj+0Cr1kqBGWWyAE8G9nGq
JcPwrQCLvCvqwh5unvwfiUmc/fACchjQ/J5ZXHy9c1JFNlxQbdcjmi/xUoKeZtfM
d/vFe1R/MgPfwCXxE0jhYFZlYmEy7zYUEp1+ySOogkFAf+5es6IvCjhPkYkxRVc9
BEuNC0d/o0OEaPHkoL3bo5uDKaDpZD4t+lTOTL385/EpOLapy9IjxKTPSr1vTL/J
cU/Zalj5QuEzdPdTzpAVWc5+NQjvryGyYVdRJ/TpD3s2bVz/yqgas0Exc7lVhr2D
Y9LY7kxtEWumEhV0t4SPmWGVpkOFNpmHqzygjD5P+yj4EPeHLz/JauFEh/8fQ48F
jwOygZ0zYRswQHj0WfV3bNdjKWZTXnBs4x/qv3qAx0uqzfJ+zwj3LJPmK6VxYjfe
9rIwH44nVxwFS3YjdvMEvOMOnpns0qWISPogTv6FDKveua46UOBSbO56aa+JPXoW
544T0+NrBCaNLpmno82VzzZzDRxlk/5/hGNWIxt8lyVnq4d1VQsANgJZOtsZF9BT
lKV8E4jCLsYW2GcrmGSeS6aWP/2aYuwHXgmMws63rW2CSA8iLeGkBP2bR/Ku4EKr
qHp1zAe24sgiafHN3XMVM/0Lb6zb0YDT3s2LPWdQSu3WWJSgiriE/n19Q9LJro4m
X/HEhgca2teVAjjYyWl/FjOLFblQLyNkA4uLJGJ/tWO7Oj4SvLulDDh7kyGIArP8
m9Z7/EaTseP3sBGsUEsl4xlpRk8WihzMEa/+8666LAq+z/XVWyyza4c2qnuK0ky5
OW0mv2KhuoLW8Xr/h+IyC8Z9i/2+glh/lUriIBc00+3YJD4mgzG0zRHB+F6ji3X7
EdTqWPRCLysD7P+m2AwbxkLS+xU3M56iqZo45VHQguRKmwY79jtuF3tn9L5yGZO1
sqCrZSEg70Q8BuUibFwwuPt0/VU60w63HAqUdujYb9WqJ3rTZh564yIvPcht5zva
tnuoXUs/ATCmJzE423OBnllyGsPoSSOpTkxVuedhTxkig9PtMKF2rIOvLbSSH7aX
HL3m/SFQ/Wz3nhpQEy3QUUlRlUBzn0Qv0wfQRMPGmOLQlyKK4NX9SWEO8Q3o9vGI
Vl3QSqCTrb1nzXeusYK7ATXI4mWjE2ts7g6XYcXKTI8vUYTXG1UsHTGa9NL5r4lJ
MZ5QAh1ScU6DMI28/bgrGRB7MWv7ICij7tA++jS5RLqEQn//Dg0J9b9ts6fu31vO
fvsuUzxQ/rsw/aVipEpo/29upTfTGNVUHCkim4i6KYrGRbfHbUjdbeYxWe8Y4g4I
TPLeuzZbA5KkAZEScU401QsYe5HrMsPMapgFJkQhFH3z2eKhomN01E+OJR1vrwAj
QSQZ5dOZMlD8MrYuB7jejRr2KdDW7dYQEtb3DDHuzrmHLbMn4AgS5cVCk520t2QQ
9kbg7qHU/gooKLU7fPoIF5WRg8lAUbewfUSca+ZwFA3ZawWsWbOaUCc2/f/WJXZC
Rxn5Hn/qVmVHKmd/QCj5uLqLqsPYcrj5624upeHB1tllLWR5Uk4i5PdMMsOXlJch
IDKOVqPZw98EyvEVe5DCXnViUqH7FYruO4Zs07ym37MUUH3zsRPILmhQjfu2RiF5
NJcHtbGBmU83Zpx7QS5tz3H3WEVv6JulojXSVd3DQDJ9RgNpGFSv3rxG+GVPwlBK
MJvwkGvXza2DkD9gp12ATiK9diYhYsibIEKgve1TimOz99YT1+kqx8U9WkDL+9oI
0/ZAduHTZ9cyytgqpGt0carJLYHIIglk+WzCW7h/0EgCW8DcGc0ISx+bpkSrOmPI
g+83a4FdUkbNaOyrVhb0tVBbNlHBQBdPZMq37KNib9bn01oybnpkf33JK3CzU0/4
kXEOLeRAKarLiNb/jE78azQhCIXWPWI8avF4UkkT08wx6kZpnGYbVTxeGJxvTZ5u
L2pHXBGvNOUNsyEmJD9BWMfvhzLjOJjADo0i1xID6fg9e/Kf0UD6k1WvMSbf9kdC
g6INRvW9iCtdM0W6OYIkjrvnYmHGoJcdI0BTJUQhRCftYcsBTSVMF2OiBBCeFZ32
mhzH8K1D9DCbOGb2c5vR7nPm1O2aivfRQLFDt8bQA3rMpYh2SVyr7nlPm7U5LAtn
aNpHt4MNYcabzRL3KV/QV3ZobX19o70DhNykaDEumFHvAVOJY9tfkKFHULjlUypG
3h9gWoJIVkgNxHxtS0FR8OymWVfngnsPZxbT6HFi/inyF0YWPT49FkoDtQ4nS/hC
3w4AnPLHziPnBqcaJvCRJkw/9k//43fXTii/6+9XJrtJK6ZYwFahN3+PyRd2TXmn
jPSDPT5DWs/Fzpu7Nyan8xIL/RWWrP/1665JXEutN0uYy5y0MkEAmJvs0sYQoz6x
kn+SU/5OWnaquiZGCvMe4In2ILzbDTh0vNnpGh0O1M9/avxb5WyJjuqrYR2flAqm
+ER2UYfxGjhrJqCMkvRHFav6+KwpP0yLPHfxqKKfl2lpbOcooM2/2ntAnPNjHjPa
fzJpgQc3Qwf+uFhQlKDzAl1teCSQw2OfKNbNO6wsRoapuxy7giTZQdX3wE18+TzN
JTa+1RDkI5V5UEms6mn5/msZQQ+fc3xCx7gFUOeK5DEsEavPRbfIIT++IMvox2dD
eNc4HIyyc7P4c1UifMlymLkzVHzU0VFtLLUbuLXbxNS4Iovzxwzk7ZN36etn0eu2
uxvZms7nMDRACvdRGfVcJjw6amxCBsyXgYmqHlL3OSmxvdflL/QA2ZAGxtPTraCc
/UsEOxwrZhVApawnRq8Uz0fGTCkIhtNc2zVyGpZnbZlIbczIDJARu7HKqua6ovuw
Foc2agRwxYi9nR9GGcHI/QOIvk9c38Q3sIUwYzOl9r8q220YBLvVBk50bfeQ9s+c
9SpSP8jn2YWAEK2GJ/3Md/dCEJ5V06c+RueqFZ4P17vbT4snEM736ALh5J7pf7SK
aIGobJi+oIwGJTDaLJVtCwk5WXDWLwodn9aPFrtr7HLNOT5bx52Rcz82eJCTQQjU
jQHoQc1ASuhLL0E1RvDeufER/4083jOjj4U7Jip74C4eguPTk4bvCEXnwG1vpWDq
GAJG84qkJbZVXZpBn92MdVr4WI6UbtriOyUeVdGi4F04qB+mf1K353ZMJ2dpw0nM
l32v4q0D+L1iM6d6fZgdMYyCkVzNyC8ZBVSLz/ndAHACRmYnI0TPa1W85Ea6lUdh
S0y2hszBxJQOk1ENgkYCBYWBdc5f90YLtnD5MSgLOao8wamS0+apt8Z6ktt2ljsu
f59l4B3LhySSjIAdhVD+zvOi9C+vF+QfY6e1Bg1OOQXA3ruZ0EgV4rIMEGq7ighx
9hSaUXQ+Cnsdei0FtLDZbJ5mzq5opHTO4fQa2paGXLJt2Qm0U/xVf/ZWryeoqq1+
8kXXV0oDJ0RbmJlv+NLshD9rRbwszOMrK4FQnS8vuLHRpSLzRijsPa9Xv/yUfXZC
N+sidWMzWz+gwDX/anUlksscFWcus0uJ85ZoOiY0Kh5fF56eq2QDpnfa7om2YP5E
00oNTlSLYkKMfL1az3T5S+WcJShdqYWZV6sEdh2zgJcQO3j84jXxuDdTuK8upOkS
4cegpKFxRROFuSSy2RlL06ZuUsQEpellhku0SrK2jiTu+BxQUaqo7PxWskd43tZ9
BpJiuLJBz5xHfoNjyeZ5D9LjfX7OWwH5B5JrlBmPBMW+hBGL6eLV1ZbLMbjXIn4H
QYWrToZBTJjX13DhfjhVO4YYcEEfwOI8HIrnO4EoTJOn0CoPv8eoOzvHQYS8nXFK
3qBR5shplvEMZ7HlBm6Rl4/fMOlBwdf9EbMB7INl2Y+j3pdk1cHQr4+W1FJLh7e8
pFPb5lSO38QEiAZtvammzQM7rg7S3116QY8vFabQVcaIl920aFD4H9RYTpzaswzL
wjcFRceUrrcCZzpqNxnc74oOczDR1d3FLTEn32jYKasr7Okuz04GIJbLr4XBFq/I
c+vopdwZgYrE5Bu97MePUZ5PbPVn0CVcEO0eohLKcY3qlP/VuB+UG6WYL4QiU5Xt
A/nxJbQmeUh9HB+9NVtFyV0exX3kPT84PNvIbP0O0i3qC2IcIcfJ6GxwFRWocIqF
GM6crR86l4rZ7Z88MBdDg+TkiT9JHGS/ydUq1qw8QhCfjBeE/3+sh5WFsZIy31yl
Eo+crM5kPnMi++Sf8vL/GDtC5gggKH1xwrHz3WdIpFVTrUxGRL9KuNvo0d47vr8Q
Iz8r/GuwfwRUV7Fj4ztBWHE6vaiGzpfbJ909PEzw4g1V4t4IHvd2rdu9FlrZOl3V
pQLcmWo3oqffgkTnFkrHfyqXa/3XYwgVu5ybf11XhnCn8GAqSo9bWnr9o+W0zcUn
+l2lRGILg/D2kZ0u8QKPPldK+5NZrfJmTyaoC/P3ToJbp3yrgJ7C3haJw4lkCZ9A
rWOwb1dsGYkDa0ya4zQU8svwebiBmxMMehcbX6QMMZTfsJhGzIUDVfmOYO7HM+JC
odu9fvY45EzHBpa0ZwefSJ21vqJ7hdAlTck+hbZ5TbFelCis5zzZOrLFaHeqaUMZ
54Gu1XywG+4On7hpudOED0qaRkYy6zadJs6htx+wgzYpJiosHJFjTYgv/HlPffjy
0nXVIgmpVVAaRVJ3y/tFETosoQ0X/1CcX0jLsU/xHQYP0JHzVJNoMWVfFJnolspg
9fwLJezIW9/nwRia46vXDldU/B9TIKC9v8TcIMsHEDU3azQYw8ppaH53jOfLOgvG
2FYzGIx2ReSblJpSoUOr5FAhGw8weHTrvBtmHgweh8gm0lsxq3nKiBzrRPpTsf7L
NuLIIH4m52GXoyAL2FBgN+HNAEbddZ6AH+1ban1JLZUrtn3+XTazwwCCbsTQhWmo
QXa97WY7X1BM7yitKDREQqlBEN/zHT/97w3PJss8GtGeMJOCZ3uNG1RAzmMTRiwE
Uf2rtmprkHOW8Pb591TjNOS0K7g3DycaIJoCr5jmstxUbEdJPoa8BOTh08jgSGnB
tmWEyMlLzYx0YdweQRBQoKvBafNvI8TecyqECNS7myq7Gy2+x9omjW1P7YWXNI1D
R1kSW22GmaGkb6dpuh1VNSdDhz46xEoQzcR/C8MaT3bVsFEzKFPhr2C5W2Wq48xG
mixyab/iOLrEC/noS0wHuznk2YbEMiC6rp5AU/PC2KtfJ8pkJGBbk0b7RRMk/hcd
X/SVu6QRQUemghDqRgmskcWBd7/XAxikg7gc7uQBz322/sDKdEeutNt6RU8jDO9z
QDS55+/nNK3iw/UCLK7/WFV8upPk42viBYhTGw/CSm/7NudZJC9OVzE4l+3ss3N9
Hd7Kgvyi0xLRFjozh0W1dUm2oY0UbnXT/oh8LJxDOcSzC6z1rAF9bk377GQMKW+2
FYjweotzGfc/m0yrManaom2NQHVqHUK6bLxY4VrqeJso6ZLkkTdambJwdX63wjLT
cnePvnBqPd8n3XzEKaExtFQtSKfZj+j+IPgwAAM+59MJM2OLFmsGf80T4XCBVKpi
z8nc9h3XrTEHqjJTHfB53FUz5jM+fgcVYpktDKwEcCReq/USxjpCqrVrS6q2SEbE
OoYKjgdiaPpreIMGNOjXXIUEj8wCPuRmOY0h9kTUKpTP3Nm5PYDlp+IMQyBzJqUv
jLxapTYvN2LeaEhpnSK8Tmv1Yp9SdlQXlE8gnatNEvs7W4Q9B3hIRdRXuqpeIG4i
w0AzYuNqb6EideoryRFNp21yD3de1UiuKMJJho2N74ZbeNXqTdv7iaEoCcz3yhFq
jBrScUhF2qz1hCz5UgSvKmjh5NWFfZRLKCQjGcYOP5aNiWsz5aNfOe/aDRr6/yTH
+Gbn5FHF6LBBSAppd5YudksLmBWqAkHPyBVVvBLJrGtHLhZt/9jA4rvooKpIL3PF
8dY/SN/beo7XOM7pvuARd1/KOPqEOMfKq3NcBJcf464KV9Ers1CNx2vxFYxEBeaP
F17f4p752DQJFGGZXphfIEI4h4tOk48kJtVXrlEDHKaDxTrqgjYBbw65B7/VSNkX
Xdvq6tlztRB3SdnbbfrrqExsgIi+6TC9Iku1cJtXG6CJH20pQP7dcEBhwMwrG24G
gfLRYsBzDnZOo0+ub8TliuRCWA8xVs+a1ApcA4hdIRiKWptukkw5X8PucEFmoHms
7SVeSKtbK0nmVFkiiQgnEjX7ih65zWOfS3KuBIiMeq5hnicBPjFJxIIlUE3VLzv5
f5cG9AG5diF1bJGui5Qbv6nDjfahYFKDYmrFza4afC7pNlzFCU/wKn3fdZ1e/NDF
cM/pitK+yzosVl3ykfMlfmtHLYGmlhNVExwa1cfIRfE2rkqttbHJrkdXIIU0sNVW
Xa20ik7++5nJ/R0qjuXlzH90bEXoyNor2DXkctiNhZ2zsF5cOHGeqBh0fJpYo0ub
jh8njtxDDY6f33SyV2nNSL0hn+J2Z9Gk+1aQdacu7qm+IwPs1xICuem7DVRHsTu+
Yxaxjv8rdCCLRnQ7EasWlAxCbIen4pYuz41w6dWNtZQbVVi+wG5Iorgi6MDb5PpA
+dmOd5MzdAtxAji8CtZf0AbJzQsKsciZVq/0V22r7YjDyuOUzks6HxQxZVM22FWm
X2RjXqh0FFCCxV7dj1gZdiEibsQQ8hxFtWhktJ3Yt1hgLWqHyle7GkjrPruCN0pm
MRcnaVJz56iSNZTqGMt3iGpQ6hLdQ5RNoQ4rXaQuL0NilrOMsN3ZivNTPpA2wSdB
TUISY3q9IeosXGWtLgFvxVemyjfFKVWza9YuOFXnEbs77b1jpWBmPxvp5wSBdkJL
srlkCDKgqH1z4OuyxJK8oVFbE2JsphWSSgGRK8Gf6V6RpIhuoq5n1BDYCEPyeJl/
Bja9A7LWXgcF+zI3C53SsF3w2zwFIAl5TFffe2JMMc3zR8TetL/CqbtV19LiB8dX
4UBpvbemRq/EzJjiVtY6eQizA+yF7A073fJdSjKTqFDPU9jiBhqOZij3WJ2g8aCz
NOMjhC+Jwr9va8kM7rfLtEpxceETJ2wTGImBjX/Cv96g/4JiWWeIJ1+CcoGRgzJ+
skr6SZhH8LG/MwyEBX3n63hk3jrtWEElKa1bpOiZBHb0ajuwFb1r0WGr4ceZ0YY/
BCKkiazUCeQjmkbC8v0Qv8SiKHknbGqxUoYiyuBIr0dOSCP2otgiUeu284Q7F8Ch
hb+sK8EfS2fWWQv9Jb0D7ttfSjojPV6Z7iM+rYutbb3s+4UgBGFgLhiR5/h0lcVH
ez/51F6J5JRzyv6l2JSmnS5xhHDjfhAPrEraYi2D+1ICROLF1xKg2Ofs7ZPabrKj
jb7zhNUHxEt/+lSPE77WgxsvCyIl5MSckfVpN3Ie6v/s5VibnChwRtZTemFlvmY6
Y1mqH5oLiRD5T9FAe7g+Deqn/DLQleAgm5bnnLBWBhT6c9qGCHZ8IueTfitukYtT
pzcpu4b67aDLeZ3GcOW2iyM2h0sCxHt7Rt192Q2mZMHPS1wg3HQZ2NcwMC1VnPAy
EAcogOd59G0KfcH7OqEfSWDx5tGeD+yWsd+WC++IoaO4AbpvFhNOEYVtyFfVrzxZ
IxM7gMt3wUkLKC679vZeMnUF09//SA2DmwLJUOuZG1Da72e8RlVmC846sCjlGbRu
BUVGC+9SB0yEJaBJzE/eBnVrIxhRHp+xMPwRyz9US/iFM3OHiFZBURlGehe+dyv/
UNNl1bZDvHwmy4TdcFvV0KRHYDSxmjEgdLK64FJDRw4d/mIiap4asSYvtAxL9srw
BDqViBBseSGlGP/iTjXlI/TThdxjIU7ZCssYbT8Uds/i38QrbxPgWnM/2rs6tXoO
7nxPVP6oNO23OZx7QWwwgijz/phvLKbpdprTdG+rGsBGsVHiyMm6dh9kG5wUgtPe
8NjZbLOKhtn1B/U+BpwdY0xNH1BhLZV8Z457xSBv9bIiUhVncWOkmpkZlXHPYtGU
pWPFC9gN/9OAtwsk0O96cfm2ugdAEIFSqBSt2AX9s7lUWAfULJnSnyw8OxilZQL9
vEh+XqqhfnFSWgoCW4ilK2TzbM66g4Ktf2KRlReUFHOzRk2LhD80ScoY0R91IG1R
cKAZIyY5Ha6DbfWIlu7RnBTPVBHz7UYmL6NRa5JCF4o3C4yW6E37LDImU3B84qSb
5MIf0zzBoh6RJhD7M5AFfIKraOaz4tdb2qH1qX35K22ncoq+kyz5B+0XdrT7hi39
8T3hTxY4Q3KRx+OBhgSviB8T8nxYOZL+NaNQTHgLq62l84LQJgNqAPIjEdLIG61b
oSU0LSIEur1KkFFde6Xvu8NO5hb9hwuWvFYGc9z8XJE3kfV8TjHQ4ie53b6WiNOV
w1v7vzReAe+aiwSrgFFeJE0UL+Ym47mfJGvaaK0+ED1sGsDMd0u0pilcOf5fQza9
U9jLVaWeIWZqG2y0azT3jv62uP+8AVFWSy6SQkbU30YpG/6wl9DSbcZpme+Qjv+i
JA+Sz+qr9+4V2R9wjHzXcpW38BZsbkmNFZwX0VM2MRfqGMJZKp+Dm2wV5YYU4CwX
AHVVsPmYPiUGpqtnnE9xOBBhE3uKCVvmNok/LK2jKCDl7dWkeaOtrlD3RpXmPLSi
02hVpfm1wT1gcKBNAZt4rewofCdNMCss6PsVc4DKGwD3JW8BcE6/rOGrfKTp8WP7
sCNi0atXwTnNK6QVy41x3FBIeMkYHIp16bmwMomntS2vlywfz28IsCj2phyBMVlj
kCgiiGZ8HLKGOMpxKfTo8VXqF9tGcPASxKP6tl0s4FR2PpVOYAndTXjngpAMq0qB
Wy2gZC23gGqZKyb0QAG/yM3Bvt32LvhlmL8P4gbH6c6iqkPXIDwece/Kp7aVhBC/
ovFjxt1t6ynddFUR/zXbPL8nbolCuG7YWgSgFlf76OrTy/IXZDOPQCU1X9AYpd+k
AK5JRo63YIZyK9zNualRsXN+TIu6k7ZmMIUxUEEcjlIYseiBGlWLvVsm0K7Lew+C
w4rCjTWsMAVZ6j5TkfqPyEr0BFzTfv0KgaThS3fn1ZsmBOkG1L17petOx2sZWzol
Xm45o7/5D4da7LBYIUhyFDVwfmnVARDGZAkHLEhXPhIJRf4vavuE2cmwaTxRlvV1
Xw39vCOEcg/ltr92cYVj79Cuny+iJsVrn/afSY6NzMH9y0hihQl3+YQHze1wLIxw
Df/LrRQLiyg4Iu8nqWQtp4rASJ9YASoBXpWf8Exs29mbUK1Agia9NYObF8qFND6F
LqXyFo640Jx1OURSCTR+o8iZ58ySNadW4lbxIlraUM5H0/reg5yO9CIpZGvV+UwW
/4hDu35Wa3adyFd1PZJikKK9bu9ow1v2c5FvWBVQOcFnqjRLOdmX4VqK3HGgnLPo
YrwYMJcK3q+pvsHK0XYb/g+LCCWQUKiEInbSJXE/DITqudGec4zV+ZkB/T+dxWYO
sheNGCOJLlWPyfHvw5qADxPPyVq/U6cQYtFlnZZ1qrgEAK/8NH3x+ns25Nn8IQBd
56rCjjUQb8OuYowXRHpuXS6mnce3pkXW80mUEKPlt/LAJ4IaHehAg/IvHf69mphl
t1/htvlqapHcd8qKyxbfmNtbzsSK41mlJYIINqFLPOmIRvUCVkUyJaGk1ZIa/7Cm
HkDU9Ejti6ANQilGCkWwwl73GjTHsiFWKIZyhIjR3Ca1/D4LZtj3qR45zw9GoVSM
5pwqT2F1IilKXsVzyo60UM8KxFULl83TNcrMotkWpI4lRBxhJTzTdhkyUk9Crz+k
JR1xjb/BjI2+kTzj07qM/P6vu9hLheVyca76AnXEQakp4C0yt17XJu8+iFe4/Gkk
aOSGFDU9YbLfQ1v9Dezo+3MY3QAhVTDWaM5Fvdkf3PXOBugMnskl+uyIQZF0iTUE
J79SZv9yCHUn4vODdeDOuJYMqfSN/3VTKpD8n1DIhigGo8HeYVDtchail464czgf
0uifhvc0lZo6k0Wl48wB8VMCkDfBLizncgMJBdmLfX9QbAuY+JFZ3FVYNBuFtHF6
VmUZ/RgAxkshEOUHtttxJYvWc1a5FBGQz5HADGaOrjeKcgJGeTCdoq+1ZxlM5LQX
S4IgqBjIuodq1ayBWsqUovTMQcOxA4aWBOCA9jhB57o7glxGccX6lch4E3Ng6St9
AQ4+QskQnBsWRikMmia+xjama+EdqaSYvEEPyJxqbfzTt0oj5PgDQWZO77GXP42E
mcjfJ7fe4O8Gr1oovqWsQgt+BYJfbjjkqS8wM3qM4efwwIbc+zg7Q/jQaPqU50EW
hjVYagalNsuuKg3SFBVLczPaEFBCkpCvt6rGtGmRTnV9yamJAKSZuG0u8NWYVOFE
FxHLmhHuyjT555Cvxub+ochQULJYkEalIwWyztHjdnWZKgf5Ojxx+Ku7Ebf7zWBd
GhSYF/2/IoQ2jr3l220VTlydJNQkUv1tEuw4u82aHEFXiZiaLc7/xnQJa8iYr6sT
Yex0fXNXRqRNWWm6gyK+lzkUor+OECs6pFDM4j9xgwccGkLeSi2aF1w0JJDY9LqG
xXenbOsb/ShlE2LppS4yZtWmPBTB9FNecEDZ5+VvJnQlVXnSwCB5Ickg16FoVHqH
dXHXOXezlTu+/7VGdqBMyivTlDv2wRIezdhviElkwGARZsJnMbNs8K11qUGOtATI
3k+rgtxA79f8aghqHw8d8mgKk6wxlco7iaYotYHy3k5GIl2BxaI5dVjj26/k5KZy
y110ThfH0HmWsH6g76SHAvVrTnNunYf5faVNql8iyRLsRNhPeCODALQGpzvdPNU1
CpnwGI3Kkvt47wuvpBdbRkxl6hy4KdxzqlRptfNyzgqyPl/hSH1gqtg0NNFBjq7q
ihe+8uT/SXpFBhNNKRME4AHI+pbVrjzdcNygeuWpQZvdTg2W5JA32vlYOU2OPj3x
47yzMTnz/TyYhbstJ/ERM8dLOQknhu6/F+mtcgasMYx76Lu3udTMo/x2JA+D4QPk
Gp3HHhXwVk/D3dbs6cGb0jy96RBk0JQMOaXImzarnPpnxO+Y33URkeIJrNiU+W/I
9XDIdNoS8nEGi6uSHhZoecv9VShJX2i9eZZxvEza+wZd+qY412iYzYcErBExTW5+
5fth8q3nxrnGgYkVmNkjEhoZJ4NbPPF/b7DxI/XqdBJyXB3ZtqqPbRylPD4bZ3no
9lYUUO3XQVtEEkMzAg4UM4T36PRxcTcV49oaHF5Ob/TLLEf4D/cFDKxJi8nguGvQ
geAUNse/lKB00iltcmxKaZhdYs4lVSSlfRYaamskpGygF2eGAO5FXHw6A6a9PmZD
rWnHfztwr241f07Ft2TjATmaF7DN1nbuB3cVmj/9canIgESHGK7gYdwx5ZfWM8bt
20h0ZDuwJ04xeEK9ger8J3Z52YRrWKg/46k17Aejm4NpPC3wNMwAnPgsOTHbjQc1
Zh3AUrpNi8y8StRc7egBzH7OLK+27R1TmjOtnZpQjKLGt6CfOprthwdDOZb6b517
saPSY84tkv2ivCcuFbtv6RbgO/Bv5EtzVXCkkNWLMMnR9MR3RORTfb9rcwZEaHtC
oryzDxMd2nfNkfmJdM4xmZ8t+FLp5Zf3TTIOUVKYtzJeFPlHn7ZRe9LVohtUutMi
Xy2J44d1Zeh5DeNnkLvr1zXCEkleoVKOdb44/vSCOcD+8UuAbjh1eMSHb7GhQVsu
fLqg5EFEOQHg/xp75eeIx9EhLKhBd5Mc1Hl7L9cUTalf2fSBDW+aMd4Hw0zUoiH/
2AIt7D/NpkStWZT2haRzUXIU53ZVkxjxdJysJprjiIJwoZu/7Hy40vH27/8D08zQ
lZMgSVe7G/ct9oTxh80ApFEGHth1fIJc8WfWoak5q26T+WJ8jCMiPIt6akSSLeUd
9CIfhTfcnNV4xPWKXVS/3X4VMiuOCRjU3Q3v3rNR/G6KdTLrGX/VAhY0m7APIBiW
YVyoc7bkI4xKcGHtkj1yosMN1iahSykATHr6y/0FcMMQfWE6c4cIkDxe4VtXtBbD
wyJ7otRfHHJKLQyvCgV1psCkRjWQxYE9YNM/TL/o+vdo/kUBtRthFAhpM3300wam
RLP86QSoywLW7piQS4MoZVI47fMzGvc3cOVZSb3QIgOMRI16zcgjDu8gR4qi8bJQ
hByjburTFi3n51Kk8FWDY4I02rCnXRxhuzNpoleD7bCGoaaTZ17kxbfUfQ5jzXn5
Be0KYgekJn+C5kgzCGTW8oHrNPrkOO4hiHc0PAXj7f4QyktN7lyTNe3IS/cx8OGW
7QKGK6ljM4jNQbZsd6nybNpLAar3n13rmIgYJNuXPRgeOECPdADMAxrdAQVfnNlA
CnH6XMfjDBCIuE1fQ11YtFg19EVBPHtU4crZLG0MmM5pGNIpbbfgX+bmjURGYRLa
uovW7xlOGAERdCgGC3Lb7ghtBFyUtg7htBZDZzbe0h9m1BpVfRvdAcpJl9Spwmo+
aCjiCNVshqsJt8UJCmwGW6iiMGzqs/6rxpXtR/aWAu/QDmteUq1Vtz+bgUNOLDym
bHRCTyVXkpYV3kC20xBwsfNE5HnlRJ88ghPv3MaKDOcGW5ZvCZVoOHMdswOy2SCP
FLzIiNIReIxVXkFNA29/2N+Lq+MY3cI5Yh7UyJQG5JwlPFHCOgL7ExIYsbtB+ZCl
Q6RW8ymh+Kar6ky2muuwE0sLKhFZ84fCJe8HV1ZX2fMWIqN1hr+KjCBQyJd77Zr3
aOeq7Gpr9wiAbm8eg2G0q2cOcGUs3yPV+Gd8078FUCdNE1iIj75k+Mrm01Ctxm+A
N8vlbUAqiSMDO3+KM0NMXOdgPOEzK0CMrznQh/zQ9Fu1oBorpYoZNgO6aENXty24
YUFpF9zDlijD1mnQCVWSWxk8yFZN7MONlPZdx2CqVMOLeQZpXv4y2C6npojVu8Uc
Pcz36PtpWlaatFhczwznhqJLFsvV+6nZy7bBwXHlz8EBRoMQKf3/B4mvLR9+Qs50
NmTH+z/qLdf2olLdd581Itve4xH5dow7qRiqH54JCF7PtLFkmYzdVwEM3Hjtl1pS
qitbix9Pm0R10KwUeoEIGp2hz810woR7a179qIp/Nx4zh4aFtadT6l2niwC/nIZN
VASEdJAG7AUBwCorzs0KqWrNisCToP8p2TIxUx+vs6cXnzuCq0O6GHpSndZuSUbm
zvWwCYw6lx6v5wFsX7oj8UOz07/dOhwLZoeZoW+1Bf7pslHdY7+2eovQ+DuDE+vG
BYZaFng9tfBQRN5o5Gyogt7urzzM1z5m9JMzRQtJ0pBhHH3D0gTyc/xaLFQftVJk
jd7QFyIj/GJYLA0FW6IusIMQclptHeDVLNI9JWajSRviLPo71+Soj3bivpafu6aY
fgGso9d+IlM+6ivcIZNHx8NA3t/rnXfYTYqaWPW/Nz+APncWu0v4RGnkrcgzIFxh
GjXGTnL5xV9E3Uxq2uyh+H0rt57jtCAxjMiYVmcVDQpw6+bDtGonO03sguYNuHsR
F1AxZ5lDcApF2oSA8u6RLCaJI459/5S9me9X4Dk500qqjrxTAlOLCoRHue0z9/PL
5xV/dEWBhXF1VCEebzXbU8fk2cg5cPpTOaO82iduu/Kj4V+42VeY0ZynCtHpQA/P
Js+El+doo8dwoDgemWl6wd9I7ztgLr2aQtFz94ER7whW14XxQrkaKQvlokDMboEt
jI1gcISPzTGRk3F6vSNJ/LeQYpMqriK1YfKz0OgXHe4sOtfqyFL0WjPFg3wZVsxK
0VKFDOPBjF+dHZ6CyCeqbyAjb080s3Ma8mBCC7UrrI10OuDU267SmEZvthPzgFNW
9+tYR3GZsSZJh0D6ZZQrFusOED7pZ9GUwL5+jS1uufwBBp/2gO3VXbIi6qQoCyzb
pJw93/BcxYdu5FEByTRTN9HgZDn6wC0nowOb7Nl8/fie3wYhAuDraIGoklloA8gf
nx6q4frJue8kTufsMfpbnuM1vlbbs/nTph5fxnUPk+sQ9ron0AY1Pf4oN3JeAiAP
X1rw0HklbjvhGWpD7JsGzyhH4Bj1S5PRopSLBpm0xhZHQtVYYvyjaHRRmp3gihwE
NSA8C0BIam+/P+RWNNgGPdRhsfTPZdvaWIyLWtlM3MQrWSmwo2fjdQ5UWxFvKSsV
un1v4m8kSLoCH79CVcIDXPE+qR/MZPnQ8VvfQqL0O6Aep57RdGBAINRzS2IHVPLf
WzqKGa31ASmxfqE+Z2rcWDg5Ti22AQRnhzklzZQqonbS+BvWGNb5MDiK3nCfE2AK
PP3eWWom14sIGo8t3bOHixQ4LMsOAXG5GPcNG0C3FsJyujdpvAivcv5sdhy8zM39
DJ8TKzZX0kVNkthx43K5YRQjM41v9TxzIuBP8RvlI/D9OTTR9aKdCdMaGpgoXeO+
5cRp3V3rjUUTB+6WLzu03BX5DDiMbm+maj4wxxmNGMizy57YCyMp9ndJRcPRg52e
bDKtWTHlGGIZ5EZDncmslvz20dzq4R316Ft+UVY7T2SMM/1GKO7sQT2bWC/F4dE0
QKhz4XKNgRL1NsvBU4Hslt9BQCmqBkeiLnpViC1EReHxvp4LSeOtXgE0KwfPjrSm
kWQ0dESiGRs86uQFoQIPAMrtAA+AODm2B8HBTRnSAyMche6A7EA4RSqI+uvD6gDo
KUCny9eYD/+MDDka282TFs11J5N/0NBbOuqOn4b0sdSgqWCZmU/f9WvnHsFuStJr
q+8tnWHuFPM/XMRjv1i5EhklzLUVh3bRH1WJY1jcLvvZx7TvuSHSuxO9qE/ZDxcP
6FJKXjrZeUBO8EOEitH61z3SW/J/AjL6o7c7Zw0Ll49tLSWUBpfuNPBWtMzlyPYY
zNEqyt0f1ioTaW2va+BSqBycHB3QVC/8XsdVTj0W+UYNlmutdDaZwtJy3jEiRkdy
jAz/mod1xWeNiHgMYLWJKWbwhJguoG3NVOaGtzEwCTme0LjSRmDZIglLvDn+XnsF
eBHIzwkWBRfGuUuKAePUrGfCsWRKIdTxK9+F3U+8lGa1YOo13hK4u1+35CO3xtty
YeY42cG6oSiVvUw07cA1NcwJHBFq/0HVgGcj5TgYRXgJTY0MEUmrLyKvsV2APq8t
tbjty3/S27W0wg7JrRJdDeGF75LNnUC+SOvBI44iFkjcoFRzKur+AOMEl7TyJkwb
jdPT1oP87XXCm0b3VYl54OBEuUGHOp3GdxDzxaQObx0sh/bTb96Y/gyKxnVUZV2L
vLoglTm4gW3AAxBXxvH3pdDUtVs7DbKLIIaVnnB63l8qljJQwRlVb6xpjD24SUdj
foU52xFdW7nkkkPT6YYjIeE0vTqmBjQlwy7nsY46qUqanYwfrLqznI2t6uMNO7po
MI8/h51CQlcD+RPlpKP04BqsOCzsKob1gN+aS6OO6g1rmTjA3L8b+F2CxsOebniF
pvQ0r+8G1/6mv7GP379677X7b99SZ56Svw67B38CE+k5tP3YcxJ3ZS9IU77MOux4
oeBjnBeHNfGhmkD6rO397aKykPj/gu6K2SwXx5opx5Vgwu3tJeHTwX7c7niIES6/
mKEcQ9mBVQ2GpwPIG+47CbYNTY1sSVY/OXXmtRnndfd++S8xyo5/fRbMsc0IvOrZ
6mnj34cpeAzs+UgB3+qrftk9WigsgOHH7P1rz4Yw+b+jF83EWrFV3TzsxqeSxeb+
R3NHgzCp7iSYeQGeFBPLBol+HXfZCVquwiqfhYkbQ2xt8M8sNNqRKEnbZetE6vf5
QxgRJkKLiuFqN5Mo2Gqmrr4dtS12e+LrywNub76MVWBp8Q/sGPs7vwMTidlAZmKW
yb4FxFEOK6Qkvivjrt+oIpPfwy1wGFvoanPfvsG3FV6KmtsWrm58Kts+FEu01RZ4
mKf+R6ZlQ+2ANieSgDt8H2VURp08lelTEPaR5aqarleI3XwkcPVkqqb1mEhIuoHp
Nq7YGbcYATFApQtdzck14dqlrcV86HEV7+GLxdP/RQnzJ+1PQz+XqozIk42lapDe
AJehmz/qA1KnP0ESH7ND0pAhZPeaHIwoG8XH6oxzzMlKuXOddIY+ju/71ONF26k2
sRQUomeis48nIYOmHbI2Ihqp2g8b4mBh5ewDiNcLkYzShEHT2/hV35MG0wMl+fX3
A9auggtgMvx56VV6nMqf/EaPD0pHHAJyx9V0dz5f17JpZqx9NfaPPiCAgPJj6uQP
1eFlldXUfv31CX/At4lkgSX7swC7m1pdoRDSZNr0+BtHWX8n1SZUc95VDvOJQLn3
bUfmYYvWAXrX3fWNAtThCPr4KRfrawFnMvT/qW+PyVuqzeDhCgBpZN5L9fjtkdLJ
vgIVwNT6e6Dc8aysdHxaSeXbovRTKmZoUGvJY5Y+Wh3YLIIPpa1w57AcLnw1uCP7
rSriAWTYGt7c4RD/9qCNvaxQOxoqtQRBmvmlXNf+SCWlSjJZXdlnHBh0ui7GtNwf
S5DVasElcVUx8tOMgXhuL97IoBcKPNWS5rpEOgQACc7OpTAnqCvoRgfeYGsxTLrA
M6Vbi5GBR1aqnUE+nZhXBQni8s+dT99VUjYyUfVAURxW3z3J764qZQB6/gtJl7Y1
T8S5TOuPbxdfA3LsQ+2Mr39EqrCXevTRDUiFtSIf1Dmj7Vald9w+3EQP7+zQTwVS
VsbwLEB+AhwEpl2TPaZL8EJAK97vTPICEE/MQ9JntHgaIuKNai5+h0RuwU98EI1A
9QwJX4T8JZcGFohUpLhdV0J/Uxt2NUbjCsjZHMBpEmw97yX9flRH3goqalhEQSmJ
ht7IZ5hevahVSShhomDpFUJ2LEy3ZJiJK7s2bW29KXC/YsLx/oK5a/84x5neGxJ0
mdlZC5O5mwdv55YWCB24QtNFl9txAl/y78gOzQyjTxhFbomVm1D/mV7fvT4BtfPQ
FSSl6jjgmDI85zbufFHWrtSr9JzJZHU+6/W56izBKsPvlOIS4vHZ+b+w/ngQuin9
buTNGl8UvZQQBR+T7S/dwxd266T4Ema4cQFbcgRtK1l7j8YlQbMN7Y4EMT+Hr6WU
/ATB/Ej70kxD986BALuw1di5YeYEx2opvzHTSk9vryzkRA/KCd24f9TtLEQt49Um
5bnOlO/8xU5bNJkoD6uc4I+YeNgM+8hEZ4vPCK1oYypSuWxkoqiFFeGtsaW2elvr
e0nPWuADpR1O5eYgcL3qw62/0ghoe4X7WnNir+73MTZbZS97eqVp3MUr4Aby9zRz
YXVfmTjrnrLPt76wRW9RWNGSI7d4p5+YxDvaLRADx2DezM29DXXuoK/UgmtTOO8q
w9kQ2XUVteHoqxeulOc5OcCM9Up7pfya2Z0evleWB47k3iJaby96sLprZrNS3eTp
xsG008bBlFBIeCiXOoqT5fuIWkA/s5ZJc7cHqvr5VCGiOCUPHAQPZZX25gHAKWQq
OtZQJQy773QwupE6FRl3OxtfsCfiH5ao7bdApRvhRP8ACUfUqHreUOBc0dAOryXT
M1qceayNgT10ZstKk5A4ke6n51/U3g9kKD8mDnaF7DvfFbDG3IPDr0KXN6SB6INV
xG0Re1GbeojSmiRFdqXMPq3HxBRzBTiYJkBQSfxCxr9MJo7Pgldb2tmr10PyXVxT
PA/71V61CK+J41vgEJY5JsazodSaH5EbSRCVivL2McZR+07fFpD4KvvjrU0oNWiD
CzlGATozDAcJtfqPvC4ghiCEzTBTRRqPUs8A26NQPr4P1vkCA8CPukGjlR4I9zMc
hHAgZRmv8PVC/2cLzzLf9PPcgz+ypEV24I5NCzLI2z4nRcmehj6rOeamqGxknGWD
8WKfuhiBuwypoa7HchtusUIU0lHDnJUSZaQu7sGnfK7UPtBp/BpJ2jpJT2LynO57
7WZKPz2300luo4FsuqFOHjiTnuLO6SV7LYSjF6EnEJ/RNmT+QJMt0gUir7u+ZPC/
YF1eJ+oSKdmQqJUSWm6RXJHYWSCiFiQSphDL744JUT6Wd8chFenMZQOvNUWlReK6
vvrvDkxcHutmKGpgcLdJEVYqCAEHhOri4J9zsx4UFqhmdn6C0tfl08LaFcldFKBm
ttX32Zps6sQn1DHz/f+mdYKYwHsL9jRIyBVDA5H0aOZfzA7j7NFayyH9iANc3mO4
Ybz9mvMxJaXDHYp/PMgQyDugkdliMsEV+/QgAEhyMtkLDM/2M5hb2uAhF2vlpCCz
NBIBZmyha7whnf0khP89MVORU+2bWIqidqagalq1JvVVxUM/jz8x4XPz2IjxCMLo
9SSSIy8NCE9slQ2nu5ZWudRzlPqyNc8LopGLxE+gGxX4E8OS8JAaos1B/oRNrlNA
jI9zligyBOa1e6EPveaSpL3/1LyLPcY2wSyzqPdkETRpHXBWW+a/urtZZn+E8jYk
Fx0KM4i7aRqBrrBUg5gUI+dtuOtAn/fYdxJFjkafHQVDTB8eYMRanWOghDQPG22V
tHJaR/mpVLiQ5n/nyaM84tr317R8y9h+4ZQygmo8Qd2MjiFh/wdlvu+yJ5bBjZDK
BpztvkOj2HSgPQbl1OxK8Ni+sTwnR2euduaXqZq79OKFxgwedp7S0ADBkO9WFuWP
L/ixDg8D2qj1r8GXnrhUC6AYbEZGR2VxuX+QOrwsfl/M3hTtyqxFV1O9Toq3Ssos
M8Yd8cZIADfJvs2tOko3pYNlPSn59vIbuocubhyTS+AtYxuM25PEqENgnb7QzcLc
K23c41LTEkloI4ByVBcfDhMYd4FphtHAtbg93Vb0AOPMrqsy83xaLf1E3wm8za2I
JRA84bAgXapzj3nhxc/AbOaDWjdHkfxTdKTsPeGe5lIucxdb1UUsvwgHlyiUEFu7
GSF5/6EBPCo0NmXtegGkcwmBMlPIqRdvdOEZj+pP0OT8btgzWgFhaYWZeq058DCx
hrSPRPwylSF7MYpcfnjp0vo6au/RpcrhkQtbTQz4ED68Jk+tACLxi/gkz/44gN53
LV+Dl3zgsoKxOgiqowCq0WSgF4iBRZBj+zh+gB/2ufol5tuvGnADdtZlLUZ/0m2+
/YN3RNYsFIkCfNPFGHZDfTUv0qEWHbfiA6Jv06LALQMqVvmmH3Sa8Z0+SS89DSkp
BOt5flueahgjzcXP1MpUeSiV8Y+0Ijl+uQm44wRyNbUuDwdbK3aPW9m7V+jutA+i
2h3aNXg02uUDLoWN+2hdMrtNvMzqR8mb5Wqbgs30cHoZvwiaVk0YTA9YPsxYUOla
OwHFD8qdD9cw62XlEsETGqnvbIhaGm4dSuNoLaFNFJJU3JQhtp2aP79+InmvUivz
IlhxnDTcVyV95qbXZ7qdVje40T3PgTflZesB/zaxMcTM8DjJ01hIlJ5UOkzLjrY3
tLxMi3SZgBY0fcA4FuevRFTPI02HRC/EmLavCjJLlFonfG8C7PANfcVONVHiesUC
SIv0t02s4GGXrcIotGea3+DpT+AqPaFk1+hA2BrszfcuC0gzCgddWDcRZa7XK2ZL
CfsZNywKBY//3kKGSYBgm5ZcjxuLs8D8QM0u9G2YYkbpdsHpquY/wGNkQWd4O+X0
J945XZ8kk5RIkslqAgQeQ3GNGlNGOkbfTHLkcRJ7OkQotXE3MLfeIz/U1OO3YDTj
hz9QoQZoh+g3eWZ+ISpOg3zyDEY5YlfCXLb5/T0zBGIge9aZ/Q+55L7EpxX2PJ8+
rMxfgHgpUTiElo9XwJHeS/rdqlqZCJ8kiRME82evyM0/KQuSQUHbNUjSXVs4nRex
/NXhVo/pVJkxhu3g7wDRtobpCBKQ40CJgt/cbt94AZu0GPuPelkQLFHi/I5N+UwA
9ZaBtn8dK2HI1c2/ZsdZrbb7AdLPl7B15997GAQzBNZVIKcPntkPxQeb8zTZPtUg
N0WPtZTHrdQp0pAG1z4ahv/LhS7Wklru1dK0dlms06iGTR/IZvWLnKnmEagni6wg
FzEEo7d5jVPXWT3ZvNsa+6xlrGNVFi560u+B6wnk7nI00KYb3jmWGHeas6PI+5q3
8gWWNftHIygbgrdJOZAbbGjofcLe/KXz39I5LTUj3cAILrIlBqcZGTUcmu90DDWK
/VmgAZ2/1eO+U1RExT+CajazaM7Tij4dCUyBf/3VDZyo+oBy2DGD0OM8c0r4n+zp
kh4fUQOaC+BfpIptwhodd80SmC/hyAzVRSCimvxA+QHy3ubmxZdEejHarllDsDxy
Bqqn3V1f6Jq5Ey2dcwLBHFkwyWL+gA0ss8lqinHvn9tyTzh4mG1ysNx+vEyzscw2
VgIbDTdGlgjqFn8ZzlWT4A6DG492m2qNVgIIt4a1u1Rkrj5+fLrj38/1wm5vHLbv
BmJjGJzK3fkMsTERFPfXc7yuuiNsA+Mxelb5DU2PfuWJEwNFESSf0iAAZjH/e9W0
HueFUJRRGvDNCBmWrvs0/JKocb6KqrAb2ykIY4BQIrIrjc6IgybNfnA03kaTVhHS
rZ1CA4t3ow8rwuDXsKeAqUxxqxCiDgDWWM0byyAfSaq+Mc6Z6UYK+AsnqxspxjI3
RSboyWJiOwfsaO3KcHJOVPs8plDhD4nJ6PEXCy6RtbPDGdVEOK9F9RXg/yfET3qc
HKJlLXF68z2kV5fasYfDX0ojEOmA15KoaFUc1VmJrPbSD1S0hgkKT8SgY0U5xYEk
5gH2zMlnnJey/6rjH8AYib51lKmt+JRo8Y0U8uCUEMiZ4SPCCkLsKd7Lw8msStf1
rNyHx0lRGLs5xcP0RMiZ37AJm7NwLYtevRBI0JsT5q3RK5MvZ2hW5e7dxugkbQNL
5cMilRmesX6unt1qWH6ELYV1+cfjKJ5s0rskr5IJgA0VObLJrPR2i7n7b9jY0LPK
M3YSx3OjdvpeJpypuKsQ+kluC9omzmUekng2TYIhnZ8ZU7FdL9zLGZ+JzbjbZrh+
lDl3IYxQd6L+r9iXM34Osp+z3h1g4MeCsMlUcIlWUa05M25aRQACzmgoJh0hwSGu
RJWcseycwRObr1tflfpNRHbjBS7K2XnAJfui211o03Nwe7CakNKVM6EyP1mYWd6I
1GY/aRnZYlZD9ZlMiVC5I7YY2IqP8crnwi+mJdQwlalVI2pD+hNw5C065Jt//224
0i734GrHu//NTEIUYS8pRLqHPtTKtE7AYsfaQx4k60lbQJvxIjcKWvXTaLwl+Lnb
Rgtub5+D+P+D2eYJww/mGaZ0c1LjoCTkM3iPuhqCbv5d/ZVkTGm1LdR0SCEgl7J8
BEPNuBKRqVIILSHM54xGUYBZ341vFz665CilKiGbD16FqUoFE2y9KEaf6CJIfs3W
V5/6FCzlAHyp7PQXMBt+bOfnautW1Y08xA5MKulAIc1oTMPWvwBkNpzjHbGsHIBD
g/CnTUJyh0DtCuIVPuJpSYbiMaSYUqpuYjHPKDDWBNQigFLZrArjid+hlujCPZKo
/lnpU4EvSCOoueNKMZVeWs8NaKp7uByau2jg1YpGVTjZUIwJjKFT/c/IZ+FLzHXC
/5f/9QRCLLNM1kqp70ewr7kwH0yEOytp/cVI6j4ePpatwBUU82pqJdsigBfiPaZI
AOgHJcLHv0Sp3nhkNV3YmyMKimuZ90OtQ0mE20+bBE5cbX8t727C99zHOPxlRE24
CcSkbVPxK4NvFE5C9xYL6U5Eui6coy/iMcP4QJVGa0KmBcaEB2HfUhKD8AoKDAFv
gqUgR/3MIIpiaeIHdo7loERaYA9Fifh0ocjOFCXr02hLWlrG7VT2j5OHdIvHAN0F
Bm1AXwOdj5x8weuxxigf/BZwObGcJtBPNSQI/rTwMX2lIXs7tEVSpdNvQdhRQbce
f9kMoaTAcUf+K4VCMtnDxmoUc8QoxEPOWOjKPPNKuvznTckB1FXvKV1VuWBggVtH
HZiJbHPQS4v5kdXJRJ6FRPnWXZQwsGfkWfGHnb1PKU4pb/4Umw0dGhkuyhIn9f+Z
e2shTl19VUF2d22wGGW6EchxkmUkt/x3KbzOftkjinoRmSq5sYZUQBvzqAQSas4M
i/jF0VZCEcqLw13xm3BXdoXiWYnVTf+B2C2UXOJ9YG70VjNp5vn+9ksICt+PwmnG
NgtyoZET6aJNIOM5VicZ+AH71J2NLHe2SCXKAOT4/LUvfauhJbE59j41B5iZAK+5
vEqMfF8HmFqcwc3TuA27Kc0WgPpIZHVUPbQtmWknmwS9wTIA+306QT4iQZEVYB6e
AYl8Hewx6zfoq8YGixuIoGdTzezaJvO51xTaHn8XTWL/hjR1O2eqeULCMq+9YKkI
SV0+ONE5fzEeGd19c6YrF9tdq+Ew7oh/F3iRP+W7QHwCLDbGa7Wa9ZOsANo3Eboh
eL17Min7OjKySJS+jvH91KD+1Ab3J9avQhfFUAJP5kvWqeXeX/4xAVmEg9n82GbC
QheZ4ICJeX2GJA6DddsN5XfgKhZCDokux9rmgo2WH+uZ2JEHZWmqSnBrHDWei2bf
o0vY4sdcAVLOhQrN4vIZ3R8sTQSGOJom/e9VSfTtncLPIquj2CEaZ3G9FsWiTM0c
uIptGaoLF6pkYqeB0IxW+Nzq+1Ys1V8iIUmI31rmxpy6xaKo8vu/ANB+K9h478Fn
18cl+Ha7dYPXLuqxYr2CLS+bZXyEbyKOX2RiWlCfy70oUjtPvMlUDEs1kh5vmEcY
59lbnDYrjzqhr6tZD+OMLozwCU8AFKk2MBodNcobI7ScvYCt2ZwkUTxx8zhp+Bsh
UtYgmB2fucgOpuxKeC7EGNaxa03zOFaZNCWlBqIIzcyl5rtskA6vXDuMS5DezdZK
YQztlWlNP4sQwrgytkTYsehbVuhl9jd0FWcrFMX+Vp2ldZcwruup25rTrWi3JWA1
czijbj9ZtiuC6nfIHWeodRsDZ1TgaoczyBiFsh0nlhdKmtX2v5NKSxWMBvkywthZ
XQI19ALUyXBTIcAN7OWlkPaPgGYoz7/Vmv6KjwaWdTNmVHYj1JoplteshlF5nWfj
H5Ca2Jke3HfbbnE6jbjV9f1tJfzuBWB+VHTuQENv2il5Wlh4mP1hNNMEL4sNiZVS
mbxhp1Uzr4PaIDv9ApOTz9dYlFnh3Cmi3srTgFq26TLkbOjlpA80tGN1kCMnik0k
wYG3LYxfi/C22FlFDw/s7S+tCJ2xGNXOLOdtTkgA+XLny33DlI9iw0RlpCP8Oftq
/tcVPblBHip3fWfohWn3XLM0XjtEop3oPxihuDQxIf0b3qm2rK/AHmWkmLU5sM1T
i6et9TaVxbrySjIourA1F/VJxQsNFjh4CUTyUv8gkOY3+WN5yjwxEyvuEa3rrFAZ
8KeTrmp2ZAFCnUYB//YwS44L3vAkDXHwyxexcfpEN4vqLy01F9KtTvP9bXvUQ6Dk
NfoweJ3wisZ5KYrWolpuVC81T+JOygt4qIZHPjfbdpEf/fF7kJoQA9ak8gYRmFRz
woX2ekvaZnGSO743XxlXcBqSZ6nKwT8XeMit7DBUHWdETKpx7CrwDfhW11Wl0jvf
Ounw/RIu+ICJxNBBEayfzzBuMQyWSDsuqlGDIBiWgHJQELLisACsbbnlz8yUTFUU
qOk4OZg7jN0lejdLKA8vJUYW19lFa4gFGK4QGsbB5HKN389IXskUR2/2+kxk+rkL
tjh+IkUUf0/3F2uEA0cHxherNHGD/AAfDy/Jdl5Ykajmz429rnZ5hSt4g0heOFR2
aeaukun0YWUqhVQGqZt9lrdbL81zqk1bvhf5kr4G9ZuYfxFpydRuUm6rpnBJuiSw
vlPoZqHlu9M6doiDjpOKeymytX7JgzrNxSzxgKYDALCb9TJE3WoE/A7FmOBZwX7h
fbLsj2CBYl+fht1spnuz/DY5mODj6VQLYPieaDhIbYEy1AapsAr7oupXhTTM/xB0
doEAZoPfzHTc4H8XW2GH+UzB5laJQov92REFjEchtzDDCE51FHOFLmyxyLNJFHf8
MWa+hjtOTQdogt94k9dQ7z7lB8QFPRa1vEE/+fyNL//HQqvCZVerYZQD3tEvsWda
6uIByeLLHRXF4vKj1SjCSdCKIgnnJn8FZpBf+GrPACPxb/n1WKymETEvQl5mCDDl
FAhbZFHMLn54iMj9mYgjTmJjTFHMm9ywFUXMYmaUSb359GGV2zbRBdgFGcx7g3sT
FE0YkFtgFl1fpgXdzrLws5JGF9HwbWfISqVZZXWysedXFkDPd98Qlzya27kT0+hQ
TRczDIrUDTKphubGHoLQz7lMlKypiwVbkVVC8b6RZjY1YDQRxeV1HAwBV/um7DnK
/4ZzEZ8FceSeP1NdgPCjTK3fFd5iid4YaR954d1EXr1ekkx7kX+XjUwpao4MJN8p
nmZbDVsAejG3llsF2Qu4Nx7nwVStHEmA0o5WCktTIM/e7t0JbyumkTl+SDKpTCcE
xYXe944dqsyt2WjlIWjLcgmAtAwLe5ksAof2Rq4A6ExorSCpbpaJE1x01kULxkY/
+VBnyHoS/xrLq+NDyvcOgkHi8zCSZT7FZuYajR0poTu0kqa3/gx2x/UtFMYkpewy
KuoqHElffzHNEUP6rhIsXfyuwipRcLEaGG3r8mKj1g7Rtyci59+wUgQ2F2Kk+NNE
HDcbRV0ZM+RhfVvIVAKwGp711OD+qLlVW78oL4OdQokelF9z0yuu2Q7FFlqgBi8A
J+oB0v99+jw+2MPVIxA6zLRnx+PQawcn+hHxDBRArkUD0iussEeAkwYClCt/vtdS
J6yewRDYNdUxuHq4DV5fpvg+VsFMr289CP0YqxvaPx8lRF4jKQHJm2rFUvEczhHf
ZVStszeAVG6Bxn8Jtn8kIMhlg1+Hhc7toFYUVaIZnW3/+orOYm9/D3U4qPNni5mA
Y4hGDD6XjHewlR8X53iVLihxBW+26UIFkyAanXbEVeKQGt8zTT1DXyIJsoCI/2nZ
0h12vbtIwj3CqSjJ3QN8KWlB2/vJ7BOcPkwQ0tv1TCTcLckCTgR0YAU6ohp2Fa7w
VPGIKXdR4vxO4Db73YOF6YHQjp2TR8dCqm2cBwnTG0HkB2qFYH32mGNSx64v/7aK
9ylp+9awmoCkR57t7PT8NkmcpeYG7Texf8nxux0Noqz6mm/CYfx8qBy3DFFQRhPr
dJq2PpMUfjTb7UbgJqGthKu3tk+GX6F1g4/i5C7jiurH9+QKolSgDgg2Zy0VHBJb
4RHOjZ2iK23uqPyk+bivTr/pK9OtGPm8lcph1xWv2EXqU+Y85nt9eOZozJ+82t2c
0eMXMoaAq6kFUpnz8oV/4u3bXZH2DnKB+rq9xW+mymvwmo38ET6SNQTYCZScVALx
jBr9WQ4JExHs8B8w3L00rOgkCrchQh02V0w+x+dMsASNY5fPO7MpXAbvgj44erUL
1xSFD0JuP6DIrS+TEhM5xEskDhwMOEC72Qb7d1EAU6SOud11kkPMDwsTXP4d7Cht
cevPKm1VkcAb/FonZeFnyg85pPKaijWo8qAE4UbpQAQwNK6i10WYIBZngp9h6XLB
5wIe1hjgWDqP3ihwPpezE5IsgDTQnTg8JIibKok+0AYnlqm5bqVRKFx2uhkO8AWG
tRekgmhttJhpZbmCQ+tzxj98NosLpjs6KiqefXfPquYNbWhtOWGwf83+8yRsUEcv
FBD3fljzRiWWTzpoKGkO4uLF6tOJHMvGX+bupBnal6v2CHhFXZ3deX3XhAmE35Ko
c2KwZLid2nJZSq93PVXtKE8GB08EJdtxtHCvdgn55dOY6yp5bcz+X92V4vZRhQ1j
t+iiiiTbHEXo5Qmf7klDcSgaL2L5gn4WJgB5ne73SqWEhdgYGBo2kGNQnfpgXguO
PDOOoph4V9y5TTjvqvQR4O5RufTgg6mbXs6CW7l6KsH/NpxnbyKWqYcq/cEAqZe/
X7qs8/+tdLlrycorFLljpuR1E3l5+uOC7cnu9FFVu749ySyzrOaLruiAVrRKMqD/
e/hFDca5BWLW4G+HAonqjeEtz2Vc3DymW1LITumyBMhO2aZ1VFteZoMotpgeXwZt
mnY9YL0jxvmkwvfvgA3DHMPc9Hkk2YfRaj5vJSN961jhyMHspgNRd3elIVq8eg6X
vSBAdKtH6haaYiPohO55P8MhIYpapPqfb9wAqR8lbirKE/7ES8DEomAo5Fz+Ddoa
WZi7qGRPyFG18hEorfNgoXPU/npE3BRZ5zwn+IfmLFW/LqaTnjzf0dmJuvgY2nPk
MisyG3PwiwJbmpewd74XdhnYlCzx0c5QT7PetBEuoyzy7fvlTnebTQeQMg8UjC2n
YnP6qyJBN0y+FXZDWnG6T4SHT/1E2Q/fDNu5g8wIRGlVCNu/XtkPsXmYPJKc8M6t
Y/TaVGMCPhmuZnFaDVNXAc3hoA4NRReHG54t6BKqhH5S0fZ6jm6ZhrD8hn7zp1c/
NaEJzo0np5F+i03mdmd/h6pMRl1t2zNHOlA+3Cg7JuxrCADcsyYDX1LEhWMVGo1v
TH2kq0uz07Xu0kkQkIFFiTCtT4lyxHl7VgRpCmonuDTrBydBmci8tWJnf/mUOUoY
iMB4oFpXh/Y/HqOmNV9hr4BtTUncmz4YXOBaNKQ+l9DTNNf4v12mJpMLIfaG8YQT
nqN2e8kupsce/h2Gi3huYHCm91ZIIFlTciEHdE1lLPs7enIUi1VLr/G27DINa+H8
jb9Mg/HR7uLbZYbu0XpeID8VXJN2IcImR6halvFrzDD8ysWXhUu6/r1xMYxljVWZ
D3l1OXWkXUmSgKr/01voWYcaWitIGFBLtlHJomsF7cqKLQgYaA9iOlnPmZl1kdgy
Q/8FeZlURgosYx+0nod62V1aMiHKsWoLmOk7U6eHqeA9rnm+jzd66/7yDJmHBMGZ
b3LALNs7mSnxh8YRkKkOcl0oe2RPdzUJF+bUwGAhO/JvUTwXWTJdRWVb1hvusmVs
xMMuUDOeQntNsanlHk8GcBnp05beo05N4eTHn09RjUeg8R5tJlis5If8uNzF+3Ga
1eDoU8cWjRGNOCnQCEwLvOPDG7Ztd/gcZjzRquO1Ok0FZJMv1bnRA5/RFgYSncQ6
8pMirJ48Fn+w0s0fmKcpiRvpSHpBmlQBPknSUVZkSGkdrctskhgiNVFnoSw8i0ro
YMJlf/YitSfRjA6VYcGssJbiYrxXCEjEy3f88kzxztsoMOXd6WM6kKhBXazWFZPH
10qYvsIsZexmP6iE7jEEV0cwRgeT5B9+VHBrwLjPwN8Nw8tHJD5WnVLBbnCHk+bz
z0QL5utw2DlbZvIHfPJydO7gGTj626JUs1QpRFt+bdB70UxFRrMCe09RYtH+ffLa
TTlejyXFyuSgX2ksBHcLcQX43q9zp/m14qKQJ5Do4LIy4VHqj4TqHogpQ/rAHjqn
5gu4DkFYmgJbM3riVPt44t6q63NNcRgX7bc4+i3wJoStrKtV0/VLOrBT/u23YWzj
PuR8r0hMR5Nkrf3p0IX/3ysbeK/eWC5dVQCJwaDjhmr7S9v39nr8wyJM2UMvwQXp
16tvhfJGPKDiPUCRhBOvLFLUnWDUkvZPM8JjQBs/hQOYN8bckBsINsv264wcOVUn
91cJAJ+tWevSMWmI//DUL1UiuGUQCLSPklJsLVsPGfJgwKdR4wnU27tg9RmBkJ2C
z1uAMfmh+Mrm+ZT31LAld9k9Z1nHo6+3Fhb/jgKsDrdVZdQwfd6Ip10VUj9xei2x
ePd62NY6Og7A+tP7J+OZIhY4KiqaoJvAHqrzcKzPJNxNIRK8YUrS4+LiyZHbeOwj
1DEuFCLTeGn8OvRVMVssCdN9E7/ZNExYpb7Jnbd8c4JCYuAuxxbTg/2uxtEl1L6Y
/JNXPDG48Nl2CYl9PAnCVPlHJYOzlUFCaxcBPeK43jDf63bIWCyz7Qxsop0p9EzK
dKoe3ro2yrONtx5zERm76SE1yc7eTjwRVcTw6xej6a0ThexADO7QJtP4qZDfcKfE
L/Ulj4Yo5jcn2VVbegLo7Jtp4toZwBp3qtHbsLufGHld01rlcrR4tLZ2i4+vyax1
MOka4B3PT2hWcVaabG4m+D4Y8xuoO+5v34ndA8AfY4ek01dBIdUsNPg2jc5ej8Ld
FVy/dgaKeTvAUZiVZAIi2OHG11ELWnvMUGR/sOEwwTYd5CXeOM4BY1OkBC/z2cV1
nL+sGaEEFnVSzJQ26jPRoKA4iEv2Pp9VCBnxsFAWTKFfkWpjvNHOj5ocU2ZXrJy3
gYtRAlq6DkopnwvhtUC7pDvd6m/RqDTzguvkJm6ClaLPGaeWoDbwoWcv7rPBvitN
/Q0rEJL/pBvmo7Jor8syp6vihuGjs5hCSkgLAdqLt3nDgU+7YDI/pD215KfXiFMX
lev5M4kL1dgNlsJIZ/d19fimeajX/q4hf0W5XPqNBCGIjo8ytVyRIerSoPHFuF8w
/vMiUy07NkAM/PUXgCYs7J+sSWz/EQUuYPyt79/dyAKEKJ4NVVYbuuN7pfOcjhZ2
pdaJwkBZK1Ud4ha+7ClbzRKszU0W4gJurgxK0+9qVgB6VngUgXcd6+5/SgnZknWe
1/YAxDSSNuBFL1U/HaiwtXbdHdLeHmMOLqZbo5iyzY8LT8pwEV/cjGGzQgRdP3Gc
rLAuvytuaGO0XktDqJC4elRCIBKAbJuG3rZRgJyUgjk4CHwVzo5G21818SNZpBnn
95JiFcY4A9FAqATiUhaEWNNpBH96TXgt59ZSBUCfQGKhfjtIpH9dKw5ybMyROkae
p8vfPzWWLdMGn4gOHcst2rpEfCH831d8IM/p6Fsh5o1dsxJn2bCtwpCmFVyQjpXm
zcRRxDvhslgMcM2cxt7Cv+nY9lB7sSM6bPzed7uBUXZKs/bJcMN5z6lWqs2RSHPw
UdVxCFgte98y9m/JQEvR6jf2lBj+RkfnqBRsASixNFwjPoFiOWCx0u8skAoNE7gp
8vRglqW0D6g+gMmnfRhSyeZPSeBskG6xJUytQZ7ChLBtx+F9hEijKy/4UI8HoP+m
sApE+GRiwoRjMPtHtKdUynY7O8ewp9ynB+P7ZKt7/TQopfA1FMit5RAmbyGri9YG
KfR/Xg0Ke/VB/m1s2Ax0WAZiPF1n3BTnApgImK1ch2Xf8BhErhKIpOIt2uq1uPnf
gQ7r8zDBTAPEGSJi2hBG2be/bn03cXvRR7sbcHTL89GmAuHOtyNSyiEKNfjpUDKC
fds4g0DZs8TTix94l5IXDzmGbZEyFcyYDp0bmTCg1aL4JZKUapHYQzDFTMdMTDLJ
HDwE8pSRewoWWEA7wdCsNQvYglZxpLlYrhlwcOocZrmsGrhSsjuqLC9XV9BLhZa/
4fhzjdEQYnPRjGRk2awFNWpIcY1cN7OpLKIJNmCroFWujXWQzEVQoflLPGJt+Ipr
aoueRH9VhOhREwMc48s0zovWpdmkkFRn8ia4frpUHG0DmMFYDQlk2vRqBuy+N6sR
bjpR51bCl38dOogLj9wOYUl45cCLU8oYsgcjORIi0JeAYAykXjmFhamKzFZmh4k/
091zbjKGXyqxS4q4sdLeNkgi2kRloVvFyjAKEMh7SzB7ifHgcRXUfjcVDTbH94vi
Jn+hggZ2nkGylqOQOEVQjZWuAzm5qzU1MgjKzwh453rkyRLW9Mj79eVS/IoLe8OJ
/gKoYiAVbt3S8tGxq8SUfKUFC78eOcdzov/d/zDiilZItiKKCq9BznFyAMUW1UzF
jgGgcIMVxNLBu0mt78hMCnRunbZJjeaYW8IeOwiq5kEOl0hxxtDLf9dnQ++yM9jr
4c+0GrtItPeave23U8igwmc/rDjcYog9RH0RsG3EGE8R26zG33+UE9vlkoj1LTua
bkS/vmsvZAsVhbJGpQUK79qCDomfGNH0ySccxm9qO7JRTcHVXASlo9HXu35II2pH
v9zUYSMFuAkNMIIwVBLXKbosA7ABBmxepuA7NjoLmfqVMnnV5sy08BkU05Rorhow
RZVgbL6HtfRl473JYlIto6cWywzcRuhpyYt1SujKIgIme9uQIpvRwrz9oR2DKrwi
okCdJAy8ZHCq/pU92TA+xSlfhcXTZ3OcbfwsbHxNB9puHtJdszjVlQ8zo2aIkp5Q
k4+VhDO9UmGwibz3tMZxZGEme+8NlcMiw+ERRTH48vEhTlDBXMZvvx6mVDH8m9Hr
k+e1l2KofGtGdwLHns2Kt2sBagxoAUw2g6/3afsCFCHARyEBo2HFANGQef4nLYxY
56pfN4P2k/ks3oWS4/blx2MZ/0yaT7NROwiyTL9DT+419ER4qbY5A+ohqZ6J05sk
TztIeA/y9MQlSKWv4csTsVTbpaYewm0q9PwgSqAgvvqYQ8zDEX+B11ZDwxAEnrVV
DojKRF+BJMlrPJZIHWdVabMYpSnS1sa99fkr2RdvcDh9bH9BpBsQbwk4+K4/cF8u
QAPsbc1is2Z5F1cfH8Q3JSe4/xyff9/U1AA0GRqVJ6+TBhlibqQlJswBcEdXy99L
IhHBC1w+tbHcAAkNkBqCMVJWdc438w2/Qx+fOXLR7YT0Nv8TmP3SupBR6AMqcr7N
PIuPgd4rVuCwNh5YhwTTQpmFIZY1Pz1QvbrkGR1gddvcoo5X/8l5rbNpjlG95UfH
Ig6c7xeTB7Y3IYBQxfSzvpxJKY4gicsuOnfRPJGPZRsxyBrnLn5zZmAjHoXZrNWT
EDgdZKpjThnJ6PCiu+M7xKqvidslP0jJMLvj9l9zuIhhXupeEpFRLPwWM9P1T2jM
qAeXftsjDrRBXpYWylD2dD9OshYqHa1jKLDCIAdXNQP+VJOs8IDNH5R96pv30esF
7m/lIBKnO+w3LrlZs7jhuIUwimIf/RSiLk47poQex0ArSLKdC9wvPvbDEvbGaHVY
+ZssOlW6p74Y65p0FzAS1JK1hi13Igb6njZ4GmiCfFU0okQBeR1t6jdmwpn70Y0A
V9EGfrKFTGjpgAXTcrwX0Z4Q8oLv7sUYYlOP1xy5mSS18FFG/VNRXd093C4mgjlV
IUwQtP5o6UuqKRNBIiVH4rBns4382AHY/V6xSc9/GgsDx+LrT91ja8maRdouZvNY
SffNN/bSJKhoUK6PgOeF33hHMJu08zB8zQ2pG6GoSy0WcfaLmUS9fH1D79+AWiD6
jNNTlmH49nX3d5+LaOFhKxh/HokVFBGquF8eSnrtUPmBCJS1YSuCjPH9NNqvfPfT
vDXxM2meLJ2fg6DkxKS16u9fCrpoCjLCbsVdtm7KnF8ozIuYhnzUnd8hVbZgSuxq
xwCL4yd5jLIP29NgpLfPL27DPEsajhpze606rp52ZITZcH5reLyP4CK2TebIUzqp
9NOcvJH6XntZtkwAfFP37WAp7nNYf7CFr2JjnHgcAONf0Kknm0BkyBpIVO2yfpZ7
iPfwDriXp5oTdYz6WH4JAvwICxHI3OoLI4cpcwi3ZQHmDWwn5vjVWJxUug1+xC0r
g8sW9UztLDTUs7E7lBcU2PyNopQzSl7ePsSs42QL/xETvHwavRFRZEJ4CHZUK/OJ
AxNpsHGxcDWpRqzF8X0MIlGhG2Km6fMN40slH6NjQphFmTlQIER3L/LK1wSeY9HZ
LfvioMVMLBEAXJTNBoRCP2MaSyWnj+PlgX21rxlf7yy3J4+naLpGlpA+ioHSb+Sr
e6RQ51VKO4cP5ogEc2CbuCgYi3/8wx5sKt2AKk8B/vphDBcmNU7n6H/hoATJ1Aag
2DC2JQb/ugifFQLCK+f7RrbVv3w3bux5eypyd4X6r+HqbiV8gLA2ga1V4u1QGXZW
sApOItcSHiFtg5vJVqqDe67jcVkPGR4l36/TLxrMW8zhz+esCXun+y4v2qC+U0Kj
5XiyyvJApdSUMdYBP5+Q9qlf7u44tW/YBvAuC8kIiWYKA8ni/u332a+XBSKzih2i
0P/DWbwtDt7gACnWefGUg+SyKHIyqvR3rUvPyd8wqrkj6RRg7yxsVB7kjeVYYpeE
SBU2PdSM4Flru+PjS7B+7Cp5Oo/5pxwLuH1VXjl4eWuRivYQF5in0v3HmXFKgGLO
5arMZ/cRyuTR2XxKC4ZhzPFJQ+HM+CYDk61J9NJ3CyJwJQ9OmOAlijqDYrl8jaPp
u5aB0Pmsds9cbzDvZfTdGgLTGL48bURStGRQUx6lNaAbe85zOy8HDjsoFDiTdKor
P5kk3whQX2pw7uotopp+Hd8lq0L1LeDohv7wVcizoBzgNbhZCb+T/ghWBIjHDvjw
zw87yHQFx25iS78r1HN/oCf59c82MXbVNE5SYEwkYqauIYo6JFwJwUW7UuB2RtWE
9lo3jVXgEfe0JAvHMXHl8BgQ1qWk23M1hjXOePgnMi8KS6Pvkpaqr/GfhvzLwLex
TP9v1BHNNM61q+J3XK35+38JNLQ0BVdtNBcElhLMlZo29aPJwcDSv1oG0nTrIAGj
Re9KwEcyi+M9soI3HKcjIDqFZO1ikb78VGE9C73MwZeZR8pLUnrb4gJtR3ajH2EC
UjJV99AvgslXgWB6yJvztWbgnQKp45ODiarDfG0ORf5ftBwdPsX6Z2Ld83wO2Ukx
RAGrVwD0m3GO/T1AcFnC/ykaWhgIx6vOzJGNTmhKcuIg8PSrCdEm2/Ls2b4XCwmF
ftlS/ztPnJM9NUdSbZ1YAbqlvibnIg/A1CpVYQw4jZ92fHoVH8J0wgpLr8skZ2lW
ygWgdJrKtcYQld0hWWEbuu1PekFP+6QeTddggFB4wAwfF2Z/wQSkfHi6XKAMRsl8
qQpQUwnAERu0aEIzrVEK45zm6Wm/6HtLMMz6C9ACUxb5jDJnGBo8rOlXLjqz9FBx
8arT2i64AdAqFEN5Kf3XOr09Kf3PQx7YVc/41Ks4lLuwtwgqineE3EpHRjVc/ibU
bDQAtgXSoY6QRDOfeBFcHAllrf/X3TXWuBHViWoQYvPHuHBSDaauV2KoHPSp673e
GTfeVDGUCgQaSBhjpX2GzCvft0B/C0pTKCMq0IRr/fyPAXFawwuCW128YoVOSLYV
d7srPcD8AgIZ58ZKJ0w70jFA1k4nUueBE1WuNImOj2E4qx5aLMNZL81+hiuRgmj6
PygCv2WnKMZ6aiFP6Zt6i38EwpzFtk6sOmixUNX8D/UWWUNZ15M4inp/hXv2gBnP
J9sMPScjKNmjvZTtPG0nCtQPFil54CVYKchoW5kvMXmypgqigevbNd0in2eqR+M6
DnX8F+D9FHd28+mCuHTYU+K1ynQbU0Xmu1WWflv1L43ACXBptjVxYkEYzeghtgmw
NHU4APF+nZr+pRVFtprPzRsXTytusnFrjCE0/JpPQ0VmttUezWYgjBtR7Kffsmgo
MweHSztApbMI/v0mFcN7am8Tpuv2kb8Qy/zn0xMt5vrEfUFkZUS30EW/Zjhr1MuZ
NJdTr6V8W1HtUE97690ygZC5gMTlucsy/i8Tle6wNLtFK4aTiptIQmjs96b195WJ
v+gFb/WZc36KF9To9UiIw4SirJJ9PuGjPC+6o56fbXm4VgvjuzAhiAcfkWmtfYyx
NBh4tcqdnfNs80JTuhtUSo+R31TBPQ59S9cu6jEhMwWebAl1WBUcVhRKr80+3Zw0
rxXBMjJUSrVSluDWv+0T1aKHS1p+aZ0o4Fm9hS8mv+oS00nywownF9u1UXdh+eMt
vMgiXZAsRNlQeQEHW98x5W4EGld3R7aqqXa3u7zimXRqtAIOOVUp1dWv1abTVzMJ
20mTjFXPQCRVXIl8pMHWa8tsyCgOiqjDeSFa0bOE5BJYuez48gOg3OtwjIq4mYQo
e4Whe9VgH/zk6Uh0BbZ3R+P1V/xKqiDCZkqrpotq+r4avEEnPiHQ7xyfgmGLtxH4
3FkC7gSlFTe1RkFXHPmzuUd5/Bc6sKfG1jL3K7IN0sHVnFOxsiHhXI1pmc+m9vGX
LxjNY2tSgHaSXZ6PGaMvdcz+cr5ZXfgUXL6fyn4Rr9tk5C36aNNdvtZWh2w3WO2/
t5tRaK8G8hF6hji7DMnQ1+cPs0T7QREdhAp0yUivgmpAn5Va01RvQ/eLbqtZDLDj
tvzwwDkfWSoVCrRSFBF/67tlQgqAjgv9+G0n3BOQYsFxvgHegORVxp23AAmf9cAa
kRfjEhA8F1SZZwi2EqhFu8S88+98XYhzcINWMkRuQ7/8jl2VBMPsXxRx/U2bsuVo
KOKRPur2NyS5jnWRaabUN1zjoUAKXbOmKOjwZZzERxpusKf5PLsEGT1gJ9tJ2Quq
v0K5fXWqRmBTs5Y7/qh+j5dTyTrBEV9j4ClxdKBsoZ1+USRBF2Zgvbgau9b/WWR1
8eipw312PMUOV2U8A1+t2TYI6eu9L1N3zwLDcVgiYIdytsqVPkNJGGbam07nm+sN
+S+XR6jnyCKHJHiuWEAqS+B3OxEX2MLZ7aAVvBsQuNm9OhoZkSyqcuupOXy3kDwy
+jy1Sd1ZqHpdP2A9Glq6z9TEfYN7Tl14TFiHvtsswIlJyHJZuvAno4Sa1zbjSBRI
dNCsPOygc5Iz1TZvfDLRfYV3ZXvZUEVyfok1XJkvJuwpCZJrTh78chlL5lVZOjlb
/wAZf0ckJDdRCfpyqUNUF8gJ0Aoy59RaLxGiiew+lbdqXs0U719u/z9PUhFpCjad
7Lfm4ODFPLl2imhyvPW11Fboiz6H0n5oa12DKX+oRt5QfROJv5U6VjmvvNIoAwHe
m83LM58gt0eW3KkSDzfUdn1nB9hzkXX3+YT2fnX9oMItiilbeKR8m6ggVR9CfI2J
C2A6IQGWIcYQjK3FJ8OP/phQcx7hMbFP1tJMN9W8Gaf8Y1dS3R+LYoBPXUbc1NI1
NLKYRHXMSdjfNqPqQlzGRr/AjUimjTE5aRUnHZtU1e6idFHbFKq2fbGWx0F3Y1Vc
pbinYgdgYZwB53LAPz5AWCLcW/V1AFb/C9VErwm7Q2/EZ2gnQzt9UESAF6BLPy+g
UsdW0NtxXhX4cK+5DFECdpRArBe1RUK7lSamoM1njFnDCWD7GV2ob84sjHDTRv1K
79u5TloMlvVnYAbqUMFZUfhxCEHS90xVuYDdOu/oqeYigYcnw1xlMZtoRCsdMk//
PkHINzCb+qUKPc6Jj/sVMR/nfcJXtNanzAWPg00HMI9VSv6LYG0HhC6iPGhbnOhd
E5QOviI9O1wuRQ07MNbOksGcI9tUQoxddk9JyeltA4Qvpm8/qRfOEctgUhqacWW3
nXlMNGQNYWqvXqIVS8SxRubv/fyr9cQwr0grdsZLLZwFK0lxwD/dku/Pb53yhmqd
VuL5qxI3oWyH33BpXzqZqdWg+sTBR/WLtiDKXqS3LleNyKVTR1Fo4YgRGZUt60Ol
rSxY8wa7AQlKEcCItmCt35Y05y0U4pRGwWi+n5Pen/117AWp6FLf3YenzyUnvBUc
vIEZk/4Y68664Ct4MbN5GtSG27CKOb3998jHoctMF3iBQbCjlKBpYfo+pH0v4C4Y
R0+2sxRNNd9b5xplQBw2s1Nr7FYhwA94sbwgIZXj9yeLDeRoND73xz5uCkLsm92c
PKVmc0U5yflrmpSpUCI6qxAW3uIAQ3gp63qQko5kQr18e+KRy7xmPzmJNPUgpvgn
/s5wwskkJ6FROG+qCiBnT61z8sYe3KfHc+KFwpdLuvF/g0FCbu3rZxE1WLO81opL
7FeUYYb8hh5C3N3/VUJDLNHyVLb8wMFirACUZbNVvwd67uc1sZKfLSmgQMbuKaDd
ajBM4gBDzHk1tSRlT2ImeHYX2usHlVa9tWJ8jS39OU4h8gokacTW0sCKLjwvzKEZ
WpsQRpmuwuYSrvLsn8ZeK0ojfiEb2Nfpdij2QB6gk6J5GZOCWArkZd47g6HGSoEj
dPrnOfJZcxnBBplFE30x5kGhXZU/nZYxO8jlDXC5SOQeIfvfpnaSRe3sPZuOS8ny
7sUJSfsDmUCP2DumvUgIDHaANaGJ1jvICxkt9mrJ3iDZVzyWtI7X34xxalY30f+I
liYLULaitpKJZMHNSmkl8Iub/rLBVM0iggs1DhTRsI9wsIyy32hWJt7ZNw/8KlUj
0Z15r7AbecehBCYXcLa98C33nDxkWTPyfk4Aab0Y3QJH275ZDumfHO5rogIDHYrz
1gRHFji3MDNQchSMREwp/a6DkbgMFB3Kezk8ESjwdK56dqhrvxR5SIlb/ZGKGR0Z
VUj4YQnaxrFuRK+bTjw3Eynl197pmv4K8osSxtQ6Fx4W/6D+T9cgcyFolm+OQDyN
WmUPtkmhwNRxmkSpkzokSC6Vby7tMJa7rpUdi6z650QWi4y7XJO1y+rS3DYRosjB
MND/7sOdYhyPMWMC+6piOKXKIgMLKnj4QJwR9Uy9o6xxk7EdX/J7le7lxbbFJrP/
CQlbwlLZLxhGA/aFkoBGbsbKk1VQqwevwg2wsDlQWLrS/g2ccku749Vmd5M/thJE
JszI1Of846HklYYcWKxcpyhc8Psn7pYWSbenCyUbF24CLQhbQc2hUOTpCiEuIdF1
0QpJEAWpwKt/2+f+ZgBBoP2otxHuWy+zHBZ87NOHIPLSiP5no8lhhy3McP/r0Cci
R9VKzQinRTikDz+3gCCR1zDzGRg/X0yJUtDP1DCzmZNqEEXXkhDMepDknF21ntF8
ElBAexRIY7+cvBBRWZ307s0azlKbm0Sh6W70eArKBN8gTEAdPnvaoqTzO6V9g3ll
dZepfc6/4gCtgTIHmZNR3jNF+YOg4WtJ9fkeRbLpQF0m9UpMMuj6YjGCGzvCpFpL
4wtiU9InJC33mtSR5eO2DoQydY39zuGuId0L6DhpjVqGyk2m32ZIq6nA/feb26ub
8C7qxAaxBcGZNjpPO6GCOv6HmYjEU53Ddqh72nnOBTAdsXOneoHe/SsY/A0y5bqi
cBURuEcOorpExC1c/3c0t+PVQDVCEBN5fQxuWHV+Uj8vHdFHp8JKDrt3GmcPNxBF
yTyturREIymXLGV8k5pKb7nrjyH+Etheysjugl/dz1dEpUaipHZaH+9p4wAE7PY0
r94zcvo7ICwLyw7tSjPKkEMLv/si9rhaaVk9elv71hFGrwl4cHrgxFbolgpQ2L8P
qN9Vja4oL9G2l2tmE80UBylJhTUNYTS/DwrzUaBC2GspcKDffpzrtZ0PfVQ9suwR
Xzgoa3Wu3KjEkpPj2cpQ7K1MIQgLsvBT3mEPRmOU/I3807RP8rkD0u943yMocBuW
U+p90jksx7wr7+dRxLLe0MqS0BzDvsfJOjPdL0XGCiB2YVOQojcWcmpP53cMrqJ9
oQ9xMmCPqaGwE6Y1DBXFN6bUoeQWn4O4BX39H+VQYBoAUT2oMyl/WYHrgo1kbkHJ
KfOQbdQqRzvrYI3OP2K+jE3MTcCtNXBHxU3x+igam8tlGTiUZiHPvF8GcNrYJ4M5
ysBsbIvFlVs7UkOyFPdxHrQXAcVhEWQpmdU0GG2yY3EKgPZMLQcY+OZYwC33zhEq
k46PnB0Zm3fFpqXwy+Ee1lsGPfubRhWhT4Zv70RwzDpQGmeCQENHAUuMx4DlWoAC
vcKcduGnNiC5V8Zz4kIAXfUP1RkwtxmM7PWLaVOYWNtHVuf0Heb/zvzwzeWM9pbf
SAqWOxEdtD+pwjHvRL433mex/r2f8TsaaMbDg2OYym6KaPMSPpQO3MRbFZHteyO3
lbbHPLbxj+10MqSMeHzL05u6DxG1yNWgRIdHssXk6CJq7W73Fp4cJ6iGK6kLSfut
dM7GXtvQPajyyEDI7nVsPc3CNSV9OcQ+fM9ay2bqf6EgNECzpyATP5MO/aHu3N0+
3BW09sWpwqeoF1Kqk8yu2oBX92X9f8UukQTlEAMQbvD9nQgD+yjDfXUNX9LE4MjS
URVtEqx7eMrtfFKPb9uTWCuUjrXeBNT5lkO/N9OZAF3qeNc0QXdEFEyc8X0JpE5j
HzmyNobBkwKP2i8bsXamsmImByhGUgin9HF/FjGikBdJUmG+McbjBX0Dz0oz27kg
N3fp7u83kkP+ODRkKI8A6jRw4wRcfnQr0/hAOsnaKsecP+wMjvhQa4Xv+wo59yW9
DGBi7HgTL5XgpnzWSN5LrKuUhLciKZmRpdXx6dhyDRCfONnUI7o2wkUbWyWbK3bd
MQ3bXlY7V/tho8jVuFRTt/p77V8vlSFu5Ca+GM07CGORl9kFNmnym4/GecE5fcWt
5UNjA2s5zOHznNxa1mXS664ivaaMnIIQW0x5y/cWxWeYle0x+u7TmO0WPtrudho4
pQZJ410nj6XCXenAJMqGXPL2mUT2o7X0+zo2vdAz22SX7E06uTAbc2ilcUBHhnQ7
N5SDmZiA8bDQcIZJ8+e2ypgSiVz2jOlhAECLHS7maP2OkISsRDR9YB3CPYSl2FZn
/sEbZM9ZgfkN9jV4usFAduPDnOhCtWKXr8qYQuLsx2Lk6TsWr/nK+xHHKs1PHAzb
LGccrK9xF8CS6+1gfSu7hgSi92c4HzrBiyAzy2qzy3ZwSx60XjISXNjMJVNx/0OS
mTUVw06skeczOfNSb7xLS+m0rLKctBikmMFkRtGWPuWM/plC2yz3+cWE/rYhGqUR
cBCsgIWCkLXAAEiH30aDzz7xvJyCkhTCAzu6rnAgXj9pm+EGcNVyq4O24EQJI879
VyRLbLjbccvNM3chUMH/3AvxN8W6fd/dSrSBUX3z0MuEspzFIDKwguwVXBz1TNtD
ClUuwB5xK0Z4lnf7cQvcQpX0fWN/0HYLs4tyj6NyQL/d+5ed/ehPYQNBvBWWKTmn
Sg5Lq6hlIfG4HJ5cLdQlUDwaOWQ2D1+UJ+eTj+dMEyh7bs0hMFvcujiMF98xNQZo
kmTk9CWlL4iPLN6bEE9oaKulT9OnW252c74N5BtwneQlOFUaXtYXqDQVtkL4CoQ+
MeKa+6HtpAVxemXzKcX/Dx1eFSa2Jx1rWtGNPyT8r74rkiUKVGgzfS2AcecfhIcL
OrXMpxmIo3br7fvDxqZTslZdmSUr/i/oajRQzh80c0He9uLTK6Bc7X/Xiradl7up
zXbYjcG9yOkU3devR/e8T7HHsOPo9+m8I7yBg7ocGvWTajhGsM7xXuKlgcy/GDzi
UAyJQM3zW41uB84rBn9rDW8HXbn0gaU3MmU6AkCfrPyS5GTCFyJmoquvtTd8pvrt
JNDsUzVpAMllrO6Bdy9KmwlZRh/xRL+FdEnfc85LqX58U5Idk1NVIRhnCy+KQsYP
OL6wgWXHHWwdW2Kr8xivXSP1Svf8BvbhZ72Mj6f913g3NIVixAivVCOj7SIPjAA9
1lshk/yAEOcvFKMYISmq+V2ehMVYuyDWTVEZEKY6QYsi2tGUVxKQ21AbkP2APyoQ
sdwQLf1F5OPqJvU4T7JfYDG5k9ZEACPibjZr+XiFwrk0+4uT6GT4bdoUWAuIlpx9
SbF/L0QF1XvhDlXTwqjesP1sDoIejtwbhH1BlY5HlB1QvcGpwnRRIYWAhwJgCafm
cPyR12m++OAS4R9Dw4reY7c7BcYzWT3F7Pst1zcx1qCiCFiS3eHWTSLhb8pXawCD
66WKTixwEUeknR3yoBjg+rKVXUdw5F8iIn52191/FsAVT4iX/DlABioQiTRpH5dE
fYBM8lYwRbQi5pEsQeZZhN2gvNW0Reg61Sv2W6u0ICQ9/JaXaaJFEemiYUKv20M/
umQ2RpqQAQvyOX8BYijusLmYTrkTz/Hzo6TaQm1cX5ebM5MwJmY38aVLRfFqTYgW
oYSJKAW7NsNAbs41clSbLTvxAOD6l1Wq+mG4zNKosqSPoIdzO08CcrYJzGNqGmem
QHiv6VKPKrWU7+0te5NJMNlDZk9K4Ex4eMFeLOOFrSiLrxhF1NcYJtO8+bgDvcB5
YwpQ4sF+mD7Og7Ka0+sfqCGON5c8xvzbRGrotLSZtvU1xNDbVx564AmhcmDCEddQ
17uFBjWW7L2RkhLovxZM5PAeJ7XNY17UASZhN4Gk+xOkfT5RljL9tnDT6cliZjDx
1cc6WX0OFRJDe8w6QGWSFFt6+Rkilknw3lrpM5t029fo91s3pAPiYQMf8X+Uf8/9
/XkJc7DUMZdnpHyHfArFJKjbwX56O37qamtsjfrRtbroe5x5g+dHtOJ2ZrqOmGnf
aSx5c4EYoOc807DyJzjC03WUejInsldzEwFHnac1vz9RfI3t8iezNrpQnlHeqYq1
yTrlIdYIeFYDaY8l7tO71E3+WUB8L6iX0/AUptyPffwTDyH8Ww26vc98wOcuVul0
X3+n5BeqnUwVUU9mY9QL2e6NyHafexryUNU8zDTqvynige7+7OvskNeL2I7JKv7z
2bEJgPezEHevSmD6q0Uwb0FhTojjXUoCFLTZNi0W1IwPpUeflP6hHqEBxVIYrCf0
Rvj0NXRIFub1xeym2TzqDPKYW0lBV9WeXJ/xHc9OJRhrPhEaPp2qmkHZCeizNA7h
inrrlOdqrFTeQdp44IbBik8seo8at7209jCsVlNSJoHIRrwEEYSMFinq2HBL5Vep
T4VfR1ffAru9BqSSmQSUIqUpjJE4mj3zad0wnZuJivg+mOPbka+kTC2GiQB4lBm9
KIJXcas08ZtiBXU8GUuvHtp8pUtgITTwT9lQZ58pYAAHGmzr1ZUfgJS1FPhcwis5
8jXRhEW1bb5bSJvaB/fJ4ZyqwOv2VkBNva4spG6myFd+weUltX6kxAynbzXfDMeX
FaxJyue3rLu5aWTPXAW4/+1UZlJX+FghHbTYP5Du17KNQSsueiXW+L3Oe4gnXqpG
+Uo0MFC+t/pfMARCvl2KqtLxbocT15c3X9a0p+FGjOS2pqgSiUQnHOOL3sq0TfD/
yqwHkjcP+PKu/tZr6jjHNo8TmFvWIhgsyu9c/tVSXnLcPTlANuRlIbcJnJvb3iU+
DSFZJUDqdLirOgMT0iL2m6Wz5EYx2gMlOoCvZH27RTCfU/towtk0rMmOpJLlkJ57
zs2kwVn3+1U4JEmaIzj1yyDBm4LNdc8eUwz8sPH5ejksIk7dKdTFC4ZmGIApipcI
q76u+VAI41iJ/J6jEKWBU9FY7mjX3i12MVnsP9r12D8DTpHarfJgWhobw5ntTJbr
vq2sjW+tD39y7CDmHfBkluzW7MghurRrNYrYTF8c90vb61GXGc4Vo8Ug2hhAhrjO
+IzWks4oz0D3j2ogFJmrRNJ7cG71lXy4bXzh7TquT18TmJu7H99UmMh1ivPrKes/
OgJgyIere3RSk9bYrdsuq1EXFpPZgc24QCt3VBczarcG0yCHH6OY6iA3MmkJ6vpA
TknhULw0lPDu0IoBpeXM/M2SyBHgjXEqLSeGF5WiML3IsKxnTPkCWNVVej4zqA1w
0SmnvHtiRbig8grhUyrjs1rLJh/thOktnG7swR8FOhXRusq5uYLErNilFG+BXZbz
RsYpsMwUTb7MOYGUkHCriUSxCyY+zT+wMorFYVvUPNKd+ZlsHifzyuRxIHjpic9b
MM0TF3P3OSUSv8wsXc/hXfCXqPWg2PwSuTTsirbLeLUWx3nqRCm2yno5SUsTozqC
0QELv/Smr+5BXSL342kk7j/zdAoSdBTnp78AVLMhLlSVlxNx5vo8rpXbLjsSdDnh
pmz25mDWluj80B8tZg69RoHv3L1qMb+R0vwI3lQuatdjHFXpIJ5hWd55p3+OSxmP
VdqjNcomVxWsaZ1zPDcvFyu92dURBXm7a9s0G7HL0z9kAl5cyqizDQTqw7Jg/h29
iEzkcUbDsw3RDBQakSSdQ3LWWJrLSZU5CMeAROpGnyJwEmPbToPSZiyTS1u/YaBL
RfqJVRQGzVmm6nefwvLRG5eNHU4K4ox4sjlprSqwMd/GCECk2EYmAOo0UaHSSyfw
S0ndkB5pkgLXhwgmS2tNA+SWOU69pAtDaoEavgdzI1F/b+zFYxQtETUHuh0vG008
o/p96TOLrdUmrsmd+gBHYo6w/Aq8Sttf8EZnsxajyfZ7c0gh8akkXdZehfnTcIvj
XLgKxW9YIW8O/KVIsNS+lAMNt0CFnJ8wIT2Tls0jqzBNnh2j0ah01nv3kikASRkK
F52VE6/ARnafoja6QQDqU3gM+IQn4vzZM2vrysb3XzENtxlzodAeGVUiCyPoTxHF
AvPjlnBkNH9aRxsJvKZjywr1q3o+W8353Uo6ZxGRyWzGD8CP/IfcETduxwTReL+f
Wfuq59WpG2Y9WHPepwZ+AsmqPMr9FATUICwvxSL+fu63Ti5pef5HAZ134OiQQL3Q
OB1mBCvPDt4ZuwS1Ay61YOdA/+B9lkR/ZWzVItU20//vIlt6Ui9BOu3yKY8cNpDl
7jZ4bz4afiQVqK6wDYIbqVm4MmV6qZTI1j7EGpOQqPZwFncWXttObLUtlmeixX9G
Kx5KiCxy0uEvUAIt0vmqIlW2WXaClMsFmw5SS9PKrUE4KesySy/hHH2gooIEkA3f
ZRFWehy43x33svkkPoDFq1RgR5Xo0wTsZj0DMnCo35GTWXkOzlm+731E1I6A1IhC
cf8+bPcFVHyTQvdk2GqoqwSso9fTmUlMW+sXXBjCNRhUjDjRm+WURDIJZM4cNqzd
Evv38qDUb4zB5LhPO3lh2CC9+A8XVQpb69EDCQojL3V1OHPjpmmGAsg8x1ukXNDH
bRtBmUcRevLR5LJhWjnxcwMTpBfTlAQo3GLNz1Ln7yhDwl1tEkEccZpprRLNNIxF
QW5+B/mGdf19hB0UfvON3YPisn+6ztFcPmLYHHFVVUsBhXggZTNOtIU0WFnYgN/x
s4Z19EfodBkq31Jpms+cH2iKBktWthhXG+xtkt7AeEN4+6QAYQDW79iy00IXkdEa
W0s6rh+nFxD3Lg20JCLy+6Hu6rX3txURogbPeZX/1EbVhZBV/OsXtT6XlYF7CUyn
gVKr2tuqIRdmyUluT8Ws96gsf6qceoZMhKtonNUwreXFFiq5KxOjBmyhsZw+aKv2
RhIWW5OUCGmO8vsj/0XFqUvmYlFFrKAO1Gj3y+ojfHKtKLbisOFpSGzlnbSm0V28
Sdurn+3wwQ8QA9gQZmyD7LYJgU7bX1K+pRbCHWfhdzfdmJJdeWvVONLHf8HVcaZy
2sDPwRQ3oU4di9pYLe4ZZaFjShKa/6C/fGSob+2gN4ARs+Y4x+CbOVxl+Z81AkXd
35REnwtrCVlmKA4rqHWRqtP2kGSx0+0wYRYmQgjnReyBOQPPIlfcINYCg6MV+qc+
eL5djbf9hSmFavdD3X6cBKam3+h3IpyBCMeiyF33ZzF+xxDuVuWPkYt5YUnrPV+5
PfMyOc6LLLeJ3JHPZdMchQH/rXCCEft1/5nps1YpcP8d1IzsnA1Bf5JSGXRp4HeI
abEZbquNtxdcoR2H7fsu8cmTAjyscw5ROFgsbk1tuJH5nX7/JA6HPDoYjt5UqYTP
33HLleP8uyiRcZlyTUaYlPMfxbSbvKsZ5ml2YcDs4ozJ/JbecaDwu5r4Z8Zr5Vtf
wDMdyJvhapGAHSRLgivo/VE+0FmeoGTRSgxr5zlkWtlBfwXQiR54OkkOX1xH8Anp
6+TVQXQAZTrMrO5yq/OP2VnVMp8DvDhHeW86kheA8fK34xjhk3W4cxW1a8HcZudc
O/WcxxxFeN7/6QXSDsSQQ1Vb55PxfGbybrOZbBR9UPBZw6H4o7g8SaUO4nfmdGq3
2sMuaBJtD1wHZB+0L+Y5csk2yo16Xc0j4bwNhfzfB6ZkcmNrtp/x4VSFnm6ocYtY
OxyP+E6v22qntE8F3pm3vHn0LJ27X8atI211XcF6SDXD8/L/mXo6381Ts/6BSMHt
hXnEWSAuX0qeEVG0ydW6cv0ur+XgNf3BrnZSbxo5wA1f/ZMFRH2Di36BCRxMXZMB
IkON9bhnEyD6+7/W5OefNKU7nFUxlbICobfcufva04BhAKaauwXoe220oURuSMnm
iiP6ajMVVqJ7oXO0zDpoYIb9DrgxWNjDCED0SFGrFL6ibJL7cmDnForOyS9H5w2O
/3EBa+aDo/ikcGSFPiOxSqv1sR/qmYnqliEnhcvMbuo16TIVUZmc/nhaA1+J87aQ
lWIv08gZmomKHJ5qo7o2dUORq/upmncy9Jo8/rVsIaXHk1dc0fzhAmB9Hf/y38M5
MJpEUgayi97np6BgseAT6y7KjxsLgvRc9kWpwy+4gAR/jHtU36PUIdDOUB6c5xx3
Is75C3h8UtI6UEKDT8hYHgliIY5nV6Blu+y7z+MLINivX6ZtCRmE4LpacGBji6TN
1lfBr1F/RH4NIDduqfFEcurC7VwiffGenphjPqNT7fOGRSDHJ07bV4ziWHlUMBy7
9Ij+kvHD2wyUrWTLTFDmoKqKFS0TDyTkwwJeYiL0iXALLYZx1zGs6UIUDg/ZS3nX
v5nICU2wAOQgt1QJAOH425m4fRCyUONR1AV+7bfy5WxZBz4Q2U0yRBzPxS0kRSu8
4YaZxlvzVfxwxsigK2lP0RXPpz8vcDGHR9Hl7hC5y5ThDyKMuduF8vKhVyT3vzSZ
Z5ynl7WPGzLF7SJTWW40XV9mswsvkJNpOh+cyZWCu6uObvrEBRF3mpTLk4SmMAho
GxdpNkjAyCCZykAz9Hi1OOKgHJ8IqShEr1iVvd6+uWWrglwLHrI2nGklkkl7s1kv
zPMC10JFI+NiVgYS9KzZOQuMIdZ0Bzm5x4POZ79Nb3ZR6rcnkZ6pMwuPhT+WydMT
+Ekl2nkyrjF6yFg0IWk0hsfJeIUKNc7yhpvGaosU6eDKF1ViJO9QB3ToVoCEaZyo
GZBao0uqm2dmph1D5+VK7UEICpXjr2+xuQowM0wouxltGwG5BbX82YZ76Bk42f1K
4NN4stYnlhSnrdSmYKRmz6lxQKgfoHj36UaDh+ahoKsAiK9BBJdGpDUR2OZYt4FI
S2LVR+es+ql0qeOCTh1rvjW3OmiYhIFzwxUchTkeJDdOtUbpoRd++z2EpQ1l41A5
JNyy7xCVSq5fIDlwto9zf6iLq5Ic00FcoAhgoxygsB92aZxqK3GkRf4fIynSdyzg
SgB4lQdZxY0NeNrx+qq4jkSVvs+SxpS2BPt7jsuzD/XFW2MuJOSC1xBOS4EKEibG
2+RFtPaOei+zYiYAmw3pFK0HA1D4/bK9Uwq+qHYXsqMqqywAS7bvdn3k+Jg4/cOD
53gNk4m1QsU+Rc0I5cJYnqOyIkpNFVzK2N6wNZ8nwj9FtdJRbUKCIB7Wsuci5TEu
G+F9thQ38wgwTXHhXY7tzxY+LcF/V5FihV4rHJFmCiFMDkJzKiun1DdYpB2qCzvf
sfldvat2/eohx0l4qgZAS46MOXJpbCkzw/Z3D/jjYnOTB2eyv/bgRDFHhf3DVY8A
1eww8jEXfwEhALZVYPA//Bk4/+FlOxZVMrZAGTh4pELiRKX3Nx1elttcA7MWlu3Q
ZUpmojvbQ98DpPS3lAq7fKFa8LsJnXVKLMOPMRbRbwpo/9oToTck4GsdUnoFBSZc
mZDWFdNtoiAuiqJyx9MJaGdkAa+WQGhUHgp/2pxi3EWL/JwNFAncVlIgugxMn13K
e9OVNGNp/h3h4Nzpi3j+Z+kTouyvClB3myLxStHSEP5apAyoLpDdhNoazdbcHTYY
nbQrmATRiC6Uh50NixIMdCAGo+xYATzt3kZUTBB4YAWDxGeKaEAM0vWH137MM1pR
IFA4fZtZGy+NoUgup1Z3an5j41WoEt3kP/4A/PKmH4bB2BEPp4gR3vRlgyRE12Wq
HDdwvkF8TucRhYjMlQ8dDvkN2E1Pq+xB7DuoQET4dO+uAVPB1ra9sTFLKalq3dk+
DI8LZ3LkZ8PhE6vvV+O6CkIi8pf06tnCLxa6TXCOyF2lEA1Nwg4yzpDI45Ssb0eT
PxfIJE92VxP9HwkgjcNcQ4hr9X8vg35NNvB604xyC7JJvj2MeNk6z3iflwBNgFar
KLpknybiT6e0lsjI5g6PQBLDvItrmtZrNwOM6+Cb/SF4j2waBlwk0vdFR9XWAgzy
zVBomHgK/vZfELJQKBwltOifjuo7eHBdyrNMAzyr4hP1xYtF/QSVJOGaBB9qRiJf
ptiG73q+P2z1raz5Pf6MOVX1fboo8/LCu5E85LXtYKuPkdvVlSLL93GrseUwwiDn
nmWQGXsiWSgpJqxVZi8k5pRCT400JxBfBHE6NQy4zM6t+OlZVPt7sOoyKqPy0Y+G
6q/H+Dur41gW9/w8xK+NiZSUu/il6fG0/G6H9Fni4g+BDb4fYXpwEZ6U0GozOKBn
N4r39kHwYKm8nNSxdlb5yim/W1LguWd2SzYBBXgyIMWqME2zsyx1ewZ1i5xrB35Q
ebyb5aIvFMPWQ1inG2kl7HyhqmDxvSGEHStiDQjLSPxgSE5/5Xh1n5kPdrUOrJnU
biri5v1VLUYW3Om9RVqiaEh5skyAukqfdw6YSu8sLgpF7WK6DK2fCBDRxuxhhQWq
DBJgV3pj09HzGnEe6i6VlzOFZLlzw+49sOt1PTRUrYpp4NSQhfnH0NLvdos1Iz29
Xo4mTP7zegBuyJ6tadRImXtFVpS0VElNvggJ6qwqxisiyhLSqPK7w33dA+lNykCP
iMfPdxAApwU20fETp2wDNwCvSY9EOytwC+mCsvntnzbCRGpFMeZPLduYs6d62l+m
GUwp503EVgS+sS0hK4PWdYJKOLi7TnzQfFFUOstmmEHVGFK33rJ9IJB+Tt4JcWhe
xXuhZAQHQgo8cTmJPRpRRCTyX8IGsagVMr1wZcc3c5vpNFdlGwDjiDacm9snUM3o
oUJj86O9Zeo/veORbHJkeCRVL98eke5CxFae2r7W0evMNXWGLEyQ8yLeuW2zDuSD
5/DA/Uj8+VGY1/CQWwICd7SeQ75jpZ2ga3ytBNgf5If0md/kBHsucN11nyQCc9AF
gM7qCQq435FObJk77bOpIdb59nO4yLsoQJ5iUe059GKuI7t7CNTNTt46OTgwEniu
wcNwYrpuLxybUZGwm7QTan2FkhOYZsH+MgQ+O5S3t6RCpDEVghK1m6flL+p7KjnW
GRv1jIQ64opYtI+Dx6MbIIH9XHpR0JIQ2Z6GPxI9nCmNtRjZWaTkl1xUFzbttMak
uHnjoY+sgNF1uKpXJZfWrsZ+Euit30T5+KKMtjbuhB85cAMyFFrl0CGPUGhL+AZL
uOAuSN08CtEbscn2K6944jMfYl5N789Uvow9ouSiJ09EffyC17DFvUlgYFqCVMvK
gMDv7ZSGzbzTH2JHQp9oME+uNIm+Dv5AE9m7TgWkYXUXxNSoQdHjzeXuU3r1tC1H
S+Fuh06QZJxYz1k+tAwdPYL7OHdEbs+XjW0Aie1BXlYmkR/H/4iSw4fw1c4kvH6a
Xjid+kz6N0a8pkq8lf2+Ji5ltMr7BaYI/584WSpIoA7/iO3A27pR7AMFG5sQy61k
oTOWw9qoCFiuU1Y6KPRj3/ZLg7XU/tKhq3uZchT2cskh6meUA21oZbhOLNK5mEsW
m+v/hS9afeaTUxYpKB1hHD7OjzghyAZ/2mIr0KRvQU5sDr6scpvy5SPMqwBx3zW0
gWC2U7cwAo8UysQzjupP2gOL3jkM81fzhYMjV0b6v3BWKCiVrTWKov9+oRH+V80E
yITiVZB6sqVyDLVFBGnL8Vq7wa3a6DfMgu8gKrzHV2IGpja1xWHYPt+1oepy0FXB
C4VF98yN+QgawVYuyhTVH2l5AlauxdUHSBVBTYSfRpSTaVmFzPlUA/QgLgAnpFLk
T3ihLbzAuNRJCw99UeuPxm2EonJ0CW6kVZ1MnFNIzaOIDaH1Qo1/LOV0LOihcOPS
ajFA9/NLSlx8oHVDgxuFnpwWfBKY1zEfnnQeAaVgCL+RvE9C9TzYpglxaz2vOXhX
yCi0mp+thhkyhrwDYhfUKpLNjrFNryXMmmRsQEgXiZnzPLgh1/MCrv016P1BtRWR
L6XVsYeyvP7K2s8DpI6lYX2wGk8vELqjGh7/7oMFO+mgTgMrg/8IUWOj1XaHxmAG
BUPJf5jDAmMFJvoXx0MAq6Yl96uR798Q2M6seGFvUEluWE6oMBviIHGF5rAMkHcw
BKn0T3oUoo7RjtCUgJr4zvDkihpy9kObiSxBG9oYCs+JlvGCRbKWtpkj1tm+bBaO
/yko+6QxF+hKm9lievSGKJAwThXdCZa9+SY0Er8uVDJd0Db/KUjmsudSNDP5QxEo
it6R0UEJDggN528BFEYfPlxrm2abgPaBRsbLsLnPAhfycJsmJS38RadiFaPtPwsM
Jj2sHPI0Ik6EDW7TS6xHsruikRLWaq6KaFORQoiOhQYsdnb2ilE+wD7LiRl8kZdE
RMjgk6/ilxXCFRXpDaiJyEuBScmw2fGQhn/wZepWEPEgDNrp6eywK54vVbYURj+5
FDrXP3gQKSitu/9uois7u2qQD8Rqdsje6081H4/sCNKsM3kxtwLmYv9K9BNEUtM+
orXW+QGThGpT5KulTt9w/YqiiSuZUc0JIfQ03tMDgXI/9sntFUYXUHUqmr8q+8xz
iFCvJm1bbjh79ep+3EjiFMjWPmRUSTv52IxOe9bM7A6YL/1VxSc4S5ZTcuTu5AQF
RuexqIgfasi7DI8N9iZOu/sXo5P2okjuAxjJDy5IDF4fF7brUaXaAuZzfGfwmRVe
l32rH2nZUQm1smjoDMtL2XJG2phCLhuZYOht2SrphmTY+AZDUyxIkriQ7HMjmYdv
DS4E3/NPezJW43O7U+w1Vp4IhEWJWYPGfc1TXH2wvxK4p5EQXf0dDq8YSxd4N2eS
x1Mrid4BaKI6MTDAvHI6PZ1nIwABPrOwJHZd2Y4nhA8wCr1D7Ljo7Eh360HXLKO9
Xmets6CtIhR3CyusGwho8qD8JgrIedAkn/rBuN95OHUaksoxbhp9rRWo4WRrewmP
ilL7HyBj/yW4e+R8ckq7DYy0BAPh4ul0jOFFTYc9fNEekp6VAtEjGq62PHpd042/
vLzjGRB//Cv3YNhZbauW+A2ChkOqkq6ISvndJhGxQdkmszfHMJTi1rTdyYRby5zI
OTQ3qqLFcOceBH3YJvF35qVB2Lwl7yqt+Qt2GPVyBYYodZiXSzfHDBHtx0Jtzx43
ZHScsN7+wHTzUU1v7U3Bgpy5MagbE1vFzu0bKQA9Xh7IWI9qUdQv9TMO4CVgjZst
T0BqphVqc+JWzv/uue7MTziYeT0R7a1LiMmBI0s4f23WkjMeSfYuSA37umItUBFm
6axJLUffqbMKm3laLMRSoapehBMvktGX/+3TJFS+FS2o+6mMrWxX4RxBYBrGcA4H
Sed0w1KIQK4MTdaW5p72EO5wWFh0hBcCioJKWqyZ4d6qTj1EDJN+lS6JoXZOAESO
I+FBRteCl/aqv1+cQ/n+VDtVkhZ0SgP+eWX76ZHkiSEiktn3+m9cjNPP01PSTR6l
y7SnToBm7NcKHKiK0hbDwGCRdXZpkrP5TRpEZgu7OZyxBN351+zRlG18Wha5jIJQ
c+5u2c3G8xaIXcl/M9QYbWMXIoc05sRMbkFMsorKGQkFPBKbN4DJkYxlYIyFngib
i2oXeNPd1kfHDsWLjM5G0uvRs6fxomgsfzpC6lpIXjOGj9Kutgugq0TM3qKcEqdV
nd4acWkD1WUueX+o/8tk+E7lN8yIwsfssNXbC6JfQxtOi4ZDF4HAFUldLzs5kobJ
e/GTtBUNbBNomufmnILEIK8V1FbZRZtZMI1XoTwG6o47Zq37xkqwuEk8N++YCYSE
0bdmDREHHgfGHD6nw5dUHAysQDWkuCy45FvSY7r+SBi74cWyNmGTKYoKSXjwIU9p
+VdR/2DdUZgc/r1XfiM0gPoRJoBv0GuOU7zZzdb7RyZaWwjDesm5fYpeJC7yPIH5
gSMcFbJOdPGzhdfvYbpq6IR3/go6sUvVWu/G1UuHT7TZvjhPZvd69ABiZcEplbqa
COEAstXiKixenEA8nEFi/q5bhOmfUiHi4xFqMZeYuPQMD7M0OXPKg/0j5cJAe0U+
r4OUHSm5//TKBXYF8+ftIM0TEv5zH6+BPetwhTQKR8RLjZeI+K0me8F435lAbZDz
7ckvoPYT610aOo8+DNj/LOxaRqvPL2XbN742GmcYGG5rolts/rptmJVbed4LfL0w
Jv/q5oP0KGcwPx9MafEstYeCV3oIo6d7IQeOLsVbOgZ/Om/0n8RU82JmAH7GwZmZ
iK0gKCAH20DHVfBAIeWuk+8nL4Q+GdYgXHInBmnaAn+gfO756cxj6H3rTKoFIjzU
QduFNSG1JSXummL6AUuLVUL4Ze5Y7s7K6a09+185Aog4jxHw2dNxqryqbDW03jb7
JFUyAnqATJa5UPsPviNsadmQ83HeW6ViTKbJElsMO6rNYQ65jxuXWINMl+YbEQFq
4Fz21yBBByxF7FzYcDedUGVKJmyrpo+rrbdIDpFgUX0T+nPH0RrvDPx2UB8IIbna
Vv5Fj0//KFc+/chR/RH0TGnLSPwlpRwB75xiQhJbD+04rGAqJwFhsQePaw1vhUd+
lKUEZAVBxFqx2HsjUY+Ybl+DwCugyII0joLyZLNavIAdGLbUCZhCaoy2B/lrnJ8I
4GOxOkveRVXW2obcGa4NAB2GE7srvJkObRFWgL57ihJFauwxc3qkkz0tK6FdO8Ik
smZ1+L5N6ATp2SqJqP4YnsRqm+nbEzcCPt2O15oqHVac0khuy4/h/GAmqN8gVFFF
x9M+xMSfpWpNNkZkofbCOXAxRPXLGEvZ1dLx+fgcgmSNbJT/LuLh0RgdYRkB4e/b
OX3lo4LeIoG3bCSikCHpIVdRq6etBiCaLTMH2cB5HPLOIjhzj7QP7UnOfM3hpgqE
nfciDqb1hBHmps9OX3BtA4b9Sa0SM4S9frC380JafgPCPNpCZGiXtJ61UXEpWWza
dWhaHZCYcqQa+pIKrLXH2oNDB00Tga9EEuDMRTYYvYSS04SfYB0Xj1yDCm2tip+j
9HlDIKeH8sWcw7x3JsyDG9ZJnniRo0Vvstbc++1VAhjPa54XMCrq051v6IkqdsLl
ukKDG/d0zqVqyxxulR0H4D68SWHJT8Wjyl0dM59F/T2+hnoyZRii8EOCj1Xzx+mB
WeQQngcczEzgwz3IFBGtCDeWNWc6Fayn6gQN0Tm7AUOsdhVG6vbWiJwUwVfyFcqP
iJERmu5ee5EdEui3Njk87t3LNcYstLxLmz2BHzoA4vIx56w4k+Iq5xDzFH1eR3lj
g26NQ0rB0zG7JNJ6Njf4kWy7jTIHiPDdOJzYcOC5BvcFTSrR3Z+8ja5fNyMVRSMg
ffT3u0t7pNhTtNXO638+ONKOG2P3UdUeWj5Ne6ByM/bgbDUolFL4zeh1uv2sZcYG
VyafUZVvwRHrFQv5iE7P34asKwQPQjEGLbvjt9TEZcmI5lXrIJwHgZjmtSymShyR
bvYj+1OMrz1Q2lQKCSPANglBp+Ra1Qa5KawN8Hdt2s/2yAhxmyylO69v20WaPHyh
2X4iaZNVCLgZbUsEHMEBp9u5fI/Hv829HbftwMYrCypDI/uRg77PTd6B4wwdYlfx
ksKvisuS1vz+IV1YkV65QjHbf6LJ0GVw7fkUBYyODaiv4zvW5xSK+so6oMIMOXSx
WTfp/K6I4mPTY0laiwuQKDbEE7ruwJe/ASDSlNMqX+WrIZTFw3ApFVBW0DfjR3ct
vIfeYrmjC6HfSwBTH8/FFmorXgKsiqeFIXToApOEOHmKCWoqZzVdNZ0B95gBCXvG
YMGdVFcFGhzzjmSDYL48J2cDuVhRdV+XIkbjh2P7BqbVhOpvLxu9bDozrqWv7dts
UzCDkekrKOC4XCp55vSqt4yrqC4lyxXGL7m9OI/B7v9UaWAWqDuthPxFEmWSZ7cd
PpyqtQLxwtKzzaOEYJ8I1o43be2tABMW0HqcwHwJD7nhWYTA3YGWHRfYo3BwS3G4
a+DjuSXCtN9EFiCe/ld8POFhGRF/PhbtQftad8pFTpOp6YdqpIP5wYq7uWM8sMGu
fXhs2BQ1NX6NI8EM0rkgZE8WsX0UZvLqUyzBFe0o2kGjrheCA8rikg1AFpyaiz10
g2o0x3ADaswOhDztJw81QvwG5whgLI6VMOZMMgwrnplpFq7spRP8rjaHV88PN5kL
Zulfzzkxrvd7MqllCEFynfFPFnF3S4M2ZE7JrmSaNK3ZQ+DtI5MEH2R4WtZwuvb0
CMshfxe7/qK1y06n7QhbV/zrwvKyZpNwyyziLVMVGtx5dWEWhg6zlMmpVzxmZpPC
aHBSIgLt7/cXm1zz/RYefHw3tu7QxBdi8DFqCGod6slwuENsv649OhpuNfUVYnIf
99uTDcTzDLAKSM+T46sStjfNPSOvOJf9X7HuxTBo3NQYKihmc+1TSDYvMXlChS7M
8TdKFZktZK5DCJm8LBwYIl3c0UWTW6Fy0t/uJ4MeNPlgOqIm36dLDVz32jdLQFlf
/yC/wHdu4HCjJBQ8SzXXGgPCpHIDuNAsiSEYYu/eqo352I73jGZPMr9BNwQKcErG
e3q2iyesWeX2Wv2oRzuU3JVNwiSyzAwPN7Fc6PAFgDjWN/E1m0NIWK+tuzXw1JRa
q6EVTfed6HT7Jq0SLG1meHsiRAbGYeaq93CqCTWUHL/VzchejwQ4jR0LDnC7xLXA
gkAnRXeQ/cwFmb519PNe9ZI4NodI8kA/tbB0fhAFWOxNAPhYB8t0S2r4deKOrXSx
UQdNNfy1XdlAMwwgB7bxUNWoBkGNkWTCmEvGLNNH+lKze+EythwzIfJeDiyWkhXN
B0KdGXcjqjqZM1nzuK3lBFBUbUliAsvPJ6cGWy2+ahm1LIOwBAcOk9+tAaN08gbB
n9oQHHGZTMsdyDQ5glkhlwDj/j8oU5fUQduGP2liAVDPxyD4yndvdrdF6OQwlaIz
DpAYujhrnqbQCV8rokTbYuXLKIVCJpRN+DahC8yHJ8lJlVYGnWrYHk6OK7nN+1eW
C21YRVggGh9Axb85Wg2I+im0BjXa9FlB42362otYJI/atOR1gNf/HrmsB8rUYo8f
E7mxD2kdDt4QPpjgr/WqEbacugcfUkdVNkDHuK3rjnA5ndRRRu95CbC1YUw126xA
w6e3c8f1zagnGpT59//btnbZXa/SUX5q/sag6Gsrt8FBbiY3tj+D9W101CWSyE3v
umLDTUQ7mN3SGH7CX+ineRQXjOP710oequetpjZ1/osguNeKePoTWnVpG++RtmFX
ZYcOFmy0cJeLOrrszPdj2svso9B9Hl53a59dm8OHamzk9gWkvRALeCMr6Cw+/Lzp
/nvcXVab/LM6SAsHfP1C5ptgIhj6/OXX1OMEMtvblTpwYzBnDqy1Wz2+O2DIHVqk
xx5Bu53F+5GnnefCgChv4ettVGTnO1Az9HeoJrN8kuyM0c4IVl+E91pa0YezFIWq
EYRfoYgseexYv3d8KbKcjRADOyJE+ukGsq7assaAdAtnD+TnS55VFjRftPy7OCJq
SAYPYc5RmNC7U8HTaTIoQbfeauT/JcXuV95lxoadPeFaYnLJTM2mBuJOVlGMGIXJ
QEo6DC/8PU1tXleGcBL9J7GW49Y5HXxfytc+hUswXczMjBO++zNR/iq6dg6I5iX9
UtZcJtj6WazHKsBORiDFnq/3fJKc0rkLlPuJ9nnCvyEtjYxku3Uz2RxCbl/fnKww
CPlZCQbzPth+T7z1IqHjKic12YpXSxcsrJdNLNq4pdURTleR2iyFTtyAi7wb2tPv
CHue0+JkHUOaYSxpnhfXeDawzr43LFwqP9+tPrsp1TX2He4ev/YlRk30XO7oo9XP
Juo45jwAL8gsZwhUt64HCCC3ruZNWx57CNKgPux0JS9gxWt7oRAwqkSuxP1mmYun
dxE7rIChMXJziibj8F+YByAWZvRLkcrzUGgJFCp5XAmXsuVw13dDlNB7ni+xzkXj
hOpmBXIbZxn2QaqvK+VvgqC9QzkcrmpqiahkrzwNh611NxhritjcGj2qpc7EZ1lH
6PZz0j5VQzkiRPDfctNkmZQhkrVhvJuBubaVIH9rXmhPItSddy4mgGKaQhNYovtx
g4O1Yy6JiIlfDPK1tnLi7wQoqrRbCuK7/iekZFNob7Qk8A+annYUaYWdzxzx0mNy
5mNfWmpyX9F9PdeuiaemqaeK7hGIwSlgoZ330T3+da+bVAOp+Sr9U4FmSnxFJ26Y
j9AQf101KPR8fYq1QldSyS64P63+4trUS2exvJ9fDsWG0mEaoQbzsDd1pPMry9cx
DYfFXmrPYGK2M/WGOd2IXevan4zoWHisFi3VmFoVLUpzN2qcVYl0JHFbydh89akv
H0HIGP+eb0eV7LluazXXH/5cjn5Xu4OpCHj0OPimdXqjVwUBBpc2xtFIdpQk+UhU
Vn1xFF0TDtmbsAu5OrGG3ylSDrBdTgggCiqguENs6vAEYNDS74QwgZiQx4bx+Q2Q
XgvV+HgVmeQAJ8SUQ++PBjz/lV9BQSSmE7lTq3qBqiNY/7PkmfjYB4F/UuLN3PUb
i6ypHngdHC502vzZKp3jpkIIut6nDKYj4HBfvBFfaGcBmAvCJvUrnuipHhrhgsxN
hq6OVzkvU06TfA61SROEMYXyc9R7/fVgnWB96cdsCRZbdR27TfI1nmt8eg36Bl23
LU0U4E8tuHO9W5m5tINj1pS65RDJ5WEK0jGY0d2zqX8w4gUufnqwk2tPgsR/Oa2q
vbeHUWLR6gAqhwwbOEGjh5quzRHuY7XCKsyBlwZWTs8wEZiXqBC8YRSPQ49E300L
W3veG6V3aIeyQw4ZSniS7DFLJTjQ6r9ra/m9M+T/RurSIU1oqQ+WY9swdvcVZG4f
j/UGNIWvZP0gw30HhFZPS2+FUhRmyTq4Z0eQTqEfrmcxuBWKvBNGg5Hd7Ne4mg7P
o+1BigJpTmBDzG0B1IUWwWaPrVulK0Cwz6GlyTCzlnf0mn7lci9nLkMSq7eM/XDP
zCcIi0/H/UgvH6/iOk7k3ecppY2NRH+Y8GCClahieS4L1JDjwpCICFu7mXK2pswt
2pbJ+xXmNskuFijBxpcz+vc3BAUzoS98d+X1jx41zpzDAKcagGjvWu6RveX1qUpi
mTs7SZSwKaiAUccAm2BRqjZN1FEC8/7RUeWDumo32aiSB+6KHn0RlAn24zf7xLzP
ZgSbPd2FJUAzOI5UB+Y1MpDizwH6ImO4f5stlTCZA2i/41vjRG/p5BTSb8pzYhy5
FtIaed1jwPrka8YONBaE0Ogr2sQhJ4sLAa6s/L+fcOt5Ur1aQxLwZrFnpP0I75fH
fxzpHBXah1A58hxixicA7RRZC5UQCVkJEDm83bSNtAN1OFWGyzwru9w6duL9DGBV
zUEiBPkq2tuCuvkQ5E5byz5qDp9Vd5FBA8wVX7IFZi2uOmp7Cn7zNpFUvQR8lwKE
btwgeDuTAZQiPeW52cGG0p6cu+jwzPuOrzBnc+V6g2goSECp01NkxJf1rlKqtvv1
MuBpU1SNyTGNNE+FyY5Nea2GA38o4wJs/kYDsP+t0Z8BHutZucsle3R4A2a06B4l
VcvxVR4mTmd/kXZUsV2LJNTH4G6YIL+EdouSkjIEZTb8+jdtwhf7lqWcD9dCmoZr
wulsmJzI3S7dyPOyrvQ2t1hfK+iQVD/7NFvftdr+s0nyaBQzOMiQ1wjoOPai8aS9
NggnIJzKLQqFHqxXfqwjLIlC2l4IuLc0oHaIw3ZGlmw20WQR3JKkH2r5fIRpYjp3
6Sa27A9a7fPCOE6W+twbOIRKwd57HjgiloPbuyCoM0uCGUxUGrXfbsnlhCAtdLaT
uEtPymg39DpKZSzDUe5bqmJqmKsrRh/eHRQMZceYHnr+ZzsSOq4+thUpcp3U4eJj
3lvBw++XTjGi43HdHI858OTvJol2j5YjwPACBdn3Z9vL4voztaI0CejTmenhPc90
nvSxjAc9NnW4JkIh9nLOV8vgaOMqv1G6uJa3o73qywV3TfKTdR+IH8kpE2/TMb2l
kwMkk7eYmIyC9/aeJ5gR3NIw16S+788st1ZSH/8dfVLQGwNhQEa3NoAk54aB3H0F
9lSpHe02uuwcsnPgzYBR9PydOTAJVOIP0K4CloPlUJ8qFoBiJxLRGrtOZvTFjYbh
Nx396p8+r5mo2tgF9UKnqY35tykHMgZ+jwlRnUyXbSjMjcljlkH3iSFqabMYWvzo
ejqd0uSzbthqxkX2g1TL1b5Uj6xIeNqdjgStFi/Ly4haDiv4sEEicbR1eamUoP2M
0UseK+AD5iueCvsOmDTDAScRlRdiljS2fIOVMUFQZRsrdBO1xNrwTjrk+H3ez0z4
phO341Lqs9QfrBEVZp/eEQrCv66WdYOUwVxqs6O3/tOGsr6MhkmruGjy1wWeLWod
cE/U2vcle/k5EoY3oS+PVgpv0AwqLe58AgssbS4R6oWPP7W0M+hVi2wL2Dn101nO
2K/vksScLPYmD0hlweTES0Y4BOeG81zRLsExyMxD2OE73Gq/+tT80GTJeTlXmPHe
uq9/YK2+0Grp4bLS8Td9gXwiuLBkLYdOQ+0qbtEKmsyhJHdEI8/7KpG/gBWQpQHs
TONQlqEs5+F4EPrCyBbtslEBEx4ufdthkMF8D3OHC/k3/SlAPK/yzDLU0JpNnrRy
At0ulukglkdHkeEP+wttwtQczrSEN//3M2PLDndHT46F2drXsCDQ94F2k7/GCvhW
9QYBOVZDxFUAOy/9mKAm1dq05dVsxVaJIi8qbZ6rspWXD36qLLoIAwX/iQ6A5RaJ
gbl/HIcRAm9hMV1ah21X9uxcbPHtuWavF/IxXjAWD932IYzHjw11344ZZ77d5Fy2
JZ+Fxpai744neGodeGDpUe8mH7sQdnhiPAFZZ7iUFJ4RySdpeglUKaRbYSWp4M+Q
iNpQC7bLUSc3NvNSptuNetCzpdIpYzFwti2r4tPxpISZ/76oFTCcdNvk/wSGd/fq
Aa/J812/X2gDOAuvunafP4AkbrjL3lTeEyTD6XMbv3aFgQnl46V4SAd55Mc9/Hx5
l56ttGlNwVfdMt5leSyKJHzVmtrdxMytb7JwqSIuZuT9QAUiGYXPfhBJCNI4Zheb
9qz2QLDEMcwm0VckD3mBXtSvnBPOz282iyu2MnbcoWNBJ28yWr7C9YJeLWijKdF+
5DWKMtDN2jcYB6efneUJ9GoXh964IFkOnQ3OY9uluM+uZs/Nic37Nx3qrc22YIUB
XNqTPl33x91iykbyf7MpWXtihDffpzfm7dpaomw1ZLGXfbT+DOOZOhek9JLeU+O4
uvVPEBKhaE8jWW0uFHjN7mbe5GgZYFaodj7H9uGWUXajEBmZuJMjnxPb6PDoONeI
pt9r1sU4IhLdyXlPvRKuK7+kMtpuqKgvzQehDRkqLb2pQdah3owRLVG+qtrJ5MwU
AjWOqv5GQJAlGf6XMX4vS8jSVDPHMTge5DocTcOxPmrwpwzvCipliz1auvdlknD2
xo2mWyAFyYXQ6F4RRWAP2tnuyscoaaKnOf57d7YZ+MKa20UCPcxKPEl4ZUurtwBz
M9DF4gfnfhpn3axZxev41RSCd6ebeO6UXKqXLx/vGpe5umut602CBTqB1luZodco
CVXcNluN0sPtUrqGlUS0NhHryD0xoLLSkKRxIXwadHToZIPELOBZIt8qwdKPXc9D
rY9U+5aeuLNsZULYANKl1iCZvayc/War5m/8CDlfiXZ/Jjq8W374gI6NBVxBeTwu
ymJjn9DPaZ0bS2TZ3QRlhNhrpdAsFxC63cBATeBtJahln/WyRIFVAXHTxXiNqKXu
W8VGxsk6JXwpI6Kcp8yFiuFd0sWEhN/DJ63PGzf6h/XYx7L32EJHSMYVnrQ4BLPv
hurGvHcOhcF+EHhLqyyUC3iGbS8YGg5NGSyqgsEOLIYNBPHCz+k2o+xQ07iIbF3L
wDEXyWz3qtdjT0WGvHMBZT5ln8kruWN9B89BDLohMmcerGWvzsGXdDF09NUr0aGF
2hp9dQ0ImtuoyedG09Ag1m263ONjym9t5JzaOoHfX1XE3Crn8379IJQqDl+CVDey
DX5/CDH6hjj1BcLSMwD0Thc79ZbcEHT5n6ez9puj40F+73bnm2dxfSO3+D7Plxv9
duoro9+NihDKKkrZnWTmBO1lNNJEaRy0vj1a+ZwuAldaR90LA0urat6zduzAQw2a
yrzb6ZjHKoafDRNarxud/+p5Aqa0bjzYtJ+FevGWY+eIzTK2wbzGVEwbeDSNVAJG
FcrwEQBcZburkH2pNyF32HppqG5jRN+6Pvi6/8G1WFGw2XABPcy6SuQoOaxqbo+L
wpD/qzwCg2Pv6AUTTZq8/o88vBH4n2YvGm+tE1CIRjseOAiRhlhF3uuPamfGZNMG
SiScFH5rcCdRXFvWL+Lr+FdBArtdJGwy1wpPuhhwDBO/ceL7dFrT28+e2Qy+ljbx
3NVVzB+8IWC2mQjhpYuBfnGDdzfRJ7GKuyq1gZWrkazffa6G5kZogUeeMT0z9EjH
9Xhxx6NuX2yU701k9QrUS3VngmFmuNJ8ozzQozLZ1gZpDnm9GKCeLTFuDCwwttGS
MomF9m7XXZFg6y3kwRILb+47iOIAcObe1u5MBUeghvjlGP5ZNgskmur7IYR/fxKJ
iH68FIVIIgJJI5LrpOSjWTia9kYVtG9LxcZdG2hplwu6HecCo5RN09U0GWltsOyb
nQu6p+Ly0mQVNptcZVcCUGqSXyZXEP6DDbM0/T2XeR40itAwxtN64i8w3JBSX4FW
LmJ07yl8GM5Q+mdrXKWs+ndno7zFxcCtxJ1FV46aMArsq0KkH3uyIN0iZpy1z8SA
ArCORgGKjqYYpoYW+Am5Pq9sq1pqySoienlk1jynZrdH0uBGG3L9O47tgSOLiP5i
yVa16urRJw/VLghPUR7S80MBdZlzcK6l8mVL8mM29hbOCdSa49LkLS8LcEQO5NJF
reV03voT2DXWJj1CVwRXIz3txc/X8DwaihnBTAzIn+CvYp3qRJ73BDVRrMAX4kL8
NkdjqmK2Ka76oEGsi855wZqiF7RMlqRP8JTgpGOFAjPLMHlX2c7R6aY5kwGba7b0
jzRiWarAr7hav7DArILkZSHCheMK7+sWwxk7S+a0zdSSQyUdr+vUupqEqsN6Ueos
fZRZRO/XFYu83FtK8vj/vLh3yaMiPkUtLuZeNTeJ3+jQ/KMu59TF/S9qUudxASuT
GOxrVSVap3IdLYbrENx0cwATio29HOw8DPm4mfR/d1CnAM7TiilebpX5rM27mcZL
3nkN2xgZoWGg7wR1+zXouDGmNzG54CU50CwT7Wc9FvlHS7vxUDMcqdynRliRV9MQ
MW2LLO2OUWhA5aGIPD7zpcNAQEU4Cp53/gvLGetK+dqU2coy4ZRqS+n8Z8+OXWHk
66wCy8ucw31XN+P+mI9HmslZplIIgAO6M0VQL6opaSq33jcq343WV9K5KtNhiZsb
DZjAnnR1U92AOUM49uiMfHwmlMlsvDQbN+xeR8d0+1hZu5zuXqiQvXrV9oiShIrc
QEjvuhZRryKNcgUmVV241y8YDQp3Mdwyf+WT/COsL7pv97KUpWIXE8lOVA018AQh
392LgqJZflq8JeASrsLGXzxwHGW/XyDbZHKUHVkZ8j7/jgy0lU3k+76ck4aX7g2y
vPhxOUz44Ro2W36AU/5JtLfbxCqKT3BE0weybeOERu0ncSH/IqU3BBbvpzl7j66G
+GDDRQk/xJIgOLJXmI60XyhBIOb/OEGircekhHX02dPsNziwQB5P4LLqYWV2qJnh
g17jIW2I+jzL4JBYdus6sac4ZGhCWGOQ7jya6gm/aft5CnGhPeYOYX5XgW0LFVyf
A0g3gjcSdw+6hdm329zZVaDkwTZm9zCP+9JiMPiHTL5HPqevcexMzxriTdAIoRBI
C5izwmZAGtnmnJrTsW8P+7+w8qYhMdjr5/4TXyZyEjeQWv57WIVpXw4d4dr9pV+t
TUS4umzJB8FBsyUyA8V85oEkbAz+m339Q3/xiSwVY0SvnSprTe8FGO5rGh7vD6YC
nE6d6KfMsXogXRnI4AiQ9ny+Uz2jMScN0Yx1Wtd7w1S+Wyg2rfFjjlKsF8pToBpE
KuHbK2hEUQ4xTFWmPXHn7Y9uA6y+6tZbaJlZSNAHHwj1/Aqvlt3b2p9Oia2QqPGc
tpaugDfCewG60x3N+GK+bElX+46NP3n55RXDcpd1LkHMh33BU9XJuVPLrZjX4yCm
xGTUCJLgw+OH6ZqBlxNh7xhBMWk2/l0zyeKYCtAcHnxtsMQlkfQOdf0viBXtXt5w
KIoFkB6MWIQvsTYZFQW7ac8XvYXr8wITImogV3SzbikYTqAwU+a4xE7iunuDdDAY
2jEkA7pb/Cxj+IxnYbTTz9xQa5FmjyHFTBfthHGJ7r4T/+8+iC+NCOMe6+2W/8fo
hKtfEZwp3qURo/sNO4LYVIOnlMCBwWXfljJK737E8u1Tw1ocsIC7iQpY+vH7VSbI
FeH95zaGh5wGQ697MgD87BJzMUZKd/IIHUSGpqFUeS6TxVMsJjLXaredusb7F1ML
BAlQC+ZSBX9nxPl6KQ91+6IfWlf4CM3FjHIOBxk+I7LL/wRkrxjsia9IhwlcM7FK
0qsZbAsEbFjnNZTWeQ0uXxx/ncVqgN3KCNP8MVBeEtJBtJeX4E9WywPGBBqWxcst
+PyGc4+vQx63J8DFXt2ju66jrH/RevxXPfaUHbY6da8JGBzzBqS0+xDxJ9XjQ/8h
IXmpa1X2AZ+DkwEp5RtYkTeE6wbnsSjhNGSSh8lGbBD+ynNddH/04B6Tnx1mXEF0
3vW4tXkYtqgeWqGVlBrSPgBCTWr1rQFgokBCO/Jnh4MIQm5UySaxkJLGTPmFfJcL
cCZUx45yIluK4Dzc6XidaG11d4lt7oe5OR5LkoQB9/vRf7F9en2LfeuVUFYxhY4i
nDgw1284CbkemiuTVRnxJV7HLiw1DTwpA+75l/g5YpM09swkRZCS410yyOE2mPLF
/VO5y0/GCsXHGCIxJ6T9bJWM8n0zztoh3hfWKqLrhUr8CRJk87TkNYoHWt3Aj1Sv
3tdiCterfdeUrAHVpOeont4mbuzuGoban4a+5wxjsJ9uHdJYtSSwseRy7bupZSve
H4WeLVUdf66+B9ZrxecbY2xAN9HkfWbuEn38Pe5o8unL3tfl3ZyOTZ6sLxYVQx27
L3yGoQhi4dY9EaeN0ZrrmfuNDCd963XCZlXB5Gt0lLyYs0AoTye1dcw/bOf0hz1d
p5UIeOB/H2q280aB+nOcQ2+Opy8AhRPgK/M3D+sPlABuJNtA1XCafaT8eRMLEm+T
+j6Hq/fgogJ/mI4eSAKXt69fy8Gz0YheIod43Iz7pS+CcE/LXXHeNIuPzEs/LGj+
En/BfOe3Mp+tn/7xMVN/FPZ8/GYG1fijiZNx6pceFwqPxUhNeV8E4VkhQDA6zyj/
F/+PiUqghFeJJHVKXBQCw2/Fa/s7N9MVebaUTYiiC5Hh6h02CMQIu7ynTb6o+Eky
RAgmfvHRTXEe7A4bIuKfdzwohCY11ItaKaC/2CuXw42b2Emp1kxJugLZS5ytP6A5
MSohsinm3D1U6AvNyC45mKnutycW8knHWkWIvk5+u02NTobqn0A3SUxiBFOAu7Me
eTaXfHvVx7ExqIeXQko/I6y9A7sZxbgldCzQ/3QJ+LOqO3POxLnZ0j7yKV8af2iu
Hnzf8+zI9NiXEYyGpEgC/qieIKVw5bkAqbqYJ2+7+0jq5wNjS/H+fBp6sqjpkM44
try2r2Q1T64OsmP2J4c4jDjvP6EpTK0aAHjC2eUrXOixXqRaPnKuYbMiZmedyfUN
VLi1b1m0/ygtPJeN0avgEE8+FrK4vsnpwqKHRnVOyz/RAFZPzd/jGxYly/WlDA2K
N9/1cVrDaBWapSgKjh9aALtquuCap5dD4B8tqn3g/Mb/J71HkMhuoze/ZPOCczuj
MPzAPmnyPHhv6IijhbSdslD2wdnAdwofREFMxIsW33raWFchwlvFh4rG8FdZksu/
JIbyrCJkoBjxLcWUAz95UoegJVM679+FMseTr80RDZS4soB0FlYsB3AmfWOqzXSP
s4lt7Td48+numd8lQ6jQK0SwSIOS6EAXEunzmEyDE/HlECrPZY0cbP6tFBcbvOKi
5lkyiERstB0WdPq5N86jY7k/Udxse9VXeq2tDtyH6WrHbyQ92+YVEEvqXmac/KzD
wSLuMwcHeG1I7+Dp85IfA1Fy/dBoIc5BV1Ep7xGbRX/AslTrflGIxdiXvLKbl63I
xT6NSbvRbuAvMqG7+7tu3BySwbSaa5/Kb68eYl2C5iW4PiFEHyMuuGdCUVZG6oDW
XAh8jG2twWVz5trHEf3wbRCrpFDfSvIkgPIbyIbasHHVAJ5yJaKHvV421PnhsQUr
ny84DnzUgez7edaEGB2yUlYfU3Y3Rn7HqntGGS9xVz9heLcBfKqXC5ROaKifXxTh
H016HkDuFG5p4tgWjloM7SOMqKJ2bJIV42hr1jHDSK9Mke9Mnl9ieJuvtNmr/3sX
ZrpKTd3fzVIoNomuHfkqdlxvPHg9v0W8ea01lwRMtxT9OlBtj2d61MGckVcY2/Ol
eUVWkk/RIuEwk5vuB+lbXPKT4h6r0xbvWayKrV1OytctzHXmN5IEC/WjNyv0stmY
I4v1KvxLzVVnce+bXj0lIEb4Wgf9oXUhKtVzCH4Y3bU8o0DKvvWr3CFqVWd7gGbJ
eZpkWZLhpy0FcaudFb5L9//1QdqW7nDY75p6zh0ooYTYEPN+2vr9reEZ0Gb4RETU
99t7NcxSD8u7ZZns/VMcpeqMU9nU1L/9pA1oNxn0If5RMQy+JtwaE2YtnJJ+JDG/
TE+X+FiXhni9NeioyPNMjax8fHf2N63YAbgTu0JmOgklhLeOaZVmKeDcb+s3P/Hm
13uShUTWmHGjFotL/SP1EG6GsYYE8/4b7tUo1issBvooQSkmr/xtSLaZkWJPyAAH
LwLw9foyRXx60dOlBDu2asqqPwtlTN2JW03C4599bvsac5w8MhG7NSUD1nkO0l4t
qm3yC4w97o9teXkn74rGUof2lhkqWLLb9e9quZ8q2LoLsheeDW7PF0tXl/lRTuZh
J3+y6wdNc6EZm0BoW+OfefGui+XJVpRhrtcF0evzCPfndNGGSYJ5dTb9pV/RHuxf
THng/eYBFJ3rbz+cCWf3RtMtkLMkZ+U7tj3HUp191kD3mPPuEXyuPgeOqwv6JT4A
hwlWSc70K3mN9HUxkvOoFhPxgWZshrnvchjGBkbfgK1oqCIDyllW8Ue5uEhODuGy
iln5Q2liq4hLQ54ASKld34gaCGk2GsFCwF3BhNIChvvnzt5BKzCyJ2ENhJRht2j/
X9Sr3PnClZMpY6KtlgTn3tKJqCZJs4dAAjIGxsmtxGk663K7rF9ZrvfjJEYC6wP6
ho4QcvtOyJ9VDfhkc+1wUxURa33d68JrEMh+MV7iDjNSVAMn/tnyESdy+Td6WT+z
Ycidrqp1k2xmmyDXZe6vAUpT0gIDrYK8KyJRcogjcagvLCGonHLP2oJh5NsWYpMI
KyZ4GRTiCSQzqkunj9/Zm3ylYuW4xjfIMf5HNwV9wAiteVfwYdF3MI1IRKLNfZ2Q
9l5ZTlbH3OsGx33jsIn8012s9t+woo7pj36vxFqYmiIVpgrcVbSMOydkO5L8KHSF
rJz+skArSdmSFG/HLmXzkVIkE+MRhBlYBJmLVe725zUIEq4p4LIiMwASCFEhTdmd
CMaOlD+vn8+jl6C04RIz/pCzfdEfOXTyUHz4cDQ8/s2IBFp9Nfa9ueEVrl2itYrg
xBxIq9QWkSVknWkb5WvSi10PGtmicd8oSNd0M2y7cQx6lcsj1sFO7QDxIyDM8lG/
+ufqjed9U9RY3kM8YLyFHMxhVXdlVyJjuwQ/J6moILJayLK1CrtqBCvcoNybEqre
eay6BuKjknyeU3uQnVfUsdIxO8eeuYV2PkEPEmTU0g5wZqIziX886dwlKisSuH/N
jrVnGLn1xaf5/wQ+URQ2T+5fiB+ya1F7vTfPFlcDY9utz4WHMpX2lQPhyeKpncxJ
lM7/lkz810p/kBp8cbjGaUB0DeJMoCZ/CnlvSvU2dFj8+MXY0syny4B0bKMi2hYq
+AweIdczuayYMvTW1zIyPT7OopgH+Ufoj3ZAdJET+Q/l9NV/UvSNWrcjyPrYR0gl
CaiFLce5FIuD5bY9jnkb71yDWbd4wTipRZyYa1g1Ynb6/y190YA6CSvFcZy4I9SZ
iyTGpmOmOEdERzhU4kRuaPHf+NsTbyy3WbS1rIdh7vRUusPjytulopFcImScniLe
Gdy2z5rRadHRIhw5wpPqdqQTLwJoAu9T+RJw/66is/ibPX+9ak5I5H9kC8hVv9bJ
yaC9MArkjA4ynatUgTP1K54OhMepwXIkQgnIT1igoY/MsXmz9Kruc6jdh5S2oGQV
zyW2QWkTA3xRaPNUMvt+4Mzxvt20E/nuZDmUzVjfrSt5NrZCKeXBCCAYSyAuyz+8
YDLumz1ZU0pAz7mPBL4d36YVV3goH5ftNb7j+BdJUvWKlf5NKy6f5Yo+mmsH4a9x
WOq+u0Umzf7EjHUixi9kNIa0sJm8zjHWj4qzZuGPPX6/gjv2w0gSnbqPIM/TACIO
v6gBoOVA9iUbPCP2GpcqQIqm2kxub0avEZ5+5VG/gzSMPTqck6r+jVqfB3PGuEYN
VJTUGlDCptPvNjKB7m5OC3HMfp75UZuJgeTOguE/na58s6JpnpKFTkxDX9sGZ7O8
aSMmbUfTn5Wx4MZIe/EJn16y5PkRmx+q2EG0N0mJN7XC9z6mdeNu7SnkR0oH+s+g
7NNpdRCtNYVF9FBiAiW8vjevR5R3qc6itS5OAMRvriNoPH2LwMOvyBTF3HeZVKTZ
q2qKFw8iK+/jdkvBYI/wyOST3uqJNl/RgpyN93gjBjEMuI4JiDYFRIwNzRtjU4pJ
naJAGpgEuaBOqhAcjJaSy/PKzCSgQiTgeDR6pP3VcPMjU2zgchN8rCz62UZyOtEv
ezfUiUgEFzSm69BPKrrRtRCT5yyHdDmB0+SnV2um7XsFRA2WtxWtDpsjW+BXNFmW
9oGz34xkXDCWUy0lVg09hz0iFJDnNw8EV5oJYztL0yyiQN+T8SuDpdd//eN+FVya
Le2gxl6aX6aK0TO+W5vK9iuPNKmpe1zZ5rr8nO8P5KzbwkDPAewz0RYRPeawbKDF
CufzbebASRB9AiA3RhE41jt+APvPJOgI8EHx6l2OyE6SPDpkXOR6ZioyLmU4nz4l
FHws0kD8sJgJWKHNDxQ2gPRipgU8+mElgnhPp0B3TF/19+Qg/MQEv9Pmsv7ycKUl
3/HkVS+t1ru20AX/56F0LDbayP0A1fCbqkHAmagz2xMwUrkd7yHp1JYVAkmkzoLX
AWxnDjTaNP4ZVcH1SxmP9HjaKhso8ytpZG0qq4NdA58V+9VuGYAjn3RvK9znTThF
E/EUg9eROgm4Q+7qgxWqpjWnIoZQqYkkwEaUNuPCpwLaVBY/NZm1flq0mPyQDa2x
eNFvSoh55kWTWKKsHsYy/zO7Wg9cRLss6iQr0WQbJULcfo/nGD+7JoxU4sNxO7eM
EjNNEl2DI032aqdjVb9e/tgnWTZ0biNj3ym7WpLuBZWnPDbenu+w9zTAgGnTG9ax
/vJsAqEePqHVzzez+8q7rnng6ZQjJLCtSm+Z+tvVIepIDLQRT7WBltTXxhrOd+XJ
C15pxmCEJAHh1YQ6RGVLqg8+HVU5eGzCNGyAR49hxFpbor4Iw/XzFDaTxN8rZ423
0yioMXTe9WufHwfqu5tW5y7naTJrDGeA+o0uHxEOPT6xywAJQyTW5Gh60GMrfV7A
LT3Oxgbgoz33jUvVxmQFLmvsmBAN4rkB6S7rHEzqnt2mufngiGmUVJV/AlqX2+Rh
SHs2nUWcJKrtv45Kb5j6u1n+tAQ9g2/YdyO8Jtl8psDlXPsehAmc74f1v3aQHUDc
C1uoIsyNOjVAyf1elhwImSZyWS1R1/X/6fy4thqJmJ0+92+QvW+WbmpxiFXRoptX
XepOAh2Wtia6TNFW+LoerbIL2FuKYGN7+6fb91A2nUa/ZRp0GIgiSYG0zRcvpXfO
9JNcaCQcczDbVRF9/HJgqR9rZZJVrBVz7LP8rZEMi72Oohpi5m/Ng8QgTB3Ds2me
WOhkLRjN+lOIuQhxXgqGh7XGfV4Xv9iVgxM1SgJBnno1C7jlHnw6a43ywgYBgVOL
D0AOq4dtTwIP4hSpqxzSGExGoxWxe94DteTJ2CuxPg1lAvxrwqsYIAGi95iy/hRa
DRGgs03svMCMQ2T3IN+S8kfNTKh+rFBo3EjzICKqVYgiGcosDsOH9tOPu506dQPX
th7VbQT0LvX4B3KE4iqgpnS4jRt6nCI88+NG9y8A6Gz9nmtBm5AsgIckBExKZkt3
53sI+qsNw+VLxsf9cPUrNnkwGbZGsnhtb0G9/+8arQ6hzKAsIZhtJYU/VpiDm0u0
3QmMAVPvG+q6sWOFQWZw0Fz6PsJGDD+kwHQJAVV74CoTWQztJoyHWmRYPDtfiKLf
4oLXsdBus+VH621r9SmYxmi9ehWA6cDHH9vEKzss7JCrnfqjvE9hTgyHn0mjrpNs
XYMrRXQ8rboJ5uqII8arp8/UoydiAMTQ4J+1LmKwBiU8l+WP+N65njAy9h7Obw4e
JV5BCCRcV3sq8CToxAqfLezbbF2gzpzahDcBtlquAIBmWutf2NhgaJodqu+FUndc
UqnOBVyOfrVzjIv1attb2sm5J77aOEH5zr84GklHqOxHfoYgJxkg6/8CEdYffMbo
zPv3VSqyciKPUnEGNhmy8LfuMzE01EfhXJcXE3qUm8u+N7JQvBSGnHBAsaMVb/tS
u5dc0FkLZ4XXFmeCXzqP8ED/eDIOM5v7aYz1MRTknnUWWIE8ZAlK3EeofTS2VGJ0
bUCvNk2pZvpEljEdOfj6RyQTefdxdA1EW9FUF7bxIVB69wX4cLIF2wYF847q+X4T
lu82FY7ZZu0GnjKvCe9G/UIo8/XoUcW4i4VqGA8sCVmbA25SiKv1gWq4Vb7liMEf
tYOhW79Uk25aXlu0FWZ6Mp4vguvt5ZZ9p3/R8Wb4LFjQZswiXNjOwr0wuDuX5STs
qXIOqhDX0+/H1O3UxnPhsNCne8cu7oyWK8IYX89wwud/Op+8gugRiQjUdPPw2ibE
Id+F5LrJdEbl8Ef2G6kGcJhjW/a4fvfifY/BfGYeAGB/Ohu8urc+f4XNib13GNo6
c7WWyhyzrESTa0WJwnxRk78Q7Bdw1lqBpOqedmrdmy3a5qTb2TEJDdznYNTJ2hz1
dLtBH3QkbMetYAep7cDGs8/yCQvYm7VrKXSVkmEpT5Q3pYvSO0mAsGJzbpz2Us/U
RMl32s9TomIxRYJuijnp3NzmQbbFX7dIPHxmgfh3OVOT+o2Mn1iiEdtjhsCEkOpC
pPkXNYyfgn2KvAjD27nCh/7BVOPTaf6cjKOfnbsMZKvAAx95+2nHdEbKqzGUhT7W
wNGU/kVmKnUlyhZ9x2xszyLuBKHAj3+6UVsXAnLnH+q/HRtOuZ7yudgd3svp5e3d
8zeJMemMW7CYBjnFCeaSacaVAbeKn0UwOOKofTJS9prEDSEw4cVkhn6RdM6r2o1+
y91a60Zai1sYutXJmnNaImgzSXqp6aC/uC837CTfk5k/eCMxjgUqQM4luj2M45S8
ooSe2xMotJt/wPigH20+H0SAJmdRaX8vS2vePTmvHzCoNKtgfiJ4zBA38rx9t3YB
YDIwwJcXi/Yniwf3i2XOpx2YEgFKc55Ljnb57UZxA73bDIH3mcoNDA+oWGhfjcGk
iAVJwudFEVBOwFiRV8QECJvG7dPBbzFXteKiKSVTt/KQx7kYxP2b4DjboFKhZcVs
mzaurrfQwsV+FslEzAsjwPs2qqNt41YV87voMBFYMap52PD4gqyN0otnE84DjIFc
+H98HmRZrSbtXgzhjxYsbmg8AmVJI/kMxtd42bxKxGd0rxlXPJn2k+jt077qFeLh
7i9Lm+q0udmVCTfI9rNKOg/40JbH3nwRor4Lzfb0yf5BqZ0RlqXOCSKhEFzO4PDO
7ldtAblSyQfbCWwQGktvzEvnKZ13Xa5xaBQ1wKYIIEL4XWGfLJuzrLq0qLEMMVmQ
N5pTeFfwRCmXytJxWop8srwsq7qiNX4DV96YhZNFsCuqO0eHeSDy1YRA8QNTIE2M
yoak3EzautlMQhhJeiZpaiqXyFI07z06ivsnjO53mtNDzxuG7Zh2GUUQUWkSg72I
ei2CLNdY8ZzBo5G4nwLLoxc7OA5uhW/xrM2+zBtAD/YHsinRjPCgeLq5e49fC/cu
U3reEuEbOqU7f3J7DQff0OXicKJ/GYVqU1Jr+6LjegzPGS7uEz3OaQCDcwKElfr8
xorRjPDgoZzgriGQyHPKcmAFOxhS3+BqjjewSBKMkNcyuxMnytdT8SMgrU8tsRD7
Vu9VuBRuk2LwExB2Xgay1MPbB2+OO9qGuxstxEx2MLrIoaFcAFCvrIfZUUIbk8rS
gKQUP3Jnds8N8XAvkcESy/xL5iLgCWikFpLtSv2llMaIF/jdUn71HRUPPHGinzEC
Oj2/eG1RZUII4/mHxzB5dlejM32EjrY0jdYaoHXTdJ9e6bptonjq0r/GSOJLPUGs
BsqdcnnkYC2O53a7nqaMDzvjnBt+rsJBH/Xtcy2fXVoEoJ8a30VqzZNGx1Em2zd8
qMsU+sulVY5QqTgt9bNopRebc+o4SeLWrGpf5mdyo6vsjtizCA//G85+QRj1JDnJ
DtboapsWfX0pJi6yNOuIr/CsSU0TiLdugMzzwKL5l4tIkYTXM6qT3yDVzE10zp9p
vGsnmN+pGIrQbdzkW26G7BT991R1P8eCMEadC4SP8WqSNJEmIOz7TLneOqbY/suN
/2O/BJMpKb7ALJepSkYLbnBlJpCUocH4roY8sO1J/C6XDnwRiwZAwZgBJiJVP6JV
optyvQAtxYgZJioj26K7RhuMGm1d8+ijzxGZ4AlmxI2EzK2FpcQARNssZwFixBbh
OcCCwYxMOmQ6bvTrDelXECbiXOHkgCy/IJ9e8HOwFWmDVYlbt9UgVRv7ViZx7pYq
WBY2qNy1HzOZ02MhBIG8VUXya02KbtWIeMNYNzKlbmjLdR52ofTrHQU7YFDdDMy+
VqLmjnTNHMexTzDsdC2GlL5hqlxrmQHomA9YrHfR1IJe3TenIjN2B3kiPOpFaauK
4YzUB/ZRvujeCG9oio2kQzcNBTtsvBLqUhlIJe9/Up5cqxl1y/eJEaZDM2BpGDyT
NMr3R9CpP7ugKN3ZxROwyFxHfWPw2XNQTlcSEQXLZ5tQ5pHDullXq5tkXrg+vZpD
OvXOjkkTmg7gU6kxy8zGNgh6uGxK6ezDGXnLpyQY01X6A1qhHnmk2z0inS4Z25+i
N47urWjIgDLnL8LA5ZYCeXQNGGnpZQO37tNHBocw/LYOIqnjEIWwVgCjpa13OPUE
zMt2qYXINs7uhqlOVQiNk1dG1uCzInJWqOjSUjXxkkmLNL0YcQg5vjnh2pn5jIiJ
+3nHz4mwe3XfB74xC4FxVMbQP99vCuBylv3FRST2XiAwM855g5DYUb1nudcU7eVQ
0/7/lm/lyJYA3EE7CJmQQUXq6TR9D80B3lrmJYb8t7NYrDUsTSgKb2BqMVG8fNgK
Wt56J/k8xyx6CwhPP+CbmVgyESV7LkS0OitEeOvyCNjoPce0uFx85bLxOgHcqNLG
0QQQ9FNwOpb8JemcYtYXIMNoQVTOnfhP/tjJoQSoW65E0Oj1UpBlMb1E1aimKg7f
QvKLdHl1gdPXJxLLJk8us3tAN7WXEfFbN6PXDTG/Qc0MVPFzRNPiHU9PhJ/irUPr
zwvgEeCDGgaM3byFPHBypeNTy8/gdjTLe7lWoXKPkMBaB0w+waBgCLak8T7aG+BN
+tOI9a5VPxP2kwe6lPUHrp0tsSF9rf5dK6MURVdBYnfvjvHQv1CKu91msNK21w5T
zHYg6kf222GxPFQ0vmrYqD3ca9XqTUcTTNbpC6jq7e01P2TDo3Kvk8Dna5539XYx
2/HBH2lFywaOO4TZFgnivm14XXhmHpcCCSgbZv6LsJ6wfbAsxwD/xuR/uKK2CGnI
FkCejFtrAF5mnxs7RiRwiWwXftLdN65gMvkSwbH2rqI72uWl8I1XrxnIYrAHBb3A
IEsRvqsKFGEMm1wfdnprb0T2/F38q7xZ30Zrh78BcYGv2tPhfmq68oZP/3hUQegU
kPxhlUleuIEBfECs3Q1dzqqlSL6x4q85NVByZ1edqBOnzHkXFuym4f04Ox/4G67P
HZbt5HayBLnGucV34oOCRVEgVKAR0r6VGYTlHRJIh/y/kuwaXXQPULzbgWC31Fwa
zIaDmi+5eTqCFm4xXDxVi5LURq8iEer6SbgYxGaOdPCxvsXCW4LktvfQWv/SoYQe
R0cooAQtFvyNIqQ6r8glcnLRl07/PfpQ85jO1APQEYosNlJwfXIxSPztqAnRtTl0
eJZK9uWq2q+z9OR6scvxgo4coz65+6Imy2PLnGvjC92taRK9UomEOTbVsC8buEXN
0FK1PkGXl4LfzZsAn1PmEnw95zEDA0Bg3kVhi0mP0LOzl/exrkgosIrd5cNM0rzA
L0RCWyr5yvbWOOvfZ+HkAXK2imne71LFMrI/Om9TD3uL7I3eu2oL6YYYDJyUTpHK
2YbEqlMTv3A6n3eEZhqjl29DvL3eJ11pcMtkTH2ZpokI3A0l9M8VGhjqK4Mdmvqy
pIm+5ypmWbIoFv1R1hRFMQYseM+qIFlIkawQoHfFz9I4hlntajT2iuoqg+e1+3Bu
/nW0WlgWlYsyeJcyhBHc5giyU5KcrblIHCDAPXAKIJSxrSSvPxt7J6iR2/rrTHDH
DhxuYPWKPFmyEsiaGCkSi8yxJbbL9MGLnVAoVEeYN2FqlB9fAvkPEfbkGxG90Mdr
CPKlLOu6wckKeO+w/n8WjBCxw5l1SUmeOWcEwDcMKqW1itQMEbJngNGLUD1Hoyg3
r31pKAgcSCUEGLuJN0TyQachi+G9OvHjsMLA88EZBWihpTwLZdF/t2+Tk2r7xSxl
QVk2MhaVxA5wggYBe6pzuDFfi6mjNclunyEjkLNyMoUv03ndWt8UAHQHeYgjClUf
MMMNVioBfc10T9BfYGxoAvH5/E6QgWJ2mzpq+zCIujeLsopl6OnErZ2OM2Q3G4mk
e0XhPMQImlNYend+KV65zSou6sUOMyIE+M9aZSc1ZiPbBtW1t3x3fInoimjRPAJY
VlJakY2mQvlhObL8sr2wLYtdjaBSs4CQB+Y/RR+y2srwg5CtM/Uc08eb4GA0qbnD
8E1GyB3Wanb88oEK2CSeJd/6gGdB7UVHIDyuapGjMaMbHiT+ql6s5XUpljRdrT8/
Bx7lZ+jZm1AAXeAhF2GoY5sYvaBkw9oDX0dCNor7f9syRSgLZczfcG+hyXRNDxAA
BKsbBQ495OIOa6JbOHJ2IgQJXHd5MwcOyEyg5kGcwS9f3fGxUtFu4GWx9CUGlCeP
v0tM9IhuKtRJuqYonmm/DZqgtg+DvqjM5tmVsCkwIOHksb9I3Na7pH4absKf7cMH
le9Su6Cu1BPowaspC2DnjibLzO6ebto8ptFdTM20br+Ic3QjXIUK8UKtwEz9K1e7
UKaetFdHXZDlXzfrULbRa8ahkK4sb0D3kVVNGXQCTKsIBLLivPrKRnD6g41Qjikd
Xq+yO73m22v9psu9Q+bt4oB3R49eoPn5+JXVlkdUydAPQlP/f9EpjVQCDZc806Nl
CstLbOkR0tuOEY/UHowhQ8xWsVQJC6tLLkN4P7bzEDD2vZ3H4k31J4eGvLL1ZEn5
6sJq5VP/c1fR2An+hLHlFaN4yohk8Y74FrBN3CMQAOxji16kHo2cJQ53EX2M3Yv1
QjZ/1HcbjkcB9CNIB3IJTA3lSJ6/mQkMjt/TtEtBhsBm9cm4VEzYoFNUGECvoVHY
5siNyCasGznwnKy4Us4XwSyQMS6LrQDmKiB7kGONrlNAJNdqrM02KkAkWJ++XvOC
nHQs7ISTGhr6nY6K09LnfxPsntVoFhwapno6BOlw45f7Y9G5bQyvQ4akx5k9hUte
kGFkFYRh1NmUOFTZkQahAObRsNuXjyNK06462ycB6nWFgUf3wL3Ii6eIueXXcucc
uHwtYvRr5roOTIc34OfPU2UORjNSc9tHDA+4x4DhGX1ZfOt3i9+aPQziubAHzP/C
ioXZLlJ0Bv1u9S5WEB9qVhvzLT2faVfp6S6kWdmcvf2n+M/r5nOvb+4y8dB9Xzl7
fY5ZYpE0w97eiSV9AzwYPqLFZiDX6MgbXKg497gPA1JKf/ZuOAw1axG5i/cRq0Gx
8kGWN9qCeQgrItY4LAjM1BAegLJwpTWPAcHqxE0OIMFQviruvZOjCsg84KQJ7Ufj
shGt0pM3t9P46Bjeds0uNaFRrdNpvgLV9+dt9ERfQCWAdm33cEC9tjuVxFyqWyFU
5cXtwu1yuOoLZC3K2mDdg1urvD+oMgw08uWIqScSwkgHHRjTzr1mhyleKQ0VWf/B
rdC0gwANK/uMSrNDWgsCDXAslrKZojK38SF6zlXVxAJHLYEV7+YQJFacvjXwtZiu
Of59tJSjTVQA/zwCjf78Io+gfrC2WjP2zyILZfOTOIG9eWQ/Iy/7ebKHZrHJ+0o0
n0Mb/bKlBlsMjhDjDBuacMu1TC/MMiH+gj/BzbxeyxJdH/cVwnBaQt/+TqBLlepM
oP0aCvdwyYO4GsEByV4pXsHjbqU3bcXr3jCeV5JojRArXlmgFdmmCuTUZ1nEKSoY
E41MVNeaajBeHBxiXDQmwcD91+tJT7zrX9XKSAuQmFJxFFei9vpv3jvnC+pkEggL
nR0x4wcg/Uv7nxJQf4anFaUUxHaAxjSboMYkwqjxvagR0XZdPRtTg9DpBmtoTqo+
2p/SF14uye9Mx34njtuHGCUfn8pSrEeuytWgF1ooxGVJuykFOMpkeL8VYpcmm5iy
dk+E/S+69dNzIibcQZ3lZFgEXWq30ZF19HOiDExQKOWIPJRvSjzyl0+NwydoUkqO
lfJJdlDRfvhcN4GIy88VUQDJCSkLPZGFOnYaBvAlVFBVRIGvm+7NGYKvXYeo2KP/
7CiTMfuo56HgdCGrtmBCDPp6yL6G9dgT+2pseoGU0HFkY3BUXGMLdY75b8assO/W
Gb8rqd0jLz+7Kbt/4V0eo6Jy/YtZDAJuVV6/X8YbXF7K9f9eZgimCEzCXSIQ3F15
x0D6L8dZbp9/x7Pv+QboEYPBtsLmg4M7NqWTKYd+ApWjLq5esrRWDIWQo0cH21IC
ZCVjDWZmT0JcaazJxeWBnYTW9nzXQyY+vnZFQZk/+sH6lt2RIZP52366L4cJqA8s
VbaRc5jl0mmPvv3kY+B8unGTP9FPWvHylxx3bnaNEJHXXdrQvCFmoovNWaNKPgHH
EXxdSZ+AP9uhBEGQRnM5JwiSylFGHWLWFri/3pR6C3lpJp6rTHClMtNBumVNC8CH
qhNe9TnYy6zxi9lE9Rv2mKaDkKnEQM+oLyEnuWmzuY0vANtqhOR3yCLLXxF9NQlt
romCFLoixR8iYBD7BLbs1CdT/5NfLRZhvmjp880nCMm9T3+VJCrMmY1NxaF7o+uA
WJnTVAfHfyJ2xc4KvSj/yB6oy8rZVPdB0Fz7/n8cSIMiPHtND0aV2J1Hn5ncoZs1
J8lfUYn+1UxJDxorvDtKgqrcZv+p3WXd6Li8HEevLfYxefAouzQWPANvddA+8UeT
ooSZsvKJ6OlUDe8XykaIQBI0ujav1pwq5u933AJA1j61dhLfjkoHhwWMVLC/4PlQ
piZf5wzdlezEYQv5UP7Cyx3zt9IW1RwZ2Nq/r3JnQtcocIJC23GjMpHb0e+pLvD0
4hjJ8JyiYYzOHybnbGebonSSMIrqiBl6i48FWG6b91OxjNzoWy5XXsYBNNYhE2JT
SIB/VV8/DBLnrRzf1uW7fVf26zAgu57qjhmGMs/Vmu6SS3krNNIDZK137UeFVyyb
4MFW0TdOahCPX8k1UE4RV1NGkb2hu+tZtaP/HECTv++8XKiPkSvlfU2rklHosBzp
+dqO5ElxoojQqfa/09lN6OKxRjpPjmWGzRCeJnqXfvXXvM3O3b3QeCblvH8YVOZV
chvl/6FI2EAVoEMNqxdUsPjnpNEj2NHOwYXhElmjnnJy6AI0H0qruvxqbsGyaMWL
qM5IjhqwPwZRj2ntFZgXuqwoybWyL3rutmVEg5aTYJr2L/WKBO7zp+sISNyjAnsb
j7/dNXBy13zs26cD7rcCo2VlILtz13+hQns3YPK0CUE3zmBYykqP91ibdhzRpB6I
0ljmQ6IHcKFoVIib1agj2ICr9t+6076f9L4Vsdvc3exHyyimHcIcVaekf96hc0TJ
vXNP46i98X0K4PqJI1nHEpvIW3vcrpbbMaIIKas8MbLa3RcSLY7z3bgiUC6zdHW3
ytHlOVk8a76898FqitGs0srpuJk3//llS0sPcaW12ySBlkbi89LTJ9zV1O1DMAaY
vbGt4FeZ94woF3VV9wAbN7gJrikYsEXES1CMtus90rfns9IummGp08uIrCecrIgL
bZo53mCI7+gq6gi2O/IuZI/gwAJF9eB4dHJfnE+niG1qXBxBIVY6jIzkymm8Ecqc
8xZp2wpS3IjKxO3ATVJfn3x99IXpkzpe+BCe4JQDr9ypt3vBQLXh9NZMVIJ7n2qh
mgkIV9baVUx3WKSdTwFcu/l8w6DesSEorj0HNz61X+QMhZweUNKPtnDBjrmF7JWH
a3lP4zbdO5ihIMxpiajbYJjlR1AEYgNwYT/HVIX9wg1d6UndDbk0Um0VNB/Mxryo
WMsXtk21AOjOM6Mbu5JMsVwzbaT/S5Umk0mOajC9aageifdqhMJqpk2t5QSt1Sf5
zimNCGWalgL0kPJZMOEkUYTZNk8Sd1uRdv1Pv8zTZ13D3iSc2GN8Q5GYbEhtEuKe
trLglU2AeWfw9HQX6MjJuvSzXkYi2TyX3pnlB7/wNlT4IQCA6BCp+HXnDHApnxLw
sHH6qJFbqiTtIx7E0xROn5m4lq6gMiqVfWQ5zhfx4+PPIhRFMizHvnV6XSHHN1Ti
C0EovpJRMaUxjjKVRma38TQ6FOR1jG/+/O8tUXOwUfE6mURX0ZY1RIc1s35YfI3j
uZ86LGAoHSLPYjreLAGErFBWma6Gb3PuN54voUCn1W9s437GTDWG8xWehzZmAylJ
uXUO+UQs37nKz3De1mfkICsyl/Lfupy7RrTdoECsxrv/E/JK45CuVG31XF/nkSAF
LCkQ7qD/b2/h2IL+T687GJWG28XbK2qJxeTQYFFi2PabzHpYiZtETQemfJ5tbQJi
cX27ts8zLjNrxy0cc3jjMsoM5X0CsUKGlG//UDLaWTYatkWylzOkQrkJv2UfhmfC
hTuupWwqVK9s2Jr7akSMjwSzWoVJPta3gTNVRS6KneK6wzp8AF5Q8NxvhTj3Nkcv
k/c1OFJwsbMpu8fTh2+Cy5o4Id5rJtoxFtkFh/IZWDJDQRFtUrgfkhpebMqbQCgz
HVnwaHyZMKEWwT347/6LqMiyR5tP6LuqayCj2iSwT8cqtIdbU3rA/29DPzFeNq8P
vnQFu3vVb/yDsCD8+4bOOfW7qjud7dzOlpP98NDPRy7nnduvOor6Ty/EZhqtKg0H
m64O//Bd9xXK7wj+xXTWeMdFcvZ1Qu7ZYzVL9R25IXMoIeEK+w7rSUiOcpP6PH+I
KoJVYGkHyM46MMmkb2bSthzjZTs3a6CLXYBrdBRoC8SHIWj839OknYiSLoXvLwoa
qIT2FBVR7OI8NAgKZjYwrZG6oe05AB0mdt3tIqiJ7jZV9gXER1Mt+aawQmAMFrLr
yYFQsOLgwMVAblmhpimOXA0jk73+1rnSbGrAPZn06JdOUJjVFGDqU7mMxj8DG+D7
qEFda3Cqj/qVK1cqwTaVVeyZnlo/9rKHe3U1Qe7J9FMkRR8/WDkEub0PhB5Y995I
8HPDTVK5HBgBBr1pDHeQhZPztwPQoz3O8Ycdgi23Jcb+6t4SsQGT/prlAbbrVW2p
HwmLi9HDe6UI94qvw/U3tecPEhiPa13aK+t0jDAX4Ysb8vP9XKtPOKI7QOkNeojw
weIdIQ4UKLWnwW/BTAKGiCGvju1U1QcNdwv61rZT7a33LpAvYYbp5lR6daNKqLCi
E2i4AMUYrpS2Jh0hdt2Rh9BJuU+ojhIhrFAKdmBvqG0kmYhg73pRVbIPrX1lpn3B
yiD4ksxa7amE3ri8fGQeEqJUWPMxFnYOrPMElhnYmuSn9uLPyfHFMtTgkowcMVKG
fkaQQhQHcZSm7QLabJGpUa6RwXnkZzIOLqEngtaoRJeUdoyfUO5BF+RQEr1cHrI2
WcA9dovoZDnvoTtyfs0GM8vOZqcpYi5EOsLX+I3CmCcYNROltg8csnMS60MIkmVA
f2kOExSFTIL+7b3M91PgElGh9mNYzKPDjGRM9+xIdSINKQtwIRx7ptlDCquXqoig
4fdDaB3aWz4oINyIDm4rNf/y+a1RIqHGljna30QR06dF/qWCk3ZGTA4Z5mXvGWGH
MmH8/1AsU7Y2J7GIOZ0um2jvq5TvZ4IuQu9iPYlvZd9hk2jdH4yer+ko05vJvnKw
/Hj6VEk5Ss2wC/6rqzaChahSIpkLSrNVdfVDoZ+1p0F9dtQecZnsRtmEEvXE7VKS
sy9ktkYYHj1w03ZmtLZIfYO04wgbc3eU0mvyEdHc3FGe8mF24YHvzzIiXSgQYF4l
bBwRyCGpR6GGC2NoiaVBlETjt6YFJIArdVkD9WLBh+WOVA8+OjfIsqLZkKZzwsyK
hofOuqZqp1pGuIiJKcKsRyxwrrqM8xvkoPmfJR8PB+hewfcgC6UFFrERlqU8hKX8
8H2zaOmsFYkFLvS/HnBJ1DFl7r6W7MPbmBXrRu+7/g/Uh4GgE9zWQaCz3gtee0IQ
6EUmf0v0TPkFfllthvi49ousOHD3oTiIVsYATvLkErTsLFOGHAcK11zoZllvc1te
dQYpFe6g/LmRV2FP6/LepUQottbn/LwEemKWYczDlJFHa/8HzW+eRRF6qTx0meWG
+Zkp3yJzfzPL2Gp/wVAugAaa9f8hglIZUUJpNJfQo480dHyIO//sGC9cY6TqPnBJ
fmnqQyg6IWyIZO20/wrVge48fKeeGqume7wpgHfO5OWid2NC6TThGGcmJmXxCL0V
C0u22DB9xIJeJcp3k0p1jk9F4sfK0XBy5yX3nfeTrTAJO18L/TO4z7MNyj+2j5df
4HRyIajyiDs1Y/e9c57aM4dlInDLtwj+AugFtPylBQO3BSxconWUrtsFN71KRpRI
Sf/aYN+3P4B60EHc4X0IjJTJgUt+wBvNxXAy5WCU/vShchqGv/RAdQawZyhOZry4
OUkqFbpHggmPC9+rV9up5NGa/IIi0ACwaTDlpd3adkCmsyhNdHjjUX0JBRfcwPPX
kEBAqYo12RzoI9uF8OU9cOL/lsXpBpQi5r//pTiKPV8ZemzuQIokwPeAp3Qr8lCj
eCKI0iPKkkYTkZbk+YhMYiO089LYu1yCf8zD5pbAzCJKVKq4wQLyFrWNCPWmkj+i
WfjFk1nafxExTVW9sV8G5qcz/DP8/4fFu05NnZniVhN0FvY9HTOhKjijns79nkTN
IGNYLbWdzoaBXwzFNo/90ZMIc4u6sPbbZT87woKyiPvEMJToTRGQ5blETMx1KZJc
IWCT8h9SUxAB00oJXsvGhlCf7ybJnG1fzCCIcG07pOKYSK4Bd1fp60U3IlY0r4iv
2w7Rmr2G/FW0J49kcXahFLZj6kDAov514UH8uJyngvHgs6+Ne0LWYA6Jy4jA/DQl
spCPQ6EbAL33cddcgo9ZhoHsU6hkIKlnNVwltfq8/1gUAJzVOVaHD87DFbISZyNb
GGykj8n3wFD4hdgO3+HL7aPMgsErBRwJPRJjS+B2ib0/1TcYAO9MCtjHAN1JwmiX
NucGb9KBfN8o3EK1l6oaZ5M1u6aW7gjGMb/EqpeM7/rOOOEMSd4XCfoDIXi4/InB
Ick880n0YbsoZZ8FQJB85EajOkxUFK6dbnI2F1DgiZrL8ajanmZTPGZi9+wNTc2H
iFG9K4qQHHcQNY73n7FOXUrFDJR+pEAACyVo/NiiqYPvVqyEl5Mc8qFt799N3Ehf
v07hFIvoNGxcxBVOTPb8DVTv7dA7vis5m1f9YyFTRUcPXebJjoOwuk7KXCF/XnKv
tGBpoKRpSy7bMmAL4jnKYInI6XrhkPYP6LvrMqw8P8PZ4mjL+TrlmhkzkRRHDLxJ
rzLkyaiXY9/Y0ho4M6GDbju3zOCbn1d3HYXiKCVN7JM+Zd/PpzHiqaf8zDRaxvgE
vuW9WIpFcZkrFltJNaVMRPHgBn/9+Ze5jK9K3yRR2zLPs9KM+2t/NN//XdquJhrz
QnqZh0Nxrmb4IzdVH/xMkXqbrVwC6q43l2KgUYOX/eH9D3ukKist6Nhc+ueD+tDo
37v51lwgspxIS7VhLKX1DfVEarvhdDO3u7QiIuyUs19gLt54Vg3dzJWiVuX2EW5Y
r7At9c+V34VEmkoTHrHpCA+qi/kzAOPLB89JSloyNSnjL2xW58S015lKCiPmXeWJ
yHZ5MkdwMuN2Ir9eME3LH5c22AxMS++fLc9EfAItsKoZuYUL7OaWTNO/pnK2+Mqb
fyH7YjDbaqAvG+4CsufGVH0V7GrpQ8l9w2YZ3uVc8F1IcJ8kfzcVsPniGA6nBV2S
n7qy+uLXgOvk0XHoilCh+wLm1IGrGjJ9n/5LykG8uMyY5RbSIxDOBbNPoTmVnup2
3+2SeAUJZbQAUw7g8rd35RCGxYE0BqJcRGLCbTcj060MSZCmF5BCxvxCm8WyR1T4
Fbywrztc1c+Pqirtw/V9qn2ig/EoXmey3jpzLR/xtXECyARi4vAQtciiEI7y77VL
+Kn0C68JAJXI6sKMUd7R2p08QFu1KeZr9OfMSI3CSJU8XHlTbMnYQanKZKpYQhxB
e7jHDxawZZiZBX6Uiq1ynWp/Ysz708PHz7u3g7LZSU1GNU/FE1c0SZw63OwuRhTR
9O3Du1VJMAFUCwLaX2LwA6qQXhlBezMPVtvnpcoRyUyV7s+sOrDj2W6OdsdYdy+J
H+32f/tiZuLZ8m7NZYF++27eTnQnOQRjIMdHDIlYNhfQlE/kbvYpHh/ab+o/IIEr
lyn3UxJ6ECuVB6juKwv3azjO6TH3+4Mp+rHjJ/xW87OmsbfZVzV88OpQuRjtxpMR
T3YwvktkTeMXBhmtRNLv0t4X/5ijlnTurufax3oqooKCNbcuIhNWNWpLjvnhkZ8a
yFcDzkm8iQmwL3oFVdO/TUjb8Hg9XbMycMH3vZ0e5mWFli+SftkHIQRv03mG767U
wpXcaN5LshnCGwxqvYxArB12+TgnCxeMdgZHupq0aRmuNctcGUzaCouvjrzOG/Du
yUNuqkuxv734Fr8v8/XGdojReU0cjMddv9BE8nIEugmjT2/QQGtXm538vGKFioeh
e6c3gJiwKJZajS1qMO26XBagwNRiOnKYBqXA5zZLAqdoXNnQu6IHGVb/OYB+7qcp
+QaNjyjGbqtAQAiv0QAmegQ1zILDANibINWsSJRJqsYOBgWIz44zG3YAv9uPZGyl
nvz9DcFkvL0OvbLBpqcjaPSEXV+7pIoM0bCEac7qPyDguNoWnLZmcgQHtSKWzumV
8/3VNXtK3YtQfDJM2+PDr3TehG0LNr7FDu9d5v1nb6bfkxbrcrRr78Entb9Xp3+K
hydUg63IXd6RjsZqo7Jp2vK6SHbWQd8XzLfRbP6aGGUCTLTaavC7Z1k6eaQwiBtK
EwagVyhqV2Dc46fmGmGA7yGXRnljFsAbJaiikm0lGf1vkb40P1QzGnScuRuqXOSJ
AGv/vTYX3t2EicS38gGaTzuw44Sz3/CUZUp8tW1kJmJqVR7dZHb++ZZ5LjRZ7lNZ
n5oiLBveYDkIDcxQUir3lQWkr9DjjrlY9zjjqbnf8lPj3xYmwXxmz7H7mYcM7B6C
J5y3/v+IafmYlVrV/ucHt8Smfo4mGpo1OID938SfoVa1VyuhZej9izb0LWOqVoPV
q8t7pRF4tXq2GgcJb9Up4WYhtMe/ND18cP4I3smJ99BiH+BU201tiZjYSqolKBeh
43xvWggtrrjvfF46KL5E0X0RlCfwATqsIfSgcLcrBk8wT8/mwGIJinhBTYKg1cUW
+m4C6T68yiFGMKM2Ub+ZxNQ6I/pXCqfhdjQMZQdrayOqX01qX444aLoNPOW8Yysg
e1lshgOzOLp9XaeL7obzcSZBrLZ3kVxPo+krw7lcYIj3KcjPHUuRy/M7wjSAp5AI
IlJPz2Yrs2Wszlf9KwgpK7e13i83e1CCIw48BPMy+5V4SJbTmg3JjPgTm5LOdC2V
/yJQz1HpF/fr0dMFuK9lnvGc0Mgzo+3LJwWH3ajp/y42TxOawxL1YY5F6/QNp6ud
464hWBoesdv9iz+713cibxnKwom4iLRkec7P2nT0cPu6wck9aQEhx6HQ0aovBDIu
EAHRp/8dLfv2qWgDZKSLp0mGP5X5U4od2VoT3A60sF3MFOAfuK3HRAizRU6Eh0dL
G2fM8DMBxycP7CVy9Le0RA+8EbIDCR2cwHgS7pLYVpG7ix7ub0+lCW/cetEIELEr
8J6nbvrlLgJueGkXjVv2hYua98KPxON8WzG2iT9o9pm7oS5MGhSdehyFqhc/MDU5
elsqHNGlc/fPMg9xxd6fUhq1aiXJNLncIjJi1EUJ4tL91hIYXvQvNabAb3h8Jl/t
CAYd44Dt3tB8OzJKh5cQ9hNCH6kUL8lxWYEFKFm2isK/teD0ehOlIF2sq1ljFW51
2lx8HnXJvz5SLYcpQi2EJ7eHcmgeiHC4TRdm18Q8fOa30KO8rwRZpir9IJat3rYT
16NyHvQfHPXF7eHT0d4foy5WZtXPM5jtuTff+DGnW9OqL3+68974666cMA6WR1WW
a+6KgRW7pKpuo8CEw1QhOPLRhyy/xYXRjA0Kyapa1dpJC3JyiU4vp+b8beaOJTgs
c4e4vONikRjBgnjxZQvzH4unaFkoBDPoo5iA1L3PaEZM9Q6e2mCvXLnp1laKaCpG
lXGIdXdfM//ww01qNNPYBRJeTcMlhIm7dSSnfuPya9jSJxhDHTXR97hPm9vqsFFx
01d+nh2oT7HSPaVylDPixkDnACwrMbQ75QZY/LvD437g+ICgm3sG8lkKbUYnzXld
FFkLyoZ18sh7g+Gy3Es8CYJXmryrLU6/WI5lyg7rS4VWYh6jNEY+dToQCIrNZ0ws
NBv5ddSmyTrndkvzTazAesK4IbpG5hDoKtaMe4MwJ/FhBqntzvcRwWtDU+SOazLK
50qEF82Cf0HVeQ3RJtVGN1IA/acRQg5GHdjzACCMs7/hiKaplMfCoIZnzW5KeRqA
76eObDnyIFy+0tM9OJKq1jDA2IUnVKsD/K2WjyW6ZViheKlXeGIrf7MJ1oS0YN7C
TPA7bkOATl+VAPYnlL+y+i3otdoxv04EM1b3YXtT5XH4AppcC63RmAkWmhd73Hnh
e8lY7LWDbvnpUTlJci5hnM4Tdm3BypWSaBMs9RDdlpjkwETWkTlPrfzshEYi0Qp0
PdOQAaMHzkgvziY+aPoYxr0jPzqUEEL0nqgU1+1eOEbqKHTWY1Lg8fC6YK/UGsE0
zdSssMN6kW1lut70zPc39T39sYn7LcltFMh1d+/Nk/OjL9FwLBS01yplhjvQ7Hai
gg4ATVigJP/nAHdwerI+ZEiY6iSC/DOCgB6dob9pn7upuHkyNllNTlTohfwBHqkr
SZ3rN878cwPwzk8wZuU0e2UdZIjaLv5uSXaKbV/2k1nRcIXdTp54ms8rqWn0RFEY
vg/HToKMhG0yEP6p/yvR19+Spn+Iff8ddCkW755rpL77fdjUBOAWcN8szlUmhZTA
otMOlGkfWI+Q0HQTou9kPSLbVwWXyGJU/Y8YwJL+g+V/tdu8I6OgWfOMUu5A9ruB
aXoSr4aCAx3OSciag0QOH3x3EBOZ+Irjz+erWORbQAcBfsosH4XCjWdnNrqZzhjw
wLv4GJuPYNXdxrQSr2Ta8p46+okeQpID5J4i9PQJwkYcPV2kgG/scwS3EkjINncv
xS5KpOXQkxiCeX3VTgpK109HnzmXOT9P2x9aPPyHYMiqZdBDe3fh/1LX21KfPVve
CG+G/WmmieW8MP3YKKd6KTEjcpYE/WOQyNNHDOTFz2n6AQw61YPEjQXAbQZWDEr+
NgIxLZqNww6iPhtw80zBXMgDvztIirACntBSnJA8D74pS66qdUdhpmU7ueRnKhnr
FmMwIxewu1IT5g/E1a5gZULaRgxoRH8Iq/1VFnj4K0dtG0sdcswpy3HCHIuQ4ePy
X09y96KZrXUfBZsiIUYU7nB3G7+PgAepwcC9EHlQoluyMzJ0pNbjrq0uP7HvquSy
mUuzzXQZXArQZ5NiUas6YRjQ6lxWhcY0/FEexpvGOQ1On1X7xDQnLc9YG+zkjpc5
LRl3gMIpfPJ45GjP2zaJykp3uLcKZfwZnx4vWQ7OCeGNcLxsj44zEX5ITC1pI1w/
mf/hX4q6Jc+SJbPbXiLRVhwNcy+lHZaohGOrnYvV6YLRjoELyqHvnosKis6NhhBp
jfs8wFeGJH0vJW076+SmlkicVTecBqHF58TPE2y/Tal8bdbTgqT71a7lZkK4xcal
M2Rm0R6Fi7WC63wADY4ZfstU9sqmzoGvuo3Koa5gvh0dkn/2a3PD8svlGY9ARESc
eWyjBbPRaQFfY+FEXDxTEjVXS/9EoQ2RYcpABfGbr4vyc4T+oG+b9Dfod0yQwGwP
tPPf0OKstNUf8Pkg4+eHVNl09e8buZ8jr7Ud9pV+L7XUVWH4hDHLOMoVwr9jP/NA
vYu1/MiULt94SGv2KdZ36F8f3aRkqDoZaco4KLE5ZbDtrI0CXGcBESe7NgRgZyHs
YcdjVhHzHaN2cLtQ3VY3opMU7VhC21sf431xIs0EiIp2AMmruGnk4eO013Gf7bF6
XHZsp3xM/q6+cQbEpEzMx0f8b+IeyIZF9h4HJz8be7MO2jjkjjNKDqzES+2wwD6h
FlDuotbdTP0RY9vXKoGAZbE2LYWbWTk+A5x4mIwTUEN3vJPJ9KwPmrqLoH3M4wBF
rOrYKj6WXQiMS83as8wB4Xpa7IEsQtxPRek2tH2FjYP1eGAU9RuVGKQI13xzhmnf
IOTam9PNvUbdcuWpTNWmOQd+oZ2uvkrtM+aGpD/Q0w0FKeMvxLA+ID3VVRooZZaG
k//iOZYQ/Ou8p9awL43rez54flbsYV6saFq1Lf9hKVfOgMR1lCCMIsQCcS1Tja+Y
DuAk58s0vzIBzIMRxUaiGKz9GQNMv8ZeH7JZ05/is//6YqsDRzYZ8rIFWSuUQSPO
ituCdaZpHMasFXn5MYCiOwZKq11q3bOGoiHKT8PSNpDJTogqUMd+bGZYNorXKYuY
5I1qPUXvzXGtJ4cblY5/meeIS7NcVBKySsOQGdWoPuVaqWMQkbYmgUXaf7k/D/uC
DyVFqCUTuIBnuP6d1UBj9uezCxB9o4wm3OKOTmLV6wCX4AymFxnja+Gg/FZAXUN+
SiMWR685HsVO3m1NJrd90Xw4bbeOp0muM3kxw8I01JRk2IymVT1LgZRXgu8pfy+f
ttzhH7wpHBeFDbioIQYiLOUupvAiEgPNkSLoQq/OAFtvmAMGF9clAp5xPzHvwoKM
O1r55qi66DlOgEjePYvl1c8gLfyIT6ZW8VuFfNpFZp/UjkkaNOqkY1NVcVMLj1Y+
95BjFmjpP2ILeTqSqPA24so1tJwUYFiVQ6heBe1IRh4H2ns9/NFxSrRcXFgxMnZ5
ugUr2lcuUnTepiW/qc4kxSFb2pBES60uo2gGHFXewxyQ5BgdWCCRbt5Z5AVaW/mW
M5fBIjhizBHB1bY8nAHz0H4QDyRPd/nE1AvZbsaKWuIuIJCEx3IemBUGM9HBMsSP
NqB5X+hWr5VyX93ltkyhpUm2v4ihlYIzxTV1lU6WE9AHpKxYKHVW1kshihs1qfOV
ajZhIkcBnD6Z4xRODksHQjwMcbBbhyLZG6uqWizThu6PF7mffI7PBkefIt3NbXRN
Qx1OrWpz2J+4yT/PDTMOO3jSaphGW6+rjTHkiVtdQzkqrk0P/m9B5/b5clmAby3L
cNcVgL8Kfw6qWZV4TE1/8Ud72U9z8E6YKXL6UTURlsl/yT10R+/BUX0RdhIX6qWH
QPcvNQP5LHRbhta/oW6ytXVhaS4n1KfYy+YqAc1Sr6lB1ph1XW1qni0R8XiEepeY
igohnqsUKnt8cCm0s3Msjry35fWzNpYPhnira00qUOzWH5IGJsm0P72z8wKNbZ/z
a48oYrvn+GXQo1l97RCbzluZpf9c9JHWbZ7Ii10AZtsF4zXTsbtYVuMC5ajQu1K7
/wThtxUiPM9xdjf8ifLEEWhSJLW/CV9NVBwpiBZvZ3pLIa03dd8eGiWWo6rRYB2A
E1LAsDL5fPqcgL6wISvuyWpJYwW3zaMT38eVS16BJ57mvMyjr6TGFXmKuddoOAvV
IxJphY5G53rY5OWYSYGfThs3P7xkV4Hfhd1z+FS3YWAZ9gGvoq80a+WCxjont3hk
GI0FUweYHza+Urvlp/fibOgtboQ4bA3dnxXOa6zE6EIksEb4leOmTZupDxkn7Mv2
vN1Dnjo+zCan2BXBPik1XwDjM/GC4WtJN5xFh8wrHjtXUnBNLbO5dbVxCj4cOWhm
s3lXTdLGwVf8M+fmcoEmZsoQHehjrfoyEEV2eAfjCg1f8FlTJ2LqnGyBm8De2OoT
HB1nBqbqx7TTShkJgO51asadZJYI9eSs5MPU5I5pGRMgDW5KPHVvbpxM0Tkq2Oli
Ezywlrti2pqAZMLs/2CDd9OcXIdV2sgvqsevO4lPPMhFbegGprbZ8i5AuKTl7uro
dBJYrKNLgMxB8ziLu+Dnn05YedTSeAu/RszICHB+sVd2N9opM+T9miSIQlE30Zzo
mydsQdokpejeA3PnrGops4qg0SF68Bi/lk3pAmJUzp7fiokRWBbA0cBfNVMRHyoO
PqVsOhyNBpJadH2+YNSs1kOONgp5NCEWN7nlt6UBVMdONsONADV573OGF4zihkGU
OP4Ulf4Mo9MposxGoZh8tN0RgZTvu5MEHEydHxSnQLAdftQtRL5pCuVi9fhq8JqN
Z6ZoUvGxRWK88yscMO9NkUexJaVLZaGfD+KYdq6spCG3cfNHcz+FEIJjxZS/i5h6
Ut5gpIXVXqb8lhXXhgUkAWSVThmtu8OO6h3DSASPeBQIh0OfLGTiRy3+4j4I1EpE
FOOly0VHvhYA7ST93mNA5/Gq3+nmDEaw1xsktZvkA8cafNdqpGimtV1II25ysVkK
VXDYzRju5dau+ZtFURBNSP41kx+5R9JzTwVKb9C+9D+dxxA8IwfqVowNwqKL/p+9
zXY/z2TA5RGty5BhP3gBbkxDXyWWPMlk12Dv5d6LNgiyVoCW2PNSBwTFysXAH6UH
FWkiFeyVVkBwn5w0GVhb0RVzzCqB5Bc1IVXnUI6DkrKNe9J5NAmQf+HtJ1D8ltmd
pSpgi8tKP9HUIsc0XX1rZOUfbOWy3QHWyQ29JY24yUKve5kI3Y8rOfSd76X4Frem
jfvqTxxF0hoHNcD9QujZTiAXmdHjd0AXyJxq6vyGnwKjylD5L6FKAQmZEPpNP2VC
Oh3AVmdyEBcdXrlGp6ydJ4r2o8o1Z4wj2duVfTr+gy3gQdGI+YfqFbSBE4su6/SH
HcV29rnKSBFrzjq6527QJThk5NLLu+Lwn3Dfxy9hH6jhykehPYfJA6befbua/dgN
xmBHi4bTg9J6w9e/QnmRNCkdUzcDN9LqTkRyMhTZwqYRVDmytHumICO9dNHUmPO6
xsXQGgA/EWM0nhCO3Ufa0gHIFlxcjcNPs4YoItEujRvAqdXt/q7trxBcWRvzwvZn
cEmfGDGf7lFOBBftqFSpo1OEQV1kM0B8KtaskbHrSTq+o0HlLQBPs4P2EaWu4bpa
IW9ABwxNDAFr9iaWSc38vgNf/czivJiXDATeIOEB5Q1Yygkve3npcKcwy/y2s5+b
x2/ZRyHgmqjznZQu3YpSCpNdAJWaYjHk2rdOXaVRtJkWTbhOqgrJBu6/0u/xyTPi
MiFZdwWRsDhaNHyAXxwzM5X9JLfRUG8uf9g8+RoJat/C192bNVSh0g6cyjepTQBR
UaOvLe0y/EUbYIjpBwuCHU5z3EI7tMEkGS3pvZMo8iC3mQVwEpDj3lxS/V2Qzcor
Q6WhWgfKBK1gJoiwZlYVp8l9WzXTDEQhFX9C2AIMEpVYLrsqn5ZgYG4zPw/h/Nlv
Fkc+0kpIplY1MfC+uZ+MLRBWCs9KcM3Mar7+kXmyhc7LrJCk1n6bGN2Hcs4Jf+3l
qR6d9l4RGRVGCK+9Di0o6y/DtOQopCYK1s5uEkI5wjL7hMjXFKdf0Oiu1nW4qDvi
jqnQQwiH/r8h9YCRn/WY5Fj23y91vwukYyTZhaD+CbQQQTH6jTYYuTv6uHNdW8j+
ZidSZmbcNLnUpJrCarmJZ3k1e0ARcL+mepiCMUF9ojzoI11ILK+Xzz4lN4fRYuy/
ei0m0y6rJD000Pj3KlKtI74JHjy231oRCwPbnmJRRa6U3DlOmQ40tmeGpEUpqFp6
EXqcNvcCC0FtJWuE7ptJD8peQgRxfe4RRgDOhaMBPUA1jzfmlc71Qbg+7ZN7VZoF
leGh0iZ6u3Hb1eH++dtmk1F+N/gcdZGh0xRKzLXhotDmWgYvbdh5AbLLprpkPyS2
iy4PsO3v2Ncai2X3GJVe90q+E63cRcEPv462pO5XqRAXi8gYHA40doX5XCZIKjTW
G1GDiaKikEeL8fX+KWd4SSDpofPMef8vMCixl+8CnCDHPFjNA2eG7uS1M4ydxZaW
d/rxWQ1T10AkW3pgI/EVeo+YT6Q2WPouYs+tLfcQy4vE5NTwTrp/cuZecpLf7zXD
Jfl38bdPCiPRGMUQbyzitQUFR+SqWkL0+TlC7rb3FTjBS+A4x9Q3j39S05Ej8b0x
Thy3gfTm7MX13XEbwe6GaNOdqpHkCVFCvM63FjJCd+d+05f4xwWME68XKa/RxvhK
TJsFGty+rUuIA5Jj8ur0pbdKQ/2U8t2suL518bXwLNbTeYPxLGNLtWdiAy7vjMZL
n4NtgN3shaNZSlI27LJNlC6KwT78z9rAIZSHvIPX+lWzh+289ypSAQWXFClkbVpN
7EKp9E4zzWquY5LkCaI3unUApJ7DC6RXxyQfyHr6Zs8lbI1rM6+ofQxvt52tCX7f
oF8an9HlMpstJgMJt8Wh7SeQWdXVSil78jZs/iivHrS9SM8x8xzkCJw47C6whp5k
ZiOzfDuBrbb0C+ppcxRb9uu5zq4UxDK0RdUwMGsCwM6y5mmqp7vRMd92wPoMz7wN
RiNgWTkJlqY6Bg7nzfCQ0Mjhv3JrqZYamDd8kd0gMW59tvW3FTYkJSoH9exXTjIB
NYRiAQQmWjr/9dfrYQRsqpMHuLBgktjAGqZ8NbX43SWBcYbj5E1u/uos8jTxcAKT
o3wwaZ989OT1kcQWTe4bAylUPg+NE77QtiBG/z+YBssnR07Oo/bS17+QCDFn3UW9
w1XJ3ys4nyZ8FxzEMkXYWW/BO0mq8oEdLE5mrHv7us5CDVK+KDt2NVUM1I62dWqt
m5+a8ol8cDWsXMoAhy16e/ofoChrZF1Uc/F5xDqyAGsUWpR4CoAAzeey7RQmNZLe
f9vst0nvBo6pQceDCGbneKmi+9mde+8OKF2koRZtlkIIg6/eT9CHYohcrR36KOo3
ROmKrR/E60skccUG1KjdGvuB3Od9Wj+GeP4I6YnBBVdd+N6CzMojfq05Aj+ePeZs
1t2ITEfggTOYkp9FXVTfRgiil/tljSzwqsfepk6uRwD1LQ3OQ0WfToizAtR6nT4z
Cvn/Hzp2F7aTdHYLYr9g3ChYNKyZC2bKrYOJaAWSVEpWpNEnvIYrg8eO1tPdoqWy
F4B5bMj+6TjGkJ7oXdm8w/dQmfioYJOvyH/0yb2IS1GiVaG5jy6I+E9kFpSm9Gkz
ZnxKLbd/QaTUhYyZ5cw4LbYpDpATekvZtIkT2ASJ2UA1INeqYrt7TYYPqEodHbcV
efhK9/+QnqkxDMScHLHWkaxtWukt9a8UpPOXiRZG7BkZlPaAe8gtq/nwTzVL01lS
601qDIooI6/0asGFotu8hVQF4eOyC2XOsmj/A73acul3Fpzu0aJSH4f7nBXzbZii
iBwxs6zEzTk3SS4dTtWKZ5wJ1PkBfyXSDBfWMgJD6qoW593EtpGC90svs7gHdvxk
JhjbRUiPfN1LTfE11nMbW2JGKhPJwi/NQ2TO1OsD3XSKp36dDwTe0iHcM2Ug0dD3
uHWjyJjKLMadZj+Tx659MP1wtVuA+gJLowvEbrLkSdYq0YtLQ4qayPemWXc2FHUG
UDYamvzkA58ihW1Ti++kYU1F/95kglCzB4AIzm+UXfkTsuXI7BkE83am8EjVyJ+t
J5BmzksMh50l3pP2BDjdizr33/VUEMUDYwuniSjJ8AhfL49qTCo2JFMiyeT4xDBs
zTyQvsWDFczl9oOW2dS2/grzT0lQVA1TftatIH7JDbS1/3myqB9gkzVXe2OWmJxc
FK5eO3/9XZk7a1UB1+vNzhJci/JbprLREVFI0oBMOheIMXw7vUXKg10x4x022SV5
i3n/TKNLZJB64fcstaYmXt7QYelYG3W37oQYgs72Aai5ROaL4LBjJPtfqrLwykVc
qZ0Pk22IhMEDFW+MqncMWPH9GMOcH8DbUaH7gYIvSLCbDMaSI8RDC39PdJf5Of/F
3qDrFKIYrXtzsoQx/iYEO9onMb2wFQ0i8oFvObQgVKoWl/ajMSlUhyaWukIcHrAq
4DhysaTwxiiq0GK1Oi3tJiqwtKhlB4zQaGnrvGb5Rhk4u6BolwqcjV8QIUxVVqrA
M1W1R1rWMsshqFfpUuptc0WQcSMIusNO0+FmUvMCaW0kmh8pKJca2i58tVVw062N
K4+VqgdG8Ox0UfvHyS5VB4FhzQm6oQkv5UZVE5U1fk6ol9NRur0gJ4lDL6YPTJoA
aqvb3hjQ1E8p/kXyrZadvq4QtfgsaGR2o3zGOyC5+kNNP4IoqY2Z9UUluGYVgPQc
z6qqOXUCJRc+QSL4Ff+t+Ia2b6eddm4Ed5tcsyMUrZp1ZNButj+ZYpfaRObpreVx
Ia+1WK0zvQ01O7Zit/hMrzo7UkEZnyODVONVCJ4T9cRGF6nmiq6UKzGypWFzOz1R
0rE+AbxK0XnFs7+fpb1JtSrbzQqk2wSLwIEG3tLSaDpFR3khMim7dJHjoH4Gl1qP
V+XrWkBApyfYJkaDFyijRRexHjYksdbuEvZgd5q5uTcCqpXUSMfPh1Q3lLMUYhpi
TGCv7RRghn8KJ6qbDTSGRJmDebtBui6eH8GB2AdWUUHmDJCPc4tcYk140pWo9GG2
nIoiJRLQ2EDRuHLefnBTTUuwUnl1HoIGUllEHVk0Bwy4xQ7DZjKE5b7DdBJLCP1z
b67Kgo8yscSz7bWlV2Q2MUlGh3VD8lpZ2yjer/UCiO4nHte0u5Y8jFajgtjmUprA
0uEDiVKhYh84ooiiZtBmeUbU3aCIUPqueev1vHvfMGjCYmkLY9epJi5TLpUpOugX
Yf4+PRwS+nvqOVwsIrxFMYexcWlvVrdHi89BTom1o3DaTGwBwrjKjv5gpAvCbkIw
dkZbn3Jfaw67CZzMAzbRzKNRDHIO4I3LlOE7i67PIFTdbqc7ZX6IS55TWdQdAWY4
c8I1ozPrfEmVaps7gjlEq0dTk2RzTZkhOxq/IO2b26iO+aEEhesOPToQ6Bep8y8R
uFXCQM8eYIruCeUBj32AgBjrtH7wWGql83Kop2rFOYQW1Fa2A51CkunCiKzUbOhW
Zjv/j+63ie/kx/hcWT2FfAESFdhNZ2K4VizDtYSlZK9Vn2oJLcI02AUl2hq0O8/k
yqILuX+rR8MaMTN69JqAHAElSYa8cre0+n7Nwg14btEgxEzm2JdzpyzOuoYDjSND
WB42a1hf5w1OqEAjFx0QCKi6ZJt4crE2tmGsI67/Z8gEK85DQMQqbqLpb+sgLBu5
m6jhsbvr1kk6v8OpRNtO3i6n/b1NUtACXudKGT+Z+Llt9VCQDaEyTtFSdLVDhD2t
Ciq+YjCcXDgtcJ2X/KS/lq9XRWRQ7s9zJbgxTmJn3GYWQsnARPgZlVxXMOK6j4bi
rMPyTr22FRee+rnng+WWqC0MR0i9WxiERgllOlK/wO1oqWtXoTrUkg90XyUwuofX
B9eXwufqFqEUuMELlSYr9sac0aHd3dK3Qr5y/1NIUyYcYpShv2foUJAMbkvz9Pqb
9TCL3hzwV4HFV3N+5LyabSBtdbrbnhHLBckY4IFNCzJcFsnL9J2z+6/aTur/4YVo
KF6y+RFCB/V6typ6gz3mTcxNQIkWZW5tgeiZJ1yNuyEw7Wkjzj9MyV+LWkLJGULu
VtHBLxc9LkNRrzZEjtqsZavxr6CsH1pirtdQHCM5BuQ4CT0d1tdFBsvUJrgdx80M
rpLTOgVgyoihnUoiQmoEOkaC+lNpKG4CXUptNm/xNZAVxNlfLt1qDjBeb0W8vnrB
13GTfUzfrUBsnWGzb62Iy0fnDCw+fyA9JcF3N3VFd3lvtIglfjoUOOB1bH4jJFFD
b/pf0EaNoRHFPEd0JkAk/r0K0RNrp2z0RgERQcF5lLVw1E4/Xknt2y7n0XsLbtGX
m3ROwr5ta5gePUv9V0W1sF1z0lIPZRDsYkn7alZCd/X2Y4xtnJLmbllCnyvR04ff
CTbZBl2kgqaIVIB3nukRCiBpkkwCSd9KPX/290Htq60d5Jy1M2v195q3JF7y9tWz
xQ1h1Nn33rNnGy75w7IPnLGJS4vjk533MsVzlwOufgvz38e0q1wDVJK3KdslHfaE
wMnZHApmLOv1dBQn0cZjF2M2VSfncTyOT77p39yBciXwX9WsZ4rGoTuFJHJv2iGE
d1nHlzEYQ6YR2PrcDDHY4kWdzcPJKoZTN/ozNEcln/jQFAerAXLj+aKN1SpB03h+
BkFjCa6mzFq1ijIvVkW4CjmI01PSwSaPj7Y3d/ZF5udvAyng1K5W2nqNemPevGP3
nhjkhtaRu/g9yKbQ4OMPCEUS7ugq0OridCQKjTzjWXapQdL+bIMsrJrGfj2kIH6l
aV4lwqlsPjo8BIiQLe3i61G/uhDzjyqueiB/89OGWadQkTCrKvlBNDGsNuuYevCj
cbnSG9QAX+KbPOmNlp5k22kxl6xMT/z7sfw+FWsOketsgfG78Aa8u/FR9j9WAOG9
hpAD6fszQTHCC/7G5A8RVbwZDvbw5QddsHxYnqTPL1glQQYUgkWDHdHdGjh+6dm9
zbmijJc24IArQabU5rThgu5CSz6xq3E2vKAUTSSXXs3xZ5cAETzkvUvuLZWf2Wtg
fUxpq/jNsnbzu8qMLBt5RsRds9nys/2mqaQ6r09TejgITGXyGtgYmm7Nb91G7/Px
Xi40DcwiGehpDNgkNEHAbQu1NPnOWzmA/COPF6ELm/urbZTxU4DNsHb2NnScZt4u
LuiqO7as4r6tcdBPNGhAS2aMAU2OrgIMiZHIlyl0qrcby4cKg2utPJyJozSfZOWL
sfdvRcrI5uc/h8dF6em4uFueF8V8LfkHssM+LHNZ3YVnF8E4DqXsQrIzAxreGIoZ
TFZXfNPg/3tTypu3qFXpynSJP1qVl8f+dsApzL6MwrzlqqOpS2UXiU9T19N+Qsue
Jv5j7esBC1mPMNONWkdtR7h1DBtjmBtlFpYR57vbVsgzIyfCawfkSPZlC7VdU3KK
QYLCDEPErPNblmtr1eD1eRNhX7Ks6Uo1WEjLhc10PpK033ZLkZ+Tq1LjDsKUxyX/
c3DuEKOX9m4FAXw/i+2zx1ygs3iTwnEG1zuKv1g7ZMrIWIly+UOT3gWTdCpLmTNv
n+c5WoCmxq9ZIroVF+zI43sieq+qqoyIUVKdXKr8UBMNCabiIYJLIs/tX+bq5wrR
GOxB1PXukzcU0SITWP9qKrqtKo+c9DcBT1pXSUijjk2F52r0n7qwtZhZJVmGyaq4
HBHdPqCAtRGVSPXwLoGQMdXKuGHA7yDZxnEPHIER/TPeM2cr6azqGVuaV99s/Thl
0DR375jH2tSI8ZZJHnSogu1XAnM7zQeaJxxfYwFLMswN3zVXpOrxrSOr7VqvR4Zu
oSLroVruEdlb63Sm9c8sa7wx/xSAWFYY44qe7vSTAx5Eqnna7OrKBlb3VJBvw73K
JQa9z/Z0muNbXwbmSJqds+hPfDIglb0IUAloqi8ZW2qHLQ5po/EQa7c4rEIeKBXQ
do20FhLOA4r1jVpkmhkQm9pQbWLY/rXTvCRWfUZ95OUOSWVLhvmR0zXQcDe7JPI3
4flwNzaZiUDcccXsPmf3zeXpb1KBSZHq9ifgZG5GWJtJktv6FUGxndAzyhBI3Syw
ZjGHTXMYyPP2tRwL0bXaFmOXYjFsqcgfWj+FxP6m/ot3zdqV8orR2s/VZEi1e09X
0O1RE4ANRQglxUGKvQCqXSaXh+LGEVjHpfO8YLYDGrnKghDomX16wiD+OzU6Z3Yc
tQ8j1E4o4iRwzaqZ7ma6d3wWvzHur1C7B+KQPwosOTWpB4uFqTDVqwOwCAUxl71I
JLOdXzx2wh6D0r4vhzEJJ+CCsGZxIsANysG1j29iyiMrfPHWkp7ciu0xJutca94t
taQ7oIxt34hcP3EHXh/eGAPXfDVaNSU4Nq2TQ5RlCmtfblT35Fu9ia19NCrrW9MG
TN9sTVdbnJoCTknCn2ZhtxY4CBn4285yybPVtyraReUms9K3sfwhDtCF06wdUvz/
DNMh+TAQl2McT6NXlXdat9lrJxt8MaqSEx+e39Oe6/KcO0+ro4fyjtrZN/zWsHaK
C+JOfUDBCdeO7i2K8PXEwbhVLmZZbJ8tHFugtM6uy+SCIuWkIXQ6KruT9bJ1A/uL
o8W+9TjnhCd1QuoO0vwPlDTkWeu/wiSLg+4O0S888elssMD3UIdzvLBT8ynVJf41
z1FCIpFmPVBIRltMeVz1PdwEl41Qpqae7zD76Jxk2z8pLjMdoB15tZpTNMEazbAX
W0CMd0li9HLcE0Cqk6sCqIbHsQMME+ZlmbmHnjOB0MgBRAdDq0t2tEjgryAWWg9E
2QiuY1dio7uacNMp35uuh1iUJp/Y8iHPuCKVpQsoeg0HpyxCAmJYsLId1b5QtzBh
MksIwjvpcNXMKZLXmmdTJducTttJiAPYKofh4nYHqGRCk4stEdJ8u/dUn9LpHMDx
WqXEc5O6ye9Wqws2FSIpHtRKPhTb018pCVp2B1g9FHQI4KKVCcendxZGpHPy8Dkf
/a9CWKgkPw+VH1zsWmhITVEZD8i2ojKs0bRHHcofSVp9CAZxm38aYPIv2ITM3ctg
ENbW0Ty7iX3NuA5jdCVHQ3ml9vBnmTilOaQYHbAOTzuXxa9BxdBdKPm/7zvd0/Id
0b7bVcIfAYt9ZWl+oQOmYjvIunMmwAVk5h9lBx33kcLnkSXG5VG3UcEGw0u387Hs
Vowz+fRKP3CN+tjAihRd94EuKVIGa1FFPfUxF53rPKR1C0OTID5AAwnB+ZlIeXjC
xB/LDzdVakLv8L4qJk+1nJoG4T3P79cn2CSWRVkM/9i8Y0WnyY5btEwzAdKu7hZH
XuIzEj72aIcz+Bnm2GKrR8e4CZmEIzN6cZ9xIA4NgoGeMCFlKd+kBE9BxKyLD21R
W/Oc8WXvShkB5de7/lu/sLnxqTXpNq2Jso3/gPzpAOFzoEXytRgCIPfuaHhlNBjs
CJJ/mlSJ56NMQT5dK0tAIXJI5m/qyMlByPNDiqazsZv6D7dRYUKaIXkAqHfW0uqT
dNHruvRRX3EP5N3y7kzPZoJfnwX+RTToUcQEHcXydDVH/V4QvVRGPVW4iZ1Nfhn6
hGp0Pn6UdhC5ydUetTT+/rqNEnLOcsL1V3oclU4SvHyJUmJBB4U8//0JlAALuQoC
sQTRzw9ocJULM0Qindms/dKVI5N3gSIwFvSg4qQ//M9pn80skpv+816E4HbQ+vqf
H0X5PLzOTUfdge677XWs2538RIl83oWSrgjCgBaKB/1OeP44d8gleiIJryqy+nGC
L8VyiL17N9uIX53wNQGtDLcqPTZ72+kDDU1VwCKMQwqVgiYtB2aIUqmLlzhGRHkm
OFMlKIID3SfOLtfC7BgizQTyJblKuk5ETY+OUNHr3FbNKekYWsqi7aCt3KRShYyw
spM2uC2b+K7ziFaIdfr9Jj3e8HCWPB7clzUa3D//SqSpbXkg8wrkWxKs9Bg2CuOY
xv8nGeHHifSxZCUvpHEV9Z62M4uYq6da6x2BgC/Qj49C3+IQOVtHa/5l4kIqZTg1
ywrrG6n4yIevr/4IfMNy58cf4ctjFNV/Ex8DeifoBss/7mmd8qyaO+m25DX/Wu5C
jspTS5Rt9g9QwSqVt/JjXmaiZGfDv6WE3ogDtkaYOX6RhvyCboGiVyTiISBUrGJj
EsE1LkU8uNkmQPUglB34wek1phom8D9fW6oDzxveFnygbvBYWr66+079VyLSsi05
X6q39W8EfYf08vaXQL84jB6gAr7VJGMpP5R28XE/g2OxOFLhT0rebTiN7mI8KFBh
kzLT7m0wcP67M+Gk55CievnuTnyg8hKNSrvrJ2jn1TPv1Ff/Mx0h1ggt7ab/32ek
+YIdEp/qn0Un9no5pGiAd9ZnaQpv7zgh7Mz5J6VJdfRpqUmWwlMnc595sBqhzuZz
FfXw/HkVw1pAqVzcsIDGWff2QO9nBmax+gtvz3kyI+rnPwQrHmNn61k8bfurlD47
81ChlzP3Xs6LlHkH8Sz+N8HxhPLV1PaQxfP73eiOrOOAN06F2Iqgw0Z7bGHhpE6Z
vuqQcYtuYUnkPELN5Y1RZRJZsTvILyC6Si+nyLgu9NEhoo7DGsYmC0VAMNm92Nrf
35Fsl7XXyHfN0EKNb9y6/0lS2BcN0XLOmxA8Th1vBkn427olvYqh4ttLZor5Yz3n
J1RNodFIfBXw0eUBFgJ6T7Ab/8T/2+oVZ11QnOxo/5sxJFMze83qdnjeP5TsisYU
cZE2KMDECAK+bL3HE9Xq9ppFbxMD/yLIUcHjgxtT8kGMvpZ2cjYewt1vknhxRnUt
rDbH9PKpFMZHJzTu9G8FbTayGzCo7hCdX+YL485ter0hVwSw0FSgVp/19J06H6UW
6bIWuumd3bPPF+d3u4Tj8GkJy8XjQSbJx4FmrL/1fQ6YYF6GVA/CgUCDxI2wYRwj
yVDgql9ENxgc+UIdeK9m+aJ6un0EjEVgES4Tn5UM9A9vlHTouPYHAhbQhqKoyoW8
+pR69+HZJa5YFc5r/JWMxhL8dJd7Zr/X+rEdGXK5UAP9Z9Xh50Gz/m+zDAJMOUXG
1s6BSx2JR8V5nQXuZtBZ1Sh/3eVXqy5/5s5yGJFPTDk0aeymZrynLXxjoQMoRGn3
y5jS3gkWPouGETSqOz8vAtFWn/YzVkQLMI4gIQCsCc3aqkRFgp7jzeWPz1vy5PY7
InWq25uyTqEdh1Ra3+JBKRIl9lM1USHRqz/3akwjpXHGoDwD1sZC9EGUtV06A2lR
HtFGg90kgCgZxW2jZikDo3Kn55ioINEWSqSNB4Ip13nEEjn/texJmgIA5ehJT5me
5HUkNDuSu836SAnFrvrLjrqL1kv54lrWXF4Y1+cU/GWokXrrOjOD+tHMT5Of1ud1
1hT+XAAUQcgs1PgKIZQfkz8REuz8I1UjBPo2utG7LD9yum6A+g+SB2cNIi79XHu5
VGN0bCuC6s2bJehPmXfnV+yKjkrvObaD/T52QqoIcP9cCwxMbQCVPCOjNjOAdbFp
PhFOyp8CmnnRbdCFOUhySXAxn1pob3N+Ui+abw4tgY06Fh4OxE3KRXEnA4vqiNZr
wS1jUd2y5xV59BlCFn3ZhG2fEwnJFqT65rc2hSbuTOQKmXErmcbPTL/3s+dkzBJ+
Dyp9PxVYGmJBy7hwF+iiSUIHi7ZHJw+TleEnK0a+KlNqMHYyvFRRpXdeFIPEqEKv
lc7lAnJuHzIhtHqxJ/lRdq6mCrSzsbltx++oTZ3HMPC/2yg4VCnu7JBlPufN9Q1l
e+0cdP07TB7MJTQKtsnaURKKHNtuUEb1/xr5UqY/SVq6QXiMf8eJfdbQ5iTqMbNu
ZToROX9dHfAq1HhflwSgXRk68L6iw6gZToItYO+bP9LIgd1ccSezeFP7/s1GK3Fw
O0sfQVzy0y8ZkCwC39Yg5AduSMrNxLZn/cEvTNAxj3BeTcDRNb6CNK0vSOTuxz3P
GOayeXyreNiAUvFrtKqo3/1kutodQ3+zmPtVEyeINW89fmS/um980GLr30qZLFQ6
jwqh/jlO1D3X50LiFDqTwxrOIPMdLE/N5ZQgaq+jRausk5FVsTVaeg01vKbAYAOi
w1kONnfPCjtv45GH/k8ADpfBF5eeAcvQzqfhJatn499Nvibr3bgiuKSRjs2IRxR5
ebiuuIdeg7L1Ct5f0m7i9n/EVn9novbIojoXRtsrsRqSzgiZ5XtVjbmmvb8v+gDW
6zW0SBGINojuCtYXQ51ocxsO1rEn+MZ/OoMaFE+0RwPlw6QUDbZ9DWlQ1RWyXVPh
UUKVGxfi3H0WezjPAIP8K1EVyh9EytpzyPPhfXelvFmb1XYXS3j0oNRiuqwHgO4G
KGCKKschv43oX63e/SOuwfBYdRr7wOT/Yrw7FRTbBqBh5x3kw9FqgTts7H5pdyDV
fQHNK2ZNra24tW09aOd8MeYNtBQbQ+2R4/6tU2DqqlPjVA/6bZ2RIJ5R9onMVI0r
M8xgK02L+ZjCvGcCHkxCzi+Y49ff952YxOqLbVdWk4WiQfcJBLr8CDjBH0FU8mTa
mE4FS2/P8zA9KoP96cbJD+qmKsz1CYSsLvx8fZvYM2IAHwrbbRN1Q7JmZphYR/yZ
wpdQkALfHPfsFsswTyPCR+C8wfBNcxbNLfoPHNzUpUUNGC9LN8MzEcHma6n7h11s
qAxnlK3OB6//89XS2Trif7Q71ltHRgNpzLMTuBks/JX8UOTBfsrkJpizjQVT97YN
tlcO860jVH6YMK9EJJzdMNKo0Lx0xOQRWoNWHSn6g2vJ29NZoasfBm2hlWUXyL6m
jOVsJKoS64L2MWCXnZ2fLkUizV7EK2zhI+GO3Z0zS+oejFjJHT4WYQLq63l66/3t
lwVtlQBCAe5aGKE1IGFCOjznzNww/LbA1Lmz86ihllRvHIVqGrwVJQnU1CZxSN69
WUMD09x+8wJIfKrY3Cu77a+2Wzdjb8IN+VPrX748ofUDn/R1YYhR9oUPHrGHxEZB
H/43QKODdFComiX8XOsOTeXHoqs7QiAJ8jM/h1ZUi4m1U/kzLeyzA/rpepT4sUJd
79Iqfwm86yRLSYBGBqaV690+LJnNarg21+bZeSLBVbXg/sly/K7j+aIZ7sDC8XfX
Ps2GFQ9Q65LSvbS/M3dLOJEJ0k2ELQqp9RtznIp82JYLOWprNi11q0zREeeWAb4J
a9m/rKfmtCLDv3uGTH45YLkgf5NBbP+c2umNz6Y4H0oBiOKFieskiDF/OYaLV4DK
PvTb9OzDkqmA7MOJ6rZ4BiiFVJzZNX9f144a1WXdN2bpkjpmL40FPjSEvpAXIeNR
HsMmAV5zw+3h3SAhYMhujprLboggf0qkm92v76O++8/jwj8u4APotK3zKNGw4K0q
/8eVfg4DttxnWcMyH6zqDag9abCQaRd2MMoDQ3bfLIhRm6nR4Q4u4MA12AxqlHp8
dDfVuyN0Mp9MAL7t465nyjCS7ACDKec2Oo2eM0666lw76GowNuUAsS2AvJTf3U9Y
CAnOicAnDQYmObutejXTWiiXkrPZgrQrCQBlIXVbRhuhfvWFKYzNx3ZmdzqMrOh7
2cpQTuFBMqjKgJjZygZlVtbusoPT9GooJp1SsZgzsEYH/DYdDfMJlNAHjNRN7kxz
Azl4q7t2iFsy5d3zu2ergOk9eUzxaLGKAowZQqPtw6AbLWMLt2cppTq7wihnNWcc
pJb2JcNJjZkFAgHUgehhcknyiZzPdDADuVWx3XIUduS9AhJvwCx8XtK90hBenCvH
nu6iSwFmAk97UMxVMT6ulNXIv6FloKqhjf2zOQ2wN6pBstTKk/SgleBox5cf0BYC
/y0VY7Ml7ZN/ttxw4qgw59M/SU71WBmSJJYOWs6gb+aLSJm4j5tY98gJxp0AYiW5
PvhvWsTGMhOtXtXI7td1Ye6AqSZlk+a7/MAefSZcbKMd8Kl07CcaYKfnUz0QaFzZ
2lcXAQe5xocAHvNxYic9ve8kfdCr4zx7hf7mSSwdZ0DVExjuuLEnoSICCV45OHJB
rW0sE+46bnqciUKF+K2HYWNieVMkaXShEOBqH3j+vM14PR3Pgzv5xN+eYZtczrwR
GpfUtzDtiK8mq6XSsc9vLgS3aXmDenlIsx1GBAju8/FSTMlcfDepOv55o/OSziXC
5onMbaau2UTq+UmlyfqHqEltNUUypEJi9RX0u5VORCrQJUoAILBc0hIXIcai3dvn
Ij0GtNkBWEGULQkZScRlSNj8IZQyR2Fzn3p4T9j+dr+5bP+P2NGGDxs14nONSNr7
f6uwu+dDcSOOPim3xngmU7fRSdCfXeKCXQ/GOqzRl8drK018+lSg713DrRcb+8D3
4nr6BpHVeug7NDxB9Xwl0bvRwvd6/BJuQkMG4eZa71gRGhsr68fbakIcn8ttH+xh
Mu1m0m1ZmSou523rbpT4OhGwWd68bJaX7dG9uXKRl8Qgg9+LCF00WwcepVYdzk1e
xvbbXKU4mQg8AI+RwfXbRN7juaVJ79rY/DUlySu8mVjQFm9goZcjBgmcnmIv1Q1Y
58LjDtaQMLLq4Ie5s/sLiY12bkofUFshEXBzjEnb8GmUNpcdaXn4Ls4TvSy6I9Hh
yxye5JSjeNh3coYZ7ioknpA2sKpVQhydY+WkFmyOn3M7Gujf3nkBoLwQs4Of5xNy
gNeE5daoHlj7d5ZfiprD0EU1hPTUmLKMmWRjUNMJDsVfU+aYcwUa9+Buy3AGmAZE
qN0LYQ+xbpfXbISS9zQltSymoyoKf6WUEyMfzgGaTkmk9CcUmJBgZl+Ek2xhafXc
IhrGMVRfUgJ+Ms3zD7i+LgkU3rGKgXX5ArpcDdxnfSSXqYzMSOlx87qiD86JYbRb
HCUALkhpG8NzveJlCSELGsMcMBkmhK6W5/ANLEaSDHJB/tQV5eqzVMKCKiqU48/4
t9Gz1qtCvap1zruNbJE5iqfUxtAeib7xv4wek2jjnLTkYordkMEM2KQiqtLVDpwO
Yp3Gx3oaJIcCkkhNZxDna3uBLyg8D3+DZfAeluYwfa+Kihh/x83Gv5Yh1fyGbX9q
H3h1vA7i3uFkHsZ7sEILXLAr4fqPbOr+nxcgOolRJs/LQgh11DQ7fxORFk8x1eS+
wFNWxErRC6xd93yOA7Pzk6+KXajoZihverO2dqHpqlh1VN/CAr0bt1rlE6dJ62Lf
4tt48L70zMMTNihxPmSYKa1JrBROOdDBl5O6EAl6upEJSnxTYKdv+x+wtqDjrjwz
QVolyjaADuKl59dCKRnVnYPgd/GdI1XF0W7ADdSKdVqMKE4MfC4kAuYYuIxMswNF
2siU4gZEHQ820ZNvqNbxo4McI3lyFCl0oNx+29DNkQ4WudXpo4CKeKHsgMfUlCWp
zUiPyn8k1hTWd2QUGDYwV7uSXk31/SrUpeEbwLhHtTxOg/5zB1qSbKd9l2UTa4YT
jOViDJjN1bko2q9g0tXbbfTCilBFWv+StsorbqNzTBcLa15ZUA1QGIrQvLdIecHC
qYqkz40AEbevcebTJIUIm+mLExs5RdJSg/ig+lUcW3fXLjVk3WtXIsCFjI3Q2OqM
yNFcbBFD1u4L9aflODiSEMxdy/vtF5zCH97lhTAsEWl70WcAmgdK5x6+SpyMkEMg
sjOHjvm5P4CIlZfqLnnrc2heQd/pLRVv4702PZcdATY/yjzFw0vjQ3as5EduR0x8
CWbcsH0Ny6peNc22z/IWHincTLEMJNbRvCBm0vZPl3qZdeSryQc1N0VzokGtbvy6
WWi2TSFPKj61Q1FKXX8m6vaLoWC1r2WkVRuTz3Ul0lgwIDSoovFS2xTAfUuI+pha
O1zqeBGqQfMKOM/2/xes436FlKwzMXvLEy6YJ5N9wWadJxCVUMuWlP2VWvKk6frq
FpYR9C8xfUB0nGH3eyDUOKwozzQEZHjtxXke9b12a8zOi7RGsU6MlsTUKuXTQtPh
ZSddppr03ORF9/Uo6dkhrt7+6Vczhoq/ZGk3Hgy446n4BA3ZabT8VdPTzuHhhIze
weoMdFkSTVPasoTlp2d/TFGTWUw0zLHnaF19Tt7cl3/b3phvj8W6xEvIdAEFZXyd
iFLqmiQWlVfd1LpNR8vOt9H5YXvYVzj5uVY/TRgDBIvbVjZb6UB10bkyv5cGPBfB
eXibDvQKhS4u6jgZSyyysq6Xz/worbug+jlbYLecPfmxj2pJ0kyUILWh13NXrEZr
pwUHRIDckSxP4McikM/qLqxDf6Y0SMQ0yPrFub+QlzyP4H95ZDaib7soI+1c885s
7QBC/eLeNZZDUNbDrqZPA0zyt2J1xMM8mETEecIWu/WwXVWyVdRC6Ky+NkdzPCIi
Uh/oXSvveJADsxO/hqhzYV7RXLWF8fQP45tEl4f1Zmh5RecHDHNXSZ4gDbWkTI2z
UkFXERhCFAHGWi/afquO4LGcDSZgHX8YhrX/iu7KjGK00PltpOojLPJeFYSwq0CM
xA6YmwNVYtu5+3BpQYt5tubNYMjpNPUPmGRz5QR2kddO9ID2CFIZ+5duZGx4dEOK
8H89K8ihWFgm72ZzKCVr55kTrZdmrpHMlMRISVg8CGvG3PqaKBe3IvKohiKrCpKG
bLUAdM7ejs3F+3LUzOa6+sjDlvx8snLXgCE3MC1GbutHfcT0WLNhkVg7HoFI4j5e
/ZwrbD2K4Irazq7CMtnQjonL3PLx9TmrUYtF8lbU15r/IdGdlempIi6HAb9iWhQZ
znA9kZgIOaEvw0Pjw5fr+GvXJGLTVmP2vaW+YV65UhsMfWIwwMSf0JKofoEPyRQP
Epm3vAhX69s20yH45At9eLtdDSX/NyaE8GjmlYi+eWfp9AzARi5he56sPmy5uScO
tr3GYDrkPZvzAYtTQYvnhLd9jrqdxZmlA+99Am4us95K1a0D23wh+a66YajaKKRU
JDsbxl3WcNNcrN2AEImiSlusnrrurh02ZzOKeQtQbOMGbWVRjF8FZDl82Cj6KtR9
rODsRhmiz0cp6r4UF92Lhajc2HOqLjoG6OSyO+toBsPDB9Cnp7zZnO01RU0h7WQM
2f4uISTDZAUOdTeI5NTkpBB+qoBvK4ITbCZbOXXIgamZGeqGD+/YMxQVfHFF9OBE
MvLLvoqC0nb5gvsOAq6ZXmyOGc8KXONymh+bVEnjL8DXvTPw/HK8pV8JKQlrtoGb
L4WHsM6Do1C60u3KeKAaPW2Xb5rIbg/dSpfWPtgZ2ce1kIDwNlJGeOM0GP1+UqEP
LePNu25Rk4tXPaZri0wwctcCi5Az2gEC1jD3q+RTYzqOh2QZulx4E6xxhKMczXVz
oEeGGLTkQi6OeNtz0vhYoBpd40K2+DT3MJ3dH3c9SDyfAMHvIwFfVWkCOW4oqtj2
saRgjVLO9ABtngWPvsK4OkU+wUCEAxefPxlyD1p32rfezyyz5Ig+erBuS+eGfaqT
GOnSfvl+SP8vvDqd8RM168ydkZD286imToALaWL+zP9rLwAs82LJzUsKuY+cToSK
QF80gYZgiphkcQfhHK8nd+lC4146jCxCXEf+GYDIQA6JfJxUm80BF713V8MNztUQ
wn/ggrEeMGcAr6UphetJ/K5ASdtligQvI2J9iAjVUM0mDj31I9fPpcmlrPhscZwN
7LUWegHyzhpWNdWng7nfe5z28V0sRFYYi7ElK+bZVh+oUM8kEShfH3mcJZ7d9hnN
YgwIdy/ih/p60r/kyN6a+mbAfYSFlKP7//YxYngbkXYZx3Gr2ap0T2LfAeU379eX
JQCH51j3iSWoVLt/wtWMn1fVWRP5jxMrznqNHcakmmmS5CBVbTErl4ePc0mngBmv
XcYe+9BSppq26VsZfP4xlYJAh3Dc8WLEdtE21MXvRNWUVFZUpSo1WPvdQXFgpVxj
x8A9QGxHvubqUXTZuuxPMwsUP33WauGtnqV9wIfRX5dVyoVcH+L9ZtzirHoOAnvw
xHHysvqah9/nrg87At3sygCI6PW+t8aCjUSmo13v7f4ipTKmVYL0WaIe81t4Gf+D
DaxyMDA2o68niIHLWVxZto6YKHEz749KG45MYuvkvH5JF5h82NZ/pVG2u8sNebq7
PyZo4r0b9BsUTfWmWw1Ys7zlPKxtki9oLDC6MJqutn/2rXBEsJdxSDjv5sbzXq30
edIGUa8kab0hACWxwgxWp4SsOqO/TamTBZV0uEoHsIybc7HrVFH53TxsvHKRGYbJ
bGbx3bhajz5j7VwEw3NO3LOuxLiRUZWbOEr/oNNz01TqY/XqSafTRGL1G8YHb8xR
J9RD1I9qkt/ohjVddbQcWMJ+LmRS4JQls7qtpRSZZJCpZgAiBsyJBEp5cKiCd5yi
ZC7rVc6lR6UXRnPDzjzerkOCcyLAqZ6g5WYLFmo7XC+J/LXuYYVqQyHghjyWKdBz
5IIzCTuW78RTUYHVXbmA332LAHyeqPsO4Plgye4h4mYAph7ZSe9+uUtcJK6hC/wu
/Ji7FqcYs6q4JrxyyKwazPf30II3Z7Dl4heLLuZDLUJLW5J/+dzCGvhiEzP9u0Cb
gI2xR8yDlvnUmgILmdWFcNR5IE0YeZ7TZfMWnF9CNS2XNubLB85bsJZZ6XLXl2Go
3QpCxG3RUY3jU5CVbjqHCEmO20VrbRnogeZ5VGsFZTsy1dj6NB0swdA4rN3Xt8as
MWNuCw/GU6TER8Bs6yeK+gqEhrXstvGDtxpmrLJA2b3nxG9ANESOW/DrNT+ADZM3
KgqceS5d5SROhB7PSDZ46S9J7TN4277WNrluOi5faa/dO2Yx41xtv8XfGMDwBReI
tYtPjJbMsQNPEgFl/gbCR+7qT/J1N3J0ZCZDMln60ivpBrVg8dYIMH9lEkg8A37G
sHYEWlEEJhnn/fUrAidXKGWDY2Mgwwem0Ao/wzJW9l3LsTRWe33wn6Qki/dRGV/d
Zb/XBFoErTwMQFrjgE1TyGamKWWl9jUuBktxG5trib3U2sxwbdzQYo9eVtr2upuu
OkP4/1W5x16c8u19FbGJY/UlbEbl3TvOS+jwNAx9pqLmGkGU8OOrKHWasK2bnbxu
6FZbbNPZjvCamawNjUmojaV+jwLgONq92G/sQfrCmlNGF0V0uNNx8FPU9u3eYyfE
lFsJCwBHA10/AQSkzkL70BQisaUALG+pPOa42TZbp7TgaQIR+21lO3QTRvC7zRPN
dOAuUXPIV+klaXnAXQ/fo1c/nUspMOEtAcNdLCKt1mZ6kF34r1tgOB9VMNifIj74
B6S8Fkid3pXXQiHgPHSc3BA7GtHq0Cvj3nUDsv0nGRy72jUPyCurQ76GOWbDU0DP
iEqIaz9v74xpz+Ar/0s/7UO14BOVIR1SZaD0TMJ58rG+/1dErrKMkEx1LoG4sEYv
Zklcdf5i7OLtTm2x/N03wto2b2TWRnchcxIpTeJp8HwTVH6AqipXBsYF16X2mc9a
7FhSE0NvAt4VCQKB37rVKJwaV52qu6ZryY/ePI/5eWL0PNkiImIquG5bZiGcDeAT
6CAom7bsW7zlV0HWsqt1aWQJ68FULi1ToAleIPqNzq50rcUQ0Gsw9hrYY7f021iV
TyUjwD9EpG/0a85S1rxwOeurx6z7N+HhGh/tt5Toa+CSyKc2bCfjOTvsOwdsEpd6
U0XaaD5RiBGtMR89tN4f8OJENdoj7H0/RomVdUzvTDs7vQPmBrfOk50zYnXm8k2G
ItxUWZ7oiNyDbnRHrzpnnsPe20O5Uk3iUVqLCdwPGgA6admERC0Gx7W0c+8hh1S6
T6bIWwGWGePal4w68SFg2BiXn3Lpw9rtnMEvaLyNh4tzGVx9+btqzYjjXxcHM1+K
sA225IVcIZHy3o7PY/i9XgCJPXIH3RkqdvEbUUMYzylgKKDNpDdQjpfMhqeyR9cb
5snQC2aKvgMy5BpnzIAhf/sGzxsvnc2lLuQf858lpV6Sr9EIkJwA6KxkYRECCt/2
ZnXOF/ZTT3TNiK0coA5qKgGal7JyazCYvnm/VFlwr3BMh9lFdniPPIyGBVqoOm03
Q2htuPVS72ZGvcc91Wgcej+5MlhtLYIV1B7jQIiUvy2kb7mklvmq7F0UTqC9d01W
IKrUraQU7Lhet/SpOGGVlDSatqkBaVTP1jhUkEIteW1BZLeM1cJWUTzQuBW5CiBY
Zu97meNX2W0KcUVKdwr0s2fQAkJY+iNOqKDFbNIL2yYlCnxunWncidaGHLXKAm2Q
MzQkB3fInnfGfPFhGAdGfPdCm8jYS1HyOL+iRb+gijubKbSy/5uCkZVnSb36C/sP
Ty+LNy0PGGzLJuGyf3tef73MfTyFfZ1nIvQ8qRsiaQT5TLAclPN4w6Fx+HXxRD2d
arh7MEEij6GYdts4k3JyQhr0YnEXDwlTD/E0kRNbqZG5MHKHYVbDpq75hpnWfwZj
0cp76SfKy0e5gHcHn3hrUl8x3BWKkGaOKETDwWZMvXqo39+qIoyqanJk6tV2dEkH
gTPmePo7z+h8pLgOeFNYIu/DsaaLK2eFPvmlA15HltkJFMvnKl/vqmzUIsr59AjH
1dpXBx4nD+32v8kmAGrteVS4H1vIhJWMnXuV8NCxgzCEcjrbbLFG78iS8uxclHNb
H8VrRC4ruw6BFI0OOlJMJDr/Z+bEgVrH/hUhW4BYWQfkeMwvh+jE6WTDa0vctNfA
C8EZ56n4G2wvnvt+Z+qB2o+KaHK60+XxSgydDUkqq8jnfuWrNEejt/cYU38DzjEN
PI0Rn1pQbhiTF37kBoyyhLNbM5Q2/wY05hD7rLwfG1ctkRTVV2aXWdEkPl+I6Lsg
1y9+IPHHzvwCyURVnohOsFow6sgZW4cOYz2QGLohWa3Ee0mqHLXn7NM29tsNcE1+
XKQAK87HfrXtLKyFAmeOyz5zxpDLFDQk/yvanhutZtXtf/k/lWYdmtDwezmDvkh6
YxqpntQyV5NR10TuyhpSm2/V5NbTEZtwuBqj1pi3nB1sRyuF80LUJGAesdRUIwGy
+PYnSz/9jA9JbfNYvBF1b3CYp4AcOdsd8l0BmchoG3qlEWM58WS2ZWWFHWC7gaOg
z70LtMC2lu5StsrLhiiTtRftQj75aj3Upohi5rl5kmcRPVPOinIOLLU5Up4EsYzi
vow32aEe7Z5J9t6Izz9PpZ7Qmvjqapm2vVH+Oi4bWr/mL2CdZTfjwvbixKE8v08z
sFaKuQhax3SNmhNZGdMfoT+HGofHTHlZ3eMglmto42JOuo9Xesz9WXEfoen1uSYC
XfODYsuCzrXz2TZreFvFiHy2dhk3vBfXkBlUwOAjLPsdCwNXX3ParHug2YMKlK5Y
3Cz+0bMnxB+yrjkE/xw6lYc/pXt2JF46xHyofojpnAHfFSKkVJ4EcerYI5GJ2ltE
Nt63qY90ljFoggy8pBznW67MhXijGnYId1oW6s29Q/g2Bv2Txux8q48Bj4qTK3bA
yoeqiAePUcctmgUAmYgWaCLCl5bfgSStZlvZ+aII0HqEu7iSrXCMwV1jJ1CWeCmk
jSvNc+PbpGqhUOtMRL7JVm1pT18lFS6/ONPBN+n7BJ2OkqH7nvQPQw42ho9dUKc2
87yz+GE67frosAtXIQDFHjFkHtsDBiN1ThPAti2o+keSz8VOUuFLa2OtNTuibcW8
EcrnCyMLHKDS8P10rNjLmFoJ1qYJgOxJ43wKI1TuAT5MotJcGBPbp1hsDpxMbxe0
f3L0B3B6JnttoYTWdecG90rm4NEmH4ocsgs9Yzsr3ew76bvi84diW3zJ7L2+AYT7
kTTV362sKJugk9t3uLbFiprHNhBVoUzuXybZpuSqDs0Ox8tHknINz6seozzVHb6H
/0ZFG/27u8G0LDtJ0B1M6MiNMv1r9YRxdlb7i4+ed+KgedtIg6V05bk4JP1XNt+3
CzMjK67qb+uyq2nj6jAoxlTkj2Iowdzn7NZp7AOGHrt6kg+UezNyK9bcRG7GjJ9z
38Sn2Qf0CMVAtwCkqoAvGhL4aJDBFtq9GOca/BiIsi15nMJpsC/9Rc7L2sL8DXt4
cWyi35zofujovPOPkCdfNnfzhXkWJzklPapmfq3uLQOT9ACZDNbXN44WfC66vpSp
CNbbUoF04AS25kx5PLPm8Z66J/ic/NHDqQ6V9pX0w5M8AnE1kbqzzBqKmr8HrZP8
O617tDAq8PT41/FzNiYN1+DQ+VkG1Y9/F7TMR6Sn+yIZx1DUccIoBzvIT+kfNxKi
4LsR9AV/J6ykxYaaehibvUkBdCg3ymnPxA4odYx/xeEvtIc12VStGPI2S4vwgGRy
m5OmUIOB1As742JsQtqIh24gcshTQPYQQtXtT7A/GR8t1sLaCeJ6Beq4SI0fzJDh
qImjkgrtBsDl8Ke7niB622/C3g+ySC1rsBXZZP8SF3/aEcWlMDKg3EIe2fJ1Wsjz
BXli+HusC/2uWv90urhzjb2RuQfsDWZKicrWRHL13P/WOaJID51QORp4+NiyyvXE
CnO2lehoEpaO0cL1wnRRNJFyDX9sZ2TvnYhHT3EW+b4MK4sG214FazqAZOuy2SE0
sL9AotSV9tfPPz95+Z/x57zE7eJFCIJWAQmcQHZ52vdHdxEcine/vSNzyYE8hZRF
FTODw/ZnWkhuSFxm5bi69j0zsCpMPoTUzIJRRCsmFD0b4GFUJrRfWOON+pbJTc0i
OHTT6nskC5vNKJ5TUg2wQAQcFQk8i7b3FyGYMy+2n+x3x0tl0Kf2ID/IuQg2AkXz
xPDFZg8DmR0j07r2UFfRSt1Uy2+iSWzOgbzGd04l3jwdGjQJ/epW4dJFLkztFQBf
EziG8hzX0bq/L/3Xl0JcfF3nlMPUUqywzTve2wjF9NpXklESR/QYJ0nrdz3zmkzz
yIfbFlXCNCN0IjE7s1NOvQvQPTrqDrygK1hyb4dSx0cKBlQHv7I0WZJ+HhxLo+CD
hMHTGohWy8HfMhJgQcxaqJ3k2GDPYz3O+fi7Wvajcvtys4X5Lin+Tcxm2DSBzLPL
/sZeaZWB8XXpyZ4lwGsdOlsaqdjP5fTYKYqf63xrI54jLdaZPP2Uj94zhDv39CnP
ArkwcZxfzkdDz+nNvYSp093kxVoPRuWPYWiZa0TEYACOEBeD1gEwS0kx6kg+/bwZ
80hVVtFcoeOqPG1iUYJMQXS/wmRSsQHlfIchWTeTqo1cfPz29mEsQwLRwKh2+Jvw
FOq2x/WyqvIFHg4B7MGkpyfj+NnUfb2Pa9yheFNFUnxYR8OOvyDN1OCNb/widfK5
jouvKgqesEGRy4OozXp6Zc2M5YNbQ9UPmJyDjhBcTPsh8wxA1OW+gExfQICu0K4E
epyccTfewmMAOxMug+WqyGH2fPstZr44bSsxFmKUlAgOLs/KSBPy6wH3v1uR8Z9p
HtI9pN4Fq9+okx18kAAWFvcRn7LQzNxvI3zcRMrqoxSogHw98bMN6wWkn1jySQbv
LaZKva4EaTFv0A7Mi7UYlHHB0ZOts3Fh8m5u80JZVMV2107rMaS29xpwbltgWpFj
O1M3NmJ0TwSDOMoeW1CyZIz1+vJXgVJRpLjCV/VFpFSYvWFO1ArEmP6Ts68Yr6Gh
9ay2UOA8bIrfTnKLBf5+vLxZ8TS2hsc/A0nmMVX6zN9fIc8QZIzp12hxXMOR+gJK
oo9bxM7cRK9cqufb3Pl+MrBMUuYd42QulxH9ul94qWPlAdaRarEzqV5GscwvSf2n
oh91j54VFWLLnHF0/D7Es8uh4vW9dkfjPoeEn/wYNqqork5A3S40nES6f4QyDsJK
uZW4sJXKLNW22oBFgWmbFSUd/8tITS7b9cvvkoEDvUWsvWRqEQYlm9XZ2MG6U/O7
OPYucpSrnpAxK+9d2ToWrh2XYPy2ICF6a/LZk26ioEa9Lwd1JBPLLA7jZMVYp49I
wjoXf+NZTKApYyNsD+F1Ith3nlytetX9SeBVCw74ILCu3YYeRNDIUXoDUnXbnnlX
lvH1XdLtVp+AuV7QERu0l9Pjn03/6uqek28BSaJrZy1FQkfPwZCr4dhIfY5sai2D
mQxdtO8S4c/MxztwAAmDdN9eLntrMmDL4MPL9j3NfhwJGbUCV3VdJ6deGuPr+vCF
TkrtW3Bdhb0dBU0Jh4jpLTd6sle2AsN0bRT+oRKA1P46eHDn/OuRC6j+4Q1enfOG
1kCnTN6zHWZy84aoxnVNowPTacLaOlxbH5awXVGirN0GEtIfXT11QTkVkajKpI8G
noDqfhVHPiBRvjBl9scw5t2RBtOYfS+kWFa8KHuwK3VFSLUMV+ZpKJ1woMQAoMio
kUghuytSZi0lSO9a2WrC+OjSDIcjtBogHaIc4os2Gvt9S4kp7+KqqJV9vXwOETGG
3K4c+q/aeWkpsgfbEqg4Y6ldZ58kWo8WpVuueznIpuul9PqVxDb69KKHJ7g18fZ6
mXpxQqiyPQdMqV9FtaS/Moi3BfLjGJzQ90JXjwHUhghPQj8kcOvoqWVdgFXU8UJL
5mxruxjufWko4xnoC4xV2jwitucp2ZK94c7F2yY8s1raCsbAjlTxyWT98DrbiU9Q
3rG/zp79VcxcQYiAWb3iBD+LF2UfCNFz/v0Gw/oX1YRXrB76UJnlTM9qwK7M4Ody
ysPYtIhQ9AlafOkiTPCn6Ms/HETZY6jZe4aQ30wEnI4dsCX9RrLJq9xbDaFSZYGi
ZxITears2aLjq02H4NL4fqGLVN19VM94bYVN2hj64SqxOhXGj6CNITLeDlOzaXrf
IBo5vu7J7mOelk1XWTjsOKMwciyE+kEJLLdkHuuAsUCzBjiGkVfEya9raGTbKqEb
qyolprXtWl+/C+wRGyYs2C2ZGaUUbCa2o/BTSkhqBUegkyDCpqHNqWH2cUNaZajB
YD1kxdXTo+NMHBz5Vh1K+fiKTPpVBZytOGhMYmcib9t/wHQTUNAa0DNQlPD7jz+N
sruaiH1s0zF2txHbQ24fZUSPC1h0/+ZsHtk/acL2quMVJYVxEht5om0cGPqlZmkV
DsLaErY4d3EbGF1NNhd8ev09eSUTx3n5ADU/LF7uG4lvdPbq2aZMSxZLAHNox3FN
m0BDxWa0As0SO9MdQOgeLUCBK/rL37VRAtIr2zxYnw1IJx2+wx3x6De/W3ciB5i0
+I58dUxnSW6dpqqsSCIqpHiHZ6myl7eQT8rrQCAkOjOUeelCutp+caK7WZqtWlxD
4toSRmP6u5Ts5Ol6Nh6+PzsKu9x7tVSahHbr299C7Q4cTCguetkqliu+Gs+63jB1
3m8PRmLiea0co9UED/qU5j4fJH6gnEXcPt4EeZvoPeyy09fe4/liFFyd6GbpBEij
cCJQ4q8A9gsdN8qHeiKu/oBP4Ns+lHEE/l41AvBRfNnudZgiIyZu85IafBqC0vE8
DtmYt4zPFXggrNXxUIRaNG4TxkIfW3gXfOxoTXggDVdJLb2sPYeAs8Co1BSbgKnk
CzL6XxchAm1+SnQW7cY71pdEKpC/5QsXlMUB+K7RLZnUaIKyK2NgQu6CpNpYQ8cb
AhOLnMi15lnCX4yPB7CmlSo51/cXlM6sjdWxMOSZokvQNF4FMyyucMwi5+5yE7JB
YUoISof69iwHL8XsAT4ql7Ve6iIcx2LZsZwwUNZ9uGSRSO634c6NdxaaDMcuXmov
+To9YgMugDTqoIYD7Ywx96zNozY2BP/vfVb1ljIITgmZgdmjGwki5n4gi6PuXM0j
3xXnw5Hk92RgIs27Gtrn2feSPeIPfAj3Q62eV51xbrusZQ6kqxAf6QKsbvd+NGYV
DCIDMBq8r4her3aIm4Dy1shPro5FFNLCR9mAs0lcCdkpxYIeYS1n6xAA3Kz1ffR/
JUC7kHGFCG7hKsUoeH2jeoo9cJbQm6ae+oBNxvg6vMGgDK+PQk0u8seT26vlHvMo
H8khfnO4CMvnGqL9T2VyvywiFNVCnwEumQEdOrCfPT7BMgV/SfIgpvhfJUsNsDNy
MrQIwbO5v6vBHMHiwlz/IyyCw1I//eJ6hivKyeUIJW9vChXYlaMGm1wFhVjHzjq7
gl9ZHc0J3mmSLG/8B0HfTlAKG9+U8sC/OC23/jxyKRWayWrSHLUvZjeHaMKeYVeS
fDmQbH4tWChQKzUuIKzYNTkMsl4mSjeHtapfhxOEl/ZKBJTsYbNXjfqg6Z+l8tID
/xY042ZY6Q19s2cMN0Ca884DYsnOvi3fWbBR/8WW3XaIdO/byBtDg+vmF8ZXx8Rt
VkWjQ/LMwZgOhx9sY9bVpN07h3Pl3IiwlMYnmzhXdE96Y6IP0iVi9p1V9wzy8n2x
K8zHe8Yy1Xy4712Dbd0yoICcGq14DR/IYditUrghdbxUAkw1gzcT720W5yGDgGlk
dmcop3hfGWA66ZwVvBeSZB+QIaAAc6J1qmokeo8Z7NXrepDDwNDQ8jrzXWPQlM+G
oev2X9CFagm2/ICs7oA7idWsIFSrUMmmJTKUtPN66XfhiZfwMbtfIyFi2fVTjyKg
tXWorfotXihJLUVBBGKDLArrQ20LQfVYJmhIWqA7HKEB0lgGXECZkYDN56a4YqUx
8OqWxL0wlxPEh2jOcK40JrvvIORrAd0oNbtiwVu4wdfceMbaRPglfzUnTrRAGrpv
bY88Mnatq+sMQgxGX+o7Mjl37YARpEUOmorJaW8jwTfefVhXqlR9DnyLezWBjR6w
9usB11JjdlZo17AfvFOI4R3Z1e+A8PWbH/b0QQ/yyd0dP0ULPnBDa7ffWdJYXhm6
g3dHjpe+lcWvP5eG3MV4eWTTkxpedw/6k32ATRUuGaM1qWMye1NT2ptjn0b88D3z
KK8MwfF3F2EbZfuWhHEoxyI9cLkS48yAPNj5hapMvczjoEe7tlNgS1j2ySgcH1r7
reaEMDVmMvCoFOfUjLcteYEvj5HgTgVOmom2huKBuYyhFKXDR/tZGRoaazBU23Sj
dbxAwXoTSKi8LePU0wMZpgwhP8Rq7APukRzPrXq4L+k+pki5ZOctpSVF3cal0b41
Tt/7kWoCjfCts8F90sw+fDQVSAZifYQWOPmSG9hJgwc8rrKa0202qj1MimOuYot8
Xf9CD2Hq9t8ArRVwqp0yOc28sUDKZqESUWlfV/80685nO36ONvdS7OrL8RzlDRn8
W35eo/CzspCQeUZVn9izDNA1rj+JfeWkl8+YJ3ZoxnkhxmA/3bSvrIwlUsvqdVuG
ihW9eV5rc0ciOIJqXyFJFQP76wYr4m4vHqJlU0WxHE/vHvEQTZtjemz7ApUvnY7k
2AIR/jk2g1X8TVDWY35eTcFORUNd/Eo1eCYlv5Euq//4O53PPlg/qwovRdaibB54
19boww8qGVnk/qkztHnM6JXvBAuvf1YUJco+EeTONm78S+UFb/VH8vDo+kjPWcpm
5D+A981sfcpdwhjdMndzZcagrnhq976xVGiaM1d8IZ/vQsE90IrPxzJ6SSvH/xyj
91rsdNmfe0DvrvRXwWiuNsxNre8EoUUKbjfETJ3X8GrPEctC6XBtbPjIhl4anuIC
CUDIGqhxWe3PZ70GqUJBLU9J3ylaj1FMNGF8iucNa+A2zplz8Hy5M5qiVVK0EKiC
k0CBN8wLs3qaQdcXWCvwWYZTX4BNcpvmP70GyFcvw/u9kF+z7Rxg/HI56fxIJPMa
Zjkno90BLoCzNK623sqO/7trs2tAjkqkyN5New0sISTfIEt+z2lpy0ZEZjBHVmXd
WIB2X4CR7ZLwnhK6WLg/KIO6Jj6IJBVNZhbpRjrzB2zKFtXqFp/RwbOwoKb71cLQ
2rQU9o2KbXals+lvmQRx97nuSvPjljRzLdoavMrvhU7s7koWQITC6wvqMKXpbOBi
DtA6/kHCtx2y+thTazBJ2FbWylvMuWqnumMON4l8u8jUCgImvkxHhK82TiuNVidL
QWqJE2YjzXgoExMA+oO5kxNsYDwkK6MXXz00HbNF+Hvpa+3MooAgubQU01qPHubp
H7gWYSGroBj1+r8qLeuXgieModswYiGBrb2ryYjk9Tliw8+J3cL9rtnY01sLHB/K
cAjvatkUeXGT1udZ7O2F1IBt54al+Iv9uGdvTyaBiFCMYV1IPqFvnL67h90+AyeF
PmV/6gLiPnR2nkDBIvmGKp8vOmBKW9+3jGghYrTH2iHUIuEuGM9J4RiWPWa4yjav
cgLqXCaphzutn1Ala0WtIUbodzRdOU16qmch69vrw8m1h6nSwEjh+u3mm3mkCA0m
W3Zt9YshdPwMYyD2kGJB0CiHHs0L32x/rrrhpJbHUOtgWoW+Cc/WoKyzO+g6uQZg
m23RkIdvU0ekdAa1J0QupCAZhmNYyIJJNr2+yPM73mtDrJu5g09wvnMVN+Txe2yL
lMTw3APTqreDMXZtWYmw8NC35M09axdezj0iE993e1fdlGSAfQkmOTb8Lv3xY76h
HEl3wYLxmk+UDCiH1eEXVhG7bz5haEUz2FiUMXdcETt4QPnmFQiLDlOH/ba89n8T
tG5ilOjBFYjriz5rIn6Cuho+i4y41MQ/iXfReR2VojEwiu2czqRMkk3T+Nfnhlwg
yUu8OCnpHgeqJZRhTiHFmHUDkjVQ+n4EuH5Aa4m3FPb1sb7gttQaPhu/xpAfbSk6
wvwb19G6QLujEXUqrpwdkqDslc2LcI1RnbvTQ7HTw6SV7UFVqaQCGl21c7/VPMyO
kYqQ+8wtDD6+V9cSLACvsqgWbuy/JB+dJM0qreD/eO7qp6uszo2UazkNyRHwquuE
a3gaK76Chu/ASRzbvgvDjzunf9C+L1dowhSQOFB3U3ZmIDay+7Vonc8QTU8YOAG2
2mkBDg8IwOkBc2c0aG0Eps7Sy4I7CE+3+rZjrMnxf8zwH0DLgHsOZ1GWODmgsyxL
crwFbCo8PCuUOOeKZzk3cAriQyIDDBUX1vS1VXnp4SoU63vBkyGaxDhxhdznir2J
NsP10zJBjNakwx4v21YSMozb46/tXp3pMOnAkg7dV1JTcS4E/vIAB68zavsB7cSk
FIiMW+0IQxSQfqqEMo6bRXHUDp2spg/wIDFjYcv4kmcFdho8pBDUL8y0gkvLwhwv
/xhuBivDFE693EnWhWgDNWndrykNNFCil7dkn2V2cp9MbRdqOZvoL6r+FLUGTUSa
DVAZHoL6+WI8PirSm/7o3fcM16DYqXpj9K0ASf90kkj0tYxkAm+kkRsleWAXWza9
fHduXqolI7IzL3narCwCl8wvaJnCJUv+4Mo02NP2QJ/vwsFLJP86eMJzoh5GCWKn
l2QjZhCoXCKeKsyyo28Y1KVvG3fOtugPItKtPt7EHRlotPeQe3tMiSmuuH94dzRm
G5jQKZXVJt1VxR1kINTMPlveeVSXml7INoizvaxS6Tl3POdEVz/Uk/mHSWEVrvfJ
fdwL7YzdQMe53JvPNaKcNqbk3oUXrZisCPPoUUODFXXO3yQ6jEb5xOTITOD1pLEQ
yzXrkSxO6uxU9fR4xsQoBuX4Md40Cc90lgExwpZ5/lGDDOyZseYJ/t1Mbi3sokwG
XRWasCciDkzXh2vh8tVOIC+6+4H85eDaFbo3DJgo9/tZ4AsrosQh1yPPkk89qI4y
PxiQqNAi6dPm2cZeDg/S1nUjMOss/Q1f2Eo2O1Hc4QUEKmcBVanHG3gNsrLBBy7v
SfUfynSd31xUx+FH6Gak2MbQJrQVC5qvqYgjwKGmdchrnGD9Z2g0Q55pBp3WsClp
J7IhyNuECRt7+zXHPCRfQWqgWDzVqykvXXa+yfxWaAxci48Qie+5c3fBefMu4/9K
vd1NhuEObI66dU/Zeq783knNJ20Glf+6HM6HjE4q2yUwweY399V8+oaP6Q2ubFvw
5HpeXgJSFEs5LRTVBvmV0c5ViBB69YuxC6u0Sx2IraA4wO1xmYq3Y5SIWnuwYO9s
KZN2d9jzleGsnhU+0Od0j4awUrwHMraIOpUbtPflYN8zec+1/voXiOzqXKXpVpDo
AIMMJXFLi2/2AlJKEIvB2djXMRZAFKDbVuKy7bzEoixJRa/XPrE+64A9f7ZrnntJ
UpbM/71wlcyclP4ynHbmBQ1tnFwfENPJ5lzRwJxY7o1JctxBQLXX86mLAivm0eAm
nANo0tsJk7o+a0oCQWT7H3QiIjGmlxCVVSNbcruYqmS2rsrRJhdL2RX+pbzbKgzt
RlEPUO5oErBH8m5WsKnSmehWtrdEeSutYvJVn9iivIP8XIC5t5GOHUWTIkpdJvqI
6q2yApgINwFfq4QEn5ov1LgH5SCf+22YANaD8OWjk90Q4t5R0whcGhlbOw/bIFYC
eipnC0uV89KD7F22Zu0UdVFMCIzw+e23jV3Wvusz5gB2LSQViQ1RytzBp5FZ3EwT
ioyGgCSQK+YsJ0hZ+nijIzqwnhriHaBDlJx4j0cn/6WqYTmeflMod27vbkkOS6Sp
5E9n1n6BneGT8xRt2hKIiXNosb9jnmbQNl+RPaG7l6mqxTOw1pJDrIIDXmOwVLNz
kW4EH+dwt5viIJQw9C9QxSITzHFpwrU4coDfGO2V0M3n41+l3/QyXOeVAuvqy1di
L5hjtPvVOI8uoAiStQRQoJSocNua4BZ/WtGmbEDJlUEmwl3Cxhb3fG6cOqtoMxL9
RyTfdkLN0TRKeZsUJAC7k1UZVQlf6UFOhF9S51kqRqZnqhhIiouDj3lMTMRxogjh
G3ZMA+MDELyqIFcO+DjP3ZNb8k5jCAl7W4IU6DBDQmKwEpYPIrid2cOmqCL6f83Q
O3nkdvwpEFVtiq+RhRWWK1qJHAiE+7/pl8UYEBO9B5zqliF8zEb4W9poswwAlrIe
CX2eT9MnCQmH22qdfJiW8gTW+vxq/t3cS949A5U8YWmrJborFacJ+hSGuG0LBYtf
tYj7IxKtxcQedsZNv/xUYgz9gLHPcE6n2/r3rkG9+HiiYbY4T0BBjA/oavF3Mgca
H6xZqtv0yfo/3QJvHgBjW7vlL4Lgf4+Xa3RaWcet9rsZGskO3QMO2WOUD79N8Up8
5BUmY9M5y5EybgnuntW+PBTcncnBMREa5ZKVtaBfk0WBZJhjIFRC0yTq3OXGvOkw
PRoWTu5xNFpV3ksWl9yvCoU/FuhkiIrVwgbrfcImi3hQGhiK76ql61TjC7ie6E9Y
kMQeeS+lmGZsUG8fpGKKa0u1Fku5hnRosCotjHL8MfyvWvpDdN9wYAM+6z/ja8u1
GPbm4P/7VhuZ+o3zEGCl953XPJAIbmx5LjEnn1RCTpuxAj3LT03Q1b/9TE2y2k4U
EdayNnU24TkdlID2NyJDdBx4x55dPVbFUvuwecIboZMq25XSALb0qE2R2m8PdvtG
ZAP/Dpud/IEx/qZLv8tNcOw2L9gVLDqblEbg+BhgpOy8pklaDtZ0Zm/pbYSbiwKK
ZDZeriLjMVGK5plQNLGl2/S44I2CL+M8yNEYZO2mckUUvpAulDR4AYTs9rF/ep7t
9fRwVnXZuU0hpcSWutvKvpIiQ1qM/fr6oRgXv3UoWW2Ep4H6J6d2FtCMnSfo3D3w
jStXzbOQXz66i9ZQ5SKOn/qKIX9COkZ21z9juABrBzE9v4tgl8Ue8CyE1KF4TrRI
sj9t0GQD5ZPweKZo66tbO/2d+JBYcv7Ut//+LZKXbroCGzb71P9EEINS/2rGDNsU
ugBkZSk5v0Qxt0THiBHMh6X0nqFmAui+iCdJ/47oebpQuv7bMeUNsSlkXZSyyXp7
9tXPojH2KwfMY0H+C/7Kz1oWNRKcesRx9GDLW7GMe3c0fwmY2BpltgiXhm/CfHwA
7PdYBn/LlCJmc2fSt0SouS4lOZKISb7VVJCZZ87s1q1BLRwE4nUv1nyL59Dc1zcJ
vpgdnWF8eeLqbrva5YC2g2NCEw+ZPau4Q6iVPF34xuOJVSi1L0WZQE5+8bxe+QQF
16oXQyqhZDPQi02MRGxLQh20MFckLkg3KpVezLif5Cs18mWauFxx9Knmfuel1cBX
dOclj3rP7Kf9ySf3lH7Jv/uN53EgJ3X+EbIbeBE9IqlG1dqlteE3WoiziVkllNxF
oGdd7oRnh1kPX44+T8kvxeOm35meqyJqWGgnlvJKZWhDqNK8h+l739rGBQBzYOv3
6u49RDzrv2dMkwH0yc9awbkln+l9FbbvLIZLXagcr4WkJVqdbOwWEbbMTIIK/3DF
e8meR7J7nhWYbXEZ1RY/ORYVK0jpWHcD11NgDIVts5RV36hRFbOsFT+uOgwegLOZ
/Jxk6ku0ZGkasVHAAgEBDvjQcdroAIfy5CTkmCoYOL32NpVPObRjyGSDwKd7IUn4
HNL29Nvx82dC9zhsShKT2LNU76PJGW/SQbeT8ru04deFTslp9TwfFHxBtX1++mhO
V0TtRQdEXDi6IkeGFC/CqYDQlm5JzS4FjYMWUpXIuBLRRBMeAloVeBr4NmJuE7i0
+aZ7QJm+nbn00TkpSpT6x+LOY3ENCfeCAhEA5IlsTTAIkCLlPXB/v6B65yxXmaoq
bJhl3fJzqufDx653P9LfsOUzq7PLDsojNKFb1J/vZlqPb9wipKQ6Lm3vrCXJP5Wc
HHlyBH418QEg9eLolbtfcc5AdgFDOy+V3AdR9IdhuTsHo5zkUVt8LT2q6+3gatNl
60YXH5rNDRUye6xkvdE3MtJFWUHbi/cxx9ViQORjW+IFEMwSaDS2L3ypw0txA+rq
3uTj6pBIyEIuKlUn8joBt1BTFye42SpBwRV3meARZ5qMt6mtb7U62SZsW0fQUu0t
N8wY0mNAWOek+uFsS1+vWmHMohaYBrAq+Kx9GLHtlfrXr5i+imGvgTco6WgmUEOA
pxi1xO1iMNJjS/V3v+y+EOVv3gns6teNx1CijHelO5FPahtw4trqk8M9p+daXhRo
hOphUXjUyq6V+mgoJmmVUUGmcn7yvQKcKAihDyyJiJTBzc5LxDAtbK1Kno3qNG+C
A7WwA82IDE7uqUjBejcmwibyUVUGlB3tzyTiJ+a5Mr0t16yR4ocF6m0xGg9fnKWD
1zKkhgTP6ME5G1xVX2Z2gcbPR8hwLBEle+V888k07YRi5jxYeJmQtgeUppapIKWx
1gqT4I+fuELSq8RapFEuYrI2Nj+s1v9q/gVgBPqkCpY6Q3OrjDgKN88PX/0itvei
Jct/GIjOXUivYLajAcFJpeF4zXq8mgGj5f8kpB+SjLzJn2p8evhmM1ALWM/eRm/o
1eMzGSSi3aqLOoXLHKfizkoFzLsIyfC4i2Pva0Gr6Zc1dSS8B+/Z+LG45Pf9FhWy
Q+pEd7aMgT8uI1ZWukrNYdaYTqkSKuPpGBIKL78oPJp/uDNpwX/bqMTt87kWSxGC
wjAC5eqjQrpiZ+1/wJZDZ6Iq+YC69OKiUqZeRgslPs+cw0JQYw7mt5iXXE69yPmf
AgjUYvwwCBz6ogfmwnNhDn/MqgO5V2Y3Z2+O7UzJT56XqPV1QLn9/U5P1ipE42e5
OKh6LV/qtVytqitSVEB+mBggZVI6R8oxnNXd5/46Fnb4+l+5cGF27YsrLpmgcXBx
wLDNytNnKmP5c54Jlwux6SZ/XOSO2j7n9doVdQXA2FrRFA/vbhqfF71BuBKGlPhO
0Icq6uBw6KZ9JmfQn0t8KU2FZVb9mTvLRxfQ3fMp3jhUljcE/2oxT2il7wJanpaT
OfCu2xIV1zlkiLsAiUAvdEXzpHXGeE0tAUeB/2GcDiq4jS7+AFn7nsaXk3IU9meM
1yd3YIhXahvPfbLqxGTrwREFOTJix4GSlR2uyx8Olpxa7j+3RT7f9AzVZGOwZI/U
0/jYXZ2+yVQXtBmELdIBRHdPAxPnUciJAg8WbGd8eXAewdqgG7zJ/A8UYeKtxqFx
izpyyauwLnQ65wZoXMKG1jclB0xi1TxD7wdeN/N9hT2J8zJX7kPiRH1hMJ/6gaMU
wTwI/rUQPEDEnJdM770kawdxUh8WGdtUeLm90rSA0iYUfAZKTk9FyzmPtKnYMzML
zXe5NU4W7Hgv6shv1tK/O0eslZsG89f53RAKKOrzsvwZDNZUf2VPkGwXXpnHSafo
1L/Fyvy/xYcXa+tDAxWTiL55ASZ31pwX62kOS1kuq2fVUvrnCByik650Gkq3dOTq
hOoy2igPcGG2jc7B+iTM0td8t0bEq26ZhAoDYJh4sPeAoPhKTv5QaM+7XfbFwGLo
Qgfn4KbAlJBk4JUKCdYnncqs0GL+58aNS4uP0mpuuEXJdgtkiuM1GK3eclJCMy77
1i5KOp2VE3ASKZGoWC7R1U5CLFzPezxuf63+tHj2UVMZTBtb8DY6WFt34NNQaVbj
qC6SwQcGpOyDfrG1o6mLxb7LfdsHhKKvmJjUO05NnGyo4mAyyBGoqHJWJepwGP5a
2fhvZH4bXMVz5xnbuL7SJ1sgIDf9YjNLaMvPkxaNPh8fw6WEaf2bximFtNnoUpDV
qOgSybmtu4Vf8mzkm3IcKYKgI+cxXUUpfEb4HrMZb9v3Qv4b/1dOQAuc3KKHZP/P
KnDbxXp8cEwZPYJISBGoNIufDOG1QBLMW90Fr0ip416jRhT9lgnVSbGYwgkUlHuU
2Q+NBq7OJGCpFFAppJ0JIEEsKlT4wSHvSx4DBs3eZDDv412/jgje3VgjGlC7E/gz
cj9Ub+zkIWEv0ffYHm1F2oL01Aq5Fr0+hRNkZqbyawjaIXC7QJWCSHRdvPqKFcx5
yhOwGxwNd54G6hpxzqUADc31BYHASr2NE7+4kwNzajzLZI6DSTl+s2/NXt6xb+67
ckaSxWN9hIMjSbWkNRiBL6aZwsV5H8u0WZ7lygaPFNGjIEfHRdhJRyiaWhRqx6py
M8t7P0aY+v/a3FpZig0sYvpNmLNoNCg1ZrsY5wk7u92pS7QWjbbQpNo4zdscSo9k
n0NbpQl9NSnGmopEQxDBUXZic9R2ualEKuMiBs2QiM091L+r6eCav9sLx0GWlfrT
r3rLKasb7790hSTLcIuSbAksYAKyDKL/e7iGJPS9ntLZDyQ0+Db6Qjf7wvn5Ocgs
iDmSSXfjfFS3SxdNItqj76DkwD7SRe8iGx8pJBQ2qmFrnmq1qV0tUuMu8lSlZHqK
o/AUH1HFeZRhZgYLL9c2+3FUONME7YrzvN83TsGcjvAbH548li+SQH8Jeyc3R/s1
hLtvjPyj2TEIVsaancHea3rS6zHeei4Aq2cYNPFYZIrVIFuMNChxD7xTMjrIcH3i
pM867XDw2SuCHhVIkpOf5s5V888Nq2iszAeH01tW+H3EtgVc48V/42hH7TWKu80I
4s0B9O4nf97Rj/UzsyU1RG1ukVbRibUcOvAtYGpkq6hXKTGa1+LlgGGhLnqTC5BK
tXJoTY5oSR0pW0cU9OsuzmxeuMoh/YQrqH5mS/DoNH4BzT7Fd79DQbgWFXjWy6wA
nBJ6wyrOwyGrQsZ6DHP8xT1Kvv2Tje6nxrTqh2cklmOmyk87elUAceTh2UDlqgiP
zQ2a7tIcsKNtuwgUhVbuhLyvaOQoJPSv+WWGvzQk/jBmOVed43Ksna/vk3qRXZyN
i1ShV8AKP0lkKJ4cL9etetahmnfoCloh43mtfQOninWC1vvSgIOBrbvpO8lGazAr
ch8cAt2PDWsBLGSPH6EqzGsQF1S780nRrT9fMe1lGF+c+RALkf/+1cW/84E2sRTf
oYHp/l3xQ/Xvj4ENqFFYFIPo7rfycIMiallv2tilKassleT3/gG3V8s+sMKlfEBU
lMltHhIjzpXE0lQxuz1JKvDZkfn2i3rPv2lBCFKHAv6X7bOd62uhrGZ9gUlbYFP1
xkqEktsMJxWEZ8puRkGkovuHoAn6tyOtZ0jUlinR8d9BPcGpAOIgrDpFT/87wCWa
d4rH5bgZPMN8ayxgNHPWQKOhwWCHyoq+FtSIk7heb8J4GRn+UJPsAFT0w+wKNLME
jEW2jzpBimoQy9CgvFsvXnmQL1dw5Ul799IVxHrAuwHYc6kQQhyXi3UqAGndKBBj
6EvRUtc7hKv0Pd0e6T5C5qYhne4t/guIVgw1YpjVGNZByvundNjmzWezIKvUrCHe
qFikfDH/XfFeBE2mcYasK+YatY6ZB9DbZSGoGC4g5hFCZNMqO4RzpGpb/+CrmMDr
MFL53DuGk+1/9J5CX7HMfBxTeC1V+bWcOAI5aVlUkNWl/jXd+HSOGcpQSrSVMsdI
X+PFG/xEU7itsNUbftCGb3LVBNRqAxa5TUXywfW94dTstvywQpAhUW6C+ID2eIGV
rq/LkLiybkpyms1wCJURM1LmBp/ZZk654Piyx+PUZnrdDaTk83jmfMq2GG6UW3RM
CKjUPJKYwDQodOE8x+GA8rTfFlSYKxpqd+8AOgEEKbAq2THcUi564Wel/qgykH32
fGVesPVG+1ayjapuV7Lt6nSQKEn56bgz6bbirqW5qGjTYeaTmzfxx3EuuDfZdJH1
WPakDH++k24GefKEvkyVkYNliyDKoVgFH8AheVUDxfc77vdK+cYZ13euOK2+C0Zi
6jbgP191sgY7xXWuef8XEqzoWYks8PMfPHTPfGYhmG3jTL/aAavSa9vYSy3nvDqV
PqUfOLXBNrtQ7cEF1vjum2cdPYRQUWlawLFR6niYDSW1EmlzcoAFl9sOzQpYN4Ij
mX280g5LeqrbwP8KSkd8pdypfyDDnYp+ssCa7BeuNp01Gg1qXBa15Ix6UHjBCnVc
2An1MzIc9RUnAGjvAW8rVX8Od27tl7SkSBEb/ltBL1ypXjepotn3UvECyf4I0Xjy
VqntSStCWABsOiK4AviKBBg+zBjuN1Nq0tOCBxTu3DdmrSnER1ISYiZciL60THSY
NoIBY2UQr5B5DJeFSYR7EYTCeIYSHHb5vgBbrFVEXm4TFzoMF+/XwHRUax5T4iqj
2f5eZMA1+6IFEH/KRqut4NgSpWDbgg2mDC66WJsLcegWj/JwaJfNbFbKBXVMg5jt
wCe0UzH56VD8j2ML0wtf++oxWTLxg00qUzgbxq4pR3dUX7XAjINsuwAxAygTHdls
c8KWqm3IE2CD16CVVIMGVcX9XDfp5eevs+7oYa/bkObby5bJTydbyIIEhpr+95xT
ix0w6ix2ap2Jr4oIMyN2fKHlCwZ0HnemnmggW1u1yuNc2wgMnNbCk1eIx9O8sV4Q
rSITvy7WT1sTrMOvyp7RsUSVkrj4m/Dz6r2qlHNqqh7S3g+uyKyHzgKFQFU91jdB
x0UkQwr4LGlvTId9jsJ2kujiC1XZTs5bcJlg7Qc6RfZjiCnPsMmQcyiKa0cyv77P
0IcmTrSKCOtMKowN8ESaGgIdsrS8JMdhQQDLrb/QnSq0zrZvDs5/b1fPQ5w9FORG
BCDjxc6SYRfXm2vNklv8I6OPrHy7ofi/xJQhTEtZm0rK9uyXLHAVj4QRJh8qEJpZ
/uuu2l0Kg6Bg2L6a56H3UNA/rtNanuYXmDdH4b2/egMcFz2sw5yPF5N5qG8T7KtL
XXsCSuCUoMLDcPsOZ9ZaUjkFoROhkqfHDw8088zMILi1GSB4tNKpHeTqWffab1bg
EnFH3kyoMScriO8NsT/RT69SMbxcK4bmnCHNfoJ2XqeqNy9lqrsW7qDh6mspPq8h
3viZ0+F0LLeCF3YEfSEB8vC1+/AK7po02rgzCFRTuF5uLVjzv3HiXmADLzBjKPyo
TZzZ1XE57Bd7jMt+l6MCX+WRZtiyOiC5ee2mSdROX6YM0O/lpb0rx8XUQ8B/sprh
zcP9DGVpOSF5ZMexSPGmp1rAxCj7w1oxyjjyI56AXM0EzjkC2cGAXVecB1OdDOXG
Z99oiD6LxZ2ATRtnslEkh62Js25y7HoBdryKt7gi5nDkNODxAuVm4lQ+QoaatrBF
UgNZKoDWK06Dt67CdODGolxByFdKq8W8g1iCh+XD7DZMmH5hu4UdyDcbYO98wRo+
aFie+xjaEsE7zfeFWpg7zqZWVh62fd61ccUHd2hwctCGGDucyfaCic7ypL0thX2H
Ws3mbn9gKalU6LQSLOBNU9ky3BiQ2HksLc9iXHdJF+3yxzn4pTg37EZd2plg494R
z8LmglvQl2PVdHoXCL2qOa/T1rEV4PR3ImrFCToz+az0HaLBzm1nssN7A8Sxfuoh
ADOQ4YiCJP5J52K+eeb+D3eHaVNxxd1Jm+Ut71cKibgkUXBeSolGj3IeB+L8x5Zw
cIFgewzwvVVgfjECLCoi3/7/h+zV4ONC6OMStrkcgLqQaOtnL5ZYVkfhfKsodDPi
9B9fwc2bnQPPKhnowPf43NVQqnNvrmEnrCPHH14F543/iIniCXLumy9S32XTcjed
spP8KkR12blt/qOpmn9mnXHuk+rdXtr3+V147N/nly7C6LgX/QYJVRIry/tbBUwp
8nEp2tFfgo42YxwiG6nHECJby+25w1+w+neQMO84Q2v+E8CgTzpYvrTTfK9Ut1s0
VaLxyLP1KH9nApPFOS9Ti+ATMEu83kTaUMBwsQFAU6RSRZabfnc+SzAKQ0O9SkRx
KNCsJAzfuK7FdsLb9YoPkNNzyt4koevnXYdVZhtazkGeCKj6Xp+iP1f18xPofNlZ
UlI290mPCUKsasQrzwSS1oIznKrbO933BLrFSv9cY0M6GRGaID/T1G5SPYu6CxDT
IRtJ1qf3vaA1v+ajYeRsjMtEbxNrAuLz8lYUr77kmwFqFU3g96/POmJ/TDDiyFyy
Q0b5dpGldxLBtYu5dchykDv6xobMejj9CE5iUmtylozSDrNuv01nGSwQ47WkAHDE
YbRHDV3xyWTHWkbYXrg663McHeBROYJHxjXwzoFshRnyo16gMaG4zpCPDrRRoQ/+
mk8WialPVjHC8mi9a9hzNJji/nNFlZhIf2nv9sTSsDJHpYRRM+sMptsJxZ3fd5bf
ac70lWB2tBWmbt6oJQTXieh5uoHh4ycaTyKAsJ05OqbR1tjzjY3H9DeWIwkFWbJg
Vcvy/dR658GCVLLD1jL5m3zjYGwFlOGLfLH2lUDSvq36qQj0TATIG8uR1aNGBUgv
kXlabpdj5iT6JWnWG/K5AXKIR6nvZnFtibRLlQcl1LMVBf471ztkqQEZZPGqa63e
jl8M3d+0CpRppMWzWLEZJoIaA+bIYVUA+ZAr42HZOfORr+qlL+5H6up+TdPfYOWy
65EA6G5TVwXs9psObnD4PnuTnom5xmPuj//KfbcVxVJJegYp03SNqRkyerVQ4kWd
wVmTsvq2SQJILywMX9dZ/Y6nHYx48gaeDjJlqJqr/l9sObH9Tj+oXuftfdZUpIIq
J3pb/tsvIg51XV3lQUVDyL5lEMiMycQTF9nGzXpexv4eIXew3c3UfEWL6rmZPAmj
ADrd7vBsv72XUICnI8Ox6gk+KxIJSnLkEVKwUHy3PZcLDuXBpf5E86L0e6iM7IWz
Gm3UcNnnNVtP1izH+gpA42lYS5YafrIjUAynDtl7lQfe2mWLXLnjDq+2MgSVKxq+
DEXNfTKtAlzxWGzZaXFU5+o/Ici4nnJYtYSSBYVrhT/sotfGrGxNu6VgRr6uGwg7
nkROqS2cpA/AzzSz1c2RKw1t40ADR5YUw1mAqkkoqUrPtblB267AJZE2Z2TFu4ze
y1tMvtPCtbCq4lCACYlOTYZDqYCAoW7Jidn7XMgofmJGPLUur6C8vCGu0Y0e6NcC
NfKvX/jjt6D3vT8r7T0Dl7FymSN7TqAa0R2g48Fn0x1OQgiKwT7H/sGiOPjSGqPh
ao7hpLpcLC5MdG4j9g+HOfwJ3BAIMXIQG0+JoMU32vFbqrPm6xqG/zvPTESplYCU
MmU1nMT7BmxCb1VS2BBOYbXeW7fBqeThkibwK+URtUiT50eTw3iDiF5VNeiGDheL
LWkGQxKWlVQxCPMlOWwYQZVUnLJXjKFMZYVPvYW75aJH0sUyDT2caxQ2copA44HY
JkpCKovED0Sho4PgWvfYTpJhSwh6sUypi25dJD86KjwdJAMFm0cNyOQZH5QUqq81
1rkruIQ2MY+T2B3pYVmsiwv5SoORPLYusb2q+PPmuL3y4/ND45L1EYio8JaDSvyM
3ECtPweFewlAXfXCp+/Fn9YpJDMRvls9dGgfhlp4tRQr6mknJIql8IDqT4+n4q5a
0s7WEMsqy24BQR/o0G+VHxJ+l5ITSQCMcLOg2zRz4ExfEVWbUL+GGgyZ5PexeAFU
k+Yi4xmN0kFEVsexqOokbnfUgTkJVXZ2GV3CpUWL+rpcXKG/EQSqh6MFyZys3Uoa
UcJETOJR/m+t20b3FmUDvxwmsYNBXQ7eXlaN3hqM181uhaM9mWR13kyRZb1QY3ek
hmKhkAfKj7k2Oh7uXmoQUoiocrfuOah6QoagpUZiKOAjfqPNJ6wyNiQJdiuciwbE
lRfrduOSaIecAUFfpPAvA2SWrn5oUTAt+tfhjyihJUTOADVEithCGI9e+6rLXiyK
qmgs/91ECUGzuaONzEyCYC690OOZ3Fbb80DavnzGUZdcu/Y3/SFHIV4IBNVZ83t7
wEe2mV638vKn1eH2dJxontgV6ZgNdzWRjuLx/VuT5fdAlqHJ53LN6MBbFgoaR2GQ
n2yfdxEvcCVDkiWWuZT9HEpHFnlrT8mop8BNSqzbVYKP8DSYRv+tGlLRVqV9HkPX
K0KLfT8SOUaGAulCgXBTkb9jRm5yGnon21BfjKT83O9QmfEk1l3Snikr+7WSOkoE
+h60WT9BE4OL6pAXxqFK9KyWGfLo255F51BXfzsfjh0jEYdxH8FZmZ7mpsgkOw+d
EDHOAvj5m4ipxADO8yztcbKSmvJMue10N4GXv6AC01iaHPwThP1+mwGE0xuCsH+5
/A47DmbbliAM5KX41MPnS/BCA2LPjmLEYDmoax91UKK2o5lOcAC2tFgsPfo+kE4k
CPsd002TfwIHRbFSz+acZThRzfS+N2U6nCb626UlWMTEHNxBW2lJRzPkHGMlcCZ5
68mSqTMJfGT7XyKOasQnBGn/N4kMrqa/HQUuDem91W3CK0zx2StiRERmVrR8ZQb7
Saa6wJS4lUsk7uYmXovIEQXwTJ9dizw/6YkmTM+IM9Y/+c22STu+sUn8lW02VvFl
Ab/ooArAltW6KDxJ4OLhMl4J89sShFqstnDNSjzNyyurBtXSK2m6Z1zvzi33EZLC
ILwvQLtC/6YYvc1xpxY8qFlx6EffpDLKVJsn4lvkNH/sp1zr98bNBEfV4o2rGbeN
WUVtSSAuSbPUvOmnH8FQAwNHhUwm6oEiYwmrm2LJXM9uamACVYFPlszOs+QoqEtO
9t6AReWxWdbCCAaM5/m0hgbHpEpdURYe86RX5iI6tBD3+cuSo3f9r9b2tyawnquY
es+ViNfpjPIXYqDwqj1I8pQYOCoaGkKdRK217iprriCy2V0UonbdC1f81hxzmON2
0XEzTNGQ92mYF5D3OL0nuwvClf2aqm+VOqoT85ri5a70pRcQI4JOds9rM7Cj3OSK
imYZ283+74mRFkU2twDy0yuFhsp7WVI3U5WeVrcRe3wy9osBWJoJgE3vU4FGarKw
xK+8LbxKuat77sUILnJMd+isOJIKVu5305H2ZDcbjl9sVShqPUl+9fd1BxKTVU0T
CyB+BBARRZkRkv+mIAFhoDOmUh17xK+AgDAMcKNGwZSanCc6odPkmBgdK9m7yjxI
i7SZdClsn/beNOOTf6lXwE1vYFn7L1aZ85pUJ7Eegw7D0YdAnJUo70aD8XYRbX1P
/5XxaGKAdHtYmGkpRQFLRelpjY/j23XDFdJsuBGvNHZ3m9AGl733/uxdBYn8ri+O
UcBc0UEmMXT7jx82qCPoshY91f/6qDI85zw8yHEhHJD4Y0x4liTDZfq4iKMGHl+N
a2pFeV/e6a1zvWBlQYs8vYcQ2wGQWE8Zia2O8/4r42+trVWo+2lYX3x8nhBPyyty
59sLE79DJ245EppzNtfslhLrME0OASqRvYrZlcxqID2bqY8uncZmpuv1idgi5NGg
i+STTJ3g+O4xZqy749dY82Rd8jZkjPfZSO/qDh5z0B0QYD/TLvX2Bmt/tdgQl+2w
pdu9DSlRnkqt4k7o3uJITE636LyIN3lQLbPhLz/wDpPoT9jE17l9eH/7sSfOHTiU
/m0QYb2PoxySflhbnjuLOKNBC73dYx+xWA+E43F9pJzXrOVbMdNW+kUZbOg6Yvnr
rBEFJ9WJTnuFiArJY4GfoV3Q7u5nFkRCW8PD4CXSKEcMK3j+AcHKl3N6gtP7sJYz
pnw5clUTiNCZnFoBavoKAAxswvKWnokKgY5MQZwpjMlTuDlBOOOq0v7Kw0k+4HsQ
C5hi/Oz18TN3aKTLU2wyXjkKLFUC0U4zzt1yqORK655VHuEH9+yZK+yP0RrCEqJ7
jRKIPLPe88N/q1E04pJiRrMc/S0X6547sJEn7G7sGh3vqp2USgGaWBwOBTZe2wzZ
Id8Y4ynC3WMjvoPwLCX2GyasrdwGDEAaX7PWzW2VrO3Nnt0bbHBWiGqOOBj50YRu
/WZUGaXH84hi48B+pEPRKxidy76EIZru5pVqR2VhccjIC4cOqXOx4SmqsE4WJtcO
oMCEB8t+5frtV2e2HE5O1utgbUlsfxB6jSMuk5Nxo704QUBQx7J76ir+tnwSVQg3
Cnzxy21qRxsJp+hNaYc1+gCJ4IZkLa1kRsLtZBeDGpI5964yYBrTfjqJA3DAUAMg
VZelfKRBd3LUODS6NpeyOObXP016IQcSDXceKsHqyw84JJBnfGuKf9azYI0qMJqc
Hi4P3DaI6eeKkGRZIXnUoAxSdRQUNRLbXTAZL+8VScW+T/QwyyJsszRlPqKVVL0b
7YKEN3wE4leNZKsfPRdrpgPXvZp1WK+z/6tNwBZ52KK2KvHf9U8wa3W6z7gHUQ/O
6+SjYIrVa4h+b6CSy1GLIwAWf15jGxBruVULanQI/oUAcg6k1gBuJYp4tTQFHMvm
D1K+9QMuTp3OXc8JW4UClKyXjsyrVWhi9zQjYxBfY7JK2xaV+oPQQH2OWyOK8xwL
llxbc/lhMLDYCi10cWEjjdvJLKLB/FuKSVUUUhi7HvcIzTCkNQ1hySbj6My5mN1s
VrFEGnPN/LQC0D/7Z7m1ruJmpPH76UxNhNo50VuvXmz8th7q5qZGKc8ohHEAGfN7
xddXrikexKQZpptcSgz0kJ7k65VzYucONFk3cqEB7UG+CrF24IE7WIa9d5nyjzWl
o6taIY/e+9oAuFCljIEiO7NllQzcmWdnNZRgEEHdTVav0fmBc2gUkLZHaWMbPB+W
It/c9Rp5tw/RwxlnQmLNV9jQt8Dnl54CqXgGqdmfVfCxsQ8YIiDjdN5DJMxPsBiv
WaAXMHTJxJufnk5604PZsXF1F+T21JBl5y3fGHGwo8RGeaHabyB+xjIAAjAxWwdq
TRc3e4GAj4GysShYs/DhGhYPEuNBigbUEA5U+g9Tqb23VPc4l8uVDcjm0U3sRwAb
8I5a35mwMxnWgG4z5JxWi9kxpi16r7fLIASh5gE4JtLy95uN0POLHaMiX4xQtXyq
at/8VgVrYnDl1Zo/MMTILhrn4G/VZdtZYAEjhFLpmGHAMKTv3nkxpwt0Ro0WFQgl
1lWvnYxXGAkIQJW4SaGRA7YCZ8P/EhlxJq7HfZxxkJfhQMTzVR9wrdjAk2gobLr8
zsL7Ob8SFFFBvBYfNrqIbU0Mfw6StXPvvmrUKjwRR/XjqH01iaqSLMshgEaQLINa
MhvwZOSVS3r9x2xptp0vQ4DrmTVXqpU8MH3/Qhk+v6p/Cpqc+rwzMuSS3985UVXH
ZvxjsQJgnENbpZLnYi3L7/90NbfwcbRa81aTS/toVnZ1Xq8+GeDk0oDRtfASVclq
fOOAYsnCbBvrCE1sw0a76kPOTbyKNo/Z2qbjYJmCnAi/QN5Vo7jTdrjTsefKSWBW
bL6vHkluw2jjTHS+aiMKRgOrBjPfKREQ/Ca/pHAP6ByFLu36cR2flGmBaI9OaXJM
i65DasrHvHp+2GXjtUpmAOOrxhH65uaXGJvaB8H23npf8sXfa5PTISP57g0ROo4U
APRTbqslLUKrmIzKE5xpbHkHmt4J2n3wIM5hotAtN7qkiE2U44UjPeR82osjuaKl
9xcSObr6FZ6g7ZfSaPQU63UP9d8n8YGECbu7bv8M5+feK/mk1ED9/jRDirruPaDj
ihnKXdrSys1fuSFvtYGCCt4DZG96g/dKfeHaHI8r+PMu0Udo8pb5ixt18mYOXnSu
ddExoH2iGyAdOgYOrcMx9jX1Gb0d8CaUooetTsB9+SGuIQWNKWF9H4Pat2t3ysUg
lPU3+UIAK1n25qSexL7MUPVckdDAMmmh5/TZGItt7hsJnLoetukk1AkQ4GaD19sw
Y3TYwQmnuI31FYs4KrhbCo7viZv/g+TmYdnZs//Op/OutnhFV8zM2F15DsBN/K3V
/NNWBNXipw6WX7rxVTKD3CtsqtfyZl3LfeIOUBNwqCCwES05MsbOdaVyYhQxc9KP
V7gYepr1ItqEOhq9unLmeJ+T1QTOxneGsTdNsdv4MrJJScavlmcvA10R41iNfatv
GuGZbLf7w6aulBheJ5VU1mhcE4CayOxUiSesmErtzeNJPvwN6vdr71uiIsAOEwzB
ZhOR5NAlMn1ZLpkk0aCsRgisWyeIfZp2HI7ZH+YeOkXhVFvgy3FkpHdEa6tpUjdc
3ZcWh5jB6vw2Ty4eXNJGpgi89g3NeYv+dyDg7PWYI7gzRvoGGLUq6jFQYxw3970m
aDosXRd53qmVUYZFN0988nsz0RDQF+SaYajRBD6bAzhJP7oRe84TfPA6M+wBxojV
4j+XB6EOYz1j2IF/jum+74wMIYioqXqW+qEwzR9L+/xeQfcAtc/T5y4RjHGQs03c
v7sz+5fMMiE16wTor1O3ASp3n3r4SXQ3w2VjDrQcQatNnLti6+2gok3fHgF9rHZP
mc7ywrT60ziVg0SfyhBQbulbsVhdBh1BeTZG5aOhUikdze7LQ8hmA+UyH5q/QfNn
6hB0unrUrO7fZv5kN6LqwEP/MW7tX8hFBV8oalKsfy76WInwni0sXzZ0EpdwN4Ih
F8QVQVG9qQZVFcuOwNZmUl0yJZMpFyAMZGef9XmrH5ZlbWapUuygBouvOB30Cyu6
VapK1GAYcDvjhXSrO3BNWA5iPsDHx7Dg3s3et454FUmOPMvQMRO90q5o0oyGwQnS
zHoCLxOjR92RlCdLtcsKvP7JTeqmBhLkJPonTvhUyNgX94nulsgzc6/BENxPHFz5
NXk6Dkj090QKalAA26waBOGQcKlM/kkBjxjjyYoP0wOYMB8u4GgS+oVPwWKIeCIK
GIC7rWCooC/r9UVmSnjNpnGX6QHn+qLW2Q9paSbJB5b9OiISHfliSoi0L6gz6p3w
pF63OKxUzBZSphQvRr9q28gTc2iFS1kL6vNZgrX+9CjxHg/bbnHKdGk7nLTgLEso
rb9i0GCZGHF4bSRZZHk/xLqrlTQSAfZbNKKQPj1Zxab6FYt8uX8ukkqGaCIB34c3
qsNZ11GiHO1X81UQDEMknPuF0LnJEwgL4oZW2KccJT6A7I3UZEAJ/TOAOUTd4HU0
FM4vgshA6bRzCfPJ50S05L5FTycZ+w/hm0eeasti1gX+7QjU3c7eaMICUN9iREps
+6xGEFpyis3k1vnzSci+rHyH5G9B5uN5a+PS95YajS0cA/AnqQSq1wZN/vE2+psh
GdTTU9merMWktxbt0uI6UnH3K+mrysQbV3fJUtYRebtsYB6+b/xjHP1pMTKj6A0c
2gCydpPnfnZ1bIW2SXAR/ifXFFedkRLTtUa7tLxszFHIYcKr9HdjXpaGGFPz0OQ5
WGhuwdJnf3YK4mxgSExo1LvhjXz6uaiBL9JYrFkRME7EEqsKBTP0gNh0C9tjDlM0
Y/sSYKPaMjiAxEPlUSkwBsxi5Cye0B5QndsenVda/9txIVUeIcnbIoQQRx0BtGno
q2ALWpMduuIN1WLAu6gVkzS2Z7J40cTdI4dopAaHSQbQgjD6mlgUVDyzMdUtszSo
sDdpqDgdGnMImyIeiGgpAVJvI4Vansgs/5+jwuzc3US7JxJV/5ceOjcuualyADRv
1W2eT4N9Br63WrRJemuz2vEr9GIWtf6fGhLs/Yk09C/uSogqhFmnqAUwiofPFTla
YJGIGQxVCHdWGVH/5HzIGJkMZOaEN4EFYfSgw1/N7jsbE+7WNWwRyymeBW4KSgyi
japVSdeL3WbdUU5XqnIwD90mTwVTyEYFz6nzRBi1vQJm5p3iZQqTJvnDKT7kQeqk
Bsijf4fG5hKcaIcbVhWw4or9ISS1/yhqFXx8HJ4FNio5adIl/K2Oj7qv3AcbtqFI
H2DU5AQYz9mYmHBgsY4fiC93qxKun3xNGANVokA2yox6qbQQqg+jKCXbfMCbN9qI
NCVchJtEryIl48jubX0fLjq2FHOtfuSqCrtQ0MF0c7V6ezbUnly5clrjH6/1x3mp
Pj1Liy4RBM1/DepveijcCQOej2vc3yKaBmRgWvF2jqY9MC1UgDZfH6OaT3wTkk6l
4v06wnOObvaA/jMrX8vQ2iMnaFRHZWvw0Ojmx82G2UNQjvR5keOL3QVtoPl2JHoj
ex4rAJRoB4s5JjATSvLCV7aSnvAaMKrX0nHw8xeLobGks/L1CKt8Pj26kNyNOJVd
8WA+VxmWx6L3Nj7WFEnwm3PECXwf35jfabinXfBe6MA/T1FbrHqMgdTmQp1srDqC
EOOxEZublSt90RTBwqsmh5XByMifakt+d/qzSFNRbCXeGpe7P4zP23SCA2UksWly
5rh/uEPwrIFcYiHu5FjsjVsRSEsT6Ud0Zs7VZbkpKQRM3b5e0FK+J6NMQUf3CK+L
249GpAdLM+s+B7Cg2cEznmHPz9jMknRZmkeZJY+KkSJfeG5xIWszb5rSatP0wvBr
W88lzEqvPU5neM2kENHX/nbqO3Z28uQ5R3siw1UVd12wTbH6J+kw5OKzGYK0zgwZ
rQiBbzU1yYX2w6ZMvO+/kpgEW0MCw38H/yoeyeHfzCGGms/siqYJ6ASq3a2rHNHr
wtc3Pe0oDy8ocq6ly9AEwnjKQcQFYAHeeNPvAqDiISoP8GrLmBV1TyAYFH/fnb6w
T1tAkmquqbKQchaBCXvkM8HFa9gNob2C7xjT5OcwNT7zrS4+VO1hSOmmzuE66iId
osManET/4g2R18ZSp6YkY0JOr6Jye0Si0EhwddYs+sF23tkKrKxoMWorXKBGRf3D
pz3E3PG5/ZbKUSWvoP3iXCAVCRQIDU45vltKCOPdYxa9zN5FbLc8NXxr7ZQW8K9M
iNLufGsxdf8nGl26osCx1IbzQ1TxP2or32xtdo9O1lDZJCsm9CJvE+/dhcqg5fyQ
GDAo9EYeXJblKWWczoXiqZcweCo6+xQWgtee1ebpHYuGXGcKoZ3G6gE6/pIqZ1bG
Qr1+cCso7HsURs9fUcA66B+smPG4YaQiz/TIet/Ha9UYx41KieQJy5rRz/cp8m1C
t8uO1jjqv0O4HM5BcVUzmTMpywnxzg0O4gx+BWL8GQEhRxtsEN1jRDJl5O0caX3k
gsUg9tYtzF5a4+jxlrm6PwgPS/KT8Yz8j6syLzQFGTvzbpwgY/Hw6QRK1rWyBtUW
OlxIQmpZUC902e2Rn0ctfhpXoX1Z+OlmEPbzCfVX+UegMe0kWSN0dKwNSCI7K2bB
/V6rG9/8stRD3nkZwOd2mNoB/OqxAOpr3++JbbTTiyyR2Y7+B+4WELbqMuygFvV+
/zvN434IRa//q9gdONFcxBJZQBd7CiTVLm0MwmHH+9VUYy6co/u+ELoW0k+CW0Bs
tzEE/GSEVrRAfz4U/zgczqjHtOCxPgXxWHnt6hTZzR80DKe/FOGxys+QWoh27qpG
avtxIx/mc7/wMRDGLrwMsk/xM1tcbzX10tvbsqmV965lOwOvIJ8G/qT3Pp9BtuMd
HCM/1sdg55+0gRnHlphsZesaO1AuUXD0bLbM0+SeGrefHGrmNmxAMLjdSdBbUfTR
KaTvURq8DMRY6Z9qK8lgy8xXwTUVcfn7GAHed7lonBiKIbvdS0IiHBKbNzofKW2F
1rJr3v9138h0+VhUhlbXET55sRLdoRDTeiPTihTa07eZxw9k8qqUuj4BgEJCxOMY
iowMdhMpQuOhr51nhNU1LjixUPM+hxMG4y5kN/6rS5AqejLUUc2uWPa52yxYsS+B
phUC4gRHXEE1pBwVjBT4+rrzZpwXVTnfrB917jvHqjH8zUcNlkZqmA2OiaVpnKj0
r6e8jb/cMPfseTlK0fluwF628ioZXMfdv6tQdPXOGlFYUW1OG337S8kvehgoR2nd
yejntMGHJ69XQRiAGWGl3/ZrEmOFtI/2dfI0n5oPuBknFkG3O7wwMRA0AlyYW6Am
uSz9xuSIs8fOn/9sNSx+f2AigAbJ+DJbiqxsmlnyt8XPveVHxwX6B40hoU4sE0bX
/9SiK2HdYzeiGsLdApnFcJcA3qaBx01jvi/362UOeEbPeucutW9NYkBzoypgUyMM
QqTevGSZh90Q30tSqsT3qh+w2NKRSoyzgClPx80s5rBrl59D30673FlJqH8w9M+I
VU2K5H+L0t6USJBoPYTYUF0Db4bt+S3srY9F/SqXYw7qN/3rZQBfsAsBXm1duPRt
BpXmh1ifwcr0V05CCIqR8ajXv66tBv5ok/f6WLKE0VS6sEblz3tbwtoEvcB8vxr6
NuoW7KWGo8tCz2rxlUSUrvZC+DIDWmKT0/LutvyPQkpSesAlZHBfwWne41wtpn48
qGWEp4P6k8UkEQEgQ23gqxv1X7d9Dkk8IaxS95i7tBT7q+PugSVqUW4CIxgggzwK
mXMcLOvUbUTGilu/QmV+/Hv7EuqOjkUBhgKwUUeGDxt1iA/ZrVhhr2kzakAgFN/O
2ZqaWzIJbCQPql+yBeV86IMJQulc3w3ujmIvIdGf7/MZoa5YBEMI2rw5yfM64iHf
agv9FileI9RkzZW6Wyj1zzdr9R0OCCSW2T5a+R6z47h0Ymbc5bC60DjqFDD76Wqd
3ysgazouC3O49NuGa0E4XpBuhQePyLF/s2PpZDdnhkkFpKWVoojwR+0bIifZW8rK
4i/uegQpNoG5f+9Eg9ANfSgZCtGm70Va5C3HyPtg5u8k5uclRrDRlaiU0pLycRdp
LXufpy935IV0k+Uw/L4I+0zUfGEmrPbSYPDxej5xTmh2bKuP28wOb9S7szJl0ghh
5fQx1Wsvk2MsRLBbr8t3XPHneNddDXEBPxWOALdFcjTw0WwauSTD0XPZSSLlpmGF
8SFWcqMZzgVH7gbe6inEGwa2QZHImRPkqnSx0rXNLXnE8IwWOdA1dk/xQr0de5dx
izVwZarKyUoqQpgoo/AjobwML9vWeonDOKIC4d9tKOggrblraViXrBQFx+SEo6fm
EgKv8xMilBWQLlgPMRSQyNwTGugiWI7QooMRbUuqhfN0pLhyA8v9AsGTq3CQpLUy
DgX37wqSC/9YQ7fXQZBi58fpXuy74PctsnAXuvYQjKmP7j8JKlYECb+Y6ivJIlrD
mAoXDPwrtE2Yj3rX5Exq/k2P5R2C2THvisfjVeWSYGn50iUtDUWTiM13Bc8wezs6
AWjczW7/Jq/atyO0ZhSSqFnPJuVC/DmZdhCbytOmHJrqWdEocl8KWjT70Zu7ae10
7WdnxhXysdAJYwyLSXZ7HqKILTNgWbz00NcDfzmIJodg9mkM48bn+4M6weoh/BwD
bhZLf7u0Lg7GPOIHT/hBFTEHgzKhLaDlbsMgV7cI9e+Lrb1f/1E/5zgm4cuwGOH9
Kga1dp8/Vm/mQ/NU75V0KDhspxHo4hNz06nUU4RfiQkffRTA4PHV7WODzlhMGjrn
l/w8UUT/Qp49y/QK+xojbzgxdIoMoFP6xrC7UrA9Q4CNUqiYqJcD6oPnovBmLMTd
bgAkAwNsXm84cKWf/E6ssu8Bxj7k3qrnVIQPHAXCeA14wiq1cusWRY2Rmn/PnCWL
g6Yy/Pu8REXAKyCM0HRZnyHh8TN3Z7dBW1Xe09r60ScBGLEYNvIKH1hkKut1KToD
52n83osKl+BhqdHzXwNYJYMo16bkzn6HaFbb40oAhFqvUMFWD4GlwYnlDP2r7tcG
Js2klL5Fnev/t2lYtE4jlqGOzCxI7sgdC+0CMDXpofLlBZEbkNM9djYkGeMagkIH
rT/6aOhy7vlP3+gNX005BnP7iP6MkpzQCmUjPdSwjAxcx6oU0fJWuSbSDlgd0vwz
F5SFF2phGEs33kDqv/BPGQU4qqpjEoAbEU6kgn4bE3NZzAg3hhf4WESfu/zNNLT6
4ZjF1WrF8QCN7xsb7rqOHnmv50RthVsHXizVNo+fI2XqtvqyJB6zQkW8OWFfH6Tj
LxsfZt33tjI7+gNEibBt1JWqIEqr9BvZFN5d5+ya/+6VJZ6iTnLethb11mcURCAs
aimnMnAIpONllm769/YglfIIVjzXsp5Vai/9I1aPTHd/auVzT22DgCTBQ9cgPcUB
+y/kh/SULRorOHeYynkv0UvN10Sgl6exHXa6e44mpZIrFKRE+IbehLgJm4XvKnHU
wtMfnDtsKpm5coGDSHoe+HZaDJG3rKbX+WauvHl8GJ04O80qhdl+6qsfKr/gxTK3
Iojl/DKagGusdHGD7QMWd92JWhhyQQmPEYw3xA3jgPhj5Qhsu4/a4TafQyAUNgfc
QbIXKs9LTgRAlSb/6o2tvVAUMru507D97QiL1XjDFcxq3a5Hn1JYOxKvanCkEk55
TAtD0Sx0LvJ5PQ4x7nrSPNO6ij60a7AWH2/8MUP0B/pc/a1IK72bjZC84iyZO1DP
oIQBSioqnEIWYfcEGiYBIi0kNZvGM/35yiblIUD/AXFVa3pphG/EwO5IVMlAmgCG
pJQZA+blVOKBF6OLBYlnkgP6KSmoN9WhJ0cx6f2afdOBhSRrVJkTb8yjEBtvLOKG
w2lWaeN+MHRcXXccP9X91Tf/JuxmwCFuqNqm549Qkreb6RL/LCLWjB17CVV0yvKO
SPfzcM65qwzP/fStfN4Krykulu+busHyv3l059exR++4MHzZBaKUpcBynzJ28gzh
rVKVbpgYfUsc+OvT6wTyc86TUru8wjSm6+koKS4otjz3wcoxzBtEjw99wPgdgYG5
BbPH8/8rcwjS2hnJBHY/oEbW2xdlJ+gRPdeS49nFwH8Twm7QHBnNPcLQbDpnuaox
mzRlQ/rZSJ1WW5QuP32WxRf4v/BmfEc1TvyhVXiUI4kn3r73FQzEcTXNZZO1Qy/W
+hXUFW6mLuzm9wxtmK2DGePwC2oWg66/yNyeMrKU1TvjXYD7S1A+OBvvDxTL+PqG
0W2ZRBuAYhmv73BbwxYZpY6Sf0nRiqWdaQ7EoBwuTERhKEkN9d75UnEbvI1rxh4F
hKLi6wWDyWhLpWOAcmkEOu21DpJOEFgWnpA0bOLQbaIHXm/NvxzWFX1rF0qg5aof
Jww8mXKR6U+D0fZAVJtMGLO6+L/JObiJ/LAcUClRsO/4Y+RFW8dHlI50YvvJ6Sau
Rv1BT8GSBRQZu7V231E4i5u4qBPDCAC3VVBh4IGECJuB28EnJa0DybA14N/PxSUE
DtPRs7tQgbJuLLESTSvT36evehX51zRipBm6GUvdIeF7rrACI0EmLf7L0H0coK6n
+qcOYdJG2OSI7Y3mpItSLd4vE4J8ZXO4nM5FBqblI9SuptX1PkeA6YAauxLNI5Av
P38stLT8Owij+dKrEbh4EmHJHzhvQS8hgml0dRQDnEZT3/KpXXBcs5IeTr/lrPLx
mFwsKYWMHxFASHtPkFxVTvqz81ybUQtrHSbIY6Bb7SdikN1OeRHmz1TQpZgHRkM/
qdU5BBwWgD9LtqB9NFtODSrjDX0Ao0O2scui9pgWQQD/uvsS0jDzKmmE5HS0KOnz
Owdi2+FeljAsl4q62+i/69kyqnxclPGtHOsDEJFBHYm4PEkfuLeP/pv0hpsM98+q
zNtTje0/lTqs+6Frk4Sp3U2+owmtCLjLa9iKQhb5msC6WxbWENOq4G4Y7/zQj7f7
Hk7IMhuFbh1UH3YnnP44f44y7cKzfMzXE40jANA7kD2tNVytlvQfMGdk+1zu76u7
4ZN2IQTxgjM/H1BmKsU5ot8suucaZFX8GwePU8d2T+wJz/yKPWIGDios1LVoXtt/
pE/W2qGV9IPQXo8JOr1bvvPuRotcffrUKJB9+rFjWlsDhzzw5CmebbxI2X083LSg
dgDBd88DfuDw6b0Q1c1r29Mz5gGOra/o9M18uz4f5F9u+ajDvgJKbl14TV+bXcBv
9NXpTGCDBf0wxhitknIAxEv0kqjfurxtSTqRFqV8/y346m7BR7HJqRutpElBHOm+
f7TKxiYjWeJ9Zx8r/Ckap7fjU1Xx3afxNbNfgvcTF4b9oi2lj8PdK5JEk2zYaJ5m
sULw1V++XOC2IXmrjkW0HeAv8COo32tKoArFIJoP57wxPiuUPXIGq7jm2vWEu9Z4
nPYi2oNODtqjCjSn9QhOoJ0PMwMvJsBiwisNlcTMyKpP54ClTS3z+q3Nd/RrRNwb
Heu01CSHFs9CEPqABDNeEBLLOUZ3pmLOrukqz5T0TeUhCAZfD4XfPGH89XPHVLpJ
DKCKciVTbDd/9qOF0Ww5KFpcuZPtzBRlWiHVEgBf5FNeMZGdpemZysqjrDQDVU7i
VRj8W5Ckqy0VYU2vHRxckL1lTJ5lVizPpntSeNBqkft4Aw/XkriC0AP9b2jejMWj
ovLJx0ZaGCu+A80ExhJhYra7Z5F28ykGsKBoYdlvUOTcXL4RpMyZ2PBee0W8chcO
STT9fiE14+Xk1Vl/JBT7ia6ml348aeFoFT5H0TivvcRtv18ohzB/Qe62v8saPipU
AjNg8/Ma3cN1oCkSuDwCVwbu01i1N+WeMrifTCaVeAIOAL5mJb8nmtSdrea+EFxn
sZX0//ddTqOkS5GrKjij3PUjn1DgFVtJM7uCEJRXhupd/phRjEH5J4y24VlGgMpB
A7kW/mjnDZGreVgrVTvFGnHllWfzF3F4MItiiSMYFCjwCb6zHKlomPZobGU9Yvss
wE+/6KM2oQz1rH0VRQIU8bTIZAZm7f5IO/12ggIO5SU4sDGsVultoAGFYt/yxYi+
+5OSit74TNDnFvzsQbq7UwOHhxaGAe8bUZlWiA7JuScEx1xM5i7h8Xv44eoJJ5aV
PIv3Yf+iEu5/J9Yc4RK6B9yNv7yU4wBvTzEbrVorNWqBp4+TFw5JPRoWXuTgFjle
2PaetA923ceMEGTE2Iv+GYYFltm4B8n/ClRT8HoxGrejQ9uGhaWRJStPThHrI4K6
da0p6N5nwCizTyXjmick8BCc5/3slch/Gt95+oN1gv5IrwFHTavk3iEUTX1wdF9b
rzh8BBsT39gj1MbWXRGfyXwciQk7t5svMx+s3mzKRYkvtxtMrC1pH58DYnBkB0dR
P4RWPhi92OXtMvpQa//uN0C2IR9rtYVTtpz+2y8RBI5UH569bKztpzqPiKcbPQfg
B/Pp7hj8kdSAt8dsI0GaBZNOeXhS9vn+X/b0ZuEF7u0Iz6bdP34l3sXJocrwYbeU
kNCwOPyUSE4TCf0FGa/HQQ311uZiLZSCQRqc+KMvRtGSrE5KQdq4evYdJ6YHl/ID
HoC1V0gK1JgL025ArcvpHeVRIpzv+fuZqOwNsQ4phZrUuUsbLvZ3BYJukXof3Inw
vZZXaNoAu3Gkj0+eLEAddvwWXOlsK92TcpHMEW3RTR1JZsGSEOA1q/b8MDHiDLs1
uQI6JW8UC+3hZAhq7/xFtEjRElqamaVkPCTMfoLbZB9iZ83hm1wgIljCGyCxVm27
p3XNbCNWEcSq9jfGxRU+Lg37hRR8OnsSMIflEv7FVI0efPZQIF+LpFMJWsmcCMGC
tDFuT2d1k5zOoU65CrvnilqeJbC5e7SgRgCDOmqYksu/cAqZFc5DyXsDjL4jbbO6
XlkqW1DKS8m2QuO5MI59E793XSlvD+M/XTwE9RsGfCzdI9bWXq+1R7f+RcScCbAM
FL5jeWCb0PI3BuL4QN+6BBXVbH6mx4gelOc53MCt8yaTG27IOZhJxtxdVH8Zgu5l
K1cEWeadlXreOJAP2Bask56+ekFclww0ppjzG1+r6QQauwJvPoAWp/xzqIMlThHU
bfggS2lyRYgMQO/dXfxllTovDLCcbDznpki4Bx8CG52HHuFRNYpqKF1AG8SMG1iH
Gq24JFrflo18f18ZwaqDrLoJ7c7FvAE/b0vFz+ZkT4WD84UnUcuW5s7/9mazrKdv
Y439g0hgz1RJcuWTkUTfFzmqh9t6/uFFKKBlHUpxmuWCRKOTMYCGU/r8HWP1h6Sq
wtvRWM8f5jjZH6xwBf2htAyrGCE6uCsCh2oOQzG/FI16Mv5YV61/N+ptarvR5NlE
DHO6wPfJNjz/eGV00L3CVA8ASV0zDMItg5h9KQPlQVaPSuwPnC1YDd6nq66prvPL
TnWdHf5/1kzcvX5rNSwcPLN1U4SvywqBams9MSNAHj4YzIl2+Da0U+z4ZuHvHzmr
Ju/Ec9FW2OiaupfK5g54C6+CrSXoUrBZ1REQyBotb1j/EWCcoj46X4udHf0m/2E/
NCsP8cFJE+sB0G8OUIQRRwPGy4Q2FdTIPMsTTQB7Vozq4rg385kVkixSWE1Q4Kcr
tuDEqeq9snsoDJUPciKwACnK2h4D48kstohr6T+Y/jSk7pLjsDmbtzB3aY9clnVl
khtkv4WIxcSwsjF9qgJFfFf6MwOkhHm3ZT1Vu5pvsIOlOV4vip2dFddKXW1iiM91
Yw8F3KYxdgNg/WXqNMwD6qvRiW07EmczQaDLltSqJbUoezKVEK1DlAcUsWzyYx0P
itwOTnDGyHXOGv39L2HEEWeDPeoFPmAXQf0wpZ5w7za3JfYzApMbq2xBCsld13zf
qKZIW0N2jRZmbFmBKldL215UOz52yw4PiCeF6ohlqaK98HAmw3xESyp3/ZkEfXjI
X7DxpSb6sXuZ10rQruwVnATNLaAKEvMEMfR0ELd1qj1qnLG6ovZNeVX+0zCTLCkd
Hl6Y1krx3pWTulxbSQRU8vahObJPKAZpYjVETIFeQZ28+SZmn2fyDvfZbe+vmNXD
QT+z/RfyfE833PomLdoex0rXyWQCL9Ui1rU1ob+IZS2T5PK0AVPMp9zm07aKSolK
+BvU5qqVIL7sQ/bDBg3xcjtN7MfoOdiSxOfrsTAjrvW+EIHLEdeIRX7b/Zv5kfjc
TYxDzXGIipgyovkXB9ITBbFh4qa3stxAR9jVaWjcdp2vGAfnF25tXPu5gx7C5JO+
jwQ1kGsyAYCavYDzWrWWokgol8l+jg5/w9P69v1r4AfQN/QatOZDf1XWK4u/MGJy
yCg/KeudV3n+jxrwmpG/Z9NXKeIxaDq+KwLyamrBVptnyqXViDuaoQmwf3XxbPLC
1vU12atRE2QQaYKyzRX2E498XMMU5JwSeVCOItgHOvmJeHELOnfhkVF8k58e8qRa
U891RWh2BZ8lpEvRsuLh3MfRMaigYyhmaeUae0YqSKCLvo0hcn199wWh9xw2z8mu
e/v+aeqh72ae8sfz75hwHH4rZo30YXouPIYWCw0lVuRC7JK9jR0JLi+Rgak0XTW9
O3IxytXSDEEiwfLZnVxO7Tuq1XM1sFJl8himkRaeVP/XthGCTRh0E3udyT6195TD
PTPW8RJbWpCqf1U4jiU9dZbztzwJyMRSSVG4uEl/Qtlo8PN8u3MPWTagG+hjJr99
T9f9haOmImps+DMQTVLXiMnRMCaUE8N1nNlNJXLbRB7vqi3EU2bbMYg7SNFtrnMy
eMYQ0H8LVNf1JJi2dPBIjtCEyybTV8of7D2fIGyHeVW+UONrkkKxvIQrCdotUKCY
CMQU2zvZB4Y36oy4DXewBWgYp0tFR9Ujup+rFhR0Shq0LyGAo5oDfnd7Qa6M19sE
PMZcVMjyJQTeRIka9ofmCVRZp9tdoM1DbpgZWx1etL0dNavPxsbf+IG5hhU3n1Na
dGzLpFi9qrB9Muklw8CVG8BtZWzWUdRNipsSrqts+NtaiLySAH8hw4HGCL4Y+Ctw
dQJ6Lan7Zeia4DGaUcUojKHGqQ5JZn3USe7eBWZQiyYCVZfTwpKd6VzyUoZAsHo9
Z4EZNd8Fg97lahshCuMKjfn99zqE5oa8n+ppamOkOO0so6sUUUab8HtYgHXaQkaC
m/eD7M8WNmVLnLcwYjd8xAAfyV8yqPgF6ykOnc9wKqWEmwTV6VybG3cL6ag7ONuX
GRBjm81i3OUGUrHSCxdOuupU3BOwCkdMJg5RISzpCE76Cf5CQdW2y7CBz+3HI51t
NH7JheLo2Vg/ky90NGP8SSfXVssdgB12OVudgPb80R0lr3QWSohr6AMKpYX4lOYc
EtCDYTwxsBqO/FbUMRcU20vUlU0t6LiC+ZjwiF1LwJt6+7rcvbJge/dZSzqJBzRW
3tF9fEoHSV+ECJoqP4oFEV22dXXHkFMc0J+CL+rW7paNzvwwz6cnV+JicTqgkgMt
vWKdfsJmO0SSL4QySBAXnzcRWtild1wACxyIvxiZ1FG2YUAgCppTeuzGIwHATxOd
4lgCOQ0ahh0RS5BmLUQsRyjucVs/iVI8x5ItPBLw1q1+n04pKZdlub55fqSh0CjX
4mHJ5Ht2IlyItUF1iVsq3GA7V8sF+EjitqAPb/3BQRV6OpjI1Rh9MD93TVGLTYTf
cvcp+JgLoMoMGTJIkNAkw0VPeNZZlzJ5dd+Gcssw5ygPkRNLb6liVbnjDJe83B64
ft3XJWA4VpLaAjK8N5tUN2v59aTqq/MJcCJG0zHApPyhPL/bO9UTYNfDtH97EnIc
jCQ08SAw16QB1/kXNlarEQi+HbUNQ0dxBWwcIW5JByoOW75X9ugyKJJOGZOZMUE3
gUmJzkA4Pu1YuCf1revE9AUxjZLaERDnxJy/lGvrc0qKa7PpnwJdUdhPfiO3ntA5
OtGp8ma8wBF5GHXuBpzeBAYdXrIbl+fcTdvmxSwF1oGYoilWAkdPnonRaVazvCKM
7ilHnwniGBL1zsuM2gV45pB9VJy7NPuEdPvvxvSGwgyIpKspU/EFJlUsQfdRX+Sm
XgaJOohvlM6ljKBfacbQNKOZNV7ciDW4Uv2jW1Oo4qRap8H5Bqx6MDIpRFzZ02GT
ZvxfG9pEwmwUGEvX3yAPc3LLCZQ4N0cNDgkPuKhA96g+zsloWBzWhaDyyJaRgRB6
8/KrO1dhhW4xbGJs8egdKqRtDHJl0OWWGhLf5ilc+P1kVA8WClY+NyTMobpTeO8f
DiRvLAiLDkLKMEym/UIHrt1//IkNs9nsxYt1pSj9NkOagb50Psz0OIUxqfrO1W79
+nYwO/4d/KN9BgLEsjyEjCzLj4ftqonrnltcHAT6hq/qJNXfsf59Zyrna74LKRfR
fs866Bg2/25+upS0SKusRnZ8e6IE9B0yaQWLchwrF0yZYRWRmXzHNfDrgGaQpIf8
s4jc92d9MxAPvMCnP0JIdwcQR+O5IcMnDw2Y0+NU4MTkT+D5wlEqhYoXQytNfp7s
MhySTPz7QnWT+6X9qy/clPH8IXjBKawaC1741HUo3ueBYonabQA2VKLv+HyY5xEh
rc/EdWqr74lA+zGr7YN9GFwJagVq2ZyOgemk0mAZfc17JKty7vgOESKSJ2WV7xFf
JelLGvTHkgP+13kqcelv3ojOh2tcQdhUwSDLivk8JZT58DGCVEBdhSSI/ztIMSXd
JlLITVVH8l+EuwxddsdimTYq3XjUsEFg/uXWQavZ00gnUOv7si4CHLu2bZCJ5bkL
lrdvErsNPwo4BduffiesVudcviAFmC+3EX4931wYk5PmD9npYabLdxBMcjhUv2BJ
g+Hg7FEsAK8oR1biWhQZWSVaB5pBBFsSCaTGiAXzqckwtxkq1cRvMPK6x9s10bHr
O0xVQTXrFiYukICEDrdul+GI3v73K8QOq6sWbz+I5AfNsW7ZgLqEjwzALZn4zleY
ueIsEi+SPh6kAlThUgrjbgLE8bDzV7niOpPshtQDAcu63KftDIW0S/NC7wIHr2l4
VP6zsJX3cPlGrwO0RIwsC6hlK3LWgcY6SC/l8+3508rlBtakxyI5fsWHYSGP9Sw/
2Jp/3hC0JipfEXz1KhfixL4efhZ8WABoTfFEcx60AVvdzHmECEY2ospFlbzrJmSZ
uUPKYUx7aMnf8SwTvTy1qN8l4JqLoTcy07IZQKIDCm0mzrEQaGCB11Tb+xdfF8//
D/ZGKU2nEH5TcGGZe2r7rFlRoV9hvk/tf6vlJ4IVAWwTPMYs+jn2vzve7jmKycFS
o16LLqOzmxTbD7KOG8kqjSs5bc+K+ZCZwqI7dyd5akx2KixNRofn7nLdyEhnhARw
J+Ejyedo8zYNWlrrb55qPKpI5faw/V8KYgWZYB/Frwg6aRtvhtLmLd1i0r6Qnvln
S8RIqar0QigJK0N1I5YYLWMJhgp0DUxzM4DVhs+fpRceRWbpArFkG+k7xA1ihcd4
0etbw8Fi6XyYffQeN5QoQYG7wGiKMbfz+ePyjfWWiqP2l9foOnZs/vB+xszn2mK+
I6a1u4cgSiCXNzEqrGInNzBhjupW+/Pp9SJ08ckXfaBNzfN+55lmVC0ZGNTJwQaf
C8EuIKM0ldwCRTAFQEjdFmxdA1aeqWt577GUVAjFeVPSoA2CTYCv6Oj6EA6Pz2lo
86qShQ/f9mZs+TdoTDYidHn9ID9c17RI6Iu84Ood5LeICMbSsMNIb1R5QSjQe9nD
uYEkirb9w1NIlX0/EFTRaIGDWgYIsgW5kcBCmcNlAokQ3fg6crFC0yF/TqZzz0Q4
Yc0TSVvDbhooMH6NMyAFmJBU2R9ZcadwpW7NNsK3EMR89fkxb4F+cryI5V9JE79r
DvVWY6AzfILHxmTZUAuZQIGJsaPfDmhxWa0/36fGmmf9BkeSGa5ltmj/5zVLBYkK
nChwK27OW94yozuZD6hPTcghNI75b2XlOU0OiaVGKDQYZUnSq97nL2urngzzIuKz
Ro9ixSb91UpJn7qrSGeJ8mHePTMpPfyNwFvvgEHtMFE0rb5yfpAhua+nZ5+xRFP9
jpdjTtjhw4LrraJqpQg/N1XyYXa3oaFbHlCTz+bD/iweFNypnE7tLHzu7fUiXczT
2yFc7hB9jjBSq0o9BOUfj4ExGGmqE09JBVAzh0YJCjesa7Hp07smrtio2ux3KZNm
A+WphYm/rOeTe0GtCn4mhW04lhp0fu4QbMT5vuXrc+gk8iFvlet47Uo19W6Iy1hC
8LMtH8ATMH6+W4kZX6hBN8B+3KiyUTcc6Aoin7950sFEKC6MY0RW6edXVsX6t37n
5kKoh6SOpnyBfzKSKfgZQavphHZ1CiZvL46yUdhOv+/8NAvrM3Vx94dsvYdtz/1R
gd5+d4TCb+kXWInay5/ijYHrkGw2/Zj18yJLkq53i+K1JzO77WHSBzfZU66O6Vkb
pfvCW+hHr5ScL9qFVd9bUDs/kpCgS0spDYX4w7fjPU1127zRg5zB+p74QzG24XXX
ESRClzUGpPnX2Sn8H1HMwAdHlE5/qe9MAcFKQ1NxElnXJjD09YMf1GceiHI8tnAZ
/R3VDzONfJ16J8Ccju7TuQMuuyKAL78GyxI1KbTAPADV1mGI/WuaG0vgegcfP/dR
BPzzRDhFEVhxc+LkPfHK0hCDRsO2nOt5zyBGATSuxhhykVxQhYnYqlK3ZF6iLKb+
K2h6ubbYoMf300K6rD8oH5fGIgNur77EeOt5DQffocShVsZ3B2tWUT92rlM+xy7J
L6aQ+xt42nO78V65y68oR/ZYUt1LAr2ZrAmJ8MyYO5qxuShqBeBcAosQFZCvqDga
FH72VUoQf+4Y8IdzFRfA6MKCl2leXStKsoVu6lenTnvBvoY3owzdTnHoSkkzdXK9
F/xhkdAlMivm+7fOq9ZBXDZmo5FXs2kKW+ICYrS2Tb1VU5G0jlj/WUHdy0Xp0Ee6
RgAm+C9auefQXFEmhyQciWiPdHGXS05Y2LBDyiyN9wfuqeuh6iDOzLWTeHr332lQ
mY+6jwqP8KcMB5fpgQVWSeHuqBqzEtj+ebVBbFHjrhuT4tk2caxW7/cv6ddV0Hob
+vwr9vrAAjQubAskqKeE3sq91Gt6skbc5zQjFHcv9bymoaq6eR64jXpOhebBogfp
WO9YcA9AYRXZFp5eExyi7Q5+xAdoO5btzZHOxpPSAMAahzVAeaEgbSAsieKQq7hn
fWIOEmrbqYdqXk55mJH7PXoLawpSzItdCWwVe1L5NMHe1XcL12It/CZItyWujCSJ
23aTpTFA5GkKN57uaL/DAtNWwCQenHlVz3DXbSqUX8PLzw7JqbUuk/z/ScjMLZif
tyTRJtuvPA4iP0w7ked4OZl6s7tIQho3hjtDO+kvlgsm+pA7O6/yOC1oP+PNGctn
oE5vRW6UBd1v7fH8yxjOfC4SwcAA4OezTQ37IFSG5PN5KFrUbKh1pnnSDrVTW2ku
7RQCXuBnb///II7J97kqWTtob/d7lSwkw8AF6zpZdmJwtZLEpwWTTCeLsFtzO52r
M78w0oirRqawtM6pove612wcUzu9eawFcRieY6gsjwtlCiTHHVAu4qXVOnSInLOq
j1Yr1xScTkL+9Qzjyq+aXe2SRy5m8R+cicSOkeW1ZI5uxuJewQak6eMeNpWDWuBj
80Y4RxBV7FTWP6H/2tXlGLh3zxncg/BUA9MsHMV0VmjM22YT3ku3tzdPLgf7x0r8
9Ts/N4Q/4U0vXuY4S/2L3QJtGQk0WZqqEs9/whF5Jn4VOnjv51tIvxsirLna/0Mu
J50ziALQg0GnRzHYblkf9xjAmGO40Jwu0DePfFRma7n6IeEiOQCa9e3+SSCziAA0
Koel3ZK6w5yXTc4xtTfTGYwsd3M6MhZUTxo6xS84VQKhZ2wh5w0ARcERgosfaTLS
sH61KqXLHevmEDi0y30GVkRf6Mw9VEvCEhO8YuLGIWyIk+1JHNMkFEMVrqMzV0/3
OoL9aLWfXVeji4MKo+2AD7e2BuYPz3Mm0dGrKqIdMQSfpAp4BM9rujg7BBm8l/Hv
5CFEQ5I1PqeO4owzAou9WcTKPxpaaMN1g611JYroCsOJ0B87lOYMoWpg8uQNf0iX
0NBiob1uOj+4jwAPu8RNhGhlsh9dbz6giHduohPXLXvgAz4Qei7cUiJMDg9CR98v
WQG2ZtpUrEb0MXyw2fzTDnxkZ8HffSP/KF6twaFQaj0zBf0ulDSgii3yCRJWJnOa
43prH3Evk916BgTscFlAOB+pMGknixISBwX2grxAVuQ7F5xhD1rGLLp4t22cX9bX
B1W1vfPpsUtn4SRSGfKLRIjIYymOsoe/29dgs4GkO7rNy9Sw+Erbu+y53dAt8unZ
tdn944mEVc4OyWUZUJGvobDbapMFAlab80sOGi2VadFNZNSUamButvKmAON50PS3
TFP7gEcbwnokzdrpFHlIJrzBorqf7kDl9vo2rCt+ym6QeaEG5oMzDp5ZPHGNfEjE
HJkmqAjiQmuwXITT7KCzqYAyYzdG8TzkXsOtCNXVWIZ27Nzn53GMyjilsZ/w5c6J
s64/MYgo/rTbHp3aX2AH68T7xd3jyUCLfkYCMc4RjqPE6D3f+kYTVGsWiFw9ofYb
RJQFKI7pfS0mtuTC++gpEubRZBm7Xip4dT/r7sJ26KsyMcVpNAwT6zkMtnj1U2Zh
9cUatTYb2Cx3gY01IEaBi/8nOCN8hF5Jeq36OBXRDVSu3BsgrduJUPvjcHXWDJd/
nXQ3BOPtK67jV6/QwBKiZ3ifms7mCeiFu4ClCgocSwKNQxWI0R3HCa5SJtNyv4DC
4i3Vb57eYEQ8KYngxDIL637XZcHysaPKJmWOLbsR2PIBHmR9Or7/UH6PJeyYG4CU
VVUL1fh4oyqhV67QTYD2GcPmXTOG+sXf/jsM5qcxbitjLpiH0AVjKIsZCyAPFmIf
mC4sovF7XoNGCUuy0UHAK8Dt+m0wJGhTOUn3EpY3vJw3SGUxTGIIjcwThhgxZoUs
4iwxFYJNrSYw09EOnUmrof06fs2uB8nbhY5CbCd1/XkwH1sHx02JUSWRUV0CEwIr
s5jvbniiKnGkBfZ4kCqVQvQ6SO5T+lVBtC3abTRrmwTffgZD4Qs4uIBKtJ2uaAOC
BXMq6bKCYWWcmk4TMKNPmFtBkLUUn5bgNcB0FP+ic+8yQCuDMCUXQTHYKg6wD0tu
IPvbD5e+DSPEPG6Te3MDnxRB7qwQSmlUUiY9sekQCNBD6sC7WX0smcDxVFHGbAHh
C0eRZV/QtwGLcnGNB6uFDIuK6dgoCb368xYNDb4KeAeB0daMZxhyoTkGSEJqzPy/
WVHQdQ0PvP2mpLLCevgHGElvo+DlRzJCYBB3ZcK834VNoXhlJQFgRhKhNtyCVNXA
PW7LQRqiCsgPjSdQy7aJbazbeR4hTZ2Eo9dOyLE8/OxPQtCzcZyjPVZMguvvzMEn
RV3sBYLRBDuZSsMoDMMrgZNM9zxJU+as+0ntpWriP8dob6hG9Yk2R8r3Jha+/IhQ
w0Z6z84J6ANgnHkiF9u/aVeMPJIEPGe8XHt/2z69UoEgmZcSW9ioDQ+V8Zh4BuRK
y1/4A3nE4QxbkHes+8TJAUozYtJVj5XIVIZFC0r0eD/pkP2NXEcOQykAvsBw6S6j
Tj5gXhTSneFE16bgFy8FEhc9l0S220KKBfFYca1bHclnh8ZmKd+RITauHT39gVy1
VbRRAL7S2wRfASgIjiCkKl4qHxko8FaekqxkNS5mWVgdYuhLIJYDj0Xk/Cna0VUY
xDD9oQ44imHKHlJ40Tv/0rFBAtZ1mCLwZqaawICfuUKlix9033hqO8Q2nUSseTpd
5OtwNd4lQ6jDuObIc1cI9JEzn1zoebmsQ52G+pgiTAWUwiV9yqRogcyeamWrFNaS
oKmi02MtGb/wzJ7pH7sgM+pTG3qTW4aAUfHwp7WEkP0ZfEpxU4a7mKtzd7ZaxjF0
joCHRGex+4FDPt7+/AOOUsl969MGwH0b2pM1EffgsNdf/2piJ/R8o2ADyXuCldVz
gj6862njg0X+Fhy7u7I5pX4v3SMZNTDHB9Sti+OS8VWJMyGHNuDA2j9S3Ru3KH25
KJ6sXf4ILfAeS/5wFicyavbJsZqCXtmOjeTzY9FG94kZaTKca8lowuIKANpNzQKx
f12vCXfl2sGCWvJgQfGn9FVgg5w4egNXjb0TXFtUkDcCXtVYws4fLAZywe3/iPp3
+C+lCUBYtkxRBnCtgkx363RDu+Pv79zitr164ug7BBtNoi4ok6TpHQo1ZiUcvDTu
gPyZpa0HRP4PBVyDhKB7NuHzXiwkZstNsjpETh9EIZCwN/jXc7XbsrMTrc/EcpoK
FRGtv5bqXMXJ3keZkTAzusb+lK+hP/jyzhuvi4oMZlTJoTGDQ40O/nKUvOcxc0aj
+VaqghBAFXqUrgDMHxADl0MAQf51K+yfUJYWOqCKdE1z5LvVdNW5gh4WC1TFG77d
Hkhb9xJ3pG1QZEYdC/MXaY2Q2DnMKVJPn5nxjfGcnPoNWjN3KWug9kNfA9GyNFeJ
KnDmnIWZpRMEnzrqimCalCWhqMp5bduM5XpwSxmqmbckAzGb2QjfgyJu2tHX9RHf
Sngzf6M3BzjtseDiGL2m3anAJ9xgUOvNt1TCylz2lQF6fYSZrQk8cCMPjcsgRUH7
4VIad9sGhAkZrm5vNBljmZadhSfgeYo0xF31N0R/ZtUhhWwrCkP1ZbXukMQiR6FJ
FqSde3nD4ifUyizATzXDjbLvdOpHlbOrOOf3WaQ34BMslfE04aLnWFnuVACSl/l/
pJ9WbQfV5OYljYHkh4Lyj1jyNY24A2viiM3rQ88m/P7HBStr607mL99QN2sZDHkQ
9iNv5bqMhs3AuzJHKR80cnGaeMqYzmd5oYxOSAEKvh2DjNVT1JkfY0QYz7kD+BtW
EDPCLYwGABJS1RNkgoeUwlAkvzJRz6NDWepyhw7UNfxDlF4SCB/NlKGfBBajDMRj
0+ONURhFomi7R3PwS3xNX+ORMwGzwWBcVTodQ2URGVYY3JpgY78S3B6mRcHeV7Hb
5bPzQOXojCIVN6ZtVmj5f6vNsXPveQNZY3TYbrAwuvivjRE6mLn5lDeRWZgRMXac
E0ZQ5Hy47uoJh+KceZL8ICqdzaSNEooNdTluYCr5XAzv/qZ0wQKK0lLCY4oXVRPw
EY9JBa94K36z9l2I1hZZuWP5AgrDmSoN+36O2r3ZDZ7Sd9coI8k/42GHzo37Rb2E
IxK+WBB8ULx+h1wPB+YSbydYAl/Eb6HLpZNavQR0506LfbYCsgYzXVHYdd4c0BQ2
6PfmCPDI1R95tewp5ArNG+lm2HYKxPvx6mSpxgbzIch0uQXSv1MMgQHfp/G1oK9L
0oVpUdijFC4vCHxDGjYvn5np/ICURvjz1CLBYQqlwB7+Ib8ioAQlgAmRqdQvm/Kd
OETY0U6jvIAxx7k2J6QuAUAz5JSEE+LpUh6+5u5LJSXsgImVxCCQ3j9tFVJraqGC
GXqMS2jMNsBwgea+DX5FxvyYS6i2ztrVvW/kDicQh9uj2hZOZ1dnbuuUvcqW2SHu
R4enekmqQCJzTFyq2KuZjW4YnIwMsjxcl5VL31SH5E9tcIm0TM58xP1mN6PixhIj
N7GboScYmCGpztd+WfR2YWQOryy7cYU0LmNQwnDgdhdWC/Qe3vslLulToWk2AC4m
aDOra7t9K8v/11tOIounFEqkodMMPFZGxTIvHmwjLXCSn4tkiwiozUxl94nr3Tti
+1ULMPbHmYUTSP7eQPtcKzPUyr1/7YYnU2GvhysizH71cvBxA5HsyZUl3BG1aOd4
1ss3OOmNea6+wLcNCs2bChWXRL6tNdZzTW0o58BeRNH/LPaYvXkj7lPLpZMSE+UY
5FCMeT8OGV5BhGaoj4ngeYLwUIF2QfOj8lMlyYBAAUGQ8FO4/MjIBx2gezAhNvRP
X/haImD9dkvkknarglBK5+N6RHsfahyDdiIeHtYMRTktf2jMnSOOFtOnebbn6iLY
HW8NmA6CDaRE4k6vevXEsN9WOPLgVFAP/wkC5UnN4+rxbYrzWbzure11sKuJqBNY
CBU3u5OCA3jp2RT3BI3ozwY1JHFJgug+ywcS/4fyfpCU+YzdHYcq4PZbATpSaiVp
V9lLBzUI9juQ3eI2AkKmJ6neuSxEdIrhs7F8idvWzsEP1cNKAEfly4RGfr3yRTJV
ISJT3VUZ4QeZBLtQwBc2XzW7LzoAVmobpW8NjgVkVBtq1n5R40AaDz1/T1hQnTwm
ZvPg5n+hu6CQoEWHHXreEapXLqfEXZVstDkwcgEQ+6iGyBMAH4Uv9qQKaxxR3riK
uE7JEd5LvreAI7MQ5NgD0PTGFiTI/476cBtSIykmVHjtT9LSRKP3eyc+usKyDd/d
Q5SdUePj/PaQ5oGmI976SnFSyQa8CkbaUTEWdsN3t2YZJWlpznjBcs9mfpZUr3iG
+2C5FqRCtttQsyUVP7VUqO0niFFmUeCjaknsSXDi9YGZwUCL/XDKY8NZekxOmp00
OH1FpMAG1tPR7eXyY82o6PDJ3OO95DDiz3B/mpVCF6PqC0AVRG6ISOPnLQ7xEify
4VAMAn6n3l6oyxounfmr8bERnCTg6PgvimazEIlUxwRJ3hEd29OgQHXLmfaLmxiq
uyQ+KtJ6TB+5+hu48v/B+rklEUp8Cxy352ur3safKla4IqPICqeHnUTH0tpGMQNL
MxH/Xn/e+VaIbU18S0prOYRodVVYCEL+GB5pwx2jrXltvthmfqRJhlOW/Qa4IMzk
qVd2Fx8xzzD0UYQgtpJ1HHu4nbS50AjRuF63ELNnGoxzudypwnINKlGhOp88lAdY
Lu+lyi/rjMM8ZD9V1PXliFdnf8j4VuTHAaFQwWyD7AfeJuQ1uvyq+LAcCoznNGNK
juxkqcQRbbI9/QXiCet5Vy53pleUvUvIRW+WCqU9m2NKUcTor/4+jBkzVQq3OBDc
EY1pN2WstsdWy1lrFZMJn3c657Iv+89ZIrFKxtPuJJjUwBJd7oBPgqH/tzuZaV2t
K33Vl1m5rGQHOY5uLoeoRns+KPLZFwJlQGIP6eNXlYY2qms1Gw2qpLcTeHrwHil+
KnS+T0aSQ5MQ0yA+y+xFcpFea5LpRBh56nNpwc4p3mLfRYkMfEDRZLE9b2qfDsqO
LGIj9LUYxX3Zn7E9ec2df5OseYtZhqvjDKC6J7mImQY+m6ePYQPYfeU+hou4/KqQ
s4AmOvfdXSFQUlQWUE9odTnkYZEl0xrVRj1ypRIHbGV+nU2s7qzUeyL3lMXhvZap
2tuu88EL4GWP3HU+CMMyfBBAvVSx60LcGlwQgAImnlEEbnDbW56DELmMvU0Glfs0
mzXgQwTBXJh4HsDi7zjg0Gm304txMdO7vvWWq/tJ0GX3SF3BxnhDIWEREPblois1
Ob9Yb/xWPtMUhC5aJiCt0MYide7uqMIPaQ+3A6CBJ1KmukbLxN22HlWLLNtYmzIa
yGCB04h7UFIAW7YT/aeAMsbmmdLhyx6pqkCOTQzojQFZp85VNT7NL+Q85rZ6Dgfk
ztCIzUMbe6uq3Id91OfpaeZXdzbK0p2el+XGTbJdPnHEeOY4g1IP3BqGeIj02t5R
rk/62WNqCdRN+U2E08+TnKoMVcYJ7nLjk8cy2gPT2XBAoJLQj6jEoLEBRZ055VCc
NdySKfeDzxBqif425Efvc4o+F3haiHTxq6KKD2kN+CzDan4+BdF3sBUEVaO4xbLr
YJiOOUQOrjbqbq/4b48jKsu3iVL+fexEldr82o5/VfL3AVhrHwTX8wLoTiopbQbf
75rDYFuH6fXJUSmfR7dkAIuAt4eWspVWGOasDajosJo8N4XMhskt4Lo8qWvayliN
FgTE+YiJDKHXzH4yjFuKRMlLabbQ0Ge85UT1AEsWOPaVDV2eQye8kmXSno24Ci2C
3/LLY50IrehKjkeFgdl+TeW+iyKScR/vbJZmnRAL1EFuYSvgDzeqfQfkNmNj1V35
lLijKNPQY+K+Vi0CcRdUY6UMyfX7TN0HhkZDcMs2OdYHmQ0Afp3eiQ8M11yHN1Um
aXUNBUl/e4Ot/HJ9fnayk/uYW0r61ITiYiOcSswh4OfuQTpkubhcSEco6V+cjfig
R3aRcDW1nWj6DIq/TOIqQOqcYh0lpOmYZVnmxy5tdjU+jASc4GpSLQULSKkIIFQj
oIDmfrg15WHyY5HEguCTHc69QNJQZZA4SgLgfW8hkgzIJRWONlDTCoBkNlpSQnWI
nls6rW8T2uXQto6Bk3kIC8HpeDQ/KONNs5w8BNyHVamn77h2AxhuKG3AdVjkOI7c
NMeNhpUpZqacwbqiPKtjsaTm0UkQRm8INIAW/v8aiCklre+MWmoGyA9M+JioC16T
ZAZeU6y/hlKsLgzD4YnSwc6yoruKuw6NhrHb41E7tlcqqp7wru79LC5Tmyuf5zZu
panlLr1WgKPSN/lWW9zM++AeiMdhCbAce1twBRRKg14g6pmFjdgP3IqwPlkQDNUU
nIJux4e5/GV+e15QK8lw5sE4R8XBiALCK6hP9CJ0Zp2onKCI/zSySnwqFCWHDUFo
koZqCL8+R6+GX10S30RPrUmzueYnj04nwcJiOYiZ4uOCUmNZrCqn4Wx1oMrtzGxz
hCJC+wluFPSNFFmAp5um5g4/d5IAXbxG5dZ7XCdvwQl+0rhoVmuts6kIg2D6QSe6
DQr5XnykZJQRvgeWY6FMiKcbh/sSarE9bogiHUJA4GKiBoUadcq1m2p9j7kPLc0E
cWPtZfOPdZzvOPQl+T86qxeRFAGYN1hen1ZWkyGGBMfcLAmv0wO7uTP3x9fuciCJ
u5NqaKONF92ppFy4Geaaf7JU7UuwD4kvEIMia4l+Y0llRPgxd5MhAkMLhNIHa/7t
emg6AWa6clMB0ZCgf3PwPO57GYM69A+f9SaKmBgrqahMkc7/mrd1JUs+2dXiGoug
9ETGZhPxozLjTYY5nASNLOwbDwHDndznHSBBhG+UkxfAmKtaH13yacQcrL6pHHAx
krd0JdokjX32dedUfyP+Av/uW4MmQTJwxObJpSZcP2gRMVm4dyJEEZ+DImsa612k
E3nSMbHRFrSNKRHxZVj/A302RdY52CvzxxtTF15w/8sYZibR49WcoVko6e4+v6lc
T5BOTcdUkfx1lTfe/fvE8PUDNvd06/qn5nWV6oQZeflEg9/ZkUPk8udM5ECYLUsL
q7kqfvZ/e7GuKGCKEIqCrMi66TbpgxHBSfXS4HCAfUV11qkIzFFmEL6wFPXL3WYn
fcLSuLWFhnhJVzmtwnPqct/RShCKwtyU9orw+HUnXOUiAn9l3YZBueQhKfExd0bB
Fr+Vf7qF5NJlwgEsMeh3vo4kG4sx4OyQNP85nbRLj+Z4peKJirrpyzitMIo4LMhl
jNTZnq5R8SlZOclKCtEXXfEFggfvEqSnpfHOqssrvMyo7aI/S2yAFKX5IExXx5bQ
i23lIYXELeWEmcTm6eUBGzwRCjhr3zvA5CU3HjDLgKcXdzLi0rL8sD2lzCZX808t
X2mkTV1N0wNYBhxYaQwOVC9T204dQwSxEte4AqJgTRCvjywLy5J04wHK311dbn68
x+Z+tC9OcrYk/V3CI+WrAHu51tNPHqGXZG8dRIUws8NiIAUFeotogpQ9ojGoEWuV
4F6C2z6qhGSYqR/0DcGdU4oLUDbHBG+g2YF/rtHZ/Fc2hMA1qJbVaSePi3vIXnUo
J4KsPjky+H2pUBbAhUpUz0VVRWPTCaOIfTHCqJVG9lfbmdDaVj6OktYI8DRKo2FN
W8LAilSnWr4Bb5DpwDVwen9t3TYU7e8LL/9TWrhkO+7nsIT7v98PCm5bGtzWUuYl
02gMlxdSmuS/nhNtzYkIuoK9Ut2NcwD8IG3JQs/EYp7hWoAMhSnQE3eHm4MRMA7X
xiP/qa5LLvoY/T4OitOH8/2AMnMvH523aqyBBffNLq3P0LMvxE1zF6qJpWF0uBqw
tgQqdEd+2/rEsQPK3OebgHybQ/w1h+i+ObNLr/W2TF+xkNQ8NcmhsDx7P0f5I1bk
seFZ62rafq3W/LuSj+UiQYBQn4/FJKZkDDwGt7IzNNO19j9nGFinFAJGAEoU4sOC
xr8TtVZ+5tLBRS65EknBuYcJIELOFfQC0jUWYOgbUizLLR+Oix38O7Eoy43nb8fv
ShA6Jb24SG7EBenmK2XOnQUduWHoHpQsv0M/SAd1gZ+wcpdC6weJtb59TrQqIM2m
8l4wH0gGhGNaYK9Dl/YcMNd9CHD78jJZI8jRWZsBQhMhNHLKrhsG9PtYtVyGOJBi
i7VQff4c5AZnrsGCZM1B215wwQ0TpUE/r8anb3owXp6JTJLOZYQLPXY0mEr3r7x6
9JwnQPwWKqk6mq88C6w2RDlg+EtsNNGaHNIeNoNnR8J+l1w9pQ5So5PzuWqXr0IU
IZ0ObbicDMJnCwqAd6gjgcn6AqH8ZK1gG2L2U6vhzUWaVdFmnatVnIRJ5H6hJaEQ
5doLCXuoa8iGlGP/SkwJ9DU5b6is7zrnLFYfolaheYc8QPjnrnSICPbTncz9EdDP
4tZYXtA1Z+ZNSVnFTPVl+TuRDEho64BK1HzISvNjJOYkEARuYFIZntr0vJQVylRb
T3WR7gQ7bDODrFPqf6B99PPTzHyPeJQMCinkzHc0pxbRh4qR+IJ37jR0eoM8abZG
/6oePsQw5Bw97AsHDGXsiCAtztSAwVfmeXYAooBzRO849S78fK6d4UjkcVd4LHA/
9o3xU5kp8Bq2fg/tsYZSqH62Fud5T5mhcwexUKn6rg9ajRwthDZs0Qtj/ZO3Wtb2
jTEaoGymUICuPrtDqCA1YefEFQZx81JHD3UisVVJStld5GwmiJkj4qXt5FYZYgHK
KrC7rdWqhcNCTuDBPOI/9cvqm+4vTGgCD8HtJ6Jf/xCVe55zOrV+8atRDNEQL/rv
BPCJuACopgfo0EtJpZwHkLTnSKWIw3sOBHAfGDyQz8hQISEjxDHjXycvYf6ri0jn
aKfA/9Ufwe8OHypNYK++EtmnEY4CwXYiicXcpkx5fskBExNdEdfeSNX0n3kITL5c
ChNvLC3/pKRLEuKH2Hbe5JpQMv/DlMV/KyX6D/RlvSfTz/XdX36U+XnDy82UlqIF
OebzHFj2X3Y7FwWbJsl/s25e3FwHMRFN4V0ZXXuN1eiUJx2Cp2kdw53/hEGARkrp
Iu+LFm/bmnUs1BSXvjH7Q7wGcs3HVO2wsjoczhPTSAs4dCH3XNtvZZ5lsTK6jItO
WsYD6wQdBCWVqu4+tsr5M97KAftSFRQLK9kESfrshxYazeS9ycw3Z/mio7aPzP0j
76vwD9cDSNensManlVLmDNJg6CNICbDf8RAczqaartiisga9PB9DHNCVYAi+GXCd
JPaxempbb2sqbLmKTO50pOyToxj0AuKvzsaU2p6GDPmkAYIit0/CIntLRzSPZ7YU
VwEkkC2+pXmSMsxVAg7HODe/C1LRuJn2H/ppbqLGrlzS2ES84+anZWoE6fkPlC/q
hZvfvkx5ttWTtqe/86aKWfUML6lPcKGchF93FGUs6/MtKsqdq4pSIwX4zn81aH2P
My3hzwvSU7G5CYD3+Rl9t6yuU3k+8cBBkSbveSrvs3ts6z56y31fDEFomQwz752n
YYfR+qVgSFD4vrOyVO4J8GpDWPzIsF9IHESmtFldoS2ywjQ/O6SloiiK6cMIRwIa
DNXxNRYKiU9PodH5T057AP70AfFIvReLOitoxetV/2nsHPUr5yPNEgl1Z3UvFyOh
G+XJayZRsWL5xjDa7J6BoBZSabstNRascfeJOBlGUDuqHFiLn3XwPCfKYPZ5kLkC
o6bYgFvLwrFWwvi9x3xynTvW00ThxzQILrsGlyjAGt9j0G3NSlPkooVlXm2gp5js
+mwySYFo1kfwVEBW6oiwGxYtP4KYsAxTHpODAmNcX0kT5zYXjC6QQ2y90vT+6SEK
ZDJ7/7FrMOh3imUqddeDQRE/RloKb1azHQrbzrBuYbxFCdvXj0TVwZ7lOuhpuAQB
m0GUrxb+S2fCDYZfadJwsWDgryH+u2wz9HLJXm9PCp4ZlB+rMSN84u5ZqR439kLp
qD2L2rhQ7HUqcSQsIGaLREHUY7Qvdnsy1SX/Cnt2U6ZGlHw0zMvDabrHLocCHuqs
DBf5KdI9+mbflu5rE6qzcMp79IE3XwmQhSc4RaR1Je1ziwrqQ0wzboVQQNT4YIQf
/GHQKO0JCM4EIzRSO0hLhyo8iPLtx2mn6An2qFC0XOpA25lHKIwehvjEQUssV+OE
DTJIvfFa86GTVxLbrxkeB57SQrvKK42283FbvFLqW5AphO5psh4GGxi5nNyuigXM
DwFhNgkNoZLBxdHXzxeyjiaWEheBI+GiNH8fin0xbww/uz3qUraHNzcHQbwf3KKq
oHIumkSCRe9csP+Df1eWbmB7DoNp7QVU+z76p1xFGbRNB3peLv1IG+SQzumg4Ii/
ZIs2oeS0udp9uTIaEfzYYnLW3fV6PQxiY9QUF8rs+qlNjnILkyEF013xBfWoEDA4
L2ctSO4+1n8U9jzuT2FDEt7cqE536lvh+EtspKLI5a7xH3aqJPmLEYz/xtEW3gIf
sDehjqhZIUAbtOw6An2gGwRUbQBHPFOkut4r1t3d29OP2exrN58GwCl/HQNz0U4z
UdWFb04BCXRmHMFMvjzKIc2I9x9mpq8V0h1xVzt345JnZ2lGmqESOwnFbkeeaDk7
KXvGlVC3o1Y8rBNTJv5wNV2MH9tzPglIYKeQJM4F1jakhdrwr4reZF/4Al+/mt5j
AtkJwHYUvPC2myzOjyJAz8SGYrNzi8/SdVF9q8Avk0VNrTlNkURaSigHXy7MjtTj
kSXcA5Ub4FSH/FVjpDAfuAwuoka2pMPSHaMbPm+a4WvsSzAQ5IudMzWVLksboOsP
C1TkU/sqUQ9vDyQqdGeHwkbf+dYljJftwMHphWj4UG+YrSxXWXN/pgfNNKIb3qUw
iE+hhB4WroWuMXkcagNeKCYzwaU4X6PVDzV3TbXrCRT5j1Flu6XlA7hF58OH9q+p
fxZFibTnZFs/6DvAcCY2HD0DpG7b0GHSz6S3ScUAFAkihLuHY0DdOxSFg7j8Ip/8
I4ttkAkTgyNTq26izjFFsD4PPTsaU86t+3P+QP3wWGU2n1GWt/olVDDp0+VYFVuO
YXI1TIhmDhC0UVWjmTn2yRMNYHt0r0mLUeWMh9oSolSSCfsHYPkLQkcckSFV7J3W
Rsh4/pK8A2j7bRnmP25LwfY3vGewtspB7Yhv9E1/nz0Fg+QAwtCebyUvSOIZugE3
/rCCUmybdQWxrkT8l6SzXVCUocJptMPk5y/wSrHL1s8SOVtgDlkQhvrkey3ds38l
v2DpWGe4hYcheguH6WW+dnq2KRORdZ9jHC6AVkcfc8ZNQD24wkJaqY9/9Ew2cdRV
GGAsMFlkq/6pnvpEY9P2tbH/6NGPvaKt1hdtdNwLHNGYzukiNLOxdj1gxKMooLeW
/RbbJ+rPFyhDs7ltailR/3MMq29Sl/enEQQh/TkSuGiy1hYyUauOa74bbqof+DkS
xwcjvKstgQeusVO7vGGwo/j/CREoyqt++3VuwdA/I+Uj0beaXtKL3+DzZUOE1uHz
1W/J92EVg4aXk0nZ92q6Hu70iOks6UI14v7SF4qdEapEODNfBFdcYpAtLQoGNybs
RQ5EzetgjjDI/qc6RLtHmS6PgX3EbXRYucvxQG9QK8VcyPPPo0ya62ukjMVvhTMi
NbiH75ZRXwM95+GNOs3Ps5zzW8GTnadpS/gf3O4INzZB8HTZVwsf9ukwTirdwyYw
cKgkGewnb52nW5CZw0A8jI08d11EG5x40nBPOrB/VriTGk3Sg7eZKFAyNwBOSbT1
GHKWeweqFXatL/ixSsGQ7byKLPNCdh58J3RcciZpekbZmU12lLlwnF9IzfCJKRAC
Fqry6l/ljhWoBdRfYlsBuOJzSO8Mysf/m8TwU5knh/eKn2l3OJXVD0oQymzmMoY6
1bsU2TJVjmqUL/49zI6Ca9ZuZH1wf5Fko7qf3H50XovufEr8r2xwcLXyD2tDrsaZ
Cb7npQjh3+ZZn+IQvVyuaF7LM5rsxUCMs9pCjws/d6vmD2v6xyNjNQamRI0odiKh
vcocXGTHSV5jIvGzXmafLO/Y1tvzz1Q042lTVJfRUPAUXxKLp09kRreAew7xcW6h
oTSI46pVDue5n/HjvhM7OV4NWdwohM5esucGgmro6ScoqPKh/NgSuaSyoQh3UFxm
BUkW5u9tZhxOXrtZBx+whc5ir3R1Axq06gQj52tSzEzdd1Z2hPVVDFjyCqhVqXQm
Sn+26Jlzp7szrErvkQtAQ2I0Y6TJHqq7IGtntwQqEn0PtNYaQ80C3ZgbPXIekLXm
ldmcLr2dz1nM7lUcYhTpdHVxQSC67Om8EK93Nkqvut1+lTh+U+erZtxtk5QUiwW6
ZwBOl5ZxV5QwXsctnykh6ENDoebnkpzm2+SgAlAf88KAm4x/w9/xjTCy87bDyHdZ
HVcTrC+b7ZBC+OHS6tRFUG/z3F9jvgzgko9q9v7rNBLRa4uYpWnc4+uVdw9j6M3M
YEGo4Eby8OYLnoiErkMxa9S8SGX2QlLvAQs/kfBDq7NBrTj2fRi0IM3Z+yYwQQbu
ColLx4MLLA5q6R/d3efRTPUNHECrIEpgeCPrTMG5jVEao66HVghVss6bpaNkOpeL
DynteEUyfQ+c4TmghHOI4MYcQNO2gykym1gseQX6sZIjqLIHOM2GK00CmpZt8Z7f
8KDZElkSqb8Rey+lMBek0U1BecnXAz4UKkxejLGZ/jjTCZR6Dulrlg+R7fUIzBWd
pwl5e+NU/pJrRWOhKnaL4REhPw4+k/6Gl0i8jW5+FicsERFwj20A6tqsM2zFx6tt
dZSXAEgZQljA6MdgSYixIenriBOfqqxnUVZ65Hca3qeElGpDagfTYZmY/gduoSHA
1a1u6rObc5PgYpbW4XjkeW5y11EohXX2GDFHOtwmrTaVa1vIBwvMg0pi8gxSAt6x
/IQIFKBD2oDvUcpI//VaZ0CBDUsKZCSR37dZpI+FC1HCJECvOAyVQryS1ubUvHmu
bp27QUO/6TUMyLIgrZJw+T3Mjq+17QzaaQ27J0JYSqIJgPMdYqXIyvaf4/N/lDId
1WrcGEN1PPYKg0nolW/Mmiw2jEYd/GloWATpI4zMW3/EseI18Ye9Ix68ah3+NPp6
Rj4XD4cDZQFo8K/qfYTBxtTQnEmbMSfnb4XF06hZ5O8EuXTHSQpNB0GEGxfW+yYK
XRCK/xqd7yEviX7C2au5B2WrIHmxY1CeMscwzl/KXNIXQY2aPX2zz+zyrQfZ/zWD
E0v+lXN00/5Zi15lgrSRwYxLLwwr1q808sMCXTvF+8MLeBIsW48mcdDtfnEZ3wIb
DN3rukZDbwggfO+3dbzLKwgNhSpRjIRaayidPFbDfiD7Xwt5a9PRebnp+52EO8Az
+HKlHCtdu1xzTvHzhvw+BZJu4ELXazVIzkGCA9yGVaMYyBDdyYn22ORS8FAHUPjB
tlYHSRl4qxfptQiwcw6i6eVd5NotlQv5pg/xgcvyidIqyL/cRgX3wtPRNrCUf9d/
agug3JBXIIortYantuoVdXqN0xhLXbJzcunXsvjjs+VWC3pjJd49t4dL0Gi8+PC9
ypQzFAlakobQVcTUTv2mAwx3/uyXB2LT0KhTJClT82YJvGKllj7gN0Z9aaGUiIHD
tpgQOqq9HhgELRyOgjNWcD89pdKI8jg+fRNL9Cwmua9DQzvqAyH5yjYkn/zH4Yt8
QJgEvjZ/ZIqPVW+cMPpLscoCt2HBheitsGGSQB5pyve4hSSaXZ0UDZkEXdE4GXuT
SFqz5nAkS9hKQCbfXLDmzOnIgkTHpj+WS7QE3IDKA+UiDvJ7GoHKzSw3QkWzgH0c
LBPKUrD5i08tCNQT8u6V014JJ3EqyiUOKd2snj7a0PF3JNyL/dtXoSQjX3Ajl2hh
909fh1Yw1fBslGAiFh7HnxAVK6Vlbw+U98zk2DgEQwVjXtficK1UI1EFAlotrxlD
tyMmgIbTbkaNuZhlNmEUaZkPgpTf2yBvw1uGlvGqi8GpnjhiykY+tuHQO8AOmAQq
AvQ4I0D6mbkyN+50ULV+oOvtRqh8Ib6wfTAjcDZ3q8GfCk9mD1FySsB5/7ZJJ5Wo
3PzwX5e5jVJAOsWCHikb2hKCiPHjC32CqrX8FkU6VuQ/+yU72+sHx20sVC9HO6/v
PzkM4YoooN4uqcNNnfCFZ3llYTyI/rn/hzjUSE1RrA5MNKGVmn0ZzHNI/0XZ9byL
6b7B5c5MVg/Wymku7dfzwsMTnEnaOeaU/3qsJ5SaIIbCHCE9bfVlJVAbi1SuexDm
86OK0cgtIoNaFNVfvX0mD3zTg4jdZtdCrk5mME8+c02qLl8GB2EROD5ZKGR8UVcK
imGBdARj8YeWvN5+NZ3MZHs8NMVStsDlCNnU2F5HG4xz1SkrO5g+70/AIalnUbj3
2uqi5Wpl1WYZhuDyITPsQgsaLs3/Lf6I9vBFKXsocN9VD52b76dqhRlNeSl3+deo
3ehY9ABelBbEssSDF8UQRLwgGYSK086WqlZFeRczWceE7cPRA3R/zbROcZkzPgGu
nPqHLVLho8cGhf4ir2V0zpt6ASpiKVACoxRwV9fBwSTjEM7Tm17SasUZnKxxBEu+
UKWP78eNVDQxDNyQ0JVNjvM+75X+z4g4l/pGWrDCUw4S4aLrthx/ZQXiKZxS6Gwz
P8TA/zWXunU3GaNZhzHsrsgq/m0hO2boXyBgzOUd9+mevSXllOZaMkjZBhKni+7c
op2nQE31KHSQex/ohLt/sT3I1g4OMLW+0avnnRdIBayypkKw7EIEtfBrgxJ8blLb
lZjXcOhEpHLYN9KLn1YV7rPapxTlUomQWGpduYUUbBZ2CSpKpVLN8xn6JC7Yy4Gq
Ik5IqRt6wzKaa5mdAP+t4TTPuionL1vheui+B08bwj0p2gKUif8amMpcP58+sJkf
qTAjvXHg/8YTPGlUGErqqIjwK5MQmQI7ycuwVS1VEF63KezHOiZofN7j3YljgqqX
v3eTeCtGYhc7RM94IsUYcM8IH8smKIzzdIs1LwU5IdJkqfGoisoAGMl5tViQp2tj
oOv44HDYWsOBQFpKq67naqcrt+I7P3KZyDfjIeD1+iDODP62BhRoy/rKHufgS9JP
L1RqLXH78jIGt1n51d4l8sDcfBaSFDRtd8v4temsNoJ8ZyCNKpNogU6T+rnEwNi/
uDX4QR0vTkCJKkrzb4Dn14NazCUxjtnwN1+fYGaSKKixnmY53OvTTF7Cj6k0gTx0
WLObi7Ok8Q5EoF7yb92874dRMJs9kXMXW0zhtOjIIxhGCB6px8J+37mrygpeIg40
kVrn/F4J/5FoU2vvqcdczfyEpowesno+/nSjTlDYguasfEYxlbBdai7mBQ7LFMHv
4zFhhdKrN2c4VUzCP2uDNqHGHjlKVQHsy/2zrPOhl8g8TlnaiUD7XjX/8ALMHwMc
KpfV6tsFKygsCUGGi/CMsVIDbnKdRZ3xxOU7U0QiOlINY0FWqbuqU0Zv4KUqEFgr
436hLzCZNKqtSafrruUndl+yhH1sXhV/HpmdXZXRUInnNxATg3/G1OO98geKDzgK
GE2JYo8XdD70y4ANaukjx0BmEbl0VpDC+E0ikl2k3D9FZzvLvCVtfllvHvuGg/nn
YTd0F45zhZbvSADaMmKdIQg6xDVTfsJ8HXMNXWEqp3uwxPHn6DT0p+7RXHXIzVxU
hIC6IBbvZPFHrqqt1qdakp/Nm57APb/YIWDuuTc0mag5V9uzy7QCccZIT2Qu370u
9GC8sjS8vw/XgiOVdSmmmohhLVhnaZS5Er6yVw8lcaRIZn2/YSSeNHFcskSWsgKK
jSYR1bvbiWy4KwvIwAY4MH5KYxlGnz0lJRugyK2SeWK5lv7pXesKkCF4PsJtpJkP
ibZPhoLIeLAMA3Vlg7pY8J02/t9WQM8UjyjYI/5pMFsMTkxbdgUtxGZqdEiYO+r7
dJP8Cg/hRM7RzyezB64Iw/jN3HY+3ZzluSJgDCLajUB4zloyMx6EKDmHToejy9yw
Q614O5LA9iqOb5tEj1miCmA69fNEQhlIRKH5PzmQO9oaVgK6PKPMIVBa0hZSgpVt
1fzWceZz1w2tCt/SHwIBz9Z3H8hjlA/OxPnPAHqIhH/sIRnCN7hFS9kXJUN2zxa5
0Q2aMXQBtlWv2KE+2GOCyFw+XJoAfClM6H4LfK1amf466czjj60m6V71EK7JO7rV
QC1YjalLbWlL3j56I7CAJoYw4t14FSSoILHvh5ryYLYRkEDL1XKdITi+hF6Bwj2s
cfXXU1WdOBFKai0ykh4tT8M5b1x3JueL8Owf6ZnjeGtpUhCq1DFSoBvqX6BaoN1F
YtWufquzsEDaNV063h53lt+x7rWtvCbslgNTb2oN7d8lxhN+sHqzVOfFBhwnEmTJ
fxhH34noWIt90xrjSH+bZtmF499OsFLPQZZU9rG2ICESKM0KIqwaDz0Hyya8D/iN
6uN9nDnnWuVPthnDGgnNZFtVLjkBZjyq4CYSVJyFnD1/JpHmNLPnZXsqGiPk9YLL
kjVfy28ITF0gj/+6befoETNoadItpEkF5AqxHrY9aPdG9fZljpNYz+xVzEBM0NUv
4PE1B8NRUVjlgNMfknnS3YQFxAOCK/jH7VoV3mr4+7XUM1n/33n/x7JHt3ny1MBK
xibvw5fBR1w0r/BN/BSArPtc+YYllQv57FiSWIc8+hfiqrKCq8htUfPVSuzOuXML
BaNwzSAtJxhtj62jfh15/i2GEk5EdpBYJkQTNj8NJTNyfisNH1gj4IiBXFSaD/eL
V5J3sogQhitFDuVK4kwKtdQJt4UuviRfoCa2zhhkBheSdw1Ns4zvmCMYMtSojdL0
UG9GbfVrb4k/+6YSd9o5peigzlGu/fTFKGwd7vGiJKeWgWMAiz3HoZhN/EyEMxQ5
d7MlCuER0CLtkLWkeJpsF2qnKx8yjMnL6zxcCaForPvsvhOWXN8q3ApL5YxmVuQ9
4jc71s+3X7XmP+Pl2BrlfQVoLPnOxL/vLYkIXsNjzHEHbrYZZmzUGvNKqQceT6pA
wfjBKibDOo/JQHG9a4WKeyCfchEno5TRTdaK/nFKlwI2sD1tebLmVauZzwWAZE1T
JluGUMZuO83bfw5fkn/Irq0YxI0B1nqNJgjvsmzkqdCb4gQsiVVJN8MuGxejtqYG
C9lWQ/d8aJaLBUD8zi75Z8Lxx7DnwCO8w3tcBAtejzFPTihK8CNC6b3R9cfWNa01
ey1BNk1Z2j2SaBuCr5ZYhy4D0eoSGLRwcgpN9F8W54G9Q1DK7VXMBiqyy0wjrscf
z8opVOgo1Mk40BIIb5aQ61bcvsk2I78ykDCdKS52SFkDfUxJRGmeC52IPoMJ7o1g
JOQExYs2PxvlI69/z2AhyWAP9fZJiKP3BjLvSbB4rPC5vyf24ulYruB2VrYbbS0r
vXoj949qzAFG1HLUwvLYwWCoNCQGqIUZaoIhuaB7j8xcQMLlbWDkl07YxKYfCsTK
vBGR2Ova9cr8tbS/Z1y9u8PwU7NRFKMCbrlx7ks/M4ePkMltGw3CTzXr0xKyhb5m
Ul4WVlyAUN3rw1wQ8BFpPcZ4ADKkM2EEIySWQpUWcFjcU4SgdJEuGshgadM1FGSb
KKdReyzoZvGsG5phyoZfbEs3nGuJrKkSc8JaLYexK/89lxpoXoMoQt4SUkEOEcdR
hJVf6k1CP9kWyAUIfWNmXSRS+oe/3YuBmTAx1KIbZT82e2/b1UpptHdkE3TFO4tc
3kSnvz3fmzciEvmSHfxcRrfcZGfvdb12bC6AiUKW06/rGOkMWQGhbFXf8vEpzC9n
jXH1tzXcmOJ7Mi80uvM7JcOkPiVjdkFKu1aIMV/7v/Qo6xU0XgD8lFpqCgpCzwpB
0p1Wy/qyEDodv6F1doPdAYzXDuf28KLC9vS+765dLR+wlFJ0ptUV22YfI6SXGPJq
ucy5FLJGTRffUqoPJ+kiHTQYC+5iJC/UIS+j3Cf+da9CreKBVGjZIM9VbO0kX4BR
jqfLK4x29Kvpft2y+bXEkZ8DJo5r68MzfLYUIP5stC5YEndm60x+3XgNpJTdXIMw
88yL6BvhKd6T7z9whmEVjus9W9jV5EJdrUsskPH2piK0OvCZvkNCNRzT09iEtX9N
RimNQkjbBouLt6Ys3dP++yQUrOF/uLx8XwG8JSTdQ9uAOP7wULDMZPnrrntF8Dem
+G07K/uEnYWnIX3TIhNf0bCBL8UquKg4Y2pWPxIOBjm0Zfv8hqaoYw1JCEG/5rjr
VJBZUI1PnWlSvzUFhZ5I7nSv5vob6BIONtBYgnTGfRQ+fWy5LicwwIhwFTV2l6nK
XE4OaF96JTog1pJZsfEgSbqd8/qO/xUgzggufKQweY+oAzkOVTAz1uiSC9OQelor
r/s5BkAvmRpgsXI04Qga4OINVT+5N2A0KG1YuPl2u/I3n2QNtMgD/mV6jCxOQkOl
tAUt2yljJAOF0TJ+ajabF/58hrZhqtH9hXRfBagqAGSjvpetrhqwbGUcaI7aVT+P
cFq+70NpidsMq9IgmJN/YvxUD1XlCpxQ/2Hauus0Zkg/s9r17rKU6iFMNFbDW4MU
KSHYt80MO5VpdmwvqplHjLDnHzpRJguJ+SqILOQziMEuSH/g2W6swHqbUpTjnrsT
FBVkApp/wNIAHFonjxGs2L9uSOW2iWA2aSDaOchbYRuIlPbjoSeXYwQNjpfDWs4i
uSXzC5DbfWooDn4EOJPXbcl62Hv0LiHeU9WeXgiiwcbWYwxGlnNAXxkFHX8AIxWJ
v+iVuRIVfsEyNAvxbQXkIilS16ZMGjR/Nhpf4aliJGc14FnmUIk9d+aj7mPHxZDR
/jI+MImyFtIYBUFtvsXMf1dz0H+sPCl1pJliMVKZSS3dyjtyIfU78NZoz555jvEU
Hf36SA0oj0ipma5A6eMmepUscXduFGiPgQneyPDwp/cRquRJnJkCR5nGP5/0PWcv
4AVQDv5gLQSWE5kEbdTBv41fTSF/LMuHlyUOEJDhRNgx7IEu3Bgjek3tBbJ+VB6P
BjHOzPqO0xcjKbCr7op8cQMu8FDn7b5jLkMirsh8uf27XEk9ywXJRxg+QgytuvYR
cuh8erDXv0ZzSgoE5w1jU3TpT2xhR23tSbT+1a0fGQC9owKNMp34lfiB84IcFUuT
ok15oYSWJqZfAECCDBkTkqDcROVn56HBI0cHwfcp6i/2X/qwoGlp9lOpuUei0E7s
Tdn9tp28cZ7hq4rMwjVUCgjS51uPeIY1V1Qale5VmO2El9ImocLr1GGJ14TlXeve
WWI61HC12QR/MTipB/ga2Rqv0WD6bqs+/7JAty8jfLMJByaDWrr7aT/l0OHKSgUs
oPiT6gHyxtravZmyUJrdZBvbHql3G3/ZMS3KnNKQ2ARNs7sXfu6QsraMx9qXKwpq
PvkjBt3zWu9qnDiBOzluIztMCRZdBnMKBaXitFQQh9GY2ZWLJnRl9WSMKncI9elz
K9McYZKYNXCjqgtImwoE4iIIG/BzY5c61b3/ASIXuUyT8+dfL2gPa0Bq4KjVVFwc
3tT9QQLzqzAAGgUhcGD5u8TP0XlFePDirZO7LQCpvA464jvqNXhMqoGPvY+DUiBj
8/CCMufipvILiAR9Bl4Yx7mn89pDR+IQXXzMjh9mcySpXybNGgRqXL1exuD8h6Ru
EcxATVJGTngMhQv5k5PzNRoJbDmKejLZ//nKf7ktpUm1fsQUtkG7qAX6PAMii4DT
J2O2AUUw26OZRzDI8nE0bkedvQ+0jupG9U4DhhrpdhPg1I9BHMYr24pT5e2Hb3qb
Pj1ImIMjz0RRdWkm97m7RbVxtUU98jhx/YkJ943iABwKEwJV5Up5EssM/xTYCZKv
NxQZlixJmy8LMJJhbonXbqgzwW0CZFQzQeUfsVY9jQLaQt78wR2VJg49xFN27+qW
w/qJgZmNaW6Lk4KOzhU9BtSNBoB2Ojj5VrwQ57uWk7lTt9es/XSI8oSQNWxKMAuf
MdAnuOYpjBHzRoIdY4CcC5Y0Ig5LbTZCnXuPsOKZCq1+V3dwDnv+Z1vBCsmT0RAp
UO2CAlFjVAonehU1yjC6j+NJND9h6lmCA2d564HWHjP6J88BvoEMsr08c7BVgf2Q
gdsuammiFk18rnMfLdLRTxXFw9eQq4tF8AKVSi6KdO+37gJSZqTkU8y0BLXpatAU
MJalHTMjIBJSBmscuQD7gDxO/j+keo81I1aTnAYYjsX2xaj1X9uUWL93ry5iK10F
epsRpzD7/+6VgMxI+/Lf0hOFTsiNvem9OSEbt4ga6aizrodiUOVQYz7QWLZFf0dO
ht4+w8/vP8ufkPpMhJnxRcDR5M4jAGxJje7EY12r2qNMiHp56/QSBJAlY6tUVsv+
hHB1bYzYfcSet1tak44M53/G+X9wOW5ttRGGUtjqy4A8Be9ZdBFmkm/dRG8s1BpS
+p9M0DZrwu7ZBXRQnOznWYT8+3KI0YBN1DvNSgPknmgLyjNGQ6buFkDgAFM+0vd7
dHDZtw75xkMfc5aa6JYPf0hrCofFPlN89WHblG8YdUHf3F8BbMlS5Ut6a8EYhvnQ
Xe0mwUUU22J8u3VrjW5mPV/r1Q4ZYMoKpekPTehJoEtEI674V8LPOu3CGfoOY3gA
nhG7bIwmm1mRAAhqvr15ligLIoHUb/GC0jd7D+1F8wXGETK0wTzZfUAS/dSBRK0l
A9J0XFbiJBCswNUSxZACs9P6ZRC9LKTPR4pPlTndN5FLsYGBBOwQeE8ADgh1onKv
qMXFTDM6EknFJygF0IVX9wKl6nFiXEePhQeQBwqsytQKnbfIb9tui3Z32rjeFWrD
K3niHEYtiV1Nv5upulMfjgSHiZzRgzS3u0/OjkVTe4pE1FIKtNkbcw1blC3/8D37
RLxGPAMA/eQhfVPsykxPZJNd7+4c+Eq2+zy+11zqJrBA8HvZZOZ6k9H+e0t60KvU
/HOHseZ5lehaOIGJ8viwFFJOV1a3JzKv2LxVlSCUBIV6YfkroPvNHLqMCidSL8AD
4003C/Tq+YkgvRht2AACpThCTiLle/uC7kxp2kP4vDZtD9oH4DPS34bH1TUEWaft
uh4ponC0544pp62AoBEAnuDeB3YVijddVG8iKBbZkC9dZAPorxctqBAM8fBPqizO
O0OGcTx+94q/smvScGtOtGcR59VXkiTUSC2cpSZsEOQVS1I241R0UJyKDK5V3ECI
VavnQYABE+/9IGSZy3Ai3pQg7+TL8B6nz/H3bcGds2aIpYySoTPNpmW7aEFsW+Fh
27e87eYsvxpBQr3qEAx2GtBflKZb33WqHP4UqgIVbvQlsW0Hh3FgmVUj1sS9WGY8
Qw7ZZY04li6dWl3xtDgTAU5qahx1TaoAYryRn+ceqXE5AQiAj11uxiHYVZtFgogx
6trV/YlItX75cnflpWFFCjC4QwJQSGuDPXyUvVTfTH4h3yv6ZJLryR9mezmwO6xB
Jw16opwdrLIkdW3QWc2VRRVFz3jOq1Goy0HOM+f1RY5TT94DR7zrVWYt4pIdhxi7
tejsV9IeY3E7MpcjXd+RqM65mfW+XBl9vBhHqnvAzhkhMtyPbHrFQJQCcmhGyjXd
2TR7UmfFKJjpRsXJwAKIbwBDpnppbubl5q4K3MP/bnLdJhsSdEVpbqkFRzMx/mxC
YQokAHWW89lRf7yjtZkLJh6Iqi0mDBrFfPBFsTByDJ4we+ecmp5tYw/EorVbzpcn
gXhOXtdEzk8k3nv6yP1AnqqMJbcfAmcnkId5u9c/TejspPhow7ZaCLcmCZL6sOpR
Wyx0fhmDjuyCWAQ1lQhlg99gRqZ8lLUrereFo+UrJKGyTsj70YSfSY8z6S0/GWLd
uhjwK+XEam3tbXTRQbFuvyB2rUMk2Kp52m67yEkB97Bi7JlYhs4xGhMXWtXP5ZEb
L76sCS1eIT/wvcufn/rmyiv98AzYma95s/59le8lVJefMmwLhY2tf19wKd7RrFdd
0iv4u0NvQ83DDNz6PUuTXWo7Ypp0XUyrQvluaBIURxscvKMqKHz2mIOJJaXxd0hD
UVVZHE5lHngqgZSEuP0xG1+KFBzkax12yi73kv/MdPtJb4NgGayxUKf3Avt6qnhk
VDLXH7YH436y9eqfgn2TX0DT5odhDHb33k/NMX/iRKPzcPy8LC3qXSGUnnbCU7oO
LhAFwRhP5XsTKVqSAV1JIT0XMBjocui0fKGRV1ThW8FSgz+wK3nzt3ILDw9rJEdY
ksTw8Il/niQ46okqqSqWlKaiACoYjMwe2zZOKS+pngP8uBfKEONnfB9O1mup4oYP
gk5g/K5uXuEaA5ff0ZS7AXt2LsRy/950SEw2qPu24wvD6Wur57mxs65pVgrte2n+
i3jPdGSgHWZiX9Z4UX5e8WboFbZdfrJkrP/haBxAj422fRBydNR5EHfnIarq2vo1
36MDbqa9lsf6lbiEcDcc2vXKLxf49QTr27xH+q78UaY8psps1auip4f31FyN6Q3p
WuI/QEhAngOOUshSd1PP/SRuc0GZEblNtvFme0lJ5SNz8bfttzVsPl9GFDbIXFbI
C1ht4/maG7P3DTLWpRwDeGl6dpMHVQPZnG8q+T9N3SKuFld12sZz3lzvoM31+T0N
9IUrd5BqpeASusEnzxIvgNYJ+u/6KKfm5rJaGvdmiVxJ+53vMadyi4KB/+fk+mtx
b+GWuPTw3X/KK1UMZGTnodA5rbX2/pMjcJa+qeeM+/JWYKToMDtG+5QJVjs3UEnR
jqpUbLtiVXBke8BDEZdekP8Yj3KxFyV77kQ/YDp4x3Yxqiy44eienMlozrPDKxhv
ku2jOM0+ce2J4Q5oaRVemy6M2YCkvZuWc9NFK6kSqLUiDLUphFzpVxm9Mn+fpKlZ
vzWLSJlZL8qqaIoOZ7+80B+yQM7WHHfcTT0kABJiTYMDuI16/YthuCQQySaZbJO2
jZ43Ahl6LRLSnD5CbnNHvh7ZsD3RctxX/kEKGt+B5YvyG8VPATJ4bn5YDn4ID+8o
ZxqTZlIvRUddd0BTOVkJnr2tXLuhKob68m82cfHf7e4rhXQuC7OhYrUH9q3slsC6
Rx49Y5oDrziXl4RsOB5KQErvI6Vfn6we+QFUkOoJvG46HAJK96tfnE6VXu8ZRrRn
iZycxMmj9nKHUIN1T9W6mq6nHPBlBqjCDk8yPEGi5xDpNxO/+5g9ILNv5yId+iC7
lZI638FZvLbZe+OIhE+hizBeitxxo2swCgO44G9mXoJbARt6av5Feqz0b1AKMRGa
0hl2gwPbZyGQoSKGWiuP0sLePK0C56B9GrG5Ms+e9BulZPMMGarnYjsshPN9jufS
uclNPpZExR7KCqS2tF6NLesm4wH1jSMy9mCcQsU8ByvsT3GJWIsinMoOGHxX//C/
xPRlJksEZKRXwAMpx63MGSo0hCCwtP2FkXEASAFp/fN7s9IgL61Y5sRIFsBcv06X
07SeHVMG47i/S9KH/LJUdDm7SLJZPRbefETq0qJkXvBoP/v+cOWQJ004mU4As+Kg
11Kpw8D0FtRQY9OuG6tog6e++ugcU+ks+7ivMQtxgeY0kRoOTW/ynhsUxZBhqUbn
P89HAqlKQGaATRrL6jLju9QSebmWYiV45lFwpWxQOtdbyIdoi6SHEakGN1LuNiEs
uZFkkkkB46qcHoiTCN03+htfRiDiEEaY7di950wDqQOG6ah2xW+8C2spWO0p0Kwk
1mUi+TSH/8rhtA3oBm20mVPR9Go3DLinG4KBko/1IKXwgib4kDplzqg6wdnBkYMe
HSliv8GndDJkjbdp6xq2a1iYL6AQNcLnSBMWqGarUes0ZJmNurJ5NvUEJZAImEum
LW0OFFY3vTRUr+o62HE7IpRo1WIc0o2qaiOJsThICTM43cNg6oQ8cSsFMmQ2cycc
Ox4wPtaXKJHnLsQEZKBWDaG62iWYkpzsSy0SrRyO0KHtlFPoNbD4JOa1r0eX83oh
GXU2fW3hzMbIdoG4YEyC0FDGihcnNQgHM2VXdUYhNbkGFcfJULtpjVLMLwZOb9qb
xEQDNITFuiH1kAmZPfiVQuVy4cdWY3bQJJmBeE0QzBjUgcyoPlUGmlY5Ii1Sgpy+
Q0NNLox9g+EVnH4U9KPMAAVZs+Lt60dAukXRaqmohoawVBHSeL1Z9gNj1d8AIzel
HbvMvt0rrfmkoBAtO2oK8/dccjfh4lB/aWAlkQOJ8c14T2TU9u6CyPbSHB8puokh
/xvMVNdLG4JWWf8pkXo/8+zVXMQtSSCc7kOLnmKbtQdO62Kr6Nx7X2cQu6kLIspR
OzsuikUCfI8W51cXPrKtWBcEvvRGVoUN7xaJE9fUK65fOL2Dge57u/88z5m18UDS
zDnr9CVp9iaulYlxBnnPhDls9S9XHG7bRsoe4/bkzFfPU5fPVdj7Dq8V37vvmnbs
fW/kh9vSgSIzdSnOTEpwbysupSvwSyMBibqADpiJKo/o/jRcgXtK6n34v/DanJYF
KMauQgoT/j48cOs01Y+eFw2vwvIiSPHta/0Ka3C+ZlsJw4lBSATVDY97/JL3uhGw
Rn22InExH/sB/ubBNXds9TGhhXH/3BiOIpsnvD0KTk83Lga9SMHXmqMIPShX6m6a
wfA/yrs5ZoUfzIMgkhC9ohnh/QgWdDkvDgvJh8spNXmPAPmpZX/FypyVxBztSJeh
EnGAYIHYvULXuOdLeL6BiaAbiXOmA7EpJPWYvhOuidlYlCR2p/JcNhvCgjy4klql
04OmY018dqlw0CAigk09Oo2Kc4L+SdfHbyQd+NuH2DWx/kkx0mmCcqOmmgpeavzW
X6mWYmmWFXyDploxYSbZBPWeVwkX2ZqlHhpRE/9ynzCSskcVWZEfWZysEpZGW/W3
mCHJUkO8+bq/+qJdWW3GXN/jTVk5olRU7L2jHRBfUDB6TuXd10UqUDZc6xRgKnSH
jcnulAwcsChSm1Dh5IoeMla5lyp4FsdomaNgdTv8uYkuiIGEhuw9n6vvpaxU77AL
PHQzqPi1RA3pfJDdO/UUnnSAGkao7tNfQBVsq3OLIYowfjThtRD0fpgL9lp/Wv4M
4GvrtQTGlqWPtburXZsXELM71Uojs8nuVuC4oU26jEPfuoYvVP0AeJtFIHiDPl+b
3eytCUvbr+KQ0EtjhUtW4MieoECkM1x6UrGkL8xcYQSaBIuJMBdnRVmYqw4+sKBF
ZrU1kJ36lZ8QsNdAb23qlmPEm/fbeuxG+kpHqxPmF3xtCxDCo4+zksoTpB0Ti4R7
7xdnGm9m69ez4xo2Ju/ie4txdSbIFIgBknRonbjIh0y2KU3zhaAEGH3Re0NV4fmS
X8O1x6PWO8MwmDwEsOVkfMr5UPk//OELuf4Zmqa/a7Em3kKDGbc2bhJ+gn7ciQ4N
iJIkm5ZbINwEXz3yEh4Va1MS94lO/CBxxUwGx9H3ynvD2BFaMnhI9pP4/OmwBsSU
HlHl5+v4X2E2nYH1+z4GvhWCDiRiNJvzEGATWSNHEWV5QQNHMdSN9rfz6kj365YX
nVJ5vVEeylhbcvQ7w0xc8P36r//25a4nAI1wkc2ui/1pyTbvyfY4V7rn8JB6eF1W
uSE7rTZ1YiiIBw8Z2r6ORjoVYeuffmi/et0fCnZrZgF4vxRMNtRGYBtPg+XQXFxU
d/93n6cEjih9YkRiViYKaIT+C51M8CDDmmz0BmmZLMTZrToQ7aGPW3JeKg77Vhn2
racOcQGf3ews0kUB+VZHCkNwDntJ/lZasvHdS3jTTewM4tQv8RVA8Uk4g07tDjop
HRPU93giYce2HLHZUbUG4xGvHDgds09IK9lIfAztT+ehAHNgNv0WKLR0eqRwBai/
FI4pp7ejrwTzeSodr0ZGqS+wkR5v5v6oYqPUCl7CsoEiKTCWBUD/uTdVMHrwUED4
SmvChHU4L/ZKzbpkKU3meBG1JVneC5oGzTBdtyw0ZDvDUDZlwY/nEqTcOKR0Ls98
1gNBDEyW5G1k5hFVAJBZd+LBmuLp8bHIhNuPOtx4vMMc6kwdDTHmgt6K5vS3w6vg
QDkTDkSuEOWX3isoWIy8NB5wfpQ9iZmjewQ0FObCIG8Nl0J2lNrLeQfl10nT188o
h5QP7S2houuaRxzCckb7LJI8Lgn+sSXCzBtKnCtI/65gNiuw4KbbkTPEG+KANlrq
dDZdQUclOyGY5I3aVs37sqyu6UzO/PU7oo4KHmQYSxKA7FKqa4lm8cj2/NYcIIRu
VZ1+pPYbSStmBtwODHIz/0fxu4xLAj0ItGNYCwSgwEnzqjJ191razpTfZHUs3mJ9
5DEGH1lgA+uDXSCdnlTXDz7Hgf8FpDcFHZ6ELWuYXft/Jei3HprwxHrGjT++SnZI
/vT/diA4NeZaqkbmoq+ysFvXvZWhsprEfixQsIbOF059Nrzd48aFk404l08f6kGs
nx/kbTjXBEP+b377qAdxunWGLl/EeEJrN48SazDWBbH2JSxGeToySRMFm+00uduW
WC7F+glhRN7TdjfQkTV3jRqiQ6FR/fURzwnrr6o+I+v4fhfQaEFIbZFDo4VQsU+a
yinGrJ1o+pw+YBu77i073o9RBXC49cauGVEtk9+I5fJIWaPRn9dX0+zbkfVycfRi
V9ODTz1VysdIYrSXmU3+FBYooZ3u/3BLDmFa6aeQwoFfu+xJobLT0/ED6CHTTowV
gPPxiXMcOQaFAYX3/nufaYgSpSBOS1Two7qkdY8FyRMQfutEfdV5Vtf1RmmuPdTm
eiyXSMe+v6HzjRGfLArXaYgmCbVLxXcy3z8xq4+2Y8OehZtKLTLMJhvVGdSQnWk8
x4E1RHa1komA5QkSXbgJjPOniRNxI7cdlJOP/tkIZYD6wIh+vQZeSCqSnRhSkwsz
nukdV7fUIxO8IoVMsm0+ApDfzrjlBpn2o2k+dWmyFXcbnVsBVJ2IgQibRME3zZGD
VsPUMwPA7zccOd4sZxGnSDa39cuoDO19ZW3Eae5p5awkoAA3I4sq9CIIjn61q2l8
l3C38FH+7rOHK8UT+Jq2GvDZFoyMzwhg7CDDHNdxnCPTZoLvHxa/Vw50tBx8pg6B
sVpag1Z9Z/DQTcGkvkq+4QZSPN9U/NU31pFoJchtCP1vBv/0887LtUdn5FxNcbPq
EkEMHy0vGZ7vFMuGZ38QzcFpDLFMfeOQH8Nlv7ckOF7CoUX9iYRvhhmAvgfSBMRK
HSc78vS4Sd16NRD4CMHQH+HzR8CApDS3x8417WPD90V70unf7MmV4u3HV2n74VgI
wCe/tvUhcS8U7c0cwxSEU3dcxYeDFImrNENwZ+3aFpcwNlGyOI9LWcdWSdTr/OwF
0rtVcmyEhrQG2K1fJpwNV03Z7VMIpHiCyZf4OFyvB0ogQajXgbzD+7ZPGTvBA5iA
vQ26vfPZHL/SreI4u9hbuiFoo0IoOWMp6eB3K+qGCKFphzWDJlIqbh5eTwQYCd0z
wnrMsGpdtWhWPTnwrPlAOv+7JbDYu1a5bEVJC3jBVgDBUl3betKlU8MFVHWMDXvA
9nEzXaQFJkq6UiolhtyPIFa34Lzy/tH6WOuKQmKiMqKbHYktw+E9Ef1sLJxYWO0L
keqZg7Qah4EYC+UXj5yizFhQXpXNmzSCLmIDU9AiqiiRG32ZAjl/iX1wA29WOuUG
DVG+TIoXXEozEEABxhMdfVOhYO4bAwaNbKmR5j6QSB0YjdVeh2qL+xqc6+G0vzPb
Vz8uASCQc5B2RejJJE/mp1+2CBzAlFqXHRyMnuHOaQE+EO75TWL/ZM7j5DQLutcW
2PTOyV0/Bj7R1lMYJr3i1EumGRmOQVoe2HT8Ewl1+ZLr/mEHL83WxSAx6Xs8HVNG
4hTVaH8YpQxBmKvo5aCJWRvLkEH8fDnYUHSHn+qJZCxMMCyFSc2r3t9b+eSXHkHV
je9dk3ZA6YIdpdRPQ8ZkPqzT7E5zvNnx4GgV4cRAGuz83wW+nWWyV0XJUwbtj5fZ
gKKZ0FUXGSO9YxAJMGTeTya1ZRKBw2LFax2piojX9+bhysy2LDaVEGufhjv0VnMT
QqoLH0booAemBdMX64eei3dRTQ8CKrRW7fyTzrCB1G3ZTmreE1YmkaULd0HixEWL
p9zZH3ZRIt6rlkK4AZkxInQdgWjqFWttrVPRmGFFagfqHkB+P4i9Q55k1F0rx8uR
VYI3HnaCvB0hE8smKpi/7MYqStjPn3POJfcyxrF0DR5GkCPsJC4VH8a57uvJpUiy
56uRpXbzi1NhgI98968Y/hAlZeGGyBKqPp+rg/OXEQ5deE781fUJjIE42+v2Zoot
fXNaefOyCQMy6OIYcw7lG+TiZTL9EDNrcH/ZUJ4Lu/ctQ8VW61x5bIOddcQ8I2tl
IFiXkwQ6b6FCcnxE/Vu4Bld1stTacW7kADrLqGNbMwSvrwT59MU7RwyyrKpCd7qo
GB/wkpl/HtKTANgs7hw/i65dDuuOkaxsia3y3U1ZIzf/j1QkXQS5mm40OdASCF6o
yPTUqjNfDYcCaTY41t43AJqaxy6Ds8qIhLQzaCJz1Y9lbo8EfxGvwrvq6kpD2ElV
o2tf1I9Q22tzvYZKjkzdNNHxyAfxns3bWkxk9QercBv5gxuOJvFrPIux+JkIsgi8
CnEyV7sdQ591h9oLq86gkQqj4m0iB3pSB45oKpQhwPIddZgmGxJl+c/SeqC4SP8z
nVgqI847OmWKxS7Optoor9LB8LL1vDhtljc9QHVGgHpJRaYrQCa2eLCJS+CfdGZJ
914d7egKU75lXiSGpSfeXL8tetZRByHsT3f1Nq8McquIFrrMKDViu7EDHlbxgDzM
5B957CBe9PlYXq1CeaAEteJ7Nyl7vZQKe4RsL8XgtWTyRRnvcK5ojFz+JIjYYVLV
wCUUvCl3fsfIzy/9uvHCbjjDdMekKc5wJP83G+lBGYkxvfjQROGv3tH8j9MhS+Sb
/fga1lEDA0ESEuAaaMzcgjmNCt1k42m6wE9ihsRpLpgfjTYnHFswwkXiLYVNMH6a
UshvISN2F/U+T4HtsnCKkUp5HrjjspM5KQSgHTkDPeRKuEwonnSd05oOlu83aXoM
vSO1eG1wBA25tfZpcJCtnQ2Dgt6GU1yxddZ8Lg1LWSpo027dInKYKMgUJGhK9mWC
tGBeFtplKmAEF1s1fbPnssoo0rru6jahm9ho5GQ7d50VDOCzQqenst8Kj2H6yyuP
U0ww68X6lVuPuxEKD6ewWskdb9xhlxCdCnmIzHKvCLkOixt88TktP1/WpD1dvF0T
FO74LjiytduiMZf9MU57SjqO9kHtFiRhW0j5XLWEqiHVMrUhcTBjjnM5PG3kmolr
DrMxp2H0ixvH2bFzjb+MHa5j2lZGw2Ad8RI8IW0ngmP6YFpz962OflHmUkZIooGK
8K7pI9dXbWnJhd9Uyd/O8Bi3tJdEAJ4Dr5bt8oFlg9lzUjebLGAd5CW6mZ/XSqLq
tL1QcNk+whu+FkGsZcaghZo/xyTu1JB6OJqMwmoxLM38gz4tT7ozE7Bol0j2Kdyf
8UMuKxJvQg4/a1miyIX5PT/1rwU1uUczZSelUpXmEShG2UUT43ty1kiRxUyFe2V4
Yt4bibqaOtmXRGbMnqjRTZYHzwteYX7LkIPQq3QVwQSOSp5187U7fcugU5BeiV2d
tz8kr3Oy3GJ4PZWm2SDZFxuCU07DCSxipNZyFX3JgfMEkuf+eqr38mDLoUdErhm9
L2RnOSPXjhgAX/gwc+lVe1QIRWeJVPCTyqiZ5XGr/DsLSyq/DMHtMOfJW6cfr9kI
6PQAJMw1V+bsY+Wk11bcexwqd/djbDMIjfCIPHxVdRn+UDX5Z/i29jfZd9ulfpIB
A/uisKWJA3QOJ+IQ+MKLUCEj+Dn+kaB/6GHpwyCvw9QL7XWV4kfGBPu644itauoG
EyQ0H92yFy53ozBY56WjrZPhHS2LrYZgjbVH7bo7VHeyTj2fZLtkS18SzJ6Bj5u9
qLvRaORsfDclySSSRXC2eZa4XzJETU8c8KzZoe60lixPp5iOUTeSvgUqpU61hKRx
9yhE5JBYCKHujlBqKTtf1UolrByorLLaYopsSPZV8IvOXSW1K/g1toaAW1uU5coJ
FCPmk8y14uIlrYFEAUpCO9uV/2cX6S2WFXEl3WkZN5IvyiS5KVPi9DTeNneRSq0f
fC1m8Lf1xZU0wo0aytuB4B4RR5mkw/Vyz98wl8AGDDmDzS4OhPA8++7+IMJm1hCS
LodnRYKzfhRjyS9oCf/NjZR17BQbV3vXmGox5veS5Ip/uu0SyP7W1u31VC5JNqUt
q9ytj+QakHPbHoE6ZCbTW0xAt/2+iTqMh0MREPuR/vhqtgWE0ELyx2WzSXCiyLtg
+fSqVbSDpJRk2S/XxaOgv3UMl3DVwPWnr9XbqL1HfTHH3idsu7njhiU/ueoD8WWJ
K4AYR2Z+tVhuL1+xbj9Cg/2yMXmiHWQ7l9nt8V39vS0+N31iwzCFYxmjc5jaK9CV
72n7r9dYydR0oB0+CHk/cnz+c5HYzfo2RqWzt8gSojtMB53FvTvScgdueVK8Eruz
HI97MIRMbdHUYh9bgfYcvvKBeoYYWqv2FcsUSQVc7O9gomkD0zMmWzUl655UtW5/
/G/288VXxjTAJM3+o9FN5M574FatA58nufQd8zRH1Ckk2eVmub9xvLxuWxtn7aUW
ybUnbrmOgG+gOnvFdKTOxiKX+dgRPdFrxoKM1onmB4AehsnzxPVD87LfMeqnN/Hv
VKVQZYhszuKcI7NBqVaS2zyXVEOi8IkhKs+hBxLhYbgNJN+EiAsCG/Xambyb3U52
AxvPSoCQSw0oXF0fnxuJJXIK0Nx9n5LEumAxOGeAf0mJ2g9FCb2da3dDdChwlBCN
rdj/JSX5pCuBD1aMHh8p/aZoIFPwFBZNxVzb7R83gyw3Moq7nUy5KCqmpGfO03Mx
q8odRuxSMj1keWMChWw0W2Mnn6pUDSy36qnUO4CCtD7ul+SGgaIAvom0wlprJHwO
02FGl7Qu1eyB1mvgrhNMj9Gx+gZ0URG5TZreNncXmSILXCYjDjmqGgSLKa4nNcmp
jZCzTD9VL2TO+luqwHUljnFruDVG7N2hdpusAN51k+XWv7hSQ5uDMYq30ssCHc1A
3ahkhbNl6V5OlG89mZ+4UKGtj3pNQlbFMbOqMZBpdXwBlybnqmu6bT2tG0JWXop3
HjVfHaoBygQw8Ss5LqRm7mbEEJYTcqzyc6sZMMI0GbNX+az8EgICm01YSLqjP0Nz
kdezzMklMcz2L7AJdLZEXyjKmOlBWXWSKn+ARgDq/hfP8L4tyLUcDqeE/rM3b7lw
8TakHp98jc9V5FBnvnSTFLFw1D08Rw6ShpEWJJkK4wuWZJ1OSQmk/uPfbeujsWUf
tXPxXMq5hnOO2QzESqGNYJ7hbOGKwbD6m05Spt1asgUcaxc/g46BAm+bMWmC0ZUC
TcitU/7SUCZ3Cx3A3k7AAU8ox45gkUqSbaXd+JjqVzsbJHZdUEusmjNmcoeLjjHP
Dl+m3MQsBInV5GxYzIB3WpD6YEVSluuz9xYdV7JCbHKO7ihElyRq8Og8PJojAOau
4HRYNYgdp09UVajylDs6ZWpdmMo9fIH+C6Egfn9B95h2hsfO+A3na25tiXcelQy3
oUMGdvS4fvwi2IZpoit3hzPWGq1BHcMYN5dbv3IlMHA10XrQZRVvGQDyo8xdTCS4
WkT1uW57XHrjIEjRKukL9WjRj1kGQ9Xe9pCV0kK0TdNBNctRe1+uxnoqShrkqMvW
sz65VLDyLGEoRCoHFSsdDqkZ2hiTwUvQYWbvK84F1wfaXocsf+tI7bKDH4jHeRZf
YngAo4LSqplcua84jwFlPVEom0Z1QrXR9huzvlHhg7/XBRCujknysR8MdZOgi/8i
8XEeoSAl21MaxtgRdMpHQv99dBOKIr+F4KQo6We0xZgAEsES01WacTeKkQJC1beW
d9ogj0TuNPmgz2tOxFToK4VGeFugNLZHr86edctxj83G4bAFR/vCfKekvanJVQws
e1Fsk61v4aWpJnUJK09AePP6ZKg1CYXDQ5j4jnfk72CqmzxEo/LtYqZdQvT1fQ2C
/z4TjXWllaNuvCponTwlwl16A/co6dPDdY8hQhaRN+eRaypQZWzRSN4CIoLoXAYR
nW2AxFm0U8Zr7AHPONh216YJ23qYvev5tH2h898IcXudmMMWvQ1SNVkJMvZqvJXP
b5qrpctvq7zYi9EO8D8AxEuSfvcaR4JrZAM43+a3fYJ7ADdEKxoeBs7LeStjSXpd
OT77OzjGRctCxwXEKVUdogcltxcYhwGXOKUAjnnT+XVG5NXCsoan2e1g8iQ8GPe9
tJQbpz+/43UzvwW0x9FCV3Ixxh+LTVUZ9F1N6Vw9+c1Zto7FcoQOd5foTw+keWhu
FraDSbc8b4exhskw+E7cOakqo/N1RgP8n4hhy4bvgqTNRNd2LfUlkXGxdMN5tXMy
4SCiNPlFkA2s1ogB/1lRluOHHh2/GQS7VqBSU9fuMLsaee9AksoEyctjZVJNcqhK
vaSCo9huQ8Wdk7GH20OMqhlMhziAyzJ27TkrpAFylRuTK/HAJkEaIZmXtbq6DqM2
CuMpv09rziUMuqboeqvMo77+bPBAvilsmwGT76RK/uwRe9mZlaAy+AtEKPofWBpt
f02mgwG7aDc2xv8/8g/9QEjnaEVG98Kzqeil/XHYb/AHTOhSGj0j4jhgHaJ+qtGT
E7rEAYhamNItwanr8JrjUFB7B2z444l60egvC19XClRz7ZxWwF9Pl8D7XCE1VHMd
gEv8iHCn1QvZBkBLQGcD21mTU629Z+lOPK2KfFSjPpOW5VnE1CU1UFQXZlnq7D78
hg+g7JPtrVPzSJZFVGb30o0rXIJzpbCLYrsz5NZ0V51b3kofdo2WqnQhDaqHRHbS
tsnDWHyQXu71YS2cMT/FrJIDaa7YleE2WscDV2QB/VASlky5vFiZdknyM5Jmk5ol
3BgVhBG+VTU1vzVL8MW83fn2CpOnNRhvbVMH9FikU63gPoB46bL1kBTIOGb63LSI
abKTvgqXmMZGKE+i3u8xSMlWg4Ic28xRdwSQm3MpXsE+S7K42+98/sfercJ2RJdk
/+F1x2v5QhpRg/lQRz6SEnm0gUZzfFGp0X6bX/ZJAkfJ9u7DRgyi2zHKlCbFAi/m
l/QYu8uAjYO5ascrP1Lsp+BJ9ba0Aj2Oytzs9xvUDiII9CBTW3E2hphiYVgkW5Dx
Z+V/ohaNmzJRb4XNos6V75fPSfD/Zt57XsURrE1r7lpIP6P3CSHBITzMmb38RHNc
oDszUmuAYZbDFCvnpdP0CA1sgwy+Lie5byQflqtE4lSZ9woxRmTHYvLfJRieoSX1
Bp6/XvdZEJYg3MtZ7kSXVhhBLfzzo+xRe2GwU89aTYBBJsP6BEgbjMBCAsIPOyul
nsuRLpsdBYqSP7ctHu7zBfNr6YmK6NWqwxxWCHb5GN3wVnAHJm7G4Q4olo1icvl5
URvQGqXDqKORTEP2uWBxseCgaQkF9Nf9R4pjCeRyPnqofv5Gngzj75Mg/2kdxd4B
96PwQBRas4VMNh6tH1Xr5soOytlzJ3UUwdS7D+dPbmg577gze8hJlWgNHwHXWFkF
shs8bqXEKeshj7GZrrKci67v8mIYy95H0WK8W2wH44UoNskt+76FJLaZMSy7xNUB
wgh9YlSF2vHpp2gdnxG/PTv8kDsvZLVZzY+T9Fw7k60DN5+dTvsg6B3hD+X1d2YR
aT2msQz2PZ6fNXQiDNwacUfsPypBAWmYh5filml9t92tLDr95q6uSVfe0P928lVi
PESRFv7ABgBFknq0itGYZvWu/ujhTSmoPOXKU5sUa7s4JRxQXzMfs/F1NV9ZtsHz
W0eLI8QHyKSER4uYLSI0DQqW8iJ2hcyTegJ5bjfin7t7X2JjgD9zutTx/PJxJJKW
0L0Gj2SXy6rFYi2D1wq3E8bNw4L8pAw6aEqWFLVyO6TMCdnL1mhbqGnPehHv6kmf
Zbzu8dayVeZBHCkUGBddOIFYYKzAfhoC6wTDfDRq0UtpcjFtYNj0tZCNg+57nPyp
Qgq2Hm1tHp/Q9fO3VXArmcTcEAPiVcrmhmVrb3VROKj7ldbVZZvPdIRgQYQqkVZw
oSB7OO9hOn6IEqknJsymJiqZwr1/nsPf2OGnOa4F5X0pFp68Sqro1GJwsiMfZSCw
aoUIrU3FBNyPbjDzwKFdjwXV9TCPH6GGw6SdCDYoAloBSnqcp1VqkrHq2Qp09bm/
mj42SCug4QU6HVz5nTy6v7XIO40VPCjHw7Sm965UDVg+xM3F7jzYZFo+L+vwknzA
GdeZlSTFJWzZ39iL9e0Z9vB7YOxBaxfe5q45Go2ElBGw36HhMgByRziRwOBGyr3H
RJ2bvyKGPw9uLVpedAbEXUxRtbqDA+y0yDP9SVw754k7QOy8la7RxX6aJFALDAjI
jycJe/Wq0VZfIW6eQeUOf0N8b7wfXKd9PsdANOVFh7cpq7i7UFPVoIkcYN6ZNeVo
W7+8rm7B0pVGY80qR8MTVpRuuVCcynmenjH11XHLxSnll5vDxZ5xKuSypYaTVWxA
kR6+d7EgS81Ec//3Xv7M1HIMOnXSlvgZ4aMyrosOQk/6xrIfnTU/9YKE+ljFLFsl
QybWx+2XpEvyxluLaYm0PZmvOf7KwS3rY+q5x0qYaV6ArW+X/D5NKMcRpTNcG63v
oyZmGrmBHI767cVd6pyg+z016LFRI8DBZwdvXDgCk1j78PVM8myBrC6Dgi8xmB+A
gG0C1iu7ZUw7a2wcC3Ai1Ro0z4u5Vg9Gi5pOfpBnWJEJGka7EaTBSwsFa9LPJ5/a
a4y0FGHdc+MUO7wWsrdguRQ5v4GA6iNGO2FDhbBEqspBg8i1llRl0XhqZCzIXaNd
ebz12L/2laZe2AH44Y7Ka9yKi0o0gAZHImFuqNYYRxP3eFmPK57Qq7JlF4OJ3e91
rTKRfiajyA87tVKw4yZN1zT6I3ias0KctkPv7mI9DqVf/4oI0GNla7c5bqjoaRuq
2nPKt2gNqLm4c6IdAChoPI9r52bsppP7i+tlv+2y364SgGWLB4LdoVfMeN0d5XBK
UoWKHQVEzdATHjsyRaiUzYoJzV8I4Uqsl0+4eKYyO5VwVCu0LrOoDbjdDFpqtayB
zd0pm1aP9NEouWJhjc+qOXMgCDBXjHbcaUW8GQDCrNSc4lun4qAECB5W+n4lvXiO
VeVCGnbPsZj9IaXWSg2wSJCd9h79aZ17n9fdPqwDXHAfdBxw51N+6NEDbrLaXxU3
iXiPZh/Gd+W8f+CGHkwsg/1k4j5vf7A5E0UIVL4y4QB60AjELAgH7tqxC/+oGUi9
IrY3nUiQRaz5nS53vXXMSk1ev7Ab6aek8uEnI3e9wlP9lB0q3pSxjrSam0fWFisr
jdDUyhtv8klO5P3pKUnvGMtrLLjVwverodZj26Z420I+nyxVrncBmXvZLOfvj2rK
9IB7n4/BBWHYRQ6+6eCd5slw0dGZVg3uIZijo29OEhigg3fDlCldu4fzZuktRkej
UsWjAx4LTNTS2hMaX6Wl7fr4mqGxYZ9dSJPi5BncaBbgkcGedhuCuq83iVEc4H/p
4rfqtJ6y3FR2SrqxTDvkghEI+l1js+KiHrwTgewQkEOYiwqFTH0OgQPTx7XGa48P
yEnnWkgStgm7MuCxYhxgi6DXDVd68Cd9nm5YVS6tZZ8qE1+NjgU+0rrIKpKbY18u
Ss51ArJR7HQVG9aRDMkqKCpI9+DVMGgsPSAbf++iktm26OcMxRbthILbpdoX9quC
LDDCsHdXBX2KYtX/p6SDc7kslVl5FInO00g8KIpqHFT3luSRZiAEoUEHirembTEz
CClFR1hyyyYuQhbxQX1XKaO2nVI5nsypFx53fjlaAHjsDszi3n9c7xWOHonCZNZZ
zCZKvQwbA6TQefnuWC2XnshMk2A4Sczf+IadvvgxZcCmBze1/5P/RWECUOXAbHp6
e+hvvvqmzypai35gD2Lppni2s9VPNonsqRATavgDx7gQMeqRfbn9tmYHuU3DQqDu
W23VPRiWoqoAag3qbywQRI2cMGqEyvKxO88UArbN8FQ2dlfcaGihbMuCf5opEpob
EIoluA92Q/JNcIoCfdxlhqjKKnLglQjvXYjCC3Alvz/gi9yWsxXk/m4jABY8uqzh
zCBadRDqEFJkyxVSrhAVDrnltdMTys/9lY+YF1xeGaaLUb/1DVBJlkBfcGDEqBk7
iqg4ArvpHkBy5ExRyPiP8YvuD/3lofE+ZwDLokCmEzlM0bhv7K0kKpngWkitLpTD
yiz78nVnLDnJwd+0FHHmVV3w7Ed09txRQ4DmlesTceaCFNdHcfB4bpK4oWwFAs9c
2E8SgukPg/SZA2WFc5jTXEL591C8detWzJEKWJAQ9oqG3PzlUj4f1VEIn/RNSG5+
DJDtaSBZFCrBFvxyIwBeSj6j0VMYx9Y1aj1OS+A4/RqH736zNchgBQhDzpKhHjT/
eZw9kx+Woeyjr9Rl7Ku/YxEga7GYzNK2lADexvBU7003vsZO57SpJn8EHH+CQiTz
FhLxdgsteIwKbFm35zs02geHoZNUytcQ9G93xTu3CHnIKrBFk7ksYYBN0V7TlNJo
uloYMGdr1ql0ucdf7gg98MuJIi5wsK9BPIOgQCfsvz65/X4AkA5YMd4vnn/wNGkE
HqscI1tg5kpym7NmCvHTwjUxq29wjx6J0L3cL1voTI2i/Aj4UVn8lVJjGRfZR/ME
jRdbewkmEijaEBA00e2C4L8Xk3JspdfOe/K8r+j0QLF9FdMzRGEPtH0Nz6CaG9Hx
sWVS/gvx2NsKAKNkrd3LTbLAPw/ddP2TrpIvl2AkOaS5g4A+q3YJpjdsbVKyF774
8fMuooFuipRFrRxjsxWlBE894hLwbqtjNFuWizZPNOnp6N7aaKhXBWUkd8XfzXSN
wYuM4WJg/oQ07WNMpIqSPodRp3uMjGCsDoalF6RqI7bl2JKmE7V4UL2raeZenrH2
NRRlHknth7AG/6F7q5NPUiB0G7lz9MgGONxlF+uF0a2UJezy4mW5Z5TV2rTNnRhW
pDZcMavL+Axq+0m9mFte3K2R0WpLU2OeKYf4Uc2xZvwIBxqwlJchJz6oXkpNAUm4
c0WvE/lbV+9Gi+B8YRUHPpPK5dJ+7GERy5JBuxy1p/+6bx8bEdiX36WcMivg/bl2
QWdl2AZkbuPL1d/x2U5ye1h5kFMXoyn+jloAOSfAK3jeLjSi5SIDUCSS+Amnp7lq
1l41Ge0ptsldRv4t2PpK1SdNc84XeqwpvZG4r+h2Qfj8SUKHQea8wG1geScOZ7dG
amTTNb5r2s2qkOFtdyyv1KG0xwvVYmTs0syKdBAim/qcSmQ4kLA2lHaHKfXiqKmv
s777tInAcy6kHFbC7fASqQeR1VdhUqIQK2NZfK+CdfynBdgFFRDU/Hya4CcU/jiy
cMunozOxM1foQon6RoI98Ms7FQyeUest/KlTabB5Qvgz7HhGshEjz3pEnVPVmS7m
ZORVveYjf6EfsBCCYfc0NsUX8hKvdFONeg3DAGJ6Smh1FABin7v0xxGsgtzVhR0R
aOrUBFzjP4RoxmmAlJdkOimXRMEhgiXqx56dionTbSd+BY5uJd5lV6Mq02OVB+eB
fXTNgxdLq140WYTF5Fv7nFE2EFpnE+eiBqykBbSUXScJuyXbDxL+rTUbLRu0BO35
8MhgozlAl/D1lyawGdQ8GFmhS9eH7ucaS8MXnUxTlJi3UK+4fI7mBvNUDV/q6nB0
5NmaaCH92chjveFcyTiLxpnnxcxZj8GSFBeBYR3QHfmLCHjOrXpG8wF/E2U04mcw
hnd366HjpREiIHDua6ZQb+VP/YPJalgglyz+ZSU4z+JmRgBAUaMkrjthtmhhSBYx
cfTgz8+SEoz9pY3dTr2S0c7pPnSVqjjqaf4h5GpzAEKFyEs/dIkaMC0cCHiMwUfS
PurKyVtGhkd7QtpwrpDk1O3iuuRM5Ln4l9FItHA9Y6F0NgWzxIGXklu7M3xqo4pz
NGrDmBV+B1YbgeyNqZ83RdBrc0DxXGETYcAacgqrUzMH38GBal6f/BMhEnR+1ANl
nFmiuQbB9O9oVcFvtc7T9+RllRUfh4Rd92J9mdayC6lU9JF3Ivjgbqctmk05Kcr4
prv1pvybaqUUoYjwqik2+onYXmHnrv0AJlMZhSivoJQ/rqi6hJP2mvnLUzS+y6sP
4sgDVQ8HCs5oDe94bY7yu0PN+GEkNZgRegNSGYZS57wQlMWvxutaXDl7XHgyC2Tv
wKbxlmnTUUrtehD+Nf7nUYTnLMl4Om4/4/Sr+5ECl0PHqUQSMDunq1spiVI3OAl9
+zsxh0U6+UHtPnTCvfUMzaqooiLrqaZ1R+nr4hWf4WbBkmZ5M5bHq/FKf0eL3uM3
9AWXVsKifcojdeKseRNkuCCMH+bZZ0cF/HotGZBIc6DwLwFTFXoCwmeazLX4C53T
7KdJU30Xuz/Qo2AuPukp2/BxBK+db1gMIXrjWPGESf5roakwGJnPd7e4pW6sOwny
Uibm3eR9E4K3IRsOVuogTUZHg3VyGfmXB0hhpKijZ4PtHLtEqgfbMlGmIcjQZ6FT
DJmoGYe0HsRIduw6HBWb4Mzd3Fr5dcu84IAf7XIL12dUl2mqvLRdu8aOFQBSf6DL
UToUY0Ovlx+Zyzn6Y9mtffsasGQhzcU3h8rltkzrzGjb23ysTCO4WX8km7RmiVf1
oFACl2QMkddg2m/PY54VMrdhXOYCGDRR4MIfIW7lTVKuzYLsuYdUf8OirSmLBW3q
INDFj+kXqABfAkfN2t6Wp7gaezXODseAfHpMaJVcEhhdyrfIbwvYmzOz+4gfvvcJ
1aVtiqiNe6pxgdYlo67ggUzlY/jx0BFfHOwEw3Ub8kFs8zkNSBfYMusPKq/xBWBE
KVtM0MHAmKEHkRDGE+ITKSa0CZZMnY1EAPz9oK/3uSRTB4+4Sv2AogpCBA1vWUpV
FSoKNxJrKM2yklSdNz3noodbnaLhk691s1d1kPVRrAAFlC3g8tqOzxNOUFnxe65U
pyXMJMyThdDUSK2NcG7FWqLheRVb1jzp5Td+y8DAa4UPbW9L+9SJUxwr+rYFUoux
ooZ4bJOFq0m7qVniOyO99VXHLRBeEYjiN+rUMvdE1C/1BkPK3m6uzthXPzs3+la9
QE7plpt4nWYWdhEzf3zFkoRLZWIaHHIztfUruXowepdgW7TzL48MVbmqBFcNfRCW
kreiY7CyaWOEFWC8g1r8FR3e1H2aQGnjTADogbiXDXcLNI8/wrXAl9DPDZnWzo7d
lZbsWvcTsoS/dMV3oMoriN8AfCNtYC3rF8lckMu/55QDjL5SkMdGzLrtGjaXpYyW
EOurhGjUD2qlvKpNaL2RQM6H2UYPGxAo7nw35MZhneFGTZ5p2CmU6r6ORa1Z/2PI
GTrhxANRG8PzbgO2tRlw1ufxxVn4CMLirKh7Pkeo5by0KL8Ju2Evy611pEH66g+Q
Rz6NhiJfaxgN32bJ9KIgTelyasPVvA6SJlGECYHuDAo4h3b+qD1rgmNeGhIQ7tCy
cR/WV1a1rA9Ohx3EbZ91U/HOeej51gpsKyI9VfdoL8+3iCep6jn/nzhz/YgmjrI3
7ffYTcwmoKEfNkFOQzlfre0XdOZAKWMSab7C9AtmI9Yg81idt5TKfXrs5i7CgF6t
k7ZHUXzmYChuQWo64UPQytw2P6gr69d/O8YRAOlxHfhCf2yMArEyXbkGxmP3QgPO
g2NOUZmjONgXQ5BFzigRGDo1/qQxfN77fbHOby7XjjtZjCK0KnZA2W3/KIIfkNed
yAA1grLagYFGvm3hH5TzK7Z+mwmwlhNtrus8utVI7PiA/bHcXoSwlaVsi3yLFmrp
HC0NCdNGEUu6PiJ2CAktbtEb9bC53ZxC613PDpuqRbXQCuk02gNqQ6Pj9WRbztcU
RAImbuEdBiONt4YQWn/zCgh71/oWPc3JPFql3d+Pdixi8/gKWqTY5sSo/Uvb/Ogc
SUzvEK06Ct9l6ww5uLruf/k13IjFX7Phch+S/Kasct5rwm6Du2wMbqyfAsjLbleK
wPaByfp/gM9ZQbpwlgCyPPxFUT1l3QmzKJH51nddw2MdJOtZfqSIUYH9hhfoaQGo
shOIyjjhu8kyLUVtY3PvlX2AqdYRbyhTm6F8ozZc2BIePhT7LJTdZj4N06ncDJNi
krSQXJfwyTiXOLIFObEsGZ0ep11XLgkLDFY+erVNvS57bAUNnA3GQvuFLaLT473D
fouEdnIe3jFYI+JR66zOCccZ8aWEVW/HXKEP6WQbmM0FEyF3RflFGRQD/Svs/nM3
EC4QC5AX9SWv4VYBWiqmPiHBpvILwaqIMIMZ3tyZEYCCr6eYhAhp3A4QYFa10Ouo
AhaOzk9BHHjseaqx3XyCRGEP34BLc3Bb3p2HOaIPyODyoXSWVWDat0XcMNIEWs7+
rz89FDTiKPJBoFFL8A/SgvgfV0RgoQI7bcrJfVCUI66/USsXBeLWJV/mwmETySO7
QOU7/oC3O6d/Hu+6altpkXJxWWOMqcillS8Sp5V0I8dlPltIlBxh89aIvnd2iyug
A4AKMZheuqju7TNT90JcGc9LYjNhe6DPdGs2GlKhnZOpc6q6+FfDZ9Qx6gyls4mI
wOw57xoNHHNb15blUf6XaoVs2CYBNRKXIjzDiIxs1Hh8HDYzsMsTJi7QivCcmTlU
onIMypgGJaZjZDhgze7/MNrIzjph1AgZlnKt/Go1qjPnGZOCfzTTHvBfI0Fg5MTc
U9TsxA3kFrCNfSTelHmNl+4uROIpcBJrZa/6DhEn3UW23OY/sGwX21px3PX8kWae
5NgKchGbPtnxWb4a3/4dl87j7eFRlQEr1OOmKvGWcguLn++Mt1FlpK6bR+aPKdKa
1NDsdeY/nxOpR9Kn7u+OYLEnLMvjhUyjw/fIkJhyKgKEKJ5ujWlwPQL9RkN3jSP8
ON5+jlg7kyTiKre8DobVqon5CRl2kB16oCgRz3g+f4N9uqriDwiL4ojfDFui7HFt
mo6l4ZRZxB9bM2GoMRIG/7u0b8YCx661pkvMaL+kBO14ItlDrkr7trTIljFQdvO5
u3GRrbQmoENoGI884AVLS9UlCLfPsz1KfwRWhgyOVrJqLeuM7YMFp3lo3FuLuA1v
85iD1lUZIVhAgUKHBtGxvPcDS9Mn/imhgfCgNu6CEsUs3r6pCoq/jRGsQgowhgxg
HHlTQ99PPqJjcjMvL5kLAFZ9Fb8ZpPpg5Ht0OxvC6CbcZGv0am3YwwOWE/ZUzTOm
CIeVzqjsqRH8CHntkaqVKAwO/cr1x4+X9TALcKQJ8+47IKD/y2Y3eRjfSfQsFshK
bBVQkxJC80OsRgVs/FNeeAGmmGbLEWpHXhnX3bOKrXrq1NM1gC1gQzjk1KwjimHF
k/5UUiQr/fSg+bPWEbF6o5ulJuqsfBe7BZce7yT6z8BYqHRgf+OMIsfL40D9Y0DM
LKr5VuoU34f2e6RYAy8jj1Fv4V6TvKrxUCcf0AIXJcyHwyAVUm25mUfvYRlDpEo4
pgG2pnW+qtUFUrd8vZn06BHQYN0iqbBxQa4TafKf2lXvKBjqcWnXjZaeGfKGes6V
ZYKc+lRErPuwwyaQKowRZVJ7r61GUOtAxrXkCdkQom4Wfro2P7fjy7/Wgg5hghxq
Jz82JP97XuBvgba4vxueRp0Z1JS8n9dklNxSrLioUqSwbKTmuot9zZb7TpqSW6dU
H31hLwU0zSEf/qeG6ihLaPR4dHv9hA+VX7i0s8DeGIbf+7fi8Ammsv9s8ogUrcYz
5a+xfKx7EqJrTudssbBZ/2LYDMR44ahdNRvwjJwcC6c4jLmcalilLlBVzYeC+4U0
AqZHfoM/PIiP/0g7ycV55fqPoRMSaDPGxTIHds5GumvToIwkV4Q6n3TJmwuv2Wr1
3SctsXb3G1H7Ou9Gek1iyY017azmvJfZI/SqEHRv3ykHz34/nvnN0KQ8bxbXOXuP
H9vkzseCrTHZU8jvkg/KMnUnkqQElsvGFdiFnFxvMbl637gqXiryqBtrdjFUYvzY
s3mEInwASUumEUA9EQrhYm++YNp6kWPl17hUoR9oCaiFOnb9dhUzPkA7dklg0zNj
swEZSc7v1qG0spZiaez+cC5nUor/NUASDHUvF3OTprnwBpPmvaVmD2+StMax4mER
iBVVbkDs5B3Zxx1sQE4Jl+8vpUjFsnzpYju9Ze5OupgMEcRYgL8922Au1wDt9D7g
XNIWgS/SPNmcUHIyZ/mNZAClOgt4XWiojbgrK8dfM5aPULXgLQBmeSSLIrD+ppOA
LIR4cTaArutJBgItsW5NGbw2qmi1gwlQL6JvF38CHec18hWiJ9gxpal7PkLQR3lq
8lkipkMADo9quqDCWvVTnfOZlMTAVh40ecKfyDXfTrqLT0HT1rPbxzDk/gdDxE8G
JT3fVIYCQunqfCDXM0xygLcW4X18Ig3kh7v8BL7cjnEvta7J076ewMFEsBCYkX7F
gEOh6BLSar55/Hg/z2dtSWB1WG0sIHKb0ZrjZ6Hp1JV/9Rr9P3UpBBtjccSYKqVF
btlgRn7U0PEE7hmLRy6AQykiWU8TxRLyijv/+ypRvLZDy4xnIdQQnchX/kbdgGQH
GmxjQLQ8xoD6EJOVR3A4qsbaB5UFpukE3sLNKPVAL7a2B5wi8vLEaTHBWMPSI51v
+UdMgkHOdKyTy8F9IiGsFKxSyRaRsRn3J1/rnU2rtwk+liXqBh+qoEigMDWj7a5K
ZV15uwHnpuR/8XbfQmKHM/mO6qTO1DrGOmlHx/uwcrlxEKyk4mUi8i972XeVGa2X
lir2DHv2rZOeG3zPmdR06Ge+dt7IU7aS9QnYuFLSdKLd6Xj9F891ShCZGM1GwBOC
s/UHugTw6Jwlab24p62mzB6uaHLJGQOgHWWCyft43/vunQJHq+jScnJ8E8wRkbSz
0keXQON3Ewy9+YTkful4et5cwgSgyJfftel4+bAeSGMbX7xFEUtY1cMZsXhNM55j
VAHR2WbKHVS0dGU7bGUW1fBYiMLJxYd/raZyOfLcLUrc/zWAxzeaMzd669djR1Rs
lqA0q/OEwkKsqGTKjuBGz8jbqChOJ5aQnaUjBkwzY73VZV18VTaxQlJz0DowL/q4
cm2qk6o2Qa5V7xk5LMN+wIWfCvE4EFW8E5t+iwS2iWI5N3gRkLaIIdfI/z+lKKnC
AswB1kI5ExWuqTd2fkk5+xCYoy5cdchhj7nsupq2CRC57oB510zGM+gi8FHf0P/h
lblVuRe47V2AETFJBUiqF3j3Tj6wW0KhkJ34smv5XJdN9RgQNxTLSGc/5X6tQsrw
nvYJ457ZyVyQuQ+rgYKd60f6AdytOr3RmJB1heeWaCVdUWNL+XMvMTWWG5PiifNG
dwIPgzVeJGDLIS62STcLhaQvOYKT1nnhwHjaL4RDSdDFXp7q4vl82lCsKUbyyt58
xpQHVSHLddMflCTI51ASv5+ALAwj7qa1tAmtNewS6Y+0MB1Xfa5SlXeSus8OYSY9
Mm/xHfJLdTnmEoN+DWVOpHsRHTdJpFK/s9qrb1+ZO/6YrrOtxVxKw+LrjlGdDxTg
5gy+GKmPZIc11R4GhpLqN/R/B9P4TUb5ExKTPIJgR3rLSnP4dXizfbzqPRXGrY3a
TKvxfbYrJaZUOTT5b3Bk5vAwlemEycz0zX1NrXVF7e8NTFgPsIJIGsIb4Rq3BnyP
cnYM0F0FvNCDTQ5poYd/InLSCrnS9Eauto0NpLaGxbIIuJd1XEelCwbNGAJy8IZt
LqvTT7OCz8oS4BjPUxUc2DEvDMACSZ60Z1/14U8YYnUlubkD2iJGP5jRzirjRQSG
7GmuC1EVKK4As39r38CXfxP/jjGRg0Iip5+E/RiZM13zOOO//hq8x4OogSzRYvGg
1KvnzDQzwkfUoS9/2YRt0W7Fams47R1llQsKSOWOwXOofGjTemXVnbxlRg08uGom
zFS3Fwbuk7IX6b2LsKnsp1CQblgiWZZcDAcJyj+8SPVap8WwNP4ZN0SLhICzQJBn
vd6vjnEr3kH/yAf4UJ9QgXG/fPUeNRs8gcUP70sg6VtG7SV2tKS26cgnkhwnCvr/
3uVbgZqsNuemE75wCLfDej8i8/L7gmITWQ56h8xwNBLD1hIEJ1QKyzKk8DqhfyMc
v4BOcdWayV03+NNCkQqwy23FJEXk5kO03kjVYQLA6nc31AepEtdyCu2f1i/aWckM
c/x4F/q24VRLXhFpRWHLLUJMgn3++LimsCo30iA5hGajBrez5AuaqCUr3Spbi/EA
HqMcHpn9k67f6FOtFHOT1Dv2N73q8ZlNz5JtnYycrH9fYNAjU1zKtsUehJN/l0nG
229W/XZLV/jMiea83juQykE/hcWx8IEjtPWW6mOmwn3lufSQCxUksKIKuWZea3Ll
XVTnl+QDTpfs4fJGnOsL3uqKijTYU1OuNtKKe9lA7Ox5FFV8k674b7ERYeA4apet
BTaPVfKoyoHYAOGXkuGd/mr6cI2lqGG+EP38Y1SBSBmUcAMvFLzdpTOWvU3JD/wT
/ClZ5kLNF87C/SId7WoHNp8s+DQDL1d2xtHVPcXhc3gdFEE7Z5MKusDznNH9iZTx
25t2nbRcUILyuLFGXowLS5/MzsyY5PaF6b26E5ZsR30VypFQW3sqrCdXb+RfoBO5
vPkcVUreV/21MEsNHOE05qICcCydp4+zzOqwsOFhi1lS/DnHM4vENPo8Q2HpD3pV
g+/PXjfiTI7IsPL89iMVS23fVFQUhFF/JimIr3fpz8ayq+JK5RTvaZuKzvOCE0J8
/JpGPGyK4xEPFUmJRCKY2xPyVp75DUnBltBazjeRT/OARlGqIrQyrFVuFArLd0x3
8COSAHGgWO2PmU/ELTKL01efBLnjmQ3IuJIu7FvF+DJAYfNeOAC2QrQmQ977HHZZ
AOwPNU6twUSiDlG6TdDU55TYMcV82J/o4r45N/p6GxCEb9sbTIpu8K+R3f+WkEZq
XDy2IUXXRCTm5TQJg5BlXcBHVKTtdofTh3n7RZCt0sOdCVuNltP6l7xMiAZPHmF+
W8vTXfneutVmNJoWcg/Qpw0OX6wgRY0mMqI+cZPgicv82yII5YHTEpZTuLlse9z4
8heUj3MQdrulTgynX0fCsQ1vxwr8SVaJY8UVw0NmTPWmvEe+ap3aksyr7rf+WROs
gPmE5JCMYB6zKl1qX/kmL7WZXmNNdJSZwtTNCR7+umYBSYpiQBnZTfwyVohtAUVp
4nN3nI9wUM8vpqUOLeQVQYAQmOZML24SPGsQbMULvn17LWNdR5NrX5SNRamE43eg
IXdGA5hjAef2BLpV78LBclRDQzFTK9zT1bu/Y2r+eSx3D+LYE+VoDYWxtNmPqaG1
vYWwhkXdSQd/pzYhjyoKP5JU+tJ0zGJyTVsD7udiWDjIKrj4Aj+xYJ/f3QgHfq+i
+Rzj6qVw15j5xfOoc1PwxwG/4xgzdLxTUp5IKvmy5d/dQqpMxn87RZxeP1Oi5kvW
hs/WEFsNMqoWrDYXWrN1qN5l0WaLMVzKj8lbbJnXXe+5TyOYo6Vmgn8GIWq9Ymxm
+Nd6CMCb3RhGvbSVRiEJ8p2/lf1squwNlI8pmt6jgSQT9zSBGHt9lCVDPt9pT+pV
SCUmOu9UTrU/pS2iQFzOlHdK5HESt+f7olFvQgbdO3VULMAZ73l/4BTmOaXhDshw
MpKzJgf8tEE1yfiKLpVuFNt4NxLio4/mNPIExxXId7prWdd0HB2ctkiH9POOWHWi
UCAuFrH84fKmlvxZMUm2H6KwdReOGYVA0pPJtSu1XTA9oLpbIf+MwRUdpVEzZ9dZ
tnQYV4J9nOi29w54CgrBt3FShMWIBEXJs8QpJsPJ0GzwFoHbYyT9AMJ85jTMzaMU
8TuaGdlZLHsdf6tTUm7DhM423XouGo/iwbQw2hXk3uvq4u3tg1VOjCWYVYy6gGBp
8WFEXi1kHzdx3YAkp9D1ql1U3wFUQXmSO+Hung2vyWe5lJzBv+oXoIkX3RS0SW5T
pQpPjLYZV/962JxcJKw8FuOaThzDGVnV1e++mFgZIxCk0TX/pi1JZcaepwlYYJqB
9/n+DI+kjFskxrpvcq9a0wRiKSIUOqxy8YtBRrLPsncrmWODl53PscjXxFsf+35q
fAoPVJ9fYDAX4HcdYLoJfGRJCh19gy+tujNUtrBT6BKf+0+zHo6WSb5w+i7Lh7LP
iUXXXCPxlV1E2c2KtVAyADLW+QjO2Pvdnqm9X16biMYtKBQGcKCwm/Un3eVk1w8M
D9OuFJVaGhsl993quOZ2k//FwHLPN4D5uuNfEgsY5KyIbSmdl2tqqg8GFGOLhCAB
G6eIZNXYtYDN8UAVO4Rcx+xgLmQy1j4AmRRXmuvEXYdMadqgWznjTsIrUDxqsM17
PeAX9CsZCJwz1wlyKEb0XSj81XFZsHPvJtAUEqMfJUgrgfOgtoSxSliVpB6/2Q9c
kvq6ZCWd6zeXABhCqfwmFviC1uWaDLkx3/za3qtwAlIZ3KPFs6P/WYguVv/2k0Wa
vW14W/GWADA//iNPCmy3wHWR+kbMrgPBP7Pb2dFABVZgud2CbOrsbz+d4W0IlHGn
9n1fjytrb6bDERLiVAsMuSLcHpVi5R5c+U4LHWRCq4JF01PfNf3sRYt6xw39OIZA
hGThCVhaqXghUnXMUMaZhLrXNl6QP0oFlmn4P8iskeAuXAcHtseN+s7jMxtQLwfV
INHuT/pcvzALJzOgXiNH/wvFQ+MGJ63Ntr0kbgM8Snxb/hiC/PqiidWsw/LFXya0
a1GcqbOpqKuav8RJZee9AGq8ulsIwtZGqwkA57Etwo7S12jdtDDABuuas2KxgXT5
webRfwyt0jS/plYvA5KWPXsk5WGUX/1zGzYk9erEWefjCMoI8AZKHoPMj0Lf0QRi
Sjk+VHtDuQzizyxH4HR6kHR55dYCpuQdNMLur+qqhAl8lB1+zcj5HEUMmuzMec3V
aijSbUGUhipCdBd487jkDhOjhnGdVc43htnQRL9qJjry8GjLx2U3Ptls6CKo3EGj
nhUosxwIKP9xFEe9WgToc7N6qaZAE049K3T/IKubZKy+9ZNMS6vT6gleFLi5cVnA
7q+1XKU0FhpqfMdu7z1DoNRmt1RoiKD+3yRfjktyTvNCOW/JCArqkmHmA7qSidNL
oFlZ1yIaIiAoYQQat9yvx9ElULWNu5woI2Zl087de/41dncP1FNsEovQPw0D49+Y
zzQEqA9vqjOnUJ2v4Egf60ClB0d4JUUzA43ns0WqzGlxwd1btnd0+F/WD9ElNlAP
WeY9pyWyw+AzVRj+AsW39OixGE2dGlGTje5HpEU1QxHWNIG4DGR/UXCA7mPCny2K
MfsUnf7TOZg+J9/La6aXKaZLsby66MMWlSwXfKwSNb5g6NGlTOYLjRttrBN/B1+o
Sm4Rm7NHpMDLa2Qr5R/9/NwTShvJbHp7rmFciFzQjWe8TWNgboi4uVVY1sdx9bZl
FyHP1WKP0SyUhnziDl5REzXG6BxaFZt6Q/8evuKO3R3pT/lEgpyVq/23V3uP0nBM
djlQaRo7m8WB0yjFMDAY1Yb+/+wTI2r790MDeC85r0R4bzK6o1KhH6PnwY3XBuX1
Oq+PSsa62wbjPM2flJrfqvH/YI0c4mfTxa0JRV+7OrGf3WZ2AiAgVG7ouy66ekks
B0HBkzxm+jG+xOgDSIAbl9GB7rK3H1rz1A/hnByjh2y1xzqt8qTj6Zfp0mdODn94
RVZmHTd7NXGvX75ClYIJu2+X5tWfeattPfypFadF4VY6Q2myE/EXIVaFxjdzOJpu
MmWnUzPKGRyGzaN5wGx/R00ecNSvgAAdxpq5c9UtYKOvL/azDkcxn5R/yNXfUTDb
+1VGolobaBwc4b5IDCESEA6oytd9Sisct7ad9SyDbtKfRq4L0YHYUAt9yDejDGS0
mNr9/YQungqMmKbn4IMMRw5KyNIs0J3tU1Jhp79lm7kWejs0pXyR3Em1p3LJpTuv
yJT6FhJtt0HIzDaJFwHOmyWZxZYPq8OFeuOSa9cTCL3Wnynv8n/5v6BOAFrhXjHo
Vpz0vv3oLd9HTs2mkPL0WVVpib11kMIIX9ed8Quf8maNtK/Rc+PW3lyU05FN+/oG
1/SN9szx+56EXh0nrjoygIiaPT4QFHyWgoZDKFp3vZ3DV+HvHr6Px40t2aB2JBsq
vKwYpn9i3feqnqH72QCNHmmC3NawzLvhlOSKMB3azvepWiwgGleCWonsEwezp10G
sGakgvDnLwUZJbcJZvUDy+2x2g+iWKebi88lzalfCzqfAlalfUsSFClv8O31VfVx
pUrJCVZvqZllkILxFrkIckkVUtzQIVAvDntQyerOxMPdVoD9EaNM981NihoWNVAS
pthE3sB8MaK5NDE5s40wn8HjuyAvhiZgm5HoXgdkLEp2FVidzImoc1jO5xwJwTMu
v+rmsX148yop4CqHoNgU6ew+deMCqWPOLGTjUAPV3avoFSts0qE8n49IiahuO561
QXNHtBXymxlytSdLfvVvxkO2T1kuZvmZJVX2+NlF9XF1qvrHhhX7ljRCQHrNvsM6
TU9/v2sH7KOIvLwiq13xL/hEeNh/77srlx1WZAfTSiTicZSBJguVkDypfYTkk5iX
jNSjN0dL8Em+v4LLe691OOUi0CpZHOAWFqXKWCKYAM4zTX3VFmhreQFMPerVZRSp
fN0Hs95wTdgkrCtgStntzek85hMrepnSnbhAft8J16wzHII+jUZP8RcprIH5uKyN
4huL0DZIYy4iKdaaua+N7jwP6RAECV3i9cvgjhJNFj0CaKw6h1cJmTVdSWFyE/K3
ejIC/aDBzXKc0vKPX/fuQnoF6C1ZlR+8n49zrTMwnE083KognpHBv9qYhsUrixXc
kizzs2Ysvkc8FX6U5q7iN50CpxxyBl8Xd8JMeOUGkTlyPT61RGSDSwGfPUnTz9V8
YkE8QE/bFXRDwBhlDZehrXDzrQiQmzmbRYYNEGevndyM2H/o5pDaJvlfpDdvMQDJ
0qkfg2V4YOtpADrKBA8Vi8yvz/17jcLWjTgsXrKgG6hgBx+I5OkUHp5+PVOnf+50
fSRcAUT20e/Tl7C3NudvqDHJXbo0C0z7bhnzAtlSAhJWufXQG+Hn7i3R790LSPrE
nEu7sjkH8P3LQ4PYk3CO2tHdjxrT24G0idfjupp1+ZgbjQDorgiTmxzFnDu1073v
zVFqBizKyhzR+th6LzE7sFKbaA0CPJWQTFNJFzMX1+fdCCRJauQa9wj7uWjlk60d
SbkR65rqRBPDiChFrHmf0WprBOj1rgei73C7gx+pyuShaf+Ma4u9OO84PwaPltja
IFmbn0HIgZ3sQ+CqvOmRqJ+YBiLSdgkli1WhIFGmB69FNBoYRJ4d1yHh9CMwRn5g
VAplaJMWIQUPf657i9H9bSXeharIVh5MbTr8S4hqgHY4oWR97Zy642YYWCu1yqol
Xs+nVsuq8WOOz0R3rwQQr760lXD0viwW+TKgu8Z2w715DGaAYzpv3C4DP6iSqcnT
i33a2p5Vu6kWuvAJzb9vhQAg5k3d7IjSeR5Vm3s48kdoURLXakMkhMyuI9fAYMLf
BdyCxZ89Ag0SbuVIQT9lIF3lHG/TVOpmz1iQpQKESs3J37gx2oGCxmqVQVTsgU4P
Ps9lLYs5hvRh7/EEfV0nm/lEqOVEH6VCgqSeTmPee3Ir/iFz/mBdqLsd9cdgZMb8
sKZtPKZRu9VBYw1N7DKyr8DrAfp+Q+WKr7yK6hIeowwq2CPS6+SDTr9PnShJZeYE
96L/W4ZWlODLFE+4NSzteZDlOnxB3olrAN4aAbVqcaA4QRz0QIuPMSY+Nz2Rl2ml
wBrhALFRt5NR89n5fDroOWtia3OYANCnQnsE5mUQ9pm1ds6u4XejiugcAHdVdR/E
EtWa7vnXOVPp/qUpoA+6OfjywJovi0QFlflRXeF9/CKFtVtijCzllnyt1lf2S/9V
dohCEC0SDeDYMl0NKbASIIElI5a406dbi1sdLxifu+1duJX0VfwZpL+Y62Vr6TSv
lMu5sQ1rDRbcU5JkaqGIbKBmxzrDO7Gla5rz93+Fb4rFSrlbpSyIDPxJ4xEfjbcm
xRy0mNnaMTs7+t3ydvN7iTha+goyduFdg+Rjdo2tTxA5qce9MfbyNYEaWhvyReXt
3MXEnt/ToJ21sdGoRcY22l6i1gMgSrl0OWZwwMU0glczsL2Ulu/p/wkCOcrDp/mG
XP5f1VQfTR53JRXdGCRBSlLmsgiEYCPnmrlOzktUHhBRfdXmADUm/nM9DaAhaC1+
bXvf3xJRYxJzBXuchRaFsrJ9IKRZZ2dWR9D3Eqc3uD50eQbOPQCbaeB80MI3FF7G
OQS4/L0PyIgHd1vwjSwryEBggUvoEfAFLt+PdUjFkMYotxFcyo2sdGyqEhLypZhD
tQ1ElmxT7nmGuNHCUVZyIdcj9qUYP0e/2pbKbmGA7/XbRI+smYlmIj/fAqB6ysi2
zqZUwcmGeXq27LvmdmgiSY7Lsl8T3oj0SGsMGtYhlQMgbWK1+APRJeBTSv3d84Mr
pTcBVEFrLUFsB0+CGW0XApv+ZjOkYIIdbyfjKCjY8DnLocvakKUC0tURKBngCTE5
BjI5xzdCVyR3giJ47iNr3bhj8VNi9T4Muwp5fdc+8UK3Z5sAvC/8QHd67soC0J+P
nVUhdmu/mq6rkiUMVBMICokThNUtB8wF32crf5g/LILgbXdmcKKdiwN1oMUPYB82
TSskWLEGkm9aN2iyupY2xBur5e7BlA4fhxKHNA1ggkQFkK8VtixMXKML2ptAyhkr
54YVhKWgJCeu34eMET67keBBqTUvzg4LuTunrDA6iIhHnt1I7A+EUY5WuNMHxCrP
JeHkUpZNMcwvid+b14FTVGob05idlAbVE8IVGur+SnT/a4h+Q7QY2XBg275nNv3z
nuiAYaDboPEOD43AdQD5TokAkYqNrtOQ5ckM9u6+nd9Fdtk/kDsOxEiterrRKrZK
0IpN4joAAbZNMhGKv3O8G78kksnta4oEtyIMkNYvp1SlIyIfVKECVZhtU+V4TnFh
8/uQYTsXVUonmUsqQ6wTFkLHkLa6Vu2Z35TDN4Bs6IbPgNyWGD5Rt+qq/OfE5HNH
2OFOmOFXXFCvj72Y1VS6mjdvkPyneWitsFtJuskuh/vLu7ua8OdyOyMZe9BfWCOa
xEG1q62JFd7zSY6FBITlb9usJbJe6bmMIEMzz9Zu2JC7TBd46VbGQwDML/+LyfgZ
hfvAYLX5XIeQpAeemA/u0GRwvwyCSnfOFhRCKrRruIa3861qIlZ+6mPVI2i+vqvg
ydC2pw9voTXg0XNlimoyKT1N6cJ4YmuGgKxkTFueQ4JahQTn6wdMLqBzQjx4YhX1
eTgmKL6HSkNt8smULgDcJ6Qrhl1cF6hIVt5sSoXbbtepitSS22hNuRN95rsgnZG2
qYI99BjbdrUBPkVyj+5NnX1oti3LONNWjyS2y8Jhzb0cuTidkeb+DRYD2ymGT+N7
zt6eMkMF9oVIjf0kFyA71flUh3wyQCvqvbXtJM/xbdQw2mOWLOu2FwXJWEPwLCAu
ytGUlb//480vEEJjPtvNvYBov2nFdaI39vmfCGsONv/30J5GkT7c4irRPtKKXyxY
hTFzC+XEYw7Z1FYZJfLqUPogwKaoNI+aeNkIpSgoKDmVp1GNFW3MhZsBrvfOJXy4
9NVQZWpmyhOZ6/DWGf7xdrUkpC+YiIWKBrnHacJEb2WqbFkbKYgChDsDuiTDmEZ+
mu6DHMOswT7d20t9q5TrdUy4ZSrFLg1YS7uW8SAHIlnJR15h9BFHcUgHr7wSFa4E
CkfdFhkoYIdCcjU78gj3BKBCMkgs2nwCH/BVoPwd0eA9yVtCLh8xQNgmkx+lduWq
BxK0ZB+1SKVMMnSSgxwGhH3TfQsr8AUV6u7riPOuXlCOky9BSrM2w+iUcLPMloiU
J8no6tzLbeR7BUH3VxegSfaRPKIDLfapOKQONQnncKFG8TENFzpjKZx8u5oFAYA6
C55JbJTh7VLX+X8/P9Xp+JaFeK5K2v5KG8Co5eNy6sfW7tbdih8jZ1aGyzlDBPjk
wv0OjRQNHMU20DUQLFvvae02tUQ1ls0DdfxuIfl7731Y8nvkOdAKDFdRrlBxOTye
PFZDLA/DXX5+Ew8VzcYE5OuVnwSi1HNp7DklCuH3S6OwmlGnJZn7p4sOBvCIjXOv
oiv2+IRVqad1intC17BadQln/FqjmLygnu1JQwG+Rx6p/U5gnSf3ZmkF5CXr8TVv
zCF1Bo0v+OsK2WiFWxHuKTG4fSiqsc8+VHge03utkOhhF47ms9T22+cDWpzgn7oM
a7hbLsi7P5Snttvj4Oo+Tdceotiue/KvThCMu93vaH4X10RVt1MRI3REAOws+Y2h
//W/uhw2lTSGb9L90AvH1z1egIPAw9qisWUh+iX2bIeyK0U0IZOKXnl+pFSZtRlO
ECLCNnlhVa+8DnKSDKd7qW/23ARSzME4f5JYhz8OIewHB37uD5V/1RwfRB6v6IPX
+7ol/DlhV8zmxmU9S8vQWZ4A8gTCFPAAUrUpMvx98jWOhkMVHUQtn99Ft+cFiFmi
zVKtbjCMCpkVmnW12782iMsTBHX6DLMu+CH7hl9IEbQ8Da7A387tjwH4u901oXVR
JOD+wvrLXMBu7JGeYOWBEPH3LBR/oAyFIXJIes+QOFMuej1RjOH+KhuL3n6Flflw
ueO9LaFpm2F+jntpuYhQ4p82CZBiynSlqdwHKItOBb+8Y8MkVg1JLcueZeFqSuKA
xwDAXnZBuZb0Afs6PRLVLXJHeUOexlAn17iZ1Iam24DvpOR05hiYyN1U+vtq8N0k
RCin6pnV3J3DTpvRVi2LOisAhwPvvrKmO8fbLKSEP4V8pdzs6FicZbs7LCM26tsK
KXfHz0/czuPt/z21kNj8yms7eh3O+zHn4I56muSxsXXTIg3kU33h827grhxVKNg7
3Qs7KS3emYvZkJf7LtiQCl/dTvb/fRYSAbzhMWKEFMASK9k9c5YoIV4HN0F3DiSP
VavVIh66aD4JHD+ll05T9y103AR3ZbJvyiu//T6utMiGNVTpmffoqvQOKOZHIvWv
diOZC+oweRfnttn2juxvTJb3OrEvu22N5ZkK7KsnH9OhMbZPX3hmkxdTGhbEBaP9
JXMkgYV67gkcV1hrpsMSgnuyO7eTc+URoOnwU2qoIsKNccAEh0QXdEOFJGzZfr42
Au5IUtQ0mocIrQzv6NmaQuuQi15E/0xTVgA6JUHDjf2xT/lKIVn1XWowcZx9bW7n
Q4LDbv4u2uVIH7wndcHv9mgQk4zVxfBTShkJfN4tF/AFlHS1hIsCF2EqJ9b+G/+d
koyyj8eEwNbXxQCO0TZ4kCJ7k7mUFJFhsZcP+0iup5eBDWuOijWaCJKqhKltetfm
X/zqBIMFzN9T7/2KVclErFOb1FWUjWGMA33YLrcLxxEs8wOTQgOa0aSK/2/g+r1h
RA5rtYqsCMF10oluXix+XqTyyl8MeWs9YGXW3c+TPb7aF4qzoVrquEqocubZE6mF
p+/WrNZ1ReWLqBwRZc4f4gFpZO84nib8LGZogOxtIcP5e9eAUAg50z+xUbS5Hlyy
Fuxdy/ihC/SJZQv1tdnvP4tAOr/w0mvv2AOeDfM0wyXbqJ5EX6ozBqRGXESWU5d8
ktNEJsUJlAQ2pQYy4BLObtDxsSi2tcFywvLcLtoQmRYMwC0heYspUqG/n7Rle7Lm
EJG4Ma52LLsMOjJ6t0Ngvqe288BsolBKJwlHicEsOg0RfFkWnBaZ6G+cELSTFwgm
iCteV4PP45Y3ztmKLnFDgNJvVP4W3HmeeUE/37X9SLuiJvU4VkIANrALDNVhx5Cr
TV08hBF+QnsVDK5WWRdIMWjO5EktCxMG5+U4nR6zG7pWsOZDc3md+f6m7ZgKuVMn
OCdivkbPJFPyyFa1QxrxtevTHzlzD0qAvQx1zV4/8+CzQPf8jwRBec7VcKjOXul0
VO2QFsCMEHqamuWudAuhbZ/FRfLZu0pErArFeDX33/mGdoXdAuUT7uiwTt03hX0X
N1vDpz+uBi+dOYlxoCSHo58ju/tZW+4fO/sEeX09TbbOTZaIoLgLJwYN/g1nF+KZ
ybVB1lL23h86p4UEKWUGR8fON/pfi8secJZaNL0oUFWlQMc3KiLcVUqJIbLuOFXv
vVieWVikrxHyzq93kmBXcHqmBehnfmHb7B4gd37lPTilOc0OLpZyIdiZSwJg9sW9
gECE9pQRoQBIao/dH2w2/r8HuDZuwKNeNSdLTDBEPG+olcWQk9gEXiOrXRfWOolS
9HakSRDdyOWLU/ZGbru8UmNxf3iL0oMbaoxTAjw2e+u2prw16em/1H+d0krgQLRw
cKpYvIP6wrPGCNfN+YDxGwsAKtcFbBJrixit+ytpnYvGyQF2+0tC0FgVONeqm1kg
2dynhSrl2pjmvBNxPqqZ2DtLz2AuoirrohwuZRJbY4u7J79zNuExnELr+wtJE14h
UgQ3bMXTRqyA/Xi36gfCozP3Qpo8R/fpbtRCP9//NeszPqA2jS9pyaN2wx5i340/
I0o1MWG8gUvjZyFVO6MkL0uePyPhyxz5gvymKaDpT9qnhluS87cu02F1jm0IjESm
PeQHJ3aNq4+dp56TU2aBxBRYQBIOqlJTNq2FRj5cesV6gNtxDNNkZlina48KdTGa
dAj0DqllyTz5NXdvtKSCbOClD3Ol7WYqnSKhC2Qxh9OfTIJKUufYIXzvXf6YWnqy
qUTkSkTQIscSXiqtZyRqTvo+w2V3mVbv6YKr+4TaufoipHooj3M16qUQJWiBYF6C
TTxHR354T4BRkjmpgTzS2ic2ycYi1bE7baNMkj6kn1/GJM6PFup4c/o3ywfTzBqN
IVpVMNBcpjjvQIoyatDoIfRAhCulsXjkhVbdwG584kyN1aLHJQPeidDNGR03zqA3
o1JJznq1/IDb3b3cCoci2+bmhuJArO9MtBBW5VaE/CFG/3PpFczjNvQbYldrJNnu
LrnVMjWOP6aVabj3+pSI4qmaMJEuihh91BO4FuPzNOF0QsjlZaRpPvSGZWOckqxH
B5X6h9CiCnKtgVCasYo92ramvqTvN6eAD/tXi/BvYciMkKddCk/syCgCucU3sDe1
WXlDcXia+sdUiIF82f8H2uRcx7CYgizybfqdNkhkUVaRnBoRwrYuZqbpDLgr7OMh
TZauqIY4ABxKq7s8c6SkJv2CXntzUr3V1Z7zghDI/aR+CED5+fgS2xS4RRh2x8cD
wzhTwcvN1ATeNDfC1ulzeeFRW4HRaMEXDOJ3Du+viKenk+hn7METES1gV+bhs/SR
T49arsTpemlk2fqk6QD9VTE/u0Paze2StESuSQOzTUs99B9yKchyVihsilfGLC3w
xiA+X8Exh5Vdc/yu6G50QGD9z5O6IVImuJfWEYsoiDhsy7cqRiOoPqk2/sRrp/in
bZKTdGf37p1yr5yWEaMwhtUWAnX+3wsH17Pwi9jXGvq7+QZaGbHhStDwVdavsUzz
qb/HkPYte2y125eZ6Akv3Qr9U42Wv6Y4Ee/iVy1UaYT66gXo7wjOL/weW5yPIDEu
J4NEYLz8cSPRvSHehLubSkYIv1b6JVAvZtJLPY6LnVIRn7UmY0nHRGDp2Hrx3t+B
aD1sLpk+/vZv/wU/VpbtMDvN4THTLTUCTYOLB3MFhEG0Sgl7F2PML339yjNAgN6a
yhKp4plRV0EPrBB9ePs8YsAwKwbniVtYPfJYz+oebN7Toy+FxhVAExxazyJuxkJZ
dNxETV368/XrX0+5GSnEXJIj4iBoWX7ICf8aBlk5h/SW4eb5tr/Z6PfgLmazjAXM
CyFuBMBkam23DKERH5b2y1zOm+iX6jwElUanIJo6yVTGdpL9O7LfiPLGH3F3eD/H
XVIF3PKKaW1pftYHHJnSHMdgZ+pvjKNQ+bHDIPO27QyFom3iRrEailUuAnx2SF0Q
9GXD2/TWQwFRcDCWdWpIiqp0zthjHl477u0f2YK79GzKFIPUvh4GPBM7z6giWBjh
Sjm+VE97wnlc+rdf8D7rx1X2KsUbE5UFs45GqzkzCC4mvhgI8tescyZrXQ+JJ/WL
kCbBUUZVHyXCyR0MRh/JxB4k56meITR3p7+a8NXb1N1/ko8JIcFC6YpfMGZftXH5
lPZb9QI7fM8XgmF/gXJt7C1dEO1k/LV9E8ZAaFmyPl4qQ35rrbkO+vKRhZUyyr2f
nsEXF3wHnhTWmEBlwpscIU3QJqxarMGYTWI9j6Djq93CR5jP++Ty+oM2z2VdBxNq
xofsuFByXbL2AEolsao1iBJaN8iW2fywz6dTl8RyUoDUMaoBTn7vnrdtAErWFyKq
Eq9ioYq7l9TzQuqcAlWjUtrvtfP4vgla4XPVl1/V6IaSnzhe6VkcLOXarN65zqO0
wsKPVxhfcKBMV+VPCkb+idUfm30y1KcOSIiq1Nqankh4U7YNrwp8+Z5AzoxOHVXA
eIsFN+LcahnelGWboWT5wyZQTpbMFG0lV5BMbnFlqL7NWONkp2hPsT0qb5kC0uhf
A+rFpaIIzOwFyPr9dLvPKK0I8OkEBReCgnEKXNZoE8Lf47OI96UbNlBGpvwS+e5d
Mu4xiT7cjse39aXLuZNBWJhWk6gV1C61+xDJCLf0GU8cQjBblCBO5VNewlyJXkXD
/fbJ6M4lM8YfHnZWKWTM0UZ+uSw1JsWg2WvQBoIhLwn8DgGPQaR1uSXQ8T0nSP0i
jkTEdsI+J400ALbE7Rp4+nNrV53uaW2U4no4ZyiBUKdptqI3B0hqMLGeqseSaGyV
/lGxGxY3xZ7hNwawHBlcxX/tO1qGS34N6FFhBlo0z7yE46KWLB6YXFouWrefDlfB
m4i6wsQWU/T2mkzdo+8GbjKHyiqmDHkHUbf4EcPb8G4ssS0MjAHF4ygWwRS0oCv1
KuyKAd4LO4/NtssqQZUQXLN42Ul3zvZgCUsiKjh1WsCj/rTzUuiakJINNEzX7LEm
7JcTyfPlSOuKDRxy5CPGlp82Piz0tZgF4CmQGqp6ja5+sqp+vRH6/BMn8zl9NFD0
GAoYLSJ/nIerJ23ASqKwYLg4ctOLrKQzT58AMNtFo5quZdCWG0wSNK6wl8AfHTaK
e1UqNo7Cp1qJd96fTenZTU1bNUwK7+k5IWD78CorAIc5sQ3dyjW/2xeqhrInR7eW
pIn3RrBqkBkauScb3xVxiVjvmNdev8A2RvY449xabbb7CZ7tUXkJa44ixsg9kgBv
aHXa2GHzy8qQDkx6LDXNdMXOGedSlmogY5l2sFeiQ3BpjwYVA8c2GkBiiKDDmmiU
9HQPWlwt34hA6OkfCu7Vv5PlkAMnf4qNcyw0ZRzuusv5xK3fBX38zs9KFee6jAl6
4S3P/GCHRQaBj1cOm9jQNLKp75Xhx9ZvuzHppKe5oCZzUKrutCflxNovuDV6u4wf
5ZA8/2SGRZFLBsD8rEFCnhdOpIfq5jd1EUW3gGcMZe2BJ+dc2wQ/titFoqE27VMV
aZFM4nBzoCVmMIGhtOzgs9inic223TLH4D8XUKpTUIdahDy8MaZqqcySKCQ1Msj5
f8NPVfvXJLGF9N6Ae23WIAKqW3Ow7BZyt9+bKaeFwyX6ZVUO4YnCCPed0d3nZ4/k
0N5WO88hM3YiDal7JRyKXsHPam7d5BSLAPX/IuudNad+dwNUygv470Ow4AhkJrLs
TEUli8UQTi44buvObFUhgzoXPwVIUbR0XsMkfDyKSRWoCpkiSSKe0K8vIPn1c2Aw
pNAaM8hb5goQQ4/mgrRqPxculqfBdpEnSXz/mNKmNzteUG0WRi2qZlI1xOuyw7bJ
axAqAtoaAUjq2G6wFITNjqIGF4aseF61SCyixpwQhOv7WBvLSqTrLhlYWI4VmyRG
Q57I2KYMYMWjHLc9FtCm9G2Dkf7RDP4wwIu2JXbrBqoQGOiwGjsT4i/cyiEvyWfC
c/7rNS7clAP+4t3bSCGjSGm+cbuB8S7rZa8vZNUwG5WNjjAcgfQravMRjEJYi+t3
ABtkdIMxWyFVfRgX0cMIzR7+uDqcFtWFt9TN41Zl8ZrOV03Gv/w/wtJq8njdGmfe
y+qQh0LWe41aGM9xTVm/TNW6ky+hYiwg9dFOLmdB2FKt9SXxH6i2kdcxsM+nImUo
dzP1GJ2pgilSvFkUS0pp3oRDuAx3YXMoW2dE5KUrniQlkIqp1FqsgS7CcjnGo7w9
tjrHWb9RijjiMZHZh3qPTDEJndKXI8fjZ3hmHuTS0E0qM05Fnia6F3Deo0CEpIF3
EC0rnWxs7hVHtWfFeOVaUaXXgi4oHJOCE+QaAPcLltaTUP1CK/2MBTfHiWfgiFuy
lf6mDnSdUA1Nnt7+6yWrIBuzIMddeM9ey0JoOr0vdR5J077iX61TaKkQdsNiBk58
A9eEsIkFtxlpkAbnbpHlVSh/daIuPfBbiUTHyImHhBj4aDqBKwzDv9ocRaJerFM5
0/d0xWfbKn3+a4yBI9Ijf1447u3ul+9Yho5fkSa0gO4JOhdWOUxH1SCwUwytWYEf
ENnc/Df8/2szUmcxrdpvxYQrT0maP55CN7Jj+Rm37KpFWNF87X5nqkLk+zOHS+XP
aCs6+zFXIo+HRQm9kc6ft/kkdpmFq8GXO1vay4zgoxuWs6Cdejk2VbJLLfYPvDib
EQPUT8s4Ajj8DKKnVyn/CM+2OQDxJGJS/Wp/mleY9ueILUbnRoRV2k+gNx2bZcVm
Kb88Xek7h/2OoewMBYa6X1EdT+YohGVLoxYIgfmfS7JdX8NF8OE5pMQzNoK49ffK
oYc379+541FgAFYWbzlKqjotXOoYaOZcRfk0od4HWwUqJ9mqJNb8FYZU+gLFD/gV
OspJwsX0nAuD9k3kLrjhsxgLTaGQb0KUEpr1j90Njnlv8eh+piZdN1+bmciF9qKx
LIid8kiVzmhMA8RJPCG/nqTBMgCQVSCsT7/+3/T828pfoF2EJyPfn7av3UdHn1pw
KFTOdjcPUadyR8NTX9f0Vh8XMfVyCch4lcn65J9xbdiR4tdnstJjPCMe9zgtjdXI
mB3roLTSTFZ2OjTOBFIvNct8x1CsNB/wn1exc6RI7mzJ7hiI5pUVSVWXXkCRM2Ll
yZqWNzWVK78nalrjeayw2GeixKAe23zGdjUEadY4wQ9AMIEYTxS2HYIKvAGd1k4A
Y7xwSuGtzRQXD5GzqqsjvFhWlzxqOb7ydFs4oNMEIyXeythrR3ltmr37GHrtDSef
j2/p4lNI8RxO8Njc22GFQtMMH5IGU4DjQ18cx1dblL6yIGF8Y07qoNdMwL5TSxg5
zXbe4lmdl4benDHDRkNL5MBdRrsZxs3+CQe151ftKC7Z6Xyu4EE+MDUagXhtQg5+
MI6ZqTBb90N5tYvxNgKU7s+RvPQC3KaOuSfI0lZzdZMNV3A/sEHJ9NTMaFzioEOR
gKzlzQxxpajHhLcMjDOEVkDz6nT7gV/yeOu7cuJrQDqU0vHZFC8u80J4k8t3Azqw
4fdJwahkhQBtAEsy9020+K8HkLseajfiX8FilG0qmGA/rEAC1kD0kMNG6Ia2tnt6
ZMADeOdfCAQnY9N9oY5TrByM5iIf/PUHZUm5z/UfGLRQN0SryJ0flffQeA7T3G2b
L55gurXImUFIbrT07roSQyu4dL8nQ6UJLLupQCE8kx82HDXzxDTf+CKJHGmeHT5G
zymty57bR1jdJeUPorMsvW65YGbbShNXbCs1m0E8uG0NNQPJkUgcC6G765Y+0sJW
IUoNkmVD446tAg1q909DU2d+fjSBMuxFaYOxTeusvvxuCFUDYSe7iHapXvd05PSw
qxvB/4hXHBI+NbNq3b7kBk60iDV4UO5AAJjrK6A/9cBFIPQYLqdDsdjc8hI8237o
BYD1wQMP0DfJ4aQJw5YODE9OinEScdI91gxW+rgiUeNklqfT/+GZw2eah8dmBrmX
h0jBEn9ryPSxLv0ksxG0BlV7XAtL+pLcI1nxsW7RoQZf1uupD8lLik8sLqHA7TgK
RzGQIYD8wjK/5CJHhxxxUJS5cjmjfD1yw/OT4Y8Kd8Rw85ehCjCs74539MjZYYm1
ZqYbiS+PtALAq1zGOdjgIZINzZFQGtRwYQYplW8nC1axzOEpTgLUx8c5Hfthw7Gm
r+7vDu3tjRj/OZxOc858FfOqcrxG0AwClInuaPx6xG51vPIaH27V5co+Dj05GkIO
Sq1lDzhFHKfl7bdbFPuPijTu9XHKG27DVag0rcTSyzzQYyY3XgUwBlzICFeU2xVZ
HC1/uBBMBBJ0uL3KBeAN6FhFRUDjW4l+sE+ft/0kOGhqDnrXNk3mbYiL1he3p6lq
z635PELlK0uhN0qmgtPjNsx4u4fBaJ3QA09VNXcckBdWjUYntzG05JjfN1MgKH4I
xtZugupOTEqWcmgvFnxU5Suz40HH4IQ534dSJIgNOXOLNpfA7v2NNqnNqohaJVTF
+E+3nYD023hqUK6ziHRTK8GNAzkk5aSvicIISimy2lHOwhNchFwekDGnTn8oC/Il
BEXk8QRbiqtNncVtddccJXvj5Oo+MC7JUkpJEzySW1eiyNTIcqql+iJ3dZxA19t1
O5P5ADvG9V6Uf/iubr0JhMupQQp9Oro8PMlGRyALFXl27te2ZsOx4lB4jIOFuEXU
fJ9qtEN5nDVpXIF3bRCIwZnhfHFT1OyVq/r2o9r5GtbmF3f4IbMzcyddJvx1JESS
BIHyMq++Upl45ACEPtV3vTG4kHvUXthyglc+AT5CTiYEIyTlz/a25Glvp+bl/f5q
Ztvm9jXyscbCXD3+mgcm1Ka4T2CkMpFL81RE8P85Uzo+oF1PZzgaWrgdRVTuYdsL
oXFchry9vAgyNd5Apiz39AV0X/7MYKIsSLkOom1TofvYutP45DIeOvwpgZDzGwlX
X78FUKg+cOXD0C23kkGt1Amdm9LergYylRFdP+qNVBnBTkcMcZgTNUsvRPMyNmb3
SkscQhi/JqTzj9NfS2EuDoNzN6N6YnnuzlouSPysgW3SxC4uNZqjKwpnpcWt/nzw
QsEokvFhBZt6U8lqLXkJ5tg7dq+8W5r+CqH9CPsUyCsSnXVA+2CwfEbHJMeFdEXi
ctnR+aNFtHwN+hQGpAenkMBehTWnNqsOwqKXFtHTOciYCWXYSFnyIhQvz784IVNX
NvWwbdJL+luYl6qd696F4SWnHbR7ImvSZpsqQgwI7Tdfvlje/R39Fbmn9QLHj5U1
JdUp0a7lSkxuxqDhTvtTRqhqmTOjlQVP+KE+jFGvS7HRqzLcfefA01DQla+kjT8E
09p9XGgxEuvrCi8SvJhKW7EUKZZslzJPMS4RZ3qtDfy5b07tUkVYshv3S4dsjKL0
E4wMjCDTdqpgYsQ67EgjjvuBHMPEJr24lyl3yokKOXqBpnw0YV+dcdFnJgVlsdKo
IuUnjomIdpitI1IhJU6Pzp57EVvJKoACpMvH7wopND59mDwKij4uHH/2ckhxYhyk
2UBZ8pdzbKleI1Xpysj4Di23pyK9scZ2zsTI2tQwPoDD/GE0yWo7OiJCpVSb2xuK
jivJAORf6+heWOh9Vo+fd0cEIVZBKQCOW4iViqgBKfug+ZkMg+qYntwtTmQeF49J
clGiOn3LJHdjfUe9yKdtWD7vAmIIH0r3e7A+zkFxfUYiAGyF1SjuE2Yd0CaPZdEw
5NaBRP3O8b4gc2xXfwumSNCI5uAxOYAMCro8CgcVj870Z2MTr+q2p6EMWWCyYFFN
L5CuGNn9yjf2WDXff0pHHOoXtkvI029TsLu5urfAP5iFEVbWky9eEZxBJovilQyZ
vN+j2DMdzc96Kkpd8JDBE5wZ/VQ/dXNa4Rmz/2b8hGue7TYziHP23ADxJITtLfXX
P2XIRrXiYt+2DF40u7nf5sIrRJ83vRDp/8qYTi8SXY1ojez/wlMR8/sBm8agPYlK
NMVrklovBk+k9jWGoMljuV9BvVVeubEp9ZTsPc6cwpInBlcu+6emF7N+0f3/5Z48
7Pp+FRgD3nvWFNqJ56KGas6No5cx9pUBLhSF4Tric7UYqVECrMVa8oD6QsPSRcPL
4U5Zlzlr7p5EKEoA8Fs8XnmGNe3KiNDrLDxY/lP/HjVeeSusNbvq9qsNnkVC0AyQ
8XN5LBGotb44Jw7x4xb5ZfDKuWdIeFimRp4xtaJAyDKd4yKZY4PwH6iPA0vFMN8S
DauWhnKzXFSR7ktN8FGhmG2wKOdpQuC3CAtDYTk2UwjpZoMP5XLrRW6bm7ITyDg2
RCTVolw0YDeepJ0REFuocj0NquB8B0lI/ouQ59n3e1negexL8gy5XsHT3goPBHlh
IIVS61CfmbKS2F6qG7BKz5AyPcHEGkdtgBCBkUSrSvw+Hf4X35L3JTOelPL4pgT4
ofWMu6dvRyARUUiiMx2e4Ru1zX5+fKzBK+2fl3aZQAp4g3r8L+PmNLABUTLJ/IE8
T/R6t5zmskvEHKVMIa2UV+VACW02thXvcw1Y3RS3AIwHO74Hlx0mg13YILG9/7dK
phZFj3AA5+Jitco+Xno3+iKl8Jr4FRjvQbS1lXIDWr2UNYyx8HK+e2qUFmo79giU
2zFDi/wmehlBa3je+LAub/m6bCb66n1Z1iC51fyRRQ5qrDS9FX5J0UBYjqR5TDl0
7yuw9/Dd+3V9x2i8mhP4OfahlW3L05azjYKdCrx58NgIkQfbQYuqUep92z/n6nML
piyA2Q0IG1jowvkr2d8WHpxtdyL5/nDncMiiSWRKlhhvAXnV8my9ONaDU588m8+s
Ne89o9F+D5jyHaLuz5q9rKrE7VNdpYXu+x8vkz+3GHPDIAP349DsYFkRdTSXKpl5
eRVN7LTT6DUWCO56fNmRlBLOtMVHX/VFCWdtQPeQJYzz0jyYbiANjqMK9FwXraMD
xte1MsXEyI0jwf0Qz5fxiIXQShqI90HoQSfFyLunHUOcJ6hkR6o0VA8/m8RzcyNB
PiiTtD23paAp1iTB26Plj2ouQ+rCNAi5C1a3/htcXY3o8Ad8CXzE6SNDdGbYGIjH
zc8TFRi+OYVdfCF11sY/kT8CvXeBVc1OndUOQoXuB++TK1Y8fe9wXXsniDbRsG/z
BlD5lkhPtEV1u7mkImt5lN0BU0lOqdB9iuRsY43+8uLW1prhA8VnGkhJQALaKUWv
4lp0PmhA6jUxL8nlsLDMw7smp9uBBDTX+WglE8do6Gj+LICMXSQ0cc67pCSDsoV0
kCk/HJA6UQHuNU+NVKd5P3t2gHyGcL9qcD8PLs1WVxgTh5WAfXSONB6VJpmKjzkB
3hdvy/GL+KJlQkUAQ0+QhM/tGlLD0zXuHuChAXCsobHPIGlbsEQmFdz01svCwGo+
WatFgxXv6qPJ1z4OI9q/9MtffGS8fiGDZIHKVMhnIhaLQS+pmSW+KWzu1he1GrKd
17ogNxAq0srE968/DYYLigpWPJVvCZwv875EDQ5vTufzX0QzLXEDD/7vKuX3uQBs
2yHgBubEZ0vvvV3/Ia45FXmWfTrMaRDEbJNsIVbqV6UIN36awMJOINY/Nq0/5N0R
xMHgvc0hiLF+SzGUYdmcIHZFk7pTgOB+tzkowqShEsjcohx+1Y/gg49btE4XalpO
7aYr+tfCVmNsIqLHPSpdpcKSpsLqz5ybxhc1ZODXSbsydq9kLzLj3yGqgK9KX0/n
wzERt8yiqsdHRTDo9GhSuMFzwim1DfHsCnT7PviJVc/icvufduRZIglhkbKtEHJb
mSxz74NdvPfuEs1ypaAiH+rjfHyCgL5sfoFpr26BMEtGwphjh4fJMC788+0Ma9nD
xm3ycOOGsddI7eaqkiav2ucnc5PgkXHNolr8464hcawZz9d1YQXuNKPqAEH8qx1C
0MQ6SZ4yLWENQk+qUECHmFQGWpcXr2YZHDBaYvrVSoVAdapMVQ4R2WGi7q9ARlXn
25oIna0QcDyzL5hDP5T7N1r561hb7QW+sxkGiNgYeWYZGCLuc4sc7f4IQIMfXllt
Ktp1BHvtCPa3rZKq3y7HoEULv8r6euBKiY1Dba092L9ztoogHKGTNPt4fv5/Dxe6
nxez6I4EsXzef81HfQHMG4Ae7/UIGaZAttZN+IDtoigLxasRPTJ2xqIbB//eIX6t
ZkCPgXrPsN+6Tn6Vav87oDQR0vN1I8oLLE9qCQ0rW/VmQNDxCPaHtvGjqFWY/sf5
K8ztWQvi+u+Jy/x2rwdcm9VlPQDNiiTVh0/0hPWwyszYEgaXxXwTaPq1Hn8NkwbK
sBgLFcCELLucu8lKsNbPAch+ZxRn4Gad5NW52zqFl6zsRJV09VldCQ843zx1tW+j
4AOExRwMVzmOLXbXm7ViPRFmkeIp7xOKbyhQKnafdRP+eFjAEWG74zXhWHTu7Ex9
WVwrSEo2gktEcOIzf5hDAATmKw1+vjTt/t9UxBN+c9ZLa+UegD5upaG6QoT7swMm
bD9P/dMfYzbZp0YAKBWQmFQMnrZn75M6kOKP2eLt3jwwoInB8PKyLS8JPsInOVH9
Qa3+30fUHzSe89Csch37naUj1EUf+RcYjT4c/FU/NSrXMC+KFLyjkQY/iN1eTog5
DSQFBQZc1DsYdmkKwPVZYcA4TPHJTUjsMFta2Nsqo/RwIqmx5Fb0LIcKbjR7gveW
BCVMdWmDzbADUwfmFreAFvEVgY/ixIxeCVctMpTWa7t1oiOugG5gQJ0gzIRmsmq3
jF3h1gD7+amouxg8pD1XhQs4UbV4yTL+Jkk1/TM6eaY/UV/kaKAPqIWn5oSaMbdq
xzgHiR7QPW9lH82w99deBeWqKhNU9HE/YcQJnZqRrzrF1pQeo76Z6dsWYllOijnC
ZZpHxO05nMctrMHiYWfBMlCdHQiDlO3C+oSaSanDA4ZEVLr2KOlRWz2/7O2/22Hm
l0pJNrVh8gk4koloIbRXiO4QJJIawuUjC8WsWmlQLwe5VsPTNthAzf/BGi5eixMx
CRGf15rc0Pnsk81YnWXTB80QVVAjoRPna2xqGaauGdB0NddwLG0VV/nMWJJUCPQU
Pjn0S2DgqePM7HEE4qz5mpMIlB1ddjf2mTp3TnuVTglnhe0oG2/6ou9oSkRnozuE
E+Ku4Y/7Go8DXYbkRW3fUf9y7ddcJ3s0DCqe+E1NAq7ZplANyNYZ2cnh8eKNScuR
6MoE7RX5wLkIAwb9kauTXREXy0TJvWh34UNC1GLq1naQ/k47wiFFGMObBCZWk3wn
wTcQlUt5DvcKGKKC6ncPllsh9rjKk9YIBDwdEEoxuv+458QAdRlAhUQgVI3tOH3g
MqfQvfPKh85KWu2pX0MgDn7QwqVuDsvt5eLbUUSPkrtl0RXUML5pzGt5CxLee4nA
sKeEOh+bK+qADFejiuEJI6WmSi3WtXcf1xSdzgt5XmRbfebWxpaMM9b/m/L9hUGI
wk7Np94/ZNm24dR8J+FDFc+1MaVPzR5IdmOozZUrmeIlEmvY8xEwKesAVm9kj9SC
Hwgq5/cburnVkKDkaFrLWXuB5TFHx1AisrJJ9UPdTJF8A7TD4SJAzGAGuJzTGXHK
aH/y7e4ScW7igr4Zmq4NYupRCD9g2y+jpQEpWbTmJCtcIvPFNmkr9eW5Gm8RItkT
NWp48Ztl0exkz32LT0u4Tw4gWHujWriKK4Gz8C7HlVBFPBlIZJakzQSsi3NVgVL5
gZVDnDU37164PAjAmt4Wzt1mhPecXxrCvu19QvioTSiHsBWmwRyxu8nTGkJxa5P/
PnkCsClPPLMUOqHHkhVPnK5OvhLO2u97+cXtqMr0d2bfHCAKsqbWjkvC09candNq
heSyOjuckXEaytt0YwFuKWSAJdXs9Gubwhx1W5uop+U7xaCAwaF4khQGUmQj60x9
T+h3WiYOtWefNZ4XuaVfe8zefzqBloZaAzAnLYIDXmwsznmx+q1DHj/Dr+syLnjl
vMHNxmFL1p8QBK/qbQluQ5ZHX6exWyrhQechuhd5J2fmWuu6YHWo2X0ELBWsfOU1
x/2Tc24du0rK915zqQpsLbaCjRHJrKEWAlFFga9svEvk4VsEehgsv8g+XN6kH3mA
/PFt4XFBE/NaILQJ75FS4DLiA26jgEf9Yumsu9D1OycF0xY3dhI44Jw8uxFfNfBk
SJpUVetY5Mv2cpThJAEQuYqZL9sPReGJmnpIUQmDRZLHV9Tw+McIHTOgqt9Godtf
pXQd0XlsgS1YZInbSMdcHkvgG9THPckYNCC8loQeUyht5570VF0vmhHRwhGyeOTm
TupOhhN7Km2ovB6hPhWNf6aV4gjeZy5q2CFS+WRv6jbO46dZK42ZIeca+nXW5yq6
JIVe7UJSQPuJNgbedB14e9Dua8NdvJl8KHWBGIlIR3/QM+Z/+Q9ITqZ49hZVSmC3
uCGaSoHLYCiQIvgftejjw4KZ4F60WhHsvAES8Wa3mARJmQL5ejyM2p9MqgZUZm/3
IPb/ZvecERRi2DBzMWz0MrIPaadG32fBuCj2vi4JdOnikhRKLmk5BWwn8H9bcR0e
yjntk93eeEpifl2kdH+bPirX5oRfPFuu0iav4Fh23rG+A0in/sDtdPoPo/lCaodD
gs9kSCS7jAEJp8O7EwtLx2d6+lZ+6ImoBYOhZxoR29fV/uJrsnqU/cAkwC1lOXhW
nlxRuHPcIVCJfAakLDn9MQ1mAH9+7AkKbtnhSd8M8AJnPCyIfgGBUf9hFwKXB3/C
N8MxtSHIX7NC1G+/8ZJ6t4sy8/BWmJFSJz8Xssa98ZCBPWmwLLiS3RlVxdt6VHOs
KJ04PKbV0m8Pt35lki+pSsuTritrenWA1LeSPoMVgLAHbrUl12RrBi0dswMTzSX0
IdtfjCogPzfH57RO7LGTSRVA+KPqFCm3fYMEPvktt3yL6pF+dnyJUa6AVbfAassY
h7CpYsOUB7FaufVnX8rr92U1erJR5qJbGYx0dnBfFXs/zxH9OQhaKR8PoXsyFGZJ
9bjfAyq6baZYbGpTLu8+OPHppGoY+zNVcpV3HaOzv+frjnvTaLUpCeGEdhQ4wouT
kbep+VOZptZYDHqvPagLpRPC0KP5dEr/oe1eNULw9QFRrgFIpuSWOf2xnF2qLTV7
MygU64dpsLmAHk3EJDUxtUMlCAoprUQpkFof+u/GSzhu/G4ycp/32OuCZYTCPxxf
zgxEmj4jue8wlI8D42rEd1svuLDt2FRIylg1vXlokTRUpXKVxKrZB5dNc4j3sQ+K
LFLRaL6EKP1aBN6V72eAp4kCNG9B2ex7/K7kNHLujcctvJV8G6yhU8IV+i6y+zRm
iuzX2EdCz0iiB8x8dRpjr7a8HoxtL6+ydgMHWH2zpL62hnAXISNcNdar0cP12avX
W+nSxolhG6+WRJctVRwCTTllefMW97knZQIctRzGRuWJLxmoOYg7o00wXDzIJTCC
Zt2AqLKTWfFaTAMfPEwhy8eTlLTt6GPstF0BJrUme+xRmFAZgUVhaEoI0MxhOjlg
IOG0IlaNIK2N6FUl2W7cLqT6vcVRK8XEqVcMHh9qUyFEfakvhIexBjis+GrC3WCO
zndGRhy4xxQ0iEHQIsMPsrPfKtjVlvRK6amS8DpQi6lQRoQWZl6KJXV3Pmc+GIjh
PBKQ9lPCtw3/rmZ8HGR3WAagOQzCZ4IQ0vnDGNpoNhyzkTYH+TPEZQeJnQFfJdiP
MrE4eGeiBhZ/eUiFhs9Y+y3CYzIiIn2Y/j4ex0QImeVhGXMdBj0G9yHSr0Ee9UFV
jh5BuRJ/aJrtJjt+E3qMCsXu0bkflr432EOdoEmruipq/7kXpv0r5MgypSqctCck
1xC+/41MA3iM8hqmI7KXG/5wP/5yizzJ88xfRVXxGlA3wa9JgxKjh5bt895kArxF
4JL3lzRriU/vYNCFkZJMOypLq2mhBcJbXa0yNpR8zDG+MjTZQhAnQVvxX2grhDgP
fd1Fx3fxAZrcMIlk6yajinlWbcEeVuzhUKFFHyYyvs7FZqDWjOLZfr0SrCrQlY2m
XGUdE+Dy9wegcvSd3CEMln+lML22VE7KgSTBFq6UTlWOgQ/C63eSREeaSfev5R2U
8IsgrP9NBe2mgnrTAHfoaR+oBiu25i9noDkIgCSpAB+jGzLZSF6AVCD3LxVmq07R
nFsiy+z3za9/ImNM/8Mujh0eMRVhijDNJxIn4NBCqAE23Stt2MGCG8PkM9hcWFih
t2ioPzxvcS4iBVHvqRWHCAV0kp0eO30If5GcHJ5EAoGkUb6j+rNO44jlzlQbFn0a
iBbBngtlquIeVirE+11WjxSOEi+/kWOnNXU+SuYCcWbt1V3rBvSzU7P0mou2uts7
x9e1nn4XcaShjYWdapdJ3B4mIqDjjqQHBJCgk7Dq+XhCkT5SwFNvqaRDs+N2W2Xd
PcVuixTbye1GM48AOGu4bi/YwH2I7Y8VwMdpFsQEuxAiJEmugOGG1ew9UJzgzTE1
Y3Jo8tEE9fyRIengoH8Jqdt3AweZlSpNOcPuYE+djnfT3K79ANmi4iwm95f+NVKW
E1Aaqiw1T1+/gKWMNNDg1uxdZ0Zg5HBWqkaHhJxNnjCdfDmwuw/kClcBBQxWgy3q
Vim+R72IIYfnMQxGhsS7ZkTdBJmUCHeowNxFuAWkunw2JshHBphAhfPKUtLxY+OF
G5JIRMDXJssgl5SeKb7PDPEvTdLJL4GdGKc0maRaosOQSVPp8onqRg9+SdryMxZM
SxJvp6PsBKLeMF4KEeBsdQqwfMSAno6FZ7W1a30ut8vKlG/uVT0rbvjXXIBActaR
G3jB4rYwZuSCB735QLrfcm2UkmKnIQ0lHM/QsQYMjETjMMturnimlp5XtpfOawXT
C5WZCAQ+dd2kphEt8rKbbcS9nvET8mK1mFj+zTtuL/7thALdBysWleeJbfdVYAsE
R/4bN3K3sVQgtVi3UC7zuLW46rMDuYUycYKaihLJkjnhrPdQLjKARpCJ384QzgyZ
0NKJnSWcEp7oVX08Wf8fzfDUy2FLl37fznf8s7bfT2NBBBXY5BXrTro0+KSom9h6
tIleXkH80SshZ6SSmZIYUnMwnoxxcq33D1rZJ9oBz+7Bm/CT6Z/DrKkn8hDNwDPt
Jote/3BDRT62XR99G77GIV9uZpK9MXLkKAxsrJdTa862fhc+VFu9+d2DdaYE+Zwt
XtMTiihXq4Y3dqVgEyJZ6835zEaM+BOcBE3hjue2u+LPrfcrKgdVPRzSJyPS0X4m
iEL5X67942q7acH5LDAV3fJURomismLJdIJfbxR17YtMJL6ZalVvd483T4xrv94H
H4MdBjJHmIgk3OKWbgt9kosOZwzhNEiWSkm8EW9ypzMymb4nXy1s6QV7pyfGV3lW
TQTzxeeAnxB3zyi6DXCK05wfZYGK7kIzCv/zA2GdSvJFQXZ6hwCu0Ekj7Rx59SZU
/1j5ROVYJC8yG9VX7vBZCx8QrOUfpexWfAzXSS9LtFXUU2lvCZrG6/EwbN0mz3gp
QvO6G4g77KFExK5GOoGI+1S2BBU2uXCepKGgCk3ZpZAwcvo7lcv5E+s9nMQUzbtU
8LsGePv6N5DVdv+oOptzUbGebxUA/oVZnENVOVkLRhb8UdDEB4rX6eCV5ify/6Y7
DFYdY6fMn4ykgM6492HQSllmfNM1W86KfuiGrmNMqxtqWlSgNNjJu30WuKiM83uI
SDQwEZD88BYn0MjggXLGbcDBUNDM/txZ6yIvqnVkiDnGPjCd9/w+hvhfywVBwWim
SExXEBKy3aW2N9GkLssgypQIcM2R8YxCntgij1WRu/0IwUDFUlpvlfpraneD5SbW
8WapTwUZcifPcOH58MrFx2GwatkEiHrXMoZm7M4JeWlhjBBsLaKi4e23DUInr9PU
ZexE7TWoMbUjYcC3H9W+SC7F64T9gSERgndmPEoycgsfdSnEpuU4INBcKsWXrq+T
oMWaXQAuNZOxSmsLg0uQRrtZJE0HHvYiNxDO3jrMOfQAdcMiqFC39QM5YFUtFip/
5AZg7RAmSDEpZ5pY0qYPAImKZk3emf3FHm3dKTMZMb/VkWLqONe21yv7TNtZ+ZE5
rlUDjL5QIK38FFeJMV9Z0YOMACN19Hs/rx/G/AaXKJJQTEeV3gE8kD8GE2tCMgxW
+0UBa6zwZKB9AmYaBVkLpRGhhCAEr9r+G9b3lfSCw1Ok4uz/Mp36xDTEwe5Dk4oA
pBb9JDcgeXlGy/MIwxVIiC9+VltPwMijMqXFIIydb9IngnpZ1uHTPKcHmJ7/tLq6
8RYDxffihEsGHxTDX5SOMoUg2ti99VQ/c89DlgA6iSFTZIp1OgDSMSz6BxVFleEF
Fqit99XrViA0yNmz0zGmB2I3soAKvRFwWyX7dQavct3zn4wsMXzx7e+kOyaEX81X
H6oaDr/rkAxY6VD/Oaan90a6n1npatd4KUVZ0uMCYY244LG/ygL8tPY7iNpN8syy
EBqCNQ7HtF8bzneD8Yf/tuDMtxlmh5m/Oaq4Aj0WjTqoc/t0NHPkndnSo75l36En
rBGj4NTKEIQHS5WiE4e/0f5eyVdlIJWI1J5WAtVRE4kiF5BeX9Q0n6s9wW8YaP2d
nnmFp5eV8bjqp8/iqq+BcR4OzBtKLiQQJvKi6fPM/iGyveEtlF8i3GxwHoWZRw0M
MJcyWd3cFvpXbNZQi83W7UL3sDSsc+OJ2QQPmpO1IWaLMsOK6HcqPGKjW9vzmMBn
VhU1Nnk5BvQmdZ98y0yO4xbLjGfdFO840nkPhtYv2eNObTPD6mcNxptzeZXJJ/Vi
J7U1drBhug+VMMAtkwnnLbZCq1Fg9ZPXc2g801cgrE2/PAqLDTnC3L59Y0vcNDRA
tre5YsN0ayzA6HP+MzgUAzpQmMkPVS64m7boqYfSLUd6yNfD2adm/0Kqzk+dIek7
HNcqMy0GWSGB/OnnpLLQQuu7mYEAnRhNkiM7zwQL9UU+kiBG+P5f0X5Vtbp2Psf7
0Wztmuh2BaFFy3Wf0FPbKwMUBr1RS5/6GZEeo3vkyrGmvfYefGm9nDDLXmQcU+VV
Vt+UY9DmuNLTMDn6qsb5ag3MCpJ9sR40b9rHIjEUf+HnzXJ1BV536b225Xza4hj4
Ha8f9JCaNS/JIheN8+rXPAIHCK7aYYnmZv61bIibjCy+EKPy02RMMFceFN5LrgvT
pf/hKpZjtS+x0oFMWrfpccOY1QTQAOlztmF3YFRR6BFQYjr0QsiUcth+mDqygpOL
OZEbLmK/uzQy6fu+9LdqS0COm4STma8xG32CnK/NKxSzu1U4WlyU4KmNiuhZKSkP
Fr4C6e+E9WCyMN/F2qm1JAfBL4XZcc/Z9A8uIGZ1NR6bD6HghDC6cEEwguXeLOq+
l6JItWKoY7so4a+XLPDcU9GSebcuP0zB8hW20boW/19rFiOkvLeCOfMUbZnnVpGB
t02P0IkUzn2QDiEMF89zmMv9L/ClGdG7VFyewDh9HyNAOfJiLJwGBgzehFtSLlWn
ZDPlX6PafSb2+RGrw39WeYFS8YY5gmUogE5iL1vL9z7zvzTONdVimmJ9q9wkiG7T
/G0x2FkU9qf01i/A/jlaj6Q8XRiWasFqnLoiRA/yJnM5ArjQWUL/JAW1ly4xBDUX
g23JUzj/9tggN/PMQ69KUNSBu/Dhe3SzPj0NA9lGWpc/g5hFQFZ+dKqaMLyWyAGT
qyGXQAUH8vTid7+ok1iJu2BJvrOVbgZG9I7r9qmRuBZxP419OkTU6z+EiXkveOBI
dvzIHNttfuiDvdlrZk5ewFdUdsdsWOOJGeKtwzOztBhcl/GXOuT8ndJdwn/HB/K9
XQidvbbkU1UmWdtIL/jhw4y2PBU3/jo3TbsKBj99VQy2v1Ccd1hKnGDhosNd6+Fn
/b5wDE2KjAXH1Jz14Q7k2IkuvdQy+g26fhrCL3wvF19JRqpSCjY1Tk4Vjgs4TCt0
ypCKI6xGxzP4kCJdbppGnA42uHqYO7Z5Y96iAPsPT7LfAHeuVZD7KkS/H5/wsVVQ
+rVuQIAF1UsR0L1prACBajvnaLHlCMlkflJGGSLguCY9bMPdMCvfX8713U/Go0s5
HuGjJLGZzWuuKfPT1EU8mjBXKuzgDwdTnhuSpkfj3Rffotr9HqLr3x22StqdPcNX
jfz3DPedp+Nxh/H23liaovIn7uoBjEobT35gEUZ5htNZf7HxHjh6rcGLha5V1nTF
57Ak8oHAo2dKVYm3tW90tFvBoIu1WsK8rLAKDpz9D2vJE4bA6mBZDFBLAZeesXQm
iYyEZwrenvpvU3ZojMSrtWXFZB4OrmdTBvJM5d5iD+u+SqdWIvyKZfgq6ZTGdevv
Ry9uPlqum02vmRQsKE/1haweAXq6X9OZhEw9zJUrgJc7RU9owXvxKLhQzACj7qWj
cXQw+OFo+EwZJPyrHsfvfp9++W/gZcktpK08o80tvbUQbHZUkmr3jzydmkvj+j4H
zrpvHCtcShXAoPabHf/9h2Ee3TjxLOBQthxPSasv2yeDUkLzk3iJIMezMY4YCuLZ
7EGrn868YSSeNINTXiDSL4r70wu3mdbnb1jdlzVuF/eLF1HQA9vUNhdVPlY48giA
Zmvg40QTc6GUCut48F8FV2WDV+q6wQBJHwQng1p+a7yy/9cNa9JXeaTUqwLm4kJ3
Dv1IrgyKDl3sRjPaS2AbmRaUhfYEUx/3ecJJ0v+DS8wD2yz1Qqe9056ZbVMBB8b0
NdKl0FCZZZ2aj8DwmlA/1MbS0cv+moqlDPJUmU9vGzVAiw8TgScq8AUb0GqEgzoR
k7hv/jptY0IOPbfJigUZG7d/wrWzphdqVjDZMb5BnWM8rlrCislgEKDvm6H17syX
g4SK3aZunUZ6ZB9WLZKOuQjv15ubiz2I60KkJzxC2nfWP/CFzgd6H7FdcNTEt1Xy
ZCMXR9mycdKvZV5h6v1PdYTlIhO0MbLRbqYH0lewUfyWfeiYL6MroM9zV3HVz8tl
ewkqTCrrA06e7CVRUz8HFe+sqyA4aIBXZh35qrD+pw+uFmwer/WXqQ5+8SGANutK
B47Nnt/KJJQHnAIzarAr3OBhfrW86VjkvVJPcHEs2GiZYeoLfawXS8DOjwKLRp3U
qTHYBt/r798YSXaWj0nwtAWqic3cOpczCHTP9MlqFKn0Ji7d9dVyOUfFlF56ELoN
cgaZqN/wbSp4FUG5FLM4FgOB03rTvgWkqmB2FnR7Xzw2IG6E0pG5jhWeVYUn3FGA
nXe6pXTHKLMQbOTRnEsUVzlTwbRUz/uaCUVB0KJXreMhBEAFk20/i+0mhRv85Q5l
4Lu/cEizc4vHI9gTeYayEeiId8aNQ0asTJznrs8MUr6hBaQsaZW98EE/VnSL2fbc
twALWA8kLE3Yp3iQgWeREbb7GMpSKp8FeRwLgwqBYqM9MQTsYUKh3dMfqw/Tgtgc
rJGd0Y1LWoKoK2HWe6YcYqBh/+dlhAajNGVita0NiuzKjbpPjM4f3bWJ5KwM8HRB
oJ46pnP7fiDxFPp1RgKmzPp16+MDNRF1e1e8C7qnZQ9ix23ybo1oq7XncC8+5fkM
rpz2MhHTfyAbuIuKdlX5xREIagTWBBywTcZsj/9Dppu8bDFqXB2j6kRySxv+K+uH
BrXUbvanIXEFKNsYICXR7KTLCPpDAgfhLfgEAGJhsTv23vNoVw3XguKZ1OyT5NBP
wM/47Os4uZZdhIJyneEyQVNOC82ihGexMjYChEPhMq6KH2bs9RAdyELDhaulGftN
walRg3kUlXqcRE2eXs4ijXv0AMNzWsq8QHzcMaT/qI4YxxSlDi0P4DoiTaLA3b2l
qFYURoDUNginhNdrZPzgo3ztv4lq6PuH7LSWBahQzcWxhlBNDX70KOEBXig4vXHh
zoO1trimLYXbvyl+H6wwL8AN8OkYFI8dC87rHmsAul57gCnrYAPo0zafQplTzLEZ
HZHn7PKhAPLH8L3za0N1cLVcTEm6Pl2SeU1b8zI1tikEUKmO77izXqoGXguyeGBI
Z7ctjlULfSuyM4t0ZaDXVflNdtMr4SjNvyjb8meIQcVothUhtOciVKmeYA44gq+d
LJ+suJyZoWzZerQxieOzmXIoC9czTnGUEa5ji6Yl68A9ytbgS7q18nvt0ll9ElLq
e3JiD0dUjXqefDiudAHOsWeK5yKV3Mbd8sMVoHkeg9uTMu2vdOgkGuxFugreVqeJ
4iIuFe5fQP3tqCd3nvdDhyZD6QgikoxxgFo6LJzNxQVCcK3Q9f7hdNtV3G0Ju3b8
sC4R/vQ9zGw7Jb31VFfysokFmhVGlrsHCljQ8vYZogD+08f8hDcd0HVoPdeuazWU
bCMy4c8ZCcd4rRQ3lXfyDk/SES0y23OXY9BVlKUHlK4NbLputbT0uXKW6CeziRP4
xYWKZxLfsiFsuUu55nYgT8fUz4HVYfNhicSOb0o/Kjyi+4DqVwT9DyJ9bTeaOyyo
ZzfB7eYYu8HXWG3OSlGLbthl8xdyrkS2Bf9t64bhGdK9LhGULCDlhnUxkx0UIF+M
czTcfbiixBC8CKe8oB4XcaTVjf00WQAfqR88bExBeE3iK3Ea1nVuYGTXor5jHVg9
LKLvaGpqGWsR/aNeMAdb4/+AuZf/8Lf3vmImfCo5DEICWFIElzIkDXF/cIU2T/n3
LaWIgpEDWZXBuQ6ExgT5rYYu0+JR8DdGg86NHoOVdzrS8odpoJfWOt9redHIfo8t
7amCsmJd9daswjUTYIenFsQtabMVcMA6s1A0uFAVivTmbeUhAcQLlAiVBloIK4Eu
U3QQMkV/UfZ3AyhFdjtBjeFb6+ZNP/qhYky0V89OIeB/qf/C6cRRaplGLQuf7c5v
2WKZerV7kIznMQoPL5shkYsvA+3mgOEYM0RgoOrAG8w+14oDLWcJOXHBJpNAI4Vt
rg4S++lawW9UP9xitDHnlxqKpt+MiZQYCM4SdKjpIqWmtmcxh5jJgFDGeeDbp/un
GOz8b6+orr7jFsJQWYOTl1co3jp0Rw6ddCtjCTvJ0Vy2zrGzgOC4tZDjU0pf9/Wo
6MtizYYBnroPHa1glz8yco3oHp2HbcUjiNkHkYMYoqjof9jqgL4jT8teWLpvyAje
MwrnN/Ww1AqOpeTNbQxwjVaevEdblqduoVMGl7LMDcy1ICag9XS3AWwmkInk3aJn
+s3qFlkJF8sKj4ElOLnBPvqHvOZlA3rGiaHFBB1TiUnm4LuW6bV33SUaLFHJQ48Q
3dPXCps1bblfZ/p4AujZJmefXiCzM4a29ew/OBn0A6IQqNgjM0FX4J/qVcgih36q
qoGA4ZwCcXcJm2NhbRT+GMHQqXzqZkPlwmopi3Q3oTF0zir06Wp+q/4VzsX8Z4vR
CX2wrha8oITTK7cNtdWnyhp1N3WFc22JaiiP6cKVosZPFYw5rnWuFTUw9BFPWxAG
lPnBlAdywDb5IpdknO1/Li0/Lptkt84I9/b8+HswKpTPLR/8Nu1LDmLVnn2/FN3Z
vQ3hmGcE+gm+nZNu+XRwbJKyJek/1Ww0HqZdRMX15A0++tWCbd9okVU0U30qeqvh
7rPdUga4QeIQi8vzgLEcN+Pj/PcZsQAIfYHAw1WpxqFPYfobhA831Rzn/P+Zke/T
NF9y109envBnfYIg7aNu6QrLXtFXpIG6an4e4Or4oglCOWaLc3fv7Lyb47Yh9kXP
Xcgko1zgTl8jPnxB/yNDMbpKG5XmIDAVDwES2kXepbVmYWImUbMfkdOfF0v+DsWG
vY+qh12vmXpa9EQW1kCgEWU38zlYDldu5VyRPo8okXros4ruasWtC28KYDinUVMr
KhGhHnQzODMLQzqHHW7ZvAbPdxRkpz8r3QvythDsA+2EytoBcTn/ksh9jDsZ7GhT
h2PqghhH7P2zi6jkzcSiz1S3rNiZOSZXvk/CSfrlRrr4hRSZE020qscPFWlkYK9F
+zA7XECpTSmy0kEUYY1qhfwPk2zE+3RN2W1gi7QSQRaQsa3EmoMGDecLXbXwIwWx
746gHFylcdmtbJgw9y5/JOUrTfFYDGDrUj+hBplZRp7fe8HV9OYWUq7ZB7/MOUaa
MmJVEbiYfTeNw2cH7yRnTd7UtHxX3oMFyAwRikX+8eNXkhJhx73k41thb25+ScFl
bA9pj5ryjDetbp2tMRsy3NkjK6RRLwqdohXwJj3ywtQYfymdgKTkVFd+NgQab4yi
h9xepX7dNK4x3GQT4qaQ6zQZwaCdQFnOAsXDkG+n+QFsyhviA0IcvtbutBg6O+7n
6a5UzvCAwMGiBW/XCjyruvT5Y3woQv3Jpwr/NqDzYXzaY9SRxi1HfNgDGzuNMmRu
ThRm9tdPI1SRgoavRF1p+ZaPrK6ECkB+MSH2/OCmmwVcIIQhjupWTcG9ejfKk4rK
TnjlVhG3+QO3Q6/CRYdoGOSEN+tiZf3a24Ek67SiPgMLsrVPe5E/ugq5aMnUDn5m
Lc09Ur2y4rfum9wMTyvgDV+/YemwdLccHrL1DkQWTnw7SXD3nLSDPoN9gTIldbzz
Lk+R25JL/4/5c2xVi5/JIySbVziM+Y8elhPIo/fQZjFAzRq4o7SOUl9gbREIkYkO
qDCeRCwQlR01EfCoUp9Y21yt5mlQ6HbfrYZ+3fhOhNHHnTvV3zRExw88f2udFDXT
uts0/Fxy/vOWGUSD04STDzdot14rv7ohhpU1DDPswHEdXcSma+/Rtf0EXqUmU5+d
M4+Z+WFs9xrgxdsN6tTO+vA8MEOeZjOObu5RAkrZfJjjVG2h7uHW+k1nK8WoudGw
PICsZksp5NQfecK4YZuDfczmaa995MJoN3Os23JBwFb6nL05Fk9/I4ZRr8Zp/ciS
uN1G7l+4heK55LnOcVzUIyn19zo1RyshIpZHm+xmbGOQE6X5iivabIhzadVAhTEU
C2GMClFxvC3Jv4zccDM8w4/4lvmNkKchfQhv+XCaT95A6bi+cDjn/jszTaBtbNz+
KCoBOfoXG70v/u1FcqWvNq/NtGnCdiD/09Mx4P6kKAhG0esPIdJ/EmnrNydHClzw
BDdCqShzTjC7RXNvj+RDQ91CxNjBefOQNL2j+a66MB5V0t3HEhKQY2kmeuPu9A81
8mhhBPSRmZqBEjcpRylm13qAdOOC07wWWtc9do4YRLb9Lop41PJfvqxDtjrlPJJT
JvylDkwZ3AMpGKT+UDaJftgWkpkL8WUwX4/5DOplzcq6dQTf2uMInVYP5MT3NSr6
ilQuzvNmLkUdUQdejN1P/Ha4YDwJLorS0N5VdxdS8cv/40eJ2YdHR8LvImJ0gfnH
YtJcLGQjE+JL+FTfHBzeaSEUcqQlBt/d3Oqr4l+9WVxeIMXwZTFcyKLcARXWmxIH
iMZ3/3AhRfleBRDxiOPKENDs5HV/FimadC8ePue8anqgS7/SJ1FqjpfGqj57NGNU
6XHZ7cM1JX4qixu4Rtz6qoImN7gN+t2qCBEzYQPRgGBzBByK+345LKGad0mHAHH/
YAfd1WxdtzApseUAERmKPexc5ajF7qIr0aDCLyrI49lE5U/UGOXm9xy+CrkoctHW
USJWRdg/d7iqbHdxPz5jJO5cShb7Ytr5HAt3SGYcbkDhlTHH0bfIpkhj35+NVJsC
37hZ58HqL7oiMKHCuKQ6X+nKD/FT64zYE6X/z73TRh1A6YCWhTfNxbjnc7Iu3AUb
2rQN2UqUo0BXfZZRTjrqn2rCwCUSjEt5sxNslM2csNOPpBMkzcGrdCE3Anp+rjC7
Q+c3vCyJ5YMOFkYO0P5L5lQHGbypEbLybJ4etO/Ul6dJp2RcbM5UjV5L7vrhx2j+
j6S6Y/HxNNay/zmn5nHnd4eFqqjDRnnR+gbhBlDfpMWyHA/TpQPE3Ee0Fri9qY8d
7x+xxBT8s3SZ2hnVs4e8cqGeA/Nac1mzvZTTvrBZgfHkwwnqDxEKIOWJd7SpQ6lm
tUluETPEwno+6+nJrSUoeJs2otCij0f69NyYrpV+Iizqc6PJWdKzNe+2Hs9JOfCc
UnQC1MWKfiF4Suw7WdmYiQ1JX8ajJ0CKKmWb5p08ZyuoAd2yqOJwCj0iTVLebVtU
31iOZfV9t/iWo0r2LGFSsG8taYM3lPuibAKPP5Xldv+1wmWqQ2QodNFD6yx8qYIY
ICRpiKGx/GCJWAR9QanwRh08wbJ5NVUUoue4brlyTbGcIykqdmBAEteQsipxstcl
0AYSNaGGuPPk6H8aGA77HwCfdIHZ28SOtLNJP27RbpIgBZBIs23F+OePw6cyBMEk
HNXpJBuNT7w4Q+xcnndTNbzYmmCLN0sWpqt2vpkBxOR8oyjQeijFs02/TnVLHkhZ
jupmLio1QzYW91bifVw9j282Zjxn2frr4wpe4aAB+KwOhhYNDszRN/TCEBkn2b88
P7aBh5WfN8JSi5VwOn96XzObZ1HgvxKdmx/kBEqWr1b4XxoFBno81vpBI5AVxCLH
1XrCY7tJnl2v0vGGmLDZWceXJboWz0yOTP1jk2iNWtxA1OPqJJf2OKskHb2SG7YV
Tbv3CbR5+g5M2VMldanNU36u/YDDwcC4QAVnVptKOIeSSUZvF6q9k2ashVleF5gv
ylppE9xyMPYYcVSywod0rdgCmbLth1yLDHueQCnWVJpt4Q9HeDRGUKON5YSntTK7
bE1K5uWpwkoYYVi2ce6i805LiTtSuzuKj7X/GPYV6QrPLWkYRqWJ6xtcMyeoLSDG
kWP/JO9I5s3weraCPpaeflwRoiwWa0VS8kVRxVwZ5XaOKahBFaE2MgpiUcfwJdVm
LYXIo2VJ5h7bn9LB+VywygDA5VWss6yRo7pprjJfpl7ZlFacxEHKLh15cCI2kSqn
wVvkoME0NLu+mzoHwOybMCgt13C1rPuzcgPiZA3zZzgxibL9vF0l8Nx2T/bi29Wb
7WOomGgXJo3Vf9c6jBhHa93/ovT4mZmH3L6QjRC/ZEDYEQ/XQUquoBygPxTNihgc
AmzUm2BUSDMB8y5mc1ZhEnMdf48dsKDN9l7sg+bh5qEePtL4Gclacxeoetzp4gQ6
nSRIgOd4gAangN1uiIvtw7xMDnJC0br+O9OfQ2fTvUgj0tFfIUJvquJaZpbM2RGq
8/hdrZtI07/DosTDkfAdiKdE0CdCb1ZJL96FuLhA0xhM2IgS34wwTRA/PbsnTfdr
cw7skQHFUPQf5S3OmN0/PQVUZTKfnYRVv2Dn7yD8G0eDpp20QBNyWi/lqtISed5Y
nYKR7b7TdSNFKZc6gVU6D/CIe5FEBHzLf+qZKB3YYZOYg+jbjzoA2KkAlKIs9se+
yYgIR8ITY6mik4ywvOCXqSiF25aj7FptqnXHOiZnO4v2xUHm+yWMqdiHOMkWcVS/
mtCFlfio2JhCyW5hJLl+6bhmRM/spn0G4rFWtsrzgQYFqszxubi1QNmo8epI4Gdt
5j3m89WriaF9reiUqempnzSk8nDifPimO2eRddrKYvJ/rfkc7QWVDptq8MPdrttB
Isrwq/ivZZgF6AlbZL62na45GH/PPF4zm1u1v88iPsZlFOvOww8OlMhTHpfSBIpy
AKWd1Fo9k13ivBnJZ73lZFft/gOomjTl3/EnPSbF38XeuuHUB2blv5NMqy5nmxPT
ZZYz0jDzlZud0yf2gzfJuZm/jS9X62Qe120S1sSI60DSkpi+ef4VC6n0NTc3t0xv
3Ho/9uDVtCK6QWygUhv4XhaU8cWh145FhXoEM9VwygrBNQIOmXPvB+11AI9GUGoE
BxW8oe9N8T76MFDais1Yk+OY1PNkj6kigo7nhwXfFllYGQgxvS/peDyOdOzt77nm
yFxdLcjL1LZ0/+TrMWuKqFH1OoLCKJleFExp9+UCC5dSHkGiVAjA5vnduJilWxR0
KFCZUS7T+OVRFsSZD5GEeBzx8gibtatjr7tZWY2nb2FlstoTk8ZnEHzntibO2fZd
X1E875uCJxX7N8JOg5shdBda/1wPOZFUbyNZ9/b5rZpCdt+OHOeyad/nPlvFQrDt
YmM0E83cZH8F8BuIv2DFhA9NdnPMioyq5Q/vdSPODS7GguedC8Pzham+do032h/u
Tq43/zwA0XH2aJ09AOoB/xZoOVNBeCQA91f/SzA+o0BaHn3+xB/qJZw3yz7YwNki
Bz4DwOBaAIconlDPGqksUr9KZgLmnt906MSF2PrbpI9/efmfIcKuHwWeKidhl4tK
uvrXOmARivIPOmuksVpjc80FqHuu81JDtDyQp3lR9/21nPwQuo5bJqeFQv6UCjPJ
8vaj6o16x29hqSglq1S40urTsNHQXNAmI+gPb28xQRiF+W5/Ny5JnldwotHzk8pN
RXj91gjSVhhXaj2GVlkXFEvZDBBeGzS/WPGkuRJ3YsGBUvEPNFI6DAm8+60C033P
C1XBNMUlgkYjcNy6FSQ3eb2xlBKDhloJvnmb7jTYrR4c3kRqAIo/Hj15Bq0tAabr
ddmfLM7kma1L6kxQQKnwae+vfvIcBRDLQCO04R5V4yUciHorj+kYYQrsTW/vSc6k
dNcOV4YpUgrI2zF3vk94MXBC9bc/rqwON6J8KTkEB5Fq80E6u1W0mfJbO9JIEpAl
HLhc+Qd1fMUxl6wl7HqfBzzgznSLNy/gTfIncw6+gjyAcfL6FpPJTSEoeXCJvpgZ
00Owsz8y2C6RsLopBFmekuY15PVRZgsW8IbJB/Ol4duDrl5N0Kv9aS5DxaUCLJnQ
g0nhLZqjkWsTh/BM0WRi3yqlpuR9IfMypjIc5Qogb3WbEsJU5mBOUBllQ9kbO8ka
6FAaGwD0ZNTssdamtAJWb4BxFJa9D9mUHL2xrnVhDw2poDGaxvPSTf2HIlQhLPpd
3+rp2pupWPpvMvKC4nMOtop3KDAoBOk3wmTHIR1bujCEHXcWdDoljwSWeiDIlExM
f8nK1yZbIeOxkCP8jAjcQkfqoNxWX1Z6eGXM16ZzEucpZ7CSNXzLEjLkfYQr+HlJ
w9kSaSvmU3Cr4FNBs53yoimpL1X3BoxOadOZIXkayB6rhKreJM2K1PM1oLDU94px
pz6r4JAApl6YA9NWXvyWJ9ZD0e1yTEDa8nqhFsgRtk4qrDeOQLuoRFilEDcnZyS3
mKOqZCSmqosFxf65zuG8aOXYaH/uGn7V7hYy3TKQvz5aeVQQ8v6Or4/6xd5Ji0g4
xj8EGmUMOa9z2vbEHxMOMjYo7JA05nqidik8NGMmU38Mnl3e6Q64WrDPHwTRjZHM
rNuAfI7VXAGqFqJhBYrQuQ6BBcScvuRYSZUHOC6gOwXdx4D3+iFTBp0D5zv7myDn
FNTdWZoUWR76vkq6k1frwQgMnNaZAo4zYqWGMGzYtRxYsSkpNV7bb7+OzV696n+V
uqpQTZ0JmU6z/2BvZn5V1o9TRlUqwVpbZ7vdDCusB/Lr8cHP2/BcTtUIb2bgHs9V
6muumzxntPuGq/LYN0VNOosX5afUT8xPe/gP6Kgr24XRYnO0/2gcZJdJHumhK2cz
61S07YuAYoiDyICZp0LHdg7438D1HueDCGtmT6Xuh6Tv760ttjnnjWpm6SiwgpJJ
CBsFsmp+splpnhoPAlt1dZbJK+Oqs6JAyI/Fq63TmD9KZt75ZsxYuovdlgmY2ZT3
QmZfDeyEFF2jYFhPrFeLGhl0cvOtssdw0q8AMo81DQbOf83D48MqvRWzHtHGH9td
rELJJXyUl1VF/W5uRUgaZQZO+SzsBcApyNUc0eyhrDhBTnVnSlGByjMgfA1+Knti
jMJ4Txeq9N4kDwiibfVgfCziAWkLAlEHLqrUxZzqWAZJfOg3akKeluo1fCVKR+LJ
Z2SWhAqZol7iG11/RQhtu1nWIXF6R++faSVBR8H8WXml5PLLnrhjHgUHxgLxoE70
z++9Nt1V/yC9mE138CRCLM7ygYmoV4VYbMdFN7ZwjXvA+Ylxaob49cvXfA3rrUhz
CVpmB2mw3Lb8fIg7IpX7TpwU6RZY2TwKESpRGPT847rw0iVTrI5vJHAa5oEMVpjx
/OPWGJnGySqiIwtERpB/PBpWw3CgniFTDsM3V5xRN/W65N2i6Z7VyNtYv9S9nIZl
R4NPECgha5F7t0GFEs5Gco/P5cGG+ZstWzOyilbiK0F9BCiWkqGMxXiwwFNd9VLL
vb+mfRPb3Wo4UAkdrjibPiO67SCwf/q0XRgTVITCYhRp9Hr0LYjs11aitpCOBuTj
7lQt9QnN7jiT8fq2eTQNJiAGn1aozA1V8iJHye0Sz1D2hPI464ZtTMK20Nu6RO+j
aIjbG9QAuNXg5PO+JtmfBAMPVaH9MaziK+Ooz5LwTndATxs1EFgSxQQ639o5rLfY
d/Q2I4gMQpyz7feL8OFhYwODyaD03pl6THZvUccWGuoIPypR67qZg1ndQo+GPECP
HGUSd9PblUn1wOLAXQDgSINbt8OapuQVCFYPIZ71dHG0evIcohIzAMoZHnf2Hvbu
Cs5/skgZ/m35JpjVw0GUhMVd7b9flQ658i3XPc4OMpuC35ldkjidRXNJ8jGEQzKt
k/hHIk9o3cKUC9l9T32EZbSJDplGBruj0RtoxqTd9koFpDht4p7d9GREdtc4cheh
ZAQzRJ0XsYkxxhSLhbYXVtnBlkJJrTjj8HgbmJN7pC2YZraPzbFKtM8T0gI7vwGQ
Lr7h/fbK/+vhIpVsS2PHv/Z0ADdmsW88BGhXtSx9VO3+qUC2+ab/ab7ymTUemGR1
5V6AigCpEryt8fMT4ZmHx3W2ozZS6yhrfTPOJi760AMiZSdCXThSQBj2rgsSJLq6
eBnxlOjDYNf9lmNWfENryuaXHsQ+RK7MT0UKUMp1MPD4cJIm89IQPvLOEUA6BzeI
F7mP3nRN9mGDkqXTuu6UdWvi7MwxxjFT7mIPZMpMfHFkljnAPtNyKIwDEC0lpxtw
PPeAxNyUuWvoQs+HnkBEjI4jXOMVNbkIL5aInk9oL2/olbvRrimZ1HdAm9ynQk5b
VMzbOgU7Sdqk3UPaccMt10DRl5f4/cnRdj4Sf6L5HrMlhkLgg4RXwASDkL0J6GLM
5JwyluF8VOMome2uRrVXc4h/4Oei3bl/XczqKrMCI/QLdFkANGE/Ls+npL6mkZyg
s51AJVpILukRZE1KZ5Fj9eHKbN/Aw7T+NUtu3JESbK2zuhzR5lB0QEqHHdg4opfl
fRxPqOwu1YuFEF7H8XeuhTnglfzIdlIFLs9jZ4F9ivRgJiGDkGYgDaERgJXo4tIb
4EgXTWHqk/EY6WQT+gOy4lMAA0hpiEriIgZ2FntGJCtcbCiIpuZAWfokggM6hItm
FRfEEuiNhJXpHAx5TBXm/8A9CbyVWBDNMs/BndWTd3p1lTqYyIEaRi2Lvr1USUsz
n83+dYe3+2JT3/RFbpgeX8ZHdv/6rZiWyi4j/NbVCn19bszN0Lo3TBO4Q9qDVvgo
DwPNwo9xJSdCzVOjCm7Y1fvJlZI9oXEh5uwUsBPi9eLgVRUlEjoILyTEEZGaH/R5
MJn3BPBSvtUY5fzveTOa/cJ7cY9PTU8jlwhkQPO8SNgwTwCaL5pgqjfUFQ8J1MyE
+sD+esRxXR4/bPSxDbsV/MVT2yBSwA8hzTMCHhPi5sYW4nU4fJjMNyRV3ggREOsk
/TvAqH66PQlb76CIORwn3nBxJ3a6ZfOE22Bo4jqmCYIL7XRYgXDMEnsuG5Kh2ZjF
7mZ1+7NIUuoassIbXs15Yx1Q1q0PsbH3zFgpH/64crtwGagI2cR5uN3W4e0BqZQC
gPNiBP4ZcXMvUS9CnPIbE3UBr3RzLc68uSb0XUI4rgJ9TzelAfSi1ITn6VhXkbU5
vurap06kDEm6w1R5SgGt8if8eapimapxzsIhnrVEekxyFmPjdD6kW52nWPMKTt0R
igSuTweowgJXDR7+gHWtHPkXpRdDfyxdzfHN799HSAwfGGjiijQM599b0atXKEjf
OJt3MfS3mqsznL2Kr9EblVqzo0gzObHNR9O5apkwu+wdlYc8Emw0A5H4SzY5e5pP
gNG2yicPE2udUAwI6dEYqAi+4uodLtAGl86B2k6rmhFCn7KoILRvmsp03yWdwow6
kF1/uq76LjlGVkxtCoxxPbLxyt55jIClGiQy3YstXYiG9kjnEGR3G+DL/2bRthyu
utqJ6ovFWFtFYJ6UjXBMhxAmJeuPYoU4eANH3igHrLVmhiu7HdHE+AE8gvYPcdwm
exitld+LHkczcRbrXz3YxEEVOE/heHyp9Fpaw2yiWsHnsP0W55nY6crjD7ZsQicV
PXxyAyXKT3l1hDws9T4uk15SwsEd2P+f+pfJ1W3teOgdAeY9Y2qpTu4rrIOr//y/
Vzkfei2bXNskRU350I4Vi7Hu/FEcMGJWIEReMBcfho8ids0E+V8CThijF1AO4pg5
ukIo5aY6wwihO87718WRmViO/6mpJq2s2E7n6UvP+4b6297DUMPwNLBS8Uwl3HhO
z4EIeqjEw5qsAS3KTd6LXWCg9fJNB4v/MxFqcjoXh2xTdG4T3BqGGafudED0x570
9jPeVv8y3jSInDev0h10EVMBpzuec0u2DWMmJSixW8f2xvWmfIu+t2ghXoh4d1pG
QtDKl1ROPoQN+RrhQA3iQfggrx+LuZfUD3lydD1eZxOjOpMA7F8thTP0y7ZDm+8L
nzlPrd5UaC+tSblbvNIvAKuQTn1JRCZlRqRURhjPz1faYlCAuXcw9HCknc8PNu9K
iO9hHdyv+H55+d66E5uHsun7M+V9BXvnkmWhwecDiZqtdXlWyRz6Lm708p88xgt+
ZE74067qPKhucVcdHetK+fW6TK3Lm2N08kgNOvd/2ZbJd1NGnjjFebAI+E+uwMgI
AilivrwlgfXbmW45dNXuBZEFlIyQ/9QXpkv5EkvGXg4BldvMWxo0cjsNn1eRcFMb
ekUFJlkmkpj/7sbKeVpWp9LXZDKTT/TRYrJ6K2CElDnoQX5cEzmC9jd7w4Sv+JfZ
QYzxna2f+FWcuT0vj0zaWGPycz8Uv6GCWB9kHP73/Tun8bIVW51zn0gZj8N0GvgJ
lTHhMRdMptpduZ3UXT1gCrXFHa4QYAf5mOioPs5yD6rOcnT0lCiaJrODmhgwqjMH
geSXeZKf+J3k+jM2vhboXElrcZFooVA5qi+zqaNN14owwJEiy75ZDhQaNU4c1xMl
HYw5AKA6IssDd43JMT/NPPj0w5tqrQZHPMvZYJs+oqnChdNfdjKadB5/GhNO+Qut
10+AXLFA01cM7AjZPIQoUAc1GItgrMQvSB8tRU9Rpk0V75lATtwIt+7bCcb0ib13
m8hWR2nDqnCkFKhyCCnRnQSSJ2vumKNqrtxYIkAAIgN9I/QGKC9gXPXYf0Py3Uu2
K55kmKC/d5jPrmp2cJXT3VVB9B/2A5ZLhw7Ke2bGcYicX9pTWtUWe25+FeZgmA/x
BB9aOzvdP2Z7beEOBSMSlayO1aLPzvliIjaQlRcd2pMT1mUlreT1jcenPOE5GlL+
A+7qYNUGuppJbvqyKoZHUss6ai56KsMaBKdKX4nD0C/vogHkRl9n7n9gmc0Fav+n
OXYuMQ+gxiYOxX9Dq38gcpHv6TU1ArDtVJIpidvQJgR/ppiJDINVYtApZuIyZf8w
2D0ifya5xldFjhCVNOgE0NORlryIT7PluXjlEwDF33EkZh9aRU4uI+xUTRu9kaWv
0j/nbBvlDhVXkvMQ1BAbazsKAEn/XO+asYpvS7swYE8dsnQK+nXjxa7KEBMY8eT2
SLqb+qj/48k1rsORRjboyVnlBGk+xprVtOklnLtX1bW7mvH24FjcynAaDt+8jP4V
DaoeGbzBsL7wUH3ciOrn7QL3CIjCNyhbPvcuFz1+b0xk1npnvm99kuVziRM1rBea
tUGy/Pe/uELgCr3DKMPdRuqyFIeQyCg71MnX00BPpw5nbVixdhnKnlI7IXXR6rWo
oEVjosjwVHxx8eO4qXpP+z2TJoGrx/ZJD8ktS3C/FRMTHaOwJ1xXn8T2ww+fdCZ+
NwROyLuV8czpDumuPG6PVBwI9o2jEyzLXwuZCc17uVaf+v7yDinlRX61VrGOaon0
MejTyHa1mr6ZlH67FHxyYojCedERhkQ/ZHY+lF1iBOK3dRDA3xCdjO3leZg3NgDi
LdD775bQssvn2Th0ZbjVg4eGf9cmO8d5mPp3xHBoKQUI7EOv5OyipaD/Rrx1u+sF
ym9xVBd5Xx4XI5pNdVCfA3SBInmzgu3v3GrxtexFsnv9YZmIqsyOkMG8/VF58Maf
1FXr/cX8Q3V0nQKDWePUf5YOY+O0y5oCFmXyWPWEEG6ouAjUZt4HoR8vAifJogsS
B4EIW5Ib2n+jT5qQBEe6CAwES7cUDbiznQqNaavf4bmQUan8boAQugnCNs9JEdnS
YjQDyStpyMV1AcAR2ltKZr1d9ZgZziif7pAdjGo8KxEFtdwLx2WlgiY/IMMu2YcN
yMxHA0mH/FGboNCMnl4LjoYa8LQjnbNy9b43eKXxKCwmpizsiIj3vi9JYeJrb4Pi
krr3eWabxZmAzmht14BkIYz1z6ZyLQjSwVntWEeUiTAzs5ZYGu0+C6q/A8JAhotN
To+WfwI3XtktaZZWv3FBIXtcE1SUX0/1loNYvFv+xzJzIUWoDGPVDW9rUfmhgORp
6ePk9lbdi8sI1Na2aZrlySTx94nfnqU+mRERxnB0+dGSVKZA+KU7ENFJ+uqBKEy1
Fq4081tlA0ZMDamdcDJ9F4eBAe+J1vAoAiuagn0UDM/8hYopGIj/u61n22kG9A34
C8zLdgva81OSkC11pwUMjK1x6tN4lpiAjMOmHoQx8A4sxy8d0FgwC0VVWbcTA3Cz
bhf7HJKANKarTW0dyMUHLCT5pr5ZHl9+G7hMGM3ftXnkxdXR+veq+k3n+QsGGV2K
Zh+0y49Ztote0Cp+bEJZyl6OkftY17aRmrmSVJhDmpSuDCSeitn03m52FOT7FEaF
IZh7r1jaiW77zyJiDN7smPiKW9N1DMLDaX0/w70VEnxuBEJW9biBVUmAwwZ4mvLJ
PhLpwRnVcl+BNu5e5ntcwM89iUpNFbX2TzLUA3H101JQ8kkWdpV8NwMH1vGtLcft
R+7lWy4nUMMrWT/lY2PmInWqeddYaqYEVEcJww+dfWdAT3PlJ3DFjBXnJ8PzB2aE
haScoj8KzN8foQVew4fVL78no+f4PI0BRnNkS7YOC3VZ/9PfM6ZH3zHcb5zg6szp
qWdPqTx3PCREruzuGQ1B9wg1oa06IBMia0XrWiZdYsIsnecuZVTeNElVpb1NrjZN
+gMLLjIdM6Q02KpfIHFBwrmxu1/hhC3PiXXpK7a3HSPJ5OJB49J33QVwQ8o1rThI
MaWJZZ9dCrU+8R4sm4kxkMrpunxLiGjY8pUvJGTVv+bPBScdKFIg2ZGjTTn4lJMg
iwQUHuPhz3cfFMEarSA4nFXuVLrefdaoz1Oh/rhv3Tv7RfxFOYglq0eGwUZ8yPi5
paa25VG4+fQieuefRJUpK/ApGsHHjoQUnxKC9O+trkpEp29xGXfpnMK5JZimeP/w
x/c/HRzt2B7W0U4r6zYDGgJz9Hsy0EJq+YmfOB2FGObFP05ovTWB2L3DdT5OdsUU
SgL/nwcSG9hZp9n6yC1Tnv1slbmgRCUuoCbeYcE5QaegQ5ZILHW7LboN62r+rvwK
UmgI56iax9NhEdMBqOu6yrsSLkQjuar1mK09o4wbh+YFrLEFAKu1GsYmI4xCMDmJ
OHDvDg3IDGGlV/u2SrSmsWNNAJ1qh2q2ElDaTtsQOkc6jQFpScl5ChOLC3XuaxOW
Q29w/mHll3KST7fWaO37EfSBUW/yFgAupf3YHKohcvQC49DOTtJJDjQXHLoJTC6s
AN2rVQw8me9fZeJmrsBioGDIrQuFjsYnO9BP+DWMhwYX85BrbnkoUbDrNglvBe/A
OllMCY6FZRkwinKjB4W59X9z+MjVV8yPyJlHm3wxg0+wVQXb96bxsUzz1qDaU04D
1tMxPdc1vjZW70PXv3dKosLq9dc97DDao8tU5DzXFXo/tubmEy5EDlgiW8ZD7Y0L
Ki/i5qGx/4uU4O2os68OSUo3NB90kRIINDhOJ8H6p1LTfwDzyTde6o0WBQnewIpW
LwPez+yydVzyEfLRFjihW/Px/YdXWWfjidkDqzm4027ymfM2xvTLiXQsMypkv8Qt
z01T+UKM79GwGAXaYnNXmGlLgrb0Jqh2dO6jnQpTFLUIvlpwF4AUCXSOXuunLjMd
THJiV3dp+tWCXVZiTVZmWHpI30DCQXwdT6ZsGvUT19KGLFAGUDAKZPFfrjn8pSRa
HiiZavDxdmraXKj/QtyinEgGIDMB76fxaakDpgnGKve+IU4x+fv/vFJHsXrj+MWQ
pAjDqN8woF48pZu+jm1HpvM2LDEMN0XYMRPdhE6ihUTnD4oaXTxrv2UvqA9vc6he
bltG1CmDpJuW6iHb8o+3K78AzeR3/uz9oGhxNj8eXwMb0nJQCgCF3VEDDjiLQRMi
VWqSN0UJZtoFpWrZcba8JPZYFyLkECJ8IFqQhauKTwPi++sArLDSiDQjB05sGHGS
I3CGYbj/SvwfQRj8b49tuQcfkMpyV3cIQwPGhn59Ps/lfiePvPlbW/rhYCnoMoaL
T56UuvOYb2/uCgz88om6pFzukOPUyJdyneZLiZnpk/qn6tE+rYzcIUUvFlimgjtC
FtPGkcHVw9+umkRTGSK2h/URvk7EdIwTU6m04SrBr2E66QnTl3W6aPD1Y2u76Sai
tcM+DZv19XuigfnVVrVgrWOX4QPr8/PFOiru6MdMdAtxmSTh2pjV/i+2BYQSKZTn
C0GwIHPtMTWv89I2p5qr7hsedC7FidWd4Kfgl8atF6nJ+s0aGixt8sE1H4TuLUVF
HKrqUPqGyWxNKIagwiWDUFuqA+bivcAiPzRww0k7VQ0zRRVMvzo/LCxAyQDsE1xQ
LKl3v8K3XaZ67TQanZ03OPd48POfntvtEpUD+2zf9VcAyu11gUONrxZsxc3Je4jJ
Uf9ZnVbizvS6zDW/ESWZlJByn9/DBykjdqDnDQas7cplEa94C5yBmpUrLjFKWibz
1jmis3WDpvyawdEmDXATSD0qY8pzvK9m2cXoQX2kZSlxQ7FGcrI1QqP+Oum84Da5
XA9lnxQhD/Ca5o9o3yIXFgUYahpGE3QAdVWzPbCvLzDe/e5A146q37cVyLoOTB7r
9XdG/A3ojyteWbV+HS/bIk9iVoqckKvDViASE7+lPvSrsK5VRali0SHEzrQ3vaLV
304lkFVSyBQDw1a8JZByk9IVWPlQTS+7W2dcr393ONs0PGzk749kiwJjDiQUUMXr
+T4UP1fQoQ4xHlPac+Nn2hQRgudJW6XeQhO0tz2q8GMejBPOqghhUmJ1gdrTCtz1
UmsJenwuHe/Mb0drue++XYPFOfWX8GTc3fjz/ASSK6Hg3Ay5AQMNEBoJjtYhWmB+
MJeyYdrYagY7rFCGsTm2Uo0jolZzzvXWoFe5gXbUF88lHWPDquSzUdplpLPaX97s
ZBjcmHTLNWQssxJ0X4XRpke6botPyv3T35TJ6XkWfaAJnX71bVCRZ3/OJ0KH6qJa
fTegcjYM09MFJxsd4JTx4PwXBM+rmBhejx2K/LB71OxRZRX1jXsOjajUZoISdFIJ
nKHpZiumojCKa0soK+ykcMWYwg1G88fNuBA8vZNweQKdAl06YUYF4AVfflF36DAS
o2QTNVyCCT7s+KDjmoV/oJreMNLcXprWsag13U/Uue1NkfSHF/S3Ciz0SjNCuQrO
Tc3yEWIjsccRK+u/eRZmy63q2Cp2dqPCMeRqq9fzBdQUyRwy6NmlpUpxSvHcxW47
82OJ0EEPrdoQ1/36cJ/hD7iUmErMjpnI0QB3BI6Usk8n3AOdi2jjTjnO/ZQkNP/q
OSutX4bfEZ7kBgXkUNIxkckMWYHZEl3f4+ozgAaupOEsfLiFbDbzhjDGh9VEi7Zo
Eg2M9rn+zvNCs3AyBCyM87DkYlI6kuOczlq3O9lHPFs5NzqezmeG3/5kNOmgg2hN
2Km8SrUZgmbkPiPcHmLNRg6TeErolZAkIWvaNtKhlXjc9uz4/CGGtYUFCHRthMXp
jQTFCwdtv4bMy6NQeQoaFV7ud7cri9L/yTR8twNLATvdeCNU24vl8g/KfW+Le70+
cZH8LTiYbJ2bUW1GP66BQrnlKyO72k0hOTQV4pBiHQ3pBe/O7+x0csmunNz2zdn7
VUzGmB0WL1oUrw4aMbxdKgWTEKkrSDHl40XP4i2lCspOtbSDa2LomioXWCfoYIyM
lix22HSCkFAfT+6wiwDX9uqQ1ybizDU38KPmF9xFY4sJZNegWqU6O89gToSz66sw
rwu5rIK0gH1xazSJsdy/DhmAV9hW+2FinraNmYmhpipn+7OxhK/5HkxJc+Tbboak
WM8ppXHwjgmIl7x4x9rOJkLlBBzQ1IFpBLzjnmvxFMMUS2W2a95ZaAtTsmj0ULRq
hSP1M+ndPheAB6ombZptLjgEjK5IMF+9O4BYBpepspw2S1vN++wbtq4Q+1p+SxoI
ruMsaX8clY7oyJEX60B1xxDvymWWKl27ED/XK1jy6YPpXrqVMwLumqS4Z7Vtc4n4
U5Ec/lGuRMNfl1jviy2bwWDWPL+wPZNcnsxNhFf+Am2ckff23f4aj9ABsNexI7OI
2JRZ5Wskxf8ym7tI/kla2j+CNcZPiBJ+z4ZQqSVQXej8NRAxqNlAbO3quoRxrFHl
hZZZw+QvC3qofWfUhJjQxUX/8ZZj6nqL+45bjgfxwUiSHE+DwVzlCPLObzND14l7
IiLEIVXNQ8L2eafBMcJC9/xVqnPKjBfCuqTukZ84Rp/os1rwznlM6jb3kCAZSn0u
/rxHg/3bMJSkqJFMU+KQk8kUaGSoqLEOr/+w6qbnsjlOCP3+Dzm+6Av3XU2fPotd
OPmkraPpa62wzIggDf+bYPVvYi8vhcRqkIM4SQCKPf+2Kdm7dfqRbXhaN50Cuzae
fUYIZf0vMqXOxJsNgdjWvCIvrr8gHPrPEoSGEo/7IJ/jieHjUenN6JsG48G48T54
eFvi5Jo9ImHnUBMm/dC56W/e2cwM1xqOvJUbPrlFxpAnz3LhEO9ADp7AFJ4eL/Gz
q0PkZg5NFsdXuBTHbvUhs6UuwbGdU3ErLU8HvXliqwEXR6KEdeqN8p9jkOhPe+8S
djMRMfnoORDO4j+3PkRwvEt7Q9MNiXrj7RjTgmG3TT2rzvNWY0r2co/XOznt2795
s2SIRC7Hl1Nb26ZkPpjks9BtveovLTmQ2r8YmAkFWSDr5+Dq2P405TWrrZPq+aW/
Iv6dqmRDhPNvOe/vXSDO4zcAy5MZ5u+bBCO1KhBxfjPexeemjlp0GTVRQQCoSqJZ
nlEnRYpA4MCXMoU4Wjxo5r3LLadxkLNxAF/6RuSfyDENHWUQmZG9HbrY6tCQ96mG
BnJiVQGrOj8ce8xUmI8a0vG26Nrx7wSex0NpvHMHYPtix3YawY6CWaghvSZdLMPZ
sffm6xHAyuhfZDpQPwoeIZghOxGXE1xFCV/l6CGc99EgIpiVkpXwOvKcppIxyJoh
HUkex5ZCuYzjicKCCrithKm2YPLunIoZXI3lSPH37v2EBoh2QD5QcYSAAJcuzn2a
l6kjy1fMdTnvjildeYZzna45TvnZ3217CKPLqiha2nAkgGubfImPbPv0UQnEDoaK
MOzNJzRUPsoE3RjpfInrJhflsE9ulDU2DW9F/JJI82huaTZaT6Bc4BKGpBvn1ZNw
gjfv73GN6BgleM3yFid02o1JESnlCy5ZfWm/aKML+GjOXOauo+AnRbYUlx6WH+wj
dEPHtHw7uYfPTchOCDwvsho8HPlWH2vjsQymO/XUbCgk1LWqulXceLezFPzBc1jt
HbALBbPc2aYvsEXT5T7kHCSArlf8RdQjwb3LBnhD/LDIvgLGvA7QaQ9VKQcr1iCB
tHyWkHT/UvkTf3E9kRbbg/0fNfzwGqBF+BXvFHceAtthBe345KTDcqCk1JdbDqv7
ScybHYeHl/Zl5k1fDLUqUsLlO66C+pEwySwZ9zbuiVlIs3p8Es8rV9ety1drYOiw
YESZ3kLFYvYP2Ry8+EtaRGqSdkvf7Cp2pwWWNUzMVpkTdHBAYsrpwYiBj+D6T+zX
FnRg1i5B7UCrEeP8fPyPa3cKQh8L8ksevr/Gno0UW5+yabU6qNpnwo6FE0e93J3k
r16R7saE4WwjXIpumj+uD09b6OCBs/PPQ0nFqsXglqFxsIkP1muQ4Ivph2E/w3dp
qH6rdBF8HYfioNU2rrlfbCjGKkJdfrcuDpXl20XZT5avgaileW8FOoKGCayF3y9s
V/7RJP6HygdfbBtuV7voGjnag6CFg9VJslFSoCGbOKY197RfdXtnXTA5diLjY1k9
nFehnN0kLGD8a6jMyL+moiXWGUay+/yLW4m5ze8zY3UCPJsH6utL/3wxy9fTaPV3
16n/nJ0ZC0zDxNL2H2JJ2iO0p/VsuPHtV0AU8V5iUmfM4ReY9bFQ42ESVVuxHdMW
DiXfgq8uHz8QAZoch0nLImx/t3FEA3pw/sn/Ufk913COl4OBK2QvlIEx3lJns/z0
mKCRW9NIbyDEd+IoOpoEahCxFNg6Eo1OikKV9v5Y5WTmNvyWcQZtQISKgfKXna9/
la2WpM+zvg47RxMsbMeXAI2hFekHT8Mbjex+vRH97wg38suvu5JCm18ciSan7JVH
b8Mshkw6ZqkGRjHG0bA5sRUVC58U/IL/b2nLp5oruN//NBg9Sf3ogD5Z7IhI65G7
vgnpwN9xVBFPKaQPGPSoh7Ratftv4CkrPJZBX8dmk1GDLSt92rVMYzpEXHQi2Yk3
dKRew9Z3JozJEFrIstCoJc6W6vR+Mhe9nBx7khXGRpQEO01+hL50XHCZGDPsC4gd
C0ZRsv2KR1nMcUJH/dcMBUsx3OQd0EGnhjc6KaSvWvJCaU6IqlqGU/BhNHvAOAxz
R3tDHb4tDuno/jDnNtGyGS5Eh9revbPbTgrcOHE2sDDwq64O+Km2JxGgYiChsZzK
9PFUkjg+uehOwEzXcCB1fR4mlxIo5LmqTCu64hZPliobJoa6O21DvDqeqEEp3OHy
45tnkNfSOMbaKym1WSPA2Bch7aKVwNaYx1Te4XpMZ/OinaxtKHFRUJrLAXUvTrGx
4tTGsJY9QrXolikTebInzpdEH9XjXaB7Zp7KZ25NgZolTs8cgZIcybeIhxvLA5bj
emutOcyeMl26O6mjx/l3qEUWUnDTPhqueVkCYLJk5uE5ZAd4OA8M6V6XZ/JXSLUY
jFDq5Qh5G8IENsSVf0Xkbcoag9FU5Ii455gLbvummqxY/Ui4Sa2JtRQ2Otqikl2f
QXYzpQPRDRAvyme0/ELmF1cGekVd8jscVrgqsDcNjGE3qqW5E7e5+MUbkfRsLylN
5g5oole9CxsfIM4GKF/+lR+8gMrh37HddLjoa6ekfXv7Chk9A/hMLUmaPza8m98r
pGvykn71dI1TXmURrWLUI/xDDtlWwvRQMdhywwYIoxUyPDe8U1pJY+rwl28cBuJP
FlZedqpXj5c3zxecA3AVeQ6RmeB0xBs7W0NMFmeNwFM7QbnictbMUDuhU9DxDzOg
qvOsuUPBgh7jwj1aqeU1udG1zirfk/HwbsNaVhyEJC5QEOY7SGRt3v9o1c2AHon9
JrNW1z+T6bKqUDQZ0rtIOOlF9tcv95S+S867Pn++el5yUvwIgOe+5pGZC9D3OAjK
C9ooTJgOcldshTmfxP4af19f6nKm3YS5YWsYCZCcZIfQ56bkU6VrnDPekBnnvzjC
9bOVu45fZM4tNFp7IM8nCRgkmM9FhSpvX8fVm8R7AtUi4r8DNI32bJGPQI4YG7Dz
mriq2rTVLLvOyyiSb7WaL6aDWPkas1V08Dit3GepdkEOG1iFK09b1aOIgDaHHj85
dGys091U0cE5NKBH0u0fpFiaQBhYwjojiLmad8kY7+gTZNXhuHDffoc8HCIksQGR
I3LZHyiC8K1rx/yWw9dBNvApQ3MTpbu8eNpIFj9HWK/TIrzeHvRwfQ1HwwDnJiuB
3sh5jPefjgMZGfXr+GU4EyKZiCfR88cJubSVbc4cPYCldvg0mVUPk8X4pQspUsV0
GL+2HPPmfsGsv5OxPQlFCWGoh+XOKFEFLiBNZmQk6Y/VW4GeS1cnqjIio0ryBgA9
WgtkgczwVdAtcDWhyFpixI/cQwDzbnoGo68ixpBPd9laVaB3WI38lDBSLjDCkOSA
d1yts3e3dNBL4lCJTXtVmYtyFpU7zGmB1egHYHn3xoFqZ0mlc0FArtvSyGOzg6BO
o28QV3JnGW9D6bG42M/RDRag7TKu9MLLKZ1v1iEp6fEXE5c8nu8mqGVRu7bEtJ7Y
mP9pHaGSRG/wTmQOy5q/dW9j4On4rv2HSxi879ZucZSktMF+iGBLb5ZNtP6qvbIn
BzvBOF94UOcDW2fqvgUbCIeLbNPT9AOPZnYykr8Ya9dqOT2oQOmumZguMkAL36NX
HfKM1ANs0gP9YsXd6od0vRUKxyzO+Z7iak576lo/vRq0u+Ti9bWeOscNNldlu0gL
yCHvw582YSBCF08rhxbc5KO90ki1nN8MCSXMPUl4x6e0SPfiV9IPTAFeWhIh5C1P
meABIbfSSSvxSWfmLg+qnaOAgQXqpncwXgPOI0fU4CzjItpmIdR4ceOWW7nC/gbk
G0B66tX/IMEZGS8ACUuB7ERZA2xTSOJYSVrVka+Ou5na7Ewy/b+nn7ZNw7PK9e3/
XZUbyd4/J4t9CAQCjuawniSSdcvvh7jG/LJVofjH4wWSgh5oYuFjbK/tPe8uSv0l
rNDTp+HCcqHMSQzFfEVwL/LmvARnHNa3a5obl+OD6Nlk4dtVZZ8QnIpML7CfxnE8
Y0sDJihOiXgX7NnkQF9LBqN0WFFYqk/INgnfuysfr3eqNAexdRlJgHQ8tJE7z0KS
B9jrhldDxJdmHHajJVftfJPYOBYpMrNueV0spg3+saq9fARiu61TCSCiOsENjvgb
BYXqnY7cHdzuKtMeByiHOOvwo8DhhF9kRct/XjakSziLOn8xC/jK2j4/Y6XkT8H3
1Ha3AqT2kUnB9gFnJmgdguECpCSE6q4pkZe86sC+imptXKhCMK34colZ0yClDh1O
otZ7/xZsosld7l0NNolC5dObBuEeEXc3BM/ISnzXuDYAb6J3xPdQUSojN+JTEolN
DFLre6fdbD5RfFJssiEX0acdseEtMaVkMqxEtmCqazfjADVAdfVgXDB81obQsrPe
Iqe1cWq/BNYTgVlgvyhBgp7Qe2ZhaxgdTYkDVjaEriNV0HjIQOmFj+Xt+NvAWFWC
dwAUwltdIkNOgtCsWeueJ14O7Ab3WBAfFV6aeUq95oNWWxan0CdkrpbyWkBtOUOr
XfEYLHa4Q7tpLCwurxURmrVJMZDpmG8Owkhzf12pufHG58AqXtGJo+Udgu7wyqds
MCB+vufZxxjIU5/FYIMJmgsOkPVbRrTkR9oFdJEtN7RUJhhYJyZPG7pGPRLkEPsC
iTj51qGBAy2AWqrU2059yoPQMqBszd1r8CcmhJdYp/8t12nJXuIshFPcAu6NhYin
DuhzOdRLeTa7j1Q7NDxygtxgpTsZ2vjw4wbL/LncC1eGT+VFYuR2zVM0siIZC9GE
xibK9r2DZpYKPhFV5Z7+FNZeNRqbIQkD7pPTrBWxwHmy73yN0IalkZM9HWhkH5rE
G9F+Pz+lnW8AUuz/N8PeWC8mFG/k9zmU9T/oeK4CNjSTdOHGgXaalaTkPuDXi38g
QcoXENNQoD03urNzuFqXXR5x3vk3wGj4a8hD6F1o9BoffMofuaWjSPXVyKq3OdXb
G1bpFh4TvmOO5ZfuxKGf/VAVX/bjj3Pk50JbzsecUZthhFBQ2x0ddFgQIwgXygry
8h3ISlISlychzq6wwnnyYzY9f+7fWZaYBPuFzVXdlYNgGDaPaqi7Qi6pFjtwqOGi
i1Ez5SWCTYSPel1vM4NgS1OgFzKOX0gY5uIE7/A6PxcXTThYIw/mS24OcgKtLE6E
T+rjq8hl49G1V7ktQb2Sqqp8eGGV4mD6cxjicGHaxNa0xmYrBiyQveQyWQhYk44o
mIXnqWMt+gyQOwjZqrk3J3xJumULXv3PtDpa8O28RCIxSJNmCNhkLbUDdUA97JhG
d/n/ceFd5UTKHQB1zJiAxo7XTlzPJs5mHrBQmrsHBw5tgFwTvTowP3POmRvewFAm
1JuXpaT8a6bIiwoCWnIZZJQBM7U8yoOYsZaI51+iao9FlKMcmYxLZUg/5rxqn3jY
/r4Me4drCHRD3I6heXiM43lqYilFZJQbOXDai8N0WaJFK5+j3IuhpxdkinU6xYyD
6tSH3EZBv/qYW0AHIQKi4EMXoxD0o1KyEevlNtxeNM+MIDwvNp1cXxl56mJUH6PJ
RTVaB8BQ7lCozQcKadLVxx6GLrXzI+S9+Ds0i7cc2zZ8aokSxO2xzvGnVUuLkzDZ
F6rfLBaZ6Nto8VbtZy6FHuD9C8mqak0IYkgpnHfaL/k1TnwgueTwJUurvzS4hVkW
cpgB3VmYGwobJFlay8xA43GDDgNIVt5vUDkL2kQALXzlxMm6qnq19VfpbwOB6gWs
CiwaYoHl9H5gjT1807dLx4i5Q9D7++K7sk6g1f5x0AIgT034th/ACFca005fpgnp
R6bf6/sHkKeP5grEuRKU1aOwcyfiamKsTG8nZGvcT7BQJLdNI1BU92iLVCrt3XT9
OZ9H+f9qd683t5aQcOtdK2eN3EneVQ1CuNk6E26idkBoUCVgdFv0i3e94baunMme
t2rhBh5TLUTk2C6Hce372JF2Hv+QhoIXqGs2Bq+Cjq8GslGkxEqXVLWq4VmfFw9K
R3l8VMcoNFcabDgxoEF/H6A68eR9rdA1zcW3Kz5BTQEbzx9Q6SMSYlOjdT2dnGV0
JCK00p9fFNmoWgfyCxV0dlXHEB7suRkTrhbBffKjotp1WsDIUQCA6MDnnrfWG07a
MRNpq0xoNKW9Dql4dI7hmqrEf5STiqPzKOhKyfUkrXt8Gzg8N0Y6CwayxZCWMwlb
toLuB35TcbwEqg3aQIuQ8V67SeWZvMSADs+gr8wnT5mXkWHfcyeSNgH/knsHLhYR
JmuYaO1aYBWbOvJQSxX1YAUL5Hmww5epU8iXxfbAigAWfFSC/5+Jy7FFoVaYBiiR
pfwrOGy77eVi6JE2cpowVIiL06rdQS5xWi1sTO9BAwn4dXr/GpwmcwaR3hCi94Hg
S8ijU9+SxYA91YOfVln2CcYtAXPwINIsmXyILnNeelzpQGZ7sq8Nut105ihNP3XS
m98IrRQD8dNo1FiJdvW8MWAVTxdrQ78VsxOan/7n5C7n7XRXtN6pQU858WQohE+p
jIefsOq+DgkjS5QOdkOKLehGazpBA3LxiyZolA9o1Rb80cfYgKg2zpXkqCgoKGx5
WBVOT1XJrrbGYMnOEetXBTZ0ExxQfmm32sEwd4wHPPSGIRaFW9aLqvQqHG7iOmoT
6E2b6bJyo/jRKphSoXmNTdqhqsuaAHvAOsblQUNQiEEbDzbm3VlCvBictvFHVIcu
scboAlUX73KEpzCltB+d94T5Owa1P69gtQDjnJbqzdf0svPTlmCezgOamPucnJfx
ANpO7/XDdcG4qXH+5xml7lTGuk0oLMZhAk/8BNmIbvSQCGn1/BEa6ENDlkgo3xdZ
CEi2ltSvRfdpQE9RFaUSqxLoKGwGPtFtQvg19CUC/bYGdXs56obQarIEn62RsT0i
ZYW6UhLrVDIavyrq3XrGIism4Suk8U+P3vPnZJzVfOtz/NTPkhJytqR+YmfK61c5
Nd28pAbOHZvQBkjFkiCG6H/FnkHW9ZMOLcecYd7CxAw8JlDEzdbmFkfJPElY4sVv
cMqGKp3QI+A7S3sgS9jq6GgbbeA+pyy3ATSEABqMwKaPLeyg45H8m/cxV5MZlUMG
8AtmMCxZoQC/kLW77yyWMRaCDZ57nryS8YzI2uFc26Uf7v30frpgaQQilxr/hwDo
QR4TV1LNqPZeMWUEupkdofYMCI9hCjJnnTyaZA5cSUlFifZU6tkt7mTM4Up0EBzo
jc2m+sW0W5aNzeIgHXgjsYSGev4oUebH+pzCe72MnORs+fuqLjAceJ8Y5OczcIJ0
jqkGPPQUIzSEB8dHkF7M5dKGhmDxUe65BO7YmQdIytASmXn5twC0JT4M7kczRIAi
V0IG9ZpIcgOSslKOonuXiGyYLFchULmwlGxrxYmHGZvOeu03C10vAh0yRK0yh1lV
fJKgbNxKat3sEECaZkR1LLo6av4APRiEJW9qoLpyudc+6hbrQSzb22a9rsRbUabZ
KXgyBnkoMnxtDO9F2jkUyXS6EBzmlE7fby+ynywoSaGl9oQoH8U0TDC/IgeFvyib
gzCW4WYG6DtpjGysrmw1h+Ng9furzDfm8WQKQxpTEvahLAqzOCpljiF26wFIkICN
rroCeBp/n5bqdhsubYP6QUqVaYRifUCKyqtKlRrHRbMvPtdAAjua824xSZwxYLSM
Qs3M+3iWKYp1U7BqzZGFdteodq6zB4V38t1ou0IQ6+JT1BpQk/vrTjsf0yzOp5N8
QxNb4e66wt98TlA7/K5E/MmSRniZe+hgDC+C4BTRdbgcC2fIraDyaEmRqnTc78E6
ynp5FPRAwpEU7MuEKeV18YU8OWYU0ZVDxjahv91flIMkbbfKQ35ScZaBXlbd0svT
gmFtUspaiM9QaCOEHbbzEzHIDoohUKvEw4Oth/5tDfs1R+4BeDCj2ntBTUkNdOVp
CS+1nph3dkhepi5GNw6CsZ+3skAx91M91ipA9xrGNOiA5H74BiXzcinbffY8SZG5
Lm+ZhouwGGZ4++/pK+7lqfRvXbDqhRUBz+Z5Wd/yklAT/t18gQh1bLHnYV5bvVcV
EeyZIjdiib54n7C0ShWgBZ+S3IeIouoGQUcW9AtY4Ecr7h/5iVAqD6G40isQ97Sa
HBS2sCzKl/QZkaLq1c4lS9ofhsskc3HxvPQCveDEU87HrZM9IJpd/THQeIymuQyh
5q6+ri5dnrqNGcBtjrnjnHdKve0DZUP5hNfGWRmRAv6MIqDe4UhAfASfNVF60frf
qlRQUrLaMCdeJ9OSNUyEnHHtvk5bs0PwrFeL2CAHTWy8+S849nMUwzfug6yh2mPT
VAUYLacbD3MOyVJ39RjQ+tLij3/Ec1jnKYdUGBBb3VvcLEdU6PXQ/4QWvk3EDqXJ
m7nLnzeMHZjqpz5QLCeefKQcX/pTWKrmHi0hU7gtuRUDjc/PY3K4SzBdF6k02tA5
n9RqFiSkvO4h9yTq/vFu+z3OHEp/x09DYM3pkb3Pb1ff8CDe9LDH9gN6z4wu7Ejm
TU9s5NeoeUf9GZ1kDGjU13/6m6vebEYx5d2xdoBGiIGQC8i5Euk76hza6kL3mttv
dhBGOukQVcjL8JR+YmlKKzW6JJPGBfMxiwrq5EspUKZmN4dLRLOjJ+dsOh/nNx1v
cuubd3akRbASqK2zSLTE7ALTDF2NzWw3LOYf5ByQo+kW5hzan9IuFid9aRRrKyQX
ZM9R/LA3lmvwIRNTHEg3jvrrm7sset3hXDa5NiXucxs68s3GTTeLv+lI6pBKyGBo
DHN1hsgK3+m/67up4gWijysluDakM1UNpRMWLXNmdoz70pVqzVgLrvpjhd5LKKoe
hM1tPg2XT61BL16rxvyPo/y3FCymcFdkSD8NXzTMRTdNRClhwb+8qhVvih22Cklf
O5VsmrPhgOGrK0bIpja3WYBIXfQNGpsbgBsIt4RlE4Wzpe9wIagEb4ZkIiPqbkUk
elT1E3wgURaeIKV+YB6lFanZEh39j19ljiMW93b4A/LqqqnWnVnNTJxl6ZEwfuF+
XFDi/LYY7J1/XLAE3XsoOYHxnO2jfk83zEu+dhZ93rv/MYzArTS8AK7DDodjsgZk
eUE3bWYHkcIXCXCNwf9N9QgTQrYDxmxK5qrtge0qfSWTsrh+D+MNgWSam8eDS1VA
VdOKXXz584mnl7Knm4QdgGbGMCqqAQmNSPgzhLIh7RZG7uuOrs0kFjMm5OwOmBuE
WXnqflA1Y683q2KcLRpL856l3iuy4FElOhtm/CzuKmS76do4EZODY+Y+PEl2XMTV
A6js2bq1zfYZw5YWxsGlVPhRyu5Zp0Iai5MnGkEfv+nyxxTXgLx8U5dC7uvTXMvn
zEP24c8jrZ3Nocg/CBLgZulEDuKYTO+xuwe+2Pvn8C+LI4e5hHrbzpc5mtxAS3Zs
P5mWDUDxt04o6GphNOmHoJdyJOJmioVU+FtMcRtSbw4slK56oSUqGGx3oxPJI/G5
MeGA2pkZBYqK1c21Lc9N3ED5v/XpQSmLl5UPJ9PXXMrpGqUZiLeQzyUTvCZGN9rb
11FVkooZIcfXilslo0o4SMCQWM5zuNRbmXEV2PZuh6V/f63R8+GgVmQMoyyhG8PU
GUDiZm+LqKP8kKD0z55sseb1LMD4QIO87ZyenCE+jZMS4FLzzCOx+LgK7TGAYY2b
qOITTdjpwu05Z+iYUced2+9uJP7ztNr+savYS4arTposMeGfUJPKsLDeNM8VHf7p
i6A+bIdFtVwJTeOyEhYUlsushaJQdSf+wX7oz2Usr6LM/3Sdi4wqR4fAaTx6V83N
x/thdaFEsFg5DRjvQrnYjSuo4MIZaYK9zoj+E3q0lPViio6ah6VPLQ1pUfwqWB7P
uJqUfcvQJ7AdhoPt7Fq/YF7ZS61aUu8oXZBV0C1U1682oEfwpdBXDyqzUcGGYYvG
db4AjiBXldeOHh6dcQfuXMF/LBhTi/XUNH316ucWCE6uuh8JCY9hkClWjU/pZr7M
s7GCvR9szIRzy4KFg1MIVAV7cvgWQ/62fo93VbCwPXVzuuN09k/AQUqByBXM/WM7
0N2pQDoZAqkmt36FXhD/lzLjeZWDHwxaDS+/ystAFi0TTlwbZJS0GDwXWgoqSLlq
9Eymchgi1y/mNg+/xzUiGcjn3mXxGHhnn34AbSNdc7rN410JK2HQaKNcOL9y/mtK
HFSaWP4h0wLyQ5bmHuoR2o4odmSQEMABySEX7j9lc3dpB1Ghf4UWhdBSoIXl9tuO
cJOJOvh8pXUz8BRerKXTYAprbjzUA8aqr3lmtaaFaPIGMb9FMnit6vol7n79N5J6
jtZKndI3+YU/mT+1h5WyUUOo50ynhe17O9VeEHqpo5lPEemLnqDVuCU/tUCrdf8C
0+uVU3Mf84UBn4oz6nIiZJag3IbiL5URoz1tBLnGOqjy2qOJCKZT0ZwikZ7x9A7v
Fcj+nGGfVfsECApWqJw97cHeMjdEUtlAAf1wU+mNnIwZD2F3T2gi94ygoyv7YfUk
UmGTBLNYNqTQKq7hryEmBjqMekvVJyVKblQ3ogbakE0NLviFkJmKk3Wom2OwQTSR
/mfmrGntErLJm/U+6Sg/kwN8BRb+oW9VPSnqrH7vM/j64fs7uXSS9zejMrUaDLWg
3lAo29N5Dk9VXbJoalpZNhr4QQ2GbHjbduUxR91RZLmth7+UIAUeH6PsQ94VEQZy
ZZOAY7NYGVD7ZLQCRZM/02q1m3p4lq5hsrZ3U3oM5hMasKEXVQ3JxiqN+fkXhBmH
/U9/oQe5zwBCMXmPm0vaJXmLluC0a2GWPDgC9vTfyoVkpi1jkWT4gHEV8SbKj+h+
FM7LHP5u3lsmy4BfDTown35kpzR0Jqt0L55UH8ZKoxJlc3rknaJp9aR6+EM9Rg5U
TunlfixHEWwfMKFGa46gTG/rYoce9jXiolWFk95h49H2fw9Ox+rm2Rm1j3rQPAFu
gTlHdB597YYoVBHjN3ciDrMJPNxVxWKHlcMNc/BleDZseQcFh8DthDMi1ZxgKVcV
bvB0zGrXdbvNbuKcIQCtL5/7V4eyNI6sKLInbb/0G+Hwh6dWJora/2eCY7XCj/rA
551vQDO2e7eJAYBEndVNhk0I2WEjU1zupeiqYcQG+Zkp+88dXhL0NLTw6Z8dpiS7
YJ++DrkrJ21Xa4RcB8FcTdxzQvFs21lYBWQ/trkeohJkLZoIGf9O8Iw/Lk97HUj7
6+1/5BRduaLVfIuBYJEJoiCy2jc29uQo1Df4+ovxqoa4C/jTbKoO8tiX1CTrZM6p
MJ2h1kRDJw5TEBjxpNBUdtsHTTlyUoP37RJJBuwl1EnlBeSQLFJapvYslBC2mf1I
PsLdhsukdbR34soNl7gEkGjXtk7STRXrcbGaym45xv7KLkrsBRumPd+W1fCX7VR5
4rCWcFonkHrHioQ/IclbDsLX1iwQB4sLDAKCnrbW8B5XcWjSyO9SbwCrxBTxRAsb
Yop0h3u6Vf+pZD3HSaVkRwimWGQJ3BNSzEOM9JAjNtCZv8RSTZXgzqkRz8hcsBy8
GGVCYH4YB0AWLjitsF4FJ0G6Z4ZLH+C2L0UYu2kwzhzBIJNkeWbLQAyJ1pQh0YIw
5ANREXuTeMOXmZOu6eIHWfi4cJwfmtfsFJ9jj69KyMx/NsLbizGJljixJCYuLA7v
U7pPWt0X5l/LELtC6sECeUtY1mQhdvzl10ZwdmlFq3B89V8vouAx4Q7/IUUF3gfq
iLJFuxVsdMKqo0/NwoUrF+MoHAvTVXc//obI4mgxOTyh6KnC4K8f8LYH4MULR+Ct
y2Bf+Aa69lEOCM8yT39lxo1lWSEPhV3h/R1YDgw116lucSZ2K4vd0MsxYRzl2tSR
SLfeRRA+HEaE59tw8irI331XT7jVqwUv+KjBR2u2L9uYovi7nstSxOXjsUVC1dPQ
sCIZxJd1Cw4wgLpVrYYC3sQbzIuEZnQJnkSawxS2UMbpqD2zWby1FEdCym0FPnq1
8ygpTEKFkALYat4ZGJgDyZfV75pxtvXYRZ+2pgfyqkC4T2ReduPObv0S7cfMd/my
Fwm/l8b6BHru7bmpJz99iZUQjbXw5DvFCdlv83sTssag6WFAeBQlc7IRqtX8VC0a
kSk8t+SxU3DefcS5vFD3dQcJRlapQClKb4a3bFDrMXxkkO1UrW9hDDu9WoSG+/vq
5msNIrj/vpWZLywiD3YnbehGXSUtgH7LX7fL5Gb+amimle+J/EL0d0vLuic26x2L
l8tzbMZ42DEkv2HjrR7JAoAjcp4xO5IVnM65X8jNwa5b88nCNdEAmIt03Mzr7fXC
EQsVQlvsBeTg04qIAFXQePpAUQsFgGvcd11MI/dBvnI78bl4nbfmCU80dtFbZRlO
TUhOpz6Te587w9brM3HVzandN7wpClwVA8ac17UyXJLf0Q4Xm2By3YxjsC+r7OFu
3helvGy/6mnZJ8cFCnbhaggPExnHr62G+I6XtCvgtnyChHSxfa3TjI/AHGKBsRMU
DHz+cGUqfV/eCJ9ai0VcMfaKin3ShqeHveTlrmFuGbaHP2GiyS30smIz5lQ86VSS
QptDXTAlg/eLfguwZ+E3eQ5CEvS8Zyv3VJEVtmsKkb6z9lXXOBTi7Jy3gFK4cPll
6MSY8tqptaBXNTSA5VRC8whXHjnHSNbKad7m909E2yzIP/zCUNtVkGcFQBlj4yvv
zCCDpCE7seY37M1JM2ZsU9iF8NHTjVEbZIR/nAomZVWT7xcDzvjEbi8ciHZafzHU
IK/6sZ5uA4Vsz0HWr9HMliDm5KuXNas8n550f9niTnd2/JJh2jWURxlSsOJmtr1v
NZXv59UcDn54nWUMjlkJWtaWIlLtGC8I9JG1n0NGxE2V+vVp1Qc6wPOKbQWHafLN
gdvDFv+xtWG4LROWEQuUuvN3WFaHTlBeSQCDdVTPdiG6HIkT8HhlCQ6cedWcibFn
G0tMAwCOtdW/ZkEXa+H3GioludsO4xsL1We2mDKMXqmRVG+OvUgX/Gwelh5IllYV
CAM4V29jVpnRBkvda5IaRnpFOOxNKt1UpvCqb4pN+QHPmkDF0NoOH2gaKsKy+86R
S+DoiGH/kyG2fFBb1eCfH1F8X0J/sXOn9/JAKcXApigedySTYcYk5KwlXoirwybl
V7Bgep64BNSaOMPCKzPSJCgmUvZJ1xiA/rxPQazJq+fif2CCULyWAw0u0pUK79vD
ULeAI+u7DRsZMEy859Z+zvwgH3X0lgW6IF8MNrgxGpfmmomAFpihvRtzK/KDSp98
viHBq7f5gGLNQofqofnsPnIuDzK4Ksx30YIvx+rFkUQUlxwcHM1aq5GuV/Mqx01X
76LGa6X/eEPC8L1xlMD/QcJSAxPK7/eEQwZlfwMrHMjBFry75B5uX9Wy7ZIhWz2b
Pa7m9iTgbAvniGiO+QXpt5/1MW0za8BA28ih4l2ZU3ME6jaMOH4p6MZE9Zm8xPU9
CGcMOKaOq1mg5mDlmVbzsKhVlJERnZx4Z2BWOcZQ5+SBZBvIxQwAk4hcauU3bMT9
1MM2vGwdueU5HzhEEN0xgEmIMp2bJRPgv1AF+JLxtAXO8HJ0gO+5R8mJeGBxctgV
D8/WXyFzaRsyDXd/GGC96oxYlh7DwPZIZBe2wlyPkmPUQv9FUM+MiQNI4KasKIjI
0nC3k44ixiFgzCwIdexOBnbW70ON2hu8P419OxnWUarM6kJOmLJxVgaNjooPdLgY
Kgs1r8CyJzNLDZMsyO0NecGQ+UGMxnNBaOpomv9mEqws6vIZ0vW6EAl1ZzNc47kg
MaILdLoSJWH3z9Mt8zJPCWnuT89li35tYX83Z132KDeCgS6AsSDzchNbS818kU2M
0p1EsuiunRkeL7fA5sz/cXfxYCX2W8hmQuobMifgSD9+5BNwkhZcyoe7sUod8IJC
52EDY0/rmz2hiEC00R3/bBZ0IEWz9kmYZZ3NdU5itfTR7vtGFYPzgvjEpb7jBvNK
rpAJtbEV0PCAZ+liWO2OxPFEltUtsvLcI0jTtWr4UvYgOvuRbjCLG1M/Yiymq7Qk
xPCjj5HQBFlRq8QeMmxtjcCo1DFqf4RAFTqf1yzMRLfSWb+/Vz/jt2jmevTSTc4d
zAVLP07x8JU3TSIL2rpHqbXtNJvYMkfFdAxs9ArNGxE2akVzCHTI1slKPvDFiktl
HwuzAW7gzYeoZnhBMtIPv2MIy7Ej4dFwxFGhhSHjWWI18eUkrafzd96zogBq+syq
KeuT68HlEk2LgGWscRFWeCgQIDf5qe6HFGSUdoMvAFuZ9qjIMRs0Ufm6+mQptqPs
qt6RFMzn+xmhBd8kmtm6ZhUKIkgVuJ1rXXrrd862ZKz+CaLq9fdlOnWVj+ghMlQ1
6x6d6xuhJDONRIBm5tsYfXYdbYVPDePKeEL5gqjWyCx4hbB2CrJoc599nFSczivL
plCLbC9arqvQa0XbVdo1wPfmUhn0BIz5HyIUQcHPb79J9Zf/De71Ee4Ihh7lU26W
6h3xirrrzD2F1sA/Hc8LAORa+6u1wXvHgTcmFoz2kuGFGlMdYaSyesfnY5FPesvl
Z358lKkueA482HOdveBYBPhcpQ+C083R35+CQVv4jv5lFzUFJq77feFdBy1VoqLE
7BoYv+wPw1AyFlLEERZeTrocd4u0LbzUgI0Kr4CkdXO9hlwWVSjFmaWvqV369LBC
oveNKZY9STOv4xNaO7BG65xOivrxWojRvrGHh8n3leyt/ARhLwGXlk9s+OEcz2h1
EV4Hub6OlBWHIcud0tgbu/FSTrxN8xmWpCeMm8V+JHIq7ACSwfbNGMnRdTl4+7do
A8nRcmiNrlTKLwWxY24WFA9kWtR2VrqLIQ5Tvs7hEfHbEQFzDZxf67JXErKFPlsk
/B2nqsTFGSpOZvj3ANfVteeym4LZ73dwuY3lzOGk5Jcg+NYiES7e/tp4PJwmtSf+
KaPR7XBRkOeAwBlp/JENdVXGZqcZEc88X8FzS1ZTeZYVDx1j/Bxdpl1wntMHmImN
UAais10cgfL/4D/fgekwDGVKWfa6CiAMz66dHu7SAq1gPGY5iSzf5CbrZdGXwW5i
fbnaBt2bQyjySqEc30w4HS39f6D+B/9/zYCMrh8NexIL3UG8LJK1qTiohe5jzxJe
qjR6+LTIShF/csXiMH1GSjzbuO8nbNxMZCy2wb8W5entSX8ryiVKFpFRcGoSbbR7
J6IzsMb/cNej9zjvKVnssE2y/a+A+mQitZPxZTKUVcXY2icXjnWawWvtV2Iip8LT
Jg69LlU6woecGAfbdRVxmAI8zWK8JTgmO7G8M9XRh/Uc52e6LExMnifFk4rCb6BT
xfItT2VQsRnDJs5s/737W0OTBIh1+p6xEK68pXghQvwmA9d8onLnTFyTNUeYp+RL
CQUYcrZ0gF7FC2KiC40qoPrfLqjxBwqpQjFhohbDUZOJ2FfqJx/wP9dv/ZS9RXM0
lhG6IopoFsf4bsPcatExd+ompVZd60sT6ljy2uzhWhIKnkR3Jl36So7LRrZjLO2U
Zvji1c35Sdgn75b5iuJy3OORlXs5i55hwc7/S304WHN9ptDWJ89BoYs2nRIlnPhm
ILC4qfz/Lx/oh0UxAhheOhTN5up1PfowwMoMw3oc56sh+2uLC8MFQrR7rar1GpSW
woA8LwMGZViqOgn4squvVjFARfZ7mhSClWzrY6fUnEwGb8wf161HTPuiIKnkdz5W
+U0Lm/09p/RvRnpMfGx9rHP+G2i9doHAC6OBouoxQi2sVZivv42SwPQ/4uop7617
8tr7OTnnjI0BReazYNt8yi9nYz0XQD3bZ2h3t0Uw/pnEuCmCbydgD9roASp9+pfa
N5M/qUJq+5RcynJo9hTkABeBUzjI1effAF1cUxGZjXnwhX1NbA63uU/QcN75MlbX
Je57aQFD3k6ZjQ9RqZv4JWczRWg4EmvRn/EalCp+93GWonNUOTfjJ2kKNhCdXzm9
ciF3gvDvcQ/7tA4Bs/4iZ65jjm0CiKXat+q7P6ENdC03NBLIvnZ8KhE24CBnLFzm
2uoLpWC0PyAzWPJbNntfdxushARBkHkD1iZ/6LE9Z953Boz33xEkb2tp0pulcsM4
B8aMDaoDR1N7kZ2RM6f+STqJsTiN3xpPJcN62OIvQEpoqXRUs23e9gRrOi7/BEdW
30DaBfDa/k8dwDw6Aw3IuNhWmkgQgzuoRmN2sR5hYY9FLjeda22pD4xDMNyGufAR
OnXyGq28UfuEUT+9MHNMLEDErrDe3/pAg104ojhyuc9U2Jn680l3dkyHxaIiQXfw
ZZnFdsRUJC0a5yerWOcNU1vl3x6xg+qeJrWW38XFDO1JRY5pg9HlyWQcJVS1L6D/
y7KKKh6K4xOgeKYN7o6KMpv08ntxkXflE514Qfw5B1cfHickDP9r7jcPWOYDNi1Y
2ujS9nKKz15ieNr6RyIcbZjxPH/fH2HS5KQJL0k3xabj2PAtjU8JypromDRY79/M
7FXkgx8voa8vPrq64YplCUA49fpuRE7X8y/KZxYFZn+fILVjfJB6l3sIMRRVaXUd
kkuXorEiYX2WZzUUmXJOsi5MCZtVYudqdu6d2+vBgVo0PusULNIid9S+MzWFMm2P
71lZyqgZv5cptwlhTqjG2mYm2PXctRb0RkhMa27opPXcpgQFe5xlH/7c6e2HVXmo
QztZq4R12PrnVBgZobLeAUEWSJD1kMooGH+4j5qvB9BEfg53fUu27+2L2gr7Svez
r+e62PzRrKuzumEk9C/Pd6V42KkfHzt0x64efqrYLGJgzot5BuZcEfLm9Ut7FAsn
6rfJy07KcoNtQkxWEdbxOLefqIHmVqDt3o5ekgCkyq+QGeqyz53MYiZpEivbvLcc
0xZq4alyXvwI7uby3jPujPHZ4bTPwhnvQD//Ku1WQzkZ/MRr8nA51NLcx8kfPWkC
Eq/r/8dCWERBtoekJKxSeoB/zVqOKs9J/RGej/OzTRGd//8CzQoAlRQ3BagZT/bu
YJ6IKpEc/hmm+Vr0LSPMs5AvQvJcYhYBSP8gMuOUSkyAM/4yY2FYzUHFFjWntwIq
EMdPNd7I7qyGFjSDKKYVhMgSrmwzcx8RX9gauy/WytHf8tvbGrDOusaXaGq/vSmA
G7z3t1foQZNXicuZDKM1KpW7exaOW1zxC1nAtXn0WCe80drki/mKA9w87MreMuyi
r9/89ZPUw/PUoo13DaHHQg/6fdjt0o7STZb9Kxi+2zLy3SONWeb4G1c5yVxK9Ktw
bRpm2UMzk5oobSHTuJEzCCgRkILghEIN9t5GWSfpdXu9ouSQqwBp/6nhhWAjZ+2B
2jGn8ywHpyzjhNdR0ITHp9G8Wx2ZvS+skBMT9x1XdYvNeuYJmZbevYy/3opYRFZe
3kWPEjsCL7CG9VOSTWLnn9MdKesnvUijRzjgpFMIz8BfACo28fSlHTbEL77aUuGX
DU7z05Sv4/K992HHNr4LhNY35x2Nlwq1hSZQW/eS6cZrni9fgkFk3PY62GzEUz8T
cN7GpqvaGWjXas+6WVwG3ceM6f8e6f1pXI2gZkFtNHp1trkGBtVexJH9WSONwrGj
qzi9Nbf910UZ/0aVlleyucoL7BlSLjVZG1mZdoJby63s2/axn/Uuf0Jdn6q5PiQY
aN7iEWJRBG2QiI0TLBeuoec2nrZCGXvOh9GtSTRvAogZzvPWT6UqMBp4LZy1jvVv
3ZRlYCJyu3zTcA8PjrO06lKBqEQWcoxxgAOzlW4egFupkk82qIJLFdIaglENVvgs
Ch6aOeCB9px48/FQKB6KGEyYj6NJu0J2kRXt9EUQWnpFLXaqfNPOnO8+XxAm2J6Q
RQuJ9zyT9GU+czuISAewwtgtSfzqI3hhjeiGfZNlQiD2CQhxDRp9KemVzy+5BKKs
Sf4q+gLbo4QrPnjR+Iw/MtMXfpPJAu4zev08UN2Uvo7ID9D2I0DtkmmaQCySvcN1
prP0AWMKWfSkHuum0eV/+vD3/+m4Xri+6KgsRHTRwDXIlty3zbGW5fAFT56j0Vm/
4MgnBdwh/hZ0/kQXGIPsDt7J2WYjxEfWG3p1rmTDIyKe9HX8uuKE/2AvbbrXr2Aq
i3w2K1DztQlxyA+dc/Uk89MWfuxbtSYiNiT2RHR/rmc9j4fYJdBPur6/XQgypkhu
KsUylX7JucXYlMTmAjlyA9EMvyi5J7ruAxkghel54tD/ICtZDEC7eMNtCGmIthVE
S6YMUGHfd7hUxQr6Gkm74hcIhrUBYa7Venu9tfIgjbREc5GpGC7EFBplZcKFCvYj
/Ft2p6nQMF8XVU8ndQBJl44d3d7oD/16egdLoki930IQBA5IVMf9lpBiRyZNAKt4
jGwWuAGhdWLHRQYYS56mNEvP69kufEeaHzJX7GQ0kL14/zSj5P2EW3RXjztbtOjv
jb3qM9Dk4SxQQ5HYCPAXV9/+2s3dJTv5YxuvYMJdtJ+4hmO+oDAAOc8VNoDdGud5
6bHduWxc6KXCUV+rUpf/ijhDCaUQ4zw3lq3Hh6U9V6SBwUc9BY3tUSI4+hASCGlp
JRS3snemif+zfmzV96VX72dQGvfs+hR+xBhQGjWTQdZ9l82qzFaWJfiITFBX0WDt
PPWTVghzshq9EbpBjCexRu3m895VhzmtAMcE/Eal6Cga5qqtgTAOBL5nr+meC9Qy
C2AnK3RuYHA7FXe2wzCs6ixbvHR8yY8YqeNMPTPLHBWRzx9XM7WpjYrfAD58UD2U
1+66QVW9g2JQdSr698F+/0MPd9XlY7xgms6zbteEnHUZRYtA9ciS3XtMsEMPRcdv
MDpLdavsvuuWYaV7jBZznov2n9EjyMCR5+GAfVwv/C/EuuuAeopNFUO2+aMeWiRL
IjntR6xtIm99543Qu8XFRAt6U6s4tEtdOhZ5SWJI8VkcN/NoFP0NHmO7j8C11oqR
s/d0pCHOEQSOsL8MiF3ukm5Jkpzz8K0xuMA50urCiL2T16A9yrUtfBL+LUWcckiZ
ttO0geJKgI+iiU7zRifFh94iXsKVi1ZsVKeJu4mcKeHFfiY44QM31qsreJeApzFG
iB9b3PK9IPpIKhbf6Dl9eWNXVHWlN/JD7YjW95dQPLqp/7xdhcuAKozdnS2J4pOY
swZeYvIwaZw2fqMKfd3VQtvcDV4fLaOxR1bLrYucmN8ThLljGHh/V/YmqS0MFamD
iizdIBNaVnganvjbzMzH1ed9cCLEVkSczWb7bnY74I28pxP+nZ1t9irjqPf4HV4S
7ssFbVnHr1snrIZ4e8AoONlrLE6Ayqw+5qOPBIJ4LuqCfF07NibvfMouMWu2v33x
sTXqfgO1G5E8CtYvt9834PPY2a1gAHxFkfmYyvWns/HKgngAAb9uChGESb3qI2Ts
A/TudFRtbAvbjLdOvD9K0butnHcAcfHDgx/qXAqxX8SLgBz9NX9lk7oEFrWe1fvj
R+/DgGePAgl57vZxG+3OfP9tJWaPeK1yvu27qKxXQeCUY9EKNbQo5nkz/DtFjV05
tk6cSFCuHw3KkHJJeh1Vqoksu8SvVjBo05ouqjqmn9Gk4D+8KdS26/DDCVEGPjA/
4XRRYLyMBKAw6UR6ISCj6REbTX0+lHWI2Aeyga8Gpi+dLDH5txGoSldyptxwAEOK
yOF9OpXi9GDAyV+VWdKD4+FnevDoDWO4eSJ8Tj1GGewbagMxqD6oxR0qmOMpSfzM
RYNFU4EDcpLZYJLq81CUkZbzpGtLR7JleDuxCaGOJYOAtwy4/no7kZW+6sfJGqJx
7HVgYcMOI2b5UR7W3t2sTx1Ga0so+bV6uodIdkXhSEmCS2mntqo9iUBKGK2Z0pYS
fLbMNeiZBMTLQfc6O2qAfpkVWc6JXldyQ6BQPEy+covRfZGEKvHdZxlzuy+bzPt/
nwtJGNrowAw52hU3daaMDAYcfwbpKg68NUUaerQ9XXUAjz9BAs9bJ05mbBT2fQFr
3eNhjkKB0pNP6wIXkrMRz7Hql+Hcq+7j6O5mfHuZzEXD5BiKoN4V+GuQP/wnOT/g
BwgqR56OcosyYGtYteLo4Zd4pD4v64wkIQbnyS6jlESKjxezTfAzFACXYz59Esdc
Ex+wrcBHiG9BwMgt1OWHrWkfllsrdQ2Eyn1bFJf2EJeQttOnLcb0oCZA2rvt4DCK
CAu+75O3pmIoBYCbZ1yFuRitKpAWKSBbLkedj4M+eXNY8IX15FDEG1xw/pCpPZGr
gMAX06Ho1iGIIiZqCMp9zcP7JGK5nXkCrG/Vgm/YZCFmCa4bqERX8WSgis05b4XF
FgfVV5944LAssSbEMSvxFBl0ZFTggN66Z1idO00/xz3qOaGR3b3kymv9d+9uij/H
A2xVkSK4gMIDLDJTaF+K3o4eVtOiJUlZp3KONyqtLhgiZ16EkX1HrTLkGdPll29U
2VtPfUY9Pf71CpuAtWrPYiEV5WGrwXm5O/7v8Lz6RGfziw0sAczTADG72jc+j6Or
I6OB1DXEylTLH7muSWMru7x0tzcxk2PIA6nj46RlVnQb55NfWhZQbsj/vQtEI5RD
oG43Jwqn/7w3x0/tnreDcXnZmGcXekiaOGRFNcNlpo3bNQPe9urQtuBbryIa988S
+1e/0O2ybTBLyVUj6UioggvOap9AcuW9Hc566ruLiTODSL3kJqNEu7yw1HmBsodv
jlkzuJwER/vMCZxHInhCiQlpKow1/SpKPgQOrRrYycftd3OuY596+pKwNzSqiGhK
laYudbsTfop8CwgtV08/80/7t31bYbHBwHKPmoJd/166/HHui5c3uy19j1rUamV/
MjtC1X4ISgS/oX+02diyYFxNzESI40WV9VYmTzz6zedpuDVDQZJlivqfbwPvzEw0
CR1wqlQY9Ixu2l2QVdpWXFEipj9g0fbmkIQCSLdO+AUEfi6gXMOI8Gm65t0nRXvk
9ZfqMIL3fgEWuXlJTcebx2IxIBYZ7YQQ8pGwg2mOnYn/JW1fOS1Fdqp32ubytFQF
hW3J7H3dQ7VWxTRqvh5ubyQTnRICETQlA5dI8k4iIs8wQoqv7/mhI/TSHf7Vn9+k
wq48bf+B8mszz38KeuTkO3xWkE1NvQDn8lTKeRg0tKNG70fWRZvrd3VIyOFD31Eo
0gGuuph1NtFX7QJWz+eJut80t9Ew+h70429XuNNwYHEa0ToRnBiuNwRbVlR9t4xH
nC0DMVgkwsddzRaJtgieLOiJU1gPrZNrWICzJMgw6Xm/hLEIj8Lg51nqOSxCjkMC
Rr3y24dy7ebe67lD6iYW66YSMxtjGhioj1zWWO+E+5nnXV6n38z6z4JlrrfDTjBO
Y8I7liNWzmRbMaPVsntlSNCp1vyxctbI39pFvznNmEimGjkV/98n9gUftWO+NFG5
z9TiJC5LX7X1WaTFLRzUIhW4x2DNYF6E8BNSY4fy4dTtrzjizLulekpEdUFBfshM
WmHzwP/qw0NzfTBdA0XdKGOB5qcwDdibta4s74WoLM+W0duLmrgtrGZwqLVW2/u7
Hpa7A0gLxHWeMZF1Z/YTwkuq9ZFxC1cTJ2ntIxC2b/AwHRTYgIqLpg1271xgHVBJ
nYo1LQI0Ku2PsNW5tBx0lzWPOMVY8uaCK/daCBaA4rIGHUBC31sL4u4Li6daH0uT
VZjep65XSzqdzsOTuzkAIxOlEaZQffUFlitBwlBVtc/SWm+XccQFg+c0q1h46MMu
0rIpLWIbU2rMYiraZQcu2aIlMJ8JUODUIOLPpZUB1ArbY9mmvvl+xNIjtmU8KDsv
5jiV2VPFgkWvMxEXGKpenPCCVx7ZQJagYKl+Y/JT7ViG5k+q6WyNtzI1m9NNXDrt
SMNbJpKMY5ZQYbdhcdbF8hWHfcfYE8wGobjfTLmZ0/zCrYNNlNJKUr2t/6WTF8mZ
TrQ0zC/+XoAzA7KtzbMcOBOIEgUi0il+zRjFDodo6ZTZWMuJ0mm+wl/Gzc92QZa0
CUD629yBTd9XPR1Xf4l5V+XscUMzvmjRbifrooLKNyh4g+8Ptv+vdnVHNEPleTy8
eioXnHvr8AMAV6MF/n/ylnMruLiTO4KQsFs6Du46Gy0aI+4y+VSQfA9eSaCS4oGV
LKOPmLQCrdQY0GwQvXc4Zb3GsFSBbn8Zpf3tgxgKULd3uYUiwgEgPvU6b9yfcyYF
vINKxVNsrXB5G57y/xCDFJynXauStkTkR60qikLjtGKLCzZ+PuXGJOKX6CFkzjOg
VPB88L442jv5vERpGcW60VRi9uqYp4Rv6gpl8NI0teZ7dAUg5jElwBstYGOYFDHd
ttG9+aNaw2XwjFYLNlD5tE55xlLHbQZ8B7os1sYnQx70hsEMAeHmrmpo3kGk4KC0
c7wNn/HQTyhIhZQja+N3Wct6Lhh5IQzmz+KMNvtvXFenk7gvaQUnaT8cWqU6yxyb
s0GWABkqVtylEY1EVqw2LO6/MmybOFcaQ9vQVhbdtJ/yXFFgZj5OOer10UeDD9v7
QEv61C4amzfNhHHOXmkaY26p1j1w2X+D5/XGlFV7KAaV+HNgCNo5xlzNind9CTaH
BMZuB7MI8xlib4DL8B96IWFubOC5AwjNCRFDqPZFlBG5xA21/HBfyVfgeo/lOGFN
1NLQQoXu65OTets51ZZ0wipOdplWDxp/Hurnc3/1TAqkNFOp5zo7Bkje8eANWltj
cbPSerhp6ZWOgK+RkRVTaoonMRtln3cS4qzSQh8rol+Aq2tju6iPjzR5J5KO9lmO
/p+dSDXl8952z0l4anPjGIOtN/wU5oDmbdwO6rEs6BcRKhFEDxPemEN2WXKMHboR
YhlQ1BNHQNAQuhvmB1bsFWntx9b2qezXGGoYG0FcV6Dw/yCkqpp6fwj7NhpjktUW
7DAJbDdUZI6e0ivCZH9gXXwqI6zr+/YeXidaMxDH+85wyZRWS4cWyDfxYZUn+0BQ
teSD4lynx95kAUbtuPj2bgQweKl6Dscwmq54Uj2xfkBQQTnfFGPsxy5ivghQw62y
EKky/D4I2bYEKVwKhWJVsEZKtl5LXs2dvKjzkemEjWhbs+/2WwkD5vgdutjN9olk
gNVfiIp8tacif+j4MWF1IlwxDBrQfgsWvw6TE64zdYWfAir9lDGg3OSGhY2epqcZ
ahDPe2FKHagdxYU9622nSOYubBT2J51dtGoeoDAKzcE2lVCmAXjWJVHKmx5eIu0z
ptC3brBaDJq0oXVyDsAVy/yQrGOqULEVQjZdpiFE93z1Cs00f+kk/uubr6rU/U8V
iwSIXHASVy5VlzijdnH4gd5r9bnmyzvfsGgPYP7K0Tz3pGgD7phMLGxfjGoL+96c
nJ8lvOQLemure8MNt22mAXhHK4+gzXwW/4/zNbbxLfCY1u8dfmo/ExQZ2rXFIKGL
XWge/3Aw2FyGAP5Qd3KfUXqTcydEfFaffnDk7eMMFMSB6N31KKHfDIWE0FQjZvwa
sbXQyZRXetqV6KvDKNKBkH2a0jfjKUSck3DOUc7eFeERe3NDk3BNNPlv9XcYbRNk
FRNS5ybEPsIBsaoW0CxOuI0RiC7rwcA1aWnrB789oz9WWI0mI0q6bAKjk1Nq97bu
ujZ6mG8P4QdUbhsBLsxafu5/cwDA7ghGGEbE2iTzL+HbsesCRZKsnyMjBxw887j+
QOf4ghbNDU4eMLUZhmevvJchrMLTqvGiSR4PMU75tT8G1I+Jz0SJ8AccZL0Td9AX
PkE90VUycz9tOG8Slcf9RgikoMl6GLHpYPT8PdyqQX+3kRUu38MkfA90wJLT8ZPR
+UG0oOH/7WZyvl6mvTUmR395JaJHlOWACa8hJPQpWEXshXJkGSaO8KGf2s1/Vvyc
eAOXA+xPUyzLlKnLBPx+b9ZuhZ4LVpHZ4rxxuhsWxU5+VXq4PG2FN/PhQxMTHsOY
hmn+Wf1OqKQW1ODRvOiPOUEdVqFMc4FktCbSiVXIIZCpQjKStMaFmTUHUz8MJYOU
UqCzsybyLvlF+L69qw3hu6M3VM+X3/EQkryDyZiEIyqkvz/ra0No3FQ6q/OnMyYp
s6AQwkwxrpr+3LqyPTa0mRUBygqnTgXguZzUnR1KSuevaweGrHKGH8N/PuPs4prd
wif3zc2yawPjN6QkJSrFmo7U+ykVChLuCOE77iWz86WJUQb7qe7asAW7GBzSEv6h
DwaImk8cE+SspsTmAlMKPtd2y2AInkKr/Jl5QG4PBWJOMDg8+12OHaFDNkPKGbPK
8qqRSmFbg2oEWCeer1MjJp4H9T7oatTGNoS6XblGmpCGfcT4t16KSYzCaYKp0rln
Zcivyyq9Up7vBryvdfziAnZWtGPVV00MzBaL8l1CHNro1+GNdSy9xIUfYsG/zKl8
zMxrZE+DphseRb/Kvqtlwd+KMvwep1f/ZbWek0r6Gg98EFKKd1kZXANXRCSQ7oPS
ZcAK39LamCFiBBORQcjHt3Wxu5GhTLqced+iCm5F6oeQ2yQvnTk6WnzM1OqmhMFX
2CY2S5JYp2UjOnpmuuX+K61bXY5f7o6AADjWHm5iSXvjfxXxZ+OUsHSYLl4DtkM/
kpxMNKFvPm+q0d2Dwwjqg/5RLvKxTIWTVh8/yJrF4iGo+gCBh/y6YEpJ65XMb4vb
X0NTByk7NqNt2HVE5KlUPrWcLBQ3edHQOGiYmcftsqWtKjtwj9lgXLTYt3gZeX5V
ywJu3ltJrnjU7qUW5y+PK6H+zktSkYWwnX3hed2PKXiWlKL7F5Gw3RI3/VZ1XOnq
xYzHr0pd3fpx1NgSHm3m6NBy5qtKLee2pKon7U6QMsRssaN/GWoGZNcB7G+pJUH6
NBJ58wNho1lajCBLtt1Le8hKbYixSs56Na6ZWkVYCq+2XNTWanmEeFNV+NRvz+dk
Kex1ludxv29uJpsS0S4nqqUvfIRd4DMqwgJpgR4WjGomtI+6BGDFp12c97+DsFYu
FupLg3PZPHPG3YDxoTnpnWtEbJIK9pc97tbhtR0eE411YtTL5XfokEudrswrr3zI
WC99GhaOD9pKrrotIwsbnsAeOiO7BpbCEw2Cy9BscSvWfFlbWRsUZOP47gqHH6wD
hNHL5fWStGk3ums58bElvX9Px/PJ98l0RX6k8SoB4oOp4AXz+cD+Jt7NC9ZCxnrX
xi6Z6RIWe7TPBhci+s97Go2NfKZ2/Uqz2fdI6F0aByJjHDx9Sbwxw4R985APEGpn
p+jeMWwayiY6CuNlL5rY8vEYarTRKjYTTA9P3hItV6Un99cN0JWwD1D1zEUMo1yX
3L6qr+qsElyZZeUQfQITtvvNYhzmBDruonxaSxSXog5SuZwvunsbT0DVOg/FqcpS
tVRp1nJwZXsQcAONVDVwzcebBPL1Tcnoh5SfV4BgjQl+0KiXV4Nh0QBPSAZAfunY
WLBIvBFX4eKBMK5rzub7Xpb0ImgQnpLnLUHNG+yNuKhWZTrUVpJKpuLyZv3GPovd
Eso7K2jW8+NnGNCimynMh1vCcZFfGuveUg4+h00U1VH7zcWi6OXDd3lo+U0v07Ul
lCXLnNf33FYD6kKMKC9/ltQTLuSQeZ/lQCeUwi3hEQaeofYL/FsxR7qmnE3qVbV0
JU6lT20mzfh9i4r8BooSKGyNwAxUXoS8Ih9fYq2Bp7aNrkI9cR8GiWsYbPn7yQ8H
8z8mLcJxASpobmpRfgAOJyKEEKMQaji/I+s7rUiZGeGWSSqku472pPJa/c8+So9w
ZdVnTRVyKJZU4JZNFFkf+OVUALC1U8JRf5f7SjO12bTjyIXVQN/8S57ISQCSJ2F0
IkKHRstbQt3nIvDzUBJ46x7mLx1VPmfknLEKlHw5/ZI1tSmBOZ094R7aKeP1PVCc
71YlubrsHR0eVqLtqZcPCZaCOBj5H8lGhZ8j40lzEPQMuUlMr//c/MP839RI9E1Q
Y+poppodzMrigHDHqk7FqcG4s7mhLOkB5PaiDDYQDH/2IkpQlgXuG4ik1mw4bi6X
twU7Bh62b5enBIM4GPzruMAV03MuQ/f6GC3p8MI0wtykFHS5eJcj0drg1YSEzG0a
Gw02boq8pT1z4ioiU2VTinCiCPeNfEOxptiAYvoCzsRy3z7XmE51OyFR3t2HG/r6
bdwsGQsYEzlHDwpB52Wb/t/4/KXvOr9uC7IX8IX9g8Iv6S3UVW5dxkwqbzcAEC+O
1ZUiRkzaRMaVreeLKVaTGi08RsVuoOEIuRuZv4fysPogrUKuL5PePsSOcU8ZHonP
L1+QZ9j2+0v3K/0pO8syIrfHTFhUQfns2pwZTr2YKDq4fZK/uyoJwJAgdsfR8aew
6QNNWq1jHHCz00x68rEACwhVDkUhcnBA+GkDHu3nu43fF2Pj9+/dLDrDBMpt6c4h
frMB3IoNE7NtaGf4QXC6MOolbfQ/zW8P4EfKb/3Rzm9h9j+tqbO7gFibbRnYc0pm
e9Acq9KmbK/OtMaUWHCgM7sImMLOqxh9GCcKGhVpQQBKVP7VsSn1eth+cmm8DH0z
qS6Vz8uQXg+ir+yknONlwNYek7V34XkJYxL/WmJoFmHNVCelGr+236P8TAY91DnX
ce2vMdbPEup5KNkOUlydwKTngLh8TuR89nrrynJxjNCRQsi16nDbgtaTsaU6MXX3
eARfopoEMMR79xY60+7KVa2yNeDWPpaB3SZTOCxkVAdRj3AACNtYvdSRJcU+kLhN
y+aNRz+vByw+ztM6/EVcGrNLkTaomjMEpKppXEgwA9iF/vXmIDYT3yGy1yUChfWV
ODwA70ZyyxOpmtdRrqLIknrjZXSDoiZfHfUE2GyCpPZtgEPlBw6nk8q7zN/eT7oN
dUzmL2snGJKZiOLYUqpCWuCqt9PTa8uJaODn4FU6w7JfP9wNcCn8T3XTTKZAIkxv
F/St+EDsTtz3hqayBova9Q3oRC71rkL4OAWuVOZDLZ5Rz6BonImKSURMb7jTLcIk
SJ4svDeLoAsw3glPVbshS+fXy+2VorkiD/o2yb/wFOY895ecHGn24f7uWDEg4yQG
k+qlayuvhr4X2eOYzw12eXBTQTA2j7Bels36hmW6EA1fDKS/zIszuKNELrLdmVAL
QfhSBlZU1ti2lfOGN0l9z3BiYqGNAmQrGnREJk4V4MYR8z3rpQCwz5rfhGpyuOpp
46rA993g3MMT7Sj0leFTFZuwKjhbDHHcSr5eYYP9rQ7XlAmo44tINA6nlXpM29jn
UIUZvMc3ZNHeiEBQtE7RAPonwC6cXdn7PSi+cpRH9IKqJioDa34YCqiSs959NTzW
etv7IoDNZ55dInJ/JO0bPGDQDnHh9EKyA03p9mnaSj2nPViDTTQmcIhrRDA2saKG
GR/myPJtcE5G7z894OcDucXqEl5CoyfhkQtUZ8sl2KASeAd9LIxblce1m2QEso97
nBPTaISIkGxVoOrG1TNUHzlruPoFxt5DSONUIEENJ+41/t6svLtlyg7pKAmrdPEB
4HywcOzQEjQKibA9Zic+unkYQvWfFu5vJwgdY5+jVtlJb/cEBxuTILxnviwe76CI
hWNQwCYjmfSk56bpiDQMMX/8Li7Ki5AWo9wXOz/q2VMSjJOajXGFE3GlyquzAVj5
9mwLqFJfpD4MZHKffHEhbITVUiUW5U3SwjXpELg97haiimQc/TVEAKGfh2t7Tcwi
a09Dq+onWHu8Cr5enK/IRetl4ep2U4S5f0cbnESQ412Zc+CFLgHZTfyiwCOXQ0xK
LtAW0OtUgMMCeHQ8QMdJlEZ+4RwoLuaocxtsuH387p+Wzn6cKi3nBy9u2XcD57bd
8Y6wDAMij2SXRTPkIXQwqqP1DGC4B1mNMaqo5CzmS/zhAbD93CIyI/7fNQYlgFio
YOZZEQy1JAoVXKEaFqBPPOQJ+hsXZrBpSimB7WiEMcZI5KJNdLBU/t15mQh75m3+
Xb3eHZ928tqLgVQBTMLBYpNeTFEz/XPRZihgXqZ6b2fONdMdZ3VHU7j978czj2Rp
w0+OUAvSs9nrBHpTeddvW2uuhPbITY7U0U1iqOUVyNBckj9UKApug2PxqsA4BkvF
2PiNsYwGhBPum7lU/iqsRnAXuA22b6oCtdNGCNbVk/X+U/ci2Gsx/2iyG3wE+OUu
bjcrroEM/onWnwyl479qWicFGRv61XSGliZ8xfZ/G/z1vMAsbtYw/pcPZjYaq8Bs
e8whhyPvdsqHRdJHjKtBOYk4dSTPz5/UF0pf5Z5RsnQ8P4mdu4iKq7hE0Pk5h2/1
/ktwJzQCrhUetnqLAMRGyfG+u57yquFup9AHRHKhcbHuXkrFYLJNe8RrQLKbKcZf
0xo4g7f4OYAYx84EDTRnJvl7iBcY9xg2qXulKRWWCJyi4Oe0DJkqATfqjQkIOl1X
ORRDjO+zHhRWXEDFf/HK4Hmsep0l8SJzSz7m8ZxPonGdMppN3bMu0RL28agOtwu3
vgSBd7MeqIHQOv212Zunym8i72ENHjBSnAiPWz0F8BQZLy39xcLrxNIbBCLnyiCQ
9tA8OAdCVoVzhBVU2j/wouIouqX483UGu2m+5rBKpjLXywMLZmZk+OzSkpo1tjAU
Uj08bpFNn2NYbcMbTchZHZeIE5WN5FQ7MA07qirFUE0WOoI0O72bW/9IH5csnjuh
xBa6bBM4LIwqFg9wbslStPLSq5RKMkIRfmSMJhpxRTRiuVDWyHr8dRpNuXf+S3AE
FqKSKCgi+iJdFOTMzg5bT7mdfdebNSq4Kp/4z89F3XID3J5B542hmtN/88K3fvVe
jf1PXX+IDnWeicGW3+9dtjQvBMNqpckYImo0RfKfXRlG1Ww84EKG9uDLYd0lgtLL
ptdsL4st/ps7wFylESHFiL9il+aj2K39zQlOYQSBPuDbmox+K6bTSkFacctG1PUx
VEs3d01w4fxRaphbTcxQHpZHE9zbWkBAfv7xOrZrnEo5EWKgJRuiGb6+y1X4Wk4F
AVW1tlaf3Sc9mPPZG2Au22xL0O+ThRQLjNyl58NTZsh9EKpYPe8VIZuPBupA+v4q
nfHj+/oIIA0hQSZ8PG5fO/ozqtr8cfGDW4IOip3Wbcgtu5H0LraqcVYAa4usPePI
KP8WmWzm9yaxVsgQxf+fQCCivFMa0aWuRY7GMGDX19NJk9jGR1T+mWqkLXYiZ8gE
YDiDDsP6uZ2pxPsvoXvpn3y5+dP+6xGwjPVgm+Syw08V0IEpeefOUOOBHsE6GdVx
kCaHjH788gfgvFHVfYqjD3s76pRr5o8BXqjBQ5rwPEpuFBKOrxletks8+Hf7ASqd
FB5lXiRSAZX4Tk/FA+4dkvEf84DOUw82z1xYs9MYSQ+pVznwn10s98AGS1wnII3N
qumxZUc1zE8A4ap7XgBBzj6PCkaBhY1ULRp4F1uwSF3pS1yNL6whc+BTzBIg+ye+
3Mc+jgO4Gig3zuFCUwfGwIOl22Z0t6jvoKLeRUppwr/ws0/It/BsBnnLvNTm0xf5
FS8XPXtB1O5buJ5ue/6YabvHJlWhRSn8V4kzeLlPwRbetAk4vKai+mPgbzjx4ckc
HZyQwmWYkGeUkcFbnJ4pqZwAPzDwX7+MEL7PmAnQ94bIqBiv434haJhjcFwQ5+AL
nVr9u/5uiU35nvnuw4EhbfQYBQf2u8ggKUJ0HGcrSGS5aRdSSOeMgLLr33HIH6yl
ZHTTuIiVxNYYSMLoRFNjfY01/6EqCn49tj3Cq++sNXpWJSoKbssVlRvckKj8DuIN
bbgEfNILUGcSb99R6IzjAk+b0nfWq1Rk+wfT/SOqqy2FXRj9zReWQuPBqFebDTfB
wkrzq++7CJUcsEAXSz/lOi4dmchv+qV3W1r+7SUi4HA+Wcf4jWoHqV3pDbnMtQUg
lLspPqxUqP7QbmcQwfOEHFlFOGEXO8FIAEwCMN4QtKhRfSYQcDzBwqUdUsikpFeQ
/MOykkSrL73nzN5axy7tjOwugG54UKy1qHRIAN/CrJXDroToe1euqQSx3PfqKdPY
/3sWTIESR/4zn6KLDPoLO3yD8f0JVfoAbuVsDOMH+Lid5jTrx9g6BRumF2iy/WHN
O26E68ceGdK6DA/sVL5kso9E7wZ8uqCq8+fhXtPy95rpbfy0w1CNts/3t3sOoTy+
X3LGzS7sbJ7BnXD2GkzeLZqBUOLdsSIGJYq2ifjwdZdCGIqBlzU2as77rGpU9iUP
PZDYyO4cIcg3L8sLkcLLFPJ8YVIZuadBNGerIaxnlJgC4kfQCjZo4AQemRUn3CoN
4Ex0xPaac1la2WGvZblQT1fI9eTvj1qxdMhp/tdubYwIASS3zHbirzKS5la+oIki
PBWYg6RgMVJvZfCvgKAQGPtVIdAMSe2hc0YYfhicI31qxNYoPDpcROBnL6+owA+O
5zg4AZ35WXMbwv7KN64gdAhVEKa2JIwvjJJOt2rcXZfMKcW+nmqsBuW8gMnJ0lqC
JFWQw+4snSzen0vZZessmh4ngxB68nD0oFc4CJuefZHAeXYOmyF21lTaLG245OiP
OMIStcPzGm7aPDpU4Bf4xj/7guWVhyEOCa1JNYBKVO8xSPFdo7hYwSbekUN2KGDl
7sLIq9LQJmxb74dLEf3z/6SlCErWxCh0k83MNPj2LG97cfqjZq6JfbX2zDamEdSj
+gSevtP0Gd2PFobvwqE0/XsiCzYboMAqcE/M6bjesFKDKt3Y+5zk7X332xfPh4Kj
FWdfQZ+Ak/SMJ5g7lNmK/jPpZArw+DiygRd9i0gfayUHik75UmlgpSvCxHsLjD6f
MDvRqdnGsTMJBDPunLt349nvWZplB4bI1w/kFFvHERmpofccnoN8F4m/wc0OF3uk
N9Bbfeom7DAjaHYKtzqx95RxrH847yMLqZtNwoWrSaNQEFwLFac6B5tuwe27sQAP
HRnZCfGL80XbWV4xzkNVLFJjlAlI7j2YmMjOzyL3sP0z6j0Gu7dZuGPc3G/rWQuN
MeOaV/0P229f55Qieuqfgmz0BhthTae47qGN2VzgnETgzgrLV49RqFVPu4oU346j
vJ+Tlp8n04qapSf9JDxHo3MdW+lQmUEOc1G1OA+CJcTeo4KFT0gJOr+8pOT1Yept
0YueoUvlR+K/sH8Chx4ghJ9jSzrx1/ZSYk/tv0z9vw1O4zxQifuG8NKUnJH7A2XQ
f2TwDE0bwy8C3B43KUmYci1OHy11UNnsOVAOQrCmjljZ2z/B+Y4H4QQpEp48Q8yb
7mblQPiVgB2i0c+1tQbKfLRfQ9SaFnfeOvpqCk6AJXaFiuzeDpdFQq8EfahOpHGx
r0gUkFORT8LiFXjrf6UJY8jp+uJnrc1I/k7uQBuwXNEDhjivr4U6wUeItzzuPBFF
wE9YKpL8AGvQplPHdktheP61t7tGluqVsr3JG//jp7G3/xr9J+qrBAXH9CsTErv9
GS8wsRrEbR6xbQrRRhuL0BCYBEM0+68wf+sB3ltw7KrG1fGv60Fq2Eko2f94uffp
VZwnnOLE2uadr8QSKdSVnYu9EsIVlYGnbuM9jaF0T/3bsRkMBwrpDQgrjQdxo3uA
rPsdZJiYOgwmF+eW4xkWEurOuyFf00IZJs8FtyOe5CLSsYyf9cXyl4NdSth76ZHJ
+NJ03QkOFNXGiRFrqlipyxoxf+RHN9gsIknSoXLrK4FAljyvvhOod0tZt/SZSG/B
dkaWLnHjP9AHrmrTsluFak4DDOn9B58qMQqMbBCetKN+PY3pknH1FcJeX5W+HPc3
TEFvAIkn2EcQohKuWc4/Vw9yCHJq4kkTbjAxCI3xRzRC7mkVT8G9u9INqV2IQGet
vkI0ZEKOHKdn2Bk84eQD1HkVcKCETQfMZZZUGhsmnxwiN7ggbmSuYfg8AicE4X/F
y4Y7ZeCC8pvvkLJ7OrvkZX6283y3CaScC3ozlDNiyhCnej3s4KgrVIRqSNH0aKOx
ZB60n51z9t7fb3AsX4Wk9XbePk42HsrZ8xA7LOnLetZtN3Z9e2SOowtdUNChqLAr
h3LPBCMbMN4lujwDn18UdFR+MEYp4s2fZ6srrQizh6kD80t+A3lSFe+3CQh2j6Lj
SY56iIG33Zze1+xmaSjuuTae8YNKmx+JOqp5rFtKeREADHC99zyM5QnWyxDt11BG
TWE+txixZztsuNRMWahuk41YNFqR/V5vJpEjgtLSVIPAHxa3UuanydkLEkebo4Aq
BleDw7NdZmJIY+r+SQF6fmA7N/vJSlWEYeNYSWcMj2IGdJEvgHkaIUXHOP0cGQcU
1H0XkEizccxOGCmNLbFDTdwvrTWEeR2c0nj9aitEx4Id7NMJpS1UUGtwtuTgtRu7
iDEGWkIGhg8QYkAhsLktVJq9tlSZaLfdOqG1Bc3S78zKPvs19JBN4Za6uTZxWMzY
Vv/0BJbDW9WgbMV6lCmG2VTBCyFnjYsUtukcZGQQrG6xhnpfg9GXmOtjaRS9DZLn
aqnZbRrsUchz5NBQauuNjzhbArROnaNbFlpogsls5/7mW7jruNfeEuwA4k6WJdZd
ki9LGiCf7q/TVEYWyMSuJaIzyOyHzgfTPsU7cZR2UcB8Ui7lHKk2CGio3OkwCYSr
Yy2R0UvhzMQqHsUgE3l+OfPa9rsJYGulP9z922gJNmQse12Cq5vqzq4k5AKMPl7W
prED/7oMny3iPxk+FMnfgQpCR1LKSBs5pMcYMSh3p8fsIMr04EHj2CCGH7mQLgYW
ap+IZrxXX464R9cLM+A8RzhtFad5f2GYkGo5ZDNSyGZwPhPE9EsMs8CKwtkD296S
K2HdDQ65+8uTyTFhe+3UkZ0PMw61tIB9B1ogtp9BEiLtt2wFNvhPMRFJG12lSswe
8K3RIRQ9ixoXkhnA1Rqp4OuK5AmjoDUvLcyVqhk9O2m55fpqpqmwTMOESKQEAl5w
ph4VLxqJp0mX4NOflaAp89FhOjY9D9WKRWx3pfg+VV1VTmFZLW8zmjOtac2dcmWZ
dzlY6w3wuAZb40dek97UNgBSLaDNYW0dAWVcB6bfMWFYCXFQrg+8opzyos15zmEG
YTOjsg0W/0ytFaYO9NTJ6fsa+1UGJEodg+0nMPfDlKtRa3p88kcXe2iVRlPRDJeZ
SuIDUh67ErUUYTjXNVKFrrzbNamuW6oTVo84IaCsniE/T8UuN+379keiuOyu7WvF
NsEYyW1mZElu7tN8ote9veTQ7cgUZoCFPy8hsUQQHwMtVoCPwL6Kh2FJ06iWuXfU
UFPqaDJBFHhgdR2aZ+9DPuglJT3ht4+MPQCe60BpdOqMCZeY62CpccArJqEHUUOL
VpU4Ff9TpuY2SWGmbZ356VIRgdPKgiSmt10bI4hywKGK6P1BQftmPsWA7d9pIqb2
u68/bAUbDAgVVwhe7+HrEoEgzd+nnL2T5NFFnAwW8AC8X8x7zcz9BCDbhVVk9oNR
WXTQ44+Pq9ui5d0Q/G7PtTaROrc1Ft7RBvLzW9Bdk+BpQWPXYCWhBk3gNy2eD6Io
qbBJx+w/gnZDV4tATjHa8XNKcQVMR5++OMqbsNr1kMVWdgmz7f80G7qTwEakgIS4
iNTchEebJrcEoJEGgPe7N/6qx7pAJXwcLC62SJ6OWQrS0TKpRvQoTjfzEgR/p22l
ldCrON2Nr4Tx9q4qnSFS9W+Vx5pOKzHrUFDu7nFGhSIgEC2zI864ZHnaRnivf4sM
J4fSjajrzCslDHJTCpZILN9cVP0Mt7JoPFbTb2Al0v8q38TUg9iFu5qfJ0uqFndZ
5T1gl1mEjwyKgkMFKiSLHcKvE+IakdRdPNzSaAvA51jQc+nivhlKyrYQHJfcr/ey
DZb56aFexSy7ur1Necwu0URVZKx/ESyOOKWKemQnliTk717MNzADry9X8kfhf1MX
aoVXM84nVsCdkvW8k4L9MAmiKHw1vbt9jHp5clgxKy2vk2sWcISK2213tFadGniT
z9vUR2VZk/QQXkAmyRac9FcZkfTTtNgH0L3hkhTzNLVXOCsj86WIfEWPDHUjRPfr
jzFM1MVR4dd4xamGU1lwi8QjdFX4OkyVbjzGHPF9iBXfbKjkv7EJ5KH1coFyFpV6
BDp6BUVXA1Rz/lLpqxFoj9hoX3em7ONvtQ2UlAcclZpvSg7qAivnUynbFopPlfaK
gaXZMC2ErXZJnPU4X5XXu5dZeEvq3Kq64f44roqG390ij8MPEZ73qGbBEbmP22I/
XOskB/9x/105rZfOXbz1zq5HoV2uF22na+ZvWsppXRDX9R1KA3ixXnDAIQ7Gu7IL
GMdgnNVhJaVC7yEmWKtJhLN/jX0hJO0TctNok75u1swXeDTjZsXs0k6DodSdxF2F
3SL8ixxwd39m+50lR94XbeEoGdWSgzq6ag1SlFaC/X/gE8V+tkZcrkQ0OBwbwNqE
6zeTHaJSo9SU/22zlGn6k1xQdP1fTer6Ay2//x4hSDe1H7T306PZmGo8YQqp+L7f
2lpDJLdufm6lBzx70mdOZ72fJc4CRsMkwVf4s9ngsEtMndiQ9TO+5xoGt/qV9LMG
KT2yUtorkNerYc/o0e3bDj51wjfweQqdJbAMiMh9LUSUer9IXaSaQt0o1rm2tTMx
A/XvCI5pExQ3X/laEnb5nf3/tNTX+WnfWycCUxu7RVBn7LDgznZXkXRMi5eYfCWH
Vpd+3bFh8I/1WKKn9ZHODHmwwTQ3OrckTqEShq+m+uDSRAhxRGQPF7Bh/eoV87Xq
RubYHTTxa8p6LrlG00xFTtgU2zLLBNAiQsLVRmInqPjIjh8KQ/Sh+V2G/WQ7BP9c
iQY0bpGuhRnmLrzI9J4O5xYmPDJacPgrVVtckCgxqbfmF/XwLOpotsPfbX4qFaxA
lyOWoqvHYognnknQlRx+NaeSlTFlDmV73Z0wcXKuyVW3FuYY9mic4eZpr/ehm1x9
JZ/UZd8hvJPv/ejHbjKckLJI4flbSdIRfLDe22q6USUA3dIk2EWUd8qWnYqVCdUK
fEhk04CR/9NRboOnh+bhCW0d/0XLtVJncrrdQ+P7x+6KuSAZZg4hoUfHL+Uo6VxZ
7peRW4PdAomJHNwvQMD9EsC6LrauW2XkkTQqsIAmfmP4t9+SJcITOpRH/E/ljbAJ
veloU3Z/V3I3mvOmEnIDzilK0/apZ/6rCSSZr6vATSOCguxIrKI2Pmg9NQFfaEr+
0fw1FOD69cW4vBKRTEAlwF+1bI8Pd3iH5nKxZmuq0ru6Vzk7EZpscjs2+tiRR4+s
f8YIGF6KNjcsAXbmzY1QJlLqtHRNt7zXDQfIg0C56Ynnx60g00Ofyj7jhntX4JqS
ro8wr05hIbhj5mfimxxu0WXzjCrA7JBjggpmBCLJgrmSouFdXRne0i+zw7P8riz3
ntuBfoogf4Kogw1H5WJ4QWkR5346Gc9hCuNb1JSqCSPix77pljaVlW74ikwdOOrU
OBPH5n+/aZ/EOXd73312ZFFQNXcoQZN1hRG8+NprHomBJJLU/7q20ZJYzO3rl6hm
6icneFo1gXG7kAU6huY/pSNazjJKVdPS8jBlsVAEK1EvA+LNfZx22+CDWq4EP2XD
VxaIM3R0JTzbBTv1oTTUfdGugyA8qSi0gtTWiWNqSkMOgFL6lyypIQAiPKd0jE2s
xUFzjyZh2MufmLJyhdQbbJBWKpp4vIDGLcX3n5gpV4L2/plVH+letZee2lD86d2r
2XgGLqwHMdy+Q49xcF8P3+l061yA2H5HXN5ZGiVb59VAS+6Q/cceMA5z3+qkGNRV
+MNx2S2fbDrVtY2f4wRJekb30pKsWGx3HcwU5e6WdBa51nQvKwVraYBVjjBE8z7L
zl5gF0oesRnQ2/PC1F5nVQrz5m4kKOVsWSIh0hoBSSa2ZTflo4P4gqaNGz1QjBHo
13+PejXEB84++EdnVaRN3Sfp4zYojJRbjyjqH+tFNac6TRwIjQv8ErScZKE5OIhl
f+VUQxPAPuU8yvkE9MWPBgTGYjLW/EtQid+hAXNVnrZemTebwYLbC0OjoV4Kr1Tr
wNbeTpE1wUSgldcx/H8KC/BxyyqEK39Llf4oY5ZaCnz7MqIC0jc5AVqq3dVX7SE5
yBff17IJHdwdVSZVJpryDhbkcGNDKq0/JaKwagZeb1oRyiU1/pgc9p51ad4UTYQF
YedJfBj2aWaNmVEuuOc1sQEd0Cgmw28dM57JTa+xqSZmrV87M/pIxOPDDZj2GJss
lP8Cqpzr94DrPMt1ELkLcJuHg16MFr9QizaePF1AYAp6ZDhoOt+Li2QepopFk2wg
1qKkOIiixqgDX4BhDUu15ibHAOEmPFIQ2XDYtPM4wcm9myoTF9AQRVzGJ/LWUMzy
pAsGff3ACuUtN2BKFhMRDYNTyEgnS5GouYl4hoXHvyU60FqDhYd4pfLHERdptJmK
IxdA5c1ZIZ8dFpWxWIwgpeSI/q7iz+7WWf+uUF9NqbNVi/qfjpnIuPgsfHkCmZ6C
dGqZ/V5tx04+5RKUTlzbQXBsAHlZh1n96i+44CGlp3ebFONIuDN9o1FPmcZwSkGS
gX5MVf7csV4e2GSAeb9fxmXmeMUrQJRgwhHWLKbz140KsYs/b8dHxIN/7Psdn8Z9
7uTbwke3EeAmiFqGeoJSYwx+nhT7L+sOYFbjb4LagJlMIVFcYe0KIqarOS+QtCGa
UDVdJryA79BIrjumDmlhQW2asZBRQfQ/vlIHxK+i9/fphNnUpWmoHGILyLLbDLZm
FMaNqbu9X0WJcIlvK50q3Sj2r9k5f8od39R3m0bmMjy122I6ceNN46HTeJOQ6rOP
62u1MbqI+uQlkPhr3xf/nBw4vr8bT1QoYGL8Da3Dh3tcdnE2GPAbPgKlisicqh89
bdhBYXnOiOHobEeWd8DYXkxnmWQeRfKuMXzWuLXSn6xroJ/CqGldO9BzqquIrOC8
0QMvlYtQvT6/BNtOAd19jMAtBJ6o63wdFT+rAM7rp+CgtyLSNRkbRdVDw0PfYpQy
NuDdUtATiipVfZPVA8osuIS3AWrGKmWBB1cQdMi1U8WBeKBL93pzY4d8ifkWJS6p
VTc4EHIj2Q6q4QtwCR/QZjiZHYDuXG7Vj5WTNretW6TJZh54OrGN7mX1DqMGrtj6
tQoMp94KdBPpOj+8vK5Rs6gghnnZQttnuU1//VErEWmjl3qDhRLs0Wgn9RmZaUMI
OI3d5i8h8LMoB1sp/KDdUqOfl4PwhaxuZotfB9rO7Awh1vIPntVfb7dlGr4i7Cxf
zc5stqgk8mdIIVnoXEJVXBgLOOrAPcUmh+K3CaSVp35iyYXmtAV/5vCjrnICIsYc
L40RJ1uoXeP2Zzq7V2l0Dck89i5i7GEbLBbxWv/rViqBwxARFiB05qnQcKs1/fNx
mUGGG9mdHJ00385QF6lzvaluoR34dGm/8NsRw2XdF187HyRO44SYKRdJhv7i8Utk
jSOjRksk4K9I0MfgxCSXjwiZ1o9n7zfV0oeuN1Lfs8K6oWKxB075Ck4Z7vlQwfoL
yMdU0bYjcnqIkiVGc8kjdma+3o3wEQhwwZogwGuNzl4lkRcbX+6275r70KRSaOfM
Bthi/wsi5AaesJPvV6pjfCFX2bgTQtMPm7AkpW5bw32XhL2VJQJm5VxfhqOnfQlo
fs/v+cNuRMkT5xAOz8HyGJJys2vLMKgaBoFS5keQ9/VRPP44SuhTF+wAvWjdWm5t
uTsU3eiZWX/zfkwbeGettdk7E1q/8FD71SezAMGCwwG28H9jKH8lpS0ikhsVfGzd
15JwxUdiSOGXVBG0dIXnAVlnHjph5RsV0uVVXIH4CcqN9YAyUSQpKgz2gSv8NZq+
md512TAWaCl5y1vyEDxWV+zO1XK99kaUhdgUE6DJTTeRXStC8ogu3NcZRM3CkmSD
BOV7GVFGqaKAXKJ43bLYR9rMQoz91Sk4mP4RzBYtIcAoTZhBBm3h1399DjjhgA14
N98BA5lQqprhVMKKFOaf7NHCV91rNxCL3I8+AtaLAzSh6eCLjx1bOzID2wlfnoY5
K6JkrMdFqJGQ94DVkwn0NTe6EwEXW4r+sKecj/9FqiLdU4cE4OB+ZEHyNU4esnuN
uypM+ngzyfUiA7VFQGT4H96REfHJ25nV8fjL5bC4LHU/z44W9MancQZiQNDNvzxi
NREw1nj23WnyLClyGWmA7+TOjn4Y15dLpYL21cyfkLdrVtqLsR6tL8BEIxi5RQIT
+3HlDXbE5rZSzV5cbRGR9N1nvmq13GGBUUPYJ5UuehUmJnCAo4+3RA2uE8GgmGBs
GPCVQHNOR/oz+H2TIvWnC/jg4c8/BJItB587eAjLwVImV2xu+UjHbuvG46fC+nQg
XR20/ZnYyMrzPUnDnVjOscOdlu5aiqnCKXVgWgKFLYGcx/UIzEHllWv53AJwvcw0
MSpZ1OyVmHcoXOgmv2eaRTwiUGDfM/EMlr/PnOSp9rxfjXAynlppmU1ippOIPB2S
zEqr2oQr8CukDEhyHF6owUpRJe4RMRNtai7MPnRq0wjl6uD/ZjvoBLcpB7O7hIo8
EV63yLgtKWZEYaq/EKX9j6Xa7t4PNdHmwQ1vuSaYtjm0q3/0W/FfRTciXErdoT0n
ycF9VrHu1ZAR+FYn37R5VsObdVSKYBvmo0PzwQhoBknup7ouCB3djNB8eyKhXOt2
KV3c/buvRa0++ujQe7MVm+YnkecA10ZmHxdXalN+Hx8jwX5bJnWhoQlXWUOjmBfJ
b0ptmQe7LRrRVmKuNTuds1TvXY/nz2wv8gyEbt2dKV6K9cbJxJD/qCw1eNonLYMd
Zyb7E3ThMv6CyFUQBsjhXmfhnH9dyMFkYS52sASTYJtn0A7M/S+Zwh+wHM9chxYo
/2ZPLJ7B9BZQxKth1thBxtc53l3bzxlQRmUsLOFoCh6L74yviTRzxSSjrFEW9k+O
UmiXYs1UTRLk3k59qFrHAyrJHRCPbPXX0yp4maiy1Bdy6etQLeW8N+0rt4KDvwnm
cXcP2WBcHAPwUmoilo2iMoJrqapWo1q5sGwa32Tl0TF8Q6mgR3L6zGEPesdTqClJ
1db+QO8xhYw98V7R4gzsUbNSSvLJ0HJgY0y9ZSXcYiUtSNvGOpc9m7VI9IZ+L5Q+
T3JnTH4ig4qu3TbjkRK/HB5KQ3Ji8lHXMfHUrQ31VhcAeC9C6JopDZUQ+t406pZ5
0TGYw1FzfttZBvBSec7/jrqJ/1vqoz70WzXfJvpSMkSx5skW+9hluNpIjjY55+qF
pzKXGF7MlTDeEbhV+OnHE+Tw0U6P6PxwM9w6QcIydThojicQ0hBECtHq6CphdbXY
ojvY7tiCBT3sYlgp/4KgG00bQpnThA1e2Xj+whizzQjgx6xzaKlC1P8px9XtaqxB
QdUr5uWfpTe4k0PdJHZijGJSIe6RWqYR1++ra5Ay7h6Jl3k7wJLlYZoNILj6LQH0
qLfBNF5vWV0z2ONgtQzMjHJNGtf/foWg7nD0/ps6sRQAFz56iJdm0pJ/FhuJ9bHF
RFvMmUSOS4LrWI9BI78WppFn3QvLXQ3WxUBe911hHqNVgCJMiW2aRui7RFmwDkRM
CbQW7ON4aIxqQk/A0lpHJxAtx37f0vPRWzZIfS9yldP4rte03/NhfLDSNwNuMW6g
BJFwvK5ifCQTRh0yn7KS22+p0SwoMEcacFx6sIJWPE18ut7aMpN/b+SqaQazkB/a
u2hDRjqMZFEshBxRnJI+x6mWy29VuWdHCVFRYw27H7NttxrkZ2fFj2U/STfdG4xb
tG/BNRc+nzorhRmb2ImBl6k7W+g1L2F4STg/vYRYod0pgeiz1jOw7WaZVwfB8+3I
XiK3m05B+i5meWwhupBhYATTBKSdGakVEe3nTGbg/C3FK89I7smpfr4N96iH4Awe
6sCpg6+kxnbUKmxAgLch2nVQvtEEEiOSTYdns/Dx2tYlG0533m8CxyqxE3yg8NSR
+cNsiTTk2kbPe5v/I5UwfoiE/MvnhQXNgOK/lynoW59+cG3y1BfmyG+bW8QiMDYd
XLzpCHMqg1Cvqybv03b2yRui4duL8W933pqbaPs4YM5TGlyTh+dhEFoxdWxCyiY2
QaICRtO4cTOgoQ9Xx9asutN0ylV1mcghPOVxWp8ckNfaxQ105j8h0Bjs4Kddv9ax
XGAIeU1rMEIj1NRfyeVMmWVDNsXNxRLDbsE+0pselgj46jC0AmGhEbIixhArKKAR
q1G92ejxSufWq78/9kYK71HA3YnM8M8CDcvnFeNewXwW7CdXPKwPsd8tIXrLbWbG
NMfeJn9Du0JuspWeKvjSGl6Dxnmch2Gliz1rbjA/ip8DBCekcuW2y4+MFPhmamMP
4PYvcTH7S2O0jBp5ZFIkbWxmb7fCnNtNSv5mWetqwAj4AdO7//osN6hrJTj9UCAW
EDBZZg9+RznKxQBPMde6NBLknDR2foPTMjdB6NqBNUoqkn9pYtI72FlIaSi1d6GY
Ov2xvftPe1UKjfht2ZeSs5dc3nq1G9QIn7GHa5BGNqPP+z8uHtF/2hjwTvzzqvmS
/enHI4l8PzI+JQID4D/37Q13B/fkmRqYQjVbJ/DiP1YqekV7eGBAQ8jBPTnpZJyY
qwmFea+NZ6jCzTylB2qHg2+KULNqMzTL2LELgVB0uUnzac7zZttPAKVN0oB5WNGF
caytSknED+KtaPzxBQA8qxdnXVuAKyHkCG3j7yjyOICtJVW4HrBgfk52gSJYXM/h
KIOx2iZ4Fyp+p63+Zslo6X72JrSWX/GbZKUhjXrkn63PXU0McOJIX4RLbUyglsiZ
ZijpZq8Vme8YvdoDlzontWz5rkDAtFnS/suEfbAiDWeR4Sv18d/keeQ6Zggvy57J
dPYLKCTUh9De5E89R4yoWvo5oqRVfsaHuT77Nmavc+0K512AMfUvzpIMrhqZrDDu
7OORO2c7VouHyr/1t9bUbtFDFLN6J4op4+V+o/yWFrEy6aiRXXOKhndTpny4xgZs
vLKXHczfXk48nfnYoYTPi7J0hxbrmbAjn8noLAZsdd1RwXICcG3i29J4ULNberGK
/U64kYv4uxDV3U7FQiN1QjOfOOxsuv52v94X33hDR1VpOjKUns1TYm+HSy34OzMd
gmuRtlJleKTfNbHPU5gJ8fs3hiyy4KfXaR8lkQ3iU9NmIyqW0uDH04OQ50xXir3/
ozQpRasWO+Nzu+XPjNdHhuCp5lL2PCCszkCW/HjdFnD0GhZXQrsJDZbaA36JyZeY
KE53/fVcvzngTkmEh7jSYR+tTgqq5x/HR1DA4r7ac55geyud1a74eWgI6doT5YFN
l2JQ7bdVX1ZV7YamrK7pOlmhUqyqmtuWb66WZIgVCeR8o5wHgtuDMxOoiv2Om8PN
No6JipRL+F5r1QbxsH5EPu4neHi9HukuI2+6Xyr228jaK+jhyQMI1GFbPz9pkzjG
PfhTvYm/HwkTNFbfQagZ+5zxqTKb/t/TPrjLgWk56NAGYr25k2RtLTT6/FtrA81g
CkpYBCXkttC2fovsb6LQAQ44OS9pga59ejsRAhBD8eWKSCeRJkEF/Eia+h+qGjhY
oGVv/vyI+XeLJE/vpu1Gr3Bx1PgZrE0BOni4FgsLQaqxbGo+XA0nMnMnz+35JQ5n
y8HwXwV4CZZ318UUQFqRvg6dy6StIysKXBjM2mtySPsVWNvqIcPVaQcjLrXO7zpY
Kpsh3jreJj/R/4u/ivLYjqNXQwBXSas+wvBYRIB8pTVIWfaEPDQElZtZJTnRWnhE
B3VGdUuxqK9/+ylJil3SyXhp6w6QnZo0OWjzyL+/QHRrDTe6EaNwYhwpiRJPgrI5
lmgh0+DSTNoFTFmSnucQwybgG/1HwCE+QwSrQHuWsLXcaZy80pM/QUfqE9BDTggN
ym1SIgAGmmj7msm3IanMvV7pwDhVQ1ztQkFPhemiwzGu0BWaZijDCy6PWkMJrPCA
ns3zHTQRuMAVnCWyLtcg/lyJ7nmn7uzWT2MR1UYIT3qZGDM4pkmrInO9Ull5DXeX
oOblKj7V4ULJ3pDsnIZbsf29+4b7Tfcxap3mpvdO57ilym9CW6dS+lMWboW15C3y
JW/zQqr94LpCKI7XE3HXpWJmucQQKWAnXt1lKXQGK1pe9E6b77OKBBD0BOCrUAw0
WFkwwx9JY9f7lLk5aby7RrPLY2I4aP+3BepWNnLcV9/RJbeHgon13+0M64S+s40A
yCMXB5bUxiVoPz64YKIsDwEMGVP2YTfiGPMTJn4lvOP0SSO9k2g//D07FIKf+O44
E1yd+CW9PM1ehi7j78CI60cTCACIpOj5IOc1cRzoQs2ax6gRw/lN+ocC313py5Qi
FnYweOna2eF1DW1vFENGgsksBTOcBKrEEJYgeYm4SDA1jNkIS316rQvT5cRSdf1X
mhyeHA0CmPcfbOUhZOVZKkaB7FyJRpmz5383gUZFdM7Y+HJgRJSXU95xhQfyHln3
9/rZy8/XASruEApkQWr6d4vWeGXpjmCTj0et1lvEAIRDV7WS9yhne4CFpSFQubTq
i9OV+rEGoREsi7P56/a6v25ovKKpwYRJDFZt5oHBUIAMYiG6y5EFLCuXRx4cDoqB
G01li0epgn5yDLSs97T1SyXg/xn+mkFl1XXtiEwhzdwR2DJcQxRnPOptup2Y2nV5
5cHdPdMSqe7brddG6bjv7MhttDtiPXvSIzj4rS9HV79nlHzVTtP+KJHlEbii2nT0
DN4o+R/1swqi6fKfEBZG2ZcwbVuPHe/YSjPW8e6vz+JKNVM0Xdxu28uT5B4/93Zq
W1upNx+tGEe02XE90xCI7AKeqmqJhoX5eSQXMfBajGtDN37DUM/DGU6ukkwnmO1H
Vm1sNmBOcFXmgcQQ0hbIH5hw3Gc+LYtDOtqaZ19GUAq8cYBS5VEqxRBPeUjH9Hug
TVM2jD00Snf0yCbHYkp2KB7jqie2r2y86QWRtWTrQIlh513OupPLxHHbiaPw2LRr
qx9CDc8z78rkhu+zwEvplh65v+yd6RP+QYosHQnqCuaJOjJlw+lTbb3x/lrUCICa
5r+m8nJMgRwRCf3igZOfEJ5AmE7iHlFkv/i0FmWFpTjGZ8BlMbJ5+TSLQJvfRlAF
clkqEXa43z6NTaUdkw4QPsxAowZJFqI48GaCKBflr3Ad8/fNoMsZ/RdJ+yCv6H14
BG4CAM5+/Qqfc3o4b7AbhWwJ6lRKgS0yQAN8AH8f4EsKkpmOMUwwAa/uK5xM3t0b
TStQf0DberE3pCVKchr52qDQfzCmbLzJ7e+QDy7bdm5Mm+A+jlUWlr/Eq3GdHavy
i/lsIO8GRVGRFgM8eW84Eb4Beg5tHyf3igs75CN/tTLQk5T8y6dXeNmZTV9cBhg9
8nXw5xrB4OB3cq1gq7rLB3B6xX/w92YjRrj1tblvE5jy6pmp9XwRx5RAuAU8A2KZ
P+F97XMC4cuKzOhfW76YmpktSPzYajAdkpaeOp/Z2r3i9/AgwyxYclLeu8W+KDnS
ow240MvsQZUDcsb86UGONjA+2lpPX/lRVERJPA2NptK8gGTvnOYNRb+1UARM3nbu
baShmq71UPBBpOiImLGtRRszTc+fg8rGDA0zDpHZMREFAkd0ewpEcDqJ0SOHrGDR
2vjyxafogJOxLz++WdAJ+6eFSyOCUVsxorYVZ3G8Smxv3m9YAYlMmKBmywizv0X8
fjP2lpXQWkopal8TCXOH3UtWLwovTbZc1TQsBgKeesJCCsCsHjj7FEp2g+HYrXTZ
CVdJyIjTk/jWEjprt6bz0XwlARe5Jnh7KuK0bLY/kRM1RQykQl01/3vI+tQizFzo
chujdzdCLyyReGWMaqBhlLMABhYtLGJUemL7lcXUo3p3vUAMz1fEBH4fIF42WyF2
/hDCintuNrNPSBZMOVOE/jyoWxyrz3wXXERBpdG+IADeV8e3WhaL+B5c25wPfAVj
D2GxjkX3693Hs0hEPt6bpkJOJ/jwypd/Tmq5spc7vukhxN/VEXm5s0T1NadzUOpF
rX6g63G5qK9DE4zjcdAXY3vGoVKFlXJOu7PD9yLb8O+Gqg3DJSUklTlj8sJl3mOU
U1xnZw+nYB2pO77iRa8Eyqpvd+4Zpfhtqwn529UQ7u9MdzLmIzPJEb65K8uTNwaK
YOXTbDtqT2BmMH2xwOCIyyOwmPpETt8k3Mhxlle0Qy3by1PsaOh6vix+BDewhNm+
t3cW8XYNQmZrh/7K8q2xFBVcsqaws0qzdCnmUV7sZ777kDJ2ezGIrwh8jE9Hnuif
pG8EjF2C+uHTaYWvVam/p9ZDmtLY+qXaUaQhxtLcVCkK/wxClzs+zQQmzsdndl9a
EBGz2yq5U1Zm8hUAUF0ZRAqUndh18EggEMr2EFJbavXG2vyU9W9ne8kYv4ZHBiyh
8V/58wBZ45e5khzU03JvpRpHD0PjVL82uQ7dZ3sVSu6fx2BOy14LyFouhfZXhe4H
nv+vXtEyQibKHovoIsNcD0I6xBdDAUR+Bg+jJE/Ot/HTAj7Dv3SMtYKI4R+M9Vza
ys5QyCTxpOcKcLOwXQdsYbpFPkfeF4t7ta9HVqSum9Z/tV/dnaZcWTZmiskX9O+d
hpxuX6lCgF4IpSOmQbr+N1qgpuZYdVrMG0Lz8DgrlnBqLb6CK8JUqol40nMcdF7B
+5DCQtB764Uyzni2WCDf6LuEIOZAAA4afJW0KenTKt86L80F0XjCHb8aUcGBiNRu
6TH1mbxaPLugGKgNKm6H2WBINTt6nC/tqqfVBGoiJsdb1tUTVHEW2lOmc+nv06XJ
rC1CDrD531l/3+ilUUL2qY2T2U7eGyyMYoSHbXc59IIlE6h2DAO0rHLPIY8CpW3U
lSTS+p3VYMi4Ds7y+gA8wixt3mZx/nAtaMEqfXca/oDbWm50nl49HZ1at1jvnOVu
OMFW3+oo0taZ24kNyQoHQYsBb747qaQnf9s3Ax8LRoXPJ5S8GaIV1Zh3WRXLUrJe
4+dNj5gUNwn4nbsbluoi9m4FekXdcLaNkriWqeChQpCe0R9YCK3GgVgkVkNGtEhr
SvHsCfZF8wxHUVyOFmf4SOEhLvDgNgDtKEemt5zW9fIPHbOilU+1F4Js3LnJV38D
4Oe7JEfN8tDcCxho3Q4EyP909rBSkeMyKxPzTTcjJA90OB3gBppwcOBQihoNYBhK
d/nsXPAKt1JuozO1gMu5l4ZpO9ieJU3UkWN+XcJY0C7x5fKQbOGo2UoDnVs6LAXG
oRzDC4qZr/PNHrjWIjT/fZH/8O3kxwDXPtngVrjX9YTKICg1SKLAwoa+PrjPIboH
RA6scdYrDm5qQwVLH6uxaUdy+Gmtx7BOM3cE9JZdyuonwQJVb7yCZ92c8ot7HI4a
f5MX8Lf9PzIl+H6Ny8qM+63OwJ7EQ7yl2Ph/18pwz/VTgrrJFYg9Z/+v0BZp2djl
T/H5s0HzVT+8MAWGL8N//V07wUupAeswRlJ+NZ4Sq1ScNs+ZX1P2aO6N0HEY5An/
YzLMGqgV+9MROSlsiUCeZOR6QljttEpcx2utclwCI4j4izWQvzRV7tEl7T6YcWbw
EY+73czNIqMeBS4mbcNT2JjZ3u+Q8VFXj5p2Pq8GGg8vnAVcv5QhdTGdzZgVgsjG
Uz5bnStlIDKRiIxtJMVrRH0KkqGCiENg4+6ObgFj8UncRq04neKEwZanZeigwRrz
LkT5nsvDZcJ14ri291xTY6gCjaY9kjBzGrsdKMlyBLBCFQK+eCKbNL57qCNiGoVr
N9UiRZsQbuPHra33JFEPT3KcpaKwB8UURRQS0e7pxCYUPMHcxf29Nkb72crlb9TI
GW1Xt1wsPmkZIIQ3JP1vjfd8DtwnM1poDVerl2R/3E4hs7Cpo4kVn0sPdujUesDR
D0b8/3CsxO+HoSY0QRFQo3kxBpsE7cG6yDilsPECeBKouXY2UP6OvMIJD9IgrXUr
IeBpbaT/zYeipzcwv6DkBV1FuIeMR3v519TWfDxpjtceIXR+yjRwfKiBYcn6/eJ6
tFBaTQDdI6XwWezXcNySnk1OnzEIri8oaDfDua9EqSdRfEEcfGOSWsLGgLQABL2E
5ET4MaOZ0Qu9YW0yFdzWWmdPVCZXhP9LYsAn2OXHVAgQ253vxkEp5z6Kca79p0qS
TwX3177bAfFO9vyR9xX/wC7yYssLyfDidYNMdwGhU+xtCewX28TRyqO/C9EwS/Y/
IpmYfKvbwZRMXQnAlgKqFa8cM4Eff40erEQwzl9q8jU3O55mPx0krV5o7EvQnFuE
qgzVznQZakd7eXOASDRrQL0NJVwCpO1yeRZIk5Hvn9BxotpaaikV+Jd8QlknPxK9
vjgKzY/mQEhNMv9UDf5RJFk+OkJya9gBWWZbIpcMd0lSJ2QYRp2GRcPDOjpBr0UF
8NbNlvMh5NCqSV7iAJR0Bd9gXwNORVOQ2kRU/IMyyrc62qP4dDqQJgwTFGWwN9SP
zO2ozRYrFyf+/JKkiS0vTf6T29JbQx5ayT4k3+1Lg3RUZi3COKtQM0A450ajck07
Uz3KkRMKEK7f+0GbsvSp7gnd2KNf4Zk/Kdm0d7bQUNiDoWX4Bn4u7P9QJJHokB3q
cQRdphtTVam7mhLTUZvZIP/TWVFknKWHgXYUmQw00CZU3VEbvwTCiFpJcEYIuQDu
O9YTefph/9spV+L48uUmLyfgzYRBUPPLhIQgtR0ktPGzHznZ7mBLh0s3z9bYfOSb
ZJIGTmkxG/wKQdjuSRRq7nnwtXPLLA/AG0ZgGaCcMvezbYJN9MVGTYZxzyW71BtO
RmCwDGTjkLgcWhLbsxgIYXpSFsvEEXs8gqGekILlHNq5WzKEHOOPoh8FOChn51s8
A+Tfy6579cMaSzsX8ert+45frVYpznKaK9g3ZTFbT0iUbDbQsvgRHU+1y5Esh8oC
m19DfxsVNLywoiVI7LPRDn1IV2ssOjR6VPjHjMO4mwFVDHUdtURbC+afWlV941R4
pPLdJl09EmGaPPEJ6woOvfYlt0+x9NmcWpQEIOPhoI3yw7FxaBvRRAkVd99sy5a2
JIe2rRAd5kTNQXyJczxgcbc4a/yzH0Ixy5oPkGEVxZae9aFe8GSwAxhr8PG2FL5/
HkArfGVU1DA5NYUP7Aj5j1Ds3TEb2mSaoxG7AvpPDT1C0yaXdVdPeuzWmwRZsVyy
t21Z/3htqRnD18UyYng0LAvSG59HKkcE2HgEeTbSY0uAkdB86Tn20DtYZK9vHM1F
dPBSw2pncqlHg9zh2RQhU7+1bt6aRu0Tw8AelExUibOk2+nFWeCLceEre+FPeb+8
J9RnOCQ2uxAobIPVnDGqF/xwnnBKmeAu+KNJCcCRWPd6UiLPhKKECVGrJt16i6D4
HuCcwM07yKNm0+nNhmnei1e+LcjAbn8pQLcs5gHx9sswl1DXTWDZwqoRvbQKD130
hd5kN1ZZAsJbnBo5gsrEg223+arJL5c8u8jaK1JItBiBNFcXxA1q2Pj8iqQuKG4i
UCHOjSRJ/R2xO55Nt17lFNWntf3uJcConfZR5yP64CRqrrSvpij0MQcSLhA7frzk
ztsbIaP6hpaF+MAJAMyWB7z56DhJJCNuJe8Qu49tF3HX3PFlZZejUN/ZLsiN1sXG
CXuhN0r4VQWYZVc59keQrySMtRCp5Cel1JtbQsyPXR1hKopxgbDxHvCRpVfJ99xN
rRr/ElpRotIcFhrO5z6CAO0YWsT/G4GFMN0omAg58LMw53+wLG13BqdOimUZWeQv
8scm41gvlbW4yZfq0/+JLUac5+/DYMRbBDYsEDHGZTxUfx3XBF8VVzMWOd8fGhTj
HdYI8bBpj9LKN06qd4/KFb/A9Ukc673r9d+zww1joEftmdFh9dHdAZEE0U3Z36Kq
SMy3cXr38m+pwSb1LnUpPBkBVvlwX0liVlCoiDbcmJfbGTonfgoEParzADWrOTM5
4M2k5BOgfbYh23bXLYPS4tRObww0RWdNVfuC5ZikemUy4Rz2GmcWDrqTGtkaRQel
G89AzNg2ReZAr0J+bS8WZJQsEYsT1G9STVAJUpRIB2h0ds+haZdZIFLI7m/8kHux
B94OwanLtNEd4/iiEq/UN4wb03qsEJB/VoAMTpC1+/ASODexFyYGO0J1xDwRl7Fm
B2i1WKaoH5lecaJefEeySFlekH0+hYE1sbfPHdvG+Yy8MhVss4h1pJNUwBshrLDK
I9IlctbQSjjjOiDTumg+vDU+ffHVBc1tZ9iLhvvVDam8l731LbMmwgDoxMJfj6n5
/Oz9ohX4gZuvHqzYdtjXmoqocb4tN3WmJ5faEEIrVsT7Z/OHSGaSj6cLEbraeGdZ
LYRpw4gUlbpxz+cb7JebLUnIj4WXFH0fQuVthwJaUgKVPmMl/ETC8Uc1acDneLLW
lW8tWcAzVK2ljoBcevJ54rlI1DAblp01tva6rFD7JaPtYVfXNWzGgt9VcH5uOp+F
GEjTEN/cxNGPWFdvheF1Oje0yBV3bSRviysiTSoOPvkqQZUgE09ULxJi+4TMe/gu
mDz0EbxFjvh6yont7L1e2Z43XDioIQjKF5rgE7VJB1FYKEd2O8jQupSgNtZzwE7j
G8hqOkkHMJG0CUHVzyhh2mLSDX3Us8DsBDfJ2VBuw1yrunjHP1vOSzWO3RIf54AQ
E4BeFz5VVPO5SOV/Dqzx6D4t/GFJVJTsXshgql7WsptVi8Q/UdQwwFvMakY7hbbT
g/7waaSIQlqBHPljGGtYXw3iLefShee1HPLs275FK6ZoGLvZpqbPO6rGgIAPh5Nt
zyZKIPh2/eV/32BmmxFkBgvRslZI0R9f+FccQyiE4qqQ9COcDvDpH7UTkwp7TU0b
r7MkYtEUtnjvWgiRu/Gqrq1ytUmUehPSmuEE9MWt8Caq2dRtQ8V+65/huwDUnwf7
v3eiVb4re/VeIoS3/zlwk2WAHHNxT+pkV6J+94uEPzyTVySaae87jXshsByO8t3G
FFolTihVOxFFhZWc77kN9pmU9NUe5xyLjI+MEtLjh/yk1l+NAMxZKvHNqaJeSzx4
B7jgMWp8L5of2omJ8WKOMsyLlaAdsHtDuCvMIGhLCVjF2NdLvzhRTXBaIM4wUuf5
w7PPZP+5EbzRoYB4z+/RgZibbAbTDStwgVzaAOehIJqHDWP+mou2UdKkpJS1HRsm
K31hvuEa1JvgN64O01ghF4zD9CiQdhPiBLmHEA5HzMqNB4uyPmbid6OABc99VsCp
kYqLc8cBD+axHlD45Q3aY6Y5AYmPw2Z8kGE22JTNx3Y7vgrINcVWosRtcLJC7iAw
iWWZAy7cJgcG8eLIQ2sbeYMdmB9fVKnu9HbXHDwirVmkP3J7wSs4S4XM8xxiY5Cc
eTmybb6waw0v5EU8dPgVI7cPLMpJp7jjIYufns1as4g4xvirrO1C/vKBHi/eNuew
vi5pAdzrMnhAl8+hht9RJt9DU6zuMM4L+0+TB1j8xZ7yQffRr04BEr/ypnsxlDGs
4Kc0LNMSsSq2FO6YYpZhzLLbT6IJZzu9dM71xBU+/6bMt0hiFZawBZfVMIzuG2ff
5TxL42mNwHUr3cYkXTUmzJRmpe5JWjo5yBN6sk0iWbcXvUrUpqB9IfmxZvtnzw+m
GBTVWZNg+DiB1joeUYsMqqTF/V73K2nGpAo4gAA2qwXzqFMYadaN0mZ8NUlanCOv
s8tsCBlAhMRqnDdSGA7W9xJ+/eysuvVJYcEdDH0TwZI5Iv3dKAIYV1KLyaNMcl6M
O/+7EjWlSeweltIPUpDBGzYN3/Qbvj/qCnPWP3UnFXmLhrU1eHkLhFSzY5b5tE/O
0c8iE8lG30OzktToIkLCrDdt3uQ/Z/HkrPg3uxCQfdX3lYbzsSdOW6TcIY/4SSpS
i2BDD6YU4Jq3EKIn3rqJDbXT2ZXAWNWYk6cWeSr+QvltvIOFVucviXmKD+qz+GUs
teuYLNB9V5WWhYI0w0OKqO4VlJ0DdCjkGPt+DBLoxSBVUlCNUSvkq6b0RG4e4Rv6
jLMXC2U2cU3zKwwwsJ0EmucKT9yrVpVOn3i5XZVLo8qPLWayvLbnli1oJSNzNul+
dwuj/nLgMPWLjllkNbLtkTXeZowVm4svIsAJkCfp3Ev541ai25RzLw4f/n5fda5b
yEoacNLli01+tTIhXVShj19TxQuo1xBOtbC2Y3Zm1aLQmc4vBxhbkywISa6jyW4g
vndboCxBUMu5pT/7gRBpCLZPCsR1EB4OI2/hXXhFWvcyLdSdTt/7bJqn0B0wFUix
VoXC/PRLgDs1NVVLcVwKyDh/ZsqDXBax8YOjZgONsGjMXHAjcFrtxeF+9Rx2T+YY
B1WiA92zUYo64wy+dOOIrM1+lWR0AwwqO/pj530xhqnQMiNsNgywdQs3j/uW04M5
SzZW2IHEsUjIE6jWyaT3idCdM3uzUWInLirunZemOzAdeiVETrTpoy3jnAHA1q9t
WMu3HGT2Lgkmx9C0j5s6fIIdAK+S9HpyNVf7hXcoeZgwG0VvKcXjj/m1WhqGsmRk
aO36ae1PFstQS7CUg5C4f9151tXRq+v+INPaROcgLWv9QBevKDhHpGIofmOhRExW
r2uoZqk/bptue3BhoIN9T1WEtqOIShuvuzv0k/PXb3gf9iV9rDRZS6sAN7s/XLvt
8nrR4ODPgjuZLhjh04ChlMTB9E40mr6xOPKA0vTNJzGeTR4j1McKeTF29jN7RbUo
n0aJGSuybqo/HmObeagv25ywQUByoIJd/2IJYdKllzMTHvD6k3BVSHhCLcQY3laj
WxpJeMSaFpYHTvdo/4HB7zZBQ3zFodLyTyWspaI1CjIhQfJMsgmUzm6rqVo1zKM8
EJ1RaT1Deam+KEFXazxLUvDIrQcbc8y6mrJUF6qFM6ngoHmPXM+mYLxe/X0DrX7J
LGuD/1RIFJ/Bc5dfiwJYLSKg2Dcyf520mIoc6SAX8qkwja348eMBoVvvPaZtoUxr
GZBqHgEAJibHdGLFZtbBUG0P6YGrMmQ2HQIsWuRRHoFzcdcn7yG0L2OUKJIBdFvv
t0JDG1Ci97zmohnZgv4AmeaJsJQwikMUjociQDh3eEpsDNuRZ9SY5r9yk87Q/wKA
uwk/RWCMTlBoib+QZH7x9e+XhYMmraj1aoiwLI6CUlMT6CqZO/O9NQ6YTxcqLtum
/uZWkQCfG3Pqs8DrFNLxcATCkO8SHMRCMYux62URP0iAfyHAJWgRO90RU7n7/sMR
EVPjTraM++HY8vUVQ8g8qexrHb7v0AhheonemXO/z26AZReYnOazdp/iRbmXdm6e
R2JEfydBXQ2pG9+aRBmQwZTdCczEvI3VL+ow1JCFEYsCGgGveDwtMCYS5XlLEZq2
YW1BCcetVFE9Pu5SXHjXUnoOSrxYCIvQsPkwLR1RFyGx1CLH6mnGL5ZDb268dNqF
4mDspAkiFnbZm5jLjSNax6jRIaWKzqwrlEp6V6LVeTImmI3voLl+/jcmIxg9Iva8
PyB2mZ9WZ42T+l+ADtPTaee1wM0yK7A6u8PCQvX1xH+2mGIyvz7XeZ0uOTEMEH8D
fMlOMGSJYKOPKjkUh+3aQhXX7Tmew0xjFZg2xQ/kfMQcqurfmT/YT8zJ/l4UsuYy
htYBuFpadOj9yZ4ZWVXzRMVH9ORuHzDSVoQ2fGSWKrj5M5+rKDngGY4i/0F+q6YI
Dh2fvpag1MgeIdIdHufRF2pbtlHpz+OKNavg1WEQmqZuJ5v/UKtEpUBaiafwR1BW
YmPxic4M8Mh4iOAxqNFJoQuVHGNXkjT+xydTOWSHHCr6UpfWF+ZEEjdNcDr1xO2i
BIcWP9hbQBy4XGbQsmvWJTkQoslC8j1jEG3osq5k1jJay7QdF3Ff7DJqgXdqFyk1
lUbP/YTTJSGGhtNypaQtCD7bSz1mffHXkxESJhfZl1IrvUxJm6YZgCkBN03vhvS3
krPtgFgfFtUeTj0MmcelpwG+1IuF7V4G2mWx+lCPKHOPwiHd+ZAFMDOpCEe4NfrB
GiJrfb/mMUYLFVcuqwyTYwxQujwQoMGJqgaDwVxo7ZOKhYAlN2iMLKfO1o7C60zV
sGVRSE44F+grZK9ZrRuy89JVm/YGILXd72W09Hqio3DmFH9YTCZ1Q01G3RXMwjgX
kswkKcfSN7uFgd/oyk31AfZH8P64gJGJQxvzlNPgCiUTCI9tuqXSUG6dLOUTQve8
34MjIWHSeNQgW0VN+vLhj2PvFVhRjufa4IyRxcVtvR+62Y8ibAmc+v4w/Z0iRavF
BdG6HeGOBKV2M4Y++OlEcI6kOXSZqUuFrdEDMTizAVLW2LRvJBsN+dHmjwCacoV3
9UbEtAb08BkAE4i0hV11pemkLOY4bQwpCeRP/0RqMST2glrjZMUECRZE0OcICjLL
zl2dvUr1NiYbjJOu5LqgcvZIXgKe6S/gtluPUkMsjJahRbn7HvyCLJ7db8HLt8bn
Q8BS/eRhOPlweLKjgJS/HzlUAQy005HvOdiojOQGAKzsBg6pT1gKscGCH63/Mmyx
OdsZ6d3ypXH/Nn1EzAHOpZQ6xuPUcfsymJbcW9S1IdptFEjluoN7U3tlCgSvQg6H
NEerp7C+Ztyohd27ENXwTyZzxENt5PB9e3+qhBLZydL93t2EaH60Nva3uwtptL4A
G5i2EcL15GS/tybONelyN4B/TasApjVCciWe/ABiE7ROtXFcLMMaGmSi0MBvM7NI
6fqRLnLClqtv6HbHYn0L3apZobJam25k3MS/pyGFQjRW4PZV8gFMla4AIAbVqKx9
p96JPS5GJr2K1MsTo2stJ4QPBLW3BX6363GJMTwfh7zxQNgSxSChKWQ5Nm0Bb/YR
8JL+PCCs/yqXni6W7qY1ch5svmOoQ3e8CRCheb+s0rA9hfOqa9bhorgsieflTFwL
48DpGxHRj1zw1Pbme88ER9di8A1+bPGBT8HnTnneZsiwRzR3gVcPllyKToB8yFGI
GBI6g9deoR49CCFk2zHQCnBT6M9faDGR2q4GS3WAmexJktUbS0LefsnCrr+RVLAM
ViRf5t3N2D2USonjnyI3nHgurmQFFLMqfHJOcP9uSN+H5tFPGNZ/BYJmlf9c6h2R
7YYgsfKFPzQrxEv2yeKWXGMhoWJO1paOPH4tyhYIIszw4eWQGGp0LMiXvgR/87Fy
O1mH5/QboWRWX7TV3yHC+7vOY5txlHjaGw7E5Wl4lJ2/pj8oL/N+vV19g8FyIojK
lasRRv7P2UFBstalPYmvzZyh5pGUwsvt2w/yMoITirfPzKEtDO9+Zu2uT0c62ie5
3qLlZRqOmTHLwMBaZezPGqDrmh9Xo14yShs6wia41MUfK4q8K6NN6EwUkueO/6mS
9kmFd6kgxexXETVAxolWt5ZEBzFswxzIguP+PJHPwrS8Vn0J9N0otTXG/LRZYJpp
XAVv2kPHufyEKx+H7FuiLNZg+zj417RYBIwLps9+i0YkrWHAT50MkTbOQkPo0eZc
SXokgWDCrwqv9oxR/zzwrHnjqCEkaaVNvGr5xvKqAratNRaB24JJBSi23qIV76Mu
2y2lJZLSQ85URFs0jHeiE1j6QeZtsFC+leIejui0SwliK/5MKIggP97kIQEv0yaB
rPFLcYITGT0c0zWboMNxDXEFFCwP0Qp93XeEtSL2OtjbrNcVqqLiiNMiRc6fCZ8X
nRJCh6s9ZSZrpq15O447nfRNFTUHIBjbfIs/NkEWS40ODCAhZn6Xek5p2fHQNnFq
Irx6oJXuLEmOWTSsbHYSWCow+5JE4FkQje+nVANMYazAC8Deol5t6EvYl9XTfCf7
dELG4d1TYZKyZ6AOKOXQTTIUaMGHeB8By7NkflvBTQ6mgsoJk428tJlYeUT91CfU
gejSwQinnN2ifUTlvmleT8j/C3bAGlJX2MlBtEXrdEH8aKOrc6j+G/4oGv3y+4JM
130PMVtEeR4CGRkK385Oi/6F5BIg8IgQGxXrSWijHXm1AF9Q43OnriDW/EBazb2q
mg9wmQmmiq74YYxmXVe5depuHO/3pnez9DByB9b0m5E8QopLLBFQed98EhEETR5m
W0jdeYCVVNnl1VyMVDldGXePS1UkcKC/64qU6uh+wlXfo6+g39OApBWXL52eg28w
zUMXtQW1e/2Pi9gX1yQalNKwiIJ2XN/mSg9l3OBRhhsoTlMGuHECYL+fvOPpP+Fm
NY+BBN/YHCco793jv4JBOW/2DEp/2g8/MiD/2zY2jFsU4PMf9q93If1UVwfvonjW
jvCq2iMwE0kH+h/Lh783JvRGv+k6c9sRS6V/IJEA3/iSjJW8t7JtswUgFWBzSoTA
m0Kmd7d0ZaIaSEuMSLIQ/lJPL7fpiLKsMlkYDwaFghrx1tPaTU8E1V/eWlWCK3vh
PxGX4ZFBWmsGT+baFaRACfq4mTsdVjfPq04atr59K2ptwkeey5t44T9M3BbiWVOL
ljnz+7W0CvsiNMkPpDn4qQXO1awPxflN32YSXt9x8UYQt9pbxtphZr2H8ZFUvjJJ
mL8uANRIB0RDqp/k7MyHsP6acfl1DDyCFBBLaD1lFxPYwdKFguZiTpEog0LorojB
q246lryq6zD7ezKAnsiEaGNQ16c2Tau/ojDLlOe1i0QSdVcrjqpJb7PW07eGU5y1
OWW2yYmz2QDaUzUpKXcLfd97mR+AT+FYrbKtpQofxbXmIzD48ApZ1SwtIBT8ZMZn
bCbtir5FTeGJPQcZcfZsuUChB3tgVrJTNLuP9eYEI2UvVGWb/63THgC/Gft0VoO7
oQXp9cnZ6039FwJi0Sm6PmQMOdncAzL4geyyaWZBVQxT1KyRaV9IAhWXTqdL4/c7
X9HHkeHUAzyFy017uHzsFGyalHvD0WxOePCP4s5ZvKYiy+4SnGVTKjt7UvHzvjVn
UMFIyePdKyJaql0MXlj8qogIk3zhvPJ9H6nRzM39x3DTPEwtq03cu1HGaHjwglp0
/+8w0ybY0kBagVLdZqv1ev2TxKofybtQ/Mr+JxqajnJRce15dXrd6rc9wa34kOKn
pfO5WtDZX0+334KfZoKwnmZFoTblfb/GlL/NOoTdEjOoAG049t4LLgLoBjOsjWg9
s+lbn22HqS5QblTZgJoZVoSbRkWbb0SfTotUHmhvY4rF7NhP0uh8TyBkfdgudgo6
QzAcd+yE89Euo4sVG5HHu/cEnPN9xFmbf2jfYjG8jHRDMJcYZQn5AzcljmlnUq5j
aRKrz5Yw+L/rLptcCHeBo9pMuaarLiYohEwIX0XxkoaNsw2TlZs080mvFyOwFnsV
aLiCTWSlQJsqutZKpZi4hrkPfuCe3l5Whz/cn2yffsRrKzdaEHzcSVD6IeKwIZ3+
V9HFRjL7WB2qISNH4bmJxWkVuCahzuO7bsfkKGxF6ckk5A4KDada9THSXe0zribb
2Pbs3Ge3VJD2BavoHnicEMfFuPhpd7OWFJD8M6Ob7+t6XNGJ03FDnKLjoqFt3GJE
lWpFkCTNrdvg+8UTI01A5vgeiSeiZnv0uXMCNU1fSff747WY0UdSAKHamDMDnGsr
W2b0PPuxqHGsWo/Xz+5jVgmZGkW94+p4tj4Lujvl5m+rS3L+dRM5G5U2HwX0JrSz
AGA1uM+z03qI1QHaMsC3Z5C/92llEZ65WZPqkHskMuHNpic3L3m6C3cmE9fhFHvm
5Es0OaqwVaGMrlN3GrdVxhMNxDh+or/wlAP8WO1wKAPsnEWCa8+Q+CBXjZ3KqROw
1UmoqWVijGg9YuVCU1n0YIoTpydERPN97ULJQG37P7XDkZqmcyNEVlJzRYpJR8LB
jNMnrKc+I38Nzs7ndAp/zHveoU+GcLuc5IfVlf6+NVEyqGiV2pxheSYZqGl0hWlS
0cQuvbsdRPpCMscE2ftO7vTrLk3WRCnR1KTNYUjc7qoVVR73CV76lV4FZU8OZy1M
++gIW/184xlAlDHjVGt3Xdk/44vJ3Kcml9CWGl4EKL9gkh0+YkYvoU6LPWWWDKZP
Xf9tCVtM9v8uWvuv0gaZq0BuP+v/6AFpfONtZQxjLHyHqq09psVGvj+ejgN926ni
c3s0M1T5W741OD5iz4AI0PZFQWUZ4AwuWXjcss943juXNfBGxoIP9PwopbbyKK/x
2gsLAyZVo7vniKVZo3Uw9cu9Vz6yk+TaW57Msf2ouAQEzokTYOFsdoRPZVNhWC0u
h13FHqmZJUhCFbWK4PrxKmH1//aLbJatjfzjO1U+KezJaRqOUMUV40TxrXytdiUJ
f+pBjRe9TlFbMqhwed1Pz9P0Fq0ig668YGMvEAo+mMoxdUapP0u8g5g+ak/gcSkS
h/DXS/Toj5rPcyBr1VTxnl5PfF4T4f/QFz/BGqvEyCECemZAP8ko9QrYGYlHAdm0
FQXEJqM+KISbvECWAVdGXg5XjT9glvmwTKWUNCnMz2f5TRULt5LC4Dq4Hdk+SDBM
+cLwfByDD9qE5x9CyW67MfW8ar9iq4Q8boIpULDHoUC+JgtKdMmxcEbrPegftNFb
CZxe4jWNsZva7quFyhgbbih7wjYu4AjcM+PBxIPx2RmR72Q5H7/XDOKSNr1ThV2v
tZFxMCuHLv5d8B3tB/kds46QOdGGnEpb/93kX4N/GOY5X3PKT56xU8iIJzJ9rHoN
rPmG4Zlyt5qeVdPqQ3zcckWoD5J8jcvjHUQwPAM7akZkiE0HphxBrbAlg8YKLeLs
2x85nAvEwinbbDzFYJNQ6Dq16Kz8+i39KgbUnjV9atnEx0cFgcCKiUeuvViazwPO
8VSYAGPLXVsI9fwiy9NcdX0gPJGIIW4WcTpY3hhouq0/GJYlJTAMh/cOPSAHuK2a
aEOMed5UD+c2I46WZnTQMk446mnzPdEmCPjqx2LnVbgSchzgYL0CrkpUo6KUKs87
++RtzMIfDuPIjSNHesawKRTEASbbBDtv6Xiy0WlcK4h6kVCmrJcQcSmprbZNZKGI
i6h2QXhdF1988F3wEQHXSfN9gfvdKRgDHsRTmUEITNwMOPATG0IwcyolRQgXlWiH
8GOQZS8LV/+oUYG4Od5KEvsH0b5FobFFgO/t0NTbuy2SOaj0Ior76SvUo0meM6Db
NuTvcUM3qm/gV+YNwa7nx7HLpxxB2nFeiaEwL0+WYBsCC4p3S431hocXHQ/zgLcl
Z9zbacMN0jxebkTdA5sqgjCW+QKBxoWDUP23SdwDHQq/g6r6jLMx9drcQPcD02xa
sRCwXD999ZiBvvUreFLUFRDgRbVpR4QmmIW/T0VRN0W6dJJslkRfxmk882J0Buu1
ccU9nVAqBGYPdvNp4EpLh7GfgiXQ1kHbd9CnRFgXqzkA0pfDnMFiyzaUHdZYOLmD
haSGe1ViSkokMyPQNyeVi+n2SIvtTZi82KHMq5j8VQQmC36jCNgysG+wQwngEbqT
5PF0LQqupgbJzk/+IOxzYx7YVlapd2VLpg/Vk0vBh85vXfJdemcox4DHfJx50reF
ZPvXTNOceV35rhuDZI66nSE45k1Ke4yqs3d3qRONEFiINzj1U77vxQERE1e3TeMx
Pq8j9yosqzn8dO/JJ8FdMU3XHfh1rG+6KRQYtPAaIKpCLCXLjysqyf2f6V2aYpsF
+XxKYkArDF44KXtBI7QDFp0SrB4zob7Nhtfjo3raU22pw2WL7BvZ7SkVuiH//jvI
dsWO/1H0u9ygJsHqG6yZ5cj1BGfhiC6oEJeZxTIJk5XD4WVB0fQ6Wf4t01mMKndr
bH5ytSDiVp7GBKdj+0WeNQYWsIyBiJniwBlsyXvT00iCGz5GDzj+hv9Z+pwywow6
Z9pjXtmGVb4U5WfjT3HIm+6hzagSs490kTiA0dkHZJK//CA50gbvxU12DwwGde82
01t+SQ0HlaaA+5lvhCftCOVqd05rUx6ayOj5oojJ5IYkjOozZ92m9nsoegVSKWHu
9d4uKHRBTmxUrmi/h5yg3BV8ETsnN0q0tiOh4ZEihx6mvh6HvSujMyXHXu/J6dD9
gy1nj+/8A+8uutZEXKV4AUOx9B2YmAknbfa3g2IC64lz2WSKowjbr8SSvIBN5y6H
Qp3TbER5dz0WxYxyFmYXX9P/Ip/u5vyGfqiZc+fMGiNDog12Cm6lQcE0IVxwRfeh
QQT5S083WJ3Iyycv/enmHRWeKovoLrCuOsMhOvgn/NaOIH8G+KEQFEjBKiYXc0BR
6KXQp9f0UulzcwcOh51yBc5c1Jvfh2yCSFj12o0fn+Zlh/PlTC9xq8FnU+goyuuj
q4zzfB43Jo4l6yamHTxtfF1pN6DCpKbU1RgZ3HsEmLSW+mT9nU8XT+eq9CnzMYxG
HLRisPF2bioCJnGe8T3jej6FXQM6Wo8o9oe3RHAJUaMPid9+NTkkOdVj4wJkc7KO
x31p0CaxjM4GnUieHuhrz7bMLJvjpO2B+XOICsNq2dnN200zLT6gZqsY1qqPtRKr
xmZhHOVTbWWKKG5l5qawc3iW4QFZuSk/ydM/x564czSlvnlxz4tssDqS1YeE3QdB
Jz1GXjwPWBG6RXqWuIKXTmhkLVZ9GUHH3bVqV0sCwDGzrhwsJQ9UuLGEzKH9Ib3s
hHaqR0GKxqkGSdoQT6pdB5/5NaoPmFajmHABNBSBaajOXL+HBvTnNXWmNEYlkvLx
R45o9cNErj66P40cNDpMZ68sHUqAcROSb5NPuzWj5F3EYcx6218LommcDuyPfCMq
zas0u2Pf1AB2LjiHTrW4dLCj8BpZjVtwvsIgqkgt/03uZ10FsJCf552JdWQSdqe9
8/WH7rOz7kiiM7VLKfOgaT1pLJqGeuGho94eq+lOSYWYXakBtXFQyZNG8F8JZYEh
TyhJ+dhLEtwV0Q9hhK1DzPvQV0L2F9iPNhgW7wXzyCJ/2aLTVXs+UDmMZRNpRAak
xVgxuLsKgX6t74IbFnvAEYSXlamgPr9Irop2tX2OeSFAisc3O4oY7pGAESA7wtUE
e+BPcZcZIj3BqPXqVioaS4/+P3TlwFWQg48KKF0mNHbO1zv/8z14Zn2xSFRzDESj
klHFw2dk49Vj5LeC8ZyqKPe6E0SP6zf3W87ybUia9bme3UFW1m7HKqMLaMRj3Clv
JEc/SdR4Cz3b/cpOayfGd5IQPQxrE6CB8+AJWn9EpWPj72YlpN076PGFKalECe/e
7vRavkxmkA6eesh0oGrKxsLu1Hr9OqrQRUcmlZioXfMWb5zpQjDZmT5CaI5Idh9x
4W+JA3aTq/qp0iIngwhlKXiiBvTehEfLG59yFCidVOPFJNJE4OssiThVbaAbB/N7
jw4m0BeSHrQUD8a+0J4pwVc8XpolzL9niyC+ZLFi0+fpquwForms7G6//lj/QZG9
+o1ga7i+s+z90h5iMLsrQ3Y4fTSPex0FAfBwrf9so0ddCYCxl3a55sujn00b08F0
E4AqM9fxzo7F7Rfqhvqa8UIRvl/mNiRZbcl89yY67C3vZ/1gdgohBr3qmVMWGdzD
XV1D242qJP1ZehQlaWykDhuR2YhNJwVsgf0O+0lBlaK3LWwqXDipJX/LjgyNFWfa
Wj9PPEfLK4WsafEABF0D9s1neCvddO+DRN6KvqEYxNfm09l1YeiIiYHG/efBcxK1
5T/Sb/6SlQV/X7D7M0yxO3b8dDsH+xC0aK4mxJ+2NelXzrM1aw3ipuQgKWkh8AfT
covUbGva6I3zNCSeUjz7FpggSWuKYA295gXhNDqUxMtd9jMd5V6G0ZHRvGJ4U2nZ
TrCPOXZHtLtiAWjKgIz9FJSLNow8k9RnQlZ569XVHMmKXpoH3/ZCxllwAmsYKNd8
Rem5IGxLIHOWhCge9TRv2Zb+qvDqMT2RkHICLcxPMHK7B6l7rmYntqxv1l5xWRzb
nXwMGqACUeUx2vpx0wct2P9IZfASCUYjlgIOO7/SqeUhRqwpIBx/pV4OQKJR0hsy
416n8pWu7VvPRUw5fpqXj2DmYkETShv5yAnWAW4feIUKrUSyDhJfM+LQgfF1vVZ/
fQ/k88cARYEFy0EzGeT1G5vA557uIjMRnE5BHxxVoXGxmwPiucl/86y8cfkfXl2j
FKs9WvKDWiWViueBjsNLngkGQR+RjBWXgzDq6GgWleBf5RnXnp4pNZ1WJESsZyRN
jDcVVd714PV3gcOUB9gNHjZMygvRxmj9e7wm/tP3dtkMHPVb7+sb0MKDAwcavW8k
VHt2e9OC7udQGQbJKABeuUX820fxDoOw1Z+UFdp+Psiodtk2gFBheM1E9Qnj9MPQ
zO4qB2Z2xB3XslY0qAYy1iH6Y9w7lSOqN/EcruBSn3QJYikRfGM5+O2kX+ZAszvD
3TS801InltkllEMgmt7n0kO1QEvu3QqElAYwhghvCJGuA549G1Y6hDpBKmj1bKOU
kn6cztRxHkJlai887yK77tGT8A+5b/d+X+0UVjFneZS9ymyRJ9I4Oe3zhnHjL0lA
x/quF/34h2BaDml6ye2+5O+qmNUETujTgWTXg4JYQUvdRx23xxXKDxbb16WygHdm
bG+aVL3MMN4NSqa8lRg9pBqoujkiIeGKdniriZBA1aq3jWxIbMzFupQNS8DsAI22
kZV7u3r9U8p1nSWh7W8CCv3uzi6FL0IXQHJd7s/JR96c6e3fLYJdcDpG8uJZ/coG
KjLUAgsmCXVv2W6V24Yxy3yKzrdc1/F0uwjsxaeAgvzFP7C2NauJ/4De88iEG6vs
/S6aaJEvLljZsCkQnHiT6i8NFvlEQ7DNv/TP0+KzOUlRyvpxeJPV5+KEULCGvmC5
uJpNIu3XPk1WalnzWnoj0oo5LRE6bTC+mqCZ6mbVicaAXsMCfg/ulPncKFKeFsdj
hQW2KIItAJ/4B3Hm+v+z36uyE6psI4WFz1WpHJ1jSfVmeC1jcVs9ZRLLbe9z0DRj
iARQhzoQ5MCccryFGheV1nOxMO01QuZlB99VStHHMtDBdREGkr5H7GAjje66u0bk
oYGFcx0whnZJjAdLdrAgjqaAA8g+wwJdvYKC9jCADl5fvNcbtAiifMR6ziV22W5h
yHCV8/B9PCEheN4ahVL/bJaM93EC5x3+RLmNBpp8cpect0wz3VM4iB75mXzOHwu7
jxu9530mgVgdNCN2Ai+syGo4dPGefnDRrABOW4MtNpCxAet820ao5eQcosbyHgcX
SRg0fUjpFBOUVFeRta5sZzKGPziSNk98U5f/t0RTUKqHvmmsHAg76F5V/fWn/1g7
vI5xOYZSvmc3ZynjtHGKAV4vK8WEpVvg+ZJBfJ8qB0Z5GePRa116qHIfJe72/QN3
zj6E4uKTCtzBOGy7fAveyxADArnxk+nFS34OiGcbThADj17Pr38s9fFovYRa/vJM
k5+lr8ucksy4K+74+PR4sDcstzhEUOC+toKfT9EC+eBHKw//vuoRznLHEv2Ughxl
SJZonUZu7vMX2mqvKeKIYekSVqoHmBxmMFP78FRfcl5070hi/YtZyhY90023AyXG
NvPac0u1jxUeAudH/2m4ZsTqNLw+r3sWvdROdRTp0Grf85JEjGTj75XiCL7QAB3s
8Ez3I+DOy/zYQhxz4npuKPUlDrzLSRM6tvY9RkkYfri7aFisskQG1LPqZkxdBopH
EmDElULFecE1yQQusaQ19yqamShHHulM8D4f1XSatzgN2o9PYYETaAZwIGuBetIE
rAEhUalIVu0kpVkDP9+cFPUkAN13WeL+dA8D0xsRtWm2qJLXq2NTCvd6czSwUgF2
95x+5YBiR7o4Q9buvmcD5lFCdjfiZXJCOzZn77C0xXVmQShVWpKzt+ukkYaWxDQd
YFVHBpjKfNPE1Ckxc1DrQawM0qZ2YJxzpP5N8FjF5AsganQ2vrL+py/T7E4xTje7
0JfisTbV4GK+XdI8E4yb40+3cvYSQmNnHcaTDt9cQuDZuY9+FjwYERZ2rdnyZTgG
bgC1gpC1GOycM7fCTtA4M4oZFQ1/lmWgtWO7Xt+LO9NfPQvkMiTIO638oi4Hq/Cd
mBi0mbc8mccExAbP7yfQxHp4ibUyRVkvEg+YkQ5S17H98hxoKPY7lO40ffU92Uiw
HHgTAorBUMF9/9UeUXoNUk9p3JJ3PgUw/G1SB+GDdAROeNWmynLtw+t6gxMUaf8p
oeLS9lDTjdU41BCrzV8rNHVtaZo8wSD9E1RejUmvHGYdbAQbJg2Cz7ucxT+p/KOm
shshTRagKoSCb9rwoEDqFnARhpN4CN8jy0TU7SCA75aHMZbBjo6ZBr/1ANviyuCm
ru0K7zWrKWgBqW1VP2lbNmPHtTolcfycHP8lnBtNhLIoTZMwQVH6Q6uyEEpKPJ0S
7NPBIecuArSq1i02rIfvVW7b6q3Dht0jJdBi7xIdUES/LaBQbU9tqr9Z3+Vc12Pq
n7XVxhEG4XxasuCUhjoqaWJMefeJZm1pgfabZE3wW5apBoc2WRaaQ8NboNUetnO4
cWgcVqkOzi6DawLfR+X+u/xoLTt4M2aKPV1oY4xwIBD/jek+2e8hV4TVLszCNUjE
XFiRySF1G/h/5UYs3bMpDRq08ldUs6hrGFm+zMSU7fUKlnQEoXdJFcq7JRDUSH89
5/uImV8irL09t1wJRa9Q9eLJ0DrohvRYx01B56QVrJd9SPNYNgymLDEtTJjCpnqc
YEoLm3xxiIvSh2UxFz7m2Dqfgsf2kOmiFTgC8yEWharKKpKC4cUnXCh8kqObwYls
qSemPelL57y/JTmEjBH04n6eRBCZVie44EF8elWgfuw8o7GKVSBTHPv65kxUN1ME
B8qH1w29OT7zzyh4MS9vZLKzW9DBJC87pxHpw1YcJllwLmc8xR72eyj5NFH+TYrv
kZ0KTc2xGDVfQ3qC33QvNKFArtLiGH2YEBj2qAycsShPDzS/otavDd+AXEL3K9HP
FvhMGEhEk4KQ3SItTDQKvPZWtFVKR4R2wJktX58hLAIjzF6M3juTn3cM0E3HL8Sa
TfCnpChQIL6bBG1jRbt8OZm0LKPC9SPokt85hMDCneMB3RGAR6mJnZYq+CIYrewo
vzmz3DIAqUrnFqomfDLyj+FdWWAJqQ7bfX4ATaggd2xzI1lkbZ8h2BWPhp3Buw8O
XM7uMI6dddJEcrB1mnIYDhlBoqh9eyNG3mLuPMk0P+Nqo3e0R3MePm2s8ytKOA/X
sfF7gEGe3I6D10x4rFYg8VP/jXGbrT5eO8fv2he4NB8V/QaMpDfqVNRIow8Leuaq
O9TKIwnwbCK5G4NisAWWbGk0h2J90gKAHGJ4xbZCQFv9tzX25rG5Jbqxus7SIGvP
jCSc8EVYi3QSuyA1dQ9OU8q6C2nn2RIxJLhHQA4QEyECnpCkVv1KZcuQYAtRi8qF
mrTBJqhBVLjnlUENTkWr9kUE5HlAnk9KiKncjD1HsbZxL26Qx8VsOB4wL/smIkPk
x10at0T2lPnUWKfYBvhYrWYVzQn3UtVZbHo3LIjI/cEDGFO+lEnqOLCG1D/VgaA9
mkzkigvbBN4MwuT0cDFNakyFWOOggTrTsZQqzdHmsmQpZ3CBlu+6qhHqCvlGAp9r
BfNAb1Hge1uC/80CYlsIY+BZYKRskEmK7IXfQKlGEFuf+RQfb0YyJvqBMfsqT0xh
KuI+xDwppIJdI2dFg5PZp2/PGRXCy/AnlimdLEDfRP7i+vS2ySucxS+3byFH/6+D
QUjM0FnS+4faHc3SKyZsZQclKGnOJTSs/Z9QvOEtHC7FJL1+TpB+JQ6M9U+OQTW4
cdtV983cT2ko4RnwTaittFCyEe56rTlhCy0kPlL5ZuLZezxfa82CLzHVcaw1hJZD
Re3RS/4vHIlzh+pYLz3DBxLocb8gt8u4PC5RMBHaDYFUw0eoCTBAv4bu9nxeVSZn
Xe0K4OwNMK9vApyfywBGA8Mk74BizWam4A/J7HZMsnryJCw4zORvz7bCeXCWS2VN
gfCyrv7GVAqdWHCIZsFJgF1M6HO5sJxiFLbNibWQAbrhsjg3N70pC1DROi4OrGKJ
obhIwOAD6UIX2aaZmRzdvJtBptiQyDVVHH06smNeDdKw7409Sp1CIXzynlUC3wHL
+Z85QYACaKr68TSHEFJUKr9wdtwK8Vgo0qlNr+AUKp439o3+5Dakb7veX6FN3U2e
Zx740J7yafSDYha4iBmdIsLVHcGzuQeugJeew3B17S9srDZG9GwLNss6dZi54620
UdQvCPfjLkr3jBlWE1FXJTBPKlv4dRY+luBY93m5VloUS1COF7OAX7KUNeEC+VLi
31WE+OgTuQbXi2Yh2ashMyZTrNRhu2gKw8gjL2gW2GKl3ifwFNNcbVa9iCbT6qIN
V7Y93wG29AJTwKj1Gvh9U26pAeLUC/eB1hKtBm/tVMsIEREDriFKEFi7d7dXdahF
Qk7CpSsofxBxHnlioLLIDTQv7x82lNtIZc+D4pwLfgB2ahhaJ7VB81BZa2k9DI9i
+sK9LOfbOB+hBiTUfF659Ny5QOgEzZKtN7FRzskN9MOCOjZvWmvnvJxuIPhnGexu
wrk8i433l5DBBrO4XOl+PoKuLZI0vGDRxn4P2dwFg19Db/Ly3clsRdi2O16cYBiD
pICW4Kz5BiTIzi8RdEG6ogii3C4PnIBW9El9nmc8Gkif8gydbfEpS3K89FoSkLff
Vs8MX5S7nGe9ARYQGMjsvmKBtXRsd98Sd/GNcF/SCtJlP0B72lQZfZ724v/ErVv/
INnxRHMPo2AoMQgdGE+UlmyTMjCDI6JYUikw6Xjmvy3hHYE7m17h8ui13fRAhp8Q
281eQgqmVZJN4Tv1fdrPVR8qOnb0x8ZUZTmnMFn5cTs0EetiLNofqBSdvr+0dQIe
qfLGqBdcUS786ppEZwmV9FJI+2wx/A6VJ5alBoYfXJxbRoyo85z4eaTDucwvpjVU
g5tL+RuXoZD48IBcb1E2ImvBQqJBHDTbVZtgwpaMpH6uYMcG+GjgohTsKVHRmplS
3Ip/gzMvKKVaUtyFXLGB2lodxpKL+4/QvrZyHF1fDMGpcT0zy9KCjhmP/Y4phe+R
ujnJOidxlfZf4KMydkEyjTJ7Y6MYopKlaMToVRO7zwbRsDVGBpF9VsH7fEm7yLvS
n/wkbpA9LQaPyGdv924dLPgKyiw9xy+y2ApejCpiNPdnV2MoLhCOb6wY9JKt4AB1
AxHj9otiwTnkzemp7ppHScvPp+MLadhkGladPcASIQXRpwYzEjYDsroCqt4iJe0w
gcoIbR8NaYv0Gef01mjgcoMjFRAOo6J/UT+ANWMXYCAQ95ZCQZ1nc6C0AGZC1iJv
NV76u0ERKogjuQO4mt2KXP82G/ov7FSatp3w1j03BwJ0KotEmlDRWVsFeDDQNhF4
n25bc7Gz8jwJtVhyPm/hbJcsSxaSKaWNICCvPeAKcsrv8yGkk7ALPN+Albf4hi2Z
KIf4a/FxWDLhiOl4xsLleqvgajclsc2xFfw+lAAan0rDuE0kFpLjwsHzHs9eR+t8
JPeKhD18C4x3GNZJ5vpz8aGGURqW0BVnfOlxPNr5nTolDAPxWnTdlrjvVwm078vW
VqZ/utsznE69BpLUwl3a7N4slhFkNU4qeuCLjaIBO42yVy1HDoPw0LnPCzRqMEVI
xgPrTRpmUMrfJHk5w6ika0oWTd4rHsPAc6xrGw4R6xAC0aVY3fsCvS7epu6wuU3W
pdciSmx06uf2ciyqKw1X18MNP+29xAwyAVbz32Kx9NOfXezg5d0U7Uc0UnCISZaL
RGnPFG0L3pRSpIT8IKMwmD49fOm4mNZFUpFoP1vHFcr5hMnKcZJZD0xTL0hd5oNQ
geMviFMwNqCFIppNEs/t/Oy3mNBwycHF2uTwU0/PX+XsYu3/maW2/dEjQr0198xw
NlWSPj+NE0YDb0NYE/t5ENbIGw/1tVyAs1lLrA1R+ixtqGAl/bjfQ78tq1J5lgmJ
brms8Yl97PKJlD8tlP819j7S0DIg9U+8xpuKEvboR/jwTWEQVEhnLX/DFLsPTxxV
36ijHs8MyVzT8/ST5H5KOReUlDkdVC0Wz2o1yoNWfC2HFOj4jImLnLaFr8BaYGgn
EaC3ae3opgBvx/xPM8cUeISNJVYkgFgaHUAZA5fY6iG6wLADcyRZ59yqRTZ/SZvk
uc9jDk7h9vNN7AYmpFSuEJI/swaOSJK4EBr+W35VHQnUTUmaLSZciw35qNuE9wd7
/LjrjhGCPuElm2VdGEBThIquT0O2w+dYMKDbtDKA7zqdpTpzQGvdqsvesjkIo9qO
tko9T03tNx17/+DeZmQyuM3ohCeqruphBH5hmiQ1AfQ5hWeIyRggYBXhALdfPXn3
HXOnEljS7bFpjcUwDLY/uL+1C6Ccna/HnGxDGJaPvmmDBdpfHkwzdtYaWum4t1ZX
Aeld2zcM0YaaYNt5u9FmJBKVer9ZtAI74aOwg29HcA4INwjhaw24VNa4gd/J8Tth
G2u43uTsMaDoD8t+5SOI5kcT+yLK2MBfdG872ZTKFo0jqyknxU3FvLm9fgV5+d0X
dhgZfaPnkDAO51VQV+ISNnxjca6qKjsv7CufHSC+sOzyDZeiZVHBTmpa4mNB7Hky
Kgm5Cp3eEs7tKSnDoP7poGSpIMfMwYOxxNv0Fp+72vI0EQ5lEvg6rj1HSHTzIMBP
nHroXk24JpIbnWQmQ9tTC5fl1gLKjzyB50hyXGb2QWWv7iRRsCXfWaVcip3qQEAZ
/1MKdCevqmdmtsjDMyXZxkJgEDDqkW7FVJBahfnddkigpJ8Dw3CZLC7LCOvXo7Mj
7KQxaOrwNV0JTB0s8HMK5LF6FwWzqTeVYD+EXs9fIG8B7XYhEBWC63Qjlc8nfgn9
DbE74giNm6a+GUhsqY8r3NlyjtEdbKjrpf6DeEWFqSmCNyqAOZhsoFhYy6w/RkCg
E8mYolvmFo47ayQ0sWQqYfEuWk0RkcwNGQsTW2KEImywyf96oB+UvabIC/Bc4Y20
At7Z6XmGgtLXsAOSreryeOzU5CgVP/CHLaDKuVr8bmiHBJEg+wYWujK9AaPdeTCL
ICUDdEOImJkPZu/DK8AkxXAh2xfvJIEVyzlosK1ul6XNFisTpcI44SD2Ki/2lPk1
t/JXYNT0oEUjaYQr3KQEvy8MA4Ii+NP1drFWjPH3VJwJsCbJl9xB+hkb8V8b3Z4j
/utZOvpyo+jukzMk/1UNG+l7J+So0pSVviTARqpZ5dtfm2BzZLohyUiQpESZ9p+l
X6ADcdNOLGbg3DauroLKY2gl8u3Ffigwx3aFi1+JeKmhOXgMedoKLBJiJ69FuKZC
ay87UQPgDojdHPRkTmXOo82xOnA6PfUvBQhE6n76OLQPwlKMH/5uEmR3z8nSmtfO
ylj1CSTBJFjs2S6pb7Aq1WwNfXTnZ0RWcc/N/U8CLTCwTWt6bZKEa8xrT3M/BH3X
AQA8AgboR/n7zR/coz3P1gJrd2FYqmWc+r0q+gtk2KcKLc4IUv+Z0bb8pddk/Yux
q7APTB/W7+OGo+6RBNmztnv22RATvOE54WC8jgmkrmzf90vwUjUiN4uwqt93GqR4
edKlZ0P55zGXl2SSqezzoyo6069SFh9/ZlxN4kO2KlOIFVJcMxSvD99ayGjpJ7YH
MG8QQQVkAl1VnjfV91C3nbLyyr5X/VKYGI0wL0ixRMmprsua2RQEqKgKPaHpR4ug
sOrTiitzq0r1Rd6PozHtF7NgIMwXT+s+4qdVyfw0qyIIDRnQnAgE/HRRa5hi7+iv
eFMpgNem8wPCOXjPqp3PFZ0TPGkhF2JUGunfho07PYeEODDzsIAspRswsYGZbQEi
JbmrecW+XZcAHBYAfXytdtg4LBFKE3bQXb2DdO7LDHmPuoNWoV+WZTvNQCFJbVVv
pJIGt4vWnZOCxKqWWLJ1Gw7cI9fB9Y1+njfROa8uLVZBLd1YCr/Rvsmm9o7TWyAB
+27F6y1H2KsqlO9LdJYheq0xAEPH8O5LfmhyxGm5TuSQFd6SQy/GCn2wmIyHSOQF
PegIt7/U4IOwIEIa8j/p2ds6vLP8BxnYOG2OuptU7SVChHkOUS8KED0oB41MEnaU
CVThYxE/QAv0oECEuG14eTNBjIE1pYFOjeRS7oaBFcMwoklgRiz2fyfYaieD7m31
V8t5ppfAyb+oFeADfR6imEbv9/ggGZMBZ9PaY4qv/9mgHfQFNDgP+tu2b07AeDzI
LY9FpxSF4u7YrxI09JLFS0BpCKkFpEuiZYj7ygzQtVK6sJMZgmzlMMWjvSJKHHmr
QDCVPDzf02yR+AUslq4OSiwfIaLmwudOed7CpEsN01iPsRaGptXlptoXMKUejWm/
ZKFEvpj47vB0VqdoBTX2fNH8eiQcP9dKwjxmqPtXJ7hs5SpmqOtSzgDYKNibkoRT
ETXIPf446FlLNNfM895Ry1OqQx4VLQ/ehrgzV0AtxXfNiRZpjrhSZKHJkccUdq/k
h9W5hQBYk3CJ0RcZ9CMv908NfAMbLee/x8dnziPJV61s7qgmfJ1KviQUHDPRmuGR
/YG6JH69/dYKvtW3bpPFBdBgyGJNAwRvg+V5nb7gC3/hF1jMcy90HJwyZmPcz/hT
JhxqupdfFizlMrPl72Bz0lQF2O3yS45O0OhWxdkRmcgZODd1sK+NoIac0FmBCQbh
y6JzQzLPisVeUcgUztw6ZIpc05JDxOfQtLgR4KAP+KC18TyblE0ZQVMzmNPMRw2U
DSZwEgjrLGcrGEqK4StZ6ZSkBz7D/Zb82rJbbAvs5/xPrPGZMPEmXqAgPAf3jxOa
usDfdbsvyHBQiNmwS8qDPSVcfNF5Y/LPt3NWSB6JMuPPj/UEWNkiuStkjoiUB0Lv
WcarnYNTdT7S2jf6Q0xC+5YKl+8nFQRYtGJ5d/eXAa6S6goCkcS5/PyqFrM7zIlP
jDgYTYM6ykDytr4SJtsLfk35DKKh392U9VtK0QGBMezQ0H/hJhfRn7/6Rl8DiKIv
rCN7oxDsCs48l2hXyzSfsubDWPDuzE/U24Z5e4RohxeEMNhi5hJ69IayTwXmGDIm
LYeyuPAtx2kHIOVLXzzMOtJZFfj+dWisOIsb8Ojd4gQaKkC+oC/NVpaRZv/Nf2cc
VupWYYTdRnZIL5/KcSOBMcrsotu9+NUkA7uAG/AF3ff550flaP1WPcQf2qxq5n/h
CRx7q8R4V/G3HmEUn+rfOa3t8na2ZRhJ2hFtXqbrH+uDHmxC+5YsM6YRQB8eni7T
shgWUrwAxAgPMYAjCO29/lfV8M3ux3LioF1sk8u+cYFQRGijhjGmg5wC4GM3leEM
nl41G/aCUj7uXSGyuPNeR/JNwcUtHWYgVGjt2N9kEX3jq0o6tFd1ejicH0FB5UF3
yW7Lk4URbjYixDhPdivTAa2ZHyJr3X1JZFrQOx4++QqivOynHcnXa6THRQcG0NBb
/xrIpqIb9IqPhxE7cOrQxCMSQjyUW2vaz2S41r3w0KreHv4ruI4XBVkpzcp8MyVc
vhc+qpunCUBVveP44IOJm1EOx7pumnoHsJ5p/Vl/8wH4kk8AU+7xchTh9vVd45F3
O43dSfsTvMmivUcXCA3Bi9ckDORxA8G1hkjB/o91kwxVTi0ITJL6atoExtMr4mQS
KAqqi6M2jwpWuwdNQz1to3e+KJ3ANVW6HNZuZ9nVXc9l11GIi7VNh/p/vXUTgZqr
LNTNJcwY3PwGv+zK3xKlXYy/5YBkd8Qg6o10K1SDFGrBZ6GDwqsXCTsFnp7dZ3z1
v2wSRuIoWTAkIS4YKSLM4fZ4GPytgSNXd8gBfPjfRY6LHRRs2/V2QFahVP7AAH0K
wiDB1qmEF8X/S8gEa9+eaWhNT/VsBY25GlvFrrQSEtXAKp2wATiWSDy5go4tgXWV
dGb3PtNQA1Ch2zci8YkVT7vfVWDdc6/Eu+H80yd7ULBQyYsg6Pc/FwsNm+ctiMEV
EkL/WzFqNfpqF7vhv69giZABu+KZ+HJiJlJUVJMUNDm7mwBGj9Sum+NQj9/B89tg
JDeqIBXXXWO4WApaDHpRiXKgws3biyVQngQIrmFk6imczAcUkACl5LxGTcaHyY1W
CVX7slRwf1hIFtj8ImQxe9w+c9bPSWK1/iHwycMPwZ7H/RaSAXhT0b0qBzLXyUqb
3frBt51th1f8mC4yFF3UVpHlGSnPwJ/JCmCkmSG+9rpDv1rmMNAdGJHncYTv96PU
LX4NE+nHEkVkH/SFCNZIiiRLzNdTXyig3aRZL7zqcZ0L1xgc7YBOT19JQoSTZgfN
hP9nLgOCUkqdcVEj9FsAL75sXZXCNq5ay7AofZ7n3GXXwfY1M9S3uV6TxCEoCngZ
muHeIQhNG3hX2hTfJFnv4cFrWIjJLmzwvuKcJG7A6hwwaJ/RArdL9vvScHIO6p+T
vULMxEge69m/5/wgOhJydZOcvD9YtABUxyFw6zt0f5sRPPD5mNY8q9Sx1QUQd5od
qHWOHH7X6OdkeK/zhbEcZrILS1/FV14d+EeVykyqbroZgJU8Tatj8yu/WLFShNRG
jxTCHyfOO0ThqQ90gAwUzlxPJoJq2KuFF8TDYAX0k28k8quqvQiwMvusei3y27Ek
Cq3k+LOfj/RrJLnrqZS07YE9SUlUTNJT8egB+WgWZaScyYR4aOYYLtNqLZmDyYL7
MRBPmfqU8HNimnH7QIcxmNLqb2cYyuyVe1e92UOIVsr1tw2u+vM17GERU8+lnoQj
n/+9vuWvxOEOEQrXrIuv1RmxXECl2EjPj1dCH/d6uMOPvnOEcWZ39vVEEdJK4Yxo
0Nl48uesR5JFmGtJSGJNWReiib8efmQA35iRaA8HcWLy6sX7etWWZUzgiu3jol2X
qI2cr/sPmfJXT9HxXmW4uYjaElNePNxwpc94DM9gS9hUMXGs4Ft/Q1gLvffXhb/w
4APDhPLvSRQfVxaAQ+z3R3Duh1H9dY2myCxLsXgm0oUBIzTvWpvQiDWNo9Wmco2K
MAyEfkY4Ik+q8MSXnf4apek4BB4wmQ2TBgHPfPDPShp2JEHjGIjpITfXfaNbdypf
Mt+vp448KwfHotitbuccugDJyFKQNg5CdE26w1EBluTooYOgulQ40J73OMkzyDs3
yLgnE0n++jKApFrrFiC8GLGwjL+m+lDzUujR4liqnXYS8oIdA9K5+KmD26GWtH+h
1WyBFPtwqMQLroZnX2nKvB3kkr90dFAQQ3ONfmNMHIW8bM0c0i52EqVMNKJrKbj4
iP0P7lRGu+BKIw22p8ZnrEM+jZl/SZyxEcjfzbfdNgYSr3SCU1zAyzwJQzncpkPm
HAPwc2rNHK0pYqzx6Fgl+yPTo9HAZaOqSxhlwooT2QPsuZhYIF4TrsnUduP5atmi
wq6CP9LzotcbQh0m94a2VhDXMvaRkrAwHbpaVj9yfifmgQ6g1ro3B7KSGc3dsWxw
dUxffxieti6RbVF+7eyxMSiENEmX6/IMGai6P0TTfTCo1BQZh8/xvxy0jH7r14dF
tyrnlrj+HWQ1AuO55HW0S5Pl9G3ZlksBZWhkh0nz35N+9gVDn1E+JNYGnPsUfOZE
+LcJ4/XoVcouEeDFZExu8EXRtEcpSLjlKP/DKjnAAVKaQu3keoc3DdD8OaFQdJ84
pAI+LgF4UA0akFjkGfih18RWQtPCHQDWVABM4pghuIL1M82QvBZAwf2XPPHN6aEC
IZwEsFku+4TfK+S74Hc1oyDXIMme/ziURDK4PrmsBWM4M1Cgc3zMqEI1ao4c/0yZ
DhxlkfWhENiZcmTYW5CG6BTaMR5beJ+Svh9aetpkYSjo5VA9R/bL2Op7lFwyk0Mh
j9QfX27hT/KbrPMNloOuC/qwNkBBmxt/+Cx5I+Gn76ga7b8eZq+vg02NNa7YfZq2
QMVYbOqikKfVQnfj9kFlxinAPzULHPeGnHoM+nj5F2jex2eDal69/HYEPQFU/hj9
Q78jD9WHbKViF15S1fdT82yszjESfK8zdNeU/r3zzwZ3Zb4E7b0hHVV8raMHzGUf
gIKk8Yc4xk39MteqKMW9xUrJGHNSULy9S3HF9XPOJoNryWpgTUZWYu/kbULdUGoi
WYndH8ImxsPDTzFW98SJQI9oPgRTZ4JeDV20w81vTFEBsFoRpiMel9RuybIzL+R7
vFZr3MnPJbmxgg+2qfCUwJIfot8/80atT5TR9ZwdsxGHpUSRiO7Bo8aQViTIi3cw
+5Y1+QBcI+6TSWmn47/+XzJwJicsRlz5XwiWnTZpqUvRX4dwMcb6YzZYd+j/BO7B
28cwOXBmbQx6crkP8IB8Xo4lQ2HpDeKQL3OxGQa+Kn770EHVii75DqyEVqfAfGzz
O4oLMJf9p17awyT4FZWlhJ7u5puXijpaFF8paJCV7+BwFAeIk1IFtygoL+jsPX23
/EMEzFrqyUIFHXQVDMwJGO3Ytk/CQnL2jzP2QCS58ihzDMxmupxiodgXLN+pb2tn
MeaP2L/jwT/pfT15SYlY64pQr2LsbO0kP5HUDFGecP0MvCwSbe33ccgLRSeo0wL8
cWqPL3zNYuIIkwJRm1MDcO6eWAoyQejZoq/1vdUIQyqBDSH9J5n8tt+eREC1l53m
/kMV8FPMekgYSFbFwjhkPkWbSXIiM9Icecxq3YLG8XrRzg3A7W8gReN4fFYm1Ofd
rkAsnG+WEnerEl2NUNUPplqQk3Ibmiu/DzR8Ulb24O6DYkjPCnbEt+8RAiB2JeZU
a70qDmSHBpvPDcvtFipvKmp2TqMd2Rg5rhAoLIMc+z4Rv57ToY/iyKf+BnbFbrhm
+3v84s/3fgNPApxBlDLMaNgxcpsrCIrCb5VaRaQ6qHa1jMlG9fvuPe4NuNUsXBom
sVA4LNrBsLZD/nEF7qoJ1Q5HXlS02ik3vpikhWB9ys7VyCSAX9p0Gkj2NTveg/ck
iP9Z3OTO3SScBbk7i+YiMHTXl71/B//rcxu2grtFdD45OG+sGs1f/oKUNHAmhOKE
xzXzazbUptDiAn7XkYC5Mce4H/svgNAjdOHcUaPvayL49AoT75tq+tDVQiNVavnQ
irl06Z46Ut3BLTsD2YR00E/iiU5KMJYSWHi/2MkyXfh5UR2IysP6D1XvJcjcopMs
aG+WqbOqJ+6HV6UzhwV4U9Ld9toKiV/uPwXkscbBumjtxv7hfCFB2wrpBku8yo5P
00KVPYuSWwhHH+2Dhbq7UAe/KHAGcazOb1VTXD616Q4Dcm/If3RyD7uAWIeZT+h2
lH6Y2LD1+oKX1fNpWYHGN19R1LlYuqBondqywFNykCJfzRdRA3lJ8Vp6qPIgpbIQ
NdaK17muM+8So2HIAzxDQ1XHFGMMsWalfg4WXSGzEclEClT37rb8kIAb6kLyhBRt
L2PzoZ+SfQe3WLFx5+x3sfrf6igLwyX314oWATzjGF4h7y3O/C0wEouSU06aMvtf
8Tip7AwESW3bABAQhGZNDSp+rTxLl6AgIjoiIhP9DCvJO6zknutu5JW7PyDE9Knn
QwPh33213SCCIDyIGcaK38edDUnem8XZkcxyOJoaSooYnGPP2uPzJchsdYfxraF3
nRDdZ7JBorqaMZyJj4k0s1DDPifTU0M1eiLBkNYWmJTbIiphmIsJb1j6THySZ1Nz
miLgicDF5mvrB/R0YtGeFBPVbGG5HgbTONAGJXaSQQQAvvmEaH5i2qGWV5EIARhp
iw6/IjEL+r+t/5TMbKpXp/5RDXoWvs4BEEo8UIDjU/JBCdwTPy0X7ASAdYudZKGO
G9wtSkDHXV5gz52O9nPMCSX/P19bgYd1gqtGrLh5YzY//1QAxPlrCxgOsk1AR6qd
dFK4SvZA25GZe1sJEw85bXOvNiHwekIIZWf8OJMlnIxQdSHk2/hPbpxM2B/O1PQ2
Whm2J7aZULaM2nm3uRBSM69kynkfK5fSQEfHYneFRFthmHU3oflUMahcqxL8CVs0
Ptvq2PfWg2dqf42TNhPLM5bdBM8tbnz9kesJrj0hdliJ5eBS7p1yLiuO17MizRoC
wlDKbVnA7pmEhWZWNonPOAoyaaTlduVUT57jrekpFXQyM0xUnNIGdJp/5GkXE7Sr
ukU/hhRMb7O7ZLlvMuoI61H9jW2ywFjcPlRdq0AuT1xlIdYj/uGomqgGji8NMDHN
GvijTEs3TVIdZTXQmJ9UVbEVRdmB29cnovPM/7r1RXe6Z9GngASXAQh4C27+LnrC
ONdYSfZjN7TlNPUlS8B0GC7jVDZhJAcdCOFcAc8uxtS1EPULAvx/WnySwNoGd5cr
YaHYZBokTJDO6oBI6eHkzsVaQNuOC72S7owxQ7NZpIzfpGbKbHZWNyKoA9oAsgj7
GTY0atGrE/1JOeDcAskT74ivJFMJXE6rHzQias9XtTNsIUnNleDhzMiXm8oj/Aun
uciWQIHDH1+Ddwe2pe26MGAULi3UuW6D759h46SZCjYW/o0B4pPkEI1tL3dw8LjU
qO33pXfm+Mw1KNePlr85lAzS6yirYrmXvcPUAO8ajw/dxoiV8Pn9lHWRKzUcZ3Ct
TPRkLCFHX9Wwy4w0xC+UE1bxPWLeAHY4Ucpt6u2J+LO5o58kjLGONSzgscIM5A+H
9Wzgug1V7T4XuiEQ8DGoc4osW5FIEl5SK5QdWXYGHeolyeh3fFqZsRpdC7pPw62Z
/aZixicrBLkbiy/mq0GBMHOtcpcuLtIo/dkCea3V4zXeUoQi5SJI6ozPhybJKUEB
0uoT98c7ATPy7lph22D6MhQUQx1ZJvUl5IshiSLwKf5nGKvlOrgcwCFEF43Ic4lH
MVu2cmwcrZumIwGw7BO9ak4iXEvJtexoPx7PFkXYfr22BgfCPkBPvPIv6ljS2yJm
kyj1wYD/o0d9wdU00k8hTOoSKYxdj6r+OaywVmwJIGGmHSdWqOse560HUh9FOofE
4Do87RyTJsl5rOh1IZDWn7ICowwJ9gnH73hvlkl+qweFE5JbYtZNeM8mGrrd6DJa
cQXhHdf05hu7pgMpr4Q4q9V5urkRL1tZdMQE1E2PC+eBf32x2jALeU5iLXxqC4is
ismfblVdg+miWBP+DhFdYlM1D/+5NMGTjM98tMQP0TINmqHLINxo/3A0VlhBCq+C
OJ1vz2SDP4DBGc91qUY4Q7ahml6hCfPMqqAMOePHq4fp0s5/KBQdPeeZikU/Jme9
GWXHBEV2AEYrK/WZCwR3iD7AwBcKtGU8td0TM4QNsLJkSw6EfiYaMF3vpof/JwY7
ZjRE6iIWdNmucS1tDF7vrVqEHsFw7CGhH5EzbeKuomB2IoljyH1xveYzkxod/6E6
iROkTFm2rMRlw+LSgAfY1VB/ayuEGRdDhyLnkd8lOElB0cwxkumZPRTKgMNbR5wO
AqUIt6Ru00UnD5e/cTWQpXPXxjjn7CVlbAnE3HttjXncXUztdqtzJTNLMj6vD4lT
awqI9OcrpR/rD0txvOV7JW3S6symajmuPdDMNzpbpGsMC16O0drNuKlIdvFcWawN
/oQxtFph3Nlcw4yP6rZZhE+Jmhl06txzTvhHtALOGqGTtpmmjPJxyosVzidUcKkz
wmewX4748vo4W8y9LFfNuW6tJd97jYvC9eyLi/184t8zz3gz9rSxbD2uJnqFP+7O
uLW+WHjvJiX8s4g/JbqoxUYdHBMqV6mlXjGHN5kJ7Mg6/xbafxZ2Fz4F59a5FecV
lNT/Nypyw5KCVnu4JaBwTH28Te6M4GwkejFLo5c4Gg+fZPHZnAb1yXKK9ZR5RhbL
z62KJuuaivITFi6kZXeMaprPzcnfFcJayahTHanFwUTpEmx2KeYIsao+GXKeCGHR
UK5bZ+nfuUCasY7DJ9gjtsaac8E7aJcgoO2oKCoYx6mCl+SaG4mrb1MJmlhdcmO2
sZxgaARZurkJMjlp4z9z5ZT2sJDFURiuyraHJ3Ah5ei54tGNSp+o55KftIJLegUb
qHHftY7l7NrQvlFBgXm0EQiOldxtMAA1/PRguHYouv9SuL2U72PyzXTuUgyxpVMH
zsHAQ93vbZWGFPC2g8Z/shPnps1dk2O61/xXwu70Tj2gKsYLDvWMeGOSqEDIYKi+
evrenylYKnOXTlMGvj0xxNIbfPH3GS+HdRHyP8UxJ5EJzCLQW8qTTOisVpyAnjzZ
NhPF9mKMhFNkU4txtKKXp2lIcufzbx6kDVrTppz+3edwC24Sy00op+sa4O0QzKH7
a9l96ySgb8gONDL0jh/4R5CDj/F1DubMbncKtoN3KJzriGZFKbzVmHB3It8fQX+g
G4KPIA5K5YGHXckXSZq4Safr/fPeiExXvCuzELbz/9hLIGhSS9EYFsVlH3HZuQ/w
Bi6BuyDwUYap7Anj5IP20Em0OiVMo1BwRRjW9WhZLNpdFSxLUixVagTwjBpjTxVX
3+iwJqLQhOzWqa8t/UqUNJ/9yC50eUGZF2mPrBE0pT7NYa2VuyF+tJSst6Kk5UuL
lt0r0Q69QQ9DOLTXiQpkzhbfhoUANRaY9zYYYKXiYkdEZonUFa7tEkrKQcdTHaQU
wUMtgJDEHthwR1iO6/3cKWQK7iaQNsfl9MO6BSyyVhCBkKEJHsg+qSWTXHSN5PWP
pm78bzTZQ07ypx8T3XTcGafZ1TFjoa26G3yFY7qRxtZ3iNJGAYKgnjMp2N7Zjcdn
iiQygE9hKzGt1DlCfxpdFiWF8kXauef+3o4+01juKzQdHk7zApT+/2iePRZlS0dY
K/MiIDinmsVsZs05r5B5YmTEIgrcZWjjKeuQHOavrFkilrbN+rsITEuX0owIDoWV
FwHAkcnd9AOhAC02KBe+Rq1J5UZPrpGpH48Zd+u+oZhLDKaVsfMJVbJbl4ktWz+h
bPXtEByUrozvOT1GgSMQRurvzBNIZ8XZ26LBXOJibjkJwQGApNyo9w+w7K8+M3vT
+1aMWumdgjuNEr589vDFJz8e87V5j/aJQFssWXElJYpAWtdZCloJAASldsr0l/Ht
iLJKFjs2stIRbq2WyWQAxcSjV0TRVy6KTtBiAKQ+/7lTn+wjEwignr3hnf0yyfuz
mOK1HQMeIroL23M4+Mpt/EISwGgJHTXGcdc2yDQRqx05i60wYfADaNU+1RSn//05
XOogQS92rcmqbe2XZC8SokxnEWrAfdgG5YLEl1tgg8dpWdtXqteKpdqV3TWzmZ8g
HAkh/lTTRxvjgM26ne0c04BIcqgqgQ9mc0sPm24KdeyQn9dRdwCy/qQeL3ThfBOb
tb6J+JeXrFDipAl+w0uagiWvVrdfWqb+dqFKhZJ/U200tHl7RzGkT8a5gdJmbQzW
E/bteOdHiL8pTX5Lhy2qRwl5TfT9v89D3uNBUfnHHZCh4wvCygBMyNHFtZiiF+z3
2x+SAxz7fD1vUGwMjRb4h7yxT5ciRjd8NZrauQRcmAecHGQ+0IFlZk1zUn12RMMi
28r8emlYkXutl1ivlcOLv0GOlc2uBp9Bvsl8nuuPjypcH6j+L8C4NMKs3Bun02I+
nKXFsswIHaQaTMNAiMli8gyh5jb0wAmbqKQ22c3G9dNLGF/tywePIDxNqAX14N3L
dsrU2HfzjXu9KqSId2sH/kvZ1OyM27hAOGoHxy5Kao5xDu3Cl5PESFWn8GcvE94/
CMA/2E9H3zpdgUOp+RqR5HG0eIvPBgmYSW8yi6hPTf7xHnRcp42ETPLCupdOLJsN
c38S0QKmzF+u0QTbUydNCNsVyZuwlfc/ViF62hG14JTwFb9zqebk0v6LhqpLdYXJ
IRkVqeeUBRUp5wzn2ZwXPPQYpLX/yQ+5u0rsVCar8udF5K3A7R12xkf+MuuqEYEp
nw4kFH0yzoHTUz5fL0JStwGQaE+P2TVafyURt0o8XSHwlH4iT+Wj8F3qM8iQle0c
aazdkEe3q0AAM7SIpNCwBsQgRCo4NYVuNHcz93XYZpGmQL2Nij9hxDWFeJLFkWox
z43auTqe4Rm8NiIKQ9YF/R5ZsEmD/G7+RduSw35knE0QRnBJkVi276lRY7H1PmYO
iNte7hvWnp69nnZwgZLqEsRjmosyfFJCQh9VRABD4I4hdmutoB8JmOfVxXMb30sh
ymdkjk1LySjFF7TyFq7UFfigw/HlD12yGmexg/G/8JL2prtZuNdLAv7ZWHiD9hlZ
Jl/8EQgUw6T3Q3q7tr9NQn2lIucC5QDhKy7nGeSsvk7e326azE33Wft+sW+EgecL
4R9n5x4uxbcVCKzfbtvGaErgyZctuqNKANrJaiB304xFl8+q/EeC5aCD9eanc9ef
QYYvCVBAhq88kBs/KNnxQs8lyecZq78D1GCbUf8ArUsHun/mZmqwNMjMQbZeG4xD
uZk1pTqUXB4j3vg7OfTkVBxNmFaPi6uAOEDUhLl6xNPtn3OHHDCd472zdQRoxvbe
c9Td254mYcgU+zjJAPzS0kZocAfi/6fr+TfYPWC9UuhffSGgEKUQjcxZlm5/6x9+
goBKzQPxUV7jpW7HAGnzHOvsiXOXstqsSNmspMxhKVwxYLhDWZx1AMJpT54XBtmb
0Eo8AtOYCZI2Zwr4+K6ptSvzjZn/ydVmi5dCbpUCWAiGjUJlKbMMSQoFSDspaRmo
ozVcwuwW+o7sUyrpt20tYG0MjTvi32d/EaALTR2HLR/h+4kkt0xDUakOuKcXTWP3
YTapB/29Ahq9POpix8iwDvLRN/9HKbWjBG6Ml0S0VreM4Ng3+XzuLUDZepHa7PAh
WFbS7SiG8G0g7/xb3T8UPOSMtuDx+jZr8ga68F8upDn3FhfaSEqS5+lDPOHgxiBj
18YBpQq22dSo1sFNwlYptGdoYjoUWFCYn5U9ErPMWLgu+BGd2OvoJXep6hMUImGK
JhF9lU1vbVyGJix4kZjt+Kk6edQLjX1SljHzy0EVlKXPW2c7vy6cuUHcaybqWgOy
uV1jl2XHqCtQydg5Y1L3wS6dTcYv/9yEQYZH6Wvv7lVyM4CqhTNYind+2wGycF1N
ZZ7QxQIUyS8nnIFV0mUKJIuryMC7vECB2+WLNUCWH4tzGZ9+7ucEVYFh4B/V051K
hMhSPVQstFuYOjtg+/8yWkusD7foL7srofmKypKmtNZ0cLRfYtiBH0JwUpWW6vlW
SMmevrINDD+4p8dLubvhFOTwCztRzAZ7EOV2kVsubTeOfWYMzytHQp1th54oyRCo
5dsPUVGR5I3+hzBmTwPG1xsf/ZpSwBhoDzUMJq/IDRvizBmbivbSx8V6LVNuvYc7
Wis7EzpyPhG4PvgyKnKCLHSGU1P2YN/h8GxKtzs7TLdJICu+s16D4Zt7Y7SurrkO
fb2g1nVcwweabUHd+/ySILrMQTRF6yqEsb6A8zNYpGGcBWmo/TnSxozQ2BDbWEcK
6pwBMTZwecxNqFc6Bc8MF2RLfwrJY2yfxApmXwnZCRhQM++Zpz4dsQ1gSYz6+6Se
GOFCaiVmeMotiVAGwVC2RDsBMT3MgGjJDKWfxKmgz9NeXeLHhRv4+doW7KxSDo6i
3+8VtPcgqHyE2LYDwp4B1GER5AUlPJ70IPpex0VYxjgfJaXS3ERuL3CtGSiaMl9z
sV47KKI6R3HoM23ca4inkEQQjYfhiwWvezBH6OGo6/NTiGdpzEIGgKC7cuT/9nI5
7p2fTHrW/x2W17dOgWfyMpZjUfbMYGO04lH/efsXcg3tyQem7C7VJ7lWQ2aqs10n
k0u2e0th+a9OC9zrSvgcbUVDiS5J0OHPQfL1LAn+0nftFZx/5wFZR8QCucOupJ82
1dsIP4AhsOUkmDFhMiKJumNss5+InHFOSJ3cSFOBDC1FmMv3IMDBCU9Mr4mWwlks
lLBVGD1GeCiro+Jg5259GgHz3OI3RIoiPrExm0SfhDcQGNd+2NemlOmG5216ceS/
rK2MCblPKSt3W+FVf+4AezUf4+9amc1kNQRelIJZCYRc3txYsNV4DcBtT5KtvwRS
Cny1UjVhqapBBqvrbgwH91zzObNSi1lzI4LMyjVYp5UHGzRStttU+lKWecF17zrz
ZkzTB9BGlJ74DUPVNu6aGu9uYqo6g0kkbqlehbPK8dz2nTDxP5OSNJKpiYvS+PbR
CoxCVfetbLnOqxpSUoaRQdBXB5qkPJt2c8Enz/d42uh1KcR0PQ92Z5rEAFAb64yF
hAQ0EKkwkVEq8miU4NgGunv1pZ2ooyPtf5/l/mO/+UEheEutQ4OOjHbUWvJmo/9A
r5J7OC/pwENlnY6iIqDyhZ7/oATDeaL2rx1E7cqmkW9zgyWFmcwLqwoNoGTpJdpI
pLGW0Xh7/5c16QeCqjsWxLSw53hoiTSJRezwq2+LLKJE7QlU2a1juAwKp81i0Zgv
KPsWCYK1c95iDv9WXJvkUkYtMqBLpLT0fCgkgnbPsGIzzHi5PDCQ4tkuMLE7IuNR
ZoG7Uu1XxSxflVM+76t/qvo04TXlps+QcO2Xmq/99A3tPHK/0vKrk2Stg6EmFMRP
Xi9L2FD6/CEciFC0NBQQ351FgXGQOjPvq2Urr0g8FJGGv7ldHLUQWjkPikSrAQ/z
FapCLbw50EHq/IlWSMTe/tOUxUS/43RC+JhSfjID2hwNdlho7uV9Fe5tf8F4FH4e
tYWjMcY34kZ7maWcKOaUvoVNr8MEqly9KC7W17GbZGh5K04EPDpgWYkEWPVTJucy
ybKJJ9qWWxljbNTeczvCqGGMhYDiTP5s9D/tJ5sqKH+4W9n6qrOKQJMzeHoHXOKC
tcxQHa5TbdC7lBLd071sZRTT1HHHXB47/wh5nzoCvwU+QxVha+TLRRrQvgRLlsaF
VHAoKIpigTFwjJvpgvbAlGafltdfMXtUTOuorjMpOZJi9X9pIoQpfjB7ep8aQUMS
qORrr53Oynj83GOmseKm8uulrzhUuXy7aHovBEt7EnkKi2C3ekP4mNM7pM8jY5oE
0GrDCJxb1CTzHQeF4I1B6ToiRqwDhULPupP7uiY/TWvmC+kTk+uO9YUevGAVt8+k
iLkZsWAh7JgYkwg5mX30CjbuBYx6SXKgeQq62WdR0ioMRQEih/gsafEmY3j2mkfy
lf0kwYKX4z+VUF1B77TZAWF9luunCYtoMIpmWzXvlm5gNPEG5UK8q6Kvd8PV/nBq
+QOfn6HKK6H9HtljYZvJtTcxTkjhD5ZSxLui5f9AyEUA2xOwe5f5Vm8/POd3D6yr
NtxDjWsD8kdPKpr7LOz82kqwqtAhNJc97pSHToVYK/tLS8gQ9gLOOSsbFi0/aB3d
PbL0fK+OjDthMgeWJPPjYjDT+0mVxuEv/c/dsGfJ86PGWrEDTKq4iYW/23RuSTdB
vkTLqq0KUQPAU6jVHtj4GH2FaWhxliE6Rcn5VjFbpkxBINpKsZx0DvFOJ1AT1h4G
UkPAfhGOc5+i5RHRXNHCrpOqCimiYiJOL53URt2R2o/pNKA1HzJLAq1RfK+WiwmZ
Ca8/mLn7ysKc7sAcvAwfrKqB0AvF0XPmqNv6Sv9wi095K3V0tuE/XLBqcdUqenYg
oRvN000l4a2Hy18UShryE+O6M07CV/mfXID1R5mJ8bqxzJsFtD5Idxn8cZw0/9Ba
nbLYebO346CBYRxFdLRui54NAo5HycrWly97VVfGl9LvQve+E9rN4gAxjwmgLMHR
xPJ59H6twwiJuoiTJ1BRRk/tnfSVQvPWYMr77i0Eml7qWFPbMa7WsBcE7T/64MIB
qWGYMsSOTJr0ddWObZwXDt/idJRm6cyYPy4gH0ACo1tnAsnEBCBf6stVbIlXthpI
4g9JCFKeJvHWxn9FjlMMGFknZOl4vDtWU/EDluIF4bq+Pf2wLxLWM3E4f5fd5po4
VjOk8Ky62inrcaIY5/COR9pkMTi7KMJUnHp4wKW4gj/woR0J3bcPxwM+qCAdz+uo
HboAyYF4mqlqYllyjhGoljCF/Rx5oW8TmacOLxWJMf/HTVDXd+atBqLCQ8kTqFLz
tXKzxkPGNl2g4M18WXoikb2ZdBipHAodOiySazJzWZ40jHUDcdjCYTt61qDPvreN
jdmpXhS1Bad6HTAMpSyp9Dns+vstoIixYeuBa33asqi7HPVKs3yhRYXBNDapq1z9
YqSevwxaAaTKmndFBzuK/2bCGy5UpDyA3in8luRjZntTvYaLJ5W8FR5EFnqLBust
3fTBEfmnmzQTLxqBziRw2Sq/pA8i8L5aZ8nw2Efyjl2RcDB6KOPZHO1hfqdTcMnE
ibeTJAtnHGYSknouaf5e63rAM9OskNi6bhJuuuzFH9nj9weOKs+ssTiXxeVrEdan
2GjouewPY0EwFWSKw6oIIGNyhGSOttpKtL2tG7Xw+pSCgBauo+TLI/8hcVYL2hZX
+DFXpoeNZkenX4F/1RWHZjPx5Poym1VkLKFJpjkD3v92RgbXI7is5A58hHJD3oS4
VyO9Y/qFYz4a/cHjNO+rmI7D0n4h+kIrmtQVHzpgwSk+xkiE/pbtppRs7p9V3/KR
Y3eyh5osQ27V4tU8m5QVh6p6JxALvXanmbBfJEyFneJ3q4RZ7/MHaSTFaMnYYlOT
264U+VA9owK+Rj6DCLQa5Hb8tjAYNiHxQPc6xKXPfVFVj781ru2fvr0yytY6saf9
/KZVZE3+KtmADve8X3mdp8wT8nFQMO5FSwkB4gOoCOOEFJadXltAy/nl7JlPZGRS
WNoJEKwpefj3Vk76SiPuaIhfzzlrEIp3HNh0oh9GUdTJF2cN3Xo/LPsftpOrAsMP
8X/tYM0NOzF+698uagXYl8mzUvqe66o3wI0kbEs0ra5YzL+1GSIiTXvOfjUSTPBq
WPaKsLmDl2J6MZUjJhY7V2bZy9+F7tLry2lg0j80CxCpzM6zkPBdvboyVmC5O7bV
wIrSg9obqGf7e0m1cZuyKg0Cil89Whtz5e4pRQBGXQ6yV62etRaeX7pqw647An5V
iZCB+FUWjw7Rc4BdbZuw13+F9BFb2EHxKLkCE7GBVvrrTy1AfP9ZuGUcbFOOTgS2
HEobyoViJ9MWvwnOeb2pTxeumkBATgXWTqskwOIE597sjCI2r4EIH4hyf2rpW7So
zjcLinGqp30hdXby7DD8yMKS4VB4v6ncp6qKj6nfrWCbV0XVjc/7gJg9hvBq6gGo
/0XZ+BfHf4YrY6g0wwvHE4nWGatH0QHtsz711bQ2bMsHpYbTMbuVhIq2c1wX5YGo
EQJJf+G9rL0sa8W7LSh5wIiALXzu5zTmmzPioDVp/SUNgYDH4wQ7KVZA5MSxYcNK
iX5YZUXtpM0+qe5lts63NoCnBsZFZmIkgba/+nq+sfYFwuvQY1GhcqV59ljIXSFp
tiRa2TdeGQ9MZIAn6UnV9EY4eC/mfzzbR5wXe7YpQ1N0Hi1xoNeI+YV6CIo1drt6
A1IjLUsE6bgjQ7XKxxKqRwyzmlyl5eMM1yOXv37NUWkpYZV8UYpo5ulExRHPmFhQ
IEOXfgegX9PHqgmmBPzihBxy2XbTIdYyjmcqckUx+XFayNAvMt/2C8AXWz9c6+wp
3tgMjDz0q6/S5Q19EmGjHqMJePvXqturMNOPeobjvoioPirTRIQwas27xm3uljtz
ogVtPYSNBZnSD+xkURVLhlh9y6SIdw8RERgdv0CYDEQvO4lYPvj6f+qlE8DVSCnw
weJ4iuu9pFEPiP4nBAktZ8JGombcMdfiSKWXw4BC7rOGc/LKI+N8KQ9YDmEu8pBm
j23K2OO8IylLcpyHJXD+JKxe+sI4UZenRh3QaiLbb9XLAHIvyDqrth54eeNJWBxc
iD/5kkqNh6K48DIVJ8DnNUnuTJUBAurhubveWltu6qEjyngbEEnh63i/7+JmdBAq
JIsFhj+MBa2xfGmkhHc9qKETjbPenDQWy4CuqDzp3Tl3mG39ml96WsVf0wmAg19Q
OuCPKOEXLJQctx8muokoGSxPQg5p66NgjOl3BN+lue6VzgeVnWWXVCW4VOYi4THa
cab2D7TUE+uoQGMGGLu5vGQSpMXldhyrWlXl1CgQxZomwkx6ot6lu8gd7304DP37
4ekE/mRj5JuSOYTiVyUZ/nulnAqNHz5AfZMvI2Nytwan9nP4QBNoOaee0eMDuENp
n6bS5M5sNGmwkIuiMJBEVL02VZvmaVdsHr99UVQuFqYe15a3Qz3PtR06ameyDR1T
xdapB37iasRywKd22g7nOQryUIdp/ZS7a7z/8hkPKPucB9jrVaZqyq07zu296RFu
rRgkclC6QFm+ymTEL1zllQk5aqC5NVJs64yV9hsXKqJMrKKLRG6ICLlDiUaAjGJl
gLggc6cS2pHPzp1GsBKXbCH9nby6o6xAYy3IyETMz1HrhQw0wQjv6IMs2XORDGx6
bDKeP1vXroOH1ZHCPB8JVYOpv6x0HEHgK4rDkWJbfo0AJWMjFdFr5r7mtUsabWGn
hTQo9lh1uZST2N+QEAQll1kdlUANFwQToaYSVYHdBSkqJaD7lIq+AAM2IJoR7u+1
tfITZ/JWJYe5JbXzUedBnhQmUB7lKVgUvA27vLZ+++K8Tao4FSjZOaNtXutGmPOm
Yw4NjZmECRk9J7XcuNxuuXZv6sgId4kjxvzFxA7QL23qYZqlgQoaMI2kbhKB9iXI
g/hhZ35rVED7mLGYFPIrmTauBC6d+4XSxnmcfvI5W3aeSB9uSB47OJOZ7Umeri4l
GGLwAXY4xDsFXIwISMaP24Fs1iSKoXMWrMIUeKeXFJIcGMMtu5VOKUr/lAExVnwn
NF6qdhJp8oukhuQpm0UAIJ0SZTTYtux1CNA7/IsOnLje7oOmI8awXBrl7MpyTZS2
XOVf50vHKVFdKVq67p4dtnhwoB8C65jrJYhkUlgwbEAcgSY9YO+6vcsX207fY6S5
O5zlV59flzuObuUQ+RvjFbPe+eucRrOwY13gpyHsvZv34qLnVV0yhASabnlx/RcR
Q1FX2SS4/KNkiBvBqxM9vAIaEJzR7xjhnSQAAJebiWvjNSuM7D6R2cQjQZVb07bQ
XXpQcztxeNgAjus5AHrDcFS5xkZThcCe6ojEouimgC7+EiV/gtiThRWIXMyXKw4t
CgEv79a+hyLQC6bW76R4Q1eiApC6Xw1YjNjUx5+oGryIlAKNi2je6ifwQlqOig62
BrRrRXo1B//DfsoEp1gU4hDuwOjbDH5O2O8oweP7vc+QMsqJ9XQkIV2q1vkzmVWw
wu8B1HB007xx5HlEfHEyLrvbMG6/DPoCm0Z+hE+drPux5cz2M9qYu9HZWDEIcRHR
4+vcFgB83YJZBWXOQcvN/oF/qrfkV+OPPQ25js9tyqb2UI3D2mgyRJEWzXabaUoQ
2gYuOoKqnaTK62hKJ9n9LgEFpw7+R6oLSe4iBmPhhKn0OOFIjk0PlHlBItz0D1Pi
zN8DIKr6IZNwTD6MF2OiH3o8d5FiEr7yghSAfLt+RCAxKUvrxspxM87zdLRk3HhX
S1BrV4EUzZROrHsy/0lIArB0GXBSlFHP6be6hrTuEY+woSG+nPYGtegLgfOMkQrh
ugiiL0J7hJr9iZJgFAVEwMgmtHqyowzG1cjCDePkVkikHPXHrQLX9AixXPSYbKVk
UDTThRJDLDH7zj2Da5I3JQmr4wpNYr4u7foTDB4YLJaTmaPBU8TckK+U6HlMGGcj
Cm3qsedn+F8XMJytAjbpBhd28oyiXDx7KqXAlyzu8aUCo2mXa/zJd4QLCyVlWGOi
raowGyZ7EyTsgze8y+r4nf3v52kb6NvxjpxbINzOyr1KlegCCyjedfRkVVhUqGzk
IT8hVxAgr0SHcMNy6V78BtRxJHd8mCOFfRebXexKPbfO/I2X50o7Sz8aggPigckH
wpmZotd5rmfOib9C7Qf5iGnTVpEsa36JUGQjBXdWxGFko5rfN1jvUkM5ghhwI9AC
MP4qkL9q0cd0loGGMMif6P6Zpy6NDLEWzgNb24neFwon8Y0+0aAuMW5kPBVm/iB2
8jukLb0bq5vPjQYlmcD5D9rNT7bgEh1Dmb17kgFLMpRewzWc3lgZhPQACLcpMLnz
iUIYzi1eyFlsSGIkXH5AHBfdmnh2eK+yEARBi2wEP43W5zko4hv4Te3Sh/EyJHRA
woarTyvJiMune2qFko874mObItfcHNgKFnumOg6AAfizZk1OPdzoeGIRBuPrIix1
BeGbusaW1ZO55R2z/YXdr7+0SHtUJ9WGZaCrQacw0kvhOmcw9zEmgaSYfNyNgIJ/
KZ2SL16lR2hW3VvjAMjIi9GlszPfgTYks7EDKxxDnNgLctzdjbz6EFtK16wKCRHL
QMTUikYASPc+OO+Qh+3sNrNezXZDQPLPozme7XUPCLu6Gjy4DYE5kh5AylvGWN0z
lV5b9mYwBWnjH64awHQskmGrUK+UH/RnRL4aYAiNQSXoVva9FYNRolwcbr7FoOw5
ZQz+g198XXG4TtDA51pJUADmPOSQA6vBjQZLsXQ0l/B5GOaQcdjAkmn0bQau0cLd
Fc2TxQd+Gtzl8xg1O0yWyTMyYl8Ti4leU/qTjc3r8e+sNKNwajulsm5j/ejHLe3V
2jJWDBHEg4wmlYi+kfljJkv8Oc3tXefrNlbfujZfn/4dZGvxBfTUB526LLCamKD+
7tSMRh9f1Kwv55J1lVkS15CTBqdXcsENJ3uM+Rj46b8MHY1wI66refbnehs23dY+
xn7k4BQWJBkgDzbB6slPjvntWsQlrrWumJ5VDIPPW73XMLcT7tIfZ7ckUn/ACJ3T
m9DtMsauqL6wodl1MgaGtjQ32o9GG9Po3yQhdb5+rKvcfwJJpCusd2c+waV7naue
yOZ7ucaErKvKWUKbkfKb4zXq6iEE+JMUbjjLMBnym4QzfIki01FVOZ1fzkEp8fBD
9mE2N2BrV5jpWnrKXyzWitRXyvzpKwColq+BLZms+NT2dMJf24HFaFXh41p2lQ9R
PwmCHU1IRuUWagJdFBq5UhIw98XStmKdbQY9/xWTX4NBoKtYatJ5LGW+J4ozdYxE
VBB+Ut6LbfELQZwGS2fDHhUPvVm/eYq3bfa+qxfEVPW8AeYKGTQ1VFO0n2ryvwFr
EY0Aur65hFOIphtJOiB3biw7UKmxtNC5CaSQLbU7TXl1LEwqrGOU6hs3gSvZX59+
Ds6FDzCwpjqHWli+COnIGWZBva/c8Ao5Ox4+hpR9mz6vNmUwZ0FhwPcEdicZNINn
QwseyKsvAnIakDN7pkWIpNgSAq6r1EVl/WRbmSN8tg3TrMTtoI/+7a2Y8Xy/rJ8y
bZmSUcaA8GbdOrkYdOVNWSgbGb4ycICrtN4F3R70XUH7IoDUDPQL+UY/YHO1lfk6
R56oR4T7w8hN9JZ3SDvW8wOSBeJOyl2AzupQqy0epd3gQx5seXbabqR1xOeW4Wzr
doBy/xSKbW3Qn5T/hWhcUcVHSxLwh1X7wAP9bl6PL8Eu2x0Sk1F1qj7oD/k1pFxA
0LoLE5udhnOYQNElqrEPnQZ+4S32EiC1YjhiN/PTl8LgscIfYLUMSiDMNgt6N5Iv
1pApRzK9DO7QaLxHoL1kcs4XbdTXNWP3DLTu4rxYNMLvChsWaPdsZGGq+ul6jyfI
q3G889LiOKtoNmNcWYzec0f36kjlWm1uQjTT7JF1SLUD7zx+doViOJXcKy4v5lAj
nljHbNhQM+9S6EQdu3sul5wy34NHQUgO0aufsYdnjW4oB9N3MGOdNF8Q73/Bsz69
gXuFZAFpjvpSTQhjT7XkmK1hLAF5lkLrKwerGfUbfPeeCxvs5b6piehw7DFnu1Qu
eox9/ylAkPwJdRJQrJrSw2ZWQAE82kIm9nvsOWi2qkrilgB24NS7tewl1bVSTh7d
b4N3J8711gu1V+wEz/k2Q/iJnGd342WqBH3Wt4rojyh7z3DvSbjx70wBRZH6Al/5
f0RO+O1ML1ay33/qvJgS7c8k/ga7tvL9D9F5KmdowNC9iuzBHLuHe4ypWtC1cbnV
UKxRdrzhDqevm41w7y3leX3ddM1YynJbxziCW6NgVOsMjAbh6XOt+/rmmvtplzoh
LiRXRwe+BZxJFXH/nXjavXA4vHgbPAoqMN4ZpmRJDhHyFSrU78ikxOdkRTviUfI5
RZUt/qp+shMdxsmR7uIGPylf9YL0TN3HzKU01xdA18UbWeu8Pm/OKmwxYNcuw9+B
fPgE7fwJ4gBCKG8tCLpEmxnJ63J+K5/NEQU8NYh7kXD2B1bcwVpHPiY9Je39Gcf2
On6i7K6+TbnPUv9xzle1kiHwOSemr2k9jt9lz23kav4uINvr/a5fvrnxB8H1B3IH
rP2L6db7wSN9OZ+kkYG1GgfBpejgRlAz8RQXwmwoGi7XBdSPAtRML45GvMhcQLbJ
acgsNfbeNj2YuLtdTtBUUFmoqCTD0/zcz5EHRVa9OEgjTM52cUrGsM+flz5rtdtH
YWhyDsSCg1Ia0yHb+bRjsxdUrpLD/WckuYjhd5OL2rMN7F5D9dgQXnyLXAt8s7oN
6KRg7wI09VLXkXE4vD8TcQRp/jXRauDfP9ermifjTO3QxCvbCtIWXuYrpNSdYQni
m/lgg0JJqgRgi9DKQ7XIqIZ9SwWkYjUqDXi2ZsvFMQ6rEYkljFPka2/9Ol3zYMD/
rgXxZpMGvI1NL1Xip3WxJ9rSoHfZOdNG0AUYP3PF/TAYE49kw3mTZaz7jFs7ILSF
D3c0ouLqste2EyKdxSSD2FrJvgpMujgz3Gu4mL3vm19eZb8R4ZMy4TgpBFKmVW4e
G/0xIp7cMouRypLhn3KFBTNf9Fwz9HtEZjOEWUMSuIuEmmb1vYudqaoP//47Ljcz
Zj6QuzDWjAgrCzqMj9yqjBXRRN4S8Zw4xoVmEu2xbKRd8b2l5Q1L9AKnYnIcBLI1
DHkijvaNSvkiQMR4oSjr6KrlmJKQT+AxidrTXbED2k+KUAgaFWnskAu/3cz3r+JG
hvi/LfBvHMrQ1oE8WM15zIxrPi7z9JJ7As/TJ2l5d6qv3lHtzuNQ174OhPCRWs8O
C5PHOpLghL0oV3rTpNlNp1qMGEmHmML/vg483fyFsqiaSdZZizFWfGXyJ++JhwFG
eoFbx8Z+/5Qwj7BgaQ5wvY3erQbA9WTNUauX8qgsG9dRnOz7JqXZYyIWmDAURz7H
DJXntT048knmLj4ryHuFLswmzp4NzKzJS06/bJEaUuw5jGUwlpo5AnhPFEyLVYPD
AzRCRHZa04pdQNCMufP6CdOQgXjgHquQyoBgFPDxiEQpkBmX74/9Oc5Yf3O6ZjaG
XGcP2C9TWQ77u/UNcyATehay8NVw9GtWFTiyr5vguNoRlyJf57i+ZmNq38pY6t29
4m2dYZK168DSdAnTkFU8+e5eCrCpiu1QL7Sl0AlGEktuWDi0RyRvtaeXjO65XHtA
3lvGqs6tsIU3riFch9wxHJ8LtWU5LH1UYplL7lHIPEMrG89v/ZW/OpwQb7t+UJlU
2eTOqEOO7Zzzk6V8/gAyDrACK75AhxBkmOn53s+V6AexPU9iBVx4vgSlRBqNGJoD
j41IFD/PvfPedpXyBPnC/839mtq8Ps0PZQVNZ/KuDS2Jlpdu0qmjdG/5GN3mNfmN
GhN0yPJASJtfUFqmMUrWm6S6tA9Ns2bVDBSZvr4NOlRs/cQINkCILYdPmnJ6uWsQ
nm5skZ8dXMadzJlQvZU8p8r0oLS5OybaQctAtKg4DrmT/B7Udw+V0VfxjlgTumOE
MFQpM69PZHZoOctEg2WXaW9fP3kHhp8PIo7lBeGzEAwditCoyQ8MOyM/RjLFxyqr
OIusqLSroLKNSTYkXwVCAE2/Dqz0JxiPom3cus1jm9XE/Iu/NV9aqW6SHcLvrFN+
tztL6G2j0nqiltScSXK8PsZL0b+XBRTSNas/KkrG7BwOTUKktyWmraXWR7DEAHWw
80tD0QjLJP/qvOfae+qEc+Q9+rVvV86ztrTbwNui3+sthRfgxzqoClfy3FHXey+c
7qf9NHI2Qo2tPr1S9Nc3MWSIXKk5+nTTx/KuHUJGmz31BPMwGitdZDe8sN318DRx
+cPwMu9/wJsYLPJRznTi71FqFaAjiFtnSj+3qepYYfUa1PhwhXC4pJnyNXS43WmC
ESrcsV0Atv+X8A/d9XWtT0GfCFejw9snZA88zNrGveVKDBvN1xwesk1OZZemhf1L
fQNTkxpNwfprb23kvV4GnCea34b7t4vXqFq+op9KrUzxiRZjpmF5YLXAcCuj4ofO
DFnWWIUDQFkp0U/Og2t4vcKQcbfwnDq9cJ2sX8k54MQZWR4EWupylGuR2Tiof81U
PyoT/bwFpQ6fseP/uuXrVPVR/9mevCAJp5uzndjB3lRpjfPO5xMt8FKm4xclkvIs
pb05Fj4UGHWxrDOj95sKCbEdbRLGhSKJ3NIhwlYe4+tcvYTvf8r40ZfuxKpcMGG1
SrO2UvTgNgkpDlFG0k/EkEORQ0xgnKkzMK4Rau/bPoztKQ91aKRMTuHuS1mgLn7P
Ls/F8M9Wz5EROowNmRBWVK2H51E/KQCR+Qn7ftlpkxfir3AG4AXv/wTbatB2w+1R
F2YRs2VSFkybpAs/AWbmSlZ74YbFivTIw78vHYpfyTYjNwaYUY1bjJIsp2NmRDNl
7cheWGkeLrZwebZXgMlBmFbYCP5lrB/ao9iy6Lb4LQ4X1Id8vuLVsSFEw5US59sK
ShPYwL2LgPnZN259ojJ8NOF+ZpdwEC/PKaiYFP/Biu/BNKuOtcAKs3C8JT5u37TO
7xKjksdoNhRwh4aNpWU1W315Th3hzV7Lq+rmznE88hJSxq7M8ftg55N/c+1liXhM
ZeBXVXeGd6j19LhxkH5RYDsRDq6LBpMS4OmsI0UqujvMDRuN6aVNX0Lk3AmuA2x0
Lue7CGzj3J1D0iM6tyaWNX9SQ0mW5Ck40/TiMNh8QOwioxroY7aJo1NOhclg1YIA
2H0d7ZUOO0XQFGe75O3QBWa1XhXblZBIa/RomCJNU4XJC79Tmrcj2+xU3cQQWPUR
ZFpZH3nYPgDvIk8t/SlgcrEhYyDFjFsD2b42s8vhMawaXulxtpIZ7Bo849pF9e8s
4/okBWc+hla0XEtg+zVEK2A25MEh9JuQB3tJ5irN4mzXU4qHNjnn+MMvvnZqjvFa
DbYCnjUnxbubBZ0+Xye+RD8MqAd5fAATNZfUgh9z8P85tHt9xz7gCzBk+LklvsNz
VV3l4fIYLONnC4zaS2DbpKUatKoPm+d3M2Q3/LOEoEPNDNvkd2c49GXCgNuuOSY2
KcyTyckJiNAbZqIDjjcAirD1uDW3ej+IffU1XtmUeQdgUgtweQyy5UBwqtycXgxO
88OTHrVcvILS2oNjB9PNkmdVNAV2UTA1NyIAuqzY25NW4mwhgba7aBVFRLMAU/PT
Q8cGJG0SHqt4wCSV7stOeoZlmrAXws95PhMg4p6AbhReMbfqnGViSKHNXnTZ6Ifn
Jrc4xrKJq5QwNSkBmIyrnzOWZw/HT1v9ts2KP7ZTSaP/nHldNvLP5fUrb4AegTIh
mCQ/S4SlcmTsARdDvApKU0R9vB4QMw8q7Kiy0oFc2O179V6EpIviIf3oKoW1FkjG
qN46i8JHr06UPnT/Me2AFTtfxPgHcI6ATvYTGtF7RBBVgZ08PGsMzmMM8ASujEIe
vrSx/qp2BZPFkhQJKhoXLpoBrsIQzyKnkBq4fnjPeJL0YCAcIpp6S/cFxONfkG2R
VboMHNZAAyK0fg6jgN43EwlFzNFXB+7U/JNmYkG0/MO+kVsC1puy3JjaPVCLREvV
7RDUwWkWugKlNQvcnwPQ3ND2OoF6g0wBg4BGeYgHvLcMZCH+mJ2y0NJ3c8nHw6ZG
5RZfW8xVWPR9LsJVou18pYTyUo0XLO+KTRptS9BcLx73MrjRMj6E8Ck663cYVQtU
6F6ImuR0o6X5qfqnNfwHw35FesY1xGZYWPI9JTNN4QxJQ5M9vEOgtbOtBijFQYpK
hu5D89ov4oxd2J83allUc4ZY2sHw9p6dYrqyqiosoNHcaE2R7xIKrZ5P2UAPhCbX
A0ra5qv7gYP+Tgn9bdy9cdZceotz6cfn1EuOUAN34yjRwSb4PRK45++ubP7Yg3IT
AjEQd6lqFqvhr6bISFRNGOLH9dGVO01rqTk+6PrtsMSkPUbwUbqxqRl33EZc5zDz
ym3mjRi0zdrgG59yyAmlPgWTZve/hWPUB4FjZ1UuC1QYAFkr9Wsfl36T44038sZq
yxk9jcDCfdaj4RPNPm4R5Qlz0ezNKMAt3zdUUX9SRihw7yqKdTBfCSiP5CRrNoAN
n+ZIQe0qGHLBYeT1hass7GLO0brcCPsRniFtdhVJvEOtoL2IMP82ibPSYBfQ08dJ
7wXXEhY1sc5IB3fdJQVprdlU3oWefLrw3MtA+v6jUqT7kYGf6eU7LHIqt0jwOeGk
HnVwbSiCCRInH9lk/W4m7+ULc0x5EZpmU+flAyM7fpAmZFWicdvpAAMnhBPEawEa
s9JRj96hHm20CjjI00QGDvuRlwetqYD11RxTm2m8mdWYPeQXurvnqkeKa8UkJyd6
tFy0cnOlBaE6iYgAszoWJ+VHif438qQhtnqNdlL7WzCbV2Igf3Cfz1460y5mXO+y
EO96xv+WT9ChVfAS6SccJsZmgd5YSwfj9cgnKD+ILmFuJagPPlPqXMDC3uu95fsP
5qMfGPkxHhCok0f8y5aq/uODqpV+I06x2TtGoKYHnfs/o2VfuukZf0tnIrQhukCk
5k2QuNEtho+xO5bC29rultLWsc/0QIKJ2B4hz2QAsiqvsaIiJ2465yLLzdJextfP
55I/FoLVmvE6bNgYfyq5EQBEh+ZsTwCSW44QWuGYgMuxHhqLEqj+AO/HmkNiW65X
8GZr+akdA6lEOWX7K6nOVyYPF1jgFvWqIdb0zbSFgCIQv0PVDn+BKLpyE0861azM
32qz3yrSSRVy3lOwH4+3fOhEvYK3X5ONm1oWVw/Xld8JUbCBSLaA74QG4QtmT9TG
qqnQCn7vDGG3NGsgwJiICjjx1r3Vsgutg687vlsIO6nJlnI/y39hftzDqGVyA0KF
R/RKmpzILLveAKiMeHvnCuELDNt7BcaMb71RK684ALCtRKd+v5JieZoS6Fk2NlKf
rymzVg9EaLlSx9VgzXZYcCQqW7BkpQmftFIU9LhRwgrjXHc+vaq7r0WTUAttGzjA
nVIoRl+QggubX1kVTRwU6s5R3eqAe8Pg/t6qv83Hca0Nkw4oNY26P35It1AWkCse
T4rcwyefBf+WqGua8EVibmIA5mKEfGx4o2YIGyQpZjuu0xGmfuKTPgz4gOzhx08B
MzA6qbgSLM5uuqrjXLwPy1NtDEjMeN1EeTh3FGPJUHxtt1jgjxlF1sochHZ1mz33
7Agj5ypLkFsI7pVZYwjMwIzmF/ETATGC6gpsdgaFBDoBj8YdALzD1hxPqcPFmC+i
OEK94im1P7O5wDns6ggrrICD+5kqtPKPNDXCsreakyHg+H+U4bDAva6SzYTiFaDH
0sJAGMxMR6PltQjOzPLczWGj8vMITMM1Se+PZMo2kvQpxvgTMtifHtNAJ98ciXGN
jI27llRewQdK+RMmhxRVgv9dRKYHmtB7vCpBkTGA+5ZGcl0JnWvq6Vswd7DTXpDc
5R5ZOY6aqtTxOrrfOWTzSlAwCUtnwqImBs/sEyr2CB8U8F8+zEYwIc0Q7mTla1b7
RFH34wmg6ID5hk1nl5jDVWis6iiorc6Tb5Gtuy850jiJaH17qV3aK370dmwQ/JO4
buxtF/qz9vPp1WKHUa8Dts9Xf//APKxopY/nLxEpntHtxKE+wSNS+6Kqt1U//5km
adKMrdLAo3zgOHHdaRs6qvkdY5Un7cqM3M8zaGWpto9kD5/fLi2cn4anV/Akfrrg
hFgNt2xvbuXjze5qPF4nnvkxFVQzmBui3/GH2CQD5SdOgjaW8/oZ6palEbe+zKS7
wtJBNLzMeqPvsSPdu0O5AsTogxTD4JSuLyAOD+vUv/efr8znjdRDlGbMXvoYDt91
E+N2nUr6SCbLQJ1a3ah1sm4HyJ7eszX6LwNTP8+E/ykHGrzT0x+6k7Is5ykgOZ6a
att6k9iBlkQ/qW+vTlExHsQdkmsVz9FHZ2Yc6ClGHc0/O9PK8DJP9mp9RWg1cLFc
XmbdlTt43Ld8niWBwOnG46FQG9VpbYMD+rWFHQOD72Iz3FYscvXzH6vVwiC3CbWX
vklmigvxDhAPthCfnRn2Av8xUCkachm75FYkyMSsPNIs9xy7Oiw4RD3L7hLQ3pty
QSpOhnmoK+Hyr1k1w0o8FhHQh/4zBDCq8TKWozyTviHd2ClHSoV+KW+BuA5WhbW9
/JUsZccfqGeKrBJtgwSzzbHC14Mf1pjk2nDd2yOc2MRCBBtpM1iqZoM+GeJUL1vR
HLsBUtwZbs5LgpJThCwfbwTPf3hOL9rDOYfYmTSxqEMZCZGj71QECaPbXWcs15Hj
r5aPuIh2e4ZOtvU89/4tOJMu1H/lK5NRN+1GXJB9X4BX4ob0K5xJVQVun/TULWrW
DjONnRsPu/GmYog0aL6DyM7Nh4Bmq9FuAKtVdI2zmVALG5GxF95JoaAxlmAq9Pqk
bE61UBwen4igGK4UQ2AK7b8tSiA6jbCgGATXQh9/cBio1xhR/1+BkxOvmjj2ybaX
UfSoo616K5XShrIifx2kvQ9gal2kdjkqWOF9tp0hV1yvotpHoPsWHgcRc+R8gk38
Q9W09wIRFQLW5qmJoLdi45XxFC2SP6vd6AYyiIWzqqSEUOet1uRPBuDkXbpYZ5VV
h9el0LBvNOePwyXE2cdzFRQGLdybbtXOS3/Xh5bdUemMtOTK50rTeNHQZNWmOPvf
8BylTknpa/ICuaW6KmNqQ9+8DAwXq6eSK+JZ5IePUTek+hqAaMnrpt2cVrigWTgB
lGIElGFYVYzNpxgdotQz1QYPJowTI0+Jaz87wQPhGQpmAZDlwjbyUgC7xwiyYMjQ
Z3DBU4KBZsE6Vd0cX8huXZmCd3/DTM7yRKk52qg1zbuAGQa9612tF9hDA/f6sAy8
yMqlo3hL9KVIkdo2kAgwThY19e9o/bliT21yP/eWTE952VBGVxmdK/7L306CTvC1
Rzdfj9y/yfOT1t7l2RAjB/BQbj/JQ7bPyQBFIK4Nqt0+pRXQNp8pMnOTE7GvjNGt
jo81WsQ9t2MwH/WLoWx/acQceA10wFwaLkAO+HSp+Lgw+U4Q1gzfnx8FVHqZaGuL
e4HxmM+e3CCZEUqx0cDUcJE4N3S5d3sxW9knzV1GxYJZqofSGdrp/skwRB+gRzr6
FqhqrQ34B0fos+TMeW7sT/mQHot/VhukFvJXYG9ELRHuZ8bx+ec3/pnRtdZViQ61
R0GbEQwT5c1HoJD6pif4UvQB6A0TlvIph7o7xcgIJvoCex8zpU2H1u89Bzajhixq
e9+XKkNnOYO/on1m7POxp6mcO6LPUbgUt89ocRqMvh95DAGfClahU+i8Yss+2TGS
odTvGplVyIdeMzyx81p4YH71Xp2F8daYddP6QafEwGxKWDQ4fcSOY2ELVRg2o4+p
K0ZrSdpJ3WWU3v1cZ0YDBF8Z3eNeJzduBMtrLwLQRHGqklTNXU0x6bcB8+ypZTQU
IP2bYoWGsJ/tfSjMP1IEdqpcGz6Bmkw0tmQgPT8wFRw2a2pNXrWRcx7YvSK8sC9C
zmcn244EXM7FDVqS+TdDtvTKqAr8mqeMPCktnZB2tDC+j7PaaECeuN4/P/6qcH9A
vtRVnkGnstgmV+qiWpKpPQ28uyydKAGrLK02Urb+oH1Es1QB0D4tAtrTcZJSDZho
fGM+Ed3JdEUK33VNUqMT43Q2BqrQ2BBz0bWJfaYxi9udsuBlKJuAXaUynKUdGpER
2bsq/8POOfc6P2XZmWXF7bV68wTeCdZCBOJxicivxuDz2uIJIEv6Hj7a/qL2SIZm
nEN2mTG4gPOOvisDtnOZt8mGVOj390q3uQ1QSfkjwqfPYLjU9ocauPmmzqclA6jt
usZAAn1UzkX6e3J7Wfq38EW/CtwVhI+lCjlgWTDEAfs2IRKQMFfrzSJ7/DhGNoiq
ZffAK/FAFlj3FVmSbtJJ9F+VhKGUgroI8IP36+a+P6wVL1CGa/jGniQgNw6oXMjD
UpxRs7EqAMmbQbxkHSTrkODSt5YBFpQ0ZXC0SF9HvdTaovZ7P9P3YcdxnOyzGGjd
ZGBQwWPJWjSNoXAaIwS5KL1/jErh910BxzmNPLNzSFlvSykSgwY6kAALju1ZcLq0
sAkGTAWF7OoicMu85YrqB26RqCbo7sDfBdYSWLm9atL7mXKjZ7xOgtHDTissVw8t
Kkaqt2w+o/23L1UItxUj7pepf0KzUTPBFszRDyA5cm33obPbO0ZK5rOnhIil6k0y
d7/o15MpaEQXjM39caKxgLT7Yv4+agi2UWfd0krWXIm+rWM93cf7mHD7nP9Y/wm1
BMysDjd/diXrY9l39WQWTgZGNG8AZgKoH0IbMdxZz74ZzrD400KPVlUSE6qHDPLm
0YKKoWiYeJMJC4cLc0M8r3aVcAs+8iRB967WHuhSPZFa8gWAebblc66otmhBUtYr
L+QtN74JhbsaYiedzH1a7YT9q97wb0JmC1ngyRwCBcfb/IATJZF4OI06qnHidM5J
4XSxJK5gKdG9NqaEe7a1+3DTb0Bwwb1h5fv4ZB7LMt4Rdr3RcgyHozThMRP/t7lO
uRA2UExLIgkZbeWucFCSG4y5g28R35li8GKBNTGgG+l1lEAkpqlCk54YgdZ5GM3H
wq5sQi4B6TFGG/na5bMJzJYx10JyCg/8bhTTWPrIaIUkc41IQfXCIqC+Fo9XUGdX
FYjHEeHnW6kJBM0EkoupXqX0BD3JBPXOAj+RMJetrpF95jz8ZKCAPyaQASwuc5Jp
HZInN5ZtPHxIq5UVpfzQGnrWwlka+A0BLxytGyhgZJEaQM6cm1Y/g6b8UKDqByc7
it1uIRKshx1MwYrGCez8NTJx6AwBUVMmoc54nT+12UL3p53Wntp2LJUqeqGy5Tk2
2l8gRWgarE2HZkY6yK5p3n4z83I92FSbnTze/v9t8YH+pIGWyF7WOuRb1ntATfCL
ccpU57zKldjM5d9hwdYbnFwZAwRauM29VvqBjeH2UbvJAN8AJbn36wrWk04fmgwK
okFUanPFZYwdzrRJ+zNSIvLnL67uNi0Fday5Zy3muxTL7jpu+L6PI3jCaGL71psX
s8Vbnv3g9BZTuqJXTewdL8ec3BDzskmmGngZRcI0zqvuaB+M5vStZ+5adQNEsoJ8
CHBcnJ7r58PH95bN1MI/saCqlDicvFfXiE0/fL7D7Uw2PIXwautewuW7Y7bM6kOu
kixi6LBrltw7f/qehyQL6dK9XzpJQQB+ay5UX8My4+jrSSI4ZagI5IzbOJ6t3oi1
5xMhVC0QVFLkW89sM+sYMr7Lm47nhLKglUZ+iLy7DxFlGJl+wl5ylzkeNEo3EB/w
lPfsNmftzQ3kjeypJuKR24G0GWLG10Cjz4j5jKMFJ6o4D8tRhZQLsMfDnlHBByon
W+qE+ZeM81YnhTgf70uiGr4pGGhRt9bhbHvVuHRR+EWINr9sy8L6rbw0/XrvOnEb
yQAt+Qrxd6d1i4ro6c0zItDMaeFWUhQXUWdzzuxS0SWIwAmPSK78Os7seVkAI31+
cAJE3rDk+XOKZbx/49oiwyG9jmG34Z3UejKoFbsdi+aU4oJzLkvWUAAQF8BapPi5
6y8jDbPIYGvqVWoWaI5QWKoU7ZQRphK46xTe8zk0253Aco+UKj9NT7axfLB/G7hr
NCOobWjKp63le/Lc9Jvfr5Bcjb39NPThCg3kTcsK1PUUoTd6epRsSsfkeIHLpZzA
4pg4j+fx/nJewCqUL77fcl4MBze/HdTtuTA8g8EeE0bzJL+daEFCBHW9cFOqIcI7
KATtXxNDvpiLFHfgPfKl3yV8EHjkq4Vc003gk14BcrFvEfuWoAwYy6X+CWiWqNbh
O2ZYrT4ZhM+EP3XDng91dqBYLOgrQbcbpsCXBI1ZDd4gL4UEYuZYgFU1M0uPW+t9
XHMlCJilc6AzQsRY5bqtHrut0NWWqgBiB41ghnb+D0lGsSJo253SFCVfWHHTgPYt
ZcjwIzu14wM9HSCR9+8jSpBAjUZmMEtfBCEoui84eDxMOpk89xznlTkD7wa+a03J
Vi0K4G61BoIqD7+HaiDnIPnqYEcHSjYclzZJDKHaSMyUBGzaBaCLHnFxkDESDQKS
o8uLGVWv03NJ1T8J10c2+FvVen4v111jPP1bK9kkfdv96Sdzz/3uwltoazpW+x+H
Gb9YN8K3Vp5fL5EFSy0Qt794xLq/YdmPxTJwI8/v/PSpFEsljmDYW4kg8hTslYjV
erJ9cx8nyugCse9rIiNZhd9LjVYnr4gSS4G1TgfHhgCaiOGCHJaM3yo/fPFbix6a
ZNKT1HV0bWcNQpgjb+ftHfWQtvu7MZNXPFhZqDl2ugXvEmtLM6q8UsFcUEJYbYFb
kO8aXuwp7IUViXKzLxdU6CgcsikJI19Umup3n8heA09hiGxSfZKJ2mUIZr8tkriO
zhu42j4aROMxkml2UMjDZnzssOmX3vzb97JOs3O+QrAz58Okxuq/HlG84k/uukLK
niGhaFzx1CfFIrwH0z5N4XEhonAg3EOOogpbunJwO8IiymOOJ5Tmis1seNxJn6V8
CVSJntajiCYwUFlV2wGo2XP86vuZBfgvtJl3XLyFNiYy5GpAiBoxpLGjfQ+/5u4A
IBDg6ZSbJweDMlTGGXdIaP8heirHNPxJaF8VwC8W6kRdFRct7yqnKFTIRWy8YYTK
hnpPGkNGC64lPRY7CikE8FGHNM8LeqB+NsqMeQEkPyOpSyvHoW4ANGud4wNeUVD4
e1OTNf42bKpLSaejVopEmmKgKWQOKxex/IOZiKcjwoxAAW77vWc3bt7yWttcGbR3
8Fa0yuwILzluumETFUlgAz6pR3E3YJylGjKXoI4hmvpA8x9uUrNDCL6YYQm8KFnM
IizCgpIdA2A+9qGXFJnH44K0PFXA/Qz3qBUgVhMN7U3yu7vSMZTpbDgd4stfqlEK
KmHCc/51R4j09IBQ7GuQ9+xt03N73YY/PHO9G6k4m3rFegNTiCA975dImZDov6EE
TD1meXmD3sAWvcoRS/yc69Y7BQ8iyu5aMbbzqNnYNSvXkoSioYnLOP5c1bgLQe9a
h+evNDHxrWhEzWGkuMlV9SIOwFMVGcBamk1Xt+dxxUKXC6NMj2gZy3BX5MxqQT6v
Zvh5L2+nZ+8UsllryG6HS5zYIEpx7rbxtgFIGIGSMARNY9uQ8xLfRTigqaH+DG52
S5UPUW2HjdprPJvdygqAhJgtvSP85n/xxJZQRQWPvfhRyCwMxVmaLU6Zl6nL1Jgq
opzOV7K3XTpUf4M0NI8kwqGcIrNL7y1Oxa1vluMTf/jfPG6oT7RP5MsHOGsPuU/F
59n6p2oIvtsV5zSbS67uuotvDMARYyicJE4MDSem9daPV3cEU8T33gy/iPJQtyx9
Y/fpvTitskfXpM6tq8YZCdiqM3CMMoFozQzNyyPvQvyvMD12xNy4va/0kJBCdTtH
IWX9dLaEW9pn7vD6JlPymr1ZqC+omPDv0hA/kl02dSfmhiaaHYmmn0HvY/x97CAG
KqtUIe/NAqCleINooGUrxLuhDV5tgnlbRTbiCZbXoh8KeLcdzys6kj5yVUTO/76n
v3oXXj74giun/NbOKbGIs4SfzqgmgBll3B+mzE0/ACmZuqmPBD/3GdXPSS8qSY3N
0BvMGHCBX6PZMXEHzIifyONyoNK7f9Jg6moyncWIREzISVwGhfViLIND3jP36Sb9
+jk2p16MnhQUkIjW0FTX2EbF9PZp4nLOf0gK5iiAjtbfbigk6DEcOqpWMU1pr85K
0qFexNiLWRrTvk24ClFndT0tLyq9v9FG8zdyTg9OfCZZcjQH0La6PjQf9l6dTiL2
jzpTgpqnpdMbw4LRPTHCi00/fOBTEZcB2/Gez/kbjKXvcysqD4zG/jkVQW12VR0B
02bwycYNCaKk51vA0J8KP8KHnkSPrBid64vz0ECTeqcSGxhwZiH+Yvz1IIfJN/jJ
ghPsT5cvGIkiceTduAQd4I/NdawtFl4JUp+w0S4njKmbLHFIqVWbdghKAOWEXX8K
6SVfdb5zxQZdyMkeHcCWodxFpm+/wn+zwBJft1CWX0wrU6wIE9YA+DO+WqziQrMM
3dfJqBUQ++/re1p0nbs0Kf1r54ZcCe5s9ptSxuAx6g5B0G0wLqR2VnyfzXUHjnVM
cn7UITaDxxTSgOmMsyr822bbQ96zchoE1gwQ9gfuQJn1UY45rcOcibRX2qamI5J5
0DUyLLmGJsb7pH5Or/6jA+IZWoVbl74h4HR56NUDwVvMpSgZrxMoQ/q1r27O9FuF
CEFaF9vNNSgbo0hEyKkQUVzYgOlT1QHkNbTuejc+7VTVnjQTu19q8kWnck7MLvdj
0MSHxGiYdWXiF12YF9T7V8pdsO2N2LyGsk2H5rF6Z6gYuLtych441bRJ64wI3fg8
WXszha3u3wghNoN5adTeEKR5rN8WCZeI2xk5GJ4TUjSW7aqyqo63HLXymGzEuX88
vl1uJiXagPPuN1gkbTenXMzERo/4ixw9JJpFuzf+pa69wtroCsX7d/7uFmO3Snj9
SMp5NoilGojljYZt1O8bjh78xbyUndWA6sU9tEp8D6hJUuXbjgClmKbEoNR160TH
o5jzcDCxkbW9V3z9/7cLM0BSjbCR8fIlrsxrZtMUS60mdkj31CXiIXV/g8+t5e8j
Rp7tNW/iJKTpL+s7mRCnH6s7BoprxYQDr1rc+mvKf57IoklIGMg4G34oMPfbzlGA
qhrXzk2nI22bP7pMG4iDctPZwFMPdikI2WucRG3Z/x0HLVT4gzyCM6CCkI9skRXZ
o5NC6lpJdKS8CM9dNHyp0zw2kxEbRslq8jOk4ak8BWPtvwe+b3ghkQRX4tKN4bmm
2DyVPEEM/Cc6XS+jhWXocRMkkoYLdBqxoycr1vd2u69qr81DnbPzwWPsCLBuS5DU
Xfs6x8N/lN6UAZGC76MlX91mQ95b8mjE7QFhHi4vrzRFi3OWSWSujXqKbPA+Uwws
bh6N2GvPNOfD6hz1JaJ4AKRP4oljDwaTcHMyUdP83RofwInBvewiCjULM7a+Gymf
fisybVVFsVVz9RvQP5fOot283X8/U7p1ozoSWBhDqFacmPTpaprdCWHkSqKCbmcQ
R7CGICX+1CqbrHTomHtr1Y0uvGXx2a17tZt67kegGQxeloGkMmHPB7uoU0p+HnR4
BJ4hEboLVSafk2sZiM9Ezmq21b9kyDWYrqtX35wVYz/+Dvj1rwK1zmd0qfPjaAoY
qcFwIv5av4vgV0JauWNytQoSFcI0nUfG8LZeOy1F43L1Hf1VgI/XC4GMIo81sn3s
o5CB2RL1YTZzpm4SoAaQjg1CjOVLsuUYeWZXyVvMQDbye83ZlOB28c/1q31Y51BW
+H7VFth4tgu8SgqQUlTMnurgdkqzfWjcrFGflADqOSa17Iw07RI9SgsqFH3gTY78
UQ31om0Kw5WXAQnzBHia08pRXGZG2T3O7BpyL8F9kaLECkLg4ukTCarkw5ovDAlR
93/Kreh6/uSR+CM+OljprcU4Nyc2clPPRjNrBUwxnuTOasNEz4ioLh8qU8qfYSE8
LpLLJ9hR8pfU9QOGHVkGK1KiujzraIBn/1Fkz69i2aIApId7fVyxaqceh4erZLEI
J8lMgsIoDe0PjE/Oq5uxX0o23w8PZs5bxQjAGzRCY/Q/hVbbHJT5aP0ta2rtnBdD
XZ+ZbBWSgsTDYAYrAkLfBplTFkGdrMHq4YfLeewYpTHZde+O/IO4e/FxcSrHw5rC
y1Z3ukK2+GJnpWeJxa9l7ZsU7kIxyZpEK1TmT+L0k5ScLT2GFTBAJgHBHLvZ6cyz
4yxp/razr6hhL6gWZ0Xx+eZEXlKoCld0bm+3KsWeRjYxC4SM0RnRjICx1hJ5mvdV
8f2GRwl80GXogQccVHjv9GHYMtGAOtvERyMGrazr3/R2WZsd1b6WCd9V4sqng+5s
fmmhFvcLLfsIO8FKEmarMGzLtlLzX6mj1Vg/+mkkZsD2D9T+sO2ncpLKXh748zKL
7CKrETHWaoG/U87aIMQ3oeeOGfBpSIP4xr1Q3vtFT86d4Wy9m1VAWZGmBpfvhlKR
3aVa/NVXwyU+fCg/MfruOskhHDaxbDw7PlVgOCcyJtZDxyxnqUkzpEx1kjFdLJEP
AIdYAQw3vp/GtLRPDtzT7kNHHTPgohAYVonbUKKhQG7yC2kJkK77wMK7+p+8/D5b
muA0vX2/z1mUDYnadJDQgQpKQqa/WjwOGcDdiEHfCn5cv8nn+avEJWsr+BgIqO6r
3h9a81eNUbRTWTSYjZyWoA8h0jMSvKs2Orh/e00v5/38ZWEF4v3RMPWfdYbL+rfd
TTGb+WJo484TaPQmguCu1cwPy6QzkQKrggEAFbme50pBrLRKqSXISLgkr7ISiL5G
fnP0yYRnA6Pz8r5V73KrDhxr8sqYBg1uBGSdIjSSVBI9l8YrTHAGFvA7Xj3uuK0l
YRvPVps1M9UGdYuWSDRMmh7EZtuQMOKqdy8jmzKhQxJvv+mvpKifFN+jQjOgJ7eV
vjrZu+hTua6zOycw8+gExYZPgHn9KQsbNJT0Fx6peWy+4vpE7PhWSEpw5trrAL/t
vHn3sGnMH7IsVU791W/f5iKNpZpUSylZ0OMHLwX4gGJ2IbtSHQy2rrN77+FyH82h
yyQgOMU7toxUBAS0lXRvbtzCr3FHex5Taq9dwi3acCMeeUx0sbcca8KHu0DBQ4Nr
GyduKl0s1ia84XjGFQxrp0ulIp4W3X37l1qiQRqDes6UFEHh8KM1EWzLc1iYhtb7
aYJVC68GS3HrfiDavbd3qY4iD7SWc89hg1P/oW2J0ZDvftPXdSsRAAdL5CDGLCUL
s/cF54wfXXFV4evJvJ1jUhJxRieQWMJYw6arzG0IllP1MFET4ocuqaY6Nf6ryIm6
QkFZh5dHjdxXX4WeFlI7iWReBkZu9ltJAnoTBSKtm+gWWAA8Zr3mk+mPDBkoVskn
W5/pKehBRSetqEFL0k3Q2hnA7J1UmqPsUk0bxvv+uTE/P1LcVCQ1tMHGrcWfYHAo
Olr4HW9+/6ABC3+VjsXGHhK+l63q95CINeQB3s5WyGf4lQg/FAG9fLkwrT3fdeyW
WhF1ROyBIVMCsjdIPv/fIcLRe8INDdb8ovpeZE8G1G0A1Z4oLImcUHpATicj/OOw
ryBCJqmhiwiEuqvRgji44mRB1TXmSvYs/s6Q8i+U5/+w6GkaAFSFGwSW4NV1UBYT
F3HvVvGO1Af0zLcmehNKlLrdjU1JHfIlzhpMddpZbWfzFVuILWhQHVqma1YLNaDJ
Z1W/wknK6oEnusbcW0hR0JRIFexcLG9bEWunMQfoJOLe2xj81Jk3ZTt4KTNXcx5I
7+mC8B/yYrqKgrFg6rVEuS4YIhnLXXJbic3jIsN94CYsX73nKGNCtbatR3yn/BjS
fDbTU35IFxbGo8eKBo3j6sVBVG0h9yPVpAjry9VYmhwY45JE8e5CVh/xKNGRFavv
Ml8yOp0k7T+vIV2Go8ZLh4rJaSj7AE9iv3+3HOJ9qZ3NiDK190obgnApGYAzb6Ch
CPMRUlsYheoU/4j3EOLEkTJzwi+H12cJtXrOk/QpW2UajK2Ad8ueuDonb/qY40mx
8Aoyc4J0yQQhQYYr0O4DLC/ws6wf4PPdUylOheVXq4xVky7w1f0O9LvRDWqRqOjC
vMBcfxGioornALB3tdAod9q26sObCMd5JIJCXz6UnFNKSr0pWt+qKIrIxgGDC5So
EQbaFusr7nvDacTECOZLpvUEPwQLC5bEAMqXROa87laLVO4uT2Eeclbl2EGL8K+1
WR3neqosIH7e9TPYe1CIETlBG1o79kgOsUtw5V89P65z3gNKSYnSxpGJ+Quv166f
j0WqbXqU9udSJo2VMyVIlKrxXXgL7I0RVtxgoAATgBxgTq4ibSMUu2pZXCivwD6d
wHvc1Cb0A67ZgfdZcjt7TuCYAeKJVD1OXakzIORZC5pnFHI83sJt+JsJKuLJ4Oqm
8U0V2qRQt8Q9qVSZQ66jHbrpxcU1GfHEXGew1l4pcqKvpDjYRLyRsZMGGCKHHAw2
KU9HZG/2dg1KrA0iPS6VBFy9crr9zT9sjNL/MuzkL1XlsjndFblmmr5fNT7GJjM+
/6v8fDsPMnuF9ixKCyMKpDjO4jx4AyfqMM1xSDkT2J571be7jf9dm6jK67BfefAW
m8pMTrSrafr7BLzdl1Se4PHpl7G/vEgjKczr5s11DbSRe01jD/g0Lkvl8JsWLBvw
AdYG5Sed77ILN+hKyCUeCrNjSSyRzYXDu6G5KIZIk+p8ap9xAVTCm3BgnCb5JyG/
NgJGsHCQDn4QtSTxXJVJUROsrxiVYPf5A4ARMGjSQF4c5Ddwbm6DN8AMwvhtJKHA
par/E8vU3w4tksmtDLhYZBL80CE8LwdE1Q07le35Je9fs20MN9yje7GAytOgAix2
9FHJwMAZJGF1VqnrM/1zhoHvhgXv81AR7wdaRgPrZxHtR5zfEPiUpWN9kH4XDxm5
pcY66yBzDPWqbAUyjhA6EI5IW7vvokIStKG+DwM7Ud0J7mehQRDoZXlvDRyg6FJV
1okHktKBUgZh0fk90CRV9c/AI0CStYCiyh0FSSQa9QNoP1yNsgJUuULAUQsrchx+
xC+z78a17i02huchWeVlXjbRPVQEd/GMRV3+N8KPqwvwMYFI1EiZN+maZXL1uc3F
AGP3dC82P8BFjM+a8meLInQ7Z8V+GFA3L2kUZA2mRZV60iQrFaL9Q8tPEiYzvE8J
bUisN/WCEO/Jzw5fN81yLlbL8LngazZeGDtLz5toOQxLWqdCyb574FBI+Pdcmp3S
qFg83OvGiRtjsmqFYHhFgf7E1cs++LECzdoa+PCN/ZsXwIPH4Xj85dyW2u+pCv+j
XYvxfkCzOKoowJwYhaIkUjUm6G9HtdWqA1LSHKglnYZYVV3EwW0bWVsZTKPxKY1A
4kqR7TsFOy+39TMKSzM7XJ72JgUdHH2w4e+1u60lNRtnmojjhY9stonnFY7Nogfa
b4cHbscgIRuJZ1ikol4HjDH/j86VJP266X366Div+mpk46LSmqFgxk6Yq4yLxYuu
7zIuggvHffq64NwYgkJnGX3L6Thre3ePq6A5LbpjgSANqJP1bn/Cu7TIlICVZKyR
nRV/+05iEpvZYy01Z4bAe3FwU3Eiej2oECvZtsmAvdEmJLzk0aiZb7It+8aR0/H0
6ppvJTf0tYSgO14oz6CkbuZP5Su7gUYVUdoPAJ7gFUTqY3hAnqUCpY+dDycCKA52
iECPb5IbdTpJ4SiQBm394fiMknceg7+C+fsD4MK3yr5+cyai1RDgWxFHUgzSgbfH
BCKBLVtOFgh8Rc0Hrft7W7xaPpPVzZoT9ELYuFqsMAZKztlQAQMeoMWpGGSWTXD3
3JNxBQ9Yc62kLcx5UKhm4RUfOC/BFXo06sOEnfqGZkpD4s5a069AqeQIkvZYnlgu
ETq8nf4RJYkD4crXQ+y5leaEVtSWhw/ypIw6ox7I7wFmPI0/u539n0Ecp/9TkSpF
UUYOlMKIKk9zCTeZ+pmlo7PpGhWnxUi4AeUeQab3A5eUCZH/9RuEP/WfbKqwS/61
mMhvzfOodHWE0uMkrLTooT4YsUlt33RlcMjpiiiOLAEKkr0HmSBcrwGTKYLhQJi7
ne3gMC7iWLWNxU+ghwP8DaTENpNGAEWZxDwXKtqKCCfbz13GE4RhFLmBiQgZkI61
eqbk2Mj69v/V3/1sENx/PhcwZIW48WXnAdWnudEXOcyEFHxwZypyaXdSkQlSizIy
Qh6T882Wu/eTEiNc4ysRj9rxq+Dl3tsuWoSpbvWwbG27l0oAotds3mL0LNDVTiOe
ShQ73dje2gtKVruJbLQBhJdgMkXy6GnKwphmrsA1wyg2//bIoBtUnzGhM/Sk0JYg
RxPbKlM52K+byqxOo4MKX8bPhyINB9BD2pJDbHVvPI5zc9npPY+Cf/32ly97dNJK
LYvx0AMi06qLsb5nO59xVDBla+c+HMRUafoDG4QXnUEhEf3ZnRUZdBQT7NyZ/4at
y0MXxyxp8076UmQaLwMXhFckApgus8E4MByhIxYJUM73YikReqYKhG454xKiBjxU
MR0u44tLHiNLosdbymUSpovaTjqrtWt6hxyrMDFRz7iE8rcqQP5nRtRFh5LijOr/
wKkGQo1+pwd7eAS/DFFts1KVgsJ2n8494TNHmADLD8E7kQUzThUZOCxMPSWOkUf8
Kr68U3R+zeREQuHJzAkR84uddk2fUEuYUPyaReOh117n1zbGu/qguPgHeKoXoNGv
F/rgt8gTqJYKzv1jQkhtsMPYSYhArYUdSjN0oJx8Hn45CV/7weo7A/Wf8iiE83Er
A2TXjrjZewuVBw4yWKiDqhJbG58wq5oTIR41+tXi3TRaAa1O++869W10O6eanhp1
gDUVFTgiQi26J0b1N4c77GYqzsQE+beDKEZOBpkA4+GdzLHXGU1jnmOlNxrts+hT
YZbqpReLWjAE9rW/y8ENo2b7003AaDf0+i2cbtQ/yPl7xV0FaiBBr+FYOw83+fHF
mueL8Zf0MQ3J94pvlj/4ExI05ZaHLFrnGYYfxyQ+35Ev+9Zg1Edt1sRBisBixosd
gA5dGHjA/RyErfL6yswOMjc9xemNCCyVp4yBeuFAqZZD/RUzTx2IqRLHvn3b1kkd
vAoTsp1pe2QN3MkJ2siTVhTACiV9FUBGQDpyW2uxHE+05Xc3Vq1vGLg9PZ2jijDQ
N+o0LbE4AvhruaZjx2gC0W2Ceb4r45r3lK0kbeHKhIVauCMyrP/G/X+6FQHgXB8s
adseERnXc5Z692qEJ+QJdGuN8yB0gxF1LH3l49xe1kDJHCb+O+egyqMFNWGxur8W
GgipqbErLp5yJZ/hh4sm9T9A82QXHf76GyMAV0fEhAIek99cEHMCTuRnZrO8EvWd
ZkcNzgbKYWiG8s3zT4S1oJgTsnsHfAPnsQfx7jaHhWE8xasrLHrk2mewRF7LgvZe
38B8PgbHMcqSfMOrbSAMY2trgKaKw8tC5l5mJb85/Cn+nXwzhjwzvAgD3VjH0yTi
HQCX4t1TLqBKloKPOR9oYmyJje7Xt4VR/UDtY8IXZ1E2DpvyfcOPhnsu0E1GTfVO
R5SprGQ2p2shCqtv80OYtkOQ8xiRNplfvTU3N4qMvGrQ4UMYShxgP3yfTb8JFC+q
ltVhDQ7ccv1S3BIti/Xi/kct3vh+zIGMtgw9d4OlfvdsqjVXA15d1G0oHWl0it7Z
f5wkQ5/GOjUzS3ze3fXEGCRCq/QuqDmirSIbMHJh8q1SYwknz1yMMgZjtRzaQ1Cb
Iv8cbg4CRd1Lz4374rsCVN3cnGEny9TiCAW4dy0rSz05FmnKn5zvWxlOETupNipC
vares4vYDTtD+Msqiln6hcmiNeiiFbXywHI8D2NPdER3rPUmCuMJE+ah7IHnYTDQ
lJB3D30QxIoz3WZi7Y/L4QBRU51COdJqfZgSUVr06JR1ojC+qIJAj3a6pLIsqCV8
jHGtFieY6VXQaHBaW0pCkWuRuvCAUHyhMqnEGIk5NiC/QskhB+OyEIVVNzrHRrqp
pZaD5cvo6t0/EpbxywRRJ3LR/LOnwL32PaNVhmu6Uw+J2++wO0bQgJx7m0FA3WQf
Rwh8bhZsBWmvMSaI3UgpnS9PiaTfgtThNsK+2YDHuxqVAQkvBGXMwrJJq0m1uaBi
dPwIyjTXa9mbSVwJ42nwh3m3di66lI0V/Dj+jMqx2rzLtytMqdhfUvbq1phkWL+E
EcA/gNVyzoTJs+c6lSNsANiJ9olBwrkZb3IcNgDMyfmHZgyzE3PGR60NRBP8slfC
89ospXvW3b2xmZ/VAI/bRwCxWP1dTmsOeYwtVjuq5ClFae+USwsiCgU1+Tt0HKlI
Qm40m/QPZukJqOQx0sN1RmmJFPookk4bUpo3fkmJe3+aUW9liJgGdzlsbNQsgHO6
Zz28k/VMVMH1WABBExG3Jhzx75qsPBrrv2Gs5hduyM1GB2xeVe+LuBniKQXFwK/Q
grriSOFzjAa1cJ5yArMSA5P1XTmSDGERGH1tk3kPLCEslhu8CdO2rI/HehffUbJJ
7nBzyNJR8DuNH8QzJsEP659MCLouIFsEAURGR8nJ5jz6wXMABcleJv6Bg04Ax4Iz
HZz0fzxH10dFz2ov9efMJtHdCl49ECZvqZVnDz0eLnra9WU71RlJjwZKQx6XhKxg
UCR8zm6tnxKlmPK7it86j+yvp5KwQCFS0IuEbdeJvyHbM4xYheRYhs3ZpGmvmS1i
9HE3F2Ko7VXBfHdRmQuABgLBRgaUeLIjl7acqXiqztxn08Xe4fhPHToWtxzvU1lG
hIzPD5CgW7sRAekdf5S9d6GY33rIbUHT5g7m4M5iBuqEYbTBbGO7cUGDVnIhu3Sj
SP08xMb/TI0MexfxtdG0AiV814DqUOnE7EAYTHtHz5wY3swDkYZyV8OyxF8Fdgd2
axf2oUm+lyT8rJb8t+do04lKcp1NU6yfpB03czLZ8d9WIqnP3r/XU5kGNIl/WUbC
qIPQdyQqTn1ktBdN/CRK0j4x+cN7W/HmZ3IC0cjhdJ56me9PqRUbeY2ym/0nGcmF
CiGdPSHmlNQQ2gM+JxMigu0DRujrVnax5vjyCu6W6+dX8KA2P2+9Nxto2ZIecIgu
5L146IhBGTUnHdGAUimv/j4x4vLWXopMJo3cLCo7/YdU4tACmLaXOBBj2zUQytJ/
7ZSqM+Xsy/WTblpT+yVHIRw4xG6rY+UOH5hIzcztcnKn0ljkCqbhOgcfDNHRTjc7
e5qxIW9CAY2af1jw0L2l+xfcGb9DwQ8mDRGanbUWy/5V+GvH6mzscEsjhF5M2p08
UN1ftH7iaMQsLN0bsfuh8KqgvPK+/OOSqJ9X8VUTUWfKf5qB5yYd89+7APhWo9Le
unfmOk4qX27djP+xc34uS2G91Ewuel2J8eTJJKzFpjMzEbKnQw8aLaoBh2iQbrs5
pbeX3q3PDRW4k8bGwm5WFFxuJGouC80MzKNPQdng4F3wJSGFrN4F07yxxYGkFuZM
A2fxb6pPWSWYRsTxxHbnQnkynuTU2CnKmrhZ//CiM2RA8BCVqyGJe5HBE2i02aVy
BuyacxaA0/Iin7kFVQG2TfIa3/RqbfJB3N0Nk5xT2ps5K3rNUPmApWAgNEG3g334
idHs2pjmpqytQJPHjZGfzADYFM2i2Y5inWlpJ3mGIATQ2aTSsgXAqkCShbgplkOO
tvMtmsbQTkCGCf52/I8bn8hu9Y3Jr0auzvfw6c0oXZLsSsgiqL8xKaHDk6vSoT4g
vya3v7g8HxZkKoXxG7vcy2ij3xvfwhg95rjzCieXFVJV947HI2rwp74YgaRE6tJ4
FD3wy2wnfJO32IBtp2PYo8De1O35xlZQDNUvijOlDI4EQkJ1V1NQ68EJ/3TlGo8d
xVrJS7qKrc7DvyKPysogYaiP+zluHIJV5aVqfshL2DbPtlkwSKS0I8+okLKfty3n
kP2NMCtqLCCbiCXFtAyoAccATZUR2AiQjt4ufCtosAlPA4zN8gDRgqMY5hITrrme
hVbRlwa3LRXBAb38gxJuPBjsf0e6QR91aUl6RojDyYN0OeY9v4Qw9AFsYQdki0GI
8UhpT6Mmzt0MQSUqAt1YpPcMECQ3LyXSPnuZ90qvQMEilZnmoIDXryyJUqr6Op7L
d/S2Kf9a0gHK9m6jQN8XklZr5ikb7n3XDy3dgEbMHMdIOCl+as7fmxXIqnFcXiwL
NOsd71f3iG7QEbUhehsnMcd4ZYVLJsfjo5h/GYWfm9wTEp9nTCNWyVEXnKya52WN
YNKPIJY0lij7Htc0w2JEcQIxNiXfdWvnYGAOd0KK3gL+7aoZpQnD61+Gp1gP0hRE
kza/UFi3WgpTyQwmOw7gGR6Cm6d+VbB9QQ3U8SwZJWCVDGHwUKhtXFFPXtGyYVYX
aKtSwVbGlc6dIcDLYmLO1M+G80RQnZp6qEYHMPqicZsK1QMKQOWUElVcRWVzQsRw
kXaVrqDxO2rOfiqLWbTobzl79LKDoFbS2ubi5+OHkNswImgC/C9hAAhIgYz2cAnA
cwNZ6myfhSIGAGx9oECbxmEjnoNmqkqFhtqWh4M+ri5uBQ5KXhxDcw+4Zfy6QrxV
0TGSBWpY9tPFC6rf43Mt5dgR/E766DfDywEAPJ0W/5/fGvilsfogcxNVKze6wB8C
ikR2KsGpB66X6idN7d0engurbkcWrLVj3yYXOURDSqmzMKiv0TRWErUWd3T5WGde
whvpr5HQbmgQSF3tGm7TReg7929MLrH0I3hsevdIDrS9jvcV8byZklfQ1qCgEVdk
G1i98KOPXf27nbH0d9smfq1A73fx2pXQF4U9kgo1+glYZPrP9TG4LBDI9cCHLWfA
m05OuH5ZYSJ++lehlZLeKlbloktBwgcSagL2mlH7bO+wf2IwvcWKE9pkLd7NhRF2
tU5F0OKuEiFVbad+uocyfbMIavQ3cer61QX+hN5NDHR6XdHtWQiDUgq39SSb6MjP
uFauepM8J/iwwGSS/GL+RbuyeByt82oBQdM/zk1iLY1gCmKnhG9pOLgBWfRlOxRY
5VfCX5DnP8pCYKnvsxUKMWFVhLVMg+Gc4WNYvkxrHbLls6XydbPZ5H3l0aoBoS64
/kukZGdZuVTYeOhJjYXHAbOQVCP3T7B/8v0ICAdjQsAY4MnbAQ6/kAnYClxP6+Uc
cudg8cnsIrgnlT9Xs0AWKb5X6JINSINKFg/Ieks2kpAbs6b1XbOhC9Mmxv150f4V
eKnps7qxPRwP4+XY6m0DjN1VOMtAzTfG5eIS6vntIyBCyDWOLA6vJ1n9VQTxvwXg
pVkFsl+mfOCj38KlvhZ4vLyNFQir/aKhE+fsIPx9EAumJSUtGVyNCamZC3vRTkdI
dLlnnTepMkXfa4liKhIVRG42qG3d7PUEFfsKPpEQFp8mmUbyU0a1ZAwGqgnpa0Qq
hcpUGocKnVo9FfDPKqSrk2f5Jt+/DUOJINaOxwSGC/zFhQ1RuTdn/B4zSJDLRFBQ
br6I68DcP/EJFvr7zDVC9FdyEC8AhgXsx2W7ITJXERi3QMynsfYRKWjggLEit7iP
IMXkjOgfjPEBQ995sopoX4cUHdL6VMQKEGb83W+e22X6EhBJwzsmTeukAhxQecIA
Hk/KUrlYsGA1Ka/D+6BVHaok9mHkPqtzzNsv9UK+8qKubBMUc/rUJlI7xg3qgBzm
9Ad8pAkdnfH7Sn33m1IN6dqbH5oDvfcZtMZlXEpTFd4mmidyBVktBoWdjXhQn+nE
ImSLnwPuWX724GN77KzIWCorHznWS5+4GeAtqERrBHa4MYRptlZfjTgDMOLDlCSq
sWdTNHMBjipVvPtq4EGNgeabJEf/ceuN9sl62NNiegtdDO+8GHqhHYiA0RvzkV4p
j2yCsAhcmzC13NpaPD2rR1EO6YqEEX8pxA6wj4mt96FW0x1e0Ot4QUXFtpvu9UBP
rhv06agOxeMicM80qnfWWRLTrCfPc0Ix+4Hp/NoXSmg+t9oHNk3np3+Qk8fsIGxF
JGvyXMOvywDHpnx4a/PQzBSq/H4HoYvsiTEF203X9iIqqXmSiharZ7mRYnVGcr3a
aloMwuRn1hwKqN47k1OaOFK6WEv6EhwzRNz33zvBOqW2qwmR/g2DaSaTYcewbQr7
ZL8zYTLGSsUuSehVE/BgCKp+spH8PaoFtJ32hFAbsn3+W+A45RFUAPBkNOdl4d4P
lB5gQ2E+xqWFV3GVF2FXVz1NNNAjdleoe9inWld1atveyC5EXSqyy8nDfZhfWkZU
yq268UTYKUCDW4+RLyVM9lvkWENCYFB8RQiTRdAaB2j1NOnj5sXkMe/776iCgHYi
uCuOEIpxjA25h9Q61MMCpYkj1gKFdTI6A/N4WyA5TkbmGlH5qV2X4VwwSzX4iNjy
a5abS97y76tZVZFo1DqpN6c1diDEsB05woSh7V5zAitARGRI8CkiA3FkapWTmCpL
CgYR77z/AuDRv1URRb9DPHeZO5OYsaWL3XVZL2+XcLbVqXw93l5wlK5XbC2Cc6zn
i+uO/aXY1wsLZLFt2pKl0FwMYFGB8565TzxVHd7vHe8i0lwEQcCEKxC1gMCAj1/P
OuZliEmTH8eWE7aZ57DF065CxixynSeJPQnWeCBkekYkFFkFHpyGmOuwIZaFu9UK
joxZQhYzV7oXjP9afdNVU3mMooWsPB1ly12XfI4EJS9Un0krUSsqqXyJeeZy4kvi
65ytrNixpT4UZxAZT//NVchjbEc8Vm5BMcL4vGE3it/I/ZmIRgSEMhWg3TPSoHY7
RPa49CBZP8Ukba17Ops66tqXBmUezs47aTsY/Y/qF91vqstZKD2aacVoav/QL5TQ
kvvfP64KZJH2ZTMbdqOd7I+cY5RkDCWoUWKcP0pkaK/STSzRZnzrsDsDsa/Obvvu
YPBr5bEWYWsJvW93nlpQPQwRmPXv6xEWH+A4hTDaWqaPirZPJhTN3Yj2IMEOlxbx
sArnf546JbKmcdU7hMUlDZVsX3aZF6cgNJoPYxrLfaRNDOTYE9M6n1EhFBbak/Yj
VDZ7KOPPclHHxwmsTl092APwQnTPC5SmMQlgmY82r8+MegymB4+IbPsOCIRqx5Fi
xt31Vl01cnWP23Iuut/+5/zR99dQwOozj6zObt9wM3aBwETKsHyjxdxVSUytiIpN
ucxx3N0+9WC2PxmVOOmWK4mqf7xX+D20lslKbmhTc9PCgSQdWrrdKwsRPyka7PyY
Vf+zTJj/PKNzqUivtf0RgrQg2+DdsqhN7iNmaKqh13HzbEEXNGi/nVdmec3O8g2n
yLjmojgczKaBaxKgc6kJ+Rbs2TOXvqzTc/kxFxmV+FocEhmh3Qg54FXOsaDY/VnM
tiLy3/bvMV0PnCRrwgutfpCX6gWhgcyRwz3NmwPBMqoKvYa99eg/SvexrtH+5Sbh
wcfj7ILlX6Ryd9+1zHtByzy4jAF95//8/5UBUUZ1+t0fvzIyCiNOH3P8ZJxt59XK
ou3g6duSdTAAdDiAE4wCwuLblqSXg5U4tHGrINOWGVpvQH8Ah7m5xMHyyBOmylwO
KX30f9kR79O04aIp/4GwUIAIvH9slkFFJelj6TLdjZfnQq+lCXwpizEB6L7rR34t
klHVnvEpR1gtkTgl404Kozlf21d2/rAP1r2xV4udWdLBdhaQ75/6gWOIod1Bs8rG
eocoLaRfJSjzkTeAqeUDUBNbFtEz6vt8WqBkYFc2JzAKHDHckOZVGGsTs3dIxR2i
YSvmtp6KP6NTENiDKObb3VeyjmcNBFQ+C8Utm3Cf/VP2SSBG36Pf3iY4kmB1Y3n8
u1X0E9uOe81zindkngppi+AQMqRbciHnS+zzmfEZrFFYPobM1IfWf8prPkXMrS75
6qOXjyJd19yzbRX7ElDZ7LISBEFdNidxsedbgTe4hCuuybKOIrEB7bDgWd4neXjg
KJdX2SxuRIC0cDbA522sCvBuyYOIeAbEsDIS0hjO1fPqvJTgDRzRN6jU8SrZ6xut
fQeWLBZcocMneHAznJE3dyZnaFdb21r3BOKI6czcspuII1ow6CpkfYdNMyv6OtXU
lG0z2eEmCfrQ+iIVBxvEviDMWwwt7zCft8rziW/foWHvYNV7MP7TPTjcUUVcrxuf
2brouATVJ3UAaF2OubMk1mY9L0AHbblXp1KHK1hcq0213JgOT7WooHgxbLfD9SOu
F8kTjXc8d4hFjQcL2aJGQhWyeHGqZ1TvSE4xRtQJlX9ZpaWO0Ni8J6nwc9hM5IGG
jU6EWLzFKeFc/0ZEkhx6ts8ECww5NO4jCEFmNTs83SXkDZWnKa6XqbP3lU0WeHkb
d2t5vCzeb6/2jozQsHztdbQXUeW29Z6M/RJM9AhjkRDaY7pMiBsaIGa0y57eKsfM
KQQLovUqcNHN2uILPVj3SdNvcNMaUdXaA3MHJ4sUVMh++aWAmcx6rnPgww3gjdGA
utuBunuAX4OByiduQ83wHW8S1YMowi6SOrEI1Ln+K3QF428dZtSKQ7i8SejZx9Kn
B4J0LrPTSSk7qvvURsZri76Q4EClhrCTJ/VpzBWjBXmikWE0RDB4kaskgjRZPV4q
wqkgVjFGD8SQVCQNU/LHoaOI2k1ZHxCEYdwLC2ZD63CCZaO2vawaEYgoJx3W06KK
h9uD4dCUk6oORJj/EtPLCReHzOitBzy4omntrgf2kvjypVksEb5kaA02AFAHtYkJ
iJ1b0mcZ5BSg1Q+29a5bF+qTxJOYguzeS0yLfXBpOaMMQxrCkALMrvzh3Nq+Wfuj
9u1wtOLc8my72BI4Z7YR4zJn2nMrrlsXORz1czSkvACBKlVjDUbFqPEdyYuAQKl9
ccg6ofXrHQb7d0DzUahk4YgrDQSbBmIfWCSBbAMTDE+IX36PceN5C9QgWSqmj1tC
y7sYehLHH5EeI0Xdta2r+vU2EhI7RJ2LgBCiK10tYu04yjvuyzoZgtI6m233zM2G
L31A/STsVj6FjSjPU9eeZ0xLVLckxkwlkez4mQgenDgnLTNGHN/SjUE7kfifOY5O
LFYWyXV59GoBDl2rRq6x+7nPmUaXytiYO4UDqAS/lfyIG/jy081y70LDRJByhQ/y
d1MquwuRVsSNCSlYTOJaRvrLCmBx5HwlOfYWjY1PSQG7u6Pe6diFCtDSj07NDp24
DobEq2ti5OG4oylQuul7NMNBKLfOJ7oaS5Ac3XEr4torlnOoNIYXBar0m7+1H6Fo
+s5E9IYR6sKI4XR780O4fBqk6V9ZfODeq1jBP3KJbbRN4OHT0pGzmKs3q/uzVfkm
kwa0es3clSq+8xXizXiaHzWGbT2ZxbGP4I6iBw90mr4JXfyTkrC3R2uAc6f6usQa
m5UjzS5BRe0HSqeeen8g0Ouv5+VqPP5ZipAqB4OQMBbklUrm6QQWqlhoaCfBdaty
2N/M/prgnsygrJMm8rhXWHYDMHmPY4it1haP90sr98nHPaDRJAo3NL85ftzqXzRd
obW7DdcurSAxQeLvk0mTN2cQagt+aLvohm8dC3isNeP96s4mvh9Nf/t9jWuBFd9i
vwzLPlKgxtnVwTimS0JZhDudzm0xltgUDKJ9qdWyU0nPYD4nXIovtUrNoQ15c3dF
rXvH1nVu9mCBayvZdtjz4vbr5l5ypcjLvn/OloeBLygTMoJn/Cxu2FihDYWDNT6j
caQqHCfu6VsENuB9AFZufrNgaKape/ZSjEI/jgLtLbi6PPDdnOc/ot1svgzsSRTv
sPPq6WzwhhqsGC7dT0QqIewCZI4daDKtEpkQp+QJTW3z9OOXOTrR2clnYE/67H9m
C2zjxtSj8Z+2UmSHQhh8w68C3b0q9l1VO6OUT43ZDfbZ5EAHs490qgxo4Ioxit7F
ayuaxjdQIxVY5e4v4YR344Z7mZ+vNOoLJsgNIobFhr4gXGX0Km4hELE4IjQ8FNES
7KrQ+Ql2O60IeYiubxBZtABzgTJxZKVfyiUR+hmMSLL0SnrMN+inVuBqyL+MhzPK
juHXOhuuPYQLL/BQor+aTscZKARu3relqtccPLgeuMXqwltzeFgGsvfZI2fNfFQF
RT4tYHa2C4bopFFliwXvbJJUAT1hpnv/kEh1NThBBo2sbBbY6R/ZIPXrP1cLqUoP
r7JL3XQMVjmw1K/7k6glxzu6HkfU1j0IPEehJXHYWkXIgm2yjkCC5CtgBWBikFKq
LR4IYye20xLN6mgzuQXmNvX3LleUtAH3N11FjbFZjpEcHHXNciMpqr2JCSlqszw0
p1H5lfrdz1fELey4dScCvJQKwC13gfWhyZF66KZqZ2F8cetbHnV+Ytj88Adj3lnl
jYcyGOxMC+mH6BXP95/S6Wn/mUZV8uP2ZHfhykP0ZzJ7BWdN2wY3v0Cdj4FWihGs
LOkvup0aNxZvaeBhP7xn0AZsLdTQterb8q7C4oPNFDf7MxyQdfCdzAEHLHH1hny8
Hw+JUv6j7Wo0zvMO3nBOPiV25v8QZQJNCM9rQvjGB88bBVrRs2gwujs0MjJ6yGYL
AbxwWnxLNxc3Bxxv3VS94cFFmKb6Naw1vvXg39r6e/TgW+Z7kMyU2VpZ2YERkcvD
Op7Xpb9pnbj922xYZj/EZdd13But5ey72Klp58h6UPvSvzXzBQ95WcZ8pEmxYCuW
s8V4QPcayZiv6fBWGUWt/mUk0+RUE9WqJXDRuxXEFn4FT2sOV1Q72FpoS7rvdEXZ
0bYDldRZFTnQE9mkp9aiIAHzTMJX+yQYZXXKeSyt6chdRJWQELsZf81Q/zbf4NPX
2fl+0qJC4hR90DjyGZES7a2+kdBe9L+cSBKNLmppLyD0ths9qkq8+TaS1CPbOW68
pnS6G4Q51Nn8EJBaMRhlNtoTpQ+SmqUQUS+QtYp2ugRBr4XqBuNq5ULPEicOfwyX
ClTUTQrMPfQo9DGbChw/5SfKT6/BoyEyVhIpI+VnrR1JuK0I3GIweG4UyfiJM5Yb
8M3mVBJHjPw/78jLoY+CdjjWiUWbTSj6Qy9mxBwpOZncgaEVu755ojdlRNGW4gR/
5q7hh1BKrPisfTH7YQavO5D2uGfFmB7h3LgGN/gB5dVO07EvUuj3bAJdP6QHminX
4bEAlzzHIW/4rjmikrveQixVss9PYQoyjTn86GqcoOeDldnP/X7A4pMcMgu9UOL8
81ZFcqvrBVEeAWboqO9QH5ysOdaESA+CQltY7FyPjExuPzMRhFUBtvVyYqDS1n3k
ODhVA9RG+AWkGeNUgjEfH9SqmrdpZ9Ii/wJKxQ/ZpEmdIPkbEbOTbB8t/7ApVuHr
K279ZiHZi1SroK+1TtXofUTUqd98mwJuRhV1GNSPScr9YPn2lO0nRcLxA15Q5e/O
o0HjsV6WGejW43mGw/GlWbjS3S2vlW7yGNCc5rT3G55n7AHKCMAWlcJ4ZCYEH4pE
rW0rHBogsCDqX/B90WsXJ+Uh0OHGG5WnLhkg8Ja1daVHi1iQnEG7wQD8ZLgJPOtu
VMLZH1fU3uUBk78IU9uamf1OB539lUHTTdQSDhL9NqpavtmK4uLwGNfZIsQOocnm
5xm0YcxsZ65xHf9Xcc0aXoaI4hEMJSsAzON29yLkURSflPwYRxnlyMkeXpuwS4OL
OqgsoADljrUW+chnOHsWWLc37BHjmZWQr2eY+4D2BuqOb9NfHMx8Z5adV+IqcP/F
//DHjT7bXOcJUdkYZ5ES99feQDNUn9cvDRS3zgPRfkVKOOcJ6K51oudpM8JRrJuZ
Gpkq9VuztpnwKUqpMJvtF/+s7BX5XDF9RwVTJqha+633ESi9R2zPiC/6Z/ZgiCd2
qyRTlZeNirsl/ceVg8xOGqtCgTxhQQpbyy9zCdhkP42xYX9GVDAwwMPjMsXvS8z1
hv93SaGIB86eRR8SH1ySeKJoGwcdEmp9Izpv95+10vOOXmXgsocGCq9IQFPuvadU
Ioihx6ZbSfs9RPHshr1Hh5oRNNSSFvnlYar0R3wOtrovJ7w5YGTR5DKV+r6cV9Uq
nvAjMiqqQW4CdxYNXBFg5Fz4ch3pNk2fIDbbtnPd77M68i1EJA3g1P0N1R58r1x5
1RskVSX4hDNdzZRMz1qcCf69UMayAJptFCNvYepWeYARBrD9gCYdoDBldtbqZO3O
/AQC9Lp5AutAXAEv1sPe9dPGen4CdScVlMe5dgyZkd0EwKDMCHeFUNj4Dlr3LPiD
9kSqVA/wS4H1dg1nAkwt8byTfxoVoeJNflqg6PjbOzMFTJb2fJKSmCwVnTVW7dIk
PA3NoVD+pfJJED8YNcx1J2YK85bmnCgv1CcK8NSW048/2hvNXkk1JY5zskxVs48l
a1THr+oYnFXg2bBWo6wnJikt0jnklbFhJJi0D4xwt8Nh7lcVwkKJ2oNvGvHjH5nc
bthoj6WIX62qGbYwx+AOCVJ4vRa3ISz6AT57tf3SjjQ7s/Psz549EzapuxCHpyxM
5gsA362JV/yx/fF9v09EhTOuiSIcJ0OUHU6XCh25svol67lJx0Saup+nW0m5H1LH
M+zFR+70lEXQjZlfnCp2ez5aTDxWU0oSxUAa4eUzz6fR9d+ATTk2e0ms7dKfJ0A+
zLbDw8FcQW+I8GjD5iM5ubUtycawDoi4ot6Op5VJM128+XnXcpeirrir/dnYsbD6
srZEAxFQFEid96D+6YIWFiXzDzfYMg9Gq+14K3NqH7kBYQadrUBGUCod5jQxKtKR
qdqKeAi/mmb7Qqt7YKusKNZotHMpsuth6wkywKy1oDdMDH1/RJmbac2dgjIZkLuv
NKVmz+j1tE26MswImqWSn3eurAree+d/2Cc/5B6TKbxrjHKUGG/5JwLSYnPtbnk/
H17KDsT045GXiKs8zl2iaWkG5hTqLEXIlyxvY8upKUowjlW+mO7fySRjRpvrlrcT
zgmT9pkJI7N9rBpxezENBNcvVTgmGqKjzpzwJRBn7d1DFg+Zyfs1gr8ttjRH0CIL
GpB0Qfer/18EogCG/fBss0H5MsvM+xWjNDlOg7ZqjLX6ZBSv3KuevqLyXwGvUO35
PxSvVx0+uEhTBTQu/89LtlWFWfwnanuX5C/9tJ8eLMinuiFSry1mQYK6/acWPUKf
CpSCZb2bpXcm+LQCAAQIAeVUPp0PJ9RpCiFRi7cgm9vC3zWXSy6ZFYG9lJP5B47x
w4r6NZUyNPCF50hVuix44daBGmjK2V+A7X6QeFHQX7ilETiCG66XVwRf4iXnxi8a
KwtivCLbrGyplrbZTeeIOw2W213zn3/TOaJETWst99oEO4N8z/pItUa0F8OOVosm
/vMIhD2rS0a/V/4Sg9CIDVG5Lf+V8wEkjsfHwB3KbhwTcHZWll0jbkLUSVXldqV1
BfLWGiwYwsI6eqWLjp4sLxJzH9H3/LqeE2Qd45DpYb9+tMUdiUlkcCNxDLg/QyYS
tAkF9aQn1YOcSgkwaCKtxttD2UsEQyTgfQ/iplkYkGk3/qMy4D/qG8xWDASWN8Pi
Ul0sgibmSP01RZB9OMp53+KWty0VHoNZjdyYDbO8gIOO8fxwUuQC1i4V5E+g/3Yg
ZvHYBCwUNvjl7vw1d4TYXKZ/juu7XM7ADC92Tr+bQbWaflcvTaVFaqJxZnd4kWzX
OYDxa706+hWAt0It33jN9sdisCzRSNEOMz2Kibe6sgM+TrYFxwHVbzuvz7iZP2IJ
ERPTN/xHIxhH0hxtPQS3vuC7oxMxDh28BkGdr/i98fQEvb3zfPo9dFVTNlwjv5Z4
TgK9OC4g2GkHRioxRPWLzYO7H7PcL/RSqtmmMQhGU28KTwYAeUdn+KEQ1xXwbfcx
yKQfe4dTrExTzSrOwDXhDU+ot1u0JFxAlV4Ehdl0nemSg1EU168HyeFF6DBLs6rL
RQwipobfdx/a8n1OGpxpE57FsCExVm6JCtB8xTdzaElTkzAuLSMPRrcvBhnZjdMO
wkyHHo9frWkZ33yv9s8W3FxmKMebayK2hfAzQh6zzS1I714RtolrgH4yyX2ePLdn
gSnYPtBkfOQZjAS/KEJX00S/ovJQDtvDJRa4oYQ5dWeyUdcPhQQDY9W5Kdef/qco
hqUH2ESF7WFVs/oZ2qHq9nIt8SeUydBgtOLplH+mEx/hp1KcCSiifJZKOk9GpWkt
CgKOPo4shAXLOEdcYiBIEStG0rjWCuvvLPq7SlywV+zta3amyc+DL+126tVfX4nJ
WGwv79RpDuhbVOOIW1VJCUhWMtZBgEwNxjPC+ZPwHCemTlrafpB64cd35U0D4j3M
3ppje19XFPiJE0ElGBVpgCzxOa+pkm4jJ/L/63E04K8V+1Y0+ND7EFmTSQcFSmmN
KaGpO6cZGtpQToaJayAoVkYLek6tShUXKm1J7ArRLpL/LxtbGCwW9OWIx0FXvHXx
A6PnJcgxzsrTIPRE9Dd+oWUjmyvWLtuT0TfcB9CL+MVtse4PcgQXH9UZ2BEbGE9A
DhqqHfJcPZr1pTpr0v2MuSeeddUE9PP9NJr/xYi40jgkDZdyCHE4B5VF8i+Mgk2l
fXFW1o2G5hm5ZFcUYCmcG3fznrrf20GZmYgD0xdCT6WlkxBSH5BQhZb58h21Dr70
vOIA4KT6mTJO+HWIb3J+/qMby9eLj33iA/mNNzqrrMwdy11XM1PI4ZUL8G2KIUPF
XTH/suRLoMXl26JoEJ+MkJKE/0h5NnWhY/q8dbPmDygcZEMVK0wV292jMXT0DCum
7vBpzcms/1FznRxhtMHfNYIPS+RfxRa11AGd7Q1q8zu5OW4rL6dh1KIWzWvV1cHa
tBNTnAgDESxo5uHL7YudndSSxqFERLxiIaOREdwhWcb5kuAGxERl+eKtVMjLy418
g3UB5zbITvtQ5o6rbRD2En6hiPQGG7ijaW2KBI/1Hk3aCn8vcjvv8jQY2b5XxzsF
0Irjjs0AZquLexveeo4iBdTDgUvipaQ4fKqeJ+USmAFv6ibKbfEY1uiP5CvKGHqt
GqrHQEbQctF9TWKiaG8tS8xsgmy2D9Os20hIlE8P9ShqSVig50E1pJ5YzRXfM9bo
G4hoifHPHOueHo8SUFs007Fco5su+viPvmOU8Ulw+vIfO3Aq5GoelrO/Kafau8w5
1/ND0oCSDmFKMov0cMJT6ca2QKvWbjFzoECDUP1AbcwJmNAr++XE8M1ZmaDvfrrC
CEJF7H8DRY4YPldEvKwsKHFsluO8Qyqg6vrCfVboGSoeXv7n1pMX8JDD32KlSm+i
da4iGA9YALkKfiRRKvOibdFjkuLvcL4EicvN2K5Muapa8di1xv3GTNMMEPD8AvBd
XA8yduAi94WJKl/lx4rkqx8qwTEXmvauDgrDjpb/eIwv+l8tPc+vMW6MIewgkqsR
s1DcMgEtHV00pLm6N6U3Eo0m/U+mk6nolfv4PZErTnW+grkUpTQeCzemNdhE3IZe
82dyZU8gVxpqy64krLLbpkF8jt9TJvHU+bdo1oeHBgsww82i09jE89WIVSRxFISC
0ZosQchVx7ZgNx0CDYF72RVDwnqADrkk2gKcE/QMmo3lOUgYOHgYRvEwhCYRtLdF
EWERBzha5CSeDXW3cpUE63PTT5Njcojow7y27LbkxZ89E8px+vn/qPikyaq7hcpx
Ut2v2h0abf4k09m5gqRBKi7sXx91xxkl/O49rLg4D2b37pFAyJwBX7YUevafsQc1
/zUIUqzUQ+vpKAzHotp0Hh1ljoh6z7S2fcLo+DgiIt4Wh+ffWeoi1lnYsryuvyDa
dQjayx0LQWDVYTjkYcUyqegRlGGPF3p+va+tRbBqsQNFg9/QbEQZBADKXIhMrysM
doBKC5nfoR0n7BbqLUvmSkFIS745WQ3o+baZdJHdUY22eF50NPAUreygYzDvy68t
tvOT3Q1hlTgbxOgVsp30hMlsbLkrQJxirHouM9m0XOiRT1jQaxW/oanPV3W7QZzy
FavEjwShaY+A322gwTzbcByk7AbatiXIqEYozZBxahMX38DiiS0H/yDvQZ/XiAi4
sDICuQU3ZgIO1IEuqKYNF9vC1P6FKGHpEBfYUKMGOMi25vWX+lRAdqTo/QDKjU2l
gv3sXlW68/h+rJWLoQye5dFG/BU4iFwOHIr3O1vUf7Gzn7PA/Fk/kD8/XSkowWrZ
Jrx87KfojOD0nMllr9+VdqxGZwhudJwuUTw11jKKnM+2tXLtt59uqDYHwtk7ng2v
6YAJXUJO9M0GO9jhapakoHKSK2HCyZBxYeYa+0YCdwFgMhl7p7oX/FcHlKnv1ijY
hjybBjDoLfTrWfnkTqcWGqR39nBrtqp48bjt2Ou4WjSSdTyUQ0M+fOFa7xVoHm86
DgPYxDaW4hWrECeo0yB8lZZ7xP3/at7knguPrdnp+fGg4OdVeiNDoSO3JQ9BnnYq
J/V62/4PImkicJOMBiTPCNF1LCNnB4IRnzprjOzuwdtUuH3Tl0MHIy3doBEFoYCh
Wl+sr9K3OfufJibUit/sN57rU2OMsIgVT8HC5e8H3IT2PN5YsEoDY6VDUC27OFTy
2Y7vclpPa28Qi2bk9yxguC3OpJFpbVZrGm5VtamrAXJMGF9ORC+kVNT0nArfkcP/
pSMbiXj4GIgcsCIAjWPenBPNE9R25T9DmcXnKj1Oo/xymmcqcXcSB/TkjXl4QonE
J7YiFrexqQROWdSTZaOJL6T2E7e9lNeX/mthHiZPwhWLOmiBxCzUWZZSy270mqJ1
eLAwYPg9XRFm0K6KI5UbUSLP/cGqa9SfUE0P8KCzcxFv+SjzY0PAQPEfNL/2Kz86
LPNCYH4E8LJKGEgoplhyJA38wApERAZU7W8a7JKUymcNyVtnHLBmQwZq9Y38/pS/
pTNr4cL2OreYjV1cD1hoYxNB4RGv+vDHnXJRGPt5inm1A7PiYyn6E1Xya++cRTnz
izXFgRrO9WOtta84GXN7JuPol3p/Y0AsNB/Kv+NyKampKUgaaG8ciE4Cb6jzmr3o
ye7SUM9ke4kYbAu2yW0ZNUdWckx3TTzWTaQxxabWBHaTQ/p07HCQ0KW4Q4281DDh
ukrtQz9hLetdFupf6OFD3AcM0IAti15ZjgfNyTFchSjtjvEeFaRPEUgkozGmHokB
zfeMXUicWW9bLsQaHb2cWeWolFUqNF63sCN1MZimJ6YTcKIzbN/14Qizu10W8Zcy
HE7NTUi18yT3uv48aDsfgrB0twg1GXwzvonbGn6fpRxSjk6vnh0w3ThsGGUPlPEC
yy/bYC1n3d6EK1nxAo4/8tRx6DhMLDgnFGPelNYmQXHt66WFdeGplJFVv+xkNZmm
FckKNdhKMKpspiW/1ThmzNqSAYhWbukji4EFn/MyCZkfCLanB410cdDwiVgS0pb3
/ETqu6sWpN6yqPKDcQ6JrdQnpNrjv/LIZiq9/QKPWS0vA1jiEhSVNbILGiXou7Ap
75Mal+aJDMbSUad/WbZhdrU6Xn1aeR5Jifei5FelkBH4Hlsg8hzjS9ir05UAWI5q
c+BOISMpmtJnHO47xWZzPNIWmygvqXzGM4vRFpXX3FACdRGP9/1lz83jY9/+Xsli
DP4tMSnENELXssx0LbEj2o7B6augiIF/2Zz3BRaTEB1Tv9aKFsgXGPOy5aV06hrz
LmLN/jP6icl3d9yVv/NPeKwwQ/7cBKCm7kptHbTIYThvL3ypuFe9HcIMKDOHCS9n
TNtgLGN4r31EkmUeGR89sS+I63U2N4E3wCYPNat+Iv10xrU3QLbnsTQKzF/CnnDl
3YVkEmlbOUw/peoky2W9bRH3lgd/UcinG/GmHgrRs866eR5Tl0crnPC1LsbiiHod
4zmEFx9yG9TNQcxt6/QZ8/3KSmvQj9TFI/0hTcI6UkkrqcTElFeqpARyIMVshEGr
yKz1B0DecdST7d80F6ieiwXLoCGJGpJnkFPkpyTu7H1mWZkXkY3KPh7CpPqZdw8P
5gAJrEQmxbXsrhZpbTdXNW+E13hiIxTuGrFMz1Eg5PAM6bSgBRMa+2xogSI0qrLb
GfO99dF83suW9CoCSjBajSCUwVyknBxT0AFdXe4Aj5EMwZdYImS9DbPph5PbRvJ6
pP2kU5GukoyEsNN9QgHLr/FwI+cZXHrcOLeOJ50Gwtpr0qKSnIaO+4A7YUpgAqZI
PcT9KbpeISZshFl45UzsSSdUbCMc1p7LO7tsJpxO90z8wbR3ziLG3fvtDCacGoL5
4XcG6MaFy1ZeLGyA27X+h7LBHr6xq8Q6pR3nZFHsD3eaRcTgl/pBU04xORngIbuh
xbgU5QWlQz1dqdPLs6NnijgfYsA4oUDisX6aOrdZsyyEh6yDjtxofCAuOcFBdQq5
4iJf97NCOpd33/UensZVD/UsettDC/wpMF/fdYaI7bfMpUxbpl0HERIOG/J10eR1
yeg9S+is55g3+UihXGQyQDLb9syMIfh9KmJfeBd0D2NNbIKm/ewURZjuT9cv0tKf
bjQ3IytmHeWsZF/ajKGQnFN+3csnwOKKokYNpyssiIQ3LgsEFCJAbdZAeo/+O3Xh
DveKTamT+UA2t4HqfShBks3qFaMlPQkZiytgt1b5+JGL2ZWoMeyWORZmwtBNNNGF
7Fnd0L2vP0U6DZAawK9tZS0VvG/04oaL/MfRVCUfymoM/0poImp/N+YoBhT3HoKz
2+9KtnRj73ByX+P+Erjd+MIfo/r0bqZJriibTzEtnQ6Ji14Wi40iy6Re2+rdpE0b
8z52DBGkVmr7LnIbt7f5n5LY7x7QZG+/+KQei8UkR37CWnONnUmczliYDK9sTN3C
dPV73k74maBoaMVcg0RtmRUxjMo8c6gfuRpGLn8XDrx2X+oeU2nivdEMrpH+8k5m
QYzQSiEN6tSwEDMWPtIvCov4goDOjNxO9Px7bWpLVI0gHSMBJlT2MYkJ0BT6dJxp
ukAQvOeBT24DJSflxABJfnRbBFo1s3GZyTdwNxFl97tN5pgLRMrgB94eRGDzxTkj
0tGjl+2e5INwFpDAeQ5HP1tlgx5kqE2pqYPG8d/fdZMyldyRrvnd6QIEfn2uTCTP
D6d7anBIEPARhS5AVkWrkUbCem3r0Z7AeORvK5+5ike4I6rkFjQlT/J4eSgplEe1
pyl7zZUrjiPXtM7ddN8BWvSUnTtWI/RnKDtRCzUtcMTdWYp3xNRet6IT070F6fUu
sCFYchEP96TDC5D9mo9mzAs3gpRqyQcmKXBtiP4CmaKC6vTpl0tz0fr16XAGGp3m
e7p7U7eWbqiNuq7P3msHX/0+dirZqE86dqSr5+RMohXMPZNqupUQfRbVi+XtcDec
YEYBZGcHcFXQ/7iuna1jj5oXmaan3qR5Xu5kqCpnJ8SJi2a9VIyW1PTur/KlKNp7
n3JLhOo9zLTf6fo9hnloaS3i1MjYOzxO/gRDJ5O+cqx+93Uqqk1rfvURfnVL5ogl
CMagDJbcSLlVtPQrSzWFXuNn1KTyhAdND0HbC27mVkvkXQnFVI2BeBs0XPSl2TIt
u1HcUvzwZky5w/zI0D+fJyGpKFuIQ4MJCauURfBTj3fKziik38tvP6JgVwSOimOE
VRf8PxMksL97hF7DFQ/C9guFcgKSoMTIIDGNdm2Hi3S5SJgKXxhrjzLnoiybfK4U
s5jsx+vPTlBVijQEzT/KetEuxpbLHRnlgJu9q0iNBUYo4V02zL4Ocl/2xr6uxy3e
kvbJU/xDyIRB7WCOc1+7g7ln0SIcFKeCWlME5e6LvhFtFurMj3apkd8wljCodqoK
9COQgdsrLTY28p/PM/5F8U5+e2Atw2OyoRGkH9mF1jseHnXg1Mb8mBux0A6w36TG
LdQdwIrO7ixxYKPogfM7pWo9Vf6DelalDMvMlDfDXWJY4kY0KLuaklid7OegCdTl
ia5JMgwrg4rrwrZ6JbdUNxE2NzCEexbp6QFFnmF/Bsb4k9tb/DlC3fKiC2poaM2R
2wrkj0THK0lmv7aWn3LOCc1nO6y5I7qUKPpXkmMvOxHJkHupYmqqkGwg0KBJ5LJ0
ntBOkzUYAoZL1u5KiCrFEoTtEk5YhWfR4vuO5qYLQ7rCFDkssmOYs5wnPviTTjuE
mXop+KBhbgUxMq5ZctbzlLnSD1BxDghmYoY5OuXlPqw3NCnmoVDzkUZDQa8lnWcJ
WZYYRsyXt1fmgBPbXXcbwzLtpVLkuz4JD7Pmqu6rwJvgX31xbZ2nEIm/hJwDiuRO
q1EruGxP66bJdCJBrowGb/Kf4vWJ5TIo3uuiyihPojznTnA6nkkPxo92yymq7IW0
9kp2lPI2+6D4fQFlQWHCsqamT7cDzZBJlatk1q4ZbYohps5qKSOL6prZjcDiWbmK
ETFSBBC5Uh4SrRyZ2sn/qvLNFfTBytc2AjhI7VjIzlrmDQIknOGbFFDN7pAjSc/+
oo4ct26uSXJ0yOzWHPetkSEgmd6OjK/ViZxGajfEXyJYM3O6FtIochco8IiyCQjL
PGMVvVYmYD5Kcj0RRsU+tiw5meA7ZuJXBaH64AafH7BQdmfm+v/tKu+dGq10EHtQ
abyOCM1kcEc7ClFaB7GoiVVIhZLjI6Y744Avx4dGHfLRtA0KT6PhOAEphLjuR3w4
KYKprCOotQpk67qbnRh2+LWvueqxuuk763Rs3Oy6W4/xsXh75DpwZPLjKjLPM3wi
uzTblzIQkELeTgvat+3OVldXQdAfWGx+eBvzOhrtr0c44GNlbl/iXZ4yJpAPhZgJ
UldbAn4qm0UDOPjTZR36izgjLGdkruDavCbt5AI6I9NYsMnenDvNW2mUJ32VoPI7
thUpLJqeccDiwwLV7ELDjKduMa+I6Ygv7WRdUG/aKe0eD+ce4JWRDzCSExcwRmw7
0OuES4Inb4q92h0Ha935M+XQZgWOGDc40u73Wg1DIABx6g0M8APH41D7Fcv1n+RL
EBBmK/IOrKPglpt1E7EyPZs/15IUM8j7zl1N1NsbF/CPHHIjXYXPT6CcmoxYaDIu
pLm1neB36KZY0kRjHFLRry9KoO5Nj9vQoNR1Sbfx/2r2zf0J+yPfKq4NPF/JmvVb
vWd9KDpjp7KgF4rMY2Y+vW0FK+PQmtoacNlWgJhDxgZEawpAs6n69TrmE6uJ9jQC
kz5quuXjeHwyjC69bnCgp5jQmhgHXSWc2cbOBynkCRjJpKwFzmC3io7X22G9CtHi
XJtm8n/yLeVlFYrw5bSqTKC5EJmBqdNDwFDPPvCI5tO5+dHOYZDp1YP4Z4Q4v4nr
svEy2fsVmZK6yQjoOTTgBxV+HW0ysz6rvtl9rt7+XyNU+1k0tbziJ51R19eRlbG9
Sz8cYtaiXLWkZUuCcAiqxJUwVRoSjTBG9hJnLJBIz1m7i/88zHQHl4zdRSLaykBl
Eyb1x7Jas7C+5Iypo6qswQVLVPgr/NEdQsF/cdQkVX0L9Gs6WFZIV9csKcs7zpGo
K6yTojax0H+7IG1yyig/Eu2uOFEg/ixoluatfWSkPs9mE464xTcRlK9NASGiN98I
gkR16/0qHRGyUupY6lDJ+z/l3MXle80HaAIp0yZ/g6IH2vJF2Za/Nk/c0tn2AEmG
4fkfvPBdF9EEwIjni0qutXOF5vDn8D3axUr0hV/LNegLZcz2DNuKw+p7c+d8WM8O
3Qpjh3kWSr03uzYgajEquxd4RMO6JohiZqBoag654Cu0vdvCOOUmjrt0000P13EV
AgM9z+tgzO8P5ThLowUCaZ8K89iOonRlSmsT2BSZ0oRghTB0Poq4QBEZXfiiMeVi
HpuK71bVbVJHCnk/PjfUnPBMnlOQMB5fx3NJRV6y+PFExzQYraSlar40u0dkHw+B
buzhLqWSJKRo6cA5djzRJch7BoG3EOukAKaOzPS98vFjHBjkHhFU/bzrJ94Cq8OA
BBocW8/tv+BRdyEU18/WhUUqn2b2dTd2KC+jpEL1TZIgcq9zzOz5KgRqPZgTxtlt
XaVEUlpCLn818bP1Mqhj72AN9DG6nyB4EL1dUkXSR+UxOl9twaPLEiPIz9BJueBZ
+pRnn1kx/Thn0iy/iFvjFuZUlCiBTMnUH3BPTi4PFViW5MScgp+7GCjHbOMLV24F
IpSo/+gCqn5pCdAmi1U9WOuGz0SKXAJ9ls/i41i4NDZFI5dv+aIrtx7o4WUWCnSK
X1byDaN4ojwp1aRvwV/t1o4tBUvc26RJCKMsIKNAc0BX5FMeLDO9+emLfXqPYf30
3rkZHu6KfVTk+ty7CfuKb9yzAJexRa+C2IosoZPEgjfd2XrFnmnutyIJP32Ncqwy
mGmgBzGVtqcbLMh28FpN7AZcH6HYKGLLPNuqYA1IF2f9iDjvqSIuEauSlw5JyrI7
VIwRX3ZUv7tsTBf1HRdAX2lNO8tXjxl2XvUijajpAydds6R6pUQ8xPJyxdMQr85i
Fsfs96b2xxRpeNu2rNBfFyO/mnXkSP3QJW3ZD7leC0fvk3YJBgM4Q4VM32aBHkHt
l5cgAKicm/mvft8xaNjtxaSA7WMm7z7vCp9R6s7EhAC1q2jbRuwOEaq371WFbd+q
sQdUDCvolxW6ywLU6uIOJf6O2e/u/r9JNaZur+ZwTNGFPv/r5h56J7BgdzDLOZAL
jheZd3dohON0ae+e1qKLVG03NClrTlgwfeYZ7vMA/dEKuwrg9lJNZgxGBp56edQj
+vxOj5GVixghxSRTC2V2uhdFD++i6B2xrr/qsLQYAqV02eVqfzRmu+D1XRKhpBfh
q+76itrqO8i7ggvUzAfZavfnkkskY50xQq7S1KJnAavjG5FV7qJpBWDkiOWbZixI
i4jdhR6l89Qo6MRBJi2qgHP+UcGGXhTJD2Yb3ejAQakUwMqi0iSQl0Pj1R4GGvjp
zfnuPmqHSXJHQl6v15dHKfMnwA0frjDn8VXkGLpsWgX6utHTrh9VmrbUV+lCWWL4
r8+WTLfCyFUmJlC9FghnsgcoDxcSjXOnOJVHjAro89Mvj+vU3w7tNRjw7xauTUez
e43mzARMCF/OB3fVUhKKtpkISv3p5ZuM38ZJQGae/QyWE35IXif8CpltC4LDgtNJ
RQIxb5nKPtT1KsxaaAQyAfM9Rhs4TSFouozegME8Ly9JRX5gr/taG9wRWN6b0cXP
KU8qiTZ4YeeaIX0J3l9zvkBvbRZvKAdJq5ZPdE7S58GCdD8v4eSpU3FNu+g3kSBH
PagBvDQA7l5M5qY+I1Wxn6TDeZrFSytqncewcK37Hy6wqNsp3MHJSPJsg9egCpMD
uxMcqdPTxG0+VdsialTtfz01q6xl5QrUcYsLMc1/iDhO7LUtZdncW7/3y8o0MOy8
2DpRBGGAb93pOcfuoYh5hnMWwcoDLZLvAb5ItREojb+ujbL/gsyaMYfKcQa+trSS
mLeC1s3K5opBxylIfPXGSdFjR4VbY1tMhEcHm167/8Nf9Dds1y0qI4tBAcdrY5Yf
Pi0h0BLRK+w3xFfNVLl0UHdNl05D35WBA0C4Sl5HwM9aL7b3oico0orSFfBqSmQi
3n9uasIjdCVN56YqAj00O5P0PEAdHamSTYTjbWiiCh0JXxpN7/wSp20HHVivk+vj
r0/+Fq2YWOfJypughGw0W0wBIQdLlQFzwDI1v0LOO3KyL7AitQhH8HFGgEuhPNZX
kQYhkvJlojm7QKI+8ACQsoTikyj2UClXc0kpLZIW7YpOvUjMFvdEM3H5SEGb6k8H
HusiNvUll+cbTGnyTal0+dGL8qwVhwKPHeW73yoy1O3ja9Wjx5clMEcoM3bjh+C7
i3GXhCOk0xkUOMgupRFnGY/rj0+1dUSVdFy+iTRZfCMkKtZNmm0hIKL3DVIRlRZV
hl5pYIrNDSn9bNRim+wASKMzFmasb3ypveVGghIznt6YMBkjJiGx0go54vi0M7LE
15TwSgePWNEoopGKXXnPz/kssJiiqSuwbawHieeLJ60hqt7JYcouf7+sVe0sRAGl
2nkMVMQe83vOQollHBPPtvQAFmq/aBZWMTdcaie1OV7xFzLxZULZQ5OUuIG1t07z
AsdactrcT+7tEprL8ptBiCUH+PvyZ3R+zM+qdiNhe+LG2s88T0IhogrAX8ztW0/g
LoWqpXkJ9qBIv1pAjIDuICOLlwikIkBEmHYe3lwiU4dGmkQ6CduP5Vrin58HUPmA
pzka9vwRD8kD3s2jkWFJ138yjBiUCvs8kYcYsu4cqn7Lhuw6kF3uOkIZMGxp20Vw
YOVo1BZBOGwxzqSGSqx69p6PU2ji+0+eR77AGKJXvsDAQulQr8IlY4wvx9mMvm5p
DNuMuiUiGeLCbp5B8dYf7oHykhtvJXqtlhRIL/AEHaZUvjrofLQVHEdNYNeMYvqh
JGRqZTl2gq+3k1EIhPjotsQtjWYAlM/M+m/NNaYLUbrcqXq1D+BQp//ugCM1alPd
GiqRyIPuzXz7Tp16mmxrit3vNCKklAnlU30W9NEeU7ZoQO4ih3imvCbf2mKrOqVa
5ouql6qKMc9MKEcSMuL2BLTIORj2QuXfSgPcWpNJgpfJjtIxG5ptiruBOEnALuzr
Sxqz6eTH5Ku7Ty4mbIUdwq8QOtRqLYt4kCihtrPn6+pX5lnvkbWSv0hiCZeaZoL6
xcmnbKfzcFE8wvCFKSW3Zcy9aqObOr8qB1GxoaaMxp3yVjFjaulOdRYsMT0JhxcI
x3egHtabbJD/hoRt0lP97f1tURtOX0gp/aK27IDTwFpuu8HHbuX2n89/2Flt/dUg
j/4jdYv3r4h5tvTHz9Adcbu8NnenKYH3vb0rVQ1NgL68Mw7MJPgEF3SYbKYQwByU
1q7y9Wm0xMLlBcv7GkD6WymyWojZ7LHIXEChRLR5xAR+kZgp0eMY6EtmHo7A/l8B
g/I3Oe6J0nVWHaS8jq7/V5iSOcCT8ZBq8dx6wO+w0PttdEpzSUC+7qznFN2TrOZE
ENDlUawJfhlUtAgVkNiw+LKogvPr4Q5oHJ9McK791ZiqwGaqA/HUT0LENfzaMKYI
9siZ5mNN4Ein0KYEoEqF/in6Twel3NR+YoAmx/95HYI857VxMzlgF9/ZMx84VwFL
flpugPUPiTQ4hIHDuhygGR4ChqGdx6fzoRGiTFitgUYZiVP0X81Pe32vnsO+an6u
EB6CvZsg3QjxbDHMAfhZvidGSboYYYj0plitQcn17Kt5i/YGUt9fzFreux+NS6NR
fhwk84c19Rvq6ViA3hz373GBf3fg2mqfV7yh2/1FIUYRtDzp9Kwn82yTt5xRYlgN
cfjYh6yaADf/G1ILu+vqcx2KiVEIJlJaTa1JLv1s60+DxzkwJTnzU3AOmjMAbTmo
9XXaS2zHuXqo0ZPVC+/OrAJA2FuDxcy81UdYh6cxsIt894OPXlNvGwMereM4fBGL
C+TjHQwJh9sJJgIvaLTtby1AdhQwcpKRAPMaL3u6YtBuot4c/gMxomm/CEhJ3BdG
XRPJ9Ff0+ct0VTupXSd4KVbr4EjIwrtmbCwatVkrkfZtZKkLZBT6xqPB9ZV0PoA2
pUgJ5FO2HwI0k0YLjnGv3LElim6Y9E2iW+hQOCY+tbFPgv4KCnKpyPWj2TmO56eK
Rwb2SEE1WsbwRb/ah1n57rafYHB9UBEHKZXMeC4/PIKDVCa8k5KCZBYrR72libHw
YoyqLy50w/4O7tbtYgM/8jlzqova5NI2p6K3/i2oaTC1aBos6+BgJ/rcKEbmmPxL
4Vys1nxcc88Xoz50H4Gr40lMWI39UirrNiLVre1r61J7/9eNDLnsW/JuU41nQwdk
1kS3fLLF424hxmJ/JmGNZD1e9ofAa6qRHXEKdsr3xM0Y6IF0Bi3+8jtjRDceeiAD
IckIz7Hbj7mEEB1Wg9aoavlqmKTkhrn0Pq1xLj05HTSoBD19u/tn3ZEvIyeLvN7S
MyNCPwQbMO4fsw7AwczEbpjZc5L0Km1IOOaEnpTm/NqMpAikdYEDwpQJkdDyoJaK
MI8Zff/IQV78vYzyUDfGM4lmSp440AfmdxQhwA9xbyL5nrExik2KYeYKs3yZkNjJ
WsiSK7fzg9JLvQw3zhpDVhSVUKS6btnxm4H+6BhHhxmzQITDUX4827/GJAnRyqm3
A/5UbhUMmX1K8EGgqiw14ph5VNeYRGGmC/V8bAbclUh9GqVDpT4AGe+9uOdY+kC8
ANvEg6OGkNOfaz46GN7WFm6LhBAzjq75xUJB+G0jBkeWTdaZTmZXZcAUhuElOuUn
tM9uQuk0OJMOXpt6R3qSTrtol4kEVecydF6QXOoE9gjqmMf6B6Q46jMlc2afOgwQ
enbWP/pHhFmcgSQ/0WA793MJ9MKrLSXiWNgNT4r5sLkGB/OuIDJkY071vjAtJCSq
wXq6Bq0axkz7xt/FfH8W6KaR/PrJ8MZBXeMRI7vGjXzxrdamG/8QnUqjFyVTk9ZH
NPyjs/yXuaE0msbgRDZ2f8KEM4hF9TJyEuA8pGnzHQq97oMNoD+tMvO6dFNQD+Vx
9oh4ExQfE5mYBPVKKtCIDTTxLHRYpRy3mki2W8E+5x1/Cv7G3M8QO4TGX7rxSI/H
6jg7Housl2JKbU/JJmARanY+8NjUxagz6r7cB//IoMmNPdt0h/09WuINx8TXS0NN
07NZKmN9xozTn+GD5qskU8Iic1/cSJYIqykGhcvTTHScud9EV23iJ4VewVspV0WQ
5nneCa9/3VjwfTzjzYLh+01wiIbUsxFTwL3I3d5O5CDsJ6V89YY2EBVSE5soPPPE
JFMdKDzFBygszyj8+NMzH69AAIRYwRYK/I2MmmIsOAb9230fS2wNVHi4jQz4uxbw
lXV4zwDyKkE2M8Yn9m3kVM04LnfFY2NriuXzj0kRe7gQYQ8yVfrGf+YfnFmYKNHr
DeXXFpeDJF6h9hRVU6BUH7hvCsNi2IAISDen1O5HBCiGQASGrJsBiMB7+hca92sE
kLEiwhxs4bLOffZOoH9zAU57lp+N3qzRb/yDte4kZne33TlWpuD9miDXUfMgaT6J
xlLdIplS6kILXjN71pboKHXJgcj4KIWEzgb+RqP2MHx76fanJTnKk0urLSqqDD8h
lRr20e0JcsFtYnjuypfFi/Gv++ivm4e0ADeHto94qtfxWwSxviRRcSqgMVzHSTDd
EF+b6y6A9CxVM+j4UGG5oQYq6WSwVKckCrtu9ZCMbABSE3JWeoH9YXxPIHI5HGl3
BPVttusXAfhbknP26YM0yxuJEXy8HYJtwME1NEN9RlAhCvlvXSZd0m7mVgXX5kjT
rNGD+ElqfrsgNEDG0K407U8XSDV9yHSPDu4V+8ina+U4kENqa/Eqkzs/wy/TXlJs
49cCfP3QF4i89XaUgmjG55bBesCMB0g9KbcnA1Ho12KBhx7yIubKszziOEONR63T
ipcSZeRlNx7GubA2YBLhjqP+RuFrhhPOq5U59EcUAvShQMyLlOP/KnSQ+aGZNduD
fuWLmaj5ZRsb+aixRHpjJUHlWKSarWZZvPIMmjDJWrYDEcg2IkPB2h+T0tfdZ045
DzGe5kZrKMFtmiCBvq4M1YCeG1dNcGKHMIqE6de/LWFky9Qx4jVz8pizHodvwceZ
yNRU51teI1hDmjL3C4imp1ZPiA5K75JRCdmnidhkomw2cgh0ChVtpmLTnODticGF
5PLakfmCok7n8WTHqRxLivAZJMxSzt5tQYZfHqvYATtqY/5BPXPdGHXARy1nECdA
rfK+REgm8wE5JjP2Ppp4m6NFnuJOwmefEcMck1FyxLsue9ETwm0XOUag8TgxOm62
PmRI+JNmAgneqJhOoZ6jaEG3XNjeRbIg3dlF427i5R1umbybIZTgIGWKL5uJvkGS
xKHwD9cjkhEsllfWQFEQTZq6QgT6pkkn4NaaMAlj2UeQTvOg+T60t82EytTdbMx0
6PQgU07EVqk9eShUv656mvinyWX7HTGsPAtbYAE84u3oPQvv9VF0C6CpidfqFsQW
9n+7e1hJiXj2gC3lB1RlWhOpG/OYYjl4aR4Y98cxRQpsuLcCxxQYepTMxuTI/hnI
QNxdl3l3oOeJeCwUdp7VKtcG8FoOrD8ORt+tRzj26jCMPU4pbyaFM0ZrM4IGIzF1
uQmvJkP7PwsejqbfeXbUTAECvVJefT6lajC2DX0bH08J7sQg2mF/NSMbQrpOz19S
/0ttT6UvBz0tchdXmlKAogcAMBfUx2yC/PukE91kfyS0mIH907sNSiKwMAf7ySYt
3pjAFZCiVoMGEm0C7cDhyNkZw1Hh3VTBlMYsUnfng0BvYOP9glFkzRtH1pF7O2pE
jYd/0mR3G6FYtj6TPlVrE92KIjxCEUkUSVk/CUGvjTNk0SrSLmstHt92075ZYg4q
l1tZdqN1KdNdQUxfVvceRjtOaY0AgGufCCcWiIOWKDA9FWp3mue5wsC8h1czXJaa
yecqqOkEpgEPnZaQ8VHHjaHX6DSTUjKIF6lX9uZTGjf2CX5O+OhD4ntmxf37QgKC
4jAOM6g9i8fYq1WO++Dasu28TbSAQUdJDp+mY68LvmPG6sWsD6gnSETfaUQ1jZuo
9TrGlBOkFBdTQwvBhiBMelZzJ0Zb3L0Hl+bCsCjwRDn1LTvCIZ9AqyJ1cKNs3dFg
KtVyMuxFjq2w2lPprzV/t2ccyS9r86OHkyS/PDvrfpUPpiCHNu3ChhqrXg2gHES7
3QQ6iYnHgH4cYdZexe6V+x8UVvwbgYFxtWuiZEVMPi/NPE1UBCgW1W2j5A0EtF+Y
kK04MOMIYsiLtcHrL3tDnUlRkr1uW1Eywq3m9b+FYxjw0O/C6riS/5tYrRMlsYKR
H4xOj3iObjAGYjmgvO0pExbvKbUbp+GDc4gMgYSQVNSZsBUWHvCGpTxDkyFJYrKQ
xv0/6usdT3c5RX0fohP89stiKVQs2lybZi5RTA0MtdWUea+xOIneKQ8fEhAK+TSK
xHWeP3XUEs3THzpg+4tri0EoHtgJimtSKTMIiiQQ8TZQHvjjynMfdskNCdoJOUlK
8hkA8gihBXoYGnZLK7ZE1QQhFMuZLqfDnDRTvCNoxLTv0gLPjH4DBVxOciGU0b/1
D0J24ggT8uxFCtzhTrstgGJW5CxxJCoNwi5cpjluhtGPb6uVU8eWG99xwYQ0jkO8
lhdY8+T3GCTP9zUzpmWTqXGNI3frUQUJBo50rCUQezoJi3jxFG1a+LTe62JOvtbT
2rV+8ZxjtqrgC1BzZa8x9Y2m9GoYa+guk5R/GhgYaGX6uRCyN/lAZCyvXQEkgPij
UniPyu+U/9xvOr9xT39Ix1K3DsZ4uN658m5lP2DOkErKzej+WP8Yav8Ff4FTAkgL
KfPCz/4/dL9sTxx74pUYTn5GQ+zlE1uszWbFJff/4olzaNmDXCQBBAnLRssSaC4q
Yir5XZadwrIoyEwAFLDC44VP3MVh4CMCEfqsVdOsV8DFNs3NfNG+frGMnJXOHsUp
4otvhHAtBKjiF7AtauGi9e/hqfa1zR6QaOUZsU2HBf/udpsHRwBlbrK/s1FBQoUw
nsoRotdFvmsQmwAV4MMtDUu4mG+T3J56QUIi5pVJGovLWnlLS2FTmWlEhjMftvFi
JP1xFurs2DQvVJvqBwle5O3URlLDffjwSwwioIayy3s6OaVVQ2qBLHJrmuFCyTcB
T4EojDLrQTaDfTY+L3cCVDz4xnxSfApZipdQoQR1GaSMyrXtk2DHUmYSXlZWDBya
74goReZ/4uzTCewjFn0eyOlnjbX59nhnnWTMHowhwCA6v1KtjgQ4JzQyFMo5IhDR
SDcD9db/i0RNkTcsC4sA9bTVbcEFekj6JCiK942tj9s6c1RWsacwlvFzqcaR2F9x
xhXkCGs101yt8CaDCSS6legdzkoM5NMVuza2/ExgjPnHTMdW2Ep5OUEg6z7w/UXT
67p0OgDXeh3rBnjWB4b5gDUIsk/l9kwbuemSVW9y9p+46VcLAeF6b7j3uzkWJhSn
o77/gxsk5cHnyUU1QLcmZhYrP956ioKkzICoNJhrdFfKej4XXK2oI8LXjJ4UEsu5
NaTsXae+IW/QGsVXcR1JWpDDVGSsQM5buqwqhGmtkbR4NEONsUR67gpng958y73J
LxPxIyzuwtHY+W8+fBo2rgidCLRDHDMGz0oG8YL91iBWuLmqMbri8diBbjjjNPbc
PXyqL43gAYayHnaGvIYeaybZgVXYNeswpEetLFcPg4uZy0HGBq+pmbZAjAwYNz4A
0OWypPQab1MKeD15uGv+MVuBFxJKEce9DmN5ppDIhD0+PauIPVK4XpEX502xMlNo
mVYY8lghgb+67jyPUcTUrRNeB+vePbhSi3g5LfjwA+4+pEX7UhX2fKZDmjdBeWJl
Nb81aQVGHOsEdxJM1j71qX1gfGpPugb4scWoHUVfMV+HTCbJ5Rc/0i5ovOBXgL3S
mJlO6CW2b3eKTses2caf4rkV4dB8XQuxFWitYFCX3U+RuvlNVPPn2ri0lCATWSec
7eUFPZRYqTCYY9v8hhLQUktrsON0Q3y4je69wx/RpOHAf61sBtVKzTBxCUuO1vOL
iPqUEWn8L2ZN/+CjNg317Qrbr0mMGLmPcefHDLfpn3eaWjK38P88qXMISklKnDvK
JYXMjX0Cp2JUaS92odRJh2jVke181QFwcpS3Ne7d4/uvTSknghr+bGoEtA9GQxq/
nwkqRQ9ArzBzCvz9ki3ZcilXZAa60BGpIiU2p5khk8aGMKjJB57TPrgrFyqUkKvQ
THOIW3sOPYuqLGduiJNpL3YeBa/eVb93I58IRpIxnf71wLVFJGweZzDg9uOtMWuU
a4sba5icJaenXplfCVOXxwk/tFx53rM/l6VeuDVu2HFGwQWegbDEk/41PhpWqW8G
2tTSskxWgRjUPo+1MwjAbf5EXrsz5BfpeQIlVPccvSARthnNNz+WnvoM7Kculi9A
fgMCQkDU31VrDOIasZHvq1zhRvRDInn7pN58zrUqJ/e9JwYhW1o5OlpyH/lD3DHy
DkL760aOofDFePiVdhKnng8lMsqc6a227nUdSr5E//U+F97H8MxV65wExF4/qwOF
IL63u0SCySv7oLjm/kqfNao2SzxCr9pqxm46cAcC0BqTcXuRw9T58MhWmw5CKOyy
uQNbBPjZZ0AOnkIgfyT/Mq8c9Hetz8xrw7ebrEbr6Q7QDRpfiJVfD3xSL8DUjEAg
gvi+t81qX/r8GwxOp7nYGF1AmoCCU0Pm9TVjvchSwckK7rm++F7Hsyac32jLKjuI
1rUUBGkCeEAdiZFmN6GGI3j5dSUIPMXUwva8fPaNwRuC7Q3hu9v+NB2FHHXoxPXW
8q7HcTzzZbun2Yt2esdLGLdytk0d5dT5RSRcv2QsIVGO8/tTVgYkJ9gFyLLaWSRf
Ooi3F4CqAQitwoY9T/tHF0mKQ7CrDhhR2St0xD05wklEPEScLLE05jW69VJp4qr4
6fEYfmFi8DHT0g2WBjm9+TmjXWfH2vLVBzWS5hiXA4S+dEkT7WYbDqSVZ7tu6qqC
rlsel1rcmKq3/phMSMxS6UW1s+C9cre1mVwHvOS30zLHoycrcfTkcn+k86yvJ0kl
N070iFiUfm1zi7ZWsgQmH+KsnajMyQmTM93ztOyqQG4Z0MurKLnynKJ9YsWddFP6
/FP66CPNMVOBEClxGjGibxo7/NZhqDLHwut60o5RcIygg6uryZhMAvKlo/jni52y
Tt3DBNY9w5t7zyIZHZ6uXHhBOkKV5iKHn3IJ9dp9byK2rU1WwXDgBKK8E3zXlKcw
rn3P+dPrrrNq8WJkSVdXuWhzs2SD/tB9uN8VvnIoCUxoQLaj7FZ+vIuWQM3hsILs
mzPt3bcWdj3RSmKzkFZrhA+6ZE9ra++t4KQuDEJMRvSWIS+UywG64G3yudOT+TLQ
Kk7AR+13JPaw5MxFTWCa1nS2OiQHN+w9rRL26zPIaEcptTjRXfeRlA4wrNTqOusp
caS2Xa9Qis648rCbfs1swUYtPQqAdelYmVOZtpZZxT5hTTIaIYPNX4SkPN3uIklX
P0fn3njK3mQjOIXmUxGMczvnqynus/e49/59w75e0OnOc1AtUdC4SvHP4G3Uotlh
dPh+xxGq6HMkqUcFUtndwXHp13rl2tXPXCN1AnmUViEshX9OUHbIkpOElzSOHbyJ
qftMSJzAoc1uauyh8slnl+d+UrpBSe1rWfoefJokSsByyfkY9Yb39PRePxuXb1sV
1w15I4uJNdGrP3Q5cRc2a1eeebkoxpOcGrbyKOaFWUzt0MHLIENIOl7bY2w3CzL0
ZCSpViBywqVU9kpxtk3VUZeSDu/uXo1zMEWDwdUAYSKIVoJVzl7AMJFfKa9TSLN2
KF/RoApJ5X0rIZWgkFnASDn2vhNy1KSvR5neXjD+Df9yV8TSjWVtwhcoAF27XxGY
a/Yyiih85Ptiwa2oSVvgvKo2OiZ1bHXUIQd2nmYrErMViHQ8NG43vNSk3YQTkWZC
pP4u1b/OkPDC0IpCJ6BAOCDI3HRFOycFlggJYF28JaaAEH+Lvj95avxCOb/82Nmk
UCuJp3QENyQg0tg7BaqI8E59atcMMix9S/zLGZ0eegKtCugGXI2eUzQ6n4j0oIuP
qZJjt38Wg4b+WlwNInQtS+Srz6sjN3ywcsVx1TwzupMWhcOnIIVlTF42LHf9PwkT
FqiifhqhPzUzhz5oQ0hBisisvFFSQsoYksDW3UWrObdMyYumLA1eYkWD+xcQNR5I
R3eNxk/wfoJSHQ/dnWyEg8fi18wvOTtwDNXACHEpahgcSGXp026jlk3OBWS0O2tT
RBox3eL1LffG0Yo5S6NKxY21if3pgWDBG6Pf/a45Obwi+r57K3DNtZkA4fsSXH5a
e9GwZslQ5S1ciHmis/PO9X9VVWRJVV3N/w36XdF0NsX8Z+TB9K9XsDKvrPsaM577
hdyErmCkKRsuqcdk5vtSnadvPSBd3b8IPA35bj+YTUkzRl6ohnbNuhiW8cHK5Mq3
UXObWcpqZKwFOBy1F6tJ6SoVojDyDKpKNOo5R/4vknen+jZ/cKyrpa0vO84ZNP/n
AB9DgCvna0eeP5rlpo4EuOQbQ1ywSThYCCbQKKIlSRbQowr8Q2mtWfLK1UwO9C6t
XnUHz63SngMQgHDgqL2qXqCZkpLXoe9Yo4BzsxgFjFyMGLGDVlLca6NqHbuL7g2d
Ch7yrngnfC9EsIm5Azyd3RB819CoIkPUOYOtiO5RUj7OxT7YT10vBU8Zx1QIy1J3
gZa415RredhNEf0T3LYzkzQpl1hCfx6V3aimGLg/m1VSmyaHgVb5hyA8/Ykji0R4
pUyWCb+JY8ka4tUixyA4SdduFBJ33A6u2F2Yh1pmTcDu8yO6sjTKxMY7+AARHPEG
xBOOgzbDMHPmjfzITw3ZwpZ9R2p+A1sg6wibx5D81xoqj62KIxTjyh6VGqAlySWM
mljKwMd66mMWEms1JFMJo0K0gbcssticubE4MOVXYG5BazzeZlKX8hKno1K11pJj
muF7wW0+Z/1LO65vk0vAVPDwnvlWG+8ZnwPcYN+1DFkzt+6m3DABtAhPS2GUkwW2
mfTaBIFkgUuECzntdEl+dKdHbQhJ6+i7l6Az++oaDrRfyIFZp9EF1KCdsmCwJAJh
tItpfyRcA0PKRYvyqJST9vvLnO6V78u9cbUVEDCNOalswQRU08LwIKxpDmELVF4C
0DENGLoRVehsOY12pUU7OCbG9iZQPIvq6YDo7NFqP9ssg4Vfg+7VrJPsBOVWeokc
yrm/FUjiPMVFWwuFwQe/bUOkrbasFgEW9LkbR3kabEVjauNRbxw3wk9Qdzo6qi6M
3iA+Rp+r/RKjm0+vopQFSFPeU9iBNPZ17a5rBFFCbtc9Xy7MnMw5DAAmLsf8xSdd
e0cq5PCVDE0DHGSvD9p3hTSSWxR9tZECv+tcfGh5TCwVKR8cBZpWsR4z9uFQGnZc
k8o+xPJOeXj1nuYKqHBTe6VhCirUjE2qjRyEyKFHoat1WUg6aP5WRis2n2/kmrF4
nUma9QSjUadJv9qUDEpj7cfVPZhEZoRbV/0oUxjxx6Dsr9EM2Jgv2URxk9ljLXfR
dR0t28gS+jkr/PGNB4FqtC9GRvX9pBndvjDEtQqO2Iyk2MeW2FdClXzGkViRPCXA
IwvjX4lmSMJsH2jLE2ARgUEP8B4HtBQaZttDu7iD1QtdgLlkg9sYfoS0eJzLWdoi
tjaBXni5L1OfT/2RMQ2bl7Qjt9BqCu/wgZdyFOhTR0SUevqXPopeflzpm3oPQO1j
qDk2kK6eUxBv751fmvFVQjg8p8hN4kBHA0KNgzAaFFrQ7s63Gx/CRh3qSN42oBrC
cBLt+HfjF7zF/EfywSNT+c7/RvD6mvgidHF0/pTqlvU=

`pragma protect end_protected
