// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
VUMcLMP51FX1hnRAC2sFT77fBLSA/+91Yu0HtCzTZFwncNfPM78tynt7zKIDxI6y
/OGYz9OPTuTCtNOWjMb0j9MWdf4YL8f7x+HK9HxJp0lNVPAvWfItt+jsAh9gZaIX
vkG5egFEqOFGAwu+4fu3BPeIFbA7lLgHCzMHG2ayABc=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 13248 )
`pragma protect data_block
UHPe8M8Ih8lZm7EvpCYJdokq0tAobGbbX8A3F6ak90VL8Q8ZvHUmvXc1OWQSS2nE
OQhTWqlmg/EDWckan8kggcP0Xnr3jE9vW60rfmV3GPfq6ktIhykzXahLkrOUe4aH
RBZCsp1fFegQpNmlTGTXp74VtSR7qA4PN4lDXPei1RFcu1Irb8Sfr/csFfGoBMfs
wp58xVBTDmZF1Cj2RP4yRjGGC7+4830tYtX3mPtb1LOOLVWtI7hYLEd/fQG3NPCS
rscSXP5W0lE6+5DlXph8anfwZgVSZv5OEtoWPtebg/6p6c517yl8l09YOQdbfcLP
Xpk9xslidmvd+DTkIfYOwQWiFvrT2gblzfHyONTbelEmakO2zML9M6eFikCGTl8q
tiqKzD4kMdMPFz+LZW+7SMEcTVE5GVLdIWO7loP/zxWyvz/91YXkTUFViLX+hqKi
9B5rSZhpuBDdLQIogVyZbdBcipSZG4ybpaZwgavm6UwwBNXr/tl6LFZLPpVFgqfQ
CkIAK0bfWfaOpD9DzU3MPJ9brG3Ep4fpAhKSxgQKtX5I/WfPzi3VRedNhqyXovE7
SCFRaEumSHNNIOomeK5Q2ne2xq6Wly/yr9abhQcbL8/rZXNkqYExBYyD51Bbr8rG
uNnDqEtpzbnxdrLLyYlbB/RkWLuEddSta/iq3+wZHtt4y5rm5wTO+OIS4LMxLkAD
Lyr4HIxjG0r3+hywJH6vqhD2OBVOS90DRH5nJ6LuQCqQJsecUbYzc0np9qOSkmm0
+U426E7GotPlArHTJCKXWly3N8eqnLxz1OogvGckFY1ZiVBVm8QTPJ7Uu6JUcZPj
aGs4CaO0IZZSfEujEEa8SWjlA+1lHnI07fhc+/EXDLdC+pz/WPFG0WYS3OVSxEf6
+KSz0j4IDJilSFq7ebsZf9JFeegPZzG7nyMczZeonhQ24/x3JoOrmJthtYcaTd+e
2p1mX1ti7+NCP30STwc5XGlZmk3pOrJMjPY3HBuzfzH907l79eLpjGSiFz/XdasP
aL3zLkAYLIjgB+WpRRgtMnorTtkJfyQPp1KCWVUSAl2707cnuuXDGUbvvSp/cqwC
Rwaaug8h+sRjMjGrVO3iJSKhK8MGMOIypQ2o+BEB3f8QGZzoFxvbM+Q4OLvjAhfE
XyWLhi0459Iy/LwCIviq3hh6SXzL+BLtcOxpFZU3gCx9OgJZvD0sc8k5xRsL6E1r
hXGaOIiRqu2Wly36Z2iW1n/h6WKDd3Vp0tqzsSD23m95Hbvaphu9nEi6G7pSoFiv
HDEdYXW4c+KE0gmO2ScfnyLwPK8jvwkG5Qr1SVJ0h1jXPI1LlyA+dyGcUAD6/fm0
RZSUFbwzNkI82gQk/r3fE01GpEz7fTRVoM6opPYqkcnpGbbMRnfx6kiKIM4MJaMQ
2dMs1vIDDQBZxerPlTmWOEt7yxu/YEeRQcK1aI9ox9WuwUXbAejTmgo/kgauMx54
qqjAMlPzxxCeEzTWivEA1838JZG0xmZIKnNH83L4CtBDLqrMl1L3BIm6RKJpCywr
Gf4e1aXjLyfBe9gH8Gqx2dU5+AU7H7mZqokG328XZqIqDPZO5s2fvFtMHR0kZiTI
xh5s1nV+PLhfym+rVRyr1dXctIiZbHEANwx3dTEycmCEXEOA8cFApiAtU12gkEAW
JpyqmokmHhFnNyMEeBXtSY0fzYt8+xvM2yw1ji+KkEF6f1XqTBzP756U9eD8oISt
/zH1rB1savrfOeD1PzfFY4PbZQsU1NMRpwWxesiMsh1Nwpo08FnwCW2G/sMnboJa
BszLi9uoYP2BL99wRQFJQGIUGYRUHaEQnG0yim/lvrMJu4W4uCjVCr9/CjQqWbr2
zu9skOTa+RplCXDc73iwyJO6KYZS4bwwnhoDM/UfMh6DrWWomMqWrns3PUwGseXs
TlbGW+A0amWBBBsChpfpmLFDPbwxULKyD3k519/ib3/o5gdMmJeRFTCc44AQ7h82
rQ+C3seMoW5iOAmaIpN1Cbtrn7dTs7JjiLlTKHH7UlGBNGK/cqDsCf6U5lTX5Thv
DkVOMk1Q3SCLXRZ7ioDGEJTBAU0XCUU3Hfw5/mi5gStszR4+hXW5PWBVxtlSWvp9
hyLYxugTzK//s2CcakyFDwIBB5VqEA87URdncw7e/+/NTGGfa802QFtBcmjBCXZN
J6ACuMCqtqFTxDV/bxg+VlB1QyOCWUzZBqFR1VVzijAKThgBL7/5oQjDGCN3bn+6
GmqAydKBXrjn4pwMCT8sSBjvubQ3Ki0ebHPI2i8JBITPNPlSOMhxC5RooSngMjvz
QkyJhE715eDfUsDIbOtro/fVZ5Jw0IMwH3L9jbYJRRmBniVB42BrBpvWMj7K5bRQ
5o49pO5OypPrM7lN9sC4OZeIG9ZHdyPvTMrKeBxeJdPBXYcxvlZbfWGySZ1ZOWuv
7TRldCzK8dY+vcYSzCjH+bnSWF6m6lRCY1HQYXAFMO+B+BbYeg3+qpv9jE4eCKap
caVqv64AhIhemjbxAw4ZlHi+SysbHeoVYM26iY899FyQtV2E8Q0OEBQJGV+UWcaV
riISKVJm8bNoEncE3x3UnTW/SMpIE3+y15JwIsI0VK3ixjtabsVTrLVoBAHtUWpg
lSPKKjzX43S1RNz2DA1nk10LnDtPIGG7oUPRq0UG6M4C3jpyuEtMGaodD6MjcZkf
JYy3cz9XXiwHtZY7Z1b0epMAvHGQfYDwr4Pco4QlqnwZzLxPfBphCAaZMdBX0DEM
enm1cFOB49fqK321MHZo+IcNOYJBshu1yudgGaPgvdwvTeiu+4gVy9G0U9QZOVr1
6pPUgbX4r7t7Er7R4Vz0E8tKKKSmwrQlTancLQUepCNrDSPVrMbhnEg4CBbZHGH0
oWZW6t2RgAgYGiTcqJzqBVppJO6+MRIO0CrttZTtwL8U4mOqoLQZblIKkgGxTqVK
NhJJLDnjWdWdbEEUyoI7WhZGbA7pdrtI9ujVdBvtdI2QOPNgP/nXBv08jSgIDmuJ
l2aQLhq4Hn7rF7CCyu8wv0ruODVDyCGD+vYlk+tn+VpOzmvZLfoPoMXYFPCYggzW
ve1rtuIAX4aKfDSEmCHcE+B6aR8k5YJ+9FzV6f1uDFBrVCOmFYqgz9IXLak0LlwT
JbKlIRXnuwaQAdXu4WZDBjuJPtUzPwFg/iC8gUsNM+UiTwpap9FguMijamaMQcWq
rmE0nUAe7j6d98KozswWJ40WiYv2ABlGsGjmJmNrp/oYRV4t96avkr01boIpbFVX
7g/81WemF+apkJ+e7tYXiCT2d98hkK3tX0VGkroFrpbbRZ1hgSbgvFYl07ibkNiB
aJVV3si3Y29cfsK8reNliEcMBC0mcHILjOI2D01Rs+WiFEhZ+3X1hTezu0WihZU8
pqUsXvj7UpD37Oihd+GWE+zHw60sJ0hxcqkmLGPQS1bVkX7jZgGbaOeXWhVri6h3
B2rmlBawGzyY1wlZhMS8iZdZpY3Nkp0erjQze5BMuHA0MWaLNP136x1ZCiYpl7JL
IPFqoebj1GMnzwwrZoAfefyYka9rJANkSBcrQC2xjXipQ11J3YKbkljQKjTKr9Eh
hvItIjY4W83AszNmS3rZiCq0faCSqxiDp4tr2P8txTtHjoG4K4jwMkarpIBpIZTr
7mdb6j4bq6/EkuBjw8Tscde5+F7tzsaQc/BUQovR1NfR2GFPjUzLALlMJYBtnBJF
f2pTzgwzLB0q1VNXaEbpfqeIQg+Dt/8OaiMUV+HpclpnxYGGgNX4fRZLtk1l/8W5
Jxrb4zldIM6+oSKKy3Xd7Av9ic1BG9U6jocODskxi8la/QZYkpRPfiXSq6XLyQij
9C592f9tJv2g/x99jf+5GcxFVsQ7raoKzN+Xd/v6oC43XgqkCk+/EngTxjG5uUXM
Md/9xSXdAlWnpberE0/xhxQTeBKt8ZJ3DQO1EKjcaK9rYsAA1y8lm+fy1yO8ozxa
pRSD1Knw1KYBZOaSFxcuss95z/DhsPNUpXdYcXJgIVrYKjU1tiEWNfWCLBPhTrlG
EjqAlzZ4yGCP3kSscacVGG84MnqGtPCTN6UnM9rnd4tcCCGm4vNXhb++cN1feUwa
g4eB18nxnyTD9g6dQRAIL7P1TbjkZeaVxwvkb+qMOmp+6wuaYk2wILYaYdZA4MwT
kbA7a8bYUMi31FAOODF0CMw6nuPS/Yxa1GA7jkC2ms9QCQXgEraJcf+36hy6jhqd
DHQCV4S6j2gF59L8AOy9TTo7lnnqjB2rfFCvaY62C8+r5YVEa5L1kXyMdrOyHRKT
Fa+UWYqp7ytUzm3fbvn1UvTW2NqF+nxWJGw9+koS/Rb9G90eLiN72QpNbG3zcQMM
CfTzImFEy1GMz5dXayjsa/fKLW6+aNaLL0UIe5d7ztSSmGb5M/w8WrIPmu4bcXnR
2xLtkL5e4/3KfZuz8KXCNnFd4vkBSHPsQKJhrOK2dMb2IP5b3zX0gj847GFuHwci
WonxJizc21MxUN5FAJWJqGs4kYI0PY/xG/gbpym1dpW4yctj9+jdP3xuLX4wy3CE
tJPi/TWtjwIg4Ma0qFUH6Tj4vzQJqLVlearKCslKtLCMneW4TtcUgCEu0kOTToNx
Udepva0pGSfUbJxB+T/qH6pJMX/QXRdbiU6wOJ1QskrTYeJbCbpaHpJ91jKVL7LK
bwr7t1gaz5loiGl4hdDcPgdlfWnOVIr6+IkROOFmODEQVGi4b8s1Gh3XFrwEBx+V
ereiVp/94L+/bUkYElspvi3LMvCtXzGUfypAz2OSq4JfXS06oGNc8uF6y6A2vtMJ
jdlnSGgBTQvlvXnsRvp++lyTqo7VFRm5kHYk4tfTw4N9n0F/48GumfiZrKDBMEFz
xNJa6w/aGKC76mLAb3ClpXRPoTMJaWzLPjTBmXggdQ8ib79dd9egkb5DBvi4ufAc
Ps6nCyy2J5nV4dF/T7XBY93cnCcx11t5vAHkyQI99NemlYlxBEH3+Vi7I5gN7F+F
LMlMz8TdV9FVZiSAYMMgvm3e6PXkB9VJDuXBHE49PHjcQ06QWGxHCJ8g0R1bqR/r
igbb1G/Etsk20RmLc5K4p9voBt5GkO/idVW1pFWX4CtQko+ltToji2Zr2A3yeid0
zBXSPGZxwEE+dbtZ/ie8PJP4g8obsAGZnbLK6+qp+DKJfuv62qodsscwdYrvC0ds
qStZf0eavLS492piVldPifyxjJKGZDfi96lYuq8l4cC3l7jrBPpCK51froUgnYOO
fjFhWoOMmIwfYuZRBMrJpTfdHAEaD0U4OVMqHGshBBaTonySP9a8/dSZ4gPDjdGa
PqN1DnF7R9C+ayEoCgo+fm+omOHWCxHlF0akmV7VxNFhS5IFZZnJsmT+3v1Pdie9
rv9fi9VXBMVhf/VYSU0+LGupppI/x9LPFQ20O7Lji3SMjFwJCC5nXq8BtZ7Q8pFe
MteakmP1SsPePwJ+UOBkVhfm6Uj2At0z7X3oNqvF4uJyyoshhp4pVOMz79MnIk8P
e6l7RqK5LXuHA7PpmoI2ac2OuI1FRJdBmYbuQfVZVgwLNKgW3R+vixckyzgHlYB0
X6X9ea8xHIG0MaqvDIttkL9SJU0F2cUy29N5642yNQvlO/Jf8CAzicxuUhr8IcqH
/tozJTKevse+P/0RJYOk3zMpGvlCj0+sYJbiYe5/pOqGAa3G/JcAiwfQuLZAjFdz
yKoRLhkTF9vlJbS8OLyECGuXu4VtldJl7xBQbLrrJ1jyJDt0sJdfEdbdQ21v46SJ
fozy/x1pdWx7wkMskWsG1scgEyUa5gWxKiPwABDQg/uFq8MlYQ34vWDcJEle9+Hg
EF3rAVpVIxT3g05nradBe4UUxfFAj1gMeV7hdZSuaqYRDaZuiWnCqeB8espUinM/
jRfPdse1Do1DuFe0jj5NWHanaRnTRwtsVZlcK0rYUqfK6dylZa1TLP2Bjfi2R2yh
Y0mVpTmnXFfaunsorZUV5+BaO3LCVv2dSrDHj5MNeCIdSbvFj6ISkW9fWVLRHvYC
UgH8Bqj+NzoStEbNKZEwCS8oQNDYaMcXhsjf3yvHppwWXn6dR+wnNqPfWncz316q
IENmQGC8YoXvvcpsZUiYCgyZ76Vv5oYEDPS9A9JZpg2Sm+rsK7XkrsqykvTXLSxj
ax85XiHPl1uQATdLWpepjsVpfM8RZhiWQVbA/Jd6vcfrWiEJ27lZZT+m9PLrO/AG
wzABLSHFpmrGc+TyrGhXXdTPz8/adIclJiLu0QWewF/zVkAYpTHghcKVmz3Qhaye
vyfopKzyBuUlNlNR0CNaG1kEIvdLtQoG6ymiaWUnk74JldoN/BcLeVIuhwqnrocZ
I0iWZVJKrletEei6CM61Cp51mqrgbpGPMaESPFeTujJSjNKys65nEgZIyddTh4u4
C3ftSoXu3VApNuaMbCpcYLe2MzpJc+YD96XFbFkXkc4bQnWbTJIobQf64yW3Xmfb
TBztOHC8/NO4hwCsaAJbuofNLv1W1k7Jrr6r0cYEnI6a8uqofwYm16YxBxzZiRoY
7KYQ6jdhzs8Jb1DkEGqd+f+lRNC80kJddEBLZ3rJjqAVij59umIZfkDr8dBEVZo/
PWbspSwbje/rVlEDMdVchO6gKpeJS+fPuWJV7GenZlOQ2tL/p1sx8BLgQ5tGkL3+
CeLcgSRrV3JnHsAXHA9PlZgXJRtzjjvD9vBxZLC7XEcQaw3H5cTgy7EloMnKUYRi
Tt4GxVJkIcjyw9tR0DkLQGzxfeJYskXl78oYRyQgECTDTjRUpao7y8evXzi+sGd8
IKRyB0VtL7KcaWj23Ncs8B5TYcVu/eUoes3Zs87mANc0dJJKxeJQq6gYw0EUqDbA
IPjbduCOzWkdKy8JH5hu/HCMa4cNQ3AfqwGhdYUegbViqAaPVDH9O3Jha8XWjQ6r
sZyl/Bigd2v6xHduSKhZZagYb5gqY3jz9thNyfBEWW3q52el86m7YFj6exgLQeso
muEph/FO7ZAXDJqJGGL97mc71vUCq+PELa4xhOFP3fI9KV53tQ+/fABDw4DdON7w
dFUGfGCmFd/rt0FhedX0pHLWSo3PTpfKjNP3TWbN8KZoUq+86SxZN/MFZRxCglzl
ffb5u+rjBdf6EXLlLVyPZbRn4+gRbyxnbHlbmBH05ZAx/3ogMxTPS9+HXW8Df0Yq
DWDpXKyvSqi1AojKjLnDBPYRg84HCfCIiLSPBmea3ETR4yyOEifqi7JIP0606LeI
XxDXdGdGWi7Vrm+gXLhz7BNlLVuN8oAcNIAbvfwiV78BzUWXMYdbJMZC9y8NatA2
rZ/LMYEtqBjL15FkvWT8GQBstYK6FmJYoW3tNS5/XNH1RkW7G045yIhjbjfJt28n
mmAXYkUuNgQYBci2+umZsVsCRI14ubqoDNFILei1eCLKzAsVjna17aKeX+o4dsAp
sOH1M69OHAJ9Ji1np5IfkuR5VROPV4MYnw8fJYdMsxI2RL7H8pkZTen8EU2EoNBa
RVdMoglW+wVoBG+QJJY+tZRadK80o9Jfx+KfsjN2umV1Wb4Md1G3TmNr+T4fbILo
8aFIBet6k6rLWCZleFksfJpvBcTKEw79IdoB04TXKMNPRbm62Nt0HFlhDpW8IaB2
Kk1dTx59nHAR0t01R7IraaEH3Sq0WzOngFcbYxwx0KqO2hnwU8KU03mvlHis7VlA
TpMp6hZuCmSMccITl5Ii7Upml4+bBYxjsO9lXxoAcpiZAr9SQ6qlch8UpEa6JvQn
vH42eiDjOoBUKD2ElwLixbENDjokqONw8kSMo6e7eMixL3Ra7IutuWRYkJ7LFADz
Z/hLO8igNTighBHyRgfUz9n4cxYptoGe7e4Q277VUdonRgqZ1Ctv0mrL8FoqZtoy
7+ljTVLyuiCe/0bMHtC/FuyQLzFGFpkJ3C9HHvjFZzwGw41BAcX0cVuKVGTcxFTH
pBjrGjPmwadpQnARgwvWFb+8XJe1NqWsbDxVN+3nrFLLY9r/4N44nftgwOEcF4Ml
9tF/ZQ3fwKhmDt+QDPE++0eKjjgkyoXU41DJwrHEmkficyNvmWz3pGK2JqWSVt9g
EoFJEQXWLTAFDnZdAJBhQeH1EINcLkOzSeQQxLUFjt1HRiS87NZCJyQN9OO0cxO3
lK4CstfxgrFSv4Lf/H0c0Q41D9SoxudONBzvXPbu2r34Opcn+D9xfRmQArQHhdxN
hvE7GdklHKI/0I7fgduljQjhB2GAXWw4oDcOpgICmo5ECFGp4m4HBv2FHmQvQZUA
1S4SAAf18SYvC4uv2t7mAWuHwdafOC8RDjSq7c4hFYjfzIGwOy7y3zmEC2oAwkKz
/jUyXhZTSzsIwdyxsNOOy2VoNm6qiLk9JBBG7EYYiKOajAE4PZyroPZd7IsUd86e
3hr2q1GMxC3wq/CM9lIr7glOGqd9ibhq4U/kBauwbWmDA2/kFE4zBZGeUWVQRWy5
k+4UFLUeQshKeza5FRD4c7ecxgLMupNZ46obPl3K/a4jUW0BJ/UZt80uvjFp2idE
SR3fIt7ZAJTyOyTpxamtb823V7u6cPTkptHExnOsgOh3WSEeFcI5WFIf1yU7oR/x
OfIPGj225FnS5j2TZgDrK1skjO9fwhdZJqHruTxg6tKaeeknT+340wgRVGWZgfep
IoSBK9fFoIs/U/BExBNKI3YOrci+pk3lmIJSn0KKIwcXFq8C35hMadORAj3K0DYv
VMEdeo/HOjhmEJ+w/BL5Pw7ZuoI5eqCwInJUDQ5+or9Y5yJrZV8S8UMKnqn9czC/
SQmNV5TvJ0+Uhokr7XT3Wb68bFvjtqFHfV0Cx3xOgCNHm/ONBw4Q8Ed5lpR5Cqfy
VoX7T24JTpxMm3z5cKC8b7TVdyqjjVF53vHURgS3NVjFFnW0BQMd2xlkLt77jeP8
P5WCqH4uUOF+wItZoULrFOoGfGjmNz+uVpdKi5bIEJ3TbAJmZ6yTJlGLslU6e0+M
UR/sH0jJ4Bc/3dBxPjucs8o/NQb7jxgtxzC/bku4oP4AR3DedJkE1QGTJiaii9W9
AEavKdQSZ3e/l+vFHwuxkh06WKfsm/v597ZjV4HYQFC4rbpqkL0aa/Hu8dk6AIJl
HZ2Jo4wZlHSD1NhLISELi+ZBHAXHX94Nc6JTEq6owW68J+D7EsQwWMU6FWQk1c3N
XhusQziVEx1Il+zz/K5X/pUOAfGsHg5DeVbBZxV+DMAuUyjxXLJ/gr1CUkNxBhpm
qtBFS7b/dSf7IDxWi9ReE5gaEqmA2ikNNnTFrVo/ql3ILA2rgcs0INn7+oovA1VY
hUR1tY66DUfDp/uX4XruVut9/JQQzyFyvwcV9MbU1zsZdHdRUQB07C4dk2HXhpIc
pbOxAJhfUtyCiO67SM65b6kChfCzpuJSmoZI/M6lPnGokeITxRkGAZkB6Qgub6sy
xL7vVRb4/Mp3arLwV5KCXggkK2YI0GoZFFqf/J9JSSDTSi0Nyoq7hfp2+/HX18LR
+2uN3zaYm/cO/RdsjuOl2fUBxIBZHm/GjxEKxX3WAfdwhidcAadv7NEysCwsPDNh
8Oc8HEhbupiClPN2g4ugJZCWTeCuYww3CmzL+2GAdmYinR8tbNiHnk/Y5uYKlIOS
bWF/TGYEYk9wFOt2jlg3ie4as6Bi8y/2dZzkvAtizPxH2JAhUr9qGy7qnObdNSIP
I+5AMXoYwaMIdvkP7XejrH5/uud8OoUCrcOtY//jbzZSRhvJ+hTDpCoccyVmbVnW
wSMpZf1ZDAtiU1HPbPBq4hp42AUDiogoALF7wxEGQptxoxj5bnzz/9NaCFe8Ug5U
BtJXqR4PEe1KypWNjdEepNNdbiQ0oMFmHQvYch6AklK+hjTIeo36QaWdbuDxttHU
lkgRl8gHGHpRzK+FV8isOXl4EWPyNAb0/2DU0s8M0oFUhOHLA7BlJxzU+f7VMQge
9yPWVI7TOdjBFdFb0B++dhe227yKRlugAnEygEl/2QbIVagj/uNlhydMbIbs6Xop
axvZnFNbdxBKislrEUbAPYAo50t2n1kjQ1BM/XhkcKoDbLlRnprMJ8wjdbuybg47
UBmVWG1r1i4ZoKQegafmgNmvt0ZU58ja+s9CLx7VEdr6pdQhOXotDdlaUKwEDJzI
jb7JEK7WpXajE/oBhlv5a7ond6fYGu9h5UO+vuvEVBYzfuNhS/ivtZOeq6UX4D7P
R/jabXbQAoe6iSyN2zD04X1sVwmwPz8W7l0ZPne/E7xi5EDJYCQchu9gjHsrdjlI
JY1mxSe+Y9xMR1BX4FJuSDgrabWx/7NISXRqGKO9rGqrBZJrhR4LUCv1cqs1u/Ke
1RvD24YYY+1SlfBUV9YLOG7dwDvzYUseBTcqIvXpIoHXK2bDqZgfHFeZ7KXc5/im
pa6Cp922lD4WRgICJLkiEtLoYv1VSrfJG5rMFhW9JoAI+P5mvz9Ke0RglFRkxeJY
0tbT1njBMSfoQggpL2c7WLXBA8Y6/hFRRci5A1LJvHIA7moOVhR6Zm57CXDvH2QQ
JOwGhiOompkxTESN8pzen022tzCancv0m9F3mzodujxM44C/2UBlaRuvVWa9P7Nl
OeHOBGboa+sNfsHeFCdJ8VjDkuRS1tO7e3DhHsQ+0ylQdgRKPO5tldO1ZGZgQkqu
+/OhDBFtvnBMR+pVfnUY3jcyAZn3FitiANzvzhMMR+9qVHhby7j4lHpgl6uNBef/
2XzXq5hbLx4AUXo5LX6hsyUlWApjt2ycfNYqJ6pl2uNhQMdEu3iIsfEPKYQfTXkO
aBYnmWezBIFLX0nonl4xAZ2P15CH8NesB4LfGHdIgPqXy7D9ZYPzJe1gmTl4OMQR
QQe83DzYIfk2H8cS6Dv8I0Jeas7aFLh0W/Jy4EMbCQjim4lx6c1sIPzDBMpoXO7z
8fzcx/bHm4ESdpdhU45fVvbZKql8reGwam1x0j5zw0WX3sws0EeDvUIo/37duCXb
X8/7YXJgSKy932SuA41aa3Tasx1+TtnJPn+hA9Ij4Cd1n9QwkWEj67koo+6JlDZS
uWy2z80fvoGf4wYosgTpjY61zw1XIrYsZ8dFdBt2jrvK17PYWda5gpQcSJtRPcdC
cKu/ODyvgTT9QMoiZWfr8qjX+RHiUHTOMXlr+fWRqEnoj5cbinfSdiUkDOVylBhI
IKxTcTIt8JN6qE1sgAb0hYVbkNZ4J2X3Wj039B4WuAENBi+eId0bq0/UMtov+Y16
rKJUXYAPai4ujVdSXePNP5dq19pYQREgSbKbPl9lC0rm/8R3X/KbsXV3lFvrRNqU
XlF/dmioHQFxIxemh04zEVDChgAgELjVKLBmwRXdDyEyKzxaivWOCMjfalugVVKo
eXgd6RhL/+HiLz2a+YWlDtQJU5narWTYC/Ksid5Dqnd/HpcW3G3ZAxKQVXTlBt8E
Ts67yuFRLma88hHBYYrY3BsPpvf+EgTeqZtmYv1ophG3t5aJnAjscMJhdn1ahTq3
gMGokhpd0YQsSYO9cMIu7jTkie6VMfh03Y/MggiMznhQ8+nkA16qdX8MlffCq1q1
194nMKJTfSK5Atr485Kqlkk7QRWS40CfLdCj8nszjaMEI25k9c8GaXtLQHFSftXj
xBCOU09XywtKY8lYnpfnaGjlxYBtRDrjEuS+ef7wgXpjLQkiUrFL2xExYs+6oGlG
0PFEqwYCEX+IWQev7Zdz9VQ8MKUj3oLY3fKpMPwWJMFnZQcdAyo0LOi5B5XLZy0U
p8Z0Bi1eJSbxnaGn9VvJTFpSYewful67k2HqxmWPee47hADBaWqPiJZHPugtCtov
G4RoVuLDHP/6MqB4ZZwoTP/VuPW3MvG3tYwnIOt+/g33QFmqDNhIf5JkWFGfLPUL
xCcHHJJMIHkx76c26Fa2t0yrgVlLWNoeaC6psf2ia0SinZqJWKrK5HdbsezwrPh/
5oCm8SWZkozp8v7OXqZZRT0K9kUTtkXnxfj/gqr43+uR3MN1zCQgArzUR6EuDrxT
LHwB6A7fkoMdISOL+1TqHWPRHd7CO4hK3oO1Do7q3BCHmftXlf8J980483IWSWxw
nWOpQcexcdCHmBn91tIekXGctqL/Ence/QFI/I1nYMcK0sARm163p9+MSf4LqgYP
sN7l/pRcUysWwSVFOGp8JXtLgMxcaZeqCn6dwJOPUNEHlF+Bq1hM1SaRRFahcG59
yATPdTsbaK5vBzOU22KE8HhfIW5kQjr2RnHcEhPXc+tzXax/MvsdNB2A5Tt7rZ5Y
iDSOkdcXt0tsPGuy1jt+/zkazllNVLQT9tozAxtn0x+lGgltcVzppcuXE4DeofLJ
zv9u8QCY4eYfehLd6LDr7aFduCcyaqPL5Uu8+7VYy16loJl2xyaOBL9v/19zHOO9
kqpg3xx8ruOqfxJW8dV7e2QhgHLghuIJQoHHnEW/+BywEQ5GmlV16htI9wGTIh3J
hzeR353crMnKYFJhKSQooxmvLyOpb5Q+6W1vmG3E9rWVOxLT6V6iSeD5jXHe/Hop
xTsJ/ip8PLYMLd9wjpvVFgNBrKvD9xOt6K0M2HIvTBdV3nOx98ihx8feKEZVTA89
zpLQ6bdclSCbXon+dIxEF4BJkufy5GC3gj1Zgf/1llXSANrm4YE54u/VoTqNwO/N
QawztdRhdZLK91ynBjM1Xuz2bUZBDTjjQePBoqqEX4kfpPsBYPLNLRHghjbjjAGI
RAtAhpADT/7m73Skt4/mYD3yu1jCIOAdHX1XppOsq63yx05buXzO3Jp67BZcXJEa
rE+ImWgUcdIztIoYH362WRoF3vKiArapjdj3wRL2IQKyMHa2a11e9oElPWD7sebp
qeZhbsPixGgkBsBKNzzfDZhVdQX+Md793hy3zWEtnIDetnoz9NjZbOS8mZr7xeuY
F+bZU27utFWEVpEBLfH3o4MemnYKnNSO1Owyzjea1fNyvBPn8jMive80WPjB+iPq
w5eM5w7NDMiJLQP4YYhey/Qku8VNj7ycov02k6JYPW8Gjc8+Zutojfgk+luxBaqw
QtEHb77ySY4nzMDOEYByBBbpwm039Pl5j+gwbd+AQ2Gnk6NzSMiQKZEjM267GDKV
bEpRHcylQ78PgWMS4rs6xDLVlPp3pkLkl6mg6pIwN1/8lbeG0gwiIEhQaWT7WQGZ
MexhSdfHK21EEdtgfScTTdq8lT9SuMfErOSE2iWQKhBpNchTeRGbjwyuRhPs7swZ
ml+iCoCMREvTEC53EeHZp7RzCNNqpLahNLyxZU798QYTYfBADlDa2J0WCqfBIRz0
tPR6zn/qnGRBSdX/EL7PtOFOx/BPA6hUbphcqtn1I0TDLiNGYK+loIB0AefXeu/E
sEcbZI/262N7eEszhEkELvufzEfT+QGQO28OpdoKn6JNlOOzyZ3QideRP2WrOz/e
E1IA4koMz79J0Ll0ft/EwhVVqvaYlTX3DMjtMMZmOCb6HM9lXhy4sdXacyIhrQrB
rNj3IqYSBza0+smLUB+CF5BHaP/3Djbc0F9QIXHjVUWKF+7HO3eXjgbfXWJ5GAq6
Bv9DWSMG6hnOHo4wzeHluEdksQTrXETVYWJupZgJseiXJULCSWXey3ZipmgZjol+
5vNrX1nogSg+OzM4iXFEfCAXjiw4msLiCxmPIwt3xEBaUPyX3hWAFpLFxYNrdbo4
BOgsH8Thctd6e6wCoV/aHtbH7V2DZBiM8CK1kvT1F41AqcU35YiTPvt1uMAOsuhP
FiCwqDEcujTCdM1T5YP3jwW/Cxo+TlsNUTEcTg0xQ0NpbNpqdBv25xa6YVh5+xlM
ciP2Fi6wsKyw3HvUaxFpoW/lHYLyl9fk+zjM+BtSBhzyZWXKtfreFUiwNcOyTSh3
/zriWa8VRaqswp6g4+ZXSXKDLzRMWngCWv3BkKpTdozN5EOKMwce6frizvn8eeQd
MquJ98iJi0PfvpxcPbSazkiT4XWcHfuUv4UbIEiY9HIu7zULM53fCN9IDFMu5RlW
yMQqGPsMDzyHoWmg4DYzp22RffYbzOA6xP1JlDplAiHhWivJzx4pCmQAQU85oCaY
4IPMW91dhnVGjDzVw+nJy1R6xsn763KCMd92uXKJIg1TMPmNpTSMS2vtIQMZa56b
fFM0qXqFAfXXS2cORh0py12yi3IWdTvyd59oY/oona8baMA+9ePu4yf63OjcuqaZ
ylX+Ux7+OWNZU4f+fdfF23dJSbuaM82g9OeiHbZdB3ganD1z11yEvvlM9djOiV4J
s6R2GCryyDH4WxnqR8crsm/1g4ma90T8qV2kcXHnYUimXCzmU86ouxBL8oWeXEpX
8uDB8Cp15do5n0RIcH/kCYkHZGmoOWL5gt1PFuajuWAVMUnXAmeHeMTYeYX7BoLB
Zl/JiiFo+bOQ7NTXHTTqb8YmHbJVoAe8EjWRfc099jQa7a82pMGbLCl2DaNesILe
nWU7+wlqJx7fKlztgBsL76mR8B/EL2EHRL8YnkWI22NffqI2KeXFKQyoxYZEu7ed
NlxX2eYWsK1BC5cOkQtjFYrnyiY324XfGo1mqJF0rWIJ0Iqi2q3g57YABCFIfUWP
VfyzGvR+66+NeSjIyZ1d7AEa18kDNb6dh8sdc/YHiYCYpdx/oy5r5tYVsrZFl8QW
8QwuISpdNW4HbZuaEFWWfVaiezzZ46DjNowhaRRlz3eWTnCNJTujCP803OgjzPr0
N/IsjzZngj5cbSqxS66gbOQ14lbdLPi4mU3J7TWd2yMhQ07aNMuNxsfIq1sVid0h
2oCoQMp6MMaiul3UMJEJBrfTyxi7LTUmAap7KDxyOuqkfrjy0Yau/OBqyL2zVBtq
aXBUBChbhBFnADK8+7GNXP6Y9mIMzAjWxUb43hE0nWREN0vjM+CLpDSV1WZgBG1k
BqqplcEHm/33yfkRhq+WetTfgd8kNzelsYm30mNa8JLEtoVMvnqvweT57jhC2H/e
oXLLKQFT/Jv1D7Jxne9s+xyJZPRzEVW6HkJV4GIX4PGlbPkvInDvLxJvcKSja55D
8NyELCkvHJq6IojldW3j8adz6SmEbOoY3DB5MNbknLnp1WO3cZ6lILhyss+Al03x
DTd/guU4d3BPvcJQu3TRESnk9L9CeOytxdFr++fXNJG4UyZl7Qv620yycdtojnkr
EeM4EEj3DDILeJcZVpelFxXduE7pZXLAgNWfXhKVIXAO74iv/lcCzI2HWDABdFOX
+ZHXgUYTr6BhGjX4KxqoYxV9ivtNvLXx2c2ce4Kcr4iopVkBb+EmRVZzvki8PKgr
w5gBn5o8HdRYoYEAYQgCLBhT6TPuc42Ng3wk1tYS+3UG73MmhCOWA0pitkG77dt/
98A0dWErUV3tPM1H95FhH1QxYme2KmI1gfe455lHs9kHD4HxLlK25KUTa38KNF9K
dg3Jkn2pdE3fvlf1jw9rMFRyZp97R9qV4ZESRLghX1Dh70vWqVMUw4pT88BbeL8X
ePYxdfTt1fJacG0XgAGONimmJAcSN62YgUHeI3FwYdUJ6Fi0lFoqysyblPpqZMLN
k6nmlqZReX12eOfM69V5hNmJ20rGSDTLcj/Vq0i8WE6hXCEhM6PzIcD4WOPWme9f
VWPtmwqB1NMVsqEKhVFj4sEqZTs8hF5CL83U5NFd+YzK4FtpPDvxowajniXyCP1R
ZVSdk2+xCWqttl2/Izf355wQgoeGlfAs+8ySV1R6s5bf0o06NKC28oLHp4q33NFh
B2SdyxE9Hdg5jeY6hPM6X3Rsz8kbUl+y6JUBkgkGRjddi4+7VBnTBARFi9MSJ518
n78aDRo4HOWg+MuKJdCIQsiNkA2siA8Tjg0MyW3mli+v1t07snyDt7/nby/YTpsO
j4y1sRlOE8JSEAem5bEErqoupTpjDnEfNExTF8WLXzpbolAZ9MeG/NlgorIClJeH
mO9TE5gfEyFeO1GfNpioQ261RkjbmAurdhqKceRqzgPAZ+4oNuvOUP84M5ssazyx
PZ+8xk0lbZXhi7N0SUFuL1Wx4UiavQzxZyxBJW1ND5lIgDVuB3o2PHtzmtENrmtD
4TuLlxSJtFoYgysAjOBCOe7BCgz+/oVfOhQVPagfgC0ut+l/RPJztBWAAEcguLGr
rHmrDPrhnW7Qfdde7PeDfbzF/1Lykm71fsSYMQusRP+TrKmnxKFEA+9XOApP+XmP
nkuRHvexPMfOxMREsN8ubrByDXIq9Fi6HC2OBT2iSCpcXkxvjRjcQhBk+HJ9Ico8
exx6WLvyKJx3qf77+H5rN6fTPoZV3RAwmxDFS9jqijsuE56siH1NUsm8cfVRSS0T
J2AooWBLm2CimHjc/5iMeUP/mlcCXaKVephFaeRp/lIH1reJLEIJTZJcR7cw8G/5
oASf9IrTKgMXSThK8IuzPXHbXP/EmK5pftTJQCRkLwA5uvcF6gEqYP6J8bxRAQom
PnAuaIpn4dN7fhgxY9uEoLP/DvPeyZ/IpOR2DZZZM/MLc7Iyj45CePuk33krko/J
GQZW4+ZXpI2QOF5B+/2+mC966cPHW9fhaAFtUyfKyQS324jY/sPqgh51qV+xBxJP
8y7FxJF1CsoxRsOV6V20Io0I5fW0OOF4HrZ0Eu8XhLKhHowukTXg4cZpCndpNN6s
86VuwjkDXUfAySdExG6nFUAL5hLLsGpgL1Mzhpg7PXvWTNV7+EnEccD76M/457zW
xQJ0aQHxG93+3Wo6P+eAGiVodn7EexNJYmXzIa+Ab337XfoS0VVP0RlE0cXghDsj
4B2cHpAQNNMAaZpdW/XH2nxL9nA2/ceCYtL0QiX7V911iqj8/+1Be7JwXhA3Kg6t
gFTc8HvZoHB1EWA+QUWrR52PRlTCmHLnpoBllO8jYJVaHQBv3mMd+e3vX3Ei6emc
emTQy3cgEIc+hOewoAdfEw42xGnzoxi46znHmVBW/xs0vg0Qv71k2bonJ4gN0GI/
xTzcYDOgXQrsduARTMU4W6UoeAPD0MV9PDxfytd2r/NuaKKEAvrOaeOserxj2T2f
JKfSiVssZ+7TqY6K6EEpKF5thhty03PaxOF72o7Ddz9UN7egWZVNWroHgTkXH2VS
317zu4M2t7kSQaJsg6PRUmJ50NYNsUCb58SxKihuhFMvSRqRa4l/YkDnWzNraS0z
cQPEGpuRliPf9eljkU7N0efPvDHsv2DX9iKgp8J7RgAG+9zMCMvPQ9KqaPk6EcmZ
4TRS7nusqaH4v9Wmp6t0GbYKDsgFTpZO/8yP7GOvVhTGspt6a7BB6X6OZ8klG3Fd
Zhu5NRerSHU4gXkp+RfMGYGyNlLMGNF7xn1zZkzs7NOAIcGriiJhAxk5sBnWmOMD
mY6QxwYs6J8/fWAAyxC4GpYkUIKDLpxbtRjHqvGpxQgNHoXRHWR7Wm3gmKOOFGh9
Om+Scv8BJhzphaUczfroksNoko9xaGlwfWkMEzdwFEQqa9g22HVbNAzHA2bv+7CG
n/I0XNt5zVLeOLVKvKEzwK+38P86sNoz7QxjZL6LW/KO/dgF99Iny3VjMvVO4A5W
c8woUYPpPGH3JqNvo1NSS7iOKS5G5hUh52lRFUfXt86SzwoF0XuIEl9H3YPS23Oy
lUgYaJSaGG+vdKJDkYDUQnKXJRhwac8bgL6/b+gKTyjQz2maE9fvRatSPlOUvM/+
uRX6hkHseNqDPL2iAkDSIQpyJ00fEAPq/Ivc9Fmb3wJXHh8m9tlzaNPPMK+DvnAX

`pragma protect end_protected
