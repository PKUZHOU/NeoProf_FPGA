// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
EdQ02JP12s6eY0muczDBppnbK7E0n7otwm/CFM+/i2ad8j62fUJOhk7xP6Kf
wdxTdjZUhoW13qRSi5vDPLXkmE9rIGkVgGWJ5tlspXlKskTFngk6jnLeysyn
bcHiQw3FDtrw+iumtqL/VWII7S0bk3NC4KrZrpszEWW65fdvlwEgidVub9lS
3tg8xUDHvBG8Ff+veCvOHWecH5c5yIuBoff3OLQRXcUAI17pRypf7Ywav4F4
KraSW17/oWk8I8MiUKp1+glMEL/yNBe9syA6kXG/Vyw/sAeLKYfTpQmNJVzd
uMkfKzBiNGGURFXXz0drcSbnMh1Qf0kxjnuDeeDWJw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
DwOlKPv7k9as1MwPIRES00rPGNH0porzaI8rT+yzMyGrREUP1LHiNeqi3Nsp
UyaR6sDPbEk46zOJx+kBPq/IEAft23UEeJqINHp+dnB+2xvEQQhuANUn1TDF
t6MBVcdqCtzo8am8C/Vby3eRHbVp3iPplFtiGpBMqbcKjE1CBjnTaM0xZ5MX
qyLGIRot6esFDhG5drNHF4Pdy1WPuyCQd7xjAeSuCD9+k/q6ZhFs7gSSlRxH
7K/u8ymoR7AbQZLeSQmDd2yAN8T5uuKZPzzbFc0sjvW433w2eqcGWdGxewS1
seQU/y126uMyEXhylrI0HwQq+h70PrN7rwK5rkgAYg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
nda7qggtc8qRGMzEPhziaIXwjWIJWKY7IUdx65Gr3U2jUAPRiM+HARckGtCJ
dCh2gfvWX6GwQ9FQiH7P2JOLyctOxwn/1BV3xLKlV+WYg31lOHKikDmMnyvm
t1QBV5mRdCBmur09p9BBIH2DT+qbwrCvwjBxCfH/zhVJoq7M3W8SlK8VLnCz
da9c/qbdw93R+8a72nT06JrPLBzWg9lTITPKlY1K47udz8XIC8vYUc8BmDR3
6KGRteGpTgcDpNnxj4EA3ju2Hgw1Cc1n+XJcCsl3KhSTqaaRQaWuX7A1vJ2x
m0H36TJYUVqQHLQ4FJ1ZfhDJmW3Vb5Nh1sNApYxEUQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
l5weCf5d/6uGtm931/Kxx/TT/v3LNzg6cyqlreY5GG0Q3xAgj47R/JneHxrR
clHRnFXYTc/cne35vjk83QSBKVOMXYSRzwu9TLjIYW3vfK2iDEH6hQZSMT0P
O9N7jKvcDjcPE+sO96E1tO6mp2a1v+PmDLvWfsfQoOCogX68kFI=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
DX15ZeMYIoW0DbnFKVWNVkZb7BBS5CVcfC9ij7VbPKu69x6/tUR1ydZRNgj0
YRqkfS3tj6RF2bpZk7dV/U3O3b3jsvxYGq2DL+vRco2JsKfjtGm+SlqzDKCY
qTyBKlo8AlIzMVfRpaMHZM+Updd8lxruqHBCNg6Pk8yAg6yHQ02q/940l/fl
g+ThWKk28OKahcdPP6TAVcJCuEDv7YcW5Kt4YD6vQ6VW2i1DHk0ycuVWO7XW
5MrkxorpuVf4hYJ/Pn6fpe9ADp/lD8gHYYvM7tsWXxw9guMeZpNYR+b89OQR
aYxkvy+/6Ya1oJc3qUk2dXSp8jvFAmY3E0mtCsxa9c/pNAEGC+OLAskzn24c
bbN5deYR9Q+LE3H9V/Md40t6pqiWKpAolCNphOY9UxC2O2Q31j8jmJs9jg57
hJki8bkB7hAWax3qEsqLsiuL4t8dI9rTKu4/GwLCoLzGnbu0I8KrCDqSuPDT
bR+GGDWkqzyyyrEqPJSn8w8MjDR4Xz/W


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
SQxR/8jq/za9nD7IxpMnMPigxYZXNa58/le1PilJozjR1QcTJPNVXcstq3BU
ZpjLIGwBLQguQoR11uZXeUf/PCAOMoBpKOHoMFYv5eNv8/rQIuXCRVbXCeqa
fMhFOPiOWEG8Qxl8VpocjLaHxbHkzlEBWaLQA53yoWIXYAUi9Ls=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
s3FmK9ktjNZD/qvAZnGV3FXj8i57L71H8PvgyLPcg6DID/OsNYYWjeYsHEEP
nuU/v9ZNZdarU3TgKhV+YMnMzKkRlsvO3G0ww7+30ofJYejyNINCOv+JdzY6
HcvDH//ZXHdH/6Wy0Q4GeoBxXjS93m+39EUs1N4cpsyUIx4hKAc=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 6688)
`pragma protect data_block
zBP9ruBX3/mGGzm9vFBArY6rneGwkyo4yQSroDHv1MO/HLCFkY7dxkDEwX/J
X8M+kMde7Hjs6dMHtij8vX4r6GAOX+I6kvbE3MGREGzfR4xrnp1bYF/Jgkfs
2DQeTqWajROT0bOedlRRKPZs27hayuB8740FxNkU+/joOuoO4VsHgi92kNxH
iAfuPCuBdSC1pTjuY8J2pGnqXhlBSP6Q/A9CDt/IVUw8A7aa4sRtux4AX9TT
ta7y5cXIUsq5/1xZ3Y9fXR/NImo+LhBkdfsBH3wBg29Pq6hMaBUnZdp4YHGu
RxlAd/5CQnqxnCtZsy0h99eYAB4WI6uhGg804lrwXxSlmrILjvWZqHd2df08
SZCSAs8ZLg+zcJqGWJz3H05qVbot7KPHG/CJkjRMDrpmvSHHNoxSE+/IENLs
5qYXCyS9dtp3gzg1vE7rwYjEVxutwR/MSpb/jkI62opnlmOrm2TLyIb7HI0y
/WR15ZIOWp5smXEVcTnQHb5f3ZxwTw9JJJ2hyzVuKBKqJj/LSJeDM6d9c6PG
d0VWzn4N4+DduEkfCkfMlTPZ3i3YRftTgwlqQt311oUYEv9cfEb6CzRcr5Wf
3wxPAq0BPBiOq2QaniDDoGLrr3vdhV1mV3pPTauz28a8X84AKt5RYkvkHqMg
K3KQ6ctWsJaEwlxLnIfmyUzt49PopbLlfDYzwjxfo2c6LV4/eCkb9kWIPGoz
YbpiqUzQqGGr28E0xdRDNOp/SHoc8eVnB8Gp8B+AzL/BLpFEJaqpCkkMk3lb
OiUZOv+2rENt9vgcAa3v6xpSnlu6H8Ssxr5JHMPgSAPL0jUb/p7rbbONY0/6
z+92jw+PH/dK6diyKespWk5EuV09JYqZohVds0oFK70ePu1SXuD5jHEjDTRf
IobLKUDs18MmdU4SG3ylgVSdE2xe1bwEkD1w8XyU2pewKskG9y5y5YKEsqgy
3nPa6CguEFH4DCCmLvQ7zSCFrdDkjwayXaGaqFg52Dyz8vsJ0aLG1M6N8JF4
UP9cG8RtpmHxnHOta7IAtAVhr2PQ4/RXe3UqPkHxtvXftdwj+uGJ8CV2ijhC
NnIglTxWtUmB5BOP/lgDpT8K7xffknP2CL5etLLLK4cCt6J9omWnOmwvkRi/
VGrIg/V0juHe3k34Fir1C2r4dwZx/3UQRTQ7Kh/gdpTRf1D+hXJYeX70kexE
hXmB95VAKi+VxlSDsL7wwwRletzjU+G/iFbdicjzH7Zcbws5QFtEvKibW3to
JzBagxBuSXu0AEKNfJ/OUUZHsjSP0WwGwBwfNuJ0nZ3DA5lg4X3MgIooUah/
EmaWN+1j+cfnFCU/SxNIHAhroKrF8m92n1ZQfSf/8Ju1giUxkZVwYDlnC9uf
h+TuHPyvdsiahyrZFJ/6gF1MMuVFA4RBnM3RoUlm2pnOFk27RdfOteuDN2+3
OysQD0RW/bJvoi5gHchd0rUqtXDT6oCTc8sF0vFng4Gajw6PMw729kpD8r6P
Fz1csDxCreJWpshGyM2geCr94Cw5CCcHTmDzzEbHdB4hefqdiRSfrbS7kG7F
ceKn6JyMlJQMyZOg69+cuVohouL2oIrNlYLJpxmENeZts8952hBr/oB+GggU
zyT3Se0MR7iHRkCy4wkA5RlkBkp4eYJ7zMGFRtlyij/TYkVd4uT8VNiK+7x4
1fszwxONhbSUpfmT07qVmsBQwHX0TFBSJedECkL5v/mzy483svCIaYZHUE7r
SgyDT0UF+Oi0z0jX6fHZVNFWnj0QUnVhsWnytLVu++GBkOpzqwqLgzsJnh5K
ooCFN18ucsaF4V8PVHAVCtLSnVFZYEA6hEP/u+C56FfrFYuXTxdA/U14A4UY
Pl5XirJWSY0nuvdBeETgHYrrTZoqaK6k2fEJjlPUcpDUXzBTWA53o0D8mGf4
FGzRLxNh+BjpOvLDQ1ZSBKqEsNbiHJ1bdMpZCMP3VL2LTDyQln60hxoZBjHa
+PZwF/7fO2LvezIFxg+UpQv4RltG0b+TurcV6lgImSWoDZbYvA0kwQlnxN4V
E52kav5Yr9eFiDQjoz6VXpCYHbeA8qGe8+MnPVUjCM3X9EbG+UWqPV94B/nq
ESjCNjALvGHyi0TsPtz3rtNaklUJEJIf50+if64bT7uuqwrKO/oKi5HfHiCs
CYGJ21uTGuxKkOQu+z0XlDQ4hjKRVb8hAS2sttZZ5oCu7qaxjtHXEoWiUVDR
x/tzPE0id909eLa4+2cASEN516CqM1Tzas2AwshpYYrUjMa4zgELkEIdeOjj
twoPDdSbIVQwpSV5gGl9FlEgMWBVM+SU87GyYYy1TwX2BJN9OYxLIMmdwJJq
Rf/FT2BWNzLbMIrBUZj0quc4oOu8pBV2gHHAt+qiREURtVWx1YxbGKCZe8P3
YmECU1klyolWLsT38tUuUdOVSHZCo1XIfACz6lA0f8vEBtVGI3gvJeeehiv0
TnHUn1iTK4zPdDCzpQp0Vse9zvdLcbWAoxCFrRfvpno2Jp+hfx70w5Tt1nLi
0AgfkjsqeKhNErv3fr1Ke2qJV91nWKgkUDG4NhiJuAiaBTuO2ixQ8o5wqXTV
NrHezW9ayd+zIfzHfF0QFzaGFQ6HR+Zh5oTEnUQFp4DAIi6DzT4kAvuYMpy0
aBxot1Mc6eWTY91iuwHMTcpS5S5WjubNLMKb99Lkav9GxpFDQJCGWe+wvGv0
NNfBeqA3n9cDsefDA9N5K571aytLX8gIVlXkyDrftQDjsDZb9YAIdq8y3+hG
w/ZnGNmI+IVni5A15CureBuXpGs+j3bKxrYuKujiYxKlKNgfwX8IJG0mVwgy
1LTudfoVlUlJHtZVZ86G2CowwTukNOJkZpLItjsZ3q+5Hiah8aDcIJRVLHZc
AzNMbb65kq+peObs59IbdD3kXAJXPgL+MnHz8ysjutVecuMIfWhulOxjN65m
sfXGV6N8C+2G3sCKO+WzoGa8kCPtaS8ZsFx2kz9yqmYv0hgC/L3UPNS8s8kj
NEq3kntJziMo0Q/8kaKwuWjPY8d+WzrPsaYTSKooTh6RolAglRMvT184OSaB
SALytsWG7swhkv7PU/v5yewiFJsb0p8kTGOjol4iHpoHOetzzC/ASTeTjJ9d
9WKCDkS8ajbOZsssfqVAvS33D1I4CasRNnptI6yfH1kNIDF7gJw8X29/LNrh
k5yf3uMjvGnuGdUgX2rS+cUOoIfu1Yiofo3MRx8YjWnOYGNlYq5g8XS49Zg7
FCTZB9pI3q8A2a1Mkapkkls0Gz7GwOk6OWSz4CaaDDzBtAWbqDMU8xvSoK07
lVH7eBfB6LnaT5HXOPUnSn1jPW4dSfcaXzb39QejXtkLden4AV62XBR+3LcB
KF4PZh+4Pn63B2t27e5sXReI36YRGKY6vJP3poL4yhIAtbVh7e5BEcfn3+0i
xM6Ng8u5V65Ih8ZD4fGEI8n+B396QpHE5VTzY47HR80L3/YrAN575m9sTgLV
ZA0V5fAisA6+LRJwPApEdFHDd6rI3CBdyTwqRuF+iZ7BmYIOae5Vw0nlnmrH
e6UJJ0hpXV3EoNCSVDdVfuhDoUciMv0kgVHYTt7ZFkyOSYLDLl/l7slARUlV
ghw0x5kjC4+vxBbBbAClSepXkG5NFgUXoFouQ3i9Dusf8s6Z+yxgrotQeDjV
RBxrRjC4Lc8j7kQd0PAKumz7hE6j/1z+ncK/3hh50J2SrxfXx+ofjTdfZBB2
QahHaeMmcMqRuYTyKwc7b3sTfTvzu2VvOnF0sw9g8UBF3SzMhG2ggzAqrdKC
JyojVCleou/WXtGeORU1LpZ5DSDj1SVQjCrTdbJL1f87mzsIqOJch1nPJ/dV
ON63F44r8d1UGOlnsogfD+rSnCYWITSDkL+izLDcLzDPWU+F3NhbxM0PhN1z
Evb3rTHOQnX6mMcHf5OOQhXm6VkVqqhAtxeQUPjWhbIO2Mkh2yiDI2MIkm5m
XW4rqBeMC4C12Sf/qcotKxd4NukBpuUC4Il8u6sx72FUtxDT5HjCgsWraWTd
Z0i5ySwtIDuu8lwJLDr3oMvGDdPFWPUmJlIO0HWCrV6XHdzWkZhrmSwlkxwR
AtDC9dPD4p+L/9IQL5J8EtnwOCgThIt+q/GGCKL3oH7XK2pv1mt8gSyelKAb
esaHXZYx9fI43aH2OjgGQyNZcDVxhfwzKZqe0dL0mZMYjTOFxw30dtQpB4OJ
/qPcC9s0s5f6YJC7VuPk4B+xvQpScjoNBYY+4RtaiBBBeuPYMgEaLQQh2W0s
J7pAK4p/dwWmBf/5zs5gsDAOSJd1Tprvo+YTtYBUF3vhKw5DtkIr4ENeXzs3
4qXr3TRwYP0dJJccRLOmcWU4V67PSYK9U1qsQlRA+auINLHexd/sBNWk6WOL
3WQoy/TMzc974+Uzz9bS3BxbtjOmb7AiMl5Iwv4Uu//l/dA7aVUi9/l8qnHh
CaiDaKrZ26jlII/Ug2BNbVR9hFCN+V3zI3L4NFhblNlU7iWVbMQLGYBzj8n9
q5OH0MxJRFSUVN1Sj0txfvug1fIfLpe0ubq8p2Ft9e6UjRBpgaDhChmkkZqn
XzbnHHx10/u9KrTNiQRakR4RQMhiTm/neDEbcTXGpppZT/Xy7SgTevQIbdRi
7NIzrTob5TDsuTpQdt2WrbAXCqMenMhTMwUWilyGe76BkdBZG8XQOq17cU0a
B5PO5fkU0gogK1QlGQRLvzAG0ym5ppkWbVJ64VKGpsOpjNzAH93TXyuML8PE
R0dGprvj1az/QF3IDD20ex1oeJM2MU267pclaM3uYpMF8gQa3OFp3MXc1x9X
uFhwr22jhE65GXnJ+CBeW16x3yzuwaQXMVn1sjTXyAnh3YsGW0WIfRkV7SgN
uNqhdzakX2hed28xgwreaqHNLoCayctoAwjyRZNv2H6QVa5zYG/dD3CI175A
ykrTnvkRn5RJcZoxAKyV5iFhgGmJeVvyAJ75IFcvEK10q3k6LvvH3YJTEn7b
VLhUEk0k4Y4pedRg2WKOSrnHiOqN5Dev/y72MtBP3lPvdBip9izWOgKSycje
NEFE7aBtywKdBMfck7s6NIYg1qu71rJNS3xZXWgiy/04dFGoaawXs1w5lduc
5FlHVtj2ifhJsyzCxyjRJlxzMNwWrGsapeQ2a8llw/mcH2M3RZ+hn/AOXi97
q6jFWAD+pV01qwIKWxtBIy/tRs+zcLjfST0Nehh1NmWcMEhdf5LnJmdjb2Yo
yFtphdLuXtk7wvbNMriwKBUfs+LS2uxo6Qe6uD+UCfRtw3wEvDWUW3FIu0XB
e2QDjgcqzy72g4NJG0AwQB0tklpTQmJ4w7N19HOFKPrAQX/Bg7I3O2CM2RV2
xXG/kegyGIMKreaJA/EioI3C5SNruGc/FL5jQDUXUey9/RgjO0ciYMKW/DXc
I2ir5UJqA/rPHUd2FX+//jIsufCdIGoLuZ9d3++KFZsZDCmjoB15OQM7zE/F
shV6GuN8KAHXclbYOVJnTTfw7vIkrSHGRGeJ7eSZfmODIzAXRgTGjheNKF7l
Q+y3ywswC3Y4+ANhDocnXhQCeGPM4RPXzkqKzz1ffgIfNgmkXgEn2VfukGfP
uKyrTBWRvebTk/y+3ExoiPzWCWWjmRLdn0S8LciqmENDs76cltjoMFEi4T2D
SdcHi4OM61BHk37UoYyhbc4LscYNk8KrsJxZdLEdKw/DKKfrBqD4a5MtTPTc
/CgNstusiLWPOTZCO1xpeMzImag4xmKG2MpQYoFHNjNjI3N4CDYoEmpSK0R+
zeYWhmIMK/Xlhnd3Oqc6JojdLnc/f3NEfHQcc1Hb8DyiREyRVh1UC+Pj+Y63
yxOmCaoWJ0a7KR/oop1ym6Z5TG7stSYjGyb7ofQqazr10uC3/PB3m5D1b38v
H9wFBcAdONTTZg7roJWlE48urCw6SFAb7T5Nih1Na1H4pusrh1p3izlnW0yo
LF4h9OsGCowzgSfKaMGSFdDsgyoja8DdayZK0P4AdZsrvrWHHxELojQkmM3w
CFnMAHaD1PDysFdElsSguSdQxQj1kZVqV2dfdsAoN4Lqd80sQJLVKaPKEzfT
Q/n/oq/43libJ6jBuo6fwn9GKpyFqO6f0Wa5LEK9tivZizGdR7fpsnJ4985V
85SGLUJP4y27NM97s85V8PXpKgFthnMDJAvAYdRkMYdZTcf40xiyiVtpxTcV
8zi98V6aYKTEFerKeNdN30wAj+/8eNpaZVdx6vZ8vBVzDFLgSiLPEN/xzO2T
Vq77/i/WJHg4V/AvGZwb2z8i5nk/XMEg14xqK1U3gssOuH8ZcsuLb156VedO
VAIaw3O2wB6zKhSJ46K8WBlpjj7UXL1kTn1paVSitEkyWAeIyL3c1xAVu6/u
/Oj0t5tpghxWf41Pjrh0q7wVTcSbbjqMwb7WQsNMZOU6/YqZNeKU76yw4kVG
lj+GRj4/uiXg13lme0KHXgEDvjD0YXByOWI+NnKBt4oHFAP4h+NUIf5muNXz
/VsvSKMkxwWIxeKJM0roKYkbr3PwQihKfOJ2bA3qvaDxUmWs66AS0kjEcKG6
VOdS9SiAPkCVFKEpoglRqGHmP2OjIatptSY6rqfdzyQjQ2q2+I82+Fya5zAl
2zQzyiW/o7tJfOkACx+tdPlR72ioZIiMh2p7T6XeFHA5TwmnQpYfANnOI6L6
nyeZPZeGfWIdqh13957OChdz65knN8/bFRcug5yHx2jcl8fYNKR2OxtDQxIb
VjzfAH71IzXtta71K0uHC6X4gROQBTsOEK+FOOPLBH78Pm4i8uGHa2vifqu8
jxselfBjiBnfhKshIsvOhrVflvXsjJRm8QHA/+WWDVorNVvTEDWOG/fK9Gwp
dm58TauCRuBQVCecZi/7cUYnZogF6JowA8YXXY3aNAn2Xv0i4qu47rhsXbNw
QpSNZkIP20K2JVAKRrxXzDP14mSETmrKlACpxgLu5tzc8QOzyYScTtWjkOId
1rWao6jLq6eYeu+FaR9KWcGcxzg+Y7gIYunmAZLsgyLJ4D++w5V1neVOfTwM
rTyYesGkiRMaRknHb07S6dsGvI8yUJGak3UQ1p1iDfJRhxTtzQg8utMUVF7R
OU36YYtep0Llh5GVUc8F9OTlQNlmC9mtVebn2cT5m6G9mKpVyVfKUgu2i5TS
lzNhQ27H9IdN7P3z6QtIe6UXO/oARuj0mxdSjT1D/nsuFtCUJU/hId7F9bk/
W4UKR9C52hfoUri3kcWeyAJMif45T2kt459jvYH03yVEsz+096mFJRIGthfI
+QDWCDiyt+1XQn8+rqkI86T0wxtfw4EtlUPhagNoGg8Z/IDW8RFLls2cgAgk
A++c0e/K9JX4UBsDdKM4mQ4F49OwUqMANiHuUyY6VqIYgW9YXrCPmm8Eruo1
UsZf8hGxgqV3ayUD3BA6LKCR78UaUNDPHe08NKOki/zLIWpJg5aQZ+3qiiCd
rMBqMlXNuqZ8W458Rp5/FXcWZBmctUifUHQE0F95EQz0DmndoGiomUUKdC9N
UP3OfzHhmqV4Ift/oeCld1CjDq+6P1Rp6Kf4+AbnKWjraIL44BUo/ZAxhkA1
+hZhMpI96jHsCGJLktsrxiTWvBOpriSPUDs6QLspoNpguaxyS+BYGVkdA2P+
q/ZjoKqlR6N9UPKZLh10olaur72QHI2+z0QQ/L6QK6RpT5/zoFpApWUr0K5q
mmaIChN0kO+QFlW7WtL2p2aN133W/MIy/YVekHzrNqZ6tTd98Oavu8fPBhuW
4phBkywJQGFd9uboL4sZzxYKm3kf4tQUYsPpWhJqpPiRw1xxJigaT40V5xLp
DaZksW/QOoAv0Q86gU80N55VHgRpD5ocJz4/DFr5safIh7/Q2xzD1uEKgbzK
JTk9cpihUDjl+lmtVNW5UN3rPSZCmynlGj0X9qzpfx24DnVv6kqzJSJkCX6P
ZZ+nPIYy5/Z1VAhI/7UZi4UOtK4mVlt+q8oJjNXVL4EBIsP3UlvzaZYDSDCc
uI1Bp5SYiiDGusbM/vLNfANGMJTeFCP5arUBeJV9NUMKTQXaaRyA2U0VS7FH
XwyzDsEawZyvHAZ71XOTmzS6K7EcXdeGBT44paBRm/74yYI+WTwuBofbXZyQ
fzNeL3OvRzQ3JRAbWgRhJsZ8y+ynq13eZlQikyO5gZZ7w8x1NgjC+xn4Q3ss
1HfUoi9rBrGiJEdRyAcsWdXQAP8e6EcguvLVFGyGQzB0kxVkHvzickfLGIoE
8ncvu7bzqNqfG7pXgkREoglVMWegQgiXb6BJvMliV1se0Xhjgi2SMnaElQ8m
L9eSp5K4JCTyEhcq2sL9DOdffnpPi/TPfAdccl/nW9j6pa7wdATLciI9zrma
gmvlib7zGn7ji81ca2zQXhBK/uiCUNvnMqCSdGPXJTcdCiDxhUxht6M5UlB9
fz0iHvZDtuW5+gGh0HUhDDtFd7mdHSVADwCdCM6hafL8ABQvCHN5mLNPEQkz
sqvloIOU5gPxOJBO9q/tS2aVqaC9029TAThLnq6LK0VoYs4D/wRmh5upYvOe
Y20XiwZN5eWYYwIBntNDHRwLYeZFp8164eGrIoIZKrxJOUrWrg0NZoMSbCXt
PUefzuiUNX1IXZVr3RYXSSG+6DghltO1f4M4ZnHtM+RJKf3RdYJoAQsH6BFM
ddqlWkZB87vEN6sT/52G9Wzj+qh7199cbiR86fnCoSih8glwaMFYimCqX/zN
z2dE28PVIyQU8PdqruD8UXEbDnWpGb9ftgHxePNjOUbdtRmiQy9ANl1RIaVi
lGHcJjZ900Ea691vn3kXDbsih1djuTZe3X84qoST47Ds1H1aslRXu5ck2wuY
fRuw7yboMIfQgmO1cGWCmPMfFSbQ6Nug/5aNb4q2J4Z2s2NWAs08sibXcrTJ
jxFCSd7zmNl1xLrYHskqOjaOlo2+h/za4nJz/w==

`pragma protect end_protected
