// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
JAINYwmdv5ZCC4jcVoCKZ37ax8Bblj0BhBTT8NGaRLGoriS/MH+iHIXBqAuh
eBNEoy8yH1+CLpy4y+ag+hlSTwo9b/oGTl96xHCqPLXsITIw/MgBh+fnii/x
d3S1YniFAd4FvANMBmR1tRKY9U1uwbrtmZ1nSJtRS2ob0mL/l3sgjSJ9Hw4W
9xVndTyyO5/JhYfUQoBErG+fJ/eBhGN6kezWzV6nAdcppvDYEdn2hnWov+XB
MKvz22l9znPLJ6rYc7SY5qN6Uo05XoZuMnKQX5aqV6RZwj7eXwBpjHQYQBW3
3yU7v1CACEIMyVDFhGeFLdRHOMhu06SZls+JdSOApA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
lTjLgShNzOgkXRwA7eC5e3AwybJM/QbpkBtxK5CeHKNgH+ii5/eWaSitlklV
X8koJQKz45YgxZX9KXtjg5WdXKC9YEdhNaMJ92CH25wXNNYdug+kF48fB4Sv
8nNQ/mJiuFOGsQwOX4K7W9Sits4fCGee19LKMa2MwpHd2TJa23Kyzz2Kiuqj
zbyqv1UjRC5uMzbCfBwdkrchyFiJVW5swM83PryYDGPQ+LVRgVGmqDFUZLdH
l8uKjKyxZJvimVrMGGp5dusEKUOTC0kSe7qTQhzahjZEyqHtqfRKYCL7JUSF
b7n++TMvpZc7nR3YyDgIlnsV0bzhND5dtfew0siK7Q==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
hknMZmXi7FFWu/MrNQgdnEwbWliPesKVX7c47QABU3NziKelb+gibQrH0yqP
4xhR4NX0ycTUNFjiEF8LNNkM7dSSspfcheqngAfuYgqTJdXXjuK9Twpc+GbX
h8CtcySlUURn987tcHXTvURIjL+Ru5bwoF11QjkMvlQBqNO30nc0YFX/bVvU
zw06xKD82F6V1WJrcWPVMblMfEjnIGnvhN/WDw7turWRR5IlxL0I6xYRkyn0
YNzlCVTp0uF2cFoDWhTouFjwPmWSb1lhoMZhO/mn+u20KrI9uVhurAX9PyBo
6geSlzEA+JXIBNOt40kJTT2JcFNj913mVSDr9qkyuw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
L5Dt4flNmM7TYt3+nNUNONK+gcfBQj176VwsLA9HQaRLRJ6vY+ap1b5aba1c
tEY+lufeNlJXC4E89Z5SUI4jFc8XdvlLKxHtIA6CaagWTLgeIXuG5FaWE0X9
yFbaX0MJBPt64zeYr8pRaKVJqvEYma3fUyPNKkW767IYrqgIzw4=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
oV4skve2C/uJXJ10s8HwLFev5TCPlhh+YNpk8XVYQgpRO9+LziOwq+5cxeUS
+kCBid0xta1tQvY3dliXHcF7E6FQIYG3Ti3pa43ptP38HWbmPZEElcSCVNCX
LaSG8AGbhlIfMc40rmzKlj7TSlHGzB3kBrX3ESHpj9ztaBO3o9Iu5eNb/ZWr
ntq1Fu5/0RL+zYv6pODDPadjJYRPSbt34omjELpJpviiVtYByvITXNFtNph9
fGd7/bJtS58m3wA9bX2oR5/bWLBRJVWZM+/pjgpbfWjqHNE4TfkqS6fSYJ/8
Arklv/LJYiF7jqmqpMisMhlrV0E8rNWtACrjq8YMFE+UG7JccAqUwpo7/uIh
eHGsWNXp2SvX3uiffTpbVRzeMawlLdh6cjrMRqVQBV+nFFSDO3SLxCLeO0Me
E2N4flX7a7vj1v0cGSsMupw/SnTK2Ohz+QmHdknCHOn8axP+4xaoKBC/dzaR
A6les9dUHFI2Gt4zjiP4DucsHw//EyQ0


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
GCuMXTgpz/Z5Hz3pdiEuhty6Nj9L+2S0+K4n4WCsTdanTPb58xHxQ0e+xvG0
NAN/jWE46ZR3eAig7VIVR4ZFcxqcKScC1A0/7bgEpAkLuKr7xDQ7BZEvfDCZ
gb49TGvlMVTviPGqpc8QC1u7Lj71noLp8MLtomcT2DDOTjKHxm4=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
AugSbj9003QJe1vOoG/eUqFcF5zn+cMO2zDxN0TMsjuXKsIrXO3vQ4CQq5Rn
zKHObOg9Kv4zKUyHsUFswAYy2ETw5oSXGJdMn9qavE3eposlFqb/LDfs3RmF
DS+eQvcvi7fsjulseAPV7Dz0tzjOEbZH/RmEHq1uRosYOmajz8k=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 46880)
`pragma protect data_block
Duo/mZSd+NrsuFYByK+DJWb3+qGJXwGUQ+S66OXN07wibwdRnEoVSL79xN4U
Cf0CosAXBN2W0lY3KuX/ooWBB6TfQh0TylbaGjVQU96jptAak1w4emFnFezg
YpuXjEX70jVENFa8EcCFkqrYf3mlDRmkSP4Cw5DACNZfz/39fSRbm4dT7YB4
+QdKoaNYw2mpjz3SzP+cA34x0KWT7cCabg1OUMjMQhw1anwhAKZdm3fLuKTq
IwWs82xWfaIVmwe6dLH+ob36etDJEYrkoYFlQ9LaP+e7L1yRS1wSui8LvDxI
A0K/cW8Ar7gfORcGqP9GfZjW0ySijQEZa37h84YsHg+kJ6upVVOm0tx3CfBE
Asy8KYCcpIG8gIie/j3puzaSZ/UJjHqcxhOf8sg8ZXuG5IMjATbO2qTuwnmr
r2CqeZnF6uRd4151gZTWMvZNA/vceTIZ+hdARG/pp8+Lmroc6zU7a3JrIqVZ
YdBQFnK+WrgykYqn094MhFl3ZQrvNYlSWerr6ibcRkfc6i7BEfsVCwaQg5Nf
RF50EUq6QUPtcF84D38jlQMTPucrRGBXckic5AHJ7QFNu90ykxOUr+nWWTyJ
y1U5gQyhJ7XUThKlpqIBRp9aBF/uw7WIPoNUfydt3+CuFBmjtpopcOsfMpRk
flkL2TlUv/NQM65YRBVMxkgi7cpT2813bvoQE9iBhDTYXEbLz3N1PX+NKsES
YZGl0MlWL1ar0WpzsZrw5mPFM0ywkKf3MBYHARYgeCR6/Zz0IZJNlfLMmcjp
mRq5aWyLtH3MuTiwl7KnPhaQakzGEr4gNqACmXJ819bJSy6iLE2zCWmFqeBB
W8mP7ztwcHr5Z3dbqR5+WkE+SaqQFWjwCRjfb+tnCQBK0RVDYkhATHS/oPDW
UviGTKeCHavUr0YSz/oFahZJQesw/7V4kvMRqJ8Biqyp2aWGPLu7jMC7H89M
KwfYevuPFF82F32J63YgzIH1HXrnatqJtathOfzjln1f4NzgVDgyyk3X8W8n
tGMJOBo8gQg3sInHMwfdAuL2AMlRYm3MBgyvWCaYBPzag6/C6GTw1SuGZsU/
nDw7Zqocy/Hig7EvPc6+90wQi/19NJGZpUk6rfYsEG7Y4wjjMGAkP5ok6oEk
kjs8uQT8VIAXX3acfJFCiAQYpMH9cRjlxvPrPvV7fyJAbPph5QYgNQPcgY9C
rLg0j0vD5SvTfp80j5RwnNmjTIdx7/pITN1S02EjSlKPy1rGRcMs9x39kzh7
L8p7jJedJ1p5EoxRMkzodSfvp7STs7PTvZ8GVvTfn7Ij/uJGGFqJ01/JSSIf
NtqPv9SCW19XJTp0ZEo1a+1KcZe0T4PpbXKbjAMk5IY2f9U+3aF+MFRKyaE9
6Cgw6DvQ/xM9Zc5Ey6YVRvnn2IT481DOODUuW0cqtb6cX55qu+my5UG8HoC2
53XrQ1NpjqdRILhXqpGguL4bAODwyMVOnv/uGz8K2aBCzScuP07T7EO+et7O
6YTi2Epm0f61u3htQstfYXb+1ZsdbOZoMqzFXlgcrq4RhRrapxoMmOyUyNQ7
rn/Au57FOAC3bu9b5fM1lovLqqnvVuBt954HEuQ7vBnK/qdKScM3Q/vfjNXt
ycnz88wTCouMgccCqi8jrdYgdu0vnNPf8oLDlTVa3sfc14pgpLruYZoovgYC
QHUvuI1XG6+KIVf8X1eoShfjHQ9A7wthQN7Zrm4fFGvQqjObyxmJwegCQFnl
flJXYLPlAwD3HXvr2rGuJvmEGbGI/ImgYXIH4qNPBpBV/wQQp0Fwq4XS08JQ
UHZT9pr0Zafr1yevURSJoTWezqKgViX7cVUPOaAXIF0DjxWt2yjDsFDd9+yV
5xnuNXB/EUtlUw+fCQJhC9Ncd57CZvxhCcxQXY3Gnah4a7xa9GKYuplmIJ8Y
sHNosf0PlBOVzuTFxtUWEgqh1MARJK/jcPFTWEI5mGu6bLrL/999pWXFFEFV
oP0SfwJRcsTHRkSh7RYkEalpwU9e6DHuJdQvlv5p5Mb2/Xhv9ceGGaFzwW2h
v4uy2K/tfoTl8Rsbs9FsGCOYQeQWzDN9tPq1VnRd4ULcWUL+QGtV+iZPOXpP
SFSTkzbBQ/Zv1EfkWtz1wMmE305Zy0JsFmlAe48i48DNGqaWYVbmm7laSSGV
qJXCr37rdtQnv5+ORt4f/pkpLvwakpB8R+fmtosqcgxQVlfQSYMtPUp21Fd+
h9ul4FnB/8cRLvB+RFgofwMZo0+pg7JQnFh/N69FizbgOmw0Rt16AIGwxUcD
wDEzgZUNekkKexn2j/3S1yHanBdDcA1LMCjqAA/WB366sxKvjPHjXbACubRg
+gLjTR3uRBBNKHXkXirntA7ffLKsKX6aq9MhFb1PH5hZ0JPNa9fyT77yWYLx
muHuWmU6LGd8ep2HP40+mK1adfQtvhqCEwjET3TUtzRXIZO7Z7gk5gkxKWKj
MSiFs6GU2d6z5u+b+6uzYAne9ykSeUzbZ4WPWlsRQkcvWW/MGagCy+O3JYJY
xdOSpfp0rbJCIlW41mnLAaQFNwtrm1TEm2+xmU1gEHbbRKj6ykV2FIT+jmR7
eTH1zYUZ0dAYOKIp0LUaMtuqVa/uc4jzm3ga/uyOHzS5Y++GnyBRIgfXAMHT
dwZDCPladFo7WSlYmERIEvLIroLtBnT2BcmQQRFTQ12S1TzH7K8M0sap86RL
22iqZCM89zUdFeNlkjXBmnTJIswdg/R3jn9L13UGr6rsa2PNlsvjYmu9Z9sg
g6hiLlLpCmrqyBW0IsqJp3GNCwbYALMdgLSBh32Haveya23v7IoIIFTeWtlg
BQHkHoEJwRPZ3GgPfko+x20dkebC0h57WM4E86PcszhGpETFUwcFxOKzY90A
teSOLMqydocnlO5XESz/hkJXTLuhkDrTt/FVhKfhPmFgreRuQmyqw8zjxigW
ToyS0hXWkPYjwV9s66DiMhy43r41cYhXcbZ76i9BHfQhvyDWj7kkNc0UdxMg
LnKtxlVXUu0Y/vcQSiUr7ZHSun3zXDE2TCMk4iIiru2otWpIE40xLyWq/5gg
iU8DKywpXgNYpTKXLjblDv5FdKQLvY5McagyYFaAvz1x41uD8CVpmKyRQrF+
lgqd45nGRRJ6+zwf+1WHuKOdMNX8k/3SFMSPJOKkAtDitMCbCfDFhpFwAF2l
cKKQ2uINKIZWgSVaEV2UdH+zw4/fEuvNfsgdQku1xmGeKgL414DGOVlA+Wep
wBxayl5XoHtzDRAPlzvAoeig9CFFII13grld/VY+s6EXQypU+h7DCWSrsCUi
ev2oRVHzGGENeWjW5T94kV6bUkhfUvQdfuUf9RlDMvm3A51JZQys0/u7dSox
ZRhcRAhnGmYy9McVkmuNbRgZA7ypQtu9lAfBJd/ZMD/MwV6Hnf7IDuAk415A
2oYlSgMxXA1XUHICzXqYfdrD5A1zAgFQz/Z6HgkoBaJ9TdbFua99T1hLGgsM
ETacoQNqd1oOkrkUn0HWRRqfaWq2T/YBGfndjv/2oHb66aKcJWavP/MFK9kc
/OF3gu13FNXvgXsZBmIhV0AGGQcw3cbsgDalj95oOMb0PbrqkxxAmo8gSlGi
+LpwVwtkztzxljLmMZ0E3f150LnHpUOZVm+7QDErml92xI27iw2rKECKmzXl
Et7+7h/NK6ffZTNsDsaoXZQWJMuW02ZDufvIahA0+uxKvo4iTQli7i18v1O4
MDGZDBWgw/2e+nolbnkwaaH3cTooJjagSQfQ4AfMS9t5qEIa0ApoqMOOgWPV
uWt9ajoqQLI4Uloh7RbbIMZc2ibcL0rB26nGl1jiysy4k9wQHwQ9OUJNzm7H
zoB9h+dJH/rbpmy5eCBYq9Wzwzt+hsrCPXP/kw4f5xDEeF3FwF8XjYzZDySz
s5VCO5Q13yc3g4H925JMK7YP8mg8PLcei7N65smx7PPpelhlVvy8yd3TcuE5
rAq/uKDVgTjR07V/Xs5wcY3C3/T9/d9Ja6UGrVeYuEa7EBIon+MPJUJ7RoGL
l9+W08jCMorUnCjrD0FOa2RWd193dSUj3vm0qeSpKeqlZ5x5yKHmocAxTTKq
QcWHb8GCK4oMRM4NCvUUA4DHK4/OAdUoYEwhorW8o9+uuuLmDQX8hj7sn1MS
/c85avFoLfpirgLfnGB4SluigySmCPruWDDz6OZOO/DeD/01Kg/kVs5Nv11+
kgF44XPzqiX/LgbeKIlAPbWaX3Rji2k9DnldYwIGETMPhg/ZjovgeEe0zYZ4
R7gs3IJixApKGzVSP6BDzPovwbBkWjCUp2rsa507Exy0jva+rOE22EGluYF7
0F2YkRGw4ynmjI2I172H/NVwEQ0AeUO1MQQ/YiMW26dRV3LuYtqswOEAs2+p
XvCzXqerVm4aczQ9YPB97jfg6bmgn6hVQlUBSPtNW+WUdYzulrJ9S6Mm/jCq
KassV3o7DQUVaPu5D06M4AS/UvFtmnnWEWbLPH7BvOYrpBj+1MoSHzij7R91
S1mzo3OHjynluyknnVdMsYk3qGFQ4Rzuos4OnMrVEf6gtexkwjnvreq6P62i
i1CJN7u2VCuNR9RB10MgN9411WWN4GV6v696g0klhwVnAtSiW9xOfY8UhMV+
+Pl3dorZ1wroGSOaiSwSHH0NOvYmJ4RFYALRdoE5e/lHVqrfjIM7ti58uQ9P
pLokR31SuIvMBCgYuOsPV7x6mjR0TR8yaJlYuiBmRYXJ2DnLszSaC8do+yZ2
5UIZFj8ADGQX83bFz92UIvLQKDWtMJ39hd7zslf6H2x/MLNgm3BGAUykC5br
/WOPEHAINI4Sre+ylLRaEMEy5UioIZ72IcgJNB11iXZrLLgflYpCkZDVLGmt
yxpkWv1juIid2086yBQHjGikK+Wy33bJje2MbLtDLiJfnEf+lEM2YEu6/UCo
esPahXOMDSmcwhJasc5w6TrSZNc3SVwZtECCb616C+hSSmuUkxEMGOQGvZUN
uHbo0cK3k1QCJdBlaE1Oqc0vjIdqzV7DopFtOoZyNPTuFuIty3fyBg/g/nFp
9PnEUBrpG7F4CafK10ogh7O2fcrsumpVofU8bY1GfboxXGDj4GkQUPCFsJfo
KCPP9wgQupx5FOQVuSu0GUENHV3CF7Vx+Zsx79n1qKmaGI2y5NhFHbrgghQB
w9BN6vfzrxjFpg6wMFCuGXpX68cmBo6Ake9i4RZfu/dKUVpJ5kzHo3KMN0GI
FSlEpf9ODJVcTU8VyZNdQs6W1aJQafURh/FsjauP/Mbd/WR/TmkDfd/foVqT
1TuW0/XjUwPjXoLVvyMpIEvAuvART9KC46NlTPC2xA9L0EGGYCz9LYhePdmD
8gGwsv0ZUcm07NruzOpM125yfKR7SymEq0sx5VhGy9Rs+GHixn54v3j1ZknN
RWvYBkezCnAYBJIc8BEnOlZ1rBvybDRdZsPIw/JeiuG0et1s1bEybh2VdcV4
KRNn6eITF6OJKCPKapjcquSZP8eTKyixKXO4AZhK6K8OW4AreGPC37FFW96C
yL/Q5tyo9NM1j+h+masJ42F+6XDCIilIC+EOOe1wpD7T23zPXZ2cBZ3O9HLk
UyM99hBAzyljABWBCR6PyrlwhZfpRPnpibFJCOgwmwIEV7Ibkk4xVE5RL5/0
njtlTGTgy51TUVTMmgdBXe5q1M0K9qgYRd+r1Uff9WBk2YQ3jHNK6q0iidll
Uoq9ozoxA7+ydEnScLfRwhJd+f+XfG9E5LpT8hvo0vXLUw9Jk/EyOj47HRV2
AN9KJZ5mEHQbZxTdpLkTvOaUe+SWYWWW9gqeMS9yKK89qUQLhacgkFfDPcME
5zjIiNYmqbC86TvCGCxzHKZMrkZHYrlj6FPcVEZ5/d5v/i4op9QI4f+WvJRc
iUDGItyTy7xZ3uAvSER8qJQuSFgaYmyjIXtJI7wQtqfJzNSBwb5xnZmveSfW
M6sucqqKU/ZQJS2MZNqUz/tB6N/w7/ozUOBQVyezZzsbZ4/3xe+8vBhnKvPr
eoBZ4xOHgTSqmp2N+YcOfSgbKov6RNUolY7gwaAkMMfTop+9gq9y0DXm6Gjo
Y2e9NaAjFA9uSUgV9/JoaKsrlCbQwhPTzx463EiCEEcXpTU/jh143IL7RSI/
k5jCXgvD4bV2HBrQN/A2/03vohUrvJbDamlQXRrWf6gwPt8i5bdK5/YnKNjk
fg2XFAmS6YIpCYvSmbVXtgAW0C3JEu8iQj4QmA5hoSFrdlshYgOg0DQulSVt
gtYkCEXGL3FuLEUfOtjV3xyR6WHb/2RAocEftrh9Da7gRIq8pb0dOdWw8ckg
DYsanXTJJlLbcjU1CmpJYL1DqMu4sha9oghy+eYaBkL2RTIbIzWfkn9HPyjO
r8t3ABWeiimHnboST8J+Fa5rvRV5MfcgAeTvR6tXuJHE9Kl6lwmnrmgX+FB8
Pz4LJTtmeqXB0gE3hfVrhDj0HAo3+bIJ+CYRTnLUmtDp8KcgZSjGLMNFEO8P
D8HK2NmBFsYWxUYXg35fv5SAfSrcff7h/ZeCvEbI4OoQ3BCqd1oHjvSXOJbn
3SPmfvvah1pL4qK/IuNrynoWo8idD7ZC0K/NdDdJyhWWs3jbiQkmezkxda1p
RYKMMwSONF4zjwBcDKkKeYwSWi1x666iiI8z/w4T6IzT2qFOk0e41w6inw8Y
KJ433EzHORMyvf9I1bSNOUx5OFbh7oA82YBYzFzKafAyhD1KQNnrUmcGwqkH
aGFNXxIppNjrbdAGc24CdenrqWutp6bu5B2Bc4dEbPrJlAa1yhnRbHtmZ6e9
5iUgcmaJDqyiJdaDANQf/ktLdeAHoyj2Wq+hhCxpcuv4AnsVQe6/2lPAEiD6
Cnz1dJ0pl4NH1EQezThajTsU6yFqEZg6N5ZlabQ+eBrYjxpHZTnu9gOSYioL
Zrxu7XKiCV9Qt8sivVNKu9JRO12ltnMjIH6678o1uWlpfRTGj4Hv3sxjhv/H
zitXAHk27JZ5e+KMB5QEiusyL9digR0Bd07hB72HFGgv3DDpMLDM1VY84LCj
quIpzm0ZaqkhxoXTAo1+sQGd1J6lbGNCYHYFqypeuNXieplF4dgMBAmF3ks0
fNfPEMJldiJK/D8M38bwXfj95AjRaGDrQh56xfCfbZsoeDnR5VjDMeb6I7jw
1E9vX5fDIklMWHjSotloHHDFzxPIabegVS1picQGzpXodoQfHQDE0yUKQS1G
DVAKT2/Wp/XvZ9ioul5WTgZIaWbKws+gymI5B5YxgzghwqnmqX/SYbERHs0J
6ynswaRA31niex8A4/ydcmphfXrxnjRMPfuKUNnP9gRLsuSCws5MQhN5issA
ruf1UxGB/N2VCAX20cIuJ5AVZCpN57oYOnlZAgXpwz1E4PkoZJHJ9rlm9XQj
m8yANP/FY2rVaXrlKZ1A5WDmQYz6hOLJfrS3dHc77l5EiSLjhER7HLSc3UY5
GWIqGuOqDNmuBec+0YSp9A7dcrHL99t17ztx1g6JHIrj6qHkofYsG0VC+ull
/qg7SSdtzEinDb4awF+KUTMHr45+dbbcXF533FiKwnoJsYx/y8cH8TIz7Bku
Yz4aYG5u4abog9g5UM6/wZDO/cB7uBMhntQ1Iznh+eKhWpQEXHuqjMsH7U74
pVOixXpTIi32qeOfmKDnLxt+6JdrmrFFf+KDyd4ux56/mFfHSItiCHb2xXik
QLL1tHOKQjpj7pv9CnLZfiQthlshQ+yM06DBAzKPYoRboUXgLVa6nG2CuZPr
zXyaNe+u7WmqzQtRjjZvBwxC/1s1J00vQgKN+QZsn6tRtVwDpWlJLgXj/6KK
8IRKWRee+vQivMqYUaisnDNULp/8uGELze0g5vpf/LN1g5rteGFdvRZVLwpF
oaW4U5zQ8m+tIskyvlGotxt/VUXM86wU1vLyQp5n7jzS5qsKMd0isI00khlM
TQ4Kam682zZQ60EC65bMw9rhU4LK7tqPy3kyb89A0dIUm9Z98Ms+gIzAGWUJ
2pPHJa4cGNmWqDyotXx5qqoR18YRfMQLr6cw5GlSpOLZuUuaIntirh301Mrd
ikAiLlBHVZjTN/ZrCp/gbEKBCVk0LM0DOpYiBxYt+eniwzB5GcPaeK6QPSQD
/gChBpsXnpqC4wRW8UZRBj6b4SPDttAfp9xw7AoRkXr8lF09zU48IWSaF+oU
mPlFJiDn3/JJCgcWM0cBALYbeQ/GrnovJGpcm7i3dq4FvwvHSTLzG8TaE8s/
TZtYw9DHbXOdxBtvsyFWknctVDCso6Jqpwyol9ifadzcexr3MKxCVB1mifTz
LA+Ioh/c0uN5eD6MmE8o7O2t7xWb0LwF/vMk/iVp/T1/z7+xj8hTsUY5uiLK
FLQ5LiVTawKtck0WF/8oURTO5uJnHqbqG7UMnwNfREXhZiqpWnkWX7z5zXG8
NsgPuRq+DKysKa7gN4yILN7kTLQu3KqiH0GfrBQk2FrIoDd41dphBw9aFVT4
Z+DU08zEAam8TZs74bkWV7NEGzSvwNDf4ixE0QDnTrE4QA3mK5j+oNhVp+NB
N7R1JyMMZJ9gmatyym+T14pBimHGv50SKIC4xHVDn0OK7EPM9RoVIEffQZyu
keEr247KmWvM27tlCZJ57Ez31ntWRXXr8kNyxgBwwdmwUc0UEv0DBJ0l7cli
uE1pTmSljADTaSPAjmMPWRapX0u0a1EkKmn7VKLooma9NUAv/8eTIliCitED
CYjxuqQ8967mK7cvdAXgvST8+wuBY6CoDnauNWQqkKylK/3VDYM8E1+TO7Vg
CsjOX6Ift4bRkWUSOy6AD9H1B8Ofns6p91vhVm6oQTCRkP8brvHQV/d2+dqj
f4hDOu22vRIJChe+UFnoR4LwXQ6jd5AYTYNbTS+c0Px1E8ozOw0fuCiILUbk
R9zsx6CSHOM1ku13IFtNUcDZM/RStDEV0kCrcqdXWJOwtKQDFlkdoi8FWXYW
qQ1JHujwse6VTGXQ9ewD+PQ3rLW5X/eEQiq3cTVUrYi/hndTEExktsSXyd5a
UU5FDz3mmcaJJyU9ggv43IsPb1CD07KclKN7GdnlQlqOvtpuvfNBidBsTDjd
12CUJ3xxTNZ/8cmQUQQ5uSN3pcb8BUE+RJ7BQLosnt0bhlhMo4CDrG2Nvs+m
Jpj+1nrDdex2Bql4mksZ5X5VOIJOdgnxX5R9Inibzwxo4pB8JY6Ca10laOX3
9fZe6zCl1/s7v4wdRCl/oEQvfJNF0R3EkRq1Xq9a2R4E125+R3IC4PbXlucP
qwvu+ySmOs1F8XE5CSJ802c08xzQVnv/jABLRzNp/l25wtpPvIwKw9Soyp0c
zKS1MCIy8D/im8q/KCHEcfjY+qPUJxpv37oVQllkiqY8P7FNEzSMs3L3oimT
HGo15vl80FC1yMxmAATT9f+DcQO60XnF/ksfNJRmfPoSbtEvA28C7/4sQ8B7
b+ytUfkWR4e/Sbszkq4Lpg4Qzmv4CqoQuwCvvH/j8tvids01ExFdGXD60hSC
YtM77RnoUWyo6wJFoowLmqdPxIwYjrnJsuU+KR+y1iVxuM+EMm01icVFRrqD
LC6R2CAtBUgHEg/RsSlhu4ydKPn5JzNVFcA/84gY7oGCZmlOxThFZGu9+myL
BfeRfdJotvqb1FpoEV70PK7BFem8xznUI8zMhJhVMRImt2ZkOd0+9k81TXAp
UypaR+EpjgK+vGeqCVoAaZDZhMx3CbF+wn2Fw8789KS2/2FWPLx9yo2S2q3o
x/O4EuORqwdAnAxaP5cQoz82xhZh7e3T4C9gE9ZMFbd+gfUGRhmPcG7WO7wA
REnEpnZrY62jAydYpFcoZpgDIVXfCKnQNAKMpRjOsDPQYxatnSkIx8vSYGLQ
2/xHl3Y/0sVCysIVc40aVafwKI3EuVMsj42Mp5kFm5unRbhwHHzjMMDD6Wov
wNL4AFHweZtS9G5Fx0PgnW0RI+9ZZ9AFHez5DPBiFAr55ktcf4hIzN+fPf5f
Ypw0jA1ARNn+yvjEp4aZ9+SkRFka1KMJiGU66wCOqIKvGnlQU9C1wdJeryK6
+ZmDPEsdXYhcEkRPI3K+/Q9YB2npdk8nynxfHc4WNmw9/pZp+s2VijHhFXfP
ltj30yg+kT701Z/qc+53VSvEAQVHo24Lll+n1W+ItbkA9MpcvI4vYhOYgKPA
5NfPRsZoDr3h49kXINGC115OQ4t2Jw9DXJOhhWsFRVg6ckl1z0y2bLTofTH9
RleOsyS48tm5jZ57xDTJhdPPanIoYav/Hdw4kXOSnm4i9G0HIAtNCoAph/Ux
06q9qhsfXm4zQLKaXhz8O9yY0Hs/osAZ7DnNrlnBo90qKbAsh/VX7+Br0JQ9
y8H3sObH2/RHu9JsbxbG7aegxiuLaF7ibArB/snDZv3KpOKYQTa/ym0iKmZZ
9QEiPwZ47ON6AASDl8CgoPR1+DXoblgBi5pYRK3ZHbSVHYOUinNe0y+vc0hu
tgkXy3QLcBwpF2jVrjHlnl+nLT+L/ok6g3pyYM5rGZY7vVeLAimJi3DzYBMk
7bLjKPlynjDodqwrS9HRF2BiUulPIjX39n16A6gpDfvEiXk9DvvWEVwWeGO/
aT0fNiAxHICDm7pcr0yUKMXM0G8yetkA2UshYYS7lLeLIWDqwj6EQjj1eLS9
FONQ9digM6QZZpGLT0pqJe2E4KixaGKGCJkcNlg+t7Fj0c8BD91g6QoxcPPh
cIx8RkRjaIbJTJWlt7/54EOOuXw7PKUgTYO1Ulazd0tbAuoCqoUfPxXD0gCA
HAhznd92PW+Y/coJQrPc4ifv44peVqvFC/x1QcQkJBSPNfgPbPlI2JEYNj53
ux7J/aaOzgpOvVxATej5GlrNW5DV8wbvWpT/6b101/ad1EHkoLDR/589pXlZ
LfWZs4Zv9EsPeH83WfyUI1ARm9UUF49mYhP7F58IKbQrYR/COJgUG0pB9vS+
ciz7k4wRVjwwzppHZWIP1DSEkgnqyQ/qzsDLu8QhCF5Hjo2B5bmiu2PdCBqX
yhzotsmsUfnKtznivJjeWxDCgUTiR77r8+Yyw7pNKRo/zseXJfDTRTWFJxpz
Gs5xZD1LLe/nZxLG+v6briYbBn9QuxO/QuTmtMrRAwZLQjjiZR+YO4bC71oJ
438GJXhsk2aJfBH/7Tt8tHLX0QG+xMgS77M2Pivr6JVThx4gucFqOqk8ybLG
+E6huJonVcyMaSUX8/jfu9dKdnW0wo4qKeD6JOItK8256a+eaol6pXSwL5dM
bZOtwEoBD8L3eMLG0SiQoiEbESAuvCSen4ewG5wWJu4tbu3820Gux7L7T8sk
AkbI3dBS+RUcGXwcePBLmfDB9cTGWiL+aTvUTCF1+GtpSWpjc2S9Jc3mku96
NkEJhLxKn5ajmIWFS4rOOIFjYo0Dfs/jJTB91MSsmDGCVYxUsyeXC5ypfl4G
IUGPBhAycqKaNRo7KxpC/jlXoKe/QTyZi9MmTL4djs2E48qRHrsSebptPE4z
jGnSop6fSa5VUgdUc98YbeFhbfAuRtL4vHg2Ar2AHjbmNxc4D41wldhnbgXz
o/xNNW64D02thJX720aNJbknofjo+8PJetqF7nzHA7DGAKp8mUWGI/7j7+QJ
KxTeFkK+mchNnw2dFd8CRZYCEH5UAsh2jT+oq1r/+L+PhTDLP0r5kcENNmqx
ajpR+cnHoQCLtQ2SClw9IVDjFuVcVgVW1XxbS6Uhfke8rIXBJsAXSQCGkjhF
5BmT1zmEY17U9JocPhfDoWFSc9euXKFx7USHRnjIkgx4buxplwhYu6BnRcPV
8vyYbr1wGZzopcF9Ef6KSwoucizE3buutgYrDbD9t1T+3kthYivbzbTDrSW1
nIym3MA+VxzZDzoYNkGUlsjtSoOXm1rlpmx9PE3i+fZAggHyAsvXMCcslc03
4jlxj1TTvgpGkv07yknQWPKNiLb2E6Fg75rwisAoBjTjv3BjOMgq2Dkv64oe
3wMbMMEXP8yh3+94Y5ul3zh4rJvOhImsh/iVd6m+G0tyDcBE/lAtBGhhHJny
h2NRG7HqoOnL1i013GTg6UakqbYBWIOQZFjE1NJneV1wUgEmlSHBv2CtwjkD
k+WKfBLbgIuaWhgHhSd3vF5ambpwg6OnzkGtqc07I8Hagbsw9JxOGrfuKxCh
lhungJToWs0AOaZ2VeN7DPOxZUU1aS/4qt8ShnG1bvDjv0h9xoIFBpPw6dLD
qYPS+j9vxrW1V3vtuStfb5bFJ2X5ncQQD/U++dec4uI8suBTbSQVSaOfK71h
IHoNwk00NOQn+qwD3UYN4fBu7nGo+9KBxxiwkt94hMGTq+fcwp3LeQ9OqLT/
8EjTgttevTBav1FV2SQam+1kvGD8Fh8/I7PNNcl8ZI3lxkXBiCxzrOw5rq6Z
5g7iqd+ftmF2+KNTeJJCwI1rR4GjF9//vAJj6jkiI0TphYeA0qgnfCDIOlio
vlSpv1x91XYLEp6VMS2GsLeXhg5DN2D7YS/aw1R7UQwkxQyJrbWWQV8dvTwu
S1De6BBZRigXK3NNb82pNT5iYO5DuBORksox9OW4KsXYQEX77bPuQ1S505ax
yi2NhTO+bBbNfHKCdnr5ZgWXYZgMl3wxxw1atUCmHFPvM4PLrl77McePPCcV
RWBqLMD3o0nXwL3z/a7lmWaoNe5qDT1JrvOuLdahg9yKX3t2N4x06cp4czqy
1UUQw7NAF/b1IZr/t8z/o6od7UQ/KWsmdSxeuwc6EyrPydjBkKsCfsxnrt3N
P6jjxdBFnJJER9U3q19KCY+N56k6iy5M3KwjTRm+M/+goLJwGn0SMT/NLcmm
IcrA4Dxr95xbyaeeE+0WXA4/bnim4RcRgIkUhBRNYNxPx5Xlre7zNXPpGzEY
0QvgspBQiz+nTP0ASxUMGtu+hBoXNUr5F49zdfZzvuRfyj3zhPe8s5eF3N/i
xwcJUfsDc+rltlMnVwDw2Ui/Px7UPiz06g9KJqj4nuW7xekAZ4KqekpeZzLS
edWiMg2BsjJK61iIStm3DepxAN91f4oUVFwLmzU5X1t2hwsFagN4LuYrgfLP
wH8RmRNIItJO9uWiGOCK1lF8R8eN3Ip90bLHQtHvlj39cuq+PztsA9GM9OWS
YbhzAhV5JFb3IZ3RRWGlI2kK0M/GBTDBl1xrQbFXRZkVQzDivJaD8eTduZMY
PyWzfkjQA5LCvE9yKBJZm2STdEvAjKVwuIZDQq/i2kg2Me/yO1Ko2VM75t9X
Tn0+8c78jPkzzbDQne4D7U2WoFj1XuEnNt+eZBxf6ETPK0+yZc4GPc4spxrt
GuqPBcLZGPTy6USBQ0BlCm9n1HcQhZH01l0LIojIg5oSXzQ3dSbPguyRhiEO
FduV48CwNOW+XEraR/ePQXN9Mwq67TBW9IRX2HlwnUw2SJDHDEQj42vMpi7+
wTNaACbk2WPZ5yu9aQr72cX7Ta8AmACGlDX5cHv/QsQSVFXcXY0TEa8PmWxh
56kB9mI656DxAuBBj17RPyoYIuCgxNeRKmaExPZ7I4/byL3ImCy620qoFumu
mcvSfhMfcRBKCtlObhgE3sH7Og/zvUD3wXN+MxDxD5QrRLX3aXZXwdfclbZt
PsDi1APBs4aXX7h7UMEpkrBwoC4YvdsgZWb+MFrrdEKG+Cg9z5RjUyw1dWML
H/FQe9XokQqJnB/mKjNqbqCmcXNYbrCFEr8xciECvk2bGkdmF/lQ7uJl4OVu
Lqw0mHjPBpEA1bo9L1AXT3F+jzVBZj4UvpvwgjSQ/Zn4e0idLh1W8S8bsgN1
IH48rxlNz3s7EQ7If8yiea8AHf5SdL4eUaEPxP8dEKdZqBQEdigR1Dknx0ja
UuKtcaogY3TCoBagM9uiA/D4IykUb2CE4/j1A3PlZ2tY1GFNfHOnGvsX8A4i
yzV0tTWnXqjb3IJaViyyj6qA/J2+4z9YhSttcTBU9E1ngXk2/df7DibwfVTz
yPbsICi0/14bLdzr8cf+Z4qHv2UQZBenzgRRa/i9iBFFQ54xfnSj6/K3Cc09
5tFx/iOE6UA0gVkFB+JVgXo3yRszYqUqrUySmGsbXqbcgskBnOBCLJn4PQpq
GJQ2z9XfD7dK3y5CNwvemdPnDtXp3RN2NX/YZdShzhxFKKSXHN2pBopRYSKj
9ZB2JxYjLvm0jnIfZWg+C8dGY7r8Guo+V0WOJ6gcCkXKSzGKYeBqMRuh6B46
GkQlreKGFF+g6J95gY94NnLZl8KikDUZHxU44N2cE9NL9sdGdoW39qhLc7Jt
oiiIcLxGaC2mJdMJpAFC87wnKzUPCgWjgfG0U7eC+fPlH4BEAia6BJpKE7sc
jG3vQIyLAZBuYPr/gKh86p8gJy/U9a75RA/a7VIYMkZXoDpIEf1sAKDZ/BL3
xOKIVd8fq5RtvaREArdC5q71Gp2PBO6fSM+6ij3WGt2v2+RgFDdpmfHDxTb9
OT4ffSPbCL6lvS9+lz5VecJ8vNy1srb1R/hlbihjRUbt4s3O+yHJgmpMsQYM
WJdrEeJOItIvHNewgZGWnxf1F1ksEXPaiUGQoPocAO2LfYH4E1/nFnXDWM2a
fdy+6io8p0mRGHYGaUYMwVCNrLvP/2Mi6DLlaZu5y4Kfft6OCQP6clc1w3Sp
BScH/XGUG6KVczN6m6Xg5AWCippGC6/w89pyTNEVVvL9aR47CJRRcyKEhUIQ
Eet7xzKgG4wXhGWvJIkqx8VjaoIkEIX9hiF0boMC7td1hRoAfYp4oKB0Q6V9
nZNlAaKSO36/DQQqtNga92rVnLu/jpcsdXHf3Dcqja3BvLwwNfEp5jA/aImN
267Bi7N5frTFeNiMwYvN6iCPELhylm0Hvx73EBCW+Vb+gAkTJTyJDUTfs7tE
zAHgZUifPTnkz/E1O0bnlTuvsaiov8LDYEHdqpe1dKRmJpKt+5xPU/8hdmJA
5WyiNxFtVK3+lnIqupeNzlRA+ep25prSPXjcOiIwTRF8IiSXu2U4lv2+DWu6
QMonxwBshQ4Rh3ofVRAxyY21Y9ODoZe6vTgrrybqKREzahrv7xcrmezw5E6S
v1cdcL1/PlWYbpj6XG6isrliNPJ775zJI2JwIc27dL9NZxOvNhKHWGl6YRf3
6uwQT00Xde8iTI7qY8sovmQxjyI4zdez5ba68xzzg2a/8+Pthm9mNMZZw+Pl
NGCWJaYnGB2FU7N8QdEcehRXjWdCCBsiFkajSN822J1ykdYIUyEh+vSRv8Fv
a3+WL6z7Ap5ZPRwnFFRTanuojnv9nx1zvpwsQKpq25BhucMW7CkcPMcwvgWv
GYNKeLeoLp7rP/cIkFVWYcyNidlhloXg6eva4S82hh5+5dj5RAJWr9SNYDAa
kWeNmV9Yn+DjhNitHMXg4wG7BNG7r0Cn7is0NHcEl0KlyOMIf8DmTFaWfCQt
z0zJMyf0M0tjNx4EUsZF5XKRvBv78mq4WeGNCStSiIKHa91Sx0ko2uhdVmF0
yrfHKAaysNiH5IhkMMwgVVjqI5+ukvU7N6PB1d5Pv/2u71IxQG74I+MpsEDu
7MmNk9dYA4yiSsofo8XYP0pvGwe5fUUfsmX68TnvNGXSbAnLsgFw8Fzqi0yP
15RXoMFHTG4BquITFeZaOpVXnLDTu2kDdfUnABzXUWSdDTwRiyq0Y79AN4GC
W89K+cl1imbFGOb2fcKYo1hkTY+LnVUGZOOpKiFilK4dIyvKb3OByrquFcNM
2UhoiVv+odrA1CYoZ3n0JYQAX6asbFK1++TLQa1DwMX/+LTf/33pDn526o+/
fB7KjB+1W0NBvcd5MwOPrnMZ4l7SkaOg5KN4iVQLO5KNeM4JdSM8u5lP1ytd
kkQ+9QGsCZ4k0MPLYzq5Fv2d2nFUMRp14F3Lu8iIP5+lW7m19sOCMY3+fIA9
orwr/Ic52ahd+fa2NuNHm5WYWTQULcSsOrEiiTIAQN7Sfep2+sQkHVJTHyI0
DBMxoYijZfZQ1S6dkwN8rxbpWFFvTMLvnRtQTZ4FsObKice4lfY/ioYKuAXF
II9ypeK4pP3LVcc1JmKGjvNQ3zMWPArr5AdUn5wm0D8rK1ckHHFNvvmQB/qN
0btIbFXykqiJDA7tsCqsqU7WfKq3DsJ+8fAQ3a2eL0dSNLsW0mq22/esgNVj
d7UAEH9q6g4DmuPP27KA2T8tgsjfy95pBfjDzTZYKIYP5r4QVcFTKa5udJY9
uU0UJEgjjodPQE7sWECTsKf1hbWVYbHfmi3kf3PHM0skli0LoPVex/kdN6uy
ObPIFuDRS+1TsQo5PocKSTdt36B6nVPmiv9Zx5IjzabEOq10dcB2ltVLtVjP
hicoeLv6RtUDpjT1Qb5+MCFIM7QfO6cFwEpZF/4PTg6bF1txX6OeUn1/nF3P
6ZBYxr102vvK4ySI6VsbqEL5tZaNptz+RVoLMBh6Hu6ybQ6XGpRRHPSpVEGz
DGhimKLrhVfhHChBR7G5nHeiGTczmQ/41/XTPAcUkNa2isNH8SCIn3nn5YwH
anosAj+tN0NoYqtJkvszrCz0tt8hFsgv5mJhVnjvarGaLnk2ohTSYOdpNliE
3dcCH2kkxVUxN/aDwPXinUeucPeUlSJrkbkoczpZBUazpnqTxA0igup0wKjf
Qqh4/MwHkxo8F8taP2hIchUdL4NW+U27EicYFwkIaLIgKsDHBLEoU54KrpaF
wonp6HttEizfD0bOICMXrp7K2aBpY1GeYquuC6TCyT2xYJzKMGjD1UPfoNvr
qmxPMR6Md+EfLWaZO0iYSNZyrjkQzd8dxL1UGhPE6tp8DDljBfANLj3Nt79z
J6HHs+akWXUy6WLNnIjXzejzCj6aOlBTcdXWvnN+DtdjNpsfS13EulM0eF2c
okwvlFDk5byhRPyo+rsfbI8PcW/qGTscXvhC1jPmq7wD3lHvsIhQbYgFIFK1
ISs4fcZ+MdImdKgbtKijHOahIyQPSQwAlkO+NI1foNBi+7GsyiuBzr7VKrG2
C0YFqy1gfqy6cxqejkUBS2O9L5cEN2iwrzb5uPJrNk3dP90FSomh8D8ZM6Kn
idO786rGZtZCq8ly294QdAAbxFksmY7M7ZPwLfyUuxnaWjvUAAN5gBtiRKvh
4t3j0c3qZiyNmITg+HNJNHIW0wj1rncjzKL+00ZYAEgrfIZ1nYIL2b6GTvkw
rM29khmspIuaEY22z+inNbdAWGg2oQKKqd90nkcxBTr13kAg5IvteHfQtODO
5+/JGO9SGMWHCkJQkpTh6rx7/XfDTluDa8HPnn1/BjL6Wo5VN39H62xjIFYN
4d6D0R5RuG+awJWtnlaA2Ss0da2/uMalfkSdK36xtiS28hwTOq8T7LdXmGwt
6WyljN8GAlTZkjSqdbrYsUIaWIXvHA+HWcW9yfwoReUyoWmqJmLHY1gXEBnc
HtnKBfkD1y+7L4jbhw7CzLflSYjW26QeJly6EsbJ9y1AA+npgNDJq3ZUP+LS
5nBEL6Ok4VuTMk0jj1PCp/4gOAcGsiJaLb119yV0bILsMCju72u5HLNcf3SW
0d8DKRH7jsW2uApWZ1qayA1R7qzIRrDowOa4pW6eHLQJGqro0337Edc27BYP
sQ4zouIlGCHvi5M/LZaXVcPkRvLMc9xjUx++l0uF6/EPMd7SrZH7WfRXK1C1
jTcFhTnPVypILdkOXURHQ79RKrPkHqQRyB982pLuslddXU8kb6g1vdvuXHud
APjwQnIOY1mrZl19KAzbfFy/+P8jSE/NGyR7hKfVMstx0Xp3dsL562iSkT4q
WVeOQx5v5l/Npg2uUyDLs5lSCmC8tru9DzFzDGhubmuegBjY1J7umsqG0zOX
zsFu6LXRll211wObdRlAkPq9AnChpo4XqVJ6k+M1s8dY6GaBHUvTnsD+i78X
/5LpKaTz0R4PjUgCU7jPtGxUsp1HET7+qEI2e9M2LHWwUFB4yoTRfPkIzi0+
t9I13kniRquHP+9n2xLi0zxrAKxa9eVcriQFoQ8aOCxCgo3SdmUkLk5DfMDf
CLCRcbb+c68S3YCDOjC4c24aWQp3ckQ0lj0T676ywcD7xRxPcqiDIfwigemG
Z2ydka/9F6kLQ7kVui7BuMMKtTQ2SKsSbS+YD0jq8BwzGKnh5etXlZxuIsDd
2O9RmwhVUaUXAuFiAcj1YcTzU52BbmL6ac7pLcBmwzMLPoURXZ6phj+Li+Oa
KID4XuauAMSn9Ix7o47mK/A3zGyhO3psokTFeTqJ0/LuxwufxUstnQrNOY9z
MfCEXJYlPsamEEf2iiTU1HB+YJnFW//G91ZweTroPYDJi2vP5UcPweisfXJj
z/DMgdKK9iMqMCLIJZ6HR6uQUZfo3QAabiZezxngrzl0wzWeJJafqouhaAA+
DNSSq7WDxlbDroBjzWxSmGDA9JV1nGdoc/8dUeoo3NgRX1tfVpjb5OD5h3n/
RpkEr/txbRW9itE5YehBY3We79XBsm5wbZ6jZAVHNsQsMtjrMyZ5IctPrv/i
o4XcsEmLmv4p/lxUIsVFj54Uf/cpv1Z2fkXJNRwnzq64nmXxfLB62ul8j+Nr
mj6CBSU+Q1jYaIwLErZzQJp7nFCsS1NBDqzOTClbtYSaezkwZql938e9jK6X
nbduLOZ0jZptEM3wmYZtHv+U0AT7d7A7sYCkxPPWPFIu7SJEGy26SHTe8fe2
Sd8mA/YNpiV3kSx4RTG9YPAo9iqHswufpMm6EeCw04fzOFAJJdr3So13SlpC
clznQONR9vPOwFQF3KpAgbYUX+Skm2aIGhFnB9kgfUqvsfhK2zWDKV+53luS
QgIECDeBFzyqdWuf0hubiOA4q9MjTOI7MtsiCMkmbLaVZHFhLCRLLWILMe69
dkxFdCcCIEYAqH/VaTVsrQrTgawsnRmG8xSeHYetgpBKmYRidNBZ1DrPm1ps
cdYOrXFkhuGWYP5Vrv2oQc4sVU+e/fkOOnYSrQ3zGR1ivqHAyOkzIzP2AR60
7rVmGLvfR6wDaewKEv8yPwa+AbbGSASwpe+37w/hSM3EAgwwmrw2r5vOAGsP
IUUgWXLJGl1wwqlwKaE1ZOnEC7940VLZ6TsaUHf2C7/3WYs/ju0A05QAqXBL
SpVL74qZXYMm2poIzhQ6Sd7Pfk367NfKhu0Zn/rDRs6WL4pCVzSKQ9Qh5YMa
Q+7wwc3cZ2LR1TpHvxe0Ap9AQp6LJvA/ELBWICKiW222fizx0SyRc4yMKI/0
eLZPHMvV2M8ZWp2Q4DPlHx2rcvxK7izpuAdbrW7JDS0vd6u7CvnNWi3zPscG
bEbjysG0kIw4TjxvMPDnlM0R+RWyb3puw4gkq9lnCAYGwNJjnyPJ2yxN01Co
zFS4C/uS/uKIAuMXG8Iwsf87RzhRBakzAHRj0lMwbPu4hou/NPfU8wqf4WxP
ipjo4Y3GIbJTChIbZ2n05jAqo5rr0kXPaX/ZaqWqAbU1Sw7pzQAgj4LuS+km
A3VKCdM69+1RhUfkvM7zn6sSJvDe7wUs0CZ+kFuTjtHGIInXKApLE2Lbhp8g
b/Q5y1ZpU7/bFEQ5uxmk+ruFArKe+wtUOxZlLe1Bh4YmMxlVZ/pSdR1Xmo3Z
mbLlqMX8hFyWnmCPBC33Zt4iniv7WhIHIM4ykIYym2lurMZWu6W9Kpen4QeJ
qd+dCFdKbxXR9iYrdBGsKFkhTubawDINLg3W18SNLepoUIvHx0TltlBMhEtX
33czjeYI+EEBjbUbOdLY5eeRJKKg59IPVQ+1z2eiheMYFCQ4D29JFBAPR4In
MKCAGDbzooieNQBPJmXbbGFSevpRi157hTCSxOToGdxRqrH+PPSCu3qs60q7
5azVWzPaYGACXMoh3Hopz5P7jMibAeVE8dKjDJ3Ek+db4k+tdmRpC1u0uIe3
XUD6U38/HAHXgnjDto5JZp6CERHjBoPSdu+tGZF+0FH9z0ti7HWHU49CMN4p
dMPqhNEN7b4TDjcLfhpjO2anuebsb4Tgf5oJr36ty4p1uu39VxKIA2mRZgCd
/XUJrkfVN+4juG6fAP3KAE35Cxmpt7q5VIHsASJJ/X3fd3fTHNRmuREEwLf9
hsXU0Vgul4w8eT34QLFKsdJivCZ5U/U2HGsuo8JDTdsRZ3m58zBH+5UfK+dz
Y25uCuQD6mLq1+u9SMmXNIU4IMO2BlZI88pZINQDQyZzOC/j8vDq2utM0Cfp
Em8i69xnt9yEtyn9QXh0FOdLdf2aK8rNPg2RM+aLPN9nxNnOvStzpVso7p6Q
oGCdq37XHIbecHyiX082rqqxvnnFFPM4qAaccOV9Mj3w4IGMR1T8fc73N8Rc
3/tGj7SPaY+zSiO5ng4HSQZF/OgcnszTExYlYgYl6LIzvmbqjYj5BKc/ar0R
6zfR5nSO8xyJyFj7NHYv2xfZQT8T61mRJIjyP9Bl4/oPLt2gTtusVIOJ8sxK
WvO9pf75ZB8vGUKszeRadmdCO3q8Tf5hafnikYr/OCm0OQR+QhjMxT2cWyXb
2n/l0bcxQ1ez04LCC733nblFrrgSzvQ2L45VY6JBYr8iBKY3kWfusOOnb0w+
itsoyC0tUeAbVNAD4ax+0YKdtRyRZDIvIoLgp7xRTFUYAtW6aSTZOJLTwtjU
IvB/HCk0fADwtnsb+G4Z4QZ3qxqeReBGZeSYMrGfghs6yzbvv8a+sL8JP7iZ
7AU9+T84D9mr0T27Jaj2tpYRuAKkyHzmWXph9Ikk5bTQ4I4HSXsaE4lRkjkQ
dsvrhNvRjEfX2ofUYz3URqObHcoyaKVOGz/+DHuPI3v2Xxperh7HGk8COIWK
xdYO+ZkZAbD7/509Wi7x795vcpZbD+dWcV9sADj98dN/0qLHYQSP5vtqvWFM
vMvOJxOshN3PD2BsJOkX2OjjgAFbiJiPoFS9rntJrvqRKdY01ySmUxZbdpJT
rEPf1Ym4DJM8hoR9OeY0XrH60Xehtkw7XziHIKn2875znZ0bTWFLc0YblZSy
fCHKX37MZHUlli5StjZiOeGrJZwdMsEHqwnfup7bjyUXO8iQwBgR6Oxhb7+m
xsqDUKGDoz50KED/LrhlqRFPOFMawPUr/QxCi0ShpRPt6CjlhxvTm6MF2bJa
3m+lapBljDcTGYe4Whth5mBIrXVL3DW5my3U4FLM+TpgWykpPMiDbbNExIiZ
J8xbdaynnMfgRrUa90DAfxJ2spzGIIvbYWErKnsm9n8GZoFJ7dX2UEryGQ3I
QC/UG8DfTPGCRS7+bte7jFFUVGcwAuglWVGfCzJ85C0nnq9ux9OaOSRcgiiV
l+9OecPGXTpPnLyoE1TyZyOhSpYqTFSdeTs6IjgUHzrxpDmed/z0GHnp8kLX
yOZaXkVbtsALROsXnngPkIjEik0sd1WzKuWEL6M8BigxgfUJonigIc5mVCDV
LPufGc5bTVIbb2ihU56KrQ5n/V6/QsYLLDi2cjFdyTeVlsJH8b394ZytkGK3
WR6dIsAvsueAEBuzQXQMRmWGAPuusfjevlv8tGLxLGZ81GLdWGBz1x87DpTu
7v3t6RqW4AVPJFTaylVXoTfe52FT/Ikf+58Lh11Ivtjye+Y6zSU8fpoF4WzC
GKyL7bDvbhOcKJV7UjGv9fOgNaLzrVThoDDCXsgn2gaJ0p0LedBaomZdtc9N
PIHGir6zaDDAonhq0NaaWgHFEr1kGabX56JllU5i/8SifAHKYqHs3q9kOyqf
VZoN2B+MpS88667j2qoWSxg2cfGnYQ8Drh2qc3fTyPwgcdqWg1fL4FqEwY1K
DTCLuAt3dl2D3rBiq5nGvlceGducQgTp+crMi8bOUFX6t47MJLiVlAwlSqUr
5F4mrm0lHmFrYAAMr6mBM76oO6aH3OsjE0pHPB5BnJyWJcu8xEQ7MBRLLe9x
ojpK3YKXQIABYGEivxQsvK8fhg0uQoOabnJD0tSur09wxMK1/TKK1bXN2L5/
uRV9SrnT8Yqblmoxk8Jk+CxOWFUAO2tit5/mZXYVu1VTqxX7ceqkPcJrDojf
4sjel+rLkZcndawL3roOqBNfm2I19VnxzrA6SccUyxay8OIsQhbZAuA2XmRu
P4jLzGYLVqWMp3YWlbvVeNjKIdXFTsfWI9f2oi5wTA/Xq0deZ+Kmi5vBcrxZ
61o1fWgClb7/q2bBhs/m+0YkUjj/oflZXOX8obGsQ2qc/Jo1lyHPYCQTv5A8
yucgu1j9jdMtb2+aoUcl/dSwN+cw+HsLUiENIs52OalgTpqrutiCNYwDsBVK
7k2zVvHaKff1uR6p729RPUYGbJUr6/5/pw8bqAzE0e3f0Gi65wsgrITeajig
96ndx+rxxMzGZHmpRphTKtOh/2TckLd0m2/4EIGykQt90mMFPPWN4pvYGBq8
Y1ExYq1Z0s5UvfxuOTt1dJsRwWg8/L26CETh+VHOz7Goup9OL51MWrRdRK77
80Yle3fSZ27SVorAhdJmUqaf64CFSyH0tcSZNoWS8H0TBpW6Gh8f1RzBsXLM
2vMYtAUbEbDj3H+FlvRJPSUw2eztlTZIaNlj40AoO52+BKxs3pkdWVROgcub
cocBwpHn520rz2MEN6kxvyjcX1hfr7XpG650eQj+8b+qWNcICuAout9rzxKD
+k3HInXayirYvGIoGkqXtsf3EFRnh5mYJgXl4LoV4spuZDu0XVTEl/TC0iC/
8KLprlFNXrN9DbFwogDOoHsdlBiF8ThZLJHwPMTHIdKc6+LB5En7QWQSo/Mr
IapsPnRuzPbaQ6ac7defK4psk8/R43o9n5hagpXjOBaS4MhTp8zUdDLxOKKi
gCSfjp4fBPEYdo9WeOYECEI44X00ZupqzrCqwDDW8sIMy5x6Rzo0Gt+Kiuzg
fkmO3CWGWGYZbKtdDMDgZB7bsCGQSVGNI+CvTJrP/2eGeOZHLYdzSbPUBxSD
9nhJ2rY4id5XhIzBOkQlcwB8kd5Z13ZpsXPLYO5m+3oY1KJ99XFlaW3YXU0V
ZE94/ENhuIk0jw6Vljebx80FkD5+She+VSRimZS6mPFc5ZRNAnBM2kXuUyhE
rMyfqYCEU2dWGNZJSqA+dm41tvO/R+teAybKXDawk/qfqr+u/mS2p8jX5erk
rYoPEril0ZcDQZgV0lRk2xde3wj8TJDJwjkB3laKno9SV0Esv+FuVw11ZFHI
0xZ1GW7WVEdZI53jtGo/h1mzI4nqrGK+RgKoYw83iU9oxHIlUVNJ50CdWFO4
1bKPAUbkUo2/hcclFzWtptgWrklm3xuiszyZ6BmqJ3Tt4VpkA6hLRyABYnbq
e95J5BH3fHgAlmPKSK/ZpinQQ+kMUfZBJi7zQIwAGuy3Y/kDEfnGvWmPtD66
aRoeVmQj3U5x+oYE9P5FQqvr3cf0mm3cWrtrgVmNNPpCEtzBF1BgFBSvDieU
nK5cSjOrnFQkKVZfqtsXz2vwJdFsjftn8SZc7UYnl1tQpnuVoDk2xIUhq6bJ
cP0eQLzb8wiDXWcruQbvXssbjHbWoSFvCSaxy+NAet4lYCJr1TJ7y0gpbOU+
UP82bco+aBxulQqBjss1tA8fhDODox6P9bPc1CsiwkhOuAAoiOp+E+xSz8QP
NwpbROfeMVVO8p8b/1Ez/VLc3tYuKSBlDYAqGnTojNu4tOdTwjokP+9g6BDY
VErKEFj3fFNRmu9Bi+QuygU/M2m8R8Q+Y5i3hwNE34EHdSBg2UFk7FqHDh4w
FnXhLcPyhLegIbYOtMH3by9NoZT1aFXqWVqj/JlisMJgvHIzuSBMM4N8jHYY
aE8VLRGreg/OifFcxgwq9lPN7K2QpQRZ/8zS6Dx+NiqoHojr3C1i0xDmX20d
sanLGi6YLyGvp/Rdn4GykJRsXEG3q1hEgyjtTbYIRsvY4q3+fHctfyFhwIrd
X0tFtg/S4dYXhixmHTk6OyTqlB8ItNJvc/PA3bOuBLgaWDc7p2gH96L6WiTz
T8Q5XIDWFPDCT8RiH6j6ALTu7gdalra7bTlSbiU0BN+8VZSTTY8UBgANSyoy
+fjhhXhw1goneeWHg5FMWuk/1YVupvxrWQB/hamV37q/dP03OX9/gGimYoUA
ieP5MnTeVFD9KhuLI7qp7Jfr8ewkvhzPL9hihHhFn7dYATVA/s4IxcHaPdPH
VvkMMKzRpgxkudi64kVLUu/36UGSFFMD8qMSdw5qTy4HH2QqwxEXPtrsw4Ol
IDWzhUHoXO7Vz6wT8op2U7KdBuz+J+b/m/s8RwMd2CgvLrT+BxZc1Kdex4O1
8uqnT4PssbVRAgvkAetdB9bz0gDbSo5G1lrjJJTa27fjYLK1dGL34ZJm+xjP
3Yz/6zrQaAcjDLKPjVGt0Lb6BGLDW3erZoLGuSo2QE6i7odhImDDst1xXJiV
z2Z1nC9cMe718BSHC9OepQkniTqhvwjIPaYeHa14EzZE9Q9OLsKWcpyphE7N
paE7Zfhl7plf5hbYBh90cv2XETmbnneUmfbYpbDqov7NMQV8kyZprmlmHEen
xfYWPJvItAQhun0BxDwmdVUlWchNOa5rDOWaLDFw2JXMDms9tCMd1+nregRV
KJJf7+2a0UmC3KmOTysoO8Xsntb0yrxMLQ9IRRmPdFeq6sEx7z3bPLslHlLe
IhG8NHwzNCo0P0qGltopWHH9kTjejmWTl6LepO181JXXcrbZvSedO1L6CDTV
sM+6s4ggh6R+7iEWZ2j+PYwMXH+ax7x69GgQ9WFQd+ZuEpSUl0afS7vW/Wyn
awW1Z88MPidvUfJ2zqaUuglh0QLe/wux6Z6QuK9fdC0Xk6MiZdgMNPXeMCfP
tZVPCzBeVJsKiED+OYzTSeXTHDazHhG+TWtI0c1fRTK3xGkK307Un77NCHRI
ExZEWQG+u25RyqMMnvZUJBwR15t4UjSI2g1+aWQhIdgRaq7cEED6I/u5t8gS
UG2jp0xtgbCU+5t3VLJ6wyrAclRRkcHyDhIcZSBQoLjrif7AD5V5uc2Wcxz8
AJmj4+1CSOW259bvTB9Ksj0E10797O+CD/ijNs6eB+A5gUqknrIw7zDZedZr
o5cwqOkBfrsSZczG+2CtBb1cCD+SmMOqDZl3XxU5Nzp3A7Tq3l2bXyFfLRNT
yuS74nP647k8xipNZw74c+etvhOXDsud+khNgz/T2cidy0gfoAJieruFpcCr
GGmZ/Vov9iSset0y2Wx4enTmfUoiTJfQfIQ2EqMxENH8ySl4SWr7bSmJ2iR6
Ui2bx+rQcOVK3ezlzOu+DOTD7nTq+9Y3vXPEA+oENc5OLRTMt/GlKD/MaX48
Dz1gORoUbyEbJO3dOgRmsyisDNsAow5f1EwM+vCnB/DuxDbiG5Eil66geiTV
vdz+tQyQvH6M1Jb6qLGjdtbMaOq67wuh1NVTFUjGxgyhHwOwRdH6LJK+dKUL
Ys2c/4UMS4PIJBZXzNhvEqzDQ4UfPMMSYDbZRbpXOWJI1d28HziCW5uTZWW2
LLXT7c8EzOSQawG6yaOn897/jpz2rjwcerJrOk/QIuub9/vqWVIHi1crO5JR
s0ds4XSo9yS/V3J2A/eA3ApPx/BmKkPhHfivwVEtFMyjmy7xLCwa7imzykzg
9brAwv2Sbq5bJXLw+unhtocRnlwFyu77Cbs2MC2VyqEyk17bkU+pwz26faN5
AadxlDKlQiKQtjcydO6lNPLcKdvkI9gDpYBCwie7M/j4xykLZ3FWsN2eADtY
2MeP6CcEJX6w2rBq9Wj6gKbDetnd/VZdTLs/18ahl5uA4Kkps5ok+4YthQkJ
qjTNM91G9eYxbfzNGIiqCsVlfui/VtEadAKiTdxwN0oyZzVZCnmSWUKREE9q
fTJ2bb7fD056dtHc2GwexrpEVBGH2JDHJOIvWglklmTJLgcHxPdxo4aKcTIG
QdoNbRlazVWTPLM0GC3Qt4ujrMGnA4U2K5DlSnFsLIdofaZafEx27TssEfuT
5QvZbXv+TDWgdkpPj110DJikSKsUoBOE2tZ4qwnvQkejkndlZOcjs7kMPRA9
l90ML/Kd9galMf0LvLz5KQcmqVPt3PajiEIiaZIEx+pnGmgAIqj1rSUgF8aw
lJ7rg51Ph5QEF64n33cYlHkEsV9FVkiAShCdOfDuGdpnoedXyqeQtQ/EfxfA
lgtjk+IBlwDmfj/0cBM0xrslxAxTQH+C8gFuQW7kg6PnW04hGxAhDbQJYFCx
l8+uJwPC/4A6mk+byY1vNmJ1id15um61L2/71nj3ErAI4b9QVx83y3F4NPuC
z5kUGoIpALFoWYuw7e3ihmVaTCAj2xRBFnQL1hL4R+gOx1AnC1yxfRjm2SQX
8Ra1CTVlJgGv0MKyrnNgJIaZMtn4WvKpcBbZQyx1gm6tCqhu021e+xcoeAmw
n+ZUyh+fJO3HpbE0MefeTMs5iMhMVkEeLy6hE0ZoV7ElipQ8JAmblmcOXcyQ
jbkXM4VdYTgk9DZVvQePUTv9b/fif5eVg0A7zAk4AVKNPA0Ztgp8Z7FTd6pm
YwZ2IcawGS5Zd6HT23gwcOF30gCyjJLWmuD1EZ1aO8k2umSZ+VwtJLXWneIK
ljwKYT6V3aVgT0PoBU2SNklJ5WCPL+OIVLz/gJf+gg951Ru6Q3GcW2zqbDlD
bqHY6c36E3h/sKGa8NXTHS5FMVBfjJtssL9HuNFamtcpiOGrBWgTzslKi7vZ
7IqrbVeanLEXh6Dm38wNBU77o7LKWQODvFUTQV9AnKux7sP/qdMYZS5uwRrv
YaxBd6on7pvrCcNf6fHLzIRNXiuR/dOqbYd6GNB3DvPL8c6YY8G9U59zU/KI
Uv8/bsj6+NL9M5mYD52akFilnKgErBvYMdacdsd3F9nIXlFJ17bJxxpQGLXh
yU6lt6obNDW/2aRud7SfssVfNp+jQ0s87F2iR1I4+zetC6LEj5GPQKvtceLL
c1/j5F//3RALZ3NxdQCjdKidFVaR+zruI6+cntqVb9zJiU0fJPqxyztSBuqq
/QTgxIBkLLMbcVANzZg/U1f2MZhTXkfoaGlicoeen+MUA7VGxKBDHPYkCv6o
a1P/csf5+DxpqjKZ6iazpyIMjLfmQdhHPYmG+Gi1aisBOxCm26kpPGQzdeZ0
3MXEp4q7ymDnEJnUf12ixr35x8mF5XYSsD4npGvH0dD2KO+QTp4r2cSnBU3u
u/xp/IxIh14v7Lp/zHJtne+S8zC1JVgKkjZqC7NBMrJXuY5+Q7C1D93RV5BU
FtaQXzcz4YA7D07iCc0YUr44BG5AriHv2GnJpFh7lWyMvHuYbS6ja2Gk2KEN
bLuIVIaJaOOkkhVHB1oybRcYGavyUrv+Ms+tFHGIEf823OYKu0dy1HFh6Srv
dTKMK/r9YN9qhPOIZnxCnKzG6srMXwG7ykD9JQyX5GoFZsNXrIw0NiCgBZwq
8OV9I/SPgDT0znmmGrRgDueBZ1qUPb9WCPY3I0bnnp78qzvIJSUh3jLqvq1L
q3MqwWhubI1seubpjbFrFP35ne6mfuWORGw/7wAYVxtjdNUC9Sl3oenc46tB
KoOhW0+jDJYPp2N6MZY2on5j61y5o8cBcgVnD5jigGk+rrMYdE/MhtKz8may
ePp7VGy74NNyYEO9npubXGUF+v+KpE6Xku46CfvY7I6/YNvMFioc6/AaM20h
avjrorFIz51XXt1ueOSaWr7FBLlSTombRUWear4cXPAvTALLoGMO3PQhEIA2
6KoBpli0pR4sEhdKReO1BcOEP9zji2667/aR08JyOr6fp1tBndNbqZdIFd5G
PRvS1YljmlHTPSuc5tmTaHYLf3E/sOI26hZTtfPOIfc7hwwA5KYb7QxzI1aB
+BZqR+0iQGiETlBtH5w2wm6y1R7UaTLIy4EWbJenO0QJRm+KqN+3IACjLQ1F
LvBM9i1TRGXAj4LMOtcP4NHVo1ha4NKv30Yb3/8078xd0XMjldphFxWCsqLE
nbhrGZjlxWBOp0zC9nbYPBPCOXrIjxNKSs6VVz/m4wwLa1q3QqtY92EbhwZg
kwrgxDUHa5ZZq+Qk2zwFjtDD5+9TOHreiXg2IlS5aB2IjFZgqw7OaoW0NQFY
pjJhZKABj7057+N8orI0JaRWeJ+wah/cpNrOKgMtGlB4EKYb+IC/NAZumv8I
gim4FLUdOCUXrtz3ZdW2/DFL8IebKEkRyJWH4vTiOGLx2ugNhCeNtFWP4JA2
93a2t9Gr/WgsAfa8NvtCpnn6zWfA8lBN2Om2ewXIvmM/q2TqeK3b05r4Bm44
KRTkvuPS9WJB5omMmYdI3gZOErgOx3RyI+LXzr/07nacAIsNagLqj1/WkGc4
TKmHD79PvHWyXgGXtXR4IYaVetNMl+igo9eo3wvLWpcTSCLp7BFecsrkLk7n
QtODGf/1BJqBXr5afOpu/IcMrGaryxYYHSunc8e9hGFwfmveYCJkNXj+7EDd
t5vcPN5jcF39A1z5vKPC71bQyBq+NfmaHE6EyvnjBtWbTrqISv821THtWyz+
0tNM67HswAbn9v+aGOz3kNlJAmsY7a+z7hI3+NAnJaPj7Rj9qdM2csl7JHyy
ZWfevqEC4wXxsMwq+KQYUgY21MwDEsqurUxagRwPZXSm2ea+cEZlO/VkDKBj
hKAf65XUHfzHrCo+sqEWg5McrGe+H8OOv79Etm+kYLal645kKQCUcbxDpInl
I1Isv2rhU0QQ7k4ydJbN04eaDMrWpkXTrPysLxla5TD7Hg0TMqstTZbOYzwa
lfxBSbmr31I4sZxEwlO/YNINn0JQMWKRoRPMz+3rgcNWzukFiKYIqSFslry4
6vskRHx/vsJdTJIlYR0oFGVsGMNo3CIUDhEQ7GFfxk8hPdrDmbi+/G6wIBuS
LyxBDBSXiEkXsFipgESBDStW4s++1S7grAn8u3m5Tdw9eL/Rm2hAPxaPK846
/rHZ1JrYFhbqjcxgfajmE+CaUO2rxqR6WmvhKQWg+Lxf5vyVzBqPWqKHrjiu
Trf4IhMVYrrvwqo4DFvfNdwVF7czoxoYNXpnztfJUePfI9Mt0+0k/5ktdEd6
lNe1aPOVittd5yq7e0IjzT4KB9MKKoEbv0aC7wp9euOGyykft97rfCikOrH+
c9YF9UMywSXbrDbl0RRKFecXXlJcWfQ4fjpUO4ss0Ns832ZynEG0nGr3bOUl
ajj7tn8yMmWFSvkyCHuECAVlKJLGR5cyOU4HlsQDAaZvzHS4KWhzK7iEj6QX
fZFCc5qcogFRJP4/X8fGV2MllnMk63kSxr5Na9EqePChqz1kvL3a5kKWDaDm
XPPW1tplc1dLhKv1hpBmAkM61cj1j6hEqY6lwTarwk4dt84w7BerEmvRUte6
BYtEI667H05FQ1NO9/jiQRM8vhok7BjgDQ+wSKiWmCpzZnIoCaRSgMeiESJr
KJBK0u2/xAstREOc36OHn6DXGafPN/0UvMoFmFzekxDNuQcFH1L+mWFAI08L
XW79mkh16W1EcgnREaxIXokszz9h99jQ4Dj2Sg3zzSLKS3+FEPCcmr89mS5V
/LgY1eOj0GvET9bHqLmDYKFHLPVjFMOxfwyBGCugTw7p1pZPUygQ0CcQcxJo
J1ctlPmVXrAgHsFTDjlPQNxbZAqAA4YSlmYoaB7r1yvyL9ZBMmCJdLowjT+e
gce0phFs9Z3jLE+QNj6Z1k9jqE56GsmpBf8njWX2twdpDZJm40Nza3cG1hGE
2mzKcc4OlJn7bS7OqUDCOtvGByiqEfNc/YrU58sMguXe1+zthJ40DdB0ncQL
MIlsDktrAmtQ4nQrkW04VUwZt5JmmDwRDPTel2joIBMfe+Q8SquE+Kbm4nv2
Jtr1eS3rVNYOF2KsSNjzLXdE36tWVgB50mXh/NFogYLiIcsrqcV12wCB0NYr
f7qolj66Cj4N5wPZUuvgZ21cYbxnOOAFRHMzirjHExt0L7bWx7ZEdM0t8gKf
EnZFGrpehZJEt2on1HEvmkwqdH6LDk4xvSaoNHgNHPiFIIqE3E+W4gz6yD9l
RuX/sv90L4v2Azce/q8gbRapKvM+wz6nC9/gS7AXpleOEseGEaOSm0X0wcdu
UxMdtTTZiLr2sKPz2fzcZ/c8Gs/XqEKCBp7Ms9B2PttyiyUVVJbFxp3GN4gZ
qKOL40DKOajNozSnRJNjFRovktSWWhsEREFhfB7f4FVjC5lxHCroTDxENlEC
aopZMlPXHvxe7LhdmwQ6C4er9WcdLOEcVRKF5qZ5yIiPx6wOeuFsU4h5GcX9
aPSAjTjxnK2Z+rLt60LeCv3ikcAWg0cwpUoabZyz5rDbo5BUN4Xc0aW70On6
ofzdjzIgSzusJWAg4D1i6K9JZs2W+Ty2NRplqQ6tZ9nbhqLEVucMqYLYW/eL
pMjjjyFTobHgNSxRBMZ9B6Sfx005uHo2oXCTrIzae1vxXkPPpp0wigj2+RrO
+/2xyDObg8fuCp3yQMJAUbxzQ/w4eUi4Sg2AKIoOZbsoxoANpn6zBW32O+ii
+XBBaV37gyxm0Sc20L4kh6Qc8cmlPG4V7gSSzq6smp2jYPrxiLk1i5b7CD0A
2mBOGuPzN08SNBl5qDeKHcFyvuQYgqOXQPMvQXMx/erdVqeWLPktDuv0eF+7
ABULhrIrtAm/msdb/1lDycBf9TwMYlWPK9maKoQakihYlQ+hwR8+KfSLnT7c
FbdVqVl0JK7c0vJeD19zn7ywPV3Ag9Yxlpqm2QzCUSteAjq9aPMIbU+9XAEM
1saj+8XSqWcrCZfLxmvESR7oNmJRa8+5QBVnYWnCaal0Vs7BYf1ZrsTfrdR0
kz+U80/joHWPtN37Al5wxkRaaPbMdN8zf2NII1vmTLDy6ls0nY/g7kbDrywS
RdA2ZzIxipex62EUtVQvT+FIWvPkIaRfOTE4pGXKh9AcZwSorAlzT7NHWBKO
GjCRqh6HXFrqenjp15//cqebRh5YkUXZZNOoIcxnemJ59Faj75EVNUjXWxiA
GvwVgb4r4ySO95wbhD/M+SJYHnD5txie6BYuWGgH6Lw0p66KG0fkrUdKh/Ri
pcKrupWXuiOon9JAnZSBq5vpZzMo4+H28R2mdzsGg8vVwhvSRmLcadpazNIl
J6k5NzbjjE7y9S521rOheTTDyr7grOGPTbomdKaUHWBwwD8TWctzTb+G69TI
f2C5dZsWtgwVcd57iXWOlpAf6F8iUJvqs5mMBRZKkv0vPDaJCu9ytmdDGjlN
m6cCIjL9VHDprc1k7DjH0f+nLGvG0eE1MKKYkW11derfKsFcW4q+nlOzdWD9
M9cp/sZSewoO2nNfrapSnZhaGvb/95nGQ8OCzJLdml9mb3Bnq4zP4Y0bU1oG
Twk1ZgL4K5BlXHt4J6dCOiCc9BxYQaImqfaOnMQmVNVfoMIIvV25DapiXvjD
suS/W40ifVbIKK0dBVfyi3mCNAJTYHMEkAG1exnW1nBuw+PuQaposTKNeelF
70CNEtfyhunSXvK+jms0cD/eG5BVi8FrCgN/tGvONptW9sk5RESOjRSehrFj
BmFjsyzNZW+JCzTK2bDMfQ7Tuljrh4OMyD5Du80gNdJAPHPCQjwrb3hM8kPp
tZK3wS89lsMW3jfq/ZxHh+9wQ9xvE3CEbdnkRVF5AQiGdcLckWa91zTRLtI0
gD+DQQcxKhgBoiLKOKSLjlQTACC6tHkqABMalw6MulogFuRHRGRAr0ivrNg8
5Po/H1VRb5LIjihvG5n2QIm19e520G1QVz9NYlhHlHNHaZ0uIF3gVz2mB3ZZ
juYaVqHpic6FdDZj7iowNQRDjcGfGb6G4SyFHut5CQP/DXFkMeOQtk0fxx48
DQabFv7PFS3x4QtJlWGDSN1jN8MlshNYP1y4RG+VsVWaNik7ry8vIF8m8bFU
ed98KNjKHjMPkl7h1Xcdp4ucUZFMyCEBcX9g2g0H4siq6bT3SgAmDwWcjSpu
BiIuQntlgGfdcWwIgkbKFesdlFDY/82z3cIS1wLL1kl4oO+p+CfylLQZCUzQ
Izz/k8pFiIS8/IX/2dvTnpWfg+9srzvXmmkKmtf0n8K8oXRtlpe4fNi8JVlj
4aOnyVih7hDzqg1f43NxkcgMQ/GgUr7HOHCWQVMB7Fked95RzXM28DlXEe2c
D88ikdC0d9Sy/+PsJr3ojlSZxbQ7IS3I/vyhNK/1NWLu6cfFYQ3OVBd6g3Ll
2eZrFtqT27WhcVmOMJ9qyE33P68t7JU7OPjfR3zEgkWLbDPU8OZaKzzRrp3S
c1k1F7x/WLTw6/zbWWxloAqKHSnKu9SxzjNQ9HJjCNZc0/orqoBKVkINuyGu
jj98BOlb64rJKUMJogFQkih5G/qZ/O145KlsB6/Y6l1WEH5SucP372MiiEni
hSxUpHRvaoUTZ0IXfVikclSKXP+DTdi4O96iUDetPYS+/0E3H8tP5/ousl6g
3wbEeFtLElcBa1HChvkPRe+cxEce+Wh9w2QOMvQXxdIdU068E8yMY2fq59Dm
TlDwuJ2vKRvDLy0arx31KmV5hoMHTyqHQXeH/bEcTrgNzR/l8qGL4REm03fu
v+7b7XI36M+PoMvyinOBHEjtyWnLT8evsrfVcBuAC6XvZUR8FHYuNGXib64m
0PkdzvgtzldvOgxkfhG6gFNnmiuvRHxDKaiUujghxu04sOGOBPQvFqN8aglb
uIJmkDS4Dv4Hry+j2DXp3Xe4McJIqgXP1hwpIQQLmxJUN8nB+zJDjudSCs88
yKXBOWH87CHOVEPJ2S4/eAV9baxoooNYYb7qNKvQh0YffS33asTRus87ahl7
vDm3FE5HACPBhnuSj6EWd2pElWgdKjIr8jCcsC1qlc4QFkdCyCRiylUcQxmr
vHUxTMUjaOJ9byWtpYo7i1adEriLuNBCXVTHOdcyMxnSPz47nZeRTQ8/uE0M
K/VCSP/c0r9v474AWPAH/fsZ+yGsu4T3CM+xc2HkZw/6Mz3otcMuk8jmnOhh
tXsjbyhAPuPCKqOHAMPnNeIeQerGzRCJrh+y1ck8ta1v3xzoxFI1taLFtqLb
yzCp+eeIcEKO9JLBLcJnpptqiQlILVCOvH6kXZRzXMEtTlQzf9Xxa9IbTfcN
zVLFNfFFeMHMkeCMl3K8Q2oyTyJTFWrQ8KRO9/Bap69Us4jcrYdAjaXkq5a1
GFrcDyPmAK5sWrMepMUkkkvlN5P3oJSlpEpDQpW2qD+c5Yz2+vXguXTWJ1HG
qeB14woN/hbbPjKiTSq5T7Kz13aYl0RJcnUGWnuCCPFd1DaoIzhBfIvkh0Ri
KEM+C0cbqaPITuRH9hIVMlGlGlBArrRG+X/+NfxYP9PWiq2xlK1ji8mfFjYC
gZ+Z0c2bzzvXbUz4lmm1N3Rza2sx82sAYIvS5ubRTDl1DrHtmOKt8RUuhzcn
LI8bhK3uSk/BPY0jT2uLxiyjmCDlKM5B5lsHCQIZJfG0kAn2kR6/52fbKZbm
Uj8QK2z4hoF7AP1bla0zFJncXNH7Rh0pqc1MlBS0Oc1GI+ye6nRUzLlNZ8PT
OPbTKm1BTrZTjHwtCbha/Cga42YiUSYnLVWVuKPeKYD3HRW0qj65Chy5yhdw
IZ+Se0whXgdscJiwZsbOdmPYS6kii1Wum6Do51NqVmW53fQenNCypsgtEhKA
vMQNlX6cpadsRU1gfSF2/Zp1O8+5s0t9wwr1riKWhbdGvnj2TWY44NFgdOVL
nO1quaMZMOEQsLjVgqvt/EaRn7lpDT20+ed0P3H5iFdk5oMYU0TQIO82yEP+
PMDfez1L3NNc3tVr0MCeR8iVIqf/qK3fe0aIrtEBLpkj2zKHGzeL62uPThRI
27c9eLM/kgtnRijWhKOer16YsJqtW/9e/GcgnktS4Vz6oG3cUg5YK8J1tDis
Ws4Veedt7KAZFlLV3LtnD1tLTN5LKgZuyDLWx6YSixkAvRh2SDSE1K/rkv1P
biVlFe2wnvcewIg3+l96Dm6HpSO4UwEdjOUGZEhtC/s1s4AT8sNzIUunTSmw
/EQxThr//F3roYjLDUz0RQac92P0qbhumt5nuqqyEeE+HGz6HLqv+QmstiH9
B5Drka99d831iXsenfXqp+b9CIQGvRBIagGVOVk74rfmgLQuge3XM0L30amM
nXqM9zLVO06hoHvFn3IqfbmJYQ2Yv1kLoQi88Dp9IgkIhmPAR/b/tIXBbb+G
uYeDehPvrTaD145E3G4z2/dr7Z0uBXpaJ6kayJrd7TDR2ITY1f+J4s7LOccL
heVZFUAJjx89/WzaQvP2SRqVQEyEP86Oz2fgbrmz718CUZ1UWs9xO1x2btWp
gs5k3bFps6Hhz816KxAb6rtjdxWpFRQoB/X3BMxTOBfD7lXmwwr++VhmTAdS
9IAzCVNH81enB+R77st3i6yyAtbKPGjnCEKPIeQ2gl04tm14TQ+TcpYz/oX7
k4n2+Cci7sPQgAsttMENg/IVQEQ2Z3K3nq3Qo4N/dc7uZBXexKsQkrxv6m6c
9AU0mnaIFaD/HDEGhcTsf7y8C5s8/P0hFTMm+M4wOEeq3boXPeQ7UTfP6BAD
gZruEVSIP3QcebIUDG876CRXHE0nEmGWbfcrdSZHKhfz57wzpvSMi4aTKpOB
65sjEyeUMswFbXD35pjnXGUEwdukaY9E4bDsWLv4m5us/+w250S27HdRYgkg
rm62wHUVBvHjTrxyGQjJ6UzUgGMIAVhxrG/8/Q9ugEJeGBcK4xr3IUgXCyeV
b/oPUIV7XEwP2RXOI+0b+C2j2Vmoz6mFVbVFpiY4Pa6RIlxSZIbyCKQHtD8K
Bq9M0TMozpUs1vGcKdUR7uZdcV4tDVmf+CuonayTrHx9edudJ7a8FqkAqAiD
fAOY8xe3ORzZjGpt7vs0sKDqc7T5aa6VxcgNPdfvWhpa9LqmfYn6RP3+Jpe1
6ljsX9vYQB7ZmuExe3REqXJa8zcGBMwIqg/SA9fSqEt1uBqlkbHNNFgLOPYz
Eku9YuvauOebXBHUQahPMU+64vtJnAOreo/ZowwgMIep499qJ13W5RhQmHTx
GAcjK3XLrLqyIRqk37L4sFaxn9rBLjoM2DFx7tuGjbJwxyOiz8loKt9nb9gf
XDL5uQB3en0qfUYhfWr9B6fBtnICZ/3+V2fOM6/nQ597PtLPaxRjVtnEdj7w
93D81xQoPXkQMhzLXkAN9MqWZAAqhBE46PnRx29fQgULAMTtV7i8S0xIrlb4
rR+QnRGfprmRtmITEkjct+Zr5wp379bVsgZ5PmAq2aYOQBcaR22ZNLD5B1nx
Hd8EjNT9HX9juytGSU1jwL4hdZ/Hf/mE+nNzH3IC6unKmqezKE6oK3zA/1Io
ufb8zcMldYnfQvOibZ1/LW824IXQ1p2axDbQ/RJoTXDJ53yfI7/UmVqpKYuw
6NTrCIByjujgVkL7OkpO2j1QK/BGvjENlDC4uqXyD43FpEubrLg0ekdc5xD1
yyks4NzIQLqm0nceKHBYnB7FdYKx5HBUWOyPJ/nZp72Msfx92aMFxnCbLcFs
lbF/PbaTxhXlTia0V5AzbBVu/qKuNzPsJrv8xvq9qEs2XZO81v3J3DrK9JjZ
Q15t4inf1rV3p6okvMaQ3TTYhedH/A8VlDLevQsS7aFd5PGdCHfMRlIcmSXk
PUrFlF+PKoEfXuVaILUnYIo11TsrGUdNtBQSKJjzB7dTtBng0JO8MrXH5UyT
MvHWEmXfic2fuIksImoMKdlqJrv1KUS6cYmcu9z7BdUWYmWs66Sq8DSns2Zx
AcblqroJ6v3s8SDjsgwPFUljBxXQzYj/6dMEuEIfZC+5nnPxI5GKPYYuNhEH
NfxK1asuRCN76Mq8sv0dHNYQq5q5JhT6U43nqY0BOeQk7Xd3eKXQoUMf4HTB
px+C5GMcu/wDixjuXIN4CYk5aoPt1+NKQOriDK1C155mCf+FSos4Q4729Bke
z6tP2JgAEY1R6VRzq6lnwgJ3+b8UUa9R0XUNPOZhcpsTc62AgqYAwyO6aCDV
ypxWfFtVmyuU6XDs/Aw8C/NBj8wBpqHLn86a01ufrmOv4STYxlKxNHRUmazC
F9Z//pWZBUkBdENL1ZTiFQy9rUQ0doLcyJzYTBWMP8vC5uelwQ8J7z7N3sP2
yKu8bqoViEWuzB1iCuubJ5vQvPKn4FWtTQMWSuPydCgu1cRuj0WJG/PbJQZF
4yzTWwD0YbFqUIVqbvJk4tf/MDq8NcsXSq7V6NZ2b+eVIYbEeTCy6wf/8YGb
PpsbY9rXbVt8yVX98WTxrQ06u9ix2i0KsiYBKfIYVHLjif0ZlR+4+ssVjZ7p
BWYBrwWESDZZSX0ai8ISuktgarGUncjd1TC0Dnk7elLCHFRIBnxqYDswXNuJ
ysjAtXKiADoWqBZ3zNuAggylKoV+WOUSoDiZwX01eN25DwgBhM1I2uslL60U
f5PTG1MDzj0qxOjKMck5bflYmOYV89PbuH1W3UrtlZxlNYUMAzhEkbwHzwhu
5Ff16XTzwjjXc8bw+tOZQ1U5DUcjt1lLMS6hpe2VFwIuT6ddNiQ7F51MN0tg
qGrKUu/21yYylZZceRqce4GiSjmVCsrvP1QTqTks64EP2s9KFsLYV4A+4HWb
0l/FKQPtQlh6IGX7clHwUbMzxVJ7YWW7sWIl/k/HeeH63K4qgDtj01WY+A5r
69UxdTgFvgvnH8C8cI8hNt6YfKwUaEYVdO82Dc/kKLTMnJ4Dvl34/X0lkFun
m+KNCG59+oEdfJ26oLtskjhGWh5S2y/mCbhq0MdAnf87kFgIF2BOlbszCN3T
0wVevCFmjocFV14lhm4lFJ/4nfc5QO5Vl7KddKUGrTS5hiRmNDfIJoClH2xN
3FY5aF9Rjej+u2VFPDW4+RgDmUlq3YNu+USZu48RephZvyDC90qfRZzFfOf6
y0p9hOk0ZsfFlnRGtzH+Jah+OYE3Tb932scAxwDVBb/p0jxfUofqPaN5hkJm
x6mIw2ZsXFvdsGYfF1Ae41blAWnW7X53iTXbMUB6sPuD0iUtJN4JTPDuvWUJ
3J9/95+Kx5ApS977fQSVdH4VOz7x/wuIU7rb4if02iQqfm+Q72eoKBTPl4G4
9/8hGyFR9QTm2tKhxn3LazpbWB0Ju2+9owRlDxvwYM4Kq+oN88fHrm0LN3VP
pK6+oOnL4Hj3VUlJFLAfZOovTM8sdDcUTbr7oHmWlz0gLEy4+XDtLNQUXDo5
Zj1G8NRrLpDMBWNfPlSrtMB1N0oBUU1DPiICfowPrTg88IW71g3yHZJkpjAH
5GdKEwVVlBOUvvnu9vI4L5czZe8Q8N9Sjcg2+3nugIywGOuBYcEwc2hYNmLW
L2OvsVV7/ive4RsnR5Fal9UpfhlHUxkuDB7YJ3siV3RtrKVabk8+fa28LUHW
Um9lxIlk6myGU13CN7M8XLgpt9feMffeWZL8HZEXMSkL0y7TYiiC5Lw5ttgr
ieACzLUVPEMB1g0n7oH8HwPG12gMRYT1LPtEJAcWj0BIq6aS2NxDJs/b5nOS
G3un6hmCDKQEfabxQ00IsPr5PDdDuBqaq2cIGGKjNBKpO/HYyc4QLIOVs8Vo
eOZpaIU55LrFcpVmiL8qTT8YHvNaLnbsUEVgMvdRXojbsHDTrPQ3D8wqkjsN
aP0fhmqo86SZw0inq7m9VMPRuBBC+flaKn07ug0AcvEo1UkTnjT3ppqTem97
8f/ukbBJz1dddu9Lt3w58cX5zbISP6MM4TOitvxdDSXN/+0gjkBkS9/5l9Jo
jNHBpHTAD9YyhCIdtJC/Wbr6xKHBEmx1kptM0BWOLgr6TikC11aMPxaqxyNn
E9knS0j3PjvXv29TBhNsM2DyKJAgy8rMAosPQMIPxDhuRrINJta1tNaq5ojg
PhMb2BhP78f2eVJKKh0/xCbWNQ21Mwvj+G/j9AHXEYxA3R+cO63Bv6Ay2OW6
mtb+/dSBou6RvgNVLXvPTZX8exT7zEBpYjCLBG+o1j1DnpuBkdBVqOezdFw5
OsHIdeFR1gkaBrxDxFCVRAEqe/bzaT7vPVcLQkn0iGnLoMUdXRLW645dzJmT
DR6CJPOYYiM9RdtC/Ngs9r/Dwxs+MMeET69/t0NWqOuJW4rIt50XZit4pPrm
Y0ZjgKcUlJuKZocjWwZV3Kl+PgJ8mq0zNG75UOXqMR1HAmqcYCIkhTaSUgZX
LLFO0piK5ENGza1rHKe20o2Cej4slzDR4zmPM68yToyiMjZfa0pNjfkRltz0
pWGA9Vi7cT/fPqFzCBRydKyiXCIc/5OqGkVvGzEyhDziigmnRPXEOpMKLUKO
O1MtkLgLHughuAtf7nJfKYy4qCrlTCd+eYKqfuVhJpI7CK2m1BS+Md9aOiyO
Am43H8N9fwJ/qrA12JLMijYLdiVkdePK7S13eP5dAPn6nLj/Jfjg02rMhWO/
1GKLofqquoxGsEIL0QArsCieeFu8SR9Vzg6T91zsXTXkwXcB6EMaOutAqqkz
rAjCIB1wy1Z5V+55DSIlMh7QET9hkKVZRlEAryoxoA5l/UwPoD8lXV4YAINx
xM5SoyD+TCgv84cAMjGj6i6m8Cfmwa2tKqDvXe8ZDbNpesfuiibrOrmXSc2e
/Y7MhpUSG04Sh0tyOwaM8rN23ouPspurmQ70rINT+sQu1wcvNhM+Wc03bU0R
mrWnoUF5Sgs/YIEh7GOMZt+dUG6+uz+ZR6f237yi0goCXsD2Q/3+M/ysGg6B
LEbMc6hwkTNEG2zHLlsQ2QVERFk9GemvRaAnOyYtEsepx/d1l8YwVqaO2RPX
4c0SquKmeG9EItkVetSJOAxbf9afOGTYIGMsLu9UM/LW7wn7BVT0NCDIkUES
yGcpFYHktEzvby+pl+Rcf8PxaE4yygf2t3yLwWDdFz8A+f1pMpF+2Lwx1qSM
0a5QVW5+tHrWFBGw15TBNe8c5bN9mYcuzK+QDNhOnSVQLyYgA451sj6Cd26F
6RYpKor3EiJw9qAjla/4Sp+VTALAyWNEHjZOT2YnSASoj7I7SwLgi1aB884K
xTLCb5jpAa+ZKNvuyqsbe8q7WGbt8aofiMman8wx+RZmc6/yc+QcFRfC03F0
wTj4fdZegy7wDFVLnmkgA+G2DPRW6tbTka3Nqe68I1kE8Z/K0mCPPTGMQayF
N1x7fWzBJTSNVuGbU9Jn5GSlFhii3cPJ3kMiDpFmY2puJZXTpkFEbbarADIM
VuglpSEi2feTsgfnLYO/+OUGqwG0bzqWv+UT2s4tISCMmNBDv1bEXT8wg5ii
NZMV0yV90mx6rHc8nMSMQ2lSDd9up42mOFD42rMSN4/iW7ImUvmsdH6zRxmr
901Dg475A2X9xrEtiUiH326YrxG8TzhthWGmg4g/25rm2E6GHZEl3lQIjWvY
r+8basi5fKl/E7e4RGZd+xOvEuIdKaG8E8Gm6GANFJU+UZfiSwSkjDGhLp5+
AkngtQtRvHuRj7t9w27MZiz4lcGCeHO6ijGQVBVppcuG8Qjmdd/DMrIMVJb4
yxLDwLCdtRicDwTD+Tbkfw5ZTv63iWPWDJF5AD0X2I97klfPgezHoL5MW80U
xVIiQderAGsxZHm6aY+JSotjDolupCfo8OXFqiE7lilTjLIH9TcoYvuW1GwE
DZz57n1b3ZmBv2XJIO9lrqCGa0eEUq3IGdWPR/rqcb6AQy6+Qxf14ojUezhd
ra+2PB4L1xVZ1W9Sn80sEF9nyQEPX+b0rDijVE4WVr01xtAQGvVpj4k+HW8A
BEPsYMi4wTHWLK523mQJGB4myLrWBoItP1ZCLAe8smBZ+TTLHe4elkVc8fOC
6pFEllYZdhPt95U6oLbyRyEt+QperzoOMX8nBWjRnJp32tBrDUMOwA/hpOR3
AJhkyab2yMJ76GFQUTMiQx+g9T/ygZhrlwid0qxywcCPWxym8kIEmjXX1m5D
nGrLqmJ0NwcjGPtZTSm3DzZo9bptp0usmskSQc0HaBp0T60BessjRUGUL1Ud
vm7dqbmktNiortHQnINHZdWu3tpzXLwhCRe2WGJeTou78lITvzLXyONFWQEw
EfC1qJeyI2R7/QeQdQKk5MYz0NRBrQHQpSfn3v9oZHDISVdvW26RQz16QHEk
A4/dBGzp6xXJY3YXrWHlaVx8HgvnDE+hYMnYOXIkQqpHlAVjon672CSYAOKs
B6rfAoy8/ud5j4++lEJ6YHrL/GbAljWLdPuMo8BZMA1VJIY5ISh19iyU3ykr
p4yU2XmXI05xTbqZ3SxHrLtRA+QRTs8/Ks/cwmQYsIoFA742t+d1H52nUJPI
amyEoyTNqo9hifQzDlyBZrCqEGZ/R48soN+n8iZcQUexRTgPSQRTetVLMFed
RA8RLIQsEU5ZWkjUJxmWCM5Ned+SNG5YMRNFo9XZ168xLazGUPR0xO2vW9qt
B112qmt+e/rMyDeumuUhDDVTiAQW42CTg6ziyJ2MSw4/s841ArqoY5M0SpBy
wJ2djxeokZt7v68eIkBO7cqFJs+Y/SDQTzn4JM6osc2AwTxrTczD7e07FDoI
MIxTtEULkzL5NG5BSLx9T/shRYSlSn2bRg0nzS4U/u4PAyrLRDXWSdqYFYJy
RdHBUMTY4LKtt0OTSpA1ZTHWcNHyZsJUcFG2fHlPmrCDrgtlqdMKO6o77ZSx
BxxbP5qz6TXi0CqVpzTOcBzYmCzs05gvogbxvB8PlWyOEEGtqa66jpYNttcP
7r4JFRqpH58DF82jKAa9voNpYaO8EJA0NQ9tOzOze8VQ9w5rUYRbeiE+Grtp
F66n4lIxNYIhhwv8LNk1zZiyZ84VLDdcAjOMmUVLFU3tTCs6oqSxe/+mcTGy
hMtFaKm8asn2g8UfXlfpNkQkcpE05HJ07RC/WlbBBEmv0LV3rVXHgdagUG+G
puctnSYIqX3sDw721jyO6XrzS7hm1E4xkll+EdtZnP68KN5NOSpUmNLgdRTg
Uq4bOvWGoIvFT/84poL0Xt8lX2TT7/lUHs5ai8rxA5FCZwLqVH6XfN0S82F7
2tsL4NfM2R4rc28AX13uTSw/HC6MpSjy3HQTbDY710r+sUZZV3+dGfePPmvX
PzXmkWTGkUWhNduwpZKsVcy965CSvuDn3qg5xcqn2BwKFPehc7imSmaep4tB
cpbGStbskc27A+OoNkVvZwnhz819NfuMvqu0345dja2ECp0Y96vcq6eyhHzG
yTjG19lmMPk6A/XbSgDQ1nfpH+8Eg05292fCSM73o0TxGWArgTayZ9fpxc1h
L4E0GR/KW/muboILwquz9JmGrf0mXpriHlPxZ+UhiqZxzxVdecUkba1QpBcA
cZvCMMvFVqLZUdX+OyK2zx7T2Pe3uGFyUBmjfvULJDQLKh08LUCh+MnNSz2+
CA4I+V4TSu26IrLAGNAyCOaw5a7NQLxdK6Z55mDs322S/AHfIVGoFGxaL73Q
njpetywW8eh8Ag1Th8obshqntmjeSE+tDxbUTSpWJLTm3tAEa6Db8dzZ3h+z
qFXcslYzTDb6Yk54BRRWbg06n7d9BblLMIfYlLL0fFDhP/Ud0ChlXBHoFeQX
VOXdsPj/woHHjdGtEqcflvRIemmYNubV1U1Ce1zbqT1Tla4mobhyUDDTJRsb
Hr7Jr4zBod8qn1M1kcgEnHVRxN6y+Xfg0wRqPe+fVeQYDsujZlv7RqF7W/KU
QLGbCmb6qH+s+BbFLq8DFlhcqP1qtdAvRBy0oy2jBW+On3OnUoAeFMZWJn7s
K2ZUbpNAmG+vFx4mHfXg1b4ciekBFk4bMUjxcqrLfO78prYdtdvD//SYwvVw
HaiqE4PdkmqnBrIijzBo1K1Kl5Rk4yCsI1KXGKC5Ury/nO2jMOEuZSRgN+zr
6aewZTCLQ67wvymBULvW+wqYMMOeVeQKgRNF0GEUAakw4Osh52CDEPrdsCf1
4iP0V7X6fJsa8c03Q4BzL3uZQj0ggjRbb60D+1MpmxfD75jQVd2v4Hk9X+DT
iXKA5Fx03315LyWHvmxf++dUsJb0199uXnO9d+rFfx4FXuGj/g2tfX+F6FqB
3CxL5CJCT0SX90IErSPlevKFOq7oF3m9RRK6LP82n1KLvCJX3dcs/Mf5M6QM
a7cAxxeq4SjGf6VLw83V2oXiFwAmyHYUhe9kcTO6GzsyWOx2BDTcqJpdMHN5
K8zXF5W3HD/MbTPvcOVDyXquqCQ798El6LkBGaPCOOj4ZQW1SibKC7tAQTUn
5dLRnQu0s2gTf3YKJzPMjLSBu2PLJV8vHeCEeTFEzbNxAEsytsW03Zv+57RP
x9c70eyN8helrtBbhDkRmot+0reXgNhbJ/nwn3kfXMp6DAKKoiClCuWQiykE
0Tyw6X3WHubVqVCyuO9Z1mdsVjaXsYHNYHcv7Ul7jyLLHKmw49/DjvQLWa18
cpUE0yXhUhvnbqy+OIK5AiM+lHsD0tohCXz0MAjw8hobeWoCKxLbhe3QQhvV
s/svEsTCnTwx8lAr7V55q6Es4gns+A9rcgF7DZcB7VXlcmTCBC9Ytgxc2Duz
nI7QNLairUkacQWOTGgKeckI6lEoFjtT1VAbeR0ad2mrUnrZ0Wnlv73NqJ0B
vUbUSxiPmPkqnIaP6TyyoLA869jfCG757sDV2tpF1KpaN9o8Npl4AuzXQ9T7
AofvsBIyi8pP+J5/s+r3DIf2ghlrBIhzUDQzaW/+v4fsd5zDXuut5gaOLFyS
SeGlhEuLUQ3LYWKwxqD91B/7fC/EiX+VlEtFC0ng3UMoSV2paCY4GxZ1rwuZ
U5ieyWLJzOGTxPF4EFIvp5RRYAZo0BbBGm6rfn2UixBxzT6qXDJT/INZlhMo
x75iBipmMDUHsMgCQtO2g3y6D3Gt7kLhZV4Y3oZDl5nLDG/lZzpLyPisDayY
BFZne9avE7ad00hphXjrR+WefN8hn15MkRMzG+GhGCYRSKjFu1B5/w37oKDX
iK/ePxuI2CsjVVA7A+3Eb57BU1yMyrVgFZCJkRWKj8VBIRJTObgcMxzDOFcQ
70Hi2XkuDD4xHZjbUkvX2c7sFo2CBwbq/W5QLhB5hS422QpZUfpfaDFwiB0t
qGCz3BzLY+jM5zgZUJaXrUypro4f5VwtUxzq0lDWFFGdpr17d+upXzOnCQk6
cAyk4YI+SEnRTpXFPu8Hz1nevutTCz8y7fsOedokb7pOqlIqlPDBS1j5TuvZ
DnVzwDgaRpCazWsKwH1zoYQKZlaGBRVRN+bYDMgQu3DDV1MkZPt7xFMZyMTd
GLzIiuEbniO4UicJfxooUlIBwGV7pBfoNFsDZ/HyTkVAZfMdTbh1C3PS+jHC
ImHo0rH7k2wo3lRK+dW5MA3wRcLWViaNargku6reH79mQ2FT6qAwB4cJVmiY
oQeTAeQL7L2z4MpKbVjhSTguMFayqfWCwTcICPAmd9+Qbx/1834myI+HFm5k
amaC5Qobi0/qfAttBBD0dDfQ1w6rFftH2nwDJXOyAL+qtDuE/8ThJObiEIpT
Aijz0mcFMHMZ18COa0wRBOUKLyfakZWSn/xoZRu/n5LLfDUvi28TMGEjBz02
AYNWwq0XYJBM52gNTIq0q4QE/uTzhgxdmRIE23v+SRH6hHD6QEhj4mbm3MBF
WHCcSs+F0I5KGKgt8zUGPhIkx35cJVaK3uE90AOeObcjO66uwTKUxv0jBAXM
d/WIXtZ6g/0zEpru56hR3atiYVNtTO7Vg1n/4ydOKCgF85lcccNSQy1dyhW9
hctV84usc3syo8OZ7XKRzIT08JzGSOBfwSoD4S5QZr/P/4N3ziSHwkuW4gLy
osGksq59XZIXqtak53H2ZDljfcQlhyor+4C0ItiKTuVtIKAGANpJQhftPRIq
vbStPnWO9i7jTzRaqw764eXxoi2BUFrtv74KC0pouy5KkF8aqqk3/uJcVbAs
x2Z2mwqyI5uFtQENpX1GWPXzKW9gVbrNdv8mJrxjcfUc5g8+Cmv1M6E//poz
juOLt3OHqO0rsjqYBQ0BeInbcpezC4TY80lVSvFgPJGZnNXfdM9qP1hBzKSn
8geQk06Z0tqVUflAVqmhMIfnkN4PB+eMPbFC03j1G10RSH2x3VQOTkmduUvQ
0SajPT/CObvvnt3d3wr+/hmMlznwjU20THm4ko04oCttn6/KiIm0+y/CkPFm
WFOQ44Js+U7pNNWw7CMJfPcNRPO04sECMnt8lEUC3K2YiIAbV4myTnmE3NoZ
WExgVuOjJELHMAH9COb1x1wKqF1prZUD9QEx0xDF4wdZocyUPd1ucAZxLIjK
BE0B7BqSHUH3D3s+FBj3MtSE2EUiZYrx+MC42WLaae5D0LzrK2SwUGWRgTWM
E8HYVPgx3jbhkHCxLNDqFc0vT816YgmojGYMARprNX7497lnLtSwFKrTolcu
j+gdkD/8K+Jzb63nKejV7jgXXEF2r4uq+PPa7o9FdnRu6KFCqpuangrT77TZ
crHvnz3N42jx601veEvdQS61OXJxLpJXkCm7BRI3x523hMiWIe125/Gm4qTK
3BOgqOsatGaplvB4zj9So5v85c8evImPaIfGyJyORUF8NWnqrMxv4m+ZF7du
Vf///bujoFG2ZmfuCEQeHXlnSMQEmj64/NuHp+a8M78r/KSjw8nEgYOndiXn
yjEmsuu3PfrvLBcL48BAOXlqm3soPZg0kPHlWlSS2hdeZhL9XEn+Wsr1yBDm
eYCjCzjLN2Hb9SNQUDEz8E864WSpPeK8xqBFSTDHcWtQGdFCiYFrz/DV1ajA
QdxaTr7wLBxrIzbBtnc++MMnSP8RIPRA8ZveVDxB+zbz1H56g3T6q31ggRRy
gMg4gYE8zgXemJsPJAsit9M7B+Bi3kPnZ6vK0YBQBr8v8ZOss5ozztcpYVtA
DQgfTyJRQlOwbpLG1z0j79/AVBIYuj/y+Asbk8gPQ6Gx/O2Oq+QKIxX2eM9T
7edG9nUG116DCNvF0ue0FMEQq/B73yWk1ipoCJ4ZQOQoSKwNSKqk0LfsL1up
7bvrO9PdCvYAsEMnAGyGs0KQ+IbnvqO13t8dJ9sXE8wYlwdBBpgTYIAwb740
X8Tqqjk+g0cN4d1C03QiZB2hrm3pk0j8BSK9ZeVBgUhrJ+9z6Wz/KjObPX7v
T220sdAHrtrrcC2reFR1rfh+kleKwYKTCL5E0QibwCU29qR/yI/3dy99DnU9
Vtxy2gb69zm9+3PAieOdBkiFUnFQMt8m7fyS6heotHZpvgW9ad/US7/YWm8B
0FftoarALTD90GU97r1cGrWjGkYEVUx4iGFyQ9TQqwtXM5Ht8dng+nw6Z7q0
dPPc5c7T+nHQKxocxQ59Til7RgFQQ2j5i2xKc5UJqrqW5sWjw/roa7XCdrVQ
COL40/sft6YWiGJ/bRNs2YPzIP+rrnDVGF6Wm/5ajSUAjf0jMQfs0mO3/WDR
jzdsAWg/n4RRC5jgsFAXxZwfPUp/2iY2ORRDdSeDzwkNZ3uXQMqkFZ8LjB4m
FZdOerAxZ4O4bKRN6+6m7bDlVFJl1N7ZmxClWTOQ66HGMhtnxyTyDhVnfskA
Qbtw7rNIWL+cLwJs+I4CwOguTmE/r+e+FXKQ4dXUWIG1tkdNAkkCBUDlZFLO
7xV1Sa8u7AML/dCA6J5NLkbPh1rzDiAhMdB/mdVCXQqfmk7D9Acy1t9ZdokD
MHsTCskbvq1SXX7YUT+DIEGbbE8kNgXsAGF2KhHcfc6OouWEFVbhWFLyvjxn
8Fq3qDLU+Lqcwp4LAny5xeULu+U8qywzBguK+VnHBL2qXI5lQl00u2mbPk2g
DhWVWLlwHx5NBfDnU1Lo6G9yOjy2Tfwnd6sgNDq/v9pVLG1JDNpvbf3WLnOa
8QQNA6eNdi4w3DJIv59bOFCpXqMi0RlVsSK34tv+JVsojDQsI5J9icG2d4GG
99Im5KiVYLlsuwjtAb7QbeoS3GEo2SvuDxaFlO8CJDekyJbfZifJN1uzwtH4
Nwfgh3Pvl1dhJusxVhMDRYh5kfCg6Ml8Y51xAYlJcNsdqjoWdrfWM0OKhhWx
QZ72VIQV9roNZjQSyR89brOFNO579xaqn4fdApJQkvjXG+Rk1nYdWpVETU4H
SF1G1ehc+uoexV1jiIn8CxvoaqIfqSw4zHQarL4/c55/nODu0GVUj3mr8AqN
kn++VVsrVp+2Z1IeTfwOVvp0RKy5gkaQ6ZO0DkFz2kAQpP+OHVv36GktEssH
+vg8MkEngFihrZV8qEswSIX1vgL3rUz62ALpgzYpq5KcUn4U5htE5gjEi2A/
xZu7dDNo5RTIYJylyC5dAE9HeKYmLia3MHr32rCTO8Fjihvky3MkKMt9lHFp
eCSTSYXlm3d1fug1+6oCBvl70MQEjWUmJZMi+kfASAm7r9DLazpuPRXCU1nt
q0ZaxO4mYWRjSW0OvSrXcW4tZYV7Fnbcrcuu8XNrauic6kji2lGiIDU089O8
YzG/paUhgP3XfraghVXWGt13I5Hpolmqe4vG+AJG8BgyQt6gwIqteTtFyuPG
jEXPUoNXy0J9q2896/60H7PjgktXEcX3Y+RdhGl7jIDnMFrYVUZI0fWy26so
GSIyA3RtrWO69/psTdbQPSS2dME5EflNKDPTOGuNEnD7NmQTWFcKfFqBdrOc
Zx1U+B1CpV3d25TpqZ3mdrtAJnEKQjuZ9oxc/WdDGodVVR7pzDahyovm995X
bbUoT+GLbCc35k8r1VmJKr6eVxykpL47ub5eBhX/W2dKXnlnTOlohHJRvWpS
7w1Vjb5wBbsWPdZgODcyUTTIF3lUGlHBbDTB1NkteJJgjXGa9hV97MzaNxcr
x4/oktQ9GhjQgSyPPoWNwkYi+tpwyXMa+//YrmmVRwrDbQqfBTzQhatQxog1
ahi9OHQ4wr5cB4wZ0FAga4JT9BYkWuFly/hvbTOanOuhRxqOESc8YPX92SvH
EZqK1KI0MZ7hmb0hCjCO0HTiOku3t6RQBxUqkCe0Qmzc3Rk2//Ls5ftgEoMv
coxFbULH34Qi65DF0q48u2JbWARTFidw91oPROKvtj3eEUdabB8N65YHEfWL
ctaWaBt9mdNhl4NT1AL2jWs1x+u/onht/1eW2GZ33oBkIIkK2hm46tYLvQCv
qqRN5IpzV/jE3fU5aQy6nRTPQJaGLfLXwSiDX0J4Honn2h9S2SGmRzJsy/kN
nc4Cs1b5POoOhIgYeLRkmVG/gzYkLsfOkK6LHIrOd+2P1GEdaT/Qy8qigAp8
BsZxvgw1G1UtmeXuj4u/QLvLbPrgiFVeumCWCZ6gi01hCm8ZliJ4o+bOastA
jyNdivFkkadfAHh65eryK7Tz4gXuNEyQYvSsZsdLl9SdfLEOwUrA5L8FrxR/
dARYRMNJnlSgauHsfXEpMG3ZknJZKqeqiyhcjZpPIXMXRCJWkGSE0qowm57k
Gz8AfLjGNsDo20uEfnPhpj/Pt3JkOJrwCGNCOvgJxb0MVUpFXLITOj3MGYIJ
fJo6lyV+/MQft1eTjX4B9P50CBo+QP5zA4zLRRn310CywyhKbcOP/5gOyGUN
y961KCxw7vEjU+a41rfCo97IZfz1BGJ2mx0/E8/NP2fdg6sfHcfn6xBxW3FV
v/hOSZmstWaZYHhvPxd7sgD0R9G+/9gfCpFl62z6RkSyrg02yNnzJ+TsdPbH
ouVkl32IjlLvj3C5oY/G/IKxfdTbaanGQIGvvHKV0D32JbX98zrf+hOVU7qn
vOzPwhO8cjYtKodVuYzitXJcNUXFZxBCeBU5OugHBia3oiDXc948Cr+SRrtr
A5Qw4DSuK18xhiPSyYRibKNmB0pA9XCHh1IgutY6nuTIUmZqcDH9bi18Eg1z
SXlB5L3t0fzOcvtoAQStVNk4tmTQbQdIizxhFwAry+Ed+3vLAhQJMOlSpE6C
qjmOquU0jNNKqJE00mTZrWpwgKgN7nXFkHmQqYupebS4LXupigyxT8Mb7+zU
06Qc2ewu0LCOd2gFVjT1wN2irmUCWBby3q2470PxFm/OA2L+XKeCyZeDg9kU
CkaUr8sNf7EnoYsSke+1iKMvd6uxYYqO6c2bRTCLXf930NGeB3EIzgtY6DiC
wVbtQdLp7i2ON3Jkdcp0/LzSat0Rp7oT/B5HYi1S3r+lU+DGLtwpwjDjJ7uG
rco4/5FUwCW2n+KaAMi0/tq2UUv36tpaw0D/qDvowrFFP3QZrvkaacMhInFw
kB2BYYb+wy7ZWDjDpReCVR/qIGeBKpd8Zvg9jLABAQXvPLDRck51pyuVKNxJ
EtuoOChlCQ0HLNtvMg4QipSj2GFISGIsj08OnfCyjEi/CykGGizld85USlOe
nFMU1Xktq/swe1e2hF6J5EzX0IyoUaryQektw5BBTKm0COQvBrsPCH8/W3EQ
5wSjYcf3pQ5X1et4xXWKfhsOx8azJ19Fmx3gjKkqRD5HK0Vgoe2Xt5cbNby2
Iot8nFr3+rqG+b37ukjJM6UmRpI9vZrF9TQoNR5ZfZkFvmfnaoKJoTxJhPW9
fEIxidAMwWUJtboIkRgtMUj6vtgcWJT7TyzzuwvQO2RGipl2Xv8x50tk3BZr
kHDIN5ZHMWF6sOQ1ThhuOuwHirEJKtxMPyItZslM+r3zMLGG1kbcliCGrari
W8+UZY3L3O/+TQU0qh16FuqNP+nKe+DhsaomKqIV+/2mOKKMzW24ax2wZj+1
idZ1CmePzrepRqaAqk5ZrVfi9R6073qFe+K11TnrXXN/zwZjct/tH2JyHycd
rD0+YlzzI5eLYiq5gpt3L5a+Tzv5HQ8EiXq0F5WZaNr2ZvYGnuGB6zxm8d4F
XjcCEnvH7dFPwc21CcH6dqhsa57INeqA0bpFCUo8RIY8zer4VEkv0jTewO4i
XA08QAmGbDBcHIQ1cxNA4AwgDu33EvMSA+Y2Kk0ixa04oji+o/ce/+/S6zKH
GdtMUbQ/mfev7V9qPVBShwCiuM7G0GyRHxf+ivUHcscWguBMWZeX/epsZ1nw
HcN0cQ/FRALSEMy4oBj4CyAKrW2/9Gb2O4QQ+53O7LColGabO9UhwjVSzYjE
2ysTRBylWVLrdNS3eY09d7c9lgIsAuB4B5RvE66mAEBJnQfHFcPtMRO6KSN+
5vL85P9Ii/cpUV8KlzEwD/bVuR4Y+gItZQlirTFK/zojMrHeX30m5UF0oWBI
205w66X2efPghjPXbEpbNi0WKBd5rmpbVeH/Ao+/J3oW5Qx+XyBzEYE2bF2N
PjnGb9c4JTaBSdYhSrPrPTLtGOsA/o0adzjAj6GDteL2z11HPEXi5V7w2b4U
LyMK69bm+rWjknMFNx7RtpZsCA4Vm1rcQOQy9Q/hTQYgzH5Fw3d4JZiDp8FG
SotwMsVoHkFAIU12N4kWM7eQVCoLbnCWhh2dB5j6ow0fAcblZ5Ra5qb9zb1k
IIacvm/2syS/OsUId9/kE3E8iA07+IO+FgqEcTSYlGzL7ywnmlZ/u0VG2RVo
XAcG7nN0piogcUnGXJpiQ3VnZMN/Q+dP9XFTL3QL9UpESSXpHZbAImiqit6P
0remd0FKE1BsIWrFBeddEzkPtkX74AdCgvswo2fdwxjtksXbRgTAHaxUM22i
za63sPc8gBDqrJiMJTSXTkw6qD44zkt5O4pVulzu9SqVLTvEURxsKBgH/fC5
cmgE+GX8EbKvzhHN8zTfgLHTFxjIAFo4eG9Q1NU29IbYQ4Q4tJrMVGsV0Vx2
Jp7mg+5MokbzMUn/2r+w1t9X9js/Im/RaR1bJ9zu8pL8tcEUpt2bv2VpbZFI
m1OfhFoHuRHe3rCWyDaifD+0esf/3VEr+nwFduEOqQAkiMAnVekL3IXQ8AxI
nFaggEv/9L29pVCHxbsxpsaeMruZXgN4AWDRlABHSrKTVa0LmK5MDx9HWV3D
krM6D77todjLoNCJrPMdhPQx3cLR3YmOFz9QhXU/I4GjCXCObcrwhWbYEEPp
FpynibWFJRGKVWPhw2bSWAwidGvnXnKHgNbey/gFicDYmpKTICYn1IefY5MI
59lFJKvNU96Pl36vWZ7Ic4fa64moa1jAW7M5PXxD3CNWKOjXpdEJS3VPTo7C
RG8FJpm/D1ZszRgInCDDFajr5QHN6//FvdFDPr72fqc14KFUSAtCUBH4YhFN
YvKDq5Yt00Q0HzUo6fD4cIQL4aMV7A+4LN0lwxDAt2IS1OBqaLYSzEZ8t7+y
pBpdkdd2qEkTvIOIKLJwfA8yZxgw8A9iAl9W3kMlQDBbT5UNYFAnOXAht8xV
9v3+KvHs6H1qrQOI+3ExA/7785V+l9ha/GfnANshJ5OL0bm8Qdl321MjfDxy
VufuE3eNh+Hgxi6D1tdRijKQ+RScAl7ikaa86uxz8Xjd+PLhqA7GjGwF7bRm
i4xiJmUV6SFuwfFUgTt7bNAwbmcCQwyrTEz8MEMHqbkqPKbJCJfrAR8TuS54
CLFcqdjVpbiw62QtBqLGnyaf7WLPUM8A5Jc4a4fRUFdX+HZP9SnSkg1U9N1c
eRmXRrtD7MoyIiuIZZ8jQeslzux6RnNcx05oYOocTHFjFOrr46MBPhGEb4GY
FQpC2gzVnwN6OrbDQugp1F1AEjZD7fmnkSu8krv1FOTtfPKTWegD+BNySZHy
ndTtx7oY0jG36zWNEqjqF0vzX7p5uMRfFyERY7nWotQ/qpzqQPzJF97YSx9j
G44T2wKMlsNdL5XFFnBAwDf8whclVfp/6vIYS1nYsA2Gi3cTA6aUx0G7HH+a
B8cmYQ1NE6lygOoZAUnmoByuGbripwBp8Gaelo45I0yaw0n98PUrOb0NaZ2X
znAn0zO9PFnUft3UV8RYYIYR/eekhvzGnphsMElWwji5WJwGK8vCAp1UkCZa
/gMHjQUuypmKNGBmKr+Uu3axBV4zIAXn2mCIbzOnBzKso5HEEnP8G3bcPeMz
FNtIPK2Fgt2jaOTqGWx7D4MZoDp25wYtLp1QuCsZhtq/9z4pCyCcCY2t4li3
otQ1tTYI++8b2YLjcK475un0JOBqPS2ugyl5S24dweoVL7pwjG56eC4vrCTE
vGk4+m68shtiEwoTnQrbywvToF4yaD7/HNfYpZe611J6k6rTslIx7UPDSRlX
91zMHe2rjX+D8kP29CuguW5a//4TQUIe8d4hIjHMe4tsvczYiEkbO7afbZMp
OTFLKUvZvudatwXklykcy4xycj9s3oQP2QxG5KjTBrMnWNLLCo+o0V++ZZS3
1sT3AV2kotZfnvxkqqN1wIQpUyQDInXAUsSmu8Pb/SJ8az9O0JhL45kwIlO7
kHhKGgkpAggni4Vl49K0lj93s6wIwhFlBDWPsRL2/w1arcxFPQey5//+t13V
IvWhZz6cYHGEPfIowAsE9knX56DVl3GzaaXbiwdFYdpao4adZ+wWJx5OVFpJ
a7Ti1qB0M3axj3cNJEeDU5JLtwPAt6dz3tSWZ0vlX4hofFVVSCmb/R4Ep+Xa
jXGP/Y9vZ/RW2NJF0DH/VbyMDk321xfqquYYgvltaVAT1xThP7X+Ss9tvQPH
lUHUIWPRx1jdJ4Nml0W3Jn4/6efEM/+ulbzrICtVa/8rFgeGLVosrvmscVNQ
ZtDFR9t9u+BXlG+Y6e5J8FQSTZy6+Ks3Kzs1GmIv/1qmONCptKKI5D6OuUZ1
M4QAfIADxGre/cYRPycMwbDb4X9brl4caU1OvPV9vhIbAwU56DeKu2MaX78g
EQoUrmlkTfhGFlOsEeDZWCL7yHGpXbmvirJmfH71sbudjLwcMTBRQ/BqxkFw
UDU6PP/KQ/o3OWZs6zIsXT3TKWGNBXyu9uYE6rjw8ynqN02NYOcVPLa6LeqF
PTczRj/XN6Jg8beYQZ6C+b1vNvgKYLRRVR55xOqtMHBFBSBN6ImCB+tSKR/m
R60iEta3TvVIfwtXXo90ZkWOcv5ZCLC6b2FBUBOTncPUYNtR5b2fZAPazRiF
hhgPwF5tt3iWPL/W0q5mtqatvyazIv3YW8Jkg7/y8xIKUvOF2GXGtWSVm46V
/gZJgLr44SLB92e9iTIbs/9jJpT6u22Sgfspy+1+hRS26JkbTJr86ZvHMphS
6DIco5x6Tk5NrTl0/dKSfTcfpCadBE03zZCmqt9n4z4mnI9LsT9yZ98JwqN1
wT6191hReNYxg7R7LXCnvH7LBBvfXiIRZZNXgfmgakZacoELjZWCD40i6bNt
850iniZ4JttpZXgoM+0MLsHNXmN1FFGLmbj16VoTS9JiZIIKOpSlEZiivLqs
ryR1UgxRzQx62Gib6U+ihIPuS9kJoOj/lBNiETnkGVZnL/KclOwvJH5GtN1Y
5aiyorQzXEkJqeX9wcoKuuJs85XKpyIRk4We7G+hmQcMbhfoABeOnoPqpa2T
Fc9V2KvuCWBBz4VqbV5b9PZGGh4HlwnXAHmA7gWFlLxRpuYgdBnhygYy0uNf
tuMO25CPke86vxy1hyo2A2hGoaS2HDVDsb1KjFz6EpBuvqoAPu764Mg6zPCg
BMsY9vD1/ZMR3oZlq4HWDlzdfx5SLkZjalXxMWEVZeEkCVItvDfPk6CBgGnZ
iblEwyIDivxFDd6hNcAE11pAB9gOHrXEmcbka40OZLH6DLqjStdcN66PQr9G
xozcG4HjRPVu7QgeEZQA3WVM25xnQ3QW5o0G1xW1G0862ZdQiz1Fk2F0gIUr
dbMPGK/sKdPhX6SUK2ia5rR6trZoOptEsklxFrJBZDCHyVB7Th1lSPP2m8UD
tGw9VrxYVPL5rCzftlG4KqeIgYv8rImoCV9V23avKm7DM+42wIiEzuaCq0sL
HO0pcTNEdCfXZvP8+gHg7TF7WXZ987cBSr7c80NmaChQE5XnIXETSNMRlPBW
AT1iV4kOML8XufdNBsekRX7xhgI68i+IqMot+3HZwAoi9RWRo3FuTyVJa4PD
SGCMN67BfvbNd5a1n+n0z4DCsklx1DkPzIFfFpuOQ4YTiGbh/cHnrJHQYsVk
JoK0dnPbmosE0iIEwB3VbfKBQ7mlkH3DKkiNUqX4xdtw8ovpUIUo+nxDWcaG
hlfEVNubk1ZXna2H64X2vaD7P83cvOQrBgQbLh/YYM1hX7K+Az/SVpEix2Fb
dWdRcfmmTNepRP2I7jc6VOelrimyL23rgk92O3Ig7AyIZOCkegBMzSjcP9A9
//bKe+TvoQbavOeN228tsjpKfQoFfKepmYV+kbKw92NCnt74paaMoazO9ChG
XYU2wKsErfVy1rFA+IZejZUY19Kq0YIOTjSSPlDA8ZLsuMKa4zqOuploGa+t
90EJZQVbASMkIYanAERZ/jSdnNVZM6hYCXYjxafXjFueWRyo9JEnCUm7Jz8w
UQ/i1l6QjpBIwpfVc+9uXZ5wk+4MWONlLDMuc/UIhFtylxUb/KHM2/sFSpAn
0SKmodkoKc14Levuo659RA1dUaEaqdj8/EYbiXrZhnAyj2dnLlvGFHlA5muw
iMjYD0XeWW5DCc/DLXWLqkkBNzISqn/qQgCzB9NeWhJGVqxThjCVdTrGgpI0
edzDZ/nNba7cKVgeeXjY+BW8p5RJ45TPGfFsq0cMx1SUmaMQpuNssThcy/rE
A8gaDaBpqCxgwyTKD09y0bTRZm4Bh3Mm4Et6NzcFpWhOM3UsVabJTHUItq9m
rKXl5PKN5lfneRROJwoeQJK8VbKRzLg7nIIp2CFARPWjX+u0dh/dX7xgDWlN
xOXmfWGdFo8neh72AykIP6wD8CuUtwUMvVzg4XwCSJQBCq1h/dMgeZi816aK
4/1FxFzNHA6qF0p9FZa05+dPndD1AF0jbuvKuueS6XeO/ZoSJQ4k4wlDX4pk
p2M/vp3NQYgJKeTknEbYFaDKrMTeuDQsU7n3pvO7wMt2T/oaIkB8K9TJSrOf
XYZHVs95NTQj0uIw/nPv6GqPMjPMKo0rnfMh7N8rlxJXAZ6zbPx4WkMNpfwS
AJkHigMA/evx7oTCBKENKZeaAq7+2sTzEV9Iom+Iz9K2eO2G9g+24P3VEW3c
f2PgsPyHqeetESTR1PtXP4ae82ssWDNLpYRPgLbyfc+DEFJtRyzEmiTK3x46
dUUL0MeSnSyzgtA8R2uZ5vLpHCWXSnc9hFr5X8ympD+DNONF6UPZ1a1e31bi
MbGWdLWYIV6BFns5ClvMDUuln+u6XfrC5nGM+xc7zjWngson1hbfYZOqGfxW
/goQbyLH7Ra/yhKylEOWDMlw5FeiHKn1i4c8RKFuA/jKwmnGOFj155UHbyls
yH/20tXEo25w5dLOU4+X7fv7KHHlGYtDChCQ8zemnH4L8xQXBxlvSv2BzLjw
Tke5fe0sSmCvbPTclZiCMWijmTBFadJ+xV4bI66BNYZVk23/YeS+Z8WdNI/2
48o2wML0JRi8vQkNiLU5kmqHmxtcSuTD0nqvP+4zb+5MkZajKe150FuZeItg
B5pCghDnGyDYMZ4lwsxkmTFfUzB5thVCnXi8/1Th04jm96B2wq5MZXjnx0ny
J5QFPEmJ9ROX/nph/rlrGlT75YtikeCOXRF3mG/K5fKnSP/oZys0S7jAmxbC
Vg//jKl2DE48aJwz92rvyirWYbUMZPFYfdaC4bGQ2NKc7gV9nN64OX5dMwJf
xNhXkl81xj0kuteT9Bnycr6/f7prr5ewH/MhspneDp+kyIWCW6JWER/pZI1o
yPkXVq6Z2YkR70ddif/ERXO5YCofyCWvU+88oHpSujJesPDNCnegMZacJ7y5
NbofcIHFkbYNgg6lzIi3a3dMe9F4csprTP43l8ECMxoHId6Cp9rLMZbF8b98
Wsoqw3yzOcfKkM66nFTgDt/Nr7G+FI58VVLQYYQN/7PtU6u1vKNyFRwrG6jy
6ZCIn/RItvQcU84ncy1HAbzkvsSgVBeptxkqKnwMRgQCRIbiDEtT4yFU5AAg
oBPqTJoU8SjP/E0g/f+CsMGn97vhKGJHhygIu6I2/IHX6bZaDQsPALO5FZfw
bWYyU7B4B2WgK0wVRETzRLk/ORlXSpbgSgSG3bI5H+P4E7FYPjYw3BKdT789
PMzHOBLmuABjQl0xha+lQtbFbuPjiA9AnDjLsrNMqDRUP59L4nWrLszkCRCt
lUH+AIXGVmuLbv17O0BxqJnw5RTTEf8k1RtlqLknyRsNVbqnifyeU8MbA0Y2
axwrwn4kNkZT2wNmUWF4WtNdS5pPdcpb5D9Kk3gaF78FE4aYKAVOye6fNb9s
COJZD/b9eWwNO4R3YwM5hVAla6onoWzwLhYagB6qfY+oKJ7+cKb6jVTgJJyU
vewRMqYhdNVW18JX7Dnk3LDg7GMk8x0Q5nI/Ii9cib3JaupCNnBhnk48xrwi
n0TnEATcYq5k1H4qq3ViKedt00Ft+6DYsa4TO+jfh3oojTbFR2IrEFG7bBVR
8cYuLq33CEiouZwVgkdSYAMms9M3YTClffKzgtK3C5cChiF8xPe0BYloJWvF
qevO4p4pCTGZwpHi1FJYq6kJNYAlw3BqoQUiq81LlMbdSC3KfclpIHLKl9qM
+Cp93RlozHzLs1EkPezyXEjlZnOuZejbNiamlYbCrAMIUPbkq9ucPRUJPFEL
JrGr8IONl5cQ37jB6hXHz7TKpktJFMn8GQfekkO0DXRtwCYnTXwohZ1ZzwHb
AASzrTfAfpblQLXAitW/78O55GWDsLEAfzPqcU26jbs3qkyRmsMq4VvXMXjB
/AjJJxqSI49h2lpwfSzgZENS3HqYxqKLlG4gmoTuF5rE+Nqc76W+JiNr1iJj
IIYMlb4VhPFZYqtOFfkks5xkuL8M/QE8psToa2J5dsrdzzAvVCqZVFi3TG+F
iOTADcpeKeCPAZBsXd5Gshut6Hm1dCOCO9SoWN5AKCLb7XOnXXJSPPSwMLxX
mMacno2WtH8xI4iNLuMVhGpl6oj+bm6vRgGak+OV2+Ipq7zdbDyLK4D19vrR
3U2hqFTKMdDADGquxnSOsK8vULkMjzgYTFgzmtZOQL1uwLE7lSBmo3WGysuA
TPdRaMQa5vkCUtJieLTF2qWRHl5FSCM8GTq+dphl2kuPk1BecMkuEUKMIjxo
6TBtwQLdhu+1L40qh7DoyU081n5Hs5ji/g0dz4rE5cNCkF0CP8vK6mijQ3Fv
ZQQMJeb5MHuBhtMyOHF3mDwiKeQSdplNR/VM48BKQylH1Lb09umFOV2VkQ91
l21jdyr53s/jh4BXUN+k2EWYfuJgyA1Ac+VOoR3NyDzcYCXANAadDsJYJHPv
K+fKvxy+dP9qen3SsV9xk3FtUuXLi25PYQOQ5IW70dK+ncIzQ033TDXl+atY
h7HoSy9x9PkU2Efj1ydDs9hUhTGPZ0aDeuENJ5eDpew5PbmHG6qc8WihpIeY
u735EVnNMfLMQ5eMhUUTDpEWAnKTG+uoRJuybVk22O3c3zAaUXWFKHiwkax7
peDJV3lSgD4yVf0xLiNF8sWUyOePZzjuxNEuZmlbMCsD/Gq0E2QTpZ+8I/st
elbdH6FETpVUh0pvJ4P5/AoIyRHxkJA2T2x8opFawhTXlSKtvtf/zREnD8lX
81EEK6jEsk1Zc3Nf2a8vmMC/DmczuuACL1M0yd+q7XFWdpVlFQInePjkR72p
TYNxILJNE4xArFeMjlGBHai8iMT3bdCA/iVepOcmoitnkSNCHcLTbcOwc0Pr
1u5pcziuY/nnB7794ScqmnQleJg8UhA1WYGfn+ZSuykfFlQMaD6b9M5Ph9Il
J7aFgkkdq9oZorkU+TwkN1goiQX55HRny5GH4H8cr8X6E+ZSsrDyQxDttwZk
JL/1ndqwuI/ZmWhe5Yuw98ueZYuGgpnMqhwGa2PO5hCBB+n7KSU2jSn5Fzsm
SOPra9/L9IYBRq/G9Ft2sDIeIBU8M73o8w5IztFMOsujrKN/knlqnkw2C54n
Ka6b6nkuKe4pKO6WPnQ3VK2LWU2OjZxKStPqh3nS+2FaqZ9pMcpd83vyHBIP
P0kHmSm6/efpduKiQs9IlRGnnDwVNkEJaDKER5bV8Fvqur/+UoAXTLcd/DRn
F3XdLhmU3daSO99RLjJ+mS6l8obzHivO7yVDW8Up69oBYvhOgZlz1A7YTr7B
YlvXdOR89wnAMyKlbgU4n5vnOM5WPEI4JQPlultV3ERP3gTvawxoZw+AxsX5
5FivMwgzuXwsq3kuh3ywrRBvoYViMs8jVEJM3Q3icj11kncNcXDbirSlT60S
BZUzWSI+KVpdWgHqwXK3yH6kgzIgIezNmLyH0qQ0QwNoBIWxhSV1hVIoiL8g
5MEEROm+dwfu4euxGWkYV/rFupG7aMO/FRj3Qpb5hLur4KK7BuwIN2+gCf55
6Bmzd1bcGNYeGL8/iNODwLtTWkoF77nLiu+LQQoYuzGMm9OMuQI8xSvx9WJe
rIOcU8HpmpyzXoQhlPC0Jj6Za4MlyipwavUYHsdkIo7I5K2wkTnhWsi+6cSe
H3sVj4y+Nfy3N7yVMWkCjh1a+5PBqRjAc0mNgVUKJoekzYmaltldz9IUps03
zUVWtR7zsC4awtl79KpsRPcXaQSrfz7m8/0JdX8Yynw4wH9Lfe4Ht+Qc0aOG
XQhiFCKPtKtbahTXCcX+zIXKX+i38ZgeVK8iz4ASQ9DYIeffaXTRkqE9wd9q
+bbvfzxfsxvkldSpY7W/BNIMVpQqSlLzu+ouHZ0p5wSrWzV2fh6lAhM8UOOh
NWTwtVfbF+deu7Kj/UHXrMqR/PJibPzndoJOQhvRKBEHNuWZrH+E2HevlQD1
4M1v0fSxp6eKEn+oCqSXRij/X1LgN8NntCNWLKSLOKIAARkhKRJhqRbchpUM
+mIzHJflbHT3s4PZ6Czr0t4+bv16qtRXMs9m20WU80Vbj4pxDKhCVpvXt5KW
k23HS/ZogwT6XEzB5RS/K77d+CnRoYbFJ8j+MDtDQ5bcAswH+iyIJhqI8XZi
K+LxjdLZZcbLrijCRCTk3G9RJZU12sQHc7NmXrHm9LjtpNyEC1wxgk0Sg0/H
kG1q6/pnP3Vv/PMzAQTI7mdyXpXYXfGtYx0jZPglVDXDaXSJUHz501M/aScv
F4PyGjqFWSya0j2LrsGlRD2pL6Euvz6oQviV+ODAKyy9JXBuwGDurzJr9WzK
y08PGn9CC6M++L1J7IIRE4/ywqFw3BPduKoA632bG5eUzmY1batQoNGg8EvG
MU7n/Ae7qnkFmDiB8R+yU28B31lMA81PVlWzUW1K81lbWIHIPY2qfbtXB4cw
D/WY54VuCnsRXH3yxpvyaZcdbyAcSTcJfLAT9xyNbtws/P4/AKhqS/qoGN+j
NyyAdbK+r7ihJi3fOTOIk+wpLnUffCv0Vx/D9d1gjBGeLiaPs8IBqF/BKHRp
l7z8g7wnC8lt3yqZRAhw1ojojqBqJFr/oroKurCzlzLxVfx3tiNqYK8JFd1X
jfG6+mgQx1RPxuOqk/QBCR0UUbeM5sZA445nZsAtVBWNYhOFX3qp33hkRtcc
eOcQrzhi9j08f2OcDksFA2EDn5euDqnZAqxtnUJPlzjRFewIbTP+qtpFANSY
ZQDOyZqjS7IrkraAgcXVOHmHdYC1Mjn8Rqrf0AHY8d/A5JD0zsIRtkW9M6dK
hAhD4PUC2v6yuaGLNXADGrxLYu8Cz5akA0exaYGv+CzBhggBY+dem4S+UrE6
cfpFPpxQpUrT9TK4d0AkzWbRVmDNb/jrhTu0/q8hlReS5dGeus23X93IIb/q
ZIjoz1pDy920+SFbXJp3/8UxKKZ+YIgf8a9Om/4LIWVjJ+tGwwEJo6yzAFvL
FCyr9LVjixAkQWD6KIRqw4hNVaRTCpRI0WMtfC96iAVBORr+catF87w7FEXX
hMSMm38a/KflJFHQ8rCxyXpN1x1sDx/WspCo1WTeh1kRD6TqcBBGL3gW8ePk
HSXup5tWPRDdrfuK8vvacjQ7hv222glYrV015AkkeWty5BYa/aLM6FyzsFfl
7UHmdj2zccXdwDF0A/4j/LBtH/YEZSKxWfbRRF33L26NxjBGrB7DWNwvp5Cr
JDKG8419iGkS13C1Flyuax6ba0c55nQDGu1LCIHzUxe3ZGyFZ6GElCsSVZqr
b0cO+o1f5inkBWDyFUg03VJ441pLPEMlEEpXfzGfbQhSTvvOJhS6i6TCu5vT
rSw+G7Q3lGGIBp7EETl4nyctEPf/HpNB1VyOlxTWLUJWLsqAcr+cbA/8JU+A
Iop8x7TpkT+GDK/PYFCvBxwLoG7cBL583+JgBp2lpfIKjtJNJKwB2tH1X7cn
wbaD/Bot/xTzsbtoa9sA9vCdt/PXoz1/pkqOvy803xdCGDMN3obb6DQaJXH7
5b2W+fwQ4r2dv1TYdgXvHK+Id9qYHbc3BGpqC1xwlTfduOZA/wI1UwE/7OJP
5N2i/BliPjEr2Yc46EBot0sV+IaMU1Dz53GLxKX5CJGimo1FHZ6/JAMUtnuV
mZQceGb2poMV0BBXfzkM0nxy9ekY+oXtkOLo3AmJ5r5BLHA3i5iLdNuPZ8JD
w6yDKlukZgY3a2I6wAA5/jcvDXX4qFeqWy6Lpq07jiMk9m0dSDKn8g5coKQI
lFsrt16DV7ojtjpxOgKmNisoYj/ufJMif6yPC2Y+kiXAc5CzDch35yaRMHf/
0SrR7dmEy9yrucbvDFFvXPyaaE0HhMYCvK7z0BS3i9dglEJf/Z2cfvfISJ2p
usIHKQs33liweRnwOqEECf5tvfGad8IPwW98VSgJe5sQj89GavXJA+OF7oK5
awhU4dnyxP6ZHryMxsiqTscFGMIUQm+/MIcmLo9JU0gzf0+b+CW6t0fElZTa
1kGBCjX45jVbPbaxbdYbTgMsQsIBYLq1q0fQ+SAV75FyZmOpNEkVZibbMDrI
pEitNECmXTwztsfYm2dALNMmkUeLZnH7TYvuhVRkI6QsqdIwM3oMUDfjyBx8
L2kuBSSKzKX1hCtkWYbYGKyShByCMP3OMqwD+i2LcmQdLHerHp2NGlRnMmrn
vx3HCzJ1nSQQmHhyBdXYTIPBwdHnJXT7IK18Ynzl0hfzq9Pb96/Tp+kE0Hxm
8jE9ySNdscyqiEaIwN+vjYtbNXZ6wlmP8zua/79mDPR8/AAFFN+mOvt37rOB
YnVPkFwNQhTku2bdaBE8Cg+oub2NRECESm/VcV/RbrSUjB6+YBBXGJ7K//KM
AmevC8TpNLsTGSNdigvFtT20T0oC8E+BOnkTFTmFQ2S+PsCS5JL+jZ4kOhWG
2qWpNjyqT5GP/E+QN5l3e3MG/IRXSvoGC4Taagc9FkJ8jSnF/mXoJWTdGP/x
AbBr/Znmfc6MEkLFA3y2TMF8gxUJX531ObBMRk0i7nryLwG/5M1R6bD3Tkyt
zyuJLSlr+EAlj5BXMbeoB20Mu+iqLA06naQTp1aOBgUH37jN8+sgFdNQvNzt
AKSF4n0u/6ZIyMav3rgROJPfimDmcuM0srQ4oF9HKUqg44Z/Nu5MhL6Zmsiy
CV+lq6aU2rD8sL3KpPF+Wn/FtVuWEYlj8N3Yl15d9ZO9vYkAyFB+FlG6LrIi
IB+acaUbbpYzds02nSgGmUEQKOOXOU0jjeDpOsIg28xBIFwQgQO44xc2ZE7L
YwuKOPqNaalEhIK+5Q4eKs+APRnGiut8qok+PVLZvnaLxDVt9cdhTzYQb9FP
Sp+HZmBIRSyabNnIzcbnkkrrFlaITB+LXm+nBEMC0MZh6ncVdLEoFAz/xMbl
q4LbyPuiA1ScTngqhTs85Bcl8Gk9ToVw2L41F7N3todsCQ9GzyyurKSTfZ8U
uULUoNEK2/dqaNdsA3ofGxamELmAY3WL3rvDuUA10xzUhBIUeaxEhs9oPefw
3GhKoOMauIH/NLBIXxYYhDprELw+v6Am89PlPZSY5yw42K3HPBEi9Dm6guyt
gk/oVlaVyA/BxXzCo2BfFfz0KGhgXD/Vf+gFSvnfYQdMqLAuMHV1axzzVHAY
TE+fpl+nn1IT4ojP4fXulApUUw81DnZRVMxflXwLHBkVJ7g6qqfq3er4iS+J
knumrQ3csWN0Pu7zc6+83H4x5wBNzDmFfsrcJK48mTFOd3eTSzjNS6ylYpBW
28DlI1/ayeRBSTp5s+CBRzB4HbYalJVOyb1WyzF3VZDMFBHAviAdNRCubxU3
L5Xowhqrj7TyqMtrFo5n+QGQ4+q/ca+htiV+2rhoVleLNLkR38zH0Y+5mPat
zCpOfFrFvzMdRJEgLhlQSzWrGEoi6AKKsUjP8Bp3B5cdNi2SGOKHPYmsfsV5
lbTWU+aelUoH6QfMgcxFxHEfR563x4Fsl3+Cf0hz+cRdLKZRuDBpJ7dtYFop
/lB9Dd75OjO9oLtYELrhnTFso/BOg9d5XPSqQaclwQfs/keRhxy2HOpj8KBI
zfe19nFPyDe7xqthJuIS9cAnb5c4gXTYlif+h/9MkA/szlgoS2t3jxGVPNrH
EY43OV9sljpY/AR54QgZEcn6vEoYsjkKEFOQbH+Ta+xOnOycNjvJQdYTR7zk
1MoRnIwZwwk4rd9UeWfhv5ya9emrJDCr2ljfkSahWGYK5r2SqJ5U67OXNplk
B24O4TGzoRhiSqEwHFqA4YWfNdj2hsRovuf2ZqCuBerJYGfgQOIVCUj3X/7/
ROExFQF0WfGj7DA+a5YPX5WOlFCE9FLQWlj9xssE1ux/hJ9uEfy2CQ3Wcsgv
mpaDkQn5Qt8ZImnL+Ufvc6wX8ZU5R9kv0Z5Fhsdnlh2+kbPGNU0wV/ilN4sS
XT7g7dTX+OOkmUdKr5yQRW/tktDfiSiL6CZetKSFI842gUc8JDtTAtoD6lu7
7GDMol6DMPkgDLqs9j6SqQ2+1eSEzf0+49hgiNJSUvIGaZCWzUktRGxgx77s
gKCpe0jRKCVaexB5o2r6AvrnUPu0/tL/5RSF4GkSBeFJd5molsTNbusM8bUm
ZCqBe34zuGpR6ML/eOBFDASGILolGIoOw2PdBRlWrt2Wo3c0/TACLROU+EeF
0qCl13Rrp81F6jaSfFiuNDcD0feqK8hg9NvXQAYs5qEBDSPCNEpO2eXizRSP
2UaG1e2ji2mB+0qOHlaru6p9LhFFCu7F9doSBXWbtUt2ojMTbQu6q+ZvqYjx
YVi4j0F3WkVxIwrC2syMZnNXD602Ig4P7Fj9bIfaIE3Eg8h7rUhtt+OmlPUZ
0Lvxsnj5d47Ak2Gb1IJR1xSsmNooyttxIssHZvA40/IpWdYQBp0l8spr7mZZ
X+PXYY4+kGPrp6JrbGCg9+KpMC0zPsa7lIv6FkHQkKFMwtf0NwZcyXKOxVZf
TECtTH7bvAMTqa7aftaBCFT7YkxRbvAmoH2NekeqzIMOnCFn30uj7z+KTWId
LEqMrQpQqJ8FCeoTwuZ2BHWHKkGh0FUh1Mz7N9rxZ9YDYeF/wra1FW31v5lu
Trndm1Lb6JDjvMb92zE7qMbnIi1wAQzEAGPCpD8fe7p1EDCoSn/oO57JTTQd
2KaUmhWxgvEdFA1A1cd35pzw8kBsp+FKdJmaocHBVlyg/9Tw7QcPgLqcZWoA
XdYFPayxjSw/XKLSN9r4u3TAvG195mT4cyBEaAvD7LrUaOEHKzOlHVlD68qV
lgwNZFDF6ZN9Lzl6EbcyeMtPUFMgD0Cn4HetahnVACUgatLw3wBxfQlxdv9Y
3fK2o1u8/W50mZ26G4j/GJzBmo6A+mxmE+g1I7pncpuzurW0b2nuo2ER/+Xw
gQ7QMPmxzDLafHUCwHqvu6NRPGZH/oS15N2EU9WGHtYmOI4W+qCiWsBflBaz
iWbBbmDxEVGsZexKfKm/n611ZSUkt9yzpWlYZ5v4EQBeatFn0R4I2p3+izMa
hgBjH9kdqqbLtmlg5YdXXJjyvlfiB/Gem0+V5uJT7Jl7bNN77A8WM17uVYIV
eCWgvGKUuj14gMg2KuXwrukVEhlp7MgIdRJFmOPgT92PvJ4=

`pragma protect end_protected
