// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
E3TTnBgqTil5LBdkbyADRNY8BLSultXHanYx1w4vv4fJTjuIsmfK23OqLAzJ
uHwiuYaPE2eJQWt9WnsS5w3o3gk3gpdCafGPMlWQW5i8WU2Xv4t3ogDxOLcd
AC1cW7HzDRmIRDgWcAzs5sN3gSYCrPw++lgN58/H4ezZx1X21ZvHl+l0CG98
dL8ufEMgwfTa0rlfyB02+Cw8capn5JApc6oGPEv1oSgovHUkoddEVoNGmCUb
A8rLxZWBODStSB0IIHBFUBRmjeZRIOCh+W36prrDteHThczj1Sl+anViqm2C
mREMAFP+YXjyj2gAfTEfTA13iFRyr6oQzQiJ849ldg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
YnrRY/Rn04LtYbzI3ckS7O8YN1nwyolDthLm8hQgDxNTh7NcaYhQLnGzP8H2
zGLeLdPgzffnDeHLZY8US6F3ukjJ1YxAnEZlH33SrixK9KEmDHTDU63oJAbP
V96oZuUgh2tZzVrs+YOkfj+LfQoSaqtLGwyaRf15bbx5DT7azR9Ts9wvsNEa
qjUsXlKUbh8DDffxNtNdtAr2OUAmw9B6GuqNEwen4W5IdK4Y6N0RbW8a49sY
gJU9XhL8ZMTj4slrUsxqrKnN9YiMh9AEvMXG5tnnVa6U6sp+CqY2fNy2KA/u
TDqQGuTYLODTMgvb0gxVKV8vO/n4D8TQx/EIKcSpoQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
BRPx/807VOU4mGqO5g2xOw9qHNDODYsC7bb4Yw7NNueqk8n9xly2Rgo6YS7V
g/AOFfONm5EvRsSSLJo+ecaoOY1fdNNzdFaMaafj/Y0Ykh+YBydBeH1psR9k
Rtyx11Rz/T3gSBetlOxsVRBCK2MIUF1/P7bBrHZ3fYSb6NwFHtGt/89YrAGL
MWHbkyBSXfqB4ds6pPn23so1XmAIv+X2QZ8HEfuFtnDzt3FHPOT1e97k5vMD
qkTSk5ZfDjtYXoAu2b+U/QiwUgvyeaSicck8/8O62OSeN/IXS4lf+yd/FYId
kLrSc4H2fWpvmtJLBBzRWhVyxQ35vGS5L9hk0jjTDQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
J1rR+xW/8B3a5Ezwsy56O+WW3NE92Y18ri5CMWMMAHyPTnFbt8mvJI1eA/b5
bL8euN63dLS+8g3QL1KF7+VClcQLV2v3G1gKFFJbIQ/z2DafLgg9fk4Vjn+r
LQH9q8vHfy1rkYbhHxNq//4Xk1JgRa+5aulnU3bwOWc3lqG1AEs=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
gb1WyQ5gv6biMCf7bf2BhUHWXOmCxHkb0OQ8Q5b23t+7Hc1JLyxv0dvgugC1
XE3sGmMYR9kTrodadLmJshywSufqwycoAuQYbm0c/FTU5iyeKOSk+tK1Q2re
86auqWfHV8BqyXzhRp3acnNtg4rdyZQX0PVcwpmKf79Zll3rtCgjXI/1qt7S
kN13k6EqxXcL94B5ddxCQA7HxMx62KyJg4TrCQtJ+ScQXK6iH6g17AqgIq6U
1E84p0Ju/09vOHWpoZNCwLZXCNPFt84YcqsrQyve84QZjhwkCPTvy/DDriNi
ZIqDsimle6kKNeSvg9p8DPqMvQIjOCeCXITjC1DnWkRPt6SfxsIzig5CW++6
Tly7ajbQZ2ch4udweSBvL8eWtubAc+eAzEs1lA/zELsjt8qVnCiGQkOS989m
0FTDa574NAhjiUjU9fS8/YvGYaPd6YqGiHzOECots0qgsMyIPVtb3MQxCwRv
1WdxWj1QFgWZvArE60OOIIwf67ejB19o


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
YP/V9omBe8CK3iEIRv6t5TCTiPX1CqQ6O/0g/J5nv67kqqHkQSdTC5Y52FRh
55VAoiagyGhIGlwdjZIWFw77/kW4DGtzMn29pwHGBwebphze6//R3Wb64XKZ
3Fba6GgaZCHhUIt50qlS8QnkpA2p9/xG9oZKw9f2KFGrnvXLFh0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
L/2iEQbuujPl8xcXiWPFJh6UL6IIrmn3NBUxwQcfzL0TjL5iJjn9fw0bJX/k
SPS6MgCbfw/UZyvOhAg3TasVffVqO1k2/BB4b0TsLkNAiQc/rZRgK+jObwyG
ROkOhg+cqmxp2taD5sL7NmUBhACeKAyy5nqY73d/GM6xRJSrNmw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 14560)
`pragma protect data_block
HeIYW0RNhcs87bLbs+FNKSTC5dV8Ylqn5G8LIU+M7yJwEvRCFAFnI7QNtAMG
mLoa0MGLU0MV6+iRS/vo8M2ZG1U0+2evzYF5uHt2asp/tMgOKCOWaiqmhnsn
7YsnmN0R/TwIMkgB3uQkQH7B0B4BRMN8xc9p0Rts7/VA9621xEQIIr7vSGpB
uZ8ym1w12QO9vLGEGGM8sSHNnBCrASPmFaDUsSDfcg6vensYoFnB8fZJ8nJb
AfmAmVXII2BM+Mf7ozmHANpf7nvYfzMEYvO4RAkY4X+ZNblm73xfTASxH0IG
3LRrxCqrh4qoCfNXOz7z/r4jeR1Wwn+j1gpnhzj33gu+xuUW1VD+7cizxYNt
PTm7jw4SdbsYwM419OgzgweY9MSwmpubsPITOHYa/M15g3a9J1LIAn4ukOf2
PYyCsOO0DVilf59kQyNqopermV8x+OzPjxwElJL4pjbdOWSFZTBRabNjifDD
gXsQhOttQcrq3wBhzeVBcr5g+gWd5TU2Fyt5tsQeAwlKcpuBhp7M7AnVwuiK
PBZMUVfszonBD+K8EiPeWv2k5EdTSebICIZDYSQIKwQevj4YgHTgF5gNBPeI
EdTy04tDPWUSIfYQ11/YQw8zMbej3SnQyEqie9rhjYQIas1xUShItaEErGk/
aQW8nfCA8OzP9mg7bk1tk+uu7OCm5/WY+Bo9YK7dH6ZGmDpPRPC76rF4Jakd
Xn2COwDcaVas2rR40DR1B1/aSeawmXwIqMDMP1RoWcXNjmMgkVy27ZmjeeOh
CO1gEac51elq7+0bCd0VaMAx3E+2tsmpvU4bpBdiyXiCd5ikJRMIoBSW3+vW
XBnEQ9nF0yHdLltVO36F3tli81fr1aoBPvmyAKFaoacrZA9rH+jAuQF6Oua0
/HUVlnjzl8APySYgzTkmZyfFa2dkLNkEA5T6hcAVwwbbXnN9fUxWbaJSWmJW
dxBtsi8X7LNA+W4aHXLhPFJw6izo/ZCM8ftYZco1DbjLe5oNhFqRqpLU6omL
GIhAlOdpoNr2JyVLUUYg+0xNSnjWr7S8lx9BVBYKFK206LBbU7fTWTd/dil1
Ou5AieMdPLNJ4kCsLqfUn+UJ4/6Eaw5/GoKv8DDqB1Hajxa5uVo5APPCDGPV
pIsXBHgc7Djg3gZ+bz6pDmyn3sq3Lc19AjYUeX8TYxzaMqIE9gWW2Sj/Dtn/
nXhg9t8Kq3/e3u5ACguthysBcuCMXGNcAoIMJXT86RWmLecveHctuwVyrqio
ao/olbmlFTe7EwlyHmuVUV/+QmZ2w040fDNppWxpd0HIphjAWa1ndzZGGTM9
YnUg41k+TaMOXFn73H9Ku2uvX2Hv24ToPL3Fl6ovso0twTXzPe7xcAz9E8mC
KNy5JxCd5I9fZCPrU0FAAPEa3PuHEgY80gY6i56ITGoXsqbAEwMd/5d+rOyB
nJ9KvQrS6GeC61am/WVvnC1irvh65Iv9cqh/M5rQR3A90F0/B2+XBzioxf2W
fwm/L8i8rIFhHBcxQYRWXT46xf9yvxqZPREqKar/EYKFV6r/FJNMO0fXkBqp
GbOBXTg6fLrIAwwtWzyncjAzwqwyvPUBVEzHZLCskPcBGp8mAdIB26T90N4v
xhhx1yxL9ABbSz2Vpk7/EyT3+RZsvHRHTHZhL+s9/JT6b4WtnAStxYILCIiU
F+nmTKkm4HMj1aqTgDJc7qm10nWOVqQyAo2oV2yWWlnvzSsO/tVNyLVIP1eH
2E37JvU3JB6+Tc8SCffh9cpoozzRGYBgO685wWCcdSAFyejCvW6Zn5vh7Atl
hHg4iBBirOdaHZrVjfwRoOgT61ZZp0mGFxIkfRt4cDSxBYKeOCacLtz6sZs8
iTqW8ZKHfdDXTgv4Hn2UtinXUSU+PLnfYQULgxUdhDMoIuBulMTfVhkKLcjL
oMnV0nH01ASmI7NcAsl1rQBjD59UtzeooIeT39N8a6wZF76aRGM/ho/h+9Us
NFy8J2RooAXOlmnPwisI8BUf540LkOMobiA3haqhTFB8M3vrlLHlRoK5AcKi
CzcC3qHgwAommA2duUa1RUMr41PBEDxFIOnauthgCIeU+S90qty3Nxpp40Tt
BdnNaHnyxprB67C2koyGyHbZ80uQNeDdfEOTlzz73I4Y2ZfyPTrk8vgvv1s5
1PrZQXOfAfrby0Mo0XtSq/gmq2fD3HUtWiBob7jjuxVkv57ijW86NAUCxNic
D9Hlb1nss6/+I/+uInF7gfBeGkV/BZeQei5LlmK7uivJuAsoN9rHk+OGA/Xn
mwPD37ru0Zj7fsamxzvilNpoD+rObRcTZjVcCSzLLw8DFPpHrrkhEU65p+J3
q8XFpPKAN4Cc+xoFIk3WjuvQYxbsROBJVN/lOob1XVvZZm3NZDNG8eHf9z3n
pwb42GNHiHVHbUgMgsyggvZA2MHjAUj2zU5/bUdz7ks4nk2IybhiCHvwxG/K
H4S2Y+WKUKeQmFBmC5LmrCRZ+SKjZ3zh6rY2FadLEZQbLGyVqWGaKSaeoaXP
woC1oRek/WTANygsJ88ysmp03s9Xp6v1EJYF3rIyYv1CJ51Wfx7lknI0eXGH
/FbhixDmXKw130igkMS/8E7jSBE3rHqAvgc9h80RJajBdwfVCkyhal3g2vTu
+bgluZJkkhjrrGkHWZZHPhpQhgvSqCbzJVj5PaJnJEq8fAVTUTDWjIjwDV2o
6L0DIRjyihsSDqbEc8yrNjzo/hPCn2+Z5KIspj7amrtx3CkmigLlx5+XN1Qw
kVpZ2XkYhNhzKLNhBYmvVbymw3dz6QFnyTk07bZFCBaroMREuj2s+99Sd5cU
RZbXi48mlW3jN2BLgVDY95fYpwaKO2aYDp6eII9t694L7CA7EluzfBJYxRgT
28ZcbiJGkZY+HbUYwyWnmQeYdMfI2FzquGIedADWKlkkFlHuS/yHDFFW6GQ3
ZPHHs7Pnc8d+OPBEEaBbMdYvnozV5N5QrWT2Lztt3z6Yegiogqeik+iPqaOC
l9+otFs+LOvEB6Vne9TYPLglfsBpyNWCBKLuUJ0hEVKQAoJoYV/68Z2SIGio
Uonz+gV0lRTggxdgogb0PZW9aCo6kVNh64psZLMrtw6rpqR/4j9RZ8/5at50
nuTo5LnM+FFfI1l+RaOHR+LWSgjicvzs+8YN8T1JRv63/ijuFG74iBtVDFKh
8MJyFNnYdB8Frksko0CqW2iFvSb1AhSOI/3ejhEMhlKsSny3UGCWd2MTy5or
hBIZmVh4449atYB8ENFp6EmnemeP7uYDK0Lbu3GmFRSqFvOCpThP22T1/p4P
VYG+SwlIVtYzG6q93HuhMNeFxbEPp8YWsSTsYOswHrZXLIWSDhxwUaD7o+pX
LUoifJRCvWMq8wc5eBtt/sKqqZkmSlhZk+PSrebQQHEclEfp6cuDIJczJnA5
gHSGWIXgpjwUvzxUvPcd4FP7VfFxdoZtRlt4JABVslbqgu3V6hR4tJsB2zbJ
CQzES+LvGZplA72Fz66LXPk8WpbPez7a8ptzcEM4cZYpYcZNyP46le+chuIn
iDKLf0/u1KXkqfq76VOFFeiBHUwwWFhEU8h4VEWvxqSPHEHAZQ5/fwrWUVnd
R9zdJyAqz89XmrKXJlj0BBOPDilnNvzAqoq/lNShFIYZGh31LG6w7NYq9kD1
8KLA+L6/hpgpvCDDY6oiVOTfGtSgmnDoxdmVPHVAlZwFnnwfbSNYu4r+iSKn
lX6i5zqkLyftxrKPMiPziHKbTTgswbiZugiDRQEYuG01JcJt3PuNSqBx5Bjm
wuc02i9frSbb5HZfxSd4aYcey6+UmNK3OtQQmTJKCG+qmmEq0fnK6fcvdj/0
aFNuEVNP2sguktGxkeDQFr2nrm0YgaVozUR91eOkvYdw1droAL7F3yqT0pQi
bGcjki3d7tzXUw4/7FMc+jYzyUXBhN7GfMoBCfa10om2imE+ze99Oto7g9pV
VifpXVEACWt22IZBxtnbVE4fT5xMnrP8e8Wnh0bqer0Afz0VIUdMJ3e4sNFV
vXGe717uDKEoiHBpXEdcHCw7g4FcJgUq6ryLd+4uhz9qWN5Jauq+xwgbnozv
2N5AKTj9MdJmgZaDlcoKO9bU0Em70+RHZ92DsEMj/VbBUSFAfiL4EJOFDoxd
knu6v9jXTqMrMVxZzW5r/25aOc8uiMugKd2PQgaWWiS20wzKrfP6Me/xr19N
lLKISwA4G8H366uZLI5zlVJ6U/6rg5g7KOAmayQQih5oTFSRL132jX28O/db
5BU0594ZOmz6vHFp+EF9bFROVwZ0+KhzDKkKqDj/Cl+kG8jhRDb/RRyJIg35
q+mWemRkuKCP2ce5D6rTupAsBds9xWBDbAF9KLIBRMnJsEuqaEkmp81ARM8I
uOqyZfiF/TZQxVRqnWLVUsGz8dff9YNzH5tw2GlteP0LrR6LH6jQGCcpAR2Q
nBQBmhsK56TP5gsxMa4XqXZlD4IQ45g/fl9ZCA2AfrId9W37I5iVHt/J0xMC
Y6n6jb8ntxly9ic6hNswsq3ikzVCtg0dUtzq4wdR/H2vwP5rTGiSQINUKRVS
xtmwmVn0iyr9HEczntL/4ciy/3OMlojxyVTCECypSU4xQ3ph9TGAVT0wmP8D
BJmtMtTow6QqcYTMaD3f+74NkdfYCFL7Nd1HkHcrTRNLEvpnde0y3VndL9gQ
ETfCDs85lVBGCVDb+NrOlklwM7+X6XCU2g1yYHIz4iBMvDQvNMmzt9vqqzTk
GO3UDpwsbfBwAEcQPhvuaMgq53DL+VSKDRFIonHYD8354j8HeLVOcX2QAae1
c6QrJt3TsXVzB06/j4zSy+nwpC1IY8aA4KLtPuaxw2Xpy9sm5osKrYomW+Nk
aOKyx85VpACFYBP1tFn165DHxfTiE7iU3AbjAfFuhRzuLxh5Z5BX8/blrrl+
/A0FRkD0fmIMT1MbYmGAf9Nf3KhJsSgsclHeTmWGuDlbVXgfxsE92tNMBVe7
TDWOHc4mC+KcmscupJeXvxGGjUGdZv2xSqwYAVg/IEGOQniSMjJYTUsk2ODM
cKNlwsFcc6KP7K89QooKEGjvGwjEpNa2rDnT1WbaoOLR3B4NaE2PewNzKG+l
phVoJb37/DfenYrNDp1squ/J27rX7htOxNbbenD5NqlsBtXqd6vb4niZQROW
1jvBAmxUhOMqmhS44TLW0yS3uMnldYQCHfWxPqhjUchnRHaFu8sVx5KseuS5
okzIsmx+p7S0wlqQ0e4iIJay/3qAFqVnLXsKJ9EWzcjDNTWFhAm6PVSfDXPf
ddWLgH+KXULJRkkZKrXqAxGJBBl0K5TM3AsjJJneY0wp8rFDktNw0SXyemKx
QmpgkqQ3dM0rx/ynoL311fy9oRQzUfezdjq6Pv7Iy9BJxUSBmxGF7l4nN6Vz
jQ89tM/nIFH3+j8xqTuyX1nBKDy0hnO/C8wY9vZTxSDLUE3cT5cR8n3aPfee
ceXewQn1E3DrmIx3lOMdrI5/XG9efGIqEOMbE89fhaIWmQfICv3kHNNs7QbL
kDizFCemB4T2KUqjATjBFvZhQQPx4ikOeW4emSAUwqsqZrSoRR2vgbW3OR9Z
c7ingV4FY1r9esiI3HKm+PbZQtzMdYruimAZ22kesc7XwybGi6yJ37epBXOI
f2/K/vFLwgYsdaVA0OAj1hmGXpmDbDuA5mk5WvHaYxrWPO87/yJJrSm9S6uZ
WUSIl8OklIe+G3pWrlXhA93jXajvPbdjO9kED/y2Hc9pTZEXrejX8idoKIQv
X9f2573YH/YJzpkdG6TsOHCxPKwhLOufiMPD7OQ28SV479AzntN8YFCHbDgw
vl2kBETkPLLzC6GUca9EDLPsouQQeuZ+R9qJofeRchfUi4vUZxtNX2MrK74w
rHRF0qmd6LqCS/2rUewlIbn+MLCrVqeQTL6TtZUhOL6B++Ag79w1LAs8tT+W
EtsYSiPq0XnkCjSPKdXysLLx/w0/ysB4Kwj68RDuvcLIpxgNrZLbCMZsqQYd
FO520Z3Ln4VqlFSMCQa35QslBAhVSlQkRMPk9Yh0cSm0v/PRpp130DA9xQtX
jekajNr+26p7Gi63S0XQj1uN5L7nbTkdhrblgC+sBF8hoO06elFIkrJPfdEB
G/UeMW4fMXrCFfW5LgkvnRbdHttngl1QNhx1TMwPfmq0nN9bfWocT7HoPwoT
2KOUs0hSLggUaS1YbOmnjCivVWA68y28IGlkihP24N3RqCNiyz2/3rDAGCaT
XQUDWu/2oyyu3I5UVBJ3c0zZE1HjDdpVZ4qUGCSRtHgbC/3MBFwU4PitBGFf
J0O4gTnnPoB4GNn0D4HiU1Ve09a3qmzeC1k/WKKxWpDP4rrOOOgyz0yIKMQY
t5bsECKn+LXYjmY/0rIRyR/8kEkmq0eYAYAtqXapZvIyqZ5OX9TOTVEAB6fn
8esugLRhO4/K5COQpxfUIFXeo464GqKG7VzCav31dfEiAAhUlwTZZk1yNLT+
aqfGB2muHStdHa3EDxvBD1Egkv9FhY9VOYKlgbBgmzebIvhNV9Bli36+gEJO
u1ioTJe9Ar40PtWWr450QM43Gt5isxvB9XDE+odaZqt5qohlQC4J+Bf9Zse0
vmah4Kp4i4we0V1AA+lLskb80QLETZmLhDOMtRiIbNQP8dZn0u7DRXcDba00
DldsOb3GqCQv3r575RSfgU2EmkV++8zH9UhAi5SSGonkrczxGy1h8x19JIq1
IE8BHEd1pOF7qRXOSi7m9/NUcN5P/IzixbnRF9dIOhF62rLP0QtDoaIUbhRF
i58OmJS8CZM69XBbl0VkYPHsNcVYi/3YJQsx/FppCdVBYmYhuQHQP71JChVc
Ava9V7NU6ZU1M1p+HRp80QLr7StKxqDqPMh6qZxSKD6+blPtvCe8+UgTlHYu
vH1MlKQAC8kmM+gQcLV1RyPFjT9Iv/KeuzSvLWBXVWf7YloipVxAHq4/CYzZ
ZUZFFPwuNeDx+bMjjKAFZLknc80T1iAOGPOdxdy5V/diVib4QZtwo1QwTGDS
/B1ieaAqsdS1JvbDnFkPt3ppao2bWaX76dwFjO0Wptj7SAVYC8ox6wfE5Hp2
Uq3EDoKk9QEXWnE9HSqTdAoFwn0SDN/OqAYhLdkIOj+Boz4ENL+yT3FZyBlS
DBDyK8YVjS/RA0AB0JBbMIfucGK3bisKlQZlfLmf5Fi5HyXicf/4l6gEI6Rr
ngmHAwbzOq+LZS/BaydpktnpQMi9dlk+qNWscWnf3fHWiWwXwJrYt3zy6NVN
dTL+m9cjWW0tXfcqkJJ86E4y9Zd5KIKZyzw/QoU7PstiG93H+L+hZzweF4m9
srlgSmq9sKq9ZklsK6N6EpW50mRpUvtpwMWs5HocWj2Yj6mUcIv3SvZTT1oB
ULkrGbzcEQDEs4m53jx92wTZlSn33upKIINaIv9DZmFuQ1GuBD51sphuMQAW
MRUx4h2lWRj+GJMQWdnlGFpcAyKRmMXrFfXdAXwoWBtL/60yBZQChZFdMgCc
Xa9GzGLVY2uoGXzNySMGkJIfINMZORdxoqmG5RVuSJiI8rEXK/0cFfkwMCiw
v25vnGXzaFTst4WPdOD2NhQh+I2aeMwFxEMI6tXwMC7ty/23VrEOP3CJ5VHP
Y5kjvSxgB9W+L5XOPJVk+klhwS0e11sfKBuLiMqiHT1hyXz+9WqLuREbmvbW
AdV09ymDFQe8s1IG2gBQTJ51aoH8r0lv9At0rFu9Raft0Y1Z1qaHJF6Suns3
0Nusg8CbhiZTf4j7zWOAnnG8LGm5vMyE18M7WwahgdZAlSJoUCJqE8LWDR/1
DQTz1Tp7fh9pxqaya7aPqUProzfka1MNpiQ+vVZWvZ4DGy/TubEYClw96sQV
zbVOVjmoxhcMi5gz5Qq86zAlYWDgaY1D2J9eP40h7+rNt9i/6CNACHPV+Xvc
RVcdgIzJcoQJQ2ZHfBiNPpjj3+8CcpvVh2dA4BagbBX4QZIIdHxc61HVVmcd
pAD8zhX7LORvTJveTOFh+1FmR/OO++AOBjggUOxkcu1WSuFK3JR31LNmYQp8
9BlW15S3+ugEhyc6uHKiSpOASyQnAIyTmAMkJR8IFn8Xg6VvXtjQC1rfSWD6
3TnUCYvwrnRssh1eUc5/rJ7wH9o9VGuy4+wRwcjsVQECVirkEqNIGaa34jYM
Sq+1td8gtcSrC2L1UhX6YC2uRZc9Gu4K9nOCK4/s5wZHoOnLo7VSHNZcdnk/
5ESA9GieY7ZRjXpi4EdsHpPi4vasQW/kxzp5eElxv7cbzZn6gQ5QfyFcMIF9
a93WwVQoiCPeYaKB09EsnBrMiZYdcHKf11CO6JpcGyp2+hftrjSkL1wSfRQi
3bLbaTTQW7CTYgR4KSa02LRSNPmB8jvbLJKETu7VP15UAHPJJG0Lck0KZRD5
bpzq9WiMNe2yZ8rodU24IfGMw64txNhI0HD4DOBMrKZ0+ESajIWVg2ulAr1n
g4Y/u0rzWU495SQtVbud0NI3R9+zmWn1cOtnJRXOB92P7PJbgG9qKTuF4Evm
4HYbFbTv3w6AkL8Uq0Vac9Ucn0dPjnswuTdWrn+u8UW/hMxdf0p9TvU1YJV1
Y9O+ZF/UTWWm6R4Zo9ulrbWnX1MOnnz6fJTzVF6sspV0ZRObi8DO/t7pOo3n
sl32kex5BEERo8ushjt1nsANOOg9Tt5ZjtD9cxl6vzcOM1BW2YyDIGa3KZ7X
1h6AIH9SC3blrxdj7lfSSO5M4YNkUSOo/i+E6wwMRn3S2QB0pIjtZrOduYY9
yhp5jd0D/aMAzQbwb28ZITsewPCGf/MOyd1rtWCMLQm/pIpYgXedI62ju6Jh
BD0kWtCl9Dz7PtkEnea/rVLMu1xKQgpVoLfFWuGS6hzsyI7HGu/9Ez0NEaHp
dSAJz5fehdlq0XX9ANGnwSR1ucl6EeZxwBgG7I8u+j766svykIeARuhsphk8
nmNOA82DyDImQ8q1MvKRGUr5J3S8TKt3a72wcX78J7QZik03s39MqfTDExx7
b1Xt2jsE5XC1j2QmPzmieBcFYOstS36zRlgnKxIuHWyEgDa2BnUYgU4j5SLZ
79MiNUaxt+hgW+6J4HuDvCyPKhHUhLudCcj2cb7Wczco8OdmHPY+ieYb9+64
biUh2vPnqoSEJkByI+xCw0IvLGTRhtE+8HKaBoeo4Eng1VIkSkMdcHfsrvub
C000HXeRsKCfgrkWJX6g8jo/IJx8O/Z835UW7WnW+wLOGVnMtSQJnOe4rz7M
deJxwRDomc0mrGhuSjCUpZm83QaxNf5GkTakYoLJ1yrVacLf9w0tkLR0AjWa
kptWNDv2zgosf4UlPhoLSS0rcMIsmEZ+Qyyu6NI0M7xXvN8vcLGwuWIk89uU
mJ/YPy80z/1u4xc/AiMV7/6p/+baKzJx+CGLY7uFNX0jFaVOQqqicdF5iKjG
1xc/f5SHjYmqOKPULbK9nXAGUY4JIljyN87WkMOh0r7q+zMgK1nHME8Z0htZ
nas509cqg2tkepgccj6ehAF7jDryOpSbZjkHPcqyhuuHocGdpBtEm7GZcjdN
am91fnHfvpjw9lRelRp3zaP4rbNYxop4FnrqYoQuYTdF0mwUw/CWdMnG3gFv
V3R2pjaVYelLgJBJcGUf6qEDDUuemaJIS9RHuTyExne4KnWyXNxK8yHr0CA5
pa256a1Y4S+1G3wqsCXU/41YGribmcYD1+g+/LJcv0RmlNWdjQaYK4WVUoXs
iHlauZfneVuPwROs0QJoYXkmRlwyWpUK5sM8FoHA/MaRwlcflnjEHvLeTufk
WzckqI7k7slPU02Y9xHJZdxjhAT7IccjxN29yia+5lEN9Zjtd/JtVPtDmPTM
RuBNNpdE0R5tAULU2FS9nCr7Vhny7owvMWxIg1CJDOMlzxc9DiACKfY9m2Be
ocBnOHqT1answNsAYSiFYNBNa+eHzgLzml6jkl4fBM1XPRB0ZECEGaubEnxC
oSYsKUr58mqyreHqnA3apC/UYV5OMFXxkHvdEmHD72smAOWdpNyj2Dp92Hv1
4UXgbQekwt1csLGAvi4xkSYvDN0py01D7D27FsDJKDpjsm04epjOOAPs+eSf
XMz7Djbtee9wczfp7vIPyz9YPKQCKibJ4ZRg3UX/ygGox3gE1A7SNSiaygp4
gBHkk56z62RqVGOJmUlCL3klIyJvIrMisd6Syu4e2hE4ilzqhuOw8ji02wQp
8PglC0Vx4x53ew4tHNlKTpV4l0poISGl1godOSmA0XzegSrCn5RfpcQk/qVE
IG+GSufGhoxH3TLtf8am06C47oTY0SNbtLKNpAG/Ne7wZJbztGnJKboG9my1
gL58SUlNWWZXieVN4ysHDKLrLE27TEyShLxtHBAD9U1EiEL7scdF/u3zMVcX
49lvjtsOOzqZC/adH2M2J7U2TR6ApqgMCgWU2m6kI6WDFhXV16HQArHX24Ut
CExl1kKWNRaRMjr6Tb0LnFjMx/xIcDhFyh7zD+F48FaMqv+aMSPHS4/6XUWy
8gkXeS2eVEZrVQ8vFG/S9X4wCPL8YsdFbz8ueq1hCvPezkEW0fa9SqmlLUrd
+ZR87dAjJU6fwt9Crlidv9yUYxL/PPKbb9yg2ZESAieoa73KRo0072yPRYah
gOYn35HJKYrDNOB8hu1wQHVhXx+o2d3ZD1uRXd+bnvQmhNCNm9XMed29XJp9
RkFdNX4txTbftyPe46xIhFoMsZRGFgRrfugFqF9MBclO2ObhoifH9HYeyRMr
Li9imBWtR78nVOsHX/NuY2aImW59CK984oCeXoGESzR/wiRvBH4+YQvYxFV4
oDeLfFJ8wQ0o9QzIyYZ/ZDsgjN9hLYBL6DJFeTQhTGbaotOl9FgW9MNmBY9o
i8KScXXtL3dRhb4MV5na8O7lFTZ11ZAdywUK+xsg02oAmsIsj+YQ5tBtmWH4
1Y3hx+kMFIuPtUKLdqnFiy5X3BU250L7XAQyidjcSPKzgvUMM8Bt9K/k0yJE
baPkgF/zxw7fwnrCJUQTp3CZQMAhdqsNC1Lb0nWY4VzjNFktw1kNG+/wO/rJ
mRqzKFxvB8XvZ0rOzsQvz408nyxlmxSZQgsposSEYs6rRxv9dS4L5+bfG5Cw
16STwwdG8ci5zN2FodsE8PAmeakmIbVz4j/bqy+TSOmPKIM5XLo1z13INEPR
EgxzFfHKZiEbVXaYhSdotdAbOgtfzcBwHXwrLBBKzQ8ONDsd1/6mnn9jIMCE
5aa3hN/tnLcQ2s8RP57tw27J5zslUQR8ucacSXT0PsyGsYODDI1VmnlB2Sdb
2EO9RAoEAYsKLXUkx3h0Ib3vLfk0ASPepmLBYIzd/gph+djkZx0Ur7XU660T
c0nsC6dNagpKnCF6eSHLsNJJw+oVC2raG4kMth5Mbf/FWueWY5/HzD9G/SvD
tNf1A3Npxs1TfyBrl8o2oMgUtZKsgbjK1MpOgwfuhLqwo0ofgYN0EBr+1dPO
6LQ4jmqmGHXYjV5u1scQtxaDVQMzzv9WyJs5wcV8CyAC8rqOvF+cTLCo+3s9
CXOscMMFxIGr4b6LLy5b8qcUrJmRmN2ly0cru/noxyvj1MUOstp3oTQfkHEL
VO6ZvWcQ4GFdGq0Mj6EbPw1FhFND/wtpQbtPhs/SUzWm5ZbJ0DTcvn9FsArH
qahVwstmugFSdYxSaED4+lDAf4t1Uuj/butmCqNg6yFXFnigpPTdnCjOf1ym
zOrgaug9pTl3GN/+0+j6uGT+ckDUnwwtRaE3sPYoy/henicEfGyuATjo6rXs
7O9v5gO9XquYAWbjkO5ps3QvOJGfE9gipXlZAwF4BhTmmxjUxW01fQkRJMJn
9KgCskffarTM2pbSx0lXR9imBibSDSzS9FHKbPu8Vtk9gq41pZsyzJdtWtdM
uoEGp5SWu51ql5jIvcozefm9uCQsydSjGd0yCcqHckEvXLCgNncYd1hX/gtg
n1gRYPBl0vS6kZ3lPLP/9tY12rpMoxZxvNAc3iXgqNHrIUU4UBNtbUoAwrDd
2w4ChKRxvI22VJvIgrSw2V2bwIB8qFRpHhYwrSOKTm2iKJbm7buS1Gm0GpsE
1lkk6nmrK9xkPTMKQEWcM/9gvsAh3yDTYgHoFbQJ1xqyiGvKCEOHlp9rfR7o
K3vZ0f+oN7Ioo6hD989MpcSrJGsBvZYtvxMod8T+/dMew5zcwIAqLFQLK5LI
4UX9FURIKA72LMRuxxVC2nb6v5IQ4uNC7XERPdJKmBUWQHkgZC0AOUzXZh/A
tCLJxLz6gP3uaSrpKYQ2fqdg7x+khVDwryyndzDsonj3iJxbzbKaqxTo0Wdq
fNRmxCn1N1xfJksaEn9idavcw6Cn/C+nYk1y3zEUc7v23ZnubWi517lIC+NF
pmpz2lM/QaSLC9EvQaC/89kInll7o4KN9YJsz4LmxzQn6F7VIuadehKuN2OL
LHjbNipDeSE965W7V5DXkRim8OfFLCbFd4SPiSy2eWHhuMlcu1B/N1IORXd8
WCEGOvUZDpcft0+jLXAzvHCBSTRX1D/QM3FdYDeZAHAYbk4GoasoPHObWAd8
Ph36vnE+BcPjKSy3LWvgmKT3cZMLmhczSnTsr97caXg/209o0US1uQzXOLC4
v/wn3njpG4WntsPvaYaKO/piw2+3GFF6aDaOf0Pv4Cdgr5pgZgQ0z2OJuv4Q
nDKYPtHExqCKnhxcIj6UnfijKP9Cf0k9Ty4SxFBjfnmoFx/avY6D40tlp8Bl
SDgYgyz3jrI7Aq4AxcmlJjWMpJRP9W/HqhypC0bjtij8Uf7E2Q4Fw0nJzPSt
QTQ/BeOwRfm93Lc+7dfmugkG1RQPiIbz6hoEkKyB9IFe3dot19M6r6NPy0PP
8SI5D3dQbiOrGirHtjvOCMGgkC1uwTq3U+0N8pMgHZ0DWgMjKssHUnHd9gSi
WiYXJnHpm3A/ua0+bAGbFTY8jmaxKO3tYTyNmeI5RqF26X00c8DoW8ohGrLt
H2+QVrUM58rpE3UBrDu+bN0AgLzbJhH+v4c5WlOzeEw20vd2a2+QthYnN+cA
f9syJPb3gaHA1s3xCEQ8OC90eV6ceO410sDMbPy50zNiUa/nuRZZkcA5gwyq
SsBd6HtG9wndi7tzHHrjZ8btEayah3Zqt0Dk99pEeyoNjAvQaCw8ZJruUZTL
k0Ah9jlVCvYTKXqI93ODdEmUmjVr8NkhzoG2Md+ugxl9xgzX4IOssMnLAJDQ
q72Lc+c0DqrrELrE8Rwcl02O44ZXbXJcAbqwYGyagTZ+zuhyFjMBqWAkU8u4
6xQK3b/R4QZxf0SZtCunM98tNzjmYJHRgKb2FzGoS7TTLqcNm1Q7lWPrPVm1
o5argu5Bo64tbX9UBydHEsVLfcxM1y1GOVziEosnbnAIvOOi00p2txTFk2Kl
GBS2poNJptnTN6CnlC69bmIrTvnpbRM/VlSL9Qely5puRi9SrNEaFuRp/aA+
i1j5tYRgVatbuY4+8NCYp6aNhdqBzfXPkiel2fBrkoIHefR96eOoLrNeqC1V
V/WUTIWKWRQQC+tDucdyBD+pdrhUY0qwomLZGVLL6FRS9enxVPmYY4rSj7tV
xSwQgg6Kkqvyk+9e6zqip9VegB+4mZhbRnMy8R8m9Cg8zgMfoy9Vy53JY7Wn
6DucpnKXMcmyb5hEaJPZzvK4WX10l0x8ASqjzOnCFb7ZOi2Yzc6XKDuW9/hN
NajC16mmqTUE3MAEljehoYDezD9MaloWttkMKLGrfdF6bfOKfYuOpqkBohr+
zBr82PV+w3Vu/ORN9zNURrtpXn3Y4zWbkCXzcFNmFbP5q9hCYtFV3avieeBe
YJ67XKHFbriAlRxjDer4BWrGTt8GhB/4vF6kBteoZHtxmjgNnWFiQLjE4QI0
SPYBij8SYGthssj/vTNPsOrx8hY0Dkb8bbCI2vrha5H6oMeC+Gu9CrNy31HA
htxQMvx6Ay1uhrMVIXtT1UMURWbdS0qcNIToCZjml72naNEYzgQVGmjJrBXz
qplv4kVp0jG1qqRlKoQH91LNqCUQ75CU2fTYJjMQoVzqVF0H4InOYSgmnt4v
dbi2sTUYLvL0rVJHpa4qHFRjGrvEJFBHr6CHSvj4XF1QuvX0vCoyRbqDis9p
9cuQWyv4LyO430JaRGdJrbFyF2hkp/4RyYckP/98jpa+j9g1eq4spQ0eM3cT
Gpo2qzL2vYIvPtGXl6xmR132DOD6RF93IdacUmjoXFl6juarE6xjCwewDWvX
AJ2ZTv3y6QA7xDDzMvWFoQdMwhf3zp+H3+97s9wSWQZ+d88v3WTCiGkTrYvu
HHFO6rbcLJYC7KMIIvfj7vrNH6+Z3gSIS0PtEdCjIGxDAkdPMUt5jKiYRzJ6
/+vXOw3bB0zUlqHOwIq4TnG2AMgp1n/ZgPbcjD7WlK34lvKKO09XIWO9j3l6
ny1ju1VvhIwSn5iSgWldPKyOh/YwjX8PdQG+ij+yjngpdIMVerOJDhCQnwqv
cZiQh7UvXU0U7BijYvw1s++4MLo1uWVFnF0Jvn1Oe90pktvpxGtqfK+n4vOH
nMCT/CAaHZUH87qdD8ozNVtu2i4C2yH2fIcnf9Gahge2Z2IHb9KTTKGZaiW4
Z8+MrQPK3nDXMV1Pdx3OFj3tZyIsHr+jQO8UeOneibfuduR6VfwgzNHdOMN5
yaQ0I5vGZoe5uo1GhmkagK5vPxuNeoi5ACsyNVMG7n1lXPPoyhULlo1+8Nz5
ZqEpQhOF0ivuoTrTt2JCsomUNq9ASb/OpPCSl1iRFWAT/FMyAZXwTIiIZXPT
bdCNy2SJ48D4ZdGPShkJ0tPvoP8viNNrHyg/ocn8lpkT7CEBpcxTm4A+YbzM
61ZWhmkcx1L1YJSNjePgZrvmdO9OEsMngoDUiDD6HSKgGc3/ICyixiaTXp1I
Wq1eYLMEG1wWYUhN19OvtFCVTi6ytFTXOhj8dILwFWZ7nZhRce0GjrqVqTFm
p1WvVgEhefR1KLKA8u8bjtmDoMfIYcpptZSpQ0+0NAGS/2uagbGrJPeabh/Y
ENOpiXNiA07KjAEXLHaQZez59RzKf8kx308GMgX6AQm89LNrRl7uwdGG6+wL
/9Y1Aq4zYR1kUnkSHbw89s+GJRS0A3pg4NmNYK9D1/YYhIOA5h+9sDjUoIfy
BYfvelYRrcd5BU8ASIeau+AkYKOJqjwJJW33rKaMp4AyA1IqAJud9m5O9vnG
fqy15MbU8ZJ4OQEKfxA6potFVwwPMO4il1CLbo+i1fZic3Q1I9Sbjfvwljlb
/XktyW77ytTGQ/+7OgxYQ3SyrzJd8kP0dkIgDyeJOUczXK618ChdQBC1+zaH
I/xYccqMi5MDXq7plGeDKQebSW20QfzrSBZpq2t/Wla1iLULvI9giBXpjZQP
oiCLTMQgxkzNPgj+iq916DPb1IjHXnbplSbSlLgKIJZztLF8nRt2gYfMdoew
WhzamaqeCpCzT/MafkXCfPtc2xvgkSQ9BQW1WqnvUy12X1fVGhFPlKNFycMn
ZiTcm8mkb4jr2xd29S+NGHy/+bL0FyN9zLSUlN7uFUB+mMji1oe0VqjTXcsX
26Z7OpDSu4CJppGk4pXR80Rqx9W6PDNggdi06NCknOye+onm7c0Kuhd7APsq
9V9m4hzDbc4it3+vLVK84JrJ7wQKypSE3RgQGkFwnwOsYfxL/6dJDcv8V3wB
rl7SBigNqfHnyTNT1KyJsuZdGhLE1HJtcMSPy+8lXh6+HGoiLf0a9iFNHDKz
6bS43+V2sUjdfKUPlkiVG5s92kjuWA9j9t9V/WPtj6yrdL6M6GCT4Xqql/u0
vW3xIBcmBk9z9ajcc/I7uCZuuzdFw0FKVdShlsmsK6FfM5rAyZnVRNsnPp/v
L29sd1Grnq0CPwscOOr1tY2YT5pcuhlrySNfcqqKZJ7Tr3ymLlFEQPMD0Wzf
IDF+7WI9fnMW68BDC02EjYCMKvGFO1NB/HElLIkDC4ldHFKLUupeGpdUA42C
jFpXuZ3WCWqavmONxnIwpGXIA0gcKqjEDIPgnbLcP+SKG2yQytLeOkcXtf4q
Z8qbfJHI+w9huzIdDNDu3Kq+LnhI7xtAWfBcR2Ddq8JmLEFZmo6ubwf/7plp
0eFnRZY2p4zHRQk79LtMY3NHuIFLTam0aTyPdWtbli4ZgrEWny2YsYx3g214
nQUNi0YdP+yHLi4cdE4zYqS1+BHiNex8Aya+US3JeddTJYVYf/uQUgzh4fK6
K7A9ZeGsGwFlLPV6o9CvfWyVMlQ8EXAZfWgHB7yGiwpiS4VrVPSdQHEdhpb/
cCuusmBaAJrPPhVE5kuJVCoBxCAWuQwLcwXBtQXzxFU79IIocdGk9hh2dtqj
XwRpfUmxdubH1Tx4urpe22Fz713PaJCyZoN/tdjXVlp0i/qQtpe4UbHiJo9+
ykp/U31/a8WD227xI7tIHZINtLBGklCV2+pY9xa5Y4LTDqt4Ut///HGKQx0v
aXxtAPTimw6udQgBylSi+idAln2XdrVik3Xbvetjerrf4ffPggwt7wXQU0Bu
ixxsF8AfU9oDvUlPj/4jDrAX0ZaGQxFBAoDZUPO9UUAq+dwUdPrU4SAlheW7
Jk8CQ7R8PiCM0herEJVlPxjx+w1QBRT92hQIWHQuCqx+gof3GSfUAE3WO0x7
SJ0odbTiRjBDGRwBlELllLQnZsilyeWIbsWHob8vwBnQ3C1dk3Z/m4oc43rh
9u0YbPdTu/Jl9Y9IehNXQB+HonZ+mHl6fiel4MNj8tMO2LlYProkgdtLzQck
LDeo+ki8fPSg0d+y0ePwwt4TCvfDFqGkWPiG+7DXW5HtBTUXdR91IAVzd0I8
9tvUWiH3hyiz0DNIUqFjtJT01DqDyiO96+yjkFIwMnCiEw9U5z+2rQYoX6zg
OB0PbAvSGMafnGxmRftqRd5taRwNV6CcMMNFmSlExKujKa0HzWTvjyTABhJf
jq6q2C2JzcI3sztBTi6LmiJ1z6ByeUlLKYghaaMCZDKnLgzWh1wYZAegfB4y
NkvRcJoiFPq0/CmXrC6SQRs7SHeMzu5M0ubqNv/xokyeTkKrEtCJ/euZRzxd
JvJSweaaORR1ddek4+qFvpYb51ESkf/AQVHuOhyXUxKE4eOnzlTSXHr3Vc4F
S00SmmMxjTvTBG7Bp5jQI/txQvsu8ki/NEh6PQhl60EYYmKR9yg82SQH3uKM
cD9cLXDXwzgKa8JoN1gDXG0yjx8JZnrb/uJJKa3LYWlT/FQivx1zPE6agil7
FlrbFsr4y9dgVW4cJXLdJnNEORKQXfmEnnTN8WKBURsP2ip1E9Lu6ULEPisP
H6c8l6Y1EWpyp7j2kVpqilgL6gQMZDjUPsjcUyef3e2261pEtCLfSKCnZan4
SDAE6TZxaNEFyBfyqmbs2MpLvA/lKNMkBQzkZ10J2viDbO/yJwD9jkYZyAsW
riepIc/8xP95ibC0kK53zXzATqlmQvqdZKeZ9HrwaJ6cUJqmUgteEZzoyiml
uUto/Q8Knwk5m/LS9gmDDSvPMw5x5K7H+oUFJS0BfT9lI1Ki9DdiH32Sysjx
mk9Wn+G/Ozzxoxr6SgCgCkycI0ZoUeqbky2+1x2zBdYiOcp7ZW7ZbwjGl945
n0I8Ckyu+BKBTaEd3s+rngso/+VBjz5sY440BJ/nBKipBckNWGfXMKTXH3dX
nx57wdWsuNt8kIhMtXGsNybrEjaH4zP/SIh4JfSfHX0IWAN85gaZD+yJa7il
uy/chpLYUCwQ+iIuTRi8pJxHkZYdUlDZMcq3W5PJJCjf3gqUaQcfLXNDNgWn
HVZSXeL9T2JV+Z+pGMdbsV85fHMrIye/9I1fa1T+fOjuTxGVZBy0VdddwwWM
lsjeuu/qbVVpou4Ik2keunJ7SDzs27OF873R7b9Emqv/j4d7mdpAJZiHH4Pl
+C1LiyTyBaffcZEzuSE9zSo6mEjxMOCH1m2VaqRuFrphLfrEIKs+uYEhhQPv
VuVTed0c8HZBTD+V4ASDcHdeuZi6rFVC3wMY9KOe4TWzND5QM41mMGrOe+Hc
ll5+aYqp2sOCcYLmqCG+4yytkJtKjx8knrs/gWGicvBOJrfFUWBFsndEuPWG
oS5ksBXSEz6XgNvp8fuyjhXLxQYmUXX7bDe479C5EB+I2MuphZ4GBdT7TWzx
yBrcxWz9th9BkRnZH5gobRvjjJxUuO4RleFjOMkTcsOc2oAIWqZWK+E9r1L7
ToR/L5sdQQj0+10BM0RnjZfmCMcVhyNDnGAvRdjkEI8IpO6e/5O7SVVUqGoZ
7hpopzkwIFZDsbqMl+7EVvjYuCLgIpy+Kf+W2rYndWKhEA+V6bSBo4+VXTRr
M4zLbSkmY2QdT+XmwNKVFmWYGXoVsOvSrqERGD+9bKPdFJsdGNWQYFxo3WKX
IQxkBKH+74YkLecWV83A3LPjstoLuPPJT9mBljW+UBVz0ymnRn6LPRHEDV5y
gSU4srBKb63+2jlI15un8GX+oaHvN2DqaNJ16sv02+k6NsxzNnMUyKFEpLJr
H3I9gMYsNPp5JX30zoeesejTbInKUtAFsDJWYVmvELvchqgnrljYOcAA0XUw
oD53Tc6ySZLxEr86uHW/0IAbHN5JmPuUAYniq1z/9k4BCuLdq8YKV9puwVlC
jm8gk7qeRA6cH6/qyWoT6heeegpp6rvcMCuL0SpS7tDCkgNQEYH7wVtnLVkN
6q4evtAo95NGNkg2ZaKzD/SMvPvfE8WfdStfEnErHY45blz/gs3F7+myHu/x
s61ojoQG1nuLFecq3VC8dVgfrxtuzc/WAefkcULTSbReO3rMDv8DjiBIq0GX
MaQQSMJOGWHq1nxjwDkhoeo7svo0IRZh61i2LExvZaLEelbvmR5xbj+aKSrX
Z6BUCk/UG6TCie65mYZPWSI+TRqxoAZ6jWv//2Q/UrEZ0OeW/HGRwowM6rCe
ibIBfNH7Mg+py37B9PGwMxNcd4Po3r2/4sGIJS34QULu0qs1BML1Oaf3ztyG
csgWdUZfPclRI/Xtcm+2SlKHd6VX7iqobrHwWQ0Ey1gXur3tNsy5M1TvBzFa
F32Tca7Uip6f0/gstV0r4mGBUARVt3DU8xPAFQ+W82Zd3/snuY9TNyVxFBHY
BjURAIHtKZsOVziceujKfOabFSFea8EN0PCMUp1C3VeyttiBCe7o4yzmWwPp
5hLsUfEZTdFvZXEY4dy8z2o7aAH0l11i6s/Zi/moNz5PJdHw3W5DSdHp50+L
bMjhaVYsYG/rzrtl3Bcr7E1j4WRkMhlOVGlAmWTjDyy8RaFUWLiaSK9Chs4i
YSpHIi6ydIgoNfN2FgDQls7Y/1Odi0Kb8RKEfngxXZFi1Qk4aA5N2oT5hucP
r5evBqpXCzONphb6C9KkZJOh7u7x8BA1Va31FTQQ6iAYUAiTAEbT87C1TDXT
AfrvU6bBMD55KNdZ6qyY+5KMil6/uUC/pQ==

`pragma protect end_protected
