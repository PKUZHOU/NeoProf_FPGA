// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
bgF/hK4mkUkpWtsh+Fl2qPgOjlEJjFJb9GOX/86NZX20HwIKiSF4be6RHjthKHVH
hpkcvPttEZVk+h+jRJpS4xgJM/CEqYxkQRvws8kx6g3Tq6bInuT8/udHbL06i5eg
QyxORJP78RWhOW0BeVBDIRpZgESv/lWzHB5Sd8BaICg=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 9616 )
`pragma protect data_block
6szYmECcdUEqKHiBL8y+zleu+cdE+cfaZ0ONKhjvgb0DcqHDCU3uJIv5X6Hy3gZg
Lw0SvT+jMd9CtiufzAfmsBiENw8iQyhu/N1jYoE4Hhk0AG/ajDhREM4YRSZeNNxX
Zt4MKrLW+7JqqesV7pwYbrM3Y3tYtGs3hdSZEPfYEEm3kTb+UnacdZCcakxMwqne
5KtSSgktwDhOgLkvLKQa7xlv99ChLlcfzAXFvazmgWYtpzmHo0NfXaPDOtzZTw61
bIEHOZJ8v0TZREtv1YYlxAmYPo2rB9ljeSyIQif20W+zmrBrMcHmh+7OGOtpnBFZ
zysEjnNQ/IoEqeyQvAvmLCcxKYqdc/H5m6H4Dwlr2WODKbNFGcAmSYDOWFRf19rn
ra0vAJEOgYl2+DcZMGuvGsKZ4kVVC1WSMMwHMOxzD2Mi2UwgzPGtS9n4aAlypIo6
0eItZdu86t1iDJOMu80+IZh2jaUMpFNpciANAjHSdBwYOTKLMp1rDg5da9rUjg5T
Uph8PEJIfe6DqQwBYeRdAsBWBRA+7GGMoG4qI1GuhYbhzU7IWbjBup2FPmLdtHoO
ooAtfT3l41nf5PDMVYyHxr464BhRDeTM+Zv4vlQZ7R5LaCzRT1lWZI73ORhLKSEv
IespE25fseTfmkOogXd6YZrfZmeHU0GpkFnua/F119cGYZulAKyceL96p9K86AnI
VB2Zu5rMAbS752IkSqq9PPUCliowLg8XGKm+mnPCmQOPdw3WPUWHDKbEEEZ/8Z5v
nNqpxzgUd/Nky9r1nr6rA3xmswh+gk+kp5vRGZp3o9zvp5a+gUUvIbRBTrUOcR6F
4KOLeV0AL/7KvzOLuRpV0OV7krvJ5QAxt89kXZqr8MIWMqxNP5u9NNmcYQzU61vN
j8ezvjTAQixaWA2AA+AQC5ZZTwUecBOX/OVo+Uu7GvUEFJiQztlhlOr1cNCLMpiJ
AaeEc7SdzmiFtSSeNJSi1T3T8ODr8880h3zpwz2eL3P/+j1TXHL0qPUxLqVZHnQU
d7m6fHoogve4dx/jioFdarRfCWLXzZRAx+S0ma3kqe1zRybIozEEGxDKC/czx2Ls
+RnafegsshNoyCSZkdhdSDhSN1JG53xQ5ai+46KQv2q9JqGIU5oz3enLs1OPYx5N
mji/5BMOu3BdW6siCbSWxxQjKlq0jtmrEFWx7wFQfgLIV2mW2rQ9l04OJdtdzdZu
SPCgdxs0yZ0Bfb+ay+qu6icQ7I5yzFuZffEWfKYkvPuEfQL52oSxkmuUE5NDYW77
AKSqHxOfT0WizM412MndwtZkppALa8RKmm3X8qpPcl6qus0aPAcTtTp0Guatt6l5
izltp7IB466gY+mEFmlx5oOf6kvQE54ruFQ3BjsiCI4zeLPptB9gswjhqLOhhY7j
FMbzICXtGFNgv6GJ7pwvDfCpti6c3N9047oBDW/PNoiua/C6yi+flYgkCSpp8rfB
KK1Pt0ojDJm5CR0q+cMNGzdJJW2PdCVAEq4ez7Z7DmOvXE7snQMkr/j+lri1qO7S
gMoFhTtGC6h0DY3YGMDn1ckDbFbQqHarhAPw4wXkCcRddNh6TGvvX07IB1o6c1xc
iF62v7yy/KJffAAKducVtfC4eT1eFYFgKfQE2LEY1WEsC1lyFjkQmPMcvfjKZVfA
1FcojkkTh1n26k/pNMvBU4tNrIuNQ8zBXdb4ScIfg+ScFlxS9Er5RWfyRPBuJe95
74a5rHs5czHn3Q8RYPu9CDHVRKSXNP4dpdxwXk5TV1EhdvqDwef2qaa91To9FVWZ
YB4QKrd7Ap8u4ofApLiXI5iq+F/YmABVYwH8hKnYpujX1DKo/5Mu/lSz8kQd+jHr
5nrS4d6Ua2diFVNLchgFGfjsoW4pTte1lm9P0XgVkF3loBNLDGf2LuG6JIixj/hY
20m6rZOjBpc1/IfU5mwBiQyoU79IubDyZxNUfvU8l2tluRjAzxwb1gmdnCjwPiYJ
VFSusTi3KItXrxkwDhnKDIkKTGMdxb0BbXSjbSJ4ddqrcpcb9wWTkHsc5U/CeEdC
4RTp0smvGw6sJqprmyKlkukr2ak50Gw14fnIgM/ntrNt84FzcD/BXaeIZVk6+jWm
iWgq2kA0RCiqMj3pRTIJDXIScSvhrSo6jZKHYrBTwnocMpDf/9gd/s8C3CF+2Z3s
DTjuA+ZQTMFaSoGzWVh7b5Y/o4WMvLxj3TWbOBRS3qKH0al1Tu+QrzMXZNKkCr8l
+bU6Ah3swKMZddmMhcAPiPqbNjFL2QLjs7R5BQyVk2tFgbEhUVBdvrztbg0Fujs/
xP/tEin+PknB9a9bYY1OyNx4lIoJZ/hIsUz6la2EsbYn6fKwkejnNU1rAi2xeS8B
p7X0AI8xB0cB/tdOUmsMahhTIt2wq7Yz8M/qtqgv1O6+gu6lNzNkTmJ41KUihOZc
zJugiUUyHLEYlyGV4fyKOw9gouCV/Yx8qhlUhEL6Gm9qnsvrcYMeYd1gPk9QACK2
iE3mxp9FFRTPECXX6g1d8S9RYlv1xHHa1Z7iPd6kG0iSomsnG51TzzIPug4MW4d2
n5f4c4Yq97Ww68KJ11YXfQlIjkVFvPSmDhASG585+F6uIOk6l5nlF/pO4GRxdJED
tp/rd3OzeCvw6+5UB9E/sFp+O9wRW8gPHYLQGfwfy3nq9wJifGRFDVQn6BwdbyAp
CapICWLEMMBLNDm766nVSsWcbSMqXG2SK/JwMZjYMH6j1IRfmZH9cI6RPJciqLh6
+DglbNGGhLgl5KG8q/cVvXAgFZouVdk4sg1Uo3Y74SQmPeF9seKNw2OzSZ43uzdy
HQEGMEljF02EClMhxhqrilUeC08t3J7P0gYxCdklW2rIyzok+0W4oH54Q2qBcGW7
I9FPfk68/EQseQ4+NabghDe6ppHns1a91IdR3mBI88bW5ztt2lzayI5Fk91mTPU5
SG0CW45nnRmkKDjffdhPzdZ4e1arZMuZ2mgXbj+DQcqPz1q/lqsweebzlDag+h5p
n321e2BWN8boBN8vkOgyGhSJjBEvg+FXxiCmbXEytRtLRiX394ZlR50VYdI/xONp
O9W15kqTzjjGP/CDGK/HU370cHNr2EkiI2J/i+mkz4PJF3Z+k7W7jrCe11cKyF3a
MDJttYA5QkXBiy+fVcTYZ2SixeL3BoKazwsFR74sshmcX/tJZELdlm/kVeXg9vCs
nnMRmdaRKT8DHmP6CFD+hvxhhzaQPe6PIS8I5r8tjNtMII+TDOhE7a8ixNKj0mII
Smnycs6SR0fiPVp/LbASJO2m9Lv8hrAOzsgh6RWyt7riw/3Xs2PWYr9r9g1Tn2nK
o5TdJ05edQeUnXUJPfMDXXhiOSRPoR644jPXCUzEc9BngeXfw4YzO8kn0xHiDJuV
mnuxE/iEYTioMebLeKPlPJM4XCvTxeuqyd0KmRbW011xM+aJyt3+VbjRgUZayCs8
Wsfm+z660vqxOB3MMkw+Uf8Qr2uUSUkrMsuKtyvI+ki/wiSaXoJ043zyjM7iep08
y/YuROyjuiD+hE0w54nDWUur5GHyuEnM/w+O8gRkTKHd5jDymlmupyjroJ1Qw0SA
Drm93RC07dttvD6JwNdqZRf8LZBFR10nUEnsFPpNkDgIq6kLgDOyr/H/OjsQczHI
hiyp1yZXSP/JrpxU+3WVDscDXoet8o0SQqX1x1bPrGK5y93QoU97Ea4tIHx4I+Ng
H2FrtyCoY2RvJ9N/870ZcX67uHgYu4Ha7UgEPJx/6AV/7xR/9W5WQKpPjEF0O85C
SmYzUnHG75ycF4LwjzZbQZetd2osrXhSiLl7e1hqGqVbU96FEAX7sX3y1C4eyNOs
PG+HEXRsk+kCvVqXhYjr5MSvdGRSxiK4F8FKaZi5hbKYR9hMGJlEZtktyiuzGNY4
Rq0wOYG1XHKVV49WVBU6yyyZ0o+QX0maBbfQYhS9Gmb4IZjrylFjVpM8AlgRvY4A
H0VrF2AtvPTEzt8yLG0Y8YOkz+c0wW6ZZVI68xHk/4VU8tKJ7koDITBZevbgbFNk
B0OqHFFLGndoB+kqDifqW56qo0QA5wVw97ul7lElIxbViwrt9+1E+eyQJBfMqZlM
VaQ5VZF/mVOerRZdne/GAwaSaQH97gZSn1VotDuq7A/I1dAaAekx188vM/YbR8yX
JAvi4CjnBcEmSPYnNCTdYMMef8QDa6o/IXYG//aFJB0WZj3oT6pOj5NeZIevL625
aS3U3ECjFrCjKZzzL4vHcaBw0jN9Gd8idTk/TxODoSYEmGmFkrGVLFXi/gpSuuR6
ZYEKEP9xFZ0n52fb9lLNKH59np5carGLUYF+pYG2/KSNXeN0T0roQEpHHC72g6tx
08GeJqgr2MZklKaSQCkrzhGpqnG2wFfdx4C8+zj1S0FRj1IRPpLFoZ5BoUxNsIYI
XY2Q9dcbFwIWgfzxUlDLWWR+xMgihsjj1HlmAMj1m/FP1iwu8l93W9PjWKgCZbLq
ht+mt0eGzZyTti35x9gld4rcivTiKyL1ZS6j9Obhynrqef5qNBGhQZyJVbK8fHbv
zaMusngo+omXwXsUi6HtkwakUKTofRd+W06F/lhnRD6DAw5KCY6U3moKkJehRVc3
HgOIGDAwcTxMrbLXSNfVpl1TdUlP/hxBSxgiA0FXdHI2HVwYWYL1kEYIhMfDWVCY
GXfX8pFsZntcZ+YMlXMa3U4JYn8PwXh97Rxa5wbHnHOia9imJ6sTjsmsPiWdTW9u
8TzZLFgtqhflCHXpj0yKc1aBuE4ZhKtgHLZNxyQrFczoyv2hFrDYXm+HNwXXTB7S
SjtUGLFVjsbLboVNXhjpb0pb3G3ZCCashCva/o6DYacaDtPxF4PtcQ1Yjw+qt7/L
n4V8GJrqbrUEsWEyywq0oB/dTlxr/m3zO+bpfe0vKQEO0/0P5gteSz/Gg8t+dQv2
A/Xkxo7F8YUXknnRzW11fs0bWlcaQK7duLw3VmHXq8ppjg+eIizY0iNK6C+vPbjT
HUGKndFHGJT0KBDXu6o4KDvsAqG4fVZ1e1gjV6mSiP7773nfDaz8tKG7j20zlI4J
8iC7DfKFKW4IQMnjx+ADrkIlzRTb7Hw35dXFiVM55Ar3rHUkE8hdIY5tIv/hJ6aw
cKnaibKuEPsM4QjXEEaelJHUuQHhwoDEWMNCeQHugJJx9/BecpRIbRGtXv8EoNhQ
eznurEPRXtnZGlWgIi2mNuWZpz5BN1ooo2eEdxOQ+flyJcGv5Kjc9LJjTdzQABto
hzqwe9nhzzake54Cfto3aYp/qG5/Db5lQEL9Hrec9X8I7CovfTL9Eq+5eLbpQ/5X
/D7OnV/HapIokk6FGfspVzF7/A+8lEd+Grlj1vQrV6nAL5zpm9SC0POf4kx/Kj1/
q4QXQOg10SrxH6HmjXkT8x9dnYj4ktxMZXiTsowEIT285gyAUADplM5Zd83e1Uz5
EKRfm6igsu5cPIxeecTTg7PdXsAhsgN7oP8NtGk+UdByQ9NrqaoBlLLhKYrQx6ZH
kRNwfI7MvQAQUy7Sz32GeN6QOlO3BDOJuCJTy/65J5PjKi8az3Q+ExGoObdPmVCg
SwsV6gdtGBmzj1zdr7hhGkwIRYK+ibATjqJK0nFl2hwOqVYsC1xQ1Ad9J9NAYUPK
K24whQb/h0oA/PLfNdNY429vDp25F+O7eNlVAnXAllyojcVO89vHvdgryJ0FWhVE
rs5Y9UFaJVd8gkBJC5UnoTpWNJZncm51nEhiMF4ZhkxXFilNHN0XUAblfhLJczWH
cZtLFPvMmfa9H3+/AmfbiI/3kgg51v9FtgUgtJUNknwO9cXukUklLsRgxvB09J8K
CT20uY5J2JQhiYrCGiKfXUKbAOvEwDXZ9HMCu8ME3s0ifabHqNonNfivFXh3+oke
wytaWrarAshbrJM5QiuBRAiApw/3vYhkadotdHfbQaWimt4r8g7PRRJFPoR0GV0g
H1wd2YfNd+rJnJOI+zlkMEjjEm1nGQ8nqbD5xGDE3Q2hZeswTa7JqHcCNMVprm7M
g10BH04lP9FuJsP8nhEc8ctg2+j/kx60oJ+b5mCcA7NRELbL9BxVRxyiU5g++60U
l7FZlLap7LQAV1Y37XVaOFGKwvJrhhQ6DMDHZWTIXqC9SA6isw+vErDEE+Hb0hZi
pkZH9vcv7WJ3hiom1Lmd1a+H53CGTqeXpBGxmp+vBHtfeybkMmcFxdZ4N2I5NVzm
85zW4dHddokLDMsZ9t7hHVECpLccsw0TknE2NSzk7BDZ9nH/9ZQM2JgXfP3cNDTg
rpjw8yVpN7BKJHZQC77Ha0r4S9b3/RBPq2RLyqXZkfwQCqdNUB9vnKkLhmKJX4wk
mNl27Jk0wX5nmrLn+pYwAfk9HKCOWZEbrNABcRRcUTCxzTb72uDU3Rz5hwUYjCmj
2pSJkdFsvAmA8zV2JhReJiVvxSN6ETYYkKi0FGLNTBPjvf7dctiQr6pka3QyiUwx
L/chqfAkK3d0JZCLLfyI8k40kG6+xQYVPdd72WFr7f8QBRosmFJqpQbncv5R7J+S
384lMJkRlKy1XExmTnCU2wwT18Pizmrz/iBQQIZTYvVE96kO3Mc8SBief1GKM/+s
jq8b6NHCHORFpxrcKH7HVvpgCyxaTmPEsyuNQR/vQP2EJNPRpYOSqJtzMLCFLtws
4b3zVV/2jDVDXNBHseecrA0L5Ez0qu9X3T3AWBkAK4+uEW0R4yjbKvGXgbWMoVNe
Q4PsDDTwKXB0O5STLxqmS1SsIVr+veeEoo7rW9g2zvkfWRsnAdmJ9OSx95ApyWaw
zReQ9ABvPB1xihYvdiA9aPTrjOn/7MsrNlcdG6nfqZVrdmRkgVCD4vZ1UsyKuRAM
7F2xPShTWUtd4Mw7CFNZAZxrUkyfJ3S0I06wRu1sk5rzB+yNi0ZF623Gs8AkxUsa
sy9xkWPKUiFCv1PvLuFaA/VJSGu05NZ7VSSw3m13BcCxW7bfTyrXTW16Ri202Kys
kuGyOCPeGZJy6dLnepwzPFAjXdwOHXrnq+mwMW3HnClhS7vsTvqn+EKDNcEEoulH
89rhDg3AWW7YCQPdbqF0KsrvPqRKGibVAHBpqV9kuQ25rUK15LbHpd320Y0kVeID
rEERcWcRMWZBjc1cHU4YCIlbIh1lJYM7gWKg92eI+AsfF2lKWa7WZ314Jc7PhilR
XqEzmxxrFy4IaU3bOG9idBKZhhNpApdDxa+UU2ztQr7eGdhpyXf9QcQrdvTh4KQO
s2R6XbvbzngDX3IkKqwqmKsrry3m6I5OOkUDIiQV1bBQBuM4RxXWKPGUo9hQkn3i
+q8a0p+hq3GOD8py04ipELUUPssCGP0X5z7GAab/WgFffvKr0QNJyUpmknCdtpPv
9rKLfavG0E+XCTO6ZeQhU1493/gCHQPS1Z+hcU5kAoeGvfHuNzMJMp3U8WnH8OTo
rqpaZCN7csg886cMKcJvaWNSVXK55qhcsFvG86TYXUON61Xq3MfV6RSusJ1eTb/q
+aqdyfN5Nzksu6iC+62B/EdHEPdwsBuvLUoL4OXPBVi7E/XZpQYDXtBdmibxlZjZ
i0SEKVnZigKc4nrdELYJqnaj0Te3goywVEvVfgwxO6aQxpoT7K+dTdTqSdkBEkuv
aRYvLyejml19TYxEjWwlx8YBXy3eyBnSDa9qxEwrqDtWnugEw4EgiLxt6I+8E/+x
VZqHVGGtQH6rHpn/PC8+KvfDI3Klfg5MFIhac0fr9xwkZ8EwhjABo82aMRsXNJyS
hBw0ADa8FBoDBJi9Gp+JeD4OiC3U/22XxsMkqzl3JyoSZZNhJHd11PGUfpapQmzw
JvFNBjRzGEjWEedwy9+f17DI+W95NQHYYZnipRf46dNVfI16sP1ElFAFqbzCiNvf
rKZJGA4da0Zwvoo8vP8T8f7AEkv5YTTdqHPgiiYQZT1k3N/+0udVTyStMfHpahed
+wTzOROTrIQsr39xTdw3d+1ciCk83MQ21ByVIpAZj0+RhRAeQm4v1pcGVmo59qBm
VclKGY1ovNEfC4ChddeDQhGxhzD63FcSrFKB8vwPN+mJkV0M2eofEx6kONpVPs8P
HBfmTlBy46MQBDpQMhwvt5fFPZISbSFSso3efi1f+N1Z6pGObKoL0ly1NGTkdZst
edjqamEkyxzgZ1sfMOqSaSPr1swJ2kHiFR1OdCTRO93OaNkyFQrMvtYAQDX6lHSm
lGXuwx0HZt7ylJ9LAuZQ1ousw9E0vPrXzMmdjg4+ag1IMdptzxtnUw03beStjPFK
0BSNPu3siw7jpYe4rTE+V8/CbuPhBcKhf4w/+qHEYwh8h3EACad3Ad6YAVKWGgcB
y482Hy1RSf4Q9D/sYeuQR0/uAB2nW1q+xz6aNZgo7Azkzc1yTCFk6a4l5B6sbsj1
9TDtUpX1Rf3xRTLXD6Id+jcLe2I8gUhXdoWURlTd9iw2OXGcy8hbXLhFKH18iLsE
AAK4lF01Qfm0wsKA49KiSpgNOCl79NGVsN0Lmh8hgero5oyfm2YFmYUp9XyNJUGs
HRnd1PiUZO4HUtyUhDckaimae+ldazocPKrOQvflR+TzC8TqtBZ71CVMWYzVEzjF
OQgPMJSvmAx+Eg+M4N4EIuVAB2hypxAF6T/0WjCc7bsTNXy3RVPeIJlMZfGsgdLf
N7YqgSZEsFKfxwpnBnWaoqwuF6X/I19Tf7+dhmb8kj9tZRpSrbzA0E0epIFdvWOd
/BawHqwHSPyibehrySy5B9xN6vJ6d+S1nXQEfVRQ+LJUjXF27lMjXeKOEAYjHYvL
O3WVtL+AS4+ej3FEHe0SZbw0Zg+trmuDOAmay5GwH7fnF9MUC6+tSFWLbdaGdFBD
bNgSVk+T7eWvMxV8yIlXrcdPbvtuKcuHF7MummgJHuPwqxCAJOd0rYYpv3lSAPiU
4HKtkGgNxpkAZveq1p4Gzzw7hWojT0MqDqapQd/EvOQiRLOaUAUpwQLJarXq+iT+
xNN5qo46S9r9Pr0nwkoYE59ENi+Gf5pNl2cBJ4U7UWFI92anv8UmN4jXKjiltK0u
9qacjwgRyUqXbmA+nQdeWdO5GsGPLTIRbhOwQx6O8bR1qd/WRrIFcXMAXUpq8Ytd
LDCO+jX5wCfw610QDizMCB1Fowj08KM2AVYnt6uzZv136mxgBCz00xXBA/mi8gWL
O9qhDTOO2dwKZXlprk8eK0FJWhggegs3huMosXs7hjaXcszfphMqoEZY6IJ5x0BI
qCnBkafQULyAIhh3mczvIEVLUUHqeZM031XIBDfDtEfvs6e+blfreubCAw12AvXM
dQ94p9nCxQmXBOpzOn8Bthsdewb9s7gu7tbpUFHbGNoQlcwnQZKbDkzOAOgyrQp7
rTO+7Wri1OyI+5DOPOjIRJ7rMOrs4N/Mv424JuhF33YcJ1POWViXJboi7SC4AkoV
g4bLrh7w595FLQN83Nki+J89KhcBHBeE9HT4bKSJeeN8l174wSp45eFg31fhQOMJ
KWsOE4HU/t43luALMv7C7OR+35AkBQDL3lOXcMDx7OSdo7m8P7GZtxQCaYVqweLk
NupK8fUmI8sTQo7hEht3N5p3VO90Jj3wkMr3uGEsNHKr1HJu/5rxHz9bultD8mbP
7QmYhFYJ9QZOdWaGii6JJmL8GQq9bLnx/mmURTt6Kc5t/K+jQZJTMAqjEm2VRNLF
JOXuO5NPEI24ntA/Wct3MgYQlPAAtOFUax6A5bbFvMyHtarb0p0n9mr9j5w8FECc
s8Ru+/1XB34jJpzDDI9qvk2Ejc+0f3Ocg0dGpJ2/tSrm3HajPFCLC5msdCsB0j/g
lisdW7x1BKj1Pq1XQ+Qr76w9SaJIh5IKEx9lvRNEXNsoJk0s7ABvFZZTl5b6A4k3
anEiACUVq4eY/3Fmf15nxxGWQuVYR/vOmiTuC6pWW9UwRgwV29lCUmwb0ocpOTVR
OvM5Ls61HbjELClVQMpETgtByU4YrtJRjO+EIrsZ4HOC5YXzMH4CpUchDgQEYLhN
g1FnCnjrEyOldNUhzipO7Jt1KzqkbyOw9ylnfLqhgfb9b+QqY7TaT7SSZHy/U8fU
WMDfdGHyQnCixDDP1GjMVp4KdU6BqlLi/iVyYmIYuO/PdaY8Gt6GX1VpWpGzAALT
j8iweVj3iRN3EtGFXzd1HcishkawX8oPD4z4Ej6M/+GxmeyuSAgFNLA5CviygzyQ
LDLSbhO3ofEV5CqT2/bgYSC5S8rBmVBHq+sVkRB6jTPwx2hsYmYn5qY+tqMYNSTI
ykn2d2D8O1u9Xk2H5P0SBeLBcZYdSLd5mTT3rYrP2MA51186tNs7NHQg/RRt+jDI
xI05zAPYycjAXuCgVhpx2fUke11c8DWAQ/yLh2UXKdkPn9adtl98VRF2jRmiSGB8
9VG2rmPyHVZo96CwRgmmqQkvmqq9L54IYdy6ZuS1hiV6jzAwqsR/6wqylBVrz84s
2ThAeV66/n6ul1ZMFd5BMiHJ2d4jxhFwms1mXVUfPT1UeUKrIlMG6cNEBqJh6mtc
BbSv/Om84o/8mB/yEpepKUoE/A6uGeyunLCJ1N3U2VGXlijgu9e9ycqPZUaXwJbU
BwcxA4nAUpd6AV99LUHGfeS6KFWxRKK4pQT7Gwjd2lrs/NEcvBcaUcKtO+74dHvA
4YmuuvOk43k1QoyzIzoob0r6PBgY9F/s0KC9iKFDChBiIz4rBShLA6Roz+pNo2hW
DUQYWF7aq2n4OG6E6bt+9MayAwBGd8ROIAfLMoPQC1TTCaB3QSrRuw3SZLbLqCMu
KsEpmR/x4HGgY61r6DPfdO2ING9GjsCfUgOeQ481Oon+yv7fnp0AloQjxbKlWbkg
x36FbFQv8T167o+Bvp0dG13MG0DeSKnPL9Et9yPGnEbXwQil5XcK9eM+vHYYh9mU
2t1d4HLfEqyN92qGYsBmPZHLH7/D+35K/TraDxnz8LjrwbwIIHscP/WaA6tWBZ8b
j/QejCDDFUp8hH0xI0La16fzeeyZqxSDn6ASgTHDfHVFgbLytQYupLapzGQfwrVY
ozshhPeMZ7SAiYoKwmhtlRe2jnnjVLZa5hKb31iN7Gr7ApC5TvRl1sKQYiILb5cs
ViuQmyTTl3QrYD+pNhOeGSYS84FMEah8F1e7TXGuTLyfiAlCM4CYsvikPknVqbqA
4yEk6FsfPTR8JwVMoKEDHYDVk5HXfFaM3+dy3opoqMBAklW2DhGtoDNjot4r8DRB
I1SMIdeLMkBDHSF1+Riw5pka0Kac/IpUfkHfIYaKkEMw5EwsCCkVZcezUmZIiL19
AKMfbhKqCnrjcUdMuWlzKuxiUUTkmE7ZiE+Eis29j1bvQh0Bf6rMiyzKqksf+aTm
Fsd8yP++w1whOflD6bKRMhSC7oCr8Kis3BhXvClVfMjwovkTWRrr0hCuKpSr/Gm5
/4GJYgN2135JB9LF/lgXT2ep3p4+wcYvew4P3jx0Fytua6znOYntcdfhvByN7ZOt
e0YFdyih86WZ2wcImARNjWl5548sqpWJw99NdCyKN1g4VdtT4OHEU5aaveG/uIl0
8b4W03zEg19BPopilXXrUpl4iWDDGOJ0+/zfKEDdg5Z16ymbki45+sxmYf8vgetH
p491gzD4tH7kbZN7XAtqVnxPAEtJU8KCk7Vm73aIRY/e3/ket8DbxRLCU+tnlz2K
eMtfyghtoanlTBlbm5b2ukBGkLCbgv4TlV0q4OSgEE70LLNYIG+z1ex7AqhINwV7
maFueiNgxbqdDwPUtcSXmAlXqxRSuKdfNxjXwxk8lrXlLbrB7lSxfTxZJruLBt7z
ib4XbZWa13aNibpYczl0BbwqWSTaBeW9wPmqDP5KDjqzaeQPeYN0+GOUmwK9SyYs
HdYoG0obh/wsTyeMe0a1Q3C9Ar4S9wrkRfc1iR0kZFObCkJbyAlGalbd/txUklFm
dchgEB40cEUF2WJPvDDg8TvcHeVwXuqx5Sis+s+xutI+v0sO9hO+HzGBAYsECXom
TFyjmBhAjVwRaQQrGIqHoLtpWaHK8mjNZ+ZckFlgaq9A1H0Ht2tKoKaNgN39mh0w
IRCBJMi/xcu3HUlMvdTH3cJbujzPSPouEb69bRKdUpxLdJnq217oTgJobFb9VGLY
EtYM9YV3ZFrC/tFHZswgzWGzGkVJXqtaRAcbqXXtpmVN8MNyHZrLzV4BSb4uCOrG
omzx9vebUzao7rccUR7+sPvfy9v4BLKQ5VjI/PFw4eCNTmPouUJpqBWHEw2fW1B4
ceX0jAvFoOAt4Srr9aD42fLIU9ey9njGOznfwxdEbg10+F8mAmyJw8Xh3MmqHTh7
sjeFS/fqEFwlaeXH6IORABIEVgk1dmwvPvqyoBCFdoxsmZc51uiS1pqcVgdAJmp9
JXtAjLx9qfQ08GimTN+ljguHPkgL4CE8ehmiYM6BQsN8vOQ9f6ZlVCWknKhR8SXW
yjJtZwICw/SkNSSRRaJglTMd64RZxCPfv6d26zyXYUTsoLMFrCOFdFt1xIVT7TzU
vQuhHPGYRDNvX8vUtJWjh+RjbflOSgXrw5qHB2HZ9UudHyeVdcvl0n3lnSMQJiSR
qNns4u0BqqDGQJr4o09JmZAMADrhF9J5RRBV65jLZfcHDO85k2rFPgkiQ/agYGP+
WJwjA9PUZ9IPyweWtU5UHmrgxcqREoAkk/CCEx3MKJgxrKQAUS0V3QUn4wwgOZoP
Q1V5kjXURvT1uOra/ISlRiu6eBUNB0Q1x/O30iy7k6wlS5HXBq4tdYwKZER02m4P
xCPY1tMfksrbkO4UV6lLfjD67Sb/vcbMuKo3PNAaM5JBWJtT4z64D3RyJ750X1X6
XyqTbD5X6XUTkQekNqmvzg==

`pragma protect end_protected
