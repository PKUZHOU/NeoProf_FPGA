// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
LXkwmD9cDvSv3YTQAsgJ3WYYLRGKBVMd1+v5YAb35Z26XmbBsW/OdeNzr+Tq
EJn0rcExpUfD1EAo39W+zULbfM6LjvEAXspwlyztvIeVRFPtOv+P/b/WqG2M
o0kvowurLWdNeyapg3Iv6NY6aLn7ZuAi/2x1pjvgxJvpNecBquUkvll0A8ov
h6yLvCERZRp1Mee3rnhH3wKzA4ZFBwTSzY8WodpljXGaE5y3HzKnaViJ3DKo
2wtUUYoL3JN08DIBhwBhUwYKZ13zMdToaaldZaqn8d+70vK8YoeyJJSb1Wsk
0xsED0WgXW8zOEunq4auHr/pK9xiFH4J8hRdhwYE8A==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Sa9Slcdfm6R79RQI36HoS336qf5hsYW7zfPhHDaLn06QabU0wMU0iKJRRpPl
DJ/MbuxsjCEwIJsWc/rP9xLD9Mx1gBG3q0km+mj/PE7bJPPoC+a6c6hYoLhV
72mWagqjkyBxI3OHbtBSwVivCtULN1ROvpUZHPXKvyeq30olJ+6psmjHIOBJ
3Yvel0E49k29/S6/sJqxu7de7vlwhY4f1AK7dX6gD3mor7kmHb2V3uD3JWYn
P4tTZmOHyUrfydoKzzhpGqMTeIa+akeQK7zl5rr29Ac6NpllYP6UWWfefVns
vcwP2POP9PkvpXA5HRAndCFDEWBe6hUrgygpwPHyIA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZvPIudORU1VHevPYL7OFTRBnGJiy0PBkXNe9ogFN0bBD/YqvhkVWWKlmreH+
D9mVZ1ugyRfsD+t7Twq8OChpmLZywHQGXFfI0gAk42Jo76BC3vF+8/0i6wCg
Tlh4Z3kjNMMn0bVFCqXAak/SR/NqsSbEQbvj2VOTlQjDonY8w0lffDc0PK2V
t/IUoGHGEGoWDf3hg2rGVnmaXF3TozT7JXOEWW2SOcqhIXJkJJZXIgh19EbX
pHyFbjVa4GqAaDRBL/mO1z3X1KfiCL1L3CH88HfFO20wvmrSX2LgbvM99cjR
6dUA3qTL+7T+09k0vHfhnulDE3IFq1veld+zU+nYvw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
RGj3PdGRlP0l8UNOWkJfR2+VndjWB/ddforAVsMwzna9SjRNLy00wik7xZXK
BrmwwYMLBzbFdtpnNXlDWkMaMobeFlwD3rkgE25MlEnWIozFqZKE6j3jKowS
usN5JEGFcGDzmkBWHtvUsnK9MVrLVbDBUzZHx72E2QmPuz6OsfU=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
PIOXzmItjzDGUoykQKf1bUSo2mpCzuEoWnSQD9RKFtwSMYl5de856CBuKHX/
Yb+D1zOtW3v7bO473PSilFbpYg5gfOYWqqVsAPKrAJ4ewfbGxVKAPgC2UWaO
ciX4EtIurmthcIdolmDJJ7bQYPCgmsj99LxSPED6U+tXw/jR0JvnrtTvjgGl
lZHkU1YMDf4VYkV3gvAYMl79NZiQfL/glop0F0EiYvwYbHtuAf9z3CyOXP6J
UCF3U2if/923hROiY9UQNDmvnO2a/6AT19jvWpbQPAYMz6uIxh0XAu6vN7Sv
7COxR8gz+3aGs9igKoATullFoViyDQnHwrK4mSeAN4b48N7LnqaXMJX+fWKX
VilZJh0vJIIMufsyCyqopj1NscE9s7PSGN2W054vbMI+LI9d9q1H4kKcg1uG
8B4RC67TTBZ1+LkkdHvpA6Wjq4cyfQW4LoyJGRxFI8Fe1fRoE8MkTJenlnkc
32JpX0LL9Znn2qa0jqPDpBkwT5TANtA/


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
C8R5CdlU5qxu7yyz+HjY50VAEzWnpNBDNykoHKNQoQXpS11RzEoVmJTsVsmH
OAZrY/3y/71UbuOzq+myaiToM4oDnQZUbanYiCfrpTnOJ+cRaF4nLWisb1Bj
ykb5Nzd3XAW7Xg74D7xilTFAOdmSR/f/DrEsym/BGICoO/GvRiM=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qq193zOmzZHHjQ3HLWw7ny1vHYTw7pBSWJgyd3k2Gt6Cy73LxnzYQ8cg6tgD
2cQKZXDM/lUeT5NkccnuX4dFpoqQsTNn61FcFZhiWrWVBRoQPr9SYT50vshd
znAS1aL5t3nF8C949gjoJAwlq3YDJllBGahaTRa2kfHUa72e4UQ=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8944)
`pragma protect data_block
xeyrKdr1nPmhv8k5jjz9sTZOcwrhVh4e9MEpecdNi/bjEos9Tplwp8WtLDPQ
hNz0+EeBHZcM8c9hFirn1s4vGlHTmJmiqgNr02eG877W/y2H2YpYxQON98xG
V4GhzVQopr6IVkhAQxN5gOtupMb0lT91gZR0YZngYYIdNrFzl05D2JuukTZ7
I5CC9TT0UWetFCmUGBZgxYNVAWP/J9sHBz0L22QdpXuE8PBdmHlTo08hk8Iu
lXQFIufrPaMB3kNJfj7QvH1BgNRTtMCJGP0N280JlsTfJVWoY4PQj4Fo1tR+
Ex0a3jOFH8YOL6a2gsMnb5z8cNlNYEpGuap3OXnBxoUFl+K00cEZE7b7CZFv
9uihwwGRfFSMwSgQGibe+CDV3yAymx+6MxykDDvDnyzP4H7in+tzqzg8NKnb
/MdtZ1yfkUSamYh7NMGeYzqDVBbRPF7NZqBEEtompzJR6xvEUbIxwB5FhnJL
AfEp1YNTCL+gM5CRIHR2Rh1hDugbnT3bjeixzg6ZQJWDeVxdQbpOL9dS3c4t
CJoRsuvMIlz9kG/eikf3AHyNU1284B6/fDpDSqxZlZNU/siesJFbnXJpdIub
8L8PFTLD0lTMnVj6z0AVJsfDoohJG0TLguJwRl2HAvHKay5hfaE8KjxMwYqC
aM3D7vjM4gcMxwZankqm1FCtGbmSy2J4yrodE82CvX4iaI5zntpKVJ5sHMgg
ZoiE4lbOUsE4oRpVIHeevAn+rSVJPXB3Ms9sVvkYyciyNfPAArgvI46rxNUp
Ks4EEDIskCECN17hol17dl7lM/mn2+si/6oY4Cb+onQDzY4N5JGKoAqQjrGM
6NzsZb3rAzKjFokqefRK+BwqiuBKpOBUrA8QKufAktlDBRQH6QZaKb2GtXxS
gRmXkV+8UxET/YuTsCp+CcXPM8QlFdPbCKQ6KKvR9e78iusfoJvu/NnTe15W
LhPp288mRlm9fHGWUBMl5cllSbJiAJb3DxVgZCjNFc6/eyQ5j8C8VxST0lju
tgo++ggrljGrYIgw1PkejGi/4cSzEwghGQvLzDm7zkQxhPWWhDxlskPtpIXs
NaS+x+DDYhXEzD7f8kHJmKqRqCpPzPMIIkhwSfoaQ7AbSwh2sFmGapiOzW1n
TXpsoUpyVBp0R3UtlSGm75LtQ5hnzwt+GX4hdiugJQGnJLpZxuliN9Jw/Z6I
yDmp7B9CR8dv2tfKv1f4AsYo1QnP1DYQTVCiyAY3o57A8VZVJ+G3NCWyvJs6
dsKO0GJhFPrqT931mC+DW0IndlZIMiPhpJI7HjDQTtxVT5XqghRbscoEBI1I
z7grYQmJPPOwOfuTQvjD//L5i5LBKAjcwo07NQuSnDXP3pFGg0Tu8CgMzzpD
ut7aXvlbEvLLDN6kSexi1OYXlh9RVafcwOGH+NQZ9i0HDi2HWPx+UAsyutMX
qQAENXM2dHqOwkIyJy4VNNCsi3F9lH7Cu6efLJXBFNSNGqho0/93iEF7vZFD
3unnvKk2arBpbfXW+ntXd09CEPp8mPnaGN9iEN6TIiwrxW/0D+BpS7y6MxKx
FSIwg9at2u0SRzOrVr6I/jI5dY5wLGnMxJhwpoDgGhXVcfdNhMAPpjJ5o/R3
pFMPuOYA8uPzifWWK7ueq35bff644zvLUdei1sFK5Nld+38LdAxbxsYdfmze
yWSl6OiaL6fz54g4//TbKjq6TchfX6PGPve8uiL2RKT7XwmBuWl/TewkJuH7
z+1/Y2I8mQvi0XkKVE5b8IrOol4vIVU6LWi4Clbk3snyNs1at+s7jlUPB92z
911aCqVKjeQlmDKsxEeS8j70O3v+v6o1E8GBsCNRY+QJF+FBOvKMgqfNn0HV
gvbpHZ2DRJXm9xix/LNlau/4MiniBUxplAHciIz6hjlsU3PIJK7/3I9CICMp
ft6RJmP+H7OXgnBdi7Zpjh5n6BVYYjGPxiD7+88AvjGPGOvADC/OHAcz53w3
Zpm2zun9PjJZThxHCrt1lRt6pxx+JvjeDpjU559LplpD/oWCv1xwZ1me+Tta
3fgVux7AtAXp6VgtJSro2zUgFP0fXY2LkoLTYSew9JXfQe192cUAMMhCZbcA
m6OtlAsNEb5FL7rT7ekyPoxN5cAqDy61l4T4mIJ1m4/Ldqr47vK0I9njeCQQ
RFz4iNi3NU1WUFVERi3jpLph899tUnqTPgT+Usbx381Ol3KMjwUOpEOYVTie
mmivJDYjULh9WCTfptkN41ih2YY3PqOFb/DfZR6gSmm3KmjhaMvNekatgL6f
6zOpawDlkP0B87vPORR5j+DB7WRwBDyPIipv7s9vz0vmF4Gn906XqZ49YMIM
x3attWVNW61bNQV4Zciwxtd9+QzLtQsY+DxXCmJpt/L5k/1eObs6X+TbxvID
hlqCAQFv7BQ3obw0mqro4IvLcQSkZDLrwA5ocwlhfIkBu+/X+o/bAOH6ZGlh
cY2dUXOATf9RQcT1oOJWppa4wXxrJ/UO2HRyHqgWjVAxFHcfwmDOdlZYhTe9
RCT8IfNoa4iHjuN5f1JFbw9SgcqjEax59GjsmFUrWl8a4ganAyyWIsh7MHls
kHh0OjdCjvuVJ9tnRHkwws+UeHyBYxl2iihI4o8NCzfSvehB4HmYs9H2Hqx2
FikRb1ZcvFZ0zQDpt9j8ZGytNYSY8bydnpXjXN/Ddi9+re3Vzw/fQRG2OvbM
u17CpFUM3eX0i/kRdCbOOPptHnlvaGoUiEX7i/owTjbAhs6KkElLjnxGkrRa
/t5TkK31UZ71whp9qN3bclPPxfEVJykNI/ZUAKY43QV4nE/yrQhXgfqYotR2
4S+Mke35L2x0thTuoz/XVD/bSwR2+FlTIL0VcG1rwjh5A7yrj2y9h2iilN2i
TzA0mcAtJkvpNjQ1ADw4tV9nx+fEamM3HdIs9TbAwlW703XYPCPz/GJlxdj+
aBl256lvHvBQ2xPeYWmWR9QgaIf/3NG+brTPpiau7/gBea7AjY2sAsZ6zc2d
efzIJ/i/CB1lP8cuXVWzdvZPjjPHH4vq914n9walgkHy0Jcn77bIkdRZigAX
zSzP2NtE+KYJ7YFuPxQ253qEGZKP0Fexi2xeNzgv/Mi/81QHiu5tkB9m1LX6
zYKIuQPvSCH52qhjRz7Iosj0kCq3ZMTj512hhGKLj3Ylg5v+gg5poxnHu2kb
MiLxqhqufzfvkXq1h8dtZzIv5Q1sqkZgE50nArCnmABXR6nnCsX+P7xp7zCU
Vt3OePp6ellUTNcKxN7IO6u9tEIxRXfXdMUcGLMsTYFH6yjDbRyodtG5VHaK
dZZNLXEBY/mjSKWLWILcIn0H+kx2yRpg3+lkopXSsGoHEPU9mgqxVWgqetYQ
Wtg7216edIGiSIA6qRzQUcjwcJFO8e/Rx8xhaXE1jGN31Ul6jHmSYuNcPJ2Q
tyaMiDsN0aYES+3I6wxXYjApxpUc2mHfBgR8JVUYhAiVNQiKbeP6NKHHl9ol
6MPb5T6wqYALhNxfONw+n0crcK9l7hU43u1e0rzFILfwTTVczeEOu4NbyZLd
RnRhuRXR5U3G+tAkt+AT3hPTDKMmD03wrFOerLYYjsVUruIVtdlsAKWkU0tS
SvCYZBRFytAhmVTBo0yR7coVACcorb1sPVpk2/aIwcq77Gi4oWjHP5+dKX3g
dHes54Xez9rylSa+LH8OlZa7TfGjdZPbnmkY/MCkPcuOHrq4YEVBSDik4bKK
ooGkIBnrl8izMRnZ5IKhAQd2IxuGmEEmEzMGpxYylcug/nRLs6ESwn4i4FNA
JFc91FhQU3UHNxLlYz/xYVqcfTbwBHhLRNtpnK5iESkZqzbtwQggIJ75NW4c
vHO5FgYz+DgHr9vV//wIM97GXaO0alnbZGy/2tlcfEwVT1ze6I6BZM24wSjO
Adv9LWhU9BbFCFq9gW0KcZjzKmPb79SZQkxYwsbBspZPDiCSM9IWkFXI3p0V
qVB5XY6RXEoeSGHstFfKCcsKnWHJr9NlaFSMOn+RKy76XfO2QZH/NIgEjsLS
gpqAUQZiAnuOEZ5DJjD7pcT7NwtXD1M6NDANK0y+pXpuIIZp6wv1v8iKxMiT
ySct0Nu3AtqGWcgplYap9nxYeHPaJYg/d8CUYRx7yKiom/RI1O/5SnVphZWx
3P/H4NN9sXS2BCMbW+OiJcM7ACN/H78TIDjPZPJNgWP6bcEDLsRV4cMdOZeL
vNp+lSagIEDR7ZEz/ge+qOX8eoJlnNQ2yPzR7qB6uLBut+l+y0RQnWY/WBsw
w3paRuFMa7vsOWjX2RbUsNGpcQReZi8Q4/YHFjdwq619gi91mjm3B0vShdOl
uXlZwchXw/B052YSYJZkACQPZ/k0gub7dJtFblpLctwZVRWr5TutZPgkCWfc
dFTYBz6GsGXzKA6V6rk+tmQlnXkCXTc0tPSwyOXmlNaPD+d0vFkk9eMlB1jn
SoPaHlirwXuzclt/aW4i8uQmO2rV9KVibKNhS3yOEu4YBwDnSQxrewyXeUC5
2ljr35fNPP9fu19U1DvSPJEosBkTBpgcRMot7oK70WGLoyFiS71yVJpw/0Ih
6T8kw+kj3tRCAbg1Ucpp6Nperz6zgdERMlkgS0I5fy2uk9rTEZ/fKEAzzhxj
x6+wCISCZ6TQX8MG3+8+jF8Ac1ik3jaPktvRlSHe/pKRoQCn1Q6buNIoVHrz
2tbK8gQCOwhOd/cODIbTQPTk7aB8XHzdNG6SOaDXQRn5H2VFp4roRoQpV3Nu
f7Tki6ntLfp41hzKicCTmKkEyjbVfB91mFpz/aYzkg/BfYHFAQ5GjQ49gJHr
Dp+DMIZJGfQOR4PGXV+owMBFKP3tuZySeqaoPzvIU2yq0aW+t3yFY4tU8Fzl
K3iEzkQ3fI/mxD2RGS9XTvEONyD+5bFkPef13lO0KpxkJ1JqiK18ZMytAE8K
FF/TkTdh04fo5rAy+Sa9g28YAr0ukcp4a7ZKdqmuZtAf+L6mg1V/9zLWeflE
c9tK+42AsXUwLDZ9fooV8w+uKQ76340xbU8Smh803b6D5dSy3vBcNOTdqykl
rRismiqMUINHSwlY4/XsgNvu3crZS95SJeXd7dkF1UKe/ZmxrF500xfS19yD
/ejPhamgjpR4FRO72t0IbnzeVjpB+L4xF9Wurq4w5X/rD1FDBDHSqBmN96vb
VvmfMt6bwPx14pTea3mMyMXfbmH5waJKzPNIoq1qa6FEsHZTXOh+0teH6nOx
Ew1jiyOpspKbFAEkUGkExDeV7r4jJNY17YIVqNs8PyhnBdlPSolGUqyn3Hpl
GJr1w6BVgR915zi8WthN4YndqW8tfrxO567b9LVzWWsRjKzfK8CR2Ls6ojc1
BO7eDSw9EiUy3WIVdAGQ3NZeGpiCqNw4nhbt/TNdK7JpdvxwmssfZ0/qXA0P
+p0YakjoY+l3k/sPZpDKJhi17iXoGtSfEsTd0goAVIVTiNRAAedVewjcFQQo
Rp9N8TyUx0oWS3+4oCpk52BVq+cnQ9wHq51R2/usWyNSwKBDR6O+yrDuZ6B+
SYMMhTpO0XiFKRyS+5FfqHy7ywGL0WKqaNLWxZj0E/dWpdy3/EnqZoVaQu9w
jWXD7LPc0IXUHGdRJjy19nmL4++JHDoEx1VFpP9wCa/ke3jJdm5/LrvneUWT
1KOiN9cAXFXyxK/ghFRVyJaqtQT+X1nwU9cOsjW4IZXuuPTQCQBx/FZ51tMu
rlQhEumgJYUiOYRSEEn28D4rVh0nMip9U4DTXYng26TVmcz+sx6Awug3UkTj
AfdK/AAgefoYZI9IUyVhmCdhOR3HzbM45DxbIG5GnJC23V8mgIVg0oHSjQvS
6nj/bc9/4Jix/H1SPQ7z9bTwNaoHAXzVmGikua1MriDADhhi7bhHoUbvuCDs
p9Wo3BK5wkSQNXqsoOs7w47yB2W2B3oadHKq/adQDRXrFkTwyxhM+Kb0LeLg
q+cGPb+Qrxhsw8OmlEYtJCoJPqttDyJGp1429eBII1bL5/PQSilm3ts9b05s
XdzuSKpsaEg+KdD2zBLZ1ZNp1e/8SPwtbfpzWBIUwUk5tEIJMv6LWucZyIWy
KwAarjuM7lh2e25rqQKDfNvEu+FL1NGdkFIlYSj+EDJRVX5dxffwTUb5ni/y
BGzRZP1skTkyIIl1duslz89aE16RKgeng6G4PAVwUnlgKsN1CF7DZgqErJny
3/AocURLR14dQ6BFCzY+ZBn7yx5UI7++rcCZRA/oh0Q4YoNiia+dfQR/+XND
xbyVha1carGuYO/Pjvx5UDM/3oHUSBFZpFSxL3nCKG4sPWJPy7tBNrrnXbMm
WO9o5GeneJLl8Gxd8NeGrvnM66fJY/h73jgp/0lETnsVu5Mthn6vl7WmR5eG
2dt0F/zVLDvMFLVoc3S/1qbstJL9DbegraJUuj0pXZ486+rpYvLEQjPOHtXn
gal7L5CdffGAi96bpXngaedrYx0HuSmsH0EWVOqPoYkG3aMvUQOAEb93JJIj
09FNOHrRJ8ITq4zkWyd2U1G7USEVldpSOBKowaNsvhy2Wz3IFnrAAFT9AXH5
fRlSdFo99yZrXj7kWh9CXbCLNpD+oqrMv+JEYZBNOnkNSz7+PXSuNFIz4O0F
2xzTPX3llWAwHo+LbNbLhUYtd4f57xwR21KNv2GkIhP64nMFZ0nlrqRDe8QQ
LX9lVHWGkSDycLCvztkC3gJVGAIceQ7K8PkykTx9RIoHQ4lYAPsikPgjJKaZ
oyIGVYEh0qQ24L0usGGZ5hw7E7ePhKhpM5pHp0dOEuAke8GIvc/97NMrxqlg
ZOyHoyVnbXzYHRjiMT0gRTdekj2iNJKMFxqe9eJlWfHQD3g17tmjrcXQLqOm
cSEurDcDMP5ttIoexPxv77XQupx032OlAWgE+tBwPL2ZWqEBQHA80FuGqVoa
JnVqj7WIEJOMHLmvQ6Ii/L28e+zirCjQbOJTGk5O/irgPynVQDJgKQYaHPZL
hXfsPy9H9q8ZX2WHtTs4p4S80ABsZau6qKD111iX6acr/F+cfHUovAVP6FYi
erSiNDltWQf4UK98sMCSsQIznirCLUSbFT4F7K/DPEhZUuCh4yH6yNupjN0U
srYpMV2Rqe+aLnMBWPG3P69+PpVhVqJSrePkbqngR1QiSMbzYZZvyKwCzGUJ
NH+yOUcuNioI4YKZC5C9J8QqpXjluaYpEIUQBnJwml7DYaqEx0vIXSI/MJVA
5IEWuqr/Q+0Q5NBgGhQN/hCdaDUrI0lRgCp9pNY0R/sBKsWVro7LOEANufj8
UDRZBgWaz4LRzNF85TUbbr/YvScLLrNWDqQa6V3vmT9yRydNBqsu/1xA6SgS
NVpDxaO7R79+L7cRApCptGWJM5wJURFsY7Ixrvmd9NU5QNKssLgLgGhP3nrW
BHp4tev5cPfy5qAwntYCd9merlee3aIzZ2GVEUPKcjV49MAhApmw3Cwy7NYR
GLlxBDIglkRWOKgMMbjM33vFB3KWWTDWrCtIUNlxWX3lTE9wXIj0uyVD+z8R
/3I8K7vzxRZdz1BkzU4FMgI4lZ9WqVkP0OuQ9DtSD68PuNx3R6gVls8TlFjs
4knGJAZhaOP2nZoLIo3qv/A3GsloukEtgKAElt1fEHrsKxNLGjTF1XU9W0wP
YQaWxzSnSuBiYfJVKzByKgM3G5+0mXqTzObKOUOKmobgrgT8/+vF0zMoa/BR
5CWKsOrVy+Bb+37snCQWCmiQrzu96/yjazBIByEtCYIyFdI8BrkZoVTs2YbG
b5WpPY7Sogf4chVioWdZK++bqRQidD8JCn9Vp5SExzpWSV0P/LPwKalfUUQv
jr6ahkzw1QaRiJlAj/tUx1KQB4Tw9jINPfDMFZs1cPZL6lUlo++2z887Z3aN
ZHyjuCcgBX0+z8HEJeI8hPM+V9ftpojLb1PWMbP5fwuhDWyMbh0jcLnCJO0g
sri3E7j8g5i3wvfqrbT4T+J0FKik2eiwtAeS9FygiLuC5dzN/hYgKsmYkM8k
H/Dok9bv2Ei00U4ERTYv7JsoVKJMStQk+z8koiRrHHcg5zmAW2lrjCuny+Jm
HG56cZlWUkOFw+VyjggbD1WA7A+L3qXazTdljZo0fALft75DJMbXhRgbXaOc
1/i6TQxcVHIxbGrgNZFd2WXJJcpg3VStvWk/7J5a8vqAZwDi4UXJPBuVtdbb
Jl0GLZ4VEtnZNYlhFerJKlOzxjRJihb2o2h5asCTz0pMyDJJB8dAkRHb/M6X
A8ZuZvNdAwnk9kMev88oDTdbblKKBp67qau7CwU3iBYgSBxud98wWfjXEVs1
r33QRtUT90we+C6n7ppk48zkL4doM1V4FnYZZJHOGRaaMVRoSokaJaX0tuVZ
Mlh8bhLXnm4K7OEMy0fgn48ZYgt8C6IXDMMeJ5/jUqUxY9iMeCPXPxUeW+R2
2SyWHG2cbi+s+HkwS9TVIya7OFociCHblzks/sXyQzRCJNYzTuhtApMFEaTk
LZS7yCVZHZn2UGDKXmKT7K2VAgxyC7CEY29gCtHIr1O5WLaJw3clJDp58X96
Z1+NLwv9ZOPBltGEa0szNlxwmkjxeTIV2N0eG2RWGELmEsqltCnATXhyVRXM
I10ypqGMVVK1yamXqHAcMXJdk++0hMVRXGMV4sQPf39B4L/YscsQhzJRHwDh
qX4kTvhp/1LQGXgDXxn7XpuaYLGhasBZYwK5NY7g3l2qCBpEPtAfwQ+e14Px
3KUN9I5ESXfSrdmPQL8tCqP1kn0o+yXRNiws5Syv9dbd35gzN6aV+SLYMB5S
L+DF3K2ndzpICiI/1XfOxByPPwP/4szN96xW4BTz6kzveQFcfHd1aP5QG1M7
YM74qYtJDzLg3CbY3q8IB5l173c1D1NnH8rZfmaPRrgBsaL2YfC48e/7ZwGS
Z9gvlQ+uipFloG/sQM2oPxcVbGe48qFtqBcZ7ebrjhRXa1s8DuJyJ6dmZGcV
V087WbKdhJyONuyEjBpok0ioq09qWNSuadfjza7Zs1eMBEcaCxs5pKZ2+og0
5O5uShbmrrREASwZGJTSiWCCOElna6GwdlAp8OhqLzWrUdIGsGTa5I40Tpkd
2DfC9JflhncfkwVIlD78++t5TO5HB5k8r3GGwqGOk99bLukvqoEg0pvDHQ3d
YQtIbNceh7EoQLvqztI10RQqbxzRwiE+ooCmKDya5LqqNVhVzso980salKzw
gGqoo/Sj25QIyVsGFhd59jX6oFYSxrFQLq5CXF9wV1AZAsI/6lv+o2/ZRLcN
79ciBnORF1+o362yJCgo1y39CmP4ZAm6pJ6+iFb6f0v1xvgKu4S9KiAQaZxc
9xuwPSA7ycNgVHFyvBm6OltRFh5iXdV43e9hBFHie+6PjTSCF1YbXm1muj6S
V3sTTNrjgONe8/gMwTch584jfbogfAkwT2t92PovhZ306wwkUyXwpivfyTSx
fXwao7c+RP8vxMHjMe8lPAU/g+uFEGd9kJbFk2opswUtRxKBQl6F8QUoR83c
/L3zZihBy5f0A7BlRzJZWRbIh/+FEVk+AlTzASFSyWv61+DJD0RSNfuF5mdd
XY0p0sP2zVzdbImIK8S82R8OD9gEnMGbZ8Jen0D9QuDQdCBr2d5tjpMnMCaL
Q53nnNcJXBXqDjQFpXMOxoWd+wskNDCKihN+/2VYM9mWz0mwisNrt0r10FBk
N0r2jlTW8wvBtvyBn+o7KcEer9khe8dX/tfGZf3q4Ks6LYG72qxqd/WiZ7vs
loLLMi/DPY4K7jr6TM50pc2JbDf+Ey9FcPRHRn7uHYREJ1PJRGpijR2Kcg5O
kYslUF1IMMIBNSvSZLjut7jr4qzgA6BFd1M7DEfLpAPfTgKdCK25ZO5/JQ17
FTOlFpq0KFrSmG8v5aCC1RtT3HZ89vk1PdegSaB3zrNzi3QETzoB8x/1i4E3
jnIb+i80bVkPHo1Cdg4WGatwcvbFoQr2kGZgX2qdKYBoQb/xqPA9eRuJw8fM
VT9qDfWqcGNCfdFS9imj0q1hmdSUYzfei0NkwKS3bLAcQLrgEhOtH89yWhA8
qqADub9VjZEVYQ43mZGXhps8OUZEV8jKeYDTTZAT3eK2aisgEQTVfapiWyym
mM+Va2oxG+jSvaR5h5TczP1GZTzgr+b+hY+sR51ZbGyrNH17b9oHzfRMbgYd
Bd5umepvrSP33BK6ssF4g4JOB583RJlHG4V6S/iXI2nF45Sy19PLBDFf3NQJ
HsfQ6NsQ2eCjJ7dk7l4IQyp0QLUUqH4fYrMeHOPx+3XuZlZEssgcbULxbuod
uLL3XXyJwHdl6lsS00aw/3APB7HVCD3LHgsPuPIh5I+aPvu12FqS515+LFhg
6JER4WK27yAO7cN04zh0RSYjF+Uimw01SlnUVfdYLnGGXMWRDUKVNJpIDH4a
CkAyjLTDOuHh/AG+TfLKXQojfbJQwF9KeWV6FbGz9PcP8Drnts4hQKsIqlLx
30MiMeFcQvgRRb/fzspwuRaZpiAYeKsw++x013jWH4WDCYy309MPZHoXN0y9
WT09FcuPjGfwm7l84lj3z6KqfKm7UdYVvNxNhXvAXK2OLwmAhfF5v2jvUx2t
h67CdsafDMEiMebIFb7AWzbOeCLG00/aMMRBR64DKE5/AwFofNUAha5CADWQ
R8b7ICiYWeA5uZmBuJ+HsCPmcVvNMNXzr7foefHTtRRM6COVBScLNYxhZVZ4
VqVADVeOqm6DoUIJlqh4QjmKtGzhDNsGcMGDKRKApd/iPeEhljtXzn/jMq+7
yC2MpJmzO3oKH5sCCMTVOIVunQm+tBk0zevNadJ5s2MPup3lQcDmeHWb1daq
zJl6Kwpmyr8GGT7wGFpA0BXDKCTlXGNljI6NKUIsmdPvgCr2sYZciU3JYGBz
ZAICU/whC96t6yTEGhVo7wXx12vWOMgh4zPmAUpxy6tIujhpETDIvmq2XHYq
hOqEJdv5mLGmFi6p0FU+GJ+P/8mb8ZMrvbqPMvRuGBkr14+2Yl1I8qHOvz4r
jCM93xHs6S5wMuIxo7zRmu2vyvCR48Yh4J/3PtwAlcdfCKUsk2zXLSlV0uJ5
fl9ApV7DsUxnxmdDwcebhAJ7lcjER4j/Z4Np+jEN34x1RtAvZJXN+SUIouDT
N5/tpFHilIumipX60nK+HHP+A8QU3m4dGKxidH72KrzWe2h6LfqQ2wTY4yqQ
n4FSSB5HCdX5zym+rkDYa+cV9aYixddT3bkBPEf9L5FgtPhh72iCRTn3fIS+
8zUYHnFXs5Bk8SdvkJc7dy2d61ijYZJYdHte/nHSJhT1HcBzHcYOuqQTuJOH
iAoU8MriY1H54UuzGIZ21J0/e232aH30p/uv7S8jPv26sltn2anEr7TQHVrb
HTyIZ5xJytOY/L1J30yW4ALitpdriTbvWgzQgYWJbheTbkLvo97BK911zglz
0cYLAHc+P3Aa1keWvHHLeUeKucBB6vuTwHA9Tji+4vqKUNiTXf9pa8DT/3io
fzAzIaKq5vmit6Ht8aQo3+EDI0tdfT1h8dS+Y9OXEYZY9sy+JLcMNo7iTX6E
gYDdGNNZQZZdtHL7iZffc+Xe5+uSLxPE85ORTWiB8c4l2/M26euamJi9W03m
nSI94aBWsG69uGx+90xRUysOtr2hr4fKbstAVT0moSfltFMH9Gx3MUu1XYJm
4w8vni/veA655BCAKiCDsLrzSstLYgyrc9fS91POpdkX8vDWtAlpZbguxAR5
YX/DzzaM1yXjpB2JtqUljkEehH36wjA7tDeCVfur0dds6tKDG1NilnDk6yKK
5o7oWkeJ9u+3evgl8gPez7WPkcXatHVHySDSQNA14e0FHw9npHRCRlcFYgxy
0qSTjWg3j0vpy0PmBRs7ily5rRczlCczw5CDeVxQfaKHJGKUT61b/gFQ5l2q
+WXt+acbYHDEhTKM6mjv3KRikI4/4yt9aUX3LW6pdLBaFw==

`pragma protect end_protected
