// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
E/srIPFCsuEV41+dtWBdV7884y2aVwwikDJIE0vQ5k+Yzf2Aa80bl/8578HVwvKo
SelFQsIKc94RRuXgEuXHBOxS7cuNRHgZ50WzS2oA/M2bU1+86qlUzGrdxcBE7Nje
SGzBIhZvS+AITEJLARBTnJZ7Y9r2c/9dV5nwdOqoFN8=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 30944 )
`pragma protect data_block
Hx7S+ycILQ6yqUmV7SE1v4s1/kr+gSEHcLhKvIzsncCkQLTl+K11K4fm4WBhQeGd
49UXPSyeFRSNwXrK6U/KU23NsJW6IuAVP1eSCNPAqv99TNq2h3tJBc1xHrBwYKkP
/k4eqI17vVmrqqlqa1RrvaCy3cZhC4v3va911O61RdITDd70N+VC+UN8eYmTpsAd
ZFSmUbH9dZO0sgqYsQW1NNddnnF5X/5bqqkM9kU/FhVum8ZJKU1iwmLze1e2SBuk
RFUCDn3RL7ZsgdweVYrK0BRdNgJv3JfXHzSeZeWcqfYgoROj2K8hCldbYdiA1nRW
M3dhXV+UHC4ZTrZiK145UFES7gLiySQ07gM6GFh4hoUaLEyG+MmJEv0K4nqhsAVQ
zLt1EhVE/hbIDbltvyil0OEpguN/lUG/8ZwWsm5nXDsD8xAo0hd2XJST4ojjhIOL
qcGN+pQ6DlQeThN+6NIDRU6VmFTzEFEE+/lzZ2m+RnJ1JM6k0KyH9Vwic/wh6LUc
7zbpuQWwCxfvkbIs+iQg0cdA4Gn55dKJXoX6nSN5pLgNmWtF6fFUim/4yy8HA307
ukIygQVN9wZSojXzOP5gWzkEnpEPYly4N0EZOIF0XTBbR0RMFFSaJenDayssvMeB
L4EjSPXbLS7NHoD3SjUEe3vKrAoC/Tews/+yk7EwdM6Dd+eGvKDQpBXa0Ag6167k
h/D5wlHLiIB3iVv/f0FgBBEfaSZWxtAs1qDS8cHZaTymLADs6zt+Xzy1wXVw2GwW
h4atTIKXK/NmLhMwc9yC3AGQJIgGxY2f3PZn8KdD8S+KKjqg3d0GwosWCAtp3Kx0
ZPp2VOMMl41b/F54LPvd2sBPob+3PmAXUnjEOntjj/Qdy5PatSYXFw4Uu1PntC+g
1KJgbuSNrO4xRUVQrinQFQvixIH7Ay/INJYkVZj5C1eM4A1SEmrjbMAjIfUkoHqz
kcvQsBEHyAw1wZzUy2+gmG/gfNGfl07XYS2f8Vvdx3PiJjVoeyNoNH5yhyB7Otfg
Tf2J+XvyAEqXGAi+yFXLal3q8/YNVMQrs7eg9Kc1aY+PVt5eL0yaO5jh1L3gjTgr
geMCrMOp23xwe0y4tWoAlOLKvfKzAiB75J7wI1Ud041GDWf38kznI8EdHu4nkWKP
/RN4PcosSr6wYsR6Uxkx2urJQMb/Q156ttAK+ybzsdlgUBhOMZXNHimF5yvVRprr
m7AGUCktJXzsUWq73IjtPVDeDRoNXlEuPS9cfAP5n4dlcBuTzRUBD0d8ztcBo9Hp
HrphALnaPNHySfjBA/qqmtW4fMpsEer0wWabCf3zV0dJUBtmCDqDvTGtBfDqHl+d
BbhzzJhmavvRgPAnj7Wk4mr9+zz/qCOlCfphxrn41QqsXpCc/OowNtc1Eb54d9uc
M4oNWIKFBSE6jPpYGBguT6cS5KWwnELERdLCo35EnhIdmxOnCOtdXcitz/qNKroL
WwkwDcnKJELKJ4+J96mHs2zPOIltDHobiALr104giQ+DNqBJh2+y0gK65j/7xctY
MRfitxzOwigN/bc823JDGlxecMLqEhfzCrTmk7tf3bYdVPfQjx5IXIRTy+TLzjE4
eINrkfEYSWp2/tuzKBbHtWCpcwtPzFKIHPdw6r7hLzLvkciW0IgIJupv8wZ9w2NQ
M/0PDDdicms9lo2xv0aDTxPa6qVHRyz7s07VrM2McMQ12CKCz1lkzTWM394rSdB6
WqjeluyVRbSgd9xzm90FgJrNT+5bmZPVdUS+/phLSHV/ADAyMTSKwH6PoyLPeSSG
IpzgzpnMpFpEukQdYPOqEPCJLZ2mOnh4b9gBPPZT9NG9++pxspPisPrI9yuNBusn
vugVI6+y+2PSOshuAzbdGHT273lS19Y3hKQj4I0OayNDBwFlDD/V13lBYaAG7X5b
drPFZURZZiYEoXJ2MGI1P6sWHtMehcwsXhAgirPrZFCNbfZ7837DrqmmiwMv+xrY
BwF/GShPHH0UcqH52Y9rN9tnCHu5IFEF93qygSyiaTZz/pXcq7XJ6/UTI0uGkEyw
ucLFD5nMIZyUX4fen/Pcl6uDSqNmzWKyAydnTb/tBmip2cC/gtbmkfWS7syyLc78
IMIrNdu3n0kBUbjL8tEUQ+fZhtbS/ktm+q3OvkjW2YWGdWJDYEQV0+Usio2WXRl8
Ij4aVmW97DkrX4WE5rej5Z0XROt8dwToDtTVwpk1oPf34MltgTDwJKOMl5FcQ4IC
a9v+U97Mf8hRnuA+LgBNfzrxM4FMFnvF1ejBq1Ug3T+tHulAxOuFJ1Raz7Elv4mq
AIwLNC7+nrXqGmuNty3F9X3CHJfdBw5liZAN+BY0N5neU0AMcAc70rJKkAOyVSFQ
8YjQMlGCCtabPvrozUYQx7rroodDyQQ7iQ3GQhf1bMvg7kkDvP8R1DXQ2c+TtNCR
f6yLAHoDeG81dMPIVJhIQTP9iTuc+6iOlXH+ssGO9iiz2RdU4SsxV4pbCEQB4wNk
9MXJhB0KOCMx9OBP5dc3AQyUiSqYlK0PxSZaOAEYPIbO0JgEJ6NUc0K/eTNAYYYC
DbB6BOhBviMbQcZHpsaWMwbsHkeqzfiWouZH7qFJ73jn2XfgIPdtgNswQ2VfheG5
JwcTMip4Rz4UGsY2d5pqVpSfjpEw7aw1x77KhnRZjstDR2paqlstI0cCcfMLei51
cHPcv2uAEoI+1b5SAy/YRT1x9F96pmkQniFcaG057qGQqHgk0uSSBR6YWwDNgmLm
PR8+fwKqBMFuHbTw75LTANVEst1ZjRG2CvfK3C/8jDCmOD+Cd2MU5UoPh82qf+PJ
TW8t2CcLgqna112kuaaH5y++0FdQwWkfrNw/OLvSXFMjnsdrC5L+GUtezWW6gqg5
cmYyPM9kB9gxFmdjJ2CkfGTjaXGPL7nWCnatlv/DgWcbw979SleSzcjpe2xqNtrp
vnvNWrLQfdbipnTg7pdMum57PEmpGAQYxJyxd2WJ3a0i5LentF4FkuOCw1meAFMy
afwlNR4oBdCquJ3gIzpx7zKYsPDcfIVmnDz6jFtNqLv5FJEVnS6NHtMXeAJzVYLJ
DLWmhm4UmInTaVHZmGlKAF+/VknTbZhrkp8G0r4i5b2m1i+Gb/h0QsvmVU2xVRI/
12Vz2jaJ1wVPQYkU2xV1phVucZx1ojXKOopbvoSoK+UgCJ8GTSLnJSuCz6QAXUQP
rx75hMa/C7TyLLlbY8UDye2amv0re9QKyqFB3Tf2uTgeo+2chgrsGY9nPO2JOKab
yVt7echew23ylloLgbp7GNPdnOaRniSdjmHfQnP6Iqf7/DntW6N+toky0KEz0/1G
mB3+EuvIH4lqTeabRZa/SiEyjwOref1Rv7RyLlj2z4U4i4o1EdK8KJFddUuSDcma
xSEhJXNbzcJdyPywdux9tc/TU8RkuQAQcomX9DBt6bfsVFDFmOVRVETWghCclldO
BLwraK7dhRy0B01gDWrvSf/9ZnpnM801zYI4gCHdxZv1WnaSYTC6CqZRa0RLwfch
1cmT+Gu7+mvWcQJcxhW30MzwUGrHqxRIzbjl7jxbrLe1++joXk6/EQRYmDIGJGdA
alt7BiR68MLmAiHKkixkVr9alqw7xHe+VtrSB16gcfjZKEJUMfXgk42CZQFJnmEK
YOrTSiw5j6q6Wy2KD2FUlZQ7Pn7K5mLnQoWwua+YgRZw3nv+XNVOVkzlR/J5G5hP
XSjFMn437Nslp1d0QxiBYjhuDRET5f9rbIO7KasS4kriorEq6Xai6uWEUfe36BP6
ciYkbwgbhDQW6aq+bT2SPPWHMp0caACM1Iw6HL4jkgZc8wuVyOWKpY60AO5krSYX
s/r7/VPtetTG7yZSy9abF4HRcEgO/ZFdZC+/tLThYVTapJf5pehHulfHLENqPFtz
4AcvyCC4cwxX2ToVdiXmT0HFeNWNMUpFtqU0hLa9Q+nCOQ8IYolUhauxbzxA/Hu6
rggrgqxiBPtHaruI1867o5Sd1hb/o20FiVLDAAbz6o/VI98++X30EwbcFVAUU6dX
uAiBA1AiACNLe9Yussx7b5F46C5o0nPZDhPa0yhHwhzEGlCd//CdDVVL79s342gv
q9nEbOTgFszCfCMykpMAmUn28fv1mGm7919AXfYVzqUSydNonylN00s1Bikx8e4N
1aPqLuxXgjVIPMouFmXbk6yKlXXwaD4+ITLMNm6UdDQFgF6qvra4rNqE0Xvy1UGJ
VLS+QKHHoo17BJYnmZKj2mSgbcywOh/K1ctQ3P+br4oDbzAIgOeIdkTcMuOvsvxR
RLkriFb4nViUGROBCtskbKDfvjGVevWknFhkgwf632XsHSyM6UUY5xq4JwXaSGto
kLaKJqbo3unq4q3oSERV4SVn6RRVsv4mL6EW5oDAkl0A3WkYWDG/aMokxMUyFJJ/
+LsqXSgwrFX6BUsBh//+Ifv/CgMseNQnrhZs2IBr3MtoqBtwwGkYFRpgk23Nk4Fh
K9W4m8Ws+3oYVLlt0rMox5/loIertcA+fKpDr2XetbiCpsfWlVJg9Ecb7eZnnyN7
8v+lwiFfVDIA411ulokNEyuxoF9WFCPfCwUhfFGalfdQVAnfX6i5pjYRm+DxZ90E
Izk+pIInclgjgDMViN7xeThzPxV+17a38ayjY41QbrgjqiElD8dHuL9YONCIE8yH
eZ/0b09jYF9LwUIAecBq3gsD4A+bTikPswz70vmBKs4M0Wg0cW+Up5gUu4dd2+lF
XHPNGrN9NHvnVoQuPsySWmNXoWtyOj680Qp0R80za4W5gYM4CkA89Qny2gHq0nPF
epDx6XKKx3Iw27jv0H0reTaQFUVA3+OI2TL4LkrmItg0soW9qlrrDK3pUwmG8y3D
8I1vznqsDMTLGkPQjxu7d7wLFN3vgdJx/o2+7Amd44WjuQo15upkmu//Wf4xA7Or
z8OegJmwFR5MDVbIXfkD386/2MNi5ydfelhnRf0cFEc+bYQ+P61M8BTnPsUy615H
bvexX3a19vEXzSIrh97JoMd7SXgBKHicHpXyW4UgATyj+iL/jdd3wYwGbyK55tNS
tRboRACBmcnqUkTNePs5/LomGvBUXvWgqjfI+3lq1NcJIpl18+F2EtkQZFWcZyxY
VA6e2sknnWQP+jBl/yCC9qAcXXVr71UBR8r8rJJBEXAjZ6OQ4b+qTi2TbHrdHPKf
rcAO3FAjE+6I5sF7nyG/eq1+15zbIjG7mJGGMdGHMHYeC/bx21eYb65plN3/o68I
Ju86bpxu2Cjw88jm4QoB5I2cYTHtMkx0uOD5R9U2ZhFg5fbknkCIvOnMwwNENnHW
Ilv+Y4W/v8RzZ9yKIdZrSTsNIo7Dfu9PnRk19i5agGyc8RBLJtu37pvEQxZYZ/LW
bHg1f+R7gIHzWImdlWgvDhQAGYwmLGjakC56ngOEc1b4jq1dH0b+KFPBigci/gup
Bn1JH7qJIX2oW8L2qAmiCi7Ol4W/FVPE0UKxRgK82cj0X2RjpLdg3htmUMX1dV/K
fL9piUAh9pNSZFVkK6sVxweC/z5VIQhK8V7pFy3x0O3CqJH3JKOeM7WVds6PxwTl
l3ES74zynNzqMWwxJS2Bb2P3f0BysrE2fCF4U83CxsU7p5fMyVV78tw0qH4xuAOh
9Q37DFxF3tVwmIruyLea5+/tzltWGLfMLggpbv00BD/mzs+meut0RunSqshyIL29
kzDfZFu1gTFYzItXxNL2whr+21G8sd7Tiv9u7rho45w2A+2iYVvz+ieHtG1dnBwU
pwzpYYrnPVicTaWHSRhMcPKdBLIVa4zwU1Lmi6/DJpXiRfSG7zrXX0A12iclIVaj
ppd4i3hXIlH1GfNp2Vw7xVEWf59cbbjmrW9zSLP1p8qdO6Fdgqw/OM3rYiNO1fTS
qDeDDPQmuJ0SHd+ybi3gjORkfP/6TyFapl+LizhUL+Uq7vN0NgCgqLu4fZWproM0
ChtmrOiZhJ0lTnDuJ2aJDA/BePXxmyUnZ3OeSNxlyBv4guxazy2zC0zutxn/e8eI
HoIEDUpvw3R5vseNEVeHBrpUzhKkCe+XHYjXoyl84jc3saEmBl+JTE9kQIK8jwmR
7i9c6M00x8YhQqYfPZEToFH6VjppE7sAp5TPJYbUo05xvWOUds/wzq6MPX+QIfjQ
Q4DqGkEuT69alvEOWOzuq2Tr6BwJQF4P50x8inxQvuqKjL0DDmSy5gwwubH7YUpz
oz7XKloY23MobgJWZt1iCDsG+s/Z52XlIarSp7Lf7v7N/1+4m5jmAD51E/IClZ3l
I0CkU8wog3JPhGOyDRKjIufLXF0yVtQVmj3XToF32K+Px7J/gE/DNTS8rfg9nFnz
Uh8Sqbm+1X6jv0umRzo8NsAOJuriv3gYl3eRtePje3pNrkTs1DQgHzg8FuakJIkf
MVi4XgwQDs4gtjLxexqbT+sHKvr10JmNTRKbIR/Jn5awjtJVn+346FTepC8C4ekw
KX9cOXIgMIoyk3bV+J5jIVjYWdIrD4TrXI+V6a73aQvL+kCmEuwfMzGPYPd4M+Sd
Nzwf7PjbkaBpAi6dtePmkf5ohTT8clp5QuCNIU/cXz5lN0N5uAway53+s9fxzCnP
rDvSiNc2u6fsnE7OH8EpUWqcSwn2BD2Gt2KRoruehUpgN2bgrpB2lTCNZWrwE2+j
owl28/Cq6YeiEWsXqeBov606HAkqxHEBD8Cdr7lgrQUiSNfpjGycW08+7zah6gea
Xwu4P/ZdpciGkkNVKsLNGFc2h4rf6dDpIOHre64seEWK4LYHvWC4gBoyFsQcQQiR
/so/HQb9g2dm3Hfa9hu7QoFv/h3e+WeV7luZWH+rQuX6Vsz4+9l7NN1ZJhAoLAOv
rHSwPeok5H60y5emEzxN3QE9nRakSlaOiF1Yw1j3yvvFsND6Fc1GmYUBlWGQgYsY
fDpz684yjg4z61NALUED90RUQeyMt2oaeQ4c0kp6cAdlucugSxg9bwhsj/iok3wl
Dk2khYyqhrsiDYe9wieDN99VRmqD9dqW2Z/pl5Xn4uzIR+IR9uNVzYd8dHsqbdTc
5jX1DEW/lNeTXb7CCLQc+wOmxacSn8Vg/1eDREu0pvXZmupxWEF9LJLpifM5ow2S
Z4Pb3rQjefCtVpnkxxmy0A2trHJVGH7I5mrPIWDQ9wiDRMzqzXcVqBd9Zl2TxscQ
sslTqdM+LpNbnziyv8jWnHD4/LwVcytKLov1dFyH1lNjYs2Hl/IoFvd2DwPWF9gB
eg3M3+ojCtEsFTNpyehjmf7g/ucSs2jo7EBobqblzK8Y79zwsduQ6kgo+T0VFiMu
ROwk825FYb1+5zsFTUtBPzaywvlFVEuMOMrP9mWXmm21E+J5Q42j7k3ipC4+ic1R
D2XrpQB7bIdl8cDOuMxCVopUa4voB8UGS2MLQtJ/g6rLBqbpt5wAXLYm1ak7bZzD
tDVny6rPHTBy99FFjBzTQpt7DRuOxaEwNOLft7f0bQfdDI1f4YBWveAY+2BsN7xB
6ptWvK1QV5Nf3JSu1hHPjMVyL4l9Tkq6OyKzlcgYbj0Co1NQShmQ1xQBUX414CA/
M2letMd4UtGNb/AxBFQ8kbQBXZ/aVOTzCE6Kd08JTfEqrZxiuN+4o7ti6qhV0MBG
kM8GKOymxNOD/zEuQrABq/Ux7b+ywOz2dxnhv5yXcCtcLGEAz0RWgLPCCmFkv7pX
iZLOar5z5A55pDPiRVvpyS+l8SlvMNmasqFBNYSV9Z92vPcO2V20iFO6YGMkWL0d
F87JMbbbjJyRAgwep8P69Mq2gitwF9Mo55jw8ABRsdWiqRNPuvUz2/9wLlnP5raY
lBajzHRZZfPzR+CfZnQ77n8oJUL/i8/UNR5jAdbaqa4BuZlgUfNE/qyI28nUw0dS
qyyldzfCxRZMzZmL7xS5W96vtd5g3g63ouUfrXNuO14usEVZFx1li/K67rep8HlJ
KvyhRttH3HBGzHpMQ6vSzoHgLUDIk4dsc2G4r25bBofADHq/Cr88SwAeEDmLbkPb
B1F7qgop/xd9t79HzRMRjD+s/EcdyPAupxr5DLFp74xRqlZDQwGxNOKgxJDgOTRn
JI8K4MkTp2Lu4S5u+eI9ssmE5jQzQBXoFXsxNv3nV3zfr1HhHNY1Xd68Ch19qa1S
A24OXjdd5GSJCFu/r+cpBfyoG/MKl+sw5FjlNrRha99C+R4coxj2ZgV1dnkYijen
lERQNrEnccq8pFXLGAQzna0kT1M16uFOXD27NvLFdSUjj9c3pweXyvly8ihu/m4W
u08xSaf8Hs+danfOWrOwveWtPtoMSH4yLwI/DjuscLOPlXdZiznNApkPKCIKf1w3
aChe6KSewnDtZetV/fHdLACiW1zZqG3noxaEQdopkydkvR4hqImY0ax6EVcMl4kV
+XwrRXmprH+rVCf1wqW62MqT+pV4RabtA1U0e+26itrVcXTi4Ke3TLhWps/RQeeI
7oVQPrtmTSX6Il1wbCgxHfScd3cPRbs8gXWthAatyQerjKNKHzDg003fwuUjch4a
69DD6fR5DAn7mZYD7MNGQtCv2uLDbJUWKhKLdp7JKyftqSKRyKMKWpW/6kKBK05n
0LfmVaL4x8TM2rV0k5ui8XItfOTMAsxgi9yAXwRSY3jN+DFz5ZQt7Gknrrf78rFg
d0mcu6WQKh+r+RqDZVf0qh57kUfec+jo4xhGKse8oT0R8ggw85i+ADM1S6NQr+yn
jwwT/W3hxMMOaCjVgg0BqL/ZnS4y2qozrLtHEg7pmFlrKlmTCjP4gP7c4BAHuBbb
kB2716fyzapSxOrF9uhYNzebVuekHgyXZjFvztFib5lTOeIjOS2cKw4Pie5NvKWH
3YRlQdSRyDfpQU5vE31UbMpeq4CVMveKLYv+u3t2U7L9blRRG/nCXoQ0HD7W3e1B
D3/s9MMRizrw7JFsmjHXvQAmcZ5/QZpZZBvHvUFriqjs0+eGJVXXVktQ9e3MuDGb
mqMltor4YARZ7GC6vdHAA/4mHg+RYLWmRxPNs1R06pJQ9xNx3AqWdRp0hVugwy6n
WNG2a/kMVxm58fKvjx59OlJEd2H8nLSby38Hr6DZuxzY0ag9IU2rhoDY9oXFF+Pt
TpRMNkz5mbnjZSSubez/f9v+hFKWGeOlssfp/qqMflu3HImL7z2PMPzEQRqDSAOh
xlqPV+A5AdIMJndaFpOyMJQN8Rhos7NPGoHGIrKNYBi+MMHQQSCmm9FACmXiY9Ki
9g+JjBbMO354QfP8bKMsEjb2NBhdkP0MJmnnBuhFWUn2LORdKTeZv/TMJ8inJH9j
6a2AZyVfUIU4YMdyY1whKr4ATKZA6tCKmxLJpRzp5a5Q3f+6W7dHQsP+jOI061c0
j6GbzfDtk5AwQdKvZt3VBQumr3VpO6ENR+7UnxZlZpJmRGDgM+Ewd98xOepTo0ff
84pHRjFbjSQkwqUq5jhYUZq3WR5vkNoRH4DlzfiPqX47O79qrPgxNIQ9/LRL0gk9
F72bPhH61vAOmZNXeVw9/rGH6CnLVtqKknf3ZaTwXFAKhBm4lh44uh5vVEoxOOO8
LLf5K/97lz2pUNOBKKxQlg/N3iXOBFSTwlLY147vsJ+/nbyQSsBo91AnDFAXDRMt
4HW8a5gePgZGqdHTsZMqVSaDIsMQ5flHs/szyx62p41CxWBhcgaomBI39W5WFKgJ
vRNJudPCsP8qA1Nt74N53LZMDUTwZVF/C/H+wJw+BePxA1Xm5DzAPLbcoPZm2jGJ
o1gb+t/aZWbtMPtpZXv+2qXqzLC0LsViw5QbrvRcuKmGJJ4syc9sU1/p0OMiVhPS
BrPS1JPzJYuGnBoRmF4iUFFOL7KB6SXAK6yyixiFObC3KsjXrlXfP/NcnIZYYrRh
hAio9LyUkUnLSZolZ20d7s8DkiQ6+2kMHkzioiNcOBtABwRLKr4gmDwbr4AcFZiX
v7PsUac8e0yEE2h+TX52T9Ai87cMrfX/CPdoLg7YV1pF2iJLlJDdcUcuiXxMhyEx
fuypZWwOvpJwMHgOjHw2Nrqdr+sBM3s54PYqHrwXWl5EMebfJeadZkmVCvkd3DIp
nXKPIp5NTdA8A7W15W0WQC0+SnqkJp7E6MEyKsnNNd7JXeuHJ97GbPJkhucKgOIw
qnosJDedVpZlMYifPFBW5J7sgHAZCbR/2ZnQ8vqUW5aCHCLYO0YhMeh96cZ1cabX
r2LJBoFVs6QEQQG5Isp3q/YtMUhANrRUUvCByrhReCbwzHlpxsVLjozjSHxlO1qp
HgXv086vNQBvO+KIIa0QdcrsCZzmYaQUGLgOv0FxuNH5pSUgmSWFKfp1VW5wu2Dv
zp/7VloPia465zXR2mgo7kG/8LlxeWY6xxOHZjvqPKaxpD8fdQoUFUA9ls9fcSaI
DkpebxonnCR3yEKsyrQvS2a0SRAFnEEgkHNQT9UFNIhE2/gdIN+RrLDdY28vUXET
q5bSa1/xnpJPx2/VnrCTRoV/vI2o72T3AcArNtevKGcuaqQq31p7VuTLWafmJPv7
r84/LI7JENibJ6q2rf/MwRcrFhqRSn1i2moSGcinW71Ib+vgv+l/YewKyK9RBTmp
hc/D0Rnpr6nhxUycLjiWMlE14KzDJ0eqQLw1/4TqX0M72gKqIcqRNEo1jaTPRDPw
mLggOg22M1JHY+PuJej9Ny9lstTzYMxenDqCEEqPr861CrYaICMHYlN+GibaQ7ja
Sa+M4CjW/knDQP0dFcwB9WZBfKTneIf3dHn7GlJUI5IOINOC/H0OrUbt5VZJpVGx
oqsnIrcTFP/pOsVT911PKo9f4dtfTzoVwhDTFczzmtAI01fHSZFojzZ/1uv4/APB
ngX76BKfWUZYx42+5veSzttwp38ukgyKX3n0ALzbFiru5+QxZfP+93WijD5We3m8
XmDqdzdMmOl18f89fOsBZ4opeIfPElaNDI0VS7Qi7f/dMf0bHKIvREAOPORBWmci
I6Nkia7qMjGYXD0UjUcq9zmiNVdkx+qyZX7EdxW2CV/xSGEsTxYj+eSW5tu+ILXQ
jFbp26YiM/tPMoUqnDVfbWGzj7LHlZphDllYK4Aja5Z+b/Xe3VMoIJZ93iT4/xSt
TQmwwrV5uZps4zw4Wx0kLzbYgXkntd4F5UoEkRrgYqqd/WPUxOMPNZ1e6ymmSRiL
U7JjQW3VPkfgPH0AmUjZOA1ttPJ/165GkmgQpA1UhiM17zE9G23wVlMb9XVfbpu2
EbRejA1E3ag35ppsyVzs2NpWj5z+4QT6wEhYvB6m1EHwT4bg2FYgPrzoba0faNqN
Pub2VE/LQZ02LUHB6Bb6t9yXnwRTXsxpMDeDKEcGCItU8k8RPzgihZ6qysle5O1Y
FsIW/my4G7eX4HKgadO/2i3TA3wsgn2R0AqTjAdSm9TH5l0cA3dQjnfiXMVysIOV
PPn1FvNZjgSozQUpvxzvCUeiU08p3ttim9F9lOWWkFp4jMBFBCmQWFowqyVF6XX5
CeLRxj3MLXp93bMkvsywZFx5fyJ4yq0ak172Y/G2ATNn0/qdHewhL7O3FAHw1VUy
gBvAlTwj6KAre/mfYfbMObO3DSYZXHNR69Qrd49OEAwmYReurjkUbAVsplsE63Ti
d2bPiy7bRAs0O45JPEzlnG3fwQBwg6QeKVGEecEEbqAIul7wZcWS/KbJngA9sfOT
tK5mW3NAw04bEnC9Zh1rfFE26cra9n0Tl2rmF365JH+NoDeUg9ageTX+9Eiv3LaD
Q2CsqGyZroMnjyPcK1K2rT0gO3iqwNmzAc4XQbpXw9wg9XIlkYTtjh3dT1bRzE9J
NmL0NZXv/Ryj+6SDEQbDug3XTmmepzg4+aHas6S3IUi0+MJd1wzzHT1kFMfkOI6i
0NwWxUIjjO/pwutQ+bnzDWlsFZZhiPGtvutbzcgf+fDTf2UgGdPccdvPvdFCo2B4
t2uj4Q3+aFmD9p9lr7TDOkCUVMTTDws4sirgQh79fYN6Qv6XJ0B7P35uepSwVdlm
iw9K7349kBlC8fXguf7VijkGx0FEyrOqYDqP7qCpJF6ZHpiHw8XulkchlATWrP9l
loXm8RZfKJqt8LJIiN9XJ6pAS3Qb1mOdY6kPvN4ChBF2rxEtQvC81O8WfXYCpvlK
3WIY/50qON7FQUhxVG1ES6H7pYEYdJR4bgx4czhwg1OWQbdCE4Yj4dqJ5rZlr5gw
spRIHNnwBP2fsNiBjbl5n1+SKX2ODhi8oIvzSKUoXsgNRfG3P9EJ/1JmMJKEKFut
AhOR1VSj512vAlzVehECmjWB0GYeHabjP26vpguw0rvTU5ZNKOa6dJu4nDtCIe9V
cOkgu02xlN7BDMvNbvgwD2+OKvNh8MDgqfZThFBjk2/iykvxh49sg/AsXzJ8zXY6
QcnNaIUgfhPO7taffeBH84ui0/V8i0R4a9NNFlRLj+cIlB4gVw/CAIM3nyMsfjD8
NT50xNjnPuY6bByYwnQbL6HD8kY51YQdOY7ybRqfmtYRt7VwAMjcD+YhMDivO2Eb
lGy3hMP1At1+ieU+freay0bf1F9xAwPP25U3rVgTV9XhmV8RJjGXzkaiPe+Zm/+d
0mKEkrBaw1nkkay64mUCxkHWULvF4BKb8U04SnhmDpuAF6FaMTuAssGQB1R5Zgcj
Lnln6Tn8tV6aofnuUIv2ve6gZxdfFMbnvKZe1f1hK8NezmuKzfIt/Ni1Q43a01Ke
oLA4GhgbpY63SsIV45DVy4eMgVrw3z5QA/UEIHrMBm/Wz0AbrUNty2I+DhY17DMm
5O3G0GlqWHGg5FUma5EM/TVGmWAIr9HVN24D2SWdrxCpyzTNTXbLLdNnYPtOLi3s
/yOwHgkLHmaZtviybqZp+JhFJ1OnlL2jEq2ism1YgWR4SEXpYtnGt5UYXrSqvWGQ
CDxMB/2Usz685PZJeShgFPwxXdpsPBBhycR76hazDfPKfeLQuhdefV4hYlhsjI4W
h1kBC+WULo3xBSF4FkyjrJ1fGheFPrm+nnPU/g80LdfBdmFkV4qIFp+8IEWjH1vh
7qgKk1KfYxBJn7z92WV7GQ5RuKAFjM10h7i/qWcHef+cuc2PZuSVhDUkJ4p872bC
51byhV0fzbWO7qardiKvPJrJm4PjtpHe5e/zs2Wo9q2Xti+Hcl9oA0EhY/nvUyS5
SFqOh9/d6pyxo1PxfmGyCAs+rCuk/x9YgMB3EPeBtgnQwBycl4isY+zBtwYUAxqk
RSC+VdLt8+bZPz10kP8/fuIPcZGxg/Z6cxMz/6wx8n47ZO8WSSR1m/EzWwf0KsLo
7RyDgxgfWFwNHNsalVgtbifsZlUESr/7r7+OKePfbnk6jiZ6iwTf62AprQQXESPa
XDFXjFMj29S5DORJ5z4hle7g/2agnSgIz7t8UMTX4Ug39YfGVJhI/ZMF3ocpjZdM
1aEYR3FiWJNUVpUapKstOXb/0TgcPgdisrV5eQY66Kdpa9fC5vQ5FTn/vleEXKFm
NbIH3sLR1/S4Q+w/sRxzgb+abMyEeieLyNikVzlLQHY73inrcn8r5hifNVGFvEyq
j02I9o//rLe/CCy3Xubsl0OgqsjjnH474slLAwmStfsuUfLw9wiqTKsgQCu95TQp
2Pc1zkNz75+zqlOwgoJFn1NZ6QkJA0KY1G/OcE0jHV+bWUnzFSXZyeiKBFTZB0vQ
QzKAoGy6BnHIaP5Vy+/+fIZWY13ZU2hCWn0LM3E0RVj2FIRZKcXoeaKL/5hQ+r7Y
0m1yxEzcE4POXsiECMi+/dVvlmbYu2agqJsqxqME5kXgBMNhnw+4ZLWht6BwysHQ
NPmPE2eF7lL5EeChJ1i8MwWPLbWnUWnhzrB17JV4hgrkGGAuu16Wwhx7idKiTqoE
F+cCh4lXhWLjrey/wnIm6Bujnbgh4qL6QIQ0fmuBfKhSZC9U5uboaxujo2AL6JKr
vb6y8hJRQX2oKwSprRMdl5FYRtaEMnSe8BmqIRX/dWY5G4CIgADtU58TJbuLkFdI
GqBsRDEEJKS5P20gSuGIlvcV0Rb52Mc/naADA4zchveMscSfW0DbzUuObYVRjKPy
srYvZQ+p6aWCfDoVthRER62T8AyZdFXFdo5TAOHyjhgYJ5XKkkbPc6udurccl94N
Ch6xX71FtWWwiizjkBYSiZnQOGWsvt4rfaxrDA3ti+gt/Qx3VjBJQPu/q8MhuQxC
XBVNa/koUPiPco2GDE6Bg/LTFn8KsWhrvYz2Iu5V2dHlZGrZhKdseF5tvFOHfF8c
MJojLDa+Gc/9qBVtX5dM5ENmgpAL5CO6hXstAjFLKPJc4tM2Tfs2GIk4/uHJnEDz
RFQ8k+18bdpC1M23NWW9uOCs6hWz8hIqZ26kIliN6D1mrkIh6GI0WnfJho8tgeud
zRqAQ/2IVGO2xtuwBmgSBuoRqYEiC0wNTyWnao7s4Lgd4IRnTOBsvzxM4h8X+ipj
yfHZZ0+q3/LhvR82S7zvB2OQpg3A6ltyQWfDE/Qvyz7dN8H27pBU9Df2aZBwkiiF
zBT1wV5gjRtkf6HSAd0I/zxVim+D46pEG+7CAbg5hNmJiIYxUBJXaev05OhDVSVR
R/dlmarJRJGMP1MKyMPmJYpYR1Ad/PtIM01H1W+FRWuUYMS6Vhzq0Fg+zhYNFvWv
T1fAUFF4nCIOPnkAb4Du/Qc1cQlrWcSAxWn+QfkNR5B3kOf8I+m5Co1XcWTMuVSC
PwhxHAz2vGeRmNPi8kMHu5FESEJ4j+IREGQ5uThpBu/MlPM0ktV5oX/lewatYjvI
6dLGPp7O/kgrmnQSBczFEqE4nUpuliizFlZZ9DCDdisX9biIuOZ1IyI5zKVDasuT
0+5PsZuqYr8+hvjB2fWLvcYTPcGVo4Qmv5cdMw1Dj+PVx3ppWIRmYW3PppXbOeUM
hXA1h5dcWA5LVf/RWfitvSs2RL9TzsgN398s8EC3OKz/Do+WYAPhNIIvaWLt/i12
heNSucXuEP9D/zOO4uP97p9LZKBzJb/4HoIMqcxNcGTCaLY2SicHAvQPPl67W8CE
ZgrZ+hXVNK1reJIvNLZ6yKWIMSOnscNgcI7jnOLPtJVqMLY9j5xkP0fPiPcfP3uR
qox5LpTM38Co6eJIagMBCCPfh8Tfdf6BFReL15CSD9T66eYcIApWmSxnD24Mgrco
GNn84fp8lflex2osLv06+wV1HTDUWoEhAvJ1fdfFEJQAOujSM9ISbL10gSNWwOKz
jkbG4jR7qUU17HRKsRlEbkwByD17VxYyI/57Cq/zK5QY8rAyFsKW5qySwqHgh/Hu
b4EH2VoUV49XjKtgfkf1BTrLOYgHGSi1c6w8aB/2QFa5IhNtuQR+BU65E3YJuJAt
+ZkZCERFpgQKbXn6HLf9UrSNKbCF8exFXfjX8N2NN9yhrpvDkHKGZK62gt2mheV/
RGkuvLlA3tRLEwEIT3DXtmvUhLFN0oyMCplCdlB0PmBR98KlhUjQJg8ThPs8S630
j2SnsDx8aShpVeY6RuIlurFHZLjF+Ij8X3YN70oFcpRDmfU7lVsG2x2CfV6ZpqQ1
4bRrlGpownXgTQAxqy3UG5fnkempbRq+/YJkKWpgmOJNuD0tJsTUV1EgCAhrf0YT
WmsUaJ+XSaLcwVtB0wQuK83nneXFcbxTjZ9+VbEolQLuFwPTnpUSoe0qA05GCwj+
zcqlFXbSLDcopLp8MQDNJ+3AXeRA01hXqxnErGkD09Pdzx3xeOQY4PfEbicbbD5U
l4C6pcYeL2LbqUm8JkaH83J4x/0KIp6ixaE8f9ivqu3yjGaRxnmyZxF2ThGIu0cj
ayeUA8S95R/jNhiGfmeR7ghBjwcWIik+ud0ZhDSE7WoqBS1xgb4zsUbhwM3KORRw
bFHv7Vw9aHxqkklJsICz+SO4cFJXTIK8oulMEs2MrlBhbDMfQ1a/7PyblYiSZv+E
xlyHyUJ48U+YaEBDvgEHPDsfEWlPPdib+eZebwuBSgYLnxZqEo7x4QTjxCSxfxyT
S6uaUxu0blJuHFP1rUdE0IV0mv2qKhEzXnWjme92iY/8ljC4N1pi1mcf9iV9SNw8
HT2RA+c6Isoms4R0VhtY7eKqq/H9APUkv3CZnZY6cDU3plsafxN3RsSVpZX/zdJI
2SaHHX0yfbeAvRQQTn4DpbivwK9xpusfmpvdH/xIAnqOgSsTSjlOyCZp7ca9I3rL
pelmrr8nTwW2rziThuhHXJU3gAxrojiY+zVCxDD5IV0JrRUdYCN+ZAdU9ti0C7bw
p5KBMYALWXcOWa8YkhtR3hnCJSyQR+fDPi1Z9tGEnampZt95irWTHyFmAOOMcWKX
JkD1DMPZY5fa87z/m9U9psKbrR3r/XGfcBRB1+Fm8bWOG6DbzLxLgQiFSNwduSsh
esZr6rjEQpsa6MwC+ORQbwWJpyK4k9B5VCf0FRnCNq+RepOV6+PwtZTy/1cOTiRP
aXE5TgC1cFcjspJACmJKkR7Srq/cLMFljEggbK82e2503xY41/EYfxwCehKMk9fP
FZmsMRUQ6fbC/y4fJyZc1rXcGy9ZIClhs5cJ7I3r1URhV20rctu1eI6k+4BUOdDl
jcBmNbVLaR96DVdkFMVZp5g9WzgcxGrQIedymbSDQJG+0CS8U/hFrjiziUXgFX7s
Sdjot6M5j7pILJZs0Y41EO9UjAn+IfHCtVMYblRFafxIcCClhizdUjM+HKm87pmC
eTuzkznC8fBcTLHvFIzNR0+6z1XQKMXTx3dTlg2UxZoEXS+FF9tE1krYjUdlq6la
dQoXn9o2xP1PQcjXXu1gwNo76VE/dTKRIEx4sgOysHg44BWUFaVq09WRpi8ZBBUZ
P+yW6wgUQUSTPhtk6A8Exm8Xn7REmxjpCjSnjxyWFqYVQppepD7FxT+uPChci+M2
B2MYi6tGhSS1oE2U9FW9RaDOLiT0HARjC9QpzQoHXFifAls7as2wnxu1fTsGraZM
XJXP0s+55rkidRubot5Pc1pV2GQINrFDUarAb0211e2i5BTmBkVgUIfW+6MtxcSl
l51ro2A6UwUkDxj+u6SqDtc545xqv+3yQ+NpUZNzNBtriNPpqCprm4yPEq7sVnGR
R7e3ku+nbeF2WhxkSXh5y2szubi6QLyXXfhqwY6KEc+JWe6jX2t6C4YZcIS+LIVJ
23miq1ckXjHMqXaeGhG1ohIj+nm088yWaX8vLvzyijgd78q5VxBEc0psQk3t5Xis
3Y4kHip1VZt2mViD1rXn5y+W8jRcrhawHysEfkJ3oWLPMSdir2sTxns2jlzrp/Mm
G579nYVdTVNNj3d8ukuMuRZH6yoa0BBk08PYW9oPF/v+N/LVLhxUSufZF3f4zqst
bvhAjhuk7OggdOlUJ3DrkMoiHxIA4brs/axaviAJfYQe9Q9oSrtlJL2I+dCTSMYA
uB3G2X4NzRSxn5KPrFx9cSVDFtF7DR6rWLuM8uSm9H2wld9TObpNHdHxBaMxr9S6
oZ4KVeqiXKYaRUhpfpXb1PzIR2u9TQza6g3FvoHfXedW7DiCIV6sf/cG+AzQ5qMK
KzRL7rwTGDbWXs5KbqhKWFL9VkYFDmQKIHLYg0C7UGSrMqYl0hnCee+mRR4Ezx4D
JM3ZTaRAsh2iJZkw1bsfWoUDdjiPSjd8hEzc3kSvyG0EyqBb7zMy1FdsoXIjaNn9
CSZ3bJFPD8axloizSrxEJX4yXKAPNm5PoGYU6NS7L54xjAe+aACxtuahF+9kNgsx
NOVh9jTYUD8ws9HissvvphzRZ6dNBfPnea2u5GUkbnns6YneYH9UaXUfB3MzEFal
W/kvQbI/yJVW/0r32JjP7wqF64MgO7kZzOcPAGJnik2ddxuZJx4/MiVYNdQOrfsj
THRuEtokd9VpR8812e1W66DVFiNrQdo6ErUEBU3bouvJrUizsEAvxHi/ikEWEacv
UIM/mCd9LEzIqFetWlfewalLQAxEfBM54iEp958yRKZyodPgiPta109cOpP0tuoP
/p6CPPF7iLaWwiqSQ5GRMu7QwdDdReADgpMCTl9bMmpKQj7bcRAp6ZSLz7zv/qHS
BIifQFD3CLUGiyMuzmdITZ9xQ9Y07soT5AtMvGaCmokN3NNm30RSjEUeWE9hcxp5
RWp9Bi706OSDU/Ln0+kEPPz338AYDxzUH3ANCQ12IdFipS/RYXY151mq89VHFNK3
0rM4h3PZ1o1TmuYMfO77BY/3OcEOzX5B0rDfRRc0klBgdZw32L8Cbp5xfAktayDF
s/wxjdwR8/8+SlVro3jsn3wOmAQZp0wCO7RO3P6uYmPb73v0wPlF1Ql3xQQiwdaU
u4S+LlyaD7QBVSEo7p8sfmsHuhT8G9INcCHcZM7W1JUAMFIeSzDhINBTtq27ZwP7
XZh+5WTyCvvyswDHsnrZvHqauELudwTqTrpjAo0N3z9tFsehPEgNlH+a5CK/SY6p
Krrkw2sFDZf1OKovNsJoA9IjK3jcWvTS5PJizGupkc0UpRVxeemIgiQSsgyT7u2+
IYDYFCcn+56rlK2yKWC4lVFXs1Hsang+uEuxKzaZSYPAqBA6fyUjg8GFOVanDgWc
PAR6LOK6TpARlh2ADPDSuqDO9wi1QGunQQGomnbF9oOcFwD0jTvnX0FvUGyBZYPC
nKWqrfCjM4U5aD4ADKL8L+3mBsgUDsE8dddk28d5YDAxAVW+YtrUz5Rc1iA7C9Xa
nhU1kk6RmbjEUvh+WtCgC96hF9/ou8TttaGpAYXROPLZqzQWkco7FbjoM52F1Y/J
doywHb8Rbluq+C3V+MaBbvK+xVkoSd8Lfz44sKoF1oEFEn4i2/Q/wEnK9429RZBP
AjmfDCpYt8hIIQAK73ZmvxjErQboNH++j0P3agdZWtNIFhEAsrOIX4lIRMKKWgBO
UGxYUUqFvfAc2gG8/Vn/fMogo2tkhHttAADbo70fR2LJErTjUK9Z9MIPd3qZK6EX
bY/qOcLxtUE6ZQLaZmpnvBqngqv04I+S7PCuIPK9TTWUQr+uv8v1aHkXYV1UE2lb
dgEBun//VRdRyQnHKvchHJ1i6xCDkRRN6AQhv5J6qp+rT0Bw7nasxR0HBhlgjF45
0gdqVmuGC2EeGbS3mf+G71S8PGuR+zsZRi+xHwmXVJN0wQuqJCKetF8tgMNeq+GB
kw5eAvNvvCtxvSAwkjfwEI3zgX+dR02q52dljV2VT+t5GGAw7j90YCUOZxBdgxuv
3gwWAouaMeEBKZ8jY054gHR0V2+25V//UYYrQWkUOBgbx8AiUIg73c+p/C3tyV+L
xgDNzoU7maeFeJuwF+t1raVOKXtKz3BcDBaqxnG2brnviLnDSqeX2pCjql3wM+Es
WRzBP2XAqJwFGSD34yk+0kxGu8ade+kzuWUH1prAxqzOhhM4u3Zi0CSD6/OIF9kA
kzkjWYQC+4XQEumaYsMfpBY3TRYnAntNWUbZBt44uXuP5AtH+3w6BEmhF6THUtrc
+li6rXPr8W3E0PpO2y3rdlEO6IOWkK/RX9gO3n8f9bv0Cfy5/1mMEaeuXlfP9KPo
lNjI4kjswc2I9unaUOdtrjScIJLN3eouc1hFgMrT4ryz8KG6CDqf4RGJpAiuCb/+
N5oHcvC1MGByD+xBt9u/F1nQ6yL7qLI4psjpOjEPz+Kr7FmlRHvFSb14exiOiorB
5VS+3MbFoOcFU2orFD+G1NfNLmZE2mnmKkqlg/jW8Rq+BF/Ob+Q14muppcapmyuI
pqCyGRYY1b3a1twVK9urlLCikHOACVgA+EgrvDZeP4vGMjEVXD+73Gedbyftgp3o
MUajlG9kaaB2aoymMWA/wDUB7v97CYnk+NB6LXbxQ9hKiTVNlJfW0avh62mwRtYq
S7OlfwzYreJxfqpu+q2oaZl23DJ3diz2PPXRTSMToe98OCdzh3IssjjRAPYqQVoB
TTU+YGKrVM8uv32I3bTdphNOZ65UzzQo8zD7ZMWUek40M/tI4gisxB69u6MhAkz/
3P+kgnru233tppith0YmGjM6KDlNbqiIU2FPf3UD32G4MWA38nZF3V0SqT/uV7Uo
zYM5B0qA5JsHzgrCnrRGDUkzjc5NRSjk/hkoCRhz7fkQpWoruTOLYlDzZfxb7UIb
1wbB0sL9qdGTpbfixFA+xJPNETFxJII2dwBvgLqCbL1WJpzb5sYJsD3ihYn3y0H1
qgIv29l5oof2uGnA9VeoqkdItafp6q7I0dqCgKVdSKkIufTOeKqs/KpfVgQlfiEx
Jdz4dxyV85AWbZeT7eWsexMneKX5+29LlQaSiYFTXGg2hT8XS+UcqVpJykwqlbJ/
ha16dynwAj7JyW9+TkP4z7VHkvXehBAYpjDfv2aCzym7SjQLzIf0nk/iX2ocfJBn
zVJhr/hpuKv1DJ4BmK8Oil0XgIm+iig+1B5lkjz2Cd1sUebvXKqsCKAbI2KReKx7
LQl44rP1TyH50MCxGneIWNdRRHXXfAHmLqzUrk1sTrjT4eK9Jh5Of5XGEIsHloKh
RWwxXRAfjXXbfudkVbdZBhL9GDGl5/FtJ9cxlIVjjsahE/aqAvWxTrdWiu9Q/la/
zSdHnlQC05CQDuV6MPpB8VF52Vo11tp5iITt68a00El/vYRqTnZg/w53zMxDeM5N
AioQ7avGABj1MdS/RMajkfQp4te4wBBw4vv6UKXoIXNWp4sJtQMp1U6WWPD+nAxk
vSlfsIf5YNmHonbVTbR6tsyK5Isf+QcEuh7IsiZpqhLXD1ndI3wDYSaii2DNzmfW
Ce4sJQc6/plCylTZPLGI0ju0KjobH06UC6DVQIDzyNeZGFjjCmtOhjxoHNa3Z2R8
O3sV4t74CAmoabD9stgSm7bn0BO2uJFFvlkJaflgja6VWpysWsk9FudqS+ZYi6j8
v794ZoZlv/k9WoLdpobGtPBdu1XiE5Dyw/E3DGPHt+JDQNmeeJmn87ZXUm1On2T7
I5tzpvteITafO9PxMSj+oIVGQ8JU0QcUVvUFrEq8vi1L4zZuXwRgn5Ra1dvvbgyL
Q6Ov8Mws0P/hNnr072MM0bpgO55wF/de2uzWgtasKBvuQmp51o8PPzqgyLhiAtdC
klECzaJSEiNANWgw7qrF8UJLxxNVfh0LX9Kn/fvw+zjI7kcKLFS2HxFBLKg7AH/y
Oh2ajIwIgYdN9f8lXx9c+HRiiA83jONeQhS6oo8uMHY7HZTqC3kA+xKfWx6NsXsC
DxlzAlAk5LtQuCeBeMkC5Ekx5iEn+atAQ88Ze4SyowjTERa+t1qrRskic2XQg3Kb
+sYrZbhI1PFLeWoUh3gdxpX1R4I+b+PWo0DBDy5qpZ8IqzqJw9vTZ2tmzq2pwqLy
dIGxZhB9wZA/vAUUW73Y+nZj6J5FlzRiYaXcEQlYqBlIisw7paH3KtJWnjB3HWvV
v+/aW3+ZubYZ0qRmKMHjt0rIVYSZ957i1G0JBnmcUs7kB3a18+xZV7lCeqTFpbhL
p5s92t6hvNtGgnKbaEMttrLSJp9G7XYxHaNjAO6Bw3/t5T528BiGmJKXlUW+Emwk
wX31UHmxfVa7hU3wRUNhh5m1ylKTLEw53FYax3+dKpzwodunwAoWqkSRNMPVh7+q
oPiXHMGMHPg5QatQTXHK9Xe45GUdyAZeJ10LuuzlQ3SdFCPPf+m/lCXXwJvHHZFt
NI0bgno/09+vvLzMnyvY2Wen2h0DYOYbIEAH8fhiLw4Ri1CpCfqVgpEWxgI8vQPD
9mawtbvi1YmXEfgkkBMB+ImJ84spaSQncedNZfYSQwNyociQlmc5CAO9KEoon+KA
S51dmy7SMi6t1LnMDreq0qowj37miE+eFE+L8dgOtNy5j8HQxdHVzkfh4JVYVyd8
iu99c4YYHZOUK1EVzXJqL5oRbeyoEC8hcNzZ8R/VYI91Cxh4FvCXJacYieBzX3DP
1LLhFLEKPn30JAMD1vBefpVtgP34UlZzIbx4AOcRliWKcZZQD0+mWhmruT5WWMGQ
KXIiTBLTL+KziMaGIY7WFqslZBwahglmhEFzuZr2RMTUipHYTd6SeO2TJ0vJOz0I
hZh2uHbycpxG0QoBgOU+4PCWmD3NCGIoZRlsY8x0c9Gh81JY4k4k2/iT5WMCy4vN
t3lABIg4DY8Dz9t289jbRrq96Jz20IB3f0oiViZ9dwky3eBbK2PjGbtwxcF11QKt
lwfdMXYdnLpKUIyjlrCoeSNNDX+b9gOhOHGDrsly13d+3fWZ4uOLnAC7k5Akn0km
RUY5L1b2MWXWzel5ZN+pV7VWZl4cuNU9VePZlnLblV6+a8nOAn2WcwOIf12yKGTl
TD6j6vXFqW1raANvS2GQKbE2stAW28sPLQSj7CULR9ZNqAy/UfXkY2iuZjI0koMx
BFj2UrBrQxoXFZlfUx54mbS3U2E3jVhXXZDf1DLUn161eGe7lJTaMzq3OPqX7PTJ
8s18G4eIb03yQYd83n22qLztdLSssoXFBupu+lomExSG1c9uRlgpureToTz5LD9k
ubnhrO0PTcPsJ29/7uE+ehswX3y2GfP0kMNK7lxDVp/FzH9tI6WbeXy3s0qsYnwb
frrz3xar6PMwjpXto7SzcVAnt1RJWge9N2LXGM6l0TEZ4tPC/RgtWsPMqdO8lGx7
tHumY/JrJlyEG9Aqj17xP+dBXZo5QM1YvBYP2cWkARkAg+BDrGzXRqs0YkJ/d1cR
71NMHp8ntdRQVh4r4LuOUbMhJXQcwjyeh78zrheHWy2tEtIuUxidPBFtsH1HT7ur
Hn+9Xbh4kUpPpW0YNwPnbzhve+s+bZueZ+gYH5B3cx5qlZoiGD3hvEbl41hFZbyM
FhlaoQBCOY9AGDXhHZmeQDtLKwYGCP1V+RBisc0svjnSlVgzYJWUHgRYZMP/iaVI
CWuxCR+cI/B280/mxQzZydg3nvDUapPi8QAf2FNjfZD3TXJhtViK5sljATjvtjQE
WeAKizxDh1FDVR9I0PD1auq7Pvp3THlgr/6UwJgz5auwu6W0xksd3gGagDfkhcgg
uCdjeAEUCuk9Ph2ffmOnkGKmx7L+gfBNYUB602iELC0AvxkYLigG4R2EA9gTNWox
/K5Y7pYKWKmQhbRO/r4nNM+4Q9i7klMJkTrEPO2+Ls4otRsITwpu8UsF0uKEhUDc
u4QEAKRx8q//MO5kaOglSfNZgKeLTP/iKMhgkkfMqwrW8mixkKIlLZ6kOEvSPlBT
BdmRcrPV6vl2p8aiivhIWNpKLRERdeFVVzIOsoQc/cTqszqYxCcJv+dflu1wmrSU
fwnLewlt+C+sSZ0up+0PKNirCSuRrH2F/j8h7if7edeD2KEcrGIw+w8Uzcgr242i
PsPHUdjdU4kmC19By2VY0IePjvEj0Syn2H8w8owp48PVK9M2Nnkn0MmoR1m6i3yb
4mU66UHxj7oD34AELFLtIsHOxgm87B+Pu+6XAED4PgVZcMtCLdnGgx06woKxhs5R
xVR/SZaeiSp0LMdOoUqilvRwQWZj9Gfgyjuxe6Quc5PNscoW9Fz87rkzx5pvJwoe
LeopnUooF5jPdIn8A6LEa5qC3ErBaJI5o+4c9MpzJ5MvaCSHHA+QTp68UMSWGU3u
pTGCky2tcNlRvAxeJ6Rp+y2EdJ1CKBuyncsxrNTJAYtryVBhUohIGyKX8SHe+E5G
pxZAD8sKlOzHfahKPElNk7KLrtQ7b5f4RZQoQkTV+cW7ZPG79Sk7+3Ekhvd9ZLET
XiSit9tAd1y7fG+CiqBTgQWYhn4Dbca5HAire7Qc+nEJHdrUrBnu76JZk9m/yTLP
213NrlVbXAHT0y4hbZxFgvZm97PGP/QAeNxO6HIKDAMy9sr8OmrEdeFAf7IBBpT1
sHVg3njffZYf8neSPYf4qoTlRXsQmacQj67/vhqJSb1yHoXsfVl3wzkTUe+25iQe
wFFDbvUnuFf1TZObcG3Hf2pCOIt5x42aZ3oFHHQrUSVdtykyr+htIBowgAmbnRP5
0DbEs/d4D8uK7WG+mmciGrBaeYp4P9zYjc0IXz6AULV1pgEEFjiRNEmX3j4p7Mdy
HMwAJFFKNdPf3nk7Zr6twwghIo87VBfp5TkcgVJhdzLyOAszbvLg+eiU9fNBxnNN
oadvmPZUGohdw1Hwa8eAL2egeNWc9+vTE6uimKdIr3VsCBLkaOGs98m9ONNkt6TN
8Q3qYOfYX1zbwRFSbXCmyw9lBYFFCO4OGcq70z3ldyQZq0UPidfI2cJcmzspl3ZO
8f0pekaK1y384knSneBD5cC1Ghm0kJ2gnDT27PBL357NeeBWMlLEuhQajWYjvkXr
Dplgiy0iRPwl3i3FOV06OzUmJP5qWwJa4UEXyJj/mp+G/Wta24twjIzOshUmP6Xm
fnFzwG9S6V8HSzTL/P+U4Zs/7EmWrka0V+Yt3KuDO8CT8bc7GABF9HlncC45J0RA
7N0o+ehc1aoTPdqpsRbWmVu+WdAhcgh7/1nMf4TK524SaIHrs5MI9dGj8EPJIjpc
9mB7cRo7eMl9xJAE7wxdT/e02W7uCSJgdgQQjMIAffpZ3d6a/ZInNFyMO4LU/e+/
yVxTRqRmvtEpSxUUhaY2aUasYWNFGA0HK1ZLloQH294S6nTif0p3UX9duNXX+RVr
WTfY4jdTYymoRmXVWXKuFVov9HKqUJTEBm4AzYsBiHDqONp8I8T+mU189rmA8Q6Y
yaku+ViF1dkc79/cX9zdX4zYj0RNerKRb1mMavTRarc25TQHZeu8bHX7ThuGSTEp
ovD2SA8UzJT3THo3LSLZEqy5Qr9tNS/3EjLIzYJ2MUAhf2R0qF74XMy8f9DpScvA
50G1yxnNfjpsxvGMAlwsTe8NVAMiao5bTE+1Db9F5D9IpjQ2eMtktlkepyROSOOs
EsxMurWPgkJB9Ycb86poX9erm1cUhJCKcImGgLdF8YHfUHnHnhRe0fNwdVmZO+/B
Mfmbh/e5pCbJ+bg4i3lnvb4KeJQWWu36hY+u1gjOeV77QKaUdCAd36EQpKYBpcNJ
If7s/K4puiDXj2X86fUlvUAhrPXuqt5pErQqnRz5NQGznDoyqeqpl9zAqlenvLY+
YEguBj3h6o8XGqDSvUPhOOeamQuOdwfod9tME3FwqhW5q1zqquAo0IpcG/e1ZVRk
AlO13sCbos/qIAwgPyfX86ffmdMNrexeOO9CGcpbSqBvJMj43Du4U0LQHp2ZpPTV
NutygTEPLMmqnW0qnz1wnLW2+4XvrsOlfxF4YLOKTvUeqFzHnQXBAspsrrzB6Btb
Jv+dYLOBZYWxjIfzxdiEHampnCPiNiwIaY8NSfqzrmXx4uczUJFqamwmGHE3m2lq
f7W4g8bUeEDzH03V9aH7ISMZmDou5pT9mmnYIKVSYmXEx7csIOQspAg6ghYd5wwV
8B5tU3gDOHmA3b77oqX7Jc0CUnFk34xcmDdjLPHh0gzXG5AGmplFDB5M6EyN3Y2J
zPfupQRfFGpCPFhx8U7EvXwtLgQvPT8jgDqgB89L4AHAm5IXOmne16UM70qF5E4u
2DX4zUA1FYk5Wt7yfwKFuQSg8lnYUiElEtHAamKN8sBiTXNzZxZGxaVHkPv8oraN
0MaKvNV0LlsbaIH1RpBTy7C4CbiufdiWLDwARdCazP8SKJ2xD3WaFJTlFAnhXLIl
QZHywFD4Hdmop599D+GUIaxHYkfaKK0lddQuJsIkUN0pIUl691PuOAzCiqdKC9cz
77oIHP8J608U/5dn3lT7lXDtJ4HX9/yMGgqIY4i13p0SCZ2CqGVxBsbZZRjENPXJ
B3/yNGI6pYi6oAZeTsFVBIem7MvyPK8thOsMweiBFauisINY4DW3NMZaP6M9XkMM
B1Op1ejEqL6Zj+DPW9ehG6D0kjbmwCit3irtX6u63Dv4a6NlfffMen8NbPopO1KN
xSDDaqJRWCDw/FQLfwh4jZ416SBNjVwrDo+KEL3V+eiNhI0oYQxr9Bz4tPHfBVIK
yw3Y4AY7f15OwsKz/drP2NA1Uuo5tvUxPo1Kvk+XZ0HUuPk+JEjxyeOAcG/LR27O
oeiI1Va77QTAniCkpmqmIYQ4RJyTu/Awp2hmYwdwAO/ciVmhzMJvIT/rzGT5Z2hd
CmEBRyOEiW/7SeHkyXgtg7+TriCgx1YJk6HAP48Hi/X33ZBDwERvwjlIwk9yUYRA
vRNa6oF9YobjtMGlXI5svsjObtbWwQfQBO9LgZ3HDsFQXVdXqB+osq1XBoBXOhXY
BySy6+QwVljmuxUYNiz9GChLWeLFB/O5yHnrHaFWjJR3qH8wMX/+ka6c2GIJvZld
5ToDMBJ8dyQegau4igvQFZUMAtxs2/B1zU2cVY9KvJV05KMFqzZx2jaJa+9pOXa3
q1yQRQPTQszQOxC52K1jW7iHGHhfHgiZJbEFwJ3SEJZHCS2xQtnqZF3G9WjM6Lk8
dQF5pfENY4DQIkONBAYpb8+lgWLlYZ3UeoudQU6cveRMImO1DD0k8qgfNGZidQK1
WMXyj6bHbEZLx2oLg33pUZo92DG997FFMIWhpMAtG6vhmj9+0Qq9sxusGw/zbjj/
EBtPu+6/XrEGULt1KkesbDdg7kyF4gHRxQaXi6mqf/jiNmVhbLliOgdhB6eHdaYD
Fh0iMCMMRf1Th+j3s3qW5vmpT5iWUY25f7cDNtwatKhz5B0tCjDTXWfMHZtq7kdc
Ax/MA/whNTLbsg/kd+BjupfQH6n7z5Hu+Wxk9MYAehSa+/dxjtNnZDKkTNf6o5aB
7ZXtnPLJNdqk39myqQnDt6buvw+vZQtrKOG64L+oH2HSicERmq/4wo/VBZXQHTuO
0YF5/6c/GELg4si9iXV6kcHg5yZc8npEL8eNBQ2SX+jn0nw2gSu3HXFNvD3lUU1k
RkEto0l05FHtETHDMspCuw5rrIlABJpWfkRPwicG7yoC9Jps7HOJGTvoWJCAhF7T
4VOOg5Cy0S84pILzjDY/fjZUM8MUT1AHUGUKJho2P2UZHC7rkYf/4Jr0pp8S82dd
f0aiPMrg4Yn7IwNCTO/dfZcha0madPNAcLzzSb66cHnFUu/qXqRLsVZYVZ0VGu3D
MP/PW1nLeGLRSYlHsx+Sg4X5924azQtS1O2zMRIGL2TIuBS6NLB2EJdXHV7YkBjG
vrWbydeN0fXLu2FqCz3ask+9dK/3ulkxZFkjCQfMDXJ+ocp6LvuaI0ucLWP1qj99
rYYly49rYGpIRuzTw0gf61ms3XtOZHp2tcbp33PWjvGLkSxJp+jGu2BAJQ2Rt0L+
klTzXO8Yr2kOEhJrikAdLZa9tY/5yCLiOCZukXeKCN3HdyIrJ8qCXxpCpyr+6K4S
j/sqpRmDoozV0YqpTHp+E/GLcg21zJUky4onoE4VRc/KxSiDEK7s7pKUUsxhDJJ/
L7rRwtK7jTTfVzurlHhd1QF9fhqTvbU7TcPPvvEWXeqoGQyZ1Peh27KNk3azNobW
r4qoOLVDULYpRn7io+Dz3tJjq6gwZLxuoNWJIb1qH8rKu3Y0L6g0DjZnVWWW/ecd
ENJiBsKqqg+/MvsfFFzJCX0GzBwwb7QSrZhurPKU8z699zRv68lE17ktqsxjgDtK
B2co4B+WeenKO7GSspN2w5yPzMviQNWOtcdPD0ly3xpjvKrWvv5SZNtgmzEhQHFm
SD06dbzlT9FuXBbIrSpkHOI7h1ZJjTBxBNDMXOhdDr5b9lJYbNoH9yifeAFyvj59
aSeZFximy/tH2DyoOqbgXmLzU1+C6I0d20/Gd9TrcNZfIc0U953QfV/LHuHaAqkb
YxRIQhLiGwRYlP8LoEAHXOgxYK2Bq6dqhvY2LPk68tt5H1YQjdk3pcVCQBdPBlrG
31+j8PEH2mQirx5+gO4VPhDtVMFRvI1lhBpdGTwnPc124x2VM7Qxo6bCrFSkHkVQ
IhpYzT9OT9TCCO1AEMfHWBmDUwPrHGaztzFyAOqfo/uSotJlaM4y9UuxDXZw9KE/
76xFALtp158nKCBd3IA5cHOnR3/eRpxzUb/5bAhwtmw90lQROCkMCORtp60+U+Lz
InHuXUnVNcZpihu+2xoTs/bi+7KzSm+UuL8QyYG6wPkwlKPHhoFo047VPiKyccO/
djMZKT7LrNGLSZcYf1PLZ4zbSWacfaIbMYkxABcEWA3TrEWKzOI3VDNT1KJ4tp0K
Ew5l6wLi9RWE/pfCS4R3kV2Nf+6QVGK2kWCRA1SDWhK4PoWi75R0lnjnbHyFuAO+
xjC9GXeggBvfiBEr6XlFfI3GiHusQvVpI836DKGQN8A20cfQXNZjTbknHHUq3VEj
HKQ/XCeQlOvFGpek+wxS9Wi+cbbvAlQlL/R5R/gS24zdwcpa3APO2+yTyD7OjQeR
JuBay8D1mgvdN7y8WrZdPhHryz8WivM1q5x9SOR3RFUm0dsPXqck09qT64oW30w4
vec0uGXEBzcpo314uRH4+O/yfWaCpZma+As9PIrdUoB5INUbCXqYO6fuM3mgDAsI
pX5r48w8kDJjh3JG6KB/277SngOVGRGmlPfj7HdYO6/OarVwE2xYasDnlU1u84bL
m15cnrdhkoTbXw3CGqKxK4mqwFOgVd8paF24NIwREyube5UHSvszzCQorDcgZdKL
J00WogPHeLGMOcV/7fLB3XKy9IHjp4TEbcNBq5FtPf+dyQ+QV15QWYZccUyzTNhb
P/8XnY90ieRGIN4dj2YKWNJSC6ENsIBzaltZsZFZV8McbDFYffxA3JNNFNjsi2ul
qfD5CZ0w1UIfqqYvxzKx0eEAsCv7bbMbQQQs1V7ESeZ2QAaZo8G8y6SYcBeQnBMr
j89ZIT56VTM3/iDFYWJBYFX08tAE2nygo86KWln7VF+jqZX62ojf8SSZlLex3rfc
8OUB7+LCwyAseCQ3gRcE9rItk/6rILbcs+MymXwXUGmUGfGfY2eXDX6GwgAYG27E
/TBMD3Ssyk4Zf38idIhQbF8gxZg8CA0aU2rj0MX/QFhZbgJIaOOSq4La+CrZ6t48
PuE1YSJ/Pr12WH5CMQ8Yjg8aYMhnwlrdyFTBkg2i1OAwBm+ZGmkS1aMf1d0uqS5I
GbyQpTvaItKI2GjuIWP6Datlr11PJ1qATcaCiC4jwq5f/yEYdMb3zdjExmrol7b6
xSzvQqVT/MhvUTUOvyw6YDS5UenvZpIXLQz3c5cTDeWEM3lA9aS4F+9YteXgJoCN
Ksi2zIwBKO3ydC33yYz/atbAjuB52hqcg0VgAqZDTpkiUKhhf29xwlYCQNrCThqt
LUT3YUkmwOvZ7igyVSba57OY1QJhOhhqZDF7mlBT6Sv96e6jRfGmTasKKqyzf6qs
eqxnCz8G8mfh/qz9LvQQJKxIYc/0JeV3XKNoAMxic4+JG3QIQUMQg+f660Va9Gg6
1Fh78gjBYVv/iYGHUxD6JaANIBEfoi0O9OeLvvpJhCYTGNpkIXvXABwTMC3xgvwv
YXfs6Otgohv+isVvHOHaOd5aWQEiQ+8msrg+DbLHKDyHHuq6KMo9RIqFJkWkCfTW
W6LSlqD62NY+Hfvq5wUMoGAFZ9d/GDB82jDEZsERKAL4ssM9PbGqrfK2sGYXPk6q
JP7gv/PJTKa8UQZ6o2cep6z4y2eHhR39r2ZdgEWZyl3yfPwmoBqgMOlw55F6C3t1
ONaAPZ7sjzR69+YXNL0vO18ta00QOe3QErN8B4jBx/ppEibCtv2IZJLY70TZeBPE
XlcmeSl/q7ba5BYre44a+mxG44C1uOhaoY7KLxNGkVkFj/DRMhEQETAuTHQ1EaUo
H19Hf4Qpn96qAs8wFYr5Y7OTOknXRg9eW+IjQNK68KmULT6RvnRj/loBdnpJpMUi
+Dw8s4ukD9dw8a7OGvP74VSJUDGS4EJ8SOADt70qsWCOzzHkjdOY2m9b+7DEj9EL
GdNwNE5RGE6gd7E4BgDtPQruSONDhbQ/PxsGv/EKVFFimWtn6yvfwnpGyaWTZ+4/
QHhD3+5921RDU/C/bEQ3eEzRKSyJYAK1AAhsB1pAuOjdG6wjbJFLJ+532PspG5/Q
06Y+sgyVaNvD8hb6N9eo/U+2F1BuL3eA8sDy0oZbugnJ0a/yfSxdcOPuyCQgkemU
Cb9gKxjv7QCnKeHqzv/uBPQnAqMAZjPSPEGfclwidwoeu6hmiJY0XJ8w3MUlCXgs
pmpBFqQc6dxRMyW0PDcYHEtW9yboU0N2Za/b7AgvAloauKOf0j9iTMk2fKXQwi3K
P/YYKeKCGMG2cjiUZB620qoJfN+5XVuAl3Gmd25yWz8XDMZqHEYeVH6MI1ZbceY1
FOVZTaKl5Ads0GfFeMrZ7l/ZzifSovsEmod0/Izt/dj0PcpRhqCGP7I0E23NfAAt
FejHte8rfsUUMk9uF8Xe7NIxt0fLVyrKA6aEh3tP0duCeDYFywELHFVS7Auk2riI
bChHW05DS4i/9uBYPTqqrDyhSZw9QlPNtFNzkD068Vmh6trXuU8egE4zo95lt937
OV4WNrL3nPzf5yfC4tKhS0eSraNNbMqZ3H33t7dipNQL4z4NtzyyeIp7e0vFrbe3
WD/fUmP/XUFj/ITN1wgPFGlCiycLQCmTHGhUYgNlsCEUxkFVYggNpPf4U5u9RT9Q
MnQfth3JY9QL3sSM0n6aWHNk29yePpxUH1ECTRoGLpeRvuDxUrYkcgQ6Zv3Z91nk
N3sVGJQGvbUGinAJdKKqsIkM0Q6yMa7OWuMITo3Lil3CEymcUZJGdXZ0K+gdI5rE
XN7Lu8wttuwYsaR7blKZJqqdSMBW6voIugEhsNs/F/Uecjll+uEfhIOKQRqNzPPu
nEtNGpObSDMGG/mVeYRKxzalCgX+jbdoNMYf7ffa1gd85pcClnxCANHGNGYz4O7F
vfyFezb9wsK1VheUOi80FJS84Rc/ZKJHSUQ85Jhr1r2CZVofYZ08F+A7F+pVxgYK
mi1+dLqRtJxJmgad1R1MXq3041+Z4PU85Tf38Iarpmbut/Daq6zWh27EC+M2veL3
JnnAhupYSX5lguQ+UsOLQhOHZUfhSlLl8y+2NEt6kcHouv+1myNTgXCv5nsEM/q5
yMojol9J88yFteIAtifaEPsFtd3rBFu3sus6X4gNrix+1MSeJEgDJfdF9hR5qeZa
x82kUJOnWc5UYtgDnYiRe30Og6dkpRoec+6OAvLnTgccb+Za3krU6Fvb9N6h2kAE
yhmDbu9zh2wDYN3Pq28nUHW6jKlo6skakF6if1LL8J1DG3QVYyc//hGK4pw0oHNi
RTzY0avwNnF8Emys3LqLxWjm7Fy3OVliJLfqFU7FHEgEf/9VT/Xhnbned6B7Lw32
zfjae7SvZwsqUfKbQr6/Ojb5HyK6PeUVgFq3VMMz68hBisz61nlsnhgn7Uip/VDC
dEE/pw+ujRYS2I3VmnqjInMx08xez4Z3+6yl23Odfp4a9/GMQBCZooXlrho8iDq7
K+LFyVI27bfxvvYfj5u4VFS0wUzhWtSR0r8AZbQMcRyFnJt+Z9qVcFUTi3enNzsp
AR8zgrGsmJqbOSYtbjUiCjJeUy+TWFgEAzNRPo1cvEUU+217i6dzWX23Y1KFL7iz
l5xFOUdZrq+Auzzs08Z87qNrujHd83HtbbvbgmlLRFUdOG+Z+RElPo+IDUnw1LqX
wV4YC6ioegXNggXOLuzJxsh7M1hqz2gbo1ADDCpthDYyyCfDKH9XIrEpN2rQVxTA
sVEVXeKTDQRnpIgg1vpFHqQ1A5YCrAytmUxYMQPEZZxguCqKOV5zKVSw6DEmPvXn
nMAMgmxRi2oVfbF+MuopMoVVafO6CDQmfbCHmJTa+ByZAqfupqw1t+8ZlANnRUdc
QKAwtrbYyEuJI/hBQ21aZEJnP5KHiDG5riQMWxUSbAuK8oR/Os7mh7lMgJvy6UBc
vVnidHPQZ6p47D48lQ/seJ8zu/oAINhR3Nek2jFIOr4LBYnIBxAKHxLzgO/H28C4
hLza1hCASQKRA83WnNedt5iGoCApV2Z2LF7GNXc55I6q1UAfg1aFlBQJvFc3TfF6
PHUSsb0K4U2TJbHicoLKn9Kgt6QIrBTh3AqrXGjnfZy6tdQyQuZwfToa6SJOrvrH
FzYDKHHPO41vtS/79gdzoeawvz0fGNUJUDnC5PgC6zguNDl0cilIW1r/bnzKmX2e
oRWZYim3RPLAt7OaHgAhBuj+/KMw70+OrQp5tGMEABUzOhfFD1riLeiphIO3OYyM
iAonFdTY/o+IrGxqKXa8dNmNXHNzIUaoBBhxg5detPFxF+N+fRlj+rTw3+veuuVv
y42/Shk9Qs4Lvp9WON/S4ofZ1rRdKkG90dDWvem4kYhn+w4jr7Dbz956o8znclVl
NZzMSX7afNA1KqUIEqEiOJzCxgR9c7mR1Sr/xKYwndPDRGZNKIhCi8mzSm3NnUVD
HnuNBvot6WN09t3RP9Sy6fpbJTr2faXRYiE3IbTv0foDAj4rBkuCk0Ol78bpsMMw
/5Zx3Q9RMEpJT8tB2k3sSZXGv/LprGeypzKXMCnJL+3QqTW4aTVyNgCbjWqpE8xo
75l7f7tZCXATyErRVMZmIL3N/Ye2ReymkO0G9LStA7LVK88Wp0djrzO+GilyMKK/
suxlyQNpAqMcJqd5TfwhxZ2vJugqtOLpbhApYPTYMmwPmAjYbX8Em4SxLwgnBc2b
ynPgfBvyLdVkDnGWaUgq2Hl2S3u8FHkgqColtBWttEjHiH01X9B4M9RQpKGUeGew
75bs9/b6+82fPZZATrHUKJXviAOsfDUsK4dcWo73+/2tIc5Q+tMHBJawhMQluG9s
5Bh7wjmiVPSObnyooBIrQxDjQxQXIsGfLlcjF5OUMNsFG1cDgqIxnbS+cJjeW/UI
KKaX7QzooRW1dh493Scrp+51dyed+gIxrAp+uRAAZlb7CF+wQg05AdfAbpFD0P4I
KqXLkvaT2xHPmakYvRdJlSdo5L+c/9uYPMXwlOFRUZ4C98yTyGSaQAlgK0nq3W5h
p1t4LUEJ2leq4W1eY0sYwWuvZux/pPpgN2Er7yAskZxTeDZRAfxPmLJJO2UhZ9Uw
AVt7Rs0v6NrOi14W0KyJ53NWcPZjTi3Nuwr+7qLqEui2WLW0SWHtdpzFEP/XEhJH
cV+EYsjJmJTs/UNXCzk4r0XBHWJtxa5qknbil2uTVf3GydLpnWyMTrxfcC2H9XJ0
SvjcQ3TyeGG+C0oagAfArnYJ2SAI43r+bHwreCc+QKKIGqsOGSc/ZkPilKK+4MJi
G6kETVrB8GA9qGB0lsqtbtGJ+3P/OpDqOvA1dlCTCwtOoKII7Uqdc5V8K18X9sYb
qzb5aZ2tRYKFYu4BD2G7UL+JzynE6cdHiySnXVl/sMWdUjppIYLSIw/qsFEcmezj
0orFVsAlokQ2BeerCzmIUQNaeWuoqxdi9hhfja6pDkeN7X7BHpGbJbY99WyWkrje
9Rx6AZvlo3iN8LmaZ6/0RO+Q/gNE/zpQNDV8E47W9cTQLXeI/kNXr7Pah5XQA8Ys
CALdJtYG92JbNFST96tIMTtbmT9fJBIti1oUgPWlj1+WOdmB29fki6yWlYq3erNX
XxvqAVCCQF9wtffomaQnJYTLZ9p8YZbOPQ8pIa8JLgbQGLS5R6KKqQlbuA1FLoPX
QvSe6pvYtn02RExMJ/JGUa5UciTOhbyZ5V/R0Ic4PC2uO+3JE7MPXEuBzsDTbu0Y
gF5MhTJr0x3q9deV/HlBRBOc9TD0pTvvSx5gNrM46XYJQOz8XPkI21Wm0mCCD3ny
DrNvcGl7FmCzOp1fmCnICtYKdxe3oKgRL8FInoAAfV1JFn3hjgZG5FIktxGms/6F
Mvhe5UCkc2wwSPxJYrxEC9OYgFxZH/wq4/m8+14B1+JxRrzT2w8rWKMSNag+CATx
uD4hhK7LQ4r49e/w7mxiY9xEZmDytPEVWUNYClwyALlPzF5FI8PKsP+gOElqObb4
8QV4Vzrp3UNsQV3bNTQbHoWGO0LUHC6lCDKSQCllrw3BEGyb6lwLmJD5YOyp/iA/
/hG/MiKBdmrMC8RU5HUhovdF0uuzRAMf1Cq1U568fLDUgIaSbkxey9Z9O8/Dtorg
NXzuf3pdc2WFn29Z/uJG5EC6P5TjsVsMtQZK897jkLZtCKcIhHneh9c3p9TqDz44
Uh5Iv8K4x7HQKg/bj6KP3rX0r0zo3Nymjko5UxBCNmGxmp9HMmHYQ9PnrrHcDCtI
EVf4L8IjdYK14HM8CE+mevWqXqPrLq3zFLLf+sY0IKqVsvKL4i+zkA0tPgOp8xYy
rxlBhg5QR06fnCST/+Kv3OdyWXsCYhsW5tfj2YA7IyQd7i2Vzp9kHsbC/EnT+8ri
5Nfe5Izu7YvWoBNLleAFuQARBf0PW7T21zZ2mNRjO0KdZCaY/xCx8OLUx4aHFswV
1AoNozFNipUTq1YlAFh9SRMUtuDwBhlIHl6ectWVy4FtVGGqrwxFBLr5UymwIAKE
OmwrWHa4Ou7YR0/jpUZ+LdD0cYDF3+XYgU5dOx2MX3JAD31AQzA73VDRAXNqTxdL
hDORpGlKS5Sh14cI2yZdLqLmwDI30ao87cxDjFOX8f9bI8Pn1tuwByqAstK7nDl6
hwHMZNHcefR2OROIgsIZt/5JaLcZmVyyGuVoCLY6Ajb4FaAnVljq8r773JaURFdq
5BxPjtUxEOC8nYuPgi1NCyeIqeyaxospoTeJJ6tj/ENIjncFwaq6XgwZTWBbVwvk
AXNnwu4jXSiWCJAC8U2B6D5FzcGjDFfV20uIPSu/Dpyq0w53zlYG/QMVWv/cdKiz
AXsw4/PvWXXo5NZ3Vib/WDwdeUBOgVcSEKViupBVqWnbCBlRoOoJ2i0rPI6xh6Je
IxXSTZsU614Wqv4n16ICkzB38XK9Dpwqa71HhwwqfCQYO/S8b3pK5TRm0na9TXzd
456G2dPImNTnq4x/y9QBzgHc7SKX7IDLefo2leEufcaZ4CUWFpwAfpj00rrI0ZNc
GPZF5tmAG80gFkHpzrp3kiJptE6b6hBQHGFpZCJljMFwj1cp38daTTfCXQhyrqhQ
fyLZIa6pvCFCymt+mT1rWoqfbseXpybhZfeyc3QoXppMHWJxYWDok6ZizUqmwGlC
M9gev1GiJcfpGtA2sy51+/W3zSiG+B4I+e+02ApmlcQLv7IsylhTkZB7/j6Tq8P6
MElr3FPO90lKXMcN+Al8pkHZ2umLU3tW13FOLU6fEloR13nOj7IflSHt1xdBsKFI
Kh4KGLv2jhXWxpv8MeT2YOeWt/D/LFtFlRK1i6EFczIyAIC8VDbubRxsHFnf4kw5
gbNqqXikoH5dav6dTaPwiw4JCl1l1QbFtWQNAX2ZmwXno5S3baciuRni/iHA13dO
Ieh1yWN6moGt93cIHMb6d+ear3+68t8T2G8oSUbMjDMzszV8ctYq4uAvXiSCAW0v
cgHZg+eh6ijjAm5O9GQA0I0TUkmpASHIm3/cy1sWagXTbpZyw6AUjuLSu4V3BOyX
Q4jGYFEWlDOmOqp37E1V1r0mfZsMQzMcrzbyxo+RNpCPC1rUOqqKw6gAQMoSxQ7v
sk93nmc3jRfscRkoKzY+aTLiMFWZSJsAxlr9pFkjo/aE08aL7+LD02e8wVKcuVod
Rcsm9LZq1qrHOKkwy0GOOuBbqGmZTE4zquYB+Q9YzFbrVF2ZOT6QDHYEVMjBvxip
FruwvMyJqh/wOUvBhQJ7+d+6qnn3YUyrgIPIOXKjdMOR1jozhoIGq9eNZSVbvpuJ
knG4nTSFEXq7JnXeiUGArdyOzxgaokCS4AZsbZ5d6vzLEAHqSWUtNApUp6J8zCsC
1bFAF9x0bifW3GXAmn1RQsaw4x6tJ/ebzbK7KMOKz3t9IxjpryQuADIGGtin69se
EFqagYJ6oRWB8QjNajO6QGIDLh8a8uJKGDobzDf4BykwaS+mUgTEE2gooFN+8sqU
ZQd7LMuzeoPLJWELtpWlqzIjKFHLzVSNlrourg/e0b/6ExtGkJBaj4vtN3ZP+ZBs
8eRN/7QZFaVgY+SJp4yXwWxKMJOxw0WOKk2nmwil6HdVz5vVSrgU8IVcovLubCGm
YExgzBXeAb8CdxY0DYZOpxYak9JMuTPPh7R63h/M4Z6GztD254D71Stzd1EhWRoa
Z8yjR644x3Ha/HiTZJxVc4kOjIarcBemWjbdc7spGIHlY1qkrsAA4Rif5FC/6qYa
xf98NDkvIE8WWn+OhlSxQp16rCT+goGO1O4imhEqY9eCgVq7nQOmGqH0Ft8t6b16
lLy7INjHFDUYnRzLnfnwrWzWBbPkTynKCZVmIas0p04iAAm+GIxqK5zQoqqq24qH
gVNNRR0Jz00MkJYOyEoaOUZtWQisT+T9newgvo/T+uCRSwb2NAzGtRq2EzY89RJF
gNdjZdcrhuIYBm2rY+uIyE49CrRBqNM6hl+zHrl3Ov2mxLJ/zKTZqGtWnDz1ldXo
mFmM6GhfjevL8xfIcVRfBA7rGupNL8iFHqGqA6G/4h+nZd8cwM6s8P75WmiR2zB2
7IAqVAcEg0yw8xi5HxBncblwavwBHZTKQ5qvOigrjGSFn2AcgocZLUc8d/0biQ9k
PYC3CbcACfzmUjxMj/7JM8iAefKKC24+BSxm5vTWiOome+k0Ut+lMZFzXe5+XkNI
nSOwm5eOYmHCeNwb0zG+5FsaKCTww+z+j2KxZgB+QAulYpMAdZRhnrF1RWu2rIeH
88k+HkZYtLNs7UYk9W65Z03GssE45cBi+IBRHy41BWnru8N/WbQBWKO6Nr3ohFGD
oL1yVWVEx9mnsXcxIXCEypYFI9IFdZkHYBgrvEjkb6Ovr98oscLvPjz1I514Q2tk
/wF7G+53x5B/w0N8bfpXYW/R+/PHOdDRzv2JCbLRm/bE8/Z1ZZJdip8v+OB1NKC8
550xY5S1QX78lb+8Df7gX7AwDd/4krvp6qveGBAWE1Ok6EOFDm6rig9FPpyr5HR8
05+UHaf8FTZnloJFRJNGMl0DUyJuLvqIca45IbMSJEBO5WcXy0TXRG3s30llkApn
Dm+kPTHRh8qV+Ss4ctFrnzmkTNQaSQloauN5JTPNrqGdX9Bu9/fhL7bZXkdmOGJf
wDImaFq/wM2bllgoBztqQQ/w5lD+5mP6luN6uMBS54TknDDd6+bw4oopRonntOHx
LuzUefcQ+PEeARPHBD2RILVLuJH6yTjs822ITYP9vSHsllXPstny+Lmag0okV48J
V4GmO2686f5SN6dywYmqSdnMmUbQyvM+HgztvoQMyFRukJAL7Z8vWjvRUsNqTnOF
auTFiJ90wrtaa78GPA07EFuQWSM7Pxeygc2hWi9tQKRcD9XPV62/oVlT8MLx2Qyc
Er58Gbj6PQZwEWhzMScNowEdvU+IVN3ZZpOYd5t0q4YZR/NQQXdGlQAeWXhIe4SL
6uDTny0a8MkGeYXVG8UvyWD5x+nBaM1OPvOZQe2wa4g0Rkk4WB7+ScA5xaGcVA+X
7kNGRcAUGA81hJIYlWJMdawJuUtXFwgc6WYwsRDjE9pDf6xuutEm4dNfw9qdWB9K
CxxpKbs8BW3R2H6P3zgpqOUgxKDxryFr0xiVjf1FNU2UwcH+n9R+i/IT3I1M4oJo
GQ2tCIRo92jHZxp4gsLanuDgNbG00aHTTqMntQBuy3A/7XcI0g1d2mym+uqJvxEk
mVhnd+pdLim2tSPaU74BCS0ZEObx+wCrIz+4hTOVU33mj9zR3lTLLMx/ly3Zs/q2
L8t+4cDMqp9t+N2E21C5yB2OPBz7GpZXIKYdXYlDYByQRhwlfZMMljjR0q4b6BMK
7cjhsIrOyBLCBtuBWwJqtzL8Ms0enP294yXAZR5gmEUv5qVswP06LW2cbhD76Ic2
LD8LRsg5qX2GGSqkx0L12n9hYyaNhTdmTFqASC3KSBImkRI7J3XT2hSPdHU08DGC
1OZOjuJEjwYS7Cv/fElvL3d8Xt6h5DC+TFZGFcf59ZGmStadTHhm84z31jmiYDZy
BD7xDT/DUZ0yet4OfYHHbXnNO6OGaZPt2GEI+wW5SnYruOBJSmRZAjhT14zbnE4c
DwVEvCiWkcKtE9PyGsKbCZtlcPRdiLh+kRyqCgQMDmMg9T6EKlPB8GeRijILdoRY
ZlpEs9gdjNefQ/IHlTUyMEsTAIkZ2+/LGBe3sK7V6rqZPJ+4sJwjOx1ylOkPwxkw
ATmYLlk4Xxuudh2LyX0b3MhyJQlWhCfrLbRHr5BnhUHiHgbfYuZQR6ZaJoFsBJlz
xrscXtFVHEftvCIVRuSr1Iwh65VZ1pHfgi/A95CXeAKbDvAWV1bTFSw6ZpQfj34o
+S/VYAO/KAAotLh0KXHnWaF8yn2DetopSyrJHsKaTD9XdXjgwg+KmBl+/z3AYWQM
p9PComZjGlF3Ra9frk6IM9UlaD+rEa+N8XhhfYTHCxcYODre5H2esGACaOjORj0h
jWTNSfXH9fQ0EbRLPN3mHHXSysu3LRHfkJV+bDleqUU8p5AFTgsuzJfYFcKFOr0B
yde6NsBDkl13eg/kc2hD6jV2fMg19eFk2A2ic5yioaLxanFJCuuEreEtJmwI+EYy
D0+OiHPA+qypmgR8hOurasWfpMj6kUBOnu3VEn/ujmn/Qa6ZCfFd0VOuxTV+x+P2
dRajq7WySQGxCEdl9BSRxxMLxRFs8IFeJbCDO1BE8JJxJHVeTFNtjg8y3OaNK6Lb
pvELsEXY1n77aJ8LmO+MHqhagY5dyk6v+zv7A7ovXsUeWJFaBM8ruS8a0l09ZC5P
l0+PTdF0343FAOB2CKL3lLSNaP4eiTEpRrjG22SjS0ywN8tzBVuoJNAfwDHhSNQy
uCKT502nsbzys2i/eFbcDLNVGFn+7UO/HrKd7EmtTowWkLSJ8i+sr5OcKL8F4pwT
kVWuH1IdAk2FiFWqxrJa7q1wH1NV2ea/qSVevFg8ZaOuOYgTEUbgpCgL/twhpimC
ERmIjncciXJZ9K9gZD5MXwW77AX7kbPT1zbeqjUR8TCLLo79wDItbY3UuTS7N2ug
42tm8XFfVzWkhyjOYzrfRYqVku3Ufrn2FdkWnlX/1yef3HKepPPsh7eF8aSbi3UD
mSiMLChgqrksCRezPrf9PKrhLt1Ni/vXeDGQIzulDjnAfe+59y1uoUsBFS2KhA1g
Z8iBB2GctHhiNS7TBW2ZU9kjIsjf59TD7PfA37aAjMxuZtl6GXAntQHgEw62IxY6
pmMfSe9C5wMU2OUF/fLG0QRfPPCX5Zrzkk/yJ0CH3WnYkVufUAY6XEaapYd6owpE
cy3+pJWlUzVyGP7o4gIsH0SoBL2FWnthxg6yIthFg3z4YcFGAAK6HoDLag+++6yV
ydk2aD0LShKdPW/XU/OYumEQq3PklO8SFtrTNoJo5ZJP1VSJJdUpki98yPJK8jr7
/wbDt6PYTqfg2x/Wtn8+BY5/rT339eT373tmIWHMtfcHsbP9say/8///LYtFHmgc
Y6yI0MG7GOrbnTzXwC9zytetPLWRJjD37GosXIUJO873a7/TYps/vxlYwVOZ/5hH
J7r4CwHE7XJNIzDghrx+/qIyu1LDlJaX2opWvqNtRZcpueFDwjxFeSLkuLfEpxBp
cp2QHVG7j8xfwGMb55UeK8WUJzdxucnB/z0I7SFfUSzOlZzxqwjJCE7je3FF8Qvj
hpaIOIZycycngD1+KjEpdH2zNl9yc//WAweshjYo1x+1GyLnfO75BPQz0ea1TtKF
4G/Gl5psIEyq7zDQeF1s9hIYCOrpIz5H4tli2z9N0C4A0JASS4pspPM1Wz5zt5Um
ATbScq8iUXt5O0UBvlYPzVyXeMN+SAYUl2qu3Py0TudTXJSt4EtL+Zn4IqayiLp+
tlEFxUNf10okYTfhRThHuyquXMJQjFMUqM3Lnm5teButTnZ+nqwkg9S8ioMEltR8
O5DFSmgx3GYwQ7L9bSqqxoaUXb60BrI1ZsGrebICRybKQ0BmHF46HC0aSyWCcECV
BdoLRSeXq7a0cXOAHb7KxWRYqkXpXeLtxAdcUH7R96gS8o7HOYPKhhduR/qvPGXV
6CY4ULmNJVGlkk84opF3ZniRCiMVhv7tzScZsHnLtilrmxXMU617kw8gvZQboVnl
OXQ2DGtEnA7uPzCogMEYtjItVGDZmiiY175EfzhngzxmYuHbBervCKjaSXdKwQod
VTei9bq/cP91zj1MKB9E0GlhD2VQ+ZGoKynDKRzW0zYBfVT4Ok8Sxy5xA1SRUvaF
X+9ODtD2tg2aT8KSfizZ8jVcP90baOXKoPmvXua37d2lCCN9dVWQz2+FtkT3r46x
aRhLStrFBd4aa3y8QFV3T8G1rwfggDzV/K7LVGw/n9NS9eeHjPxaROWcT8UI0v/F
nss14sn4rSmBTxvWFrCVVVhX6f7ObTitLdXRrka/MxJS3Z5W2U2+GqNMDmYL/jEW
QTWBrXf+NZAm8nHZ+8ZiUe8HWOWxOYOR9Du0fWbteGOs+bzkcBLvgU5upP1BO4K9
7AOF9rbVHTmXrYeD1F0CGJzs6QbwhOh5MXcrXUES/oGceJdioVkByIanAHVT2NWl
XaTL2dUw7OCYGt9r4wd6cOzylqRd0KF+oeuvmJeTcUismOWyt6xMCswGLXgpa43N
1d7xCpC9DiLZg4AHf7XIgRb+z90P4uNwXoaddtmkF8YHl4Gl5yf4nSFffEMzzudt
AefheViwfaul5xPg/0FaRED67A6byJp4ou5Pk4dmIt2MBG04Xbd4+MvqI2ZSeMcP
TlE9/oFVdjwC/P6rDVHiusuEWQGoy+18kqQ5O2b0TV42eHOJV80XKf9AOe25XlYC
XnO2n/ErWaL9V8+YI3gpChY4pXJjmPYxzETYw73rkparsHoEv8uN6SBz3oFhZR6U
4yowaktP2W7xUpF7MDHqNuO5m1jNh8doKY4eESkQrFf4KT/cXaDtSb00BwQblDS2
h+AMVk928OiEGF+FM0AE7bFz/atKMPPUtVbm7y1TCy8cGHY2y1YCgae8UWPOReUG
gANIV4FbY+/893crwJ7UeY+BbF55jxnJSiepiT9qZT7WLDNwuck+JxN+hmdlPAWA
6YIChkcgUNBzVH+BXwz7q2zDI0lsO/t3n48+HsB7L5IB0a7r5S8fPx/Uea/rGDyv
6i9VbCkWtPkUsAVY/NdG5+yliqAa48kkv/sDLzIuE9aprNl7rpuyOB2ufF6aIICM
lz3yWnxkBV4CruOJF582IVwbIPyl+fMVvTYqNdV9S86Pz2dWTi9ISjW0VdOjFA52
SrVHropPvUmQlows2U8dS0948d/Kpq4NLbUU/vLRo/IQlGdKKOgWOTMkzhCSO16z
m6fdhhYg5bENhUIagT5GgYgTv2lSk5BnpE1hSQ4nTe1cZEJFVERfaWCzMwqYUb48
IMVZ2yN/GEDVpZZWApKcEQSGVli3fYm8yOWJm72QCQk=

`pragma protect end_protected
