// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
2uZFjAJUcq3GtTyBMSmyl8nv4tjajd84zNbPaMQ7EUJgMRtPgAjVvJTWbvEE2f9x
BN8D7tC6lEq5xSuSqXPf2IANAmPtsc273O4nsJ6P3eFI0DEofWVq4S9iq1d8OoXm
BGZi7cZwft2RNHeYMbTLYV56P+qp5CeSxi7Ed3BdyH8/61lvRzrPew==
//pragma protect end_key_block
//pragma protect digest_block
sBzLqM17thmM2wpIu90rzQ0PKHY=
//pragma protect end_digest_block
//pragma protect data_block
m9VnI1Ggj3DJerg0sgbnYssXWiEd9PvgRPuVOyNdVf9qX7A2ChDm/vdYVmMDzg/Y
s3eOWkTc8d9W31qqJI6LRRZewsABqyRMXwdAZSL3mXjwAaI1759MZ0t3Jd0r3sLq
n8k0jxuJAvRMlYmA0Rs2ncvum9Hc33mST45Xp0CrBL6NHOvaFXRSk4vs7yciVnbr
wzAfn/xzLj3Q4orzwAwXoaBamUNdi6UCUJjNgUtZHeS98THRe4nKSVkgMtZQ82gB
YUyu/vntkoCxX8TCuCVuoRXKyfgV38zGIfpsBXC1K45v/NUQ/5js5rBDzq2nOba7
52fJFoa4v0Kz28+Xbt7U9fER61wGzPmbZadk0Yi+YusEDnFklcX72Jjc/i5bTEC8
3RTiU7Ky8P2tNppAe5w6XqPgi9bYh6MtWm08rt3JSyLoVMNvTxEtCfFua0HXfekO
DQsXLFraPZ5HQHSiGDB3yqrLLfgLbYWqKfYtZRbUHvdbeeSVu9Mpg5pRxtJ1IPFy
BwyL2/FnXGbp0T8wcGs/6YXrLrhYbPSAbC3WR/i/FHtYtbf+XqPub+3psSTVM6/E
WWY+On479UZQXOL4E5Hn5X6hiQ9Qkwhnzt564GOtvylNdMpsO07q2c4W6aDarz+i
i4LG4p2SoD4azkyytAwM7m84fWGldwhYsBRWEYtZI9Q/MQ2zSOpoLecISYHA94BL
O6xXvegM4zfyPJ8ZVstfVPo0mnr/ec/tq2ymoaDXOZmslWTAht1ywZEScsSgQVjm
m/bCSsnrgVKAGQUQMn6n/R1TWE18yB7/ej9nA3etqcODqqm7tk8pRMWjTiystUqu
xaZtwqNZ9utVmHf9MtDQFpjt6HRB3230zM6cILJ3Z9+SaOzLXJ4DH5uZd0wEVO4O
KsuZ8O7eul/tLAsZHBASi6A7p7DVTPCcwbua1fUclLtYRpuU7/+EGSQPek/Fv//a
DPFI7pEM94xP5aI22+0nDtSi94RL54DTxE1hqPOo3UT5Ls7t4j2aVEB2XQXILPZ/
e34SDro6iFM27e/RDnEZKx2b9/QbIK205cxwfsx1/IgS7zXyQPEYYO/wk3PUolGn
AgMzr4Wa3YHJeUUc1nd0OsYGjexTzxxk+Ff38QeJJFmP2cJw8mUUpaahN0ptGUw5
dsDfesB16j2KTtHRfJyuaiuZp3yNPDjPhH8v2SxPMROTAMxDGlntygxkFCfvAoux
tczm7hZLrz9DuTnFgl7C6X/iFEW/8cnpGmzNcgxsE9PkbInm1ZuQZwuU1evwa1Ld
Js/OEmMBLqER3gHot/EBQMJW8ASz32Yro+CXaQgJpXz4vDXF9B6CycikqhDJQ59y
JPsAGUh6mW8KoORSwN/nLR5BnzeQFIxrGKsFQDfBH55m1gxBkGm2HxZk6VyMGm7f
40DdYaDHTHlNwdyzWSfHFp25d9t+F1FHdHO3LSyoHa38aWmvbW+SlEG3SPTPTrFv
ru97SVvDZ5WAjRgo/3KbFPbE3258wCNdm7MwHFjafE92nVe/nO+BCRkY8Fswqxu1
p0C5OO1juuAHlj1HUA8Sc7fHUXkZkn1b3ciVIcH1PVJMp5aNLmF+1WGLdExlfQDn
1HBCbRVUW/7Fi9pEsqtTYCrx7BUd3mwv8owU5kYebYufg9Ax5XoqHeawER1644pE
p8Sz3tTvqP28fMp23zXeFU/XYTHR31b9+c6gROOr8dzfzXMUKYFpsmfTWP+ImlNz
6dLzgtHKExHLhzsdd2SFs7ADcaflQImNsoThKV2MmvuwHVNRrYZV3zniCOG62Ad8
ug7fdeavBFJNuXLUzmeLP7wd15AsG4gG+QI/ONVCLHaNwOSTE1yGHlxXbIBsmzXG
HNbKB3yY6ZCloR2M3WpasGJoSUUtKM/U+bJNhPp7nNkgL029LTveWwW+rqvqXEce
CbcocGoQCpeRskDo36/9/AUemO/0Py3mz8QoX8hEsXOQgEeWFvQkDzRAr5h/BNLI
dWO+g9QHGJnrUOFR2hfx9+l4BvqMN03Ke08/AHZf3pdsy+Y7ygmzhcKuqUjyhgVY
LZ3mBfReQQn+QxIomLFXW2MuzmzPQMRWUzi/OGPycKv8prTp3LqYdZNKqDdb0UGt
nhKT5970XV3WV5ozGW2gOXlJVOjA7/n0LE0JPDsn2ohvs9ZYk9wXyKwYPLCZ0Eyc
8upFnVdAIF/Ef4bUOXotwNXZ/dTWRiF7IXku0AAbHvoznxT5wtGUNn4am6svdISR
jScbdQyaNe52fXifD5z9kEs00eWUyjt8bnZeF8LpsrrlZRlmxqM7PE5eJDb3T/YB
bpLC5SL/a7V00B7kHNY11ujbyf+wMOMqXiPKk/bBMW5zbzx345bL9IDHG67qPXcB
mAeboI6LU3OsyvpxIFD+ugwQblKU2uZ6ZPn94DLittp6vq5GPNaZ2Os6PTY1B/DL
34cAAFzvkaknWiIaSJ4NgtD9zShJo8ItuTbJB+EhMfC+sSKsT+W8b4CINWgNO398
mK6vLKaIRdX8fpt4IivyLz7lmv+D5yuZmPZhRCfYrGhtmGt8hQ9IGx6xo4X4Rofr
gvjjpBMdDi5B+CBti6MV/Z6K6MCttUvf/yLcyREFlGdxxDb/CKyYpyTMkfM1ucOq
WzMZrUApcEdJ5Z3p3Y3JGkt9FjBepnbpFsZhPSl3K/MN73300+KsLeIJthNY2CPg
3h05AKDrImV94oDtxidDcdHjfo0qDCMkk6iXoblX8RkoTHFoym//bzKdMFJwkwYa
A2P+KdTOo5Mn8+kZmrw8h+I19BzpaIk4d5CJH9mdnSRlRRHd3B1szXj+Fz4ZYYcm
3eLxG/8mpmWOPHQNQuD7wv5OupAOorcTyx/Mza1nMxu0DNYP7n3m7y2WSprUJIvT
qW8G8UR8rONPSnzN9ViR49HXph7QVpcnF3ezh2u0IVeJ7IpDloZBkJDKgmrCE7Kx
FW9NVnojTEqYFYtZd77muhvrxVGQboY6vPcO5rBPsAxmfGngOkSPUr1ZcQL/1qI+
mi1ku/g7jhD+On0jPwxrA8wG9mHjZ1rkm9ER6VXvwOYkuvH801TOjGCChdm7SJL/
tantjP7N1MONKjDfT6KlLYQjknCqz2hX0tXi5rx9poYGjJhxQT8k9VC4jkonyThs
inmYbZ50VWDkWn41hUMFZjU9OQ9Kn7nl68t3lCh4g8Ehdk1FtZ4ezWhvJtM09k4K
fcpvm001ICO2oxUTWdROrZfGbViwnP4yuUZryU7oqojFLqbASyJRgkd6qSy7E4Pi
nzEFh/IjmfXB9ZucBBRQ4N8yU8YZCQ9KoSOHskWHbvlrzmXviHc/1V39VTvBI01m
r7ERrePOAjMlivPDXq1TPogR6QDpo/CYTYNB5lCt4QwxQSdHsq0kMN02dhm+6H9O
xrpg7bCQh1kt2P45axRvm9EmSJyKhsYzk2pbr/G77V+WcQ2GSHn5iKP4rLwimeBd
U7YrteeUitqhjWBTF/AXbp1F7DCwe7Sattfu2LFTg5+lH+gY92Mcm3blVBuHYIbj
WkkJ2AOmlY0+ibWfDYHsBvOsVdqttGwO558Vq/KIi3UD0XyQO9+8d3z/4Ss92AWz
mNY1VKbyN+Ez5JUlN38m8kmTNWREobwWhcLvVVHdL5NHkocpoxeaLfKM/rsn91ZJ
86lBVWMgP4grt5nHW6r8CYXygzeWhoAiak59tasu1GmxcB93qdTtyosLNizi6i44
XkQtbqN4nmcQ7W1ExMCeLw6d0c0DQvL10BHKyQtCS4kUhJzJO1K2/G8Pii1ujreM
P0L/tkhqQoIzQjmtNkAxIEEcWuZ0iU9SLf+S1IMax+vzuv6v6dCItKDc3AxUJz83
SOaN5QsnUXblEuXfaiuL6yYLMARb2GyA96QDvyqZyEVpqeNs///W+YLatJDPmAGk
K58JvXwRzrBJBmd3CXQAmvJ20PsBucXiPjC0WsknLZko9aZy1dW97uI6CrI4D+o+
71iq0+TkWH7RGEBy0IRttiEKYPtUaHVCm4L4volocJirFHcIldMinGubrekXOe96
3NwJHz4xOQ2tOMYqn2AT9dHY0KiVAMzVesrrRZzgF+2bJmxCiLgsr74ep0l1bB3T
mxuRzyQ3MBPBFl0JhA4PQi9aCpv1yw2NCmIuKiFXuzpO/0VhuMx+PAn5USrBTtBF
7ZMBvVQS3OhbmlHI91WYMFDkEY6roi+ndwuMpSPiHyQvi8pJ9RBLsyjHppQB7Y4U
KlRP9FvmzwfL3FEEWjr0I0HhATdgti1qCnbcO8gGUV1bWtLoEdIqADvYFDO7TUC5
I8X/Yq65qYObRbS5EGloYfhYWrZHvImW8QvNr7QgUK4UFeYdqzOebR9q46Fml8cn
3JM3nYtOaNPNa1RQZwVFBZZv3KMc1A4X/zdVrCB68pUjrFBo8jPkiAPFSuj0wFcX
vn+P+kjMsgYqpqU1w+IrRUafUUhdq3xSyyyOiu0Gh2N3Z9pBICRgZrfCtxiJRW2o
sZwuFg82LUobEU0vJlpP81zaPLFONfGyACjllQhPPaewzH84qYC2hZ+0f1rMc9Xn
iugw8zUfsjugOXk8Vck0g08hzRt0YOhS1g1RuL4QIgnpgjG19SD3yeIHcfCe2mUM
WmcKju+0ITNlGw52HJyZV6xbuZ7gL6i5PMjHdt7NJ2rOzQppr2BuSgAgNBPDXgGb
Pw2RF2hVSXwbJWi+ZwKyj7td4EsdNvA7F+kKYhMYGcQrxC03Q3zrwBe/DV0RH1RD
/4Hi8EiGKfURVqDOaqjYACCsGtDN8bUkNo/FN5/yVZ5RdDOIlfXaJ7AhtshRMhdL
WzUUW6uHDYpkmKMbN7Jw/wFmQMecCNn6JgFpDcix7RdEv5wVAfy4hOWVMSbdLx5R
5z+dLmtqTtUq+LMHym1zXYnaREkguz8M00lRYQ59dYkQ4Zf/Inm+VXQ+U5G3TdvC
qrf1Xo4NBo5FY9WFFC2uJBg8z+SBLJhaWIXS02KAluYLeAvV9TaqaIygO9U5G7WK
qgUzhCjolRWA/r0fRBci81PiADUe6KK+BU6L+8sKagl0dnpl1YT3v44OMZ+s3EzV
ITOwF8RwZXG4dZJMgRYfqHylZafHEONvR0qufoHh8Prb39Q9Ae84evjBPRWRPBMG
UKSS5ulqSfZ9gg3ycLCsdhmma8bXVXO4sSu8Xqh2tM2wAb1KXc8jRAcm/exCoXSp
57b9JMupHvXWXREskNOHw8jhxIQffQmwiA++utaCt6D4Gha19GAc1ml85U9/YNb6
B57gRcZ52QW6Z1w369b5uMvhCNsk1iAbXOJsW4PFU/RC5zT/fX1SKABJD4YQ/b+I
hAbzHkbkJGFvX5kSN8I0+tmWtGjZ9jj09nS7b2p7J1OphVaOKYB1snfxd/5vOJpn
g6MycJBcgm+wkUORff8or8ofPa8U9rufq1NAdedfhe/Ssv7+Dh67RW2wjpT/ie4G
3iRAlTllzLyv4Q/uSh17Xn8QKhvzOhTMZX5mbp3qSyM89EBQcL9PiKUq4qWRgOjD
BLkS5PGXveSwgH0vVesWSkYFjFZCiNYSYyGZgEShByilVWrky+0y0qH5UhWiwDdf
W33mEOf3e+uSSf/acD873WYLKQq73TleoQHkRWfvCyM/XzGVVrXw+F/TBndqaqNL
o16tVYsrdscAeAYH2FAz3pGKI7asd3NT5bjeKdbi+eDFrk68AvidjFBZfxX56wDj
RIEVSmEkhyLHp4wbx2n6Qd7W3R/DXhFAlzXmc28bhr9ejtzhywDKbSZiaRvUEQzE
L5y6RuB+UDjuhGAYN+3dQjzpY30/hkj1MNXFSTTw71ZHbICICMmRgfLaBpFvLQw4
ErJ3Gi6fWUwZttTHC0vMznwmv4MqKjHG1q19nGXPe1NMb66wHzwqVAWEKujeJsKf
EnucFncUV6OpWPIDZXZj/2SnFo+o4uwsLEYcDeLZYM2eR6Lr05Bwckdbb04gGc/8
Aw4dqg6j64lKDsckqOrOutP3oKPqZ+SqIL65JZy0F3HOYdwowRzG6hkrynW/hLTF
AslcUcAO6aCFNNcqrqzqKdDxHSRTYE9/3i1n9xbhgj4SALGSMWM4Za5RKq2foy/s
GwJ75BAR71gNZKvSfMIvxkL8V1G51qlGtikCLTao+r/ioy6p0SswcLxiLwAdXj1v
T7aNzV6cM5WarRieiETkTuKEVVRUAOXcKKwjvCJuUg6YTcRXn1wy62r+3yJbxWxG
cnaspP+wEbnpPuUrGIO/KHAo1SFMQSifPCBwZLZvgLFGeXEgAJdG2KsKevo/erVp
3cmeCf/6LKwrwnBkV0hwsTsP0JydkQMJg8oldrfrAYjgMTEojTicDiT3WH+mrsvy
SQpPOB78C5nAm4md+FePs8iwXOoJofl7pvNzsiLNXicdMks1cM7Ch5OoMtnIgoH3
J3RSbhrEieBdQYQwZhfZNLQghmmbRXhDF12CS8YtkFnNaGxDd7a67k+z7lGwARYs
Y9VB/tbF2Ij+LQIUohR4rNT+3TEkFkfsE4KsjQ7eJcqB85MuGTmdd9RsU4E7npRI
S/TArOtqwxbvBKZdJIYc7iuFVd77KMUS1NkjvUaCCNTVXFBsOjOxEUvnDbrms2uR
mug7+k72588LSDXGo2GVCMpFX/YCAWq24ppCmFd63VYII4R4YaMSttjd2SMah+et
QZN3Bbnn2t1fejcG7ogonWJCMTx/GqfmpB5nHKPELoYaT+089lRVA+QmwOGx9x3s
o1Aa9XIRgmXLFAARsL+q58lfFtiXS9kSzqrVGpog37rRIVHsIldhrLxWq+PFoy5S
i4Mojv5ZfQPiKIcHaEKUqvysqYauefd7ALbzGOO80bMFr3TWt++9k/kPirJXLtmA
4Bixg0zscd5H1TGH8EqsMSJtDXZuEimBKq9B/Pw0Z/JngcSdVNATs1CJevQ4NW5H
jlIVZ75RAYs8ntzSZ809wj0qs0pMK14X/N0iAN75Pj9vVHn/UBxBQNS1iW4tTpLO
8yNbuGy4o/ISaxmoj3osmcwm9Y7XwqCST3ojGinRhUlurHhWn+6Orzpk/BNOtLQV
5wub9PNcGwZ5h+E0qPO5ejZFecj1LfNW59H0+wzVL0INQLrcuGMwfFIgIe+8iy6G
z/zIVbVwsWLWFbPCadoUy1sF1B1sUwhWwjvX1UYHEHf4ChmbMwBJ71JZ33p8mbFj
Zr3PXquPmOL0NJC2fsxciotkc/hZIlbp46QEfn+TFEv38Jy/E97S5Ynt0R6wdKdi
rL8GL9oXbS/pv49YbgCjaZQkGlpk/JsvzOzcZHEEhRi+yYB11K+S68HslGPrzb2V
suz3QsY3nfchAcbcYaKAIJvCw5Ab9rnEOEBjI14KBh2eI4kAk4PpP1EjmNDrEJgL
80Pc2SExNI3cR2LRC6cLQzMGqltILnwIcoBuLmrdK2FdLp9VkX47skrAiOa5kgH/
yFGX3uC9Fw80/2HQEDu+SUCVHPYu2VKSdA8dymfkUSz+hTGsytt5lUX49Q7IsLSI
xgIeHRaZOKFHCLWBZkSmsQFzUY4kinNDG9NFxR8KCJZXYtehVg+pNXLEC1Guwwlj
W9Lck0SZ18alhcnHULVHJ/nWbZIrKvg5Ra2YvfFMRisCI7tPWiFsq7FdEsjHAPms
DpQmwPFjIfJDCpvMJqEF4T8QS9vQqgO8cLkbfjEdNWJ8/CW82/7WykT4HyRmTG/+
Gqw8WDzYjHSVdxN2CBDRSsMBc4DZbZZZ2a1Tfdz4RMnQwHsqsi2mIGbS161uekav
SWn5WAlQNPAIh8DiEHafXkWx42F5i0+Scmy4kkQe3dPqMnYsMGRmdrIIpcxJ+n06
ZytDBQWBLUHpI5En4txCfrYa72xh8e5D1WA+1Ogn6G4tvASrPhLOZzviamsGjN34
mePrduwEnuC+1tJoyGrWcndMZnf64YmxMeASZuTwbmaaCNT6X30H1viM0Xl0Nsaw
M/46m+TvcGlvhR1hbqFJaEFnZylfFDdsd3AeISugMRbTbwYqLbsEBVcuauvePe5a
HhnWfOMQbeNylwIUcycJ8JJfkr/PGjJghyt3ivyPncZ9wIgQ6osB0JFnhT7JS7NI
5oc6KId5VanfpCNH+Q+jxFw2yxgCOSfdfaZIh7scqXa87im7m63MQKTSIQDg6wdc
8a+fkFSUBY0eSdHKSu8H8vmqfOIuduD5O47g4SIVyw+TNh12uYupprCZzX8iLtYa
6WIxl7wKyopKNotnFLW12ucdOhE7NiYlqasaeA0E3CmDy2uuCGbP/2A+lSuFLxkm
0rzjjZi0IN/K1bmQkds9Yt7dKeeozk6jaO6LCePgcVIgwxeA46opKPhd4nmq+Qzt
/UXJ+ytRQaKWJLh2PxEG4f2t/kNTnAUNOwSV5FdhRFAI4HPkTumTHsU1dX1xTcvX
m/l1p9xZWEw67M9d0/r0hGREV+rkMEktV2qX2pbmXw/WqVOBOotK8RooFU+/Zt+c
ycKGUle57AHfXc10rMKafm9dAa5IkEdNutJ9PVhUc5AVAWqEh9vBA46+tW5EpN5e
KkGYe9wEdGmnQPaJQTlG90K2MkcNFP20RLvSj5o6Ng3rBe2B9WuFn6GO0OobFcR9
gVeQlUBI3caVJfXnG8Aln0WW2HuDebaoQpfkLjAptls0tJevp82EpGBDPax3maUZ
195S5aYwMAG0YHKrUDWfInZWB1OhlE4r/eS5c0e7QqINoOw5IrrSvmiQLbOG2oeE
CPWMYYC4xjK4CBShCsQiACQLhAFEERzIjH0M5XyhgP6aWmrN0AlLxJH8Uoq1FfYq
slbNFPdjksctIPvkoyLnqbNhO8+cIUOkP0OAQm7pPdrFBjdpbAB78mR8uatQah08
Y1aouDFfjQg/tmAiXQD0KeKUCFIuMwJ0BQJyI10vWbXHevcWPkNBVvZnFtBCAl6b
L7zQLfXfdWwJjZlyhWCvcd9gdz4XJYc157Ask+PT/P8wK+qz6athQpt4AQcHE2k5
0DnCpM6PP9R+s4+PJ0lIi0Cdd6kwwx6PrSDN9//W6O9hID7NOD1aOYFS0VkyGZKF
wyFHzW6DmfLFJwv07eC9cwcI1UqaDHUKF4Txw8DJHeQ3dADiBCwJtDkkUGrOrodU
2nMVuyipiBCWXZzhCUmBV1ploqwequM0Rp7kSLkxx2slrBjoyw+AzyvjkVLvDFLd
GzHI/p4bi9pWKsXF0bUjgfQfYM4FHEGHej0I3RL6tQ2p7zOkTRnKCCS7Ffkozxbq
J8DE5qEsMz5fEWVzhBxdKA+R3cevxuYLb4OsYVAkwQMaI0WCUQUMIKB6wY9/Tt8y
qM1XcOZKRl6jX6Juzexln1gEjXpQ8CIsb9+54Mwz25slqdwYfZbeeyEuIJjtXhFi
QrMDgo94H0pYLmQIvBHhdxIP0CYjq1jAEVKJQGSaakET0W1pBqrBjJwdnOJW2n8J
AtfLYW8S8/lMEdNT6FyJit9a3SUDGjv1f85ojAAqRmTDstORNwoZB0iZJ4yo78hg
8d2eQQpmf4Z+8QypJ/b3JE7m4JHGIVTmIZA+EbQUdSyGNY+nCusqghvRGsJ4g7nL
S3MuKqFZI125ZjMGpmBKta9aH5ANTami+iD/6+TF2tW8X6Zz+sKl8PXopoVarNg3
UvwksGfaAFxGWlFXFi90hsRQabje+u2PSXRJZpn52knQXdIL+a5xtH46L7+1fKti
w4Ge822aIzENKGTcoLO5ekC3xM5MyUOgZRiyVxN9mpPGo52MjWgMVIcnQ13t0qfI
kiAHIJzzmjUU4x167oVPK4rAmhMZZxs9CoDZ9A7emlhByJVUcw6QVfNO3JUFPq8X
0as8blv2rdBtsW3qB9dxQijy7Vdfmhw0eb6Uzafoj0FBa0NFNAVwi6jC8TFQGSKF
BU2wwaMqqITEblZpg6vpyK7fkInxIPP0sr6Igzt9djfCDB9UoygRFR0M+qnyf4lE
CD1gRv5ZrjuxiQkUMC58RDZcLFzSL224WfVbtnSyOEPyA5VP4QSw46SxSlzhuJ9Q
jQqP5v0jihGNZMhRzUEjTYvX+KAosyjGa6qmArJhedvIfIdMc2lFPBGvXdHJ1z+c
MPdooYKxbOwcMbRUVBRo8GrsLiVpiWrd/kZIQynT0qWDMXIk5Zv3+VPaAKVWorEs
bbCyTpsReqz2gM3Pjm73QtxswlFYaN4Mu/K+nNMmTNZHp/Ds1aCyUvMCncbMr5bk
pP/pX4PQ+JCmrQcdBcXZ2dQT1+bh3jL8NLjfKpdTn61cSXI91B+lkYb1bwhjPI/5
XTGq3wTwPp/i5lsf5+BOsfKCiWNlTrM480ci/Pyw7XuVmnqa08G7dkBAUmsYucoT
PAggK9FBxKXZTQYgBvZokOAo5meI7srAbmt4RVe99MElmzJz8R95oMdzgckc7BrA
OrRlcpMmXQIgO6TcLhOnMfAQXzfOKS5IORJu8SCUkFxSO+0+tEWi+0DU+aajy22a
Jyr6s10lYQ531PfkRH6G/PdTedvF4ECmbYawDxNMFpBE6gSr5rQUdiK7rtCi0z5q
kCq+KTmHpo81NkRizWfDJDHg8EZ1gVatPgV+3cd1BXaDa3g+W+W9uIbiIFpuf7MH
f2IVmLcdN2tQ0QL0bhj+hMolpbFansH4kTsnxiM7PN6qA1c4Sf57vCQqIB18EDlH
ffspKOjMi3MNvn3IMwSwNEDyjnxfB0nJmZy0Ay/Rr1jmq3NG/c1xstVbhW0zf7gL
+rP6kPeGUVlCJiB7N4GOiwFZ96kMDghJkXZIym3V4KSis5HIWVltQ9RKCJp9BJSY
GiL8nqvsEvfuAqeQ8kodcPTmxdLnLbR4hFEYtiWfys3xSq5dFLlE8CSgX6XnSnEv
z7rOHWDqVUriJiiQB6PDECo9+dTjP3Mphzf2wX5Fqab4fBdgbFf6Z6Wp5N7ssBfU
nbJkzHhoWGMEyDbNI1wt/2foxxRmEAHyHF9ivt7rVwPnjrQ9IXGyey+JUl3HpIr1
yxTF+ByP2plpYyeFFcJPRWG38WeeuYE8adbbW9kliiodyt3yiT7JAdJ+WfEkh6e6
WTosgLES/T7hOAGQuCygeiH4WuYcNTggLiBKEfqpz+iT4OcxYmJwvLp05L91FVfO
kmEiIwxXJWwH+1rpm9muMnHbuo7qvj3TrgqLInIdmf5GA3lieqqvLk0BWpv93jbw
EPx6jrQKj/IJ3nj/H/k1N9d+c4FP/RZpCVJ2mvpsrZxO3LDkPlMybiuYd0tBLJcI
YIJgB2e/5Av9vx54iJ2lzdR/zMS+2X6IQ+wAx3H6cbpZSZld7VR5MmojNfBhi/CC
Nc9fd15yKtcDak36JnTom5PbArN18jAQ08KvwFyEUgjjcRZEZylVTL6gM8yAAfkw
8chYwRSc1wG2jWU4wSkUgEizYOIMYP9ns9k2FDIBldxS8Y2PHBBY/yw4tqZHVNTm
A0DyqJisFXHmgdoU0VCpj651Ds9DoXintK8ps/cr6066Dq1HV/mef0rTWss6qvwk
aOivqXpc24ZefyUiTUhBXTOfnW0y/jcmjbfMyF0z45T36jRdJ9nKWiq55vAwRAjm
hSuFlVd0jooSuOTdPYa48rYqDi16YFvzxB7GhxEK08FjSHIC0DcWR4AZqlDaoKQo
t6kduLxRi+/WqTp7hUt3nz+h7aGW3hUmvcTV1ExJ6hy0gP/Sd2J2kPTlMSSEO2i+
K3jGwIWKuS5ataGW7ESFQkwnjkfFG+Ab2bhzUiZ3MXHnPgYEVUypFTkI22SC19Tw
edupc1i4lWElhVcYDuJZbHUw4xjfiGrHWQZAvrteYxIZgtkTPLlT5ocKzCqvcJo1
hK2dhd5D/cItwLrIrSjy0T2nxUCafMyjFs68qo3t1iyhdrcl2IcHTm3Q9IbWgRTR
RzZ8xQ6fLuNwu2pJW+srOo5CbH2/pZoladqEGrGhmQ9hN3+n7vRFAUY8of14zgTF
4AHaoAFukTh4CY+yaqlbbWtUBzlYI/LqRsSXycffheKr/LwNk2g94HRI0GXRTZK/
j0IzQQpUfx8wF2ouuz9NYZcmivdH92QnrFfNJYlf9GmwGtORQvPE/wEsXPfGz+Sz
kQY4llv8cvEvcY0vcXs2VtTiMLoypzRiykxwQEsVv3t5BbAQj88cjPHKxLonWKJF
JFYF1uZGdQmffcCxsO2Y0FEX6s+rADxPhDz/vHPDy5UTsYCcmSHk/r8hnXJwCXbD
YsmAXnx4IuhBl1GNgSSn4aI7zh+W8LL0R03YdM+1+mHeOCGtsBICeuyhPTnIdbFz
iF+1dP6ZYAEFK6NMHqYhZp8vBvCJLwWotIzKo4KpGS56lFNfXBIuYedv4882GVAY
DPsyokSAlDO334Xb3RVQDyVRwYi7gfdeTfy7N+doK99tW3JYnyhQOLhrDAz3wMgt
8W6IJA9977lXUATWDeGlkPkS9mnzokTDzIncBVIYrxKoWJFMi6gFQbvIt6gCL7Rb
xevCzXl8koimH3Xioeo0nYZPxnqs6ERTBuL/5KCFVs6fA1bnrJovRjZmHo5mkoJO
3ygK0b28asiG5GMi2yF6XNRKs47ycmpTpP0mrri+258E6pai0PBINMU5d7ePLorD
uhJsziOfIYazUr9W0CvoOvV6mZB34u1cgd8ThciK3XO5z6fOgiAkym3TsSjpxlbc
idjz2UKBpWLnjkeOZUNO6SpJcWjcxTnpT20YVSucRiPQjxjpOwAB7MY0sGyveflu
1VD0Rcxd+xrKk01tgfpH0AsjczloN40fy6HMa4UdEnrvcW2loPW0Bnmm2vAX8XOt
phZ6B+QxMRdotbaFhdD870YHYFnRcJhuNwxF3PcXyP2AwgTW7f7Rjz4aWirlCRio
ygMx+0cY2h00g0D/lKhTjUNqrEMAlBv6GMYCArL6TN3utnP/z5uCOOm0zlgHmZoC
vLD1ATqx0h9sODORoWtIE4EoGKzfezq7RkI9MHlQghD2azpv8xLufggLuE2xQ1mU
M0VEMeVeO3uYL7UC7K0ysAnZKs7k8f81Xkxnedi9izCMj1x6Rffi8WutHwqAUItO
SWE2kSQ8VHvyt/tj5Jz2Hd0a4qRtKlUgM+1OwICbV3kx3od7wUTQ4rcxHGXwjW/v
tpBCk4InFqWf12wfTPfSqLNrdGCIY5yIJiFDXieG3Y1swsPomc/XjvSK540q5J6F
+6AONPmhwTpy47xQ+CyQpehMa1OCtJpeQXTXJU4gFcP37o3HCw+94qgYrx6OmJ47
60G6bLJbw7w6GhjMmGeeOqCAwajZoFyrbt1328kWLwEPg7W71vWC8tSlGZHed3tc
2jifQmOjbF/u4gwT9UKDIgFH1TyUJh4tpgeBVguxtFmBX4P1V+uor5HTG0S5okhO
vkNRmZNXZ4vk3s/VHFyS34cLabs1R/AQZTZEMxEbyRgn2B5BSDZPZH/o8kQtJjHI
ZzrTc+jtKJCpa4ihrZtGjO2tG67lniNpU5xJXADzTTKHCzLRy5TbHCMZY7qkFkAg
XJjWtNNshCbFkLYlTKCU5l7Q4dkdAW7Do6GOkHwJwhboeXD+D50airNMjw5g5607
FV9az5pYK2izBk6pDordIoP8FY0dsoKmz0lxp2kpzFhubsm9vLXD2tBxIyOlGIUN
9egrb/sen+t5Y7kNlIr8F5PBU+mg6+hY2DE7d2MNQpsxdm++7O1vPw/ooIvY/mu3
ffzjcuZ+WzAwO3jhd7jPb9ml5sfdOsJ6Cl1K7B7ez69kcN9+kI1kAWPRwjLwYei6
bEY0uYdRl0M72LW/3o2dSkVeQbUbZOOtywfPNjx4CeONmNQYJEOMeChzzIKM6XKK
DjYA3BTzRNUFuFb+PbhAaR+Nise1PcmO095P6b6m4WT6UzwUgQJW4ieWe9kmZdn2
47KkXtI9sAhbKR+1LqP+SSg+hNWaiOiugXIAVpQWl7N1XQyhcl/GSxJmTRekrfD5
YEZrDNovgB0waitmYRe2DcUgP62qMbaIcQ+a7GuvERtgtykIs7UTv8mUzAF/Ug5N
EtfctCR6JghWwjJN4ZqmYqQN+rsy0ddtvEV+PXjc0yicUMd8U4P2ZqIS/Mzkh7Q1
ohnvSctRfCQJpL1yqmHPuy/0tbVe9RqNdoKHdTJqrPZs50zqkCWi0vS3jMMaEEhd
qgrk4KAssCIAs3P5pfBKJr47O6Du8oZ1UbwdmWSPmGvZzEW7CSupfLo+zQMMfqVE
MlGrAPuU4fAKyBkjCeI14PT5IWQrolPCgw2BbvZT0Jdj8054SPXzxnnXOUJmlbpg
b5C01SOCh/f/ZzJFZLMAnQxVXL/IuR8T4xMFo6KPTTEhApk8XTnpyZhHKnug25PO
HY5VZ4yt5ZwjcrpO3im8g+02QLjBDMia53LMcsj6uWVuhBZIz9WnMe2/TVd69S5w
3sAkZnHLoeG1jCez+AERMXpeEd7HKnfuOyeU1fWkRG0r98r40zda46CLUwdX+3iP
oPZ1yJWp7iEMRjVjFwBGv3jYJVoYgTD3FSnLHec1XRcAX9UvkWYHlcwxSkj6AEjY
FBb6VzS+w2jHCIvN+T+XQ0ILBKvM+D4E4CbdQFxVI+aDs/bInq8uUuVLSm64/Mf2
S0Z+ANbOkDEzcZlKLlf4AudOJI/ytsXZ/1vaIjzA9mHTIhAio+9RNIVbNVq1GGgG
/NiCyd/N78yvLfPT15s1hosffltPBHO0LCm1spulbfCvU14aM42bw0ary9EOSJR6
JmBG3FXZ68j4mp5bxZsHBPao7MQuBbYhBO9d/ufKBGRLtRXZeQTHIrn5PRiyXzwd
1Y3J3QdKDz3/iIY5fZSEYXgUikTQkD/bIKTWN9Si/yGLvrvpv1KQDAle6PebHCcf
cakg/u9Y5t0vMDsQRmqMuRkFJy5BaDV11H1kOLiGfgNolGMm9wr9gnjLGan7JJ9o
5bzR6aF8+gXtAr6xQQztoC9Mz47MWdXmHii7GszR9hfhlDdLGpjM9AL6/rX5rHk6
1fKzpfLypiwSCLouGPVdtis77WjHP21OFBU4Bp8QFV39knqZZd+5LsyGI0fisoem
fQ0cQQsABDmVOc+9sPzcWukdsm7TIVIarVSuSSU861cIb2buTvYWjslZWvI+NQc8
AX09vbsYvFq1QtA7tUF7H4/2Oxof9+sJyXMltvkf1KsBVA6CD9Ze2bYMdf2te9TV
UisFk0oJIPazMdZUL7llHmqBxGyWD9dA7q/Jst1tzp38wDYwbFZa8IMfSo6mHzWz
PtkMlul9lGhaoNc+bgXQikIBJiTdEa1J0vrpG1So0RdZtJzlKj2Z9iJGyvtSBEgq
rkr/hsKoHHZ+KUh68dKlJ+V6mConSR0NvehgLvVpSARLH2dCK3wMgAI+cyBihXHe
ke/BLM8IBZk2hDf6/mjgFsb6dAiHK/VH7/9lIWvhdd9OJWfY1lACpd92neqwDADC
MQLjJuD6+twc43vxT+ZNT42SohtQUjmsWPV5Dpk+hTJL2vBU48dx4ITaQNnN2bZX
jOhyQjhNUxYWDx0s3CmPm1ALT+wWCGeLTbmOCA35tbQGnPboUEZ+hIYTR9GAsctt
xKdiMQzZ/+JdImFhBQWIMH45YQW2GFXiNNFSOjgrfemw3XaGqT3e3OHPAkNoRKki
DdYSjvRWFMUb7bYQhC84IdfVrlQ+5fHrqOsBxXf8CqwW+7aOhxUgU8Wiqo+5S4so
h7ccmYmOVlCrDoZfJyZjW6V9nLeNqKAl5GVe+Kf092kufPBv0GCeE/viAq4TvRTs
+aW7vbFAVO4c5X6Kh2zMW9QBxnHwu6Hf6oUirCgEx2P66sl0Q2r38jT5deNDo0Td
724dAI72ZzaKmUk7suEIX+XRgmozx6OSnFxL3v0Ou4iKf4pZH5SmkE+vVlutt1Hu
hgX7WpXQiPJmeLqFMOW/F+w8tnbOV8gk7RqXwgtUrv1hu35V+e825bnt57ySdCpj
H5ryd555EiYXOIuW8+aBHcdsDgDyMGx/+YEvB3tYv1/1uGMvWOk3I9raNqrduVlf
FK2vTzH2sP/AtAD4G41T9faFceuFAgWHB5iUQwIpUL1RdlN+O56AVTU/ZhVFbFWq
/HfTbehR3WL9KfcOz37QVuV21CaDbrCaV9zyHN4zpjQO3HSpYKatA68wRv/qy+bz
n8DJvuE++91jc8lFKCJcbwNlZ6UqCYkeR9A7OmiseTXZckfKsGmTt1bb6x3VEUu9
LFT6yOreOVN6k2i7onbdz2NGuDhhpCJ79YdhslGsEKUslaMlcVF+49MQBfgZPGiP
xywY/BjRB6IChwKonRZw6uVlaJ8nCKJKNobufrZ9+LVOqMGiDBf1F7zaVUiE5u2p
nlY5Nw6eYafeVxw5sDMy3HP4C7Se1LiACOQHFIAhAer3li6DCQ0dISf52gknDWyj
/nmQLBqB0up1ZB1zqGjVw/WVJzUFhs/1LIa927lQQ2ZsmBmFoDQt/KiyZNiXVxkg
eIs8fYup/Q9cUD6nrrZxH77pF9rP2Jg+SYCwOPkR37e1RxAb0LfCTslJU/SxcyAF
e45Xx3467hJep88O5dQYJJ/BY8UtK8tfWiEQx2Ip1XpVHPoJoGlvUlkNlgFmycJ+
TPWNV7XV5Wsi8SAgfK8r9B84tDh2kNSvzO6cx7OKMAfE2QlaXHggUmrFW1bHsEi1
Ti9v27HPjMCQiaA4KrIyEYdLfnYT7CZOvR/yRZcU1CHciYs8VzYQ8y9gfTDnnthy
HXxMeV/aRjt2b/jaQmaK6NXkgpaR+g7j1zXgTHyOjiXCUPxRIJgJ9yDXPHf3VI42
iJSMy3ELZlXmr8uqVXEimW4FB6Ir1q5ckg/5Alul12XL63P4do89QMEGCI32BFLc
C6KLsPnCbaJ7GVhws9AOdUZkPjbe6SEVFyfOwXb7Jwh2bgvmsb0dNuye4deyV+Pl
W7sA89uVKmIVSg15IClYMdPsMC7Ox885tg5GNJSFvPjoq4q8XUIgCp9M7UurgrIi
P6TXHKRaJAhwZKMymHgBERDOk8tcjYaWstkPNOT0Armj+WdDwVhUuoyk7wPwGHCy
xCrcSPjqGf5K0J2plhwjBQeQB+87uAwedGVty52eoaYoRtqyhznEdZzCHRGZrd1J
ZG1Px1Mdnf5880RO1kfun3E7eG1XaYUib2LvKfmAczz8svUUSrEd23MOYN+ENae+
U4iXXZ9ixzuJkTXeXR2SzDkgTpFhGygpA45xAbpVDs123XfmCJeJMA/o4uzyoCQ9
4vFrIwuAeDiyfS2SxTCZW4ag4YkLqZmJi0P1qf721ZCTKYlFm3qBQxg/ENrwK7q3
7PuRVcyrSZKn4SjR2ESqRj6pTwbDyp9rnITQFsCGlbDSKc25YlbS7m3ZaptXfEau
fsU/JRYVJ76K5S4meBgUHWEeE25KZC5yyvyuPt3TD+SMdr+2RuXfKEW4fDOUun/3
e54XlivyfC5djI7GDOIlVF6i+ptQnTR5K/RcIAmPaCBjwD+P8GY94OpytVFduxaV
O2peFKp9OxmIe4bQ5mgzUxTinIjycj/54Xxclv7zjWG+sfBHIJynhhr/+VdWEY2X
l12HopFJJCTYY0lf60Zzxxjf5RcfrmVkKArPg+ISW1BAMkY69AURNQGyiBIOqbln
L88DiMcPJsYssTOqQomb7wtzWzAjRXQ37GSTdgBY04I1JZBYua0mGdFN0cl1NB5w
E5ntH6K93YzRKhpq5crwqk7bNRm2LQl9bt1hI8dOaRhOincqjdfZG5/Yw7FxPBTV
yPftBXKN5NSDCAjqBVDkxvpeTx73wzs621uZd0avdqsb51Y0FmIFQGUxQiA8gouR
5Gr2x7mJniKeHkSdJv+uVPLvKpz0gUpJLyUqRSEM6oJ6GT3xAEcUZd/lv2v3n42I
EiwD1WQNf652h3KzF0XY9AocOT8aqexK0Bxqpo7i1yme3UnHKdQDL0XOQON8beEW
fOjt4L1J0+IpaaGY7WN8QsMTsEXFhR63IRyvtzM0DMg8BZwNk3KaowoUMGC2sK1z
KoGEBpIos93OwT5pfjKt/B2kpRVXD5pyiTrz2/5eTgafRBWcI6PCuQ3SQjANfEEC
vprCAxtp6qD/R3Bb9uO4bUNJ92N3U0BVIa1DwbQBaDTTPrPQvBoGGAAe5NqDVzBF
J0beDIrKR+iq0rAjVouSDvSxVbcYif24ipuimIn/xXbhVYRgxq48T0+4Fkvgnsz+
VZ1ZpH5DA1owiQq6w8dLMAJMaqys652g1MYcTsSOeOSqE4ThDtSrCg6A0a9SPUsn
Q+RJsb89JX3FkqhKDMA2CNxGMz4fdMr6Xu8oLkSxbrUgzwVcXyP0nn3Lv0e45B5Z
tNGFuD+dP759G5WfQMUtWwKwFxe2xz2CXPAZykvpfMgFaL0uoJRY1nXghL+5W6D4
qcJd1sxPmaR+JdTYHZfO73Rl1AbYTeQxlRr7mm8fVzlQL/1GsVO8FTyC9pKa6nt2
xbqaLkJFfn/j7i3ZBgNnk/AHYm9JzS93Ym7l4s1dEKXRpFggN+3Ix6LvEoSGGKMk
hHw1O5JmrZN804ikV54TA7gZy4RERdLvfX6X3GGuxRKh7nkIbuclBpe/wHKkMV5e
XLQm0StaVcbPidsSjYtONZ9pTb/QBgLpyCfbkQR8r25XcfOo2eJ39rOb/0GK1zpl
BaQVUACmHJxcy3xxoAteIFPL01GVRkjiBWq6UQhD1s0mHca2OGx1y3wLS9Zf/Xbn
OH8HJqKGA/yLi6ERfIp0uQUJZ4cJlH1Fj0xauIvstq/0acpnWAx2XTTT/K1JkvTD
/7aPruWkjq9mXcQ0X9Ye6QWeoqluEl0T+p4tS1WA85vJ18+FGNc/3pWIj6orZd+Z
Lml5F2Jcwg0yKTwJRqH8KResQifclO4TwPK/yjQGAyViO1I3oqxbMgv8JLo+dGzs
kvoXmuugj67Jrv2USShdE8DTYSSLpsKTxPBN3xPekBF9W0nCCPPRkPJC267ccsj6
Djebpd45srKPJU3AXu2T5MAIXXknOFqw/wV/Ra2kj7TU9mYzYznjdhToPO/L/eWk
d72CY6bT3lesMTHiM81QxdoYAK64+apyBohJcO2YG/UTkGW5U/0/LbxjSfwn3qG0
hS2vvuZNMl9QrS28n5nU54fYKVn17huVmKINOEvC+bfye00llIOAV39j6oseQ6xc
1d4cIMzRocx5pZnjRulgRup3DOcO1/zUEIvsuoWba81ucuYyKeerhz5IhwenOQWw
PhITqeVqjRB91+PEbFcIr4ukCPM9PJrk8XpjX56n33pIZcNpvgKnWEdy8TPJhGCj
V4Qk7ye4gVgzfE/nNnB1U+5lqsKDvFv7zs5cYQ7JC4ckjYJ/y3pjSYoWKk30rdXV
gYhqSodbu2afnm0HCWCBtHazpoYt51NvYIZpwfhfZUVgbEtzKfx32+V8p5touwHj
NBEvTeOunZIoULsIlu+pTISgnU7XuV1o0aKz2EPRSDdb4jve3ls6IL7wVfBOj2MT
INKniKV5hUa8zQcylSOTuX1heysxUn6yEGiFO+4Dl9ccO5l1phzp9TkgN4VNJj3i
0ePw2+25FPIss+EHbMZtbwURRW3rCbFhu2HeT3BfNaWE5DnLWz/o7gasZnnebMAz
2kG6YPzZ4kWQvtvJWCrxEqcxNsbhJvr7H9Vfp/eevCHgxDScVESQxbcyuBXuo8bD
nZW2LNH7Gmk3CXYAv0OGKxZlSgl6HioPLRzAm+C9zV95ci2MZg2B8BrVfiTzZNAG
Ij1QSW5isACLwg30iIr8dGVNi07c0K4z3wwpKFmb5sIlKSzhOogKNgF1KWDe1PI9
CLeGySD7r84f1N1HeX4dkzOsZSPD4KIkxJAOEBpgFpLxMINbhAOxZx2P09cKsXts
nL7r5RLVowPm5rfESPFnRpjGVOR4pPbY4id06notQfsSJxwyjFLsuHNdj2Q6zDZq
yHw0m+fqA+RMgS4kRQYU6Ed6sTlwWDrj5UUkWze67cY3WOwDAed2QVOp0yx3Zv6j
CTxYQ5zg5r70f0+46x9AC6ZoCFzTExpdvJMKgWK/879I4GnPgPybaC9R2iREyYQI
wo6n0tSEiloK/Sl6HLB0R1yMLZFfzPpBl2NOHN+s+QKmeKr8Uwt1SS9KAIAkJvyo
J1MN8/iVPNvU2Dpl6wgDgPo4FVepaBZ2wAhKrcUFrMwGyH2NcfJaBkKeKXx02dtx
kyeaEX7nEAznqGg8uo8df1VfWyIzMMvSCS93UDgeOCd26huSE1p/KywH3UTRMlQr
ofkYPOH5za4DSqbGLu/lIZQIOQ39aUn6qNvznSMRPKzeBtpaoUEjIOBkt3pEccin
im7En5ILmXFt0Usq9Dk1weJW+zOXDCtgv4q9VdPEJJvsS+UK6pBlKPh4rOCQxCFY
+fSjKJVcr9zoxDajQz0fUXd+3YFoyghMBz58V+cpAlSwcwRyF31bMsAffiMv/aEw
0Q6EX3H4MwnQp4fVowJLq2tDnfgfEEQgyHRT5XwlJkTu3AEHSEman/JVidEdoe8Z
UdRSKCvfZyXGcgF8iAUX/ustZxnUpPoS04jeSy980yjNRyEObEE6YBKIHZ7HIe3w
gZxtrpHyrvL6xOUKEiiYeCgBdTbwD7ZBavKYSrRcc+vzlIBKnC2CL2KwoNE3IrU7
UJLOGGPN4VHn8Ut9lp6YCG24xy6HOyRYimIVlDMckUtX7qZEFuEf3UKgRyuRFsEm
eWl2h5cpilHq5wnpQS5LUjqhCpXiSZyYNUoO4HfBmT5KpYpztiLuW/JsxXOvWefW
18Hh/pOao8tw5c4LoBEcIH0badSL7xfB93fvBHpCu7z+AUY77wYOn5LL4Pu2SbdZ
+1TVgeDj5BFCg755z974Fvgmsrf+jCabjIJXTjqqX4I3+5cYL+kIW/EjVWMLpyl2
GhRnu8looye4a9Wt+M84Kzh1oxRxh8ThTIxNoHnwkOCyRannOhta02/fx75jghRx
sv0w/uP4bvr+a3t+1+wvBHUvSsr14JkzsxuicwEVa9tBCneeZE2W71aEE30D57iq
I6xdrpvNZGTlK6PgrJ3KJO28MjLTMr2DnPAjhvBJAxNGJx3NOJm42p7ElyrQe4ku
v9/wtucKdWUnhUXGwTXb7DHzm3r8/Rgf3ixJuvuRiHGcvK/ryT9BzOx0nkqMHJat
tZHVRyV122OWC09CJzDcGD1pVK+/+w6SFBY0JoBWC+doNpIz7A+KeVn0pLyKOg5m
i3Wo5VvW+RUZH5qULsOwrmdJ6u7lqsbfq8sYSb+cmbuQNWG2V0RXrUGL75oadbje
Iowkmr56WnH5xdjCv0+evtF/Ehf3ZsvBYcXgd1jUcCsVMXUZJkPZZUkZQNooIrtn
9iVux0UZQffx8/kqWxLq+dGNNrXmI/HYL2Z6p1sukq1TsnRNjlbA0r0p95+v36Ss
n6Cb01YbKjTuFloB27Zyh7HaWEZlUQ9fCnD8YOUY6GsjY14/tVUZhfahXMQtEsEi
6f0J+Fus0+yLbh29SPfJT+ffO2XAUm6BcGiUd2pGHn4Q2jE6UZQ5nbcVM9pD4Ltz
bd4YhZTLbU+t/VR0gg7MZg/Ozg1RsYT72RNbtfitNVJLlPjFVhqQd+QP0XbHu5wW
1MY2zmtHMeeFkm/fLbNZKBiyQEJwzlOyrk6iFPbXEody2R5DE0gdkcxLMTAM2foM
+/UNFB3xVQ3UTrATS6cTisFb2R3ofQcF1OAjcMWIHNXPmZUQvXlATuCYHBsvVHq1
CGwKJvamCdEYvW62l5GZtXHA10HDB0rDoEzSdfjUK4pF909Pct0FnhPRuXdueEsw
I/JTeLNbuUSw3hpoIQ96ZujDeubqIZebNwMN2i/5VJ6OZs7f5AoWmUjGwPPatfKi
zmszt1e2RqWcu4X3tONOHLueFydC0JlX2zvKdduntI3A38uBTvLBuKoyu93PKt0F
ABPGKd9pQsNPeIw1Dq8+coKidcX3hLL9CMFjh01igKBQePBseZoLQzFEh3TSAGV7
BKNdtl86xCQxfbAhy/CQLfT8tPos++nDcfBXA4rXojhx5O4QQuqrDS1tGg6nSOeG
/5WGpb83NMr1H0h597q8iYXV+RFJtAX9ADtGJDtNEwiT+Ic40bqyXphFLpJVGp3E
QWYHxoZJxMAdeY1r9mkfNlEnAdI5xtCa1kV9no1/5JSVrE/UE8aqc+JUjdwjRJ8p
csaponz9qjV80V5AgrqKy9d/PT0Q/j8dl8rQ/3cKlUDX/YD9mt8ijWqv0OPwYVTr
bPJYEv9dlupM0OHuHs7wItrZOx1IJd8xsw3HHsQrVOWmi4cl3YxisZjF6kCBhUFf
FrFvzuibPlGVp1RoNB3zfs/X2iRsg5EqaiPO49T3qRE5utOTJfFj/bX7crA2aHgi
MvwTQIhqWhDK6cOPSLzMZrj8JplSiah9OyUuEYdFs4UkMob+7tbO1Z8O7tINmL5H
lKl6v1uJvDruhzpEXfYygFmz3/0jmSImj343FcJB+J1SI2GKjv4UKiLA6v6zGGMu
A5zQaCn9gZc8tQDxDogeBB1i5g4WO9tqiFCHcNTEaoO9NHJj2QUtpElrT9XBn7Ly
qqIxz/IHRJEemxefqNaCOoZ1RqOqZqFjqz1q22luFbDi6wxHjy8cil4P7IZNEMR3
tGroWuuJHeBrT30J8wQYusUbUv8t+dTZM3QWPUoKv7aejWIZ/HAdGpVEj5ToF4/U
M/xKSl0vAz53JzRRpc1GTpqVDg5A1s9cMBh/EMckgMq3CUSMu1Ih8VYM7KiiBl9Y
Kg2Sua73RVKRg1JnH2yGkm12jMXClZzAWP13hdTOqxmvUvOAfpLHieYyaRukJDmK
0RSG4x5VLXnKA+J3mViWLodTfoE7rzrqw71BHVLgjkepVoiKcdg6/0IWWBifzq9Z
c6YZ3Y+j9NSdUAg0YJcUMwSPBLZ7aAXqCSOZ2mXrmavfQiIEncx+qXzzVv2yhUu4
E1T+dngWE3uGBMinCyD6TXYTaGvyH2+l7ocP3N+SmCGxHz8eSh0skvZEA+EwIyBy
9h0Gb2NtYK6pEAsuFuzGqWMS0uzTiEfYer86npeqREkWgNjTtKf8/irTCDO8IRgo
wm62k0SZbKb9YXr4kxRupWcoyiG8Fol1FtZsdvNjU2mzC/uXmg7oadjhq2HcW4cg
+5+3MwG8QSYiUa0x/aEZK6zb2XrYIRI0nw6XZHVstp9M/7XjHm/SlfUpsPT4wg6A
JInqDCwzp6qRlY/xpCX+jxLycgzP56LiCy6LBiF6F4gg2COjXp98dg6hpUZkTw3n
oeYB7aRUHpX3jUjvOkWZbFaA79qzVup+KipfCYnzFEwTTHSqVwwZvz3FP5fxLsY3
aeHSoS9FNKVOQNJn8FULQXMVC8+GEwFTh571tyMFTGC8h3pq+RprrkGZi8FH9e0D
7Fx2TAS34mUwkDkB67ktqsuHrP6kxvJUWzQvWZ49GLQztydcDLTQ41tBax7GD8eA
ugUxOJNeM23qXVc4/CsjcZ4h0g8mTrrGB/jdHqQKlK6uy1Rd2xbTslUPKpcteX6X
JvtZUxQkF8QlPNqIEzykhe6GlKy01TV+wQoViEaARHIRNt1x7l225G2+/6I2aaJn
HW8on+jy8UXVixL/NHSTksgPR2L39HtQiLpzApe2XR6Jx2t3LJdveuDpbFqZbnE5
p6RHFOAbi02n9MrP+YrGD1zQQutXna4aWx3T/IA4oCUcisdBUbFFYqTGAdRa0vOK
tFy7D8HFCHgwdOTOQ5nl27goM3fCAXf8DKrLMNdAT5mGPoeBDkPNzYzZyuUTYYvC
nV+sIDOJNT10iEDiT8z4mbikO4K+Hff3F0+vb+ViX0BPC7KfGwrSm3ENKngUvxzw
0d/gItD3kloAWW5hWsKYD4y/U63yYVZA1c2qSyzMBiKXg+lp/7KjLfvTNCFAxCpR
8bU475kN4Ioz+1lgcaOR1WXgAsuCAhLALShwXOnWkvjb19y8TvaO5Hmkf4cAGqaD
e34IKz9PVLfJtznNFv+zhfVcRMP1UeF4wGif1ClSJTpFXXOU63nXu4a7Li8HJOsA
wF/wKM4cS+cLCXaNxEI4tt2G1dBKtYt+pWSvpH4fNU3uGBYTdKHHBYQcSyk2YAvC
JLQmSdFaiciLMuOKihRvcEl678fWzYNme6IXgxhuLoR7ojYPOpH6soheW3o9VH0e
mu2dcvN0h0GKvM0o1ne8R7GIrvPEH4qBxC7QLJL7oBhwX3e524M0mJPhoDhhboo7
JFNuC5vZBE29TNQDl+ym7i90IlCHJ3cYZD3bae16+itD2jjvSPp0ZwT5ohpn80bR
ElN96JztR1KoybOY9rCcbvDHljQoAN40FWllH8ZlojadGuP57powow3FvVKwGlE9
jtQyXaAPKUenvHPm8jNmh0OAXzOexvraqFZmdGwAH3bbmd3Xfaa28peyzak4y68J
Zo32QfjdDwx6cLjU+6PokpsEHlGU6eXWdhbn6A2zWU0AWF7gOuMeGe4JVo8TS2V3
QvBUISUoGXaJY7A1wmYI/1NhByiZ2QwayOfeMfuI7uyLet4PWaklZkIRhV929N3j
IICJi1/q6E5OgY+VJac9L8Mso6/Ck4olX2LfUg6pIpdizceev5cIKSB4blg11bH4
msPGiAlMlQt58bUeukcP0idrnodbIxEPwPkhXKzMBCZlJAXtCO5dRVX4URZ/Utzx
ZV3MpjLLiC5Cs2H5j2CfMMVmf0iSQ49OQfvxSBh3G/xTYZ50vb3oLsJ1VTk5WF45
iN0GcDPH6oW9GHoQ8fa/j7Eg5Ko5H79x3ecwlBvJeLGOANkMwcoWriA/+QTcNGiI
IFobKURsxYZlVcRNExVo4AjBo4n8w1WtVMN9NUlnFdJWyjrWwQj2Uk0nPfSMJZcW
b+Sb5o4RCjAgOM0kvTe5F7yNPTO11O8IUEIPIXZsZtfIri+Q5fdRt6bwSP1X8crl
oEj+AZoe/pLohDuifyWep52ubCQA/Ds3l9Bte5lFQwSvVhR8kdQI//U8h6axzE9S
Fl0jjWF/wa9q1/C4k2Kvo0tenhre13L1eD+89Q3myK09JnAtuDkOqFMlqhJDdmhl
zVbe3hO9Di3aWfML6SNfRdVAOiSe+h/fHMIeq6fi8HLZ3gHPh2TL/o5h5fzkQ+Vv
kJ1Hi9ibzf+C7tGevmnXJCgMphjqLPpJYbnz1aDlcZ5AucxJhYhOTi8XB9+AJFxy
guedYmUXvtovdS1huMLZhjh/5+rMEnaAhBzdau+8L9DDdU4U6+mbAbqGa2P3K/wi
u0VvoA8M+nUUq+4CSNk21zvI/ZtEHgxc3329/ERQ1gDj2yOgqo/SakjmX+KtgG9m
lwNE8wI45ofiJzEi0NpyvlTLMGhGb5mygRN9pzjgM6swg/yfy5N/GUoCUO0DvsX0
9xdqiumO2tJnMperoVph/Gr0J0ov36pcV/u1kLCFFb5ON2xWUJWMIEAKgF92cOvt
30YCzkTsFFWcU4RDF+sFeX2TPQCMYlkaYmQ5mehopqsk1pMwCcbSmdKFTcoPq+l5
K2NvlFmfy8R/2RJwaXONDaXOfXgu0ihciQ0v4jNCJA/LuThcphU9u6P4N0Rn0jpB
tlTN0YxuJTcXPzA2HlaYneFHfKRpCN3yRXwWxuNNGVYGZRFDFVmj/9obJlGTBA3H
QIu+rVqwygwkPNfz6NbyEsrr12xC71Amta+g94fzCrRDUuqDdko48bb5tnbaSAQ8
2KJaOMi4TQQgWThAtgL6zIOv9pbsuq2+voDcSBOo0YpdgYo+xU3AAYC0MwKsv+iB
QkG1D7r9z3WSv1aj6FcO+Q2VUsruMfmyaYqxR/VdHbFdlC5jwPaEVVHZdObnh1nt
5eUBsXVB98143Cr+myutE7nT6ofScytaaLqDZoZjiQLlYiPNNN6TK246f/qdskpX
YyRgXgXxprylgt6jdI6muCb2aDN01o6lY/FTstQ71UW4bgQouZYehzn9sljDSRx0
983CxFpYXiEfQo2ag8NUBWK268DLhawY73Dj6ajZ36dODi8lQDtDfNknhldXK1eW
gCUGyQD5xoWp76ofXUbU9QHQIlvMtB0eDqmT1mOQIe29yFDIu4rwjK9nbn6T2G0R
vw05fhTJoNsk9D4aIM5rZI+Qz9mhEhZMVmBxPMw6sn76tR+OEnrVwLUJtkDW9ZHh
bSEVKc1nYdASOgMTZKe+h/GaNkRCQ3z69COH8ozMdQL0tQXHmbV7K6itponJhk7y
MfM+X/Tjwv75Ai4SdzFa00g2lZOrvG1YwFC6kGksgo6ixo9RdoOsRGz1Tsj7ts/j
bDMjGOv76qjDy7u9en/7S+c01O2gRyuChMVJG9PtTx710LY2V0srchLK3BMcNGU5
k/R/prEysyLp36Anv7Q2ry4Wsh3+10clodsaL4q0/1dB8dn/56A/hd2wqTIgVqFQ
TcChUdoeFI0fMNWmZ3Gvnw/t9qvT3Lhz9QCcKFkxBj/wPvDryfXWaXHMVBAFg/LN
ZnnRyIsB3EoTREk9e1TtwQNP4npcALrERYVR7bBhB35cSXc2Oa0gL9IAIiO0ciga
hyrKdUUheObkqAvrH8RlAd8jOMiTIV+2la6wDoRdOjIPb88rLexXcICqqMIKKo4J
9JukzHXpPD/ERAHOKA0XKXKrIUvvZtPafyeMnV4PvvQs4EGMfu3sWiWoV2w0eNcx
9u2JhpgMfmVsh191o/cOeyEv3o3XqrmaN+kNfU6s57JJmY8fs53QK1AgFo6ZXwXB
c8EjW8T0eJOdUAxtuqg07ez8IiprEm823kBpTUyXHj9HAAeol/UokOth7Aqh9iWh
WjWZc5V3zzbEooCQwoRYSib+41VworbdlzHE7KMXKs2zPfe4pUjYerkI6Y0bL43S
pQ0nlv8narvNtVh6IYUUpCKQI3D1bEniyqvcSaXKRL+RcZlQJENk8PDbUUVhMBJr
27uM05HXdarUKqt8a2CGguxXDVebzbm1R7we6jP80E2c7D+mo5QC8fjbH2tW8bv0
nhxvmKpuP7NJo7IXzpmxfXyPHq7c16CI7XnpXiqouV8OfmDnj6njCjmtktc5VdSD
Di3J6VLlu3TcvLLgjxjgXtc8nYSIeOOlW3e67e+mfMUzDUGasEDg6mHqCLgf7JC6
FunTQTDl+LhqrR0iLQmHOjoOyMuSqp3YNh8Whc67TuCYGRS1GCStDPyKOYMoowIA
yPM1sZmlDGgPhmm/oxWh11QFGKisOxx/7LV8A/24WuKsJil5WfsS3qAc1vGq+4tf
xIg6DkiL0TLZVgZD/NbFNQ4FXmrmcnYQyPlZmvU7LVKZ7sZqhNluhoXAhBpkokkt
wh/cimiKP5LEAbcQwBk4xfGTI08lccHaqSQv8AlJxsNMCIEZhBAzC7ZrIW7HccJU
gfaB/6l8rkRY2HowqgbcHETFas0naf3V3T3XF3YXEk3a/eiQDlb77O2U37n/8cEW
n9kYszmjLN1cdfDj6nDJjqLeICxJqVWj3dRZXZ8b7tzNSFSUSB6XIavQz9YFzBP1
6zPam8AQDuLWNs75uH1WKUxQcxXKRhB4wxq3oQTZLnyAJqaMNptJvKvTAgM/W7KG
HWzDoQ4wld4yMKC1GgfdMsktzGfZocOMw8Spny5gb37mrqaTg7p4ho8MztDrWScU
e72CFCu7+4wWOwPvpn1dlmubk0s3CoNgzFuclCgG4gNRZSdR37t7ZbNQELYnAcKD
npyzvx6Hpz7hxWuwa/yRZHn1zguGUOkxw/x6k54ZarZOOrSV7cE1quk4hTAp5Wxl
4nuRLXH8stLZjxgpKrtSzfsIhc2CwDz5OeDeRZFYUQH3lrQnUjJqn5oJL9OIOH59
FB+douldACYSZFb/B75BkyTPMKnybMQyc+xx7202vX2Q+jnGzAzNJSHuk8pa8jdg
2261ZSW0vgnVjz8crOd8Ikx+QGp7KKQ7sFr7n0YhqYdC7zDQX0OG8bdOW52BBO0L
ceHbFbWwuK/LpyQxc2loND6e23RZKqVgrfr24qpJYFhi2p73Qg1u699L5y2x6wc7
CWcabAN9OUbKuszYJcYANnkznyVAru7OyZXOgXUWf74I7vVIS+lY29cxzPN8EK1E
V3JdBmhuk4+m68wxBvWQJ4khNbMCpLUJUeRixkQbRSP0lYe0kgHmyK8Dz7VRUaIi
rEOJV7ganhR+5sqDf8MI/VjXXOZeuvGgZo5/wcqpx15QdW1OABHhjJW/fZ+VJH5d
RzeDFJnk9+MXfbGqdeMAJMuDDDfjc/2JRTwTaUrqfricjOAIOFni7xL36xr3a2Kn
U4Cqx5YA0S8l+gD9mSS24ioAVzgjv9cVDyhsSB5Ndlki2GdR9i3oieS43feejKoE
9HsXLn0K20zRxU71KoKHdSwNEbO0p/rEPwtTrfJkEBnphV4AOxd74oFjfWCOmK8o
piojJ0CC9qcM11HhwhUY+NCiONg8zXLKvK/S5zL1EpeUFhIRjRfM6kicet7FJCHU
ZVV1KzXWAylp3hZdZCUQWc9hgvGAbpYm5gGWJ7/GBVUrnWnVLaKnoooliqrl5bdQ
3XJuzFCmdx5FBweP3TCAmO4t42JNp+l7gse8Ncn/f9HTnypiw6jHX5b4DDeYTGZj
KJtqRJCWOvJ2zSTCn2sxEqnfkwHx7M0nwKplNTq+YMikbU5gdzwx3ts4Oi5yMhvD
vu7hr9lN7l3URXj+sx8jX2SBznikF3Di2062g/0HK9zXgnNv/41d7H+A8BqfeJpu
Ns5uUwzFHK4rAJqPgdI5Fa8VIT7hvW1WXPpuSCHo8qmnPrP/LDD7k7qn9G0Iwb5G
tklFKuougALspbedldgJsZWrgXHg07mqQcYaVRnlHCdUsLO5BVdK11aD8ZffRlmp
xIdgDT2u5FTQtkcBBFzZQtkcm1MLppJjV9Ei1U0NKAjXQk5mscRFcIuPFqiu1JhO
cqbB9LgkZ46SmPe23CEyPtK8z5m49TWLz5ugGt1FjizUu4zNx9/jDUT2lwMf9yym
T8r81rlj5gGpvehR1jcDts5+jGhAoDr74Oa6oVl/Xw4YIRS2xLu4IAviyqNsvscG
/v+ASCF1xJHcmw4esUg6rzHfKsvRoSf1t3cLwuwPBCknaZm6hzxDkEDVy7Ljbrqu
yf5/sfnRdKPzRRQTBNMzV4TwI7SwfCh1Yusa7MX8NbT2O3nMzABn7v0dtKFWxsfv
H7p6F+C68jEkezrJyP+k+T81C2B/+xQjQo+O5PeZvYodyBjKa96RK9ebtNcubmCy
H/8QT95XW+QWvg2sguMne00at8heb/QIPzPf44c/1gI3W03zXrRpCGJotxsm0piV
Zo14Z2JtDyT4RKGOBmGoaZ/4WUp1AaaDAbBiIvvQxHq1SEQWEpP7LXpM1h+mbRb1
yDMfIk69eH1t/8pzM9mwD8PzqJoVjuvD4lIYSN8KLP4Q4xBLT13GRfrADQhql5G2
n0mXzjZwD6YXfYqt+hyyMtpS3gdsDzVqIwjvefeQyqvaoagzyKq7pkLZeaPvAchK
uwj5G98zd1rZsoY95JggzmXfRjGgG1xp4LibQzM5zviBd/ivgkrJrnDzNyheHYpT
6gaVBbyKi1wN1P8yDVo4qoHAGhs2BuJ9UcyutvZQzwF9pLXOgLWWd3PW4k1gIHRr
MJLU9OM+qAvd6ITfAX/4dxBZfjPTGpIqJPQ8r1mz/3ZjQzh61qIjSaaZqd+9WiNL
qNStEIhAwpjHOATpWooqtVItwhPFhJEuK1RJ8oeek3kRT1pVnRgxZRbE2IOidDyO
/LGtAqw99kDaFAxmokwyOV7zCnJdJPc+GwLWKj5EEHGy/4N4wCwvGbpI6FNu67ze
/FoFazyZG0fb0vk6UQoKZ6P+A29siRArL+TdYarskEQbi0z76ZceCEEm7nd2KV/e
m+oqhr5Whz2R2cx8Oig237UkBFhNeLevbprBTcmsFpoqIc/QLKYVJ9i3E9Z4FV5h
/0e4QPm9xcDXJEoPLD7didK+niifrcRhUY46k+OYHxPrIdB4RL/qXSbfk+ITUZ/h
pxqYRyVhamAHWJWz6yjnAHqkoRtzeOqt8RriVxeK1J+bNinupBQTbPzZrNoMj5Qe
7UDesGNUyrYRsYUiSL3bTH0Sru8Ll/IjCKuAXxwequ0YTIBAiCuf2wI7EAZwgpjd
30Ru2bCVBNy11vR3/nSfrOgfsygeKzCdmXFDvs0NHM1xbAPTbTWExuHFiNB9FFx/
OsVC02+Rf4/m9xwtxiqVzz5i9RPvpzKqfQg1m1A3DcgXc/Li9gv8zGJtVBcJQlM4
VOAoXFU/7R3whI+QUjsFqxyc86Cno5xYH0cy7srgvPDGJVBpnX4vLICryZ511qGy
nT2PI0n9WjqFuoG7hWT+B7FA0V6E+kvBt5Rszr4UMKrIuMr5AM2XM3BA5pXntxDg
MtqzBarDqllomPejwSx07jGFBe4QHBsDrunTdnmrM1gICOirZfk4RdEbRirrrV/E
8W5VbcZ4Av1inVEVzbMi6+idcwwnnveAZdAoR5y2i9feZw8agXpys8fm7iJpaxLi
VhPx1PZcKTNppAs0y/XYv3CgTt++iDzC0+MZc79Bo9V7pN6MdXDhnLiKxlgnRtBJ
NbOcIP/aHnT/N1JLUQ6WHu6mzpNYtG15n9Iz7PD83m2bvvxlilm1Uljk6ysfFYCY
21TgPnAzU8nK18FrljTiApcJiy6rW+5aHeZJEtiRik2aDAhSnZ1OhvBijdnsS86A
aa9kFxoN7GGdzda+YmzTZC9D6OBek7+Fyew0K25Y21SnQeL6HKtal9u7n67vOgHU
2vwDHWDg6fY/c0hrya6GSrHTBIBpLnJtZmhe2bsLzcAyItIBQDb+rHMOTgMFKfHu
aR4oWn9qPeLnQWY719OvoW2j0nqwhJkU1L+13F5y43UY6v6sLmsGfzGAmVRBdlS1
RKalMHCs0MIyISKrvuo9gJRSaxgslKDqoTcGn8JKRniyPAiM2JnULCOueaqhZdzB
OQWwiypYzS6gNrlLXmLgHXpyI4a/hqGLxDft5rIDEWM9w8sc+9g46vFe0DR1yLgY
hFD8kBWgOQMYNIdGjAYlUmx/BAu6P2+EAnn8looQp+X2buYrTG4EG2Vwnb+MW1Na
xDuUctKxX3jb/CxT0CG1hdZzrMGZ0O3e3cZVI5hy0eJzdTmaxc6O4X+EUR/ViEUL
4cUhMSjOk9uyjlTEeyNuhxOfwcA9bj/IZZECIS40Na2KzypXTfQHVoz0LgdxrVBF
A2ApR62uDG39+tb9kaL3jsfjTVajKkQ20+6MtIsmfay6I74PX1b2KxD/Y4qq33Jk
4fWC1GHy/V4us0z9nFnleEZQT2U36kCqhbx50iY0lslUQuCcM66BFrVCUb1zfgKJ
qAXa73ITfMV9wnhewoSgOnXJtwYjcutyCX00Ln4ZpKw5OD2Yp/2Ee5zwKUTS0VhQ
MtRu6yet/F2e/WByLmgLbZtWsesPCdhIm15K3vznChtl2A0nPzpNUQqGUw0H43hY
SrJA/wcDrOfq55i7kLfG0blXNWrheUzepxgxaZKdhpVpLijb6WTILNpfLpdZqSL6
TQZ1tI0pMBYE2HA/Z6SMgh8gpc20MKQxBkp1gpqE54YVsct8jXJQrAxMcnZcauL5
wIUhMYhCtNob3Gzo5z+lqorqa8lb1GD/6VOLvcE+L/8mNrt9qeuo3oqYIdAjFKZa
jbY+00mf/WseqDvTmTIw43b/fqYcwMopBbwGBmWaFFIbhOp+G31tQSi4aBMogwKm
6Ez8nNK+n/U1KRPFSs8y5w1IEAwLTem8aB2pAOKcS7jNOuA/1BXPLMljvbkUffIu
B2BIKzc/PYkIS/Y0bFydmNzf+DPYkj31XncUWEpeCJdSnbv0cCLmWpvo5mq6/Q8g
q8Dzex8es2T8xCNdmevl0ad9HxL6Org7lwJ3kBs6LwTWOyw1Zi8JeveRi4n8TUU5
LYJJJwqtexICbgZzZMj+aty4U6VDDcnk1JAvgW5QeC+vJ//XLvJaBvpfB074IqXf
d8moDiJ3L/y4pWeAvlZLu6mkWiAvDWISYGv3FvZ+9Ly0tSx1Tppsf+3nWZxMclCn
/TA0wjwdNcFoDkC6mbG25HErLg/sDoTkzEOhyx7VhMO/0xJNxWTGmdkzBjqzB7iB
mzcSshWk6z7vxsMgj3Q8nfSIaNwqqC56JTtSuiGFgPd5wO/82LVCtLdofzVkHp1s
Eb8EGov64Qn7ZeHsV68O740f5AuZFDIxXfMhLJQafSIf1uQEMOpmkKIfiOrRvLgW
7dCTfZolrL+VomR78+flkgO3xVwTdtfKEomgnEZflXKrQX3ACAYVPoKfzvGXRoky
zzSOY/QBPyiFDMIGnykf/J7aDPV851wgzL/hKoB2C2+hx7ERHOJ85SGi5ViMKUVX
EL4c81AKPEre7pjFjQqTDWjMiXqvPKMVGfs1H4d2Pg5GHDZM7g9f1DBlx11xIXJs
Ch4KeNw3KqAsZijzLhGj2UJlBiFn9GCbtzhA6Yos7BbMKuNjm+JhgLCbHIP26Vzm
c1kdCnNPebHkbxHxSGDFEOwVdOB1Q935u3CQUuf6zpBNDFn/rWjxaTD26HRn8uDV
KJGXRu/TMmhNejxuQ6rjO1hxHAQmj/9XzmynHQ0cPR+/R5gokakrDKQLwMCaD2YT
aK+QexeW3H4V8pgrw2Wyrk/8GEtwwqQC/ye+i8Mv2Zof0dSJ4O1hPFdpdJqO7TmY
nzL1WCn4gXfDRr4Wi84+IRc/2Ko7kUL64hn4QGlHjGkI4LwWZKZLyPA9UPHlzl4q
gfYgvFIjiaAYuBAICsF1E5pqRQAFa2ZO+C3srTSj0O5Iza54W2Do9h7qzrMGCheN
QnecVNRXzhMWEBiYn3XW8LurSCeI61Ow/kjmKPxw7CtUbhkzNfVAj2DtbNGmE+0N
WuP3Uq0wiy7B6Nw4NeQwCUstTKS6uHdPNoJvSeQoyjBridXS8BYWcZeYFGPyk25X
Z8Aq9mFHu7fAjXhYDpjtIEJ03h7dubSRGZW+dmHtI6PbS4lnwPtITu5xJe/4Erhr
k4KgKK+WhtsEfiNdODz5fnM/gqEfkdjP+RjYtxBduVe/7ANSeMOh0EpTVbR/qSxQ
NsHzIc3G16VFbhAjc8c9aVWXD7fVvjKfY9wpbd6aQWm1+b+k2GLKKmr+VxyFe0t+
bAeNA4CG2T3s7QA2EQVps3nli5cVk8RP4I3WBnpDxd+JDFGtM/pYu3cYyS0nsV9t
jd84psFiJqu+UDSn0PLcWIYl+OL5RlWxgGjC3V756iynuL9HviXpxbX9yaJDc7IM
Bk0n07vdkMtLnitGPnOSNWhuff8vraNOc8Ro0SqFoKCR9Q4e6oJfzudCU1vXWTp/
AA7TxbvyAsFlnTdyFpsCCceI+QHMmVj1AC9VX+7/8NV4+kJ3+x1Y9JHB2ju5iLp2
oqZHZYxM/THSKTpxFRGOuyNWX7Qm/mGlVcVYyea4mg2BRivOOa30n2Z0nbVxH58G
VWPdC+wToaykGm9C9e+vPESlnGK7E1vMY1FvotsgDGC+grKvN2K4vWMnbt38Joyh
f5vzdEoD8ecVjQ2P1MJOwE2LOMipdAoGjn59lrSXBoWeXHUgFQGRClWDp7pK2+SH
HupmJ7MMj1ucm0ygdMNWrJI6rANKS67LGWsmCWOoxeMpnr4ULtzHakyuvHdL8GXh
IMkVmBfZUmAFxlvk+Z34hJRdTqVaQDPLZpbmcbpFIjAuUDt8sD5tYgpphfMLPY+N
QWkuRpJfH41tE5Q4yRruAUX+NWQu/x2zCloqGD0j9FGMVvqzTOBG3ZScrXqKOPMZ
BxWoTIMlOwxSoTZxlpxqBjM5mR6lYzKBZwRleDW1SJQFburNb8A6MbOeJDrduRCc
/IjATZ4oZoxCU9H7Zbq02Z0ntTDTivl0JtAixxDMG01mPAOx+yxK/tMEO1BH3Bd2
MHcNMia+yj0lAAEGk+n4cD5fz5uk1O1ADcgKifis/yOPlPCWgA0Nc1rJeZO8N9u3
P8xyS71UTx29/V16KcJwvBNSGm472uhMvtDMYrlRKai7PSVNpavdY65ZDkoOkdHE
pnkIs6egLBcW6qubC/wqrYoqRZZBiJRprYH6mAezH9vHuXCfNV5MatRAnIhsFmrE
d1u4TtJliuG72YxOfVorQKaQ7ADn8r/zVZjZOZi4iyvRZggqmv3fILgYR2yER0iZ
qiHCVb3WPo+l8zJ4YWu9XPqfaNYeRrg+pOviA0UR3aChHqReXgriSirqmIhKNq08
yC85rqnI06CALBTH32xDJzMyrI1+AKPzjBbxTfLyBk73CASEsWy0y9VVf+xkEkML
C8j116pW9lR0IMFM1Ew9dq6OhaaQlPhC7bbAyWyV+hm8bUIkkGbP39oepOb4J47y
S/aTDg7Hi1Y9HeFgpAb12+XUYPJpaNwppVXGAKAw8+1g8K+mCrfIyC97VUWbThpi
w0FqwIsiVVzATkmpGMZ9+Dv2Izbm4MIM10IMhE/Lhdgd1r1WhMPtFfXk5GItFGLb
WEFcC+pVcYDjb9Av3etVA07V3iRzP0GlTjC53ylCSE74e5vGfwZnmSRlvyBO0a4b
xJaDLPL//JMKmEIIBNyA+SdJoKbkciNfmEREEb5+anbQmY0bQQWbl8X1qelMxKy5
2XlNNqrWuHxdjubOd8ZUq8GlttdbxylFYP6EQF4QakIrrK1Ck7f1YKtIB2X/pbs7
XyAmEXG2SiOho/HuzvPIBiVhZLQ0TB4zVumJ1nPCxULiWxm2V3M1wL/Knbccl46u
ZHxIsRLdVuAMRjNSlnQfKHdJfeap3kpexs2OEdgYAi8DHJaYDROJs2LPVWzsLN+1
OD/tnXXRMUbRCbpESun1n7esvk1lYdASmLiT0U+p6C6mnHFKRoMveBuYm42LQxxB
j77Ax1Yc0+Zfr1IDbQptjG34i6rbsOuxTBqb8V67c2wH3hnS8TVBUOF1KeVvC4tq
1RuQkbc50Km9rA2BxBzuYzU0PzdozPTyzrfq7RSBWSWuU+Z8DZzPPWw+/Z5QuchZ
h5mdJtNkiE3L1E22L7yyKz271XtD13V8gyEEqixwctUGj9s8dmf0iL9Yv3SHJrXH
2mn4nuidkzWVNk6zDKp5SgTVLqpzAr79iNBzW/K0LTg1GAUTYhvXgdMvIQ1BGm51
9x1PYWZRbBeSNWAtJpOlZQJ+yo3wOw1XpanxyHuN9+l1XODIwgi/HDSRBB63ZAU2
M5uCTG9w+0+RQtA8ChQCAC2C1mB7HH170mJ6riLJyWM8muI5P0ANjWk3/mJiMpWw
OMOGHys7DCZfsXznhL93bbI/FuFkAfAb62mGTyx9bjmWemVyfY7AzdbzdIy20nHw
fiiBdCnXYuXkUaZRk4JeZ6x6RS79z0KO9QW2pSl46HUnIGZsbZD2jHrq98T7eQQn
zio80uAEQVC3tnzeg69Caw9yyS2LNMQBo8prx+jN4eb4AG4Opk/9vKfNgQGA/a3+
zAgOpIfmkY1JaUJoOpYsRnlworygARXqW7jGOBImcdjXYca6UX96IcsLATMlIfnL
C2UFT9wcITerdHC0l8haTnVGlKQdpweERD35IJkc5wFtkw2KeYWHr0eZ6yb2tTU3
v0X7K+ya9zNEY+5jUi6kKC0prVmLOa7hIsYCRh3XhVxkzWpolnXI0EwMyZ6ZoRWa
gp4UpmRIIlzXMBj2WelAAL4a9qhv4g4NjmpRx4/QRRk5jqfLW0+mLqN1aSI72e7F
24gEuBFLNzieshRM/6G+d8Gu4VRM/sGs9PWDO7Db1f2KCw8ZGSee2e+uUGtB/dYP
NppBNBfC0nFy4b3nD9Es9BeQNM8rQqmgB+PdSjWE4RXQ7FezRkamQBA9dnkdj1Fp
XXdI9zXUuZlkrP3eBcIzUPEsDh+w2Zky5lcdnIE/ggqXfgk9bhgFVD0lzCtPN6kS
DMiZiw1BVFa+16bAQEJXnHKU6RUwUlI//5jVafdGd7mk+bv73Da49A7Q/EQDm/FW
wDpk+JVjWgJu5VDSDrP+ABrzWdpcZXiJEYkhNo/7G0QdTcs4gWkxI5q3nI2GOBOh
UHvykApQhaUpFMIRWTl0fSD5KKaytoIWhMMFvAoFHPRJvfbr2T4vUu5ICEz9ORlz
Scs4SnC2Ce1Nr5kX2rP1tms7KuzFOM/mqTELvYOAuoiYRMZl2EIXw0rRKi5xJShq
HJszWRq7ooFq1UGBbER7hU3XL1NYlzVZZ5WUJE3T0glDpdDKQgLSZm4akFUoUKtw
3/LCdJ0gjbYA7EFhjhjaoUedJ0oe86rn9e9T9RIVtzXlCYfOEV2OiuttAodHKeFM
nQzDq/QbJL8ULmhiSxeoGXhyloIOfCmbpasiKw4WjvkaAa9QG+zLUY3If2sJpNmb
JClBISJsENZcec3A/OVCgcsVuQoMqLzDhs4SMMmhiGUIvM1YndtLcyIpEz1M+9uD
u7N6VvQZchYoZFap5MHRLftY/tIkS3pv7z12mbqICbGTXtjXScNFDNK+NEBcMpbe
zyzf0IyPIf0XhIFMu3xsBpdQ/LT+x0TKj1poK8c0gTZClCwIyyzn2R5OwChgcUFs
tgCEw2WJghjmTCWW08ghpMrgZuQYyQgFiacBn9YLE1EGlB151cCN403xFFy2IPIL
4A++z4GnXiGwoaD3aLOUJ6bXkwQH4y2b/sS6f5Lflc3C1xYD6AE0rDdlWrUwL89u
4O+x8gwzAAprapisDmJ+We/MF36c2dcSioGNT9N/yb+psZY+7Z/E9PoH8QtVgGDQ
wfRHDW7ginRq5oDIpB0K5WsPwKv5RqsZbko2g6zQpCFIVE+XvLJZHmR8NHa3tr6c
cpv8H/rZUk7MITd1k5zW78xY+c9d8+BIOPP664n4jZsPPtxfCJ1wl7WzthsGzxmJ
pBtnvQlxBjJEU8X38dUvg+ll28JZbXK+bv+pnzMEpjVnWJY+Wceq9uJLeWtKYt1W
qGuxzKjouVgQmYvMaiK9IJIvZW6RL0xKcpkLht2lWenEv1IxC77041csh4s73/pB
hukSCKEYtghlUuiqpLmpr8rDLZN4037TiXIravGTZcwbrZplVbTUieuZnScc5tfV
bjcBnHQ2xXzAybk5VKCmTTZKd8Js/LW7KES3mcYSX/1SuUZBax9VEri+uz/aIshp
0KJqg9WQT1OWl6z+OvHXPEWbFfhMEv1N318Qnau1l04YGRnoMGDkyWN5SHBqpL6S
dLK5pffaSiXJEDf9fiYnaVCg086pQuu0cVV6eDvRpzbiiw87nNpAMq/5D9JIeBKv
vWuQzeB2gGBixAx+SPMmvGeKBJ/Y0LOKLeL2q7DHJ0/VKYXLqvq22SkuWU1FpzQU
mbN5egPnDrE+iPXxq2+slsI63IBIIvWVl7EBCzjTjW1k2TaocEi4Aqb8pAuP+jz9
SdRq44mBdgHrQ+Vn20uevOD96kg7ZaV8npqhElHkTm44SI3Vg6sc0+70T8DSKcmq
EJHlwRW92YxjosZXWMMo7OfzWgKPDhcgnoJzOsJEkKTDFZm+1O6WNR4w4VKWKwn5
5a0rsI1OK3WNbS3Mq5f53MTu62eRay8kDaMnTMdW+YJ5bQg8pdSOZY2DMlPp0SnW
jEx48ydgeN+Ox18cU78TK7HMah+Q1QqpeaPQ7X15qbkj8gNV73qfZb4ZwYaV+CrC
nNnRAqy7OEm93Vd3uaaA+7zyGvkmnhoE3LJo8Xui+b2A7Lb54fZEq59ySBrBCBsb
FkP8Rl1t2h/1EC1DGXCCzXxXFy21g+Lh3SK/rdm8PuxbtzE14QDuHbqyTjzfzgo9
2IGsnREp1wnUA7VyVYv/GxptAa5kGtYMFFwjTXGHje7yWhvyTbqPZM86o+MKhdV9
91UjPhTWzizoufbyMaIJU9YAw7EJPEXGLmVa8sjH7bh6YcN7BPOj2093ZopY6Qn7
ATKFhl9qDM7SBx1Jre21BhLxesuMo5L0HCr6d4veOGvnl/7f5aZDBk3ob+Es6hDj
FEE9qOL+MpvZ0beOB7uN1gGQokpeFIocpGfTs4bwHbSVdxiiZQqdCcju1NxEDIkb
J74KfcrDkAVkZzncGqwR74Fox1UmYnXQEDIkOBZ96CvwGNdhI23h3y+bbhMruPyJ
rVGLcdvtnc38IJPN1islQcWgkZOHYoqjnWJ5m5WOagqQK/46W+/rSW067zOqVEpf
gcLmX2IYgI5f1PtoQSD4xO5fUxPH7zc5r0joFmi8NV/oEoOFf7yvepibY7cnSC9g
wN+R75CQTghfHT0be1VqZT0w7KDLyFq5Eberg6JNVnDVkzn76tFjd4AVnpcnaipN
rOUzFypQB1zCaIu5Lw2lfhReQ9Vh8SA3fVaOZDH+TUVzJf4h8eWtq7IZ+MNMMblL
G1QoBUq38NUF21c4W0nWQrQ0nePZkhRWMT6G8/kiwkQ+nHxxWOLUsCsZhnxSCEbt
j0nW+WER5aKNSHvasnypNfeLvn7UlVPpufbCZVN9xjWhVSwK3ojQ6uO0Z+3C/BL8
UsvCcemf7YvELQHrPKJ6vZ6p1ZpAVQVonYOR2FewlrrmkHRFcD+2jGp/6xC+68mN
DzdvFQknlcQoU87Tbw2UmPvWOifIGcvtpWiX/x7IE0wG5gONOExaYbwddVZW1Jbw
4XnFslS+7lHIMnoKke+w7xGDHypi8IT9nYm2WrbOvC6rOGrjigU08fbr5TWPPFw9
lbkXmk1oMTz+Lygr06ArxLj8xcLoiGXuapzJwhcLAA4mvjxUvw47n+/LuFmHX/YK
T9SG3N2Uff0y0tk76VfZZm/vRfo3SxJ2eX3r3seXZYkyX6uZ2OC3VdEN4QFF+P1w
FXvxqG8MBGQ0DcvDMdjHm8RDMobOON44AYfhG/5aqUidxTVynpf7dDL3VOn0I5hP
RSobV79VnHsJFPMuJja7f/xeQ8HHRfSJ78D7f7GRT3mMyggJaX9wG9tdir0qwTiD
hRRUg7UBuwWioxK9+6e+F/T2p7dtPPc7EOw5ztXyl6CSqyQB9KX2HhSbfJuUgbCS
WigTakSBV+8SCUbYEyy8eKqd368R3goSwjpugZGYE5kGtIO1dTDgwwq7Ya4dj7Fe
68avgVwz/eIYKcVo7jc9yIe9rsBglp5XCgH4HuBbuLzb+8ApZgYDizLAq0yOqJfN
Paxpvm5tF0qGVxsbCvHDEWz1F67F2kOemJtHV1+TjqLIiEsNtbR74n0RSb++TFUW
KbJrVTEqNqdJH+Kizi3MxZAAR1xoURxUfw3QXz8OcyzfvqE1F9sVBBLEVgGUruLk
EOZ05X4n9GgqmzADczDeYhhh8FSOYNiAcDJ6HsiV4PGeujO1voHkwYgqJDeJ/edn
3fF3dnrzv+ivatWBWYs2BvjFrEiAMiKtH8z60Js/IgfJRRLL6yjgQQWYbfM3OOjA
poC10nzK5hUiEbhRmpOoVTDenCH7hmuqHLJL6kqPWry4t5HUUrxn9oKLjFBdvY6a
rF+7ItKRjZIcYRb35vfvddo1BZ3ohG0mFgqcjEQ65aDAXXut6qaPs5s1T3+TyzQh
LCkEvywxgRt82xtUK0BikSGFDg8otR37hutX+JxY2C8yDND7vyU1HQV+Hw54/ofl
OfTpSD2bjEIf5Gdbnfqy00lLkiwBz5bJaTBAcvX/ln+CRQX0r9FkyAexTH3skvEg
ZDMt86rn2NYQHlvQI6PezOfRkym/ZwLnriD2FcR51eoq10bqETfcLf3C2hUfTeiW
XuZEOrgBHJDelJvJLcfk9w5qLcVg6RdnHaNWgTplxxPyBKcQ4S0u3EK/f6I87oXb
mVLR5K3mAhGMT5xwZgnS8E5EfGV4NzS8mCbIlQTKCzyb6IxEB/6ZXkTQQN4CwKlI
ex8DE9zyyaSFHILboYrp3bVl3EPzJ8CaAEjjRFRNXEza0VfECNhJTP5Hw/fi+jvU
bXchEseZR7hJTT8d4gyZc5+XBQok2JjWW6wbQ9V+ITzHJxM/L3y6/F2d2MZxqATP
IBE22yphg8EyX/EK6aHnaGIi6yC7Ou8N2p7NglbaAXwg1+dzKND1+Zw26dZsIcDu
KRcHzDkglVV097O48lqT6njkaLsKc/luvwuP3nUSjsFAKm3jzpThGWjrs/RfigAe
OXTADSiu2gGthAbBPyy2VLXBTF78fbWmQqQVokx7FzP4ksf462LZlT0t1GJGqvoz
khnPCodm53srU7p6h5F3YuI+T704/sTzhhN8BQvzx2SsvBLb47K1JFjwx6Vfj5B3
5gTm4svGIjgMugH0ggWrQnJWc3TcAiwuWKNK6I47Rx8hVKPlrOdO1psxFDHCQNFc
6jxLVgzKoJ4TiPV4vPcYcIczdaduOTOtSp6sP2R3mvALU8LdZUrBq0v6POpQQxeH
whBZ3GgVT4xBENxMIYa36IckywCHgfFssbt2BiYxkZ1LHXG/FRNb/vx8SijC0oTS
UxicBsoVP9CC5rFNuv4XjTO8Ci6BK/gi96mtccSbCdH8HW/RDIPv8nP4EBGTJEEz
qR9YbmaLw21+YPQPqccfcuykX2AZ4FJ0TJNzaq03AlNdzL7tJrKqTL8CO9IPpkZ/
KC9Q4YtvzlD+7/fk635PUZ27B/tXnYE6UOK/Wm94jYb1JidrJaZoMN5jhyqDU/8e
LUNk6QpsU5sGl8jLXYVRRLBSqHMmD5N5kG1HTZNtefPS4ob3rGKuWwns+c9HpJFp
ITwUfaWfW3OlCJA59bB+DGS3xJvkhB4c2BIlcmCJyyPEO1sM7dCfHQSe/yVbs0zr
8qVDgPVlZlZvCB93NE4Gd0DmPbzyGKrb/rtHbmdSY/+wPhThtb8yJ6S8CE0hafJD
aS6KLFQdbP2naLrq+h1bZlK8Num6lu1NmxYU4iET9v6BOzVWFNAAj8noRUfMqM91
hFwlPdjzi47VGLTxRcuEE9vVq6zCUyDgUU0iOMEnunxIZjrK4YqUb4ED5EpQWmtb
aD3LhB3qJl/uCELaD+rI8Ndh708PFGC6p/DfjN7Id19LyqqpHKKl6sGGI7IGyQCp
NSrDqfPT/XNdhC5ybVl76D+CGV//TDDYKhULdJbZw+cGud1ud9gAYIJVMXeGwviT
3nF2BaZjzlb7ybAduhoF2TfA0yVHwkKH4FMsG7/3q7EHjGew1YrlzpwJRAKfFp01
c8WdZCSBEqHI22VvLThQPt9i5L6/P7BUGXLkt+v7fKcoEkeS4Xfm0Fe8ij6VTVIn
uCzuyB+xV2GnmXKDpijcjIxPi6EoBv1qT9R+5yrqpKOA4/ncUhXbza0o/Mbj8eMQ
BM2E1VP49YoiXku3J3g8lLDjDqmRPtWufNucB07HrSlwb3iU0pO98h9T7YXH0JWI
pGGAp1f/NkpPlRW78ZY5gpcg6Y2ioKJBX1lCEAAjRhv1TeEjcjTOCL9RvErrEBSj
SWu488ozgN4i/ZnvW6aV/fAjePPbjHTLrlKq5oXN3CHWeBLRRXLtG/cOxQO6vxq2
2mCQXFV/H9u54fgZhONv6nvwwJDqZvmAMvMAdwxh92MPx68xAbm1lVOti5QHVllo
7kPW/DFkS85cwlAiuYiyE+KoVgXnchCZx1x00OwhmAIAEfyfTNTQDwHvnybd9OSc
E7BHWJ3h3UvmT6Um/K1vsOVQ/BWnLgwWlxmkC4rk0xr7c5DzRCvUHaJBONqh2wE3
AjAwPp0WWxTl9h/4wnBoUv3KTOMumnN2drcl2DyBlUo96JAh208rBBXm2QNcIcuN
vPQR9uLc8xRTRlhQAxjBsp18RedJNEKuNVPBC+VEnMzTNtHswz0DyySfSaXnz3CI
z+8VIR57VaN46rCKbSAH0GCK0BHOO3xYfrGGN14/1qxl6vq9qOpNi3IX46E+prBg
RMHg3BWzpg0+crEFyjNYu86EiIiDSnroySjcZFgbU73kVh0HkIkyLPKcNrABn2PZ
RjR3hkhRHLlNZNt7/eDTh9Frgl7EdsENjxXrUlM/8f49t5Gx1DlcdM8QIMk7vlSW
++Bysb90UPkr4Gse3HSinW+1vGXkyLwAasuJ1Qapeyai7yXrejHZNQDwMLJl+Lft
+4fUe3qdAUkNXl/GryImd+5D4Fb9FmcXpN00fwBX5z4wPpn/b+/CTpn8J9WhDP1b
yETT9as4Duj8q2v6thZEHG4tkCPO+IdqgFYMIy4mmA4V3g65gML8t6/j9EYlg+p0
uQvBQSzx72JCsF6vk/xCAI6ZsJVnDTnBJSWMtLu095nQ1tSsBRNe47NZHuvEoa09
vrgNjZ5AEyZwbpQdSMILb4HscajirdMCKo+Nvj9cDtPpflTYo+d7/wtQLv3Vferv
bTDLKV2MYg5tp/0G5HY93oPAfQnhr/K/yNPU1IyZ5keB1EBSyyQhDfOHmwKIb1TV
nYr7Wo2dyafLXjYYV4xSzf2yPNoWEiQt+WVRdIyH5W/EoGNwmzvs1sdLGIzIxPbF
Mi7Pw0//IIwl2osGcM304CTu3jPK5tiGu1ivyLPZlOv1747ugHtYAfZvO7wfgJ2a
Udhh9x3UzaV8kOs2XyLbrjo6OTHXqp2jELXHlZ+L8+1HsS6ldyQLmFQgXDm3wUd1
8uj9wpANDtrO99lEw9hAsS7hRZHTkgnpN3/jSXw99jGHkCsQ+zcWkGzcNc4o5U+J
0BC4j1DFCjRh56OOhfQj9PJgRiyNPhtlKZVIs6ySoRIDell+KZ3sUsEsk/j/CMS9
wn+i3Gclj8bBH7/LC20EksfU3hsRQHJMUp3m9NukIhFfv7rkJF6VFhyEZwKIGc+V
7Cdvkmr0GHTkD7Dp79mNT79tk6T7UWoxLUMfXdKUJNQNF98yy84odIkRJxhmyKaC
D3uQdoQhlEZupvPTt99CO5otX02h3iXKhF/3VAhJHmElvcti3KdwiwIslj5ImJ6b
RYRq3UwjqFmHIaoSPPij1K65V2JMw/GPJYUKS/Uw+o1t6ud3cmOsXlG4h2Z6unUh
VNyUNwPSFR0tH5CnwtmOil0TUohtGss/SioDH+eT4f7PpYqiIjzGTvf3pC2+DfU3
ql4zIrMVjEJNqSM3YkBdXkJx8HE7p/WPQvMGQvVniHNnIySyIC2Ue/iGG2HLnDfz
xrb5h6BnYINYD4S5gHkghtAqacBkA8hdQVUMeEKae2S8z3cD7q6EzaKT0gWe1QPD
giSLTeZedrt4GIuvP71aAvN05E+bcSacspAHq+C4TJvuKIwAhH93xR7wrwZzMW/K
rFP1hJiM7qq5VOR4289wRdq/5lFmurHqZd6fW9fHPq2GeWT9B3GIi3BSgp6PQXiz
jzkuxp4+Cix2rfn//g9Req46xsXweIVdUhkC6HyAAFJ70SqMnMcjfGOAV7L2qkam
W+1NxGCvGAyEitoUYOZz+jwnjhM/Ex6ZFdPn/qRojroX6qM06uP1fb3gC8xWfgLu
OcdBFwFtHbIwG9ojmKc22mTxVcUf8rIJl/jJcKcfllX1vn6cWABFjFzqfbpAfIJF
P/qGIZQz7avTcGnJ1AulpdzQGEHBLfAB4vg+uETsJT7t8JSJtE2ovZnYAFXCa4/X
NfJjI4FMFiMxnLlLQISK7SDw3YLqBbu8iVv9Zzan6Td8YuJGCpL4jm6bAsugykfw
B82g/gwqDHIngl6yHI/yN//zG0bMqfKw6IgIqPsGRZBdSdIV+roVpLB9HjhwvJ1X
cJjul3J/20ODIkOkum9k/1rtQUe/r2vyTdn1aMIEj+qfnHGOgFiH+7gpN+puH6t9
i0PTs3vsjmvnLEZc5hZbiD4ENRvBLEmyz9lU76qv7h4uFnvO29wI3yeoxgzD6Czc
OIrG/KrNIIk1vn4AC1N4wJtp4OMG/dO1pdaeSxZaG3D+hLj1OsJWjLt4a6hfaBUw
1uUmVqNXYxq6rwlb1aDEneM6Jdl3EGnFHVUN0PQDdYP7XbO7okA6mAN1FgvLEV0z
7v9DI9L5l5ONhvJ+OEcoyVwS53naFCJHyicfxjd2ne2K0kN9Rpnp6bIbsn85ANRo
/xlU+4Z0tBbdfxNoftE5DPPRSYTzPaOzNroBUy5n0RrPMk+5JQWFhgnGrjAkpYRO
UTXTL8cDHHVAaSUMeois7ugxvxg0fgoYq4Ce28wYHfMmc1Yv/M7SFlzFQTdaG2XA
hvYbrTwBRB+PhPSKIQtSlyyZUEgkYWanM/HflZpyxd96iY5qo2HzcxBxB5HYIqKs
Y0gJIV8iR4R/zi7DmBxeq1TAawwBAzhnEZSY0eQFHJVohk2kkk+1hbq5wzyuQqwc
2G2MkGrbmkqAfNbxUMHRQrIu97Wpv/Gu6bB7O+B2DJUD6Ycb1fOImR0G86V51V+D
3K8ox5VhSgjvZcP0vmdm4Ba3hkDNSpmR1HgcXGNgfN5/StoQcTFQDXHV4IgJVOFD
BES0xPH+QFu78YFk1PTPleuQLIG6oZV7ZVzTG6C5DoIuLyPBr5j6DWKEc+2sfzGi
gLPonqmFlxQcoMEQh/Qcdcq3c6umzaD2BfBlwDS5mS80tTu8CByLAV7YIoGImnWV
DiKRTQE6DrpLtVp+ijhrc0+bmtX2Byv3qDUXCsuvlrl9IPfK0NFl3j72HR5Ye46Y
d93VY09im5Otc9IeXcf5nXlYLDUDQPWUPqECE7NcqtQnzd2VoE1TfXnfN57whzM/
r3Bh0NivQ42fvTn5sHHm3fRLjGEdOVGRmlifiU8VuLa/N2Sj2bq1Tr64TANM7FGu
DBTfxLKfcV1qlEBLM5w7jVkQultAmi475eP1SQpXckMD60fswJncq8DMvO4JhLht
dyu/db+5RfgH+wIox23qflLaljyX4k65rxztttdz4dCzHW6uiBRD0DpVZn2zgZUe
iozC8pLOSBPp7fsdVpfyYg76ZK1FmTbIYMSoHFqXuyGuUAUxlhZpTQ+msUNk3/pU
qmNL774n759KTS8/SeDsF56VUgiFHSjN7W2xw9lrGr3bxX5KbPeYLy8q1Raep8Ec
pZ1j8aicV5pHa8eb0dmV7dYXhD9z98as2BO+O8B7JIr2fL/3aNpWplu6dbJiSZPY
GYLsdof36RUb6lNAxbNNtGvMmZPgyqKmdeilEmdcyhp/JKXjBFW7x1+qCGGMWyEJ
wG0YE2CJmw+KUhn4D1duynNBJv4ml9dfhBEHptTKZ562PAZ6gP6lm0UN4syZBKfI
/JBfdOQddyEZAcyl9YV076lIVOAGb5LCNPbZC0+6Bj8+GIEyo7VolIZjFsoUuIe6
HUL+IFqjx5QN8fGK06NNBWxN4udc4/c98l3FdKF9gv7kGrHuF9Ho7sub2XdAQT08
yNJfTLL4aG/tjOQxCPWEvWRHx7GNXE5RJxapiQX0KRDb3oVw3/CSpVhmUZ2LHjiR
x4eFYQ0TyYFuOUo0eBOmzQfXGbz+HCZWuiCWNsmQYdqsrJ+3GrswMH+FLNBn8K72
or5zxCpRlXwz6MsEKCcJGSd7pTgaROkSTTdCRDPQuDfN3zKZ59wS/2aa8/MWrZ0z
FcAC2wLCeSaXAL6fjBRrt2eSmTVtxJQrvCRT7keKjjoPMfsNLFJsOaU5cePsCFVZ
F+7CX6VUHyjXyyoQ9o7edn5Drkre9c3zlt+U6mcnq5BxBPnu6gCRd6z8Q3022H+r
/3XlHAzMdh0p54q6aCnzCNag2QBS2YAbSZm4MHykx4gS8uLIUO6ReEuNu+rVBSjr
InJ+MYICn8ukN3rpXTAiAmMCGUwevaAQk7PnkYUfWWS9pfUWKZdaIZdxKH+Kdma+
coGLPnEBGmoiwH2IOrzcxpWbvEIw5gbPblywSGNJesIQpZC0oI+Mg0ai/37RCDE1
ItTptmaEIIzuTsMp2YoolQLkv5NKBdPrHWCIA7NoIBHUXZlDlsKrRBZDOycz9xl0
StdmqLXM5ivjHk1Tz0CMjWqmV1z6QtqI5FJoYzmos9BDZxgAHWDvoP6IfLtAG04D
djz+W8c9ihFH3ElMDOjesKUAJjsMzGCj6sHOZmwFAF9cPKhqCLS7ZAPsc4Xrte42
X8dBtrBvtB6Umn+T6TXEqeEWCV7We55wCmrfnmqoJhZB2h0esY4YYMUhEf3mKOt7
pwlNjY1LMLAg3R8V2N4Px918a7Ej+2iW00Jby6eDQXF6/pFgN+5OYdK1v22iawMZ
K8kV33APWk529vXB8JyqM/V82xJcGsWpGUKIzP3B/3nC/BFqHf/X6zzw0qzFqzPi
75FYXNnI1X4Ctm2/qCPP+Fvr0HLvkJEoVfef4rPrXZfK2Gi5YLcWjuyJZaQzfGQb
A/JG5q63ONex92kvK2iYPS1vy/lZE56GuYhC1hkHHjCYTan2u/FXnFdLQp4+mv2L
HShz8XlkaIpZjWqWWGyTA9Vi4ez5Vl/bomPqlV/iT8TM6rXxyjv0+BI073VAXYFS
ShBxmlSZaYqV5k4Z1GNDjhQeP6sfjdbtUVOGB1q2+dRjcm94Vf7c4R1aFVZcPc/N
HtjYL+cRshEPfGNq7QuTfz/V9/hK5xd/sbIBjq+omW8pfq+6fFPULHDRiMRet/Dk
THH7DAt7wzqvoyvElXVyq8g+mmjxlIDeJGGg1q2Rny1JBt1k0QyUzL40s72aJOAz
2WlneOg92JU1UBAOmqiaLdqNBQht5bzL9SSbz44BZFS3Ic3yL9ci662VwdMUJs3B
swUuzrg+3w/8x+MGIgEQ90II9Ipg0EFcAwIEdejiDFMmPU6w1357iCq+jq2AhJjo
Wc3ayE8DSNjDbqrVDrNJp6HCYFX7ugNLej/WkMRSMBzT8CmKGSlYBcY4DFAVQOXP
P+BC6JBMlU9ZqwwQieQK7RTeB2hsEVA3coS64Nxpb0SynIbuDaPIj2ytkUYCwbiq
M+RZna5uJk/q6fEzkNqhcygemAZLmb0xU2Yx5Y7nzIkcAPoM7sx3mTvOyOoooTw0
n/K59tC9rGigubIxsROiLHGCUcJ2K9Avrzhz9ohjB6e9UUT43PzXfKBnkYPuCn2v
GD9aVxYyYDQntAgtfV9pregawnO2B416GpL10fUw31RNK2qfnYFV31X+GmYySrMg
QShQ+ca40+L5JSI10jU0pq/IOdtg1hR+8PJI/wPmq35lqjDIgVktz7lRcTnb0Kxt
O9/R9k7rFnPNOxFCx/eRgqacG977nhsspFpr23CQlg5Bs5t3Jl3cmKGt6RXdOAHm
M5g9Na8fo3xaX56JeXOYqtgu1EyZk3ywb50SqjW0D7Ru3UdUV7i/BnaRFbeCPbTj
Puf6+qUX6DlpaGAfE8XWW4ScxLa1UxNNGMX5mrMaiouA6FIMnn5Tut6rL9ViCMPA
Tr1g5gGO4S9uCYJMWqRrtfzF9RIj+ZLix3wsW2ktJkYUdex51rMYYs6XFbPdjUyv
c3kKz7lN95KSOZnoC2j3HfM80esdhDnL4ALXti6eAI6xoIu9WlONmSV6wFzYbdlx
XPznbo7Ubds3g+wwxj0yTTaxn7XQLxHgaAgtsBezloO2/az0Xz59dN4CAe1xUlHt
W0t7vHdmXm9BQhPV29DY0KlHs2WOjn+TcKgz18vVMG8gTsQjMF1eZrrwbyR149DP
V750aoDZr3+y3QARgIILltQc3uFOz7QSQS0zx+v6LAiVwO4BTvKRTINUCXJo8RTg
v2PQFyqgVV+SfzEqDcbCjeNgIi0akd+5V1bFOyLqw9NIBAlxutyiRvPiZlAnPx1I
q91t1pgdyLwPZDX6RR21Q014yoKyUjVGfmX1m0OWL32/jy4Nskn9bnDoJdIatTlc
ASSeQHGklNMsrOBdRy5KblCeYR07MUhMc9NabZLNuvO/yUrimIbyhRsHsSPd8gXq
OaMxJ7zZfPffdkDMBVmi10icto1CNvVcK8JaqnRRdw5XN9b0TZ8i9vzVuMk8oCA3
fQm/uA9ainp0W24t1J7OvKYdSQLqwXtSttkMadSR7EZpaCoYh4GsPNm21gEGAQQU
zpnEm3+cXYf5HR4C1UWHpBcvwECsSEXeKNCMfEfLxva071bGD4EmJRBEqYTB8DbJ
skTrlGcs+nU+nk22lXMr3HOSCoDAcojerCOBdRTCKIwYCJ9dGHzpNEx70CffB5VR
HP7c0bk6E6LLAWWw2bxOQGRUv2zW5h/6/Cc7y/sBhJ6cmPZYe4BtEK53sRcrsu5J
7JNYN9ro0kK6zWwmPRs0nnYun35CL30YKqaZgKLpKp5ho2xUh2QmRZ+lA9v6Zqej
H4+8csUR7rodhu+M9NhdDmLrQfuIhlZao0+IO5KGR/4OEgXUW2vLI7b9kXgAzASy
/MvS08Yd+al4snz3XhtyBH8qjoMabxkDwMUiqw4owpRPd+T3noTOBQhe3/546Ndn
fr4zEE7XhHnfdA+SWP078E/aWszSHbct2Mrm4in3A2EhdNexDrQN7pt9P7tKi87P
q4tqPc9yrhiD1Ty1tEyYb32YkYKblEz1kIZPuTZYEl2CM1eTPgpM7NtRNi7Vf/ND
v2DmkuXuS+IqnxF6WKrzLuO46Fo9OYeXovV+cuwR4JeGvMwSBJpq5jpLd768QCnf
StTaAJweeODLuuBQGmjmLAHwf1d97Ct+wskzMGVaoIjFTrcVvamh0t57a8GYV/NK
/sWyUZiDiPbYwnWTyOiPkozmu5wCcGtiPrwhM3jZRSPqhUHu3PUMc2fGClivsViW
Ds0WeZVOpTiQLd0zS9XV2NfOrtQnto0o3SZarkwpRRzmJbOjjMt99h0pItrfXJK3
BDlo4/xEi1Tu0TwlCgikRvqu1SaMoAK6QR4N2mZmUxWeMrTYuSMLWy2ALM9PHjzi
DFFkvDaWyubw5T/NnHeke46oH++e0jQlURudV+tubcEG6Wur8XfMTGOO+TVCNb3X
DSUaVCTUcheJldYLZSluIPLB3BseNJyYnpQryUwThDpYQaGR68NXdDFz0uIdhO7v
qpXJ5dpXhqDZQX3fed6ryCLhHvuaOhWO+mAb1NSuqBFNDKXBJFaXyF+likfF2X/J
pyCrvAg9FXS8fGR3DmFm2HU2dcfbt0VsxpNfk9BxJ7Ej4NsYRzh+KwLkO5GzzLft
sHwEbb/abJKHG++1aGjUy5bAN5403vJv8Sn/73AUCnvmIxtVUhE8S6nNwG0NTy+E
KbtCaIWxbh5Muu4qD5AA6nX+ypL1TMkHZPykSrCqUP/s7DtfEimf0pIOoYwrm5Sv
k9/g07JwcaI1A2reSRHCBh+JcYgUeNRRZE+2iaIorXhSKENqXPvI5+Qa8gd6AukN
xZ3VHJZ0nNj3n03jW1tm+8zVL24O/hjxuaIJ3zvndBgPYkyepWy4q0GWCp8HWTBa
IhBDAJGXmgqjhB3lgvm/tzecMU4M0Kk29QRpwokGlsQeBRg4FD4XYvudLW+q17r8
GRRsMuF2sZiZXvkJi0fsCFM5c0WeKyYVTE/8DfkgRRdmhpNAVdL4/LdfrWriw9Ef
11IKZ8JJcVyW7eC5G198hMM9nPKHAl2G8CDb04Lm/jaYBAfvyT5uxGcw5+tKekyt
SE7kj2g9AU7de8yeH428XL+P+aBg6VBKx+132cBNaTttdCF3c6eepkp0UH7w3coD
3sVuXrAqb+KVeJH+6yZnZXHvaSRR84NtogQedljkmBSIGB1CM4qoWWGDXuGVSMcD
YSSlla3HNPRaAL33rzh1YQZY1eLzdpnYsr7bPGSFqHq01wSBOKCqziZw15q6G8lo
GpX/Ju8lx8nyG3paO/S3sWdVCCdv2J/+P/HWpdH2M1wQD9Ia7wxmhPjzQbpsnyyJ
WbAzzzgYtAuMRNJfi7OWfcDH2VVNMDeR+RtLURzfYDlvT1hUpM9GGbprOta9Wd2p
uHFGm5+MpE5dx3QkCCOw8Z8qFG2PNqdxHqX6cNy+LhwFJLAOiV6TitbEfFY9Iw33
7aM5M4dzaWQ2LE+add9tyB26P3cBoQCC8AGVLWtzcveoDu4OESXxpZOcwgjpF8bB
zX3I1KOKzJid2gR0dFFw6B7gqfh63wkt2ym1tp4+eO+mB2Xz8aCONhrGLeoaDakk
5xdzvktjZtnFzrpjCv1xd76Y+ARUKjQyn5Ox+37HcfmtHLyilx8fQbTlBBlxhNZr
8GO+MS9g7h3Hqc7UjhjDILigENGBWPnMvHZfdUkGtharPhVGfGJY0U1rB6GJIZ4p
p/MOI4mMlkzlhutwd8rl6+argoQDyVzHYt/QHGyMWZ4VMvHZNLdchnU2mw716aPW
Wr10eIYhkooob0x4acDqsiZ7k/USW6VUksXwPwuWCOaPVxAzg/LY3Jy9xcPLtemH
1NRqXEJi8O/EQP/HPdK3ZfTvjzS5WTzlV8So5VTrTOc9SZXvOvqLJNL2HZHRo0Ms
UFHHYg4gaSkH2PkPosGKW24vnYtjILj26iyZB4ePzr6EheIu1HmUuI+9X2G2t2Zf
qdrIaIDybYYNFmmdDpH5m1THKnxiAkG50q6ZmRsjGdxCZwDFqqRU0zGO4TqA5+6N
rJ34za4yk6jsMvidxpyzXoeXfZZaC1n09fwnW0YH5uOXdvZFw7oC1AnXc+gbPzGX
DwMmYkDkL1axAPhE2FzTnLREoaJI39//E4IS1JdfoRl9evPehb0o9S6yASCkeGZM
DdB23yx5o6O0F1mdhq4HsYYQI/Hr45cOJoFCzlcdxYHGvGjXvHrMgo6iPOVlONyW
mfraf/M7+hdcah6uuJbipqlUJ9YVG64fYGg8+p5wauX5yeQzgX+BKF7ZvfvI2sut
gXCX2l/3/b5LXfSZfuWbDr6C1boCcD9zdRLUl23PIVrs4a+eoeAf1a7+GugEDzhV
YLcIgdEz+n7iK+Dpe8N9YrRlCG+TDq9E6B9g5xG06tP8CBJapUEtRr67JqLmijYg
WI1EBhL//brZ9UrSM0U2Tb9H1zhEyNKLp/8BzRczXbQBjevyFiI+Wbgq8qf+kCVZ
mCYW07txoE2vyPvI6fygO/O9apmndqv6xK+g+v+YmXdRBi4QNx69tr09YRlFOszk
4jUfikFyoiQlYxlvAHEmjvBOcs6FtdRdLbDvQeutLnYsOqGIDY1EewvWQckIQtCl
FazqVCoEQU4rfRICfcfoNcDelA4nAVrzGm0sd5LzGivoBoL3Nr7ZSAOq8qhzSjqh
eclIB4EUAUBcJilGy4kObsBPopop3ce/lLRpr9pyOfDN8Z1+dECSjdSIM69cmHhb
ZRz9qAQUyUMYus4nWEgC8Vp7+1HvtWaItHW8jiU4zueo/i9ycVR1jP/nTYOcMDD0
So0lLvLd320BidC7R9YOoQqUNv/a5aLSDNbZOWRPAQbIB0uiF2hb+LkvbAR8GSHb
Jb9ms/y0V7FaHCSbgqkE88t2FXaGRSEB/vASoimyXtALkViM05Q9oZ+zO6ClnOPv
K439u4n3ikJs49s0cSFRIjTy26+SugoswDGzIB5iaovlFJwnJaZVgQInLM/OzAPt
5OiJXKyW75L9Kk4OoRYVijkJAQmWkCmVRbc+/JYnVwSsAHadVCJJtt4lT5BPcKJd
d/Ft1EHt/gZMqX87Ox+hMZ8+5rhoapulOmz3EkFEFygoo5somZY2PO87GeI39Sgk
qwt4Vpu9AAqjWW02ap2EbXb84iqLaE78b+jtfXAyl6Jl8U7b/1BS0ElWFcHDmcdc
+bH6afexh6cO2bdnzkNW9cCzw9A0VIhIl0uKyEBmWBuMBJ8YQ76fV2lpWptqHyRs
RiL9AhAMpnDuNHAFAwLTQD85/nbXz6DHfizy2TjzBtdgxC1R1PiSQh/w3rIpbUG4
ybnsSkePnPhSJq/lGlRCeQRBNd9tHxqEQHuYUt4IyBCQxJPOY0hiDvkVXTJLs9vW
LyeVrDZ4/1ZaYcJENa9gRvynIorw9wretqWSKepxHXTIIPJjLGUsAISpsPQs0kv+
SDrEpo4e1X+HiTjJHxykAryq4zQshxR6/hBhmlWqZQDkEass1r01D49KYh1nUMKx
qyqkkcxeEE0sPvFK16Wz/oKOuxAmSSXIgOprwOSvAHqMVo+8KK5BcJO9HjLoXnCT
MlDC7zNHjYsKkAbl3fTEWlZoy0jz5B33jGWn3DmAjb21GvYWAbTvuWwk7v53shLA
M/QpQmwXqVeS243inqXkmiF2y81l0Zqbu4YBUAwSjLni7IJaHAJcj99+t5Dk41OM
das/mpPBG4+SsLp9padK0TGHfMMQPr+FsyKOIki6P1WOA6ag+gL7nAstOz7CjOCk
/+PUdha3PbKYgtDgge149MzGRQmzB8MMS0W+Aca4QvFNSlLepQypnJi43+di9XAB
iUHtvWjOZtKd3AJAjllQeZnOdY150D3SGwXbNPiDXPtQ6ohxBQDENgm5YnmfYNWd
DxF2tgwpIeGEjNAujW3GRhT0Eblkua4CGe/MS9ABg+KB+pPmOA5moRi/RvOIvZ8E
+sDzkpiUYXJM8OUSdtTa7kuxINTl1nenwgkOxKl5hW3pcmTVslXSQqXtLzOH0oxY
Viv9nwkutbmGDBJa20v+Y2hTm9sxCi6oI87m0U5mR97FYaIYYaxhPesIdh81UjlN
nP3R3VW9qctAg78muUd6Gn+t1j38D9OOiEaq4nBCvzm2ChHmIdjRgKI8Lf6sFC9s
CvkFznyrWP3qPdqHncwhUVOGuajlpHej34f1VyVOVq4mFXimhT5AeqU9XWrXnkR0
Aslwlq6mjhEdHWWzj2zHdSG3k5GZBArsNYyN8ScjXse66fdDkyoe24vi1Sc2SdxU
owkXCOi8VzGC0d07nFcTrurTCbbKX/HQ8GuqNlYBGEGGJuoiKdn2TDVIKGScFR1C
jIUHLXvN7RiRPdhZ/i1/xyS7TO5/ZA3hVW8PHcvnX+Sys1VHsMmSPtLb7ZDQO7X/
b9plHo9DC2EDD3MVggMVBJYPlWAhCTpLlc5NEP0Xcmr8/xLOokrTowBpEUpqXrrL
tyQnvNnMitTJWsN6WGRrWnnNmri+k8RhaJWQeSnOBYGbB3E13IF26ajXxJGME39A
qk+GHlYOc0HADS3T8X+6PutqQA0WM3JH6CI0EgG8k4M+yyhljIyX67Yz1tv/xLhH
wfnd+VQ6JrR/Xe6guwmYLYPhuQNHogWhtpG+ONd4pvVQjw+MTqJ9yxKuAIthSmhx
1dvD9z1OBRV6vgY9sqNMkdDGkY342SdxGtpNpetl45kfrRB3jbiVH0/Kj3OEGcFw
J6jT0neu3ITVw2kKOTgtCQlLDjfebGSXh/Hgt2luYmoYwDJzVg+mjPo8FeGdjfrm
VU24i3rElCtUzDJ3PET7eZqY+q7wFkyt9RYfpfHGk/67RNo4qQA1VZm/SBEx3QAI
cykrjjzAyTscRA3tHjWlb2KkMDtCj+JxZshTZdfkTZPj3H6cmaDmegFWa5khYF1T
kwJOGOhRquTg1ACY88MdCN2glT0e8jes1Fc7TXYUa0goA0wweVh30Bj1YleSlyT/
zpSQX1mOVGWOMmJ8D5l1QA+rLVG3iAZMshLCiGQr6IOdy4ciCU0WDmlVFb6qYGBw
mT/PneWOLn/8Scnqb0Y6RVBuEwK7Yp8F7ky1IndDBlrugvAh5ycoRn+1KV8wevDi
/Ff4eWdg/uwC6SGN5d9D5ewlvriYLY6L/c3UzS7dpHl046Rv9bQqIweFbalzXQEN
a2nKLpOQj97EE6q0mHm18NP5/6zIzXZt+eaNeo8sKEUTSEO4CdW5D/FTtIOr4/3E
ZyITsmgBs8A1iUzSniS6tys2UlUUef2iBXH9sIF50zcNgmtCNBIAg+bi2loGr0Io
WLDpq4nXD3YGP5aJU41YpgcrPLw6CFIhKapMbzA5fkhBhLlABpMheiN5UxGXQ2es
lTPe5bBPpmuhx5pw4nJDe38CTfTFFdT18yrBWKBlj3E3uLELP3T8oyV/EvZ7NHMf
R07kJOom4vE1JR2aAKOEkNjF8ylaiudfOLeZBohP0M54YlQmAzWRRQJOz1Pfd46q
PjbW/olZLXWKPKS1mrIIxFIjOha6ddv5pTuLWFNotVFIsWaCx7aLKO1HxLGQjOIx
3jJBTqgLPkt1bCyb0bhCZqhQ6Mw5LlY1tWZOp0OUynHGXbzdwiT+biA2p6R5r+fT
KkPFqHLgTmbYBoYJCY0Yg7a4qJWYNI56RZrquqd5plowmTWZgmJEI4V2eiieYF4y
+Eg0DgAHPKOrxIhTAJ9gbsWWnV2ptDS1fDfSQFoNgOfrR6a9eEhf5+Lq88a5K2/Y
1pZQiC8LoYdfI1cmUZNwFiYRed2ubVHPLJrU4E3DhadPkgxUBa0eNL7rfI7U5wqv
P1zNgwCpxMMMBmReYgqvo4xRiqGQLtxNz61Bhq6r4DqrVisU8X4fITq+v8w1Nclu
y/IGaygEdBqPxQvBLaJgba0uUhbrBwe1Zv/QO7uSM+rXEqECFyXXeSHosQDHwvPt
6JYsdc8FnRAd5GuUSNOT6ImIqrIlBR/RCfMafC7hs2Ybn9I9TTfFhMyPlQw3ggGD
ilEVYDiGSEHuaRe3ykyguHDB36VM+oQE8tV0AA9tJLSKmlqa92/CRkcyAJOmtvw1
GZDKEshqRY6KKl0WaKmjk3NOGKapugaA5bKFEESzV8UIxIlATJfKpBGDEcXvOcAp
djNrZo2bdOmoxo5AO1sSxDkD6U+8M3A+ilBzMQIdkMXOOBETlPMV3w7QEDYFDUQX
n3iAPsBZl0agAhJ53XIkp+2lq9GS7yy4zY9S1NHzP9khUE55/u+WBr8nx5o9Ykq4
y+GhMhMwE/TH3RfJnwXHP8HdzT7m9BUai8vJvRw6dJXUm6PNBRnrk9LQANCcYaXh
LshDZexFBEgsSPtKD+ChtpOe1zcbh4zgPZjd4rXmIphmo+Os1GPnECavhfhRiQ+u
ToHrzN0q/KQwk934auoJspyH6fPaZwBtemtZSgJz8fj7hIjv8HtAQoguWGQSrtuM
li6SCkS9ql3eziVzPKHTJMKzxJNDRvle+5UXL+04eu7/GM7aG2vEc3ogw7L4hnrz
e5x+f86AwrY6Lx/QtWEprDIJJdHB3xvg/VYBxKqbLpfPV+fCdiU6dOEoN4trGJui
nwnnyJVavvmDvhc0MrnR0vD/+cu1Q3SW07tT8guEgMvY2fh4P0LWqwp8CacJS8n7
YTQT1Gcc6fmxhdNjuSDwbNa8pij9hZ6l0QK9ECdvjJ8KaX2GiY6sDaGfc1nHHMq7
vEJSbhDjQCbPXSUxyJQMahX8aefAAF6CYGj1bLIUWDIU2qp47Pr0vWcqiYCSW5v3
706eWGBPApfHZ7FDVgrkzPqhjfoIUailsIt3YHLLBZS1P0U6OqEjwGSTHj++N5GP
J6bwkcdrsN7ivKvaf7X7msgm8GOuAKbJADOw5RUWoXAEilit1uLgU9hVP4cIaRJG
DW7GsB5yt9Rq5tYNLVUvHweI/u1woPp7ZzkrrTR+cO/Ouqf5G/VMuRfGrDbyrh0S
PDn1Zvl6mxTMsqusUlITZWLUF3sdG0vWWihe0yk10pb3roBB20XpL31st0Dzp2Hh
pRwBEQJOHmQ7iLSaIqOjF7SPSPA2eer8d3sERQJ4YxaQyVgG7YoA1u6ls3iYXxUf
SdtAJV2mB1PM9DJF8PrZIhx7K2sFBwcRZZ+5ReJGuglFoKRhzwoPNLmWd+zQV65v
PLn/8aa/dMQgegx7YUpegVy3LT/HZbNlfb7L4OepOBdQwZpL1yrS58EfVMZeJRT1
mUOE2HSph7LxXXw98QmJ+rm/g1j7zZVsXd0cB6mMqzKcz00q+0/Dnq/Bjat4TfZH
DKSAih83I7SqH/tMMG1pTGXDCHijlVxPsVSdRrh0UVbSLatSvuA/2qrGWEhSpTIX
tCLStbb27pMya5t2hF+r10PBivz9mFLIH4XMhEkQmX7ydwfDx9H0+t9gwUAnADKb
OB1nu7pEP59zo+D41pkGuKBNrOojAq8LfP2dRBvbD2uPn/KlR1bvxkSCDLZzXosE
neN6HGWUr76azKoHXCBPaItXaYJh3wnej10YNjHk8OIFKlMOffCiPu7bsMMWTIWN
5TaPRxhmQEvKL65yke8LnZYY3XiKilMRw27PWecNnY15wP5zYmtWzhZTeX5RIFRd
dvMNzGoKJSYgcaxeR4Bt7RozXFnErd+8YwTaU1IOqQ1VYtqAlyds7S4+3ba5Mpac
BYWj78xDQR4v5OwgSTMAoL6+NnFCWwPpUPfymtUHRQfqYkRChf6/EGt4RJ8ZIpm1
sLLNWDjmkeVyoU3jYRryrwHBV6Vs9tGTD2ybxrEJQrUp6JEUE7lMDLzwk2JL5fl6
Ne18QMyd8FXp7lFFws9rcHhOMkvq00H13xsqoh3yRYQ9f3pc1ZhSuJVLT3nM5GZf
ivYvPzQ2aRk/+68zkCKaf+C3iXdYVr2QPTBUlarT2W+THjbq9Yby+xwbCDgBWgNp
TcegnsWFx3y1u+14Y02p0PtFKaUONW0LPoxm4R3m9tNK1K7z0hiO8/2K5QJI14JZ
BoPKz3MrzrraVdYdyz61GWa0YxQ5il6ImWU9cC/iLbRn3fKiSRlkth2Cu8XeqVXV
HDP1W590phpxHoyc4BOQwi7EZquXtc/r6zqZq+rM7KTUb2vIn4moIx08aXGuAOvv
GDe9pBrv7XBCsGI8odub7ApwZTYEQpjHHPlJMcSEQiiZchG9joyPaZ1o4g3iow8U
/NK0SoMf0kvDy8GhmAVddcA99WlEc+n2AyiG9t7C/4GKOcHqTyz0GqJ54mhhvS2y
PFU3xFaiyg/zHg5MK+sI+KMecs9YMvt3KSYnx4Nw2xBKGT21MODJjTy1//Ktu9JS
lfYh/XYcT8lghKdPjjM4yuhDDBMAiNz0c7mMHjuQbBUilOxlAozejxe5quNBM/UE
mfvnQc+p2r6wo5CZQq0A/oY/tBy0r0phW/UeTEg+Z1yf9kU8lv9pg6bApdWE2WcK
xcvFffoQ+E4KsHmmlZbPnf7i0G6XE6eiWUsDzoDcUm10DxcODQ3iJ1rV/HCQ8lGC
X/1cw45Co2p7rJ7m+z8Th5jaHrRf54WK3ORRkTBmngCj0jesz5F/htl+POYu3+M0
/Tw9v1alAGrB7zhQKjtHqhbVzIIgjMBRzJgUFdZ1WlYKijGSf8Ib6VsNuq5nSGlV
2rRiJDHVly9gcsVHKzYjmztudqJZzErzXiL00ARnVnED6GT3iSxszHZ5ZX6OXkxB
O2mYDYTdmP1+zGlQkfDzW1r7gm6sW81P7piNUG+x5bc94FGlPS7WhfTMyNkQZP8i
wvpRoGxfWtnXlej1b1wdd8vIAO7p3UeM5rzS+LhxjdFygpv0n4coon93bsLufJG1
iM4VCkC85O0CxAFlOHFU5j/sczZigVsCLRcNU+wRo/g/s49AK/GP9qXOB7rRW8C7
rWEzfZf3FVFzqrJGtZbBMKPSlmJ3sYPH8bWVZSsLkzM0OSMzPgY9kY04jD7Sv1zU
FEpEPzrKzA7QtYWmksK/NMQMHmnW1ttxwZBpc6aPI6IrVY4HzKobrh3iBLKo6B+1
AQOkmN0WioCBAVzlsTbU+w9TtfaCOTIJ+ZEauXzD1ifPL4lbxk2mYvC14kGeXFvu
BeAWPdY9PX/kD2oC6EXxwq7KOhehXdGllaTUKe2Y86J0aqG6UMF66o/mHVJqP6A0
jVaS+XM5ci6eI/fvEtHdclStpqOyJuS1wdum25QpGFW66zq6bV4sMdV7pVowvKzi
MO5XrHhYgFvKpWPlxnJyYynM3ozZ9eEmRPD4IAVe6nVQbT+c3i2oVWaxXtMmgdAM
V9WnMKEwgYuzIEzgrLlk1f1xkO2qh9X1oura2f+jJ4H+ewCoEreIdCincrpb0rIj
p9ubT/A0IQcnBREm5RiChAWdtYwStXDIOxfl45SjxQH/H5FhbAU2EV+1OFBxVGZH
OfMhlimUWHqzARKSwFQt34MxXBAOU7IVaFWtN9HXivdi0V35fMbwgjRe0+kbzGbn
qnpCA1Jg0Df+O1PROebg63NOpoTU5EX6x4LZPUoY62Ezrjhv6I8rkIP0KrYOhKZD
es6oqBx7UjQykjcSpPEOzRXn5G7SFDI+LBFN3Ksi3wfrZJTZnjC7xP/s5ft4tp9/
5X4Z1qGsPnq0a+4txXLsltmFEP2bhggEDmHJ4JqTZLwzK7oHIcLhxVxQG6EqDmjz
fFhYM7YnbPc9Nfl09aKxMZrbUkYoO5or3MzQKZfmpaqbANQzq2Vz597tiNjTeyTB
Cga8zeMBqmxJpIFlxDCgux1rIDRpQReNXxtiJpZa5K55BGtJn5ouPhQVpljaUwqq
O8CFvBQ13WRU61J+GAjoJc2qPtnX4KtoffPTs9A3OKwmwOKXy1KbXlQq/mMLfnJL
5vu0KUCKPTQr+9HHbiWdCMTiaGViTmYDa0aYxHqp66RWhx8/Krd3FY+E1cIqJYP4
xMTcB7re2CRxQPX5F/N0nuLvVOXUYknxQD4AEE9AGr0zUJRRKjXxyfv5cS0EFhnV
xTTWyW7YfyxbbDUTzoyixi/WGZPOKERtrddkeQyA56M5XLiNOFCZLuCftMVlgRB2
NhRUntiNqRwmTC8USmeTGi0f/cZ6t8BKSMOf4z278iKohK7jlPofTFclAqAPTh8X
HOQMHm3zaftKcR5+UywRGAUmK6wxE8hDF9TCMOexK8XD0AvMDTeitqUrweCri30a
1lBfTjuIMCwyDuYO5uABWERQMC9y2YMHjLT5BkLiSh3fVoKHK7tGNHJA8I1BIaTv
l/rPBSvcO6zlcRhzad7DHBenupdeNZTYwfsqm7HnXpgTE7UFVS59DOGl/meLQv4a
Nu4sATHFgxBKTpHfIPjMk8OUV9gQPcgs3dve4uhrjIFLvSSnllYa/vDJKq+gQs7J
T6+nnbwc/3oF7XRqjXa+W5DZnMqWBRfN2pc78neeZZQP2j3o78hn9qYAghOc/LiN
YJ9G7051RjsOlUK+nSFEfzRSRdhKrDW1hbT+LdhEVhs0ikd3JfL46qXJ5UimRilo
6oIuOChGGnbVFDvImcFohmyMnL3jyM8Y4gP3QZGjCsjXRuDbbyB8/f7bkBrpddLJ
S5PPZsctPbBx876UUI7KNyvazIhJ8r/1B0cVGcQr8BCZ04cB7l0JiD+k4mWxmBgg
SAaQ7aEpk3w+89S+OCOV8mMcjswfKfkuufc6MpeTzVZBUi/ADyAFtwm1XPfsyQqF
GjZxf6tesodw2kyewkOrs3FL0sIvyKqF0wBVoANZ8tIXfObIMOWtQfXn+2YXPxnv
LJpibUKLPEK8jUIUoE6+V2BuZMUEGck8LbkH+HKYozIiVQqT3rwmnUEQYqv1TemZ
JPIH11wMLwbvJWDVlBRSS6vS4C1Q89OQ4HTx9INr33pVEYByYBLWrswcXLaryKlz
YrdEa6Reel+ECxId7V8c9dGfaTnbDkJmEnE+Ys3DXt/1+TPqyf+dAwzjOTcp1nux
MI15q20CdTPd06bOx6vd0zKu79y4cAaO6dNNQBXtIMDKcbcMx4e6uDf6x9LVhsjC
ydH3BghUKCMgC2gYlvpn3zxpUDuUyALZ4bfPnCAOzonrmL0WeiHQhFm+/ukN007n
mOO1CHWnXYoTHPEJgV5zTdEGQc+cvt3XYoE3uXX4OWUYJZ7bMHsG2M8Z9B8euTrv
gu/MOAqDGHMg+TVMx+0ZPmF6zZFizFfrFc4Va6QjOr7/a+mH6P3FxNpHhDz+08Z3
lwwiunrnSjWzT2yovsDQhp00ztRKGeg818RAbfFNhPhQwc2xAT3cJYg6k126zmsJ
wyLp7LihGor5uzV5bXwG4uHf26gXnzycLa9T3GETOw220mgh2AiQ87Bvc+dLbIJG
aLbIlqip85cCCIuggvs1ANgena3TPY1Ef3hWksxg/7b8mCViyDoPs/YdU/u/W5CD
iTrEJL9N0YIcTrG7g6ugGHe4DTY2NGeG2ITx3Emyogubtu2HOVR6U/zUQWTptFs0
8x+PnGxTqdRkUuUFxaeicGlJpacqOyTUkJQCXxIYim6O1tuGxsY/M5pxigNWW6QU
+9cnZHcMG59nNiqhOGr8/z0R7p7aX0ZBWo5qW9J/4H5UcfIVbKKwdiUUCdmXKW13
Nz4635XANgUeIPm34/ggbP09ktHO9d8dzHtf4pyYvN9CWVvs5mMSYtB7BwDlLar8
cDK7jhOK/rathTwdDaLClRtfC3KvERSa58iu94BKpvaZYPaqPbst2aVkOtmxr+fS
4QCIh8jaYwXMchrCYL5uU3tucUaB0YazfRoJk5PVQXQmzQF1tw0LV8I5acJdeZkW
ehdPUlzKilKU3YF83sxtLzdWd4O8wYMvdr+eZmDzi90c4n0gl0cUZZWYV6mvj619
1hqZp16lwjF1i/dHxTAkme3y0yKF0B8YH/WMAawoynaYTxVBPiUQcqHS/N6D66m0
L5W8TxvBjznrCvnlqMq0jT4ZMveXH67iood4z8RvfvBZOx/enjdxsA89CXJrgvqi
40yAoHZnZ4LvZXL1XfgOe6ZByBPD2UJSavwAYcfwb8VD0U+k75VSJgNCeUjaJKcM
xEX7+WW1t3TDrWdnZuOtboPGbItLIp4HuR6lak9gTcLl1zKer9EVln7i/Fmgp3rB
umrEyc+bTl5r0JDnNlmAHw4aGa9foMB6BSmMAy03tuK9jbk4OGJJBuojOuV/PpFM
8k4s87YxlWEtP91RcL5Mf281DmV7VcbNzEsdYZsGdrPLXxDjyT6fpfit4CG0dwaM
KhV+enrs/9RmzedhQ+aylI8Gt3e0WwuKvSD54wggtWx8m1W19vq0U/fOp3r7fCC/
tC4c297WUDz2F83lRaG8IfYlJh9ShLVOJ/yQIHt1RzLYR2l5OUDBHygrar7f0Npk
6ra734wasOFIfwUXL+RPAqAd5C8HZrA3dLk/Pjrw+YyStgoWfYRZpZi2BB2+f1d2
mMEPruml8ofXL/xl+mNiQgjADPH3BEIWPKY0UcorvZaudZNgGLPSj2m//2RaExNc
UjuRBnRTWCHnnzKl0S3vjaT5LWG2KBdO649ImSV3oBfZ8M4IevWokfpSEyqjUR8R
zdLqrrtta8bl8olojH2ESMAYM8Lz45/ZVrPGAUZQLkrJc4priDZwY4w/n1gqWISL
g4blI9NShh3XFVwp3KmfOWxTWlx3ZypWeZjpiRClHe6k9IWg22qBOvJQgD0hdsRX
PgyprHWBT3j1D7PASi0BuoHhPJ9kW8hTmzk9x3nJ0BbinSCWqkNlvH9BHc8FU226
DVmSLS6c1NAinDfVrsT1BzDhs6wEOa8BZxMWR1CiFVV1zC7HYHLttap7v1AHROtB
4ZtN97ejxcSXQ96W1bgx3Z5cQyywt9RFvha34U26LfxtFeECqMKkWpZ8Rzntpxmo
x84RI1XbC5HnyCqQPwTwCV6t1/UlOMyZBUlsg4u99aJ4puRL8g/ZnqqVXUvyNNIY
nWYXzdIMMdhpWaGZKbkTZPhCZ/+eEa175nMEtBkf+hclMWHlE7psiRlFAtpQzMSk
G1GKPQbhZQZH7EhgIIp9y35XQJylngO6ZZiqBwhOfc12VCiYPqaKm0hYnqfHU58/
1cAPQq5/p/e8YYnIEvDWgHRExOVvHHn+WJKZgiAJ2jWsuu8uO0SfEpW4gPVqwegG
qEJYHBJdJIb+cz0RXTJekgGB325nMXNyfdDva0t0GB1YxKQfZOIsMTi3QtmRsx7Y
UAv+gclRIiqKQ/s8v7di9Vavf4LFrjoWgVWKo7jLQd0XhVhuVOjpvSSt2pK6DgLb
pz6NYM/tbIWNwC3kJ+e4w4NkuA9/D0Jn5vqunyHyV4dkmfc+I0uafooz0oPMjn7Z
suhioGFOGVKdfOSJpneDhLsL7uMrZyFJYcKJnTYX0mBvTKXWETbCgR8dLquLZw4O
n6FRSetit3zLgSj6r/qMZWqkuoKoahEASgd99/XEdyPR+sq3SaQkajbypeI4WlAq
rbsbA4Ov7I6pxfkZ9K2q3oBUdv9HDHQwLnjskBMABl+ZC0X05VGKL8aPtLMSsfeV
6dvLBjaiDQn7AFf4BhUJ5ozZNMtwflGw0p0aoOcAHoSqjgIavrbpaQgHKtbBdxPE
orVPf9IJPr8f/33XAn9BpGMv0nIHSSyxCqqnoqZbZYYsUM4LCZHD4Qb/wX2y2CFb
ogqZh79JQYIw53lvM2aPGXl2P1lyATu1IFYTR+hMWyqYkL6VDe1k7LLhJlraBvUH
eI8BUl2wE8A+o2orulZPnW2ttw+ns1sLnSlqqIgjDNj7wXqtYi18vJslooo9Wn3a
0/j+wufQpBgeNmWHja/aSDRQw6N3ZJz+UAmv84NiauHn3hnCktWCLm2pFOOVTwNx
6Zm/x7t0+3Lvpl7MnD8kPdUbgmIEEsH/xYomyDY7oHqQQCqvDXd5MAAK+SGfhtPt
v6noh9RAKqjuM+80QHxQ1KKT5iTHGibQA17b0VtzaId+Sg5dNSsycXMehYMwL6bW
uCB1vpSe4pE/cCbhki1Q1jKMZkvcdpVf7h+4Hdh+AgsBYOhqgY+N10QStjh6U/8U
eeH6hvLBx9lXctaSmK1vWcXgWjtbjloVuzcSiTGAdLjXNPCrXaXjNHeLHrCEvju7
oF3PzXo52mlFoQxFHMmUeLHDMgcAEbwjIrHiiPYJzLf760YwvQBd/KmEIj5S6UJ8
+EQmwCaod3P4IQB0kt0DlWwfXfZdADpkordpnxTrfTfEvvlOOWzRmfnuHm6pDi5R
oScM/Jgkdq5BBxHYefIbCIcAbIwmJrt9w/FOs9qJ/U+eXWxXMONd1CMfhVZCpZHD
Pu8RVvclcZB5Jkr9lEHnA9G/1ilBfK/LSw9TGEOtrxIt7smLS1+gL4Y11dgnll+l
1xj6MhVVCRs+f1udSyTTzbRv7U+mSopmWEYfMMUvt4g9dzGtfU8jPIYzq5TZnfn4
Cg+Mc8dUKn+K1clKjL48+pKHGDDIuuMsigTswuh0a220zZHo010rCIs/czM4U63G
e7AZuymqzaDL0xQGPVb675upA0rRDZ/5r3Ik5n2QPZ0IT7yxRM3Y0B9bMH9lEkPe
rP7r9Dy1/p+f5KeTtBWzel1VIYv5b6BBgDThvX/vzMB1o0KEBkPDqKEQFrAcvXC7
akG7AlLprkij6FMx20sLEn4zPndRGQO8PiAyVJzWiLYTzNZMjWGRB8JZ7kf3/PY9
i/88wFWlljJ3RJf3DXsUgdDfa3DAXoDSWW6CnJ3BqkMK+hPg8BPzhNS1UTrra+f3
IsiisuFidcRSYfp3ndG+VEgHHS+YBBRTmbOhA7b2oyE0JXNIKI2ATvXsjduXSvAr
mbMkoasuiyzllROeP0vBFJp+unq3Mz2CJU7ilsS72MpyQFhOwO+GhzSMAEUVP+ed
mNAiaCBiwetF8Hs47gtvkHsBjIXeB6U4pbbwb3bI3mCtZZrNds3I6mEu3hsz6ysv
FwskJpMws8DuMfLVnAjHpMMI07qYhjKUjxVOXlBkax2PFxp4j+Dzwhbm0plxyh0a
ExkxSIzhvtqQN0YvN/bJHiGOM8w/7O7OwXZ3RFP9JpgW6YIf03W9r30qqmVMqwhi
crhHw+Qd0L4UrocXrELWcJISZsD7LGEm9iu5wAQ5LjwZ3dNn6Dxqv/f/Hd3s+l/1
SMgotj3Hq8MFIXd4wmkMdEheeTZNg5mQVZspADMGOnBqJYVv6/RD+q9CVQsgkbms
/1n3ZcAPiaf14RMvopBRmHpUS6KSOrNcY0iA+afRRvHEQyVZgupnq1V7GTj+9sJV
zvYY9IOTs4n6S6iTj9m6/ewuhNUnAR/8BfNTHAKq0ARoI10sawW/df2Ft3lrdOcb
uRlwT5mtee1xEgxIyNOYRh++NrVGH4QekzvDif6Q+mSR7KJmZKyBz1BVEs7aWZ+G
xlFEkvVzNrJDaEtC/WFP1n0b5/YMGt4pZCfmQKO431Qk7woD8iYe6mJXhRyODzZK
X0pYNhYV1rOrrXQvm8Paj2FUFz6kifbWLmS0mxaP2n/l5oXQukHZ6mz+vEjjSHQI
EfM8WBfdhvQXsBoPjq3gZMPZ5BELDzxy2JlUPwxBR482gPD2kU0HMPkP5IKciprY
altfS5TaFNSSSsGqmRSAogHvqf/ZvF7emhr/Uz/jn+KXVasE7FAq6q6xqTZDxAu0
yyoex2tcFxoVOwlxEAE6Yn18paOKabs+QRsi/a/IE8BUpo9DoIxFb4zrWaO+Rj7+
KM7L803MOlfn9ubxFrCEFYeJwniw22KkcoOTpeCNQUpvJDoqi9RwnGAdhkQn+e+Q
8EcYddRIsVy53H31hLC2BFnvzXlXhLUcw3j+QKKX0mbyxZQpEB5QAvmdL+/UIDSU
8GRBtAxREEOqybIDRUetX+hYqe3rTY7d4zmBvncsWaj/4+425ZF0gkmFRlzx19zY
atEO+ql6TWHqGewng3DPnkbgn3N0da6OGNOInVvXxmnTOO+WOMXYhceb1m7qdpjx
6+w2VtwxTLS7DS/7kABitfyKncL88JMDnqH19zeJG6onAPCZ8WUYSOJ3c2eTH8CR
RwzywVXri+mAcloD41e+nU6p2PrgDVCNEVTtt6nZuOYyVjDupmcIm3ipPfN08P65
/0QHfn+NLj5N4Y3taJ4bj1G9Q0+/AaBznrNVjyiaw1EiyRrvNkxm73wagw5C2yLQ
QvrV1LmR9LJ5XDYjRMNce0iDw5BvOhCXt6GWIn80HXWhFgYxtx0FD6mQwdPoy7h4
n8GK6I/3OwIBauxXfwE2c7xCxyXkafeHxJxG2XPlPqWhe+fqIiSuxHqtH5FGoz9j
u+2ypYqsPAgm327KBWAdgs1xjqhbhExHu1NqN0egD4YmIIHNHUSlR7NbBg9QbQWb
svnyxlzVpw2C3qhDmSV1ynmcjg5dTYmNweLFEbvoo7NiIWSYz/HvtdBgBMrU1Evm
PHeWU7ijVc24wpAl1SHQn7k9dG4MEvVc4D10yWDcdj+DHQ8uL17+ElFlm4IBZyw6
w32ZudK8sTUz4XbsbAtkqacsZx4nDOKKox/No1l6zuZBezsSanVsu8UGIO650PRa
gUWp5O9UxvYfq8YfXAJxu2fUDNP9zkqfKEcpQP8Pj1An/ADaJ/7do3/e6BIr2+AI
CiSSBl1DGEzl0h8qm4W0XCWgncvBF2O19T8Ltow3CPzO3tEoKJfz0fGDBfaC/mzG
o3KHTzg3SZfqrXenjHd/pstmadBD70tZEIu7k4ad/sRQv4VQ8zf8JAy5fNPsYnQm
WlK5OGmE98a3nNo015Kyei7ntRlBr1BDtjZHPpAt+dRvE0JRD7S+St1DgAaL1jeV
5reV9o2qAnAQAnrbGudsOLRaYKwzXaxuevWPHLyDouK17eDRAK5O1Pd1KHLdSVyU
MnNdQs4kibyZzFsVOOYg3wp2jFATtokuOBzG8JEWY9pAlOKAPozcxosLoaeDZZGd
EiMh86GZ1IxxoNTgknQIr2vJK9eicJvXaK0KeIbHARLQ2zwcjfZe5ShLMZL08CcA
aQ/kZWFTHF7N/2yT6f8zcG6i/lzY+FGHa91itigapIMvHxXR64/3A/GzRsVc19AD
2nor5aEWzClOy/xbYnYRYALUDODHafDuEtw3o2Q45WCKoz9u+XzyEU9SBossz3Sn
MgRDqMHv9hgtWNQQxZtRz+ZNTL3tjEG0CzlydwPDR1AFOTweaTNuqKhr9nDTgVgU
6wtTS/A4hdxWZqXMKTolZ2sFQaItXS6ft9THUbnTnq7kr3k5Dux1zO30GaZNgPfP
le5Dx4F5nSawqdSQU3U2bALtSaePBlEcWLw6B8ai2VHwBSVGGwsPTzKdJd4vadKk
RCMVmXJb0koF0N42JbUIMThJHLjnhj5puaXDdRbxooFVRWV+jfAEWlRgwLZ6iltT
Ro2a57N51QkKvg/fll4hZjwstXCXaAbJCPGqgRFWWEDIWJGojNLuaDzxcdmFpayE
W2C5wA7zdc4F1Pf2qIUpH3Y/KdzLd6wu8J+LE1Xl7r47oit/0QABLAEjFicLKQQr
KyyOngO1FVg1J7clt6lDjTeBTW19UByqKGBh+aDwovUaDWFW3UlX577MiExq0KGy
wy9zfA2BnGLzFe1mHxBsWI49ndMjz2t8ZPAWcqL4O9jcjnvg0hagkYVSm5ZmeUYw
oRgNGjOTZKLjBKoEBS4fJaiM6KT92b6wDtYNGIsJQ/Uedai4mKMu2ZM3twVyjWkK
qosVyJEkdtMC+NauojmlMdJDheAjbhqEagEvlb/F2QOJj0sMVMWvvDyO3oedZdmI
Yy6jS/xu/EtgteHODZ4m+HMwmkWuVA4n9kas2idRcUExo5jKQ0pc+x/Lf3y7BrPj
u8m6lSntxzQI4fece7lOHVxC+zGTiZ/o0vSfgCyBHVNCMiuK+soipzU4M8B3a/Am
z4jSEYPDRyGGzJYD049uMzyGSTJlSIF4HYmEZK6bIs77bL0wim99CiABmOC96t5g
Idy9anBDjG5bpKUqO+k1j8w+8ZTLhL90BKRPeKsCHGS4u7nOCsjfEtnY+SWBZloy
mmNxOOEQ0sUmGMCp5M3lwLnLi/DNl/Bc6iBmteqr6eLaDdXUjIUO8yb+7JPEDq4/
5a+GPWwKduOYOFvr8VXLBUsf+9qFRtXnhGj10GXwZizGKVntnKFCA275qL6vLTz7
B9O5qDIx6XqXDOrQwSE7XVvXvTVsbSIdw3iPPCib+24hAA0+JybelJmXJvKbXgDX
uvgkX6REkkRQTiSDu3vqhChTtsdZJdaMzmVeh+Z6TYWARIotMavPVQTLQGgyqoW/
xsNivRbquGbYYMzJHhX6YYh9w3pxDYXFaTDFPmSwVK0V311Rf+gB43mLrT3TqZxS
Mlbh4BJigAhr0Lk/eAab7WrUksEnWakOztwpXopuOgNu2sv370wNjdODv0lm6XPU
A/ihCG6PkklOyFEX54f/t7SIaCppdusX4DVKy0BFBEbRKW4jY+PAxFEH2vHJMpLe
q97/qVLR1hnEmxO0k9Ue/SRXal4DPu55y/UQra4RkT55p9rLazk72ZqFYpJNDyxB
MvcF4l4vTNgrVOdPLhWZJOsU+ePCqBv0b3pPFCnoxFW/5ViyvjfvyAp4x78bvX7N
NWWNL52aJosYaPpzYAH8pGQWTR7t8ECjnUgE/WLYnQwOfZVxK/S2sYBx5VObE+yx
HLzD0OMrsHTS0AsQ2/P7F6dk7T3kEXlFy2H6IeQmntO8maM0YoZJEXh/tBJ7sbuv
IqRoOaHWdwUF7ITHcOwMsgtuWhh2MUT/BOMjoGEqEjBpaPhh3tMl3Ot6QS3BXJFy
r36b3qRYXL5t887PBqKcrdCYYmNmMkEqPopD5etVBdRpBW4tHbg60j+r9aM9L65w
8DRWUWTs8rGhg6pO79zxeySwnsIIR2D6w4tbqX2uS0KNiUYftMFN9RTsi6PHqrqT
ZASzD7pIDCEM36T2facps2JO7F51oniJj5tUN73/XMPg9qO9lzVcBvk6rRNmhEg9
d2h2QaVmB8rIsp1LZPIre3+zBmIGEsB0Uu73zOHGaknTjAPmIqM2mjR/ysprQwH+
zP0XRNJKybGSQIeNkHnoZjxZJTzOvP9TKqRJG9jUVw0ApuWfKejPyYxTxoOVqBjI
cNsprBdLBQ7XvVEoiGW07uszm4H3HYnr0m6dyw98StlMTgWak1hhM8Zw2LhOZEkU
d2XaVuL/RE5ruyN2VHjqyUCJCzoSAD34PuFsD3Lc8RJP7WDAS3pOFao0uodWeKAi
9Fi1ASEpBiK8uCcLbwePott7eMxRmMqcalvbYHLSahAymPZDT9xQHkVTdWG2GYm2
J9on2beiUeaPWDJxMFP+XWbrinzXlI5JhyfB+jp5GF7l6vhBNjnCAC+ZvSWDze12
CdL53FJWdRQ8KdMVbIPPXU0iOV9GBo7qbNU4ZkHhpZaPUdj9KAZPEAK4VsO2NX1c
yQvCfzcIIb807Du5rC70b2A6VXHVj9CtjNMtz0GdmmkGBvYKqy4UqmNSc+OvIGQy
7VLd222Wj/1USKFrMZulx3tCZUmy6wHfnBSwd76attXqR0axfU6ocT7wdGviE7nm
j8lX474iU620SXkyXRptL35VxEseCQfefzFFxuhAB9lLgumgLKxAQCdXDlXskzvB
55DvhHNpgHDlQdtjHuniDd0aeuRFq+GAX/rmJ3JKR2Txr95DQFJtrCDkxKNpz517
0hSvwYzbopJYOypKG/BO+si98zbP5F+JyGCJiH8/hTNOE1Su+YamGcdqyOW4cb78
qZ3g9T5gGXJ/X9PNnomYwbw7evWTN3R1ccXeBNUOpQnNervfrPT8NZqqCLAkINCF
MUpiso/avnOVg/y+mZnGIkgTRSvFUlyl+C1U2MFx1XXJbYAuxKaqtdTK7b3I0fTD
bSel81mAy+dWA0ydgCP1gmCwvR4jM2X9ae/KGTkyBSYAZBMy8RAYNZkZvH2ra373
ugSiShdg8tlNPHHu6DdbIX7H5tb0kyFYlwQ6mZ418SfT43/QKJQ25sVGDlLCDGhn
EomTJXcju0FBA3W+8B4Esj4yBE4LbwsIQUBI/Av8/6Lcb0iPhyni22Y1RB/HgAYT
3X38DpYD373AT49pmqWcDq6hb9udZwim8rCsp9GWtymJUoC95b6AubwuIKvP25W4
MIa9idopx7nwxLXDljOn6dufd/kCRGlMIIIkymQzlYK91bBXkpKwM3YYFHyxNDOk
cr14d1CySLP/sZs4ZqbcfQC46I7TDypRDS5zvLAwdF+9dO/8Jmzmyne6sw+mGT50
wByutz2M3eLrJKugR7xzqWeqQhknygKrBoAwgkd9UUmbs2REbpi1w8nImLgl488w
wUFVvA+2IQuH5+WKNdDIPC6aHxou7gD9TFwqPpGVh8WrbyTwaSBIBg0CVOyw1kro
aukv7tajYl8evrzdYuYG7QlKkHpqbLmUAY5Phf4s5NDKiY1EjIZWTQST4kIngTbd
/V1RkAhfDmtNj7Ba6q/Pb/7V2YGBa5sSYdbbkC7F9B+kCLdvAoyrR4rvQ0KFayBk
fDigHi6l7FZipJewfJh76HiLHgTH434KW3KQ+NQiPO9TFYr+WebAlUexFt/9edsa
avrovKezo9O2HP+qwbBvEQVuxr/RSOhgMbPddizVLGqsFL265WRooeE1LRcoz60I
bD+wZu0XqA96Vnmkp7o7IYDwaJZLZPKvWdw9AtiEJwKXtvkTxiDHLekiRj5mD6CI
fcmoy9FZ1Hz5kZ0/r+xlUiZiCS8yW7K31s7UbS8vbiECi31HGao/qxP0hbLtIjjP
VUw9Ztz+AFQkdA5ccqA+yhFPsfSTWuYZdoDpJm3xMF/QWLlgFYECF14fl+9AGP5y
EnfzTU/ShnVlr+gV+w0dOD7tfZINWa5oibG193sbtemJpROyLyoZY9IFlDNmryTX
sA2npCmK6S9oLwcWiWgJgepx2Phnh2Dq+F4mq5/I/d1ww3zRMI0D4R8ggnawcwoX
bDSTAINpIk3cVJmTUyZThIjoPxvwY1Vs+7/DS77swg6ydbUzqVSWXeHDoXaKN1x0
kvgE4Sh03rlQxLLJHrD9Nu0ezoc5MBAXaVD+jN+HSHZR8vsriyJ7VLyzWn5qLn0i
UJeXgOwrZCPc2Tq7o5nbuO5rj5o3xXHiYq+g9z03Ct+hDabA4Dkp5MF5FUmMYY9Q
oqAoX1z/dXptMZ2h4TnliLbn0c/JXJTO1yKPb7BoedPeGcjFdJdFcpQCNYKoBfr9
IfwqnqieEwZgbSGrOIEbX3yYe38Q95yys6pLgL49wNt5Po4/Tadb4VxGX1Gh57LI
MlGqbobxfuAapHJmUyiVHrpfOYVL3wq66F62Nfg607tFr4Bpqc3xUMAmKuqd+MnD
iePBqigxAO/Qb/mKrHjD2rq8lBJ/DMFwopWU7eQ3NPcrOrz9Af0XcO+wFWjCaCT2
9dVTdwBXLtjgB1U7PSO9BNO9PUAWRDY+2PcqHoQ9tT+L47LGOi0JNcDzOZYn53CO
fvjEqNrHXPVZYBPm+Us/tnLGa0VqbuzplCgh/47HDfWQwwJL1+KMFyW5ezG17JMU
vVQ2pfKfAHZ4Rldv1evHGLymhf0DufVM719ya4GKtnDEC8BJmGpwZ8AN+oUukEhc
RD+Z5Fl2li3RS9bOBTMRdq32srBnewImtLaVF/rXIhp/5XPkQ7WG8S9K7InMwjez
y+LlRkSAfbQ1EvEXvIM7wZU3bS1IpMv6mj6420eiieVV8sDSg50R7dqiXWpYbrL8
caCYrNWDFFtnS9ugDU65VnGoF21yV5hs7I+rUyJm/Li3lMBHg8L1S2y4kKJY8AJF
ZUuxRMZ7Gv3urB0lUg8YuJD8Og5DcupUmuxgvlTctTp7zl9WyozUtZcUfZHNMXDD
/lqlICP7iwYIkSfYGFJGGze6GjtFptse1aI4H1B/qSfuANwk7lt4/+nIaD3H08M8
sTIyzh27FBiZoL6jGcgxRnnIZMKHgeUDNhxc/qNQqxf98aoAqXNGYDMLiZhRG32O
0nc12j+0rpySHVDh1FPeG++9dDOwresO/NOPU/ad17Be5D8CLYrp+HUNtipURN0D
+YVhouigEqPGy4cPeTxqtPIBR3psWlZ0D8vOG7di+VjugDOPyp7/48jAlNjKaW+S
XmA1pvuTFWRO7rUGvfvb+Sr8lpGU0x/vLzvsgahiK3INNejn/gxWtyn5n+gPTb9a
k/o10Gg/4im/a7V9iyoCOy7AKqO7JZVAdBhb1zuBHSsQezUMUKOwcYPwWZf3L50S
SEk3Z0TdHdvMbnHboGHLDJ6fZ0bIK+pujh7At9LTv+sPMDuwjcrXe5WIArpKIl3I
xbt4MoMO2mDvPTF9kG/pJSs62d1dM4oFshQ+NFM7UWWTWsdEXzpqr2lNzEqvU3rt
uFfmehDVkmr7B0ZcpDJAAIDK8PBNx3IREVPsN1QAfDIKh1yNgsNQKtYtq57l4SqA
zG5ZKGGQipKtSYN1tkM4nY+hi6631ClgIQ0YhgO1jcwXtl4o5stgWiYjzqbyhz6Z
Oo1O88jV5iMexsvRfbvSkVmBqT7k4cqozf6ZOkxBVEHSkQvbd+8mgHKJeypMef3k
1hpJeNGoITScc/exPUoZ1q7y6V/A7IZ1nT2k4MGEtq3TRVn9qwrW1xs7QRHmDNuA
LDgL+S6aefPADFYbKDiXa+7Vb7CnWYE9FWV7JnjjYmPlj4orhMICpgUwPIVHknl9
/UQapmgSftE9THxolYoUIgHX3vf1y2Vs6bYdnEHsxgmpDrgukUPIbS4YFjxbhuKs
DqFWB+xLuNjMtR77RPS96Qp3SKUUkG1Mgh+j7xws8fAQI5CYzSvuh6Ch+fEAjjkD
0BZIAGKp47KPvODfowES+dTKDKihtzdAq0vIUnFKV4OkMQRlvMDXxrXQiK9D/LJb
uHTRZwWMNyjwAkF9kGit7XCCZltx7y79MI32ecoRhEpznuNq9BMunbo4LFEoCViA
BaX1XlhluhfKFn1tsGck5qzzYcNT3H3GdQyf/DLvh76xIv4hhh0wxatajnRJyFCY
QLzXsBaYq6l9NSBZv4F16ZGc0KqrL6gIyHbWbfWYhfLstijYjSmeSX1Qw6oXbbr+
/Uh2lUnZ7zf9p6pd9ay+ljrhXptPz6gu6sz86t9fxB2KHLe/+i6I1Sza3cOuJrA6
Wp3Y3Spw+XK4+dOnQlImjkiPv7Og10Pz5ECoSCX9Qtd4LdOh3k7gcJZgUDjQNb8a
sbJ/WL2Q63ZcLHwe/YqlRpDelNAexX8yQezy9ciV/Ea6fMVIA3CZseCLQuACHmsQ
5wezIv5AqWLJlkVEgR1WsfmV2n3+izyXbIvro5eKbXwsn2+W765QvaFXeeuE32H1
fLi0BiGOZVLTRApmec3k1hxa1aICW/RPxrJSZML/wk6swGGpJV1RjpQg30Pj/hr9
bMVbmj6hSSBDpvZqstRbc/rXhZgT0H97pbrj9QmDqQta9iyf0jMOEpRNEbc6fThh
8eBGPkcCypfDe5YHFE790s62zt17kjvTaWpSGyKtAn6W5JOvUHL0uAhMBnboV9FJ
B4sRdSfwdXKzYL60++r0lpZDtyCpuU1pALFW2deRlihnwDoEs8PXWa0DSYZyg6pH
oVW09I06IUZ2y2nOSR/Ya0LTMLZ4wC6aTCJLWo7yVzdNVfINWmWhtOXqgBqS1qoV
7r1gp4Y5fT+qDXC/fyX1BTG0gMDXoRIC2Y3yQZv/R+uhqQ52O/DPNz2bb9wspRLL
KI58sqggY8NNQ5xowtdYuG/BtzkqMOflQgOfe8UF5M0O/Aa5EFW+U+Z21G+zxafp
M+y4y1lM6T/Z6hYJ9T75IdnFh508wXReZNZ/TjfU6cPEVeuc8+h5OA1kQU17MUiJ
MBsVDcwb0i1CYpT1gbW3Y+ckNroWKprvFgfuegZkiZ5qhaMnaE431KHFBf3+QQJD
b2GziERfHyPrPegHv/8hrwj4xxooQiXdX7DIVHX1PnwSlzRVboQUeQorRi5Fs6Cr
DYHZ15eAezar0QMONEk9xPQG3Qi0CblWoyMH2V7w6c6eU5kRlYWJsfAzhMWbzCM/
hBk/xZfbgh7S/dr8wYo0A6EQs0WI68YQn+XEU/BoNy0hOGtpnWNIqQbFzqiKgB5d
vHKa/FWbIYYLGSyPPcKoC8qwucq1y+mBulLNDqnhpNIwnSH+DqAhTuNgz7yIMIf/
MsR2f3V6biRFhFGV2pjKuWH0ap7kEfBPkc0WSskTZPuDE875nZhKXXTd86Ye5mac
CAnR8HVgBE6s4hYdEPhDkRYFrwyLpGsgT3ukEOR+OvwvUTwQuiE/cPcijJd9M2nf
6OIbnVLA+bpx9DuUQzvZHV5+B6yfpctyVMaM6UTvW4Hh6VzNW5SXrBjvwmRMZsaX
g//q4BwiYLNafpj34c6rEb+iSFyFe2pTPVyleTzxzELLQPAcPyjS0aKPRYKOeUB0
vO6VCODFZ3dNtKZAE83KzYLDVPdyxWHZQMY9PGdOOCe6AmLhmms8U4km4ZMpt0BP
STul+5hW+4yzufQ6GAdDxov/Treu2LxU5ni5mOqz+g7zhAjq5nB4WPKMeTfPeDFJ
AE56CdotqsiCRnujKQhi2kLF6v52YZi6Ctj+6/HTbGxnst5BhNDmjW4IuNIXfsYd
xKJKg3qYOGf/uNp6ERs2CA5rbvYcD9EDyN+s/nzSiptPvaFfrZOnwzZIYiNeP5o6
Xdp7A3m7c//qAliUkLWXRv0g7sbZjcnAn4+cnC+0W/+/9Mlq5j9S5mrpjqAyOWUV
mMxSoYso3F4XznUt3pHk7T2AXrZKD+Zje0shtVmnKm82KHLBThta/B4AaZ8XAPq0
T/gO95551Ss9jm7Wqi/ZojOBp7RBStoMcUe7VWGwTorPThu1QJDglgHPj1y+hmXu
GP0K07OKQBTruZdTd3b5GH36xV181pr5J6USDqXtb6S71EKpGVzfpUvzeM68iOa/
53oJucxn40lk0kCXmMeH6wUuiLJdo9nNq4OMDlKDXgceFXbRnIJchvO6EGFeCXQM
4jPGIo6IKRQOGpZjD/uv0jR5ix2rIH15H+zq0yXAdUcZuruNQDYKEAindhxW4/Tg
4fpylCD1MGNRnVSfgUI6DBQGaXde0LL/r9CSTgZBr9TkMEhNthH/H68EyvD8oldT
vV8W4tx3ZeKJu0Q2ktfGiaC+wwaoXfb/GWph2Qu85+uiSoxbgF4e1POJMfe48qVT
dVb8+UwScbnS6m1oLFcMd7rwwhGpeqNE7iKd2aiYYexVvRDD9EhBG4NVPs0acQLN
mKls6perc/w0r/3t9TtPpQ3Eh3aLiG8ltYMefiWs6kBZkPE7izuowg7WE3hlAFO+
tT6QashszsK/A5myclTrZdLmf88bUZsDTD1fGeTh8YcWHhGhg8e0Ec0rCbMaG9ks
qfaiLKzrUHjgFbDXzjzUKu/u44nHI7WpDjMJUC4/tqIjaKTKYrgOQiQiK3UMb0iI
78/oyJ+9pwybbtxP1Mz3Yidp1Fd/Er/WUoNIx4RqxdGeCoMBnWLCJwC+dAxqM8Cj
PRbPFSIxTMyp17w4Pn8aOXqS70ANhZWZQa/7A3EHX/gH4TQYxAxzJ0K7G8Aw7R/n
/Ilbj7nwqiz3BMGxyIqaCVYifskGm9sBCMSuTEQJTraw8Wvh7sxezkrqS3VCK6bH
b5H/gp2ieg8x7U2Q0BmYdaxlFPegO+EwVpR/a1lxelGPeF9IgWH+ygrqBVQGq+HZ
Yhew29jy1BpeMiA5M4PgFjJZswsTDa9KGcQNcMhGHy/MSMPSjhkZ2PdeXRQdjNfY
wgOkb+N4otWhSvtAHrtOnN7+gkFZWFwzpjqnFJX+yiob6BH/wrmdBwRJyLi3xGk5
7ijWg+0xLK9wYvuq/CdPCYMXcq+eJNJJBWPsEeatzLR+UaliZlRAOzzSuCxCaKyF
Bewu/8HhL3Gt/2kjHeUCyu7t3+Rofj/Ao0MtFKZQKWmqay0ophGvZ6NrCm+o+xS3
RQYDMwX7m/jEmzvCiKfSnQoOPnAHkpwzNCqOqhUV+p8jB8WtW5MSQ6Dpobep4ml1
MUCQJgCHLylwrU+k1lagwz3SimiduMapyXPRDiiO2x7Oe+UbQuVkj+959HU0tAX6
gUPTjq1Sh/TBgss7bV4uKjOAkVSEGVUmAkVncutRYu+arkcaP44AlSe3lPaMbVMp
MxY6aH5fP3auV56Sc9/R/VTtRu9+85+QP/0UxKebtlJ4OI1G+JjoeBlQFhxb41UK
8O4jqlXoHwyDG6/h6F0+NN3t1m5fTP0ChyPQlVu28V3jQx58LmH1PmYe/FWxWTgJ
4yMJrujg9QKOhSvuqAaeVRl5DJtC/t9Yrg8Se+0bpuDLSfNdf2EMgzA0LPQgI1Sk
Y8ZGVn2UMgKJZ8tqSiF99omtpPGtxAgZclqcp7WFG2kwxRDNwN41kaeFF4nXTFXK
pl/E0mq73VqgxiNGQYEr0Rt3aunYMvc+cIEotzWI0Th2cuHhq6nYaa5jONL9yqpC
y07TGsYhlXO/DsTEZRo/GBL9hCnIPq0+h5J9jXIpL1EDFBtds6pdruc/kmYyEeTp
Id416AJAZMNWczePnXZqiYWJb4M0PDWWQaZHwyjTDIhao7zUweUlbhDGGS/3UE82
qBRhwQF6O3RxbATwz2mZnN9xG05D41BdoClbORf+cMg3JfYM9LMspERAmBQMQt/Q
lPN9kkhv2fFeJ7dgRkue/jrQIs5F5QGt52QOqXv4FIpw7ueNG6chKk6TFPBGguFf
UlLJIWsAy5qCN/bxzG7NBtVLpjjQDoCWmwlvhu0CzoAs/XIp6k0Fmgfzp6ATwL2y
Nb3j31OIDHQKQwene6fS5/A8S5MK8qzTMl8z1oxRG930KxFbI2j/nJrXoltzuwQI
PYUvuuEziTwKxHwzOZ6+DV/0xMf/ThG+9DGn2jMkyAEMrMuyyMDWnOfaKNeLRnpI
TL4nm6RTAAFsXYrZuhFrb4NIa+GqBKuMjJqsPlWZ4I6SoLA/GSV6Ltz3VkQlzscL
sih+jFj3UtTBgRNM8sqfuLCChwv8YLEnsp07DfgwhaUCsH16QkiZlHAQzju+np+t
PvHAcB88Wea9oakd4tDCt2muJVjJ3UvwEYevcHryPeYHvDglcKBa/umDK8TwXySa
VSssD7V4P/McgDIFbLh4AgAcbh0t2V3Bk6nelYBKZcjmCR1ZA+QIgWeq98qPynCO
cWIOeUPvVpY22pnuURJfODitOfIfM8XIi2c+aMU/SCbV6wXYdskftQrzxEA87aZn
QwrqfRYUcQivr5N1AgJ74Xlshj8Hvw+FI4Lk2DtUm0jrUbwp2W2W+aG5PultLlTA
nxM26cMBzPW2kQtL1pQYKZOdStxSxOBF6ZnH788Q6tezN44R5hkhvbiBVn1I9Rsp
fQodYfEwHuFuyt9PCvcHTioqP+IcmuZL/sfieejL28oQhWFIAWdN4is3+eUfHjza
+QJL+RaprCZLUsggX8s35Lcj/rK9ZrRnu9pMdyQwt/lDtZ6FAaynw9/AVXrFoGe0
/dozLpYehGNoi+5YwU5dPQqRADrdCiBPumyGMubNPzGde+MKaeHIeJZep77TqGeG
z0WOKdG51OEYAVbFZc9W7is5t2yHKui4wnDLwd8dzfJIYOwSL5wKu/QtlctnyiUV
UdnV/hHGf56DWGVWWDvNn8U8p/f4s3apQzpeFqoJ7QWgiCzSc8tuxgfs79zy7IUq
RhHrfDcDwYAx+cCYS+Ytu/UJCYLPyqRuFqPOFo3R/Km2xD00jKr23KvUsnsVXucC
ovWj0EfBmhi0k+gqnCeFwjT63LEORInsnLYuH9sy8o0q+K9zbULIVWC6rWWFQPJp
DR3ppLsf18jUuWmXC4cBD3y0poX8oNQpRErMTeCxEPAkeeTy0IlNRNpUunhRl7ag
fIK9NmhTD2rjYpUy6pNdHquLEYXEMDs/XSHOCJTuiWpvmPMtrOmhW5mcJYgURyWH
Cpm0amtXUPS4Hwv9b1JuJAapvMxmvVvcuPN9fY1TsnOMMSyELddgy6qi/V2pr6Vk
N6iXi+JoaQRIfivY8S5mc3Lc6Ch40cac1xiQ1l3pHzISkefANGF7sMhvCLmWWiuz
bQMHhvunlSaivceD4S0Ls36myUS67R+PQk3K1AKH51HWPV6DzCd/WIwKKKeXW+AT
z3a5oqAQVkbUOnu3T6yJ+AeH9IZRfSkACUXmXF5K2HlIRZGsU6dAF1R5herg87ck
NXsaa+M4OTzPM5b4H3Xif1CJ34EyPOSVoGYkygK/412nsgYdDPmGd1cgJm6sY7WQ
6Z7hwC4hm0GjapmW+m6SSOnmnaTeWY0OVCZwJC8LgVRBcckSxEJCGlKkdN93UZPn
T2qUu5ZZ7Q5FBJOa+n7qCelm3oSnI4Ai/N0q+OA0Aed6An7Hr5FXv5Ev4lu72D/N
bl8HbIvYQ/MHnYqhuR6Rg0EH18ZDyL68fTF0XB/po0h2iqlEdQgc4qq++Tpn6xqu
HtIlZNKsMgBv9XdttHAnyWViP8nsqZU1AXiykc60F7hTskJE59cT/Kl7m+ry1uay
paGv65xEZUXwFhgYshbt0dqveoiGXG/gySyfIx76Vf5Xt4x7OzdsEKpCXjp+agbP
C0XvQG9KJ7tFLwWkDbU37DcnnktBkUe3fqDRTIrFy/HH8gKdeb2fYIMrY24JYFvZ
EHEPPmX6Y6YvRMYNC++AYHQSxmHgkvqTXRLJXkdAwCdDmaEy+wI9fMipA6xk61f9
pwb/mSWr7whQaAPRLbA+FUlPjKVCQuTJWkF2tRjrwfQw07TBxCCFcWR6p+PiWB+8
btUFBLbPP9nkpcTJwE1MgACUH617OOiMxswoKBPn3toCVF8Y2D0ZOLXcP53zTxV8
R3sQ9dJsOrnqyoLo5FSP9FjcMo7dG03w9kaJ/BKb/9v3GN95rinNjaQ0Biepw0dm
RZ16lUvBlM4PcjWM0oUY7w4mZ2VB1xrdwyPqkuxx2uDtjgT1PF4kdIbjM14f5xay
gs3hxew+ykFVZes7eO1KsjbgK28LaVdev5uyjaEuomwFtm+Ph2PmwN2JJHY+jiJz
jphKl3n9X4XICmXHbOJK6k2wtI+BuZM35iU/8OITRy6QWH7kIjnGmeZ5TMmZ73Za
9bNFlsfJ+82OGzFx+CFOotPb/J2gtaTsWtxJQYc0XDHvPyhHq2YEj/2Ic3X1RuMq
7ZutVUWDt4V9RtKmgktxmK+Oj516MNw3MuFMPoW2EP/e1js9zAAc580XnenLGiFh
jH7xSv8qXMQhlqjvmxOj6TfFaKTPizuCS87V+t924304zSxx5ggxWdR3nlztcaVb
FFCDZ0hFiIcNE8WNGKLFFrxVWl7rKUIfBoS5ktTNZnR59gp4xfDwHcpMZvfLpY78
gnAHjnMuPqa0tZzdK2qwbY/6Tr654ockrNQQN7EG8mXKV4Bn4yZbj1ezHqyiAdpU
dd0UJcIK3RBKn9CZzoB96s/6AqF0Y3AXfo2JnPbFWiwuzJDDHME334t33hpyJqLz
nYMarK8kGdSMZ45KJZFwIaQxKtr3s8ol3VaxM0HHPH9+zDfW8LhcbgAOxOY+7WCr
eSbMlL4d9VHQ937cxV2WzjNJlCv+kzKogoODVb8A5UKuez56mJCgTf5TekwADt5L
WbOp+jAhxjjepKK25VA9aoBtjX3h6hITOM75tYRyTN71k2xh6eMB/uAoDnzISDw5
ivL5QNXnkpTFs54D0OWZX9dNizEKTv5/UpAsKQH6GMAV+QPpEEc91UmJHr7/c9Mq
yHlnoDvqEFTnsC6FE6wjFxNftCiqIxyYjdD8veP/HVUT+NAYPsiDoSZoS779F9c6
QJNwDQe+zOcOITNSC4399BxtwGfBGSivq/N1obhBGPQFS6QSJ6SXJRDDJPYrKIsu
CI9Eh7aySRj7t7g27mJN13kyEe6qn7ypVXHKfkRb3py4lHfQfmOqH5oJJot9qd2L
KQ0rsqNABP9kvgl2ib2yF3Vz3axI+b4TiMlxjwA1yBWtEO8a2cl0X6ZnTLRQtxwq
EDrsJyf9E0KZ7NGWF3mV1i4AZwePQBd5F6w6Y8Iu5N3JlXMwuz5bzUbFFNMvz1+w
vugicuPNvY51bwK4aF3S/y5XCBv62l4BGXEkQpRYz2OZiiZQr20OSILny0AjJS6q
bAfdd9sobQHPPY8RfW0CQ5bSA2MNBGAMIptyVI5mYwX/gfkgUbRDG1R9YEBR+dK5
26qG5m7eK7teY8rQRMvH8UK+IzAtZvYPbgBLR9erldTy2SmySNnmfwK1Vpzc8MTr
qFhOMbvCHmgBRL17nfvLBtVQdLWome6NqfOzcEtcMTxRZkfnmCydYanRVBgkOdGT
84J5qiSQ2u0vZYoeVGXnuRdydVXiMT0YYU0ufgflm9dscgU+KbVuHwquUNPDkGxO
g5SKqmSGisZRJJQDwYEczNi3WSPcoQq4H9tgP2/WXnObmVMyVUAb2oelCLRzH4DW
grdYHBfENtv76HZ3I9QIiDjCTlgjQciQFfAEn7lw0T44VdMBNdOy0yxGBrhg16xl
STMCD7jUcaQxoM21rFhRs8igKvgSH9vuHb2zXVq7ZCged/kv6WdOSGaFAVcs0afT
+rfO62UjwMs63K0J2b1vYcGKQOgF2sFL3Znwa3kL8ZuFnv4DWJXpcxMDMKObsgTa
EVSce95Xxv9J6VgQsTIMvXkmDG3AuO3bJlzGwRmVcdSelL7Q5EylBSIw+NLNGvOa
Pn56omD6aQxWodrCBO4XldBXD03Xdh8+G2uN1WTeAtSJzPv3Kfiv2xmz9mkFSQy5
2ofi3wVUQtxcxNcV0lxQBcrp8o6rXo0U6aNvabnPfftinM01KbUP0c4D2udd6U0X
CjN2BJrjm+syFz+fxsGDcAmPsTWkm+gLI1daw8AhPXPd7EH0OAqFRM5gz0A+B7JZ
kNdESQ1UukOIAqzCXk6bUuy/PEV+lhiXEA34Yopyq6qFDoXUj7+mQqHdH7wxHWCJ
mDlyj6/xB2U0N43ER3oVwEuTF6k+mHpSSE/9ojlaokKLP2caduoPrIPtBh2/5esc
a64zlVNNxsGASOLMWT91Q8niFFTOVTNOCj+ZDEFTKtVClK/kNiOjoVFaRP/5AFfz
2jR4iqzPC+cxX+E9LKyBi8vhUmiDxOV44/krVK4sDcUfY8yfDk3kdaCvrQPi4dYk
+FLg7LYZ1CQyOJq/ltIUdXe979gauwbjo6I1U3t7gn3uzRlDuAGjxyf3TM1ZVC8s
vXQ6W6Y6H2NDo3Drw0fLsMzpFcf1Jzlh9WXcev/MGJ3w5VOJlIQGV7b8o1rat54p
4kx0XWLPRZX2NFykhDOXG7zwLpXnJxAyYcLocMACDaVo3z30y4p+CeflNCrSqKk4
evOkyg0JlqFiX7pDAi+UE0toglAq6ChBiyC3F45zYPU0iwd3EnweDH+QpU5locgO
Pd1kvl/clkr5FV0OzmvLQxcm11B5siAQILAzB5hlUn0vh25Djxo95ANTukAa5ozS
vvoC4vjYZoRhS4qPtwRwLdWrfil7bfAkrE+6XnzI8QV1uhpwgdglKhZT8lQw3JCw
I7EAQ3IuVaMqyg3TZuGkOyS450QNTim8CKk8DQiZqQ+o53P4xyJKFwcFzy/qtCTl
YfCKXxfS47s+McSc2syse2ng/H8ZTOCGeetjDzqoRC89Q8CnCbfs6tw5zLHu/MzB
JaNzLJDHBRfyg9JLxhTodlOfTrOTLq5gxia+vjPle/NywEBobItxhjgWxcgi2tWT
EcG5JJdjgwT8oQUpq1DvXGQvBYSSlfyjONOrDHEZXMGNpeMrVeOjsxmW9BSsyL+V
Fq3CLIF8mFWQOOfBmXpK4N+cH6gPoxKIqvYDE/ix5Lho3fuEnmovbKm7OJtKRs4q
6GWN/VAI9f5Oo0vDBVukAXhL59qDF49mEq2smtqErsWFve9416HJATaz927Kb17C
47FqKFZbxxhpJkkvzRtOsWraRJp/lEN36DMlaD23f/ugmeTcvwwSyYwJMqR9tpPv
fBmlCSONIHpEGNOQc+MXQpFLXi9+4Tu+5qH/m22ottk90Yu/o5QuMCdMcTdTcdn/
2T3D8BCitDUxjFh86CTXQKSlpz55scN48666iI5cUADsytA0Y/FnaLot9WLiDL7U
51ue//EMM7QX1A30itt35JuYynosybHUCm6oUlZ0xPceHpLJI5CcFyGtkR9gUcTV
2S7o2G+obFOMbUuoaKm9+6EOH34UyFnUJwf3G8g0kYhFn1FCa8qedn1HXgxRxHsT
gv8hb7npEllO/yA9PUPavi7C3KDnhvh1SQsmOrx4ggGPDnKBIkxvBGiKQhNKYr5K
Rt8hU9ATDUJF2EgUWAabTGQYnZwMLRTvx/FYDBOIxy47FDZtAmAlWrLmtQxurQe8
Q8tUz8an5zC5FQyXXUy/bQMmkWjvnLct+1CNZ70eX8lnau/LWcpHsg2SLtSpM0Rp
rhFVkRxsE6IGPCUYY0MtvkjgkkR21N4DR8DwbZAHhya3XBWScxNTp2nkHKKm1bAV
iaDsBEh7GTL+VVJsJvle+tEi9xFSSs3wUC2ezCRMiSApMxG6Lm5IUPCEvoH19cDM
byEYtlAH5Dsjq3+gbUH5hn8NyQErv/Eje4YOr0Gdy6HlDIAJST0lGx2pi3xCqu3K
0iXpMRmVWCcTS5PceG9xm/7DDWYqesF828B/O0TmLIBAYtc1DGAkpUHOYaxe+g5q
Qz4NhpqPbKxBwZ5qPiYD4xQP9gRFWkTwQ6YfnY8X+lWKuVIzDj87LsKn00eMpV+X
v/0SliIk6xtg8zzUH9vXTOOaTi0BE/YCjUXxGD3kLtZY1HIHZ/fK2jdYMwzTxTP4
Nxmxtm/bo2HYXCzt274hkwydAuiM37p48d/K1Lrc1ol73YLXCC/tpGHYT01SiXu0
mYcELGGXLFZOINQu/OzkrySrwVBHmwLfLbQTIMhXdjvPo6erejIqpI1cM/SMf7fE
QQXno3Wj9JLGfOki/Cpu4t/0/f2tSyOKOiCkG5pOMKOB7x8ZSySag10+ttga3sAb
MSLK8U9SIxHJ+/9XozYHhRDQNZWpV6pR4j6mM+/cByXs4BOp0xJC5pBxxPwgxVmF
5KC6BYtBuICF3SP6xJT4Z7Z8SiBZ7K57dM6Edfzl+sLdhhDpKqwUraw7xgJLxq8e
Yv53OCj5MY+4CCES16lBF0UJ6jc/7HN9lyfCr9Tk++DYR38eFExR4UxoH3AqVoem
2J2WDTaTLvLUm3LyQKM2wxZPDT9ziDPUtsGu4Z/ZW2CScMDfZvlRmuLBN6hGcLtf
+k1+Q+4cMcEjl62SvLXhNCz6V9CPCQHU22SaGnuWsdJg5zF6dDnlkU3eqPWWqqav
NXW9un8Pq/NHPDPSx3Jw/WR5+AKhObmPWUfkhZ4ok6S8uAsYzeQ8Z9XqqBdeBzEP
1/MPjafaoGBf9ZCKTBFy7Ngsa1tldgUzumo1hmqIk2cwO99nJkXvrnSbPjI66/Ic
qc2ECuJHmT9WOA+znn5WUmwM2zuvfxLCnyA6a6aLbjjqgF5Nd8gHETviHgyijOo8
HeDb9TSLMzIPR5YLRkZbUXetw8nNmax02+Hrwg8MDz9buDURPkXujpwNPWRrzrkI
0MkgLLSYla6u8tw9gBc8PCO2AnydOajo3JsLxykudQF0fg3xTN88/Sn6s3OhXA9L
p5+9i1TmPj1j+fpa7bSFsO/BSXcY3M9SvQ/o1IBGEfLbvc5RvZ69q8SSf4Hw/54G
0QYi8CI08UHsTt5O0UhdSTuYloZlbYRj84OQSiVnTMFD+XzWxm8wjSbfhBDwe6Kl
fMIuXLqJHnU1FFG9k0ZA47L6WwbhcFMwZnE6DukWXjQJF4JXJxcqXXr0jCn5MBDR
9NyEZv/0W+mxPFMsi8GK6xwUOj0s7jNvBhS6UFAaZ569SOKjq8wp3kyf+Ncl2hCu
UFLz7qpBlyKJr2YGMAtFpgrT9q3ZHKdc+FFhDP/wiKu+1aqFsfXsC93WVROw+m4+
Vme3XoC0NNhxEem6hTJ4q1HpTr7ldfrRGRKlXTIHXbMUgHGW4PmsY0yeyhNGdBxN
uVAPofF0v8EHBWKiDQ6NSyb+vM3fBMnwwGJB0dfXSb3AX3CyFN89IbvHsm/FALtY
UZggrY81FrpYLa6uLb0DaFM2Y69lGSisBYhmCSIaLjS1N6TvSKtQqwImzo7QLcFE
BeKJhrN9/z1a3donwZ8GZznCeCOWlJFtJMlP1P4ABweM9F9HmKhVWiN8pxgDJ8Q/
VjHyLtJriECyaOJyzKZdOD6Vge49Y7xKidYFVdxDXBj7iG+TJ0zYv5xJBhI3+rFL
LWTfAarKYshCr/FI97Yv1HFyhGDb3l3sm2w8kqeuXNHQbuqitlut2wDE8pB29H7h
pgbQMfMoDTy8Uas7RXriht0y2DFlTHNc5R8Yb2k6FWMBHmNWTLW2ikZ79kpRzaC9
fsSiW9zcA75WKDXwIvwAYFQQzg4fyJPaiPyFlrNHr/HP14Jim1P8hhvk2S8zSVe2
euc+SqQDB52KyzxP3R+pGXIcRyA2QmBdriC8OC6wFga3+dtq8Mi7gZM3avl+zNk5
Y6qauEohhUABIyl81oCYlMPyGUnwXfLymw0x/A7nxLyZ5vFGt3cvRW+KIK8tYnS5
QxbxnqR1ftu/+HZVpdWa6s+e676hOyBvv1QvxLYlSH/4IDSkWFzbblfHwWvpKm5z
rsj1fzVOM39y4Q+MtZwFs/9c2XOLN862SHFC2i4CYO8kuj87fCcWZjqqHfWuk8In
vLYNYgDiDucw9MHiYvIkuKAkL3D23dbqHjOx5wmIskUhLdBva7ltLRgbD3yMYeXK
YRFK0uurnN+CEIECgVv4b42Nio0g3TGqPwenImWvorV3wE/4TNhQnY6I48x6uNop
BZxJ1H75aq9yuok3UfZ+t62BxuFt+SdOotacU7iRwXuhuHUyLvn7xZaxrJB9hjc3
1fEbZB/QCwW/Qy96A3Z3uOCpb1PnzFHVRlZYgl2/9WnBqvrsFjSViXhtIRj/8Pyj
m5g2TfWVN+WFI6Ld3eCSh+BIJKbP+smj6qnMhsv+yIavwTGbBsj5So3+4nLkrfCj
A8IivTprCawMavWdDFLS+FMq2kezXl4bv9PH3cfvo16REmWGiXiEQFXiHrSt7s89
gkltVG2EzaWHhGhCeuS5ttd8jKzo2IaylnJHyo/1ernk7mjiExQie3nOM1IhWQxg
XElkeJttxxVPj3RLtC6y2YlAdXCTEDmRBRah2cLQYtRV+r7QPzhRNwUOqTo1IR5C
F9jKGPvOKhrR7y9QEa+NW0w+rW64HeTP8CzXX3lyN8nvZKCktQWtio3wkMQUnaMU
vF6OUE0MeLn1H26xoxgPKPtGyaT12HZs2KWhohJHETrMn2WQB30gf0eDv8IjtxfB
ODr4YYg0pMguTApTXGJ41pqiJ5NTzDJSz2koBKivjQBSrQCJcDAEGLQEZN6biGLq
8ZjdnxA4UtcSsSnP0ynOVPXHd2TpNk9waMNsM5PyHehJmbx+obwr292OWUpsF09/
S2r73CM6FK0skROdxXuekNVqbx1YWuFF2XmyrnB2y2FCvy4KLZUmgRpUmxdyXBbu
lXRhQDnS7Z0AlDm+mdlTSSfwb1dAEgqLyWzy2/DYs9dKfjkePFfY6GSnx/5SZgVl
6Wa+iL+AlWJkEIyWT7mXk15FFNnOihaHzZeCgx6T6GglrTOux6el2KqOSnmvzKI1
Wpw3GjfsD4GWmMt/vdJYdXaXoGIXfd+A0exQ7PBN8I1vU1YSpJwzk7TOBMg+Pfsz
F4H+ua6s7729Z+T1xjmCSiQ7xWWtopM4RPTKBP+BkRyIDFItj/ekcMepYCEgF3O9
j25Bzg4Wf4KhM8zn5snVIC3ymh5WK4qObXRtL8G3t3X8cI7W8RK2ABo3Z6b/WxO7
TCOqoOKBoD7NkTFWSSSVn0Eex+eEWm0Gy1HOmwmVrvTdM5rx3rP+uEleRKFwXpAC
30jgOsezqa5JqSw4Z/imwwxGoNeY952mlHX86MOJUbXdluu71R+IS+PfRqK7xY31
5xAvQfs+DgdL0d2k8qkfG0Gy5hVkbhZT8yuybza87WX9f6cJNmNEgKReEiqtkuwX
4HNBvlVp80j5oNqFtruGsDJmFJJEIC6bx8odJW8e4EZF9Fy6OoHDnYbsjQDRyg27
icWeeA/6D9o78ao7nw/KpcPMVd31xscm+V6ecfOAYMzUlWYXZp6IDX2FXeOFDjvn
SC1rIaTBjIg/XJXJ3xz83QhqSQGrbMfd38QvETMGfA80OW+XDDaoXt0IPq6Su03Q
wC2ZclQ4wq7CqRwoR8c4e9DpY4YYKy5fiUE7+vuw+TIyXyL0qb/Msw7HWCa51uzF
yIVagSC/b94jI0xLRKcbQtZbK9F40OkcEavXkOKVxexfD1KkTS67igfhkeZvBUOY
knx8u9O83pHSZCezHmMEBvgJbqTt1SQlaR5Ofe5ADh5VsfASb+gvojPxXiGKID3N
gwqjpREwk+7vMp7QY6QoMMFlrQD+gg1fNUDicWu6er8M9Byii4XO9A+lfGdjlU3R
M1rGGxp2E0xo/rLOqgQq3+9h7EQLTGVq3GfxjvGU9obp//3qd60bGFr4rkeW8ydt
/VLBT4XYVHDrLdWzN9tWFMkn/QUHdtIe9A5vYzVphl3A3RAwab0cUbIOIDiJyrEP
791n8ZxaCAQtjSTQ6c4EHZJz9BbMPpExVmiSKBzghj3XdVYtunjKwSpspHkmwVg2
8/wXf2fokGBNTKNPyKlKi4+UfSClA5FcqeYNSCsAe/eAEcU7SoJWUjOelV7jaIk8
cxMFEELzOIbl8xZs+eIF+fyYIysMnT6cZldHlxifg2qnMnsx0eJOj/fsQantwObX
OGnGcWSll+1g6YnfHJ9g1ohHJcpv8LZ+hFio62DVIoXiFZQiEcAQQNAZ7fyLB2Yb
s/02fVHlVRcPbBmOWAStUe+aKY4dhysBPjyg1VvSw2Rz5bbeNji/kgWvo1KG9/jY
08qqhK/nEZZ0r6v0GRPDWrvDkCYzXel8j5Q6QGXHqSQeGCqtSwws2zt+WVtPsuOn
WOJjzjXMYxkxD2Y+0AYX3wbsbfv2tOYvPjQ3InvAOFBKmGMu1ZhUEYtyC8qKWslQ
2qSRVQxTZtZ2uP7mG7ukxLW7SzhrKPRCi1O0bJwtG40B5ud2/OL9mCd4mYyDB+Fv
J1WgMQ5mq6N5LVPIR7UOB9qpoHmDwvKBdoGdC0iA3a7OwWuiyuBXbcAh5wvtWuEX
Wp0dc/zpDfIKTTDdvOs28ba0jekXMZ9gZuukUZCR0T8a7N5kCuePCPs2XOueieak
uI/4cK9eME/0wALOC3YCcvj1h4bn8ZuGrT95qDDgdKptFAQmaJ5p6VUMsBdCvLex
FafDVsCLoNpGzvu5FV8/SCCarHX1+qsRoZT5msUE2MrO930jMynSNbtO+FXrAMqd
xz1or1SfsW36xezQP9fa2jCLc4m3PkVCo3v4QuQ7OR8TmVtEIkNaGwbEDrRFF0AO
EAah/dz8DhwVOCPCzzdTSL1OILrlGuDgeOdliw6Ucz84/0TAMH++A6ek8DgixqQf
eihx4nRXT0ayccQx02+OzjGGeiABaZGPrzLJN9YN6iG3dNUW7uraZvv9ukz7rTC1
ImGbokJ0qP08QqtgdB4cSztUpdAysIPYjySsr8UbEvxs4IYk1JETpvVISf1e6/xx
0IMuxJjeZHNIVjqSPKXMMAyiwabvmQ1gEOqRqXXptFrNioOJBXbNMMVlM/msaxWL
7iy3c9VdCeY8lDtqjBUsp3j0b0GSsNDv65JFJDl5bySu2SqgYg3Cad2iJ+Ynkp4w
GVjVHfZzNaTcdJUvLXD5od6lmP9BWWMnt6oR0vOdQv9JKpWrofh3FEiGNSGfsayW
AhobUrPkuLv/zsYw7ypu+PKvbL36SoR+8olmYpFjjkZD5YwfkEu+AP8mWSCT+m17
KRNT1rEVjULo++KKrfCfpNbdiKdaqbGm+7rIDLMb35mJ22a2WzPYLUwJXgDcUQeN
wZy6HA0cJCDuOoOk9tCF41Viu6zCeB9YTOYq6YZCy7cPKpPt/PZu06x0hRdVzJq0
PQQ6F42dXiLVAZD6b8V71JoOdN1KWKhh3cy3wbxNUWbTisP1aBstGYmqrR47BFgJ
Sw21dWIwPFbwdk5K360tWD7P7Y8TElz21n2IwbLVtqUQ5VlKW/ngLo5UA45pPKWO
3RMg2/cAtpw5UG8nL7nktblc2yny7uwEetUts7S5cRAB/mXKVINkBtiy8QJmEcPz
b2oDXXRdpC7td/FBAaMxiNSXGTH/ROAUZzzdXeJeXi+0+ANEgzt2wREO11By5jMV
7PJS6c1UThFK1FHL/foUKeowkZlVgPnqi+wsr5sv5IklaEQMYWWRn3uGDNz/RPaF
7miN2nwxqLFRIKsbN53AdD9tRURHATKyNlzKhZsCjBolbxpfQTLR4UZG+0Hf5cud
ZXDE5ltwXqcNmuDG7tBLmzsuBtlf2ku3L6fS6DK2KsfNsj6DKZ09RDgBeGjVtmFV
hqiyGs4KFnvaOZJRVERJw8C2KVCs5lvoSuu04GGn64TDnUvcmRzvsgZPQEQOov+w
CUGBXA17OMu7UQ4hHapJ+GPnpZdoDJseU4MiSpQQANOupkVbxi/jcesHikJBVb6O
h7UjyL7YNcucRwlFi6xCN/luNmHozbs9zDNW8+Wb2JfyUHdZxj8T6Y1Ra7fmCYO/
NsZVJaFUFFdc1BVxwGQilsWg1SkpTigpanNQWYbgLaDHxIBLGTrbYDpt2/1s8N+X
a9oFOUg0R8WJoI4R9Wlir5cUf44mahcYkLEsAplGYQT14ECI0Xst0zjfej8sY7sn
wzsL8LEB0HhZqrTuxCGqekPNBFhuXVGdRCTFd8nFQOycCh2s54RX8u1eS7fq4tf9
IFTwV7QvYN1YRAs9mHm0PxyeY7yU30zIENXu1uY4dh97lyRpXbdXt28P6JpYsYgo
CYB9SKXNRvdZ3OwUlZjrN+KKlVf7ymMWBm6WO5FKL4dwAEGGPho0lx2mC0jdHrTp
hDXQI6ligFsfLN2a32FXa5yjiZ3NgtBiQ8TOfr1/g+w0tTO0lQYqsnEz1EpSyapc
9y1Wr0iLWzCJvDwiYfVmKsnGTTmj4rYbBg9YCsRu7LbpFC+WvFoM8MmR6h/Ee4y1
gglefp7titfXNAgPWssH8z8A3BVrkGWXyuYrFnnCPRLQSUun4pTriY3LTxesiHru
WfbJslxQ64A6BmuB45O63VSuJJO+NXHyIfsBzDoQerxtbjQmxwMFM6wuWoj6/vbW
6gq23LXULHNtawccSCnqFzdSDT+QrZm3+Fas08XuGpVH5aItL5MV8xyzBFLN1kEB
aKOVSP+3iAjm2uP+762kfLx2hhCb4kz6oxr+1muIibcgV742AEyO/K3UOo43u2yl
A6KUGL59vCQ8iLSD2mSEDq9niopLK3ajyp1ah6G0JMchXspC8KrxxwLlLoi7HlBU
CI8i/UIiX2hNHQ3g2QHSvewEj3XFaCSiyFdpyqLb/SU+UQ62Vw03bUcTlmkUP5GU
7+yzfHqlGeClVHaCNAAPpa/zTQDd75KEwZoojnuw60FQK8iCjSa5U8zcXsw6zYm/
jFaqHsszURJ87ObGmEqfalDPK658aR2HFXnZfM9SPndDAYbetxaGseaZNtX66WEF
o1LmoYpyO/8OC2iRDdk1MS2aQtBnu48logl6whVLBR8oKd8SpAXNX6+6ixN2z9ZJ
j/dnnOjqlL0X2xWpfXywoOG5BzKRuhLS0FcrMfEtolKHDivXa8Z9ZbPFqvDvbKiN
7EF4aygHo6sHWjwvCJnCGacorOzSMlf7ecsZxs44c+93bkU8toejdHcVKO5FYmzH
aItiFRl/8EZuDcJfAYbjQdquErqAYKFQQlHvj9Ugj99ZPkluegNbTtdu0PGX3cP8
ZM5OM1mtwq/Qtt4EF8U4ZgVMmC5PBB3o6K1GdEI1PDXEc9KeHBt88IHcn9h7v00W
PnsELWi/lW/56nJNZRERVFjyxB9H34hVnGOP95ps2GPr//jpIdjOT13z5s7af++1
ABgbnyKXRoriw2ZrHkBpPddsIvTnHqz5sHxxsZTECDNF0wbfIfczdq8Koi4F18YZ
6cCC9sy5y2ygCXp6grB2vwmbEJRAtn9aTzReT8GKNaPBgH1d+hChuHCcbIOUhLu6
Gi61HyQZpNsLsJLk8P0w03VfKuhl2Mea/IBNHaZ2ie/yOMmlm/KLnV22Wuy3KZhw
8qSYwqZ8rLmOqztVyt52Dd7h2BYAYFl2PJ5wmgRgqCxgQSDsZd6W7zLZzH6SY8E0
oqyjd2z/NTC7aOvBJqWNsQNjr8g0TZCJtT2ksNOUznHmb2YRHxsrWR/aYwbTgVQF
CVTrAWEXW519F9BrNoHO9yhvBaFx34mCOYh/f4NbkCrRIi9PtL7aohUIvveY1Y0q
aOo0sLdOB8swoXjbWF/nLJcmUKpBpm2rDZDpOp3xiSUX00FoaVKJQyUrYh6FPlsU
j2o7V3SLJg14TKx0Q5YPVb0CuWLCwpmFDTvWCQeZKKhr6hrg9xXNKze8vv372qmC
vS656Ik2fSWaNBBjK056tfSijmiyLNHsRooIXZ+x/CA+CYRwaIx4SS6uHHztTXzr
PgA2mG7AP48V48Ej9m1uVBPxsfoP2IH5dMYjTG6tI58RfvsRTEd+AVApojA8B9on
ubCeKd/7dlR4ADJO7BTUBhrYAByYSNK5GJEHb9dpn0T2bgN79HWp8YI5FmpGjpSp
vGgS6xxsQs6/BUbwg5vxm4IJRlkr4Yfxtp+xN4Dolqy6CMBklGy3bWdiM+QRnvia
vQzUlpPk5abLZreUu/ae3yHeWe3FQScupExqvloU1P3Y2c0j0hmEaw2vTQNvqALH
hIAO37XN+sm+hTYkc2hFNH1zIX7P3JnFMHDnLvA7A1R2cYiUPjHwdjDBgUebJBkj
oW7nrtyEGB38ADDheuSfmavyPxDvf4fG48MN8WvPR/P0s5SEmPW4f/CpDRtV2Pp0
BjzJSBMj4ZVea+WQJSj1BUpWO19VwDDdmEryssLENOHDMoxlp0AmtztEo/PtGWfD
g/LmHvie4uDTfnozxrCzD4j/zw9P8Rqqp0nPB4s5c3+KtumFGwV1rPeS06wA8gD2
Y7y/orQ/R3sbj9ymtkfLxwIQl1iCkwvgTHIGjxQKFPtr2T+3CRCebQlarYKvLRT4
zI3H75z1b4Ytugb2DDcNQIegup3cBXIt3tgF8utqb4FvqMIGBO+fE5j35UpviwYt
NwMag8ZPm2W9LtuJKhroOmUq//C3RLYqwyK6R9OvmHuQMNgDWr+i+vQfb6Cy6TTh
v/5S6oIMm/2AMYn0ESAwromYsUm+bJQxsmbRhp/+15DU1VmFYpPzn2hKffPdg0sr
HMW92iST+nZC5nUf5uBmD1ZF9xeeaEo6nofl88bZO+G9/EZ20+QYqfqn8bO5myDl
HfmNmUmRKTvxLXAtKXFlSIV9Wg9NceDCZKuQDnaAQG6LaClzofI8ecooHuS9otJh
I+4C0rw99CInXIheD9zeAq+uY3ykVENUzUtsDV8IQG/tiQNGSor+EhkBrbjM5HST
1VLnSNEX8cqKT8YCCG3wGq8j28KNZAlwLoiuX8ge2VRMo+gWGMkWaP9aD8oWD5s4
8kMVopI6TyHMO0nbG4f0XkBLKJ4II6Xnxdo+/RfVmpAgaqMw/pAbZ0u1GAgToMsD
r/WxCKa4ziv4y9qHQszefwPb8zUE55NCCU+fzvv+TIMlO6ptrh5DZY89x6o6GPWB
GvvRO/hL3lKXnrnChiQngrNf0TxHc2dpdtBvLCr9g8ZPsFETvTXK36njeor42T9W
6FJHwGE34rOsNJuXTfyvsfme7asVwR9SdPWXQwDhBxLA7lP+RUAPxZiikuP2PWvh
U6fQq21r5WC0NVzHXhcTsozsG7vbWJSUrSLplXJBtuAQPIJ6o5UNl0L17T1DE5sk
6/Mzu1UtToJdyFZI/pHBkQR5Vf+G1kzeNFOSpmzT+HJGiSOFRrnhgbcIP4uh8ozh
JqwTVRGqETEdhHMdkOHd2qE+3auKiqttmCjfui05/vVETh23C7A9NocAChGZyz1c
HWbmWaHxMkMnMYyzmiHuzHZHeP5L+Zw9dX8a9S/mT0XeCwmfD9MD1wdtLBUpqee+
yLlxyhk85neQSiXJeAm3du91Yq+th9tYVArZiZNkeXq6H5Y/Kb+q4NL+P3HIkWhg
0kNC2zr0eOyN7WmQZmPLzYrSVV44BW0I4La2mkeAYwkEUiLG4H+75VsvZ7uMNKmL
s+Yp9kij9jiBdurqWObZUieQ5GP9HpnNgK5jQ2vd+U1E+OCjP9KGav1mnd8uruNO
3oHWwwDLYQngyD2uv1Ran0+oTpg1YUAGcBXoL9jBKkY8U0lbHTP1gYAulPYNg25v
QYyv9XGC9GhMm94taQJ1xXnZh9tLHHRN1OFwyTeNx4rIQ3Dkumr5h2Bn6meYpNiR
sULfOpX0S3tGcRgMzPCNYy+359oEwn9D7GexLwmxIvexa2RAJHh9tC1h8ztHWI80
IwZK1VoePAkDoofGG68h9i01jrF8Yh6d3Qd/BTa+ELip3x0JlDdA9rNNmo5s/ZWU
ecxUXfU8IFErJ/NOSuxL/i1vrwVWLm0sV0WvkHg+RIF40ivLT7Jqnd8qmOOWcRx+
Jr/woU41S0C2rYCS9cyg9EnIVqhCpD/qhWJvxkh8/e1JsLRRsbYXEWLAeVBLPTRy
+HOIuMTcm11htpqOenVpXJBUAHHT5yi8gVKwA9mr2X+dVUCnk/ryA5VrEBS2gVoB
8TeSjk3v+qCNHJFZF5PE7qiRUd0TGZd1WtMlWBdYlzZJpqmZ3Nzh22flOvbxfEbD
0ntkEKrzosOFUBhYE4e5g1uc2+3xirAIwt/U7WCcOEvhpWZlftpKoM7lx4ecyZG9
4k3GUH2ecp0n3RwgsMz8NU3H0WwC69Az3oIcfifXsG12ccqgjtZX0170YOVdVODn
+rLUXtu4N0dhtaSBlYN4uiwGuEE1Mx00E8Rn7ivqtfgxWE5wU/PXkrLKiIRUBmk+
DeUaiujWDbH521I+cXgTOCgL2VXRtiDEbacF2MGMQfrRUcEaGBXkeB1LLJyTueV3
8dv3jlOb5icKjmYQdnrcfPHfad/sTEvbEkjdF8QPoQxLWHxoMhSyTJdVk9fWaiAA
EI465iVcijEIJ0xsDrP3o/J/17eOdpVwLUHmEzAT0peSkXDNMYUqc51pXueS1VEv
ldEPpcmfcolUOC5WSQHcAfGs8WrK2OUWIyVM6LpInxhQP0RMcuDy74n+9PVuDYXY
wi8mnv8+gwYqUTy6ziuk35RlzY0EQK9qfKm5aMx6wXDqE6A0QuvfkFELTnkJPcVq
B8vDG2p2HA4usYUCWjjA10DznEf/Tpej75j/Crq2RDTTGDbklMwAQ+FdvVwWWyz/
XgfhFhUolgYsWYIV04DTqIwywEIiUTfpaKY4ut2Tmii0TPPu1/sDlzq7ACwFtUeP
bn7ifhypxt1idlgKaUxXJue+IkKQYVkB5ZqQANlzOZ4EtFYiIbqDkUdIb/A8EpGd
3HESdpKgo/LNAcZ+0+4k5nk0Be2COgNTq+AqFjeinQTDhFvOInOLSsQBowHOHAhC
LWZBt98xz8pDe3oa0vBvQGfT2OHK+FX3eUdqcHV7FaFCnoP6t1ErHXNHIeuFsa5o
17B+hso+CrS90dt6kmdqV5LNvEh7xGgphlgTciqCBJZaBW3wsSDmEdgOzXU4sUGA
NSJbQtSfkEwLUpXIZA6sgL/cVHA02nOvtij9yqojawGhQqjWbd1j0IQbS1Zb9WLF
ToBZ7UbZY8Rf5ZwBC6oJtOS/XhIR2UDe4rVVRvX58P3ecKD02iCBmz1m5sXyM8tM
e9zlnf+pzsMjr7/XMdYjabhOm+6XeJ3YRCVuC6quPPlTVTpp22aXitPBtlOxnRtv
Gm1ha6t/jCFP3G1qqIKKEivuEa15yIPhF8gHLo6XGwIVu42qLXkIu33M8qn5YYxr
+YmRIW2kacJ7SbcnejbmgGGupRIItpbe+LRkYFiX6VI4gcjTpnkRWHO8hoNlHrBl
fG7xjZSd6j+EH0gg114zF5PjiAJRyojRqY9Du/gNTAksy9J4MOKmwXz0t+J042eF
c4SH+L5PnlXFkuayFGVbnra1GitjjDwGxVjBgzYR/o8/z7dSLOxp9VdBQYtCMasS
yGPq0Qsn0S5X2emac0ezh6R0BlD102c2yJGiQnupavYIPbOdsB32U3kkwH5nMntS
WgPk8ROkf1Tj/Fsx7hLHDpnsNqYPwB0NhdfhgaD/vAj7u4sogebGxzwnDH06TjYy
1C7F18an6boumL3pKiO3P8AwX9LXTdoykCyUC0vFuS+6FQJhFRsEcq4JC+wnFbeq
c55AcJC1FMoM4p1cqL/raWCm8t2CTwKovMW0+qW9bFrWyz4J3JK19OMZMgVzyfL5
CiN7EjcKI++KNDm8jEHuBLnl54MPdWkfTg0nr2LYio7kCPyx/oZefs4d+5qAgwpK
nNy9dB7XVBvOk8TnjqxTMjJbmHokxVbQUrfl0CkVDuOAaMp/TAAaivsd9cLhhKf1
CnhNFzIOXKY02mRCZ8fQp2gx/1mxgtO8xwy4i5FSNlOSyQ91W8Yt0ft2F0gFheVH
ij6117cBm0S9FwOEVs2lWIA5ks/JsndNRn75at6IXj4It1YNxvUzUCy2vmtVXCN+
Yeh69sgmfemjEkbtKYapmVIN/xzvcBu90vWisBaFbL/t7YqIxqGUbVRviCO4fpaP
FpVeBPXOnHdDcf8DzP03ek88H+fuHWxVdPluF6uuUnioc9VktQXBLa29MdGW360p
K/z6y/N/n33Pntc/mYje5MRTVug+7O2q+eDKDwORSmMP3j6SB0QWomL5lPfiwjOn
BpvGVZEunXFjS+551t2w5Z8oYZ/0ahs6NJRkU7/tOGO2G1nuFW6ymYf+Skotoo/Q
XUc/NUTj+nJIv6TAcG1R3EiYpZVyGf3hy7lPwvImkhzpIirCR9BvKGjpa5WLMBmm
q/wAbT1qobWdKb3zpX373gste2tZ9fichHfaElSaH0HsWtE1QSTEfYdKda7g3Y5+
+8Rnd6yYkDPnv6cLt8Y0rv2q5kmehG+0uKAPPsCxy2RFsdgmi/laltlQtzJclScN
/7Tcp9nxCEJlOtIx9vb83xXXqax04YRVdcJTGoFyEAULvQxNFvYv6LL2sDNtep74
Q/iQsa2iVv4f/D7QOyGKExbnvUGYVk9Oc/GvaeZaPx0qDp3Fn7PBAvn2xXVr7khS
rVeC5NUrw5vbQtuFP0hWwhZCbqh7gtkf7WZCuh3cyNu9C9hEOqDYJdygogzC92FS
MUNOgggbH5MlH44kD56/YfOF7Yvt2GLIY8Ga9QtyNR2DuxHuL8QpxuWQzqFLokhL
tgpyllCqR+c49OSTYze5nAgX3DfeF2Uwr8ovingIc7PKezjg2WOI/IS+7NT5f09j
tPL5oy0RN6X6Ft1lb42CXYGn90wAzljcAU9o3U+T8rqg3wfHfWHSbXjvyC+JRXLD
/2XTBg3zVuZ01U9zUz2tyjC30ml/yZDt0SzI0t+cKZB3sGlAYTZztxRx5zrC2f9k
yBwfwjuosGIQuyBXw1C7Khb5TWo34vbcsYx04LTxIQFzJ+QfG8UduJmd0M4CXxlN
D5vWpHWQdZta6P+OkoetjRYIxMNwvBZc6swrM6K0jfgFn0YF3KB1+S0OksRcDCgl
4yt7lY7uHPNtdjrMQOvbRLHLEABiSiOdXgAnJvLj/AWDO5kGPZGf0p88RtAWS/GQ
/7VYLudjjXK9Byg7qs9FlXpj2QDJdTSuiEX9e7tsNb9j/95WMYBRRwkD/sbXxXBj
eYMl3Fr48zvLFBjVcNhRtAKvTcFPPQQm9LPwlKHmTcfJInpuvJe64SD4VCYNaWEa
z8fHIG6Da/mvL7w46jIpnDwgnyGLXJCAZp2qkzWcKfQWUYX36bSkX8EB4othCxxc
/0YPnvPujEyzl/Qsq1MRCL2PsHfSG+HUpnN4qtmN89kLB2MgfPtZxLUS3FQUwthJ
0+7nuRYgdDpwifTULiewZLXKIFZ8XXdpMqsGDfoP+AROFQWGLbHpBIMA/T+CdRCI
vvssBPXVVzoRvbx1Mp5Gzt8ystWNo26JACBpe7X6TabvtZhVD8Ej8wBIUVURaXfb
UgXT0BOS2BqTE2IHrdyvtQIWGq72S4QqhZoRAI2nnrRx8g/EURjf3uamgqZU5vgX
Jkch9r+ZWrVoroJJL84pxNn8cNxNQRp99bxaRxb+F2S44EXzeBvImcMoHVXpETty
c9XlbSNzrKbkbO6RNmXedjgeNZAi2n/dqZXhIkkG62SXQUtMp9s62TNBK7YwY+cU
tK4dTTLBdnPx3ttgZV1gzl2usLXSsHKs3GD4vYCVuoUKkXsfSW0pt5byeilrO0TJ
AH4NVMvISq8QUMftoOA9PVF/2BtqbmsuHmfSNmE79LLQIVxAo84EuKkdHj2FcZYP
LWCuLUqsenmFd2BsLewzdLxOI/aTphkQfJRfxZWWxTr2+0ARjIOziBSiVjYYvVXH
c/cYSt+h+FrMxTdaME9ebj5/r3GmM4+slmoHl+cm9Y9MGef2t5UO9V/lcpoBSJ/q
QymWUNwPVB/H5AfDqMdoHU0zNlW7MF8LSEuRV+2F2a6XoZePFZE82WJrrGOScuHm
SXEpFOACGT7ahCCHfARXgBomUS/Tq69B/tAr8sCSeITreEnP+f1dxTuxAGbjU+Kt
VZZbsxDs42iogD6eRijNLWfpQYr19upUHEt7eWRIYuX07F4s3kkxhYxRv09KJrd5
G8IUo8xhQXYMG2rH77S7Yhvht1oT2jkvS3fcqEHGoaafyTc6JPNQx3HZ4wRQ7DAm
aBw7Yfxp642U1saiLchF5iawQDWnXsRqhDeyapL7iZ0UL3rOdV3ncsBBF8+eJlup
na5Xv78xRpGHlf3U+fWnW2ijc77T9xalBWh5raZJrMa6cfj23nHplyWRdVqIPg9+
fWsWroWwdt+aNUXKxgJOjDn4LqCsuEvAwfBDGpSrLBZTPdoV36wrUGTgZpGKLirv
6cSIaeYNic7LbGaOBGP88b6WC5tPEg5Efxer9Xu/ar3lcVqOSlsT4DslKo1qaGAB
cMtlrW9mlAHBoR02X+3HQitDi9GxJPAn+7vhej5XrmvTt/wbuttAC6wQcB2T0lbk
QhwJ8e+6Re7PCM7AIJEUeaH+pIshpALrcHaDBAovBgnZo4B3JTBO2Ox9imfLw91n
ivS4rtFo0XST2aWzLOth+wfI5W+Kte90EaJfxyPTWSy6bTk6r5bm3Z4BHQ5xO+c/
JBwuEOvhbfXrFiiVv3MS14pHqiuPija2JZNKDQ+Nnp1OfY+grv5W1PvxhoLpfqf6
30ricCFqc3JEiW+koezYryH8T93H16kD1T3+M3FqRTVlGDD+rY4UfdCiKl0c9TkZ
6kncjapODRnP4aKWWiVx+kzrTW+ei37CyalsniO5DmSFhqG8QZJPi3ivPuCnrcjp
H/oR+Pkcw2RWkYo/UycIRBed9k3NbyWiQClPz3mYJzu6w+eCRDhFm6p8iYaXl/dw
ff+HPIujibsmyka2DQp1s1BpT3nYN2DYnF2FduQbq/8h8H/xr1ZZhyxh9+uPNXWb
WGWiDH9M5jZBRp/64UsYFIOG9nSE2n2TusISsR2FTvzdkkRfz1W5msACt6CJsZcK
qAq3LZmdKh5qRMIJwh+29DcZWutnpGbAay+bsiSt4dylYQfw6L/n/LRGElOEgN2c
rF/E+R+rMLZ6pyoIvi0LkE+pSXZxAeuQ82oXURzbG1hthkZcdycnT6UWVqyo7tbG
Xhr+sX0rf5ZHAM9ZMTAKO2uYPkmoWfWI7Z8JM74cMf05UVzhn9qr8u2M280L33LK
1qj/KRE+TAktmB6rdwM4cgrB1IgE7T4quzq1NxOMh6dZdIesO09lTYRsnJP1b+6i
Ndh3bqLm7tssg/iB2A1qtcNuLYuYieFvAJjbXBmsJqDQO7Q8WM1UlzNA17ojXwUy
IgywWTRYDF/BbLHhgnt4+U52df/T1igRu04XUP1+SsULKpBboRYWzB32Dwg5MzTR
+GmNKnEVlxvalkYoNfn7eLpArrRR81bZiTQ5jIvBG7N9tYKlvL1mBgc662Wo/ZA2
H0TsOo34hfIpIb7+JAGUnGCt23Zbrl6spj04FMY4nr6aiHUDl8PMPb8FwEqUwbrM
AwMcetCoK7D+Y8V+XeLH1z4PJgEQUkyfalhpgGVXf1pt4mcZYPSuBfY13d7W8FZp
4vtmPRf+woS63HeMobmFPPujSmiagcg4WLoZKW1ES7s/Ldp7p9J3AGO7TVdBuV29
7nulHr/JbcbRSNeny525ZxGM//hllUk7iRpeRxeLNFfcjy9fQipQj2xuV3vEOYqF
GaLE8gG6/KXiGVV5esCD0DQh61Z5JaSllA553dIX4e85rJDfngkyDbPaGm/J30Nm
JBp+ZldVEYP5sXSqpCfAly+FR5W+hztGaMe916KjGTkRA4Rm4sSomNwQqEnllAxv
biFocYe7wrwo1vjCT0vqqc3x/vyP34qx/NLu8VE53iRMlp/tIqZeJ0sDv77wyn3y
f7AWap7eIbxdDMILeiyXt2e8tMc9bJPmsackoK8eODs3fn5hQyttJPU9UJTtbwI/
IWoYAbkJWzsOK+YqJCGOJUSMxK/qA9brO1Mkcl3QHZrANitrsZjXHuVIKBj+Ah2b
yxG85M466oo5Z+OBrzONuM7XVBtabD9tthF4OKMgYLPSaiRZpyUoZnAgkNHzcqMB
f4swOxTRelp/edFWxlziFXW1NONeYHVtDiZWoRbtvu1YYpjESa/O5y7k/tMOQvrU
W6VsGrNqsla1HjQA8/DKD4PrP9xdJJA91QGXUe47eqn0BQs5b+PypGlczEB07uhy
aWMKoWUqjgSVyuU1G4oh7DsgG8in5g/neQ7zK5RFxsKzgicAEBkb3PdfznAaRmf8
BpFs87DhgfQjD389SuAie/IgMPJq56Q6zbQ1dws5ush4Kpz59o26Ttjd7+2i79hn
Xstgp2h33l5s0ilXsu7Wzc8P4wtas4POTHHozdzzkxFwaw5KmkeIMTob4JzImYp3
K7CItTldLSW+PIiDQAoRRhOgvSSxLHqhjEmwNXhR9Rf3vFjy7yeEJHGSYWtCI0pK
iw1ClTLQYtb9n1idyjBaF+YP0GVkkOGXLlk1lvXNuNu+rRzjlVWOUoYEmZDdfmjB
47pnxhAvRyAbSye9/gNUhHK1X1biavJy901vBoXveVDelASTho0vYRVvvSKgkiEX
FK9APAXGIh2ZeLAZNJaUUXzkApEIp8sXKE+NwuWBj4nf/Y9eNbQSkN/0BlaKD/X8
6v5sdD/f4GfxTFzqXDN81jCs9rqVoGAy2SF9kUckYSCTZiB2JcOZa7os8NJyDJYK
6GGF84Md4QU4pp1wBidgYnF02avV3z2ZUExonmoW5JRbqQzYdCLxZ39fylRpDgVv
1HMc1jz+xaavRMpudO6bymQ5XDcIPvpCx3OIW1u5QOTHgbAf66IOJf2NAj8oRaTH
/AP0Pt9h85pm0dX1v6yXG0OfascyttOnyb1HeuJ8zz5GfJw12JMb3q3fzPX1ncoM
vuciEqrg3G0ITzGPn4hw+H6Yc1k/BwTe4Amm3kJV7Xb6AZnW0j4GVDToTGQB19ra
whY4+LTL79KryB7RKA13cSh9syBcXpGWaPtn/8orLJ2njSopYgF5jRuwNSOOdmGv
+A2qS8sTQzGa5US78KK/8lioO4Ee31j0nCp7oE8wgzj52Af+bT58YONtK72lCEmz
wWNypiqtWeTP8T6e0mF5HvoH/HlceG+/s6xlbqQA0oCT+1QkXhgftbIugnA+jFo8
b8YpgAkWPdP+/GzZM21ib2wrWXjiOXb+v3dNccO6GOPFpDVX/ZAzYQIWKP9nsvdg
+h3LF8t0Kp9axrRSVQxIrsTpWbqmBkxj+1xGklxFucNDEwIl4pucbGLMrU+wbt0F
RdymXT4GirL48wBO8VldvE29hVaGgB8xwJBCWYSWdVea5GmUiR/leeSqERB7espR
9Ur69rogeW2uhdJGw1M7ecqn8cDByr2gy33E0bNIXrcxw+7lN5wMU0/bZC5Z08Y7
tzKVSnFSbRvH0dFJWOJtueKFJBSq4Xd4JstSwXIh5JVZnumT73DixHz18lfbTZ3G
6OK//J1zxz8As0QNxtzQMVm/5vNtxD/pv+Enp9+AND1vIx7GwLya/7QD00mRaQPv
zJTAXZe8wp2KML7N9I5qzc8LEUlEDNDzUzKjDUk6UeyRX6JW/TjPztrYh7AnUeCL
e0nVMlYl0Cx6SCS5hh0qPBIchTRgzaPWj3H3VE73GubbDl9EJJU2TGkhhaGW3828
BIJhC0eYNPJuAUVdsEVK3G3SqzTRcRXGdvao9uqgB8x6Bb+GqhluhiEJsUt1oz/G
WrooriJjy7hKTzVQz9PmHSuYTinwwnvFuyWyuIAYIJXCznzKW1aAEqiFGY6yqp5k
6YficUIFjD28iM4IP679ezZk1enj3vj5sWS8jj8GKDRYyDQ4UaZPHNqjy6tpp6Vn
Y8GUFQFQgLkocXraD/ryGyWwm+C1zH0vI+r7AXMxIbD6KlqilGaZj2qgKG4tUKOO
bP3WHg9E34s440sX+M5hUE1Tr72s1liGULJ4PTv6YAlIUU7G7HIxYUuQnQT9V+9P
arJKgKjtcwub6ktBtNouVEgRAdWng7lF4IzzKU/ORJD20/QrT18I9GSHoVhYDaEq
3bhvA96uh36RAYpC68Hu8kVrYCDpjTfSK/kmg4Vnv+Q7bXj1gRZPZSyb5z58Av90
wJaiXB/aL5CF41KeI+kRzkQCs4DcvasRO3Qw/RePxBJvzWdRrA7zT19M3IYLxtIt
mR6sx9nj7uP8PwuLW3Uim9sZUBfXJKQb4r63Vyvt/T7b2YLDLibvfYaXqL3N2tmP
y2zkJLmmu5YdZyGZhRrIIwLmJhQdzUF2kB2lChhn+7XMSM8dO9juzgY2qEDeGhi+
Ev9blFOUWo2dxESFnPcbHFSkl6M+r9Wj8piZJwlgD3V5DqtY62RS1q8BGs4loxsC
zAMunmQNmaqb30lg+G/6eL4V6EsXvCuzZ5fg8EjzP9OOyCtdr8ptK5m5sSuSoHwY
zAHjv3KdYnSdQIm7EiWgK/mhG6X51o+IsqemhiV1uE+GcmIHF6xiT/4N4xEchF6i
Gx71QlOzD3GsR4Dtvc63nMzZluYJEPu9rF/zJjXsQOVT+fnS8BYQEXOBay+E3nSP
cMFBziaVZ1RywVohTXv/s1b2OvO5RHZtdbSwvDmJc5rn+AjQFVkwfz22Y/yg46tG
xoI1X6zzLbGttn+H3dykGMnZ1w7n53/9RdDm1OHe1iBuwTaVVN/Qulqpp0M804CL
Yf7cQLLhnXzRBWR7M8n1vnWNgT+a/LAKnCL0SZ6D5pUaAu65g3zL8tMDJGH35h11
IWXwmHgeyDTNtIaXOcexbxbc8wmBfEVFJLfBLbCWJHrem1ObMSF8G0mfm3FxUCPS
NTFIH8uJkeB3RTMs/C69eI322wNj0XInBPpEJ5el40hQFkrscAMwv6SJNwG7cCh2
ut3yEQXkuCUcBD8kC2xVO/4ykFR/lZ8+QXOz+Y8sOS4sT09SYnvd8u7XV8Rr2YL/
pfnDAMC9Grsx4eFn/6uCXgMHXBRRzeqBLwGukYayqgtScz00QyXBlw/Zvy+Ln8Fe
NKZSxIT4gp4Idr+dgrFTOKoaJkiFwHgeVJfdQ+8E41ycniaWtQ0T4pIRiL5rbI/K
EMwtZTCaDV2BT90GMIOQ9OCeftfe6Dx/dQnhNn+QcG+WSng5o+Dn5ysK6jfrihpH
XBoZnhWdwJK9gC8fZ6PLiM/NGtVVmCTe3HZpq8nG6tqEyz1sgBEn+wyDg07b7Uce
HkbmU9ctFxY2MIVpPyQV6yPFoz8xa8L1FLl6GgobvJjLHEADRYpsjUpmSh/5fROs
zmCdfwIlolJZ0LjT2abVUa7OUs+nmp3SP5jESjTCnYc4ROhPqGHUBPxXsMyN0JCr
nmyaTJlivIWW+r+TPWqpYEs41NL2kl81LLxszO8Ib+KbR52v93TF0A6h9u0yVo6B
1FpttKddIOL9KNgKqPPFb4TOxv5eOzdomCbZrxoCS0vIaehMFBDcMi/8m9b8Z3xZ
6S5IEwykCnvsrtRNlggBS80jKJOmSJjYQ3RsILG7mnHuxK0ej5k96+ls4vw4zWbN
ZwVVdW4/AW48KIAx/82CpjqW8HV/3pMAkv136JJ11eEqJ74jrYkWTLzxbAmI2jub
DEoUUo/44yQxbjfrtOIT97fb1q7GQZkz5/bE1G2jAa0o2It7Y7vUlUT0H69GTFYg
mZKnEAL4BMAF5NuLh9wg74ZNg2YHir5cl4e2bgK6hqhVub9bOwNbx9IQVd4WEKY4
XD4ottbWIX7Ivhen2aCQO/tYKiKUef+g7s8EaHk7V+uTtnvGNWt3EzORh5zZMCiE
2fJgwYU7Su2YX/5t0tCx972/zn/h+YPLKK9zJohfwf8IznQXjYgnjZeglY919gC3
qxWx+fN+RjkGne7JEROVeXABLm2fNadU4bjRZAQqNO73SMXzdvkYwWnxDkJfXNEI
D64Yri4qt+OF3QClgrucz9zZmzXeeZhSjkUPOropIf+hDMJE+ufHmftRGbnDGcdV
gtpFkIxUdJughiUEMVfHnzKfQZMhrFxD9HKr1JFlHtZNZotN+7e3aAn3o+ISiqos
2xiq5Csb22aWeDgJ+BcAX2Yp+FVOEIkGgIC67ueTDfi8Gsm3XlDRusLWwdvd1KeE
wVWf8Hkd89amnRixhBF1f+2DR7D+gqIuC2t/Il7++gydvSOgDIobroZ+v54DocV1
b51L+urckxF2pAPfh7klKsa18SOD4SRiolfatO1aGLAHeMC73YOV+zm9/rmzLlsW
BFT8UzPpdE4cUdmp9ckgpRH3cv3jVKEgjVDvKzRqFtN/I/XaZ7CJQr0zKcDHLf2B
r8gM2SoxEyo+c2jCajRrhVXoHl8lRrg6GpEwlol9EhdSveE9TyBYI3xXdiUBsXvG
3E1dC33AHZQbVLv2k+jYNZw69fjgJCWVo9wQ2JXr3ETu95VVIYjgbIFJtl/X5M3A
vuz72I9mdPY+0CMAZAqQNGrGJrAOnM1PW7lHNg5CGs/1vWEBXkZ47q3rvD6bdlBi
nq1Sj2IJm9FsFF1FsDFKYO+WjfnEyEoPB88bq/Ra0cWIaaXPv/SHu1KUeWPl/rzf
Li7S1/vZXDybPGDsMHMiQE0m4w5lVTzyLTdh4dVJXeskta3gBZ86DS/2wOsBQR3h
T8dPomuE5s2dCKx8SM6nUZ3TxJBGyqcUgtBsqw/HdXURe5/3oBF0p4JB5YwanmDH
IxWTqW4t5KjPCrHcE6GJ6iUcyiL402wEcCWJkq7syGD6PPg1D3dlP+QjpnZmJVSo
B8aWKtmAhW/gVvn+3mxWqnGAbvSxHTW3cLmB94WgB4vkANpNTYjmguZTLMqcD2/9
ENB6y7ca9dSgL/PzIPFYF20TBaCWajNjgqMJuJ5IrwL20vJNmFglQa/CVq1Tq4HW
OhN1IPXVp2og/15zF/2HNo1UiommuwyENMIf7WWlDB6Da/3xipiOWCG+nBnZ7bm5
vPhsF/MFNSqTywg9Wmsu01yYNWfrrW5u1KWFGqW1uCyqgekR6jvluKlmcr6qT3Z6
xX/ovMXZTbC96JGmfnx88HctNwPhPmg7gY8UcS9rC6qIIFkGkvwNuf+4XGAWmwy4
HZUbkZrKun44Miu3nxfDmBql3FsJ0oHv81ephzSzig2yKe8J0qL25wPBFGLLCKdc
r3bKpuqK6aeFxs3z5LSWrsFqW0QGZcOFQAQ4IRFyeznTrV5eRIolJ1nsrtOG6w67
wUV0wXT46sN+ojK3Fa/3NoGXCFA2yYo/W5zaGxbtV84IMe5oBXQZcKkHksPnIgM1
aXZyaXVS4JbRZo4rLWkRoL/i9bvMami5D4UWJAYmXFRxwHed6Wg7ZE5IG68EEv/2
74C6rP9Z/jYmh4W76FKAzQOkjNuloMrd7c4+IHwR4FdIlc65hfftx0cegFlqt2py
Ih4BalA/3mWTlufr3kcer0elDVJnKp6ulZ6xjFeCWFF8i0zsuVJIJiE+c1GzsWyy
T7TCPd6k8fbZoe4Xa+d13EwHTZylESFEoBzGC1XcprSq+P2aeBPHFsdzEdbniG77
Lc5eR2Lub9kYcdbj5eW9voUqHhA+eZjLrWok7DlRjTuHZV/rwX6mda7nkpwO+ZsK
Oc/5xeHyeTyY8hLxE2h5/4f/vjkaGkXz3weysAZatgwEY1rRt9QAo0gphlArn92O
a61fU7S9kaF9ztCIlhjd19DBdPl7jW/LASaNtXET4fyd9A9xRkFo6Lnsf4WWpCsq
8uz58Kmh6YqrTncwaqX5Jrj/fFVCum/InSq3pYM0ZLA1QCxpNSYHns3ChoyWDKd3
SGufhU7PLbZUoFXVF9sos7+KwobIDvl2gegHhfH53COI3AzGGR88dF8Iy4zncVKO
fc1xX56+JJihbQPW2e4va5z9z0Z57lgVIksdhdvomrVMyk/ayxunji2HNIEJJBCA
tAkCLM9YPwjr1DrgWaAXUKl/wcfv9FMWToG6p2gcZnEYh/7hDRD1C+PS8688Z3Hr
2UbRtWs9H5GJ5wn2aIL5YxJuwxzwteZn7FGzNWJjzCX0IXN2FwNxzZ86WzB2as1k
Y2cRKfZ/DHM8F/Rqma5av7teB/Sj66nr8F8hCsWn+uPue0paqbFwI5J28ip2MEN3
kYMkfpCJ3WnHltYVx+2rfPZC6vy+rC71vE03v3SqcI8XNu0K6isCD6ZkvGMK+7hX
G6JslIsp76tMK+U9IF+T961QKfbueBWWZ8N7HEumRsjFHcWeWXHB7PTdNB7gQ/Cg
UI03KQZ1E1SIh6BElTJ7WDDCOHJHN3Bp+3h41oZsBCFIONZQu4Oc/G6UBiEUYM4s
SP5pAq3YWkHXzjvvOFUpe5NXYmFpe8PWtbQMlYQ6tAkwFVmN9eQunGk5elP/Su82
BAMeq6qAAZohqz864RkNREeT42aZeLAOHdVhgG5rw8+9ij/BemUkVgTXZVhobOIm
MlR+YFdfDuX1LvNiIfT/s2EqfbHRZtmONwztT9Dbi7Y6ezkgGFS8nOHmGFHNb3o2
MJEdTN9m8I2yBWvPwxCJ27Nm6IxijtV+YBEu6cAnDDcC3VFCSQqhhyd9enOiWHKx
ZoHXjJLg2fimht0EWVH6PNH9ejQ/V+5nRLlegSbHCSt9Znvnd3d5UhrpLfk19Ohx
+fe0e/RA24fCKzyZAsDMJRCM8UMx46tQSEhtyUiMDxeTPb5Qe0Jr1cz5ZG8i+IwH
cycRFPxig4hDDjHAFBH/lKhX9Jqx1kaHRSB5vUHikFmyAIrWd87sqyiinFDp6788
sywdfvMjjCcKkRHD+y0/iCxEufLwNdVfMW4LqlY/K6+CJWBnkwZU9yGIfSzOUlQz
s1cXW+qN2GuF888zHCsGLU762x1RpfnzIxQGXpbVZoB2jN9mNMOU37ghqTgjfoam
u6bHLx+JZ5201VwsYMIeVHuECSU0ehXmwxImyg7DAYTo3yjDxBjHm+ZvSQ8l8GYV
m5Z/MTC6MZ9EtH268NvPLadZPXiMjbeq+vrYVPri+Lfe82gOthZwe2ymMy1IF0Sz
KThBuXUyTjNWj40ysXov3KehG1law1RcbrBikVl7mbfpwL/vOpJF61OZJDoJ7csS
GFcHAvkQV3+hJyOvb69XInd1pW+Ah+fcJqjM+UZH5RXwgPIFa3OAweUIl5oI0beP
7cL4cADeaPs9ppwDJQ2QhBN4IFWK3qGiXOzJd00ruvwl53H3JYWbDHdUVcGLTv7S
n1C52KEgFWQp/d6NIi0lHlsM1XjPoCZmVW3M0fHh6/KxdB2P71mZMLhUISQPcRsn
Y4Piiw6Ts0RmDxcRuE6oVfr/VT1dfkoensr3Mv3aViN8DYC8RFdBXn6RSOvsM10w
2W50W1kQI2OSbJJnLdIK+7f05xlEuRZxgYEjS2LP5RhBdKl+a+ORaj9OomJye4LM
ozJ2L5e1lQtzstuBJ5uwzN1lvBFrHudwH567NGHNmmqbo2jfHaHLkYA3BXm1vqrb
oFds3LDrktFkKovHnFVhLHSuNfbEtkfhaLE+RK+hQt6Inn/8LFmz3gXRQ11Jo3t0
ZPH5y7CEc1YCr1ORj06LgTMxDjUWA1wUbV3Smt/LJrljStK6auEC5dscq7+iugtJ
MiUNrSSAQkMfSapxcsmgyR9R97DiruS3wE/Ox43bYjV8akBMrL/pdJagyCladoZR
swLwLEm5kDYKyaSg7UYXt171f5jxcCHiRVv7+THIRqZ+fDRQTMqbizqHVr/W0LQe
pe9Onm+q4/rVx6s8R6dLYNLLV2vgw7Ji2KpVNk4h3gOV/7QtiHcz8LmgyiJG4xdz
p/YhK0NDVGnFVIlhkeXkoasxxKIyNuBbdrmqhyZw5P7wTYL0ZaCGeSfauBJgmEbd
QVTtA6XZ/WyOfPiygGkYqEw18pEUKpH7CiQ0rGazEUuEMqY+UXk8qKP+ZWxp6t7U
ovI4GR4OfAkB6dwekNtqP7yKtSUhZbz41T8mZpZNQUjM/SOSx5aH917U8MmJLCp7
sTwk7oItbjzxSF9cuZa0HZ+3Z0DFKu8u06ImWazMxGFsBjvbCa859aNW1dA3iFcZ
rtx0exzKIhQeqjzzks/kafjPQ9TvX0gdZgxyYobTkXUjgsMVoR/U/YIoe5X03fdV
tBb+LjT5FCNaA9Mtp6dWO9E4yVXeK2Qd5GOTj1GSfAivOeS6jbyL4O/nEMWFW4DV
/8SN93I4aRnFLfJjQx7qeloPeYhmlB3jf1FurWgWSz4QWzfI6sHs0ZyS6ZgkqRTB
Ib99VAsrsY0rfnUyAzFypY1H2xnMv+j7+yVRjSuCm8Mji83/35fRJLeNXk6iFQGz
3i+QiWsApoVDPmubFShGBC57ZLbYyUA8Ez7XDYWUghtijWT8gvWMndOKKfPHXp15
x9PGotV7jfGfA6OcOPn4VEdDi8W6xNsDXZJOFFOCbdv8IJ/pFrqto31L6OMclh3t
jVAujutAWjqb1x/1Um56QLMp2pogKY+tE7x2f2ob2bpRB35GUvNINFDtW9xqiKdj
tPI/C1FjAzw4Mp2WqCWb52RWhrM/UC0OBHVrk5ZPfVPO2YMgtm+Ys3bhtY4UOHXd
Usr5ke5FTAhIWIEoQBeBnyDVKrmR847+1I2UM5IOB1XoEADxptb2+ZfRHwUsOHKH
0eNPmvmuVvMoZyVEYu8vyNHqYwl3CXexbPDx8gaiTMqMDP0ULdWr1OML5FLhs5Nu
ydki6FDJL66kQP2VlPpkF7j7h8mfIJ9/qMA7Chkt4jLO/ova5yq1JS8b5rQQ02SS
+HUJweJkpA8cd2OAQZQFBDZ0PqRGd0y08P6qH/pZcqUcEYuzTwOHqbuUOjyRjUUb
D8RZeXZ3FJgNNHuPwTL6c72YZyF/n4cj2DxQ4xgN+tPtB3+6bMtnMd0KrQvwdg7V
6YWXiC3o32v3u6SyKZVACjvDr7vF2HnRG8hV03dd5Xa1X5dacMRA4m32NMztYLjY
pKC/gJ3t1lSbL3Q6zA27noSuMAIqXGg1GBQtAN5mOPCAGZ3wu4B1wZua7eTeLv6V
z0J98jTRhir49bq0SnkNHyZiJ80HV8qTDyfQNXEmUJp2Fqixqu8BOVEKEqReYtvL
usxkvekrQqGFuIimm7HqFX6trOtJTRYs/+APmgRFkyt+cf2r8zYxxSnzbVpk/TvG
+QaUemN3E0GJ1t9cfFqUMSRSmFKocgLOUdTLmO86xDbwSbS3VkBfDsk3HmSEVs7e
r062Wc0M1tkODq3RCPww9DR0VkH4c32pciCt5oiftTg0EHEf3Fi6JLUs4x3UczJN
plPUM3ZLZygbGwgAnD26sDHZIKiHLlbZB2I5U9/zT8yngmnB5mmKKP/UVjeFGm/h
EMrYM5KrjH0fSvKJc3UW34mJ7/SHjRA1nGy7KDhcFDqy336QOCchdFGtYEShE2cI
K20d18eltvit8WULnllblVAxsyUh/mlyZ+u0OjThKEOlgB+zXseIPH5uEbu54rLj
mJxgml7mFbbypVFA3IIIUIxVSZaQzcDIvQ+A4f1IkY7IAIevM9qvL9p5sWVPHonI
DHUZL8K6urVeZHeryJZ8KRe4cFoGlm7zOxviDJK35xbDAljXUluAeXKvZh8OFhSV
LxENE+ZVVceZlZSLgomKiq4PRckN6m3r6yhJnxw5npHT+IqqBiQ1ltF5a5gUxeQb
PbYxFJ1NfWLl8H7uKEt7rq5+XHLAoMuZZ8FVO1cTPHzNMsGo02ZsxcUett+HYSx/
mbp5XemSCU/qxiqF/uxcKGD7Uqtyh3NEMjcY3nDQdItCwbWa7khaHZ5DA2gXFK9T
fhTDQtsomolMwocodNKD+GRpVwOxIy9JniVkXYifrQIKtQTxhE8whttzHxdzviRt
6U/AzvZD3ZAqcJtj5Fkmjs4fwtwj5uSBTLIfHmaCxosM2mPCLBm3jyDRUy8TiVPx
V+bqjA7O1njnySkZNTS/g6qpw9dZSLWjxDjQPcrtV+flmkYHUkxog6QL/lqVpPku
Ms5a9OEupWwdf5G8nNHnLwyksy1eu8DtEKFUlT/hFbDo5im24vHf1OxNL+TA87nk
OM70qrFv01sN0G42fq/Jwkazicqn3DoS3Z5YE9zzBLRzDphkPuSL7DRMX8efGNdY
+zOHir76Svmw0uKWY/rvshB4sq3vc2skqGlbkISq/0UD2e6+fkGN6V/xaAiBKmg5
NTuuX7kL032BFy9kUGFS9rcuedNRsx5DRiR2n5RHHQgb+VjczAwJ956woIwmC/5J
u4loAhnyGUvL38nij3Q8r+Zr3vPFmIFi7dQjvwgMkQAK90ZpXzlYmZA/QHpMJI3v
mPJROXR3/cih/c7CPeUSohnNRQOGWDJQL/7qubi/AZeof2Ylyopj+gLkFFP01PJq
u3ZwKCNuWKiWVvGI7IY0KE4kSgjCB7ogkvMWBOwSwOyJE0+S4YJeFfWaRccaycDE
X1I1Osp06k0umo7byUMHVYuToshM2c2XsU6Uvs1n7XC1raLQhWey3onos1TbNFcM
b2Pc/8M30tCELq7jWBlqiit2wKRURvW8/VrRb76+dkVYe4eGtxlkZx2y+iPaNAKH
Fe+IXOIO8XM+bLNNXYbZjk3aazxooRSe/Rmsp/G8ScYhxxpypOQtx4GIvZYOvFnq
7Pvg5I9pLpAW+svROA/KhmoX6+fHI+++xCQDHO5XvneBRru5JGRBnpZM5bJsxcYu
A1S0SN6f2vUKWGzAgnHVfV/J6KOpMKSdJmVo1fpSaJusi7UHs2P9z9jOj+ZKwM5D
VNOJK3DhimyhPSfBwspKhHTIjZYXtdr0Bxf6NsEBVl9OhxMxXZ80/cQTOMTogdWJ
7X2HrnPl0JYBSGmmmi2ndjMl/m4GIA47r3cXO3f5zaX3rNClRB86+H/sQjOrSq9F
+Vzqc0O2PdwMZoQAdmTwGUjvTqaokzaOIVe4U6NStR4iO3W3V3Nih8JTWxvnXKt9
kC7BSRSf5Ypsal3356qcIaaSREzd8kczupJFUoV9BvEmIrcZCxTewzUWA5dPy9nq
v+NFGWDj3drhYiZaT5EIXgXS/My3NgEq8nvg+G86KCdtxEzWvdUdMogy8jtbCvgp
7TMK1Xyrj1XBdK9spTnlZQpRpsWtkxl8CG728Ku5nQmLIcqZvnCD11pTh6gFxeuC
gpqLXMaL0NvmtdPgf6RkDYSBsZHk/dkc4kVMcKq66KxyEE+YUJEzKCUnIF5lQL6t
oDKnRU+Xtvam+7jiulFy2OKdwkUJA9OTgPDCLJIRtzhuRUSjdSLT2Cr6rScOLDQK
A8WCYOoDx3R7yXueNlqNo5odJm2LUoMNnhaFmCdlURt3CRYBmOYsRq/TKiRYqHRo
DHkGJMVa+DTP+wPPdXeijRvVZLPB21a1Ym9cGXmUWNXLIkFCBXwktzO40bzV5jMG
vuhytdgC1PW66Cx0FZlnxvL4WmbbbDCFTPMJ/0IjA4r4dJ/m55Y7npsEud8Kxzv1
tpYBQ4QXqpFsqPH5LMlwNGAzJDnqf2FUb9han2HlPQdzFsWz2FH+PxmgW/1Z2i3V
QYbp2CV92wHjY9A1czm+1CYbxlpV0OG2ml2lBcK46yHfoOD0phR2ckKJLGQRK0NI
yKBBrLee5prSehX2Drgmq1hY3OzgqBgevVtrfPjFz9JlthHf1ubcsawhc56I8j12
0h3PhtBuzg3DxT0nASqfnOv6SeHJmCdzNQDKKqN1YY0vFchuTPDIBhCNyVjG8pdd
eSxaecRXRGz0g9PTkm/1XIp6mxc4oGt0rpl5q800EfSRps/AfDhb6/gbqqcTsABM
0Ti/CjKADDIlCl7uNo40xAhGfX3lbPZ0/CT2s0YFJcsZrNPl5J6sIEUeMAY56fP1
B4FbpmLSiSptz7F7yy9AhyoJ2QwQdaUZfcsryMqDtb7NpdLscygkDi6wN1BXgTva
Ksa4/cUcxawaeIjJmF++Qk+IUTQC/H3YGzMTZIskAEUfQrFuOd4HSTTo1Gtku8b/
aRH9K6MnNnNxTF1Ki7KyP1IE5txDoa2HJxJd5z4E4gSAID0dEnoRY6e/XJNKkSp+
M+MOhZTcb45moM3l4LS00JgQwhBo5hWKfljCX1Wxp/ef6M3017fmT0/ht5191Or1
BRIhjfjmbk8dWcHu13oBkteEqWDzKWSV0N50fammTEXbt7Ei4Sb0NIPgBee0Ctyq

//pragma protect end_data_block
//pragma protect digest_block
nddWY00UhUqbiWwdTsExaOU550c=
//pragma protect end_digest_block
//pragma protect end_protected
