`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
UCJYOBoKGDHrA/qY3GWHhpMF7eLzWE7bu88fx8Xxiq5okIz6QZPIayZ8G2e4FMhR
Eu6jxFhUbV+esYNe+PNEjfRJBLw56ryGbwvyr4gABjD/aI+d09EfjXSNKHGhGQWt
0Y0tSV2e5gl2p3LZPTNAQwB42XeM8z92jbo1P5UpjWk=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 10592), data_block
le8+bttZEqcXHAa2r2kEyNnvqSPK4v4eYjOZt1rizphrG9NoFBeFgf+8nxvKFRxz
h8ZlmCTC9NB7o66J32A/n+yhvTcnzUu4IlPOpGO7bJVkvFmJAcrL14il5QwI1nF4
adQ0X4zys0EaHOhLU3lCmXwWs5ddqV7I2Jt91l6SxE3s7NGyGLSzv1hzWtMMLUpd
tT/9lY38sUX/NhawyPGESv9ey3uVA7ZIHvVyh3bGYimkvCoxNwYNGskk/xx4PbvM
qei0SyUuXW/xxoR1Z2/lBkG4Uq++dyJMtrJ96acZ7fxBk6Q9T8KF6Z0C/i4exTsA
fJ7OIe5Mi7knVei9/fVO4NE/1oue59BR8KA4+CKZpWvBFIu7oOX/HMwf+2GOoLXb
9tB0r7PR8Fb2iJC0ofeeU+cgnt9cDsfTMvejUmD0WDFtujw6kiYaH9BE7ptu6oO/
3uFIxi3O7vQwgvvCOzKMvNSseaWD9AZclsG68p9UqHv69uu1y1Gc/nYa4p76j9YQ
DqbM1tWfwKSQV9RWjuSKWGsEpdttb7tCTbJCoyl8+VnmqhNCqbj0iJCuurnP1OGd
ArmBmKN6+Cma0sUC+uctB77t13Yu4Fm3eAyYViySyE5tcb2TaG3sQ+2MmLNRADPh
zOtY0CPeOmFC1YkmBwD6RgrIqqZy53X4SnecdD44ABLF6N7/pbWJh+5exh5MhFRu
BC/IC4AuuwfxlrDona3FBL2Hg9tT8JzFcqesdEnMA/2C13dfCTRl0CHPYRDmqeMd
/fzdGab7Nni1gmfmcF0Q8SGjyYlRcQNn7LCWHa05lT32Ug5D8dE9n/dKLV2hKg7t
EWrZDr5IJA7P9Ew5dn3CJ+uhweu0Abklr99yN1RMfSLjd+0pOWXdGIJpdA2OUOcR
fb4E79M7UK92EBK0xdbSbdsX4Kdj0R4YdVEcVnNUBHwMe8NzsinVlRMbMMSC//2P
XrTv/BJl6dgIzPJMSoHpYLw0tcQvQDm+9yZXtENj5H7iCnfyrrpK9p0Nzc1ETFUd
5eE0Mi/C5WNzEZOv1ca7iTWkYfQAmQYWh0MklFwwKzRWDybSDq6+wD4zeX1VRUyn
woN50zrHsG5D6a1RMmBQlBjiHU/hg8iQaO2szbHNeTIPZwrNhqaCeIJtt5xoQ907
uMKQZxQ8uONqxct+RECpsV27dkk1kWy1AKwKmVhnmn/2enNKR1qeQ7XvE5iEzngV
CFtvEUvhaeuj8UTvZC/CxSI+w0tmxYdMrstLmNI7q0C0nGuLKEyj+SC4DMwuawh4
jPSAqnEd7T8mTRSfLDwzd1pxzE+T+VUKtxM4f5Qmzn43H/wx1xgI/yPPiltGitDA
f+Dp4k4uWvQsvrfAqfGzsOzERUGG+VNqZ3B7uWcQeAateGQuM6JLhn2kWNicTXBZ
yotbnTHEk45OgbwZnmuSZxXtJ9ptq88Al2RDhIP1Kzmh4PoV8oipcW2Ee4QMyQ+Y
HcdY3Pgj1zk99BhcdgmRvXq6s2WnUE52kwHxp0gw8hKW+hEo8TGJAYBUjrHBnBq+
oFmgCN5Rfig+U6yzakPKkZiGP++mBPF2fZC0ve8M4zPw49RBDn52pm9/efAdkC3w
HPppMeVASYyEDZ8zfQ94VyaAfhhY8m/aHVABlJCvH4fruMwMUvxyfhjsSHRuayYQ
/WEyDsRHfcU81s8n21R7HQDbdorE5KTLbMsJt79iUyAGY8lvstaYvmEUkGMTIEYv
l3n+E8eHJdEWXKkTNuxM6sifMfFUOCOUZ5JlnP3bouNrvF3no6VWUWW8Ut3MhjwG
E2zMCoYA3X/poQqQT4n5K4SxeSNAvh8aUBrmFsuhgaYPPk4WjoOdquWYeYoWf8+b
qzRkFDcK1iNQypP+FOe07Vm34fR7jvjn0llyw89Y22VfbzR/tn23SNhmabb2XoTt
6LOsmyQ0la+ADQHhyDYDZPNXOUcLl8MuYY1/dpCp9eBnac7d+9jR9nggNRqDXfTG
UuDUdoFaQAO2CwC+QfCqHOX6sBpNmuRjI+KDkrYzvYnWv2Vv3i4wzuoVUspEE17k
5JoB+1bh2D30aIbwd5IJDTErbJvb4SOy0JF8GAyZSoflLd/syhqsG8ECVIt5r2Hj
GHJrWV908QgJZJhJ3w9ET3zCJVk2TqVpMwZjCQ4Ek96s0Oi7Bj2fcPzejbJamd2c
61Wy5fNZzKTwINleVBdDwd8jj1aD0Yb+KBxHJSlSCKwlz9vzDoykkU4VFyx/p/Ce
xJ1TL/kPX2ZoRM9+PXKBIOuMZzSib2+oms+bNlnbFy2m/LkIJq3KY5UukzxpglvY
ZK2mHqSIBGbR+twQhK2VfJXnfzOozHbdxI6PM7eEd2YJ9YsI2c68keCrOa048Q6f
IFs3Anbe1vzHxFwQAmhfdkGVvP8eIA8uJI8nnhOA3vJtADFUHGODaAiJ0FpwjixK
C72gCnnI8IZTvnktXG1v2QP2A9niKlMmJNb+UxDcX2uQZF9LiYq/hfZh7jCn46/B
e8jb7Qlv1pjv6EGRPCAx0NPZER3BL+aN5V7L4k5i+P2q0BNEiHRW4JXPopfZHdsq
uc+aeuaRRcqPgmGRIBc2XlMkGOXfwU5KQ3RQtN6DDZCkXK7/ajNM8XzWIJfm8aRV
2KWXtYLOEuV8FF2/jI6wEPpEEe4wYxFEweTvK247vmh2ttI3EFgxIUV6BPXf5cbO
aKpd8vp94oYAkzKcYzuXzm8N+E1+bdauVDbTOmFhEof2X8FmVilJj6VygngtHWxM
wDiPHx75xsM9CH5PJn1Q4vAonymRI7FKGhzXPJWk2PAMoaguBZKuc9DOOXmSr55O
tf/jh91vJp51Ehw//lE68DW9SiaI7HuM8PHgM+MNCDfTRLSzQ1W5mCGFvudMKgjt
7hFCXzMVolXp2YwPZ6hUHPo8jvqgnZvUaaU4Dh1nbGWhXPzeLr9YXV/JKuJ+o0W7
kUk/15Nk9n+EQhg5i68jKx6RHDHR154w+kUykxi0CoQUla3qPFnEX5KBbGto+3ef
Ubc/OQfFeA5B952V5zjwAFujHb3JzQZr/sdI+evMN6S+4XiFtir8fNc8/1AY0lhx
95zUs9EuafjiR10KsGdnyQxjfWnLgkQlB89fOE1qucy3/GNu8XXwq7ccQ95mhzBK
+1pIgkubxCmxnZP5/fUOpFqUa+Jkd2CE7tZanw/8TOScs0mVuWWsNUlXwqrc6kPz
Vj+YKx4mJbZt7XzEWlb4x+TO/FIY/FvhfEiLnpTe6baMv2FmcVMjqvs9l6V2+yQ5
dwdTD4UhwesEKnKGl2n4seklBFzvLzyAvEBR2qsH1xuYsy1tG4yEGuT9XvWX5y6y
MlP0tPm6ruoRxU7O++udZ1yQCE+lkk9fFzXV+hrsItgG0+1yR/+n6MPGHpdSAQDB
WD88tjml4pgGWKV5zfW5YRfUQKZls5G+GFWc4tq5CkNQDWOTH5yuTizJJXoXh5Pp
srk7sV8ZHbxqZodIn4tXMUzs81nrYHlOQd9R8l42+M86AysX8VDJ9DXepuo3fqjH
TuwmtAThZap7TC57pTr66vdrBcTZj1WN+HAa3Aub5GrnEmZZPet4b4aFDf/gL8By
Eh2M17ZTt1lY1q8ZX2xCquu77hAQ1MLRtus7MPQxi/nClo0IfYEttz4+lKZ0OcL3
W71EH9/pbQ3qjC+u8Al397bf1z0M0FB5Vg0xHa99VJONQFXJVnNSfVgVgD/O3r5/
s2HBkuTYs3hffZIycIECGfIrZ9CSU1RwY1+bBx4GqdTC9aETRLOu38ZTd//Se8GH
dDEAKFF++EwAlxc0UP971cH79dTna+w0cF+Lpn5Jyeo1nkqxQ3erOPQrRbTEzKvc
6++2CCOff8JDRWOwtoOmdxCuNfUUzOnn5ws66o1V+PTu/icwsmCkc8qAiJgx9g8o
8ceSzP4XcZW7prm/YC4a+51Fd5Jd1RNb8zEV29HFKNDyYLmXJoChYv0AtZqlNBKk
4CdHsE6rXFrL6vvf9UWuZeRzI3zTm/BZTL1RguuXTTMuEyqRhtjBPBi+oC5sFmOB
FYEO0na5NyuGuXcYSqsKoC9WceuV/E1w1SrvdC/iu30PEIBqqa44CIT8JsOHqKEI
IQjzmp1KpCyBk4EA1osvy2UqsmA3axFgmlyTVslj2IwwZUQrBf/RdwT+D1317cgp
xndkHfBJGm5AX5B14106cmTvLBZixNbv42m42++ZNjFW1fYoXpCyvJGIq2Bossyg
V+o/mlY3zvpoTaaTmb3EePfHVQoyXme8BYmzfZizz/8eG0pNG1g1NCkxRF/Q+/al
Ed+0U1fe3EJLwxxHpe3HzFlW00ONaFR/nRuir3oWwB/Ba9IOs0tYZzo+BD1DB4LW
xpgqXlFIZyw4us6l8GK3/ZpyuCUAQXZeWA0SkXz+ff6INzc/7oUFY6I3lfiTKd+A
TvvC/jq1WaO9fgzZI1LWXoKZwu1UMBb6v7kEBf6ss4Ommx39k8UFuVZ9sH13FByj
HNM6ya0vJNjLqDGqn9qy/bBzZ/KJFVeklZVLd3HmtW66xz8tmPjmkRbCsscK/oT8
iUqOizlr37Ba2fPyM38Eka7UV56XZHg5ccvCwWoVwMCN7nMfNeQzLl9SoFsFYRVA
UNZut7R9UXlHX4TdwiXzHFRu+ab77DPF4I0c9O6Qpe4NsAgg26ZkV4psUlUklWe4
u085UazUR2ETj71YkOS3pjxah6lBEOHNxJvoWyxqaVia67+9wOedKONd83mEDIJ2
YmmqjONT7ntsVihqFmiL5eqLESS/VaU0HNzROSTRRBxQ36fcPYRylPS6wWsAiFO3
MxSfRsclptRuYmy/OVCTADH/QGIWWDnM5Zh3KQkOw/5NrQq81fcBWWrq3qpqEM48
v/jBXQmrkkAKK2L+viHkUNkQoxV/pDUj6VFHVCyNPoPgEcYJqhXn/DqBNnPIAg9s
OWNXIlYGbvtt6cKitdssqLa9MEALiLp8uSwO3dDxj+AXWOgp+/HX1wGx30BvaPup
46RvfJ/knQDmLcbL6ZFp/RmZ9NEXiep6RmconCxzXGpZvrHTzj8XFet6hc3pugfx
rwQ0ogkqL1/e+3bjlLwGRD04xlYbVwsOO3wFf6cG2MLjsSrNAQ9MAhhQ4sqSHapb
BAI+w4vVasDaejl48oCo19Yti08RxR8zw87JRFUJJIaNgTWrs2UBkfApx6cII/kT
lC+yZlYvbiCKviZV9tfsD509cHQ2URjzc13I4XF14hA/nQMnbV1T+bkXnH28NrQH
NIpeQKgxtZbNp/AnzNJV6p08nZv17XdC/jOV5Zk8tH3r2WlCnofXO6LmdRis8aIq
IU+yVqWB8vn74DhuSFaWWH2xzp4CAz29/2/p6zAyQZ19eICLgpqN3Ce5JI7rmwol
KY99weYDVP3tEGzYw02TYH+w7Wv55+JFbhAPGIAAGQoXz7oXlS9r+pFmX5fSj5A3
XtZrghYFZIaKiaj91/zMkFfICFc+6HGqOI/fD9R8AMB5qkDTbBs8w+Nrm1CHZ/8Q
EJUdssZgB32E3QsWJm/NXyqwEXqqfg8xq8aRD5RocBg4B0PED18nKvo2UpQN17Fd
5lE0BZJmFRd29nqsmQ433q8gv1gBE+dXiv7f+E52Xphki0BqJ3yFqckhttWSsaqb
BX/uOWFRm+BAiuv5WWuF+fOPqL9l6125hI/JkJflPQ7afY3FrsUwONNnMwyhJfdw
KZGUXh9Nm+PINOkx3tTSUjZfvtJpI4ZcimxiWhd1PvvTnRRu3W4Ei+SKEXY4t6Mf
SOEdNONTJMiFHvrLWOuf2hFJQtXKOzv8t5rXaLIOD4fiv/7ufW8gnL+R/4O7FvQw
d8GsDsCHLwBqR7+w0F24GNYSEjRUuNlS8/1T3wqh1WDXLFO00IC8ih+ln/h7651z
cTdvzDjkHzYGP5rvgAZ2c9JqPAlrciJ0cp38CDuOGOHkqqe+6Z0/HjSJusbsoKz2
O6iu0Icmpi0CMERdrYfl4CG9E75jYipVKtkvfZgA9tFXjHRZVC12FvU08jqAULkT
sLW3VaDb/FeKtgm61aFyMG11aOg8D0Qswdp/4PviAr4i8av9unRkaSC8ajPuTRJG
vc18iJ218dRLdmptn7Z3Qmo4NAuZMJXudqk8KkdLtPJyFEcfDs9JWkhIzK7qxmQO
m0P9YrjIZ0pMh8AO6R/4ByUMlMNt02ftzmbLC2/w7lPWehM1LYyPQtbkcvkiSbZS
OBPRtRmTgU7CbRa926jRdy3p++k0KzwweMtjzeRlsDyCpscev5IPRc0SQsGIT3CW
6hBEUV71Il8hy3fuxPV26qRmctIFrp/efrWFQwCEUfZUms+rVpYkAdsdiF9U88rL
uYCIc/BY4Yv85Xy7Dvoj7eIozzXAVDKWVt6D8vsayk6iyB/xeO1055bWXI8PDuyg
rYK/IWD9fj+bLAYx/LRUVSUcv9L791F+VYkukGvTpyUcV4hnyldOPsOtZXTZUmdV
P4kBBqKwXyRg/Yk2BRcQ0n9HKM9isaq5VhIqNBrI5Dx+jQh2XZtyOvCLT5p1wzsF
Dp3lBuw1chAWR8etrnfuUt7xvQ4rcHUh8Hv37MNmNvikeouiiyLIvn0Fpoaw2IQE
jh8UL+ws0QJRf4ztyJlk2h9ZwkSUbECkVT3COXPojAf27dKSfDx1Og2LszrQyh9r
ZWcsQtAAGB/XzhnsIpTasxbWjREA9mqRm9xo8VQfz8BVpEnUnxKXK1Tq/DGTdWFp
aND0WbqNhotFviBLH6UwAH5Z1H3WEHEpn2L4EB8fa033qwoSRZkb+TVJW/VdJc7p
cUC/3HLwNBTaagqJzLSkZTJb2Gjt7EPa/ipxflcroNBxx7gn4d65uqirEtmb7Gq+
vWKS0iwTlUI5ZidC+gM11tPfGSfj2ciB40JGloldAAXCy8v5i8OiUoSdtaL5CTMy
C4V9PT7K3WJCPo/AZ32g/zxKxh5TKxlViwLOXYuT9cSSQ+addxRyF7UYr7mTKh3h
0ciLMghySFG5iWDt4XLGgtnFn/B7IOEeq/9/5Ts5Ufz+GwSvolvwPP7htIR6mDVK
KStryrEbr0SLbBOSyt+REywNAV3BfTqQMmgL4XJ4T2LyuSH8PoNPYhVoU/NmX9Ol
iLi6ZkbYT+n+rKR54VSR37vj3cHXgzAlUDKZCVvOqo+T+6BxLlV5Bg+lxbacqHEb
L1RkQR7HJFeHnq5cLWRVJhVRMc8H8aomjXTxz7MJzFsAnFnfNkIkiUmWzCE1vvro
lfQUGoBsmdD2qkY0YlQWLSb0kCKG9jEjSAU4kqRiYaz+dp4PI1pNYAQVltCsPyUg
Fh6kDsmPqUtlsnn5yUgYCfZOkKZHZItF2K3Ia2Oa3rCjPJUuHCTI8ec79rYMR2tH
lTNsuIphu+kPFYco1OYI0g7jbuL29YkOtPzo17ZitZfeowRgnQa5vH3M8oHvG2eA
odvd3f0VtRNFvu2VwmY0y29eWPEhzuHhbUJSGX5cQmPzxdssus8oR3VU9Rrj55+W
74n4QLc8wsR1GnqH1FzPSpTOxPEOXVr4qal9OflHbL5CQqvXx4in7rq/HmY6UI8Z
IhC44vehqyUVpgvC0q/RGSEP1Bzbkdh6cstpgWY3r9gIzFLDW2173VcoGWZmrkPf
0ru8TPkqTd66Le9xYUb7p9fP5AfRT1ONPsx//8ZAZPK2AmTaHX705B/4cx/DJpNH
ln2XSznAtOSXm1W9V6Wj9UiFt8mNihRZ1mKtZ5pdUHSxPo/qAdZAClMe+DEZvQIC
nJkijW28nf5KD+YLZjgIKGCdWWDvOdklSZpNbHiJnZI9NMH++Y2Qypj5WnQ6LhZ/
wJjiv3mG4dFmg4FjtF1Q+gY8Or5mYl+aJr/5G04SxEI5CiNXkDuqqvhdl5i92KGb
bBec762Doe3chJfuVkvtqKdN3BIF8vLu0fdmotPBsct2LpsjZp9uhd8WWjeKvaP/
ooX3iaePd2XvGdYJUo17OMXOsYCm4cf/thvjlYIA96Lo9sg5Xcpr9QNIvV0DLbiv
y5JCmr7IlJhDdHRcrvc11peEu4ohtGV8VhlPaEJuSuSf0PyK0I1GEMGUDHakgwQA
KvqMQGXrh1zmmxt10FjkFb/esGRCBZW1Ic7+hewGIv7Sspp6x2fm+EOUIdaQbQuG
Q0f7xwfNtTHFZgGxrHAbMAbho71JQHD6+ZE4AfEriacjmHDJ/jS+f1pqSuwBiMgy
+u5sqJLD7TTcTgtwjfLXwhaKvqZJNrKnzcptRxoaoYCrJPBU86EjWg+DuqL7LurD
vV3+Qfg6Skl49zmZYrdNXWoO5PuvOvlvHqiEkrwnyr4L//v8rzGWx6XvP4QasIcP
DXXP3b2B5Ct3sVtYSyBTrYsTDBa/3YjMaLRgwxxTpDWWYTgjkdOF6r6lhHCu9bZr
M/e6s5ooG3LdWL25YupTn8Y7QDN61i4ZWdshRIqpwCXHQk6OU8+InQpdd9Sv1Xp4
iqTEb+mnIYcV5RZo7AnmI8Fu4i9/qDJu8X65CDAthc9IB98+VccjECTqq7jV5zvX
UzKnOqg+Ll5655pTaDgZRKNrsb00aqOUGgHNXC+CB8I4vk1v571msUXWT2Y2xeqe
vED3/qbZBspLy8PxYG+oJK56/hRbZJFV9KXwOveJEUDmvfZ/3WpDn9pLCYv6yPBo
e5m0RY/WAgdKyZpM0eHd0Pvk0w9KdRwy9Fi+pwtRZkOe/aK2M8hc45sbSv0S4Pot
HxQm9oHEp53S04A74s8ULzqpaAMwXVQNjivOwy+HK2nGtu7hRluU/OQ/4hl7NR/A
Frzbxw0o4dXKpZUv/3suDYu1DrZwnHx50Yawj6RjP582ZBkJQwODsMw7dUUAT1iY
ba5X4lmlfVfZqbLFtsUAfalSZe4n7f+cTYNWOmsdjYUkxdqzrWntDRv90tUd1G6O
S8c/0Hfc1N6BLpWOs6iiCIAqpKjqSi0Pqo5pxZYTh5n9Yr4R6OtFYX5gs/ZzX+np
xFIaf3pOf+xC32ermkmLud2OT6vd7n/dbgXFcLCZntwIkKVk8TH8DnPcui0PirsD
744Sn3a02RmA59kZymjtmw8Slfeom/LLul4yNawapNfOCKY8rGePSFOWq+KMTjDV
z6L2qTp6to8ZYs11SjphejTgtICn2tqXYZzqgQrtl0d+pomzjj+5qjx6opHFpU5e
oeDnkC6EvHIozHqDLGAR2mwGQRTngo8AwOy+QwHwZM7kNqycBI4cOGUXXGIf8r0M
mIGInvINkaJxiqNY3rlsQIB1JKZwadh50YNLb3zeJ6FNjIqbD8AXl3r8K0kr8tJO
U8ZWBlLv+07wcGt6nlUMC1r696r1z73OIQfcCQUohZjfFf9cC9Lw6+3LHPMuuXSt
/MHpMgaRvAwn/kQ3ZmwXtWEZxX9u5b14Tkp8L3y9uyG+1mVPjsIYzAVho30G6WYM
faebxS2tSue++XxSMEi/vXZFiZi579FKuoPJeO2snzNEafdoPP7CHAzqs7zo3Q7k
irrZtZXm++OqacxTZ4CFipUZDrX92ENlIoyIy65jl3HZ1CkILSSmY0i+54mYrKaS
6mfCYe6HXgpOQGb6JShRDePYBNDwNBfoWyASECbqts669/nnRUQH+OClVOLi/JGT
dcvg5domgaXkMo+GjTAn+c1KmCECE2j+gF6698d5ZPIi4zjgtABhKwIS/LcNdHHa
EY3RJyrPD1khOLWA8PjsP+IlwiVEIN95miqgbZpFsZIiYUUHWGfJM5mrmO85/R4X
pRovf3TEOJjBXX2Gm3RA68RGdSJ09Su9rzXGKCMC8brzUyOX7cgVS1eOrZOoSryc
U2aLth5bTb9IXOG78O+rlGYaS1bnODJ8LsyZQEqGlrkpDMRXouvEuUYZRNTItilB
l9fpE3nM4N8AAzs+UPx84R4iumBx63Z520tTvzcRMXrAAjFniv7SazfqtEkNqHmG
vQR0fhNPigsjOyuXrdE7TSzZulKMCBA8qDXDWl3Ut8+t/q8p92nLobHI/5OZegrC
VDswcaOJx8Z8fpNbHPwVQ57rt8Ek6VDqKIIdbq8T5WrdXS6H4Uu2zMDWqpcrkNJb
N+gSTwILH23SONwE6WbIP+EqthkeubMv+9yzGY/ufEMzJcIhVf1FSrPaFBvhb+me
8SlUaTE/cA0KvxxniHIdWiinRRuDqTiXEZcqzWU3mIlk9z3FqUZA1agObjf72OiG
ekg4YSM8h1sl8sgeAonUHjw+K1VaoFiAc/HurnNmdnb4huDuAyUSdoSRI5k6x2On
jHSb2qOq28S+54bU2qlmJOUFrx8hArrZCKnm6bvCvomR2JOZRNb85oyduVC5X37m
Xnfsio8PIJzLjuAtrY4wnN4V/0j5pGySAPSwCB+K08pp8Cjn1mhLn/k1Kpb91dyf
Nq4p06LhqizsL05g7TnoLKy/gaHiL+lP1LySkcim9pxvRg1De1eV4V9WGT8BM5j7
EEooUy0U0N7H5zm4AKoqNNWoAbKFJcP/zhsgH6cK4RB5uONTljhocYojr4NrKpqf
dJLWms0Re46Ewwz1olRQAcySb52yYt00+CR4xbqYC8V/i5jSjC7IlhF06NiEHF6h
f8uZ6CvATD1jpxe/FgDbZhFzHVtsZt59YCJUXSnG3j5+4YsRzZSVXv+bc00DFb97
zl3TW4qkl3QQWkhzpA2OPffNIl5FaJlOgq119X6N9e6b8GarNOiC6rzMs+85KPEH
Hj782LtJ0Uw/HcBhLy6+RtkkG5eBi6K5ZERPFVZClWOWwkuzE/WaVth/Gz3rjuqT
ZKk+JsQaxJepwSKkJwdouIMY7hHP8dSDdkRo0h9fQNH8h/Qx2dn1b4ColKwb351x
Pwb4N4TCiPPBn1yfrSLg+AXjzT1wjHL9yYG9RTblPPGrJMWD7/JS7EvkIiQzjSV9
tbPUT8JwjBlU1eseTHQXn7q+aEQkJKkAdcosuQXAJ0Mgvy/2rkFC2RC4p8trbQ23
YVULJmnD8sTldCgnBkqMzBFbRC2N7r+ksqRi3dadThAW7LPuWpHnJf4DXafBaovh
oIG9vioqMb32IAbByxw4cMEJz97ZatDVDjiBAp4r0riPb8Om+9HeNZJOgY1pDmEm
mw8l81YaalHr4Zufe1MsOChqagAbmiAFG6fFTEVATdE5wxXL+Q58k40TuG2VRbn6
coHoD+y9tJ/VqSyeZ8ME/iL3PkBIu9STUkFH6P0qLxu9xbRwrgX6CDpUsYpAHwCl
nzZGFY9QGuW7kRJac+IZtNhsHf9v01tPYY5XPAeZXaF+CwF7H05fMLbYI/EkO5Oz
qcGT4ooIKiW90RXpg9DNaN0yJ7EEqyQnBeMPqjl15MsPyBc0IpREK/ji6fbmS/O3
sK8znpSQ0I1dzIEiNS2s48GvcyGs8KI5Jj5bP0U/2H8vKO0RslGxyOkl5J2dimYo
yWOYtFXqnFFPJn5gFEIBePfJ7Bx2b43iatKU485noFiIn70f1oGOV806sgLLiuMh
lY0iNo8tZALqswuTxmIllsjCTXBU/2bVq70m1hqqdRxjf2b4yvUbWGFdIClJYoTm
/qu68g9eZMeV74v2aVpqg+KFnFD84VOpM5OCxAwy0U9I0+um0RfBWFlOmYG/28Jj
Pu6h9Nl3LwqQnu02ig1nS3nLVRsFFgbjem7dTBOD1dMpc2Pu1QD8M1N4GIWMeFFQ
ZmEhXAlavgmCNRCzrm8RnZopWzIwayuqLUfelxoFsTZ4bUMgWhmep8LfhyN2eEdr
CGc+4+cv8j36MyC3pw5Vk/8R6TFEZ+Qk/ZVgFiYAScSv/zVWjfmE0EgBM0aJiKPN
R18/y8VWFoeCrzonvVZRnac0YKMcU0y6L9did5rLPJsIp1bNuTOlw7u/Msf3vQCq
pvvMl91bQXY5F6ydxVPlIQ0BSmcmmwntbaeUcsaVH9SEsm+ZD6uBGww2lUiHrKPc
mqJ6B9U4lvzGDid+D62Ai83pbeMqThVrGQHAw0AUpTrSNV2z2ECe5dE+aWkHcJvq
aNXetz7fuE3ySknq7ZxR2h9mH3JVFgHCmUr0+oWI7ulF+AAOOv5SYVZgxwCLD/ol
d6/9mEYKAyL9Mc69+0QeQuND4fSA1XGDM1k/WTpfpK10ye0lda43ucVRu3U44ZIJ
PN6+ih/E9dIMPtOppqupSfzPi5SrqeOaQOx8voIcEP3Xy0mqmaDk8wFL+6Bvdc+V
7lPik1zay14bM7qXTQNVf0kD7Lh/cSUmaxdxut5wihKZK0n4p8vWb4pE5gZcaX4T
nq7sx4366HP8qBeTStBf5y1JQd39TQLgKpAG4HSChY3IRryzImUDVgb0bS8LN2WZ
9bYrLSfXwP9ANEqk8lYVHC00hVNUTA/f5Ax+uqs2LpG2UCm49PbB92FTr7djQHgE
5Sh83YPm61tKE/p72HK23ecf3tp2hQIYlQY2Dq5urov5E1x4/trhCnzyrANtUJpn
/cLy52hZcmNrZ911syslP7xlW60OTTbX2nbwWJPyi4W1hCw8Yr7gdzX5/jWqPY7f
9OQ/c7QQf8Zm/3Gh/yltm+jZPFAq9VAo8Gxq4Y8iEDVJReuRW6OFqIVfMLkWzm1y
227rm7u+b4tJFM0daNAhHGnDf6P6tvCZjq1y7x9BJGrSFCAP8G/ELsnl3dL4YdWZ
xSUMNnikq38feDGVYtBQKVLbaTvHscQrHGfdsGhR9sfvakviof1P0GN1undWrEkN
V3CM2YaA2Z6VqmTaqKdKwSIZTgGX+hmdAd2iph+jpGczMCPAwhvXL0wKld3Nfc++
YvyQU1fgiTY9j9HTvTQSEy6OANhP7JlS1MmfOouYums/jKorn4nDcLOweJbsEvp+
ln4sgOBOVOIaZxYhV0NiDsxx9jSj4hBI5L7OVPB+LXUqiNwIVzh//Cul/DZyC1fP
20L2TgTycrVfABcisfbZbXeqzvi/5XgHkLA5jpAOYsCLnS1H8+ofKtuC+r5Y1cvx
fFPEZX2zpZvEAdwVh5Q/m/jQLLrmmpXnTUNBCXMGiWyaPvk12baIF59dy2URUzjD
SonBFFdWW6nPgntB4W/U0vmkHHvxM2Ja34PTjxPVPglV+MyqmlAhrpY5Qu6tgWJq
laSSmr+veRqDW7r/avkMXT7lIWIHwrZr/IP3Ydc4AxrntGUvPSeRJj0ctcQIGwqj
m2AIZcI/MDM+38nFfCA+tcDOPkVvwjlx6Iq6aSyBsFJbo6XHSuxwUF7rWcMvj+fP
a8CUu6TVLBp98lKKRqunAvF/5q8biOHxExKJElcJ2xv1XQvwZ5oTpL8AdiXsvHrw
fHBzQPuJGZI6d200OFRVZep2qHzHcwiQNwnYMPn4QFM6eaTC492UPbxZMpyA6LJE
MvWPfYtOjXIyr80AI4tDoJf9GXtDdOrjEUxwwMzl9dB9Rhl7sTT5lt/GOENSskqG
KS7ykJGPtnlZEwzQgYN1YYydJ5iLY44naS/jPBB1h8SUha+5Ho7++l4cdu5ctLbe
cuzZ27bbrNqKwBPNFpnLpCoqiOJ63orAmlb+dmCSowBH3EH/3Tl2vn2wwtB8YJoS
wF1khgtM2l3iSZ4IXQrzcZo5QLvJjf5yq9aK+4bVU1E0rLeCiQEvo1ganfTU12xi
kFH/XW5T9Fqog+IgAC5rCWOAr9ivZyw8+a6ZzpxtO//WIBMd1+fQUkDzPlnMCl+A
UYeqRkaeM2DuRkbrR5TvGU7xlKFb4fDopsau4EexjUHzfLDlpPRVEnsMlnEDRiRk
bKrntTLfckobRdzLzCY3j6YPxmrYI2iWWau2eNnDY3s4YqmcVvq112gk95leA/tF
Z5Qu2DIpHwfZ0kPouOpSR2R3BhCh/K9gVl7Ck8WwdzWXYbSY8GPlgevP96CE6ZiY
vi7DGRjfNJ3eQnFYYyBVHKR7XnxZE5YJQFrze/P328ApmT2KTntf7JFVt3M89E1D
8cQ4rDEnmOHQWhBhhUnIqNFxTvtiR5y29lSzVkRiusox+JtTIHrhCv68C/DSFl67
3nPIQLnMUevTMHEBP7LWl6lupdXf4W7uq3nZXK3FL5F4Ybd1uwtaj9dpeOIlDhqw
DQb3J0uouYbPMlWTkm6pFxzXIKWMDbvTOBf2BfpbXbFMxmIw7HxmbhqLbbVtFltn
23RZtkCjeRPFWK+pEFStJwWC7iCsSKcX4NFa4Y3p/CM=
`pragma protect end_protected
