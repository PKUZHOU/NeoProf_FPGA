// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
cWrOuKTtnNIVJeDhUalOXhsbbVgq3s93rv7gGTZZBvN5gywCeSAOfKFyBEKRrjnmE+AccMxve2Kw
n7THr7Z/sMI8Kd/zWV6nGnNOv+l74vTfsdSPRqLkYKOkWHz6FkktcsSAlvAgnR1NGYdFVE586l4h
f4ZDit7sSdVuKFXLOIBkJDGo3Zr+Zr7v4Gw3bGrJWX7EjS7x3cjgcUZBAJSD50WJbTpEAWLDhzvI
R9VTF55/jTVz6Kh+dlDLKaU1+QvTLPSo0lHB8p1krS/Y3npAlX6Bu5D0k51ijmKr8jhcR0DRtU8I
JIFzcu/V/b7/i8kTJP5uG+SrI9V8QQoBB1bILw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 10336)
bn8jHqtWR338cjewAR1UFXGOx8nOFskttaKI4sO/MksH+O2bEv704EaM9rCQB/VUMVSjFZIQFU1d
RzKUrLvVg7LvpDQUmY43UanvM3KqrbMew0atFQ29HG8FOONx6IojEq0zeuOkx3V1KFw5fYKFLPUz
clnxO7xQh8dqLBkAj7bEsmlrWdf7S68cuPo07EYG31GCChU6dZ1CWDGMpGBT2Nxqcrn0/21N5Lsn
EUBdotpBkQY3VhiMXf1gQbXcHygkJTs1Cy9n6jb+1bwCVt1bk4o09C7azoFcCLvnrPyknS5XEsTJ
HaBOFjnNzcZeyvVXu25rp0HBb7x7+XZvgxx6CuDXlQPzOkqhj0MHXYClvZGg40+CJ6byfO/PQLrV
SGnfXu0bUm9k5Ifr7RgFjkIJLnuJ7BZ/Ix4BM2SzBSyTf1MpIKX3ycI3lKksSJjY+lDy/0xASXpd
3X7HKWQwxBNp6wssGfJdbe1x8YqsBnHU1hQdXRwNmgeKqGc8wQViSbzh4ink27vgdQxLq8jKLyLh
GswPRxjz4jYZGBYOZm4GYBhEbGkedQ8xcU042Oq/wYTStR9ByfezXbUh3ppMpoOQ78JcOtqoKiE0
lP46w30FuEPNv0TIp+2Bd0ITsWnSgCymgNotm3b9MHxZmguj43aGZfa42DGybr5+BFFQb6cvDyoF
cun3EItoc9mg/KNMLj5Dyp5gcFb4y6wTwXYzvnW+UxlDaSisPpk94Yg5exp1n8Tc6I/btFR0hNpb
yGNsW7+CUzJgAaWqoFtps1INUmTC2Qr2wEXRkHTa9ySEnAD7YBuVzhtwS5cojF7yUJtQ1OLbfnTH
iQW4T51nSoaONSLWdbxDXZggr98xFXOhtuKF8/A9a/Gzod1wafGJvm+Uz/mU16k/aBR0EXHLG19U
KDCSM3H5G5esnXKFdiww+qqsiWhvRg9KoD8lDag2cGAMJT1oe0cWKIRUo+yQZ7tK24zZFHeXMD4D
A0R70oFsRZRgsV/rpStPRNwElTGFPyOFk7M89n/azv4mfFx35pbLj+iDX1AHd2o/QtuWcUSP6CVc
yHY9r44vZvZgXl0zaeHYmeMSbasK/eB4LrNheTqO+ibXnbIwuaL7q0qp4NdnYDcqqIkLA4qASFh4
x9Ncevnt2RhRiZs5Qf9rx6xFnLSb5ftqEuH9Z5y0+vJBRsxMcpsWT+0JCxTlvAHkdkFPZXUHWFJL
RV17vSpnLG2XySSRhCgLMdu+2QUjXnFMPcK1H2QQPeKsCSBXzOnhfCPj8sm6VtE7cpzdNU8aIp0z
VknhIdcEFBREPBx+8izX7alJeGsas1K5nXtAE8iApEFaI8kghWpWhJMFNoJM03UKjEGoNYleK59+
J3KGVfYy/+NDNca7202xcf5Xs1lZ9G3nmxbHNEsoKva99NIo+qRQMteWFw5PEnyPt4OJmL3wjmsF
SExxbD+SpucjyENUS+Swbl8VoD9Bm1MmLlgMhF7FKiMh3lCbhpmIAVFIkfiV0JWOOLPjQwIIWluh
h6kP0Z9EDh2rq07za0lyqIYBPQT2nukn+UADuzzeuwBhTKpkazDg2g7s86P8Hx2RCST359jkrOuy
+RaQz0aSQAjcsZnukxgDa4lni5Kh6oIDkJT1J3Ea9xtKINVf+TqJ7hEsF4C1jU0Jwr9WchbZ0EXY
EI/qTMLNeFUomtB96Mgn/GO3AvMOceMZArCeJqPcAIP5SAclDlE91dCd4MZZ0fr32LLUA0HyFRf3
G8o/aCFt43L+4V3Vqg1deTT3CraUUApDFntd2llRkJN7BDb+enfppmp/sTPr4Qogb0v0ctbGKrHe
sx0Jr7ePj38R+GP4Hdvw7qyQfOisLESV4FHZ5V4SY8lOk1XsO/fMfu5ybTNmI4AWCzne1/yEBXk+
QvV0C1ZtYZSB6/dtlRbcIHpTZUUWn+BUXgXPNuVUv5ESVER4R/5dakh++bfagiJLUMlV+BgWjiEC
shynwJS/ky+2MH421eFj+XaJoQnrLhJU7p5vGQuMS+kHn9z4BS7gqAoijqsKDwwHb+SbMyi7Vbl+
7sLP/wrNXVPAmxfVB61u8lrbcIK8zPIZ4gqkpifdmasbHzDQjzM1NCnJslAYwYfci4xWxB2kmGvQ
TqQ/XoE4I5TOZvXtU19Q/sFv0AsLSKml6U+pP8BfhjVLUY1AXj00jM+YqSFOJ0Gc0XFjn/GnMXJE
DI9/N8Njeal2YMGr6hI8OWscwoWvAfALbH37X6T06gGaUsRzCB29RehRCcCFFTTFFHfF1Wu6YW9r
lL3kzo7B3WYIRXZC1IpkwMpXKQhe3sMqNDw8zHpEfkvqrrBbFicgHDZAtj60p8v+wjhKL5a0a0Z4
eTm1Rs3QHw31WkEznNnQ8VLo1HxQtXg1FmBIKR4oSADntsQS3OMMJdybYEObFirLBy1GOdZKs2NB
kxbdwIpb4KxpXOD7BYLixwDSbI+2QnTc2jEP3FMzdH3FVsI536J1MsE9lEvYJ9647uyB828ifdbX
l00gS0kZMkS+qYCCL2NpjftuIZAejQFb7Zkw0wMeUGgcqaVnOwXim8A3X7vawlkvMGULXSikMHsO
C3zGpZ2+VaWpvgZZmOoLlwdr/a4mZCoqWpgsQ9zbbLWc+KaBRcy3qVF1ECw2+HfmglzYznoVWC7Y
qISI/q/Np/KURi5WL5LInhgLXBqg/0MfcXWIpGx2a91gH3BsfTus4xi5D0g7M0kHP9g4e1s7D4Gs
oQ3YbvhBn6jq1Ve75aZGqHsnBCo8KTqB5S8VXkoqmErg/bNQjOHuMFQbQfvJkay6GXeqiIcoLFi0
+IO941x7KrCw6WqI7sL3feBHWkkfCU05vBygc5bLM+lUdhYcfZR+NHK9ipDrhk40jvPFdqHciLvf
OZvPgR6GBrF+IPH6xnuAUU6fgpOuaPxLWZkBQwcLdSkuQmed8HDeAWhLv3DIisiZItV0EkAmCYdv
YEiPro90250O83++tGvXSf56VIma5yy22mtxNDBSyjPO3V6ciONnnWXNso+oz+2q908QSNS4oD7k
vrIkgoKOIBxvOmfhONSQo5vwmaJtBCWWHlbqhYvSlk+CKBr69lQZEq4mIyFJxM29je5mxs7IA51c
ZhbXvTkl5nLQ10TuPSp0qq94lNZMrkQK9mKg7kfIe4+LJ85cTiKoC0/UwyeTiX4cfGFG9WL0oovH
F0nIKr+znIURmBbYCIW+mS9gMUalsUO2cfZs0WBvfpPPIePedb+wyCVK9SzYXHSmxbt2qzF609yJ
R42q1cxtyl4Osv49kb3+AVV2GJAvffJLFfOZOyUKW3xqGlJgBKGIWbOw+LYI444+E3/ilUMppatX
21VitL2a9WO+JuNu4fHhDMh3kFJby2Qo4axuzEpgmu3mBaebN5XFlpex9mk/sVAi2vgX9lJZzcz+
nLHzk0bBOmkKS5r6zpviJ5UiCBQItztNo8EINYc9SHsiDnOjMksqdvRfWirWo1bOvXWtKjRzEJIm
6WrbX9hh8ESuhnihyzUd6iRQu//mq2UBQ4zRT+vmLGKCI4bbJgOnx4Dee3m+dOTGsUqwrHBn8Lqo
9RDoAmAcgeMK6N0LZbXsS7jUCFOQBIlAyj6Sb2CKIQtmx95dxaGqeDFuW4izWtKBhFKhKF8hwoNA
Tv4FVv5prZLJmkjQNByL6LHaE/5cerR+GiMXWq348U6rcLPumS2APp5+utQcO8TlPYmsDii1A9sA
OtNYQnGSI2bGzu+S2NVrBPcFvllzoiNggFpO6HZsKK9RcLCMM2iaKLqMJDtUAHGYNN5VPZANOQX+
fBp4ie9CLdQxeVhb+3d8UU67I4JnOzsYbEXt5usQubyWVgaoo7ON/nP/8V3ETxqzEP2DwTdqFxfk
S/JiqmzHwx6QzSjHqoS08pejcNt+ScVEjz9R4x36jgu3GYyluksHd27+pXCYASMlkRM3CJK/x2J4
VguUEt0bOG8F5yKhmGyvvoZEafrecEf5RSN47T1dWy3XNiGmdIbtUrI2oZNZ61dhzUPN415Z6Qaf
RWBejp15HABlKAmqd8CYp2ykvroR4t88lQu6ITrZ9pteHM3BdQ5/I7YbX4PVBk5O/jE7jnJbgcMg
KF0yzKdxLD2qjkd9LBTu51gEHtlGkGPzylYuU9Z21KqH8X72yqta+C9SYnIOl3An3k1ILvgex9xT
aV+v+hR2owciV5V82HTL6UN1ccNB83neNO2sgfmCswh8DRTH2eWLiWm0ANa2lm1ZhZTu4G9wTgew
ivgQIey7unhWChnkcfztARVHbKrC401bhaK4fmJMSPjL8LpZG/p2ZHSCSyLiS4aaYdCsAOGrMrIv
cDsFSGlKdaXm6cPN7eU/9I5bRslUU7BWDpnDYEyGFWdxT3lejdfPBTAdnS3GP+ymblXpae6vBJhz
QEMuyGDWFxAdyv7rkCCaiJXzs46zSZNavozCI5K9sta76Z5Ijw8TLmtUNvXhRq4MX3dNCq34sSTV
wyoKLF/xrvFEtn/J+6OOGL9hb8Xutr2+6ehnz5rukCKJlotxQ25K28+YvXX+DA2knI5s7so+RG6c
Lf8uRjLw3dNorU6OR8D+AuPQa3cjsfg6Ty//k/X6ToAM2HFHdWfVkwTefBU1LXpxMFqh0Y9oR27S
1YX6ySNkPQ7b9ltEaA5CdjNHynYdWrnhAJHKJi7bcopZ0RisVnDvDL2SOlkldtKXoAVxekEWBm5G
dT5m9M4wHyc1mqRpUxJ9vnhxMXGd+jzKfuDFEU2kG4gfHk/I4NKffIT4C3OUdWxQiEQaBa8TDAdW
shTeL5tk0gasWHcTO6qahvlgzvsGs8+zLkTxb/nwD0FhqfbO7LoFzrkQJB/hYaKemg9jwjSPQVhQ
A1lXZLKqX/OUcU3PxvzIJrzVKyaGqrfSnHLCZk7OXhc2ZfHQPWtbiBgzHvksu36/pHpjbZnSa0Uq
Zu2D/cGgRkrX9BYMQ3oY3r/uDPfrT002FPQfGFvXJhxSazDl+pn5OFuHFE18ibCh4XnDIIeOL7Gc
bsEaBTqGa/g/XBOvyFP58LGormtbCbzHAQHCbNft2EJ/Lk+NiAw/l9crolpZqfmXBy2EFUvKCMDY
AaRxX8TOEJ502Who8R7A/bA7QSUidzKvzXCtf80fWFr5pKahvTqVScwLx9cJxRJQdr4jnNeYMiyX
nDjCpIVHc4b5aFBdCRDPgEuAtQKLJa3MzWcJ+PMZGiZNNjVlinfT+IZwsyScycrh2wTMDjn2hJtC
KfViVe9aefooBJc3gWJR3CZum+kcaXx3vxFvazQd3kjsxYOXoxp/QkLLXZEXrsCQrq42kfbgiSa/
2q6ocYYSUZzlBNVhRxKTb7VROl/IG+afzlrvWyLUZPzZg0YvPSSrEgeA/blWCWWpiPTQs5Cp/fd7
B9e8iqxetpxun3bVZeH2v1JdOIJjHXm7ZwG5ZbqGHnQt9559q5B/o1f/yAJOu9oYeFqN1xAWIkSY
BFk+CIjMyK2Mht5DdBIJbkM7Fvwq+9oW/ly9U3HtXIOZga0l7Vc+mzqR1Ag2iaMHZTmKeb6SlgJU
4pUj73nm06bU/7vG51C8cyvKTq+DAApIFZaZZMws4D9w65/3Uq2pzguxNz0cmzlaqB5WtsciEEli
3msqyL0iTyM0814jg/v3DCHUNWgEfXFJiNi/WQtxD6C8CMBiS8Lt0IdCpoRQZbyje/8dX9RYdXzD
WexdDd5NnTrnjEvEUrtOKvNXQKXpdXGjHXqNcpUXCJxs2KNbcYopuK4HhRDlXcOzmfPnsr0FLp5C
zFFofrWb/4WXJ5voMp16Ox4yjj2pubAlFQxrxQfESDfJ6VT0Ro7QT1R88wzIl9aH1CDn2cF/khUE
BcX5Tw8u8+W42FC/0fRcYQdwhMJWN8KA3JpMUJjHnRx3CilmvlJft28LJxxZaN7Sir9vYUUgYakb
oYTk8Js1cpBCZ0IoGPE+WydxzuM1qF4LCDe0KNCarDDkhhlOMOLmr+MdySdOHzWJ1GyeuFww8RR8
wT0AwOgkcLL6o4+MZC+CL/cTi87QWq5Qg22G5D6Ok6MBGkgBc6LQLYbrUD74AgYxsHT98nuJ99JY
WNQjascRNSCmTtboqDZfVA1TnsSvpkAZvI/kI+d+s9Isee/BO6Pbih+tMHd0WKzs46POoca+rGBb
ud5uP7UG7SXqwAymGa5EwxX7vpOhZSa30wq3C0VVPlgjUPf/jBUcwp4PUhUTSckW8JB+8yd0z4x+
3FlfDRMEZzkNiQV7FiyvXdRVu35BoEO0QPdOmqENaLZCwgyKXQ4IzNuO29SqB+qelnYiZJMH2uTu
uPAnsdQ4/NEsEPfPuUscirfYDXkjb1Vn+3HYFSVoZLXLXpDHWJnTwMwFF31/uRb0H6ugce7Ld06i
34mHkF2+y9Nopv682bd0r1uo7WGsnUAjSbn78nt3I69HnHIi8L2xCxDDizbHEQ03/YA/xsaGKRVL
3/8TNRoQrxgTvrV/c7SRI8Vs++tmmuWxt2n5nKQT4hXRKLkaoU1A92ahzM9WkvOLfgQ8HlkpAkcN
Gdv6zuJ3LyBn4MBj3TsTHWZb3WN3JBnhd3L++WdfLe2fB5RHfhDdcRQoZRiyMHMvmFeXoOE/f93S
FdO2KKd7rr6W9qrDi+YXy85Pp3By9jWEXdVv+2vuer6Ne+z3mwoNIcvegQ5Vl9opFRYi5mN6WZ3c
DdT7gD47cx1/0Bib2Nn4vN7ibTt0UbYBf2XphTVp3J4EhlootaJcOzsRhLofNyPk4Njm1KRapme2
jiYjRBohb/LesmaT3HPK14HKXRLOGd09adkerXlticUcA/7RM9OzL6g+F1yrz0/80T0IAehT19sv
wzop6TeSrnKBRh5aGQ0bi+mUR762jbXjN+aafFddiMTWss7OrqiTli6+364uhCzAzrYogmTVtdWb
W9xGJRJ1WSU2Pf2vMs0K+UB+z0btChYPcGtH9WeHlI2Qy9GOi2Hn+Hf/yX8ZrU/Yv2fAsRpLrtn9
0y0fLTVDKG6tK89kTZrwOH3E0Rb4PONYS3Nqlh4ShPWhibENXT2aCX5zPfAt7NZzrnOruk+qfFQk
2T4Dj/9XY2atTj/24bBVYuwDl7SI+bqwiHz8jiXWl3HCCgbWWpUwC75/ScqPDPWQTb38VQklDWjB
fXUSDOH5WogByuBPbt0lWrek7VtJjbBRdDBYY2Ex6X0P7yLCplFDsV6Xv7yhHBdI7rrqVRwoxGT8
uLeIeo3CCac5r+S5+qZ0D+yyjAOCYLMEmMGI8sKuyGESelWIHO7PSAJAm8fdyM7Y0Ml7XmJIIPmH
LnSBzQZ+1EfJ1rHx4tBChxGBWRZqfHK3DnofxrO3YJTC7vR19KnxvhQClYgqaImlKRBvS6hSFncq
HLuokEbaGhyLRb8MdmAT1XfbeNj5Oavl+9sYbUn2nyqY4Nd9FhlIPaZ02699Xem6r8pFY9OZCnRq
hnHD7rZ/HvEaqZfXJf8Ob41F9+mTSii2VW9V7H0LXcgDkHNi32U1Y5xPGuo0fN7I97jK/iC0TSdN
VSJbFF+Wc8u9nC3n9kq8SCZfWmrYVygvQ25eMZvc1Zc+fFN63a58b9jO8MbR27X0oY2U/4nAVezc
h+sD94+li3TfeHxsR/HyGHlhricf4ENF/ZBycq22ttuiimnwvWtBFEWVnWuptj0c3G97i3x0lpAh
HYNAEz2N4JTl0Fa41n7N6XycLRU7zj2AzReBqmejQFbFo2WxSUb45flOFq8ymP7epQL6Tnl9+h9Q
2shLcyqidZyE73ouvRcHnuQNtcqLIfMEzx8ypaAg2J3pHiSbRzh2xgwoE/h2ax8UHjzvM3EHP/MK
/mIPSTwUmBhULWFVij/ucMQYwQh5zhHPFfooY9xoEFd4dTUoESNf6XOpdbfZNeGgTZs8VO87MnbS
IHgdGHS9pTNvybsThS8PkNurZiTcqs42nK4t85V9kLI6OkEwkf0SB69Z21RAgtAnbMlEHkwH8S3Z
s/e9kzhSfw9CgCl7v3fPtB8IJDllQIGENdCW/9dc6P+9y4u11wZmKs2zlsAjRHtOxl1qVzpfxubo
/0+I/bT7IprGhyY7UUVEhRc7865dm9sDrkwt+AyLuOIez7KJQpasPI0L1CibJMtS/HMX61k6/e0o
zc7Zt4MoO4h0ZJpF/gii3Jhp3PA2E9oqqBEL9z81Uf2b23ddXBusn38N4XDX7PK36SM1TuOp4hgg
ztOJzjZflXNomryFi/kvzGYB2OxkZK0wvd1TOwj2BUZOlTptcl7V35qsr3RnqsvUEH4VkDPnQIge
/pimedNVtc7Q72uwu/CLnko7ne5wI25cqjmMxRPy3DwubC/SPtEznMwT/j9QabgV3Cr5sWgkBA0j
xU58CtAryWszk7dENIdy+qYv87yK6H2xs+RauGo1D7FTUPv2Cbyz0k+a2Ym6pXuFo516wzbq0MmB
GMFEY/s8bwV9tx9RA1Ngtcllw3zLyhpA0HdkKNABNmfShF1dRdhG+3jPbFrnjJRW/uM7n2QHBkhn
5pVwu+8tteP/ZAOQT1+aSpiGz5hMfftcElw1U38g7oBtO+58JnEVNQw7zqCJX8wo58mEJiVd+7j9
7l1v4WV0PMBX+acg/J5t5ZBdhRDu37+W9D0nijngmihpQXPsq0C6FyyWyU3/GaUNNyK85tZKizbe
teydNrS2o1rHZKfk8p4d4xoQsk7wCkyhhKuDqGsDGhs4mHZMQawt2sYhxdNLvMvvjqfViI8zDqu2
mJZxqLQF1ngUVZqyBoXDmEG7WVrvna6TzXVb4gkklqfLeCvxRqTTApmkh6HC+FtUNdy5iiOHKDJR
yGW0pYceptj2HsSNbJIRRSPpyMI70eOw4FcmiA9ZumE4HrgJxon+/P0JVzFYSswQeAYCzEfYxMIp
h6fPDmm6tLi+DEokC8OuznX6sXYZYF6Z3upkaqnUg8FYobHZHT+e42+xGM4mEYCjkwl8Cjw/kMC/
hEdzbm0Majw056xynbxfiLgEdGBz/4D4Mg7pjhQLgphO6hXn4fZ87jp+xDiYr53PSJbMjQ2S53La
3BoMPzCzAbFUfsp7nsR/vpWYl17zNiU52LNoHlm+Hl5Hr6jm8arpURJZ7ErqIuryLnXT544kEXMr
gULZgvnYYNuum8SrP06j9ipbkK+sPTb4bvdqexIW3Op0YEDaovkNQi/Ad+M1Cxz69fcybd8fMRBA
MhYzJaMXCDPOq2ZrPhG+q8B9oPGOW2KmTZVcup+Z8Vl+no9utWu/SN4IzHd3sVDiTSFiFL3OAeFI
u4+1cLOXUnsw7KlsRqG7+PbSly4zuVvS8PCUwzCUz1IEH/Gtts6Umla00vdQnZI8AKRRZzc+nOv6
gDIN4/I1uR91WMnrV5WOlu2Ad1zhCuvM6FKCwGpjcW9W7C3H3v6AZSh18OTqAnyx2DDvxwaS5A7I
M55nkifR18m23TtVzOr9JnSsBft+m6WL3HrLQhf+LpUM3lArG+e9KFupIOAlfwq8V83ok2CqBwRG
Z7Nc6FelfsOHsREPyZj5XK/WDQtMrpFPJ1cA6zGFJXHOwaeJIzN7pPJxXQousEp223IHvKEqrkXC
QgGbcnGkuzpW4VJf/Kpxh1dFaWEKbB/PI/ghO7usJsL/2G/nfWejF6rSHzPJ17i/swqZv/VjDCxf
BgRn4UzlT/t849gllXrOKY4wvv8nhpINKCqAjtzr0YQG3uunaycsZ36FzmmeqMy/ZcA1xVzvykYU
hryf1/+cHGzBrXw3T8lmj9if75aVwKbZCUxS+h+r7dADjwruAW3r5c9zMPLDMfPVwwOowxtM4To+
FJ6hSm53BZTZBgxASuI6itc84hJFBRPsPnwlTyoZmm+bLEivYrpeoxrQrk6Vj9JitF6yhqEofB3I
M8xBn1zffY1Xsq9f+uB7e7YAeg0OnkgbPPlmLJyaWfceAZlee/G8yBrbxTCMpgIgAfWyjZuw8QHx
5sXcWmu2EEXEAT3FfP5oppuJCwFaQ13yGII7J9nSpkK2qwKpXtZnLbHklPXAXYQ6ldjcdEnWLyTX
Y5l3bTnz/LTahCtSiiWdhZgJukKwcEWi0zB2D0fwovq7lgLxZ4TrQWorsIppxNPkXOQwBSQTO6EG
ckVIKJ8OPLJbWLmxtHkmeYQ3PUZlMCPwA/c0Wta9d1icRugyaXb5ItDgt00Y+i8wyO06bkes+H+T
xCKMwfcHopMfduLPUimSvlvySuxxpfRIJH7G4MeN0QAuMFFOERzjDhsE3n/w7aCp/EySO6ZjAAMv
3AkxLNInEvVcI7Uti7wWOJOwEtHAtDLtxUD01fovPKn0QmX4l/i70ZdcjXtxNqDY4ZNH+xJtaZab
8Q39BkxnfG/ETcaQvITNnFzOj8hyq74GGPGyty4hnba4Fuu8QU55y+76IJEUa1BTTdnVGnxTyhml
SY8Xg7hp8sWFxNUJnc/JxgaopY2UH4aevJwHaHquxyQ5JJu6HEzUdeQWlukfKHby4NlGY3AnKa7x
db6ptyr1x7fxTxSupjwcxQ96DX1fTWjr5Vigau+vW8iYsVImP2k9vTdrD6hhQ99wHnSZshq0xAUE
tq/Ls/oSnZ8OEndGkMLRF4JDxqfYoohEEBXeQTXI4pqumYZfP+SjSbW3cnj1IETiWY4MSMxArVVo
S7hKshm8uHVDpTTwPJXPIh+hE7dqsVE2OfeLdjAD+ogtpiuW5aik11/hQBhBTDxrsz69qzMnswKN
eJueIS9B1oxCi7mE9LMb+gJ3/aew8y5OjTEkEs1z7DAZoT1ajLDF7/IBRQWUy1ey1Hr2qYgY/oKe
RbLJEd7i/xHbSYulo1fLL4Hh95b5Hx7cPH9eT6gMTqvrM1UTn8cAhgZvWy+B6GuLcGna4RgfPcMW
6v2GOTD9nho1mMwxn53FFoYfSJ/nIwHG1+arBE3YDcL/sBHvdKh2Y8gFA3c+4KziAZO2eJskvXus
fpMjtO82R7BY47STrYAh1Euz4qS5R8Jg8DUer5xthJKcv/O2ra81OYsSYN61ddIWUSJak7eilYs3
O1xdoDPCJfz5xyiKWhL877vPzBc8cUgHQVrXndI2r2vW0VaWpV+5glOyyU8WdH9xEKbZ16WjgIZJ
Lv9RHfnldc9lub7tEqjUp8tuS77bMVoYI/G9WE0R+3GNcHCbc51yCSnwiJhHZpHCS5xXZv6JB7OL
GCLfv6esGRMHJg1lvfHgd5CTN6r9d4jQYTnAt7McN9FzUPLGN3pwk8Z8a519VgQhvI6jxwLREo8w
HkE9qLpuBT6nkpe5EEQMGLaqBMxQ4KArQQ2HVlqcSzQwOTA/Jv7smUPiNZrvw2ZRxlEKqzBrY1V8
HUON5EofXYJV6tWx+BVpldkwiT0cvz09lZzNH5f23GBQ6tbIIikEZHkZ8v28P7iVLEZ5+88qS1fI
p7Zn3Uzb5xqfYBF10MLVHS6M0sc99nkrQBl8fM1FnyQYU88y64/SzmRB8nSwqBL8TheDZI/e0oTi
nGVIoR3n+XZZ0/mIxLl0ZxjXkGc9nfav8l9+SVMhMJA24dooWHI8Ht2MBi+N26fM1ZDCkMhSdFE9
iFINX4bqUJjCimcDscOLIrCfnpdnG27UAthjICt4qdP7ueLsoMyMQEYV9XbnrehKTntgb30PFzrV
Ka+poASQANzfeiEKJEiGrPu0g1edo6nHaM7xmuBWkOB7dWgYYQIGSZpxLXHZBAZuahqLFcmNIYXK
CYPDvS45ZT5oIkLulJcmkBGBtCeAPV9RE9nuJQET8MyKKp1Zv8BPiqNa+BJ4Cup7tTvDZvTbLnsR
muRR3kRVnYgo6txcR0/fHZNm4Z50BhM82hRDhLpqVLcsDS5LCyi9fKDjQ7ciQQbxhh5ErjXBauL8
zKkD13fRdR0B+AzsQaKj70HGcWubjffrfRRDk+pH8Q81lW6JNP2h4FpcB7pNqUcKR7q4UnPxUBeI
WO+TccfHjIyGc1WKkEKphene817X5GgIHGcHfhnOCT8Glzdw/sHnvS/YDHsY+2aGYBibQtiGa62t
JQLsd5vVdURnqpO8woPqr4s7SnKgsGQSrtw/vpFDDE5WuLSRP32JNDWyt4c0jlNQ2fiZztbwmQLm
Jvq0Ml1l88m9Z5gtAWKQKKHKJBW0h2lT9/2uabUV5oD4u9+k7FrAXh3VK9WTdjH9b2IuxiAjTxgc
NfxltNWRbNs1bEz3QZvLcJoUfRvnZzleyBVYG5eT4gL+j+yeA2HT88U7JB94zVeE5ZekLP6m/ttf
VrAxD+RkDF27KyePwhrneNlYAPt7E5DvHwXrzhm0R3fP20AGPm2tDP2T+Z/lJxx1d5BQ3chqlDYA
Prq5MLV7WGXK9OSU6C16+NE1jhv9SJyeoM28RrUoEiVaPP2cpW8ce8th2QllNSAN2S8s0nM4WEWQ
UFj7VhCU3Nc8zhU+cAO9Q03jgxSSl84epo7h9gmj0y4P6md8QY2fs2TBGMN9LRaGGghVHMgYBpfy
Fqb6kmFxvOgL2LIvGwDcrVmvlOiXOYdBCO8bdeZSdKmb9E0PtZlvg97WlEiAuV024LJe8BT/OaER
QXm3dg8LBsIjW3CAcOKW/cZMLRq5Cu58xwlQvFo7pxtZkxoanmIPrOimUhCQr+WLOXtRPb5ct1GV
l58YNJEahJELhUuDN2EpSpS0NsFiJjVIFk6EIMmRuOl2ZQr8R8dDF9qCRdIsNeDHt16m2qYJUia9
ZteL/xr4sTVihjOzYjhOL0vAqUAc6y12/r5d3/Le0W5Z7miKgfy8zwJuxgowEFwH5KpEa63k5fKh
cGCQG1O1lNAMgwSdlE2JCfkn4SsKlFBmatTz2JbkwQMbx9m/CA/juHR6IQl+KJ/+bJi4nwhQGERl
gCOKb3hSRy5WAb+ninO7TK5copIqGccAu6fgTPaceF4J4SteesSEy87jDrWyK76Cd4pF/gOA3Z7u
LkvT3IvxDcDOv5eLv+8E2OPhvJrCY18ovo0x1vVYC/t3QF8lYQ9CAmw3fbOnEByHiOBbOd3kA9NL
lY2I7ntvsK6jewXczejdETzylmrdJR2fuoxo8k2ezbZp/URSTIiFjiM22eDfmRw3m1ZlOLB2upI7
MskoqQUGBtSzxL7Dn5J+RSRQciwVhzmBAh4e/G6Dvw5c5h857hRhDG1rI+tecOpaY2lNnRxM5+rH
zZV2PaFt/nzrsvdRG4QJ66g7+QCO5sK0vEsW+mCxVCugXKChjogRgNkDv44jhK51ujV1LekYVLDV
vOJSDE/fU0CFuQcrRvGziTQmVgdb/OhINHyH2snOX2tlW6gfmkD9PgoRuWy8mkF/LygqC7fC6aaV
eaO0cGD0bGG/UTSGUVLSN+mkhrtqpP9LBbG5xNFAU2l9UeAc5zpzwrflZ068mUJPdNwvfXczv92T
cCdInM281YCVoC7JNgPWp2cpgTZAAK5vQEI6aJ6LtQ3ApQWTZ4c0nEMQj7zhcxuabScPoq98uMaj
nXDvBMU7MQY2vItgteK0h9WR8D101uC5uH6jmHJO5vlov0JPNYQ/uACShOEjG+bwAR+EPbJhGwLG
E2k9o+328bKJ+BWw46Vz5hAr9FTHz8lDR6xB2y8ONKrS/6aSn55cHUYv6deKUQe4fJ3pym57KXvV
9wL1kCcSu8MezQfh+xs+WUEYAlzZRn9X+ZXGxJkh3NhQtVVIqrb5sn0Nx8aiLxUnXUgTJSDTH7d0
nzfieYYabtJEz+fhFQ3S44YIbBfDWWRHUX+vpCewETfRFg5Js6L/jpNikSC4WgmqvoREv+axPpoV
WGPres86hhmIxboZNODm4ZRi4g==
`pragma protect end_protected
