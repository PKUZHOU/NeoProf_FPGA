// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
JdE1mFDmMI2cu65Kvb5W7SQaif7wFLzd9eDLN+EdSd/8HYyKx3ErEA55F2ruFHEz4m2KC+9n5CL9
YtZ6iYVRWCwDvthzy3dTvq56/8nLSsin/NyNFw3ojrYZlMvc1T+yCfMWnQ7fWkn0+QnN5udSGmyv
kACZYW97T6uncDkNzLsy1PO4Gq8oB8VWlngZjsuq5JqzW1W1B/I3Vjm56urpnq5xettA3ManLhjq
XmcqsCwm0Rd1Al/SuupOLLyP5XSKbJyYl0rNX9Qqnv3Ufx1vZ+DPyvGla64Bhvc6po4+xfBVJbo6
cd/uk85VOzFOczRlMrk69m+vI7wX3YJ16ODSIQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 9616)
04usM5xdqhC/pnysPnvAbDukXuLc7WTZMH/UKZxhvqO4t9aXuEK52G0ZnzfSXwKjBG6xeQySAhqx
bLlGgrp0QDvDDDB2R/Luj96s9hagyNuhHQ1o9cF/RQ5w3rclKsArHV7ZRW/BQnQ9gzVRRyhsx/yS
qKOqxdRNGndyaAXo0SQdDFovigMZVFEm1seqjy9+bk4q4K/njJZZl3Z/jIYyNxAfqIba8waStvYk
srrVFCy84/ByInbP3dSIdatON7ncxo88zNbS2LqlhW4rOIV+2JUt03PeJ0hceJS05RHlyPEbtzND
99XP3NBXyw1Cna5/v0hxl0E6YDYtKVUWrBDQll3jzWIRBES4xtD50FKPZziaH22CRiT9SPeMWiY0
YMmx+Z9oVq+H+Nn1BwfRMfn7QJhDBZ9Woa/Nd4wD1OnT7Txrt2PR7exFLPrt1ODTgDMudp2mj/Oi
+BGO2Qau3hfYmO9GxXXUxLILX+FDTrbU9ckBrn63l4KWcztc3Aek2jZhMRCoFhBT+riv9BexxmZU
MA+N/lEXGKArUwfqT98qoc8gGLLZQLWOAri7PaGuC1bXfPf6apT9ONF9KwOJNjGDKKvScb1mZwi0
JmQwOZ+wgvwVqaqQkMtNP7LKd5dJIcgB4QXBRJlmz+XSb0qlKvoESFC9QL+vBvu6t5feJPJ93cdk
OYkAG5RW+TV/LoZEvmnEf+rwWMZqtICphWi4lUCZEfEuRTMy41dvBGYmLR4UAXocqDvj3ojX8zza
5ZDhOVFy0RhWXvShRaQOiKHcGEAK5Rkr04ipqail0+4Egf1xjjCsxWdB4SWGBYpvDPDnBTC/EgpC
uYVzpH+RGSOdnzrR2v5HelOK1IE0N/i+JQFA9RiZ3Yl6SbnJsZrlEhDVGSfLaO65Hu6YZWGBdK4E
0MpZVY1jy3xeFpxFGjIxbSCyOyqd6+zfoq5xyRRqnjaDqOUHuCkD7dAIsO0j7aQYFOIFNoODrCfb
3T5/F5w1oJ6wc1DT1psxWGC8KtTkmnYCPy7ONS6sS+bwqRNrapshOG0RaIeWyDehloETHtS4wcZx
p6fayX+ovalbuAqOpIMIESr756Vic8cf7xj8VeIS8179dlrPjDJB85THEiqC5weVURo53iUwKvl3
+dxTY21wkSSc9HEtB2MHroWdJbS6q7FPczVjt4uKT8vrrtmJE43mhS8MNwNlW6GvN6cF6IyDrjgY
e/K5e0SwKPqBKUsCtfX6qB09jWooO4NXiYvB61lmyFZy/R1CDYIfnu/c7fIveia7YDTc3byTVbU6
egPe8NwL272UnTLcrYQYfYp5fnEsPyHseY3cLAdziHWSKE4PVRZFqMOvU1YKsySiRiBANMcLnTLK
GeyV2s9gFui/uUIA+MiSzIj3JFe44RdbmY61BhEXBQH/HDQcIsiYQgiQHoKZv1irEEi1ZcKlJT8T
JciIXhI0wKxBBQMOhb9yjEQtQ9MOsWBLZx0Ze8EscyX+iK82a5iCMbpb4kEocfc3p4BMvmMRiEaP
W6Heh2RReHG6tnQsbT8+5ussz76MlAC/nMgqJM2fCMSZq1u4RxnDbjWD2ZStfFKuSkI3chy09sGc
PWhOgoL3GizKre9iEI/7Nryf19DNst1prP9DGoJEKKqvfRjw+Sun+iYxXjN2ivYP2eyG2Bpd2Oc9
5p9XEAS2QNqCDWGYY786Apveev7aldRzhMS6VtaeYSf2vGKV5TIGAy0eJqkwd6GB7fPQyMkTHQB4
3DTlvHiVM0GUU9AgOu1+ZVKdhoa3JzChs43/OAmN37LdPPMGzTkj/Lmdtpiw95w/EytS1MI80tfZ
GO1htZmuSC7ULVYZW/RsYXcECpiv2pqvKYDKd8PzkSNuh9WPKwlVcrqg4ogUuh7vBeOLOsuCNhrA
D8RXdKU7wJrl6PDLk8ifVBRKuNqS3F+yH0FfZU+m9CNQZ0IciYZ2E5Pj6Zbzeu83thsusKCxKCm4
POMKdrz1wMbOrzhAE9y3EqeZsUkeL0azJRznsuYX2zSGyyLpLTvzHq50KkCmAmgklwnCygRj3DsJ
ZIPgDL0uw3RrI+hiLBJ9lbJbJ0idzryyTj6YF71oY1YwsTw1P/ujuAkYJZfBZSgEVlPHUhIbM5dJ
hQhu/Ger06WDFBFz2tPy/4FTzeYAhr7wBOn/3gUQM8b9uISc8jQfWMMUQw9ezk++bUQG+esDzFU+
WkGzUl0k39rIeyjqVvgWLh195Rc4X5j7S0J5AG3ivXzqDktIA3mP41gEiVso2dtEb78Ft34Wy4s7
UUjyTxA057ZHPTj+h4hG/bEAyLgOR4Y+GUAQ63eOMMTvJd5bvw2FPbxHey9wEE5O81yWLnrXQm7j
IdxJKgdxplBHD+TFLjybA3iflIkIEnu1l6dkfGsS6YOiF9Wm+tOPPFmS4wACjtmtbMdvjskDDyGR
iJDAeNh6Dxv6JhIO69O3LqczpgzARN7vCFHO/wNFSkxuizMx8m7BKGiqMiIlwwFJ65W2UI6KdUyI
YveOfY27/Nq4m1w5pcv/a1eAeRNSwmfiA6qWOIiswCnpUIZNGrS3dFl/z31N0lsCxkbI9tR68xG7
i8O3vfn3gyDRchZNkFvMBDTpFaV4LP9zMdf0uXWcNScBdzxCZX1I9Fu8BRA5Y0weJ08cGxl3LDzi
W7vpWhjq9zE1zECneZYt+xG8+NFECfDmLtkSSbJuwDqsnNIFr3IE2M+fxtNXcBFDI9dHRNJ8e3fq
AS+QmGOLFBHZ0a0jgbileE1f5HrvFO/1L7R4dPH/rlARwz2UBb0Qxo0TsmKDUEzat0mcaJjpUoit
2JbKgfHqtQRenP7RNHTycByXX5jTUDqwgcjwtRIPDLLevR6vsNaZcqxCK1fbxbsSlzYi17at8Ufp
tr1Rua/r2QL264i9+ZZn2rq+gpKmsn8buaEN8P35nSmVDA/atwZjzAIGku7qhw3SrW1WJKsp7viP
dQwFTsnRylaWWeK1Kkk2R767GYx1kYXucKF2/f+2qQ19utmKmh4l/Vjy1eg4DA9CD9PlEkoyEZV1
cubiYndLAQUlT4neew7LBDle/M6O32h+W4ku0AKOsk2NyNHq9SR8hm63KAPteSYBFfI9AGnslu5E
biwVByj+z6s9J+lqJxaKKTm8zy8BEznraViPXJNpor/V6cyQgmNe8pBLw9IHB7pkxPrpoH0cIMWg
iJCGUa5KEwcYHapX1Fy5iT9mTOy4pM7gLBZk8nKzezXZ4iyZJca+HFED6lhoF/CCAWPbGdm1qSfc
rRhyYH9hfDNWryXWGkYmaIou7lAZqnBhQqKbM8v9OWoP+CEf6ZeE1DnvNJcZu82c2ELI3G/iGOxu
9e3Qz75xZuuq0dwL0Vk7OAFl4nnzD0Mkv1OiJCe+i8lDa+qTnDX/Vuim4WPBnD+mAW+6tFBI4EZF
1MlIC9eaTgKsH+7IIsjgourrJ1ndo1r+2d/5UFlQDTgKFByCPtd/uOCVjHqne6m+7Rkc6jfqbBSH
JGQR8+7KnFzmd5hm2kbif/QmJT+XKHiDI+Ieh7WC38iWxMo2fwLYSZDW7kCo/7VHhgLWWBokHm2d
VKp5s43TklCjL1K24lzK/6xhpXoPcCh7E7R4dOgYG2X6/EgOW8rDvfWJfmX7FxOqO/vTtBmwfiop
Yup0DzWJs2LJXhR0x+ztxw596LJZrKmPamzNV8t99lEp8jBSnBRTO8Ej+paAhDuRt5RIQ6eZaEie
YlRfodNyBpaSDN9qSsEEm+NurlW7QAqyYjIeQ6bUfptJNOYUSCFhmGQYg/6wH29l9lONn3KbOAlU
lusRhtqts0RfGkbbo0hj66Qsispr2KZcoKx+Ekxuo89TiKoVX4qmLUaTlX8lR07O18mvnNKE2K5f
Mj/GVXNUozoY0RsRxQfw6UjXsmTIST57L+B7RvOf74lFEJFGSG5eko0IPgwNnAzG4tRpWAuNAtN2
PI866OtRO00921HGoFMJawqN5cqmqSW3nRDLkEhQVAffTJ6g2jQH2dzGpoCrCt8i+Y8n6sb4na/K
5Otx0udZUdSWsusRlaINH2GP+0XJL4vC7b2LWqOA7f3tgEyMK8iDgu3VwGn+DtRmhrzaT7OnvBjy
qJF7rmg8G7EXD4uYW4OMwknIA15k5HL77az8XLVoaKhWQep29/C241J8UNJtKfPXfBH7MqgauIin
eR7CJ8NvOnEh6z8qI5q0PrAl/MUnQCAsqcomravz4XKkrS+KhmUmLp5OOJNRk/2KLxrvv2u7shjt
9v2h4kfjTAwlZTPgsZjevTgScxnJeDdlNE2E+FzNZ4zRVx9FHNWNboeujVdffrLI41vkV7F+4cqZ
FC36zOn689yRa6gw9ofCMnnCie0SCjaTtMuatIwKtSlfZS3qzfnqPfbe9bdeln4Skb/yanuSUtQq
zssvbx6KWxXdj37x68UqmYsn7VCczSK4779KkB4d8YWWxo8EKcAxP1p1flY2etvksA87aQ2Maqir
ZUagxyfdER21OISEq4YwoS9OWA6mmAe5MZymjdlEyTctQEEtunqYGB6IZ3oQ5x9bOEPvZJq3SqwS
EJlaFbZUcub2HVMmKTzmEyyC7ZH79uYd3aHQL5M3RXztnzfA7fZxa2A/Sc0P++iiQf3MKVpggb5g
NLByZxlNKNBnlXQvXUfuKfx8Zm5GS3YwIxLwXtWxFiD9sVBS9JiNoVgoKCPuVu885Wfs052WQSaU
r9DcoylYySulW8uby+VvmSb43BLonz9NvkWoSTqRMUQZwLd7wEEBnrthHu3LkLNwSF0B4LDqPIJP
F2jpvJjRMNn95n9BfdurrmB6FKo3Y/2AiTwoK9dndD94dLi2kXCJqsJ64jEPp+ITLXp2fQLfDeaj
J1Ge+ycVHlnzccdDjnDMmbk0WWmjGxuFVvgQ5DgvJ1rfh1dhyKeVXMrWJAstx406qdw75j37yg5z
pTH0ui3PGIMLyiqibQFQ1YeqYUxeecKm5oT82jJjT/1+dOdKC5vBflKSlQQKEatq6u+gQgfLprGV
ab3gR71Y634dNxkFw2dYBMKQJG4aHFzHWv16jI9u1noJaqQeM7yCs/RA9fpme+qQ+4QzHT9bcZ65
TAxPWMgTiSS6d3zs+XUXopfxLKfP2OTyDJUigaXi4m66n0NYpZuzy8kFRhIs/YzXPdfDa+TovHmE
t0CVCDYJ2Tsn2YV9wWV9+zhTzjaEGtqCDCLdbF15rphMAKhHnOnowi60tLdz/VlqOf1Ladwb83oz
ua8Kr65meQkE8JMQ9II1vchp0Z/dZIzg9waMk0lPOpMgFXpcldaAUtIdGwAqy9Xn7ug6J6BTA7Mc
0v+9LW0XrKTHZsv4yrTQE8NLoLRD0334wdllObra61SL5+OuVXe2h/tql/jSXa83d8iOGIS/X2dQ
O1hWFVKvyzMxo/RRbd5naRKMBm+WOmwHq5sedRtRPhezSaYnFZ9IAg/bUSnOfn1LaMj34MhEO7iH
LPdQ0vNbbGkruqrk1jUgCuG571RQuMWFeOIdX+Q0eU9C3EY7BU2mZAlFCE6JjlzfKzNV3iieWrNI
eSwDQUsSTTSYX/dxEhAxPTEc+uRgK9Kc7GVB/8hmM/eBwzrH1Bt+KWIw0z+Y3qSFqGXpjQNVFF/R
zKdejckR3sgjSpWv15k5M6NtKdBZWq3b0W3GbWPbrhNL2Bqks+eJ2zkDLh7d2AIPS/R0KGH9OZJ1
Xj5sU8fpxCubL0z6UHqqDIEJvHu5hfbSVCgXSHwqRYkgA7oFEwkgy/PaBR4fP26nqM3n1CCg38Ua
GAYhNJ4qNsOoKaq4ERlASydQOr7Mu7byTdtttXluHZk5Y44mLcDSCI9bQKkYY1cO9FOGYImh1azz
JajUxF12HdvMebU1FI3rLkvfNuEc0k4++wacpBdHdvQe2BLwMFkpge/S0EDiSDOOqya1bZOlydTA
M1yHWuQ3ePhggeA9zeWptTLMGBBUNVmwBCY8Sj/Zxm86Dy0+2u3uyShodg41W8N+adybn5N2GubT
z7PFbtr+ASrWbhmutFh+ecYGxy26P1IXDHlBTUCcRMPcEL4D6KPnXOx7JxkUROceHeQor6hTxu6t
qXMqaubcmFQv4lpRCmEcQX8Nj5u6Fvi2V7V30zTm7hopOEi4MiyAr3ewdoK4SYL2uDisiZHNLjgX
t+i8FlJC+ug4IWlHDMD9vbVd2XYa8j8mPduYHRCH9LWo7R8rHa3/A5yIZ1Hp/KEI52qrloFCvTzl
mDBZmYdViFzsLStYtnldJxPCpH/ZFfKguiOQuN9yiSk15lHpHbV53kbAoffqJMdEi10KM3tp+Q8w
d5TAXIfnvwsuvCTADiP+2s5FBz7ERaXMXdN6ZddmGkIq9rJR+2gtm4huRdOodR0bSoJyv3vtcZjX
yDzrUR3VxbYFBdMEkl+cItvwpBsGSzL9PDpJ2hRp/EFC6/BYMOQJ2lrijaY8UBGDYqHvFD0Xl3qJ
+oTqe1Raba++gnI+b2iupcB1pQgJHnZKNa0CFmC6Rv/FKt+x8uwLlwiEcMx0LZGneannLEV2sARb
XFna0ww73cQu+o8dmJMv/ER65NugugnmG/XOPtO1tovOYa05Yu5MN0JOtfSWqyGs3/FLd3NapTZy
GjOfDt6uMjqgOexLkc5yLex1FzvZAQrd7ETpewe3KCkZAVXdYHcQy8/5uI0yPIxNyWkj3+9tKcHv
PvldKJec78vqfzbG7h5/3xJCrStojxJbZu6TAcQDwHjvE3NniFpmUNOz8UQwKCwuBi7926YSK/ks
zfxYyePWSLDUk6lYgCYj5BirNTXBjNM8Sqr9uRBs5SXj450SPif5XF7RHsWc1fVmnEOg3qfoQgRx
szRBLqJ4KZiEmINuSt6HMaCsQwSMQb1I40tS2Zh53a2uTfds9nsKHnyrdIjgSedginww6oM8q1I+
CPyygnDXSYwiXJ7WD9yD0fBu4dImoBMedceouN9CpARaxHPoRgGeNTID6mDM6pQ+NiHlIr+Wj1vt
LnGXioLeDN9bhlvavvxh/3dotwq0BkR5U06+tiX4jwC50wktHKcKVutDURXuvbVGi3OL0LLTdOvn
H/qdhFyFs08GMujespvYdYmKPad2kQyzetOdrnr+v/wtEB5P8+cKi573H+l5XUlwMwiTQbHk0FDr
EzeUP9kO0tgc/de9mXbmPxiDkBtxfSqiYZ8koj6uZrog895LpSqwaMHK4I5eM0hjs0ZhTPPjqQiC
sUnIzyYh6JEkg8VwBdRmeyav4gLTync+8jSkLnx00eb7D5SQdiuIz+eKWmuAIbXnXByGa9x+80Eb
Has3WdC9NMUm6mv9LnEz1CNOnQ6mJ+IfX8U0iAVQme101FXDDrkBewNuKkS5LIanFxVprI1ndxre
lN5BMsgPh0hRBsZNZs5m2+jMfYM1+uo7UMEvEpfKUUGE6aECyNNYhq8KpsME2lZINPZ1UU0B3OoH
babX3CtKDycDyqXBmRI+NHN9jaVBJeD8K14s3uUPXO12pLdDeWuDh5nGwZ3UJnd4JwPdWDhoBCex
FHLlBxzFWTtm04y5pxVqvHltpsIey1HgPaPQM9i8TUp4MPiBF3T5vLmumfg8TER0+ppHIuDr2M5W
7QGKMrXXHHwY7moG4goOWcQRMxWqM8eDZG0bBbpM9offghHFOuR0Jt15GM0fhPTMEpIWQhXJTmp7
hMBoFmPFg9GdTCYONAnqxkpDkpB0l0U8vOhkMrPVPq1K2C66ymIpZH5iqFc2WirkBOpXGnDfcn85
b0J1t6HOy+6hw7z71b6+xiaTQIWjYWaiOsNlWXeueFqaVC8+eaiKZ08+X47PMq8grHAk5f3RQe7y
KIMCA6t14KGNG5JS1jAoQzLatG2xeSNMHD/gwTuHE63FROTU3sZU0pFHouh44GlMZPzEsTS4QLr5
8XgSMzCwaQV4OEtDWJ5AqxwGN/RpEmdQObIBfX3ID9OoLqXQTBPtweFKqT5mK/owQAiAYNOABsEe
lR7SZ/xI2iZdkqyUBq//7LxN7pKbQRqcFPzBU4MOWyrm96iMQzSlebutQM6wCSZw5RmAyhNMV/FE
rF1U8P6zwjFe7bre5oZ4Pc12rBXEaVuc9dozx24PGkwJKBAjg4rk6RR/N86/HBnoRsn4oICDqd7I
tdor+iIKzoomPz/yTk7+q3DyzJs4dP5lboMNKo1uNSeFSyHb6ZVRU8AsNh/xUWt5ricklVROBn5l
XqweV3qrUaVekA3ZvyYJ0xa7rng1xSEI4jCTKVuamJKPA0J/CEnmYUGL3f4A3nB8MUBEIEwF+nxE
CUhu3mutMJNroYFL8ILsAl9xvqn7rTIGd3XY/lgHVG75xYh6JPKJBjVARI8HLEHNoBbw6cb4VP8F
TqOn9JxVXFH0hkUpyHBC6q0pmqPNkwb7pPK3tTap6nrinXCaK7h3cn6NDDbaadzPZoXxra2wXJ9D
BsjQ1JEUfPNTwbWnR0BHFNC4eMVtJD1K3r1GJK/So9Dj8fIggAm0UOVHwdNdCrj8y+Cit4e9vVzQ
q/2O58J9bzaHpXXxx9Hs6OrEfsCpsdf1UUN8m0/JNccgWlKT8ipXGfJ7p2zRttbTZIuqQq3QnyR4
+rlUx1HlOH94voXsXCexTzq1qm8wvqZfYlZAormk11Mh3gxBKU1sC7WV+A8CyOufmghjBVAWzyXu
em4kET6QwBOio1z7cMkWUi5kndin3qDq+imFz0RRKMZalmSHuYd78RfrlriEf8J6cHdSIpVT2P/p
2MK8QLhjWAby3be74qbr3+FTdFwv78MQCTQzfCstnP6tEqhFiT1gHOl5vW/rv3/CI11TKfDaBER0
nu7K22Ve7yYFEA7TeBP5V2MraJPr0iPAU+r1DoZCw1nOa9I+HCVLz8YazbKNQkxizNAtvoAsBCrv
kxEk9Iuss/mVX5Td8EYJmU60Evns1xs+2Qpu583vBke3BZjy/XoUGV1PKJZS11EweAPM9arAx7e8
Ap6DvxM0gxtzMuRVgRjWUafjNlfYot6QmCJyIu0h5QFikYlepnEkgaJaZonFSGx7RrwBG4B8+P4a
4XjTP/8bJiAr6I/NiwU89UXlWyFOoNVGOTdNAolpFk85BLUS7JB4KADoaMra7b4JPULAgGUHxZr+
CsWpzWmSQNfUrlOsaXTvUN/km4iJ7md4qbk0jgLINNsX/v5zh20z5HrI3BKo9kjFqWbRIC1FnzZ7
k8021Xy3yqmuZJJp5EuyJD4oXcDVPLrUUC+C6vUlMQK+RP5+c2Y9wggPYjuPzx4pSeqg1KrC9m7u
MHgYfzjlFUAn0ecL+XgDe6+jXM5kcyjs5wfCDlwJQQ/UiEnlyfiw5df0AUmF+jOQZLR+7aNzNo/X
FOzNcB5QNxOz8lWZ0/okWqNxznYRppRk4RZTJJ0Cr0aPUWskMGOJBIIA3DbikZhiavJZMF0PFeBu
10c0Q2/Zv+wPsxZKEFkP3zXBrbdc/26JZZz+Zif1Calx2bzuF81F00yqdz4CbuhEc8QYGy3IJp06
oedQpbZhaDz7lkGqsA2ociLBFj7iawskt3VpOOvBfzCa++kCvnkblh2bq4Cwmm7P/yJZli83iHJD
irz55g00wxu8JIyFUY3gyIdNGkitA8RvyNg1lEoRxLJk6yXX4SxkJP8mEBHo9N+/l542U+M/tofT
AX0rWWIA5wy7a8xdqofZ65T7f536eOlXYofWSU6n7enhGNQxwkwuuJehjocw7foBOFj1UHu+3NGO
OwFOtNqGLBW4XDtd117hNzP5Y2P8SRrSmkULOenJhIFdvgdJF65XA0vd+KEpN0x6O8w5PG0vpGl7
W44+nQTE/Kz8LhNzPohugMxakpsFmW6THdeuFX8Z/LjW2FJArpjAIy9489/9XFPy2GLqQBlyMDRT
ftoYWWZGFP2pHiUQ+O9Ek3zpw5Ga8h7Vv4B2egnTCAep8fbYMCpGnBMmUXGuKgwSmixfVHSW2zXS
7MWQ3NbdgAkU+TPpzwEMe5PLKO9eY1jX4gdONKq7HNThvam1Tkehrf7LyLXk8E33a1Ir1NixTKUX
SWLNdbr+Wp4okJQpCXAR0lNvt6appf+njJuYKgAlS6pkV4q/4dSyuubTRImtm6cNqPXfQHWv+5em
/59sozZB4O7OTi6XwhRN3ZQZqa5935niWltnkGUG0NO7saK3uFwgZSsW6vwLp13BFEGR8waJmKTN
qgx8euSB99mkoxMdUTLLeb8Jr/Mu5PVUWRGfZkpSTdMztzGC6MWxHNHuKtD1hNdeuq8dEfiR83Va
dKrEKTgaSxngpTeJdsyGBNQabfQWHBElvgBASLjaWW3+MAxC8eq+Ye/6v3SHlovstoKVlBn910U5
YdhMN0Oy74spcX7h5u13obCMKAlqJkymjuAYyTWllvxFzdhmPwDUXyp3s5BjcnKG9NnXnx2J6YbQ
VbsHyJofD5Nz4UetDNpVy8BSsZwO+/oZpgsnbsZE/BdoOyqZOHRKo7MgK7ip5hD/K9lXHq+3CtLT
Tp6cJbRUOeMPbzKvpOoEsIPKG0R0Imr2sYIsRhnTJmGoOe4X9TK2qNWp0ZeknogU8Edt8UHA2jXS
vJM+IwLKjjx6XUUZA04IIXwJxLg+sRpxffT/1BJYVe5o27k2VtjcklRu3o1MXovx1ejy3niiQW4t
6IZkKeHTBPCLGq6qOtbt1ElWEPgZRkFoj9i8DOPLC4vCY2gS9Cz5dlGo3U6+WZIpzZmWHUOh+WH3
YZpIGdER2C61wNScgklYHpJ/RfhPOodiBwT3tH2gwE08n19YMcTXTwQI0cXR0oIW3QnhRIWsEy/9
m6spg6nnMIqytscXMayjFykGdgSkhxApANHdvVMwqf9pno1dQc+Y2fNaLlfhP9er/NjuyPugDDl7
QG+SMXzbObsqr4q1oxRzHQVk+r4cFVO94O0zzwnT/n5jKtZG942MHimonppi7q3PJh/ZOcyaCSx7
98BzWVEmam0m2mYNtNXgja6zmtfHTLoBzDarHnaPJyz+7t4XoXL3G05AT2kfqkspFyoYABOPHVTP
/RjZCrYL90OHPEPHA63KSsZ8HOMzJOjWjGzDYqScumbYT/n4NiVsBt2RhTUlsn3qKOv71SVoCUTF
667kzdbQacCJ+Re+/CIZ93X22G2aoHd7kPYAaB4psVxEMyA/nlqjm2J+2Vf2fCOlwOFK7+B59Cau
fh/iUgQf7RDy08RjGVVc7F9wgP2m9zedax94Eqs04ClY4tk2Z2s7OJkQJ2r9I7saRkZQjMAOrWBT
1n73WStlI+bX6USDzmkBfbJiFLwZiytMWNO98qw2oe6+YdMbVYpfKI6V7bRs5SX0pInbeswKyPcZ
ksAzDWWOPwEnzYE6Oir+SDsuqTJIOHuMUFCsshlucj1k5B7xRcrjOCb5xdZT9s/8IO/KmQZ35ZHo
jYpDeses+TDcvCpPAksDsisi7F9skaUfEGrprpHRTR4kbhk67r+423U5BO064iVOVHh3shH5DBcy
HebB1Q17sniiSds7yOUBXd1O18MOvdRJouopkb7tUjLdmCxOzprdvbTdoKCfvuJBumpMtrn4+M+X
3VSjj3VaZqAHdnylD/RDmQ4BMEN4xaWCdhQ1RmdNAk7us809cCH/diowN2zzsebnleFz3x8Xt13U
H3DJI/LrU2ZGLVGL80k5YB0OKUYbHWxRCnG3sSVfhuhC6rKFZ72DH/PAkEE30+dq4UrKAxPptO0p
ybPRzDmczlFf8KEzD7p+vfgAuJg9qJDJIM2Vv7ps73QQ9ivuLESPUi1rLTaO2L0eFNCtHvfcFBRl
cMy6BQmOWcOnyfW8hgWUYQAhxbcXJwTLlghtxZgGZ8XA42NdNoTmfKcd7vYplq92wEVuv/GjwJdS
RSoPtXZKsPnpxahBUmwFxAVKJT2E0CYSN60xRIgkoHK6FgatK8djQ38xfgjbMusinhjW/kMHrUw7
CsZiJ7PKl+B4CmYRnuisRejOFEqMG+bz/jnU44QPLGdStMDMOiPf5N9laOcl0GOzWERYcBVkESRP
O84E4DZ2p5g/ZWLAuc0ki95xgwH2wd2fdNn00Yj95nMTQwEM5EUYKSLEcVIaEqRo7e5nYXiBQojw
uPg9ch8wNaLdLOYYeked4KUSjwnDrMAkmTk12ADtXEVSUVEXCnoj0XKnEPdvjD0o9IMGI6QV5KdX
VQWMSAU4Xl+peOdWXoUbVHaVR0ktWIpc0zoj5veNeUWJ8SzB5suaf8Cys8equBLcGvnA40CrTFnA
8O9V5Onb2LqTzX92B3GsNtTAPZAYOYLx1VVT+LdefPRFQ8/pa4iw8Qncm0f5togtXzouExwBY8QR
rgp2MPzK6dq7dLlXzRMdIMd0t3s8VSb8m063qntaSWzx6FEg/2jvXpXn0I6aXHkcHXhX3on6/fJ2
Gsrx8Md3OcO8pa2cdA+vmO9EMhKeF4HqRP0hiB1Q3h5poS2d0ikYklZ28gMJZS7oLw5Jx8akG32I
KekIbCNKJsK9HYkxfsAVkrSeELoDHgGraOix5gThDh5+2apVaPmMgTCY2lt8VzgCPDHLobF2buMe
Fyjuj+0f9ac1IPpkV3/slBeB6cQpuu3j7x++lhF+wanjQDeidpS4Rlw3AWvzDZOJy/Rdmikue9qX
6oDB2lUXKs/8lECqzXirgZ/KOEW19Hjpm6vSF99QX9GloFRJoozc+9jC1Y0l6FZLiXIi+TMRgXMi
MRSX9M4MsNNTDdY5/12ByLD2uHLYKLpacqAfIKdlqTv2MKgwH4pWWvGemoD8XNtOiRzKMH3BhIOM
Eu5wBZMXpRh5OXWchVRCwnHoiWtP2XHqAUdm0BSq9aQFL4dWBXnJHw==
`pragma protect end_protected
