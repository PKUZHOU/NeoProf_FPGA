// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
DgNNcY9/lGi0Nz2ThD7ycqTH5jL0oPzLNyLDv8scku0nC86/5ZDyFjR7oR71zByT
2V9BuZ7sIUmaSElA5FMS0pQmjLzi/OqImPwcfhWpfhw4CKrh4SwxiKZ1x5dnY5Ot
KGL62ygCSgRyoT1EWejwRauV8klUyhEB2hWCsaJeUBQ=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 20000 )
`pragma protect data_block
fo/Zlc7WSklT34VHAlDu6vFMsjIjekyk1u0E1gdDmAE13TI8ivb+KaqJ7j2o6iVX
3yNX9WDPAPS4rBeU6dgGXPQQIZjmjnFmVYD8ky74Ky80RkOObNZtS438zVo89CyT
y/WX85q+RfKBo6nAwtuqsgQq7VSr0Lvoojej64vdYWEG3gcXRmmG/aQv6fuWRwLy
t57vVFT2AWMSO1OucatE5LIowDyCgWQwZUS+kq3CAefQFVE3sDdqL0Id5/AyhaYW
EZH1YNM3aUbNCreISjjhE6pkB/BfUBjlhXpMIz3CCRUAjsqCPfc0OxqNc2f1ZPsu
MdgEYYbdEGt5qj/maLb+YmoSaZGWkcoHSAHNUoJhQKcU8KMcxPGJC49qzjuWKEIp
SL6T4C+msEOzi6A3gmQPgHXcLeHqNUarnu9PUh1wqTem7HJbNg3SIepwAkvyR+jj
IOrzUN61Ndui1QFgzRpxObsQqjdj7OBKyC+Acrav3HwIwWnU+DsNDEryBUv905vl
09fUOnk92t5ujCCuHkIjyCPN6EQw2PEMO5r5kIWPaftOhUc9hRGqPdl1hY8dX0XY
NXjfR8mI7dg8i6Cr+w/NGwI7LYoVAaDENKuwsCFSkZyGRAmZhjNwF++eFCAsS2U0
V3l7De/J54jEaQXsTa1yxEbU3cSvWzWKws262rcax8GMpH9gBGcdSbcf3eOLk0tL
CVAlOcU9tWihujXobHUwK81bB758jN1w6nxC5cddxu3pEnGwsgVbfQG6lNqzTZkV
Q5t/tiXxiI0ELOZQ0l+AQ4B+fOiQJquav5acAPM/L2vLGFntRpV3Rc/4nE1ePXDr
eezrEM6aJ3Og7OQLsivMu+m/rI0M40Ewxsu2HUrv3Dfoifxuaa4X63/ASuehSldK
u0xl4dB3U2glO+P8wOCL7KVB3wm+Kr+uI1hWIMAG9Ao0LtOXDF6MlJugZq3BWEnP
jdLQfk+rf+2uQrhMCf5/6grnbTAkmEAELNgoFBKMVbklf4niJzcWbjgXABVugQ4l
KPBpqKZ79Y1z7Ax8m/4kww1CSpVJUwnI9OGIE/p3FVtx5zRkfFapXbLLBmcQbeuW
eEtR8YFYpYJtld8uf7levUW4FGCsuAhmjZN/agSQiT6XKpMhkKLB8m4tzmLIRS/4
166h32J4EALM4RryyBcaoSxgVFyDpVs08oTPQrFwPDA+0TEDdVRj6yJ0/RKPR1tE
IkSRIN/kuapprt1yTYg0bMI7+xXBgNojWkA8HdkGygDg75NeSAd+hPYPCzl8Izk0
F5TP7IG/UvU7EUmnG2J9NbDiKyRTdYmWhonwHiDR6oFslmu64L22JveR3VB/rqAu
FqA/dtS5pLazecv0mR74U9mbJ7z22ARRb7sMicBqpIrK2S4VVXt25b41Zpm3F4ni
BnwMIlC32hcS7S9YTiEspCbA5fKJUUz+afJwYN5hSGm4hijt2QsVi/SFqmzEX7uq
CrhZGvCqS/xUHgKBCY5PfX2802jgEmJ+Vq+d5VBESpYHUDAyTfWl4j93XRuuEM+c
8zv/ksU3k009a5wZSdbFoXcAnnCbT/aOJR3hkPJIqPPuYUCB8FVtzyYRxoZcAREx
OPFEi8kCDGIqQjwNBntLQxoeRS5ttQt6eCyZMEEm2tZOb6mrczE1tTPgc/7v8qcm
HqixKYq8I+eyKBaiQ0qAWYuBtS8pk9fnRgvPg+L7tghZBPSrhsUUL6yxurWl0q0Y
najlukXpxlWITOe7UinBWGmp3+Gct6EGAJqVG0FlWMDWF8ck2oGM3eof/S6ASr1y
SbP12P8SGEWy7k3Kg77VgHqStzKrT80LkYvfJTTBE0xgQC6DKm0rn36cNMoo799b
TeIkv2u/R1FlVt4hfe83Z0ZiKquMYXIoaKHaeGsN3hMyqF+4hNHWYMJa7zmI8+1I
pmvXpd7yLjVf5+/4qm51kn6NGcSViDtxodkCKtehdAno/b/wi+2C7QV5NSxezckh
NZUvo24FDWkqnyrD9mKYTdRrltjPnvFLVLEnvrRsLdmsP1za5DnZJM3l8yhMZ2Vr
wmzRfJxFG3X183B+r9sNea5iG4ufbqoDV2l6fzxsG/oWDeiUXdpV043TAlasEQEK
Er/fYscnHjo/QIc2aL3pQo0FVonyiYihbWdzpI8c9K0pQqBYVDKCsAPYkY0EFvzR
El6heIH8xBPQL4yOHvmqQ1o0ki+DxJoncOmoaWOM5hFfTi5D66ZyENKYb/s2v9Qx
pkxYQQM27BhCWMbf0NpDib/P8LDgUHsaxVOHoI9inZQdfTXeBol2r26rdd1Amro9
2VqRMKDUF18aSh2E0+zjWvwCJ3QORngEJEsY5rLlvMDeCPchSEiGa734KjnXhUVY
Sm+VB9BoHmrGhBB+vW2SxtLp1kaxa8iiAiQJgKEgeQsFkR0NOiA/tr19p8bCnBj0
uBQBON/IW7+qiWqmDKjXQLcU+pZJfTwqWtXCkPfDZ5DjjUP4RYnyhOBXNTEadL0y
uA/KmwmVKHlq6R9+hXWq1mqLmUefQv36SybY45zyRuaGpxAnAe/DzBRvjtPPJsBS
gzDx2xTCY04PjDeQO3q+cYk3Rq/KHSDXFrKhtvnOoLm3sa1A+KRJiJW9SmVSEmxz
s/GSKnnUWlc+yGYOed6Ku9Gd90+jJuwZGvxxJ7C7C6SV5H898EltthQwFkBfWP+5
rA06vRnxTaXpe/sPej8XBPAYp9GhJo0B+U9N8wyav+2li3gu9xUXMnxVrTMnDkBm
ZkhJUaQtKR1tpI+5oid+VQ2tMO/jUdJVPSNeJWjhtbrhKe1U7BctRzrbfLH1BIBK
OeGpcycC+HqeTEwjxQqu1FFAjaZswvpz9JBZY0xY85t2BGtAAxqLCCihI+8FyGCg
3EPU2P3Z5sFjMxzqW47KYMlFB4OO9K/rEf7M+biinI0Bl7E6yHsAeoDP21atxn2m
NGviCzrnLgfLbClWFunYMEFfKaEshe7K+O/S2L3ftUM6tFQG2tW6P1Bq9lbhz8U5
WnSiuktkZLtzuIyeXnvLdGhRljeZ/46LCmABmA4jLsBafPN3KPd9Ix9ydoTMK/Uj
YHTVadHnPRJ/Wfi4LzmqMeBAr0SpGUkVlnbZUc++8Pxy7rhw87H2gWPC/PxnbD3E
4xZEyElivrjAvbk63UtGv4bMpT7oa3DYg+6MNeS9zIL3cFHwToVFDFBSvMzVwCo3
eKDkwe5laN6r9U1JpscsYaYraHK8N/hYMUqH3tSwFF4o3829N0hLHK7B6Zj05UTH
R4vkJZaZ0aJ5GFE2yPivOKyMEDx1tUajkNGDZcY2BcdduSVZj8yyJ+Ef0iEAw0/J
yXZzKBva8tqVAza3D+SCYJNak2LIFQcVeq+3BDgJeq+THPVYTkoDd75pxM9vJnQC
7oMv/aGma/kUSnvVLhQ5FqRsWVtrS/OW4O+3z96NmhFavsh24ugExThjLJHWwE+m
CLVwbubJ+MHCY+aRFLdQmmKq4iODGSINC421ReGwY/RP7WIvzZRARw2iA9GdOu8i
ZIG2nf8Ch4PexXBBYVaynzMClkBwoEu9d10vPT7kv3xPQfylo/GYRcHJpoobG2im
hKlrIM7pz8rxUJlPZD1hhf6z9B++HK3NDHOdcTEQfuai8OuZDxuBG8r76aC5BovL
Kqm9bohohjsFUCjS4gF1ZopsTIcNX4euGlwwwxpC5aApuw+lYPEXAeFdVaM9GBte
fv2p8WvZpp/9FWm6md3HpzJF9qb1lE2kYbgdw9WnP3KFO/qzwHRQ+A2AGpbH92p9
48pvOCiBi+CtK9VAwUnle/cNzurPVjPJZacZIHXN966pyHxjBFAMNbkwEb+4jEyL
4jrvJMCC4cMBBWUPySTrulKwXqf+qO1QIkHU76wbbmjHN/b+Sb3qU+PiqtPa+5N0
wroOusMU3yQ0NYBJLtinw54kj1jXcXoFjkpeye8sOs6hDp6rIva3FPu8PMJD+/j4
y2RPihSMDBewiTk1vde87diz46Fy7SHGcLm/uR5HiNY2VZ5YNyzOv2BRjZX33lRH
FovE3WibhT8oBd6ZoHWeWJcU9bxdHs15mGFUCLZTVI9s5kSeV4Nv+uhQGJzf/MO3
S1JjYQ19hcnsYJt/ynPnw1eDeJElAlJmO9emMcNeZpj6/4SDm/p1x5blsO/LqL/3
up9EXCnunfeTPnQBsFpj6qGgtakRKS5wEst0treWHb4jWz6ucX5cH5ZcnG/HupvD
FRkcDDHnRtynn9hPaJbtH6JdJTyijvbaoRBgW5ZbezUpTxn+ByhASyZLtNpeSaNX
Y8ihaXE40aHvZOqwxzpezvoKmKNsAH8U8yPXlL9Satr7vPFogrOQbTCwDcHp+dp6
ZvctFQAxndBvmJFDSXlF9YSKvoew5tPkYinGfh9WjevO3sVf/uhLIwqlrj4oTT6u
DgZixCcyitTdXbPflT4kMLfBnQdEc6SrZqe+8OnWmdMxb2fFYhqjrQjot2yTim+O
8Ck7uvIFItnfufQ1SVg+ukfc4mx/dOTCkheMG8wK1u/Z6rG06ileTtYuhsXjXkjO
4Vpv6GoEFQCWHZ4deUQnWhUpWEC7h5fwDyDncdi9nRNF788Y4PGyHQHgi/YbNHlP
jEMjkHmwwEp1grWpkJD5AvUZa0dMqD2QnnQILrFpr08+mjbzaZp241XmSvWhihKG
k5wD73Wj+yvp1yWSxAZs8XM1c240DO8wcgKwysIlVKOn0E5zN8rcLP7g6OvRFunB
yG5wmFnxQSKJIBM/J7pHZpiQqg0KTI1D+MRn0KTlqkNXGWboP3Op2YOSgdieGDxr
jXxiaqSmYEDD2CvLM6/Mx+gE+rjqMp1dd411x8rDi8hLK70ML49nZOUZxlX8H50O
iqaSemwdtIeZpOcNACcVC7Bhpj+UA9xhc15nMmfty8aIuwUBnpF75Qpsf7LGbeVc
hdhk1/V5GyUo+b7npTZerkN0J2NaN2fys3FxF89kOclBXudNq2QBUVXo+ERbf9f+
5jkc3CXJf85ZHBPyzNukfxpWX6LiujL68+uZ3/MjNYVlSw4bK3XnK8LjASbF4chL
eVW1c6nraL1YnhhJijBYNSF4XsWl8dkkMDuIF9W1ASD+GkwZOp+GxXOcRm3N0D9U
/OADtV/nbpHj474d10HhEBVoh7DqO5iTUBxwJrLsKsfPqzx2aaYmVwkrEtuZLEzE
QK49QUOBPos8KIzlcAUIOy32cXfHefS9uaDDu9DZwGBvhsMq6aT5FTRz94Ksz8MU
4QRNPD+/PaPKbUGv5Tt5duPd7KvVbs3hjLuH/2boN2h5a8iPkIAbz5MMypTDB6hu
3T6soppdw9O/1x8klc8xvaYrG3mOS8jO0qRFy1je6cNbWrhDrT+N74ZKjoiq6ZV8
r2PUm+QoTrmij/GC7jvdpnVlcIyDXrfyvdVCRa1uUJ5Jj1I4QdZRFsbkW5zeK/J6
qyce9d2quUDc1+v99QuAAK5l/zELc7WiKLogQRJEuVa4YcejpAf9cU/XsVHHMPM2
NgL2tL3bz9i+LLnufpiviSm0NJwEGqOLiKApAxF8h19UOepvpylq4G917JyDy/gp
0I6IvVduxfoRBan2ZLDWNykmKMNH2EOPnNyzcOQyM91XnXEmbgWrEm7ZsCEYDzFX
uEdSb2YxwOpibamQt8lyn+rBKB1UoadhRXSEKb0TGEUShPcmG1/dVOg2wG+MGSuJ
Jx2bQ4AqKv50kgLVx5XGifxIfJvMLNnl6hN6T3Vj0duECltas9jnYpgWSpudP8x2
xgcs6dNpzJ6NE1ESZWSGj1wl67uihlYdG0/HWRFVk/0ocXv9yTMdqcoW+CGgsnuP
2QJYQyHhf9if3zGGkUECSkLu4xURnupRbiVSf1tw1L/mMMNgQQ8r8HCrnEy/oB/F
QJxqMtNt5oe4uPFHrUtx+HxrPaBqS6rP9yoV7iBZZm8Jgpeg9RUPNzFeo2THjw91
OlRyLc0DVtI898Xe1Bo7t4/GQf+8Dx1nocWzY2D2NA+BX/nG415dszh/nCGZCUT/
ZurpkTjl+Zx/QQE/ohh+PgyB0xaypYAVBck524xD+h/qjdENqATh5liiXuEbcvbT
073K4qwFHnP6auHtkKeIIzC23urI/U3oqiy0UwtMmbvmjEV29VxTBu8siEd0hZpM
U7DVdaYtqoJ9D9tieDnTD7RJze9yIa6uvK0TinOyvqvPNzbu+uEVPqvYsFGY8Bh1
3KWduBgRbGkUkceP+8WkYIfi04pdgXZtBXlL872Om3HJcOES8hW9N7nF4s4iPmyO
M+e/qG5Zmx77Por4cromrFMBMgzq79UlbeImRpKIhOP6Hr7WaIac3YmW64x4MHLW
wgptsIS26O46xbgfs2C6pBeXCyeS8DYNd9FWN4ZpFRnunWTBYxVj2WskyitIx8vo
Grerd2hlTdESmeyx1Qhi+ICzpXEuK9UA9682I2OXoklqggjt25KWZNeq1Chg6VkF
XTgUSbc5qem9GZupanPo5QTyeskOQmog9JXhZsON2IwUjOfV3v7tgbhX+oIXinI2
3Rqd6J+wrH22hR6+2XoKlovr7eQ8PdULfyaGNI3AaVNvu5NN0qzgvWz4bcazSGjC
vLF53fChPmt2mrqQ0D6x3eqZfmoIz+wgoEFB3FxXUTv777KgTfe3HizQTd1f8kPO
wDAGKAYAx/Ou9gioNn3BEMhVrdnejyHobFLMx+keKdjB/qK3qa3z34LgoyKMrFj9
mhQKgCPoMVcA9LL8+AmB6A8r0eaJ5GFOq9y7CaXA7FNb37eeP72CrvI/TRQp8ajT
AeQnuQt2LT0M+hlOff1QrjcA5vY5EtumgRp0dB6qRPY38LuhH/XHZzm8xN7P5adV
afwG2v3J/5SUaMbzZ2vF/1MWY8C5iRyl1PjHvZuuJ10A+qj8c8Tsf1PxIWWwoABH
f7PWqIXPXYBnPlObhFKWUPH0XbK5bjHX/BaOPaaP6MjsMXZhE6YDdELTIzHlxK8W
RADGPpozg5zYx7Q61RnwssoaL8iZj2MNWPKwqEc3OGmWvyqpEeTtzFdcV8Fb7U8p
4+m6uJ3qns55RCpizvJB3U/7bNwtAELyuIpQv+9XP50zPLjARGGuMsOQXN0Q3PO5
FRC2fsfqgEUqQOiijbnmWLhkYfeMuyu+nojqxRbOOEkMDk4Jbwbm2LSw3UcpZB5F
7/6mD2wVvUIqcDwvV1aNXzI/PH6ZTfa41ujku65UjxvWiisvAmCXwt3xDtD98ocO
QlXuN1D1jEaQirfdnPz8S2yTQdR1kYTCBVnwQHiDDB/1ZzEYjgHjYRZULi1CYhAK
I7CbSUwkzcsLjB0lpYvcKTtOdYClw7CGEzdygKxBBcbfplWevF7TGtyynQss3WK4
kYzegBK2TR5MVrPZdx7VxRe3s3cXdQHyC9zpUtMmQJqB58JlDzyU8MIhcmWhNsgK
ftqy3H1wPM6UgpBmt5E0pCIWrdM9YdELAroqw32VIxvO5dC8jHsOC58PVpkCDIGZ
CCAQflEuHpG453A/W3d1Ls0oKIT3Zc3UZrrf15AajssQOWM3KQm3yyZ4uGXRh0XQ
YEvErBwE0X/9JRnuomEhWabT2AnSgKUae7quiVcPznPJWp2BHze9zhtlAD1fLZ6i
5Plda38rP+IcIJsOqqjd1ZYnO5hogwX773/t552SZQm2//Tg9TsgOcTr564+ZokC
lHwVsp3QalQqpVqa7nxjQ3RITBP9LvtUVPfA2Y7Y9MWlpoabtkRlZBeHVpbWTN4o
x5HoGFeqGcw0pp07TxLSv+BjDQ7brcebVmYj/x3rtJEq6WNlFMN9zPgQ2JOTzKvq
bp+gtJMOMOEN15a5z/TQQ6Tpwkfz3pCdIifUiJZB2DwFDad8w1g7LgVAf0E7aLIK
PE3YXE8D363takMG1s3M3MLIlC5shKgswlk0RZPybVhN64/fMQ2A9ixwO0oldyy0
1TVj6PjcyxFaNv8tc+cLTpH5SuwNSFBVc9NU9ZY5ofuEU5jJdHXBKUHSQ+Q2WeDo
BeqyxZ8VF1bYF2oa/pWhwpGNPRNNOTfNLJvpXY3Urf77wszw43zCcD1NRMYtEUSn
2m07am2hWZx/FUvijCQ2WS1DuSXGs43E3cBOUIrKnJfOrs7BbHX6wr6BNN/b6t5s
hEOqlZwDgHZg+DX/IonEvWIF6VHb5yFNJ6u5UvnCXKNWpMmB3Lv8K9QxMe7oc5fv
HBaxN3ealQc2QPA4fRPZoZPM/K8UlK0Qg+Q/FJB5oM8VjWzmDfi8yPsiovRQyuF/
Xawes+FFnqp7vgNws7ZuGD+pueSYbhzJ5LCnpaBC/plt0BtIXFMzuGfMHs6HD7qs
IbRjnLEpgEUgwPAmc/xcROklS/pOncFoe0tCxQkdgCldRBz1TIPGqzdmiTOhNxLm
BNdMnnWNXpVCrzzS5gxcu45xKUjQKy3FffOJJnG9SuggxC/PsMVSxREpnPp15RwD
8LcnKGUgNsjKeKAC1V7xcuytocbLXxsC/sEDOpJed+8OsfR2FfSOJMRevmazf0HS
f0z+kxyoM4SOhtSTdlFqPw0gctTLiJ9fna+eRNyZ3t8athpBNdE4yo4UpQjQk06o
vtzbLpc4fznNIk1xYeYYccOpBo3ytfHFZd3ebbUuDgNmagM3L3Gsllfhzy4G5cjg
IvF1sMTrIIu7mWdKC5VaNwuCjsnWqAECDvk5xma/plcaM4OFBpLazL/twjArh5fx
8SJpMgqItnH7HvsyDBxlfxtN6ZPMeEpfej0rsxrN4sq4SUyVvFXp1c4jb/X52GLa
XacVHohHksW1b/AqOSCoVXY93glDz+4BiP73S/VYuyCcfyVLYLx8resRP3r3XFOz
252MleJWhAah0boKQ+0PQ2BrPbLNH3Mx8Be9uTnV+K5aTyeJVlhsNU2Yo4a3Qk33
a4328VH1vgWkzM4B6Jy8OkWNWqKGOW9Epcf+eJkuQtaqSd9FC0tnQ2yi3P+7cyyF
a3yhAP8hR5M61Y/1GFY+AEv/J390tShbMUGgGB+gwExu8sX5hvf2aIbA+28lGQR+
vJ/ko0jZP04Wjz/uhfGsHQAGKWUorYGO5fNRRCW1/tDD+wvJGtYRlUhwBHPl6LwV
sOYbA+41xEKfmp2VOAy2q326PqKZrVXr+Bm7W/84qmNknJGVUeLAu1hDNdo0KKBo
5vO89Ydn9Xku5MV9nI4P6wGzFQM57s4qoIapKs5ScFka74+MmEKxrPCjmyJkGjWg
bI0kl9Eqh5Q2uj0RZHgHc7BzyBLU3/I6cJkvmh+b4jpTas2RQCOyenvHkm1vIWv5
PGV9k1AsluBuEoBtOlqxyRWZzKKued+jTGzElsCYc91XecxNArCj+tO/Y3R/kTo3
MnjbYoDHda0fMU7MxWpb2FrUnVINUI1tQzdqhAD5dlQzWpwwcCqaLmReSgNa8v/o
Hh2YD3pWo/1TxAVUSHbDG65+xd2npGQkvZz8+J5nDEaFjNBZtHT/j1L1pdSYmXLZ
cILP8oJ5ETRDzfF+h1a9yFuouX9Nj1dud2b6+RoAwvppRDv1JWddqVQ6xW3yY4/Z
zOcqjr4/akY5o3+SSU4dd3uDqoeNZw2bz2SgR+96lgqo/phfjO93Nvmrp3DlNL9p
DiAwutR6CWAnBM8w9GsPc8lYP4GEx7kI/3GymCZDABsgz/QXVR5cPqi4Emwg7uit
PLd4Y3Ghb/swA+AFYhiegLIawmsOUo5X8zs9MeOyFEYZFq9ozq1/h7a3JtgYWiH3
n7w4wGudXfld13Oqx5GT9Mvz/F53AP19juW+jmyleca4UVOOCk8A7sMy8IOM/JhT
9tGhT9L4Y8ojiL0ZS6nGHxLfeYFBmnEX3JxUyLyZ6sBoZbZVbvz7hap6Aay7twIz
XAhZUGqLDrMv2g4gb8a0eGsjhsmBzrtQf+jJ6fu50XWtRAuVY3CucBfYSJwxjixV
Rh+TsV1IMQ/Y0NU0+HwaBW4Su6wbRKI+I/9MLNcThwg0b2CskhpCy3wi2MBdHV0w
3Y/r86W48pjVbvP5t+vhKSQYD4FhP/9FOeHrK99sfkpE2jsoRJuVPxZEb6PScI2q
1zKe7kME0Djtl/JcfG3tC/l1j1P/hsWj7V5ePr+BrQ/hKVw6OIC3px/a/Q9MxOQq
lypEiBQSEG7Fs2tzjDcZw9Dyjsnw6tErD6C3znlOsowbCSBlDlKqR8vvoOJq7I0H
+1uuhCyg800YGtEHl1niIW6UzSDNrg5TEDWdbPrIKvB4ItGWVQ51Q26vDfUKR3p2
8TFE6/mzwpKoydtIVljNOXmIIrO7rixJRkjp4tf0zX9AeLvqDSv+DBqABVyZ0VE/
usAWB0lhB66XzOv0nsvIs9k1D1b8FFgbThkKDCvvQsKbr7VW9toQzyvWuZlpP5rL
w7FDSczd5ZerGFVHtDtC8yNkMGTzcs+2+3NGCOw/r210ekipoOVMhW22xksjv+OE
6yjgMhIQ9kt0fjLpA8/aBb8wfEneeva0fgHMRuPKrQgHXzcJ6b3MXaeS32MGlJvJ
khqWl1RLscXzkqcq9YT7+CISfbgaxeXY6WExvgRmjoovxaGzVnUAnHQWaylijE2G
YAd2CyDWc+Y8FnD36LEIOKPYtuP0vSiSDjmuHfzw0AzRu4LutCmFWbn9lAVVSL9l
9CyBrFuSVaCPr/h0g2Xap3LfSzZyOBqwqSyIpHv0qPht2NlD8oUBQb/QWada2qxD
aaea3rEPWlEqQoyzkdR5kHwlc97f2viOkX+UsDm9xrKaOvmlTvoNp80fefDkjVBs
dwnL4Y+IyDH6aJaXoHldSpe8BZW8rC0aqX9Gl80qvHz8WL+QUvQbjhSTUAmAhIPm
JNbhverEZ+IuYaZz1Uf6KYEuNHn3Z/puwOHfnSxjtfMMK7rFirrK4857L0ZoL/is
kDfhGXBn13PuobgV9EKCRvDBbeSxv3nwQxhcs+piye5ppSzT2SRbMMxn+gvy6/DV
GuEdFEtg9xGVJvH68cxvXzqfz3ejFf9ZJSsY7IHl2CSvwer9KQz+fr9X51ZaJkxf
O0yAJa+9LNrECpUUhI7tdtCmiAjVZ3agO2RevThyaUEIn+gZKKWKaxe1TobyK1j+
ZnTCT7YV7olnQ2TvK7XblMD9ytAsrurU4vZeRGcTpmArBE8u4tEJ/hN/zOr0ahdS
R9+4n/v9WxYr57gqFeUHgCiQrc16ElIAIibm555I2Gxr6LNzfNkEZKZSejm6Hjpk
IymseqU40wE674OVY/onkCkKB+IGRWAPTQ6fzWyJlZYLTmyFBVhmGb1DJe1chBhU
UBttgRPwYtKpNr+qOSabD0onH3ATMzp3SlHll9dMuPoic5dzrqwM5Cs1GW5kogde
B/7J46VXkpbN5bVG9CqPfLsSShFZ+SVjpoZRr4gOYASYVvV7AkZKAPu0lgdYrmYs
wi6PGJGhySaah64sy0hjfxmgicP3HzHuol7aRY7vbgUxuNUQHkJ/Dw7hVGyWRQEx
u/ZacJ5IX8FPdoSpr8INKZb/iBChiBOlkI3Lq0sJlxfFF3PCziHEto4gtZRnTeEh
SdaLoFdU8FPNwaGlWAByohSkcBmr01iDEy1CIv+diUR0FF+n4261ukRNZkK9mGr/
TKM7qYSTyHm+lolnEJ2ZvfejKUAQysJEwBlmkTgvINtcJLOKrZa3j2cvNrwfTzDJ
RNmFIDWWP70JZXMdsN64nElrLZx382jm18W7ed5ajK/Ry5qzhNKNy23NbWKzPhNe
zrTLIsA7oNBsNpdrsHRZbKpwWE1fgQxZ5OUJj6VjPaMC4MKTb1vREkxmdOmPz8gH
MlXU5rwQva3WY7jCn2inOw3sEAGXw2E2sdw/tefb6Y+QMC2Nza/dEX8tNSHctZhp
wxT+z6hcZV+GNLD4Fdz7gqZeQKp5n5oZH1VxmqA2VANNZxsOovkx2OGDVc684sDF
1cAyznDHwXkqVlmwwtjJft/X4Tq6De1hs8dbyq1ZLWeorB3dDIlTvSpCIa6s397A
xhyLxrjQ5nx2b/8szBMdPCaWLiwp4OgC9Zi4nxq6yNAb6fiOkVSsUHZyWRdtCDzv
hFLV0qiZqi3QZsl/V9HDIkx7PNwGofmmASWJ34WUW5RCag+USZGV/iigv9K/UhiV
7/Yx1fqQomeq0GI0XTIacJj1MVX5KXdsquG6MR9ON9tzoB3p8MDROYHdEVbBUzSS
ECmtOlrXzadTsXpr3uUd9/+7ZC+S9P72cNJdxCALmVhhmZd0XrAwxKavx/jWWrIW
tOxcX+CwU9aNrJfNZ0keHBj9MgfIUhL72zmcsxzY2XmPi8ayam9X+2A1PcRDvD9t
wY9qDa0lgGu9iv5wI630U99pNgACDWGq454ZvOPVEnVb+uG/EVAat8JjXg/5aXpj
/167DH85vHej1mZdg5QyVOSoDEEmBKI+Es+bjj6WTCvojyY0ccmpSJ7qHTA/gECX
cqygtqCt3yNwFq65zakYWpnUBFI63+6qlTTzpmI+valMTgD1ITKVrkm0QVkZkMto
Ne30pH44L11Q9PJ9LiwsVOSRduc0+LJDZW0lJAS/QvGnZUjNRJPxjyhvQaLKV3ta
L+NbpXTC+Eo27bMHAYusTKXRk8iGQVx9LqE9kJeVbJzR3OcCIYhPhQCzfVXopGQf
5NhCjZwfYkRdx2NMMggLSJu7qgeczPIT8AsBtU7/l4at48TsGt8xCepAQgHVBmuC
RGMg2KHtJCMCEBCqyVuhzMgH30rdx07h65O0ut6DNf6nXEt1b5tm5k0kyW09dK28
Wi7q4GdZNwwuxQLLpc2vhCHyrj9XZH6KE+App2peTDBGTP/Qb6+Z5t9ecjTPnUsb
K48xRQcZUaFJh5Pfo8c45y+FVkBzvXf3KN6+BA8dTmjMfz/D06Nzt3BG3zfr2/D8
DFZyPVy4dertGa1Y/xD5vL6HMkTRwfe1GePCdmynGKKnY936IFrSx601ED0FbTHX
RSCupHJzBD9YT1iGQIt08RASE4lHHxkHcneR9JrBk1IR0MMb71IALofvZ9iP/eMs
6cln/JxAlUbZmYX+JYuYf/gx/zSdIrFvsB1kPYdrXsg0rI0iXYQWvp6QkKO8qqMe
AtCNw1ZDqpZp2L7gGYgmuMYDyyY0AOIoO8F+yS9X+mpBFXJIFyHLwrkhwqWYCmBY
Qe7fYy6w1Gvzgppj2vV6kx2EDNHIE5FOuDs5o1uKEJo+Jo2NUD3XZMwLrUW/qFy+
sLJ/AAvx59y/1D+p+yfmbVYMoNIH1UEaFnLWQpt90FdgynkivOnXdeDRdIkPAWK8
djRFHJl1s2Ge01kRx1wdWB/PblUULST40cuxA9mkSFx1Kjmb6V+TirhigVEkjPNs
sWmkKTdHTc1QCd6cltTHIQhZp1W0p7j6l65rvYwecP/FoNA2xacx7fJPg05nmMv4
sWKN21op1JnSV6eWRQojvOC4JnYjEuwPYDafwk0LSeGjATTg6sEVPPcl66WeFsIW
uuIKlxHFHadjSskuaYUGVPsY5yQ/7OOFfq0UniU029s3uq/k/kl1eKTUkZ/0p/E8
lk1OL1nrlp3FJQlQwyVqFde4mVrb0OxVWw/fp0NQ4L2fvHbC6jzV0loEc1Acmxw4
QZLp//xG4hqJELJFcr1w90FcbOR1tkfsLm7gBH3ZwZczqyB3vUoac8YI7PAWKFOv
+26IAfYK2hZykc6R/yfXmNhI0S7iQw5soggr6rafnYRsXcMmY3ZUPjSJV7tbDdwL
vrH2By359AmH0kjYbOmrgr6C/YqtuUCEygbzq8IJJdNGDqo2s6YQ9BMzhGfL23J9
qt8bpoqxPoR40lnSubAItbeOPsunu75cyaf+8i8byO4uoTJcaMlciqIdRkPjPpg1
xyrKZU8DybmA7nOKFBvt0Rm1yQ5vv9IeGAVTe277JF1hFkRQNxw2gpbUDZK89YUt
V4X1sTIjSlUXWQkX85idIvWbt/uWAyy9YgBIZxiMOWCQIzFGaD6bHLZwhrhSX/4B
uFy96uM8SEXXOcNbQGIPxRB3hvBiQdg5Di0z3uKN5+yvnglLuh7QZk2wGqlHE/qN
GJMd72Munup0/lQb9ZHsKsaOWnT1t7aidQhQ36d5NBiFb8gMi0Bn5U7xx3t/5XFn
m393i5XHuCLB9F80ZHFHyYG929Gs8PkgY2E/CSLb1cc0aIkVJYIpO9Z8ZtLLxf35
L+0WphHTFp39IwJKHLgTNpJ4xrbG0IqwVS+WuVMzzhSRjRBP8MjPE2hZ/WPZ1bpY
BDn5ERjQXeGeffz48jhd8bcZH2I8+Mzfu2KG8lnp+cxmygj9V8HuV6pFcKKygPXo
bpKV0YiNbhThqhZasDPKN+fSpTqbPJ5B7hN1aTGhOTYtwnDJS1tCQly32N9KK8qL
RmQz+jAu0jHIFgls5W7shY385WJnA7o/fU+QxjkTE4mK8NsE4L7U1oQYit7T5vQR
4vl/SoCLsZAQoxKD0BwBrPXJWyty5fuDL1GWMoThzib+mV3zpXQHe+rc49+w7dqg
i94CsuyB3E+TvVAw+p3/M605slQIdkuTgMtnar+73oKwXfomacQ9OZvumh/G3z43
IGJqJrpg7yAKEswfXzUYu6i5LRqwfjg6JwBQqmg6lnoPPHU6IXlf7cs3hwUbBOSp
jmUQzjiQx8FCOEF7/v+BP9tP7SUcB19t2vIw2HrSeCK9hpjso1QbywqU89pB20i5
TeOfzE3OGll/Wj5IPKbb9jHSegOOYE4pZUnD3FzpnVjFMoCbCyXLOcA5FkVuxYgd
XAgWHCm/9eZCrmNFvXooaX/r8orqdSMFwod0OV41J1OUPKOMniK8d8xy3A7nFCFP
aARIUrZaKjxKryya/rI2Cl15hrWbgu1jfbAEJOODSB/l4bAk6cXtNWsAJoSNZL9G
Jk6uRPg+be8ZZtIfTr3QJRc9li/qKrgf7GJpJoeyxpid30mptbII0iZAJphnQRMY
UA2CbpAME72XQwDgA/+0jfaLNaHEDf+CHUHDwM6GpqPD1HoxZL0eRn5+XbpqY3XX
TcTwkD2yOhxjXG1zIatLI5sfFG/A1sNruwkpZF46BTc3/cv/eLd+AZfHblLrX8xP
9dIg5tY8s5eiKWU1ISsqpFDApiG+qw58dYQFqdAReLO2DedL1aWva/8YgN+Ml5GH
BpeptSb9iGH2Iy8jNT9OpbDMig5yogstSgDIfsy1j/0VMDWLFmhnFIvxv8LUKWFG
VtqWPKp3Tx/xbm/o9TLE6IscaqAJifpxG176q9fDFGkW50h8rthLGRiblKcSZFF6
Z9hVkfGm02FQojUx9shGLVbuHkrEHcsrYhx5UkTBZZhAJbdXZ2tT1JkSl8tDtnGa
jDj3AlWGpZ6ocgI4o2665EBU7pxTvpLgy//JigK5ry1j9rqpDMoKbKpD3nj1xFyf
1c3+xTJcnyEQ0GdUJb5oPV2M664Xtdlu83tL8tVGiGsgVm8b5XdsUsyc4YMt3UC9
57LBWpg8Qp0m29XvDr+IirSXMtyqBg1BmHGg3hGVRUnZJ3TXrR2LyttYeFH3OMEM
6S2NeMrQBLvmgE769KlGv0HERrLMtGy6Kyl59jxihGIHU7Ee9Nz6jMV0Uv/xSYva
08/0gAtQuVJwGGeyjzCFRs5IheT57dtTvohTKCZ0JkCJmtZxOn67wmrREAZRYAQ8
yFIedbuzABuNVSVP6folQOrce1a6t5yroxhFrCXlfms9aH7Dtbdow+vVxej4w7rF
bysEKylLw6NpFLctrve6JHyGi663AT1wXmgKvLp+21AMWqLktf9NE7dMndd5/Pkt
cHmqEL7F97Fw2FdfMh5GBDissNkMWUF9aPWFT15SP+/7FFK06PtGochcdn+bF8qx
xp2orYdoQgpTP2wCkZX2ac/bydw2JSFvVi6C09hYDqw7lk76VNjCTDIi9VjiBC5r
L0Cm5ykv5j81SJPVa6UfKX8w+91rnMBvnsqI0WpKmwulUcdBVQm00wD4yD2TvdmE
2rN6snyAbyexmfyE0fZEbQ+EJ5zu4coZun6K3s+K5qtEeu0K63bzmWcsw4edUhP5
3XAtZsZTs8N6ziChURUfRoevO3y3ABOQUf06X9JNQfK2kHXYILiPGgqGfWZFwzMb
L0eWpQvpeOq9LJ0my9fXare0H80PUGRiSk/cT7WXL5QyTsSH/pVrVMBq2kFrc/9p
NGU0Mk/k/NZjfp2khZAqSvtbYpLPzW1VeIfwu6lySYAnOxlJ4bctZAqEHGqw6QEv
SjvyaUfv07u4pEkDtJx/9HXMdlDMRjf8++8206cP5ELOKL42jC3gxB/2JEppNhm2
Wx5/ZM29vUqP6eEZmwKvaAxl0r2wEObkZsY2UCa3LXuMAjn9pH88lTh4F0VjDfRo
ETBWawCo2LzWOfBowL7eEA6IAlyA8mg9qn6rTIjRljRFZ9Psv6zUQZ6la4uIDorY
E9RAphUXxIPioBFTCZZgN5x47IrI/F+BN24CrZZA8Nsa45A5lGpvYe3sPY2dChBN
uwe4ojav4L/paYUcGLbAKKvMOaitQ5fFgLZ1HrThY5LT1Lo5ZR4YcVEAUiFwg8mU
+pduCOWovejSYfCtyJWiLMlsSrOn1ZUh5LsikGBlDQX0g00ZWZCezq4pfWQJ8Kv1
m2aBunQtItvP+qCwJdZstViRdjx8J4fxm2xinkE8nYibRnjvbWZkxg8uUuB1NVlN
RVl6OYVy8lYZB3QZxAPpQOxA9c5DA7daYpTW31ycnLCRTCJzudY2Qhfggqd8pK/U
VluXcz8SXN+Oh20SQ9Zyx0Wqm8FEO6OirXfdEO8f+odKGEEmz0zCGIvP9DQbPvzH
C2xphTrsYtT3Ezxhu/qPDc2F2zALsS0UcKyuBOZ/xNUyUoE+Bq1zNdvtDdcJgtLI
Gz2Vdas26rLFRfWRF8CZGr6OvCN6gH9wrWBsgnoIFAzk/UMwoInAbMiBJW0URTbK
G23wehW0MJXIk+PfDETz9pyVZpaRm8AP0ZTl2ToPxxiD63pVDpSlnaXR744Q7UP1
niLkfHMfsgqVP8EUVnZ5VgRHH7G1/iMYje4fyPHIhOOp9Pc1AEC+LvqYp7PiZiYW
iPxYXIyBQbcDv4YBKJXdb3GT8hQa77sgPP+XngB3nfT3fJRFQNimv71mqTrfVDbL
GQaDoezSqpXaRSTPS4lnDC01t1jhqGHv16HATWe7hmshZIZbSLOH9sNQ4PCxARix
kfv4TEhkxcmFlRKV5ON0yEreLa3LPqpStbDpRlZkeCkMWzRQYT1OVjCLpwJQvHSl
ZvxAinxMBFHmVCYbcwfsz8pRuNwN1bxIx9YSHLz6yEAjvbVQM00ygWxSCMpj5GNu
X98ndMvbyjE7tLmeo5q9BhaJqI1HETlnsz6cAntu/s8eAixM6odqc8qKcjLoX6LP
PV5LDad6NVsE8scBoJvclF1vdNroLYgpC7tBxgqUu82yOweMdLNklJ18JTDHBvNl
XwqUH1bujXefTOjnE8P1lZyGBAVQrfEVjg9cXhZfkB2WCx2YP4nsuzwpN+VZs42y
R06EQZD3TcZHuBQrZhVMrbWFeg6eUF4vZZ1o/PEXUf2MXXXce8QkxR/LnF/0oHkz
vKTK4UA9UqVrJC4+iygDg4chaWZIj4MbVgq1l76DSNHXQl9qeizJQzipncEBuzgq
9aMs2hrx05G2E+gZHp0PqMUR/0RadAC9/59dkZNKdcVl4jazybetXvuGRbo/xkQF
twJ5yBG5XMFXUie/soFVYYNLhgXPd+xt/bZnuEt3J6VM/1/j1wevfKC8HnbHd7uv
LJ3eMuqbjiJnZqSwlAygHkj8K3tdE6f7MVv6hZUX+VHdBsMbAmt9xTqyqbRfrPHx
g2cdgLQQ2dqS2byDd2louh+CQYRJQEVa19a3Gfr5anvr7jmfxkKXNMh8xdpusJi8
PLYAfMrWrW01ignKu/JhmePYQylYPsIzFmKhJaOdjq33hgWYujEoLDfWJHDZjBXU
OzbWTyVMbqQEhVAtFklfgXGEsg4bn0bCFP2olhnaDSnIsGVvehJejZDIO8mldf/1
T+KyqkXuBrA5WZPDb8Q4o+1E6l26FwNbzYtp7Z7I+SlKFG2L80KCNso+XxU8YxhT
1gMaUHTHfWIRzn1HWkt7/F/YyDGFPveDDn/ZiucwQDYy/eqkJJSz/nQE9u2qkAMW
4yVWk+6KnFRY9HR9vpzCJFNgbm1tGZxxhsv02u+jJysH0TrrWctACcnrR4jMy5S0
FCXRqAZmbQb9QlDiv2a3UM8BDMNCXzhSNQziRVzbfVPRLIt9i1gmrxbJbAruvA+A
wqunaNTRLxgM3vafimk4f3tK6Kn7MokZsTE3F3bAwOqx431O0LUpnQeOzk1SMS83
veLMJ4T9ZEnWFM4zg+pOPKZp5Eo8O8wzwdNiT8ADRRKJD0pf1XR1HG9C9hCrttfy
Yc6tjx4fa3K1dTMyuj5/R2GbpWUV1AkobpqDTdcfQvWIDKL8MfCPsIxgmg991q1q
qafH/l8jOm9ZGLIQbL4pI0qxT3DDXu/3KrUmKIxOJOhi+djO3QVYZIIG0g3yxGVU
6Vd4ViFWfhCYTywE3VipIMN98xp4FoxWchkF5BtQLm9+u3pEbt/OgR+sGqsKt4k2
qBaf2JPuNCG10wd4EFS/p1ssfK7rrzSzffefvhL3GWDjbR6zo+LzWLPz9l4WVDNT
qWuUNVpjkGBSRoOSivIy+R8J+Gyqq+Ka8I20RnnLuHRdhOWCMPRlSFfPdsDm5iJ/
3LI+lkLYuveppE9+MQRjFAFckLEoViUyG1zgSx7MYdPtl9r4dknRHkgzyK65ta2a
vnEg7dNLZRc5UT8byakPZX3kkqWv9prQlaq45C/2ArlQEifoCw0vQTy707ZRJmCE
ukXbuBIpK1ons7e1o9306+9brEm1JqJWemAktwpGBiUYCBMuMe/qu6pr5s2kzBQ6
OMl7jKOrBmtabB/1gsO5sHcI4kDYD2Gzv4qRsEXTH/wQoKUg62Nf90byojy2roGP
VIBiCY6h6G84bdMWkzeVydQoOl/djM14dWKMIO0L4/mA7VIKG1dKgBZ9gT8J5yMi
b8cFB2EQkbEW55bfUZ9mad9pJD9qelE+cg4kcLDZ+XF15IJjqbEr7y+My0N6rGiJ
WzlkuqFUFfvpq01f87fX+l8WsF3v7QRNsCwt7ru5D1Osp+/3mHQtceVa1BMLOKRr
DU/rt9QQ0Bc6zfyRkolhki/zRdU0tCp1sr5Xogo9DcwFiBPXm5bjRzD5FofV2cr9
yy1UB7x6b8KhE+QXVZ8y1qCF/AZW4wgWgjxsaYkLExKoCWi4EVJyEXFimm5WNDVG
NJD00nh53/7JU/gEkawlP2NRQd2+h6ntg8vqA7kZDgmWwsbUsIfPViZaRvf2zKfG
tL3XCK+SGqL6Tkx72UrGHuZ7hp/wywo1gOMAGirjIrQOZIv4iidCDsVj092+R3gw
G175sCDE4FhLleyCGtMs2DlJRumfOIwp3ES2xJxPu2gZj+FVb1izCFH/NiGTR5nE
ZgJRikPM5bhpFLJzMsjFZLiaB7ha71QrlJ0MrFoer9+Rs4dUrY2UGM2X79EtE8MR
ML9HmA4ETBqATDTVK4Zm6CsFEE1q+jkLr+pnQyyqoKyWNTgaKic4dRbLv4+Q+dlO
/eCc2omCs8Jciwc3nDS33xECh45cDkeFuav1M456ny2Zu6sf8wpH37XdOxYXLTwZ
1CLnRQ7ir5zZtUV8njC+NEJnrtjbxCklJDQZG1UheyrA8onR3I3DfPl2SeNGExpe
WRa4I5aSj3mPfsiFUeBauGDNsxmkSVGHFPrMt3GyR0nUZzb/HoWYJfeIlo9NGsOR
SU/3SLXGdG6duMet5Gm0UFok3JUmOjgW+BiziKUnQ1c8+i39HeLbIEnCgTJkXD0K
BYYxxusaorgHhQVt4+9pku8IL0Rn+z1OPFpMdTn4f79LY6hoKkjszHuF7caA63ZM
N/sxnnGU9h9zgWITL73SsI0QZlrYr6yHq3d8iNlRkHPgxUaSaa1s437XNe5MEsgl
SPrteAsm3ZQ2ULQzjroNl4fHXF2OaJNUGejh8jyOelj2jkk16di1tG2hFnUw/KZu
BhAsdDkhJWA8BLZcE53pbGTFDkfrCIg1FYqsDpDUxqX+qlu37igpw1mRkYkMRfln
gbepelrrcrfeCq/KpZUrRAA7qbBsZqm77I5hZKCFMyPN10x8/0SmCa/zjEGuxDc+
ziJKayNUsenlhFHzB4+U0CNl5pirbz93GZK+2ecRc2ptOFqt8MkV+qs+kLJ70ldo
cP8ByrHIhbQ3AgVn3ihJKbPiiWyWXegTtWkd1Rz0gfC4YM0I01vuwOW5WJJfxfPX
qICvPXgjNyEk+JSQ/csSmdKt0FgVE+INcYhTaQzmkpOH/SShsx8pqNbo61FwSdAE
uLK5yIih+7R8XTrC1gcSRFxUZEhd1aDYMABS8ROvLHjHGy9k26nZrPHhdyU4DSWG
Uz2kdWZC9tORokpSDKepr+1O87oSnid17paEfQ87174OetVlLOoBF9pHky4R6uWo
u7nkXXrYiMjVmDBUrzuxs9f7eR+1q8dKWTo+Y808FU6l6Nx1sALG3DNZebknSI1a
mMhixhdcx2SBfvMok7S9wX9hS22SMEn/yYRvgiZtl/tz6pVEf866UE6Ae3/RvkUi
GIzPR2G6oCXe41e8coPpRSqSb0KBlb7WKqjy6LO0e8DgbzKhA2iM86ZWLc6DSZY0
zm8u8ugI6fYVWYgI6P2M7REQLYce2ktoINGrPLJlowN0xAE4qjuj5GO1eqBdMvSW
zkvaAsGawIbDEw27565aPX1RuJ0Az7fZOQ3digcWoh2pJx4TTb7jhW39agSC3HZw
O2GmJ2Js1RXIeTgOPspEUliurTxJUdPMT4zjTL13pTSpLItmT+ggejn94VRKkqIF
gTBTH6ZiD4x/RwcvONiXT6eQvqKAJQnHPxl96jXvVm5xGUEL9S9TNRCiGusgMNKk
iMhfbkgaCbcytgosSe2wTWTZdzj5SnJ//tKJ+draBYpmJ3ZZlhEE8OO3qvhV4vZ5
Y0nRxj4l/GdOLhbeT5KsjlkDM3lUYNyRP+NuIMR6iPQZjHz81SDHhWtgFbDk8dHh
BG3gdo6F62dRfLg5QatFILweYHiifKjJWtU8s+6LnuFYCvLUrMr7+60ifT1m2eGo
MqWc7mOaA62n4rWk6mmiefU4GF7BjAtiwikXfCbN8w3caCAqjdPh2I5NDkUd2L/3
uwis/hmZ5+p7d2ptwP3ZEtAitB+JTbGnP6/R4mO3eBbnPEPERXiz4ooZ5xuxva+r
2i45BIsDLpa+SOX1HPn/WlsKRaF6OcYxpjLrD+prnVnLeST7sj/2iZ064ukWhh5G
S/icNp7Z8El63DADnKQYDxPiNpVFCJFCVzDF2Fzwiv+AIPEBFKOvXKtX7a1i9RC9
DpT+pbTIoUeR6G1Kx/5wJDP4+S0Cl07fNVosGW7zhrqWxm9LEFHAfFTjYbe8RVyR
dO98QBCnWh5OyPTv9fRo8YdutpxPVrPHNDdC40E4ct68YoERhEdCS95NdTaJhpS1
u2eeXsjaCEjnZCYBK6+D1DaE3e/mJ5MFSNWU1oVZcUNv24eqfEsHHM0HifwFmkTB
iPrWWdw5887N2IxpOnPmdcxWQKe3zrT3UTGvehG0jdO60+3le8Emm+Ra73ypvkOS
hpiBmCTIWRRbD1kZ7rNVBswjmARH/XF6SonvukmHeyHG/YNzyOzD7kHxn4EQNFS3
1chgpihP2looECcscCARbbWgOybADqM6AgioWNfA530+9QM3Vv8+KqDwCgWiAqFG
O76EcXF40JAKSVHv/G5cqp/NNgeAbXGpbKBUvxxC9eN2mRX3DDWJ87HbKlWJCwz4
2TfLSFmCYZ3p2KDiJOH0UtozTbtC2lfcCuWmy0T2WNjDZYWxoyopISXaMVBBcBsS
g7VXYTkUg8pwrtH41oOpAPwa3KlaUdJNIu7uqZhYt1f7vgejmfwJTx+Xoa3mlOGs
PWUYdsAcupyvHOs4F3GJWBj0RC94x/hemuhgcieh3hYAotc/izT5uQQU1KBKhHU6
ixLXNEZjnkqHR73jeN1WKMWcVnD2HtymRcsHdo1+ybf0WxYexjUgKKJMGZ2bUrzS
PE4PBf0wQTfFbPiczitZwlEBEsqbzf33N7+LEyuxzUSJeXp7tRCgtkGU3RKSJTQF
Bozcu5En+GGv0v7S8kPpYjWxl0HykpslVNvU6B/bvxOCW61q95QuYw4QQC+5fdTP
EYh13OfY2A0NUg7FjZydbJfrbCYc5Zvw2b4VeP3F75swyszTRqGj6iYfAeSG7IJM
UTTHvGV9ekG6p4golAGJ+S3103vfMdZl0XirLrt1NuQ3YuVEeejiWFDYrslpZzX0
7r1OuvxP1omTt2Z8UkzX70XRRRjMGarxRVsajtfOk/rgQ0D8dGAUwUt7zDqH5voz
0K5sbHSy2FrXJj9CaBVmXvsizj3QBDr2d6LWHoLJGkPlhiHwJB9CqK0vJm/WUNR+
ARzaXMzWXYXESTIdilDmkv5S10WQMR6KVGCruRYbAeSj1kkfKmYbqp8r0KWbqWg2
Qk9LzuoF8qWuyCvIyDpugvqm64fMzDJHYsmT8wDjO3niNTpTzCN3etRXRWYaZv9S
lgYQn1htOPli9fTAgwnEeawRG3ZIMmA6FCcM5P5GR0JNgHqtwUnmeCnGBB65sGHX
vKoN7IEoc9Up+k7eEBcsebcaOmgR5Nl0tnSX0PY4RUptDvgnbaTzZJ6RTfvEec1f
WQNIoPv0AmKxjgyh+z5stMJpNGuYnuMOmPfdimHB7DZvedVYgCElp0PpbqRcpVuO
2VZXPc6EzWllWlLO+eDbPMCNo28L4k0kZDQ7i0L2gG0wagJUFyOfFtcedgVIG2ce
LCXT0go2RrYpMhp05WBiLqe59C4dUqBF25M4txhnF1wih1VZAvkcMX+mLEh7kSuf
cGZDbFR2HyeercAjowVy/ObDQ+3SZdOdCgkTREARD3S4lybWl7/Mz0HPM7RaWWT2
/9kRZNulWQTsSC1oE9KPPBrbXFVTd2ZrvxIHzmZWuFfhWgVEbCOro0yCeP453C+O
vWlpEEMPG55tzFFO1ru5E1mYqkpL9OtwD73lTLmudlqUyK5Ap9RXb3k6sMyvmCGF
RZA8NMRcDo56zbWwBCjjAuc021UzSFHaTuOZeTKeXz0J5XdSG6xGV536NHvxrKIE
ecllnIZWOfmX8Gt4uc+UUP4hORE0T5Zz9b1YpU6yeCcShy+UlqYfvOwi5mdhBmLd
CApBq/uEk0mUTlVySQzAzt3q4VSMS+N2J5un18zxmHEz/E4BT3EiJ1zqo+OyhKjA
WYSXp0jZxapyne0jcYc3iujkporGzZ5MwTk92RCzVzSLLRQ1TYnoxEeHh4y7w+Hm
G5Iuj6uqMjln/YLSsoGvYhZ1PMKwGCFOYJrOmYolEEmHsicT2tqj3aZOnk9W0xLe
rWtcTqbjqN4tBE3SyVqlzS72b3aaB/2iH4+UBX9XJ2jsWfJluaty/YdUaQ0n8s1V
trA3qk8wiAgQgh1nJb0oJwtCx2v70YDmTWDsijNIRDu08U1oNFiK6N0Oakjuf0St
PtRTgA+M1lXHoTknrmNYfBXlsrSR64EJjMsOFEbvXfmiLKehuD0dx1y82oybu/M6
KPulAgnLg+qGvJlYO5KT/V52jMG/7Mq6GkzFDQxGqE8euy7+sfJIBvoMFX4pgU2V
eoscTAUycRWjWAhh7BclrQNEdNn86n/vh9jDHMebu7s0tz9AARvkoz3y/tXWq0xB
Ogq0netnUPWOJZgsOrqd5QyExa1+UQSgkEledrVvgHg+eiQdzK7kN6/p5zbkixsg
AJmt+qpwMQBAMXfAyiubW2hVM+T/nG0izxuf62ArhLxq3nCyddVU1FoaB5y7kGei
liK0f3wC32JHeRCcBjZ9T+LwXc6Nb+z7961PoobncdHw7Dh7k5/g/U/wbBtTbk5J
fbgwv+jSjHEPTLEtyTO4rifX5OMl04uviaNTv+hCDXCk9OaAYS3WNAax5YM0irfh
auNScZKU+5jdXdQLLsi3fjxpEyFlrvlywUsCP6UxNXK1ZYUyISEQrX9d9TcHaWAP
tmwsgS43mdZe3xbrivWaiWt3BVtJdyFG4rttfVIhGn4A0GoPiAPQUcJ0xZqrua4w
cLhB7IrW1JuxnPlRQguuVB2VTwOrLQ+2Uthqb7lbI6O47YsQXC1/Cf5R+YxpYvq6
vfLUw3LboPuu5HtaaemDekLxeS43c/N7T2H3HsvMIMxNTYA3dFJhdLY46Ht4PlVs
8l522eCyyEkd+l8uPSkh5bZDXD9x0FFg7dTgtSi3t4jda3t7G//eoMvSk4RLEZpp
MHFLFAM8sNnlHP6tNao+6+hrJhIlKfvrNhK/+66+dMRQqbK41t90I1q3lVoZmOF+
F/a3haMn+Ya4Oli+LtaG2fo3vvUMDF1bQkcULERHjmlQQjNNzhlcTQwQxUM9r1d4
8IWdsEviNHhR0oBsJpajJK9J1r+mwpJU2X0E7v1j8jjxG0E+P8ky+f1UARSG4hU8
TYwBd9bK+K3xoqiSTpJLl50vNsN3oJanQu/hnER9kxswHJzIceI7Nj/ngrInSxST
vpXP1uOPSVR2XhW2GgDQZtf2Q4y+Ovwb0PRxFbAWFQUzIVq/8WbFaDdN/BbXwmSB
0Isz9gt9qfVJWELFVTDqDgjDev0EHVK19ePEKaH+ooMSssiyYgSyssDVjzo6oIUC
YtVuhyhRyPEjci/TSqdelXJYbzGJ9NRMS69Y2aqErqfIPAg5ydjirEXCu0f2IL/f
bgVd58iWDsx3gf2WdOZLOl6H+xsTbkXxz51iu/YjCV89j/QYq8kQzHRrNWcw6qNK
NWmu7PlhTXIibgDcY17Seej5EGoBeOewoySNr55875kwL/ifrbGyti1Z51YQmcJU
h3XJ5qJgXuMaUIlc9ZCAbOpRFyaPNhmXIMwaFaklHQbgyvL4DJtrH3h+hGPGSkjm
qrInv0tvPmAvGul7ATGLX/SjfNEB0EDSFWJ0sFAX0v+Hepg18TUCJVeZsfc9xNOA
zGSWEtkoBrXuswkL4GLnaHQMi887ND7JdbeexhbvJHo1qT+wR1RODg8xW/PNst74
hVi+y0hsKWhPqSUhLtYSb1+atGduZy/RLW4cGJ5WFt4qYa/A8/cwQPplCY4Zlumj
/YE8OBsm179JOYo1CG4TQdUEbiOem2tmUyyUGgx+/iwoI+rHss1lUEVd59OnHEzc
rdvpb0ixMzGTfK/ekjc1On87yOTy7mZn2E5axqBpRHMjQQt/Lz9w4kcImz8GpfJJ
ahdFM7qKzeZO4tSJCiRijll6au9UcXpyJaX0mwz3CHatY9dDJRN9g5Uaj+6IQbPP
4xSGe3C28b0lc3c4K4ciMx7azRzRwoo+hUALMMJUI8xeDfXFfRfeIMuYCUhVtK1t
cSXArcGIs/o5mu/2MXg8sMXlj7P1atC+8wyIu9e2+6wPjYY1e8j3UMO0dSrbJK9p
ZG9DvVbbVlA8M0mgt9amBhKsi0MCXsRQydPtswyQWS01jW7BISm7dZMPEBbNA7YZ
Jb2Yg+2elIKSGVUymNbUs1xVyzruAQfKVw2LM83ikWWQRjeJmuZhhSkZ00mrbXCr
d8ZkLMmbEdiEB78DyNYebz1soO9hGRj5+Ooa0gRUnbEGuGpn5x2RPY+6n9yaV0Ol
wN+w+wnNs/jx4OG6JjDghzVBWjSGPg6Qwd9MxZQ8ubeTpUZVF/aJqftB1y77uv4A
OGS7ov/B+WBpxxia7IndvnG9PRxQT4n1DuzcW47qFjh7/F/kT39gnzOv7nz8hlhK
IrB3pZq0zqHt3bsAEI7/MFPRuXePg0cIIwAQijnUOr0ZSDFM0FIoqueNgrWIeBlU
mDG1Z8B1TjhQNHftC5cGhLk10GI413QliU608MlvRDCTsgODtDk1yqEA5LRPqOcH
RGR7tQoofeTy3ITd7icjtG/74pB9/bqA6wTrQeWobyphbyopvXK/c8gIoPcn7tGI
k/m2awcecAjdRwstnGnw9y7ADLZTBa0HPJ8RzmOYBspWaHCjQnBowc9E1tWv1bUZ
kvxFHQMGj7mXsKvuF6RXwiK89WLP4+zMoGi/aFaPDV4ncfJPMywuWxfkL+0bfK3S
GhvBF1gngsi5L1GIGMo1KIOC/FmPMace1xj1ippRPdUTSObvDL4bqzdRRHRZcXDs
c0xml3j1bY+bRmIlboPk2B+s/mrf+cIQHkIQFBM+PNTu2BEVGCtlH6mmiyNGELFT
lAoP4bq2gBVVQ1oe+AEYEhXeVreto1YDa6CYACWN582gERIbtsL+OXQB/G6SQJVK
/zbNQ9NS7DKwFAh7Kg54XKz9X07KOiCll/1DSMwtNSgaJ7hcLgvPFkrqy0wpCjsX
h49BWN8v8YR7H9/hRuohtBmLnG7IzFTa1R/bBUKUy7FGpb6kDnhaEBnjvUitdanp
ZkzVPGBSIfPthON+flOyJm+/ZdONhPtOOXEsA7DHO+/6yQIw7CJeCpnBK8phBS6e
ovr5TTIgpL84bOkLqed20Ut31Aq4FPsOrOxPz95Y5Fkx7cgRoxv77nllXK70R8OW
2uiCfBdb851zfb6zn4YvEyfes4cK3d/ZB5HVbTqKG2Ea2c4P5r3T90895HYTQxQv
XZVaWLUmgdH/87gqAbBuwjgGbS0qxAqybEwQ7webgCA=

`pragma protect end_protected
