// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
RgXo7SgqLi7PhQ1DSE49oRDgBhqhTZKLUwFoZfppDT1ToJrl2QO0GdyleeVBV1oP
aJzMB5YWdGTybHxg8ZSgbZETcWHhSy38pQTPbnKSfZi3DT8qDB5WQ9H5z/P4MX3E
cgzXm6EcZM/ZSwsBAy3COBLJJDv1dfbVCpNIi1GIYGM=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 76880 )
`pragma protect data_block
WgeIuOj3MdONSudIY0QRTz3YbJ9Zin33jXWHAhSwE6Gd1zNNahim7xFXcNj3I3mU
iXkEso4mEA7iSeplbhjSzbpUVcKvcajF5OYbqEqTm+WT3UWzjcUdexBLXwZ/8xYx
irhwTQCVysMVd+N093gnFGRgo4V9PKpY/Nke36n8nmAbvh0TzKeuD1IFsSCH/PDV
C4TE/0z/AQI7vJXzubIYhUqb+3uUxQl54y9Lq1h2EVxRGYgnY/mia5g0Z7eFL4Nt
ZlIuFJehpAwJFYRx+2BVEpogECK4oPpjfLgC0+wyT163DGr+bNra6A3j3gkkV4b/
onhDHvPD8oQlfg0fMECSIYWSa36RTnOLLoY6HYz1gMNNycEROka3m3JmvHknRHoQ
iQDZOWB5V/sqzSL28KmU82oBXSauAB/WSn2nJnqHk6xB8S0qAoLcJjEL4LLTYe8U
Il0iHGYDcWGq4uU/+L+9GniC+fOuv0PHYfBDTmZpVDHb5DljZJ/N+oiZtyzybgOA
ehY63trD382qL3sawwGyIVS8ZaALpqsiasiCqxPqygm4pr7zBl6syAZiFTf6OjLO
dyM9K3jzrUYLz1cWka5lICuw5RG4im0QJwEH3BouErOS9UPqbyqvDgosCfIkHTON
3rnWCKmIWsDXlN5l7Y8LaOjAB0sJHQ2dhV74mA8pDeWSGUJWjrEmlSumieh5W1eP
R8ii2GpLyLci+VYB0qi0/xmAJcW+zZaIprDkWoDe77OX3M7OQBznt3B41xGZZoX4
nHa42/q6bjRmAz1izanIF57tKRK/j5iO4fdJ6GRHMLCQHGdLOc22t74ddRFE3KVB
CimKqQkz+NgACgWBYa8bcXl2ZXZKa1oYgtbeA68SJYECQw/Jg7M9vht94WZCVmd8
X2OJqZKH84aOYe+AwgTR0LJp7JlbysBski5hwjGoWMkpaG010RYZrEjcjrQBntaa
0Z7n5+H0GWKgOTouxcyY9Yu+BiTo4RP9aUQHdYHNcmkLPpAZ5tVpnMCTY/w9zS1y
E5hmKm/zfh18h/1TFMxUr/1NCkh90JlR3rCiYhydMm9QnzCmCz1C1Rt6YpACu96l
3lEcWfi7cZZafX7oVop7Tz3qfeA++pW2TkAUey2dKRmz3Pvg3MZAUNK+WFqaF68e
7nvSvIAgxs/l/O6BwNdqvV+Wg5Y4vF1+PIw8syE4qMkzaqfdSwk+iAY2NcPCHVl3
0FVBZY0O/Surj0zVCN7pEzpbi5R4AQB/5VZAtQmzv0j6AIGBDPfbLjT8pPy+/OpD
MoKIFYphcIZPYKufzGQW5wfk/fxgRnz32YtxMkjvEXg3jU/2YE9S1dQ8hAeWUVQk
fh7C5MCzV8/DJCyqqyxFj8d6Ul0upowWHnD1iwbWU4Uh5LRwcmWbxAvIFUg4B/M7
5Fx1RFKH1yJKwunCsttwheEWXh0vgERUjL0C/Q2kHwqBRUk0nBdEjxuYqB5tBRMV
Bka7FRbZFEgauKLozOx4hIL9ybNO36B7Jg6JaHOviH3dRtfnbWBl89BNy1vgMhE4
kAR2OQgl4PtttIbBpxetQ94PD9GPdrQEjwKjFuKsFHN8NHy50sBLk4C+tXGZbhLb
/I0QH6xJ7Dvj0LdPLcZiSrCpuo8/Ap+FgBQd4tKKPUtFTgPIL2VBPRh0Kg8O2Q38
7KjpApob9DG1gGDGZawM2mhXmhfQHikoJqILXyw0SlFghCazdqJj4Wg6F4sqyzs4
V361N+Ifn9oRNhL4MmDGxE8cW6TK+CxoLQQipxr1/wPHSngue5HxDS5DjmYXAwGG
eDxaXUu+NeBrYwAyxfNWJ0QlCf3UG41yC4DrX7kVeNT6PiG87x28ADUFKSZIjQtj
XBiStQfpWWNKklo0f5hZBGY2PEdwuy5+UNr5QFYIDnzJWQJG6VU6ALMOS3XE2BZU
CpcNm2q79RkB15DjBesxgv4XQegtBLxCjflh69w6d9bNAYmVGjjRtWfX4mlVulaJ
n90JCY2ecjmhI9+fIl9rhMYr+7+aogBR4Ryzst4V15nrOcLNVK4QuEKu2Ga9AXQj
2xAB0bbJ/UWtjw0L4A/ZJpipYC0CTXiNGL8MWmjmk9DsBSxCIrGIGgU1RQPqCTMO
meOCJtXgaLPv25vVE7AlZuFaUo4Ao+ZGRnAjvTsrErx1v/u26hdSfXR4/HHDSoWw
fuHltoH1D6KL46ysXH8XZV2szrzCmScY/4skMVGGvRECDpZQuro+8+AcMd2xscdC
L/cpnwvH4o3FjVCcy46j+sT/gcBtI3zYJaQk6U/egd7BIeaFR3OdR8cXuhY8fiI8
gir3crqTlXTr3E5I7Jox6C/l7SC2TvhyXS3z0nhBU1rpGY44pwBf4dtY5aTn9BDT
3rsXEVLAv/0jCVlwBty9evkxa3KULU18022XVNl2T8bnHVEC81ib8YG74sB5jMhj
tTCqS3SV+dAMiH2LaGRZr1rUvBk03aU9rYQQoy5/9i21PQ4BMHGhS9zEhsukC74n
CvUP7XtHMkEdkybcYMAOF4ZDrTl6YHjHVVyMdBzy05ER500eXyPRRKX+aTxNM17t
GE8oV57kFx4kMLh+h98XWtt/3bRGUnopNafvkJt4mapYyt//I3a5C/chGhhuA388
KtCu8fYXF44sxuHHZ8/xSQkKpMS6GXDTLJ8oKdftWLfy2L+MzyBanQDrsagyWKij
IkKYJt01JJaoXwoMGnvfpqtG7Y5p7eJD8WPeVlzAPNH2Qr/ttDlP5ZZ7TdYpqXDo
cDLMoEhyv/j1KBc5675+TD33aS2+0O8Ayg51QaKCPBXUjUeRg8FOqLeHU2fNtsLA
Dc577nOwF7QHCpwga4hBWeYnaQOAK0hAFtgiov36/ja8oKfBrRh7sM7OrBtsWoAS
SUCrggXtL/mASvVZuZyyrGzRy6894FdAvmeCJQ1jLq++NIAXSl3RbPcwaHEJgfr3
bC1NoGcwDA8hL5EKLPndfv8xvKAL6QEa8bo7uHS6v4frIxUdn+FL7/frxjpbwkGC
GD6VezfjvoSNH7Cxla72/GRsQi0IqZ0oI9pTSKUq1lc4hgJJvqIg8j8G1bpA+3wK
ev1FeH/BI0oENNMQ8n9BEO+bqwHMHqS/nfm69C487BZ2ojz36vCaneMwLfIS5LP3
C4Tk4UwB9tNuc/9bkVVqsVm8Ynzm6Ogb7E3o4XOBHz1BrKO7Qium0B+7NWkADiwj
i/b1t82vA4/4F94GSQWu+st9nkdNEN7BJALhyuOxLg31al3f+w//62cLo286k265
3SiFNYSs3fp8keFmJUC8nMoj0DkD20Jzjal7tWMOptfC4Qr7WTY7S+C1KFv6BY9L
/0FvzCndXdouim0ZZNRZdSAb9Q3Jds4zPgXjzM7wY7OXgUShcBexuqH+MG64vu8b
3TbJz9f6X/YBNh2W6tznzlLfQszgoGkSKPnoRcSUulvbMqpwnm8yix9U20CmgQny
aH4xpZf3hjJEW7S7JWmIoViX21YBVOhqhR7R2ePtJV5zT6FSZIxPr9ZW2DBzgUWq
9V0lDTwu1xElGmGFqaQ3cLToaE4lWZ3budf4a6ZSJAd4sqt7eadCF0VsXHcyxIXx
xjUehGOceWq3LPo5cCXvfpsMdBlDRIn3L+vJe/uqGHfetxtlhVPaAr9fWpgbwMO5
YnEw0y44haSvU/fnKWTwdx4yWLKBVuM2Gj6whF4+7nGq955rE5BQc65P0yeIBSuv
dmuGvYhGF9qFPrzP3u9HDrGH0Sgt7nAeDZ19boGyVcv4iRikB9HpLLjdnqSqPtP/
qlkQv7g3wlYIWB6qHvDl4M+B+u1USUk1D/5UxvAvEdr9OUrmXVBEZrDcwCH+oEIk
BgmZN1ehHpYEA5qcm7Swq1aSCE8LumunMHQeKbaCvO6PxdRi8ZhnNONUQamRc6pe
vFFfv8U/HypO93s3e4DigDpcOkAh8gHMb7CR/OxqHowg0IYLbothB3StIb3iBwwp
s6IymbblPn345Hdg9dja6Zi7nN2BPZizV7vSA/Z1A7033F8PWpAEmcbgkyVM29pV
3/HrMXtHYDB9h9nkIQLzNP/dOe69iBmHUtCx8OmThlBoJhQMPninsvDvbbz5wOmd
H0qZdiuI71hVBit467xORs3SqBWloRMyUSxktYUEUUufjpQ+dTyhSY+3NhogJfRC
UPtsj522wepldjSAKrH1eDkHdTDsTjtpRWZ7OJpfkjgNgDuksHT4h+C1R0y/l7kH
97OWv7bVo0aSuRFXok83yCdLvPRaOo4S01fzJsOqL7gLPXhSud2KQWlei9efe+Ab
oPmKMCLRjqNhExkUds0wYJnX11vMFLNbPRX6DFWAKKGjDs2OA3cwVrY3LxYWZaDN
2J8OZh6XGcRP2/Tp/qs3WXWJMWlrNgckk6zNdOaLYBqyGFDtSGmDYhn/om17zW0j
0K3ULwvkfrh9ARpHmo1DmXE6L24OOGK4pX9DBxLJ3TmAoiRDTpbqgcDhZ6gkuJf4
5yjOfODFEBRGCs3VLeVmOMc2pheR8DZy1tljtnGMj049QJs6NImXywHBpuB7SIAz
dfYFNnmVLb8v3eB9/Ml7ptaQTFQuy/3U7p9cUJnnV9qFV3INEnv14iVXadbEoenH
G1ItaWzIqc4GjS1sL4o+2zbfxJj7r9coQA3V3hpd+0qPAk4q5jy2IFVxbY87X6/5
ojgehIdro/7cglUTCNhvczT/7iMhY07hD74BNLsOOaYZ/J7lbGGJWCUDIAOP6nCk
7K4BJgzxzI+jAQG+sMljYREQoC/SuClECOzVzD4ZSm6oBByAqADgFNLSBOiUe6UG
hx5nzAPgVM6wPXI11bFsWkWTphy6RXb6w8Eduw1+o+Uvd/IHp0t0sHYSAU81Gg6T
DpnqW6nZymYgsypJ0d1Y0JakMOq3ExvJ7/Bt3aUe4JvjdBSiP8aa7M6fLOZ+CDIX
hpjsqDhlyMt1ujXnsv1hlfDtuTwcF3f9dOAnny4qy2VYqhEqg8idKN9s07DeEQi0
y9N4GKmq7PlM1RswrKy09PjrecLRR9jCY1KpQgWagZ5/TzNU/gcvJ9uxavUGeAh7
o2hoq9KownFBlbQ+EpxK1HBpAmNuTUm74zu77V5q8tN3pqbbzT6QD3Su/moxTg7z
Ngta9eiw1zh9yZXUyErcFFB3hgUzeK2Vljahdv4cfK53tQA5pubf/wAcSHw6RiLt
93f1iVcNrMG06sF4GhCoMIzHU4DjDATxeMSkC2HnKq1fEJhNdEyxdlwbi4L9AAOO
l/WGKG+5dtnqxftyNzL5BW3UPRG9hTJvAXrJNcII2z9b+SR8/UsUjb68Ghfb72QO
q6USr3+nb4eKXOf4P7qSlOL4m5dXYhp4m9oZGlTw407CQgeRRBNccvvyaxdj/pDi
ykcPKcVT5XXTwM+XXUXKdUbgFmnq8JvfRzgRe0SsLwwtzqe/l+YLkX82ue5STPHE
iY3oiAbnz0osHYmZV3xNbCgNmesWQTXNedV6CG8AkMa4dLZES5jrqtguWYWc7Rn5
9jZxBK/v6ZXHDBgH1ijltAX8b0pJhiWXrQMJVmRwwcfMaOSnblrzrN3YKwJ/XJcd
ILSf6a8SjmuynF2TZ9JGZlE3/wl3tcIqpg/0CHhomcjtkyLEGWZvcvX5RQTF2yq0
7Evu7qk7ljX3+e/bnmYB72mmwlzVE8Nw4sbV9KZA/d+FPZgTSZMoKaytgxB5RhOB
KOMrq06yHMwKT6d3CIv5gBrp5kiOCbuOheDq8yDB/YcQrqrDfJ4Z9tLGDzMHBxUh
52We07nRzM0hM/dhnW+aXWzulsfCKw++5psBZjZyX+QbjjcSy3wjyh/MT1RhFmZ2
8Rz8ohLkqjD4zKWJDijBqzzkLk4HZ/ZOPMRQOjl6/y4UrZyIc7DvoMbZ2XmZhfVJ
yZ/lVCb23FhpaXbxByG9f8+EH1EyMfgNX/G8GlXgUA3M7m7Sim3kM2rpdjW2Cmfw
zdZZY50CrAKbR4x3Tvd5bkdZZCqxREsUAconoYaBRvno25uDZ37FLOVucI890d3J
xsETobShHDite9giNEdWsiMEoX7ftlM9/EyJjZ5UMt6JvpEPvp14tAVgONEGHgsC
kQKAmevuSlwlVk3ctJZ/a03/lgmco6LRpzN6srqrBytWxEghflZj6OXAZn/t4NiA
zx3+y6ezd6kPXFxtIrJhw77izgtqMbPe5+h1c2WWj2vMJKDu4M9YbAP/ko78jcIf
y38yw3DUR6WgpLSBT12r4+KsmknUxMWwRKunVznYHBgRBOsZdzRVLYP1ngHoy7Dr
a5UuGicFRRR/knvgOF5uZDVed+cqJz5JucVC62q4hEwzASz7aHtspUNRksBU1gCC
ODtkznf/pn5YusAWwPzhGIwT3Fzi0GJB6Y/27tqfSsAK3R6qaTfIEwOe9C+17l4X
7E6wtAGJI3kpUtEN46hloB/VdMmaSRN/suik+edUktizHdynn9LLP/OLRvZJO7XE
UfcV6hmkEJEftSBVIM9F11zzU9EfjIRQMyDHj17/RBPAtsopX1oNMpIYAV/kaP+k
Qq2jd1UFzS4nBBUXpEfnS4kN++GLPA38bA6vZh37gdBk7Uvt5D+UlCwSjc0b/83L
Qll+eHi3t2brtTrmXNNf9+ztswHcmM4VhPzspTunPFXbzbSuqJ1wD9Flv4QZ09Pd
0+tdYftYb6EmyVd27XdNclhqnq2Pde1ilZkC3TQ5CV/QX7ZhzN6PpTQNMxVFP31c
aluXWx1nBxK95ywuaSUuU7eoT7xOMnUlFEobmFUDt4Bk5IuQ3oF93ytNPV3w/3BZ
q7fFUb/93OziCHof3IYGLZj9H74hJKIiPVMiGXWORO5kDqCuE68LRNvnWej4RC+C
AY9e2xniOrlexLYGLuszqfYstN2ZA7hbCu7/EIUjx4ZVbHKmvk+cfgxb4JRjcOw8
J3FjMtWLrD9fyEqA+tk0uANbce54K2WB5Ik8ddRHNpdUiUVASFYkktqoJPkVJc30
olqk1qHcyUZ0hLY9bqRU+Ss7jly7UPe26M9mMMMLVTh13NHBdPDve9PYpOGKAg2g
R5atBVT7/FqFZNadk68z7UfxwB6NiI9dj3jX/Xk27LyEz+OyMwJPc7zfaRZSmEjG
sn7rQr2p68fxZ4FCOq1NZGOnaOA9e5pwR23VOgzzNLuxpqf3Y6O9mkvvcIb9bE85
J6Mu27Gu6sbHRARTP38uFLo+dYV761jdgXbqH5sQgToPR4fHlzFqiVtTqw0xcw8Q
VdgYxVOQr2AHXAm17MZwtYvBIx9wApvHlmYSuT5HEg1UOdXxzwdIYrixid8pOSmr
wsh2z9pikwKWlD+dfSDnmCgwPgQuxQezK8ZfH8Fwge+obNHgy2yMmJaK7wdEpD+0
3tvleayRK0BHdO7CWY5fqzd3JzPe5SZkofxalDWSU0KIYxno7w1/7th5rypLTHrW
ENY8X12VlmB7QTvK3krj1BydWqyQQWAL2RDYERaT2KA+1YwlUTa/4q2bJCvQSkef
SD71/PTfAwdv7D9Qe+kX60l160WpqJO78YPSXFsjQt2GA2NxaJJJ25CeUQVuZ+lW
7X6G/QT7/k1ODAcVeL+VRjWrYiL+nLt1ahTLENT3T1KFazTjoHi/CwsYpRFfR9mm
iCyTdHSAQKl07eTSGsZK+6vYCcm00xBSG++nzydUWixu0b4m7yStGWfLYZnfxaeH
HYXzmTuCElW5w1jy8tXWxZ+vUev5x6FUqEiu69ersedvy465sTpeiB/kQHmGb4zH
/rLet8LxstFfOZ2THFjt+jAAteqXpeVCG9u279XFWx4BqjTIJCv9ZdpUYJtA8pho
PKKEzEGieDihMQrArGNfYGgtp/IgqVb+y33UcL0IamDtb/MAdKysx5K4c72XoMW+
qsiGpFiLeQCkUEZlayT+bQrK7lXKzuG8hMY3FhKH7E7dYaS1xFmKIuR58wp9SJcQ
7fwnoY1ThzrdQcjlbjSXZzFgoO+yHrNWhET0xPhEInD82kFYu7VZqM71cRgcUMEc
ytXFRItnVwjImGwE7IVVuZHf8Aeuo8pRi0rK91Ww+kXvBpdFhDYx9xiXLWeqm3X4
8PeERh90IQ+wA073I1Mo6ak9D63AS41AColP6C8yy8VojvqF9Djls8zCYzrAza3K
1iMcKx18i90M5b38RTZApaeDJ5V96OyEu29Xcj94xT5mevr/ym0ufZ77NiitJX7b
vnRjm0Bihyp1SPt3ovCRBBW5Ft6aaru2CPYRNlHiPhAxszVXmpJ28oxPBj3YR+0Y
8O122KsaigavIJb4fsxC53YSNlPokUTNi1oer5iC0O4vHVHJnRMBPe8X1jz0zguu
xljJ/1pBpUQl/I4ihiVSWZqQOaFi84AEToAZ3hwOjYVYoiGHxTgDvdXohJBdKRaZ
WXQKDhw2WBnNDuTyhB/wTfTbQJ620rEz3uByR0HqQYcLVdR5mQD0SbeE6cMyfJXT
jm13T93N4rInaICGKybzJaQ2YCl01+SbcN6amysrI8EWOUgl2MRJmjlkKAqdMkZN
cCeEz3vCajAW/+GfxSfaUYNOS2AuzPBYJdo7v0ASgtu1X2/RBDKl1nSosKnaD/qA
K4Q7jMfAYlv0NNVRqoCgDVi8rEykkroVcTPCQ5A7MByP9ct2ea6KiWWRSnBsP1tX
D8wHN57fL/Hw6JI5UHF7BXkBrnHalymiCXmok85QW3LEy9SUCF9gbhu/g/rC73RH
j027xSQvmKDD2oPB3AiNmxt9i+mP0ffL+uqEqIeK8nf8dUx53GZ87H5I37jQ19BB
MXYRyUQJ5EDjod8fkUfmGe9Gs2wwWoaHft9QiqwvrBV0u97WGq8r3oRtkRjNGqKn
6IBbNrJe/RgkpF03FJb+ZTEb9pKnsZ6DQPAaC6DDocTh8+14AB9pyXDqBiMW5ZI5
Fmx94UiCJUr142XE2BxMKw65iYZdaD2zJOtNP9mLIkhpsLgqxQk0ERnXkVGCIYCM
GuN+10I+daM7ulEkNL8nHlnRvX4fVdlWoHBd6bf/dCHndlRGmeGgK7N9uVQfd6uV
rTwLLdXQrdNz3kWbKWS2Vii/XK91f6qWtRb7wcac8T1jy3NNVnDJwasJexqhtkeN
McNZbhAqAYVlAbBD8gLE/7Sm3MxAahL2Ig2HruaUaojI+q+12jy4gBvjCgglOzyv
VzkLk7btS4KT8VGKL1tbRywXDIu/5gOjkhaZf8hUvvHqNE0vTbIusn1VDae1r+tz
arf5ymdKiHTVojD515m1OWq3zLqHPNiq1vbRzWetr/9yOx1WqTBvMeNt/Y6ioz6K
WerRl3/xuEJVgWf4hP94ZvbGnEc8ML+i9r4emSEoeK/BEY2hPzlQH9MSensTieg5
HYeX1S2Gxnr0qGYqCjcQXQTmDl2mh7Ctol2c041ojfl9kpU1RHO1nAvBUO4Kgvyz
NQypnRSnCmAEcQrt9eKmqG3wTGR9vapCrgxrTf2X7RR6R41FSI7S4F8phUuY9N+n
Ig/H27Efm9LJuNwinCepl8JmGkK4EVZyDYICJ7bMiXKc8Uw1u+EmAWGV8GL5C8Bw
tnVw8QuTvURBGUf3HOPAGSVczpbx7136HVL7ohpraTXKFWKQwpE/tDdeOivp6D1w
JPBR+U//O9UQm/CRQHluD0sSlQfxeIAEzSsFCSY5VioSqCfk/g3BBsPEUfgq1TKZ
XudIC/c+0sqjJTtRagvLMR+vjN3/h24WxeEErhN2aMG8uarX0cjmW77am0eUIb5q
A9WdN5leUKTZV4iojbXWJSykmyM2aDhXfhxbwoav6QnCVxglyjCpy2Gni9IVG+HR
nOBT+LnUJldLeGrxAXWdsCoYInNHdnq0s3GIBXvmCD5g475cfjHKLtpVha8utO7A
6Mm0kdolM85W3Pyqaofn//6szaN7WZv42ETcTzqjMJg4HWsRrpDd41O6GV3gX9l0
qCEDp4SY+YR9Sflbon5A6ADEuvc+HuBt7RXLFLTOz2VKElkDbQJan1hoUBTWGG5T
VjZ2Y+NoAj4ZwSV4RMYB2ZRdYhUudZ4tZdB4Ecu7IkEvuAjqfn3weSxkUFW8aOTm
TvPSeU2mrFsKQr7cN7MuQIJG8AquXvwR4VP0vowJ6RnEZmT7OTegBmalzy1X/GAc
pwUvedgPUyKNSuB8lQuoc5G9mbSZzEOBVb4ZedhPszR8jy+LKGP73SRLqxWKXqa6
hVgjv9mbC8uB19Dah6us3A6cXJ3ftWfpYQK0kbc+ae5GU8L2MNO+96+HPzCc8yvF
z8fUsiQ6DOASCA03I5nz4vY3MybaNI7Q/fAss1MzNp6d3fZsweGi5RzFulC842QK
e0F8FDGqyC9x52ogtBn31dFYLymUMcKZ7v77a7QUxuHXvHBfNSqRNMDQ23fZrgeP
s+IIU4Qo3aKY6RjSsT8LM+d0r43kblSTJEcMp4FJPg2AsAnjjg33/7/ICFgIhF4q
Goy+2I2ByoFYaea77VTl+SR46UMxFCsLd5SEtn+7o3V0UFXlXEpvAGiTOV8NY9H/
4ltYhvUMYsk5DDuvTab3r0nBs+l0jn0nsAaV84xIp6JMweG0eyuSZYxjIcyd1C87
0wxkbrSVGxHGzZPRXqhHGjGMsCih4zPhYLl+DZeLGKTjFVb6/CPdjcc/NO8sPTaX
/Aib06L649V8ZcZ0Pq4taOvcniFbi0bNvq9rXinknrpDCXk4Pi4ewxb5oZSmQWcs
cTslBEY/LlMxu6oGcH9viss+rjQsmlUTj7qy4MZvTqYXOcpl1yg5AVwr843A027d
GJT+kM3z8AUHtVytWHkB+8896OOK0uA7TIYOI+VBojg/ETJpTA9UVLGxh3dgTBEJ
s2YoYH4mc65JgKCTVY9sJV3SRLcKY2qe+oDLpVnoFClKFnAMfLIxpLEDyhS9J/7u
mgmqX7MXDAwuHExIe4PBXh1b4z4UdTPoo/Mz061f4QJ4U4EFnWLjYewnS+WeMdGi
yBBB5l2m/l4WkzB9VHlLXgwbt7lY+UMUqdCjESNNt6b/mQaxukcjjtbMw8DDFDTC
k21WGBjxmQ8xMBpPiikk7FewmSKeIP8SH3VA3Q+23Ce0WA/+4clrJEI/i2j3/x51
isb5zfeDIU/rOZN486zppn9pKPqPlAeTxOo6euf33cJLmj04bVUAQ1qtsYfeSZ5K
XwG8z6i7TxPeGkb/fa7GOOydYWvt9GFQL9SWJwE9X/rvQ50IJUWX5ud6N6M4iJUJ
s1h8WMTi/6S17+XSyMp+k49MhcRjXV+7WZF+ZqvHU4M8tVBIPv9OIcilp7n8cjYC
qMBXs6hUxOWuudlTzjDojvw5Yacj65sX0bFKr4m1l5VhDk4/H2CYIO8TEB3cqSgK
CToFB1IQW+DXTjj2/4OQzYhXfy7UuFkFuOCkr+9zyzltVBQP92sgsk45BQDLAhGr
KgOibXyNekWDqs5EB1RlYvWvhnguAWotV36yTvEZvT3gLGq+q48ZJbYri3kczu/Q
YlFKk9z4q8iW8comQ9mYeoeueUQre0cFzMwxJeyzCPQdxbfuBF5mgkRuVFzroGEV
+AIAkvnXb0ZztvLBe8ljF1jL7nY4prun2/dwcQ6NQTZ0Lozz7dNQn3DAnsQE3ng/
BmOKjhpwBwnWLwCAziiApKZ5PRFu/5z7IpvFIKk64AWCTLg2skXg1bG739NTr4fa
gA/1NcfrIQJDDASNwdz1mo7ItJ0yLNRb5cz3EVMTpD5JtRilzIHMuLOvnhIGaZxx
uNnpX+3PEEedDw/vKPIKMSfi+yp9fe0nhINgqRl07tfK+dhHYdfXrWcvK4CujxXg
Bbjgwo4pt3L3HAJV4nbYOKge7IFEi6qZMgFqyYf9XP+ufIWppcZrBh9W6upNfuE/
n95eiPvRe/6xvqxF+Xv+vuEKu3jFdKXjvrJloNvhciE+EI9GCEuVXz83E0N1tX7A
KreimodJW6BFUGwThHDE7xxZo6oDTAnG4gJYhghICLHJzqT6vQoBCk4N7MiJDcz5
PbSN5CYp5JjqK8R3TKPcaajO5rDhDBAnroHOJB4y9w8+MbOlbkT4G7XG9ZYd63gw
lqUfXrNs02x0ltXid7WsoysHEEy2gyNqjN6Kitc57bUZfjKA5XJiViMoPZeIqLOp
s/3nmWkVq4aAH6ldMBsWMUQDrvzNyaEnMLcYqZeqE5HTPJK80P6TGYkvAcuOb1I6
mzWzvsUOJw5zFX+vFSvGqGfciJGnNNEdlvZ4mBmtprSmPy8YFwck9xjB6mtqHHkj
H8byRwgn1jqPX68TPjNoMuBJrYE6xZ5SLyD6oiZEQU0ufa5GlNuoJk56t3ncXKhB
mfZaIgjGziPbZwtN5ah271sKb+64YtfGwgLf0PSnIOCqH3/mX97FGVELnMiPZeZe
sNpdQ/iBuCs+34NSMDb+AU8X/SxIxEYWjzfB/+HEFY3sQ2G0A3NzNWyNe6jiqGTB
ZVuB8+oW257sbk+rVeSkwfv98pbAg35D1Ea7fJB2nZCkl8Ipen6bTTyb+51SdstC
mlP2hzpqa+oDtDpO1hTwIrMZURYIE3GPAXGJMpejOl0ThUrb9MfsCav9TcNn+vEl
aTtjBLzKGuNjWZcYtA9j7SKz/JHvnu0DisDiqmWPXm+ULqOKyGfj6BWBMl3WAz0h
AMzKB7kLV4D3KwMMBOF/iCtmdRoQ0PBpyjqcZabbOzgA4Y7C+v26tm/kfn0ekhIk
1yGgyc76xxpXa6qVLPFQxBghHI5DBsv2Q1bc5/KmLU4k1uOvD7iBxnLF8K/0yNZ0
8X6t4yzM9ByWxTEvBGVVmZjnO9KhrooXstj0DlfTDnPA+mURST1FayIEIZ4H3DRP
XgbdQ2I8yLqAH4Y4n71uvuH1mYkHkdaXhZDHI2nBiyyN5hwICdqwGn0YLnTj2A+T
Ol03k0RkigpvODFeI39VCwh0JqcFJDt4XPRIe59nnnhOmH54vdy1iQ2Hy1qTUPbi
fFJJh99JWPd4Cg3JTjfytX303xTJvbd7o+q5TmSHAG9Fqs1HxOXrw6p6oxvJ8+8l
jOa45IvjA+Z9uGuMUmiID+Lc482qVJITWdEovGyfvWONtCAyaDxwc+dMhTNPuqfH
NrdOhV2px7YGZC9grrhoWjSdMRbqD8ZSWR0zFXFtqCMRu05Q21JCGRoeZ+V3wjPy
UgpJRqg8E0/qQzE1GYtdm6O0kBGfhA5oXrbPACUZVhyHw1SteyXOMTofa1YTk3sd
8g8cgL/OGIqmi1LA46zBWoH4HQJ7ztk45nKQz0qojwl0RY/WZAshycHQNuDnw483
5aCz+NBG+J1KjgRIpjNNekJjeBWeR3zGYn+yHVAdWhfFvdnoYT3r1Js7IFdUU/TL
QBh710FsU/K0gZnTTi0tQzxhT7aLulZzUKplC+BoVXNWsOVMIOesUrFCULPWGjOP
/jatlL9gVDOUIWrpgM2Q9Nu4bWRUmp9fF13M7dSU6GWgV866WEYjEYa4F2C5ATER
VLSTHIMTrKwNNV0Z/ZRu81zUVvKuUGJAvndwCbPHCWPhEHrJZ5qaAoKHHPG78xCF
erJOqS2T0B9DdudywYBKgyE0v643DqC8CN6rfZ6lUGtVKP/s2GORTGti7MeNXIh+
WMoLN4brfMHZ/GqAQkLnR9Ttr/yBc7xoeoQ3zXB2BeJu0jQtg6WlOQS1L18Qn8a1
XQiGHMO321GbBiRhIqD57cn9xTCP2vj/w8RBff5lY4MHsDdVn+/P9x7xSIheHYf9
1k4WgXpxu/uVr9JguQqzPxH5KETeaBORtIiI5SMwLaSuvg2IeCMBllKd0JWdG/rU
yJtIZ8U5S7Qq0Q/MzT/ar+Sxi9fBx8NCNwIIhXepsgRCu14VoQuZDZZGb2m9NRXm
DhdfQ6MeJ7EnTDzGAiCsNClnD2OPrpleWkUzbT4GcIZ/wzZ3BYcFnq83bEWERwB1
cF/EC3MqK/6AvvWOSW8OnEyoiVPNAOzfUtkIffdfKJOc5pcttfqYNuu1GRXtMGL/
UsIQ+www2UBYiTU+VGFG5IrbSMh+i1ooanSxKrqeFX85qgq4JyH9qwNtDXKldmc3
btJrKcrgcs6fbaJGQKFV0Bvs2HZgieFq0zTp2RGGfXIwt3DhLgNC2zipj060qif9
qNrQoPvIJ8/TXRcpy34bA5YO8WwFG2yw58Y6XXCTM4ARAJqqQ2exJD9H/vp3sJHs
PTb9vENb9/cJwE2TZJCbAskrP/KYeuIEelZsGoLsT6RUFsWGY+Z0kYEJVoD/chL8
hcrW0tj0VIBCH7FIHCtU1iWvRPiP/v/HNvH+UrJNpWi3kb5W+qDPZln6YRmrsmGz
CW+EdDCXfqoU9tgraGQ2uKJiXMUbf5xsSO7NRc3d6PkjKq2DmAOFUZQfJ1dJNU5V
O8vhaMLjNFcriQErJABHhEwonq3C8V5xJHvW8n4A7aQqoIYvRuPFcnBggmx2pcTw
Dlr0Ik1GyqbhUXmMRsBJcPxmoiTxPpjNJx93s+a8MmvQF7hnCmVRQTWrXh9bQibg
zDxU3/yJjbna4fNWCqUqvGkzFZN+el0wFSsNqL1CduNxTAlbcpOgGTFtW34q0P+n
eaXvnOkTjFzrGe31+YlsrjjYuxILZhAoMdrzNkIBqdxr4wEemTBJZWaMU2XmM0By
buQDs4r/1SY6MZMTuq6I7hLX3joI6lGwH+jrHAz30WQ4updyZr9ue+MmfH1tBDpA
FTV9fm8JBCPi8x+pWQC0j2O6/vd4Z6ZJCiJjE8Id+VJGuTJPsihErhmVym8ukK8I
/QrKYiYwg9xaidRoUms92fXQ6oWj7Ko7bCjCdBMZjsaM35mn8xzM6yR4r7CWqBw9
EFu5k5cjGSvY2YW+HvmnWXItREeAShJhkzs+CJ/OsYrbeMoetX1NohPB1BBq+Pqb
GC8BkCnCHQ0iD6h0Y1M+f8xt1mUE1lIcERY6nPwJU7ZNAXPV/N6sqp3KvOZQrJum
UYTZc5P+UY343v2DwKEV9tjoxk9cOau2C4eH8wlF5iJap47z8KGhx4+BMKhiEQUF
HMUuNjPzfgNvcSG78WDoyXzVNWan9eyWjcM59/0Xp3ZZCRSzaGdW0k92WwDd6394
EQR4F00VRo+sV4E77PhhgwHSxWBVD/cj4XotyYF8chjhRJEEA9MBJ2ae8xaPMyxh
pzPnAZOZYgLRxdSXutWfLaI7bjboZGbLWdXCygo9S1Yl73HJGJSidMUirUt8LpQG
8/472CCIi3MIDqYXHTt0rtT/ai7pDuDGK26a96abqpLcn9iqsUH9UW+X3Vn1hTbA
HLkWyEdf5jGqqCbP7506npj7+UwXZ1oyiPeVO5dz4D66R3YPN8pNAVLVVPNf5EU5
MYSZIsT1RHc+hrsoKt+n9e3n2L5WJSm1y9x3/XRiS5ZWyE212OHXcAGl955gGjwd
MOW6B4rdbNTt1L5RSaCgcJiIFKZwmmtYmH8sxQFmDAekh5Y1n7DeYMPTa15a849O
oE2spRjO7M+oCsBiYSJR/DNCkQeqhzYHUyz28Xp6N4Hg4VgbXbrDy72Dnc5pTUK3
D8xVBYa+oP2BMafxihxdjnqJG0HFMF41pbChVFgRV+9wjLP5SpwhWCG+xX3aBFO5
RRUfE9+X0kMjn7tCL+Y0jJ5uxzfXGZZlVK5OKz7V8H8Jvyx+zG6sxNaLTYyEHu+8
1Qt5Zi+UXT+XrvGUT5WAV2438KuY79dUP/Sbqzv5jga5MxQnGIXpTyjUWLRtpeLv
18C4WR5KMXoyyKRwy4hZ9og2oOHYRhub2ko1n76WwJ45P0Ybfpi3iHe8MD/Nl4+l
TgUujBbg1GXNTmoN5ceP/skC8nS3DrrdZ0z+tpiOWPyZ5vP79MnRUlipa9xV6SrI
1VSvjfoXH60fxQ5V7jeXd0HWE2ns8E1wIRR8m7xB7fb/7Actv3tw312esUglqn4S
8mmGLykdGgXQOeL6LPIIiAD8uBC4eg5ROQIoUBXljDaRrv790LBYMG6T3b+4VBVk
X0vCjTZY3HyBYbnZYJHpA7iKqroeAEpwPdeL/aKbQCPd25LdcSb8qOfHfkMa1fhX
NPqUJK7xJSqSIAqfZMu3YLWpkn84rkmU15Uebvwse6qSKo+RfjeRu9qxC0xxXbxI
wMo2BShJUzFW4ZXVy0qsF7WfRCd5Ry6SJTL5kwm6ScmkJP9zmr373pMR91jJcDMw
0AzfT/4RvPSQjrpEstIOJb0uHNCwo0OdbgUGe/XyzmEEIDc+PfkqRYK6XO/ygzHi
sIxJbqX8R0961K8gOI4nGyZeJbjihlFQjtCHi31J/SWp3m6ZV0qTuoPVcVpomDl3
m7YRn/Hd1OU1Y4ZscU5WewUQRBpcoF3D/JA6HnI01Fg4Qfsd1q0y8TafN+tzYNb4
28BpmlBQNEYal+ImlkdTvP/rUrAbyR/Dlxb8l8Dv1FAfM+HC/uC87GHydg0nHOex
sKmPiJuMiHqr7i+l20fZ09HU3UV/mY5EWeed/f8wjeuZ0S5i/4bQQn3b6vtKccn3
wSSZPXEEm+TVpRVS1E9szZSAq85hghaStoa/2+AFgCH4xHMFV/hSzLa1iQZfTSEN
okiGECJsjx3D+gcB/GMB56XPkBSXff1xSbTq3H1CNFNak1hMvcioWvoQ2kPp/E5j
A0CNcz5qeJG+AF/FtIlImjJuqOvV6c56YBHwx65SHFEj0ymIivcyD0Jenl1tTGY8
HzLhmrMPRldfjwuliNyq68kQAxtEuDO5kJ1q+9f3SHQ/2Y4rLNOnSQIje2/kdH8X
+kGjmQLyzI9cXdpRHOQ1dWvKwEciFrWJ+nnGdscBH32PN6ZW/fsGNtGagXGjIojW
iECcWS7nGCi+BIndpH3qFajB7j5wd4xPEvIyQ0teka28Z4xSJOAdXhqLoL28XTQQ
de/SGuvGxj4pbgEnNfkSMxq8H2TUZeawl+6YwbS6cDg0NVnKJLbOjd8WvmDW+I/S
DG92RotYqqS4RoSDs1ey24P6Z2DtXc/tXSLmzpNFExoeQx+mCgiQuNwkvZdW5uz9
80UFUFaOGNTPagOCET9W0IzI4Io+M9XlIXp3BmRt8RVQN7Sf6N6vZNPcwk9BOrqW
D4Hn29CzQl1sdbadvqxWeqTvtHwlmjGd2NTNnNVT7OXKvCw4xgpMMdMQm/iLesPo
bGQXK/yI/+98rJNs18kfqpk1NLIRta0/zzEuztWUw6U2V72pJdyy/qHV852VPH7E
PRVsxEJSVagMkhzU9Lm2GEGWzM44fsj87+uyPswTLWa4zhbLbSeWStGlrB8PQWW2
ACLACSNEi2Z+uUzpHaA7b7E4A/9T+cNngLNra/12t4/KwGyogRjG9sTNsAMAbeUf
H9mV67WZ1cKyEfg6l9KYzfwhcBIpfG53bwvaa+sMN8MLqbKUsyLHmADH9FYYkQVT
wx4nAx7oxaoKBJp3F6D/MEjgI2X9MqA5cTixb0nbAVfvMEDLH8H3uCPRA9ysmuMp
k1LEQL0KmXcqrkNmwC4Qa+q5+1Q5QMbtt2GP+D5jDc1h7jgKlX/glWHKiYgF5s+H
EynnIBbF5d7pJ2ddqCBYatTUCzjuj0zB3bqZpJTyMCA4eCWZ1xzDqX/laXmg2pAL
1oPU5p9PehZ4g36zViKtD5bPMmDgoaCOPTpESiozzYeV/5POejR/e/stNphuQsco
mglqZ/l2V3YYFP31qOECEK5LDz7sPeo54tHIqrcKWm6IpYrqYiJiyYrM/FuHhNWy
IwWNNrZ5tQZkTh1E87JcFgVb4C//RqhJ9C/MggiLoTS53yVvsCPBYr+WWbdQEIKa
3lYdqHb28tMj7P+TEWdO9W5DFXP7lVh+VZo2uemYyHDjpOmrBQg3lxk7Ocpu535e
yCMWC2+aUqgCcp3FmOIweteVSvamRH5+mVseb5BZxAmzZ84ekm7CRXCJLScLiIQS
j/1BhVIWUFRWQEcr4JDC430bw0yFTdezST50rYWV3X3q/q+JHDuyXnS5QAQHyqHR
I4OdTL02sN50CU+9HJ0tZDxJOJ+Kro/sS+frmpIA8qA8NuadQs3aPR/G2k+hoCU1
kX8fcFUumloNvoH20/yR/D/QVE4GMOOqH6vEgTw7a05K02Ycl+n3bIrN74bP9tNE
//9RV4r0gQkF+alOoUU2TDBLpVPMSRlDWTQKmfm2581zEHZlPTyu+B5ifLHUV7+f
GxKmzJW6wFK/GMeNBGGACdZRz5dwSiuOkAV6UHuk42/Oc2KgLFhUtFxtKypm2lBn
7c22N8h1uY62OT5KK+eg3Gl+sZKZ3+HApwTwOkpVbexkSHn+eNzmeuNzdjCInvly
tovTogRHVLOTud6646pBu6FqGmP0fR7zQaYs2jywzQYu3hkrc8fkmf0fLZ96OAs8
Jj67/oUICmT+vbVsQ2jRrJSgfH9lMqrf5fKFZU4DshDp+6C+K08o02prPuM/zas3
ZDL17XGrQ6mWb73dlv45prSMQZNZtL2Vhr5CK5npQ6uO/W1wOzowloLo5A/2ciE8
VqCsmN12IgDs/+tdnFWYxM3GWYxBtafJJOPD9zmGmuNe9Jg2GxXfqSJI/1HNEykg
0R34RZuRfO/UZXM4mv3BChqK7/WzweVkoZvGr0IrSXsmts83JpOMYk2j8oT2Ch37
9iJ/K/mlIySH+nME/xpN7xoIMWCy3EGmvB33QeXk6hfsbPjeOegjopDVulsvB/fL
6D6T53d0+Wi4ktBU15SHPPeeTYWMOOrDZn/HoRPKF6oUhXQaJB1a+qb8QzQScRHs
EuyL9OEsxJwnhHF4M8SdDR2FBgj2WsAfqjVS9nXTt+A+8sHCg+Wao0PTOfk0fdc6
rGkjYR1XlO43X62qMAtWe25K75h6QtNNKnd70jJ9V704AFomRGgG5k03d8yFbDeF
2DpiQ/2ELkdJPKhnmo4vWExbDvoIobRSQMq2aeJFe3DNyJOyXs0a6QEHfF0M/vuQ
/u27OxX6owM6jXJSd2B651Lfm06F1pzaDrGFplsbx8wfhZ7d6zTs4TNf9mDrabAE
R+iS+6XZx6lwtcQvlmJwH4mnOU2g7w9r8Uses8bRSh73KTx249VnfcvYmt9dYOln
O2JdzFp8Mrjs7KmF4B0GK11JMhR7E8bPIbhkv7Lg+Xx3K2m/8utz+RLOsDr+JuLT
GQ0UoGunKYloVB0av7qfR5Ex3XfnUoRGLa0KdJUszFvXxTfbAQ/YHGQEuap7hhGe
28mZpF1JYd1z3ErrFiDZ5q9W+Dqf4o9na1JAURfJRN61+CpnP82f+t7NIGuv97BO
5yGxRHCXqUO7DqCLtPSalzRFsAkM6gUti2kPDw0gf2ZXsMW4ElUkTYxq7KEzJN2I
oXwD6cvulqrpSJK0wOnPS2lf/tHEmXPdvIotJTR99fDpt/h/fBm2NevQve1HeLA4
nHfY9JSUNsREsWUwOco2WVbA+stiFF8rt8O/FYIuiFgd/Ocj6S9A20OThMGtFV/c
eCYL+aMjnfFU37fisrO39NoSRzUaN7U3C93Rw1AOu3cHT9VedQpZdz5P/3Go/S8L
skWvUKo55AjXMlM6i4P6YmyNSgKN8dulgziPmrx0/D9nP+FMvXGi9HGETDhckqp2
tgoWtwx6aIDJXi0BeQSEqbK8nF+0qyEgLR6NBgYlHOpYRMp9GcH+YsQ9/b3dhMKk
tRY5DqODXhmxu7ezew9Mr0x/Qmt8A9z3Oc8rFoD5PatjpQGBr8Ktwt9zrGQTCIrQ
scbbrzqnBVrh41IRonlLvJkp+Z5iP+n0SIf4G80R+BW4Cap08EmbpP/Idld05zf+
o5MRT5/dI3Zz9lWT/6HyCFqxDTBKQtaFxSjz/vilq0r+kVGDKCaFhqsZXT8C7seu
CwoDPd31iFawKYrj0PkliYWbLcDT9MLdYPvvGTqz70HdwDB3bXbqa0/e/cl9bQ8c
BhUeuCYE/WGiwLS62/paBFNvu4puvAQt0SeAaJ8ZPvMYRs4XtrvKtxmjtSpbAXdC
lP5dQWkSKCPoG8JigaNjMFaZMob4P8SVTM4Oa8+poGE1O2NIV1Ebi8z3Zgp5atNh
uHPEqsExxtn9cDbn4LktjaGae+CmLP4P+cdIhP+m9MWVX7dp/D0jeFE870IFdGfp
ieRFzhMQVylhJ/xB8YF0ZQFerD3NjjuGIWZ3RmeUp0JbWrUgFh4+VeLP8nOVIEim
01iZf0WIMKN+OshW4iAvP4w7JmiRTKYWxC4vBkqmOjJgKIlCJR67FxMRZ66FTcvE
WYJZgWkwc7anh2i78EBnmL+V6dQe4VERM8rffktAZgIkl+YVIYnOCMx20BnfaUkq
MT3t4034WIT8uVzhdgP9x/LcrMFkunk2rMdfAwbOJ/HN8bfs4xe3hvn66QcU8Gy2
HrXSIpNJDlnI4C/bdEU1IMLV2YII2xBVB8aIaC9IzFGvSPYU0MEAdYqJ0vgfSdGO
VerKufUzl0ErnAuL//0/CmuaJ8yo/GI9gayUrjQS/ePfRW8s3G4TwKSTqZB7yOdn
dqHWBb9L6A6ZA++1q9A7nvzThh2YxYrvfYit9vA0e2NTY8wIqNxhBRdt76yYAo/B
OZU6OaJGHJUoSBhw/R7O1JxZqjQs2TI5WZZsBHSx/aXsHYlSjN8pUstkm6CaXvWN
LyyWwRWRw0htGJkFhAwDSjZz3vbOXCM5k3AXcDYqimXEZdRbpUJCi1sIYQgGlo6/
J5oISu8uoGIMdLv3C8duvaYDxxin6jlZPjt4NDwS1IlzFu9p9KEPJfB7tO7W8DEO
GIF7Hqgr2VhFu+OtwrJSjIeQ+vgwJ4952vCJhfz6rKInnf/5ET+48ZpOTFYru2BQ
TOkBxDqBG+P8/sglqtp9VXiXyDwI/77CLV+6P/HutgVk7h6HO0lJ5ABGy6l4mUbi
lzGC8I25pdSX8H1vD+kZ4YQXGJA1Cgt/6omzzoS/Vje+m0Rk/jQRd6C1cNcdtsiM
oua4k0UE6l01b7j5t/zsLNTU+kGkIJdySuWvE+VfOyVS+dnEfsb+LdlX5N9AEtto
sNeI5v+IWYDT1CLRXAB/xutpL5aoBzG3lGSVa67tEKMyJCqc+cTZwwoRchdPIzRJ
+4NCtHL/3iXMT8OWVYyaomAAwXO4ZieCuZDClVW/z1lfesz09Tg+fFJOMbap7/JC
9549TL3zo+w22CYhXqtww2K5pKP1k5K5aN+0PsLbo1iGYm1z0FhLBrBWIb3NZqeU
CoLLpsQc9Yfmt86y59r04irbNLdJYYfGO/VCxoRU5p59y/s/v/hnZXnbz/GAK/cv
ACnTkPJWC0PXoudypk2yBVKThcX7VCLG6nqXCWudFd8OgGcqlcSwkyCroC5CmcFZ
1Zf95pcutlQoeturLNBIH8HXQXZNQNxdMz+7QXx7nRbWzcUHamWRdnK80+0Jejk/
DGGXm2LbZIK9TTDZ8NHyEp2ePJKS8K+WxLscEgxIb6KXXyeCzRbXJK/Ja6xpHq3l
Jrx6/xz2pVRgWWdmh0Nv9nJDf+pmjDWgPPKfNyudoV75CV8Zyjtm+WFd40z6vN2u
Bg8IbUEUVJx2IBIKk+qBBnGFxEkqCGtI0UXv3yReg3YvAxKqdmZvlvOuMLj1BoMN
jY6lK6utL+IGe+xMrc2t8gbiBBIe48Zv9b6WxeuU7RFth28hHEcIwBJOwz4xz0jJ
tmOYEf/7PZzB+aUmvUushnGR/zptjpOgleppQ65SPlJ9y6kQxM1z0sYM89yV2EG+
HQpiu85+QjCcKnujrYXibdEGEpvzB4eD1EkUffo+hHyZMlEe7jBumYntKR9kvqXc
S22i/TafW0CUvKfizQFCzCAycrs47ug9jVBc7EcXJc9wUuztS4h1Q8+HdlKFvpbP
h5OgBFQpfywupEueqeJIPZ/JiFMRc7D0kW7CxqxocNSCblyS0/06XFxRFvCrWlJR
W1TJV8ShJE6r/r7iy7y8Rg580xhsVqPfDtvzLmTkh6MPtaKdWHzXDdWM7GShDXFP
9v1snQjViRqWIgu5hUYKNUSuNAeNQjGD22JhhQXZhGfOybrGaldPVtelW9KhlVVZ
Avub9rGsHnJ4SQT6hJpVSK3WQ7vPSttb2FjBt+4Jc8qfIiaDMUUk+vOSdMy3y7oB
xoQZ/pL+5fZYlmqbEz/xyTa1fJJzq1VBRoTSLDOr3Ca0T9oRQs5abAe7YFgxCvuc
cmU9CCHlM7s0esEnM5XLbzlFxTCrfax4YLK+XiujpHG8ZOjWdvQeB9d8AJAvVqtg
nhMFJ41xgbwVc1ulT1FQ3WTha0NPqynC2tkWWJXBL0IkX4Bv9X0FeBwpqNVivajv
kdQ+mp16aDKKMOGNLiIfpPFzNY3oYw6ImqQFzCKKyBsOexWQGXNlSdGWBa7EdD5M
ORAMz6mvbFKg1eOMEUsCL3XizMlsZs0tLX7y6MGRo+m/fbXjsShs1UgA9fPXDdT8
+t+SnZF+hWofjOOc8lQWtwBjq/5AEVPEpzTqWd77KY9nXZqHMc6p7lY+y68KrhDg
wddkvqTrXXTTxY2b0cjD8o0l7nKvc9Tjqz0HzOo6AmEmk5I87AKNP65dszDxJIK2
Yvq5yrRRA7kKN0DWJA9hhNOfi8x5VEoOgS3NiTLILnggmms04WObIVvaNzS8lsjR
2oFBUPM/RXvlxZT2pS377KtH3QiDOb2EdH5lOs/XFZZYmlQS5CtoFGjh1nNofWm8
YozeHDCtw6IDN10jxvE1qXbwrlWyEUmIWfPvvXOkUAfUChL50iHaAgWe17aPErIC
wIid+txo5BN5bfxQQcGNztiUiZfKYDY3IukYX5fuMm9pPB1D828hjlJ4mlkDmp8P
MqTja46OK9aBSPN5pFhwAtA0S6TW4phPKE4HbtHlrpiQM8RDPBKVcBBuyj0xSb48
RGGJIpuUOoEfT0jklKJJJmg+/L0dRPsrKdV6T3YQmAQGfQWKSXTkYP54kTCOstSr
JItIVmrRyTKBAgYgGv1T/F65rbcQ60eM0GqnsVq+2T0tpytlyp13GzhncKqschQX
Q5CaQ2I9QoH33alQt/ilD92ji7s9+Uli3uB/0uzAXA+yCIxDxP2JVsQkDhCFGaqr
KyXatXjtKbyr6Z5/tqGqpNm8Smudxa7Rl3Mf4cECCnhs0vD5XY93z+ViTWd289N1
MoxS6BlAG8KVq/Taa8fG5y7ZXIgwD7bL+f/qEIHYq0bS/wR1goxHjpAEtGq8whCq
Ec+mEaOB5PHUYGwvsns/pc0AtaaDmg1Yu6+Lh4+PEgyjo/v1Q5LS4lUiK4mLD2tB
2yFwFkxUl7lKkErsXTf+hr88q9BU+LJfGreDmTvpe1NP2SPyWWnGtdKFWYAwz+5I
HAu2f7H4xyetHAAv5jUBcylESaYc1tcoHGjn/D1ahwmWnBfJz4bAeeRd0p09qvAt
EnPt6mIOOKK5Fo2sRc46v2HwNooAWhibcp5Ai7OusLn53tdw0g1qIVwGTMNbJtu1
BzwDYEk1WeYyBcwm4Kk3YhPe/7CCzsDmkzVpTzI19rY4gv+Cjj7Y7GkNCn89+M2T
O/tGUqrM1QnDjm90frnJ3TcsVR2LpxMQK1pIeFTqXARD1wiTQBrhDk1PDud3vyom
MfYNmaN14aH2SYZt+CKISbkRdEIm6lurKxjzRQrI1Scp7YcmN7aTinpgQ+lACfSd
iEIx8hmjUqvHx75qlj4BYLBogDLs1QSyJhiM5PoK0zwZwy6kXdI+Jm/XJShi/elN
gBssgw112xJAF8CtxtRQX0vJH0ItEzrterxJ5lJUfqz9tJn0+lNS9t9dQ/Ek/KTL
RkB6EqM2Ere/SZaEABGPGjW11r+SbQilT0qKiRu/abYuX+KXPkIQBvcnLcSj6Bai
KI0Y4np9XKfAE+zsC4r7I5rE1u4p/0d63ScPsbrLr8IG21ltEGSxQGoBUUc3HfPK
hyHboNRxwJ9Gx41ohh3eTVnCkakwJ6v2GmMR+zVYx6NAJViSs26GSNc7WwbTrZ13
eyGhgrMXAipHwj3dnrR+WK04nIjv1f4tSVbEG7U1RwXdyDrB6rDsXC8bt0DcDG8F
BIYKN9rfjq6Al1YlP3uzUFPFuV8Cyzcp6+M6BWyft21zIlCzELpo2bIs6P8nLknj
cqJBnoV80ZuvzRgDH3bwkIWF4XRWGPnnPl6OazFiAnwY4RMvnrwroMPAIBncSyln
OnIa6WnI5635K2LiD7nAnaeLVskR0Bgx67+RJtGvY/12gq0Cge0Gyi480QqXOzLw
2pJaLZErx0MgWSWkUB+PryAjwnlsecLLi8olKYmkxyTpdP2rLB/q2dqAiacS7eTH
Qz1gD7J2WxLcmjEVcst7Qhwk6q7SYdiOisJok9cLt4FrDGji7g8SPaLwbOhITF2A
nEKBTMfVyUkJxDBxgk/JAo1w6JE0Jv0Ae84pWAlZg0kPPaEaKEz5iuwa7lLkTKol
dBD63eR4c7er/LyeKHEIHSE09dL2BOU8TK8BsbvfoAtoJ+rVcjtDayqV7r6jNaul
klNBfQUZKzvJ/aue0LS4f5K4cVtPqJ9wsFBR/GqVNCT2GwfdtoLk5UEZFByYUDRv
SoXtlJjUvaWOIq4n1locPFGXBNK7lJx2V/qx0Ndp/qVSn59dE3Ow4pQ59uTq3BAg
/y4CUxIoVK3REPmvTZKX5JjHifhwJFUrfDeIiIrZMjJP88Wkb7ex5NFexnXyW7dr
55rvous+2uY6QGQaAFP8to7unyUnwCjU4PDQBqDiIiRxk+MFvNIKWPqQgF6im+Df
4m8FXcj2dZ9xuPpgKejdBJkuRC7mkhcEOZN2kFU8naNU9dMGLGMJLngmlOSO9oRf
M93qLXNATdxkwDsY3tCTTlZS88VU0zncz95PVIF3gZwrTVy8GOwyDar/8GlkG79L
d2Pm9EU1dHQ46+++kIDXddBOpKu5liF4JPU44jvx2cW/wiYJJsm32JClmIRvpu7U
e1RTQF+I6sTlrjOlEDPvsgYYXlojV7JsXUuzWZjPcdhIoKFZ15SLHcq/qeQqxQMo
k4Yvtul+Jl8uC2qIhY+MjiJgilwUKzL+iO2R38EOQSrPnLUxER0pXdh36cu+6dPl
9AC7hnjrCA/H8lMEC0ASnAd4vK028U+ahaMk++24nNYUKpfSihuxONoI4+YF98z/
sMRwaV4QjCAHx+aIp6aW8Uxui1gkzopibN1I3oOvWlOBi7oApAq8q4/rHvKpQjSE
gmhMYNWz67RbB9YhKtPtzr/KmmfcyHl/NU6+Li7QxbbFpEKBx+MiVZnXHeTwu5a5
nvuB+3YJNkjfmMJQ3jYK8qjfHVvOd0ldUXYx9K3l24V7EqoyHxKwjQgWj/YsV+O5
CHajFr9RPMp3A1IOfXxh1s3J8R3z7uJ7xahb6UF2dLzueLlmwsDCZtpbZpBoMOkL
Njx9W5AHCSjdvCGEUtObirMbbktR5T6EJKQhJMr1N9KhCx7zGb8LYXvK5CZ7/6q6
jPODNVc9Ko+QX3X04KOJrqn/AXW10hVwTU1X5lYMO+YDcL79vujLcoURtY4gHAB3
4su5FyEJMiyECkDa9+u3gH2GbCSBMi+U4g66RA6HqVC1d096WOnnUI7sJcH4PXRc
72cYxt8xB2gTd8ytf8dIbCPdCWA7wW2iem30MVyw3DPhOHGOpce2L6bAhPzU5/zZ
yeg7xXj1c6Bch3/hBHidgScE3zaqrKz9ei09D9z/la5T0TTLMx55ZE4zt+py7V0d
HLMishxxyAIQhwonAxxp3+LT6IZ+AglMzrDmAcH2xeVWF4Y71TlA15JshEn454mx
JatA41gnchZra9F5DPbP3NyqFiICVDgftH+nqb4RPEncVWsvsrsTgaASeAHLIXGH
rKQwWF4VLQddfhZPIaZ2cOQqSUnCJ8umKymlI6075jsY7cYXXF85PE575lB7dzdf
CD/FknCmIUaQ5um+SYsnR1ucFsXRNB+gOnpkkcgAo3nr/jxtTBPMUVAidcX3xFQ2
YuTR7lqXHtGOHO6foyAJFeLyrzfm2dReXF9TedUEy6xhzouivA9kE/F1kTHoOjD8
g3FL1EcIJhoTw6Uuh8CoOHAb0mUIsjZkGYOzirEc0lfri7euwhTO+50/n8Z0W3+e
JiK+B1NXrZFhbKf75b5W319UH1+RhfvbOGGH8XOArEk77INEILtjDR+M4davzfk0
DdGqgbvQdCIigldIpOKlealyGL0nG1t/bnEBxS4a+4IglyENf1eP8zca+EnyHAAe
rFOEaUgb0IjUXJztVxucoZYV2QS2vT1qoAZeaGGSO0kqrwCYQOW9PZ+jyjXWKnZq
QoS82WWAVHi0ms6ksJjQAtMeBCeNu7GRpX8QfMrlCHDDK5jOaBEj4g/j8ZMtGiaV
O9E2Ym1Yes7/6OtfPVsogPhO7bvaz735FAjkzhtpu6eOZPwCka0KDuzxF5MpDSMv
+0OSGtYe0VFGf3V8dAJGJ/uJiOtdc6FRaCTbV0VHOo1rItYJZgvTtB3z7PUMN9t7
VigM2DNf8+rZ01MMk4DFiv1wRyIY6OnmOhPp9XVp2FRNA6zyzpyWu60ur1Cg9Q+Z
7XN54qXz0HsgmsCPRzZKSlFD/SNKEdpYIVafHjS93dJZ4ODJfiWxTqYOBKnE5F9b
0C9yePk5cMKOzIU3algXB0exUqQ9CPRMooC5xuwvxzPUbSJRFUNgP+quUPbSqE4l
p8aRVcJ1v2TIe6wnUQUVZ33BNDrm/AZJPvLkkZdhv8beL16yoah06TwlrTHNzgF5
z7ceLfJwOWBncLAuWR+ls6XGJFjmU2AoE+maXFrpkOyD37jIKQXGh1Std0F5VCNK
UER17m3IMz6CEovZYMTcZHe6OmSS0YBg/6DO2RuZ2i1KTj2CO6WOhuUSvD4Afar/
0MbDt7CPrhBtN2sLxsSmu7ar+r/mhaxilM6dAqxg6tYqzMJWBSadHwrc+jLrAHlu
6StUN4fhtsYeI5IM8jpzmZdw/AKjyBm8VH6N25jm8fs4pXD8h4zAiK1fUlxPRJRW
5mw16EZH+y9jp0jtesXH2/Ic2dIgZiYmgGLXqRwbHUOfDRboIgn9Ip1JAZO0cG2y
6lOlRKQxHdiMX6ZAs6h92sxsiSnNFN2F4XiB9vdcFyH2m8L09VkihQcCnbhpoLKu
euQdsDmsLyqZJXk1bgFaVNpK1dzX/DoYsQjK+DwNR7PSlXCR++VqHbqkG+yc/2N+
Z7nC9DveKD/kJLAbSvTJXL5+xXLgvLn3/Sjr53wyT23oC+sTQ80CYDOWAoIdLxzC
g86veoKBACbfi2xOhODDvs64jasE5bh258/rzrZ/2y3oG9pYZ6xu382BKcfqhXrQ
wGLn8OwyObs6DyPInE10nlM5jMpBdHMs8CJjmwiqZ0+EvKDmRAv2HlyHY6GXdIgS
1AWFobG/sjgUJ79slricLUNz/9R62OgsvCvwhct+OpzzsLdmap9RIaZKLxEGmr/e
Azt1cp1f/DWTf3aBus6VfhpiSnTBFaxJKIUtJwZ5NafEwpgB/WlNniTLjfNkbYIp
YoKLCn+DZa9KqxK/tqjUna4BXXXQZ60dYXc8yl9b+gz4/vxpX2ARbHqNR2OKAB5X
ZbtC7H4+A80K9ZNPeNvWrESRpvQH6GAbG+CLpJkYGN6Q5Wpo1hZz/6IBtXVXNxY0
5250UWNYb873RHX9LZW91ZuG/izaXEJtdTBK0dVR2XjLUay9RkWaNGoc8JvfT/gG
bsFYn/sGXyEQkW/FjR++vYvhHiIQzoxF6bjW+L0PiZV4OIMN2xQhbva/GcOqUaop
JGvP8bVDWub8a5d+/ngtonZit3MwJWSwl0tamN+1Ns2QA3Z21jNL5Zpmav11fi5r
+/pxR/sb/IlzSGX+Eyrc9C4Np7dA3s0ZE3ccF44bsKFiR+DZrieQSqh4q0mB4QiV
OBHEECYNLlEQKDTUR8iKAQ5qnwUyNFkQlPRn/WZy+rMCT9j4zfmVBXn1IaCpK1lg
qBacuttWSjqucgFi9ypdg34JymeiQvgIl5qMVQhZejQN3E4Ndam6kQQH8Z3rpSd7
OiQT4mfTXCQwqCV8FVye5mLu5TKPCpnb/z2CdcMA0Douus1b2E5ZE6V9KMTx09FL
ovsU142nRqzEIREr/yJeDHhIOgirBrEkbbbT3kwL1xi+cPsxeWw+MP9xdVm1jE71
QlAd2Hb4Zotppv1wF5xS6GhcML2fjk4vGXeOqBCSiJsLg9ti9yd3cwfTdUgblz4J
bEnkMVjcMWyN18+p9RO4HPPw0sUEnYxbCHQgZT8DHCatxamAV1A3EcVrP3z76f2P
8vvXKAvDUngaIIsD+Zt74YfewDTeBoJyrX5Wu1tg2JKjzQET2zIRk855eewEqqU8
M/cEftXeQ1GI3vnoUf6zrzwaf6Mz+x6EH2Wr2mEJ21ukTrxIj4E8iuLrrlkHTCR8
OX6mb7j2TT6NO1fClbKjnWrxHg/UluZpRQrB5///5IxeXxg/a9htpDTrnjuhfTiK
eAciNkiRzLax4aBqd3/Hw6sWvtUD3sQOkTqmOoEM4XhzG0Egqv5z5ZjE/C0xGdVg
FkBju2naAvSJ4GMqhQSl4qBH2hJ2eNTEUr5nD3UE6FPuOH4mKOpjXYqhLBzpOx1H
I/LU2J/CfLoCj+5n4IScEhz3RBZTqBUKdbBU62cVUCk8nOcOW158EtBnwHcKCzY5
VSDX19PtSlsVR3KL1DGFdBc9bz2x/XX2dXULvpLPb1TTKzLDrTs14nobr+hGlenT
/kgHl1ttKLlTJYSMFhSAkAdwYnCgGwjoUmUyrSpfDvTtjtfGm63jCWFtWDSjjXIn
OpcwiuFA4AD1p+hFmiH4A9F4Jz5CeJrpNsOXYOrZlUWU9miMpq+00eSLDq2I14jT
up+RL5TlIxgIHuo4Y51qaPfZnDx89YuafLiMTz6TopQAIKddHIfm8v5ImzdqQ2Wd
F8O1TduloOqRt3gx6eUGIJvE/h5mo2zL0//PGSfn4k7Hz+g1e/nRLXc4MvlpgzKy
Cx2KKxr+2UNPBC5z4keDNvI4bMnA2YkP4K/zikaWkuLYMtyIgDNfEXp2Ro1JHHLI
TDmjvwMtez7xhFj8ZL9CJfflRGSsHM2wzSjaN4azPhWYt/+0Tf+sg9N8QmkxDQri
IWa/W6GRAAaL+NwqtLFLNolXtYh6JzTi6Db6XeSSN1YEe+0IOP+wsfWkW0meeCHK
/OzGwpSa8zv+G1VuvwlIlYm0g/yTQA/0sf80xrn62uWk9CfWH5iH1XOr1t9B/RaL
zbtlrKvqpU7MD2bagDPMVXelQbbIdTkdcoH/ggSDwu5RPoMiavJIKYYWfvEnM2i3
YBOfMu9y/KqOzMrUu3xOMv8houT0MWsgW8uDd1BIC5/vNhkiC2CLZxaJMyhSTCIt
Jd4NFMjLM4qPN1+pEiFRSflXwLOyibrzITKeiakDEkFIbXqfVZkLJABVGpshpJmi
ucCvbDau7CNoZm17SuIqmPKTzeHlS9QcnUTL3Ffks908rinsFTcGsvzOS/bNWqvv
RVpNrmAyQ3ucpoKy4RJPjU64bl1SJUAhlqD5A08Y/pfzQZxid9LnkV/ttONcembe
g32E/TgJ+uxIFESCkyPVCdqCgO8ss4IfR2a0mscUEmd6OopFdxU58+yCg/n5nPzL
gzOnTPZNCUB95pdPVa13Trm+vKUnfMWzuwhVeSYGs7hcL+p3SHrH0YAqsl7gWqdo
aVdLDJk67kow6kII49jrvZnEUujKEBjVm09hyxxgMv/1AV1DQyk+DuRJKYzuXPQ6
VPb+fiyi8FXWEPS40JlnkqHUVP9HsaqZKv6p4Bk2z2MSOG5tmbXhOEimIhJF7KHr
bs8k/qVu5Q2cm1xigrnzCxXzZY1nm3iryEkqMkM47ISOWmwFo0f3fT0g0gpX0Gss
fdMy66FidtysmQrlmFtQimW++saggag+3maUsDwTnN5p5txsc4/GRQw4NPm+Hk2B
2aEFHFqrV1a3Cp2ksf0oBE7prtjNu161HMs+NhKe/N1RO+0cagq+12hpARCBRGzZ
ABbhNPE7VPcpruU3Ga4KSNb0cnfhs8y5ULP1EDrx4JJHUe5ibAvzxT8wwMM1exGE
RTFZ9KBFCSP+cu+gTQCbF136tEXyPPFxz3ryy1DTkFHkCXeOlJaNfPS1InHVT9nv
IbkE99ABT8Tj9WYd0ykP82SDBzANRWqB8dLg6ABdcK9I5KeX5U/YWDE6Cx3HZfSg
48PDaCkEqiL1OVarbc+2BLzrVpeaWrOvFSKDfQGuCFY/+4WpaPIgz3C0DW57xPgJ
EutNNIkBgkN4LS2lZOoej8SwciQ0Q0GJncaPMRJXdR5ZpsK0Ak54LbSmnTolN9Oo
w3m/NStJDRixzs6lMKKbrzeJlch6bsqUDsbnz49uK9NchHzppE1RyEpo7cwrkqWm
XdpoueQHiu5y0w1gPIxKYJ1bGWX6Ai0CpHuwm2D56RYBbIvmxyKuDZU8ip5PSUd9
NHdUAPJBAR7F6QCKYXA+FYWwsjCQ+0yiujypNctsqabdDx9/dF5E5u79R/UqNa2S
kY5f1SizFIMoALOYoF3DHRph/IJsNnA2BKstMxy0J/O7lkaAW+HZOj3NFArTmUnI
m3zmHUGOpbceCUniE4oqyLW5wbApDqSbhiAb2j9Q939TPiTk5BXKdsQmSVNZSXA4
UtgPN6rGR9ef1nXquGkPE+7tMdm6khsUQJRqszVlIGDRBMGeNwklrgvAl493nV0g
QsYOg9Tl5laLb8UQ2XyjcZAp9Vk79nAtNKo0mJaEQwVwaOKylT7bZd20wrBKtKt5
/0Id0voNYdeWqjsTBgfpT4LXaQ3FVB/Paz7vHf5ftYnLV+1YpzXq/NCMZ4wcmlb/
Vor0bCHlLsLkkOAkZVK8crWWgQuSOgjCztM86bAsMUqMzNm+UdMw2t3qKIOrMgdT
UFXQ5aW53BJyHJprTjhWN/91BE7oBeRL0UPEcozw7FVbYutAhm0qhiBVeYYgpL2e
QZP/iZO8Q/8OB2kqRbcBtOxE3ExmSM1Jn5PwSGha8iVu92bMEWpS14r/R9Y9FRob
GzD7s4WNrA6tX93H4P1YoghNJEmVMrqU71EeTCxdBawNDn7QEW46OBUkEbEZXutu
qj74sv5IGdVk5nYYlsw6vCzqiiGD4TZ3xA3cvve+4fu8INociJ0pARHcCAQOTRJK
TtiNkbvYfCXvx31Uc2vqvWHK3Q0rc7NYgNYFzMNlxlnDNt4Vv9xHH5kcNp6LHXSN
a9fOZjFUy+YQzNTjZpOx2lNEL6DRE+mxtpVx7R+UXNEVMPn06kkKu9W7L7h3fiXK
I55R5dJ6pepOyU0ONpkZ++ltLrTHf/n17AJ5k6S0EBLTo7CfIQB5OQ8SsW58mhSw
oebMcKkJ5VlB6Ere2d3rG0JYlD+3W2PQo6gob8YAiQgISI1aknUDzzGnb02bC2/H
GVuehX/M45cSVtLOBDewSTiyNDrJcQD1MpYQRTuZ575XgajDB0xP+MRazRoR31qo
DEP9F1+fsuTd5XWgaLALtCbGWVWPP3EWtTEYn2d0I/uGHhofK1HO72KLgxNceJLa
kvj+Xi7cNJ0A0GB8TO1vnmLHbYwxlCITFqTBb6ICobzkYYZCfpr6dAsOxUARTqFa
6ZCU52k84jU/FI440akbIJT4uDm68PEofKrJ0kFZWamaiz980IHXVOMocTyqk3eG
NxPhL8hjL1XJpm7MI12AHqYOZ45zJBTygD8C4GCukPwO8GYWqCqcGdtf9YfPDQQQ
0x8Gh9B57V83A5l5zQRmC5XYXGJapxOJiwosS/ZLRRfGmljdIcUryHkR4SO+ZeKp
BRpfTU9NJebTdHFAO/CxP+gQPNNn78PHAHMqr4f10Lnb+rxWgT4yvoyNx1ITp2z9
8zZlO1ZC4LXgOLf+IZnwagfk9vqK9AozpxIgw94Ym6K9jc9tdOjNq+/QYVKXaz7E
AIq0Roiv+tCByQNE7Py2ksra79DNmpRI1wy055Bef3ExSn/9MHmmEZbV310O67Qj
sSS7rYNc+0vvCD0gRfXpH5FLO7debeZEZs2evDrCpkH+hv7o946duhyrP0j8gdHt
OSUxIQGYs/el1FAe6w6YxQQGtxMxVc31jAqdDTTXoLqBCtEU6ltqvv+H6YEiLBM6
tXKM2m28ugVfnAvUS78Oyo1H8j+1NwfbJHI1pRFPydYV4gPWOKNCZ1nYw/xMdzVG
/Sf1PvJiI1DX9PEXEUJqTwT7hGI1iN1tw2IStceAcwYxuHPuKdfgX7ocqtbjtxj0
k/Hke/Wh3BDjWFjR8yiZAOH+3R30IEY286dZN3wgasQ93EbyTI+RxbxSsEovFAWI
3oNddG8qw6YJx70sJMEgcSAXEI8hI4bjxlBlKy4nEaxi293GA28fEcJQ/6eRX0KK
nNSuMGbkzbd6L0Hmfxhi6wiFl0cVdwKB6fp/3SZzm3N+V0SuoYSTyxjNf8NKVlLs
zBMce6F9wGhpQOq8WN0TtBDKadqs5OjcE3adEoc4EMbXhwfLTaJShzpGRU6eAR8h
7VGlbhL1uSJfHQb3rj0jycqioNa3C08Ew3+HrMr/+4YTFZN2zDl+lOhGdf6f2+OY
D1qfzLV8DhciIZ0iUOzKYB8aRvTmUdFpNwCKxB0WY4o9Ado68DODAPaRXwlmWZ3B
VHWWmZTyLmeouQdHVUa3gzDx/sqoN6ih3lYHPc+4ywEyva8ujs/mr9EG2glNiKl/
snM02d4CMFcPHsJ6Jk8dDYIqKzoMwY4ClhGnxeJFZi6yRS8CCEjFSnF+2vySaJkB
ZgDfZz/8LhaKJxJOnf5M7DoYx2p+83ith+PA6kpwLRON9ceVzXUdtyvzUXU0VT7W
Me+KQOh4sT3NN/tuqToXcSoyoyhcu3ZxguEUwDEf9KmtSsqUUeLHILR3AA+M1yQE
ieWOVcJOoJkpdG2CyhAGGv6+DyH/fa4RpKVerHCv3j18U+uRtppqihCJPyaDAwcN
3EzuRzoXdCHf6EJttzzhVAPsDiBjXc1E3UUUr6dWWUa459xgdpIpkpBpmr9ZTHmd
F/c9FC38BjhUg0L5+nwOMiMlBkUB+/4c2onTIxzqDwTlb+1NUhHW1VNjyLyGgY68
mvh6ZLZ2desUgPjUfCKbfITvJxMoZ+bt9iJo9RYOPZaiQmiKaxhDHGyxgFtz8H/b
T+yeL3BY1wlL4Q1I/oRjViB15aMRH3giaz5KnPnZjv53YAuTFxzfpXFnLPnk9fRf
wtzPHrAzzGpevaBrlHk3Lt3d6mbyOkU//pxtFag0fbsChVEZRaeZyduMdbtUjjiV
FxS8ohySXsJDSBfW9oxnTm4Vt4cCe07YAKgh+X3sOIAh/FHXP06x4BtRQvfh9mgD
jsKmM5AhKPwObcUuBB6VZX/YB/xKla1TJfsBfXyKnUSnp5xSWlclQ+w7GLClgWLD
Dnl6z/GbGomcwZ1DStmdq42cta4l0ww+Y/RZGEaxmHoVqJc7UH5F6WEU+BV2HHR6
FQE7B3+EE/mw5ju7rTzdXuPk5KpnXu3VS9C+C4t7OzLUtc9XvTT75Dh0ICGVHJvJ
WV5RzgsO7NcSNQlRLOj/bmtWF0tkvWfHjTR4NdD6BICkxUDll0Uq+kcbdt1rdBWz
+2i+eZeqSBnXPB7iQyw7GeKyjpLteHaKKNvbUNORyA5+hr6sTfwo0wb+PQf21Lav
uVfYzJpgZtnbRV5WQqemw5MTgtT/+MQSDRvk1GCb9vyG7brCEBbzLz2VehXrvATu
w3WTYbwrqdxAycI6d2f1jB3XXZiVUtqtFNUqV5J5e6BYjEwVdGSPi3NxCQ6bOeFq
8ULa0pGyevU5HRMUm/GJEItCQRLI0hKeqTfzbd6Gt07SW7thJETeonNzyTaKoWVz
B8SEAp0DfZn7Ku3J+42GF0SEAbTMYeL7wxq2jPUkekOmu0FHuuCPYyC3DI7ccd2E
1pUaVWvVnDlk0YzCpXTLuX+MVZdi4RzSEHzme+JN+pxAwfcvZOXh07a/H7f2+f0u
VVViV8u0QkvT8MFUTcCijONXjBHFt+5L4aFrwsmMhH7Atst6jqZlM6jRCNpAIdVT
Yk/7EPOhBxAZW+doSXkHhXSDQfGG2/83RwHCM9HEGtfGDGX4dW5gNdTF11X4TcAe
7QRbCC8XEXF5rnoFKl+A+vQF7kPO2PofsMlbRMJ91thy2uzY/coP79Hzq1F/BKzE
tsnamUQDYnDnJ3UMmtLCHEkSs8+2Fihy7g9ub9bncz4BdsjzY/wtu48uQIXnqIWN
Ze5WCUGF4ILqrXCNf3qd4IkR/2eTuxuzQFq0FUfB5+kV8OW8rqJ19eX/I1lFvUDC
5IhvLp9Qy4ZKMGCm548fmHDAGRd/eYUyudiMMHN/CK80vkTwIQTyotZkpFgzHRjF
6LXJpjH5W7XJohHvJ1NUawicp4bcrS+xWK90amDGa6f79nKXyP2hKVTExEvFyDqJ
sxxIel/cvnwXTefbNQKx9UKiniBSEOREm9mzZTKpAore841D4ko96Hny7LdQYiUQ
MDNtOqeWbWeTnxJJCLCE1cD8jcwBjFZMUuyO7XdXn+qyCCR/OmTad6cyn8/PmqiH
8a4aD2Gv4waMZ1gl8Na6AVgzwI+gzsDX4Jl5nwiKhhyTbgwGXa5Q+LXQz654ZSym
8FEyOX3RnDyLmJdtiKEA6IMu70GUn9F1+9JPxFGeM0GLgwD2k5JPXS4KxshYTxJG
4ecHkKMaCFfF3bLyNyWffqiQsWUQCzF+hHwiItxVQrKQpAkiZgGW//MSkL1jk6Yq
I3riY7nmCws2VsXcr1/BRfNleP+gZFx6CU1TUHC4iJpDGdsnxie1v34k4KXTHkBx
cxBIENFlknRXJRrNEKy15mDMX6mVcTzvWTzEOAr1EP7xmg9d9hWCgplQ20Uw5djb
Kw/PEY9THdw01CjgDgvR0FJlt1HkzaQGEmusggBXyH5X6zxNdwdHRGPz4w2h3F1O
ByRgd0q9dLHpUshv62AKWAzAYENsy7LCTEIkPodFuu2Rvk2j4bmCJFLLzxIysmLJ
yLJSPGsLf1bQwoVF45+8tfRomn3rbFrFCf5x6+ZQBALHRvQ0d5L0PFPnbkc9zgJE
Tfbnty3tn+B7Jdh9faiSAJYPnbkI3VmDFFB+pE+lulKNSE/giXVD9cybs7mkMC3/
fGOzqnHSaQnKfSWanNJFdrl+t5lZ5xVi7MgsttkBX4X92MQ3AefepMxmEeyXoIIh
gbx7VeNAtPmUn5NqiqDBk03xkTbcWaARRVqmc4PmMcfsIoYMWRcjThYeIv625iX1
OPstWJxkVxaju6FZLnrT/WWtU/fDdSZC/D3WFKyIqzWmQ9ybB13U8v8nne8HByw4
3pIaCSt8y2U43FugYCGDHVD/048p4uDdfcv/GilLpSAi8eYll9tPoZ8xshhzv/II
mKSypwEnpmTpCW5dpdNmzlf4Qok9OSCvs0Hm5ru5wJ1DPw6RRpx7xHbynu659L/1
zfkFJYiUIDSMeuwEa33Dp9n/QkX5ZUJOCzcP01OSwBU5eBPtwutJPJBZ9XPL/jMj
lSzkJlRpZW0fpgiGutoXLeNcbszltNfxiMNz9bgc/B4cps5xpZHFPNd7rKFIv7bf
jeUBnz90vGuWmwLtUDuokBu8lmQtk8Fx5orvsA+zlqUzBXPm4qJqNJS/2hpwQ1se
g41pmdCU8cHxa6FN5aKyi5FYPuIB6Cj5f9woOIOgpcE+DA0CRebLaM6j6kZJkab4
WUR4IZf/uJqc6evcuSQAeMBPHMab0o5t6fqELmP0FsSBaEoyO58+Z3mwfYsMtJwX
nB5UxpS846vknSUHpqQMw8szEib9bG51nzhTaHxigVEL0Szcv79TBGtJgGJwMP57
JnHtnpZuqzAxbqevEfjLd3EA/UWmEDTRW3g7cnxBSGVDkzMi7dDy1aNpJOsG7FZC
/VfAveDPxFmuMtyH0WhrJVrVfDfRrWFHwzdMooHD+oZ52O8lik7BwnaGxd43glWF
PjilqgoP5QVPkVqu2kIcXVaxs711URiXWOgPcehqp9ZzsM156LgbqRyP3k80YML5
Uajub6gAu44fovLAgZIy33dyIuDK/XmGJ0EM2z4tmDRLCAqKjGZ3OYhDaSi6Cf4K
BnwAnzpItS+QGVBrHWa1fxu7SRVXIVJqSO0rYl+bJFjTWi3fFmPwrDpjRtZTPgsT
pSGNei8s5gJ5uEVnUwHi+ErJHgKOSfwJL6gX234VAawhIXkS6jy1/8dxbFmGLfr2
LeZWs1arFLLYEEKHnprxFCWOT08UGMa2gutwM/EOqvFnHEXJeHGSnh/sS5hsgEWv
gqaViZz508Q5sL2e3WVHiUrvMgh92uY+VkvfU+PUYbYnq4kGzL50aR+6RTUxEHXI
XftmICugyupCt/xLgzhsFI6zs+xDTrrNV6NB2pj+NFxIEDU1TkqQoCGOwnOSA7eD
VoJsgAqLDDzuqPfRAsVqD8MxE0It+IAM1Tst53BuounD4zta3oGrTiCkfksB+0QI
OeKN7KmtgkpuI22kGCWQOUopqkA5FkDX1zne04PYIemtQXUpgTMcFDkkY4Pm3DP6
9Hs/fGv+YFAY0xRYHKNPzU3ROzp+vZNrLDPo6qeYyTpfdLmxOyYfzGELCNhKt5RE
Z5+6ZoPNrV1WmjaQdvm2HpmAvqFsMMqHsBSzHiVT2eMcMe/3jowB5+1CAIEZY4G5
51bsUZo0Eg7aGYPfK64v7YHvJZH4nMKf8GwHjJmhwstzk8cHH78l5wg8Bh+80lhL
T09tQ4wcN6MgSR1O6S2pzQZqeYnnbxNIfmEh2GZlbHF18gegbAYXTxkVQOkqeMlX
IFoujYXHsOIO6aTKlR+y+cXpC5PWbNL43k8Tfn2aE0A+16w0CIUqTXINrrg4m0wp
TVUx/3A1yIp1cw/mlrWk5LVblkgzQkwEpl9nyCIriCxLS3PXdU9vV0fbJPvNzER8
QFZznBjPF+tDwkRcdKwCAY29vp4XOBExika5A4O3ixZogIntvt76/tN5tXIDNCHu
ahRVstvXi+JarnWsaEF7Dsw5tO08AIUcJYesjHeR6e9/jpzyOV3KVMhw0+p0IRk8
I27Eqs6ciMy4MjQvYUvOhaAshZk9qSHkwQ0HtfToU4DdkTy/1gvV0/HwtFPb3v05
Tc3OMgxTuPnMSYBbivBeipPCf3ga02Bw2Z4ccEZz4yZk0TEW4Fwy+g+GGDp4zXo2
sD2rMUZ5MVqNOZe0ftTU65UMLjvmg9HCr9V6e+XCh20b2BWpPW7Ngs6yeuD3tXt9
JTnfg/LzOku4WMhNy7eO4tplgu6IbozV+aJ1OhXjHZYP1pXHTX2i4eX2ak6+aYtR
ujPE4vTVJeNumkQUeSpfV5krJ4aYKyRhMS1g59ROXMVnCvqEH8qfps84GnpvCooA
6h0ircoOQ06vlt+ho5ZmxapsSRkErbOXaI8IJFld63YbqE3pwSlwXuywcC+VGkL3
C9o8kHPBqPyBpGXwqP2w5lCKTzjsvp7iQiAyQaIbRSvnx46Ybl0mPnNOKp4UX+1+
7+90CeyJkHc5YfrhQAb08FeT/m/XyJvhTcmnF+Fv7wB9pykPFQaYKidxzX5lRtMH
/1fG3gy2tXfI5BO3E7r8qIHnjtTPBtEnTynOy81K/vYVPp7XcgZhjSui6niEycjQ
uL7Bjb1u8zBzuB0BDpQ7yibqSS+eGuu18x85j+BVfIr4tU0AXA4Nacwzif1mYG+z
z1OHwdFdy7cNfq2wjAhHmLdP7ImOiODEgAYH1jCZJcSrg5n08yjQK4RBnbs/NkBF
+qpBPFOYtOVzsN/W8vRpHhQXsLVFcP3GB3zm/T17lbetS1ATdNixigdRVy7rZrnS
gF2dLod0fjtWlNv3B7JnFbi8HrIHSKKYX3bKCi+QKrvHdxxESB+4u1yQhwmI00zz
HvFIvxRcaWi2toMrsFiR5E+xr50AhY8HIinxlUgf3/vurJHy/TF+q6MQWmGvZsvN
/0F3eyysyQCXLU5zLzT1beGzgbJK7IUGEn0A4Jzy74xBaajW7u5xMequqRJ2DAgv
ZcH92GNLU2lAi0ckICNfpNtg1Nftb9Eo+/mVuYyg0VwsubjRbBu/HSIamhUKUQL5
OmEjLXol+IlYanyPfs2615w+IkunS8uTwmGTP3Hj47oh3lsP+39AuSjDYQ12qXPU
nSDy6nTBXHnFgxYo4SxxnFadXfTK801/8yR2+Nk59o6oY5ngYSuQJ54IVHMYuhuh
doik93A4OdtW1ST4QfLJWjDhZJCV0O2PrMo931Uq0W3EXFFJIIbrdkcW7H8YcqjW
HcVL4ACq+QL++H7UPy/BF09IYZJzlQjNQmlVRglyX8yW1xALlPPOr0zI0RM3ta2h
CxUVvYXqmktcqBIGrJgA2kBCzu8YJUgQ2jZxyJMGUpQH7+/++o+gULyQZKCyOyfY
pCpj6fwJbZ2N7oKj/IVpIjVKh2I0VvGvyZJOdC//lAmxuhcytD3LREJx7vBbgIZ/
LRl52aIE0GgkaY4UAxqwwD0fp3fLjl9l4ekHZgjrvY21GCrTlhAiUT1KUE06N2lT
33CeeMPhIQ/bUrMwa+5zPE5Y2Vn0LCau+7MSQbu1uRKm9SxG1iWa7W3siuP3/ORe
4boOVUTHKc9rVKbfSh3Ezx1fYAmftwjilgCLaSb3kxOfW6U/v9PDI3aEBI9ru+G4
DAxjqAy0aTcbpJ0eVQtUQxUFtNuBY11+HjPdMD3qLKqMt7dMA/7gxzXkyg9m6rr5
C9lGrfUHs3EaSwAJO+2RP65JsDX86tocaQ7O8OFD4Gzewpfk7mH8VPpni7o/t/zo
kxE4qQ9UvfgseH2AAa102sFPgAlCB79KgNztBBU/T6twxZzCPkSYnwz7F1v0fcvh
g+R4CTeRcC05zrTcMoxytPtIdh97KFwAxBJma8nf4AXNgB+uzbJ/j4Il1XU8IOfh
YSJKmiRHQaKPv1SXIzcPB28gFd4CbmGm/d4MiR3ZPoSUnFwX8GhuJv6T/xtOp6+2
fPQ6G16PE554MNMt7ip2Dr0WF9YNrPBFCh19ZTXaGmwUVqveQYGt4N7sHdYjOnd3
3elEzw1LUPYVeuFGk/+bdW9LhQlwa6Bp6/kS2lnDgWxCubmOUTC8HBKPrwOwkrPn
8P7uyUAitB7eyCJJO/VCvxWBUOCj9EaG/V1WhSdIgzjHceo9gCPHConYA+oN0CoB
QFhw0piDXdU1YIgIV9dkaY4dQiDqxPWn4Hbzdkwa3W3+M448cphcoeXoimIwS+g+
tXRA8M2IrerdT5VgiZnyCL01W1FjlfZYQTwYklyMxw/9GR9GF7yoE1MVamQ8LuOF
hmccNPcA1ajkyoySgAD3cNsjDdQluUbVUh3se2sO2KgrsSJli5NBOWiu+PnbhidB
aOZEQFIHI8HBSEYNmRBrDwCKqFlSDdz8BywElIc04mDiNMzuLYD0DQwswy+Mt22o
rD/eKDG2x96fDYUDbjK28YsiF+4Ml6aImCWMWPqZj8pITIBRdROqr/KmRnNp7RZm
KRxLTIXwFjZUOcel3yWeyje3xSrid7o77PJ2C3T+RvXwb0wlWLuhLfgkthnvzjy8
coZr1KZErJ4gxFNqqs9BfTtAsZNfuKfW/wG054LINVT0q2bK3RW48K1zej5DADPa
a3p5OYyrSYTw0oAvNuYkmEZAsrD0OJrVEbhC4/q1GchhAEN4OqqfFlKTQW6EfkhK
KeFHloH4EXP4ybOn0DDu59WsQugjjfSjLU7Ny5mBVsHiM/2DFbpLf1LXsRA4M+NB
Pat46vSLGOoYT6pjh/aIZwU8c208kwzypynMA+AIKrfdUYAaTpHEJUbWtvMTP7sh
bLh766cyTbVhEofUnXU4vPazNvuQsbozzsQ7qLK1wpA6jhv/WuAT53LuKcqAEhyT
/4SvlUgocm2jVriHXnarwJqAOMFD258mCSN1VTyZuyWeDcDDdldzj6duBUu2ALoX
vzuo7oF7VrrHR3vhucXQvD1Hzc3itb/MANIs6DSGiOsxwGfsq0r5om3Y+EdYvrui
BVayZbma6axJUsRTueOcF+zxywUit9JkkSJ/JKYUs+p8enASu1Q34H2dPD/KfjGq
mbRz8BRtx5Yl6DubXrUc/3DrVlq8ZYw8nuiUxXXioq18vL4Cyv+URj4+EM1sZEL4
VwZfxuBO+QMF+THakawV1xn9LjNKkYZYY+cGClp7wO+8f1jhfnzJr2aHn8tLQbIp
ttal9TZOjY6c74aw6HRUhANcB6k6M+/2FO6mZUBu4LOafSB1XVqLkl5/97D5lLDw
MKZbIFmOVKkErg0oJgL97D3qxCMjgpCXswUvnfMG8myJxtdyW9mDBNQLKvz7fl38
hbRWLUGT71YtiPwEyYunErYg4yoiE7UsjQpInMmoqk6e4IE3o3Gs5+PtOBjIs0Ax
818x8JrxM+zzQQyrhB5o7MxzI7WigMGAXvMjefVgEpTdKNAbgycf9Qhdie2XiZ3O
L1szwXGpPIsJUHl2X+M1JOOYvRa73kJPwV6UX/KtIKBl/UeNHndzDfdMw/K491Ta
xKcMtZqli9x5+nxvHpk2euTwCV1tmr2O8SZsPApYzxGZ5y8qwJ0uklepGr3fEnOb
T0glvMINtx0fpL5G7p/qS0cp4/gJSMKU54tpK35to0PJ7psOY5v/dHmeOublVk0E
e9SDdFoiecFUBVvzib1H6khiJREkbHBZ8mDzbOTD6S4iOygDqwgLcihddB2M10KU
5pSGP5/Z2CiHKp7cewnXmvb7zapF9v4mDRDlEBnBh56uM6SyCpkzbrGNxDqDvLCZ
yXwWYgRagt9PZS8Of1FwprilHEJn28Bo8TfpymGGLsVxJ2xfNQaCIuUNs7dzqFVA
J2S0leAq63nqHYu29g6ggw268DNMaL7u9AhSOMXEzYZVU1EgZlyEzOD8fMu3OqLE
swoKeRtcfn9Q/B7ZLvtQDa0A3pKSHxLp0VbH4sQxASiMWVuKdCGUSU4dUAkgDhV7
rEo85b7hkiSVgDTg+wLuMuJQvuaDaMhsdIjtN6jW5J5ZC5pavqbZgKkFSm6rF/ov
JWPokkEaCJwM1PPaxdQErN8PT1KJy1UMywoTaZ+/oQDRfnj9ErMlhzrMlr1n5jts
65w0wx6eeWN8MO50rOqZPIwL/L+Uj9Xcd1LYBiMhZJmPmG4MjvX6LcmDz+qW0XvP
JaBh0Wo2iqgMacJC+Nv0e/NOvitXT+HpRpuG1JJl3m33GEDINq8pZSHHVExlNOVI
ShWHNLiHE3k4VUq0SfBj52orWlCGmwfUnf6WNRVsPBLEPjE2pPiA+ZvDvllGzyWQ
F3ISwIUlLTl9H4BR2hQrZ9FyzsM/sEJTOsZZyArACRFrLvqRmPVodlaUR1aplHmn
ygiN58Os8mAYf8z3ScX/hEsiz3SY716/zyogqAS4r5gSVoZbo0L4OeAUgw6pxaKw
iGk1Trj+Gjf4rdz4USkBqa5wYpDLR5f1ZHT+O6jb7dWv0EAVjyXWzRNuMs0YBXeu
3XIs26457g5fN41boMk5Eyp630dMoiTVNoy7fMvmwzG7cwVeVSrmiJLKDh6eR2mj
aLKhg+6A61z1NlRp/lg8zQdI+sSxMHHbde5+wrEjrIPIpas36iuK56o0TirxdWnn
PxRHFlNtUP3UikbhI6mwBsus72NUMv/qqcgsWEMFxLtqcr08nTrIug5EYO5FE+jh
F/s9shLZfBAfnQNXJesQZEu7SJhmEI5uljzcAGKWk094Jeddgn7CcWZSvxGHv3B5
p5wBn4Voc8d/DamQulXHHU1XHLA0u+nl7F+PVELqObrjc/hpuoclHzlCX+7U42Mu
FdTkr6gtNAKDer1DEWAADaHCRDUnMXlG4afpQyC4OgqCgde+ouripZVWmKfwvJaN
cQ8qlk94P7zuAsOL+Xfr6r6frX5TgltAsVXsQe8827MasN5WaHc2/7hI+NlnENxC
ZwMB/IXoVq1HQTSZXWVKvYcA5Dqn8xK99zErGN1r/M295n1ScNsye8VPgHvPAuB6
amIjcINFWc89+mTAim5MnQLbkfVcN6r5+p7t1Ia3FT5SdcIGydNFEvzdh+LJrsc+
r+VoOvF4/QuOkXCy2nipqQvTx1pmsIhAA1MB+yzo4MbZP+i5FrED/DSdrNmy1Gdl
DN2t35Nv/W0bSCDc2s2sI6ZffjIQ3mLB6n7HCO3om3qTv//3vz2fzlz3NLuJq4Pi
olzINIuO+eJqcGfLf36FfrQqzT1gMAUVEm1vNx+uTLxWTxYiOOnuZ+tjwy+kwzsG
ZeG0enq/KOvyUy3SM1pwdAPl5X+hRrRCj9pHp5yrvqbDnU5WzFvJXAapDjx3FPT1
dFHDpnuHubwPAB67N+fsufncGNsnzfEjonLlIADveluIEvwKKz2scIVnIj7VB7DS
hl2wXm2vyzYNjJXK87QdQ8BmEQYgQebQJyEMYMaplqvC3XoQbgY9LfBGb/dWZvpd
vBvM8gM2gWpNNpCu99a2rp+/CbgI8uqjkIIebipsG67MNGRA8ROJ7TFdWkKScRP0
2cdaE1fhE5mZKUwpxJrUUklZFSRuasiGFhga3JsACzkjPm7NKtSDVcnccBnD4FuO
3RD2RlR2pU8YsnEVAO647C/mVGSBP7Un8+I+nkLboPlYmHxRxIELUoCfNqThcW/b
pYUz9s05CPxNFe3Il3ARkBwEl8GEEixgvAtc+Sgs4106246vP5VUnG2LSV0aMm46
q60iBxprGJrSpE4HsiZM6BmBwbrWsMlqujTbP2PfGbk2Mj1x0uCOA7xO+8ylbahY
HIfFJnQ6uyJxSpROVOy8Qqj1bmqbXMhIWq8sWPppOnfl+spl+V3r4LrWCmSKR86j
x5IB/hLyIjTr/lL9eXQs1y2crzJW0QLB5s3My43ypzR+ugwdF865q82YWQPHvHNh
IkZTA9HFJS1QuULqVOMcn99ExBPjYqhAia1WgIk+hEDsVaJE+Uo8z7ZOPlQTqUik
jHOetTiAaW4N8yik2luanyJ09E7uL8F0oHL1KOH6jeNnhQ3tdSmf0x8zM+6as+EQ
ytupM35mOXhPWYq4+8WgA0JY0YOJxOs7OU9s6c+mxXyNQnO9YZuZ/+DYuHyrj8Am
BUQoTRPlGGFHSr7gaoS5VLSYOgPQ6HXDHM1cOybYsUNfR387/cDo6kCGbXK6aVNV
TJ8nA8wXGDG7i7AeJ1D+Ch4QWvDsvSU8NIQNmiZZOMEQwIvkuBiPB2WIru7ic4Py
QFamMaAIPpt5nBx8qo4UBJvLtLR6CPZDItgnyXWjuJHX9zcKcmxnjuICdT+/ZxgM
J6vGUttIDW/WJRitRiB+7bUNzPwQJdPU7e2C+XOvKfyu9JxwnzySnipRL5W/8EZq
wwl7BjdFYE1gZ3Kef7FpZAyx5W0BlMfUScaaGudzrGU11WD66uL3tplnFCD464gh
8PndmHXK9gImJW7GohLSRc+VWVait8lrRiHoY59C+4ryM6nw7AvXeEWVDcfeDWqk
UfOgzV9XZLyChidRsCtTEK7en1VNitjJC08FjirQcbYlIAP2bT4WFYZ+ddC6TTxN
5LVe23TuVL2VMBNDmwNm8a1rn6ii+G2p4XqqwtZh49OpFkszAIjXyVv3UIDdyFZD
0xPljMxQc3LHm2v1nG+iRYFUrT+qDFArmzcd60+HvmIJnpioeo5Sl6JRU+v/56yk
RwzfEohB1mX+DgZoVG24/azobBXWTnVHltmSx2UkYyXOsZPWLJasXU2C/B7P9T/P
a7ghcgHykjCUOIpAnXiD2YE0dMyVM/RcFw/7cniz8gys+I5BkX355QgPN7IxkK6i
ytiyyUgs5su+5fZ2t3NigUW4vtW9o1dYESJJLUpKLr8I2TcKYe7DMvagPwYOIZWY
b3rYKJH+9ZMGX7XvLPwT1xF362phthu1epb4EP8vcz9xRXStFjSFJSruwNDRgL//
Xgzc/m7OXVfgeO91x6dYqqkq6HCevnEqHk1DzflA3Jf+//C5+N7rhSm9Yr9qLTa1
AGj9GtQDuiBXQWBNZTdms8bBrHLoqVT8vXohVNAsy+iwEQkYtDEbKjCc6huShBSf
yEhh+6EymBCjdviUyKUKB2TwTi47lZ5RqQJ3qoyqNmiHwBqokFn5jpa6XP89mE+4
J9xPhdz/8fC6S/kHYPrfvm7l8v+QeKA9A3wt/k1iomnUCayYMS0qS+hZ0qJ9BCad
inlcU0KV9wAqE51Hla3QTs7BCbDFxv/d2F5OhO9CsrywJKHMacmbYjY3KyV5jtJo
LNRgAM3psqLVRvln1GnVzwpeYBgrVkzwghlgYhu0XDGZakuYOV78GBiMLsOR+pRL
tnShJkHsQf965Qs3UoP34KO/nC6AmO1N1UYGitidMj+msJVUwwyKeW67I3RZiB6V
Kg/SUlznFdBt/HqkuPZnOEPEHmsvzKMrhbri3qVbFj4t9fn5OrrtHiiYx3yYkxRu
KuZXLMIIzzPVDSCXaYoHVExeoTHs9Kl2FinJ49IYHYv7fykJi0aQplUTVXHXqM5Q
W+r0QDDxxxHhsmI6X0V7TR7Wbn2t2lBTNQEDY091IceBmXnvtHX+r7NI8glu26Z6
O3ey/TA7ch1Zlwc4KLMhCtiZ7QVIQXVb4+nyOV5+jaF7Ibrmg11BEDwOYT0zP7gF
tr1VDOz9KoHuEsyO9tDbak3sDp+63F3vcyosqp6BvP6ERUih/SRHeRd1RCIZt7Xn
ZpXpLlXHev1+TSI5mqTdEhxmB5l1nBkXuBc3oRVx+GnlqZ/pR8nmknoNb1U6IAA5
1qymCH50tnbzOgsE3DiX02yJ12ZBowDV2sSk6Xu8tAKLJhKP5FYU4+KHKkxNRuss
h1JimFs78lD5unthTMHUGAVfW2K0tjcCqQbnx/SLVE7sY6vzP+e57CS0ZbZB8zcW
94f47+tWGJeFwpYBUzvcaNokWsNO7Gdxw1X+opoM1v+GeM3wUo36HwyWr5ltrUrE
G0CvhKYM0Tn4BKqwfBebE+ZJMi+CjBvq2NtpXTdg1UCR8nyIWoozTnJ68JmTgRov
z4AutifJ7l/p8hYPaoLkDL1M32/3apulZldiLzgPFRFAN1uvrghAY/0bmXvruaw2
RFNFNrsQGFsma0Z/pwvrowk62Fv6hJ/S37MEp2kxyG4KPhBou8ESfBKUJwBesYro
zVgvKD30ISk8Apu1CuO45SzeQs9Qg2Wb8Vsj0WVAvFwSY6lm63MvRls0dqGfynDg
16sD12CK/yLHQizqgIar8k0TvdQviZ42qxeOLJQU/KzWjDwpCm/gbvDrL4eD9wYn
8hlgZOdT1l2//WWwWb73GiC1S2vsK/9hXLrU5dI/WF3wFc/lwWpb8ZxfxfsMRFx4
5vOJbSiE+ZerqZ5RkzbApIPtNP/leklekIUmtFCFmillO/B7B57zt2iXfw8dtLyA
ZISnu4fiQrYMO6oxXVhHDVGUxBEWA120VflAXXjTIXZaXi4u50riihP2T0heLSSJ
rixsxd7KDDwOp6NpCWH/YHN8VKWnMSMXHmxZrsZOz2glJX+gPkaI5zfGbhDLF4tK
dgAZJMlSjHNIVLbBzT8TeVbwaVXB8JgCDtragZrXTX04XYJK49QppVqMsemjHI4b
pdizHHlsIYewENw/QXWPnSYtqkspS0QNpXZKztPNTo5UR7Wkf4xmxQostj91w6ts
Iajh1gbPquotYhAd3+0GAePm4wLhQmTvy2qgaODMxKJVt2IHhItP1a9srBi4fU1z
taYShPXlcbPo1ePJThglAU/byjHT5r+ecdnA2WRxxvLfEZn07fk5NCn9kinxWBki
nF7RQnazGaqyAwRRIAXCkfXCuODXWFErzohgo4FdvlLbQkXyd0yTQA9oHaGJkSrr
aWIAPNewUAEUkuwKvCcUQi+aYYqHmsRK41TaTsShJ5vYPEgofo/vBe6yx44pTP+y
ujUwg6C8NhMLpBiMoOUUsn8qFnrP2T7btG2dplVas/z1EnAZ01U1GhBd+NGAAVu/
2S35rJ0d58e+vvXP8Nwfj0/DysfDdhCpCRVl2gGwYhPPbOsDaRRkanbMHXC4r8pA
buLb5uwHjD5FApbaVkjPAOMP+uOWtoQhhv1owBvz8QXuzwg++tU9hhwILU6TsORe
k1aFeUJjt00eYtRp8PVk9J3+8nwSCOte1jIovB1Jga9tpqtnpvYORDG5aKJsx3TS
ykTjA+v0xqRnRZZY0UOpNel0LczTyKLu0EeYvrqy1hu+loSf5ismej10Qk/nUTSC
rJD/ZcMZ/mHu6J8/LpVEE8VYxH7+/f84YHmC7aD3zhuWucPeQe+hfVDvr/XuuN9P
GMJK/bUt/sHjLEwLTDAhHSg7F0F4Gf1aDXNET4oerzilbofeCOaNhe06ypyyQkjr
FXiFXmeCs8j2apmja7F7mJZ9xvv4ZplkxYODxhyvvYP9K48YRLn1JhD2HLyPwX+V
uKYE34GI/YCzLJ1cpeW1GbbhyUlEZwL5tYjIWyQL100UvWTsAnBaSSW22EK6yFH0
/scmAgCULAYM/jVqIutDo6QGCTDdlKlNANAhpIcYJXMk1NnW8uMD7Sgwdor7gaDx
b58EkPuktbAU1lnSwa+NiSL0KGd7rsq7yidhgQ0hdzxUN+tBK8V9rzNpHJ7yEYYv
BjKTz1e0AtF5fiSuvRURSmHY6WWmQu0csSITA+00hxSPWlM15FggtDqacgQZzEK5
XZ2FcJW0J4ECgCjJZ0yMR34copF+lFYR0Lrp2avB16aMmfWFN+v4VodPyfaFxz10
//eLVmVP/WtwltHzbU+DDIFj/4mabQZNoCUYEyDB2M8rv7Xx4c9TneyWIGH6514v
3DEn17o+Ijaui+5Wb4Z0sJ3v5BS2gl9iQFgZHUlD65D1r8qIidW1+VT77z8ENpUf
De2umzAkgtMa5wrSlVRSFqxNHyXpvAXIAeXfrx/bhWJS5wqPjdCfOWXTHs8bS56j
MsqVALI2ZG+gOdKz9ddC7KqFESteXPScClGkcKYOldqtB4YBKpbHyB6gyID0o9MW
iUFJD7v+pJu0mzcTiOdwY+2RbEB6e+QgVR6uUySDh81sg5RDfD9pCFq1bcHI9S5U
ZXZt4/t3pv7+o7BA+EEfjSOrzZflTDHfZuJpipXstf0FVr+JE8pWhvt18/HdH1ot
SMXKhbphuQDwQsobBMea6WSlqaqwvk8BNkySNMoizr3aZCoCvz5w3WLL6tmd7Wtx
v98j4mAi5+Ujhuztob87OMzwYa9irQzHSZIRldYAADW54J4F9HhavZh8NAgmbJzV
jQkKGdjNe4zoKPH0BacuQYDnLVO2sCEPVurSikrNCnFjF+//hGOT9KBXpRNmQG+k
H8wdkvkIWfPyWUmLSS+dngWDc5lweSw0k5BdKjI2rk15tItJDy18N2WvzeCJ1BoL
6MEM226g0nEfCPR8phZQ16AmtqrQt3sl4hYQTJ6d1IFq9xGNBccx7zsVB9qyRylz
DB4KViJTjmdDvpf1uthtgyXEN8BGvNhf/i6Eq05WFo8LQCA1MWXthDqTp2XKjycI
IohkofekSwq8ZF4SUOvNPYE93UEowpSeRMUpOcq4GTy0IfA5+OwP+68+/X8DZRPl
2vg7NL98avcWZ3UBxtnn9iMHeABrXvImb1HM8V4U64ZBWGbfP8dmWElN0hXrDuR6
sIjcxAI3NSNDpExLCZWZLpfTFeWcyO9LF1CrJ8zV0d8bkHS0RFaZ/zLSkxN45geG
/gUB6A5ifyHj9XrDPjIjVuvORQYtUUHtizN00jRvC4pDUcizL/Y+v+jxN+0AU5+Z
suy3bDX4r0370f2Y3Bxt3XRj5EMfrAr245fyLFvmq3uB4EXM2GjST/w76F/1Nz9+
d+qiLOWA6Ch1d8r+PItCPDdreQYMDylpeOTVOEoT5ZSmEU6b80FipB6Yf7yzbpTt
Zqe0i/+I77zgsstag7SQm0sLx+69koCLr3tS5V5G/HSM+CdpTBjMh3ZoDm3uvccb
G8clkVMpHzgMOQhhUN1guru+9frl7nNH8ibK/YSWQhdkN3k8C8AEtLb+XmvaBtGw
lJAyvQ6EvKjmj/untjvdqaSrnYZYVs87iGufT2CcWwCT9zZb08x/hCj5Gxy98RpU
XlMYC1zvkxFsjNckWXhkCpMdccAzE+VUkz4zisALGHPmF8w48kBvLF7vk4ZZAzbx
PibcFWYB+VuWYbl4vx++OeAIi+4wYPJZ64EICOmHgj85YXgzo78ymVIJhlt/Sq2B
j3uoyKB8VplYac5QhAm9AdJfJr/Q9dAMLal3H69pTeYbJe4dU/zTzDUMFJgLsxIE
Rt6Fry0/7rcfx6b4v2b3fpMn7mh3Xqmrce1kAgZByM1pquShlDuvLzTscnL491t7
DSiKo0NONwWjNC1xPW/IWm4Iq0rtGbxRv81Ox+XUrPKcueqY+LyHGOuJ4UMVKTwQ
nTbeaEKD/Fu1sasT5Qddy+vNLj6jDR9bdOmCQ2+JyBb6B2b1C8yE/2R9w1acVrXr
wfBsSemMWTmJI5Mq+VYoCuxMkPy+vwvImkpnZcLCjd+DhYQfK+c6U7ehRLdvaIyw
JSw+LcvYh8B4ALto3U/MjtNwLBLFoRDDSPaO4qWxwL3CDTDOD9sdLi6u8Ookq+o1
fImYhB3qQLwAQ9FMGVljcQLwi9yrSjSfYrN3dtgE3tpnQVy4emqnWbHkK5lqxI1+
GkLXluIvUde6HFFeOJVWZJzjGy6IC2Mf6rlacymgkBOQxQeRkGn+rwmZTlr6YXUH
OG/H+cz3V7K0XMe1jUQHWTTX2BSMG8HdzETst1GFX1nGbic8hEt52vaTLmCHfK3r
mC+DT6YLcUY15bs5pQlQgOca5Mf2TTndF1YoB4pWc8+bYsk3a/c5xdX43qKbpa7E
qV9Bn4LCsD2vGImcnkWpEdqFkLu1Uv4F5NqS4S+rm9e112O3+LdMhoc3EH9CLsi4
M1a2fWY6+vNukV3tp2Y3c4Wu0XgFLMcxWGouZWXKrSJ51CIxwFIza/sJq/+uqccR
ZMnxKSKVmeFPQ+rSF5J12GH1tsI8LEiUIi/71etH5ltWaHtAghtPXN8jwVx0xK5M
D3LcodNFlcAVdDNU/FKhEDMECZo6VAncsQRsztBb/AHQvwaD593xcxabpOgros85
Z5jyA7UxI6uVhtXqcIG9ULVnldC14h+QUIVUmcJ6DQwXdK4bBnQJx9Hx2HANuRlo
uOtVmBLw1/ClByMDWzFkJqdTQ2X+0I1yC4/5xbuIaYjEpEJs0rk7Go+JSswLEH7V
gsaxpwBedGTEWPeI4JKey10GhEROhHazvoPtNx9NhFnyQkGIAJ9AkiiD6w5Mvsd6
RJ5fybzc1d3fUKxNeEy5erxuWfu7e9K1KN0xr/HyzDDABi3UIb5M7bsrQJbdtnEk
xjwTyLTMw6iYmW9eH5CRTRItbt9nTtCu0cZ9VrM23wpZF7PGPEFcvewwKoTNVDhc
8ZThBZ0907B4CIdS+b1R6AxUp3CwgUeZojZxDrWEHPEzdaikSeyGW5oPG2d6Ti5B
9Urb3wPUHmXfdX1yai3lsLRHL1ihEciaLqYHpdMJyivPwC1HIuiY5CpLu0QaKyzv
Z9xY/vMefm36L3aSUwRamTqURr/XfKbkPoAny89mM2Al0XD6DeOXGJFT2srglT5U
1IgN6IqwAkvPKnAFbLLvQZxqHvqcU6M+X3pElsLzHSZWeao52kan+chudrjrdCGn
E0ZQkfsnYDSsjQ5uTuFdAHuiH3Hx9mz4L8xJ1SMQmsi+sZM7kCsBy8hG5hZIp2uC
1+cOTaVRWEpbsoqjU+S6LzwxHC94HWhsd0JMgA5eDmm+4g4oEYqYf3IXu6OE7QJY
6PIPNV6VhVdELBPMQ1PVQXr9cefPzp9PUUIsL19xfaKLILNqzfFiz7emZWIk5wQj
s7Dhmd6SJ35x2wUZ3wdZO5V6ynT8jjss7TB5AmTm84V4ev6Gl0ZmTsfVnvSqTI/R
ZhuSMcECTPblXz+vfacXc8i0eRFp1aB7EjXb93mRF9EPJGtf73S8rlF7aHzzq0iP
sX1HrlLdHOGkrhfgNshTmYjhh0MxxfbyGQnc+mOxpyySHQ0Uqz/yoBp7CWPBMhpY
/tfrDfapqjVBJ9Yt+qhvKhoqyxhqBOUjEbLbkjQeC11WyDCpNxJWKQbuNKGAQQK/
QFIv3baHMmkh5fz6zlk9MsAHKzF+F8tYfilKmBQ56EHncjV74EQr66zhR35eZhfT
Te9VtLzDVdVgmaoqXaPu9ncg/z+D8vy1VltdVDDH8DPUXEu/Q4aq4y68hEqoaH5h
K8vkhkbEz5fELpVe9q7uan86sEupgO6dPtHjWseiX+xnlwaKstrogPemqUTc1r3f
4/ZsSYCKfnPS61TYOiZwEN3wwKw88U+LhjhxLNMEYFeL4D3soBOfUsrOzd9gCDWL
EuMED2Mi8p1nK/6Rzai6MILrAtW+9R8KMCAk6VS5WytxhWsjeqOAQGVn4Bbjfcv8
KoOrFcCOdGHMxZGZnBzlIX1ZC/6pftOzXLMFF0V0/N3ge2LkI6mOQ4dVQaC58Tc7
NcztEuQKY1JPbMSLQdt7Vn2ZoKxUR8mL9P9FOn+9ypqubfMadP/u5V/VdDnueKzy
JbrO8kK8BJTxkbY5OVmZcbAXJ/c6ZxU6zulgJlLZEMiKoCT/9wAYN4up+dL79XoO
A6olvHTmlK8+UyA02M1aQpbQMbxvLmYf0xcbeKUj4kRA9QB1EMV8dpj5uCRRrw31
UxLdeZcgzvCPIma7lTUAFRatnPbbuOB3bJKgLXWseUGU0Bb52/sPBFJ9PeSLxXwg
Zi0xSv9GLmG8gKd+J2weLz9dIQTbY5/4P+DsqNMa3HIZ7Dv/wtoZEBrEruHVzzmd
Wfu5Au4IY0LYD9npmHccggmskrMJymPdQwntE2Enq2eV2KL0geqEtkp2qSKDl5LZ
SH+fijcWBsh/yPsnuCVenIRK0CeLxyUCCFsSgF1mr4jLSlLnjtZ25lf4vHmShZsO
iV6WMGNC41UW1ckzcslv2Upg4Eq4Yupv4DlODTr/58qWWdfphekada0SnKaA9Md/
4SuwV5jKghTNHrSkOoAsibh3G+KfIJ8h7XN7axAIM0jP8Z/se1VYd5+QPcbuWJE3
RdsiPJEolEjibRpD0I1xFqyrdPkvexTh3Vz2QKMIMn5asNkGv57857Jcuktv7lzB
4aahcpC03cOnGGonP4bxDLAmYc/RbF+tsbxT6RyPp+pl+8r9ci11b5J6oCa74vlK
Va/vNdU6YNrMigr8KEwDQCxkL4o7TdKGlVk6k5YK7CAtQ1dlYUeW7wHJ7P42nAQy
stKgRgThWP9Ek+tlqW3ZrNOoBwBueQWEa1ZZuZJ9I5TlvOLpI7gr9DbYBC/F8HNh
YihkWjGbHcLbqdOgopWHTLzDH4P67Bu14I6rtp/zSVi2KgO4UMR39AxH8C1IrXke
WVp5xCxFBZNWWo8PV8HwgBliGeE+A4grkAvLM3l9cgK3wtlvsKHPGTBuOiUouO6U
oVhih1irdpsry6gPSCdlInMWn2S79knnX60STUN9ON6FQ+mJxlr7dVOhMxNIORBD
zCIDO810pRg7vYDlkV4GjVrzsmtHg0Q7nHw1qC4otmwy0MkEn0OM/HCk5hSHHlfv
/GBjw3sQ3FXMs5y4CH9iiD3IFTs6AFmrhv0+65M49PUXQSZrvFyWTFrxg0NNo34l
QeDlN7goryJYLfFuFU7NvShIWPc1bjtf/l9xH1mk/pcnU6vgXRKVPV211h3C4Tyn
JMLPnFDvxvAUQTsDvO6tfYZUdjWrWjvbU+uY3tPwoesiJhNv4zK9/TaoILfp8iv9
FrHulmHAo0IJVI2U0Llns/GjktK/OQAqJ2ooDAZRJ/G1/pMRq2kCyh6AB9oOgMv2
uD4SlaF+hgmUhhtMa5J6ARwUaF3lOAXZgxKaZN5MPp5TGhIxZ7i26rOiTM/2M2Gz
C9FUlPRDwQZKY7HZXwTMmfRa7/69Zqkone2IfgFL+sRrOWvoX40NIk4hBALgdpPj
p6REvIDdvdTHoN2KbQKkAQyig3IiVVaFN/Fd+rIFM+3Xp24OXyWAMw66b+CLpqNk
sfV+7uYt5s/o+DeIJZ2d6NMPlg0yXDxQq0SlAiEqEl5o38qxKAjm+mY+BT0aeRmT
Phur3HKsBOVwKcgl49YpBGcz9yjuJ9ER4NoLxTjdZrBQY/0ccle0iBUohndJs6b+
oIFkBT8BPN3rw4j1HUGB9HAMYiFBzwdWIS5PGd+q80EWSsW8N0VtWCmKb2hmTgKG
0nizeHU1iBDW8/acWC3ZfozAcBL0qkNwjNprmPSUs4JgXqDJN+gnKDSM+FU19oaF
19yMZS70NBXlYr3ZkVYI7JkCPTrwI9cQiRHXp8JfU15Se1/lAKzFyraAJkdfMqUp
gzKyqya1Wd1pknF5lCRXpp1ttc0ie691lQ3nqcpYRKF9oYuYM+6+9HnUPa4ISjVg
RtF02ne1DqKQdh1SRc2HRFd1xSeAI/j7qZM0RXeqqrmzRobuZD0F3MW77Mu6X04k
o/WrnBT2GOhs8SxhBVeIendAUs2B8wkwx04prZ9gRuvseQza2oPObpakNebCF4oO
1UyrJLfpMfX3P5YAztPBXQuFoJlNo91Sau3ADV/TaUQVDsKPUj8Dc4hht8tgP9aA
XZmAgwsspXQY7+P3Yxl1BIZxJmM2QUoVx21mfdvmTlWBoClbd+BtuhMnKZV1v6KC
OZgtfDTbDUWy/4K99g7aYeLnqg8qjTS3sbSa3RpT1KYTvqkFAIgQ2h85YxhCA4Od
Ar8mO2h0Zi7/zh/sNkK8KTamsp1i+o9FF8Bb/xGXPcBfbmc42u1cBt7Vq+quCwJV
uKn2Ju4sDmNUGM9D8552d8NWONXZZmscQVr/SZaBaqlVo5rnxJeyxHzgB1skCdCo
2Uykklf+99ek666mPrROU2sAguJC77dtiaCdmnxBRQ/RnZx458bZXi5+S2mfsE0U
WIYRpbgZxD/6QweCaZkM/+0RoPis4sBtz09PtT7oYcFOBrKoCN8uTSsLeRPxwaNe
bSr4vTYsgzvs7/5Ge9DQgMUc3v8KaLxjR2OjyMAugK/z3GFg1BSEbFBo+yLzGubD
ge5jfp48bSNZSvy8Js8inXP16XzdVTcNe1Ac7bcsLuDmPaJRCj+gVGyrK0QW/lXd
bTVKJyqUf1lDsdPhz/RkNyGzh7lLLYafTboZYP6Ydaw7yvmyBoS1DjdEtm7AteEX
ZKiSbsM75tNCMSC9ZvvoCbux++MjQclpDA6p0amHabRFqq9XGo8G1s+0aNEIf5BX
x1YWX9UMa4hGhUiKFAKGQa84iM9J+TW8lXlNP3tqGqo6Wk3fI0eEIwheOZ0RVBet
g0aTNA/80mKabWD0ydYmpZ/mjMUjlTvhzBFmo6VsBBGEF+rSM5PeGeKT6nggz5/M
KRaBO8M4yt5pvv20F76M12Ny2RfMGRbJc4pjGE64cyo1rp48/L/+JPm08y2Xawmw
FntA8FRdx0+drBHQkSdNWcOYYpDkygIy3oOEOtF+DgB9210zWNRW6QsuQexinDIQ
vJgwN92Cn521tERSvL5IZmCz04xQTEB4VyrrLOXpbBIDYvpDukeANFrgJejhUEt3
6sxKCOYXbtbIK15r166qxMcqKr4GpIt+hv+MkF5DdXss8z8T5Lg6gYbXz7wFsdCG
X1R2xGF00kqBi/xll+7dPDK+a7HoconN9MCsjFTYG+/l/TF6MXmRZgFT81EcSPpt
nXtnAU5IsImm0z9LgPRRWeUlySWmxbN0SuKrtuRh6X1RVQPngIHIVvjTrEGBOnQh
Dumah9RvaGdICXwzzM2eg6cceAcQ4sahHZ0d7j5brISnB/lxAM2T7FksXngkE/q9
Jz1WsgKzaJoc2FzrZblWBcB7/IwIG8htKsicu0UgLpYADSll2d+kOLNcFFO1I/Od
YEOFYmhTRThsPnBZrSXbWD5N6eKsaajkNueckwIH4wckUbQO2/FJqWKK8BiTUmfC
FQNS/FwkDu3OQiuWxkhcKKl+TPQ5q/twmzuPVCqD0t2//Pl0zQ74SW5gx/AVjbuI
a6BJL6iIDHPZ2QZtApT3NRwnLkCPUlo8xxAVdsVI10IHmkDaGLEQMNnBJ0M7TYvW
HT+/GqN6/pxiWkg1+A82Eft1G6kDuc2cgKdO76CbmuVqyKQq8q5MlUi3m2SfWkr4
nEhaC4ka0/nuaNWcrR3nd/ZqOZAnOHwwhwLa9NycWVQDr/BaRXy6KJBCEmOviMUA
Wji1QqN64LpdWtyUTf3+l9+aDuGBGS3wiJTfrkbP6gfq3Hp7+xMMRyX8yucMVGYM
TAv6xFweI8vlSbQ//snVNqj7agK6Vi5edaBi20+tUwbk7vQBu5gy5NHKH5m4aqjt
QQWuIfSDjvqk+FVhQCHgsY68X61jCS5CVNfoNLgpu54IfNdZDQOuamOL20J2dZ/K
bO15DZuE2/csTBApV5g/DHEX7cQIDHvP/xFlLRf6TZw9mO62tNZYkNbRHj2XTPqQ
KMxv6o2AHRnuHV3CVU4AYmEtqUX1FpiQya38AFPQWdVNrbsrQJLET25RGbWTcEVg
h0KWn96zDiofmBxFWlgO3CmJyTYWrO27nG4Gr0/2VXlr5EWUh97Zde+L7hrjWrZf
FonfSQ8pjTBH9DM1a0ix1o4qC2KqMsJcDJrLu7itexugPNBR4gly/BvxCnt+GHHi
albEy3geVQ0tv2nIRLUt2qbX6BjRdOUIXejBdSvH2Bam5OEv5KCvWBjmimOw4Kol
tj1sNG0CTkFkeJBBYvrsjBGiRRyst0+SWv7MOa3HkU5SFR+W2RJPP8pAp76ID45S
pWYHcXPoFbcDiKlfscaqQNqIOus8jRuc4L89rwEgjLobcYXQ3jo9eLdToOWKUbNz
lRmRciKLz3PnIqIgf9wSaT+p9PpDcKxTXPsy8dAcoy60gtDUv8g6dp7qFTKNogfh
j5Eh/sfiFX+JTMvfX8MdQcJUE3esa/RheeRcBBYGJ1SfOLib33KnEtLc5c9r1FmD
5zj3vXJ6AjIXSl0UH+FAdzULEysJZWrek8mxQIETYTHNUZrIThGfPnhnwMFqKcNJ
PEsGFtzG7w9Gk73vmXOFx7XWGZ5590KaFTiFoh3Qc9Ep3MUM25YTrtTAuZcKFpMx
kpTdT+W75lMFP24U0XNRKQUdlVkKzfXHXVxoDfiSOCG0FS+jFoLCKvcbjUSCIvV7
eKwMGtC6VlQjU9Yzq2kXU/Sw8NNXxfjbZzio0o2ZEcQm3nALQZZY7MY1sDQVONef
ZzNd2E7kmDVyF5LIEUTMJBc1HzmuQH16N3pBsmd5DhaFl3e2vqs0Pgz1g6mcA1ZL
6C9HwvG/J2sBGBJQr0hiVnoYs7IGrG4FA69edNAn1JeCOGKuToG3YldZ3oocz73Y
MHUVEW3pTBCq04UBbkqoxQ3+CKNRGnO3BQJMy4yih8tC0hq/7GbQ8YLLlb9VGwt8
D8eQHdNz778wxxXijvOn82ZejIC1+iWuM3zRumQX7dpyD0hWFhyBgeZ0IBOzimc+
Il3yWxAU9/dboRO+ueyLZ5nBnUn+POu5gv7rhG2g5+pvGSHB5xzwAc/Okdwj4Ajm
5eVZHSWKz92kp+OHArTnP9ZDedg4TiwWo3IdnKiaNbSk1WdWKDJ+8jbQ9Fbdw5M7
3FnqmgG5nrYJin0llBKSAqmeozRK6suDS7+gI/yTcy++DXXo07kEyClFQgFsSA7w
PGMmOyIahMBcnen64l33zh4mLa0gWcL2HdHf5bSkwTvSmCfNva0yfZr30rL6ty1P
oTzM0LKTwb+9ovBM2lWZGcFO3FAae/lG4VFfcvJeAKhXgI3ChGj/ft65TO2yUPqM
1W3Fb27c84B5ORf3ipTF4yWSBiXKZkvw8fyYk7SZylLUZKH/+ceVyfqGdQ+f0NPS
e+esKROZmvPG70zer+1F9Bzw2IVe14sgOVmqDVMnIQzSMSyZA4080iSHc6Ev8VXG
atgnZWveWvBZBrPxZqc0JTlxL9mOg5QT02I4/uuaznn1GXdUcmOpweXvknUQFLwI
HNXxtN7Egd8qkYqqjq1B5W8FAmDDyLUlRooyNX746Ut2cDAQj1AH/b7ugDRyFHs2
Gr+20ry2562W8THr5SdHN4U2OMiiLKSQVPEEmsUA7l/iqQs4f54hyGCTeSDOEaME
EeibiDCVk+eZJ94TabcjiToU7HfCZFWylk+2d6jNXfks90NatIzCMfWJHnLyNgQa
6iVYBbZvw1dW7o2hXXOo4WdO5OM7MSDmUe4ntYZOksOeveq0Oys1rAOJi8dIpA+M
cUoaUbI5p6hU4EmjO8qQAZOKxaz+5M7/WypeA50kZVivUEk0eK3AuwGlkpzWhBdc
2wikByx3BOS1g4Uofe7Cr9wviQugs+B9UxSh9kF4OwfdDNSI6JmlFTN7hLD4OBLL
Q2A22Vvp3hEr5UppG1nPgDbZ3F683SBzwQ7A2gBxhnHrDB4ThMQ0gL6MrmjP/Ffd
CyAvbhbUmrAV58JS/KgiKFqcZifgRrihSua5s1C1iAGxBdNzKamB2W+mM7VxFAPt
8Y5TR5rZBm8U+BZUrAJ2ZIvmNy2gTq2vAEVl4Px39CfYIb5pZVdug9gxN0e4kHGi
9XadhWwiwR29jM9vq8fjTqBjRXzKi1z797BLzqo2/VB6PwYe4E1yx07fZQPdVDG3
aPXHaHHyIfKsRQj02YbNn9bfViNKAEqraDBT5nevIgo+mH2Qvbbuj5ICn1AxIrJu
K7og9Wd80HNrMTjcqBUAyOr6h/wGrGciVGhIwlsU29TP4FjR+j2icySuIQmw9m8k
ETu08wF3QvG0bg6ZtnJijWT8fl0Uv1TbORhJ12y0hg8iUv2KFpaXj+2/rwiBl6jv
NDMaoEtoQI8/Fv38t+Z6DSIPYs5Xw6XfktbDtcG1JGot/vVJcT6cSjMqnmT4b6CJ
nTa6dXzRn+npZi8dPAESBfiLDuDee9sKsbFn662t2ch8e1xjA7RsSPVR0ztyeMSe
myMSQuBnYCWjSyQret3rzOlnPcu2Gl9xHHSSIHk3tYRJIGd1ZKXulrhn/oGTaQb8
hRAWmiTjTm72PonRsmDzDOetuWPu22AN/0wZGQo3WLAWdWlEQkS6xXg2dlpT/4Bm
lTpk5oZFva9geFK7AublxyTMjQ+5wINdqJOmT7UuEoBu7Q64NItTDzXdOYR0gvsR
dG4Cop3NBtvm6jbDJytN3VOC4DP3/B25GTPtvbIjldHJVOmGOxKQMTuFjBTTV6tn
7CwqTF+lrZ8Ld2x5y+krIwivYo6TK4zRqxQz68U0vVHoXOCpd7AO+YsjAvtzxwFN
gcHypzt8cZvvziOUTbK1CDBAN5CJAuNIZsyodZ4tThKUCW8hR8uJigGf9qi8yPqy
T53kZCQPQQm7Tc0/S8+R2sDhhUcS2Us4Q4WrO9G22+xrde+v6z38SNuIsjTA0Q+f
yp/Cn+s0DXhP/9NwEZWbtJ3GJ89F8OImDnnlCwRSzO3UxtWQX+aaBdSw8Ui5NIGW
C/SrpBstmp9r8BEEciHMmbcT+0xdhHXL7NK735rQnWVnVWHJ+0P8Aj4RKYDNKdaL
dSw1Bl48/+si/nF2JpDkxyUbHJBkgyXT5h1kbKcxPreslsR5JONr/tlmkhfKlRD6
RBBIGNVi35Uh0Xs8jFexZgLfLkupEuZSOyPCt10QYIJkd9uMptLZWt+JEAwrMLt+
jE4oKS7LicCX9pXJfM0e8Xbg14mEzzuJ33FtwlII2vmotJL1pRhMuuWpqKe7U/4q
xxoy2+Kom3pftt+5JWEMQ5lEHafn4YLvzDvGVGuXy6LMiPZo2QZdrFspdv7dXJeZ
NQFudK2nr8qmWG2h+0K5OmZKZOr5g+h0hwZdjZwz7Ef9qY5/3ZjLLVN6/sDIIhiE
BAK3b95igVm/BOIOqjhg34+l6IlnHSIsjZzpx2SlRRFbscrs+Z3Hg98A3i6xaVsG
EVFKrUHfavk+h7tGhPDMtKMvFWiVNDXa+7/4NW1BB9rFXPbQmwxMW8Z1wFzc7M6C
l3Tk5YLu2O2sOj2iD0CK7mEHzDjDmFqDLu/5kRXrEPr/uIDTqm3+iepETgwhC1Fn
MfhnYLtfFupeG1eM+5tvCS/2GnxWzg0U5WjXZjX8TpJz3By6/mZVdijlMegaEDpQ
6BMgz5KYXJZ6htN5Wr2QCsR67ZcSizS4LL6XGBni65GcjPttgJK+pAyMHzdVnNF7
lKr/Otn9aFCPIvkajSA5QpuSdosqZjW0OPhM4F1B/00m1zGtKOuUOVcLDvBamtMz
G/qieII1k7imUeOuzrbyk1X0JygHUKvFvOsLvRnmHEJORbGXDK6VWUa1Cwbrgd8v
zAlCHlEnkIEuuMcFVVnQXqDX8iKQQjV9fR04Wm9ZjR84EyjclG9Fcxh4gbBkFkBD
w4DNCAvcfFDgc+JKgCr1O89yOPCzAdTGPA67Hr+7bHjZSgV1yr/k6OdGzZvpaKsh
v3MkvO3DtX4hd2a/xO9W5noIjP276gfGA7AH6aoU0IPWKK3WZS15t3FGVIyitBNv
LCBcl0dPk7IGUu0yPG+vtAWR89KozLpWxhsIxie+0LRuQquZO9wW9Ejs2+p8taGq
DGnnY12o9QaJAPkqzIOdU9Qm5bfSBivCWJTh/1Anw20aPLSk1ENreq0jnBXrjily
rGhGqwG7bH7Y5tvh9fB88mF8KyS+eifxZSvpPjrrDPGLR4MDD70fvbPhXqsvGR50
0b0qYuzIlgkEgnAqzWW4OK/vZ5DpcJ6vylC05+xvHhATp8qHdLmevMxFiZKGWk1J
oK/0vQ5rGV3jPeew8NWBmMXDLj+AAZsvj+x9rE0ppF7Jl1zITrWnlYF/G0dRXaXg
3oTB4gMpvd3ziZKcXr2DdiSSd0rJV2a6U8Yi0EkEojKgKW6Y/3ALPwswxXOulYZY
7FGzQYPKny1Z+UQzcEcIUy2L47KTPF9ioS/ldfD1y0SXRNUgE3+8+NzfwfeQ3tJ1
udvIWe1eNgMpcW0LN9K8coxD3V1kjyhXxCjL4w5b4FgaL0IDbSgveNwM8U/jTr7v
R/WE42AYtj+1CNpdJFmnhy/IhZDfpQtZ7F4mYtqc+SR2khSXaBQe7Ql7kgRFBNof
dyBsmHL+J/YFDmTDal5STvWzEpHY46NlvBZtdEALvmg1ulCwWA3Y4LZQQ+pxP7B1
Jo5eIlaYi0bgQUJLXstRiQBGdVqzUksu/1KGclMycktrA5apWb2aP+M04RngVqoD
C0M+s0WyQhTDNnbN5cKBF2Ie81XtcKJkS+eAl+X8WjySiczLnV01m+Lbb2J/2RQd
CuXGh0rK5KjgfYH3hLM2JoZOAbGffHL4qVK4kjyIUkbOkagcehm2gPLG3CsYKx0c
jzfV0BNyRRzXo3RzQFttgStAGyxF10XtKL6AoUx3o0Ao7mpbbeJW9MEF0ZuLE5Ge
jP50N7RVloUFdRXjlxufSq3evLz6dCW6Hdy3gHpzusz7oqddKEF8srKSCIf/xSKl
MQgvG7oFlUhlXyzww06e0AT+OxUIViHbNlrr/8Uwy5j4cDK1y32CRhZ1rIqq2r4P
k9DrgTK6QPdIY253t2XZTaGVnPrAc6PrWGowuPkjUHU+wJ3qX76zEMJzbBt9CW4r
dG5BjKkQER+Yjc4cR2jn0ejuTfXVbAE+j0pzMD3zEWTIjGZp8Hf0nerGieYcM9YM
2UAaS/fmyy1NPyzq+Q2b18NIYTG8WTHXqC2nYURSsDmAsmW5I6B8k4JHUcIAvSbx
q2SxJweWeGnW1AXY9Xa/oMS8t5tgZDa1kNckxFUMFakpHd3TPi/ayqswccm6S9v1
CQMWl+bfOVpSqdW+BA0CdGqjblivUV2oCAtJgJJ9jYuOCn9fblrnO8n5EIA1QP/0
MittCa6s2NDmmXnzu+y6TdWLOwjf+2Yiup7BQsLjwsXiR767dx6YCCJU41Plf/wW
7fTxEHymbWe8T7QhXasLQ76y1dEjS3V8WlSl4JEW2h9Hm/pw8aBg9R/JMsvgWmrU
QO0yJXnjJDwE3bxsMTu5anphFzTQ0ZNcUeJ4QCzPmt2qG1S8bTx7+9SKJUeOylvY
G9/mwWfEp1pWoHhECHff8GluTpG8qXWJ9LZd0ISMM0PF6DvWrvK++P5zvKhWXzjk
tTE2Y4Zfk/8JDZhQt03lSbThjDaVS7iddFELzmPZtbJETHVnLsFbaJk8NIGmWyzB
4icV8kwP5PprwQRXsy7M5DRCdLWaBFzkT3zfaOfTkd1QB4hA+fFr0yJhsC8UUf83
P8TAo3p3Zhr8U/SQ7taDDjYJWr6ZAHrz0QvLtxOqzRPVi2HFK/BLVXXMbSFX3CsI
wv+1ClgFlVfzBnxPE0KZuYfgCD0NUI2MyXrZswei3KETSbzlucyePeKH0SK6s/Hq
vCKqmhGvUZ6w0FLFDCsaXrm/fb7HqksyraeiNr6ddMlYtgj3G6al1aT4WbfqUjmG
oT/xGhdXt+zmSBavQoJ1YdbCNHGI00A3YEvfzUU/N+hNT9mK/6SCsieFIOSGoNkV
hNEj9aP0YAx0UyghnVh0pkkPSRdCwxyoBf2+Fwd5usulSZxopbt2poPmOLOE6ci/
IqoB1c+BMP5+HBktUc1tfTw7LqGGR8IVe0rUPIoaZ1KBXgTD4TGYf1RVK+1r7pcn
llU5BGK04E1rSluAjLa3eeY8y9BkNE2Xp8DG5Q5STm66oPA3MUszyKPyrswq7vYG
EL1VzEKmmVWpaaU7GLvX1WRehT3ILn3GOmkOo1Ygz2D0TxLKTHEXUBdhAr8RtHfC
6rkV/3cPNX9uvxsq+xD/65gdR/8224Xc2URBz52xTz+Ie6YBUl+rAPFdSL+zIyj4
qHlkwJT1AEwkYXyWojw553j2JCvyAAM/INNdzXEHPWZ4Idd0oaNlGqIKp9/wpLBg
CVCHaELRoiGDoWMdCBT/F3chTtH5dWGVfwnJvd41wE21NzG2ZogBLpTvzV9jJLX1
QzhV58xh6DzqkLF8T3NwCHEEB+6JGzernpBgEZvM4iUkG0TriseE9w2yN5kIYEig
cm+BndKokECPIvHi5aE5McduTG5Net/GsWAgyhBluF+iTQJ7vp37agwhD7sX6Y2h
5yWFEPeXqrzcwcTUwYXewBiCK1ZosZ1AjiN63IjnCh2QTdKos9O10G/3OuVf/i8W
cU5V/ElSc5Q1xo2ce0n1L8d2c1O0RJX2lkt9/+6QMD91DrpGHIy8RXl2kLHREdWM
g1OiYgVrq+Hxrn26NNM07MhVtt7UR/BiM7wmF1p8tl/RZcxDyDFV02Qp75zMBkZ4
lSiBs8TO01ZvAUyVOgf2eF4nFxfWdzt/V/fr8T3Knp3YJhOpO+AXEMmovb0kBV4J
LboHQTRCYWNeYeYFHfyRJ4eOjF1/B/7E4X8tXc7tne17RYmvJH1lmEmylCh7nV4M
u9j/pFY/yRUmCZqTq00qkX3SvOJ4uVPxf4dIgvdQrI5Rf1i66YboqLkdFRgNSwxc
WZm1Pd0chZGkE1QrNUq9Up8tdAcOg2hITH+ntc4w3JKbkbtq7CmTVl+cqKno2FTH
8FxA0E3tWQpnB07ekzMACfbD4ZXTapCgncCZraTJnHn6sjthJAbkjUNhXFevLZPc
LnEO45NpigNhS1pw1nQW4WAmvTdnnJs9GYJQNy24vsGuG0sJYxjU+2qqtTBI4+dc
wOTNprXK9l6JsKI3xeo+/Sz9m1KGeFJy6vHJPAGQ7H3UfiD4NAgfUzrU6RMkMUNL
GAIMOASH0/fkR0G1KOOPC+3PNNG5+TEnyb4jMfjyn319ZlHdjCzqM1gHZGQdPEty
CAlY3gVelawegq4oeHYmid/WO5Wf0+WPUjUmXuhJUXsnzEEcuB+5oe/MYkCOL9ZJ
e3O1BKMzh5G9UvkGiEpwqXrF1P9B06lyCC0AGsO1Q0Ct33CUg+ZUuBk256q/mOGl
4LgNy/R32ABc7Mq/yPR3T6HMwg7UDHYhByMfxVsUjjmo9ZmPuPva0qgboCdDBzFe
ga7uOPjqSDXh5fZydfpxcVfycRq6k08Gz8FIJ/n3eaeXJ7+bN2ykjCykELhJYZyS
YxiJtzFSjdKfKhCxCqQbCePMbimQFsNBUCdazKlDpd2jpfSsNuR2BUUufnfaZGxK
SJ7JLcLOe6XiAzFtuH1SDSplPjMVh0gd10C1OhfutT/eGe/q28u8JB1xyaiXYUBH
ocxThFthl7C/HbU8EvPRfKyiC9cl5s3dAWhwAiqPVm9+fBszWS56QWYhPtNWg/b2
L6rq+PjP3ZjYTmNWdW5anc63qwzZybWDaX4C1+r+aCglC5jE96xUwdGrR2mamf7m
j+YQ/z0MITWG8cx7h9yzhAgFMJMmpzDz1Ydh0KUUrM4DLfnNYoJP+RBkgRd5rf8+
r3T2tyxQ/r8hZcdLcqxK/5h8SGP4Am8jqt4Z523YkcdUdeTmzz+O5p5VuN9N9BW9
wx77epzrbQ5goROY9hgp/LSCUObcdhN1nApLcRsIJWgMWn2bSF8lNkwKPZRpa27y
vfUVJrN8jg8zWI4f4KuNBYgzafiqrNOjRfDOEJDe/DCxAifwHjxwJ+e6oOcRu0EO
xGl4Rdd8rN9L1vlyR6N0zu4SaRcywT5XKn5zZXGh4Du583uS5KyHtZIr8zOYKa8z
SP66WQWTl6TGJBWokLlNNtAwDshzfDq+npFn4bTQ5o/oLx7Khu4RGaZBdFZSDQcf
sLsa1qEG4vcfvuUkawOG2w9aXnqcdUzP8H884R6ToDv9JX8xV8bSr2c8BJw2Mmrl
Az733w9M/X64E6uwGecuXFDNiCsPdVEm67kM3R1mqJY6R7U/JDPHn/z6ZJprQLUw
lr1rWXb9FHKGlpV0nRJ3ZmPV0iQZKt9o1N0f16bAssB+3e6M6yOMBiQUT7ebRgB6
WVNGWydwOSURw/rYR7kYf+VgdHkxlVyZnQA8D7EizcUbCLTYhoTbQ5Lhgob5YBcs
FurraGZGV3m2GVRuiuOLFKWKK2VP3JEuRIVaDaudF1TrHk/sWLp1OzMSg6sKLRWH
GzVIVqhRxFPDY2L7fhRpgAgcCOHGOMrvoyiuQTs5GHcrXxbO/lIyG77ATC2d1WxP
+a9Yi1qEBJ+/AJCJkDWSXrvbeRNfhA8030t77XgzkCoEEi3CbhYiTSZ5Ur+ZNrWY
E6AMS13dv2qcCEd0rbUwqfBroWduHuOra96+jWQvXKC36SjV+oJVT4sw0xZGfvK8
4EsfBKJ54vbYY/SHb6WvuD2XC884dXf8N93hTIDzkv1LmvX1ZEXFK5RuMR+N6bKg
XmGHsmTNES6qildnVrn6IvVpdGkNUHa4mRq7I2gxlgX2Mq8HynxREfwnq00Q/tVJ
5HVpHus3j38joo5+f1TulrZq49kdv+TN/Ev4ZTSRummuCnhSss1+Iz1+fJVKJ3g8
QfJmh9CJs2jNOM3AwD1LxYHXS1vIJKoAmObvGqQ0RhV1xUNgP4ESvDTSnwX5Is1N
RXRZgUy8v2x2cmQIL8mEBVyj9RI3GPIGfWGNp3OQ+jlYDnLQ0xX7RNUhOgOPGIxF
+gW/3BJHG4D6fT0NH5Aa/HPRxkwV6xZfGO3vkqhGXYS8yeJaL2RbrtL+X/Z1H5dC
D7nJQknkZ63zUNB90fDFYx4If1P2ihhSaobx/i7BI5wxYl/ApYHvhlmNILgaYHtg
b3gtKiBAQ6L+yQ507xDyteKdSziyHLNczTE3Xy/3Kh9EkRCEp3fVqxdPHgsvFz+L
YiJY8uWIX+4hhbpsUf3+KkEOcZvgP11mMWZyg2JdCGcAx7jr09aHFg2suA89mIdj
pEHja2ctCc7az+JfFet6FDjxyjPqDqIKJbg7cVHip3xsGWxorqXapaB8cCg+Cbyq
psyvo7Qwr+jiKH7tWmrjzR0bd9gc6GK4+Jb4v7u6tPm2llBWT0urf4c1v9iIopq5
7cbYJxsc3wYaZfofkp4/denZS8qrV7VAe55WNEPlU4239D1xYzg5BTgK+0NTlS0Y
ps4X/pQ2pIz0DUrP9m+okLwngWcDvdgSyAcK7isLJwaAvMzff4dlfAEqEMU+kHjH
VLaFx80emZSjB4YdbLGFFPKmsVhw72F+wahFyMCmhB84DdDx1Dhz0I+9mSRC8K4W
1bwqqPvtDXma77T52xtza1KwHYKYfdxLLZEZhq0S0SIkaLkVPJaqO5/e7dJWtO6o
7XDwBU+ujam7Pke0j3CeE1VHk8OkqS7HAh28HFR9wg3UaiXWH1yNULbBYmqqqzsg
k7w8MkvXUZSpIZIJetarj9yNKPalDcT2WHWJZ9h7kTx6F3uv4RTVpPNwyjkOiARL
z23SgGO3fNMrVlZ5W8Me2W4gQG9ztG8jskUzIkPEXPVMkoaNQFSsL+4+6MfGZ5rt
zRcQ9BL09IPaeUctU7f4zDcuL0tlty+nk5rlLm31YsMXwZs6J//N5rdNACUAxl5v
3+PnkiRsY3cKoFnKuFo6jAsUStIQ57vyprI7CigKXBQBNzjjhvKjW2Cwte4to+By
IDEozL85LWfOEZk2J3bXBYGHLseLvEZIMetU3hAI7t/eB/8VBET8RfHnvQM92TBn
SlUTbXeK+Wq/G4IvkWmzGxvhq4qOQ/efKhZiyT0m6PfRTyoFZ/mMlyaHn6R8Kndp
zkXJV25MUj++pLbG0NKkkYfxuO2vN8L4bvPiiS0iaF+qlgq5Asp9cGDO4ZBi37fX
I1MV2ZrwkB/uatKypA7UBQxQhSJ8QcWWFkRN38ogzyJSjgjD1lL5MuRWzyZm5Gdk
itdyqVnoPR1N1IkRgpZIuyljpRY/xgN0ZXUcfF0Wg2TUgWB/HIg76A0rpxd/RPp3
1S94HBfyRxGH6tWMD2FS+JLTYm4+ss7VQYtAF0uabo+CeNvB0eIEAHB620rEWHJs
Zc3qfWESWFDJsEXdK9x/FK9us1gZ8XMop5fcSKSpRlnvLnaDdewJGUejcxpvFl0U
HwcyML3665NgjxyNZ+7H7WwNqxeifDyt/N2uatG5vfbQQb+xJ0Y9HuEiRRyPunbd
WgTjBmmB0c3BPiq0NQ7KDKjFhkBeixK+YEQrRlbTLQDs/0uyaI40kVJZtSjViD8t
OtVQH1zBGUw7dfk4tcq+cLduIyzmPgKGzLSP/I6mbbLsMM0PlaVZl9UCjhU3/5KI
uPbYZ0+jQegq3pyR1TaQ0BI4SfLKmjw96y82jZVgZnqD4geS5lNKHl95mr5mGLNL
HJHYPLYzldbp13H1rs2q6PIqsW1v5XkGv2XtvX2dwT/9YPLz6NRkwqjvZdH2ptBS
4AWy3MFRSApQkvmuh+7WU5Q4LXmy3f69moRlXoe2NIGyp+rBjKK0Gbuj9FtzngWb
Q3S0fXAP53sFmzgkac6OL5SrPQYsR3qveZ12jX/uEhcTfawRFaS3eiA+LuBJz2dN
CbEKs/uV4PPxiipL9EEH+vwAz8i6ulqO2waSyi082suRVQmhJXhXHxlCNMdqYEXG
8csF3H1VANQ6n/+r5Y7RQK3Cns41AUmMc7h6HO3zUzsyY0YTMF0MJe+IY80f46Zw
Yi6uYxU1fbIRjLdSwLxxi4cwaU8dBFChypIOJZvwS/qgAHiyN/RzqWNOhxrjWvzP
et85iREpBFpVwG1VXZZgbJCZcr3Kf3NTxpPmLM0V6zH1KYUfdqp+/pW7suQHGeY0
ejo202dvR5zqwvZgq+RYYQJLgcOH5WU+gGg1qlgcW/0PGtcVm230Ux4oY9LE48eh
Qm9PHGCqMn9eJ8yReq3PH0unzUZGBew5VngJaaJvDeR2A7xurxmga1t4RvFGHT/3
iNw7Ua1+ihYfqGBVZh6ZFqagPPbNAIYSPdOST2XmyrQLTkCYGrtdzDTc/Cp/OLp9
O0QVNzz1iEVP1ntk+gp+RMc9c3CgYumlKyNF4Uo6Ra7wZp7MuZ/AVKAzHF8hUlXI
JiSDwKiAFoiTYJkl28zVJiuFGFO+XFgpWZTfoIF2B0hLwa+yXbExCgHOgK69Ob9G
NqmFr4Q+52+QcjQTaing8/ILCw21Kk1p9T4lV7eIjq0z3VBrjV/MAb9eFa3avGdq
p0qZGkLKLu7q5JfEELntYtH6MXD6ARvOGOtqZlPM0/Ytko2hapQofdGbbz+0KqwY
R8MmSgW2yb1mxol6KksYSRh2e+23EcB1vqU1anJa80xhENwoW8E75K3QFmgfHLgu
usmf3IRbvC328CfVZIXUgk9WtSrStyly6MROJMoTDcLhkadSD+m9h9hA9Q8ZWGWZ
mCOf2ekeVGO4QoThpFt8RjP6UD8ZK3UdgcQEVnDPer1NPL5UbrXo0yeWxFtUgcWV
s0DPyVGNOVklBYUZumO0KCrIkJjn5nc8hiJPbMSyJ3og6tRAkZw4RVI3EaBwvG0O
CwPF0DPgX4i5SLdBmnbd/VWS5XRYx8Cmc2iQwJ3Xu0DymkN0RBYctwtvENg+WZn/
WvH3DUM4U6fF+fYoCLtUgJlkk+VtfzHvk/31qUx0IQNPhiqvq9333ht1n95X+tAG
2sgo5WOxOfQTySLXlrywsYtz2u9i0NEvgbU1Qk8RPiuk/jdIMW90TS+HJdRfCtfH
YC5vVM/Ph9dNzfTBIx+zBZ1pjSHODovEA8WNZT/Tdg/Kf4GagLnv9phn1+/VVLQ5
B6nn/DmeGDnVjY0cul4mn3J/S6af6fH96W7JfTLGb/IsLWzM+gU5qnmDfaITtO6B
BaNrzOMT3AD659fI0soZZpm9EFbG3oBKhqAvxIw+Hce2qJu0V+X8p4Y34Cd4wdad
IDNlFHOMb77UhLy+RMyy9zeHdZjWK1GccpnE6j5ghm6yEh+ouFtZZc3RYEkEH6PG
rgbrT89jDrZggWG+yih2nfciLx6lw1vMc6K6kLSPfP7Gi0vCgEsBvZ5BgH7H/yzz
ElCAHX8Lq3hgywbfuu8S823MyJwjeoafx4Fvek4u4blx3lqgeXQbTdfiKLaG/0if
vg+oCtxpXvLbC8ZiNBT/eTh3cnd039n+d16PEUbSOme+l2335rs3L4IU+gnrFT4W
jC8ZUFpl/iom3c4gxc8h15YVuqvmzAfhp1470Qda9Ra9dMQObtE8+7/PZvHyWN4u
9QrdjZEXBSPoFYk4qz6ADHFuds4sD/xA/VC/RYNJ9sise4YyeHmw6ewktFwQD0Y9
RlJx9pspMAojB7CNl7GNlKiVF5wYOWbfocPwmNK4CKNIJAHm7SYOEfC7Qhb8Q1MI
JvzyGeRmP4+0tP4e8dtnu54nXOPtMTql+UAQW4JNRLPUuM8O+SryL1iWX7Itew9P
vLPKwK1TvITyrJbnAHn9tGO+2hj2YmTdXRAd2omc4KNB4xrrsCU+zdIonJcwv8Qu
sEJ2S4/H3mIgXH6M7/39M8s+gZyB71sxpWjvIQAac6HzX3bA+ErV2kuZBYpC7UPQ
qODANIfT2NqLBKsDj28rxaJgMotHuaxBhkTUUasTKq2AXoIYQEIvJi8dwwDqeEoh
HHoNDxcOqPiMWLNKgWkUhGd/oPFw42+MZAL5scv9+uJOLfoQaSSNVITI32eA7NQi
BRaEAXeZndLnMY0P2sRAhUBU1OqQCPQb5iNYHBUnqIaAeARrxB80qRbM9BEw7VaF
XRf1R7ILP30T30E5oC17Ee++ZPundtJGNuY389UHp8qHujmER5vP5F3DOjqbRJTE
kVNL8qyUupE3Kn8PLwJY93pr9maEoqof4xGdYjg39IJSrwu3JP8mxpXk08K/czqG
XTj+40CbO2vgMh4/PjeXamCfGrF8QSEof6ALXDkwbircLkGVxYI2ZFbwpozcDcyO
JyFGTOwAPAsIVC7welHYu//MDPibmWKUkvCCN6l6CtbeQPuGaiw3IOqkuc6R6tE3
8zPuCuz/a1TwcKStDtwmwYLa2iIGOyV7dHfDhNhm3EwoYwt/yRW9B7116QWUCrsg
KALcFFO/HyPV+dTr012YVZWRzoS6H0TyZqYqAop3YJTIKjFaVZIiehz0UC/v3kUw
WSRoU9rYIOoW+wdfRunXUA69JdctCNkk12W2euGLaVw78oPzNNsTdt5xJu32Qf4/
7RqW4EDLSUVL+muP6hOtmrO97Adzn7OaMExJVBOu2R85dy7SPso8plCcu9kUrBxu
E7K8Hi5paQiQI3JLKroEau+Z2SNpeTePeDeYGC6PSx8aCPMfTT1E7mF4i9V5qnoW
tg2rSLgELwUi2/V7YORcVa8ezK/vFw4brNdxM5EB00byXxE8QvmrRFAAD7gkK+y2
uXUFAQN+EvPk7TgczCCXmOOfNYSoVTjlPWTT5hHeOUJy1loFPghq+obq7g0wHneE
HkJAEDL66poJGS1bixmPgQxuPU4UWOIqC//P0ogwFb7UtP5xOB5kapQy19qqbGUK
SK1arS8RCSX43VqzmgxTpAc/3gyJAG8ejOBNY/h5jKCuJx208aIT8qAuQ5y3nUsi
WlcwEDq3dxOU0/doc3DqCDpbpy1KXuHT88EJ98uylqlhFl5zhE/6cqLK052ij5/1
/2M4pZHZnCMpa4KWpzVENhbC4j14PD8mbo/uBoSbpo4L6zXlWvaMUQPy/YDd23xX
D1/uzLKSlFRijHvpQnD2Hs/VXPw9unjlBPRTul2JecnDBVyOCwhtl+gcd7yXDq/t
jPruH+gwTozbCfKsGa1K8bl0h6Aq0K7temDXjjAffLVno3tI2oIMKCtLV6feRBUF
H9sdF7soRas1fE7MXE7/6IRmmPr3MojMcbG5H3QltzP78IgT4Ofq7ICkdGKOugum
NlGi2fhzlxE/uwv/R+PlmyWvKuvGlN1u7zU2mS0QNvL2BKXLV7UOs4JddR54cy5g
YElGsXYImdxMTufhkn7IGccz2qhBemFdYOQ4qxR7KFlS5c1lx6SxEC6fh2UP7ZR6
fK1EHvjRdHPZGSCRTsBSmdRR/F9SfL0RFtW3sGKSvD49o11AyVEd6/z6zPhpe4gJ
Wu2oDkOg2qfAqnS3FsRZ5LBPBybSqs6gA0IQXofyFZSbBw2bu/CVvLxgl/px/FHV
U9Zf0w2wKoGy0XTmFkRAdEdIre6xVmA52BYuz+tIol9nBZmd3jZ4uLrpMAnH1qab
4YI+2/w3wEiddBuFLhOcmd19VmRE85PByYmwCJvPtDHr9AtAadg8XPmhVpEw/Rfq
fYdME1rYvCkxC8k2aaum2C/teoopdGv/4y5mMsMtuJXMWWRGqHdjjD3gMNDgOHbP
ziv/XwFGTojBN/rpfUUfDogIckQUs/B12a/VadML9yN86wVYbUK1d76sAgA6WW5m
rIawZetQ/dKRey1XwjvvqPX5rRQG3jaAfCy/3LPeQ3PHNGCWGz3/cgbq0adtyqkA
vaIc3TPAxGu+mbIQkp1QAz+7CZRgfkCetO/D4vqzFx9yoa70LxSIE7W4hAJxZdts
fE2nrQV1DT4GElcbwnM+ZxPYWioWoHvasAeXJ8ZvSk1IOM/3msA3HD6LNYfU0P4J
h4Ivek+jL7L7LS7KDjPRiHW/yYjiLXLVVgUTRt/a+FFJNfjfZFc7IFQvUfyQZGY9
dqtwSaL7jLCJcbZcftbumixjqZ9edgMuObZKHvbVdgq5HXbtRWCv6uAbVDBBlSyM
dFihCAQKA8/QH9EBa+/AEi8xepaYE8nyIVpypVS0rZFYcOo3h40+6ChHSPqSZvSw
Oy4OjvOdcxCW1VDi5sBzx13BhDjg6VTCE6yZ7cgPaXKuxzfLFww+TCbQd8DUD5Bx
Bk3UrGNTdQO9UjTrypAN1/jZ2pV2NLB3wGEasBL5Zy1nWIU63JfSlCiHVQ64cKwZ
WSV/+HO4cpcpWunPa1jPynbiua47Xuc2QfAquLDAKnzn3YsnyAxE4EQ7j3tZMxrZ
OBjzwNTK1g/UM/bKpSLV0ASoHcmdOU5gf8Mrz2S4M4PG6WUp7LLfvZOmByt8DfH5
svJcK9Z+VeNbekv9qkCcPNx3KekZ04TPBBBIARdSMVgdtQsZEG8d+x7Gfb2/vyJO
VYLuug+gUF3hYWaSxNCIZ5Pg4fLUbpEyPhoLKMQdWVITaW163S7s4mMHwhhJZ95w
zlFzfIwHl/9TcxVqdvrFalZjYdBQI7wpri02nL9sSwgqJpg+HI3atuFQ1RUK13vO
pZAaWrtexY5e/xKC2gEkZ8LdR7FiWY0wbQGTQqe8O3pMrnpjjDYDIfvJZnhiewZd
JtFIdBhYfy3drE+HCHeM7vE7iM9emZ5uCj6dCY+0IQple7lCuSTZDH+WY7+xyMWa
+PqZ8pMnPOrLwnm8BCMfvFGQgvKQ/qeMWreussfHFcel4qDJIbxuHM0QpZFUIps7
c2CUyaYGtVn8vQnDSPrtzODwDB2aOqFpf79v+EWqKql6Ov4iRrG94mUcuf4CqDvP
lG+PT9EqTpSi5DanZT5+8N3ck75hICrIukziH0u0pR1sJjW/CZVoY5xF56aNLgVo
HjVxLH5BP+oq+2e4wKSf5aZL6FwJsXrs7NzZPOZgPleLtcKAvxaJ1LRxgge8x+AY
CJHxxRv7k0tXtXhuYmxGmdgq2/aVJjJliym5vS2jSFLMKk5pZVRmCyHTfwm4TAOk
JUwaYkQ7RiXH1IUHA74uqaocPMRmjHl93QJUvW465yKC5NZ9gjJHdtp/aBN37iU5
LvVmIg7HKXvT53HPeUoeeYlERG82whLO7L50myiGY2ZYmdeYs5zF6uqlLqxstco9
YEDVySy07Pk0YzcutZtjVuu1pBSDOP16zHfxIKkPHa3sW3Bt/0uSotP7I6V7yOvX
xvIx93syvlQ+hmUUJftjq9Z5oOwVIJoY3OoMakVaULmQZi/EVMH5fiIFdOZCneG8
HdojnAxdsBrpZCQEhtUXIfgxWXZPUheEIC0YROvSXdngUUnrNnvMUVyUzlPCwFBw
0datw6f+p+WfD4Q2XGKOOlSPnGRlPDFrUKIAvzYKdSZ5Pru6fhZ3KFCKf3F+OxiU
jhjUkorXypf+ABad+KrA492NGx1HJZn/6ops3Y976mGSCt6YuX8bOp5vqIk7VsuC
ig4aMyuk8VpLqb3CQSmgC7mV3Zi5/fpXJzRoA6R/XrPLbbQ/TnAy7pAXQR80PQNi
e2ZACHBsNR7F9SRg7pl7C9aPqXSPIyBVooV0jigRCjSD3Juvs8RF+Up1c/Vwb3/5
kzgTaNBceK9iC39+LuGNUnegkofVGVlK6Cj3imr1t1g682AKrkQhInjnNkf6KDLU
DSEC82Gti8ekRy0vf9LyhRpqT8UHxvUGD9RVWXoHvClGS+jeCk+5VIO9zqapj9vr
Om3tlB8oQOxL8Xq9qiEhKr/k92aK1sLcKljYMi6WueoncTLQm+SbZyZqJ5m41rlO
SwQLhwrnqx+vPq52zvU+qTfmEtObBUpvzRgNGPiLOqh744jniK0RJylnlwEDf8Bl
hbNGKTGeshcSCYFCoUf6VSg1t7SXIx+dmhw2p+dHUFE/8lqICq2IWxo0oogTGGhQ
g77uIguoXIjTDRFc/6JJQnSUKhCR+peflp5oAroPJ8z9FPvbCOvsBvQf8Qbo40PA
QCgC9tZf+hGs4kV8XrynnbM1oVry+/jiUuZk6vRzNqroNGttFooba4WgrybCwZBt
MH/2D9pX+nY/bM47DJxLhu3f9CnabhSPKXzPpDuIRLtH/3JEyZXB+Bp0chLGvvMm
0M7acz/bZGVJ+co0nPZ9U9sI8nd/C5AshxsqXwn+jDe9L3jd5FFMyUtZSKrF70aV
a2alu68S9cVPVkDWFHf346gLcV32F99MAwNsBN3TsyQdyNY7QwkA9ZhfMKA6yaTf
K+3I8+i9v5INy1uFk9IYlmbhprs9v8A1nh29iQF1UMWC9DhSaujauiYNSnbZ+Wtm
ElRafDWF1me2vuUUatwrWZ7JchjMV7sHCuDiQmGV0u9/0G2lcHnvsvq94Csy5aSV
Od/Y+E+5ACuG6ZCtNK8GxjfXETJ4draLhfD4bEpLMLAb8gAKoPsP/51LrFRtwF81
KvlaP8swYJ8jDDu2juYe+aAbOWPp6ATgjpVl1fp9HiKkazcq4RKgsS3wLRYCQAm0
NXysTpJ8egtUiQ5vJ30SPSqtwMQbyoJiDcN+YTX86aCtMn4auxi8uLw4QXDHUIpw
BIx8EktU6ooymcwVNqQXDpFgfQ5vKFOfxTLZPOhYq7tcNll5cfoSmWbc012KnW5e
tozY2iTZ2/wvotvKQoneqd+TSodxMyJIxEG+Y1AeOSCk4bj1p7xKyE5Z2WZrJ0Fa
37D9WcG7NuWnpyqm2Ug3jM6cNtNKDvHpoo48WF4lEP0auId4eJWqncGLi2X+JoLi
E6Ec1VZ8DCddu07lgssIX7MoNgEu69ajP/hIiUnX1uAjkIrcxLG1kNj5t8FQkBuz
H2FQrBgOpoROw44Z3ZJf5Y9z9KxXoJFp0+QJGVDWImFemZ481YUsNrzOMKrFTVyu
Zqdd0ehFqPENsW8wtqS7SKrMY4taWW7RIA/nWBaR6TlQpQE++D5+w2vwcqgBMWdH
Ut73dc1ThBPplg+mW1wLNlRGVubiy++GQUGQ3PrtfKT5k6j2uU7noXWw6WdYV5+l
jEb7p9ck5EqzW1LsFe4VonwK+pdVQo5fFo4QlZf+8O1Kx1fsGUH1ITxjuEcRcsfG
pq5dF+DAByiv3XI127PMnjFfnk/6eYF62loQb0URTWc1N47keWdWxGUtbLNgbWTn
GUHfroxQ/aFlF4hb+WfytSKgzGWhRS2r0/kZQIfH3G0kydnLhGFTdCx5SoPsXq1Y
m+nHbXL/ZlFhUIJqsmU4k7zSymLChSXE1FawUlngGaJE5MWGBohlx4D61gcspYAf
R1+I/Mx2Q90exVq2c6gDP0c/COqLhvdkDDnPaRlqH0aAUyGhs0kXv4Lh8qSBCOli
RrcjZifBAsD1CRtSEekjFmwrace3epSJeM4OHhcDiSMMr126dH7MQc2w2l608L6C
FLWX2mkSpnWyNFfat8UItSKV8UTQAyueGEDFp9zK9flZa6BAuiALklngtOuvUOHg
nhAhSWvvh8Apm8erPT3mcD91aTHanuF5iIgtRRU9LdKVwnMsxRVeb9Ch+vqbdO4E
OyLl3COLUNuqLsW7mHlOhs50kfaMygPd5cRWxlrNwN5yhWJveQtiHnfF4nsDER6j
MVzYfXIZtjhwePLYJOrz41GocIXXZMK/LErabcZK9QMUnKdCr+RbiP+TpyTToD+J
AWA4OYva2rMsxFeZFR2/2Q0ubBKFlciTgtzM5fkeNtQmW1bwiLwv/IN4/XLsLXUf
L8uNRfmHbd0L22CzjKsnxQ2roi7QmjUp9ThPhEOhowy5jouTBaYq8A+JKatZpSQ/
kmfDtXpJTKGYUlb8zRhu7W0nln2fTjYzN+YkKJseHOVtWMp2hZV8cBD76SmUbfXH
ySObnfJxVfAY2C91DPEbslO0gC+IHQoO5K5QOx9K81oFoBSapGgmCMnXo2KEeV4Z
JzB6i6OkdKU466YqDhSmCi+g0yC5d1kyVVf5ABzOGggSZStJ8dzxUS7Ma1FuoZrh
YpM/mJRlqa0D3OznzlHRPAhnq+37RwcZC6Xz3UeAImglisMSdXQkX6GyCQ4W5xZ1
GH8PGTwTytexbA/FYXOJnpv2N4hitYCKeFw/jKafq1uR+m+5dibtjPpuhqaCtTDn
ra8e30V64gV+LQYX4feiEK3KCVLZBkQaYes73stAcYlEmyIEfc9s5KPdBi/Qh+DC
fImoEcLQdJnAmJsiyNVJYnOfJKp5uXxSjkxbdPI46H/ZvG8vjpjTVt/U+hPf3GxW
TJgJh3cCGXcOPKTvimNXcVMzz16miJzDl9olOLsA9gHVfe/w/esVPXv2i5xmkoN0
VQSnpGa0Zo7O9A5jzJACYg5sqOhdzO1cKyqApfwHAfitYtVCIdD8IW6qdpGjMOOJ
+frsQvbfvXk3vyfAd7XF9x2hdSVkTJW8AWXAEviB1/hpfaB1YHqvPtjxeZUo2RqV
jYT/rUZJYY6kTr5+nUzgololsauU0QBc9dgXh43fyRT2GZCZ/1a0m/BGYd1hJhYJ
H37YCx4ZB1R5QyxzqdPpePemEfQftFyGiSLQ+B5BSv/EF8KIGDabrHs7dGVqjAcN
4rq7d8Ox6j75xuF6/ge56st1NgUgMsHoaj4KnmYc48McCMxqjpoMde3qmZk55ecL
k0PUDUvhQH5iZ6hmfP5bMNWW2AqBwR+YAAcvAdFDsaZeJCBv0a9K0IR6QguIk/3F
HH4raiqiirogp9xUeDwDNdsqE4Cmo5VkXjfVkrsmZ1J2OSFwPjorSeFJJqvUGxhj
3FsLRWQ52QpPPUryid336NjqcnNqK7L/XOwuMy5ii8shrWUqzpwUJRytOwVMA7XH
e1fRsWOrD1FW/NwgGmYveNKoAlpHO/95D5xUtRwxE0YcwQL8OY+uomim3rWSr4Xz
ftuM8AzAkMprY0oxndV5FR/CiEfl0rLdWvyGsQc1LfmC+ZIhv/j0rhs4NVWKJ4Sp
McZaCl26oXTtTbKBLo2xfCT2I+R4BQb7meOrlTLW8GbxJIiZLPmvQufpNWiiME0o
+HitqIhapj0jO3uotyUQ6JXXYHDkQ2aW4WILvIL41YGr7fmmszb5QqiPtbQ6OTTB
AvIsnDRjTz+Ih0KvD4DtiyPbmjJ3VP2Eft1rryvnpT+1AseLshu9sTdrco+UnsO4
pZ8wVrRlDl887zyWozLNRc0T9ZNkJdSRKSkNCArQ4a8JCrKRjl5CS3nVc0Zf6ZPv
nWYNn6nNcH9Hx+y5bm/J2Hmo2JDmfAVBad+yA4vsWsWBB0NavXd3iJlxihX+Avm+
zXyxwHnbPLGdx9kOMiWBjGplfxgTtpeef6gEToAydhK1SVez8NrDv7ehhWdH10v9
+3PSXyM6Y+rzicFIJc5GZukV1fQff2eX5X36Obq+ZC6HSSz3dkFg9aVRadWVnbW3
AX229nqsDZ42u38UNPMBZ4KiOkUtvIrObw96frmiHkOvtSCXd1sSbKjZKrMUj65P
dVNJ7NGYx1w+GGsp9LKP1XOkJKTkCTYxr9aTdn2oERFQlo1e8XiERApp14d4ADPL
VjjRhIejurei3IkiIkldTyP8468c+lYxyfKYnG74OZZ+AzNstwMBw1/Nx+m+g1Ge
7tkIWQomm2Gxpl6kv7DbwzFjNagQ4h7/zOFwqgJtSYTIxcfdAhqQCZ15SOlfMcRf
oEit5D2xWLd3rI86IWBes6UkTYUrihxtir62YTgDxaoP2F/dighFI2dWh3cmC3Od
wrZJoClObovPHBhynPEYcisUO+0q/lq+bYdJgilu0D/lfvPU5ljgjCiiejZqqAk2
i0Qvr0PCaU8npAF7Lo92IxNhiw84tf4QHXMcMF0pdqBQqedxz5Rboe/GOy+W2SWB
yK4oLd/lsF12u5+8UyIHiiQoBXeZUFfzr9z8sRMQvEtd73qWVs/TQ5qgdfwo9X9r
N6uhS45n0bSWk+hW6+usar++Q5ethVUA/YkgjItOtzWxmkOkcemQSPx9+395pmUn
vkSbjdaskSOghTd6d92xJ2GNL2jhF3YJFXOu6Ywdy63DS9ipeKcDhfc867w5JPBE
LCh0MtKqp/RqjAF+7Q0atKBgIfAC8P6zZ8HARvEnZUb2zA1G6zsku72bs0ffpxsm
nRKMBliCRkCp4ACGcBxIG2v0wcDYMsQmpVyxFZJJ5V0dSs8FBJAUzEvYK1Nlnv61
fc4aZWyIAPS06aRxze7f2NbXlrVIPesGgoQ3jvVpC+/OsPYywcLVYl+N28XYGIdj
mWls/jwacrzSVzfSyFfgAqXUcTNywGYQSOli/nc3kc89cSm3QAPdMqTyWk1z9Xha
huvmTFeOPfSwdbuj0/8aqfsMPIhf7y4Mh6T3ARW9sB0fki2mt+YaWmH1LAGyGODy
W1KhCm0EAdvwT8fov9xirrpfkrwC++B3c3GkUdLXAoIa4L11fixOGuckwYXpJ7BN
IYDgJepBtsgUEmgqsxPaN0TmVDBdOj0GdP3w175L5LnCxKZ2FcSJIa0D0DMIOf+x
Dwj889l+v+UMVKvkHmh9EsyrAdpf3cujFEmyN9BQ2IuIIQRqxN3cqwgC6FOL47hc
ZpB7m0HSjyd/ronS0k/WLS4eGk6uGtN75QAgXuk9Il4mqDsWupsd/JKee4gMSrRq
4wkVaw824deIR7xIgYLWzfKE25lyq93CnuDnzIkJwLcSyYCKrmLz4oHj9m3M3M+d
LCf2JVXpkGiTDdVI7gSCm0l6IbeA1OE+EUeiwu/wonAVza43RaSc4KiETgjD8qPa
P6jkHlKkckqwO/QP7Aiuuui6J5we7Fuxk8dd98Y4bd2Ydp5BNJSxIZsnTY4o4b4h
LEkOsoMRjJD5ANNbqTJQwznvYD3MKDTfORZy8UJPp/U4XstNqPvWNjzvxhA+/Zee
WMagrMY2fm5TROpCKivZxLauzC5kQKDdiqEnC35WhVi6I95KthF4q85DGvWF4mI5
SugR5Iq/h3hL5ji6NNO/xiwZAn0JB7xF1pP+CXSV30Ls++qOFWDQduJViu3nPew6
eaWkTv6qHUTq5kfJ5oeFZOm7490410LrJffhmXJwWM0BnVM84GhBX0tIYTvirdIs
F7KGewW6DvaCmr/Pw6wkr0aS8ULb5XgeeXY2TMpMx3QzEfA0oj4A0FoQvdTjlTFz
skptUB7gbZi2548nFYa0h01hbJWOoHMeEhySlrNCd0BRFvrA4zJQfPqeC9FlEhoB
OILP7EmoDw5CvQeVM3dRqrZCqLX3Z0VkmaBH2RHqv4RnrMjKVfVNgzupuSKQ3R8O
Oa8RRWYYoI2VRjeguZGuO8wFqKohXnIrqXjDY+6EWnh0pCeKkvQ6DpZFVf4Ux9Cs
rgmVabx29IzgwaDSkae4wuiYsd28Y+tUZDfDAoR+/JTeA7gj5AUiHs6JAjIpBi+8
mR2x/6P2rQP1Q38vAb8dSaTRqr/8nze98J5xeBwdj0ch7ByM29iHsXDA1egNCNGs
eIKR6/sX+azOe/EJqr+p4QssTdtm4TBv8WF8O8miOOTeE5CtZBbQGKjwvEjr9Cfj
/YZUBNevfWsLw9+um/CWeqZRh3LzaAUz6Vl4YG2mPWyHpa50B2EkhzW6DYpgB/w+
nmlJ0chM/TNSkqs3SIKLrPYvBWxR7NF9tvrAYb68X6gPjWtHMKG6vC6khY8RDeUR
6zYmtIYJ9tZRAWmFru90XYYYGRsxsIgzGXSii84u1WPDjK+zhCXNfTYFZ2GRByH5
WWq1PJ5f8IsBX/HB94NiWQLmPSHeIFAl6+WawtmxEBl8KTFVnoDHIKWNw6uf0lab
WAi/yaaa5vlEWtquAKubhqTeM4Cjxw9B7jxvktm2feXmey5Cu5c/GwIUI0vUMwRy
PRhgI5iH06VqpF/8+J527g/5VJYwkEl8ObOCI/y6bqzUuQf/WxiydGQkq984QGAy
fO1vQjBlByH+DxO2Jl2SzOgIeiWbftDl/nZ3SIojvW71TFHHsBY8Rx5K+8LiGOkp
HeLovpqIGwbIbLnBplpNwXc2HlhP668CQ9zzwjB5L+0R6Jal++wh8FpKtCubMgl6
Baw98ddBQMma7upL7Z6lL9I3bYAcyqnag0ogjlGYEwl1NO/jtDt2eQq1lAFHz5sU
tn47gpLCTmkkmBHoEv8B3nVvT3gbZaYtfCregefe727LUcxhFq38/hPrOR5ps4V9
h2Q5zx2dNlcB9oxUt2103XnVhfYOKBkiyFPDyTX0lLiCTsRsWhB/ZozDogE/Mi5V
ojLv1T3b3T2GBxvmJbkb+3VicAOkPVauvtpbZFHUNAX/Ini7lwKJbTRH2WywZkkG
50ul27R+zgOWd7W/6VKrZE8cC82qq+AaHal5o9rl8CeDZTIwVKLO1CMkTFn2CFE7
gBo22vyLPoLwx8Z9/X3hWKY+GbgSOR01C6KKDUgoB3vQBza51puDLbgRrvijAes3
spBWz/af5aQFfJmyds8al5c+5RtD6iM3wZaeUtGpkEmsIuqeinxTT9tDjfwU1BOb
54wUCiK3zSB/YJkVzBKWhQF1IL+Qo/qp0FjoqP5TyoQpVtlkqVd/ma2U1icV1w7K
M0ebDmP4R/8O5HAj2TG6tVALV1iBF8JDVMT4KrH1eXh7Su0jQGAxkK7zASDOwyFt
y55KqvHS4ohuuST4nDkI6IGOz22s8ibF4pQXHPEpgtctEy1wbf7NcLGWlS3e3XAf
ttsuqh9FZiZOg4QrgKkP3VHaYxMLE+LjgqJevYbdqDrXksFCbWGp4q39rkn2CnBw
BRKz3FfEpAcOeXIHpgRe5HkRoMRT2jF0g3tx50XYPlzkvBhVosZENwQhYR1bABzz
TgaJsPBtyCTyVZSGAk6+VikNM3g9QPARdiJizX3RHc3Pk6wipuKSUs+s4KwJpRaB
L4vY9W+GsbnIEWmqncjWE+lDTXz4UdtzVodYTITiqMnue38yR5C89snPjHHRaFFA
xuoX4EiAR6fWnvv2gu/XHzaf6P5Ave6S82QnQC29o1NKuayoBhmK897Ezd197qkQ
jWB6JTxRXsm4sPmd24DCluIXviMfPhlO6Iv7dwIa/jDoiS6sg+uYN4Su6PJxEOUR
k08FxpP1qA6XjNhnHKbcgkG1rtqYzBFaLGCv3MDtBKiZkcVDLkL1lXdcig4hrPCz
fMHtptcHW6ccvrfM432Fxe15QdiqQekksawwrBTh5Ch03t/LT/JOSVcMRs5FrwBn
DN8ZZFG+LIdbX0IS0qrAVKLGxq40WbCdRCUFiNJj/Yt7K6LF52iyUwXpzg5VbQwE
4CVLs7U2zwLA6ZSQBsbN/Yvj5UeQaKEq2KWrAFBodS0O+UAzgHhP8vgLoifuNgyK
sB0ZRWDii46FC6rR3sPyt64VXQxCeg6eL8zGoPHVLn8Jt7yUT/eT6B2Nb41A/YUh
r+17ackd+GTPAv0UueyK/KnSGkxLZry2SLNPXguiuR205eKd7STSc7dv9ImTWO0b
hf+WwRqoKO5VE8W5eqkrN5XaxiMxoXbrLRZ60CPBwFRDZ40GQm6zVFmU++K3cfxl
jpYSfFLb8KmswiH0I3aRMV0DKstwZz8VIApM3y8Pnj3T67FqkGrb6MQtMX2Xukwq
MqyVGEaYdV5HyLICDTQmt4E1pTODIEFHXUwDQks/a84aOlwkwsJOCgJBw1ngOqhp
V84hFWReulAzhHA7UlAmhipTjPKiKt8j1OTJ6GU12oqz7SpsDg0QDtGcsvPLZNaT
q16Y3fzhyRZITzpegDqkYrP1L0oJQAi4yVtAR4kpGPJtoiruFFuy1Fo6BwOrsa+6
bkwgCWyATIc0A/M4GQMKMLbpymE+pLLXfCTdPu+d+UtcYi8zKsrDrJ+xxOFQL3jH
+HpgDVgm7UCPgYFJoM1857BhlcbVc3JVV3y/LZzjpzCGu3tz7EOPbdjKlwgT0oo/
jvhbGf/BZSW29Rf6h0o0yz5JG60hmoKn8++zqavs7V6Mi++KHaAbAL+/D2QcpSlj
a6nmDtzvqRHuoklkduOq5zQ9BpothpfPLL9NMUB2WJFW7Lozt/DYvQFU8uL7PUh9
KvNx0+nVQ/aLrX06pxtqmhV5rVxwxnN8L/vXt/GvLXHY3LhuMlfxvlQUEjMoNo5J
hzArOturOfuXZ+fo+9EJgJBFmTFkD9XAeVkTc7cIe+cf25yRAxOWTqLECo56Ptwq
s5wLB2qI1r+lwe/9eGzcz4JB9bAqwj/iev7F9qpcTA5raT/7tvX5vfRKJ4YmZpI2
8LJ8AW+sfVbPbIKAQvfbCt0plWwJJuBLbu0RM28VShFPnYgPrrjYOWz66rxGda7E
1uIEmAl1CHke1/ESnXZaBSdlCr16gOsFxeas2OlJHB3Wb2KI+6cJFkgX8EEsRg2w
7wxyRiCBbA0sgPPNd1jYA1qWt/sj1H1xliC/66KL+SAKK0HME+mThWFV+LUSQvgI
9KHu90AgHQiXrQ55ZavFuSiZ6+f7c9BQhGXTI/fyNXCXDqh8JwZsU+LA25c4wrhL
afhuqpdyTJJQZIa39yF7FS/u1dp5Sc5xZ6FProseEOlnqRJQFseBM/j4xiFSIS4a
4T/Iy9/t1GGXl1PHITWenpypP16KSY+4Cv5QIWOUkOhQJxicL0HdJwWQj8OtVNYx
c2gAHoe68TuqQHH52vn2TtmafkL0BcLgDPumP5YqdbE0qVS5IYjBoLpEI8ddYCSP
yOYZmkWGaup0q/DoaDI1JRJiYBUEvmL6d/mehSX/ltkv/e+l766qogIF320WE5LK
wAwZ2KkPX25X9TXzvf+q39yhioCk00o9U+e6P35vJ57KTQj8dOg19ITi0pFfns0F
JopiGt8aYJYWyElNVdddsV7CqtmZz10KgNyfVRzLC4jy9Tn9duAhryXcU5Xt2d2/
G3VZ9hNC3UgEcNmDqbebagWWAAQjqHCNQhfq1GpTSIPMTSrm2836tofYwiz9YL45
oOndokNK7Z8ulq1V2TMBkv2UHDcoO3veT3bLX1jp9qp0ozXx6BXV6kzBLhDmrTel
tXFamuC/Gggr7QSfDx4bPaWzz9GpivUs2Ydhg1WptKCojc9MpMPneeixZ89R/KLT
DagTPC4hfQOA3Ragp8aSUnnigukD3Wp13lRVRbuzzpeNNkV8jiTtiNDCEV5NNwlU
tKjImkPmnkqfcia0pNISZ21zz6azQjuaIKiV0faRHlU+VzLCkRV/UC4a/qEq8VzD
hG1VNiVDOqrod3K4a1aRzpna73LupWJV5KDhDV8WGLuknXgIRA/z34Wf03faWr5T
bj3cFGt3igyknEJkQ0XftaZ/j3uCQZyrvljd3CDUp+ptJKHAab45Y4A1x3deRYEI
vHLY6Ul7x4TVAfkhLvJb+16B4TACZdHATYHJG0glSlcXL4oEbGkluX8QCerVZoWu
0rJAZWCNLk/0zzNSgthI5Exp681XvQXxFDzarFSik/9hc4BhlqB9s4A3VD8eromf
92sXMYt3usiOX4fEZv8TxykDLHOqiUfgiZ4VR4Z9vOeep8wUAKwHF9XLVkhYlFxS
K4UCx3KNNgoph1QoTjfgGd18GhQ2o3nTdDSbxh6CqNDbgTkATilWee5CTcfjeils
KQ1ZVPfxQe9PcquW3ZWBPbk3jEpfBXGdjfOkL1hGZJX2JTBxpy2BWSZbNlOtVAVE
IBRa/u6XMefw9kfHb999kY/ritjH1eKAzeMigNJczIZJ/6o+/iy2OsHwr8A7zbfh
ngrK8S2YE9d3cTGEu4LvU03ysalCEi+mlZI+SG7PVGgbAPTAdyvkU0HWl8DqPPrh
XS7vY1+4ywy90sA5yI2ueM4t1WKS/wnrX//8p7eoEwL/ftL2AoUgvINiAEAzE3ki
DcjVzLLwxjjRitfG375T+j/qoC7fjsnRUaYRedhTCsTUP82WWIB7epP/sKYKbRdW
0OR+8ayBViOWMbN9E2HQxYFZs/s771bpHo9Bht82olk/HnzPwcNpp6gb7EFi59wx
/JP8Ps7b39YbKuAGev9nRT0DsT7XNWSoRdXLccgBswpqJRvJv87+VsOEClM3qask
t+MWvXE0qBA+nmAUEqc3KnAkr6iGoXF0A+yKlxUB/hWbrXJxjn17MYzvhhkZuVCx
VlyWcVwM23ev82CqZcqo+47yujfBpE0NoW28w7RHfzkL/3SGAMft1RdWXiaIv2wF
ES043t65GV9lspKraMVcTh87O7NoYhCnqTGYd5Q1zpl72cFhVnbUZFK/O7ikKx07
KqUHDLf63rkMyvMOtA++wq7wsxqR+y4S8B0iihvUnZFW+7XUn+Aqfmnfzd2wEaxk
JMtWBO4RvCkQyjUOxeZtUPvp6RhM1LpMJMmBoZ6LaU1L0tzRjsvhxkMX9AfaIyIb
KPUGiqHKxRYnc0EH2h9yZfdi9Cd7pciK6DZIssjpKkJU7uwUF9aciHy19HKQLW5H
ysVPVRYDFbNwvMogZ8HrI8OCVJ63lon/hlPlf/umP+bl5RGC/89sakmSEBg5V3Is
mKy3uipSt68caEfpYUoElOfmY9BcFTksXc7Ysd/nzLyLKWbOCZVH7Gfd8Us99RYi
4TOxBq0utSzH41aj0Azir08Sj6kwozRtz+3HyyXfbP2okcmHHgnrBMfqIthXeEwj
3NcCEG6imWEZjAxju4Jph12pYvF/4LIpIwaGpH49yS/fupNYnPp6hMdwDibAEN9F
HnAUvT0Ct/zCOtT9YM81aAs2GxJf2KhEK6hvfB6tNSLBGK5Zw10g0RLfQZwFI1Gc
+cZGdJBa6bXlpXPZkN1DPO7mHtrwppbOdk64Y+nil8c7z93jdPomEJGqsyveJhOx
XPWo3oPP8WMaweZ7Rior80/o15kWHBIXrysuhKvUCIp91Gv1IAbW95KIdkIgv9AI
YFWpYzHWAwSWvH2OxZNsIhIrOnoR9Shew5dxvJQN8f/jycGwZC8/WIO6sbdL1tFk
OHb6+8B0F2zoGHZN22Qx0XrCBEUxEPc9LcffYEFDOQdfBkKzNMbpLt3mXanCoALY
Eeao75BJ7j+B4WRMJkiohJNWhj087TiZIhbjaX3u+KbrwwORbIr0mTGLPuaoY3MX
Hxfw5rcnyOnlApZgQxUf/SCv1+t5ga0MxqCWQ9qq2CyHO9C62x24l4QcP2d8b5ox
oVO//bPKAC8Y+SAm6yEABXy3peBqjN4KzfNDfLHcDljrAfH0uLLWRAiAEVEgvbnR
/1vXEhL7xYHdVGhDZCJ0Zw3KFORaxd6df/KHcFMwKXFGuldm4mUe6t1Rvm4Xla3O
C0Ko5CJWV7PXoA5yhg11fLbgh74LdfTlrLgEpjztpJCvnQeHug4ejl8dUUEcBytJ
kL4p/TJLmDLM2cKAWlN87y1sZVG9ieDy8uOB/Myu6P+qhz6AVmwskUBVQTbZLd50
FNED6FvPq5hllXbmVsoehuM6n5pN5gy1n5TLnMS6JWIAEXk8GZKQxQIv2GvLIOZv
cPQGrxHbZ5DgbKStLtzzIuiLbjU1oaFttNMTBIVoQ1cT5oLyvID5e4bz1W2l1RwW
bQ1E9bWKJ+5eTHyy+RchcujjG5iYLQscQ9ik5Kj014gC/H1BvDdD2RbGCHd7ehTg
LppEpgxXqvzraRCNQ3Ndxn+dAzCtimwNtCovyb+EUaH8vaUCTaAcJD7PYfduPCz/
GlzVii14EXGbp51YCjfXIEh7fQcs+zjjl9OsXxP4kaCWvsNJ1H6p/Odr3XaUkIPq
m9vGnJiqY7dLVYIqjEE+EBmiDI1GNgqi2G3MJMoMO1Ych0xVvuIIVy7wJRrLrq44
3WVdxGrhA9bQ/JPw5rISrpUt1EjuE/eBQSyxs1UoSR30SrOWMeJ/SabtOalEQJOB
PmjCdvCnntzjnxFVFTQauu0pcWvumeKrZW0YzrgCR/RrpuxOnmV3OvWpvjEf03cs
4QN4ATs+QGNtTlXPeYyXnkoXk1rmy44UwSdwXbmPvrJWhK6P2737+Q/7MWf7GK7q
IPCITBPEj00IHouzbiB69mGv7D3kLLWLFhz3GiawOodmJssdmvaQzyy4wpzwn40u
F2mydKyeqLlV+A8lFTnVk02v8J0blrk5QqOjfON/pvGDZ8KiG7RqfL7T61OshwxC
tXwnwx8ItSVGBJaDTHuWMrNAxCQFifCqowDzcuFU8JuIyT8vTmG8GQTaKbcxuVX5
lX95PdfFtpRuPjbLDu6AIWCGWTHZkduodBrG0mt2eVc39sj9ILtlGXk+sZ5A1fmw
xSU/LtvsgOzAjrey4UqTnT+8N3jDG1vMOFeMCpxtkNeTm562LHapWVqzqqWzA62d
u21xobIUbbLJawImAvFMSNsDFgvX9Hykyz/F77jx/z674D+JQ1V6yo5G6AuIMUAp
7sqHaULgBFhhgpowG457m4s8YeKNISKtVjs90FhJnjH2YvxE6CMmyBqDo8FieN3W
FGlDBYGn4KvTqfh4qfqSJFpuVuBZEQc6LrREPEIH+5PiR3/hCySKILujqcTcOLUv
wOWxMV8wiylwut1LqiU2igFaID07a17qFqq1AnbSCXIu2kv4QARfQCEMtjBZeQDc
BLopgbdxIK9YjH+LIJUkn1mBylBKelDvNZNRbz2Ru1SeuVBG3xZJHlxrsXjwuIoU
mY/Hpg5Vg1gJzT/20b7ZlKVPj5qvCSbEh6IqfCRCIGDQuQXX/hLIqw2RdL90MT6s
Na7iDizvFeU5/aHtJFDPm/wnsFvaUb5Ln1AC/JtnkQLVSQeFo84/LM4QvIGiSXX7
PIYApkoZ1Z/JKVPae6TjSn5LDt+5IrTy8LFr7Z3xrjA24X1rkBa5D0ooZCrYIS+f
BJ4eE8Po43m5xOObrIqN2qfBjcMD9J4YifjGvZ7pSy2V3qDzEGzQJPM81dkxtygk
cufv1CPG5xm5CGKOC+k73NRWVMNYl/zclYQAX8qtGBDpgX/dAxSvZTx3AjWF2wjy
wz7ZkzITJ3oK/BA7jsCKZb74mf2R2sKkqXidAUlc9F472pR2G4+6o9GeeyFJe95A
uerfLFG6iu9VzSyPgpTIvjeSXP2tPXDBcNYxF4Xj6hpRhDR4MBDZ3SoawCFB74r1
BTvRz6cfK5+MkyX1CC9gAp5UqvNPGQILSom7S2jnaoXItnlgG9mnA/qOhoYq4TzI
rus8OD4guHkqbP7pAMoDYWCIy6dzPbv+/bPyqa45E/uoaGp2vtsJczjWsq2Pw6PF
/aScLVittlUsF7oCT1H1s7TP0GyIazdJ+12sOqZc1eNsS5UfoVVoaWOh3OAto7GY
+QJCnCmhSZaFAvz8uK4ykSeATQ8XOsSOl0Jv4WZUlLc4PhsTcoYorrrzneKXosoC
zkMwa5LPHomfdnfb8wyx1hpTvaZnNzrKQVeVLzBM59Upo4hGrHPlCASjpuGQWI+k
xPaU9oUwokCzfIxK1ZT0H00khdAaRWK/XTWZDWUTlRJZnckE/VlcaKr//nuIMO0S
9EzqnJkGyHgn4TKlVZKZ+yJwYEaypmsNJSINNZNU9eXNCiXwt6Zek10wUzYFPFgx
lyJecdo81fgEEYu1b5HLYwELL3xzMb9q/2am0yfO5c0kadEd3Hurso73/6AgP1FP
ksPCI9r43qFeohAq3EsdWlmQYVhFgi3kFgKf9bveQ54exFmHBYEQFR9YIlgNK0Dy
5wVTgVeNIa55gvDZmP5LYIZLM4Jckko9YAEoo458vQXpWG9ZfORzyk695He3kJk4
MQTJluEYporX7cv/9+7RCPLdOQXiIp1QoakpQAwmzvcavz0gj5X91G5mCRwiPDjZ
fGqYDqDKuW7NbydXM0+eLOm5BkMjn2VXPjL8bPl32u2FeIKvC78LYIHPqM6rk1Ao
Dn9Fq60HjDDoClf/cDpA5ii24vf496SD0mzizTrrGL7MOmRmWUx4w9VlwB02GDo3
9g33zeZVZ1QiwTe7u9uQJ6+c3rw8U9qsG2Yy+lsUgYTbMDC4PY29g3C/G0cWTtI8
i1pjaEJya6ljW0k9wcXYB26QzLXyAsxMgZqfx04bgycZuju4Ha+oKkxHSHsrUzUM
4fZnrzZtoWngdBdK/v7tyf/itT8pU68xj0V9jXhtQhtYyXWeJsSIwR+4sDWOfbx5
jWqWAty9e3/NxsrWF/8ki6+3IT8JKBWQGuf6BK2b63toKCulI7/jT4jH/U3x49nq
XUbS7Ej/lfYzGR7Oqd9uXJUlgSYwrOYP6K6MrTriIElAqiQJYCI5U529uCfyN2Kh
3SupRduraMIBCOAxSJltIjEEH93bkJsKus6yVEKVLbObyRfHEPQk2UZsmcgq2jGK
5ts9NZDLPLON+W+6HAokipG1QaztdwJDdgFVfK1KKKGqY0ZuYFDurhFraYfxpPIx
Hg/s24ZAbPKApGA+3qyq9hJr6Zf007cLxx/k8PlJux8PUsovTSCjUu2Zt1iIBBmk
V/bg6+mVIS4tNfLSqwtJZuMZiJCVLUn0WmcH4l11XVwplifcIOPSmvkbr52UIV7Z
8zVBkV6sA/whsTN21J6kS9K4Y/uKwjjKGWiTjE6MgaeMSbTuCZf/dYDX/lGmX9Mt
a499JT2reHv+F1dizEBPprQpb8bRN/PP9a56WKADx9uZPqcOhFlmioAT/V5UGE6s
pshfdz8MaO5L4pFfZaSBOwm4aMHeFVUZl87gE+JkClmIXxrEe7B8FToRGjdsRzRd
gYJWI5f5GvOWfHglL7QF4Xj/nI1YtqXSN+QTY5qR/NWnYiq7jxCfOuNkvMfGuh8I
YsvT0wBhfjU57xW1cWVUhYq2Y5c0h5Mw6ljIRdOhbxVjwOJB/PEOUSpAvJKe3+sU
lKi/zVDZgGlB2qpjybuxnU/N+tRcZ5DNoZVL2neqy0tF3sxNI44tjz8pLByKrGiR
faH3PGvRG+MiwHuq97yV4ZxZmEKDbQ66qmZUQVGuL6s4PNkGtf47A2+WhebE66V6
LNkca5ZoUQ2JjpjBWa7j5y6d5Ryt6ppWOxcUSDcLb5ih3KJlaM08u9gj8K9jNAnr
buJWdR9CgH1Eiqrh5eHy2bZ5YKdWPUe8zf8KX/m9gTLr1jVVjQr868ar1KRpB76o
vk8NaBSAH3ZnNC5o/Dwx8qDbIWhrQKAKumVuMd6/3UpQroH7/FQigmWkbHDvm10K
2+56EmEtjC6NNPPPI6FoA/0CskI3Dftcy2FoFFGOyllT+bFT3o8gbYC9w8Ge6lY+
fhGhb4v+HzwT8lGEaTm7NMwFwYeyiHQwczFLRMOP3CzxMxJC5K1f/7EpzWyHfdCG
YLnY+Tz2B4ZwF7ybPQhLFaB7OXApMGi1qUmCiWaf/LLr73SsurVdA8qEurMOlN4q
3X5Ta2KYsz0mFCiD8ZcRg9MbQoj221B4o56Fchwmgd7fVn5ZMuRyhbRPGrxwb44+
hQIp6dSm+GcgXjoo4u/xkS2fn6P6vq4sgGY25ypOTv5uOOjgZicfFhDuDKTa6dJP
k0AOHKAGi7vvaR16xBossWP9eMPOHxNqWtL6q+gFas/UgJOy9meJQ6abFxGAtgDp
pOcQGO0Ql0r0mZ7hbOb+envZerdGWILvbx5rkbgu2ahdJ+SVyvdBfEPVTK0VrjaQ
Rqg5+4isvAELz+92MwG3HZUdYhWSyJaRf2yn4WkPK84yLU71zuUtf6FKWNDYiJS+
x8OlvSiEx6h/mZqVTFxzLfqoIBSBgXpPApYNJ0mEkcyXBUE6UVD3PY2onMGUWJ07
vHtsyzGL9NKdPwgLCv6YksSaoc5BJS6Zl/rSffwewBDFHUrH+tr58HK/grwObTeB
BXZMvbaccUow/3gQStYbIcFdhagZfoFxRPu6hiVjM4lzy8lsyUre46++UJH9sfIN
jiZxLvZhdZvF+8Adoi/TYSBTd/p+LQAuAxNnjl7jM164+gTnuwOA4STfLhJMyhHR
/dpW7MOW98e2tdO8KOeT4/ema/uPZFixSORtvvXr4zYAAax1kj4K2G1PoA0NSC53
NZ3ylLDjhUJ0oetcAOw80oifgahYPJzuqXkw30HDeGjg6OktLYpN3eQFCnzFWuER
2vDbf+3XPp4xyykG75XrPZ1P3nNJ5r0EHmOauEuEZVfrbD94kN7sqN9lU3Fxr1Rk
6+iLi88IpLsg9b10MBjPEztegsncQI6GwLAhkWdIXJKl+ETQ2WLnwExpGTh3FU/p
X0Qa8qoshNrsi8X7qGI5LxmVbU4CBGmB5I5oFzZFztAdf3A3B+qM2SpUFxp2sep1
XlUWbyXZFpf7MLZISE76+p9x5gJK3iyzUuGCW41yzUTDTgPcGvTb+KD11YToB7cr
+bWYX69CF7JeAXxIs9b2RPwYpE/cJ5loisKXO0vXB4nJmd5l/5o/s0A2zDxJOGyS
/LdGviHqhGtNjyDJjfkJsjON8eD6KUdShRGn3pkjZXXf52KoTZSJ2rRRJ9WaIcAe
SE3EGeKNSbiyptzv7QF6q9ylFxopxT4YDDJ3a+S06tZwZmSPTTG9wNVSMYZ0RHPf
wl4nrvueEFRXKMxuPaJFc25v4+tPgYEoFjIdJ9XIutmY83m1fEE790hJ2Z0kV6wG
rS9hwrjpGBN1/Y1UcVLBioNFvbjIYLh6j+9G7aIbErP6P3TjXOrkfKHeQlNaYCDj
CX3JubCso/JGLVI50OIilrJFX1pQVtqNmcbXA0keZiyDKoQ12whQRxcnGh2CDdZs
W+TQFxRgg8TKuuWd6YvtrVv3d8MKt4Qpv191colOdsfxk8rqj7+yA99jfKWK+Fgi
XU/EdK8eaMrE3aU1wS39dW9DOVdqWHWSt7ibDXR4skM2bCZkDtQ6kUJAm4uNuZms
rftp1wRWs7osV/HLlIZD3Lj9FlLTcktdAAQxUVDfWyJDy0A8QHFLvpw3izvBnPYt
ihgDIBkqPwenqz7p6YIMiZKgFwiz3tg+r9D+0d7MkgKYS2CLMD2vri91/Lqm37Y2
d9Jxp5wVOg7jEZ16O3kTPlKGx+RASWHlFFAt97ggwmcURgQfHIaj9UOReAHg7MX8
oGWfsS6lSsYUzA7TkGKtmuMCKhT4xB1sIIw2qTkstkSXTQvcBYZIzhMx/dDIaFTd
tdo43hZlKHqfWBHsUnx08MSYKLux7PGH6SzrcpcRlTcoRZ+eO1GsUrrdU6D2wtnX
6rPUaCvxpN3Rd04XTCRqoQFyspPLxvHwxPkNHayYoG6YDRzDxO8O0qY5uthWflTp
Wp3MlOAHXsucwh8DLRWZ4wgSzkRjL+jgtuuKCxhbjRyF5STyeKayVCKZAU70FsX/
MOoeag15t8juEm/6j+KBnoUIS7pp1TD9AZiyFZMjrr2g2D/TUAHNnC78ACDgqdg8
ArN6gliHcVQxWpfDO8EKPbV5FjnhkTat0STOJByxXoLfHEdt0fU4L8FefhfQrmx/
kNVMOJOra1rZCi+MwhnlYl1abLUxH0aYG9F8/k/JVFPXSg2lcux1vbEC0fk53cgv
6xMPHgLn8pEgVrclzx16tlBfSxoTzz/PYUcQ+loW9BfxUgt10vEViXDKKi0TOzAd
1xwXV0TPigwQJv1jjxtSr3cOBPSMqsxp/SYl4cKv3odpe7I/OmrzP3u8Ayb/njBT
v9tvttlo88sopeW+vee6MQnhYhA5qOaFzTS41oTQyrvs/n2fWYx5K5nl8aRBh7Xr
LZ8WgAk+palDC9XwVS+CK+8HegY+DaosOL3iKbgBkX6pu2g42xplE1EVQTPnfOl6
DNbM7SbCfYAwTF90rPlwyyci+N6XOjfp1h6SNDCSIzdyXNneFHuBycefTUzPz0fU
l7IK4jdmkt/NsthQ5aZxN7OBOGbbLZmLIQ7ya1ZoeUSM7gSBYWRls/0qkOfYTxVw
BifQk2Lf168HMQZBYid5tIViir7ZSFmVMeyXoP4lZ8LNddUO84cRUC+kRJfZogOw
sfYXbIrF4NO1oeKVotaEOfD9MNWyRvmyyGmX8Rc88vZ2GUDKhTNCVxpDPaVxCUdm
jIRS/npX7/3Of2/nPWoou7+dbmhPhFLZyE32TN+X99nkI/ePUfd5wvxg+xNxj/mT
ssdMZsFWH0sxdCg9JHrP4C07ripiqNcYUC1/RdG95aQ+29AjkvyJnXFz8QkYNJ6G
1AvgPMxWhXFzxgfjyxFyudgJd+zlzTlZeuIWgVjFtD8Oj43WFrBNMAA1fltHrZZS
jQnMseWAB6LYoXAHFM41mgFMhvbKqYepfCVXu4fskqUt0A/yM32KhIqdyS1W0Exp
PPjGNucsnpSaiJhswBK8yqc6d8wU9fIDNP3GrQvus8Nkg9JjLXrk8ZQaxOJ+ZRIW
KVA9XKeYW0zANCE8DRzMFaaz5JR/YI+cc4YLN2uYITTSPP+AzKKQQb46ewxluydo
98PRqMzpPfeX85UI0g3lC7YHtdZ+gYW9HfjPcwr922SxeuKC97cjMsw0ed1i0x34
gc1ZMtD97BWdcZQ6P6pycGrjEY4/p8fGfNHbjrDAUFLWCBg8Vtiy31+qwf6BC/wj
Hj0U68+x9PfWfSLw/np40QiFa7zMh1kJZrHSAfjq5IALXdlHd+PxpV4E+XbtH6wj
CXgcwD3mbwhoJ9ONAdVCD4E3+bHV88wDURu28KOu2atlFvG/S1d/vkda9T6a1s1V
mUQa8ia7+oXdCtd8FPt8W6rIRUBCnWtI+kwnWTjl7KHsj5P1XA+aZikWELWBKTvU
Y3nmDIsmv5OUnKyhwyTRkqouwlkMEOtuDfAbgmUOtuJaG4GnNVghsYF+E/L56Ll+
6GVaC6HOWkWy583crHV5QqgoY8RQp2vjCfLT2HBQ/hbn4qO3OywHpiQ16eVqVbBA
sXixbuFiUP3rLqpEZaEyc+pirzk3VQXktJ8hjL9amMBDoNHe66VMC9GEAK3VjscA
vXnpQF4wjXTZuueRzn+DsJnFGQ6QY6nzaoMo0dCTeXXUYo7FtTHLpSQwi+XHEPmQ
CqOyfOH8zTBK9VMOW5M2hQhz6OyY0ITG/X5Ao2eNeFnKFpVWibVJATsGwP2IKnCm
jLelfo0JRp913jiMrYP6Tb7zNniVc0XT7ZsJZt4lm8VExJfjKzE5o00ycNg1JS1E
s3Iadk7/leLWpPXr90+QcxU5N1YGFOXlTG6Pgfk065v1/Wq4d+zsqnlUgWLIWNtj
DyBpTrks5KWW3qAG0Ws05fBodlLIOU+WME4zy8Q3NshS2woregR1YEvrPI/qIBn9
z/3siP7mYOxKR9UUxSmnM407aZU5fZQMmfUVlI8YBovX8tOnB1/badY6Qsoi8W5r
LTQ1zqnZ5kXY1Ihasoajargw2KMJz0/PhJdCvUOeRJ6HAYsv9mbD9KNt1cwJ6CXb
QC9A/XWooy9c56x1BKebLKbRhHCnpE8jaCJiMi0Km0SitZtiBVB8w+vYgTnVg7SY
Fz0K1ZaYhCFeHr645uM2c9WenltH3xXf6DzSTD4YKo1IsIgbCr+MMEPJqdnTjY57
zfgJeWGOmg1XCGGd9liaiqBdgcPO7S6A+Mrefb5i8hTmYR9xzL+8bLXaL2yVLQyR
dabNV0u69UEGfNfYLF0zOEpGZ7sz0TpLph333uXDaqoNyfhmChPJDn8MeNwhjR2W
/LDgDHefEnQqUzL7h0sACE07efHTBEpkUPXk39DX9txjeu9wMfF1sEoFye8Uw3/k
yN+svW4bXDmKvXONpHivNWO5dCNFRN4HOjvluQRrmGZSYdtJuz8p46yTOIhnPO8B
ciKLeaodl1SdEEBbkbfrXct5heWpNRTECW+8qeJeCwKbShxZve48/YjIbqYlA7nk
c42CK1P2OW4/DzZIVK7ALMJ1gZ0max7Wfxw1KiEzV72TOqyEbM0Z4IxBUKY3zKAD
9gmLLYDpjmx9x1h7c2FX/GpkoohdkNnDsWsAQxtGQ6eICtuvZqJ3oqIYCWXbvfof
kslDvdIWViIEyq7XGqs2cYBw17HfctnwmvMxu5PoDsu8EtH4d9Bgp/tZog8EpNyD
Ftazg5LpVU1lP+Qsa/XGFskFoVi1lXTTOHXK4bsPecyr6KEUyvdkT7nlqzL19iT+
Mu4vhUC0qPPnD8dFoF+UtY6VIejlRGPHOA1Kvh9PRfnIb1d645iQQ/Yhkj6JIOE5
jKfah5BCjOZ+OgQ5zWIBN+rXopuElCS1K+QcZq/Z/D3hCakPLGrNGYSiZ/ZCuXeg
au6m2+OWeTElxsvwQ/uyqJWRQkMo0eit+Y6fROAbHOw8XDpchb1jASuQlU1sqrvV
LtS41uFC/YkKBoQXDXIBn6jS0mZ7gWnglpq6K9TOKZz/GX3OLkUSo3IjmPcbaK/x
0KKAx4a70gxHnyZpS/IUdt6pGcVFBt68EKTog6e0nfusn2nddLOzILscUEa6tobn
XGzPljCPsNYi7jdXRYG/K8D062mF2jlad8B5LwjxDC+4nv+OtADjyoUSye/Unf5K
u9BY+rpgJS6YGdFb08v9Z9DAvLNTQzkeqd0pkBtAMUMQEhjidoEnoSzi6ggiorHv
63hijTvJVbkn3WKmtAbxeoCLA1Ul64TV10a6PpbSUwNzN/+kLvGBCy8d8qMFXdOW
OM/RzXIhA7dQJ1xYhq4lnQ6CGj/XOnVwnUSmSds8bw5oSFkZPH3ThjqPj28AXwSG
VgtHYLxKPPG0eRg82JIgW1+omV/aWQYRuOpZaxbSyBrnmtfAP9zLaw3tXZK4IVEa
XhKrDoWbZ3xmcX/1Dz9qmk0m8/Uoe8dBjV/rKeRSLCeqJ0ujpiSh6chgEf/hIDFY
ZNTVosgzvn6Ibi7u5zyKUQQJFmqf15hqi3Cn/KRPaOsXoxYW11XULze7zSyXRKbu
6EHNsbFWOYKD40/gUc7Gxh3Dr/X8CAKZWzHW9kG/ahchGjApF5gY2AUxgv6pnNY/
vqF7km/eKDCQPQb9ojHW4ngRwDwuOdVinSIxDH94JuIbKojR0ALfdeARtPb8Gocz
3Du+SXx/y+cUMgWBL0G52q88vWrkQaD+ScHD9/QqCknovsviyV+rGpQpfHJu73lj
XVeuGFp0y8ZV0j93dP9QMXjQqN4KG8r7j9VMAlurExTG6IgRZpakvL2qIv73fAe8
pQbtGKMcYfhppfXTpMzk4ZhSpCGjRQIWNrRqNcKq6qwNjaQXUG3nVu8G8s0QGsGq
N11k+utROQoAB0WBnssE584wrTW1IO1FvBEm/ce4vhFPEfpaBolysB9svpxgXeS6
o8BECZCYsXnnu0XLYhXCvdinlWyAAaX6peggAiLXEr6jKHQDusFhfzlGRctfmP7P
HTVt+5vRhb3Dz/J+eXFDaiJKw9W7YFe4C68oL4njVzT25Mz2SCe5FBHpRal7u2E/
cZpbR6OFyJNzpQjW2gKhhyIvzNGfHTsJVkloL7qcfnjr32k8RH51ljK0lgo2BROR
WnIcjT/hiRPQfw4HZ11ttqIWDsuU6mCnBvrxp4E9J2ELC9cife/pfCl6KNFEwCGs
ypmtHBHVA8w6e8oUTaDzPsMbAK+PTseSJGNGTIvSOdTE9j3RNcQMZmjKsm169cZ2
YuwUzLvTErb6o6mztRGCyAn0ALRikbiG7XoamB4EPXYwe7qKry0qWYvonNKr8yx0
cClNyQBGth2Vxa3h4CNH3n5lM3kX6apL3pbH9JIjC3/qPhAfwsdkeApMUHS+dPZL
HEjm6ol1jOG2U+0hWjgLDfShl52HfHTCsUwvf8+6b2nclegD6xos+f3FsVeCG8rO
e6nemFRD82t83O4A2+xp+t+fHIjYQ1JnZ2GE4n1+OUfqciYpFr24SHfry6vgONn9
NARHLfuRG8OFAsTPhfCVP3yBGWgRC7XrJYVnyB/jZaew634Fd2Bq+EKdsrdtSkRG
jrvSTzFmabV+nBj7q4A/JhZrn3/hLsO++g6hCUYuFQaxc1ACeLkkDXE/5y442oJI
c2dz3g5/Jia9HoekiX5ChkigTUI1ptv9wXJa7Jis1ByXY6N9tuIXm+mFkVuuQJxc
gLdqKV9Sd3l0kV9S3qrK/Uu9bxizHSrlEk4M7P6LQPcOXFDJZ0iSrnCh+vhY0mmL
9xunPQkPQxnkm9/gYht8RlVyDYK+9zk1Iyfd5baDMhEcIERyawDRex7PSejBhk/y
nX1i9oWopiDbNqucH1v0ah84DPRjcUfJyYpDHSOedrwl9bEjD4uJ+8B+MuhLPWqb
c3jE1v9MF2ulorH8vwigOj9cKSFWhPOiqFXm746VrZIwii5w/vis/we4K2AsbDlW
GtVzZzlY9Cpp5HoWr2iQ+FW9RKp6pAF2XQE7WL3g88S5oB2WKmw9aUMbolTASwD2
jE6ZoyheB9CLwPdguFMd/peQdLbfoar4h6dEvdD0dLvjjfw375pQDLg8rNvzMg4T
1tJPk2N90qQIcDmqOvuD1h3vzasH19eeZm2QHuoSkvdWqlaCbhPfY0TAFgH83FoN
phm/OP9SfghZyLm9K6zbjVu2uxq+SOB7zafWgZTEDJlWV+0+FYpOfqfSq9Hz60LB
mAJc+utQc365JP4bIYyKohLdLqxmxyfJrDDUGW8S9dAPtRR7qf4tZR44bIxtqYuH
LZ5z+BH+bQs8JNS58oowdrrBUXBi5FKLHMR/fRMW2XskvfJiCSyNYb/gVvGw7nCJ
hAIRrh6sPCs2qcn8w+QkLNulxPuTOy6IadWzZhZJwTH1oKvni7LfreYseQOrR28s
PwLgqJ+SP5JU75cPCY4GKtaNZvkAzAGeZAu0pX9FbPEoy0b/UQYrN3XMjxWeDyLq
lLQBAgf2HzeWGKjgol4srwO356GqyTqosZqWamqAZLVCQNDnakisEBvx4wHjZrCb
Z1hvGWWaYCDOwLZFRtkOpV3cfSkHVPlIv1Ob8+ujxwUtIOAKTxKruySaLPkYqmk3
v0J4xrKqYE6RsEm4XrUhoOtvd3T+Mm3RZ3EUkuk7tryEAfTnunrEN3OuqYxIm0au
cH052GKMf88siVkwMwUqUnSOFIWICrIVi9g0kS+MNGhGa4y1ufQ6UzKvyKi8F57q
R7Fh4S0CrsW07lbeZJo7qbesBVbJ51/dDacreXmacv6F4NZ0Dg6yUGV0F6BkeiM2
skLPP/0m/OC6MhHkiiVa9S/pSwGBmHnk6qf88/w4lxzXoFQHdKSAENmntYAVGoyN
oQ/exI8Sg3ods0UKUdXN63RVxkbNepQUeBEUwVPOffcH67aecc5Gg03Aj/WCSfto
BJ8bcnnzze2DTm3+Kn7eqA8GXueG3oWiffkEjp7O276IvK+N0wTADNzFvQm3wRbF
RwEzA524AS/230RNw3Hs2RaYlVR3JPqqkG0udPXL5fLwihc1pvwER2/k+3i9eqgL
ZwCOpyrrwjYxPnstplztLe65d4uKUiROgCTWSzCanPsc6OXgVv0Zw4f2wvX0R5VS
yk0JowravgO5vXre31W2yHgUaW9vQNOQGDVrm6MXpCys+crtW2B9w9rNk/Og3+v8
nG2Lulwlk3o/LT4XJjgyF4TeZQYTpTbDjRWpR+e1se/lQI+jLUsEEfyTLSPmzoDq
zRe6gZk0jNBXJKEFCnpnZeqXi5zDQ0qlHgaGlvEMTcWOwZKtkJZScNRcq2Y5s8uU
bx1ptkyMMWh4SQYUMFQUcif25UHJwbTFnyxBBaHiYVjk1PBvauHx0zfiM0q8ruYo
3i0EyIKPelBcym3TwG0IFb64i3hkHRwCwTkUP35GYBYYw2fLZNNLEGAThlXNJyJg
Z5fmhDHc0o3kh86zmNsqwlS3eqP2rUiFoxC47B81F/EENj8IoT4DE624RM+GMZbM
hYScdAhv11u4YCPDAhukqaHnrhvMaqJzrjqwyBAi4yTN/quM0foPfH4FJomSN8/O
LMaUNbNySuPR5Yc6+H8xW9Yc5+IyFk7KAHpR5OlPcevqHXPPckwpby/9kDTtqhpf
t6Sb+EMaLy3JtQeqFmea4SFvX+i8P88mNr0lOMBhs+Mwd1ucdpQCYbYnXWMDpsb8
SGu6f1haewrnfBt8a9GFvlt4G2O1neSZfDpgzDyQRwcBWKEjKDA8sCXfeHk5Bim6
5ClFiEA0ElvCDuH5GEKrrhVC82iYw5cwLyf8AKDqIISf7KOHcIlEv3lJG0QTXIlL
fPGsEEHzpmqh6QF3TEbcRQhGLJSEicfTyzckSAxVFrhG05/VuPUKJB4uuA6dGxoz
3pRHXh+w/06VnviMNrTbtS3jj7PJraF6H+YctzLJ/VTkEEGUyy1lU1t4f/uk7DKT
H1SRwyvx0qWxXf087XGF/ZGe3eAGS738tHhywjwwNQ0ZSX7kZAf38QL98SF/aUaY
lr/86VnL+FCYQ7ygsgX6delXs5/0IxxP8rpAPFNqh9EZmwXwn4NJO3R/sXBY8jxq
zA5iE5/yeK2Ewh4Qeb9hEnZ4qJ5Jek1OWtcCX3QKZsMsG8Kl9VCa87T4WxDuPFRb
gAk6gKx9eHHfJuObFF+wDoUZGkuNQ63EFtsY2Vv19WVAHON6k8MzWmjmKbSYdYaw
Yn3xDTxzsXnMm9fZNQM54ktR1jW2aCCNJgQ8lulTFbon6msdy1mUpGCNbK4dRZ1Y
25fUicilVwMOFNR4gFn6+j8cJmGUUb9UGCWN78R+JSYtS1nMGPpa9/8YnJ2AZ8Dw
nO0jfnuiQXTYSNJnYDkX13d7lpUKPOqG2RCAFhfZTnVL+tkjYm2XPbYRTqi+aswX
11wcQ+I10iagUngDNP6l52Rg4NRkxA6t9gb4eAGru5A+0Yxnb5TenY9TqHPOziC4
chsV3PHjDagUlsbAZSsmdVcubfxSQPQKeQ0y1YcFYdrKplHF1pA/Pa++pRsCiuEh
9GccjeZMNAMSqKJkY0Sfpjqyl5T41Mlu12J7x9tcJojPqHRkLQu/YF4kQyOr5mHV
wrRQVgWm+7DbdcJ7WmGXg2FSw2gOsTpX+k+ZbA233s8N63vuesmS1sF5C/pNmBXE
sL3s6Hkz37lA8+HDSlKmuEQyUQAUqshVo0Yg3SB9GFSgzPuAr8m2stEjJJWWhAnY
3GME1Oqwd9Q5rxstTrZgA1uIpD5SQI2VLNHJvmQz5NfvLXgQLtm0YobZQ3+tNAGu
aAvjVhrZlqFGST+boiChfI6IYxekJ01OtxJfiy4Q5XXXmxoT0C3tGwMYstJPQrRf
Xj4dCJxAN5a6rlW3803uQmH+Qq30/Wal89HQzWtI1z6oikPlZp2GKSLc7om1/hm4
fxgylbtpauzW8QLLU3Erj+yOOCfuux8Wuh+qEBXFj7MQ2AxpM9tVpl9fNGinFGoN
ck8RQ+6MqvBHQUTHnKYRxapgIA8PezWQtqzkLpWPL3ZSrCI7JpEuqz1WWkux+OD/
TAoa6LtX8Ijous1NbBegdfJyozXVPqWY7wfM2RT8oSaRBGnGzDNqA6DZUcO5TvdV
zc5o/bHkH01ZOwWg11SZ0IatryX7nZyu0PjftKlS31f/RgebsE0DrKIbFZd8aKyH
cnDym8qbl3m8synxtqw+Wwme9uw/o6XIcwosfEKLxBliiOy+teI9DCfUOtOk3BWi
BINcnyva17/4x6H/MrSpAxzPb7TCCjm+hfiLxx8Yd9GizCoH+5L5wqmbked6Xdlc
bQA7VHZ+uokgNsUP7cdqfp+9fKZ0kXNrOxZj07g0wAtafa9Aq0m74O3uvvoN1wrZ
IzKWN4gSFdsHdxQmOJual8vpSPiAf2j5rk2SY47iX01WpwVp5nZIZQs8BJf4MfDI
w9Q/RDAy2bON05hZFbYiy1xv6/ThnqKXmmxlgF15TL9Rj0MVRgp9obby83TUusB2
5qifSZOoJarWNWf1aOKxduS3OyYrIZ08Q4Km1Zdhbe/mlgokW8jjlIOV1Od7FGOr
y5h7MGnpqr6LXz2Zglid5CGxERNQ8yKV/tDupT6J5qdMOIjkDnt8aSgJpAjg9WTO
EolfXQJ79CL4HCJJREw1JzjtSVyvn4Lt5yHpCI3PELEl+BZO7HzALrEurRbooUNz
QOpKWKOCQ2ilJ1jOoedn0QmyyekHq1FC+Gpua33E9EsOJz+Sw9+ZkW/DgMLs45vx
LhIm7HMF7ZvL21Wt/1xJcy5vyguQWNOY1sZDAlawOTAmPd9IsU7DkE4/Iw8yC+0y
b5ptVaRytMsmzaqKDbgzEt6lTltS1cx+DMH49i0LkeflwYigiLQteHsINZuO4KPa
Rdb5yfA/EgsK6iDvmh/fEKd6udQE2XLHem14wY54xaulnU8j8LslJJNOR8erPDSY
q8JvTEyXnHB4sYvtQdP42Tl27yVTycYWlOOCOhGsH0mtPwNutXbXFgWXDnfSejyJ
APSWcxfDELdWSvhC//8nDKSLEKZhgPSCsMQAK7OCRKTGVjrIXMfYXMMOZNfIn0O4
A8NiTERTmaOF+V9T19E4i+A2Zb/kqbRr6gyhf5qdHK39qWBAHIYS21cYK1QUYMRK
st5zIe7GI7qx5HXsPhQ5ID8OCq7nB81fm8EvbdJJnSZpxvaMfOPFeZLN7tz6DuqC
6g9BpiPBtwUZCOLtFfC9lTY26tNAAojyrCry00dkNzFhRi5i5Ga4J2caW9w2wqls
MXrx8WWHlnwwJgrtMLcJj/npyLXYlr7joHwYPn5PlLx162TEy6KN8ohBGFSzCBRO
QPrfMyOaEqejl4l8U92vmKAvrCoFFklREr5/DdUpPVk+FmYQw9OYjKNEvGvRZzGW
UjrzS/bRV+MU5yBVODQKgqXfsMWnnEmMGCd+VT+weMqY86v+UHGaO377fDJrZumv
bmfwIeKI6ZVztaW0KIjUGp6nh+H0ndUHoUV1jjGVTdPGKM411UXv7fVeu+G6O59l
fPMb3I/6rfJ5SgxvGruy8Hgqv27tbq2vMlsDwPxVu6vq4yuMf0AdDQNDXZ4Tfd6T
DgAp10VsUyYCFb4+LGWpN/MrMUmFk81hmhJcng+zcXK54iq6mBnKK5feunxQcFEP
ZiX3AQElNed8c5FLGBsFqvHmP9JE3eFed8bbTXhUXTLsAbwxWXK0lc7peIAwFZ2u
xPGNhyIWal7YsGJVeSaiO9gcbUlpfr9BncWZhPGT7ZwhZez3WqsgOZlgVT2zQPzC
OXpLyFnUjP/MhA9n8uctJYa9F5DkfxHhQu1y41qWdUMDSfX8U3LboNBfTB7SjFkG
XAqIkA7y9uu64GNde2qlysSsZW1gBcs6iMU0juF42y+i18Kdq80Skxrr9E6lig5u
TSHloJY8dWZhDjswNZoxYR+LZVMPvNFxb4AHVr+E168s0GOZNhmxP537TRyHD7bS
bqKsuFKgEXNoj/eEk0iO569jq2penxn2CaMmGqRFJlH+NIDRLqT1uLpuGbHz0OKV
s/Y3Im7WST6Jpi1EMQVnbkX0Tst/fLigoCQyxnx7fnaNfvJifUp4Q5JAN0ikWRcB
i6JYIMfglDobNK/6AOZfwxR1UMFADVsXC+081B8IKgfznOsU7A7lmEhtKwj2UvVL
MqMuHpZKmeDskGGK5M28sK3FEIkfhAdtnaJH22PMBd7SDVIRO8Drk+IxD0aRowPx
nLPRIKnKlZz8CI2vzHHJU/vTyj97gS1YSV4qdxibpIL1Shqb+2TcNIE3R7fWXP4a
qn/f5mNTtuKHtOv031eUQhuYG28NmQScrGXu0Bad3isPMDqThv/8DL7GLAcEgvD8
RCg4wmGJpUoWfltlvWsdwLndyvW8rfNRktZRaZRSm7ojXKTC3SVk49ZB12D2Kj6D
UzazLWigE9Zr4NLdyWZdlfhPuZanOPd7W8cMPsj6RlkRtqU66dcC4N2wYTU+8K5f
JZDPjkiJHsbO8waWbVf2e8uE9NTYj6uo7YfEUE7EAGqWp69XjY3E46kEugOh5zGV
5hfUXwSs8HTdNclIdZR3rRBF44n3J5XbvHsHjvhlL3qwKbEKSee1ZLLjHUta5viS
OkW9QWep+JafTyeayfCDcQ2KW4/xN+ctJbew3N4S7ajWOd5nxJBje25ouxJUI4mf
KCgYKeUlhVPl6W6cQCH1qSKpm01EsC7jkRjpGGuwY2hcdma+IVLrlQHacps9KOav
wzwfY3QUnDFrd6tD+rtVR6SWUxxfo9plPAZEa+ar2ifUIkyE3WZIVoTKS1dHrggT
+qEKlEHWCY6Xk/R86FZf6WrbFeo7op2Fu8wr3Ax7IbexyUnate7FHzd6dwv/8RUC
IB7K7BTdHWQQ2dZsArvgQWCuphaht4DMxPO5asNKyf69dI7bIKDnoohaSIdHv2++
Wg0DSeGDzN/1sNZ342Mulz5xS0UL2ySJE/m2uhpb//5iJmTET4RSQLM8nLR3tPFZ
mVK+wIKe0X6dHj7Tkrgk6DIURb3ccMQX133wXyqK8l0ribOxKP/VUlW87JWM8Vy+
RwfcnVoanklbxvGQGkD8ISkM5e7HlEkv9oZDMkUTCaWXbWSFHudzAPT35LvbfD45
6BcYttpeyeRDsvInCRmDTZw1Mi6Yao1X7N+X6Ia/cxHicVuH7AOVN+t5tgrmZI6x
GOx/wu3pseXxhFrcn2w5LLlheZyqQ3gcSCopCSVRMOvLd49oo+aoTaJys2okMD5C
WnymxY7gclgkmPqbVpAd89XeD44+gIgx2ENkaBZN6XylRMpVWUw6hnZPb7xj2lh4
R7iWIN5JEMyRPj27UIrG4Ve/sQI/lAGOmyQhC7uKM8SfGLxCMrAGBIpwYPSzcxd/
AgJTlsYZlFCBHgHjHF2y25yz/+wNokawKG/H9cXyvzkOK+t5ktOWW+cFrqW9mpUf
ofIO1eYX54R69N3hjrKPFHiBooCf/7LeC5og5OYnn2mWCqT/IdpLiu/MQeHz0DDl
cyqY2PFg8w16wCRRlExW1DW3npFlSKsyRMpRCFdhYEtRhol0ntwdrtXVR4sd0m0z
iuWUTT2+C9+FTN9yc+DQs/r0tCrMKWC7Sa6KOlFFysuSS/QynhVt9WbKt1HuWh1N
jBjakxIFyPq7vH3CUldW3wHUObN5SkgFbaIxHuav+GWKpG9Qv0AmJ3WLlGlqbHzW
CHpdCZ4OAHo3ygtOhSJxGswwgzUIRdMwasnUvPkdMdgCm9xUysMi9Ul4nMCxIUVN
dmca4l+/zAY83iedNJ4SGFh0lG5r5T24VU9LHBEFLcrgPgh+v/2hjDt3+oaUOc5i
6zNr72ZiXRu1bPhNBxmWiy5qjO2Jvhgv8SDkv+dmXdM3XW9F5P13wjpdNol/96LF
M00I7LUt9WnBHZfn2wfKrRtuE3VwpEB9HCvo+WfkNu3U/VE3wnaz0Kf/k6pw2nfp
doc/12YA17SoSVMXZoUUWN/WLb281uPDSJOV3wsxN2G1xHed9CG5hfYe7lS9GTQT
C0jNQvGcKOC0ynmVK6vhkMsms1nZ/LwTKqiwg1P76gn1AoI/wDc49NG3d4b7N4L2
EbrJbMqq5WYnsulD7nisUNsUCRDs/RS34oOvjsY16c8TVa+/L8hwwJjYo9D5iJrT
2RsxOdEGftqkCEOcbnRdTXnHqkQqbcMn3HiucTCtoRBbWRftQd6VtFUrO2bUWlEg
n0NLppcwMZdxcw7A70AbWDvrXxf0XICDz5xD2+QrTlfYLrmhyYoy34BwfZ5CNOYK
9ZfMrisi31xS+IGRsfaP9ITeEAJEHr5eS59pOs4ibWGh+/sCU065UxihAPHj8Kw9
1b7bcPuDYS/+K2jReTYbYqo5Mp3wy1ie1VtCYksO8YEkFTGcYQ24yEc6IVOKrTOu
kimzvSiA8KpBFHq4MPh3NTmKs5XPuYuxeRjx0LVWpP//QWtoKSRf2ZJ1zTRISCMM
SfzrCvAUX4ZYPkQyxHoIm1awg8gCMvHTha6OZRF/fT3nm+ffZMTkVgnjpSLSMk8S
pXLuKKiq+dHXl2JvJrgCZuuSeUF9g4U7TxTsGGug4XJVo8VcCzbOgr4YOvQE+33o
DrG/jbYIBw9LN8b0nYuh1bpPSGDts4hFYEtVjW8P6XWFAOFdNEUsAxiaFLC1hHsK
rh8d2sJqOjOyXTC0CXJlYpBYtgIIIsboDpCpQeldF6haZewBXy9zXLS+kDigmhSD
Fic0shb/ofsLojS0UAQLwN3N5iIDpgDcwaSlIw6oWcthAdiwb39BrFchBE+1GMrw
CTXWUYHx8hEJ6tmCSU1/tevQJY1a3FnEnW0yxFae6l2Ah8nCffLxxX+mOgOtFcwL
wgUh3FY/UwiSDDTo7Rd7/hu8ZjcbT6VrXS5BnsSjbgRGlKaPaztJJL/C4EytQt9r
piKud7GtOk2WcNREFrpNauZdIfSsvfDpnllIwiBqjwE/4bD/mEyV/SrQX1WLwtec
zVKpvLQUgLZbbXIIU/3IvRx8KP/DZfObQf5snWzEjV1QHK+Peb1ibPPLphm0QlU6
yxt7h0Ppwid35gYO1H1o8IDDhjCEx7tNqSIqi87gmFFdegpLfE4EGKyeJ26GwT0K
3cSUYObn58AhAjd+ii1k2uUwT960kFSu5E3XvS6SNJIQ+gneQSCusJT4VFsTtfxg
A4gqkt5rxyosanQ8pDjuq8qPqBkB8tXcW4T7fL4LqHY1FQMWZgUNg2XnFLrsXuZu
4sTdkU2xZPIrfTQxYryWnYLfCf3wQ+iwTDRJHQDxYcz1sriIsBfgDD9GP9WplfXu
jLFxg5XhMbMMjbnYHBhbaBPlLA3H9Dc89/DiJQeYqrugxAAcM+SujG+BcvVS3n7v
qy+JJqouhR0KYsAQ8K8Zcm8SazY3/Ss/jj8osG0C0UDMPvOnCjEn3Ufy7+ivDx7r
33dC1OPFVQKhKVVFvowr4xAEWKEHG6WfJwbzQTcKJZSPI2lc1q4TYd2s4/sp1h0b
MM6ptWp21yrWXh+lMgLW5M+hxNOLR7SkUrqE/zx+XKKS97KnzHpZzcwALsV+PJgQ
YJc3j7dV6JUfHMNQjS/yFYyT16B9tCof6rrPOJrknv9RT0dOvOZ9s0Ds/9CALZWR
+Fjv55gfJntMfRz2uwax5RgmT0LR7ZRl/ofnEPc8LWaza5TpMbF5njn3PwYBTiKp
y5u9ggCCJMoKcOwl1dsD5BtN6aVk+H1tF3pArzkZRProzggTdIqHdnhXgmBgVvy9
g+Q3ogA+aL5dIL831OIbf5u3gYPb10EeiY1l38LQPGVa5jxPDZHoHKM1qKP6hzXr
Wi+bU1PAyc/EA+ELLWVZAPdvis9cjvVFZ6Z0SaM8bAJ9+TDKYEkIdt4w0mJLr4QD
EtNS1/wMr5H4k7SZ4Bm1iamk0WbYCGQVaBYC4Ede+XfRdn5eSVaiNlZbpLNfPu/u
8mrX7dqO9KECwmSGo5tM5ibxYbVdxEUzzy8epmq5Tzizzxrv0j7IGNyReo8QHGtV
HeTgChryVLNkgUAlZuxRj1kTdFxKRidy8I3ba/JDShGbuMhR6SnlXYKpHocIS1gc
mSVdlRpRZp5gDV2iRz7py7cB4XNHBtpnAlXJKrJThM8=

`pragma protect end_protected
