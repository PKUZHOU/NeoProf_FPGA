// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
JZNqLxR9c1TTb2i7y6fHPgWsor5926XofX4pL8eSk8keWV6MI17EDC3VZsn8e0gn
r27A+9M3cBeXXIW6p2JGpchHDIcDq5rPQ1E27OdzehLDeHiMc69xviSrT4maketz
A0NMUzT2UDpfOYHdjpMZCk8GkWz+0vBZcfgsYJzXqo8=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 29856 )
`pragma protect data_block
UWLMRAUhQVcvsfsla9POcFkdMzpoNnZ472C3IX0EsxY8qi1CIFB4ssOv5cfj5o28
Zxwr0ucyiU6vExTlXhN0OQG1tPbttEVv5tUTSDc2mGBI6sAF4Co7zWDrYCSmEq0E
zCYjO5VwkPO4BDLT7dc6LTg+5BBRYKYnG/AFgahkjkLX2VGrFe+xUX0xstKDz2tF
ZnlCdzbEDo4k+ysfFsKNC+n1HsDgFw6upKDPGDLgEc2Ipf7+GlDwgTNpfsKjOrUN
easMfBGFn3pz7vOa9RcpRxXK1UF9JfSczAf1MreJJNQAJ+pMB9ZEx76miWYRemDs
HeLj3KFiU02vqwhubo3l0HpEWgGN2D92TgIHMU+pM/LcOr8OBdp5yThkvMC9bxWx
dEuzO2TwCS+Z4r0cOQQ4aJpBn8iWmDDl+k7i4ZO3c1eCDy4/HQ6VohFhjJMJK5LV
old3SIgjPL5KnbjzJuoyby2M/m9J6IwbVOde8tkTW8qTG0U0FQr2+dfbQWkoX9Dd
7dII3srJ/sV6XUDC4fOz2jTOloj+Q4ETfzGVecRLbgjGFhaswJcIKYPRTHkchJ8Y
A+nxIX7obGTqhmc6x4bVwyCBFILVcpKzx/OCSBPsG7y0PtrtZvj8PqayB35tEX10
tdQmSa4srDMiGkUpAFuVpVkDVzOVncrOP79SrNqIL09msswyIKcj1Go13JHFUd1+
Ehgd+LlLAzdNcwZI7pubW7PaZEXONfwxN8vVIapJi1uyj0xJnmO1uuFGARMezujq
tN7T5GFitc7eEPE2NNnOQAK1blZV7U6sfDb2wWgBDD/agCQ3kCAdHs1v6WUGUEa+
PjV91sjb+NQyQGIg7W7r8G4gOMyZa/FIqs2g9kt7ff+Ev6WyoYegfvTyz1IFmp4Z
Z3Vz5LqMUQBAmmlD72kN3o8ODcjFmP1bRlz0QcK4OLX9JztBNrqvR0uWVhENX0IR
uCHI60tJisY0aUmC9wN3qF+EjjggxfeTaXOehP6Nbki+VER14R7bQvP6AgTyOEPq
cOIyj4qjx7QLdXFuHUXG58d2K4Gz+nlzY5mRIW/TtrmXspftMJp6ze9VD/lC1lyr
mV2j5Z8Zw+fgLHsYJBC5r6tqpva6G+jB6amrSPuK9igNR+/PzHeIA1qOG94prQd6
ZYMx2bJHw1l3wMnzPTuaDHsDoYlhu7e06AGZMExQiObDe2IpDpIAcXzP9SJRT9Pt
t78tosjD1iseFf5PLTwhFMvYaMrwMoY0jwXihLVo5S5DUOsX+hDmcGa43QP4VYYz
9gEyuAAwx8qQuFhd+QKhYWRSywR2tmwkQqfnU39JXDfipJnwJ1MAKVFGmcmpweyI
0HI2iKKC4I3S6CQsFvDDi4nu9ihdRr9ZYv93omk2UsKMqpQrQ42MvBZa6HcnYq0y
IQBNiMdyhZUIifa7/FjztpyiO77p6UG1u1rto2BBiEoXSeWM0c7l4fAuqDbjQCWu
/tAvP+C7rPdcL6ncLY/hzmx/Hj2MWOONZmmEZpe6JyhrVl1/9AGkU8evFHxVfC/T
PjTTcAL7wqP5bzsIDsjiM0rgrkdX0DctOlSFinI77UGCLCm9HBbDJqbIQRnn/3+i
8hUcYD3j+GLuoqJBmc6VNdzEjhWwoWS+vkF1lAZvB8uXVU1Mf8NG9VXCiAiZG8Q0
FnYwbcM+uDL8MWNkVDyNOib0BtPtGBLNV6cBRCqix3TLCTpUfqhOV9yE4cOiYbdw
zOh6YKKo/odiGKj34rVo0qawgAc9YN6tMglOiY9IdCAuEmxXr6wGarhHL+yT0AEX
csE/OYYZ7q4fiuC8fAhjau+QxZEhUjy9F5AA/YaEdU1qep1jS3b1R20tMA7rcxoU
7Ez5OnuYzF8t+21twcsGddsFD5fs8K5E19wL336rELJV7w3KrsLiLQR6L0pUMh5/
60Q7N+EF8PEWSEM0cJSIroSJHCv1yYka8rDLD6D3Xgx7ApMFhYQbgVYIoiYUgvfv
YoHosEFLQZUZRTnYduW2oVzbEvWVSfefB35Pu6rbG2qDeMCtitZVZZXE/7QEYbo5
sxweiFufTJ7VXrA/FBx2nr3hi4OnD5hn5pQ4NB6uFqGenfDWUAlawilUUK+KNNBT
XHPHsF0SVkUfg7sAurECt/oA8UesrnEB2m8SC1pC+zM1AOAXlkbGm7yugFby8+qZ
dDwpAoxvosDWCoSNnmcbVy1TLz16nQao3sN/qKUX6DvIiTe6X4vMdhcKQIuTVQTs
S/PwqyAv6+cm4fPkZY8oXPpfNVYIJdlxKok8liykKWp8MVefDOva9ZYVZTC1TNTM
2Ta0OGr0xRYO+ZtNHuA5476igI8gBrKAHw2mcEGPCOYg+EI6csIVY7V6QVXsMuXR
1N8XmySA+eApLI6tshugQ1jxfzW545dbYqEX7ybnDy4+abr8cCSP+OhSZmx+PHaW
L1+ShKTJimWTiFyD6uqlC2hSA6aBOPF6T6M0UUS0OiKgAA0zH6iI5giiQk/YrU6n
jCTBntC/BS/qt5YEUCA5PPRSXmEH9MJeRYjd5nXZvdJ8bihNksjbzG5v5sFseZJn
qw+H+n+ETa7OKrzmoDUrDtI7e1fZgAa1aUJyIVXzDG4YVgEQj567gPmzcQntNWAz
gRx9S8z2ETjGlHQRdojeJ64iZTEKSVXII1oe6D7bZYEBhJ+59K776DF6Zqyw79Bs
n6lFxsM7J4sl60uYTSh87Xz1y6g/A7mMKbJm65w7nfelaAih8DWph9dQ3gr8LoIN
rTyuS6w+8ONt2jiD5k7t4jld7iNQX8p7IuiWdtlqExVejOkxaQwAIEpqD/KysAo8
iER3gSbgzLUgFVY+dVjLqZuaP1OHK7/8ILarsTbyO3n8XQbh4usDWrVgGPZNyoS4
W6DaCle2QcYkdTGBQVTN/4uvm8gBT9NtrjdC7PU96RrgC6ZlzUFjoDV8i6uX3QSd
qY+lVrxqIow5aRj+OxUto/UFA9SAjjflk4HdWCniaF8WLAbpxagxSy0tbITCNxXN
IPFSKFsd6sdIQzgMrcWEeX5TP8DNy2f6WhWN0H2yS64ZCxr6SYtvThp/sICx7j9s
RdKcweDchBixePY4Vpk5k2DHtUbZDQFyQA1uEc2Xy6LEbsVUk2gQWnv2cR+6AUbg
glDTz00x+ypGcRqrMru6T6+tQH6s5d6j4eXDoJb6TE+i2gdy/d3ylOVcearz3pq0
uEi9aW5aOnPPNHp2qBZ/u1rB3lfrwav24GJD3dB+dGGROAiwifd8QjG+cfy3lOb6
C5cWYEteQOxHyIMmUny9ymGYDHti9cg3/6UE7itJC8DnNSOHhpmdNRRX/1C50uH3
uq4vUmQe/RyfnOModqapY4FaHTUeAw6fO4iUflgZgmGatB3Z+kSadaDn1UNbUUg6
ATYTgnUwHfsMDFGPlSZchOubS0SoQVaJQvoDLxLyHxj45SyY2SRXYCMrRcB10aOS
gXDVDmVpD7TWl4U7bQ8l5OCc1ucz2ZPEtN3vw60AkgMG63brGCqHRQPqvAEYaL2o
+wmsRrgLydup6Lo1OGAxhhsUDF27p7coopdQdcsQLbWsxgyQUXM/vstOTzKfepDi
dTKXy464hEHkYl1BmDRviVZhtnwrzDr3JXqNY3pSFTSBJscqSPxWji+RWSIFEMOT
cII9VODqJVJNkaCCt1Wj+mYJFDJ692Ukh4Pa4fAl8CR6T+byZzQ1qBzMi3XwFdPl
xO+P5rmkTuu9a+25wM91CZ/1J8QSH63Ykx/cD9jQK/fvOpU+kG6QWyKvNbQWxfyr
qZXjJRqQ4/7VdKCRiJTr98CXO8A00WNIB8OBmHKxVx2PEptgPMNOcPNdo7Fz7N1W
0N+qk/0WonCHhcl/bLjqFqHAYbw4RV6zLN1sv3XTjvpn+bDSm6eOA3SOcP/pDJNn
CUrVL+FE3Szu1PLeHTSbKZzpwpmdMPDM2k3iSp1qxuB8e+iG3RXJUjAdbNHd6xD7
W7xLUT/LYm5iE8BmmeWv7dhVAgGXUJOzv4OrSR8Hn40INzUutgTN02CisGjMjEyR
fUSviBJpk7GpoJ9ww4eA60SaIkfTyT8oK7PGU/Tkg8/9Gp5U91gG3yJmWNIEcfTC
xs0vl5Xp+ouaIr+BsFXZCgYX7vtdMkvRg7sfdIK3vQ8Ww+UqaWhrc4wEw1Xp7j8U
3AoKZper66eDLx/FudmY/pTRJS2GNVtZugE136GyiUQwhImE55vaWKbXcQwY8+lM
NADmZKgkrd37OwTyHltFqlEYybmz4bxqTFq4eY/pSrhwe4t1Sj1zTyLiKyuyLs5f
ePBAscveempnjnJ5CYSqDkv9mfZXI7bmsrH14y2YZiUcHO3MMWFFuN6rFexlZztw
fad0YQKIuqUzcTU+8ewiTItgYSfZh+ihMWfHY6ZqQXbhPuYV/vXImqt4iKYBqBOW
/XfutLrq7AWfBLwR+RrHD+3q2tUhlBMzckvudU7NbD9CCLwsvZD6cq99cQqUX3uQ
y22zj6GvYUemc1zQzzKqbKdHzHCte44oJPhjYgKrwu65r1YJ3pm757diS6NvPzuw
3ehyatK9ScB4xHzWmh5vezQ0QejIgPYr6E904GWuHZfkFlNwigwopR6hfYIHRSmr
lr91VKmj2+xY7IuO1Iq4Pxrd75TPwFQHqn036xSbt8pxD43PJnZU3+Gv+LhWMnVp
vqHe0GF3bdeb9o7Un+M2B1eKKJ2cQ1QLz0gNwWnm4kvw3K4D3yhQGyErVHxQSFBR
gJMN1NyKu7Fz8ohgbGEmvfwDLeKqOqovGlv+rcA5HBQQ9hH7WMTkW2KfNCBNL0Hn
L7jt5IqIjPgRf9QegoOocnvieTYmeF0l5KuHqTN3SHVSqpjYeM757CFLF1LWDbso
0wWhBsfL1sM8Oa59Q1mu0RFGQH1qzWMj/WtWUVz5adOXKj48J3zmZzsV8wsmXuCz
b1vyEo0VaQL6oHp3D4sPs4gfGfZx04gr9ClCbKk9SV8wac6uBL2PTPue8VbODuzc
7SXrl+mdssi5wKJTShM1M7zT5iggoUzmf2znKTH+ceCf7bFPtj656DP9B5skA/b1
HRhrthcRUcXn/Eo2uu5cI6l8nzM805tm9WbGr6m6k9Y6VvGSV2D5BN0UdssYDQUm
cB6V3m3/w4EgKDDFDXzYXOxj16OLqoOpcUmLzdwBVawnpEB2goy3bmD6Di74CcAJ
Lcj4/hSSVqRur2WFTeCeex3l0CdZw/lHNVtlqaNTMhJJ6EP6vBHaVySq5qI2Z/4r
HcFhaxEOFBCIin2qKnqZ/i+sCNuqiX395HFB0DyEnmZ3EBCKgUx+nTe5Q9YM5jPM
OH/4kxyYmJ3wfuZy2nsI/fQEWSMz8STdeWdhWTruszzlG65ZZQqVRHeH9GlrsiDa
94TffGJXipXP8zM2GAJ/D43vccYGMzchzUc9weKSuDl5MlLi7PNtqge7SILIPq2X
9IZ0gwsWT+1CXqAjgdIa9nfb7qjc97zw+8bVRkPbZhQTDI1zwt5mHXT0I8AJurFw
2UCxOigLBD94+1hwRGj4PEnD6ZvlOWNmuWXpOvlCxN1tt+1EodnZEW6/OOdNoShY
Z+xffo/XqDSl8v5Oycn9ee5pNdt/K9nH3XeAhbiUdTzebXqNtP4k3l2Ipgc6U9EY
DS+i/eywbhEtSkNDsFlB+NRPR78AB9yaRFI9XIuwjM50noKDMhLtGGrEIrd9Ptc7
aPHU++dRqPdstgRnayKo5iJ0dWLUpicSk7tZ+HHiBJiyvs3nr25SkYGWeio5Wy6R
yh71p1ICpWZuloEa8m8t1nL+W2kZs7sBHIfHEayqalmRrbIDmYNZDFTN2wqRTnjD
nBntNAp2L4mMvQiGsOh04b9Af9ylzXi2jGztgR9e3M9sP/WU9D0SZWy82TBvh0Xn
RFHd73mQet5uwk5bcKrzr2yVqafUiBSyvt/3D9wqULGW+p8y1y+v0tWerLhZvh3s
ZtcCg5pj6B8v37biWeTD58YUFf9YuceA0sr/cbhf+Z4ojtZq1CWYMHdEA/ZC94FM
OwG9Kkb1ZJQGKyWkhLQML5ICIAfiuT+YpsMZaypuNVB4ihcgBe/a5RpsJImRDQfS
Pt9wDAFzNx/COkU3xWG7B7kJ1LrNyR/nleKe205IR0pPKyz+RoYBHxqsITdUEEqM
lah96P9snBMQoPmJVUMeInUyf+N0dVIupIwOhYvv9Ryg/Ztp5qmD/z1wjHWxO74i
BmrwpKWpwTECGHJrR7epxVhwVMVnWO2YoRDgg47SJDqnvV3dX1cM+qITOQbmqVxe
DF2G8SphKT4yxj7iVVtn+I0iiqeQsfUbEbwki5k5uJ/Xbwc4tgnrpIFqNPs8Dv5b
alhN6DKhbQAn3uBczOdIX2sImlHrTxRu/ZGviI1MYUL2eyZV3UgwsKAK9VoBEl3Y
gHDmA5RGS/7hJOO7uTf6iyY2MyA6mhTF6hlJ67Bc8Vj6HkYyrvoasNGUpeO3GeH9
inp5Yk89UQ4Gjp17YpBBmImu+hZacd8tj5O4yZHP3vIWFMJhR2Kuuuox/2IIQZCE
Aqjm221EhpGKJZY529z5vC/waN7NraQOP3xmqsJYUkTXNnrULdTfQ4YLRBORuGCs
9ojehwXmY+CP7t4zP7UpB8b8+YfXm86P0FnpyMlvGaaUToqURqdtMu42nhyHpBAb
hVEZsRbrWuolUjU6ewm2sulaN496qQ+3OY8s6CJAxYhDMkSUmf7fsXoTt6sg2LK0
6j4jbdJIWA8dnioDozlVv+kFcG18/9vGX9ottiyOp9LGvv31Y45etv27JIY9vY/X
EppSy3J/UnezvGGW11A9a5JNUyatCxRE9UBL/wpXZPr3gB552QA+4g4ybvKnb+/t
NE0uVuLkOuJnq2yQrPeKiHerLRm0Q691G6OT+g7rMnWZP5JBB1asdZnHdk62gV4k
C7NkMNIPT7fmAw8QOg6ovJfVrWxCl93DCTdBJCDVimKwEbRri9S5h9saaZP4dVVV
Xc14pMzURiPGF+BKTC85qmn6N7jJffoznNpFXTARPaug9GxnM+sZTgYycriG3I67
C0/gkCgaRPeUiIwg08TQ71UrLqcfB8VDHJMGpZz6zG2Z3D1HfUarBXMiZ+n+IpeP
2fGAb7M/v3J1eHjb4SgxMqNOijkqv2Tk6pp3zhzNz0PpBRL9KFfCOn5BqmdnzWyI
XL8NrzmS3nw8mQpuFVidQS0UjDBrPAqAL9vU1ANGL+YOSM28IbXrjVa4g3HKwJ0+
qOy9yAOQJbTOUS6ERXBo6BL6jhc1v/REiSs1pixjDfHkA0esv8DNTWYb9KRMNO3T
90owV3rIyi+ff7ilj0gDaGKxPDBL4X29aqkhT2/2y44n3ctAwhygLBHCTk67pZ8O
OnZ2JrdJ4IFGm61501AuHPo3M/mBXsmRJH4oLmLF8D/nI9/pisOEtKgPNnPmxoHr
bIQ6yt7SoQ8se4IfbC4xC10c1Y3GH8ZtqQyQcWlOGOV2DGKf1l0PGe/Mm/1UYRg2
tN7N4+S/wV3NMH8245ZnLsRP79jQqZNEfnjuu4Q4j1MeN4oKW2I6N3e1VD0XAPct
dgQ2CBnUNunU4F2NNi1eHraIZCop6hBlWTCzkmYgydIDiejMjqkq3PSMM7jJJ8iH
4jqRC56qbjT9YgVB8+SIPpmbzmK0SKWh1Rk1ZUaFeQeUPOvfIS8WeOiiXo/iEGqI
/t06e4aL5QWqrXw+yaLLOcIQ1w/JbKWaoA3HRfsz5/o1RNSTxUrvd4LlXsYGOub3
UH16NCd57XiKUFxirgKh35LYvKHj5uplED+msI5X/9BarUa9UbcGn+WGC6eNI/Cw
i2ymCZWLMh+L01VBg0f5Oyt+nBbUTLozg9LYqmI/NCUhQlMsvaJAqUbw2EVoLjlI
Wc9ei0Rc/edvJFc5gIfU4hyfyUTKUfPdM2HGdl4uoT/ebgHHYtol1gN7B8Qssbyv
G4CzVrAzV6j3KPyAXLKzjJ+D3zQbK4hNi2Q6AEWD7seNZFOo6W7qlxU1NfVnOrAE
HhPaNU4l/uNAwJchv2qx3kQw0DamDleSdYifnu4KXudZ6XqU9Jkgc9WlEodk3jcI
RBqEVESCvdlbWU26ouVlJIPElAmnSw9CYWjTEG5a/7K1dq9sMB3aq+j9qipDRZuC
RR1CqBI6wt2nZ0ZlZ2DjdcyaWVNoLWHngzUz5+hAOVdv3+zXBObmku5wXsKnMqO8
bkMUILBPihHQmZ4p6TSa8y0TlnaW7dJMz5N3V+yvHYGtkgo50oza+GShLwk/G5lX
Zdu7rngviM8DUmr0M/zniZFb0Lbx+KXqnQdeHxRxRtX+jp0wavT3kSxh2muWTZeq
smN6wGVLdRZlqoveUJtLQqiPgR1TfpLGnlXHQjNsw42Or2LE/CuiXEuyf+eUpFuY
FFbUVRhbsKpwS3db+BJtgvK+IS+BNybvvU8PjxnPWIRf+U0VKTSmHFUs9JhGYMP8
HybcVrvbrdQwb1PGP+ho8IpvJ0/5+hAS5oNknvRsvkOWfbggq2VVir3KyEs+BsDx
aAJCZCGH0W4IH1KDvw4J2kozjSVk1POI0vSwmg4g34MinZAxjARcAQN7UsLdoQTo
is/ZIJ3OF/XYyFvbsTP992guZaJYpH3VW3/W++brkXk21ZFdp2Kpv4JkZgITJY49
VWt1BqW0yybR+DjQO5CeENv/snG8TUX+reVGax5gxVbL+R4dzmEJPl7q5dnI+jWp
TGqWpCgJ0GSVnX+32AKEKnCqWO4+c9R9/ryGVlhxnoPL4tuVTt2mK3vOPt7tqpJO
7oaSMJNFyp7B989RsphqH9f22jh9d8ZeD+8ZoTgPDFS+Leaqz1MkmatHiD3C8/wi
KlC79TX899wdvXPe6puL23mXMUaxnl7VkREj39jZTIi+jNb0HNAr1X+mLIICq1ps
LHPvWLhIaCwPvcNt4rCFTPN2aytyLvhCy0MYozOhzCMA0VufrBU0WGDmYgsgl/bS
4Oe7ocVC/dM9z/lJBe3fq+6ILQbqtba6qBEZFPTa/07Um/8HOGeHbWllXmqMCPEB
8fpznj+eDpQJI8jNURbNeGY/UkKWE6QegLUJdotjD51ksLRTlKuYTkJbvcPZwbaQ
e1l5mgsZ/e71vyq3AQT0irkp0raLZRznxyuLQavgoos2f+6gmn73yrB5SlYQHh//
16Fj4lI1orRtmDelKZe8CtouhM/hty2rZwu4Dea4HNh33dvMFYRp5wqEk09CrGai
xRbUFn/H4fv9P+wyXyV3N7n/TWy5zwoZS0e81sKzTOW9FR457sNuu0VbM+wj3dFG
AhC/wpZungZ6TJUoVdKCeIs9dt7puRpRbAC2eeWw6B/wtLOqhEnXguThsyNgvJRY
sgjRRETUAKzDNZitEO2j0VbTusbkhL48qh8YuTUQKqIu7YhJ2BaTNuntsP2jZLzQ
LxsX49lAqtS362Oh5/HVJHrFOlYn9NoxtEyOCWI/DGGY8R+D/wn8G624BYZBFhpO
clqBjBEO819X8HouzZr0uYiZCFNfyRbIruuQesy1maItp73ZesfJWPLCb5U9hn2q
lStsQl+y0Rg0Khg9PQB6UKojGoPy5ixi7dpUiw/NrmBF2boM7ZZr/c2dU89kB8ug
tMx405yItztMh0wSzuYASFZ+PSAqqKR2o4lumgmrXaJCOybyYFvgIpsKYTp7SbjF
dMoJ56QTB2UgBlGf9X57Bn9HUlA0XgP0TtZbscNZA5tu5PbwwkQ5xv4MN0ZfvdXt
4qNCeufPckLmLNBVMdasAx0KWTnAUcfdl5jd8B04dE1hTEQ3SrrpFmQMlYLFcdRY
GV5XpRVbBf96GjZjhnfWwztRObIrvdwbgre98t86v1dgjaXTLzz5u38QmV8sWDEe
Ea2r7TGFxnqtOLXuQLLhuZI+BrkTmcys2y0ykyNg2Y2ZlYj+YQitJPrmluI347NB
7+CkEkmelaIjPawbiCOf7Ec/pmkyXhkM8OGCSn7S/FgxqT6pVlQxQOyQX7z8NefX
FHCYXzXgsTlwFwgLgjVTpTuVYI9iaNo8JDmUr4nogDiyRU5OpM0UbHzyseK/Pqpx
LnkYleIXt2IzNFTXwuYehYFEJfMK2Uyr3En3SosTqIdOu06BKQCLJ0VJaSttVBgg
41vWR6yn3KD+fstiCPTaLAWVXWDZdaThwWrYDwglHaP+PSz2z4N/JlWes8e0TEv9
geMlyCtC6g+JGFdGOakVqKPOIy8LvV7FaeH8jbPKsddeBRyF76nrL2GnbOvAiZNW
Ix/M3Ig+M/ma1RTEejRizzM7m1WGszQARQyR/Z8bGvGtTTO92bWVNv8xSq9QTyjc
sdktZePFQPGJI9bRE0ysOwXbhu42aigWeBgdvHJhkZieYeFqy5pf6UmbcxiAiF1v
bpsn7v6JfstKxA3IW+/EmRn81hNT3deZBPpLb6z0vLQk5XRjWM4yUVCctF/hxN8e
9S2euKR9UHe9XT9xWxLD411xO6UUHGtADzCNkdTv/BSEYIvbFDDPWAeoSm6htGXK
E0G0sstvCbawHbYkTuKoQgrIf/uiFL4h//wgNrfcnVIRgEie4D7iwJWcn1sgn/Kq
RNrbA33ueElLSsWf1wEkD+qCnG9iggWLl1Kx3CXFIU2zqL/TU5sQ1B6AXd802Z3/
KTkYTvIY692J9NmqAFr4NSU3/jBK91DiUMo/rQAOukHK6PzzMbPNwf3136ga+USy
4sHOaDojKkCUsQXqfEVWEXjq+GoKs4m86jvnFwBbsLy6PW11Yqy6HEXI8xADMu3s
IMzZZBIxaXkt+5P4bt004pEsASgKVmtFZMuxC3yWgNejYC/jMx4mI2xCvpZRjSGO
nA05jZJTkHfjlF7tv6nGdwim++jfoZab1dEzUM+Tzh1SqLeHji/eRLRAfAY+qxxJ
qBmCTwvsBvFq3kv5iklrvQlo7By4WOWyRNIBPdWf+TRIxZ4RChYcRB3VRHaAgZ6/
8OuXkiuSHWXbji5r1b0szu2DIp2gg/Ck0JBm0A1ACACMji9Unkz9ulj6Gly2X87X
ZOET1BrH1K/nWVKk5qHsDzs2O8mz1mXlax4l0DiJsZ1ryaeQvf1/sHn9NcSRZfo8
LyW9APmg+dWKzzhCRxkErcEcwxl6MX8zM1GCR4JiIlN8tYdbud85riClEqqZLVQz
VKqaCfo7HSRDPXfZBTldYo51Ep03ME0KILn0+xDWSwLPcG6yvEDcenW71K9zB0lN
dG3wPNxPQTvbZB1Mog0VdpVgI+22E73XwTc1iK33lWEUmIApMPPjFI34TF5A9kkU
cWzcKx3sJLP5FZftlEI9Ty5rlWTXHzzQvNa3sKKjwxBDJgmFsO4i/zWlQab5IzH3
pa35jMqbhEQed2CSLdzV6lZCuEGn2M0qLr6qSC9rlJVcDuFObdQieMXPQgp9tw5S
QQyp2N4wJRFvRXFbj2L4oB8Ojv0zRy5vM2Oc9mh1ykCiiQEIGS1Zjf4btH22RGAg
JE/9JEKkgXaNHVFbhkfO30NvpSGV490gBRlV4qKvCZMHEXP6kLQRwil+zcZA7uMz
xDvjUmTPNCKeOz84pAg9PRRXIxphpFMFZKZTJwo6BgqVCVkmrhT8bujr8Kgg20wt
LNTuPeAiQhKNHuyAoK5PewQRLSBZPUi/8UxXM8ehwve+o20P3o5j7a1ukLbGQKLh
XM/e7NXd6LblkaukrO04WAQ5jh/NSTJ70mzNcBC8zi2AxWES+64mIPdkakosTNeL
j8BeuB4ZldxsJ/Il2dO1v+Onvr2qNonDX2amUirPMyD9nyS9UeNo47PjBzuWiCUR
xcE5CZnMylXGJgplDlZOzjnmLyzVqrDe4RhRJhYfp+BeoDPqrAxRZQPAfpRrIKT+
B5SCjCi30k2ARSRlbAyu/m3lYIXwir5uzYRrj+Xpu70UwXOitIZZhQYFFbjugnMX
MJXI0IyWxBBVEjHha2qn4qFgF9raL+vTHHFQDA1DlbwvTm/kD5oUlH9WPuELt5su
6NwXr2R3hvlsseTBxwejIznb+w1wOf9Wcw5lGuaCNAtz7vP4RcM7C5rtwKWNhLgr
FscOt8p++tUmrnGpbjXAndSzEzakUOfrqipsxIOo6BzoGTcC1KMZM5iVPKrVzvwA
QWE04W7ff1xu9GjGp/CpfQFbWtCPDVIlUiLlHjGiQLzkCzw8Hzfe4PImlPZgNoRK
fXpOD19ukGPVV7EUCoO0LvcNzNcedNCnRIhpnvHGaSWzPFtyBtUe/6dGtHo3IMI+
iA4mN7EubcxrOkZJ8LteQuBYOaoexOYwuX7MnWKBXd4B8fYIRdRyuPB4+gmN5sqc
ZEwRbSzLBz7K/6wmnPMhpYlvH83YW58b2XdaqB5cGO4sK4XwG1zGzohq6IRPy6xJ
jBqklZua8/Rj2eFbng4kr22SpRXqiPPgdHrGCQg1ncmNrregL3jga5+Z8eoCJYC5
W+Qg4+5F8mFhuf3Tf0LRB5V48nWTbyBcSMzk65on2uWM3wR20A3xY4FyKMBv3lwf
SE8YtcHgB9fow0o7i8Ctu4yU9nExpEIzo+s5oadeZNsS4DpdYFQ5Q6NUBy4/x5PO
Lknd1W0UAlhEuOO8D3bNBKL1gLNH2kLO2mrtfgJo9Dmbq+TFnlN53jePLZ164VzK
0FvhtWUFR0nqycGyRoCO8xg2KJOOQdSvPAyJ/8inpQfrotsK5xUxED9bn8MrG07b
x2C/x7OcXf1R++JOe3DjVVlMbkZoBNaNfIj1HMNUOMsoR+F/9EiFb9WGNHpW9ahL
giQmPsvxS3m9T5uQsuNpGu5U9ZjamD1rdn0sCPbdDJHHQ15rfPVc/pnYI4pIKfmr
Kqtn2ZD/TheNrGpHibgXSf0J4mgJ6YiT/vxGoLODHV3r0gtOMdwdDaUGBaSUX8pX
kg5dmYJ/Ut4BA/ufZddAHY/puHwaoMca/ibI/v58WsmuEmHN34vGBCDNMqodvfkK
fKjKAoHypyKgdes0yfP5pZ0diGd8W4UHJIefcujLJnlDyFIsi3MziEd03J+A9S4I
tgWaG6atzXq5DsyjvNeYfkTewn15ZWjP6kNaUjThIJ0KR7kt1zYQPcASLqeqRt6p
6t6SsIJ4iBl1KDzh9D9WAm1CBc08XJHJSgufS/qr+MtBkREvMNkSOI6WfR9wdCD5
PF3gqe7tYQ5P7d0H09DIDi6lx21y0Gcy1fUD0bWD72w1sLGIjxuNa+w1Qq8xQWqm
Rmmqqp8UNOwEK4gP5zgvgMRtH3McBkP6CNIj7GImN8S/6NHMGJJICTqzuPa261bc
ULHwre4Np4t/E+yMU0ahYF5oGehGG0xtQSt7ISwnVxIOrabi8S8unQxovHFhdoLE
DOhyGT6Hjsl+RukCKX+ZmXKs3m+RS+bZbkuRVC6QcsboeEpKbKrfUERy+ZAS36C9
d4BM7SGvxFfG8gjGSOk28EDuhn3Y9jlBOIpWs4YRGxi5/sFfyyrBId5u2hxc3vSa
Mf/lBD5BBY7JLefF5aa20yhMqYoU6OHLDUC6Ef2Z9Cs4/MUrcUQHfKIOnK70FgwI
iT7YXsyltN4wgOfOInB1xb/v4mRySDyzNHsQKZI2d21pHIPcbZL2vWpwvwTSnIqj
DlDQfZnAYBaxRPKu4ChAAsRyv/Yox1X3eoGEeTWIHGokD+6+c3xSTcmIJ4MOKopu
mtit6YsHScBRXpmmB0+sRb8MSkd5Sem3dqBOmulcx3roEvFslIjC5dG+UM1a49Ci
fRxLtkTKzN3CVgKdEja2MRSJfBFRZc3JIFSvCEQOLp85UTZNkK1ZRkRKgj91rB7L
SQzjCOQ4JTvJQxWtYcvmeECchC7negAJdtxv3qycF7w9P+L0MxYTHF8v+yYreRIE
7WQdsGYAQjycswbmUcWw2oPtQH3jDWzXzoF2S0kNcrNeWWZRCWj29Q4si6rsf21G
hYSKNwNf1QqRUN2XQyZHEBTY8QdL3Gr2a4KO3qR+1P/NTgFLjBqMbn7N4bKMxwYD
kL1hUh+7bnL7yedQNjntW5n2UHTGXoDsQvD9HpVS1jx1r1ybwWuaS8AKBKtdF5sK
6JkotFfxMwpEOdJjNpONSHadBtbslPsyu70PhOyd1bKrR4Cn3n/8/keSzugrCg6J
fWJK+0h4F5hbN2zjpHhNFrqZDTLEzZf0DP8ng7sSquOqHsfhwbS7QVOZqSnZd6y6
Hel8LAPg6Yt1CYg3p+Kh0uUTrMW2sHFq+aD3BlzyqE3IamiQF33vQ8nqAUDPp1mt
UEw6U9IKGcqXFdl8PG829m69WssSxow4V1btmQjAb1y1cZxioAYqa2K2zLd7geLP
/t5/i/rrxJOhixuhUfsW2HRS7R+W+Qy2Ap4XsFWf8hdk+e9So0q+urskew33F0/s
Hvu+xrifeTsBYkFXiuXJCpedSpx2H5RizhPlxwsfEBbGcgOMDUeuYu9HG1h/gAcE
HXNU0L4WAwJ7i2U5U70NST58Wi1naZsUM87dPpjNgy8n6M7Q5sDZLuMTcXWcwUd+
YFE7BaXx0mYqRhD+yx8zuD2Xwb0Iz2JBS1/RjVVRrJGC8HewoMY3DZsk1MCIGw/2
hfSjEc4kbhGKmGTkRl+dhiOcuNM5EYM7rsllk2s/fnVAD+MHXzUMkfSqWa4xHcan
Suf2R1NwNe/gCgg8rdDOxp7a96aakXH1MbLNUDGxoBuwqjJk3G2toUhCJJSVl/rI
dSjw5OQ+AAcFr0w13fzerNHhvIcAo7OUdhXpOQEAzO0HuCTsgyJKcm8MBa/12W6H
x9OgSQhinlfatyA9UTVQ5qabVOLSYdGRw/c/qK6Bmc0d0yWs1WmpFPZHSxFKI2+H
EmPz9tsyPgihzOXvXBob0hp7sISsJW6+R3eOGb7q98TSwqx35jKhIOGMGFqzszQS
jCmNS/Thq7ml5RsJm4YnRIV4TQQc74GYfmYhxsC4F9q3Hf2zh1jHkYOLVtfHMOps
o+/RLJPqtQyPt3QeGv43j+9xAwrzmJQ5AqJmVkEQIm8jnvDGQUuAZCTjgb/8njgW
w1JEb43/A7QuBvNrL7RzeKR48OXdiU+sp/ha1JV7+1MpgRnvWVEQSgLfTdpPPtov
qkGGucvzm8INaVCSMfS5IpDrUxjzWjh0DJivXHQF/+0eZ52MXWF0nLVDko8GX7WZ
BTXQM5swC/0puAYieZCb4tMgrAvNmLRQlUiwr3vppFxT6YLO1nPzrFwlv4ua5w+B
g9nxpyOTJ0/iiscfadXWc8ECM+9xw/7QaW2xO4hrGpTK/gYhKml1RejdCyqkmuwv
3Cfe/YdtHNkGFDauCRiXbmIfZXGmtYzhsKgVfIfbsBbVoWRDsqnJs0Y/LsDzphPB
m0sN4kb0BrmkwQT70Fmu0V+qGYVBFeUlijKztm3HUXOGshIEsXr3LlgZr2NMVP5u
OJjJ7mImet4xHJIuYmpStKvqYDbXBFPU64TzzmXnhtBkVwKty18u08chc8q94AdS
aTIMR2Lzeh6hlUCBuxNlh9EvOMsab3uw3ZyGbGWdgXaYDAl4IW3REz9Lg555mCqp
IiTSJlU4gScCwsQytzpUUf4v1P2dK2ThgsXb8Y9YPQ7evxkKJ9MidC27HRyUIdVJ
NCn3IFUpIO1hh2TljYLwwEwX8M3l/2vRzONgf4oCk3eIZFgSiGNk+eL6ZxkshV+i
Gk9HIPKKE9FvC5AquH0axkPiEDVFGojhJWa/n4YQGIQvMv+4FEocTnMSE/b0IX+Z
f8v8rNCB47zwvh17pXQ37dF8wo50QyFfZC7mURo2KyUxDt1zD/cOXo8TJopfKWb5
XRzCSESDFu39TrDQQEAIoqbpDieU7788VfN8Ji87BzM1/QfX3eO2cAfi/4s1Fl7X
1PxFNoqJSe+lNvM8wjpfWUX0L9tfu2XJAq18ULwNrBTAKc/dKDQuhDMH7LPp5o5K
njdJy2RdDek2opcICyu+br3oyxERrZx0b8c9NAfY2vmsCTULMh/QncNxcuVxMccu
/81POBBOJWOMAf+L7i1reCNj38ffD5gj7uazgav+SLIpHRCNH6/Sv3ptYTRxnykY
QOCEKIXenzxoJIFjgaSzW6XWAT1TNRr65/i0rh3lp4vlVHtzgaGNNb0iwz6+r5+B
eGA536oGKu8SZwOsJLYlt9slUS+pNlncx/1M1C6XBM1du1g2olgsTU4siId2zCAM
pP/9wxgSzpIpjzji6wStArCpx0aMBFSIZRL3ifSABVdYsu4Hl/qLR6AAW7sgSrkG
8t4nHXpw2JJsPvgGuRjWgScu1T/8wE0TOEhRHmQ9bGYQUAQa2CKYIfde9OLFapUr
QCfqxBHk7Vc7O9YCFHOf8PDmbqteHa0lR8wH7Qic4k8cEW64O0hNeqnpbsVptHJc
uf93a9u6wFOIoIaIXi+dDGCTDgminwS4kpvPD184gimiX6UIUBuPCA5P58OMlr2Z
SqgY+gEopvzB22h908kpn+DUP85A1lqIK06g3rOO9nfox/0YOORCVcpbJICaNivi
CPzXQvKIUXjmOawceetmZbrLRsTiBoMwoXpNsYQkFLXPdJtfwvHtttnuBr+yOe/g
YOrs1Jv+pF4LF6xFdFC83fuLbzl0KHrfFm+mbsdskql9zxLmpbfm0sv/CYNf284R
zoS8rHpGNM5SfXvERv4kDAkw9Rs7R2tUb/1ibqGvBdo5uxNCaywYg++YhxmLXNCd
dRgKLDd/zIaVvIzELgiHYKl33sbQBDOIoyYBx8OvC8Umo1k4UaN9sMVdZfpLV2aX
1PSTRefoS25iWmjjEbIPXUXwVosvUVegOAK8NZjjVv7hBQFNSaLOzyy6dsPBnGQD
1z9CDBRg82/T40CWHxPGD4kcIQ5evNxijfNeskJDXmGtUNntvXF8rDsgtDaR+h+g
DMAGw3PWTNKgr2EqKcgVtjXVzFyetoht1AxQXUk6vkSnDcAi9nShPcEAaWUJpGYb
PFN2sAV3WPmJcnIUy7jIuJbJeAtYblLFUlz0fWxJ41UyTzfadjRbomRehedka/A4
WrGB9O+l74PqqqnyocODQwjxdOlJPU68zsK0eJaaCBobyIpLCEGHLLzMCGQ3867R
aozPBH84rsnknnm5ikDkz+UON/pnvjxZZ5cTZO+XuY4fQnin1TTLlVGEr6244o9U
ksfehzWZXYdE/vwRbgr2JK0PZ9iOElOR45eTzWaSnZV3QSBnJr1ukZODUZVwJwPG
n233PoM26jiZ64ppD9gKlFibOOssicr10QGJb0tqloqXI09I9GyEoq2QHd5oM/db
BxfGDA5B2BWWBW7cVaBPi/euD/mzunZbQWLOYMVh6Ir9S1oH/Jvpg+yUUg5sh20U
bivAWyxCippAP6lSGjSQF2oPXNDvdazXUAchYHhpt8uikCTAPz/OqHMrQ4R+x2q2
bElgy1ORNS7Eb/VygJt/Gr/nmDRgLKJ+vzaUkL8s/b/9CXwH9hI2gIuyoX3CW8Hh
vMeVVf9dqWvfwIZBEda5KzaK2J8vOrYaoatI/k6v2SofyVX4GyS3/9dId2azHrfW
l9yy08J6vzlnYGW6NidQvfAI3MBvSLeaUV95WaMsbZGktsbIr41VCOugjL7r2esy
j4YNl7350Wl9yn8JgwJokE3OuHZOgCiKjJTWvwd05PvaRdY0y6wIt1p+84FDMiij
1Eq/xm8Xg3lSU2cJGFtvWshpwMM9PNPHs/xs/8W5sw1gffRGYBMU6JnlOiPnPCPc
kr+0JSwN4Udp2qtkg05YY9rh1sGPptmv3hVNLREy34OXSwf7nHS3N0NVCluP2N6s
t6dalHPY7LA9X2bKXePFLZkHpFrKaKFGfSTL/sxlKp0hWK5yecJK+oRJELCzcRy4
AGv73EHQ8mMZKie65Eq+6rfkBvkFeJYK89Gyws5k085YQw+nc/sJjIcPjrSRfRyy
O77YPe4Sy6UeeI++XmOiMOjO4Q5o0zSo+N9NzXSAyNsoTOjCIu6p3bOYf6T5dm7r
ATZSbLBaILz7cQffBBQSZPpCo0CiO+cnbCNDsmn59de186R+ZuoFZMoVdlLo4/sR
nInILspaV8RDmV7s9LEvcMcuAFhy7Rh7T+0Icem9hn2we5JzrbqUpyM3ZFbAZQ0s
9gr6YBlPrHf5MUSs9itqKBxZqTYnFveboL0vM76nkfCRjukZxqh2fSX2rdrYqTxn
tGtYEmu+srlyLusjq/dkMz+x37hHmNph2WW98qFSWevkdX1ZDENy4JchMI0ZHV2E
mT5EBQNAERtlxfYf8uzItaOjZ7EurgxDUTDvX9ApYIao5bkRGr50KMb/rO4XQ6Hx
Lq5Y02AfxtZyc9VbHDwEhg6lZEcdmc48aXxQpYaDlYUUO8AefGGkJvYDBzGWxhPv
0x1AkujivxohjgFKEbTQDiZT19XpGiaRbXEnFuy+STBoc2u03WMravA3bZGk9BJB
YHXXeRros7Hqe/po3Z95+X2eBhf63brelPhlsWSN5vyuTsVvEuzUWjSAh3UvyCjx
cvPlIyd183TDmVLPKTDyJOMm74NyZZGWsUEcWxmm8sM7YEIh/2HaGpy6Bs7F12MF
+0Tf3a+VI6XXLQe/I6UxPoEheTQiD0GgsW37sd+0HnexPNIHEdRH45b7PsPgXvoj
piilTMUm69q/6TAgvp4V4oad3cEXRow5U8cMltOby6BYjJxbSRr7lhAn2tSunGcx
eUruXx1Ifb5H4FOGz9kJCXAJTx2omCbAhaNzFHKSTi2oRC5L0+9F6wznSJafYwtD
J0DgI/7okxdzr7QI1sy4UwsIp/L2YsP+ItksjRSIa312lrAaopngxqgjpYCnMtdP
GKZNzJzhQnCCqaCe/o0q4dHOZxPpAmtjhs3YtZ+Iqz+I7SPP8yStJaT3qCUpRS2C
9doocMR5HuWcSMt61itYqFlYI/0tnj1C0NIBQ8FPmWlwOENyBuOvsBJwJWlME0+7
DRViIM6WfUjypavJqVzti865dKoQC3tdNYJWS7C68z72UaSZPWyu0NApt1uCQNSW
K35qp+Lwe2ZMXKjex27Zocxfng3Iz8baC0y4wSPUAEbj/SW2+nrk0GrA2cVE/DYD
+c6bLM1cvsGoyGAcGz+w4bY/Kk7L76ktsLMjLncy/wtqLeDevylJ8GKGJlbGSczG
fZ1Bm33Akrh9JTSdyamkK4QDG7MzgQH8+mjXPEqGKUiv7LTyTH+IC58hfWm9uK8t
0Z0KpOx9yMIv8vGDiUfA7Y2ZegdabRYUtJY1oHraL+NeG+a7LDH6vB8kXlTKCwk7
VivA7+6VS4YvaO+GTRLe9EpLJAhJtUrB5fA+FpsJW7vaPSgcSm5RyQAjEphzK1uH
HXQn2PSU/mOnqEicf+jMDeIIGpkVPluJzUl+Z3xY+RJh5dsSR/7CKZQyYLRVxQRr
yOig8ifP3BZl99Aa+sbkmkqN+GSFPwHtBCl/W3ygA2iSQ5e4OCbHGPw8aTAeWYzU
YXmv5eDcYQrgRY9u5tjQS2UinBpM3Xrn3VQyEr51lF/55H2QZriNwF39HctlPT43
ebizX8hUzjeLSAIhsO2b2PrJPOw4K3xSmg9N3wvSZpMSZaoDuIge0An5KIEfUTTq
443p3Mmvod+T4gmphC2vxSRmZsyqyAaRu+cSr3fDGvOKQWU+6bPtp876V9JbejcB
aEw3OP1QA94NOavsMH/oTo4opWBQjM73inNWS/BWLsgx5PYKfFL1cDLZLXLU9G9U
a9tO7e2rpSlicy9DOBcp1A5GayGKizwxU70BhwjR0UYOIbNYn7g6j+1fxAwweaAU
u3V2hpBvypRMZZOiI2lczBCMqS3XN3TBbDGRFau1QuCx8P4SwAKySnBbCoTxgW85
/m2KsDbtb7TL1lypPF4txfSNLVfKdiT3TiwPNQ4AFS4HIZ6QPBTJ1N65uVr+Go23
X9kZmHoyemt/IeC2ZDM62uVTzzn3490H5+nN28oR0lQKZcr2AakLwSU9q/05Jr9g
WvW39iukMZtGuZ6jiVfxmaQchkzBPEMCGlMa9Z6uathgFez9ZmsbhdERVTDsrkax
jgEMMjTWT1BdU12hR8fpvtwXeJzkmxWoZnVRIxFCNI1ekDd9XVnS+DpIRfSxD0B3
P/qgwZEl167kIKPieCM7ZM0OmooWiNXM8a0DQLWSlpoUQ10+K1XwCL+I3Xo5wC+d
hPL2IOSvtPVeo0zMxx30GkYIrSPafbvK2gk5yrCBiRVaAVz8alStFGdB3Jp9m75H
o/S6nufmSRCKvFUFLAcmR/Oxc7qORuShULv4GwFhz8KK2xVm/BYZFw8MuuC32IOP
aV1J9zXa54S4teEuT7iHY+3QGg4mZ5FP8n2T7PuG/HfRonD/g15InbCci46n1TnK
pMxI9qMxcq/cTaI3RRY07tJLakT1ha+974CYLonJ8gWEpC/z+BnOK9bC7qc7oo6y
tWKUANIQ5BKG77t6O0m3W0PopTpwPFeZcyenwFKxaTnpSeE22LpmLbGz12c+QVKF
4KaflhZ8EnnllBR9Lh1kS75d9hcxLc8Ub48EyxZ5/+PlmAmabB1pOGrgR7MhOvFi
e/giGP62U2ih1WXo4WVSklNFHWBKluvYrX4ibh7SvoakLPnOqHixU+cHo221WrBj
bb4m15lX9wK1I2m2Olb/d1MxEMF6GTfJAxUiMS2bBJKUK2BecU0rxgbGB2itw39D
jSv6aczBQeq87x6CbEmLIywqANWEvoox2/tAYYt1T9lsNTakashmfa3kp52u5B5H
U2VcKiyxUf7Y/bPcQ9lDjBiLY/tGIfJJqJJSiBJgYhxUYIYgSPhjsbv+ZGFEJryL
fp1yz73cJFPc4AyGKzQWZayGMrqL7KBqVdjqufsO/+TZSQ/orcWa1F+2Hj+I2YYi
J4/4r3W8myT/3+DZt/x8Esfu0vAYuX9wsxckDuiBfmEyh8EOAAsAeN/HI1foDNA6
CXYeOD/c77mahC5NyMPIO4Vmf39lJ8esCKB/JnHIRXGPNqkUwuvR4fXZXT+Nvk6t
CImckZTSrqu3oBSAbTvEkE2BrwCm4ab1/nYLisH5Uk3fssBTdEDsfd6De0/7T/EL
5XXq/eDwWx/yhIxZpVs5P18LyscBelYm2tjKOcOe5jCTvFP6VRpmtEWkISY/KXex
JzUQO/o/9BFQU8drA+e6O/jFKxrqqCuvN+iQhTiSQKUZfGTerXvuZb7wCBH5KGCf
9PZnn8uAZe5M/4c0qc9C+92mLGTpS/gaLfVIeMLjfeMuZpPh9insSdoDks5EUG5Y
p1WZAnCbaKr01wTPMjFHQD7nNaU5nNYP9enF4wAtlOJM690Xe0dMBTJ4mmTDtjiP
TCGlXT1uYhdzI+3JHOmaPPTBapGA/LOeuf6jPucsiqOAZBHK1wd/ja+MBz0cDZYm
5FFWeHycuMqeHNfE7rSDPkcp8lJxfh4jF14hT09kKuH588EDnuLUxtukOtyKXyto
cKGV0zUpEc9DD0qXoUQ/KAw+tRXbred1mu1RitDRsQmSxKL11jAY7WnFh2OFOaK5
1ZChev0NQzfUDsR1vRE9RvEsY7vykOERG352zxQ2K48Dee4vQBb+BrMVFE6NA8Ce
MKFPc47vwcYPV3w7X7N6SjUdGm/BX5MjX6JNirh7NSrByElM7BAd6My1Dr2qh6ya
v5H9XmAGgZLCgWXN3/pnX9GMxDSMtks9Ot0/ySGu0dw1j2ToZxvW1Vj9ZDgM/T8n
dc0SffIEU2h9oDGhUojtM8KmFPet3eUfqYPw9+yzEVucqi+LQ93sQVAjTso6HuCe
Awm4fyxb9ySQnbSjWS0rZZthAwdIzwZrVRiQ9M9fPW/Ao8K2ro6dP2WNBfuaxZj9
KTooaG7gbiJ7i+1jPx8SY66BpTeBd9UBBxa2bbHpEQ8y1/2VFhmBQQ5m+/WPs02d
rcr5KHiSUiLkcPk4VEILwl8qfKmtrycmfUwKkCItXJh4MlUMEvvUHvfNh/9a1pdG
l9F4VPrjFEu96SjFbPw/ilM5L64RiIUJFtbEjuJqMuZ0j6GCFo+aaXET9/Pabkpu
SlmfypjPDOVmBsPQOs7c22YOfxp6xuGZzCSC3e8j9/n1lScMwqkhlLOkkiKHf93N
g4PzK+7E3GbFw4sPdtM2riZ8DwPvHWQwxGQV13VyD6jQ3osSTgxOCPGEhRux2YVw
banljdtWk4mEh3ZC/MS2hjp3QAbIANYfbdwMqHa3CEnCLHnS7cSVVjwTB5T6VPiv
1hjgD36+Eb1GjjtuJeO8fKnID/ec4Ddmf9KcAfMvqp5mjbaBjh4JWsqaTvxJIk1Y
FJFwOpttq6WWS8qtWAXvUx/X3YV9UiOL+pAAsaICrRWqNUMfhYl5SkZSzem5Xuum
X7G3wA1Ymn/t7lJTPaJeBCDI6F/y7Tnot6/xfkEU7IKb/zXAlSZ3B65xx4qQZUZJ
J3P4gKdytajajyYtjuloj0Es+CqlEzM7QyshLF/7sOPwQ2cD3Uy4NmCWucAKs8YY
Fy1c3QD3qc5jxClM5jqIKaSePbTUhWChMq+CfokjWDMwow9/HbLanE2gRJ8WivXI
/j8O5IT8gXm9qZA9dMYNUPk+nveBohrHgeij8/8qxyI/k3B4Jxro1sz5gED2pwld
SQUskt0BzQGqQ7OtS7NCBFe5z7tMVQFG1UceV3uEIb7dhWdyNWdyEv26+lJHsDMC
moXaYpYACa3MaxGD93vbzMlHO3/nCUJq/mi3fRHnZbvuV7mRYUtIlYvYtJP88zBH
KXi+WnSnl1XHwcgZUHnwjrrUOji0QL7QCu6nP7eGPImO61FMlIivBJgf7HWb8EOO
HN8UBPUwRcrjmDG8wqj3FSunfjRqIU3UgDIVKv7hYoxWf9kG49Pe6JlDAcqZhBwC
0iRxBF7AdnbbLnfld+aK/O96EBzs6lgaKTM/3fS6ioBrwZ81r2g5Mz9qry1nnvZI
aCtEoGGu21RkRGgwhlpFKEtIuHhcWKBlmbJf0Dd5+3jS3qxnNndSO9qmbC4dj9ZI
+UvwH7tPywvqCi0ynRBOwd/Ur+LTb6UDLrp0hL3cLvHdJnAd3BPVs/6mb1VzYAOG
r94hsKvhcNY0MvpDAnuDJzAsZhmXERwvl7ADjaF9dd9Em/9p7pnHib4XWAmLD9ld
58gE/Gk08jHo/JZReajvhhYJ5xuWn4TwaZNG+hs6VGma9G56GLcLHfXxVtYKJQWd
YczDs38CB8tvYB3abNkjlBjgwBAJcEQ0vfZo9gmznb0NhP73gurs+ux8baYrcWQD
m/IBLdR8E8a4VEQeaiC8TzC+Guo3vDv7HQqJK9DaJ05D8nNLikiLY3H/5Y/4FwYa
W0WVImlRA+vfqXXTcK56GGV8kxpldcE/NlBiHNTSy6TD4jSM4F3bRctcJwoDLbq7
44xJ+VB3cK/Z0rXSo119liR1nPdH+hg3MJHPKXymGCSQid5+R9HthtWNxnebpeBx
5CphmLiovxm8wHwNpv7tEUNxpft/Lg+YCaSIePe/Qn8zKFLMa+d76LET+B00okmC
YhshsKjgv6YktoFt7TekMfyXnN5RMK8uLcc8qxIALjjRSk0WZOjHDXMiWVAZdUo+
ka2I5mlVy8rTjZR9hc+2Xlx34Q/uorQxOoPSwnhHtxTk+3Txzp1Z2tJw/uV98TBP
BroNDJHveqOMsdMps30TrY7SxtbgvQCuugNzDGB6/d7fwU9eMxVSpiGTHVxH6Aue
fBR5Cr6BCRgrI6Hmtv1amBR7x+1S4Wiq2xJaiAGJpLRGG5vxxwnYMCIfkOwZNiqT
qO0zbICHdhXR+tf5PNOSyW7Tx0cUUSDJ7CEG5lGy9Ko4GvPYD4G14MKhXEYxpo/x
vooE4sOeGYS3bU5MKsvF7hxoH859jUa1G1aMKMYFAfQAa+7AvTlajRjheq7cAdFS
U6ZE4OXR0lmUzI6+kjWmNsW6hWQOi96u2SwA2/+/w24TAncUtBG22AJZ8/99ww5L
qPepqnmr0EP0JIGxWU1Omy1Q8Xelmc8fUPNb50QemC0GP8mDqygBRYLW7CEO9Wd6
wzXF3nv+TlDZi0hYDapPIw9tw73D4Zzc0lvKy7mWDbDX082rUS3h33FpJgoMeM3O
hMWPQ3SQBvahYMpB6ARDSCoW3W/AV6ZRUziaDmpcIISB7glues4gjXccHfFCVTpw
YC1LizO61YkTyI44malVup2BOnWgcLVWaIjRMBnItX9KmjmgfeY5g/4B/FuilRq6
STvl20GIKa8wCsaTSZF6fN+xWGRcWueAODGwydv5/deOcu6H4PkAg2amVvj3qeHs
D24LO6KEnVCu07NGMMoFvoKuE1R8eBuSoZmyfeZVQAcppV3XX0vUSg65KawVJ7Qh
1E2xWt0aJdIendAAlyQ2vV1EqNI3aIbzM0g5AfHOqRXVEM978C9cOppiqNVNNxpo
/FMQgr9XnLF1zD8L8yoZtM9EWK+cplJBKMAWUHpzdCHB11MuHGjVlCTOsrGVOVe3
nadYN9GVLoWrqlbeeivj5JTh27Oan2TdHIar3AUIzc0Q0CgDNpn6NVT5DRQ7+Xi+
TYRWKK1pkYMey+zTu0S2MK2C1XZ26hkuWBkg5GFhgBojpNwU/B5VlqJD/p5OJQtn
tVQA8z/eaaIkFD33yGw0yOAqfixJM1wzdVKOtx7ffyUa4j0ntUoIXl04M+sYgr5N
6S0M0pSLxBlKZ1f3TKJPho8VZglo0i+kOO/BrxW1WcFemfcII7wdTTnwhioWaa/a
8cNA3489iwONF3eaakudlSJn2AgdSzsTCUcpkhYFMVA8T2qYcSPz3FvsJXPyxIk4
ldZYJLMSgvRNEtfJmtYV9wTNERgd52JZDtLf6LdXUKrCAJCg+wVbjtxkw5lldK6A
lVDvH4xJhA5RIQHZSD72MhnK1CjYnFDxHB47xIuUmAY5m788RNAqD2DmbG8UV4z1
ROsOwX7qFJk8lb5cZxm85IobliijoQ9L4+68yzmoiaqrmrCUynvrG6M4Odj9+Otq
WG+pGbayeF1mCVOHZlrsZRk/lTtdPUXfj+XSMG8pNd5zJnlpBmhcMIvLLpygUL+0
6c6ACsHyCAr3Ga/XaVDyrUMrU5YwKDJVj8c7SL87ImFNkbzZcj2gm4fF1s83DDF8
/lsEOhaKeLTPEVfXycWgiWqzY1FM52aDNOz9ysT39oAapA/H7QSb2WCRa3QBxwjn
E9PjzQuwlfzH8+4LhgzT+sRaZn4ToJBIKjHa35NzOUU597uun/5iSj2KUwKeLdWy
By7uOY46eWQoTKaJK4eE+045hUQbdhqG9hwU0EKYCaPDr+0THYSvpkt9xD0h5OCx
IjzFdQRvhzSdb6olo+Wj13URoTfxJnKWPnySbwn0ufp/+t1NSm54r3PzHVv6GIR8
UuF9J0Q0lpfDRE7Km76Vgoq/BH0W03koUyqVRKpmLVPAxnzB/2MWdgMx7GrMr13K
Y8MpSoJMcW/LQ8LV7U/qdJEWon5bVzisTZdQJnOEXJ8hqSOhqHieEw5pIzZ0/nyH
qbfx8T6lxONyPM9GRukX/EBg+PgfLgUv+JSw+2tKCakjAffZ+RS/oJKuZQ9O5JoJ
952dhArzvZMjpHj7f+NfnPkhUn7ZOxULlZkzSDgOxy6lN1GotbuSKkXFR1nmoOvE
f1/5fadjBTp+gElkYNeoA6h1h0ZHJhP6ETESlJ3iL9V7XG47u8TGngdeUBKrxUfT
bzIBhBlGpdAN4ugcObaVikOWXIZStWcieDnzWiA0a27I7n5w5QrwZZfgZKGRIzPw
jeodbEF28I5sqdu2YwMSotmOVidEmTKjnoEaXL+zV63tPBYinoW+EQi1XpB1vpmv
riA5209Cv3EN3We0kxxc1d2z7LUDnyJiQl03znsy3ptdFZ5mP06QhMSNC/GvIy0V
lnp4ZODToTmRmyPEaHR/xnmrEKedzOpNjW9tRcr4WVggYp5YzOuKE/5d6PHcHXMe
i78k2g1iSFvzegCwDL5SC+7/AALBt92j/R7qWr7XdV7udzM5fk5BNh5f9pFpOvnc
bZTfCdXaUijwVmdaTfvs1BK67HsxnTlOZ7LV2LUW8oXPWwDwcZx82i0F52/SJP5l
vDzc2Czh3XIgxjxlL3B0OzOs0b1lpMJyncVTHQR7QJvR3PwDFsAIJjfZ5iwXqAuT
XBQoU7BmLXVCM1O1bPit7GtO5uWKWe+IqihgIxaxaTsPeYNAKLwv8r8HkK74VLvi
yqEzKQgEO8vYx0Z6nCo4YGaM5athevngUwjBpCGCrKk82qYSpsgE7plATzEbD/ph
5TvjOPecxV2BQELiKkvGlG7E9GaA2IiT/ug2WXF2t6jO73H538DqGKM0M9eJpQQC
v3OUJAgnluJnFHop9odR8ZsleJaW4uUjGq135bNhfamgko2XxiEZmHRztu7x1X+B
j+r48RD661OpC+1vFrJvrtuxn5OxpreB0MzMvZghY06wlXq2ZoZWNOy5qecBK4NR
mkC/EFHzxxqO1kFvjCyhSuoU9SnJ6hfPdwC1FClFKMBcgTj5EdPSCyYWGgJUdBs+
tasgO73GRZoXunGWG8NaR7UclmLHeg0xZVxgJq2kc1RI9YMDP33K5B5iiBgqHXIY
1HhTplmr6FlWkxMSH7IxsDzHDW8BJ3getCiYy7RKGQQ9B5HjwH3hkhHczsp+B5Yo
YnqBpDBSqGFz+37S4NZFvxKbw6R1qn7Lclo304k2SWYVprEccXL8+gqJsDFV4EHi
QD/FxFqv7elpFIRP0UW4HsP+nFNSAfygoKGHB+vk9xvbg4wqnPSpd813zxw13Y5s
2nMHrU1wcefnWo1LEdx/aTooQeeV5u1Q5pElf4NHCK4vuDg+gHZdluOoKTDsexT/
C0uXu78FI0bzIaQ31stXq+vWVc5nNO6BLyqOLKmbinH/fZgQIM5QZBrRhTuXZ/WR
enJfFj2uaQ/inW7jef/kIIu+R1tVFKazXa+inaRRsapQTvUaqjXukLTDaPZs4Vlt
IEH82IbbNGMiMLN3N/vtOmVdg4wEsBrcqs2kFzLTUdnSrauIyu92X579IVdoAVfY
/ZqsCXNm9CV7EtTrflAii9K5LnpFSUPQuZA18CA6AsuZm5NzDFVVbBBwMtquGrSt
uL/dPaf97WXPwjeR+1FoaxDOS3PF6e8IcA9jIxw67PcgHvopk4zYgccHQt63Bwil
P536Z1FHq673JxxOs8UfbCfdMk86FAhCVpMMxvFVJ1S8EwcfbW2qYS8ejjpj7cW6
Rzg/eyxeb3aCYWimaKNsZrlthzjMERVt+Y0OI/eO3sq9OLdGkpEuHrjJ5F+xfvYs
bpiFkQTYdgQg0u4apJIN9/pMLDt0F0aUTkvmEdt2Y5udFAXo2/2B4E4yd0bAGOuz
Spj+MR8f96gNVLw3m7TB3H6VRQ7jY+1WdAGc1eyg4DPW21rHT37YKzPmrXZvHtlG
vIWii2i5xcX5CpL4xhIT7WqACAbWz9/F4aeMdCx7h3CwVw035F9BMJiNQJo1GIo0
yQSSLHQfT/7QjfEFxbP2NNWVlfX2bf0TZFWG4dC1Z0ukXlMvf3f2fc9erUjv1xov
LrPBcpIe3ey/azegWptqQbAzTYHdq74CbuC38lqBhp5XHjaVGBVugJKXcyXXzSIl
HePDteEEXdDAHpNpl8jdWsvJGXgNYxYl2dzqcpQIkimlwhOQIw4TFVpPsj7xQ7Gz
CDEadhmbBRMKJazB5suVRDQQr3hQ59ofplQial7kxeJ6YYGcc1j5AI1+u8jATBKr
Q3s//g6XSW1Zm+x1q+7GtfAFZBAFYRp8MODMwk2A4lJ6jj+HF+DTBkux9stXT9lo
GpYGAlWE24s7I4hLgvc/rD4in7jAWGSgNlPdt0Unel/aGxY6CshRhHcOEIqj8LW7
+VcWqpXWT1hEHY1IpbsJW/SG3AX/fVGAdQdvL4R4Keu18R19phoGf2aFqsNp8+UC
0eJJjwyvWUtaRcUCF2wQ1nt2tBwUM6HeUP12olmcDOK86tjp5QdFBcOYNoGDlVWi
VEmx/aPPQsG0/IP4fQl+T5DeNackCqs9NIdOLCRb6jboI69jGRl4r4/CjdnjvC75
AjQeKqPCjqsCx5YRjQyOSCsSesQjW4NKcsAMw31+Q+w3E0s1M22C/Isbgpj5mG1X
nMMu39/KiNax9G3kks5tvZaC9uEpLX+BEidGIAqtnFRedMuNIkTCdBkVdiQgJC/U
xOfhvVRMWfWzm8W/eAlN0NxJ28ifQY+fBzGUT+t9C2fIUZPeS6xaMMctOeMGuscR
DCa0v1Mv6BvHSD0GcoeaY9u2cNuIhr9u1Cfom+WCSMBzykWYrUngNBvBG24rKLhg
Of/Nx6N97YY3/zZjUbrj/JuejoFo9p+F2V4smHRktAZ0lqovY1g/hNPPyqXm7rDO
NMDkAWmPdDEPBVzXQlTimj6qxPvjgBw0f6SX+LU3ZdlWAMzAX8ypmqY3tV8G2hEe
22OlQlWx8FT/qNGmUT9pYlMahYOivO4DnqMp2ftizSXuNDjUwiRYRK6GwNnzC7Fi
t9AhIXej53SewKBj5ZRRIuFVEm6Qu2NkUquWyg3/6+N2Xke2HdwF3YEA7TkNrs+Z
DrrVX2UZEbSdQwjwhjngBtGidALmn+9MfiwspUP1vm6CgPULkJGtRHAudgnRjvoi
H6S0u5SQC04YvNGiXUfwBbiM71F5PnQMjCirk5xwMyIBPQzacTuLC9/dY3hovwqC
eH2P4wK0B/HHb6tDx+mHBr1b3XMXCzt6XQW5ext8oX8Fws6Z5DC5Wk+JOpZey9+K
6c4rnvyicN/PUfvBUdblxS3IsvvvYD3B4uj9DdUFg+qwe4KU/LzlFftaSpj926Ql
9VcJIYGyHslb49P66Mn41CsqG7bQjSyMKI284jAk/knSyvy9GJqUV9vp1+DSJDpu
eORjcUuIFHtJ734Ww1Qmmw1J6jhX/hL/mKBJvUJjhtdkHlGKtH6t/bpWePp6FQ98
DiY2Wpbm7cfUWUTA052gucddH6OT+U8Vnj5F1BEiWedj5aUJsaT+hQZwks60unW3
u0FjgMRN2ALWW8WRzVuyPbGf+v7oPI9aSthNUYP6Uqt2pQLxAMDrOaIyPwhFbmFo
F11WCGn8CC2847kfqCvzh4nCwctNwxn1u3OpVVfQHsdIyHrdmJ+0BeK2F5a8Eybh
lXz5uXyKacxFNRfghD1dLuyvJqNCtVlYs23AYhx4lzg5qrFXXFaELdnDBJT/QWCT
wxthCzYeQ2u0WJQi/6blhPSnajYGaHzHIFpHDjX5XDMqtvuze6Z1xP61ObjQipqT
uffa63Wp+qyl9yMuvh30H+dkDJCpJfD0k7KHk7/IoyTF4dPLSoFEcJdu3EwwMtVJ
pUPTjmWYsIuPTKLfTGvHBMh8F3XH029dUb7G7nmdmZaY9bOkHlulSc7SvRwuOPSI
+z1wfKOhqQxL/jVt+N8yq/SxRSD7jbxChM2cg7HTeYfplfDNM0p2KNBx83cWhpVD
01jXD3yerPvVq51yPIlKMitgU6n2yvxNhytHvPk8kkGJjAwuo4ZcpGB8yfPI2Zau
ix2QjS3Io4W9vJvdkBaMtr1M7fkMrSs1Z4dJN1ovPr2C4Oy8FywNZ4tfU9v6tEMv
fbV4YmkI++UF8JQ8o1+11VJYP7raoJiwh0/47Jx5MoBTMSiM2FaPmr7VQJgegmzf
oPq3aN6zNr7H2Iv/KTSHGsxo2gTF+IOZsO3RGy5znbzpsin22Qnd80B27YwyZw4c
fhRuhj49wGCcUiJ1Qh0jqN37GbwdlntVNvv+/moEbieIL2G7Spmg8xJAEFJ6v2C6
DegflZzDkkBGFEo/4MxahA89A2oNJuDh5YGqPC4KnczvJ15iAAWenChv76qb3hSL
MpIcPoR+rkK5zXDTKFHxvg9KaYatVH0SEhsGJ7bm5BHz7SmEK0cnjq4VCS9j3qdb
OEeJ+iYW48lZs6IWjNpUADYgwfIiqmD+WvCYz9ffmr3h1nFKA+P8k+3zkn9RRBmF
oemHWAnOOD4AYCZgjZqoFeuGzvrxB61FQHT9k4EZZ4mD+NC7dIBpDFb9oGRLHMHv
2OQ89/Ys5Aa8JT66dDEKLjSJp1xB8WnaE2g0XHuD8n6S8p7+0baw6/tFweZKnLMY
W02vQMOVwp8i4uqs5uD9RDk9KZTR+qTxseT9s8uIih9efPm834GXtMaLdGM7PRMQ
It4txDd9tiGaWCPZyYVbmmdVYKlBv2tF84jfoBxiVK45/fZYgXZS7KUteGF8yB7+
F2JcXGi4ZzfDdmiRC4gtKUsB7Vl/TEvDpaONVS5l7/Vx0qiIP+47Kh/zFFm8k3oO
v6Im0Mu/wc3GnFJGZult0Vg2rpgsEXRoHpah2n7gWM/NrkZirP5RuIg5DFjIi/WE
FTeFjfVkWb9BUkpDVLAlTrargHFo+WudnrkSlOWV99AznifxcmZ6BXgTVIsl1f+L
c331ausgqT0N3UAe3D3/R6Z5J8cM5Pzurx90lZGZBjxiPWVdYFpNf9KHPCcYjyS9
Cfjv3N9I/rbD2e4OPEqPlawM41YBC3rk7bwuLp7V7sWCGWu+8T1OFNvm9U0ZMVEx
j9Gr0CgMat6ei4C7KkiP2FGVZ2Qw5lEc17a0Y5A9Ikx9/nkFNB6Fc9aRTFZbAXzc
MDOhWdFhZKcDgOM+Wii+UH9HJM1Rr+hXxo6imf1U7tS8WJb+IyzzIjLMC1iR/SkC
UWmKKDHwl30sH0iM4SMmfuPDTticQbmzfbPJVVENNRGqUKjJa+kYmlMDK+nUg67K
WOk4CFJA25lGk5+KZx109UsavZVr3JQqZ8/OrrduGmJ9+LuxEAoe/rmzVRUYDcts
eCeOsAohWO4fMSKABVp7qT4Odc9f3eL2TVbijFJnPoGZNbfYjAGeQb6xqZTZJ3oN
pcwMJw7MJW70ZhG6iGRdiPUo3I1ghAqGTTWOAZUs3IDElb4ybVU5wdIIR+xDbn1C
S8CEoUP9HDMIgdQSRUisqG5ohbr65alnofsh8sMV9wiA3zwPmms53YdDZeuEcPs6
09KsBikTP00YdEFR8RO3JAD32hqV5ijju0BJS7kzJ3VYHDmHYli6tK/T4CaoC72E
kjxSVHwgKOlzAIjSLgGnohPX/TvPkJcIhp29fY+UGgobfS1KgIH1zwoiNBqJvKdP
4NRkC/Us+lPxFhQZVwJUvFDftHITQ+3CkVPzeHGI09qmiWM1LUzrWxk1auJfUjuJ
fNZYBfZgVwA6W5I0jlYNwkOpXPfPUfN3gZdsVI7qjyLa3aGOy7MKT2MOf030teXy
w3meHupE0Rqexka7z6dEjgPovzrhpUrUyd9RkNfcFHtAUswwCYlDB3QHycj8e4Bu
2TW39PMHzYK8vy2Fpa8rtkagb45CeClI4dZ5Bul8lJGyj3FQ4WLDheBm59MsrAIK
/mBcP+fZVDf84SmP5ks7w7K98BgJ3ku9LGFxCvPYGlLgQ9FMW2OosxzoNKV7Z/Jx
tUr3TJ7wWQIshbkPzeWZk+XEHM7IzBcKDrOEYk590lA1eqPKV5NEYTs8Z5IACo53
Y78StjIKiWsjQbCcG7Aivo0CLMM7iJ7VqPagVtrb1sVp+unXljvyGEWOg8wY9Q7Y
x2gMW1WK28nQ2MdltukXyUDZGLlGxbOoCeszMhmWo8FSHArrmM8pHeZgG+dogRn7
l22YNhu/6OB26L1opLieSLE5SvOI/ePEbDFniQvLobab0iAjKeDNtV7S8erJ/CcG
8+SIdw61o0xXMjsk/JAHvxWUE2o03kuzDzM6qW8zvQkEkuoYBrjAUOuDbd7wheY+
hi3h/CcYO/sctY/XhcTchFB12up+Wb8VlJThXUUdq+N5XwviRqbR1hHdBURKm1/p
RR4v0e+lEOI2+6leok2UW9l/1KAxMLEMgT50yU93rJMGMfqzD9O38K07DWEl2uBW
hkvzlXLeVZhtF1cjBx7AdPhmiyowq67/NeXLwc80DeM3gSurjBnAg4VNx1AOhRZJ
wug4DUsUtaLUG2NQemLI4WhV5NtSxA0kLqKYXNvM5LUUU+hglcCVRgpkVuHzIWih
CEbxFijT30uOuYV6I8yLf+lmUPq7+i/hBqCr3mwjn04dK8RvfTeid0QBiWy7fha/
GvKP615iYN9t2k7XtF+wdHOBL0aNwyqtKty2lfncS5OBJZhlqyotSRw1YnNu7Oj6
VItu5TFyedYGFtWtsarSzbZVpcn1GKHYJp1yNZP9ebPvLS7HKEeuFjobdxoKwqZY
8t9og9IePMvz2gt1hVtGYWiJTWgk1bwtstT2ZuE6lkYKPYfB86UTJy9zDqLikvNc
0RqI+vl9NqpdGvKRrChnJi04fILNnlDt+1y9yRWtETi2lHsHpNjY2LcGcN3jBYRj
qCnCm1DX7VmNb12/5ILq4cf/cb1dcYqJTFAQgedCCaoBOhy9JjBo25o7rUGE+XXf
wk9mnd7dZiYQSXsPVLABI89KYeCl2s/AiV/tPROHZAzcbQLmEn3Bab//UxdG3vz1
5NCisrBLo6An3MjRjmjEbmTayVAj3X0mPmWee0/bo6xnuc0BSa0GiZY4KBre9neI
FkEABFWemx5IhFcgn4d7fHcIZUOAn/53eMdgfYlkZIfZ/CJIgOrglDVdd5voubqn
5afNNhNrZvIOVP/Zz0OE3ubIkiAW9OGiM9iNxwC5BeV8586yyss4VsT3uNKZ8Uvm
ikZ9YrmYpQXU3cfG+HB0zRVdoTmKIA56beh0G+Kg9po7UziTnZaJKT3uA5giqg29
sKJiHoczJ5BEFRxEBk1fH80XdFWlGrGDrXX5de7ImkWDisbx5eRjRLRoVZ4lVFcG
p5+/v3mAJF+FVjXKEMk8NLq0xyn7z2EkisXoEOWjv4rlj4j2YdXcyGQuT2EuR/Mp
n0dj7XP/zkjwGPcndMp2RT4hI7M/2ymk/XFyK/cfEo7JhbnWbcWCaY4OF8A3c1du
85rvL+SDUwcbNlK1OYXmXwiCYsmPqUkXifhf+QzRzPa36RplsqH9b0G7Ag0jckV1
F4Fi4yt9kEaw+MdZvqigUGaEBMIKhhiQeiCqutCQJGtw911t3a5aW7eYqm/KF3xd
dlrYez9KHx7olvKNa01Q95uArv77zW4e9EXGW9cJuX+lqecyYBn/ne0eAn8Dftbm
cd1XaTScusOmyWsBDMd3J+lojP2DavJdAE82VByGTdUlmWQHrk0EBEXmBgf45Nux
JjBQR/kQKjwG5npLyhJUdAZHDwMXlUIpUXVWPWq5Aj1IPOgrPsufhU1lLaE634e6
gRCcNlSwVw2uMLRL+cX3rgxtH976qkpkxck9oO2XHfB66ZbNIfXM4PqOTC29kp7G
iusoJEZpjg98jcHvQ80MDqk3KrETGTTH+WMoqQ5wP4pAgrqVthqGuDwZ0YodbbHk
I2LEXhCeBychwKKVjCxzIWIo9KFulieVvfNGSsAYLOzqZyR7/F0G/S8cJuO6a5tA
pbb7gi4iXXC2BVxiu+d4nmbJQphTC3gSfm5asdJ+RyKio95pXrGEIUAHU37ce8iC
x7997/p8eHd4MvHUXRagt5W1Bn5csoyToZPehWZz/DpKsmhAjy4jM2Ti/6MpzAOt
BDI8YRL796dsUARyTxOb+jY8+jWEG87Yk958FdzQ6V5a5Mlq1TMKgOHTqav2jczv
FflHU/RjTQhJ26iPDSqZc2e8CPXUwyr0PRtwcX/xv8TFH3ZSCEMONBtsW8qJYVLx
w5RUTGMNoY2nlrUCZ/SQG/PWxg1YEnTZaF+37xxCcPOioqGD+jTWTxC5OTxZpNlk
dLClqvLrIOixr80zagsTPKUKALjdWVnm1BpLKEry0zdIhq+R6wGsZAbZcVgwkrmw
AonSqWoNGHw+OCrYUpOFzzTMcPexs7Buf7qNhxK20JtDdYVj1l8baIAvd87Xycnb
oUJKavwkUkfhPMsRL4e74XvZpGVknpfjf+PhjDtjOCrgexh1X5GdLRt+7WS5U/qd
q4BgN7866LvRr0Z/GhFriy4Kl7qAm2nArVBD7nfXLsEbJZmiD5Dsk8QfGbRxGl5g
EVssGBCMd14SY8mfXG9EA3kjrsIYf70SphHoOv1mS9UWYycMLLhMHcr4Fo5i341G
uKva4vTfXq1mLngzQxx5tIqDd+gWORa/kthrBUKoPjvXoTNZz4KVBtJOopac6PX5
z8z/GxcAC1pzEHIPSU/1WS31A5BzBCByCXiS2ElEV4nw9LulwdDEXEFbtejuicLH
BdY3wCHOEqQpwsuVpaz3WQjGonFy69n21nSn9louUV6sptLZuQmh9InPXKqJMLbT
S8oY+9ICMujjCAVqOgzC/hW395g8geu2lPyZl89XN+F87X3RH3B4EKG0Wrb6dgtv
vrSrgVowPMryXN9ZIkxLDUkZUfrOXF+8kIVs9iuxKRPR8UrwXxD2Svs4BZSj6EFZ
bmu1sdXRVFSQ+jNR1KEHvyxR8blECtt1oOC6sq2s/beZoTbXjzsQqamxW3RlfFcZ
MZ5TECqaM5c6cdOmTYD/G15qsj+ycng0AfnrHkUe/zsglt2kG2A0/TuNaQlggVym
hrdfp2gPfYg0xVx5i6vMZWy6R7RZrSFM2/DdOueVGQrpiz0SAMiMevRmP1KmkxOu
DkEXfajjaXZS4r5EH7Xr7Nn/vs395u2TnCFT/0VlLzkSAJS4bOiIUAGGyTnzk1R1
7K1QxczVBpsvbKFe9jNAUmHHFxL3kQRjTcerHixNa24hns8dlTEFrN3nbQ9jf8Sy
F+gGjlnJjKQIZMGcr05ZpA4RffGaYgQ431P2vxLkOAJp3MGWnYY119Ua8D6oLkAW
TO0YgoVV7LsIAKitFIaarK1fUjVwF4ccGc4UKE9FT7Dtz3EJgnszdybgjh6BsqHO
HGolvbw/ozL7r0DzCHn5UwGo+2zPP6IuvHXf6mPoGsnvzePcl9/tSFNU8AKQOYfQ
SWSh2iSt94SLGG2DKey1maY2krCZZAup1u+BJYBL+u8vM2i2trP9GtMAgoZeC6Z9
aXypM18AcpnB79iUdCFgOzLp7YJ66ffNCs0svdupC1tZ5zaiXWoq3njDDivp8r0W
XzgzOQeyWE0acK+opfXFaTZRgBfCJ7yoEW3fI6ng4yeoXDErP1laIJ69sSo0lSNn
gAJCuOcjMXn6/y///VGfcFHDghVkw0s0Ewgu7pSEs1WBsqZ2fO417MkBnbyeuU6/
Df13roH3unshzvSHMYTXuSAUPpV0ij1Zf6OFxWHXbDozy5jrr+L3K9LFE2e2vy8H
EsUpL2VYyv5Hv7Suy9lwZgjazJObioZdUhHsipJtdXgM71tQMahZsZPnwqt7fC8V
R9AqrZ30+cjiRlPwfsT0k/bT6S1CwWPeHacZdvw5mSUYp2v3/jWn1pD521JgmBaT
3Hqlxe+Mzw1aAs1JPRJEBfFCHSVCT2PQFBUbV2Gy5cddbjWFcHomKnB7NvzGb3/u
JOleGTO3rh9+QiOW2C95BOYdtxvPIJUvXi/G7qkrn97tKLmCGYRrkEIkGOa374+G
RF3JcRur74HGKmHZK5EF+rpAqoeNwRvrrscAXmjQTzCJKishWF4NNfZlJAjxMa5a
ppHG7gDwlizGJqxR2SSTIewiQqUvjRZX9tPpov0+O7al/IU0jt9yZ4JQqDCFdZHr
a05nlF0lYiN0VUffFK+VesHUAbIw+R1BYV038jYVbjOUoD9W4SCTDIFIK8vvL9id
6eLKKU22rDHqw3yog5VVZri2tAeM7FGAM47ovxhbmDQpESe3+est0LOykuBiQ6WC
ZxrLWyK2evSnPNOFcqyZd3aWlBtG4kxDP403qDRoUevyewJPhmACSvb4zQrUHaNW
91hPUsWpcUBpEkh39/hXJMrccFCfNcGhAlhMfQ6FdTZ/icuMCuF/FXMholXUGSMG
iz/2W6adWt5+XzvfaR3pgzuLFG54v015PvTJNWQJRQWVGqTufVnXLV3MPVRb2foT
eaM5cKbYp8BzGVA97ZG8F1jTwkI+jtIoZ5eN9L0e80Lupg/XfSX4awBOjLn7dLFg
O7EaUR9gAa+zrMBeYFLoV++Wma2v+B9/ujFOBJktfZeMTNSFqrnXfWGy6mfEDhZH
YW1HUfT8sOitiIgoAwYRSKmeMUD7swPS4kO17RLzurZ94bd1Rbz09e3YCHRljPrJ
Mv/B0714gwAq54TmGwlgQ1pziOvGxkrfqxNoxDTPR/EHFwo1vD2XUx+UdUC5Wxkn
ytvyia15UqVkiIcc2ghig6M4TgqZv/mfbUBdcHoh+p8TFIzkbvEAZTRsuR5dzJGe
kjwUhvnyDBOnni9XjpB32b8mZ1aLzBOkCsZCKkn8EtN2zmcNFkWznzCDdg60nXMs
XRfdm/MmD/2qQXegSoevv2dttfAFpwLF+aWOtDwrIsM89ihrEeMm4dvdiRGuoY7l
Y+on5JE+I+47TROWdzyWHyedJUP4RjrBfROsg1TyVpQtIcnqb3MKh3hjKjNcuvgn
wopTbeeRdwBEtmqRe+HCHyDzLATeN6G0NT9fDKhJwV2jFtjfV+6npLMXKzFHW5cZ
XXmGRorpgWVU1kLvkbmfjqUCwjTofJ1NcSIRKDQuT1ufL65xIucAwr1YqejnvcEl
Tx8zLTObHbu1MYYyv3NaOdJEHk6wMxPsP4+iJpRIpbAVLptm9mO4pResVzl03B84
8h7nvwe71ViosQyNTiDFbsZCiOTOKwO4EtobroCZa00nBH2Q0b99x9Pm8Erw7+Nj
oH8DrxUmytMD1Ee1mu8WWN4Gv/o2NyzwVkxR4aGKlB2FYjobTB+F/dGixR+RI/HE
EAftCWxzhYVk/l2bVLUzxspHjIxGUOJ/fVyOaKdn7/8+zenbGiYF2jWD946DQulL
9yW9TqaaKD6/l9DXQAYwxwwduHge5fm7Yi5CjGpfE5iFCFtJ3KXUXE+3HjCdwIJA
OGo/NqQUtcsGYc0ULb25+GEL/ERxDR+v9I2n5nWwspL7Z0vnnDYO2YmsRab6cvke
huybnBkTLQIL1QFJVEJ7knSjUWXyPYf43wmBZtw2dM3cQzDtOYHPAu/dkTbkiq70
SLzqjy9e82fttB9H7+KLcVNgMm/OUhiLApdj5Vt1HtDPR/iydKWlNaCekpKFubGS
ELgXyKcbKY/89Kxk+1+ezV5koThawEZkJYTJLrhQD+BodSTphE/FaF19H6dJ0gkO
1ezm5jQJhcERx7TfhHJr7CCjkpB4sYI82KNvEa+4zMotE0ZmF4coY/muH0aNFzEc
qZPNcpvt0VtWpdHi+wcDQedi6bGwL8xAN5SpPTmHZpxpCpSTfETw2t7WGTkRDmpW
rboqt7cnGrZIqZv8Ax8++6J05DuVEMy8YkN6/sUgBY/HQNnfy7KmWlAM65qv4o5T
52sMgxZ7k76ZWlUCRFptZsZomsbaSBqxOLb3zahTx/p9G0JIL1qmxnOt7amDTq1G
rb9eVWmFVbykMcr5tMX2cy2ptoFDr8gx6waY8iCE887kUurUYRZSH9MDXrIdgcJC
Gb0XSjoj1xfEoV6JhTXEgEuAsSHLT2itnInoxi+cyzycbzwJiFBMBkOgSQ9vUTA3
4hZD8zqK6Nu2SQiKu9zN4hort/EX1HFtXqUQDlEH9ix24hQ5aVEsHMh2UVAHlcB/
yP77P+OTUZaasgm/C1o0qeL+UWkEIuqG4zEH3XrdLmch873lbblqcEH92hw+FeOy
XuxXaQOaLuijHcgoebeD3J92R/6DSuipc7TiDJR9vxsZ+uUJQ8YPlZ68Lf81yw95
UxCqyiUc3IIpKbCMX1tjw/snqV8ijUyJlZ74pCkqLG+wqVqFeKBhYPuwPQKpm1vZ
Nz5NONlRuHxNCCBaRefrc+xLVYIUusCFcYd9Yim3ql/0FlAKIIYIgqnllkQbWXDR
EErqA9YPevlRxEPvuUA5GB50/RV5T9xWiIghU/JvX3z/3Q7BgmEO/SC95XOfDKbK
CTWbKermJlK5LHzcII68fsBDi7ZeloToajsNhZ5i1L2UHCIZ/WhjxoFY+hfAlWv9
NA4rSZRtZHALlpNOYa5kFPMD6l5w9qguKNoKULgwfZfWoYOdHDDQEaxIhuipNZv5
RfZfZp+CAWHNwhIqS2CvLoutfudBpf/LArnfTxXj4S+apHOcEb64BbptKfZbz+rZ
CyjROumqMEQi/DFhXMXMermMGVrTY/PuaQs1bxoH/+7X5Klb3veGNdfOTmOvLdqI
HpvWBqN4LsWt7+HXgrHfX8DGBpKyL9pigZrppC4oAToYT/H/M/eH/cUG2vY2YD7O
h7elW1w7x2D1fPLwe7yyTBGSViYGkyafno7Kq1liID5mSJiYbeJp4YiZPqwDxsrv
RW8NoGmE8vMekaQngvJtt3NG8T3EGycKYfgn8H0ZOtQPsEUg3ppO4S7LSlGIxyuF
sdUU8xI+kkbX35uco3RmBw15We+WDGIYQb16hJNJSTUEnmqpV2LkZqzwiS5T05Cq
ly88qs4jMxKcOVR8aHYqmz4FeMNdpKkKjX0SyLP8NAnxz2KyPleBnRBPfLxRQcJI
WpToI7abNqoJAeOP0cRcj5hARQO8IeeeXakTLu6/nugnP9YEXSXI8g/mnF5E/ixK
QorlMxTFBxuqRqr6aPOIbSfJbknKBZCijrN7CQPZD0gbCc2ahym0FpUU0EmtAKbL
IAllxGu8a2WN7U6sIM7h7abwYQCMK+IFIqPLE5EE/Z8Or4q/k4pWi4fD9nDtsexQ
f0vGJeli/8FPRl8YOVOeD2Gwybr36mjPCQA63tqtxBWrOQKA6e8huSfWcIFcibjO
Z6peDmoGS1AXP0dYcGiZ3q0XHXHhYOANkwiLeqAv6Jk/yudWava08N72QuHKEGwo
wf40d8WtmlA3QLk9kRnp2DevkdLEZAjF7WFKR6Lvc1z7hBjoQn3v7NkLEtJJeCRR
ZT4szh0XKhWaJ14uLEOXg7o8ERyj7yfDq0N0YNlShaiWunuX+ZlOl+UrVqbo05XI
5DxDTbmB1tI3kF1zyUC/bFZuTKoPOX8xUgYCmU4eMBBeuP2+Ky+B4k3DxKvQp76I
wVtbVUxgNZ4E0IZ+xJc2Sj9IkwVZpqawpWNH2Ogpa9q3gHFrHCfGQ4FPY1KBIunf
Qs/x+4jeRvX46v7VKey4EQ2IMjy+sTPG2kfJkjDAA4/aoe2WH5+KsSqAcLwYSDZ+
1yXC9LS08uTUtpWpHAPoJppk0lFxiAvYVLUr3yvKYwWp31ieUKzXFtNcuzVhvQnR
pb+e1rvew0FfJPZ+LKBmrqPYcP9bv982OIMqAeebF7fsKX2qhYB7hUGggY7WmIoN
Wslxu1COS5XMWZoqStGz7kpofZuV97G3R4ep/N6n30/z0Xjlji7S3dQIe/nIiC9Y
S4NnqhL1GSTgkW11wnAHWR+uZRKq9i229gnMhAXh5oNZdmJ58GKfQ1hlVy1LXW34
C9XSSx+T3Dz098ns24xSTduJnX4bjTAgtGte7sxFv++exv8W7Ui7iXGmJS2SYg6E
qJXEXsGmze1Wk2HXgzrRkmyxoNxrJQsPq8xwvZ0GcbUvRgs4iKw9e0Om1WKQXKGD
B2nGFgZUjZ5yNykHgo5hdG/m6Y/PFzrMfM2j0MgOOuyStNNXRgxQ1JoGUDCQ2pqP
DjL/d5neK8IjTRcEQqynFmTLYcMGYHQHm+5FuTYtrXG5tNMp4dg7NWHsvbaxvXhS
EW1Ba9mQ6DiTRCUXziXNTjFethBO7/U9on4/6ZY0AW5bgcVrrupkO1EmF3bBUeNJ
rfcAgwMnrK+2zHD3TRYZx7CeVFnbw+J2ykr9yKZJWTcTPPrvLVwQ836ijNgGPgs1
A+7aqYEKqQ6iHYqomy8Jp0seQOORX3zwlzLtsWhJyjjIKZ9yc0/hEDys3Lh8H54i
WgfQWZ0SbDChrFqlI8jUb5z/0g0Od2bDAIU0ESnvopi9OICCvrHFShMqkwVF3JS9

`pragma protect end_protected
