// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
CcBV1c1twhWjJF5xjj52nru3LZHdEh1RSAcOgMvUuNTh8zAvnvqHkOaUavMv
+tL/SVVDEIT80Ed72sH+06t65XoSopOW3xjQLjW5H5G2RiasWE3ZUtY8uXnD
7uyGrLsHo/FNueRyYXTQC6HPOCAehcg72h0yD1glleakmNUoG+1iSqU7ifEn
G2uxqGNLw3WSrWs7u/RjMD7fAlJMCdX6Wz42ecSamnTgwQ4ckOwhlKdzeuHR
uHAHSVD/HO+LvMsXtkpXhdryaoxvyUPSlIWw28j8OquBWCk9SBn8M7seo9kG
Os4Ju8DMDUFZVqilp4nFnyheoo2bXIapUDoXpC7TFw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Pxo0ptneB5D0uQCMz/VTy0IqzH2Djh1FoLskQ13Dv8lVaiA4hj2/9cvcbBoa
sneAzWQmxwrGZPuLPT7ZMD/4o3z9hqYHlmG4Y8fQgAvNbOcDR6i8gRjPP6c6
T+EgBIpgpmVbS16lv88zCvbYc7XVUcl1I5XuYcIELO1VpjFAT0ljDLyyiWUC
9+gUlHIxJHye0fk6l4Qyone56XOE0TPmQWgzk9vieDVaJb2zWj9/hEcTVAOT
ZBA11Ae1AqHb4T+MqM1ZTMSguW6lqZ36UTM2KCQexE8EnlFtyOilOPCUfRQX
g3NBed+NGDQqVEA3U6qt2sKYUxr/r/vSTuqXvRum9Q==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
T1x2uxu/Lnzjms1sUeVDmTAyMJz0w3srTXGodoRUaV+mfIU/FQKkZLGfofRf
XLmm8WyNP75B6AdFpgtO3m4PwVIXddhPiREwy3TS/Ptl0i9JVc41Trfk69dF
lTTGDN35cFfC/UuyRmXRB6Gj1pNF1S+0/jMka42p171do0JbVhSWDIVawKC7
Z9WyXiz6fos2DASZDFNd0kgBOHaaSKM4BmuSvZJv9Gx+rep1Ccgs8bY7Bi/Q
WUuexhSv92XQvdu5H/e0l+jFyiEpE1VK0vrVz4S+BzNRqO2ab0q1bhd1Z6mo
yb8HdU223ovzZm56mNI/BR/j5ViS6Ay/2gzWKXBwbg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
QIb7S7F8qigPrqkW7b+YmbMjQT7hiTeO3xQEpSvHhjPDrxVrDMrN5aNOmFSu
3yWOEKYv43ybR0HM0xFyA3ykGjz1vzH/3whi0iM0VnUnMSEZmScBivUkekgl
iVw4wOC/gJ4k/u7atn/inDQ2euZAhwYc3633Fh1rnZ8TckT6EA8=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
SVAnSL8tpnAPT1XLsauTcA1uDeoWqsY76zgi6+5cXbUv5W3OSoc3zEOxvZoO
FKPDGxaFTJBoOULEEVJDRSfZHVYc84ufbiytRr8g1qRC1zgJ8uP15yEx+Fli
ypdZGhLks+EGjdZEHJneIbFtvc+fqwV+9rFHeHNEjCTxgrAquY9PkUNEl/MI
JqiA9UdN9J6sLIl+hIdbh9JnagUuXIhcdPoTUkb+n/NBuSMWpbGBpkmteKTG
yMVRTOFwZobpFcziTAjxRKzjKEKzdH7Inxmuy4ceL4riBC83ehmr1mRf/hmR
vZD5XfcGrsW1XpA7kiJPsZKETkWarZbI9A8np8+DOE/PUNBUtVQ2KznH6miw
dzb3rbBGs9ytlbKcOJR5iSn6MnDfyJPkcV+SojQy5cTvoU2eBD3ojriFJnyr
1Ym5Yzu+vwbdefvOWaO6vgg6dMflZZa9UNnwhuVqZLGSM4S4ZJ5TmGy2LI9z
sDL1w6gLX7zt5CZgzUpQMZFMBagCpwxJ


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
cDfj/1GhnVzDhZUfd5TTcB9WdTbQxRqbghEghaevBalJPUO5O14W5lmOApoH
OMxrg04XeJAm0Y2g5CvJAPC1u/sbhfcVK1GAH/qpmRXbbDodsuYktoli/ZQt
ijdFklaJtfYrorZnqUJZU9C2a2O3TyMb1juu6GFoXeXf6JVAnsA=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ejgS7U1egDIm7GLOqd42jrnUISqkpmK+CdOIV42fmiHLIBAacGpgIzJUxmkP
/aDJRuDq8qDEtQhUIbx2UdEvoXaWqQFQWCdfOyLs+/73FQIqRsfuYcgTZybV
Ah7n5OMCqqjagJqUDfU9EniqniL62rfDo/AGBjOmTWRwY0t2cvI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 18432)
`pragma protect data_block
7WoSY3IbS/jHomm7I8a5Ew1C2+ArAjrTHzGSp+WJD0H2hbgMvz/OYRFPkZDY
tkInUcDx4ary1LOJ/QtIl+5or2U7JMlDXOEbXixGP/iGrV9VdTfjW0mkRyA5
x41RNIvgxnojBSeTHADMEuu4tR9tBOerH80gwYtrYPuBiAFQtsd5xKnm47EL
egxv6HETa23imSb6HHksC3hHU0jYYEUvck8GtvTCPYIlRvu7bDClEKrP13Ir
+Yok5MtWAy6WnYc51sOwX2dmPzELnt+cuU4rbfzhs7JsSfJDAx4ioUFiQivg
I1DA2wWVvjStvQa9mA2DPArwIQmVeJQ0D5JUirrXNMoXcw5dNWZjUkctF4sH
+YxBDZgiMoNWJxRZAqABrLbB9apJxd3UwW9v0nuK39d7YxYZdrawJQZp+Mmg
QQSK09Z/1qqFZM8N8zngQRQpYUWxrwq4u0aiK+ZYRy2YBvt74zUAaxSWnNY7
RoVAlqMEjn9oARRDEf0oyhCUShLi6btsX5t35OjQO4EJLb1QTEXPvNDA432r
saoD1FMJZzoSRv1VbaqmdC4Rbif+zkfQybbUg1qdOyHcooM3RDeTrsfKM/bO
pQBopy0rm2SsbivSJ7PFdzmdB5ojCb/VkNegdtT3uX4a6EvmcwDFVPhsEe1K
foXwo59kYLxMyu02ExxH0wR1qM+IRO64d8z5nBzeBtoEaMQlgGO8FCaNvKN+
XL9SgvZ5sNys++/bBcrC5F67QktrjghpuUxIJX1Dtax5RzFasJcuICmcIIhR
PsOJPzRcxzVOQRpdVZ9RRij/MF/od48BuFhNlvN+INkn6rv0suK2nVffxo+S
Lya/y3e6d6Ji1XtrepfQTOqyKyVQhGWycNIROU434xX6H2zE/T8ViIezSAOq
iwiEtN44jizKj4or4ISPrxkVAOCqp1WhtjPJdp4p2GJpXJAbbuCC5W9iMjRH
WzTZcbLV/g13FlsTlh+v9Mg/w76uIYQNCX+iXziHxHY6eOrT6iMCUp6gaMkT
2njFD/Gyfsf/rQG3lpvWg92MD3SbboceBW3kRgWwaSUOtB+KWhLkLvWjg9Ro
D/rewQT86DHR0eJY8Q/OfHdci32FFL4iEatw9iZdpH82x69U/zqd5BO8CD7O
nYGHr+gprBeQlbW8Dzm1kSwWT38tZuxkyVvn7gr2k5fw3bzlcznnz//Nob0k
KJDalwP/L36SFE6apFTHZpEFdln7nb9ZHFaLUxolcGbejprzfYFtUJzfFMym
8L9CqEqWDNNBVYMNDLSdNiGBQhGFb9N1zQuXBb165LnW2ypU0W/kDoh6DpDp
U8dKvUFMfrA3ZL3n+vYnUIyQhT/TGdUQ/z4SZo6VMbl20c+kh1/0NrEnc00b
r2Xyh4pug0Use/Pq4jkfoJFSm7HmAyiBDGAD9lspc/vjmJov22TYr2D5htHn
EDHw3n6wg5cF3NgGCnAX0PkdSYDrzdVVXdjsumNX1p2yr4uOGvirAwLFF/YI
At4fm2TZGEqUoXsRZUyJU+PFZt4dymWWvhWYVzJLY14WJPI9t6ByYQS9olup
bOJVA7b+b0x+DLDa7Z9QRjcCQ+MK/Qjco9bfEWlSe2bPcfF9NkBqFnB0sbUN
kLcwNB5DXlDprS86kYQmBWeOmoAv1fq6tYr/cap9oSE9VZpCcvwUSKay3YNW
xaP3R+3pKLAfOlg3tFPMg+bbH3e8fcUMK8cxmIqAeYMviacrmblhmV/jbsJ9
kJiRPwzk0o3xz0KfpkDqzbPjDD/omzzEAPFQJ0/mmro9Uo9W+t9x0CW3OlQa
PtgG6rpqtBMoE9T8W0yZa+zIIBjUe/JlhvZHobjxU7Yj41ELoas2jPJfg/tE
qv0kJmRMiDGVGVRG6Rwv2KWu7mvA5rLiEp16ymhh6xVwwt/g1IlkQHUhZ1QT
sB0kYqFuBcO8xe+eRj0aPIpHN/I3J1v3mieLcEHo+dPrdvNdR660HqhfGblf
xOdI1YoX6TkbOCxNFyJ7vQBJKG3XLXHPLTjcvtXK/pqfHKS323qiMSvUqAvp
ShXTGS7QhEoi9iP8o701Lnc5o9ejaxFeOt7zPs1lZmqEv+gUf9fF3QTmqeAW
4YaYOfxrGQy4V4qqDDdTfN5Mfy8rt7sucz02cX3MeYFhA6wfVEvTWcUItHpb
3VebtsziGo2oSI6KyZX6P95drexnZWbuZML0RW9+4WoG/D/F9vHTYMxU5kG8
oKDVsHTZZTKKfAPEzuOxR0pO00mb38KAMvERwMFoSkTrUeF7qnYjT0RKnfnI
SXc+mnz3kg3OcWvToMq+cb5aXWScO1QsMnVPpMkUUnFgLYG2q4kLkx88x4Vj
As7Ao5UaZwUQLToHyMGdJBhywuZ2kh6ULBosGhx3/GdQOq2FpSYkg5Z5rbL6
n2Y6Ujz4kNA0TfpmGY0rMtWpMklUS6/PzPwhYycYpNoRsnLctEVScpTmrKBd
DgR4I2g9KNiT40aDYyNzpHzBFHWeyC+2CVwQwN6KjZMcNMswODFiFVTAakZn
av8bPcmpH5anlKhNj1lqne0SKCcgYB1qsZQyisYIFqc8GJLMixUOOKZ4VuVM
8f1AnSZBnBAaGQCp5Tz2ptTH9wAMbN8dpvDvVPqx5CsSt4j6NVLfEgQWZVTQ
ubx+AE0liwg8wm4QRT1n39FGWmA68+GmdOdKrXEc8MuBTLdIWSEamvIFJJkx
klQ4H6xAdvpS6LhJb21qFvM4bQmMlQRpy6puDjoIICjwlbyW3rMRNUdbb8kI
ax9x3279J93jOvLSFFpeoBO/06qrYHrB0Py5XV1a1GOamyqIBKOfLaa5PaN9
TrzM2eCkYzq8b2TEyA7ASd73javeoCu/BFpaxtrlphIZhACm5qTl5QB6p4hx
hUfeAEWK0FFk7+QYTmqfW9Abp2WOxUvuvRX1nmOfzC86zS4V9jmkVwKY/K+s
JnEeP8Y5p1g/I7qNhCSJWaWvvMqgTjtBY2XubXxMPjru7gJKAwAoGF/zVwTD
Zgd53E+S2V3+cUYRzmGHM5q/DUJ5BjdyMVhcQrdN473snYUlhUgmbJ8lU/mm
iedGaWdskNOZTc5FDD3TAyJf9ZloHupqkRM7XKgBgQcBxmzIHPSrC0Z2gWdv
3F6EIC3tdFqtvQJs+u4T05yGXsE0FZ604pvIEbrXj3liESPPL09V59o44rac
TUxP87EZYEbeZJ19XaLjUM3ckeNctMj/O3XeDUX4qldxql5236U+a8pK26wN
YPov7moFadMBzpcj6ld5YV8cTnSpp9zlwJMtDbJhzZFU/yS4QpOwckLtN4oD
hLUrKV/GbSoiq7qPlXWDlBzgEo5gu69v8qXTka1azATFBhfNxcK/UtXAOxab
bQvFpcvjbHB4r+e6+pdIRTDa6r1qPeMbSzyYOtzYzx0ugzvmHBEYRUnjUNgl
3F5kSKTrhk+B2dszx5NgNscb0OM1iOFhrkPbT3A95D5LqWxlXEnbOns/CSj1
izA7FNdbazbjBW+bL5G3BfquCy8cP7ZmFbRB+zRR9u/OX6kVmCTmFntYjy3f
GckQ3K9RNg5lLIT9UXvQtJMWzyuWX8G7oP3iohG3bnVA74nsgUJ6iNTL1ioc
M/U4NreOt5i4Q7FmxhNmPUjfOIMiZRScUHWi26rH5AiIp7fUtRjcaRhBItx3
fYGYhITO906OgoJXtUW4XRxuLuICj6RkMKimdzhY3eVx6Cy/IbMZ9nEfsbar
k7cLOL6MHJMo7mcCM60OEFLmxsLd+Sh6DhP0QjAsNI7757vCNxz5XzZMHW7p
7IYS0vJfaK01gA23gQtGMrJWhyGrbI3plaDL6D5OXtsjh4MbeKvIBwzU9xpa
uIGC7JrszwyZayVLLhjbev2hHreZsHGcWeFQCMGuzxG8zL8AZMyElozgkimq
jCPvehCF/seFxrbwZRM53sef/G2C0b88WBEc0zu+oKJ8ReQ585xG5/len1NE
IqTkgLEnyFJAgKEuF61A9L6GdIX8deM48p9hob6kWoNjl/2qx7+4IIN/2IpM
gbZaHP9m7XWbqzZWSgNr6TSVblp4lqiubK/crcurp6kOYgbTbbsdlgh7Q2f9
Rqmueu6Q4kMzorji6NUOOGGAzHTL2/xssR7wmcrbYDqAPTGVHXgpXWT9Tvg0
SVKwR2/rowm31uP5ZbJa6+7n4MNK6MYfajxNkxuY0pCzzNEvZY1hF1WWWwnP
AAEEealGxt2QF50rUJQe9x6jxDfPEH+Z3KUu96fPhkMdBKg5BIeYtC7FYCm8
F7c3z7DfWgfXjzFpTzD/6iD/IOYvmA/vZETzK++rtM3tSlZpbbLkDYJDuucj
rw6E5agJOvr0YcuO1X5mOL952grDz6AL++c58S1yXiG1KU1KIhTxko9uhlZC
l86uih8Mpk/N5lp+ISefiWwVk3J2zPTCaebWJcJzy3EsYJfN6UucAO8Piki2
s3eih3XilhlIBVTaj3VLlwETKwBLoxsGbyBo3HwzQhmCXK3VHnsNwBOTK37L
D7igkrJKELJiT1QNSvDbBo6PBclyTwYW8steR0I2hqn3SEGfgAYt3aW5SvZL
CgsXRAawfrwAaELwP16Hc2ar1MAOQr6RNLRIMvvggNdOselulVAxwOH55ObE
it65tQVFBrcpmBLBV5wLVypBpS859APMqwMjXqE4hE9QgSf9zMZtVbJHxhqa
ZSWQUST6AzUD4LBFY+lCbcDVo3MWXW40s/XtarH1wNSPGhx145AljF9wuSvF
3gamb1U+tzpPEoUOSZAjhO6AaPHPFwEyO5JqJ0sdMd8N5o8n5Zn7ZEmfMt57
Za/0iV+bxQvY+g8G1fPwXcFBu5Zd0z71psdw4m/WqEKFTdcYdhyofZNhM2ts
ddo2wozDXhtQSjOT2VOBYXo002bNZHgNVnQsJ/vBBMFZ0Sb7ruOjbOf0tL70
zrFmQjYLPA/cpXUn8y3jEpyKNL+6kzXHfelR+krJ6bBgHwXG8GJQTbbxn1ei
YC8dKngv8ewViTn01Bp2KRomjRHG4XfeeHr4dLThCPuz4GnrAbxzX/kVpfwb
1zEVv6hrh8K4mUEQlVz4d9+EZamVM4WY8LCM8LE7J0aSf84+U9UG7iPYokZ1
Cl9WffnvCeIjsuQ6pfjFv6HuDDk6Q71mtc0hVYdTLNOGmsCDxwgC70ZzJn/L
/ScARqs7iET5L9wOm61uH/D2QeTfEqXD0Z0+MPoZcIgMpJWmjpf9JeOqMFrN
+zqrKjk3sOgqIDRZ1IK4a5+23AaP/+kGxuM3sAWZtBMct4gwkMLy1WD6hNCF
i0AFu9NtX62rpz1b/EmFqmqkMUf2YIsNYveagDq2HqpoAVc7YhndWIRVmarm
gFv8/Pe+V825md+U9pZEhlhwB+Ut0IzYTfvteYLf3IPl2kcFDhKbCGaFupG6
4zidXTHV3fUhUU5ZN2sXhdhEhZXOe8yIaVavUdbku/k1S5Z5/DUYRWmlUrt6
OCaTgYLFNzbVLdyF3wPjBKmc9EOb0MTLNziCxn8mq2llqLsjCCoz0iuGFN6d
U1oQ8jeEKEZ8q+0JSj7dno3FafJZz2o8mbTM+Bm7bzhYfsIDVMECx4eJr1C8
5vkDWVspnYjBtj/CnORNZB7C2dUyGU75N2dhfwZnlA01SiKbkathz+R+eo3z
v+zghsxVNw13U0KCJfNKwXJ8UuJ+2xFocsRtt8xOxajFTgjrUa7KMfPwm0LQ
lRfRQHaw6olTTUx3MTOZjiYJS+JYpgi5Jf6wP/5Iqdxwwy4eHofW30sMlQo5
odfXbjcLrQ5X6FwO8B+SsIUy5VOYQ71sSGsFpL+zY/y2UNOQZDZDGr+xNVVr
O5g+xSr/FgGndGtIN169Ktq+JQue1wc2QWgqOdOlAGABZVYYZN/dCtlsKOgl
mZdwNRa2Teh4t0CA9wGgFBjutmamxdBqpEp4Qo+4rKaFxVd7QbEHPM92iEYk
9cg7yfWGF6EtjRxw6kOe1Vtx5ZDIsRgcyqxucVaPXswXfkd/+bs2OBJt+WVg
oZVl6yGcbAw/zG0lTI63UMaVM0DQh9z8wX4sQ5aFlyy4l1/rHU8CZyC5Wly7
rKs2UnSEpdq1v060efsBJU5DhdrnGzZ/EQTmJ5OR2iFmBmbk6lbAWVy3Jc1c
tr17fCnc+rl88QbbRoGCvlsXMHXGKztXfFlvc3q6rhk1OcspWNeiFJQB4aRI
i3XUnTy1RLdYjmFS7Xbr2ELEfV33B5NCaBTuTncrNvB4F1YYnoc6rMWHKYIY
ImpmpCM2D0kgc9NQIW0GUrzFE7YWJBWttPJ9jL3YpvoPGeOmxiI3/N3wstKy
0rjdIeN2LO5SnaSusOls4gBtRg08yEH416YGm0YlSczl6nxWjPDdkcNWVCah
AxGO1bbBPutxQE+Sn8pT+WHKvJDpgPJi12kr2d93TIhmgETtthFO1riKEXvX
PnstqSOMYerVowMihlr21ICuVgr94Fdg9Q9RQ2lgiZtl/dOQJeBph8y9q1vw
cw5LZ29ipjKQlg2JbjXwVg2uZcKRuvIgq7GPW1FJjuaHD5c+gn3rshPEGjlI
nFbD3FX8cf99WcULip5jEDYv5ZuXOxQgmm8algH5VligPCxe/1IyYUki2upj
WL6AYJd8dQw8JHoGTzmNPW911qw68lHbzV7S3Aut3ox/uijVySzJdE4+KpNW
Qkk7h6f9HoNkYbqAdg9CeAiRsBpTqbZ30OOnpD4Te/a3J6yl7JAQJ6F0umy+
90J93z+kUtQNg6FixtT0IR8mZU8ixAu5BwqWtTyDWE+b8bq0e/L+17WSrebn
b7tq0VzAQPwk4p+NQp9OJ9btW/uVT2c3ug1sS9YBxVyqOIq3Z+TSNO4PKE+Q
t0V6XDdsl/StHmsG9fPemzkK4sTcrvwwVoWnVSjRgTd1GxGXk/xuJmzfIfjF
5tflwQNX5tNU6SesYphMJuNVW8CA752j3QBH4vIZkrxdsrgZ4K5rKpzgwjth
8LXnTmxRthPIDzo9dPSuk3y51w+kT2lAfINeeP5nvRDo37izLoHj+GtMENZY
qvFTa6u9V7bmdORxIUMpkH94x5n53mdoiRpYc+8GELRT8giiFFXFC7EJjyz3
HzCLH16X6CH6F50vffhJUerLLQM35OR1HUoWEniLDs07DA0OqdNyQtKvsNoZ
XxJpCphhNl2vzL4SewcNLHJ0JKnT/S3krqiYaNL2N2ZhXenYtc3AmvukR1dS
osgDBg4UF/vX7xPFv+4C0aXV2t574pndKuZ5ABhBXLiknuCnIkm7uog9iiY7
pGtgS6VF+TkJzfgUZAIi1FzgiS3otdmK3ON56Agvf9xYll4gSSlztgkDSEAF
kjg9plbgq66Feqsf5fzERIToj0fFILVDbGVLqo6H1y1mV7QDZJAyFNsiLt+3
AU5xO87TlX6aDFZhpfFvNJb2DYT9GoiuV6SuBsZW5E4OERgyYOlJDWgxALS8
NSNP3az9+jasXoziXNXgDRfw9Xwmu4TtRoBEbbgHL6c7p24u17DTctvIslTI
wgS6Jenb9SI/apZP3hxl+d3q6f5fTK0LCt0uFG+Say8Qt4wl7WKdQoLjhlJg
ol5c8z3Rx91azaPM9uIFa72nSfKlnIFjvq0PqT+LhvP6+C8N027ezUSOy69/
du0fLUwg9Os7r76V+bMD3wWhEMtSxvJXvztPQAcYM5ZseK7pg7wkx2OEYDXt
QrgNFlGIFvucZt+tYEyPszByCAR/2buOi8kf0U8fsLIgO8FvdeVlPkjhP7JH
KLM/+A6h6GfJe9NnyWS+BTbS7cKqJMYu4kEgpJTmkpk9/vYHk4vH4uYWE1CK
Cw88BFb6G7VLSyDVnNh1qDMKrtZI75Zt9ln1rSKXOMPzcFK9ihQNknT/H3NE
YZ+zG1HBybsqL4eEnuRFXJ3bBXokRxppc5gwLpcMPG6f5JpQZKc5/8AnBql5
GDYNGpZeyCuhTK1aTi/leiofGbXYRrpeLGP8z467UUdXaPXRQLI9e0buXCJX
aNlbzwQ3vF7KGiVHrjn/0vMRGsttAOQDuZ4JiLDJ1/kSrcGVP5oYHoW8Krfe
28vyGiuRVonl1jb8b6iczSy55Aj8QOqqaYcNhX2tl7i+f0uJOIbLKp7fJf8J
13upfeYBTlXHCnmWH1fjE/QQNMJaILl2ZDtixnc07YHRzrZJ33U4VwLDFRST
6q8KAJ2opSQE6VYBtAeyy0QzwjmT8NekEMIwTAOOZ0I31BNz7pmsxSUX8KSI
f6xpTs4YLXh7SFKbXvJ73xfSErihoqZWs2AQOZQQfNuVPA0z/wrbRSY2gHia
1MFxuZvaSNPALBjPopJZtcmwjJHUSfyTHGMjWe2K1kpsyLKCWnk8lyEWjZty
LNsr4GV05msonHED92Tn2AsGcyVRuL8UVoaqgPgE5OAL+Z4It190BvrdThaG
YQxT7SNrayYSwozJppyl3hnYmMjn0YOQChYk6LaMcZrkcE9UQN9p2JXZD22y
E80xP0ClU3ig2TgNGTvs7R6BX9xXzyHtevQCw/AabAtw7DJ3HMh37h8dAumn
WizBtZsPpEkNo9nIU/iLUCpme0ZmdLWyq5Y0RkBWmEzY8YVz6/9wxWBDKbr0
1cDAEBptWBdqM6/EqRft6qt1sYoO35HGKuOzIP9Pbh+oY99No5c+13vq5NC0
dz1nLkiefBjrzDPP0QXJ2HTKA8eppEiJZCri/gVuZsSgYp2lxQ665D6vpfMD
lQDwOQ/2qrgHbNAV1cfE2N/I5mCO4A6C57h5iIfw4yrH6MrpEu8w5GMgWigx
J8rnMjhR5+hv32/daWWP58HI7rLezVi0IDOlOZ075PDJ4Z/yKqXgp5VqyLoC
6nGv3Wvv6oQy3e2TPPEdfjR5bseO+QUc9RgNzf3xKMOwSgIKRCnYPdPO7Srf
c1mABueOpQoUcQn5XhPynYG4EF4Z77ZxthA8fIu6hMz3xEi8X+QizhAI932c
BWw8hBgenL6KMvCMwlTFjYrtBOINAgMehGAGyglUXYjnRLWqpjt9u8YeNVkN
1wS2J3o52VcaKk9yRmgloYQJhjA/NHJRe6DzMIA0KKMu8RjBb0UySakok8oK
YSVCNB+fiVfT+e+7RIzFRUIkSKAhyqzDxfjRzVvfzlU36osuEIemMNBe+aJP
Z0OIse5F1V+9jt5RONaZGWKkYLNqiJrcLIjQlCvd9zdR4Kp/6rhKCgeKiUwj
QL0r0WAJGf1MjfCjTRgxilR5sP+S4k0oTEBsTV0BBHezsVGSwhPX/fqBVIMU
5kow+8nAX0t0iX6SoIHw9JankUZHt1dWZf0EBMtQEwLwOoxA8yV2gCbaVGgw
ZfDIMsBtjfO4wvIcjuee59+JCUx6cSJ7p0OVrybdNoTq8v/VWSftaiHvG66v
oNU0DzMwkOgblgN+JQJEPmhTexAP5iPAvQQXEst1CPDDKZ4uKzmpdqhqe34N
qXb3wqkhp+mcmZ4dVDHfILknRF7Wfpp9VbZS2eZST90lAc2L8uqQxprJb7FV
G3Zrp6CtoZNtvKjiQpcG4Fa57IV89sugg9o0Jra70sQJbc900o2/PBtZwtTm
htcJPu3Ngo47I+RAKvpeju2hX9bu/i2qUOQMzsvxwrAjTtnRa6/piOTc8EXY
qy1+AmHYwp85YLrlmBRYIb0EtxO/i9srhVAzkrd/IHWMrVj0zVPYMy4yoauT
LLYtWxrkFQNc89V+kQeH+zFlxZrANv1e0oURF0YOjI5ZrvEWMK7o/1B9cUKe
rezqetYraCQ5Zp4FvR5pOcOzqKxhEt34CRPlw4+M0vpsfhmpYY6tCbhJUetj
ppuLQDiO1VKGJrhDk0VyX2XJeAu3NuLW5zmGCba5YLHpEqIBElMBcaSAAxY4
S8QkVEBqjhReweZRT/MJERVZ3q3RTPA1He3k7mlLUtSn61shJ9FHYffqUs51
nVHmwtlXvHp7Ei12vy164SUUrHYcD/JOOyzDkL32m69PwOpgS3LuUd+M3U0p
svGFq7lBDSbWa0WwrAP2fhZLHUixSG1snoN4qpm58CKv9gpvOBpPqVPEhNNZ
dMU5pW7DMtCefNkBSS3zOOSneATrS3dTVefF3QB+NdKm+BgeSTIfExS8mV6f
WBl52I79CixTJXPLpOv+VWwpMZ29MPtijSrOlin+SXuYoOeB6NrLj2qT1ml2
gcdTfJGqgbGM4cXTjnEWQD0Dt6HjoYEICPeRmeSx59S4r0oNonSUl5lskRAK
9nFR1HQiYQ8E0yqhMbuWNTJC9xy0hxN7I5Eish8B+uQDXK/en7tm4r7ffKtK
QdmaYwm32ZkNZSbm2y/uw7NK2gjH3fQhv5TDsrxN9bcYEBW7E7mBeQeqBcib
nn/eXgBjY4JybwSqEXFG8kU4DXykS3cM01qEgvDm/Ydp65IHVQC0pYBum7jm
sar4O3jjV4iAvp4p2ha7dZrRAreniW/aCbKclOCRRULkuHpRzaENEo9eRS6I
YVuuf6+6AJWMPnLpqcud7YZdMcjrBLBkLFAhVMYri3SbgrBnlf7jUn2WFFQ6
sJkgA4aX93P+Nckp+JaOw64P98QnJLbgwYLluBlDRCeAmfvpV9jLJAmJOQ8x
l8oxRc/x4OT6JCxfdvuw32RWH6AzHQatwciwAS3nclu1+rhwEedCO4I7rDi8
dyuNeKXFGand4zNXLWB5eQSBtsmVFU5oKlAMO+++3LKx1xs4Eagpb8d7ioNL
hp6ouegpqD6XJ4MXz3Ikk8j0GHj/XBW65odgUH2h1lf8IbTWO27J1DhT9PNZ
aGc3JITB0DmWGqGMyOowbTvtR4FDzJo54gzwm3G23XPGny+Q5i2/7e033X3K
lmToQIuTPmm8VbvAsHDE9TJS3hhsFLOWDRKKoMZUtQeyqrZMhHTIwumzLBP3
Mk17yjzrMGENgMWZMVUI6VUNjdYguTCnr184lyfjBGzAvW/cuqatPk0Vh5D/
FIw6q0ICywbAa+/WS+VsvawC175kxoGCQ6Tm276db7vun3OXwmmSLkEDwiZ9
296zea8z8heK5crij4gDhfu1hr5ANA7soU4SG4BXPaxTvOZO27phq4FvwZ+m
tDJP1LGRXL2B8t1SY9rAmkAr6XG058eoWLLmWi3TRrUT0IW8n8fXbtT3i5O9
Nz6OTeiRYsiyavbc6NDROAp6kW9eDI75UB/u5qhoCTo/9RwUFR506jNkvYLJ
2vi8m0oMepiji33k8JfE+7XJLfuTTxto6QF8OoQ7gLYfbP+aq4voGykBL3eV
hWrhRnLyB2OSshVjmqp+YFZ7ENpMLX1C8tHt72QKM011qq9gBSnH4C0XCtkg
Cls1lHgTWVToJ1P/xkYPzkpsKULPyQXHU4fNX41GDxrLkoQ7qabT7YZlWXgF
ICROMIPxSZ9NwqJuT+mV7EJAT4ywEgK8jUvRLjttNBJn+QonAKP5RAxpej4W
Cn+Gip/sIQ8zu/Ygx5DbhfiRgSOuf0w3VhoKkJ3ir9nfiWpuhN4zgbXXpOfK
TqNS0K9G9fFc0VXsyo4w46/wW+KdcSyGLgmXYjdvR/wwNJfwUSgRQQBX+hV8
i4RrVSdojGeT8qap9uYNTjnkfdyg0J7uxr9H7vQhbNwSoazwTaEfzPv3dOdP
74itTARXSJJ2YZEC/w1DJGOTomntxlrjH3cA8uMWLkOF10c5anNkz6xmuRaW
H6pyV/NrJiJestjKF1j0AoMBRtyl2rGSL4GQmgF/stUxUgjvADO4l0FPKAHo
DO4me4YMB1cLGxBhW+PAF3O4/hkJ9Oc93m7JHX9jveXaBDzmZRu3N10dCpUT
iMHaqjpZ4DxejDKwVagVRp3eVIz0Zr3gOGF6+VwL8PTYaG91cEslLy3XSK5Q
wbnE0wwDyK5mIYjzOFnQiBKGULTWlh9GLuMI/Ntw+yiKmaRdTq6R8JU5Hbmn
ZUTKrrQDB4VbK/uIASzxu/xrer5EBwMnnOcjVpmeEG6LCGMlkr0QDFHdF5Ws
nBOJ8fjQhRFna5O23RyvniEnF4Khx5bn1dSg2LbAbNIQmus3Or3yKgfp8Ogr
NBH0fNGSDwvyXGdoA/ZkNQckZCk9lERi5TvWaziTyugDg/O44vpQVSZASNe0
Dlz99gfTaw4yCDBViqRrunRtGvZPWQqlk9W6PfQ1sZnTw6WYJeDj7TDKldwk
kHCDHylFDD7hXXvm8aBeSceZ7VmCF2z0AVaFRSIGqSAhTIhyQTsGFRAvhA6n
OaLLf3/QCVcufN3yqmDezEuzDddoUBEYk7g+rxez621O5p40I1xEOcGNCsTv
HJEUJ9PewKMBbCo03XFs6TyeCuEy75MHtLEJFjiwW2t6GEBpkH/nUP1qUgta
eXNQPv7812Ep5Z67g1Lq90jM3BIlix8jY63Yyl4jxFNnabtyNjrS4gCtEl/r
iQH+816rRWQY2T4K0bDOWrpBiGHhY1wRDD8evFOaL1rlPglgF5RuhQgfyZz7
G4XQRo+vWm6VQHFPM1KpxsROM4RJOv9xcuWEKQmSn0LFc9/glEupPxs33LZg
f+gVyVgWkLcqmQAUrDy/Oj8ilt5ho8ng3YfiNiHqpqNoKTPzTjo274SaEerY
kxKXOaYonP6AETVKR+ioBR2Hl2/F4tSXG5zFGEeOSiioYWQfVKCg46cWRbl6
cXRkC2dvLUf25jcLZfp9FSKug6RijlVBJ4JJNcwPYfyxg/qlOqdNeVKAAR4u
mmXBbyNbUtrzEhFWwsWrM3yybqEkR3UyrQpEYtiTIeR/oDmkLQSDLdaDb5MP
hexRjlJe0XPBWNNY19Qi1RxGqhnYyahS29ABMt2y4LEBbvlC0Nlr3B6WoRBV
etuqO+yh0J83G1oHQqNm59aQwgRARI0351I7jdlz4TsLtjwneym9CDpzAxBD
DSWK1lu2Gy3ukflbyq6vRGg4QfDhu+D6zoBnfmQTpzKYJLvGg/MNEjXqvriw
9FQWqyDDBayyb0SIgc6l1ad0C9ideXPC/Zjg3FFjXOJbmR+apxMe1TMKpNks
Lv/xz6eZ/gcjql/kW1+8RU24toEzYHRBO15H8ByQZYDhR5CMeYh9YcmAwK36
/merMjE0laC+N8Y9onIUgpQraj3DATlM5Xb6QKZGuFpj5voNUG5GMSxtXp01
7/G/DjnqamEIaX0YsX4+bNw9QP3TdjNIdkPBEbq91qjPtvo7zPWFsri/jAns
bSa96c4HFy4rqBOshjQ14auOd0mY6Iu/ou0qSNfjKSaYSqG+Ltdgcf/CHRFy
uWy4m5ZdhfbLAukkg2/nVwiMwbKPZLtDAuHZDTtigIJaXwWE6BobO3rAORBF
TIPxtmw5YeFvp2V86gGnMc6E+OyHlKiVnxe2BLevuSiw1+MvCKkK/g+FtZa6
Bf1A+P+0Ae3pGhz5XZSPAjovYC51XOCAcX6zo0DHwOyLUZiuLMF09hlPtyEV
L+EgILchcxyxm/4g/rhA7QybA29b0r+uMbubmL4MHxzYF5KDDejshKMnYQ1W
scdPL+tCT3ZBUtI0dm0Ho8Itxs/3HCI1+EYBkyfSJJafhvn5eDsWZNcJppkN
nvv1W3Yfh6DbFdTTt6NcK2fIhNgvETnqHO/MQRmKtvhswjmrL0oaRgBqgjN9
H8AL4YHcWJQCGgOV9KzQS/RXaXFnuANEjaYbaknGERvPSUFn/nXMh7q4dcqn
zPEo5Y5as389A30fcXMjwPqXiygSixOq+WTe25dpwZe1KDr5MhjMLjezD4Og
erEzvM/oX6L/Su7tbTEt+oNYQ1ausajJ4R7F5k6URTcqKC4btDINGH0yyEbl
1vXzmDJRMsRsBZ6f5FiYpXbg0vofGcC0JCQaUlyj2V5eXSB5of7E8ymjv6Vy
Yljv5B/mRaQ4hvNntuN1ezBYGhZQIgF9y99Mcu4EuNMS0jwWjraCmE7pBMCj
2YYPzj/eCuO9d1x8eMHN+my4fE/4FZ6cMdCBqxoikl1e5LpJNI3st8l80hRs
5K9mhwqzIblnUAcTG/GEO/WlLG07Z6jj3Lyc9Jsip8UzHnp7qmsOE7muE5D9
NiE3nHJu8/MyGETxg3qRGKnmL6pvE5x0F3kmoXLfQcuCCY/hffw3i3U/pnJo
8eK/DK57kFXVKns10wsCSUK3/a2XrMdFLVmh4Kgelpyq3fzpdZdrY1rfqEDe
bIdfJ4aWMg+Qp6DCGsvPrS+2o6sv6KZzj3XzEI6r51mzmDFVU+XGusbDQq0y
0E+LizTT7xZ56j5NxZjV0jDotA7jVYzTFSx+RWVXPKHaOg0kt7pGjceNmaPE
m2omj4WFQoFmdT2Cd6L3eMbOWn31Rg1ADy9vk11dSlyG8Y36/m2sDShl/CXP
Mm4OlXM28R4n5cj9GNxmbSKwBvgx1LvriGZsm3v/f+On2qflCYWPCCmH8D6h
hSIaK7JjecPxJ4ocRuLmCHxl0OWtYB9PiYg3UUdcubBsaz9mcm2gG3h7rFsF
BG4ALBq0T43EOm2NX8w1ukJTdVWhq0xZszWWREEykxYfLG9shMfpnhITJjdI
Z2J/FArywcybjFBHWl3lzlNkQThas2+kEyiyoGYHYtlcOgVmG9KilFXky0nM
oMTiBLO8P247iQE08oSxxHUhCYjC+W3YWlJwYZ9MpCG6ASRGpAS5WGUC2G4c
EeDlX/1W+WVpw24iGHWP1+ZunOkTf2DW+QbWjGY7stiA5yGMRvOC7WO/3cZQ
rQ8UfwAl6kJ/WyLYwC8R7Wk1Ufgk9qpE/QaljrvteHLj8grsItlU43vatu0Y
lz54fLN52ebQ5Ewq1jpEXV4cEvZRsD8Z84TMRP6y9ozvooxSQ29I8Zw6VQOq
+BLwvEN/F8TGQV8noOxNSklRMwfgdMpenwqEa+bPd2IpoA6LEUur7J1IcCzi
UjdXVuN4c3NbD8J7WzpptmJTHHvdxEBW1/9KS2vU02PPxjqo3g/dXZ3spOxp
x0z9tz7tffEG/er4lXN0MUUeKlDINY+HNQClT5m8+/Yji7vA7fdqJJ1qI1hn
Pkzhka47evkfoF91jnTtXoRhrBgitAwar7wUDoX0nGQFaYHxKHPbk6meVzRN
6UrMNDW9TO1tqeuM/CV+XAVmXTuuEAcikLh6VKCAb3YmsCOyTRVk3XyezNwe
FRZHq0nd0iSuzKVIWHh3Ux7pRAE8KsVoE6OnLs/FKS2syveE/6w6Ki81kz+m
i0eV8A+Hc+z37gVwutXxjA99E94QhK56JFWkxcbChqNZdNyV8uplJOo+Wzwj
QBkQf6/gbHSa1A7NxeNbrv4iRSkKPXv09kuiEKbffdFgtKght95l7JWjlA73
ndGTvMHbZWT72hwjam4LB+Kh30yjlB//cWuNgyn1Zx4kxqP7n6DyD3mTl53r
ivIMpAuQYZECmHhezf0LFYIy3kW9JmZjKISR+fqHSbTXVg3skN3/+/025AMd
H0aVUpbDb42ABS7ziZaRxYDFdA4jWntKIPkW7KDmogKDiHwaN9lDQAA8yaB5
SMClNw/pXwAffKJMYISQYxilMadzc0kPqxhE5qVoPBeQbCzVwBO16CPv0F8z
hZU+9Poa/zGRZNsE77kHljY4CJeVxNscjrJUhvZpo8S1w2AErRBIH+DI6MiN
LpIukrTRtXAScsbIGEIn7gDqBDsUq7MkoP6puD6NNojWirSmOH8HUatL/ddN
wvxYnlckwmY8a74KBVwVIxnAHcVCa102hQ8OAKBvtMszJBnZpMm/LU78aJK0
hzUZ3qH7mr5auvUr+xWu1q2X0tuaoK5xzYXvPQinWdqO/9unBznUIw6E8Jo8
+zdxAywS3tem6QHnPHcOglC11C4YP+VjIvOiT/Tj0vM2YtVOvsiGTp1iOGUf
VnKaaK+zQvPeQCA2Oz61/zssIthaWCb43jYUU54y8XlW8SMzB8wv4UKblHPE
k7/Clxt59sqcCrFALmgtCEMWX8eczJp++sO+xrckt/rTXXhZqeryYU0z4jjQ
9nd3zOT/QuJ7UUA8kQNTVIE2+DNGQGrEoAF+Jg6v+QlAcXZUwmw/H+GP5sZp
dTSP7947i3QAOgmo2uP62ohEhUgznv6ioTq+1McBYc4sKddviBc/+0CUaE5k
/H1eqSKgQuwdBk1RgROOA6l0euXectwd+0blxqv/i9tWycbncWJEUMHMjdwa
Imwa3MJvjMaQqlNmqblu/KzK9XVVM4l/kqy8s+pkNJPNdIQXFx6GvebhUa41
Y1nS3v8hZG6E7bYt/z8t3OB/Wl6pHGgMl6qY1Il+W8ExyV2COuo1OFYWvVuz
kPInrQgQBVlBG5Jgaqr2CA4t/mjfSo2a5Ix+5cBoSwxM0CWs4VA95YEXtZFb
bVn2U/DAYa8BoJBRukEz/4fkgt8+XBKFcvyxV6LDzTU4ZP4sNdEuW9MjAaZP
AbVsnU6luriu/ytLiIDl41xG2z02bqUrZBKQs5yO40LjiGblt7B/OruVQQ2P
zDfqvDn7aa+55cVHm/FqzWBkKcINP9aHIj6M0Ea8oLMasMQpcKa1s7QTQ5cK
G6MyDjEIvpA1y0BmetHnZDLrU8F1qDi7byTIzfpxdeurOPg6VEKV5eQs3VYh
bser8mpq9m6uBtZoiCneS/JDLqsLXPZ+K6PRkr8YjWdNHnNNXI8CsDxm6oKF
GJIdVy/PzCGf5lz4MKvaW4tgs9Qo+DaF41TD9lFGULHHVLIisx+FHgusbCFB
8YojM2zhdKdEhTaQgFjxNlABdjIqj8QWIKbT4BFmUyy3kWag2bxoTRUdE6Wq
WFRyU6cd+aPI1ZL8Cc0qngES3GN3a3STfmTaYCAy+wGzsooYuc9zN/LFXPn0
/iUndZpuUqHQI57JWyRjkfdBc7z6cK+zwuIykiMBFA+atrRtDimR0szp+ZwT
nbe17ySM5w89Yy7OFDMNjEED0e6kS/ApgLkh9Lj4mw0/gbxnvFMow8kpPDK5
FPqbE9f9hGkCiGhzcimzhMt6VqMSd1OkNm6DDUN1QTF6FHxsTSk1e5aznsPi
KOQ1Xa5jg9M/Xxc5FDrJbwYn5e8e7kGqUNb5seniTS6DrzVef79CeZKg/8fn
CLji9kw+sU7/pSkfgO0Y0zNEnZTxOXojEIszTk1Zrz5Uy1M140hI6gGiIxni
3jcUijzJ1KzBpWe77qdjjKpVEjANeP/4e9buR9sUVZSP0lgZwtjDos2U+nzy
WnnkgEf4s0mHJHIwX1+2T5dvtO93DhaNcR7zoyxIWF4+vJlXAn9jufElsmCY
b414NDrQ6+TdjClmI2NkPOiYSJ3sI+V4SOT4c5EPyW7C86N+HWVK22l9ouHw
II+o6VzY6EqPCZKjaOzsZUNqbmVIi2vNuVAAh4LvhXJcvA7fRbzCK2Gt7fRX
AwCl+dHIH9HgSTF+btpwm5FfFuEiHoOArDY/Fs8Jt5J77lycpY1L6rFPSa8m
MNhkYjRGIpU5w162incIjG5I8PkqtOnujIEfeDDgYzDOGjt7WQLpN5pLLHBp
Qv6Jwu0rMZmlLP4LPBl8yS+gOzDJYUVXQI4YrDN5Y9nu/0WzXhqZZtVoWMUX
WetR3NUtv29xiS8LZvIgfjWKjpnXEb1lloPt/1V1pPkM/5H0R2gNkEhzHWSr
yGUG+0GqqMbkvqJcv1LZB7VLb2Knc8WLtfFbxlQ5t7apd7ZeZ24USwcaFNWN
yIxrUw9FY7RloI5MRSFxj7St2KRK5hCkXmSPVrM84kjpElNczsiqLbfoK54/
Gh97GlLrlyuQo1VO8At/ceoTW+lhs2o4sVSQB6HR6GRNdpo7zus2YSHu9CvG
VIHSQFQpcLInNZPlLhIYiKhD4+C+BlFQYPK0BvN4x1i82ioW5NVU1iF57I8n
R+wq9/gjLsOiin1o1sqcjEUdaNtpTnupN/X0XLYdYzPUs+TarIy1xyIzvLRU
Cu838cQdgd+3Jfs+5xls08FYNRrMbFGHMFSftJ/qPs8lNTdpxSQNHJDVIYkQ
cZ5xoiSeH1uH9qgL9b1E/9gQbW1mvWESCrJDjQ7Czo7afFGDN1ThcWwe2kVH
5V0yq5sDc1Ie+EucQF7H1LaXn2OVaI8xSAn681lDgamcIjmOPVzPdLd3ILi7
pFqsy7GQrrMNIA6/N7QQB1OAxiApWzXzrezfrYcVPLl+wCbkwVm5QLR8Y0Q7
ZVc8omPpm0BGYRASmRoYJmo8kSnEfkr2QyW8zfopw4Nzv3UG0DVCpIMD8dqh
godkJ4gFqIbb+pPO44TEj7lI3Fjl4BEeXOMl2LQOTKbRT18DDQzFM16eODLM
BFfDf9YnNpVEcCRuQfH8amXoy19Yee5OWPWtR33DEGk2VPm89zCTCRpa1mSM
I7cDG1YcdrZ9dWnxDSbV4itsn5nA86YE+1evBSwGH4S7vAjWI6L/8hRZ7qk0
UAj0qC3+nVFNp1IyVbGyLWMaCv49bsm1f5soajsEBph+Qxc/5KoPV7iPK9LR
KbSi8nTSu1lJPzFCegBMq4vKD21ffVDgoJZMZocapBUSk/wgnHnlgZFq6uL+
wh2n3kzHBlNbOCGkMhzFcj18VCmLbm5toS9lDS/5f2xh+fvhH3wfDKE8CsT/
zvl3mcddbm/ItFtnSUXLUP5FBE0pI5lor3fJA3+P1YgKWam1Fruc0NZlx+15
oZKBOl65ker8AMicTij/0rTyWAVfPGPBxVTnGeq3n/fnnwvrEjhokeZoJ+bp
vLHKwZMs3WcSBKSGOO3w13r9FoGPJCBDTty40zKyA+D8umLOPtY9grb7dxav
z/BpApLkBHJ+ghReQ1CfTxHI+1UDdsUo+jh/kPXdVDtRkHOkBnje0UpdUQqQ
JTsD2XRTmM1dsK4N8GSOTqBfCdOXTfjetDkhK29OVkZa5OViBJxdXRCzEVil
kQCn0gsbP7vftG9+DjnL4RsPRy1b6cUKEJ9coDU0T1MEhlRConhQeM5GXdSB
Ipeku22U4Dlz+KVVB5u4zPdVlhO7hJ9K+tTzN9ZQqx+XUjfqmsBPLuGC5aL/
1vwqz40FARKJtFdIv5Ba7Irh636EKFPQd4ECy5DyOWgq5WIPWj5mJwm15CG8
3EKBM182V2Pct7uYUyBojL1pi0/0A88yHEilkEFBjcINfJ05Nv3MT16krOcA
ClLOeWG+bX6ILD1+dCBAezq0lWIMw3W/9puT0ERzZ64tl42VOjIe73/AheuL
9dea+nZ/UqrstNe7zdSp6xujMKLRxWssFYFM5/LrteVIZqSsismm4q+mOGMZ
ZiTnqBCvFYf68z5xL1lqOj2v+Et52XobgapwQs9LPRP3dfa+tJIREF7oFWNA
Kh9EnpGIUn8go/1+Vcq5a29jKQY3MpAukh2nYPWbC3hu8wtulZTXHPALyBcS
kBwyXJK2fobl0Bmibs31EPkAMbzH0VHctO74jzcsTmVv6mO6Ym66CEb/J9W4
JW0leJir7ZGP04JXZDT6DNoKmRaxPHXmmWCHpqsmAekfImHaXWl0oxA8JceU
9tkqU8b5GNWBSLRSGo3hDk5QDUNy8B+GLSFjzXfFRdjR0PNTnM8AZ7X4dExn
rtK6gBVleBXz9vPiEAfJnNVONN5ulAmiR4mrAXUoebmvj9ppvdXCjMCWNa4x
mmjXXign4bCnRpzX5UoYsCgtrsY1aic5BVAPb9Pct+U9gJqSogMS4P4/UcXC
WJtvGmDQUNvkorXCQqSgbD7lfo0uTEXECGkew/rQjSuBVuyIa4tiKwakTAiW
99zHNRJZEaqvL8noMyDrMleAsIQ+o07+QnO7BMje7wjLbJrab2B8xrUaRO/k
PYT6a+0JEypk+TrunPDvu9IUHuhz3bgX6v1frPkszuf0uCy/kJVDDELVlUQh
ntptJK4OKmGysJCFTumHVdanYIV43v8Vzze+cFPYp3IVOSOQ/JlDhMfFXzql
OxkWd5M9U6AzFHehSt5rvZA7q+X8l99WXsG0cKvS7qQYDAQa8GemUX7OEiwN
8ZRImdO5CKJ5GKf3vA20hGRmEEJQKEwNjyAGBa+6scnjCERBv0j8AgUYdo30
B2lsVmJLuNZpI8pN6mdjuiVJaabTVVO3c0B8mpEKXf+6R6Hrh3NzVB+7h7Hi
9ujePFxhE7PmQam80QWbdJ/yPOs4w35yUUpaHFlc7V1Pl0ETmaN0lmDPS0P6
Xp9v3eohd1HMM02fG/g6jWB5v552sxYFrJG1rsxeLs2vUiTq+qcpnT25tUqm
uX4LDUnbEXTFtpEg0sPSa1wn0qw3GXdWimy5M49b+lPgciLmnCzkYt/W45D0
IRvs85VibtvVJ59ko/w8uDYRiKRSeLXdP+a6W5uQEfeVAt+1P8X8mO78D+90
3e+gsfwojXWDXq0M07mYf2SxUYKyOjOhELXqtgpp+2C9NuKGKvRQYpZZ+LCR
HtiIJXnIctosU+YWQ4vZW3YFCIVlbN0D7p6WotZFQaACOLI4KfrgyhX7jF0r
3RVHZf8X24/SugrHqArGJgPRi+kOdWUKfbSlmjGh5Ad2ffoEw4Zwx3O6v+lE
aszfwVhv4uN5sskN2lYrEC8mngPNz3+m9/N5/Pqh9rs63XzUDUJKqmbSWR2e
ZKNC1y/J2bdGzKcN9MyO+1d0zhXHpLVE7x+TJUxLdSxZHI8e+wJ2nTcNTLor
PXwMMl8FhVCHMIxZrwGCROfDQv74jRr+NFudbxRF581CrsAPmW+ZS7KiEfTl
55vqtXdLn92ip9Tm10Bt0d+5oYfXecdEzAexHpCtwjH/FuRrwHC/F3K2XN35
Bbw1QlWISnqdv6To6Yy+uzD3H7QWfDe/xR6871QrskNGIVq3862p/ngllC1H
UIaKybmgat5yXuT+V7n0/qI42X/f09uzGtJB9p4g3yepkbTQN3FeCRBDHDvf
6jzBKPbiRwG6WrOGnRpgtmD30pUJyOzu+V3UASrLYhsrdPqNpJP32/H1KMEL
3j/bnCRGTU4EjmgH0XmECoiR50bcvS3HOydKZ8FL4/TKtHbNRjqddyHBWFe/
c1O1NfbXXhMME1rWL49IlE5fZy+313Rx3keIZznV01puw+O4WEvt/7uzOjzn
BSIG4lpTjLSd1PoCSPs1GP1xhUmKyDmx1NLDCMTd1Fn6sIqzaVviof/AP7Ow
h7K6hxeF/D6GxPweWd28iH/Z+vc9L+cuNJycVlFGSBsbBPNYCybNPHSelaRW
cdNeqUW6Hl28Qv4Zfc+1bgnILasshvqfqBE1no1Xsr502ikCEVlpMu9kYnEZ
ceqdBmNYYqaUoX8oKR/FNRg2jHnOtmrZmVLhqrZOToGNTLZXHVjOp4g5WcJ8
+4Vnx9qNDyXD1yQ/cEXbQgSLxy7XImIqojNGYK6pS7bE3teTfzt7B3R+ulj/
j96kGztPlFzpWsnUJ7g8/+qLJ4U+SgjAus+LeGgToeOkBw2XJ3USAf8J2L34
AqA1Ov2Gf2cSs9FtqKbZHzcnfwSRqr+s2BmqARt8Fvc+IhyqmHk5T2eE5wR6
06B6gppy5XZCfcqwwe8us0heIqX2V4YnpVlP1BTVriGG8MD10D1iC4uzIiEs
r+gwf4fGU9hMVHAWF1bj2Ayj9Pu4OSoD9DIzyrdNrPYD59o2BDxMt3w27bw1
PDEkdqTZYHphYsU7ys8EcANwnhmGabrXrRmoTuz/yGEy5H050O9bH1VCJYGA
VL0YZTU7VFPKBYutnbfl44sGBvHeIFfcbs2SkBJ8cRLlpKnDp3vyCUMiABng
ppx3SzDZj3Uh9XqdiiWTbqDQnQOgUl/uNfzd3pmZeIPHflol6Y/8yGwoqiHo
QUhOpEh1Twc1qE9UmXpSEeX1RrSEVs2BJVaVeXRPb1xjrt1Pxq022ceWUXTx
KfiusNyHxaAMMhtiklnyj22OF/D1aaQDmckEddQLhWaM6vWoAbT+gmWULDzb
5wBbVXrVslEj54vdOHbU4LZsIBxax/2dAH5hLFKA14Aa1TT/jXtssq8vI5E1
YVqjaprVPwWGf2v2ST1p+l+Ex8B2ikaBw9K54vV2zZ1cwY9MIX3toW9VCdXK
JpAbxkS6jM+AQwA592FRqjr3mg9mkyPBAE6baG3R7+rSHMmew/0QN2mOVs86
b4mFrsdKBILt66XqtjlOPOCddwLY5DLBSw+FUGAc7hQ9wqSwwX9TRwXRO+SY
MDQnBEw+UOy+shnsYC3E9V+G5k70n+hU2OjUhCq6yeg4zPpVq1RbOm5iu/Se
qiJZpycq0ZB5ldV5skawqPmOuMH7WFZXKpuduAGAHdlm/tk7n2Y6UcolPkw0
rThDzxSK4NGutCRI/9N3H7uu+O2UjUyH0IWCJfhnVD6uzoKDzXsXrPjPcgki
M3i579N9Lgi3ps6H83W0d8i5AYy2CQ1ehM+m3ReEsPLOz/sRS+yLX3vvBjUz
iMk3IAjfdCGUl74wkF9rm+UzxW+iKA9a7iAE4WWM2766ReuthHy3RIzQbqts
3TcT8m6BeHUmh30GwEbnUeqC4tT0UW2QHHOyHmh1037YJPzpojCP/fkpdwRS
Jkhz5OJBQy76DfG9qoRGwvPYCRkW95Lq65krBIDr7zVgvjeka1+415ZKZ/jB
BFs//DrbyUxFqBuJz/Txe0nC8UTEYKQfh6rT22aSSoghvlO+vkwzFhllqE1/
1rF807SvvcakowFjNzTFlG/SmN7Pcm0aARpBMP7ywLDZQjP9xCnSmg17NbGZ
ll+GpWhA1BAW28QZh0IbPBR2pbK0A3UbUfY79o4KrNXyjdvsZ7DhwtfExq0M
LTyNmYLCjXNzUk/kGyO/r2C7ez/r4Uhr9sv/yhh0Rce4kXmsBxdUSqK9DfKj
SQM3Dm2n5OTN4nE9xNbCrCVmCKjYYv1DhTSMdQhXQA90RphGNnyIWM2CJh4l
lTX484FXkt9mY0UTcfre4iA/efzVvWRWmnWglMF8tUXk6U7BJAHDlX30mQar
lG+FrsXuAf4I/dSqAILzy25kPMGuItmU92/n0MFIvKjjvQINfgXnbffTpRjd
HrVBVj0TWE28dioTbQMsRmVpuefNCv8Uwr8JsjAnZHboRc1xjHW+JXXCvKPh
BAlTivF0utq7P5LWIYpe3c0y5FUyXxKJ7fw7d7HUdPpQMgiB7rWFmaTZ1TZl
nGq7oLZkhpr3P0hqQG6A9hx0C/kk7yK8AJkga2+nZ44k8vmqJCtqG6RtsX4V
JkruknKaTMZhWaN4HXtuJnkRDsK3fKxgmEXtGvChtYhNdXR/214m3Pyl7Lj0
wtaU7FXkL00OHtJLOZKalcLFaq/CtHE4l1r155wbaB70I6x5CPUyhnJqhcm9
TAv5MCULHPkEweoG8Yn0rj63jRyEW0jX9FGTaJ+ThEPx2ya8tSPh1JUycbjy
TzsBJO5IOvkSL9QBSLBZ6/iDakMsoyZi45fSPGP24QhA8XUboRmwbzIM4yOC
CaVZgq5RKTbdnlFFW8byIqoV7jLCh2fsrq0z7TjXuTAekm6nsMz5ftFUVX6Q
2crYXfXmOR1pinizlwH4NCAbcHtYQ3Lc9sTVA2PurAF/s6tN1oAJW+zzWE/M
o8EFzFouBqxEi/Mv20iMsmr9ud3iIKGY4WPRNZaJW4QuRulug94k+O21PabD
Ct6mlQ9gCjT+ZJxCr6p9kIoghCcbsYTBOsqUUwjlfz2b1GCF+mEahwqzOz83
NKFvPrTd+bCie16cPAxLgBTXIX+l716UaeMmJRoZmTgb9rRcIgypa6UpVykU
reexXxKmqTXyUvx1fALMG5bSY61FtWuejoel+N/g5hfJjhJOc1o4lVeEtDPd
mgcHYIdPL9Dy4WImdYvpRvr3X2VUmvtcvFAkMh5ltDw1ZLUNGjAaFmsoc1VK
jGEMjIOJlDxw1WUiEHsqAHLBFIk5sKGOUI8up3wIgsFwDECMQ3ti1Nt9kQfy
gG/xUOPrMtv0uV8D18lUlpA6CrCAY6urhMpumb6sEKr25g7iTLbCxGHxGXdu
Jd9pnBShSJTKTwKGNWagNrmOkNHZfkukFXojHZBvfQHfzL8m5pTYAaMH/WiN
kAHgAkwgYnrcvD3We39qcZEGKQghuMkqhWuClUuIzHpTzEPnTmUmFoJh44ss
c4aztuQnKGx2As7ir3on2IOK/mKmhlO0G0UkFkgZNoB3G+vMgyrfp+MmGD/w
9bYC5b3Pgg9Du/drnysmluzxdHcc8bumP9PU8KM0qDCEizp6pEiPD9bIRYX/
XcYDmWOydu1uw22lt1wA5YmGRy0+ixhSidpMPuLWpKXq13FMQsadreB/36eN
CZPtR/CKuT/vspv/t308nFa006MrGpCNropc3GqDFzf9EM9jjiG5YXoRb5eN
0pN+QA0q1U0N/7EPiQvdemzSip63BPdla55BdA1xhl/YhwGxcdyyaNaKek6Q
YH5nLq+xvaXgM98QPDCSj9QXsjqrUWnvgvXgps+5eBehYBwPKBtY45k4+Wir
Uhk9vbRgAoFr7fLUz2tRQbilCc7fDyW9PE6crgNo8yoM14d2wJjczCyn+nnc
e+javXk7Nhpd/vb90zbDY+aiTg9Up4tbpRHclU7GXALuOy1wvPVUErpmT/Zw
I+iPM8IawRKcR0iP9QQyMWllQNiRD/Zpv/ZICAWgQEG4a0HGAPuOwsClKGF0
n/F8iYEHkEBET2t18k25NzbGrCjsH8cfXrPYPuZxGPCz5sSafqYV2bJHqnBj
Y9ZLUZwetZiT6KLIcY7hmOz0PsGqRL+6HGer

`pragma protect end_protected
