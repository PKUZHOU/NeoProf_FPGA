// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
o7cuasg8d99GJ/4E3RJIEM1n7XaqH1OTsJywHrUSntPIbm9Y8XD9l6hT7ZX7aaOx
V1iygs7ToghDM2Xg+OWsjBehxsfvp+hz9P7ULb9oa6OCDKe8fW7JskNohGrKQaJx
qFSqVKPkrosRDP6/mQrtYL5qRcsh7Y7/otYjYugxBSHS4n8m0e99tg==
//pragma protect end_key_block
//pragma protect digest_block
8Z/hi8pdYygdiTaCREO3YErtx/Y=
//pragma protect end_digest_block
//pragma protect data_block
sZAjr3dMXorl1Nswao6QN2b6fUIBo88AxODJK42dg7UcgvC1UVt1xrqTnZSwa4U9
K7NZUNJIfPaoGTGQXsWpVTpKD8caeIrOKVPqKs0CBBIqUTM2LQDSqQIgVm+0INeo
j1YOMGTQ0UZktthjD8TA+h0rTZP999KH2aX69DbckPJOgvr+DFM34TOqCBDa/byL
5jqXcYVoYYaE8zLsGDbTpYyXmQq7RJhrFDMTD2h1gd6HA/jtnUJ9N9uvDfFeHJpD
G+7IBHdQX067005ML39oj1TPbELViOdU6Pm8helFqbyQiRp20QQ8UjbuRafMCFp/
sG+kutaBhssrKm+IrOd5IDQ8Qm2IbAoB/SG+63T/cloUJvWWS92BK4gN7UVkgc4+
Lc1EVOVdyArLjqzQ2tzSDrX5K8R4EWlM/jMVhbLLHRIBrV3eJTloTm/k0fLXpvX2
mxMfttrr1xylqchf71ru8JibWWgGXbFUsQhgjKausZreyS5H1aVgtPEWTav1XAiS
vN+51bNSkTqKlbQIWdRgHRo6DVpsGdMJ1/Juii7utW6aGs8HDNTjaKOYk/p1fW+r
eXpqsoF12FyectVhdmK0beOLb2Jn1sniFKfx0G0h4eaqpNIvSFY6m/qKaCW+7Njf
Dl+6icQEVdhGIIfgiFhYF8Bxg/RnsZW8Ym/lCvI3LtKCzmbx1Gd2uvb78r4QDlTl
PHqMRiAKspmfAr+5luY5DAHiTeBciDBEY5FYfbgVq3Ot3wiDWRwCzQ5hlgChTct5
w3EuxZMmZiH7f60RvV2HkwlVzHmSloaD5uH9QnGKec0PkTFt+RJMP4vui/Omqh3E
rweITsGpiMc9QuCYTl/UpYYgAeoKjGWZjuNrbqnNq8Rh1/hV3TFPqBVTD3zLXNmk
AykdxhjgbicWB/n31KhU3gXgJEfSly382JP4XGi2+4Si0MnBB+AVLpqVUgf4toBl
cKgLX78Fl68919xUam6vcGD2zwB+2cQ30ty+rnhSFITe8WYCZs7XwsMjWFFhATyy
xiqkGu07GxULIrJXn6137Nfzr0aDVe4aLoOyC7NESuPY7K6b7BN3GeSbaW0qtAjA
T78vTsBq9qhHvuQx5jbyxLFKLQU76m3cWgvnhAjPSMty3V24donZZdYO5QFfyhaR
6O4Y+forAlKGJ6Hhgy9kL/ypM1CsDThtNTDywwWywS295EQbnAqQEyGLmTHm3pXw
3l+/XV3VKCeVZXh1FX1uKENfccuKMMCNI5tbqJS6DceqfIGIbBqTXfN5xFZPhemN
SrzV4GXC2PzYfiGXhEAqP6ARPMk+GaKDxKeIWE7lxzzr0oDE2+ewxajgE1wN7+4H
36jypqtGa/EkqdfiBQeh9/pTUQIF+9hriOAge4J0an/DJEDePB0i9QevCHj2BiZE
iQA5YweBZVFveMdUaQKcsvSJMtpXC+UXSnFM+TsC/oMMqxTb/QN3s580MBZ2Y7Ep
qdW5EcdbpM0Hcw9qZxEEMYAJSe+qbnAVY54MQFKPJURg7Wb7J0EONp6h8r2IFyWv
gfp07sdVLJcn0SXsVxxWksNwEFaY50hNKt6w+CjYIQ3vjptxF7n67kWTFF3p42lQ
/+LjwiMFmC/cSkGG8xDl6ZftrrZZJTy7JqwpFS7aMVjHWuVeCyLJkz7Doe3u5jMo
zV/wA1KuSR1WoOmNpYAw4rug4CsJOd66lgXOYe+6/HS1TMixH67J16TvHw1qORmW
nWsmhCRUauS4or+Gj4BBehLP75dGS9PIPRzMcNdQWO9oo1OrsRTRU/WHXRn5Yf/q
KNOSN2pX8BHjCGNQJklMdmqvNwyhz9hyM3zfDxqhWXdY0Hads8Rf5DxOtyBPFyMs

//pragma protect end_data_block
//pragma protect digest_block
LVQ+w9XKAjUEn8HK2pvXH9k6eok=
//pragma protect end_digest_block
//pragma protect end_protected
