// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
18MU8TfyoCcqf8HUdDSg2QnuyV58DLECUX7PizIjATrUmp8smtlMjAF2EHJV2Jt2qj2a8FRFHFL6
iQTjzUX76ZpTcUZLs0uyADE9DmkzaefOGwXbW/1JZpUgjWYc7bAIO8Y3PobHuhSR6w046k+VBmtU
1b3ItfTjw7R29ng9ZyPlu7yQMMa+fndnKGWeIQkpTloVpRUky4kUZdziUA71XjHb64QRshJrHSxK
bNrIR19stG2FQBJ47z6buquMF8Td7Pp4nVXNS18lEVn7xeW/tgwwqnZ2ETjv/SoxXREyf0noGzIe
riHR2Ie8fIjzY9wVCxeKAijJ+iMNQWo48Rl1lw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 20000)
uyofViejyaVE+9RmT5AFQPpXelZFOv9KXS3o8vwAMcE5OeNgzU/Dl1HhANPPgibQNgtr83o7P6/m
wYG7dYLKcxn/Ke/u4p4G8CeFMz5FNRLd+iHk/R+4sf49W62dM2Ana9JF/ndyFxPwMkYmvyqMeyQL
mGn3paD3grmF+wpRHDt7PrsGBazFkJvbruDoAPM++ulOFBXicICBD2HJmYULMvDY1AgIs4P0HKsi
M9EmMhDxXs6ZjBxu6EZ5KhLHSO1UpI0YOW0LcjW/7ZWmGkALcioaRpotVQeGr00oJ6UaWB/auA+s
jnl3SYBUSSTcyMFEK7tpXKAMElV6ogWl+CgNm/BcvmJAw8/I0HnZQYFltD8ljIs/3h7aPHSLQylI
aYVHMeSFJyDTvb+TJL3cxBCpprPR0OrteO4NJ7qqQ6eZAv9zrq2FpyubH/nIYModYKjfPbhE6ha+
uCgmHUh/l+voLmK1Gw3BIwUUf/Vw3FGhOxzwK5JCXJ+/sCJMbLi/FHBXkXfYZN/rpo7D37X1HXbe
gC5sxjZ8EDx4InxT41GIgH2sErZLwlMGzwY/G49oYSvrUjOOWLYm1Yw0XT8Z3NEgFsd6+czEBIdl
Y5dq2jLv8IShK9Hy3ruHfcTGtseDM/iO2gFmfUa00eLhgqWyHrMGyHQ+7m0xN/vt48KiCZ5NPJmL
e1X2L1LPdrDi3h5+nk0c1bJd3jKElpwCEONnvVDOJ/w13EsQUq41TowEYU9p/379nP9sxOlu7Xqq
iZpw/jZT4MG040zq60HU93V4/Y7s4YiZFb6EzKi0e75fnunQtOpq4ZH6yuYmoSpUODN/vDX9W534
42BHbdNs7Xcc7doXjSkY8LJ0UkfhdKScYPpCGXVzPtqZfcGvZzgdjm9/bQ6fPzGQlvnJ9w5qjomo
Dg/nhJSa9RJ038BCYw8tVvgqK523QQ98G5hbiLSAkBqLKHDhBuu+daRgfpOzMTD9HtBdEwpDPOZi
qTTOAw1pre5rOtyn9tbR59idFe1robUNoM51GRgI7zOCNJa2gzp7FBGK76nVzxjyTUmEMMdyFfPD
23cN/rxBVBTNntEqI4xN9CpGoXZzeYvjog2SAmhTuxLn65D/a6xedzjfl+up2P391Ol/EwYn4AsD
HmQzuAqdWAamNDmNWUSWlM/OK8fcwf9gLKyuN7z+VWPVD9v5AIW7RnVD1lR5cqPY7YbPjjB12+SW
wM4tRsYeZBDeliA36iqzuorzRMZHzRNcppwbxstp8XjFlNsfoN7/RiB6UMps4uQTTDqRudEQ1PVR
FfoCjinOPfGdCsbdzDtcqBmBrkXvLCMxPnWNPFPSKeyJdgecAuTDsVGUh1k6Has2vuXfMVZD6rka
Z8/GiCfhc2ND9JPJ1xexZvJzOqCYU+c8poueWq7VeOw3+hOviQx3A6Bbx25wzxc+MNa6EnhRrYj0
in4w0JkFjs/dunvuaCljvV4Z4eRexbI8bFU14NHin1dItG4tC3iuic3Ue6SZ67jo61390rA993Sd
IFJJpOn5YCcYg4qErfqVurlCZacdHKu8yGB4AdkAWW8km0KpT7NeoShs19GFUCv4NGgyF0D/rTKO
dnqWmCXagyV6XYjnv8Zb3TjjKQivr1lrxQJHYhg3FvzRiKmlFPkX17GEoqXz6df6zo0HIN7U2Bym
6wdzzYKTOJOKTjzAVd05yzNr4dTE6JUMyne67R2dtNhnW5E5EfiB8lt4s2QIEVbmmSB6fu8aIZ6b
xat2KLiy0ZWkOxj5WljMavJRYvGrAaTm4mYT0xPI3Vgl5OuxgHxxQQal614pXJa7BkVuH8ubRgR8
JENvxLo/j6qTohASO3bbihH99fFjl4TvJkHb9+zloyHX+uMGhAbhx7I4T1rDyn9o8bkYL+4RyKMh
25Gh/8DBWKDZUhQsFHWmBgCz/4UJr1eGSyvx8XFLIgDrqiBO3n4XttXTZKrILd0MF00TKm0BO9YM
AvUN0dhvcGBAccVbIK9BTFS1BytPs+Eo+0wOgv4I7aDRcZvqmpdUmm58Dq763A9FAI2MYNVIs8zi
59Cc14lE21a316MMxQG7LetrBgDaQNt9OFSYyttYEd8tCLUjp8ur8z0I1plju+++2q8mgtHBFuKh
m/9tSlwKKv9R3Htv68EF0P4qu69FaJsHTcz8qOiEWQcEd7UGk/S70nB+3N8DL6FeQpx6xNzjVptO
Zhhtg4BzfX8xmULLhYJORYyYC/E11G69NlAqft9NqWMpl3xJuan8v4D20uqqWiHlX6FPGI7PWb8q
c33Paa85l82ig+llS8qlfGggw88Rsm5KqcVc9UtzQkbuk1vQq9fPah6zJvPHmPGe9oydjoL8329Y
x/FW3W2RBmLEycHT8V8uQg8QWfASOWggeYWuUU5049MmmxggTEZszIAB7Hkh4fB5y7BwRdRYi4LW
azpyB40cXRQwU5mkQBEfUg9Hvla4JWjkKbQH7AB+8dsLzMVp/cbDqqKxH6YHDlgdD6cPGNQAAhuj
XNVIlx50JKJ4FeqoQvbea3fSb0jya/6FEcr+97xJvF0j6C0tV/92A32chKWP+4nXpzIybZ5zCVls
5T4Fz1+vykECiDC8dvLnvRi3cMI1QXiQ6AOiAAyo1Un3eu53/bBrK4u8R5MaAYsNapYvwV+jQKSo
WcRkoOvYdMmMbi/K+cc9kHLrnFlNwHgdqXiadRZk8SzonPgXFbG2jfedwS8rcDWNBeOrTe6fS7ry
4jT9+j/tXKwow/DNghFmCTKBedMBdYI2pqTtINZtJy1bsQDKnoGJwasWEqHMdSCXk+5wlHEoFAPz
yGOG228/u12JQ8/TydBHtusnETjIA9w6E3u5tXawv4BSnV8NLS8mCmsSbNHaZFz/owl7E+AXdQxH
iv8hqXwgRlIYLEan7DMeENvg2Ea4DdAMPb5A1Um71mVDW1aWaDyfIiWNfUEA0NMZ1sQgFbawH4GC
luiPK0ELQcLuWHp8N4kM3C4UdDaI243AUCngSDlxHWPxIHquAYpmyClcJN9E9TrtfzQx4i4ghyov
wEb5wZMuPnGjfUmfaFi4O8hxIpsMm/YoUEG3pqqlOwb6ofrTVrlgJEo/gpUlzUIITsKTTj2gk4oe
RCfgwOXslfeTHa9tEMciI0QmWJFuXHuKL3D5RjUVdkwEJ8ttOUn86/gniDdqxcaXhZHnCh+eVa9g
Ic9uP8bvc0Ody4l/hJ0I1wjR0cV/CgJCOL0jFJXxeAOcn9wE6T4qNPgLSYKOqt9rTEqL8LZ9JyBz
zMEBiYN9I/UnBF2TP7hZay0MgHxkbSwewN4UTTMH6bc9hngjZLwAa1yY/6S37k6YGujx0+nUszde
04IPGvlZgaLXURd95JrMlXRjAbJ/+E1G+vCd6zp+dDImMrePlq6ZCxtNvGTHYTg+BUIHqUOHdnH1
gUOdYDl9J4Q6NAIA+5fHIiSOWKBXw2VbWR8rT3f6sTq6nByO2JgwKoSyPrMnJcwquBNGX5EyocuV
sy0THq8B7mUqgc5dO0Uo406TRFU6hSHEca9dV2nvdoHB417FvVoyplxCLG0nCn9JeyJrpOk8pLBo
XZdUG3bh+aD2MYk/FMDOrAZeQnPAcUTIoghAJZBaS9B7gYd1IdvrHP7xuZ33kH3OKHzkd/oHSjg3
ha6E8nZHyPc58CQlaegcalOXYpx8XqxeBMunAmmw8ejjjXmg4V8fBmg5sp2oDQH1BLmloZ24ms8t
N5WNTu1mNQ79g17vA4YZ6BbtvJcT0/tUJ5C4SLtTiq9vfXn8LPTsx8L3vPWOQQwKoMF+WToSWDBo
25Gk7Gpxr6noQv56BJFeyM60r5G6mIaZAvwNu4r14r7z67ZQpxuAntMt5yfjDN/QL2Or1vFnUALQ
pj/leppoqW91xRl1LeLg4L5BxxZPq2ubKhuN0j+AEWGH+Sh/i5X6N+JkrETowWw9KNPn15e2KsWA
Q7LwPJ49iNAHGZe/9l0jE0Zpu+Jn++Lv+9WgFO2fhyNu1dyY8iiFg+R8s5uQUtBoQ5MzAV/eByuZ
4Hsn5er3hAiNppu3AGq/IHryiEnEYa8WZXZ1ognCQ5hS97dULPEOMdvQoyqQN63583M8fv1EU6p6
KuwhEiPi8NWMOiXYWRUCujCUPHTau1s8jSj206qqbi0o5j9BYtJT91Xdz4a/HvC89WdaxI1uRCbo
sLa4EAG5pQ2VCKXDr2ZDm57UZU8WzWdLrKsKS8Tj/qcd2duHMOGKjKwYFJio94KTQ3AZGLnLeIoo
BfL7KLAb8pad8KcK8IwOJrdbmWVpZPL9x7/dMtrFP14LSF0DrJeWBIQiadG2SrC8Sq3ZHmxq8uc+
W5YsAqQ0vZ6t5ct47HuhJC+FqkGW9m2212zbZlitEnnUPZy6W1sJleSC2UFFlJUoHcR8QDEboPlV
YIspPWUrzhsvMXneN5NZKj5KrOTauiP68qP1PMDzRmwlpjzN4wnmMiazU9nagb5K1iQIFyHfW52e
7idwvNLoiuvsBDRb1izgPwiGxdLMf4oSLOd6xtRLzNQh1TJ77ZZeqx9e9ZiA+B2G0IsEfELbGcx0
xgryamaLqTU8HTSzDGZZGLufaV4L3Cj079I7gBThPgXsSVUmzuUePMzQI1hpEVDY+d96anRLyMan
csrVe2aZBDvqRwHgiYtGlYMvftbkz3LyYCviB1miHDICOkstxP77jjYOjKh531/6OWPef+v4lAz8
1uGXheaV0pkPfXcbhVuHqHVaMT93RyLqk4yrR1gh5PX5TCYpB4EnRPIEF/40n4CDZ37B68TQaGCO
tsJZXbR9FmcPeUkK6rRyziM/t0B8HqEVRRmTCpBMGmMSBjrhmEy7CB7sFxrghl/zWx0iJke3fzik
I6Lma8rV8O/eh0ZXGeHBKGgmtNdHtnO0afSN9+R7/wwEn3U5mlmFjgnCsBIPJo4j1mbLSdSfwO8n
3KEFwKbIg/KgB8fp+2or9ZXD+2X/D4RAzbYKIV61MNIr+Oj5/ndDI63KyCj/uM++CXCnxRXaFzuC
44OxTXBJZxzZKurpm/9mfluyoK3SC0XXlrw8aXoEpmSiMBKw4O8xdkVMwpaIplYuUGe9FR3aeV78
/lrFAQhgQfZAkGRmCOPNnv2cs3nrvhQSdr9ZH6gwMMgeRttqI0O9ng+DvdwFWtWcKmF5mbn5YRUI
326jaX0RYIsYb8pcmj/5Up4RHjnrbEfYVg7GtH04qJJanWiCbT+PKYurdwCGRKUg2U5UA6lPrRhc
7ns+5QZCIIPKUfBo32yeK8nqRRupVkz/uge7J4hQFPiXjl4bN/xK9ZQXWWpHvceZj0WXENv5CIZf
oxfLSsuWjiHLJ2MgwQWFB35y/6SIUoEm+17SdZMRKZtNLqo8Qv+jfpky2QK/dET0hGYKWjx6vGeC
iVwukOzpfByQzkqjyNchgEOW5oOQ6I+yuanPqmTiHBcsgkPnApmklb9TOdmwsGBwbomMRT3n8aD1
OW3qMBnPlyI8ITjSAWhVIgdG2Miy9zGn4nt7idRKSZ8viHQwWxxnk6dZqZpCQTTniTtuZn8j5l6q
Vb9xZ40Orngko6eUDj4eOmmiiR8/pUikFzHWfqjVWNPop+hddHCZPbd2qlfQ9E7b2yx3k343WCYf
40YnkBbXFOBnCkvwQY/9IEmgL4FAO+Ty9peiUQrDcKRZqE0S98N2kKJ71wwd/4SJaCgEYVLOXa2J
w9i5gV5xTjtdEBJuRJZvJc+TldyBXmBHlLoEVPMFqV6dXYjDX6XQbFrhHEXVl1FYU3pWy99hBhzH
B9e5DY0nHEhq7rYD/jhc3OWSX+B9LHFx0QWAWM33gO9c/CPvZSL1acDrI5q9E2Pk2OhxTNsLY9Dv
9Mgfs3e/UtgMpUhkEHuht9gGPjU785uV4JiMLqB75J7DiXDNtqBDAxItJpytDdeg6sNhLudcBfhf
ck6IOgsv+rMLO+joEBWzbGsSR6DvHMv9iiD/qYIATQs4yDXznTOXOdycY+dSesNVvNCbWjEcAu+J
/rbaaa1ANZ++jwD3wqH6J6ICbys7DPunM+ee7XSAY3WjwdS35VU+BMSy//HRQZk06tttvrHsbJyR
DPzLmTYCQhI75WkKdO1EFcyLPkKWtX93ijVlKTBy6aanQw7mgoPG4/hmBOCJGxK7tp9rr0YhFj0n
s19rgVAH6xCjJ8GanrtqUdrMyYwusU6B9up9agAzwrIi8PUfBXBX4FP3W3fnGYDvmTgeK62rPUMm
znWnjXg0Wm+k1ms5GS6JV33lYsdUeCBdMzCHDOsasGnXpAJjj2U1mfNWW3VImvNxT3xRrfokx4NY
G0RgGlKmIiQlWjp9fm12qeFXoYkaydlWgl0Aojy1AaZrJ5qlfahHf6r2paZO0242nRuIjK+pWEuO
iLZvjK9h2ill77kGglso7h6JgTjzMAtD7B4wZP+SEs7XRMkV999hZ50V3nBk8doOdHLJ48UHLXC3
xlujtil7OtokR+BmkHRhdkyZhdQQ/+PQq27kNnSDFEtIFWVNTC7ckgLE3r1IBiSvVt/YuE02iwB8
EKxPzRi0JJLmfsUnpzuPXSFygaxYcdn54e2Mh1hZPYHwiFgAWX5gz5ul5c+kYhlfY9PPa9fYJTGJ
1cLkw1a/e4GxnlQ6V0iDclrEVW4g5ywo2naV+FAZTHwFhDzVkYDEO6V4wfYb0D0XjsFFLdUpk7qU
TD8Zf53Byp1iywHfe4m/1e/yAx/IzxntXeAI15UgJVi2/NqYobixdZLSUaDQdZo6CT4YVrBYR/SE
Jerfaf6yTxg5Ly5OA9C5+C6YySIux0MDgoYYb8QuQ8H/aYs8EN9eM7LetZSirEwdV3jMPcY/+GOM
PHzSpIba43C4ScFM99cuBMQS2PXgTwadBs10uu8YcLmIXdula2JjoSTEs3N05a27chRwjzTOgcEa
EkuuNtvrDaq/XxmyA9HOJDfW+T5VmjeczKNXAyx9SYsYRk4Kbpk2Ohl5MsleAl7ZehifVqETz4N/
tp+Kf5k+oxrqQKdnqewFcrurHOx5lDtY9cinicrGdXKgZfauL74+4Lwq+klovLsxPPhmJ/rzNLhp
dYnF49lNNwRKlU9r2qKPdQg02rc8Wna6jtlg2ScTeeDfNwIbwOw3eTXqk3MAeAY7lZfb3nkRLklE
EofZdoHkLbXDGa1lCUqV3D2YBquEMBWnuK5v92e5Bt3Lc74CL4+02WslfWdTKCQESv3MRXRJfJro
7vdoFrwTXy4lK+vZ13hCyq227yrKRFoaS3TcH3VwwHlx+NriXHlJ0LNcGWkdXIq8nRnWWfPfelM3
b1x4IYiSt/GnCiA7X2krAsg8U+KxufBCv8MOyGL17GXnDoPv+V37uOc2qQh4ONhYP+LAGoWeVjGs
P8pubu1PWnMbZvvZAPyrglvsAeQTNUUI6IVtjLdzNXDaUwEGhok2o3DMpUsbhJrsrz5/jyaHU01v
X8+mY3luWI6zswIBpM8wsl5/G/hAFMHfPrrid+pmzxFVhrAmXNr3FdGJsPVAUiF2G6IzKRyvrzlw
60jHPgQplnSUDQEoIIiYewhjaGmwjhyeDGch8HL+7797tL72KqGOqU7OgpCvBDONRuLAL9plup3v
2hu+QKkJBtpLIUSb9KEh1i7tqpbc+8vTDdNaPLvE/yRyqwubzOhyAPWOlI0CiMqxsAZA007D1gAj
HJ7RVemFpwPKqb8LS+ZGn2y1NjbIb4dgTgRuXanwHT644eZIKe/HpWJFgKLJjifBxwQCiQSi0OU+
VmgyjrVBgv/gLf9GvceUNzGLKE08nXz+6BiS1chHE4yjdGHVYaHVYhLcBureMbfrLqNb0HUKV4xp
nsplxcy5rntlVZBgnwB6DxcGxXNfwjuOXOZiQQqyuyp1xSkUP+ilHyPEYwEWd1BibTdCX1lRd7GM
t0bXYf5p/LxUHaYMirkQClNGp8zYau5wYyPUlw6/GjQIK8l6/vzRX/5CebN20h7y7S6fQ2aAHfum
4nE4tcz5U6uKZP+uTpIaKB972a4olYO1tKFbaxpJatT1ac0eOiAzHqn0yZH+/3LNRKWkTtA9YCaT
NpED2n6WFzg86cGMjw/LVYjuOJjCYSZfc1o+4Rg1cWQuYsYftXWUBI6ovzvzFbn/8fqaLMHNAMp2
3DjsATHW+eCgLsksr13yntJNCGtftEGGtuLKjC8QfEN3B0OeXr14BmSPcgSpX2w+hYQOuk+wY+tL
mZpDhrDs7QvPDeZfGPzzSRiirzPaWIVQsei1RNIIjLcdA5LI6F9GEW8M//1fn0ByBS5Qj32ov9LV
wMm1wsqb3yOFcjbuz7R68M3Wofbk23XGwsP2iiOIshvBykjkYND7NAkxIBq5+DlPKU+V8FVdQix4
ETtAbBooFU+c5BdVvIQWciySmlV8/VLItsPzq1lLHFoPn/eX0Eab4pBs5UtM/dMNKYHw9yFZdHTZ
ND+5YEI7uUpfu8kYKjfSGKeEDOj+eCqP1A/W7xyI8Hg1M8u/8XBunUJOIC3UXzpkD3M4DVeD88bm
Hu22axTM8zq1EjL34gf2ljcDvWP/tvsyiOKPgcZ8YBnHFrcRUZZM4HfKYp1IF1kSEl0f6vJamJDo
6JrhPhjrooe+WJetqZVOagVZu9iJW8RRpJfHH+X1WGAp3+K/t8zzO9+OiIVd3VJp/vX8pMkwpqRT
aGE1t/2DKYDSKVuo6yBmByk4jPTJ0Oo6Qf5+3UQ6ijvdfbkZBqwGATzYNYlovASxDFxgyHzQ6ZQK
bumXi4kdwYzko8oCshKyhzPHhM0tKQ/4joEmLn2MwL2b/FjOzAj0c2I9e+ae7luF0gM2CrJioO4w
scERqYZiUx6lhRL2gtuj60f7z9rGSet4pCYxUySfXZrwpOTt2iR3ACb8UeFyyVhjfCnfVEJiCo2V
Y2M2DQB9O+wIAvye80QhwSe/Y84I5vX9+LBd9ZZlu/vx4plrFHaeAMKX09CKw8AaFcGCqSZJvI3g
vnuiSRtlYmpfFiRop9HJYxasJIoIv2/byP8w9ILPK4EF/dAEwcUJZWSURHSto1cqiRGqBL80OnzF
KM2+K2kPSHMiOrS/ac+yAH5V5N8hIt1SIx/Cvk0++iIxr5ElcXeSOPOogDnNyOF5MlFtzQwE4Oqt
WDqoOYpeMirY3FQZ8D06NtUUhyDeodHWRAxiS8FLeHxE/AhHABJC7QBBHymevlKOTO9haRtMCDYK
aQ9kCWZthGdoo+2wLS69bzwz7o6KytCQNCMNH8Xf5g5Y67pANg+U5xnQ4juUDCUBzufy2OaIbJIa
iBj6cuc1NtxU9Oxrhi3HXer2LKRLZGRpBBtSVEgof66bexRI1W6Mpmwkt12iXBKsIejXHOuwdO1U
KQANU5JxRQ02MB3ibUHfPpPkho2/t4SLItwnCcQzWyK3f9NGTlQoNuJr9V6edwTESw2g25BzS6CL
GaqOsjJIEyGsEhh6H1WjQLk6U/i2HjxGtqsHQtl4VVwkuDWokgJTInBgAEXTMMIoEs0jvSLJ8FqA
SYL9e0ql/SN5iws91PezsUQbHbsUPCpiyeALo6nnRAfkNAlK6sW4aCmCFxuBzMxv0djsFN9O2SGo
+SHtaVjZd1+hF050bbojg/nVKsY6Ki12HXZL2pulyAdjjlVLOHybBJnYPQyKXHDeprXaCX4L1X0l
I2D2m5blguZdxehYVer0QWVABvBNb2glTx4mYL+0WFeHMNBjYZ95GEZj6GoT6Kc4ybt5htrk55aj
LhIjG/lSKwjxVKqyHQot04GZEJZkGeUk629WxvDxjY+wIyXv6LUkJDNCMIr5gXlnZ5WyYSm6X98m
l/MY/2YTqRAJmLCbi6g6SW6Iqj5LucIiFPv3+ufqtHAorlCmALaIXU+iG3s94xf8/ioFi8QXgDfF
pt+V/L+Z5jwggxj2faK114tXg+LL8q986mGncuCRoOr0ocI7smJ2qBLQX9mtrGFv4BgCyiIf2QT3
vIPrSJ7J37cGMEYL7hmIcU0JaB0uo6NyuKr650ZfymNdf8OUtoE+cHVIOSeWZ+5dB7wRWlKUWPU2
eQIsuJ5VIrDCwdj1WvOGza6307lY7+XzIPemj+hgPfBmgqgi8V6phYa5ittLAaWHa3Iq6GMGMNa9
XXcH+4U+YHBFlU8VSMAfjjRgXx5IsVWWy5K39SSzLqOetqEBhtP5GDy5tBtGfiu2sED/Hq2UFG4z
ao2ks+qre0jbWOyQqFo6XIXNIRsaOxjleujh/mxGmWesuAhyHDIXqRhDD5ZMMQgiC7I5Qpf0nX0d
c47zgDoWrukKH07zlbsC0qTQB8ZCYEkSJOKFDaglpgNgXLqqjCPO+9O+ZTki/uiiXNuIWI99ijUb
CCO+WOODb10cJCEmGn8+kXsgElMgL6RYUmWeJ0JvOK5dOUyQmpX9069f8GFXIdrQXFz9eFLvZrlO
ym72mm97Im0lXNJT/P1H+LhAMa6prweFk02pZaWKGB7ik0MKRW70I3iaEB3GP7rbgoQMkpUVfjSb
lFNdnI+QjygK9nllBgqz6QeaWosRGCAj5M5HXL2YsHfgJMpMJXaWU5eGZtUxwyZ5ZU81hIfs4P1n
vhwVar2pfHM2lKUHop8RmFvoPqYU/JcOp+t5q5uXSsi009AT66A+LXF0lDTGLpO7711fd1h5IqTc
ZYR1n+INz0mlYcp8sT6zh42E0skHtNx+q6xldXI5LNTfyCndOLgY71uOvyAYXJFKc6JCiCtbkHeO
erJAv7J07cNjb8naPcjhyUNKe4ZiGMoOT2DBo+S8vl2gUvdwbu92pX/uEVk6q0EBu9f5q8dLz/UP
oaO8NGbHTvO0FdgRXhABbEiHIbas2Kv0H7TwHlteLbN2OoMMCsO27Arb8tfsz2CoxqxHIzSqqWus
cluQrFmHTYuDtazluyN+33HC6QXSeAXWUi6xE8kC5jEZXoZx9ewppOviN9S7MeHj/SaYnSmvKwyD
Ze7AFB02txHcrJQgQebZXadiw8CMzs5vgiL7avKPK0wtE6aIOyTC2kNAgadI8g6m6pdMj6eGYVXM
M9ky7R4tcNCQubIhMVZrUcVDZcp+W4ERYIJX2QqV1YCnxE/FpcgcQ5yv8HQ604klmYHPz6ytuEAX
rhPGRSbkjo29T7+ncfJm9fq6Ux37dUu5WsyK7Bfgz9eZdKJKD//nLusybkrg4zhjWp9qpLmq8YfS
mFRLSOEdw0vIAQzX7IeUh3Y8Nd/Qa0RwkkKTQ+2iOXr1sY0U9sz+CRv6RE5YQ2eAkXg2yeOhcWWm
oVwkugCu57tbFJ/t05buFSm704p68r2Pmqye3Z5V1IiZ7ZkG8O3ydJgc1WL1h25ITmwBg/o8TiMl
PnDSpTLo5Zzf+z6AcIhimhk15lHr859Z9r+2zBwJqZOL0zPN5eJ4wA5tkyFK/ouLksSJpIg+DekA
mLUhefDSkte/iQ2bhgzTo+C85Cen9YsloGiER8asU8u0W1zDmffr7HLFxfzSObxMAwI54T+7CmJi
3512bHzJhLzIVMy72nvlzTr0y9u/wDTfYAiV69zT89AdETDtmEWXk66mm7FMrKUaiGKXuu0TWNDT
H9Tc0oCaJZI0DfvW71+uTzb8btEuvQ3b7ytCl/ijGx4b0+RghIFMcVVOoOouznEc4FKdqgJY+a44
E6dhcCbyXXqsvDKE8GoVDnVzLQ9zCM7wzROXwLSi8xltgHVcbgp6KD/96sH5UWmnek7bWcGa4Yvq
bz7pYvcLXLvm8kM7PodSQRoW10L2qqrHI9Ji9mDe3DrClHRMLR/ccxH25LdHRpzCmQiz+m01D/X4
VtRkRIUQHW4nPnCiC6ZURfiHFS/vnl00eWq7pxlLgBpNTLjZfhfgmeBIpH/zDW41FPe1z8zSe0Z5
oNGJG14GC4F534t/2HrlkrEBH1Zu7EvupcGEmJKMXMzPPbfiYC9qSg66QlvtxX5Ef8hLD97n8Scd
2TgsyPqMaK1mKhM8kIo2/9NjcEc6cRq3FdsU8TPAnbvLgd/u2kpoCrdgw2DCY9SGFlW3WoCoxCiE
6/US3+tJIsTLupjIbq55qoP3G7uzfGHdr0IOHX5xN9aonC3V8d9vZiLpPAXALOlDqUW3/GqJ9DSj
AlLG224VxBBVcUeeP0+c12hEQsDQBTL8XGCh6yLTloQn+U5zeUzO9YrYycikuV1j9Tx5x4ewgP2W
fX/+HfXBnNJ1kN7kfxPDehOChLgDjk/IfJr8+WCj7IQGPalVty9ax5vyzM3LO/jhrL8NfqI9tK2E
LwLb7O6Z0aOyeKoyQt6G10alwphNF8mepbElN6NMHUrbJlVtnm/AyXUcY0qPZyfor3PYDVnqHX18
Hgc7SYyrbiRE0RZ/dEIN8Hc3ntPzgJvf7gIBmHBQ0A6S6m9mxxKlbOHMHQ732PqffEaYZhQn2OJ9
qu6yXIbo0rlM82PZ6nSgYEnFwggzgs18qGNTdgblf/2HxkZ/hMfCmHVoJtYSU/OPfwKlYINGGPHa
mJEwV0xEOYFqCpUV8Gmmx/CC2YDyOwusGQ1UysRUsZInVM93oYXZGlZ6CEbJmw+grk3ivfDi3UnH
TQV88QDCwiJaTgyheJY0aaTo+JtZ11eua8WTXJ+SJd5ND15heiKvwDKRV0b0iOHJEr77NkTVsugs
OaRZk+g6FG9kdQpyeGs6RYDwKEKN3bxofSTcG1kco3qnpwL+FjA9TS3o9KU3FLbTLSwrFYVVa4xX
31WEtOa4W2qCM+DT9xB68KKrUPrZg+cPw/B1SS83LbzfHXJfS5PznEJnt0j3VdeuHrBFpTZU8U+7
wBglx0cAh3bTAybZynr4i9rwG4bvooYxO5LpWryUdMTRPIGNDUwzkm4PjVAzRhjsvFLNWwmJsB7g
09I87rBF9mE434tB5CrsrxBO9j/HDj3G7j87tiKu6in0oJr6Glz7lGxJd5gMQFpnb5LTjX+hIAbH
Hc5eusmGl+wbysNtEDg3P6Z+aorIo3rDNzG0DFgFLdPlvDbjRZKGMtS02x9hanRfVViwsU+vQmel
jADd1EZIf1snH2z/UvO0J0FMMeOXsUuRKovQdRhOAaazWSEftEHgoFPbDRsJfemeWw1e5uWYjqZm
DMNVcoypsjznEYQPMjm0cKfqekF0A4qWPGJ19sPL6kKdfr9h+iZepxZLztnczFT1P/WdaJ/f07cE
BO2XfLQUfCdaE/iOMCyKcO5ioqfnbCXZqkRg+R8Q8W67nGCFC+RiaDlgNuborD+uU3AO5Bxw9nLx
Cj1UB53GrRjlZjBx4TnWpnWWFf1t0x5EB5cCGKkvi+7ABbiVtk491T83dF4bCW6JiOs8iveXB5JN
hapmsLdLDyMM2YHbixUIBDSvC9CnxdYW1S2+2nUYWzOuIiT4yOhfNJ7Sf9uyJ2hvEgJxBzP7KSGD
UvP5GPsRMNU6UyyCBGLU2dJ14lsfqMQTw5UuY2YoHSW33RTY5GZA+NUhgtlwi/43cQ0Nqdl5U9QT
m4JcjHH4FysAwUf6QKIv4bu9Pe8CdYkKhQzXnndPOGqhI87HsTua0YnHT7/55lNzFBqr4FD0t4Gm
4dR3xGgVLY302w3lcG4fLZN6Tc0uQCJBWDOHmjetSC6RfMvHDWmUdLApjvo9uFYCj2rG3CvauDfE
jod00FRzApMW8Kyg2RXxQk87ytWBsRt9QYsDrNEWOX9XiRD7S1w5Fy1zPhhEuJ5GvcmrSTjCvOOt
74kfA6TYiiXXd9LNlq8U+FNhgqPDH0ZTp/ks2M7DLJZRbqGHDpfRio3+eOZMZj7Sm/v75egdDZhe
orfIdNnyCgapKeEdcQynkMUnYw+xx+jo7FA+7QmCL5S6TN0Rmfp6N9BwsRFYvKEPFmG9CKMBSyEY
MQm4xAnajC3kpraI4KNbQOJx5ObHUzObqRyA+bf0iMB+2sR1sbZg0qJJ9d+EmHpW57w6NnLA8Ggd
kygeEa4sQ7Ra/gm47qfS4lOeAClBJ/MdXPoyD7rvbjm/mFkBL/7k/1p8eGuMzd7XWSw9D41/j+kO
A6Tj4TGp8nmW/+zZcjyQEyQNyXMA71pM0gOizQDQKXIDjf/5cCFD3HAh7Dht4GgSVicwowXfxIxG
MWBOqVqXYt9WtJpVHw+oAeKlbO0G6l2VY/vDV+HZPUtyTFv2Os2us1iCim6DPMvuiPqqA3cQkjg8
VSAxGlUKMfSRbfp/e42JuTCRJa1gqkjW26oAkbD8KoP/RQPq2fBGt3lK6niAEiK/ptjNNo/Hjsxt
vz6Ym3Jmp3jkfWAOE0IbBhD1MZ2AOwadJTF6GOFJ2+Vxz5wvxZlf62dzVr40f2SHPvNhji5ZHCPl
WUdKlZ7R4k2vkn+uTQK4WlCoZGolqMjbaiDAcI8O29rA+X3eKDsWNWQHvWQ/ssNMZL0pyt3oaauM
u8jYW15kXhBpq0FqsqOgDp9JW9p+qSdQ9UQIzGj0oZqjQg3TFe/u7CfgQanuaU3LLqKK5NIHcFV9
ByUovs4A8XOkBxBfFNCe5eq7Pz644GKNLunXGHx6C9l4zlOErysSxhpCnDHoJ7VZSjjUoab3SzJT
ayZkAPqgCtxmBjFCOpac+H+Xe9qIlp1Fd65Pap8uTAs2mozrpj8SeBxKFogDQZTLPoFb5ZbhtkMC
G+EWdKzNAOlmDhRFed12TUW2OPGX9GBcVgE8tkk0qHz0Lia8gNwmwcbz5Qhc4t/eTd7Nl3SwVzIw
Or/Ht2lafoT//rjRrFjQrc+W9z2cC4xRPvNGd9PLJFdFIwJZVR0TZBsFk6DcIfNWqdvqHm4TXUoZ
YK1wyhQWI5+pTYwORBI83w5UlNBR7vq+xZgAlXxj0KQ0UmFcBTki5MLQtRpm8M5ZHq8N2zprfIpO
ge/LMS3NH+DQzaC/kmFaiTEZJ/0tdWdejADv94dSzagAtcpDP1NnfQcaBDYUErcp553mytg5L2yZ
zik9kPtH8oISy5QQu8dHTjUsXl2fpSg+DwVTsshPHFKC0YIh3juak80O1b1unw+hj3yw/PBtu6Gy
li/XlPHzH7xNido/xel/MiTqeQH9A1fRKOvjUhjJH7eild5NvzFoxm0WUJrQDXUmLc+Ri6bDlyFu
rUMlAtEbRMhfcIz7dfUp/8eN7gHvE3FtkClWb6rxXwrbfwbJ0PN49Nn2CMIddsNZSO7mUXLt4ppS
UJXgD4HnYOvFCTN/9jORESSK4o1sdNczSrGF6V9e/2mdpHOCIfg7bowsC4HCWkt9cHBqjwII3e53
+0S2eVB9ug4rYo5Zw/KO4wNr5N+roQXqFhoFpdcfv7QrJPrKb+LaM/NhFz0TOP38elnE90GFPmzp
aJse4dWb9brcoAI8zln2oBLbfGFSdXqJmFPYgaa7tb8rbdRVKSzprDxfZNC1V7bAEBi6LyM/UfUR
8DWy7TUBgVm12JKZ+6oFD4lG4Tk+o4m3eOLi4wNrrhYxDQHfdS+OYeM/3967jMcVm/Jcj+RhN83e
hGehLI4WXJlrA5HZylpxVk0peCsOkPOk6jWdIG/LdaVE7Iw3r7s7huK9lWfG7+7icV+/5DHCicf2
oENG5z3kZ6D3TzNrJer9GwOfQ2wyGQnHFY6PLA9eLc7lP0y3bTsEmJIbQ+or3rCH4JIHnDa5Ok/6
4ir2dlfp/C4V45KNLZ/0a58zFQemCPeFQk9ji+xHcDb47/kai4ya0QpXRfWJv2O3Xjd89ieXfltf
wR31M951hFE24knjGx1Z+cvirXkIWMAARXic73kAKNoYCYV2snuQEVMNlI8Vf6n+tQ3W9sFUA+g1
7QzRMoQu2YtX8QLuVwIBQRcdPzbdPr4kEystvkB9uVI9rTNPEnwiIL00DyZ97XoceQl49UN0D916
IM1VCDahTlx6jT6RbHmBE43Dz05GA+ZqQ+SczgfYVxy11f+VvpUpP8NjkcAyUnBTWQyZ3Nv1tUaY
HpYNk78IzKAiq9zOKUaIZQ12Nvcs5L17wV4EJpBrKI1ebo239Neh2MWcn0P5pWgbPdUzvl9xqJT7
ZjxonLBFyM9HqBJ1YYQoPX3Pga4XeDl8d3IEj35nxl7U39d2AQ5Aur0az6TtuE/10yoEODdChXd5
eT3lzGvx1Kt42J5joBOrNnCP9tnLyHcUNezzQ4pBlDRHcDCTFKZkpFN9EHc0BXWhWuH/X5Zs5OEa
uZcLLnm3aeQoejT+V2J86mFt0dEGeunGkjYyYaqtxiUXIfXbXwlIzWokAgTPjZNOp2DjIuOYiaQG
dDa3+y+nCdK5zg1UOFEk/hhqrTBeburZuu6ecwoLA+q+WfBMjqCAvfLQaoSUgAi/O+BBMjIatQgF
dgtadiK+6CuYPxMv6jn7gClP5dv/JGtjhiVGtiBp+gUGqIVY14CJBXmumHXfaNQO27ssowropPBt
KOT4Zmm7NArhjORauBATDaALAQnC7BIJHCYehvO0ThFA2t1+mOIKOZEOY2dXwiA8KGthWfgCpq1p
X2DF49XYxIroaxudNskRgTu1/io0EJdI35LqYW/BJZhJ8htRvIuLjHX3wS2+Ra/VOTrbjPkCrxXN
vw68d9pgPnU29e/G2+oYqZ2chGbwLsr9TAU0s398qsu+S5P0oDcDfv0XCAxax5t+jC/ngwYOlbSS
R22kSg1/RqxZdoVFird36AuHMPwm8rMkzIXP3VRNMU8FJRPWSRNG91pM5vTjCmbAbETJHcApVDOz
cB1SrZMMCeOCuW9t/htYCxIB/c0Fem0bf3LzQR1llYJO1ZjgpRGq6FrWQVwGlCfNmKMF970ZKBBE
tPus93HOQgwj3De2anZajMQrphoo25h/xejHy0cJYonLEGjtgbpG+KsDTNi2nDoEoiG5Q5H6dgoh
SDuuaSWvRSOTrsvp6hNBxaHWTRyftiz8FZEp7LUgAaadOw9FrFZoVZ6AoE8IpuFfrJEb825g0/sP
XzKQ01Hqe7A1UoylY/v0V975TJ9pxzlK+FepS43C6WHqug54h91+eB6BCIn3UsNFxDrSBvK+zTPy
qFZad1PEpk2/aSINJajatJ9nZWMuBQ+esjznEvpt2M7uZFVmKGL0Ste/otvjswRQo3UBOEwKG2ty
Tcy2oP0np57PT4tzpPJVqUCY78zFk9fHkyozfVNGH5y2I6ndLDRarPRExfvA6mMepd8E0gqJ9bfu
8lDQTI+0cCB6LTEVcbVThzj28r0ah8mY4bHywa6gY1UVqvwiNpLKSAerzmfw+ZJhLBkG+zQ4qsTc
tj5jyDApLf2mMlrmcEXiw0sFC14hvIpPbunZgN88KsqQSUD51xTQeYMHauiBfBwObwfE7NmUvgAw
fkbMNtyKv5W+srRgsdI7NnzyNMIL2ePXU4cBER+2z8kmXhyjlNbOU/RynWHUM1SdIFI5wIo/+6FR
i6Zobq0YbLt0VlU7Ff43zV0CE0CkwS+SnkSrtkiLHEkfbxaq+3+erLp3Qm5rraNd4lUPthofLBsz
ijAprmksdM1bXsD/6lO4uUnQbfdGbCbQJggva4D77ZiuIxUIiNwNGrJ+B9Vmr2arc1v95iaSI4zX
kK5I7TI/X/HiazbNK2ug4k2blFXLE2Z+47x3eCb7YVaRh0LrtNx+ukt26X2phXrm0DUWcCuvuVg1
TX9b4Gacsl+fSsZlVCptKEa4BezziOhV4faOCoGipcuCOr4W6gnKPvCyBRHunUSQd5Ddh/oSszVi
yyCrbJvm/DWBC9bj0F4bpMsPGTJZM9/jRnt1mxIB8mgLt/gZMBl4pwdIXotbrD9RWHuI4TGtUdIj
T+H0b6qPuuesLXIMxL61AphEAaEzNKfkFGAzTwjGGpV8XhwkOJVB7X1VWxtwRffQIK3X/+Bu3Xc1
SkG7b430L34JFZ5zJjy+dkVtbRHWTz+9cjhOVnkpYHlZR8o1cvWLoZelPPgu+2hy9Cfugh7h4S3c
kuK/1NYDdisw1ANtnw66IlUwqPuNEcU0TwdyXl2boRA2A+sGTf+DPE9nESCa165Sfe2NvvMOkST5
otbGcebVl+zd8Lms8OxuTXGo2SIAp/0LCuEIpgd02vZtMnLQtTmfV/QRucpdugkB6s0jvO7u2TRc
wKaaipvs7lrBNVjdYcgB/QKwSecBYWQRa+41EuXjkukontvhN5PvvvggyHNzV2owNry4fUVKyMvV
totm7CF8QdnFrxW4Bt53d82bAXIMtq8zci5UWkdHcUP8axkkvdwfYt1FtbGLK5Mjz4o/LgqvG975
e0vVmv9qDtkOrHy3FMG9VTJ5nomyRzLZAlZ4NT/9Gpc/OOWCWcG+tbD354HMS/0bEL+bZamUOFmQ
AzTp5931BwjjKEpV4W65nTwf4DZCIRq3FZRC1SNhyr+GcIj+dWGcrp0w54RPLV697IGstB76fgze
zPdy8YxPDgMpmR8GWkqQTY1oOKDfYY+WTu6+oA4WoIfT9uXHfTT9giZMmMAaEdG5EvNl3UeSalBr
e9vqejPQ8lmGPan1KquQwi0IOGnIpRNGlL19tcwn0n2oAs9GaSy+KhqEYZzJAmT/i1gcICCSska7
KEyJn1g1fr30kilUA77h2u6QFlqfyJbIAv/9gbhrAWdMdFatrd0rwxUcJesC8PtzdoS5T+6Eb2Ht
quSZc5XGDrphKUquMTlLqEg53GfM2fZOx1/Z1HJqz7TyElWLTJYFpY2YSj/cvs06ZlqmMY5j5cxV
Nl3Erp3xnQZzxwjv7IqFnbzn/E+9CYR3hZodQ7rHq3xqUW+31FpSBKVjnq14PM0MEBUI4ld3YI8x
vo/WvHGBNkeyEgQ6lLNzMQzf/ofkwzELJYcoUHoOfpEMuJJcp7Pg+yboiNvFUjATLhp2HR6evl6P
u3X2dTCH82/unaxW00q5JWfJgQXnjLZarABX/KfuXJzNzfidf6yH9vIMHCdorMpfFq3SjpKtRTez
nWpL848n9k89J+MVMItoDk0KCaBd5YcQEDrVUHPIcsNdezm+YloIWQO+QFI3irsR4YHyx9wPTtXW
fuI37h14nN2F7/hIOEOJM/rcUxns1X2L504zAQvtPm7n8FJe4y8WB3WAAvCY72vhhmxJimQ4yNye
oAVy1PpzutEfLMVbZi8kDdTJAoFNQXsgrxHBw8mvTAekO/PEzuohm3qF4V+z+4l06XTcX7V+vP+C
ZnawqycF6+0J/uIBsSoSXww1H/KGJ8Pv6KVysw0/U8R6V3yneOPUfSYuT8J9EnsqPJKBIMw4LCX+
Nt2zO6MgYu9+ZIYNWsb/gbMM0WOIzpGKjL0s9NF0Xp3krZPVbclEWjE1lh7u6ZHNzH5m+2DdHu4l
yhO1y9DBC0Goa6vkKUaFc+L0t4rl8cJdj6LDZjZSzWXS2uPjF8UJN3k6akcv98sI9dUhLwvDhqp2
NT4AQury1sEJVA1MjZATqvDfyV/IIJi4JCSpluUxpaxeNW6L++XAWMqIV59CmzarP1+pRNxZTgqm
2hatNWFekJcC1DkCb4suYGALOf8KHOmpZoA7w9CNB4YcZclfXFjoE7YsjLAvwi30TTdFo1gBTKlJ
ci4b6DwkQ7cEBmR39fQOB5BRRxcr4SWPIzuMIHFQlSLJhVZT9oLS3uVeVKHmcay7sY7rfeCYs8Xw
J+EPMO6WB3hrFbcVlLGdVGyVJ/IJFvA0rsABaY4uejVdEZazKTuiQP1oMwm8XRPIu9HYGdNSDceu
350ExXg01uuSDJUdJ2XEmPORTdY5az2SVg9TjWqRnNs2ixo0leWf0n6bBEeDr8h+RPzxv3ne2wZH
w6bU110rZAmpoa1PFTA2SH/nDS9uma0UjfTqWoCCkhvf6bEXRpy9VsoXan6jARQvRS4gZqVLGCYP
2hY5WLTEnOI7e2rQuUVJoTksR1UR25MN5ZfTInwbfvie0lWk1ygZ4FbPPA61o3BXNqHy2rabcH6A
X8Zm5KatV/UKBAJlykqN1qG89AfvTN5m9WuUCv1ZlQV0u4YZhuVGvQj6DuXUfvT7zT4YuKTweOeJ
+eEL9OhQB885DK3VnINBgzJlrec8ueYPiXtjWQdTP1LPEdsNEF8cQOez6OCQOdbPGO4BZqvo++t2
guMeFNx3RJVIBZPxfOHCX9FJwofiGBhzlsxGifXHdHkov+g1r1yZX7db4OX6u0DHK7NnBu2bVOR9
ffZSwHpWv74vF6FHNkTAUIo9XHMhug4GwCbZdR8kXjKEMmGuhOb8MKIct7UzQEj46b4wALN4DvZP
3id8Nkw2vsEUGnDx+M2IyIzOmiGSgleGaSxFpq3FBQqCHmZ3obOx/xTKYF/vegjWM3jFtjEGe+ov
tWMtgd5lvuv06Nmm9J+b+U3E5AVPo+xgRVM/2xQgkGyYJOpJZHxBuoRgMI1ioEdvTB1/YWUrOa3F
qKQxWT8LInGF4Rb9jYOBcoYBIojH2orT3RBYHK66WA79gpnpUQLr8JzPAbOIFJ6VT7sDxVIEHW38
LnJ1u5ZM3nM96S8ubm3xVamB3HOz+oPGxcvERKlFlzHalCuvxb/OAm8jK3WKEstT89sAiLJNIGRV
n3HQSg9isvY9fBMV9VuEoFt9GZC5Z//vsUdtmLCW85sjJ1bkq/tBWKhf3KOwSW6KaYkfU2guaeHp
xdOE4p34pUPh+b900vBjT+LrnIHA3G0NqJBGGlPNfE/rYJ03UuBecrngFYaaNnr+aK9eBnsRcZYH
ofrTsmCYUV/aTerQ6SsAzQQFLjuv5Z3kxRZDuc03U+BQPTay4SlxJojV6lNKGK/vwnfkttZ4UPRz
AY9g6T6PSZI2ZCYENcgHUYZzEro8mFQ7zgc3QADsJjd2/SUHbBdxEd37G/ad/SObNnv7IwQi5b2f
tbo2wyb+dtK2owq8igbLiNBTXY7J/T050/eBNAgpYTZ3Ai7PIvg/xjwFZE3zMvZ82SYTP6v0hDEg
sqvtLkY1aB14rJolh0fViJp8rrvuCrKpyv+PFa+udKVxTfWtXuDxHGizXeW7Vg76nZZbL0c0YaX9
ahObfPN/9P3KUSsUmSZUtuHhlMT0zq68V1K9zGLzEp1NZNBz5zlNxh0eguMUi1m7jP13xulrphf8
H9JwZLgGfiHZfddikK1lE1EGqePxkusInr4GEUh9puz8NwkcHxyEOh5B99OPTUHUqAzuZHFqiI8U
4ZrzhCMju7ywRdlnhnVQzy+R/b8JqCUaxlTkm7/cJE4WzVqIUSzB7ayQ8rY6UOwXp3ku4Dw39cas
amMiYcmn7Wp1W6KzPT+x3UUtpqa1Y9i98smS2J0XcShTPda11JuWuZtwUu/9OP8bqyiA2y8WFgqC
WkKKpu+PxuWCLYwhSCc+SVVIWKHde1Bgei1Jck05O3WX1PO2H80JDBlRH4rt1FuifeWvTlEQ5VEI
lgr1ldjJAUW3jO7vfx2EdI6wyb5dyz77nn9rX4f2JJzHtXVr+ODV7NUOhkkIsVsTNopLoJtI8db0
WDbP9CDHAiLNpbMvFuGeWd7n0fgYT3GFitWaAIJClOYHqA9T2cbR1MSGjvfT0FRIJNqvwNta1Vj+
DxLNaOZak27uO1JxPwxCuOdGdyRGqA1j+gJvDX99TXksqXCqNsXLuC7G+hcqM5ODAoKWRd4YCT5+
RIiWQhcVv+/Gawtx/oXmviuI/MIpuREKd8y3G711ioxWt8A+Ceg7x5/sooyidUUvYQGlif3tV1Ad
rmMxYLcfuFj4s5fUBKcEG4YFdmVonIfvNI3aoAwpYOsDlzIROEdjA6hEAwGaXx4oVjkBdpZ9w2WE
GaqkyUcM3EmKl4nquoq4jCsvWgdxrvEdTnKhXc2F/J/jGGr1p5YQt6dtL83kksmfk6Iee3u6IgEv
xVP80AjEvFfxYPhJMqWocDewHEzaX8P69ECS+PWdUlz2vshfHGB0LDluCtFkkiqIK0FXkmobsw1V
nPMjQbozGGIqhADfGiF+uU4X00kT93IoDFTiflQ8XzlGezlz8DG02yMNp3zUN9YpJsnVkPioqlnX
wJv00loqxb6y5pPY7bcDK1FhqkmL2tdlh6vpsZ9rN7Ej9imC2RhdSg4J3Kc5KCxjB9VIEqgc7Fl8
W5OwrMxXKY6Vkk/xSHyKTdcN3b1Oh4nFxbD/rmEOtBbQsi4C0i0RKvrXWTVvKUzcIWV3ocyU6EtJ
yVqPB/XzDq+hDQ+ZG6whiRvjyXqp3q0Re7PpwJhwvDlBCMioeybRwTYUyAqme8DZYHFmH5di8MBE
iGSM2HLstBSiFZnFua2TAVmohn40a6SKp4nz/8PN8cHG+/buPc56An+THkvxNKfhZ6MHBIVQJMLD
Di8SEd1EOdEg8w10CtgbSq1Xg2i0/BXKYn161iQxtQ1yOAw0gMcW5pDA12hvr7nQODPEkwxyB5Yh
tetj1BPBD7qxt/gLhiigdE39mFFaKcKVfvwDzlN/NqSpp2xxiNrhF9okBjRivvisSV1IzY4O6bG8
iO2Rqoxjy5h2khbvUu+oK0PQGKd60YpzfIqPwInR6OdihqXFDLLIENKRxW9iVMRqHReKh6cMnpm9
tUajf6COp6qon3p5C8m10Wo9IKCYudtYZ+g6cBXIBWTJ6pIW+frulyZOLUHwTBIgMW3Rnondt+Fi
nMzJUiQ322q6akggIjWnu/5Ro8e1ZJIfBWeV2NWLM067ASDnf/5Ax/pxESIiMsXm81deXrcDFQf5
5YGvM5vzliJDXDJ8B6KuBIfx+R2D5T4SKo0sJdhV64I7MuOJnYFcMB+HWXTtSUwAf3RPCGzXpV6Z
+lI38deLnbxyCAUgUp9F065jJTTgs4VCvH0co4W4Mv3RsFCAmnAnetUND7l8fZOPC36azPfga75y
edWqfDBvQ7nQlDDTAnhpGPS4qYV16rXzIB4MtryKwzxT9/HcbltxHfM91Jnigf4FPsynG0H3vgmv
/vK/4cC5edrqe5WFzyzL4wqHMAZ7So8SrR8jtL71BYXQb6DpMcx2k1mWl3NDgGKXQQ+RCHhg65Sx
Tm0PIqhe9vxlcadTAhKfFsTB9zo/qWBh/SzVI6znMy4zpQ1hO7cYHiY1ooluOcopyWIDdm/f3Kys
ejQy0YheAD5j/U7PqiPdj3xu7CNeFllWpq4/dBwjEVlTV7PiCmLtxVvc+f0gDFjbyblyl7aqE1z1
FSRXvVK3k86SoChJaKDCeVnak9giUqdWwiDDQjmV5EPpfBbYoWevS/TBGMGKIX47APGVpxgqry5W
BFbOZFh0e/PU245ocCgZRRpscXV+kUpeEfCrT+yn17eVV9NWyLGh+krKhZ4kLKHrE8FQzLqZAXXd
Q1k3OdJUYKHGLmuy0RUTFNS+BOmgpDdoi0vYCRNAIw726DYSzPqsgDHZxTPK8bLW5ogzRmBAA6aw
9852Qxm1oVlbts1EcNIVv0edPM7IBI/hXXb1efohrZ72Uv+pKAifa9a/bGh+E3yRItUtqS1B14I+
edPvT8+LXL+7de+XsVEcbffqdsrsekyYb8wm0i2VvzL2S3sDXT2M54AsGBS7OuUMgGT3Le99JC81
DbZ5NhCBK1Y44IJdTyd8FyN6hcuMXG/fwnDAcDSOEOAjdtSd/a0+KkthoQH8OyhWxzNpdg7B0e12
xJXJh45bRJLSkWmK55AH38Bl0QtFDY5Jz++HUg+AB0TC2jQ2jgiyK+8uEpU842RDS3plr475URbv
IZ1JuW+BsgFGSLGT1VrVeo1mFbF7OPB9TMRSHbM+FwtBfd+9YzUR/Y7yES0I7d3xQDY8oh26U239
0VN3EjBBuTdb8vd07D8d1PIXDpjoEY30TJTiDz7odOS+eZpv7fIV6A59bXTxtd5VxoIzL9wyvkwh
zVelgzHhFjNNHp2AfHhMYQGBX2I6kGIPvP04PaSvtdnyzVZbM/uHit0oodhzbACB/ZCgJhNA8JA/
2tkDMf7xNneDgAU7ccJkqbjZq13Uztja3h6uoKgnLUx+6rF/OMkiu1fUY/2VPxqEfuBcC/ZsARcy
ktjOvlBIIA3ElhZ20gXLDP/kiyW04i6fzQH9I6i58yztFdYAMSZWP6w92ADgT07+gxYyvC+UWsbc
flBCU6HmPdMguNMxzplchI3AItAHZxDsTn+OBYeVFUo/0cupMnDT+bb73/KAOcftf3Hmg8vvAvNz
Ra5VeNoaM3Fa2b4K1kV4RQme3LVnoXopFvP0+optTAXRNCBnIbfnAH60ylYGg3Lo8+I1Hw4M+fks
hPOcj4BPRCKJFsXEm+ygfBJgYyFacNKHRoRZvdtq89x/a3zgZnIffXJ7BsewBEB336UwjpkHadiR
XjIKv96+G0hH1dfPxYMj9nLE/51egjF4azvCRvLKlG1r6aEzc0KhA9wRdSIrRDwtgyMvjqnJltdZ
oDWscFFG+65zD2b1J3WebP6hGo1gHCImnOHqnDRcnjDkSr1v60dww2a5wsR6miEFF0mNh5nSzANB
hojPOJ8t9EzNJByNnrZf16qaUeFVZq4JcnjyE9q6yEnxRz5Bknm2+V54JoswZ9vn/oIeFgUk/kdb
Lgu3HcSW7M+DfNSVkrUdJCgGkzLXJdBT3hTTmAfOeDYJZZD9r1ECnPmranUIytCfsO1ak+rqUFLk
biXuXHOWasD/ndoGVrO4LkiOeFhgOPF8LK40iNsdCkgR4G30WeQpJKYy9Nif8PXblZGO8TF8rW6r
qMwSFvGOvAIDTU9SrIvTq4A8vj1FToNOr5niqTPB7+XFdza0S362GDgXp1slLQ5szCqyNVJqRgTo
3be2Ri+wnKBZZsJ68/0Vc629kWm1CjYy2ZQ82461rX4suGNFgLAuIzAHkA4wRx10kkxtFd6Ev5+S
RLlkjzi4nxHSL/9r85m4MRRVbPx0Xjmn/ZJ1WBMDluy8+cCu8lySRN3WTl/ylQM60Xwv1vDgIOFi
RYIFmkACqyTt54GxSovG7WXGP/bpw3izouFDTrMPIAJEP5yxCIrORasJDoPOhUNeh9S+z8BAn5a0
hKs9ngsOBwuiR2P4guuJyRFJhuUtf45dHEyjjm8qRSf8KPEbuRRt8HE+4Vd9uMXbcDjL1PxPQKEC
5y9jG2JdpYUvesqvxRRzoJnVJCcKXDc6PpnPCrdfFHH81QMBC0RZ1t/HNTzz6TKkY9Ab6KfnonWW
fYo6A8yOKfoKVLC73baNYMn3+2iPAKrv1b5prayH62x8i2BXGswnHtApfit6y/X2Cr8g1bpSkSWo
Pn0gEijT5bikfnQELJFlgorsXrFqikLbVCo34rOQcdth5tInzhy/BEODJ8nGUjzgKVIm2cpnF5hj
x/20En4MGoNrOUZJiJQCJafWekWvlWPO3C5iEsyIfQHF1irjg9wPu8iSpIKpLQ09H7SvW8UdgZvf
H56+qKYHmNJE7+5zbFDDkeeXvqQwI7v6ZkyszRkOlKOIF+ohX0PqB23BDnAG2bh9+UMlmcaFM+T5
pCnuTPqjziSZU69n0vO75/Eu1DRtBrhEAyuZQdrxRFqpjYH4OCI1EENkzT3UVY/NqVsVKSOLISIR
XIcXlz/1NrSGTCguDhry86F4ZdYjB/GblcRfrU1I+vWVZappC3k63phRETRIeg9F/yNfLzrumY4I
II7Wd+VpYRitXOKsLjY2kVIfiKb82sifm23xImR9fhf3hezztgxJmlbFUAHw7OI9OERMYIexYj/m
dmyfnf75KZVuJek7JvA+FJClGeb9mVMgHSNwW3zBMVRAMJ8qcytbE18VGlyEKKawU3c0HoMw2eIY
dWUp3jRBksRtbFV/fmTyUQIc/ZT3HoZaDxWpdpM98xons0qe3moMF98qkU+GxuQBvuIYz244eUb7
7HNEtzkYHbZq+jmZDFlXWsHcKKTnhqIMkSNckeDhIGbgXrkC2mBgjfpY1MimdONJwM1pJMKgKf8/
eD0z+AZE0KSE6tyAMcpR3dYNYBbbm1TW157GnQGusxOpAlCtjW3nqcB2LnmhNZ+1VX6ep8ZQv91f
OHQ53qn3fAgPj4FOcaudETBZaEn202juQr2tqgiubDxbcPpOKgEg2IRVw1ip/DgI2pW6+1gAFSAG
WqXNX9UkY94dMHVsJXJX1hwjJIWbeW01PsHpDFaKKogJoLpy72mdpBIjDBiMaFr+wEf3qKn0Foq5
6pZ9ZS6WpQP/dT5YP+Hiq1YOguey10Grf/t1JFVJHURj2bYFcBJ3owijtXInTrVbjQ2MmAYtfK14
rqVpLO09CrmvbzqWrhjIpCGkD7Nd4yHteM0zwEXff9SdajsrLL6gk6B87DMTfznu9A6GpKDNt6/I
9f7DlxwaOF4xW9Xv9TbGfQOR0DY6BgGy+1CGzcl1JLqeEt0usUjPV2hgGTefXU5oszYGesTrnOyN
aJk9rj8/gc6bDrwnXP5wou95ZTXdTA90wbRPsWJjy3EM5eN2zo2dqtN5pQCEFVqPotyBXna1B98x
RoFevm13lfsBev3LRgjpleBZahPhvptbquXPI0z+zkkrJUXs2kqPmx85VVImbc6CeK48xHLhatPs
5g1w9TpI39v44YoNsEtSq1Xf7kN/fHmjvw71m33iFYFq9qO/SzOJXqenisidgnuWKUeBv+Ve8g3F
eP/Kpr3nAWTdcU2o0MOfYed6Dd9ne+YgSGcHp04JoEKuMkE/cqgC+CzPUIgeOLqlbBKdkF3RxKVt
iVRexKUxjEfy9OdHaimNhusfGG47Erwd+qzy0BHnWSeDTqR+Ug769fNi5nOoY9+UkmXgCSu3ZcfW
daueBepFA+Uv/2HnYktTXYRnTGTAe28fIPcwgFqFihb4t1i9LwVpLfE0ntfaEoA7mVE=
`pragma protect end_protected
