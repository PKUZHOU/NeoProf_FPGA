// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
UUWCwarV6xJjKqoj8mJdefj1OFpPH+e1+ApS9dvu5kl+H9XHvHrObTHXPP79
bQG65BKQL/qlj7ZBcJqLLMerGGUDXFtNhath2h7e+kvWOFAf3dOBOXgj3Oit
TjpY1x7BQ6YxQuOaJa9DARFGoNkHYDVyheH7LdKlKQKoUQffIW6WsxigpNtG
unzVUsups9CMcsAB2dCg4xYQWbxhFT3KzyELq0Iuuzef6RZAKrMFf119Dom0
Fz+Br1N8d0DTMnsNDprq59mnPb7PtjhTmOH3FWyCNmL7VzHM6Js93x6lAv+Q
CxfdzSNk/buCCiyIMXwxWGM71C6b8SRHBmODUXbVvg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kNUR9hhe/8T0/tAO/6+R0PO/5beQfLY/WAdZx0nzAU/+DpuHTxLCtou7n683
XcRhvwV2E4AbRMObTK854WkDOmkAoGttwz8mJ3rYD0DQ58VCP8G8u0YGsp3b
ZhvA11x1DKtAVyyeKP6jg/wcjOeNNlP2mcpkuEHYXIbABaaZbacHAT0vEXpn
fdFTwTn4l/ExmCy/95al+yvRWt0M0DX6YjfHR3iImWa2csgCBWfXC1pP6+VO
HY0Ev+S/OoJizrx9mLmuwWR2rvZGPYQYBfxc2doX34I6rAoRooKwVdcZ8M+U
licEWZ8sCCp2QjdIVPaow0tRVi/IKcNFuHEIxWiZag==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qCTYwzSygJva99WKomwrWgcyh2ZREHGczGn6z8kgPqLkQZzBaHQiMP5i+uYT
gU/CRgEjQnpw30fqbI33NoIow5ZCs7u2JJKokXdDUmEB38+mVldzMBCOViGy
LuvxOd9kb0pX01dzq7EJsubW6SY/T0KbQl7PggdnlBhQYX1cZzE6rJz9OnAm
O1fhj6WHvITVpCZDbOGAk7eSXYZZMDWT8YgwgMLuU1FYYAdfP+xhMBcFwU0Q
61TogdULolXZG5Wdd32rAKx8//Kjxqjj/ou+9ae2BVi6Kki4IMH8MWSbB3dj
fwEXit5jPQT7o6DjobMKsjy4es1FLgYmvyIiSaanCg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
RwBD7vSzWvVdMjUEwUYWMNO210NSe0f3W1/AcdgzMtjtgKjtM13XONdE+u+g
Gi1EQVXx/wGoyyg7gJ5uFGYytEvrQeS69EWpr7Jv6tz3IianjsVCnVnHiLAT
l/xA8QjNK/Ojp4NeEjATDFs9gmx3DKkRTWezl6TXX90iVydXUFs=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
px9loyU9AtG0ZEpsNb6dXb7kOezGUw90BOV+Dc+D3UEITx79fynV3zegoR1h
KwzQdGw3kVGz4jtqkojYhVOJ7XCA5rC/VMOGgK0JhDL76nbjHvS1G4gfszBB
pety+csw2OwxdbRsPT4Z01aveCKuzabgL5G4xTykhh9EFW/bck8E/hZK0c32
IKzz/fnsUbogE3nBAjD0QSM38zEsvlpdmYh+FZNjQF6OJrTriKpSrZdHY2Gu
huyEBFH/2iVw6qA6eKpyl9Kn21NlAldnxW/B5IORZW25iKxUCficvcE1+qjc
wV9cbGtTlCx/Elm6FCOMYB73f+vWnmyP7NTVmiL4ZdrtYJFtJDdtZ3CsxMec
+t6waw9kH1d428oVklnmbNPoZEJyIrp4aoGQM3GFtrKkH6QiOeIozV/B0LHA
HTkXulKf2xs2VNdVZG7p0Qn1T7vq/jztt/GEscSB5NZGo1by4M/LUH1RxDwi
rVgwjutaA7vTGaLuBcgU3sLJm8Jyu0xF


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
H13tYcJz0f6XGcY36vW4Y4pf181owA1SfVB1GWUtQ0F3uCbNSAFIMcM9rGPu
L9vm/t65faxW1lTV+B7ZOnQ56n/GPr6+dDdOFUQZzc0oFrdDF2dQQek0E93Y
YyzDsdBCWFUE+NQFsqKzO9T+9Q4G/sJ7L1tD+zLgx9uUBpOBomI=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ikNCd/1Y3ax/hDTD2DXa28sqpwI5p4pMj/B/uxgoquQ4eqBsx7wk7im04C4K
crQP9QGcZ7iE1aSgICZbiMcXeKID2jnzzepSeyiJQXWJG+YwEtCz3puewnFR
pCtBETpLYYoOPJxlpPCx9Coic3+DCrWe9Ig/FGEABrP2SV5X9HI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 49392)
`pragma protect data_block
J/vjyQnMAprYmhFsoLIlLTiQ3vw+wdn63UejyJx5Z9hIcIPnM1ZDDlN3LT/2
KwqBSyRlxOiYjgw3DM9vVcLlTr9kUbjYwngvxqxQ9YcBBbgikW4FDbxu51Y1
GhvaxXApEZ4shrJu2Lifum/r2pf3Rye3sRCB7ulViezXCoVh7iWBDZfAkDFm
Y+bixwZ5hBgh1gC9dmBXfrO7y0K8m8Bz4HcTReSw+ZtATJ4t9/h4lKnUQZyP
sjz7TVttbR0Zyh5Ej6MIWFO1ZaeNRXHaZPQG+x9CmyGYLG0+u4MvylAZKSea
Oa6wFiT4G9wmSG5kJowmQoYj2etxrIBsmWftvLSq5nRa8l5zEUCZp9Ct2SQT
6xnFs7q/sFbyDL2iT9i75A5lN/raaTwc/AGd/wln0CmHrtqNmMSFhAotB/Px
XEav1NZfkV/UfWAYZGA4ilNXCnb2EzV9xnZRaAtRxtsqjsQTOFCQCJwgQkGS
sSk5GQ5D00LsCVZmsii1x6SXU4LxdXkxgzcVOau0agk3G00kiq17C4HFmNRb
QStVYQ6+PiY/66SIGyP1T3wVdXKU+phuz4HGkWyqGHfync8UjXEdqV7AwCPz
ZVs9JkzWSiP9EAD0tX80UsIA//1g8HwZ1vUPBFr0QrW+x7r+rM019LBv+cVy
JVOJUI3P51+IaE9ROwafFSdS/1wWRoquSMVpejmks8U627maZWcwTAtBslYs
K1caJK1jM5NRQY1Hq/cr4L9mXY5WJFbl7JV6txP0DFDMI1RuyDvTNLYr0L3q
K74U9XE6YaSjh0WG43AEX6a9YpOtjzyC0bhcIFs7lZTTlUUokOMMoy3qUEKd
YIsmYF6XHt0Pi0xFX4Mi/0B82DjnMK54RlhZSb9l7LmuYMhGh7m+XR+H3cxr
8mYN1fh8kMOXukBv+QK2fEZ+7hDKnc1EpFTcbySGcsmBvuFZGBh7Bkugfl9U
fZxo1/shOnnwIEB24cMiKaOGBq7a95wM8UKophzUHWo9rPI7bDNOxJ4aKUaZ
KtxraXCzjwj90hdnDfYqvg/boDb1Qsk7JqDRPFLlCoFpwu8aBgr9bCJcx4tA
fs+vSW7NgrRXppkZAk2wwhzyApvprCZspjfg1yCFFXNAPdCzTH1l+/WSPKg5
WEEDNINsdCTtoPo5cetuldLX9lXkVPuEKkX/jo3hC0Wis4sM+pRqr0zuKQ3S
1vBmx19JmG76xb9Z3AActz9M7xOqhm/VChndXgxOE9wGlV4UzXWgsCnPyFbj
IEUAmqbkhMeDulN/b++CBS/rK8vZic9rRdNA/o8PP4VUae9N5wYAIO//bAIc
oMeu8Z99LES+qkx1F1CtzPv+aeD1ntdpdky5Upg2nfj+ftt5OBqX7je39PT8
GGr6qepFL1utodA2xy6Y4o11wSez6JK2nLRBkvHg+aE94mGypqRRpYqh5GeY
rZhOb1y1qTy7t5M7N8gD+PqBKhNdUUytxY0I8w6PWVpSJPfy+BcuuBGrFrTF
tBxn1LaReIxKLZSBi2W2557OoljBteb69xbaVIGpU0+Ho8cBPJpPzXq+2n+i
KOwxZ5Oq21uPAFVEwy+ysCQvvHcLeWvg5ABpKyhxYfO6U2RtT8NeYTKid0Sa
A/TMRqlggRh5zDzRsCuid2qcqljTxAe0sDcw2QWzCibpJTpd0jfiMBY9WkGQ
D2+cxXD/qFD7GiObx+79oesGMlhRF5ZMdkTZ02Y+yFKnJXAS55BtBhf07Vf8
CY4gp9ktqHLTZi9vXCO8Um1Tr2GX/5wqPM7vh5TjfMA6RPgB/F0Svsfju9Jv
n32W0vWcdw5T9K8NFmgT4TrlfyafJr+u/vHfDEcGbPNZfR8utehh/4CrryX+
mR+olE+C2T0pWQfu7+j19a2zmhmHGgcOjnPB23l2w4nOYwwrPKnN+P3TPKhn
TTloYR4/Jjn8QvrKSU5xs/EIdQ1HdhgK4dZVsWvAml3GH13WJxItCa3a22HN
AvxfttqzzMpiR5mpSUIvTGSDdJjtawblIF6P1yjXOXpQKCo04vka9a+ogO9n
iWlTciKKvcS81SwSjUa5tOhzXhu5akncVutMDpr50pMNhibrNPaSUmzS53fE
uA/4Ni81NgPR9Zt+z3dMdY9gflC3n1rSpi9Yzh49eiY8PuClfoPowW0s2iEv
+vHAQrHEkq4yYeXdGMra/2BoM0rcmfyVjo10YA8SijBbbtDzpOtgk4UJ1Bfb
3FdgqNUIRR2dcZzC4/B7YnPVZDWtp7PQYQfonLO4/2BLxQzGi+YbfhnQto05
96+zfjsrKk+iJ+NCqVd8ooE0H0OeQZ9quNN/jzH3oKT7ViykHpSIQIYdrmj/
cwJfCnx0494kJDunqoqFG6xOxIalNrH3HwEjq0/0vJLt+sQJWY3dTkI1WQlG
INKiKVuXLtfvaZNURUGtvSyYfOhPqyOApZfPxw+tgFM4OEv94xP5cPTWR21d
S0069dK4o55BUzulUHAZR/JzEXQGkzhRX37aOVJZrz1Q4Hx2FMBk7GycnOJB
6TkrJcCxdkhpbpst2MDeMeEUZIhv1KviOh2RfAtmjSc9g542ITizDCpb/GKl
TUN/ufdC+peEsvzBU2XW9Vt8P21zlwi+kOl6vfj+tJIgulWY5zRJTCLrr5zF
SSpTIHN+q9XVIjUbkSwPA8FTYPI6ksw4U6MYpbyhTYQzdtm+i9XKAXkXZCf7
l/mUndLO3LtfOaJ0HUwSD09DRSOnFZ+zGpXjzHkU74QCCDnfibjJI1xVYZNL
fj9pLLUsCwTWhjNTLoKrA0AcE0P661kyNgNY90Gp335jGa9TYlO0q+hujwH1
wQ+hGW3L76kRw9grNf7NEKQ9RegK9TwYHc6Q8P0yrGvSUTb3GTziiMY23xrd
E2IA5nj0Pd+vpl5uDkGUBu51DpNeOuY9tHlKX7ro//m8MKZmSQwkSqr1iiR4
UpqMd4BXLbpNxJCHgl33TkercKayaKXmhS8ppuJ/U0wKiLYWpXZDYjE9XSBp
1lFmbsSNwM8BWECiq1iGqh45xQV/JdWT42li7m3eeMm6+eZkdgDrdkDkHRcQ
BRkyntITAmu8utD2Rsyno9T/ttVnAtCDZ0hDHh/uiUtm2mG0EYbM406Y2CoZ
mE7tsPRX3RXCwlHtHSPhPLmoqbVGCdKi9C/Q4ug7bT9Sca93HtDKmV9eBzyg
UwxT7rS0+c6HjHma7lu/7e4Cfzqqq6RjN9LGGrl7SfnOBQuGM8Kje531dmD/
n5gEdMW6soVRs15l+DXOhyKwU6FK13A3T9X5xMsJeBLR20mZEyd92FFPs4vI
4mVxNwRVySs/hOzgB1SXH02CCE/686gPmH6b0hePt5cnQFNMrrYH4LWfkrOj
EvJJ4RUTeVVoNHIEZQCB0o+6o6cXqoawMa4gA2hxVz0XVQbNRZMrvd/wQNiA
FoACgGU20LDN6esyGW0Hcwz5XNdftcVX0WHgFZnmYHE+EBVLGM4c8rzFLDKZ
egsx4wP7XXZqGR9OE9+RHWod93/OKF32w9lwsU5bDGHR6mEmBQoyph/Z83Ng
W0Df5+Sy9xZN7D9/5TWaI+Gx0agaHFc5xzrqRsD7eKiT8YI410gC9SmYyTc3
HcOmLUDHQiieQBvVgjWR/xsKZigJuUTc/v0qpaRl9crlaBOvEDGNZC3jqDDr
ovOIcDsvg+zPu4C3CUUshNiHVGhaCiOpQr4xVkSCcc/Y5SfGfcKhX3mna//W
5MsQScWLWhHtwcyZfnf7kBt0iLrsc9zYlGGadMJlNCKD7MQu3KHLh/J4h3TQ
AVIcK2AgQTV5W285aYd+UeIRs0YmMqSt5VmvGfddPsZ7v1MNNvI8IyCV10pl
XslWJAUsZpCjDgTVcxrJCzFNLxmq+Vz6uVCyvYsMCQvxMKb+4362i8GA3g3J
tO2ywSh2XgP6yhaW/jO3tBzJ3YggNF7qDeryhybl2TLYkL9t/hNH+KHUCdkQ
VM4R7t0S3KTC/H6jolSMZAwZTlVETebJ3E6gnSGS5zqIkgpa65EJuLfLjU1b
aCX2+I/gBm7yBC7zgfCGEiqBDfBnqr+xFrvN0kIQFSAAMCQOIGVP2fZLW5s9
UD6EdNptF+Rp3+pB2ksnh/lHOij0rrzUOOeDyoTJcvRunDuqhcsgWwYFNrH2
xmxDGbxHcY8ily6qH2u5o/cR0K3KrOBEKggktJptJFPdKpdCyTzFVaLo9lw3
EK8Ro75p24vxm0shFLivFVqKjKd7ympVwrb0S2PdoLRcKvPwviSIIVgw87E5
8ZB8og1Bvsb2S8Q7ujpU5dW6D62fAMiASR4giFH54RydVI9qXCiBQZZghemX
eMaT9dri7lFaTAh2dCiGvvDVQP+Nkh5nRmVTXasFG0TXsmc+C0Ntm7I2cdCb
YsPKVAuY6CL1WyBTwls0eo8UVLbmpjY/f7OW0vqWziVXQxZN4GAnPx/DcUk2
VbufhHPEWHFUQl1TomSsYsjrA3G1lke01VCLq4R3RtPiUR9Uz66+sqFCTTiV
SFh4WhkPiVFkfwxdOpfiwq4Lhc6YWRG0hPReXNJZeYzOZDXNz9ewjCsic7VW
LuhyIKfpcBARBRzwGGa9SuNVVkps0F43VIPxgGo1rbcIK51nAuUlmmKa61D9
2wURuFewbcn3958uLg1s+GYE/5tbgWj+gCL2L6VNW307gg+gMM5hY0+twUu+
Q3wdU4acPZ48e4sYQJYfVRPiXssbHGqCbba+D82HPZQpxwtWPusvlytBFBot
9VzAKMt25SOpp1nPlnGBlrAGZRl1pXoeEI8/CcoF5pHwZhmx7beA0Ck/Q0Ba
3hRJ7/OxHwv+FbjqMesCl4ASyAmtiSW6nJAtOq85LdccbXC6ZgNhFyWiWcgu
9DiMzEJZSfKNlCi3H8qOhUicrAc1WI4v+CuFUlfUbvrOGe2uW6+J/2yXueal
p9E0kO26l4amp/ktD8BAwAn/ZfA8yX5wDV3uNu+ZgBoCl+3CPBnXE+j5XOy/
pImfnr1TIf4WQ8vWTzY/xBiS1RPoTIh3OsPXZlunFU3XnU0g7Ab5ilHxQ+kb
1n8tDHI3HR4cvHW38h1X0kQhyt2Cny/2R81u7QuCngqhojym7DyEbvyZfpuD
ENSIe3igbbe80IpfdpCo5Ihd4ALSZCibGs+mz0PNOZheo8auKS+oM+dL2n/I
U79wSevgHFkf0IbTG3AYlQQwp5R6sFQr4TPES3rSlp8Zl2ImqlDJHkEF1K2O
03oHSDYFLkIJd8DQtUYP2u4gY2MgzC78Bycsg6rGnsMUqQCWFZJ2VZuNuKW0
c3/4qHH6FN3X0/OOsD4ahXuvgTY32Umfl5lTmGmZZk5xBxSWyJAArr4skVvV
jLrnt9o3onczUhjJ8C6PoJFfdHb2G93LLOlgjTvUStMBOTfb0rCgSX5wHa7n
pKlYuWnUSZHShLKT2fKX2SPSJTlwqkIgayyDj/RkS+ejZy+YkC7+g3PZ2tP1
aKzJlFp525jfS2tBILxVU9Ywux/HeM+a6V4ECO9vEoR/RLuT8MoDkTk7A+Ki
jONAirFndYOOUvKb3WP9lu/JEXES7ADI5epuN2OaIKq9Xmu7/ijnjMdVujh7
GPT1uLGRuOjYFWZkE3WY/csWOpMTlbXQwEuNI9Y/eMjAm07kqnpZv9cFEr07
J/PUaeVgfBdpHDkmEYil3hp9tdxdNCQpBPhqhW/XNmtMgMMTy/iKdxmPdVCS
sGr6g81/pHuLFcm5hcGUhQkY+5ayibyuMlDtxfoW9fqFe19tHxU7PqRAjjCi
AHVJqCxlTh9bOADMr/rUAXXXklb3cLrBclVfbTwlpj0vrSPqKnvff0k1187j
ZtxU/rpyVOlnGiLqH7IqDYLgrWHKTPajuzm4ve7Jvg81MWaBxVD7p+RSze//
9tPJ3s78WsoMcdWXZe9/LiuDROt8jLkggq4KOdBN4iYQyY6a70H/kv2E9nAd
RieavHq6SliyUDl5GfpJBSFzk4s3AJfDuVF+y+d0xpixuJYohW5z1MAWEchm
gzEvN4vsf2/5znoZMgggqaENJ9WkFDRgRK7ebrcqFhPsOFjF8ka7o9Ut7OFJ
1nVE6BTKvsNpdAa03GO7wCJ3VN+mp8qsmpDZGSHSNGBcLjNjdxRekFifqcLV
cNzamc2y1Cly0qV7sGzYAGG/yAqIsMlR1snHgN1Y4l0QNFg4xPLinqtkpBLc
72qSd+OLPkueIIc/xzgGHnEiADkGbJcf/zyURji6JP5vxY6XD/pbZhXrHP1v
lKpw+ncmg9btZQF6yRMzI5WaWlwVW0vMHP34ezrZ5ecvm4YDoBtz3AdzqGLC
r2/o1TssBClFO4i8QnjOfmrY0h5DhvSy8JDN5PZyNtlH1QKKjl13Ctjbnhsg
xze8biMVZN0U5Myg6AkFirrxaKsK7bUXFC+ME48WPqzFlOuknkicquCSaxxA
RYrjqYmJX5zIk2T3+qonINzP5tgOWl2M+ruuv0DsSz/szr3ENPu2zXWItfNC
mujnReT1zC0oyER61BI7ncCVGyqx5aG9/EyCIao3fzyfGImj3813OcXvnhYu
zEt3hTD8nn+iiLjwilqCdWkNtxEeD2+uWTiRAaq+c1QTvZ2P/LMzgJnE9dGE
qWdvwjB12ws5Rw4tYjgHi7DA8M1XPVs679ynAtq4vY+upclVggNiZ8kYTNNA
SNPVpPO9EEQhqWuAC/b31GtqZixan7ckjoC1Vwm6odNEN3kqwaFBh6QyfBsk
/nKniZH5aENeLF7ixLf3Zas7uUuH+G+Z9jaSDIxDTFL2L0hU4YjGzH0FY6GX
eABTzFLViSg9Mg8BV87RBpwLGyD65RJ+Z5Pp93a5WcqdbCCQqlBbv2WREvs6
/s4qkeQfWtPcm7q9D2eybGmCJIBKlByCAU75GJgw/dZsOZbEx71jKZgfl6Y/
b61sO/6vOrl6HQHmUjUK2ei9U8UnEWrab7+czFUVxId9OzgKUBrEHcRGcFTm
qyy8sUg3EHQqh0HAg4R4K2eD0R2StpB84SDgLgVXj/NA0eJqjDb2PhXOuuLa
YhrDPdM2ZoZz5fAAkPmHxY2vV0WUOcVWJKQs9NmA9wcIFIKO9I8t0EPKqx7d
6DNiK9k6dzyjhJgLKq/Hkeu6tF7fSLLtlj+m9SJboKBg5nsCU+mkxIAwlmFq
F0zYt/3gLAodR/1ns2Jc+Goltp8UNMz3QcGvlGv2GOXFuB+GXZzhQ2pYrP7R
v8KtL9YvjuFssT8aJOA0x43TTimEn12O4gMru/tmbzlFHh296wGopVt2GoCO
/cEXjiQC4LAtqDbohmDVXyUFevXicAu4Ln5ftTu6rh0uPBJa9Q1UZV4Oxr+j
V6ZuGALDB2VS81kgdC+3PV6m2zkblats+Hwr6KdqI5zcXZFEvE9yJs09Rinn
HfYiNM2nJTv66fPGmuMg1zcidv6Hp8i6K7lsM/VRmgugJOb6a8pHzC6JE3A4
Ly/rwLelmWMinQB3PTokA1nFZn6GyuP6woK9PHOs/znn2uU0dYMWSkvUaLFm
qiT497Gq6e50LfSMoIXEytQ3FnrgdcI2RHmHBo2g0WL4te70KdFfH73HnDSD
CvgcZTpIuvC2mqgPVFMaAeHcvNQA1lNZJazPY2j4hwG4Bt+wzicWXtMcKzoP
ory24/XtJ9XtRBn1uO11Di2SKJS3neElqvHpXO+SDZ1ixp5RlIi36WkgpJP3
d+8uUaw942bMs/ine1sd0oqexBKjYcGpKm3+w1TuNe79rZq+qEsBC1FBow5C
hAUpB+yaYTym3pIsl8b938CvY1coEpfgesUjQwyFTQrC5cKbImq7srucbTQe
XETIn0rJ+WfFoetSbKnnXuJ/cTEOw6QNFg+JEWe9/PzQ6xCmQJYyLNMZb3dm
qBbOk15hB5A2S3KVDYX6Yw5oT9pwi2ByFH7yZMWxmU8rK6+DhIJ0V2WL6/7W
AvIWTsuSl0GWBxvtAd/Lgcy+xpnbGIyZ26FEBONGym3U1nLPIZRg7xKHrWxG
skHjznFTAE3KpRagT5AdRwGG6GDOXmxyFROXVPVnFWegMhowYuJHTEgyfXRP
Dr7gaRw2mQ2drs6HLwTDf/UcsOq7TKosfZEJZO9QIfk3AymikY6Gp8pvXlvG
rtsnlqvdouFyzyH7ZEg/Gsjg+1TPC0vJxio5cdGmTL4JdnkH/gwifaJk85ih
3Z/34q7CRA0FHu24tPk7ZglXbu8ilXBlCJTxUEkiUEF+QyzeSWVKJx6WYzfl
qlb8OQ6MVzAiXOyhNsyJtFdOU3OC8LFTj6Qoo/OxQp0BXptv4W9mS583UUEK
brZpP7FLtSM6lDv6yHcYaqm1iL65eKAcpJfQRvuM24IusYY5Uwi886gF7dk4
e0Mhy8I75jAiwm+jD/pdiRDsGr+sK1Hc3hNSxvAX48Qc5f1b5qUOGAO+X6HV
mzD3z17dgESmtj6BTAYEPppPcObwMFpN1HxC7zTbuXI2pDbDgbtUcgb6Bp+M
YvNwGHzsl/KXqKbtAJyAhhDhz3lwwhH8sr4GVoTbz24aChqbgySC5pL1NkPF
5bPF7ZXDJydohADBDMjjb5L4/1KnvvUMWz7QTXTT+hSN5ZdB4cuOxFFoq8cB
828BB7pJLJWf7opqeaQ7PMRKKlxJ1Q1b65gfx2YbhALRvVIfSnidYG+sFFuv
JUEk/UMdi7Jydqng8uGM1jLAqghHY5SPu+PkN/rnoe95oTZfqI+r17DxefCn
WceTaaPpNiUVtXzMgjMvAl8atRqC76LqZiOhvVmcjvJO9P8BW4a0i2acLlsj
A5mukxPonOx9S8dbpjwBppFQPCEVeg82Ns+1b+8NvfGRUem6BzwlVGLX0PIx
irJ/xNXShg1/RujyTiH8wz68pa/eW0IROVphwJLBkLD4JtSwAM1XkxEA//qo
eH70RNVaaK42P7Xe7WMb5xWRMTh1/4gK7WgJ4QP8QxYXkVFzkIHRv+HWC67E
7Yu+PyfW41EgGjSGr92HhXPH15E4vi9tsvGl8UMejqicg1koTZqMFBsvuysH
rIbXJKDxubZON9KvbftUsDYHBZEgoMgS16/Cs2Wvj8kR+6RRJOl+Xpt/7PV8
4GvVeEO1ZBtiWjVtloaGUWN9o0z4FND++0II5zpRflZ7WqllRpxcbCg1aQLe
sB6dMLlKSHVeWuH7X9iJRMHqEjWlgojZPLG7JESZ2ZA3LB6WU7PDrrh+bPeY
mltE3Uid8VJMvge+kaC1xU9HiCX+VGE3RPIDNNf3zGypZ5rQ8N0LH+K7C9lT
jUkygbvORCKeUkSk4Th0w/e6NT0zoHs2k5WxCeb1QN+MLco6iT0HBt7sBi1W
hYLNuQwIl/kbB5scv8wsd1EXgEWjICXQ0mLnN6bJJxcpG66lFVprZssCA9sq
9JdkMAPr7lapsW/cksLTfyQzY+NxS7je9R5h+lWosGvyn4bL39vY3ewQMZzb
ubLUifhD62QBwecYvtUYvdTzoDz12Uv9NRkCkitnJi0B56cGmJ6nHKykzj1G
OkyL/mq+HyANuUAn2Hm3Bs0PH/2qHCbNQJpffFt4QvBCht2H3N9Vnp2KPZje
p/Pt5PvW0PlMkSjikEl7bspaDGFp6meaqed1ZORdWPNAOfgesSvtBTPdZ/E7
h+xt0jm4jlcjvDStgDSDplcndXNt99y5CuqxPFpU3rFUMb6PIpS/QB8U4Ix1
evh6FeLDNhCT6g+CuzHdZzdNndV6bBkB7Yc2l6snuLMcqr3qdkXhdoriaH9t
UNqWd2Ap8s3gUFyGzaCDrgJmSJkAneVza5fV/lTP+55oCjv8x8IPAZ62F4On
lZWUSiyd1g9r273ByeIy5NYlFLCyQtljrCDuSZc61akpa8qphNbLhXX6V7++
tR75smSAmVQNSGq+fwibaefvj9iOh3OV1Q2CC6tT+DsKq9kh/RVhIp3RyYPA
YqiFUnjdjuvOYyOEDgalnQVi/sS0cCDJYrrslL0J2qt1VMlZfkLKNIMnwEjz
IdLaF1Ue/jzhNxVn3BbkG+xcujb3zNGU2dTxa9nq3OTVAisuR5JeRwDMTtua
F2P4B4guhtG7Efge9P5CdmELW6OWMG5JVN2JOzVR0kRb96jvOV/7Ctloe9xf
SSFQRk555LtvQTzS0Gtso8RQwEo1E7uaXq2TEacov/DrvckNb9vVY571wZJ3
PrsuMPgXkBxOjXeiLis6K8gOw4LztPQOmfRVTnFxn0yIxx/YiP7WH0W6Hkuy
pEae6VnUlPMDTUeY9i+eyYHRT4kScOBfrgCdSaCcu79+6fxvLsk57iq4c+wy
VAVnBCnkFxe2Qq/Gk4P1T9qkqN6/JSCImeXRyXM+I3h1N8HmPz1R0Hcpadgf
m0OSDmnqNC31yAuiTAWoGVjMe3qAoegvCRLbKKcnzIOlsJDC8R+We4Kq06ot
WGJ7ySidyL3flV2NvosQ9P343h33pqgymDfMdegibks7+dHsWgtXEmgRjNE9
i2yJaG6e/cD77xZ2XrTomQ2emIQKeXduClyPEjH4ahDj0n2VeLiLojwnWGkS
BT1ybCjPtdwC3usoHkg6aunywEmlSTHb+s0axE0p13dOTFgtbg5L28ubO1pz
RXzEE28zK7JrkUPQo+ZGX7P0cQarX2lD0ftO14K20Fx0tTci0dOe4c+N5cnv
cTLSvMyKEb48B1W5p2VNNENfXoJwdmid6ZDFq9GFxgdNSIsnzWCJQnDBzm01
OZL66WTzEnCWItq0JD/ZQbizX/0nH8tmXYXSj1Am9Y2Gpc3YBNDfnAuOPagI
v8zieTFHM7xB/Uvta+8zuUWjiy9nRsDxQ56clxmHvm8ir8cpztW84sVqM/+O
eeJVtxpxjZ2tREaNxQKiPPsVsDqPwkgia4RH8W4PQhf5sI2TNahG32qZsZIc
GnWpBETBxA4ZVkGMMN5hF77me0BOyoBT0FkRggOWcB/52xFZOGVenrstWSJO
a9sLXaLKP422oG1kNyxjIK5S8ZtfGCe8tP8Ie8ymzTtq0yqnvcTPLDWwg3zl
QYwuShPV8oG3rbP4aABHMP9vaPtIOAHfpGp7MsgKg0eGdV6tG7E3U9YMf0Tv
K7JaY//N0yQgqO3rnCQECpqpV/tiJQSUCoIfJldSPCSStvLHe883qdi+Rfnt
amLK8sN3H4105emmU6P3ip3k/LwkaMJunLKUFe2FiAawClpvGWCHfhaedzym
b92g6V6Hjdg5Yt9QPi056R/5NNxZZKt2N3eKHhQyDSTnBmxqwAhoa8z56gz0
nypxY0oV69O7iRmZN0Z9ZWFuA4ouLJrvMJv8nvL6b7Vm0t+iRDffo2HGBb2W
amuH+XJveJsC0kADp7BDJNXhOfFiJFHxtLLSV+SkbSo26XH5BEM7enkw70p8
B3DFoeoORqzRmiu0A+QZut5Hk4CxaJQAe3J+/LmoNYi87CqTsuMOjQCR49GA
aXNoTomg7/ScuZCfgc7K5GKj/TdtQNhePRDByteBA2K4lTK2FFgBeobbwp1C
glVzHzZoRZnumgl3alGTFYF7F5fSA/3v7FfjypM1s4vxbPBy07pxlV7MSdNZ
FyvQ+rBXZzihdSJhy8kD2OGo6CJe7h3TaNvROl4UrsrUcBu83oBFZ+SNp+yo
lygOpvVNgWQRiXtSpgfDigsDM3hC3T1RgM4S7nrI/PRt6+HE9/ioistnJOA/
eX6dF2zG1BA+PGc5RDd0td3+BDEyKw0yTGIMYd18IBUmRv8ep3Frysb38m8z
TOt3YyQgmOFQB0sKuTwU8X5g2+qO1hvZu+1zSJK21rOxThVG1vPSpbi9uPT+
PEUOfogRY8h/y2XYCG2MbLxJ+yy8b6uQRbC5CEaHN4XFTouWRY5MV+OKnusJ
V+ZfoZE9KeZoauZ8hRYb65uZeorhUc/gICGpqzqL7cezFjnp7xhpki4dWiD6
9DaStKTpWgmOvOhAWbV/UK89rK/8D2wykSXoh1wGgvE0sV6C6OjSGjVDY2As
r0uaGgPW2pcgPbLURIAJdT0fQvPsp4oWa4d/uFzP8m5/vXCU3Hc9X1AAd7YD
24vRlpr8Ui0SUhD+eQCy3ejwbdP1JwqUyB7uKzFHLSqwkkq6XpYdhZj+whXW
YBL4SKaxL2F0fcQf3EtpW1O7hlp30P5rVr5pwF9HT93c+znwRp8gFUEjll+z
6cF/ydttBHreNHjrsdnzttQ9zwRrox7w61ErMxPG4Vojz5GAP1n36Mh9qG+h
xqXa8pdzxX2yXWmgfVJh8rm+Bl1NKn59KXw3nVNQ1HqV3X0vxdUHeWebVeoW
gvBDmrokmPdIW0hAyPYlGljbzfa6rIlWKtfjJ+mcHDQwXBS20FGoHyWwhHo9
i4D2Rsz0r12Wt8ZwIkMn7CCLEowShpzhXFOskcRpnP4ISIKaF6XicHUg2RJo
qrxC/DSKp9elQFDoAld4/TIqdWS7SidrSfs1TyfkMKkAZ9HpB3P64LWCv/zy
yFe+xOgGVm15n5Of5aqPMDKQ9Qj1IhXaPsEZ7d8obRbBGrar50ZY4KPFFcaL
ZXQw2qZMQuz6p4ST//hsLxmqAmpH66EDZ55y8eybLCnnVHhlKANNycXCWyRh
bi+ZutwWMlgzlbSXYQxPwI+uk1OIiz2uuOhLcLnjtXydXWzJTlQORMWsxvAG
gboeP8fJ6YcNeEAO+cLb/Rn1ygc2HjycoUhZdvBHGxe0sQSgxG5ys7XDVvZZ
4UfG1ZyRpNayZkKJXVixvMFJeuXHekxEThevBBjaPmXi60bF6oyhis/npIoi
8DlX4usFqJlKsbdth5jp5dm1Vnd2DS304t+S+mx2z/zu9edZ/dztzIo53cui
Xvf/RzEq32lQ926vaFpkMEA6s4HWkOuYRAfYVk2DvIrlv11orHzSa29KXa9e
AfJY+sq3CnHW+egLGg1FenvC7SeL1v2BqopsFmq8zZCZLNft0cwVY/63+PL4
BYDcjNPdMvRXgYuwX7qdglxe+S7m5rRmZCWeLuKEYNXE8Fh5Lo+/Q4jBiC7R
9ydLqQFV5NJWxCyc7tBpsHcY24MQLRkfFcGqFLkIym+Y7xT62TDA3ASYZKnR
hyFmnngXr0q3ibWqL+PHx0T4eWTuozlwPNn260nrAfvSAp1Yq6pjvxBq9Otw
FQNjWjUAuedLXE+YRmBREqfH/YyHMr3QkzJrsYEmTloV53VYXP7jSdvpb/E6
yX+DdnIhVKPnV0l/8Wkz8c3+dq2ouWNrDfRyubLszbvlP7qqFhQTor90kpCY
XRKMGdm13RqSTnAHQu5Q2YaHNCW00K8OHpLOkLjAaXFa3coRWwG13v5hlXrz
iBo+KRV2iygZzo4ZiTeGtvphq1DFrVHbYVMKvOEXrjQ/AVFySTO8b8dRFFlP
kCL4YPOVyZw3xpoj5fKySLD3ReDrL+M359PtfBk0P05794EOqBn5bzgaFH/r
3Waygk/Nzn/uIiNimbVkTo01idypwrkl607q7Q7RFKPnVCChtlJ30vJP0f50
vE2jVGSMlhQUKPTE83F+3Ao3zGGxvEaftPpFz409ATpNtQ+/FajgRAVZg42d
up/tvzKfiIIwotwR5roe8HNuaZy6emgJKwvKfx/irb0FBWyBXTl1bdbrHu2H
naWjmOuRhPNKBlAJd3Lz79Fcy5BZ3qrsr0Z0xIwPQK7ds2prgSBiBLf8Dmbt
bDafBhQtkaPoB3qFClO3NDGXygTlp5Dd1bn6LOHRBF1N1fk6vhdfUaiiW9VN
Js2wNG6F8DM9L19IdmAnfOudWiEIDLrgJv21p5L7CuD0m8vzB/bIy93Y+r0l
ZMjNAtR/UP2gSVoEny836hM07ZVupN/LHqsACo3MwXA0L7+tzWRlpbA7H3JB
MstyJ/9McNiCKve02oWCEb9OvBVlBBtZFHclKPvYqb6xvLR9+ACxG6Ls+2qt
mxgTTKhn/2B5RqA2zn68C3GK1JzcHkZhxYWdn8cePQfYsWnbDatJxk3PMTxl
P7WUqMCqzAsneyHo0VHiQ4XXitJUn4lvxAMSVmidd0G48blKjw9dCfTWMsiD
iSwFX4AxCM2gyiQTplOBYtOlnqr45Gne/Tg0TNLoYAWBA56VBlcOKlh5/Y9s
0edsquhzC5hmb/9D0woDIDvRm/HzBz5Ghod1UYSosuEuq7JTTzm8wEVOmeuU
xGSarYQ0koDPRLFIKOW52JZJYZ3gmhGh6m6uQm3TcrPDzve8hUTIzlhoKgAv
PkIkBzDa5ja4ZcJRC4Qt4rKYIAYZHmGvtMwLRvhm8dgUXFGvOiLgs4Ghk8Wc
SaZ23MZX23noeeaIZ7k9BPtllwXrvJsu+TgPYOwPIHM3oSXKqaaYKBsU3EXh
hVN0MIPcCuIU7c1xHWq4/38HSM6Pl8iqCp94cbYYUYHqDWQ0IiUr68UQPEWl
P3QrDo25S5kAmr3vd159HUdzzK4ioe0HDtgqQTINvLUGsjJWvvhakbSfzfKM
ZsxoARVbaUmI3GDNxtPaSg1Pued7Z6zHT6Ec8977251mY5du3Yn7i5gcWvHU
0D55qoQHnv5YVg5cFF77qAr3kWjuYMDOVYrYVzqvrUS5KPmFZZrAuWtSz/uK
OioGclV/CP29xLAwlZQVGzUUPm67tRHB/9uZ0lvNyF99Z7nbrEuksXXia6mj
0dLBP8f/eCHNVVDfQv+fGaNKikLOabc2cbdCHvEoGEnz2e1Rhkzz9sxTxGua
WQ0iPVAhelUHv4DDzrtlIik4n0hKj207+mtgVujv/WvPolKuZq0eZMH/Zljc
ogckzmEpBQi5k6a3yxk/576gOJdMbThiNyZ3tKPfu53Jh7SdmJt0FWR/NSHi
puLyiQ4oCAZxJZXz+GdPZhglfTl2XiGxJfm+dqau9fucnkO2vUGYD32gHv5T
8w0dmFakqBMmzFui6S31w9DhKOVPDkEMIH/obn3xp/GE+Ag+QXmOkbZzyW14
PiWq/1hV7t3Mi+7ZPHbHDgYZ+M3mtxljElS5qn0CO7nOkO4wwbJigQfaxaXz
9HPXm4P4R54zW4DvQpPmrl1l3XdEk/q3lLcxeD68a0dWIJ6SYp1ACm5rjP+w
P05L+rsQ8Uxfpg58bAeXC4TElDrkgta4ey06GghfuxEhyIedMXLWECmfr0Y8
6Z0pqvGeYUhpdfKj6ZbJBQi492rKLDnjs88avpxVm+4uPx5c6YW/exBg+wvW
kiRaevjkZoWzEwTETUVI1Rz8sTG15hRcnDnab6Zl5Kk+K+BjzIZiDsaU1S90
+zGa2ErXNFjVBC31nuISWyck8Hij6646IiUwuMwLKTCsrXJE3SuV+s8EcdoY
nlBO0hhewAp+c2cTVKpV3v+YsRGuv+qhOV2ohQN9SuntZ0UfgKtZcBW3fY/0
OlfDZofQ+yOJ5PGEGCJmoWZbqVoQCzaC/5NLmmh+Dwh0ckxrvR7NTB1oGVU1
G300u73oggccpbpqnaeKHfXEXaxPLknPsFk0m89I2klQqQSCOkxCURgeryjr
y9q0GxBb0bDSo1tK2snMbQfocnxJLipKqzdN8DwD/hcqf5tHLZxNg5XpNVWR
TUzvjFRJRPlcbtI1JPkgV10mOoY1SyMkStDiaK+Jj/upEKWbNhknuRrfS8a1
MqLJjztS0bjSaZpemy6MZaAv7tdzkvL8RhgInLiH+p8du/g0lw8SGs85pyMg
1FurKZlB08iB1e+07pCtC8NOMQ5VFvgO4Wwkyj4YQwbt0XkTHvt0hDtM/cLf
cBsKuhhg2FWN7j+PmxVN74TDjA1vifDzZ9UeASUd7svcNshuvhoeAAFQGLTJ
uSDR9ap2SWSx6rRl847cHVAR0jRR56o3mUPZg9Vfwx1Dm4Y5qRNpN3FaSlf8
Awl4nD5JPyFShDhNr5AAXXB+driuMFGOOyu6hx+AZAmFUFzWt5lM2ir8Uew/
0EEJtZqHPf324VgvK9TJD3kNc+s9dv0kw7MDJbN32TrqiFDN07tikCeB20bv
0nrfu4JucVc2UShlHhR3gzE+JQNKNxOfZZPQAs67f1JosJewDuT8dieIMmp/
7pqaEQUpz7ivU1njGagBYoQWobAHa2xL/qJoxmGYYJGmlYDGObD6oxCMbcEh
LMqmGbg8G4+ADbESPDGWG1tNp89dnkUhlb7VwrcA04Lr4oaLZnfTMJQUmQXz
3hQS4T+30HskeGP3Uq60QfxVbO4muavbGPSf3zXgw5Ihwbk16GEucu+335u3
s5j8AR/ELwS3uaSIuxQWHTOSItjkbHbWUMOr/IpEeuoCK3sEmEPxA4Qgjemn
Bi1EQGKcLMYboJ3JVAfo6W0yEePJrC2wxke3og7B2nd6UjUZ03t3vclffGnO
s/MygFWAk3Aq2hlqCxXJ7sdjAU6boHo43RygJM4k7rKndsoEWIyV42z8CRzp
RCWgmq94wnVrcwPaLGntt/QNK+F4ovWbiBK7BgXqUAZsI5hVnFlrrAGi8J/I
riraLTO8m7Cy3g/QxH0gLd+50NoU410En3sLrdRh+JYRlA8x/gfei7fAelne
S8U4IY8oPkNH8/ga9QQeMSJZ03uKhBwrv65PfqABHH/zG0bFpct0n8OV1QTv
+M31K2fl2aioxuhCXzu33zWP9iNSWyhLp8rbxnrBVLBplMtnq6Wbt1yTIYmj
3avLdtVevWtDqi1ug/1IreLYLTu4ivNcvKnuue6l6TmWDlIbfwImQzZdiw02
0cdO3cekOgf4D76p69uoI3i5ZNxslu2arv6lVaYnW2+sLw5OUYjoi4U6O2Af
inf6jUwK3z75IrQY4YPMS0W3hKs6/1X7IJDVp9AJKmYTvpi21XxE/baOk9Qb
M0CFhfglEDhCMKI/+eOtzyrKHsvTYetd2sbG/fx+GU/Llx/2496vRg1t0YPR
6Z1UyD546tUpkMECdYTx1/yykKg1Iv/qWMQhBl5mutU/KJ1h1F3m/qQdYlPk
l1827YIvmvxTBtykkheIIWp7/ZZMqa6IXjfPFedz7Ej00XjswMZn7P6A3I58
pcebvBcQR5gMWy/7OWXPXhKV+OmyP9h2tMh6XCzp0Idna+u14LfpKzrHtM5E
BdLcZmDyChE7Cye0aVj+Jm8eB0Zm/aOnEpkm1wGLnHeSjMMft4fRCgLZJvMu
7oLNyLw2iHmMIGMkgF5ZI68ogQemGnUmeiArH+wD/2AcJAyeBnUvszamIMO0
YUJbnBM7YAnpCQi3R7xBTPhR+654hUxHbdjJd+2vodSpCf8UA686Dc8ZVOK6
CdPUAi11yZIReuM9AE7X6BWHE0Y2WVn3HFGoETXbyE2586h/EzFBI45ipmvn
Bx2ZoVu6w4yn0rj5qCIlEDoXRCIap47L8DH0Duz7eQc6TG3Y9L8OzxB0M01Y
APPlAf+UUcxbMh5E9DgGZbUc8HthoDW19CIwp8U+E9s2PyvHuvqajheibfv9
I0Q4MYgkfkRuLgX03dtBCWGofGsQr32FnMOrX/D2bn/FZG+fXJF/daRKxPpJ
M2nvfAFsvx7XI9Y7tIvs5pMAeEvY3XO+H4v3U8f23RjM1KvpAKxYlBpyQf2I
pcbPON+ByRLhuIyllnyDLru1VknPg1o6Bw8dewzvZGg+zhFMk5nImoTFJT/A
0Q+6CiABQT1eGnCOy79lREOoTcMzeEY2BA0c748P2cHHRFCQ91Aaj1kdkurJ
2rT4xmevoHfPT9fBVPFCWLvn0xOlJ9ZySylIXdA4PeBcdFSH1/nj0zmQmjal
7vKzfdy0ZG4t7Rq8su078GUnC+hgBf/v5TmIeLhO8IAF6MUV+fwaGg45hpQE
vn6UnU11yNt3ZMRWYdWfOn8/xrePvry0I1XlAFF/bcI5SU9RF54nyD2jfCkd
YTEJ+UlQH4ZnwbtbFw+z2Su5K+Tx8BgIznarIHBhejNJPP7ZPBW091ISoX7P
kwgMQjMFHFLg+N5fzVXBkqc6hZuhpq9YlbDNMUY8xkg5NsyG1/PWA12nbBXq
aR9GQGa9RBH7UWlaK1Jr2cr++5+8cMa+mTjDY1kGvvhhLofgw5T/3d+RfTfr
VbcF0q4GwPbHTI/Qq3LQZAwGbPkQQXYolrEdQHR2mzDwCq8oXO9XWyLYWP9z
grUN8sjXuiXn2VVutxoR3q5w8TK32QeGfysAjaEudhaw8HANqngO6db9q0hM
WWq/hS8oBHL4xWd4lv87vSzVrJHuKrVemWmEY0egh4Es8QuFDt8e6IpBTW4i
+2KTqWqq4bbdilwlHzeF652T6DoSZ4VHgJitPKP8Z2uEkVhfKQiiCVzi+tDW
4rz8Gb9byhjBjQssoLvbqlEZnVI1QM1QjJIyhUxI3QhxyR6F/zif9XDp5C6d
zCNyl26T3Tbi9jyLYhHIaob1mu2/YhK349xyGf4kIOIHSWnDESLbXlFhg9qH
6VzC10L2ww0dOb9V1r+BDG2yUvzgNUI7ogIwAHhlgNDhZ+PF1kuP1mguGF/N
L4YIVkBS6HIdIrBQKh+r8Vu2kKfnm2ZYAMbRkasonkvvyCgMTy75ngDWZgtb
GekXF7jJcIx6T2sOkD8FvYEkWrKcEHFwIPBoOQjSH1xAEOjdLmEZDFYkzQuD
052YsSwBEiyRHkXW6xGqS2Lq6fEzqg/JOPzZm2jklxcNtEQhe3umeHbfpJIu
385ly/VqZYIgMHMM5BPmNouL3gOfdy1KnC6znz2NSSMfJv0+UghbN2ERY7n1
Rv01f3NSZ1F+m6HTptuHBL/X4gZ7cZ0n22FV0r6MnLYKRrOn5LkvYDNNW3wT
MqILwhNN32ooLUFQE9VhjmXbO9+v2mW2zib+3r2FHxJya+slMWuf8wnBhNOZ
327XDlTm0k8udCDyD1WEfubzLiCArggdXObZFtHj2QvimZLSuht2M3+fttGv
hWvdrlCnwwKurJ4qrXl4jvpr1bObNVhcnP+nPLZLfYXzAx51KveMjRKMvkjA
di9z9y9oj+DbpYzFJpxpsb+KY5Y+qQQDdcelV5WL4EOlOzQrk/dDsJjrOBup
0wktkE86CeDm2AGykZJEpsVUnEl+aRdFnI0EQEGreyfoV8veSeMpMoQB7K+i
GmS+Es8fzsjjzW6UEjb5ZSmRwHaAaT3fijX1KHD9enjQRYGGdFTH4rjzPfhU
njIqh5XXCLrVGJN6M/6zq6ObKOGm2f/itpYsc/hZqHp0dFHS+M9VR7+YFWnR
RlwzwTh3x9paQTC3GJKKvAbNaB2BH2FDd6PBpv+6Y/b8CLj8RzLVV3OW0oHz
RPFZ23NZzB4TpnYnAin22/rXcvvVXHWvjYnt4HjTYdatkPWsGVRoDigdrBvF
wO6/pgU3KKsyaibYU4FoQn29LsWDQtflql3m11Af/PrNVu7gWlVFLlROV5p5
l6qBndiyIkgCJpB8R0I7sv2Ctn0kWgD1NsswIn8KkA4i4yTbGiF3yJNgLeQa
gx0PTj+853pIL5cLi1WQKmpQuWCr0kXx0IZTD+e8V5CdqF11R28l8zN/jbJk
WG1quMwCXaUbaakbO0N7EelTGhpt8h868PNU9GIBtAqtc/0B/dXdmTTD+L7X
i+2PehQv1qACliHwLsjLq205usaCGghAiuGOkVMI45p+UZEyu4xqgvicH7HW
TzdclcB5eb9iTf4pbgqZUrSqivqkKJEnj02J7C20ozgAWCedGyrz0bLYG/EH
BLWt32DwacBcgwfaz4HTKv2faqRMrVhOXTmdTodzM5APubvMEMbhBxqApLLy
A3r9KgAF+PPevmdGPyEdv4mi0gLVa2pec5Irsl2M/GmJGaFsDtt8fNgJyrqT
HTS5H5NgzeD0JUM81OA0nTN3m6cVqfL1S4+o6TyArRBgIZP665XQHVODjbMl
caPgIUdyjmqKyg6U4uGUQSIcOl6TKDMGIGwjzOjMCjAUtEdHaQnwJF0SrWZP
5gS6McV25txiraz952EhMKWIkIrt2hZRQQmYCB7kTg66br252PggzqgUa1qK
So9ASsfIfb8r9zlyAL7SYLcPQkGjbvVmEogPic2LXK/vi7vwI4Y54lxuKBbS
lw0aMpiIyPEyurxVBorKaBhcnH4fzeNuEdsONQIxAhEiAlXJ+dIJyuJaM8v3
NexGlpEmzQaJ0YyDRTU4z5LqNblLmT2C6JpuHURfy6nT/ZWh519vUo+XUTq5
CKxAmvi8qe9TgKnZ8S/xMHTw3bPkLyWkd4wPjCWh0DACQFf57WmG1aumDn5+
JbTnZmHyXUpjl3MQB1SbcLT9bwICIyjgh6HHTa771indKMrkEXEfFjdjY8a+
SfNFJhi8GGxIhxnbZyploVT8gImbJrThKG+D7dZWzTYG3DTNcDMNRWEtLhVX
klVw/Q4NSFsNWdnDkw4iIuXuSVE3dxpSwQpKY9v50KALR4p0yrX+4YizlKo/
fLk6zRrVa2qfMh4BBGBWrG6GxavwAYHfOWdQbR856jSC2iXxQ88zJ2AiiwZj
MByKdcN8e/NHj4zaBrSq0PcqYCIRC3/zFTl3rueD24Ly8ZJWVQJR07Y/bT/t
s8LPK21UjvB6/ei4y5TxP+Em3v+MjnWnDF2Zl4i+QnrUedTiQop0hC6+SYJi
Ewusq4jLOv9/x6TzOYEgaEwDmO7HsniDS3s+26WcA6zaE7epSOuPygYC/qg3
Xqo7BLFE0XTA+N/LMGrqFCHvwlG0niDsyA2x59VTesd3K/ksd8962itPlexb
hJwHE3/dCMUfL2polMMO/yUy2aNN9AR5ayHfSgeuXw/MbG4iGA8LMvCHPSuS
bplmVuYgsnUeDB+aGvorQXJhwWjqf4HARl5RyZBvBdfBU9Muna4wd9c6pGtC
0zSJUnW0IKKqEZcgJZdvKGG5uPGMYNVYsis+4jF+WZENr86/ONIufodmuWXt
TZ1XwAiA/Gsk/kF3FwSLpwQ1WsvebNuaJWazTnls3cRzoxNrby0EGomUHHTa
rBEn3UvDYx99S4jUgUACXj/skj2DPN7GAtIkCLG0g2B7rcx6mewV/N+q8Tli
qcafW8xtGgWztt6NfgqAUmBFEEiLpMJbiNdJcYZi6wpvNtzHnlpFTaMBA8Lj
Xb/6DvT7/ElH7GYxo4DMsfX634ZCwvj/moZLyUiD3OXvKNJFCtKOz+7KjqhU
ocJQ/7J8FdlUXLREAjORs44ESbUG7WZ8unLJMyzbeYVezVRkB06rjS3ou7A3
NgG2njyP2NiTBzNQC7LjU5NkG6a9kGMfwz/e/QrO+rp22JD1GJpju38n6NkL
JzzbrqjjaMoTefyYsKcibKoKQewnenUfeR6GDxKdIZlxGalpT6YPviH6T3W+
m7wtUxQSdvnqxg/wclhCDVm/x2LotoTt6SO2av6P5wzB3jEsET9dEEfqCs8W
DvIeFq+NADdjle1oudb6vCmBJNdJ+Zs2itKajxgf25e56pX7G6N8wa3LsWdR
buEXPBPzqHjL4gvJRmh8MQq6GY+mEIFSsYhNNSEcv1mCbD+0/q2nEwynWwXc
0SS79cQNc8YJtQ1qCuNuK+D1iU3yepDpYb/4C8U+sWv4jt8Zl5zZzpLnf39t
R9zzdgO16rwbhBCkM8Mk0yfdY7uZ8sK/4afVb2rMhrb3oEWhgmTlqM5uvpAY
seZwFwcjRYBso8gKS7L5GU1bsDThDWLYaKQRIxgVA1Mw2UVaDTsQFDCnM4eF
PNykp7yJQsS0C6sDFWH0q1/lCVxUOGPCFTM4xsFmwMROvZ009s9/3sMQ0uUr
svOZu/TYACJoLSiyP8cZVMe01wbsexrKAn3LBk+O5Hg0N4Y5r8o1luv6Ivbu
jcLLUtw8cuBmhhLw5Ggv6zQkA0yw2wyvkm4RFIhPfYWbXWr2MoEljdJ000td
do/KJjT1X17oCt1ird6XuvKQhLBA8ra+lIWx/T+KDSZzviFlk428KN0L2dZl
yvh5YNiRat3YF1xbgZp9IJsvL3p7nkIDkklhi4+D8cSx70E7Vn7IBsn4hTCC
ZOEcOR+7J1yMYftcK+1sIioivtrJ08jFGfd1aT27BCePHOhNiGFR5WG/klcA
5Ru4vkRgsnq7wJCn8GXe+iR63cndWgiw6APMujinIIcmLDrEOX8IGbXel8bV
LfZ8W/zrxWGUDepEqHRvghB1CQiI7mHVCNCKjgDt1CBx1z8FFirN3SBUWL9z
U0P0yC8ylDBvgm3Wx351NIUdsGrygcjo2d3vR/XygrFBGtMmA/+97Ga7AQcq
CJZW4j77MML7lsqt4oEFAWui0mMyGM5hZQu3zp0hbhUhnSAR8TsfKs0YUMfq
DieZu6wNebVr6cPQXTsOnZUM0hYm0UBubClfvfWyqnFRaUvj5ouQgrJrlAem
pI8z6KB+Yb2meNlPRboIm5fXIqqdJF7BrVvt79t9dVtFg1QIrmvjatxuHlvg
jrYNO8r1zVfwDOm53GjJ+R7r1+FnfoZz4CRhuAdlAdM+9WWuZ+MM8EXmyt4S
spkfC/ozMV1yiXMddD9VkUhL5sTQ7G4JwydQkVfb5gUNq8UvC3h5DEzyapqy
0QRnL1hmpjdKkIedAPeNcb9UW7eQ299W0WPFXQu2Sv4/BVSS0W81tOTE/63A
XvALfsiSfwRAr8QxLczhf0vJtOMETzH/tVbHFLhCHc2BmEvK2oChsKXPhSDL
ljNnKbXtF8XMdxKAiRrRpoHhsbpw7DbCiKcVV4TAAfF72iBiq4XKNkKptAlp
rYRSoTy3u3NJcDXSHK2cPzeZs457QCW+gHkQJuyUdCISCnUeFvP3bWf+YPzy
Z6OYE5gmasE3hkBaAetI954D6HX3S1aub5tyiqmgwlFnkmZEAk4YIr0IWCfD
eR7X0KrFjnYep/PGilCv1o/kZXlGNimGzPiG8uiUWEI745lFLdqm3Y402kkA
CkQ4PedS++8/XcSoU0IbLDc1ZtIb7Ply5YYHuy8t7u5W+o17T5v7IfumgYP1
zXpQyQtSQ32xpW5SVF1JWToAknXIW/+LRXgJWLbmQ0nmDdaB+VHqJGd/k6q9
EZsOxUXv7ts29ulPzVrIEXoLYmAsjyR/rh+z/nJ2LQWuQJJc1lP5uSy/xPWm
rwDmC2yFukq33KCc7cH3fA5Lm0o90IhJfx7fVfUVzxHSzg8lco/bultK+Tnq
ZBWzfWRYO+NAQWwgF4Sxr+S53YlZi/byGpj6hL6akynDAoaQz5A32iM6Im/Y
8NSXOh+3rRu1Dv53Om4wUqBTDe9MQO7z7+tg/B5/W7jjrdZxHaNUPzsjwXrj
aL9W/2uTJrmrPn7R4eWyaD/p3baSmzXdnD/NDd+yLBMSUXcPfcJ87MQiPPPt
CXfzTb5eIyXDIh2Fal6QSj1hsZaqaxL6/xixzCM9989kpSq0FE2neEDs0rPK
qiFOW5u6i9dEw4OCfk8Fkoqnzcs1/EvpoGZeOX2M264UJ+JvVJ0HsM1J2Zuy
nE2Yd0ZVheV4NNmXkqIWtduOdtRT1L8+btqq/vcMlqOMmIwaPfoPcg9cry3I
ChGp61m/rfHc0AMLA+MpM1JsQm72euujpJYHzeYdVWEj3dmJfxZDkYhEqEGU
eIl4h0zSrqVl3/Ak9hQL4HmH3PiZzZJRA3iY5XEAwDYY9AXuU2MNXcLuqnz4
5DegXQXyRGFOnFjc2bwH1unOaxta8BpVaERSdqGlxVTeMmjv6xmA3alxzyoa
FxvuinqCuybYzg3IJ6wj434v8THBT8FS4q4KkpdiMX64AxD1sYDa2dIr3O5Q
Fmx4hxJ+FsVzJiBKirJR18/XXirGRoOrVwIO9nS+E/G+VdIBBrT8G7JJibdf
gydqa+/6aPUNu9Y8DI88Ilhxr1grbGm2zR3eQM51Aywopm+oeDr1WhIuJqS9
ICT/2/BWG0DswqHK5oq8DwkicaKUQHm4SFJvalMBwkjqYVfJLRLBBiZ3JRtm
0fjsiaN4dozNnYaBZ7IQHIs9z6JbSJp65OP0V4rM7deJHQxS+QuUfVSzDDEW
PxTPJZZqKlSYNMWwrVancfpzoYPlHq/hHQLv+71Ah6C+t8AsmFYE94Fb//Gg
eDnFpdewtld1xK5xw1UEIDZ0DFWyNAUhfGwwa3q/fRP9W0hZEN/g1Paz9BDx
QDpH3c5+/nxMcLywIjF8ipp1ze5HuSuz9wffWz2ohpKxuIcj7T5gVh9OM1QY
JLfRFKGmyswOCk6yxM87kcnMI7CNGVQBoERkxEmjhNYeZw/h4Q9ZqTK8h6DZ
UT1ypSae979cFkX0iSszWAwJKlmxIEJKr+OMOqbrYDXFrwhhMKJWGqoPvPsr
UpwS3MGDcoUMSiPd6JJXnS0l9Vq6Cb3nhZoKn2Kt6yaWQuxKwvg0sakDzVGB
Izy2SzJFQmjVfLTo2yJzKT1HdokrU4lB0tpSCKwMSPVmTh7XrqFvvdrplMD8
b0zwcXenoMh/ah36k7iT/8jgQaGu7hNTR9w0XIlBVGMmn9jfPt8772pgqd5q
tckmPOFETIy/JmK13kAwDJQGHfUWbkYtvAWzRbjuwL6glT9MJUv06KfQtOCH
9FJbcNJP4giyX8ZhXy/hABFPAwVMpNgZ2K2NVnXMkH+yf6i5F9VPdJik0Vlm
NRKd/jdtAZouQT3cBYUNAyo4O4x7MgbcL8zTfrLlTDsYcG7au9pZFVgdwzEs
89vmgEMwcmcXVfpkOT12rPNgSdSqd3ENJ0rPufWr7XJCZs3LCpYgT4F3/LmG
orWWcirDTYCtIGfToZ9sC6z4zx9xbzmHuQWDALI0EDo9UEiYqSQNT9Xybus3
xbtoL5z9ZQiLjqbrVI3auJ+PBEZcIWhkoLex7g9tjLMAGfMPpWwqWeN/s6dD
eazwqtdZHixH/uSn+GsHeIYu/drOTo8mCn7U4oeYSoA7TNShgKq7utARBi1D
BIigaouq2m7Uogge/Yf0OzVOnVjHheLplnsiuQA99w1mu7+JYbY4p++4cyAC
aa3Fs07eB+cZg0fjMJfxx/opC+dr9Dot0DKzrPYGhfzmqwVbxHIrxnobEpV+
bROUWCYX6EliRCYOXp/MlK2/4aBp6I+cuJ+JDUi1G2xSIC+N6BDLgNW1jnyO
wwUAhh5SL2JSuxnuRxMMVxio+UOew8DUKJeBFn6/buBGy0S68mkJ4IdMLVWR
h5JNjawL8qhBC38npZdDnwhtN6ZARytWOJWC77jLaXvjV8VlZ/XGkfVj0vHG
7uUq4Ppgk2OShX18T/U3MRqZsXtEX69+A7Ymm9QYfGUEkrER1kLMXaf1JveV
yxxbfGr9yN2sjGKR32h1cmlFX1qo389CDeTdJIQVuthcuDdgXvhOIWa5sGS7
ANW15CpZZN20w8YTcXKKPVBN9feQQboBv3Ge+1HnPhMOeaPMQXuRq0Jc0x+J
PQ8rfp9ilUpJVURsPOnIEbFrSf09y1DWTDm+J84/CPuaRY1+z+1jy4m++Ea3
EyefUHVoNDQ461JLI/3UwcvT+g/1MT6Wm2WVNC9tGt15oqKH7W7zdlYIAV1r
mG7/8l47SElTe7StxUEiEICTzqqOCgu17c9Ufj1SuDRtjI0BDYP4NGeeVrMt
+hgrKYRvbluqdTF5yLJ0VxWx0s0012gRQ+jjo5CVjMwk+KPP3bJHxiglwvF5
4fX+fVvTOJvY5kjWYIh7PL0UAhEhnEe9FI4DafaY1C+FwHi1DIUGRHI1f0hU
76cTOvJPIR3kIbeYThHpUohHZ/1XZTrSY71Is1igliYx3b5V6C67RXwKfyxb
x7ERCEvyrsY8OUQuAWCctXcRXoxld3PVAmnft1gHPgHI1v+I18mIvRijL5K1
w1Jbn2A2HevJvCL8LnGEuVoOZqodmNkpbGMaXRiRCd3e8/zug/EJ1/0zPdCJ
Jfdx4obLGtCaP8EQID0IWU+P0XXD79zZd0nMiMzdH+6UiLRBp/FPZtDhAAPC
yifugZOd3N+bYdwcuEnN0vJDkBZzlynTI3ivQMwi/yCOqjTb6Z8D0sk/IcgH
DugzbyxWtAAuaH+6Uj0q8yt/7NEXo7WJM4p7jtcFCcES3FxoZ3lPXFspDpnj
6C+WGQ8Nx9nlYIs0li/wLoXDu4OayryriGv5HmYEdXDvNOeJ0/oK5B8ZjqLd
h8pud3mBHbfcIdelBc3SCCRWdsdZkwfGotlBIFlBGPq4nMy896VwsThZXIfp
JLvwUN+yqGz+QCHZ8O94OxN4up1s61vAyVFEAETksSwDJ8q9vBUUMxfYwsdX
Lqc6So0NQr9Ot138VUWcWxznOp3Yk1Z+ykV91VdXgg7RCJAWj1nDXn3IOcS6
U5V4tuRwARytMsGV0L9Gs4wtKIK426ngY9FfyY0RmAy9kpB8/dR6PyWM8U2C
ZB0CM1k2tyulDaX2euFDO4GCV0Lfe80/KosNL9/hS4pgpovvY0XOKE21h84J
U00kv/SblNindodBXJR1NlgyK0swkFfn8/ah7JKlg6f7ybwpMegQu3e+Bg00
krPrL6AOIgR7iWbqbIg8d+BhHkFyFqeqNHfLh00y9G8OizwlyWsq0urECD83
3YDWXVoGIznJyhunhtY2k2jCsAePHWIMSvh0pG6fnA5bh89vL0brYFSch2tE
Fi192JTYpRnSJFS52j2+hoWSKFn4zJIR96hmBB3OUk2w6H9POr5gHfJLi7yE
Le1Wc9i6PTDIcYkZZQXxgXUG+cTqW5v7hNO3XuClnyoQgzOXJJ85PNbVcUDo
D00pXoFcO/+ybEHMjfamTU7fkh5wqmLyY7oV5h32WxrpTTGXfNUbPFKQi/5V
Z3Pwq7lBqn0rzIVaQ+1Besu2ibELVzvmyBDHMKNdO3/hWQ/czQRkoGYNjYQ4
9CB8qNl+qyL5ws8lvHhmbjBkQsMirEuzW8SM5GHkCVjDoBDtzUEH3+RvBGUE
m82hTu3efOl7NMfNI2LmTKqz0mF6mG1vgnUE1CLoyBB7D7OpXlfWqF5Vihb7
CUhCQje5O7oLlUy6cStYhtJWSthYsswT0xs57GwblXRSTaLXTfOmDq3he6QT
GPGZL1JvonYJ8P3KAbWUO5zsuvtvTpO7hj0vwD5uCGiqjMaawFo1yVZe9jjd
IIs2cDk8TgrpX8is+N1oH6juZr66vAsYfkXX89/bjwfxHgnAm3qDnJVJ6AAT
vm5mB5xToYTNaD5FnEYw7D3efLSPh/2rEkKXeaXrgm3H1nLA6B/YEU7aAWJG
dz1x7FWqsHEjqDzG1cOPPWV2wvVdEb1CAg6azpVWZnghRj7F5z4bdpBj/nJi
wB+Z6aIc+EyIxjdcEb+2pRfGAJZQqZqHO+Untks82lZ18SqSSTQhDJyWCCFm
N52hb683y1r9NGsWUFUubjCuvNJ6LVz+73tiBxMC/H/ndUdBRdZ2g5dEyvTN
NZ/P9HZJV2DkC/Aj3Baw0Zqqo+WPJ+hOjvS4vSPZ7pqKZqBwaQ5rOLyXtmJE
unI069D07YBR1reVhNaaARZ5Ue3+6jq01jHsg4aYshgWszG6AVOjkCqbaUDG
9vZNZpXSUUPl96yrTaM1yQO4Aj3nYQGCuqXuf//gHWFwlXwJdxJJjQsom3E8
iDNcXdlzOIk2BK5RmmvNVghUbfQzzO13iMhhBpUyyA9auy/+xliNKkR6flx5
uHhKYWGxco799UXMJOmXo/roGU3vK9/sdH4CVHB4EXP1YwwbwszXGo7S96Bh
geBoV5ihGA3cY6/CAKjgyGa2kUNU3R8vyOSknIA13fK4ziBqpSO9lFngDNYd
F2qNgZ4niZbBFpoEDs8vQ2SF5Hr4mz9l6QqYLPG5ImfeP3zTNTlMBfaQzlf8
7kRy/mjzQgSa9/gOFk2+sOw6cTx6TnxfoNYZ2J+SvAmLuHfzvbjLYiGHKY+0
u4TgAAAe1Fr8PznT1J0OhDbTw62aqfco/Hr3pbYz8PPyAF3UulKAJ9+v0mlH
XEShp4j+bAmzGVXuJhActTlWhzRujrqVkgjQblBeoaCBoagSHMUcCJvxfvNM
ve+c9g2q/pcylmYLdFeqSNxhbR2tyz78QvOKMdpjQ3OyuGo1bJnIPn5iihiP
m4w3SLQyRx5YtJEBqo6Q8elrz/lbmwIAx1QCTQ7Cp9If72rQy7ilEgOcZeZH
wHXIV2vBGoyxG1hJOqNEmJy+ynJ5RGHSXR2YWcSHwd2SIYgsNfwoKeGINYs2
cEMjzJkZcS8LO8WGfN47m05vx1McdsiQx6LGYk/yJNB2UnP/SptLw9q25ZPY
Ba/M0YR2ODMuTDOFpToza7U163zI0nILEGkomYuziarzss9+J8NO/A94I1d/
e9OKB+ErvkCetYrD5LJL88kbiRhNaKy9Tckkr8Vb0vhxh4Mb/3l/gi/7PCRf
4C+pNYju1NkyuL4X1aqrh1FzuPde0NK4l4GunA7mC4AeOnvheJYZvj3dPPhZ
g3IE+JoMltgEBMCFEQyVdgtTuOpsdL65AGY5uNj8GrNN6LfLi7K3SfTkuk+s
xRWfBrgLkCl9hUJU9bPzyzQ6xuTIuwxv88vY0hor7JcqBdn6JDYWqa5amenm
HhS/Iauv7joCPIGs47uAXOyHaWdQ4nbrubYWVPUxooTqzXBTLkWGb4hzxHKE
inftrp2YD6rN9OGOORlppYzEh2r5JsT8h7RbCqcXrvDrRjPIHPgkrr7HUKhl
yDBSEqv9MrsFJhM8CJadgsKOtwFAk7XWjmTqN0FlFiud8sFhZJqmtc/Ku7mq
K1VduKKCnaTWy1qfFKasz1+epWtPtChOopFmi3RbpVs1dW0aZzrw8DmmZaZP
VXeSFi67Ys+PkT0BaRKzVR1UqwjpZqC0sVjM88dkyjjBNo9yvvqXFESEaqYd
bwDh/3JlQBNQhZBllC7W+uJE2r6sCIKh7gdENLWwMWa0h1BeEYW2HQ+rukcE
zVGpiZLtnDcmHTsLiiia7rX9sYMfvXAOeetRXWca4XOImudXWKsgQvbzWmZE
TZs26C3BYcA/arnbd7Ublv/kyPOuOmfdydwhmoV8NVZM4NF91/XoZWgKCvgE
6lUCryOPi9IkRteK0z7m541TuzLUZHg18gvVvP71Lf/k28oiYVT65V+JMlWn
970Ir0qJmWovi/wmmlR06VdlKROUoOZUciG5qe0CRdlw/dAEY3bEVDE/xO6J
9Sbua8gFWnS3lQ9SI5Joa4sHJu+pGfBLMcix5sZQEIZcXRZOHM2FIFv5zB5d
gIeO7KwAEtpScAfv2jkDhfBTHXxw/pzr8Y6HuBiFtHATdgR7sk9Vnrqeai8Y
9+aWBis/RyP7i0QNnOF/aaKoaPSUrOdqC7GBae6c0fiKUFKx06T60qYLPWPV
tzJYZqfTtDPiK1OiD7EgbY64atueHBJMhJD+XunYNxQjSusPLuzxbx2OOzRB
ER7mRk4TF/QG0aMxoxKJdutBrxt6p5i70sTl7Ijou8AUU6+bOp8E1jiYkyRu
koSm1KnIArxxin1QJ46zw7iKQv69Y3ZTpODIS7oDkA5pLxOw9/rMbe59uFc2
u6YjNV9dxxTZm/j8LEhZDLsbZks3JSjsIn0IAEzoj6hSxOfwMXK8aCe0LTFJ
fj0EQuGNoI4KOsY0RN0rVGwMz1awm5EVkbgTZ4TaclTOgKImBh2F87/4LjWG
72QWI9N9ZmLdAA3Rt0pgbLvGUYKiEzx6I9m2x4Wr16VHOymdUAtyQkQwNkBo
0jNgcLRxsGNl3umOhLJeW8NoQ6J67Y2InqAl/Hkwv0L144hRAz4jbAmfnK2s
c8L7syMeFm+qxYw7R95QBNIVAyZcUfmLuu52bNixC7fKpPjMEF9GPaEbL+JN
pu5V7BMr6UQYHug60IPbb8adO2TqznF73XD5XDAt6c0nPlkKWjRp7uoQFuJe
RMaLGGOB0MEqU6LSjsx/mSjIKEP4EFpyIIc1eoIJGWIYcuHX8Z75WrTva1tV
yJEX6LTcnq82Ak8tJqKq2L4Lc15qbKtG7CTtBVXHtmZXXZCoM/JCFWLCx1Lf
jG/f/J4zMPIp62VgRjMpiOXzoV6hKh9bIyjmnLGiEcMf1zHkK+S7xVkPAb0r
oB3lS9YzL2b5z803rjIBHlF3Z2YjDp/mOq4g7iBW6z+sxXG2TTe9XTmMH1FM
/7//pJ5zDYB+J1vb1RcE47HEGD/mN+gNPS97B/Lt625xXKXb6qFCRrChzyEZ
mqgRIsa2WerlfUbpAlAFPiiTgREAnJJxydYneX6s5VWp1haLXLKGS+Nv8CrZ
RMZW93C9QBy1BONDWTwuEVko51pgTkHJ1VAZYc61uBL8lZ/ld8aCVM2oMdbi
6UaqyPICXjRPQCt3olTdRD9kOTsOfxNHEpFc10XmJ+29FmCfIRKYZlcrJj4F
IEyVULA1AEZ7MTbSCFaZnq5vsAv9l8eFzjBbyFGnPtmMeNlyKT9fcnp+/8wH
Bvkt/zrtV8lLQM08ICQurZLsShKeAtEYWGLBM6f1Qhtkh/YieiTvdi3ZQmVU
Rtug7gpeDw24+culggQOGOk2jsC0Gl/yEMh2rXbb9e1oSr1apY3B9K2efobJ
nokO7ou/R0dNCDIK9ckwZEcgERqS6ViWI1eRTkbTleg6gSxWVIHSTM/iM6qg
mC1oNnU0oqerxOdPd16O0lMCgqHRlzzX7l4Ry1CBVnXmSciSwPxkCc9bqSYw
dzNWMc/8KA52ewBghu1B6snMIUCLgdgO6E2Y6jHCrB4wwFiuvdHl/cGV/7wi
wDoOR0RSp6ZtRTdhF2wkHnkvGFW1xd3lkf8pKwe5CNsy7PLc+mLZgb7EMeip
mwgBerKmevM3ssK5x/SwJ3JY5sLIR5cw6c4r/lupEYPzOaSGpTFirpVAbU+i
M8DXHCRBl70YzBnr4CtSy1TVWnsDeIqhbyLmZcyxP+GeEVS7liQW22+2nwyY
XNcQxHD44Agu1l1fpA8gaCCHdD3yPpD2jQTVVSwUHw3Nm82ZPffTcf/VGrPj
MAzGB2VSEi0CMPNbu60RXZiQ+I0hRqFsIkXCRUMT1qrbM9gAGwcVp+ZUW0Iz
LOAc3Zw9o7mXcSg5Uxxf5lZdXUGlEmk3EbTx+Q1hhLaFost7WgerSBZI8ywy
/L+TLSGY7I68r1mFo9rZSbcHfZRWVpsVlJh8eT8xalKWTrDB1iCqdJzr8PnA
zcgzoBjgjMMdw4mRsGTsfu1GJSuCj0QVNRW4Jz0CgO0rZvdtGjkjva21a9v0
d9Ihv/R93Et4++OuYWFRykgp45bL70Isxx/1VdT/l5tGN+S6iGiRuNomAipf
gu6JejVHIj/slMHPh2mrWwGSEnd/DgRlX3uMu1ysU7joW0d/KOX38hfnkj3Y
/BhTunMwHBJn3RVfBUK9yH0rC6KKp2MOQ5OWmupk9iYPcugmOOgYT9s9ZXWw
iQkXpCLwiyrsgi8hths5QsrvD/ahtQcVzVOxNXJfjvK5FZcJgKrsSDRU6N/z
YjMZZf1xel2MdoarlOX44PCcbijHmAZdUOX5TrpvwRMaEonuhfjRX4zHZP4D
pw7ICGCTmGetDFZQFsaCDnUyWM4IGRhmmgMuzD/My+di0Dnu0JyZ6RAUAZ/h
q+gDDx8jWU8qk4PNMN9m2d0T9rjvllqN7KCF4QKsnZqlUwrTJ76zj+VZNhQ+
RIQ7owLzj4Gh9eODVcwtLc8/kr+jNVACzVKhg4Gxb2d37+cxIHx1F8XHDIdq
x/zfIBcZmeUAgplTpvG8lqOHMQa4ymlpO9fTIjurTpWf0/SXmp+ohgcFrskn
12cquxMetR1nuvjOxXgNJkPMbeQBjrUChat1MZWgj0tDg0gRLfDq2+6Zbfjg
YyE1zaKbp+XBCqjuo1WXhJyMFe7H2AI4M4hofwB1gdm6nvc+TTrKqvg76UVg
RX5zrnLObY+KFlzlIQjVf6uZaEFUImBGiEaF20is8m5dyEvOjAhKhDsDJzeS
y8IM+3AOw/zVjQ6sFSROlRrkvJ71ij/jPYKCFHDcdCKdFeAgl4QtvQKRBaYa
2EuriHV6kZPn+4+ftymaMZAqszuHkYbyrtygYz6OIFPiSIB9j26AMeGcPfhm
V6J6rgJ1Ubzxb1alow3rsr9cLzwfiRsoUtrhgU4XFTxsxgXBhNR9QV1uEnoB
yl6BbmdLFsaWBq3cyMgX28iLA81r0zvWqC44LosQMBh7mZflDx0MfycMW25d
Tbiq28oe+ibU2MaigBQxKNtyoTLPUFJN8ZgoakpKmmQLH3UWnPwdvju40jBm
tt/Rx3ItlyX7bktgpNpdt/6vBxnbM+DrLqRwCTNtxzrrx42cxXLdFJt1H0Nw
Hihz/7CIehICtAxXw9jPrhgzKE8ysM3HTcPLGocZPZH2k0JGhX/67K9WXkqt
qWk2EcRo/nRaeWlJEovP3ipfGAhX0gV6zuKPS7Z6sKk3sUB7n9asNPU4ObgB
53vWo1XjJTDSF4aIqSufn+7BhpBTAwMuhAHen5KeYoXX78WpftGl45TVPqz3
+fHhuKI6e4xSnt39Sj11nHkVpqtn/47Od1DWKWPGD54dlCvqTrDvvqjB4Vob
RAXjpazfUD/quvg/ffHJbAgRisVZ37xEBYAuBchdIltuIvVLFHjx2/B/OalR
gCNsIlB1K14qAhzCYoBuoG00Me3jK7/DmuQ2QMI50KMSJYY0s9tOx9qN2kK/
vyq+KDLWdRg9IGjYWRU06J0IaLQOmq2jacx4RQAnsdUq/HhlT/3wf2SOQN0G
00HK8kwSjks76gFB+FoGJHc4XtB7/VgG7uPpZUo9fXnTMkKwCzeBMeKhlRVB
G6mKZWUnNQotIBTw4XH32jyiV5eJdNyrY3mCGaCxMdpC4H5s8nK7vGtWbzVE
oZikEDq70vacvNgt9/VgUTnFmPLQCryJJCpea7CgnbdXdig167HWbpip1n8V
uA1epYdFDNaHfNw7b5rDomQ/PlxqOVRwjTygDOI610mbbdYYreIO7k2/1dTd
sR0HIbz4sUS0WxfJhkVeQiJMyoxzOxjZNNijopOQ6jEico3p+X515IEuvds8
O5NX+33a6WaF1uQ0/1ytS11mYjyIuk+qmcGm3IOomvyxiVhi5tZCUYDl11P3
TGNreXIt1j8+yeD7CyTAjt6UrwL6sLk/3nIGHHgccz+H8K1oVaCN8dwqYt+c
fTPolltVCIlDiIxELOoe574AttDLv0fvhxHgkbZQcjoGpWxq3KsCd7dyRnzk
2uP6Glh0NFG2TRSXChENJQ0IqXAwqo2JntKx38khiPXmYwTd1Xxn+D1lnB0y
WfMC9fwXU6Lr4JyP2Ewa2Zl8nfAG/Xs2V3MSHGkIP1MqTxwXieFsuDDxBT2v
3WDEk78ty9pGSiPtWjPUgQcZrudNr4qjcXqT/gpQxfZz/Fv2dGe8Dobbq/l1
UBB2gOxqBOhk3HxuqRiuGkT/9vt7Wr5TFEVaNw/g7v+xwNkgHnK2g+6QkiYf
RSVIROMrDi+YJRRnTyJDgYPYxpEzyss1OsMrWWGk0wt772UtJ+Kz1oCdY8Mm
4pPrEL+R+3x9c/Q8j099LoqUoADL7pTMZeMLDOkV8viGkYOYHEpx4XSsBJ+P
Sa+9IeVoS1NT9EBRc7pHuEXZDvUsz8xgzcWlQ3VNnC+KNUZ1hAIqfvisIBks
F87ILT1nhP0eH2XI6AYm4qsTQdJ3XmbP5eeF/1upBh6Vy9PjDVWjTLCREW49
CUUlJo4CTHIDNXLBVImjz/nb52XJizNs+SUd2K/EdBYNScM/vCGZjDPqzwTH
pKCarfTfuKtqNfQI/M6H7uWd53y70CsNHC/e6vnnuMw5MSbiFsA7iO/DB7vO
mFzW1uQwfoAlI++SN8o1o/DTsUyoYzZc/ul89+4env8jdy4v//fA8+9rUx3O
pLRko/EJ39wPWLLQKKW48JgT1q78ve9qt1DdeEmbl65nBcN3sskc8C1p2Kyj
nwSogfLRS5aYQCRSe/avnjQ7obM9Rign+VaIkhuF4yEuMB6fAFGtyJLtIlGW
Pl9sfk+S+wE1wrMFq6L0uo9fynIgJ0OuOIXmdXYjT0PAZjcZPisqhTDdfOBp
Jp43HTgIT8RuZvP7ixxboFrG2dV0uhWpgDtpz7NePlrqr5E8vJmfPmaAhEn5
meeFFz/2hGKd0vdtiAy/VJf6ohdyOln0bDeJAqPM/6IskFlI6nVix37mKYtq
rUXhHvRsDeHl8cwAbRJYMpAtjjN8I8CjlmnEqCn0NbDXj6sLyJmcea35V4Ze
mKYWRS3GibJJLIKj6IatY2yTkuvHYMkTl0669tkTrOGmnhdbCfo6bdqkuTfp
CSS7T5evxOYYPzeHaa68BkN+5uGn7zDKfoYiOAYdeSXg4gz1WaWhyKifsByJ
si+dLnPH1PLdjKiGM/pvErS7JOCPqN14U09EMZ0L9CXqYRCQWzRg5ZE3Nqr0
cTo7euqynvZDmbNj/oyXHSMgHWG6sr5f+cSfYRj1jTZvW02rT8/s1n19Bqt/
SEQXBDngmVkrOq7+h4OiaNwyivn5f9WVX2fxCiHLnLq7ORDgaAh+0hxfOlyK
A93G9/PBswbsJQyRhBWBNxPK3vFOzr0VWpvbgYBIVmC4J0Y5eb5/sYZyytAU
RTUTw5dhhHdVLOdxlAZMUqcWk2snYwzrJj88pauPSt5yGejzeh5r2kx22SmU
vD1f+yoItBAZ3Yr8GEo3SiAqL3GxIi5Iy9xOc6j+N3hLIop2Vqv1ojgnPu1k
DnI+rONY4YqEdk1SENcj36IdvmCQ6hViOmfNP33IKwdOm7cDJsAcYCCGlSio
ta7PIMJ/sPwFBC47JU5faTK1wAoMoRNJR/X+aCeyC8OUsl4mrGja3KWwGuSG
k89uFRO/ajdLTFQSdQDY8wZMVIrDNC1yn8UIrwWT8hzBXHC2jZIwKTYK5Bz7
Ycqwj+32s/wQWBKfZ2jJQDzXvffNs8eESaM2WZ03vpkBTTfOGx/88iYMnvkI
9kFFzr1Hr8Ml5RAG1rRNXuRxRiUQMDATuofyxDVUhUUByhXMHKoJGCmjQvIU
nG0bzKWOT6AGoD7FpZbzw7tUZO27OK50+VVbvbVdUkGqkSucxVeN/em4D8Uu
uvFr8NYJ1sb0AEiT9FoKuGDk9OEFKSWUqXrNPhOm3wfk7ny5oxvMMmGdxOUQ
6PtFDUjPx4NyATSr8HPHKN8vajB2SNAUNZP9FwCMThavFjFJjiIeAqdktOMj
s1uxfQ9dWP1zaQL4JwHuG+tDQdWQhSfSKMKIDv7jdRErqTXSdWpViH+WQBwE
VSXI4CmVJ5rT9U72jd9edisUC1xKwJfxSDMI312dNNUlMb2QVUSX+XazSkfR
LUXasyBvXcRmIjDOrX5O4prM8aH3DJSDIwxoCZ2Nc5ElH1dbGfRSUIbCWTX/
N1rdcHh3FGqCubrG1oot16hk+IBBOlgZhivDl0lyZfpagPV+tnLKIKvOfOn4
qR61JIl4QIl6NDX0yTX5VDRu8za7w2fjW3ir+hptvwlDE4L0eGhvrNBvWIyx
5oEe3gmlukg8CKQTIttQ1N6bjEupQyXzbx9Bw0vqaNXnt7wBHdHX9WD8Y633
2ZEjminKIsxbOx8hK64GRt39KbYDGkqGU/RBRgl3Wd7/+UBNDiSUplhTPwCf
gFyYmAvD7f1YdK4dpEtZHxqlG35UPXg7pvNNu2xTRjhCMeeQOP4sSZEvpe9v
stej7WlP5Q3OwOR4qzl1lVynxYUaMT9lMhmnX/qCuB4jzHkHW8C7uD35shGL
7tyq6Vy7p3c8Wp5CVsG10dg3SeLigPj+DQeI4u2YOxdokpBEn/4Vwj6uMAVF
DBL6vsvJAsRekxbO5SmgUrEy7zYe7EVUNuRiC97QwDMeMbdzfvulw+hUiA3i
lPSQur4TId2ECjC8rYlANv1TcbT8mJebZ0tIX/4eXomqi2tAVmavaodM68Jm
GS6J5R/NMTGubNIwo6C8/hA9JXNajDYMqIdES0iPXl86FBVH6u8SoLYGUa2B
veENr7OFnIC7cDFRa7/HJVuhMM1PztcKVrVit8yJoCYglKiFVC37JXD0kFHL
14eMa0sX0PqsXlfFkiRK53yl/gAfzHaMpkNcSRnh9CNC1kH249dMdzVUp1MJ
rC81ptxNR9N9qSHa4k/D82Znj3Guoh1DzbGWMN/Q+Aym6zYwY/PJD1wdhjVM
QzzZfWrQ7gXSnfv/cD4bed6ZVL5ByvAw+GjmvbphkKNLyJ2KnEvIL/AS8YA7
UjfEpl1wDV+B24b5r9NzKtiUR1yDs5mXcP6oC5JsvGDPxSpptoinBXUSwCpx
9czOqUg1T1fwL58FrbmwQ2sEbyB3PpcCwtv0l1Go812yzn0bPuOXPo2qukuy
ycon8pS590gqnSbo6MZwUZsr2VE+nigYBHQWGOwueLEeOpGErlPA+ZmcGe5T
/aiKwEkgnaOjSbIl9+Z3u23V6NxcdapmJOxM3Dsvj/XS3rylH3rGDNhxZs/R
d3Y7IEBfFJHZIn0O3bJLbhoamHwz019jYA08FQHokywZvkAXf5AsFvWYIovI
j0sIwANI5nolNGPMnlixeoftN12VomXjiB3vl16ETeR6RN6g1nvcK253QsDf
1d2kxw49OCbvoo23Q+RgLdx9ub3+t7tek1tkeir7mH73fEyAK9nxeQSa4EuR
lvVLFKowP9bpIAGd0rM8xdeKsE6qtQcDyeqSQkqKtP8AB6No/3h21p8uLSS4
SVMbE9Jn6R2UZZ26cESTEIV7479JF5N07vKhT/EcowLSPdBrA2R0e6AB5Kkf
VmI4woVY19jBHhmFJ0d0S1YR5QMrK951hWyhT0Cu2D3EPO/zdG+X0UfxtHtw
foz/pKicXKffrBV7nVq96GXCwGlax1YZqj0oL9Rjy9MxWmhUl6qKQcvUz56x
NC/35xX/7Mv8SwvbrH6U1EsVGuv8Bx3R3mK87pgYOwJQhKeuwsHoFLbG6n4y
a2wd6IOGLV3ix1hPdzSYs9GOAMwu2+Anr+o5WNWn0tudXUhxLNPW9c2by1nG
zjZv61UxWT/KmTGk36wRRThId1JF6gbpkCzT3nQxRT42zbXYnBSw90IH77pQ
f2h6RW2nFGiNgq4Sb8e0machYO6q+oB2Tb0Fy8U57nj+Tm/i6GuRaqrt3vRL
CSs/1+e/O6gW2pY+OC9SAsw6ys88ETWuS3ZYtfLNLKgWNyidrduIc1AuLfwj
VqQgh+trWmzggbyXKGnNYtgZpancfrL+EHQePDAs/wDAnTBdyKgkSgOrIdOA
ezHqpYCTTKb8QUSCUwYql50ntmnl5D7ws242tL+PyLm8DcWgojqeVanmoQ1Y
YeU/aQoG2dqJuJmDZcOGf+DLTYfguPUDW+qkRaWB745U/HaXAu4Bm7CovjGv
X3XzkjQ8lXCM2YCWw42Tj80AkJ20wYNmwGJ55Tj5z0eKYFdg5knW01gsWmjg
zYU+9DMO5OD7q0vpxvFZSGVzt3/uAFNTVUq2NDZdMkey6Qd1D0hG2LdepIjA
/sqIKsoDHontL6gv++awjxRGGPhajZxTyOcHH5IMAxTRmWmtYxE7UMg+pv+/
9ObHYUkJtOSvDPjFQa4C5xF9LLtqtt1rQCGHH+6i5KKutOK2f5fRhBrMJQt1
wbmtv7akFRp23SfQnMlCqpQI2g+QgdYEzALtu23wELhJpVsR/U189+H2XLN/
cA3IhaWJllO7o9av4BRv8FIVdzzQnKlR0jgHbS6tYekm13i0TriDGDacncDJ
wW4WKLJJ8BdVJYQRd3jlvOVeMb6qOp6VTYmDSOFJfsqHyLv4a2dBkbraZ0Vv
EK3gAzG5U/c+Px2y2a9ZzGji3VkaCrHBD9PFb1UbCEREj+7lLzlIOyegQS2v
IjYuDLG6sPllEd6TOkqS5+EBWh1Gi38WoK0nNQ4PRxjog6lu8h+uBuGwReDg
xB/hhBaxJ941vnvZvtRgPitQhxAWa8icT3yVUNnKbmozfpX0X6HvUtgQv1u6
OpUU0alzgR47Fbow46vdRQMnbdWNhsJja+g++ciscGJSJeegSiZ4WlzrM/Ql
POSb4iTsVu8B3aawQzd9bkshXJ9s5BVXFnerqKjHXH43UV33PR8keJumqrBx
kSqo4XD71BVVpyUmssmDLtdW0y70imtPYjsXTVAOcLgL/Cx+mtmXl0J666pu
5BTyrmfQed2NINWFnyi49hvjYqFdtR4H24nwwAWP/9vUtUXM4tSLPLAh52d9
JYyH85ooK48LiVBHw/M5DecLtzh0Ykp00LJq58ha/tNzlEotrx+V/ufbT9pi
XBAHDGVvqNM9O0UxveNa3766a5E+iTGV0GH93K6qGgXJMPfhdhV7n8SSEFGe
vBQrT3460aYCEZ5Wx2/cIAG74Cwt7RGHqMsF9Lgtyvj4WeayzXOQswU6ZxgP
jV5aUk2SzN/3I3KbHdelXD67TmgLCaOwtjQzncs74I7SutW8hx3mH2zECdfQ
RKAv9sUInFasLMOSkW8P9FZtgU2eOLELAOBKnwmaKW6K8OJiogMklsZHorne
OqXtPSDFWxHm5tYLbT8VXHJ8ySxw/ehq5atDWLV/qw5yw7DGhrchnNRoOjyN
orYAj1ypF4qRtlL4MAAVj5B8+PdJ4hXWp+WXFLovHku1qWB6JR1JHQPOk0np
ymtoxejHZIDBUOprav0P2BfD+hZ5HrmG6CF5JPU3bdvIsxtkHWShFa4P3og4
wQ7oW3/dXIUuKjpXRUS3zlM4dKnMxeujXoghRexQ392Fc4zB5jNQdByPRMzM
FPdXcsDPxI5w0b++GVXhv4powcUPgexMfbNwLwmbIHVGv+57u03k+KjcIlup
+d2Jashvq9N9hEyzxqR6pCnsvRzgK34S2StpN2FI93Glo3iFVeid8NY+bK/1
eWtlVy7O9WbL9UPVqymLPTaJRIOTBMvb5Fw49t62bEUHFimYrjpSFvHcqjnn
ppHPUjEfL7sGTZUD9nRaHQv8fsRh/1WLMYd2ns97WtB4s33XL9exHkBbJlWf
KuCmMk0lgu2nlemkbz+aYfg9BnNvFRmz2O+fGoXiH8FtZhxFc35piTJVkW9m
mA4Lsi84Ag/ej95EjMOFBcrvAVt9hUJ7sf4aY3rPGLVja3duWUK1icIJLt9S
SmU7fvvl5eloS8T54fZIAwM0u3LYS0VWeedXJ+r2zXxR31vq2tmilD7o1Ymf
6LvEMXSZb4OFTpWuH4ibIUD6L5FKzbE8k9ALoE0/duxSYp9DZ758qt/qluuU
Z36TFyC37eXcyYFldCT710ccGAgAfi23eJYQE4H9Nb1tzjNtiFYf1iEJ6AKV
/sjGm5bfjaBCNKPHz14KYuGiVy7PTxuYa7Rn8R/kWFU6O8vtO9XCQE0LYoq7
bJeqa5PTl4dDRvDZO1S0BhdVsXCnMCS1g+y/FjI14eIityQCRkGFGWiHD4RJ
mMeU0d858iX6iJUV5YEkoLh/fWn/nYeq9QoO6WsyxPOVpcFVm+fOU1L3uHzn
jTp0r5kXr7KTWr6AwDnkxICsxxbMfqcdgw+7t5vdoVxdQrBa+B8X7EGOUCE2
v5zy8GtBneKYirwvaJ8jOGmRc67ti1bts5UB1PIFV07HpdVTrdGcr95n7Edt
/pmPQRHlcE6YLiEG8h/mtMLk6Vp9YGifcSL5jHRuDtah9LN33fDJEeiANPG7
AuK6hlxb6Vyd9rmdQ4sVKq8ZomU2GqSnXfx6SwYE0iXeIqOCxBApuamGOiTx
/330kjRyxfX4Ea3cfOMyjTy4WSMllh55ls0vrL6HRvfXPbPEYYl16PiwysgD
1tEM1Nes8d+5lHKKGAsTBnv6ZcTJhfY13k+ROumFMPfd1QZeId+rfHcah4SO
Sbt0uAX2VmLkobSK4j/f1JhCfbL7ST6ZTUDXHtwBD9KaznwhK5kFQbC+I+jG
5buldu+QeDVv5Rp/b4e8D2uMARFmLU0156LbtcnAfIhHAXQ+1UDMtoU58+A4
VAJVX7P9bLO2KAdY5lf29EO26aLRqdl8XMZyedjZydGtjHph1o7rkzibKDhE
ZHXZvlaUzZYTV8Syn2y4qD/pKvjgfEUM9BDCMx3U+Ff7TcjAz10L8pQqHsWf
tEb/PeLJEWw8Zy9i1uQ+SQocoehxaF+Ll5S/5E8m2xq7HdpnRox1HWKrdFhq
AJLVH0lb2sG4XNeas0bWTDQYagauK61Z64/JA8xrEDTIMT7+32BOjF17AmGx
H2YY4kRrat6cl5/s49X30DNTxjTD+ND6HXAzLxjZau2UOIA/XtbrwR9/MWGh
QTfYmi2sB46fodt6tZp2Qe4XGNI9Lfn8akmZTcSSXIcTa60JA8RHhp4FCYro
+8hGH+92mvysSFv/3uMQz7JONlJvy/5id+JNyq+XqtLurpZJBZL+B3XInlAq
TWGJHu/tpB/AnMOaM077zV8k4ZpeNqcngP2pQsNq5ej6noY8iRefsYmnTazr
8Y05kRY9+zLqVbhffKJTia9S+WTJXDKgdC/0spmO9X3EqooreZS4Z+dShGbQ
anV6Sdps3eNRcHYmK9i4ZhDJ/MAPXy7bWVU23iUgn3wNp7ZycbXkvaBmpF69
Z7qVVoSPpsbkMfI3X4d+rxVofQEAda5hA/ZqKnRBSca9+NJIgL4zj24vfj17
OHgU5AMKLTHgSbhiy6dChqsq8sknmm1VdWFvvtbtg9pdvo5A5DLk94X3eWGW
zkb++lPB4IxWTgKekm9Z/kjapIyP+VHhl/kue/xa74XVcKhL1G+I0d1tWesw
a84ZQNdqKd9BU2ilM9fZ+qjAuexaRVk96bNsP2n1ZDc0lLskQ+z+8cQTOpOi
wJtVzJsARxQ/IAJjFT8RSeAEoDPWKZyPEydazE1VMYoEjMHl8d7yL0BCpUyW
QgDfjkNl0Cn3swklvqORO98EWCYK5hlcQxDHP94mbYhnN6W+2WKnH8wIh2nv
36mts38DgHzcJEDN0TtM4TN/zLmf7ksT7WWcLMjs4FDogPh53Zd/f6Zmobik
O/OMYOHre2gtZvsrjk72kDmvKLj41yDtLUVZkr/nhBScHyifZAhfR3E2uH06
38t+TUujaxGuH6M+PgoM0GMRIbDTBw9b78nF8DkaNQ+NxMOsPX697ycZwNy8
X+RiT++PVhiLhELM8owvVu+9NPyWW4+ekR49Hc78gBnRhnayCRAr/B2/+fbV
3XP9+Th1UvksD+2qh09fMul+QOg24KI8nFXO2NiSuRZmKA9F4YpXL89mpv3u
kcqzhsOYN4/CwhGfxWMbl1tRFNEJPdfdvcwRlcjxBcxMSOgGnJ1f8SSHSoZm
5F9d6/DcWLhed/Rh/DHq6gBiKvBig6wwFtbB/Ge/rgThmifsGtVjXBmj1CxB
ZL4HEko3GZ7Ml03kbndW5Z9j+kO6LW+koUgTaovLrnFA0wANSvgJlk4az1uY
AgvtiODEsV914Yw0Iv40cTNOEb3Z87Wj6t/hxO7acNZ8rB6P+ra7uokC3hku
WphmTSReMd0ACIyB7I23Any7wiBgnMKz7BL/jTZIbb+Wew//FyLRscvJ10PA
ryyQIsYj7anHPpoWU1GYBP2V9zstsniX5xAMpWzqSuu30W7pYxFGcKZAe+d3
WIu63WxjA6hRQkjace+LB6JtMHs1q4TmkcdHGqJ23Y2XEkshT0hR881gkb1P
AFeYyfoql2lYv9EPhxM2NcpY78Vr6xtiMQ/qwXilG5R3nQYF9xBubZb9m5Qf
sSiL5a5a/aQRJ6aHWTrJEvpCCSQVBRIUyMTC6nRXDx+Hf7XNt+rrnY0XdFju
X0vi0dLL6MIiFt7z/ZlkDJRDzrTcTmSREq4seVuFmaV5ic3P08Xk9tMlsA7p
6jzRiV/lU+7GbQXA9KXyUN5c8mO2b5QxBqlh9d4NPRBVyggH+q8ofN6X2D/K
3/p1++O2YJEr8aeKtTzR/mUzRfLncQiNTNUhaQ8/55tKkTKOheIpPeGUg0pr
4hYdxLXvwm1sDD+L5FPkwmda7+8zOTGYaHeobCufRISV6PGeKSus4WItZfy1
tZgrBCn12ygv2stoUArWBww9zTl5h+Z9iilB7ez6UYYYznqWGhSIivL4xMD/
RysYIDTXyK/dxh3qxoUAb/7uhQGCH+v6BgTQljtFSVYlutGY6oAl7uxuT5D2
e7o00U2R0HYWkxGWe9dAeLhHpPkT5q/c1rEp/Wm5Rx5oiku9EPda5YOA+Rx7
qRtFF5JAjdztG88AvGvDxM+yujhLnUkxL1cl2o/qD3TLo5IUO5tyntkW8fpJ
VZYeZxO7cb5Bs2aeGAWwq2NVNHM/0ZV6knkAoWxYFlVkkYVd89YdIXoU0JYN
NVf3aZyFTMpcxKq0k4kQrDBxdoI/OojHrJ4Z3BQZXsXbw+3dIHDMYFDVxilD
Mp5nnH7SSp9pem/1/RRv48ipNUtI+y+y01Scmsr9v2a0bVgBCKFQzq2vQIhP
f3pbuc5BAUGKhL0qZB/Q14ANGcNNKnceSf5bC/DstXBNbYBQ98XXNKUNqp7V
lmP3ggIOjFiTsXQB0e0Ztcs7yq83IJXATWtHQqfyYI/5GZI/FWIkjtF8L1v7
q+U22lSlSE7Qz/dTXINeatHA+v4vGlJgJoEOJGL6g2BW2gBwOVbd6daQ9Npz
2hjqvFgXsdXokYIo6oGhMIns3+KbLczvNZz3d8mIPsk6JZRw/Lp/3UUyD/xC
z8LQC0rHpmW2XFkPI2uGoI3AubVraisV9StM6/x8hd8ymk4W6tmoib2vRKB3
X2+BhoPf1BdtLPBanuHWqQ6wZlEf0Cj2iWsx7EUDhhr5wW2+Wi7YeJ1V3E0R
Y1Od9OvThN+E4iiYapKeSBQvuJa7BzSaoPqry58bXWRGjKcEiT1zraqaVdWp
3fQ1iwcvBlo+505KhFs4Mevjwy2DY41ismsRWmZP50Gl4j305gJtKYkTv53r
Qqpz1UKkxOc4SIH/68Cmjwy3nD6o0qt/f+eXtD1JOs65/wEGl3M8dKWdDFQr
ZJEQeKayz2RmNCA2ec88t8pRFKAfWa70JEF+qRUn6EOgOK92AlDlbDyccnNj
//EkCJtkX1SphyjVEJNC9tGZO3XQqQc11HDGRTe/UJkTDTpJmXYrnkHiNoZu
kGr9K5GUs1pvZ5IkSQDX4nINOLqm0F9EhL5OfXRIUEQyRw/s66JgJ2xMZTmJ
gKxlbZluOdDulBlolR5M5hUPZKowbsusU46bBJVLb7Xzy79lHve7wL3iIsPq
a4BztXTTZh1Izpvz0cpd8xPU6cMh+AVN1l2uU4pni0/0osG7E3592J27Qvxl
KLdxeErk/rezcxfZ+Fp+SnPj7KsPB+yGMWU7LPiRXOWpR4t+5X1cgZligjVF
7b72KmY5+7CBWBuH3qcNWhg/XeIULVjUkPLW6Tfqdk/Hoqgk50EoAIZDuH+w
b+zAv3+GByWl3pXIoJlcqek2G6z0f3yKym3Gr0QZJ/AqrCkY8Ybn9wwZMzJ2
3b4yWNywSsBzWaLRK1ItXmnUjIsK4e+kFSr5EZpx/g/1eEMKy9VnzlnabVom
5mLgraVuvI1DrFLRWAOHMbJ4GUvalnWbSosodgU9HFNnqcqoGvSugvyUNS3h
DdP3+1oTDGtfWb1vSk3ExshZUkZMZFSvEb/QGX8D2WwuImAzf81IzxN41pXt
dE+geUBjOAGIsQEo9ZZc9E3dx0RKs/vimN/REUFRUN7c2SF8Z+Y+IJhElhTc
96jgb4VJfrHRfHHYSN3bxny0K8j4RC3F4NNIQzlE4fSd3OtPnDmvIP058s/i
scCuR5rev6CahhPC4Fv9vjthh0UDY9HzYtSFeo0vNircw8zruCiPwtQAoD8z
hFgsxV8rVZ5HIeIQG5ZsQq+7ZeaA8alkKPRfKa17dxxqM7GmQFZ3qRt/y8gQ
bptjMalq2sXczMvXKjgot352sxcPY8vGQXBLrUnkhYqRRpIrdXfs6YixtmIE
q6VDFexbsJWp/nXcCRSdY3o8VLNPEtHkr0AZ6Ttv1v7ICU9Mu2y5o4HDFNuX
YG8zANMd//qVz1D2snin3D4U9epc1Ib1VL+GSeuGC1Fp7X8eWTXsOpTER1B3
mjsRohRqbleaSIZn/I+4xIUMLHIJdB+YADRusOkIsWtI5Rgf/z3SWvO8gjfZ
xMF/pIs9R+rgM0QUxY9tFUZruVbjZouCyg0SFMUwK7sixZBOzeYmro7T7vNe
GKt2Q1g2Eug2rwSzytB3PUA1zGZNIX7ozczBKk+idprEbOTIs2rW87UbwJ5n
afGldpwPm/IjXcd/26EqxT8g8bAVYpgyxkPhfOB8smQbaRZDnkSY2JR1XwCz
z52mOE8+PCuL/HDQDRwoTQNmBrJ+WxENPsJQ8CrGMuobW2LF/7NvzlzDOb+o
4QK6XziW5pYHF953LzcV0FCcI60v1LNJ71wxFf7O3aUKtvp3wix2doPftYfs
nlHrWfjvEHFRjJLo9IjiEIGTs0tjw8K2lOWZcOpzxr8zhYKTdcPUZQP96x+k
hI+RBqxm7V0/KPb59lWmJ7DveO+zlR5egbW01i/y2QIt6HLSGcY468PlH94Z
ESnmakj8Kqc+SrtHpAShnCCtkwAAg4vOzxmLlvQsCBb5Dxov8dRUJ7a3fmi/
3JJleeEJEelzVE36KKllZQIqBkuFQJq0sPriC6kDF8EC2fsbEzwfI9zmY1VY
enqcmkzVFiY5Wrd2LfB9KfSSyHXC+Ym3X9NcIo7ngM80uB88vpkyfn6irQRG
hMJ7O1XwFUYESxdapZmex+FXbjbccyrleswae+PHm1HowZbwPM03ynj1hZgq
vQgV/Ec4kztKp8ohZOeoHooMehjx4BFBb+iYV8NnMHc7B0QyAOD0dKoH+AbO
T/rsJYr3S/rSYPDkC3gdFW0/j0U7DWrYdA3oQiQ50FdYfWvoWIshFqZm8Yzq
t1tOnq2HDOa/Xgv914PcYjQoZAV+TGOkqIIqWWw0JUOcycUlw284PeX8bilp
kJqK8+hIQlB0igcp9pWfXeVcmh/Sx3UD8vqXkCqPeHFCwZQXiPC7mmssslmX
owPEvAfpr5VGT/wO/E0dwEaVJ0obHe5cL0BYH5rZRWkCysU6PtLhQfhT79vl
E41HcV6vZF7zwVOiAfiuCW7iNfWKPXJyVJfhMM0DwS/E+f06bYiPcjPMOCwy
j47/aAGXukcWkS5rte0Sf68gVm1mGTzexJVUhT3HSDZza5h+a9j5p6uc0b0W
VxPCke/FdS+SQPon+C8MvTAJ2ws+p0JOze5lK1PqY1lzt6xGU6VsqbiQ7iYQ
JObtRoDqlR7eDZ200xWQFvbsNctV2/EWy8nQ9nD31ZC55EWA94oiF1pLeNLv
YXXIWvuDR+VlvIQZj6x5IpjgCCRsC6fu4s8tMnMqc9fVz+RKss9LKz76K2Py
NKlMXkNxcOulIOqyKCo9AEo+6t/REKkxmWRuy3DELxdPUPaZAthYXNaHAykE
bfbPUrNNVR73MTl5oKjum+QQ1q6py3d26NUVqiE6OeoMPEhP7g/uccNQXN2v
speeb5dCDOleBQIukgD7X5g3RszaAJKpiNSTEvN8jY7CC64QBch5eyvhbiz4
8zI58IbgeXduBs4TSR9gSO7KuFOdyMnxrkFN4jgfvoin+zVgYIuiWUwaUnR9
wHywzGp+b2QDwLa4yZbCwcd+xV/Wz2zlIptqicy1jXwVSZYLTfKFgMYnXNxn
ojCT4XEA7/TIWG6HR7j4wKE3eKdB0JmrE6om0LX0mSilkzN/4DzJC6+KbAlf
czjSJydBviOXz5aWKn34zyHU5BBzGeQML+uI3z1zz6Nj+RO7h1mpv2v7tXZ5
5ynmHK2cQ4qYBGO/3VSXCmWRsneR7lwitu77a9/tHDWTKjIhsoaDkOhap4jR
7EpLWww9yvT6HcRPO5WwExHg6bZdFGqABEDZz86BUwK29yEQCPW405Q+vys7
BIWJG946COQnpLun+8Nn999TPvr/1HVp5G5xFDNVclON/DHWWN3u7324qa2s
TnRKLA9LrHQyh2iYGWE839deviyuGfRJQrtvGdq3CUYsKOC/3tVfKbHW6ovj
3yP542ZgLBkU2EcLnVDz08Opw/WQBP/W8zxmwxgKyUlZ+k+oZKTMB8k48HLt
bGwRN/CwmABcOpWBAUPoGYMlZkK7tBAW8hL/knC5/kek2RzyddObA1cJaY/A
5rzojwHAku/qs8Z0/5ETdUW71ElykLoNfwELGwAbYz5QfHmDzji3L+BzqhR6
TAuwe3ixatatBpYleg+JOVYBXjOCHZo7BW15Ru5PkvtSmD7sAPS7KExrTkQi
yyRHhsVDwGomUo0bk+wAw14lBewjxDyVHfGzKJ16WGj4nlu4RWIhXZZ98hRI
uoVIJTA8t6V5QTZFkJTqxwzfjSiR6S/Vg6co0M1SJ175O6q1XnuHvXaYA1eM
4ZQ/U2GgHLoqJs4Woc+Hg5758gcHJK9mmv+pOaPzYR+XR65ZwyaZcaKeO99N
DL/YF0aMxzYTexnyD2OZeUo+Y3pgrODL519CeJ0DJoXcxhxmhbcq8sMY1J21
RKVWzi2mSCFefzlq4F7ZTI7obMFyH+qi53zgQaH0nMPvDdhRqu+ka8z1HPIV
OH62mhFc86q2kQr6w6qfFVoSHQjUbehoW8tKvJ8yRRxYxCCA+EEjra3fTYkk
ItJnNQbwBOY7Z+TQrDeVnClRbRGbjd7cg4rEKASeb61Oqck/Xpsw1koiQacA
pk28dZu0WxP7onx6aMy0NOqUD3w9XdFG172wgxpZVNtfQd74Nr3aWqwPghLB
xTQZAw1dFhVpHOKC8PlTQks0f74nRlM+Y4oWjzr9C/Nsmgxz7PbkvZ8LNh5O
GTydFF3w4yN233iCO5IbCYL57UumUOjuB6+H5zQ6XJi9cDI2Hm2n99/WT1QT
1bDj8ZkrBJ3y94xIPHL5ZyGTvQCTurLIN//yngGlo3KsT9mildNR6Nmo2ALW
12dZm3XqmBnYP9l9/tIZL2BW3dp9qh5M785iHJIBo4UC59WcnCplnLoLa12U
7PVUdB/ydUe/uvCZqnqtnO8pMZgepsJovcaF1OBjTwTJJKDuYmmb+7KXFfko
F5mvEOfgj4uX4Pwx+h72KnfrD+cSaJ8wiBfMIV3Wx6dBOsgoUXzYwKX6pzRH
8tw9kcisa+z+Siy5RJeOpGkzNOsckoE5soGevWC8lLotD51OwxICLRhN41re
syf/yvHZhjA/smt7ZaZ91oivAjIpFT3jr0eNwmzVJRr7pCu+9sELZH15vxCX
EE3IbtDTUc7J8kGIxQvGkI1OPos2wg39sbC7PGIXLMiQJdcu994RdHTN2jh3
8xLHrHoWsesQfa/rtfb1Yq2aaSJlc7vT4+53TSLDYwgfL/qhtQ9y7Qb/Q3XL
8LSy8FqX1JiIBlL9UtXkmcGBTXfzWW9/y8/7uhONbNjVk3u/fMnSvVtL55k4
BYMJbsh+R52z7d9/iZujotr1CME7LsfjZEylTP9gyMVENKKqyMT6zzAfLsEq
WYFVZ+jb4HS1BrPaSxHDI80sL948o7ksCBD1V/+q8PH0Or2+zqhGc/c/DtJx
r4Bp00q2cA1mGIpYWUUJ2xajaEYAHXVDgnDvNiF2AQDEExzUAiayOxlND8Tr
nEh1H/HNEPcakkQkFnWg3ZEB21X5e44OG099T2c4TST7p9TGEFtvqhnby07d
ZMhJYAaS01gGXNgUl3ud6HnjfK7XZ/Pcp/eFn74+y7wLU1BC8pVtltJOjLUI
b5pYPsDeVqVeZyQoaC1X+qsb8Rmbl5c2LuFCBL43ngtYE9d+PxwpNVO5Pv1I
obrpC4im02VijuyCkGWx2k8jwC7mGUIxGx0U63quFOy5TAB01rpZQwSl05Zj
fIMT5B6LsDFUbWGWQNx1KtUVTyf3lCM5t/YMhUlnaEtc5bE07aSne8j8sdcW
9vTob6cfDd8n5OAHuIickOnL2DzhA1CUWOgRhHw+CfVpmJebMTW/peSBSCTK
/PwKPLNb6LPUxUe6zmIP2QotRBFQgk/fwtOPvKsWgU6uKE12pVb+YE/7pDSr
1di+EnRDVa5loQaxx6fAWtoQ7fP95sC3IW38NNI9cahotBynoeNc5u34b79v
4n7T4EPfKNqUnhB9GiiM6+a9lMkW+xky3/XwQiTDT/adfDOmoiM8utyexTJm
S6z0G4G1M4CgR+itPLYbC3ziBYB/yVKwtEqd4AaChnzZ97YVE5DKsQeGMKus
f2/NAatlkNFGbcMw6ljOVT2S9K6q4MmBxFZD0yvJTrLZf8rQtP+N3dfE5zTE
tghMrh5MTxUmL4s9xHEvAQ2+nfjByVKUrwtecpH7Yy0pZaq6et5Y+nJ+rkp4
xaUSXT4tM13YmLXyd3DvOetY3HJgOWPzgqtSYwOyxTB2r4YOR7D5LNuf0n+N
7apaUZZfnDtvYsjAR6qwj7w6foIKc/7VwIMWPtbo+sewwT2/i7FpwkRlTPA9
wYwOPUSXt0pQ5Aifp5lAcFtWtCeTjmtKythm7tfCdD+kKXHQysm/cp3NJWOW
gn4Sh+3KtPGgvGk/WmgiPRMCceMqcF1MZ7gqYHpQMeuRjjVXJPnBQ9jDPyUL
2Bk/Kv9CaYa9X62zCP5IGUC6j2R7unWL9T9jyIxwsdR3UUQ+JvV/sh6pRwFh
ovCi1O+UTyIHpPH6xY1ZAuBXCUIlJhnZ9Bo9vIIQ+8Ii780myMkoTokbjQyx
jxfJCAGiwcz6iMyB0od2l0zavK3aDj+sSyuWO1HG0/t8RekqWBxqjatqxapc
U02tX4EGK8fnJzBRLafkTElF6kXcvn8VOFAy/PygeKhZ+aAqpR2ynZFPMWvy
tloax01yReHebdx45SJlSIy9jm5OHjVAcjSXWaYsoKKAtGcpj1fFXkS6IOWd
lL2twlw45OHD5nHZSciOP/R2rn2yLid7rwoViF3SjMZhySJcXHSRijkxqGLr
hVgaXEcuvEABxyQBjZZxnOnlkxzc0UPEJ8EpLENdMEzc47kEvlgHsO9Xc5yZ
q/fTV0SpJGlRZGRJR58QkBhFGA/qSDjprL6wkIL/cfcdtAT7rO7ViAC7RWp9
KH0SBuoDe43GPvk9cdjivr1U5S4c4/O0AJEJjKeWFXUKooVdFfF0U7M/x5Pu
6LW6WvKlncbQcmFhiZXWM35nZGsg1smw+QomNtvSxlH6Br/nKzsAenrcL9DF
kiG953K7XxjjWHcV9x/vh1Lq3cvQ383qAxpgnhtUC+0Eb+6UGBzvCPDKZMGN
rWIA5wrHhyyMpDE+kOOd5P7hqNWm21BkdSUbNAq9u8ycrfzyGgX89eyXQldg
BzEwO2r3oC9wrMaYw44cKKkyBIaLipFRyQhAw89UbLtSubYbNWL/WBvXEw+r
kDHFK4fASPrSWcq259+g9LV/1gXgSF0psVS1wQvqLEbWdwHz1zBhC8NYaxdx
7yHKFWWf6rJgNoIGfnIM7ehgfeBWnmnJH/ix5L7aaUnVPiCVcLGrCEhGLmXg
OtJqRuG333Y7JQ0IciI6jfYvVEI3oOEKo9C7iVcObquW+59N6foBVQxX7vPq
FoVG1VpmF972r+N2D+J0P/l4JJVl+oADrgcHN3AaPEk2WwU/5+d7na+AaD08
L8d/Tk99EJ6zEvUtQBgg+Ao1yVjsVnrtgKrKZO+3gk2QO1BeZat1mA686qgm
6+egyXbVvzFCoKFqV5h8B9ts1YqsE3cVDltmuTm2s13IdUWsSTIUh1e9yCdZ
8Ukkj4oJdFuVofmJNpm6thxZfITkKN5bK6mbZkxnJx5wdsJznRd9NZHede9f
ipdJd7VkwO5++DhTseG/mok3QA0VzCToMdfwcyIDkwB1rZaqK/bwnhQ+rrui
XH8diGFY8L3MP3LiSODd6pL9w+9IWTRtgrNL0SLvUlkC3eKXdcQHPsCNDZt+
tmqoc71wxHlY7EYdODaeObb2UT2i9NfCjz753mbzpb78k1TajyVRNjasXaQ6
dBt6740bf1qf+Cloue8IlF6geLiuITM6siHzMwpCw8sDYVsQLahIaSjtApzq
CXXEzRQxlVTWO57rpar2CuWBIH8psoB0mGXcmNv1KT8ChXaUQvWuZfjZGq02
WHqjC72s5XnzkPpK6RLMxR3vQapo4e4GEWwRdcdGUWlxJASPd6TpqJPQnGoK
3P9D+9lILzza63I9xz1/LmurBotxZmuRjCmC7Gmf40qk9mrEA4neyKn4cj+Z
i0Q3oiY4N5aCqFX+4ZbAJ77x4nD5dhPtgy/lU7NMLP0bXmtsDzVBhBR8CI9x
HG4xhIF5buSZNrwbSudgozbdj7OYBDC+6HBdzpthWukaM3s8Zp3D1/2KJHCl
MWuBajFRBAryibHi2McP8Xy6tbxhmgEsTzNHJfEwGm9/qpwkId2M5TKGPhlF
XKUJNvpCzxFl4EzyzCEisy5ABT2rAz6LPu2L1XzqBTars2FQfIBRbkA5YTp4
HqdIn9yjynZTSmhkB8MepAtxmtg9hJJCU9A4LXotu16RkpuxJSYc/qw2QBgS
GcmGG10xbGjH670DtiZM3yLaEZku8kMzeBcZ8ijnq6X+cMESTiRlsNRXKVas
07EjA4i2KyxNZUVroPhjWUlEaWK1KrK6w3PkFu8Uexbgqu9+1TJ4brJhpBF7
zCkNGyYGRBg93WQEea8//Yy6amnT//jA4jjWApi3dqlfwvH2uwPRVPMPL6kl
no8njrmNWf431Q/VhIMebMZKvoVFLIYNOZxXG+DbGfpooPtGHgO5hijBvSJO
bntomQ6tsayGdKbUoOPOQqNc8A9asnmgCb8vp2ZQKs+OX68B+S1nRaZRkdMT
CR1AcbpAbGhg/DwTKHdG2rewvHbpVfRVT8ucLD4JM0ZuEc7K1bgGLWII0sYY
1b5MrFeBrvca9I10p97heZQzRbRCKO6GNmkyIcoCHjaryJT5aT/xRa6RtxQ6
EwvvGvayKf2j6RTzoFnq3W6ecDp/3DviSXlmfragfsB12nb1FvF9nFXqQcOc
V7INE8mlASInpdWpCZR2RT9WnpwbM+gwckxwdYAPX2xUhDzWPguM63V4bWEr
wDnmtMLmCcl6fk6JFIXXpCcekfOklqRsCWVjRWHWq4S6/ervgEYaq7iPpYkD
K1TM2KcdAmVEWCV7GNxHrPd5r32UybXv9OjKBoCj2mFxA8YpI6/0Cr+QEvcI
kQMStYvgJpF9fGcYhUqqiS0F2s+ish6RIrKesOIN9ZFMLZOTzmxz5Q4jeCom
NivkE6ruRe+2N6j3FXY/JZUJNfMiXJSejmFFgPfVtO4iSwb4WwiKZe+o5t3v
a/dIlUhAXObhyDTkHKxHdDmbzEQIX00E3ypkplbPwU3PVg1U7yF1fk/Wr/tw
4XTLd/9radWf4WXmB1HHv8VvxfQ4DvdKZnV+98sIuOOm3+bPqOTcynLCdQO7
wCZb0zBx5/FT5gXDfvjpPFhrrjh7RrWKD6ox5DFOaMYF+8m0EBDRz1uWivdm
7MPlls9DuBO5f4frEqAlEtabmr9tmB7eeZNidVzIKFRJbKrErx3QvGQNeJQO
n0PcXdp7ZkYqpiiiqVoyzurktA8D0hw+gVh8dqRnUQc+W0EtfjD9ccpg1cna
3B1a0dl/r0CwYME47TCkIvq2pBTtgTWSTkwKCQunn3Z9BXOvunOTXrVYlciQ
L0gQhCovTSE1+VOaKVvuPxF+tjudd/x5s3z+ieOF8nkVUldxQhnJ611OHV74
NytCew1IeEJugB/S7I8cfONSFZ4GhlfBWQ/yehMylZEZWRRWOV+ySHsggeAv
DsnlcmuErJRP1huk20jbNA66Qnpvy3YRwjxibrSdBOAUibd3MjLb/kSL4J9L
owh6cH5q6s6NCnl+ji2aR1rRqQPJKxoXXPLSVf5nvkhaG1mq/yL8fFjNzk6R
0ZlGmuGE5drXANRnqMdkK0iTsQ/Auy5CMS7HLgwUB7aPWZT/rw2ndA7EuV4m
fEVMhsVk9v/qlf4XSTPZW3qI7ocA1aQd84jil0Y7dX+8PMpjOVK7zSUgVwyY
EvWru3L2EL8mucU960T1uVxMM5ozQGOsvfgtEkSwvHPWuq/7oyaqOPQUrxan
qLCw5ZWMFL+E/1CY0mAiXRmFsakCbLtLAaCFFDwhKGKKnKlL0OX8SyjoZ0pr
ESsd+voZ9C6byXaMSxrUYMONMVIqLNQj0J/qHiFLpBAP0zep1s/wDbmF1s6a
X2qGOn0fFa7O+TmRmmu4uQo1b2/69H60fDTuxMWwRKzJQv82Az01kNR5ey8f
TGIoP87W6E7Fjsl8hqsY3TBTLSK1a5QPgKp7bHobBnDxPGe/b9jDEyVBMfxN
VbyARigZBT3Wl0m1skKz4VyL7jWhAMNOcFcnT68JXnKWVPYJr1VYPyaYJtzX
x/6Kt9lbrciPe7sZOdYDUk1AZmE4vxDuEOfliyHN37ogr8AM1Z1/m/cOOjWy
/Zsnoc+hTWuevbosgMh92t6yC7dDl0inJqSwrY2NOGkXaHGe1J9fWtyuWLAc
Y77rzzbDZM66MDmjCVyGHaYRDoXkOebFoj1P7eJ/IjMlPLi/g6dIgvBxjBC5
x6J7Dqqk7F4SpT9OSsnwpGXydeYE1G+4JeybpHYCSVZJPpBSqe4xJj6D59nT
L+fynHZ2Gc5La3LDckk6KGw7pRaYf5ie7cLkrF5HMd/FdFoO8lSHONargw/N
SKTR/tkW07y1A4NGQ+wZxzExG3/BxVrv5RXrAppYBIw8aEZQnn4u2K+jBPI3
jGA5cTXlfscTrA5QZsFMsyTP4xanlN0WXMrSlb552LT5Dzwq+x4FT50kIilu
uzD96WW9KYG8hrqse4Br4sASd5sgMg96FWqPvWN8gYGELbjj7KdOg5cbAWnd
4fNN35W3a1AHP7bEedDmhU7n00HCHkoJrpRnrx6bHLNGkDhtgiYQfkk9BlLG
sJIycZqwVkVWUg1jWY0n4kgt1+u9sqqq2mW7pasoBXTgEzu5PnigXKk8w16m
bj/jeQLOqDpjRk3MEKHAGSDWbtvnaTUC4eraIGLUYrS2uskWJ9vKOKK7VsU+
btJh/MaFQFd/HobfGGuRL06cKxeIOvsqTKNwml+99BAH3JTLKUNANRLJtzt1
1AWx3u9Fnjdv7uKtb6c8zE8bLJAhG2G2h7V43/K1Srq2VQKKc3daaxB6ofJa
CgFzAHIpIJjesatflc8svSeDpnyrXl+hRbsX6A3K5+XsgRvEbtnI9ndhWJIG
9bQ3T68XJBIae1lgGFL+AIgOXvwQVjk5Z9374ccrIto7VA631adDrna3TpqW
5uKyqaE20J9fI6XbeEoper5Zjr7RIILPuRl0i3dXfg7cdms8xlbsAlYYMzIH
jrXgSS6Iw5e4AbRdi6RYqIMyzK365QSqQCopzKFNRFM2FFm8d7VB8039JT8t
cNp84sJwL28/HDgfNBJ8bN296OPR79By+gLssnB1yko+9GTzh4k7xIHQciIK
A73TpcyXppk03Fk7UuA8+cFXXkuU6Q9knRwpTVB7vs0UEPv30aiw7LeamgEV
/s5IVYFsb7W6/X+51pgtCCBRUbEiBYyFtG7eQslqBdvWZ0K7oAAMvCF2p/RL
E69sIGraAUS2bqbsEY+fzQEyg39u8x7wPbencmjOIajDWDhOda8XuJhFubaG
WmMeQPLwt9U30U9zmtMBEoowhEcffbA/kOoxEDeRBATFqEt1i7VPBRSYdREk
dfKpdO5NamWnqFfwG7Gv9G4zBWTP7FPnOnqixflovKmvgiENQeSmhA2YeBKC
b/Lf1F5mvGt8h6bjbb0zG3heLqUv8o/1SDPk0sV/5/XJQmabPM++f2bvVLPd
FRCvqdNKXfH5K9T/6A3sIDAHLh7kVF/SEpGbcLaMy/zbfCrPXy6U8iTe3248
M/JyMYtqJygwCdQsM1QNdHGelWVKVGAYY8cXwoI+T6JgrPeut7s/e4grYCeE
jw9G5JpmExXH2w5qlJFwiF04/aadQywD1sFVuxr+MAZIM/wbXrumlF12SL0h
KxqMaKi8SxZYgzByHK75NLnzzASMVZ3rpgXbygBYZAg4RdTLNu7cXCZABQmo
c8oNvgh+97QbSES57JlNq6KwtYCvBU7L0qN50dC6mVcCFXtbCJeBHJxe6/hI
NVISb+ZyiFiqnFGiR0pTgVyjnOTiWTyK1BSTm2xUXUAluRzQ5/Oz+YYPxCbe
TIzyUb7DEHiTtVNdSiK2W1ur3ZN4K4OJyqtd0jbbBzLvqe3Gpn5tTTq5MlCO
KwE0uKS1kE7X92tb/qu5zJ4SJtAQ78WoHjVTLUfEw+Oa4q7Sv9/x+iJB31NC
EbDXaBN1tivVKpHW00TtXX1S6xo5JZ9VC1vydvS95KcgO7/V3hM5kdkCMdvB
oriDYC8VDkJTS4XPZJkTrNTaUf9zMCXStzAJJm8WOTqM8z0WdspnV9XWyoLZ
sb7lLgbEnMvN/D8Rgp9SHoNAUli4NzeGy3ngv69r3MU9ZLi800jD7jgbsD+M
ZSsew7yRm/vGixXDaVcWxzz+0tmBgitPDut5kQ3MaRwcxyGj/iIh9c0vYXY1
7GIzVknKZz0MpdNpL3wio0/X8hgkkegbCOMEx/I4+MfJtOmkvYKu9+N9x4MM
Q5p2mh2gIDj1qTfj68/6SZh4tBvynUfffXa93jnWSUse1q/rsgoUapN0HDfG
9gKHEHuZ0ULuPDCUWq+kPeqpCUY+n8gP+dO0YnLRSth0/K2EkLXBUr45X7AR
eupG2IT1lj8cPJtR43uHlzccDwRP5yhIVKbK1fIdCa7ocgRRLvFwmZRcz3+l
cN6WvmiNdDov6ETTvAnYKkk5eRlokyTZcQcMP1m29g4e/2Z8X0U1DWwF4RlP
eCVMJxhQkz5yL4pqS0AzvjfV6zMAiI+W9HlpGlHR2TfYNNICAANWoPj9b/Ur
Yw1D1iNTOm4ICXx1+X418UAM3zDlz9/e82EjIX+AJvYmgyVjPDrnATkr0FAB
VsWifxUULUgOavv7XzK9uczp4WQ3U2JZm5EaEGjzgH4wYu1+Y1Q2rVwsy3z6
gu9cqdMFqggdfs5VOG14Jyey9JC3bG9LxU2/Dpnnkg9seB6x4bjGzPKMflzG
DilIJgAIM8JRFjXipL8eD/L+9HQC0POSEhuTBTlw4F/NCgcVBqWZiQJqYKIF
dMycegSANS5CfCYU7ZscP8A6hOIFXFhJHowbSfJJcwBufzdz5FvGr8iOhwWn
gIrJ99vXIMFB4zP5XxH7po2nF4KFyx2uBLzVnEylgyXyPXseyYnJaVgqhdRu
W9g1lHq2xRBLvNMozfMngcfLoIZXItsKJfgk1y4Mc2TKwgThKT9xxTE18tdI
5aiNPjKg5tu3ZaEtyv+RNO/qLTwBv3lnTtgV9R/RkTvkWJg737HYDLjvEQOo
ocvZo56iDmSgxRHKzxjKUJozckjgvnZ39j4x5eyte1SB+0i1K5p4nL9eRudx
/cjHonvQkcgqgUGdyCdod/OM5NETLQPQZPLEp/5MEZAfnL0vFszlU7cbZhV1
uQodQKunnu+xLrVZxRBMjvWWBfT9nawNeb9O2UZjSTsk88uhQ7oZBlLNZKL4
3tmVV3N6Ez2mUyEkYcl/jZXr5MPerZFwo3t9uPkbH6kT/VHjOFXhzBHP6XUt
+bsVxGCIJzQlu0MBUUFwuxD3vA5RuWLo6UdrOdWyeeEUqJYKpd/j6b53NLEB
1/UwhjTEIFHtMu9GLlmUASc0lhySpDjLfz42ViPk+jBvfBDjsfKVNyA8Fk7q
LBngNWP2AmmjMxtWpkzMvFwuGRmdQa9bddc0s2E8SIwGBPGt7aQlmEMSLtk8
+wuKYjdeZhJ6EZZhdltZB0yfFPuh74w7k83/wDOEbLLg1DwAckwtev8fOGXs
RnMr34YjQRsHJAltg88t1c7kzr5zvsGOnQ4T8hEbbEY4a6FgTRrjAP/uxoeY
aBZsOlG7jiz9/CZuElvHX4n6xIhDnTnUZClg4H2tkJU1YgMaBc8azAUykUvB
WE6QxJhKwMzejGGbanjWTW49ZfSB37Z1fIQYCXVf3i1hj8EanrC9yAYAh/tL
1e2Dwr2PXa2xdrcYoWI8GweeWYtJBbGSDtbsIhw/iCAANOf3TiyZ8t4mxRM0
SmlEEq37Drq+bji1qAnzAHTBmjT/AhrtTgzdZ79CtlFIwzIweCEXGZtBcQ9t
1GMl2+PY0lu/hEZ17IRb0AGJMmnvFu3yk8T1mUaZh2axMguX2uVlZk8hI9vX
zZhyKmc+qx5oE1U1GRANt0j/xKJgsC7+I3FRFzsJwAcb+xEJH9uuqUcDdtDv
7qTen1oold3R3cClnYWv/5GNElN1NYwurtsHlXmAXBlJyBx8iPUSiJXETkGx
f4DyCzxe+oNKKqUyOqZAnnYI80/fAslR0b5rnCUcR2Fo/BPkQWTPrKVYmLIi
YcsEyAZPsO8siyK4AnVYRIYFge+qeryj/d9zfLFoLDIXFLXzpQR98fOZuIAO
vfD/EHqJ8TLwAfPONUB9+b0DoD6IPISGY/IBu8Cuh8QyRxpoWa9ILUgXFyAv
HYgDLRRicGiQb/ZmgfGcS5Q40OEzEA5RTuavF5KwXcBAcHPJDmzQU5HLHJi5
Gc5Y2FFFnJoIG4IFx46Igx+2SYJnewKZBZ3qnM3DDe4mDPvw5Ozz9Ue4q6fE
7CgEvDNNtmInvOLlyG3h6HeF+aWyrWdKsUzaBuapGYnmWZ0IsYtVKpxq88Wg
Alt1pIquPrtjRQ/cfipfa9Jy+XLyBuADIdxChYTmks1+t/u6e75NL4PiLGaG
8M8B3WbAZxobw6btgCfsXZPz70URrnHSt6kCo3YGGVIPYLzLcoGw/uJHqGSt
3n9bBEC3GxG8KyDdBc/rsDPJP30cFVhlxWmGGX0xTLIsdkgBpTMNCnxsfjnS
YiW5R2DMtI/zGCS7MqIWhImS/R8fTb0wysYZVK/ldywmnbiCxKZG02HtFivN
E/NtswW5vv49Td6WdiGmmXcZg3zoCX1cug4hxBAPydlfdJsr120tezZnSApE
V6cSccm8qh+ItFgxl0x60X+ineJeBMa7w67WdWVPFzqdqrhApRKA06S71p4C
dg2SEikeQfNXP3wAwqtcpewNBzjyZ0D2uLssAm5sYkvafoKPb8N3PeX1q0nV
htHCrVwotVhSP54Y7dxU/LC4L4z3pOkHcZ1fQK0PfLxnQ9M0oRXVXsYZyuNo
9/zpKzKBM/SD2PHuJb4YBs1dxeNW4AuOU4eJFkbF8v0i8rToApkJupXEXu/Z
EGW2/b9SfausYDHD9mv/9udsw3hLW+OIjC+zKTpSL1MnXOqfYDGMSNAHFROn
jn8GT/F/pqYI2GIKfpzc2WnChwiO8U/wEip0T2jtv1T+0UsdWJvlJUFIhDzy
jUe16csAZRm/AjiF4ozDoYLvawsBsGFD3QWUPtl/HHOcTXIUBu88J3kVGtqR
1onAJqAzcywtxGQSK1JkPF5pGOcPvKK4+C9wsNgdbsmrwEjnDRH+0SST9hkV
RocHMou30JJ2HHvUSVv4sEBtVDERDWZoFIKvhYYNewMuyZ2I7d1+9pBIv1qT
nv2551i6xHKilpjidnBT4ur3KMCLoDKY9nzXYOD+t0j5RboZNqjhBWf9HHEd
Ec7OymbqF8EI8oHh7oqhVG/fQlr+9pac4UOXlCC95R4bGc5yNjT9aFixC7jl
Bk0RVK04mnn6fPRsiHSatNrYaqhCergqBp+CKnUpel/T7zzNeucfeAfvvGyi
6y0P4emKMDP1GuGoP+3jzQ4LB5j1UfOd64JbH9eKVIfCwDXSaRdnZRjcdkZq
+ceDHYY4W5MoYrITH1qaqB579OOCuebHPPqhdjkJQJ3zmVcUeoyTKP894cLM
7hA2415iHGcFtS8axa6LXEYz8PHQCOS7iqZPooZGrJVLuEFSUkWjsogyRJ2K
W/InhfbmrhxNXzikY4Fxm2d7n7zqNGqcgaUloHobG9MHRZU7TlZCJCXXIG12
qkUsIlf24obistyGtccMbWgpqS/eln1pLFzUoQgbIjMKB73kqoSzYUrDYcfU
oZmIsGQvKDEKYZRhKDS+UZb+Kw0QOZFVjUT+b6muM6r0rdfq4/wEkoUnBmfd
haeeRQ4MPa0QtnXjoCjI/dB8VRnoOGlIBLhUZZ50m4Mh4hVf4JqSfE6MogO8
lz39tzk3frPGeOBt+AYbCbBL7cL1VveooGD1gn+fp0Wh6x3ZjoFpAQ+qT3pK
Oc+eLGauYvTsgUYNNZPzG3f3UXl25mQE5TpRleVFt+lrNJ6TawJCeXQkXmEN
pBpxYTXIipG5chnQ5mf17Gjp6pok4WyYkEL2LNPQ4mB5FxPgzO3Y3dXkm60m
/obELW/IZmHBcsnScmUm+ac3RBf4mNB/dttbacuBzDIqrPMlIPkDyrMihxds
s/xo6niv+pERjTZUTSaYJMVsl4bo9ZwsP1uZCxGHRGaGBPjV9gb7hSnejXZU
vA6GldBVfwpQ+bB7ozHg6//Y1jK2dis8LoUVyKgaRK4kyEgKULu+oITfyUA+
BT83zd5uRdGbDzOr6vclNSZGMwv2KuaK9v4h42liMqct4JLaTflfg4ho5mkF
WiiHbp0Kg+GjnOXkF6FQzK8QdXsZf4DwR3pA1ybbaVhjvZefIz10lwqxndRg
C0q2kiFwWNkO/lFmxVEhJpNfLu5nLM0XqOhBBGkCt4n3MpxWUJmhzVq3ttGP
nteFTvgbzln9jB5VM/cyQjUzjIaNMJs/lmcLX1ZsbQ7zMY9Q92Oj9DjzbZhW
aq2ViPGrvGg/f809qLDWP91Q+4c1YW1OZIDNHPosizmuLKCTGm8lh8u/32ir
SBY2Ltq8DAZDEvvFrEBSBQdcrBWSDdEbUyNdIKaaNJdW2i2+kjboQT+yMjeg
t3pTskr3edYpi4/KpAnmWGx8WrZ5qgw14Qzy4INKDkMSVMzlZvhiZ4CAY0d7
DJm1HLPFgW0SpQoWEMOOPxCD3MhGAk4L9nCnbOhQouU9+/FADldGgs9oVHz4
Wwh1CuNxwKfBIScrU6FPgQ+gcd/jJbJsmlLBB5lLYHtcmplI6Rp3HcZOjX+P
+6eDcsrY1uHM9kyScv2lYCARjYlJSLfFfC4a+M12c+g6J5DOUakHX1v2Suqt
uHpHrZFejA/5IUaVRVFn17idU9RmoJ/9KpcGOWuVi8+CHpBcIrDRBNQXA9cJ
9nmZcwTXuVqCpKgPCpmdzW8rXrcg2s+FJ21z7laC4DLf2PKq9kGLnIHRPdJi
6vX1R9BMkjs0GL08cltPw5NFzLhS7qmRESMWJjrmsAErRoBLtH9+7VlfU1mq
naYOLONtWNlcMCbxTRSSd1UqHmgr6lIXXsal/NLW6+8OFambS+2EsJ30vesG
NTEf6FXmVVuPDZhXwsIU6a6HuYfZcDJHnH5vJxfxxSQPylePme/T/GmChQ1+
BCHYnR3xV6rU9mjKOKd/4bXW2fmjpJjE8rFUCJ49i4B6BGeYiyG25av3WC0C
hjvFUKYQLnWMNI2Ja0c/pfNDv6c4lAOkhnYEd5XvPcOEIbPbS5EmyMfg6fjj
Z/LGWsvqMbdXCdXpLQ+ctMrj9hZFNNBswVTA8vbTc5Ox6i5jE4u/o7wWRAR9
A9rwGZlq4AHCo1+tkLxLBQy6hgoFNxClFejrHHXVdfHkHXQErUuYOcoHSU8U
WCXDp6xtmVCNbTjxZbU8yr0RvnE0flDiddnFhl2EsZC9vZqhrXXosSjsok8A
JNDSKW4dQHs1cIvMLAWACsV2G/AhqLBnpz71DKpQXAAAhHeTBOrR52JAwwLM
gp9iOMdTkZcZ+HSDUsxiFIznwqsqpZcpX/SB88wpfWM3Rn9NBfgDr28+vRTZ
tqf7i/mTHY04swBASapSVngsuBll0/iTh5F2w4db4EnmFoV5pbtqUO3cCSi6
Zsgn9A2zC8B0LSNqshnlvKVHRF901etT2Xfx732pr08Qt5c1MY27T2MYw9jr
cmcabOju5SG2LqrrScSHsEfZUhEG7ntfdAmb7VFKPi8Lb5/6ubR+hGkc2Y5A
SvrZDCzOxwy5rk9vRDCOlLq321GBogzTTVKlk/1EH+foveb4r7Ss/cjv4WzT
vq5aia7E0o6hHk83O3D53t8QJ5ddOW/TO4vxxA78ohc9nmvH6/WxZJ/5lSwb
5qku70hUNkYS26lCPTIYQV5VBIneLrrQ23x1U9LoDBhEy3yYu9U9pH15NZcF
wtLsXe1gUamK7mA9t7gEaEkFRmP0nJDIT53uY5mMzkjJcWNiLQ2CQE0ebqW9
TfmRYK83ys3EhDEJPLkjvo/9XWR1ttZskL2uwQifKyOwovIzIEwCp2r1hJ6Y
whTYgpepE03NxgOyhSrJX5pypffQu6cuirQYzM+N/3/8jlRZ//BKPq9yvUEH
ya91QcnjI2sSgtjg099ny0y98awCs91VpfJ9b5WZoF7sUel/HL5MzWg87KTu
otqAQAuN5GxyVQBrFcYol9XsJH0EcZJ67ixyALAl0cw+/FbwNwpUwIH5K36F
y0jWDfNHxQwZ8Xke1eZqKI3BtkJum9/W+sAb51o82iziXTN68sjtUh4a5Aox
0sjhrR0L+GPxS7lk8w0nuH68Za1fLqbcNPUq6w5h1A+0iT37Tkv564OuIMcl
qGiGZGeaOGHbx2GXwEKLEQGdUjiNLrz/untngU6JxwPgV6huUsveNurKbrFa
drmYSdul8CFZpkVkKB2b/i60jNbqvE2v2owzHtkuxwDVYe3Db681RGmxP/0P
4u7nN28XI6oVCrElrzaWW3oHMVdfI+7UPJgHqrLqgI/zX3h/Kd3Xm8VZ0Obr
9ZIjpVBcvbnPfFDy9DW0xoalP2M6b7XIWrJTFuIWoX5TzikfiC0izMWRKMKI
XOGlyTs8dlBLRvb4zt56kRy7WGN8VqsyK8G8YsJwRxlXZfkQtP/hsR5qlVM6
5yy+7YcjtlvWtG+fxC5k2WlHY2Bb9JEiR+FNw1UfR+3KxGVHNd331RGD+B9F
thMZunSNff0y+52aCSWpEvZl/MBSZ/9/lQTerB5HOwvCppPYHb1qjDL5fNoB
9COQAazfZCCcoCHP2rd30T/9bCXmF5SF8zuIJwevQerB3NgF1hYid2LpkcIG
Rn/d85UpLFtN7pTEYZByZWdHM+lBAycHzcIr/6Ixs/bhj7PPuc2qrRnObobD
Z9gbzH1wZEUI/XiPjwZQCC7YsTN4G2X4OWfKSFh94m+r6wA5z6mOrkhKpiyh
Le72ifYyQB0gsgNVxN4wqH/OHOQK7EbX4OOtrjsx4jpULrEDnTUlMqLpfT7n
e4RJBtukKUDuadz8d8Pzb4kvel+hztkwWhjWkN4gl+j2KpPXNqSxMrkmFOip
Yxw5GGseFn6yJEOEOCpvmjQmucdNkHsCGhhhUE9zgdbslYNDi3i14tyKJhex
ONM6G61pVuFvGYoIgvzXKJV/msjpILnr2Z9ASVTwnl0vvH23l/YOt3ASteu0
JEJZD5d89DatupO4oUhUEcCU29bXz/EiyGZDYGCtr//ljoi8mQucKRuXr64v
yo9kQdkxlokt+iciEBzdiYWemcyIc5lx2FLtp1sX3yuS/Ejgn8UbMOmSHdTo
WIVMCq5ed7WoGVtcrXcdUD53SV4ChoZySrGRxE1CrOu9AXoNMKLaaGWRTkMj
RkM5PSQ1BAJIhkO9fBh+uJOnsdl88HpeppmwRfZPsuT1tv0N0hefuNfhJW3v
TlB0a1NXKSjPK/T5uDTWdjA6qJSf/S34NO22aXUIeVZNJOhsMR87hOx35iDp
tTIpS39DX/eBULmdo9Hco0Sahzy9Y6n0gyxk4XxSLOC8KQF/FpYKA3QOILls
UiyC2X8zsKTvScSNPUjV7M2ZHU3JDiz5ZTORsgGAXkjBhdZ17kSUhGPSI6zn
bA3NVtXT0LdxkmPY5Fw2raJL/rMZkvwEGIJ7sqQPBfe9A/r8HxgOIYvKEugi
2ZRYEFVA24IcDuxgzTy7CiRtW1ZEZdjnwCjYk+dxOU713DXUAr1TnO0dRYk3
r3e0FMOLJygHckhxIljr+si2M2hcmHuInCsXHPcQPtsRcnNDheh3tBtNvvFz
IFlElG25StLivH7wcPtqnRVFmXIo5tGV5YqKbmHy+ynU4Cii9+zn6yyrdLRi
W4rU3jwcNQbYUxcrQXmPjuwLM8a46JMDwFCvErXjL418y6Uy4/NPOqYP3+9m
pP6fg+bo55o9TcHWs2edFP/GvMQveNLAIoNMu5VXZT/MVsQIxHuUdookzCmB
R+z/Zg1+XB5Ropi1il5mHSEpv3iV7dKsynA/rM5ugLE9P8d918z1ufjGfk7M
UCKIxsxg4roVFClAx42MNjlZeXQ5G+p4Ugof52opcpEfyLqdnH0wttVII9bO
ITkvxdH0BJW6sHinKUUL7YpRHNyDQTEDcDZGXET2h83tRVd5KRJHVzFQGLFO
SV4nGIguUSWeillwTJHFNIKYHru1CORCEsx8eAVaor5ixnTwcraAOuyP9iX5
uXJyX9q1cx9ERF4YCIWWYpvESFAwUhkoFqV2B3NaGnvq/kiMFHgnA+SC8uLW
Si4aGpo+lafvrHuKoPAmjIL0BBvSk1x45oWhYA0gpakAriIMDVBssrC8H+wY
4uPtj05V2dLRt6Qv58AI1ONawyoNIwOGg0isbo07sndhxoO2HKy/ZZDh27s9
rJFKWCu2pWE+RGIza/1ANgdwDsH6NFXgcIN2VIZn5xXkYtjDneimbzZorD02
b/HgTVn3Br0Zk+yqfeiix6eBTRQj0eUffa4+nfm3m5fUJz+Z5ngBT3k3dc16
/YVcgeIrlRBMbMlVEo4rJmoqRMAKoGUaNXlP1IL333BkdNWvIXtwuTXFKNlU
opCBSmtkkZ9A5gQkQndHLiEjKB1sblUJ88aIgOLZ+nGfb98+nkv1pOBXwRRu
ArZYxeQ/CajKkuGZjBOF4s/THLzJpc5Ulk7eAnUVQ3Af2o62PTAnktvEjmmf
HdlxGL7lAYVuFljp5G29AeExqm1niU7S1seSsuaso06wucOWg2x9Wh/DdlgG
ea59Wi6KvxaI0X56HHiK6NzbTt4D3azIvkyIPBkugr4A0jwu++8jiwbozKl4
07RjJRlRhL6DwLfOXnLCp2o0BySd2Od+8oqOkZ6f2Edx48pQJ1/622v//9vH
GJDZkanYoCEJaecUMYHpNNRrD8S4tHXZFfHC4hc5jLxJFDVyjAhwH1QUrMsP
C83gpP427vFGQLR9tbV9BLafA55qT+Y6fVs/Tv+Vu1PE53YBpIdwCeHBprNs
bM88hTzjnM/hxW40ZgNsq6R2eF5U/iLzbxlYLcRXbgd4P/ggdt4MAvQTKoCm
UU0PjTNstjLnQBSyNCmO9tyxIEVH9sfiPse+L+XbJmbj9Icshg4QxRNYVGSG
9Y8jZ/R0++GVX+YEqVcVqaifgPZnTw8uRgytUvbFPgVCSsRVR71l+rgYXSXG
YvdRtjb2T2D+43xUbKbZ3oxxhxP0MVq1qfd4TgYZiDG7hHI4SSl0j6urM3ho
GeEt8ZdJp0yPbPQGYYf+MWaUf28xJO0JE07peS/wTYfkT516B7qNyceo7aZe
0UmMvxxVD9ThY/g3Phq7pgahTpSpYWMRRUjp+3MVRoJ40jr1+oUJwXvXpd+x
bPds5J4ZSY8vIc23XhopJWF9bDAiK0xIr5l6SfQwG80sIPfIXRJCEZ0ctI6H
hYLZeJ838qOsf3hueyJ2jrdnon8StDcvVD8pwVUFHET1K8oRC3Me9CkPuWSy
utTbbyl5jGVlZ6VH6Q3HvIrRR5U4Cok+c0NulMEgYNgEdWeEzJwXZvKDtZKI
kh5toj7WajNNHM2z3eMVhwudw5hYURkP6ePObcZtUZySQlhrHW9avi918WHu
rWC9TfXFeAHGRtSka7hw6a/9j4hQcko9JPgJUJnEMWHr12CMN+cpUll26JXu
Hja3gp3pGnBJTE5PfcYK1WgsUa8jw7+2Gx0xcfmFeFQtC+MW95rVRBULWYRy
b1jNh/WtJ4973eQp0funAdwh8kVH9wrkWY1i4awT80mOOD0kepdZRLoSe0J+
SYXN7h/a3R3LvejtlERguA4UV7D9qoc0GTrcbhX1MKiJKCJq7187sOVg/Wg4
O32QNYQpOr9OnkvzI5ovWMn0d5c8GP2m5DBwzYSXRaCGdN2v2+TbjBLgipvg
VCAX3PRduK177TNZ3iuQDpOl3TiDrhao/cQeyKHOqiZdSS6GH859FSljvTNN
FQdVOPYEQf8AKeiULHCed4s4lP25Ef6He6bE2QolEYKSLcK+rCgRLN+E8xat
jl8pqXy0/PpXCDaexnUjDs9cFqLY6yxAm1UTGddvOHD8QyZB0hDnho98oEUN
5sK4Rg6lsnpYoPq24NZgZnoDF41JzwjcNsSmFAc89AyDlPRJ8hbjnvBmgkC1
TpJ1L1QGdNHVgiHdlyXdxEutuKgmr+1X47M22G5v8/l8hV3ZUNHkaHjrVUXc
53Hv3Y439dt8oDLqg+oi38yoH8HwDtTTGQ+D2LwPPUTQIAsnvvam0xQAqNcP
HpfCY6PviUISNSDpUSUN8DTATg5fuLh/DpecmXiz0HB3YuQpl8tgJ9fBd3qq
80qRvGQVUiYIbkcJtkvZvQq5mHf9Jc1kfQ4bmsGGPEz76K7CoBrnmQh1pEx2
DykfMxZKchu99GMKIQthqjWsDsp9T/SoCnZ3zuO0rg/yaWbZcLls4KMxJrfb
MgHfEECa8avzsC7R+ilm7dShDfCq8d1Z+CQmumDq/FHzQ+tKVds3uZH5NqOR
ZHLLqPvAxxvnZJBy4Jty650xVGlfTuqbTUYcvDVTN8uFSvL7RWJPWDf2D8Fm
oiVuaAtX71814crKzi0We6Aidp0RavkWmik6QOJO3mE+8J2aswZgLImp0oxg
Mj8pJiTLoK4ZmpwLdQ3cmzuj1OR7xazMbonJPIG5L3eyrjsIFfaQ4UNsC9kg
9X0pkNFD7sy5jU/LwbWTMCGND/yI467PpKmEbBpB0vSRCm2cACQgFdsc7QCQ
/4uFkMBVVX2lxLL/h3E/sjJDH/Z7jUGVw0SV3q5XUVHmSjBLmiE8kK4RIAkk
7L+xPCHzy+mSEGnubypHbHAWCIAi/vTdbVHv+M5H844mq1z7dFx+gtvOZ2z9
cyK1UpLs790j9Zhweubq9mnbxSVv9G6S11E5Nu0bFhrAAMxlQ6ofj9Cn7aP9
VGFPSrvwn+ga/XVodFH0ut4Ypq+p+H8RZvOa+q+HBHMA6k2HlxMEXCZpIXBI
z4uEiiIhIIldI9o4rQ13+UukLHUG3O+fd97nLipZHTsR0F08H90oe9b2nXlg
dBH4ZrRKaJBe3/WxOGRsJIAWazzXoYnWCPpDyOuSmwUKHVt7AtFQRKxRqZJ3
SbqzKPJQPvI85RVb8XWGuhPBiOlRyyMH+P3ezIw5jkjis5hPsHW1j40d0jw6
U0q21ptMNSVWH3hCqKCo3NAHd9BBlmcc9NP2KgT+N93W9XFOR4mGkiNa9xmY
hrcxreP+mzEGR6Y7Ufxa1H+5Nc9MiAfX3wRYY3R8MTwdTrlKDfgW+QXQElQU
QD1KqPNOSp9ucBaNDnab5ZCRBkxBMr/y9LS3JWcn2e5gimgsf4KWPY5jGZPe
Wmotm7a6WurLDdDKizq1r44gg+cQyV2XvyL0v+rmjmGlr3ek9BOY2MoDui/c
3CP2IGKvNpN+NXoP3lHWRfUkA52UFZl3Ac9h2VzIBH39V9+++cNhJa7aBbcE
YO1aAQqrXHUnwlqg+vtJgL/ZlLFYK02LPTdDQGIdzMXyUE04reEVfI82fU8t
vHiYLshizX71R5e7QLu627fDTmdBz5tPYwk4oqOcIpgZEGrjdKHVbgRJzPal
v40CPykx8KG9Op/aa8ZNRuwoLxPRXE+g5Tdnb+CIWQFf0ur29BKaV2dM6h0K
nzKOkf1oLqvk6mj057lyXvBETwE+sfFvYZO9L2RX3UdLnjbNyEAeY0KZ9z3J
e3/Gz/ZJCwl+lTaxOuil9O+D8x5gmvpTrdZurGM6OEN43O6ie785xH0NdWjt
cpnSZcOdiwYZ0d2UtkFcO7QEodsAgaw//KyIqS9CRdAPDOLYe2aKJAbQLuUF
IclnAnIvgpSuMJyfAVYlV/a4NJiAIhRrmA0LQDMO81/IVxW9IfaX1QVzLcEN
3Peyz5Qky8bET/A4VO/T0GHlvBNJ9drD6hthDv36opfAnt9/FmChoPOl//RP
qv6UYKWIeTTpYR+z4dOIfvWJyvQL9syJDqmS

`pragma protect end_protected
