// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
crW92rF9A66UZC1w7epNt6/+NzGoQR3QjeO7KnuwhuSMcw1RFhfamWRqEmh9pLU1
8Sqz5etv9jtqdzYBDspMkmtARGBpMU0EQv2bEvPUP6fH+gBlY+Z3x36e8fdig2Xa
lDLaeSZwnaS3e+wHAsMpceT3OJGF4UH8Sr3/fBsMiSo=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 5936 )
`pragma protect data_block
l1SDqKqOvF7M3EvfOdCNJXSb13ahnpvdreQ7wtyjnOZtXMdHb6bDLgdxLdnS7iR3
xZb7gWgpcnqKrR+GZwnqokv/S+XPXr4qEdCpQXuLlGrUJVpLDzALoPIITvKT5EPv
vAkRQitQClhQbruIaXGdGKpakPXLRCRR4Fe7r9Xn4hY2CwbWzLGWHPg/FUiffOam
6U6rnR5O/deIj+BEvqalnuUBIsPdNqQRSQtvzgwnPx4M7WunrB9lZmM3zDR91kjB
u8Zj8E1cA83I98xvM8JsKd29jQ9iEz/pVM2TkgHNKKJ8HfgQgdLx4rGVAON9Id+J
82roEKw0QHjxDVKS3NRwPWVyHw3r7XWZsYVvWHIbSocqD5uI7uaPdDkAZTf75woI
RYj8ahrIP4PtlcWHWhiDZWm38xbE67l0ppQdrdqqAuHfW1PVhPe0p/hmT4srePqO
Bmh5n+NFw+4qATFtqyk4omvf2jbKoW6p+VNNWHZfM4MbEngcU8fOeYPze48b/Odx
nFvuKMWzJX5tXXzTGawKi4N5571a1osF7IAavxGI/WaMFdedO2lQ9d6DDlEdvh6B
DrWj9yN7YozeeVZ0kveONNHeavemL3UBFb26OFLS1XoRypshOq1Anh9fAuBPvRB/
ywH2k6moiaHL1JZgkomZBCyAGFPXbvP7AdBmsPbFBZCa/+tlD/p7hsN3JJjj57ef
nAsDupkNR9MFQJaoS5iClT31lbSwPAmQnp6mFcRK4f9sKnBppJUOoJAHJ8vm+mlv
W72VncId59SEUvnbv232L8pcHPKogj3lMGJD6o5yFLX3uao06tJ6qAu5tFv3gUpp
waIf+k2zpn7rMkV2iiZpSp+tsQyrEdPKNI8F6dy9LIoq/v22l9RwxMGcv6dgmJBj
lcUPCbRhZ41urO1LR5ugzb3y33NwZfNFUa2uRsFnVSQCiYz3wcE6JAnC6YefftCg
nZiU/3JAp2rt54C29Bc2s8Qtdy1YG/ZbThozHzXqONPwjtSOebgnCthYduPrLkNh
zUdBT6NopPnl2yVYeUidYncxW6SGiEgksjy7+xSsCRjQ5kJLgyuQAP14A2sJ+eZM
IFV/c0UtfbA35taSLRoIxkKizeKwBqOK2mVy5i/cWrQhemb33qAbZuGp/vyUuKFG
158U1iiKNrHHPQFTp7S7dHHRfjYV2+je9JmlpCSuWuwo7XaJp22W3Ml1kydJfW+B
jRXHyTny0PCnEPi23kKMiAxlcH4u7BGwaSC1YnsIHKW6MEyv4qJ35tmOpQ5zuPNc
6eHWCWy5MSDWfxYwroQjImqMaQGWVcH3t7cypsGQtUV7Mi/QrCUUHbSHK5zJyaPR
zQg2IdlbkQAn3um1ewcUlpCDnI+GqWbiLpMHNCt1NvrS5wTROLj6rSIIJwq677r9
FA2LT1Oj/Jx1eih63tQ89qVkz1bwh/h9EAGx3h5j/qFMLHM9pZR5HDs1g8cmEyAA
sh4k1QCXIh4iWCxmkZinb/bpKwtqD4mRX/dGuhN2VnoSXXB4OcJHlmdoNz7VqgOC
025shKDz+r8GYOWuENhLgK08g83ZoDFKyGDDEDdoay7G9/FzD9pq3QBBNUxJxhyp
7nzW7tD6AbZvnMrOBAJv7Tqjl6/K/XWFdstSCNCFp7aKoQcfHJXefsKNbmR10GzR
beM73MuT+VyudMvT68mzdsgITnqz3HCz4cf8amsGGe85cCTox3GVddubLlz5HzUa
eMXI5+JqDltp/ykNntCnFPUcnpBVBXZ9qrxgvp2ey/7/ayQq4Nb0RD0OLhSqYFMd
eeXx9DWWGp+7YsVXtmrHmG2lI9TUzxJLyNsUuvTombxodtvnk76AP6RIioiB37xY
nj36YQ9Vlp7iFmMAj5Sp8wXnuovBJMgq8Z9DXLR84ZDEFSq97lJ8lRhwLgcbdv9g
uX15uDe+/l4Nesnb2rU/RB4hs38ch5VitRYhSh7km5w6nBc3yzwsu7h7icSgNHU2
G+MyYVmvydEvAJKAuJZejDEJTOsWT2FTso9Nc+SjSoa+9kJM3PFalXJQelNO4VDE
LEfU5hTEWrXkr4X0lkoU1yJMR0N2TP1vVh4Ok3/ZpFPUFNZM0xnD9qXvuAlOctFU
BqJBv50QztrpnPNxW8LMp0AGzg7hsikL+6sJtF35I8UT4mW9pIGpuoHfGaEo6C8v
bpJTXTInO6tx4Y3v/zDgQxXyinRyQkz8U6TCPzIRbEml+42ixtRy8EfgGJe5FqAB
6NiL/CxH4j1eDIAwVET2XYuuhcC0egNkfaszrcmX3wunsXNNg/1lFwBCEkuke4K/
djWejZbCe4OVoo/gYQPtjmmm6SuQ2woyG10jWXF6IPr+lo6eFHS/0QOdfz72T6CE
k4OGnzXXaF/OUynnXtQo4o+LaNhnPIGRCwkTP5juA8Az7By8/ICkfDBoKd/Q9Jni
/77Yy8XzkfYRIxb03VBPs+VJaZUfqiF0mVocE38/cW9BU2wSLbebytX2CZq0ZtvG
vsOtzZQbFWVybjzUS1goIfVPwkeuFNDXrEaGRUiOU2pKuDJ3GPHpM5xL6LiYdKsD
5om4O3FMWeNeld0HckbsOa1wobT3bEN5Xw8goaZEc6NX19J54qJfV0NitMhtpsLB
nY7FzjSavcfEf45W7MhEqkEnAmF4sOw0Deov0wawsvxgdi8AmzBb9qhDfoqKRJ8P
fI94D4yB57xAiFP5YbpUpEUbA/xKjmtUN+8EeFurk3NyJOicH0Mq6eHIb665yCTS
PkreaekSiG3Wyit+ZxVxfXYeZzkzIGwaLDrHTdH9H8tGDT96J1rC0clcVMrLhNsI
QAQ+LwK2UlzdvhUObcN7gE3aocUdbYFk4SKtkgAihawTHW++7J8TkhjJEWnONnHb
YgK8FveXj2X2vMWqAIslc1+dmLPG8DeIO01EWoAmaEYhAWlKQnZXeESe+RepooRt
/kTmojt/Z3/PjEUALSOUD2Oodp4zIELhoDOyOULsuLFfQWmuz6kba7W90Zbdx8K3
mTa8YoVw4GWaDuSuM1B69v96erdEFRu5hh0Yu6kHhSFZQ4CTL+zFvQ2PUYPmGbPS
obR18Yt+vUP4WzBf1xA8bhZc9LH2r9VuC3WK4kenHnRKOjc6sql+pj+HIsE3dYSd
FnPZwpds6/uHFFFwu4z/B6Yihj6IOxo2BgG7sBtnRU1CNP9B+IwAsviPmVbhrTcJ
wbpYcmxZIBcv+chvWjOnIm73Q4Jyi2chVE/yZBZjkjK8gbGlvDWvFdcakX1jZQFI
qMbK16cj015Jtz9+4N+pr6DVLzvNJna5X6Uq4tMZ96Iatg80wqSERTk3yntdvkPq
GhQPhMCCYPX6tU5fNygaY5B4FIqXONvU+jb30uYCSn5C3+0RuuEeiJgh6igyYOoZ
bel8ZJR9V1DqtHPUQs6Y8rVS9Xm3/4BZTsDYvadoFoy46Qp5gxad4mchV8XhKTWK
48YOJpkpQAJb1vGGLoDIb01jLquemr4Kv/aS22SVmvGmjU0MMnk66HEr6jshfCjc
W5F1BWRpAMNw9W6fvRgDLAoHnD/ZA38Toxwizawgnzfo5TpWYithCUlMa4FMoYdD
zFot3tt1KlmIxwOdBgsOlBBVHHzSaCOYQlUH4E6+G//X5O2qdLM6zT66oX609CTx
T3FIHLIa/rNXFpU+PL8KldZI9YB1TrvLMpdX+lYx5n+iDBrZuTZ++QveZQu+LLjz
ljwXLutevz84+5MKo+V/I+zsUN1697egDZgsF3VqDMdg5OIM1gBXceTe66NnSKpp
IUB5E+LU3NPpvLrbsVjj3OGfEZ1dJDUxeElSyfwbXFoVk7N84buBswcwCG4JTQvj
6A3FiD79xEY5n9WhlMJ0o37mZ+q0dPhIKyr8uK71F11Z0TJGvGb+isH2te9qPRa0
04LjiVA4RLreIXPGMLi24XNTd5lZL9ezN8B2gCB/tafTFaB8x/w8i2Km8xCrKesK
XNrfYY0l3sGBxCCafykn8uM3/XO7WXPOkL7m87mvZ0XReyzaMNnIWkqG19Buqc7t
iAoleL02yYAdRWbOqYQ2NWbi9ujJZ2ahZuF4naJ40bOU634h9yIWC223Kr9t9Gza
h9pgiJvknblaAkeMOR3g4wX9W/weVJ0CTBGhjO6tBKQXtkAp02kscbdj3jE35Z4B
b76CX6FQup9/2p8pPsnRAGFzJvL2guaKBZ2AEwGDTa2jrYgcdOtbAwS4iFag+h8o
6DB2TPnj8C1wXrQG4HTjOBMpmOb8b2vuE9HdG8TRPcBAEt1maxGzjFRRoXZBNY9V
mxMfoldFotdvnsTvjXNMrTVFkXk1xBtSW6bIRkrftsHUkbcKtkikZ3dAu7Cmd7Rw
CFuRKEGRyaOoZetNmOqWmPt2QPXoWcT8soR0TX79XPRpFv99SAAkv1QjRlJes2D7
M9Bb7DScdiYJpZgyuE8+pf+emDLyFNQ3Ku3LhwobZ6qVRw3voO1FxCcbkNf/v/CL
hBrU14DpyJf6VjzGBZh2D1AvQWZxeW44v0v/Xa3fHQJ2AApWt2O9qVwD20uiN8ok
HBkF+nOX2UAgZh/+YpDqRbgjDhkNaJHUE6RQqQ5LV5SqKZtRI3Z7Uc/ZZoj3mAbL
PtNmAzzSeYc6CBzKTeY2RhEVDjIxS+A841aSzQpam/dvQnI08/cPiK+lKjlhdOtQ
8sMTFOqAv9YrX9KHTcrKHHQSzyf9QIP54Lrss0fDO2fFd3GiOolEw9U5/BkZfXIt
jcQWUZDWY/xtZS3mZKKfNCX/gJGEemVK4UwVwHiYCrYr/CO+b3adhVbvxW2RxO+T
w5axrLGvld0UW5OEQZqImtQJY7qEynli/mlBi3heFfGPlyhqKDcuX6D0n6gel8Xc
LNg4jAfEhbPvR8zVndJtxvFOm6codSX9WWxDPFCfGQtAegjNkZsit6rU87R4JfGO
R4IY4yx0sQhpY9h2fxwydWbWDSHCjmZRuvF0ERTpor1oMS3QGcE01KV5sG94m2fQ
p9NjIhRJWq/KwCKXl4erRwJCRohPzPcccxFelSkzmmlhE4VjtCMXq2Z/x7tt570L
ah/s9OkbeNyRtufkhrpp0Nw/y/6mYLJWHfnqXBu8ll/aIRaMpstFl0v6aDEfYGbN
b3v+1eFZQvlUIpLxqFjirMKW5fQICjoEggn5Ol7GxqrRjFqQmg/Urnt+MkrmVPts
8mnXQgM06j3KMf/BsxUiGaIPLYqNk3wCsThMW+J/ukB0ZAfO7wPolqhLUjrZeJ9c
grcn+iuoCuCpR5i8Bmb5xESwB9VobMjW8Ko2+wrf/F+/u18dchuDzEs4W7V0xX3l
i6GIUqY2tqhVROKl1pDfgcCS1mcqEK/nqiopTSo756ChkHNFlt+3vBXzr+Oz9JYO
IS8l0q1IowNHDE3X8JZv2tFT/l6l2VW82l+H6RxV54dFZVv/D/CG60l8fZk+eG5H
ip2n79MZDMxbVqDT0IFBPmR62RQtFI6u+S/H0NlpOKqLmjjeqt3Uw0fhRr7dWkQV
aqadcsFpi4DHiZJbPaoMzrOEXrewJl4twWD2chKG/hwRfOUjONA66c0A/+v9yqWN
Q9w65UmGkdknOQaoNQTxBqoHZ58PsTU34MDqAaX8FTc8MgIga01exfMbDZDETDy5
iDvmYZBJBDdcBxx5hyRmO5oHkRZwliFQZp1n3VJ4pEWsY06T1wm4TqTME+UOJ6NX
WYkYu4t2laTkhf9sbk4b8+ZRwv00BX7QJ3K/crUSWqa4nkhf8H0ljoFppwiOqBvv
f4OvwrMlsS0sO/DtnGCF6s09f4IeuzgwJeNsueWuarXPIMo0l4QLCjkBAp9zF4dh
Ikqq+9xPqKyxFB1r6PXe+oIal8V4cjDkZaEzjPzE83GQOe/lG9dAWpP4QMNk3TjL
Q8D9qnyNoGzUfFXFt+K+B4ijtClp5+/USgUMS3AAUaZNIZ9HiZbKQNdabowbrwoC
UzLW4ktG0WZswCduu/7Kkt6bBcKxSLD7fUnyy0nMYZZ7LxUMn60ASTVSqaNPNg5f
5mVGO7CbUjJRBKnqiDWSyPbrtwgV/28bv5aKPsgXKDhhxC7ZRmQ14v4YX0AacBtY
sbjR1BN4VankRSLQvQLiyL9xk3BQzZVdt/xmxp9/VO6nwcJROCor8Qku+nPPyeEh
RrLODn9MEwcXhri974UFV9hxPrRsbAXE6/9cZKO4QrD5VPm5NvHwHjU7BpqQeHki
0bI5+eUN1LTqi1kfAMX+Prv1HftegdScUnbrk0VZSlZrXpcOePl7x6aKsXMb9RR6
MVkGII4X7E5Uy/FQyCW0ncNWQZ9RAiIrWoW4md9NUo2I2PpspVOL6WKIIIbXbtD8
IKVfW4isxY/Db+Tv6zzeasHtxPOx4I3ebeNP/f/IDTeGfutMEqF5aCHZds/Vut1P
nRwI+1gJOVWsYbIp4SQrUq9ujlprk9Ce7ssGL8jvQ2IZvPz+mwNRCUWXb0wWRVjh
EwiipHKbOBrvlzvyGBqvazvYE1Texwohvj8I/6PU25o6bG7oup7smg1X6bfirbwu
bn1ViDGBspek5EHfbmKyIic4hX+HASurQGz6Pcx1pCNzUpMf3syt/eg4tpuemxYi
IL0X5yI22u7uBk/CefmuMZGctcNq/XIGs/uFsIpgFPcANbPc2+fMnnzBZJNqt6Is
QHAp+2e+n8SxL/L48H9djS0iBU54dBZQNeC60S6DxYJpnVPHN/ONj3UV3kRtTVsz
loxAvmqrZ0VFmyS9cnENHZX5UfDxxQKbYBlERUHaPnYlwnrk8zyElyRjg5p8urRt
gmbosLhXXo5wt+JdO6KsmKUP7U0BpJbeW0HJXZXEH+B5bg5D6f5kjX3thmBXZ6ya
yZ2duEIJySie4nFzlMwKIKEx7uTROMQVOca3ZIGsPcEuINeaHxfhIdI4WQBfRatH
NCrKe/RbUKhks3AiNsZJhaFAmz8fAPE7YowZDCUwVf9hXO5gt+b1nVAqXPeYdUmo
V4DNPLyrH4P+nLYOLf3haaP+J0iKSuoQlfNVw16Hx35lmmePX2R3fTsIzulUPIz7
hn+HHYu7NsaSeNVj2mP0bOETlQfZ56ISyQtEYpPkr21qv7hUBjPZyFwNdlMDQLcS
MovpsRa1+ZujNUjyQEEMyqBVtzL3mG21Oe2xDxq7jse0ozC0RILjGH7Uqx9g/HJ2
9uuLaJhE9dUyYz5pCZVBmjmRcmRXXqXQiqHO935ul1dIzjbosVUXICriPIrCf3fV
kVoc+rFNTWQL5Lb9gUgXwq3mPoqrbhqmKAQOYIB64Dn7x4OrZZ9Lm+QLeWjUq9bM
8uScb5fOAv0ZFVd49qDNpPmTBDarI/F6RteqTF5SFXBzKVfJYfwqkioIsS3vQbqN
Ij4rI57DFkC/V66O8XgnwEUtBJuYtcpue9mwMa+NCujAM3UI8GkZTU6zmKcqv/zk
aEC6IPNXNHm3Bm781rfWnyBrG3ga7zbARL1KOP9CnPOERIYFR43AKgKptQlvJmpv
PlORiiBGXcg0D+cEN5HiiyXQJk85izOfRxUAFfJbdJK2n/FKD51cZvg2QKx3bbKv
1ecEDjZ/zNLKyheh9vcFY/iTBNx0woykKF/eMrHNm2s8RpC0xGSHCteSnnzR1tm3
fuS9PlKGgbVCiLPJiE/Ns/Wd0T/0ps+QHt4Ug6zD577uqB1E3V1sHD3Og3fRTaay
XukEZc64nOaxQguwmpm54Tz7ua2/OuvlgpmCaqkS+egMR15eKLdkKkF2qEG7AmHV
UandPdddE90deh2+KuDBZyXb6JpUJoasYDA8Yk61c2U/Np94RTY9fSEcKfMFNBse
YBRtoTbdV63UdZCpK/Z36oktdjtCi9T1n5Y/DAWLYz97jdR49/waqC1sdVNrJqeh
XJ6JZ0HRPiL7H0IElVfIIEj9k/fVVfBrQcWhTGtRVwk=

`pragma protect end_protected
