`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
pSXFFe7+Sh/+BH6pNruloDaclAD9D5vfbE94Krkwi3vz95s3WMgLJRY2kgJEn85g
B+NJ5+8MjAYnQUjkOLoC+cP0eZd2H9GNhjJxDXCNJNkgm5ZB4VQhtRp+HCkI7oY9
l9RdbiQzieD69DoTnlQIPjzArkXf4bCtBnw1LTS8X/8=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 8624), data_block
u4BO8mQrvh+OShWRb8r/SLY1kvX5gQT4mY+4WWQlBfCFmT+0jKwg4ctHY+KkcgHq
VWr1yBX5ov0C70fG4jxfIbERf0UePESt0pgE+sgjzS9h95u4Z4INYb6vcnJU0ni6
mwNAN/8N4yokEX0ONvr3NNTjNq+ujsdlAj1LW3w3h0REdnQc3rRACfNp1q9s9/+k
DjIIpQGrsDjcgxprmZB1xpELAEY548ZYEgTQJznhKnaMvlhwz7VtWHnFYFNs6NPf
pucqbFO98cxYRyAAYu13cvIlo97SY7sryLFR7XeeHW8eK0r1YjzgJcUfOP30v09i
87hK3fMHIgctHFiCHUCaCPE/L4hTFtanaROar+1QF3w2NRFZ6iFTbsUMXlPQDkJO
PoqfxXmYIc+NZwQ2bIDKMZGT89Zmz6tg8Qgt/l3zSHFH5ZwPF1LMKQ39ZREiuF9o
9t+Ecnq6jFNj8Pr+D58QUx/uYXSCIDhF1SKX4jLPTgCi35QUk7p0FOAJnymmWmZ9
hxaPsfWU4INSCJJnj/ge85+4NrXOTSLOdmv2WVnad1C+iqYVjXySok/ffqP7rHkn
VKBWg1Wv6AycyJLKn6wa8xmFOnIZs0O222VcZm9Nmgz5C26IJKq7xYddYLtzh/ih
Qh1hmxz7SFyUPCFXqtU03ZsOaSEPwZQWlAqI2FNBByuTBTR/8488RMpnSfbADaZH
C2ygEd0YEDHbS4EASD8BKbs0X9xkMQyAo1FxGi5LZFsccflNjehOVCtB5duMGvY3
5ko2FZvyHVqVYQyKcqf0k+WuIZJPPVg81kO+icpkMquBmi1Q1D0H+8NyGNz93zvm
6wxortl9JIQbk0Fh4rS5ob3ZZi9eWgOs5uzcNeNR2vVMXl0f64CB8OMoGNvmkDyP
91LRhjp/jSbYyoXXBK8NlLR/1aFLZWMt+tceUybgaVfiT9EesDnVurhWcc38Dofk
fdKMas8IEgodMrh5OCcbDO1PIAJACFmUR4KIzGgnmLgy0BrUWznaEJMClD2NKf+w
HZSClPvLJeFPNYrJ7CcPPmHPdbvgwTXf1HWaag7MY4yQ+3gg2uvCIeZbyUtDKSE2
3++NfzBWw9AuHLMNskj7Oz1yvz7sgEVh0PdFNiLEdn+FgEH81fGlSnDNtZihdFr/
StMdNEtY/COdsZXb5M+1wsWHefKn8ixKWjD6OrhMxAC3udOAz1Npe4m0W2RUHcUV
z3raobbKW3SYSjaGh0wBJ+atZGtg2R5Faz2mjUD3iS6gkvc3H+t0ohzLEkGIo3xn
j+mZ68Ndnzl7B4gm62TBMRt0IQDFSkd4ShNDPZPfJ5oMad1mZ1tsULK9sWCdULxE
F1i3Kh2BRXOp4pmsFqVjxIu8wNPF1RLibu3Ui9guJEKj15ZQyJcd4TFyDlJ7Rp8d
FELMc1fnuSvmwvepMuAbMquBDbR8eida2UR40h89r7buOzefCWV36xM0MJSFWadV
hOfR5a8jrI6jpPGqKPmGGoJSzczvha/RN5IVmlNn8ocDjJ4uZwTha8XnKeSUhWzI
r21NNl5oMHZGSSn9WuC8U3at8cnZqxuMHtMRqazSx01nJxW9BhTBGlBSEKT3GTL2
MuUGKszYuHZm3tfq+QHztgFu2ApZHZ3pVEyfxe3PzrKV1u3iS5qss8Hb6/7Oytz0
zzVHLawRsj6eqS0zX8FIdJviZ7AtVCg7OTbPVRrfzi/yUVSlYj/MDLi6EO+ssDgj
RDFgibpQX+yu+fdJ05BgvCNSRaZaCsxDOMv3OzroS2OtBiVLbUjpOE/hSBM8XiBb
cc7ysREovcWibNq+wv/DMG8HyUcI2XaTniv155UwpzR8WlTTe0prMDK6cEPNQpe0
8xXmbiurUKD5msOQqZO4R6Y5AOoqxmX/oJm69Lgn67V8z3CotMk13HEMYM57W66g
+1gpHSl5tK3r4pmMbWFAckFr6AlpBvRgG/dkwZYyNtvxTQBjIAWpe2qXJrUO6LI1
PSGfM2HIKSDY8ttMqoNvLtBVI98uwqmnbTFLS7CTHLcdl5+wk7IXc6zB/2FehIUI
QboCRtIc0pWn0h2WPr/Fa5ImkbWkwoCM41oYtsomx0jRDd84yVEPvgBAp50X9n58
Sm2caAJyRDsPCagpVTFVTdWXpc28b2UsO/ohEHlaWBkNcDOx5K9cIdMVEmIgKLpW
cLB4sZC6ZvaBT+s0O8jzP7inFeF8JYwFCnPiDCLaPbKzdV8DAD2t+iBEdUZlK1q1
yEbGkqkzvEULkcF7v5Qb+uf10OBD3amsHgjXXiVSKGEIfLXpTBuuR+wfTkMi7o60
gCKESBV6yzGBePudXNCB1UwQ2fIPg9JIOlf6FE4uaEd+P9woWZWPu/6NminqGTGp
ruRvmHfUb7NaZnwH0IIbt/6TpMnTfczQSnT/A/ihWz1lwZddy+EONk7TpCDznR3k
wxrldqABOThUXBFnffCx9PO9fx74pc5sYDdPa3dcbc2hgNF36fhsrmIIAn3KyOqt
QMl/i8hb+xWgkgul+WOMF5dQoJR1YLLPRJjEhCZbhnEIRM4sE4rGeLpLUWJvoDt6
RoOFUZyR8jA3ZOH6a3ERz4RnOi8MjakK3LpmlIEMXTqtFTuko13RGJJMJC7rkQcj
OYopQ03lLLKaa5kE5+1Jee8kH3Sw2s1YJh98FsigcBBre3AlH838kOwCIJZdLWhA
hUDsDSFbPfJv8iWbSDfrHpKHI/RhTWDTqMrPxuxkZzWzT/KOd0KNNqK33MzjcPUn
8e8M0G2FcJaVSSI09y9XUrujY0uwzmJhV87qLEGQSg9YYlLBPPhCDwW9bDE/PLbG
50cFEoOI8vSgtDTZkFTWjnx++ieMZA4O84XT4VZ6GZpZzhth0for4Hd9+mPuffzy
qmF4yECCmVKdzpNARMiS9O3bMQddUQrsRWexvLjYDYLa7k6Nl9dpUaAPvZLbPG4v
VJA9tR6CDuHbqABrj8NX15bCwZzv06ML7LNkbLxXuocZCcPLPJV4CnSwlKcXMn5h
T8zeOisfv3Qnm7F+S2Z+O1Q4YcYR6ueMI1V70sqoM7RaYBuY94JeOPP0v5mrV3av
NXrctPHXF/46zBUec3GcQ6aNdcBzvoNZTAvcvg/w+6F81DjRSs9jOEPkFNj9JZfW
inAig9kEFVYCpHPJqL1+DxtZOfrvCVN5MoJB/cycmh+X84G06hZBSEIe2B4ZxA3c
iwcmW6aHlsj9dUKYdj/+Ya5GDH9OkPNgxXPWHLQLwG7tUZi9Roa2PHATNwoxwLUc
T4jyJZY2Q1RNUWEIaJicSF+4edKpE1nVEG1DIuD4KZyZK5lMpUjcu+d3Kf7iB6k8
MmK40Q9+nBe9duFdpHg69CLSY5Mnc19Dhc5X4ukM5Q6Y8v10FB1hD0wCPHI+jrcO
+LgROEdr7DUQlewZkQIIirHgBINz5YSshrjmXZE0xf12kDR2Z3jLFF8lPrlUPHfR
RsgrC4H449A/NJJliNjiGaEOWKes/5db4Wj//7T3lDNWpZRNuiDXxAu7YSr3Rb8U
+ln+AD3J1xM09WV5ekotI1fji0Go/VDVQxvGBxZV1Qk+0XSiWEunEUH8HHcMnMZB
+ivPeJomHlBO407cv0842W5eFCg+/mg+emSFcFGsjEv4n5QvtQyHS4utZpMX71mI
4SnRz7eJv3Iqk2Wm6kG1WeqfkQEw2NyE+qOESUnzwiscb2yyXtlq37fraBZnNM1+
Uh17nzwmkgg06CToL3oIarCJ+THYrEABHsgRDXMkYxlyNS5of5kuKktniXtRcbXZ
CguHGxAzvG1bRrUdJicXf922xYj+QzoSfQxWi93FjUoXrbaURGkgo/kwCWe1V2ye
jGaqxmpaWYN30/EjveRUpfcKcivnyYn9IUaLE24GwOaCRF7LredanWS8q1d7fovI
DMlFYU1gjLlNUD6NjsbsjB1yvKRdfPKjMecRU8Czr70+OUdzqOK4hzzmzJJhtnE1
tFLvnRaXYiUIjQnrKn0fYDnietKX9O1U5qsbx0ooxBsfknVh++SJmerC+S4/SK9g
UYHb/AZxXxO+RpHYuvBfCZHqVcm8QuqhoxTuYBJx0yA+KU3vHhYzmJPIfb4WWbpy
Y8KS37JFmnQ5w1JtCs54lMj1M9t5g3vIOd7eLGUHWinvbXpLF+ETzrDG0iQdkptW
6BHrAG5QQ20aaklfx5KcwsqMDJGUlBr4ISKmnzBREJJqeUEdGQU902x4SspK569M
zW54QarEpHUk91uQucn69hDDuPwIXINczS/NN0CaUBEM3nMafAl6xzhT9msSwDn1
MS5WK6ZEDF1VosZoO3ZiK9Uo3b+pMtyMO56h7y9SZA/vlNllf34JtjpqSzmGa6Mx
hDtVXn5dSVTrmwAM8G/b0wWA2rvQH/yjzkyfkQ2Ge150ArsUo8bH87eJZKC0yjPG
727vvd/EEx6NPhWT5s2mScIgm+owPdltNoyU0ruQU1hjvSieir522VcFiucNkBlT
N5L++US4uKyqRCWjvaAYMx7pr6630NRV1rHSpJA31A0AmUGHOn/8XeLXbUBLgVs8
BbRYZBaDoFcd0nnAv0sQa2Et0MOue9K5wtG1JUqKYaYJa6gp0IDaykp2An3v6SFI
8uvth2b7We27lBNEiMVpjHBEIcRv0n0KEWyyH2p7Vn+uAmOQACFETlHeGWelKWqs
B53yS9bs8bBSqDd+0OX6xLV3kc6EUuWQ9RQg9TLo9VaoQGK8m029GamkYewsS4yY
UsVwIsmKSHsD/mPwnMhTGXRZkonH7rX5snD+cckZ+RD2lEJ3SNJ8f5Po2rjWTbvc
z3E+lJ0fi7td7zeWIynANY0Z7GFFJRVdTeTfkXp7YlYKS7Scgkcdd9+wQVPMrr40
qDUIvBEJ8iExnkn2Q6PHMuwCpIHLW8p6FIYSur/kgtjFBHetEmX1dUf0gTZceRTm
cdJgmOzdca5pDWdHQY/vCwwe4Rl9HkZUkPeqNCaF12qQNfcmUJopw62ingL0dyeW
ntHYXVFaREhWkl1M5fouoYxyeKOCFALImz25cerPw8f66LkfFLCIfdvIKwkBfqjj
DqNA9UqpkgyWg0tEiGrBBNc+VwOE6bKnjOGenoY5Qbt3b9FfJ4jyJBycvIDpNCAY
8CjbyWECcpcpsJkCQnEQHswrYf2Ko0kG2wCF93geuUyKkM2vcP2U4FOAh+NFqmyi
dIdGceapgQHgfIwpC8I6HfigD3fczl9r2K3zj4DYSy98xS5IWwFZ/WzMDCMGOhoQ
elHaYLWtgpp0PUA+GPAKqTxHsa9RtJeBLj1z5LWTNEEuqw1DWoECRdGMvDDMTxja
SeXbD0OUaxgYCu552LAkNlTftLh15ewmSzCEbm7CQ4a6IJMKyYgYCpX1NqwFcMlq
yjJp/IHFUGbRSWGHndflIs1t6etzMJkzZFz7Aa+Q0bDs7nfw0ETNthLcM9y5WpLU
L4B9mLin2yMy4IjJCVvdcU3kRZUOyj1RVr7A5hqqxZqY5wgS8EKXkuzGUAhrpHzu
2T97qksyXH8YkC7a5YnzKrXJcujL3GHKXnhc1vP/vt4rCvbwO5P/pGxk2aArE3lV
LyEJvTNphHX5mRu/e2N201BzTNrUrVKBtoiQXJ59tBVl9C+nnhvXXZ2v9/e/Gx7s
Op8NMkK6CnYuEkl9yoWoRx5GD3sR2qBrlPTgLMaQV6o9h1UZ+VJBsc84bQ6C/EmD
7U3sVGz+TDWDHAkoS5oFNCLCEd42TTscoHkleW3QY9C+YG5W2dna6FwRsgYMkvWv
yoeiOiLzR9sOV04mivPhDyUyrO1z/8Ra3Dh8VCce7TVtbzk3bqtyvr8pCAwxQihc
9ELR52UgeV0zPyAPtJMIv9d6c6z08zpzy12WinTJ6I6crxLQ44S2vo2jTapO/2l7
q19SpRqzq0pJmyi+5ohk88/UJnYWFHbkNJWaBCvmoSYnvlZ86OxSfAjS7/YE3Ph6
mpHONbYwj7whO6xt7lQHFuseYgHVZcosSCmh08tBihPyosyrvPW25muUf82cihy/
1KvEFMlCididvjtfhRw1Mh9NVCEcPBX3XPKz+4CKWfsmwoCyANiXH4pHtjGQUc4A
J7MTXdkIQrUhHcJZUQRxy8AZ8fi14+Kmh9PMw39zDdYTsaPfF2oqroVTtt9J8b4n
OCsgt4KVZpIVLmnJe18/ksU8IF1sOsGii5jqy5E50d9UvsyBnzI0+tTp9del+zTV
/KbPGrsDohM6KeGiOKSOBZS1O7aDIfbqgykrLglw7wjr4fpViklmqUweC4hPWKyG
KKp0Kp0+4P7d+PIVQSXEg21nWaTkjRmMLtNIdbcj+I3idhAzdBQQl9BpWoFiEM3J
K0cpVSP9zXJVT7fU5cjP+UFFLen+VVXxuOXRcVfrSfU6UPv8OAkVDChgP4IdvdJi
PPItbHaf+tg0Kx+7zjphkOYdZyJgJLotUc0LXtTN/tbj+iPGV6di/PSyuetAISWa
LfWiJtv4IQT59rRvy2+zuXLxm2Th9IFAeDpKd+QRluFmCulHQ0VA+cdCcNtq8oMl
i21u6byUDBFzlPN0PqJ7/FwBInJxBAN3QjNohbGmaKUmqSXTnA6BDSbGPUXP1DrE
0KuHPzv2NF2C74yYaTF2/Li0m3lJBqI7HlskTn1dwrlcwaw3Bxo7vdHuq7jUN8v6
WC3al8S48k7V9wvNIS23qdHYKF125YidtmpEefE+KNxTaKudZ5BzAPL1oij6foyp
Px5ihwahogE4kwRnVtqlbFCkdw3wrSU8zxAs6pW+ZZKkrxPopCqJU8KT9Wh3bk5R
oQICBQALW5lGhTOdZLTgzBppEk/z2AjPoAuv1iFO1jDb1AzrcazLUuW0F856I5kY
cAaNYs5Ye6YMArrWg6XmSlaJz9ondlvVsHwId29PUx47bGDfP1cfxk8SvpsBakcJ
WrjLetEPlc+fDrYhhsnX951LyEnkXQMfnTMPRKaxBu3RkXZ9qm+wLKLHms2X7/Yc
qr2BQuDC+6uvzMo4A1AwDVofF/PDmRRFDhEN76sVwXPKXimtk1QE2+Q/0Pz8GJtI
pY9fZh7R+USPPW0iepxLSS9fOFcw1vmDH8TcMUiZuNOoShc0DcWvn+8961FnBbWG
iKzAccoAQEkEURE40FxEDvyHYwYQ10r3kewGV2xtu19P5sFzlFbo4OhtX8e+Xdhv
FbZutVjGpn4pLpqqeR3ZPksP8JkQCubWCz5/9DhyC6PvWymxuJbrpak+F4ad5BZP
4liNWn/v5cHH6UU+PuAhTOo8uVXVqhpj0+hMth331NZy92/PXYXwDwy9e6uhW9rj
INYDepVwpktMcbxQE3CqlfKAisCL16F4wOGWBVrJxg444/lso5EGeOsZ6QA2NXFh
1CBqdEUGQWQneJIPBNk6PCF8hhnYhPRYY5HScdv/IXXeqNPMGvYFoNomioNs3aaZ
yAhe/h5BlCKbvm0vTcKsKs5gRkuYULzQyDd4ZzeJXdCgeTHfY4hfPhHWolLZ2Aow
kLfGvL2UKbBizhnUr+fRguATy44xHrBhzce/tkQXby26peYG2ovnN0wGrRkoGpPN
7/tXi2rOfY/EEGcKmy6WDlRCmIXD1nnfPfU4x0aOhU40hy3IiCn6diP/v+GZ/RJs
60FgtsQzHZu6P/seytui1DeuvrLv3heW/CY9HPWUvEZ22jyKcd5RmVh0FrX42qcQ
al4R6JHOwW/2H9EFlRkpYqTPuLIZcbvqiGY+9/HI2jcKjQDaiK+0M5gnfTpoUF0r
7ny2fmrRSAKaTF9/SdKvzZno2OpcyPRwW4cTTgcq0CXju5Dvwz46AR9m9BgQRE/C
ECY+Efx+6I29bIfhxejIT1FoKZnrwJzlyy/tnGTKQbjKiCmsM5D293kuBZ0lAt0A
MdIw+N8u6cnvJZQW/HXRNcDpmZQUGWn0fDFxdzTtj3E6Sr/sH6ihgy+yFKJJXbJV
AziayxEE6oyrgpdxnF+BxFi8pApHQEc204er98cF//g58xWp8klwCXC42z9nq2Ct
unP71yJfIMZoOhW+ggcbSLJRvVYizB3yMsXlU+O9JRZcobBUHLHFWT3BmwmdYtG6
FZ9/VxQ39xpAbNFd3V3ADlS8fCxNhb5it6rurWSd7ON7UiUawEtGsHYjRTDEuATr
Ss+XqcvWOF+afvylP7cu7Fl3xbOoNbWJtz1xg7VRufk1rm52ug/mJ27UpG1nyb0U
gSBGM5gCMj7rW9ZGWayveXLDJ5UgKhFr29F618XpEenhGH0Z3TOIK23ELP7l9kKm
DelM4MNH9+EPwQyjMWEbDpPe8mFTMMn+g9MPuMaGtVAezp7WfSI6yysecWInIIpM
LnnKcq6U+/Z/OWKINW3O14X+hgC3U7Z9ZmivBM9Rb0jwWtWBhkPF3FthdmLYfszi
nrQ6YYlpH2HZW36Hbey/5a4XtOzwrCgsiNBAa3PD6KG8+LRugjIuKfjtjbBJcgfl
3eTP4P0QvimIbzQT53W/jZOkmoeACeD0IWrx3Yn7JgMGyZVycgX6AWPBcjFaju7c
VXruI0bxGCS1RjSMhT5T5qVAgu4MG+O98IPicLE8q26r74WkXgfbvvYva0QBx3QN
EZd9KKRsDH9uqx5UNPWMkuASZkdPXg8W+YOc3m4uE8PGZoCJOEk5b/W4rncbKg5W
WfVZJ5+sDqntk0z6CGod8fR4rf1mIyPaX1qT5fyfTVtfVrt5ac/up3EoqV+vr0Z1
Z60kfbpmQ2AIoCMyPJ5jMPTkEHPoNty2tAvE41A6H1XWPMdVUvBGTNP0w5scKS4N
3IF92f5Ijo5Fo5Swk7duT04dR+FVRBXnq7rsyq7ePD9v2Aa+f/7UZGI+k6jSSszD
3aZ4TgVQObvin9B85onHfZeN+dQtcA6lSS07YdzeQ0CfNbkdM60nTcHirl9Q7WB5
C02tG58yn5xsVat2r954dnWJKfuEnBaU1QVXNtHDF4bLrjnXQVzlODcpqOX3XzAy
QMe7SDdQ+cD90rcsIHRSSl+5SrAjfPddbNAgh7vfWi8eGVmyCiuqFiVTlCtTPyS/
ldEprfXtB/mHyOIH7QuujjacirpreUOpM4XBCIHWnY7ktyWOKkRs7UkMtLMnMTb3
ox5aYEJ8h6mtVi50MKyUU98MaqIALRtO1HMtnPOMDY26ozDpNYkXgJPHPlNe0y31
GKxU80KgZWhBX/IvZXCD17s6TL42OQRLYMQRfDpOXejF5bknoiQNcFm8VlvNs7kU
vLBUQr/iHU0Er5xJeRb9PRq934mawbn2ntvECaDBcQO3XsLEtz856dXnfBvFZvsp
99e7OOFpspnC0fyb3HeATFoG2UD9svEhsSVH0mcAaXTb6PlqrH72JvoP2hTXUa9P
PIIOEBUIRmWiFnveTbGiDfp9/iiPm16kbjC2yiGvL4uQ/5jUuerIkTMKF+2r+jDD
UoG/diWkxZtLIxXDJm+rYyGTjjgtBB08uZbsVpsgpErbbUZeNp0VGzlhJUJYJSWs
kwaYtte0NuRFqn4AV3ErCdWn/hRj1GI8jt56NAOsVT2lpjaQFSeDJZurcJuiBHMI
pr77n+NmxNfxNHfCmMj2ZkD642cUoik19+CvQehuHRUETlNlVDqszTT19+xdEZY4
dsQ4OZh78sW9wVw2OwLF1wvpH+gQ4Qq9/oScWjocdB+XnTk36yfmdnTETxPx+IXV
WXXih0gWspXrp5EnA3ZATprYDbp/KccGDnjIWv/iZSWJigYFDuWNjovcJmuHrOS5
ySjX/nK2Sf0d32U++cYTrhy3wRNdphAmrsqr+gid6DPXSVKZsoIk5jUESiAmGE8P
V5OesX/cwUV6r3vmHB81yWWtqHEKCDE2BJdi/mgKwzRkDgTTiKfy2d//SLDfZYad
lKY/Bv4aOjcg2QHbjWULheh0tKbVS0iExz4caQcWILasujzm6ewHdTC7hJaqyqCY
wX9UAzPUgpFAtYEMQdtHqcXfEwZmulaT8bkUNDmouYAyvraZ/HyXnqqMmWxIHO5d
2DEp8dHxlPf141hiAUfefN74HTtUnArru6kyrfCQs+zSKH5b27dVTLq5fv85Prob
CtYSEtMqFlBl6o9Cz3NM20Br15xXlRpxJSykdt1KmB9sy7UBHtrVGCB+UhnqfJtx
mN8XZWYsfRnq0uFG8ZA8/pFJhFdIO8M/BsJUuFlAARAQaiZrwnSdLgAB55PzB8xZ
GkoYXJAwDFcvQGr0mFmM7oMUB/+MeL/Ua7mUWpt4spX8PsvSwp+hJ35jR6oBgN83
+Awgy3kEcHWa/BU+KDO7GLSTtYmfRqhXSG0IDSKNXIGTnMGaX2f53uclmb3GWTrp
KthhwbuIXUsSZCiZtyJoTZx1xZLhJnAcyvyr7aKT8oO+10iKh0dKOy/32PB3K4v2
f0Vn6paDocCP4FNU9v8zwfJmsZTPYV5T5f5/z1pKQAkeABuerynlUxP0tNA/wzhV
oruRROx9Zg6tCXfwq9+6DvIKAtoJch0A5D/YZHyWok9snnW03ayD1qr5j0PBECSx
xzM/xEmCOoMUxf1FWCP43nQ4+PEkDXZn/YJDyCX1amBEOA1TBXl8ufXy+ycgrr+X
RyiLr9sN4AwH5tMCru0fxRca/K05aumL8DSZpSEI49vSD5VZY0fPEJVpVPNS8Gya
HWUJNyyc3oD0m30tKC8A4pkLd/sycYjtX0tbZ1UsWdtvy25AYovQ1HpKkFOxKI54
hIYBPWXuyb7ATTCBmftEhnyaEWgcncpPV0r8J72HSnQul39sd9ZcsSTE7ikcel9W
c6WqMdbyIKZmKjEpR9DY3HCnhNf2cql7+U984+hKgfdTbgSHS5vnAM8pfCAQboE0
BGS8dZsoHTa5VAz46aeBflkqHsOfpTk33+XC4ZdY/QHvPIPY4jTW5hFp/+m5WfKe
Nfx/RxxelR/B4om0uE4mQtIhaAmQuXUo30Z7iIgMubF+W7JouSVd1ol7qsDWriR/
cc1axp2UCWDCKvwMVoVElYBNV6HdHy8pD5B+4yI5eV0R9+3onS0Qk6+kExppeIWc
2Wr3O4olGocgT6b1zca2sDwaMtPMDP/jcCQY7j0H2VkEalflREaUWA9wk6Y9S4j/
es8EhLSP0rNKAozBz53OVoMwrG108CaR6u5MRbCewYuImZdQSgnBAVmN0i8MPDfd
VFoLd+yCCFfiC5rs8CVekRnUM2K5DjTcZrlhLz8X6D0XHaymGMPF106fWFc0eEgG
ZFYUbRTlM9NIdONvdTXfacsfiHY/p1iZvtzK2yrS3c91x9bplm4aAQqqCfD2ozu6
hhPktHGhuczV2C5Soo4xYijwfWixIZ3eVxxMk+526iLknx/xnDvyg60/MrL+wvsB
nP4mSQpjjSY3S6ofiVaaetW5p0YUSLgebvjvzJTnPxz/FF9TQ5NfrNJAXqXTaGdP
RJrEKjpuJInOndJfIvG+VT5Wwa6uoEG5boNOEoeLmKsWBkv4NS3/ZQwYcJoxBzxn
l5b8GVpofW3SWxD3M2lXDrDbNKW9om/eUZ4Ruj5MLsg=
`pragma protect end_protected
