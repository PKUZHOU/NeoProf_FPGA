// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
0gYpJyymeTG3oZBiRezhVgisSPtimcRyg6jnkW4icSTX04LC6tooH/ZHMSFNFu5c
Kuz5faNinUHywW7de8MK5DjfOLCpSxthE3xHSyc89aeORyIA6lQxw0bv+66NYGrK
B11AoLcYPaRlIjKMffr3rm7bFOVIJ2rQOFIlyivqX87S2SCmn82uGA==
//pragma protect end_key_block
//pragma protect digest_block
GvoyL5wShc6p+E5pV0OP7vdt/4E=
//pragma protect end_digest_block
//pragma protect data_block
GjF7kjOcGKFOV6Mob+lvTuPSXSDCsmiSV/bzV+qD21nenBYl8PQN91KizCAPfJ1d
ih7fwtCF+bB+EySoMXi6lqNzM/mTdCOyY1MXAvMqeJP2zuKtom4D0c4ZrLGoO9Eo
BEM86BnsTW4g9+nuRR88VXBdAl/BZWE5OqIDZlWnnRw6a0uxL6QG6yPoOO4oIiTY
0qNk/wyC2jHhy4dNmbe51h0oa3X0G5PaK5OeCM6bisCMLmzLQhhba1Ar8/zWb/9/
CX+/2rgIM6G1KK6wh7jXv3U0XmtLsmaOkFYVHYSRwIaO3uA9qHdoSLH7hjJ+phnJ
O38RCcn3ZPglonRinCE8s2jKLRWn5EGyrDkWnasNs3anQBbwRAgl6+kk3UpbAQ+A
VuOjVB2QLCzM5IDOHdAslxpdFRJ/MTpRIsKgoMZ3IPk2QGRcaSq1GNOovHF6QXQV
sWteZTTirP8yaIfGhgXcev7QAbfLvI89nLuCnyDYD5/OFF28p+KrdpIliAOmmOeE
9kXmUJdpwU+6BP6wD1oWnJSDl5SddUgRgFJYw8/czqG6Sf/1446mAUTSiz/oAbvB
5lTsEHLXHhnD9mhBMLqRreBbmPpXmIGwqJ7nX6NEw3ykfpBMcEa54wyeth9JbYV/
u63GebrCIOihHbElyEUEICGGv58nwoQP90ux5sHwNe5kxOTqgOzggHvrdMg9z19U
DZ0V3tSwc1Gy84CXdJiNy6xxHb66kf8OBDweBRviildNrVYN9ntEZWoB+LFlBghm
9PmHVI2oBbnZjaQY1NT8IAyZ+7cAOGVQHG8E33hdfEVS9nB96khn9/7L9KAGkZOu
TBei5e1C+s5uWKa5sn8dNOkyb4hX/9RGmpSy2hSW/0tjO75oAjgz4bLQJQ8c0Tgg
/ILSVEVODCgN3AUIoDtC42WutFKPSUx5pCgCPwkttv6fIjGJX+Tj5KstbFdX3fQK
g/sApJduM+IoFkINjTupymZmW7dn89INqC6/u/yiIkLy38jH+7QRAB7FdIXD6Jwc
e343ekPOEG6XutJloWb/qLNcK4LXPdGmmSrE3nj5M625rgX6tnkUXyov4PfibZQf
L2eY5oB5QxWfyxS/85hdMPf7SFXbcp/KUY0vuc/VzSBOMXJKn2AHsuTj0Ff+K+vj
EcnfgNK74NyhxOgjdlGAxHtW18VrODdlHs8z/BP8gSsnoOkZXDOJApwZGs7DDGhr
1Ijhsk8Y+RmZRrJS3uLtQIv9b3DvKlJh4nXLnI7UHgpX3nH/LwsxqAt3BuJQsEKx
PI1ywMvX88BTTT1IeNB2dKl/uveTwOOveh++a8c+nIPEd1/ECEqGU0gD+MMrRrxx
/NkciiTakUXLxVhm5WTz6qVTTM06PP16bPCwVLGoUF8OgpfMh1R5cTD7lYd03lFO
JCtKjwIkfFPvFEXE9sTpn3K3MtMHkBfm9cHUImIB2wvMlQ1MiDT+kRqH0lzm/CYt
Wm+LCQ30cc1PeKVn+9cIL/ErgU2JUHalJoyQM6SJgwIuxg6L1QAqPhHTyrv3oCzS
tbjysXbndPGH6mOKkl866tpptd9GMH9C7eqPCpFj+spdGzpPVBp4UQalJroQ+rr2
O89ZYsBN8olYVkymNgJBNJ767tglGkkk0ZL1TUbx047/bKiW8k2dM0J9nmiTPeTX
mZkeo1LWwX6NybLMpxrgTLEC1BbQ1VKT2dTE08GTPRHbjnlu82p/gGH8trXgKjoB
kR8N5ZzLQ6/Q2gAnYpCH5CwXqKiAF7zCAigVkFjaE4OWQ+/Is5RPG2IDTfU6kNDI
b+VYI9UGgQq5YgjYvDAN6QEogfaT7RVHFdDcL8LeH0ePslG+YQf/wfETf5KosLYk
L37sVW8jt1vswILLqc6Pp2nQAYbyYqJFZguY5+L5RGW8xrYxcKwHtmWIIyl0Y0r5
nQUZD8wZjoCAD6bIFf+bl4Cp11ZLlFpc/zJvN/Kw6YEvrMQzcGBrXu3vJXOf3ItU
T1A7kxsVKKh6hFjXVhLio/Q83vzGGcRRQ66ohnjCjTI/tYfw1pfgmmKuk7ggSl5K
9/9wGJFKXvsUn3PSiw93jDRkI3rJ8vJZpjiNxcwGc/jGr4H2R2vZwq353rW1qi+2
rvWQpYkxAQJTmcLZSSiCRDYoZTuUV24kC9FxiD+gVVPCwXlxau2eSVXFAMQV6mvJ
FT8wZEjorvkQr+QUeX+ZGZsTnXYKz2htrQKT5tJ46GiqgQbIzKS8Xs8ANZYlNsRK
Ztu5vZpUonqq8AYhEI0pK13+bi3j+HVCCUSdF87P2k4g0vMHeEYXgecEjIKKhbRl
Hyr0n22bZUwHJrNQEct2lOpJr3RyduOIdjsQJ0dPDgDO4ZYDjhjTt3dvHlHuMV2D
xry628eTVO+s0pgMnqpUfT0QufC98k3aCcxDbyPK0jUm4UANTGzxtAKvWTgwQYvI
Oa6Awu0798oa8fiyibMij/1B8xvPPsCexOal+cJMsZqrsZUhMbMKjXw1yTrhY4vs
4udXRiSgaOOFryJ9epiwZKVRXSOib4RzamUnhtB1eZ8yij+QyIZgwLxaI4Du7Rfp
2SVOAvJbLd9ZFd/D+EKIwrIw9H/zl7oZb7mOEIDbj+GqxORtwpHFXie9yX6NgvI/
JumdhKewRiR9T9JfSdJRWojnAmUQhL/3vvS8XDCvpnAW/I0s/NRWkX0oESbW6aPh
M13KupMCkcOz56hUdurXBWCHvrsFGlj5f8isExMosEmsbYmIYG1aOmDZ9YTlBVPy
rZf3iWPqCOELjVBvelhjGkNTeBxDL9xd9EAnjtq103v6yRSb0P+vVhRKhyV0zMsQ
dLWqPlcHnZQHP6a8adgh3aG/z4tCyM5n9qYSNbqvcWRqMqkqkpe1pfbeZ7S0wILo
usmaeF9HCwIUphab/MLlrhY8KZagisGUAMWH32gVsmfY2dftarbM/a/E6uemOaur
ljziDSUISUnRBlZV4SC//rW54Fg8551lgHBd80xzjMtRLt2kH3iHn4pQg+x8zblQ
joCxW+z448u8S7aFRWFa9XxRpNlDD7f8cL+0i51tHeuOUhfTm9+mm7/2cULuAY2+
413wMeAfAiAG/6VwsvaZ0WSuKmU/+s2o9BhZdx0hTNXShq3UOey2OeJF3BhM3lJM
XhyaHmujo6MDYrfog5CbstKp8veJ5Jr5WYm3pqEITmIiq8SjHD1Ls5KcfHwpbcxk
M4ydRhEt+2Nw34VVfIDd5UKkAeuyJlzv2X3P9iOE+AoJ8qJSdKKRUqNPG2PGCDwB
krNkfu78CCGR/QTHsL5hf64YUKfmbUi+g9oi9aiT3Xn7ZZiQ7SWvHMpoRRKvNzE8
b2zd35zaGLnRVfUYVR0AGy8gflErrtejD5nDB9rVw0cVeu35UUSGIguijaI0gCTl
3I/LoWrkkZfh4Z6xEYMlaAwIP1GMymvwZcvQIgp5Wo00kolkvnAXPQ+0mCjedFiy
KiMDZshgLRCPoe+aancGD2pWeAd52gF0ozyb9xxrboN7DuKC+3dlnK0xsD2cGd5v
gscWqwn99SSij7ww/THRBgD/AD0RM6Ll1znAhHizVF9dYjMugrYi+6eWByIJOuZW
piz2O2OrEAkWya2fi+1BRQy4OTxuJHk6zgANMW/zavoTDebppxWrCRTAZxvLHLY+
C0ALgzMxDpPHSWM9UwfPnVHuNn6djMaKHAQ/bf9MGvoDfasm4f0HU+c7Xwzx9QBO
M498/IRxJhdXq4XS2xB8lMVijhmEDFZsNq8umPOgnI1VvJnQwiSSZVykuKgS/GeW
l4QKwc189piIJMqfUO570DFfZfXe2DZwEbmh98gDIMkfhOgHdieb7IFUynJ2jKEZ
1567u/H8dOi8n6gnc3C/LIbExSbNgp+5X9CDTvm+MbKzEnwhbwTwPHQi4hNvKXDW
Q/ZAEY+yMm9lRe9I126UOEM50A+BIS0Ty69r3G00Edy6LeX0s6u0sb0UZgOO2p3/
4Lj4nyZfen38FbA/ojzfdIG3Ds1Ovm/5Cpg11dhHeqtM9ifKPqrBznqQHhe+Vl6Z
ERKxtJ7SqRETPv2pa06KyWaNA/GVPq06OyAeSYiCAvLyDaYJhCVUzoXe6iI4RJ+o
7K/PBTZqcMzCVJk/hEGLtqHp3ryYasHomx+NhuAGWpAT09+clVNZINqAMhKoyqcM
0HmF2BW8PRwOjmx9SpEDUIe0SJrk3s11pn9Hcl5sK8LAy0PdeRfFzQfP4iroOBTe
KJy+9/yPWtQ6zlCOmnmAdC2B53MMttShawQ9nBxkpzRZvLbj2fTU1QcAD/JYZj4L
9KEUzHkB+bQi/0QswwmnW6V9q4hrGJgoglQJtKDMDDi4sHyo0le4WS7DmEgZGP5O
VhNUAp5iuya5Z7N+h9A3H46kAiVTPaQGZhEBTYIL+PX5VPmLdSYRpxeLWwQCAaHB
ZEjKpZEEf0gK1M0jMAXbGgRHttQ4OZ2/7bJ3YtbOZRIseS+d4EAG0m3lx9ebZdAU
jc9KPSWNNQwz3Wt/Z5MwLDMmQiHgVnkDBUi+lzQWTaBuf6saUj7XBtKaWWROUSuU
YqDSj0r3WVVMyu6+BvL36g6luA5LUOqBMUNAPDzWX5eOgQK3tg5ni3KLNOHSFUCg
Js2Oc95lTMGwcNbTo0Bot6meb52oiuE4knPX4kbFlOBuNjfQ6Dyum2QZqUwG1z1u
JWSX/+F2a61+9pKcNMVmUjhuadfnTlr7MH0HPfYt92CJ/jAVNwz8uUCr90Z+Ef0F
8OuA6Dmev8PehuWCiQlL7Qc0ImIzN/Ht7sjOf7eEG77dsXXZSW2aW7mV3tNAG4lh
bXSxVdJjucHFvr5xLQhj59lMCpaApjd6QQJsgvoPERqkwLRdEVwWs4NGAldQh+/B
wUmcTLzryRLCYINkA5/CdpATXuiTKpFzZMoAkvTL/DatC0iOnWTRub95XTB8KvB6
sb7EV9D5SV5jywXFfczAqZM4zqFXEhwmvzg9Zl8yHVmiqe1wrqcX5eYNBg5SI3hw
cVgLF+IfCx4ks2LQsPl2gEnDDYCUw8MTOnNyJBOw5+UPrWbR8qLESUZZEVSnZP5P
UUmfALqsdadI8EgcROyIN2lCzF0g4Sderz23RE+u21kM32upA0DQg1XD74Rqh8Da
PYT8lTsBjyJjJE5iPsXk4axFPuwCVK9rQHO84U1eUfuXnkysoXf2J62fPAfY0KH9
az5wxOxrUbm82I4JMDkQeW8CYY9IrQTBYzu+D18safFKu5lbMDbdsPd8fZtRUFSD
t2Q3KRkIVKP72AiRLNyHqU4PBWhwNaU8bFI3wB3N4m+MEXUkLTTtQq8i31hRR1HX
c4hmjLl3Xr/Ry0LIp4kkT2+gc+YNjLQnak73WoGqyn+36tgTG+5l2tvjmxR+yMSf
P72MrZINpEGtBaJEyJ3wzLGey+YngJRF3+pbc8nfKb26b2WWgtutSgcC+nYrmeI6
HcPHJrLhnzEX5oht47Ra7H/6GZPrav/F9delQ8Bdi/v7Q6KKjNHKtCUz+L1ZPgV5
hPT2JuuJOtuepesHGJcpH54EcV3UAGUSPzRURKlXWCU1ozMoqT521SThAxuLqcdy
/nJA3dR1dlcD651hyQi79Ii2Ac/q2Y4JnVzHjv2LPYELO6an0GrpQ9SErdn7UwTF
RcvdITMUgI6Ix6h+6/e6Ux91B0qNObT17nlz/icA6385pEYkAt0wo5StRD6yUoQt
IgwHzlXe9Sibj3j8gtwpIgY4M+C2cLzROIDwS61Jukvh+oySk9+go2ejUnjglt8L
xB4xlp+JKvYV6GiGeVkzHkssS6nADXaxgoiIt0hSw9yl3QGl7jXZDX5DGXNQZQjR
hKonibo3NDy+HaQt83Eo5ABN7wSSSPv9OrvDYKqapMKKxsdcM0b4jUxkoiScVgeA
67RE/nDgApENmPWB9rQGFgJB7pl8sReJNTC9mgZJT+pX7jB+mm7YAoo/2VmqAIUn
7w1kCTp1D6Xm9R+h3S10F9VGoDZTiBMXHEV72pkPlDxamhBvVZX0vbW+qOlQxKss
uuXVW2UxpyEYmZyzUNDar2aioqH8g9jRH6IAMbg03viJYSVvRyh7eU4v38/Rq8xj
XlitN0uDKSbizbf3IEI2hSdThRXPrOKzpVftyq26qfN2vNHCbqUPgGQWLkp9Loai
jRdSn1tsNQMYAoBwm4jOvf21++LNfL6ScpjMmWzOtkJ1Ko13NVbvX5UNHDPFTkJ+
wkBK1rWgFvdtmBZTXTnwkP7f0UKieYBcWKd44spGYr4+Au2RhSGASXnpnCIHC5BG
eqQPyAelQEjmTJPGnZJSVawoQzEnLneeFjXgu6/7SZuSIcbAdm+CfX5sEaOOge9/
rbr8D43CfRd+q8l1T3YWixaXDCHOsdPpBXh/SHj8oSPFm1ItnIgNplMfWRDXMker
vEurek9phVoLU7UzXVyiFJHgK1hvUhcPELVs0jNdAV6F4zoOnslG1R0f8WRbBDPY
uQUH2pT1cgX9S8LpGMFATBjM/SzUB/mf4gzra46lC7+4IuRBVjIFCN+pzeVd39dj
keMP0KOWopPiw5AvrAE3exiC228hDXOk9N+ioz7FDBlwE2Zx0hBpph2V/t7rBzsL
MBLUwN2h1NCA9vGto0/P0K9e+w/vEJMtisXiTOK7Uvx8YCfhMe7wifFUATnt1cXN
ZSE32YCdT7NPqBZw7tISJzAfMnw+M9zJWRU4wy3xU5nkTL9xR6ZIjqfQh6JQxB0P
JHXe4g8i+FlfnLWMSNImEVObk71wdbSZtFs1Ei5L2nKPoJQXtnSxOOmWjGRpLulk
+Dn2Y1y/0F6EbaGr4Ft8ibJSj2qVrSjjxwRLiUY63/5zz5wZf+g7vMhA815J+W1l
ho0GywirHEjqOQWIKTk6mWOnFyN5VgqDOCffPV2BVHYy5GPq+IV1w8JMmfRwr51K
FoPKdQIl3GhNlXG2gbJOfTxJsEm/UFF87UpH9bzx3i2eg9Q+quGFWsbAwZrFm976
nrkfnoTW8B0WNS5/FQAE4YLs5qEisJBv/efODmOYIM4mEeb79qJKdmh4bog72lb+
heXVq6fWG2D4pkOzv4vbh1XehrH5jU8aOPXLbKAA9u29yj4arXZv8xFgZ8U8bAn2
ap65Rji9KJnKMe19nkJNoEu9IYTfGjfsqbw60qjBiRzx+0jWPwNNIQtdx2oopzR+
C7IoTAnb/tAkqMVyOBMDXQJKm/rWPmhcqBdVF6ZjmBdDOGdD4ZebZP5rFP6NzbrG
24vqbGf/FzLFAwGWMJLWvsEIpRSkNjhchCVuVuF8qB5lLF4pfRzXY/vH/CbSGAzH
JHFn8AD2ElPQty8UxLROI08kLe2iuqYur0KrjDD/hEGARGFEXYN8UbaWjFChG8mi
SDUgIQp1QUdxK6n5qR1M4gfymTaw11jwl5g+MiVl+Fsuyq7/C86nQOeRTN5V+lG5
Qmn7jTCnQ8sVTWJJwf6PQ6xwn9ek/lE6S7+d9gnI0LJeHDYPt4JcgZVIF/ghEzQ0
viQyuCF95UikAQayGo9Co6wLxb6zLRshUxYAXFRgFYl3wE298LtEu7QlCyp5zHKj
yCN0RYJ3R4KhxOyrwoNQreIHnc0o79DUL/i/9Gz3aD6a5dDd3kA7EL4PIlczbaxy
jrkn18yKC50k/+A0vsFgQWaNwAj8Zaq1MCJ4TG8O7Ca3X/uACW0i7NpQYTm0lrhF
jD3TpLiDO47ewU2eeA1quozByetW7T1AKTclrn7qr3AYMDxoUQIgW2ak9vPYnEyD
4RRjz4mvdExjO8q8KqnoRm8vv7hmFtVWmmeFh93vg6Yp86+GCqA7N0G/9X2oFkXM
R6+4je3RTE0x/uixV940O68TPF7q1RyL63c1h7fkD+7umzKpUZwgwgeB1wggl2I4
7Zytu5YVleLSfD/rifc8txJCaut5f8GmJyAepDcL3ClAsGeiMaLjNtaUjBLRDtAu
nMOZWCyUwfBVI93QxKMLxLBwwN0oriP2BpAznE4p4rOOYWcJW5E1t9PvSUefeYYT
7Um7UFxFQssI2DqheWCG59qsVnaUc3W0LMnkkYih1nWYnJIersMMqg/ABsGBqPMF
oiWjkIwI5ynJCPP2T8CQcq58cQSVeilNkM12HVjKNF2chdCrFe6JZxPgz7tM/3rX
kMVFjLSPNbZkUUQCmwlv05Mz+j0L9MVt3YTt4/1nOogTLHvBqwadzohm00+tca9+
y+u+hXKuej4qcbbVstlXGO1cuZgp4khnKdTZ4kGaSJVLF+LqGz/O/1AYMc1YoM4Q
kODRjWj6kBBJhKIbxCF4F+5Vf3RZSaJDzF6PjvfU1u+ImmGZytggAgoEyfKdP8Pf
690VKIGJJsvv6KBLwzkQMfdUC2nDjYZlbkNgRP6Lgj6BVS02sArC3M7214AWQG8i
4Yy3FrkIeuJkLCOeQMAsC1+Yv3fXsK9Tgp2Jx20AqgrRMNRw/OXcQsPBg+KqC0PL
/FZb+53vrQRsBjjj4yWRWp6LgJu7FQ4+2Z/45DC7M/CpHRB4lY0/4FrCSRqSPx57
YqgMypSkCLLwIi8bAIUS6QFk532mEPlcT8TvuZsp5RMxiK56qRhu6nkhsUURcqrq
qeerV8GqBhX30ptY96kM2RuXpXXSd9WkXdQKmRiTBVRFqPCHyRQOAuPvz08aMb87
5mEhZp264uuqeq3wcB6fh+Zh1HWB2R1GWZacml2XEc6lRyNDlKWXp4/E9rpXSGc6
cLS3ukfo+Xbb5UTd6chH3PC2zThhNDhOkt7xUmbyszE0bGahot+HNZ65k/6GMExF
cAF7qXiWySE4BT+9p7p9m000FO5r/uJD+/uMKFYtc7FmIJia6tSzjplRw38z62kA
BCBdXKoB0n5fY877LEpj1QDvKYNK+DauyN77cpRTnQBdvZHv17GCqdH6VbMhUDls
sjL+bqiyjz7ROMviStIj3KzXOC05i5Uc70oQ1Km8mhZ8OXnc4xiBXFLWEQe8NIG7
93MoRG0VqF5TnQWTTTwEto/4RwWnic/SLKJUlX+MZTFWdThi2xdJwa0LW+eCuFxI
WelY3rswbcDQk6HDTzwY0Yki7Ir05KvHZ5+YDOdSfdevVcjBrKhVRLyhispTbKM6
vrdC4jE+y5S1GHt5wWFfo5yc1SNVg0mjjSDm8uM/a8xCrxW9Z+21d26GToMtwHKy
v0o1pHgnl4uowAHCiEvcOvOl1ORX0KCkhlZJVFbP8uDE5NkCyU+j44tZqZ4eqjRM
KEDrXnnwfBSUnKWlJaE/uJ4ee7fhGtSoFVGsCGvuHFgS4fBkHHDJZ1k/noog33HC
45QGSLXEF3cv3ztCo5EEdO9VDNu7Rl/SdGZ65MFWQUqwbhuW/zwJ8oGeA7m3z8k8
GfrvK/CqkHPDGKg/sZwz0TCrKIiqz6OfYYDf968WnndpmsyWtMxay4z1/Z077o44
j755XfrBJ6aafh2BtBFAWGd9ZjjhnNrAf+2OprYGFSs54WKRH9rVKhf8ZCqgLit9
yi6N5485vHQ+SZI1I+Lwm+T16W07VvNvN+gG6z1fG0lDHeq4giaf1N9nh7kTGUX+
P02+DLRKzUKxmTdv5m66ydG/q/rYPSPD8HZdYGdeGq2fQ+wZ/KIQsSDy4mpU11By
8pv7uQAQrxm4A0B31azRt62vfYKV6yk7k3bDXv3xTai/Tup0YErp1kbEZnb4YBvI
UIra5d6tJceR82z03uGZekxqPKgqVRdPcbUGiCggkgVaaxS4WWfr3Y63M8EXnw2j
guF8KY3Re2bz752dBXtzZc9zq4umZtcMVkEH7mHk0MPWkcYbJgY4UNcEX3mds+bz
+7k09H4wb9wuXo8mp/kKfA+2E9L7tpEADf/rDP6JfJ7rx9O2PGhy7VdGT42bxdXn
fOjxz00pjpqN0rXYk8gMcoOaEOwr60xfVw03BemWLfHcx7iL0NWebduN1TYQY5CZ
xMUl5z5QNM4p1/oBU+5Uz4rY3bk6P3BuA2P9A9dFSFs8MfofUkxzDdGZuDUBlC5L
clLJjd759L8hX5r2ib5sMLytc8tyagLb+kkdaqapuBnihvNuEpdDgTjxYQHX/1HO
BOnYm0jF9WvTYJL6iMRYsg+WmQYDqHSqdoCOmiR8p1hcvRyfVhtfl8REMcW9oJrh
gg6muGL0Wmnw6wkqGZQ/bONyTk7lssDs5GbwsdNDsR8SGdXxlwDQtvJVF3EdxsOt
7Yhwio0KHEbdmnPd44IOEmeDlI9Zb8BF6zEcTlPQJEvu7Z5fVnuuBUcJ8TcW1aF3
x+S0+IxrTp6PeW722Jb48OTfPeYTfz1+VuYJkBnk766AbkTpH2IZAuoC9LGzmus7
rwECQcIDXVGXv0P/pI2eXmEvkMRVvglOqfXQArERLabsRnokvv7zz3i9T6XFYgJH
zFyQ1vVo8mZwbfCviXvZXTXZ54XXf8NwQrlz+KXEuHU29y9xdGZ1U6PA8NCZqiW3
ndaYmPQ793f40iXkXzBzxzYqhXYz3ARB+F9OPt2qQaRmc7RgEbdpO085WBtxqYoH
Jb7ClrgeRnUN+t5rvl5a1beCFrGGuuJXo55V3IJggQoieQbRfERpHEzs/jQgmDi6
j2J+zZSeQkwPKTzhhK//KIFdOs9+Wgj9FKfXnBpGEODWhZz2otYdnX2JKWB7UTCM
j3qV7t4/R4gLWSaoN4lFl4jTWbSRhke9/VX2xJMLpI0YE6j4xxXlReNYy5JkaDEs
VQ+deeAtsoz0ZRhoM7VKt1Y+e4B/RHoZ5Q8W5Xthyln4i8um+0pAZYbAyK+w8u9t
DoD4VtksW8uysEh16CBi5DVnd+8qrMXWNyNCpN6bRBM5IyvnJgTFd5g4rq2C6+vA
S4gfyiB7Dv3qqFcwqxS1dA7dLC/XDytt5nWBetcrXAsQdQKncVxDXtc9r52mliM5
sAjOnjBjshh7+jZs8Uo/0RYcOpLpupvSh9BeYkQzKfE0aVSVx6fEXhy2pH3djSX+
kI69Z9Z2u1mLBXK7LhwTbl1BhqNCEFAcRS21hoWkXNBIuQ9hut/ZVDMxJztmCxL3
Nb6rzETkq63Hf6TzGTvCtkSz48GN6x0vAaVMzXoFPp1dcGdb2Rwui9ACpK3IZi2O
661CoNQMmZEqRbS1WwvuKk9yne9/cNw1kYi4tTS3N1bQnLm6ciTXItW1013Tg1NQ
8x0Xc956YV7A0nDn4B0NhFzCJQ+aNUDykArDmulWjitMEqXTcziTP5nFuEqWTCGb
IpUGfSmHST7qgNypcNuw4CbJcEwZClPvGmcWINlZ/q4IzjNXkzioYfFtjoPd2yMv
4TVrAewsX7D5GTk4wIWFWyT50sKgagvwMeurkx6l72+VRUKyQd345f7Y0VDaueYa
XFA2VdqmeF0YnmeMA5xosLJ1sS8vaGfjrw3zwtR/+z38TDpPWunXTrhMJ8TUxAzc
kxlgMaK0MJ6rPIqHTH7fwMTGr0ETPgpzjX7ieEC5KdU75Ui79/6FXJkRu6wBgtbj
Ux919d4OnW3Ide/bo9mC6iNIhx+j7k/J6btsuigfZ7jSv8XvrU7PVUEow7BhSu+E
JjB8Sgk0zJwi1ypFnEdbop9r8w/YBtsR/tD5EAtyiV2RR/Eou2uRUgzxChLwr+BO
+sz9ZyvM4vkIun95t3Ivxk8qqWzVn1DNa5IbHrPJwcjTPeqtHnpZ2h6xQjS9PaMM
9XDqgoNH+L/yrVMKDuHNWxL8W/PzhBCqV26GGUAdGgHqB9/y9S1BO6MEvmrKSJCw
R+8FctQkPuOiWxBAR1hnWh0vah+l+d5CEZ+AQlGbQu8KtqXf0vTRAl6FWy973/5j
iQWkVP5Qim+v9ZQdWJR+9bu1cG8YdEyw/cKxv+qzlqE0I4brxsOnsA/l2ZWQiD+8
lO6lW/YyZ/Ugd91h8bUI8GSKxCW+QiwNQ/ma08HWs4lGf4F+vP53v0yF0jXUYzVt
K0xQhjkOX28ErBuNTBtmSRDMKjq3qIT+Ipop17qNFaweE2QVMYsac9wjze/+FNB+
ZR/Iady9btpvGihXNQApAJsSQOfNAb/G5hlfmfRMAaeq86zSxFQToZuIh/6jB+FR
J268pLIMp92iqXo5WCcE22e1F8p/2AJ57lv06YJB2uLRBc1+zJBaT1GN/JmDKcJt
4n00Tfk0js7h57AH/58FIA/+fg6lwOiPW3mlBNIh/qCuBitvHC3NN0kHS3Ih55ua
ROyP38iGaXI3MnXTbPH5LGxQg0NkHm2HvzTUL/3gPfJdtfBZPQo2/QjNnx7LeTTS
eGgvEfnTPzZ3vj/wRhAqJ832W7quaNYxuAVd8wZDEu+4U7sptesT6+A3CEHZB++P
GKKVUYaghqfx3gPuewVN0Jh72gw8iq0GX2lmzKKy3wVbVBv7Ncv7J1PTpudWGNQk
L/XFd9ir4TkzcXbkwkAbpv6qn1A1vNEzpsoN9ysQG4jd9limxRphxU0TxodSxXPe
8Itmaq7qn1yK1ZLinFlreAX4FQH1QLwcU1cpgSTWKL9kQGNNmfCMUGFkNgYTviYR
r+eCXjFmaweRl0ssDF2JFn4aKWmEsUqTeoyIGOCCHglgorgRMQ8Zi38bowJtvvyi
QAwa74Uq+8x9hUltO0aXbiuP5171fvAcW4YNtFTCvyusXmh1qV44bfEbmp4Ko0sh
K7feOoDCW5hUZykv6a1Voh4BJstXiahDu6vIFre9g5DcBOMOOtjqLhW7y/KpRfa7
JzSKS5b6N9v2ff4YuNVjXkxpF6jEp6UkdPTZcsflM8vQ8Nj/anI9ZH77qHahPhOW
9WL79E/LDAKXgw0afDfb/lMDUQGMH1gGugb+7KFLyuePRyQvm3WOJcpTbfFW2QYo
0MNMPDz7l79YtLCnowliyjbFjk8OQKfE9bXn9jpdQi8WEepOmUVpnsmYxomQqM+y
PUA6fEtKSMiphZIsUNh9vvlradCTfVKo/2c07tHTUEzVBQ0k42z2x14k2d4/r4e5
OjRd8KJkMdwm/2+oniDseJKPYknjOKcklxm/93UDUuvysH5dqbvvxpQg3n6Xaz1m
9jTw5AQxzpVCkpTumm7kBnnRUCVO7eIdH3dChNxwo8cfEedOcPcdRtSQjxqCdt8M
6goDS/g5FSEhL8lrExZFiCy7zNMcbBboGmRFZFw5TvuDzUeGiMog1YbggM12l/O6
38vClJZVNfcfUvH7tiX/EmA+6zopb8Zqg+CTCfXLdBNk70HBxIJo3CLvyUNrxE0w
J2mD4yB3WbOzHzCqy0YKwaF64iizQGgIQYReZcWUi+Ysyc/UWQ+NmjUQCDzAPtf1
Ck/FEsKMQ5fQ9KZkG/GgjEFFqhGhPj9oY/kW5ZrKrhtFLx6hx34RnRf5IqRkzkn2
7sWBs03gi8t/hfRwgsYqYxbcF5tjtqqpNKMYG7md/u/aiEwGakGkHALd1qoIy0n3
1ENiV2uAhSrKtoJEAF865qPfRgsPMEYqhx73HBPxs80qXtKbx8N2lfIC5R2uxYAN
qDca+7vu0wjKdmzBjUeq1rysstckg82cnuN31HWSNva/Zfyy5ceuqWyO8XWtoHKc
xyabyorY3L0mFNeszAHmZK/pfuWE/fKgWsxemOEOr//M/0JgoXZ0BI4Fjg2VEnyM
an4PijJgvx8AMo7WsBCdP7auDYIrFo6uwlD85JY1YrlDzJzX9S+18AerYT9wjW4Y
qYjY3zB/kgIDO1r/j0vzUKHCJYDOP9O2QVOnFqkB1KUDBhZpM3LdXw1vNQIKlkdS
+D6BCxt6qJmxojBOhutbENI6d8ZNh1gQDYQwVkxEogMl5WVxbLGLyIgJXOrr7gBN
cQoBl+OuXOgjbuQVHco/UW/d14nvaGWZEyO5jdCtECGtFR3DJKWvYHcLahfA6hZZ
QE7bs/5D2DmnZJeIsGmCiWFGjg+yMLj4oIdZTAY9lYNjopwlXgHvyar6z/EriR0M
9l/vqQUtG2s3PtZ0mjbgOvyfA2h2Hybxwr0eS+TJYjEA8XQjC806Nyc0OaOe3DkW
Bc6vqMn8NrDKZvAg0DSVxXD2YIiZ+PZWvFtl1HMPuAODoLsc2bJfT7oTc7CkDudL
wHkR1ubsGT3dI1Z1YrBo3q1l2dZ/lSiRriyV+nqmxjTZGVQSd2B8K0tuj/QTrHep
U/HQd8WB3DdhSpp7f9mpz5wNoUiMTN/z+DbK1nZ4dpRXySLnyTT/OW5Azul1/24+
JdnGqaar5MyywWzAhQPz3uGs5hPT8rWWCfMyqO7B2qJkewA48r8NW+AXzV039WVw
RDyRvqpvJgp9eW8Y8T6tCWAEFQN0TrTVtfwLIPwlx6GWyXBWcIIk3uBJKe4pMr1q
wdu4P8ltqucnPL23Y+MpZP//fRkr2gxbvAu7IthhmgfwyKnCXdHnZOfizo+4p+DT
W9O5YXiHsmgoxjE6BDo3VYWVUQGQIVVAru6YoN222LrIsKkN9YrDSuXlcU032Swt
GgHl8P2m5DvYNEixKg45iWupnp3KedTsItjKt9Ww4Mvam9IIWWoUTBaxVWw88IEr
lX7COE+kFABJ9lU7tPgjm6CJ6EDZy71g43CYNFHbOadtJzh7iboOoJQeWKGoECWp
g/2qDYoKBW9rCfh1GvpbvOpfF3J1nRwjfHL9YlHg7sOrOeovr0YTUdqxjJrmfUIw
NPcmrOlXmEoOj9/UM+6g+Hu+CiXi6a3sHtU79K59aC2FdWRJGw7KUSPLKE7Dt8kv
KX6i/4vkAuR7qxMthr0lKlObB1LLooXSGkXlIpAXPJO1RCSSzFALGDw7OAGWseoj
ahhZJfez8bYPQk4hrzTp1prQKXvKb5wj/CSqNCpNUmXQ7Csf+i9FhZTc9GjENqlz
JRG7PvEe5lC3Ga/yPF2AKz5vkCcUjawxMcXXNU8JTGsIO0WIb7ZzoUYy3Jqt/V0G
V/MHcDp/dAfEJDjctSvi7k5gjyO6DpCst/AQFL+pacDaszv2pnDPmRyoGn2nGsv0
FEhQ7yviqjA/Hc7P94fDdB691GQ0zKRaxeBZQnlr1Gki/8hc+3IIHIPttXJT4Lp3
fN/uwPRF7NZAPxi95VYwwN5+qIJDzf3f3KyxRjPi45iXTpmSgUDWLassKlKcL2BM
zkRm811ysC7K6fB/JUCBpdBf8ZlHTVzSnt+8StT9w/fspqDKy4wsehIhYnriYFnB
KqO39aneJ0TSSv0rnWSwyNeRSQLtSag1vTE8kZcnH5Mi1q10189li3Hfx6qnTK/6
Qc4f7HyJ9qOFgjfXNFTMyHadqJiwCiuzlywEmZvTbtYQNwwtc1RuHkFI16E0Oq0H
L4tn3zrNnXo99THoNzlc/GWCCfxV/HR/ShRiOmbnBVkFz+h4dgtfXfytKCwCXm7v
h8XzSLqImvjF8IN27x3jJqMxjpo3GwQ9rw0uHzDYFo69ZHRAfeQdo9GeoWC8ii4s
0mmWaD1LVvQif+LrJtdfMDjAjIZnUVhMsFcHpIw/BbR+34F3RXMF2KktyRJiov4F
ejmFCLgT9XW2mn2PIwPulZfIDuI/pWXcYykxonhIzWllYO+AI2TrzprQ04CrKFce
C9QPJjmVm1WGYDug14DCi1EPksP4l5NQsu4KjPsSlJSfpOx7D6CyR9dvo5JdDc60
kcoqe0yjlrH6dCZSmpU5u/Q9kJtymErRqrQItGfDwBiwZ/UiaeB5LHc1wRgYko94
IYB6qnUNeqBl8bR0CENHov3EHMB+4qBU3VPbA/q90P15JbQ3WnmnMnyb13kG3RYv
sxlpaKMNOZdJcYj7JdkTvqiQnILRGHYUO13UfG7S4/lxnvf7hqpJbJXvQk6cYfpZ
ci8lkhaRCL4oQU/SEZn3D3gdEQbFpWmnqobDuP9oX11O4a7nSrWf9+vS1cbV4ETa
gH3l4sUfPT+OgvId32CweU/GWbC7Qv6X995G3BAwAedHPRk0CosTMxhoL8JyrT9+
bAo3NBbD0Z21Oc3O+AjOA92rBFcEFfq1fmS+6EmAXdugaMSBcbl3YIo591mJC0H5
M8zyvh+heKQ2+2TIndUoAvVfa4CzNxH+RuFmjkf0JAf0pETdvL1bTQrKALuD1/J3
4Cw82ML3aYdcGucS0RwX49YTOtuRZR/pzZ0QHlDZULQ0YVTF1t7JKrjTLHhuwkDp
j9YDinzul0qa76aHCgz3mm5h7LunI6Rv7UZam/TmVMJ1CmYwYwUIS9uo0hhHWHzK
vqCtvaiiekZZ0YQyr4mQ2eYqkn+oUb6S04rpCBKz84xsBOovwAG4DqrIj7utHAaO
+3Vxjvxigw3CXZgRyhBVh//Sa/WjSrEbLNNAcbs6IjN3rWsovKtujDFad8PGYRDi
e+hbS9pqzSJn1X6jCcKTFrSGvYn7bst2IDKFDpywZbSMW9N/nJIhn0i6EHAhfd7k
6h8bQXW2isa3z+B17x2Vbjbp8gmRQ6GyO0ADKe0281vflpgcLooexmcve4ihlk2R
toWVQIn8xN+19QnSgmDsLVf+y9L5F+dOoR01BlX1RHzMUXuCGCr/Hy3Ni6TRVOOH
uFjIny+CZsubfL8/v/4tj0ThPz0Q6pjQTp6DvSzWYrdV6ufiE8MPY7HzeH4pp1+I
euRUGJKSoFk1k2pGATpSO0RhUDcTNklS9fqnXqm6J/21bo4mXluGFmGiWW8rZZyo
aEQPxbkr4i3+be0o+b+OPbqxSb2lPGGK0yX+ba0PUXp0wLwW5BIqANZ+A0xCFAxI
iBd/g6gIAJTh19g/5FIS4WmYg59EOm5pps+lBAah1LBVfWD0Z6cwaWIBr7ZQZrfC
Pf3CtEXGm6OkGGllTcHT9uFD8BGO+jhWJKwzxKJ+ZPMMVAvJKK76ltc61wngSxlp
IDJTHadcx7YZFGX0LOb2IqPhJUV+2+1En/4htiAjoE4uNror/5pr+HSPpj+dFgkC
RqvsU8BJT9C0O3PhVHKMQI3VF49g6GCEBjUuK0H7+MEuzyU/9lINPm4nPo1LxAgc
8tV+bGcE0G258mgR4BGq3dzWql4n6X5ZWIxh8W00Y34Pb8JDx2LqEwU99ZITwpZM
yYkrti8z20xcR4MGZYXkQ3+N2cwXZHXfO6X3fUaq4Oix73a6MkMuvozq2vMshBMN
n8SFLKaIKot4Qeyng43Klejbsg+Fcu3+TDWbdKXoqG9iFNhLbDX0MPzQBG9vYmRs
vcbcAe7VwDLoIWG/WxZSkMn4f8C5aDDuc/122Ui0T8yBkrpljSe9G7MzzeN77q29
BI7BYQtJK4IGuF3jLhHnjtZj42CahxtZgxnIE5qgD7zjOhyxq/jYbPCI3dOkvwGe
BzdsCnyvP7DeiRVKIPnF+O9wJ5JpGzdeM6Ha8lasWnB26kgLeDhGtSc8T2lsMggk
v2mWpO7JC9o4d9FjnpDcVQvtCFTUguX1K5vs6r7Oo3KmzWF9rqm6qUQBB6gpBzyP
GXX4zdm2kW1vzxyVVreAkDfMg+GZ0akFJrg/NpxxrgQkVPlqv9X++EPcBrcuvQNV
GFnRowRlFS9FpegiQRusIDteSqvCeQQb7VMoRt09/IuO5JLdlm/e5KjREMri025p
gjGM/0NROFoWaAMKs4AaF9A+3s65ZX5T1Quo9lqXO4vBjjKstHeV304IGmRPek3Y
L5Dz0ivSSbeADWoQEUb0zdcWQMJkFd55jp1205gfh/StKyVw/BhIVcF4C0QFs+0y
u/XkyXkJM4vjyBh+SoUSVAY7m56MrkFe9X+r3DUOHiEPia4Ye/uxtDSAm6zbnG2l
j7EwnvQMzd2E5kGdHGRhfSqh7/um3LsH14NxG9P4RXfLOf18yzFtIo64tkgj5m6K
gipzV3uyn+a/20XipD8xSc36SkHrMJr0NoajOk+RnjZQvyNFzMxKt5lBFK1Mwho1
M21AMgbBVdDXzYYVxU298bj916R5a/2EPGRy/KDjKAKAsDSTRpePlECSvgGGZZw9
qj6j5bXS8nn7Ofme6ZYvg1anzagyAngCHhXThX39QzLhIDXIpRkgkFQpFtUAzWp3
ivG5dCRuxjg8l6yLwWvQbRAwXleN+UbwWm6CMLMfUrRXqqLwbgG3HzWeCtJPWAbZ
9OGJWLCJmikPKtII5Ybo/L3pGCnwAadZKbAytbAkaxHMDk3KvL+usssTtGsHnIUx
XGFiWtKOok0g7DJE/osD90zt63MQVWkl8hOW4uOXnYdbob39amYObFC4x6bLb6Tg
oLOWf021CcjfRlSuASwzCqa2Lvy52cfco9Pp4A5k9ERFzefUL15AdhPdYnxH81Y5
rxoJ46OMmXsHovyuJzmKOHvApURnXUXU2psBr4aNG20a+2I4yEdoC4bBPsP6xc+q
OY08I1yA+TDAf1mYc9juDnvKaWRn+Zuvnvfb5aMXGMvae6GmkpoHfoSD7wWAr5Wr
oZmn0Gq5/fZEP8aVabqR+pAQpMjH71kwXJ1xsp2Mv/j7WpAjJieYV8zgV2jwERmR
V3xUwDE6DmXFLnh90uLUQp7IAtU9Rlp+5rcTVRG7DdJpJK4+IGFfc/SypYZZpCzd
0PIX0W82h/EfR1MPcg6J4y6jJrEHCLZwpKpOgWW4ecGZHjrpfywJQqvvnaQpQWpn
b2zpse4z/QZ1K+abe5m+IXNBmQiaweKBpRpFJTi7Dtts6klJahuPzcws/EoT9DmL
X20/RNTl9foV9Yt0f2OB6uyuXQK03h4CzOeTvDQw0idgNKH9aLn5zLk5oGbY9LmU
vhr2xSHBFwGSRM0mnZ4AXRqjJhNwqknppOM1rhqnZJHdgmrCMsdW1QlHPDnX1E2t
uOB2PydZbMFSIKpZBBxC4vS93hcurNtkMlLaqTVC9jbNQdCFW0nKblmsorLApY2J
5ZhCp9+qk3HyODGH5dIOFnM1oG/QFaTqXzIDcTkQawKoROmdZPg/kPwx/f0bz95H
HX82Sje4YB2M4YvvihVm11QaHmuLbuA1HWKsN5fk3Q1tcevbSISZvFpHaMKbJ35P
qckgd5jlNIZ+3y8KI2et5mOkEiaCg+2SQUlPY4jwvAOAXLYnIg6fUgTZKIHzBN15
RQtsfHytmUssUcvvl4btuADd8goJZ7o9NBRSD6iWBJdzj4IjUsucRSfhznq3dQ5H
xIzOh1xBFaN9dhc7amOHCt2xZ1KL+lso7gYCHRb4345CvEp7Nuli8vnojlQqW+y7
RLwvjxUsuoCWD4ZK3P+caqvOZhyWlDPV5i+M7yIxjsFJxwmaBAGSqo080d2kVmaq
QdJtCmCD/avQUUDXYg7d6fKMjJQ//hAIH982qu+6/tXIgCsxm4LXNIWpfaBAQHAV
24wE4SLPzrsGfvbVfpo5CDL9z4p/kTLcUm52kzlsi+K/apa7zj/Te9V1tqTGnFK3
GyW8xHKHGarKNaxwxC8Ef01ILMBlatwb+N7OUBKg9805qdQj5g9xOdG8SkT8OpUn
o0h3s8kYSlPtghGmQ5EpMmInI1kobQh7U+/QbHLK+MFJz/kV3W6TjkAr625G/MIT
Sg0J9/JkyeMHuGBkR16mwpbEfEc6JtOIA0v9LNE/wAeHoHlIEex1AEvtlM7jeLiG
qLuPjpb3vURgl/YB+L2v5Y5VRQIzRBBR7aIyg0LFCVS/+vwFJlRlgZr16fxbxrZQ
iP5/gwI8Cj7pIoqk0+P9Oj1/qd77P5v0dsLmvMd63F84bFm8Fu1GOGQE/JI9Crp6
wVgCx+mhMlVkpSlKVB9zLXT2Px6dhkHDgPaABgtoNyd8fqP4H3mN22FeEaUmBaiC
WkCRGsm0GoxNVhCwbw1EMSP8RNQBAyNeJ42u5K82bnZ6yVh3/Yae5jP4lnJo/MEP
cjdYfg2QHwM4zLZcc/wK7jD8kXsV5O9E08kq31VhDQs6P7BTy4s/kSJCf6PzQIVa
KRdJ2O/VC6JgnUiKmQt03DvnXu1448BgIJF2bI51znqogHelhQ8Q2SjmE4R14itu
zcROGckCUFahahtIWrDbqyuyfqTrtfMxMGp6/z34PtrDN+dkdGTVyV7gu6Qbk3tT
SeLz4kZkgsOfMfUIW2KbDYCmb99ovuitE6VJWky9Rot8SIdVByqJL60J4BpFKlUL
u3uyVtYz/MpsjunsMBmPeCtth1bEgCto18/RBmtx7+/gNw/yVWBVoO2o/Op1unw5
OohlkJP/7ObjO62mljFNqh/fs4kxoXGAsTx81ZxWKICaA0Ch8tPr32rGPs3LcYjw
TIxOD4X72hndCOhoecTvKflRnnFNcbalUTQJ9l94GYjAYk7Cqjd3dBiemojnzkKo
zQrn6A0PJwQX5v53LJBoi9RGZKNEVCtSTDpDAX405+koQMeuHrBdlfKfA2hf47O+
fCLDdQqsYSpbcioMGyO5F7H+bTbi4cuwgPuONupa+UQXEcIjmTWSTaepc9iB0COq
jy62eL3N4Y9Y005Ba6iJAp2aY0CVplLOOS74bS6kPDsxHo7OEFid3ORGow7GEXQT
7n1KAn148dUJbOO68Jp+QvqWXM1WkFk13T8KSGH52PKx5xB6hXTgppElzOzTDRmV
13fa+Q46RiDJTy3/Cn/8wUwrkiA+4Lsxzcb0FYH09q99hBnF9Lc1LeBvDd8wnZv/
/5hl61XJxvJA2yzBlGCSCLvsCuXrq2ABHboT+eJdwjGk3K6fDt2vzNv4x12c0vSg
1CY2KeNQLkuqkjNua8JyLjS3w7GuMK9BjY9+2yZQylnyGCbFvNv0BacpWMgSu45D
NIrEIx40Wopy/yW03hLczEc5okqiEoS/Q/e/JsQbJTih4EUT4+cJIpsd1SSsqDrv
tjHskwGCZCnJHLjTI2g8EWggdjsaNVZf1sCzRDMRUbxHX2e8/QfZfQ3jRo9Tlu6m
emI+hh9qwCS2wLroaUSXQTb1OkhCL6AAZK35iVLCOURJF6Jdt6REARqcJeilpZ7E
s2QH3ShIqKigLxHj4ZPkCcah6KISQAs3K17N/4nJq8h26Dj3AXrkAL0ei/r4gVFf
1XAICgYHS7xNe1KbQRSzeFEku7MAHfJYrVRSvJR3btX08b1Kp4pPInX6y8Xc9E5/
be/5Wmk/Ed09hP2ibrYjXCsvx64WZgxV8CfBl18UBSXN2jowVvJ/fVC25An7D/J5
gRGbJdVaS6BV1m/q9lB+RbPsrx/uOOu7NIG8GTCK+uOCS2Z/mmGGh86K6WMpcOmH
3iXIB205mmg/NkzzDPbnP/8TCl+ytL2nlvV+y9168UvXcmdald6AO6vMtO1QHTgI
cAQsNYh/NFf6hQCXkYtA4Xr2KNrERMXUWrUaRVYHo+qgD/qdmjUJwxAT15ltG/J9
ETpwDsZFPWtyMnIEmp0BR2/fBgp7kvzT6i3ZMdvPnE8LWVC5OHy+fAEdXz4KXQWq
PKbqc+ZHZnDrIGKTncGRAA24GGB3TQs4NgrCzome2K2o70Qg43JEgprujKDHwwPu
szRUYXs5WWE+0QLu0144ZOkVt98mh/ohY1kzaSfUn1npPoqELDkpwVjwttRnwtCJ
qtPYWxSAfWwK8HCJFJrir6IbuMVF1f1F6lqtkp5r0K8e6UuW8Zr6VKUkxhx2MCMm
U+LqyQjFjoIAD2wWGaODq2yoMxi/F8NQUDMo66W7Jqm3c4eSl8WjdPgq5JjlcVd+
vKn/C8iTxQ10LrWjjJwtIzGSOmvbH3vdg+1SWCmzKbm5yn1Dx0B9cBRG5FrLiHV5
RAPmRq4Zq0kRl9VB1K9k8AbYysbM1MT1Fn8RlMPjAWKPY1/329anSHP3KTrIS2D/
zp6pl3UnDFWUgdI7wmCEx3ZZxMY2nkQ9eS60zBkvT4jlww+Im1owWbSgvcN6+fdo
stvE53z8PQMV4e0bdfxUMmN+3p30nHEWcTiLcMj8pxNZATV8FUbAnZ/1PNLu6gXx
DGxeZ3HyffaFkxA2TzsqpNzOuyiPchsxybniax/AW+9rct9VoV/V11G+u8eZXpx/
4tOOWSsAMrllF5ejU6xgyX3nF/4UbTKUGPRXfCoyS9W/wablEJEMgdbHej8zVByh
LClWBIq+fmTfjOX/UxIW+t24Ic5S29DKdDX1ir93O/2cJMxnRYmgj1xG4xW8OoNa
+HGzmDXpFs0KdwympcXrTaoDOZy6G9cKMlJ5L0VLPhc3+Afsxa4PXRDPB8GHJpWJ
oGx1bEWY/Swfqv9VVHwII5phyt/3ySFrXjJ9Qoo+oyDTBc9YCrHC+NJqeYDfboW1
jPkReDR3rZGgtZ2BSmIOaEQ5D8TyMHeK2N8+qKyGNuQalsR5P5otmWZqWxZEN186
mIIBUXJ09dgYCVNzBLKk4tZYFM61FyLuDTB6EbPNzcCfxQw4OL8U2hrkMWqmBl2F
gcLesbtMn/bziYICP2IQ/7bbS6XxCgoyX0JfpLbkBqMY9n/T8hbC4FaoSYvOqM47
Z07WQGtdprY7LTwyuoq9R1e1yqOiX5OfKTc4POfFDcouqNuSlWf03aaOG8uCI7K1
3fI8Y/uV3YDTgZHuO98Zyb9bG82AMN51rldLCtCxl4MoZ22QVXHJWvpQfsEiqZ/M
PPw0i1XT98KA0G3Iq3Qp0veL5mXydLX0l03u5xXXSJ0e9f9O0+FiC2EzuErSjPat
FoOlZL0vOhZRkNl/C3NC458h9MZfKEnG1TEbhdFNRUipmIKNh6oyknqs5fuckFJq
fq2Cvxli1UfjHUpoBVXfuqLuSvpnjdgNhLTyGuHAflsf2SwsvFnAYaUlnQJcl2fp
u+a2JIFBe/wgi0Hf4IRwFv/Is3UDNmhs9rMVNRDpusZBi9qC4gdMLT1lmYXnA2RO
BAO0sE4BJMkluc8/Hw6eV1/rKkezujlgMQvUDCFHDm9MNzxGee5Do08tW7UDbLwR
pULwCW1B3s3ljAfDFx71JVyq50djKPrca6Gpa+qz7mNPb2lKCc86LtthSuHmuDoI
5fS+E8dTCpu9JmHqXXiRNTPRKiM4LDYWMuPb9wrVChUdEJUaOY2eQ22bKUB8teMJ
Ex+e4FugKRqVvZs6SmvrKf1TAjqZop+QLKm0QYcNeTZdfCn3+nqFUpvaVgCFMQ1t
v1ihwvGsiOWbV+Fd7z/ODq7aKz8jRV8JsKidx0Hjzw/nstMKJ8Sx/9JmJtiECWA7
xA1Jb5N8B3W2yV1cSnLnhuuxsM6VgMO1RMUa0AKOAOcNi62m9tYyZYtB4cWyjtUz
2dtrmzQFo+R4q3rbA3Mj6zc8/x5+OfaYAgbA6lP42nFDpUr7F4Zv4SO6/wpmspHV
E8d236l7UOqe4hbLz69VvKZ84JqdbV+kzkozxkL/mi+6V31GrKYdDkoM0Cc4IYDz
f5mxozKCHQIAyXqkQns+VYrMLGtuZXClIdfEJyofY95FhDZZ1DCdRJMVnQi+96rh
I4fBPxZIYzDQgtnJF+fotVDI6hKW9CAsbdRQxbSf2LhBB4etUOdSSoUEpQcMhNfF
19BWhm7xpteyYoM6U8UfTox/JGi4OlQU0pX5oorw9EDx2/vhSfrKgrMcMXwVt8NG
jRs96fUHBWSxU0DFLxOFDPEqxGiAnUo/0LlKvJASBMNGBa/u2bXePMrTd8bbUCKy
Lirf3+2scXTYV+kbaUKPq+TigTA143EqmcLd5C3XUMw8R85vweJtcVWpyvsCftaJ
Jx/eev1GggMK42eu6I8oIe0M23Ctqqy5w2SCA4XAcWLLnVwMHw3rzfXPnB94R1nV
7YSqtqw76yQXnmkOvbxrGuosHPjpQWqIWLLuF2WKzqllxKe/b95337We4QUxDeEu
bkMG8HVy0IEMR14k8Q3dS0cdb+UFSBRQvr1PdxWSeQH5IqdEZE8JcXoLuf7RBbL3
14C3W/L4DNQevX7yxYgQqrMm4rnEkeXM33ZlTmybwo6RtkNIN1pUP6a6C68ABvJ8
EZl5kLLC955h2TMfTXWJ3yfrjg84ujjY4ILStYsxZDuySB4LJ7//k6X5dhT3K7vB
VRrEwBiXgjOOvLSd/hR6wc070gU8AeITgrrmp0dqV8vAWuOWTn12s6LP+s6fid+B
0kBWbJuhs/lQfRPbmsoV+JyC7CZ6asxL8fRH0bysNUeL5Hk+dhXoCERbQ8ulZCmp
PMIRXaZgE7ib3nJ3zaQwgemitlpaJ6p9iOQELA5c08u6fYpqkYIpz28ii4W5eRaZ
MiMFSxVVe5eL3UsEmp3V8m1NRQdZeqhsuXVbWLfLZp0n+PpvjQxwnQkqxrWecunb
0ouaYZcPUoDEimuWq2tXjCsxNQFpEcaqkexQ11rAtuGCKYnTo/8z1V/hOrO4A/b8
wX2c2BGTs/7B+Gr5cEQAoo0T//8vZ/qXT1RtPY6tpqeeVQ2ltVClPBy0ZmWZtSc2
2d3UX7aeI1oHwKjPnIuzbaCVa0H/m/mm5R6ll5by2Vv7EZcdSUunGvO/roSXsKhq
By8KNw25Fw560GnP7cckRn4BSKv9DagDVoVvl1ADig9GMsJhSUsKFBXTBdPaDEcK
23XSbL1Aqf9IYd+J1ej1GAnryyk1Ne7NdcX7mXR1btWvhvoPhTssDPiZGRi1h3yW
I1R8ytQktTVKpsCaELdSunw9w6Z1+K6NgUCkHSuz0OKd/kMDjEZz/7W9dQNHfive
MpzBJ9UEJ5EwXSbTwdKmRrCmKnxPMmyYKf8H65LnO+2KkBLMKQic7YobGu/3YJp8
roDDJ0Mt04pe797wmx/ykW4OeH17KWQM02duJVHXXp560yriFoy/3Ocu92/2FoyU
nXl0l2gF2ClIw8HlplbmhUOKVoBYChRNy0Yv3vrEZ0sxzdycN/+zxpWAESbdW6Lf
wOHSz22Xvvp8W7znucwdyuEk1+iM/5AlYz+I4zlxw6hmnwxjskmcxqXFXXuihmgF
1DQsT1udSF+B60fr6DkZNO71ixsPrjKshuuuMMZc/y5wAmX+k4GMGNDndxCHoo9t
yc9YjZaDbMrexM/7bR5KTl7SqfeEr1AEf5V3eDkas5zpLXgHAWyZma0TxqG4GapW
2E0C2BlBdGiKl+qGd1FPuOQ5wzPWga9SMjlJjKOy/7oAH27hUdNMVQ8mTDdUBgYH
UyimKoxdvmApFAr8uJC6DwkEe9Xh9257SvOENK89jQkJ7pd6bbXAeFCYfcRji138
4lbsQkjazi7zGQjIyxNJ0jlgglDLZk3iNJDt9/6xcG7XYElGp3kZg7mbZkCST1oO
gr7SLUCwBaQIz4H1CIvRfn+ubFflfiKmyM0GgLKYPTEKlHOnX3BXw6nfFTaxE4nf
XZMmFJEH+zWbqBMBFpPitiyShYmgM0kPwvVvU0+AW2M64KBnFb/oWYYuswhBMAEQ
zmfHS3sFnGretJRpyOqZA6GNa7zf6ySj5YPa6LRW0JibDuyk2LYCR6aUpR6MlsO0
4ec7PnFWIWjMR/QXa67FQD6uTDeEstCXqMufmpgf1QMAxHGnxr3ZgQ0o3r/rOXW7
O80ko1F37BHJOOrwp2YJt2a7vMTEWNzdyyS8tX39ElthNSajTo4FOdpwIF2IGjcd
Qfcbks9e+Vc4RwxG1Des1MY+7npBqcYucG8xIUfPUh3B+KxEcUzxbDr9w4e2Ncy+
qSZfZnjrxRPO+On73PUpCOIs4eXuYQbb5x/IakdRsC5+QkOZYHQ+pj2OdXrIs6cR
qyOuGYHNAoVfx5i6gvLD3qx6Zb/dWAkmW+5pYbCTzs1NYlFCpgo2vSOdTLmdW7Hz
6zYojCRMIozt1vjJthmvLp/o3fZv0tyi1HS/hcTVJjHfg9nSS7obkWYNx68al9gC
1kuIuhERdsrXe7YI7B2daTGgJ+uRUEsIxRlF8wnYtnU79cBwoxT5865Vdi08CefD
44+Ii0oC/1ycNzYuUx98lFszXVuJCZ5ckNw9PuFwltEqytQOhwPkmIP7J9rBO+vV
DDLuL/B158/5gSevdWdj00QsHdPrMfI0uXn+DvDRt3HxflCbIL6SoqgY8gqrP5Hy
q5pNOtbaT2oDMI6IFCrvLQekqswT/8PLPoh+P1qzfz5S903y4TbaHjkbIJOpdXX5
UkM6BtlFH8bZb6QTJA++qUyWwjQ6FGeSew7Qfjx2pOrNOvds9H7BHcizc9orLmEg
BOiuYfv83c8r8KUJ3feBqUjhLCnbOWF+9sOl1v3KXNlvYRoQcWzlxhUFOZiJoBDn
LbmHSODhCoaSql3d5STMOle8vWybQeiGnVBDZl3gb02p0Xvuw0Uw32c0rMecCvYE
vxYYJQ9Hl9TEDZXlNHz9+QLPjf7soGfkHBavnW+JVLDvw9fOiH8JzulXQck+NIYZ
Gnq4a1oH4XLIPY9a0x+ASmRh5HggKFR8Bcok/qwXUiPPXhGv+jUykaJGkud4X+B0
cAj64VTcpEoY3xJ3PXIOhof6PGEV9di1EU6RVRRHAlJvnXR8jzSZAdyqLtHs0npM
4AtYG4oa3HteYZ4o+uT/ovYI8qQGmRtdfL+1AJEE7+gUqvA2Z8QJTdMAZI2QigEU
YsmRk9tlnrMLGetn7isM7X9DAp5KoGBgfhLjcuOvKQDvp0jYSnr1e8+mAwbxwZsh
ncyjb+rTEh2yHLZ/a5HSVoG/zdiVIPtp3axaq5Q0BUH7iny4n7y2DaHGYqf2Bvt1
KetfuHemXQT0Gu0pKL4pn5AffzKwY52uPeKHpdnEWftLm9pFXUTCQMw2ppCV/b51
3Dt1hA5CX8ltr29h++o9fS0D4P+cwh1mrM7Hpk5PaDWYNoC1hOPQjYsM0q7q9joq
x9coo/e9H7nyWHwDzbi7tuYhHEelI5xvxSyUZZ8xpHI4cOaUTV7KCFIhtnIuaOS+
VgSEljOmWBOfXIUBSJOYO+8v6dBgz1uxvZ4tVWCrbwJdJaELUEjrzfJyIgOH2yWZ
FKhDgFASUTKnFzw5OOvWxHh8nCMAmJEiedYESXaleEDYnnuorR8kkZn6j2JxJT6s
ifv09txbZM5kIBf+iERlw84DgqYQjiMGKvnE4i3488xz3xMzYEvD+a4EKiVxMXjw
M72aoZiohdxCX6B1XLCtb4K9KNHtRlyX2lsSwhrbZdWBpbbPLYbaQ4adiMdhDEtM
RX05OHeeLrN2HrxueceGyhpn9GNoY1GY4D4ovouOJACyU49TgGj7MIApvcs60M6o
2RNklP2PIfDZ5QZYbsGQZBGUywWaMEHIkXdE6ULMYuVw0KljrNU+LapP0K/OeUAM
zDy9ExV7wImX0BttcCzMEXVnqj8NbOGDxHiNFiV4NmfAb2PokB3W/PWMXyxx9po0
7ELyA+wGeto3MOPxkFkoDwGqN9YAYZX9/pZkK/9hrNuQ20lPrQZLgpYo0ofMVGYZ
frlG2/+vlvQHaA94gQbHb5aIqLS0hWJ0L4wynjQNZB4cM3t7jqkuNCNmWkUVpqwY
/K6UU8henjJhjnXC0WrXMqXTK1L1ezc1nbUZsoG4WWVqVod2h0VTB2P6iQ8lAHo7
+x8GZjHEya8bT/93vLeWVY+zRNCdtcBSKMr980N6oEwLqIBc/Guk+suQYe/8l2W5
nh6vXXKr4+RG92d8/KxNm7zdNY6dyLC4P6qW+ZPwpRkBlSrig1HNH3dAFP+HIQkh
CClZ5qr29s8sAzqDCJDmLGctFz5+ue9vn2TDefmlxkNsYrl4W9oX7m7CKv41GRrI
+Kz56ZAbZAop71IVxTU/Dnz4AT7WFFgI9M79rqIgPWzRUdBBnECQok/cdplKuyYU
8O9k9M+FkcfoaCbo00LzrRo9+9fQmKs2Y3bF/5kjYqNEsIUGA6MiE5s2mObMSgGd
q/EcvlzBLK1BUcfsqAJmEpJsLlat8s22OHbYC4RxxHVUXjdJXfS2k7LSK5abCrqn
AxPAu/kyhMJEX21WFodl8axTPzDMJVHjSOWWEjpx19dDvlkLGt2fWMF8p+ZTl79R
iX+jTiEVwnwG/kFjLuhQASoGYocLW0KlfQXMgoHTmq2O29V0vDYhVeLxzMnUOtLo
F/kMHAes7TsApNQdeoe8+gI5WPm9xq2Pz0jJg1B7zw2DANS4b/gTsDGGtWizteKb
6E8F9OFekq5NGiE55jLPLupXbLZux38VGAc60xInQH299gikZxEH05+gmAEh2x00
63EsK2IGB2wtn+9y9njSW3kfIkeq4xUROB5+0VUiSSIr1ZHfwK4FhEbTuzfaUHem
xdqwc232Rqzb3xh+4cE+C/mwwOL3FVtnTYF+0vDnmufA9M9W+qAW6KtlrinazdsC
edSh1QTDGW41VPfh1H6ejjNWJ6d+qYO6cHJaaCEKnCeU933bkB3FrTzbqh3c7xfx
H5H9nFw4dgww4j9eYlHxeOzuXQDqr2wLssQbRB9YTRQHMzcA58mhn1KH0W2+BACu
C5HYrGlxfj0b08AfCxVKuDDuUOBw2SUWGn7C/iRp/fo6/aK70aDNbCbBSADf1hRW
O3uRU5Qf9edWiwrhzWd5kXd5sNns1Zd717mpaD6b3XMs9IA5OTBYqBjoD7iz8Y17
TWI0Bda0jQX4wHp5vrfINeacjAz9C5MLZ5H7+Z72VjSxez3/ZjM0uvTiLNOq1muT
F9itAQfQ/BRqyZ4sX3A578tlejt4dQQm0sStnGGXuPXiQLhvuGFeelNz6b0dYnlS
8PqfevwIEN2KCUlh13P8lTw7N62GST8KKcAHAYUH3M7g8Hj7xF8kV6gF6hrZysGS
knR+mRMfD043H7zHqc16Li6oiSqxiJRTFIqqIRg8Vqwe7OhBlHRASoaqMFDRwR1t
uQ82vyWbGRrPkoyuZlOxxTPj0jYtqhzaEq2flZ4mkF/Yn5ZJ4flFIGvDFsnlunfd
PpAtEb//URue2svIppVcj9PNQdhw/hGzlsxRMs8lGMgAgpwqEXZJ6TGlBA1ddCmY
uaJ1p0sw5guO0RN0AsU2DCpq1EX/VWiI8VpjVgny36703o+91CymKexcdl3InAV5
kbdXsVUQyMk/BAMK1lESFC/xQz/IdQO1sjdibV12kKgQ+/Gxqa+jIIpjyZ4ZphCo
kQhgZrOaJ0YLbx/JX/7qUoruahURflj4kIs3O5wNgbmqWSZnwOzFn4htSvLJi55X
Mt1mvK/kICwvtTBOI5Rbvh7mR/AJHLU7tsUfz9is4xvA0gGsWAvPE8Tn8Ddh+hiN
pXMEnixBP7qvYVvUj2YObgm0JvpQ9Hf7c/26L73OZ9+23PEBin4WO2NNQE8V4Wt9
clSSVciMs74H6o0//q2VVXMcFxi/eIC6kel/3hJH6g69BPh/cDkdFBWW3t2kRwwb
U0lne/S7q37qi8VsB48EjOC5pvDfHVmfXAjPyev/2sYJerVbMiW5vVfEMkJ2IgdT
Mrb8v2m/FhGztk13dSpb2P9nDT37FBQKYHy5M6oXEQN5lxOQj9xH/Yqx43UjCs8F
mtUduGnMATgT7Gr5ZVaQws6yzIAAfz1fdE8QKZKFIQyxeqogK2W6Lh6FP/H+buy1
XOKSnfYFWOL+VAOUWunsT4vrjyAYqv3CxUk8HP/532Z6erzSsvXutlH/c6qJKAq5
ilmE/6kFX6eX8m4NqXwaYS1x1LSGNMN3a5Gn+f36o5HiHqQXWZC6hrq+zpHh2PRp
s+i7T+wsUoQm4RsYmylLKgOWtF9Yhnorx4DkgA2hBbLbNR+ScpoqCeAewP8qfhoe
+PAtHoxlJG7OTNhSuxnw/o6WQONt29iDiwjUrtivBZ06eZBM+04djgqRCAb3udfI
C6PICSLZEZYrpTpD6JGXFOiTGsekSlQ3mb3DGMBqaILU5SVebAW5uXyU0+0n8cp5
rRw9OfhTSPoeHsF3xnJ26LhwwBPF1y5LZBBvae3IuyumX/cCUgFr37+Ze2w5poDi
qN5shdSG4XFSgMyx4EQQHE0zA0aAAE0KUi/CqwC+E2kX0Wt1P8Wu0KIwvoI9v1DG
m9l4Dm2V3aMYcRhPXWLvvdJw5GTgryNlQGQZtELqvj3EZCptX/5d9ywc8+J2F56E
Db5K+DQHSqKKkjU5dXtS38aSq2y+HjMNGh8x48cl9GNu+jbPHJfBdrNohb09t29/
0ZOFpG+Dwaa2SRVtCDmATIwJMigviJD6wr4OkqenJDUSPetOrT56O3NKFDBlZ9E9
XF2bmt6wUu848ZukKpy347PsREs/coyQ+CjnQqJGB7eNRqnNxDCYnJ3J7RDcDO/a
vAJ7gRVCiPfntFDde649KdyXFRguyvuSzcuxNwhTWueJgxABvBQUSENw/PLWG/2p
BKIWZwCM4ABPVhcRX1xEfnvqV3UtPjJK3I2PpTi1S9kFTML1GrASPBYR4uqV6E7W
9bGTTSPiWRJkvk/H7vfNqKu/I2NusiQYea/7ykHcCBdqJyTZBbGe0VflOKMqpdLp
nbBeaM3cxdsDT+AX3VoeobcRUbKNwIxUajKoJzz9VxtlhI6ga5aHUrmoWeJreeCc
E//RSybsy5hDSiaDkdwFqIGkiYDX691ziX+ogtKY+pp7FXArnsGSsZR791BQhsti
d0u70F6EeOh3oX+GzAMDxP9Ypa0sXxYrPWAwwAksPLyY+UDP/iObgpv52ABCazT9
pz/alu1TvxFwf91ueu7EhpUD7hFG8FDZyVRbexdVRjayKE1iwQLKQTAZ8sa5ncbn
Ac2KN8bsGQB1fyBnkuqJRBqWBGsHUG122P8OqwysmEXPAKG0MuqRaoUUzP69sLst
Szsd7RUpiiQgiWs5FbfZf4khMbjIoFCmEmq3cSdnlnc/4QOwJB7n96JSu5Goy6Xe
L1O9dO6PPWO2n47EREBGQEStcTdp3X6KQ9THLXoMVGBM18iknndPETJ3R924e3aP
Cpt2epeb1TvZOD5pspiCz1xNOTnIryKOd3wm2rBzK6fG3Obpz1dJQgNF3UqjQvdT
gA9HOjisLJfwlxoNxCpVNifG8Y1c1/6+9gOCzIPn+HtYsmGdlfEv1CGRbE4ecb0R
TYUyzSZDtaOXh2+EyyWpMREuiAzBmHfpTj148hbGEiFRZcF/9Me+267iDIkmgcoW
AQYv7uwEZSXBLr0IgORrgt8WyhObvBkd3Bhe/3YkcXRIrwgr+2oJAH4w81eVvc9X
ryJwu+Nvyt4GZN8nq5m6YwLn/n0cY2s+hj5OovagLVKX81K4FJfmhH1zrtG/41Og
q2xvW/pq9sV06Ff+bQWACqtRjz7KUOreDp5AtMF7X6FGRFJJCtyHPk+zpzSPyfe7
pH5tEgDVVPcn8Ot87kTHOpJL8SFP4JgCi5u4CZy0d/dCtb31jtfWiuhbYDeUDzBa
UFlAG61QqBzO4yqfJtkdQ/eRcdn6Rp8XvNzW0kmTQuZpKWjnpgbN6N40EeSRBbOM
hbe1gGMf0uaSjH9+B+SfS3vbCTE6gGSeNnUS6GQccc7ufWGWMHOC3sfhyvYTwCcP
9VtOa/hpGI6sJ8UhYS+SnKZwLw2JaTEmmuGTQPYxAUvD1ShpAfIEj6Z+NDSuwfro
2Xe7CIXwguWfmRgzXAYdNf7cNoGd3YqdNYnoHE7wzJb1OPTr4/kVUxwNp0mdZpEW
sMOqfQlNPbMVVdGIsCLVByftbGXKAfCpc5M8X77uVdmUa0HH4AwmjCQ+UOxyApV5
IdyGFZ18p6ya4bjhhMJu2+PExbSFrN5wut4xH5WL7U+5nuT5ycFLmOgz3OjgtUUm
P8TjO7OMKKK+ixAflc/Ko1Co7OwksBjmSCDkgd4QLPZybB6N94i49Q5c//HXWTos
Wfvyy515O1eWOvNGGui15+msA+cNLdIgdkhGEe7I3UOa7KyQXz4ZYxT8GyrnGGFI
cWqeQf8t4KOxUS9GC9lCrAF+09ZHuiOtG3rlwelMRsOZz7fj53exz2qz1UQIv59B
qxbQVNw+prc1zPn/qbOY9VpqtY44JfFVa3qC0lJofvboqf8Vbk4mAjM4pHcFOxH4
pS44D/1j+FP17LZdUrf06qVb+dt/o4msRu0Edbz6qzZnxx6oclNcDFtWMlvrL/iS
KyY1qxEyyt1LREbDXHct1emCVB3D3YUAjJHs6OojrQYfGotS4o3yc+S+ctG2mVUC
FBHXQcyBOfKeIc9P4+FOKKV3BAu9Z1DJj0lNflCVq31TWR9Bj39WEBwIHXAip6TN
49rcOSSofP0+lp/md+90oT7C+WDoCkbCf/1ZYnzFIIpQojAj0acqL+iGuxVIaYqA
+eA/DhRvHv88SROIwP/ZjI3CVaibCOfp0b8XwOR2L8w0t29H3WX09riKSYv60qbo
yc0jshtMYROk6gSuRFHdR5szbCAD6N+PcB4rzOrwwG/43XjceDY0AC1lM9QiPBRQ
DsHl0Trqu/2jI0Z/Taaeb4rEuwDBGwnBgw0fQ7Iv/tyWxs8voP2Vz21YokwPI/5I
LQdsPJwPiW3iUrcwlLOCQWRXNKbTmKWnTeh03wyUqmNay/Cc2xWALk2483tcM/Q/
XnaKFS8RwAMX0oEKmP1balultGa1Wgc05OPWAPHGCjFBhGghMNEaDyVFeGJiJgIk
m2D5SNKbCtwepBcRXOgWfwttr2cxC4GwoWFBJwKy48/va5UlBexBMF0odwLQoTYo
56G4TRKWP91x6ycEK1qyV08IbVOZH22MtMpwt9+KSur3gaNpaqEs92sl1K3ARwii
SVYpiwZOqkC3aiKnOBH/y/o72hK67annY3fz5+jaMmDb12xIAwX39vbtYhyomhU0
UFMQxDSDOv4Vg5tQz5iu4Z4h6GpW6mW4g/jEiIDRku7arXh62DxCPAKEOirBN5LR
ktZDq+sUhBYBl1ipwaUOcgr+oYAOhJn2e4NpYYgWqmWKyBndQXWrwC4lmaGjsWqa
4mWJ1hHoXX/dpEZAL8ZMMR5lQZO9mK2Nlu26GiFubzod9LQDJBxZxZZfCq0QqPsi
BIKGkSUK9C+Kx6Yg2Qs/N5lNeJyMYs+wv75sY5B3nnlYbghCwdKxBkKP77ajaQ23
TAAWvJQ9SY4ku5AkVIxoYlsul/7FRsT6T8cHDTJ5gvu8gjIuKnzN+ytASiBmefRU
w+8K5e3RqtIzVFiNMiAphEi3fuHDZaI8cvblyEgXNprCgnA4ULUVUR+565JWQc03
pSoOJ7r0N54Gw8Kg89OlJpxm4QEVQodTDnUhXlFciko7qG+myImVZ+Hkinn/DKuR
j6ERFIW6HfhLxwC8D5ceMVLGZf6CWCSts/CNUTgiRW/EPbQG5chBf3y+NuE3aWGc
L7EImPC1RDv+rIU73F3AlEvy5ThoqvNHbkTMhvfZDE1iYM/Gj9ZhQAWihAiyOrY4
AOEh2bAA9ELnzwQCT4GE+ylDTm747mOjVvbHBWkt9B3y0PELxtD+SidRWUZaxehV
Zl4gIykoTY3OOvrhAC4gPgDUti7iTp7V90qs3nNXRra1fzoGHFe7lZNn/hmQ2QNL
FnTH43p0oWgEmtF+K8MFX6m9Fm9JDcrLhe7vbnlGO1C+GRFHe1yyh+g7GvxMquNQ
exmYUseOu40gxKc8Oge941r5wEFeX8MeiGQUKWXkC/T32fLqjVI8L8UoFSQXYTR6
8eUULT8OJkjFjKnDCoq+gsPheaZ7/k+DzIbjuB1+382cHnQXvA7jfTsdkVfHS8Mp
fx0v3KkBkynF3eJIMrHqLKOFAdBbdJT5D8NElPz87QmSfLdMxVIXxkdiNChy5MYj
KkMS5z3Gy491D8+kruBgRhZEVHicRkJkcMSGL/s8DKENe/zRnLENvEZid1ewMf1d
nSNil4cfUP26mRP1Bl22YXk7hFpW7FVNeKX6XAdqAqweFX6hqoPPn6DOqO7yb27m
Tx3kNXbcBQqPFdmkVs0PvS2pn52NcknzbWl6BsFGgwu/+vUxBN3RE40UPzsJhoZs
iIQEgRuu4xS4HzTZmoHS4SLMTm4rM72IC1RTgiI3c6iapmBThVoGIf6Dwj/bzEbi
Jaj7HiVoaLqepfyPL0CNX9s3swS3vIpfKdRLLB2Wu/4vrhCy1cHcV4wnYRZK5xS2
3uba68dj2beCQAs5Uw9ON/vp+bOlkUIvYDT9aoM1m4qB+12zIAZp2I62NWFD0Zgs
uLSYrkGp+tZql447BFq6OjYJFUqJzPXaR6jxvxkD/ohtWvkaefsy5vl99TJtg/1k
O5rvmQf+VQfgSp26DDQ6bfVorsvQsKeGRYQhDlHA5VGoK1NtQjypS+YDwSNaVvOB
Ka6jKVPFn+saJykJ0HQpfb1VXctxvUDvDRmihdlVZ17M69TooC9We1U3rp9crgoc
aqA5A/NJQA0FSviv2kwexPcbGERfOfzHds+EPvT7kL0JA5qlpCGxlwUhaPUszIll
lPdaWaTF8aDtyEZbQzlfoti0CM6rYTZOFSiUstsub6nKUW4YX1ztW/vcOWSzM5zH
+5eeU+ex2hsCDQ9GoED8sPjfFF1wfzFiKm+c0oqzanlfrS88F3QtwyGOXfMiHYGs
Tte6VKYNpNNmvP0G9H34ZzeeinjPBzyCsAG+zh5UOvbgHYv8ARB33d/gxuEcAxux
y53ERLFHXbArvK63Zpa/Ge7oX518RMETs49qW3VNoMnjBzUyxIhdHjJ/zQslb43F
iVKgffo2jm+h8P3zkZIVojmbFNW1S4XkXiJ9uBcg2SRm6HFxCpJsSS6mpx4K8EjJ
csdI3YiZHM5+KlNzS+i/9OjxA0+04RZnHMdNqhxyPHgd6ROcdb+XEkWiD17D0dNa
HuIO4GRNfGTF04L+E/bXtihAa9IImLM2VO98Q8uvzvfT73olLWU5vG+1bmgMwz7S
hg6WXFQba51fQjp5rpSR4CkdlUo6SnJOVk0SWT9H5sGx9nTiJ88sEMwZ2hBXU4oW
w/JucgOhBY7IpQaCWWudGbfYHJa5ycReltt2Ffbz9CzSd00yKkDUvdH6PS5eznf+
o++f5HCNSxkreBfYPAXvqSOQvvUXZu2R6Ym2miceGY8GsAWPQjT1AQFgpOqV/xr1
m4hIkMIyJRIKV+MLrhNf3FIVFBwsSq62kaERIa89A0hJqi7+sCeVf2LN3UMXrTy4
u1PfbAJ5RF7MHFLq6CSUcjnIX9YI/bIureRyY+So431XQ6gV/1rqGKhVZo0CU4qi
t0dz9guiUuMA9rtNmG3a3KnKX9kupZ5+JOcktVVLcNYxIeZ7AMezkthESxQkeXIx
pdOlSnK5PQDR5FDHjFtFg1SrfPsIwlduwSFDGwHz6D8FQYJ6kIweYnCwICigo0w9
raDG2DuthFzvmlxhYtdVwPC9UyoD26tWFRl/CULcuecgkjT1LiLCn7FCrAylMBNX
LlydGQRzydXhpnYPSscVN1ZSBRQ/RbvOQqCpYQqoNudalCdL9SbCnZLtFa8fjYCT
mk12/rntz2uyHd1ID4TwfWy3MaArmXi1oduroaINpBd4phhtSGyDXfG1jJ3fq49u
BgjVZVQA7GAwgLI5mJuQKWPfoHWoc1AkhRvsTd5ZN32sFd9NEvCokhd4pKs3Ti43
GEIOUlPrMIWowFnA376bfDBl4z1D/QV2qbXsXvQL2kHbVBuS0SsUunm/iaPUgbXB
BRBgJwA4miEOa4vkNJXS4WVX/oQA22ysuy6b8BCmO95S5MLeVpeUPNkDx+DKdoRv
VGmliQcJPWn3cmYJaWDDlCI988NN/1Xw2VMtn8Q2aQJsLhpWxrXCAruqQFcrnRbG
DsHLw7uuc0QvXTKBiJT/FMsDuEW1Z3n95BBfzxHpr5EeIrsPPDzybdqSP5/dwFxn
4FEMdYchWlcN3hsI9upJ8G885LJSBn0Bdn1RI6s4b7JIHGLZL47PtahzMNRJmzZC
5dmbmS/qhWGD5khu9R0ad7x/mvXtBYVnCSJnaZ1gRBWRaqrG8/FrSfgQpNj321ih
9QJMJZP44g3wooMh3GHB6a1sX1+rPNPw+kjNljlnrzeZL9ekj/sAdB4mqQrAk80M
3A/3wgYyzNSubfJCkpb83KgOhBmr3q3LAP6ulr32TNMiEPJ7HyyxjKFYoWl5HfmI
eMF5C8nnjuenFpLGHbwNembVSxnozaPgMQPplHaWzUahlPQuQhidizzjH9PyL+uv
OeXNBXe5ONvHi3nb7n191LdfReoLgTSb42387wFowgvA1YCpxnBIRCSBK7GnHc7u
7qjWzIsiXzXOTUST9Tq4Pi932wwJ12hjLNBEHeCrT5xcayemnK7xVjS7DJRw6FAJ
OttQ8Jn1zTtWmxCvicmhHN39nWLQrABk0w+CrQI9jSGyEKefnO0V+xaP+qBBnPOD
xFBWzUWsXHx2YWDt3cTh++Aq5RiJcp0QLzBbyfWfJkUaaLfYAeDHnbjBs2EMoeGK
knUt7uDk1kUnNJtpvRonOY/HbLgpNwBejA7fQXuByLJQ2+rPAaKRFDpl1f1QSwFC
Lhe6BNWGNBZ6V8xxVrO2fWoUJk3dxgEBu++vJQNJwqOynrbbJZcd/bypo0dqhDdG
zggE+R5VysOqlrdrHYTgRGZDHs5hih4sBdr2wZZLA3EF77lDRxHGj0RiRpsfmhFK
DoVZUyiqGtykm3qwxAzI9pxiV4mi1Vq+rIaGt/+PaqEyuqtXZKg2dpogJTAdaLfR
nKf0OgIrMt52fFEt5HBQQ9c9gAUjl1VSAMu5NTRafrbMKPWr1QwFA8SiJvuizesJ
MEjKTdCoPLGLgY+FZ9FfE9gguxlLXeXtgYNLMv4kUEp3KNXxPKyiUVYC8hfzu+cI
V0SHNW6xhQwIFyGw4csNj2ce4lTzCvGIXs9WPuV3yxsxrHkMrIUxhOk01zxarTYS
4rY7t/RQhdZ5TXWcaN2qxPIDKpofni6vP/nqZentVhYnTWbHCTk6KQTlY15X5B31
TtoLC2m+pDMhfQEIRuNs1R8/n63R2iPqzftMif1AhqUdcAKpCKivRwbJvER0uiVm
ultjP9cm3HEfEjFO4fSSA191o2PZJXWYefhJE/TwITKUTuSGVXNOvrh9v40Qgrmd
mAFWPCF1LzztBH6lpDrQiHdZ4Isce/1ZNQSG2sO/Z6B//D8ZnFE6rhR3tnXtj5Dq
HjVbItmWzfUjdfT6Tk2c6pfzyn46me8dQHAfHtMwj2mDU+V52Ca7SotkGj1Vltm8
H/PwOl5/OZzs/KLk/OIEcmlLT248yKvPclZiBSUmV53lmTGGND6JOOcIIOv2cpQT
88H8jIeUCURoA9D04bpMC52RYw2htYhJePOXMzBszxrphNTsOAyerxkm9QUj3nNJ
BUTtKRgls3D3iMnc7KRl78tGz6yNVgoopqepgoPrwIlEQhUbki2AHfW8JHSwVqvg
lLHURRnH5SURHOGkxRwMNxsFuPLCG2kApT5uI5f03RNU58LgjUjdBecesMh06gqL
z79zLczV4Pla+qOnCT4HnLej6N0e1kEjuxmQPslBIvjbJwFxJwPUBDdlo5ZIX2Ex
0Y06Womn9XKHleo5Lw1PBMzUR5O4TntKBMjm+fmH0F+PVf3bsmFUaQuJhrLE6Ivx
e0Dw2hKaBOOVdhs9nN6aGzU+feRrnrRr1OoIvStx0L6/UvpCLY2XJMUnQijWAYKz
ECImwGx6En/ZcNMlyUqqjXDXTPLgES1MzOQ58pmQZTebiJho0BUruZmDcsX42Y8a
quL4fCudOnUu5M5fGX7rQI1jG9Gd8AHlmFa8sUYERr2/Mty/a1OMzELff6LZQpqC
uOn6lKLBPGizbr0QeziM17EPVoi1fvVdmarA92HHdZI0ZpdMxcOiogG0KQwo2AVE
R8tJBCa5QY2C55vkCoc4q9j/64azGQReGKXr+ZwHIy8So2vxhbHmE1T/J2js+6sv
nOnLddda7GdiLLI9wyYI0+V6suHAR+54hrqabgIBZTn0tE8d4/+uHhVnw10QUnkk
NQRbbomnwpfyZDtM7S21fQd2WTAbi1E2ZfZe39oURgywtuYzXjwPp3vAD0+U9Xci
Bv8+2kwW8/DmbBFy69Z4CuonXdhtnHaDrEAUDvbOWVzCUsFAUt1vXIrhP2Mh0S0E
movU3WAbeAxhRQThiqduiv7g6UIcqD9D5Gm7KhzwuEkWM8ckEXh1z0gYyiKWELAo
HT00NCkSqoQDdsvgsqabpuNUgFsMNq7dvhqkeEcybkoTc9T2FD5Ub7jtVNA36b3e
o8zURR6n76I+TwZLK+jj7+OUKOQ2i58K1I4cvZhwL3l7DSIPrIXBIc4XoiYwHfDX
6WsraFwvRxJ9G2g1yg0eRkDLxrtwxRR1BpKFn7sW9fcTB2UfqFPXfqZjTWsKcQWj
T+PooXSsLLzIO/qjfxNCy8ntPcQ17xHYIjPWqzBcmZjTGQYUZrc10vrvDArX5Qe6
8jY3FnfPeeN718lhBHPUgB41lh9zLBy2XNJRyelH0Pzpg/BMzVOLLto0hr+tT1Ef
XgW/+4nyPsOFXeVy/HPDIF5i2V7ZR/dyE7PoQJP2h00+tKyPKWSDU91dE7Lb7dcj
EB07MpFlFddZMo11c0DkyM5Nx1YTvNESsHeeCxvpSjqRHAI/1+ha6UH3fH0sVOlk
zG5ys4YsRpnQ+qa21fgOKPiEg8FNdlyPpJMK0a1X3wLFICZZK2ot5KjFEptNUu9B
qotdT+XiLLinpOQDL44Y1Puu53ejtuN8JkKrTQGr2DjT9NdG1PsxJhT7FsM1F0Nn
Epd23IdJxuxlFu94vV0DtzyNp0vzfV7bsOnKv+HCtUtfOQvhyTIx8F9x/32CC2gj
WlTQCKs0VIJdVf/6eL5EKfQWWlR+3tBbtlW9S6aKPIuW8JDXcBRmR+pc5EoIV+Yc
q6pDjtPCl8wJSnSfPjOlG1Uig9yOoPQDl+z/5N+2rb3ZsBsmcI16X4RyvrNya2cn
40aFKIRWH+j3S4MU2R1dQ22qIqaKIrS3h2qFKb6IRXW9ZjjGa+3eFAFfJQwUZ+0Z
yfAJgljEpt+PfzKhRNzOFebRjdEzF2reGAnsxud9fLWX2kxlmY1p/Ipx74HnECow
KMVUHtw4SokjUPVhb4l4eHM3EyLBIofy608QChvA6jZV+HZ6CzWpBH1qfMUtVTFf
njkCDel9pCBRkMNAgr8PeYxpxgvj8hu0aoarRv4/LcGQNabm3tth+xMrEjzrsvUv
WqEUghtAgwpF9yMz06GgeWXz/s4KxrZFOYvEpB7o9KRveZJNeUwKJaV5+RuEgx3X
/W436DhghoWdE6smaiDD0p3ImaEaOYinjnZt4EqcN4dq3MtZ+sUd32WgEnP68sO8
aCWHgTiVlgv+slrhNyHzQQVUSxfiJjdAntxpE09JkBWlFgRUQg/y0n4CUEpFqkG1
sUL4ku4rwu0bP1QAlPCEsv6XHKL5dSXXj+O4OKcCLvJfBzG3FWhMiAlgvi9ikK7Q
5NgqELZWgpHKgr2T7oPpETz/LaXtydP4f/H/Dzo/35LKn/E61lkE/IKObDcPS+fk
3OhjtL1qJPM8Xq7LVzonCJu4pEGRAYMGuDARviJ0ZoeaZUK6dQgGdr82RmSa6LuD
8mZSEyTcadrfp3p1EeWckbbYpByIS6uyEMRQdBVoaVmzW4Xd/8QLvZiLzeKu2Arp
Tr20eV1X6yZtBEeXzE3BIGYp5yEDTLly3mLnNxRZiQeR/RUoxvgQQTTJ9VyOhks4
wCq0NL2oXf+ozWx/+zHevmYDYjV2REE1fXMoljo8RwxCUSd6Kx/jxmjRRal7m8aQ
X/OsUCbIvLVjkuB3bcUqrK1G17Cxl1eNtTWmzYTxmKTKAIh3oKweNCQqvVIWqIAZ
++x8wZ2+c6Wr+BzboO3OR3U6j6DUx0te5Z9W1Lzl7W7ZqL1jEJyLx1hQeVOaMTH2
BNmhExyWWAbF1//zgfmOip88wdUfOYrcRrfAOrqwjTWjVvg70oQbMGjq40g0uwQ5
44lleghDuqNAUJ+qG75JxCrtOBywdCxizDfs7iBilUvnD4NqV4j9l6xFz4YOBISr
HS1jHr1OltOF7/CqrM8o6Glihx0SbLlygY6JiB66gySxGBdM5oF5jX6Mb2YOoLdR
fHFJkhrhKVrrluQMW3g3XKDa9G6KJxD9P2YOu5m9Rt8DG7yKe4ntXx1hFFl9OJT5
Gee6bPQvKl0R1OtrVFCnOu1r7ML8xnjVSQDI4+Q+u2l61LeELD/rE6Qvnvngxl1T
X2kNhJz23FCPYYiW6KzbzLSP469MSPPLgH/YKCxU8XrzEGsZI7QX1cLfgqYknAOa
Sn3Rbs2fNchp9c2hjb1sTDZJRwGz6lWf2hM7l9o0ZTUvFcI6rOAbx9LsI0cP4OQB
thm8iCklnvVb10xmjsviW5FzQxC+ZraJFkP6fhwAmZIcV3kmXYdTm95NYIXsN2WL
wSri4y/Ote5cDRwwrPcU6W5XTU8L9OO7gVqnIDeZfwyTJ26+6sRO5IblVxi/PjMm
cVwwwso4qapa+84i1G0tFcRZbOskMhJQ5RRd4kNzz1pLjpxecqI1VVlkKGeq/uiR
GwT8It3tgsuMkxAZOAZt/O8GR2EaAqAc+PV6l4kl1LJ2lPV8wrZOJYBEWZwT5hDx
v+dZe9d5TRxroVDrD5QRzpDkVn0kUHVpJGFyVbulmavq4fYs8QWYo04bVzj6exJc
UOblEniksLQ5OCKc2bDplupPI65j1g28/BPrBSBBtXNvcuWOs/xd2SFjPw5o5ZWe
a63xgcm7UOPrnWy0vMZ0mAikHN/YCklbIKkSiBPKKu9q9hIu+a621Mq8uwl6pry5
yBIvqn5eA+p363PygJTnkyjequV7RN/qV5GRYhPTRM9Pl3GLTeZl+NjXwf+fAl6+
qoGiSOIBiCVG22Re7d0EFhkPcaTbZ4ytMb0QUNjredckCI6sgcZuJPQxXbH5pe8m
T/OWh9wo9sTY8GKUqvGJkJMh06vKnehb7u41p8fyNmpLiKUPzcP+zI2gM5x5DuSE
2aDteBmog8NDGX2xqpnwsq+gpJEr0PQ0gD9IFtUpvX8fzCLtckDXCsyZTYAfsLwA
KxLipSz0/mUBVEaSF0mQG0A5YX8npuM3JmrOefdBaL9sZi1uIoKRZEKbe9+zjH8r
cKKSRNbtQepazSCUxdcjSZBLXf+lgwpKBby5amb3tssULPuqDhdqKj5H14ST8oP8
XxAB7J9P5RKZomYV6Cc4SYo8BAVV/eAtFfrbU554nAiLvvTSaKIQQFOxUGi5AvUz
m6jVJyJ2B4uXbdUCee8o2SxxJWmJesyXwKBHufdzvkaSmWVNSwH55VpFXgbA4qLY
vBVsgD6LYvYIN6+o5I568HxnBbxtEJCmf033vbV5vc21mQQeCWMjuawcnBz7nCa7
0Z1vaG6rMVvI80NzJtjgtw5EMGBBLeR0osgcsjDjv+Z9JtV5C/aO0WNHKCGaSWkD
sK7LF5Mas8fe/EnVhwTib2p8ZgYMaLrGxMH4grQFnGxStHYUR4g1kTx6AIHf6uyT
Khkq2BNA2n/2xNqL7bRhuJ3tVg/UdVO3DV3Eeg6JmKN99euFEvyaWmEeoVMCSSkq
a+fyPyXH86023HyfpIdvX6wIF7waNZOtS+Sw066aeACbts/BL+8JZ66pLRG8XwM3
lrwFMCwox47pAGyvS06MsYc5JIeCGqe/xVg9GU7zFTcwqtZJHOtG7qkP3UNcA88Z
aokdMPVUNrfVqRal5204gZ9ihK+l4xDyM/AbiZD8Q5rpMV62fW/lcuVQQVStE8Ez
Q0WgGFfmgeQ3JQj/DiscT7/XyEUSi0jEiqPUeZ+obMjKJ6q3O3CM8xXUBcM8QaLi
KOX//UVI7QzEBCJcIp9Ia7z8kM78Uop6CEDfxtSfJNNBOa5UcUI6crkl4OhYWCPI
Ktimz0uI4UdaGY0+5Pzvctm7eFrurzduAGMQLFTe6yX2yt8djZfNhmtD31NAR3aZ
Qeue+6zjvDWw7UqdteGuRLcejAgGLynTkWiHWsNCQl9q4WOuR0nmeJpWuBnjkP5f
y+V3u5XcepcJ/qzlAREc9hKPKmC8O7+PsxWvQnouma6qBb76IPVm2fHDzC0lIiXb
hk2v62FgN3VNgVnhrEaeU9m5PmXr4kyetUvjr65dyAvoPCepYLBBlBVKePOCPhPl
ca+GfZ9NuDC0mkP25twK++jI/M/e8q30Z/fppQAR4AxgMlbd6Wll4FfEavSOB4Ta
JXxXbPjmzXD6wM8N8BDqJX8I7JI/kjaWySD6giL4k/8OjtnlqtrMDgdl78ygpKwR
YySsQg8Yo0sYWl87ZuHwMrwgSZMNZbjFJv2SCV6t6mrfrNl8YU8QF7gKZPEFV6bt
bq97bRPpovP4GwyIQW838SunOXas/W0ii/zqwUdRT6uHJ+/P3bVEIabQh4+kjKKI
0NXrSXrCZfjNXvAffnDKiklAJcI5CbBo9COolbTlCDhdVrftdWnSWuzY2vUhyuRc
Pt5mfSs0OZwzk//hSMfWZZ9ZRH9I2ImzXZNAZBbzeH61jSZq8YygId6E7Ll86WCD
VuSMfrHWeWPlBrJGIdbRZ5O097YXcTUohvxkTLvAduIC6S0u25JwBHT6TLNmhXfy
8q+D9fsCmRNfE+LuB8SXfUa7IJGADnMf6Uq7vk2TfDiqas+Fl7eCZZ1ERorHMbnj
cQJ7dxqhZnYNsHG5gmHfEVgPosBk/yT3+Feg45mbgrufetkn/gLiMxTO7vgvUd3f
dL910FDSFTqUYgTD/lqA8btmp2XqTq75OYOLBKUvl780Nyjrt/Odx/TWdSEtsCSk
QpGqxifq2U0pkiqnU13D4wwh8Fh0gP4r5ywFktc0/58XStYE2/UokH8qq5cM7Uq5
wc86jDFnXVIf4ljeVw++J3oWL9crAMivmufFL5T5FPGQETzt3IFrINKJ9p9Zta0u
caz5eG+8EQdKsqCCm2ZSChvezL6TJHQyBBWZKr+6Q0quzq2hh5MzkolDvc+VAP3E
gd3ZgHokzvRZ4w/zuuSJdGYUBh13DGF0j7dKP+fDlcovKl3rz2/DYghmxfwYZLGc
BdYlFlDc9J4JfImZbIMIIy1QCV6O9fpCCd0DLQXmGV91b6PtJXhl5q6geH0/BbsI
bRJFDNV3jOpyROja7i3PLO0gKs945o+iOwFKwY2ILat9ZzC8FWJ7QyE/z0QkFqY/
WY1EV7v+g9/ThHg3arVnRAvec802ICah2/Dskm43+fDYvaUFDqKCFs3LGEZ9Zb9u
H0NLguJeuAjZmbOemf0bljzije/9q8eKNzwaiUJbhjLZ9/hqNlVisPMAjGkn94kl
Ya4tt8votIU4ssdCf313I4Vb0UVdT9JUH56MHbTyb11mqjSYcMAyr+oEY4MwhIQ/
hY3uvaa+PA97H3wyBtVOfRYj6v2KtMzc8f9GC0E82SkKiapvknoKVOHydTyk/1Xn
B91w/fszpZmsOnhYo9O3qppOpoL2H7HrAcW6lluY5H2aZBMLEBo27xyxDRStF2g+
9LjVoRbWPKaTdb2fugK1ngWxPFl0GQ8HKr3sluonK47ekc1ZcczQJHlIjBmKl3KM
ibiFnjBpID9F79kbjrimNUvYyRXNvP8Pttbi5bJrBcf0QB4iEJlVptRhfk71IK+s
F/IguP+sBYbyFiGFyfNm0RdTnFVeOkCi3Tz3MZfBbsHzdfBwiyANihnHem4QHEBe
Y1Rv0aXGaGo4NgFpivYcIP/y1Rizqp3pyL/t5k74rRflfRwEv0BDX4PaWTj1ylSt
2uuAqtB2wZtyNk+PlwCtx1kfGUAmWcoOeUtQ6EmBgbr5uqr6HE/uhRVElQj8FgsW
K3IlgboYPrcoagBqoZJg4B3HbqfPQUDx9Vb4TPXcj/RF58WtprCdVWyLDe1QhVLD
0VoVGfeVxvZ6AcB5HuU/gQUAJSEfO0G6pK0DHcrdC/x4hPmUqkN4jrjNcoGIDVQs
Bmb1qt7yU2CrClgS6pfEsrDvxjEt/ntC+XUljBJBCuNMLvZ0ZgXm5wYOnEqOxAl3
3FhR/qdYdDAV3vPBe5m80jm/vmhvYuXNNv9/beiwQxNYW1JwtaalYxwfRQjr06Xc
R3cbYdf14p7akbogqUKezfJ8/9fzO7IXlcZwd7+LuI0WVrBco97O0RxluTV8QSHa
t9LfazDXC4wev3y54BzvtnebyPAGCGEEEAbTtwFeqHyVraLYq6mPIAN1a3PXwliK
Vy1Zh6Os6OFHhlBv3mlTqs6+cYKe/KLye0up9Ei8RVQgTA1y60iTFfvtTodAL4Km
JSoFAujtscyivIEL4i6vPTmU6pUdhKJ9RkV0XTsV//jUy1nRmw3T537H2roBJlQI
LzNdk2hOQu+n7BQIBuu04rH63CUFBu7ctjRMu5I6xfouzwt+55kKDHaNZ8h1OqKp
I6vlwSjBu0ffcB/1Bre/kDpJZfxImLxmCu1GSBnk43Lof6WqFyvRTc6vgdRWxr9K
k44tGCydvrrzDRvVvnbdcvs2cQ9NiOk5KlubZ24eGc+uY28tec7dfaW6dmpf8+j9
r55Gl4T4pVh3/830gRMdU6BgdwDvHjAQitSOY2DvgOIPPjqWUY1k2tgHdgpEV4p/
Sjh1kfVTFEm4DGmLNy1kc+mAtvFmwhPU5JzxKG1M2Z+ltGSW20PWZPLPgPQqRC7M
OrnJ7TB278mhOQw6xGQ3GAh2ZhWmPsAhWf8oIAWUwo8ecLpBnLcLX3di8XvZ6jYv
Pdgd4e1Q5fhOHKMmlRIFl8v94PtU1Wg3UxNx7dSRYbufLjmxCOjqbZHVE7lT3yOs
17Io1Nn2U8UQwBtO7IoPEHmU0xVBB+zDStAlsEkxfXOpwjoH9xkE/mPK6LLC/vha
EUMfZIp0ptx2mdbJD/kilV4AzzJM0VsD0snORu3Fr5Xhqfc0x4hc79TWixd4GfbY
UZSAoyZ60+FAArcnkrjqH80zA6xypfexUuIdnX2FIDxmPPzOv48S+Y+19VCUgJ0f
nbnsFjzif3heMnxJ9YEq5hMH5A+xPNkrIjxK0ZX6ae65osfaMi2ooWdH6UYm0Y3P
4ToSmTMsaDWnDwEI45Javf36SKtUmiX7fAHTNTXf3pVqm0DVtW3tYcBKQWBGgPuP
OVRYglgKDNhblg9kIj9k0f+zEQ5gET9+6osLeY1l5120Z27la3XH6ppLczsdhk4g
FsyriehFvV1+JfcmKrMcCkL7SA8EMmU/Hpp3jqGHty5Z6LALvIJiwCPocGmCaowm
ykW+bg0yBsluM7jwlKOzbGsjbXRWKEmmugmmF1H6pAU5nIGCGdRUNZV1Ns9WY2Xh
FQXSLbtIRTIERV9CR1+QaSb3FuvdPEwhVjlufg9SepmKZPVCQQLsp/jOk+uVe6gV
I0F8jMjOpyZ7WfB5cKWaOpp97LpzakaGMw0A77iunJcf5154x1RYP4WuAUPeqL83
zvZhF0KxtU5FMO4bNDxvlx5krW9ZL7Y/cMzYjStG1DzOHPpGuAWsavm74HUecWfw
ljFKgPNKou3mZr65CVNikBpEwlV+p4WR4CSoEdMcSqFqDXiXMLt5DBM23P6H4Gom
4ozd4iytXTiphk384Ps7J+7IQaXYsDwCzJH7cG1fUL1gu4XMlqdV+zcTI5K63Rpc
I04OrtdvtWSW/AEWFEyqRyqpUDvdGQWMdizuLk99bCp65AeO/iT9CfpfGNeNzWU9
WZicspzpHekWtQ4WSxqsZWv0xPmWwLxMGHu9thMLA/8CJodn/qbYPVQ6VXpNPWLt
SjA3CvhBaL6f9ZzQKmUz3hZyNswQd4+rrg3xQajS7xwxB8p6nTEumswAD2fPfbN5
qsTFN/KN5s1Ii3Bm9JZV2P2cv9NmQOlwFniDpkIsqZONZ9Mp3Ow2iYSb4NZJBUUs
yralZ3PnemNJSTTSMYALPYsnjBseUOAJ5XwK8gVS2KlFSck5KYuPNP5hAT/KyS9n
5/LAuf852HWF5Ev5SMSWTSiWR15bR+wfzGHJXau2bWAdwMjdKP/RlTe2DwxHZrmE
7bGvIyCWyHAixrxBE2HNOwaS5CRluB+mVBIqxIdyMBlWUmKXokVsQGTrFfsmbDxX
OBQ0Sa2CdGX049P6tMrw3c3iM5X3wnyDSJgPFobz32SyMy/8yqVlKaDNvrb4mZ08
/qgg4HknlBuRed7K5fzZKvSxLYD7qvN23/+yVh8anEKZC0/KGYVcN6DicGx8drOL
Jd4zqa1asILgPqWBrywJj8VSpOa9h832H83uTlrbiBcfJMp0faEJEDeK/bMgydUu
Q+nHC0K2IRbPsWrYvG4w5qM73jaIkpmf5Z57RtmP0H7pwzMwKIUgvtlL8em0NH9o
5NKfb4OdIgzkOuYeKBEyA0FehJoFphu32FSgnmLXg2ontv1v+QS5B+7H9HtTObzm
cnIoqj12NEB7sDFngs+L9Hu+kwcpAoE1/DZ9qsbbqzMZMcSHArtTpRaGRzsgzb0d
C6icFgu+srIcO11RF6E/cj0PvjLP9wp8AViAZZB39drH2hS0eleCNRQzCCYQFZUS
7EUSYmZny8AAz0cBteCy12oO1daCCUb8+X6T1oA257aTKiFhLY4aIUcQ8qgafRLY
i7KuZ8ovU4uB5ttOmlzCYSi379LOaanl6PEz8oCBsa47wTYkCakJiNpFpbwHjuhF
5RQEVsL0t59FwuIy7+Id1c8OT94yon37y/VH87EmqkmbZqGxSNuf8uxMKkTeM02S
3Nx6CfRy3rzGi9D44qMmJbymrfwrAmSxGH2rnB4gHNmI6NPZpoLUs253zjcZLqq5
HPXk7740LAbTrZN8yG6MaNNQHAxQHHybe+KXBJIE+6OTiS4dv+smXtDLjwTSBeMD
tHDuYsoox2WFaIl/jaZO8y1HZ6mvlgwRiQBBEveXfqKuQLi3RpxBZyr6Xua1HQSm
kfPJZDczWAAoLWlDm+o7GyE+8M9kZnJtHLPoIWa81joO84yuCMi1ejPaZszTppdT
XKHFZ+MK3vKDsLaGAVFWCubnNTS2tbyPTKWxEP0rGEdF3qGRBbawk0xDkwx2oZJQ
poD5roNkOLjpdn/DJofwl4fFJ4rGgUcEOAsYGpG0Gsik/z4+aD9cVNGCvDBGQ+fy
yul1bzkEKyousjKh1h6H0xRz0Wq7r18qnFoJyk1UIUadafoeFkI7zDCYRLE0+YLY
v1uasebsSYEunyW/j6MKvirq2sxzcknaXYRRhaDGTPPTKHZTma5Xpwc1IiB5BWhp
j+g5vtRuPcRjDzdYHhUk1KWR3il21vorOtzhTj5aqS4Aq5enyuTuYiwKCAQyMIoi
+tzUMGU5b9P51xU7gLO83S98xd1A3DW6D7BjQ+JnrdD1It1aHu7c0IdCNQDcfcgE
3NF8R2HrvWJnvTP3IxjzIKr8axo0ZhmIApnaytNOxBrUD0lVrvRv50W8XVnxIw/C
P9gfTgmOoik7e4/Ja1HHljYiNqCRNA9XwC1YiYxp59mFJicHHebRMBo/qrUPSQHA
4hHoDSEVS0TD5SPgx71UeUPmx5FlyO6lIqllyEzJTM5nAAU7/+b2FpcJEfWp5uJZ
60Qpyk3ywNd0qYgKsVhMgESS9TZljPJOV5X/gVKS7Fi6YxUzc9Novhn3AcWqVaaj
j+Ot7Rp4L5m2o36QjvFcK19j24NQYoGJ9pbUaqoAAi5qHpjb8ew+uhuOlw9LmOYx
KDB+8motVe/5Pl6vpgIWj8zH32g+GFQJFVth6yLOQ1HUDjwnjpvhZJcYdM3Vj4ID
C2qrN2fRfvMVX4ADz6kulLZmt9Xf/qSw0hcjjgZyqU3Dwx2ehxh9ZW34AlYocq3+
ZDM56eoGnuFXivRurpOZMAXJdyZzATaaoQwO0TnuEBoQg+FRVAf6AJfw0LsREX3Q
Ak9Rq22NsIoiVpGhrop8nPOkviGANaSCTYRmdAFvVk5470GOyUv7JsKtVSQm3eVk
58D0ubvLesX4TwPK81SU60EZjMsSWexrevEbfja7M4bg2BY/o+b8lofo8ZXz90O7
Kbwm+z2gPndON8U/i1qFZ04UPbm1deFDnwM2sMqZB3kZfWMFu/lVt6ifx22aEw6J
ay5jsKxB7F2l0YPxg0Kuc/PjT9E1u329TxMwZMruQRyeGJywre6HF87CVV+SQ7n9
BkSO8InRemHJ2D0xMgzvdMR4gQVlwfR1+A3MJ1kWwg58/1wbDNfLrFDFHFVw8MIz
OVoZQ6cF+WJFkZv0ZCLk4zIZcSVAoDb8jlkf5ZVuY9rNo+Yk1ZX3BT3kbFeM6qXD
TIVtFvowY379tlXKpSJ/6bmNU3kEuytWGzMQaqgoP0puL0dn2UwLHWe7o3UP8aYw
FL5IFOesakMMC7HG13VnI7tRY9SS+NGs5Bt4jaaKCTU2kg2IaqwDi4KPHLA81Aaq
TNPw1dRjdoxMhz90iuId3R7okOyeFrmA08TIcVKm9jz4gqJkwEp6DWkmfH2o+zgP
YoTh1MSFYpBqFNY7lMLKRfDkN4FvUyZapkSTCGtsXldbw85wbIZzLQGPU26ZK/o5
9yp5DFz9WuzBKTRgK+Lpx6ExtkFjTf6dV/ogZiJKctqtP4etaLaMUYKLY+7WATGl
UxyFvBn9cEXWLg8UgblDNlLOwRWzaYOiv7vHwXs+JgFo/NJmqFVHO2AS6tQ88bzg
wYcXLasZcPEvxhqIyw0GSwLXvk4wHmvJP6414XRrXXuPftD7ARyGGZChypMXd1bw
eQRJJcweZnA8aKhXqInW0/z/zprpaSV0X7rkt3Kn1zJqVhOib3b3tVnMHOM2Mi79
LAPR2mnyHmu/fkep2s4d1fO0ZeUl/b2itlKLeONXrFu+ywfj0/NqdepS5TI3+2jU
1RdUN8R9DSPL/K4e7GL/spLwMTKwqCC/IdnzOT3ePKH3WfomIm4Ee6XBgJXmQEeM
ypqQAXxiqppEQLf+HG1tC6S/8xoTbn3+RyG6kBB7cmMKevv/hE2xSAKnuoC8Fxom
ZzFRevp3Zgq25T7UqRE8/6xVSsngfplZoEqcExVs5vK5Q3ojZrCsu364kUm6Sqr+
uu5UTaVYtboFpU7NOGTzSkfk/pNKaN8e55JovG6sBgARU/vDpIQppCsCbScUf70f
w9rPj/EJWm81yjBEY5KrPCP9TfK5sLN29Xl4TLbH0yRMz2EJsK64vOcPYLwyF5KK
slNHaf1ugsSaILDhhW+j+G3ffvmUjuZIC4pjpz2VNfiimqim5ylRP+v38qOSxBCs
fHt3FOSnr8DQmutGJSW7kbw4cMr7wRN/1ttivKZRbOQaVD6hCjHoPysoNZmkMpvM
ojAkBEvXeKnBgtdKZEEa4DcXgNMMwqs3fbXuvNKr81OeWSO14uVRXHdVKRq1WLfh
4fv6GSlQqWBtuXy7T5AfhvRayuvOFe5Qs4uRbst5IfSSsbjEv8c7O5btv0gKox3V
XUxL6yTNRCe4/XF6eEXhr6WxUkEK9nXYdXlwVK773fC6PU6mTU8Oy6hfop1EjIgc
XM9GW97kWp7EL76PwkOeT2roR6c/wxAcVJUNtjTNhd8FEXqbeBiX2fIvZgJwBuKK
3r8IW8uGdx1fOZGLfUR0BZOT2LEiFmJMEg9ls/oxkknT59MHOTUmOMXB9UEXF6oi
55vFqJMGbsEw7CJ84qarZo5L4/SETLQeId3cKNpJEUfFEq4s27kedO4bkQyvGl8K
Y2U8TGfpiux7pG/cDrUVZmeXDF5TXt1GV9gjEV8IQhVapbjnClaPr9cdbOeiM3ZC
h+GcV0eKYx3CGLZAdo8L9roSAZZQeE9yTldC5jmSKAVx7kbiIf2LYRVze2EA8cvT
2M+aTqMqiFw8ObX8Tl1h8JVcKfbfKXdtBNwhY3G1uhR2o5+uD7I+GZszXNT9QlWC
/B4ozyyBaMDlLt+8NHvYKz/WyN6tzXPg7spwIAJdLG8aS5sKfB0BSuN4wWpIyb8P
nWnlGBbUMSZN+bShQY+M7HEVQ5ZARhtpFQNA0qATg27/YmpDWF4mS9Ppdgg13vbf
F7y3ZmKHcZMG1vtmiV8DP0UxgT1Xcbdv+bVqwq57G4UF0S5Hk2lg5eQ4ZpiZjsal
OVSeFVFbDGS1yg6IZnM2FPzt/eiG49YoH/Wk5w14R5Gzdvy+SR7ZGNNFyxyN5rRD
g9didVwlDeD46qV/F2BQMTvIjMi+4rgX6Om81Ect0jXRu9xDHz42hNf/YtnlKQ2A
fKTgT0a9mhG5+KhFs3vHi4EGas0MT2UhR7d89a7XrlLiKOWkxCjN6LUqwZOY30jw
K+o7aLOp1jpB2xJdZfuNTDq2mpaNbxkfh6ysPJRZ8rXQEhU5faPSNKPMCGgttaWR
dA8vicOPq9YtPGUL3ExTfO+jE6D+wD0Vfm46ouDSfdMs68A5bAsVWcqBrT9H06hM
BRL8i4zdR6eLFp4Ah5rIJ3PQLOKHZporz24jAtqfBtrJYJDEq6+hT97Kyt1kyEpC
AQ5kqVbCXrOSXlWQr5qyvk5Q4JOrWXXwHngljk9FzbBs5Sax9ZHPkbZM8D/MN3YY
w71yrJxL8uKOv/wZv/RpTcvtXjOtiajmIXd1Cum5C/XK9Tg6b6Sag3VJeq5arXO9
1gBWXxLsc9S757Wlr7Q4Fn4qhHi6kX2SNl6W/ClssRR5TAkh0p2l+XRt03OtkRpY
sq+YW6QzBfUeQejgLXxCTX8TQi/uvFTv5KpP5nGSz1qmbtFs/XIW16+WusKAtPjV
4Y1SpexmHJWuNdB5c//gSMd1x995+cKwFFIr34nAg+WEqYInWDIJBQ5TkovCQUCa
UayQOR7JgzsfDeC0khfO5/Wrqv0BvImcQp/T72mDgKH95yUbMp6RzeWhgToG+gAQ
0mqSpGC6jzVcBQbF8CdkCiA+yem4hzB3MC+naFPFEQHkIUZ/sraAvrm5/KDYwrdZ
b600RSQAlXF1y+kjQk83iN9cf4NWvQL0KVzeFG40PQrKjRSPrhmmJ6eAkGhq1b4U
AK78pNX2onCesxArn+dvisMS6FMPemxF75ptLgyuK7RpclH700lRekGHpzx+iIeY
Sgq9MFAJa7h9kWVGJusdelhnXArWZHKr91WshgS/lmImWq8owvKOtOKHkeLSe6xb
I4OJ54SLqVPzQm+RV7qI9grlsDUgKjR6RyY0D/zbOFA0O1uMBUe8q7diIhjAUDxs
WeZJaUjIU4rYJw/myk7G8V9qSeZpSJs4etK94PfgzyMs2LOa+VqoZJVNGWQHevo8
2hhxjtDTdctA5BhGqdI0KCN8xtX0fE2z4XrSkINSrLE1PoTmIPXfJdL2U3LzY4Pc
RUpOzLbRLe/sk5v6hJ9eEQIxbE7pXXRuTGMz5oeaFRjbJQncSaz8OtQEqhM0ax8B
oWFElRaq9+OU/d7iIbdVA6KcvWun1nSFo+GhCa7zMbrbbiMQn2PIxtvciFXsK3Xq
UqPlEfiZqOPVWVXSbuCAIapVnX+hMANGG+2/Bf2dqyE15eV6NswOjH9hj7gXzzsF
ng78usmVXWCFgrgi8PM3EBxFGlS64Zhdvt97R7z5hn9UJ0AHR+3jtzMyL2XuN9Uu
MFJ/qvugRmZ9/k/CFfNFmPX/miaNDzD8U1PSUF4EnWx7Avo1OHE5EOSQfl1OCFxM
LhX0d5v/eJlQe5vw5DKLxPsI7YZNHgpK6g2C6rTZU4lDApME9b0OVT9JZuiQFOVa
RXXvPBW4GpZsDq94//4KsiD4M8tF827dYSAgvAdAcp/LV2Dxjz+JDAZ/aAdvsACq
VuBKeZoFfgX4/l2OU9ZxUgcITitzGOd80ysBDkzq4vbHoLwYSAB8alF3czVyIrxE
5I+Gu2AVmGs4sVv2zBb+IcQ4EMNyOHcTk9s6IKCPgvY4J5jBUWQkv6NOnwEXtp9b
4+gq1X+Nouf0nAg7c+mECLsiB86RRTm3C5F5YqwKE1x8IHCmg+8Oh7JDUlhGDjLj
QN99Nj8PfB9NyKxEoq+/bUa4Zqhye9WEh14Dpe/U00GFfO2EsgnzbCGQuYTgnG17
OPQ5WQ8vHhONE5vSYUnxWiS1SCkS5uTCsi8ddqAAoTMtOTAQ1AQr8bDdK/5agjSk
RhfSSDhiQjWchX36IwIf0gRkX90aLQnHXqqy0rqqz+g2emL3hvdUDn51veGTCWSw
8RhNQyNMjpwpRgeU4gXYXvkbLwnwBfp/L0qNTgE0yQVpOKcyArRu1xZ/6gM2AR/Z
PxA2QxL4v/hq8a3BchL4a2Xc57g1rLTKEPwQyUgeiamgF0wIwt9tKQcIoAl4uN4z
y7gZabtr8+MC57R1z8Bl9L7tYRpoW8fGRD9IufkKbTQrfDN0HQ237kvEjE5iU9Mz
B00hkSWUv/5AMfZomAe3xBMNibMPe2+34Q2Ma/PTdXFcgM6ycJdpbb8hId2Yo2hN
011QrcELS9+NmuEifZ9WJ7+X7AGqCRHSmslmSeTRvO1IqCUsn6DCn/LyUVl5GVoU
yr8cLWv4EozzQvkk/kieMKMcGzv4PA7+c5HwHmklx4aTMdk39CuDWXzVqez8r5st
4TlLHthWySB8nHCKC7LlVumhNoqh3yi3kHTD5z9aqkrUXiOUk0ZXWN7zquv+xBl2
nstSAIZQ7AdEEU2OTJtcQYi83iz93UJlBi0EE0PE7bFx6aoPmo1tOS/VrsTt9C+m
HKv18U1watWKEcqyE11mMsNX30/+PGrLck4UinzK0GmA1l0an5uYztY+Re8uTE5S
pW+UAHDrjQXrpSmyQzYEY6mhkyRCOq5a1ekDXRVDj63jvGuw7rTiMgv+9zbe9G0m
Iy/XQdiDC1JRJAQSpllEo1jPfz9NtDbYBkkYm9UBI3GAQNXqrIGwO6jk92q48Z7J
nMCHmB71NEoqgEu+WXhqUYTxkvNXaKwi9VocfpkTuxO08CTcVyKtAL0GCnllAWoH
QBNigky0qyceKUtkn2POuWRRru11PWiH072x/ounnNa8HRz5O7aOfNGVo1APBiva
eqaxpSR2PoCatU4p3YxG+2ma6cjDdLzg28E23E5S2BtpRwoGFcAPhO+u5rgYp82q
mU0Ueyq7Lv3knyw+Y9/r48fOfOyL2e8xUXPXClTeNyK8mlZQnBWLBYGV0/c69/Pm
JnJLm3AU8jFKhdUewubfTUljVAMAXmUYC6CytNH18jvRxJGJNuAK6dyR5ywuWCjD
6Q3WAUe9rxXLXe5vrqXeMeTU3wfdllaA2+4bskqsZ+U6fvV1e6FfzaOZXSJe02Qq
e4BzIF9lo3+WLTT7A19nKcrgNFJaR2quFLGB+zlOD6cumdP7/ECoZcC/1H+VO4d/
UK4iY5A4dF3O7YCD3rU8ZDrouSwpimoTAT2HMFRqCFUlgSXESNQeD6DiWNvBE6dH
zVRNy6L8XHB1VYh5jRM2wUcq5D/vlNF4N9D8IhSpQLY/sFcme3LbU6pZrJgrdXDk
Nznfp1fY4u28tHIDGMvqnMUa5Oo2wYz8pUvK38b/ennl63DfQF+ysFUrtLq/Xq/H
VBQkWI8qvIjbqB8bkfGZ3YzVX/SKtruq6Slv5hyeIT91cXYvkDXBhtbEyajWen5L
jJ/K9LUB/DB34VzT0k+s9dcyicJyCWBdVr713MLPAMB0OKzjcSiqF3XEM8UGzc56
qG3Qg+8TOrcX4yET9HEyqcLVokhtj0s2ztUP0g+l4EnGtDyxBkM3muN2pm26hoXb
JeRMXBHoUt638uUun9bMiwTMJRpiu4WTzzFrWEmClzjsXNPeDw3OmwWjAE+mRqHo
YXOq8MrxYWud9jtbEi0BC/bBeDnpa7a++OhWv/CEKgqXG07BTUlwAMrHO3OAMubf
nn/JL/l932l0hTmjNLCY5NHweyXMgF1c2OkmXcYuNLVyZADvBvlWzrWFpgoyYMjw
b/M/+twXgFI/w/aL9nQLUuIVXvDtMszCb7QbP3g4OhWXo93Z8cZgOz1V+EQ9lBre
g18eIG0+9sHPaKFxDpPJRk5TDV12l4mfvCPQsPPnX78nVZzL/nZMrX5XHmI0ydy2
4w/M7OUQ7sKxdI5CETaDnswi0REJoXjtgDKViJC6n0peDo4EUZ47qhbHCo5tt+dZ
MdfU/N/KLjNQzTqXrPExY7suKj/rQ1IRWoi43Km2dgy+0zJvja2mDGDFG702I30b
EgQhc7X2pVFkA7TQwNeECqLSDoMSFKDovmfZ/Zf+WDkHsWap1/fMp8Zy/pX0LNJS
xxF12MZnmWBKB0lLyFN02mluxiIpwbsxnOnOEjdmXE2j0FRiZ62h2zWUj7FKz0IQ
U62O8znyLeHkJMJKjqJkIx4PvdJnEhpMovRsr7C6gGoh/16Bnxu8oaEKzeTE8yYx
ZwRD36EHIrZrEaJzObW95AZj6VmgGw1eAEI1uT5QFFxmGxNa1hrjCmGI0lAK1bwF
/ZTyW/nErvUFPC1xcNN2SMqMlEKH5Fp5DpO2C1rR9sbmQv0UQoLzqYuKFqMwiM5G
MgXvKgaRdo1tgBwjTjjZQIhorTpn5Si2+OJNd3u8iFrL79CBM2QljRADjF0njC3h
PAA6IfOOCXKRxFjOo9W7IW6buCQHxSp8aOc6V3lKThLu+EDloKKwAbfZr8TK9lgl
3Nu1Uy+DitjI8mRueS8/cFfE2rgtmKqwa8NwoUkUiTlH8UQ1smeVSBnNbIqq4l2G
v5xcppmnnIF1UkjTDS43lI3Cudyh8257xuVK7GivWDYgipM0WyK309avbnXNBU9D
1Svb9kpmvEcvcxVqkH4RBi3cdxCZJgZOm6/t5eyuzYNSVb2TW8wjx/5vEvSfLIyt
0bg+fhV7OlLwCyDOF84XyyL4oerwgLYoDCthu0dv0IS8WLXlCaCSjzC3v4D6piLp
wMLIqr9TXFt+M440ykdfg5G6N5WlHRCkXSDP+Z47AFz0kdUnLsi+w/hgjbFbGz9o
O/7Al1Z7i6r0JLIyWIczW7ZQ8vO7u10pjmmMqIAEpLq22Up0rt3KFBRzjUkmogII
lxbWlVA7IgqJudbSkr8+y02dez/5Q4iVjBhhkkibbYViiILsHOoNNctmp8DMYNfU
iHt1SA85aBBkwejDAs/Ua9AaX6MNsiafrOhZEN9s1pImFPikS7lkZrje1F+m68Md
EytwxgbDJBNC02SD/u1//K5Hnm5lp6B55P0f5pezRsP7fpkygkZSgu6xuoVomxoC
r/7wZdC9GwooADZzvzsiHc63fHg2gAnI4UG4q/+cVb/7Z0PLV9fwoPavRBX6ZrB0
2SIhwz52Jjp4rk6rjkKuEuX0R1Wu18htZzsam5gbbTz2JaLQQEEbGfH6P6mnT3j7
cPQKZyRDo7DtHdPwHKNLPPDUP2u9M3kg2ztX5Uz3vWt3yzgahI1doLSyyLrq1lFw
wBHYUw8/0iR5P23wLdwXZLK6q6Fm7OqA4XJW+trTK3J38W3qIAHc5RiLjBQA54b1
6bcYFl67wfR6x6rrcq2Le9FZRa9mvfVar7fyROFPkVm9P5iWqL5yI4Hay+kna+6t
OTWUbeHkaahQqmWD3FAmt9RY13phyDictdzLoxssNYB4c3VaokyfZnpLuq3JwP4S
ZdVatwyInhK46fCbRdaGGxExh2DrfYFbj9E3j5beDr1xRDGC9Kz2HiPOEa1Lw9CC
ZyEGQcp/zzd02DkYM7SfCi+yGJzog59UnGb+T8Y8R2pY855qgIYmto9PLsvtAWfL
DljuKVRVlbs0IFeGIbmmS/BgY9596+YvHNwGd1UDzTZSlxr02wtCSfg8bE9NrCiV
bNNBSW+igbqsdvpkEv88oDJGo6J8DLD9F3BwsI7HXo8JmzatZLNTvHQj0kml84tM
LjsdNDzy5xQmeOe817g79Ktfht0JeVIiDbIergvPdbSvC/+SIFL0bzNC/A4/LZ7H
buEey0Y/dVLs63dyuTQDejXubSoxqwEJLXoKkiLgKjmt1ZT2aFXaZZIksfrwdJCL
JENrlJjngNoRJU1EVRcASGF+94XH/Tff9EC1RcUH5Ylq8hsqLPi+dUfVL7WmOClm
bNhgK40Dlly304z8svNFk0erdxUheYTqW23Ve+lMUeKTMhhg9zADPickFk2V0Plm
KSzbq8sUNWEbxduUGsig6tBHPPMIrWx6n4fE+ZLj5Rci6EKV90vnp/ym+ITEp0bJ
d/Iy6kv7WZUAklYjfiqIxHus5sLILSWh2KuDeX14yOKtPUC8bYIOlLjqmEiRzMYa
BBky7//jxKN7JzRO8XpYZmCKyKx90sRQ09sOt4S8sYRDjT+YJ5Xg/wol3yeGeyms
fMs/fhqo+epwKBNlVr57mPjuELaGm0oUxd7fPj23S+kRXLwvxe0hWG8vAiiEbDQq
BAFL0B1+Ooz3fmwrDLJkyB72ZgI9P2i41i9xzWt3lEmjzaOnvOgQGGS3P0dAQ5El
giC3vqO/iZUk4wJX7UO2okqNcQtsY5Kblwi15eSQv3eTjBjZj5oDe7tlIlyHotx+
1ozYlf9uLyEbwjIm05Cijb79dRKX1RmayDD34Ma/gyfJw0gjynOIdMqX6HaZGvFw
tt9hc3XARcKSMiGEFtZWARgZnYNfKFBKGAsME+L9FdKtL5SQQNF4FW1a0kb7uh4n
aOJC0oWoT3YQ/waHAZYB9x070tu7lVOuBx9IA37Bk+WywhoiAZZMDv7aSKNwqAE3
SrNY9Np8itwjAn7Vfh9sq8Gf7Leo4FPZjkQV1OysvWXZtaJo4WLB0Sbictlyx7Gq
gVfGdZUzNv2zu8hyKa4SNIKDQVl6wPMkteFJMBL+YqYB+MXMzrd5CWVjzBRHGykk
AOjBv3Is4HqHud6yGyXM8U2xOlklCOZAaT7Zj5q1TYpFbgbc1nR9p8/KawCCXgNF
HCKGvM78MV+S8/uSKKTGdl9tds2n5eVwiMefKOm4/HvIo99a6POldNpjdV7IGOK0
usveQjZNpAYj9yxd6sbBa9QwMGx0ZrHMGRZxyrCPCSnc+dp1dO2fCs6/akPcSe2V
PYim88wvP3laowVHcLyDTQZh/R+K1lxbp2f8yv66cCVtJAxGFMsoptSX+qkw/lcx
sNYvDcyOq/d4ELOCYJSXRsJJ7QKZyDLcFQGdcK5UoORu02L2wscQvXtbC735Akkm
Gtnsjrme4s9hzZiiSt1nfMGnXNYVuChGHmIP/4R9XcoBplKLjkSfl5wNCBs/zPFj
cHhTqQNu5sbvNzyx+KP459kz4hRHWP8HZc6EyWNRpzO2lcf+TygRpViOAcVsOQqw
SvGDmB2YrHYD/ahmNLnc82rvW0tJhP7HZva5PNG5Ml/Una94cVWQnpp+wRBOcGnB
80AvQ+p/Xk8hPU4ylac8ujJ+gDnz+RWHB21zaqKCOkdq8qW3kmiqCCyGgHtMx9wI
sh1m8b723qnVHdlzibz2x+Ve6i16FFL+KJ7UNn9VVboAj1cYfK+rspnF7ejF1IZU
B5H8xKiC/Pm32TWaTMOB+/i+FvYXmoEkjn669XLy1D7QhzI0oRnRRPEbDR7Fn12e
6TqLD5AcrGQxvufiyGj5YTXd3PXOx903b6fOsxzkMFPv/uIBnwuqYokISZ+CjNd3
lInUL+gj5IvzPShT5UL6I4TqqHwECFDaM+bs45ZAZXPZK/8JmK9W795ceONvTdOU
Bnm0fhE18rjgYXx+lC98JlmZs8lRl8OeAOqRoJbHD5qeacp7xN+wxrQCWqPbSOkl
BFpRRlE8qGpxeu6k6hd0lu4CUzLFNzDRlW7imR9QO8wRBDwKLPNCn2Jom1kgSWv8
+HyZz1DosFDC78Uw4yApbxaCXlRw3vc1N4GGoOy56spUcC9gkfw4PCudez+6fc7v
QYDhpS8f6ILchcwj46y/4/0MY1+v4vVfwn3J85tq8syYivULx5rEzrP1W8PY1Jfs
8C5btTNkMVhUewov18BLYH7BP2ABEXMpPxBLLit3yPyTiW1egiQvcKF//CCmiOIt
nmua6/jCmbZvMpAxzuSX4zpW464XAi2IgrYNnMVTPfcmmPwsvxxXOnEUK4CrOYc8
hqq6mG+p7fXL67LQjh7lh7LgBVcvrqhdAyZ1IKBbXLUdFCezhZhuV/e5EQ5qnFiE
6azAM2CXvfAx51Tz1yPOBrQbtAC9Z15vYeJIN9HfJS6AUCb+v0aM8sG1NfSpa7RA
tJscTVcE23nbWDAnxg3+ab8/tQB2XHHWVgYvczelJH4WMJHYe/kdBooBkb1BxtT4
o0341DbwTO+4/dJzsga5t0WTuMuUhUk4n+j+dtufwnWsMJ/nNZofCcC0TAkY1k0c
Z6yOsASj7VeNGRyW0r6R7bvvVT9RiUhQTbsdj/FBFUUSkw3LqvyQPC697WqzAyMC
Ol++/htIEoirBYFlZ3OeAhMcveIzDTtsgaOEFzW65WB2bsLMh1R0mIi8s44ve59K
5KxSJPxsTZGhldyhb16iVpqktA1ryM1Ir0ltpZeSszwSB2d5FXQV4ZLTSfHMG+IN
2C0TQkXvgfYkl3zjux6cqYtp9DVd3lOcYf8M8Po5sUgjPSGn+Q0QMK5ulZHKWyrA
QXCZGwtnGPd1xvrJ8EUgqqKZAhz9WBpv9G3xgsgI7hqTNr2Y+RR2FHPhU4jPc2ee
9Hr9FJtfCtBqJGV021WqxjHDAW8jp/URY8NrnmUCa/8eU/XQOo+K39RL+1XKIKSp
9Oczh1zpPv3PlK+P6x6gCugNZ1tXXePSehWj/G/VOmCMWhViwFhJrNCgbMBvDZtx
Kd6r3ZXGr9XSfV/zU+StKdvqcfIlLwzKhMxzzZp4//bqamaU61FPM8K4J/xyKgRz
Z4yDp84VNiZLjfDe4j9i1eFKaXuBtT2TzN22FyWxW9Y9yMTrKTlQK5J/mA4zcKE/
9R5ztMwQ53mrzmuZDPdhHTXFobPyuxjAr5pYgVDW9qzKzV5cbknhSwYn0Mpold9b
ukyTXZb+6sEGUCHczO/ZSyxt5b+gL9T7PZzQJ+7Nz/0VCNty4U/BMxobu9Nl5ODI
KQNc2Z/ofs0p2mfl9y0fa5+Av1WSwrmoDy5limudwUMgW9lGtjt+XptEXYZWhtAz
DhKcE6RALLdb6GY3f8VJEoDGjSqt7RWKWvesilhX3eZzoXG9wXFiT7K2hRRjOEl6
UiLnYdp/O90OcKmw0E4Acwh5ZCnCADAIS6/aGMFEY1MW9dw7KI4pCD3nIm8yeRmK
2z/cXfSxCl5jwS7oRs0eEEI7wzQYZR4gwaYfn6lt6Zh3s88Wk1u9rNtltq/TDrB+
6B0Cj1lB22rpme5pwHSuOYZF89bM5q/mYCAXkwtJI+7fFc6Ib1k8RnsFjhprmfJL
tgzwdCywTRUwuiuBmtxL2Fio+hrOI6ffgyArbD02gdW4HIgklLVH7pxv63jYm0eJ
blSBeUX5hVtVb7JHmB2aynQJS0Vb0cQngczankkpmEc0JGS25nZRrwBKNCgOB6oJ
2M1ch7qWsvXC0WoB+KBrtnpRCRGg6N7ssRq4xni1rECLXRdhzcF2LNpMPj4gOnOL
0qW9y8lnNQNuEaOxKEIjtTkMR8l3VpnOoVoHM0TfmtzceOSxK3aODJt8S4E7z49k
blH50EbCY0a4d8j66NEZgkaeSmoGzmQnmPEXn/SqACUjg2USc/b8OasRDJujPtZI
bXMev81WIyHkgJaPOdlQQDgTqh6w5i/JdT/hayymuJSBYC/a43jyoVTpMlKixOqM
nUt511mMFgkj4DD5/C7YfeECcTeL6/ojT12Kr346TwjSUHnt0/sidz86KO/YV3O3
mkNbvSuNC0wjPz4BDAgE1piU7g8R0d2Mu4Vbh11zhBOL5Av8EjpVIoPxVougDYTR
SG/QfQKmiiZ1FlTUeHpwuwFELzB+kl3UD6igXZMRnC3nqupCRy4dKR+m1D+g/qoK
/ErInBLKl3AMv2qn4mqg0spWSkhteXiBVMuTI9u2An9l5TBFYgDJTRjoq4H5t1eH
nQyodwdyCMZhH/2BS1eQLuaOwICUYpBkZPdWZR67xox2UyyrjxI0TJGrwfFUOl2v
aooHMwjbPZFsfIXNAB9amskxA2/mAD3A0UAmjY+mm+OR66MHdvvdWZVC8+QIcFXV
hBz/NQvJ7vuoIxPBEax5baODUa8PFG001kdsiFG80q/QAKEW+60U0+Om9ho/lt1r
t2A5RPs8J7MUeMB5gwISZ8Bcr84wof2IsHexpu+zqZu+ZMzE1Qm2VFQRBu7l30WF
xbg2fgesbf0ls+Kip/lEo3/zJVIbo5RWlRHwJfwsUGakekOpOFHvOCPQ9JV615vR
1Lyd3Ew1WHbytJLT4jEPM9JeNH5Goob46LgC8KlIDjHowMrdkm35QM9chGdQ7Unj
Zuiq/+pV5CVK+OX/rJxbeCArs6baLJYXHJZN3xyQtuuO0kvTWFlIGyJUDfICQFp2
544lM1gO1FX8n/VNgt246cdi1MZ7ILmcylxeboxUmGEMtpsiJQvPQaOA+r8u5LyE
g16mpEmOpGIHLQI0PETUGCtdmZz2VhtGlbGCkjL+GFrfLtivzhv7dsI4Y/KZgkTa
2mezPC7hFCJIUV8Vndt9V5hb4qmbXNDB03iCN6JtLtaipOIOcpFtZ7ptVPMCpJ5K
i6frZ3XBJD9h4xuf+P/nc0FaUEaVnjgs/vCqZHXB1YOK37jNeAdnxVMFkB3p7MrO
EULbNNmA1Pt1OYp37ajxOzub5pYCF7GYOhRRmdxlpa2U17NleGkeo6eoZ7cWTbAM
9naiIJqfUmYOxa0/XRFo2p3f7qJyPbLcJY+8+K9eB470t/rFTzq9vxpBg0IRs8Ud
CkPgUDF0XuT+FnwbgF4JrDLzrOj64kfndSsjEHH5vu/h2G+R9me+U7Y2Hgw4tb5y
Ia/YBWon7rxJkTHXz7jnjdosilCThTtMeeR6ZE447OY4uHxM2BWBjcFDNvA3pcKy
mPJDDPI6P2mRtwGIDeG0/DgDtpR+gZ4m1dsx+6PJoFpDtPBPGtKRk6FVdMpUlIPu
lNcKLVoB8MERQKPPFDQM9E+lliROXkdn4CnSlxVwXlHJwsKbjsLQZA++OZBvjjA4
SLX/Yho1lMWac97jNKPCAG4FO/fhGgNzDeUzGOof2s3/2ZHIrZ6ksmm9Et+iYr3w
TdxZqzuE4Gr2UriAGPzHwQTR0JvjBFf7IC3cfQbvnwq8Q/NElrx6pf4iUCg9ojsW
e8sT4LbHsDIqiRitK1DF8gyx/40vslN3MdTjD6UjLLzKlxvsgGYGH5MlzxvJslk3
wITUfDNCRoMFpxQF1eTtaJiqw35SKDX9YdUWuyTidw7Q3NqiI4ebOfIFBidwZX6f
Jxb1DuQGRBr4bFYjq2ivzKkRfkgCiB8QpMe6g1/9RRaoYCjTNc8QRSqF9Payrm57
qZurrcuAVjppMCT+xlXMgIZr5YlZ+npvjz4Uwn3ymr7tg5h+/C3aCI+GsmXPKj8x
r0tsCwlZQE4xGowsfyNmyb16UEW3IUmxO5XsvGXK7rBsyNL5e+Ki0p77lfUGBPzq
Db5tXWaG1v8xn8U5rnJrUMTnjTi6SZO/yLUpID7mt9/ULE2WzkfKX4iNyyuRuYEs
a1T4x8S9nJVxjydfYQhqzQLRK4yTojygw1/DUTOnEe0p+KcHaY6RPuQtWzFBq8Ur
YMrJXnzp3yGMFA5kXF6HQktW3+qAxHEyIFlLoP6uzNKXmNIaqSpmsy0tLIhx+gtb
a5BAdNieTZxlvQ+r+whFqhCo0JmpQwvtNDiU7QPDhu8NHw3Ui95j2IjiF8dtar5G
jI/YubGunX7p363NrGmuTiO2xQNrR0G+hqCy1hb5QOF7YNId/toqmkf3hLQhZs9p
Yn/HttuI+bffgbEP9dQlo8HfopvkEKiTo8FGiFtdyEOHk0CCnsKV0OcGgAnCTZMf
5aho3eMRcSIbb63kzTBv9aY31w8Os7HE67Eaa0Et/6iKTKk9YWY4yrkeTd4Vt5Dr
RN66i0ezrOSELIbfSNOuCY6iSPkv9SHsAtF5RUqBmdDYDpmVsF6YE1GfBRvn/cYQ
0fXdTs0Au4R+sVJTfv3MTXRINhL14bS06qAjrIKcFT+zTYs8k/MmDXAClBhvAILq
ESCCh+EWYIDbERjISfcBLmkYZjJEmRLw/axQbg/WTYKGX1wW60NKzoAXriyJZzyW
MLMsMeqS2wcpWbi3EGp37CZqWQF2S/bvYZCcpyU84eqSo6BZ3Rcu6hikuIQGGzFY
YyyilxDVsYa/+UB0fg7SS3Tlp9tto2edxka02HRAR7qdpm8upfRBLdI6Vs0FhXte
tb/UqLWGvHTlOCbcNucFQv7dSZnSqRsLA3ZMSHbfaXEpv3X33+zn5N9rlx8KYBtB
kOu/76lFtDRvJjP+41gljH0h2r4DTA5Ckf8LtGswsCTthXhltLV1u61nUCtTUwF8
HYXCaWvT5tpH3el0eaYIASx6FnSsiezrmY5mdmM56E92I9uzrCw6w0+Hx1+hLarc
/MBxcZHT0o+hcrtZNkft9AJlSzV37XCQSMsFHClVTrV1jl4bdFvSxT5dUPoYscDf
H8sRnpefTUHFywWp6j3W8M4PZx8eht1g7lyn/QOOgDomTxB9F2BCvWpz8eEp0iym
ruCStEez8a7uKyUGdfwpNRQ2ulm8H9TwfsX0O1m5IAaikDruJs4Z63lkU0zboWJn
mI0er4Z3KmNaB31CxAAMPVRYJuQxaYtjsEYRIVdHcRfLYBUq+aOdwcqBC5At0J/f
NCNIGGhJd4qLjJ9Ask9XxSgB7FyIi/Yxn637Wf8aaGBMtv+o8uf+orWFZoY0u3Sh
Zxa4sZy26Bp/7Jcj66O6pVXJTAfeHS2XVYLxS+nRWjiuUP3z9DLfmdECunfBkwPC
qioAj5kifJN8ikdPhbXvJ9j3/+/LxuCzNsPqh4NL8aa+YFfqqkjGfJPdJdg7lwu3
GqX07ItUvoqxj+M857b4KgXoLTP2MAgbJ3wzLHKPLcMrcRbxgi82UQeCAaxaSn2t
4emHJcuwVvhCpYrbhenGkQCCI1ZFLMKLDbWcdwhTclU7x+8whIETloVtz6+HF+Rx
WO2qVw/guKVp3yMtdA2AvaKjbSBuyaX+7fWHLKjB7t1hiVuV1SpvfBAqGsfLwsdB
uvRPniRh+dYv+lLLn0CgAFYrtiRoO5oRdSP2RqzCGoNtEiV7yPh3Ch49X3hg01/L
diujxhdNxF3nFWLKSQxNi7L69EEAyKBEUnMJQwkjfd5Tw64LbeGyDHFioQqA5l87
z7naDKgqBNh+MXF0Q5ONmq9F0aWZG4XUnLnZTXrlMnCh23GUQ5Hd9DQkdfeS8Ucz
rU27s47O28MQix7QxPn/Tuj+j77hVwxmspjOat1YEd6WQjtw9xI81aAcQ0o1WuiW
Skm+fzoCX6A+NxrMXr/4rAprWg365VWSFDn43rufzPxcPtS8b9uQbCjyrls/h4gk
gaGGpf2zNRrOXPdZV3UQzM5awcSX+YT9guggIv/2F5u7uoSXcAjabnCXZxt1h3Gk
fuohBaray8GbcgxiQBh97JOe84A/UJxFX13MhTLd1SKJ92GLwCGQIMwSs1olAS3m
WfqZ18nED03LOexskIpttX+wk5J1PJZh9oKrG+xhA/w7ZAEo1UvgKAENykOxm1SH
Ic2c3ZZkl4lMLV3n3TuTPuiO9ruyPblpnMvVEjh47ikVvc8oXW4TzQ1haDS74H7v
zbu6UyowceLzt+Zc23XWLvUB2m+XD6goRX8x19AUSv685h+wjoRejOFd6MKnZdId
xOMy8aBj7UO9zz8xjwYmE8eBWdFGRuyEoHYqmLbZLXBMONj+AI69NZ+Lh5cOzmb3
9SEU04f2C8iY4CSEAOMHq8RiV1yPRQGuXZgEoCrJ4UkhkNST92z5yrbDDntqBwjs
/AxvSavRoEdABV8SxVGHk5PG1H5gxJWmuwp0vfFZuth0Tw4dk3hQl5VZLoO2qg1s
3hB3aSR+qWCrM0IFgDljrq/wboM8TqNFRE5WhWbuJDyHvVqAc87SZxSovIagM6FG
6ehcSzAZu7PX33NSoFPs3eG8XgQKVJBqXiZdf40kvlIW5dvAHao0WbrA/fVGmp1r
8M7T7WmKRY9Zx70Lmsg7viq66mji2gtPyzRibCS7WLLawg5QBkrzcDJmr9EHEEjx
IgETb0jPQi4zF0oY3yG+3slCdlaRc4HMmh+fZlyVDtdCNdaNgsrUU4QlMKDdpV01
z6fFjT10EldxT3hVIaQiVSdJ9GCuf7QfaNJ9mufzwzKK1aBs7phuBhq2cdZZ9i4G
j5vYJXuXnetllfOOs2mqL1tA0GpyWYnAxv7b8geKWXydoXOmaHFTudkfQ0sTjQ6T
TDydS7bRXeTeaEqOASWl1q7ELVChcg3SxluMZnaHGqTUsgte0Sou8pNb/x/dpK5O
ENR0IHA73lGVdQfWsqgpfqNl96cQEGc+qoVdGdtsuwWJb7qLDp+/KtO6VS6TeOuO
QeYtVnHuyhXDAjziwFgSzua3HV0GXNq2tvSJ5fDYQhwEYyUY4wGDSR+BA9xqMZpb
J6OFVYhYYn6BER4IH0Yi/1/VNkAndALEi6A7acW7KynlIOWmtAhxAuy4WH/Os5y4
uNH9C/KWzgVy67sXY4i9bh5/HvwA+l/s1KxC4Myyz3V9/2Z5IbMgyNie5PwN0X7x
4Ot0WOM9jf0f2Z5F/KQZdFZy7rDhHfwlYP6j5l5xOtZHD0h28a+SXKklRs9u11eh
FP9Hs5O62lemSFAYFYoShGWgzXy+8WnLrtCJQcrxWuJFjSaobNq9vpJk7Md3DYzx
sSagp1SgauBY+M98Vv6ezZyywJQeO2H2tmHxwERLRx4unpGWTgEKb8fSKKp/cDgi
6JuUtRzZTrJvr+RnRtBrKeGGMAezHKV8355w4+WFd4rAFc6vednNOFYMqlEOyRx6
Pz55D8octLQh/r+wWehzlaz1fBVIMM6qLTGzJo+qg7afm6iENYjueDk/vMwtK5T+
KuZXWzQKCsGoKabkvujMZCHJTtQcqSlEkL1LgTNMAfVoBXoHPHrL+M4lC0ikfpir
zS4qt3i6+8TATtesNbp7oeT8oHq21jXBMyMx3BxZNdVvka+3WEtUGbVm2QFGwxJQ
vPwp1y/8ai9vyzQO9eyONZOf0Lh4JRU1agiSg29fLKVEUxs+wpOI9MJAtFO79SHe
Zp5f2L//EVfX0/Pf9vb2zKaSd3ofHAwm4jnp8TMUwZUqn5Hgt28kCC0cqSrHXR1a
jSR1Rz4yo5W+X1ciExmO50ygHNrvRVlJAFSFaB1YnQR44MZ+j2EA1DsJB1Yl+iqg
N6YfUYRq5Tbxvn/4nrpvnpZOAhwgYaU+prVVGgWgJUvjY6QN+X8Zg6ll8Jj2Sh4q
CaRKC4lV90J06vgKsW96BQ595YuAuadq83nW4AEstk2eO55kyNoREEBRsXVrInaf
i5WV7VOsr2B+7SbSvUY9mWCbFeDxsncYS6ywkA6cAMvTzx4MNcA2EPeSm+cDHFQH
KI3rU3Dd5xyMQfG90cdDb1naAgWXuRIJgIM1f216To3/KUMPoz+zdIdU3Iu6a0jJ
9SdVxRfpdO1ZiaolQE12O0QFU7RqqnSA1ZzDztXqACutvVNePMVrlRLiz3+8W+5T
PCcvXHI4dMg3Dv9wDiVeJmbxYD18JMrT/ze8lm0ua3mz9AOJ6DqgeKcSJnF0eh/L
/hgiMPa5vv5n0wAvvO/W7zTRog/7YcRlGVSHBtAdkXyoZlQJPb2Su2aDmR75PxS2
vRTDB4ZsI3KNAPM83+YV/BRQkLccEKnPnnwa+VhRE/da+fkCMkc/phRJw3x+le96
aiOwgLGzP72gv3gjcSfuChMFOfBCC37VkdoT+DcLPyS9peYPTquLG4HH1vVhPEcc
7bys1jk/cuCpQoa6QqlZImrmhDLLnXJz0bR7XpLa4FqW+CXnEgo1Xm215q0R7HLq
DyGXKrnGK9UcaVJdXi7JVITZ61fDLpyZ5OyAZueuZ2YWiw+WesVtZp56vgYwNZUn
bSaAdbE40yrOMHtiKPoLRMiJFkK4n8/WUOEFRtExw/OuwRoLWRpkWZdlc+R//UpI
VQ1Z+x87g9arroHW82aT1tfViNNfv0gTekOLHCF10JwOGiZUIbnKBfOciZJ0KXU+
u+LPM3BsHoK9aw3woIza5lgVp21wslXV6i/Tj7rhpt9E03uiPA0hGfO3NLO5ma98
J4g7JY/AcRhcR8g5HYK6cQryxb67iEtbudiM2Sq6B6SheeuC5/0+4vHvGcaotZV9
SvOotc/689m7caI+/1v+QFGj8y8NymcJnuVyhAnbtBTVQWFNbBsbu+uJA5nO5jGk
WAsr0wS0cDWQLw5aW37rpzBFVRz+JcQwzcRgDe+2GQhum3jd+cjkCU0ndu0GhgDs
yamO1f9dUs0QQeUUrCs0hHK4vcIincUm5b6B0VN1+31HvbpX6Rkj3J+ZItBHwkA/
UV+j2C1crS2zyVUKqbbnfezs2O1F664tq0dz5yHpM7rzcigaNx5nt+cbTVylC1YM
IA6QnVE7WRmAKW/WcF4eRnhs/ak3PODwEIc0Nicmd+SR4A62fQQ838/eCMi0OY+o
fKJrfcGSMy7dTkqu8gR/3ABpetyFX5wzCwNty0n+fqNN7p8er0+Cz300EILqpiZ7
VDUtZVReWJTG5Ou8N9jZ+sNvC7tFH7o6SN8AFdFoxLFZDKrwNWJgzlq48x1E1Mdm
PhUcBcA4qlQ5bp/L2uULUA02j3KVib4H79tOiKCo6OeKCAxSEQD92P6/BESUA3jA
SVbG6gSjMU4s9TFgNuWJuCUAleLZ3D2j+zRE5dVtr8qH6b6xaPx9/OcwPG8sK6Ca
B2pebkG2wEX85oXf0hwYp/NNJLnzs4VTjKhcJO52tnbDi9V2jMoFefwNR8JVeAuA
gEWkQj8xq3ovmCKWqyZuQyrAIs11MfFexWKGqbO2syINguC4tRXpmPweWBhDMwp+
hyT7Biy+sN+uYMn3rg2leSi09TJ6AUpvV08IJRY207X1ndfXyRfBGeytihBAjbi2
JBJG3lIV8UFXMWUntvEUCNevBhuKb0JGBP7z66nruF5zMci6YF/ejCLrkb1lOeDe
Q2K+vN1prcmif0lPpPdismDBE2kFxuRXaD5X+i8BPwinbh4l9DUAdH+t2qnWYkcL
aWezhO5szQGsuo7l9xCvNQddjOpIvZpVWloD6OHg6tELGmb3UcaB61qer6hJlCak
gGDfL3QtOfes+dhyqwqGAXNgea5zQKmPVP2tN7JrtXvnpNFs9FjSVHIfqo5iZdv/
lii9CN9zUUS4zPVesLQjjAVJ4BaKqHlG+orhRglShhErohCQUbsgx+5UKN9/5Drv
S3luvtrw2Lr1O6sK4DSnU6I72H66UBtwlE2rFhp8FZ1TPg4sAW3BPYzGPm98r5I/
nXOIL3Z2w7y9mOb9lsM8+6ETDdKGQ6IzpdWkDvfWQGLZvt3I3/PveraSWveCd4Ty
PZslucYX4sClTQrQJVVcKQyIDVp4O0AEx0s4Bf2x6icM12toWSv2/fWZFX+OoXpM
NuspIZXXAblWRpk78hj8RoEGPmpk33CD5i5Uo6UnbHsXrc843gj/o3yHsrPZtwco
IYot8m9b6EIXRQA3zkHRzAUOrD14PsyP4Y4jLrX35XMwzrBdGmsravy54RLCdSO/
QR6r4yAV5XEfcny2JF3GiGVaFqtCOaZPRc47B4oCNT9rKIIvDjIy7oGqmVIUVXLb
5tti7xWii5jwFLYjXBGL6SDtgpY98fGk9Iu/CdPL0fATsJ3z1odGO1Q0y8sn8YKh
0P+J8A//KLMbdlBHXs+m+2zEbbjDY7HsrQHw4YpbQ7X+bWAwuQNZ1200xWpSHMEN
nS9ijll75M0P+UH3JTidLcXpkkZKrCDdelDJtO4O7Tbj9lTRO6AcPb1+pKVoUwei
DfwkYLH1mj8XdKc0M0iXXRTiOtYzX02U0DZtsss4UnKrE/Cb4qk4mWtTf7u+n9wa
sJOj6aXkdhBT7AYKVPT8FTQzToStFXYk3bdc9D98QJcpYyykaqxeooaViVpv5TfZ
Pvc26OrjhAWy/ckINJsOBgMBqsiE2ESJ8HRFSzY0kYo1eVd0x9XM9laofI+r2xFZ
B+4eIv67Oz5OvC7rjBaxCgS7K/nBKZW9Gmd5wsbDcGUzW+jhpgdQ2xLQPRtG+8AK
apOXzgCBjryndaJxE5DXUg37DOyIaka+3UN7Y0PKNZjIdIjkpkDQvnhzG4yJYr51
k3KgpzaLFy6lBLQq18WFQT75Nac1bmp84yk2xEiigBySGsBZ6tl+uzmqg1fZkU4E
N5ArodtJcKUHgvV2UWsQGh2ZtpsmRexGzlm9EWZpjc0pEfsCObicbJYLXcssUdRy
/8SDxu8aiaaGN9tLDKLbSaWI6R/ay2Qo2iWVznOTXKTaQ8QA+JfYZ2lxt0zAJKHc
LFbdoP1RhqRcGm++O7upz5Hl6L9H1f/huUgiiH31wMVZMOlwHcj9kpHQm+vai1hv
QQgiHYsrBh1wLghwo7cxORLdUTBlin1rOZu3EK9Zi1hj2O3qi9zjhMSsLml/+uhh
0CJyehRkoc114cfDVeIEC6Y1B5NFcjZDTY4OX3u45chODvaXfz+W6As7+PimRsYt
PCF8gUke9v0fCp/4073DuA8tnI59gYvFDSPrH7gJrqr7j9SSfBw9HYSNm/rsb4WC
2QRJIsw8Vq2s2KoJgWp2hi0hWStcreKF0R2qXw3f5zSe+kPa/AXCKYi5YlG31tb1
SUxbx3SyuPuVeaWkmPRHdcSvskAA90i0Z7QKLsjGHruTHK3FVS4u1aFcgJH8PWMw
OyLi+cQxL1R04BmDxlSg39LVtgWXc0IpSotTN4CQ5tdKUK0ODM4B7/ZjIn9PNjGs
FYu565yOwzCPyLC6ABIfwZjW1FQFq4yy/4GL10dgkQqqw0MU7ovWE61ySZvfgQGS
SmwymYouSmPhJMtjh3mMLzbR0R8vgJ8L+268Pf6AWwphgcr8gNkC6bblB4Pj/ReI
P7sAQo6x97Y5vNo2CCp9UlvwQ3c6Jx+YeNyjAPuKSMI62Qpt8AUopzVT73+pgGun
zJ/bGTEVFxaDf3M7IhSP37nWlO7IMGrpKxeh/QsKTjyaQRPqp0bOvO9IZySEPsSH
qYchPNlNgIebpL5CuAX4MqiYgufEEUJJokxcL8azvR7J2zne/hc2ZlZ7dbDMHSst
Mgof0DfflePDbZPj0gxWJlUHnv3YF8VNUl/nugV6qkLqOoSf5pN+U0v7vZRwx77/
S3+1ehfmXsi30vzWEFdUUTS8pP2gC5DOLnEbGUdnXmF6aHuxKzUoecwpJGSpqSi+
D6FmqxYRUccbXhBhTqmiVidNnIeqCFBrjqrA3bsbx4A3X2LUd/41lCMYgpA0KpHI
rRTkRY++8JNK6Nj3yeab7C6O9PwWTouy+iuV5E2LAMx1fEQAznL7Ph5k2cMpYtdA
BKhpWTRtTPhJf1sSsu4MV8bvMB9Vg/jLE+KU+nm6Hpp+aXF1TYnIBEgDGSRIs9ZF
9KExj/8qKS7y5v6EFx0Nb5fSYsArL4YGBJmPItOsZNqD9LURtTaM0krZGvn+WCg4
EErEYpn/xcRumzcwmljSDzGpFzletbS/RKNlK2cG3uNzxUwvznm/ZKTCtb0GU8rw
YGygi+XYbkhqUkWrD8ZSMOSwSj6X6hUJJ2C6r8rog8Ig8AsCEz8mk/eQDbUVqe0d
DnhkeULazr1Sq9iEeqGl0AWcSzKnpGk84ZINSmiXx2Lm7EbTLaH4XTETvSS6xRFc
CYSzk2MnR9VypGDoP/HBWADqixFrTvm/pQp24DKCeaYCmIFtBTVEX3KzH90CwaZA
D3/sAe24JXjptvip7i2YLHgiRwHcniwhDYIH9c+ir6yRJDeiwWD3N8qD1lM/gOIc
kuuCaE2i4zrRFMQMXf0Br9EAGTHCVtZKa79oq7b/4SLi1ZbGJBRWDJxw6jg4KXOg
aE/h/7lBVKCBoYt2UN6WSlx6SckVFWkyPYJnosRlfq++tfbF4UmziL+N1HKHuxLb
c6tHg5uDM9Zhou4ihIH7qT1YGFpKERUx9bScmDLLN80RMcbTuCPvippPQ7Bj8Hyu
4egtZmVo31xjW5LuqCCordu327qKVSzCRARKfOReyIOGXwIYhpoETXT8YT1/WRZM
J/c3Cw9m3V3zaXbSpoA/uZEhWmaWibzE2O3lu8eMRzptq0MQ2zKjp5kq1XME1vS4
SiQZmctffVGUbOxlcyRYqBC0l3LdNOa/PFK2b4B36epXN6GuLv89vujrJr8HW4zs
v9Hxcq4+tfrDlsnD7GalT2Z/G+4Zb2ToAnqbyIQ92Zy9CN6firdkKXaHkD2WI2Lt
DWhzLcXOf3THYf7a2cZNuYQ2hiHnETu34U7cKd9hrHLAuVMs1CrPDKuVazFIUExB
RDgU5wDrD0NVyD5vm43viEtN3wYKOiA2g4Pf3Xefz7li0aTEugoC5R9yOqqIXzhG
PFZyNY6MYcFPacGPz1DmlOW3HyN+Uwj8jlvnBKmvxYDOciwAAO/dv4xdYbtuLHPL
aBjj4hAcQQfOcHRqeEy8GNsi5yJRhzeCrgSw+w5PaeVeTb+sT6zkJHZhcujXFjVV
TPR74/JmJM9TA4/4RVgRrECcmkyaon6T3oBx7G7xgJzcScHp7SMyHXabRfo50fDE
flbheCrbR5jodBF38CMZH5Q1gOVgTvFdaRYXI77UhT8rXnnfZU5HS7cMP9MPoGmU
3i+hDP4PG/tbqooTVvP4HSwMRVYjbWaWmHi+Fsuenw3DUsRgTA/Ol4A91bJ86Rf3
lfx7t236StwdQs4PHU9TTWwq9KtA8jhW6REdq4ly3kUgf3L6Waft31qWcK96rv9k
uQJtPL1mYLuyN+v7QEo4356KFbuhSurquk5wTzAnoJS6HBm1OSC7B0KR5ysi4utx
dkPhvyREFVfAVZrjUwSV80THgK5eX41O/C07JNlbuzR+fLryNU75ViTwmzuHb3jQ
+KC1QGTVVEvItUsmQQ+W2dujpueDgwwMjFoIUdenNAu8D6y4wHkNTCmGjbYqBUyy
91auTyd7pDTDcge8vVHcaU3wH/Jv3+jmD2pumAHkYyvoZ5k0YvEaRwK461XYdz6b
30D8bkA6ZB5LadjSMXulaA0twulCxNU7mtwWSlTQLxiN/NU0sG43DbpsZYjp+IiA
BYz0Bb8Dv78QrP6GEmxGzs1I6MoUOfZHGtJj7uAg9AeOhhpKksi3f/pX+dAhrIAW
8FGSAj+aZKEWJ/GuLsfzQJGtcAivft4w+PZZbQBvWKNB6q8Ohh1a7bRCiRh38oWw
F9LuMHnpgQFpwdTfvIc4wUetM/vxuRq5NZ+9LlM0iBl+2tTunWcdwVj7fc+wEf8r
dtECT4l3z7UWtzUt8hd1tn99HvH6Txnc5BGpTOhoBt1qWIIix3usjOeGeNb+uuE9
Q2JXtrbjQ17le8X+7Z5apamnYUJkAUC7XPA5jN24Crad+GVE4LS3GM51sR21iv4G
oWfNm30Wbqumqhky1xeQgMuI4p8IIQx+n/9uphzekteyzDsS7uLt1rZvyyctnde8
BWu4fJpWW+4sKDEsdU+chnZuzW6QMx4Hoxq2B00/6NzQ0HI7iDSmuyWx1PTmhy57
rwW6sPKBc9NMmeVGJZk6rrqtdIzTcXula+L1b3xg5Uj8qepzLLuITWE9WthHWlb0
lT0ujhBDLK7DHQqMc3FJPjwttze15S+O3LWP/8jhzElAnsevqCszqJarOA5mex/A
nPeRoBhKgYz21ZeZ7qUcv+xfNXjHTH7IhB7Z7jgLwoFXDOqu/5WZR/6B8YqxHkzq
8b2sPjvwrKLYmb4lqIwlyzO98zcexy+hnSAE6Y3+G8aw+/GL5Po/Ql3M1ZmAW1bZ
Cb1XdtPo4xAzXw6aQP/gJVSlw34FAZjQVYa9Fxp+MofqiPXsFuscIU6pvXPGLcRH
qypRXYSd+2FSvJVzSk+ubyIk142ENsKHghOTt0joQ7qKlkHsIEKkLX3s9g64XfZh
j0f2tSRtNBJjgTWyizB3dNulzycG6k8ftqUDsAWWviNGGi6yhsSZU5J531+SRG8P
LcY6oU1JH5D7USIJnBMcOOEZlyDPu5+VS0T85+XvChfEhnE/f2hx2Os9JgojA4xs
FFHtI6UPyEktHFcHi5lH3NHHi2H4ZkA/q6ud9DfSsmA/9U/aq7jaXsG/wzTZHB4p
YMK77T31+n5ycQTIvhVjf7ic6rk67k/sBwimKVluXhhE6W2b8jUzx2k+a3l4TtVx
ppA2fd44XErUosw5KyEFNBDonrzuWndArUP3iKd/YdUY2Y5+sTH+3DWPHDG3Pche
b0WUXV2Bb1rUn2Ahlsok0YPL52NCWK71G/NA5tcy73u7iVTyPjxHF1VpuVFvR1G1
nl82skD5LZ3hcHfSnTVapiyxmJF+zGV2etY6xFry68YU8mT8i5h/35LVGHaVQcgU
hjSd1KxQf3zPU00HWJhAqW/e3m4KUfKnJsa53NkLqKRugrfMn/1KnS8YlT366LyW
HcgtxG6lY45skmSuOcguP0yCG7WTFo3Yb1n/QF589ScCjBZoFbBx3J/ktvfeVbX2
P2L7gpQQCh6TIuQYyebmkCCqB4nXEvRtbp1+N3CbNFUzg0tK2Y25jqhFLDRhhy13
rqaC08aL/PUPGz3HizDd50TaE+J5/KaECCkpzE1nNle8nnhgwR5tJzGxg/N6LI8J
DZIDvT7iUmyPzuA5ZakabtD/Pjr3tGtWET9SAgEZE+YtiPp7lEAp6dC20KN24NBO
9lgVgDWBmCZqmV3T8qlkzBeAu515UUcJMaxswnxzklcxzFwZb64H0GrqR/06fH8K
nApAbv9ECA3/bm2ESwCrbHvPfivqLx24VJfQWp8jhbMuFVwNoTkTZMM5ZTxHIE9U
unKgqu3keCYz82mXXn3eks9gZ/kBW4qQ1OPxnzHdSGNKrUa0vHZIEw43roRYhslP
2bOVesqRF4QOtsyVHe4DPTsvXtFIAEGLAUUpcVE3PiPsqJr5mgNbq6PNiUP+FQj5
iSKMytMk3Igkh70Ycrf789ETBoIFhCJ5GCuTShbyWWXvTRwBSP2uVOUS5UVX6n4K
u4G2IX3jmMtTCzL6/7fRuMxEhfxVhdl3OEIFI5bM2IK/JpLDBijQZf8j12P75k94
7yIW2BjR8aV3eKDuBM7QGW+XP9ES2mBTqNroBgrePHkcH1R4Wxg73fjqFM6Ele6A
eWfqx3I52oaoJ6j7WPAPjN7YwqW+HDjDGKJBwAJnzZKdBwEYQUhpDfzMai+fy8ZT
OZJVjypy6v/3jasxt9EHt+hwFG+s2CfsnbDwgu6Lec05U2u63qIAancyus2CrD48
HSB+eZwMBH0jg1450hoKi+Q7q41Yswr7kR0Pgc5zcYNuYD25gtdRjaTmTwhAcJY5
N2AcHbc/kefmIeyxizu8zz20jkA+Ue6fGxoApjAXVkGWkRGZlAG+IUi1dYVW+iOb
enxP/XGbn9mzzHKRY4zGclpzBs/3CIP9/gfvWfSOGoXzlHwrcyKh12FiSR5Rft6b
Q94jQrg2nwRtnjwAdnVYfodIA+qZVEGUZ5qP+qVofydUhmZL1WySjfI8203xm7dg
oL+y9K+42PAU6vtN/fi0MkgAFTC3KwDmQ4yikMrXNTEEuxbTo7dXxyck6Ngh1fsu
X8H9YzieKDDX0v45LZTRQA6Lm3LZ3pB7fmZ4ok4iOcKE6Xgq0nwcL51eGFTqgxKl
yG19ecSHE+TNbDQnFC5lgFUixeAuQMqlpBTSkZmyNRTWo9Z0tAL/V4akVAS0sE15
vLlKML1HXj5VNSSjxUi32DIBbKfs5RiYZE7YJgtXGg9p8kNyts0CU3alSQ73dVmo
F3PbbtlJnanV/rvnD7x8MPVE4p1BeNr3shk3NG9VGVytYt0vJ8NfTROyaUyVFmUz
dmudhMA/d02yfS3cu79pZlKMyRjcfY4J9Bbx8iCc7eh2tRF3EM0zWnK4ruTk2zk/
jn/WctEoQL/SKr4CLjbM4mxhkucbDwXTtREb2PtBgS7FntVCw97b/MoREJeTXta8
XUitkcfeUU5BTjdiNiTrzXQ4fZ0FujxZN3a+EfvQCMh+mYQWAF5xyrvosA+VdX1h
RqvBatvmIW3izOKe72r2zys+XegTIEjaIIsnZ521BkHLNieXg6zrcyZpIq4Q1KXG
ZDio3ub37Fd46f+ZzJUmbWhs9z8MYFmk15a8RxMEC6TgCInjJ70ofFdqdlhJrbgd
HLYAD6exEldkM5IbRUax5V1BtNXSkUj2RMv+t3toeKLKMWwF5wlshs03Dm7/bmRD
xEJ9L4mifZdatB97VKXHj/BQ55x3LzW7QwSY3ZeXFVjQRfKmAObHg3/WPdQJbXe1
YIKm4cyEymmZnLYJVxflJEh3VCJxaEXbtPTpD5sv6YjZJgtWiURerewV4NPLcElB
WhUB5GgNoW2kAvTQVaCMdwuRWNfw710rnxH3a6jNJ+wUGUesfpBbBiIU39dOclXl
8aMEu8rO1aF7XGoBfeTz8MiCTx/w4QXqXZOe/KK+7TRTkP7gyhBFI87MCtykML8F
3aRTvynhrWkuI3h4Z+iH8USbZdq1mBgJ/S1qUOLEAsjMeUEII9uUA8ppVxiyQjzS
qdC3eeunbRPHncqSjKcGiMa0MD15YYNUFz4BnsiYgtz4kxG/OaSpqvAYLsJIVkUW
wI4PtQ9q7a6Qlg441FSYDRra4yYNRWsd+nNVJD95Vp4UcZeUMXJIbtOtcIvMhlGK
II4XuZm7KPzrn9lsWEtstUevY/QdUoN0wM7nbYKne2lwa8pDf2uFsPCcNDSl4o13
QUMtAOTCcuGdz79df08is8+JfS58UKsMEIGJWiyVuv259r1H6FcbQLQ1X4tuG9so
6ldai99ixFq3tLbJPEs116377OLp8hIUl70PE0N8WKUTRWjOc5e7OF+Wzx2yLWvx
agaW7nqzE4oRiVEuNpptcZ0BtVPwtcbPMhZcWSMgTlFAYnc/he55bPIK6O8Sn0ye
h80zRyWYnAruXGbIXIHgpLSesSejdLfafQ4MbwMxhObwd+Pgt1TkykhSqEiKGk3g
PuD5nzOu5krKG5MMpmwvX/ZeYttFN69cWLvxakcoHJUoi2dvI7KEGRQ2SqhXV1Ca
W21DOMMxs5ChllxvgU3HbVt+v3qit/Anu8qxM534Ere7MDNNvebSpgUepZeLSp9S
jjoJdixw77NOkQeRzNFaLCfpNseNta7dhG9ykh0ALmJ6qn+xBiHL8jvOyzgnlevB
nbGT4wliPhwp8FmFU1rOmtO222oZiXBtLqc8jbno+x/WG2NuY/MGDvxH6iOlevG4
rka+FGLEFdxyC6UtvQ4PVkqKJu4K1HrepQxM5D7AQn8dLI6bgTzx6oTE7aj+YArw
1unSC/CqSIv1ubCN+mglmoEmawugUu8rJ7+tK5JFszRnedPT6kFcZgQjuAkFym6t
3+4w5nyI3/UVdRlr4b801HamrOY6s8ETUUu+qTDsTbhnWs7n+u3EnR27zcNI/xC2
9QgZw2RjZ/BOiREkiUzjPHzBB9alry6ZXjZYfliU+EZ4QwqaJ6aBj9IUE6CMxDRj
L9JNhaBea5aMfXS+NDh2sPM1TbcimFuoGR/okqQDQFrNOIkjtdDtoo/0X9pDNlzV
gHKjZAkx0JOJhUKdYiQD1hOgubBrFQDag4J4fbqINw9RJ7hjBNml5eVvrfpJuP6G
rtTjFTGi4VMCvVaH5DnENFuNHfLK9aV5k/K0W/h6H5F3xBKz5orPDtI0axy9QUsJ
e63nKGgrn0RLk3oYaRrgR9UcqZ9Yshy8xjA1CXRH7/RG8bNtGVQ2ZIVDHryB92op
x9rJB5rIUvKcA4bzkmy/7HAZZ6A7prV2nGXHyiKKbrk7hjbMOH2o3bfWKfqrP8+0
07g+R2k6eWTlIlhBDVtnFOQ4CPVKCuhHvIl8EvBYCE97tq9ObvVoh1+JsLq6Mjag
KL0n6h6sPLgtXchNM3vxri7xTABC8xbCwTR3vegKmWCoH9cvBavA3lX5Q2niKkQ+
cwLSeRpe90xItXwbliVVwkzXmqY4dfpky2BpO4mEsELO7TfXsZCKupFnuWMUTTx5
lMVDrMzrSqnt/cTgz1nH/5yqM+U33oK1kn2wFSkR3/YG/kQF54t6hDDf35ZaGG+8
ZRpuS1v8mYRYD2M4szTBonXFfTaDIj+mD8YYeT8ay374vebEUWadUMJpSiNnE6mh
Voq5OIWa6t/cFEr927GPsmZowydorEaML4bTmOF6R1Y5OHLdpG0USFv6+yIqmTDj
9p5EhRqo/GXE1wrfbazpqlpaXaq/kCPGeYhn5cO31a0LkRi7vEt9sB/9bYsPMt7z
pUBGkWsdfnJ6LZkWBpER8dhDmSdMBQTtJ2bmjzc2m9qOno/xeWK4LRhQb0VK4JGd
jjiuFZstjNvHH6zET3GenH3rXOj37nie2pOV/vSFaKvpDESmt4OURILnv65PdJ3v
nKGl/xQS/yNZESo5dFUoFZRWNlBKsFvhqVghS0C770mX8w+HyU8DQ19SC6xAvgda
QGNJFnrMqopyTVRNasNgJdDBAhiraqXoJZBA03Th+QNPIH0Oe3hwhGKnT5iEgsQU
ufifO2O3BsLpJEpN9zwIPcRCf4kaduRWjjHx6eFTB5+JkIKWX2B8u+TT2c3TQgdh
WoTGNo0tiFnhXh+ypt5aKuvbEre6MY/q9Cydd9prn/+r640wt2ZLH96E0GJ8SnDs
qb870fAF+8Mra5YNUSczdVum6wxK3BHy98zfyyAdbvbqTviUU80UKQaizL4V298q
lOz1YTKjm4Myc2QD/RfMAiEcUtmudT1ArRG5gyoaXpWlJRAqcSgYMFMpTCH6LnLV
wZTjEqHRxUzJt0Eod/SKJ1KzHEVKiNshF5t0hYA7Ai4wPJHVmFxNk2vqV5HWwlgH
NLDgRw7FLS2+QZk3ssBmllC8fvGzGCNSaeL8U+jCP7G4+st5/BCw5LuojuaXNTqO
Vodkowk3svgKXmx5Cy/Z4rQGl6ShUtc79DxsjCQS9y66dM6OiArgfrNwqsLbsmoM
eKvOyt4rwt3USXKB2ZhbEKL8V/ASBL//S07FN03OGtYanDtdi/C6lVUW5gs5rfuv
9jq7jfL3EsSFR8MajLgxaQqrkSyUw++HJLUYqz+41L1d73M2QuPiR/dypVchnP3D
TLZAre/NcgQw+fEEfsYP/ObKHnSz5XqKTjP3FyW0irhsixavVImofKy9SKTN550z
K/AFw4mV0OmhmjaPPVlMZMnF2SxQuzypnwNacP2g66DHTSMxz2Rs/HK/dHRB4Zo2
TmR6dFyQ6NwPSx2ANtzvWlal3SF5FCHj2+5hFy+ZGXLov0h70PYeldUGe+q3Jbxt
VWfYfJqY+xMBv/58nvS1XPf2G0CorHYOrJAZi8Qb67ME8S8W/gyK1X++2O1EDpkH
UEYNGR6Tb+1mScGb11cSYZsvzhQMvvDT3rzUwHKFKLnBfq5TXGtxUSk+6oPMhMaI
ap56o5sUL3ILpIK4uhLzdxQ2vf+3QIlwdr9X6ptibx8K8TRAUbzsshT+thkbiYWe
qmXNAjyHaphGNVtVYBqZPe5vFWldtVcLFZ8sJEL3i7o8NTSy9egttqc6B/MjtsqW
8WTTkCDlz55al/zDzAXAZ1EAvzHDe/xm1nlC2ernpgKeqz+mvfkRwcMv8P7OuRYP
mBE9npYlbLcVNIpdBEIxCJN/uwh0PdCL+mI7RID1g81tvsrBYShlzAHeIyIrurzT
C52IX+MF8RaaDEEwYG227TQIzuaN3Ga7XRxon+COckFW24JIu6bqRnGlJLFYL+VS
gBrxoPZGWbfyaB/wW2GvoYfPo9gO3c18juVnTt3yLHeL515Y9ZZ5I3piPisVfhyP
0sLFftAPoJVDm0lLzHI+EasaqhCPHq/2MVYKqnL53BSEp5axSXKBthJGiTzL08SO
EMTBGLVlJETfV6k5g5ijgXPuidx061hacC6LVdbp6yxHfFIoyg3W/mNh5cMvgeCv
Fk+8SB1WAAlEKNHP2FOZSu2Z/z3QT31X5VtFdFLJvByMQ49ifmvZCbpMeuqKekfG
/AOWFLtlkHuMBgBzy7Htrr9wDzhgNqOkh0ga9iEYm77a80kMcrWcX/VPoBtIp6Zp
B5q2XZjCuu/RE8SslwBj22msc4G6kEdT9z4f+KwJROdEUr42wWVwv/EpkmRFnqq4
e0mKUbukD92CJC8msyN+RiLl0hfqs1+q/6z3ZHE1KsEOfP0psIy6p/ade0pFywdo
JEr77qUhpMhq/3HabPH0030UMzxQv15WFEiMrfl6ZLroIgVDdrTrtBeOcKiLMAdR
c0In2hFwioJ1NXz6LRwKpmfZ4b9apPERDGzMJnANoJ6bJKJ+8cUImdvQXrh0/OHp
NK53IaPDRt99NfeVWc2Fjp4+Wt5l13VawuMigLB5VHPmdGlyYGUbUg8JMGUqV6Od
GhuypgMLJDS+/rqpCiZrEUbZy3T35nt9dN8Dp9elUB0nXmdqZJQqdY5x0LhKHJUR
gryaEpRDnRmR0+1ImjH8yWZT6tW5C6xKi0n8Wsp6777qBMpDVLldCI6s3/c6kiUw
Zn4bnkTaETkLg8JRoWCUPm5a+hL/jZN6kVzJHXXYdvAwFpBOw76P8K0DDBxtOb1A
MtZxxaNETpaN9MTkLQ2Yuw70YAZjIYvGeLe/xZCMbQ0aZKS1pJg6GYCpgwU8+Wdm
gzz3ybjC2jzjMPLASEfkdwE3j/ihp1V++0XiAI2yT762dOuObuCLYMN8HftXHSPS
fqX1K6zXLoGRkrTNw+RcjQv1y62MULLGsiDY1pTmRruNzpH6zxaVCnzvaj6zOexb
Y1CDgWlbyvCbnsAVP7HH7mAMWe8TiEeABR/4Stz4N5BxzV3+eD48wDzNoOuK1iFQ
j1z9LfQk+ufBvAEuJ2kIBQ6aA/y1ZUoo7XmlWiJywC9cdDSWKz1GqZ6aZaQmY+SI
IbhHtL+tPzJvaS52i7XpXXLPxXOT2f1Id7zVtySnCjZPIVLbpZpynlLK0ylDfEy9
HhOx/pmCmhggLMxRTXEiL52NwgWBWODQt8bodpe3KpMgl85aSNaW/zkAXAPbzxC+
VkmFchX4gb7zm6II1F/3oH5Idj91Gz32Q940Cz7vR/4VnDkGJdjXrOdxsnGywl/r
80Y4UCIKhjE2ErxDS9ky70VrsqveEfjXAnSYk7KYuFhMVkDPqkK0dtd64+hIss3e
ALGLHpIbr41i2VPGKY6lmr7Rhmdyhhqw3/nQ2KIqLU6ttYoaGWM8a3BjZH7RlcjB
eA7yz/lTNu8k1qOWTT+d5iU7YUEOZtIMRyybI2LVgN6iJvEs6zrEWlo9sxk0i+RE
rwBfDXwPaKJKQVqfPzJAL/uI+zTTSn4t6cHdu9/CmS80YPvemnINgFKQULiQvD+Z
Oy0pt1l2qi1bolfYrlIucMcxhzfR6RqJpZsO6AwJMu8LR9ReQKAIJbfW3Ei87Q9H
whPeo/ov0HtaLbHl/aFjQr17OYW4wUcCrIna2wZ7NToArIZTq1X9/qUDTr1E6IrX
eEFxIshj+A7twgAGNHxDi4MJlw5sJq2yJ65tYnCEzUssRewFt5xtlA61rfnVnaFf
qYQc7uLTWXbV+i8d6elDdvIdASvEAuTZDGWbz2IAAk9HA0CtG6LB96WvpaOcRmYH
zZI0Fs6aCdwxxWh5/nbVa2MAWcZu04D3uHPyU6/PS+G1NNvZ6/Ix6EVxSbtnpQgw
GghCAieudI4hNcCs6rkU78EdGOm0wabfRlyYE1SGpxgvXl++fgybWsCMIUP1qYWB
RFu2124vBAlCb/wilMdT0Ia3C2Oo5d7+bstw+blEzdCH+jxgjRg9CdWbN97FCSc6
8oGRBq2cMI+F2mWN7Ssge71dJnLm12k3JWEg1O4mMrS2h/H0HbZdSyE5TZrjMWV3
JXEm6ztpFezsaFq50whaYqLvi/kg31UNKVz7N8qVcMxQd2qbpMYPaBRUDYIn3NLK
cXx+YIb+2MKHZYDHqZ68cI6bDjO4fv02PgfQGUvFOHRXMnQIhrCaQKDe1w9dpvpT
/mbTuZiD5gtPLOS4YPyksLi0G2/08OZA1ArVb3UL9shHoy4pSx2q3sWPYPrQl43V
WJ4818YY3FZvKEam55JnqSTJilCq2zQxBmFMuD/4yeNItYDrfwU7xxUJoq7BY4cW
NIXoUGA4pS6CzPSqzDEEIRqeK3GqhcY+US+ezm7mNI8oqRG1/gCgKOnIiLwprIHn
JZaIBjb9+kX8pyabDkdPLUlKhyfJIq7hbOyCMfAHJuaNq5T9k6BHIRfr4Dah4Pev
TerLzofT84UQ7a9UQQonNaJ+dYxghSY2Qk6KYtS6JUsADQNRvT76yCJXGE7d2Eyp
z0lFKegpG5cz03uqPPDz/ld71DYeKJKrK+2cfjVESQI+yQlVxdmGoh655wzkPK47
meRBa7H1bw/ZSw6x+qkYGXS2lzDHm3PGRfvvSwBzPMgwz+rCSgTfXXGxFrBRzS+j
2RaIp5wCRaV6wlOq1JyRfbkTFNYrwpJwI18XztmoWVjrKojK+v6tbUhtt9dZYejy
iEgpRZb2ROAbOB1MeQwVuDrH7fnJCt53h1ApeTk3MFhj3GDyatL2KgASovUuGeHk
2Y54ppgwpYAJW8/RlFZQwZpw5EDK/cSic+KuVXhD7JncXaKZl/ZJrvepU9SDU/CO
FJGkmuCmSQtG681gGA88af4lnmHa3/0nEskUPnSuWIRnOR6Z60RHijjMTVknquI+
H1u1Be33qNWNtxL5e7EW2PhRCcR85Nsbyj3goUWPR9u0iKK9ibRPwpTeXWgpf9lB
gRaHbffAoqiTfXzfje9CQYwrYj6zRq9UakO+ic1ZQCm2LaXJSgXbQBq5onG0lMYI
41JFmd1wWmBLbNOwzzu31+KZcSOGpmmVMNVhP59QPBMa5fuyN3U3veh8Z2mdb2k6
1rx3jqrzXu94pCCSQ0mx4YVDrr1utcle995Tb5CXRumIeABkMjCtAGnrXr/ZbrOX
Od4AEOZYbN7Vze5EJtmp9VJ5y6pADrMelP8QHUXl0ksx8Mt7TEjDP9UFf+QO++Xo
k9xY0U1jx76K8RC7he2e5dPPCPRIUivzLQZO10iMzrKo5X0uPX9+QKXocflFDs1D
2B28CW1nr4db0GEc48RQLkvhyciXmw8Yb/hmvQ6/2icjCoSOxXkhBSXBclLfDpZC
3smAuzCZ17xJdTm4zsXxA1bD0ejd9daZLiGMRgrORqeB3FbcNlz2JmwAuz+5wjJJ
SaOBEydgChEPYctkSJLmKUyamECMlccsLQnQmgsBl3iHur72kMrx3fztOeG/Av/0
QTK1ul7g/+tnCL5yabgsJBLfxEEed0IPnpwRzed2n13EAT11CrWUwfEYClHbYgwF
IkXtq92q8WU5XhuYXkd5nMDeqduPcapBhL+iL6btXG06hWZqbpUQ++m5oMfRpjt6
dNgAYb7B+xg0/vo/xSk7WZgEDAgxPtKEMsB+58+tFpMQaJ9J5Kd8JXbGhQIbUr+X
oSp0MTu5yTNwri0mr0I0m9l804//l80bORbnNgK1qgNQxQ6gLZo+NF3znq+bEK/t
zvN9xXBS3PlgYjee4YK9VU+bvnprtFXp736alhAXVQXZ43V5ekLkbCeRfhVGI54n
m8LHV3gvGdivejb93r1UjSN+K0vNg+JOY8LvcUagEz1ZQjZcgeF7KwXp6WO75RfF
NRs5GoxK1n18LaWuwv2Jg+UQXFN6HR2Ige5YtD1V8ViZlwTsykuKF2SW5B1GBwnV
KFrp8hg1s5jrPwCBStYA6eT3VFTWmF3iRjOMdecQjp9nWY3v5g8rvDM6PjkpMqKs
6l5K596nhirHV/pK3JRhxXNesxpxyF+7pGaZJ4PM/ZIYjjvY6oOaWCkiHN89rIjm
DCJCfIbhkKCmEHbIEMgKEeCstvQ7NZnfOwVbaE3cjj/zHTUf3J3GLTL9UmxphEvn
FHZEnp9maxi31UQsXxd1YdQlVUXf8rqWfey64GALN+omE5j8OHVzX1aU1Tc1BRR0
DuG2n8SXCpYilmKVulo4S255LvNYBQ8RhT/hSYxVIwrK1+I0/8ML9NLCDsAykQeA
5GDC5K3TRNkMXCPDkgoANeDVOsy9bD8d5eOn8OC6IMkJiSkO9S5qWcqQ5KyHS6uw
dHaxnU5VHmp8wKiYUHuNFUeqDqitoLH3M0t4OeLxOS4E0kJBP6Q4oyjojTdmGUre
9UlmjumdZn/Owr38IHuhEjB5BtyoWMJemgeJTIVqMwWWbP4FRqu4v1ncl/jXK8rI
OsF40VcRVVqrkHTAOnIOper01DFlPQFOHMI/X+zjdXKWIl+COupwjFdxvoqcUS83
/xlRCL8rsCl2uZXFTmpyQgzAwckFkAV+L/M+P4Hd5QPZ+6a4FlqAHe5vZFrvpNBd
lvsHHuwC5caclCNLOxR1BwdhlfZzHunKRmhcxMS0XnyTzPr/fIn8ay8u8yExtELw
6uQD1ZSlEI2qdeZzJE1BKLEICuENqRUjxjTI07Ej71+d4NzWFfEeFx+95GIJ3IaI
0KT/Hv6TCwsTkjKXHzdlT3ubKsmQ8r1yi0rHnrg1MC4wLAGwGIpuyCZxGwp/eMdv
QscAiy6tN0QEPuderfttVe6vG8xdkEijmoVqLPHUWpY6f+NDX8W14QeXXAF9OnIH
wqKjTl5+pnTLCpQ8whAyr5k3gZwby8O+iX3RqdlJ88RiVPVhxdU1S7U/KfN4j/2u
XixaIFzTH4fhgOKHj09o+BBmKDZT04QxNCq7O/9CLDqQGm7aBKxV7EzQ7wQAOAoi
ON5HTekw0EnHW2Gvlzes/lr1ZK/OLCUBQtWKkboflN4QLKNjF7p1GRgwjMttSR+5
BpQ6M+9KQrLZXh52FKW9i7MOCmwDm4j7P5FxGgRf09iZBIIncLmmw7XFXlVc7XAk
pguXpK1uB62wz8d75W++7HuSUNYU4YFHoggGshGvs0n2uDYfG1q/4UH3LFqIkNWe
V6owUaOhxsP2c9V3ybOQL/oNfHw+D9a65pPAzPQJw9xdhgGhUHfnbC5VLjkHaLEd
395JmerKpZBlj0t3Dzqqv4SN2nBz1gEH3odh/OhYknURnLh8tvsTgcAn2ZY7NyJQ
WCPgsX9zt1IvXARnpGKr3qxbvquXYPdSp0NQRfWIHNIqOk5bLVuOPdDmv/qtQ6Uh
srgORXk8D4wV2K8Ld84KRxcxXQ/Cg07vQQzfeHncVjAuxvd+K5c69uK5+UmmQmZG
HMykes+KT3bj3VB3tq/DcGSrje+dHPfozD3XInft7QI5tbbvxJ/eUyT5DO9KPXNK
nuHhRBlkWlPg/NGqnrl7yUX8PQJUOa+L8BGmscI88ADwOZdD3BASn6STEybRZKEO
0MMxljWVfljdnH4ePFl8WzPY+MVdR0dYeKex+WPx2yUoBb/LgaDVrCZm7eg+1pI1
qD+wPtmVgip6e6sO4YCNc2Y9uHU9KIK7LMotUTYdT+w2DukjunabKFGc1bsgneGi
bcxW8m1YWtXJdu/uhbMvAZxnPeTIqVoykLTxk1JFPG8QR61y9gGjiCBWZxG6Iuhd
dBuLAKkgamYGU3rgdjJRR7k6eeTWik53pLQseFBhF+NHPvxc/2Ji/qbOeb3tHJfM
63uZODPE1cYicl9XKMQGrkr5H4SeHqiLX2hhvg07bXoaqlqE6aUk4l0DvxJ/asza
NBfkht/EDAtU63q7lAtRHURod3/fZR59P+czDy0ccjJQ8+SXBpNWn35a/bdMxM5u
oS4yDv4AOH3ZU9k+MK5FiGfhFNhW8KkrvtZ95rZl14Ltv3xz4NBEyGrgsqRBiRC8
UNIgFNZRvSQWccGB3KTrXgwB7VVjytgvqJIHDaDd6TtObrMNsYy2IIYffs60jD8X
UzEEILc0if0gEZOxWBYf6HpLDwlnjciP1wc6Pm9DfbrgIPh4/93enGwgwrzje4Ut
JKZjlenJ18CjHDvLqNiFf6372dk7l0HcxdPxYYjEMZ4MvQ3h5AbY6qDubZgcpBA5
oT+mr/mQDcOuLILQ0rSvBrGoP8y9aIu3hLEwO0sSIapKVKVtTx/8JU9+2O6I2GvD
9JG5l6J5O5v14FL1dR8KbQxpDl/EvvQzyBi4KhXhMFB+CBQoxR+0+lw+PSGy19qK
wQaOYqiZQ0XvZUuD4THPxu3OgzIgtOW3peOQVlm73FJjlUuiThA+BrEFzYoaBdPO
Ih4htkjGUdHd37nSXx0tPSkDWfjqEJmX2FU65oHWk4r0Yq0yKSkLOSMBNwsOnH81
83EsRtTV9bY7xOQHdevYwPHwba11PBgTuley7g7X4UyQ/OZJdIwymqI+5vz0vUiC
k7qRi1PaLQxPmC7zsRSZ/By26/rRp5TACP+OmMGwlxYPEuWE/o7QWKnHZntmBc8B
1j4utjBeY6lmKJ4K+sbnKl8D78F1Tlg5ubjGiKIkNKBPhVfC1d3coKzNBcp740oX
PqgbFWtZ3TBVF6SBwAy0tozpWJOqAG/HLvbQA+tj1R8fpTgz5IshkqWcO9sb3RJs
mnLaskyLuWu2nMDCtpMf3KZPKFFcSC7zDqYdXrhraRPB24wpFEaRgXFXuO9kM4QZ
DjH0zM5UjEwUxLaSN1vffRMMCuWkZbc3gsNxSMlCj4P5IEnKOemKYBsWcNJX4mrU
/H6qxn+3XW0+spQsSYiEXiO/w/CySjPL4zWfD0qofWdlykg62D46FLvL1nbDXRmb
GlLKeXyrAMx+PnXAUFqXgMbhVdjhOsbP5F3XQI/P4o96MlNyJcTG6oZEatzFqEbB
b6sHqL3XM1huZZP0N1QiC+ho6QDjNvrFndw5Nf76UDxL+8P/WA16PE85iwlvOwXW
C0uG+vWIzHn2vcuMh6Trqb3wwvWnl3zaZbqkFNXpFa5N7JIyXqlXWJDOp9EJE4C+
gtdN9r8MgP7LQYmSUxxEZAHRbh30cXg+NjCnd6MxhtJrgMJ0sFjpn6MtqMQ/EksW
A91Zr76dxXmOtWiP6Jep49oZo93mDrrDzz4ySrq1DHpvI7jRcNvfwXa2lIoTzCHy
Q/Vx/Lwz5BfTeSLV+o++L8porcI9kO03krpR8EpWB8AO7k3zsVvdyL9GlCHe99hZ
NHCtib4MJzbRzGkdVvYd96oFNdtoh0NsTb6A1tzcgWnAWPKvt9e1lexVqWL9nIB1
GC5J+m6dcjdp6BJRsuyWKVSOFZ2pUP4cy15exW37SjZ4C7u7i55y14nsS80eIC9I
hnMM5WSLIQ3OlhuraA43q34VWn8jyAKuooqPFysOeXSfCBDDSOWz+9xB/Az1AC+U
l7bu/Mi19Az3/2P+SOMv0HN+xRXEo7IZucAkjmxQJWTGgIJr/LAmFnIFx5k8GyyN
E2tawsCRRo7F7fgJLuEY7suUkyHXho2Wt6YCe8okM5yXd0W17zRr2vtNa3la37Nv
YE807lKdjDh+5r/vDmWfTIZzW3yRwswGnz3gSdLUr4S9uwUJapRcywmYg1Qr6UcX
zNGGdoLSMUxG9uW/FnDa1eXBmRROGQCcDMeRMbWEd1TKuZTbHsQzTYwdx1rez/OQ
jHH8F9if2rERJlYq81Qr5t6/fXcCDvGDLHsHW12J7DvdQVxjtM6apqZ0t4l90gKw
ffzWyHtHayd80BoKUbu47gpUQb+kqObGYE8yHV4mD+a+6SVVTctYyI3j2vosukmV
2Bl2Zxru7edGq1A12WZhaXcnBoaMLjJwBwLDU+jt9vXGioQdbKkddZYuUP4xhx9p
yVdICQk792SOJHcvQAVOxvEbkbLFZuS79VXCFw1GJmGpIpxA3qOV/BrT4wti+N3/
rJa1R6c3WaJ8Bm5eJTNnAYpvHv+FQJ/QX4lbE8y+Gk2PA+ZO7ii5BosKywKGhU1U
IleJrvY/XjeySGIiURr5hHvyHfnO+ZDaTLaKeFsKo9b5tBG6+AnI4ajTJNwLG4sr
XoH0A9i0hwTVfPGzUrVNVWFcMZBYNWxWVgh2DBagbKYDBEBsj4oOpubw/8EctTma
0m0MM7NNvOh/+v8/V9AijnqglhX6G+6ClWQyAYPiAgUZE1eVVOnpibJqjBIXpbbb
XgvpwLJe8SjRQ0lCTwtsDQfhCrX3IXE+Wcng4c8sCthIFPHITYVh3kB7M10gvZHi
GRSfI+EoXiNNjoVCyNJdGHlfzDPQc84TPxFD2Y4K4k1ce6zXkLP6JNde0ETG6AS8
9eestLzOM0J2tsZpTcB3xBn6yoiel/7DK6YkqAczBkppmWQgmQ202xQMksqqpN8Y
GztZ4JQZYK3HZ7CPN3TzoRfTqg4hyzkHfwxYEXyHpbRWThTGFAHpyW3uIMw5OpHJ
4Sl6YhUbQyXkvqs6xoXJRuPb3DKqWmg3Xp5smlIUmZCu5i/d/PD0KccoWjZOShjg
Ep6ne0CNFH5d26jbnvzZqoMyXWtEQi46zObeKZQF7c1hU4jq+0sOmXug4lZ2zUZO
UkydRZo1kbWTpdNEOgtPRWmPJ/CPP3RFM4KwQS/izFLXKgmZ+s4oQ9vkfGDh5r/k
44w6O8RsF3H7gbcWM4s2TeRuNK4otE5vyGr99077ZdXhOUm1voafAJ/vHziRgZhr
ja/1kHQ0HoCQ6rlZ1idiPYmBhUSa8lgh+l3o2YQl/LXibKkTDvvo0AK1uaDGe1qa
H1CQnPxzMsyp3p23k2RE7/8H5rfYOMsQN/uH55ySZ1nC56JDsdyenhs6GOzsvlYq
u+Z4EpXnvHdHPNlYYnI/Qj+yuOjGNF4ZEUaY+kdTMfDaXyrSRZoAUJs3SfBklvkg
5zC/JeBDi8RlvFQwNRA/hxJ37Sf+/8fpiirtITTA/O388E6v7QXuxYFAyBHirefC
LKDlrPvA0RvUklWLxXQ+piXT6KZK/ZgJLYfc6CnnyBg3JtOM+QjsZ41sp+wGcBiT
9+8VLSrX+fErEl3ygoh3hXsLyq9wRV49IuLkkcSXAW11Qu56ErIBd3OdsCBw8wBZ
G+0mfC0mCtzKev1KHPOch6h00k72FZevnbbK8MfVVvGm5cMYdvaA2jXcuRJMr8Ei
JjKXXJQYeAk94rAGAeNKW3Bg3Uk2W+YPVgRAoqwMi76PU0RTJxufG01EgRZVJvle
4Pqe2ZcFn5hHic4Ps+25/wwfw8od0KMbFJLCTHmDXmvKPBBmdMimiTvo1Q3Gqb8R
TwYaIE/SxUPnRZl43/VyIVH9LS7lsiiNIm46M0n757HsqBKlKtSPWVW2fs55Hz5n
XbVWjYa6sh5DwF1SrLGztntNcLX/08joowNiXOug49DCRqSWuBKES2u3lwY/277I
oFaLs1MiNfhF6q2SlKSTiR7JIZVsy3RRGa160HzH6vZIARkFn7m6e747itOYlg9y
Qfg1b2izWuRcuOigMztGWz2oJMwXWYK9ufEeaJWa3Pjbopx0sUE5IivUn5lohirr
MvKadZWdKabCqYxPqdXOIobWVDiNqWw7QTQ6vGCLUUZ62cZdc+eFGuEaKYh1MBxP
1+gZW/bXs4V/+T2iHeCLyf5a9CCg1byHk88YLBVOMR/uny5Ddxg7nMGZTrgyVRhd
PHGJemG3+XKzfMqU+2ZFsUO1AmFW9OsJY4TKuSXuX+TrAOgmCa9HNFrc7CdU/3cb
VNCDkHCUVY/F/AVHxYAXjOh+vHUBoIO7hOZGd1W13q8iOR29fgLy0tOUzyxAs3YL
hqQM8TFXcUz3Ey53jv0S7oeg++fHBm8dVgquWAvRPCuQs3rNYqH524T3N6z1IzQr
2apz+2kBNl2DNDa59YYPCojjAwzTzm6NnMH/fTxMUklguPItK8+ayhddNQLnFCIk
FKbyDUQkZiZoqAyAcYPfDeRigl9/rLUdqxdD5jlhU0AQZ1yLfI1UJj0OxbzYK3+s
ews7VT6T0HOBcVD47exU6Ao2PrJMwgLiDrb/5YVkrO0/a4MY+mOhqfoYxxb1DxEo
XyUjEecMKemZZ7OY9DJ5tufalGGrximHMUhIH4uwIE5/cPs4tRFk4IO9Ie+jKES4
Pg8QxFu+XXuk2qL01gH2PbhVqx8ugRJ2Hrxt3JkI6Qk4s+LFCWBF1NRu/Q6HNPF1
Oz+Cy2ai2PhlaM7zgDXGB148euraglAOP7WAqDBR2doFrl9HwVKXw7+U3xkmXEbK
36JFB7iQsOak2tndisqNjWzZhriODzUxZcziQcf0w9zkRVjubIyX5I75KnI64v4N
pnyz7L5NW9JJReMDBNnRTyJzHAlb+RRDUkRte2rXQ7LVABUOCC/MBkO13T958VGT
I6KIEPYJ3IcdmD1L7oR+U+05jxjIXVLRzWXcx5At980JD1ufCdHXP+vxB8mFsYAM
LXbAgToaYR084LTzTXbrlJOG7VOdTXiLUv/MIx3sOYLR75UUehQzTQDrqQ6l6FKU
ohhbxpUXlGfQ1j8HR9ECI7SPFFgcNkovOUpWm0icNNVuMNdvI3FxQW5RKPvqYhE1
H9Vch3wPBg5IxHxNB+9hPzZ8KSiOzor1WVv7Fg84e2Qq7vSosKOFyfjJVU6hoT9r
RfCg6UW4NgHDUX1irkRp0gbbRJk8wqaK97JvG5MyNLqhFjwcLbZiBp4uC2WiDeIc
n6Kk4cpHcvC0LlHxgSU/r+Oi65xWbzOjN8rYVS6xGQCFo6vfYwzDQjptXh0GgbDX
ufIWHtMHjQIA5OJNXToMgC0dpTdBRbt0khPKIC9Nt1JWTJxriliDyvtYO5rILqHK
oTBMdomj4SOZeHNnJU5ppRkBVVzpqIdjn/jAW7xweQYgCg1YgoUeU2+/DoqiU6c4
S1vfS2E9BVMt5oVL/ulQoMOesGW56i1sRv5Xd/6YmhWbL+3Pwrc0sXtlb5Sanc5c
AJKuFIZB4RPzD/A4dBraVruU8O37OrVlLCrKORua1stB46TVTEFNVROP947awpGa
pYh6QmAjygTAQg13Y4J6X6SHIymmi+SAyJ8DeGYvvRcz0SJYdCPFFKzj4uM18nuo
X1SS2tS2BscQV9JqCthf8jsDQwIwuyq0+MN6sUbXT08dvLqu81uqJz3CqvJ7h9Uw
CIuMm1vusVanGgqs68V8SvPbXybyrf+Hpvjwzg42jQNDCSoFdhl+ZXwDKBhxdF0Y
wEXbbZWfRkN2jr1/E8EArRhUCtiYS+ReHJUW78jgp2T/dZ4nTeiFfbstT5XLjyLz
cfNOpOwju4szJli4nwO2b13xyDlAmBkTGdwmaVQbZw3QcCWwvjD8ylnKW6ammrzo
WdRWyKQsdnMoOKPAsKU7ku4enAX/ENtG0nWGmJuOU5yX0vCIoZNhVxEVD8L61SQT
hk2RF/4yaW/4Tx6QSFL5GKquf54GEzQPoxgbg2ZF53JsVkWIvJGjDL7vzKCLcWx6
ttSLawcLq7nJ3Id3bZI1YRIEpu5NKBmCE6V2M+M8q/5pXMgepC0EDg5SHZo27Kox
6/T8J4uC51MzVsMUYCtgbrkTuo/yl4C0+/OGETO5DWf8zG+/WuUxImL+RxiR4JLt
O3DpNv3JZ5HoRnlKFxRX72OWqCOHl6v0ZkrcepospIvPFXvn0vltLJb8vx36VkBq
Tj+j3iD09xVRKA9SSTKrv9b+OGZUbNwIFuJe0KNzgiiegsn/Z0ab+/PGwWkC3iOB
GbcEKB5bjvfBazCNd5obetHoOhKlJ5rl7j9vR5q/u7MBALUovWSrICQ58tbA+uI/
3WDnTzKYsRfnBHWaXS+OLi1/G4kc3G85XXgvA3sidpwDY6l+lctNXS6LkM3hwefm
e0YD5F9M4T9C+xXMeUbHZ6m6rVfp0OfjY19M3lCvhla1aAw0R7AF4Jo3KlUSBhFz
sbTi9ekYDaQ4ty34R1Qa/+r5TdcaRMNEw9bodT618hlRtEZoDlwPL2zZVoEyhFuU
JngQ5JZecZgS2qV/xE0LE4zjUsLGgkiHikNVus2C2Wtvg3fc2hrHbgcM5sVitmDt
z2QrgXNA5/Vw6RhWDbZ6MNHMs63UpfiFXYoGpHGpcVZtDQg30wl72lA2WP3jDoKf
at8J0U0LaFQ7Sa0udeBxuciljk7mvl2Yv/4vFbcRecLG2vs5N+y18i+oT3Qix2V5
J73Med6GYIaIC9H/RaanMDbmcPYa2OLCrJaCojrru131r59IzeGSCgzAbDFDROH0
X64ZPRGQzGLYodAKe/ZeWe/5XyliXMwOrjxF6c3nUhBhZONYuOVPsRvdZ+nhokSw
I/L+JjB15703x3wsphladkWt7PewmZPWYyvx8PFzeiwS4198C0HO5QgCmiH0Imxq
4IBiQ4qfJ9Dv7joNU8cIfeeLhb4DTUwSRrbEPUP1I9b4hpVh9U6KdjyQoyW5fSiN
mJc+jzhewDdGrxvro1poVyc4it+7Izav+fy3+1AJRPV/TVGnzq+SPbduY0avBbKZ
pV4NBBCAjdxqlcfLy8AdMIdKHens/Ovn/PUyawcVKlw/IG4wfyhsrZ4dPPPJs2zu
/uYcyOsCELBMd3+rLfeGCQiYPxud4qToCD3JfGtCYzXncSeyB+6sQrOYPuof+uI/
QJX94wskijFjpT5v+XVSY48sH3UCmlG6kfORTGvEucUOKvQ986Q5Yx9/T/iHkq7N
KIk1rwBOKoPGD1hm+tnFOV6Y6K39bGmMm5UXI1oezgomrshmPRE4eiEQTUbepYCH
sEYjAk61vUgDVk2HEdLAk4PZESYaNFIFymNE0YiLfSoHHA98Aucy7jSptEBRhq/o
HjZpbk7k7BU+aF3oTFtxkqjJ5GXbtlIxcim0y8PhTfOcyr3OkiQ969HFuGSk0CkK
eyGFv5js5YKeatDf43h0x2FlojTYST1W85n8n64/GMFss+UA/Dwept08gci8CZVP
KLBP887oV2rxFtGEwRhtpWNKM9qGYXXLp+7Xr3YX2DvKEMp8sZazO5ibzKg/ZMsO
9DRYRUIgANU4P7mEGGJJEpalOZU8/TSE7E15sCt0kA0Zr37msMQzD1ptHkRCY/RP
e0fvfNCuSwIuEH+zTU+onHQHytiY85J3imgBJzZzFSCtTVN9qncnCPIprkweX5Ei
XaDxqznNeXzOzrLtIjcaFLWUqkRXucA8aMfzj0KdH00ovj9NGzrDBoqWcWsPRqVJ
wz4Y4iiplc+DEJmNvIKaAORga2n4FVIZCN2O3uXnEStEfJLG8b4Wp96dFGilB9SO
d32iI0hbTVshY4TMJTFlieZ1qwnxKaB0tIgjsGddnXgVELhqowh5O2gJM0PRlTND
MCiGpchvadEIfUt7335adB10w+s+Ir9Vl5Qwc4eFah88XEzEz5DdtY5ddgBi8sf/
2Khns7yeIeRvMiGeB9TlwgekJ3l3yZ5OqkjKgvcZOdNBwG3reokDyGCrlnNhebVR
bBUuhxu+iYOMcwwGBPqbeVxM1266zjh4qkMDvamfZltqQDKi+YI9J1l5qoHd8qtE
0brYxH48V4Ck+Qy+4ir2CgXfIc7zmEVkgbGmegthaicXv8pkXBrajEZfm+H2ef1k
kEYmw4yXuvxpKh1G4yTaKpzl7cXCvsCL+JnU9/peGX0dSc7Cn9TKr2xmuVBMlwwG
gCe5iqmg2KF3MuIgngC1Sg35nWkWUVLLlg8oyUcPL38MVuiDVkOHIJhPyKnEUKe+
jrU1MCyCeud71ibQ27Oxs1jhkJuSM934nztJ0TBJjQc22tnpNB8tjb3KLpZ786OY
d8rmjJx8yiaNV0v3p1+vAuOiWzF85F3v9T+m/obH3OssbwIfcVwFB8awdz1dU+Rb
FgRNFqDcYrbzJJ4qKbNniFUB5Y0z9XbmuSch2k6L1jYeEG1Z0Q3k+0dhCdONd/As
oCv2l3YM7+BRGojYsHef6veq5mZ0x2WK+7bPAe1MkZLn3W5Lx+T2YDqMn9XQS2nD
xsOtn7C6JY7od5zi7wEo9LJqWMGe81xXiEEYE0YD+PUgIIP6v3xglDGLpW0b3Vf1
AkTmmkKoL7QBzdYcjwJfc5Jj5Z7IWSIkp2hVut4AuW/Y6rrRsr8oi912UmP4gzRi
9DCE+HDYLsm7eSYOM7IVT8Itvrk435YSg04hpgsyBMBbvs0zhbf/V9CJc0pPK2/e
umrRH0VOeixZ0HKYuP7v3N6oP66Cg5y8jVlqazpQcdLEDi1BTiCthujhatoZ1kZc
Ug9/eY7zG4PWKnhbyaKsiSadJn+IoUvUb9zRNv6k+wZziM7RlVvj9+CDAS5UuBAs
edmN76K4NOBVg3Wxxx8bOYM1N3B/k/+R4K8kHLjlO92J1kHbFOkORBoiwbycJLPe
XLHWuO2t7bdqwqkYEgQR6jg/ZQ7B8HDiyjthY+R5J7sVg79cR1M1xjX4CuwQp53m
sWU7o5UfQ9PtmqDctxYnz8R2LwRtBvfGl4xrAuGYK1Ey6RC5FeKPp1z4N+nG7cbm
B7jbAKJOZurklL0Bev1gditwyLZDmRb5Q0Ll1rKZmLy6GEP24MPfC1jh+uvhPlRP
trEvx9Pjr9kjN9Tj9SfJDBrZHRRWqEdhTznAxrl4B8Gc5A9g5gmpAGN4SRx0cUdt
Bl00qK4wXxB6kq3I/Ia2H2mL0CviYiORNYrHTIsDQgd4Um6F/wkWJQC+3xlV70JM
GccAjlqlaJ5lHALdiKeKB1Ra85mbS0+bGQigdGLp/LsLmLizUgpIQnfvZGtG7CAW
u8/Y54YSu2oddvo6byiUdUF9eiapegvHAyLdj5hmjwXUqXOaWOZE3bcwDQOQ0x6w
2jLdFf5/QGJ93zYQbz1LznKtadJJqltE9WVMNFOtwYF/3vPiEc0WUa3HTmWgi5Xo
Hl5nsAxcf5CmvIKmIotbQ6O3IHt1LIKc438YaI0NQ5DQQ5yi10U5DI9ff3dI4AFF
gManBLso92J+Ojl13p7nM6SxtStGNE6MAnP78wEvHavwuX9lAdAb4LFK72upr1Xs
ZkCrHtTr0op8fCDcb4tCXuPz/rs0iS4kizxrNRqMKT2+zwmFBmDHrTuvB3MtcxeU
Iu3bFGWmB+JzlRFXBi/9Z1Ek2rc70bHlp6T7vYJC4WPyaKiMLpbmITwTb2aaSoRW
7bkF0uT2DC92OMJ4/W5V3Cz+KB5V1bQf4SWM3mFmSJzH1/LmI40GlSqbYLGp5HBe
pueA+/nS8K9YXw0nw8nfgjGobkewUbxUnXdYCw1BY+j19+i+a5mw1PZCfg6Ovr1y
tHKPNxtLR7y5RAlqcLa3tHNB/hjU9BUvv0Mn7jOanL2k3amo+MbmhjWpmfsWUys8
rH1cEZCXynbMajRYm9S2l189FBim4MSu7xf/pz49M2KoutqD8fL8D6bpJQlnMrNi
BNWKluGESse1vzkqYwQa+D4c2vclECOKD2DbwWxuu7B+aaS0V8rdEsaX8fAZ+wLZ
CyO4XaQT1PQnr7kqlwfF2t7gnTHUh+tOQyewftoWomh4OptXTUM0tdpKX1t9ibB4
JddJ1Gv5lMAqbJPuSEfvRvE2hQ0QCzEvK6eHZ6HkpQl5F45ZiUP6cpreQrmVbkTQ
PyUGHFqic4hBrOxniz0SGw5GHZIrb6OXyrAvUNoUkSPEU05I2rlkexVrUH0H+VeF
EvpcCR/SPeNDIQi8U6mmS3SbZpxk9gqeTqevfBaWUz+RS5ZDL+UJ7aI9F1yrHcwZ
7V/TCIw9kdPB9Nd4icR776wVNjE1TJ3nlN4c4FT23zwB8MpMpWR5S3WSPMB0VwlC
YqXKekKje+IJ8c5Iydao8ShYKvIB6Bu3C25rNR1XHysuU1cDGalWMsNZFhiPWDoh
2Ezise4GmYTLaXqrKQMHfjBJz/hBtIky63pbgmLGCXazHjgciQXc8aMxZi7mYpJq
nwmdt3A5iWDGfrlaWdesLWZeOCeygUqB93Ls4AtxqqUh+MPcZMKMgIT3sVaINFN6
Kaf2cwlQ9Epldil5lzMH+68rN465kHMQNbE+J9rUusFr8wvC5gO+Nj8dtqmkS6Im
Jhxulw3BRmB0xoU8tH2WWSRDbUvwZi4r3lktKi9/LuPYzLubLnAK4XQvArDtpC3+
aJTU0eEb5KGm2U48KX+XhR/Q6AdvNjlAHdekmzpz6LuKwsGxAsdrg62p4beBQXjA
NzqENOFz+dUlo+Pw5mPVtfWvxLl7E2XqKkiGlkqBlejj6ycueJEXjQpUQxQDYD4w
kKO04CkJ2Eja7pQaM7rKjNulxQVrl2iJpUY4njWKPsUZtMCeR+kyXGyBmfPRciNe
q2Hwk1F/6blZ9MNfMnFTT6yr993TbCAhMOh3dE3lgoPV7sDeMHby//CrchTHpPHB
QPkVq0DuE2ssd9vBjRrlOpf+xa8YVeEli/iIKDePBe6S/4pcUOIrjKWjESGnbod/
+E4o2ahDq7NxFqkpwOqlt+DyAOnZV3+SQqE+EQZpzr7hHc1BITLzP6054SPWWupS
2vtb8aAt1/+ddcn1CpMDk6bwK8rN9TZYtS5oDtiTd7vtp7WCF9+HsLz2x6H25Tdu
k3yBXV0Tg+c+rRjL1zxVXy/nHOLAqaqMsz2WhVMUy3kHqBwQktYVJfZ0ZeXnZ/wG
t88uo1Hi8tiXTRqb7Tj8kM6GNkpdaa53x/iHdpzD80R7hqPp02L/onhWjLOcexTc
aFFktowVHBwiLvTZznJyBVe7AgUJZdq2q5xh21VyQ/rMZ8OQ4F+E3iyWgdp6TyMw
8ZWKF8JbGGuuYnx5Isgk0fUlfksAKJlW4i5Q5XaGVfxbh/KyFpUt0hjibj30jDze
+a7RYy5FpUfm/xxTlDcOOB6rxAploHUAWNbuWwkbTmdZobakY24fvBdp5+3RhLZq
2W8o8qglqF9Tfg2JaG8RoRZmUdP2NN/ORxqAtrpLaAQog65/bacoabCdFtC5TC1a
jVY8YpwQuzUu+I9oo+CVv9Jd8P2X7bcLBbwOWFE9mAh2VRwq0CLp3y1dqGDs+Hqm
/+ydF+5Kh+cv0oSstBRcv4YM30Dy/JrzDzSW3MWA8Wf71iarFAtLN99yaEVk6Ug7
BkCWogHd7bBLeMHxfuccVOW6hTT7hacnRD6EkDJfxnV1UMkoA0BLtXIUE4ZevSMY
+oeCJo9hnLaFBGD28DEnLaS0K4lfvKCcjIEoYx773aWvK8f9JdX7Me0kdRGrbLIy
rpJAzCvYIEYhdZAdXEJUJHdEQq2kfsP3t5HLbUqIQ9YGVRjKWDy7Xn0asbVe5tes
eJBAks2+ppdiy/86IMbSx7RXscBAf6cLx4dsGlyzLzyTwWE+uL/FogGUMEqD5Yk8
6WeFjbVKY0D1Y8Wzh4pHnvJdrywclN5lhxp0L5CntytgMqkZGphE4txHozVE72bW
jYDXHCR11QWLuSDd2/7MuWjPVY6n/BkKKbGbtj5M7kgRIFU++A+fTMtf2N6mrZxL
/9C5IdVh+DaWRrkyXqJR7ygX+rDXvxGHhiWYXVYQZwi6LTyQSc7PabH5YV67cLpH
SAJnDxatbu+rYm2S+eHiU/VmsPVDHeCkEgU5GVMrQm2+Hu5f03CmWO9YnFhvFEdM
TEltu1V21KPrGCZr0EiKfO54exTOsbGabZC95EEz5NgPB6YUuUgYRE+nfw+fyHVf
I+PfKy1Tx7F/Y2eCfskz0IhYhmx8fcv9ACvLDyq+MKbAHSpBo6fmbKS6s5/71JOJ
KMT+ekpsxOj502Dr/8ijlSQHT+iiipGN5rsbYG7+u4qxGqnrPM8YmMIXytVQ6Rw2
J0pFCcbPfbtH8uqwIksKFRuP7XbP5PJHLXdktDgqztTzBSYpqy/zQviKZvDTsE6I
1OIdXTc/qkVgV7e3AisokVclkPpP8kKyGB+BrbESNeA1y8fQKF0n9dX76p03Jkuf
uPBEEJsZjCtXP8ZVaCk2P85CRRmDfxkzwUBc6IcP98TPv7uBrh6I5O8JrRqhF3rw
z7188mvHS8G19wALvg43WUnhw92gyjkrVXKDuYk+f5GW/OSZQ5Z0lhPBkI5bpg5E
xJ9Fgqd/XP8+lHMJISWuPLvy8ZxQJVqnvKIwAjK0lz54YKXDH3LAp2+9COZxfafL
ehs0iK7cq8vslBh1CnE2Cw0ihyuCLoWecTB/mMeTp7z28Lr9JkpjFIlR7bwuU2Md
4DX7Aas9bfeYEz/3XHi+u2jjIVqGZOfYwqwsUQvbrQ1SU8GmcA9cB9UifZ7yZ+D6
Y/nh82yhiVy6AJIj5rDcDh0Jyu5u8ArpVt2tWlYMcA642VNHD4BHPz5MdrEV0wRm
R0/lGuQl9WdtYWvjTOXCI3CPUogu2yQU51BjIc7Y2qyQRSIZBWSLsfY/tl3eG+gA
nAm5HK8v9yv2nWQ04teQVAkM3RioX1E0V+/8P9dPIegLmhyaZlyvSdlGm2NSEShg
fCOENhQlSp/B2T3x8KDm8dUP7bHt/j8TXN8YdzjQPbuBwaDZudQHvdQEk3Oe0Mnv
jrvVRrmql1RXu2R7Sa2fTxSv57ucq7219jq43GxgqRCr+p3BVS2Sue9JPC6691Lr
fsEmUCyjIYGEgJVlWERZLudaQjLwdyrcc8rBLEZizrdBKhmvpvFrGBmJSHNpifmw
VbKDNCTqvNj5wre4YbSxa/lgZvgMNSTWwhq2zOdSquI039SIdsndeEgA9P6mHgsn
GbxOaanlO3gpzZW73BgxKguHsXNg2i01lbkXZ4fRhj+mzISpyMWzM70xavF41def
aWaQQ5AdE8dhDdlQALu1UlMkKX6aXm5uJtE4Bx1j9rXGsHShCwNRWqgZvAmSerC8
/UYgkJeWU04vZoeFahoQXg7z5OmIyvM+snnQVCEWAVsL6kh0DTH7fvrZFFTdpaHJ
jzHfAHEwARyPbH9v8Doj+BK0f3mGjaGIFBETur2pSDDhF0K09fOx9ogc9sAHdLng
Akd6K3WQ53s8tyge8ZrYDWrnRPkaQl4hCa0y9gi8EI6FkJs5eA6Lv+jvIMUCEbSR
kUkH3CjQVtzaZSBQ37NkoCgz3oBu9iSjakYOR+ZhKDLLPgY7lTTc1k8rleX2ujxH
N2hEA4f7NVDUh+SxCGkY2WQNn6DS1zAy78AXmzKfXKzcUtzthROzTUsmDn5UbtZO
1m63xjxc4c6IRpxtMcUNaF6mBiRaai5KZKrmATY7RKT47ZQL7QQE1/NIUmxh23JR
a5qziw1Xddb1EQZU2deX6Q75LFKJswTk8iGj0Lzzm7FfWFolLtaQ2vpsqETswPlM
7WczbgTHr2OglWs68Xtkb+KWrGgCEqgX4CQRUWXpEH+rxDQxBtSIbHOkGe23EqEK
p4INa/vizJp8jxQhT/7vd+nthOvoXGhQpgf3JC5KAKP3cG26vGXElXjYGQItQ39K
X7shbpANrPg7MQgPYUCPR1Zztkffbr0Cq92FyVfkmB37CSku9viKWmBX41qb0slv
P0aVpKpJ7htkHgXusn2SNU/cb6VunQSSRFvjhBuOlbCI00oelYYDIlZwBc++YwPm
cP5X74AkkT8HovH3ECCQTCRoKKMoL9r+id6K34KwVi5gS//ChKZpdkSt92SBEtBy
gKuejCfpYaeIdneYN/EFJBUnXC5zx8uTVs0RlapG6+RfoebnbS66dmI+OY2Yzy1x
IV+PdQZiYVG4i+AWgiiqHaYPNNfaWjCkSl7M6hVnRBn/+F45AjlYulHFUzEgW/u5
KhJ3D7KKaVWFvlaw4OZp9c+LaeTMW+LcATB2nk2sXSMlAmCGbbOl28T6Vhq00odb
9E2BNfiCllZ/Bdg3iSf5hlOExmboWlXldjgEMdpmxmJw3Ga3zaBuSk9XtKAdx4Rh
eb7VjybNs1mOR7rfSmSQ84Gl5dibEgzR68d/w7JrdxLed5k5vy8xRuoI8UGUmhRF
LOEO42+X9g8hIeZt40MMa0kkI9ix6oAm2AOdsXWRX0rnhMPm0z+cTXjDBnWA+QpJ
OFl2IIzP08hWYMsnSLHUlYbpt4uHDX2bEwHC+eOCdlX0uDoC/FqkGcz9MinJ7SX6
jeftTqojxmcao57AWFvs89dqRfESBO3dp1lvI6d6Ctgqn98s4Wjl18/pyYAKyONU
qlkoeenykPjtCy0NienYLCHr2Tn6d0Wab00JR3WqFIW7G6utqZShHicN+EwRr7Y0
c6DYmN7fQPBCArofkCEDkgPe34gCVVPq6W8NfQx9gD1ilAfhf3IiMi2FQBSRpXSy
Ngzs2tkGrYUkkpKt/oP894rrSjJIxXlh1eHIqZ/mwtHpT4bltS4JE8ZvhJDXuE9I
Vq/8NkEll/ImlB/Xtd1mO3szD18OpU6CPorQmSNh+Ayx9018LYAw4XIWiHin5hhA
0h/pof8fx5Nyqjye2kAsmRgCQrLa3gQBpdb6bcyOM8t5YwHHKOZsd6UYQn5Kofsa
8PJsLBgmHZnTRuCwk1tqtIOXtiOx5kqtxeeCY9WFUH1PCuoxoo9oYKdHxN+Z9yha
n3kc/t94PrF0ZFZtNHa+TTqBGP5pkKwD1EkgJ7FgYokB9OOVoAYAJedojy13jPbQ
29iN3e1imDHRXUhh1r6Eqnpx9C51NVVv5tAiOUol6xG3YlK7PB/Pm7O/fgkxF5ao
48GeI6TE8BsWPNnvTF37XZp0WOqHUfxybyU67UO+Yp1/8NNv8jYGMLQl2F3IXPOK
Q9a+fiERkCBwKEQBlb/dccxrjsAs3d+hhIy9dJzfJUcN5mNFbK5KFekWevrdRxfg
Ix3YM+vm1B234lkdlP0ZVFF6WS3nuYFYplPswPVSBm5tao41XOlItI3fWbpuwAMc
6jhwoGcktWxMHqBu2/mvnspcGuyCwReUlYvZxTxbu8H5z/YzcNjY9TglyHmKQD3h
J1YKYR9r4RJDqfjrOLMLlm97GB2ehUnclHbrIaxg7kD3epRqfAj7wh3JdnA6bjTU
M9r0+hR3+LfN1uNIYbR/MAUw9VyvccSTtlCFn5fQR1jDKtTWdwSCjpGbH/+D/LYT
0gBJdulcFsJxzjhxS8JwqsbK7ZHSyxmTo84gBtJ5oZvnLgRF7BRQvkroMtoedVeo
SMQAm5VuhM7Bgwh096qe/EUUQowChCPvPbwWd65tNpnjfwF1jlCWYsGZM0WGNaRJ
q6GegpB3pSMVFlNPm8RVIuj0mf1sm07sRGaxOjo80WlCsbdPtJA9fGdg641Gr8SR
UnMuYP7Uw+XgCsiDZ5NUlh52SJnRvNFtmbx8lH86hlIpKSLauyZyEd1MNRJho/6l
90/5PdifSPHDzx+Lr9IZBPB7wfxf+pjh8Ie37b4RL5rQ7ad+J6Rk6ErmmhsXF3L5
fo2+F+6jdYNm56PW4Stev2k9JE6eUdwyP2nPdb/SVCDpt2fTbxngaRBVdEPPGpMF
uFVTdf/zWQtceQ2EkXm3vnmm64/yYfWc23EvfS1hq6yGjlJf2Ss7yPT5mUd8xK2b
mIsPrhGYmBEmzzaRwquKYpNT6ZD+2F25KQ9QZ1y7p16ZhmK6KAV7unun+Zuq0MDl
TjGw6sgJvLmqvyRZ6h9w3N2aGV10GMlE6DdRCSWr/iKod8kJUL02TLB9Ji8erIlF
xrToMmPr/sOLqdWfUJ3hgBnaQ+heEvmTxq0zbrWLMHFgY7a1VLVT3kcJ3ZuLBZxV
x3eOx1PFcXlxWXRzPsdr1vv6goXkCZ8Taz95nv8t+eDJ2a2S5tk9+HW1LByGMuXK
uCmrcU+EYw7S0bECnU+2lxU0q7Fj2LbNMKn+xFs/OMv1xjS1K0pZKwCbecSiKWzl
6oSFm3uQLzev3FQ97g0HQFBcsRGyzzitieeQcC+LPCmkoMx2YbP5jmidL3MBBKBn
Favk1osxyPhMCIafp+zHcNZNzP4oP/AJwpknmE/quzA/aBtKSx1wrWS1UEN+un6E
0y8e76P4+msYT/2DJE7xRORVW8/Xgl4Ec3dfZUfVBBkb2ia+5A9JTWabBhAOYDBe
1f7U6mvFq+FUdyI6xdgeFulGcP8xeCbzpBAUlFH+fDhvTKC3qxdDwyKxOPf2AQgA
BdKLb8x7QdY1cZfYQvKHPBVF9pzQd6gVDv2cJQzFqGxj3v7vOZ86tDwRLYqKXSFQ
bhJbP+tM+AepsaeqEeg0mgYGQA6k9SCueoWmJEsoGwIWaHoM5Nd2zKO7aS4s5myV
/mhZCBke73nm+Se0C2Sa7vjIlrcfcmGCUDo5getN+JMhdutK3r13k0+kxJV9ZzTa
yKNE4qN9A8Puyo8wx9sZgVc4lujcEhIq9IJu6FVgx5CGjh2fbQr7Z8agSwsi8qL6
MM8v6CDqksvcjkw3CY1gYpIlsgQPlEb1DROG6MRUEhSAjVtGyOcP39G2NRS9I60c
jbnMNKGfoSKoCBBpPXTSnP3e2vEuBZ2UxA/ERjXvUubupg3wg3GwkJwTfo0BrziS
9NCWVhDI6z26r+caWK7GKE2yrZXCZfKrICk+2lg7A/gyZa8SO8AQGFjmAybqPJzM
lvrfxukwTG5ogZcTTA4JQppXTcKDO0uF5Uc88sQExGV0qcspw7TxODzNQGdd3vRi
ywcbmvzR8UTZBspRPQj5BeuNcxkkipcrJY8lJ/hQlgCnrAR/F4Jvd2W2C1CkDW93
g+92J9wME/JxqnK36FDZd50cgPnf3DSl5DBAX6RuyK8ED7UHLznDvTDasqH1N4dM
FtnHA6/RuecwLA3tEkoXm+WgByVwjCJp1CnICWYJRGksVd19ixWoT3zEjzZ0pGnb
06mWJCZH1IwhZmiL/MvkAmUgRMlIJ+rHhKp4xD5v/oD16RhgxN1g1hjmnfq3ufcA
l+BnoeOD3nyfp1bcehAmR7QXSn9JUqgoCZBFcte9/JmA59y6AWVPUVnDphhRJHjT
KiO/t8guGB9CPMpSUWQRl8SmjgcRGNXaUIoEHMPRBFPVcB7dDFrSpbmAKhafglLO
KCK+YryzG2c2crmRv6ZqfjOSyKS8NemCno/o0lcfu4yh/tXpOh3SRyiZ4AGzxQgO
RrakZlwWSbrnBccn8McTxY73Jz4Vz/i9DxJN9iOQaSaJEHsuSXmkGms8lY0NSZxi
KL+zTVrkzmD393A3dDJF/1bVaADf75+sfRKxl4Ye1vJY3Hx8bjsPw30yvWSIbx/2
BX3v/Q/uGquKHUwPSelShYPetZwM8icYjvRLk9dRgP7Q64vb69xmWkGDFiASeX9v
E+H+qsxeukbgjgecE/v/UVPqeIyBYZb6zows8E4+9uJdWFP5QSf7dH8N6M0VLIA4
P6iRnamjR2UEO1Ss5+slFqIt6cb9gJM2FrBrxcc9EzCA04noJEojeFE1lY9jA/AX
bTnkeQMY/zsd8HmsUo5xKCAOAWo4kQrYst27Y1MdXoE7VBuplDwFK21/rq6aBAif
J2tDfDnll4AnYggI/w/qGhfSWCfbbqo1rsUw+sSZXJNf8n28MoEeWVbMPwwl78EI
1F6dBudrHSmTDb1Dv6PDdqcHeHfgmWQfBtDD7MH3Nk16Ny1z7+77qtS+dbwU4wao
mkRrZwETNO59zwrvXdj9V55z2KsqY7sU/gOMDUMSqZ982CQgZUNCtN7sfQWMSrGi
ge95IvJp9X9v/f/2SdbYtBq2FKzmLPXbzxdhHCkyZKIDHG8B+fWjpGu9enoagJb0
sxB1Ms0BEvFxpmkh3/cW9o9IalX4aU9Vfg1HsNMR1JWrIrc7cjRtIpeZeP7hgeQj
pWQYVoh4V2PorG0qlIjzjWZ+P6V/Sx3qDwwff8Tvs1lhp0d+k41+lg0MT2nVlbOg
PbO1rW76j50hpD5sjWLzA9BqzMtDi1+/mwCw/baPE/IdFoltEizg9YaDLNfOCCfQ
ze8L+Y18ltMR8fS21225Qbe3dLKzj9UCY5QHCDXPKbzylz4MgaSkZ6H5KyU5evZo
r0LdCNZGBqWAQU4TVJrhbZ91kYwC+u/VI2HdnNPbiin7HNko6k1BLZ37gHI+ELyk
98sKoZXFxQko+hQiF1328ZgntVLJKk0xB9rn2G15/y3OkRiSRr5/ivLlWKyzKn1d
/4XtEnR0hEZcG+usIgJOJ4lfEKpUJdckelvM6Nb/It7RCFRE0ggSCwhzdD6k7uQq
dIQBdXBczjz33no2LgMjkqWSJZopql+p6uroe8VYlKAkqBt1IE9cCxN2FTKU8Ycr
oJQD9HUhCK1lH4BV8pnsZfi+7v66N+9Q04xHCk6AtrCozMMK8hmqujNPrkyLw15o
9dYUq5eJO/zkuuuDHTNDeiuWZmAyWyZ3L5tOMUGOcgPkAmuRitP3x+ReRy6qm8Tw
epCf6fFFTFPnobPSd5lkaWY135/wbM4AsceFjTWabykq9WMCWvTZsk82KzJ47HZd
9UfBqziM8WpvoCU6NWqSlJAxizzvg9zNlN8RfJimBNg0AjkWtuCB9JDi8vI/fD+k
KS4VZdz1ex2LX+LOjVpmK4yafdbGJTV8/ppbqYvDFwR5r/epMSM2a39RKd3nvkHN
NUamvfJbhGaPVgAFWzuuoq8stUoek7s50WgtPrIMBjdq/fH4/pWAvBH/dgDHhk8f
bcDNS5+vExhKMCShH7uOZXdRW8oVrACAXzUE9q4HgDAwpdBwQnUZW8Puu2o3BHUW
jzcFBZ1lw0SHgJgvgNUkv6VpxIuRSb7+U+uTDs4kfMaKh+0PD0Y48vIJkgUaCgNf
HMTC6OFDTfB4fqWY1RLGk2MGj2UvdnVX66+xynT45OCTjjQedvyJpVu5Xg7Anfmy
qdf3DsVdKPqyXJWkOAXOudgnEm3/CDK4/hWm5u1QItxMsEYSVUkfbYS9wUCTpbNZ
MtCB+Y+MJrQs4IXXNJu/QXqaXGZvOdBGJRNi2j8w/9G4GnY+jF8c1qLpS8Rvhr0X
b1jcNRw6GEkf42F+fPROBFuox5qkWy46xOUHaYz6yk4kVn2TNxcZC5pf7xwz5F2O
vdDkgQi+uumLcS0fx1czcID13H/quXYdN0yE6Klbii2nnl3bD5TQHzLOoBK9ObaN
OSvvRFCVzGxuBnM1t0WpLjTmAFhEMIEH5k0zS7zQoju24fQ4IE5ptmo+AumIWUVJ
tmkXMLPxOwy00/au17mSKKTnguhDm92F0DksCVY32nKqozzzKNle1ElPwujsh2dK
SS4CkNbFNTY8WizT6Xs0cpUVq0aSsPyQ8o2Ht1SApNXRmT05TAvA/VD9DntdMoGm
6xYMjoyPJZ3ONbFFiRfWCgZbJPm1a6v/SxaOF/VjgclJJfK0RJCdIXExDb7djD53
WzIR9jtIDl7dhqWkYJM4JWKMOMQqgmgzWJec/tIpSrNNcC1uClRk4d53JTLg1qTF
S+9bYZCHACNmKlXvx8U6h6gBckcYiSdz7/MTCUu/ClcWWd5z6zOipUXu5QamSoBz
vNTii7yltRe9ZvyVTrwQ0SFX9e+G+dTApYLufGkzFfrKx2PMsIt81Ro8R6XF3sUq
cc7D3o5QJmKWk25G1meB/3E446cgbXlvMJDby8+g7xgPzrnADOExlsW0EvMh6jb3
7k9WHm5wms1U2AYfvGdimCaHFmrtMCG/Q7rHcQLsC6DRrZaSHwVCQBAtTmbuY7uQ
5rWGZWTxEWfxFy5fxafj2384ryao1ipvGT8Mvxv3Iq4VDKTPwuxoyFUAI0b36K0U
87zI48VJLSKjVrCx7iG4ntym93wPTFHfP85xbzM7+ejAEKsh/wijJRHXIp1jMJTE
kxdck9Sj5iDJPxybd6umOulVm8eVDb0aflOkPTVx8Ih8W42+HPRvrOIs7unDN18b
UaDVzNsnZ5BYey9UN9ePHf+drTxCkMsJxrAALM4dAyEOpvU8EQsMLT0ZsFnTTsYb
TuYkW9PWaMbLJpxSoJG8JVfb1sk5OgLrXNOHDJPUxi+//e7wBinEfn2/Y1gApoPL
pjtA5Zxtrn3OumKmvyAebdoVPRmSPzdT56RHKFhWqoOlDltnLOiCrXbY3BPAvaxT
sZEwUjB8Yz2S4YMaeZM5RIlqREc/0VB8CTfyS6aqfPIJHtOY99hhfvAsFpa1JRqr
xyDSzkiVq5VNimPxgVE8Z3A3xdhI8nA0+hkavZQ0YjDe3xpvdlvwVdtIAwY740Cd
E2IhRMnHlxu64xsBnOBjDDNf0n6CmD7RKg0A/LspZYQagBGedAjoP/GW2BBeIDDX
ou+SjX5a9vapziJ/Dxp5tnv72EmX0xnTeWWa00mVo46ApiCz8N8fFq+WHjhSHdJR
qS+p7nzApydV8KortAkvnKtrbtLPuyUWDcQarnXvNF3XJruXyBV6Ybemg4S5enQq
k0ru7y7AujxggQ0rl0t0pdbr9Y8Lv1t5ZsgSxvRHcQq5NpiQeEzfkkiPO+cAdcGs
K4lsYimqtIeGg0seFX0qvAzZsILbku+mmizY7PEBS7OxbJ/uAZU6TAkV0qi6YlqY
/RVFb1TtaGo1k9hsZjIpVHrOTPcWjhw05S3eDajGvY5lfdPD3k8Hjij9UIclQMxH
6EVLZgggoHfYZwzA+SbrXZ1fZxiS9pGQtvJ7evTvT6RjrPhJETAecoClmk435kEF
3b1krAx9+2nV9wts6bPCRPLaa2adIfLVDOwgu3IsysnRpvPI4+jova/YGoL4FkU8
eLDBW+2FNbXCj2x/FFMEegO8Owms/Ws9D2yB+aKbrQO+8OdTmxnYckMHGbSZPINv
zqKNZwljAbtZqvgPe+IJ9SqUUhXnEpDLuBZNfIGnzub9ZrC16R0ccnBkJjRmYUPb
271cob9EWxlbuBYfAevk4JVF2O2pEwpo4d/a9y3S1pIF+6TWi4jV3k64E5GBGKM2
xzrVVqdjoz6LKfmuHiouxfP/M47sMkvY9Tc2d/JEPZ3VRNkxoerTkNuK+rLHg78F
e4NNor9VjDVyfRnw3FbBdR4k06gqggqQs9H5jbxeE9Sve4sPr2QPEc96ZFIGWPiH
6sPAE/jhT6agUQLIfKrQm4sETq8jMUf289x+an3xptHcDPasltCpDPf4RBLbA/Xn
Ez0Llq+rWBAuP6o8+rVpPESSMfq98wTKkQrOJlI2hW+6TPs24TFrGQj6cc3soAWB
z7uilALAXa/Zb9Et+2ypn0UETGL4/M4C72YvbAnj7MfDcQb3HsRm/NlbNtCKFVm5
kpIqBLiyXtW7GhDcK9kAwUBigdb36zVVp6HX7MGgKFypX7+4ZqJMRDZ4eHQJRPMA
DJTdX2q9EOJYqSfz/PsrDwpv9qQP8TCCGSFu3KCVOJOEB4m5hq6Yfu6HBAI3oIje
o0vmqxpRzk6rRRYS+Mwz6cSty/zENaoBVMQpWaW2phuNTT9NgjPv/AVB0n8GNUpw
7tgLjcOC6kxxKvIWTS7nObQVBO8Z4b82ftdGTjU5aZskkTpSfXZwQT+BkrU5k4Xw
7+0AHRWy+BLcYSdN7udZT9QcH+VWj+Hc62vKc5JKGya/ZlYlW/pVos2//dDB+72H
85A0dNabDEOR/8rnQNE68e406RA2zaiwZdlihOozsaTfUDre5H5FPUoFTCS32yoN
3jOT1ODUPMDpTFXBpFfc/ciyRSqpH1MkLGUTCA9vmFhH64KS2Z3quJPZzQ34161Y
lEAX1TqvYB7o/ETu+T5kg/jKPXdNkhpzyW/aaP8TIefVuY/Zy36ppon0fGVCiyGR
z08i+22yw0rCWApo4XtvHMIS5IwkHGhsCXDV6gAfeMw6lpl9yyo23bX9/OIMZ9xK
jMmW40xTiF30A2qkC9LdClJBJFXKnMy7HUe2WY1Xz9mKIuH4z7d/nlq0X2e+pq/p
VkZWgi35KxWAckgDRdR+1h/sG01bpiMrVz6rdAz+FUKRrTIkVpiTeFwTLuJAx88t
Z/mDg3lby3Txl3pJX4IpC5hjDAWu8dEkQltcgVizsoNJ4j1Vlxx3S7MYm4S2yU48
XnwoiXKMgjSQfFCjAbiuwjai4KmfL1Kkmpx9PDeMymsCLBK0hflxsOkhYOY03J/c
QV+NhB040+Aa1c0/szeWR5+nWDIK0T7oCITE1RHhzalFRMvB91xF2CLZVJmBYfoq
v4W3LyqTW3s2k/fWcyVnXvxBkX0zUYcHAtFK0fCclh8lTNEbLP/INEfrc5YpMYI8
F/F5c9HzeyU3cbrSGZm6BGXL4EjtyXlGtBSqK9X5P2d2cWttecAas+pHMsMAUV2u
AVHxOIkdq/kLBNDQAX+/CIK041f19M9IMnDQ9S7qssMD9swXaaOJgJg7hZ+KC945
eE2LI3mA586kFukASGns8hHDN+E/9IIdBL4+NYIyWI4E6VcD7dtfPhCQfFiBaQp1
rADLhNk1nSvte3NuD0+DpNzaQLpQf7u7+kt25fNpyFP5g0ZpNEXRVM13As/VUAVc
jkkRiU4ew31KRzxbcVZBM8Iw1Q4GvR/OluCIVyFMzoXjRdeOEqOzNn+Wjwm3G/u8
RJfvCWrOxJS6eGetRwNhYzmvU6bOYhVz8/cnJVhzUHbKbukXsZctmLXVh0cSmtYU
KWLndCEv/V0+6tiUMEvsHR7+biDlmAe8jKm0lQlMijC2GSm7HurS5+w/F0ZfAE1o
BAozNmhOm8e6FYmjR5zoZ1kNKz6pYS8rPkjEhHxAAiVhck18mgRosTTcZeOj36dw
ltTGlAdSb9yXA6qfWGiuuCz2/YLP+KisEgHt0kzBURrVyb0T15tjvkCG++mjTEyK
Hix5V8ORl0V29wey8Emo4ioJB8ghTq6gjAfphcmi0Ba8ss+S+tbEI5hjawXRDYTZ
xEUrFlhotm7MMtrjch+Tqp2ZYbr+7ieRmPTd5fAdX6mF0e2HzG5OR4rP32hgqBa+
lKt7R6JPWUGl33ZvTm3Emq2BG7iCOAOTtrLfLyKHCTXJduCO9f3976f0+UYiikc1
frx9mnEtlRt+C6zUgE/DJ9jNtxmKUxeNGQIc+bttkwp5vM5T16k/U5eGx4Pa0eky
6AR4kAZ0F/4LeFDA7EnFFZ/vR9BL6l1H0lh5DKGvoeTkedZY+4mXCzNo95TB9w5p
rYFOUzAmkIcEVZ+Y2tsI/d8D669fMrQ96Rryjie5BLYBuUeYzuhJcIl89u12mNYt
A9V/d0toFzULMhAsvABF1gliGSr1kHLU4+R7IWVVbOhNOtubSeU5JtA34KYLm5eh
305n/xAyXDJSNEEx5p4cuM1Z7ODCtw9lRHAgVBTReBFWXGR7JaV5s7D3VLpRJy24
FX5zEU49PcjscGKM6Wtbge9SkG1qn3I0UZ8+fivUjXCGvHSRtlQ/hakYMileAg9C
p10AIW1IcXz/Haene9/XPLc3vkAB+y1wJihI8QD9ca9lkYITf0cZfBBx0H20gZ/s
Nl+dxPT/GTVTvzQLXXQys9OaKz37ChF4/cbBVzxr2XcqWU7I0llqd3UJXHYnKwyA
GDFMDZgdsOvKeXMweSWYzQHBCV4YgsNfkLT3TxnJDBTjCbLYIvmVnuqIo4sl3r6m
Miix8Dn0U5S4o8Z+au6dKD2XQW6FYDyC0S9GsW5fyFBTI/47+2tLa8lVUxmELSol
/OXPszSwo8qOpHDsrWeFLlNyfY8Pb4/5BKwYu5MDa6Hvv79uMVNPgAA1s+f1m8EJ
FAf/UYO4aVu4pEgAXp1npwh3diMo3mcTyv/7nhUI2EmXwDKSlHB/FjmFPZWzaKFY
W9kb77BB2jUHVFVrtuis+bqxcE51JSwPTUn8GJsJdwW30FGx2wCUl2QKc4JOHUKb
1AKdBNuQaWvowr2ndwluWvDsfwns2XBSE08xxlAThyfQPaahmNK6KddQnnEtoI8n
fLwmQDyAy4k0YJv1z9bl/N1/jogtlYogSOfqTbM+NqsV4l2IYwcgA5PzZrsJyT7c
3iWR8gzj75g4JxiLf8StQrh7V661w9E2nYYg0BctVwhAHlSEpOqFwR10nCPnhgGt
8UoZpAjT4ULdjP45Fdro9V2LP3vOr4ru4uAqnfOywZldzCNJh3nkCzXz0OWneDdI
sbOEmIcDg4U2V6RZkVDi43jKvH0wJFXXdakbNVj1nHCI40FAossfM2nmnL2dmlOF
Zw7WxKTKBG1u1ctLXoJ41dGACaE6vJZjuCwVrfjLOp4DhNCEPY3ON/XyrdQPDnUs
LoyT7+2+3t9NRpTpzHDjpdi5tJCX5WXL6Hwdm+iwIc8/TCptQuEhjmA+sq0hawWz
obclI6M+olTTioNmpdOlaGemoME4FoyWxGv2y+aeUlomeUgGggp5S3Op9tZvwvnN
1coPtF71iYtIywaETsgRIiMQ/eLLdRzakOow01Pn178/lU96ju6GFi9ZGiKLOJqU
yWhPkc3JhjGLK/u5qjbt3FGRhmpa318bLjZi8jNo5wsjbMEHigu8snqIGX2qIyvi
vFanGasxbQrJ3Ig3bENOFJsAxjlrp6PkKfs6plnGZ2HW8EUhIILOCx8fqi5mwYGr
es9Mw+NzFD+kHWIZWmDvrrpnRLFn1YOLEt4bUUr0Z2jrqhN60SbqSSZ7DGHoJ6Xg
3jLjznD3m47kdIip5gQDDZ8kpIk2zCam0kqgcqd8r6L9AsS/HcmYUynbBH0LUBNW
zEH2L2Dv2/3CXoldJ/rbogQrNbBRlnCveZIXYAzRwenPOmfSMJaitCoW2OC1y3IV
ju95c3ZsLt9h6aXA6pqMYSiKzDa9nZ1RXPH0bkuqS20tibA+JzEHyRTkrQwHzo5K
7pF0Egc2bKSiIitvYZKJrnq2N7W935raLOo3ZOzTUr5i5H/E9C1U0PgH18WaPSSw
3Q16z30JFBvfufk+sqPwtHiYxZA33hwb9TcjNY+RvZxWEz2ruE+njZbBQuAgC/uq
6UWlmQQCnIODJ6lN/gPxd58b7FZY+yIUOXsRjIpS7Z8iYFRkWqu/n2jNa/ChuewH
3FW7g+DtNXw0e6G/ddYvsFxxH/iTOTJf7fMwgQZ7ktWuMvx9evs8agaIj4QToDVj
sq+JeFjK8b+SO6WB7KLrzezQ7vIUi7lV2UtAUNiCguGPGJKF2kyS7qVIGNm8fBaF
INSxwHYSTpJhvRm8j7M2gzOYdpomKVwaUOAg1f8pIfII0mlbIc+on93EyUGBrs/x
ESeJoGOnlIbuYwL4r9KflzwwKmwahtSoeKjroewoaW5nccHwHXzIFn9HisEySyUr
7M9tPY+7jXcB5y3TZJ/7rozaJR3bs32YGaxS5WCOK/foH7JXwVQe91pD1xilmwsX
OFifD1mCTiJl0JfiN+1i+UrgjXyO8DUwEAmD+H7xZs3WpDEyKXpDxz35uzSV+FK4
i1/IpiIoQ5s0fM3/wFbyGiT03DVRX4IL6jqJ15QQeLhXsr3sMC/5NzUaTwLjjbpb
xyIsLhRPvvh72vhWNzGdJlttLlnb3O/wBGsM16TzIuKqK+mD4k9EkD579TV4oY6Q
VzshYS4C6zwTPcSUDWhGX3OqtPsr9eR/PVzitAoNtF6HcqNG4j+4t36hoaKSGDHy
w3BKxAPFYur/k6LfP7JyaM3zgVPqrl4OP1vERn8bYzKcRPpYfdfZ5MI/DThJMhJM
Y4UYgInjHFlntvJ3ii5CbFh5tqIk+VkpgpqUc4Ajp/FskXYNIw83GXZZOMBVdwnM
9LDuCZUkjlGG51M9HRSDvauK68Rsn1im1BF8opTGNKT0wgm/AzKzWTJ1IqCDkd2d
w23XhAp5PG32ugaD6zVyn0DYCdHRkRzNfGWlk/w4Y4Ni2a7Hx1g7Iw5coRoVTjuQ
P5DIME5N2xcftKcW5rESWgeawOSd5px9/iPIih3IcSF2f0K719TEarRsZXdlnjw5
PFm6x+B8P5K1nSgq+vY0O6DXUjgKC1Y3iAH7miWLWgdZx+snAK9TP4Enpo1ZJYvL
axNbsHcxkbEGGipfBOpZF40GWtKTR/Axx+4WQTAl2ts3TQ1+CRdFYP8CvONXF4i1
zZYox5+58LMGZ4gdaZp9dw5gkTQwZP4yWIn2O1tAMChHRAWVEoz+0n9q/cbPbe23
kY9Xz+YhVmPo7XDIl7QuR+LSH2Fb+lO/+XfndKae/sUPRm6zwfSpFnl3DsLPPX0f
/GPRYhk62ATU+9V/IqpfIseusRb6IkLCAeMHRpCHEaG7ofZGs2yIpk18vTrSD2YY
qYGEfImXSEueTb+QZa5lxEyhYnwUKJXNuOkrp6kRGsfxQGNOAv0CUptrvkLKkEOu
1Rj01WUMsO5DbRUxobmEuk7G2H9cV0qKcGiEajuyqEMpDmy/Bi/jLEj6CT7mCIcA
YtNJXpwiMq2qSLNMRznQI345QAxrELDN6C7mzlnGQ/edQ2P+ebz7BtR6cOL9MmR/
n4WeAD7KggOHmd4/L9x/xJJWWLdMdtbyIpOf81XQBtuE9sfRrdBxYePZHr9cNL+y
KT8cbirjRzYOOnD2AMoLVjMr4rZKKYl+KFcLmKr2o5y+pwRxxmPFgQEy94dXiLqt
YG48Ku6pE/xhKcDHyrENRjmFKDomh5O9di8t7IYRRv/w8+lhafKGdtijFulCM6wa
074RfW3D2eGHii7y5fnvYqFXB6YptZyg6WhRUZE1e/7lFpbQQDwGXDuHRGLdG0Gn
DAAFZNcoD/Js7NyfxZjzJH+Jf4JSYKDQ5CvAUakOizbiOwlafhNuxIheIYWqAuk6
5Yd1kC2lRXuaNVVkGabQex0QPP6YPKaVtgJD2zLFY4l1DFIkXX56FhqFOmOZWmX/
NlBqasJtmZ4ScZp/vq7m6bpv+5B48Zb5pFKsg9nhIGL0aOn28ays5NZtAoS3xBQD
wpZvJKaYQw0iKwpn1JqasSxai5G4xemZbo0a6Dr6dtKiB8rbjEGOWSA/imvWrf64
F17Lt7XOkXlhxk1hPxRyVE0C3Ar+ZOt4fSStL7kgXQwjqdzUxax7RFFs22NEsAkv
5w4jH+yadNFEmp2LGW6l6vQnXcjrNve1VdMLK+bMTD6PEph9N/y3VGEvoBK+GbIC
QkwnyJlfk1HJ7ZPyazD6UWhiaap8h4S9mhof4NjhaRPDGKPyxZPPXFMqsi8TkJV0
s2+xGW92DRvE6yIsGlcwLWllDfh1O93emqWzHUprpgLLpi9+ceau5KSDha21M7xj
DaPZLcvtuPavl1xgkTaQAAWlvqANg11axZ8Yg5rb6XGcBhqBf91heNlYNtUxBwI3
R8RfmybRakiLMIdS/H4NGCbhh3LVZzBI6fVMav8hWHbEHBUUVD9FvmPPFudXKbE7
kVWyXREawIW2rMcFC1zBG0xziYdCYce351KBbtIGXoEeqK8W+2ERRuL7bbRl7wFZ
G9LwOoTm1CdrVwaHojtkZQhJCNqHnB1b4rr5zyLfCq6xkD0Vhkm4NL8YagUeb1pR
ko/g/3PrxxpWa/k2jgD1vAkprnLB5gQykzAV8tLQardokT0HWynPTGKksVliICex
wlBs2N7ySmFA4ThH1Ddc+auPf4kn2NFL/ZQ7SC7r/mGxdW2zBEJD2gZMpwmHP9j1
1lws728lwZ0F8JDn7C2/skU+suJriNlUsb7+M9hzYODa8UljrJLyNNxS9APr6wAJ
HN7dImw7wBtQN+48GZpTBjFukAtz8cmzTh5p7z0aEy1rugXLEA1o2Fgz/nnk5QiG
P34ynjlJ59EuAKwRo/FdevUQllzi/nl/Q4IA6Td5NYgmNG2r2axkPvBr7kmoe1mc
AsaPioIxIkRTD1I5lyhKg6QGIT+0DTsBv04VTXqTq8nGQFIt4VgmuVOMji8p/qm2
NnHk7G6eh3D9/BlXQ0uPv8KR/be4kAWsjNzZ5oEWe3MCmqCZMTDvbo7IjtV0zoSY
bVOV34xIo6j1fTVgYpB8ypACjKyBhWhSMeB5AiKXoTS/z8fNSq+bnlYYbNsxX8Ja
m1thz6I9N7zpH7LV8K0lpIVVyC4ycyC4ygs4cQrwt6dqYIKzGM6oqLe3vWLpruDl
xweI2+b6mxmzX5uS7QD4gJiz3pdS9S8dWkmcb0LVfNKg5X3SDz02TE6ovmgAEh7O
rjstLQ3or3v7cz7YfqLzPhy9p9tM+PRUUE852Pk0M/7aGnaWAR+YuUybnp0XvQCU
mDqa8IuWQUofkx2e0iEbOsZNviS5GYRrTJaY0UL8VNHLOrlbplNHgKXyV5ONdxwY
9j0V5ZH/6QE2NfcDWAmmrI7AVO73VG34riUiok28lj8of1CDwCcStOKSu9B/ozi5
QdKnrQ5ykxgpa1FcEXAhttdUbnbAJAuR/Ytim6XHm0Ld3Fs9fejjlfHcwqmeYdQi
fEBt+OOpPtZ5WipGbflPcHxQj86Nm76b5f71G2bIc6bgZaZeLdLvd+syoOEE4Mu4
zauHXrcEnHcHHgY2T5WVRZvMJ5erJNXMVCVPZLNnYEBcQauZL2MifH27zLdxQ8hI
cHf2OVcK/+uYGaSA+yqWArUOqC923zzwIHZ7gEijONS2Un9hvmjL+AtP6SjYK7aJ
iQ2aa2xcuQI1JXput5GfQ0EojNhvAVT/A+u1qYGoElD8BxEJiLRz6bevR/7wH88T
yEd3WQE/KgIDanxhenmF1662lMVnmPMQxSpKlEMWvIaqs6a1nb8DX42oXf16bTWx
oeYxx2DtJSYXKQJoMqCtZTKGQezwEMc25XHaWVjzbIKeqOgItdlI2B4lgtrO5YLO
6IV/ncL5vpFtm66PjhCTN5qDc3d6OYYgUZaEcE4mk4cbegfbfNGCoFjUGQ6xPPNl
BzZDefGYY7nWK5rFoWyuet/9vPLJyGj2l/Tab7pHigvIvAjpyt7RFWRF91NTZ1/B
hn+ILAARp/NM3lPNckwYAzHJEMnwoDwyH+PHX624v5cuUQKu91IElfoFeE0m31XB
kXLBt34YZqRJAJW8v5FehPUxFqvVsJYaHam31NlfvStQtnIxNpY22FFNxJSllnnU
WLFRFW1B6mEuY4mJOXZrEAr6KFn300TT8U9XzglicU+Be/L5wFfbYFlwXT1FuOR4
YBVw7JrhOs76UWx6JtpOFsauDjbQTZ79V3gWXK4NLFxnMVqBgaAKFu6/6RNMf4OS
C9Lbh/xSictSb8tn99evsS8gis0QaNh4Aj7vqxz5M7HGmlrruTpK3Rvlb7r87t/x
vy1QkzT12NeFiyGz3RL5Ok99EHdi1Ubu1P2MZRk+PCawNqtBcusk+7ICqQg3AgFL
PCAaPjHqPIrej/oiBPxHUiCG5df4s2Eu67MV0b+RqDDjvtutYhPgUkq7pVwkniwe
wGJ9+AAI4Pn9CtqXIRx+Wwfok+vkYCtMwSzjC8jj/TR+DTefPKOn8ikSGBoc3dPf
pflvfzAGcs69BO8QycFgVw5Z1T+Nh/HKJtTHO10BnZJ6P266X1DUUqrY7mm9uZxH
f95c03hXUFVBXMK2CvPsD39XA2L9oH0lTdW40LT6ZfMyNUYbg0UDDXQBsVobExCn
Y2RNLC1jVOj9DMQSIRtTuPsP6/V87Gyn+S6r5qoQJNYztDATntUZU3Fkb+mRJFME
MkFEExX1mmWuGmes6KrDdL5B5mHzxmKj4BoCylQpUUUFS3nIv3NqDsqxsmhgOuMN
aoHKnc+bdzBWi/Ob0J5Dd1bLlwsOBjLkg88VW8EB1zqfThuLGdUDePivBe7WG/ZR
X1U9bajGz5d2paG9KqEWDVA5M1v3fiJX37TjeNsHIkxDTlx6RkEI7lbjYp75/yPr
pLnp7wdB5sfkMmDwad/zBg061fULDzhHLGrpJrjtlxCHVa/QgBTBI0YYnxmgW5jG
X6xC+yWaSKNErWxU0NyYsFVQanD6SIVG0w+kEysemozVKbzHGlevK6cOJ7su+wSy
91Sxn+XtWE7dmiAtap7yDpHq8FVOg+m653BaX3TflzJ+wjWpOXuVIgYarFUDXtfQ
O3oOuev+jewTbnBvZpM/eOZLJ9N/h3usyFjVzsU4Gd8nPDbQXC2IDb26DP3U59pu
iJGo3UxBV7X1a7uickjv2BG5Kb+ywekbuOSImIYoEhoSdDn4YLseNCTuMn+rKjfd
zGpNDUbWTws9LTGc3DsquWJsijx/nsE7AlJ41Zg9G4F1F5uRcwGicvRt7Euj6b+h
W2W8eUlJ21tvcra8BGxncmiD/roX0zM1Izi1SsguGu2IfiP4wteLWdkuxbdpgxRs
ATuifFJ6tKy02r2GpVvLgteub7q0BWk99WGPjjNxpbMYTe5abOtr645QR0lJGWoY
09QE49tM7l7f4zT6i43Xu1uIixHfdiqvi6DIjdeSmKQG8Zmfeq7C5dgsZHQ489DD
HCwZ+KiSOyLO3/nBEI5Oot7e3GjEbTXv5IH6tUUUoSF1ew0PkpafKW7u2L3momJy
PpR010hzIwNvA+kzNyCYfg1cpJh6uKQOfNM7gPZhpU547BbTwQobfZiN53qiVA0k
UEwaTlEOkgKYuvdkjcePxFNlI2DvlVotQkiCpExuFDyzs0qUbwyw+B656g4j8Diq
JDV4JlMCal+h6u7Q7d3ij0Sy5y6ZQkfLY3Eo26ggODw3dOxFhQSxm+nFpjyoXtRW
7OAZwOwMSeI+WGpDO3iAmlVmg4cniBHUcz2Tlvbqa1+mhTwltPlVBmnmuE4rgfiT
BRl83ePIkjbM4xBxfG3JHiNIRSvhRpV77dp0LZE0RMA2EqcfrRl/BpQtVJRaEZ8Y
oNU1O8sGFLqCO2sihBGHSYO2q70ueUpseldqucWfcUF3j6wD17O4kcqLlQXKv3d7
4GC7AIJ4YgeC+hk4Ae8Kw/yr0j1/HtQGNZkeIQM5NvBZWg2aIc9Oz4NJt1+tChwc
Jk71ILU9mvmqeFy4DJKQl9SHquP/S+Bn6Z4PCNnrV5adljNmTxvvwdN/iSFye5Bv
nqiOZAqI4DyPtor44b7ewIA2OXqNSe0Dme1lJt0LOiujduLh9pr+udneLvR/x626
IEMZW3fyISP8+atnrZyMwvZeuej351UW3kFHFX6Of6Y7c7ksvySFHzAoRHW73/9q
JbHfjgnYMqxN1OKzmyLhqmSlgAVGbTHhOiGD24k0/qK0hoynr3dLRJKCbkWYljPI
B5ExyGlXyq2Ft+Qgcy+Wa4/IDkNNLSdcCm0Kdu1PVq3AKB6z1l+dEbuNEXYxwVp8
W00bWAXXTfgqx38vrKbe9vXC5uoS0FluCUn4xizkvVK93S+6MXfX+oIQ52FwDV1I
FSGg02bvVZlaqJUz/0defUhUVg5rQb2NLJby2Qb88slECz/gM/q6zfJi8n1pRp9n
R50GDq8bxmtdnNm8fklaTziVcd9jbSiwGMpVaoTuO/vx4RIMdLU9qsalL3aWTHSE
gsfqrVWsBfZ2mOYbfPw58y3OawLxdDSt75srlwzNOaS0gw23Oi/9hD2SMXx0GjPm
8M9C+knxldnqSkfx+GsbstdidTryKLR1/7O7+mLk7LJdtyXOZj62ElBE4AsWyBlm
wFWafo6ko698zybEDRExTQjUuehswkRQ14kg0gnJ+Bf7RDfHEoD1utEOnAa2pUrs
Zvcx4SruCNUhyyagR7Jb2EnmYRAH0o18cWgwqe9BjehRE1PD+2SyRYSfbwf/GLNu
jQ20FNY/9lVcn7I6xg4VNg23id5gxeufb6hBEaP5UNAMoqM2oyvtfe/peX1wtK9a
mPoscLacTkddPZVhoftto1GYVRAXXLTP3+Sqdsi7A0KHidGWnVY0TrfbS6FIXTK9
pJvNoi6sZ/x2nkwDxJYz5hSFtdoFDeYmatrOnt7TmY1l0s7h3IItn9KijByXktVr
FsMvg01nM/d6jullSRo0mESVh8GG4Ox2ZukPeaCxtsWM4laRcB27pWh/Y7YCZSM/
MAH69Yol21ATOd2kfQq5J8NIuQBmknyesYFKnqGkXMRz+4U8ij7hR5g7czSjL9Vr
m7+U1Y26UyuMWax/0u1dUVFIO0EBxd+sASjjlc+Cldcat4gOtYcqy4lh6YIpDbTX
nXSb01UucnHbBqG8e/5eHwfPp0dfNER5tIbLsZQ+kDRY3pIicEuREE/gDx2J3ETq
TgkdE583yfQNx7CT9ioVHZUpyZU8tVnhVydkcx5Tjn8rZHw8MYYQVHOJWUktcidL
UHa0uK37fJ3Yk5lDB9blyXE3BJljr5Y8dNnxUxcG/uHb2DoR7/e1AOYqWDigZpfF
NfZ3qMP6sSv1JocnZs1b0qTyR0/lF8UbDbCmFBn2knsgXyaXmDfSSyJDlWB4pwsb
8x/YtxmLKoKn4ayjteMtbJIpFm83bUCvoQ1+2bnP74G8jKxY02lgz96w3eM4pa/u
8FyNDJJ7herXYpmMJlAXV4xIFTrWZWQe4e3stOWJfm41qm//fKypnveCTtkWC0cV
SvgFXdxeLEYD4GmHH/uObZJPK1MT1gYHN7xdWsmUzKRIpXlk3SzvpdtIV6mNT8Z9
RPLySkKFgrpwo9eV4z6fpoJzY/f7HfcNR/NveD7xz9qUqCd9FuJdlUEaw2WHRAaX
SBX8dnrPFPF4/pZgIwdrRhewl/cmx6yanEZ5f2D1dcBUVwEEfVytgvdB9Uqe8gX4
bPF0bfxA7rFA+XnPiMEfYTrAb0B6VFFNCkc/2n1Bj65ORaTx5Sh5DOvFqbSeU5ls
nuXw92z2NLqEOsfjNWCZVfvaAaR3w5q+axpexplNqA3tcQaWVi92wxA7A0wDx51c
xfuNtfY7eUEsT9aRMoLGRBkiMUcirjdFRcmBFXuDRChXpI0Ghpf6QynXEJVuqsHm
HRBwPuIWT0iVg8ONCDoKJTFTCR8g0GFzSugvnyeO7Ph9rSG0kYMkk6rKI8ZiC+vi
RKdTkL4ZIvBMLdpjK2lx0fcqb7RMJDW77n6Bo5BPhuR1oNZi6R3qMxvb6BQEpUu2
ZYaUyxgRt2vg3KKS1ljp8y/CfskrX6sg9Sszb4a+ewmjYCR1sKWGEyIH6Ssl+O6P
RZJbjXuux5jJfsuuc/FB91vE7F+KTeq9f/4wWxxTMA2SyaH5YOeV3fVG5Fy7V7VF
gQziijFAlUYP2psfcK1vj26wkkrVb0PgsyCipLZwNtm5BnVpHH+TIR5jmjPgm3br
6NiUf+2cX4R7NNxrupZpJbFIHhR4Wv2qT80nSVJus23kTuCqkii/FWfwqLG/6BzD
kbH+8DlD5ftX3DLZQIsGKLg0CUAfkG14vm1cmBeTRfNnW3XwDQMjbKIdQ4C8GhtK
htJYc5NAWKxJKhWbmGG1anVnKumAY1YNTv2V7h1f6+L/jn/Pa028XMJi4zJWaxca
vUdZFie4f6fpaEWWhpQG9KvWqvXiq8XOfRmAEXUVoACEm8rQxb/K6rVuaiHi5E0r
R1XRHGQi1p4UwtByykTI6RBFz3ElSuHU+b11bw+NeiqAGA8496LteDiJU64l62jf
hUGVJDBjxjihZ4uB3wjQcE2M5N5VhKscv5P9VvSClg5+h4PzS5p/gHQ7j1THUzwH
LAtu0rjuvT67qk/pdjXZ2Ux8BeVZCf52FpZtS8KhavoeIkjrzUqKTqhnm0YukqPJ
WehCqmft3Yb75Vl8UlN3MN7SQlepsdJOo6OT27Sh7BBvIPYgTgLMnDuWEo8BOr3o
mV0PiXDG57kuQluvX15l2vkxWbyem4qx1e+plLvzY2JVRIgYt28RD+qNrPbjSFc6
TiEAgs5uU8e27Pj28V+ZvUalkq48a2fmkWbIZoTfW9j5odZ8mqSl6TRWkHXXToKE
GSeX3jr9wM0K4UWZR2yyYk9Om5eV0MaOwF0cPYiwABWzrWsg6EMhN/N3PVhC4Qvp
GyRs7BbntnMSOppOZ6EVMLPn5MOihHoigCcTgLZJMh0yqoaqHQfMhp3OrOMGUjjv
xCYXP23h+orBChkiioHtW2C4phk4yzg7jT97Et1/U+vmeVsECNYgB/vKQgrLoZBq
+d2DbyufiJ8GjLcV5eSFdo0ZjA++vj9vRe/bPB7mcbyKipKZFr6y7rnpuuS5zjg+
SeSeQMVBxD2rpi1mY6R2SoPjGXJStgpNlKllJcCWARhbw8O20SfEJFpmdRWC9LbH
EXtDcwDLAKXroQgHB8GlCkVftcaQ1VImaUO42YlSWwOfuwsyruM4wB6ZuQVMdFXC
FJIxO2db+vrbRgeVlOfqXs5IkNws6aimMFHe46ow1kr4h+UTKjfEDg6ps2hIZY/p
NoQJFDjHA7IRmu8eR77VfV2cmYhWdr4ztwk4Nce3cP+54wQPrTHHnnFvrNiNuv2c
sdunv5gJA+WpbqFniDRN9KgyjOKM/QoHm6xPtXTJrsTj5ABnbVocNKygoBJ1ERoO
YwjwTiV7xVRoRve4e6+3+cnhB2xhSuHrf6HtDwTbVQKYD+SeipriIAZRRDbDxRYg
oRr44Ka4lQARiBUcMheBsN9eDJ95EcJM8RfWPicR8Xfi5Kuq9wEgat2JgJBIO359
k5Eh/kvD/mGQLDbbbRJ0KOE1OfFVL4LFLAb3FgYdyNXS++YjBLj13EmaS0vGU8gr
fTJtTtxjmdbKEyxBZisYoZeT4W2PWJwcMUulczthCF+QvWSnxzovJrgwTGoIbzk9
9QRrhrjz0sjWuSPDiE91D6av6POZKvPaW6MrBEzG7LGDfxC56pvofvRrshdU+fYv
SbKDiUPwcHp5SVBNcsP22g1oEeIKd4DpnyaOeWeB1RxM/g3cPYQGTyKdMEW9hqC7
Qsc0EeP/yujc0/tuZusH4wvzjOt+wo5bHKVcMyeInnkobe6nm523mwTy5UgVEhny
nasMj7Zgj64aHPnzk8SYG1nR7rjBs5w3gHrBcnCWQuXByWR9FSmN/x5GHJzeXvyp
T5TifKEToaK5uTViNSGRNhEKpcYQs+GrnJD3zKHKfz1PIIwz8+NYWJIAaBPOoYA4
KyqDcmf+5UY7wngGqhyKYsUdQZkAu6oY9hQh4EdY/FbvG+tMt3PaJhNsTPyDNw0s
d6ySou4/P/FcM5WmHskomyGBs5vchN1CGeYgAVZ4+OkHIahTgEeklbe7Cu551K8X
O1kv2K6AB8+IgesiyYrfkyDFC3WtpRLOqZprcs+NQuOEg6YwtwThfIwiDgrYYfPs
ecFs4PHlNOW7X6AXyVz7MR+IxfZqfJDl57rvrujbZE6MLujhdIkdnMwYPbfO1q0L
+hm8hA42RrRUaZ6CHoViFw7w4KoCLC1eBOfPW6wrlSPSMdj3U+kouYTgRYQmbx56
sFFXUaSzUNxZvp6PPzD3Ip2QI9+LZngmcPPlK8SF7jesI6AA27kBADNLcj3CV44D
wt73bqNT5kuJD6ZABoyTdRX0iYGcuhcaF4WaICEZ0m3QGtyO4FDYjhTodewI8Qza
lZPtu6+6nxQ0RyO2lM4NrtO3CrA1skR1/tmuVaOsuQgDt+QDjxsHX3MEuOLYi7f7
YUOuMAAzaA+XjoTERzbEz1Mh+G1xij8NW/veEcDWmzwRayhjqzY8eEJKzH51g9dj
1irI9u2tCY5jxm/m0cV3cJVHoH3B08cMvSkMv6t+aNfpBefVzjr51veU/4AePsrY
fAaOQpDFJJpx/TSLSCo6MP1Uf4guM9guyLnmUVt7PBNYquc3gTI9J043Wq/j5Nke
NfyiLETV4QJPeOuWHdgHPxrAYBnXoAeEO8uDbdJuvrwMAnU80Wy7EgFalc/dnPu5
KX0uIyuJUzNiWqSXt5dQztwg7m3oaVjv12gak19lbVQ9YFWHhbG2Hf7QWj1PHn6S
b4qBMfZKk/7dfnYIMns1Rou35A7wwhjLuiXJ/3k2b0kyfLmkw1FW661i1bL/6UYc
r5bfe+mNWefOo29ywXESlRcDolLWbE8FYW8Y6qbs1wE9UG1ETOuhj757rEaCDd7L
qLAdpYEUH0CEkQv0nn0A0z/KG/bwaZ5FpK6dST8Viyt5//3uOzpyrM/vZKW31cke
CMpr78ZgvDvTGZX29l59sE/MHgNF5y/umMHYnkHoBx9txJ3aVZwev33v4yysifOe
STu5+C42YvJDNL3xa7N4m64nBUSJxz9ub/gc5kyFhnnrcOq84YgB1j9Yvw2HLppO
ddWJt9imeO2KnQIptejxDT8VsXcm/6W5BWWsaDbMXHxfRHozYsNTPx4rhBgUfBgj
Upk7ZLVhPniwz9sKuOPSc6MIj0Eo19uStlOPYUVipip7rn9RHGhmPWIE9avhGtj5
xdKcq9JDh43Hvq1FgBQojSjaGfGCaHSTQA74GBTBUCNzcjaY2Z0SAnsQIQvkN6R1
OItP0sR4Wnxh6jgOLwvhv+Zl8ZBztCdz4kkSdf45rCFy4iCqrWXvOl/6TQTw3MxS
l1RFceDTqc/HC8yagdCNRxM0K3ytOk4mA8XB3PxgICTQwbCiQJ1rElbtn8OADpPj
KH0h/hpYUWcGvKxCKILNGGRI+YBQ7AHDOJwWal6WV4TsljRtmRqGs/J+8SnEm2tR
zCbJOJhKjDZyoWpes9PNtIsN0gS8DPmfqDoMe66dqytM+2D+5ErRvLBQelCLZN1z
thnZLFzKI8EqHKrl4z7AsJzKvo30ZEIJm4eK8B8CaYVvmWZVrVDgxhz8HLzaQmGH
tFXV+ekSZ7zUNQTDBef/mKDGpsYIU/KBrX/8z7fcCAzbqBBie5Q5dl+EnrmF4Nh3
9IsZJGnCWBd8gnp+a2h8nbVgqAUYEz4L5v+H84vylmgBOWdo7YlJiLWVO9Vg29PB
Zj0SdM7yB1luaEcS1tOePU5luBIYRS5I6AHkIJvFgt8+33zPcyT2us2Soe+FxQeO
9gQDNHi7SibB9H8B4bgPTcS4MkWIZ+xjP80bt8g42KjEjjnavysXBmzqQdo+xUix
dOPENV2H42T3mmQGLSxQggSztznLXWk0PIzt0UZ9AhANnpCio87se7Tlapgw0cAY
/rtrl30rCbMKeA1r6ulORYwvixe0vjnM0TSa6THfq9XQzYuLx77SfGvGiaOPvGDn
C3rgOh7u/5W/ffP59gCVCMeZB0wixSBrnR+vAzrVfVRiOkbx69QpZgmmCScaJLUB
6B1fcGTb6H2jE5tR1xHjajv9z8UU3I/L1UIl90ehG6gGvsdhsQ7h904jdHjciMRP
UUs69Sp4tr/31V2hkDLjowWHuKlPdE/0f2EO/ufG5vDHmCvjKPouDvWsY8gRFhlf
yhhyYP1rKCmmlNbohQk6Hcp7pBJsKplUnBmLoQ74hEvTHGpcZkKRzh5FZoU4/atq
d1+o6XekL5Qsd5f5WPcVFarg16kttWxFkS2ZuxtzIBMAQm4Y8xf63rvRMT8XukVr
rfo9GSyHX03hcZ5v3g03vkfZbsfKF45wWwI967a3zwT6RSyuoVsi1yQqEc0B5yhE
MKOAo6PCtwnRAGTWFCeOlq9fQEsEc0dWKzcBm2bz5F50nOEJu1DzL9Rf+rzwN8yD
YqRiWwov7bNZFeEq++WpRqejYTn169BMh/6TDNSk5fq1taJ74Sc7hhqsCODUwp7o
XABvVTixteVAOKLruxNNQDQSzW9+reU4xrnHP0yQLFKOXVQY/SyW9byCvmaTTsW+
1l+CqK0TwtlU/1DzmpiUh4aKBT/Nmk95KQfj05ztEfwNlySAtwa2Y9sJWRObBdL8
iNEPfL+dUX3PD6CEEwPIS4pnGaMz1qGKLlOj24qviHsDAfVHRBiXgxjdvf697FtG
5l9KjlervcdwXtE0xaet+vfrCaObIJaXf8DPsCqsZkw5H1AlDSbZtoER6CF+e/tm
IUAs3pHDV7ELz/lumwS+zwcG3T7e4oDCktYyqvZmiBYrcbgb6+qMAKrRhKaaqAEr
BSQy3+/AsspAj3vqXuyJCKqM1SB/6LajdFevI2Gz3uvcBO/UV8O5jd9D6s/JlC7A
mLQIJ7FnPo/L0/uCRe7geo6fmitznRkvC/YkV9D/QdKIC/gD2J2D3pYs1KXTm75L
/5BtpCQboVxyqqYed87+oHe6fAR/ELPjvEmnnchbpXeDk+ki6cTlho5URDyY6axh
mTz4EO9t3sV8ZLaz+w5BNnjA6vVe3x/oeGdNlzcDrbLJ7cb2LpnzVJbLAiTrGCP7
+hhmQ1QayLAczZR42CvCx3R3z1QmNpFIK/IjZDiD19F9g9b/ac4gf727/dlI6G1a
aKotv5PIYZh6ucf64m9rNlunnKsJXZlUSzAludf3kl76sehOMAUpeZMYOJV4BeAZ
WmGrYSj70B8z9bR4y30Xw/VbLNQcF3WzFuIA//RqbF+IH+L278TL69Bf/5WDu0Ow
4xQc47XoC3dinlOgy2jhFssxMuu4h6YKqR3caW9wpB1iCd1fCpvQ8C/N/r9Lh1tl
kulynXoDwY5M913p6SmsoQFyoOkPJhwLkpovyYArblJp4yxMSpJLEN0xgWEB1YED
sMPEIzABHDCE/LCoKCYXui6fCC18iqq/I/2pAdxDspRxoTK69bs1KK5FphLAORDJ
DMFi3PlPjEOXnbJa+97SObeDln7b0sNfStzyfmNb8/1pQupGEUuvjF8ka+JJXwrD
2XYYD8zGxaf7qQYGQhpKTG43gx3D1mxyGRIDL8nODmqrxWICctJqVcd0so+Z/AZH
iGYRWFOF0bEow0WrSb3ZhzOTIWNHcmoaLYr9DFiWL6v/z/k9CDVLT1f4mYJGtVc/
PA2GVeiRuNSf+RYb/Zy7JGl/+2CwpxoayYRDYxgZiQCrtQlybXGFqGi6Uk+gR2SL
PzvvzeaCdR/cgU1TB+fR9x6mseTZgsZl/LirCNWxLpAoDw4ABhuZ8G550YFrSCL7
lXMjtD25ZF8VxIZGlklEow==
//pragma protect end_data_block
//pragma protect digest_block
HOq/C8tMxNV5iOAjIfrNwCYCVmc=
//pragma protect end_digest_block
//pragma protect end_protected
