`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
J6s2YXU3DFkAR4CkIQdAjxnU0oroTi8EbVY/3FjRFTQksLztugCR0+oTqC+0iAFC
VM7C+hLVbjDjfOb2cgC8hSI+5u6TvV3VFxIEzoQVP7i+igLsOXyLU7NJawDMWfVx
3hKOzCnEqYKmJpJ/PO9yai0AP8IPNUBdLZTObPccbyQ=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 8576), data_block
5o7DNCVdq0iPbkh0QxMViJVGaUCEnMG5r+uWEwesyzxRKq6LXCTPC9whLlKRiZhi
NcSgF7Ba4b78IdBMRaby5Tu8scVU9p5sMYo42+J0LWe+TahOeKOM/8YmDvrl7Ogn
mh+6lHoZRiS0Ub/xUdPBqpku0y8dgQ1atKQOjFrSsth0V7dzczCyQLqqQxaIeEdH
SZH6oisHOPGmj1MzO25eaYMyoWN2+Z4OvoUWaxmp35yObkT6cxr7wWOTcsWMcw8e
tmi9mK2tR0shCFBAS7SvOGztSRXjB/uW9yZrheh0fXk5IMZwx0M4++eG5f+rkvJI
ImNL2YjBlJi5BAhBKlYnCBHY6TPdVZIf8AKldzpk2k72C7ValENzB+1xN+TQQPy1
pFQ3NP1QhnifFMqaf+9kqM00KZZwqN/44wOVEwxdjjikX+IeP/o0ZwieiKshjOXN
5Zm5wT4tBcngKHcAgLb3fQz6KJGl1nGL2hGHg/qNo19enoYiesei9PbKz6By0sOT
DyVJi2wt33d3UuWDMJFh4yQzYplMzjIaTOrPh7Z0J7uvgw9hRp6w/d5PcnmgxTkh
PfIhjorTeGRp9LOLF2JR+FZHsHylmWRfIrR7B+S7q8nR89tOVelOQMKVEZtuvtOx
lJrPeeDKv3xFt/jNPx7A8ujkN2rLfSthKtQJGJjEju0c/nIOUcl6BzsWONg2+l4h
ZqBArC6cyELIpIW/0J2BXrVLkN1Q6nC0i1m+xTXjFWkolyyeACrN5x/TTzWCy2GC
qRNFT2gFFHMne/VtMOeFAtMFWbA6ccy5bZ+84fo5bY7VbmV8o5I/EPB+MUA3KzC3
BwnPvFMSqGUpWRpOhoTNIneGhiN9MzH+Pf2ts61BhV6DZMcD3ESlpiT2FBpdeasq
pUhs8vXxaEOnUDmzpaOUzgl89zjyntPmnQiB8g7KQZTa/5SrtJ6f/Us5OTgMMb27
O4gPzWaGpuR7zDlFPvvAXUmrldZC500Q6oqMa6VE0T/5U3ATzCMse4A0o8a3f/zD
nyq60fDhNVJpD+h3X6TZG1ke5fgP8dNKbw2XOGbsnJIfJAwJEEf5ClYJcU9zc2RF
GqYz8Uvfd998cGi90YUlbHvw986XtQHR5Aa6EU4wDG7LK+i94tWNxA38l+/7ZmFU
f2sF5QmFWoynal+FU+BpQ6CXB5Z2M0eGSKgyEdgYwGVu6KAVOmwchwywr6c1TUKT
Gq6poGUjN+31f/eq74GqON0QQEU11jhAtdYnjpy0nHEVl9AQpdBnZmjz8V8cIuYV
SaUeKc0KK0wmHIBJ9e5bXJVM2aAZ4PgPa9p5EvoBBxCCjtZJe5kxirtuC3II71oS
ku8gmSP0mdljHSwbZkb/L2dhRvXXy7v0ocRKF90BafGOhVoBF3rNUCbMn2I7/s1M
IN1CHae3JBaifTTitWFQeNPW/WmR26qhPr5o+VuIMEO+Fb7ERjlpct7R9qVnj7Pi
F9BlsxjRxzwwZdgPTWbczMn1raxW2aF8GbnUEvDoRIdoQUp8xfzGZaNaLDY2thhd
QXJTUb6Km6786pn+XHbWIHZ2AKoUVkXqgxhXL53rYR+5VDWdsOqDXC9XiKHikI7h
KsU7YHmulejHvSe7ai17AuzVf7BfdO7P1PYArDzNRHfiNUmB+9d4baJICh3+1tPn
jmbvry9OYegJ7W1p93NXijmz2KF0RsTu7b1mF6adbRubW8Ijo5mmQsI3biv7pcb1
MT3uorXPaC55Eksfnavjih9tcvcvhvs9TBnlfcQSJFYWwqyjm7XRrUBi5kk08OVd
3hGrGRIUMx3E+peB9Fy7GUukAm0Roqn1cPSMW0uN4Ho8n9IhP8JOZaPCwuLsxY5G
rJMA1yoCliWqVqpKr+2P3tlPyin7RHa82etQc8gfcLr+7s46MRQ21jCmgLOzvef2
Tx+XTCeLpKTc2t3bxiba/9Sw+plaYqn7E9dul6++y7hOCGVxOV1LH/Gb5Tm7YbSW
+u9187NglLPvqfMjxu140qEdiHTaW13eQ0dzO4nR3J77VqwMN8USx7EOKC2/hvJU
/h6tnOrnjqFhXrJVDhDB0mfuL1sFsnbHz0WYLCYoMJUJNc0HOhu/fGf4O2WC8ZPc
vcDL1/bwxuKDJyr+g3zYh8P/wjHQFftjYbG8qMO8dGFZ+aDR66zYFVwJaPa/RPzo
PS9hcj9yerQeha2A5beRvvde0ol9f+XxsWPK9L91A+KK3x/hxUPbLkf4JImZcdKE
5l7gHVU47xgzOi2ZBRG3sHLnyTBR9IKOqIIIwQSg84KT/5+AdvuBzV7DBoycsDhM
JJH1PAsLi0mFD1HWh//hIm3pR5d2kIhFdSvz368T1YFvszJnbGK8L0ieYNgMmwZO
jG84r+SCDUMd74FiCjtGMgvUpU5BeMYLmD3UZAU+sJ9JBYOnRhpqvNqF5Ztc9G2/
DicQyhpa9Rh72cnVX9Ab8GHFoSUbI2eyGbOVJgF9gzNwQLxL6Jh8zZNPNZVmCnS8
b33guipQ/EgJr93hGqh7+zfFufA43xcK6iB2yP8QQBRONhp4tmXmiongmmEjBqCq
O/9CicAStUKRzk2FtM7bMFhfSBVwMeyArM1pYRzHfdFuSYVfSJkmwQFXRrpoiJ16
eQJGSu7rehwraNlxYxORjhuM0JyWb2aJfbp6VFaOVew2SC4Qc5MQ9PnF0DM9Zqva
j3pSC0rLcd1JsFoTR4vJwlP1aFUPBSAbIXKGxnTSLcwJFL+D8OK+8DSN6K79G9t/
ezyy8O8gGcJxZlCZm7eULaS8hpUMAyhsfVZIZc+5Gfr1uYbxEvXhF6oIJJumuTJJ
2HpdFeThYOJ3Nn1b/wDsTKGUfKiVTLo6lm9vP/pM83g6uo4wWn2dBSq4VzOJNzBw
sr9gYVUsVs1SIqT2uhi78000Z2AejepzucFWfAcB35eyhQunIbC7Mvv0Gt02IDpo
xrvvkBvnRawJCN/0CvXebnKTGmPuPjBmCxIV8RbHg4iYXxTzl1NYHo4IM7QTuM3i
VQDYlPqd+l+OJMlw8LrEAI40o0HaPiT12SrlTsmosNgHCMvf8Vh9LoMNesiIwiwg
kpvHexOc1l2oU/k0lSsTVns+FFO+LH7+InSgyVWaBHgs8ZM6zX+lPZfAIMKOpV8m
ErK48dh4umDVsoOXzIgknLM39vLHOcDDc29TpC1iS5654V8aWaHI6uEQA23bypgA
fyO2rLi40np5uDW1jQOZR6/LG6lrmrN4U1+xwaX2YrtpCtE2oqDGsbKM0ScylEL6
UHPVCWqZ22/KgLbEepwLzevwW/QiBbMQIQ09XX1ncqMkHs+v64T1tBh/YEkJXSom
YkxP/+v66OKEr0XF/s+bFzRrU7aej1HNXHXk/fA5vTuHEGytIi7hALCBG2YxFwhZ
Y4ni9Qotl2ts0E8IA1h5uViYDV6vla4s6NRnWqku9PMtkyb0m0ZtnBW+V0b7QrQF
CzjY0VWTlSQtzN2flZz4q9kyTEocPN4Y+8P8jp+31awiOOILqmdgtCWBBEiCSwJ3
yM91Nf9Midfphu2T6qbrfHw0ULuEqUVUX+TzrId2AJl7EDOK9bhtKwkuUbmEtbVi
FPvQlf7Dsb9geflH5h4b0+r3VlMPceNk8ADVjRQaK78IeGA9moIIfbC4NDFvZ3T+
O9u8T/kPr03bccz/t2fn7IS++xomTivi3eEuHqOij8HfIv967EqHpv6tCCTQVrim
wVQIvvHyfDuon0SSYmjQgfzSVHoDA7vSIe7yHwBGKXRtwctkYl04/i4r5I0sy4mc
PTeDuClX4EQV8DHEiIBmbDTKnbiZrQgKiZ6yetbkI//C/BsSMTuTDIDeTGxkNO2j
LeJYubJ9/piMmJ9ThnAIJJWNppn1WLCkrJzalTBphottTgT6ir8Gy1BbHqjM+5aK
i94GzTjGNlLIofy7zdA96QRc9KC72tt8U7OMxwvEhCl3/D+irctQsbL0mZo8wkhl
TzNlERV1swwc7G1YbKFZf5BA9bCfsA2+EDVRufv/imj/xjWQvR5FhDIqAw9wD8Fy
KdiDeY5L/Dc/zw3QCsnfHDYv2LUy+x88K/WqLrs+dxwRm6d8g1cXNtQX+FQHT1pO
jiB03lPysyX0OBQ89Iyy9xfmmTXZbmWz0FrcDvnrkqHswffNhv+W6usVb9/1CR8D
+Mc2bhbhwPVBkkT2pL2Xj0n/IR1aYNch9C/Zkb0XiM/chcY1JtOyqL4zvCPFj5RY
TdfaFZrp6enqMG9KmwziFz5UD5155BRMvJud+chVmSbfr0Xb9UaqM9P0hMYf3sXo
TjUsYrbSlApXxL7WE/s/j8lYWBrlPbLpSeUYQOfcVbHvJpC0labrN+iN28eV8+bP
QM6v2wB8jprfiUHVS1X1r0sFEzjUIDGBACF4eI1RDK8DAD+FlHzWh40Ab9y2EH83
1fPzAFBrfY2HSYUasBiiuBWZkUrYTZRo5prcyItb+uLo0poRbMPpCF84VRmimL/Y
rR+NY2jTUAfIhv8ezz+YW7PVkYqU4gFDCd3s8wOAt/GP1vEt6y25oY7h7RzYKx5y
tHQDdxc5Q/gK6ruY/Q4nlpUrajC0AsI4170p4Q92ODLLEEk29qz8LYOXvYlCSsQV
3aalTz3U/5BKl6hDD2ObJ9qbLBdBxskl8vl5fkSzdj+nl2tx70kpxkZAJgK9Dd7V
9i5lZgwWoRbc9bp2tBnbzhUyikEiuQ6IRY21qpnRRW2gWVUZPuDPi6G53hfl4C/E
W7WEaFOoNl0VQ2xU5r5xDrQKmQ1JTyDG6F11UPpn9ZkcwQJngevPEiesKDbb8neR
RenbybUjaZJ/I9EEWWLpTcLa0r3x+N9vPcw0kGJgPzmsQyLhVCxjDm07yMD6GpI9
CXMMSZCa0OvtSONSS8vx0WPb5Y2vO8gseJU4Ici1RkAnLyj50Z6BcYQ5sR5vnDpD
fRMPuzIIN3x77PPqZ29/oEOAPw3anLDLnVpwRJAcVEIkO/AlMGlMdwVsla0XezXo
S/WI1ydoZsRiECgqD1lZ4gG5qrIORMaYrmVRQI5eYFZU2PKRB0Kj3has810nD2ex
rihEfpl7ftToj9/HBGjRudBty14QYh7Yv6R8BT+3IcmBCtjhQSS60byo3I4Bo5W9
ajUWLnz+FXJ1rOIjiV4ZODyr0pEtKvkaV/WeIYpd5EGFxYgSTmZmjx7B4c853ort
73aIXjowbF+0FwfeWN7pIdajLOm/BOZ+zKWMmSSP2zhmYyqymRgftUMkAgrEutO5
eyTKR+AA4qOAzRI90NXF/o2ccI/TUjiwqXtd+rKbewEp/AkEUml9x/yT6DTwx03j
aBvNDU9OSHjjq3SZlEL2WSfl+wdR7ncC1x5DtruiZTNBtV+L3uEnmRK1FdXgw4B0
MuBvMHYjUkQFAOq99q81ioVfD6pRVgXhInAo2kcpQhKd7I2hMF1my8johDp9Z4Qz
GJBvPQwvT9bbFB4c9WxuR9HMEDgRv8hX8YcWJd0DILZXuoEGRvlC44UDkXn7sg+F
pm/Vj8yjK0jgxewEUr33renTmwqQTE9ccQ5g70btl8vwyAiWLf2sg51GM7MTJi6H
cgaIT2Bgzc99Z3Qtt37cEDfKU0X/4BH+m3uvMkXf2OBRzQiH5iEE+o/heFubl+OG
zmtKfdf75ge79jd3pSKYUyHt1/B/oZdxGoziqvclETIeu0jrIHz3YLe7Q9UGlyH6
zSn6OLGy6kRSkHU2xYEbf9TJMliwdm/WivDECJZrN0QjoPKgA7mcSbHZlqdsfT52
g/6Y8gD2aiRN8ezU0UE/3Gmi7T49fyOTeg7V44odLCaR1nQp+Scn0BujnFBUVnQk
YKuUHDSu5QGOFEgNB8i/DRSuGGCMhvIQE+yMWT3EkRyhPWuFibt6Q06sxtZxw1YF
q2tKaVMIGxxytaKE7HWxK9fKYu6rGwqORFT9YNf1oGYWfJvJnBxNbv4c5JMQoEyo
icfxk1q4kYQhQI8SXOz8vyzBZ/6Q7Pi4X0fGPgKLWcsolIS2k0aJFcF5YOe7amWi
RBry4P5hB+tIXxPQOvGDGw68w7t6IuInQErdfu+jsJGqSh6phJ8VoANKRij7P3kG
IsS4QfHi9c1/KP6+T+6tzMZhEt2p4thH3kbp8mzkC73OD7WxeAvIQz1WhEvw9ZRN
qhm8de0tdjX8/e5rEwbAoJECXcsZ6b/Z38Hy8GGEjL41K/cEgAZ78Vz4qkYGTyvo
e8gIDEoea0chtpLuYmw6olCJFGUijb+EKXB0k6AibxWtawKIiR4SOTzpYGA3sTWT
qpPMLspmMWJ1s1LWoJzbiuzuN2GxROjM6JE156kPkybLJq66B/KS/Pnrge1btKM1
+NMs3KJo5uLdWKKhkXgESp56JfsthAgJ01O+M+DdbcB7TMONlLa8rFIcw5nkwgGJ
2/RiSGXKiFJg2eHHyegO/xdVVAwFnhmkZgzGBiJ9AA46bnKz8NKyRtBBNlYg80bB
UVAaC/+E7qY+iN83cly3/AE/opzj/SS1hYHUSz23n1rcfrdWhAQKk0KuAScTszvd
183ZYn/GfHK//Ke/KfkB1CczEixHbP/hUrkk131IpSVvmeLaFB33b+6TxlKTHAzj
+ODUTqTItycPCtsxTfyq59cjleYkpNhlQqd/lnwuVgNGTEh3HXvfEue73RlQ65OR
QDWUqgTD81rXATwJp9buszzYTB3meOUqaaTDiLiqx+Oj/9IuMBtZn6HiWC+btYTx
OpVfsdGo1qS7ojeeMF/LtFJmrJBDI5Ds+tSHtw2fYAz/p1E6xo+WPir3uDq+1FpZ
Si0W1gJ0hFDnQVheikJUCWOZg1YYcg4EqN9/a538kX7PftGTOJF6CdWEe3ScZ+u6
bFwUDdwuL/hH8ulckSc+n3n5NmcouoGI31/bT668rLql0rw4SQqPMiXNfO7ix5me
sdzPL90Gc3IEauZ84LyxWkOyp5fML0Ygvr9UPewmvBv9YokruwaGiHaIQjCLDzKm
X7wLWUSscQSpOfkTJ6PcwlIQiOUn2w/8Ja/B2qd/rJmOeGZi0MMoVdmvpBdcjGVx
QohCUpgYWD+PJEhHCNyyD/M0+fMwctkwFwTtuo4wgEPMcjFMt0mVeELvIsmROwL6
pF6gEiF0sHpo7F88aAw5mSZu1SnFqzsE9446gzC43c0lbH6cKnykGiMnGLZrNFJm
dydjlDgrn20epxOjig3IauQJdQjI7zVAtIXHrV4TB3nE7zCHRtUbrQGlkHwzeuCl
aKRnNXyoTFTx2Bs8Qb9LIKr5lsHYC6VN6GoJmMw9+hHT/81wL0Im8NzCg5CvDSEy
qatzZCTbCtebw/R7NQnkbql+gU/5pRKYoLD/U21HuTf1SJ5eED6BjX1fqOY9ScTS
xxXr9iArVtJehtpfQZG67dvwmD+cxRPIWCH74jMmVhygdZ0O0SkOOcXftAk8Yo3U
dO5jQLEXEF9QRNLczlOGQm7bc+x0lNN56Yluq6bb87GYo2U/cCGSkU4/MeFvZn/j
Ry1dxRkwKU43A9kQ0BfqWtuNXRlOaygQNIBHrq22yYLk+vUcAGyE6+M1sIzc/Ksf
B0TksX9zIHhMOgndCRW9r/fPkoK+RJf8FRouWTUr8N0blztK+vqCyLMO6dKZtkyK
1tDSSm7qP8bIWleTCjLNABFk9n1Y4ciBOGOj9SJaX7CUtzUoYzR4HWjsJrCbWl5G
7k+/F4w9aUJ0wDRNYxRabDivyF/iqa7eWf90c/vgBYshxNZXAZwM7aHLBD++DU1v
hOZu/b4p21NymgB61zsYfoLV5DCAi3gnXM5/Vcbady4WAP3SdKX3kkWZT9F8Z8XZ
GJghRzWRvlcA+Oq42C7/BkiqhskRiN7J6dVesxFaVlzcmSF6o1PAe+h9f2B87tBr
sqvbKXTvAZdmWxaKrEBl1uR6dRytZKtbSw9iyN5eGVKTNxi4CJRe5QkmptWkWwa3
WMElgGZhMChsuae2rWTQ+Nx/t5IzQtHNxnQviqauuw+oyn3iq5fS8xXUgdfZMEWi
kpNmp1fQUFeiFKlsnAsdYEFS03KZ+jO5gC6KQ0rPkFjWvSY/gdy7AXrfgXXHsycv
d5xQ0eUyMt1fIn/L7O41fbR3YSJBUU1ENl3pRsRO5Lz1463/BSlceYrBcCGRKBV5
sp3T/5ISbhQx8nJT8xXALjso3bSLk8bQs/hf3Ss8XdbImTDc0YoWjLAtf2/yd1ed
5rBefV4HQt4krPaYkOk343dq4mrGBZaeKy67NX9EalKP2KgM32YOx+y7Fzff/FIp
h1WYmxMemPG/i6H6fJ57j6aNh1ecEtQyEXmpr7jCuMuaHAVcC8MFkd3oZeJ3dSRR
fK1hDitjI0Hiqg+ADBtniIuUGFv1svKW/tYUAcgE4CZHdZNwOQd2JWpi8KaxJ8XA
ZB5+nnMg2urMulDjoUA81nOz8e3t9PrKDLs0qLNvT83+6kSO81HnCFdP9yiQ6Jx6
XFH6EkF5o/3KMwYNA+YsNzVJ/OwrLOcROFdVzfwi+4SrZXT41/vwR47SNavziHp3
rMegYa6w4rxqWSdsXCTtlPVjsn8MYvesQaKzXQC+o7T/VOGKZgmTGaUAwtXmlP8X
3qBsG4L9kBh/yqLHHwNe/xTeelqGxbxXCH6mKJYsAkHpOPR2boMC5E4PkoaJlOUQ
9x7iSgF9/jT9yxeYqF70Bh1NXRbm5xy9WmCwVMnYl8m+cksArtHGxCTu6l18vkvT
dms9409eIn4AZ0iGFhf0EU1S8gx7mZhs/kdodr8PAL4TmJe6RN6d6LDhuMri/CeX
HcjL0usWlD7im5h+DYtxHerKakay9T0ZikqaRUB4I4LsS2FuY7yC2jYvSmZUM7xN
pPO4QWO5Sh6wElzIjdD04bICaC0pONa735k4zGO8kB6H8l1XJGd9wa+yOkX8RnZX
3isMTOLjJzLjzW6N53v0960EWldKNvcz3CleGF1i8eJhBfFGeDPEpyCqIc02CsVU
86RRg5sWdNehQRA7rIO36gTdmvRl3oAzGUzUf819Cl1tJSqExM/9LpWhaE10PNrW
XmngMLBauOHR1OW8AcBio+y9/LWquOXKdOraoc3klnhkXceJdiGgRATu/JyxI3xS
H+83S14QsfRLIBE2NuGUKwE6Z4MwIqM/9H9AOs/iKTPXUBeIQR4ZdmwhshXtaXuu
Nl/XVBBXAhrU4uGLPKJnMBY+dvOJo+cv5bwBozrKfyGsJmCABHxeqlJxfrV3u1e0
j0RNfpgCNWCEmI+E0BWinaZwgcUIqPvOwrJZzIGTC8x/dsHTj15V0Bml8uKo8gRn
sBGSsQ0Vxguw7UxqGNaqwelIYUXSA2nL0Bd7AQHTng7GWI+/Xnep1kMvk8bt7cAP
/KUMMTeuQiEVy/GJgr7zdEBs4rLsHjFIQaaZ7VPUwcEFuokUXiWlAweqYeqG+/dh
VLzhT5oVSUeSpMFvDUM09+owSzYDvebiMYs5t4VqF3xnPYx0z9kQniEPGbFHxbRu
5zkfuZmQSuCuIOlIIjWwwJ6777LIZJzUZfmIlo4a5eSJOn79GIYJ06MIRPpaQlHg
frcJnRwzUXsPRQgTKXNHb5nijr300x/8W2srXaNvBeFuSKNERD7CGqwJqXN0ZCes
yVBrUSSEtlXgxbrKEZLFgZaUQb6OUw6Oi/7EuvzhkeHdyBsy+N1y9AANW9prFbvg
o74YF5o5+m19QKSBxS9je9YAL5EIu0mhTiAfUil0msWgTxhoe1HjMWyVdgFhyTlL
jpUgXKCNFSG0b3tOT1AcQLEw2saf0UXeo6TpEmI4f49ytQlxdrRs8vn5f/pZMuEv
lOhF2kP2kADfth+Z3BRbdQQAfaHfOJfqkalMxfRCg9139pqSk9R3NqBUw6Z3wZH6
82PaYbKRtPfRxidnJ2fNa9o/df0Uowc4IN5fVAIc+2ls7wJhs/O2uuJS4fJtG6gH
DlnQN1R8zzy6cDo/jFcHOUEzu64Lbsm1wLYpvL0KeaiJ+uD0bv+9+Wtx20UuaXc3
qVvlFUGBpLv0wYBH927iW6w84xFkal2/BOJ30rEoF2Zxz47t2E3oOzUgM0FHcIUb
b7KCTlwUb/+srHCTOco9tROngkOoU3/h0hTFcwEcwdgvQpnvRDlIjYzBa1lVC2GH
aB851NWoCTHkluMlqU9fZMQat1IeQiGeo7OiMQU4qoUc6eLilLHccAREIOzymwJa
YEukh7VWbNDjPqvHvFDx20rRGHf+XpL6vMlNSFNW+YMzfP9mNDR4k41sUnv0dVal
QAOUKH1ssTxx6kMJ3F4m3PfQdlVHXLOMLEFltF3PszXGtdyGuLHE4HhDMOLIirqt
hfctH3acsQ7QdC7n+fEMhdmNioteT8Ghx5Ku+TD/Ebm964cc8Mgzxo0mYcwLD5jo
n9lauGDSn5Gp7EfsJJJectzrH4bWXtLNkubMB5j6//lOP3U9wd5EgNuPU2SNsalP
HGyWyVhOEKaXEEHKE6XHSnmLEl5/61++JzUKHEjlXLUDrkcCLvZ8Ch2rDqmu42fP
Emx6RCrtzSJAn1bs3VrUcjg2S9B3K01l85mZGYqm9e9ChUU/RufmnmuVQbw9FCVk
20QEzxw/1POdoM42TiVsHATdpMPqisb1ygtP3S8jLK8OUyKMWA3bEj6qViGMk4ZW
QjprUfRLHukch3KUP3ag0/L59YICbpOHmB28sZfGubBJ+b1Qq7xxYNB00F+J2Mfy
4Flv+ROUYfgrdh7zuMhHGotjrVRI5oJSzZignRB2VOrgkydn3oeWjBcjKvvXAnlN
+D2V00UJN95tzhWr3YUmN0RQn1jO5+wlrSEYDkYaA1tsRCs2KzofoZWmp3/hZPHO
ihm5CbRPLEyvtoaAcKLDsk+riDVBUi+FFb8QMbs5+fDXFzvTlPnYI2wxAe/3crrj
SlOoSXQytCTbbxoKn/bZltn7EnR+eEKqW+uwssam3FD2+G29J+fBtW3WpQ55j0sC
dWWtVZ870KNd26Bbipahv+sUPJy6CguUKJTOqt9VjqtawpH+d52QjmQR11Ercflk
pExcYLX31rAxD5fvQZL4vVxDkIk/3L1RmG51e44AZwvKI1Z/R1FhZOWyJDk7c2Un
ElocwufbUOEgJ++6xgQBTR4E0m1a+7n0LWdDdyuQQvm8UdWQaN47o7aodsrepKlQ
cLK97zI7wyz96UHgRFsTlUFe0Ygfwv2RDC2FjguV0kCA3Y028SlyjEcr43pQFNjg
0LKmjzegNiqHtORayQsYQqkSOcVxnvQyl0jUou8+AVwt+2EYqgjXiRVln3WrIKz4
jvFd/+hMdWa1hNDJvjQ9SRv4SAuQbr6L+X6b8waZTNw12doTqKENBzRHd1n941a7
VHAY328GmmyVDYyHloWUw/LfFzfIyBUamXU0Y6vN2hfE4ep0d/Xs7aM6ef5pPBNH
3olriTVm1Aq/BQFihQIHXeF2ETfZuXAmaVPfilod0zU=
`pragma protect end_protected
