// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Wcjo01hjhifLLRGDibynossTLkMCP0yO4udOrPm6ea15KsxyoZ8K7RZsgN1q
eineS05Cu3SVf/W5Brp7D3nAztyEgilNV1bVPKDvtcvzUrudhX7QHIkpwNk1
G7Uimrntj0ra5WVzYPODzd2THkZo4bmciKYJvWqSSkfPSMzZPGOwQH/MEtv7
+YETemXh/wJ1qGRnmuCW0QqHIh9CH4atOQnc2/fOMuO5IiN5wq26BJkVbVvp
zv27zRxSJY9tD5PGm8MuUpEJL9wBhcQwdM/uSrJc9RTihuEvf+SmpiinAO+S
mclJP1y73hRUS9q19rYcf1mo7zskwkpMXKjjVk24bw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
LNkxnBhwKFYdO4eRvC9D3SR6whD/EKul/5bz7WcFM8A1KjIEVW36q00uAqhF
DUtnuoZ0xN1O51TPS6C3P9dQfyzL2YxJqd/gPNPHYViLh0Y1I0LLv+CQ4XsN
6UEVOY9T8QkyMrnSgSDhwYTJCAdzoEWx/XkOsYXktATnDfcxFFRGKe02/1Gw
TlNp1vhEOTaemnpkTcR+nsrp2tsUIloFMmreVinnfCvJxPxrgf7S4JFWfOQT
r/pnNmmjrGRBwwvuf9L1ZYzA8M0NVt7vUQL+Ld1AFECgHMzNjVJrXHy3xKoj
u2JIJtNJZjgbkNTG3DvdcBTM6S7om4XYtcrVPawwIQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Bk6pjakVQFokabSAsy6U6iTCbs9jn+ieHWH04OrPc3yH5E5AF+hIyvl5D+Qc
Vh04bbudpXzcjtrJgBKw09Srj8dtx5rxsPIMHyKgBNHbrI1ZN7gcM7JjxKwI
CATqgCefFeOyAsaQuIDZJickeilbcGWsYJPuUdvXyWgdxQluB4S6O49jvyvz
IWAunkwwmPDoAuRzVjDcUsh93xG6ycYeKpu3vsEumXGa8YnYhYBIYj2voBiF
aRrJ+DvtpmQ/f3Wh+rg2PjlQZ1QBOAfw+qRODIDav93pbXkOX5mJLfh5MwR7
M3TT9tlHZOeNIGZZKGfuhLmuc0ocyzQ7ZhERW7v6YQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
rrf64rr1UjkONSldDxpnWhpfocr2Zh2FIbAxxja3x4drBBZyFofLzHnMSs3j
dyF9jipytVNsIh4xNfx8H1cIO8LU5vctMqUWqWnak5+IwbvbcAYpRZH63wAT
rtcUC9AKvsbBurkv7bsQ0cxNv+Q2w4/Qr5WUzlosxZMJpQynZF4=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
sHuYgWJ3DzhHK12kz+JXHiLvfWHBqaQqnJAKOEiNO5GRwFn/YCtp25R85S8M
4pHaEYp95A8lxo0Vb8FcrZLRuSP6bSaxrbYibLrNPczTGf5C6qBPWKIeFPCC
74t+9uFghb+hCtCNRWnvGuGVgyyibTVeOX8rlN6llZ6+tFjxvxA0jbHYh7LK
WzsFX09UMt3D+aCMr2s5A49gDyE5PxIC+1pUVsHrIZBcPI90e8sGhLKrlCbI
HjClEdeOjWVg7EKY/nVAzj/HG3PPyF/8EdEcdEdIfuoR/sXCTR2seQb2Wbsi
IntdpXlgQpRpm7r/R9OdYrhMWVrg3h1puVPCKGN4PdW5FQtrx1VoDVE09t85
Op4O4EnAaXvQJDSlFPn97wY67xHq4hpEGncC1v6bwcENuVLRpC7Yl0XhBlJI
8YHxQSqwk7rQ7SAoWbhGByp9d6xltDEwO+7O9gCmt6ZfkEK6XFYJe9l21z9N
ynl/EEmf5Ux+AMXKWCb1Nr+FL4cL944N


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
I5SLbjFLcs7nZYsCMgyvcLflgs8FJa9TleXNOkzYk86aaAX3ya2f+g9midHT
OGSj112Wn2Ab04sWHk3gH8mso1zriT1PhXY3b37Lpjqw7+vuwFxtiOjXlSa9
dQJKMtegbevzwBhdm9WOvGLHU8AGRycx+4gnvq3BKK++8xQ4AY0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qDUr1vQSOCHqEAFA17I8Sytps6ulBziB3KDC1z3qVk/aieALaCU+MXS5WHGD
IvfZqvYaISNbgc7uUnb6BugLobhRkzKpPwDQSGqyhlKZe0vsyGIYazmzLnfa
mDcjliyvBot8t4HcRgqzMP4WPLyF1Rf5X37aX0AbuVr8PZjN55I=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 14160)
`pragma protect data_block
GblrUYlIC8nb1Z4pa69/usenHET+sZxUJ34wPcZfWTDT3OLLt0rfYj04G5pV
5//nrKcNrggH+FJ1lB30/lsaqhgBXfs+Bu5plRebFOcUb3155hkV9aldpp44
4WOZaDe2o0DSj7nHUJwno4ptZGg3Nd2FlDZUOEro3cfQJJG8LEEHhDIMqkjZ
oC5w8ejhD7ozA9tlEGANLjQpmhegSOzA30qgFwQDq4Wz1Zgebb4JxhwjRCXi
iY1FPn51NTiBAZWjVQC32Ve/jyU3cpjDBwxPPJqm1Eeb6OakylBkoLvODL+f
pLTkU4bs6fU3+3pR3wObW3/JAgjgD0vEZ3knJULuqNJG9irsLpQlhO1H/tVm
2BuWBUxHQpKQ89M72bCRXQBOBTuE4q0vhhqryKmkq4RWlc98kGVar8H8jCre
NbIMStRKOoo5g494UfIJwuD/EmjwAx8wwxOWuH5IuAMdm+/TbbpjHXFFfQfj
HDOn2xKav16YHoMSryj3iI0cOe54n2d1vyOB9GSyPackGKolE/ItFGdCQ/4J
LR5gdKdlCMEwXHBbcz8piDjir2ZYNHogebPoTtA4HA3BRGgus+wdE/wgzZKP
mkUuJEYtJF90vhk2ehlY8Upxnz3d3g4J+bs6DuR5ZrTzGbXptz4PfkUKHFll
DDu4+KKyt8MFqWvPtZU7fSjou/O/O30FfV5kNItpLvj/FwVfpIEfVsyWUa3a
37QMRQCqvpy9K+Iqhgs1vj6QVEhh4TH3fBy+9k5y8k9FaGJbilW8/dmSdljY
g9DtZ3oOSrmeW3UT6ZJq/EIGAMJ8m2oW8Gk5fCNbtgy4hTWgWhifTwkJsGfJ
pM+BpqDbgOeU8RmIZgGxm39WgBMKWVOZFLdKQPfj5+Q5Ci71+UW7CwucZMC4
xOulq+u+AP8zWbLXrxKQ/blxEPyGvlqQBrU2qwuM4Keh+4iS1bUfjP3oS0XP
bfqn/f6OhSuaF7FfVOQyIprw4c2MkQPHi0dBYWrZ3OOTOacnN5m91xd4hjSe
GQzLVjSpsELro0qoircRY3R5pKFvku8eTmfJiAwbpbE/fe3Y06BkdV0TALnk
NErxo0Wt6HYmI+/KeYeGhNAI0qxW0sJpOP/8cqvH2GUiZUpJdzzDRqHuxt3V
1eWwFLUWfnpaBdcWs//IFmUxT2gSYSA270qHwUkaHUcd5dG0r9rfOSbW3pUh
LPhofFfd3oXyBLnUIW7SKP/GISNi0UJJ0pyjH8u6FKh24c7SXhgITzPBZcnN
EeogWfcOQC++ugbZkH5M69p2bHjovPWL9uxSMed2tXLoaR3cy+VN8jMph+4B
Gy4zqe50qLXMlD7Zr2QcK6Vy2psGELmmBY1aOIdMTh6Vj6xbVr+w7vIVjHJV
aWmRTTIN6ZV+hT/OpgQb7ab5/3YwQHLkSvDTaTuNZbCHDtjtoaFxXtEOx7Z2
i/iRGWzabyJaQdJGP6Ff1y9m05dkH7991wmgMmpbztqD+hHYTB8USPAp5pGy
OyMbTJ4tj+VUrOiBiBmuJVs+p+EfVxMevcfQCC3n0f8Qh6RbV612gZ6CZPlV
3xXI296Pk37rS1+fl7kWa4X4FJnAnsxiVw3bCFG2aGxSjnkpgVEgq+sDaD4w
BanhYziMoilIm6VlxcBhtYZigrsxHUEk/t4cowmW+HBaKX6dzaNhO6nhwrxl
gr/D7U6Gp1OqDgacMXYijIAuQmVKqnXfTdaF3ED/Veahd5ioSSr0B+WhrXDX
EGklR4QFyxOQlmVSb47zLvLStqK0mFeAQERYIGPLX3JOIpoNIwcdnCvWB9+C
Ni3/z4ghN/GCErxuFlUH5yOBqcI7wyTVVWn7WHzB7lhg8vFgWxdaReEwtZXg
C+muzMXupxbp1diayAA6qp63Dho9/99LNXKdh7/FpI1ib3+Sv3PMDK72T6N/
XQQsILa7tT18pWg8ZiuPE5narwY6ZjS7n0JHVEbtEqWjxsbMHZNmXDzUqn7M
clQIHDQT1c0Fa7jOEYawm2ZDx7fkukT4Anh+0fS02Yujgj7GZ75RVhcP9b+K
H/Te9/i5o8EY222Yn3OOcXAB1YBXyV3H0bZBpq4uuZ1OQPXj+0sIx7kosOBk
LCx2G2/RJSVnikgIbRB2o5hGevd6KHf/ynmBBa53pq+tb790s0pyu+TCzwIU
DjSTzB5D+ALLrXZ34xOm3NZ0msWNLkMqBax9fwB6zEldf5wPAHLEHxM6VOui
ziNs6cKLS3BBX6OtoYLvKXVm9C/9yPesdR5g3vvD400iDS/2jEwG96WR3Dlj
BKH7aAMohPtmh/xDP1WOJmZcd6A3GYDNEI1zQae95FxL92OHQY9CS4yAg5aj
egsRS6WgligGNlhcjxsgO181I6gYF/DOfhI687enamm782udHNBnGSv1rtWd
GerPAKHkkJX0s6JrQU0fCscgsfzuk2DtlEFLSklOlkJP2S3LWKVBikREjwfY
i9eEpH+RTIxyoIPxr0+/8bLpzKHTOMsJyM85T2BMp++AN9hsUucc1C6rZEzH
LEQNLAG2/C1gFKCrCBNx4x4zRqUqux8Ey7RelN7fPbrDLJ0Yrmb4v+e6DXjL
bekmeuTShpDc9MMWSZRhnzzrvzc/KB6AZpnBlvrUo22yiIGpBCYaJVmDssWy
rP/q5njA+0G9zIXN/FAIfXKZ2k5nnI89L77pqeRVvTljdV6QUYyOPAguWAm8
qmr5C1/7f2+hWqasU6h2+Kka+xYg9khqtk/WwFWGkn1Vj8gduLBs/kKZ2BpX
DU2luRiLTdY8i7OXZIYQG4Tw7qtkAqT3AyzOv+I8fFxHuhMMJI8KYu/ImVLr
nxJv8lqoKoxHfw9opn1WQsOd8HmGr0MnHBkI3mZ+m2h7Z372ZE4KLuxi+FZ+
pR/zaIZNSH70eCIZzfZzbqger3KuRck6xouIuTFaQLXuEiZZyqFK5D/NWt2D
KTvr2R9S5WVe4LKSRi0rKwcIS9Q+Seoq3U30JPHecxCPbqQp3aI6TAHrNfdE
TuiTyqj/aZqTo5mS7OCpRvBQ314ATS4dfVgk1LNQ1rUrSx7ef3hTiFkkVt8K
hPyeg1rpAqvaHLnvfqyCvhguGoWGqwuJbsQdC1jZ9F1c9KCJibrfzzCPKJ2B
dxVgdVS7fXDzHDhdDwy5I9opqIKI//py7JEUxOy4MvZDKTUBvfGfyEubKY7P
xup8yYUnqkN+jjvHDWWVrg1QCNkaoWuSVjtB7gxTmAHO0hmHkwyezyxKp3ZX
sQWAADXW0LEaBFA9c+T03mfTtnDa0HN+0kjylgb//K3PTnfXZ3uiPQc9GZWG
Cq7RTmInyYp9T+EFWsADoZZcYwqrIvEwiefjIu8hvNTJuf6XkTtWz11L4So5
qWu1nM8qrFNiGjSPNQkV4+OYXI46fOIb1+x7N/vnhxf2GsoBIdajUcOISnrW
rvy3XDTKkJascXmyZhcGo8KMo5in3UcuHKZg5V0UILPzqcbQc1ugmdyKi3kB
iPW0z58KcI+OLmsABg9djOFXoFGM8lSOxTYUFh4sykhp9LMxzTXP/7TAo9TG
eurEFG46yN3ssv6KblgNpQDuglta1yC05g24jkuFbt5oqOfNFviGWlDr7PDh
hJssGWmhulqOLV/oG3HBqvUnHlybMCy6dcH1WE7u0hRGrkMk0mqd8xD2V39g
89TPWpf7P9EZqzKqkzPWjYk/x9E3WVNaYZo6/xVhPxZK/oFFipS2MvWFgr3h
xJnpVmjazYwFp85INZ4eRis/cyVxP/v1ACPnKoVTgC7aJ1FkyQRlimzeVZbZ
+fnOp3MqDRp7IPQch3smlsnV84MJtKGDLYBV1FEzhWdNmX5T7bKrGNPMGhzc
3Aq89OUPXuIPdYAkZD+46tvO+GjdDYKqhQeWTMj6uxlzH0h0VoFS1T+p0wbr
LHe4frZxyFzs9S9KrCfafZXkqqxQEX9DCj0LAqM6Ug7a1Q1bZmazvViU47NO
EhsDIsSHvX52Kno1xeeLUpWfA3pPemmup9ImpmgUX3cJx77TOk3kltVZASDA
eH5B/eBJ9BcuqDLfobxgHPUUtfNy3IN/uDh5Ve2orxcvybLy8owff0QPpdV+
w+AUgdWPmgSMcTqfAcQWZeNvBdZApO9X+WX1jRG34SHW8tdc7aAR9EbS2VT4
9v9hhwRI6t/hqJimTyS66UypR5QZt3ZVsRJwOVtZmex9Dac+RyIWyRW0LbrT
/q+dKQ1VenBLgU0OEReRIHW1Gx+FHxYafMMAYgZDzjkfn/VwpEDwhPgHEqnI
SIPIAsqTh1t0Q9OjKLoXviLOIo0XrgXJfM31BESEMTiZsApafEG+ZZ6YWGqx
Si9myhSa92+4j5bhn1nB9wG6oiX1PLGkGvnfi+bcD+LbCUtHfCBd1SjTe77/
q9/RGrpJgIdUF3aAs0pDL5N6DAxrRCp/k9g9yrHTQeVj6RprrtinUjNRocax
pRJLJ2go9iucovNb3AznexeWzPhjTxdki74xMJEaFsdjcqsgbNSU2CANUo4B
s9ciTTQ39hbjAI9gBAYbV1fUKuYp6HF2GdvnzSt4QjUpbNHcUrX7uQoxfhLi
5bamrjKcCgCsShaJSmdLdpOjzuktZD5w6Elg22n9dRch6pRfZ6Lb55y7ZxFx
I5O102BkdwUDc7f1c5lvgp8+r19GrJjkC+Mlx7Sm9WYzFHCm+vjfAItaxj7K
L4w2J90EP2olGRDb61NHQqcsIn2mcUMkzE8jAp4Ss6WegLaniMR5L7k5enxh
J9LxsObe7g8mCvrn2UeEQeSNbQX0/KjzmbGW3uZxM2lE24IKD7CA1uOZcGpo
kgjHCAFI1sz7/hiGsUNSFLjWfZ6AcTAOTd79TBKPXar2dje/m1mhyu39PGFu
926IHCmi8A9vJuJ8CJCwTHBGGw7aeGusZzttPybxn347GuU5sRf9N/VoHrbh
dZS/5r/7m+afK4xxkF+lKausN70PkkOhpY1sf5niwr1c1rQDJAYHGQFMXZ+J
zaf4+qzR8ZqgVz37L1aFIUOfZz0nyG9DU9JjTw5XeEHRRofjm+GP4aSkzhDs
wsWxQ55/x/nI34spA2YX8Y7ZdpNljtECdYL9nbETXRbaplU2HbPSDC15DkBx
+3FL4sSsFVbTM/hELhF/pbJtE/3Z9RIhpJfQ3FNX/nNJtrsO+HYh7/hj/sv3
8eJvMZuhWYWQasH/eLLSdt9MgQqXSmRxSIr+dTEe/pX1rtAm3wNgEeHhQG1H
kb9Fy+7FkVFGCD3LecufCsWZIflJapgIoWC2h+nNHQ9rGeN/1EaO1GgaWoCq
G9A4na3UZulV2z/MiNFu/SzNGX29cMy55Hp6yGu6Bp7xQp5QiKLZYDo9ytY4
xqZcwI2MmfpKupp0WblGleKmCb2UeNzM6z0GPphHZDKYO2jSB/NNJxgOGlj7
r3Md9B+Z6N4hHKmoygis5kzlU5R3C0sl/a07EaOTS4ceMxRkF/x91YZ+rMVi
yuZ58tfwnZAsGNtqLVJ+RgqvHyhxJfB8myiB0NIABjlAaaNE0Uy6KNMWixti
umlNXW2U1SIRGgkEWZvnnHNGbEezlZ94vnVxZim6LZoVwn6YVWLxMkDyl7ea
7Q0LKxkXl+nV4vAwqapO3ltuQkwAvkGpd0NDmYedxl9HG8iXnXlfoNAv1FkY
VxZqm9y3i5xKjkdTmMRKIEtGhm3631TfBBWDwSEK9+2MphRxA15zsox52F/G
uyiafJbdLQRehC/mdiQaAIAqMl8JodH+FubqFTLhX5+rVv1g6kCwJa62a4qr
9kLgSfZr3V1Ofj5ACC8REUkSdTHtyNJ9LYxKCqKMy9h8SslxzUV8wPUm/gqO
DGqh8n7JiArf+EeIKl0240/fmPBX1gtrHS9cwC0nhBbV7u76tCoDjzm9yiPW
oTqyVYcn680WO37e2XU10ArrsehKtllprDE/hPJAoksY8Mb+rtS2AYGUZuCy
h6sK2L5AMLc9NWnOu1phtNWMIk27lEUEfSb742bo5snsX9rYJ4v7b7DKOoWa
gXsMoLmjxmtWmQXJ0FKygwkFfIL+c/dRdo23J/W50myTOtEBFD7XaLd5Bmxk
TDKj04EWCGbNaiUulWj6raHX0eKpo5kF3HszW1Fu3pEXxXTSPt4SQnfS/rLv
NyPch9xng3rceXwCgaHfMja2HdhkH497yqY/9ctQcsc397bLQqpCElWjRqxS
Tm+TI0lrsx76SFoIJuZDdNIBvmTipBOYxX4cdkZbg2N6ozQkz1EguwD+MqAJ
GLr6X3TuZWW0Lk+No+VLJRAQaxNS8nuyG/6yWWYt9mY/NwQJz3LElGhT+xKb
AzmqFAjcndLF36Z8eeG1kZDkp5uURXJ0ezprwv8wXrVyTawnsP9tY8w3kae3
iE2BFjCQLyotBdjU6PRfvDytaFuR1i72947F7IDREqh+CxwOEWipEhhTE0T+
NwznEhdMshbL16krM8sBnvtoIyaLcKbk5Y+RrJP+nlBlWJAe8gWiI3686+Qo
jnsg52UqaduBpnhHXZ5dY0kJwbaHbPtFK+WnU5NZKlAxd2mG1U5guXcamp1h
eNfDE5chQNwNAygNtKdts1FNG0KZDEuXxr9WdBVRZwki4sLNu90mQp6Zal/c
EpRrzSfzGJCrotbbSLCWfWlpjQEaUiKVc3idrdlrngpE+/fPgXJAYGcdNKFy
JAJXKnY59nyXFNMj+Jek4FjM8+czUApvOu61PLpLGkLumATdfpxjKd9hBm7h
nSpWLnwKBtL49ZuRCpgEmAkaYmiqEIp8p16Qfd3W76kzM6I2X5VxRJOt1MaY
pJpuSrTS4KOEooYhiBsLLfAeVprxi5sl4+SG+YEW1B5pW8nI0n33srRmnZZk
E/JzslNebuozc5jTK22PBDg9HzwqWI5wQEItogb+/No/NF0VXhi4SW12iFTm
YEsMoyk/ZENvjw5EyZHwg+VFqRt147hhQYcv3HuXv2dKF5L8gskGcwkEk4vq
cKro5lRfPwXW085slg+uM/3/yHPt/HhrZ+JXaEk99/RweJ5NcPyEBiCxsJIC
tF6DGlf+TNSNae9LWpJC/GIn61U1cezkW6r/OoBTnqRuxsIUeGSE6O1nJHx9
c77GRXgsKoHk8vAoTdTKIbNzu39g1ALrS/e+CbeztlSJYJNqUyASoiCsVRRf
dchdufjNzuCkR1eoZjCF4dAeZG8gF7A9T+TUVpkGttwy5dbzw67r037vFe+y
oXWw22EQz91JCdwJ1xUfTvfy6Nuw3EPnNT85jBwifL+A5pl8VzizMYbz9yF1
CwlKwnYRqnIDdr9vk3mTEuHwTAWMjBvk6IlgQ9IN5hAlcs6/OJSvGpxeJ+zD
wlHgYoBmJy9I3TReef0LngjR+0xW3uSWFplZf1397KMRZMAajd0fqcFdJJ4i
qeYpnlHJJVNVW4VsFiJKgAyZ3g/G9LzXE/f7f1wKrfxeJcKcFb07LU8qx+gl
rbJGfFXdyyKXU9ldrontYq2hQbrbtRkemYle1j8aYofGERCOO2xSMk2W2wfH
PnIxCEHGTGLu7RFSeIZtz4diuGLQ6SwAx1OqSqICmoMUqPISZkLZczOFcz5W
SwL0HR2tJc3PMsMhSmCZjkh2dnqr6EgCXHCYsNBr7rIYEFm64259/jVb2vZZ
1yXs6eilapKVWtfKOwmtZRqSgVMMSp37GWsUh79Oouv42dE/RSXxtCtNBs6E
AQtXQ0h1YaSzsB4H0ufvZ+0pTiAzYEAaoDPIv4WFNQUb4FghhO6nVVdGFhUC
mXB3jtAAu0EgnsKAcw5OD51GVzBCqFTP0KNlkVV7zqT6CLX12lkVU01HEUQj
yhIcfNLRIxrinGeFiWS2w38beNUffzumCnkZ3mmlqbNI3EYY/8Kss0Ihk9TX
8AGBqnrqg13HOzKp7hKNBfOYBxCS8tP5gDWfmRmwsqxyIY0kVAYDm24W/ad2
e9T+k8NOiKcqVU5T0/0QeKYmbLb/UkdMmy1O0SOW8Fqfr6tPwNoy46uggxki
su8gN5QPZQ9eT/qlHPaxTYkyfA/q3ULW+NNFmicAOvSvgTtT+vWDkKk/0RIt
hhomhpNk3pQjZmUTzaXOaoI+mNR6Rip21X4mD86MCW59/GUFUQCrbiycyt0R
16KnBzDnpxgCBoAYc+6dg2b6rLHG8UQu3A+yhEz4WB4gFMbpZQQzYmRDHeDW
f4vvJZ7cIf1EfFtHFnCElvOW1GYdJXlzyjFoL8hYCPGajviFuLM+c1aXyeTL
Let6bf7nQDh9Qw0BzQLvh/EP2PIAuO37WEv7+fZcdYEEYWiTSGpU3CR5S/Jn
/pubFdow8vb2WF2A3l0IboffXORMKhY3aD70uW/9uSURIyjGtmd4ea0qzxH2
/M2BWAPeP+h2NxU0uqkOhrQiWoHzaqSyIo+lUTymY5W/qVhFjm57pksJMj7A
HQaL68a5L/yOz1Y0+3AWHCCd44t4vyo0UT90h89IbrlGXtN0dV3LDKyxzzej
RmITQqlUs6FbpnpqyC8zmaJA8ve8i89OtB2O4DA0MTI8Sel+N6jJ/Ve6VhiO
Yyzf7yZpgSQZwth87aFM2TrZuCZ8uD69setWxI1CZz/RUAYZAnHhd7EHiJon
I+cHH+RS+bgCb8btTdPQz33J6JBCnmZZMGEeBLZw8Ee8a+YHzH7I19tqVEN1
/3bVO7KY9fmdI4RARRZgVXCUC2iNViJW6+fUNCQDcwn5JhadJ5zAalQTl2/3
PH4cZfd2ZqhDu7JTEgw0Rc+VUVyfIr3ULeN+ajxHJLgpDdifHTNG76rc/CAp
K5K7QyxWzhzxlT4fvARMw8W2/qWXMY0rydldYNTBzqJnuigUOVVn/hHUG/oU
BMJk0qgqyEjbs3UcM7yJZ974iF3PiM17r6bxUFkyigCFl7/C0/OKv5tK75tp
0fC55bRWWCfv8nSl9YeZ7BcthwBeY6HVmY+IdEF0bbe8qoIR5rgatvnOsmT/
zkHSjHIEFWwTRSGHgdIvH0afgzv+b6vOfjLQGhkh364TVGHfzWkgtibSu7IQ
os28NLejXTp5A5zI3kl6E7Lc68SBm+D/oIgn1SuXdy+0F4ScaLK21qXhVTKw
XkK7UoMZVokBAKh/iVLC8HvVTjWgv9topBMjm0CvT9FQfBLSXXZ1PFTNDKpo
5Hz5u1f5wu34yufVvkkBGTqoNStKEvWdPoczRwhoBh1mC6mgRoYKrt1jr2FQ
elKxwRPWOsLvPUpLeiKM6fRyIhcGE3g/aexgo2TCyzTpshEMOYyQ1kGRkl/Z
6na9+1nGMXdLo+c0niVAtUYA+uXLnxFy/YGzX4no9Ew0IiiXaK6fNADdhUnD
Gd0H5AkJp2uTsJdeJh8IfLmHLG/ISDood40vuwo5NAl439OXaixP14JNFVQp
kwlO7mZwpy9c1aVPMPHisGvKLTo5MTCwHzoaUAVPtIMYOTTW8bGEDuIqndn7
TLRZN21sPJ1m5BuNJoFpRCbpLCexd8AGa8KrVPIlaivHXZNBdA1d+2RjmbED
pHrY2SOXP1w97xxCC22nbSZqF1GHuXYqAarN50+Bp6NfCtZUT69uNHkIlK8T
k/5p3k2H6wLZ5YGdBp6blOEcUnDQm3689GRpRaWtaZLMcKVXFmtzhIJoWVd4
XBxHnGGF9VCIJMC5bPDHNARIAGnh2HrxZIpb5+tLQpYgh8tPgNbao41KKRqG
nrnYyIYqO3PX3JbMP2Ue1mAgmLPF2ZHPhlYvvW51mduDQqh+bRdExmimCGK5
VZs9X5DosyLaOaEbwoY2LicaZ+GEOzMBgQuWLubPSAA7wtp7cQUcfAGBv+kg
a6VCLbOqK1WegTADbuqUZePNyIfv6v5vlvy1/fkeM4058AAzQq+buLsQF6RF
myt8dYF4VeyA9YuiTy4UlzGO67Xhuj4/9KFS2sCQLM2vPBYKDmcB9b8uBuuZ
id9hAi/vlV/6om4eWRnlOlk9ItKZs8LgGjUa9njSg168RRwwEfgPl9plOXB0
RM5y7QRukuia2X1IjBM/vsHFiDDdePrMClqi6MV++Imp9S5DcdTt3KZa3hGT
03w52XlHxrhLDH4KTQxc+7JSqWmmPssDwRSdUoMjjD0nHArBR2ziN3llzTi0
cZcT4E7PhcMZgfKIk4nyTCxWl8dzL80YGUReIDAvS9N7CO8KN3ubg4gMCYTH
i/7OQ7Ho5a0NIL+Gj2gtkyiniGw3GJoAn2yyZ5lL2DJGk0vYXnp1XWZVET5U
y089DQKyu7O5z7GQQzFzLIHUdPb8BojpmXWqKqxWnQWgWpZPofFdru+s2gSG
SBcHNE7DG2dwpDMg/uYhj4F/Fw2KKTduT5LEVTDsQc5g4CHt2FRHOYhAkGR1
NrQwU2hE98xq6j5pHnddlZzcsAweHPcOPCjbjUa0sutuQw5XyLfALIN3puUv
n8uD77klcOIghPXGOk5V1treaszj+j3TMJzRL9EhiXRZZHBPE9xPrsbHkffQ
rmb7vQbFoOxkcSlUxNd1YtImc5YdtPoIasRT9mq//tH6jKobp0H+EKZvofZm
SjuH3V9uv1mD+i86w8rEBh9CBg1eKXbKywgkz0PuO7LFpxO3YAot8QBKbayv
1T/DcEMWGcKP6gdAUI4EQW/hOJyrnMfVne6UMnEdBbdDhZ+jRdkBMp47ps+P
UJup0H73FnetdrgsuMWahP10SYW6sRFO+KHYK+nCtOgVz9l63oso6Ysacb5G
o+ShPWJuSjYBqtnFoXB6P6ZDVrpkfbT3Q8Q7K+B4A+184Jx4+1PUHAi4RBfI
BiINa9z9R0mPkXUh3UI8QyAls2TVSkpLp6YLrP3k9mTIEw1IVHprqpQHxDNY
ZHXM+il3GUQ8GHsR+Zc+eDg8UKJk6S3mE4R8nKSp72F6S2JjSUSqIjyT3Tj/
oO1vK6ieHxLTF+t5LD2XqdV8QsdNayb5Tpj9tXhcfqrskcOQiuBIxAWjH5tZ
5DPPM6Hiee2iAXO36S36VdoSriej8aupFZAQbgglK7r2BrZmJO0WIxLlhj7E
9wiOiTmi3512Is7fohuVKspR42MdlG8O1R6iNB+OFn6HLOF2zqK0Azch9roR
a0YHqHebNEXrTmCXwEFmT3Fg8A7sI6r5gH6k3ZLCEaAQIffmXwgYiQI83qgT
gN0IAf3tV9aAmvgIBRKnC/XsA86Q7uGzeIt4Uip1KBO8KO0YH9G/7TqhNUaf
JoEunkAUI1R/t3o+RfNKgv6sUHx+NFhLDkUJ7m6uLn6B3rrqfvm2vVweyuc+
d794KATXWDoKWRr4iW95mh8JY90KN7V3zp6McyhDDnUuwrxhLRnqk+IXotpX
NNaShXXhR8fmdlp5G1hh/EeLiOAV9a2NE8PVvNKUU+XlCeBLh19CuPyQJnk2
AEujhTGxmFv9Ofy5a3rKcmS0H84JM3w7Qy/gPQbVCXnNYI0VSw43Yl+4WXDQ
w/w81PofSJ7U3kEnyonW1NlrFZ24K8Ncb3BKzVzlpiGVbDp7jHvUr6m/gSd5
YhoybTeiAEs+BTqmhVZmTa2wPMZOmtyAGeo2HxDVR8A482Uk1aimrhjAuT85
59ghlg0/uKJpcQs+Hsr5Me1lPfQUbA1MfJoI+ScV4Fr4n1uL/sN+5BEcQeze
mDjbwWrwzclMUz9lW63OGjwa8PGgkxQwQP8QAO1sLWeFcoXkJi9eCenGKkgI
zotFCAJAd2mUQKi+tnwMknVMD5KO27ttfU1G6X39+lruSd1DFAWzXipESHa2
ZuV4mvsakz7264Z1ESkDVnqV7TEOj3Ayv7MZ8mxVUYyXmU3/IRxFMGVUYdWa
KVHa2xdQ5tvKuixCgdrh5a2+vkcgV/SCv8RUYyn0MA2jcqqbJPC3EJvAUijx
V+h9VxQAs5XJQQ9OGPupSJy6m5wZlpBui3pWyWMwo5VfF+6JzhwEtX0vQvOy
+tiTedh0sgx1gX2yf8jDGKZuGGu5O49UEUepElG90nZNg8zeMjcTyDuGxhwx
KpbnurEkegQsvbPUw46KvjB1qs1HARBH8e4f5LJAFjTZV0xc+Wjp02IVBgaQ
WBQMOkCILB90vAH3nLvPqxdnSt622fzRWmt2drtSkRCIs52DCgMkg07McIl6
5N3byfC2zKs15CG7TFyu+I8/gV31y4AjFMoxA/LitBArUPlr48j8GC+j0lrN
IiZwZ1djt1uvljbOX4/DtsiM3M/tzGjfzocTqxzXB4JWKF6kuqE2SYVvdIbD
xMpMXv29K//kfJepntq7JXMpQSE4wXptRuhGBUODKtNwP5zUEDUMlfZD9GyE
DZkzBasnt3gxQvyb0rwRsikNRDzpl6MIyO2rTkerGJmRxU2EClDHaLs4fE6x
A88bhiqjyUh2B+6OJ1xUTCkvEpqakSjIWxOQKhzby7sl1LFyYJG0iK+53TPB
56On2OWfFt399WlCa6tLYiGFQ/P+VwP+l/Hr7QGZtu+wZ0CZQYfWeHi8znKb
O2LnHZ9cT+FAf10C8AIDH2xkjrpae9nNcWwsrjI8DArdJFsiZFR8mCCdIH17
vMaV4PK40DFtxZ2CRg94Eoa6PZlJ5JotiJjc6NBGyN9WucdOl/XoiVClFqbD
lHGpaMAS0WSmJk9xpSS+YPlCdJow/lhkZYF0T3U9HedRqW/IQRvOU5ms4Pxb
cHpYiiVrJheASxlQ3fy6ECCYgqq/AnLzVEIjeoLzVNKZMCxQQFFGJZSdnpkC
9bMJlA9DjRldm2K9PogOnlEIq48tgjj5oGGlU+c4GUUjClQBoCV0EbP6KTtk
3WTMsQ0AjWUC9qfQEn6iegJKwZuWICdG5H98Nxnyxz6NkdXqrY27wZPsrMOo
Y4Whwkuakk9TYEgSbpuw75akO3GZXVsqdWV6p9wa8/7jefyHAK68qUUUEd/0
5q/PY8/9xvglSYvv1mZiKY831MbrDaXuZCvaPi84k7Ddtp3dAhiZcnPzn2pT
FrW/ZD0mvjuaUjVfw3tYZ1cQkdDzUTe9ik4RQH19tq1PcXhTQvB4OOlZccZ4
BlDc3CE5fL5hKE/rT32Ip6L9S0h8+bcL4YNovoAOm3VEezfnPtrrO5hJYKAQ
F9841x61GZeAzeoR/5xim4LHVF7ma8Fm7ydazHivflqv4Y9W8mQ9vdDSIbJ1
iYfMMBgPqyzS2DqKTutmoSoEEvI1sCc0f9V6j/aGUeeP8a03cZJT6cua2M3K
ywvK85Z37WwkWsnJYP7t0zgeJrIqqCyoOuCC/DimWfAZ6KJGActh2+MERPld
1f9VDn/3gCTE5lMEFW5hemYkGGy65YRgi+6m23cMv3Uk+Mt8NYyH4SRGHshl
nw32VQ7SKB9sNOc/TQAwFA4HCMkOLYBZdStxTwEBUGstcPwDKJ7M0ljFTgnO
gRoKSsgT5Uc+lmUpNBHWaVFuAps1U/1TBEzj4WErEEsOTOW2VKuzt+t1d96q
R5eAqp1Uuc9wpYmKDP4m+gSwe2500kSpPhOa7BT3IX4nigkokXJW+4VuuJga
seAtsvdAynrLAvzysw1OA9SzdXTXzTFEV+mJ7FmRMh2pB3RXLWRIZ6YeDw7m
2sh6In5XTgmwoWauXLdgTpsP33UZDgaQs7SUlsvd1+XM4ZwXkgoC5eteVA8T
1KchhRvHC8JVavquyBohwqdVAIYhDAohKFxJpa+GnPg1Ja3WZQXBCPJ1BAlZ
dimfih8DXU9yzkx0+CJ0UEgEqNlyiDIAtfZSvn5ziRFnTMVarUSQTgRmk4NS
YCOXCeHx+FS3VxS49CWfzSZfoUjgteBg85tBcIjMDkPSF63+FHAct+gKuOyQ
YPdFNqPriPXm3O/+CZTj6oXb/n8l13cKENPP9L3jbmO4j8M6r17GQbH8ihWW
7S54MXfGrea27OdWC+BB4Z9V43Oe6DKbOvbSgQiiFDSuHd3pHxwo2htbUtoM
gHMfadd9HdqWlDug9fF6s6ANKQhltBSHGTNso/X9mOXl7lESf1kdckkNMDjf
C7fT0jD5O+XVewZ9sBPCRjyjGZ7W/pqwjBu11MmjtDV/dJlBEA69ogchJL2y
xOGzik9bTLz6nz1DtFU3Y12t9rK94iB7PZqKiFWs/D7baLSF0G6q02sO1UUC
5vEjazHM3WYZf/zDSsz3TkD0EOKkJLWRCHQppKjmT8q5YaqyVMVB1Qj5pWVE
rRUYDP9jlY8QBRBTad77TBJPTEM8bGk6rGqFJ0tfiwgE6Mxa0KbA81lFOihA
DwVkYqvhBNL6fQ/mZ7ocLe3XN9myl2SLDldlz20nmwA0EkH5Shyd9t9kOIc8
zk1iS8Aa/zpWDYQZmHzaE/DTmXgW85PbQFeB2uDerfvX8igDxsYPDozkLPYY
7ClCUzdOq0j+WH1q4sSvs4pmIXBqH/DldbyZ0fU8HvaJ+31UgxbTaKEdL/4l
hchzilByw1ROb0T5eNdrnc/V0GIHVYWRC86G0Jf+u8nt6HOWBKEYaLWKNvJN
oRH9XMDLlCtlWUXSGeiTInqzgzWd/Vfwx1Me5jWz/eNoP1OzLVJvrXja3OPy
E3s1WzLcgOzdvFHf+1m9IJvTYNho6qQ9cmjhgFXev3D3QJ3Uz0XRc9/zLs0e
98B97hxkwuUWuennnsx8ny2QwSxyfrDNRfXzLVZPrAdWEmWwLzZVOClPj+v7
qzVSDod66gC3hhuUYZE8YTpi33eHu0W1O/KUKN2ywDE6VpClOD7UEjA0xpZi
QQwm9bNwvZT85JzlVifqCZlbIZR0RCPjeWttNHXmEG8nbWe36t7KI7hvkXjk
wICmzKbvEnhcW9QUTGFvnO44HgDp4ZvXX+sJk5KQT34Bujs/aCkiiBzP5RlL
kpQDEehuM6HjsG0rSZhivH50d8XDsfKVa7BgXc5T+NVRHEPq7JEhJewku3tm
5IVY0i3ddJ+Gy9gOSLc4+c0TWnE4uvlyfwHN6KBN76A9Gw4LK3eaBx18UaPJ
1c97X3CHDgL53jPAtP0QNeg3iy6cpqpHEEXlTAwhhVwck2K0XQ5tc/u8sN3C
ikaWZQ3blyzYU+zaWi9C6F493uf8fFeQEiwOLw1qREsKYX2/2Hu5QEWuWBKf
Qm5k/5XQdatj0cTS+9Pdxqd5ShRqcpbnFeRn56JUpaBgrwQa7AcmJtl7Yu7m
732iUTo291BiUQVkdm+oj58+N4NnKx3Aka0TWSGcCmNmrKMR1Rpor2IV08Qe
CL/acsWNVCG3XqYU/jEewemS5P3+1tnoomwg6Otyullj/R5hV6BNSLEFKBss
qua1EGpLb2Y8GJAQyfCrwInjdbJs9QMKbfzn9/++R24CmimzESnmp+UOpduK
laTq8NDDb5Lz46w/qOY7gocxVyQOm57lWuWOFYx5S2SrHqC0oiVNEUvjGc1J
g24/Hc9xTDN7b6bFR6ATizUJiHH2yyD+ItuYSCCMcv3UzWMJLVt08+1gBmw8
hlKL9syfEjnfqRsYxgiGWK6sG+37VxcynS84qaXcxsBYAGEVO9qDO14dQGbn
Shtsm5z0K9rrOwCIcwAaP6XBunp9/QgfCXq7sj6TsX9h+sbMy4izupC3uqlS
BQOMXt5HR8UWsuUxV5FssCmii4jyDOKTTRojXZvfVcdBe6u6psPA11Wg/r+/
Dp6yUP3uzSpVHONyMgmWowcSwtlGgJkWijtdFFDi7pIr/agwF0M2JyxkHT1Q
W66CkG6pgPyX/w7xleBufq/lmuAycSFfcoRyAt7nQk9jPZWR8YBDoYHtGAk0
e1iZaHoLoan/wUzriyobC18OVX0mvpRI31PZy8mhSNyBngz66NCH3CfBM+sS
xVMl1L+pTPjLF470IX5StKK2OBil1XezR5Nd3dx/PPVvTgFjl+OTUkPCCkyc
634fJWrJIornSROYxA4ofiJpy6lUFuB0o40PshRNFiO5rg1Auk6WRJBFDBKv
QLNFDKi5eL0O3Zb4ZJHjd6s+L/IZPWe8zFMWkb4C8WthdIC2AuhiHRufq/le
kFnaYjaLxM+ySsARD4n5Q2rAFPH8jijHyMU/7eP0yZSjnVXYHpn7sDfvwsTj
EL3QxJnB6LIWcXovJBZGVCoHyspiKvuJSSSmjlVM01wQbLBUrKbQkQxUjPag
baKnXnjeJC8PRFDEgKdZUKGccDEaYWqOiJp0Lr6A2r4k2B3ctuEVEClX7YIt
YA8KRyIGzto2wfeABcySubluEclAisEdeCvRUQRt03QfnL6Nv1QZsAp4ET5Y
Meallhg8bZnhzq33ugrP/VVHUc+nVrnyoBFpRlAhm2Uhfxc4QgHhC2BPytvC
YGjgmBwIiaxWy6GvtRnpue1Sw1wUlYbFQujvigBf2gFXOknMEcpXhiWWPvYh
+DuYFTJzgwD74mr1Tzd1XsarQyawEWkcoNq87+OuOPHfgrlV2Iw6rLF3viSV
jSdakQD4PG4AQO2Opx61QChOuAtlaVXpzahYiwPGF54K6ljUuHZGZ9RQVq3Q
AbnezAUJIhgMmyFGZuU5gejLmjtmoOEEa7WA41pn2vtLWgL0bUWPpyDsN+o7
Z90bjRo6Km5EG/cgq7Cx1O+zhpxZnxoaFEH5AgQYelMdItsA3SSfpianmORo
1Q8XprqMa7/DQLbRGo9yD2/9KVNSsUei84yJ0+W21X9B5GBUQDcjS3fHaUoJ
zS2fXS4pt07lU8vwl6D5WMV3Uq3NtUbedTD/bv6DbHeLAnJZjJBefGQ0Tq9F
qWwzT/jRod7GDsy7azuuJGnXvmQ3v8u4+meFUFvW3kSqzcETZp1OsnW/xvTq
fS+dUhovDiVKc6i8eKB8GK2OI70vEQjJ2q115Y/4iEJ594cxNgTEYy0Z3lb/
NZk9R42U4gc1vrenVf3sQVUUtiSq03W0GUZhelL1jy5Ufvq+P/cnO+o/WpKZ
Gnkrv+5weRjGbk8Lc/rdwLlGGQ7yRErd7Nzm06EBufP+jq7UrF8jNO3RBlFo
uoc4dUHMqQSvyN/U0e6XqLbmp4WrKCem++hPH70h/lP5ISp44Bd3Z+Fnkcw7
hMkZp7Rk8AKOfNqmh1Qqf2+XmWpqNJfefrwZF3kcLg0cY/wpoX6fVn/3PD5n
TI3ZMoTz87oZ140ssDPJj89aubbaJTU854Maq2oDBzsgrcBo57Iju/RXIWhv
mSwGcvHiQdACRA+MWAYegSud2QxtKz1uXaHoWWTkyrKVJIrya0OhPGcR6oFp
e7qWcPfor0cX2GdC54roYTRqpCrZztDmTaLQQJyalqGxMN3ZGiilZRLUJIa9
LjVJQFGR/J2iHi0FmSwfOAE3GVclkR0xrs0ONfhYHwBk/uCTCRZ74YyIgF5g
nCBOX2R6B1peMg8EqL8zE1bqJ6ot8SluRqhm65cHVEXqngyKMRiT8yaL3uOt
eEIv0/jErGHvSSlUKwNgeDxaWnHUuIZ7uCqge4ghVhhVV7u4wH6vRggsom89
J9z3GnfVAcUGu8bzdjvFnSdeYhmBr/jhjpo6PdTsSfcZhPzmAMnpA8giTB5D
GJij1eYkhh5Cd0Eg+ZhfPuDpQWtxALUuA/z6zckKxxJfX1fL9NJbEmIFcEWd
d09p5MebhmO1OXSg/PkzygOEzkLlEL3Z3jW3F2Ldepsyn2sTRTPsKHdFuPUq
+3kVQ7NEKQxnl1xourT6bsTDImnln0quzAwBp+IlPCsJV+JlEIF2YupjHHSF
1C01UQEUcapAQe6O6B3GRlg2l1UaG9YOkMBmNBcykOHG0mZGLRGBxmU6uVxr
KEGL1cjdCtH65BBZbJB3uI+wXXsDSFsfRUEW+h/1R4NdOCpQRLQ8vUdbd+wf
+LsSZFlKhAVHWOeC93gCkIDLUhnE+1a5vWHY78ZjiZxgDc5sH1Oh97NjRZx2
0APbw/TozOaonv0rytwgo8Byn8uYzomLMh4My9xUWkh9jfrSnhz0uasIymp0
HXi6PMMdPSb3u3X/7mo+1IjuGUNPebi0P4PoPWlwDE52NqBIUVVslQ4pyiKO
8HbVMHXL8HXoYCkAFZckXXq4XVwlX15NxvHmV1ALmRAKDI2TvDZNZKqvM6Hn
WGRCIrieJ8lww19YU8BIko3IPVvUQYJcYvXJW93QDfObsLFLM/XWUpqhKGvW
PmL+nDhJHMGO75s6OHtrc5t2x7h0svqMKMI4Ii0BM7EicA+JHwUnjWZq1sSG
lMKACMXsCbDGWUS8dpI3K31DcQbzQ0rqELA3ic9819IvffJeNhgQ32s2Pcqu
MQ3sLm0CWdS9ZHgBXemgcEyFTK86wumeLXOBVA126OIDcdJRs46b0xG53MCp
+p4eDiazFE5FGwQ+E3yGCeYNAZJg2Tm5qENDuFmIMF8OXvdYZic2gqGHBWbN
r45bHewjCl3mcagdn1g7lFJkx+Cpaa6bjbBVEOAUuxppEI3x8tLRzZ5wsMNY
kzO5Uv+K1y8ywcUjsXRbcMj7V3sjO9ZgXM5kQSENVCpDIF2jCcOxbG7n+98x
NnkpM7M7YgqAQzvplV0qvmkcfF0sQhzgFeK2lUN1rf7va4C6098lB7KN3g9u
vsjCI1GRdhX7XVyJ3ARfaTHaPAJ9/VrXl6hRaiB7GcuWJ2cGJK0z2mJg4a6i
uHfHA0eHpici642qKXMFA3aqRkGAtHxohTLfHi0QLvxmbq41RXR2HPDoi1z+
cBOV1LoAS76bpHv0WkqKXFdmumZnoYrUU8z9jU0G81XQU0IE5BJJx+KPaJTz
dG7yZwpdy18PKg5QFyVtkdDcRJVeVg2/2N4fxHuPM9WQm7TBRsJPJafPu/UH
fwAisW0N0PM7qOZmthnHQJkitgKUx/HZq7HS23AcLRWY69eha/iAgw97SCK3
Rj6MJrU8DQRoEMzMzaGHgAB4j0KsTDThyKLpEgjYpaaLyWs2Eb0zPBdVFu28
M7aaaP/Mta/MG43pM3ANhwXEJwHFeyrCqqlkgtlvOTBAbXLwwqx7cEgY0+in
+9vLdcoWU4bh7GzZ57IhOviDIsDwxn1L94P1U74N

`pragma protect end_protected
