// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
T1uHlTWqcMMXvE5uIueZIA9O5ss2BkUDFqbgRVks1bVMA0DKDiQQr570vXZy
1LGEU/0zrEk2JIQW1kNqJR9BHncR14NTOp1rxBBx8c5ZAgkZGIBt1N8p6NCD
5ltWK/yAKdmgVcyC398Ws0Ux8oEiCdPmCdVWnHG7/i8XgSHkkjGfMUIHIhWX
FKZ/nkAs1ldx02MDC9v2BLFu534Co++Cj4VQS0rPQZA44vX3ww+g8NDdOeo+
zg/SJJykHQCNWK8/JJpud6edu6DxTkQBkTTtGerGxov3V/ukqazEsbCiz2Iq
v0evZv5MCjaf4VPbcvyY/PSfPAHK0oUqPhhiI4A78g==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
OxyncYZhRYGWyFJiqVzalfgqmHksxcOqo9kxOa0kmVxotStHrytqO2QqMlwK
LjNKAq3aOFqfJGTZmi63kHpnfjB5peEDYeMYfslxMjvxVzuZcvq4swmgVDf8
/u5CZlcd/+p4HkroKgMPj3TC/w3j/U1ycdLdENJTm30ge01sQ3q7p/Xt//Jl
el5O4G5urqD+XPS25zjKSoZp6uJBUjFnWOtAyt3tkunNQHxh3JLyLDiybrTP
QZ+ZpiEU6NSCUigol9E83C+F7nFO/QjC/DJYaAHqh3SwGcQ4yHWMdETBEEMv
NpcL7lPPMQoJHsl/6OzLvonf6kZ71DAXAyu6m3nDXQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pofT7wsgX6OUvcfS1ZokJkylE6VGgMaqTstZJnlQ990jJd35Vq0KD0uLDDPU
msL+reJjcI6z2bV/kpK07/lI8SY7TSEdY69KQOxGMyYB7mlfEi210sp98C7m
Yd2Jrt9AMV9R7A4FrgPcBQal7f2Vzwnu4b5DxIH5HbPR9cThtpS7yzvwVzWu
DXGbffi7FaYIB/a2EX5K9WVtwNiRZqgrkn0NqcE6L8kslBFSIUuPew3nzYKQ
46S4phto4yQmpN0Erpzw6Du5B3oDyV6MA4sJBrpqFoeatBhgoNpeLux5aITp
ppSky4uAxemhSiZYLBAUqN/T9DpLUoTI7sNIjtu4hQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Q16uic+Wen8R4IhWz9+WVsrtNegQQUKcDi3a47uMUpEN4tuil6bSsHtk+n2c
AgXcTWC/5AjAtHJBBznr94nlTdKefmCR+VB9Jwx8UZ0hek/asa5cdjKQDzhW
pkUbb+Av16vS8TR1uHZQHcWtncIopttdtSS5mpwSTXcXWwVVp3M=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
mUFv3rPmUlxblzdoO7jijR+QjWLta5u8wN4P7ogUW2OSRweTc5vbsXhre1QD
1IG7KwVenABir2TbrBm+d3ADF9wVNCEDUbjqWRjmlcfmLrBfI+cGfS2wJsof
yIyk2cjFCngbrMarNMwSUVqjhs4FHkjWWoka0tAldIjhdsnbDqMnK8KKxkCf
tN/injVxE6mWsWZnqSaPEsTiW7Bpg+Ws2R4SkFlkuuae069N+U6D961qEwzA
/G9esazj8PNQCRpcNUTqQn7PdVH5ACdK4JkJrsrEotP20NUvKOW7imkvdwqG
HSq9nEVVG4HslLEHpkHQ15YQLFMVzi25O1QxWHELen/O9AzjdPIlxxEz68RA
8TtzgkpsPoOYK6vIPoVctWjfkwcNXKyBbXPeTG4xkJE+CmbErYPGUOAd6BdA
IX0NoS5SSAKF+2usQfnMmLDgxZnWF6PEJIc1Gjn+oHq/auOxM96Bv0TQ6uUH
TmCrcfgITYz6vkscIm0Bkf5ETp8m4MIb


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
aIU7DPhCxhay2AwkWfDDbk31B+tBnjz5cCMZcT1AGFmpgfFuxaWHzgj12YzJ
aOiDhGRFqiG1x7stKNQi1ZKPoCgFbn/2G1nSd1+3dN+Qd6AE7AIxhLo31EFf
TXwe+bnKoBGkog3XYSfrK+SGG9FLA/lNO06jCPUi6PaImyNaqYw=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
A/GjEm4f8iAgkpFOtx1UrVkf6rhQ+2jYYmwN3FFO2rkQqKFDvKVpuEZtlKNq
mVADllnnz29VDyCK9PLDwofjy1zAnztMCzA6ibGtjWvI7eyP2JQh4O+6XVxN
S+lwfxLnFJJbIjoVFViUNiURRjvuA9QEuDL4CR+J3SgWtUEXQ9A=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 22880)
`pragma protect data_block
Qc/jWcmveEf94mz4qdsdsPnpmT76SDgID7HJhXXn5Ehfnsne6aLS4w3ctDx+
kNH6iBV6O/dDs7RwO9zG4Goi9ls9GKOp0YzunKF1mTmMv6v0L0OHiS8o9Q0t
djvtGVvdwEh/r6ByN7IongvwWCOPvvASqFl6PFv2ejT8pfR2oZCrbcwKpJBX
V8gqvBjNglzx7Mh8qrpLqP4RELB1al1t7XphbcxAukns+4JHiYaFnpzccMKB
FLyqSeES8AmeWnn77ieZAYQXuBhKGdxewonh/yetsYoLVQsHIyOPRbYY/K9M
pziAtrOZ7Ddf05KmXKo01W8JjdygNaeQoKcWyww2EBHPa7kwvv5sKXQakYub
WRBPFrcdHpDBNbBxtkhlneO6lWlkx0mnWVqStpXs2PrhRS1QmiXoT6pvzC9c
ADU7sz3Wzmugahdtwj+7U5FkG0SighO4csCEbmtBk4O/OE1/JDQvWHfd2LMA
kd6CS3wT8RVENS+t5Xfvqib2Ft/bSzNMosad+YuVZz9n1IYROrnCHOi1AtZ3
Nto1lhvnSUTFO2TECUmg8IAJDHxvHWOMbY4tVY5le+rCOq61KGw1fVR4BJZ/
qa4hRxpbqtOGviGiAVQa5sTyMfixmuSH/JlIUeoZ2rrVBLox9VJyjJfNz76W
xW0ishxYYU0OYGunT7FWf58Me1/EEijHr4PxOokYdTUVpXJCPWkf3etHpKUJ
hP18c0TaKlroDwOQSJRjv88JUy60LO5o6ePJyIaqYo3TGs+2lo7Yp7InpOK0
eHCQCyxO3eWYpgd356GPyZ392qjVSetpCDZqlMiPWOe5Cw2bbQyE+ceUOWlW
SBLajXFLsli44bc67qYTy4lZa8oj7FZdsnKRho5RXTfZb+4ske1e6s+9ldx9
vpufVtKjYYXmO/pyHOdwYIdOVyzlWsMnfEBbD/aVUMX2UiHr5009FiFa4ac0
Dt++vvMsq7QaiSoE4cr7AY1++oDq9I8If4nKfnLgbLi+ShJVnxBC74/uOvMN
a9HhMrZ7af2pAG5+kanHBc211uXSL3grKghrFd+XxRZYAthUb2ahqLIA8Ot0
ZPKKTjuyqR0u1lUK3aHB6Nyu1g7vQfrOaxwnh7b620oK6yxCURSMA8xpQ2ZW
79bwkIHaWv23kUn59WhTTppQlE61Q9zsdhAsPjuAzqlgj2igZ8bgoBbCeamS
a5lKPaSebENq03oZBMC2KXv2dN9Qmv+dwV45ra99tS9gypVJ+j1n7f2GuvoD
Hbg/JuD621D0po+QIDOojsSlYK612VMWrXQFIWDcHvcu+bFmjM3XgiqbMX7k
qaUXRr5YLSDNM89odUOJabrG5SOKcdOntKFNnyETDvnj8HRue4BxWSCz+LVX
LADv0rdKHs40te6+CZSyxk2IqTNC4pvrt7v7t9afF0Me0Pu0NRZ0LfsHlxwT
r/vDISeRNfXkqtpTKOVC3WNKQOyzZJxkwt8Xo+93WISY3J1xYIwK0fNwVlc9
/7R0XPX5+JZ3hfnSQqtUOpeb2rlGAGMNEML/4DrFL7RbGYYP2BOs8b2zZYZa
c8Ro2baf+h6S5sw7Hv1GiJgpCULqr7tMXH53dC7Vy5m+bOaGO0kHK3gAv5d2
vVdZCqbi0BbtNJsewRkfukB5s8gOPXbMGvSDpbkJC70pFtj2E0otTZoi1spu
QDcpzf9+JoX3jsrEBjWPIlY/sTYCVR4/heCHX1toxHKz7lzW9/uxfEOK72p5
LRNfEOT465QhnYtnXp1kDenDJRvfihthnVtavmDZ3GN7e3Q435tN/lPk5PCF
AmOcQ0mDhc7my5AFwOqRgYYdIPpZrWnuTR2hfDk/CGwc7ux2LFaeiw+/0wSq
3tSiP6yR6T514LWukPq8lz4LvimO+ce7wVTHiXg/isfQ98kj9cxyj0iWFm+c
BdF++EzuC8sXvugMGrPT2zsAKfuGtZwvQfBuMz8lMwknexPdcgPkacejitjq
gBu/rzMiRJn4zFsdf56Jh0ZiHs6esLALLBZge5jXFfOkhENB3Sp//TLTkcga
+hs8IiKi3yUrySfYUp/M5vMFr4Ib6g+LoNjm+la4OxCQn8nN8MDMA0za6Tp9
+OHmEhy5BsQSJAftyCA2UWQG6BFS1JfxGci4jOuK4R0EaEPskJhJUokxc57t
Mjb9mxMO+1NSbRyLCN2HsT/Y4W7YFAA4+FJZxOixSTbb4LSYQZbipxToNNMu
9Kl+njXXuNKjED8T8OUo7SEMeBrwRX+AlLnzP3lZu2pOGFkooeQ0WcZyM7le
Ch0Dnl+TWmreWwv32tXv8RSZ2t78XchxegHA/+ybBdXMJA6RpWFkEZ/JTuEf
z9wwDs0g/fvG1v56B1aIXUvpzusN/rJq6zy0N31RlvLG7KLDFuvOIS73PY+b
li9ZC6kFev2TToQL/s/eVacJMHOx+YBG+xMQIFw695L/e+MpV0xrqjzWcZor
aaAIZcu2LqT5LT4VFcRIcq4rGF9Q5P9lSRQFpNQjjyVbneycgX2M5n1hCuJr
c0EB6+QSOvO5w3z4H/Q+GTGN0VIWapScizUXVSOvb7kF7RCvkXraOFz0dAdo
JcVRPICUclUr7tHxX4YpdzHIKy/9Sy+/zqOI3oSjwJq7/OdNIJOVv7T+RKX5
ue7j0VFmjBwBSbvXvhYeO7iGtkADYTh3hIcMND8xaLJpNl8Snb34Pd4QmSGL
m+6bZRhuVOOwLtxVs96Bq6gSmWO4hntVckm0YhqNmJBTE3geAjnTexGBRbJp
CP900JPcdleaBscuoV6YuGbok2JZoElxIOg3F4QdpP6K15zm2JSkmaQAMLCH
48uN3y/tmUrzC1v8sfWQz7ZDI8e7pv680HiFPrJ4huVJ0QYXJjiTTB87jyad
f/NnbxzgKqeffseQLcDRm4AGaVDD7zyvl/TfwHG3rbp1niNlq48NWzNSlmrU
R0V9SJD7gh/UxvMhhCmC3yENzVAIw5kU9MYrVG7jd9SIsS92bpYb7JpT0e5c
ongfDJ+Xa4mUSN7vQu0HuyMvZDiiXSMVq8I889TFuTf8AtmFKsATH1vpQXsT
hm7Oxy+nx4w886aWs7PXFxIQspZRANqDLW5qlzXvT3mmwqwcbKAE9oJdQT+i
DuGSffR2CBoVkKgC2rMDdjGHaQnPMtDfWz4T3623/rnLlVK70ZvYAJZxfGOT
ew5NLJ5+t8d+daHPVJ99uiulnVxlKucOVpuNMwlhcVcMmIwzwhnFSHn1IdOZ
BmueeKEuFHxcHaHJ9YUJ19YZ91+r5e4/nHzQHI3LVnhw2FaeS4BzFcmbA70O
6rE9h96VQSCGQPOOzJpgLzkKWOfUzs8KzT71f0e7yyOsrmnE0ry9W5vXq/Qz
q2MFWSqP9RKjTezq5cgfYeihOw49tWhSRmlQ/tzJ93DzqB8/x0+cnW8qV2l6
lqML7c5bTHbcNoUpfVU3lkDZHFrKyT9EUjuyGIIFhRGU7Vk02wEkLAODoz3V
+JxJEdUe5elIKo6VvsNXnEVR1jQFTUIhJnfqMaKb9dLa2l6Bg77eO63kd16f
99MXhNSXrLpA+v+y48n2fPEnv8/dG3R9+2vuwofvxrKge2YTzV8GMtT93GdW
S43njtoLYpvX4rYv6s1BsoZVcINWCypDWzVirghscYDzVMlllkZihrDIWsYq
JW0+/Ls+GwYnHhXzuyeAZGmOZUDCnaCbXvcobC/A8VggLfg6QhzCr+Atp0wF
l5xjpj9p0RSpKcHdZ4Ei7GwOAyNJOtbsLsZKMT5AJUAcs+9gzBI2slKs080y
BlomLmbXZ1rImvfS6pEU0sB4fAccrrgq+fe62oiJeuUG7ccl2MEtThljCsCK
DPKKGnwKt2n8tOdqXczlf5R2lOLn4UwdWZETABpa9ts94ss1rpqPOpsCJuBP
ru8KVmxByoEw2S51j3tDTodAXLzjvXqreyx36lBZa9mH46cwe0u3WR5r5KPr
qMEaBBMsqNuA5DSOmew9CAWxErHPG7c/hWhFdaRU+E3XP9CdoFBm5edhXdPv
h7wXKAc48fVcTi3t5oVncSHAycuwrhcQHn5FV8NjkhPvQx4WTOT/Kr89kujm
FxdOH6P6DMrqiLeRh1B2jqBrWc3YD3NJxnbZo0L35/QlWXQg4VzlpQ1+IqFu
F9J3a8NA17sXkogLqbFLJhf8HaxR8ewMfiVmXL6r/ntJ1EEWbmWg+OPC4Sd/
R4vM4xA2zdM6VAZXXU7OJDSVlbdMf1EsB0LS57eHsm4laQ4OKDMEaL0n5q4D
C8gdP1hWTlMzV1+8ipwAaiDaaUROeXZuNmVOWklKheHqm94rpmCzJS5VYH15
sv9rQG7LPnVzWgZ0bF0C8CLzZqiM02KFBg4v1yBS1QetC2oiNwG88lAG4WsX
HV0sXJi8fCpZMBlTb9RCwaf5OWOy4EQKx7jTYHC4RT15kTa+hFVLImFopgC+
ejYEp7xawmz/4NT1C0cgx7bq15Z5VD7Z1RpkJ8QViwQm+gWtRIoeQA11VL5Y
PYgc/nPRsK6zAmfhBwyQNOjQ080hqQ0pyr1sM2lfXyPfhFqYYYLk1iqW7vAp
x9IpanMZXKKvwgU4eNsbkD8eIgwndsn7Q16YUKGNYGr6PyvnXgFTaO/wuCm1
rgA9NkSsaE9/vU6P37LF6XgyPTuH2MyCHHDi37026DJDfBD8ow9p0hSiDDJ5
gVVQXpIpn+mF5iKwwBvopi3qwCbxS3G4FTL0VM8Wew+Zqp87Edvt+d7tt780
IuJW5ExeAdkntRg3mUpTnssT3rfc3JrN99kRcwwTfSUx/OR8NueKyeGatB7r
x4yEdzQ0D1NTzp565ToajyzGE1QolarlcmDcDeu9tZXU5AgZz/ug0RXBolHT
PRph3bSMiu3DzyqYMz5QoMnTGYiBJJ60WB+G2PkJGeOGA6ffapw7HnqUvmDz
6y2fKINGnpUdgFf9GXyOhZktGWT63s4Iq6e6yuIMY5a3goOwBJ2XnG37Qhro
W9A2qALyT0AaT6cd3q+uO1WPon9CecfMVNiqM68WBUkBoayMdmnWhZbMnz4/
9VxY3hQ9rS8iwj3NnfgY/8weg6VPcrJl3hxeYqkwsxpKMFAT0nrQMJJx7SF+
vyCCGtoY6d+Bv1/OIqbBdr54tp6j7099tCbw9ahXvk5O10JvVOn37e0ib7J/
745uVmniIz28s9YVB5Xq1/0GADkJqdVpTMSBBzcPBYeaTjEaSrLjHmk6jnop
vaxHJwK3kuaDDBENEhrvyZJT6SP3qQ+qVLl9miAC72XMLMh+hXme8i+QwRCt
TFY7j+KjUP6GKhonNXjivBoj7JKS0J4gFOUTkwhyZ/M2l/NIBbeAFAUmRqrc
LP0PrfCA/Epwetm5ExmCty0hi5w43OTuIwyeFhoiF84zp5TTojni1WoxfWYd
yIKyOfC/pQisA/voTv0ipaBqMc1xtRmtha+zZnxpaYySYM/GnJKLpAGttI+k
AQ3sgeTiljiZQUJI+UfGLyJ/Ux+xVxL7N8qs1nTyKycd0ZpPwMeaUGN5PY6S
41LiIr4XIA2ookp+H3WD/5ZrgAxw6BZVsVeftUS0qKUC0M48tmxz9dfj2VBg
qhC9ND7EgQo5T+Rike4jxacnlyBYZwiNq5Ukxeiz6HicCu3c69ZehjDUqsIR
EzaHkddyjFugIoZZ7jiDNpuTKaLAJD7Mit8gdJBSaLbGr+ilNJ10NwRLsK2U
BoBzzunE/FHlxBzWCmUN+lP4bWvLVfEuNvrl3UG8qSOf1N+ZnTkLlTo7QLbP
4KCTCZUe71YALOL4xMZFaA6L49pjk0tzllR3+OhPViAs7pWtiWXUmY0T3wop
6txql3CW3OLmVgq+0qWX5bVUj8WGPO9Xtt7PH6cpyVDCfzhlFrUPEhNjkVvn
Oea4iN24lBjy/x6Hev9rQtpujAvu5/1SxbhtJW8uybjNQnwB/ZmPwPBHQIo0
zGDnNwy45TM1kehw6dhk6KHsK+pFsUXx4pwpNdZPVwIxBc0QjiQpFh797oyy
fp5+ZJNRaKss/xvQ2Eua5WHpzfamH//uwAGpkbY/YtJQIC6pEWmlsdOfYK1N
xyhezlI6K9LFA/VzivVUhU4NqTom/A7pv3hPkFYI9WJac0Br8E0dN6Wz8EhN
b20ZzvHrKL0vnswnMfYlNfF6BqW4yk34ZgcWxhY0RNX5e7ztL0Fn4n65QUkn
2pfsJ348UDZbxdAdY52phZOLTdJZLAj7njm4RVf9zs1Xf+6HQWfMTgidMr5p
Tf5/oSLx/fLz1ksS3fGuztvJA3z6WBPE2M+jtpDPZwc0dTeV5FapKm26WoEd
YpIZTCId4254vJecC76A3iCEstij0K/bhkovDiULx5GrdUn1nli0QGLhjBN+
0UGTBQ9qY+C799ExR/n4iS7jR6BE1m7o9nY3LyW/CdDTlbbjIdj3SQGHDX+8
Hq95j3/PwYdV9p0sSi3eLWtAfP8LjRB24MFrWpAPFI5iWDUUjTKzbehq7l3i
0L3G406ksOfNJSEWvlg2a8CpgUkPO/7gihyDz+g+zOXsrCPX+BPe2L0PdgQF
3xjEnzzkLE7m8HpGadXaYe6P2QaQESm+i+bXv/3VGT3DFhvpKWPhvLzAilcj
u5JeRarWtvz+w8ArsbCcrAJAFNlaC7zAJmfwiFHFB33XkWP8Tj1niGAU4rJ0
luy2uMFF0W8kLWDY7rP3VyJI8hpdGjnvVH7whJdo61/Y5Y2izI4vX0nqhuIp
zOt5QaOeb/N9h1GioB1SWiXfGSe4CbWvZZ6nuQlxiyqealC5sOmRUKObklp/
YWmBlrOOCCrPkAaei8C+jvtcbF0NsGJWvs/Ikp4nUKxYQIwl9A4oaOcCC2lv
SVrwWT8WzqdqAtCd0E06oyXFeNfID2wh9T37D8Kx5UKXm9/S+DIfdjW0P8Lj
vzwSM2ZNb20mDTQScqQbLCXHVo0b90XXRsXPdCgFnD3raTY37HcSzDdU0T2U
qUg7ILPf/O4i2v5LjqayoM4DsrKyE7Ds8sjAMn/DzAfo0Ta/riIVPcS6ILUP
EbZERMwUq0hcls7Y+WQcLz6grCP4uHiSGlLceLlB49q7aEpuNcJqgcBz7YbG
X3CC4IWQ2rsRzNYE/9EnjUsvebsUfRfZrlfxv0BlvCeOl7i7lrkfPdWtaNq8
45XZl9yBDAwGK7lgSbd7H2EkV+PszinfuKU5OJSGpgC34AutwQP7e6K0aH4m
eNEoefGuPqR1XnyZN0xvaJr1vI6SsK8JZGjsKf0Yetl6BP2I1UegNBeL04ba
XQJFbqa7q2qmU2Ni3fpKPWfa7nIsmfEVl4vS7kC41d2FkfXetoEa8qG9K+3H
i06MdAVPTYshNYJ2dnRNJF61XU8QY475i+2CZ9Ye9S/MhbzT1C8bqLytMScT
RAy8Vjp9b4eIYxRLbR0+t3oqIBav82scfBH69vBM1fJdy9LVDhwxkcGfYCmp
HpHIO29FgZOLAcglDZaJAALwFqtaprojdB0hRPKcJ1k6jm0Xj3Co38SHQIav
y1QE0BBGXL7q3o3TjPuuF+9SKDQnSc5kmAEkKj9koYe8nbLuIYf1XXLggf/5
wBstbqcM7rSb2WB7MYeeMphD3bLU7J4hrsrW/eTW6cqLGTgAPKbbyFHGabAp
K8E2Ax60FtMAxDIRGRtGdypxe7BMpizk9zJkpcJIjxwC0xCL98a+uXUsk4Iy
mrjQgKIaRJot+TVqe2A1sDdE05TzE4JEZh5o6abvD/zHG59YAYZo6Wu6qdSZ
HOOQvOkSFFPwmR22NpeYhJ9OiAiIX5ndXmRiZAY4gGlMChp7EKkZIdR1LJ+0
E9KORgsnHhZCiUWIKKna68HeeHGVMoy+DFC5oNFYHRzW8zeCJ1rqEV28xAFR
UTjtKT8VN4pimobhC/FyMUwStI0IQxroCHNXlUzy52USakBSwfwsVrQ6aTrq
4MxwLGxnkH0iqFIqv0F9WSOHzvhdXClWg7nvF22BeXG405jRBUcBREDhBc5o
Hd30NRJyYH//zoGJ3vweOP+bTxdfgiDvyNoEuUn24FyNzqrARoV1gcqHoSPP
/wCb2QfaP1orcZGaZMTf1AcjsVPiDYYzsxCG5hWYXsKMP7qardDM0UNXWVla
OcH1q6TyBVcomZahYXPI1g6uMmeUuIS57O5JELnCWo8s/DWqKDbL9b8EZ3zl
Ay2Fe+/R3wR3p91MnY7teRkay3zsjG/WA/G//Y7gv09j0K9VvhmdwQM1p5SJ
Mn5Aj2xL4Xi0UDKA9c8YHpJjQkHBzpzYEl8S0ZI6jmfdQVoi2ZT8i//pf8An
M3z1hLfF0rvn2k1eNfpQxc33nsLR6KMEnol9WlKWA40JZQi2T45yo9d9+Ibo
DxtLx+WqPexyYkbDfyNNuZgUaIomzb0nbAKICUakvatA1jJkUeVhIf1E6WXm
Z7L7i+trhfcaJoGjY+pcILT7IO0Ei16+ASr1lCY3pSHloJGB/mrbdSwkm0g6
nOF5frEV4/wWZ1DobM0IbwkxQ3rFhWESvrp/Dv7yGOoZihnjhhFi9VVQLsOt
yIZd4Clqwdec9tt6VeJMUA+CDFDl/JTX6UcSrLGS1dm+StZbQ+hzD/zyenk9
N7uQV9yHkBsay+r6feeGzu+ClqJzavYnoVa393BlrSDM2z8pOzbHnxj4feUK
rYr7z1gZzAkLv3otblfYlGJFc3Nq1XCwjK1Jxqd3jcoZLDGW02+LTROzAAZH
WOE+GfQuGfr2oyrXM5ztybF+GrPws9dwRo0uqQJvO++tFEEFsJvxgwTP/Jto
Hs7IUeywqHqPFOEubkvNZPYywrqdmKElD25y/Lkq91IQWfekmYUbV9mMBtah
C6K25Qzl2GSp7AS0evhBRGjeHLUzbsmyXNyfZBNX6db0Ta2o0qLbzde8Z0xT
Pc1aBjnxyro3GVdEADUG0LknhO3rswg5gsUaXiomVpvk1X1ilV+V3W4NyZxd
hzhA2il93WUKC0StiC6QIMFLIBdw4RaOBlxmA1SdMrccKEgkSQ9mIaWjSWAN
D0BoBOzJzNfGLHfMpl0fK9AXeIMVHCG1Ca5a4r+FCa55emcJu7cOScTla03T
mamSH+t0ZM3MENBP3ow/Qk22ydbqIBtzprSJKdS7LTeKZeAVvLFF561o1GV7
GwxT/eCIJa56vrrjMzQcCXqJf45hfOYoqrNxEu+vdnWdhzMnGv9wOK1n538R
ZTttPqrCFPfa+QHWOHWzF9GWY0zBL/sH6lRT8FXztlX/AX+NDlJ9VzOIoYBS
xaUeJMY54r38PcB4ZOVpeOoahOZlov8mL9F7wiH0GTMLvRN3D/cQeufj0Lzc
dhIY50l1lh1ad1L6Kaopgiobon2vun9q1/geqb1xRYq84IPow0oVrRCZaBTr
+2skFB9KYRugwcy7s/HQgshdzw+5onwNGqUk0E0mqA3zOuNHNCXZamAgD2ZD
ilvl/4/3oI5LbHrtyHtisyo3eL2huuxAbZPY0uimVusD5bkcnTlQ7CjzVDQM
oAaicLdgB0WXH33JYp+sLUA5tHoxxz5SuosQWbhJXXu6KM1Cw4vxc+nNB1G/
xvu/NCaxrdD2hn1+UK+/e+Bw4gTAJzIXpyCN8c8Itrs/c8go/Lgk5R1+8+Jj
jqfDiqTxkDK6hBSMLk4kG+m0tqprc7VEqp2m5c9kqdM12OJCxnBVu9hxYs/J
6/lKfPrWC+oT7DLRRffechjI/JHFh8aAtFckaj2YLQY6ji5nC9OIhAOQOdNI
5Qq0kbpXaxVbZQE6tkorCX/zaHhCuGVJgERhItOrRGwM05/Eje10C1kQDoQc
avDeWud4UBVODrzzaX75c1CZpUSU9snkgH0u50ZPw4q3KEzqts/EbCOAa9Vt
lTjVnphyR/eTq/j410oSGmQcVEB2uSTDZM7fiKrkZyu4aQo9WqNLEnjzMg7M
brAGnF5zz7pMG+hn01TiNLWuZYZPzhUM2txMKl6/1a+Ye8aq7WSjJUe5mnvW
YRdZ82pQMX7d3xOHVQAwLr6cz/1/3bIALUnu/nAO2uG/lpa2MLTJuConMFyE
iYIJ4KRb2t455evQ8iVbn33Ouex4q9kQTHYDu4TYYNDw1UaxWotWGwXqLi4b
yBjNU81IbW/Agh13vbpp5BsZLNBlBEbF5zexeNp86nZVxHdSmHzTamFzySEY
f2uzVNnDDsXv64HIwC7+Ct41n38oy452Kl/PrYNsUGC6dKihxaEhrIuWk+2q
+FxbrWr0TzTl5dL9LxPnZeKDtv2RI2DZV8FVhTIgtjkA/1o4ogWTwGjIxYUh
J8jYLf80iXidSA2yoHOClrY18bl1k38JlW4us0s3S9Jigg+drFdQbYpipshT
zh0MKA7sBmuboql6hHXt35n6bnN2759qEL72vPEoszFuLGNM3kQb3kJULV5X
vQTh+g5AM96zbjAtbQfMX1mt56jjwPcjcGr0B94WNzCNgrcs8aslInuoZ851
7tXh2DTtz7kqXyGtNnjJkvrNJ1LbExqLxE4AHwX1xGf7ctWg8CsC3ni0Y2Rz
y7vpf5QkCFrNHRvpgLO6TqRjcqypXxGLMjMPJaF/rOqTwaOM6tKep2hvDNgH
u7XjwgmTnD9MmWlTKa3q0+xh1C40sZ1u7I5ma8WI5Dmi2fHD3/fb62CcLpQD
/m8HTVWFVa1LnAMDLUy1UyRnY6ekz2TE0o+OBD1uvFAx0l1IMRR9Kf/EjkTd
8b6wrPYYMbTqca8ngeBOuGBWyNb39TfCNMh9cIxYTvxoIQy6/ZRhAgzBXEMB
w1C1AsH2ptxFIEbhfCY1AzCSSGGJ0tQEi+w8pO8K27dPSRDScJJqFJs49MwW
jH+uL/o6qtGzsYk5Ko08jDQ8BTJH/eD2G22+1pAwxUGXUjR7eH6m19zc4Dga
D4SLUs+fRaITltMv4oz6B06aCpQAeileACfHm2fuh/W6gYPZCrU3QdUU3Ha7
YR+R6Y4pFrSeq8Z1W8jiOgoNrWfDTjtlx+QguQwobxuwJUMgxMiCf7FlWoO/
keb+0eNp3jp1r5P5IfiO1R5mcuxevAmlrgo3EM6O7zLpb4pDQFfqNHG5RE2I
CHIA7EOW6SkAQr+A6Vi1wlXdKWh1DJEPN2XB0Iv8WZDhCHzVtC9C1dTaBN58
Oq5BAfZQjGWoQgifUdRkxJwiGkKEpvT5LYdxgvk/L0b9IfUQmBfHolcQ4pRv
WQasIDOwI8vIvmH3stajShIcA5uCGDGV1p76LJLPb/lgRbUA2aSc7mEwUmFA
Tcf4bwWzh3KYlCkFSlVZ3C7lgrIfyZMF+Pt7iYEunser7Ut1S/bT1n03patX
9E6WgjPPteiiQxtzie6dBZ/8yV6Atpkcn2TG9t/ykK9f9OASmCNRtS+mskfs
l6D5qr3ns9YwLGcT61kbxtM9QxILAqU3yKWugCP8clopmWJ2yQNwSEABomfv
xyJHrWDtQJdKD4tewXsOsEW4eD/eXgIXzQfK0doNtEyPlHQuE2mb8VLGOGJl
v4WfnOS6rOwfMom/9pjyKKYgDayXKoJQuaWch6/uxkSnZ9KXQoZXQ+awXMJw
mMiBjmsueo5N9vqTemxD3R+r3tDoI37wGdVCoQJS6pmqgd8QuefjPQ/hQWbs
GP++R/QNqJxxHPuoeonpz1Q3zvHbZGEEQcV0uL5rLiihJmdOxzfEVIToJ4Qx
RSXL/GEne3+7UvdQJ7NCIi6ujMOHeOPUL6Fgcwkz++i5mRu/EbK7YvKOnC/W
XtTJKBd+SSzmi64FDuDl8wBMLN4uPvqjiz5efSGSIKcWfH6W9CedNrr5dKrh
CpkjefLqacWlIcUtWW6XWDGLHXctcXczarC+8r7kpmkknh8tbM1IzJiLVt+i
ciDyuTj9RaGbO3oZ/G6qs6NFdyk60lj0Qqi/JxtHV2qY/diIYiE893OvWJVR
eVitM9zRUNsPB07u7bWVu3OG19HwERS6zT1GTsJChVd9q8cNJd9J1psfSGwg
9z9ZoGibnFiuQJXkmo0frWwf5g46w7IUOoXq9LOJe5ANgwyCxc90oAti4dYK
6+nvKJFMJFVCjU0Wbnu881bHh5rFbTOTQ6MQI4Q/hySUxGFnxrNkxZt8jp35
DyycDrHjG1FAs0gh8JqXHPRzlO2B7borv22M/BcuvV3bX+1HdqLeRnxxjbeX
spU2e3PZCDQBrx+u4baLihzTqmkbdKRWS4U10FsXJ1R+0K5oKm3T9D5ysl+P
Dbdjj5FCf3PC119VPpBv0Kv5CiA066r1RD1GwHCQINAtxnkqszDlbrzAAhhb
mzXd0oEPOeE0g8fqmAGt98d4sSfry8D6sAOC1768fgGqg84q17cqLgI3Lsun
26a8mz0y/RfW6+yHnQxDwxe1ruO4oZukYftqHlFkA6SSzAJSNAy6agURmVuU
B3nAbIFHoxw8ZE2QfCkCqT1Pzl3BUUeU86Zw1I+5vNhIQ5bExzJWm+YuK9jp
X+xeFBbes0txhc4lg5M5eLMHr5msLcVF+7SbsGEXj3P13kYsS3f7v3Ose5sG
4pEBXZ8KVAl14wfaxA81tKVh9fAWlOfaawabJKtub/r9JTADowSNAkpTS4jC
r8yK2A42e5E9jitoie+ptjRW8FLzQYJzTMfOXjIjkUsLNjZhtD2mLF3LL1iW
HoyDWQsKSbmnVO9wdFofTzBywLfcNTXCcCyoMgMfjjsXG1Szw70N6Mp1e9Nd
VHw2qyfVsDZ88StM9R+St6iiMZneP25L9xqzAsro35uLLAvR+HFk94tWs7MB
enOJqMBngbMbfrnEh8KZaSiXIrx73ZW22UKKqkjSTFQbn3TejvqSsRNs/l0K
Bj1LfV1QHLq7Mb2+T0he1kO2f3+3XzAyHLk/foIe7vkBOvz0MXZfJtaLq2bE
RJLvVbih/UrBfu7S9rvkiTBOqW8Y5bWEU+w0urGCxrG+5zkHAH1G9B4fPkeG
iLwORrdsDrGkKGI52TdAEB2spiVEt2kIIYJzF7y/eho8sj5rl2rMuEPWJUDP
kI8e8uUSGuCTt8iXJKUHzQ8t9DfMDoML/Zm7ApjyvpVWsKaREps8TxRGLxWA
Z0ljjfKI9omwdQHqjS6ks8pBGwszH7NVbNhAg8KYB7NRYpVOfyIKyEXSYBvi
i/T0qNWUfWKNLCWz++WuTimHp+XAKWDl9RFFR0ambc2Rr+A0kFvE4ICt2QS7
4pxo/AIDSa0BkxCWpD3bviFBYC1wsTgbRJLnKNSo6lmsG3PP6e12L90nSA17
xwJQ1pnXhorwgwzR+NzycZFP9CEd88F7ovo11+L9lZLafcQMYLaqdyiSPHAv
nvtTbfbY/oAzrWJGZpdtIzQfstU1aoZjDkFOYS2iMp8BVauhkLEhKnaIcxAP
aoNQv0z/aDZHxthVEedakmSF4FyEPH2Gd28KhCh3Tq7g7LgeRYtCZUOFkEJt
fWeo2HNRhnWJi3+bFDDpAu+4D9Ex1tk5LPqIR17wLqGDRjC3GUpQVupQqWSY
UuMchEpnDTJk7vkgoP6i8itgpk2bH+ViRpBQiV56TVhbM316lGH2JK1MjQ3P
7J1aK4ddiEn3S4shXYp2hXRzJc/LZr8JI6jZss36xNv8Fhzb5kH3nbP7Bn5d
LzPo7BbwT8vvq4rzSCcEd8U4AzigmJ/yQANIH9ZTaGv+3sWURoFGMa9sq9CO
qaWDv/49299Xfh8beHTVLA9jt0Hs8WW9dOc/RJUejmr1v2vZk90hLLdgkAKV
ytBJ+WmRF20QGU9Z7bF+7DuAznUUanLvld+NnqIAfKgmXjCBt+m86KcNZYLk
SVVqtTt1MEUY2PnABtDw8LoCjcoA0iqdbfdNg+1/RiM19qhO6jgBA6FEpupd
mjxjDyPfkU9pH7JYdL3IbxGOfKyAAsSh7M/gMx49p47qV05POeYexruB9zdR
nwMlUCmjC/BlQQ9NxMIGtuWfpIVF23cuQzBMM+3MOtxfGDDLDj18DrJXENM5
zPO6/VQq5LK/p9+wCgQERC63+VXswbl6yzZvgunILPXEEabi4PHHZmWUYKhW
mNPUskpAiYh/dPTYemBswoYGIYjieroHpU4v+3wayDSmEjEZjzP/DQ47tG98
92ABBDYWcwEUIcV0As8l5uPZN3zqAc+gzOLzoNRDn4YHT9G2D9OASauaqeUR
aO4a4zMakWb/3AuOTfqdLNVqS3ygHaAh+RTqBHsGQQjbsarw1uSDt4aU6KCU
eRTA7+AwRv233XcXNNpoVbNi0A+8rOh/9evZtRjDFWMkWhri9zE268pxe2II
UgGcJ685vjruclQpBbZGoeuyM7YnKOXB4F2S77HR/p1BLSUOaMEp8oB8LZdX
yBp9j9izNZtvFeSjN7sqXuYDqK2lh6QVp5lPTfKRmY1capC2HFXzzk/cTWrm
A82yMA1TPKUvRc/smSGKpLhkXiQ5OVZ80s8yW768B09IOlAIO3wYniKZNnoq
xBB3H7Fc91S4JmRbB1fFru1+XA1C+GuR0IQXSJY8uqm/sgzTJaAIsWDNKzG+
Fk3/aw8Gzw89qLrkQ07DplmAuFtpADY8Awt1VgELHO6+9VtIVbtaQX+oN0BP
DwQEZTc1P4rTYC6TH4f7VGA0+0jhFANmOr587XaIo169vTrf1vzSGOdrJ2kf
GOY8Q7pKMFjO3GxsWC0NQWx1DXdb/qMFY2JQjYT+MhXyQ6HQvsBFNIGSPZFc
0mBUcgaivNxLfm0zrgCDKVGD9pQnq5O2usKk7imcfnsgHlUWu6qNvAvk5kz+
xGrumZNkTWIukcCJDinAxtMqDsftLmJHqzkzpOPqbi51RZAQEQof36Sr/8Eu
cP4Bopi3WPM0dykNg2HeUvgyCJtxP1rnZWwJsY0beU8eD8fCiPVfcoudjy19
8Vac6JBuAwQXJs8Wf18jv5nbRC5M+0LmKU/uYC/+Lwaxiz4WVz29QTJJMAj2
koYWWmP43lOzk2naW/WEU1n5sda9/KoxKJBVJnmuPQLnqd6kn/18gJyJMaQU
thi/Bbh2AgS3W/FIj1IvyzoFlJYsMme2O/7y2Su0/TiIQrIW+uwWW9dv/NIW
HMYXRPjLpx0RUUYsqegY7QneSbkQd9G9EHWnLkpJnWvR+PSXVtsFxyRiy6Yo
bcWgee/2evFhD7dLFL4ZHTDBEC3BaMNRJj9i3z/Q8SvLcBnquEM0pC7dSNnF
gXBMj6ckKC5bHztdLSkxJUT8uqLa3PA4TIKFfR+3TUQKGlveAkXspPICj9LB
yGUiumdmLLbVywv+pIG9dukNOHxjO+nf49tV3K3TG+92QZKE2S/YUBtvUo3t
mfXF59BbRJq/Hl/I9/K5qkmEKzyqtZJvPRLWQWujUmFFX6jVPnZgbKkzsbKQ
WqXwBCi53wAUufOkan3L/8+kbvBVNgHiKV333brDxUBAk9GfMnqXcucmxq18
i8rivrwkq0cW4UUnxahvCzm5zmaN/EmMf+YeiBuObBg+jdPBYfO52aMi7iA1
Q6hUJr/Nk/vpe9CiN+rD/7EQC3Xa9fwjL1DzSot14TH7P/nKjtS8mKwgt6k9
SCJYpzz3E+EY0ROyY1lRZ74hnMasQ3bQq9Mk8kNcPEc4iPHJeJjWARgo3AdW
L+X5MIbVDjdo1NypFMhXKS9kAN05IQz5lhQWOYRyW7C8dW0CvQ5ZnT3yRPuw
rls0ZqQine3qaD1K4vrWcrXTnH9Mkih+4Rw1fyfJ4uyW5j1IONbykstwzSTi
A74QRoGjmXfO4Bq2liWcoxmCdGMNwfA2EitQHnXG2g4qWfif419iLIPKnbLx
VQ4/0uygxYf7aLM3FH5lrJOXqpy4Lw3+NY8ia9IzdeU/giH78Ro7ZHdP9c8x
1A2GDyw5opeqJVrkH1FrrMjEZM/KWbtjtR1EL3ijqcUqq3onTEpkiYkCh8RC
7d2GJFB6Q/5SSEGn63XNzeYBV0jqeVsfqqPfABmz6xfvSnsFmoOwsXM8LaTE
jeplJ4My0DJjRHMUNHTiA4Vj2/UtgTs2glE6Gdn7ow6n946MI8mJd3kl11Vw
RhG5+8kqgUWYOIBNosFWrHecFQLrEPs/ysM+7kJsyD4KO1hFrMWVYahMVvBe
T4QvcaPi6PWaEnPxf23EAxdV+2zoKTdItwQ3osXXk5BKM9VjVjAYXAJ+D+or
jrPapbBLvYD9yBf3zPUNDLAQMLjnU8DiQtFeAOAmjqGxknJWv2RDDQnnE/I7
XpNOJCSePtVg0FoQQqvbKlADb30WfdvXRiujY2tE3yXmh6bYyXReaN1FexUy
J++nWj7SYpTyMWEfBTv45CcwS4PD6ddhZEZ0L42/Iha6s2XDrj2FHnS34gNl
q0vtVc/0f9Id4/OgPaPMrXTBRfVJRZS6uGYhe5QaGOygTHbIII3WmtJ+YwC9
BmD20byErSGWsTFkpSjIYj3v7HRhuUklOCMog7ky0ADSejYCZsrcWTSTL4t0
xPS+D/Mcyn5Lp0++zlvNQDYQg1Yc9trv/HAsoTzTpZApwhKgPOT6tMq4/il7
gn8OUq+WfZ31d2WfiHePxXBowa75tRbA58pCY03euF9siLA/nnwamjmANCA6
bT+CzLFzQ++zdrcaKiVYqTxzJIHFjEKLKvkAf+YNgnI1adT3EFW66RpxWLs9
k5ExOJh0TgfDhZqQGtwEMAC06akv/8FETGfx9Uz48R8+0KR0VoulLgRSN12e
9op0feIM9z62Py9mXpQ+1iwZA35L9aW83eY0rrfd/ApzIEMxR9oSsyM1u7xH
ib3PVb5wAs6IGbMCaTi2ABNacRIhAEazoy8m0GoLNlTXadbqdP3DHEEOTwcw
ZXx9irGt16UkmePCwAK/4l5cz6vtzAp6W+a4nWm1SA/Bqw0iFrmwqzAFb/oH
uoK+YacLH2CieGtKyx5M+XOzw/rR9BBBcDpwvkCFPdQXrhwHtG9A5MAdirID
4EQSjtFtohbEwKFUXbKg3GFW8E/YyHM/ivakoz4tK+Hwmo+SQq2W21BtT+oo
LSpQ3oh38xxO+bhiv6VnaiCQEKfsYJa5/QQ9IptYo1yCk7we8dCH2UYNzTDa
6VyHQZ/BJ3C7VNmXsPbPgt4xpzeKnUpwdesGsy/tECmWnmRfEUk5V/P8D5du
jFEbLuzdEUUhOwtSJagZTvnKbbOqFtU2bKnI5Yht+zBk4u8pSLuRr85iA7E+
14qvyVj+LCF68Z+whk/ND8veQqwElMGI5v8/YBlNsqsc9qkqVjouWIHGqMi1
iJvWDFmYYLJfUwmI4JWbjvwkqHMbhUFdBT8k4T2B5YQwjpcbLOyJ4IMX9/tD
ApVmqc1dIU0Uc8sAmDLMZF/Nq+yxMFhVSCUC8N9u/QEEr1rrxV7GnhmJ9Yyg
188K5KkF0H2pjnWT8DxWicxcOyohX3l47p0Grb9w2pr0v5gVNrm+jjFh55gn
cCAXWtgeAq3ym4uy8YvlrXcfnsGT/66P/4bnzLYr0sqbWce1ni3j7fygYG/O
GJRRnMc5CBfkAODXSc43Uc8Qi+3+dqmTP/q1pJ1soFc9g5vzPIDS2DFrEJVS
BV+JSV+Wv0YRahKMK+h4xC2XYIlqKcvzHWj7lBIYYLhRMfgbtE6Ui7YydeLl
U21z4+kfFGvf3dU4slW5A0daMjWof36ytPl8F+CaOzzj4CbcoxImY85Cnrba
25tSGmuR47B4zb/a44ko4a+LBeNYve3lksz/xKULgKbi6F6/KR9aaCpHvsJq
xAZuDfC3H8GVEJ//K/ktjamGZa/mAgkS5H2KF2mY4909BGCfFesttZFNdfyK
LPlep/wP+VZ0f1cA8eoZYGPyTwLfoh52NiElOoKUdJKBP9O1puFcYcKNte1f
Xe+hUmP3RmDoJm73LiCp0KlcY2WcbATBf23BstgLoq9pywhBxrG4+6rlesXi
CPh0UuOrC/DDdryq0B1YZlaa3WSzVm2AiNdkUbfB2AnnBuBgR4bsK/8Hit21
oxVdqJFLUcoco5YfJdT4piXqixmC16Yh6BetkBPHMDTOc63/rosFbCZJWonv
xWT++Vdpm7NmIMSn+RTydzkgEB+94ECZ9hfYiO1lwgrYXqR3H4NDMYd3ZqXq
PH01YIxBVwa14QBPxPzXZGp9ruS3+nYKdaOXJ/1EdoBfAddP1xUA+I9GEnqI
M17/fghLSQ3FKXGXNKPx7imcxRS7LVMJNOa+eoorwCLde6CDRgJ3z0rDzk95
SopPh0/YALDc4ZyxA/HXWj5hX1U9SnhN2jV8kghCkLVhYEA24jpKE0SM/Y5X
XDNChTg26nGOME6r0svLQ++bTGPhSpirTF9G6SjEH82fTOpDkPnxqZCw6MGG
AarRFF7NEkptiYTyjS8mVNlkBW+GHOO03cbZ+GdyqWjHpAMi+lUv9DKc+Aeb
0+yfAiH9kRoAATBTpl1tueciz9X9hxAtrbfNTNeeku08KZz7wOTeI2rfx0wj
NDFksa0VUecmmuSs5cjbMFltdlhI+d9Zb6XK2lj/gC2D/Uy+8Q6aUb4qXOfU
5pVbv4p2dQCC+w9vf/ymePGsS7ssQ4VI4xQ4S6jLVW2Wzv8N/ke14AotzvgN
870UcrxKseu6oExTTsulCaL2FwTCg+SMZDLgT06rZBrX0T5y04ZBVNi/xaTG
Uy1/XYbThsGz26IaXyStarBn2onRp8UcDpl+oj8toyA9nJJLbEX2o9ByTyf+
+64uoR1CMVHLsw2o/YrT9b6MYD7GxXWzAKLcJiK5/yRVoqa/8GlNcdwktbMr
W29CQ8HFdD71ZFn42YY8Xx8YKoMfIxq1nqWVMArGTpT7MlpdiOITUTkqGU3C
aE8IJkFY/I9557ITaaVFTQkB6idRDfzEuZQMmvXH5vL62KDEL0MDJn+XcOz0
beaVIaW1cmJrzGDAHJbgQgEZNHrlRzxycjxOwwLBzAIJDF0eWeEny7o2w5ji
AmbK1+OA++tqME/l5RxlkyC9R/KZ9UCiImG2Xk0t7qmClJLAHAM3j/0etY74
hxwg2BEcrRe7CctzWPRz5AJ2AiCNbHJI/DaE/YC+PTS3l2GBS82YDdXOI2xa
w4pSTULr481Dd2uBtkVe3O3YW0q7VUY42LozHWg34FCZuY2EejInI3Sy0HdA
hD6ruOLg2i3n8vcQzDB8rsiAnYfi2uUI4l53S6ekgBPUCP1S1IXOisI8fGQo
tkfvyPsJCsq0B6K/smXuyXGenDRFs5Lu0nN0aC/b3dqDaODNdfG7k8BoLVXG
e67EzTR5AWBV7l6OMOMap36dEfZ9EwGu5W8IkJar5IzbJMZSCeJuWnujc+Kd
+WmkUOcvJx2YuHCDZo1QdzEuv0fsbqh89XuvpzCfTwpFJkwfA6Xo4hCV1tWx
zkiMo8rRudNSjsbvla6UZ3MwByZsnWTmsOjYJhGKyymOQbk2STKfT/glsy+D
z6rQ9ChWJGJDmcgmxOs5x2B2YW2TBA7CE3UshCp7FtYvYOo9n8NStVGtQY+m
Uxrqz5k4bGT8XPwdLZszPbka9xdlJD48XxIS2t+cmpH17DLRZQVA5B+LdXdq
o9rmZjC5xKWhhbW8BdxJr4z3I8yiQWiMPC/5u7Sx5k0sA105ogifCW8uP+BR
WhhCklmRX5W3c7troDoi9CotVCQYIFTCdpbULEkYx9bqJEmSYcRrnW/sNlA9
/6Q9oadQ//Q3KDXjDyxCdu+YeEvuzaxFuiP4TbyZ1r9W1m9o80soC2IG5qY0
elJS6An/DkEyeTHUOzyQNxQcJEoi6OoLfdRcJOmkS3SNEFBNbHxYh/eRNVJV
0bTtqLt8MLNSBGSLiZz6JArSulKSBsRoNRNkdOoqPiij4Xwse4VCIgWhdv7Y
sg8ex2v6Ni76bgVpPgzbDW6rcTFbk0huJ9/hWrzQTpPTdc9z+eG+jm7E2hH9
bghAyocwLqYSYRxmXkZHH8UqAwd3hLRpKiyE28x+FgFYjT+h5MfT7KP+xFen
7PIgnxpFgdo7UiC7Ik/AWMAWSwuyvBiBzyAAatNa5SOIz2YdHqXX3SNbFBpo
jPt4N7csJ6CF9qjDWvQjNEk7u0hUAjfGXOXZfE+r1leHteNHNRmCxV8Ohq5y
VPPED6jQpVTCHun+6JK+PSL0wd4Uf4h8UiOoHEqa7TmLfjEcfh9bgG8GdRDZ
/6pu1HiVDQFCvMHtpmv5Ai4o3l65ScShr198Q0M7mf/t2tODyQE1yjXkpF1W
n1Rsq+JR0hewx93puXF4zMN6LOKpyYYlhJsgipDNugbg9qCTupFfY+KEMy5c
S242ZAXbxTybcpI9LrbTq+BBslVcXDKXAVDqgB7xLMIdadEzY2QEUr5EFdy2
T6WKHvMTgi+NWK1Elfj6L+M5B/mkJhMmzOO8N7sHHFKdrgO4qd1XIN251bjJ
KQw/JR9gf/PPJrd0xMoVBwvAkkqwswbKXq8kEsLxYY6tCmDf4TyMosyGVKFv
uP6nQTMFJC/Qlnz03RK1SnR+X1m/AcwNSsnvrlYOVguy0BpDq8lQkwApg3gH
7emtf4ZSoy7rQ7pohzqikgaNUJWVsPuc3tZT8HoRjh9Tn+vs7VZEBTszCHJB
QO9V8TdhJK6iR6GmOq/totTPA0omkdPyHmeeq5bQXjFb03jiXEMDJg/2zcvZ
uHNjztSx1sq1+uTMcKoGa9n1n4fpCWTVLilr+QCrhIkDmffGVK4ZBbIdYxCe
5cm7RYKSgNtrzbaTZFUwgnJQsZzIZVhWFimkFcQuUpSWNRZcqF0jETcYF8Ba
LublEKvPAwtR98UV5Nso+rxti8vj1J7FtfUQsbDQSHTrtRjWV6d9LDeKzyc/
gFThOk4cCBRuxkPC/IaCcZLW28diX5MeGUJ5soCG4buU2pOP0Y333WELakpp
tescxM/GfeC95YmxmG4c+J1uYaPPsBqHSuzIVBKau5a2iKHmfaooVZaKU5+F
V/XsbhoUZAjfxaQ+6+Zig3aDv4xptX2z2CdQN273DGNlD1xoQ1WwOk+JfBOz
y1ovbeepWvC5kKC/xx552XrPbdYd1Ckc+gKmslGP4gdCkSFJ6tiDmcVv5lE0
MaHQr3aZUdz521tisr4Nc1algEu7fYpb3q4SeeZwkm+IR6dGiIVTP0hw6Qsk
7ALQnEXP063gkjZ2ylk1qLuykgIad3agQhHnRwK1XZfXVXFOEidWcLQaW0uW
HDQSnqj9zBN0NhxLJk8Pu0UHhIWWyqnO8adwqNaHaAqsA7XajroYs+PcNgPV
nbXn5ynKgRlmc9uKz3bshh2PcIZkrLTgp9No74K+p4qemYVGHxjBQALXMKPC
YuYzSdzl2tw+0hcKC5XFZLrmTthJpLkCL1RLDoAiqL7x+W8wuFmlZ5Kt7Xp7
xAbuPPQ+xLuGanYws/qjbVQvDHNC6+OUmAtPEH4YYbWTDoJ1WmFPJrAz7ky9
5FaY7gLTmNDrt/USZPG66v5Jw/0uLs1oDH432hpWt8dATE2tl/CZ1EHRl0vO
NjEvWGKV0UFrHxP0cgtBPmY72qE6yFXh+3bDWXUGI6aDxOjb9T6jBtWs/N6I
yfFJQIEK/3xMQujtcRX2vq30edcYCaltyYEkzOewwvaS3289WwXc6NsW4lFr
LykjzqrhgVcpbkcWtPsQDRxgpCY0ruULycfgLylBfALpBdQTCWaPhid1C8Oh
SsE1jFXf2HVRkmB4QNHKf+7wYhLneV6DfQ8kCI0tzXa3mXV37ZeGlFAofewP
xfx9k02Pp+nx3GfRe7Up/gGvcZf3nGxOMedLqDO8hGiHMktZ03Zr93BVU9Cc
cGZ64u1+sraWa8G5Q66xeOSgvVrV3zfE347LXJK09PRIfBKFON5XhFLrRvto
9A912M47xzXlmMsGs5e5bF5UQ4Z1cOix2/gj4R4FdwWW0dwQ4GuimrdYM9wN
QFaRVsY7zXh0p9SeYafoesxAQRDeEu1M69TbsPxbqbjXrLXXOapWDdxEWOsV
I0t13GcLelI21ChienTLCVV97NfjYnuZfIho3rgDCvH2eW2pfLYC0Lio5EzI
08Rcdzn3l3/cvA1KcqkYtq1SXiSl8wdtiNDK7rpdcDYxAzwC85IJEtWr5sDO
Zr0Ml4r5DgqF9SSGQa1LbyXw+2hQjcWtM4Ctz3YRE4L4K01pr0p7ZcfFmfFn
fmG1kyqa6ICpILqNTk3frNtRmp7MkjLvIkxWCQ/H+PglR8LxjkWMbBb4CmS3
aPzOlFM5YPKkFxMjJYJX6Eg++8ZSu4hfkcKaAntTfQqLZjoEpXt+xUsm0VDi
vdXV+1opki0/2rVkq9FYgeKQS3JhOB4Qz9HXfQLYDd4bomuoq/tur4dqmqmz
y8veMQKibSu51EyPt/U/k5vvAAtByEaylURbQjdB90STDQBsNilsUImHU9MY
DzhMrey2+7oK4CGN8zAE7SKW8QY7rNis4p1kFO29KaOAtniYVrfd81+Cz94P
0SVzxqDqELodKnPHUrQUJ/lTPsRxkt9h5NTRxMUdR6Yd4CMqEyKWV3n6flQx
S+CB3puEDy/DirYbDivAz6/2zpCl0L2MOkvHFQavjddQ34woq6ozteD1Q4nf
S9uAnQeifs1pmgf4DTt5A5ARZM9y5CCkAYxfqhMhCczwp9Zd+Bce1nkU1Mi0
+vKW4l6xGfse9eUJXueb/ORr0CUH8OIzfsH32TZYJtbJUCrG/Rgg3ELBQC4B
X7uFaWpXYbisOzl9ArfoLsYOJV+qWiPU1vFrttiMg5Oyunpta51/zMX6DfW5
q/C4dv+QNtIuVjtXWkFl/NnMo8/C7IPVy60XypvdzejkNAg6XUP7T/npPVOT
8gAYS88EtO4Hc1Y+tCJ64vR6nNtv0CUdRKzpo4c6wJ2hZzvEdigc22WjZwl/
/pEC06RiYYGmzawsm512m91lDlIQfPigklE3w9ST6HalkzJ02XFuk5TRjer9
F3/c1QMCY0eM0b4RJB4K6FiUXZJzi4dYTxYiuZClASQUCPyVvR+IFb/a5Spc
OVYydt3i5G8kCIaaTRICkWomLK8r2oiDMNUa3DR0QaLS52N6ms/MsUjmOLLn
uNzYXjad5EQWkJGu+20XyxHQEqWiQjpr+h54PBuD0R41VdeGtMCniYEVujF2
3wsCbSFUKwcCX9v/hLWVOtPq04aCPPQJ/uj9Z2ORaS1imzUnbD2PHGwRUTE9
oxDH5rEKBgXV/x1HVsiaVmDvVtQ1sXrKlGqLP/ftCP/YaaO4fjBQ+NWRB/1B
av4x8jJwve4SlgSA76XpW3pf2gqw4Yp3pqM3Rdt1vOoHKUkOxc8NetWwCng1
uwMes1gx/s8Ah010uvGlE7EYl5lIf04aq3BKe5UHZiuXNLaCp5eag4d3thQP
3dGv2dtBbsZe1jhOgdnwVq2bI9wcatqJTfcjvYDdsLrRonsvrE9sdre04lx0
l2UQLcB03X3+w6igmlEDnYDAHCozpMTYdwe0K0I7FDYxxR4JPwaNfdHcBEAE
crSlA1mhoizSI01xZA3ihgxgSD2Sm5QoyOBHc9YGvefPtadKAE1AOVF9eTZJ
ItUSohqSkADDQOks/nLgdAZwXCGmJ2yReFHvD1DKyZmvxlrepECki+yH2FO9
XI4pEa10pWiq8Nhrk6zosV6IRYn0gb8EdEWBmSVmxrOvHPhquVVz/xlCOn9h
nCqTU6ezPeB3cAPZb0A+MXXUiMLlLOWyIIjAniBNqq5Zl3ddjCyegug/8x6+
0A/s5uJdK5fSXZOvGsGbvzIzhj2O5MvVsdtV57cM0LIQNVv3nZmK2ZELO+d+
pDbvW2sA/V9qiOzhUUCuRXLreUnG76QnZkFxWerZFX8OEXSBQCnoqPdxqwQq
WFLPp564vW4jkkguqK474p6BA9wRmnzwTBk41D+DXXSE3Btz998PZk5rWH45
l+XdO0QeBSTfVF+dTzoxHLBb7RBEM8EOzE2Ml0WIZkAhwKt6Ws/SbCCbcAk+
TYW20VqlnK3IYj/meWezsZNaB69PxFJwFVSxMpXmzv6Mj79JNUcYxfhJJT00
H1VQBt6/k1Azg6ullwykmI4kTXXA9onHOjy7WPxdhcGq7ozakDfio1GzU0in
0ya1vcDfb/qGBqAWw/V2utfhhqWC0si6PQo1dN0GXpjqjPMcVuXlmYEVdm9Z
R65mVddqFtQv0K7myRN22lfScl4GVWYo7YM+xuAQUGMG0ykAzzuD04/P/CrE
N437a/IZk+9rVQ3na+ntEz9BqodXdBuqwmhB+JlQTuItliDA9N6+9dlQ7R/Z
2gDu19l2bnKsfe2fRUxTpjnx1zcKwnBmeEDEPVa1IDKhkMirs+MIwiXWqX8u
9CVmzvwuG+k+v7qHRvdKVHLi0M1HrGqXdL4b2upQvtvwaCCIOrExQmhrLG7k
OuukPM6nlkW+yeKLymXWDb/dqJZ80+au5l6M/OZOQZVNH90CPym5oh3lJlBJ
A4fvC/gtAHeuQj984/5/eLaS+9CYYls2eLAovlOB6rrVom/6Vh1my6/B8B+R
NrrGnvjAvoGzT9nzT6tyQtcaCnL3WByLnOu6I4GLK8C8puCAxYRbHQDJGw6e
1xRAbEkp3JCuNtY0WQL1D911TlZ8aWilDe8cOoTuf5LA8vf95ESYguzDf6JJ
9Ls9m/GFdlcRO4dGG3gR55hAjXmErTwsdjVx1K9Fxe9sACq69EzzO2K2jvmo
/Ql/MXvVsewrnE9oJpmZCdkFTe1kP7aD4dS33w/j6QiEZRf+ECaJ2vsodJy2
7E7i8C2MGVpAx0Nb84BbInqZVqKPDZSQNSOwOgT9cNcHECBXn/oDhGUdXAnG
ONs0fBfzKf0SuVYbNMquRATycqEhMxY8efSvBokDJKPVgM41ggbkAa3ke/nc
xyKcIGeFDGKGyLzyaKAZWZtai/wO2ybBA4WRRodwHs0etCN3L6mRTN8Txs5n
5zbmcRbev4sA+OH4H4kzZH1QOF7RpL+gVpJHT7rbNfJFZkrSvHpzLA0+1SJE
i5YodcTWJPMMJybYOhTXRwb6qpUVsRR7aaDj5pmGM1QilCQHLefNWpgv1Hwk
b9UBrMpO/GDtBl5+lRz0dHDZ4gtELNaBnwdbkjGBd6vhKMIcCpLi6W7Hpe7Y
tZt0WDb/+GbcULlvsflG0p/H+BQSyBeRvxBkHqXMnxmQEk6yBdt0yps1ZCOy
pJe0ggS3Rlhxh0uJ53LFkNEpSPpLEKh6t2eWRVAscdXtWzuZDBULN/+txhEv
/J9ZA7BTlDl9HWMCXQuGmnyozj6uN7zfJx2I58JU1bCTnpQHbkjhoLFXZnAy
2C5tjdAqNkf9KsB1PQ7ZvDZcHBprJjAyzXkxT6zrpRPAlk4s6PzQ4WoksUDE
1GQzhGbsq7j7IrfEXsrGCMCZRfEmjX/5Xoee+rfIbfCLo6/vc1+A/N8KkhHb
OpFXBPeyMJuymO96HcwavlJpcdLXS8wtknAITGO/Gtc3csumKB63SDOgIo2U
bOmxqa4z6xvBZ5/5WzYrYYJXD2OR3bKeBKAh7wBP1zPbJ41vCjSWiBP0ArAj
tLz5RURK8GQwMgqmkljeDjWhnEnLZj6Zgdgiz2/H2azkqPku6f8mLBHSUiTZ
Ps5dEBypUP/58EBlAWALYIrn+c/TQDKUV09WtF2397MNG6WGbxNIvzFZ6hND
Kq7p8wXe6F9TOzDcB5Mlr7kndZbm4by02/w/wX8SbviHkGDbN7OgszQdR+w3
u7NUDsS2a2lrPd6GjkXASwkrMq16KSThdHCvnqf9pjIzQQvjmup6xeFNBuDK
ZNCupoxI0W/+UaUNuT9EcDbhE/D7qTe7KbQgrN3UpLFlEPm0hbIOCoPtVJmj
O2vORqhFcnvsiIiamCLvadmC4Bvz0boIcKWCm8AZwS9r2oMtV4HfbZWvENM9
aNKeM4obb8XcXIPXWpBqN6lbm1JqOYvpwlJ9xmo5KynIKaa9KPyNUkYYuMKG
j+K+d2OWobAqbneX1LCtQXZv2jZFsjJicCseH0srLxgnfNpCukmasMnLNwDA
vQcZxqqf9lg+Fw6qgeNLUKB6LT+oiTUJJey+dgLImirlO0xuDxqiuPVgo3Ub
F8AJb/hugccuKhRazV3PXOUDekhc4b3YCAFPNg0NzEk6XhZIM3MY3yku72H1
L+rkg62Msm7KrWDA0IfmueMpgdp1wbPqeNorBbKqVFpDxLI81N+CiOyoTK3E
lGVB88lY//bulhDCCt1ZwjNkoH0x+rbSWI9lkgdy6BF7Gdv9eewPnkEpbZRW
FgkPosofOWDPX9zUiUzy8ddEQkq8ObpY+x2XW8nYrzhsgaFZmlea2Rg+/fwz
0pPaRDNqw+gUCjYq5ZT8om9x/C89/geXyG8ovWwVmg1JrqWsJAqN6a/E0IFq
mBl86jcMCxbWWkb8+kXr3mhSsbw8jQ9nCOJ+/qMbP+VikyCxuC8VShVtu8x2
Tr+73OV4T8tL5b6whTpL6rINw9gmA1fAcqdgPkUFN+BhdEnscS/5M0Gki2vt
0eirjUoQ90+01IuhFQ1eTmocDJgYV4jBFmyQ67h39QakJ6W5oV2vAm9KAkgw
fTi8Xru/sE4OLqvXwWk/+hc0O9OxiAQneiQkbxLKxQiwU40TO6zcn5pxofmO
Z6N95O1IXJbbJS6/Hf5hdKNJ1MXu2tYXmAFpLFXWtgH25pDqI9LkaZue9vnS
cPoZCQh7VqssYj7d3DGwUsJ7q/GSVySgKIGKaiu8IYW2LKdoghF7C4T3OXlP
/5gc7Zlfkj/Bcj8qbqf+5YEE5O4RBYHdCOV5Lgdt199yAZ/KS5G9cwCi4wVX
fGX90y/2Y+GZFbxIAzKubM64mYU2ifOWanPenTt6b33obdaC9/PyxcXUDRpJ
sI8PMltYyELjwoRikEg6fEVB2PB8h1qp9R1Zd0Owdi7XIP2nogataw4yEox4
7wISbFw4EMY8JTEtJ+0mMz4Mi8sTOIv70f1io2HMRiAnq2ncvicXOUB48Ao5
LHNObq/Oj7kkNNnOH8VXmh8+MJhwnGXSbcsLA/okxoZL+cTAITVJbtKNenpI
mfPKeJp2PU1uPM0cxV5eSO/En3x1cyVUobz1AU1zZQTIviuMFjeR+1vZnlk0
uU8A0sfNc3YwcGezyDIHKav8JGHtmrKT9QwTtgK1FOPKZMYJtzepQAZfUk9I
U/KKIJL6xMbqKqSRXHmKVCVXm8SkS1KQn8ro0IfxmuEMz4ujpe7Og36b4OCU
zuswmc63ablfeJ/ucjCJljbDDsMazQ9UxlaY1eyukRe42XOUtCkO8v9s5aXK
5VfgRJfLq9sRieOh4Kvrt/nVyih+XZmXSeJV/MoxWnKcsZr1bskwWnY80gMv
BZRQwz9TgIMMVBVc9BJrgEzSYKgM/LIJ7bOlnHgPQnb86navZhGYRpwRAwpq
pDeLq+cMgSjShNWLIQIivhs03wk9aZoRkPywUuMwSiVjhA6haLAaekBBrE7X
zT2ofYj0ajTDhnHyMCEzRlDtHQRoPIJlsOTFZxbBBtfQVQY3BjGwVD9ndgUX
j3WBZt3J3W9L3Qfp6+4SUsLky+p3tlYQPHv2UjoZGnG2VzKY/xapdXRIu2Lr
omJ0z2XyeoDr27ngJnR6WzIf10Coz6X1XcYuG8EI/WCkKhjmLgZZ9st23/CO
U6QEcr+izzSPzQDWsc1Q4yKZqkjSih0NZTPr5ZtkAER3OYnv7T5sWE573EBn
9140ciEZpYGLbIKPd5A1O6N1rTFct90Ph6VbRx1s3B2Q3DbqBJxo8Z9BztVd
7qQK3rhfdoy0I9bAEIdDyAy62oM4P9b+Cy3eHutzR45D2m5Lgmheq6lPshOA
RMp3ezAL5qjpWPAsZX3dkFXorP/np1OUERKLJjjcbEAwq3tJ4Xb4ClKSW/rk
I4Zukku4ecBrEOiY/AxaqXnUpEGIX6w8Yh/7JNsCPMggSRIhwqOSbUw9c3EV
cmfQD3A3GZZRwtYOwKSejdj0XaOTSEg3EGlri7Q+nOZVZlzM5GTvAuLb4OEk
4zrMflzTtX5knz3MSOnsfKiNSAJvcgAgWwDhdYOdCovUuIi8rEy+/pbSy6aB
Enkx0HhQ877qqHEJpsJxDghBcYfiY03DhsTtB+d0VrPmrdMQvcpzoQhMVjtl
8EDDrdFnMB+WFQPDwSefFkEzjItFWKeHEGZemAFRQro5252cglz+vDBoOuU0
jcTfKBRUxigq7mlNadOH+eW1YnftLcA0cPJ7MrAe3ZCYSzAOstIma6wyEWlN
fvk12yT5h/wtegZdUptraKhHaw+DCQjBlWTj25LMh52paDKSN5rWJ7VjKlD4
Z5BESVEAE3QmRmbebwnpMEk5u0vTDVNGsP9EpXmxtA1T66eXn99zn1NxeL1A
6pUyI9LDEB7risOHF4y5hcFiRVxhsfE+QbUmgfDopeBneDpDjo25ZCzxw79O
TajUtxiU8vO4Y8/7oKtmMwKvunoO8QXjRhKSRAv+1hNlGweVIHfU1IZsGpZ1
SIclCFksnYwgE+BuKGHktPNCnVxteFGPEpXwRAq6MnV8avH5ZK6G2ZoP2Pxs
xIWyvu4lA5pMtXwiH2afcERNfXFC/saTlOgPU6k4+9OIjB08e5CTn+t7Tonx
DScgxet5oHCLhEh/o7XmrzLnzqaxqT5vxdN97s0PkLl7HILynoVge4dqB/L2
Bh3csfcWyqvaSZw7oOC3yMl2YhJLLSQsibVA0ux/1bm4YNHgDybr4wdHJ2e7
j/7895EW/lZXnjNkkBjswv8gbvKIdun5czKTpVnr7i+cVayGd+FR89mNol+3
ZpthA9TqcqTWyAb0OIIRDWYldBj6pEKkeGxjMZBAmAZUJb+nEOG172vTzkXB
ZKELOuwsOrcmPPAM+wPJx2EBUrm4yt8LjtM5j//T9+DDeir3BY1Z9jHLJmxV
ILYKrxFsEvgEx5r7+baRbD1fMk/kKdTZiNV9H+H9Zy8WMf1SQd48BEoo1MHP
YIDQZhZLdXuPHU645zCD2MpuW5tC55vtwGj8SSKnNPgij5AYN+/dP4SXXYp3
yF3/Np2g2RNGtthRbn3JSdOhX4erXiWdvq5MK/h026ZvCf+4r7N0mLwO7nSJ
RAmk7YflgtVv7GBnz1BOjsY/nvGRmSs0YbJsgOgNVjw1yxpjPUCsokbg/sEc
AT9nEv3d/xeWRPasJkUxQJn2CV2Z0qZcdnzeeRh/AUBa66bC8BQCSOiy2sOR
jou3FcAbAo//RIIBwk+ncHCN7SYW5MbDWk8WfLU7VJylrs4cM6AyZ+F+nwNI
Yb4LibhAWjFLI2P/Lcj0ZYoztlBlELj4QWORcIdGRH+isaTBjKk6rYAemK9y
t0mxzBSPQ16dtnJ4h3Q3J+3/7a+eAcncDdwqz20axPy7d+egtFX/Bz2abSsw
DVdXTAp4Gd+L9S2e6WJcRq9LWt56J0+qhT3YfK8NF2cyoUj2rPX2Fpm68VYJ
pKRzOvxeT0iM40nxYl3sghW8rTK4JMa4kzlzad5Pqz1WKe6D5PHloXiTUb9S
M7KzFtwEp7Pqe9jxMUysnrMoIEC57WJlDGQS2vENiz1zyXgkguxhkIMsGNdh
tn9D5AKBHUvltGOH/Ifm8df7qGjmoNWyAvPdtp07j8pDrOh4SWQyUwnFdp68
iXy15OYZkd7HY2G8CyxL3uNXmoGzUzH5BD1+CWtiNPMnaerk0TtID1aN/6xd
mhjEcbcTI2Dt4Nu8Pt/nlxvvdSLSa3WCPCvZieUzagzt1Q6L3ZOKzY+vCsYF
nJXgev2R57g8DlSm48AC2eJpZ9uIYIj8BKzds3SpDxT9pnd7jZtlFs/jds8B
u9ZxMAFkY5A/CR2yS2IO+XL89RqUr3720Q/wYDnpWnHoXQYKtQKHDgXqdAtS
C/oefFXz60N9T0fsTNUts68Zf1Q0r7gv+wbMKDFxVMuaIVuUrhGC7Nmchj7b
L8UCpWRzVRtLGfFaHfNREmftlnUV2qB/M39uum9t6tO1j+lL7Q0o5JBC2ir+
4cHtUNjDlt+m2Dm0sceX5xO9wTiwOCFIo1cOuAtA/iGSh2ry333jVxbj5pYb
UlQhSOy+t3NGA0TTHJ70dF35q9dEE0ewHxG4ELCbD33vBkqL7QN/7CUNBn2s
UNPQB51TL65sU3MJdb7qk15mXVDepvAWHnMpHzJS6+QuQ9UvoUrDLPuI7BHH
XO8OoZRSSOJOVZdhIBbyCtqUvIeABvW+wbo00Afiz1/mFejSKcJAQw1N78I5
8O6JYGeqS6NHc1xadQMNHVE+L0iIFtbOvhSbPgh3S0S9P5Vr8YkCAGW+14+S
mleMUplyHxDkZ+0FH+Aimu/rT+wvweDOXc2loXEaEetis2F0U6JeUtZk2c1u
KyVuctpk7wBrhFbTMHPskWFAmm4kUrCqPAhb96xHnfcjEprKTa45HuJ8TJ97
RBUstXz+IIDtNM0sjTAAUEfdqysqHwQdTWFyRlMwP5jucg9VgJAuXDolslVF
vgYseqHC0l1ZqiMNx4dwrLIIjPUm9Zy/tbdEOGvmFDqHt0qG+tAG5RkK1Mpn
cezFLG6LIk4w72XhBIF8W1jf8s2X0DSBVohygmQHnZgcOA/ZfPxqGTCiqCnr
m/thjP1fTO71LDn+T5ic6Vqj9z6MarJcNFIgWYqneHlOQwDayzLZ7WWDSQ8K
ZIljLsyUVk3Dsk0UVffe+Dq0ZoU=

`pragma protect end_protected
