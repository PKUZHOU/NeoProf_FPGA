`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
LO117rqEmbDpUJbbyJT3FjSg5P3pUM1PLS0ZCMcR2BacXV5LllbAivSKMGVN0kt+
V6fFGpr3BwYNraa+QTfvIGTwohpxKQ2aHKLM96VC0NJglrgZD11ZzZO7wAL0mW7m
KIOKOCJTfgP7LCd6lbrpKfbaGwuiKn3PF1a6c5JwL24=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 9696), data_block
e9T4pcPJFKBI639N/SPuJHyliZ/ACWV1d1qtjxSqBw/C3Ug+v5Cmzmj1227VS5tN
QNlO7d0nB4RkwpG8GRrz95IhuU+11D4YCwrvwBptbdY872qkz07ZcSpPTi3EVRCM
2B4lNCl9S8Vwr1Vh9yeehtziniwLPyVeFEBxaC9CHpPUz1trbjkCbJDZ8PAsWsgh
DZt/LDZxjuh1EcFvUu4lis1wDgBOaCntCjT2YEYs8w1oPKkht0Kn190LPBOk9zNs
tCHEfsPwQ2rfrn9ndirGUAquwDv02E6kP4/qqdQJ063knlrUSZIiwBQvWcEIm6D1
/MxjVSpz0/9W1KtotmOQ6+7yPUXDmLDCbzxFx4oJokDTVVBc7xMcTi8Qm4LLe2S+
a4CMv3HTtxKhrDTL1DytQAS+czhiSpCyvKyzqmE5PbmCLBPmROsODcP9CM69jYAX
cqAhf7XHo8jhgafVeKE/uBS/4pM3VD448b4wqUGOj2iZAkjcI4lORqoyXHmWS4DG
XAH0n2whiOUtbvU/G1dtvsKHZqSEucgL8pktVgrUxt4YVCPvE0DMmLSkvgFQWC/U
D85qZldSGaeO12a2jGoeG0at9M1cFvVcASiPoCMwjztVFT0cXEUIaVNjIiEYZ8fb
aiawS+X3UB1Iqdd47F9/RmLzuglzoceLLwbrfr9b9Ih+EImcE9TIXc4ywUety0XN
xi0wrS1dTNdpUDXm6baoUf1GSe1aed7h1JSH3BepCJQ7lfS4nXc3BnADhZ9ytYM8
FV3HnG+QlCj6HwUchCBAoRXUWo3kwoV82nzVzgXD+A7QkDBpiwswhfZo0Pmm3gjL
nBgvQTcDfsBmyPxn8z8WKbToVWMoHmv6cms5AmBF5C4XWdXgWvHiXz+/8eb5KzwM
RDFFFS+oCUtupJNo5+QgzqovKW59C295SDKLax0qPCcucgTx0xyr0I8W9ak+U7BX
RQ2qDsLL33fDL2zOGzPhDt9GXoxhZQiI8NvxnaACfvLXHoRWUSxnhIduZx9TeHmH
6SaU3zkTc02+E6MPSMViKqZOGqm0ucnjjJH9oinuDPr/lffN2o1ThvU8QmB3RMnX
DDXwkO8cr0p9jHUFQ2l9RknQdyl6/dbVEqcqgqgZ670anCAPwUz9aHlYfj+p9qua
1ubFaD92Q2V03nlbIr+2FqoS02mPMJ/1uf9g0bauy2tN+aWuF9awNC0Cy0KkJIl6
jozeGUFAkp3mARj+l/6ymDKeiLLWF0hI9MUly9V/EKfVvMG1bWD0x8BqxQnmX1Dp
nTCAdNAcUceLVDO9Vtxy98n08kdBOLXFMtrC6hqfsSGIgtR4yhoNjYNXkgCkkAIE
DUn1RgMgnel53eIx5JZT5R62QvAbjtqu8S/luSuiB1aIpma9kLS8jrMekpfALc98
juNN/7lc+r8/2l9XL6TWfQCATegXD/cNg9oEBBZE/yVAViQMVrJTyKmdStyv64pO
MlrJjb2p/WD2zePXaInUCW+CwXIPw4HVXMBwFuiIcU9osQmHTB9EDfnWzbiNMcbP
yd4FXIfX2GOcW07/9JQOFjpCgmlFaTUeClKIV/LIofVCb3WrffB7YFdF46kWD1La
r29iDZh7TLSWMQ0quWMY9qravx5aziuiAbVbQAUpN0kdO6gTks73FNB5BffOpZvs
ztvIZrW52HPPtQmeUX5ypbn6oJo/DS8clowagS3vuL+jT1QnS+IWwwodz93exmAE
Vkm2LRPQTDIP58t6gT5JheP6M/scoMtQ+O/6EAF6LRAqv7re1srvzZgSSmDfULVN
c6Irn2kNpQC8LWvxiIkIEuTPSy0S7W1LREgvkCRij/467j8GkJCl0RSyERCNsobx
QY8oNXCyT3d8NIZO1qkn0ZUeV8ilO5EPP4lY0E0n1wh+SlwDCN/poxBMgPN6EUKx
edtzyxBXLYai3ncYi5QOOpJ4Z2MeTz55bF/oXy06EOrRUgl2F/tRYCGNhd+mtiD3
zCpCRsZYVj5la7NB6A28LsNg/0Kh8E7MvqvfALfIkhuu4jWZbSdX2sIeW8UQFg19
mrRhKnZdYV4crco88b1dh6WLkIF0Tb+gZV1HJyFszRSR4n95i9LQ3Lec7XhV1q7Q
8qcXiAD3rjF87Xmppotlgz8ucg943Qv5hidjaRnnbJmEnWXbBkBRISLuFI+Lyb+j
N/m3BAiB04puSFcle7Mvv+tOvM3OpT9jsbm01k7eZbtrtoD0AYLwnQ8HhteQY99/
sf3x0Pv2oCUIQpvrQxPuH+MgDM0/rVTplMLzAPTXbg1FqYLLTKQQhPJNX5eqCYce
Tz/OZjqU2cLApCIUe4omWCXduYc+W4lanQUGM7ZyFUqQ/gzM+52BI3etPQHsearS
lVR2FVagpW7zFv929zdVC/+DDXOq4pzGPOXNZJOtEkzo9LnKynPiT1ETksXAUDvg
RsThm8o+ybXxpSZL9q+JYvHLq5Jv3a/ZA/0E3wh586WuLfO+rfYbj4rr8ZCqnaFE
cgUMU29PNQfP0XcE7HWnATQ/7xGJXq0V5p1eQYf2axfSubSYzLOqDMVKP1eOvTI8
i5ziSvMhOgyrwV2R4WcGIFQweJT0PWMOwNnOGzA5nSaY0NnFlhmHMENkUQI6YS/p
wJbHKeYy8sdXF19WnwkCfpyR8VLLDoUI65qIJcTYF6HOi4chAR+H58RdIF0ykLo3
LkUmVI6gHfkAlOfSLBSDwtk3sCJAQK+GZUgkzk07UZ5XL8wPe68MXeujRzYQ1OXx
GrF2mMl+7gNYQZuNeNMi9zYiX2M4Siq5neg20kBA1n7BqhpSv2KoL4wiNsBX3pJi
WlzhYj5ICmEu1RxtGi5KYJ9HVCL7rpSzINdS4RZkTrn8NWqu9XEOgRo0cWaSVBrQ
Rw3uQ9TF7Y/riB791pEpSYoMwgIrRda7xiwCwn8WG6/Q9mMkX6UZOF7FWITxW3Vv
+8kwLo6TdK4zPK333o/icAmzYbzwLQyUpwLSBGNqzFbtuv8fzyL+/feb0QeqcdXq
nDoFMMJJvG5f0CVLs828QX6pUKcH2xfhf4Y5/kxbEcpejA/W6aZr5o35ZKqK4Nwf
xsaOQPTNZiujAjIyB9oZgf38acOj4xWdjKM0Xh9dSMweJOf9sK/L+1VeJSBZfYIL
wRG5MWGT243frxIdmWk5bhQ9shzRloP7j1xeHhceGd2lGky2sSQv1SKV2icER34L
WzOvi13nyPx53Wt5yrdfqRfA6nkRH5AcolF/P2kw1y7hAf+0ZrHnojHfFl3h1Elb
jrpzVMJ48GwcGtJxC3oxiolD0Vzz6JE8BduNML0+asgkaUIXEpjFKGjNb+43Nbcp
v2eV1433LcC2LRCx3ZniZm1p86HIUbkh5m3FmlzZtaVGxnlKyaC+IUx5/kRG/JIi
X/qyRMQLT6725fw6Wx4aECfNM4sihUx4U66ReNI929+OIDnQFzA3+FYx05h1TwAo
HuEIgqm/T4WHF+fRZH/usUs7cuSA4oceamwMJO1uzXGJHwLQ2np01ndkcKFQVXg+
reV0gkFbvSbcWXx3qnp9u/Cnx6cEOCdEBqWNf2kPuCB9AxelpUTu3KmHXE2Znwss
C6hlsvrk+ubuXwykvv+R+IHOUG5d7rP7g/vfJSTv+gTYXFX7th0lz+w7tbZQD3bC
LxusI40mqyCZWRd4fCFxTkEm4VEYE9amA5QB70BpBJdFPV7VBqjeLU6N1o3e+ccY
vlo9zXV5r3UjYVthcv3R1Yway0Frt156rjo6S03agvn1qswu1oz1da1JKO71SpdU
QEx2Cs2ZbXprK6jor4+qutbXHF/z6W+onqvFG35nO7TVchr1Ptxn9zuYIXCGXo1m
Bz8MoEVc73xxz+Li6u0vj5CcSaQ2nTeOWntbxzB1GJy1e8d2PN3V3cpHLgVNdeO6
JjQ5XPf+w1h1DpDK8RmuOegwtUy48yVMsQwG7zp73KxLp/fGoAAKkFCdIP1wHw19
bqvdkGfXVvdAr9UKuOVRj7tDex5imRVxyRFCby2iHh+VIardwW05OI2+uz1qZ69x
3gSWNTTe8uvQHWMZG2eqWxsoflpn9Pn6v0zwIuPWNJYxR64hTJmr7QJNdmMz0bDn
5VeWgByYaKbBUXbo8dYurczb/pwmLPFOs0GVkGrfJhaK15uJtasuGqz9TLQv2Svh
rH3NU3yM+Runig9NDsHHf/0+vEiRTQa/bh/8EmYruZiHSLmC6fVsiKvhUtWFFm//
EugUiWpcO3aNdorakrE7w4g9ITztpn7rrYQreQ8C5SzoEN39yrDzskTwIEwDDOAI
fgtL2WO6UrePxUWIoJOCEHXC5SfKgmVdcT8piRBua/ArRn/ejgTlGXTANcUlHyhZ
uGWZxU2aOT90+svTSUilgDWe2wZw5aWvKwnJqdqT1ik3s+OoxEuUa7YFPNHjzGLw
misLF3w2qY3m1HwUxrdOnZlo6DEF/GL75zGpUL+sq93sWKXgPF8c4HEr+uBJTWnt
ox6WIUueP1pT1cqjjGODEjyJTFHOt+Ev/MZo7QVBCaK0JQADReUsMUcAHVFIUpw6
JHaSHkJz/7CmJpZNYCo6QdKmqJberyFnDSasBxMH91EDj6M/rRxeqxiMt9i8oKrr
k5JdPNR/YOkLUvfiXG/oKtSejG/wF1KsMRswXbo7s22jH0whwxS3Wn2cjELG/5I/
m8eUO7xEipCE1pkATqbg3nZSgkMJyAKXdipZLnTR16FKQ9hgDAWHBUYgONSzrrNI
G/eRyHBaQNUhYceqiCVIwtrEJxxfj0wH38fzXxyXJwdBUlk0ZxmMbN9vLvTv1nxm
poqxflZ5ij3n9mBLVEaE0gTjb89wNzGgHzTCtzBm7W4G1ent5uLAtIFVCKe+UMPI
R9Mz2lJaL33/nuD0OgRSfE5psvYZ7h/CFrDQTt3QeVY56NemJCzrquG0MJbf2INY
WxTC1oSR489Cw1N+NyELZ+AfO3wVQJhQlCQ+3ihNFIFDvUWeeZ+F0bMGmtPRM4n2
mCnBSQb6PJHWRZCt3O6WJWaMBA17Mo1uXCBQgg70OnOAFs5dxCDD7NbjjgkVQQ7V
t9n1E2wJu9exxuvhj3+l2IyBWBcnkP+rrR1UIxQdQcJjA4gnnJYS51mutoFtyA24
K+OSvL+tW4U+pTFzMC+iBy0MVtg5wlT1DiNgQ/uz2FHDY/dG1I3fsRVhPfMLd32O
mCEOoWbYM1AP27OCBRCkUud9LSMcKnQG4LoFkkojcYBWuiRzjuGj0oI/J58jZn+A
UO1ApC+BkM3k31unaTZgb7FglVdvcb2lpLNZ57trwXeKSnkGGHeOh2XaJg5g96Sd
/e1bU8psL0Fxas3wQtMbanM/exm3rB77OCItDZ0m6CMazJpjBHDoXB3+FwXP169Y
A8yiOsuDEG62HZ0kjNiiL5NI2JwuKAR/2MizE+Qao3j5oYXzOQ01Kgh+F+Ivt2or
CZIzFI54nfdDP3fJJdfWm/wrko3TMynQ9FTA9GQpoGb6gUYTcV3yCSd8zDU00sHi
bQ9yKTlzhu/HKoK+zGnQs2Cv6jmZvoxigcPOPcE9fvfwva6b46XNMP17CBbY/zo+
WGWzLVdzj9Zn9V0eQUXCeZ9sClTz6++JJV52Ybus2Uzgx6lxszVJsRfFJIzj/d1g
MOtdSGSfqSEPDvAmYHp37rfjBz6IdiG0od0iORnywSMPSE7NcE/nKq73mHjOCfWR
8Kz+TnTVPnSeIHUY8stydsQ/t285wrErPqXiwO3cHupNcU4/QgtGgEzRLXU8vh7e
Q7fHMSmLhfdG6GQQ7iRIrOtVs/9jzf/TuUKVGDOGtj64K9N1kBluj63xV7Mb8qC5
BLlxOpZ0sO+efFfeeeMPQd7a3cp7PceIO56JkKyCtADeVTsTi0ZTogwoW4BE+qCc
UVlZ470IR8QZxP+YzEnAcPBeXzAwrhjG1E88xDWUAIFGNG21fGdisX8i7lkuqCRD
+idfqaWMgA3rd3ZmgZdpJ02jYnjwDHQQm+G+koxJ7eUGXXfAWFW263AGJ/rWgE4U
wUgbuOlyZVpmZACakONk83j3+s94Yj08ruMary6x9+pTu909xW1AW3M0jII6jn+6
OBkSK5MSNWMtKnfMf8r/+UVW64coPNjdRTTDNZ3KJIvFtXt373oUw66bRx5Fu9yp
uaS7eylzqqWi2tFjf357f58+jPZZgW/oNEBPk0tLYgOdE13vUVLLH/ifkyR/d7oH
ZmIo/w3rPiD2bhBatgMqGK03bK1VoYsZCWfg1fro4uA8D/ZkB8PmHyIRL5sJH89c
e4ztrtStXq87pjaoc6r08deVjuQyqZa9k9lRBGjxP4j/T5xVuk014K5BjeuKa8S9
7bDQfRDphklR7saUSsz9YnUtnksuMCDAcZMXlEdc/xdu5ToLImkI0BltILVyPSRA
vd/0iNnxV28TPNgvdf8hAxE7DZmz10ZZGnKnRPO970Me4w9PpfhxVrpOFa3xqw2R
D53bj6YNFcd5jwXFG4vorWww4FTiYzUisxDRqELsAm8fm7gXAPbSRgZQBXDwyuTS
r/zzgmqYtHlEblkHGJt3zVXUCFRyB+MnwR8xN1LxbwmSL/6rNcBpvQcs5Il+OpW5
FntZsXORkYnScRymrOMLZHajidxTpXueCyeGwL1NPnWtlgRYVzdM+21gRZonIksR
lnvfwPb4TCOB+Kv2v/TjoH16JIC5D0OepI7mM3pLwTpSgDhzaRG/pbtbU/1bKVw2
rj2VRpYJwt7C1Vly8YtxXVDZOZPTmKd/Ca8yMvEl7pMQd1Bfrl8Q6NR63Flwwb0E
CjKG5ejD/XEYsBxUvCtinUgEHXFRVodwghRNrU7uy7StY/Xs5sublLnntHJA8Ina
S17yzRTKIeh5nSZHCiv6Ahgyn3ke09Qi6ELkX9jKTOFKJ3nKCM3Ws9Lmzas9OGD/
osaoSr0rTONPdsiXMtCcf0Qx57YFwMsJFE16SkIwJPF11wdqoP1T/h0yoKAHTB0N
t0xgNJe8rKQC3TJB9JbB4cAMcc5aAvmPE5tOHMLv5YVn+PKYKn7F5Sz8VxxXoptQ
R+l2lB5cAY3+nPWEmyM3/3iXHLKwNIYPR3wZOMGkWZwjOmpNk/DHfCXVpxBOLMHw
o+TFMXBfLWuhBxJg6NwIX83fPfElnyt+BPRYo4wYQ5jHNdHgdf42TcpZEew7lchx
qyxdcGEE1w7Q4dxXp7ArNxRqSma5x6cJHvz1lQRD1Jd20KfyHw5ZN+RdDHQOcip+
X4DVx65mb15iW9sj5vNKrfAhiTlUf3I1mSLJ83WULsUTRN5C5/UF9LTfzcC7jbXi
Nfl8vxdsF1uN+wYdT91TzQiPOq2fyHUdelEySwtvJmSPjf2Iej5G2Tqhk8boRw6L
YUKRmVUAgoVh6AT7OxoIh+zhQnv1/lLknpgN2h1JZCQrYjNuSVsLDSpO5ghzkfWA
4w/lHu0f4VXXQ5hcrthlkPlW4S8bE83UpFGAS3+ozEZRsU3e6pBahSXGRlQ586Mn
D73C+zubAE0vjDIBrLbdEysNnKJYzyRvdK38CSCOR9G0BmMdZaoqG8uBrfS9N0f/
184gj1kVzWpugLt93XYwcPm41WdwM05fwfvisyxfGaL+LsedCCc3meo0sXWbew2P
Xe1TYFN63edK9TOAXtM3AfiBc/t+oejLfAtJbnlkH5YPqRp8DBd6HBtq11Rs8Dmx
G89bydhRwL8NnQEquD5lwah+df8B5vchLxH38bOJYHCVPB53aBRMBiqkz9KQPv3I
Z6wMMnnryeVAeGyKSz70j+K8oHKrJ5zIM48atJnte415avCJ8HyPjPJTJpbkbzJv
YZ9uXVbVVNNlSGcXSt4FCgf80K9a4UBp7QMyuulQAueRytoGbonutt1BUxrbO5iH
W6/njPRMXnKuTgvqmrt1TEZ6KEefv2VZkZX6jj2YQx42HpfJAnNsdU0EvyywoT/J
/86jpJxnHf044HNdrBoi8zyPiyjDWZVAcTf3owsAqSXzrql12cruUaq3xlsAFUX7
c8XYHHyWMx+QqXN1LqqNjk8WAPyk1esh4mm8HBInxaaZepvikfKGcO6nRLdiU81n
k5KZiv7WhwlxZKpEvv7SW3P8NpUpBzKeZ6YEVMZ9HNpNUpjceNCHRBDJvsTvhC6p
Ltob+z0pV0tqB6ICLmGSc6Mxs3NWO6+njseby0DndBIetZ0PyBkDaAXNCXaYAuCK
c1G1lJDKeG4ihSCtbhwb375A/JjH/8A/7giUHoytd/GAz3aLhTGs31b8a2hbLmXe
DzKu9xdnVOu9ouIK19YJ80C187a+TN+wZOi/+xGZlxwseiWsoE+yVPJ73fRXUbFe
vgR3oyMCxiqtuv3KMcZpTE6bqeUQGhEdDtZqw507D/NcAf3bBOP9OZBWdGuMFlBA
6PdzSKl4ujxJZ6BMa8OZLMca3Rc3ymTUQKFXTs1ZNvqTSNH0O7wONBNCq0WjRYeb
77MTmPVPJ3pY5e0sN+gff1RIHwiEepBeJcpslR2ztM/ovH6HLXrQ9NFAewoLGhB/
TvgioOATCg9L5d8HV//mFUJu1TMie12bKDmFJmPWktdC6HwNZYgw3mx54Z4Bsg9U
oP+wFY69yOPHgRt/wR8A63+g/7iJuWkBKRBA/2e5CamWMtAYHumUqY9J+2VMLQWk
ik6t9PnIO7h5VtlYf6txNk2MmGncxZU4Ez3HuLjihPgALjZ1OtpSyx06/rVYWUlI
NiorXL6zYXybHrMbxx/00/B7TuST2h5dEN6GdFaR9r5aNkYwopE737yX18LtDmVp
P64o+jKyN56j9vfzy9qtrf7rWwnrY0cKo+oPFIBZlJt+zQ8I2gg3WvUIk/Wvwbur
JEb1lLjmjgbUcwAXrxD/gHNzqZNjLVCIT/J2VN2l0RyIlE9MC5O3l9C5wRGv8ebE
h7zGhjwRbWqfr8Ol0TzBL0qHUUOu6OVmHrc14LdUroGVkfkz5MPlLFhXzaSmIDHx
hyYxhtv4o5BoXcwi9+8SMJdg4Hl2VQJCOddGtKbNukR8dsEqX+VvILHRzeqWwwSZ
8GN9s6rhePwk/hne8ERFiv2MXdk/uoadxWNQ5nncPIMpIpXC6yeokixXHT3S8nZC
sluAFXRD5mUVM+QqQJvoG4QrXlW/Z6CKzbr0KCCbP9/LbHKgJ1pzMnrQAA9T7PFo
muUmNEJc+PZNMc+N+IH+C+EvGDJQns4AgpbqhYimRt30CVjTbFwVW0PhZVbgY2Fs
ARDSBZWZ5j2VCnguPEPnVPntZwsaGoj1C8SuTfW/7b8cRr48ndHRnUdsOLhGLejU
y0NcbgDD0X26QrK9rlS6fInqbcJ2Bx5E4mN2C+fye7VJ2apJAtdxSjPJa+9DYW6C
pMBQje5GiZX/7QmUrrx9rnS3CcJ5n7oF+t5IjcMrH+9zq/EcpIcT93t+I/8WhFrb
h44dXKMHCb3rAMPXShrxo538KDjcO7MhS4ELsbEkdlu5rkBSJ2th2OLBa0xbxNZz
vFtCPcFCkxLTqbEEYollcwvWEis3xnTRSClpFn8fiX2Snz0nEphI5wSWfY8ld5FE
fQplWB5Zc9YG9V+BkXNjrIB7kQjTIM3WfxJpEAwalq4MkzrT0uq4gQ2c9l5zqO4Y
jybEUHXDyhvutaWYocaL063wXu3LaP1FwhdnLat17ezcg3pK2qd51FRhxXPiNpQu
SzXVnhpMHLidG5zDQM+8+5EoB1fdHnBogLh3nUwu2XhRvHWxaNM8wuSKLMiUQB97
fwL2HyrVk274FbLs6bxiGqhaGgTYt9ilVMl3ATW0FExFhzEZSBN85CqQLP94eqTG
rPP2JSr3n4Mdoe2LgtRxzf4fqsKCyHg2+XLlMKtqDuMijMLPDO14QNKerUQ7yaOH
9i/HjPzji7FPC3blZ7KOQDfH8bK+BVB5RjjkV+sjhmL72fx8bVTfHMdlujxMlalE
pfKTuwDBA4nc3aP1IAhwwjCoiUf9LwfM7l3Rw2uNLC4Y9UDPuZJhLmhzHoWEVFX6
G4EWrSHfqPwvy7hPArs4ikF4ngG4FZ8ywmfdOwnS7jNxGAYM7HepUiYQ9XIS6zVa
2/cHVHiGg9RvnVMHZKJ8rh++ID0U3yb4DgJ7LStYqxSFAs+67ml2I/ieCZ99jRZK
aOSIqH1NidoBHpNiCcg9Ao6i3v/AXkBpOTsG4BJY/W4Hr9c80eUmtR+c+p4uPFry
8UOxWdkZouPjPe4ngaLtrUPlJWhllvldMne/+S3Ptt+ZYXGd79js2X2jejxKqKFd
6rE1BsGO1DYdLUAWqAg5/fdZ/V6OY6aP7OJy38WuHNJBkftC21mYrDOUBZMB2qAm
CoTInvYfdK+O9WdowMmkbkpWvCh8B18L5QQqItKaqk5lpQoOcrlhVx0Srmq4RWCz
LtwTcE2hpZQTdCXM8oHGqcYbVfHFvjOJ5TbuL227YB2e9iqjdNlv7coN96bGVOJq
5ySUe+0P+zEOi2V3sWBy4gV1aJHlzBIP05bh0Teondy3c4adTUlD9QLo99GTGiGI
KVSszxdbAnWbIRdjk5sEJWjm/aRghS2gYSguiiF3WZdsSqJrVl0itgmuqdG0NWyl
k0YAMV1qz6KD2UNq0Ws9frkAaBkRsKHrrioPLd8NIN98AsL5fx+kGZ2a0SLrfiO5
G94q6A2SCuNg26q+M6CFUcr5DQl3xrNFsHHJ68oymtXobEB5xhMQFAK4BQJFgSg/
XPtrUteZZDgT5N1XYdNgSmtDeX525AIStJDRDQy6EDFgac+V6twFrz5xc9toPs1d
2ZmCZzY0nNH1eGiqYUqYZKcNjWIQR9ckkd+XvWg3GFnP+YULy2/zkdB6oFHFrKof
xecbTLLN59aBDJEUw3Ui3cGcJV0B9NbRpTqkmdPoVRNeP/pQZnNIAWVCXoZXygzL
NCEbg6UuJKeLlrFWVgVM6TajaSGRU7SxseTJxCLpHGrAJs4JLmRtfcP5RbplGNil
EjayFhSIwkDmBg89s2dhcHU3eXE8oFbB6m57h6YF9q9g3Vf2G+YTyeuNKJHP+3j7
7bne8OdhqmThACaLh6gxpdTu6LJgU+GiuqerrhbF/S6QFz112aGQ5D0tpdvxd/XX
orBfjhaP/KZr3EJmrrI+VuEylYoXXai4+MYXMyMBXFAlEyzW7MCFqY7cAhSCB6Xm
w7Sw01RScvqP+WiBe9jqSzWF+EfYX+UqDYNksTIFDqgZs4apkNCppWDr1fH/dj/4
dbaGYa0MmVzJmIOOXfUiBGSXhjC+cLNuhAS0ncnyCF8OAcCnwhWu9I9HCdG8+/Nv
8XjF3YnfMSOFoDHxYY6c3YdmbBfUXwd9EZwbgGZ6rjSRPPS7M3Ov1Fn67vKV6SnJ
J4d62SyxpzJy/tk1c4L59Lnu9IOIVdEOZ2lfvHiTKWf40GZQcXaatyHoB0VIU6r4
IAuEsxRJcznEeJDTZ8SvBrcGGmlanVkhCZxGyJQ8XxzIe8G19DUn83fcjNrfBaxX
kiuS+icwRxp/txyVAtv9TtySAR+sdFvlDCx7OBxao547mFq103EsAryNg88QizUf
fKZ9TCdzxS7Z3eFBZR5FEmYTGsxew++fHQ53PX7BeEwlfBDN3bRoVWZ7stEZfdpV
wfGNWToQs+jfksxah0QVDhkzvh+tU2AB+ShD6iNan/mKwjmZnQDYAgAkEJdc33v1
25FkjgT940v5LdSkaYikvSO40Z2cZHQCJFph0UolJPWcNJlFfZXzwXDvllYyBNXY
5q9UthwMWC9x9LP2VB5O5tvhxYKy9oH4Jz5Qx/PaXZ31vsnpF7xD6wcEoN5Z4+Ab
0ymIYgh7OvtfRV5D95tFVqa5wLfQbXac2bN9no/5njxy6UlaeHEV2qkXcdlusyFC
DtZNU5YlIEvqZT6EMGmnPVAp2/lyMezo3QdWwz1EPeW+dHnzFBmYk/aIk4dT26TO
bfUV6cFSvfkOSMrQ5ZFi0inSedRD1Dz+OZV1CdSxwRo2ibCJ25bwJOkjpCcBWKJ5
i8pwY/cNeXOk4NiWNvQKRaESrdanQqB9CORWfZUMdoDuy5RzxfBqd5QtxDL0hzhc
dU0e7Zdnamdu5HUcwJjaF3qSRARoSL09DGsy+ScNki59jsbvAIUB/MOyJlzRH18m
FhpzmzptqXJ7eP0ux7U7gXLAGFbkmDlwfMNxKcthYnIP4jqX+S7qTZDARpaYJfyn
+q2w6ySXMfWKTnJhSG8D7MOiR613VF3uQKv0sUZFk9alZyy/54UlnVIzlVk8wr19
2c4z1UE0nhTIG6OVyBKoGBpw3HZST87b/8TNOCjpYN1S+34LxOWmZr+jBUvCPqNX
QlWgnDhVQOB6biFaIHpVhtBRqx8RjvuWWdbkk1kvV/AT6haq8+E18LY0dzksEZKL
/I2WNrZX/pDjlloHvGa4uHEuM3eAUwJj5TFLhHBDIEHRKqnIRRmbAeNmvEqcqnBk
rpULQX8J7q40fxQsRIkQIL01oCnlo8+Wq1Lkn9XYoY6FHxnkmjKi2bCVaQKO2NzM
FQuN6XHxc9zTpyQo/S9NX32uSkSA/Hl4fpP98Iejqtuxpa6iCvEIGndBaiQtcWje
4cjIlqBW1+Ujr8S/aJD7glHgaFat8Geu/f9u4sMTZPuB6BAxEgqLqQQPHX0try8U
MGMLzodyf3Ll6RKSzDj9M6R6HFxoTo9AYbYt9XWWiWv3Eil/PjezgUmULoMsiwWv
FvWm53b86/mzc8qFzyKQxc9y5A2H5S8CQ5ctACehR0tgVBV5TDSS320tTn0RY9zC
Z4zf7pIa1O/rCy4mofPHu2qMcr/JKhuqA46VJmP+1onTK5w2dVs8UNEnfOAZso5r
trtKl40hyWOHENr6JLmqHo76awsDgEAoMRutdLPi9+4abzj+/UBI+pSaSGMvaJ10
jekJjrNShjHLuNrtXaoNhiklSvdvIXT1GYTrMlNS/YyBSQSGCTdhrYO8Ci5Yq1u1
`pragma protect end_protected
