// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
BVYH2cnv5AktE5Vli0q6tR0r6CMAnKn4GDOS5bmfxwaG64ggsJL6snWBEcyx
xcX5gyd8IUOCxzv4AqhsRF/NkHVn3WY/Xhj+z8USiLZS04i7z2ni8bKT5Tl/
G0ojmGqcB97weZMG6z3HOZNgZFT6pcAwJeUbLt9scER7H04o/kbnWcGhNqmi
EHM8XJftRcEIAl+McJUhclTiF8Xf+VBjEt6h5kJkXoVRJsduCd1Pxet0tMw1
bcQxdedfgA+E6sVpc1gAtlZNNfo1P8lxk0eaam1ZOL6x1MNqatQQMxzF1+qb
UUMd//m8Cg/06lnSHso1VwhG+nfR6D9rYZEtj9sLQQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mgYTA3ozwozptD+SijimzRk3EKEGrTrq29+ICzkEtvXSrYfWesMjybiUbv/J
nqRAkNxLvk7HO8Hbt2XtycSHpvLCUIqDDQ25dHkwXBVHSxmlFL83kfXUmuHe
V+Y6GuIDAX6lYpXhMHp1NIa4A+2BJ2P/DDPdpx2RhzvkHLpulaBz57GVuuHn
9OUf42uEr2L2Yl9+6bW4JQABkb7tZpLQgp8cef6/Cp1Bln4nc4XMv5yKOjVB
gLm6C5XKwSK8B77pQPtp8u2ah4hABduKMQRsPtF/ygmxfJaBzRyGEV//5bq1
P9Npisl/5l1djoehe4d72xbJ9LW2Bzc9iIgsIHTPJA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
aBlz9OqWphHG1yCOq3aOKjoUPpidq4SzJBINFoyn6NzWzFIVbjYFHbYYOleL
HXCrfu9MyiNVXQbEXr09CsE7EKZof0JUT0GUG4TMp2Y12dGZ9coCpBZ8HaxE
bE69rhW5hrcz0dvqpQRzZa88UyFPt+n58lWBkXT9KJDo9Pb+jeZiQkiU8+/2
dxiYLrGit4GYy2xtr/9nyoaJXTgQeAhed5TcFeeK8nOIsG+L8CMfhj64x0Rg
iZfp0t9qMCD2qNqKu0MZiG56Ay2Ztgrrxc55IDZx//yq12HKTAi8HLyLsx2K
/RIZ/5ophubETb7QIK8lF9lJp+59GAsnBspxnDZ4qA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
NPNiJUaGOa0AGOjsrSJnVnPSvySkUtONXGzpHY4kJ7hrNwARt1Cq3D8B2X8H
Q028yNRH3hY+zKFgD6ubgDICzXwl2Adg6LtwbipHrLEgwTz6n1HxiUVtZf12
Vou/Jtgi4pRtevyCrsy7mngBvlxvD+SQGmYia/XwmSpOczpiy0E=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Etg2wmFvGouhBWM6oNfjPUz0Z1OIsO5VvvGKPi/fTUvXgulkvQHy6cOHw6u2
9tD70LgqCzVE8PAr+TsOHsvqeJtcdkh2pVQGLIu6+Ziqh8gathwQVnkOih+6
kSC+27kDLqMW1Rb5uldubV/HCMayTiVcbaxPxXbqM3YfJjKCC4SDRscMcaOt
zpQt7Hfea2hm0FpAEKOzuSAFkE4y5lrhMnEWJWRBBVlNOc4tasZlD8jqMG9p
Eiw5UYH+nvyRzflDfnYJBloLxoheTWW5EiSTOiFrvjPxlPqfP2+HSOqLsbFw
ozTiiESjX/xiCIv0TnIWOYASbAhI4Blr5uNtvzOyvD6NwGHBI8mEms0G6VnO
Zq7ApIvTfek0GrgWEczBByS7RIAxPHDC+KGcPY3bexN1W8aprqX760wWbkKc
hZTTeVl8VBG5gfHdVpZjWyrkL+ft69Nm+5Or09K6vC4pYw+xARpFA46ZPAIN
Ux6DdE9z1oDUTiOmKT26x+SponQ5eO+F


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
GEi1VrQaQH5d3dKYtXtXoIg1bvdT3i3p8AsXLC041MEIiNcfdTqm9d5bg1ms
fBr0LJ6iWOB3lA5who5ZNNHv050Ygx1Q9GKLTSc32fV6bLP8cJIP8lgzja21
PsMbh6oJ9+xhRAzeRdbwlrXl52CRcM6YYi6E2RX6dUYW9LAo9lo=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
iM7FtpXFJDaK1lONrsvGFWO+P5nQgmNE1G7QUYvGh/EnynQo1JPjgeILi4v4
Y+TsmkFDQyloP9FbDu/W2iuH5du9STAEYuqgpZ/s19JuAAbgZDWJ1LUrdLYI
ooTccwLFjEoIL8u5xjHNwcXHfDaq6pkY4t6UD4dzdsJ8BFuOJdU=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 30032)
`pragma protect data_block
qnfa9EDjEMsMG+4rbY/PFmKD37j/WGY6sUydsM6L+OL5Z55CnEi9+qSo9BpX
MPPsR3hzT6l2HfZYoMQ8gnklFYyXcP2VbWcBRmdEHK9BFn16hy+ulxExUQ6M
EjSSnwvyOOZLvl4/5uF4zvSTVO82fa4r5l1YwpcSbi3FxkYzdTjNHBjaBSdU
+TtMbBLr4It2BnFJqoQEcw5pvbi24gWL+SI4x59WWgt3qX+u3mcux+GtFX08
h2T8UuaeVvcbVip5AYkc8t2jsLVoHYy+Gy/zNlD4ZSfWlO/Jj8CLp4r2Q+5x
1XL6zrJq2gEP7KF+gXbroRngmy0M6ryq3iB9PZV1oK9zg6llRMty8nuJeUWV
c8ZZkjY9Pk60f8u+9NtGrxWWxcTXTCsJLyWEqmMpQB+CHztP1NovbCEaGp0S
H0it9vcuHC437C3MIZ5GlUMqttjtDN2QALSoahaCbEVrZn2lZxqsXdyWMY5V
ktHpW349UQU2DpMsaamcMZ+mMdYJxUNm9t0ZEKcB8Gyp8t1qrq/YYHPN9FSr
mnWQzEqYXoWut90FwqmRhN4tCXm6ssP97EJ1f3WcFg28qJyDJRWxtt3rSNnN
f+QrqwIn16W124LFH1WArrgUvaJafRDNz6gw/d+CIVWtEdyO2VVrcdDpzCGD
CpiCHDfpXQp8RNhqbn7ECwGRmtUMrVKhRuhre8qWknsS7mkkiW0WesyXomWn
dFOMQffF5OQjpUrI+B8T42r2ynR9+3otfZaFUWEdf1KqG6CGkjx+dFx0SABL
kCEvzBYn1GcR+ZtZKY25PJ1dOEph2vnMFUxvAxEwtltn9mupq2yWYsScv33j
7Fj4MF6X8UDLapiLFYa9ruAHZAJ/obNfu/nSa4OeWBcdL3l0xhmgg2ajxc1s
6fipy+a7Kr37ivhKoToMA97h1llzybit/G5GouMIBvIcLxWcrtktPcD9qjq1
DfdObPc6pGHo1Mr9oO+B/BBdildlx5GEMJu9EbYa0hDsgeAmGv7cu425GdDd
dnNI7Za9Z+kgZ6aEn4KSmhOo4ZZ4MOxsgnitZ5YrxQbeUcKPecb07N9B5UHu
tGGcoWPUdIYg3naLNc2CgYGQA563qmvrLRvIdaFGC6Uqywb7gHiEoLZQTP2i
Aq3ezmH16J2SB3y2WcSRXhpS5q7W97gdsQLS6LVGYpTs4tPMr+C67FAht+6C
SZMwsw71pWMRc0OnLVxQdp8cPQfmykdoCE9aS5FCkhztJ39Y+TNgTUlTyZV2
/FMddkrYFX/opAUcymfDwb86VZKeejj74AMsfIkzUzFDwO0QIG7W/W6ppVml
90+MnDC4aZEj/juZhxa66zV+oaIOMm48npTAu8mikgivviHhyx8lPgLHHYwV
YlgJfsgkkMFQeoHb4eS0lLcWF2JDCx+hjCbjkH8uW/nm7fpTLrdt2lK81EKm
V+CAFE5dKTgnUngr23J7pUqNevfcE+AkXRQJAXIq528owZXi6rhdPwVAjLLS
cy+xDeX69/w7Hf3Oy5CnhgUa3nKGJW1MNIS+63aa1NzDQofh5DAWRzxs0Qom
Rp6hWSO0SSwlfFRXlt14RVw1JEDK0fZ2vusMFZ3LeBkJX8L7rzaZzqP2gNAE
iGXBTnfAZImP6r5RqoiWETaG6C440zgK9i+J1X9ZYNTw3z3EZNomsdk3tqqa
cQJ2PX5QpoEOsyILVExjx03VvCIyx4hKKVTw/HOCpbvqOQD9ygm7Z3dxx5sQ
vIxJY/WSevBx3Vhxt4fXM8dVd8NTdca7zX97aa27mlRn2LGLXkYFWL8Ayn9s
FaQnbjVlvYPvhga+IFSIpEYMsQEsdaWUmwEr5Rzktdj/vT5Zzw1bFT2bjcqA
J9XnF6R+ZvmB7b1cnxB1D3J3X0avJs0x4eZYkjoR1JcIm3iDZ1JbiIgsYf8s
0Mp9fSInJz9xQKA3/u+MNFgYfSftJQ+1vYru07UoVGj2W0ViTIQb+mx5yJrf
cKlM7FRFrBHYAE9YmBtyeuuef9+d7ggzdgYOCGRlGUJ8lwH8rEg4SGNkQ5QZ
tMXYIRZ9k8Ja/VcWhNamEr7ZeJLIGNdYw7guXbJOuY6Di3H4GviSqEpuOuB8
cfpTOc8KAzw4nWrNvKXMs15SHm6+VRz+B6BuIi1IeNPaV0Q+W3I3FrymIChI
v3adGCTwX0uevC02amhhHhYQ/xaTFn2ABQ/Vpp9nPRaLiuIlfbqNQA0f4Bcq
zNropbIDkakLvrHM7O3JRKKi2xJ4UMudFdkLUe+lZbBjsUN5PYQzy8xHwxeA
eRyNEMQD+xZVmoiBIEb1E94UIlZh2q1EE5/DLUHW7DUpHu1elxJL3oJofGbe
xj8DDAB9tjqErj75vBYGnRdAtFfwYmghghEZbiLp3CDRWHbWNkURjxQlRibq
LUqk/0wrPvLb+6ud5b3Vbi5piX5n7REw0gDAUfY+t14bIO2fqQt2SNlqD6Wi
6gcS5Ha4hMEtF0PG34+ma9frXvqgaNCktzooAzvmycXOppMjghh1mq1APT37
l2o8vbPn2liPgVB+vuIUubJ4kuxPu7qIDVmfgOD0+pzUsGJTbyYhzxQaFTrz
W+RppIoVTUt24KW05vcAmOxB08ZslaJvw2XNIrPwqHYBlgE+QiAHEVUVa2h4
Ctbz1heBZxihtA1gedVWXIpxZtz3oro31KdvHYL+rSoz4pffAFwDZQ9HIsj4
Vazdk+rasKOzHuqIBOxqrvPKUhwwo4yyeGmJcFZkvF3wI+QWt19/wTmf2C8X
LidUbUnuj7SKuaht0TuKvIpJ/fsleEGF3Hsv9kWvluXf+dQXZ46E6yuiLrZM
ACySUP3sRKZxYVI+fxII5w3lxosj866c+HWJUgZxEntp4JwidNxl951sh21f
mP1l9ZHlsBdZdxhTBa1pxV7PB6q3tng4I3eQzqUpSXvzO87XKXUIjHk1upER
eU61BAAAWf2FOIBEXMR+D+VPDWiPbU9ysQGJL/qNDyRfxTKKetukg/gKxAfo
7aIo535TSFJkA51LJtfNv8eZyDa+M3mZQ7Cystn+jmR6eDSkuh6kmx/+wm+v
jZ8wp7jvyejBbbNbu+inbaH/k0Ee9RkRAbaVipO62f2/+uwEZikaVBVwmwJi
vOygbOkNhIDyU+WNxEucKKZh7h0FSpH/KPrmOLNYEMshlIHjY8Jz1f/1knDj
Sjp7C/kUjiYv5pzh9AjqP1Qp0USMHYMf7ERgGjmOFrqpk4R0Nx0Qo4xXpPee
Rg8hdHva1qgld3ABS4xaW7JzrVZ9SCcuPFGMOBemb8Ht1uo9Ju6KYZtfln8+
2l7u7GDwFCgfQ6T9gkh/HCk1jWfd8ep8xI8tz5ed+2mqYMSbXjYAiNCp4l1w
a11ZF8WRjvmTis2p3fbtRAAT/JxXTVD501s5FrgBoznb8d76vqydMJEvrX8/
4Sh73+47Gcj+bpKTSohoO1yfp0U6FTkOLSC30wYXTQ5TAd2fwBBt+VFSO8B0
hN0l//G3s5KuV6mfYaOB4H0Z/hNWgMapxJk2QXo3klEABwqmE2EAPw8B+rzj
w6JSrpDQRHffa4M2IBMQqMcFx4FDd5YgnonfJra49NQHUrFjqoNN03Sr6tIl
RS5tNOu5t3GQQjvgrhiJlZIX0qCDaL5+UEHxNc8A2chOZ52v2vq/35OGBd9u
9H/Hfxc8iLDhR/m8NcRiV/Yib+725rLCfEP71uUu3892rDzsRkTdrb8//sfQ
VBqXz+QMPKKYvNNjvUGbAD3asajG7O8+KwWqjule1khEMJjgKcpnGpLD9npF
BVVJeDxnM9OjNR/ZG1mjNB7wZc7ae8TSlj6g10KccZQjGRAQoXoJNV3VxjsK
lT44B5YVVRPDRlIaSE+VUt1dqiPzTKgv/IhRk1zwBZOz8oWKUlsI60DfjJhy
JnI5hM+Flb5wcTNUsPmhdzMa1kdRhsPSasWRwA9cj5v6w7tedHWP2F3jKL5o
qglNfZgbz3h+F0dcib+CEMZcrIBFFi31kZI7DH2A/di6+ayryJ5Fke2jNlmm
TYoSrlCEJh6RqTyvbux3KNZzEaVxcUu8ieZGj8MohKmiMP5G+68vJXMqfKfA
jaFV4HteakAtbEspWMhcOUfVS5LtcoDOSa2yqjfPs4FN2zrT+DGiZyQTgdQp
Igxvt5wuwP+KWly2EFKtTH5c4yIIhzhwCZVzEUzMKQjEeiFRe6gHZvJl/JQb
FigAjv4ju0ggV/Dinm+Kv5dXyfxC6Pns4NRoR45Gp0qOewia/GId2C8tFuxL
51gBQ+KN9hW+dySyUtPIsMwzXmPRW0k+UVe2ZYFinjsRbXCxxgQcC3ZS38Ui
4TAcJZjcJvfh5XmOHODCTOBukp061QHhDPuY23LCvIVj7Ioxe2/9wtPg/den
fg8ssVZ4nXpR8KCGvkNfcD80teWdisF97+VhJhBvmSFvUFavlQ/iXZcG1sH5
DNfjngpB7K8mjk9xtOlnENUMWN2/qsEHEDCDlNRqEmkgYTV0QGpQE9g7nLVg
jXxDkK+yazeQru9rbywfVykhC8lW7/DHlePEXp7BKZ/HfB9246Vq81514Su6
sOHvv2XPQOKPDqEJlu7hiqJ7NMhZfv7ekh/Zeo+UZdj3v8RNCBl4qky9adrx
lGK3ONVzlFfWWIZTi7Onr/8weWHnmpPWLQDB3NLwYCucbn7c1r5QKSqhfdAB
xQBnBwbJr4NEfLvC7kmUpgsIENoY1V9+vYaTy9HywTENBwwjmrwR5S0qQ6cs
PaN+VHfVv4PCmxuyTXu4Ea84n3aYAD5V+qzdNEjRKAsr1Mq+MNqS9Q4mKHTL
gNeOr5u9+qlGmXNfcanzv9a70Qve9gzyo0qCMPXktQ9FgoVvmiHe3CavzDni
nJPYGfbcSeeJvvprwQ25xwBp12mA+ZqHYfdL6g05Wy7keqfR/i7fMhsxnwrS
omDO5TUTaLeS0qihAyknxkItj/z7hYIq++EopB9SQEmO4Ip/QmAfhI5rAb2A
G61Z0gVJs2BlWOgV3WJ5tVkL5eRcMzmqbLoqmj78tfu7RMojAA/taHpu5CXh
+ayvBq05t4CxYbZggbBvGsn03HVhQelemb4pY25QGLcl1mz16tbKYLPPA5BK
+UqtHg7gTUqLQpicvw1DBydhVZKh05WzzSr0Kf6RwBYMJvlfQ99+qq27OwW+
NyMnIlF+IvxtSirsoHxS29OZYbYzX8n8GoaA5+ExpycK3xv4Ypsa1H+mL0Za
Ior0z3zRMPeM3a0D7WeAcOvtWua2uHHQqsGQ/BbHSUm8LCVH6FjS5uUx/1F9
4vDwWO9RrgLTKNw7wvrj2vmcoz2PPnJ1dxODo+bQyyGRH4yggmOB6OPQlmpG
gEwCjFANNZurUFmVJkPNgqFsXbccobP1wHNXjMdMvgCgsfVyhhtuWQUDpdpy
fyumxLDXkf1vvr82assCZFyug0k9mp1bhyr6PhPJmYC8XlN4qyoRKSFRt2kZ
bDBfHPob7Pqlw3l4FBn+UV7GA8JWkvjlFzua31bOxu8EYvoes0HLZi46hWb9
a75tSmH87zbgr7Fm1RuRv9+5G21Pp2CvWbeaKPM4dvD3DkLo4An+9qRChWCS
mVQUbcQU4BgwEqATzyB1ONShmfH1fpLUsNJCVMwfzUV329ah/DdryngDz/o5
LgPA/Ozn89WSJosASZ4DpICHmIFskidvGpMXtKZ2L2JGHGkdZEuRGuQ7Ji8+
fjAX+J2lYhI92hRU6YFug/ubZj6ifDysyQ2gFObem1oaGMNn7ECvx1OBVVwr
+fjgrek6bFd7SWEsaFZ4LfVJZ6sOIh0J87RkJUsFInIPa/Vs+1xOtYUi1k/8
pTtoPCyA9nLBfuwmfu0gp05C6TD/ixe/f3Sux07oGJS6mfSfrPOoHq6ukONX
veZH3wJSBTZ3dUcUppjZo4eVxG3TIfsgilvi1cTw01DAORwqjcm30OMs8l1n
IO5vMkW27Sh1ovi/U2tet/5x/Nm115gkT0QRmD+rbLMPzPFxmxsx8cUCBxAR
TOVRi7CNixr/YaxvqRBOZFJFYOQtDSaDrt19l/ah8oyL57qcrJ65jNbg2sN1
TYd5U3IcH3Kiax2UYHdv8mc1dpqlCATQ/zhvDtBXiFuYvN7maLdoE3b6sUeA
68buoEEOfmCzUc8GWRa3o6gWI1pkmh6cfN6pbeufp1lzrf5wZXhRqzwYU2Io
qUnD3rb52n5Ma9pZ9rUSeiVWfYQR3PFBNs39IKb9Sxeb0rSCVPLWpF8m3kAy
R4cwd1K4Euwo7Iuz6tR6rLRoWNwlCqeq5LHZ2fwPpU4Xl7gsIdhcb0J/RGXZ
VaW+pw8aCtP9ljAZVz4kl//lKIubGiLISAjv9TPqy6zd+8sgmWF6RwmSRvUr
KGSMH9fSUse6f8JpseM2W48vFYIVafD9jUubGORsuy9b77OJ+Dg6SSlP+pJJ
5QRk7KzzZigQ7Ks6iYpoK7jzsdBd4g1QOuq+ooQz1z+E05ftCw5LqQVYjQ18
P40smA1ZP4Tciw39XQ9z1O2gn7hy81gq5U65nr00eE0TqTsDonFuCvu/4oKb
PoR1ut7+Q2rDS2JDtk3XGg9VV74sny9/AY+7derpFvhrQMm6q/f9tiqy1cqH
cuUxfpPE4ZR/QqkQLz8L4A7BxxOt9yzXmLYNe/va4WEzL/bBHE4+fXRQ60DH
XzaAGTFkOv7EtusV94ujNy2S6CHpIBO2UYbvXLDee6h64c9BOHPV4TLiznlR
FbBSPoJP17G9G2+VZ5AIlJDFlQucNfpMob8g17tfnPRRb+qzn6xBHomabjAn
i5aIcksVIM7UQozJRM/osS0zmEjzQ/ghzvB43LDuwJ89Q7pLfDCnUwM7ebpW
8KtDY9+U3vSzLmnoZZ397G0RASJKJOxKjRLJzxSHfkpSDj6A/3M40kAChSHC
t92SEVT+tmhNpaiITqfi7DYotRMofRvjdeGM6uwwuJkQY1rk5nojWwyBdOCp
/uBfbSO7y7bTDLSuJZZBX+OonV2XG3ghWFxHYIs2CVMTAkR3RyWgVZoEJ1kL
iOyXe95Nnrp3+YLAoRWSWQAPyj4/Dshd3WMSyPAC0MZj5aAvo5nnL4KMcwYV
sXW3XXnUlvZponf6GlG0w6RTDElrJ3kNvmx8yZ1AXVpaYnVC69hpZWRQoRTv
Ho/JnYcj3EV36c9HdnAKvV7hXJbQCNJjmUKx8NSp5DyaAyc18IHrVN7dgA0B
vrUzOT1sY5KtG8hyyjy1TCdnu9vfvOOVjs8Bs4aTRSnRKeiHBAHQxFtLkzM/
cKGHR1bD4kPBA2Ddoc2zdH3hJdyuyTBFF9UlJRyGShecscQqmhj8kRdSa2SV
xP2F8qPwc4zfahXKlwfEsRrvYRTSC4yHXlZkZuT6VQxnjGMrUrfMDImkZqCo
WOBv27XIVITHVzSlGN1WmSgv8kkyCGrhOO69jAhKDCccCHpGdjJSqNfbwEIo
gLksbTn8T6DrtIEyg0nkzJswpChbwQrwR/VlWxQ7/5tjr8QYmEPfwpINwu3z
y6BVr/LSU0TmSSLa41x0x9uKNEWSp7cW1ntnjqN7cg996oytNeDoA9+KFsI9
bRVIzvaa3wqKrpnwcw9bl1K4eBlfXv9GKXZVXuHpTNEDNTNKsWm45AKYENzV
RhrKBYD3bXWr+2j8t+k6x09LN+5iyzT2ghh8Zvb78If802eCSUcRuCpQJCfY
Oy+f+EPr3aZ0ojfqIV+QHqUzPmdIX/L8ryg0O0HuF433HuNmfucIHcXLo+MX
+lTJd76/CvQz8ZNOxLRdk2wmM9F3TCnOV0lGWuT1KPoSFRiCuBvYP+ldD6bk
k/zRlDk4doJXDPG8pDfpo0NsvhRiBHSxM8C434yfe0XPWpMAwkn6BqCPOEHM
2EDfDTKTZPB8rE4bcabaxH4ctFnP2BmqdpTd4z1jowneZRmV17261SRVupqk
tcu0O00sxbFOm80vjzamnaSiIlbaI+9+CN34KX8rIjkckB5woKlgvQOynaCK
pJQOUNZ6NS/HO3kz0tGVwnXrD+ygN/s8R84tveaekW/1UfwrlvfisneGznjy
o1NaXDUDgGRpfn7QUMZEs5P0UKw0qejOVN6ktR34bi3ddcUPz4gFDmYDEkOX
MtKCmwfNA98iDtQRT1kO0IZWjtV3BHTG0E+Cwu7C2VmxWG+GaQ4ODMR5Ievo
PUlGhvmi9vpGO8trxuo16lyYRJ2I+Fpmqg+gBmnMtBfjZ6TBodxFnUAo7Z1j
WbJjt/dXI5ncpHvMxTFvfpjCAhTmxSFYuJo65zrAlle3KtCKIXRtVZOaPvcU
yDvGfeBX77iPK4OFon1+IbEsCPcPQvjAlCwgq829Sxu+T4oNrX2q2JrrcjW8
x0XHtEWV32NJKLUo8NmzjkUvPIwMiMCPnZN0l1ANfKEm1SsS5k8wuGnYMArb
Zy2jeXy7x46crTjt/4GKBRuiYA6LEsCSgTFgG/cDCp4kYQt8ZaLaiCCi4Kop
113cGhmuoi9MJrv4/JYsPAmvAPAd8trp9hkj15utcM4dlFNvJHGURJbyWvZl
8yx80Ra0B3cpbU8Rsmgm9WgP0B1kG/cmjOSEDnrtxw8Gon1NyGehGrPAzZ0x
JXy/7SlZ8erOH6nA1EAFORnsgsSD8b3dqkKgfkElQQq7xHbc8E2KgtkQ9W/m
5CzPyhGjVaN8pkqvWxuHiOcu5WEJL7mNCFwtF3MoWqW/7A7OusIqo1zraKl7
BZgz8tBaSLK9z6lWYGJnP7nRtE6wgMClNXxTzlYxSHPeUND300YNAfgo/tGU
Y1y1bo1pCY83R8KujNAfwo8iMCHmSIyOeSw+vJ6F80hWZIPFoUOb33yLwqsB
CT0AdVorIwLICJ7qHGWAr8P80unp0s86vuu1Dfz/empTq9HkrPOB2yv6k4dL
mIH6RV7CJPH0BrrFeB5FD4NHn8l124MQVxy38V6NoHCKz8Qklbd7mTdFrSwy
M8Xz90WsUqUFavbGDimbAn8giV46hBovUWno/iRU6clWG9ULGgeMfRwnIP1k
uC+/YFwJqm4zJMZsbs3dGrO53sIBAkDNsL46WBx6zmsh7nJ0HQz+Uh22OtAI
x2eJQsCaAzriJrAkRz72M3h0LgCzY+vvNEUIN1eroV1UrqbKTrlDbmFY+kvS
Gb436L+qf84NM8B+y+nQcXaDn0CpXJJvtveHxvTD+H69kJVK0UxlbtjVO8X1
+Z7yx3HrSdLevcc5eVbOKYaJJYv7fr3DmVo/6VtKwmfNsGNvE9j0eR8tEOcu
2lp0rjUPGLsEy7P6RXTT7n+lHgbdRBSoir7rNdQkheOirsn1BDPY/l9HMRRf
b99iwy1MuwWjBNJ2twgpH6cjJoxv1PNBxIkNv2rLX5sauEsm3b/b7Xkv9yqE
z/W6cp07SHq+XbtcJTsG2l+Ie6JfRC5/a7Jp/++oIcF2fKNX58qKsN5Nv7D9
6J7WjE88N5l0IHv8cf5mUvICbHDMnZW8zfhsuKT5grVAS+uWf0qVlPHAzYIV
DlrtWMHCTB4ENfiCE2BEM57cyo7dNh6E82B6dTveabF/o1sdsrMRHogNcSju
s7c7skeO2RHXoNQIpa/C2h0eq061jds5l/D8JF6E0duLRGoiZ1Y0w6au8VQ5
U6SJdNA003b17UvHxA/Xgs5w8uBvJvsO1rS8oSC9bx4q70tiN5ZYu48gvUV7
RkouKk8G2PmjY4zltauU46udDNlxrvUn+1sDIKQj4PR7V+0c0I7ZMpD4wAe2
UyUomXd5aCvozczb/JB0iCwrid/YvnOvOCOgoWrH29jHyyLW353lHhjmY8HF
6CImwbiUENRFjDpOxt5kfpMejLQCBo9TSbnaMA0Xo9QVoCtDXXAyBwE3CNYy
nE6rDFs/gC1LmqZwG4UZVYW38PaIJwoLRHnW8gT886smYP/uajOtnQN2egFW
zEYZzgrBfNwXYt3vm62H9CKhC1OqRnbvnzvt3qwn7mnkPYaWXO0t3kqgfwMg
H9C73ZQuRpSdplo7H/JbUl0To4kPjK0o1a7yBdU9RiO9aecXSLbxoEhhOQH7
QcnVniAQVyW+lZiaNRnBndZ0VUmFBFPLgLW7qfgXQv2iWn2JhGs3AYA3g0co
BOllbpzYrTTREKyPF83NkCwGx59LPlW/MlqGsxsmsy7gMMSwKm+gYCwvzRED
jT+HXCsx7GonDk9Y2MV2qwWHQzW0xYEoI9brAZcsIfPepNPeH1LRqVR7dVSJ
gJqpFAiTWkSmwoTgzq8dFJdfvvGqkvWB+3I5wOQs2cXg5d5678P4iQpJgeDX
KzeKS2NY/6XBqD7QiFlbuKh//6SKypKTuZlXOSL1UTFRqr9TvqnttsxI/5Xu
glhljds1MLnpclopkN6FSeryM98ew2Y5M4hiQlyTtm6BxrWLtReNVcI1v6YG
lzvRhMBGlgtXSIHF2Apsq3+b9YYUwYlf/NIMQQ48h/S1UaA4cDWXgGAPtW3e
9OHX/ehE/+5g6f8UJJoTPTG3K5u/QSDrAWh+e/XzwSQ9SOT6vA8K8bTZngxf
fhKig7ySPTwNnVhxygCBUO/WU5YsTUAOAHLSwSqo/xnD5J1lA9MxyxTmv9Fg
/hGra/kYk5UEC1yJ4aPfFNOnGf58PGCC2zQQ4yqym8Vxu8bOYjyQxFrm61xe
CU2zEYFfRnWlskQbqgAsuirtr/wkG7ltwkX9zQHUqxdSuqFnwBJazrjYEtmv
KxrAZGkeYoEKAMu1D+Xq0m5k1j2mPh105uiG79qzBX09eCbwjstMLf6LOhh0
7rwrclyHVWE1sOLXIPkdKuii2MNL6VUh05yB2y15/mQSFVbUoUtHuZxhuCZ0
OPk8mm1akbseWiFL9In5iS0cJLDzzmJkEKwAqYvKqNcVBJi1ysFYuU4lGitY
8RQc6jZxkaYerIItH5bLB4t6wPln5zkMNgu3+vCUt7iu1SKFWDj/mC6vsIHt
jqrqt1lWCQuTLYGA7/8tRWL88VjirGYHpl9XBW7rnU4dOnZnZSd6V3l8DTJl
obam6HR0934rjZ46MoDeqo+rv0qUe1BbRuKYsNfdo5EWoT+SWXQI2K4jSqFh
xwEwvdL2KiuF10fni2bx6zAoZhmCqLHl1o5YVt473clI7p4f8fQAXWa4deSv
Q21/40Gbph2Ur/tqMirYv1a8cVtMoEtpHwloOpTiOTbbJax+G5pv4yRlk7l7
MAdsO2qWBNYjHFAS+EDb9cWkDLSi7D0nq9Co70eZJYqm9VYgWpRoZagR935l
IiZwt+j863IZxTG8Sap7ua+j+kIQhPpMRNxaYa7s7QvtQtqPZBxwFS3FtnDK
0B34lLiWucOiDhHMdy86uJkwChzzqZAsKlDxzx12bONMFzLwwUXqrvlPBWNg
h6qpS6fxxzF5P4LePDY+q6t6C4dSyLXSaN+Y1QUBFJj8Tx2YcajmC6aw17p+
VmtPjCnf1sAu9zb10D6yuKifXLdfk0BlUHLO4M5y4+oPaknawt2Xh+aR0txN
+y3iBFZp/md7c7hJfZMRxDONyFXVAft97RJ3LFvF60drbrY5L1ea8coLLUbJ
kkF9/PRwplnwhUs1XZ/Xo3R2uFaZxNfZttTxBh27EVloorJBQkvHzW4nx/dT
yDgdKVtlY1TsEPlF/FR2/nNqV3JyeZTy4mFyDEaq2K7F4q1aAF51yRunysNW
j9B0vCpBRq225HMSskWMqe8O7U0MzBM/PP+12y9MbLb9iWobN8PZ/jXKtoWb
LWith13kDj9mocjkBcWsvzpqUyYpEKjf9+9h/XDD9OYwHWiT03XyUMEaNinb
zqlA7z+u4Mzfgt9mZzsjeylNJZuWsERcYfXt107wXdvSswc4/cpD9+MzkpUf
yernIv1JOuFN+IqHkTr5c/gstIWhUtgAlK70KwO+18flndRBeo3cNxoeTfXs
CIex0qdWGhZOQBjZMAj5kvgkN5U4aONfnl/pSATK+QUp1RkqhHw9ZIoTFnaJ
FMjpeLYA58Qr/Rv3+W+l7jhqePmEcAY+DDf2OZVrvDYCZP5DHpXFg0BYVHzQ
pg0FEZHb6rJ+sSKi4wx7z7DDU4r4frm3JH2s9Myu6HyO9b2Enq6v3H/cU0f0
WFsn6e7e/lC6haUz0FCmU8Ug4movFq82FQ6hQi9gpU65dlRDmnqm/fYD+bju
Uge7zJ8HA34TYFMjbvg0BMjUWojcqcvbqDpRnb3jzsHJwCKWEm9M0MzTL2eE
PxPLuiUjadhyXOcTlUPxRI3xD4FJNj5wHhTg13mrsvhbRweJ6/blyjcUlSTk
STOrNmkXToyXjF66yJRrnLTocFayNUPhrbKqsZgmX0QLLQASRIZatgSDKmJq
WghnLEQEzadMljV2IO3uUcZ0DhkIapA6BAohr9YYbkim0L5l4x+KQAlEyEO/
8unTy8sYgQZor3/TQbkM1h54ahOuxCDlg2eRr1xCgisNVNwFS8Q82Z9FcxAS
AlKyHeRtIO6hEjH/D3Kk7tsw18zsaASITIq4gjdp4GBHEysWiLd7su8Ek6jy
MrxDpT7MlGyZ2KsibA2A3zSMfzbMsluUEmvWA+ZBP6ZyawwHgHm3ZZQE9uOh
RggMnMhHTeHY2mgwEKFz3OwzuRICb6Ht44dvtryZaePU5gSnBlj57wgqF6ce
Es4ttC6TZ+M1xnCShG0L9aWxXjCjIrzRdbOe5Oo+xf4dXfr+kJprmvPtX/5v
GCFsSn52S+ThVtEyZDEYbgaDcqwPNM0kyVEtUGYuPSxtE+6cBGTatur8f712
nvREOF2UY0Nst3QMf7c8MYvfKOG9O6UtnkR86BHugUy7IYuUZ6CZ6MLy0nAo
DcE/TdUHrTZTxsT8uP8QYy1bsalEe7peehfBuq0Z3EUgfAHYsQvGlfIasWrX
knfts4TwdRGHMMFEMD3cdWP5N337vPxo5Pa9DvcbxsWrM55VHW80Y2D9GuS0
pUqKziu/NHXAnkkMqoycLw5einRYyrLlqiFoq1erXGUZpcU6RO5Cv1Zlyk/9
KlrZsOFrdvBTx9JZhAJ4b/OmGWIJcMhMxfSYzchozIyDB/NZDByPAl/7EIcQ
UP5WCRvXnx/vNS49RhY3zrezLW4slVVun7y1Ty7/l09twYm3YT3EeSKEqupV
Mbrlodnj7I23YToPv3FXUtvIhYfDVHufhfgh5P0BaG6lhpbYgNFraZCYnh2e
eN7TmZq0RZwQvCRtZb7bm8JmU4ijtGrgXifgSxJJosZzK8utWp0kPdcyaY93
mA2LhjVOBKZNs3/LEOcYeT2xCmsEfkpqSI0n+zVpeDhnUSObFBUo4u+SH34R
2CMdmHq838YgG7MPEFEjBdgEGgW29BB4pnuEMmUVxrvaL8yU0OiHTpLMsNAl
yWHZa12gGAtMC4bCLMNEtD3Xx6qjAZ8LBmW/wFkntpsy7UEF++/D2YTW+7xh
SCi0udaNodIw8GDobTufnBuScLyAB2C4VjsKMcjBTtDnJwOQdfGSSkMveH7b
hTdHRY51akAQdU5ohVbN+wvRqgyWtG7ppr7CN7NQkWdNDpnCyXkszwsLs6Jr
aLoE5bgxPu5dK4A3srsdFiz7iu1vJU51ooE06tgheZGBco9tHnxvuDJJELEO
jUHeJE9iqMWFC23bTnbCWwldJcsBrNpywNjEr5/2zmDPOoIvjSuRHlYx0S1A
ncjzSbmDcQcSLBhUllE7QXtBLZbXpMb5c+u5YFjZRlaNj9c4obNwEqm77ElA
OG1oPIC4CUHUQXWYKxQ1iWKGPbu0IbehryLGe3CTuNVGs+cb3DgCquE7zC/U
3BskDVtAu1FSdAZEakXtwMqYvnx8g+lOeOsrHzIvaA7MB9Vbb7Co1/8YEtmo
0rYPMW4R1XBrdhrqLkdjb/ROfKNZz9bWTdMSZAdAIngbQdhqt6pkAu3Or09M
H29RvwTiwBntQURMRoOXR1rYMJQGG4nkIbdA43kMKaY6JJwjCl2dojY3qJ+p
gQmUMAYVlU9lc/+HlyzhbTvu+eBpr6orSdfqU8zhiuy41Ck0Ihq2iTSDBVuT
HIAMlxKA9/0M6/TvtZoQzp4ZJoUgsZjSgkwNI+ZhqPwL22VpsKOyf4IFdcJG
IrgYctUEyeScF/gySBZteQrKIhXcxuU+5kzy4Hqofeuo7HFDXhBwFuNP1D8u
75vgTlbKwdDUlGlfnLFBLnOXpcaFG4E1kJyK9xmySwQtTNeRoGNyR0o+F9i5
TK2c1nVLTvXPn2RieGvR30/hucaxTeb3bAfAPHB61K7Xjtznykrz7na15Xl8
uQ8zZEXOEFdc0JNqLzRie+EtGSiZMOOSwxxEo0V0kZe822TUCcCd/p0URm6c
3XRYHLYyu7vnocB9tAB/kWm6UNlzjIxZxGQPSUT+zHQS3q7aE2oQbW8UUraE
wBenw+/hFoQQss7dsfI6C0zRHShnGsZLujTV+Z5yRn3G+RgsGT1lx/AjlUXC
Qge+7PYkSs/2UqWdAW8kX4004n5QQmIABWo9w+1BeEPCrMqU/Zn6qHF+I0Y9
4jB7WrAzJYy2DMDUXEg29mfju8m9CtyWvCsvTFSA4CewlpbuZr5D7YuCHsDS
gg89kAN7Z+vOORPlSaHy64jt9IvEQL3+3aLw13vxM01MW0A+ESp9yLOhSKGp
DnbAslT0ndk31OLu9iwHe6/8H2jlhsRuqmEzLmhuRIvWgqk2QJV/jm+7/F3q
PWL0lbYrWJvZC00KrEBi70vtsFZk12zm83eE2IQs6zl7jFLaUKT9nM70GDyh
nqXaR/FhKp5OLggQQ8l9mCMjt8pXu9EXd6HJnRZtaAKQIOg0WIbFET9iwWn4
jdett20RTvXdq8PQ37YPDZAr2FrN07AbaTHrHBJYpFplLQxMhym732VsZjpg
/niXDNVarUlLIbZthzmkOddF2ztweMuSwbI6dNrBkeN4lM+C9QPCXBRcktp6
DmgEuG/m/8pCQNJPXgJjI0Ri9ErM2+27X8qhzk+05NMnRk1SLHpfeV7JidKe
XtFO2DvfXyNn8DkEfcOsiCrUHG+WzIZe5navTejn64cXW+23O+bzOqjw2WBh
JG4EEkiVPxPM1nZacXZRiRlE5Lnc6t9FzmSFOJLRsdZmSYydW5a84SfSpI8c
jOiTSO21sB+RpdT9fgB0M+x9MMTosnKyVKPnMkf3lHdTlUwranm74YvxMOQq
uHokywgOHj9cZ9Us4rNWrul/x+YBqHElerYUGWzsaptyYefYw5bcO87VS+B1
XvwOGiBl6uVZK02Q2I7Np4AG9g1oWCoNIFiT4Efa3YIOc4mmzJke1bn/nZBK
pNUIFImo6kPQGgq36FtYXC/tKbon5PS/FVEiTsXYPx5E9CBq5yzCM0eomAbr
Sr1qnvlr7q0zDKF5OuK5/sUxSdvoT4qdolVmlzaBPFBtnMhZknlcQekOXggD
+dcaL3LxK+Ps5iGiXD+RIJlF92sl6qRmpkpnQr3Op1wv6RLQAPp9gCGlDEj2
U/dmr40i0BETzJ8VV7VopxgRhTf1pTuIoxi4a4uh/KLZ052xeRg0ju04R0kQ
A31rXjUIir7lT+mKewnbOts2eyDhmcs+txEIUS8AnqiFPVIhnapQG1AiZELm
iU2BksEj7Gvmw0YEnBjYSFtqi22HC2EYie4ctkhDt0i6aTAAtDUw7YC+L2cZ
wLZ1wXEFoSjglM577AS2uWebP3UCZJ9tSZnQxUhOFm5hqJ+ajNJGZyKsubzg
paajyhdZiwzKWUPDliAp7uO+4dDPnwTaMgE9ijbppYoZdKU47gaXAab+0PLh
xdKOUUGHgm9WF0OjSp52PeKN52e7bbIQb4hAm7Rko6nFxMlVXnvHsFopY2TH
YO+Ou3CzQTj0SlCvlS9wWAqOuEgPYnwxKkHMNwNQM4UFiSI99aJqkRh9XdVP
3OZDlz9XT6PKW9RJO6l0bx5DfFjQrsCjWdGLmI19nu6yXBAc7pGz4tB2MlJB
fFYECF2KlavpEx7wzQfe/O0RFlI15w7AyqrMr17M02KSa8tFLSJctPu1gBli
w//h2CG5GGincWD+xrvxCgtz+7my0yWxgOZWtpGQ4xMDUGNKpCBbKtP05wRl
nMjWr8HHHiMHJuPRtqvu8AEHrJtZaVRb/Ya7cYVNBihiQB3PkMySk/2B4IMC
g6H1Pjvax8q3aGVy3FQ6GkvzvAwp5O4gjVkvaPLw8/9vawscyoVemZnVSYjI
RdFGSZwdQwy+NKXJrhDzT10el3VajMjJQS/ISepiJA77blGbCa3uOhMe2y/F
h7MktAPM7I/AkraKHlfuC1Zvz8JzD9fIrIFwcFZ9KXbF9fURUKzhAsK/s6Yu
fXZ+ncNWhB9pqDMkhSiasLkCrwkfU+ozSZjuaV6Hn12eXaDXzmvRDH+Ra5RB
F1IiNtWGFbI6tchbZlsJxeL7b3I/ZDVOhp5HIwhAZWOrWPp5F6NYpQ+tjPhA
EcYjy3uf+fOgzFe41wpGDmLI+sYnoKlBAavn8uH6AREBwk71tAuAO6zPGGMG
OLEVu4S9i5wQI8RLBPXqKOnQ9eXrG7iLRodZNe5KczPvCqBfGTHWvXYrQpAx
1kiBzdLveLtri6Jylkw9JZkp7LfziqHFAQfWfZ6vkPbcjH9WzeliZ3JgUpYR
7DI/jVV7GZbZbdiGjTKWI6Xh8mwIR17GX12ayryqM8Z+oABK/nLULNi819at
iNNi32TXNCaQ3ethiey0JmrOwy+1mOQkrJvgiMLK00DgdycioC/DLGH7XwaK
n8Cp5sZ895DxCyieCyCgfN4SVjZD59s8Sw7gzIR0LoUoxtXou74JbwhulGvv
M3YNaieKpmQ8i3Idegrz0qwxESbis2BddEPZloWQgnIAXPE8UY78CYr0sA0S
jGnb+3GtaCHZjtxeLkvv/Xn+WkqTs5dlUuIIfOLV1AoAFi0kjy08KNSPAvnh
izOX+G2aLmbLk0v7/LEPgoG3Unq+6AT9vMbWfNgv2ucUAGQ67ujVp52lY0bj
/Eo4oKy53PY4kyfgS5A77NFsDH0OEuTgICKTcrpqTLwd4Od8Ab0sCUASI9H+
3L6DnOIANQf02R7evTdvPLDI1/bJVR36chayErfUPjMD34LYBVIRgCwBXgvv
KDibp9IUByfYBlSllpveGrU1KjkRQcxpKG4ZwScrCdjToBdKG4wbqKB2niiR
8EMSxoJ17KvzpQHtbV9jf4og4/QhI4IeEt/5/+JnlU1P/hnn3R0S0n7I4AT/
uuPwQ7dABiz/ahn3J3ZRhGt1YYa5p9u6WdsplwMKoGwvCS443/YKHiOdq3f8
nTqt970zIdVDMQHRWw6MBhnEynUgHMbPHFeh7nvHjHbZlfD/GfcHLFiqZtGa
tFfPdQhuaZ2ixj2XIg9lzS07PIbqsT3mx6vm1XZSpmPy5rBR5lPDs5iR12Wd
sFE74lzbNGre6EtSv4wx0Bz8+9fwl/YyAxgldxBlbustiVQM5vslNtiNPGF0
ziV/vudsMj9xNyR0cfEbX5zWC8IAR9wt3fT3ffsdQfjgp9Kl20plhpYM3Mg5
NaCxJfUffnyvB+3LKvyKEnr9/BnOxyN38AafRsfV870mgIIbwBGe4wuYNm5t
ti5MxXWZ7KG/FKW4EwCMyP3P41ak0dJF4s7MNfM6aDAeI3WssZVr0SSWurlF
7tXbiCDFs8PPDcXPyfCrksTXRCBgm1WsoUSN50ipCfdIGUSfMPs5YPmeSgRO
cS/ORnplkOQs2XDDKTdntbd0ldsU1NL5hi/gcqytjKlro7DNrMoZY9Gf80o6
bCkdKsTu9TXHtdiFRDvWEJ/Fk4wdQGL532M8O/Cawcc9tGoqLkUt8DvzUp90
QWFkMdv5RlQ8vyi1R+9IAU/iJc/0dhrYMrFh/vCFUtcZzlufz+B2ihns2Owa
zt0cLM07VKNLItx0krOybv8jtH6xItmaQojFwJyej7qrbkZZDztVyk9qCmRK
xK6AB/0uVskmskVFDXLmg0H99WphrSRpV9UrnX3FstqxmwOctsSXnHqPigGp
pK2dT4NmIGBnhFS7tOAsZn4gNn0EXJSNFzUVXi+kVDAii0gScTyfdDqaz6/X
8zQ8BpB5gLEHI3Nz9+/wmPwejEwol75KLHnAg5BJvdtgf/Gk5NjjtmyWarOX
nyaYqclkeQ37ONqNE+zvBQP5fRVjWVznSL+nPx7x46yf3j60ROz949ZyvGmf
pcuMjfeVG5JcbCPjPpz2wzbRAOIRL2YRLKej/x9+80Jv3oAFf9sG8WBQkgPa
MEXyxYgIjIXBtaOXzm9jEMoWbZsyCQiCDqePcir7u7Gj4o7cq7kSp5sxDbKa
BOYNO+1unY9YBXe1MThgGM3uKZo3lDo4kmhIBH0sa2Lux87tJq8P+mLTyk9P
J9K/He6S3LfibWM1/s74tHbqr/G4AQGrJGTurp/eWfWxQZJIzQyefBUsC+cD
7lcTplcTPtYkI8ti7K3QdLgZd1RkpNkxbZy4HG4viPJUgx9s/acJIbl4ZQCE
0A9/ExTmoAS/MHEXmpZVWGF1cAr7ZTw8O9bZU2+vy9w1lWUMn/IvT/jrWog2
gahkCqjJTd0ADTDz72rwCl7IfjuNybADGMe+5kfOSBZ+LFniJ1KF7IBubkzy
KHiLNHFJOHKWSsfYLztb9AU9KaxtWQ9cuIeCg3Rha/+Vti9FJxPoq8YqsZMo
j/pYpfkAln5wfBtSQvP+SRmuCg7RKh8JqapRed82GupeLcBc+XzLW3yc/dP0
UIceOgsP7hphMOgtUdYHUqYHMSmGdxqPtkAsntjnsVUMvEsImUDX685qTtA6
rqCbAJQEPu5EOvk+D6Hv2K6QnCpdGCsqD4kJIy7LHLe5L4d1LnUzlipplKfo
QSiJJOg3SE08c4hc8DHrgRUuLKfX/fIFZxu+7XkpHee7aKd4lx2cVP3GljoU
OSOJMOghbKJ7yrSoE7Jn+ioPAvYjXHQR/GdFASF29elsrXHXvphrC2HRg43X
EYvph9dDDX3OzeYxOL5rIwbV+Yv10Da+8xQs+DWON4KxkuMa6ZpyEnHVx/wZ
/SsX4kChI2csG2Xdmicj9MwVVi7v6D+HG9nV8jw758Lssmr05MWouT7nBSXo
bmNSbuLhaVR/E9E4YG5JSYgfjh9Ixv0/QUwszpg/70vgzKGnq9ShA1WaddJ0
Uqhb38Sn3zlp9WnO0JWylXpG4JxyeWaYdGBsOV0ZZMjhi51y1CVQ+kAkmcbj
yoEuzlrPwIOLTjdY1ZeAt0vby2seiBB2RBJmlVZAKW3I3gS15ZxH/MMYomRq
GLX+wZSNFVE5Zxj/awcbcTa34rI31iGHPIdkgnRe+kAa0sRpLOPB8ULZYoTc
KRO+ZOZZrqfnoq/jHjXHyc6FYJdCjY11FJwmbwZBaDXIHAqRq+T1x0D77+6r
86ig7TXxxA5Lv8bBgAkI4PWo9iiEC3FpmC5A/nRllDcaFKeysLYNXjQoqmSl
lp6pBA1kQlpl0WO9Ti8adZYrmcJ4rVUjt9tvrLNN+4Ny3z53dlSK5HUS8V9s
3lOYOyt56GZ2TlsEZRpUtvsfYbnSYR1Cz8r2UXGkCnn3fq+myNP/lIxkap5G
UR4U6VuMpy+jRIDEerXVUNG9F2niclLwM9bSaM+eYQNEOcMJCplhfsggFz/h
XbTUEJS4+NNPNiu1gytfaNpOtTSC8DK3IS1Ge9d41boWs/YqV6RAbl5oHYCj
XugSa21n6kTynORJFCHF7ri0uhqmsCeI4gkVp3kiGx6NPrJyu852w40Y0YGC
Yb3jTljKBe3TXLGyJwX4upy3cnGka3F2KEO+lrPMQcZjOPoUTKHkTkpsgfoX
Ke4jZvSYGzjzDLUMJg6uty49X/mOXDQPJ4nF2hkLViYajfQc0IqHPyjpenlx
8OZGAQr8UNL7GpBnkZwLwBieR4bKq2/M29wY5S1s8S8YjmRsaC/WqA6F9iu/
V5ZoYiqC39pL2HAuGTvj2TUppEOga9HAzOGtht6r4YqC4DTnGMYHDYGnbCCh
SJplAZwTVAOZEi3yQelPOwjaBZgQoUlpROEFfuYyzRXYziEo/eCCVlYE5mM3
lMt4S+ZLxd8PMb4N72+AP4yDCYTpZWZE5hRx//Ho0Bl7nMKEijb6kB8qGF1s
rOZQqpAoOgW6soE1xt8qK1gwaPVI2gzKKkC66G5Wid+n0SllozDHCMEBRX4d
YD59ONFKZRy/3yjWtS/pbJhEOTS0NLVUMPFo+eSi1noJ1Vlnp23psftj4sNS
82MeyVyHyChZ4RRQq/O4DxdlX00jgRi0L+etxGv2xQarQ0xQlXb/wA5b4EIB
7y4vEIpl3ZCVQxdMtd91+n9GVJsvYz0thozo31mt2/JXFh+Ftj1t6CK7ey7K
IXklpHlkEdMAhLHmCYpibjS367Pk8AjtuiWyyV5FRp0zToC8F8Ko8bEO+nc6
LbCCr5QTLvjY8mjgo9Mi22xgg3f+iPnaE+FBOt2Vs+Ql4/cDYZYMcAu9QHgI
J+a1TcuLUQSiYh2sGAKCp0Cc9cMjaZUZqFKxAfXQK6gu1hd+JeS9e0IXIXXX
xjS07IdpCsAyxbofAgt8qxqf4GjLQNXamRKU3vcSmFxZhIz5wwk1xs+nJujr
bKwKqNYXbT9KjQDLd1bKjjrbkiyO6pXfrlsIHwwxIjH53FiwxdEhArMcEpmL
/WkMMNMjwvmGfFIYifTnmLgM0sYejXZowew4YdVVsfYx+n5Z66gwKo/XHGwM
5Dto7uhbmOCblLz2Sat+nqH40ca2Z+4HnKDjG/wI3Gd2DkUPH8HQEu4uS8la
tnsns13iSZUTHefhUX6RmGewU9VSiHTPss2tVkNKhP9EMvSqrnZ+pFjHrggT
9CbKuvzgDtRKwVXTcn0lrt+5zV8G+2OJty/SlyAWzDhQx1CYRf7zTHy6gnkv
k9WWOrCvgZ6oXfaZvdVO6Q/EGmAWOIDybAq3yb6IP7KshMHSgEc8hYXCniit
34sjGe8qGXVtRe95o6r/AqhBeZauIXeYJw11WWggEFsZbPsMSJP4W8T6OOGx
wFUT4VLwtLgWBPmaw/gYug11t6e+CEITZLh3hdOXGkxTEu+7TLixHH62yOpG
KtX0qRJf+TDSoYqqeF0S7cFTDLW1LaPmePziMcptytmgaIvHTmm60CIyQUZO
0xbptZ5vzZ1n8Kwfw5l/+uizTcaxc14Ba6Xzu3cbQpVF/1JEKQBUpmRLHnoq
Q8YPBvIIB4g75SAW8uMiv3S0GPzoyU1eqyDY8UGm0Z8s3x/zXMyBxvXWoWpd
8qgcbbLv2kFPGFUdDlEpGVIrxo7P0PKcKCdeWY+vSbPy/jaFC5vZVnIbXanZ
sh7YuaqNCmoXpT+W+EQ7U8mLeYjezeztAyvzH0QD1YEMN+ZL5NwAwtpVTsDC
Smhy/Sj0SmfebsCmMxsGLsYPkJqW5TZRBrYq+V6xMFXTOphPPCaR8vOTDUJn
8yLQr+6JJmes4csI+Qi0perB03oz4kzYd4lx3Da3heASQW2SAVBh4nohl86/
7T66UflpRSUD49/TpkyU62haTZUxp4ho+7oFcDx9erqNgstNklprLiPNdXaC
zfa0Yt7wwv6C7FVysJZ71wJ0UxsCF8tab5IzshLRb0+f2mQYVNmREWdq3haY
xl89d7HdQuElEp960zVHNt+sdZj5HePUlWY7Tr1WY2Sq0sH6xTm9J3QUypQZ
kQ4n28HAHhDoZERkKousRJCm2W1pN+jF69sTPZwZ3dyT94abM/x3mWCtYhz7
ELkeSX5Lilzoh+NvXHZjjkrrTBOMo3NCILNw+FsCeecEpe0EQsErMrumTAGo
+/L/btj2UaBS/RLk2+WHHFCrEhcUh8yLT0aiURUjZqT+u6DMkkWNcPk70Z3i
ud61r/7pZcIsXPOGHwm9zZVNXXc7drzLgkldbquIOhWgV3cf4/E/5pf+CpxZ
nTzzp07fVw3IVr2V+5CdQeodfHhzEbBGytTu9VKVptgJrm7Ljm7hbNJ82IRq
zFBAdJUGcB29LVA7Z7ucp6/s3XsW3nw+W7PAGjapPfIKxsTj1ShkC/O2+QXZ
6nObePsYmHb94AxAwp0RtgkfrzsSgev6bhinAc2GHcp1CAsXe5wUv237PapH
eGbVsyTUFtHy84PFUGbnN8XNV8vXNWTtpnkL775oQgIkMKj6CEB2mTI9RY0l
aht6pGE/TeaeyVo2JdVbRLdookRlFkiLjxAPceO9vEFwWvQgC/N7bu9pW3GH
mWrp/UNWJVICLUCfJo9sPHQnK0Anh+mvgVBX6MR7goGP64+9Ui6pHWARCk3r
yKFtOYGLSo2794dbrmCA1CK9fvv/Lfe+Uhvzyfn2iGjV9M8/sRDXIDFcohdV
ljSLdxnFNlKpjSNBXr2OpTd93SyVuqymCPKFHIjX9QbFO4SsySp75LqveT+x
wWfm+E8SJ84gC9EjSx0T459QiJ+w/LgkKGI06SOU7wJZNycy9xGxa2h3Z+na
UM0lC1IaJDA1Z3D+gTylLqF67tdMFnQTVBmAkRcOy6VoXKidSlgaA+5Hb0Ou
BSXLly4AubtxxSRbjOFmPrt84rghcODS4WXCeU4oxSh1Gswv2Id1iseXB9GZ
3q5cDJlni9DCG86vMYkNuEHcBgbAzEac9KcIEMZUXIQfLjWo2FAhsg8lSpmR
i9Zh80M3NSbuqeoCpQpA+LgJdxO39fQaN4v2G0PLWH5wX5EOQQGjjfTb/uJa
puHKq3Kl7EwJMgcR6QUX8zTGHkHk3Q5eIucgIjZ+eG4J4EQj/NWrO7F/xSzv
ptvmb3rVRFPYnJ2NEJZRukA/sf7OUV0+gf0PsHuDTvjhDoLGmGLE0Vi9c+/i
qa3tX7UuBrNlTRxayWvkmLHmabqZjb2ZowEnf43L8m97WNwZtdpLZkc7UCtw
v1q2yckv94rKR1VpV2JQbkyoxa3tovHtUiHe97b3NKstw2//32H4k6MqZGHG
TER/Sp/hYSgUzqoCPFn8KCS/DnEFOhbLnj68a5MOQCkeiaBV2W3xszLWs4FQ
37y7QqYNaJrnECAlKP83lMyLrW1bOE5EHBB3JsFoSg/DxXDqSuepkzPfXatD
vUploxOZHjh5+K4sLTtAbMwmsI2OntYcslitZjzBxy03ShBs+g4J9c5QgzVR
NRCBd8GhczfsIf331rQ43bwjFGytGcQjC2xAza46jh33WDVajId+GuyrarBe
/ngqvpE4plATX3MwdulZp4TlR17l6/OMxlT4didhlCJ7FWCsDSNUYyongEpk
QtrT3Bvxl5UCGD3nnSx1SHYRnUas5/UxZkKc+UFZaeZD/GbXkiQmZtruSCvs
0DTxwKHxWHoghJtVg3QW6LpubmYEdgqWRP6VDaOnmhcL+WTI0AXirz6JX+dt
jWQlz8+hyHkLyYrmWcotNjUWlUbVJl8ceOWzFSBp02+g6Jk3yUDnTysu+X5h
zWs0KOmZ1ywCPiUDcqDeUj1I7cqtgBbZafcXcf76QUtD17WeCkHJYiHdMe+v
IOdWSlsZXkSideBaRqXouaNNzfp+A5hgDiYrSYp2EUR2W5mzYW8IEPEcbwsb
9lNrZEfIf4AaZyMWJJVQ8NQRix1kCE8B96l4CAPSluS7HeYobqLxA/hD/CaL
SFkhFDNpk6NouebOGu1x6h45ShgZEspjAoOZHL03c+jlOxnOkrSlnyMUBF/D
In/dpgqQ1O8Ydfy/cxf81BRwtJCoDOSsr8AB3KXTRLh40BT8Ayt9SG/+ZvJZ
wf0d8knj4vD5CwVNMpGfFxTaAuE13wOq4Rfdf8s0KPOVqSVPomD66FeMBqOo
ci9j/57pxR52q38yynFm0S/bJ2l+FLa6BhLrgS39yH6uizatxX5drSRHbQEs
0prAkT+r71IoMWAZx/1psdCDhSbF5IepvPueYsZoLMWad8LPR2t0xGJcjZg0
3ma30hK+apRs7JgcZv9uepoWceDFzaH9N94rXzQ6mD9hb/P2iHtOzbit5/uq
jkb7zF7GKntEfiuYhvI/QlWvST+UHqDMUc9eA+2DSjpwvrt2Xa6Rx4JEQ8EE
giFkcnBpo7H3yWyW6Tpgx+9qszRCsZMXntnxF57jnZsY5XSXEnL8t+PRlPHm
l9lMmV2zS1Yr+160UKrOFBX2pLcaEgHiG6vJr3VNHWZligSkGBFdo+DH2VOG
VWTM7d2qzQVeCjRq8tiJxMo1SCAi3ZV6wgKHNbCnj4B2UJmGg7OkrhqgsWhM
/1fUZ2HGdwYBbFadBXuMHOxSCgoaUm7xeD8+vnJ8NqFsHvzXw+7P7cZEv6EM
7zrhhHYnz3qzfNNZ5IVDHduP8nKvHf4vBLGxt79+3KsIN/mnOtctpkkQSJEb
NO73ZoyCpvALSQo5TPGrNoLkwxJFHET5g/3afl0yEXHc4QjgmSyxMAGgbM1b
xlwOlOv/vtfW8kDafEDB4Ai9trq4oVIa1hZUjYPQ2g7WedKvrU9UgYzWmJd9
zQNrDzZA9WX44QUfmzRjstnmf76VAM2FBYj4XtF8ROcnHRhcnzPVvSu7cOrU
irTl1pAvMjemwZ+QuLNG8WdBTQfXnecOZZCZ44Ac90/rAIGAEsXXd9wFMAtQ
npNvrCRym4IzMycp9H2pEF/jcho5BYaRQAFNNuEzR+NZWDA7bctdUc3jDIZH
NvGJU0mGnDl8RDp2vdbXkTCYTWXg7uyBP+gawp1KwVU2v8yGvptvcpj67GVp
SwKqABw07pqYT54s2vj30wSZNslM8yEmDTO/lU+NiN1gm4CAy2Kwur5aBVYB
5v+YbKu1vlCC30I9/K5V9nfBlZYzt5eeOZuwt/Y31HAOZ8ZkPWwF4s4li94H
oP5R4IxU1V3WICFrFOvtLDwwdHjd/5t7cvObB3Cpt3MjPGDZmoa6rIdvJPnI
674pxIHzX2DR0P7ir6NT1PdqHByipS6BGZowvxVKhQDNmZLuPuLF3eFVXk30
TsiSn7IXH9mr2Ga1aXknYUKxtuCjlqUg80yPbzkpM/UGYmeY9OinJiYcK9WB
Z7rvK5xOUwz19VMXoa4VCwqpQrMmIhTK+Db5tUz9GaA+Z4yIG8S5lhvZ1d7R
3prF9/9iJ1Vnhg+EM1ikgWs80nU2W3KlJlITJpIhrgjZc86+SC2Bp07O1kbN
It5J9BiF8uKYDjyV1pDY0UjM6y05Z4socJ7xPSAbRl0abElwTijaZdO894bs
ZuYRTuTctwLkdolp/gDvXdWKyRXGessAjD/C19v6Lp0pblOXidSH7lghhxyd
wCj0LGzZj8+mz2rn+WXfd+tNdkay56Ty5gw4zFFw+Id6Mfw63o/pzVKrnD79
+FjeFF7g8pVG9J7tw2gdLcqArH+7bWXd6LNQMr9nNYk+zU6lXcuwSZ5WznAK
ZVGsZjbiKmeG0WRMzYNW27NjhGqPCwzRxfWwgzwhQ2gdhZgub462ShYXFu/H
5dlOueRUBJAMlesfI+DnfivKlbw2TbxW96svIfuoRzBhBMQd7scu5hzBnO6x
eFGitNztA3T7kt0UZbA5jdlH6PvSbKLeLqDw8D7j1L0uBENLGuk7avkaBRKF
wbOP/R/AN22iLljA9/qAJ9SOz5oNzpqIbfSxO0TkPgRhh4qnFU+hzhUswK/h
w+yTwd+VyUM5aJbM2o8JBTAMk69xwTETFAV0PZXmT6GI9OBtLPyCNgEGS/5d
bETuDaPCFVMcZbXkuyE0Bo0EaUHAvWTZOKvMtoI+lUkHCGnYkrxEtXmWSskt
DbkOlvOYCSYPLRpSIDlRXnWR8KTV9jTrNeyLeX0kvrmO92cRYuNAad0r26rM
FMv/2W6NKTVMh4PulbHgpjuyc6CY0hzWJx/yh1Rj3Zy37S6cZ9CP4kZHMsgw
hUFCQrxLMb5ujdoAa5GPW+N/HIT4/ETGDEV/bf69n9eYE2/AbYR8No2UZBzD
WIf/Qo3Aa06WoidrcnnAOELamopzbZ5huqSAonV37wvxQ7ARs1iHcIZlM04V
9KjagtXyhCVMiyiW3KaWxUHBZRJ2Aw02ejpJpGdUsb6Aqe4dJqwL7at8uw9O
afbogq03+oxDLJv7Ym9Vy1+DqQ+1lpVEDtjkuSWMI0xQVssKwgQL+N4Z58kt
KfVexwFMH4eJEvYX6k4A97Zwjvkj1Uu8hPIP9XB+qcMqWBRFIJw2RhqLg97f
dEAN5COIXRxBG0rAT/2+68VZfrCFSS3fHRK2kXc5APxZTE92ezmvAU/lQnR7
flyYORkGLB4Fn1XxBJJqRoxKyQl9AvAUW03Hd1PtbnebwdFSf9yFpxJGC3SC
5OYkGo91cKvCNkh/FfZ5HD7qCdJJwR3rObjj2xKRqTnDs2JwPKt5Yzu/1+tr
ODtJpmd3A9/nbv0wUcCqvO7QJwZTg73071WYJffP8uZ3yqJxD3SZvdJwEBcr
KRToqwkcV5T1RRaACNF+9qDAot3QGvFiWlbjKQ1F61yEd4FKO3u0e2o6ftSU
A6R27I89Q7XFTqxDA57KJ8XS1kRuJV+qZMjdEasQFBIguc+iqmEQC/3XVWAA
XWzy1sACEYQhBRhl4ZY65P84sh714byLq9sxtpARP+cqnYf87lGxzUcVP5PU
MIUYdv5oTzMvDus/C8zhjBRGnJin+8e4k0BZfBJVE5KaFL5ioXd2IcCFpse/
8CSghn8DB/2CGLNq3tqC2T7oEGL5j3taOln+ZlMuoT8zgtp6OmoPB2J4hSED
vxuUfqD3yN88Ulq8RIRmbWOa7f/+YnMUEbjRxxwjMGp0aHybHZWAt5bjLphS
2xSsmVYddaxuO0tXfMw2ZNjb24hlgtOQwyHPQuwFEfq9tZF0zsBYBk+3sANh
7PBe7sui54Y7ostrtxsZ1tPS4xxF/qTXYFAlOHrn/yHTN5Pkt0NUGhY9WQYX
qHWwvSSrBofZDkkyW5rWkM5nEOiYgpXK5OxHGZMetgAZs35+/lntZ/W2mVlh
iCseYnIcy6BXIF8bLP+Uzgg4yRYqctFjnQLTeCo9i5xKtB5gjiiVuIitFqoh
QiFn7OJqX3IF4sxV+DIggsOLrGB2gzYznya+3cZr3c96aUAHGFmf0ZhTnwj5
T3TqsVigsqOK8AwR+EZJ/50bC4SMUHBgf0GWLYgKUH58CghKL02jk8Hpu+K+
eUE+WpJiv+0dyBUjsz/10bEjKp9sn9iPWxTR2KJvBE2JAxQdVsIu3zbpCNOD
qWA4i+CapmcZMUM0kK0FbMfrpn+t2BnE46bLmfYRuVxXD6KxiXdTexC/xJXE
ireInYM57Yn00d6GkNbGYt407KcCIanPvmF6DmSWDT9x/eZ+6T900dmvyggz
C2nisIxZjwoVPE/euX9wEAgby8a056vqKamIulSlsS04aA6htM3sHLy17oQH
rPLdUcoa4IHaXWjPvY/dOwD8jstGjTaADn4N+ZSn8SXQgwQk3ICvWJOf7s39
PWWSyQUiL+f5F732xyk1xEU3m22syyr1GZjfBrWij1ATSBHSyZw4zy3G2UA2
4wEDNc1diKWZ3LL5gDLb6eBhoMlaQaIG2qnoxc7kRpwQHvWNmFy9bA+KNRov
4X4eNDzFA7iZlBlJvLQOQ6VjHJRy94SPURP9qog4HO8UP6XmG7uPe3/LlCnW
0kQmhsjlDYkoL05yPpqYrtGuStTul3MJ9ufUZKH+Pa0onYuEowKv9plY4snm
TQX+pNhAUOu2YVZaG6uDdTlbOmgBHfBK4QJ4j22Bcv7gGkuV8Bn7L1eCikbS
RrvsTyd5MDhaLR8dyRa6iSc3aBqUQFCt8RpA2LGPCuOPgyXKqxPux0Zn/lmw
P7g67X+HLZkntn7EldqipGBOVpaML6QGtn6h+jyAZ2tKNf3eKhJS55IbBPCK
O3xVMwSiUg2IqXvHq+LtLHo039zgdPtgI7DMnNtGYbGdAP9d+nHgy35MOnU/
jCdbf6LWhl6vPQX2G7aMFJklWnz2mNYRwcl8Tx5FUztgBmHPadQmvA0a/ma9
hAhk3PnqF2ly35yqeLS80N+l9MVVnRsJzSEaKQoHrEnwB9DIvyo/aD7twWTu
kfWGlZfGqB2dG7ypspFgIo8JaA4rM6xvtM/Ek39rx2fdjiFqegEGFuWuHE79
8tKG0NyMd8TeSsJdi+xeu0VtOvwIVRWlvj17CaMwONZGAIF2aY2OfvPcqgf3
0h7IwWkKBHT6wxmJuALmIbjThFBn5f9Rgb7STuUBXmYM9Dre7q6fH8F1tnd2
/Nj17kYwqlCY+FLj1ARE3EMx7MTbugU2JlzBjaE6Mf/X+6JBRnFSOMfYekjS
iLNZKREzNsJBIjAazLO2jADgQUrzX1DQIz2K57YGLkSMkDGXXr0P2gxYmpPU
q5FRcmWfKomND81NAu5yNPL2hdt3y6enhHzR+djMLljqyczc+F2adYkqvijk
OU372uJA5pQ6wwAnvH3VgV3nxzjNgsOyB1XPwRKSVSFR/5XCoGcbPQjsmpJv
J+j7TGskB1gIiNYfCxLnl34Yr/N6ajhcIwSTS1C9uB4YfPz7x9682Klbz1bq
PQaRPOvmjTt+LYS6aPsgujN4EStef8KKs1swEYnm4vJVXQLIQ+ebSje5DjzT
UlvfQCiQS5DtZi8NJiVluUURyAs/Yw599STig95hb+nUIPQCnkGW1tNz/FcC
GOuXRbOjdf/Qtco29FCCMnWY54FYBlQbbJHMjLuVt9Lr4FpZyeKVUL9YVy2x
fZzrqxqmLwxiGM3nNZJjB/SclvaEwPOAEbBkSM1zyhiTsymVOH34cHlmWhje
B4+GB3fIO1GqvzHxA2zf+qL9topF6XgPiKw4gqA2RU5qjapPShv1QTTtAtsS
OI0LCjHH1WxZmXVAobifT0XENWAOQuysVqcONcyIncyGbjFuFTvvZlxhlXpe
ZSq9eLkVTj2c9Hy+1YB6u8A+0NNqWtIO4AscGrp3Ku+IoyR2TK0EsRlQTDCC
N73EEApiyXybqUTkWv9ahn+vk8tlF+e+jkKcT3c29j3ZVeq7HSh83Xf2s595
az8rtWAEf3e4IIJ+RtBUqFiMV6APnozgz/uiDdLtkZuiUWsPwfwpc+OBvIYA
m8gpsYxgGdt0FzAAB7aylK7gSABXzlApuMm1sK/glDtRgiLLxTKF1MKGVhDg
dR9Udamq+Wo5ySkU085dAgcATo3hBrrXDC8A1fSOity9uw5JsoYxLM0I8lMG
NR/pCpRypE9zXgAnpk/+Lk9KdWchHJgLKtwEOchYA9HAM2bq9ZTvhDcGJ0Rv
2P+HyFguXz73b9cVmhhc5QxQQsx8Tjek6RpceQAX+lQhn7CPFIdkb93kVjRw
uYYrici+zwYKkeYe7URctGnWeDktuSb9DqIosjN+8mleqKW6DvECqclzYZxO
/A7C7tgRw1FNoYQOlJSax0x8IUEg3zuxSj6skcfnzNCQcB/7LyBCdJfPkYfk
l2ckPPuBYqIoxhDBf3CSkXZIrcuPGtNsPBqhwwvC46zhey5cmKTrDO0HpYgY
1s0xkAKtaKQ8a7JlYP9qzjMer7zKr7ZZA4XFP/Zilwi4K3AdMNFXp2bvAO2T
24SwDvT5xZRPDC/dB5hb8L5zT2IdBvXsbMK4Ce3fCeYypeIwwjHZzqk5s4Zh
NcGaptZ79kfkNLmAlwpYv1D7H4w5t53cu/PYp1jj+8JYJ5XSGZNL5SKRrEpn
D3n94AWj+yJo4iOx42WD+QSiDZfcVfsqN7pIXURKrbnZJlpR+WFHQ4c+lQYI
bnQ1anvnS1YsWRU27XWMUV4O8HmSVRxNs8PvQus6TSODvEHlLrXXI5koM/ND
aJ+RKPXsnjw1zkYVVtSYbaJvtAHW45RT9sHscZ2WdS/TZ6a6mE7AIlJRpcMb
KdLvxAf64Aghydl1jT03u8nG+iOHUhBcHTygQbqbX8+jhPkdOYBOkQsM0HeU
NTVopFRx5QXgZC/iGCqnCF8ACnqn5zoIgRiClOPVEGmVa7Kd0GfOkm/IuctD
M/EayM0e0r/mufJpT7tz7h2IQIHjB85WGsA8KTrEcyx/6PwUzEcIZNEmo/oW
0Rt0jpVYgZrthqHd2YMPjf36vwUWxR/BubFXCuM7dn3XPA7hr7Xoj37Bj0In
FKUYEWpQBOXEGt9ZdwsgDreb3JP9l6MyCMSRUBbyM/nFKkSZpTr6pEbrDP1B
QHBjSKJh50lPXTSOSbdJyj0fpIqA+mrVXt7yTRUsiGWjg7VEK+vBoXHG4bQp
h0ZuLQURbuldj2I0kFL0WLiLKZ+Ch2bB7ygbvv2PFs1/BCqnNIk9n7gkFTTJ
BbuxwPB03nVekiygeZmQ+cqGubFgtX6qes+hgT5yo/CTnF64ZT7uN+4jtLzl
65aJAa8xzmx1JMog2bUeN9QfeXP4jQDoI4Dv5YULuOcvSbLl8gjyAO1deHOs
2ywm0hKvsXz9TspbrpNI6qSLE7i2MOIHv9UgXJvcUavRNuGdg2eZwNhaBEX8
pLgs/1SAMSbsjqPdTg/HTJrEsYFYORB+AGqvZ3fotrztGAQWbx9lPMqR9xmj
IdGSVhh4ytt8sLDsOnl3dAYKhJmEHfUr07RcFtG7nq8OoRZdHs9GUK23BduZ
kpPdGs//tnEG4IYtSZydmngKNCCtttbvof578BTqaEYdltMXrbGNWcV84VzA
N81OyyG7kcO1leHsYjjPzs0T/L3uLnVOK9w5x5wsqDa3xAyG7QSycT5NQI4L
UToIcklnHyAX+eJcwOc4ACKYHR7hDA5GnyDZfXpnC2hHfU0Q1N48Yeokbq9G
NE+6z53CZRi8Kd3UlKOV/IjOSonDAXsMBqzf1oYQzY3s0rchtXJg/QpejAB9
q8MVaV5ixONz4IYFt6/lxIUt4XhoCZ3svJk7nR49/tnwyQC2QGPjsmi4bTxZ
mMHJuughqo63snSvCiY8ecxbNVNrwLQc24vyTll8yniiWcWjxLhtIzi2PMtZ
OuxK3P3kdrE083w1PnLTjP3psaP79ilbz/O0CuJyrp8DmvsAeFjjLCYl1zPW
HkyApaj61+z01V8YG7z2KPZ6Ac+qnZgFwTIl6GiqN74V1RXuP5CRQBMfbNxz
9mbiFW5O3u8mW2T0OKOuVLfiZVkF+v7X6jzQsIu+a8ZqSUEEqq1cnAylFxOP
s93bs4SSm78OxRAIBSHHedixYlVhbbHqNtH6KNfPJEB4W1X/tilLg2Q5eNlR
+BvPYyEj2g0TBWSkVntXhN809efmyzCf/bZD96DkKRzmmAR8OMMgSsqAEPiR
3tC0eK8BLuFau2JeXK4J2lYsMHd8pO8llMcDYbIe6E84EHM8LK8N0Yu4QwDl
xwb8pljY37+rUCZXMfih1zWObX/XE71K3RTGLVA+Hh3vA5FtGs45z/kNHjgt
jAL28EfFgaEGOD6JniYJmw55EGtSwxcOy6iKB79E8xO9esIDn0w0oLUvY+d6
GfQdaeCh3OnMxK160z4tMoqNY5cEd8PjhiyvexJp61qxTFHsEgBw8BW5hgxd
U3ubMcPpE3XZfNPSukJt3ZIkS16gpUVK5tpy5tOrqw9F2OX+Pul7AanN2+Kh
9Giod6h0DKaazAmhSTMfe9+Fmd+qRyx9MVkXsrjxIdty25wwnBrwJm4u4aZ8
KJMAoQfmPwKPcEKfLJmdMW+Usy5L2F9GGI/kQ9c+aXQ4lNwRx129ioP4wQ/G
eygUMDaYA9eZBqzmcoeFopPOc7lxW/6bSCBCnywu7xMTbN7qbXiKRlsRzdNy
Ch1RxFUdWm8i+0Br3LkvWL7gcRK4m42ZMRZSbNzXUZOw+WFrCM/1qBIxD8ur
vzmJ4rqMBnyxxOuHlTUOkIcOCT2zUiXPZdzOTkyPw4rtKUWnpKAVGAZR3svR
qDq//sCbxWjWM9sRxwmKzJ4WqburDecfq2DqOLr8QR/VS3Ycf2X3htHJfcDZ
iZ1jwXN4UsbPonXcykN2DyCvapQqN5Mb4VZvzSPC3fl7kv6lcqd7e9pqDIJY
yb2ih9jT24zAor5ecjlN3cWsTmoHqcK5c8nxVtYq57Zg/5T515prArAc9xE0
yxXo9yhPxJcreuLBlmAcL4hI3lx1yIes59IZMtv/tiY0jibBpoImj+OpBwzA
y+NvzzoyjMsInnabQwGTVO4AkBQT/nTqy0W+Ws0zlx5SITGJXIe7uR38YWP8
jdw+rf8OK31RmNoP9FpwoUU28Xq595pBw8IRx2+mo5CSFNcI/NeM/UIhYspg
OA+SlkAiWK679k4sZIj34yT73oQVx2A9UpZg0dJBNtT5GEj2u3cvjJgQI9Ly
tgy7fb2kM4MU2L46bcJcMskFixCnxvl4PPduiSH4UyZdwi4ey2tNNEKSL0aP
jr3m0e0fGEEoV0aQ2YhOpvEv6KL40hbX/Jf4t/vRQKAXIHv/R9j4AOFclpu8
G/GOV9gDs4UgeGKGquq49sZa7cEfmP7KjHF4k6p2zT6zIQV71dU1RG/o7IBR
0z/IX1IZFZ75CfqVVbCt/CyN27SXDR9pAjLfse3gF9wmIkThbq4PKLyduoUO
G6r4BkiEkgM6q8gK9vWwpF1eIajAyiHeGHKIBkPCuN3QDE82QK67VZELuqpN
+wJINGAJkyeV/Lrc9YL8FdY9n1twJBlir85H7d8wRSdRMrBVwVWZI3nz/mgi
QGtU64ln1RAZanQaGb6taUH1peTRAp8Un7iOjRCPB6oD6PKW6wBOHB9HHfde
k++hwSC+J51QWeX9kH38IYVm+Ku3UaU6/Sa9xRuZm22/IChQg089INOYnh77
qHSgsZnqBnFNLis5baPnIqFNEa1zN72opQ9CGYXAlmYFdz7Jp13nYVXCSCvr
72M+s8lMrsqa8AA7IxgZrtf1/Loe6CiHgoi9JA1oKtBa36ViD/QRgPGd0KHK
VmDH7vgiE4jSIC4o2hrwDw+8cqJQwxWKgBrg5C1XU0APIv0jQqMeLs92WiWO
BiyCdLIVowtKOKJ0DU5cIoJk38FpwOC5V/mPXe9zEe9LZHonk5d9nGFWR1hw
OZajn+zpEf8dRiFQx3YWaAa/OLi3IvYzt5cB0RMZJbOADqnntkIZPy0IlsXt
JvaxNxHOkrd+eIWnnrOwhqgn6IXbECbbXwgdmMbkZGfFo7Vyr+JRGNcLdZhz
85eCpuovRPtFOtIQhdsNWY3AJo1C5OWHuJPzIx5jwoHRio/9HV55rlsaDG1x
vsG1GFbwr/le1XfyRgLlPMfabIjJNfaplX5Ke21EPPjFr9490BCY63TAHLAK
03f6xxd8nKKrXVJFeV8acJiGSFAq+up0tNVZw0o/h5KaFK8cotyBZvGtRXLI
rTlTdB8KNMwBNLuH8/MfU0a3DWJ6v/m2h2zU8s/zazI0gy9OcKMKYRSr5ao+
JlBeHav0h/9a+/lU4qRDMg/3Yoe/1g1vd7UizsG5NiBUT3Dz+tDf/61Y3Cxg
yxyABvg08nDdtba/DKNadGT4mRxcgPZJxf2E+GkqIV3cNtNijpqle4Saf6Fu
UJd+rzNAiRrBAnXwjxY6WDqc/SrW1si/ulR0LWI84B43g2izwLNIvgZO9g+6
34vER1qy3SmYJ5BuIAPbB+LpLgcGRRY3KZPo6vQUx+sFWOtdxHbIq/HfmQVC
zuc9x6IWC+bexqNb5oTlPfwgJWBipisXeQOy3qaoyJxe6gDMIF/cNy7aHy6W
JXMQj0cYr5X/7XAPMtVDcNFuwHrsQdUt9uWLPdFEuJ9n1x64HrgcP2vrDFsy
qeKiH8lmOD22RAjwL6kDcK8i8VHGSLRKtOqjkq/ONvCytez6ds4bxoqP8eHn
+mBoA5Pt2aWurWdcA7mi2sg7usYqFDadfpewhbdWevDyGmGnRVf96d67HBSb
o9RZmXzgBu9mITVgBEJIAxnrR1UYZfZ/Xl5GUR+di9II25+WL3dAbd2Yyykf
UHY/+zuHNUHO9lvXgku2xhUn4mPjaK2dq4Inkz3kT7PqwtF1V3ojMIuj3Q12
l3dOOFbw5oATM2PJkese5YKL2v61A9RUrBUjP/dMPuU4n7Cp9QSX+eDqiFTM
6zH5Ao9AHCvlw25IwPTGMOGT6yHOvuRc8wHZiSozf/ps2FfCbMCy5x2zIs8S
DXDqT0gmJiJiY/AUDitBMjqPHY/PTs7TT/ouqQ7aLLVP0t6H/5r3m63runPw
CMi4ZNeIyNWA6iVOj1pM3GkLViqO4pyer0rS3tD/2NVUPZNi4wIabgElxLr9
nQK9HIFs1RZTt7nc3syXlsXu+HhiYdRrtKEQD8X5u6qIKUYHRD9U4eyq4K3a
eAiUmlb28RHr718twn4Blz19W0nGLkRPjYQWF76JyU1/6+JfPHCRXbnbfBBu
79v5DXngroe7v8i7M1oidAe1OqeEfqGVwnjTAcXdlh9oooZnpJGbvKEeQZvC
gi7ZhVAdNMbfXRm5CzRQTIgMhQD1cfRoC6rUVwJ27ODuRISIEWPTUv8xuIrk
UHvNErYwERztcK/6eJul5qjBV835BUHz/GfsOLVQx3FeSyj+/fTJsciOVoRN
FxGuFZ7ARzPP+cjAVa1Cw+qwLHwPVsu37mZ89gq6eVoeJQcLROBKVKNLhO9Q
+OIPnHf+CZQJIXYfVxX7mBrTv5ZDSjFug3gQtifx3G4o7QjIytVtOjbofgYW
guWrvSLNDThFe7wntkevTHQcb6k0g4DReoIXmbcBHukr5ytli4P+mSC36yFc
dP+k6K2q/sSNhBA3GxKRcgDwA7EunR+jW32WWMnWEC3pgm/GPZb6g6nTRfmb
s3BuT2qYdRiVxFROD0RZL9HfIAOO3VzOPlNtETvPLCCyKrI61Fh1mAJ3mrYd
YiP36dHYHfGl2oTikmIVPKZ2vh9sGdnyQMaKWJ+hBK4HfC+MMxZVOnR7wxrL
IHRFoJP9879zcK1THFFxiq/zgHpqu9X4Nm4mmL6O61Xef+YFDSy2KfHpPpI7
G156ajjwVTKpYj2CouJDRsXIG0k+oiC/3oOQkJasR/Sow/TzXOMHBUnufFYN
0l/nKfgjqQMFM5qwbhTmRGpzsFXO89ZrYb5D19jVm3tALjq8ew2BjEmG3+Px
wJBO+mOtibAjgjORdcDNZRavmkiiLthC66GRMBnUEzcRni9yEki9qlH5wR4q
OtiepFKLxlC6zBpRBigs1f3PUCIzwj09fiI0RHvLXTaderS/RwR03YUjGeNJ
zB8512soI9JE1tT+sxa//3JdMGwdLJ/Bl99GwaP/zn9iQZ7YglJC3vgMnvx8
esRvJ6slBj7f2htH6K/9xye02vOYvdusRcRPMrqe/9H4H1ZJsfLJudsAewq8
MgUDOV2pidmMw9/HOg0ym70xLO/MnAWf1zWFYicQYZtDze3uMUu8o/xiImnq
L7NUGpLRu1ohNSTgN4fTYYgCN+RoabWjRuJGz1oKYNAwb87m+JaeabMGNYA1
rB2uQqAbM4Sfa6I9BtG9F36awYh2okCIo7OsiYqDZWIMeYIlCVpo5Y1mBbBn
gF2iIdHQKwzGqbfNIEEyqpK6YIw+cpWNGHXbUDyzpIiJTagv+XQU/9owZRQV
wKk5/RPCOTrJV1levsOr49f0Pe/Bj2iIG4tUuzUIN1C7wN+ZA7NVfQoCpiFB
Gcq3QoC7SxlNk78AUQQi7wWVNAa3IMMLxln8pAecOlT0llHhAZINst/NVlke
kjpND00PH/IzDIgNiGIRWz+BuKUklshL0LE9+LiUo5yu2WOQEKwTst3MWJXw
rVAFQTuSnM6QjFQus06AeHanjPBeBaGRGBpPh1q6f1BLGU1p0vTp5Vx/cdXM
BYFSQTe96HGOZQUNDgPAsDdK1KVpBNHNaTA3Rn1SULQE7ym3CbuMP+nornNc
5IFOhX6xHcjt3nAOfD1IDqfSRfolk6mL0HADcN2TFVgzNSuCmJmN2iwSXccS
z1VwPW38QkeiQN7CLxY3Tkb7OuplSWksezG+fVqA0ZdqWHjld/cSpAevhRah
g5PpXC45YptkhcZ5eb3adODyssbsRF9kivt5DEpe1sNbLKWsy1o/vYf5Q2aW
+bhRMye+q97iTiSYAy797FDFYcPhrMwzCxQwUig2nV9QZoDj3WiNVATYqd02
2E+P5J9qR4b7WENGVfjVw3YTkJE4N7Nie19IsDoSWGCrxXz3eoKLy7ayrAH6
FJtySIpxmFRgYBeQWxhJjg66UXF4Y7Yn18ZOsy1VdUW6yVwv50Q/YqT8Yky2
1DUSfPvzzCZxAElZXrcrDZTGT0G0BLj5aC2KMA5KbLrZJouqRsgvV3BhomTM
5ZT4sH4XfBiJcgskrh+YB0J5AQpkwoCKnR5/bRkfl8E1tE9qBvlNmc/nuQYy
xXLiZLak++ESM6mfiLIrhko6PKHQQTcwMZRImkHgNZ1Fvl6XH3qATiV0h8WW
pMq48qSUlKdS1qT5z+d6VHV88dXlTIXbBcQUVaigNd0I+ReY5b+BvEXhoS7D
m8Lg3EH65U9pAuoNJrlxdULfX+jADKqmmH5kEhicezBq1OGTzk6x0obKb3tg
zEpjQi7J1d9T9GTj2LXWBfTmTNq8owk+qArTuOqztTULR3yGzem4dACRRyKO
YK5vbwp1fAPbbwkY9IQ/U3heIcM2na1bYhaNeTZ8pJ5MYunvH9bwpVHn01W7
tAy4t5u9WaGFAnvztnlKhqs4lpuP/QDexMYRu5H5NXjNwmdT3G2qc4low+ZO
p+GxRHdx7vPNLZ2Y8zvkl2yIdlmdl6NOqjqQHtbNlHaMt/5ytwlbZFLP1qCJ
uUwQqspVt9VT7WANRRBCjCftTXEcpeNzuF+ayjRxs2zmWvVT2gL4nkZpGaj/
ztOnOqYWcY26UEEKgG5muIv8d8Li/KVD/lJUSC50iuv6OP8GsiqvfzYp8/rD
o4ygecaZcLgu1/Boto6n0iErHAojmeb5VocNN9+dspplte2U/cQWx+/b2Th3
FHVIv5EDuUp0K198QwQmd+liMf/p29bIkeOnVS0rpApIwTETzsU1P1q8PKDK
mnsvrEIswCYxBtwMXmDAl5YZ+OpN4wPYCWCdyd5jxsCZTAeEaHH75dieGhcb
HnfjS6/psmvSo7e3DSAxlMqPaRFK8Z8mCdqGuYX1NuAo+91xF25qk8pnZKso
URprTcCnhOlXhDYwjWj+q9M7h5eZPs8QmjRrDpA8eeNmoMXm38vB4rY/n+tn
igmnt0tbOWNNc2vXKlv5zf4TMDn4AkY3hrNgSxDWRpu5at8gG+EYhHlgQNI1
ao6eKqu+aWYkHeL2WUpcBuyeRqlVSQGYXiq4xiDSYjsqWPzHKLLk+xnEdsEE
TnNEbpqptRPh/6vSbxUTm4WEAXggOnPg7DCVaeYRr8jAAA5aQHR9RvEjwqLk
PFZYT3Eu2UjDoggw+ZNMPP8u/uKImSNzAp8hMuqKo0wKfQzz4HSxIIltaP0p
ciJHkmQShEQJdExwF9FJXkOGbTpJuvaPdHu2ACw7BCRKh+d2MiZ5FYgIl8d9
L+ykajsWZf294tJwDCZz/mimOTdh9JkkV2vQbG9zMlwEUuZL4KV+FiCN6l74
qaH5WSlS14hsp4Yo/kxh40gb5Ch14ERxRv1ngFzlIcRxa4PCmy5iTjjGZST9
1DCoMtOqp+bTgWNPH0l2QFqhr5bIcYTVbvEeyo9OgTQL8DLsfR/HYdv51SHf
fbxTu44spJmwKjfQ7t03tMCTUbXU7VkgBjbnvCNYU1Aja4XbYRBCCW+tNTql
Dkpqn60nquE7pb8Xp0UjwWET5sOleKHjqkR4Ct2QAgogqYQXs28GP3geMjYP
h9s/hEPVH1xeqUD/psfVjrDYE8QGxSIfJm94wptMEYcxca1EEyvFpzHEF2Gn
L5v/UmvRdBh0XEgH3gWfwa3kAo/VMUxxXAHHQ090sO+ZgZsrq12kCAJ2EMSF
MULA1kJ/bauqJgUCkerQWCaPTF9HtQzk96obXssv7qUcW5TGUSnlmXlZkG7P
ox6E1k1AILupbNrzU3iyFMuPb2/ShtmcybF1sQSxb8sIglKLTG4PMQD6I5KE
Xed+1RSnLm9U0XCPJ4QlHEFCyoTBWwuOzFBlAciMIPAOVouX1lxtO0gqSeep
M8mcGRN8PMz9nZNi/C9OtrR+setudGD+XoTwatZTlCJS5ds+Pz1tGdkX5x7Z
Xm7CFWTlCIXpqCMop77Q6BkkaussEsDzKD//TtNWqUUu04Sc8ZsFAmFnMJzx
CFKXWx7RnBaMMqPmtApsBBvAv5KaUFJD6vnsSBgUx/B0Nhplld48TV3fBsm+
M7Xp0VMoRWiv2iHYE4efqgJO0fwd/b7Xw6gdwU8GWh3WBouvTVaFUVjtGeXh
lfSQUkkbj7G8uBoo0k3YQlnLiTWhXG/PR0zA8XX1MDnLgC5nI7/Ojj3qDyxC
2iM37h4zb6KoolH3K4FKtXsDOWCWJQBmYkjeKStjLvB2Lwk1Xm67KgifOIhc
HTwxy8hZUv1HTIq+W8ipBlE9FMDvjpulEEt9e7Q9EnB6HjcBLQ+IZ1Q8D+/T
xGh6xTHjjkHQyIItjNbVVMSC3iOlRxMkwy9NZOEbb0xq/ydLmZiPzBLpgWJ3
XIqmyxaQQJRC22qvYscoh2fvuiJKt26pIL+NiM+gHplIUj2zvgbbomn0Ikan
wDOm0Uun5BD3i2XmFRU6Y769sMUF+ce7Xx7BdgZg4VCt0iqwWFWCVhDYuEqT
xWXfqos8nlK3SvCapMVaZoUVXz7afxk5O7vDLoyAsvTmOdfUFZA5BKUTUIa0
IljYO8Dl7PFy1OrthsdXR782wv1nkQb909Gqjclz/oXcJiMEi0IriMN05DQl
xus27FwjW7Xqstw7PSmf8R3ZqATx/tf8R4TNHepszIYuk4qBKlVGYWCRQjLH
YYUyza1WHhwYPRT1a5ZC8IT6JE6lbSJ5NQ8ENcjw0qQhGLz5bpwZ6BspkmMo
Jmbo2haQydIrwYloFS+FlMAEf+RvmYWDBMQEXB5dI/9ifsJD0VuWkzen7dVs
08SuwNZX7zGZEN6/QurF4tzA1/dJ3cldILEpJitRsJlRJqepGOBctD/1Ygz5
zPLyxvQqvLFMhHe1/ZJYpnL/PlqUWcNADhk6d75/3I38xFnKQ2QJuBPcoAnb
KgbthT1inVh+hiT+dc9LWjnGwmPhvrk86hxDoFdCSZj/+yoN0o9popY8wFBn
0wci51VDGYYKBCjY/NRTXLrPPoF5UiL6s1OEr+pqLLmeNjmYsTnyfS3LCBbf
o++sNjkNIkLpBiTyCgLQsVPBMQpP9SekCfCiq83ZR55I3QcngfaQNxS+dphG
TFq2agWXLkTVe06AMrPiTl8l9umiHd6TWlKBMEB6Q9T6pV+r5uiPnW0Dz1Eq
gW1tth4bFBeHq+E3wHtz7c3equ7hKbF4UzhhwlcTzePjqt+ehNAgDgf00JPK
EshtOoyuxY5DRkYmH3sIQl8lfelB+WIHjdvJXX8p2ZY6eLxHUUEfaKkIBXY6
FZDq0YAbqdmFOmb+yQM/byU/kLBjl6hFsCPm3x6FfGp66VZVQP7tlvpWbnjf
pTUnr/wr/6y1WEsyw476JPhnsTEpjvj07U6/SE/K0TVKH6wrfL9MFUXcKDVh
z/h8Z7KaIFRq9M/UX3UKFQz/L1o4cnj46hvQNurhN2LToyPPPRT/o6UWnVnd
QoVfiEYZ6Mv0pShxkf5or2750QXkZNoRzHDIoRdLEvJz9Duq78Lu++4mYqxV
T1zZLYOrFJHhbOX9ozRlJoDUkkRqckTuf37DdGfPfXRhFQKc3Pv31qWww3Os
w6WFku0HzQ/bgf5FZnzCsdkX8/OyWPuTi/qo4zP2I08SalziZgKUT9b0I5mV
1UZ0k7oR/6ePE40J5CQPp22+1zei7QdOlZp+gcOlSwpi94xwgzB86vthwVZY
X2N+rZi3Lv+E8ku6LUDNpq+s7gKzOJa0DZCYI77QrSGcCjuQ1ABr9cYeX90h
EBtEtrnuA09+8Ol+eL5hYyZ8RVTpCZnoxEcGci/84Ia0Arj5cqvhgmrNEHxW
BAjj04Y1r5rortMquJ0RzZSQiJLcuUm/+35P/lVE89SPT1z2KrshgzpElWnu
pcUIX8BrsOxQQI3Qx6hzNeplkxOFTi2VM+fCZ2F0I5VCd6ftgHPMal1UtjrE
e+Hh5a5zEJmXNV875k9q6yGO7osrnKhfx5mTiU1jZlVj1VF5Qf0cBuMRCK67
+iLwTbfh/GoOFjoHV0wXqjsQs2/lDSUqH9+CJ96sp7ioM+zYpVWFbDkdr1HP
2ILadiDD5hW2h6DSn9ekgCg=

`pragma protect end_protected
