// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
xfVvmJ+qJA08IcG8qb72IVxwBcqJHu5zjVuDdZPUvHB8GONyqQntl45gMNKK
c1ynDnuyvVKDIOR27BrbakgTn6KTkb7Hbd/57JqBkVvVuewZEH7y/lqFfzFm
nHJpYc4lULr8Ce5ZIDxAzvgwRVrNiXjIwxMNg77nlE9m6Vb5HYQf07jPLcLO
Kouz6cIM3B1rnpfYlcoLIFBHSLpYOMg9bbzwH7vP9l2P6NIuNns8wVfRdDiU
QbADiXjP0daQqWOHLr5l7JgP1hpH7c7tZXpQrtAv8ov+QqEZ/+VCYAgudBcL
RP90hsyZpXWRhrZTIZQErdsMGTvOp5+/bKJq1yQMKg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mncZdlO6LedbM207UN3lOXBfFHs0/JxvxWSEYll3MNknHgQRaZ0NB9skE2ZC
h0p2HCzTq8n+bMVD296SGD/Mdt4B8zLzOAhNnOvZT2TRvi6cRLgN8gEJIn3d
mOu/kL8zWxfbsqx5KYKipUp+Wl054zbBt/56rVwbCPyDUIk1GcIiKB8clAUw
0vAACo1sCJyI7iq/0PKr1bom8iT2dAc37KimnbLpy1UERumdZ7y68x+dOjM0
s7rJmHcpZgZ4AVC6G5i3CpA5T3wROulSckNQyuQkYZ9oY2/rXWy9p0vcP6E1
CxAY0e+s6UM5wKvccjTkaISgRyrQmf7ZEB/GR2tHhg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KDN/2el2UFw3KP2oQwdNKSsD+WDzqVu/rW2Lq/NDoymjFJFFDywAamTHyFl+
bqtGgQ2laN1/6pBeOaWrFbLv4L3F5dDoToDeWulUc6vYqU+k06jiRpb2wwap
ZZU//AyabNONwq1gz/nMJe4E1VcOX4lZb7nqJ3/j1CPAiVjGoxbX/R7O326R
sQ5LttsF9jt3Y2kHtEMjzJujruhSmxDdiMGOSYAoDPYSuvJncr6SWXPg6en1
TbM98EOS6sH8DV2k7SeMdAVrNX9giKQM8jZVgbGYg1WUAWbBKmDbUB64+Om8
gIIRj3ATF1eb2g378bm8TcMp9ytq50I1SoXARLjUXQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
WhbOLGpLsUuNn4r1xOc0OCA0Afy/Xw7DHy2SV0g7ZZIh0c6+wD9fLrUbJ1xE
F+R/5OcTEqv7WKllkXwpNUI+KX0KCMCuMp9V+kACc0RgxD+SVyHWLMWDC08I
yhOcLcm+dm/C8PLY0VrS5I1QZHVwKh2BW6KoxaDDDYRMNnMoYLo=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
PrwItTpI5UKieNS7jsILJFhJv5M5ke0JsM9xO6odGfpP7t+C/iCkpKrAKsql
/f1dioAHOkdKzQh8zRgRXJfs1otH22gOd0CTZuWkVUMETEg+zv9EwWyEz/2f
CepNEjvpCkpVSi74W0FZP1RQt7Qg4ecSzllZrByBjK1WuRarFLOZnOfZky+E
q63bZfdbexEVB18IXWk0n+0Ky+gM664VndyyXBAPd37QNA1rOKyiuIyMB35S
UqQTJzFjEv6OHvB3SOd1eLRSj8vC1zLNitYKcLcXBXWILWqP8QvxZYDVrYNo
GASwO4e/olz5Ov0c7ESkRlQS73rf4GVlqVbR7nAhZ5UqJxndXnkNGNKw3eb4
B5gLGl9zl/ntBMITH6KiHTpc2ItnWx8aHtsV4nu8hMeeHbixiMP1WyJBLYGp
yzYF1TsAG4B7x0kYu8pf/PVo2Dz1XvjadT9MoYpZagD6ZpcKA320DVxbSfBT
R/s/O3vRJW9VR5ZhPwgZlcLsAmSnRKLR


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
k0K/SEcHvpwptXAGY3vUSzAKPCy2133zv8mDi3oVdjvWHLlJ5iq+qnwe8Tm0
I4RQyBYdRgWfOPL6mw6SyFZjaR/aZ+54DYrf3lZJ/j5UCpglpQlMUFEN4XeZ
K6s4aYYtxvpqwtTDPBxxqBRLXQwZmADVNDjExx7arJGbk9HYoBo=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
lzN8Z9nBSujzHTgIpLhgukfp7vJUZ6TkBYl0DD/LMmL6cRAu+VkSLKAL5Q5T
3FHFZH5WSvA6ghMoZ8J8tI22BMKohJ+1ld/x4JHLq4xeTid3T0L4qRryj0ud
pcYt5qHhgOGd8TzW0pCwOcQIIfb5LesyUqK7OF+2jvkh9KY6te4=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 23536)
`pragma protect data_block
0500vqRGCtlzr2Sr+Lfo8gxm4P+Zy3syo1kPXEACjAq8n8DvJXoo1ODACWD0
BnzEDw09zkrphaNTL9cwX+PPaFQxVmfjSDuknoPsEmvWJ8Mb9Jpbv7af2myz
eb/61vtZts7vh4t/Y5nDQoobMQCAg09x9rjomVNPTU5RttV4rt5q9tV3r98Z
f3PtLpVu5vE47kE6bJ6YFhgslSQmZfaBeyHoPFRbZ35WDNHJ8qWcVTMIQytZ
Uk5ZPQ84WseQmV9cIuY6MwhT8KUAVa6zsKFKYKv4dRZ81UODWe25/7X/6dnc
G5DlFisEWWNOA1XZiX1arf42obns6rf1o+rDxGuVc4KD+PRpyBAvuoZxKTh3
iCA2yR1GhccFfbJ9KdeONO0jcmLc1DDI0f+Ll4RyRrHqbXOE8WYWMT4ljvQI
gZ8bk+ImBI5tPUNBwnq5fT7XyRwPzQcC2fcaObyx/pqfO7cbwncbA29Js/+1
OgY+FALvVwwgR0RiG8L0gwmoPz5YDJLSW0t/0E8hYkqDb8duxsH5Kio4hkJK
gwItkIpHHPLKUEw3NEeX7AOEmbmc4eYntJdCj4HfJSKR5Ht6djYA76K37meH
X2G+LrRMJfGBz7vEEx4KWQ9ZK+p7o8JMubpsCRW5hStNkvsqyrwbXyGDIEXD
s1mpajr3z7dUt1uCvQBPZWILqC6Hi0f61vxfqpk3AGO+mTSjLGew0kJRHwZ0
6sBl6m5ehnV4blAAVq3qI2O9n8vFjntrRhFIo3ioN2oXQQEeOMTIqC+6Qn0L
SgMWFJraFvgzdLxlbA+EUig7rag6OStvu33REnVQCZh35KutvKlQE3KwGPYY
StETMWsxTOqCC+0rqdhVPpmX4BYGGBhganAnLanemBI7WL2ud5gi4aFaj29Q
pwsjzgkHeN94LpI323wplWVAGitNmd+ikSwHfFBemRGhLK+yxDSJ1sti7djl
y2+yd4ZevcAROEC3ZXV8TcvonTzh5qJrVo3fBUb63FHf7YcLAlI1BKARtRkV
bRNz1u29+c+D2X+4pndYUoFhAePWHMy6HR8M0zZMDhQ1Er71PjhqltPXkZ7D
wIT24gCTSgmT3hYgNbqKRILRuRufP2QawppE2E82eMzEF3dJwdIE3pF3iO/d
zOeE5uC0u+ZeFAZgefxw+vR7DrFT51wvGrS6S1VuUhEvBEEq+4CiF10I1rbS
5QMPcgemSKEIEf+5Zn9PYITTc6immGM18lCllVtKEf7kUJLC3L/M4JceBtvW
5p9oIs96YN3YFmO/zY4VI3j4k3dgFMVIuS5ITPkE667sKcJQ4mgi0eVzY5B3
yk4Q2KwQaNe9qNmpnkrOXfFLkyvBt8JvfOustw5XaPBcbbRsmCec7lpTVNM9
kivDrHz86NFcQL70CJYAHFG+srpLTesiu6KAfqZ4iczWySOaEedd+SrJPygY
B1+tAPNgBCTJ9QgDgmdyqDVwcD++9+vZOyy6wGhGDcBbij+VyNNxIxpQE7S6
O/Q4XJoIczS12bmUKm+MlwbrBIOgBRu/dH3COyHs3YPFH0jB+qKc1Tv0lHPk
lPBj6Rtrn/Fhzzg46t+WUy9vnowV9x4aPe+aWeAUTXSYdny63Bj4sh1Hamj8
+jCI7iUSO1/6IH8XaO5xMcyUVUbmIGai2Zp+omc2UDWPsgXuC8g41JKW/4TL
tjPSNvL3t9deC8NvymXW8Qk1zcpqqOuPevPGXsfwntBk/MJpTgTuu1fE59L2
IhYxW3PLCunwg/fP8H+FWhwJHV/HXjOR8XfMTevUZBZJVgvSgZm+T9KAA9eY
5i6lp82AhDJGHIFZKiMAesHN6dzlKFmmYr/LD4dcJs8iyIQJ6Fh2bVqhIIkt
Bh7N09MkpIRBVRl07bl0cV2KmfkswmatrglI2Lld+u3PU5EIEsYU+796Zr+j
px/lBpNbjrdpSIUFdvQ9XmCwN+HYtUgJgHwUyqJUnUx6nzup0s3qyMb2YECQ
mEADNPUQyA2j4dTsfEzP6eeNxAtUWus0KCCeoQ2Y51ENzhCNwzlVKgOtUurj
FPqyKE35iKCXAW9TJ1ldvjSeuSZWhTxxzNbbRvN4kUkB+FDniAVd7Nl9jN7T
p/sMc84u8jmirOEsHUKInKdADzb2w6zgH6jPYE27V60t/yUTA77UOQsSnydq
zHTscctUd7MX4IZZLiyjfw+hOiBvxNtSMllNkB3DkjsttYQzuFcKRhp9b9wu
JpMoS3lyMVfiWjlD83V99fVWHhjSDEeTQAFTw2vjl3I0tp6mz8BBkejJO+hP
2XTWyBpq+PBJUkXDOgEpBi6/pmHqqWVEtY1sI24v0Vd9u2yTmIt0QdaQ3XVO
8DW0UOYZl755M/SJB/hAVT9q/v0B3i6c6dFGW14hMulXBRIRZQV3LqMjFTkT
ERJiW4PbEyrcb8EzEj+xGJi/OZ+JeUdKaggrVDvivof0TTg1AixL4FoTeUUc
o7gvJufJFZJVznfyOFyu/uF1jDAV10bUkf97lcOMaLd9UXtttbxsYJZ+NiVg
eaXJS3uoU072dLbXMwnY4hKMW+49EYVyo9O842hA0fFXsc9BMQnLHuA9D9L2
0+YFRCve3r9Nag8B3lhjpsPCPPFAkG5tLjrxbREwrusVq3AG2DkvR+RRisGy
CNh9mDfnv2I/EUe2LPunoz/E7YCzSKBqFj20FIapGKm2sVvwVPgFERSgEldg
dC6HhnT9zjeL33VTgR041ys467qR27TmoIke7wYDDVmoP5X6RQt+OckDLILd
0pCi1fJ0FOyHiBo9XxYAi6wZZpo9ebp3UZLaK0NQqdthZ1NFDB83axhHQqx7
J4d39TntfRXMO7RSbcLOyGBY6yCFVXHZEwkyz5iO5sf8OxgIUwyiSc5BSjXZ
XIYzT5VZ3yIxjnjLnpW1LWIooZPzzY+lLQTtWHz+1Av+fkMRxPUsJ3oXrI5q
3Mkrugj79q7zT4DhIgkcxKmXz1TcqVAHJYiAkTHqxMn9mI6BGgaqnWsg81vY
sb8YZPUJNYNkZhQf4mDcBOgvezss5uYfP5AvDFmPJHmIme0BVJr4t+VPK8uU
iGBcM41iPonEGnFNSXdvCiRAr77OqyLfkfodeQ0WzRHrDnrkx7NJ3xbN6Pqb
+sc8RZU0OYMMmXBDjhcvcSPVpqsbQcia4vWtjwkw1ggpLCpXhbgjQEQObeYh
L6a8ogXURu/sf27FOERj7VftStLVWqUOENeTqPGmGDeK/ciEbLFHxXGGqShi
/X4+mYfB5pu/pjWvRdX76iWOK/7bGXJ79EoEiFIQHmvt3/h9h1fPQXDrdhuJ
lPrsOO0NWHiczxGvhqhv6bJI1PdI8wapENteegiMoacbjHP/W2ewlfi5dqvJ
dYkJZZN6epw3nHZ8UWUobVTVP7D44CIgfw7jJrK8vIZBDyuzcFhqYsCl9Qz/
/5xESbOJHnfAcDCatIYRC3JXtcZ5AGAOL929nh9pdUmWB+6kc/LBcjT6+TGD
6Mam9IdIJnQw0Mg09FN556Ha9+2U3M1x/C6+EDur45yNlyFgNWstrPy2AK2i
zeRYnj9CloXFLLk9esVDkrvdbdc3VvFMYxpSDYnJnveqm3ZC4bNPxywmooXo
WPPExo5m9FcVmU6KE4/c6XSmxvf/HsFq6ImuzU2fwVDirbVorgasEFmzjSWA
amA2c0/xypJQzcNlOe0Vgbpmg5USkYUCV8dhmF+BeXEr15zGVRhRCPyMK9Kz
bI8u6b6Ft1tk/IPerIYhH6GuZlPK9wD5ncLgJxACng68+vj6Uj4E3LZuR+S+
Zb4boTtf7Gi0N855WoaY7HBnp1zA4b94nkIbiJBWlaavsW9Ia/M44dbp6NKs
83XMo8KXw10EaOp0iJrHfCD7xbPxsb/OewiPYfS/pNWxUbe0heIr16TPEggB
YeeQHhvsxAbJsCAyoSZyR6q6shO/idXOuerCmIa0A4jRYHFcakoCr4+8UO+D
1/tkAO39J2I7qA3bAVwIY4zZXB1Cflg/l4GDy6fgzgPac/vlM3JMkFBe/orf
UQwBfj/26icNeEwXaq9/0rkqm4jUvqnYCA/rBPvODhymV7MfT4D6QQw+uMO8
UpnCLplw2ta24oV08tMqass0j27BfuPahjv9A65cxrICMejyUPSO4bb+4F7U
zl6cYMsYz2q2RpN3uWDddH3w18i8vkwOzXRGHrVtkB2xk8zqA6Ax0/4AHipG
qDfbneJqkNt5zn13660M3O83gKGh21p8EgjH/Zt+qhSqZWDWvzcqDKzeoGEp
Pro9/z8kMTzCnll5ap/JrSbVRBXcyqAiqG/nOK0Ize9sKt2HXswYz9HKk1nq
XmHIlnkSpyynoQ85skspnxK60vit+q01n3IlYH2+xaWrO/xVySopjToe6cUM
7agmresknucglCYt/IbejqhiEGDDFptGi8KTNQs2w7VZ1q06LY8fbZ7sOpMv
NQvg5hQlmrAqcNPmHHtjH3uOVqEEGJlpSrO8nGTmykuj9HtT46y69Cs+L/bD
KYLaMzxA5LG8hJFIfIMz0uiIhjahdIq18xWi/JLBbNPnwUVcsa9ty6SF+m3i
o1CfhjkEaaO1icLfPyVV4s7GxyCqDxaoP3xJQezzA++5IyoEvVqbUfeE64Rc
WVQzH6fXhKJ2p0RenNOa2buOxUU20eAZXCgELPxQszT9fsMg3YjMSU4zYyXS
zrd0+OKLpGVrAY84KYYLz4i4T2SURo31xjf4jZJy7DwrEm3PEQOQ5h+arvg5
OpSWa/58vxM76Ae17Rr2SBEFXdHv/H3vu2h+ibtMf5SgCQwshFn1Xbd7nmU0
v+2k38mRcoRK/yEASL30q7cRkhQ0h+XzDMjD60RhjnVyOMJvugCQq/9a5yaa
P5p/sj2lwKuXOhocBJF7nhwCA/XOAv54cRMD/VgxudwLLbkITMc/XzbwmgGy
r6uAoLDp2WujDNkvL8VfTyVRXmkdD0XkUMMAklQtbVZ31AwpPj9kOFWBfzGY
yeuKHI0RL0zSun3XZGeKGWpiMQSw6cd3l4IVXOjid/sHHtA56pbeUVMw+uar
86YT8ka3Jp2ftTq/XqRmvP4kkJ/5dXMPCrRXv/EYby7yMd/Jq1DXmMQASVoh
edQnKa0Ezik/A5e9DKil9gv2cgSUJsmlxrp8Cj6/W7HF0MKKnFPSNkU9t7Op
xEHePDT7Vuwam4l/vXXkAh5xdGFNQLFbD2KoUXk/ebkSZQCiVq3JN4n2wENc
oxeCKwu18FDYA2rsmeAUW0xiDuNvA5B/NSiQxR21bXZMjwrflvDhfQe5oGmj
HQW5tIbjjlWUFiJw7ZJ6gLkXAFC+w4a5KQcKDe0PS2fvNFUdAM3wX4DarxWn
CopjOBgy+nyNnge/+ymo1es1kd7dr3sPLvEQhYWsbv42FJcYFeEt6VSl9ChN
wYDRgTteGBVOiqXBqao7QvH7FrJE4G5bA8ovHYjcYP7VJr7EBqB5TJeg/dxC
ONDAB78r2T10+SE9zmVDuTpXv0seVZbDQPB//0rW1mXu591G7PgvS2FIObAM
1VAchEO31sHFulGPbShU5mPCC5JG+nI5IP5pGcOk7Oin9mdtpuebKDaTq6D2
hhPrfsEwivD/4th6RsehSpgCyEXrvzCYyHaEvjmJOpAoKnhO6GrTd+qNZVSH
+0cXeNrYqmRggxQ40UmQJhvKu8EdJoeki/1+E9R2NOomuzwGrC07SCL8zLxt
h7ITjq4tJA1sYOcSnEJ7RRwmWAzP/j8ls7n5dopTgGzSfHCpKQdfdxD92WGX
f9gwcgDP5e17MXWx5NAXhfC5TjcXKc3b5Kx7o5uf4+4W/go/oQ8gSFJLxYJf
2EKEoIAIrr7PL/TC63YBFEt0qMU3u/78pXn55oM/tocliv0Y+/cxIZPh00r7
CIukFELY9m9IxZA21prKQa/SGHQOzTUA+hE5nLGL5GgW73ZK4FGC/Nw/c1vc
bILl/WTNqg7f///EJ+v+dtPuK8ZKE8GmozsgHGa8Nc+MLtXMIZl+l7GTJy4v
5xUmuc/HOlkS7cnKTkdv38jtBqYvM6BfCqQGDG8AqS+eeER9IyUp4FjhtQs9
cc10QiOes8QvNtHlV8HgKu02Vehi/r4naQsPKbaT9EdVVU55edPSjHdllnIF
ArqGgYlpTkZB0hqzIDx0/ptUPb1UmUzCjTg6qeyHGKQ+x0B91OG/++CpxxQ/
UyoXfnD4SwdV+TGJHpJkbfE4j9AGy3rTsyqMzimAlSNtM35yUAQXfKRC7o8M
7Or4w++zbEm5vuZ90bry/g6aSo2koetIkzF3efqM5/+9tGw6kVagpzJ3cMwq
5MPl82SMy2IpI1H2lOYVWxWtuAoXQUk5LvPw7ft+Pjul5z3uhwXsP+A3cVy1
CWP6ohvecjR07XLaOQWA29t175yQmcqQrmbZmYPHAcxMLs/3/t1hjFxJN0XA
mC7bUEOoqSLfy3imTLcY7Ca4TsyxPzRx6GfsgFs0upZDoIN6PKTAKyDiCzox
zK6vjhXOY5GYAgCz2J8oXkX1oN4A9ImXCgR/EPZ38k26J+T/cE5dLFtepkYD
gJ8mJrvRh8yUGrZRrFTh6i04rSzVd8Jmi6HeSho2sHKIiosTfM6zN1gnD2Fr
juVw61t1kPVpM3T8Utr+S7gz5fvwwhrMH0DMWveQ3zLkNZ4vrGpgVubFZrC/
gGdInWsL7+aogvauKrG3QyKVpSD0FYO1J7kW6if2wcKqYhNN52ld/u/BJ2fZ
P0O4HltbIG7L0m3wdnGJ66/dU1LsWsJJZfECNLgddWIZBAZPa38v3fJfMJ4n
+7SBSxA0eyVaRla2YA88fqBCp2Gxs73bOXzUPgo991N8//FUz5COgLgcNT1c
JfBdxVft6aUH4sBci6UVxjK8MLNKpUsNZLaS/2rGvL+TS8/iJVCaI8MuBENO
CADGWdRWrs6AtjYB0CzO3NmBAkEXhAu2JL66CkoliISdq0BEQFNo610eZnZ3
zYyot34sPdngQEEDQBgd/7rQTw3/XYIJ0hfhCOqUV6/qvlTgOvKZyD9EQhZn
9EirocrJ9oqZ9rvVDvz9AbpaeZrbWqwBbngCYEzzf+Kvl62uIrLR/aLybf96
s3K5oxQCVRHMREHGCgNU6XT4P+sCBJenMJ5ILlSWZJQRNvZHcq4Ve7UG4UMu
TyhhlwLOX4Rrb6QBkolwy8joHxaax542IrzXpV11Vt3RkN6IQL7vl3REb7+f
K/BUbgexQHW4fo3RAav1p6jhOTfoC9TRwR3iC5SjhB2xod2mU3/TrfFAB6u4
+sSlXM/hq5G5g4U6VHVa9bg4NbRGertseuo774yAgAJ60fqJvGYrls7YpfLM
fUi3F+PYLVumKWNP2MIio1paHEB5hIoMFwaLNsG///bbomzTk3DkEOQyumz3
ggx+RqxTlndEdQEqEJp+17rchAuGfHTsK2CUs109uNYBnCRK+Feka9ctVaL1
+2XIf1LEAwzfVOW/R1XdVksKAGi9TeQqweRrVvvT7uwhZlbqA4Ku140o+Aju
v4thd0M95NsjYHXmxcZUL3ohb9xeNdOjNZuG1WnODGRxxNFcfmgl7ZwMr+Md
3piR5mjAvCz9qBwym5uXtG4kMVBvtKlq0kDFVBaJdGxyfw9Zdwl5hFRMCIkL
SsV+CMxVn2Tuij/YHRuxmS7g3usaoaucjivh1aEM+5rU4UanNP3E98uDNqTt
thxJWbgtY9KBH3csIwtyjpv/YxLzzzWRVSYxGFgXQKO3kBieub8L6ci5Hw5B
dHC+SUSJqfN1Cl9ozq+Le7wo7EpNZ3YlKIo94rC3LkPe8fu6WMRncAVEv+1g
YMv6fkprH9oo8/MZkr3G55lFJdRM33HNIPWCCn7kmIOUU8YKv8lLh4gLRCkZ
LpFV7GKLizTVxmLUsx0dkg8EW5jhg8UfzfJMGbA7nAM+DN2eca//Rpw6RFyH
F2jbiecSm5oC+QiYXMhZWgZJCGcAiS3bL1/UKlpuieqHhsTEW5MMYXawdc2T
LOc3BgAGfSZj0EDpumOWjmFqnVtk3fTrcNBlzFAR5Ypye85j3WgAwLAG+q/l
EtLNDiK6DTnKOvP7/RcbQA/oYJSLmzAH69qX3OpYGkbISQPrABBuMVco+TCk
ISCxFvFvDa30m3oYtLntgC3RQoSR56Pwld31meAVNCUlP6JK82ebgTlSOtRz
NFHN5whHqkm96OYjH7oZwPnxa1SY7hW+uQ5D4tEkJk09I+ljA0+lPE/VAqT8
sv36BDmhwLw9LKLdD1JGz19TvLSY6uPk6LmwPdi3yf5pVXrVz97x1PaBAIP7
fl+2pl3ZMgT9HB5EkrqY+SoZPepvx6KAgJi/wPCreO80QL1zM7x3V+m9DRtp
nL/HFx7aUmAg9R6z/1u1xZm5ACsCsSoUnpuWTCIqNw+ooVSELTsb+wMS2HK5
49cjkrNtWn9DjkN1GNrvoEevkTpZoT4QXS64Xm5ltOBGhxZKiM3e1jz080sD
GF1X6dB4dAigYUTpJsVj53VopJzljQ0df8s3yHERBKCzh6AqcKTpU7qqHoB7
ndAbNF/530VCm5OqjqXEOEe+id7Jq3h/GN59vWR9jR9h5uQw9L7fRzADxw/T
Yvx+6GZfuazz1WlVUIFOMZeVRP1nhSxIG33FkQBcAzbx1OO6SUF/KrX0V+Sz
G8IaYj93groLhDVNAEu0PodUY9EcrKU0el5VgdM3ptK5YZXoebwbmXlsipDS
awxjNkFmHzz41/aGbGWz4VWo3e6JM4TXuzwL+WrRIjStfm48JZYI03iNDLuY
OwmV60lBhDT677+CMg0X7nJpX8P7HCl9VsoyGfabyI5CaMQ5y0p/uZGphRUZ
kM+v4WjHPneeBRtIE17Y5NYFG4id07FTb2oeK4QapLR/xPqTV3gMf8oZqr86
yZf+Su3jmjM1XD3mQTuSlKkeVaw8+ZX/JKjRN2XPQuZbZ9vpHvLeVQlAN6wk
80qHeLo9+S2vNWLNxmfDyAccQz8yM3WhUDiPe27ZNbaIZV+IFLeLSrFXnRY2
W6lLtziW+V+t9I15024fAj9zIPWdU5xXmoOw7nJfigv1+AjUXiV09b2W7P9g
LIYdlwZQeoDvxtE1V3Kxh90Qn85Hx7uCZZ3Mf7bFqmQW3CburweFMpsMDNkm
UvEmomq8iCgnDGKRwDPlSF/zDaT0rMMvMucvYuI2tmOXP7XqzskYWQhse4uf
UZY5RlJzJKlQ5qQ7KCPSCfoRPWbEX1J945mpJ4KU8r0ANHfqmKO1qa80dufV
bkjTBVcQN7DxbAjyiOvxocKkLAjAMH3E6ncexGI9iFVZtf1sO6sZoJ9EaiOC
11hbcZC2OsZN8+Q9EwjhwE2O73aGF4mY6OGH1r3L/Ff+XJEvAhOpedIviJk2
d2D/kctGqzxrTRpfUbyntQ6a/B3DJrKaAfsjqBojJaUgmeMI5KxsFk6vL6LU
16D+SsCWducPb/Q9R4CrnJ4hRxqEGRgih/Scdc8rsjYFm5RuwGIhKIp6ix4t
oqnBj9b8xqZ5oIZHxKn8be2YQSnTf78c7rsNJ3wWd4a4XMPpgaG9oUzGfzKV
cmyhvAIibTZhFCJ1Z6FIcjgzKGaNoFHDoiFz3jNm6uo3YtHkcSTnZIDHc0xc
8C+Xv2bAPH/+Jm66Rbm/eSEcfMXPxsL5xNmJzn5w8eAVJJlY8WoCWaZZnBu5
N6Npp5AfogZ6mer7/hLKrpTxmmDlV8xdpKj6S4UOtD7gLdkM4gVB6+49E5cU
R5wQq7/EsH6IbX9zV4eQxGCdLBksh6/yJmly6v6Cb+vG034SbLqCKo6hdRen
n3Fup68nGuIaCxnXGb30u3+KDcO4zOhvfCcSn59ds6tn+d0Kwhfpxr1nHU+D
HicJ3LG06Nsvaee7ECfplBPKfXC2KRuSpnYYo6FTpvXY6cVfB9Vagz2D8pOn
+WNyhmfJWYnylxM5ch3M82+mIKVCinlGE7nXwnn8mCWYo6H2eoUvWUXQTUoZ
1HDtnSUAd1agD/6PN3oO9vmCKyS6E+n8PJdwHk6CvxRq0OE/qHzo6vIsCcwu
kd8UCyD/2KF9tMCFMOZgKse57W36ShuThIsq9BENXWiZ4wsR4qkcUU+2u52V
/kAIez55N7BlgBH6I5hkkOU4SXTmPDdI+Y9dLsqR+kqlOSQ5pkl/i/KtPJHn
qd/RjdJ5kjCFRYZss18DR/076BXq4Z+ZTGYijbo6jnVKso5aV9Hrm1PiOP3w
8NZnYfjRMvh+WZXekw3OWKXFhIgq7zB4synKtsA59gnVxbhonn62+EAx09cp
w6Ybd7Zj2eKFn+Hl+4WooUND1XX2hK+Jk2KKFuscZ2p5okAyzzptKZAfuL7b
BZNjj2UNfRynBNU0eJgPCgPxS+TiyKknx2bPlDLveINvbAEbvvB23Agu4Efa
TMVZYsm3FJEN4OO2mNeJ+l0z/B8AimQwBqjCCrcl92aSu8+qtkMEUXUQY205
FmeDjjQi09MUKs9fUo0+uDw4wv47XaY6G4Dmuev8/U2ahTUSdRjVcYeWCsgn
hOp79xGCe4N2b8AjpVff0ogRmosHJ+/8dM+e/JkjQni1vvzjLgnXzaJl3qnE
28LXHuHcz0NGo65JrrwyXILTag6yk1TjHgnDKXEo2mGnvTtTpk7nMbRm0Kvs
NJW5Blv5CDO4ibV0R4RZ1GMwSkPeXXRCUkOfr46eykqpGLJg12A+wwJ3EpCd
6O8rnWyG8t8uhRw3V7x7BULOZms37K18S1KjgnThh6R4+Es366jvUPyciplB
sFy81d61tj5zaE2tDajNZVZzV3NpwVFGTLGmEI0bZM6YqrJyfS5Et8b6FUmK
0J2BnG4scPjo2vAk+lt2r+gIYpYMOLlWXqUlZLFDBO6kIujYvHDMfm1G7+3j
AmiHrFEA/zy/unuYApI9JOgRDeYcvS7pDTgYJKomuO/HMwAJpu7gmH8MYZES
PuhPl3nuveOr1N+LkCqlgVg9Ox6eYNwlW4DQ7Z1dL45SRoCnnkVMi+2cO0Gk
i3T4WU2YFWgrp0h7AHcD26ZPhOhxwn7QRT7XXZt8ersi8T01efiLKXS0NuKJ
HKdhNQQsS7e2Qn6pItfdB/nIrEYM1Okk7shUZHVq8vcIwv71dPcHklo7qXOg
Ls4TN+he619o9EE6kxJBR3+gSQN4qaXmEEJWYFSdz/LZ+yxk41Nhrvbgu2cd
A9HXTHrJe+S3+beZECDaByfv4sqGdeJsxOuxgfg49mhPHaLMCudxfSBSPB5g
ye3nr0JFX/1o8i1iNQSTrpXh8eFlz2WroTmB/tuvwEwSSP2umbuRCuJfs+Lg
JbbHd4smgFdUhwF5lSkKG5ywBqMq/HHnzvrugR+18NFOtdeWW23Y5BnR+9hJ
CJNat2sxv2zo8q7+I4PFnAy1IGKo74pjmIruGCDXuFBTF62YPmvCqM0Epqe3
fM5NjFLLmW90tBwl/GaidZCn2cLEvKd74rEDZ+ishdsh+uGqcXo2y8YF+SVh
DHNexPWt7MPF43pyGFD5MJHgmKsA5nXGSxXx9b32Zd7IN1JhsTeQnyq7Y60o
JIgIyGKAqxebcc8N902S5/wFjpZgyNGgPmBUZoqo3KS78lIkSmPbcB5eMeu1
txh0vRJkhT1N/26mfjWCbYAkBSa6vJEZSWBO/ICKmWnZ5pour8hyj5WIynky
+z+2oEX5Wp0YPGCvtZ2PZvXdB8II9kQlptBhE0E8vF9s3Uv0UXKccMrGv4dy
eyQgbEnU1z6vuL0QcFphfjdCbIZR/inJ08rIat24T5azTS2sFYJRB82pkFnl
HLuz9n0a9m67/eGRbxDNJ4acy0Cq+4WeNAT3tqEjweVrvl4avi1X6VRbaeGb
eRMt3pMBLsmDjyh0dwWr2TDFdpSkncIWUxfY1zqf24NPC9l2O4Lj5TB5lwuP
45pfDh8YPfnMl7EWodsO05ke852qZ5MaE3OT1kb2JkHt8GEkd16weOixjZIi
YZCnKQvfJ8fWf9bd64f06nYeH9NgAx9zv1x6xko5HU6FMFh4/Nr0vuVrRUsi
lZ+ggFr8qP1FYf6xRPcQeZzpRMFLQfbujq33bSXkp0m4rrV/GvHWv67pGTTb
tByAC8IeuTBn2mxQ0m5HEPJks7z+Qlgy44hyQJoCw3feeCn3PRZolJg1L/XX
akp1z8HuyrwVH1MmKu0C1pksP7I60791GDuhwNW2siQWjbNsn3etyf4G4n4P
jan1yyTAuFm8YHgdS+62grJfcs1kUfOVw+gDNusdyu+c8UhmLZTnqC1s0RTD
JAPBdTHUh7ssvSbzIn9vPyt05IbuPuK9RAZvgf9O24TyFZhQihAsemfii6lV
tMEchY02b6lZw//V+XYwakDyq5/yY0ucD/KD8IuhBpe+UmzdS1En/LyLSCbO
tn91tt0AjrAK0bd5dLq73fpp8RTZakZEhGQ0QZfc9Or3/UzdyMY7GAk02YyR
fqVUEoV7qTff9nLCQD60plUnG316KGJWIgc4uyszK7WUJ5Rd0L5uneb/vYpQ
m+nhOicxI3GIHJorOYszmSnmMUCYv8bLhEYpFtfUoD8TmFQI3bxJ66Z2tK/e
QaeaZMAUm15YVJgA2px9otmzr2MPI1tk7tp2GWcIRosqY7r6Fwdcvy9SF5bi
THVGjHR1Knv8jbAWSx/Y+sVJe8UamnleBNsNpDZgFhjLb3iUi8hMl5KzOMvf
upooatmAeZbpaOutGBv9Ps2bx/1F9C7Hwtk6i+e038PhPuQXJJIy/toBXAjI
Y4z2MdILcCgDSdPZ2Sr4N22Lj4cbKRGZDyCS0uHTwxAvbY5/8sliutlkqxP9
0Jwr71xcu1r2lQw45EtQMke67GjkpBTbsiZJYGkwA5rPjC1cWj+kgx6mzylO
BZ5XrDPPNA7vWcAwDIHVM5Uv5YILiXjyCXflf0BoZoCAZEYx9G2XWFShSD7e
UKFq5y7i981NmvVuNFDkoGw41V5jU8rX82tm1BmDCOwAEMQR2fyDGrtYDVqM
cC6BmaB4Y4k8VWdxdLgD0G+ogN9s9FVFKQLNJ19HTzAbr2TdpJJ/lVTHU+2v
toH9U5xjf0jpK1Gi4iRabXjKpJ0HKV7oEXtihspkdWMhi2quzbkvZc/DNHdE
LNIiTJcNb5057xT3W3y8AOfI5G5KqVTBtrk0T5FOhbu6gZddKlPuHjkt3cUZ
jzU/XP8DmACBgF4qLn/Ff7O1k/sQsrGWS7ET1SkUFEPvYMtQbkJHYKOfEMqe
Ck2FrWZVfE0mdStVQsoVlaasDtiwBu+mzoPfthHQrhqcQYTo9fJX1e0GhxqK
m1KBWKr9nn4+VoV7ZW+BuJ8e7eeAkImjwWi+fkOeBXKpbABiPMixXTJR4X+4
Y6uxv7rOT6RAECeLNqagZGnuci0X4gzLy8Z+Ogvdb/vcHHOpRjKZHYIJ2oEd
82mAa3bISgiBSrr4r2Nk+nVv1N+m1WSMpl/ZGSYdMZVghiYIyU/IXye4oE6K
9EWwPZYa36VTp8nlfqdoosYyhzrorrvCReU+MJ3+ZlkheMAiA+vl5TCeR1L/
0ATlEM0asOpCj7UtgjaOaqJr9+srN0y9Dg0xziOy4WzhoD1o7Teyln4bRcfx
axxxBe184tBtqB5FQou78J/DPlh3yQ+uIitC28f6kcS9evg92E5ry1nju7O/
gNpR7ByNDFbq+9MDwxe7W5cc2fz+7CU6C8Map5tSNqnFYpQ6BazOUJ3GLzRt
4FpKXWQl18NRjLC3YQf9dFu8y7RrD0CrsUka0DYd1Zlo8o7IKByEh3XUB1X0
Mz6EpAUEBJsEbHio1yaOkZhRMnptdSr8O+6+lwUOTsBEMcz95ma8QXMwGYu7
Hv7y/Je2jFV9InQ31BDhe1ZUS+k27woLR87z83+W+2/PD9QJ2VD4DiA4XLx0
GtE46roG1EK0ifBU8ejY2gew+1VCP2ucvO6CnAyxvwB7SMEcrxEqVuaPk5A1
F+CUj1amkaqJ9cTBPObDz9l45Hzt0VZofMLB/NXlQpT/Ux/Er1282ZNU/o5X
NKgcpeY4iThQB2um93p0IwlK8aCHepatoz6gt6+iZ9JTqvDGJ/qd3Dlkkdxp
zXrHmxdQjDD8vhYGflgMiFj8ytijXcmPFwC//FUZua5f6CGrUHDGmNkplNeR
etyC42U2lWWR81GkKzl7l2EEhsKwunqFQkrjXFXRYeg0escRIkohmyJmex7G
nfTxsfAsEQtKGvi3OZVqWDeidkOvQVWwDS4RTNKlNdLv2X5I7VzraHUuCxba
2b8VlHMXBq54phXHtgqRMk2hbxrt9Ourzh96Ou85wF4pkTbP62EY6s8PPCoy
+caVHv68F/Nzhn/3w5UE3DRZH32ZjGViCFQc7+yaY3xGzAiyUsNmmrmc+pKE
oVGmXpKE9b+wod3TL52NL6o08hLQe2DzNGGOl1q179z/X2crZfvGYWxea6a9
s4tCj46tiahfgiYwlP8Sl05i0mPQ1bF13SbHoOcLRTloijB4RvSptdyvnlxm
8O67ucciAjJN3w4VAnHkcbUDogU/uNWPwB7kwDbygMK/mF52SuGfuUUHpgXj
0MErNSJzsVPvhXOalKrINrbNUGZxqUpdtK9j+ocCl0xcdlGu8RhVhn1AXyQv
MZAe0zvQabSsD91lhIAOmhgLq0LRe0p7oHpjIFQ6/KqNstaCl6Q0Rldfb+GO
EAcl8EPl8gWs/puKnq1TwE8B/DNRk/IMmfNGId8JGF6idFSK7xSDGr85cHMb
M+UL4AluKgAFT43q/frHrRYy4ZGUFwJCevETRH1Jg2Fw+gv4hp/O0xetIILQ
ajheMzP/Ebhqz9PSvQKxe1/VG3gf3IhHjUREAok3J6Z0w13QOS0/u0f498zf
1opK7cZ93YlJXrxJ3i8aSu22Nfb1C3AeN3ZCN0s8MedLSG99C0un3ruPh2oM
E+S0ApJCnNPmuQa+0qySFGntbM8emy6+4xWjRyUi94QdUFD7aqntdOzAZCIV
QlW4YCWe3yt3WE7V36JRLqNFRJXQGND9G4AzHlTEDdhaVPlustabUBZupk3O
bWrOG3fK/9ZvVchTFFuRdbJyHpHAWBvM7oA01BQ9e0K4hUuOnvoHOIA9zCg2
F7l7F7fRa8Ysj5UbDseQlGxgXDYNAdHAbPts/zRv1QapoUN1zs9TiVWbO6mh
8cD0fKoMkLNc+MlXVbvoWlXtDd3/e8oIhB2ftuxPVD+h+aAh6ia0KWw23J7V
0hz5IYcyERmUj6eUPV1Iom4YQtwD08RprZ2ice/bVbRTulK8KMJmbY0Jontz
hvgLO+vtO8E1cLmTFIy4PEV7NXesw7jriZaIdLCy8wX7fUW/2uCNWUT58kwZ
jmg2wd5N8h0RK9OLW4TzEgKiJ44mxHsUSdzpqB1T6u2UVN45CcYUdlZMj8EH
z9QCiGj6HnT77/YEJb26sYuzDkElF27GuL28TESYnutpFngIW4u0OJx5sWle
PujvLk+LrJR8wgqZLXP+fglqi9maolOilEAiUO0jOV2Bqka2rGfr6DoKtJOT
rTTqm8n8mBnL7GoOJVhCe3XQLSNgsm2cMgWIo5ZVtYC4SjgrhYyyuWsYqTHp
YXQFTDXSr3teS5aTtBAd0WGPT2Zaf5EirfnyjqGld9tpg84EL6TfyS3nD6la
rXvJuVpY5AsA+cKV2M/1d/M2Ltg5LRGSdcmNY6wxMuTH7l7NiCUv7LbOk7L5
G1LS8X7r/iYYkStXZAwAsBHDCgRvmJnfkhfX4JhDz2eC4bNjGok9bMKXQYSX
2B4skx0XBf1c5N0IKVK32nJ/PiSGWP9P/4MPEnzEGKEYlouLzyan+GxLZhxd
+qnp5vSIoNm1Qx5aE7uhoO3bQI6pz9Bimpi9GYD/LeZRjSrnCKk7aWrtddJu
MgQkMAImBTjW2hM12Z81Wqq9OomT6rujaNN1NMarjjSEl9z7Vg4/QLgLdcCk
/sDmF748vpfkzh8rQ8JH0vaCCIbzjA6fbbiXFLkA4jSbP7ZvAZClJZq9RyPh
3XfhfYIgKtVkiNfsAIAn77MN5QveeQGeTQQctrbJtTWMihFJBnRPDc5Hr/RW
x9LlM8HqdI1lWjeK+aYPhmM4/U5yZWpkkoSwWFooMAw8Gt9NAG7uASCd+xxB
kQCY7KVse+HjEfTP2qUKYgA/pKKOPbFcGd7tsK8swnekysXZc4AsykfKq4Ho
qhU8OLT53baF09DZNU45qj3XLfTtlNrzO81pOwMFCzdPXboc70CF3NjFfo8z
e/yA5UUuhVRDUxogbkiQR+nUTHMdzmfWar1yzuGBU1Q7/wUr68SU32Nok0Pt
k1uXn1cxBY6SLq4HCPKzgYneWa4rVpE9oLcW19QQkFRNR0t1rpdm6Up4/oRn
SAB/XQXB2winiAU0cjjX0z1pn6RMFMCfYKFyeJPjt2Ti0PUUeNjCSUyLC5zS
DmqEAxYUIIvzOYSxNFfIxlTSbLAd4T6iAKuvge+K+M/qacoQlprmZd8eezH2
JnKOFCu5ZT62pw3VYbTeS+1nfbqEgLe6JkV8HgKeqVnwjVmYzbxP6/8meZve
zYE2sZSk6x7c/Wd2Bx9OmiwtSI06TYR3WJQ89X68bGC5nUO57EwQINWmz8VE
+tOOeLVevk5SofD9asEpJdsJB0xaDkvNJsomwA4QVuX/Xzc7EC8kkn5P096w
89qpSfPX4fWgM6QBWc9DfxbK93PZ2rtkR4gFD2qOh2IXGW+rqdFzbY00zpOW
pN4kGuU4tEgKTcaUu2zhGXVU8vUAP0Bbf0NxUzdOa15dkLAonzy3rkQXbjYD
6+4G7JkpDFqgpbrlryda30o9Cz23AV3Vi+K+ZxtRiby125IcLZbXHwNy5eHI
HgLCLoBLxxPdkeo1FKaYJ4KUJuFyqwnaxUduBH/OynbF8MvwDSoyu4jstt8R
Rq0FLsLh4hLaSrPKYn+ZMhb0x80hcZprmxuqZioX2Ew7zVGnPGim025RIBey
09gv40qIL96dx3nZrhbNJ61jliclnmsNyaRwirqhQoviOflSHZbCBv7pz/4z
4Y5mDXgpOz9DvMIe3eJJGw3eASIO5NHPC7nWIcBaHmu7zdJU8LorJpcaUjVQ
7rxSoPRyfred1KRSO2dmAFyOMPUW76oNSDhF9Rwc2eAuqvCoaYH4xQaPMFH/
xFSnrORGlTiAFugUhTI2FjezeW5/fWeAr5YFmgaQHSO08KnMptwiMWQ4rgCi
BB8KQGzuDl9/RCS7DHOus1JxByMGRV5TEsuy7w0QKiJJ6XfFYS3Tg+pjmFT1
HbVC/VjxMKL2JUPHH8xkY9+43IrQdj0jF9RLraBW0LaY6h9f0krLRTCrqsrb
/44kyreuuajqGmuFzeoweOqsHMNUiQYbuiHMFAGgccI33ihHoiF7bro0pLiG
iHtz5nIghww9UeZ9qEdHowfXa+QBRjORPQ3sXRyjZl2WJ3VcFBhDvy/Hbv9E
TNzT0GuDACUIdQrhZpk3jCxE0xO/Zypjysl+xR/Yt2sD8Sml+AkwTtlTRmQc
E4Wvlqi63vaxKn39xvO3+VyOW7rjEXewBrjcicCauKY1+aDK2L/yIKOOBCV5
SWZDkGOfZN12NROUTjoTG5l2qDemCgS7YREaRSGOu1Ox/m39fmosvKU4OFOG
QJCBNs2ziVDoWj/HS3oEtJmN6IiWhhpBzb7sOptJ4grvpomMzAV0NT6JMvq3
Gng9OYq/8HJzBud8JpEIA/wDky3kIogaa4WiumKCa4UM/vhiHIavGofwWzbK
c7WS2OrpHHNUReVSwlIX+ahyv4xX5EI8peam2U9qfgDw6/LcitKA57kDU455
hc6hqEDiYFQr39nO8Dr21cf4WFXQ5pFFVXe91dsDmkXDDDsRno9hq66JFFfF
RfbfKa/P7THQqYCCKi/X45lOh19Ol1DbYBHrPR/YaSVYbxAD5gp/mDzh6Yt0
jn54+J8HXTjehhblL4uFbzZlVVBejq6Y7kWvCQe3HiXLqf27PFnHbEiTgpqm
sbBG9/W4v2I9CJ8n8MDS+7kRjdd9gsxx/nkWcH8Co/5tkjzVgOJcQ9ZTaLF0
uR1wWr4fMhytoK4ZzEs6D2C4KcyutLX9CCpM5bJByJewD0CDsH2lEtEfBGv0
Kg1luYNsucOyFw4Hc89zjO7PLxPE7GVHjoOhA6Gg916r8XDgOzygt38VxMxg
jplc5jPa5LR07DdBNC4nkF/l7TkSzimSRKu2V2X8lL/ttilL8kTYZyofSdaI
CuLY33SFCiL4Iek57IUySD+Ge1beLVWsrDQRTnJwdLEICCT2TDQQlw55tCr/
hwrzx8NTkyUKfXJifKmRhnzQeyfXljxFX9xcqufCKr9KNwyyPsCP61KCrmgk
g0IGsg12oUp/uO7lLXxArrg05fKZ56lsBgQWKRgglC356NqYdPDTOpI/kDNX
mE/UO/Moa4bLxhHhaKT6Blq6770gMuovZWbgwoPSMYFLK2qOqZ9Nt3XYio73
e4LZdfBtjP3iVa+SNV120ZgaSbbIYMV2+pyEjls+NRfVI3NLbFUcZztBhLgQ
Clsl9O6KH8lzurfrKTMHlIO5B4aiiZ9wNWq+UPATYqY0B25WJhpsWLGKaSEZ
JTJjVAZ6OUdH1rjp86/yefw6/hVJIIRt+ypC3EYVGTyib7wbZOILKutnqqIh
LV1yG9vfnWoVmpJ/PseABVd/JOARHjPQDd757gL23hW3aM4c+8pl1mS/RWd1
ONJ6RkLlrFiscwXeMwvoVB+yd//hOW+j37YTXMW4WwESCvJtoiyhy1hCu/1k
QrcvvVyfe+Ss2f8f/56Rz1G/oLULkZC9jsTLH5IqdEPPniOxmJ52PWQlHAxY
ojnhrmNXdDIpF41aW0DI/FJ6GttreHiGIDmnDpIt2jYFMxyS+4WJxsS7uXMp
WYxqLEbbcIM1Oa7tVOv9Yz+meTg+XlVM8ed0eGYUtcCt/ZaDS7AJ16oeuxwL
4Jn39SrllLVsgRvrK1JjzI1+vJOOv+9vmk3CKEhqinHS45SsXAU5XJnNsAd/
vYWk1s1gSwFdGGPBOMsHA8V+8fZjWPI14C4Pr9Va3X6UdLzTCXQ0bX47Z6Zo
rTpaoLxo6bfeTMRrw0HkZAqT3SVIfGV0a8SVEhXI+8CW7j1iRKdFrhMhMxWw
reKOTRN0HpIh/Q8P96VLKbERIVR9f1unrdHtVwltLvQYYP0qCQJHpU3RBWn7
iv2Ubz1RTkQOiOgVuSMwzyG+el8RKgMPwcC0Z0AZK5tvgYju29t9majB8YD0
RLni8t0uqJd+hTWaGwL5UPqky/G0Ah2HY0MAEgLvgxdtShHX0aLJMQbWV2Tv
9qE7ZNVOX+XyuSeRZpbThnbCfuIf0zUBL7e9kqoYEd7udcC81BzC2ManRZfP
kbcJ4f54GynJmnDwajgrMeRdg5Erb+bl7Fob66AKNgHFr8gS+SXGpzIdOcdP
voFdwFsmc7h1k5DbTkFxTIGNILq8qV+phq5NJa/wOKB4TEQDt7I+uWLIx/qn
GX35EW4AmUMD8Vzya6lDYedAD0joRMkHuUEdUMLeXFyB3Elt2gGZpTqXZBWc
y/wH6HOtnvPT5E3YO66VdjT9yKtaLnyQa9vdVgVmbO5HWDBMXF0sYEIoCR9t
L5MUfFzgJ0dsERxuJDIntadTn3OE8/Kp4dDuvNsfIi66rEXujWPXzNiSarIi
7OZyO/TaWb95iEsfY/ZKTu17OlfqcqJGJEekQ5ZUaieu5gr4sH8zSb2q7EFY
dsjweACToYwSPaFTTWIqofp6RSnZhHW9KOAntpEZ+wq7nPQMAneI0f3lqCa6
UPD3SdG/JdIfWRWhdT9uZJesksMna2Ds8Fe4L52oI/sHtfe+tMM2l6pJrzV1
a7vO7X3pY2coKj9yHJDKFpX6Cw4EdIrKRPWkXlsk/WB7JiLhZnncs98NJ5dO
V6MmHZKbhCtKHeAEN5tDSwWqDrNzbNH/cjyK2hk0q7x8qBTVerlqQVa7sS3B
/JCtFp2sXUql78KUXPvwiB+CWZh/e2r2Ifp6Rdk2cdCIzaM7o15D4h27VyEg
PTyZ91EOorp+FdqjMyrUShxYplpHxyfmM/iLkX1oXl85Ij0ZF7uAQtQLvlxX
m2haKhtzHsJFmM4lXcrnSI6MNZdPL47T6St7Ynu0+lrtXxFxbe2Xnwwnz2UC
yuC58uijrijVwnaiPxKwIPfwM12TSNTPkTVwhpPzOrEmn5o1lxcJgZBP7SWz
aRGGV5HivJQ9ALadbNGHqyNEhxIxhmI07w7ZVQipokHVAeuZCj/mlQ2xutCz
+QtMHCBMEY5ALC6JM0UnPmp6f31Y+NODUsgNcpW44X70DOl75t4eVa0HaR0o
kwMfO6PkR0ENGZCI1RZfrE1a57cTWBc5E7W6lWXMXc5GMrikHOZ7NjUnD1PD
Ql2SuMw9MZdk5E87KmeuU3DWS3UhKv1UmsPn5Wkm8S62t2+acv2gJDIQPSl7
Ywjnp1fSsjW2u9kU2xbgE7jXptnhzSZ7bcVeuT4wC4DD6APvn48gdHbnSDqt
vcydOvVsv+FK7lR7eMVhDab3GCOi5Euc95cNnZSQLENKGaUKvLpr0xZekIsR
/iw/1zcFuF253wGkx9tAgcdKKOUgRtAioH/wc63oa92hK1En6Foh+QCccMfj
gJ0o232DAX8J4kYdgEviC2m80E0SjD3yF1br7w4vnTd/gsZAZJa75/qhs3mO
yvxVXS4U4VGv6u79lsSyl+VXLtpzOYjRMkfBiYAk0AjmBuCCXqcnis8WJrI5
AF+nOcGxgj31kmcoN5GSYco+358Ec8X3xJFUPo1TOPfOTpjG0APqREQxFzSi
LD9MkHIdUYG0f9S3Yf724NMAHIN35SQfASgCBqkRG7f3MITGcvmp1FrKogbQ
H/roWJzey4l1Yi2qe9ZVCvTT5q4Hymxz1mLUJYB31IffrdpSDUY5+7f6XduN
EPjJ6uk098UQd1O6d5QeKi2t6DSc/QPUb2YXdj9LsgKDA2mc9J4jWflM7Ktl
7Iwhy48ki/vK1Ld05iYjA+SSy0rDIDEe5OC+yBtcUn1q0FbbVRMHXurMNQOv
A+mPRoIgJou+zvU1OGD2+3RC4QyUrzAtlsH6mjWdAB9uNTz3snTWJ3Y+5Tn3
FX5uViIiyYo4U4yxinTsgmMKOIccORBx6mIlqcs0cSHsNyyUT7NtuhFU/mwN
LoXx6oUs5iQeoBxl5ryxO/VH7VU+kSXs5qxWtk1lMuYNOuZH64FAHMvN7gzI
x2MaallQ10mzB6tZJXKRQKoiuiiU+jdbmxAbAk9Pw3XcQyZXHr/M7bum7FDR
79mAJHVHAgYb9bVNEN8MJ2BMdEEy38xwINcKP12RHYyBzqLXr6p1B49Mlc2B
pkkBCZK8X7XyhALrSWgE+i16qwwqvQM7JBVlZkpDI69jApA9pSib/vX4k79m
Pq0kz+W1ESUnrWPEXlmAsZYyOGwNmfyRkoOkYPxftqbxvowHJRBjnJIGfRbW
XmY3oribQnasDgwZx6ZVAdTkurisicJJr0E2oYUsVYz9+gGLv4bS+FtypmwR
rXGIy+UZJ3iFgC3YNOM78OZ/MeeKm+CBMTScPJAKcCskE4o/ChbPFVd0lrVD
xqoWDXuSMs7/U/TDdVdHsREdMerUTHFmbhH3wvmeIW0RvFf199Onn8PTP5S6
l/cU3LzjzkPkIcCr+moYQKTzcJusT0Va83/x3jtHLCW4OUXP8dTkbMKnswlY
xZc0bFf6P64tmzZWwPnbuWmIufsxQPL3XFihBYa6xF81KCxkSEQk3XlaJMsL
Bk4YhbhSXwBcrr7hUMfzrQWWiy6AKvIhIlD53GXXmd7zvVfEBliDGB7ifS4o
1q2v/dNQ9qHiBW7XvKhKdfQZAAu/wp5L+VrvTecuASgQABz7oJdUtgdmx65T
ZhTpWOH6OzcBEWS7sgydyMN7t5s8YaWjZ8tJ6N57SAo1dInEqdCXCty5aPcb
wyjPUdaK0opQHqpMV4K2n21V04KcytPydzrz8yeniHS4hAqYWYjyEnptQ7dL
Ja1oJHNSXADBkahJXw9bAZAACh77JrsMlS2k5HI0om+kd41MM3QC0DF0DDaP
dtojO0qjHgbv+N0uVrK0x8WrtqmXZ5becNWcFGa2dv6yqF7yzrIwBttNlp1v
TzlQOS6XELgVy/SlM9/2FeoQgfmzLrVuBBMFFchbbjSm8zOfaR+8PzEpAfWG
O6BeSlVjY8kWcZIvMT/sI5PfLrB9iU9bJcEgo4V5O0su4gCdNgiC7GJtYd1N
uNmHlP5+Kva2El37WkgIgoB/fydds2XvDFFgEWnTiz8dVjAql7vn13EiK9HS
IGb94KQTeiqAyK1TIcrzlNwMPB1GK9RbanI0yYFTGUuq+EhkdsIOqziwrM2h
9vQE0ptgf98xhXtKnwSVdAllylkUlFiYnhFPmzN+s514mk82kEeK6C9PbJ/C
HO46ZTp3guOeoo2c02yN8G+7aTSlO0EXtu/WJycSCvJLk9mtrn1lM64I0z5h
gJKPxXH93uo2472R+xIxOCO0+Q2R2GBcOv5+JS25zjUltW5a6zVZ/fgdpVu9
e+ztBjcecXJF029Io0ww2H/DQn0NQeR+/b9YOJlNKHVliGMWnCdbqA1H2AiN
2/Eabzmmdsu2VAza1PFUmr5qOD2MBGxVFhgtSAcubhQKXURDkJ9ECIl9FLL6
JPWN5y5QeMcDNDZUzWQBhhbVRProEpwag0hW1TA77VLqpRJ/GOZiWK6YSvU9
l3GQ6Wx22/Raxv6SZACkrh1w/1mXr0Pe+S3RgSa5VhNLrC66PNbaXSq8yNSA
1CRtqqeikGjv4qMfAgfAwRy3EtSsibLvjZUQ8BdMa9B4pAUQ90mhyXlpjlYU
Gu1Sb+TFtkEMzgC3nqkFwZtvAG3XOi0OfvShKlJkgdCfrPaDSJHNUrgP5i3v
uPSQBaJ12TXkqzibPdF4wXQ4UP9VOUFU/n0MrAmF99lEup1MJ/sHUERqOxfd
fY0VI+BJClIWhsh+z6CNXzMGtdaHktGhZppy9H1XtBbqaGb+AwzX6haSqUcy
rUUnHn/nkSSIF3SXHHDdcCAZnae5QeHu8egnaYxZUf1MMo7H7I+Nm74awjxn
+0yiLHgNgeFqFXQ697wSUQJwXZ7h2moqxLtMYR4MS5vH1KaY9xEeo2vtarC/
iQmgL0gi1V+SmFhA/wqgXfzaHdHN7L0fGCcLlTLAF6Rkr57a/SuP4rZxd59x
L8DNWA1f9eqEYQbdvlWN5qePGqg1wKSt5KfOtKwcwaHBQ+oGt7dXVEEcJjV4
sxig+8mVmHBG9qLWx7FdMAXps66xXt1K5M9z901axKNWgF9GkPeXKARshKi/
PxUXp3NYgcm3PA+WI0pTZal4IGBhsAB5V7/3La32nXohzefmmbgTfN5qu6x5
LdVyB86AH49u8Mj7uz5qtqeuKIGIkCJu9v49MdpA2gKW6az4z2/A7ulzfvoy
0skfCuagE+4wneG32DZWzUfLdAK9Etkml2iQAkynhI0PFcj1jQkDAPt8PZAA
ibMLM23ueCW3FmgAjPCmRKc1tO/NMxnb7TpfjBd/VplibTUCxh/nmvEYRwen
vkWC3Jjcwe7ZtebGClUZ7odqytjDbW4k9Nu1n5cHHbzk/+RIdcKFtqbcBzDY
kCDVeb50cKL53Gc0fiLxXImrgFJE0xZcbQb+22vjLSh7p35zXuUgkOLllGB/
pfRn7TzujZe8QycZP262KtNixENt99jtbbALapTqqqJDA+sr0FTPrfHcGO8W
YjH3HxzEBU2ILBLDlqpWhK7rgkmb8rB5O2Thj2Ss5cKAKxPl4BgZJ5iE4gqK
GMLEbf0dtD60qler9rozjEGAmTk/kfehHVFp2X/z2coNBGcE3lZi9zq4GVjP
H2Vj5l7RNFFKdeUqWK3BDschCelEO9vUNGRRV/nlCpVkOrA/b8TeZx37xuqq
OjW/BuwH8ENFpOjCcQKDRG3+H3c4s/xYfONG+oHlT1bCqkjMboUAcsP16bSL
QWqiqchGlgLAsZOwPDiyceW6jwEwx7xtwqOHjPwx242cSLB4j3++FJ3MMHl/
eqcnqhyE7NSCylfi4x0vb9szAX6kIgT0uosQCd9yBMGUTf/SmlaEbzb0dmSi
JWIteRTOEChhygunkQ9F5A3lOmvmTN2oyeknX2GXB80+3xBk880H1XE4H93j
62YqITTKPzlTj9OEcB8t1+rQFEBlgHWA7iMUhh3HhTapxMV+q63mZA+REv85
9rbeUwuRg3uv2rv05D1mp67gQhlAyYUdfotwqilQDeaOtUoHuazFOxMtCuqY
JEceRKVnLkSfYOWTf/niB0yEZ/wdEHhBWP1VbTkQpcsj2MUsXAmg+z7D8r7S
SlzSjh6sJj6XqYXrZqLgFGBVDQWcacMl6kLuhRhi7UUx4i84yWDHf0BQ1ExY
Eecrf3+fdEyMg7Z/V1E2E4zFlUu6e9M0nNavobqE8SWZfN4oHI+ts/To5MBg
Spkphm6S6ZrOqISBDGRiCI2tIv1xVy0EUnSUEECIZ4eQPXU7S/7fdSZt+/ic
errZUkaI0Xd46MSup7KezWFM089GCoc9oyvsPIM1j0t9Rum2w0bkmxSEHJDp
YnDtRIlCaaPpixSJg+aDBtcqsGa0rmc8CZFDnqFUJEchG255YzWvS7GauEv+
UsjhmDCZQEszwcS1if7x1E3vb2BKEsCeWVQ4Mvl5K5Yxyh/jMBlwMSPPpMkT
GwCujiVFpMVgIKq4wB3vnXpbhr+E4wUYHKWfv0bO0oqzRaqRbrbWoP3aBEOD
WLtJDGz3rcQY0vkFmus7kdCvAbw770f/Kgg+n/8QmPPqHDPbu406BUzaKO49
O4cDhjpaFp3Bm8T2pjSeEV/4yTD8aSCCh2tuNxgHiVhx89rrxwsdOGMmEFkj
5Pb5F/8jx1V1LS8v8fI+6vhXLyPF617TRhWfYAts6qknbKESKDpOxUTuve2T
jyp2SnVusTFZdVv9lOyFUBw1w4gtjwkseaOBKLp+JUD8CmjZ3rsCT1m00dfO
WD9Jjeqg0QZRTrkxWpb+wE6f9YVEs+sFC/Xpa6dKXCg4FaCSCHxm45zwaN6t
djb7LLXk29iMCnE6ItwughxP/2M1fPTH06PBFSOPbJ541lHCt5ogUE4IbpI2
lLXv2NPIV8C6Cj3/6M0jNCD1LvNj9ta7fTVIEfvtYXyObSEWeNKNWfgsFcjT
lPgUlEa2FQ2tfAoF6POuSbPcJRUjA1SgiR8mlgb7lDTwY+JuXS3ItDTAHmRQ
cWuF/tNelFYUpc1PTEtFYnezwgi4kUJhM41v8lr0gDprX8xsf3wIk1CtkWNp
sQ9c5ZtLJOe/J3NqPVV6ibrfBeT/Un8PMZNHPlc38Lw+bkdPBlC9n14nXq09
Pi0TgkeMt4b3Akyaf3IhRe3EDBzMt1jUxoDqldbn0zcQLdlJGkEXsbeW8xmm
6QDfl8kQZW0B8FLGMV3ThW5zPl839kKBIgfuix56MZ2SAu6EiO10erjic+6e
A42wFnaalTcvxa/+pYs2nFJYvsAOLplllLAun+GrWM6j2hQR5pdfhjR8EU21
4hfbLQpThWCQGK1l58BFUqbvWI0bn/RoeNxuDJsBD+aKZ4LswI0r1s3ztPcM
22gGn223OYpan60aRAM6pibgO14w3hYO59eMh4H8MOuXA4MopYv6NSYtOFBx
y2FJxUXZ7gvW68PSSxnTwBcn4GxhAq17PX367ujVpncwgjNbIzXZncVn2o46
JeYbumH6qCpjgCUb3hIN2WckKq0O9TiyMpM13+em+ExOqtrCi3xiHi9s3upl
pYUAZB7vZjYkGSkEteoCfXobLbWK+872ojbeETg2jdw7v5T87XV9SYtoBhON
3pTP6t3+Gl8Z+oOVtaoZrxvWWsaZ50Kouauy1TfQQdqP7x4MRHdvgM/qekVS
wi9lZ55owPvNclN+F9kdWIYaLjsfbdIQjy5iREArIO/NxDEwxhBY4qXZnukb
8BGDEloEaz6MKAHEPV7l77yy1hozq+Xq63JNyjvF/ttZj6bHBufVzoO8id3f
TpNThJk6xknq034JWI2bIbfG618Fjcg7nS7kWgLOP9YFeXcXqE+g5QRntPos
NO7I85Nbnd3E0s+LdnBoSOlcqhvLNs4Mghp+rs6GepZ37xD8Ggrgz1/z7JVH
46FP93Q2qNiN6spNJ/U+mWoeKqY0iaimvpV1WoNop3GMUf432zGJoq9eQ6Np
aC1bXs4A4pJLmlRH6Tf5bvdiOBBIZCcrx+9FzYkoIUwMuJ9A6d7GGh2HgwEY
56CPrUsVXL+rIPjXbXL7n0SatxPfGdQImNb9wxjp+s7BTOk1kKZ5WDF1FWCO
Nus5pGwxiRFJHRWzbN/tWp3tWLVLHYlALILW3YuXHl8olhXGHEaYldtXbifT
KhY6oQbSLsTeXC8gNi3OnwbDMkUnfeh72WGxHeWTuzPbKa0J+0RXr6sPJDTO
rnCRvg1e8K/p/x1VoEhOg1hGBNV6KEo/hHHXB4hTi6u/bXQJ1LFU+aUoVDQ4
SdcfepIxg+8ctX29AVTCGBMfpTUfz9GsTn5C5xDTRjTMGWvZMLeXWaJRh2W0
3T94UQ3coRfVYEbbB0VKEGZUJIwEE1U+H/MXZ9f7aGVbd8D5jjN+OpnFkWxe
KEcBu0kn28HPw6F2gYoKcwwYDsUY84veVImmVDPoiJjDPkh+TvfTsF2qRaZ6
L3a7Ez9hR98OCspNXnyu+AkA6TG1n+jiYE5Jgllhu2hPAiC85/FWrj/EELkB
075nnSjiG1A5zqCJFwWKCOmWIAsHeGIB43XCXgrQ0BpUDNz9fCXrCzEtqqj/
f1Fcn4pTHs3bes/L0GuSK8qG+pL2NRCB9TYZArJ+4UC31ypZ7RrE4y8xtjBb
l4DKmFgGwgFNp4YKqCd8en/d9O3mxoPsHB2GezZjM2u/fVHpgj76klDivEoz
MGAh4CSsJrFh+gVHs3OL8AMJjv1ewNMvIcRUdkHN+d0yX5rPoSGzxnmJTBjz
Nw13p4uCJZ47427wnXgNkHi60jpuka+26+t1dWd7HmghGT2ZJnTCd9OKGE4+
6N0m05evfWelkdJTvrPY+ZpsGB0U/c6mL+GBqIni5/2Oyal1lN9no/XVH1VY
vticuwappJd7Q83/nQ8XSf+h2+hlOelWqeZzDAt74aJDxnfUtf0qlW6141H+
Q6NnOTnu2tdUCRH4iGoJJLF9CiXxT2F1tGd+Z1EkT1NNu0VnBVQmBTCMofGG
xfEI50LQDOd6QHxpVjafiyw6rB/5xfKGEAkgdk2r1Ppu6AcEC16so6y0tNgU
cgSn13uSlGUhfAj9jxPtsjQnrXsxP3IvWhl5j775mYHmbl6c75pDxVMZs771
N85nA5vRO9s4/bnBPaMR/PHno8Qz+71YIZ/zLv8OyzA+/trZCq0sjnTy2uyJ
ow5C4p0QKecvq+uqe3eiegST5C9rM4CPld22ZPzP9VkfaNM8KpnQjn3BxjJx
xYuKh1EgCJCirwq8MYPmD03Yy9jFhnTZ1daHayks/hjfU9LlhnWMW+5/j1TV
+Z12XOWeyJ2kpzC1BvDPY96iyUAuC3khRDEG56UJ/DWsMgLyYwLYdyPFpfay
9FSLj8mPv9nekpx27oHrhU3kHZ7DX5Xu1bhzsokXorOfxc+7HQkPuGKi95Zn
o/IECM2t1mbg1MjfH4CUgzsC1mVCerKEkZBP5geXmB0gqbT7/Izl6slqd/9+
zTLBFfoKzK2b7DLCGpMxoMfBR04ipFxsXAzHZ3h0E+L/OILwCvv3GK9kCn21
k8zCWYyo/1P54UhuBL7rggaLq68fIHD80DRODdvTCnoO+J1+p6bX6DS0q4Ho
ptd14awDkT8LS1j1IS/JVU5ZLnhiFodXmiKtESEu1JuOBRP+5Sh/LGtt6PLi
gafzZh+zo/tu+RENmt2njM+5Sk1JA8ZvJZDBdEapUQNOSEFv3JGxALXKcA0E
Jf53KC+BLjp0S3i6+3OUU7yfkaGqlGSOkCxdEnpoOLG8tyahmSQJ49rTGsZG
BwJ4iTNbCBcshNjWMbFnessTfj4URNpdf54gygka6B6oWfaqD5wl2uUZxb6l
B5qxGKM4jVD5atiG+lYFasXJfFSB7E3Aog+FJveZBie7nThfcqLNIUZoucPh
bpdgJC+UABj3eziw13Oy2zB2sS1qmqRJQtps5rwYwIWvU9WgnuqruvBs+9HZ
XNJ48Her8wGNRNt1ajmN0EP/td5f2f2pUUvqXHPr9clXNHtk+aGvkxnb3ocs
jScqc3jw74zxTxQpDUWXhpqbhmQTNQkSmScckwvXCIbkGuH7PFvYTZmcsOCC
UICIfikPcEDTGa/brttCYgDwUgv1bzWsWnhL8ERFQXWC9QN7dV14TWf9Z7yW
GHbssFV9zA53qPnO+vRd4A1jcKIefWwj0dycskHPUYB2gv8I2NLWWlkSBryE
l979X0AOPi2s/pyP6s5CHpQEC1jpyBqbRr2hpQZGA9Wna2BQktpzELQfxauK
iPTrQAngDe8Su9sAO9nFITZZvNsqXB/UKWXFNmQg94ZtGn8IqhvKNh7ghZY4
4ZrIHEAuh1SSQvUnNHthzM+a5LWaLt6zpxrlf+fk8HPTbm2iyvperAqWHycz
g7Sx2Jkwo/rIvx8CTtzclLZUkgjGeFPwyLxili/TsJWtIPHIV7KqTrvDek4Z
a/+Au94ypaTnHjGc8Mv/tIejjCtlXAacHLTSiI0T6flqm1fiWh+MQl0aYQae
5c8oB+ZLoxkJyJQkgakR2u5lzb8rB647z6qoZkg9uL+A5uu8j1UoKtBMgXXw
vaUAPjcpWFAYRTocJvQ5wFqaz0jlqk+e8OdGeFFTauGrFSogzUt97639HyHg
5onCgL8wisRMGTtyF8MYsbWwYgpI4nDtXPoegl5yjQ+BlG8b+WY7gxFSxaYk
YoRpJdJpu68WMbUI3vWPznoaxFtdgwu2kONsV69J7bmNffnfv9/iXD5ada17
tX5+ZCdT2W8PX1qMFMwOdw4xHUfU8eulmmnOEOhHDrrkFITiLLxV+Thgbxjz
D/o+llPQxvKFRiw6wg47XgJx9Dj4tvGGESHMre7zQxcLCaN+dNsnwSC9Cgzo
ft1PMzcqNWJPAtxLFf38kd3v7qpkGFbKvRl9B3fBQANZenDiGItK1nKbe5u9
l5O3aMtB9lEEuFG/Pekj2oxVMNGFgO0HKWyXC/s0c1Px1L7QqRgeqrMze5iv
jAxvM4929mdjMQgOtYC9SizBPKFmYIVko8RScRXd2StEcY9iaHpE2mr3G7LY
bPIlzD/ash66j0P9g7HnM9g/IRQ/rZUdOOLJHAx86va32kN5akPrvrVrmG6W
BzzfE4M+l+PTI4Bj54g/DTNH1ipMrTkDv0WsRhT060PmpJsAQhf2gX51gQCG
xTh7/+E5s+Jly9HGxsgK2/W9THnksG7XJhL0jGIlceAGpdtzNNrT3SaMNcuC
dz8eMO1sSt/8zyRljULskK8LPFzx6/FMiBlOzmtWJmXD4xO/48pyOPa65V9p
6nxCcJAjN73J3umRGhBchI8eqjp5Ck5bGKyxsKR8bk2eD2QocDXf+3BOh/6M
wZh4mUMSVNNr8oMK4iWjpWJ/Z51NfMFZCDZAbCBCcjRbh7f5Mtt1YlOYHK5P
W1fEl7SxC1S9Jq5fV9CNpiFLmDTT8vwRWGVT3ZnhRauRBcn+yjWjvGUY+N7Q
1yjXr6fF0Zk3lxtA/IMYp3O+UOxGlvEUeHCFs/aXzXKygEzjRnUUi6FiZGte
SzkWxWnVklITsnKZtpjPfrPOhAqSi3W/zo6gytARUQkQBxlo/kCHUnZ9ipRf
awjc2Kw2Q3x4m6Zzh6nsx0mzybvkpbveL5PRB0QE2Baj3yot6lmyeckT9on7
LE3JGXDbEWC3TMTXk5ZjvXUfMI6xaDSJMs0KvMHGHsmPSwSSxObJMxgvZVvb
Kd+lLfT2p/bHpflXeZNyKABVxEW/iWnHL70E/KOeSh2RtH24Kt+6SDZTZpCZ
FbXhgVJloMHMUy66vCUf6v1pFiV3fPVsvFKx5XD0rbQ1Beop8rxkpnzDWqCx
mgHmox+b3gBTfV5uOahS0Ud1FGXfSR4yOPKCbZ3dNNWuNn6y7U9J7Zf1zGQa
v1CjzrBoNnDS3uOx6rfWLNLoZlQJdrx24h7YsP6RoPQNF1v71Xi3C3ZWWjTX
vzJq0tYHXopCJqUW5CAP15cZtboa4M8uoeOutfeTC3nJlI7nbxoAfJWkfA3M
mY/vhIteq4t5OzEnOeKVL4sdmeE8YCgiGyLwb6S5y5GWCPvr7bKFHi/JLPDg
kX75VZsK2BjTwlVXM+GZ0lpTi2/ihiKFPErSLK7GStRcbr8Iqd/wd51BXQZM
77YoVXU97nRWiI0sK1gmG2anV5OQyHOqSA2thMk4NLt5WosYJiMk5d1a/qeM
KC72vkD/skgt6lPMOVdShNQiuHiwxxuyv6XW3Ym4+IBIqdLGZu2acO98zZWU
/HNZHpHiE8zqhv3gT91Mx6oaFzQsUXy7pPa1lV0j7hqIFEj7W0x7Xn485g7/
3uY9zDK9unw1GFoFGeY0M0D+17KxXFPP0GiULmbJfrYmXwM549xPIDX0jTH1
wf7F31KRoykaUlV+L8K5+0A6drCd5NOYXOwx/MhSQyubKbzgogXXansVacBE
/SnddnUQhBBuBIwjbA404QhuWbEnq8wLOHXiH4Kec2x4mawa67C6qGJFuiSN
j3EzrWDew3UpJJf4LGk+y0mCadTFQPiJdFwyyLc3KZDsC2eJe1bF8n5lam11
cpVb6eZu0yPy6TrS1Pu6/3jwEFwJYN9/B/u4t5yNixwgfAgr6oISB43D+mFc
jG9WvV98+30aLIZVzrdM/8mLGSKQltUrkNlNOwBLDQlZdqPYz5IDSeQIbT8x
oTp+m6FvTUjhQum9y4Wrab5854SHtchJbiPis/5zDdqs8fze8krUiCUFxv3l
GZGJY5341efmArovFP2xFo6w61aJfqRmsyPEkLApVMc8GeVDrmQN/+Y/K+q6
EvwggABSciwqEzzOHRXGQvHGJLSX5te6FQtT5Mria4Z0pmmSzAvSKoNCCjdq
8v9D4fgr9CFuaqKXShzcDy8Ki2VcCVOBtHXK6mO/LIF0CfhmFWspS4+6RTi5
/1UPRrnEPjKLTAm/5QArjKASjECmdGbHz38Wu1D0MpGBriP+IXXPipiF+Ax8
QylS7ExW+xVfuFKpDe+7ne/K4X25dp/JkCBEskfZH10H6pNGfkoPv2Glcdkt
OLctL+rEJtJ1Yv8pBM8uePMkZriLgdaf7f+aSZioyhYeqP90SDkHX9yHgxoT
4jSZvj3NEtTevpOMNe9tMB2Vu9s7Zg4foEFtfw8hWGroiq580a6rPYRDgzS0
UJBcnEMp9RrekDndGLh1E8zNDb465nwlBpTGT4YB+IUM4Qr/wXYlHWo7czqK
iQ==

`pragma protect end_protected
