`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
qja/Kd1f8M2d24q1jWQY0AzKJeL++26a6wCW+tduG5/rO8Vdgxzb8azCQ9IxJZQi
rGFMI8ArCqKaB3qoeNKq1a5m7Q4VGxLhl3MdIhWVNFX5MCudATL81O1bAKbPPmmd
131eqmkq5AJmxo67rqdbst9dzW2lyhDXJisrgeHZqU8=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 8736), data_block
Uz2VnSA0CEfokCP01Oy50qj3JmpEm7z0gVnPzlSeMM1XT746ljmFZnK0H8rxAvaK
HnFeSS3uDQvn5Zmyk4ZphljY5UknEMZ1SwfYJPwjgXdcCMO62RucztAcZ/FjKbpv
7c3ZCjxB8pnzvsMvnsF3L4L5XcF/N9cWln3Qgn8Zb6+BYjKzCp7BFMgxN84bjD+C
0zk/C11sJWLxut/I6UTtw2y7JE1xy/sSH3EujoqnFd2bNWzD0aqBzUMJVZ8tzTHD
+ANtubmDYJzunLfLdexFOI+KpxmlNsRPs2upHbg1aSRKuSyBQGWxPUHcl1Fx7Z1M
q5tH6Yy5mSYQSJ9NOH5APmsfzS97MRRnVji2qJZwvXCW3wd0PhFnPfxtA4NzktrV
9jxxaxcAQ+o8nwpzAPaOqXYEiqCr9PEcG69OA2yDK2MWw778GTBFN1n0PHuFYICh
f7tEh5wCEY9kRTMf/ewt1fgG2yQPKVi2YJ1iEGXSJnXmv1QXwOaTwFVMtCzXRGSS
82w4ya0PTYSGbQbdooiy1wsgOk2Tgw39QnqMVNZfjd3HXy2/c1/SAHVTiadsrFTW
PDLBHYFQPrYMdi7YewwXWgflS13shcyLCC0nTnLpt3/rSu6FMJoPqZ0nZqqVT9Q+
VWyqJcupvc655YuYSJYaJdLnhPtmnPmEMzAJXE0GZYYVhUvpeSGeU3ijcDrUtzNM
J62KaVTiZYMBm3g9S9BFcdcQwW7hsOTJzzS/w25+bpkd99ShcNsGkCrWre+wrdBN
PFHzWmvYEf3vPbwXk7O2GWM6FbDnymEFVSEjknncy8Fg6XEtvIYX2uAH7EDLOJy6
P4dVKvCmJebPhZjvcpFKnO1T39sLD31glyj0M/IP+4pMaNTFBwaTfzZn6rzX/ub1
NbdMzVihujOJFzamLXqN2XXdzeSX/VMRwyJAZE1E+IFiFvxYqXjDH4gryC1a/FW4
DxH12H+W0hEJ+Z0iBirSxlcCgls+5pg5j1VpqMJq4hBecug5HnJMMW89XfdPZoAJ
8eT/i8EaEBYliQcQWq6yr+8PZpT0aRjRlnAX75LAZxLdG9RPqErFY9C+TLizj3Ij
/A+lsmh5FhG3PMgVfTH21DdlYHzXaqDz5VJecy5uFU6LoT4mrNWZZ+uxF08H6x8t
r5Z0DCiuXjIZKwSQiI934DIPXUSITeNJ4rarJAR6GzQu1ru7RdR1E7OBDcjqPWRw
z43/XSs8piqbC1JnQNkIyyKtBvFjv2UVHd7l7whtaAX8srLSTiFSm0MA2sjIX0Gk
uXVJQG8ylCYPidpKny+ZP9KVwUAD3JQlw3aojyg0Tmdy2+aulwWWjZw3geHNhGPj
Bit/9xMk7uwnjR1rUU3cGl6+lszfsVmbxTJ1M2nTnEfCjri5HjaRW1V0zcCs3/Ik
v0HGvpEDNvNk3TaWhs9zXAubP9kp4KMHCxqDySNpKw83GdrH6voqj2LwAq4cwIhW
xPos3C7CpDVibyqpJsxO17KjuWRXkE4uCiYOAL4nofY+O5dMSxzLHk+elbKT+mOD
ZOiSN9cKkbZjHzy55cflrPEFR6ipc2TUOwYk4EAtFK7a0VCQ8j4h0xHF8Ia+wvLC
/rBNwRtlN19dronVxFAEAFeNZmr+bmTh5yNpgE5OG737k9WqnzODILCUv8VwN4zl
eX70HBi1+vxtnsFxd5L38YF4Exl93HcW6SAgmuNxmoFkQ0HH+FO7Ps/LcpMQhp+E
qxjFrtWDz305tvt0JkUy1Ucj+zIH2T7PPwq5oEutHAoASDgtkjP8ys50MNvkUz82
0sbRiotcyZCEemrRPWtUo/mA49NHYqgTf1HQnJm5KHBOL/uOQu4OjN9CRcQaBR5S
Q6rRHpJ5dVqaGJFXyBz8XDeTuA8bAfBhYWBOLVPwkcsoG6bQjER6z9+SKdP/7jCn
RiOlAQNPdaLt2X3CiCLkB1mfpgshpLnwnq85GAsOlVhC5RAvWREwwgjuvptOrpg7
0N/iHazzh6UnEx7P//AzGEj079UG1gMXETpktIaSx0Pa9b8dGZ5ZS7Dce5SQIfNo
kOyih3PCj1DuVj6t/GOCQB5I/sEB+a+MEfo4p5Wt9WWPFZHAmT95yApnLAj+ZUNG
Oqq+RRilLk4MkodCLxKfbNwIQw+tp2ANzIioh8996oxxbL4pZiJ2+BmYFJrzn8++
OJ7QVH7rGm7xOCVbdBxz/5GUQfazzyV9eSNDKu9Fwzs+zXFjdu1uZakTB++MS7/h
fywiDzoIgQTJ7orsq7MoZ7Vx0KRH24ESLbrJENqdrKMCex8Mo7B9pvQ+fNYK8xp1
ZDxr+NoXZzrnLlaVUmJJMZpJVTfWa50ic3piOqeHnVHdu39+3OoQpS+rsvF9UixR
pSRgiWS0pDORaub+bIyOntd9yxbZ5Vgh21D27eGJPFbTlbyQLBvTYPPRKBiBPKiT
4rBohDcrXJA7bNb7yzyH0V2YRdhA7INilANY3hUSFWAQlKiRFq/xHukmUllJi7fr
6Tw0h9z62S6hjaykVVwL2sRy7psZ+mLgx6pov+FLrpMS5k4MK8RbQe1oyhEPQZU/
YqsOPIHxQpWCF7NfwoW74P68weNRNoAeD0TyhOXnohs5hNK/M89iOdKcxedStOkc
Xqof7H7BZJs/bOJXptgX9p9tV/u1AmF7RpMJvZgIUNdqODuzr6eAUnHnu4Wr9bMm
jUYTUWan9dNU4xgG+a49V5qEYPK/3TCLXBIx1l8SrXcK1k5KSLsr6BDs1OeFDEEj
68fmrXeb4RQevHUisNMRKJbFbIQb2FTi5FMTSOksuDqhCCOSRgeuTgrTFIsuupDZ
t1ZEKeOv4kJj3OYf64cBQ2Lt2jfOT8DuOiUpp1U+wchmqmOb6izrbEUj51n3H+zI
CTkUxZu7sV36JJ5NfbTVObTmt8oJ1RLGT2VS7N5uwqHl9ICxuvunZE5uCmDfYu2+
ioHN81xILoTuWmhYtxah4WGg2C5GyYRyeeK4V8h0tmG5eavt27MAwrVH4Oi3kiUl
LK9rDULDuiudKm9SYJcNdrv8/Xpq4ah+MjVr6ZRy0OVNxfw5sJM7kQE1SNPs0G6f
P2QIeMwRrnrlWSVXeHl/TpjUY8Vr4YKoE9nNpojY+X+m5CZFpRSZRLlzxkldYKXo
cXdbTCRDvCuOZbxbfRcMgCVMsSK2/imKlTGIFVJNxJ/Funv3mO2PylFTLJUSNPZx
+V4c0xEgLs5fTq8ZLpTiQwHp1ON6VYT3A9gtwLfESti8x4ab86bHAG1kemxCqT7X
rN1UAfs7+8V0Tn/+7LGLiL5hk57GZLHh90YZIJIe4W36IWyj5+CjVWVpXXdXx5ys
Uphfgbh0k16BxZ/gpbH+G8nE7wZ6JtwB4FiXHhjipCBw4BGYEZFQor7/bKy50h0m
O6hVWmXtxUshLzut3/lWGpQyM9Px/kvT3AQ+4XEPXMhc+A0J4ZvQyvVccd2JBXqA
+5Xl+RcxJBWS1WML0C3yti4/WlUqVHXe+eGCqdqalZmRRxSmVhJGNHixDe7i/fQg
3WK6y4s1zB+KmgWEMOPBS2gJeaeJLMIDUu7YJh9+0lulmHZpRa5RzIW3UjDZbzYz
DA5EPvP5QABwim4AzqFm8mEw4LyUBpgjCuxh+15bvpkUiLmCBAHf6Jgg29QQuFLg
HFDFRs4GHSpdX5pKHTKjcHP8ANq8G8raoDsuZ0LCmxlKVZRn9wHOJV18SAEJheOK
wWkzu1fFKZ81U0CsvAcwWRoADTKTwte4NdV2DWP+L0jRCorDIyzpqCtAKqBAzPWq
AmXM6rdoq/WJrpjzgAEe38srb93WitOHdLvAV3vMAXlgyrqKORDyX6PhEhGmGoLM
NnobA7L7mKYo9/Nv3oArV6/bJd1LF/9TrHau79Mdod1CnFXXkRe6K9AoXVUxaOAH
JGLc6a197NhxMc78iTzh8LDkR7kCl5l30Du0gOA3wY4FD5R4bkZdto71qI1BhOHV
+aBWr7z0aI4xS1SxCd45FBcYj2Tj3D5pIFtYmQYcFk0pGYDpOWqLv3W6LotQjBAJ
8vx9r3cfLUdB8VmE1wvsUOGGK6ksQXAFCAxThZR4YU39Ok9CN8k0z58NT1iyWnXG
fkSaBZwfgnB/VXvqjYKW2kHXH0ubn9MaqhHYzCnEpdaalGiFFlx5iPmsK3Z72e2I
cDVdCcurTvIRg1BcknlfUEBwu9lCHvGzHxK1WR0hWSZvexUx4PeYwZKeUd1G9Mg2
73IUkWFpb3DjNmkr5L1QxHRH/g6o955fd4oMn/b/x+4dyZSXdCR5QxgkyVsw/Vum
49qlpC8YbuiUH0eiF7dANca9JYtaGaY2lzWVdy5V6Q+oz64RigpjkaWJtCZPx8FQ
X8EbR009a16f78f+lJ8X2AIygDcd3QFuIdsY1gM8q02innynFnXGu5Ksni+/KW3n
N+brij8FoRmIXhWTUvpIdfo0KphLrzw0eVnb49wLhnP1laDE0acipIULEGmojiFU
qcNSemt1yT/RPlKjJMJz8DmbXjmBYNkZc9lZyXKAmd26xxwiNOxrFy5Nxxe/7zGf
b15pJwJZZGYEBlcaHd9itIXZldACdGECPYkWefWOYKh9xi68e62su8rYauVy55/l
CAxVGLXhd10Ofu6Uxw38lARs8COCbPGzdja1kujKmG3YI3iPT8RNzI5Y1nfG3lj+
Yz7vqRAeVlbgAsIQbMGWPpPqCAaClTNVyHTXuuJrWrnv14DLzGm2NUqDDbQHHA5Z
P9Lhwa45Z0T6ELQ/QSn/0UxZVMMw31l4QrAuSevwYYt6DqZhiHkWeloGssSmrnAT
f6M4Toq64wiNjrXlqzMED8k+IGC8hWYESpecuyhZI38o+Ly8MTpxZoC9rDcMIBhU
rzh8pUW8zTOxOGTksx+hoOZkDdggoj+Bt3C9QpbcHQUMqO8FPlozrYlT8LYn2HFu
Fcvv680/v/NEQLaEOaWYyxNferLDN6lfmIqEnMyxZK9tW2x4PqiOEA951YNv6Gic
lnGhweySVs41PErQ92kwgY8Wurf5NmviIArnaqxhlDuwMZuO0bim1b2+L85VRiP1
iX6+v3gvbkh1diRER0mMWAnWKDy5oJDPzOkVQ8vcUBjSn1vVxYOlsld4B9TPUTsP
8B5RT+C3T2DJrI2KfmHKX8dyX0bfj1R8DcG23zf8l9hHi5jgktaYXgCW/XK/nHbM
rjbTfHMj7WKBq4E6iYq3zqF5kHCfFsZT661UjG1X0fZB9YyHZxCE22NUSnaIkwjt
Rs1B0Lyo8JxqgcIZhRmNpqKWCDa/jaHhIYmEc6H4lClm051E1RYui075cPeVZnId
m87tPrh3GOSL/tGV6b1BpRlb5TS3x1mEwWpyOJBgvma+W52hJW5So4F4kXVyYm25
1ngzcxncSSEgqaJE0kOSWCWHgbBD9qTy5ZJ633nC9R34Om3AIH6q3qfETCHmoxva
KJjhdIMEXClmMCRs8F1FiS7ixhXlhI/X38xkMj6Hq4tbmEHXJs1J2Bv74pcCh4sp
Z9DKIp5sg8X7kVZyITU4zJUawpkC3+0VKxXejpzzt0sq3D4DLbjwjWvwobitmJZV
Mt2TlA0ue5WaOJj0gsqXKZeor87jRdSoBVkDt+q02E7SmmoK72MNMly+AcxKYHIx
/3aDSwJHpxHW8gCvGKTHz8Rbqf8HU88YiDVDGeDwILb77AjCSLOMerNQ8sQEEuK9
y6oBHpsfzcezDHwgzUORdKRcPlEONSPTres5mFpgdzaoJqQOHQFJXO27oqSdozi3
1Z61xhIereIxgszuqGcleTJ8eBOeRg6Ld3JhOR5dIYPf4DoLXSxytHztjWk80UGS
KqIL63jcRjIH+nqMXty8Fl3BIDW0xo9OxfJB1gju0fL4CDCuFB+fsMLDzCaj1O59
HMLJkgfMSeeUGgqbrfczBajBuLgH1lDzu1kZomoHDPG/dWy4hvzZmSfceFzqXu1e
xs4VuqO3XP6yqnwcp1MKg/8dlOSPEH9r8Hka+vXHIJgU5Nk+LCpg+TgrvcqaljTG
J7v+xrZYWJelY5YuK2aeb6OfDGa4Ym82RGESR+a9gDZ6b/+BU45POWIzKOjl9PZs
SBjbbRz7soj8tvE4Y5I1vl33874jRy67WsALWf2or0CeS/fUmjVdnWvSWfGTT3R4
t3pvvs3joScHI6+b56qt7QQW3b45IejLO2aWJ/OJso+JZEn83xS+W3LPuLMq2TIJ
zjfi/M6kkWssHy41dlcXEXVi/+tU4KwK3NaVVzhcvz2XyZJFWRJdwGZPZTd9/jVQ
YpFkOMA/ElyFDYqzYc2fV1HGN152y5GlU0MDj1PnL6BoJEsFPb+ZTjAYO3/k+W+1
c1A69tOaBo9XlYYYgFmjn+hoCx4YOUdHI2CeG8LKS+W3PRcf6fJOw/i7cEabTzZy
4bJDW3Kz3oArEJV945kKFYHhb57IUu3Ktl6Es4PFXuouNSdp74HibkZ57JJ8Cb21
jGqmovQUQJp6ie+UeutLodEquJqDhLR9FfB0qsSfbfkRPxtZj23ZGtdpiEA8lBg5
nNCejNQHYQO6f6afwaIyHAO27ZpUzWfHtK6rXTUW0aTsYtMd4pQhhm+m8nQC7hvW
fiaoT79vPsqB8OHbricXwyD8/defgjQXkSXN0cl0v5qSo/4LFFznUsdljJas+rwG
6+lBezlR+6HOqgx5rHbIwj8UUUH5oYGW8r2+9jtufJcs/IUHfO6dWgNRb6zO9fmq
RuAtl5HZWUce48g6Fa4ejGzMWJAr/31qtbII0MZEiTPprMO25gzClK436rZn9M+V
PLw004z53SOc2fw7ZxWN72LyfoRzvGg7qUPAsTz8ssnolw+TZWUZbNqAeiXjFWpZ
v0l2fZxASFV8HkiUiQIzH62dp43TBDvrz2AxiT+ETjY3/a31c0Jo7RM7z1Xw39cM
VzUg39GDHSCPqiLw8uHSqKO/dO3P6xGrJCn+STwmON6tFTSdN6xAyAkUz1RSR1by
OJS4fsjJazalRiKpiRU4bIaY8nM4Wef2J5xbWjx7mL9RThXuasBHGj8jTtPRuoME
WKUrKFZ+7R4wN4DyHeGVfIru530f/ZIH35CU1HweSodQBnZTc/bKtJPqmrvtwsz4
yfaYjddq+DuVqeOBILOoqwW8PWXK31O5XuerfuMzizdQAgHrdxHNWz8O0t1ooIxC
fEVAISXPjhL/bdLR+oX91JbjCDwYklLnziw+Q5+bZvHV9/K0fHNXQtbT6cEkwhzm
1wCpI8htDNjwjZQUlb0X/eNWegBi3afNJuAGwCWsoSHdFEKH9m04vKQWDLYaE2bA
88BhUYy2RwW4u79F5A9UlljziMBzNsgG2IIMSOPwkk5nz5ejQFctAexVjptToQa2
0PCxasMDdWtxl7dxhIrS/JvjOT9k9g6bBMWP5XtmRijAGtfI06MPvF1DVucq6deZ
d7FMG1Qo+4IuRdvwf4KMwZkSyJFyc5e2Ycp8PsQ6ockYD1IFnAFSlEe8ZgHc/eD0
dUJbbNCsEitri1LgwCU0vgH62zKgIVDqvkS+LNzqUdNsv2cah9duz21qwSDPl/hc
yvDuDnuTXDBY58XXj/b+PNjmRutVJtXxJYgEWGMLnQ4V0Hd74AqRIYfi1bb8YesE
sntuhVJzBWvulHFxRwPsgSlFLWNKuJy25yQmLntjDggtoFowNV14UEiSsnbwZY6z
uGASF5PDwQiayotZWGekwOdJNi51G39drAhuAxO8Ujtkasaxiedi5fXqK/tka6pi
eMuenuOt6a4fQ85sKWOhLgRr0+MSCRwrmLuxmy7jfiHNuD+ZCGlHONAQoCIrPGaU
stn7tXFcbmkpvselVxuwJUaOZ03OHy78ZihDeRTdWMyEUWK0qYVlZ8Sb7u/Elq68
PtX8bz9gF+8vBftTb/Br+JCj8kzMX9u2JqZQe5zmG2BVlSpFlUkreD8D5r4TKZ6/
9J7Vy65Xm+NBiMPghANmaJApm9kQmOMr1gJ9azhBdQEVi4K66UwbRl0COJYJcnCX
XbHtoxHY0uplESkxyoYuxSUeoMKO+I6+FR2S91oE5WpIgZXZDdrVwY1wPRqyqlan
MxWKy91nWn/jj6SLKOYY0jFpOY20j3OVHzSVVlffwrIUvBqxmGEuuvxIEZwJD+lZ
x6j2CsR280dpSitOuUk6YUrlLwbesASY1Kxq3V6vGZ8XC/m2CG+78pL6Ar656t4n
a9SKhLzje2+z/42uwkXEjNxI8Kyde1vd0SkUwx/oVCuG/+yWHdGxtJZ0H8NvYPkY
yPo9BvH2e4emGEKhzfcEFB5u8vMb2t8VanFHvkVIQbYrwumJLjz/7QJCJ4aBRMiN
brbXH7tYwFClDWX7U7UF5yXm1UHrQRnD4ZGxu6SPxfhn46UlHZolMMsB6+N8h7HZ
mMpknK9z0JvI7CXmPsOt/0THXjOeoRph5KeNVWHpASOdLaptrSBNckezp23X22lH
y2dolw/gWeIR4XY/pDtyDBa3hsW6Cx4L8v9b3tot/PqHEvreXaJFxGMMQO+RIzAr
TNs6nnfik/LgvzpUHyK6e5iySSYodKcMB5DPZ4XR2m/D268FUAGYuAAg/EEvmf54
qMriwpupxcArJuMzaw/OkinRb6N+1mHq25mkGsPE56QLosm+71WvfJ6O8R9PkcSB
/waJG9ghyBH87CFt4Dn+hGOAJshKuIZniy7nRqDTpKsbApBVDwL3Hx6CQoC7zNgK
Po6Ynn+EF9Lyw+hR9FCWJjYupWTapXE9T69B6NacZoRjA+TvdaZSvI3SvtgkvKgM
KrTl52edfquIwGEiy20Gn1DPyZ/f7pJWbrPxiNylONDTL2WbwIjylni8fN3m9RdM
UQRff3ZtfsAlrA03RBg/4ryXhRfkBddM9JFeMDO9h5LappNemZu/AjOh0VUL73j5
aVbpcNcfGi9KUavYNVjyMtc1KQawRnwdAOgP810u8tnBQyRi/Y13zf/HTU3GfrM5
V35a4K3xihYwv6FhyqxWFlkAJxMBrWozk15Z9T6z+IfyKxxX7/MW5w8HCiYY/1A1
F4LW998xJOBmCjyyiBFcnVh6vKOHtkLlW4VpE5z9+blpY3YKU30+63Mhvvs71jXP
WKVOarjTWWnek6f/GN47g30LBfQZNGrZvFO8ZuyR8335W07n5L/yU1PHjqbQpkq2
GojuBs4sQBPGTUmA+OmajiruFWhmaUM5fRsQNealukfwIUDofKl4m7uJENcoqNiZ
mVeb7sVVI71dYYbZgwkhBVV0hJLZzICT3nnUaUMD1KFmmz4CAyhTUnVx28JNXnG4
ZZGZhq+xdLBI4nb6exAn166c6WPTehDIdneRiWyC9KrK36aouqDx+qa0toDmDmuA
lOCsItsJZ5OmsVpJHs6z4lvYaEG8zY5IfeG0by2z5O/8EBrwXdSCDCone5YoeXBF
5Kcc8ipaLvXvzAUKv1hTzKHLT5nqRVNEem+UyZaFQ9ho1Edi9XcZR9k70mXxniYB
eginhhMpOf+MM8jNmhrEag65RkY+sI5+uutanFoy3t5ZMo546++FHCdvDA+EDpWd
0naJdi7ysvEuUckQRURv2eBWqXIr2RFZpk6M2QL1OeVRasAopLbPk4BtI2SwQ4rX
lTRScdJ9iNvdeUcBdt8IiAxBcsaq4f1s4XyvyUCmNMX/2J9HzwBHYzTmZ0qXlimI
DTvqenaw+hN/Pn7VyCkreKNeCjVgU9KDpBmXZnR2UJvy6BjgkxWPuLWhJQDsmQEa
OOqQYXs5uMNal9Pmt5C4JvhBjbHfKmF8ohWFtoWjBZFAXMZjk9nh9ienWe3j9HdQ
sCMVs7OLv2O5EkBEArQGPxbrj4ZbmFW9svbtqDIYf0JLLQrLrJG3Na3omnwgGfiz
AKSBjX4Hq1gE4zV/CPInoZUz/Z8XTGNxsK9rnJJr7p7oIeKsQ4WkOciYbHRnS5zE
ni6MpoXnHVGLCfeW4Mj2mhKEJnA6G6LWR2isNhJQYwTKanEBfKyT+mbr+0cmg9Qe
ww27QIHRoRXtYJXZszwPoHyas3k6iG9UP5RbfWhNBY3Ka/GIVxyROHWv5h/3RbMk
q1u+6JfeFHXh5xDkLbzw/YCb47shjE/8ZcaZFV98gWXaXrAYoSQLrD6JdsjZBwoB
Nkaj3+MRtqNEAYAf1c7CrbIj+v2c6VxEzeHWX/jo+4Iwl0T4FNs6EoCBWJWhaEU3
mazg9cLZbJVlxZymIjvrdJSGAWCxey0+dWirxhlGV58ArSZRKP0PWApIS7NdfxGB
f4pvdzpl0dVCV8tM0mGWF3stz4UFJj9FsPbIVy6pVFF/9Uiydf5lfC+GK/DlkfzP
V9DZLGZLlCCFvWIiRUQ2qOQ/XuSqNTjAV1palwD2JNucjSRxKsXb/dJCMf/U9JOT
yOeWnWfj+XpHjgo+jyTKECXN4oopXkvmVbd+OK9fq8IDzwsfCDIxCpjg1PPK6oQF
N4iSSuJ1DRAIbv5XTK035lpm98Gz9kZrzoH0T8WI+VQMdHdf1pE0abE7soF9xFmx
k2CvOlasM9odh0zim/5+tkvVKFk8RaVrrYcQUlVgua+TVH2yGBbxXvJklhUzGO+K
Qj6qZuCUTF2VkHSspCkvFHdRfHqET5hSIxoxO9JSS4OJjro3ZxGNpp4mTHS3SfrL
Obv7BbykznT+OqYDX61B4z26vsdgTXVJVA2+Rq7nC877BUyfa4+f+5Qo6kWyiGup
tNJg/9BR491ctPOxGO/noTtdkz+SPvwnIiGzROXME28UBPPQ3frM32ZesN219mYg
qNZF67X88LwewJEtca2lZCSYmkLb4Z/c5ARMOgqjCRj8O88K1EQ5NRT2ZtbYUOzi
t5WWnv35xZKxLw7l/6FE8Qm/PcWmp24rN4+suIBisSMJICRwZg/5tMJ6itSg5reo
C9p783O51Q13iddsorP1mecUZTzHaiweKe0wwVvwlt3WDVQmH2UXoxWDKAUc8dpu
vbpxIXJu53Yn3NByiWGxknPTwvj70OjalcdNfPF3uKBXXl4no/jNx5kGx6GoThPn
nvQXvTC1Y8Xa2DnWXjy5MYWpHQkvPZslm7dfiImVL4JSFLrEYvokKtjG7RdHueEf
8mRB2HZYbluzLvIK0ZDaHe1EzzN8sJZlC7hR2WqLCoira4Yl2HwMswncNLhgu7Dp
o7c1i34DnCvV94kRXzwZOw2TF661vG+TU/8sj78Hac3tVOc4t7LXgD0KvNKhOQ83
2EUtpl+UZXJ+5CSGsU22PbD6gd0pOEtz0/dS9zuliIGvWx0jBe1Xf2/C2I7ceD2h
9DVvr7uB6TCuw7M9T9SzWPwwzptwn9wwTRfQlV7Lt1ZPyCwHMfJtkJEnBPBmrQDF
b2QRB2sjdkRErST1O1/VbHaenn51jhZ1Kwoi6ZcB7m7cMk3fwecudAy6agD6zNT+
nMRYk/ZH5AfooAKHexKa3CrlmrJTzOEeWFMsbejVdWiJkf1yy+b1yoTqz4uODdNd
V20xGeUVHatl2jycGp99d6hdgcWd2yjudqQJXaUvYTtQNRrjTEgacFzRE3Q6PsNB
BoKYzreO/++DtXQ9KIOXRpoA+BxFSoTggsEPBUqTzjQyEY4hrMC/eOiLU2sngNKf
zustFO3nkhhPPYNdt7xOUAmMkRVuvSmbS7bZ6EMAhyqYx/uxpw5q1KgCZtIMjFtU
`pragma protect end_protected
