// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
Hme8ub76alKiNVVLkbqbWEZ1OHQ3yesTTZJSl3l7sOWacRWGcP3mquPetqlJ2i8sBg6dMfhOLBCg
qvVRQcrBSfIWSyiNPPeTA22aHMF1t3lnPUHZPe/jrCy8DDcTUNLFQ77Yr2l8q+AId3gnvKxQvYwE
WVsGYzJPz+yG3KURQUS3+i1GKJhzLs5UiCc2nAVNbLIfzi+7dqAbqDSCTcSI9xapYByLBuXbz/1a
YCaQ8TvCX1bi7IQWqq1UKOp+io7qLQw4luKaolePOxXGVf2EZi0e3tF+GxfhrgShIZgFuiAHUVSP
QYBYSxHCGwFnDgtRtPAP7z8cdNA1/v+ACPi+Cg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 6144)
xX+Nf3ytmVPpQ+muRzjdA3N1QHKiTKi+NhYby5tZeJ4EHoWYCeyFjpfNNmONvcodyWSdaD1jJl9e
GH+RAiJWYmPknhEhh2MTfwMkARYHw1uIKopDqFE4BrxstI6vNhDYN/C03ipVptGVJvwrMlF0U+Ud
p1zeFDcBSCD6ULh00XMrknD6n6PsRlk8bCHjXM6rOg2lr74TTySChI5MRpTOLNZTXlDbptD/CIoU
82rMYClzZLYPJ+kLRU36ufFaFt61BKYBMiY3rqVJ8UEOzyLdMLln3T/wzNqhmRQNAwhDUahG7nqi
yxXBj0xBVFAZLCDBal8lsUiWUwKG8xz5tB8ZFHms6lmqOGkq7sA5JAY0ft9pd2X9PzzKArEvrEux
q87s632aFs8+dLmr0Dpet4bAsTd2/TMI1NdUVleObAlYmAxqnz8YfhiK0zFIp64NZXdQgH2udjJe
Lss335O92qEkfqYjKZE1f/WoFB20J92kzqEnP/kJ553jNwvE8sXp5qmwqj2suNuFuX/YrYAuXCSW
/QrBkTvw2LKktfwnDYbtdxmYJhWamXs2dviDPsWeBqXTVT27t6rVr73fCoe0AcDUVYkCSmPNBi6C
yi+gvmY9+OrpH9hFNP8vtYgWpMrohSkTTN1dPpN5qGHnQlcx5MhooH1jb35vvsIkOt4jAl49HugQ
xY27sbxDfGtk7VgSFqgZFNHbBCyWVqrHJKyMTwnCgdOx9A721rtLSan8CqXQztFi0++IKE1DJwiV
ICFtQPAdFlFSas56pY8DePYafUSoihGG5es1B1SoXbWlv+1gJ6fqBNzaJbRCGo9B7YlTvLrTOAYq
bFyTK9YD/xLJ1uu4bKXZQ5zmGNjSsHIb3YP4oacBSde3Atv8JPR/GrVcWoDccn/pTyMS018C6uuc
Gyz/27yJ8l0AfI5jbwGAb0Hy98lZRnYMCeNzMuTmypqfhw1GyH0yX/SwixNXq4FCRlxgLtYtdmUq
T5Fj+p4ZuzOcjV17KeToJdsuy2vxmfRr0VQ1uP6TPm5Wczwu18JqnJUNHfzhVJCmwMmdPAVrYRue
QOxHAWNvfOD/hz6tobLIx2lXMKbW5rMfzdNf/u5pXZBManGXXM+3UpOJjMbEHCgOpzcrFbEDdxLM
HAyAmhdjHQQOtPNrVgZG8wNiYC4aRSBZDk9Fh3DoeQMIhro4LTu6KJ/myh/RVhOIjkno57gr8eU+
fQDZ72/IG/jGFbnOJxYNWtHfDhLyaBbvRgZFkQ5Sgn+pMonjgKD10UfqY4D120tlGJTMs3rTmpnL
D8XdLgv32Jm0lFp7kbDjHUCNIUHSnjDFci0tZeS2XvA9OLUTclr0UIpYphVsgnGstrK9PZUMp48V
YFpI4PqrnGHbfpZNLEOvhEuZoa2wWZQU8lE2SJPtjnLeUY1Ub5HIVmAxKUvu9rJeA2gpN9vAn+5U
rXT1YP0c7o6CR1ifxyX07Q7SpEFptRov6EbqeqetnHN2VYZrdoMKOUC82uNKcYBLeHlDbevZ5GOx
xcVqbMAnXIt2IVLe6VSJWyotWfeS4F8vyOixgGTVZSCI13cwTfQgz/dPsKBIXakweQfPXav4yUty
fclqi+T/PVjccvb8O921v3fji+WjtJ9bH4J8qJlwrZkEHt9Mlr65NHrkRQ/Gh3kYXgXtBWhc0O5A
xoUO4hqImJ+zeFTvJvJk9fPFOSxDueUBQtSdkbDsW5ZAS7paHptJNRnREKsgFekbcjWZa8vbqkA1
W38j7TAQszvwazf954rLPgFYadYChLJdtunUOjcTGDb6++Kwj0SFyD6nDB1kJrGtqXVQnZ3eOKIm
eXjpyulD9Ob+qOH1TJ58rgXq+4/hnSMmz/v8/Mvpj0UqHQT60c+EFodaJPWyIoTCVgJzgm/LVH+X
NOQxCT0hOjN7HpXsk1FOieMRxFS1wiMFxBK0oMGDSc3HgyakQaODWE09hau2AbA1yJ2nv8oSa3Jc
O6iPsnqOev1zTE/Q8IW7RdPFyyM7rpTuc0xKxWl8sceCeRBU9HKo8H9RqXQyINnLzC4IAnRmcMik
m5pPjKNpMwwAhbwlY/7H0psuv57lCebeel4gVra3x8ednIQFTCszxAvYCoZT7tjSSU0RinvW20qQ
N+rDfbqaIJXZEGGjloqypQ/YiIKWwjnhVi7Q2D046JfoTXtzKDD0HyHKjse587zC6AeMYEtCA6qF
dPK+aXJDCEx+2FR0wFjCZNKNVsHX35+ZhO6efUeyoc4m8jRncgNlxEfdyY3bZu3OWffjEs5H+Wz1
x5LU6QKeyiHHZcUbFBBEpJA+ptPkCh+yYS5Xx5CRrhxqIdsvBOd3D6D48wA3lj3UKuTWxl+9C2Sj
TsGxY1yRpXViHJrRwX6y1PztNQBA1rCwdLRuMUQnsJ6LCMDaPgL1V5s7GZnjPiO0FKCrz4rhdKRW
C4rk2RZYm5q77BdGyZqEUgDAU5VSVpJlI6k4Ki8dRqnowLXzo7l4LCWHOeVmEzMRoXV3ZCi+7u0z
wgEp/XYcKFixrvGxyMdTErvg5pRN46CtSwx9a3AlZTdh+ETNm7O2AWn/1bGIWywaaRkv2DslHR/n
cQrDQ3woUvUwDefy13i+x/EtNu/3KuH22coJwN2eclnYgKOKKAkSEDrT3ztOvTsEYD9M6lW2Vk3G
Zkm859SqXFaSUafyf5slGvRtgcSpD4ebKATME1hc3ygYN3qRU3l1Foy/hrO/EGfmQyaconDCvTbB
R0isJYLGbVIO5cmqZjwgRcu40hnKFx7e7yyTrUmU3HZ1o1yqHR3M4CqddoVPzO3Bvo8xD7GdF5+E
0H7ewFazFM/ZyLeeOdiWnnq4KsCYGnYwKQrb3eyLAwe9L2+PmCS41Cvy4MJsMcTagTDYYTYdLMD2
R19rxMm/y3aRp20gsXGwhULEuU7yAAYpg3UJJGWD1kPCtOJPuI5XgH4Qb0HK2ErfOuDNpYGPhgaz
P8FbPL7GWFUg3xFDwExdegMzhyQKLVuDD8iehk3vKd79awChWe0PEkLSEacANuDCy9UFFOOxSywU
/SGveIpJFShG2IKMxm9tUxLS74CfHExzu4F6cEuGs/fhD+p38lGSD2wea7Q1eMVtuJ279zU841xL
DVGbNZrM6pR9zVlOl9w0YS+a5ScKMCm4/V+8BUfbjgRzskGPrVzyW4jIBAfNVhHP6RDt8ZyAp3B8
CGn3BD/R9AneSMonJTpGff7zx815LD8p3uBxhLE4gFaH0R8rAQvFHc8zfEGNLX8D6J+E6Ohx/sx6
9PdfZuwgdw5bVe8EaoMMWw43UU0tqnO+b2Y7c0RGoAW1dPr0REIuBSafSia2BwfhGRyHLHTAMw4u
cPuvDvKqFu5DmiOZnIBLtFHVY9AofHxudwKJTrTfJzc3wfkbSyEYk4Rnc6PBnJCRP8xb4TuDZr/C
XvO12uqMXUL+QF3wcC+gu5LKDNZfH6R+k//DkHkL7OI108HaaVM/7MxdgzkKDFnOuXG4QsgCzsNO
ixfeNwwZGBSJaC722H2vpiG21xPw8JVCYmC/7gp2ls3/P/+kQ7YKU9qIKIW5hKSDKlVYmrP0bhxU
PR7n9JrM4pNIgZde7fEzrhYMxsdVXwK/QHJgNXvMvXgZYxOYdfceUIjyWkzaBWgAFT1xDRcHoZ2o
hVDit2Recm+WIdviZi0rOgZ+pQ+zEBgYONxPRFcJdMw20hRn7PsTtHzgR5HbwwWsiCjq5iUVdGuW
lskeu3YbwsvwFWi4jNqNfct6wxglar6a05Wf1q2VPhF9kka7GWD3o8Smwj7/eIbVuUs0nU9fssd2
JVqkXCrZ86QXwxoaytLzPztGWZ/kBoE/U6TfJAweHIKQs5DLe4kfCIhimk/1bFM2KH8JY4Ngfi2m
wfpSNA30u5vVKcccztBt9yXXkqvMVq2YW8slmomiu83W8ppCgqmMP/oZIu3+d4B2Milltu4yO13u
SNC6LmaCBAnDCo8t/V6ZvKdy/JihDtkhTA7BZic+eJ8HPTAAYG4GNztpUYMle+dfDqN3xB/H35rn
1QJy3MsU1+t7wo/7hOsaQhfMACkvCPRZ6sCDZpgEm9HGlE4JbZ7EYl2nB5I+BDh7lezXp95y31Dl
KaDsmX+q4VeDMX3ycBgD3MWgijUHHKAjWLNb/NVUDpqQE8w7WCR6z3OmG/LAxhO98MIhSsLBh65B
VxstYTlFBCLljYLhIBGoCc/T+aynYZAlMZ7OlKxBhtfVUg8DXrZmPql+ITbNXOy1tZzUDSifqCNX
GeAUFBEeqsYSNqV0vkqnQ7q2CQf5SE9K3mMaKshUv7kP4Jprat2XtqrjCtUzSrnqubO+v0PTWuiR
/RRSxSznojqyiGIKHAzp3nuOjmuby27OQEyD0C7nQoXeEXTu6V5m1+Jz8ijvdcHkqnrpeBEwZ34/
W4LnhWTP+huNqBxQWdQCEGw2T6ZsFilUK9XM2UOUGp2Hh4sOq5ey0rZn8rocInj4Nt9Rl5DWpKAE
YJ3mpTWMx1EZ6GIQ9Gw4WDNNsOFvrnMdiPS0pAVBELfYHZVfGOn4qSMiTXopSnOo24QTkUX3r/SQ
5LhRhNRgkKMuiUmeITQ+xGHJvJddcgSqhFTjYVhE9xK6/Q4H1/4JoH4QFd4TrteTD3D4+XNdDYcU
HcmyCxp2ONuTG0PVbvy6uIc5oRpFmHdHT6WTXlEdhYm/1jorLKLmupOx6AVd1Trvm5wZsx17wdT8
lHRd20UKhJqR6FTYF4gnSV38dh2w5LpoRXsqTMVsWc7+QkwRbdEOl7two3LlLTGofn0z/hvvHcEo
FtF74N4+D03I60gnfXzoKefKIo09vlQfgxxFhG9wPd/ZoPcQfrGFhUpiqJb2iNvQR+7bLyGLG+ZN
6TygZq7bfI/pYU6IDKy52kNfYH07oE8qAgNsSaPWKBSR3vv7oY8SYhoZq51IQMJcRMRmOeIwO8AM
c7XgUhMMwfZhFKD93tKNxcQ0qqFt/rnvhBSOT4CJeAUly44hGQm/PyfkzuXji6IBERwwDktaoZPO
avSro7BOX8yOZPnak5X0dYKkH98xjsBdkQ+5HOe3Q92cADoLbB5uQNzkv7VrcYUwyf/UBIVt4OxA
pooxzhpKxCQpvtmuKFvhObWmAHjmx8U34Vrs0Y6IFtQgscJBusjeKAmb/TAjkcieefTlnLY7YNIT
WF5hAAeRcH8C0V9LxWdUglP2GPokf6BuJsxQwIDsgD3MxY4ns2EAhdvNs9VZzt10IzP3ZkAXr+3x
3cB3K4sP3QM4127HCklTGIbOHpQz+uJNEXuU77ri6vO1oUj6ip8TAq7h/0rANJttGTWKOwryTsUh
HlfAnReU8360rY+8UjrlIjN77cIjbN/atg0YrQGNm4RHNNNErqrTLy3OVjt0a1ur+oZnFRtwr25a
Nklvs0EvZjtg8HsW4Wambf5ZMCGPWMsQsiFdpTTGmXlwN0oYqxn6/6pnZ+GsGAJwh9JV7FZp/mg7
k6Znh+ePQBTUeVaMa7LjPCo3Kuue5ECqtPYGKuV9x6xodd2c1LiKUQN4ggCUKiq2eKle5mGXixkP
LAnqwnyOVhCDOlO0XHNemPOcXbAm0Ck+oyLXlUypfDKVrOH+SnTv+AZeoI4oKVn0L9141A8nmlBF
J+pLiv+Pnf2BlDEXDAMdxnpyq0JmgPRGG/xhiqNvBpfcvKQxHdeWvYZWMmuOE+nN+oUJm2a34VyJ
XNROSNOiY0rAN/Ap11qXzoa4WsgUKLt1E93AIyDEfoJ1dAft0kHf55Sp01OZuzyE9dht8/+OKfHb
Clu8dvE+CvkUF1oTCf3Zu9Bm5Uzy7DdTFvsz3aLO0IVpBmTFFgmYvLv2bIpP4jSzhNHF0WMNIdsI
RyS65mz1qJnrTUpqvICmG1y8J4mruYa5yTQdqsa0ysD6OJs6zUAE+TaGOTW+tjDgOAUUPUQ9AbOc
6ZqRJvhaoIdRL9DvcNPXqH6fpTBi8uiyMlKhmeurv5u65U28mJknOND0KMMbhgg74JRaDsVLI5Eu
ZXpCiJgfW2pu2NOk1sV8Z+IQi0QRkCxpOkRNHsHoNvS5tJn30iqSTYJ4jr0tBJc95f4NnoXYpXn3
WAn3CLnwuFJd3SDRShGvrCI47DEiLB3jIYEaVqWoKVSGb9zYzfv4MMJkiSQV/TLlcN1wQKDgbOIW
LqgmpP41xKFF5+9zxmOE/INFNGHg9uR2sdMhTkNA+bg8yN8vubyp4JQNtnERbYywKaJVC3pPqqGg
Ju4mOgnboDiO0x5mNav1XWTbKIxr6z6uBCCuRYrZl+e88imSLGfB4WYc4YspEexh/82V2s0o7oAv
w6qWxOM8RSxmgf0pmRy5GKoUliCQbMlIyMLi18izvMHDXVIQ2fFKJylte1zSLUUAqg6tO6L4UKoF
s/8mjEHolrOug/M+lPXu0V1uPa7uEoV+vZt4RHsZjHnmj7wkRjXMirQ/7duOBIC0YUF5Kl0LGY4I
N3Z2yEtgfSjqoEGMJPFA7lL7kOBwodVF2qVi9tMgdtYHw0oJ5YwXPWOFY0EJ23r0LYTssSrtS7wN
EKRNaJOnw2zEi6BG6xb+iKxv17PYpLmnBdzsmYf5tDbKn4JoNVfSTRS3O2NUYQdY9BxvXzRQfjNI
c6AITzrQSwkeCKUkY51q8SHVHpyoGn+BjhfEfee0O+GcJFn8HgqFUDElC1xGe0cI8d04eU3ggkEq
f7/yQB+KS8blt0S6kxVpUz6gDeyj5Y0WWRKfoH0kTqXgsynrK032nGbPuTAdt3p4iFUfDfg0sdva
NDdt5urE7D1eAo/Z9P7gvwJejFUrAQhKq3HDj95kENxRGS74+m4Py36YaEN5JmaSFY4SWwAI6SCY
vKFKYIIxw5yEluEr8fXGWtaDlpA0vjmwYS+BnkJy5OGpIAbjYZjTgdofkeObWJydmx7F5u1H9fdx
O7ZsVMmH5sydYtxkJZW/2KQaofUqsR7rsTn2ydirr8HcBfeo8iC737NxflSUcuxXX2oyADLrVEwN
11I2gJ9h60CeH0pk2hx6MzFJN1REdOS/QpK8eurg6u6BKbX1YaN/mEGv43c+WmOGy+EGZ+SruNp0
SQhLLDhIELPRlsZCDdmnvDpmHxwjLv2GrQVNRUENY/au8L3tc46AzoJ3thZq8dAwdjj+FXMmgv0N
n27PoiyUHV+GUTLSFoQJhx/q3dcBLZba+EpZqGGN2IvzfjJKMV+7UewsEHAirqw9vBZCYvlsNKI5
kyZ2oa6SMVotyen2dnarnzFvUqrR3mW2FVjaQcVm3LPjFBvhUWJxrLnGCJMH0mSIwACHdH/YfteC
YHxBKWvUUPIL1tRnPFIchX+C6W3BpQtfMqZNf2PCJWVIelOzFdEpyimtIOSbeLqnsKL0p+pnF7jv
QBOMwEzXfE1qRv0PRESsSe/uzC/VkYuG1qFdtW9WYdBlDMsH0sd8/WDQpZQXzXLVQZ50Vey3eK4E
UiYQ1cOEYw/9+jtAf/cCjXX8Vel9QwLMZmiwdRcIW44okh0FkJixn7ylf4zTFxqDdqC4ZkKhW555
n56cKQo8zB51+tJoCoJw5e2YKLXPQkNMYcT5SrJwPG7JwIeJ8JrMMnIZvaAz/8+N6/ThEPLGWeuF
Bi70/XJCW1/uEM2nnlczW3UzYpn2uK1hYN7nh1H0uLCsGq554eUY/YarTRF+u8IEpv6YWfjLqpqa
xEHyeGd8O3gT0UGTqWMskZWIFUZ4XwT8Rr+u+Nf/t+ZG961hJpgweBhYoz5KYyd9BWymojFxqYLu
wEc65Qlz6vVZi5dr+RgVrqTymTGFmcEAlJQlwcUTO0IHp3etBVVUCcSYcMkN7euS9MPNpDxeyJP2
Yj/d6v3Haw1oRIl0cA8j1TGKYnFKpjoqh3B6sF3xnssC6PmKpqKT2vmUO4hByL80tbOucOjDUCKe
Vz0NWJXpnhkeF1Y+4dTK6fw5d4BRTvHt01B5Z0KSdd6HbPUjEBVvkSUcV3Ztt9lZ4JI3yr6rhQPg
Ri1VogJ4URyRdjnO3o9pBecI+I1h/1poAzJ30jT97JnrjR2/dRFk0GiqYkv5DwldgHSv2+4FO6t0
NGesebxzvg9XqDCed3sITgEGAV2MA6M54k1S8cTSLR0WFy1fFOORbBZkRX49mVg2RKP5V7OzIIZS
V6DeaAnppLSnoCu1JDvFS4o3SvOB925/bQlAZEh88MAB9S6ydjZ2iGzlx1pz
`pragma protect end_protected
