// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
iHXiOnjeB2+/fgJdG2j/skUmy0N552oZFc34exBQuj04SI0TDRCIVFGHLnzgBi3j
ahGzoLx7THcvje1lKvhsflxfLGhR7uBuMUYzSqVK6P9LpswOdSBnmvmrs1ek7M1o
baEPSffN6SPt3i7drhnlVtkFY2R5UNoPF3dGPjRxmTB17gmaZel+7Q==
//pragma protect end_key_block
//pragma protect digest_block
F9c/E5nkIZjHHc2HEIrdjQo8e30=
//pragma protect end_digest_block
//pragma protect data_block
Xx7Ng7jjoPwvZDZWdkutF+FxbljBKGQuKPvPWK41CtXMBpeJUZDofoAwFHEiWfzp
sPC227fvwpcxFgNfA94JJubmkJ+2e674V5hN7y3goIC/mZxCLGIo3dxPNXbL8XFn
/tJPN2sE21S1jbQb+tgb9SIxOW4GKzWAtf1x+grI345ebGzTLFyJiQoC61YeLNe2
Oc06ld/Ks6j8xkuYU/+E2krF1aCUlbP7Vtxg9b+CrbxGCmY92g/Iw35fvbTnXEkL
8Y0b/Q8SH+FG7jYiVKza421oj+Tm93p8H8MvE2cX/05CGWby0FJNmuBtyUMJ7T0C
yxEiC2l6DVaVLNdAKSajCMak9XgMVFOcQTg8MdchGHqYS/XfEatijfoBzWF4WEUo
39njU3VATGIDNSnH9y/XHB/kozCqy0Dp+74WIgf1OWD2qSDBR8i4TYjkmMWfgbZo
cGZ0NWSK77dmq8SBpCIUlAqxCSyxn5dLh8GwjAruXnAL3BaZvrqy8ap2CVqaVmWj
ojkCwWfu58KcAXItn3tr9iNQ8lKkD/kE8g2WLSg4Xu/DoO6fZ1Gfu6TZgKVx02Jt
YjEYa61R4C2yVIP5smnexS/DsNP6icw29vAA/I/6Xf2x5FY1CO+5hZuyQ4KBP9F3
7JbUdJ+L03onjvkPi2yYM7EcPB6FzcyA/D+JBMeZa2muEY1nVew7YZe3/6C3erdY
iC5SMMbYB8KNYgyGjCv8TSfKbbCAAdJ82xfwvbcHzapMG5CcpwcTc9RnS+8MfXbM
ckpcCL7M71t04x4HbRyzkqa9k2/YN5nv5v6v91X6priv3XfApiMK/nEs+Vg6aHqR
jONuztwObezzCmCFxzfndaJXB1ezYlzXUajIO8Sm7WZsXJfQ7XiR3Fe53kl8MiZV
JnVzrh/R5CuKs/IiJn1w/spDvE3xjXFyd0QxIyRdip3NZVDiFzhKEEXjsioBF3Vm
42MLfdk9k8etuS5g27jB4Z0o/jLMhtsIaLbbb0ols+uGCbfumcCC3EvBv1qyOnwn
D5U3dE0E/x1zzbuJ8VN2RFoc7Ss8LIw2Fubkk+zaYlCfMwYrKz3MZLqShQrE3EuA
vIMfgCKf5pciNLvK6ksU+iwpK+AIJFQC5K3dnglyU+deRKlLPX9tVlv+IkQuNaWt
BdxlX9Cl/NqGMW6FDerc1HfIDAQ27vZSiNmykYxoVNNoN4d7WA2ofD7hL7h3CIJB
H+eg4x4ca04jGhsYx6cJezY0Cbdykv3lfDcnAu6dx/mHiZGw/T4UiH12M3HH0KS8
AR4BAgnMu215zRDscpAsSKjbkpa3rgBlFbiuJMlGI/20QOW7+7e5WcHeH6eieR5s
V4gA6ITTjzUIEPRYOvI6GHtpoYdGPKy924WjzOLkM/fRhW/3X0+JHkEFwEcvoU8K
xj6wAau0Ls/xqngpxBg6e78fR+DTt2i9voYr9fd9WmWvf747SXfsDuQlDFMNsE0U
CIkjYlXCm+mpNnn6KjyjJv1vyPRfan2waIpxtBpVxaycuF34P7jyB3BDt8gatFmk
ga+GDpjJqOXhF6JM8g+bIu3RLyedlsn9V2hKmJ3dZty2Fv12XBt2JvaipC1IE4U6
tJD1BuDDAvHRGujZSL7DEF8TAQsOF/Q/O2p4b6bIqfwW4tB2h8jFdCk04B9OLl0v
X3PBLCaAoPrY4WMqSj+7LDQ1Qco4lnjTurLlnO2SoV0A28A2YhJLbQ+tomu4m8jF
7TRbo3JIvpgM7O626W9mdpNo4cjoiWq/56xXNsuXsVklvEetj/3VeUhrwy6rXO4c
meChAJAGw2ftug3W/PV+X8CgG7HkZWowFKUYOkeGFDvmgsb2i4ZM2JFd6UEq3hhI
7o6GqeNcMpDmxo2M1RIaX5ZjFqzWepgOi8TkYjShGZxMs6tfqN+Tc+Kw27WXPQZ6
vidSAQF3dJfUWPWqk+Zd1mfIf7aChzW0fo6djb5LOS1hQZSQd554RkY3HQBycSHZ
GTr6+APfAUKqlOBGDZthCEFibIs6ycNLAPQ79sVh4TSa3cuB2rgrPMBQmN4T77dK
zmSskQXedWwI0brtDMsXM2jKd9QX6q6crbdZ1l5Q7xgxqwVAmQ/AIWG7YNxNxtOm
prCGX0riLwqGkF0kpCxOr5SbcGcWUzlpvYieH+ztw8FQ5LgJ/Pmp6tJwVi+2Ebdo
/wyU5IGREOCq4wCAczSu9KPESpWMvEcAjZiDOhicuVQ+MEvezk5Vn2KG5+PTBjlr
VKF0mGfikXEplaJHf1jiCjRJycOzYntLTYpKDkh7sDG+EdssnqgJIVUxbwe7Oeih
ZM3X4ggZUR2V2rNUEl0FSWmdW16GQmfPZotavaOWJUT5GXEE08eURGHs5Xc3hxrl
koVuUCZi/gTQFLh0AD1fWLEP7clZBC2o1Aorjj5MuXT54sUqvD/63FQEnaCDl3fk
znLVm2m9bYxEJkQ7hasw1hNPzPOMT6SRkui3Z5/y8d7K5eN9kSYnkZtI1iY0/7YV
BYeykNm2aoa5psr8Yi4EE5mkS8MkQitcoKO5ULVdKgTxChKINKQtqgk/FTIdYNX9
WsgN2f6FX0OpHHzwCP8qlkHybJ0vXX5BEpaTZ+q4UXATzUJr/TaQHp7cstIRbvia
rfmb4Png4Iue+Z/IcaYv3nWcCH2ve6/OpxANPkPenKGN1sY3gkqX2ejpVvvkU8vc
U7U2ixGqrf+H27sgdFbRxjE2ZltSjwtpgB9rGjqok82w9SDTsewfETSuoBH8tzTb
SvO0xGec478P/ny+DuLp9urv5lr03McBsybwVUEUcm62dhw1z0uTtuzED2bCf+dV
yLDK+AjIc2xcgz5kBt1qL8QMSpN2OKAKUP/3byKgDjRtUQUNy8Hm6KBo96iH9B6b
om3Mdspj0vASFZrydndeNBVZGMqKvMAvCRMhmcu59QykRnbAH1qJe9fzUHDGJCS3
ZN8BrRqYVULqIL/LooQlT2nyaLMumUCAr1KjpWIKfsvCqHrqb1PmuutOrW1d3HdF
34i1DOK+b3tMGSixxIOpJZ+/+nok17GsAlP9YI2l9VytCdOdrVIZUxOiK1mfbnWP
KYgSwZaj9jmKT6iUXn44pl/0eROFOGsfkSI8PS+Efu6EiBoKmTP11IpsfOktnKpt
Qx9gUvbqWmw1fGPhYkRgzrQSQtj6LaXP2ggNqJVslb0wc4oIvUCVvDxW6BYnKjAS
2DCqqx4bNEB8ykH2EYotsilh1+1A/lhaJuaYmTdDJgn80qLewEnePlhOUdVlgLRc
3GRSLPqqFRgwDLK8iN9Vy7nyGRo0c6CsOPiu/033xV4srerzm53u+MymhvfQ5X10
OQblXN9f12yyjPZ02D9oF0hgkWsnmpxdYKJnlHL4HyzacReYgQfMOJIopxME823a
pLLWQK0m0OVk1gH2GShQ6YQu3RYwyyISUl+PA9lfb4HWo+y459K1IUUySpaD3msc
gVWwzDIbKpZ4vA4mrc8HvyDUjIb4A5AZNj+zdPrReAPEo/AZJ7HsRAWA7TbYSO/L
d5jq6AvgQvPr8+te/cOwIu+q9O8xFaYycxRInrFLjUBlUdBvu3MMj/ZaJCWI+Ixf
pCyb4uBOKPxKp+k5UHgF0HKGgUMNhps7nLDc+qNaL2dwOlE3OpOh4GpFv0mfiCbM
3KI24biZzPgg/AFCwxPB20qsKepZ8nxv+cqkbEjICAkwJMGFX5Hf8akpvYPymxov
7dqyceAeIoAhmrVtShU+QkkWQsU1hhWl98Usf14BBA+2kKazjP1aREYmnCJ3gUV5
4bCf3eW3o5uZg/0NAGmyi4aRI94HWB2537cg8cdw978LgScxJtmUZclE4xj0U002
1cQy5sXZ+3twPqLQ6ZbgFx0d1mKtFj/qLpF3JIAfydMbJeQhUeZ1PCfNm29BZARo
FmJNGSilak/tJ+0J9Gu4DtyU+OCGZN5zgA52GizRhINMGZn8z0bQTZy+VzH95m5F
pZw36qCroITaZx4gXHRX4aVt89CzeJXI5AtpvRLtdbNLNz6gpspUv3MBo2KrJuE5
R08/81tbJyUow2/2DlId1xgyG3+MybVSIcHOQkmoSMrQVVek9V7EPUUJ/qndo4Uj
siYfk9eXPUGiF/aKnUWtzo6CqsbejiS5y9BeiD4BOhNKCO5CStBOqOVWOom8LhB4
oHViPLIIUIWC6EohFw5ozlm/B2bj4gJnWXny5+tJW7+c383b8DpLKSXL9/uI2mFl
esKjHrzMM0czN86T+psZ4naLOfdsGfmykJimKBzmLVcwB4IT1OPoM1nrgy/z69mu
YDpRH+sLhDyps/tME1PFmcIqBzy/RzkOTnr2VkoPGYk+mhdTN2Qmey3tEmmhK42Z
FnI8mXNJfsjlABazTcxTPFYbSLEa3fgVbQNhksY+ZNr/O6yJWBdKkm+c7otQQMEO
aO2FnB9zX2YLWr7lw1717VpTiuHlFSne1ubOKo1gAjEOIJS80oLuyhzJFLHahEKa
KPwMSqTSLzMC+9kt8SOTGnFqbfGaXEnrmRuTQpWJe+qCW1crKpFYnKNo8kIy3oZ4
CT9DbWCPe2zCu1sZ9CVHTTM1p8vYOfEF2O0OS0JfHyKLxm1tEbB2lDlsmqLd9LCz
F1NTgyjgNM/Sz9q4M4wF/djUzUifi4RvlSZ7EFh2CGZgL3UK8KNy76tWR6eHO1z+
xQRy8utbpvh2UXr39eDbnoaZtXaXayRd1ObPc9AnFdpGXr61H4rvsuny0wQaNrQa
p8Sgon/ouYY5IpJqDHeF0Q+hHY2bFnxdnQofYo0p6QrV4b5lT6U0T+1t8rqREWRR
uvhkHowvKFNZjn3xdzpOd8y3HAe8bWKUKQqaBUM3f41yBza7lsI4avB05jKJeH8q
2X6o3s5IXcDPmbsPBsMNgC5Cbqbjt04mtPZxHAwQ0+AdZWMrl6Mli588N2TA1qzz
KkghNNHC6qKBMzZn2gCtrFBs0pTgdEjafyxBALNIvOAs3nPuceWlBxosHSeQP1z+
wyGOT6XeekAK5VEHnZ92i/+vEhqxxcxgBIY9SOo4Lm11wf3f5ZveGD2zs69Azf/L
ihltioSX8gFPVeYY91uaxFXPEf2pFMJlj0rdgH/kjGU6gNlGqCJC9k/2UIT7zBf4
JHVIAvitIr4MnVjbWjVmlcOVo+8+3Fj/nKk3LvYnk0t33tXTfV4qPxvJ8NcqlDoU
CrhwkvhsZbdYgGp+sGxZ8LfXLBmU3QMZU15KDi9wFPuN32Fh2Cm1Vaa/Kmt5R/bJ
AS4VFy0BVKO4ZeSkwrpouyoi5618Z69jLi83r1NiqBn+N2WnuAVW26atGMDTtpEi
ahHBqVblXNymF5EKgcBv00QhrCwLZg5zYOPpkCAkCmx+S3InRLsI4yNTJe0THKyw
M9puo73/Ysz4To837TQWFpHKVEXkwpCrDVo6G3mZ4RmUsAcNnPXVYGD1qRQwdYYK
eRx6cUx+0FgqebYNW52lIIwP/duqODU02FiUjq3N22JL1/jMIYa1J9e+lqHgQ6MP
P6/bNaa5OmAmc1JLcdvi+0zuvcBEv6xHo96mK4g0zLg9iHx9UCgiVC8/o03KLRq5
AX4OGCSZFi/PuWnEWrBm5JXrXcslmzkQ6PTqNbtOn7ZIDjWQ5MV1B5PbXjNlls8v
5LdJ15hznvfU/rIG20CshMlQQMS1KDFQZIJ4K6M5zrl/E439/+WW60CKHU9/Lz9t
XPiFHU2BYWnsrN+dUTKOwOJZo1iwpuqPBT5AOUu03aiZ1nGHWga1zwflFtKSKSdY
0Y3l7fTYk/8VAHzK678FWxOh42LGAkceb8W4lCCYnZXBLJ52frpVgw/fPm3VNrBh
UrkEU+p/FXqGxXbJ+iEC7gcRIf4EG9GkhdWoX7Ebvhs8pYHfRbb3Z07U/sKFnlnz
JR+SuCzvYC55A9EeKX4tqWwHF0kfSQbythzufX4XGYBGqb1eiDUE6MYMJcHOXYxA
ou+zCRxjPKzuRPoFHMLAJD/0ezaoaSsAUZX8ks7zSv+IgKoxzrxJ1NZm1iEi0ksM
tgCx1VS1jYM2kvJQSGZULezSYEdlosEYqTPaPVBUdQmWwViy0iy/9UwGpPIGWjje
PK2nkjYZPKnaXMScyodz0BruVazxhe7XRn/oYOttJdnLwY+Usj/BBr9+pP+pRARr
Wkaijc/v1SDaRMn4qUIr9ZDhE01SiFgCNXyt6jJ2iiBImkOu0PPq/66Yy6FWRK+5
Rpkcqx4Yvy9o0gS3HrGAKuEda7X2m4Ja27zd2BCuUAYrw9C+bJlxA9jT7Rrdm/7Q
5F2xqjoxvXIvU82unOktY+vFkioJ8iQ1Tyt4jz/pvckC5BySOwR9R/oggKKsgyL+
coefQ4d+cmhFxmGek8mmGqfaZSVtWFjdTuz7VY9RRFaDvSPwBZ2W0w4ZVpA5j2Da
mzNAT2ydUaJreTwiNnhZ9Yr3m53aGMc1NaIvhDq20gdkbl01dbqOrsfvGnIvCpgk
7osUpBDo+22Z8QXZvu13haeFK+u+Jl93BUoTEk/WXam01nHqvoPo/K1VtsVngMT0
Qpd6paphh6Ue/1rkuYZH1oISu6kNaXnPN/mqPUVULDu0s1co74NRnYdLCHBsgY1+
eOYVmDcJahcKDO2+0geXjyOrACsk3Q4wtCxDE4truq2W+SN2FGcVvPupD2gYDKpp
YjOo7gXJ0qV8Mtu/FhX7CsgiKhJ1zyhPdXtHxjoOyczWW9pQXIiZLMvWUZ3d3HrD
8WgjJiBSL6ZB/uzX2Safc3ZQgKviqOwpxZwVKH4RYZvqvFrTHdhbiN9grI8avF0n
UF2bEogspUj2vMDrijh37VmCxOHXGT4xCAFF4LjzEOjO0Gs1wN7btO689birZexU
U3BS70eCc8hdwJhVFVU0FZt8mqUvSVl80nGhVyFDlYMejrNJ6LCBdWSUFJVoFrt0
BS65iv3hMGyFejcUDlLJVbMN/iUDdD7aiWlU38627vKYZ7zRrDTEDzgMom6B1tQJ
OE8tn/QQl6WDKXdp8BuvURBazvudCx8TSvYRTIhf/pyXxMBCAftMErPxUtfFSNcl
lwpP4eq9wroWwjcy1aAsWuD+akA4Kib7Wp3+GALOeCY29z1WbSK2K9NahXjguI8u
WYhexeEsxzWEVwXehst4E8QSW9JUbLMRI+tqk5wg/YHWbhoGjeIZ07lznms4qFFa
LJWI7+97BHGWxPxbqL2UAL4M4xPBIzvn+mjlXLp+FFbXJRI+o8fam1e8jkdPaXnM
jJge7r1JjSd64imFoEDtn3uJl/s2gs8O9fUsZ4n0oxp+3LkaGjrTOO9Dr2LUOQ56
wdtFmwKVyw8RygKr2fDPzcMGsjnAxz2Fz7QGI4iU+kc05e6EUeg6qN0X0HYOGOj+
19++qw2WM17MLL0JnvAuNR+eOdDQiu/wdkds2cYqQUCia0h3Hl5b9QDjIn619mN+
tBEOuuWHs4/h5L86SElnEtZlSGrKKbdfG8l3yZfpSwCLp46s0gA4Uqe87zng3RX+
yCeOc4vgFgLTBOXV3+Kc5JW6xoli3DXsxAPn1iknjAvFp2vT5WG6u5vaykxND1Qu
kEVZzNJoHcJGPUfIyrCpWgby9SsVVXkKAFBYdZ1DZ4Ey+x/ALlSMa3p07hKcZBhi
wY5MalVMmiEBE2kKfxXAmxJTuVeoRI3kxbwTLn+4nors4OHoy/Z/zV6NwXRL/n9t
3LiRTt89h1iYTjU7QwVIeHg9RmjLBGlDT9uSVPs9ca/z7DkNYg9UIe7Q3ijpOvEW
vof9e0qXn7/sVLGSnMypLYIfMXRP0USlUHMGClWOHE4eOmkSN5k06LS9wF3GKaPX
eBc67lVJ1Drohr44svtI7/qScehQANMR25VpU3F42CQPtgIVsKqGX1HWhMy2/QDL
tpsj0NJSzvglaYJ2pcrb6ToNaxpHUhzTZPEPAaN7z8vrFxf87D2jVXh9FeMTMOgL
scgIyQThGSYAMXIp+UIanFTAgJVOYqrWzlHSf4rzykIO9y488KiIOKh+yE33TucI
Xuu7s6kxY6FXwQrR3F9O6jj2wcLFyaB2Z6IBB5HJEdUqpPGr4MtA7vcuIE8E/feM
MvCaRBy1BfA1N7zzyLbmycY1U+tUFvEOCs3iasePDuVRHOXEQjV9LaVqbfFZ8rOg
3l2pIWvKho5p/3qaEs+JGG1laxbmQzI788FJV6PmjZt5kjCrBn53o8Q3RdlHoSPJ
g0WB9Z+MCfJLLgSW61NfX3mjGlQfMt7N7AjSZKlZnNS6KIszHWgKLXmLYCduZRXu
CtdGckDxPjx4HkIDbtigcyb3sJpvF+6qAMnSi/bgkFV2JpDX6esEEsnrQ2Yqd6GF
pd6Z46/Ay1jR/5OwFrrZL3/ynIB0hTFBzCkqVccEoirPBiLWT5FsEtdz92cG5lNe
c9EKjPU2szLIR9/IhIKM9daruFKf14bI6mUqyAWUhqW+PUqdgMa0CLMwC/bS0lfd
62jAeZggpt9IxbmGCZ/vYY4PmshFcdeGuCWTT3K0Rwvboat/ypiPRynm2TP/w/8/
/kDjfWDQltSJkF3SaNx1gcu+o58F+rGu/b8eUErP2FTp7Ma/6Chak/0h2qfydfs1
+IuXxnsV/m/9x/bbQ4W3p2ziPIvmEogQCZ0Ht1c3Y+LrSw8lvROGCuUjqSRzf/wR
qNMMGXB/uGKf3XRCmnCIg0gnce4WsFgwUMGeD+Y/xmqy5bdimaxCIE3H3iEHPDig
PecnoNkgBH2eNF6svRoFVdZbjntIck43seTugojxYkI5WnmEfYpr8FRyqaUAwWQ+
YQk+evExK/f9/AV+ewMwDtxF1Do3NyBpLjjRcItptKuVgSzgFLw6QROzv1rK/7Ac
2F7amurtiq79VuY6OOzzQMXTMEJMHj8wga9BiCcsHKjoWr2RWjGznYQUmaIUxPIT
0D96uTXGgZnLAKk3EoAURvK5rlW9/15VE2eaKhVrV0c04001MnzrtvlSuBWEQoIP
TE32vvY5yA3iiV2hUUolKS+JkLdtYSTaFwIgS2JKZbtvU6c36VqP/mcsJYTvXVgj
RcZ2WDKI5Yv1Td2bqP14wVDIskX5Os3BEhwzNdLV0er8Cw7jnoHTTsApZoYfGmR5
CyNDRu1XGCC9PVC7ZwroqUOT0YQwmBQar3JLfdxdcCIns16MpJ6n/BMxR314qji/
sC5gB35b7tLRnU0fjCevTR6AE0Dy3OaPWR5TVWVL5byebAbzELNPThO/tj8Dy63g
zLSnv4fOXM0deU/eFbCkLgnVzZkti/+xDfjpJp/KMZUICSOoqMjZ/y2I+VSkXsBO
eVDHCzjxfwCRzjlDanPe6pU2zfy9nmccmfpFyEJWVvZuUR1E5q7BDqq76l5xuiCI
Pivi9lELd87eeQIeFPLE/v7cok3SqHdLYLbwSvNi12qCR33+StuDLY9ZkLVsR/ae
bB5R0EBN2utI5xTm9SazP4QTPTJWEuSXlaTELbGVV3seH2R0fJU5H1KDOuOnOjbr
iX4PfCUpjAKp5blsdY5Jk/ubkZMsh5mcX9pX+G0HhEIi/2QOhrqQCygpQtR3QvZ/
muBYyZFPvb97dDy0TFPLQJvv41GSPi+wDthvg8pnYCSpwtlWfn0Hub0TceScGB5U
mDXnqyEZie9Cp0lcn7fTMQNcm5G8c/x4U8gH+YV8ik/d9WYruZTbs/DPLQsSDGrg
SwSgsmozVaLq7hJXbEAyOPVmJoKgkNpiYZCeKi/50toDctWno61o1EyJK8S95uyS
sixmlAMK6XPuIDxPjL80ThYk6lYF0rot/RY+mlE2fWnkB8L5u0AhAkgq3HJ+Y59X
rce14gX1//DxpT1AyKh/naOUS2e4v7T37bL0oyNjr64bqTXswtRzDcuhpIAaBLyd
R06r2xIy1E8Dx8xLh4k8I5G9VXsI5orASblSvXp79dZaktazKeZWlZ1XX/gCQ2kz
s1i8RbeRXnVGDngB+oQxkrtSo0OnuPPynrnrMhjN5Tcpl3bN/YWk5+y8IASCmjE8
O6Cg9qklXiTK50P/sUTmq4EClxpioB0mVdBLWQCZ5OsTnSpOXq2+1kks0Ck9KuqR
7sGrMDm4i842LknUwjGQVg9Q4HKg8svsx/Nmi6rHYS0Y5MW4PfP3IrgT9AGaTQsp
v3lb8zsNmyx5bSp/VLLrkoCV3oJGBR/3DHSklF+afjDLlBfVOEkxlLCY8ofriu5m
HShCvAwQlns+a7YRaHwDmuXyV2VnCTBHRRJP5LPyMycLEh8KD2uhl9Bla8XkhdDN
RhHGL3X+HhBNmQ0oyeiPCYRVszMijjOhLKyftM9l1IlRefr4Hzt4usKtXPCOA8Mc
9CjEBLdf4n9a8LtgaODlrvqw8k18VrX019KDlN/zn40dvS8wwqbFClC0QiVtDw9r
2l7ajLXq++VotSHJs0O4VugeoUTpzFzdSUQ2Eb3K+i5r2P54bcpBEFMNhFoaClwS
9oBU8ddL+VEwXAnV+mSASfXMflR2Ln6FdJtfUqQ9kyRWkJlbvCAnwq0AkJZTeInh
9VHF9ZQKvUilwpRPDe6OP+lplNcoJwN+FXMljmJp2BtyydRIZVueiZNzJs6CiU2T
5Sn7GbyD0gPZjxL2GR6/3TlcuLheVdLCB8O9hYqPLvbz+ES/nH4l/Lu1+nl8oRLc
i4yBCeJxUHhDdc4+mjO+M+ohOc9sKNqg9zDnR3CnK72qdhuADs0Eo11HyyA9PsDo
vhFshQV0JBlJ12Q+jCXmNAEpTaBBnmkg5bc8xBSjxtLXVfvZDkq+H/sVd6av5ue/
H123HfNH9clVk3I4jaRWfj/sxlqhyU6g5Gx7MmMUvl1EL/Ck0IEM90cVsgvW84Y3
MESVw2WMtQavBiUXJAh7cv7xzEk5msPq93rv+JsHZWejeHEbi1fNVxDods+GeSJH
j6B3bKL6oM/3JxRAs6LC2/72LOJlURzV3BDKqt8BMdT4WCywN4M97byaKTmQg1p5
prKj7xxpgodj0iP+pVY1cuzp0XUKvJNc1St/KPx0GDnK5uM5tHsdKMjh0bUu3I/n
DStKROU8PkbS25Nlu3GG7YGwVlEe0quv12cG2IXUmifXWRWuBlV3FDA9+bi3XpEn
mW5Ck7U4tymIhKGavjNmhF6gPCnGP/tinQI9eTE3hQjaqnG6dNrqSaY1V1HLUrLC
ccUqWpf75p6Tm8Q8PdqPYJTMMUXZJCb897nTmNhS46ZuN8XSfWtADRIXxLAFf02T
s3CXlfdhhJPidsSISPRHRHl/1d4nBrJVkh2EHW5kzo3NNuNb/4KuLTkiulobpuuf
tX788bOQZoby4FxEgbPvlj3lgOtZyGOduR2cloF2dfZtqrj89sDoKKqRQYYnoodp
OZDtA0CB5LRB1TBuKEAM0h57GdmcY6tGmwfuLJjQZuqXLuAq0epbjVr78/hT+Lr2
kfej81hjFkEVw1ojNVzRr9rl8Uq+bBR/xahsKMUQxkDmB8+5C1LuZkQY0hxJ4fJ9
tM6IW11tvug6JOWTBNplvX3Xrqf3GM9N57uPL2dhnJqKSMKVlRSziTmyYRlA5JXA
H+URxZnYkFddCOUqbmrI4AJVW5vrXlTT/lagbZKD7yG4aqrQ9gy/ksYj5a0/Gnbv
Z3St7aYTj2bRwUbz8DSQltoUIhAG1sO0xOXxjV75XhY7FvycAxd+BuLTRnCnkJ1Q
SNR/cdFNQR3ayB6COUWgpxiKnyaudFlnolLxTuLCi90=
//pragma protect end_data_block
//pragma protect digest_block
jb8X0lcG/zZ5KjoKh/mmlxrM72g=
//pragma protect end_digest_block
//pragma protect end_protected
