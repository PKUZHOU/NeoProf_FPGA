// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
VMVxYn6hZflrfJs1wKbNTFLihe/6TRFcoOcQKWYZj/kvRZJMCXFJTnoIC3Mov42x
3kLERmoAoBp2MqH4JXvbOgvj7XrICsG6xfnge43yk8eT+DZTBGr4Qet+QWHS4Pqe
bLSrGF74lR4EFnYfXa0yavrX78RyeOox53uul3QjTNDhP7ynGmgxyA==
//pragma protect end_key_block
//pragma protect digest_block
/NT0WwXDatRFBXInbKd3rFose0c=
//pragma protect end_digest_block
//pragma protect data_block
YgBsOvUBBNbeGC8jHl/f1ElIjOLCp8w/BqP3gcYZuT13ux6ybmAuyUs73LXGlX2s
ARha5HX+JorwFTKOenEn0jADYSc3by6nMAi9UN3ZwlvD9KGZYWmBp3pVtqSVGcp8
5ZP8Vh0RvIJhJOAZ2MrekA3G7e/5tkDzr2tFJyQ5nLy/BsyIWO3408aqyg6dl7AR
IgG0uIJF/i2mcKh0NVYRI6UgIrEKXZ9XjMOyUK4FHlbUscbrW+HxguWkiEclgtDr
4yIelX9oI4NY/JqBE6EGpReq78ftW8vzFMyqYcLfrDHtxv2N9S90RL1Iy84om3jL
CVcQ7wXFWx8gWNNMhZdBspmhJdrfD3zXN+Hz02Q3G+84B+NFTJeVq0+7WeHIIlao
9zhehnzs6U6SDEpIMaoOz3muDtRiHDH/3BgCT7MeMz2DpX33oiTdSi7hSrQ5THi3
EZEnKXJKfx90TO+8ea45z/d/FZkkFtJBlsEOFpCQ4uKIPH6HR6tvJJ5eAQ85WLzb
9fiUeiORMgtNSBqp2P4m3oueKdtGw5veYohTnayJZvdBpub0Dt60MBE2eDbEdteN
RuT+EXRxjK9NbBa1d6O1Z4iLzgy0wpyZznHL299seqQiZJvDnTyjOUs0sxrNw2Bo
ZdzLBLZCwCed0YG/+aNKk1DwP1uubIzxeH3KasfwYW2fLKwYAmPQKzAcNHr6nZYi
exMdMQtDCFTW5ooNa77hGtoaMcLUINSMjireZhQYdCsgBxuRFMoXHGwZxYLq3o/M
Rv2UZNVuOOT6u/GuyuPQdBRI+2RN0ZptGYyZIfQRnt6TsOwn/aFrRdPsuPfQJatf
JgwHUCQdZkZIVCkagOX6ZCBTtHaeTeKfRnJHv7/yUWmS0ixY5e9LCY7SlkZh6HwJ
TW11qeXYkf1amkZSsWgxkb2mFMs0UoukM13d95Cxdi1nxzgM0PeLBZ7CcyUhWVgX
IiVpL+/swuOO6Miiw3jH0pM0KajyseogtNVIhcpwq7v6X6GK11q4j+WoubhZuK+S
o2J2n1S8wxbUHtZ2rqXbCbFoBr+czEFBbaM0NMhuy4ANCqckyFOvPN13/pVdAKeN
VZD+sAxddntuRlj3IxBNsL6yC8XdcqXSzUAhZNdkUx5aC5VAnl743Gwe2/+83wnG
JdWlcR/sIZ31ImRjiCc7Q4Tn2Cp/aN3vnenGRp/xIH++HO4I0k/dUR7ToSsK9oO/
J4y7nTcJvZMAOY5pd+0GpFJCcwPtfasiYtnjnRqM+2hX6ZlZGbyWxZRa1x4/Kyky
OGBXGGqv9cEtPLA34x5LKYdw4NT01T/1il/8O+xdammHed7UzG7e+Y+5cOvsCpfT
HpaIDs5LoRcgPg6aHBjIAKQrgj4g+ROLYGjYNRmxENykqsNyFx8mb9pMdcrGWg7D
q8ImfrBzTraIUSFubIrxvkOyHDtNLVuugB26blqzjQN4oZ1KfqlvZW4BZD6bCjxj
Goy3b1gqTktA2SRGbtry0ey2N9jX35ARIqTPeTGn36AFxEzmbFJRCcctO4sHIN6O
BrjktSys+VSXFqFJce7ZbGrvw8YDYVXSiVT1q+6CHwsm+wJi6ZxbnmJ+8uxKR+MM
XWj7Bl2hkKdbDDig+vVjA2Up8/np9kZ3b+APsiE878QA8aKEyzB/03uv9Ov5JJuC
QunXC6OwiIXdDQSGFnhspQGq2/LeTEQYKWrefmUUNI3+84Clm3PF//WyVBoQUT/T
/87nKbJvYR8QFq8QFDFCEBLLoO0x7h20yHhugOEApDiuewtv02CbRHVynf7NLluw
EBSiqgbKTEFzBICjQixFSfZOLc0lsffY8ZTPN5dKyEeYkCRFS+C0zcnUu9kq3QiU
MuIreFjM59TjdiyOhi4MJWoPcKEznOPBcyHN6LqAYceHavfBsmCp4E8hcM2eJ0i/
bPTbWfNBQEObfQMrTgk0f/p+WyXauv5drXMSMbux8rMkAWonOOZ/4+6sez62DVtn
sC2jWXMjeugh1+Lxi8oYEiXG2Y/26ap1fZa6fMKax33MhDE3GC4ic8tL1n0Swt3V
5JCGL35DbJH053VgPydus+q66mEWKM6XDHGr31Ob8+Bzb4nZf3tANo+rJgs8vCsC
pauiMGodPAFZhxsbu88lykGk46doRZ50iYDtNCYDhLAemKrSlZqnC7ap+ymNbAA/
NhadrEC/9l/HZ7UOEWq4uc6EsJHInk6ebXomTdbUkMT8Txvb7p6MFxEhIGAOMpBI
izqxwJQOZ5pWQ2uZ6iKyP4zftK6z+3wTlcYVfGK6BhFYyMQhMGNq9EraRt61J3Hs
8lPm6XtqY57STTKZ9Zu7qhZ+emWXkL9DxlqBuwQyAJLBu0aUv1610zeI99D/6QHM
q/UaNFI35jy44+QR1mb40ybz5H8BZVIB//UwZm+wrIYi/WACY+yiIb0ejvPIdkvT
Pf7Jgh70FZHfraDzgCAWPZiuzYZe4Y2Hy9jEEu+/k40YQQj0wnTHJcdy/bOSJESi
SNQwuZ5Cp1NArvsLZ1nojKy5hpDkWk3sfDR3s2Kbor7Kpqfr1lHuDiXVzKHlQ4AY
dH5B8wHmB7whuKaGEwHCBGm8reu1CAYphBqaGApqyQuD5FAwcx9n9Gzp4In9i2/n
SypvYcq8Zn4/4UIz/pW7As/C094ptBeYTiY9mmj+uSnoga8Gweiy4shV8v6l0gTj
+aC0M1XCD8LbuFN6En0nQKiv43ZodmEdIn1vgNCG5iDNrwAFf71nJ2EWaRLFJ/JZ
aqF3kxPpK9mx3Eo9CIQxltx9oAH0vzCpv6GRKpJbQZTNNxhxN5eWSF8QWK/ZCga8
T0zuXlhWijJbWnnBc2gxx/uedm2VM30jexc9mThhUHfOhei4XAg6OseFio6ooi0x
d2ShJNz0dGRJ9usn7R75upoRz7T57J0PGDcPdewcb9aMBYczHZbNq0EkqkC2wyGe
0M0KZMTP2pTNnDgQbwCZhXBLxypLlP4CB4/hXCGV6sBfEQqHW/Nc2QnPED1Yhm9Y
vZc2/sIKBTRg5g/VUCOdsDpV3D9A4YBOVsSGr+DRovpyLwPjjLgEsUWq5TCRtztI
lChwabqrynGl+6C67jfAdqlrLJ3fVj6hN5Kx2KGVHZ0daalAaGJ034PwjE1ziLPG
090hLrab7zrNHVqoKzhjd2SFnncwjl1jO3PCHrpB0GD2QfClyYjTpQj2S8NEBfow
Y8JWbz9A93R2a/i3xbwCDNwrM+7GZd3KNB1lQ8q9I8UcudTYPh9gbFTadFofgnhD
oABYhnyLRuol9/A5IV5jX1PQFaKfmf98r6QtXnYnnhqRSsPdVWMU/og40KFOelhP
+wiBdugwlg+j1xvpaKbhiwrZPizS4rHst+ne7vkogot/1sGGVOFstNQycZnApNV0
IziFs1UomRbOjWztW9KQR8APLn51v4vBUvnal0gOLYamIGpzztNSG/MrWG7LWBoC
hixp97YAzPyDiA8zZUQF8alFNCV4DeW+n9XV/olEgW3Sk9uh3AxTSQ8i/Fpn2ToX
7UgRImAjgUGdIzRAuUBTUclHsNBAgDgwEr/MWo+lkdZF5VkyxrupN1e5vpMJ2ssV
dj2aTeWG0EiihGaFuCVdF3oc3wKKOz7Tbs+44ge+trFHO2/05i9GZFyCPiX3gkrw
Ffe+OLMqzc9S6iUa5J518vwNGbB3ocM44OdRpzw7g/HyauXFBmXxb9VGmsP4YTfK
xCE2lQtHpLH1NeoxBn7NyRSyBfSx1SmJ2sqoqs61ISt+PN4Fz9gjpk57p6EmF4uJ
S5p4Ea5AHbuyg1+kMPFcjnYzu4EQ0jtszL1427KlB5YrX3j/olr7OvTq2WNsfFJR
1FfOE8XwbDSOsDFb9KuO4Vw4A7vxLVzCJgmZByoN1K7TBKHu/lw62MLBSF7+ZPtF
sCM5HI+OhvLefwPj2FqfNuq67T5q5gAZonNblr5CTpTW/f8q5PdjRXUu9XRd0QVQ
UUYTCVfXtRRKaxjz9KXMJ+OByMncZwcHAsnBPwF8rxDIHl2Kj06Mu+oWSEsYth1b
s1OQndIvrP2HkVJQzTLkWALyidYM8OnE/+z1/0lVQFQuFBO+/SisRFNBMKgJ1nki
8LLR9TLAUd8N5zGSaFXPTtWf9Lj+79ZOJS25MoF0N/DvVjPxyxKsmnVhyz5ZOVLa
4JJ7YZ3q4nJHZtZRemCAD8k9OjNoH481cYNdR4HvgZjx/nh6Qs7u7YJmZ2Axo03A
wDG8quRgs9Y/MqbAErqwEa0O4BP1XCg+iYah5kOe5XhTzsxjQsArP1C8gsS6X09h
nV0k24YjS8pv3s+nQrOmXmfwnZ5vUoMnNkgnNbX22kQjSFc5cEx/uknbdlkkLD6q
iRUIHjKUCUpFv1JH5Csd7czSzU84+YS4G6FR7Q/+79LK3VGi7rqOC3KWymYOJmlY
AZnblyycX2TdiUXQmDmvZeRScohXrfpgtJh6zM1+uAasWfZj0ywaCceoVBP7+9TX
xKNgSd4tdcMztil2oziwAf8wcBiYyKZtBtWKxXR/sENpZkHIUBuIaSfnuobSrdo3
l34N73+5A29kEk3hOIdw9guKc6JqohKaOf9XF5g3cXtuFlVtyniyxJNHhdIY/HMz
b9NF6QwvPcAipZ7T6I+Qi9KaSeqsjTFV6zGHveWVac3CtYRyW4S8wovVdsnwUa9t
cESgFpdK51IMgaO/CHLKICMZ1hZdLBrublRij1WuTH1OlJyzzY8+Swayt1XAEmP5
8vWT3iAlDOzPL9XofC33LFw7PxUdjmmiODL3vinzVe3UC6ZqaFBuM0cnZ/2qcnsc
kq0/9ZkOr/TpNl7BfTPVLdrKbbx26YrK5nUEWz8n6h7KL2SGbpgepUHvZgZ0AnOD
Pk070GxErBw4Vud3Ex+KFHjw03Ys96Abcor+25JDDxUjY43FSgB7xpVcffRDOr9s
X+6kdm+HubuaRCcoxwqfyFBSw60Udt4YMWtH1bLVYFCiw+Sp4zJsHO8kNQn3uCXO
v26G/G6jchCAOqlGrY7Lwf8KzvglA+ST536AacHXTcYzX2b4Q89lieVLv3LFGg25
BJ62lt9tzS25A2y0AKRDOwJxyPJW5ZZIOQxlsrjl1TnT1bu7E4Sb912R8M4sB/AV
c9oCPeiVlfdep/vs/aP0InQ+ryAhbkqsB7aJgzW6Y4Zj/RS3dSz2dM2ZRQJj2uJr
1r07b3hhVIQQeeotSPEVuD5lt54KcDg2C7JNt3HuLU+mtvO6yozPLnHUmsbSevbA
pKhpZdyoiDG3Gsp+p9FmAGTyfoHtsv7J6F44G00i1PQUqV7107OYFXWKbUbpieYf
mGixKX8dTGqWabT1j1dn50XjF0zO8Q+S21i1NK5I3PZNaximr+HaFNremiPxl1El
3+fNUxVd8mg1pZWGrTNgEwBPKUKcDzZMGryVNywER6NtspZIRLtlRz6yoVb/PqUj
QKSV4cN0ciMASRoFOAtRFNErStHmHo77ECfrX9VEi2GiloPXNW2OAojiebuw0p+p
8sc17HzN3yKEtTjIrN4AnYKdwxr/KrR2OD0NstMS8t5jHqdo5IjYpRTqsOnwaOFx
I7PHXbUsy7pZrHrxFidaFubC7bGjcBebm+Gb6Shm/lv00UyYdre+YL1JYOo2U+ZM
Q4ILoC8az0AyH9fR7WjxbfD8a4PIaXL487wAENNXLewyC6rT6xnRl6H/8gSvCiWT
C1fHjZ1K6MUnwUeOeEB/0zZouvksSHrnj+mRzcad9HQrTecs/kGR4gHGhHVTO6GM
EQ0ILXD0JLh8NOyW4O1TEk6pwaMmDxw4izvb3z7PL/7QApCH+ArcYB9Kbhh7z1m0
stmd6A6AW0aYAqrkcRa23eLZkWJzK2v4n394peNg7a4AuriKoBws4KPNksRQHbjc
1HwsN1nbtmc0ujhT+3FzZ7VkwlUiyE8qiXGb7+3J1tJcDI2l9qBN4KE3tffxyrsh
rT+oRa2Gt1jKmHwnAPRxERlTiF+LXluBjI091CP+G1HBPPyfs36ats3lG8txAhH7
d68gb5W6IVbom8bW0EprVfjuFM2Dr+IOYAm9NUigQgNxgxeTQnKvq8jbNEow2ie7
SN4crvc9aNCLa5hqbuaRJ1RTlM3YctK5F/UkhoYn4+OoX8vRmD3nlmGzc1UZD8fM
ymH4thIfD+lA59Qd2R6h4NWnkDVd9I6dWWtZvYozd849a2W/YDYR2whK+qrmVS+R
FE0pMrHHvtwJ/Il0zW/CJlcPgyM5gftMS9d1S0an8lWyvmfbPNb1avLxzIKCjiuD
D1JZTl8UCrJ4bdy0Tdcio8jIlI447cLLydueSc/N89Q8aXirwrSCzbXf1l8fHEcr
heq2Rp32qZhPy7TlJifmVApwxPebIje8O0Lx5YgY5oClzBfe8EsjkjnAW0uY3wk+
PzLSJKgvYrKrtcpmOZVw78VlSfLD/K9uP8fSfQD0JDF9s3iMBbqjBU5KsOG/v4cc
gZ10QqW181VABV4OIf3v0wu0bprOxLIBj15ZBHlP5kRL1YQJGBKkfK96v7Ha2Wdr
h8EDDuPZ6rnd44YgikPd154T970Zu/9HjCH+5hcMGhVcaDQmzkwG/zK9CJWcAZ38
dbVZYUAecPnvn0NsaQ/2D2ywp/++xe37nPeXK6g7X6wlQmjf1sBBF21yjSj99l98
lIm3Px6fzyvsc35kE6ztbTiv+nnd2JSQx/nG1HLA20FxhqnUL8hi69DoeksCJueO
pppAoNaXce/Wf9Mci5lKvpKql2CmvfIRyFG5Glwbu6K3x6upmP6fdaGyk/6S6MhE
747i/zwN7OVEsJ3ivwCwFAxOhVpysSG2o0wxGH7n9njvYN8OPWOrcX1J8Mz5WaiJ
qBOZaFfXWhASoX4hHi8q2t/i9zX8MWay3qM2gTdmwg7rubJ+fBsLd1csoJ6qEoaV
QYGhjsA7tPb9zNWICHneLp08+ILfgbr+WzjunVkGXZ1iMRTHj300X5ZkOxfgn0S3
tJ0ijQ/9qtJY3XhAAP45qOTAPPrcQXHcfoAfsX4QLo3wlqknAY3OKtM72jBN85U5
aD/Bk7lKUyenTFF3uwkCde/tcgsQDVsvfY8HTh2Sv+2VRCxBPHSrbYZdoASuP5KT
JaGWa0CyFlKSVfFUKultAP1xgRuG1YlvGE3n0RtN+TqSeJad1S21OeFcY1o6N3/t
btwc062gcJk5pD1SS87v9yRXrHTpsJibouJoTVW5CkFewg3jO9f0xfjraUyGDCat
THy45SzC6RMSG5+DYxJZ5N8ReE43Oa99YskvZ8+GUPU7qEMnUhBlGtlqAJ2qCVzG
ASKOC5odAjXB8Ss4W7t+K6DMCA3Jmd4MkDvI66xkqD7RSYQqSUKhqqFNJ8lJse0u
QZyoeLXAkeXl0LvOQ18GPOdSDAeTWnn2jDbi6wcV73Of32BP5eIDzjCutv9zjRf7
wk9dg5D7OlB2ihxn6MoopuUeOxNie1ANms8gbCx2lJAMUe5/uEHWOShpCAvb+oUQ
kkHVfIG3D7ASFzwVccAnnJUQe4dJWEGWRT14GM6qR8VeumJSx22EO8pyScay9J/6
M41x9pQG+Ks0p04HzVAslSutn+q7VoVNmSx4J3kIZ7Sg66hfGJm7WuJKspvQ283N
7iMCcJGkp5JsaXE+wUDoyIzBDCTgTSuLt7DXdAw2GSEpuebvjlPFfsRwY4MZa0Rl
u706Nai8Bbkl7FRcMf12vYRyh1GEfFYrbUj2M70g6c+8QyrQVHCTdcxWXbEnKG/f
ajndcu8bSXiPi944s/xDHKd8uaQfhKx0Zm16/cFYGOUpo/5W5D39/7cuvLOaxZ77
13xMtx5kJiCWXEHhdvEYalOtB/corDeHmwuu1OQT7og0X4U1O6BJGpFoj78ldfm1
f3+f4qyhcWzQKzjsVtIcgRa1ehmDt5kExVUrJNbkXSA9ygWBHYtz69KJqV4JFizO
Bwhl5GDjAFX0xQy7+DXyqBnc9xWgDOLFUFN9r41QSq5yof8C00qas9x9I6LSnoq2
nA8OEeENkvb6m2Hncij4yBJgHUWee9Cy94mJTXel9M2N0jx+zpe/n8Ik1eNwRWqC
BRmS1qc1R4VZNPhxbzG7WyYShDOz4JeC6k+uwZbwKP18+FTu5Jiuh2cn/q/ENIxm
xYMZTAJBNjFPmf+wk8W/CHH5/jkJ873IYAOD2X/fb/jf2myuyJdA33mI3sQ6N0U0
qfqIV2lnZHRODtfbAKNB+hhCdYn/J6o8JZODHbtfa3+TQy4IUc0yqFuwVoF0tiU7
PvvdMBFk2/Z+Jxee+m78gQyJ2086KOPs+HbSbmks1ElwaVLm4Sq3lnQgTCTd+d+8
uF/qkvOtOfKR6f7SIVoKnv52EIxRFamvim505lqnNO59Zeqq3RBpEFmsVZ6mdGGs
2h+zZdQZmISema+qAvM96+b0aB3VyenC3txPzYE9OwD+X9Dy9LL55L+tsS6fceZh
GVeY0U3Y6nmoMb7PcOwpCzx3xGgIXdwP00+IZD7I3UTwmtGNf8EexVje6cH5RaHg
FuF5i55X2wOeS5WqSu+MnWD8V43gh2uUzKf65NvT6oRYcYVeYz6sW1ho0Mka6/WZ
fgvZkMRtOTSdX1rbo1aMUzU8MVJtAuSLEkdabcn0WwNiU8xdelxTH7YGn9TFCRaf
ebEoVjWcr2b7UBPOCyTvsc6w3KcpyB8BDvcnVbic5q+QL9E05RsfbxXqb0D5O7uF
GsscJnOeTPqZzU2X8KFlUDlI5BFlYfQL11uSXtScrunEIuQjfcQOIo0sTiPIhPVW
Z7D7bvdD1E7nrTOJFQsGvHq1MqbdMFHGnJJbDW/hGmLe7pPSRWtWKZ871wYr1KX4
a0QSszbsTirShAGSM1CjuvbD4zfSwb917ojWUKIevhCMVl4VeuU7Sh15iXV0eavv
uBjka98mwaZww48fFJ//UnHzNny3ASiuQpP8Nc4jQMixFnIM6mzvc9G8U8XIuT2p
2CRGfQOozBhxOUnhXk/fIKC6+bYg7GS6smeAgl90lgy0ywpv54sqw5ULR3YaFhtG
+ttIkbMQfpt9Uk8DqoMRt2L4iaifIvxoXLhpCgwQ/V8CAR97kTDJ6WPZynPpfBFr
h6eiv584rKAYeVeJWpPza5/5W5zjBEdYCpcaMK0zsywHkwfFZLBOuSS9DJJl3Kwv
0z0RUyfhZTsjEEf+pM6MwUYl7UHA049MfMKa7mbUdRMidi8U20hO1p8HVu+wttSF
3gpgH3KIfMa3o9YSAJtSQBNM5Tg2tys/nUCrHEQz+/doFaYoq5ltdkP5aI3R54Zp
f1Wj0cVaiuJFCJMxpZuPOi8MKd/2nCDLKf3otcc6hpj5Diubpv/sqbxLrfrfwLwu
MnFK19i8N3Mk9fmyx2H9aOS7ncLgvm7mn6m0PVswXw4u2efzTiGN2buCBpuac6h/
YAsWeUSC4vrGUfnCoFQ0zNLJKRwLKRiGGA6bbHCXNpwUOPMED+266ZZuTP8fA2Hs
X6fFGAFoEk3DO9QsxgUlNPeTPRSJieMuubXR6h/APIPh0KBNYBmnrh0oxSeVrf2z
PqlFf8TbcT0zBask5l8iLRjZHR1Z0L/8eOz7XmUIjAiC2Vr3+bp5oSSDXIPdMOzc
dOD2lN/P9JPySqaxj5571yROqOVRYmVqnqDx3dmnr7SNbi34p0GPgrTDbnuV+rWI
tD4Q1bL4huTFeZZmWwkfsSiRT/a6wXrIk/IasXgCqO5DnrK2k7AMJ6k4XE2iBwvF
IhKlm9xUQFF6aSzNpGknGvSZPu5wgyldb8hA7ub0jAQPq5cMD53puJd9v8S0a8pM
LL50iE35GwSeKI4fRzf07yJlemdyrMVf/y1aIV/WZTP1tttpOkQ9t0h+olkxucMz
wu23LbNDnnjh8KE1pNmVxDkmN4Ydu+PsW1gglPCGSE0IzjD1TCHOKlrHjteaHVA0
dN9MiNaofW3kjEFFPs/pyZs22FZJbTmiB30h/THbi98AeDmIPAYo6OwSAG05QQQy
fGiayOMcRL6O5LPK9MSR2mMc6a84jnnTy+cKRUiK9SA6XLh9eY4T7LPcV34tUdKc
2jmpnkauR0TIT4qMUwxBb6RrRLI7bLBnChaSYUzOSIs3VtYZNpW6C69nSrhR6+Hd
tYSDyk6Ft82Y9Z3rdar5ybJGXYnX7YQfyDIxs0POsuUi0gcPnSMkp/0aHOQSuMeT
+lGaK3oNZ7380gqCJDZyPTOFmnvkVfopZLhSi56rI+Uq3xvycpK3Z/0OltB4EWoK
el4a6N6YUr0+sPRKwpBwsBbp4/uUe5TbdGVUnjxuC7aNB+gvo5JYd98PIDbZKWIy
2jk6cPq7g8OKaoP482gIxiJZGFXtd+WkulGi8Viu3ItKRdFEZjCZjuMcc4KMCCuX
GouIZMJiQ51aUd15v2JPmVq3vIRsFSVRyyH1xFehe6yWV+R8mkuzgZ8RYhYA5LNz
iGmCJCUtoO5yt1L13qy1zSLuiiBeZEFILeVV6y9aNdWjKvs6Z8dfM9T+zvXQtwJc
JtPaCVppk9JuXuxVmi1XU0RsF1ROKKzInZzzlYcxyIGbBIqEEPwicX/gZ+OvOTUG
OdWdlmftD9RR0QsmOo7Z5hyN7gGfmZTnpZF1jplq8YGqLVpK4d21NZ9lt/+NY/gS
c0W6MKc/lt0qGkNHNXb87kozfmyjbIxhzP/WQwHK4LzeSnTfdw+FJcX/Mv62VhzL
3GEjqnhxyVTEm0MUzW/IbIgqgS4NPVUewHw6K6EnVLXF1tSWzcQsS8R5QbBfr7Um
UBc67MX/7ednSuxrfiAEN3djup3Tj0InSpnywDB0v81jgAO2ZQIQ5c0sgfx1TOwe
oK8mykzKShdjjrnLJjngrQMx5wEpfphAcw8e10CNwdDlc90IXaHBqn4qlFgl8T75
PWNyxzSAClUXolKyhpY5lkbrfd3DetlJca46JkwXpCGVvvT6FRN+IB35kVd+F7i0
vrUWYVUAEl2BxKy7Q2yByT7IUS7Kcirx5HUTqdPObWd3O0ZepUq4q8cO7u1v7aYg
ow0V1HxduA78bWLfAy2fsRlCnHEP0UbHelRkTcolrBeYJPj7mM7K03rXdCdn7Qce
BZYT4gAYIZFQMIlpffdS6O05KSwDEOKK4tA6gnhzS5Sgt1kue9vDHQE+OVmONaxk
G/A7CzqD5/MRGc6AMowH2EIWC1DVWawUD+ajOZAhDYJz5sQVZJYuXV0qThBmI+RC
V7g4DXQlSFVROhTAk/U1moI2Dtd7QVHGtzRJUJPuEsAHYzvcgGkkLTjbbqcstfBf
t1haVf9RQO994eIFyNfRW4z7asfc3PPHdxR4ida2oyWvjZOA4yOU+qLi9vt4G5lB
/9eipNWu4OAfe6uZHwQT72H1PNXl6vKZqvpWAH/fFSAaPpFvs4QowQ836E+yQRSO
630BsDC3dRnX90mPtiEJHbxfY/M6MAMeXz57O3xmD9BFA+3cWzSsx+uSJy2KXsIX
nb40Z3Dl4D76yoabhnc/jkhX5t/KiozWWwQz6YqwEAgAECA5d0Z10H74IOxetRF1
cQPziOPhlyn4wmGi0g5wH6r6nJUk5khD1BZCySM/qQUT0bPRAWSMA6GDwNK+ibOi
84CVucJJwgwp/RyF5Ze6UwKSJEQeuv8oRX7LJ5ZsFsQ5efrIvy5lUBtMfmEjyiV9

//pragma protect end_data_block
//pragma protect digest_block
gt3Yiiza6dpDbzLG7RlM7qw/s/M=
//pragma protect end_digest_block
//pragma protect end_protected
