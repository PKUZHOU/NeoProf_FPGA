// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
w/qUP4n4dwB+wix70ZXLEPvKFehjWe6jvqdqh+bWtETPG5OroYyYqUKFhX7MlynD
foYwTLM9D2AZvhr1CTTbghr+bNz2vI/6k75HFZmTfPaFxrWBH6VQxsKJvAfaYpxQ
WBb3gqTBI5+GRJNAtji1BDcNWFHq2k+mcptaKU5KZns=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 1824 )
`pragma protect data_block
6hdJJanTUr4nPMsEaQ0Gf4FTmQrz2shmfvioBn9EWSkpP9AkMVhsMy8aMMXmKCo6
aMZmnjhol5NcqBcuO9oFu+aVMNxngqmnUwPI90Z5toNZEOgvyhBvWdLr6iDuveKt
tvOFYylxZ2tlkiB0wxeXEXUcyx2lPStX+/+MVgRMJ4A9Kf9SvaL/XucER2Ewf1Wp
l6REhJ0Wxt/4aL5Bg0nkQ+z0eaIJXvuoKLdfT9v8kf4vsH5RA++vJMIiIW5iFlld
FZaRzu50KUGcHzQmCnHpBOTc+6uhmn5GBCCCr4wxDt6beUl21AiWSzNoim+RerUX
VGuO25uTS+VjUVMLLotjwWRDCF5XrRb7sobww/L0HdDAa2axB2RwZhHrN9+khGoJ
DR2k9i4QYWYEW+CBbgkKq53kqsuefNDou5cY/vSar7ReHGYlosWaIuKnCr2DoINf
5jp/49gVe33ahpsCT/X7g6i2tF0sa+DM1eE5kc5jAV7ae8nyXLvrra4lpbLbCxtF
5SzUZowZp2SzpkPTPqagGPTDIW8R7ye0dOYYYRc7Oa1QzfaR3+REWWmPhs6gKBkA
i4oGyDqNqc39cR+Ldsa6XMvq+svbGRBiUlt06TbanGQ7ZSP0SWTbQQ0Ne7uQx9h8
Ffvorkj0KdBv5l/u8li46wsgCr/tkm7Ke1BhqnVLxpjs7xQOMyrNK1WPxFOD2e5v
mUmvrndTJs/ldYEQZ1fkJ274b9IjwShA+1mpYAOvE4lcybIBp5jNo18b4BHo/zVa
cz3nQgbAcTi8QsdBNDBcE3cNcvhmziYxHdmDMEpOXtO+FQlIKnB3wRqzf8jHe25C
y2l2o932tevqhQ83hASwxGM7ts9OpFvUQ7HfNEWCvf4SPJqd0RjynKlfKbjUJUms
VWXydmOjupOahy/suk7V3AUovRvbHOXHJ9v2nHCr32xy45iytIPw/GFdd4mupUD2
KPe9qXvkPQ66fHIQvc5ayMsnMnyI1ui/rwQOhsLvdTxvTe1hNeJIGYqXSRt3N94E
iBvpEWE5uEcdVX4PES3YoIpCLvCaGKaAREf3FyUH2+AQqGWmC+wAX8slOtofjpq1
tEjb4qAR9H09Ws+7sxnqdOy7LxJLNFtUURNeBBp85mtHtgEHNy14NiAlOpGAJgPr
u/7YtTWnvbBETyXFJvywJJioooySlnEGEMkvrmLiaV4GaNFWVnnw/YKjsKXA1Cmd
b04MXVa6m0qpE73XWHR4kV/JKUKLwL46v9KJm7TolWXCDiJwG1WBJx/BVRvpW5B5
+zV7SvHVT3AEZUcigMROZuMxy20h8BonFDmHKQ4DDV1qBrtEHttvLR+b0eacfGnm
RVE4X5TjcQVFSZzmbHesAracUepQirLddeGuewRpPDegjDZz/DC8njW5Ulcjhkg9
cwKPvpPSSK3Nu56GC4LnErvTuELkRi0ybQ7uetsamfA+7znP2H8lQGQrTrh7nxMB
Y+xWIQrdLH1h6RT+7u8mFD6aQAYPFJyk9wr6UB8XAUZZ5Ws5IEH7KY0U0DVDrbRu
ThHJxLYwY+dJkviaJ8Qn0kbXUJV3N7mfGHu5qIJkbxgl42o0CV7vsvQaVaSEdLzs
xFXYRinK1mI+A9E6SBKogyhXCdH1rLh/S7c1tVqnxOlknrx8nbYYlkEPPFzVmJEO
9N4fTjUOLxveo6w8+X4tu7VgA7rfo5s5rdRjNNH7bu4AdbxB2bNyWpaonLv2EcWa
ioTMNXZ6t+FDW+aufLKP3wAJkIwH/LnSeM16GNlflepQ20GXlPKE43idwA2MPKfk
S0Ammzy66PQIbFpTZNZ40II7eBLhB86fTDchhc64yAhpswfMONTsusDvexd9+n4v
53wF5nR94CCIoc68mS85lMtEoHMKNi+acVl48n1UVAxTBGukPxx02UcsM+qOOk6z
Q1bzrBekhx8/1CT706eo72tsGklZcx0D2S4oVj0shXMpVRKfFHgc9iL1EoMj2rsz
GtNVOHlD36kQQpCsmriA9ly0e3hdEn2xhcT4g95NF4tYBy9Zyr9k5sBSSMvpRqAB
pAtJ0OGjwJm/Y3aoCZtiPuqjK1M4Ah6ZOSMjqA+WWOT6fpcT2anI7yhMGjs+oF0Q
+6n2/aYZKxzDpnXt/zwhYpJhkBHTDy42dgnn0ZYzPcqL5VLKAyXTqITEA5+yZvn6
opOOMAZL1WkJyaK/tlld1sJDi44fwW676/mtc/QZOP+eWjOgKdnWXkbVm2+99UqM
RkOPLzhLGVygkXdStwcq9VCgxzA+0m+7aMrww1t6cDTpjCxBc8o/17VhU3Q9zT1+
riAcQ7c7TVYYqrGWRkm+ZlnifBwAlzijw/2P3OBoTPIZ/TCL4Y/0UWzIQHbUwh3q
c+g4wCD2oW0Xcqc1HzLkOZIlv7Gzu4L2JJ4XqO8ypHKeWQmoQUgZzSvUYWCqGh+P

`pragma protect end_protected
