// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
xc1MK52yo8YqsvdV8uClyOEVhpJQVGoNpZXsu3VYexaNnOyd1DDdxOYR4KGtDN81
DZbyeOJMdfFj33vzjZSGaGCgswG4RaORDwziirhSbXdZusvBS5bWjdbVkO/ZuXfF
612j1AoDKFke2NQKdsIpH3nKe68vPHyVnBwgDtc89yk=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 1376 )
`pragma protect data_block
jSCuNwPvN/3Owb893x1lWRR/E8HVH7w59bMZfXdkfS31acJvjUhHpJp2CDb2TqOK
e5XuWIGVaz7X2Ix0EjUYs/YntiXdBlMZSNI28qeQE0+sYP6c703A+nGnAIzNhemU
7zZwsxOnCBf2j12KPS4H7EImnsTFZ7+vBCYTS493qlLp+2tSjyjRhdL7vnQBrlvj
ZtiTM4Lo4EalZ3ErQkLT94bfRuQByP4NYLa6McKCbU+HDFuaYOzfYu4pYSJodcqE
yJiYPbA/a/oQxkxl1Wp0B46Pqi5QceGtsgvIeuYHxScpyqaBuy2aBGEHKtALFB6m
OAehPYjFULZ7geY5tPhi8F0DmC/e4YRmbLYIK9sOYO6/zlGn9vP2IGLdF7Ebz+yc
9HwyYGyaUwJ5AxdWNwRpGfOwafvzO/TKixhLG5NbTsRh5avl2WNJqNm+XyvwCPRw
Z0WQ767eI4gk/v1TA4sO27htGYxlmEBPxe8OptHCYP3tgspdlJcHH4YYscV68Wyd
/wU24ADXKEDTvjdTeGIYpchsnbCgyws81yio+d0TkJ8b4pVtxiLFRj6jkh3auLvK
ngj45e0DDniU3XVO+R0zuZAlEoWq9kocTxQR8MkePPH6ph6FYrzZz3VTbyYYrYuY
KS9lUVDkkXZarywl8QzfNlQ1EgQHWxPCaWQh1JI/wlsiawfV3Iw010EHsV8g+Ghm
cKSL1HuebVAscD9dguqgZj4lpbOrA614D8MuEqs0Z24dcIGII7QGiXOD5gevTGD6
m3+qVXzOTxXxmeyKqrGpf4Ubyg141/nuzwbeM+9tIm5D7iCOUr1btH5kGB4iCTO9
+l4uKZ1EFIRNqpFsPyCUpe/7WRKQaq+RLk278X6oUvySSqlEl6AwCxZ83FqUltv9
LyrhrOS7eNPr2PNYCZ4Y0+8PjzAjmaSURqEPlDXjZFXSz68aCancAvE7BliHWyki
JCugl60O4lGz3txSRra7avqZ2P3tj2fENUzVa6fgprOGktC/SDeJWsALF815oAbt
cg4VeZmvM6huxJR5uALPx0UQN0lNFYDlC+JqJkgL07Ejd6kXBV0blcc4bX7Gxlh5
Eoy/FdvcntI2te1A6CBzPmAXs+74NMIK50VlryQZOylx+VDW99rxbuc9hLmCLSIz
5lDSfwGJG33wpaSiXz48VCneSWzNh//ehW3WmF55KHX8sZ2/su+Un4fhvmBOf377
T11TI9PP1KAa1HmBwgzPreXA4aVH07XDZbFzM+gOv5OvaYJp8uMJQgwc+UvXfBQI
l2mXlQxogJPQR+iBimB7zmYq42Tltl0koeN6SLLBJg8Wig406LQTepOepVwtmS2O
dCMUdV1UVEamBDvmQSaNFDiqTCSBvAsK1wqXzUoD3Vq4lykQ1m1jl24TGuAvDyUT
YJQ3e/OWcHMBMURWA1QS4zndvnx0QvMg1vMoVEqU3fLDJD5OCvZvB+jEMdSsx/VI
2TjSvrWOkAt1vDv0BF/Ge8NuyiT43MEhnBWJMZW/hPLy8kb15YHOpOhPEPjUsOBk
81miq4e27Jh4tOJbHM7wanUsLoS6v6ml9EhHfu+Rq/MKw000SV+rq/doD03/26PY
JOAVcRP62FCPHICikfnmbWce2sUBw2hDtT/+iFPaPUR+N7VNHK70ktGaWV2NT/P2
oDu7ECfTlgRcfxpUYJ/WKwg5Iv42IFlt3E2KzYLnpO7bmldrPpx+JVPqu2pSr2FM
MZUsQP9Q/12/AWHr6k7sAhgTVm80F6b066b2NKXGhFEQkh6ShpR4AvuNYGid8PHy
B3xK5DutBUO165Lwudi5rMEo3cmftvHJexG1qm4NqJw=

`pragma protect end_protected
