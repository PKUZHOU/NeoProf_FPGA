// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HTDp8z3JrxvlBZztkoii+LRkRC09JgfwEQF2Rk+Mio/iBv5EXVtzDLRvZQOk
nVZp6wxKgS1esMrJOFGWPBQcvR5fOgK1MIUNKfpFta8t/aPVOa8e4KVurfEM
acpEW4HD1ZTZ4wNEyjuJeI2hJHZpeUzbTjlHIBkDhpNufGUxvFTADT3nZxO7
gd7jA7VONQbzkgBI7AcQGewMhnN49mcL0lhuV2C1Z5+VKjhhoc0hLC8Uh0Ru
e5DRzB/uJRoL1zFmXXMCtnTrKyqhO8W23SZKWqy2BNbUTS6L+3CMXqRf05MN
ttJ5aS156hfzcSYT+MLGojzlMF6vBw4t0WfmjsU+dA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
MvsA90+aujuPgUeAgLHZTT7ZpjMccfQnIMXSXlc6BZUWwSDcGXk2cj6wPO3y
YX8zTmeXuL/M2y3iePh6r/NQeKuo7SMNWDiPK5kZSpLTYDMKFXLeknDHrxxS
x7n9uYiefZoiWMsutWH4L6lMTFb2v6p0tXiKXEJeKLLWVORK6svFyGSaGro0
7TEwg9nMVp94Ylx0xOe9ou7VkHpdMqyh6Cp5PpvLFP6fdlOPAu850Pstn8SS
TNHwlYwsnVxs8YuiS3ktgdEzfBUVpLBNVCWEI26VAlDUrqI8ZNrdG4Nq0pxO
y+AGqwGP8XB68PmDQyj+y396MrWn6hjY3unRfa74Ng==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kkIRo4OoVblYW1BpylpSRd3WtpfqDQgd/xSJIKS6GubLQFqR40HLMSYBItti
eTBClvm3oaQ2NnwCurqFMfBmH52tKol92ClOvV7UUakbHyAGp2eOlN4uqRzf
KVtfIN7JC9Dnfp0hRg8tieuxD6DyiRJHttfz2Q9BSOLp4U7xyNQ3V5GW7OWX
mtRVsCCfjwKmFeY3m7OworlzbLoiq3PuDq3rdkAvtdca+GPUtYmFSNWLryEC
A7fBfp7nVKw+QTet5Rqm5p8vbEMQYA/KdVFuejgaCjfAtv1JIZF8bsKDhhgC
kxb+oJx25mo7caf8S17wsC0uuvN/q3lLRjG36UHIIw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
mWtrUp0k/3S/FOe40dhD06b+HTVp0CPuvw5MCVYXlm4z6mDGz1gK9K2e/1b8
/5pnaFWmuVjDT5n8IO0gSfr12iqsONeR/IFgZgV3H+FazRiHRsNnhj22caJx
EG67DQ4gFVBM9dLvYz5axFR/qMcOjNKjiY6wZOXV/bVIlzPiA78=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
bRHtMJJFykQLXBofDfrbrDVyaecabRIpo0QkoqIwPHXf08NDxwVUN0B3XaNn
MqWeAMgCBVJKGof9nA+kA8PnYbfh1K3SwY7WnIWCjhQHvlbAz5dSeZktrBl+
CbQgPqEHNN94912zqwyW6HXgEJfQNjtC5RNV2Fsw8rkfvayYiYqu5xhQDipO
ZnuwO5pn7jYB1JGEMeK19V/tzP2b7n+YKD6ejx054reCxwRT/LHQNoaWLt5z
AI+gfdUqHE7dRPKsHS/s/XzoYe6NognKxg7R6Mi9Y+2fwIx5NK5A1ailZBzJ
xISsW6lVzNb+3DMOlXO4w1tIdN3Vv8T0nRNaaDQRyOauaYNLMd+v00HGd94h
oe8nM7gHFpaVGVADRD4QEjLebfx+SxvEEeJx4vfLfgTWx6zGrUZj6Lo1+vNa
zWtNvZkf+Pqj5b/6GM/wKzViIx3s9MgpOcSp5tZYKhA9gUkcHcJ3dWSYAINV
UxczqM7YR0CLIqScmQyndEay2k8HzpAP


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
NGwb3XN+V34N2p8NVHPDAV5BG6FEUE3yyVHZp3i6uo4V00DkC0kWrSCZAI9I
EKuE/0MzVkaTf6SpQjR3oKunYDXVJ3WeXUQE04IRN64CkDrBFxmUnxu9uuFW
XPcWN7QE3ulkQB21W4W4GQ5zQulSXEORoQFhgAfqsL2/CB62uQk=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
soyGOruC5mUWQG//QfbCuPKvE5JRwP+Wa/Q6F0sGt04eBK1YqBWP87/oFBUn
Y3MSaHjsjKj+u4LaXK46lqWnvORIqY2veZ2LYGZIyUxLgFaWT6x2y1xi3qQs
IACr1OKuTDYsoAz90jbcJKt3Yh5N4gOPxwikvSXigLIZpaSoex8=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 6144)
`pragma protect data_block
TrfdPqmA1QiBbnDl3Dbmqi7DRwoToSpzQHQq4Km+elZhqdqT8qcuH9u254zg
Udfybs24otO+OlXz2LSMVT92A2KvlB/cz3ccmSaaKGyXa4HTcW20dCCPm6zH
T2nDrfL2dOPYz944UK/1Er9k68+R0PYi2cJq1LTLET8WcnyubOHztD1Wr0vT
TcvrMZCH0vmhxG0klQTnFeE8BRtuH0IyqCLWPQRci6AFlEFlyAgYGrUOsRCB
Cec1Nry7eFLMrtToq9A7C6O89IeFJLhRRj6ICFWC7xdFp4ZgJPtPt7enEpkO
pvFGeiHvLcONuYbpb+JWcObuU4LYYcN7j7Sgoq7W3WXSmJIzJeTb5v3MblJy
JdJHy6LpyW6P2MclqJJASmaZzPfe/3S2KvHCUbqnGElIu1iY1aguPmsNGeX5
tF071BClmNPttOk+Xgzx3O1jgovTpIhOUGLsbQ7rV6urzs54C6Rg4/br76QO
wIrAuGoI3jTTd2Ifxd+FLJtkXKDe+5EybSslm8gEWqlsK2ec+pyuqv8r8uGz
Rw0ohlagLU+O2dsOj2lMVH+N00WrD+1sObL2uwZIrOqbkPIPjE9IrxD/hfH6
cDz5v4nEv3QlCwKeo7g6drN/pgWO47+zD5ZokUqhgXh6a3vBYwmXBg1JGFtv
MDWxjZcq2fuyOfruuSGvhV87rvuAUtj3pQ+qF5/pX3gOpcNpoqNNbEwI5Sle
m/7R4Vamf8Ic183Q5qQAp9qixFSj0ZIklMemJ7VoN6sN7gIJsr3SZV8JBnr5
tF+CT2+oy5+gunMCT2eyzeo8YyInP8AvT11AqrhVOg0UiL8MncvqrgGtUO4d
s2WctwjPcb2PVF4uChgkqHh8IVwfXvnIBjqxC5YlRnWq4ScCptj3nrE8PbaP
JF4rgdASHlr5O/Shmchobq17egtQyaU1KFTo2pH3fSwNNKArVBpwoZQX5QJy
xg25UL7ASfFlCAoUUCq0OdbKzB66MS3vlXPQ2LhaJrqLiZCw49FaNY3gtDLD
qg2L2n26KPhUuJW7P/OyDj5GllJ1Wc3+47ImkioaF5s2urg5RpFCpr0tJJ8z
227MQRq7OcAiFQr6q/lupPxuzDUGWST/EkgHRfPKZZigysSQIifvDmStr0n9
aa26+Mf6IaoUStgAGthlmqVc9SpDVM23h8673StOcQpLwVzkVhpQU5HgQ4Nh
xtaJZ367pZ98OmS3GUHnRWeMZj3HItCIKZBoCsx83BrEWSkH7bWozemer9za
HF2BnQ9TceHN/pLqZ0BWjLPXeK5Ma0TXev1jedlgo6I+Wt+SxCA1CxOHxcuc
JpqLexXd6ovJ4to25C4OYTy143vAztrdZbnuR2NaJnnkwbNTUreKGL3eTipm
Pd27uCdfIZMw41Ag6ovOyhdo4kNN36Lva8/8OS9OTXhXgsk8SS/Km5zH1X9n
FnHQCHsBL4LJWm6oY4ZxRXmjoY796ppPh/exA91OOf2L+RHj9HR3UAHIuFmC
/CEpmSoNFNh3sZjCzng00mZSh0XOSL3+jZD1t8MDY9PsjbdSpvSRKnFpjL3p
CHGsVmRgqbC900V0+wBE4Wa2PhhBWikjXjyWropbutZirisS2dc2yEoU2YKi
gkvoM+KxVgipUT4VboAOsdLCpkqlDwQwVYcVcocppgksB8eEQEKwDtiz9pqi
/X5zpEhpwTOyOnbEwOIDcQT8AiALbV/tkkj2kBU4ByJnTIE4yp24oWq/Bzo+
uPs3AbRRHRC7LSuEZ7GX5DBKs//kSjr56aq4/IaJQ2D4V2sA5XYi/cRdbBaR
hY3BEgOJ84ew2fpTBF+07HrQ6RMyQqN2Wp8esbHDnONXQ95pxpfoQgWVWZlS
oA53Si4cP+cY79zIgegl0UFDbjS/Q/svU1SzCrPxu3qvlyQI8l0yR7sn0y0r
1xfUGkARMEQ5VxYXQEWllPSJAZaT7C8E4ycMjK91HHYfdwikEHqMXpJ90ubS
ajIX7jGdCIxj6+pj3z455kmFs+cUzF/T3jYrNb1jQKsC1EbM2Qe5ZJo1eC76
+uve/T2mmyDjJbCFISINy2r6bjcNw5XNGsXVSLwlzHYoD3SuQudC/HFCiaON
KPC/dEd/+sox1uypKHfS88Y/uc6hqROLpcxDwA0xfDlClNFn7dsqP9gzJ9ny
Fr2cDJNysxf6QtsqOOKsI2qtvGs0Dh7l7d3v1rIq8ufZlqgDYKqfwmwbAeT3
r/4zxdmExGcSOvLEfAe1iJA0usjzz5FyhBtJS7xp1VmVxixdoiHANxKz1ugW
ui+DhAc1PLc5IXb3kSr6zYLQ3+phR8GuZxNpKcMOOaQCnoNGc3E44XRu7+TE
ed4RJP30vGGhkY98MlQyTqPlrJKWtK1+RvvVBiEpiUOXEtny6a8Bk8nYTrai
yFQMVURXfcY+XZk7Ntybe+n34s5kMX3kKSvyg+ABccVNw5lVwCr/6WlLNSOI
J3A6hmTxyZL9p27+Iyey7WdVcR8mqKA6fhX3QgRQhHA86Ac0rP0cTT+3Z+93
RPDVRUwXBtfezPphqMjjjHz2OSJx8xzDwiYjPUUtfmDoz6/D+fjXPqK8fJGJ
vHBcr2JKtGgqplmideDJq3m3l10lDSM9vY+XMtohG2kw8tQzSHw8zqrNlZTT
EsehcKdzkcT7l+cTz28huzxqEjXQhW8Lpe0+F72kMmTboHILf9yLuIU5cw6b
WWSUm+X6hn/K6TPbDlXFdJUL66yF2mU+oJN46JRprSyDMatQP6W+3ikAZqHS
hhICQ/ptASL1bdcyGWez2W0YdSHXPoTSTg/NkeqGIPbhJonvSNU+1O6BLLxE
A0QGfJ1KfLiWAD/nhEd+ptM0vnbebovcqdrfospNY1UVe3tIkqzBFvliVYeK
NGov3D54Pi3TgtwnCMc6hsdP5oV5SjFXyzOXohK4SyoPFNIEYaNYjLw6r/Cn
X5Go0+rpBgOmweHVUwiPOnMJ7HnwKGWkTe3CmA0b/u0gPMnHDXt+UYNTWnif
XnDjeFkLVXj4fW45HvnuI4icYdhDu7noj4SA8up94Nm/XTDJ7ATzwoylPHvB
mQFKgk27un1MC40kWTXaxAeMWmmAyHrpVg1OehmiE1mP9YAKyuRVUP5bdbv8
qCa+sWMv4wVcn7V0BwKPBuh4Yg/FaOLK/6d8crKTlbe47/YQGweRGjB+jbDX
kUUuMm9KLU8JghMYHBp3ryDaJC9xrde/ZQ5MO56aGJ1/byisC7T4h+nLrrYa
mBdoi4fqThJiIXuPI0ZdybNL4z6z3GH6yy/6kA93yhQMtQpU7eLeH1x0QJ1N
Ngfzl2l/Ew2bApW4WAVEKrZlfJ56tT/89UEWJsFFjtfOkVcjX4INA/hzEpTd
4tk7JOZpV2ZR2tCigiD/l/nimFH0Nf6KuylVMfwoArLeVYJnAyqiPu/oOjrW
mk+fxIrH1+w8em3g6G1jgiIc1X5NRIvPMjSKYIR3EpiUymPoD9x83bvDXuOy
WshFj5sTNCbd/Fu/ehcTJuYtHVuaynUrVSjW58nCl0dxContSWqUokhGB/1A
uayctbD/Zb7Q5WKJjIzh9ACDxMmsf9JnyT8Xw5bUMwLo1JFbTqklk0ttYSyP
5gqrrgOAY/+J6ldKonNlkQ79QUJzTv78/mvMoLTI27VQPrwpUMoGPZxiamQ/
MqfMyoD+ObULYSY+K648uzu5sdhZ7TFUxoHQWpmKE2bwK86oYoT/7xy2oi0M
Rdg5kIr7HHpHpavhazEkbWbJA4Tj9dKzbNh+kjJp10rgDSw6NOjkXdedf8ah
Ir89pMme0HUcFJ1SWLfBROb0MXh9Udi0bZeaLVGoWn9vlnvrdTVKUHnR+4E9
TuHayYc2rvt2x/w3LVXtviw/M9p4sVd5LB8d2zeeG4v9xa4tzQny0doGx5UL
MuwdNIHjq0FcYmoQunvqx/Xstyeogt9KATp4Yxsjm5IiK5JXI7hdJAGi1ltB
zrAa2kRKOMFXu4obUwq4c7AWLoh9OR+j5wDVWty4vFW2jmhynkgRYJq77e8U
zFrLAaiJ0ZC4Qw/9IisNcNuLIzVufWiiVjI2iro4eqCNWLKE94Plz0zYCu6r
uwejc8pYPMRCEIgG8NGQEbBwB3Ru1E9jJtS2QQzXvlDGQWFdqlmnb3rBhcU5
ERcfL0Q5B6XE0c9vgvxQ7E1//GhGQrilXzgPGaL3UTNiJrkcFFZyxIusSJyC
ZlAu6XtTvx5DKbC1GvssZLGarf76ZzYutl/xDvTwiqIJeBsRE8vSEmGJVptu
yBYn4cFlb4mQ+1yYTHw2QktjhUpzx8+xp5i0+oI3M5KGsm0kcDnMN7xqOvQy
UXuXRIF5Hu03a+yOtm/DpuqjL24Xh6wfjYtJmHYGMEJjx02DbUPLpbGctui0
ouC16h/yO0q0qGoLwefnF/2ET6wavjGBYSibR6Q/J9ygecjUVnZtqG0CSUs0
1S8TwlIPZjC9CM0NY+muBBFNBlDoGl6io9oE4DnmRyqTnnZLhHhk+8G5j4Ka
05oHori4BYbn+9wROaa1vI1vXBkjxILdi54Fhx8cHn9ORdrZROXvKpoxJGjL
On4gh2pIJB9/nplI1ocAWhKDLM2a78KjcvXjtJKhdzQyN3DpEbU4cpYuJ/Gy
s9FbG2X/BuqEY94nvcCQbSYG4aP+rETP/s43Nmm2qerMUMz0VqULcd2nVjL8
Msr+n6HS6fA3toiNRvRjtpkpCwKpHXEb/Z4w+vnWHuspZrR3Hkx2XQoinYuQ
BwxmuZYtGDiBqovs1F/UDAv291ST2RWF0+uOJEHZlhZL1XAEVEVttRN9UlNq
ib4WWS+kyN7i01cZ8McXwOfadWO5A1SEqIcIpLvsb8Ga54ZXbUqYGYxaNVIT
rOpEuBHZOGMfArJkTpCgjnCsAZrHDO9L+jmh1zPtVP1MZucJr6N/oDtrbwLG
tM8MXFVU3ARKcX10ALYp5YczS7o3RmTh1kT10iIp9t9dVd4SRSkv2tNrHXS6
dDf0iU+XS0MZ8YMFXm0pl598gKduO9cXnsKy9iyW6wyf6GHxlSoiVTwjz1C/
EJ1dUnagL+D3GITfr/1fgM7RX91NkgSZYKjmLib7ZIYEXRZRuI3dsTyPBazv
bFEfANmgmoEl5X7EBquM0nc+yCKK+MLSt2M+0P+6tFVa8v9nqeflJHLYyJMj
1EWbMR6il47vAdHph6uHAqy5/s5aFlwqctkazBdOg+pg6bIIkocj4/zLNyVl
H3TZiqWWgRTuCTS0FAKRUJ9DiehFuD0T0i9yTI1wW6RusQQTLJNai9qxSEtG
iVhzf4EnUdX+rrIP7quIal+ybGbCn/JwPfkrahdi5vsPOfOAanVsOXrQ38dJ
VIwOaqOmxVf6I2zXIVZHTUxk7Vj4WXG2rBBZH2UImSQcGfo55hea2BHsrVSq
MtaNyzpP8QxKnyn2Q/SauvaNijIwExzzUgtOohpfo+QQHacXQz6CO+50SIth
A1RxBppe8zxRYtzoWlgo2xHo590hADOWovE4vS9gL28fVBqtd6F6leNJzZNY
aXc15R2LdRuwxnyxyWoTd8grB74yh769RV17eVQVqoDctadJcH3Z3DP+zlvW
xBPczUEPamg4lDht++VfqjZeCGA251L0afH9bKYQRoU7bql3RsKSpJ+wuzK4
xqKcT5fxIZRdIWMdzxDLBDAwuU7J6pTVRNsn/aTVqKTDru+Fi2CzhTRmgMJB
4VTZQPBSbpgXWora02C0MQQYZXuzuUKb9aNu8fceQEEg2kkp6IEu3bp/kgvh
UbykeZVCQZUcOSdKUyfN3D4xGdygkQCQjimzHCZC0UfsSSrUAazYdd7OHbVv
A8kB/kbBBKmXOVUI8Y1csdXIwgw7jvlPsoxA7FioPkkRTI4aKpRLMVir8yqA
eJR6pSWiuozFjeE//0h7am/+j9p31KQSsRQqr0vdEcqiGyDN6q6Wog1Ab9oD
Y5TjO7C6CjZ+KXoHmZuhL63Hgbz/Kuow/igW5SnoX+H2mXJ8rDpGuC/ipPFX
jkw6FEFuqkM2XtwGHIMvkEHXQrnq9ysJaGwcySILEvPNC9YHQ4tvlcnvWHz0
DK7QKoZWnsW/YRfX+L5RuRQxzocNCdoMGvHxGsqYZabfHTWQTQrDDlIeo160
nsbsRTpNynJhpBNxB+XNwcO2YMlXLYBP8Ofmx5gnQvePtiZOaKOFCWugnv6n
FuAVr2dJBK5E0ibKZRcnPw8ZgEazK1W8MvbPeIarvUYJszY4FUROSt4R8ntQ
YM+Tthjcwst4DKaccl/NtnjqRv9TCCunvwubGaDbZWrc9xV8ozHsyewkwvuK
4fjpk3NlM5JpFXDqbAeoruBQvijGYyC3EgZdEacK6GvMUpwTvbNkerc5Qy1u
CIa5Z72UEE7iaLVgy2/4JfRE05iNbUTTHBCNnlU00gLiX7Ml8i2X8+2ZQw+g
N+aZ/5ATMJyVDPAr5n1YdNE3pj6xWgXdmXyQrgqOUyp08R/L0nNsHOuFBicb
yidEV+npXeEgbCdOrEszt2s7lwweBVDFgDSnvnjyWBXVMotr/subA0ytXxKQ
VAwy+ApSDwzcqMxKUnMnu5oAPHWaV0NgSt55dPWYIz0AsRZHhW3H1Ys0b+fV
CfD/pI5lG+6seyIIi6amsBQ5ULelFjOnAX6A8UFragdiYAi6oIvFUIqH8aaa
y+z2cYoye7fncnBeoLJmYg+dSSxauoDOyai6y1+/Lt8EEyebq/6ZhlNg2/kB
qohjEkZPpq/MHg0+x4NUMlyCVQU5BfliZTmT1BxocJNzEc6chQdmSTVkdqhR
Fo5Fq3GvABJGh3876IbHSDqPMZzXT73VwVSZ6x4p0vNjlWgnjcipcLoD3XhU
9zi7PZN9N3gFJtFH9fB+Cc4GW9VjmoEkR+md5g/sFye5FEj+miLOzME8K2C6
2c34Cwc7EL3NflG6Dzu26jEENOV3ctKNwVoMcZPJ8BqKmoh6S6ht6veEoF6J
+u8LaA20eC88CCzW/qXZ2dtl0VQeduz7mic0iusJ/7rPuJAJJkWXqokoLXQV
k56M4eF8gBcEB7xB2MQZQ+EjcBNgqicRBtOZpJRkRtsqVLMGKqC/VFq/wyEC
HE87ORl0qHwuIt7WM2DTfrK1/RV/IW3p23F3dcRtUeGrkQk0z7RA/XPx/ZOb
R72LiQahZD3/YbkuUAGhIelYedGhISGLtgmbxsXv/kxEspHBV6uYcZfr1Tqe
pFwy//1+iSqvRDcyJHnhOdkImfyAKOhFhDBHV+uyOw+miHYgG23LTIpujWYW
KQCg1ROlf2+AL9dknsZWjhKpnyEfcV8MRXfNnu8auYPB2hGtMTLnA8BRCl7R
KHxQwblhw3wBzycYtcyPKg+Z7e5smBe5Kq3ZAu77BlEowE5XT8iSIv2MaOSv
gFx/vgdNGwYOe2d52ATTUsz1AKDxDYQ1E9ONghj4LqGm7mGyhCTIo9K1TddV
klXqXnIua07/kbaI4YdD7kdrMcy6cIws9Sm6bVFiKTuxNzYS2r0BqsMB/70k
Fdt9iylUiqHNRnRr4EbPgBS+7Tzy6IqTaotzLzxA5VJqEa26W8TeilBpKZd6
VTrDtHfOufKwMQcKmu/goGi7047fQcP0OMGdXIfPAamRjIk0eb3seuYFyc45
YTB+H/d69er3Kr3FfjLg/rovDDUSPN3OPT/4luB27hv/48UB4GcLce0r8/IR
G3FK5tybd+Z3jHeDcDR1g5W45sjaGrUQblBNUHOsJmYoe1E809sPP3D3y3gu
OCrPkvmOMwBurwRLHKfZwRs8CMMHroUPPWB3ugoP130pjvPc0TNXtFexwaD4
aDWyqAE1LHH7xpE9gvxYlfSK7ylJREWitGJcBqcTPBN7hzsbi+W6AXxeJz2X
byKI51QuCKDFDXP5RePsdxqdjD81cfcd5bC1LuWCSjuMAsIsyw57XyG7cE9e
aSwVDshjgGll6ir5m2K+yf5Z68sHI8flNP0IdwIPRs0Yv1RLUkdns0y0L5/o
PnN1w5RSISQJqBdgeR7af7WbGXpDpRPFCdVmtZ7zVPkQgAxdemP/tafRziVa
FSMnGHtpcoszQmeOkgs8K/cTd9tCW0mJz1VUki2N4mFc2jrT6JTkvZFWGJRF
eJ1nknpj//AMUdPxvxpl6S2a7qGLoSsdDDg6wm2G9aOtmvs7ku2xpz9/K2cT
v/KzH2Zp+V4OCGf9KSnx/ONFOEkxUH+x

`pragma protect end_protected
