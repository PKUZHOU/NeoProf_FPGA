// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WSlyXX5OZ51HxBrrIynYQo+SAG2qfO7sLowDI3Rmf01VjjPNNkpFGY+S20KC
WxCpSMhsmkex97GxsUlZVrdX8nkW6ty/ADNVkvQ2jRCnmPd3WbNg0VpXKcOB
gyaUUaOGFB1/RU3wSM4p6+/7VXXtj3nxSnlIApm4myt6M9PgkWNoViIYbZ3r
HoeNYznjiqpzeAtlVnHoz2KOR44BQmePCr6Cqjyf7uLAdWH9zt33aN/h9ay0
TKyYAboxmLI1NrY6KR9UjIC89lYVJiwQaa/lMHFPTBJwcidSqNnbbVHjaOFn
hNlbRVlGBokQi6A95J29KeiI+EtfQtfLxIqU9/fr2g==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
aD7Xz9Vep9RjsKSSLxzaf6IC73dyzjDZax6S64cqDC2yo2xhcgolTdw9lkze
Ech47QokallHzfE02uyi+0AdM1Y4vJG5GR6+8X2dr8y2PqvIqWt5WkjgQ3Dc
HjXBRUkwiPfMv8fjs5jHsBk17q0UxWpkOTsAXvMt3g/EFTaONew0BCiYEevS
12qPbC4Pb07jOtWzchets+53wkHBC0MruFZEQaA9OsuoLnxSO4FrMgDQMk2z
HG3+Z+H0JQ1XJ454iFeuOX0Z0ZY04olKo0iANxNxZ2jcBn3vmQMl5Wzt8yw3
WKqxbULvbRjYT+o8bEG1xfFnPBbozQ4wSh6J5KeyRQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
dtg6+UHW4JdqXlyKgr6hCWoIfTobOPfDcuzDsK97IloxDjqLaPFnFVDneahV
S22QKB0RNahfIol/e9zSrXrSQwXE7p5l2UCSHSdFqN1SGaeeEniCB/ioqZQe
7BYxZ/My1z42fZyMpNFOiUaIs/nurOHF4jgT7fpHbOxDnWbxFDQqlCrXlWVg
0lz2Q2e0DruzUySvbYYae0XwRdyrDSAv9mKamwZmcRvw77B840R1wq8UILpF
EQHc+e57OyvjV7IRCLLpnudX8xjSgWPYCCyd1w9TG4fUJC4iwYZnGCGi1HVJ
zrZVdj7RqUbQPjBqKwGNuG6pJOI1xsN1T8qZpCAcKQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
HBNZhXUdadqdpekLbDTFznc8SBKBjtmROBYPbF+TUY3htrvK0/njImmUnLre
a6ZAI8g7UHPtymHfj4Kp3/YoE6qGMJcUAZJC45XIvM3028VI9qSTKhNm+1Gr
Ub382a31Sl6lZWtOwqKVjSrHF4L1toTejFb5FQAwW7KSmcfw7Yg=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
AiuYBEWYevYFVTb6C/QBQLzyOKqIZsJFyarT08yfn1OTeIjApFJXd9LGI3wg
CeMmNnWaqx4XocYewaOZldFdf9ORjLJymXvnj/haa6UGUu2urPx1YmNfRfps
DHmzC6Z1gBDY2B1wOIRF+Gp5T2/2mIs2X8P0oruEUcs0azSFjSZnkVw83vRc
QydbA8TxqXYkDnsOjsM3QlidJmvSAZiEMfO8LqWWXtrsXBztOBtj3Y/VSZUi
kRG2jz2ENQWCyRLBpNM8tSfCzRftlo7JLzogdF75MEhe18r7gyhEF53XEQSq
9+ushVcXFY4RhBNjnBW7wK2hi9DPYJe6u5rEHb7euamCmcZGphNc5Pf+9/pl
h95j4rACWDiRtjAweeESh0Ui7YKui/Bgkw2tEHrmWCj3jQXjdRnumE5x3jrq
FTB4XTi7tkT1fiY144TPcszh6oG2c1gz85a791eXu3YdmyW30Qiu7IHJhyKm
zsxOPMbv9qiuVHObTTkbGWXMvSNlzk69


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
e0HnIogAYYOf3gPxSTRn28F71xqACgJ+QgdfIARPd6dRPMge6vOdtMZSHsHd
/GOwDi9gQOvR3TIjiZUDTyaLvNixdfp8KEebWOPJieGqHpvhB+rWGsfh8eEX
Y7PAHBSryGdD5pgpgpmMpwlUqO6UMa+ORvdz662Z5BOAIPjR5ds=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
MuNVqSUE3MFag8QNESbRgrz6ZM7R2+x/iU4jtwUIFaQqAdtxfRbu/S78Qmia
++g1kybTiLs2bHsUePDKvm9gKqazkPyDaynlnPYyTski3XKBNIP/7OsZBhhZ
k2WhD1un29CCbEFYzHvxvUfb0h1HTPJ5RniIXYRPFCemfr5NU68=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 15744)
`pragma protect data_block
JJeevUaoldDZQ69nfsliEYyOsZdrAUVFRo5kjQoCvN7NEeHr1Aq/amIz+iLN
T+Osf/GbXn5qOU6JtudadosZqzgmW8GNqWPnJm3U5W6gM5d5AAwXNI1hAtVr
pp4/D+aUCr2KBqapOiiBPEHIt9UqF+Rk4od0E+4TbKjt/NLvAAbP0SNNA00U
dK4CFQUXrKRKI/rnq6akV6klMKavn0V4JMimSloDUbZkVZ9pYnz9rgZXSeXp
0O9hGWCrY3kTBq1G2gbqwofGXe6O9l48nhurYC4sKLDd+H5IDz+K8CAaF+lS
lLOJdIjxJahW8beY64RYMHY/xWSu92DAPcInfy2Gn4uDsJhCOa6zKMtkCaWM
EcjBs/rb7S3SCayv3boJ4kKbaM5s1Z/kdXk6W/2sK9Nh+wS1Fyons7OfWhOZ
PX4RnmN2WHuiMFZ11VjKXIscwLuh46whDrQuEKJVUq1vPotGJUtpCZKVhUo0
px0VYzQXOHwV/XeGsZUEDyFIuTshPKd+rxD0n5DCZ9UesLHM3sW+HEQyS2XN
vUTwJl6Rn1wkccyBmK53QbPJ8TNllxsYRF2CyEZ7mCnCLAzO4UhiENwuS2jz
vEfBGPW2IWqdMIoqko8ts/yGvlzLdecE2T62X0UMFUa/Taa6ZNL/gKLDkNKV
MJ5/Gll+WO3lyf7zRYczgMw36/UG3PxDQdfTs70llFLtqtz8QXd72DcFzUq1
w/4tk/jeFi6Ro3PBcwyT9Asvi808xwmrV0rP4SNpNdpGRaUMVUKhqLUwTZ8o
RnlU76lZ+hTq5wknD6mZFqUF7eL2bE3Hktrrl350icRxq1wdJHernc0Zp5dO
FZXfE7aT/5G8nEbgHsOCSLiEhiBHjjV+l5r5lH6MySzkl6Hr4bpl99xucps5
zNc/iSORiMDrWYN18zrvk29HbW08/3jN8EMLXcn8vtoU7UbXMCVFTftvgOZm
1+/IDqjSIbE7wwTR3JIA326SooFb/ltfvBzmQZFIW10cXu+5mkt8naFxngDq
4L6JUvCl4ZfcN1ZVvtW4yY2uVobuD+3acwD9CePNbMgIFrrreVsCxTtWrcec
2vLo/0QlSarXdqXilIq99FsIXjkU52olShkfcjY7r8vyUphDWnuUnhPiGULd
Dgv2XBe111Ujf3ZtN9+r1bRvM6sb0s3RYcbypDuiJp3efSdWT7HZYUPgfOSm
bnAmZ0nR9wN/IynBMJntcv6S25K8vD1VkUrzFEJLtUVDmSWghGRY8TkiUIk8
7ShJQNixQ33AszcRduWFrcUzHdULeS6DPoCZWZLdj+CvKQdJLw1gMIi/DLgF
3YHMsrmDsWpSREnRo0Nh0yPPM8Vowikv7BZEQ76niXm3dnENV4ny+quFC0RZ
+5gq0165zb8xdRxrZMP5urjR42CmD3o+2ezSYxxnK04XvwuThLiQdLEvMnEQ
ysjiCxAL9yw0cKBs0/I++cRej7WWzGXDWjIsTmzYHkSSZKm0hdJXVF366wTl
yAkoZqdeR5MYiOxvwB5HlGdPf2rjtFvboP4gMpiyNuZAOFyyF+gMNQRmFc4C
G0lXZPLQ4JUL1QZs6MMXWqiE5E8Ha0/KzZCslzOkJ1PSeGXpzGru2nmDc426
z/GDkXViyJ2l8fZ8iqL1HLeZV2AjFx0UmMxPUSeXYyzUIkMgzpsvQCQeorNa
Uje3uEwEPMX0Lr83DaYRFtGGIVesQPNrhAc9C+edgP3f/ZNyl1kcGmoDPuOK
GeVvKrLBIjdsoE1IBvixN7vkHbNPJf/SrlAN8TsQ1JKfgyUCf2Gqd35cqgK3
7YYhkUrfjAsxR30uZqwu479QwXUukwBXQCjB+ZovQmwx3dSXCll4CZy8kMcy
UdZnnoFBtqgi3sIVRUNNgJ3LImPlMYvMlkyKqxr7WkstxqyAlOo2JvVhvkDn
1O7GJfBL8WY/gCeLl8FMyDelO8P9xXy5D4iOYkqCH24L1NlGtwGRkne93o/l
29fW2dJV5XRKp2FZ+NTRO48tMlRgX6MljgTwMVPz+cw3RRmq5f66rLXRO8oA
vleSWxAVx600QTqJw4ueDyjec+QguzN3dW0V6zdDI6qCOY6d0jb3vdZv8Fue
5lp5g9d6n6v66nuz8uBnd4oKWRXHalon7t1KEQWGf/DhkmJo4UhJd3gMiJoX
7IvXxbswNK3Y5KUjW3yz8xYfzva4KNMotOC39h0b4ZC9iMtV8XFL1InA7cNX
bxM1g3GFlee5hIe4bCUxR/30e6GtHokHzHI2kzpNmM0cWf7IMosYXVMaGUPZ
tRxVHoU7XJMAC/3oBUphgts0zCzfwp7954M7oTAtmowHI++D485gekOPBDsL
bMmBs6zwvxsKiYPCSLjLKEMxqehnRnu+4jVKHkPHoJ9zPTWPe6/W0UajpS0J
xMgTlCmyfq9ilBW8ntiorQvhYilnSoYeZenFG9zsrn8q0Rlh9sAAHmbp+zhG
qKt7mZT/4CoA0Au6y54XllApXM8NYZb1zLCGj3hIVGnixzsvpnNC2xH/KZmv
DAqwZvka0oGmEm+J/FgG9V2I4QAf/UIwUwdmfuSSe5iKFe7K3FilXMRsKI78
Nv+yjLzxCrNO8bKWnikSSRfz9kdQIwbrmG/Xk1ykX7QFDaQa7Q5ImDmRQqln
Sl5f7uBl0aANusszCAes6oefztAUDNjUX9SXEnrNpWbv0TYvs2Dr478hXz1U
IFGb0i6EmtIOa2kP48DjQ/S/mZl1lnm9d9spUQuCWus/yYspAZ0nC1o4x2pa
iFQenp0v63A34w2NS5HOCkojwUCdRpPd6cJUz960AXuOSQS7EYsYU7OEH8KR
xYd5Vmfyxz3xtttaAEqGTmLjpipjIVr/7mVy2EdDc5H5WLtUknt44rcGr8HD
EyXeJhsdqZUmCJhCELV6dSz6kHGoQZf1RGjIc/2UFPKjMLx4IXGyvDWbjOzZ
aknAoyptT7kj8LsNK8YOQNSDy7ivOPt2YaD60HMOtRm76kO/xesjC90001kp
8im9SH7YBWidOaxrdbn25LpKc+Q/BSegWWJ1RJy+Vx1x0nHUMyEyoZpqndlj
r6WHetajUQAa4uPjoyHg4UU6ccbLECsCTc3QGiO18A/RAEgN07d6NS8DwzCx
ED2y8OAKnyAtNTjPNTaBvoathdsxR1Yr/bobjeBZlFZFNg6S7qMRj3ZpqjUw
dmYz594aP2FdJOSto0qQR6c0ddxfuj1wlJB5hOeysXUSoBHXY+PzoPmioyzC
LjunGR8yC3BuvVFpnBfNHLTupCVRMe1OG5lnkRkCP3Estiufv/5slOGP6glE
PRTMd2ctyiVbiKnU0MyK+InuvNgxC1wnQLQfEzI8tOHGkT3nj/K3rBWVA0IQ
FLLTPfT1fRdIMkRjH2wb0gpAvVsG+BE+RI9LNRafxL5WPkx0GiDaT6zf5X0K
K1DA1U3xwkGlsbXQAG78+APpRv6KPP1Y5r1/eWi9pRLr8BmR55LMiT7TIyvo
Gtl5kEk0CokoyNXbF4gkc/bHnZ46vbh4+vDcI+TUY2JOeUq9Hd3lDShdhU59
cZUZzxqxXI0VYJgFsyRRe2O0ZYDIOWpMHLE907vNCiTjv79AiBUf6Mu8KUm/
VTuKNYJtKu7MgkXErtwrRCgZXbYI6asMa3mRuwuaMwlV4hGQXRR5nt3+VMIR
LOxioORKjOlJdNaJi0ptKo5J7hy5c6YJ7VBdY0cD4SOYlSerTROBi2KmgQWk
CQywX+826S/R1lKBUMwuEUJ+v0iVWBfr9WHy4jQnCbwKg47n4vICA4lFfHwX
ecqugbWcr2IedgY0BhC5bDJJisJLiROlVVUsqXgYw0/IlpfVerhptsnB3W77
t9cGiJGKL8MFdUQeVvinGP/lqBdfW59oQxc00WlPyghZZS0Sf7QPdU5AR0+l
H4cKVl3KXdiE47GTWCzQkpY/5h3rF2U+mBwNDn64oxIA9MkTTbZT8552OgwY
uxOZ0K3ehVoyO/3k7Y4NS7jslCH4VSFXsZMjLRGxzd7iHOKPQHuKUKz4ZW5b
d9jYq2Cqpz0KmqH5ArZu6maXp2aIR4eMgdv6Vx77NJD87ZaVi8LwM1YHi5XE
sAGG9ACm1P1KzhN+gYh+LgHpaFyo4JroKKod/wSIgJwhaUSUCHmTwqnFLlP0
maWTZXAA+W4vpGO9iOA/693U9Q1+R48on+1sEGkIuIymElsSZesCJTyYL0sj
6xgfXf+7K7x+KLe+bBpMsRgvxQyH0wdneuuDKXSuYtV+bvgqXwHKemULCBIJ
RNXZUAcJ22guo7oZKmy2xU/5xfWOv+/VBb0KocqyrTh03IFsMx9CdNaB25py
8tNt+T9jHLwe1KPY+DqeZaBBON30dqnz+cmRqHYGFS9Zl2OWW39QeRrJIn13
jUCCCssZ2WA5aKgt2jvJPQHyUmJ3abygigawf8kHg2TJAWT7D3Qmwrqb8mKp
g4qbhH7yr5xWwxAs/8e8qLw67v4z3tyqWzFVj0xqYUV2sIaL/7rkv+Y+TMX3
Myb28sHd3/VB31NT2q6k3ElgtxT/Qp942QWk/d2j8RR0eQH73q/QQKGxhMvN
hbUOq4eznhOwKdwfHHxyP5F3HOQO6zqaYLZwYb8wK05bTTHxA1D6JHcykDtS
pzwK/lHTdnrL0BhucX4m4r4qr5/k8IXNJiJyoShkmKA7tyrwRe5OzOXWKRTK
4F9JNkZky4RhZoyhBUJ3/lJagCYZWW+hEbRt4mktzanF5J+/QlRjI/gC1E0U
V4uxNoPhxcliTzB95nrFvgVRMz7WADGKd00kDBHjjF0U7HUoO1MiStC0NC0z
ZgJoKZfyk5yXhHf82liN6gjlFoO0tBllCstBOVRFIw1Xtb5VRxX39CbdvIek
U0H6mU/1aOjywEBdLvIsXE8U+aBbBBt0V6S7t+f/pxuoaY9q/wh+zvpdpor0
9JzZwUgU144wAJ5rV6muKqkLvB7HOteX0lqIzNPcj13F0sqNgyqgHTGP22nP
I3Cef/kwcd1oDZJv2WKFb+1rPoBGZM40tYJlfJh9TzusKUR2vQv/JfUO7qcS
DvVfZTM9HQTgOnU2ANReD0e4FhcrM8dW5k1XefeWenMJ37iooElJU0kstE0L
l0hBWrKgurShebhyBZEIbdvfjwACIzDQHXBHQkcqBbvTHF2NGZ9AZaKhuWyb
KGaM0rANesiFeJbTzZ9ONIYMOsc/WbRqCo8hHynOedToy3OtYDL1O2sQ51DW
3c66HRuyFCc+dUt+JAq5A7vi01qrFlt4j8sTUA+hnbE3XiRlGGIEI6r9ryf1
BqCEJz1CqypoBX/MstimqoLTXsRLxmyv+adWTz+E0FfQb7JRjyFvziHulm8N
nbMx+SUJR2iXrOFsDOrhLtUcI/Cjh1miBFFqGxN4p44650JT2gtGJvHf0dre
+Qi1woRaM38MnF7tyjWnAenX/ftTBmfQcG4AVjTDyzsY4K8dUPEEUe7ugnN2
uSzvFt0WGJm4v13tcVjKw/0wgkKf59vjbp3CCZI9mMgg/RvfFEjAgPqQ4MXU
z5f1EOAJwuuD6ZOus1oYL0/EFnrNwO5nOFwQHDWMKj6qrkgKJ1zPcHRUfyuq
V7IJBR1STlH2FRCDRe5gEzU7NQma2n9gcfqUvj2aaICeI6xsX1rnJIDGsIPJ
cL3KJlG/fmzem84g7aj7wmBdsFJK1xiuxOVrI/TdN5Io/alCc4eNzlaeEY3P
xpSxqDgC2N6+Rx5W5wVvIJrzWOio1QbdKa0J2VoHh+GcxJwYcshhvc7AOGRx
cjtT6bSHz/ioa6+GO6aHUklHnr1/J+14KROy+/sMADn7KiD26yuz6JXhRuyy
lzX+lHXyOaCGWaI+BFJn9fTIASAf2+vUTdHCxxk38Oubm/FbWupPDNwPAERP
beiVCEmRtBhpb3TI//QzjwXrwAD1BYtBaiAc8Z3GGD+gR8Bzme72Hsszkoy8
41HQ+uztDaXOy0V2ADREqMBmt5BFzB12SCFr25eAIwjLhKtCIrefJWlqOdfD
6JiGkRTG10ESaeuXYTiiy2iicFfiiGzh3dzz+YOmytLpfHQyQEw5dRpM4qhG
9/4SQPItCqeMyv7w9jJT4AxLUdab/it8jnSf4NZ4cdox2Dd+dTjM6xQXCXe9
mDDFujX9Dg6B5vvykGmnf23yKQ1MGm2fbmE63COX0gvqxgX6m9k4QWnl/iUz
nLipKFKkxzTQnayPpwtZIl8nvJAWEjdwteEgeZ4oiWQ41ulnb+hqKZhBIkwd
4hoyah/nHzDRJ1D6OEflJ3wVZGZRrAbs2Nwr5rHs4U8Dkl4sWmP8t0eX8MMO
WC2YaejWTUP+7MMfhLWsDk289y+UjWTJO5SdPECmQ6LoXZHwcsbDvMkNpiX7
B4hJvxVzZ+wmFlOC4FCkAUaEiVvpI928GM7yWUvYjYTZinOUNqEKOgER+88X
Cnv4RuCsIrWLOAHc4xj8OpWfZRzgdvBmzpNEpGzzbcoSYg/yiVx2BOZXxHGQ
KA1kqoD4ldFup8RTQdRJDvple6+mer1mSawqlr9s82zXzdAnUoMo8dhbTPFD
DF1a4tggR8M6Cixr589ucMXaerJf/EmI3cbYZSM5xgt6KUPAf5wFEhtW+s1Z
OSx1FIxL01o6wRZgFEVY8RXUZVG9uKPlTBEDUoDTiz56LPiprb2R1obb4oKq
+gxt1A/dFr9HpVlLjZYITcTCBGXibnE8eKlCvGndolvBP3N3ocwd9s09U5MW
Dk0dufncj4l07zumUrCp0ZurDKex9pd15rDXJCa6CjJjUgjY0sM2P8KmByVi
CYuplbL1+6VXuGOTknfxDcsw2xXDTF4aQZ3czB1ltu5JThLTfGB41qQAPJ8S
ErdPRnso5xXMmT+dcJ9fjrKGaAvn75YtZ1vDmxOgtFp2cSOZbZmTcVkJR3iW
kCL9HVzZjdjKR6WOqD5X0RyLJPpQbuvxSuIAZninoPdfSarsDJ0isA+Yk9+y
9OnYvS3xmpJg2yJhhuO1eTumEmjc+hV6M6vdQUENTF/UNDNJnfva8VB6etAl
DD5nw9pUaJ65cwHXZ/yf3YiaGwjPQPWrP311Frx994KpWoUG/s9VtYYxjy8L
XSoarYodJvS0rYVKxIyr11/4nTi7kKW9rQwVendx9277DZJJX1ZlADg5H/5T
wngdD0EqynCQVlzYPquojUtYX6Y5S6V1M+WLhkJN5ukNXhbfOcrv+8S53tSh
uZdv92HKswtXY+F5H1qhvmqkq1mHipDyE16Xf5gegO4YlxjMr7/Moe+KN4p/
UDuicQOWBf0+sd9NteO4sfihHrxD//iE19b+jp5GJ1eA2yD/BSHzeFfwjGgA
dhfPtBOcnJ2O7kEANECdE2KLlCeyAKpWGm6kRq/xk3oW5KYEnMbta8GwEBV0
Z7MBlr9eIG4baj8udbgG0l6Nbq6FzZe6F7sF06NczHbdEgnG3JFCXZou9gMh
5ClVv5ccMTbjJIWOTtUCUwfC7modF8KYD1nvgMZdn0/5cDnjpv+uMlh9Ik8s
W3a+HvrWUNiNU8hNUqxWYGq5qJmz1haXHjNnY4JG5SEwtnusb4bwyrvkJvzl
cuuvccMFrwQxapTrNuWFZkkQqtX8DEgHugx6knfau99ZTXOM5PgqA4iAm2+B
W6xjmIuomuZNqRsJTiVlWEYO8ivkVgTD82v/fBiv4Agho/LAs1yR6l4TPoTw
z3L8Oe1M0W5DTyfMjI41qAMLzeP/jaWn+CKB4Vb3Bc7nZ6bh5a5fBX/Sg3AP
uvZASqfbtJqRValIVAxcHvHX1RocFUY+e6tgJ0XdDUinUHx9OzeVeqay1QWo
aVkDvrru77BZ7gwb59BC2gz9Jr76qYWNEKXULJA2uhclnNsEYkQVA2X/rW/b
gnZ1P2bf2e0p85+tL/XGYBB9M7P6y5Ok8sbUrdVF9peiCaDViKU2xsWs01Zk
4mmlWVVYg1Q6STW0uLwwimpLGIv1DJO0jWrWtgXvGtcSQ0fnXXMOfXCvawbF
n2EGwqu/p+eTatCcocrzlC1lsLaUycaNGeYmqoa/CtZ/0vPKkYPLgijS7HCW
GwZkBLw3Pqnxnqc77nRqSlYFLMiyJ8CWol4sYuf4gbzm5YArXu8ZAPyC4TxO
rNQP7LWMPU9Kz7x9HZnawIHs3nu8OHz7VFAJqh0+p9hzGh73uV/SnriiK/qk
QxY2dtY+cuqk184ZhWWvYbyJ9As9FklwFqYY4+sUz2h5xbAq8uX3HeqAeirf
+CciDQ1jsGMyZ1OVJMamI/1EwReowAwMo7HlfuIylmiDcrFacQYqAKfz1kpz
nmq2H5t9BbX3mwnHDDVSLwDHBYIZcRCZYFNAk3WdBh+CIF8DfZ3Kr+A5T3Fm
gJ68y1R06FaJAI/mhn+MDbAD2etvr0OGfjx4sEq9MhOsHFQxdboYleDXNnNL
lMRATl8xcQ2ihtNuO75wDJ8sYxNVDx/f0MucfUsSETbExgSIVvgXlsj8zfS8
53rJXsQaNHmSfg8Tp9YRddIz/lqGqP3CdyJpuaXT7v4Q9UT3BwNxHexpIE+m
OX2R4uEhEOGWwKBC9eHUBC7OSnA/YvTQg7SdXv7bQ2UjocY2kPxG+/c+0jsT
jpE7eYM6hhDLroDaVaqVc6uqg7de5sqy2WPCx0oCPtV3QCjihP+m2KFwR6FW
Hbi0HXmAx+2+WVXdK7xMVLcj60SArgmEJr4vlUFghZ+7kX5hHourHI6CFG7V
0fCJSAoyQDGaTN/etjrHYRTT7jgxe0xNzRooXf5DV29eeUYXDBNgYYwZCsDs
sD3qDYlzSj0wljG/ffuEGm+8/BsvzTcoI/y1yBFZmRlG8OHIaU+GUCVnI+cx
ncRmfR6Il0SvqrP2Zm/B7Otqgd3qfofaNVvVPPTFZbPi/bRJokMYstI9lgQ/
zxgWyTpSV9Qt1BKVni2THJR5Zg2PNZ5W5d7O23oApLYkTcnZsz/yNmuHJXPg
v/4uS6safpzjmrqbTJ3KBkXhF9Q6a2q3UHo03SnIOi+lLmZgw7dNQwP9/vyW
I0fgg8xo2crT+pwkS/3T+bP7phgXW8wYAN2sgVTj0zJxoCaBf6DJjE/KzvSR
8VVOCgwO11WozZR5Ir9X/FR1w0yc07W4w1rkTBA1ByraOXQN/Tc5YZr61o5c
LUtRtxbruVLiVQvYvAK4XiHIKbIVJh6hzkkxye5U4lWea3c81XtxEmcBLR8h
+rS9qzzVce6Gj7iDqs7IVJE+2CHj5EyfgW4ytY8BzrGDYOBH9CbNchDTe3U8
dLEeJC/XukPtxJv8XI2BMhCAhIalN6sYDVsE9bzBD+uYnPRWl7I7j504i8C+
sywBqa56JzvVhu2x+2UVLv8SzT/v7UqtadZp80tBQNHS50hzXRBnGk56FnP4
7xg/eUjQ9NJxD/1fF+q4Ll8eedzZEpXyEfosqHK6RoiE9vwloMDTL2Voy4ic
TsykXvVeZ9ux4vOy2Ah6zNkZfXrlg4zG+MCWuuMepvKT9upVvcw4k5VPFxO5
DuopdZSyCtPtozMxhPitXyO1k4q+1WwU1MCRIHfbGAerZqI/TAXhnM2xEZg5
fB1gVcn6DYAOU/nUGjn8GMon0XGrpGtY8jRWyE1GZqE1BHUTswb1hYt118Px
arNmkg1+X7M4ztYIXO+vu6r0snLzEbS5HXXPF+Q507dHhmqvkA1x+KwNCJ0A
xD5lBQmeqEmT5SPXI63ue9+DiACSOGdUIcS/lU5B8Sh3nokcvUbmX3x9rhAZ
/kYyOjU0acZoBfhdwt2rQgvX6TUovNCOAnr/XZF+n+e76fwylBmPt+VhF9+S
5PV1MPNmgJNoNgIRzV8zwHBkivRc1KT/cbd8hxj5e2HPt2nF9l2txLrhLRRL
syB1RoG64CWRRotpiJhGCUJeHenKo8Y5su11+SItMi3nOD/0fOEudfai0KVN
sfjxQTe/DA2GqzvccBdXQhFBjbslAKpdChgEV1NsUA5jrZrLfmWJ+wuaB5cF
IPZ7fkClwyZIbaR5+9A6Jg39qX/22usaDuHpY/hIHV2xCf9TIT+t8agatpfD
z2KC49UoaiZ8eOu41ICBM2H1QPikpNLNv7cXNOaJTlNoxV2r5ckdJEkS6dH7
96h4duKIMc0O8zk8yBVfadNa9BSyWo0vKw1syrcNKJ9Vkj9EUCWrAYQeuw7Z
Bw0/WIMvqnAw5gZxM4Py8LFchTxZwqP06hWSv2tO217LBAVeqY1YC5hMkzS5
O81j/A6I+UW0KOmwc5DBT+Kd/Zh8ZRivuf9PI43m9x7EyYT2WVThAuUnJhIn
MWxPKm/HJDnm+yd8WTRJNnfdRZ4aPdRrepxH8pFbzesDZM8UiIfdMMAJ74Nc
LzkEjckNIIlveBmplwl12zkKA0br0w9EkZcBDLWMqSJN281yh0LrPt/zDPNY
+WJTtEs1bY2jqfV9e/zJMyOSy3VuBnihwhVnNDdrdN0fEsRX4DdgD2mH2A/f
38bKqdc5iVaVn+e6HSXFCpuFwL/pXzegnTohEOMPfTVvqUmj9ucWj1xsVqck
2lUatbOocbQSFYpLLDmTm+Nzu0sThNrTZYAWKHXkyj4gMKxiFRHlanHgriWo
j20SjfqMgFvRYA0kkZkH+0HJwa/ado52nwrnGpdp+PvvsqlDIueRXvv7LN3t
Ec/Uv+yRdDtyf2m8SjkECvIY3N3oC03q4Cq8apdNmvYdjBsdVVtj2aim3qu9
wVGkWjXVSBg0um52eq/Tri8sQlrtCrocN9GNSM8vUtOimN8sTEuzvTQrC5ea
+e5IBhPQW3EGbtpOSDX4AzEx3viOd2+EROtHRll2vrlyok2zaNOJtSGv88Pl
BI4Z4tovAo/fe+t+nLyLCF9CdIa7D6HWIpl6b+tU9024UPlsgymhC/eAv6K2
lYhcBtgQy9BjH1t/gyz10DCpAsA+/4kE5L8LrEpW40llv9xatz0Et14eKhp9
QINNy8/V4rd0a81r9N/h+pEAPgbwpcOxLhjpcThZ42K/XP929HiZHiETQsmR
WQkDDpKcjYZ813bFP0KgxwJbYDNOtvNHWUzNjxuYU/bzSV7FUf6mfdd6JnuI
1MXRvX+GrhY1zrYa7cQ4fNsh9MqsXzN87X/PSKhpnm9w7LF6jWB5qVOd8dnE
pTJxXwMvoF57Lw+PZ7DmCexy5IyuCguuvGdxxVAmawHIcz8NJPzPs6luG8Ny
2BCyIhMCXc7eHNpjCjx0H/j8JBFoFug5gndeNRkOKtHVgLbP6zZHJLUGBAdP
FvRe9c+2IoEqxqxtd+GDOEtCOFWQobiSfG6yxpuAFiGzI+pDRY3OApzq0er9
QG2hiqXNW+z0/x1QmX/pWpAOo8TxyvWEZSm91JtZZG+TB+/5eSOA9KTNULys
XzwIuLsErZ2erlhudHz9ML5WpDligQzN2UmT5bT/GAYwvEPu9ZDkEgN4itdT
r11Ov10hGvx0PFsJYd41BcO6/qXCDTDBT1pl5QYAt/PDyOEP8/C8lvfSj4Wx
8CZr6k7lnzI+8fy0ZRHzSq84ki0vkit72eqXD6ugoUCihQkAPYrPbk4hIYyN
kFdW5B3QBOnEqM4tTs0ep00+3ySJvGtb51MPPfz1tI2bGqmqNk/KaTupNqsK
q6g6AhQEDeG3F32cQtVoPPbODol4bbLlnxZixhYHvNI9cAtzUQPgLCOPoEQr
ReqMB2kvq3/G5jKSnJW6GXgajzyrsBy0gDtbSSl59RhMK9nrwybtoUpoNSJT
lbgCg9dTQjLDPBR1RMQCweDdOrnuILqKy4f23/OISPGx1/S3Q4jdpolW8YBF
h88Gen2ZYSLKPSMDCJql9TNlwaJWQFWJFlDr1UC+X5yyawClILM+xYXZapm2
BmEiYunA1o+zCYCnyR9WXg1zSQ+U21PGoa/yVer90cDrCjTLr0xzPaCxZ97J
hPUMcEX3SNNBZqXtybFhm56ebfPCdu2Dzq9+r/CgDpgO0lkrQc/+xUrtyohY
dwW+NChyDr8YN8PaIkPFpWSjqVBpe3Z0wQ+G1bg5MIHGSZe/mXekFLyodDeg
qpGQ5N4fz9Os9F8kk+Zog5lZfkMAsJef+PEf3UzyNSPEsTOIVRAqST+0mOAw
TAnUDKCqEBHtdywZeEmonTMBA/wlLpcH6JtX5ZnrEZWIXTyZ1sjCc3xpDa8C
UW9hfQ0yg+Z01x3oB3KxrtdW86DTqJwR28TwRrJ3Su0cmadQeWuE1D8i5IHd
kqyULwbg5lHrcZp/vjv31HcYZA5cZVFwwl8nfxVGAGLHvfL1xlW9qJxiBPUh
vZqwd5ATQi5ZKokgAgjwykNpDIYYC69qPGKDmlYppG7qUA/fYr3OV9QNs8Vj
VcXvPVx8aIgFISwu9cTyYhsIu1ksicwpF9a38w48gsYH0OsXwvplgt1Gb6RI
qpeR8rR5N37jSu5LoR0s6oxQmWdwugrAWKXvQy3dAp0JfpVac/5alzJb3R/E
0kLq2fRPIu56wD7vJ/00tbpZIDGwxOFKQuW7MfMF3nXidzkgp5vbn9w8OOaJ
/A58JIkZTUsY0Ck5FVjfN82kuO8JHJqjdg+/okTb9m7TrpvZrIAXQ1Jo+cQx
09K95ZWfBkTu/wsZIJoia1YVBDvqvKhzb/HVLFc3EwKn5HP4NJjFESGB4WHE
DCt58HJCTW3KbJLa1k4EHnuNf0vVf5CEwW1cZ6gCEXoi9EnXuMq3mCMKxaJf
smxyPcoEKlUE3j6ows7o0QlbrdBmlErT68I8YiTG5Y3oSEytjO8kGbasRGZt
ByCmYS8uCZ4cueHXTtbpijOZmxmrtVp1vvb6YLR5DxL7kAiNCwK/JXc6LU88
afdmb7IIyefxBJ8/Y+6nHIboJ4vgaa7ODJ+p8qGhB3H9dctDoVzJPHYaMnzW
m5IkeVFnxaOLA/8zuA5p2i6b82AoS4uTb+NHgdvSLIUYUtk1YiJVByxmVYa+
kor366pMM79Ks5Zr8T4aAFMQ+uuh0FX9ffDJXke5hMnq1x8RsZ7slSlmRNzj
mt69aDe+h8kA2zcCrYaf9M3XRQtC05zehOWnMf+fz9/XHs823ktd8etdopwf
nf+A55DqeZJK88krc5xKYhKxRMNMzYoY8vyo2zSUJcyeiE+duDlKaQ9zEeQA
VHIalyiHabytLBfIJNjoqtDEovawN9ufqo7nG7UVueQWb/dOmG7gNazjl+5+
OPg7Qj3Payjeq1A0Ppq/kCU/mM5VsgoovxGLUT2Yzu+4cWB0SLfBglzw9c30
fQWmHKUM0O0VUAwM8cufddaZJKUPve7Zz6dBToAAAw+ORWFz6NK2hFH43G0o
j0cAvth5CAMuvrMyuKxGUltYQ9y4D8OjH2YM1ts2zMdsnxWmnK0Jmk8uYdHZ
DlMkSGWEg0n1xxOJtqw5s2mwpsRJcUJ+HdowbHNb/mNfw303QYYhbaRm2Tx9
542oWW1qmqS/m9Y1CJsLVZbIQqojX59XPRcmhMtLQ9ek41b2pmYQsNj+dYtL
vah7D7a2hX0C9Ln7wn5JgG4KhP+qP8YDLC+65MJY3YhOCeGDhscMsAsTggcQ
HHx62DovnjG4GVePjLheoc2O0HUw7qwG1VyRXUXqarlOedlEzTbKO6KzPucb
VIDRUhBxoluKSnaMUQjsNNmwrRvqv31N68nGm/DkHRgTxLiVPpMNXvBqYQcI
0Gj7B7wGhBpF7+NMCvrKl5Sjx0cm+yIU0E/S7Jr02XLIz2goDBS0XA3fYnsm
Y7+FIRBSdrBLtLm9bo06n6k5ZQVFl0rngH7HG3nPprv3zmNhEdVbQ1kEqxLS
aG7z6qT6vpp0LfL5aOPo7MvsHozrzLoNh9TpFwpBNpCvsU8A1mh5cNMAvSWx
/rxQGUSey1SWpWu3/m++WPNy3qf1r2K1kSA4XNki3WGdlKKbG6nqI3OrQ6EK
SF+vI9+Ceh2QD1OSrQQ75HqlbUG8bFnzXLln1JAfSg7reXjXLAHmen/5ES/H
5DkBJmfTa8IzCAScZVABEsrNHzkMLLdNYyVmCBU5T+Vql32almHdPaDqwyRa
Qc930ohjUnz8gSq34nNPqilLCLi4PuhE509J00oRgMoNDYORO8rJ33ciMFbx
0P+eFeimbkEz0EFw1LSo9hEc7Eg8i1Rl/GaS5R8cMA7DNqrRBdFSl5PmBqEh
nx36vNwgU9DB/eX7pshu2ZwNTxCLcqefeFeOMXHM8CZbHU/rUKbFoFIWjkYm
Vlytm8eKgWa4dNTZ85eQl3uUAwkwkV+2o3E8qjZtlI/3QiTzm7KLS6Fzy39w
QkOzLN+bP44XO/rueQcY/8iEhSqfI99pn9/mRHbJtGjJW65VTNjbWtYQReyE
p+K35co2E5NvdnbD+XNHGqw/WMROdu++dxID4+Hpjq1jHTXycCCrRv5OROXE
3v2373DG+q7d5J2oFxn6ImURFhjolQKLgldk1Ic8ow1CxgmFd4mgom4cWNHs
8lxSIMVFwy2zDsTKahk5FEWZdiJvTORqpYVvCKMe9yZWqaHzME+AG2uDFYZE
Mo2vTqrPIdbCGBQyvgGHPyJcYXht2PRl5QFZ9tRlGdauPNnoEOgujjgzvI52
VHnCDETGjBiV5CcPpTjd0QqOWjGsNCMww7mxgNjmwHYjnxEdqmj5C/MjFhmV
uvgN+/KlwG/P4vYTE5ei5uIm8mDO8mhSDSjlEjOMzT0KzQX9/C9WHj6ZcOh6
lwF4FVGCsVPkF3rHAeFeYeNvON+MN2+Ymj7WfDf4IuhxCwAdF9z05eV/dR04
AIGd3QxuHIb6ZpoZs7vq5ZGegjttIKKO9wbS/47WgLavzIE/ZXx9OxOQ1/1U
IJDS7JhcfKnIN9piCWRG6Jhp4itbClRgrka2sOD5JKs459FC329hQNZH7tjY
zPSsR4myDYv5MP7dju97or36TbgCEhKTGOpMv5QlGRB1X9b8mNrUtcbw5nFy
ZnatCvDMJupkYp10jR+dsPZYZRrzrPEY+Z1M+ERyA8TDtEGGe2xUYNetFxBV
ZVaATQnbQA0ZPom7e662TAtGmdd9cjnCjb6TuA67pfc2f9KZjAGlVh4zVGYT
zB3FmegzDhnXjBmifnkvnjyrhbrvJNu7tGlF/FLdEFOJ329P985E5RleHsy3
4Hed8shiz5jNEDmkd9dDjeR7JJTnKNgwhHTuk/6vwg2t+iP7iLYX/6BQziu/
/1js4jyCpD3a8eiq37jJoi+Ee8ZyD1/YDK7AtD9onYpr56M3oj+hYm0nEtc5
HglLWsSMHsbn9OfUH76NqjSeHtjWRAn2BEoQ9kNgxh1yD50lkrGC0AxOvwvp
SZtc1kS04nxWds6kcFD06RIArFJdF6XUCu2btozajbmrtNVtD//+KtAQcQSs
WsXhgVhEEqEnIB0xyyHGW+uMeDYiFCXjSO0BpoZiCKRAWgAZrWdwvX/WDEKY
2zHx4na3lDAmNHwn0842pOHarLTnoaeQQTYGcLIXpNJ3mf1+2CRmKIX0xmAT
5u0kfr5LuXW/6YXOtg3E59E6hWXS1Tb2q2xjD8QeKdbg0DUzhYCN2MVrvF1t
9MaT0lOwwLlZ1Z7RMPtaIq/6zK309rkJNjDgqhHdbxUmWVVqhJG1FOEjtQZx
+9li6mYn/6+BYCYiuK6qehjnSGHAJN0mgIkP55sV8x/3RE/oT35yEiay/Rxr
QhuiDA9UmDojH9Tzg8ladn/7+mISKmN8yGSiYmpLBAWqRD0fCce7mz9AZkJY
82bsqKiCSDtpBXP6CqhhTMogNj1HH1IpDzhEbV22kFhIQn+waUxc18b7JF8d
7MAoS0aEuMG4fbq3FiWzbFM2Xhk6vvYpO6NpI8+A6YNPBKkViFyDKNqAKIa6
oXDkM1f7OiI5uzMQV1lMmJhFmsaBeipkvAFX9Zr5g21KA0dxqgDr9g1ORtaS
VutMrAQ7nrX3XhFm5eMcJ6WsQ/K9DTv3TEwGLuB8I1TnDIiewbVwqWmVoOZk
+E1qYQUkkoPMQqlOGosI1Cayt1gZgR79rzbcTTnxQ19JJiRU2Mq3A8XUpdpK
CUEU0cSDeyyF6C0WOMg4cjdpz6MRvIELPfeIlqisahIM9lbhIQ2dcd5xmNqW
4SktUQocYli9mejkgoyQK7xSCpj2F9H/SFLIkNUOituUWMzqTM225V6KE2oC
mijXLo5pIAXxLdJzAmIbeYP3qbaZ4yeS984Vd/OJMY2FJ+KLg3hZ3TIqrsvD
GkAIqcUIgS+orrH76napw+Qy1iU2WfaqyW/GacV4dq6cTZX2oOhdiLg/HkoV
/jzemMT1KxHoBe64t7DjK4447M05AsJMt7U2h9bb03dx9doJ9+p7lEHln7Bl
3ritpqhixyMgY/lTSpK6pbSV0m83RlwCKiU8DGu7V4xAakRvUAdz7kNPjYUS
M9ZqS6KdPDNWRogKr2l/bEnRUqOrViUx9hJgIg0++XajVKlVVL3qyH++fgSj
KhdHXZZItmaFhZI1gYKmkd716MSiX9sKPGk+XZAcuHOQbc9xwqYZJ9er6D8x
Fow3FmciMCTkttkJl0AddkqZFlvjhOUHISY2W3lyt7WqMNFkqYVAB1NkZLQ2
EmjdwAMoJU2+OT2TUzS/jOFzjmcpg8xMG8JhbWjmQoSaVvOoTUMkqOMwRLZi
WBWnk1yhVCdo985ALKkIjB9UakdvIdhONju+AVpVaFSDonnascLwmtuA18hW
csO/4+V28TAdL7t2aUQxkT31QFrWEpqL0W6KEnKhQN4ZJSL24KJRmdB0aRBl
Z9YVZ/zUGa2V7zPbTDvmvpbVGYBxiPM4iUxDe0I1HmgnbXaKE5bNOrDFnXo0
PHmqC9tocZcTOjUx7Q+hyxPsTwS/qHs5oNb1XZG2OWql1QPFJJYow/l78Fp0
2xisE25YuYSYJh+B9xgpGvKRdnmul466PfX3GL6sQo6FQvIWSGkyKm2SXPXL
12TtvZwtrLl57WFmN2pfI8ES4UWzSlfhJZ+lo7RALZQdGf8gGfiDgjxrxb6x
zR8Rpb6lGgbQpIy5eh9DyPX7UOWHV1rNj/wisLv57tmpNt1Vo2Z+P8zfhoC9
g/i2GHCsayg21Lt7upq0VyzDwR83oIlpDfCRqLvZy+nxN0MlsO9p6VJixchE
M97CirO58YeVgABjpeNzbVI8Xoz2vXk0GoTQuOURROFC6jOt9LFQDq+QwGyp
dIfowo26bardz1B3+aPQDHTZXAjtqkloiVNIiICxQIpDOOpBlNfdp3xw9Svh
XiyPGP9+62hGt2TyghR4A4cSnxAwrHEi0+gYA29lEzogqzX8H0rgnftJTHax
WqMLt/1+/V8C67JbuE7r+JE88OjuXfO3EC4PxXdqMCt2BAm3BvdU0lxPMI3P
VQ6F1ambrXcFWPOXsAvLfcCrgS2F0M9KXYL6HceT2v6zwu6Xd5gUgPg6oLVF
h9PtSCu5272Oypvk2jX2CZgNiCT1knxS81cxvc28o2PFB/LKIkL1S5i0Gye7
GhdzSR11f4XW+WurvdxE1GBH1CQ1PqnZ2Msq6kUVhjsjAmCQQZJvH+3F3dAe
j3GDsdoidQbUrBRq2ixb2RpoBwelICpsMczyRdprbkVuMqpv6afgsS85k+/O
C5z+D+84mz37sMvADK4ONeKOM73CjuRKUO4+UTtt3f4inTjiefo8/o45R9b8
aaWYdKh7U7+h9aJRma43WSHKiOlUd74yLgwy13zzdfNTUOqCF9Bf0mVVdgWc
p3Hd7mCqYNstCbBFrkavboQD8wJ4OjD1CfukAQiQD4ldyZ/LfDuKHNI3Cqn8
RCChHwNysa8sNTwT0GXt9eur2aOu1KNWOHWszQcOGifmSTuPmYaFD+/DLDe7
h9HKwThd+1NESp5JIStYVdhi0wOuaCq+nOtyyrFwSo5wsH5+YuGLzuppXo45
6mEyQEKre1L7mCmkVpZe2PTO6MN99aqRvDsBe28mrt/cww/bzyOgjFBO7DSg
h57N7LeoS8NIzs+fHNsBsH1C0bJwcPAmjsLR1QeWd/gNnY7iFDahM3OjbraD
Rsc6npD9/M91+NNV8drH3xYlPAOhOTy573scdM0TS1PNL19LOAWU3zaws471
nchZpwoBOJxRfzWU6Q6+ocpZIdmXPd0n3qTHcoGDLKxUHciLlACzIM6hPYvI
lOO1tzG9WVUJxEV5/ztQ/h21pJT+KoLp3p0K1WUOy4vF1FbI32Q0nGnaDENX
2Tx1vTEl6vDOQWjJ5qIkYs/lyngdmu1iavDILfAN+Qdg1S7RczagNZMwGRQQ
9rTXDTz5gniySi1sZ744uLkGzJuPlBdFS/I10NhUxa3K+Pkw2XyLUK9+AI4e
4vFG9wmX7FVkKIs2IyAHaqBDJarMHxlaJrLmEpnAdhBa8yHZKwWpBsNtkuDl
h7cMTYlIzR2W+dtvYNSuy8PI8x081N10cK+9qsDud54bTPz3eTQvYAEKR/O+
EpDuLyDlokv72xtwYnoNc8cArzX5+4LKQBUw9ySkZJFI18vVoOYROpK5ZXav
sXGo6lRIwGkSrhNibD4cxVVRQziW9WW3ELwHFpbToqb9C0WAbz68xtFK2kWk
SECIE6a9us5qVf3+vPUwbM0y/fuB+byWNbtbI1L68IOrzBaALsRjykK7yyjF
uarv12EATDMFN0hPYlJxFFIQ56RHOkEeIMId2v8W2dKWIrR60lub6HT+mpJl
5UUTHLdn1LY+Beh25Xxd3AzeaUs9eMpHW7v/AJIXjqsePGDYpJo5ldT/QKPE
u5R9nZzINNVI4Wr5HQoZEWc8ApuVu9nKxhO4bKwm5QhenTjcr+yoo9x3g4Bh
nuYED2vkTadIFQ3210PDhi1UDAoFfHjHXxPj3ZbxRtMjUDEvn9vsO9GGxOfR
D+zyOVhrXqduSTse8UtBq43f9Y1rstqL8wGLuUgixZkHfAJ+hBNYg+zs1/zW
KnIaHJ0WvrPldGZvqlzHs4H1nq30zrveeKFcsoCqqEyAOkf2BuHGCVtrzPoO
mn3beDJ6fFLZuSsdcFdzcBYKGeaUlnUsk2vYNLACuQqQjzWrS5ohkkzjvUKg
TSL3fHStDLBIGhOMr8iNXB8wAw34SdJGfLcHNpZ19WuOWp+vV1cuXZLCmyBq
DbIvvCYW7aSMx6mV8pRXEj4bDpnu3xrmbeOhM81Q4ndKZR5aNLMC/CLAVyr5
hkBDSayL3HITzc//Mw1WOGHW1iSkL0xRrKxJPo9baHD9okFdRqwFYUA+zJwW
qeRTdVDnO+UZWd2450HM8WJK7Y0Ac3phNu+PmC7PS1Ib3Ceu87P9uAVneyXb
LNSfpxdC266STTuocgAybEHob4FELttXZGYfP51lVQHItjKBTq3DDhAVGwB1
0IHiz89KTgXEWPcRk8HZqOIco3nRZjI4AVmg+qVq77hCPgL1jx1q1TejDVdR
d6BzxvX2ODf141rAgBIjbzydP6+g0ix8hxjtCysS3O/hZ+JGQVrAHznPeZu7
4vv+hy5zc7M/e3nZ6FMbPQ5LgxUp05xk4wXqX3CwWicyAUSTHnBZcl5KhSYj
oTpKaNQz7MX58LYL+z6hFVTEZ/XKIyXs0djYcL/28U/cnyNAPS6G3grq1Hrw
W9CBMba4OJVQGSfy60RuS0v71dlOghlqc82e9v9elSji4EnPPg5YTqe7o6kW
spQJqYZBXHM1CYkQZtaqruRZ/iFJEXrNGLw5xjnzWE06uP/zyu4qrz3JeJrm
xaXqGmsk9KgdeLtp2mHnXOBHx5ZG5J+AtbmQjvHgx32ZTYTgFId9FVcaQpzy
wHjMo17z5okAgjT7CDjT4g1mTHjC/8rZdNBrG5F9hZ42C3eyGojOKHUSQj68
cSOmppQZkdk/mOW6NqQ8qa+3AyD1XWKgtqG57jx6vKHpHjU+8uZBDVX4zD+h
QK/dX7kNNh7wgG7DfmAE4rSx+Sx82tDNQVaXTzlCrpwO6sd1m4ydwAEFatRZ
19PHwu9Gzg3dufhEor7VyPXya0RDq2cPTcVTn7WBMNzVeVMdAjqhFOWMsaLs
J+/it5l+3X75M5DOXkpVgwm/UVeuWrOXQFZ4AX7mZrkTsbK3LqM8hDJN6Woy
djGwaYNx61II1FA4QqbCxbmfq0XNTmhOS8xNIwsbxAn5xZKmA9niKA63P2k+
NzvGKxIxdMn3Yr1ajHrfZKnUFvYUA4fdyxj94xernqYKhv2kgzB+r7hsI2xr
YYum1FTFKnVse02ePnh9d4DjUM5h4UTNiJIb4+S7p9McEEYQ3HkfrRxE3FLr
I2s/z05eh0+T7ODIWt1zqK1dwSZuznOKLzEVLLJ/VW6/tANLcQLkgdB+TspV
5frFVqQ0WSxp2uWwBf1X6zimzg2vIHFhxOMQs/7vYQZMWOLW6nk4qq7eYA8o
FJEpUlCTiKSz4o3ZE+QEBn45PSaAkknihQEpFXItR73X+N20XHiPTrBHjPVP
cI/Sl8T3jMPkkW108y4WemSpr0NJ2pAgbm5y4ITxKLmUkyrT/gIcXNht5sAr
G+2LJhatiJMLEOkJjupXRBcJa/9pSQs6OGTYCotfJ6Ht6h+saVS0qoVa8moE
KCqwIhjVTFYdRdp+n/9jOFClAQHdqP+RdXl9mGhbIt08cdd2ykO93G/qyPGx
Kb6xvgqAGY40F3HN+kxkU/qxBFCPinxzspIYLRHcA394O8CyARR8YxR4j59A
BysHzrVcM441bGeG8dyyWP7h+5cPS47BdweS2JadfMon4UGeor73VMeoNinS
0IbuL8vyIyvShn4w8C014XqbsP/ptGFokHVk2Oezri3IGe2L7M0nQ5LQgFp6
ugGrjgIuZM8cM6xzly1No2pClDQVRXI9rc5rHV9SS58EeKfqZ83wmiFvUWkv
7LH1eHAi6TcRr/stEpNBxQGzb8cpkxNGEAbVmRO1/n6TevTPhclLjiByVdir
aCLi0a1WC817JjQL3VLMKUrkVjB6C0tl+byoGtzGzs6xsBgm7tjHNcqtjo5/
oFOaoFU/Cv3hXZ97Bo7Ujl6ivzfM/qFep2ajmV4rrhCQdLleiZd/LrOMYKYW
XOT5wWPFT61AvnyBrl6Wixa56YLgKiVIx372RfF/UBGw0i5T6qA5

`pragma protect end_protected
