`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
LCoxgRPcRaNKcAKgfU6TauTzZZ78LmbdBTTHTEFfEPHKFv9CTqllL33O5yAQ88gu
5KRhwK1zKxZzCWW0XvkH233fy9BABkcNjc38gCBzLlJBoX6eaMjk6hjBxBE4hSFj
VNfOgQ7Tuuut66Ck0WN+C8ktPngcSUKTby1L5doqMrs=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 4032), data_block
Qu6n53r7d/x0MlXhbpmbuGen2NRUhzaDJ2974n8vgJXjQXnrnnEevlPhtZEHoIO+
jGsW8zz+c9M9ubd/gmyI3QU/evt9KSbe/y4KSEfZFUFwohLjkhoza2bflveUtJpZ
FUFsbvbuhFz874h6LxKsoNRwDoRgC9q8/2arfuDVuhaVxjB8DktHENOn7i0domUg
xETwAjhktA4Axeivtyf6XMy3zDJoO6r8mRRP3l6Aa4w4ncylcCkhC/dy+eSxfzj8
vqGEz2Hh9TCHFaoY6jsGkeoRYK9k7pflXVQXMfHzthTOdZfp3xq5dO/7vfpbNEyz
iAatPGn49VyCVHrMOfJzrUIrmkiHPQmGRdhTKffbTQBi5U1K0bKKIJBdeto5Jc6c
6tw0MTl3jKmxoe8Fjm7aX7q5kOKFF76UOSxGCHss3/pQc0St6QG5hjlBhZ5rG8j9
oacCTgtH61K/i4pP0Hjmq3Cv0WrjRF68rpUQchO6ZBGTP9NDLtyE5pkQ01XwGPwR
hB6o/k6mfVzdvcKM2SaF2b/j86xbRcH9MjS740VSExUPAqEaHOYyDJQWxVHyV8tS
P9t4E75jD3/m2N+sSu5Ti5bHQF8/F7yQfvFgAFvZA1xXtJOa+WWe8Srb8tndeqCI
tb71iNlKVY+aZALEqREYFVcsqZUW2cg8X7+yPcAoPsTOAo4ictS4sudoCt46HOeK
Bf9x3VaY1VPDOXnoKRv61o9m6085tlVUbetcpBCHvFh/hFtAUJsgrMMg4oFEcN8g
LSiOyFiE2+6PkpXNjzsW3PV25etZSRG2VnkrRdnfIU4/X8ZEGILxfdywyjUsJ77d
NHFlhVTKjRaL7NGPRr8KVoHLY0pHuCPqcON1gSD9R6q0SDARHC9+0cVFbEhFbvWD
7EFq4l+/oyuBz0lofXg5iN2w0AtZUP+/957wKnG5rzDYmNYlrqOTO+u7DDf0Y7pB
8yjkxK1F6jbmiKdCdVkr41i/kcatsL6mXz2hVIkUjd+qb6Tx3cgEm4u1JJ3C6ljB
ANBboORKYb9HiVTl8lDtdP6wnqOm1coxwBSRVuIfO0eIzEUtaWr6vVw9ONT1n85B
U23VNeF/yCF51ERABWmEfCTZxyohhDSRNRNcWMbc9zwJ+rJ8B8B6e69BF6OOpDFj
Ll5GGVzh1IjaiTJneOUO3aKxXH1mVeLyx3kNg3OPM8exCzLIkhOy0V29hxgChM1i
fUX9mSgTZ0SSeUkKJsnxajJbENSTOQPeTgsG1z14eVEWsFLGwqrNMwc9o54u62ph
XUykZo+5Rdrtads0JNY27dBWXpJfnYYl547uqWR0MaoLKg7p/t/26MiVaY3ao1J1
hPDB7fUDKJx2MimQZRE4PEomY2qZvNA10szFub5cjpVqWbxK+j1vPcVENfEuE36x
V3Cs3hedpQ6U1CUertAKXNdZefb+lc7dsnrOfUbfY2/HXEzMzPpXPj6uGyqPfAYL
ewIeGy+7q5SWjTdfPRLH4WZSNpju7V8Ts8iGW6BJobF09KcIbbtD1CJsrHHKXBfv
HLURan7qGMBnBw+LjfVmduDPre1JIDxb4LPGkKjpJ3Z0kvPEGkSraLc2oULR6oiV
f5bTG8nyEnnFq7HSz9khGfkXKisyWpRx8VuXbGjF3NdItBpGGMei+bkW6X2JGwfi
zsxsWzzQosCxe3V4xsRSF03FgVlcGybac9cKJJ6vVQkk+d8QGzzaaLHXkKf7MWKY
3SWztV5Isr1PcYhd2B8xDFARTZyf1XaOl7wcvB/8o4XUrdi+AOi6sEbz1uyOCW4p
CybTCAnioVrIpdqhdkF8gOZ4+M2upycf72OX9u4fWG4t+HiLhb3cmoq/s3g9veAv
gAG8iN5FiYFeRlyLa9yK64bN/ASzhIjAIR/s9pSBb+JUGRqKcNR/Z302eTLe5Pes
orzQgxBHCxpTGnh+eLIcKHrTTWCaYAqZ6f2R9ZuXLpzhqMdxU20Rmp+eFichXlmp
PD7K1ORpw0O+jf5F8dCSU6Dq2icjYrU+nwxyCLh/otRWtzwYEmJsjCQ8F2oFt2m/
65jMM7BDG8Xpz+XhE4qZFs5XqifjrQWhw5Arm0Ii/ZVjJqnDYPxxSTa+atjGAHiW
l7ZT5GLW9ufp9wWWVXyO8IHWUPz2fxSWAPBNQX20IXLhOULsnDWSnjavapNeeGT8
ROyzLqUU/HVX5ZvbCf2Lv/1LQ+wD5sOd1qHYTXx7r04NVF+hflRo81ekG+5l3F9+
7tOCJRVEMMWZdfBo92CrYO1TmEOR6WOZyX/dW7ELX3fxjUU69rdXQVOdvrc2TYy7
PGHLd+C3ARDlxWZYaybML6A4kaDGJ6W1WjvhXvJG83QlGTjRqK7UCVLExKeRf5BS
lm9KUWZMHKUB/e4RIHtSpEKbJyrqsif09/F4zPjY+89XcNGH4toitAQjxbap+WlF
DeSCBTu9XYqvVMKzbJ8ALSOD5n6ePMim2TsfXIQW6sKOSx3EVvgfUWkCSHLXY8E2
dsA6tXrZamdamhTG1gTXxU9Hh9AgJEPhRPd2WLjyQFPLkaRScu0IOmf753klxeO7
3ToMln9ebnV/g0pomi5Mv0BYxdeGGdOKrZR/9w7vPeZktKEkkVV5k1yGcXZ0xvk8
vUrIo8FnB2SWKjLFuYLioi5EsGEnXYcbFeyBoQCYAP5PKJgEte+LUDj9CjXsKnSD
uW2rc9EuNMz+VWl5S9cMkAp85GjQv8Lg2Bc3N9C8UwgYrnid7pccKsYX9KN4yDu9
rvpaW+TAnk+LSHfcpA91NuRJB9I6MESH/LFKqcx922pyXRrC+kC1NT2S0dGBN9Sm
OpdD9RUbnEJmDgfesLw3EHRUCb2NDTeN4S+WD7VeXqD137cqdR+V64pZv5HEOT1F
2Zr1bGlnIsxnbMgUwTtnwTPG3koHtDDopra2a8NaI1ARi7tSxo5VuQqaKI/GWI3i
M6RU+/rpiSby4bKlbopS+r4+eJdXuAfdyZkhIpiJOe+ySpCK53RQnYza44nPfMqq
7eg+FUYtwvIOLngCUJfEgsg3MUC6fD6WlZbPWcXAHZ1+PXX0rOIgcDGuEDGSEv2H
PVD3Qc8CTTvOSkKRU9wlAGo/Qr4jv/di1/hqDJ06VTdd72aptdcAYau8OXly1pyE
qGbo6VSvEwVw2TYaMzBj9KPIATmgicGgnmSMRe4TUjn47STpvnLWy/g5GNNlH1yV
TXjUvBwyteS+/C4Hly/m5BF0CC9pXT21mZbg4Ivhod4dweDlg6BZ2vOwHEcxidk9
Xs38CFXWpVwWGjXQJtuvvNgldyNuVjUvzjmiXYKTuHYajIrf1cqd0Lt1Eh82ea8W
YgnNREDYgQetSUdN2/OK+eyRqtIXv6U4COTjqoQtFTdtpjBLd4uVW6ANPPgDcsiH
129WEUD5CAOZ9xTxV6wIHvhiZdzoZAFBKnfukhFTlHRoI31lIT+QSzs0H/59eMFu
d7vtTdwCPeZxFcY2KksPodQhN9c+RuYUdl1vOYJAzKRbbhZU29SqpuFv5RxjwST8
0Shq6zihlHZ2DmQicBdsBSflbuLXaNxleXxOTtYCLE0nhAt5Wn4cbuxoM1Jv4F63
WnBCTgHvA1vdILbEFzeIB0gnqLE9BqZOq1kk8VGy8dccIH3ef6qYLRqwbuMmZzlb
XeiggR6VhmmnbtPvJNB8U+3/K6m4UPrgT9GX1ft6GXHjj0X5ehUMz7v/JozcucNo
YxqFa5u8DlBgSCKJ5AfNsmIa5ABFLI0XSyMdZRU8E4ncTi2F7JdfMk3I4YlPBlzn
jS+o1mMWf3/P6ydyiYvmfluHFMCK6bY/kOLIAanvwE2OGwpS6sjBefOSn4BCD0xx
mDD/L9/v+6G9Lj1/4AYjs7edL4HAo+5MDb+0c0gK4PD5jAGMcNAqIEyfX1FQQba2
FyXJqE/Jfv5mDnZFwprotVIlb6joQlBQfr0o6DcSSRAAQnknAxs4AtyLYbO91rqR
co+i8Y0qrIouFMey+GJ+82Uq3JJdPTuUtYCNpiIuhGKH548ABpBK2iTx9qeQLWOY
Eamt2nnnEu7UIabqRAWZZ9YXHMOVouo2JxC0XNKCVsSr9318mERblrYRmpM2gSGS
zeRukWVrQuqWuvi0tH/kitCfNNhJ5I1lpBxfT4syCji1CBa+NM9MkOzUUgC6Rn3h
jiL/gsnrAYuIYh81JeerB73O0STbyZ7bFRQCMBxWFiOPofC7WYreCB7/GFXGB6Wr
/hucg/b8kImDISdk2jh/0j2QODWHFbnoMwkSnkof7de9DbsMO3z5OgqGlQhVu/q6
Ai9tf1NBXYMnLAsfjdcOo570K4h6zYMjd7hYKKfIPXC50wHJNTHxfbW358er5mt5
LKwuZh5/Q7EBuXhqVpgm2l7WZBjAMbGuh4GP5YjI+vAIyaQzsuXKGAXQ5ghdGIhE
dvjhs+Ol9tII/MyFqYi9NYKarY0ZLGdi77SggVt+KoavflNb0t7Kz7e3iC0Q2RCQ
hi4MHN9FqkeMo9Ztbk3ecQEbcyTWaqg0IY8AVOzthzS7ASpXcZcapzq/ZybQ2xqU
TBIukuwDt0cygANBcxy2RRu2sGHF20SgyGc1U7jzS9fy92a67DdGGd7wkPa6spgM
zLyN3Ve+4L3PbQR0rMGiUJXcrSjNhz8BRbgK3s/9NH4ZFBad2tfPpx0yNlMhQG4i
dcpmQ4b6Es2yLhlIg9SbqM0WuV3himiefHlFY37aRPkRMNXYcgV53J98yhULahhW
0trLleB2QQQ6nwFFwgAoJ4+2AbVqHFQCf9w94qnR5AJb0IRqUjMA2+jzF84Vv9yu
M+ZI0T5RubDlrbM7Y6ERqfm/na1bQyIj350Z/fbWiiT9Jc4EToT2lS6NqQ9fuICr
e3MacNwGXDuM/vSM4mBYp7oVGOSSjiVo9YfNvmFdOxK5A+UWyZTpmQftjnuRI9rQ
CKGefXBau65BcmohjB6J2Br8+wQqg2Ubw0o//vEblFepkTHBY+755n69vNIeLNG3
f2Tx25uPekxKyANdatI83k5ljvSo3EQB0bQpOnhhB1pODK3Df27r0GQt7FvmPmIy
Q60E292nL6dINFpAhgtn8Sm0raWT+H0I9+KFOmYhu18dD7PH2mc1p0kDtmd/kmh9
V3MQFCAvPMWbTAcOZWQCPTxgAqrHgQEJLJ8Ym3384kD3+wBlxoeAERRrIndh80nf
ULBsN6OWriNrgdB5cYLWnZGK5Z2Z3O1vo5gpzu7FBY2+2unlHhLqqHl/MhQrAPgg
HUrFkAM3maa0dhq1Oe19mSN/dDvueq3kMZ9MzEeTzS7+rfcpzJ6KWvZDW2xIIk40
AcG5EbFSp5KyfU9bz0EdvMZGH4XU+lTa5pbnPitPVHZFGohjDxKtfpbXU+b2j9TW
`pragma protect end_protected
