// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
fLnKltq2XRQoK+TrdWJ/ze9fbG59mEIOtN94vqzRzpz+VZ4nVO6CoA3JqqSVnaZgcd1ShylY51lL
iRz1qJfNrW9TAgY/++vll6fnlt0up+Ce0j8QisB3ArjLokmh9kYTSi5rK2ws4litkp6voZ8V//nS
QyLwDhHhQlyKNoxOWJ7ywS5odqp2VoCAUAH6jENQIEI7ZL1qfDQNFL/O7s37VgN9uhrlTleUV+1T
Csp66lpjRZjQa3qEBIgIJcsmAOB6mOg8QQyi8L2WwMgasrpt1grwvyAIZ5OYWcxx7ny8gp0jbkZE
dNmgKGgpxiRHHIi+k2lOlVLfOddAs7lQTtJmFA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 22160)
XTZ+TipQPVFrKJrW0cYl/3vXh8MO9nvECXQwRGIwrPJgs4CXvjqROnjSudag6nt/MT2lktqndURA
rt2IefAyEJqj66ELsvg+SZw4hFwi0eEPYoSvJ03cgYh2z8S5Y9Wt8dUUGspn3GuEi3Cz7xWV+w7J
rHxJ6XZeulX37AO0xpv7WTiv80kz7mQKHtnMtuUf76w+xftOUR89mNo+EI2MRGjDwzym92XhxyAu
vAyrfMBfshScgBqADnwtKVjk0dMLig7TKFlW+AdMdkukFJ3ZlLz7WoX2YIZJmJ3fjPI/hG9ow7oP
8OSr4FmGjp8vQZZ3mLRVzhNgKhCSmcuN1wOit7C+aMa1u5GJhvJIkWBsCgKkBfZt6LPYAPo/8SFa
Z1IWiLxAvXP89HX6pQ7NHjftTt7MmOcoPP8Xjt7kUhcC3PpwXjgphGjLYq5hFvC5hSL6sXJ9gGvQ
/6bWhYlMjB9eo5YTx+8HDAo/7TTRA4D1rKSSnjobZ5GZlJS1mnQ4ymzM2SmB1nJJ9QPAPuNx3efe
21lEgQZuZWKhj7sKDNzmT6lKfFaFIHJION6wdRTzWi0zFyPdVrr0EbcAO7H3BIaq2ndaz8Mq3k+C
zkYM29Tt/6zZdj6zyn6BYcjf283XLs0EioXjDFtGluh6iCu46LAJvGCZxABSDSk6hhiLkVhtV7CA
ndhGcyvHInRL7UrDqQC3aJqq0yOw2hoNZ0SjykT9KW3O3k4uIDmGpuupaJnTHVWM+vICSsWuyfta
dBrCd0UMOejxtNH7aR3A5ydL/6ee1KN85MExTpUez+XuyM9RHgMawTe1cxgHTawOXxkVUzWbu72h
wmiPCmtP88i/VLLj1ggKvOXhxt5tuh8ykM1ABFIRPhp2ZPIz1iOmaYtbCUXu5JdROAeYP480zsPL
a7C29LrFujQOQFBVF4i454UzvtXcnXCiX+z01gRVfsAawRKXBGAtG+GpKP03XavltKvHDDNPQIx2
jEkQTHbeWh3VPfRDez8iXpQHKsm9HBsfFqSXpCmsPHraGP5IQed2pz4dSv++jSmSYaLlHLaw/+wa
bmECVp/goQxWeATcbRlnTfaUgFBREMr6dau9UAXB0BzG5y85ykHEX3HhSu8+wbK+c45IanI3CP+3
3/zdpqTdzXrWRir2iHYlvgcE+260YX+PM2hJOiurTuKV/2HfHOCwk4ouDLkJljfMyt9W2vSQWuO/
ARUKjrPbuIUSNAYPd8IeZDaTprlsmXC7lTNLDSKm/Dkouf3CxzyQWrLdtGglwOJP48/7wJUdHeYY
creRSqfB3Wk55jQlEeBqOj2+9wQHr/T3iF2/9kqqxunwiT2njQR7B598Q8O580C5bJd6VY6C1Bb2
myTo34kPqw4T6ji3xScj7b1WOei32LBiKIKv5ZJBreSUCyy4gjl4n6/JhN8t2YF3kM0b4ojaaDCq
Kexqx6O/AHp4t9DuMO54tqQpdLKVu+oP2PfNaDyqQ9fUuG88UmspcrOMdv1Pe8DEQplRfyNWsf6j
o3tDmpaJcFzEactem/EfpwqE9ND4xne2eDRbGUgiwt82+A3yvq3EPI6togt6lXPlxsavqrmgKWIv
epY8fhSw3EnAxfmFH5eaweKAJgKrHH6Ega2EkmUa4o56IWfoxBbg4t8cYppzi7yvhYs5xJERoQLx
nlj/ki93DHcHhQsarF530oC7wk++4gdD5cLN3M8my5mZEflhGcMzE4j0f68XqvtOdIbFQb9XbYdF
AgrXUI17I/tcv+npjP2z1c+RxGRUWTHInsWHyy6DhNKqFfn57GXxd2nqvldu2FZMAOS7CecT69i2
xz7ECzP8P/6Lo5SPy9U9XnxeoiCRsX7VRY9UPqHEsgTiNC5TMpFZtmOzetZSJERxDhWpfGaa4NIu
W8rAX/Ibu4Rt6exa8Ccd1OgNMDdt+0KWFpThFZTW2j2TyQforyAmEr6ShmhVqbrxT92e9T3JHs/L
+wywyILMEm88eSAEQ7MmecZV82MXdsAlSpvrUd7dzN3M9L15KmcmToIaP+zfFirtkY4HIiLSVftl
aTTg/Ob/jZ6A59DeP1OZEXUwgsSeysO3DiRpSwm1laqXnhOzc1bh2CFNQf/SeYhWoKOoM3zCSApB
BwE4GPAs2FKxTUcu/37RHKX3Lbj6i76ICp/obUhR7DkQzIKj3BUSasWwtGW5D2w1o2l1aYPHKUbk
n6L/WNBxuLlEDVJKbi7WcqsicMUhi4VWPQSjcGJvtQpuJcIVw6/4FB8uZiyte2pGe3+44IeFQRu0
wxH0CDWTkga7cHsvmG7hU7IkBdqrnOOM3toQVCtl4ZYaf8BVICgDxLGqigkM2TJf+F8l8OhpZHuX
sKo9WwXxkH/huQU+f2DZ131M8b/8QDxNkQtYicDPSt9D8+04AC8onHJ4qdVtP/7pTtVBGkDSmpwQ
0aJ7HGhV0sckAs6800iIWwBrNYKs4PRFReVxl+aJSTJVNAisaSjPrS607qfCaGQfx63HMgHUeCiL
lb9PfbkJOfqMs8Yhhp3R/JYiLz9Mg5IfOONF1IFBZMTgH62i4D0LqtcZyAcauWmZqxLft+sbM2A9
KUKpLBTO6q8ALJ56bA/TrGeVsVK/hIvuw4l9LHcM0oB7g5mNZ9aOKNFEf4R6s6PhVKiqjlzdAKz7
6t69aGi/ATv0DokoJbu4iOc6mOGfgm09dj9OXD/RMxCJCy+MXouMg3sHkmmzYFTqt1eHHUH6bJRL
Qj70bwB3qRrW1EXP462MrNxtL+x90tIchtol93pAlxBrPk4umvkVXBGJYgvcondpITmjvysW9g7+
RLW2A2EfKzOu5n4OajOM2Q7W1WLcQC1vVggIOM25MrU6872vAoqJ1mMyn4m5qYxK/wCk38cFlb9/
/WQ2s/EmTtnJ1mLNPx4qY4SosrkBJjWCueprqXUORetEZG5clPwIO/10B+xWbMEHgoSkt2j/Aee4
doeFKsqLeWoKYe5uk2D3hcXBNXm0fR4LwY5jJEIK37GFUcZ7i5cd4Hytru1ZGuovArXIYjnT/phb
Wg54uJh5wvOMuYcZ0phf+f/sPy9XrsMFLjeGLa2B8Xd0W3M2YMgVnN07gj//xZ2t6tlIQzwF4STU
3vItEdCTcD9jjfKpTwbYFIYukh2IdofA+xjuWnzQnUQ0kuF+A6mXyYAR71z6h27wmmFsiqNO0cXo
R8dhwX7Q8O8lsfCd1RjuAMVlDLbMGiXGpntcqd47GDMmOJndMosBQmwN//dNlK0zbNjWD37koRCY
AlbK2OYafiDcgzHpV4I3tqRqO6uPlrv0snDp7KjGMxspxcfDOk15HJ4SE31DTR+ATJQLaQYA8HAd
WJ+c/xx0DhhTLc7RV+wCJDGFPOhi2C9f8l5erRyXAowQjWGzrKv1EYYwQjEHT0FpsPqB0FcslO2d
qzBQ3DZvpnLUEeIVLGdBbZPYb15/ofAz3mHHNeyfaNrb3UmbCaOSZLqjF59xHVw0M7XtyLnQ+58t
H2kzf1moyEjeJvY/5XJIeUI137HVgMSYNj+BNj2tZMx6Ga93UI1asG1xvhOppNzATCgZeEwSVWAy
RmhpzAGRF6lLcOLhNP30VNWWu3koo2mzQagm0ux0O9x3ohbHVw71n41yHbr9fkqO3eGg4YkJLbJf
IZMP2SLDtxUCUqPJmhimM1MEL+fusVPVvOL4uda4eihFd6zxof2D3DuKiQeO1akxmuAyDuJViiEY
QqDJ0MKiFYdYyHstMpHDueP3WkAa0is2vH5r2T6l5xsfPE+p7aZQ1A+fi1EomKCio4SNGbnSRSL4
Z5LQYpJBuTMYqtJbMI4bZ9VKnvPYffNcZcnYVGtJxz/L0xJg3l3O7ZOhbVvp9xhOHnwblNdlIxDq
o9T+dM2peNHisOX2Mj3lf+FjlU2B4eEie9/ye2+GdqxrezfuwbwgDT0CZAWWjCnLY6nlByF0P55C
uVyofBodYNHRVzqwAf1lxsXcQwbjG+hYLgdO7C1of98knAf939OJkLWe6J0lCUwFZ8bjNk4DLOyt
Dyoa6G2gizMqznfdFaoalmeUhwGxbdd31KiY4oJso51TNRb2QDa7BYenOBr4oKn6rAnAbiRbbeu6
PVVsIPk6guI+0O2LuyCY6IgmGjAkJqUSKj6JVQMVSep6/OsIMdnpLNpHjVRa0yKfVpURgBdelLd3
ixLwhUOq7XnQa2klnJa9Bw5HcMYx+Z0PWCnuDlCKbhvp6d0mV1JIm4dluE+KWCOXta6yhfb6VkdW
VYHL+2kPm++fZFqwXcaNzGt+fGpi0kh5pd0mgFRYnaMKDSrA3YWfY8irIGUHrqlWAc37RaU/RgML
+SN/DoyJzECtuB3zC+cn0t6PBZSruefFVn3OiHq6wZo5A23rYv8DN2QBqJGdjYDnXi/YWmdKLY7N
bM8mgl3vyymVHjGDdp+LcOi1WEYaFHnSbAyTD0rHvi8DWke4SBZle4r3u8yM9PkkvHYt/HWUTfF6
dBYJ9jZ4cje4VCwMa/6bYtniHjxL7EZwFQVZsjTW1MqobpxdeLWr93WvkbrKcqVRcfWjFzNc1mxJ
MCB3ty98vhdbHJHsZ72/2I7Yf2UUTBMrr9ui+ezTUpzKbDvExCRvtDB+9XkU7LcunbGWqMdBD75I
zJ8/s+I2ajIMOkzWT8goARdS5r2rMcVOnHx7tNVxqB4SdRzDbdJkyHnm5T42+yfNiY92hk7zHks2
1auxWAjBELlrWwUdRBorslCk9rJ5BB9StfKL5a92h/1DP/hWeFc2mupHV7R9gsvOPmGwjwA8fffq
djAceXjdAxFnwY8v4/7lR76uFhSXUcOKRgzL/cA36xgoAG/tvw+Bi2eg/ePoe6BCUgL1zH4cBjHL
fraX77mklBJb3910dhCOS9V4yxNQHEih2MEsAdyH8NSLl+cxm5qK+nKc2qSgBj0AcNWB7t9EYiDb
LMLIPy9YOUAauDMgMjNAdS0cm5UvT1PPvlvK4Qiz0PQ8YOpsIv1oluki1Y3rB1FlTZO7BX4ujHMO
c+0k/5G/8Dc4OVEmN2vXk2MPQRJs4dFlYWR2DwpOGb6rQmjiV8taFKLfj3Fkg8/ubffiP13dA+6f
waAwbvU7qOA14mc3LnIQi5o6pnawZIzMRGxjPMPRrchJsi/WcjSlak/fSEbHMqGycszRt0ldJsiP
klPGea8ls4PBu3ZmdnFB7ACffyVbr++Zk/Z7FGHvzS7T1mm7HT9TEM1sXPNjgdq5RqrTmt3NfcHV
O/VSicsS9SIqXLHHX3fzYzkjQuBfkLLkUBDVMw/pVHMji6QEBhtCZpXIKehKbzjKx7atbwxFLKfv
7ratZWzNEN4wSJ2/Hnri0Ne9f2n8pQQKHuBBRchaPC4OdCTUbckn0l4P7Ld8d/SOpt7m+JS260jy
tS6HteluSFc4klcKJo6PtGeLWN1qqMUN1rf1SdJUg1mW//otgvpIKj1KnsmldM9nBkPQLk1gHM2I
TurmfzWSuuPW0Xz2xlC3k9RnFiCp3Wt15YVsHc5Zxqk04u1f0/Od0y71lXsClwurxF70kYHP3Csi
TbL7pItDY2ACNP4xD7G2s4+OzJUxThG6Y7hA+ZVYLTZypfHFQXjUjqSTKHIs0Gjqv3Ga2vFu+1H/
uT3+BEOQHLrsRm9oQ/m5FnAcngTWG8hUvlUaVOqi5SyZ/J7i1CB5vODYlZMtfd1/1glmWe4iMFe8
MSxgimd1L0Ri4zjNYsENShRnMK/Zd2VlbN/neQ2kg1bloZMqE6AmgJn1owVwdNrg1n8LC67EriVC
+9bnyCTfkaNB/dp7vOwH6gJvf+KGSLKRVU4SjI6VDSZXIw/r/bv/dRVJ3LUG7vj3KzIFLjNzHgi4
iW/ueSg1rM7M/zNiE4RvWvKLhk5SnBdLF1wRE8TLcD8lNMQwLLQM2rsfHp1ZgKW96SYjSnsnkfgu
DsDFy0//JYe5a2h+KGXYWaP6Sz0uFVc26IKti/Aob2YfVxYINtYY8MP9zwQoQlaN7ppr6FpU9j/f
T6F132inUi49vtLuiiGFihOH/AEiT2CBsrgNREOsPIYq5mc2p/SyC2aCIsLp8t95RasjO1tr39iU
BZzOvU0y/qkCiEbcMD+bGmRvyCYMF7biConewPvqXhVKP9spEfuiU6dS4h7+0u0Vh49D5yqlaBul
UHsX+616imW1x8XSe005KGxa5Qq6anUuNiLHD7/r1L4xsUqzWrgbU6H7mt1GjOMw1rwP/enRIHUJ
MZUBuk86OQ3TXBVPb5KkVc0hiDvoSTlArAjd7Cis9UOupELwuYD5lBd8hllPYKtQyeMU3M1CowzK
iFreaAL8Catbu8I4P65664SJY8tKvif7OtnY9LNvd6durimJ3wySsjNh4DB8IdoXYEZjNfXDxqHJ
hwsONZxLVTb4gqMJpw0gf5tVyQZIFIo76Q3k+qIhjpFeS49elQA+Dq8B/woUlY97oWYybgsz57Ue
VQONP5lF+jo87cdRUty+poxSl06C+w6ANxKUZ764JBomLnOhESuFSg2n96AzUuHvbYHgcL0+vxPj
EjerKq/j1GBOECdH6qTV8MJXpNpqTyFBSVGMjdNeAXddByQLIudCzOuy0ntHenGpRLwLmTGWwGDE
2cDj/lKPJSfWTUd/OdTo8TpA+KhNolZk8fs0F8zXeIKF3xgro1Wn6sIz4h2TBcDjrYCrIUvHKy/6
Af29s6MyFvVQo/krA/JeZN6Eu41BzEPR5z9zeoqeJkt48imMg0nxtZcfkJs4QQq8wwb63kQnpLJh
3EvGdiAOU8YuUF5C2tbN7OKCPdBrvSZez5/K4uJ9/OA6tAwDOmqsgfWF12QXkw8feWIIJNjCKOpM
sDAJN+q3pkCJ/Klfn8g3wVSsCr/hn2J1aKgZyig7fdU7+frCL7z4yBChRuOzeUn9Q2IpEn9I/wmP
gECJ8xHTCSEjM4gJMKMakw3LPKTtrAO/R3WZHYPQlrflcOmr0Lqv5sEn9X6gW8W3tBU3mihsgyaZ
VjnapmPXRpvNnbp9g3FeQXgwvVID616SBt4UBv9IqBPMTF8EraM/NiCtoma7smI2jXoK/teoWGeq
ZtcgE4tPDzVIHDYGGzV5g9xezsrmJWhkz9P3OP+bTxg2jtsKQg+lnNzGiF7q232q5FlAWAsLmqkS
eNnfZdchHQ+Ms5wCAhrO3RYcx+sioGB6pF2WAeSk1HwKYBVxrasy3zpJ/jDa4FiRP+woFOlY4mWK
7O81cmGPwYZAv7v8tvvlE7mHk9ZLn0C9bhJs66UTnOwCUYslsFl9uCahZpmHoogfPr5c8z4CH7Jw
RKG8CEp0AUaToc1tvK4NeH672Exm1hRa0MKPAKAQl9nM7ZtaR1pwS2/lTRS5VZgmN/s40PK3uCt6
TW5I/HeY6flqgMSKa5jJMcJBEv5G8L9KqTLUxL/SDPYAU1jlhzWtMZ8BjRgNvEu+Yl9lDGGrPJrX
nZ3yNkFzvZJwYjwu6TvAZAT8JvbHtAB1ERc24cL+/4cg3fq/qd8hQHaSA2JCsA9ua2b1jTCoXabz
B0yFQ5yyB1sS38IGd2j4ZGIto+GxmAfYkQQxJtbVrwjGGU3mlsJzhGBfnWb0LuSv0TbLQC+NUJvT
SYC11M+8tgw8i8IL9cX1lBjRPxqOviaB1kxtrbzlLF5C/PcSM1D/N6XdH6idRwpqhaBfu9Fn7L9n
um3QuyIprInjAnMmZBb75Lcg+wS0RmTZHkjc1MoSA62XZq4EkJyy19b+wVkNYaLllfJJXIA9c3pc
IYfxkPUaMXXEsrFcr1mgaFNOvlSTjnWWlFlSucKYbsD1ui5+HnTQmfbzDqlj8Ae1ZoQoAvgVjLpO
vCRmxZoKrTYtauGEtS1GMDj8Wg8IKLgh7YTA3m6Ggts9n5Gh2gVszBBROEPaajB6BDdiS0ZYPWNx
XpDkrWX3YTCzIUbtWi24RSRu8SWa7BgUVWt90mB4V9ag7QmjD2cy7cMUiuXCyHEsd1cNiH6COM1T
v+3iu4miXMlBgMjfocAxjMtEShsmFs9fEPF9qXTrrgQUv0RAxGMm6PuuTIB6k6Trnimq3RckegBa
vOi5Zv6jC6kJtp4+41ryvXTWA9cNR2u8nv8nutrhQ+vN7hz5lLiAzUBKmWnBLrsoP4xqRTE7eH60
cF76VrnVf/Pnpr3Iy6GIzs4grpFV06gk5sA+PV71O62RybXxABJUzxUsL6zVNz49jdjKvf4DmXIT
lxFNrFpFvhWgxhAaWZKUVfLY7Q458dBhaRsEl0vcxxkEFUSjy5k5fDfBS6jGHd8TKY1Xo9sdb0o9
iw6/a4W1d9ETsrVbeYtBPgYSjqRtnuE+6yIK6BVGbp2vAmQMV2haV9WbShF+j5utsfKLsp6++47G
PmDPEzH8/nElJ9MJ1rRH+47vFa6ii8EXRRinsDmlIbydYhhonp9BWNSUUCmV9D+bDiwdIBD7SJ7U
RpTmrVqtDLt2u6tILP+92DBdiqOwTxK3RDEIuz0CZ1Y2Xsc9ogWKO0Lg0M6PrbtrHAJ5xhpck/pL
LrYZtbFaJQA/P5HOsdGBZv/EroZKkTvkPkTBp6jAK70Rsy58CrVWDtroHbEijp6oXCqic7/szljx
hruRUoPdJF0OVWXA2W5qo/i/i7QeOmiB1jEAXSMRw4K/oUtSl4MvqPv+YCBx6c478ymVaCjO2cm6
Xsxzn4pJ8HAkDB6yu3iUFAf91HsmzqJZNP6jUl9KU7bi6v+sML1NEutMMkZwJj68NrEPEtLhAJUe
Pg3Oj/UHunJCu0d7AcCXunhO/MmNQ7XFbJyUBSjhQqa1CHvVvkCEX4Rr3l6YhW6G8RuG+4Gz8Emz
drrInjp8d2u6QWhaCbT+Dta/PGxkjfpsddpXZs+9PzitYOjYHh2BP/0sCZbWGFOyDWUxFLMvU1II
9JQJxYkG3JNvHikCY2903HdEXfTRufGEzXuqvLKeAp8sLwu5HqAaaxaBvOZPGKFGLPVuo0dTQwMg
W4JbaMdbvpfrv1/tLdIGIupEWituekyW7QpVv2bliKrtfr/T9UYGRHB/ZLNtjv3xims/KRhOlFJl
ne9ToLjnSN2SoCQbHiPNhAq4vcj13zt7rwA49f4bVvshzt2Ogre0hkp89ivpIdbeixDl+NmkfAb8
dKuHfi5ZmWOesPqHMnIR1kHQ32Kk9UbkwqD0xjxMx53Xr88zfKgG66+jHIHJoUh139ZM9XwAp7Ir
ucG3tjimrL6UlmXaobLORay0bVukAJWbVnJst62zE1jVENPK50nGUlsg00+8SpYDNQj36Cai/QZG
hwlIZBzTgqQ7XEX8GgqV5dqB5B0YqQ5jb32cVVPEAqjvwovW9EPSS76bsm2bQLtnQgCrgU5SGeZS
QYhb5fL5/T54wMPJUuVnuAvzzUBYUXChbW9gceMeGaB0pV6Rr8wXArMMdLlJT4UQZNSsogRCrWW3
BWiHhx6wRiaCCJIStIUGTZq8Qqkiu59m8xiRPMcXEDMpWwa3cgHfJmYjKNewS9CWk0vXUTB32btp
jtABpUvZ+qbXirQzI9/VqzXDEriTk3/tTpJokaK88iPfhIEzW/INx4fwsAcPYCH/rb+DksWPo4gC
OC73Q6s4bpnvjEzqgsko2m7G3MD6lDJhi+Qr4C5UMXYTOBFr+gLSXB+LqBrFnlxI4vSwBPWX/7iy
6eddKOgeRkLW9pULiFptzLQEz3Jqr2NaHj/k7wRrKIO6x8alePXZBIF3JmnDpOUYUBu9lQDhQ5Jn
HzZivB18NujHddXum1+2WkOp1VgUc49LEJpt1a/Aea6U9jasKD0iijuMsLTAUwZKslNIQGLUK5mg
qzMPDqfcsNu8VQ7BqHUQ/8IqqPO494DNRfYTbxpIdLLv+K1CfG03cdrgrhiaZkOvLAQXS1qGIZTt
iemA9weUbN2TN9iJJxpCuCoqChcbROfiw+38o9FsjBlpgKeLp4WMWORmrfOapAin7D13zS5Idnm6
KF+tFhfzAE5CAgD8n9hUa/7MbbFlJHY6niLKYoy7z2lHr/cWeoZc97OVKAG9Wg2667kMZf/x4Z6S
7EyXC+TxKeVJP4ZSASUcTEHYZPcqqtd1Ekhp1x0grcfXEHNvgZmyx4IjFafYR7ReaM+YQLv2WVOp
ImASgj6LTXN5U0Mvf63SlbyhK4J6P0lC2c+i4N8o1xOk1sXa8Fp92G8UEFbLulgihIKacU1GIvTJ
Nz9vustZ9HGODRYR7cbcBWYibj0MpGtLls2ufJnaPP26F46dTIKGRJkEJED8NU3a0r00BVImtSnG
G5uFm3IVv7iN3VPJULlMjnOPJ/v1/lVJT6ITVjyqm6s30G5kGwBaiaKQKEMlaJ1MLkRLK8j5B1fg
Gr6KISDXDJLALetu97fW0xKal0hUGM4OyxAxBnOWsMpn+Q8M0R0VdOQVjoMFZFXvofDn4VLZMOnD
zxF3h932GtTr9m97DUwKfeEqsTcIPEaxJJdCXPeF5HkJV11gZkteVYaDUQQqdixA21086WAhaPj4
pzfnW0pKtrMnuxqF2s/NqcY5GuzRxIRonnSgGdSFIZ904SgSjrH3tGK8+5SR9zRd9Qgr7UlmJBHk
J+StQmLrGSEVMxHb1RCWpAflzuZZGDn5JSdcyfORyl0IaavgfTJGYedMWnq88bjq2HfFcB3xWwAb
TJqwhFtR/Oes/t9e0LlgcCHKFgJPZZBWn12xZjzVu6z1Y34XCLUBKW5GL+mDTwsqV/c7W5lpCaCJ
149aP2a2cx2w5cVD4AsGXfggdCGsU3uPOROUCGSKRv8b1h6m3/8NXq0dsp0k1cLYISgUsyHQuMl4
eQHIVytSD9gQIQjAhJQwX14f28EMwfZCx7zgwqZiGAPMP7IPbGPiQYDIju/EIPPkGFHgAgX+wyxh
ilaRhNIA2at8xhodt8bVzMbxqFPOAtR76tZGq1eUwbJEmkcnGvqenKZdP5cDmqfwthBbNFn4v/CS
UsbZKGJeG7w45QuX0tSWvjD6AYkuUY8QoZqgtMJ7c4W2WAL1aJguB1WDuDzCvP4q7zCtlN8kzV4/
yMr/ri69TIw7MN22lMZCKlg8nTZCOE/76o4S263va4rU1/rJHLm4QKWNbkA5qFi0pgCfr39ybwHT
eNynTY72BM99G+ZwpAvuF8HLbIavoaBUvIw423t3cI6CCo4Utcv2G+wY1t5rdapfxrsZxyPC+/7m
OrP78xv68hxzSzpa9PznwcZI0rd6POv1kuH+Eh7kmXQB+zw+oHiV4arfxMU7gaUvhxJiBoFB7RF5
/aikxdQ1SH1zFEn18VnMxNZWncPp7H7QrAIGNg2gtaNUW2oHRV53kW4G4pge5/f0HeNBByAd9qQe
EEZ4YAOMN0kAkEo39fatqIdPQowzecb13Op+9CMQyMBFIeMUJLF7oLoxjhQkQ4R3RJ4hUhKTMUDT
xE2+xfsexsOjcw/SmjfTMT81mPoZstKqU7VFUGioEFODo4WqAKEbUwuF47wbQAGewYHtORTlo15d
s9EadthHQAwz9uW4K422Ws5XRzwqI8+Vx5YFswTrhATKF2XKboBZFHG/t7CBwpKHan0y3xM6Clpk
IiW1JgAEL4Y3veGDK+KhEaAtdwiuZVWiGxdZ10+nCFGHfkyMmWbCIW3Dn7Q7waGf1Ft5cT1Z6vs6
odE4dsPcHdOlQC6nErSrZAUfH3TXEmLBkgpMNW2+t2kesEpKA/oFvh8mdryJ6HqV0SmSuW6RAaOe
S1frbnmkdrPGn0zAiyZyOSrsL/BD3VMp/5CEnOpkG6gkgIjeDyauZYnUYOjsT+ekJssZFo96b3gM
n61tCu7+mP8EF5N70VqvQ2sKfbL9epwXWBgXcQ4FVeAQQoF0ItX0J4SVHEUy7cVBGaH3BG0Evo1F
kimDlPvFZdZj83nzXUmQDU/2Pw/iEjrhmMwuVqvW1vMsWDvArYObC9KZVGgrlZR8BlEiddhYCfFC
mxx28RVBW6zySRqHb4tofV23Y0o+n8cHY+419E31kfzrQvawmIONT1KRumePeXo/F3xn2/ALup2B
kNjfahG9bTzvxKstaUowsVvJfKFMG5avNFU7ZHTESli6u3YoOARugksbJb8OdhQLxqKyt3mv/dRe
UXMQQ9BwO41824ulNF6UEAFh+/UAYQocLGUIzBBwn9HvYrTo76tXHbcXl7jPKJfin+BDxvWy4KT/
fNHDwpuWFB5zUlLfG14V+YOVPLBMTSl807ePoB95LJiU2S0umRI6WfPpCYhJEZtEbmOd4F9pM+6i
SkFeD7eRLRZe5DLQKtl2kqC8+btv18cn1KVaJOc4FmtcTW/6jpI9Z+Bytq4S+inqkmHhhMY+Xb1g
VaxiqGiAjQ1rYvDFkJHiMixXxE/qr/KwTga0f8xfyp3LSSYKoH3TktPKreOl1mpF9zHlulCDqQJT
6AOu0l6xisjAJE9gMeZk3PTcjIWJNzS3SJO599m5sunJ12NEmV0VTRY1gtW/yWFr/cOE/VwOicM2
xnBjJwPa6BbW/2zeUVNYXHrDlV/wNLoysoedZ2J+M6BMN8cSPsNA86jfpfc55iEh1Kmytb/guz+5
rvozloCv1DgqBfzHP/u9MO71WW8YmCpPz16ZnleO5+7lhgzpssSxh8W1sk/EbJqYoFg/ahVofdNc
lh7A6PydYm7rowqCD1bGAuZSVJLhJbPwpDPSUG6zi7wH6VUzDRq7gAiXa3iWBJ6MANRefCdzPdL0
FcqPwqrzeAyh3XbnQNzkczDfXHxEZji49Dw4VRmwAJN0elwU1VnZ+gCg5obSklwmqvd56eaDVkKb
oJmhxgltZ6rZFaHdTHWMFkV7PANVTZCQtv+rAbVYA9ilQNZwBzs6ZCn84k/YtiWGk/ImqAQC2Lpv
6ASWnpUnsKK0HeqNRnN8TASJb51LwqNSlHYJw40m9Yn8SrpXVeQwdgDgkw1+sRQ1Zn17Tls+67Qw
bHySfHC5P/1bw+P8cJDH/AtcdFdMFXHhDJ6ikNFuHUTJqMFRR8gojHYayjHVI7FZJRQVWq7bfNok
gfZ8Lyk0HRPwr5RoFmAoxi0RYIPgUbXy3YeJ6pbje9f5hrEw/kXCl+M7rjx2cXYFu+fr+uomRzfv
BKOjKlWt1tVPXKWeeWhva+Xre/dBQupOHkBL0vufEDtGdFztSqQTwY6EP41z0DfiFdMWeEQ9HheL
eXou3FcFeXVC+keh4Miz8ztJFCUxiSrGe3JD3D+P3GZVzHczYnAY6+U7CZu3UIgmU1OgeSnib590
BuioyT+dnH47MKrNvnwRePaTma9YgAkIxQ+GsyNQRk2oKVFwRVdfZFBTTV7IHD8d9QVVLX59Y4JD
XY+zX/aJfYH52iRr7KRKHuRWA+TWgAioQR7VzaErbvFEkVta6hzg3YF2yIjnQRc0LQ8TDLxNE/qB
waF2g6KD/+7HAkLooZdUymnGGd2NQG7MtifqgEE5ZJv4/R3d8zePd/AnUqosY8j3U9D7OXkGaCMm
2KLa0S8EJbZJVvbbDSNuJWUmKrpoX8iGFn2DUUnoIlZLxgJEoqIoJwnrKOEe7cXzPT7HKD3Miw2b
Sde8FmlASejdbhBfP5sBhbBAYoKhb5yK3lHsll39h5hsp/nJZ6ObrUXz//TaM/KPOBx2yrPNQ7JV
DIkQMYvEra63/OyeNdDYSgflV7/51Cy82O2/yXgZBXX2Q23yE5uETFpv29tO1KkpNZ16VHdz+xVh
KaJJokFh7lWUoZgZUe+zBwQy/TVkh+9EnkAJLfeUrHkrmCUWiCzlVgR7jIuhX4C68FPU4901Re+B
r4GCg4zsadIHDOrmqoeil6SaBpdlrKJgcKnxzmwF9A58KQKrDvyVql5PRl+FENQZXt0sAhSMduvO
vhXe23RVQxS3ltc3kVBjb8Piz2ctABpHFPzb+mLY/y6P/otSd5KUoarGHBQc7WXV0WMrkyzlvkCN
2mGry0sfwWqUqJe+i4oeBWQyAyY9n1o9+vFVz7ctE4G22ve7DsAb/rv+5BeDrsHBXgcDKH57rMUI
G8nbyoRMZhn5rw3geqOU652hRz+EaD2jpFnV2RL3gh7T2vfkNZAoHHwaYU+DcYEAwfVEgtZoj0vO
xZweun+tkhe/qmNYF36wm8/VDDLHrm0GbXnZRPZSgMlfPHpPsyvRL+PJoypiqBYz9DunWWH/19kj
doRm8+/64jAGWYf1cp+FvIXTjZAzlEEMS7HTFOV/ZSHawZk+kVJTUdD16JCwQ9MQK1AW6qsxsVVp
CggaxaEPt4D9Ho2oiCa9bHQhXZHjWOySrjJHm7VOnD3IBg44hLRQGksiMFqFxRI3IVVRBB9sV1wk
/SrFQQ4SO/VN1JEA6NtSO3y7O/UdwQhbwWshlYZUFz+Ql1ViOFJmObvSvcxV2/IX/P1HnYKUHAAM
MWtW5BRs6qvYDnwHCX4kaH/XsJLd1gOKzJzn25BOLq60g2y/WlBGyQcGhgME86+S/RlYpwA7zxR3
7Gq6PBTIS5HtMcZA7q5v46awu1A1++HW/sjgh0hdiuLRuEXeBGWILD8jC9KOzabSCuzOW71QXRrU
ylcvcqbJ6mrVbAX8bD++BadwSksZjLLgzqVjeL2FG2SOlB+X+tyLOi7LfGZsaDwnoRSGw1PaucNl
7q16lRKh5xIdd6i5Bb3odtqny88CRPzYAeI/MljcC8mAhP37LkHVwmfsalO3GrPmiR1xiqxIroUM
2YFCahOWryPBpnTqkE8CN0a9RymMtg0JMu5Q2hqjVa5tPYTE7swS1mbZPkTKu//oNg628ULEQlU3
dcaS/btKtXHXDqnw/0Z4oaBARLsVAMvsQiHX5cQn8o2Jd+LL/RFdbeYLWa471IhIY6b9IJ9lCWw5
+1fpiwJRJbJnESqwrN+HyF7LkE0EE/RmqYGmseCggcZnzDZx0sdeXLPqfG+/Dk4AQrdGrVqgJQ7d
xjbh0khAUHC6N5vjZjSx+5/5ZkXT2GA4fbu3CLmN3Xqbpgn0QOL2D16uCU9DHO3RNM4VgKbI1AyU
xtK6qqRPNr1qrPeTKQg+qMlljshbzk6ZXvF7eFjasbCRUj3hZ/rrGRXutuzycvsDvnDjZPxMrSkR
FCknJA8jPcN9gVNipQHyCJMxF9grc87oIoiezU6a23/fVvAjVUi/P31juvfhe1pX3285kniU+ysR
/JMo6XeFrj/9QEv962cf8x7n5WDiN7OR7LNImGqHuQxOgARmohY2MmqdE8IDjOD+9SJhw/c2UgYV
wkIVt6VcHNEW7mV/MmQHGSDsCvTUz9hyEHiYuUtnuwvAAaWDiVbXao5+jZoZFr8w10JFlvjXk9jP
SoKp6MR2qNyIkHIca7Nkq3ZrZVl/vl94iwqF0uFHlwLbdYj7nISNtlmfw2hGKOgM9eA4bR4TwGzx
abWHFS6oU8nKTmdnf+21R2kFUvLl1C6XzaOsoa1sfKhEPs9ONo5Z7bDpsDaq1BW5ieZFzpvPOKzo
6WVj8Mbs9swQXd9mGc1xuMHdsD9dLbd1K8lkeqqH8AReCRZ27T8UhCop0goumSD5nfcaPlrUW9G9
eC5z2+6+0Mhskp5tR1w64zctI6xyBlpzEy02O2hVOeXJslhWy5DRoUG3mhAE2z/K4OiIkB7XOYWp
UOyziL7ePIRESwlC8DlzpizzSZ9QDStLbuM4hFkMLnMZPiRF09Ce8B+3ycZriL5u2VVmwXOrBF9L
IivZ0UwSIYrF0yMNqlpjcCVFUmYyclbanfJQVZ0+vrC5IHbnGvUBX7aVIRxFcs84ub35uWPY/eeB
SxFRgRAUH4jBfDFX1eGYju45FxS6V2Kf5XjxmqAQHEYLhS5NYlcQmWzRBNnXnNDgtpmpzVXKZ+Lr
tei9siIWyxNhHUFapxlwUScmp46CXGPc3Bro68NYN8ShXYUY3+KgcrM6R+Kb9umHyVBlgVDwl5qJ
qMyFAt1DL026Xih7n8vMRcRpHwOjB3TusA3XIpPTiAW/Kyw3M4eelr02zFwbZnbHpIbgLlzTE5AI
+JeMs25LD7UrMzZUokrmLqNulGxNs1n2EHrxCZwr87c+nYnroh0PfVs03b6f/tQYkDmJsD80SE6M
3vGDTM00FKpjegM1j3bxGR+L9sqdNeuRiZdJjyD+NMcDyzaM2u8r9ELWdLB2yYfQCMqL3lRZ7j3Y
X2JkyLxFvolj0yirAqPlwnpvgyl8GDcGnExJ0VRmx9GcotaRDCjRCsWeaDfLGAFAvaOr02MHxfC7
ytdAj22NDHNhCwkT5k1c4jZRh3LYU5mUImgVKb1h518ITzBa301iQAjK1yLuRYjnXJ5u/07leZYS
p6bOtnJp0s6RsGkvchqaln8oTkuSmCWvzRJwyQSPphbM5GYvoHQDcgTkn41Vh+jzb9+NRhusg6Je
ZQBX6Cme8YuiIJrmZERcyvZoE9J1n8tfT7yEm+Eq2svW5Pto2W2xJZePyzsF6DMLcIFOmTiplpBn
/fgudx+MeZld3l+ZnYu6D/aEWiXJf/XHuwlQpCAi0ioEcBE/JfQzX0ulPBFIM5d0T6NnsAiZm6/x
eN8ZNLj6ouZHwQA8wR283afEOIAcwxDb21R8zHT/lPEmfzJDZhAYXvjNJ64qrDDXNCIRL5xin28Q
3EH2PUa54ypapx+uZSBr+bVBu4WLVLeFEC0feOfamRAZ2R8K/+p6QTT90mqvoHHVfDa4YaPqfYch
t3byinYUFzifB6JZT0T+ecdDzcMHeWqr8ayoGt1cuTh64Ht0dALshYTUWizDRnMC8ITo7GU1rDCU
d4k3x0Iv5cU+HVzsH6kDU1ih8aE3VyYfFBv2pBEmMFNc2DzBBvjuT+c7Ix5DNxXXZGArYkyM91Nk
XTGJQlmobvsByPKjLe2cw7rnswsOpyRfLxi9ZsJOGRmjTxMQMzPEh63heFmeRozQlNj1hJPk4tMP
jGlxHMjmU68JmrQhqxb/iiXSrAoz1DbV7pMIthlmfR7imuSW4WsU2AdA8b/2t+GGTizzJtMX0Zxc
EYw85lBhDB1DBEN83BbzK8ZrLuyOfdjLGkaF5x3sHX3Przyv3Kb1kbxweGqWrEdd6q4sfq4Ts5bV
6+1E2DE7cct1U+c61uCVPySnh7mCBSXcJfwyNM/ENxdmpKgTFuFvHr0Ur9MAwJZjHYhqr+kte2PX
/vHJXJAAhWMhEhFd2+cFyzz6WZ+QLRkcFM7j3xAfo4Xk9B5g1FVBTOWcYHbtfs4itmpMUP55bus+
zi1wshIrudfakRkxKPD8XzXrWi9mXfV/9WaahCEs4EFEL/+Bfq4FYkEXxo6L4oMdSlOaLjENx8fq
mKnUJHCic/ehYrh/dfRPatwlRh683zEFYBHaErp0mEgiRIvjaaEgPkTc2i+riNebxF8GZBWt3mxt
HOyEDzj4Vw+HilIxxPHEE8xv8701696jDPPiOJDg1Wv/WV998o2jnJIFsE0f8EE1r4nG8Pc6xqYe
7bHQdCS+gyFfJ4cMkA/ndHZHmlANiWU0oBYmbyMjq3NynflDn2I5EeiCakIPFX0YfaatzZFk1m28
MbUSUeZ7tnbs9w/WBvuQLZhgFCCaBZHL8LPCDg7T96CdG5aQyAwyXQVTnpn84C8QYOWom6MwSwk6
CsvZj/iKh9pdZ0xSkb79t2HgcihAlhyOijLxzr1Knx2zPZipIbu68DdzrL82wpjkyC39TE8NO4A4
3jDrF53bhBxew7pMmizRE1XzMtyTcQpcbf7F1pxpFqNWvBSHk41cpeTuVeJM7w5bGkV55Lax2P71
SHURmFspGmr4twdcEjKws9KvKqlScwIsE5b/yJ/GLRDBLb1JKOuc7fxo879wsAt7u7BC//bZkJzI
zLLHW5hBYtBB630m0d+B47S/eVrzv91R4FXhIULo9cFYqa+6vERU/EEPh+BJbdLDEHtzKRZ4GxJn
uSqurZ1IrYES1xrwUNIPTOYPXyxgIn57JSt6ik9VELVznCIMTv8o+9TLI3AxTdxliF7Bua7yiqNg
4KLJjifMWxSJoqdy8f1MKIRLyBUc7EcwDvcVMn194zBd4DKbNDOqxiX5N6B8bYrswNfgXlkkpCei
p3bOtCF4MVzScVlKUUcjvtLOjLnQVw5WSCmTXDcC3IbMd7+EHSJ7gdbObpU4tlfxVcNBmzsy/uUw
725+t7YH/9V43RVepG2z+i+j72Dq7aezQQ++Zica5Oa2TqV30LUldQK2L/xbZ5awbO93jyZsFv+L
uj/sy7hQcYswoohdFsoOM9QlTWN4Q9k6W9cBDqZDHtzJTEihvjF0Gs1Na+5cNAYzsqHDiW33P4Bf
M8jxKmSRlnhrbdxTdLoH2Oazn/h1+gvboDlp/82KY4I38NqMIW3vfVsZtY+YeSJYN49JU4+KJG2j
dZJke+DoA8qG4S2DW8KI2OFR99Za7WXyLQnAQLY+NMAEdT5iKxcgnvs5jhFA6OZYrh+UVp7OJxS6
fDcOSJRdV/foq3CPMSPwuUUJbzlHaLsNcmHltX4vAWwfYFQzcjeohYN8wtmPWzQtlHY7uifyA4Xt
CGS8uO9k+kme/d/NSCHoppsnm2HyxOivz8/nc1MxW1CJKE2xYZlsKiAT56zO8diAt8Us9yy82Ln6
5HFGtlgNMMRHc4HtkljtbwhlUQ5nZowv3dKqTDekUisdreiYkskm/cEMFlqevtMjZsueZUSFIyO5
Ht7JxybFOL3amO8nAZurS3J8VqVOrlmCjFY4PGdN57r2myVun4vphpUOPnW/gvs8C+t7xSQYr9oZ
7E3bh1GyMNjUoqTFwqr/2OsCCYhLOfnwFd0IE8KwE6nLy07EzNizUibf498F4OKa34YWkCS81aaE
8PNLD/X54EUVgn2YiqmKvaqF+F/uHXvoNxwACmjsW4bRmbfBcBgToyCylPNhF6UCwrPD5SWt546i
M1WVHl/cJVZejswYBTEQYTvi4GeqmEVz6lYpDuEpw0kF8S5R10/yLR2E43wPS0h8M6q6rhl+2Hbq
lwwntDKLYFmTs/KnCz77TSYxdQpKx8iR16z15D/ysGMea5+PXa5+GHrKZyAHhsUDLawdu7U6Pul8
RAi71LAVnFUkUIi8lGukryCqRmxnP6K6aGVaLZZSxzNXfu5hrOh2/kw/ELW0GpJ8267P3svqus9J
QcRGbA73rcMkzFCgFY1YRuNW7m8yl8cZ9GJkNxM/9UXX3Oylppg2WDo10zIKNs31LpGf1hQwQ2XC
SiJbBTUUyAZMlXMYD5TCFBpbhs+wdSgs9Nzlgyj9Hzjh3dsjw3HE9wTJ046LiquqzO1gvbFeh9qz
gxJ1HWPi5O/OYVWfn/k0fLXaICcgaDupPHr0AlrJEp9Uz9Zugd5fhvCG14zEOAONnlXQqtGMa+AN
kf4slNUZ2aai2zW2nnhQAEmIG6btBOeX+hTTkdGXovGoeyGbG1ufh7PPMIZSZK7tsysy/HqMjQVg
oXAn2JI+69GagMs5cBpriLcSAzjz6D7XLIubvGQE7OJnKuQ9LPVFsZo5yxY7KRNfCOo6OxY8Aq9d
6AN7KFFJk+sl/fVvcuyZs4zDKyvJVkuzu6wXmf1XguvgZnFG2XMrv+EYqsAMWaMQxHECtfC4Spzq
DmjI8BXd1BNhclts2u1U5koC5oLUAX4pSnRNwknG4CDdN9J+ey0GCAP/CNgd9Fp5jaB/qFx4YwiQ
EM9bQ98JV6D1SN3Zr8AUtMzL5dDE9dfOL8YttznT2ZXKxRimvv1c4C9baLZEdFNrIyyyiDDGV+Xh
h8ZShnNO6iuGgxv7sM7hANrneg+AI5QvrpINEg1xvD2nQcUFN7zt1KijrK/eH7tZyaEIj3fCiif6
I3yQiRylFJHxmIkuTrGjk57ZtbOTNMM5twtCFElIwy+02ewX7lkyHHipOuwZHH8+V/0eCQMy5nyc
DInabGRQYm1M1GVf72eo5sjdEY57nrR1ZkiWrNuwLxH7mslNKBK4WPJDS4z0JsrgHwLJZcQAK5Ty
C06ti3d4J8fKcsmBGRbVF1E8dCdpOrVqpvw1+xcOhn2quaKGlFVq8MjCHSTbWJju0lW2o5ryEf2/
IrcBI3eFvLn/i9Ovno8igFU3UYfy98O1XznuJGY3GlCOggFmPH7rj9aM5Yn+oZteCyWwsy+irTwQ
YWPGqn0f0ZQ2NdlAhochyaovE0hPYc5frQLh5HOiAu0uBEJvFownHAk14ikxM8G+E6NNJNo9N6t7
05+8y3fvonNY3aTyI1IbVILdcb73zwqIJR68ZROJW63KAoT3bcP0PxcQTqAlpghLdWLJcn06Nd0h
bgc2I60Ayk1P24Ki3UiemtoNwyKuqqdmTv5BRD1HhlFFVt9T+H1teZMnIKOVanOlqf3sLfxr53BH
sLHIJ0aVLl8g/NP2gAEl9PjY7keOp1TZ57UxPOUO6Ewg1SBQjNBTpR70XTnQAJV2mne+Gl5ABPil
Lc9UTZfJiYw7K2kOooY5/R02Yx0WYs8BYyoP1lkXQNNVtveRuCivSpCwD0QgyATNGO0akmrGwl65
ClOBZC+b1ouxCFGmnuF86TUATkMQ/pHyOgc8FRrWERmDxEQ6o0h1qnzSEvqYwSiIrXYJiKvYlVz5
HFX8zrjVk2dXEXmSANYuwJIxa6UOWtVJqTCT4FLyu0+DvQKB60K9q7eINoMbGxklwg9X5LQUtpWX
NImYs4uJKLo0X6w5LyGVK13yqnVIolVUCiWo0P7UqhVsWWN70Q8rTmOKf6FOSCRfw3HFE6E+6fCa
6+jq4PAz1LOFadaHYxGwkvi1r9C8bLHPRRMxcSAq2HyoDtBVF+tSrJwdc9RhafP//foCaj8Osnkl
4i494qXJ5Mw24ZjcGxU2+7T5tpiUR7fsVHJjdmJPu+uKHL/SJVy4zTz85uZEngYQGPJ2lq/deMKx
MnPBfpi1EEEv4hYkZqZnQhe3CKY0u01Xy7A5uTW46nL4JS9bNplLGZI7uqAo8829R1+0dGkcEsls
d97oCQRnYwglhM0bGyAfnQKPSzKVXsN+23AP8adsT3MAyHkYHENCmokWhOxDCchq8uYWOpJeqO5u
LSfErlJbhRRinioafzJBJs/KkLcAVQqzyzvqUzSfunAfjepsoBR/3TgK3fxS7K1YPWCl/Chn9XNx
pjAU0FN7iu6q5oKNC1s68yq+ihoJlxHtxgQK13dsDm9Nnc7BA7eZcwTBJLI6ckC5ZP4wO6xHi5EE
afUK22yWr85V5D2UhsMOMLG0PT0UIbr90VasCS15z8M7Zt9XqWNgiGICcN3Pjr3zo6gG5tVvdtWW
ZVRIMUB/Ey73Lc0DxxpXz4g+zDrxKuDdsLTNCuBuUNb8Ug4mqol45hA3wPE2LZOg+ylBxqhWJh5A
LRTQFhk9eXWtn7F+wlOg7+WwdJCbk04PfTTqQMB6xhXq5jm3Ysp/jJPBsxJKNCqkolY2qgUefd/5
UpC4JrcgLT0PQKgNto5gxP5P3KAbOYk+DpDvRKoKZQjx2rO27UBKs/RlKuuLVMrvSLd5xK24XIhC
VPTQIEKxA4djnVuDmtglzGE7glL8mqwBvcDswI/9wtv5TJWNYFOp8/plfaT3XeO52ClpogEHMFix
WjOS7pKc2/PkC4s5rGmqo/j0xC9rTvxygMZwePmqjGb4sW6P1uH2NiU63ZlQUZsEDPjMhftUMT+V
1F81+jdWTwX5TidNb71mfCa/kKKcWRziMX6GBxmyFB0bY1acAPNpeG8+cxOTWh8LZ73NNf/+dFg7
Pq6Klo1dlMZl948+HKTG7vEWI65AZUkoMfakque+ML0lZffw0VUHy2K1U7+py8kZK4zdrxtw7XIz
6R7DMbnHV6gMzX0fzoFUIY2e6RwC9VqJhizf09uYb8HE0PlK/be6XI3hc/QCcx8WbowlDPziUX9T
QEhnLGnmAUekWpbCMqpDclOSLuFYqDtS+DhNxBjJzLRD6+fClizX8MMW/7oXs+6uyRJWcUzlX8av
r9rzEzWkP9EaoLz8lL6NWr7V7xpXz9bjj/t3RLSHACinKivKDp2fw4xihSa1Z/xUv/3iT/xrUbq6
mhnHLArlqv4xOZuD/EeCVSbBfDJ27myKSC25TsGtWNFF+pLGhaEMBvFkIKJBgfaswH+xLcOVs2/P
WMVxtdpUa2uSj2u/u0OjhGTxieGOgKWUX8VntGdFjLY4xEMoDXWb5G6AHVYGtmv5QTDYTytA6bjk
olzgsiJECxvzeEEOHr479TmsgOjv4gsGfLmV67uVtdj2TaP7sT0aiZl7cXBQi5sBqrp4gMvp6LRo
E5k9DWMFe4p/8rCpZ1NdGNl8OtTtxTIf+OycZAKde6Ma0XlujMQf7aORpmUGQ/0H8hBXdTVHjoMA
5cpwMANPD8Rk3lJfnDRhajF2gpN7HS6TVxOW/9WUhoDLMITgPoAfbs8d2iImyKcrrnWgDhXH1UMs
xyvDESoUl2jPByHvl9ogQoAT27keJiirQ2NcUO8xGqDYDQxfPa7woTy0zaFpzFJiZ8DtAbKY5Ra0
S4ieUPC1HkHhL2OKen9zc6eWTPoyd0BIIcK6GpEPxobTYQiDTaZYbYA5J5MR9/ZnEenDmIaukGh0
Q2/QfMSVCxQmVZl006AOl/EqRQEZBxKSZEbLqvm7r1ESegryWUcO4CDneZOwLUk6b1XYouyDoUeQ
fZloFFvcSVJDnOCdo3mRd2mIle+9nB/RKvdHmLfdzYgrhclcoHUWC5ZPWdouf2WF80w4YR/Z+Unq
avogtq5rHlDtFb/DiOb+BMXhBBiex3ewqtfDA52DT/ltofi3knNLIcp9uLfYk/2ufzKXPYY5GL53
cxlkuXNWlou9Zo9w93OOVzqQGpjDT+DdaFx+c7yXM4xnHi/CUvtSrFgALknWd7cH7RK1KesKyifT
CT8bD78OA+wRzmhsUXIt5elLE09l1KXgTA3cKcW8Z6u5E4bfIPZqIqo9Eka17xip7M3UtoPsngWy
hL5GrwOIEUvm/nM8l27Z/iCS2Qpm6fDwELWprIrpy1O7u3kcByYmvf65KKW8SvwRUTrNhTQoOvQ9
y5zJUuMFweTcThm58X9id8InL32MnuAHbBrF7vLjP+v2ld8KPM2BYosGpunbuwgc5vQP1WboEFG+
XuYnbk5pE1gUqlc4hf0VpdD3/fZNnAcNuH3BOGQSUUEPDUycdFeAjlcO7HWucFXnQTYD4dlBPdqf
+x+f9C303As6jrYVAQZW4fvOklAG/v1M9E7B3OK+dKrmUv7U1phlXVX0LrkJb9j52aNX/0xa3oRQ
FMdA3RKS8SVlVtivyofHVdTbheb/N3/1PERqL8nn6z8PQ7OKagF9cRQO353LRSMxrR7HaM6LI2Z5
LzoOrknZ8gKwE1cd4nrLJvheTtWb9dIyh45ycwfJcp9d1b9jVz155wkbpXxmyas0BWIgGV+iMGIM
JB0C+ppq2M7IJs9e5ATvCMT97xFLUdpkyjfy9ycdfXU8W/y7bux/nauiLyP2KQTi0AAs/I69H7W7
qT4WzJ05qZ8mijLSmyDuX+YuREpnHad+WhyP/rwdh4nsUw+9pkapdz6VXmRNDb5I7AJNfkXkvfJ6
+KMUJdRBXxyFhEUl0axZk7NBqVAu9HFGwJUS3t4w81CDAvNl0JWEMMmgGoxNmJiXp+ta7k/ERPg6
6r3OH+pY9HPvHo5i7fioTKTMgbraPJoJpMpylLbDMha7yiAoVfW/w9gNhOF6gU8OTxuFOwc9inRE
mdXxvq2zbevkxZozTHxFUlfSzODPBBpjPlE+1boqPlk7yo9BVM4tyKouvgCnLWtcD1bCpW22+KrB
HjMerMWK4NiNR025Ll3TucZqGygvIpKNYUST2pzDJzIH2QXZrSXCypZwo4yPhKYnzmM3x5uUsuTd
0KLm2XqhsNTaDL/5nVxDt8XJJe2HQcqiK+mY1E8HZujdQHPWJ8rdL08nwJ/3FJOiHtOrMVNWWGSf
CSCCDtc6686JAd1mTCTNwkERMHi5ngzikUdPoU8vBRmbZodgWE2n9W3WHT8AVU+nt/mYnQnXKAq3
si3xbfAatoWIpEPDfM7gvjyJhj2H92z0UzgBrPjVIPnymJ97heFqbb+KFWfK1fvTjwsWN5CzZszS
NOXZwT7RG7DcA9wEONk0yp5grR5I6+mdRLkwJqOE2DJAiosgNBHnbTZgrS9waUOTkO6il0qsOr87
Eo9OI6KDpv5THeDmiEX2PZ8gtL+CsuBjPzG66XygrL1vJxbB9Uxfng6h+ATisBgMsxLpI3wgcV4S
TK4K0dMxkW2HFjuUhl7ll/iAr+2uaI1AvmiWmS1ZmukGS1fHpTMDd0+zVGliEWdj8x0DAhsS9Wei
DO0hxVD7bBrpgONbzt+f5z9IVZ+w6yF1GO6x2UY9d5fdZeJpN1FU0FL+vQMxkgjsCLuIwOM9AH78
fiQ6uPVR49ddxbJM8WTYI9QoGG/S6XSKNc/PFOWjslAx3aJoW3b4kq0wffo+Z8Ov6gLOpR4MHBNT
m7QMQ7QPMEr4Dui0zusmNEElb3RnH458BVKLyzTaoT/LMI+0URQ8ZI8aopIgE1amCZQmGdPN+zm3
GFdYxgsMXHBMel3Z3Lr+iPqgfuzM+AeJYnbIHH/YUeVgpgZSy9Iw7HSGwY9ntVpg2piYzpFJP109
WS4BpX6TaDh8to2vxuJ9LhSsE3A0KGKfkSRA+4dfQ6kyvjx+IH1F2vZXpDh+y26Sqw1Xs856nOWC
eptIn6kLgNL1i0McLqy8NkKe4ucRTGQWqJj4BntmYlI4k1zMtHKEV3lg3FS5Xw9cgNP5UcWzbMEW
u4BbGC8klQE+Z+2v6RmVzqhH3+XdoPcKSZ+sBnyuupfy6jJ4KkQaLmPjHgZ7kqMvQ8y3Nobjzzz3
9dz5YOiwntLwSIj0nUlHjU8LUUCwowlwu+XHjcmedrSgqXf59+yYxkdBaJkczD42FdKNJ4MnXem2
RXEPCOP+1JDEmz1u1HXrVOp9Q35ULLwyJClxN3RuPvnHNZlmX1Vi18RLGhlM6gGqER+NlqO/cwGp
2BvkZWVzHDn5EpO53HMiJrU9dxulyV3WlNZ+MrZPU9XiLD/8otQYiHL8pFQDRUoKSUJd38UNIHJe
K8ZhFGOCqmCm7BMrI8Ll08E7OHCGl+oQUmin17cu5DANsHZm3xv7Elv7JoGcgTyGlB+WFrpzvCD/
LXkPEjOyH+ZAbO116KrODWiWyF50mOnVIWIX53Z07ahhl3rRiZt+I/16DQrz0eUnGFBtWRXKuYl/
KGOlfgtEV1Uz0uph+d2GQn07D+P4tZXtPxCLAfNt5281x3ANTuEyLPTBuu+XnoXUX+1nwWx3EFha
YBVVGSN3ggZPtokolmbf4vbk3mduzVjmve58Kmz5EygKaESupH8OdyJ4PSb9ItyL79DiJTkS7lJy
f43KGzLlxV5/MrhHR4L1aT/wc0uC20F5M2FBNkINcQ+4LZ0MZoNuxmEOjnxwn5RNldec7yv/7/HE
0xYlad7a38bCeff9scFWoJAQHPX/ccjxQVyaSXvws/0CKRegxE5zkrDBuWyZHDbfhlLC3o/u52bg
ncy//6dmJvob4mglTwhhgbt2BrhI6EDiGZfX6JS9N/4jSq8JD55V4KPG8Ae1Ae9FlxjsUDYWLq5R
IJQ56ZMEdCqft3M2frAcTrOecQ6yiz88Ve6cqvT5fw9HhDf86ToPXrNWlxDgokNU2s8rUEPTabMo
DDlX55YP+FC9N8qqMlhQHLs5nMlFT308hqdamI9DSoUaxzx8Up+qs38YCYbVxnjpYGfJhkYIK1OY
ArEIcKw0EfkbEN4heNoxzstScJRg3lsB/zkpiVi2mWch+PytrSOapiO2dElEx4fuUpQ3ZDY8gdU2
BaEI7ADfOKAD30YnxBTbvpnHATVp5QGZcaxbwUjkdodOfukL1OG2fCCmyTLQKt5KGad1fpA6jNkQ
cPJW3QxaCx8fLIPZb72IqSfDIAaZxmMmJ5UQ9LDt/poSCPDqTootniU4SH561TtTmjZhJ8mJQAdr
vqcVmW5nki/YjdMLUqAUdNi5zKvZ0AKMJQ7fXrMkK7UNIPkksW4HvgYbsuq5QXLlC7Aw6kZAUC2d
P/Ihyb2KZpLAcUGnu25CYWjJGtryY4/RNKf31aJns+6rzh4fsQOnl3Jfj7AIy5tGe7SOpVoOVEzd
bstvkd/Kn/41VeYFpg/22awGEWlyoJ4CWFvC6XDgyPYP3C0inlX5jsC4azI2cv/negl0u+UZ1v10
me/+dDqAr2JUaQ9r2ivI9J+2lvzYJUoFPiqls12Nqz2QjumtKBQIYiX/VZgQNdOtMzmeLOucy72N
QqHGr2XDUiF7zy0OyPU9EaBqQIXJeBNzw8pT0bmlbYzkHE2s+j6pgY/4ndzoQ7aXs9q82HbkKba3
YkIy/tuZUVw2LnkUA4iANHPICjNS6kpxRY75qCsJv5vwStXbPclhECK9U1v0OPwExmP3HDeg6Fhh
lKCcB/N2uVKfzS1dv3TAwA/Inf1+H3ox6Pcy7dyEIyZQEfYfNjmsd7HMUXrtl7gHYEa+elG/4eze
mrcHjUI6i9ZS4Ab3ymMGSoKBQCVZ6qdTptSmADm+LxROzGuzx4WM6RtXK9nkCQaSrTLRM2UF3ZoJ
htkRbPAS+CgaFngWt2i3Oqxm4CGFxFixxfGiVBkFqdQE/4OwWAtPX7Pk6weIyIFL8SCbGZZ4IlzY
7crRMLxkmrdfpVl8bu5AufMuOrABJtqI4cF9+ULTsSaQX+8wTcttzEVUxQXi0W4xEZCdtz//AevK
hjFwNrf2jco7N3K26NYfSR2AlblsJnw6A9n2Gzp4pAK0aTg+fl2qIWfpTkbPidsCl6NX2GnhIVSw
lu9/4NbyUkzsICt345W8+RPZeITBmq3zJGmQjVCIAuWV8OTlGiPDv7gFJ0Or8KVBCjP5Y2/6XfnZ
9KuK9i6BOgkoKrJEtdNJH2lMcOqgNj4shDBV4ZomOHULXD6cvg4Gwj4jlMkvnBN8mhSAx1Swer+N
wqGiNeoI6uRGAnjLadNgoWze80MUgQthKnT6qmQdVWi/cvt4wLFbZvLTgNJUXijDba16bgTOe8yt
ARvFHEWYRx3xkgGApyBfQ4gg+EAQKkv5xCP0QJZa+f9VjsPIbU9vELyCKZttAYP596qyb8lKRXi/
XpLYrLFriBUb4yJKEirEtYuCSuyhj/OOe1yTYiySTFRxnCb4MXYCq7wr/rVNG/97AvzqkSfJtmh8
CQjMS9g+D8fUMSLJvJ3UaAlrGRxWKlm8mLedssAT9kY8JLQ31NOgeh/y1FKQ41Y5JD1OeukPEHVb
eMd2NWrXBlyEa71kQSTSQ6XLbeO98/NxS4LhPqMgCtTffxtdaacnDj7y5un1fm3xul6yT2QuQTqa
6296ARo9rUodKqeJ6wC09VBin+rAzskLrZjjjVmtmVuLjv9UIYoP3v2i2xcxlaNmHSV5mk4ztrq6
pV0kNayLwvKS7tkMiAix0OE7lCAl1WybjuE6Kn6OndmmX4DgrnFONjRCGj7sGkNW0QBHuQPEyat4
xkwYwFDYl5JzMCwyZcDrtJ27EyUcthD51e2DKSwqcfhQsbO8ej5G4nuoHlbuPrtmNHGKZb69QiSB
2mfw9vDpQwMLUwlrto/9G7A8MGXJGT2hYy2LMxiSDryeKS2BbN1hYo5ZmBsiKkNcExh3ZHc47WA3
RS4ymNaK63Nps6GX0PepwaYktuekAEhVv0uLyu33PIbfictBGV6X+jrnSMga32oRLzawnQZ9ym2q
f01DJC3dnve/XGDVg+JDshFdFIJdU3kuR+VhFht8iTa4GhQCxoIOFDMNy3Ay0HxoTMQCQ3bWYtR8
vQcxJUMA1saTVp6z7PvmEYVIER82ppIdh7cJsvNbzgMuqaesOSsyKHDgA+R+rw11epD4rRbgevV1
GZXnmxMmO1bA/MhKt/oTpK0iEGTpjYEs23DuB13lGUV5lXOK6D+NtKrsxZbm5f8F1riE9Jg4yIjk
rVkFr5oMVMd7tzqpnjc/AmGDGDlv2Q1miqWsyaZNa/ruca/NW9aS/ul0FJv/MrPThmp74yTMKB3A
082t19cZoFhAVh2Cc6KfxIfnVbqenbXc+zxFL0zo0c/OHInW75rZol1TRel5lSTJ6ckT5TcuV3Wk
6MyAlyN7nDW4H3XdjPw7GB50/I3D33oAGj0zitMqaZLX2dfD16qFxNDrA57eY+Qh61qVVa9bRINZ
VBAxRTR1vk9/0mOYhyHA6EIPrJkNWCH2CtXuipKyWWpdMS9mpJZeolOJInHTd7x7WD7eyMlZtGPT
v5IOSSVz99DCFHEp4m0BA/X6Mix2TawR0srts/qHh4kRGqndfJEqJV9OGRBjPge+ZdSNP5GtNboF
LgiwQ5JV/78XtsGh/nCzSZgAIXXwuUQBT5bn++O2MkuhDb+UdgHoQFqsjIg0WYXchT/Jwjj7AfpC
rtbHcEWpFswxC+N7TdsB1Qa2e4HX3DwH3PvEQYh4+Y9SHZCPtRfBaf7NLrOHto+jdf4WszMtY1wb
7mkv2mQSlQatnpMwf7I2Oe9Ccnfg8E9S1DjzH5C2EBFE6lDE0FAtybeNAUbAethPX7c6h3h6X5m9
WUSQhigfJzvne+UMRLbt02G1nhvf9/L4wkJCqLOluMvJngqw/XucrGIhdg1WSew+uILNeZaoyucd
UNJ4AOMloRDSoJl9avpGkKR7n9JZX/rMv0aSEsNApfaL8zjGC/ejzb4sTl25pHhMLd0qJLc53ZgB
et1L/CQgiTJHNouqVoACP7dR4Eh9bTbDE7LCuoQghYozGOygFsJIXKhj0Vr6/Xry5NNYP15m6X4j
k9RYA2P9t3fFB7H5cYv9aV0cMhmFlc2u11R/ZHq78gbRyVSBmpplUTYZv4FQSdBPZALvtLhHRlFH
s5sFfcJo4uo5xb72T+4KWu5Qj753YT7teaVKVT36z81wby/g2OB9a4FoSnjAWRQ8kKTbi8XZjaSI
nXPjiACmX4q2JUS4CEXXZubYSl0epzv5l1alXQHC990McarBaB1X7QAIVzBAe9BQ7Qm/HyJ2au1X
UYg1zr43SY/2Ujb6mPOqEhwk5cB1S2WtIzNIk/TnfoSDF5avUJa6e+RlC1ZbtEZa5lwt6phHbEyR
VGtymt9GvGb5nQ7SDHP/G70V5z1YTkriuviT2krmlLS7jelQvh1I9Jrd4tuuqK86ttxTAN+PoMFX
SbaD2J8z1yFxM7E1NUwvyZ8Sn6eAq2jZDyqleKHfUuNbZPHeOC9Fwzs8khJ0E5AKcMBzUXpEcb13
Y8Gr7R5rnJOVbTrYEu4k41URBClHrVDEAKCL00QzP298h6SrQXd/WoqD2scVdHsSAdrD9BIfkKo8
0f08lCUP6dK7NvNmGDgVkz0FmLH4+PEvUi5x3NlssoqqxQ7jYTsnei+57Qpan6TKCH8tsIhgrLsY
OBcKpDE8AeVgBdQ/2KvK/xyvDDxv519uyHGlm+J9AgHp7H51m55fNogbTKwfdWsfjpKpY5VIqVP+
PyRTbHE7VLsEFSAvQP3cWuPG23/wDUtIpkfcKuRUIWFVKjVH53ey1SQFFYqNhkvtEhxuJWIucxYh
WBhg26MuuVGOrJ68vnGxcQm0leHPvBHV75eLGAGl77BD4Ag1Wl3C7T9XBjo=
`pragma protect end_protected
