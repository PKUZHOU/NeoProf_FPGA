// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
0v4+sY0rkqCPhjurw8YDy1STZ3ctg85cum87eV+ftJZr/774HEIwzUo8YN/PMMYxwNwTWMKK8Tum
VNPj2OeZgvZK8HN8WyXVYv6sIGgY5+bXJWNc9s73hATZodNWNoEq7wqB5NczoXAOd/p6+X2wR20I
x4yk2B7vwVD4J94LsSh3yPADhUT3g/xsaJDJ3KzjUcLdFImjeM3yL0Q9PvpOYhxqqVLCz4TLpL0D
LprjCIzM3gDRorzNol+/JAk61HBr2aBs8t6KwGFglzZ73zvWyOds5htcY7W5be8CGbLVefV3cjSF
en+wlTCSuZA9OyGyPCKgztsRdTa2lKLY4aDGrg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 46352)
699m3T8yrvm7HCxELnPfYR8aXBRZZEihsHfeSHCstUoWI2kcTw7uB2ddl1WwxcqiaDc4njP3S/iE
PJ0k7btng9DqVLrUAgZZ+YypJ97O79AFc3CCAuIZPBjqrUk5WOHxXpJGHRk8AzTboD2zFX5GxIrS
48clC0EnvWrkSDmpTRP0/kKxsNGsaGmJ0S2OzGXoQKwgO8hUSf8iffsk+4rtgcTItNLbDWn878p3
08a1HTLyTHP/hALRdBGXt546xjKFvFlPagyZc9GKYfW2HLcJmrIAHFrsS9n5BRypE8ABEOZHp0Il
3FTtpuKK/zwc7Aj5l2yDP5wCXG6t4FQ0BXs78KRvxH3RcBLIM/WnGkLLDUOd4Hke0ejbfCjWNfhz
v6WxDpQ6cJebS7Jut4n8tsLpY57xARzTf2Moo8SB0+qh2L/+JvCD2inWF4laiKT24Rbh8cBHZxLf
vlV0RJ2l6+PHdSaaATQX8xwpxzH4GEqcgy+yvRgnKik571piMmR7xzm+rIIIONTccwgaLkKnk0ap
9C4JmwhmaCJYVoHUWwpRtpbuf+b7OEW1Wmik1c8q9LfXhWPslZ51JnoI3ghW86hIMCDvEzdFDhVj
E2pNlzXgid0+WOPOKODd9NYD7WZep1+OHUTifirVvVn/iQ6ucJ/FqFtHX1ezOLOTDeQYKkuIRpeR
QUTkHtcmQTzAsPzSmdhLiGO8NceCHlZxsaAypvIB+nHz2FftiJhxNSpGkZQfksgEurnrnOw4MjNC
jcosTOGZ+u9Av/J38ZkP6htB2Xm0SSCzyNV+iUO1T548KeVVTyM506i4nXuPiHgPTEeRpkLHOium
dV5ZT9C3fVxgUAMGN5mt78Mwdt2DYrORS4/rzw2AFFWu3dPPzaO2UGXk1DcAW4j0RM1GZrMo2aaD
nCp8Uu5vlXzYPiVHZxVZcXpjdmimpLLDJSUhRxRJLAcpm+IbqAhidYlkWbL0BVM18tjqTEh0E5Pt
tDP4ASVqTVASbm54CbdynBsZ7r0an5/2dqOYKcoAkcG6ZSyz3ocKQDHG137tgVDA079fD8udr7c5
FBmn1TGg2M0rEyMTdKzD5vJRITyrLAYejPaOvOD33JAwA6Zke3HNXaj5NHMUS7ISNGoLgHmi50ep
oH6rkcNwqBfjvRzmtKwYsgXCqAdqvlVUIC91JhpN0Q0geuyUvo1tAMi+GOi4rm0XGmIDNR47UzA+
Dfl6lubazw/QfqnUuoDDWe0oaPkhfZYWeLyipHvqE1MX9nPfR4judrhwr7fhofihGBRwyqPNS7CV
DVSw2JGVlqxwyahCdxuDhAgy9DgwHO/1q1db1S5ObLn9KUNa4eVp08yT+d7Sqy9ClODALmKkD3ea
Ol7ICG1GTsJQUjSaxKuKpxTBXO2wVjd6MWpLsEaU6E6aQowfkn2L7kl5ZZ/6orMA18lCnw9utp3Y
tHLWob4jKtEuDvrusv0eT86gb5o6s/Za2C1yMdBxIdOIKuXz1MXPXGO669yp69beblFiLGXUhx5F
2CwZ/7mLk5B/dNMRpfGIL+dWRzzdFinfTlcMMEvOASBzhIbD233YarDudN59zjfa7bG8fTry5VfY
yt1BjVUayJOol6tlTVtsnkxqAeAMXaH0biAZ3R2WS6zaX+cfYvyohAPZPnTbXgOZ4kKXDafg1/Zx
R07qgQAiaev2LHLuzx8hYO2x9V2xQ49qrAgTtsSp43EHRqE14Is67n051KncyNQ26T/p6WLLmdwr
xZJND3a2zdshbKmn9Qy5fF3Zf61Zwk/bQb+hS3J2lroAqRu+Tbr2Ajyx0Fpw5Z3Qa+PNaXHtR+1N
Pd9O3OJtReh50sBkV6TMMNYnNP126YM8O8VYU92xH2zdy/0xgSedKuqLaS7ZRrnaU01iA7Oe+6eN
tntW0tNf4meXXgO8/9Kk3z8Gk7mx77UpBbAWxNc5naxGHXsqIEho5g0rPnj6jKDQJzUyVZDph5e/
epyR203HhfBj1lOK2ePOGPaUqcutuEiKmC06hOnP55qoA7eCo4oSVtNG9T0F1nfp8nNkQyAo2JnS
83lXrKTWewUQUTDl2qN6RdXZfPnbMWMCc/hLbZzRls2hPZlqgd1/uue1GkteyqzDk6xRS/0+MNZq
7DJ/yydYRfFGEwgBg4z8f0/ZcKlW3NhAV8gCzRLWzoGV4ChLVefvv8cy3midhU4zeoHVTlSq+R6/
UpsZ1S16jXYSDjerYR9udhzrObop/OXqjHH8NLMdQdUr7iKT0boStnSznjGzO5dXwodlAgOdH3GJ
PXbmFZr5Iht3Ygl54iNHCHXi3/z8xJedJwmjVQsgkr1a9MW8xIZBB0DzTY88Bjpqc2Pdz9t8464A
i6bZrwEBRBMKtMj03dHOt+qTOs75uHxP9ooBaIWrGnzdT568HX6Ue/q9R3l6S46v88SJKO9o1RJj
RufAVgkGtf6NRbkopNo4uL5fpIc+HFsWULJvEtPnoVZnP2wFW9PUZSte70GXViK4jx6wo94DOUcU
FO9WZ+wQgg/DI6j+56FTpuAuv8HyIoVg9e7wZLzP7n+jdkpRXx82vuBzONeDVJgLWV4AFNqffJrT
1ESgeR7VYE7ayWeazZoGHDLGo9dxjySSTySCV6p/XwccWLUSiD/MGAf4ddVbCLF5WU2Tj1SEQZgC
E/TildY0WvyQZUgDCSIzsTGT94J4Y126ikEp981YLpR7nKxV2vAszZnNhVB9YMbj+FuPsaQeGm//
1rwl8SrR91OiXnM1JetqQdigdDYdLEJ8FQhyp8EFusAE9oOprrGPn6fNyh6S8mKCXsF0qoZcwf7l
EAd+9RWIsYtnnDLL8knW3LYnI1/hi8yJlX9gG588ZM9DaVs901AD0OhRfrJH9GRPJ5eHozQScASo
fJM79OOzlAbKIInY6S0K8Mcu/T4Cfl8HkPk/vdX4MVlJ0OOhaedAkLqDhYOqqbZv5rCex+dCb6Jf
q+Gi2dwbN5COpDye6attb+7aWYgOE82OCJ9+OXyGmW8scUvcrMUzEzcZSv4Ft2ZQvsz/uqD5RAWG
dKF0liQGMVYc6IJBSNGYQ1EPv4eSkAgyWdsDcm2sTZ+oajfhf0P0F8ZiIG7RANfSzkTKTOaOVkim
DJCLLdhB7h8VzMOOohrgzpcjB7Kn/OOTeaJT2AcC6itxceml4eZSB6rkvMedYB+fZ6dMMRCwRdxv
eHYqAM/A6yYGfWsfia5DWReI5AFymMvNLNRYRl+llOrb6qTJ1Y9xUC98rrbzKXlvuJD5PoA71MR/
v811HYRkhmuMH1eHNQHNDpr8Czu6drK4Pa96T02tV950Sjv+s2gxY7R/A/z4xQArMct5AJQPJiyA
AEUQCoEXfBryWuz1DF//iWyWPAMGioVt2gmjNdFOnrIRQNmJT/hz0+lqmAvVLe2qGeL38iVczpxi
GNvYNbMfUlrfXfpdxuRE3Tfs5s8oRt9VSF4euqg1b9Fbprt8qnJNsrAl26yy63o5lUhsrpA8H9I/
4E1XKR+KUa3gBBqRuD3TdwPzegx3DnmjvMjfYNRAiZTnCB+7UzGFcsOhACkm4AQah5157b3sqC2W
sFh5L1gtSU+CutAJ9B36kc7rWoFb7O4QIuTEQCdjTG3aGektUxG8GEo1krAGp2MWqK4UUqcuZjvV
BMxkoPS3VMuSC7UdDtcO66btLlsLXujJvE89wlcnDLIi4z+6cux8D/ljE8zuNuKEcj/hgnR1QeRp
L+wJi9tUezypEujUyxD9lWCXu5MOa0yqtVA3htAoxVqg3tq9W4hEpQ16nVcq8tAcpupA4vKU13iy
XY05UdGeZAi8/fi7WaJ46AwscPDTsDqBMwWvarTeJP7sfyyLee2q4obRLZrfk0QcWRAznQ9cy9oV
HPd6ciSnvaLiMUv+4I5poeiLL1C26KGjKK1doh3C9Y5tSaaRcaaTmpkSi7ElClz+c0i8TGtjcqdn
clILX9RMuqvI9CmKTsnkrxGPJ9ZyjJUj/28X4fE8yAipVFPQCNgX79J4I0ST+DtVVWI+aZwV6itM
IKBn6TjBJIAmo+v2zBKJtdzHg/aEE9PNX8gJvqlNXkiZX+hKgAVGnoQFp9tTlJARJWH5W3Lux5uE
hHKm3GUy9bPEhX5DFAI557ivEsYJJ7AKQWk6dfM1uXDF51fhEv4JrgLQ1g2ZMr5Ob2oKPQJNfW3+
cn9Sks234JJR3Xebh/gyHyO3QzwNMLWuL62J8uUlllKEHURJl+IeaJq9y2MMyldwMP83odqr7gNR
8+T/Jb9IOnEIk9DpUHmi1ka919dHcbN6OLlHuDpVxwNPnx4fPYDsoiqDdpepfn2akMdMPG8d3ked
Do8qzp5Chwi60+96jMPhel/qEZPQWsUgfEa6xuzRI8MJ0BiC9z37pN22R5ftQKnJoDXB2PIXqFen
6XDjg+zkb96OMi+Gw/j06x5AY0L//yJrUeM4ZvQPrCzvVcxQDYkg71gGyIbBVV++wvdg57wSWEMh
/BDsWlfjqM4VFcN0IqcQEPIW501ZZrIQdIAv4MMtsX0Q8O9L4M6cTG99vKhiGPFyl1jZpuj/IuVP
Gs7GU+OlAznFwKiZkQN3OWNka4lrzrSzNpQDtsLR6428Yh7G62u1Bo++ufJ4fcR0qMnves+38II+
k6nhtth3ybG/xrUAFDogmvHicC2PI+PbYk5AKrXwL72sPP4Ip0pwrsCVk6r8UomjjQqEul3loDwL
O7qSD/MuaMBw3/ubcL+lOea8lWgWq4wmIKro+3oZBc0adV39E5d/ybl9QSupgqcsw7sCwXMZaFXD
XdcxmJoaxHibLC0llJIpZQDEiQdvE4G8+FTTVm7VyR33bdhOhtxu7d2ZInCbz8k8CE7yDJ+z7JCt
wK+wiBj1GAFBMIyd5c29k/FNDMNedH/I9dtDkfVnYkG3qWU1rNk1GYytdSsh+zWGJlW5xuialen/
qhfIVZ+uCrUAS3YLCPaaNMfWdZB+Rtxe1OaCigXtpHrAv4FKU5cIHie9x9LH9texqE1VWtdkwfJS
Y3lUvGnjPsl+VnV0v4HIhr6WvCeuFFAVEGsAggQjqzktM4+N0GSC5HJTYCnrwDYjZtPXhG0s3g+4
UlQsBttbfiKqaj9AhnhyM/N5wj6bnbsOTDmg6iTe7ogjhxUjdEtY0LYNgu6wWHWmb/Zrr1smRmtn
DucQy0l7SFLS+wXrmeOQ4zKdv/GSYY/V7X6grqRqYhsPJfWXCY36mvOIGQDdqO68VUPeiiSXSYYG
dorR4gH2R+5cWtQpvBtxFzWeVOfBeMQJXtDjUvZCAEr94018/a1TAKgCgBJ7gbsy37OYc20WJd/a
4Xl0YAKWZZ58KMJLlHWSLNYtjgc9DAW9/U0iRw1zKnjux3T14JyWcpOlxjygKlttGJVVZ5qCXv2r
9iHzMF8pRhcsCcmhivqcJlznQCpMU6wMRtc4m99Q91YoFX3CElbxdxMrip3WxTBUFlJwcf9rI/pY
tY4Q6Gsucq6jFG4s+WIQhLKAwrz9BA8Dm+cW7MUjh2mQuVnqFRZ4bI3JiSnFtzGnA6ui8HW4W6HT
GmREMVDgwjkFi8m+PfV59EMsaz1CmV0VM6Wge65scIdjPPOh/qxB3pho0OB2uJ7cFHkwNnjtWeYw
AhRSI9h3Hz6DN7pcJ4sHYTI2CP+0Si5X4NlAW5jDW5L8pdhL2m7UajwR3pp7YLxpX9qCPosrdUrb
i392vYhogQmfK08BfBceQg7r5VcCk17H47GnoRW3p26QeDUfhsd1kB/Sg3glrxUBwwB12MBce9ue
2UeWQtXUlLs1yhF90oIgMyDvypmRweljcR1Z8nr+/ogr1GuvZpr35yD22OH9jx2dOcLDrSJEijcF
4cYNwisFYjdaNWl207C8HbzwKbUDreccfUnLMeLPeuhvm4QnGsIaPLqtWbjAEoSo4k1mnYHi/SXW
wcLZqVh5Q6zE1zIOUJEcyZZyyTr5sG6TMOzgFakORp2xm3EVE7D8EUoh50zOF9eUku0+SAMMS44T
+9HoulD15kZTDecx5vJj1Htjo9q9SpXF0dxaGMfFSNbr0xEj0K2Ph4vdHOsI1yVk7dWU/DMkWJ+S
rYw+JQ1HSqTHotx7I1tF0V2iWHXs3kKtSOCoD/DYy6+22Mo599o1ar8PsmkQeaWWrtQ+QZelDM69
wp4XMT93mfCSlTrQWnankky+4KmqgWKfm8j9j4iZhNgAndZN8ujjsi0wmgmm5yptZnq0tafqEydl
tH5H85R6DSvTwd0czHNkW6E7qE/A+Flgi1odCR3oensn0BK/jJH3mKkPvGDYCQElCj6z3SREA64o
pGy9ENOS332FDLid0tNco3oBZHXhi+KhsXokPfDLALYKVyIrK4zkoBGsJvUdgpq+u4lOKQCH+Yhp
O0hAdFARgW4rPwc9ZxnFN56OrazYXFwzjSI1/mCwhF+vfjq3UQ03XrtPfDltX1/3AyN2z0b+m7cn
0riqrr8Zkqsl3sPogY99bO1WCnU8QRMTrt0g3YWw6Oe4U0ljwuSVUr7KZIHeOW0Z4cxRQj0OR0Jz
aBb0+b429WlPVKSir+VQwyR5ivKpbaYOP37tPFu9uyapwCEsPhmwfNzJ5S2oMd8t7l047plFKv8U
h6tcrIUzKKV3RmJMk0hnYIpicgb8WPzzn4WBNFieoeuJGoIKrI6AitVufrhV9Qqx3QH+hwRZwpqf
hHtW4Jld++21z3HKf20wPAOwk0yZWlTpGw9Q1L8L9/AOvnOkngOa8njcXkGzcxXWjQVrcnuOaTXZ
7AJq/OGmoETPg0vTs0yhSib8ACKebm+Z+30yl4xkfRYq/gal3RPRo0qp/TYsnJurCT4H2Kx0PP/B
eTEq2OmFek7jlJ0R2ljJtzNZ8vSIaUivskl6+uDiUg7t5W6eZxQT3ShvxK77SSAYe9ollP/xR8oo
uKeohkyD6vVw+rus8N61RNNFp0ugr2+Nrv/780/cXOu6ew9wPzowNdrA5XbUqybjoHa34dycABOr
q/7Z1W/64QSYbK5UXD+mx2w9ZyUd2In84vPnB8eCxbzMnl26LX6SInYEoxxwxjz0zWx3iEmI5Umy
WrQQszfbA3mB8ijwcVKQLwtVy6IZdI6/pSYLKY1wAVmcdmIyJu0AgZRz6XmMgLTh81+78bC6WS5g
FyUYDqYSWhmp+JIZODtl049dPCkLjcjsB8LSVTIxnh0oGznAg8B+zSFv842aV90MNJMJSujwsZj9
odrxINQWfKvW0HHa1TYgHYq9to5oVKCBa8oX7K+48+r255uK7K2s54LWgb5KmxpQCw0ilznEX5LL
gDB2g6AksnAk+ZIxTFPQ4ug1R2WDdrEy0xnPZn6K4y+qh09CX4JXZtq58TyTpQpjd+z3uykJGV2I
KR7vXbaAjFLVrs6Rp1tBj4jc+hMibrgbRHBTE6KMby+OTKZZRer9H0D41+5tLqGW+8o0dDPzP88C
2xUmdrm1uvj2kAWX5qu/x+7PJZA0tUfoxVgKzWQ4fYkUMHya2VHpoNLEL8zIHa5b+HHqAfq6Tk+w
YUbL4PlQbqsBWJkQmiwwQTgRaLx7Cuu9g61dv+0tbr3+fBkNfcdgrPUE3+qCiEo+Sqi/XE0r1hL/
nCgBzen4kslFAx13weGNtGPb2iQtvbTLRUz2p6XvbzygYloCPeIKPTuJ90Vkd7LrKJhqOJbeNC9w
ildrnnrrAIhFWl61SB6XlPyaEmIJ55eZ66eWt2yw4iGE4ZNp+N0xl4AgjxUH7BG3soy+I4eZpuvI
Ye+SRPj2t86TFnMmm2th6QqeCJB8Gq0tIkKl+SwARONDCugPIiVSuyrSOHWivacAR3o0b9w/X5CP
/h9ymH6yG7u7/DJoNs0AEM5NHg88VSY+m511HHME+d7a/sCB+WPKEa28HoksL7It/BaTknOGfvbY
yzSG0got6hkSsAgqBXbt5BcwBjOWfMfSEUcJS/vjTGipusNXs5Hc9aBCRwKZYVjEucT/4NKZnNx1
Gb0sDKBev+NirG3CblpiO5xMsQ2RGq8bZ6QUBTpWyszoHYck0e2Z2gEEYY6Hj8NVwH+1+V9VvKK8
jAPet9vUXFLnOAo2l7e9fsLHMzhsdpsN/FPuaTcE87+C5+ok4qWJ/cQxkFL4qXcP15vNigrMsptm
/Ne82W4CpBobvfKpJvL2EzRzbiNcddH3u4/WkbCcXLEUO/Wn2jv4e4X3m7WL7HuSFiWA3Z4naZMx
6CD1wBvan8/N95WU/MdyVooZZImdjzf4BI7vzl9F9sCXHq1A8s7Be2+wc8GmTVs5h4XaPhXrXJ6C
toYBjuXhV/OKuZ/OenXqVlHteExTEy5EHRmbrtiJ86E178ZRu5uzkqgusaFwl6GqNR2nGDILfhSg
FWicqRQ0B7gF9STXfk9VDw9R8UdtM/Yvhsr23W7vBpjjK9oomQ+EHKWQAYl8JJ60NbNKjclZUuyY
/K/V8b+/D9Qtil3JagmBD1yfzMgegKp1zNRuvqKeCr9WGkLdkPGjkP8hKTYIHYicPnukAFzn5Eyd
/swL01cShRPFNBAj7FWA2Pvzh0PKbwpfIq1NxHMsUNpy/9RnRcnhRUJ6PiWHkai6lcQPJP75P/vQ
lg/OphFJyucqnwT9f+sc/K9TbrVXqvW+ManHfMnK+e9XtIyGTiDZ6zq7cQ0DtxDRX7eADYgsXMjU
TyRA7Rvm3i0/ovdXc5Ihb4LZA6u4GiZlj9/zgquFmXOBivnp2k5Ihss2dGVpZxx5//fcN0JBrpO3
ivlTMLzXT6f1l/ldyeK7j+2ZAvZ6BYpcgyXMgduqpL2g6HC/1CobTfPPbVnWoI9/aesEmFWlobSg
RFIaQXH/mj0l71EMuQHYs8lHEn9MbdkCe4zsap5RzaHveflFBBw58YWs9PbM3QYkfSa2Hr72ekBk
IQcS7vLdazoI6PrAsGXx4iW/A2DcetmbdGGufCy2VEQu7bKrab+5KUT5tlihADwHdvdl5RrzU63w
dCNGdd6s80AMLNcBWYqm6FnOOafzwKY41d1gmQRqDR7NQSsqF3ETK9IddIy+cxRlzQvswsgcxsdN
0LW78mULJzLszouwobL2WCU7Cumy2W0fbKeRBwTONxDr7qQfqdmaw/ww1BwzSG++7H3NKcWBksOA
rXiEBvIxOGK+roctx7FZqYNqbTqRW86dVH8yjJByVkO130/Xrp04zRV9k63dW0Qc8ovc2CRxKIvR
wZG8dlfWS5YbMhdBWahS+92hCNv6gjG4zcIHhiQUWSZ16UfgAeBdBJFovASAaToevv+CiZ5sXM4H
akIY+GKivO+66JNUjGjKQIKGBUmYfQvGH70fIurTWklNYXf7CvfMaZWwOURLP+PiBpjtySp8GXMc
IO18JNlfQhnEgGChVH4PdI63qBcRsiRGGb4oxmrxb2+NAPVWsNJ9Skq+xRRzGeGiBt5tazLxS9us
CwICd1JzJtRFuzSsWpByC/Uf6ocPk3Fox7P7Q4FzB1cjR/QPkzPKvyShN79IEQniYbzeSxcqypMY
PEr8ZFtWXPF/CF4ed0uSjp2SAc3GaeykcE6BehavL4yrm/Mucxs8Nyq+7+VTlwc6Ad2ekuvoz501
xzUUmWrP8c5uYCPNptfkPhsNiVEHju+VoLfyex0Ns2QXpFlFyNOkThphWlmEQuuWxvVXeSrodD25
hnOC/RhfUzJSzTmqLGJcFOCS4NjLWK/kBKYRvNIAkPD+3BsigspJ/V0qA9nmMQW8wITim0tg/dMP
Q6ogT+LQt/VbA/3YaxIfVGZ7/AiHLccvvXDUnHC9hVb359NSzITZzfQ7HVxf6a7GcIxBD5hCoXQd
QDmDP2cmU3c0Ke4RfJvzAG2XG/aP4cNOkOJhnXE4NZM7atfM+JCFZK4gmluA0KX7tKdaPRgozxva
L3CVCnKA4TJ+6kCm9fAwRNhrR/fi5pnSj4MoaSpH4nlTKoBtlZVPUGOASG+G1pj5JmNo6Qd1TNyb
ix3VL5k05WVXucQXtTkNf8riLZx7irL3We70ZOmpU5rvdht6ZA6ckPGTSnB6PPg5NIpJ3u/UfBhZ
Kz/Gj6ctrvBEhKkVnEx5oo9DjJWhpJAW91zM4AcYwnyGprlWK1zJUoQ/CuLr06aqkIpz88UycZPa
brB+6ueYzbdys9nffabVqRePT5cWg3biUvPdyid7rktPByd/gqg1KuptDYTEFCJZahFVU8r3dhmV
7IQo9Vqx6OwvGPLZBJ1gHBNf9XYq+SmnQY/DTfG4iFTFHjMQYUKgZLWCAtc8rF4iwzUe7kPEzz0T
5l2qxlRThb0pdBBMqYOqPRiz9ln+auT6taakV2S1I1SqmtlvPGhMRM2RZpYO1RCzO6K6H8F2Tr28
REXX7DsppyFW3Id1YbiRyEJQ6LiMcoLmc0Hx76iiDyGtdAe2TEo1Mhwn83OP2uUuwEXyaOjqCDDe
Tetbmt6VJvSJRIK3kqPv+WVIlrwFPMafUSC0eF1zSiy9C1eQO5b9XvDcw9wPO/oxCEjqT3Ayl78y
1azsJ9V5TJhcROgJ+b42d72ZBaJBCzJCLS04A00AxiFl8Ij2Cav2Z7SLv/3PzIicHltktRl+Q5lQ
1nYTIUuvhbxqfA4LQ1xIMWmbzkKHccukFOvw+3sfW5S8aS4ZGlbosbMiqgSIzt2oK5mdseAAIHDK
w34rFFfwemMk40oQOAKbq7cz1DpFnR4BLJPiMX084+cqRiF0hjXlun+B5JAjTzE44I9lVwBKekfN
h03Dl5I+3E6PXfLiqd3IeZkgXHQKdnPf2TG1lKgKbTvQZsZd32oxesFamP/3UVAFC2IX1rgNQozK
sf1xqTr3v5nbUOE/odecYmArDGz++cQpVwOWE/8YExUQHOXryiM5adZcmx4uORZgEbEiI1wN0uWd
0Yn3AgBWADwW+GaORsjghOZqWzTVRL0BPdgjCCNElesX5VUvxPZfFGEpFw8urGQ83cSHdFrFnGY6
uviY+Pj0xFMyZnDNHa0U0dZx9oApZAp/7TOGPprpbg9nNaRAp28MCUV51mcX/68TYuwfm6xbI27W
UKFHvfj1gSg62eIqvo7TjeikWCltP8QMN1o8VPr6n9qFsrsz2iVUbFKW2LoMSSOsY+cN54H5Vdj6
4p5Sgt5E4Dnt7NmAUXXRMG8XbGyn1kPfxYvgnkMjUilTKZ9dmtkux17AVm0dCSPUD5S3iUc+mlAr
SWWSZ25ZNA4Wd/TM+t4P6ggpITkIlx1ZmzRcYl78xBJCLAnApPjo6pNvlhLPQsqSPslqSHsKAaRU
Gyzcy3rAYXOllp/z4GaJyoRaGc7FVm746nN8rCFKVFOPynlfgy2T4f17C14IDdxOMAVnhj4NbeIl
XLrgjEU00D3GWNXhrifWDkgjU4W9Iii4ygVQN0sgWq3Rl70iDPX4LfyL0cI/8a5sdId0pwN8/k6Z
v4Cuw2dPKSz/vWLeZIwL1m5pYmQYyNKGKKLYtqhYo4kflKtmY3kMd6UbyJyrN9gKYVQ5CIDWypES
gyYhhWw5cJtH9w06g6LTcU/APbMhbAMGfc3rUHsH98TPfwvYaYICM8W5ZUvRMbjU+aHcGGTJYmDu
+bBL7WNnzSW/CV/fh4jUCJHxlcvNY/wF2LVMCi8/3NGjd/8a/oWKsxFOg97YKiY9reSyYIy4WwXD
CFXomTGJPQa+iv41ffxTy9mBgoWeA6hdIZQHm8sUu/Sk93KVNSmNCkKse4JsI6NOsqQawB6L8d2V
3kCPZfll5UedgWYYVOXBSwTykGsrL71aRtet/TZ7OMF1ItfcMdJYpJKjLQlY2JQwFsg2DEdtG1lo
s8fLyVlsWoobrfMLP0op9sH7a41M+/bvTlLrgDwoEA5CBhcvHZB8L4gBpsN9HtCkp1cWIGEJO8sy
A04Abal+j8KvtcrfSw4VAQRRx6uJ1pSxSNAb15lUs2P3HB4bDrG6Do09WR2iqLo1xF82UyDAbtFy
Sn4bvUHcmM3okK9/5Qz1tUb5UIWpQlzgWf12KrtyajrxA1YKecilXfNlkshrkkW2Huzh3uXhyVcJ
DFFGLGNogG7yJGcMrfRJti9/mIs9OmW7a9ewst1VluakDXBLipYuGQtV8MtZU2VRdvwPJPc+OCGk
fUBmY7Fs+1NiVBGncr4gWGvbtvkWMeF+Vleh8yAXiH/tu2afCm9q+WxT877Jl2y6sVWPfhX3xkbO
0ClUyO5WMJN8yEEMz0t4wEMOReaC0IU7WnaY1XggEivhjUSVK8BD/JnnX/tGqTqHQq6AkwUCe3co
zZEhG9k9OK4/hcQEOK9kj+SzNBLOwWLLvDPf72lwP5hy2DkQR8OpZYT9M5sH59rDUVi+Tn/JvHyh
AKBF54XRjJYvWjEod/mRsMtgf7TzJEUbB6xEV+aEo+/0IhZRnfSRIc9FXHfkZcaaXK4Slfq54PEz
MyNPxaUQJqAEklFq05C8qrZEiWy9sWu1UWeQoz/rXU7MRPZA3yrUw5AM2e9EAuH6y8SOI7N6yaat
DwYRPkiJuATG3eg6jHY9QiqRsemiocq6eI6gi3QWXLC4vLT6aygRyDPNJp8kxX42q1a0slEO/tn0
yC3UjTfoWWbbUY7v6EWzE8kgBmJDRZSPo9fORYr2srfyS7R41ylaQbVqfYatEXLoNOtJOuxppESU
w9wZGLMcMnJGwi8QM4kQ0gSLxzakHsLVQrqr/Ko9QdHeQDP9KnhXLYV8aRg5EHXFpc4aUvZMfmqI
fiPki7GdUaSlr7P+u6vZysUnk4gDWFiZBEr0lK4Xz/txehL/5qlZqzcZ1Z3+czfhbHbPp38nkdbe
GPWcmUxIqXq2Dms2ElLkWLCQ5nPUL0kh0xaewfYYUkjT/yu7uwkjfwcIr67XAn7RJYkEooXefR8F
Sz/wymACBra7ftTc1REElc/T7Da8HRUGKTDnkqGqb0ehUon55ZPaEkew9nom0YOTH32abUsevh0r
D0Y/HRHd0utfX8PMzi4ITVjYoe7HlO8FI/wQEQrWYaKZZ0WUHzp3tErJrefiO4dZutSO5qvsDGFS
dqhs2wAZnkHFXW8wE8QBVWoxPV3oeNAC7/Jmfo9LMKWvKfQlPP2YAwmZUG2t6IGJmy5k8HegwBpD
t4hIOPiOTcLjlJhNOyvK3JxsuG1Z1GQcOuudfed2FLbnardkjZddnzPqWg+4rOMwnjFdBR6I1ZVE
Q6W/ZKuFBn50Rh3+hUMEy9CLJ8HARnRAsPfde5ifNLvhbgvCV/ppGCVaE1LsYVQW4H/ZEYYrCXyr
Ltty54FVcFNCYJlnafThEWkDSF0k8gVhX2gEbrFyuEw0sXsHNo+GB1P6ty3ZTDJbQEgvKQ5Es9jU
kaQey3Qw14VNASn2nvjwlekDWQ1yZhpDMgIOWRF0IQkvefwIbgyxqjXhLyNvCO0rEUVqTu8uG6P5
NjsQxH0TTdnEtIAM4rq3ePWGcSQx6A/zvrJ8DznX/2eZ8Deol4aquFowltYdXVHSH8053YQJnx76
8VufQXQWkQWQplXflWMGNo6IPVA8zfIXMGR5oUEkzhMf/Xi16WWMeouZ/05KCi7oQD5TXDbmCYUI
Y2l/6XC/JJ2TyeKcUfun8WtNqE5qmtCVLOvNbEDOMokwrdCFtvdZaqsDRBndE2wPXLoUdYs+gT1F
9yKOHYVdf/lChal+Fav05IlP1hHX2ImzFgFydqVBEOzFDWBCglXBvmrr96j2y/XN3I/B5PWz+u0D
1wEft41Q1QGLHQoNo0fQw11R9hSkUMFFI8VU3MCsCWXWIYNzNNcqfPag/v8JaMd1Loz8a3GWbTVk
1idag8wcRpUcN03LPvXBkDaVIJnE3sGUpi4lgLs9PVRKka1cq3hyJak+qf0Lt0MEsXNtcOTf7yUm
SkOPb+LlSwnpQLCUqrREli7wJqyH9Ctp+ZP6TCKJ2o792RQ1N1WK5SVnTdjEQ27gfju8p55CE3V9
xwKaFIpzhG7xYZ8vEgYH42yMzw1YRE+hVdWb/T4JGlwPebRzTrh7pEbgOg8V/dgJdN/y5leeK/s0
4jgG702ZDU18u1iB/Im7ykdfeRwVnVlQ5r8w9UDTPK4/EADWCUGRn7hlS9fkJ8ee8XUzIIHRU6cM
nup/nt3LzKF+oQymGwiVHY6zPEzlfy6tBNyQwOK82jt/sZ6omPTGo6X8xDDfiUsgXn27CrXkjk9Z
f2fnBQQxq8xANgbXTmuwGDG6wducg2aytZHjwZXXSYp36fs9Tdhp1Me8VZ7XHgjH4qrybnZ5P9Ox
o/2w0XDBYf712quuIgNXzyknsJ3r3MlVXncTbThTriov5NnpYqEY/Xx7V6wI/JgBWpzOANmVswKH
zEUldOw67tmo1xobYn6iL4hY1uDH42ugJjP3/ZWPFnRHfhGaYkSGoj+w2+8sUgHrthd6vBpz+bcP
qOY0dhKQgNTAxwmp+l7/EG/qYpGdeV79MgRxvNO5+KTovKPYB1yHp5oJWP/TOBbOlr14PMlvGX+f
ZmAiZkcVuirbTBvxk6dy4lJIALv83+TkMTdq1RQe/MWpsHzijbLmscNinEI/AcO2AYlAnGFCsqqM
KrUne8vIivCgnjN5FVPVS583s5kd0cTH/H9xrOxZEhJaW4aRTyWNd0nMD7qTcfeCotYrFJNv1faN
QRBl9zQCq+puMMnKw3GgVAW/22VASGmWlkyKsZMa6uWwNreSCidKBDkWq3XxOzBNPzTS1OnOf7v8
/gfJEFqNN2cQCIru3kHihbHz2oPn8EAjDPX7uVRR1p0jYUqB0Y2sDQBwtsO8SpU5HtVyEVinKBxY
hdBaLQ5w2BF9Yrp/daiiwZjK7J9W/g6XLg0fbP9sO0iYmfvn8Epz/oN5YZfkgouJBhZe7BfB9NEL
YhabW8/NEQyQt0mgSpOYYvRuuEGgLJ8Ou0udsu2buEzHjZSyy4x86c0Q/g3vWDKwRL+QqT/sSK+q
7DQo7VUoCR+yVmwQVdNgJ1abuvysWqbKYkagPDh4bytsWrV1GKgTis1y/fuk4HWhe3epPVn7Lvgr
/l2GrqztmTpGKpOOXfZaw852ZYghyUXd9c+n7UONb7Wys6uwPupuvzm6iFgOq/+wnBYyt9RcEF6s
Y67CVK3Ze6A1QZ1+XrOqGu/i9Kj/RdgzpMy7iqJ2I2DCVLnL9zcYZPUHYbH61wJxRdheVaVGZ0yB
yjczlAEz534WGIl4fmZQMGPw8oGsVibtOZQSaAH9G+zkqFVrG4HCkjULRpQjftIYGCSVdaKqNu4S
zWRjpx98QbBeb58yEhL92aY2/jmIkcN0Xzm44lDZN8fwPIWsLYCR2OhxkiRfPtqgMDecxa1psmJJ
uZdhRcTWWUhlZ+Bl+Hd7WTlVglo8X1l2J8k40Wn6KaGxCqAM3y5DPE7wjj21Ng6ZEGNtjxbZE+D3
0ssVzrNVHFGamUWgFSRRC9YjM0Lzu8kRNrrEHlEXvsC53JPw/is37gu5XqIFSje19UYajEl9nbQA
YDUgdoeyrFaaUBMq/zAIkQ7MnhNhmD0W1mflriICrYcxZoZnrxYS7f2WbOuAl0jFWwUnGjKo7j0n
NUAQJzbgVDJHsUtAS5eU2ZFVyY+rU8NZeAZhV/tpN2UJh0U2JVZMVNnF43rugc3/H83aplvWzvgY
cl35wENjdmwqKno/ws5bwoFf1XkOaLJjhgj9Fd+NRpokN9luyJOQ3rxzaOjfw8Gta26vFSDPDANm
qmsVbIxSwXEUFLIzZOCyLx/jJRQ0QLu72SylJCqe7NxZZ6MRo+9yFZfKMvM8NjJf8hrXE/2R5/vQ
4TknQy5MBLOsLEF89nwVhwF07SxRsQynhxHpr/OOqKhZYHxi/TwLuFAqNufZrKLyc0VPFhw6QUxp
r44DcEMHHGU/1fGOM5mpLnlHiKlzwomJeMU8gLKqtMC3d+WK+OAeiofz1gaiIeRgmnJsckS5kr0m
CxdjzydJtkaygq/zUHzwkfFmJ1f48qc0u2kw9ibxKxnPGPNzp/qYGMk7ZwKSt4gk5hpGKmzECmj/
LxlTydphGV0ZUNj3ZLjze/Qu61ISwDwrWJK1EKic78jLgrYHd7VU6Dv85KLAMNPTCufFGMGMwHXb
f2WOxeIcODbF8cx5BSpZq1eT4bfenLMh6d8HtFobIHBwpbEQh6zHLXZnaoa9LLNnrctCXr7BbvRm
tiFrMHQuLAS7MmkBRRjhBCMcMUQhMScZgfyupbE21y8evFXI4HZ2hPWqhmfKPyyiMw3/Z7bAkc72
mQcc/bvhm3Y0n5CgYY0TG5tMRwfdr0Q8G1yLJu85dJx0mkYRm9oOc4cD0qqbTZ+ocRH9/O9wU61J
GqlMo1S01KETUZiSRwodUo+9oI9qGWvqsxpbbVvCvQG2iEDiylBm0X7tJlvsOB9pGmIulqJt/yvY
fAlWvLMiZvXBxZGq+F9R9iEOChy5iwajQFmPGvoMDq2uisGf+yXmQr+0/ADBkLUSr28AoLYy9ZL0
cq/0Q+weVo7LxEWpfY4/hDL5iCLF9eC7nNlXx8hSX28cy8WOIHaPmesxSioAAtigRcMBRKIpjypX
EimKJsPoQyK0T6CVMNz4gGiOR5RfVVC4T864VVPa/INCxq9hFad8wqoknbxWPguXaYTh161M911W
EH9CMmn9DPciMdBdB08pUEtTUKKphyTP8U5I2Zfjym+gOWWo6LhlF1MC3bcUQkzzCV9Q9sPPKB/P
M6JJo7EmHl9q+gFyS0F6do8vbenS3v3xuARsVtVGG4onp3rT7A9SN6UAunv59KuZxIVOEdNXljwR
zE65uU+F1XVZTgAnZn0Z8ogJbosonDOi8mv4fiJoUtAvd1Ub3z4PfwADApLst5LXyUr3QO6bJNea
nZV3Ol6XlSiHyd4wNNKYjIF7UJRtb/bvFR4esg6Dq/jCryMvhMYi4qfqJGWGp9QnXADxwnm38GD5
fcn2RhDPwMhl2oECca1gKTK/sA3eZHI4RPIOgsDfg9PK5V2VDBS7JGDbn+5qQGA+X1waDW5DvaWT
hPgfwwAGVCcAVw53nGxLOoHN3bB75UoYMYj+V3lIHJo8q2Hv8zmrlcwPiVcnEUbxUsrs1SNBjtaz
9wT0C7BZUgpgfrEa4eZ7lLg8Son9iZj3Di+51XtY3WJDCKy6Dqfl54Wlht6qI3k3QHqBwGQ0RKeS
g3GXn5ly8hTznehsodyx9ZU8SAVyDGP7ZrNNX6/9HEjJQhYzDBwQQ4yvMit7FP8qHjvM2MPlCPN1
kLhBbzCtMHIEJQYDb3ujsPm+uiTrotDjj0RLe9uOS08MeBaoP5Ec0EYdCYXUG4DHpN4XhVwMvH6P
ZxRbMT2bTRVGs+PdvIb4KxTgj7guZqkcRDIfXXZo4JWNRWtNCU5iXd8KQaPW/o/Kf27ueMmNHTOk
VN5osfo75Tdc5Ev0t2RggVKaPx3HnJKSXRM22IWpvLzO4P1INXdMXI9Zhg2xbifCUvmLl+zJP/9K
ZAlU2O85EaZLOhcbNOFadOsV2Ux/hAJxC+wFcwvFLTXxWVpmOKFM/slHadFVfQnf4/sMEJCediAU
2EnxWD9e7EufMxdm+aNtnyG471+DSdtFFGT8u6l6SoQ37errTfmPjZ1xv6KLgiloqAMlC70gVQrJ
EPqlousHk867DZROO20pSHkNpolh3HEjU6CRRK6hqGXaKnfxFHfrYRC/zQgSA2y2Xq6sIBBOU/CZ
eZqsxMPVF9U8YgjI7O9UBhvINNrl1xskpLg9xSKB/9xZFpR/5oIcGVZXCN9iM4XNC1lkCvcG+yLq
deLwcpVxjC2QqTS6YFscM4x4/DHDPPg46MVQBpLKhT17+N0UBx8h5ckin+tcCoQBYWmXL3v0cCSw
T4q/C+Ig/wgtAC4XW3O6q83wI38Lzlt7MKSqPxNNtie97YJqMztYTAK0UTpkX+aiCJ7NNA6IpuRI
HlOKcmoyM0DH3HIPGkUbKxjpLOqo0Tz9kKWRIvtXrbJAnogycCvJUT9TXu3+W+638OdCbWZcFODH
o9DxTWLngOf6bOR5OnzVTiHvukYwxKnXDWkFtAjNrg3604cxDuobPH5xKbyMbv9HiiAayWdcNN8K
4Hod7+kxSB1KVvXphBmKAl+cUpIRX6gsGTPb5JyefxsPCSJE6QW1cbVauASKCoxxMfx/SWlhNECe
TPz+VWJT9yzEmPV4bNCTE8vF0cI9PB5P74KkgFWsLwtyTk5Z1Dba1FgfqU+ml1fx1rBaqAhkAPqE
AuN8OXBFhD8xnssS149xFA7wbKKzbg2rJJJgWQPvmOxHzR5oiFXOQRSYIEOZWmZHuKmWfHAXGGMV
0QoSRwyli6gS3WS8rPaKLj2WW2Bg8/+HD8KxlsH4vcjmp2WEY6o83kvWpZmVfVzZrClLpOEUjbzV
2d3nLFqhvAH0mP9a4zYrvxS3i5Jfg1bvzzcVx1gvYwCSacI2zSt411hvi7nyg3P9KDnQSyrZByut
JwFHaS6DJsbw66iNNjAWudGUNuMhf14534/T6rpZ15bfoK6qQH7HaioYMUUpFbfedmOeOF8SpnHn
Kd9Bmk4HogrsHDxtnDuFMi7bwqsMK31iVELL1AyKyB8joR3+JCeWZu0twi7tSsDYSFPbUipJzwwK
vltdBmrt5xbqBW+vA1VLKvnR2oxesRfwb4fes8obaJ5j3td29I+JAIhmJi00nUkCd7f4h9ZeepVg
TfF/2JZ4bUEQdCOFWqhbce1bpNVFVdMA+LDK7EkBtX33hvCPFoASznjY96vdH/p1DaBYOn3X0Z0C
TLRQmURJR5a02yx+VaxEYTlCrnQqky3FRHD7KTHOhGdPNjEK3eXKte9GxzLs7V5ZDJs+BE2DTXZG
/l8QknMCahuGkftYqGHLTUK9GcFzR2TYm8DBvgPVHcqq2KwgA8Lm9z5cfMaqs9P3b+0eAm6NXqqs
SS0VuuklFx/4izy5G5lEBYkcIL8I+JyOb9Tj75IvCzrJYYt11XwjQNbsfu9q/xCbp2UetYnY1FsW
IlU2cd79WT6gN1atgLCvcIwgOaDfI7ZVTPsC5yIh5aP7v3X7g6153gOfoS0lWzx60zm9RopesOvl
JufMavfiLWvr6gfcSWlnU5vKValBEZcGu+cH0e7d3lhhoqtEz5ZFIz0L09LW4S25tO6RgEkk5QAk
GhBrNxnWQIxTc5kZaVBm1E59+C7m/npYMn6aSHMpwPjiXqHjsREaQjEldA9aWqe2p1bGCWDE03O3
+cunC78wfi7s2ru3lalI4tPhUAaxqQpBJ/sLl0MGBdxkgQp8YVmCtqoT6WyhB0eoShqf3kokYfIF
1ThSrfBaTuXK1c+LVJx2nwxKzZr/MNbQ0xiFGOS3Yp12dVV1iTrT0cVVM8doMva/kW3xQTbOaOYH
bFvkHXqHAvp9LlDg1EN78pfu5YTOLrlSp16v9vfopaIYN+UDsztYJ892NJgbG8ZUQaOOfcj3f+R4
q6N7i+Y5Gqw6Jg+HeMwqXmKaq1MXGPvdt2vxItn3P6UggpW0inRyUHs5azs3yCYtFInt/h4PplTr
YiQg8q9UVg6EfSXILXkEpNXW3AmxScLExhxK7TTQnnG0Do1KwzN/TQKPYcKar69+QAQC+loiNOb4
Tbg+/CGDhPEYUGJ1uNK7n01M6jM9oD30rt2e1IgMkrS+EdrXelPoKTl51lAQqbcdUUKQ1PSn9YVg
R+HYZYQENrvQ8JOcC4TGt1NpDFQiO8e53wVyofEZM/oi+35vDpcKildLGTNc5TQER75xIgQ6mUbV
pE/Guff207WeY5RVOiMwiNShdJ3tcYTW4lppkFZqRRtZa3zt7gJMjr3540vXFx7ujpnYMK3ZwB8W
c0XlA6P+CtTyuSFlTgOp6XervtnLvXLIVtSCLQvcqX/uR58sH3xRXj0rnozZWI8LbHwWAshgk0+B
rO3BrRdAaxhLXT5iwDS/3ePtU7SPRjtEgQEue0xIEXSMZ1Q57cSkUv2y+YePKuLfdZ4Ul/jHJrQ7
+aGCxICpo6097T3vxKB/Bn8uZsUPf+uBhV+d3NCrw7BzYrbrB4XuXwMiJpe7/QB9TTfEx9vPlIqL
NzGuAfGXAcjgjDf4Ac4YXV9OD9MXXgoaK6OXfytZUvc+BhCAPofEtqyLLvZzWYJVw5bfa2gkjAZh
Y20mBz/q+4Q7U7fXhYc2Q7um74mTbmSR2f8KRvzyBv3M4LzcPpUmhKL8LMp7IXElu/rmZ8DuGz3Y
5JXxMj7m67k3Gvb8jNVGraC4maci/E5pDHg9T1byUpHCv7TncCCZ7f5rDl4gRjqGsmbmR2vdNGhP
JEb79/iQNCK8EUiO8W+FpSjxuAryxbIBDdUB0jHamPGhyAo0nkyuCI/ltlDGaoY9zKTKkaWp3Jc7
7EOgchMNcDYMf+qlhp1A5S1o4Ng1NokJzbts952djuG/MZVUOGAxllJqVpeSonn7DSJ9EYv5p6pn
MGhlwW5bxIWtci9vFIhUo1yuZtMPoM8jJuTBe6SWvc7JqCa9nEDrkY+4Roq5YcXU2kz0NPSCggrw
RUORVmkJV9NEr7uPQsO04XUWFpTKVI+XicnGxXkJRRvYoEbzTEpTR4XdyWV60V5atd8GLP98LVLD
uOnlwlbpZnPA6dDV90t+biXD2Hvb2vMKepmCw3tj+BDW5d4bB81cgGdobyCZ3lvKpQqoT4/8NN6Z
0Cs0zWNW2I/vkTsgwYwPmcOLEU3TpFQSGf1f4609/4lnbxBHn/859yuPl0tg2wep7qFDQYZAqlcu
hyFS6An9QGI3lAn5x/hGXuJNqIynOgo0knft42reOUo8kt7yYIOfVj/NwwVGYkrQFgTmz/nWc/dP
YN9dDAkj4lL/WzynbvKsPxjpeZIei7e+guKQzNirnkmWblZBWHRisMkxhbFvpkaqOBhMwAWpdNLs
/nH8IP8eTQ+ed3paBliCEmaGhltcr6OJEkQ0uC5mFTCzQ5AmFUR/sUPJ9rKISx/FvGA66zkrdvn0
Do5abKXZh6JHJeYu1JogVxMK/GPdZ2g/TxLsaARpAhpcUx8ErQewT18xPv4/ABnM4K3ApSbLP7yE
On8iJJrNKvgwNzUn7UKXt7FMrrMEJdQ9yr62g5pTuB47KQzYkhSzT0OPs2BD58/Ik0WTDHOOLKkf
QBxBS5IK2Jg7o4sk9V5XbHSJZVQZCI7DVMbJrbA4/0tsYEK+MVxq2l4uEr++bDion6HmPmKHlyog
/cEZsy/iO2kjsfDcCt5f4lXdMX1jWZxCosofqCqhDWagHkMi1MaSA7ewVHqUUE5RVEI/lB1jvMvE
v0A8RA6UPZOqBbtxaj7WnSqmqTqj8yHY4Jth1YTJ4RLnHEKv2E9x1higzVam9DNuG2Kz6kx6fdve
yOeydoX7UrdFzSngltIjKzxuBfWOXOBeoMFcAu0QldNF68n5CdyZBb4DbaDCr0Q9XuPaxTuxJeG1
F4pRNBWO7q20zgyBoG4bvsxr2indH91jHgtytRINqoN6c+7tw/ZZVrkAJBC07UQnltIagDnXCDuf
M1+hZaG0fdF2jeLSNnjAPcTE9uBSlpHsO23hx+vgIEaYAdw6nBCxjVbIZflpgVKaxmKhuawB9Y9F
UrEJ20XqLtEQ8BzWHxo6oKUfUy0sB8G3bMTeUNSfeFLrMNyKYB4d0RyXTzB4IGtyjbC+KyR9n3xC
JA/z3cmEQY3UQ7hpy7xNtM1h74yTYiA05zUfLu6Moi6UsQirc40ckfI/vHf8TQhiWe25OmvOyjmv
NJlKAXZiicGmBs9r9+6tQQ2HJ6uUjCJszh2LTzHodIlaRYrLSBotkHcL9tOCcWx9QS84xnnjFg12
uE2DkVwePbs5koZUfUqePhct+Utiulj0PGHA4UtyYJVhQkhBf9gHbJqyqlXalxVEiPIu5on49Gm7
FgzvXQvazHj2XVboFJpe11CHUMcmogA0zFJJMaUvQN7qk+34l/yb5Uhp3PtrJ+ST2J1cK+AkIr7p
j1tsJYNJy5j5dOqIMfI3yUBsOkWQj5k0DBvVqmua6h+oTHHilfiBdjUlxtrArtZmCE59HDnUZVt9
DD3wa29VHE8XMIUGe9Ge/Mn71cuazYY1YII649wNMW8+u0Oni5GzE9XtT3zROjVY1I2L9lu/2b6L
9pM0FUQuWVKH/OAzPkyqNpieMlw5wRSWEuKiX78l1DfJP9+paJpiOzOVL4YX84BLyNtB0i4UtLlh
Fql2KytUk9L1RNsJjmvr1UScHRU8j44tMXJB6ZfiAxTj0wyrsM9C4/UM4jFN/9ZYIO659GVJsDig
OElO99fmDwWnWNl71WIKwhr4pvvtGd07+dzjkg4R3TlnBHCAjpQ6jRUOkw3HdJ1Gyl66r8Pgea5J
XCayuKeEitDoDDiJzWXqUT6r4CRkQ69usq6oxJ448zPgSM5hoHoBQUZ7RBMTUGMMbm6KtCGeg765
dycOZrfIOoqGcIRTdbFJY+pDbEF8JKdNIItSe/N7A9fzEHahvUDN6TOzJKyUyejD7FSfta29e8K9
KtCYsHuZEpZsDV1XKJr6/X//Xu35Yp6DklYiBede2dXj5iUyD+NJmQ8wJsUmEffMlLRTwbJUPNE6
upMz/RHrrzB5yZQ8YRo0MfBCNvgmIVo9Kw+P2Gh98Uw8UejYnVulqMl5VH1YU0bWb32Wwk+MR4h7
aNOxXwHwu69bLT89zNy7wlTv++Jrb76Y23d6NRavAHXNAhuuf5ybfNH+DohbsJdlG48JbDrzm4rQ
gCphCK0/0sh15JiBy8PgExAEVPP5LQr5osWCYtyyTXoYvxpqX/iEMQz1FNtrRf1gi2zcP3pzA2ls
9Ll1i47bl3USQinbVP2/OzK0cqBkZ3UKjcL8tUoDdmk0ZYjyr+EqCVM8oO8B1nGedojpu6xmF6F3
4bvXDhd+4NcfGQDvH4Fqmv9hiIBIbH0Hc75trPuC0ikSUmGylgl52uMNCaeMmW1VYtaH6D+kU6fC
99mNMiJd8AY++gA30jWoXfgznWhYsJbCUx4rrXB+JxkyEY5su+9wQW0zkWP76M+sa+vM8TivY/ho
PsFr6nuybrTsGR3e8eRODQlpi48EE1z06TAqIGlrhE485ugaXYlAkM5ngTsVASareE/1ciqBqFL9
lpRaTzrJIBfHDFjFgOXEbkCDbxETqcryZQiSD035AM+2AH1w8Udm6FPwtVvqEnhzdQ5/MVIQ85Ly
0ikRrcW8sqXKLR1UVYEMTwW/Tq8a5xSGcn3/AQK4KLMWD6FkJNweAasp5ecWBRe5gxSsHCn42K9F
AxfNghhXjmFWLTvp4/sQYXoPELDM4lHXq779ldgDppgi2B7fFk/Jr93NwzsAjbEWuD96RmEGj2sy
ddbeX4NSzHIiw1LRwIJvT/ZpxfsbcjSOokhqnrbselmE+Y0QFD1OQ9yvq/brLJRJzWGjP8U5dWRH
GuHBcLJnKLaP0zYJAd8UGnV+EiSTcluIaA8DBlJFAw6MOPdIzXabZYkZjNouRDeMvehtOCBocbMY
KhovPDC8Dh+pkUaWBj2v+EvMNKeBMjO40S3cHstXuxLfxgPct0fpx6dX9ayMiRIMLDiyYXOYBuaB
qTaLdVaBk55cr5gY5HwYHVkzsbqhEaCLP/NB5kUsADrH/VfnuWSuSbdmMKIPoFq+IFiWfF24x260
X39+YdTZ8cMCsniBifqBbHXOF6MiGwZCU2vaMDYrDyXKjpQVC5WAxVKU8ieIbpmx3R0d7LfFB3Wt
r0p7mZrhfTEQRA/464lC2RsT120u3rMehDRDtbHpzhp+kOSryNAQtVMc3eVuZHYhdE3qGnt3xxZf
bjMesJX6LdsfH6nw6x8APDJr3KLMXOsUwvxJ0OHni52hBjH1aKYuxmHoLe/2Ki7SVx0GTjMFrVpU
UEISTRDCYkMALbtRmWrJqDMCJvrrvlx1WaDAMogpzybrrphXgEH8y5tgtCYmSCTJvHJQ3ZMg5Moq
3mJPZsxSDek++X3AtpmHU/zHlOkCQ9iERtGkA3liYGyj/ogRCNgCGZR12zwoi4Kk7ajEDZxpCxTH
QbHBOm6zMWwuW1NCC5yB4tqF578Sa1BlQBqY4ftuDUAYHG6G619GztLIybxHHE85tkTTF0RGpBRU
33Jq7gwyuzNDCZrCHJyn0JSzZNDbV0AbleapfwFWJxaobHvLmdGNAt0l8udetliW8xaQaV7xMjkm
5/3zrNCnIWUij7WcVb8r0KZjK9plat4xBBiQEgBmacdB4FVHQdFlCtjOwcukkLCbZpL5tZZi5pnm
BQOVLG/nT1vI2lJcunKj0GW2+NWldWn9ccLwJSaat86IdPampG0rdUfW3RDne+2tfL2lFZaZ38HD
PLF7GeCOSKscUUgZP/xquJBLDyN+U3KZJ4UzyfiC6/D+EcZ49ARwKEbbWVVWnDl9shgBSoyZe9DK
sSZDcm51M+b0XozvkMZKTj30doN7sF0vFgx6EydT/0cQOm356aXbn/kf8jhA9ajlVDaJT+PxroJt
2wU1agYpYzeHzMbHXuuxM1mFvXDjk6IV9fBIIrljGqnSNKiYug991xZZP3CFZPv7mPQuTwqSeuvs
O+9agV2+z8PwjoLPTkyl53AWx5AkRZ4/aT54kRFRD2OE1DtOt5UcmFhDA6hFVTSQYNhfB3Ynjag0
68EN4sweGqTGEDIaSrPHmuNz7X0NGFAqp9CYZjk6CAZwTmtmWkXyUs5s9oISFCulHVyDsAKo/RhR
+x5OuDA4O1YVHyRxIZuWQoX5C0A1PNYUx0v041MO0uqIBpBLVtryDfA2rVCK+NnI3hJJ1dT00GvH
MIXdvgQHTYHagfbEEnhw5ytXC5HSp65wwYIcHFKZWyPfPwonfTxTlcyXjFAT/6VONiuJIwMnx6+v
tW/+41XUGE0OWvG8jlqgAgPU7m5sJpduYHHWiz+mEtYq15AyxI3tSmE03e5SzUCAcDuPo5m3baVG
2/0JkBVd0YIQoziMFOUp9wbTp/geJo3ssCERZn0y7maB14la6jluEZRN3iQnaQVjvrVZ5cJ5eAp6
tzzlLj0jiYaRYmvN4aAel6Wox/0ZD40ZWVnEGkltgwSgCMfk47uBadGd8di0zc0S6Z/DX7uupgzR
23MFrTkwY79+8Qlfi8dtmqZ9xLrYo8bQHvfUIwcfjqEA+9B0dZiU98xRQDsa7P/ih7b98rN0lhO2
VBeTIXqEcNp+cn2iXKrQNxziwEyETKicix5jneuKA9gvS4n8ABp2gew/rMlXfFbY+pddRdHJgzPx
9GoX95qVe5fAcXIUglrJjx8x77JphmmMHGUEgr5st4dPgWaSCEXftFfmKwDkrgwNeqXsm9PMjHxW
R/6iP11kjISMOr5hsJa438NqIJPFSO/FdNa4MmG0NiCnAN8YTtaUCqOBfZA3v0XdcQVLexieHV5a
VCfCgQfLdgexac7Sae20ODPukagZs0SC94/p+lYAXWMJpzVpr6D+ocjj4wTi7Ny0FL0ppla0O9E+
gskgDN0RQKzpS+gL6RVJuzt1M2f/iAtAD0kwJzRk/GI4re6/z1ASpj6tidsg1aq9HMllZi9SMnEd
rk2+EES13/TrjFH5GmYsL9ew6bFJ6swBp61KJd/J6amhMM7oR2IRjHj+TDb/8a6WWVdZGotlXgga
3B/srfULqUa26if6WCvMctUdS2dWmeBh0LII8SU+08TKwi9R9GON9T6B2zGJ5IgPHl3gITtvKSTE
3tMUtTt2aGmndsSrgyX16VTg6ymWG6XDZ0VFPWwUR7jdYIq89a/s2e4RAycQd67HkupPOEDpv5UA
n76NkaKhoccoawlyGyXvVF99mjiRAvqDakbnf1Db2YWXOPK+EKsWva5p/J/Q4BDNJOXEyaFZvmZt
NYiQ8fw4UUhtJDaUqrKch5cWFMn4pn2T78cHYqbhcY9MXKkuLfqBtvcQhXVTH5WW0WCvN+E6sT0R
Y6Q9a7H4UBZ58uZ1kfQ8iVwTSVI/ifqTTkcsoyD/bmTmUQFFLnbXtmZ/RAcoN3CWY2SGZLAiSVXj
BpUMJQts2tNNo978ZeDFaAAQBLEVP0OQZof+9uxwYYenGzBSzb3iIJVXi/2DlEfzeTVL0Lxs2Cab
A61x32rmJTY7WkdgaFHzEEnVuJcgj2QUSwhuNV4TeyfPC/yKkbsMmezVd3SCxEVT0pYBAPOs60fb
RiAScWRBnhM+C7dMBhc7BoPn27hqCQA9dJFmLlrOa5h0f5OPOdugCsXmn26PJxDpV6J2hfynpJjE
A/lqXSpDVUcI5zlfwtW7wjAC7ha9cjhFQ/w3JKW58XLomtsOHewHQiE4RH7pZVlOh1WoXbHUBOWl
av7puftHLy+UMivRV5VHVRGU3cNYue2MPMYy3f8L2tJeaCsIDQCDwSV6ERouy0tCd187iytgegGM
8STSOwh4byj5nKltjKthR66+4Of5KOt7yFm9ubO/qP9iaR4nBteKRKXtXr3O4xgOKI0UtFBBUqJl
uh1qK2veKmLyF4JYv3wk2pmx2V/YpoqBWHBf1zKShtABuoXzkUrKnMETYbP1PsW9pA5SFnQjfrFd
yxU6BKMFFk1LPPU9amE0Dh3XMmWmZQE7zadK07A8oi8P5SbCVX7Okz2TGuuESzWJi8oo4fOD3Or0
DqntG83jO7jHT5z7GUZ5lZmWYhc8QkgZI4xQWl8RrSahtIqQsyVaYCsxLhD6ifxckdXlBN6Vh95T
+Wj6xBB83GnA0OpoqkP2HQ28880KQwOF3ZuMFQaz+nJg/en7CrPQ0LdGKH3iatBMwpKWOzs5rp2j
lO5rPql0hybRHfnLDEr4XQ2mU41FWyV1sDqCzHc4NQFd5gNDt344lTL/xoFsqevUmY2o46hsl9oe
s5vrhOWaWMUxzu6eBjWhN/VIUumJLkkEJZISnqQW6CWynMtRguY2+PjK/ySd9svCzk2o5uL2lFVU
QCdyprQuk04hAB8OW5fINRy0YrX3RkQ+TNu7MGJAg3dLqhRJrEfmqTv6UXUk2oAkqcDA/g1yYBE9
NiMONpYY0ONxUtLmuUCxNxn7qCBbDiXrosgy8n+DxVdS8udk0ViyKjojPwyeaHO8BzGk3j/WkZdS
MdPlbOrrGZcRrriWS/HrAM6LAbp6mRnVt3ipdBupJe4uRmnBxRN85ZnRmzJO7FbWXQrB+6LiXR7T
RQQEEwXHi7qdfEhcZhiQei6pK4zhr5NTFxHmVSCxtycWpoMYfUzjv6TfC8dfp+D5uw3tTGb4BKaM
19BSk4AmN6x4kKbRE2uuVGEMjLIiQJu/HqFD+As/5nLG18Nm3o72J8z1QpjwsaLhrE0P2bZhiPwm
rFopwMFXPgSsOqJugW/piQD6TLYakI/9SzVD8+bp2lerqXrXJ62FsFtWPucrYBeYnYbQwCWxxiCf
M0oMKa5GuNdqlqMkQaSUhNXMaIAH4+EVC+C95BiFIO+7zkp5Zdr+hhcSQkzGCl6dRv25KP2dBB+U
XpruCul7wW8tyTkd2GtjFikInlckA+xj/hSYwEg543xXXwGhu8/WbmsyOdUuBdxXFPM6AM6JmHcD
4f6fmziSup6XRlgFGQ8Uo8FLYXknClcaWej4CFu/yi10eGqyg+fBp+nXqDupCQCjyTPBN2ZtOQcF
MiPLNciyCjQromtGJ026D8oeKBoAsraTUe8M3bEYEWqZyMdaNm1EmT1DjLwzd6IAMJmO1FneVP89
MBqsgegwW0yWJGstkuhI8/u/q37vXbJaCBdYvmyJf2E3UruKovDlmLPp1jLLZ8hlAX84z2/YSbLA
mtt6C0y+RW23/gMJ4LJ2Uks5bWorBGhVvD6VOIgXEbBR0M2rcYekZUmg/Qj8xKw+1KtU7ftHGkx9
filhHjIgf2++zrAt/flUuFLdEEckzQf7m28oS6poUYdIq8AcFhsjpzZn8Xn3VhBHol+f8HUhNT4p
QmUKolIK9uyWso+whZwLUkrW2gpNeK3nRFe3e6dK5jyf5a25pVM8hS9puaAes9PADH5iDP77WT8q
0FG+M4cI9CIMXrVs65F695y2DdE+lzpzyGCsmyfKVK8khjiy3P65VnPz93ufsyJpK8pyqRs1GKzN
1/2S7DdTtuTtgH1prRKYFI/cU6oEZhl/HOVI//QoI+Fk55wmRCdYgw5ZtmZOPjiEcFdS1F4JHCek
8KgaJ8Ds29+71mPMxujsaGLlF2tiWUfwS0LOvdo1w8eKBF1t8GXXAxY685yEgbsTvf5MeIF7c1wl
AKDRRqk0WaR7zzfUgBhDgg2axzW2ojhZ+eqwdKCLE0g/uvwNE0oyq23cEQzPjECSfvXjgJATacQZ
atXOEJuavESsA1HsQYXIRv0jwkAedCeTuT8K/ieRBdLz8ss8+iV97AErE41W/24oroZPsk7PqEI7
1M3M9idPX2uI/1CkwHkkr+zaHc43qe/v4d8OWjufgKpOWC5/4R+WQdC5quHz2cCUMNfpQR5AHq/y
IOycL4/Ods5d31DO9v/FaPb5MyLQMD+E77qZbgJ7ONG4sNxzuvHPW95wrCbXMLdaBXY/A6ApluqQ
SCPv4/ybTbpLocwL71yr8nsxQ+q7N7/w0hmQzmfuhaNuj4iAkJ8q8JxOS5ldcb5plBJyuDimjt2n
22Q1asxGrV+Cs0HfGlDWcGORR//ZJOhKG7CV8ZkyIAOE3GzX0UN8Kdkpqjwwk0GnQX4d4RpmYa3F
gJAZbt8MX/c5lj02LfT66qA5lRH4X/FBKTDiYQI29wmsqaPbB9LsZ8DfTF3W14ubZt6Le5793RWv
gl2YfZDBv9SkYyZ4RXZGQ6KJc9QazW0c1dCemrUSEZsDiF2QBJ9w1wEUWk+ID9FCFgj6kDBy7V+R
RTLuKnUffaPM/6/4y5Edq+4zer68rmC7vi0kTFs+MUFeDBibcRMGLPnEa/2FIMlroBysw459Al3L
c3pQF5ygpCBBRwMVDxahedHn0d8/6IWUHereYHFSK38FRtbuiBIGcetM9X5/8VFUPv86v+bxzaOG
PCvxrXXp3Tp4Kimnv+6Ehiqcozms6jnvVq0fo5hqPC+ES1DRO3pPxQfNMHrdWrao7I+aFgZkRYq0
SJLBI/RD8pTheVzvBPIFmhP8u+NR+bG+Ez2Om7LL8yYh2zdcNh1UhF5JzZJ6H2bFeYHFJVrT4Y64
QqP+x9K6zBx0BV7Pw++N8l3cio9kgIeXl6LoMPTfMf39AarLtbSbnS3s2OMeVCEsi16P0eU8v3wH
fFruVEQKH6vIX0KxoAkR53q7gUENeNKN+k2zJlbgCOCKk6o87hnC9fJct+P+k4nl2MENRnHLleU+
lZUv0U/BNqUODt26kqCkZN8zzUuAvXdeKe5fLG3VIqQVxc9nBHgNrbwOQ1Lw/OfInjPsopYCPYkE
0bMdX3dghE6T+h4f0na8rsLcUEaLYw4oSly4pJouNWaSPedEyi95vKDh0Rf2N0gx3bexBL7+DGku
46Vc8WAND2JTKVBVysZuf4ISRHIcRubxcE7SzPJckRvGHwyvZqjFK/SsvQtgZTKadDJ+loTR0muY
QTuSU8oD3dt7bH7+28z4gAZ6uGwwwnifGR5x437nT/DJdsHoKy/Q2cjRSETSNp0IWwuJiS7vAEhk
MshRi7kevbnT+gX00RqJNjsR6EOKFu81v1/Mjhv75uf2SqqkKktWJdRP6ObqWPpdY+PV7P7Y1W6O
wvvqufXVbzqxgCm6IiNtV6YVlSDdnblkgQY6DkPwutiAH0IHrDBVKag0QiYZC+xNbtNsTTgwqvHQ
m/dRG2Txr6jd/uedNBHFaKhW36Q9JjIONzUYMK/DH+BZc7nrVeABm092bD95GREMGMRxaEha1z9m
qyZqrDwQ1WZ52cxCzmWb4EQjRPlEk/V9BLe+e+SIFwt6xxKaEyRPXvzloZEbnJMcF213GdkaAu/Z
i3W34D8Y6KKLkR5Dn2M8Ry5kJX4GoH8zcMbKH8iki4zm+acGpxoM/0KB4vm9Y1AeobJY/DOc/uMy
VJBBIYpkjDMhqo5nS/6zTYkdqLYkeksE7PNaGDEshkFEp27ylktOiSqUWu/LLaOIt6elh/SqEhzN
PZC/KNaygMGIjNYfxkNc9vKXlAQBXZZdKoHvcv4j3hfK4jyKALA7vkElmeJnk+P31IjWsZhJsgJx
OkhcNvbcuDr2zMCVNJTwGb8QZDdMDQX9NII500zRSdIqlNpr/Mv4gO0I+6HVrqlVD4uoL+bD0DAf
NeBUDjj1tGXxbBb3zCtaxk3UVDvP3hHT2PmrB0TN6euanzGIbRWX9blGVscve0mgq/HdSgWLzlEp
n0jgD1kv6+5fN0m6BfbLwVifQQth7itp2lnOd3dIB9d0lRv6rVYGBoNnCmYnInwuKza//DoXczIM
teT8PfT0ahzDjh1mqKHe0nGm6ECVGHX/HA8hdpUs06gJ1qq1TeLmjBwofP2+aiaxkifsrGhB6sxo
AG5RQwYy4c/yYyr7t4C48WLdwqp/SYN5X2V+zgjMl59CdiWoAHJGPPDA+kxP19i/XeqnP1ilkuo2
js5AG9icC4Wm17/6i9W4T4RhfSo8v34FkiltlwhwsbTzLhXv9CevlfKnx6oEyKH7RGHHFH2cB9G+
XtMEK3BXUC83ZTRUsKM9Uik1TIJeyY1ceJvf+Efrl8XX/cJYqRWNB3UGx/fpbrBV1tkAh3np1kja
6s1M8FMdrQYn8GihanQ4YaX9DklfkoXYW9+IMHO4t+EA4uFLWU5QwngxrOmZsgJbYmYxOZUQGvTd
h3e5Bl9lReTj30TvEI1MgAH/QdFrGW3UM/oTDZIPxErNiW2TJL7hUibx3ZsUGVBTbIQsf13ZmvFH
4leU5SEU6JPeebciHLeMLN1yWIkixwPJmigMHhZPCT26o1wf13eKN9fTWIQLe1GhKG+QVa+nMHNy
HWYjGE/1CLPYWTIKWvDv6Cs5TPYeaH1kZB5u+SRafl6Dwk4vh/TC3hNt4ZoddZVm9FtBwqYi+nKC
N//mJ4b+ixpln++JoDEe4v+ZPhZcvHQ+EDj5YhuuYpUPqMf1K/WASE/Bwf7m3YYBpZ9Uu49DOn8I
OMPQmJ9dVvxLLmjaAPOLS3/vkX/OA+yxZY7BQ0Y6GQij8Aa3I/7JfNxThoO5UHvrMYW44BZlf/bM
rj5Mwd2aV55KREGli6fb4cIG+o0ewKCQX1ZpXU140uWRbWnJBRbtQ+L9640iBdwambgXxlRraSEW
uDWdAX8+dAO8mFyVJawSzhPJcIZmfFfwXkrKjWOlb9li3hNpa9+G9MCt0XPJbGp4eY8wrRTmAvRI
KbAjGhFWH6gq+WqABwzacsD3U0fgVkhBd3g8FbLQVR89hip19iqfddI6oFe31uCmqDe0LYI9oLJA
GrucB+OPhdPjUzTUb4DQ5I6E/rsE6au9InUdeKD4mVf/s+Q9pvytIDsdiz+0uEzqMLV+0FS6h6ie
HAlFp5BQw7/3moxogLlte9TIdvTcgNEYyv5C43fKIxwatcsi/EjOh9AMqhcUDJAk0vh3ze3gPpWD
cuR5TJ3mrVo8LO4xZyEPourItROuCq0s6QHa9VzXWxTWHesOMLvy+s8EI5/CnSL8TjPyk/0PiziD
yly8Q+ynqHwCMmQAlHxAEUHZ/EGirDAI6lO672N3WdGPZjv+Z81rHwy2zZhXtyjgf90vSJEG9kxi
EkX7cnWJy7GRWqTHeub/66J1PVU0ZP5wOvAmtJ+PUIM3/+WnZl1WXKngWx2vBApZo3+vaAGktaly
z4s4dDohwqzqZtzW5nlJuji0R5XhsbVeSDFO7+fJ4tFeg5Gc9AdQA3slW3ObQN3s6Xu3f6WCFzPT
Mpbwyw+sHvKmZd+5jnnEKKQpycVcTJt20qj5s0UlJ9B3ZRPMXmPns+ksRQQLJgyzYF6qDU3yJgI/
25HIbvtTiOLtDVsxtSTRrbe9Ucuiww3HBRhwpcolZP9Xbg3YxXZryyMexhVXCmSzchO1DBV/Tmz+
NJmdpWlYpVEX+SJEORvAOnZBEcVqrp3dr8/D2eTF8w1ivCeMUb9WewzcftjJ2hUB7HcflP4M6xTv
+L8pL18KFiX1esozuWplFBnVjg15liq7VLetDyrwiuemmPvHW0E2d4ncF3z4yZEWAYBdveTE2I2y
8malP4eYoE94umYPkHCjPIMBXbPa7RkylnR3eAAkCtrXthzf9tBzSJudAZT0q3MVyRFToLFfWwnk
e/7B9P1J/rwGxtuxTZpJBJAyPBkND6EubO7NJw0Zh0akoUXcvyBIyTZaCPBqBSPjKTllJQNsZMNH
5r6IiF9pWwESLRQAEhns2ec/mpLQEG4TP2dRrDVEAZcWlzJ16ZkcU6CUsuus5ubExyhMxS9LW4Vp
zsUIaGceBPjHAbrWC5WxxUNUhmw8sIivbVEV4sMI4X/PXm4Rr8YmDdcwT6/YevwcDe9BRa2eGa2F
kvecplhvfjR62zNKiqSBcT2Kb4sOFgMG3nkg9HXUzCbt6DetEihytx5nPB0ZgvItwbeQITivmFFj
icmeA6b/39J2YBU1iRVqCrAo2B58v1nSw8M3vks6rA1XmzXCtvpRLknDehAHXm69uRtxMHSA8Yi+
G/QyW6TaucyYVum6Ewis/r0M9nfXc9FgkPftLJpe7lmu2sjpQGnbu53tcYDhV1ru8WXykns/pyqU
+T2ZewIy1VT3pVp6T0WuMVdTBjF8GPI6lEs5Nirg1KkZeVvrj0EtGoPS/v6VmBxg35+KnHA8sLmK
WcBXxGfVDzOlj5x2n1geUFGPXjWWl/1miccN/Z+YKt8sXOahysJztHhJbZXx3uJJPEDmdvduFC9y
5ix+wJ6axXiq+hM00COtZbKvZFhJrnwwpMLm2Ec0FFwiUGvs7+nQ9ssI2SC7pSupX8yKIy6Rveuw
Bd8VFQAQuyczoLRUMsIdotXTCF2nqSSrMxZFqkyCHxyxsL4gWTg55Xc3qDuk4S648va+WuuubOS1
INhngFwo0WK+7pmbhRWNjzMArkHaJB2WCXEteD2jE+00NXwiXHJy7u9L/wVfAUisdlCJWtYV4BLf
hHGmX74AUqW1YFWDXem6B06JZ8wGTdZ0fOg+BcFD43SMIKKRDRL9YPbP+RG9fzSGHeuLa+FM279b
jFXKOavkAR7vQDKPwEbheDuZXODj4kIzrRwaNR/5QtwM8L40k/BOq+PHNC2sGE5WY0itXYiWDL5i
8x61050UDgSk2rOb+5KL0lSGO5thUGS7jca4cxduMgqEiUwLpRHgFFVzoQEFfZesIAcg6MzgArPk
MueCxMQlaf1kRd9WsYzr/fmvskAKFZa5awyksNSF/Vx8ltPib3eIVX2zXtB191fWkUYH/i32zQqr
uXu1Cb5etWRg9FwhwgP02uayACqPlXT/lGKU/MM6VjoFQKO4KMQ8wyP1KidtJtiZOHUAXtJE/H42
ETSdGyTIl+kjRGC+BHxuSlOq0IKvCCKMzJByqrmPrzXoTCwHYqnCmarMZjc4uvS3Yb8Lv693F29D
UBm0IQXTdoNkULFDsQR4XsWHepL2mApiteRNenInXl1jsKrD9fdvT4OaDoJ+tipkpsqucTXH3Hq5
+2aKyG8iLElnxNsle9RszbNNG93/SV3zbqP9dZRZy+JHgeGiu3H0uO6bUnUVppLCSyJlG7kqiFXF
v0QLD4NlL73PXXYN3bCdIoPPvkLtEIrUCH1CwQL3+wzseIWVV9ptagafxNlW321SON9H00rq6EV3
J4MHPCFIvwkb+EoG4TOYORri3yDrFOxJWuOoAWWXMWvsOdtwAHXOmhuSWWRZmMp+Zaoow3P1zpgp
RogHjZ3yoaAQ+ITAqJ20ofjYMYBEktVYR8t37+31kxM9Xq3GIAs9CWOY9vG5EkNrFftzKrgbTrXj
d98VV8euCROjvwsfKhMZWOaiCKVcon5vQmzEA/en+FSxyTk3ENQxQ8DsInJRyR0w9I2hetLctwRg
d+dRS/ybguVZ2ZFrCiQMGOkoP4iein+7BFSOL7tZzx0X5IzgMkVshSwGDR15uElwDj9ZMwMrNuQ5
I3MbZdINq3fqIl/dSENATHcVzIT65XCBtLF6pslZlVvMjVqJXB2JTpi5XXgg3dbKkKK0BdNNbqp4
hojZTVkviN2n6RsCUOmr/H7ZaSnk+uPGrfE5wb/9NH41gvyqz2DNEiE1URIEbPyWG4jhaMPvcCUi
iNC1AJ2p5aJX+0ma8kijB7Ks8/aDOpWqoyrzVvKSMCl9DzGqy2o1hsO1ImcU1+a15iEQ7aeaCuYT
KX8b19IGWMC6cgIBNK6oxAVJP1nfvwtw+Llt/Bqcs5Hw9EyGxbeQ0oMuoQOtxj3kDn7DKhBpr0FL
5J9Dq2yLLp934BEil0XSstLhClObUcTTnEnUcd+izwY30vNeW73bBwe0FJQQPjgMV4ha/L9XSqJM
xIEgmDvqyNP18KB0j82bN/gHVtTGyePa3cDKwB3iulJEX32MnQdbHBrlf0LjstHsQBbPqmAWPQ52
txsAiB0FFFqFKltm6PBnfrAX2Pfv9f44wuRTPBbt9jrLoacEGyz8+CCDtpTYnRBEF3QVRZl3oyeJ
58OgE43OsUJLPvD0o1MDW6yWO3yR/lWYz8m3kw3lfpn9k9CxDMa2uOz1ru1/sJTZaVVMxlVuoWq+
/iagIED9vNlX7MSsnq8Pi/EvVirBNIhcQW0jucWmXfrEFpDpgRPvWNe+iUlsQHGPN4DYKDtowrNg
ea8b2yBhdI2VEyvwYBvpoHoUJaGrzkTgadn08mR5Nki6gYtJKUY86LMnOLqjMXY53jjTc6P/Vkav
+8nu4cowy9Vadu4V56ijbath3DcoZS9GDPEM2OXPdAvU818SeAKxDME6h6nTerfh+PO8hjyimwOi
a7zGx+LmZG1GEFNEqGGDI8RtXKKzF6yVYXi/FUkW3h/6mad+xWA1Xn5vBieitvIU2Su8m47WIuIq
Hk1YZpvcacdgxP4JFUa0QL+tdUg83qb+m1atbTxmuqVxTi1IoJTnIud6dUeEUnm6sJEUAe174HPp
TA47ihQOv/ytt4za/Np0lC6jKenvULrNWyfKsW0VrpaEHqsUvEW7/1wYPeb1ff3+sO+rkhhJ/93J
r0NKy/VvxMPfHdGCR+sG1+qCQusvQZ7kr1kbCBOvIy5s9nyuR4wTeCxeUVccgxRT7jR4Wg/OtkjL
B86rmmeiqgRkwcM37nJ4O0byvwrlHazawhMVzE8KqhhFdkAp5zMz3m0AKpxcQvpn5i/kDszn6WM/
5SJCFGzA5hVNHXOeofKGy8TmKx234F34Uu7fms7DsF7ZD2XYrgXHlt4XsO9vpG7gUDCp6r/gg4OP
TbXqT0Qu42X3TNwEBf7BTXpge5tdwAcAuMp7IUSzThuYz3673WQ0olOlTTEP+6S/DujzqTaAAWp1
AbTaWY/C+QgxvfOdJoGfHpqpZDFOaShcA+AcyeYrr+AUWn7oB3kaHj/K+P3o+1374EOnwtgEmx76
c9lOA/U52MuRd9/pDrEK77xjCh4lcso0FZtNiWyAGUjT0xF1R0CFGvZ6p2v5sOmdw+TofK0on/Ky
q7J6ktFO8Bq4q3GjLeeHuR5iiRiAqpVxeLdf93XWNFZbT7JddunhFyWWyYFkEsYMncj5Gb6IuiXZ
HF/OmSK9L99luVoEdH0/iuDuqehfNCmgPnEaEyFptXROzKCvVzBQ0sAHLoViSagyutC7IHe6wEfx
VQNjl7CnFKLKRfK5Wu3HI5wGaEVKAEF8Dpahr+duSjnoFebHrzvqMu0QThedBKUj0jeBpPILt8jZ
FmTUJT+QVj1HhBclA6+0Vx7VX4+5t0UVuWjZ2wzG8PDV69KeLy07fUmn4OXdAy1s3Kr6SH7q0UFd
H/x9WeQWm0dzilXRyBqgGfQ4/6///f/qRoc4mv0NIYM4uRCuw3UHK5XMzooLD/LNg2heMDmBz33Z
aClp2Ov92uwOfBUxXPpdBk7oUtozxYmunUI9QWgoIcdOtkJ0DYr2YtTTNmqHOWe7OQPi+vx5j6DP
OtXzH6io7T3vxg3WPd0AHqfBAMAvibBE7M4u/RhpGNtYioyA+HF7/a4vpY6QaJmDC27Tn7btHSnE
uMYja3sZkbSuek29tqspHhWOk58XQW6YrJAfLwu5qjlxbacE281AJx1DdcGFYHW5Q+rze2LfEx1S
QmkW9A0kVLe6BYa9IBjEG1zTwKVjmFFCn7rOoIlLkhJ+ftGfMmRGjsM1r4/Oj2xsN+lNtnoUxawF
ppUWqCyq2ZFbGglPg8MKE5YHAKJol1G6W8yBl0EUFlDJSCudE1nDymeibGurRzS9iHK2/YOf2P51
OLIyRapQ9unGLup4kP0phZ/hKBGFbpIE0FCooodpEoTz6QVy1Xr67I4464NHOsUih3QqDnYs10Ek
P31RXPKG4M1mDFbu4dHn54ccunEH8AWeBE0Ij6xETaBMBYimp3ngjRxGLbZEMdh7OcsOljmiZzj+
a2DKvWj+avw9P339qi8jgxZfhlpormDxz3PPqc9HvM/8NCW/X8gXv8e19jywPwiw6d4xAWk26m3K
j74SOPAnXbk1Bgot5PorE0HiOdKZDb8p6vMxSg8l8oekNuRRPE9LTT8CrEKp38C5qkaSBfHU6kqM
VMnuleZqsB9GTp+Gzj2Z/oLPqejm/hLCb10JG9O+fnDvdmtgcXaoHsUKVoSu9x1wn+tzxrd830Mt
WpmDHFOM8b772Uv4d7xpIxQ7XGtT9IstkmXV8SRW4cjHbSWO9ioRxmBiiLlgsxg4z2oXMG6aVHU3
r5AiEpMuVZ/yZuBeoCE8rJrqdXhyWhaUZpe+Viej5ScY1EsAUo0xMelntzvfFXO5Sj3TaZY5TD0u
N2lDWoEMBKi2PzJYu8bZ1JNfgeNagHEVXJEo7tSOsZ5QzGjOjntajKVPwNZHU9eX4jJAUoqf6ZF6
FFlrKOXC/5OoRNQE5VkGLxGaEeZth01r4psmbS67zAr3Q5UGfrLom+duILXpz8LTxw79SgXDcvXj
Wj7VNReWrCKmS17231GYAB5AExzsRuZb8HEVXTygxB4HWBJXkIPQSKWhz+em75zfnNd1+0JMK4vD
VRrX/kGO2ZaSViOSVdkKA0tFmT0//Q4u2oES7AAaMzve04ZYgo9BGkrAiccMSx+4/wXjTXTsBsKu
RgYN8sWDfsSur2edgA294uIKNt7pyYT3HnWRqcHaRXf2mkQmczM8Fkgv5Ss6utp1S/iVUEGXkzmU
Sa1+FeKLVj91rfRpuPSrF0AGx5fSOVBaUGMYLBAGY7xsoptmsCeJA2l+dk8UJmcmWv4tjydauTlw
hn4NZr7yIAFrI2vPp20CTr+fBR4X1zGcFhGGXpYHDSXZdfVri4wcZOIBy2+PMMIfyfaVbxUY/N2I
1Nbxxk6CtpTeT0ONmO1K73Q2I4L0/ZC8oHcnBfu29KcafP/ppGqUHi8FsxNb4rs00ZOhg07mwQAH
HHBUN20D6jQG3KQVhXF4RkDx/uR4T8rNg6onGpY+coef93YBd74J9tAVaEuPrWARZjT4kZ19e1bq
wtqVX+tKM7IbDSFOSt/4ZHzkfGGi2G9ugTMwVbH5HEKb3+2nt1b6ZyQO433iEbVKMEt8pHIB40KZ
e5BMf23VGjmZeQ+nuTY00rWrHhqiwY6rBqFnDkBjeTP/u3C0+P1bgJndQBVydIDnsnlYCYyzTAx5
8Hj/XbdRRES0ZnHehSLF/5jeiJDLZevS7bE8/Rzdfxw+c6iotP9hJHakXEm9D8/0GDObAofAKIIj
6nzvil+JXrCLh0mbW6RgBcZeikxSotLIZT1aOdUdY9KhW0jMjUOQFj3XRp0wStgE05unU6eCWmjj
573qzlbo9Q/8hhEZZFkhUWnL4yaZxvLwMop/rroILEcHRuX5jMeGnKyS4z1WaDkAKv36odmpVQNj
beD3HDDac/93ns0/7ZVDwZvCnJnXz3JchmUq6VGW4zr+KmNfsszU21OI8ov+LGae4GYXG5VfOpsc
1AKDrlL0cnqQU2bIf1yRQcDyPDzgBuXZH7QZ5C9ppbhj0ahwX9R7pNotjXDzr6NTlOBHd5PhPjSs
7P0XtOcvSq7nV5Icxxx8lUhI6AGMWKkVNKeni/TD3X5yVZt03SzsZi3PuWoTWBeP4q9OyVf3pQff
5jC61Wpg3dB9rdVLHfuv97F8Uy1azjKTQWBHbvCQHWRbFM+Wp5LTIv0GLJhwLd63rkSVv+LUsr1b
yHwVcoqe7Z114FKUOnozDYhdcMsnC1jD0TUGnt4OjAJvY+d4Jh/3JAaxnhi1G4H4PL99xr+CIC8U
scTNmmcvdxmFraVMNUm7mwNqJHqv3C7V8FymHogAnS0c2i9jUQCN9ve2tfNUKET1MKvaSYVebRRH
u9pIAgrX9vxFmEXj5kkbvzYyGBdZ2na6dDPpG9BrTcaH4wRwzlBYOP+NleTI7MoKNv1hlIl5zogw
DRSlrQWRej2GrO+nRDIhuv0t5eXdfx/uiB8kzOEdA2Ls+e0ZpU7YGl9s1y7x7PcGpAZZUPL3C2cb
I5ToSFmLyT4y7h51I62xLRSJ8Rt/dfPZnjNZWZI79xsFjFYOUWuZ8yluC9wjTPPAsdKV2g+y7OzG
k6HecJxg213EVfHmKSMT+xg9S6l+lw70RWwA+L9JAVDiOEbA4TvEKzaLAEijswLkitFpt6kf9umL
CN6jWVdoWIiqIjXyn3d70Q1CYEE3Y5y4NG5BmwJV4/BaX8tihx/jAGnUMyRqToWMOk4Cz+rtH9yp
iPpabWjpcUPYBLgrGMJydfuPYTUZE1mW69HEY7RwCbf79tDDXq4l6l7kk521ZcV6Fvlq63nUvxBb
vr4HnrNNg0/mA2gb/Dtwnc5ilTi+3z13Yc0+EBrI4yjbmtwaNpAfsOOeEZ7+ERGsQAEg2zhx6ep1
SfrSoom6LKOWtelSOD4Mp33Ax++z4GGyJOtEeKxcdy08P56YJLJQGxi7Ph/GIci3/Ei5SIZ2HK9q
8kPr29OvgC+LZDpAjKBKhBgec+8p0W8udIxydnpdMOWnHizQyxERnBshcdEuG2nzry3e5mK+GAfp
8cSgsXUoJto2a9/lcNFWQQ2kAE/BWrmuEFdwA5DE0UUbMFQsOiWooTIeSJDwl3fPfBHOrhLnvVoZ
nepBJDX7KPkGa30U5tSDrWPVCbVFv/8iVR2qb+909c7rt76oRiM9sgFtHLHQz9S5PQIhcBMOCm+v
2BLL+tt+3AewX8L+D77LZR7iyOrkKP1miP2jIyqTlsAbmj87zl8spqeHnHOhtu5Tj1LCpOxTofu2
0t9Gs/rqJ53MEae56N/CXMm6H3j+WJJLJQTYHWiwOqvk5Ruep7wI5GYHubv97++Fa9esf6GitVYM
2wbRaQ9aGgJu9te793YRrMtxwTLQTeuCh3AZt1a0qdpMxnddaD56hRANkPFHsC3LOiGJl2bqmvmo
6MsWTrSOST/Lr4GPEsaNkkSz/ZWs5TmFi2fvdqYbhgNAIkqdJfpnLCIE0QNbX47TATFQ/NJ+lg7I
XK9oxbn2VX5Uo0EX61oQxqpw4kkovfc1QCHXzub+pJt/9B5fRYHzSM6AfQ2Z9ao/kB7I44NYt8gs
sfo5wT0XqTCbMIZm5j3qvMv1DFn4OEjDSWpkaGPfOesU9tNrEmwyVLC1QvaAyEph66um6Emo6N26
hEGYlANu5Y6yHdr+OYMACQO0eJhqAG8Rw6/6iy1du++cmvNDj91gjOMcu1aeuHS/2tMOyc35AfHr
UDhHL2QyeqaZBWz0Wlo/Otn1oBwPUfkYxPLNM3rpVx23vBETsN8psjBQaBAD3cI8mY3oc5l1N4dP
ze5Ssc6a2DoSAGNTMMd8X4UoBmISR/1GUaj7Kdr2D+AQT1QxIblVAUj9YWJEBBp6UioWBDa+T61K
7vXN34pGDPaoCU5EZ3AahTn65rK5pgW7ebhPWyu35dxEj7I9fzb39uHKj46iKfAZwTsMszU4ZWTm
k8hDzdbjSZ4qHhjeT6dUedL04uhsNyKJ5JGS9EBLpyIri6ZXnz32+omimhk8n8TcPfYkiUAViBPf
hEpbTn0yY+bHe2cDfK3Lx8aH+y4sQr7+12OQvP9oaBeCjedSCJM+KxxEeipvfncAS1x+02l/Uk8C
aDq6XLZwtuoNlbH3WBddbywiM7UI/oOBiT6n2qfs27pWPh7xk4OQ24i/uTYanNcfSq0gJ/HHP+0g
EOqhVbeNqnx4s1E3tLxNWECCCzjjTizWx3RotJnIIwVrkxCVCBGNBuCEuMCStJCnPrV+/B+17bDP
XuKFNXbPcv2vpe6IsYmn1zl0Y3XzSAm9FUsnS4KYYOf6r9iXgbEBOd/m7/yLvTW/uDdT7NBLSUKV
NcLsqaWhcx830k9hu5IFqCeW8tcQJmfkRtHWZcGvCCCSAORtoO68J5kRU6YLQAxu+2+WAHXhZM7s
8G/dwHyr6UwaAw42LyqfLjTfk6jflt/in4GOF7/zoB8x7jkRCz/XeMRH6K3wBEjcIEKn25ss2umv
rhUgHPnak36p9YSDhX7ppAVm/YyHdty6Wzqggx7M40QaMvTp5v4R/bQHy1DV/Lsce8wJcboPQtWa
A1E/SU7FQkB/c7ywkN2588K+g7MKwAGAT0zTy4j4OX58PMKlypnDgq1RqTLdNYXcfmN+oVt0HRsT
b5CNQbo/fCc5uXEgW/liK70Z0zukOyKejBgQkYJqrMMar7gcTvxlzw6nTIX8ttqnC2clG/Svhuti
i5T12wUuk9NNh81eHtZyq+Bhxs9J0M9uxslAnmQqPgf4j3oXUMkrT4SZPzOp2jI4s3eIA19lnMmz
alL8HYl7sZOi8H3MQqCqR8bdNnPgkfvCd//eCYoZpHNgc1ti+8pC1/o2MXQ3LHvjs+ecwohu+x7U
fU7y8Ns0XjwvZvx0yTcKHXqIRl9g1/QjqN4JVLbBRyMY31xgqutMGWxo94DVKTcTInfGOOPIIuyh
z01NjhkqzsHq6mWglJa2djjbJ4m2a5nHkVEqT6TtlXzMVexN3rbdyDplJWYHjjIViHzk2CFRoKPM
q88vXp/crBE0TAM9s10Y5LTt8TjJJWKVUOGkF4qa84IO+0fd9+GRJNaAlIaxUS4fUM3/kES4WvOa
emB7sNSHFscSSerVJ8ucwv/NoSUsPAxxJQ+dRuQaWgmFCoxoINbur6Oj/Mh65ULemMbQv9C0+F5Z
/eEHMKFRyPIAKuZK+T1iatg+LjKSa8WZzGcuSEcH7sHb5zVhYYdaBANuXG+xJ1UPEhVkY+Mwbdye
CYNf1mxUmxuyg6HQ1YTsvKpaCvIwJ5wwMcEOcJpt0JGrKxxu2drJPYLV3IEwQc1dzzbOXY+gZcV6
QlZI7encKd1j0YTg0KBv/U2wOnrzvOfIaCynAiJGXTGUTknUOF4gUUboCtsxGoMU8E+wWuCl5OB0
rVxK6DQPGGOFoMf82xM/YHUMLVmAINug+TZgn4+W3lhP83mvM628BEu8Co76O+QyNY9D4js11Co2
x35RQl2aWBtWDL9b70Uis63mCIShjd+6mxHkcmfBIwKyaLgNpE9wbhm0QZmLlqsknM5zhHdl8pQg
ib3HTNr9QBBq0ndk6sHm31wfL7bkgCqPdrWBTotu4YernAr+uoTcgmDSaCn6+BBmxpX5YUgOmZse
jdKMQCRHmqQjGThu1ZiIPgfmoKWqKHlEG/xCEAaVrPSCJEh6WNDrCK+OMLH3PHGCNqc6+05bHTV9
niTgBF7lcToGevVVM5HmkCnT7ZPpQjRaMHYp1oNZJMEsNMHjb+4vPJ87x5v3y93+PEJSOMuPLTv9
bkgnGorNgV7JvLUQ+1sj5KWlPrnMFXaZGTNchbh2ePYY4869nNcB0sLaQPzttoeO4SkPAdmJ+ERY
sKs5ySAXdVf1n6PVcQrwmpo6eBd3Fmvfss1qBihpRrzPN4olrsg4LvrAXaAi9IWGF82DAafP4kf4
KuHIoM8nnp2cgZ/Mbr34gLxXEUpoAIW044jp+yLshN4PoJD31tBa072eygoqNLj0LqJW2U8TrLTX
Ja1AH640yOmnoIdxqi8kxzaqyk5vXA+0YGzBzSph4SQ4ZXYIlt3CX+TVR0CQnI+clKNOHzykwEDt
DUoDGyAAVW+zXZpRy3C6VLnJMJDkoo2qFdVENLTiNXz2cUcTeFyEW5+ImCPXtWyiS1cCAbWvnk6L
SqNaI4LlMPwDvouhY95iCNx0zugY0sqcnxwRLtMsmeqxS3K477V83hat1tIDhZZ8u03/VxvIyeza
bDwVifRX1zRXzdMwzKRrQ7B++CxJK+vtS7FTSgyC5HWk1p1SN79+4yx5uTiVNz0+ReSS4hP7HGz+
kOgvXN2PSfSGds5cNrs5lx0KHbskavHCSxWCsUh1Y6FGAmYzShIKQNCdPjaGujmYS8yp9Q0Hyyet
L7D2sENcYZuI2udBazT8VtvIwOP/hdB8rBB6gO0XwokifawTCiYT5rhn8Pcy7gyRvlpS0z2r0sQg
hipjocaP2mq7quuv2s0XhwRkWlcluXLDc3Wb0qFILS844wTv5Ms/NiGgSfGqNUEpcMNgjD7J+fZo
6+9JKZ9lWPcZhC/8bYRVNDiVVsZoD5+oZze9tO6Gw1065EGMLv88cmYXU+U4lor4c5JCk+HTjQ0z
D+MSi4maBhnWKRp85lAeDUktqpROcCTC11mI3WfAsHLHGLtpqOevOn48Kgs9Tffg21HlE/PAj9Yn
nzM9tD9mRq5wxnMnD2G/2pNYyi4C4M12zKlumE46M4l6tYeGn1XxuuIFiiiQKpMRuGN/RXQUAhCr
MYBgbPqGqYHCKzyVNof32M/V1+YzpS5Z/yFzm9K2LFg8sJhYpeKio5IOluZtbSUfml0T5J/Snq4f
K9NJKliDBWC0fwBETjvGgakmkGrzK6+MUo008HkNmGKpIEnY4Z2WiuQsjM8lsR2ulvG1SyCrqqaQ
KFVynWCMNfUvMlh0BlYdVMFJmzQ+E/4N5rJNotSFUGiS0GdHSEjDV1slfR54ExjUQEk30OXbJIYI
vRcKD3b+On8D0hb0rPCHxXluiJXurPKx83Bq96BJN8m0sqWtL5mPG/CL6Va7oW5OHPpSNiOZvV86
AUBb4d8e7qF2HLE/yXehQzVyjZmMtmrGHgwsKw8BgxD24cF1Mpf64ZwCs3WFPmAq/StTqiiLTImo
tIGq57t/zzNjPUiEw50Raog1x8GfDmW9/EG33J9RbqPyWLbKl/ESJuoQ8ihIwm9b2nEoJBSpgISZ
bbjB2jlPtPt8roIANr28INkJEtB6Z3S9rVkht+QREaRSUqRHzfld+Uhpi4DIEJrzS2dnwXnIR6SR
bNMt0AQ/XwG2Zkk4oRL8VlnU/Eg4nfplCE1GtrwO+CgzRHpV5uWVVNvMP3eXbQOP5xEDT3UDVC9/
qrNZrpaKSt1G+EOLW0wfKQw86tjfM4MnMRfd67+/uj1DVs0NNwIzw4hmm+dWcmu/6gJX1BgDJcmy
FOc3U/+F9TXNtk8ipeJ2+XZDUBUlnTfusAaea9wC6kLB7ZeeOdr5zKLHsStkQXCX/rnpblBxBhLC
+kLeRWHhJr9Nb8tLajTvS3L7mQuG75zRvCZKHohVEQe+3Hn7A0IyifCK0sU/Qt22swu7JW95Cg7Z
jxvoD7EWD1SyvQpHFubbuz/jCQqMteiwxIe1N2mAz0lqKfFvdonueESWHi0VyyrT+2Z6GB6A3pHz
vYYOr88+BkzTEm3dW7E9j8cS6rtha12GMKg5Me2sC7NK8GbfJEspBjUh7dBiaFrha0Rc+ejiyvs/
KZXbC1XCIXRkyLNWHnmzd9k/w49yJs3QrL2959zis/AweYRuT9tVR9HOhwzMDvsmZJWkoXgrqo0U
Flfle3fjYsERgCYdT+MfQCMMiCxGawJ/jYrZq54ii2ajflQlXDJfBuaPnxEoIS08OFjTCvvCjYoU
tLZ+0f0sy+2KkfN9wiW7rgO8dLsLvnDagsM39wNSK2rHH/OI+e2jkqIQrYlKtfbYi30EcauuRDek
ecB+dNTFrlQ9rgKmKZL39przNe4KHx6aMoIuLVDiqOwyBwqdL41egWSR2K3AFNhMUAWyudZJU93X
H5dumpMo/0m7XG1d9wvm7/7cTEaFQej7nymGS04IjTFS6M1gkrC+aLoUDEpZUKPXpeM/ME9wkdpk
esR6SG+ago6TVIGxhl76pAtT6RlDB1LqjmTvx3AaYUYDFToweaQxjmjHFdgi+jZdfP5WcUkz+V12
fiUYeQwEx0qmUDgbnQkzVb0yD4373gDMy8Mmrs4LZnEdeb/AvBVfrU6MEs7DOQuOhz2viKpSiBdw
iIh7hqCrA7JPDaZxegsVMhNz5Iw1lnlaNAT9qj2Fn7PrqmOqd3wcvUMmxT7e5QKIbUSxfDNhGhQf
q664/+iJkTPBJcd8c28KELbNpbXaZBihxkcOs0CdfFb7hc38UD+IlW9THvcKrHrvABxe0zxc3IFc
GwLfyDtdlI7JVAGb7b+W0/QVaUNs+jwbASOd8Ij3K+QDqwqTBzcBzGOvhYUP84XepTxNliWGFqwl
IKm3WbZEZmmEBqa31sf0CfoNCdLTFthL5T28vqLNt91Uv/fapVz75WZx0PQb6nQEGOH7xxlnkf0r
40+DzN6iyps6ql0RQWnc0EROdgi0/eqBmliqIjtcwSC2EsMrUmyQGPDupdcctlaZaStzGFMdEwvo
uf8S38t4ksP9wrkdSdZTJ2oiaZkR4BJjL6pm7Fp/WMrb1/KUQ7O6oK7lmntJvIMKKCnNXkvmymYN
GCqQhw7nqJPK9DMckRbd6I7DzZXs2JyGEWxzqAlkPj3c0l99BE2kRQSVAAw29NNRtuJcTxDm9XF8
LoGQqSMgpveCX9nG23tgYbnyEIxXkvuOEZKzkU9L/naYNS2m9D9JCRrjP3YbS8MHi+jwe3FtpfBi
9d3cV746IStr6K4Cxt3zLuVayEZ/IG9iJ7G1E59TAIg+hSeFRxO293VyeL/1roy4+O5PFTUFfGBY
aYbVJ76PSRyA8VLTer5LM9SSvioP9U+aXUs6CCN3J8jqLgyxv5Bklv/G14NKj9Cm9QGpZQGcnshs
a2vKLkDb93bqvI8d8Os+CB1RruENTWlS/jKT/NQ3lkw2i2knkkOxlXRJvhMeXA3lKJQ1cn5lrtcf
fTHCsz6evwdJmBRidSscGcwhty2CMappRBjnQuAZvot3qu3iP7RW66UmM/FYrFzPFDD+9rdsV4B7
VnsqVeCOFLnWlw1nXzXHyXEf9qy31T/cwjBFfEMGmb4GXUpQ68cD1ptodkx9bP+pBMmjd6nykmn1
yLJ+5mEBxMyoR0K8g3EWV7tyhmakoXs8OR4LTMJsjzxorg++dOCc8C85fzCGV/MOMEuL/hcWeZcD
TM6j/NoykE1AQL9VH7VcWTI3WsVvd1b2m0opoZ6MIOyW19xPX5o0B4Le8PpfcBKxrJjdzDWtpfBa
Q+W6rvj6Ft0P65eSe4Lzdb9rkVEtyBzFiCoqZWnKeWp/NDE9Pc7zMe8n41Smykj7oNL51MIfz5DV
AU8dGV84tEPS3VWzZQuEHVVUJ3EtOLe1SJyi3z9J7H3juVVOBI7YQUALrSSPmV+e+/mMBAoexbYh
4LKt9jPTHo5zkIXKDrlGh2GY7EhGhmS2kFS2xNwKfTsbxE5awU4a3kX4a6CI2gt+8imjtrN18OIK
dYUYf2pK5Y5rzDfLNWxBVoYWTOhgtNqR03CZXbC5Dnt8BytIkgii+SCN/mgSW4XVgtFSPibx2gTD
OoJCxOqqNWswbN8iZhbOD/L4OD7N3n43wWv8mtNHn0XcttCZd3NuUVq2xIlu8cQ3muSKhZy9VQ6l
2XRO17m4+ZohcCeP7DnsRSHHJkwvxb24Kje+WZmMp2oHeVaKQztrrjiNvdZ8YixzXicq9HGqz3oa
oMlDHf9iK1AT+6XnrQkXVsdF6+kF67MPRj93Xr2EG8StptrgtfjU0kj/FoptlNxbkbnLpMvhrLi4
PCu404jnfTvwUPFHAE0Sw/h94eons4nTHGFskkPT8eDcaOZTXWFa8uJrHBkYuw8KE5fAs7S/XQkC
DhBgDvuhYWY931BB9AgZQ9GLEg0mjOd/SNfd5aYgI8EKNZvFXmeIg16O9E5M0SxKS4biN8wyWnr3
YAb3n3GOa2SZabQnVnVURgrxh49QM/JbShNG+B1OZCzRAl76oSKnUugoWvVwv187LqRjG8rbnKMB
JHpfrT4g+eBW89zqPAp3MHAnV+N0XJDhGr2kBsjfuIknrZy8kRDeOlTBUwINYRCcxVgQhN+HEFvx
r6LDxoShuy7PQNpghxBtJYHdVpQmdgoydESvhyO9aJi2NbW7D0pcLNVJ7VE4sKeRKqHNUBnGIeqH
G7CLOQRTzp2sH42dbCRFUZ47BzMQMsxN7nyXvCguQYG7sezd/GBkiP5DZGkKh3AwwFujYZ//5uU4
FlTaoTNgqiAFKC1fEW3d4RPiEYVwQteDBMqBL5IUUkxo0VFhYDYkvQUxWxvRNJvWRpojaq/H4Gxd
s4y9b1Or68/mWx9nKFW66F4MvT9XRu9Mt1LxCe5wKvV90x2NGyWCWPaanaEMnet8HYye0wZxclHT
gWvtNOIs6ZMsXtiMo9rLkq2Y7zsSaQwoBtXX2YEJnpd2EzI7ZKJvwELB0Z2Nb5JqPepK3xVOqOwA
il+WcuzHMSMGmMqLm1DXP4Rwne2ZIJP1nCM/9LTRsbpIWHYTbqpo95AVGoKgJR8Y5AfKb/EutOsh
bYHNJuSxzB2Xi3U2rRTLvB4I1qARKjsgBYqIoRZtMhpeyS0VgIZ6wxlmv8Jnoq/gAxM/5L3UbKuY
kILAJIejz8dRoyB2U0rBbuvIRriDC7K8nUyJ3SUDPDrXjUH76Hbww5txlkdzh48Ri91kVd8Yl2ol
PWmJTEWKwu8ANFi8w5PS3kGEuiDzXg3zKs5dTnlOVta2AFgNLbd5FylO4wjSqtC3vKZIBfn/O3+h
GnTitAdYN7RuVqH7r/SzvcaVCDdaDucdJeI/LxT1yJMJ+0UOvEvTSGjdbHmy4u+a9aTkT7iVrTP0
CXGCKDhOsXsplm+NnYLBZd/XegaNzuDcqRbZYF1G6BuuQvQrl7qR/k9mktCtKNV65Di2QkPb6/Gr
uQwQHpZhcuZC5VmoBpjfIB5QVyrNwwNVHB2gOyO+lNaq7dmrC5LD8l4odYu4i+/mtSk42NWMJ9Rk
panVF8019BGQuAfKaqNzmXQunTj786ePbdqsCAOzk8cwUZOEezZcccHTnPwqROPCDtknIA+i0TzD
Lq/lnpC0aRqa+IZSZoAFrF7MKQ7AjCmh46EBHSPowhs1YSd5WyF1UlC7et2qtrjONelSQ/J+Gv4E
f/h+80MsJh6Y8Iy0Qdw4uyX9ZRj2M+BULMqEjHHTJ1LXagu02iSaPhKazueCoRCJGPmDyLtc4Hm/
6taBreIhWtZa40OAq9s1NWhjreRelQMT0HmKxr6r1jsVjkCojqAGOQu0dK/twAtpef5XMgq9Tun1
N7/YdBvumyL4aG+qaWP9ITf50OJn0dC0w9I++X9D/mO/oiM2seizoM/7vpeSh5wjJlls0BzSXGWF
mKi/XNq63UMlVIFg32gDMxwBEZCANcyYeyKOp3bxBg/vcmR+1PqV6xpDOV0oEZHj1UDaFjqhdFiZ
1/FWDILBlvJ36kusSCDWDBnmRHcqPgTce8U0RQ+xfQcaALvhYpDFrrq9s7xpjKojylGt1AToLhdh
eLfd2eV1US89t2JJsCy3BhmNluN4GaDaVeQmIjwvkZaf8W8pZ5lDBwPjPniklFo1V2JO2XTAiMtI
PHlowy+MDshVQH+/QJQdyoFoQyvlEw8ID59sdmlL6gzPQLB44Uash+jtWlKhcE4ES5yZSx27piOJ
BxozekHdgRY2lEupn0fh1cRK9kKSQDBCL9lJ+YQlgIT6CCD6pagezzcrk80wLcqy5+sFJzC458Mf
kGAlRZaLepoK5QqWteIIy2d/3uPA1rEDVa84fr6X0QUK4ym01tat0GOpnZSgMbG9iQYdMsYOHHWj
LAU1hMvfAkiiS6hNMzUwvXMYqgayef690OeUg7YfSY4g5ALCrlgBc7O2gnW/bpGCpt5MaGKAPJDo
Ba3KIY5K/kIy2YvE5eAxUCnySG1pC4ssqgYw3B/GgfF2RhuB3F3HMblUrkC/Pv4o5lSzqUIqPVcA
JwbXBfl1ciWeIUZBlVUPZH5OseUBDjupgQBnJo6lX0OAqjHXNg+74XrPOmEjYUw/vWejsCMCUM5K
8PQQ6qs8mQogyUxlVwK0hsu36ghuBxPWiEINcPIUyCIeGCt+k9Zcp7xGE23VTbuEqB+Hrmn+33Ju
gWStC83FuS9Z+zUMbV7nyEVCpRR5ckujvSn417MQKOdoS1ig/XOlbEwW9Psksy0bRTxYatWOsoPQ
uPXFZBug4Fk9JPwCxNBVoRwUnOiIJO7lPKk63PKJE6cbyNu66iUWLnC/2GLaFdkEGuD+it9TkehE
7xNEQDOSSNbRiRxnfdL/YkM5yCNMHJfZwBMxyjm3+p2CknrBXSg2WRo0rGbIo4lTnraiFW6TN7/4
+YAJ1GQdKoKYiK1DhxeutKMIoC6DJoy1PMavUfMuHuNni4zaRkPacFiwpojrfuWdqlscXZ3Q0q2W
VhTBp8Z+u1t/zltRrbIPcvp11eGpoeHwNNZfj9AgA3tKkvQemZls5pUH9XQ+tj6A4tB/YlxK0uzq
uXxeRURLi+7UhgIFgamPqNQ/2qZp3/TTD4VoHZElTn0JJAjh7wlcHIE1uD1DClaQcxFD4gCg+FTC
NREPHa6CKa0GnqoemZhlni4mRRs79sXznx3Pb/TQxo2FprRDbAiMPEZ0EoF2zrwFdL4S8Z7SgttB
QRSkKx2D77oMVEUcf6WcmdMlxfaKqB0DNz5oHf2PPhd168sFkp5pUndrDTHsfyP6V8M7WT//xYps
OhvOAp8zGKAvcmmFFOngm59Q62Q0AAGMiNWsujZxZ/j4TmNj5L2BqeJekMAQsEaQcLZZLotpQdf1
/LQXbyVsrjnPhhdNfJHXGBtxvljtfw94VQLi9hrrsYMtPhb6juBvHuLx3Qh+cXbLHSQzlndgQWGy
Pjasbq9cDZQPXpQJfr/igPIiLjyYE2DWtbhlfR7vp8+4xFJ4KbJPabRUKJsEZm5F55PqRhvX9hLT
FiRjlmzhi3PTHuhlYHXv1Hpb8TEHY01sgPQ95PCXuhC6GEO8B1qPcH5ScO6K6uVpoacBPQyC/F82
/Wc4cxxoWSxsycNWdPyxV96+gdrqRkuEPk+bqZjby+y5Egu66K/OtZ4A1P6R09ArUvMZBE16WfPz
C1bqeN0yprKE5yCC0HRTFijspLDD6nMOASTIgKVkKg+e/VtlRj8m7jSCPp5lynyBqCQ1gc4GWOLG
Ey8xNgcKOjHTFJi53RlRRQzpoXZ6V1BktQyToGQ7gs31oWM/3VJlpFwhBEJZzq2YfgRBXxJaO0nf
7YHTTj2Cp1ymNBe8jlOhU/hhLUxw1eXHHzj51q6TRKIj0ivPJxel7S0yGp7R9g9T+jAGPHLAJ99s
dOoQCU3kz80D5QIo64gPYevDuV03kFtJrbG/oMUfxjjst1BCUI6pCbR0uGYnpayOqz8IdEeCc+9M
lr3KxcYl8oDEFZ5MIdQa7z8DBCE0bJ6BpDgI8uTYzSPJJeoLNOubxJNLj1zQ1Vdm4mppx4Mvxn6s
PGJ9XpvTy7CN2+a+6ffHziOB1U52//g/rh9qFixOA8Gf1U7wLS52iJPeQy0rk9MSeoo8yRgJkC4A
FTfiYWYG+uP2wanPXgqdlSxYDJv4TgVSS/fN+LO45M+l2do9XUGjPzPggqy/YDFf3amU4S33hSO8
2W4+Js4DeDEJY/LVqdSHzFI6+NT9gCFDePSWu/NKpT2OqE8+5UB3pyKKMd7T5ElMTFGrzyRXk94g
FgKNoaGLcJuZAKZeyAXI6an50EhvUQAHd+X5aZmIBoDEzfj1B7A2liacK/TWMpj+FbIllbg9dfKh
VRo7flnV4WoOn43FKFAZhTPi7bTXw3XWX99R4vC+hcQ+xNI3ycWlt7M1Iwj3dHMaoa0X099vFDy3
MK7AyonUzyJHmJPh41oE4kNwjvtqpy7KWaVof5FcPfk5O3iu4cOlbWrzHCxWYt4yyEmHwickE24O
xbTFSFmDRTpcprvczPeIt7WwXGeqrv41+1bzgjrdsNBfpMMoXYI+P7UQNjGsDruVrywqLayPuS9O
N/xjLOYOysPL6bCw/FTwdLv7OcvEm/WEBWTm7LvdoG++rUeRZRu3AhglFYpGr37nbVtnV6tvioVH
/+ZcZBz6nssaXHMRlHF/sjBluc/lxg/z/4wJJoUAjoFj4celvn7V4fUk8C5pt/qZDcR7wlgFmdHR
AI3WfIP4q2Pv8RM1H+s7mL0DQqhwv8RK9BK15L/m6FaeoPu3gXM7tGkHlRicf7ZSRmDWnYqNOluf
84TFnLb+CB+hrU4DgSeVb6IAW/S9aFQ2q1zZY0eX3X+ptKmp4jNG7KFX2gH2Gfp4mdJlZwWOiulY
v+FZrPGpyudeAbwxyaJTe2KoDaA8Nail1D7rdXDJ8pmwfpA71f41B6SnqXNoNcWmojzf1YZQtCmg
+0yfsXENOQyKc6sPJSCtBoNZ8ePp1n74LEwduiWAsUMQ9+Aew0+FiY64ls5IoulA9w+eBDuhFZAM
TeqGdvWpbVPFp1TFlEpaBMzOxV1EBgLTwiDvNR6p/fyxv9f9X9YupZ+YoijxNJ/NkLNYO00cQ0z7
smm+1ePvpfuS/5y4ZO/381jnW1GLkFWDKRYkHjRDZOTMN8BBioxZ/mHW8mnjyTJSdO+7rna6gq4O
98dXePB14MHp57D7/15QDIgW9fhBhWqtlHaHAQjtyPOSor8ydixGriZ9hj3aeedXXizex0WqYwVz
Y3FtIES1JhW2UI5U41srIAGoM+V8lCCR1VhQIt060eEJ9MtkGL6Gg0/BGC4kG5yhGGkv+RQ9LsW7
2mrkxzPVlWybx+nq8KCKbIbVbSFOs7dY/mvGS4jCA/MpVMi+T5Vn3i0yIXi/96AOL5HzRKADv1BZ
Dl9YCJtZ7nQCfrZB1jNZGtYFjXoZjK+2JeTVoEucW3VW6aIBGzyErs3XI0JtR5Kvzntwjk2f9LJT
wddZGaU5AcslxLjsa82ekKYombQCRqXAdjhbomQ94BMH7liXnM04ZaLVqUAQUPCVErVAnYAR1MUS
FwkyDkJClM4n8veJ/IoufRNU5z2SPKF2YZ7kEP+2EzrjbA/jw7drVJsTHXyVfie2IAlJWBd9p2H1
edLubf6TmRqJCozivNHjTvrn6VqVYxoeYwGI34j0R78ddJEJGkwWnGVIEJIpOBtW5A0NOh+DyhZ0
rIqDzhkMGVl3EgoBjnjFKnEMJXjbTMe1WB+9O4zvDIKXye16Oyf9fU1F9l9QSd5wuDbNcZiIMLpM
1RBIpCE9AydqBbLEWryLLIQ192AhtuhBFrfJLcaNtNv0mz8CxY6SUGR+4KQvWEwQMslrlz1yku9B
mA66/gU9+ZLLAWRa4tT4AyQjSuAm69s2wJH85NTjpX355v7ix7DCBY4d5u4Lsn2ZsLXtFW0jYv4N
PiQLUcR/CbYW0bGFCO6Mw/8JroIfOE99hYpklIGs61f7M66dBYirpMxjOPaugpu70xGgOhjLKsPG
PQFlC0KEepFfnlgqlQR1Yk/P9f1D7umSd7jEL8YVAf6YqShKbtJ2FfhvRegvmd/nfogQYUG88I5g
x75FWj7E6b9E8Cl+KXXZI/ZMo/886IJIoN4tqSasOMv5qe6nUS/RWgPsHb1mZUe3L+JbEBvrfVtS
Le5ipRE50EGwmb23kjwKzTFQF6lOEedZksAD+GASqdL7X6G37cukuos9QMuTtyW/yMEZlPS3P/cn
Qxz9WTmUjiPJwINaKnVwBq3LQkdouFtJIBt4+S386acqxgYG6jgJJE3mBqL+hbzXHycrEKGFYJhf
rv+H815p3iV4f6TkRsTxnL44bgLt3KV0lk2jA1y3FECTq02kJjdtbjcSfxgNdmFqi/uROhKklkuq
6XLs0XN3zZYuqK9YR0z8ZMS2QFoJKgD/QBH8gR628xIuSzpvSehVy2+BNZ0tbY8UWhSMMXUV2JWm
/ITa6NDzJqjrJhHyiSL0QsHAesSbeL3CsG2SdRQFwG2mKNoNckZrXUG3yJqlzc1lpU+ZL4xspTjI
KP6GiKrb0TjmWnTwBbfJbz40SAAFfkf8oAxL6vZO7mcrSBi7o3GlPrO1HCqVoe8fnxK1SYpZiRad
SQNQzdL+5hN8MS0M938uMM+svxNCZ5rnsCwHLx2DBIsQ78yBoRdhEImxgW6+Cye/c51zH1iWE429
/K1bYGRws35Cw3KZsPt+zNbzWEpvw6lNfB2Bt3DWaYPWL7H2jb68HJPY6dDfa8cqjGtoGT8A6bWl
XmwE4zkM0uklE/8SPqPkFB3tj/Pvr7r5vNCGbfFWWYKm4ZYPcnmfFHIMGPpyrmnrs02Xkgazr/CF
QAWT8G1qQyTrd/ASfHhH5/dvX9CZmlAyx01cd5n25ZWhiXCCH20rr3U1zlHZ90Ho0pVu1FCGfO3u
W+hOtOIT4l3qDgvzmKjXF/Fw/JF0degqvGLNsuO4g/eZE/RRe2jjYcQCqhU99HSf0NOULkUqIbUT
K2HEB+4W4wBn2kQpEaWGkF/3A4bVRTb2EVARMgvPE58eoFbvTqtjj2BfX2eLVQig38rzDu5p0YmZ
cuIsWIqaWyHutNZ12eWp1NI7235wcYUh+rakJDzP79QTycMmUjLngLjPcOScD1AdS3IBb+D9xv1j
jk04NOiEIGDolpKUPN5+kZx6PA1kW1u0BNvnQZWdesF9qFnHfneUghTttx0uf6AosU5Ckc9AiH4B
VefEpyp3LD8BHCOU/yZ7eiFhzOJURG0AnSnqyGUtaPg3HCBhOYLuieMhm9mlxKrqfSLXr89FmbPo
O9J2GMJvpZq973LVRr0gD/by2Zy1GYnbQnarmHrj31Mq0QHI9+++UE4EA5SbakoOwBTIHupOdN9C
j222nTY4hvWe9ppQs0tkkThSBTRDyjkTXyyd9B4fmXEcpoxG2hSCLnArTPam8kcDK5e+MIID0x+L
NhyM3zpQ6CR0bjx/i77USuFHz1j+rk7FBB7ozuNMMyXm0HQS/kyWY4kQl1lKeWDCMfV4HRvzYtMA
psijcNWxtAt6yRHbu6W9m16fRipJOA0W5yTkRaFSoD9UUXMkPQdI+BVixmXBrBk2aHVgMs6nCZNz
FZl9lxSn3wxVYr/GHMBzJMt1BrefnQPjBjG3OI4xbgMnixvoxr966d4yEDkvLmo57ZIQHg09QLWB
ZIxyD/NNO3+PcJvyjrMWYNVz44P3Wk8PoOYJaLFcUeQlHN/zAzc4m1TyQS9tO8B+DW/Wd37m82Wi
jMZHsEjJYnprwTgooXMF/o8Ved+ggou1ZpIHd6Vh1AZDrFC7aQXoPV9lFh6cUY6GKA8M8L7Uf9Pr
R8HhwjsITf42U9x6pZ6ewNffulzgTAktEHCF9XQZ1HbaDIlE1T2GvxQBA9lIAyjxN+H3KoJxkCmD
KqNLo2mLsD+POMG7xL18PTZsDLev0E9kOokLm+a38+H1ApOnIkATdA5vemsEcwRae8uU5iDKzlms
ntSzr7yomzSQ2/4EyL+Vc13/+OzLRxrKcOVg85/elqmuXVtu55pyJjbUomjMLjsI7puRf5pPZmxY
IJpeE/GfYMnUreVXf+2l43K9FCZUS+keUWPuYmrxDZepXueSJpFWFBJ/C5hgD/ZvSHzNj6p2ztot
WRHblbiIa+ijOp0G0Oqnft0zlaVMLFHU7bOgvnz0H1lcDZyBpLH/QP1yFtqt1odXQgrsOlaQIP8x
wyiODmbD8Rn5G6Vkys9xgIq1Sxa7eKp9TRx6nZRSt3YAVCZyr/IpuQE3BX9oRxohRJ1GXzkHtMQn
wDpxSVGOoh+YfX2mOr3gRf78XxTHhHpjz7lOWmLoln8/UhJ4WbuEkwQ8WCE3KmueMh8MpvpOTT79
ychM7yKNyMvvBQUeFfPvpQe3ou7kqrBnNruOtlMavh/8XgN1ZImFfOl8fFs4HHYTN3iXlwP+C6F6
I+DRAhN9FPsGO09zPcOuRKMgn3QU4QnN0ouesXDub7JCTIkduMMV9HRUfl5/TRu2dIuGnxYbmVNy
QfS+8JItsZFKyEGYlu+MJzR5k4d6gYYCCBtejyZ/LL4h7tCqY215P07sN/NnssR3LrwMnuF93RxC
bMeaTGm7oeOzbmX2KNXDQ7ZAArOTZHvuNx5wH4u1eLRzomywPleO2NJV/iMRvPhM1IHDiPtudX2u
NTDoAZG43sUhiBGH7J0uDZeN/4TzXOefefWQkrZGjTR642hdwukYDdKwGJTQ4kAQppjyKidyjOf5
+1NXJliwNxjNjvyZvFPNgPh9JQv/m9rF/04bRh4HuQS7A9tP1DZl8cK8Q1RqreZt1KVYwKk4B3js
5hEWS/V7fHICwo7re7yaQAF5ceu1MEGu2jm/RGa/ekaMkgHk4ml9t7xGeJH+IG5ZQJUgt3jyfOlP
HepoZe3N9eOR2xIzduKy1nC98mjyiRR/6ZSEruKntL5g0CB7DtmksqT5ufQneChgMR1HQxPy0B3L
hgs2IWRD/jX5eoRAQLZ7GvhnvmUpT2Qgtq2yCQbvRXKWckQjl0PkTZ96fmD84xMWwG7nATlbU9DJ
R/UXeMHY5zuaIhywk55lbreNT3W9f6DyIVB3yLO5NIGZNC1Fpa6sYepHXZY98JHfGREGpk04p9mu
0NOYBLP/eDsa0j8RUbvXeiQwJxZkc0sgt3fr3zGfx7QKPkxCF+szIVrhtEATRVMnrmOo/f3I2c3A
D6YiPkmSCbY6q/8XwEh2if2j9yeKx2wRr4+QMNpfhAcj8fvoI5PHNWL5HWjunXcnO2hGLLVBPJ1U
nDxg7cR+4pNHEZdHMxb8vgzO8KYG+S3LalrzlpXDi4wIYXoyAh06/6V9V3OtaplJujeZqs6ehALH
8qUjVivjogwHG1CkDjaWkrWd/h4359JUe/vzP3b7UxADJawUwvkAlyN8oMdLDmPy9rsa5DlmSNNv
5Z19CvPaqvkrVScPZVi09KchQyCsk885Q9RIZw/zn5Mj6+tQgRR9OCbNLp/K73tdTHLL+R7dH3xB
Rg+k8kkGNB98CjrFhxTUdIlr0BFltN/Swbg07hHYF6WFoYri2jxmj/nSOpWDA7CV9KJyl/bciXZQ
FgeEcgWJ6KUw4xU3Z4lsAI4v5UwoCQnsDtRfaIuXR63iC+PGr02PKv1JEFWOslxOIOiJ1GSxtA55
yWiRzPc93sApR0MTe0ee5YeYMbvEkqBHJdGxzQTCJfvbvuuigBdPxwX2f2rVJ5gXDOibcgQCjquv
6IiGq/L02IyIL65fHR7jMrncpcvHJ/r4S2Z+QCURSFmz0JVikhT+zw30yHc06xpMy4CnJvXTf33d
Rc1HHlEjZ4q3uphZ1mGLRr/Wyol/4AjzxS+B2BKRLoHkgYLpgeuydjE+R/xXX9VytTmjb4e2D7Wu
f0skHeMrA+sW5d+TGYPWVuDRjqs7aB1GY4ckTvgheGsjTd4RFyM1jB4auuFQftt+vGyRiLefxGjK
IiWtSnCfi1+OBbZPcwvfyhJfeAr5HhEYYkCzBZapwWfTfwFBWp/mkrU9P3AmH1lxTKRFuy8zKfX2
wxTqEOh7qPYLSRdHf5UzzyJLNzDP+oPpqdNXXHT6ZjxKqGpxczSSZsbQyBLw5HdPtTIv1GrJ8qf5
s5PtiS2XDLZj6ngK1Q/elnEB/mcanC3EpoaF8dD4pHzZV6HePOMrllcf+tUT9V/WsJ96dleHVELZ
yFgtAcag1s3CagLzzqm+kKn5Q17xhZ4BE3yRKajKJ/W+uTb2lPXZ2a35L1yMnyeRVP1Wov0GMUGl
g/8x4p4X6B0A+25IfkPvHqALIPrGolLLZPbW19kQzpw40c0DeFQCf6cIDcPLcOgXtG35+MMbQ9RC
XUE0yaCv0mXrV/WBZDvRkyliIqUU1rMIhmINUltO8xXeKMPjwY3eQpvgkBwSbt0tLbwjF/0WIEja
9yDO6nL4S5BlJOOrRow64ytFmxTs1GvGiEzfWWgzbn8lbSAOMvg0d/LoYr+XpxC9ZnwhTnhFh9FC
UmD5PDfEOWAYSd8F7KPEm44u3zpjh6RPNJ/rXthkPGXDBwf+cTokqxh+RLoNYMGHYNPYN9uET7jd
f+wKPakLllDLf8FmquNdpVQCr2/qdabLwIF5Yv5iiRA5OVN5EUx4KWwT5/lgyplBLRF9UYK3xpdP
UhrqvnBNGiKIE4CBRJk0HGgZG7iEqAl6snLIlPsMgUBkWwYgVLCrDvDSzEA1kjHaUOzJ26nKMa0d
GchWse+UJvNiKBTI9aQfyayQTND4pQTj5LXAOmekpo5r8nmlYsBXd8UnCnOrDULyiDAWc6lwKlnn
dkI/uzVMeAe6TsU8TH6UPl7HtXZTz0XeG1/itGCQhC/REWi2OLSWLc58uewoqZcAwG6QPwAU65Jg
tQgem1O0f7/oI9yDtF9Y/sm2q7cv4QcOYonnrPct+kCTrxBVQ6+jIb3II+1BXSlpVqg3LOQVKNNF
oOZgWvFxnWtlkM3s1QuMlTvuLMYj8e0cDGzi3E2omqPg31ktVVidgyFS24X1JDJ7rf3eYjGq/gMf
4plKmWJl9MY0sxeLQJXBEAYUQEVGuCpslo71PxKpjwqDgoUr6brOoY6zqhlxVlc5F5KLSSqQzmUi
Jgl285s6yl+y5nDWGScITkYyxGMYbBC4a/2AsnzVumaU80fot8R6rk1FgHiNbBEAgJ/scXJz7skx
pF/fjJtPKk9YFsVa+jfBDeOXJb/DPvHhrqwO1tmM75qxU33RNhQ7pIdH41KnbJhblxM8E8JsjxNQ
/PM/OjEL2Cv55kvFE/ZoVXjgG4aQxz7JisovDrEJDIM/3Pv+ovPV4WLiudEkVv0jbicNZRC9VB7+
KeLV2FqB/f/QKB4My9pc2/R9MrblyyRSj8bLIG4WSO8Ddb+2KkKesifhfIQryROxVUCmra0bv76P
ramBzNE1y4Y+5cKE4FRP/ZcrNXEOmM5alUodmB/D+Jds/fUvNfyucLgl5jmLKzD4vSZVbmj6VjV9
iLgLb0nMhI30Rr2if3Xp30ov74UupMTeroDHhGS/8cMQhVYWmuCn9K6WbOmiCjnEJTHZH90VNCka
UL7MbbHU96LpxcHADyQGIRcNGnx9WS1q4/9a1fM+MulA9pvafjMjI240XC4ZPlTyO3nVuUp9+dU+
8pYubKrWi/Usrh7YVNST4qxEumoc+HiwSPn6baXz1QBwf3dOhOEEHaXoY+2EOCJQK2cqUU6i5uMY
phoAbNNaJjXTQkbPhVSq6PRBdsY+cVoFhdLsHmXXpibToVUdqSrYtvhXKlcLLg63IswQ7T5h5/rc
xpFn5o8KGsqKDXKsvyTiDL+JVa0DOzrk0Qhkh8r3+agBqNTjfZOcTSA9TOalLeJjCLNPEutTgPFI
z3F6IMPrBX/H8TiQMQCZxjqdQyvUIqZ28HPrIxRnK1x2Fds7lXDx7jtOXazxJoLkuO7LHijEXLMX
OkJh0zj12QRKd/pzMzvtPR2MhMkiedltbV8OvfySeglIl+OETw+Fd6HVifVEzfrPZEWS5EiWXpwi
vzDWGSrll1BFY6nrxM3eTlvhyjQmqlvc1TQtFBbOdpRAwbhgj/Mp3AQuaC+7aSrpkzw3uB+0G1sU
xrVzxee58i2xljv6uaX7X24z4mV0k6q2SKBQ1TvlU2LifmaKRCkoYo4UUFSOHD4WQwcScGx+uabA
N0SNRSfXMNGXxZB9LNeG13BlTSrS0BPvn44s6N7nc2Ijx86ZpMkbkYTwOAxiXA5p6VtxWJddS81q
hzSDWCUriml8vsdSWZOjss3gVjlhf0xzCJLhSyyJ93xmGIxOls1kxdicLIQijB08CFxXFZ0uWBlk
JrH7Ss0aAR7ToeiXG5jqEs/qx4mVmPCv4VdSmr7BoY0bw43um8OCn9PMe3T2MZutfxJos4qCJsV7
C7d/cOH7q1vx6lcaiRO0ljfzkaJlpUtDJqo6J2oE67aXo0z4LaY78S/SVhRR+XuloRtk6Mz2dM77
+VPHGA3bQDpNnME7dDwdLESARycPlLSYePNgzv5k+6KOA5ROFlVSrNuYMJpByUuahklPgBqYGvyp
XN7GqJZxFEKUjw5oucz4wzfEaO3pheLXMkD0Zh9ttPq6ibLidzZNmFccgKdck8AqkKEJ0KSAL6Zy
3QRzg6m1n47pjvJ0rnHn23Gn7IoLEMN87BYs+IXx7t8BLxShP0AAlaTrzp6lXF4h590G7z12B7r7
iGcm5wghkPvqke1x/LYZL2qsPQgcNOJfvbr2ZoqH4NGLq/RMkWnS0ODnUJLUTWEjWOnPZSyZtmjc
ZHZD3abdywk8+zGIxB2WAEO7ykBiP5S5sdw8YJpV7Bsqg3j3+WuhTXnNOaGgcAvk0g5+H4FARogl
us46hlYyQDSvxjgZH76qi0tAINStMKs+cy2qd1aSdpcKx5TZXrGec2e3l4kl/WIfy8YJ6AH9UMmg
Np73jm67G2F6Dfy+0jIOHSNznkJ3XaHXXlA979BfIkIwei1ajFaekdHj7AvBWXJnK35hGt/LjbnQ
FlcHEDEKDSpfhj7lj2/gN8O2gPn0X+y6c2MELnnd34VW7BfWS8/Ru5yqbe0kle6AhCMxxSovV4xD
Nm/Vu+v5GJbSXaqHl5G35GOm3htXPIdvubXgZi9lKbi2Up7Z3NSGnADwTHM5JjGWjSA1Ty1/qIL0
3BTAYUj/tK+p4DA9aM/lh4KP/wVwenSBLRTtb4rZtSXiR66Tb28E/MCVgBwqiIe4Tcq8EBHiW8Eh
JmWMvMOt0kWbnKXTB8So4LcOpwUBGD1Jpb1O3jXSErMXGWCmDAqwZgMwW+ad5+DARyC4rlwV2D33
4VF6s7OIf9+WhDJY5Upo5huEkN8jYQRhGf7fqB9im3+41d9nY+zE4n55xQnjBVNjpSDtxhBVFAHk
f9jugoo/LXktTtJyz6gDkvJRzZ3GSGpqw6g9KvjYYxAQzcUFHwoHeCopPmGKJYD3rdU56GvnMFlr
QmJcfdo8MhY4x9kKRl1BV1YIGNSb8HaooLD9Fc89vzxZbYhnGSnrXXIcvViyb41T3iyLtaAIuKo9
xpGftFqTomnZDKxfM99ubsoMQ49nWe/pyf1L82KqukypnxgnLQT1bzpJshZ8AdXOqQporaVBaujA
Cc71QTWT3xC5ix6gXJWzKMhBk8NE23lIAYU+yw61l3UC8VJiXhcTOFE9VL1GfMJtsIE3/F/8NU4y
lklLYnF/nqWfbfh1XDYvEqZ5ZKfL78LpiqrP9cZDxCgDZH5ThtTHVduE/ueyu+BET6DZzKWhs6fA
9HyxeLkwuHzBn+MNoHIkZsBMZ1Yv241i4pjzHN0aCNF7zXqM2cFo/DTSU7MWkyGf+M6HeCU/ZUDD
xasgJEDYSzTjO7cULiOBdCY6xb+dN0P5vbYjawhZddj86Mex1eFRIPMBEty+YdWijs3X+uc8p3Hu
jUGJG2AOHluO8AAFoL5JACtQKEFVFx0BvkOaFZxzOxMOk9IDG6KDQa9etME8YwG5yz/SBK9oMsqQ
qCaOB+/oZ4QhcxobM5qelYWL1ur2klbK9vJYEuFDtJbXkJyp2SlSW0GzAlqFr7SZU+NC9mgBxP7j
J2eqpSovIN0FRr+LTvSm481v7p/1pVGKrvbkgfP0m5V3skFxAsEDioy8E81HLgkxNzVHxaLlnLu4
O9PeRp8p4r6NmQI+LkPGzhYPAe7TKs3WwQFh8QIpmNXxxkPf1+EITynnlYeClScYTL8RFYk72W31
x6BEtOKcKuk1GffGjfvnjWgwNb191+7pVTBDyo+tkZDvZ5sAvvw4yGYAfoWWdlP1P6dS+tiNR5ID
32pqKWdHDv/5huI3KB9lKrbH6UG+SaviG8rNL+llyQ4KdZNGa4OzfHWq+54K7I4aeLvz9f90/+ko
kE5A6xt+U6lZRU3aBrYhFzDBSMLMp1zYwB6B3EoO9Mp2w3g0bMIZy9+VcbBiVScvCSEm8KMH8BwU
l2dQWMJIjePSkInoginf2vTrowSCtLNG5dEHYIbUoFZbj/TAm5CeIsiRMW/IUN9UXs9szXppahdq
dg5YfeKrqULEYsY5FiGW3/SZZV8HGUSesMRSQZU0KAQAeT7as2x/6UeIZTbRWIVY48dFD5QvjAF/
s5pew+JFpunJp9QeUHYQxG19zct8IwWLkEAivQ8btZ4fHMnvxvs9fatP7VMeF07PXDpSfK46+llL
tuR8nrdZMnSLAricP1L1qHF65lAXyjDmzu2lPUBwUlOyqcVHcnU6106KWOuTWNUzzIl5MZX1FfJ7
Nzpih9kx2c4vmvjofuE1OS27TGgnQgFW31iND+zkHmFiQmrBS2tMZ/VU7RYH7r5uhG1/xQOfg/6Q
xjojJGQhviTSNL9st+18AVhFa294hiS1p3C1pAiRhBQ0vniZopvTYxPGWDIWoYfL/SMyu8M5UaT9
3El0ZkGaZ6Il/sZgfIouEAha+7Z2zrjb9H/3rI09oO1mLxhdSRtYreY3DJXneRpWE9LJyoBruZa9
AcQQmU7ikJavimoug7pHlnzXCatCHEkB9mYAWjrEgdz01p4r7+WbcVxyABn0EHlTARECe2zASxRj
20u94E3aacTuC/GYQWBjPfnUcWxjTVD0mGFjl4Yaehbbs5EdJFWaIvEFaLPtBh3Y3bPBvWsYMyYJ
2Z5jGxd5FoM+URagV1Mo5FkB/nxWcVLBwIkef1dOj/eiF+BS1PS1mYhiWyqqiMHP91cyWiRWbCEG
Zthxk3Uzl5oUuABG4nKxwtZ2o9+6WBBbywAzsUuZkOhoX60QbGUqpHt3UqQWTob/mpxrtaSGR33q
ACvoAskwIhljsZD1CpSAn5RuveWiq1jXzhKmuJrdleNvVAfdxaCfUPvN2f6Zy6GN/+PSfqjLOIED
safQIVW23LT9EkWEqt+D9IslxMGTGpijl0mdBTSAo9dS9h0R5Ve4IAUQc8AKvDAwMcQP3pjvjpRT
2Zy4HqiYbrk3R91h9VlQo41SVPeb8leeQPzpVHT7yYQTL+QlpjrF4CKgPXemXnvkFpVhVHAkiqWW
o4HHmrnVT3iye3yxQWhsS4t1JTOXf1Cbs3tlf1l8FN9iwXgLfa1QtTEOyQsI4tQ3V7HnXalFs10u
YNxEShrQFH2Dup8u8i5llmGly4QI1tW+VGFzvUbFoIF3bnxy6i3zh7fyyCppf1buU+7Gg1R6HfZM
YHxg94T0+qm3a8sFxU8FLTk6nsWzYjyFAFKDZjnOrUNLUTfWrNBIEK+1HM9FJQA2cVLgg4FRdVOw
V2VWmWK+bNjBYiDwJqXnzqwWEF+ydwrfWu9ifURBigrvZCiDs1xZ8AV8YhaDAxaS7G+vEoypjcxu
m4LF/Ofe43LDMXrAHH9/m9yk2AO+vwaq+5ix8rSCJ7RhuM2z0PyaICZJQwvCQkaYrOE8zkVphgop
4wc7FUzN53dW1Zl98MNa5kxUCvs37swCaYp8d/z/sI1BcXhj9a3f27cXrpDvcI4iTGpY7WgXLPJj
PXxaQ+ahmb7S/azrzaH9boyElPYWVSLqvEFOaxn7RI7kCGFnN+/D0BMSqPN4Y/E7XHlxG9j+krQ8
rTFrg1iYEPCmOk3U/1rzas04lJ1WFmH85a6eIGadyzv4yhVdWLaiK5ZoQ/Iuyfnri5yO4KEZfonU
EdIlJbPF91Y9qXs7TYKW1oWw0ZuSjCoY7pcGbjbMtFHzsoILtfFDISZWaKdpyBi6nCNpDLblQGTY
s2GXr+Ern9fuERbcX4aMO56mdIIMRdkSPjOm6KfkTbV2QyhM2cb1Pnprjw/C8s4vz0oCiObJIzaR
+n4JIQ4ywohlYks=
`pragma protect end_protected
