// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
tMfaLE/1g+GLi8NexvTXLCDQA4TVL79gz+Ez3uWXHAhQmwscoMTDS3CcvavsF2Yi
RP1e4cZGYZdNlwmtgeUQWxwClHrvVHHnUun9kBWrl0EV4iS/PcPa9KioZH1iz2Aj
YX9fjkFioF/uBQfBe0oPQkidUAV6iecwPx0bFyfdLEw=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 26496 )
`pragma protect data_block
eaDp7gRMD11WNlqjhAuSUuO84se3jwCBBEhwvbuQjP4xC/BSDE4PZNbiHL3q4Pk/
dEIvGpGY8s3hAoJ3sCwhpmJGQ51vPebkQDXkgUF/gX7jyoq5KfYhpIc/QaBJ0MLN
AnqTLJYgz3VGyf1lzpFRmrQayobWk9ZZxDoHEYGNisSjhMsvlibQelidBqIq4W3Q
e34FHO5tML3oluGL9JM6fCCOlRZ08UC3AKYHTQPDG0K1AaGfTDaKYu5Bf1ltAbzG
xjJV9ygZq7dNTOV9XB7Ixe7XC7qY6tcUqVGc91Hag/khdAhrSbayFPznv0FRD6xO
M3iQOy6clQdn/wb0SoFbVNuJrL1NW6nKZOWt84N+IskYYjmt5acO2Yqekv1tUY1L
5lJG8B441oebGZKeC5Jaw1xoGl1R9leFoHgaDOdhwUvXtGZoyMOGCaP0EZUmMgyM
AqEy2TqenIqdmsH4zW+ksFj+/dAueW6gBSyGmA51yYaf50v9DUEQMc4uTBvKh9xl
tqjy6Dfv19tGTd//A013UUl38WenIQU9WeLQGJrh1lAg7Vatr4qBCYLMG3TtYuUE
tNDbJ5iSBfaH4nbeS8zcLbEDC3OX0BBqIQucmEu+bTbQZGotMBLRfXDXH2vRzJR9
b0TQvmvk6gd/qPhy1ShvPcTy3NNYdQR88qqR0cmvvcE/PtDtMMdEebFCr4Q47xAJ
MdhfUNzsA2rZ+fwjZMNl96DPpY5iROUTBIIP67CyjFdmZpbyA8nqM5e8TS240Jn1
SEeeFYJYnwQnr8BqGsjbf4qzdTWPGcR/v4MtpKpnJ21vpW3o+WrG35Bv7/xu6dm9
s2I/UeDVRYRgbees0KeEiWl+kWoT9GHAZxutaJF+jbZ20uai8YBahgaVBaQxYc+w
90pS7sJA6zroISVDXWg2FRkD45ofHDfc3eRSzma4ZHX3wFuSpn/VK+rbxP1t8iS6
bVtxKpyU3IEiuMtIlrRodqMRRWTR8ffHIx5m3EkncaD4N2Tk3AdISDvw+WbeYEvW
1YMgoffyHiwkVITaCDudY6wkz26AikZeqmvVEKw52xWD18Jv1W00ZqK2Mkj5rEaB
t3pi1UiIbjbqnYD2meM4ZVabIMfIBdrJVj9vofd2EcxikwT8/NqP+VMSUXAl3aWX
7ParFSB6TfCl5opR3wVnqXql2p5kS6pTqzjpCULok/ECh/OAIjcoja8MJvj3HImJ
0tZtSr75kqPkKaxBmFifjCUz4+tA93mdj9/gtUAz33NkRPqLvoIkmyhw7WDnvZ8E
rSTFVyRhPYqrs3VJ+3bxVGlW6ELU6OlDIhF1kcOhmD7npbhkMIUDlbkHsPWzt44k
4r4yXb3UGVXOqVEQ+4Gj+BQjXVdVmc8fPUzIroBHmno7vKy0rR+idH90pSThI5ww
ZWFRvnPdsMn7tigaEKezUqJCujPAi1B/74/OFcHgs+Rv6QOEVZbX0gffSuK1uJth
otzjMSovN9AAsQYcx28RgQ4vvt3hdxseJBYZDLnFcKLuKzFQWzNfogDhcKos+N1z
uW7fMdRYJEpO9b7zcElKTiTjSIGRADzxPplpiZRtUUPB7hAkkujj8847X6x1CfA7
L31JdAPkblb3qCrfBMBinUjSFgUW85knQFHF5WorhG8lNoMHPYsyqnFWwgG3Kr2S
jjg9AVI971FEDaasgcfT2RB5cjs7qoDlzhCdszEKgHbZXapwUJqJCUz8zHgD6p+U
GJj7ZX0mXcCn3diADhumRBg2MRjv+Pqv9l7MGXWxwGS4UAW5Pgua1G6O2Zctg2Gy
8GzLaGLxpEh6/T0U+/W6DKhI9BMhjKUtnqOXNjEyxIEvzyz5V1MqsilDXPnxAk97
nN3WW1EZtdnMXHdouCG1BqhzTQWhNM25ZS6AQaDAf9QDuApKWE8+pbvcVuVUQuLV
3B+jsWNn8IoYqc38jPOD7Gf+dvH8qiJOT6lcneNhA+QI1vCj3nUlDq65PJSVoZru
/A9O3DIeFiReBt9QTTrOiotjzASQQNnQpyLtMth+CDaEjWNdroB1WyTV5N2kfEkJ
OsGFb9B9DqvSIWGxdkJlsmnsL+Zr+LaPDnsrHda+EP3dQusERf/o89DrBhKgiOK0
JKwTvyl0mo9Lqrf1KL721goTESWHesCEjdNYPUDjJRI1ldGGEyqyW3zNNPHeCtGd
vXlbRSBLMKMzR8JKFNhQZOErZQRHJDRoUmhTOQbRo/Wf5E9RL1JbL1qJO4uJm37y
eAEbXSrhWn4rP4hoTVyMmMCdnh+uCyJP3Y0GWHJsN9lfBm/hvt1HbeSEmd+lZnCJ
ksXR0o2+7xC5bXXlhsNFWWM+4W0KLgCd5N6aZFWw49f4BkeTpz07cOCZn1I57VGq
Ortxtb22sNmIMu0kbbPpqZ5L9UdKOMWTrOdMQD+K42dxuSdvsezMWQQpooFVnL7C
jLrOeP2wkTfLfcfShrjJcOjbdk+3OiZiJSn1oiLktHuXspZc8D9OOCSXv+PVAmrL
fYB04LqjsPbpplB7NtI+SRCZBCeI/TE2t8ggdOtQEN3JhvFqXrg5213zFy7qEAiz
EuRejxb5fwt7UAgID9xMuZtn8JXwEawLCu6g3F71mZlaspmQXmo8FpOLs34H3pGR
ciUenHculYKr+MsHbzY8BiAGN6nf4WQJ2rNnEfCYKNtQN9xS642X4prv4oeIkNZl
OCB/4UjUL7nmW9uzAJAvV4LMY1Pi1P0B7iy16ytjtjWYAmhIeHIGSluit2GybJqF
kn4cifPc7EyzqLnYDQUDLrjNzsUF/2Ub7ywP0GKGlLtdxjZVluNN2cLQvyUhM0Zo
I3oZrSYX6T9Vt1WEIOeF4D7GQFSx6ibRN/5R/uexPPZ5oj0LD4ms/+Wasvnx2Qkq
6vtLxevWPmKgbFqLuhAsIsU6mm3OeJmHncnb5rKoxsqeQ9cKq7fOTKML2dNXeGaA
QsOlysY0vU/7ct0OCVFxuasjE+q37hiJXcvGCFCPx8uRVCt058IVXsl1Z0TxgXNl
eo/jxOj2Y14zmLWSo3+tHkdkHG9OOglXgjM/EWRtT3dEIZUf5QixXyFzHHirkq2W
gy66MKeQwELU/mox8rGMyzOgXfzcx0NhDPZycY0JyWMSvtMr8dQlOYq+/92+e/ar
RotbVHJtcMG4yCSuYHmXw+D8t4hNSNXAlrEiSnQcisixqKd/ErOtH3VzHHY65SRo
J57he2qq9Un8aJCNiXx1EXJkq7fp4tnuBqplbhCphFGOjzgBGSNcKE+IPdZE9a7D
o2+d6x3/xHzFHFHaVscmGRa+VVWBGTlWPVODNkMJYwt9ZkucLbJ/JUEkOPrd6zTd
8DeSSY4SmjYd59kfjW4KBppSZ13JUtQKR3OvheTKfs+RVqjoC4AYDyK3ehUsPkLH
pC7IZ1wuNDgWByaZRZ9r6Xfx8RLV/s/FFue7b2J8vkNgwce3PCTDrF25GdYLrJNE
aFJXkRXB1JTVYn9tNND627DxPRAdXyZR7+qZHKsF5zEkjglu9gwNKLSsYvBsInBV
j4btAxSdycpIjXPbPZymO7KYe+T69RLaTSXi0YbKy/mNCC6JpUJF0u4RzyIstMcR
91tRyqEoXTAIzUd8iji/XV02OnniebpMjNtwBXqRIQDulu5Yz7Y5HfTQ7JjsAu5a
kix4vnk2ZI2CRVkkkPVK8kjAa1mpo7RhkPT3LoO5KFETRYupuTug96tIxJQ/Exzk
Zf5rnNbDE5usR5uUSzRwesXWvLWrHVbSHwroeFRM+1ZGxpZeD1ZirKIaj4znHmc4
RhDNdk+Gff40TnuRxOQn/Yn9pGavgnohQH0cRvKNP44sS3a/Gb2wUSv1Adqf5gxO
B+jZ61lGCE68OCy1xdrLmGqWGa8W32IKMQ3H/Bx+dpcUZSeIis2GN6qPw3Qlw4/Q
Q3Qchj2tXdITrh4Mk+lhQOo2DMaS1eEFhShhxvVGFl4yxrjf7pZnIOrarksHaskm
vHp63EXjiiJk4d91nLF3yciJ6zqSTDJOR7dskjagN9k7dKlG6DjblRnxrmfExyVu
ml6zFBAZZowhjxhtbZn2q0Sn7cI8ujJIrCDJOQhjvm8nJUyCnPKq/BzkkN9CaLN9
YoZ8KeHNDY5ZK7uREBUOfTkbhaT0Ouf9hksqJKTxhykrK2PLd9g6jU8cSElbz+0Q
A2/kucaOvte405kmq4XxBoLcinmqXBG4MDDHIIb9wqMAflSvZgP3bI46f/AoFACn
+t8vH8VtE+pfsGCC6tma2j4fu+lwbV4fkIUByxdHjpccpL0wlFmOQF+bnYqzpyXH
vCqZhfDBibxYRH/FUZSuMU6DBDU/GpyVc0vqmLVJWM36mIe7qJiKXVa/qd3iiqvj
zCrq/kKuWldYkG78DfnMEqD+QJ7M9Uv+WhRcF4qRRRTmI4puGv5Co4x2qCC7EiNu
OVlR+hHoGxN0rY1ApmdYLQiu38Jbu79vbuDFn6j5rpfIv6kdlKA38GAbM7m8OLF6
SE3aTM5BtA8p/KWDkofWZgvWwZD7aVDiY7EObRb+PL/ZktDFdNoJiTsC40Xj64Tu
sPNP8X7gvYoc/45q3+CGX2E8ra5BtBWWUowAs0DHVsQm9UTnA7c0JGGVhxuJlWed
I6Z2DEpk9VqrAxg2HiqdKzJpbG5BX88KdU1ItpkdG1heUQfx08hpk3mfG8RLzI+C
2GzbQxVgPMsa/Z2oi03Zp9OGzb6dljBuLYW2aPNs5OVPdiY5HCbm4m4a0umLxJqS
it5SL47xGdhbGPRy3oxjsdh2+Y4mTvbfmV3hCZerlcYgjObB166RPLVwJl0oP7ii
FfQNZaAWWBnY3tnr435LDjycMZ6wQ+PqIGaDgxYoYxoLuvuG/oJvgUgTtmWBw0OM
LDgXibY08GNooPQKIpPxiPUiyZNhxDndD2sfTX4YGOqACzqUfNtda1g2UCRhFE3B
v2pr56N+nMUG0kFINo+I4EvU4yGT7czGxleuXylvugQdnCiOsFX+ciRK10AA4bS3
Bt26J+UGW6oRtiLqmMgaGF+McyxisSv9Ybe558QeIe3mcebzJmQZR4MRE26PzECt
31HTkKl8EQH0YDKh3rIxt/KjB1i5meOk8YW1/797YbwLi5+O712TT4huMEZHSGcf
7XfNaGj682sRs6ktXd2qOZiDij6aoKxwk3+nCIrncll9MZNyKfATEzfWPS1sf0Bh
Ah7YDI0j+q5lNzoxg57ty5AdjjLpOGb0ySKHQpUqAqfh8nHnbqyvtg2YlCArTViz
44/Qle5zMWohKTQnhY3C2p4Sc/XTNosNyurMrLeMkNJGifaE0UcOucg+Ihbc3Be5
9cbssCxXj9/8rQXUGSKlAQJQLA0RDjIbStus/VKGyHcg01D1PxVt09e/p9eOEfou
2eE1jYCW1m+nRHVWLaEVvSucYxpvJ0HHXh8jv7tLTb/PSXHtN/lfczmiQgyJemHM
2ASXPeRUkZ5AxboP/THg44TrH3pPh/o0Mc9YqeONYih0b3J+DtAXWUr0DXS+rABB
7WlHzEzry57EXHXjoWNGHiJ5zCkJVPI+hVpi3WCE7BJvxk8lybkuEGDEoYu+5Noj
khUxC1WmidmM+cNrRD03i2z9iJKIC1a8sbj6AoUE5k7bfhYTS/2ftxImuwQO3ya6
geE2DLpFSBUDetihZ4sMWrHKzv+LTS6EMPPDdOg8uL1qyPB0rvaAmHMJhwL45blh
b9i5oKuhEFoyEXUH8NK0lviv8JJfr7KaaDI/tOBGgSyX3XECmNQ1DMYkO8ONSTjY
gLrkTusgU4yr8B184TCgOCjRmiacDHTeG9m7+EiY0xuz+QTE5ccz3AGzD1ZVHYeK
KNSY8m2IbGoZYdyBg1PrDMgZ2/ERND+Ie4WtcbJ31pPFntBT1R8Wodotdmj1jMfY
NG1NXz1S7S828j84JO6fjURrOehqdksJeHyBTBf+m8lhk/34X7gUkl98sn+iW9Ut
g+yap00EsAWjtYDDGXza+leDfEeQOt473Gm1mV4ioH2zrEQ+Tjcq+7w/+dLUcSbn
U2NrT0p51SlAC5DprG8yBA+hsD1MvqARzHg5eDLB9s02ZZfcsk9FyZDOjXeaEQe8
IeTbmoSPkvRDJZSzvv+Yxxdo4oD4sxABv2xqIilzECua9N/sRjaBxDz00K4IMuyf
rCacW2C8lZ4sQIwbNANi4aIZ4tR9eiHkENmn9kzAbfbQqzJl9uhich7DGLH2Id3w
GEk4RE6qrWdeH1Z8fxcLDDRLnnODm9/DWU51CIko/+X5PBdNkF9CxA10FOkH3wZf
O3RakNkn4mVq72D2qfSp3sK/sKv5+c/Ul0VPQ7Tj+caIGUNJdo1C9dm71zkQUcjf
mzXn3uD+SC+zFj5J0s9aMIO3RMHErMFCFy8+dOPorNS17H31+auetkg4hQXALNxZ
ThgCDAG++3SeuQDSakV1/HvOcNwhjsFpQyZOBIF8N3WemESLGQ/6oCGDkCSEmEsM
OOsO53MVDz06rqV8ht7mFOzHAnG9ALsqYyt+lep8QQXoNK3oZFM93lOgjb7s3O4Z
TIpZZCrZpRReINI3cNZ70PY4cV2G1XT6QZ77FwT8YCaZpoLP//j/aFXfYPhGzqEp
w4kwDxycJhVRGGdwMwtAYKzOMGq26wEHQSLHZoSxFeUuxcQEgCh6Gt06A99bGXsZ
PHIFCgcHtfRLpWVthLdkn9bfL8DFI2+ql+WJqNCeTCyHVELMkJ/Qa69GNM0yDvQW
idcL6RQ0vkIa2Kj+n9qUycDOZEJty+WR0/yKx1083EKTnYBheDFwItB2N8JZEt3s
F8CGxdBs9lx7v4yM9EzwH9JqutbNZW3v8+/23119pUzwKNzCpzE+bU4Y+/B3EcXp
D6wA9lOBxAvzR0A+8PMAsOfPVXzxekdALDOcDkIn4iD/eaHv2SuqvwDwsbNyjyMf
4tMiaQztdze5XrXU1cly3LXi5VDPEX2EbirwL2AKKPnqxPDAHZZjwk5QYE34SmQF
3/2Yd5W4JNCS+P+1MI1FEZYtmVyzVgj5RNnqkCXgAGAtCuWHMuZkn1gmoyYIpHhy
6OKC1gyZp7Q02W6RL3A3ydmdxWWF6DbJpRF43kXKi0isqpnm7+etnmv+5elCp0zo
HyLqiOLQYu9eHpGIZg0wuABEznOCgDbkMJa0N01Uk7WvCdpeFmYzOtKsVB83t0GV
UeX1ks0CKzEizD2Q4QEBKTdaq8SHK9k/YAP76M8SsigjRReakXZDAkB8f3Uci8sy
2mw02OthsEYgGtA/gqGKWEAXx0ZdCRtiA+EdMAhX5bbP0viezF1mL1qm/mSccML2
XYGP6lcSZpItLcFWD961X9G94v/Zj6TVHlzNdiRIP3giGxxyC633orLQ2r+o06BV
/BGgg2T0MCy3yGbWtrMEv/3yQ/fq+B9y2lasLt7GjtdaN67e/56owhwG+WrU8EQc
I1l41z85XA6hMjMpk3bvOqG/kpiv9RhA1jdsyHoC0XzEjP8D8IbbCxw0JezMdFka
mEU8IiJtliNAtR07QL/6OsZrvPEvj4KrPI8cqVmo+c/ctxRs54YD8AqWoL5aoahL
wacLqU0J7dwoSc1u8E8jftMBRBhyWLM93WuworJLgIHATxAKt3C1RqYntbc0fpWk
JL0MEaSUj1s/zXb/StTUB37pUrelAtbs2snet0ywPXADueoiyNs3JrpLFnBSjbSJ
MnYV2CPx1biogsQsiLFkTptm6GQ1M7WTk/C6bl+Bd0QfQXRpdT7/CQDuJCGYXcpv
7PQXSw+PDep8A24zp8VPd56TdesA+4ZyTGtSmeesUsN6T+doNdDRb6DCuE/XMsk4
wva6NfeuTxR9YDbvluM/f0ufVlQr+E6dwQunxadVUnf/W+iADUXqdMiHChhfP9vu
N6v9/V0umGdiPqULGXu2Reot0xgeHOlxjiw+aZThRvXNyxbPJi4sh2NC+RMk7w+W
daivfpRvqBfBi9LU6TiS1rglphziUZH3QnelDo5nGxYMI5zo9da53aV7oNNlrh7f
oOYfQ2jXkEOqoTbNg3IBed4OuYuaS+zP0xV/5QQHeeazJhsGKdcbtJX7B+pE4DaR
cMxjvbPiwqiysKjtOTvumTeIinoYoBQbYe0xN8MB0O1sjp1PKFNw2Jt+kXyQXbUk
NQteOSDLEjq9sIT4Nur3CIzfoJKt3H6lALH5yy4NtEaxoO82bvl+eGed0m6WxbKt
KvGDqtEQnw06cFcssOE7u7nuHcVGOT67bADua6s6f2V0AUWxaAQh+w5jGjtdMivA
CpFjXI8fJgR+aWRb7SCq1fmFmFIXBeI8C2iZ5p/m+AqvD+Bo/zqAohQTW0l8JGgn
A9azzYlOwvSysg1i/5xf4I1eOpkQEV2EPpOEkLkHTgsVr1DQ1nQb2aV5XE+ZSzUD
XgG01M7dIiSsomdszxuiFlypk/GISqxEqXUdbBhGLEsX+RIxESAv4gWwCu+wqJAT
O7xXeVr8IArM7EvpXuW9ArUBlSbrplynJvyB6G+zsb3u1Jc4Mes4h+rGVg1hRL85
e4UXMjbWjqWa76VkOibg4fbTgQxkCM/5AjIfTBXqsSzoJHSh8npblOnYqkuv1PG5
vGWzU2YaUKSFdDQquwQMMOMT6UfGUoNksT6n9yoZNtomPyvTR0gf2xdRRS4zpjeh
VJkQHVIKkQiehbso6+f60sbCblFdj4/1/oCtyQZ+nW7CngN8yLOKoc8h1PHBPQGm
yc1B02SK8ZOIFBCKyG5zgG+kEGTBhqdlobksPnZpF4W5DsmwBYqBhaB+9cvN/4fX
1+tPcPG1KS5O0ZEf35VU/enQ1wo+ZFseYwQMrveZUmJjNOIB62M8iZhXL6AoewD6
idDwRBy4AtCD6VRxgNXpAuxogotsLzSRMk4nXuzxtCQhTk4tm9zHec9Mw+WobA/f
Pr8eic3yOu3ONNdfvw0G4h9K08G2dJYpVBYMPj5uBADPC/Lp/ZjA+5uMRlihiamX
d9D1aConbOv6e0zCtmxJX0s/ASshlGlq1yfaaAPriq1NdYKW56lu2RlwyXxZcVIX
WHNh7sbtTvrPhITegYr1CfLhEgoBOC0BajGAuy/IO1yAwie+IoFgUEbrzd3MqoW4
wX4Pq+mWUeRnrHRCHk+16nBnL+Kd5Db7w7ddDJ1dUvg1l8wOSuWduKv/rNelKteU
SQ04zY2QCpw4tT5Pr2UwBLYKn1UiI0jzMD9tlrJvqFMk3Y39m4C7faEl4oqAozS9
Dwtv05eriCl1vWisFZ+g5Frm6WaJIQHu6BY29T5LY4ApRn4RNvbVchw4nJWfbVuF
2QmA7iOwECh6hVUAWOAsoGX3H0TMFPPS1bGrq1UyP1rba6qbPHLHjEaNSG+up2AF
BCL4Jg+ArZCb4/4d2NOOJr3mWsKUGWNDe5o9+LFy5Wqe9++a97Wpt1gKtJpxjDZo
Py707Jxhxx5/5NwtfQuqHeXOHx1qYkWOjJLIyEqtmPmjCmDAb2APTtdOi4veJswm
tR9ahUasKt6bXh3zHnTcC8pRlEWQH5840J432DLHCAC8prkeqr50SxgtCpYExoND
3riyu6w/xifN6yFHxH/NlFTt+dWsmaMuvK1gl/SJGqcAcMFA+gvYfdouRR0IZSXk
Dz2/n0GP2c4F2fbUu623IeY6QlO6CakleRJ5VWivmRGia7Bc2AtEjwzbQRan9UZL
CkjLlT52wOg9E78PPxzm5T34FXFs8hc8vL19E6OnYRi2cmIsvX6hpMNWD7o7dJlt
2+MQTQkiE7ToVH1m27Ox/J82DoiQ1pR4IgGkDh+zBC6fn+IyA6VPvsAK6JIVP9YN
PqOo+c9mk8gp/RSx4eGipsKsoX9lHbIkEw2Nga6HXwXW+siAWh9qkG3idqec6XHV
FkszlbdKEPNMNozqFoyQX7Wti4mfXjtlIQCfj59N3iOSFSeZi/BIvg/ZD8PyeHBR
CfoIPwRnr+TLcGm3M9R7W/GBHl7cN2mAxEQnBdoUnv4P5tfIqlhkJ41+rLrdCOUC
1Kq2PH8bshH+P9aMPHf26jdQAdhZkcTu3Fbvl867qiaU+rW5ufS6cPMirJurVI8w
zs8pqVFKVkIbB6dYrReLXji8mGCUsWyIyeRtkTthXRnyz7Dm0WewsH1CLd4oWTuj
iIOeoVRFAbqwRt26leE0cdI5NWmD8w18jT4Q2p6LwTh7oHmYDAqtxOA+sxEB3Ug/
9SKnclVHKcPZBuVtEHyDdUlntbnJaeryOgXwNGs1ixgW8gIxHd9mAcjjCIojJDjL
WEZWlweTQZvvG5uqZMjDdBmwTKMTCl3XhdOu5ouoIOn05DO2s2VgUlSGr1fZNl/d
aJCqnQMFaaF5Lgnf486/EUAWytPWm27MOHAZJwZ20F/jEE7C8dj2f3UdR1D6s0Vl
EEz1VxOEHs3pWVb1ivSqbQUiCvaCPEvcnucxHzujoYFFE/IAeguuO40R2aqP1OqG
SiGSIASy2R6YaMfi5qoSmWkKXNeYANgRBSiGxxN6l6KkdRkNLxZRk5JHvMwsW6k+
+eF5QnMy8t4mtF/CfpuSEj4GxERVrb/L+Au1PbJZAhVkTzdyZJszO20CXKGJgoKy
yk/KkRsHmTReLamEcWnPjYoEi8xdaoPfphNNF7nsJMkO6vROxLDxC/jzMaw2/W4q
+Kmr/DVeReWsjsXgn3G00EGYk6TWj9H3R+a0guvD61MMkkv636xJWpFNvcDUG1Lg
M/jUwvZiy073BcMBhbNI8XhbM10uA4/yJwy0HmjUH0/BSFphoiGYtLJ1xHnlJK7B
TI0Css3McZGjW0AfAKNpCJceOf5mj7TNJG763q4fHHBWd6CRX1idh6GBOjc/ezCG
BnNMtFTwN7/3wKCZkkqVugfqsOwuK8PJy2sW7YIJAIqRMIiTa+yv3yyiGXZ26eOB
XLiA8vXQ9xPiuKkC15QmDLUKQ27pH71+kXYwwrbO+KYun1V4omzKm2DRvSH/13kS
M0lTpNVtUkCuzCiUOejC1LmlNBV4aM14U1XBRukDPPwTZRKBEpDsS0OLuo7Fmmx6
KENz9K32eSF5UC96lfby4H24GFpfHiufVeNtjRcSYn+Q+7JjakrhjC0LWMQT3MR+
wHdjvNQcwu9wfFM6rcYELXvZtqHtUHXnCCO1VxZlMKpjk+qqCtg3qnKhHvtPumTa
Fv5NA7JHmeBEKMk+CTNjsJ7iPTEeyuxX6eK0dDDYR1fkQpxrCmGMzg5fwt7aChP0
sVaagqIoBzcjpG6frTJ3fZ2+vwGJXnT9vpFSX2a1YRr8pERXpGl1glYir2AEMgiz
kREz1LWWjr92meMYhFr+OcXBAXT85h35OVrZnd5h4cnqDI6NDFnauOUuyl/s0W+/
kMynlZPIagqv1dJsCdBZAlk5pQ+GZSXmwSrKb8M7Q3Dt0nJT5Sq/0cImwTM8uw93
HVV24M4L5NGcBUbRGcOrSjZCOAzMext98VSJFk2Kj0QUxq1wZYe6GBgiGlHiDGRx
noGJh2nGv0JZYsvb75PEUBhYqMvGh5hihVqsI0J/K4WdJdc0+g4dXBOi43Svqvt9
45SOUOqkvL8CsS74Yj/hzpdwEMycYqYNEbsneZExW71FbPzcoorOY8cswYEfX2JG
iFE5VP8edp2ebMtH32cE7F/aZqR1JT+OBmUG0pX3APApas91ttKDe9mX/PcLn9QE
kktAbScqbbvxHbVytauwjJmkwgCTtE/roiYh/HFGbw8UgG4G5yjVOAytR6QXp/Ko
gwQBqQA/tBY0r73VS4X1RvuOVEWqx+km2MimYLU8+p2pul5BFGyo/EBSzhEjhmXu
VneaTGFakRt4aBlJl/9rLkUMWXRrOoqHE0jkOl3JL4iGNDQpMg/1+XdOpFlEiOve
Pefp84yWtAPCFmdkRg4pOKM6GCEQli0GlWh8Nh3u3J94PkYyfm1C3GWvjFSGUR8E
F6DqJm3iVhMU6lxWghKxAruwtBTNTPii0Hd5GB7teZquhm16FZdbg+bPkheX//cG
iUN/9gpoDPylVIxlRj1w4cg54fw+rk/kVEECnin5iLS5TKyGnRFTClJAJjtDk9r4
ihhm1lhFAG+L8LXMUSq7FBqcZGKUq19utpJje4Mop6XlxED24OwX+hFTrRY2fPvK
Z9CXVLzzS0Ah7bD10OAF1SXlcpaXIifBCeehgbW/1Hs2qDfPNPeI2FehRlAJSg9J
5wm7XA/1hdsLF8cOg/H4GxbPodggGz3D26MfJrNZTWwm8VSDqi6TQBZ2jbzb3xAQ
IDHRVEphJH/DR676QeInS+4N2ZRxkwe/Dof8nOKyVusKWjZaFs3L+yfVfA69B47H
Uh31p+eidg1SgBmlKCWuuATTBUV88UeEtRBNH/oUVvDbrXL2Tzbn4TVZbo2pWUI8
epUROUq67UXML1xinQRxNcLS5dbSCzlsqPs50SIOLbd6f5kGaJAc9JyxkBwymar/
7axEFJANL2BUL3fFo/aDfi4wwCMnKM8bJ8iCbka0t8IlFGN8XL/ruODe60x8hL/Q
h4M/pZGpmPfEa03cbexxzo9a58BQ+gB+TuBTxfMtIiSsC/8UDXb04Dbb6MJnDseI
E7xPRjMhWvNl+B7GK7CkN6GFSDBieeVJzVqpvVhcpaxXGDvYPHwVgltGKpnmHdGx
wqSKMHRJtzr7Z7QIfHlSH82BUV5R89Flh7qTJUV7JDeAp50s1o78G7x09FHqoC+l
sj/FLDu4GSgHE3yZB5s0T/RP3TBxkqsKClw3A2EvHRQ88i4FwnziZ8AwmKbHVY9Y
eeh76K9Pi9/IOxiZ/hMCwLE2biENPEhpmPeqg9ctgl6iTZAzusvmeK5cl34wGmAs
3nods/SwJyQzytVga/IbsfQKtrbLAbwUi9vrqOXbtoije0lAaJ/m7BFS73PblE+W
AQjM5HEzwQQ6WpYyM/ps2Gik/0tfapXBY7ia21DyohTfcj7K3lRJMA7C8Du5kD02
hW0vjGqAnVl7/H/LCL1aFw47Aajj8kxL9k6ghUzEh+VxFlN7Jd1fjlzqHpx2OwJW
ByXhiuDSpkdZA96FgNWCjY6bH8vW43Oez6VV4Wr2j2KYyY6HgciYIZCgr6Ew262I
lMb3EMiWZtljHbZP/vG38HJjkDpGMa4BP6M9tW8I9pFEqdMfII/DSetNh1ymAnT6
mJ2jgmD1AePHUbQubrMAi3Nq5dilqGRiCTJ2NGHSjW4OMtpHHxyufHuEhLDr1N6I
p4FzsPKdRc3LngdXKJywiq5jdIj5iPd6/4Uu5yt6Xceex4TS8LgMZqBzUwe0EV7m
DzA3z0vsVeSS5NfqdBA8GzyOlzMvEZazJNfMPPQ6dqT0B/upbWMlapofg0DCLOQL
VXxoGeU/xhNpEj5njxhe4q1326LdpbC72fLt8LjcUqbWISoySXXvAdG6GgvCw97T
MhNIZuk3EKmUtWSCMCSHhV6Q2A0rtMUTbM8sZCYAsFMhRIS17t5VIzx8aokPsB49
q39ycQ6gsNNeUErZ5zLBbcu3TtGtBKSaVVfMZAa+iWYilwxLYsVQjR1GMEynYF7v
E22RHiqYhJF6E1kTHidasYa1e9KJgS94/HURI5Bpf5r38rE8cfKEZLVmPCG7szTz
PwHpI91MSV0KFhSWBmNzmVlFJ5E64yicEKTsIJ0TFT6MVNswUZb9/jEoPrZCUQoU
7tvvBSxK3aSZhIzk1K5tepeqMrLqUWPSNmJvq84AReE1Xh1Mu2HTmv0mnZxJZW7C
SpRH2dS5mbqaVth32aNhRFgf93k1OiIAwT3WIZ3z0kWcl4lAGIYbwXcuE0A39KoI
ORliIEawKX5TkJfL65recWvFS0JsmWLOh9ImWSCap0EHEIb2iWcBsapXzCiQnn8m
RZ2k7JNTd6ZhCiO1Hmon3Z1HxZVwirp2DzPFMvc00YFl01KUjVPShykpP+NDhzUg
+MiII49vX1pk+CnpVEMTTuqTIlOfJ95GK30Vbah2ci7z+/2g7cSr3Utbr/KzqvI8
Wh0I5MHzGzonBlK+w5UfAj7otce85C3YdMZQ1kwVEFJIER/XoQIyFO/MC3xyLLiv
UB2u4eznp+YSW7HT94hOoZ9vG747o7MDUW0dzDGbsR2yBAYK00MuWX0ZFZf31/8x
Jd3YTGZ99JYs7eHQjRcnPwVSd+7F3LkOyv0Av/dmqZLa0QM3k4HBfITr0NSc8Q99
wbxJ1G/5Fy+yd/J7GM1Ex1t2n6Ll6zp6yjuMLF8YybtJRbVN7UsKVyjn0dgZFIvo
tl2/obq1MBc0FwCFvjrtM2kpDf9KRFhIDr5QBQB1LpMED+z3353VoiUidaXUb6Ea
7+VEXhnHDTCXUmjQ+xdUCm4r9ZVTOBc6A5sd2tffkfKRjlpXiEAHMvLpSfmR1Vqi
qY6B2yGaXOT8CaLPZpyGPqUxm7426+oWu7XHog2J6hGTN9QnfxCJQ+Zm5fqbzgig
N2FefxJLeUiw8gWd//TNamojYPaI+RiY6y2fLRC1unGp9K94d/wLBPxDJXHY0Aip
IX9oju3uuuNApIoGx/RNppUHudXmxMk9FChxpa/n5z52ngrYdUww+o7NAuq6twMm
v2PiaSAaedQutEyufZJFKY0NMD/xcc7QMIUWSgMXxzhH7HeCtj/sy4DL/PPTPNHp
aDiEOtDrDIxREQs77+Vb6Subc7Wp+B3alUUF0kkEsCvYOxyWl7Auk7O7+9YHC3p0
LWMLqtUAmrzTXSwIzuq+9tIgaGh+Mq+O5YJMBw1NXoqk7fa0HYNTgr2BS3JQVmOH
pbLaTv5Kz8WbVTZZSK2jHdYxVNZmYL6RDKTM5JXtlZqrAyfZo3Pu/wVz9r0CBvV+
XDMkNYdW81gb9qTYFmbY4fEZnfDV6cT2bIPLmMpzKNzMAAa6oeSBLRzgj57em2VH
nymJkeHpBqOU7OE3qeDdLc3hQil1cpckm2loolngfVuXz8UjvzqJqT66iDM1/IsD
iTmbK1byDrQL4eHgHW7ntdyRfW1gD8sD78SJzz0S7l1Q0xP8o1FU0z1x0/knuMCD
Y2jQitVEnahNmYwtH1Won7nYgxINXi3lX0J2NnzYvjqVyg7Se0TKw1EtQIBQt7jI
VyuB7vtRE1XV7hf41y+9JbS+iy9f6gptFAo29sQ5/BQsi68GY+Y+kNDnP5NihrO2
0uVWdeNQsNoNTdl5vNbTEdPuGbySDtEZ3AmYPWVt6atLS6Pl1M2I+8idvI2Dk4n5
4KEOVQ57CH4y1MfpUu9odY/VVwmmLfapzpfPI6+oW7M+GVLGgzhnF065cKZu4dUS
KRN5omB5G+6xfbmis2uwDUFQGJ0DFC6of8O6Wzq+4G+DE2GYnH+ZsciFvezezZBc
zB8o6/AmddZ19CQUE/VTjbILpGAqf7KKmAy9jO8HKZUpFIpIA4L3opNHIPpeIkms
x9755g87U7l8EWuv2JCF8ke3sTNJ/B52iAIRWBt51qouIycVNp/2C5bg9wYMPIU7
RvaCLU6vsyNFssltOGLYebUc+pVLcaDVFFqFaZqlnFvU/KFFNSQ2wyhoze51nV4K
RS9nTkfIaKW6Imb1UktiZd1MSgOYWpESn3kQ7BBdDDnkOFYA0LdpsDbJ7M+5bTKI
z2sF+zUjvM8I1UrhyRlgfafSQ6YPey9IcJTGu8Z1Zy0s7/YfUoWsh5hvgsz0DMqW
QPRQ2wKRzMroW9CBKoOlD5Sp4FJ7gBcA1A+/Z/IzbkP3qrzhgsxRtcAZ9hiEu0sz
0UWuSoN8oHs/56+9KBxh+s0HxEdpE0fF6sd9dAC0V91nxl/PGRp3dgX9Zsd6sgG9
Yos6bK0S7HU6Vr/OkUAyoLI9D2V6g3xuVxCdDRa23VHGpFWEETa/apRlAXefINho
EFRDWCQ1kkQGJitkuB4pHjUqToeJfJTT7+8UMycVKXBrIsgi/O91p4/18lUaP5Q5
xgWr2VpPL6SFac/cyUvAEQswsUofo5G7T8cfPSif88VCG4f0TIDPM6r/38sR1TF1
b8v579GsfOmne58clo8j2ju9AQAykfooc6kgNafGWCYdOm7PgbKqImiuJi0RHcMd
EIAC1OgkNh9R6pQYGaMu3/1rCPF8mjAeKmsHrjnMTqsY4qldRgJuCRr88PrAW2yV
2aCrL+FoFmShvK/fTI2GICHkPNHweIWudf+uZFdGmaUk+msxhsKwfzbulraMhJz9
11pbNG/Bzg1VcwqksWDrKcwM8ZAJRrI5mvX12SZ5N6dHF2sqHXvxsQWafeWzihDu
kDi7J28vji3b5Xp/X+QFGKXbqlaV24/Aw4nu2aKUbG3xFpPCGfIS1ZBwQo+Cx9T3
tl2AXkDCdgKoWhVEHmkbnciaPYdJgci6Ezkw3KEvMw+rqVaNLhcPdrFBYAFSNdTk
JTmfrmjd7J+nUvvtat7NcztvWpqIJ599r9xiJEOECC71RUWKoIPYX6784lv4nUgd
z0aR0TuBkObIEcidpwaqHSVshdo/Tt68Pxu29mqBGegl3SusuRF6hwAQlT3YeZi4
BNcWrM/PLxOajOodAxZ8yav6D2XEIciJmpTUmSFuZidWTiloQrxaMWh5nZe7Mgch
eDDf3lNHaymKk7NmLNxVnE0eI/B87d0nHPkpEgU7cikj3OVlw+ucOsjO0tFFjoFs
8jRFLfeyCzqlEjJiQ4PFUWBFqpZqO+H1q3q2CJBzreH3bbkAvcm4DQxYBJnQnhtL
ulI5uZCh2GF+EqpSnIZGnzLgIrqoMTHXLyUOuvHS6fLCLwJWuUQL5BWIFjIN1b7a
3I58ZOJ/pheFKeBlHSRkdF/t164eTvRYy3BngVfB6WRxvNfTaNvFwaKbPrV3/9Ua
IYiEIBkNRbD9Z0Ux/l7MCp/ff3gHlPct/nFpwNCUx9QHh5FFJooKjEeObdblBWBP
imCXsevhRFW3JuNqsDqUGp/licZSJJ5pYls5ki5aY/TwtEhraqiv2hSGYu7fCt2k
XgGbpgX28tmKfnNItKaCo9FEFcQShQ1akY0P3559qZp0O5LfiyTm6G1e0NMlA7Sb
MhPqiGbP+HUx38Rfo1quci5/7/VtP6TEfmE0U9KbnlI7GrGImewnpOJdibE7ZTJD
d9Si6gLPESKgJApy1agErxxuZyyK1B8FuHKKWF2goZRFO/ZlWImANfdQ3wD+XBwl
FRppT0PGd8/JG82L+x05dgi1Bm6wNK1OL0QfhNnUEC0J/iz6/mxVhAHrXiG6zT/W
TGaz85O1cx7OveFN1Tf7vsIfaU3UUcwm8c/KbWOycNo1QsXBAcL2AX4XpGajygNQ
uRh+ex5KYpXOb/tkVPJAlXpy8qzSy5xcVPCk9vVzlZ8BDAIdKVwkmhyYVDqMFgKt
vxAi/hfZIZDJIiWml8Z6oGDvaakZLGK7Nh2CWJkyGdSPiwgX+HWKgiQEK/ZJrB/N
TvNdeifPJyeYhpexOm2oa2rGEUzAokTGfd594bKjpq/gB2HRZ39vGYDUHp5duvyh
njLBQenctkLyZvUtYmvcIOl6w8KZImm+wGiHEWRdNSnz7pl/rdICED+hWiuEQuoX
GWFTC+BQscb368O0SrF9G1/8QCmReajlaQ90H1IZKvbL8norGrTXFqqYqmV5qipe
EUOdRKxreRTDVNjnpHOreCS90D74CNE+dZgNXwecPUQ6Yf2Pt0/ZuvkcbutyWIqW
2sGjrIB9YA9E9AiKsLsz1zmskf7SHJna6NK89D57XAkuD8jMMO151RTjtNaf3yvD
N2xZmp5QdJtX3n13TXvMKq5+SCNHRrz3uNZMhdgsWe8fklWaR//6VVZy+IJoNUJM
nqhptbB0XvnJBQ0X4P+1tErsFOYtl/mCv/uqWX0ckn5n7nx2/ir9pvmy5Sp4o7/3
Adg8/vq7v0mTYZYvDClJNPPWfZ8PSSLp4N+gjeYwlHn0rucwMxXy0PVz94SY2eMF
hFQH9zhM/dmMUIdRbXxGMh21xV4HCXdfh+HTYoje2AHVdjyBLY+zZL2NbdnWHUyp
mL3AUEntZrH3y5CYLt9+MpKNmUdzWvA0QYMUFzTnri52KSLEhCKpTNr3v9PEJO6T
biEAXky2IgA7Tcwkeb2P5BPvjjVguF3B3szYdA60Fyj4Fl3Er8BNEMRw8aRwA6pl
rOdxMlaBvbt1LiqCzLZ20xJm7lCQkj69qxSo3LqEKIR5emiOoHa/31PnY3/kmzM3
yZeT8J9A68x/hDiNrSC0QXPhU+B1hk0gnzLa643WIOvnlpADd1uIr0wDstLNClux
EZIA9torEnYgynEqTeICApLnLWK/oKLgmI50IbSYTuEFG7BGaTl5erChWcv1EfpT
hRKpZ6yR1i8jd/nX2RfFkQHJu2mXvDZSKHPdV8dAyaznMqrNfEFYaNJ2afzhvGnZ
fd4CUM20w2Im4pg95Qm3VqiWUTsCBK8WDRVHA9CJjzFkmfQ1iqFAJU2wzOcZLZzn
naBA/GyWrhsshrIR0gKbW4POiQG1/Ofy7G/w9Rj1gjH8f8chbtpc4j1fnzLKaQeF
svcdW4XDC7sNzY/+YVBeZ5kWQvAb8MS2zkKAbCX//x0mcJyn1cHuM3kI3agxhiH1
zeA133UC3y8+zJsZMsbU5v7r4w5yEMQeQUAqP9agdaJ1ptyLYCvZVCsN7DMl/Qvn
luLcma2H1lW4ouOu9muf8g861n5WB7mE8Ot6PBktkA95CVBnAXYKmJppnhptfuI4
S+nRmKInGPfd0Z2OjPtIeaqjra2tG8lrZMHrd88GNaQ9q7r0kxU+cviWMg6n83Hp
0/xmaznYkK97wjHFqYspoR5OqnuDqsvGrEN2L1yXHiTeCLD2fpZXJu2YRDOhuG8S
IBfUwU9pBQknEU5owmz5PAj6Dz9zyLP8Cae63vQmTouV6QVOYiEmnRifh43RJ8jy
+ShEfdOvkAi0OjPpFgrohVGurvGL1OWGdQTldQ1+v+o33dj14fnJzYjEvzOm6PjY
pXJitJEPzPOd0sLBxzhRjCvl56XnQ+pfxpyufNJ4CrIWPICbT88Nw+i7x3pblukF
krmXtmksYX72Ti2O8WNh34r9KgpidDKRJMenQQ4lnQlz7I/GRqKLfdwqK7U0RH3H
xzgpEGzaMGSQqXJPPIIGAZXlLop7Wljpb6QBJfsR5e5U0jBKf/znWggRgqRyqrPX
0ii3gQwrGkWwAV5TwM9bAA8v0EOX1q37LSQ9IUrsSUcuS/e11NCeMMrsqcw1UzTY
nTVxClFlwggYyK3MGq6SFYcnHStfHF2zQYpvwDeh6U6CjgwEKpAkeR+1zoRyoeyK
ud34+Oe3Trkz1pLBgki+n7ei/0YfpCV1ExxxO8Dy14Zi3+AXzXsINYy852q6yx1+
Bcnk73CpDjt/CV1rzIGd0nhpBfk4lmLKYm0TlUjrNsxp5LezbnCJcMkV8MfacCEp
k5xr3GqVyhJM1jK3bZJ/k9OMlfmn44w5xbIVgG5UZN/T+YV/6mHtoAwVa3UNR8Y4
7579fk95T2/mf0vdszfWazSMh9LkY1242TRWAvvepZG2trcdaSTqquqOAEd819Lv
qp0f3L41ulweuO95aKo8K/dvRiUaOvZOUP6tKJ0fs0xOhRs/8xjXSxSYlSjBvRFR
PHhjOtD180bFrzXsaTuy2adPifTHLUU459LiBosscc1Ng8lomHDiGGRj+QV9wAP6
GuR6wHoMM6r8+6zwDzADgl958/MDWS3LJgibYQmgXV0Dbhjh2AzKOsLU2/6z1yat
b2dnhioyQWjN6PDx4MQnm3IqaG6kJ/gs+tfwLwJByccj/uNvoxiLqXRlVGSUr3kG
Ub0P2SQppSiT0mgHUfiEEdoFWraglblfKGT1EwIDOECfdseKFVWQ6gzitcKm0Oyp
oXJiumCat+VHFyAyR9c7f9BleyDC2mvHc8Ls7IntVnbLI8KzbXAnDa2DooEr2UAa
1VAIN3Gfhx8B+CzoNmUvqe5kvgGKb1T3g2k6d/ld8VoWDL0nQuiayFpkmLmEDW88
xJHAmxttn4r19pNShiQviiw/okggKQ1mGJb8JI1i/CK7Em/zePEIT/2vjE9wQSgQ
0DREp/ADBdXZRgfDDAAYPQGuRu7BNwqdBPI4NSuzaewyY3uWOWp13C3dtyVxMDBa
7xdJQzQnYpcw9yXs5ZWLW0OVH2SKlZ4/VC1bWv6LXVxjz605lI98K5jqtrZ8ncXR
oUvmRmFUgNzgrjQh2YGXNhUn/aNRv4M1WAh3ZVLo7gBMFXSnoril0mTe06Dbavs8
KDIT56w5WxCiWZ01f7h9KOIQOcxFA/xpyEXK06FBUjfhwh2Ry7OGVM4EmbqyT0Ni
RWVTngLsHzgebyXsFvr7gx0hmWmGAP2q32BOM62kuxU3Hik7ZcB5i/Z8g2xR36gN
Z5tcu/QCrsWL2LGoESNKcd9tvCC/Fy8aaIuXbhL26IFSr/wlg2NS6KjjRy3APzZR
TolLytUPiNn6CaKa/Jrt0j9Lhj1qu4iyGrg51i0BiDecd44N1pAL3rNstSb6CWbc
IObA4j5B697GVlqyUqTZCJpPqm+o7pb+bw/Z0jbZv0rVFHuNJ4fSTv2B6dv2CedJ
1JwSOAMNBiJiPrHgU3GVcBEiGcH17BUL8/jkyhi623MPvY69FceG5TpHGUw7lxYO
tPXmScsQXZFF8Z3wZsLQJWgHr+g2+gsSQEvvKXNVKN2YClJ+TxY7LPQA3aSDybTZ
CRH/3WTANozw0NKrINlXPcGV3OX3OdsZ/JQrGgIphBcE7Y9gwITlCffxDxqjmheV
lM0SzfPok3gTlcTQr0uKdmOl1sw5e5E7Zaa2KvYKiRjA+6hWvGP17QA5f/NaKJZ4
JSQY/zRQHLRWngzoiQ/jkrs90/Ws6oTVcRIyXsMtKgIYwBpYe+idghIUMM8OxUFG
LO8rbT96KttRBR5aNM0THst0BGoA7XOu9jUux8JqyM1tQAhpf3TGRay8KnM2BlYw
2KyqVD35poi5N3Va+YnfqN4LT2pkjnr5FPo09XqUNEtHQA5lRPedZwwr5Cv2NFz7
cY6snSaB7UL8UXhsaT3XMGp6z+DDUBamYIgMvpS8N9iXb2LeyLf8bJGNzvWN6ywF
dkjOTrsvUnrgUxcwC3+yk+HqLcVk+5rYxN7BeTXywOcuIidbeML8wlGXLwySsEie
FwAIOFvRaVJ+IDIABMoIb53jzWwY3gU7COATG1lPEQ4z2wJ1jhTQM5w57I/5MQE4
Ur5LzpzkOUGfshnN2pKomx9UEjhaNkUSePh/cHrR0AG4dxfdOsEhpm6XszZM80k8
AGNi+VNdQ13bGrr++BnNoHJuC+aHBXArTEkIhMim5YH+R9KiUzkjPkcssd+UJ8pP
Jo02fjEGFk2p+dbPYT+tpdqfLTCcG9yRMVPMgjRpWi/sbGaS7TxlkIrtx1E7j9J9
di7oIJTl/7nFNikMasDbnewFo8ffHHXs4SK0JnKwB2/4LgDpvvitG5r4JuibrvJq
NhStOoAOMWxVCl6acsldIBqHVMdh1aSV42fxA7lUAMWbDdCKRTs0HEPogxT16OI0
LC+4c0UXc1lq0WT+WXvnGSRXvgOTuXbZhRIwhgUYv2j2GGqPbun7IsyDTleEwpba
MY8oqDnyS6AMCMAtQWAPGon3wT9KYGzRTToiJUNGySeHqTSUhkVuJf1NBSRlBZ5x
3YLMjYAzP1OU6pdI8l4QNsmcuvzto8lMsw0O5sTNGXK3rdVLfn95c7Se0wwjT1Z8
yrdgjg4iubUyTK7XxV4bfB1vG4Djt9nscDiWm4/Mn7MHvECnttWYZFAwHICk5FP6
2TcGq4809CUJ16ViILn75sOfHXhPpiZlB12sFE4oW0kqt34IsRy8mj/q3JzlUQHS
OARrrOJ85K/Wa0/bATnL0RKGStATNPFDRX8tvrjadvooO5n6ZW31Uwt5iXjf49dp
DHIXWd0Bew5SfrjXaziwhrBqyG9QRGan/VAUOGPBxIjp+2gVFLc+CsONKl1J4aKO
lsikfNtbQLjNtkGx+4Av7gITH0Klc5sPMP6pADf1QdBH+kcT7fTGxxzpJHK8g4gs
XhsLE62NpudcTtZ3xOHnxM+Agiqw3X6G+Dig2xLsFhTfrto/eV3cpzxW2kG6QODY
AjSyZzM5xU/PG9LrV1huQL8wAYE3zeP/nfi2L85CYEj2qCfvvkLcOlVEY26bxv5g
dIGVM09ve/mnwPNKphT/nXyMYuy+XVMUcoCGAaQE5UuWZaMEit7wxunlMVRl8sCi
/eMOwMcvWvhVuWQChmgFjdPS66IG2wJTM15xQWoWG70bTSeRVv9IdehqoC2PLKEF
pMtWTRiGhNZrUeyzp2Z0JOUo/iLtHj76qO28YQMhpwNCYFAxh8OAiKbg9vo61IM2
xEtRRWszApYVizahdF/y4k8AOiM/nkmtYSmnPRezAujV05ZN/TA00m42iyI55gJ7
Ei38mSoNAbrel7C4eZBk6ca4Rf/IcN2A4hAm4D5HM3rbNxnldNXc1PVhwWRj7utv
G79BBjY8zl8oncT4z6ABP3Bb+A0Gk5J2JCAhTGWQmD2eN8zMiqTywcDYFUlkBqzL
rFMp9xrQi/AcfmWUsScsxRuuTY4DieriR/dBosRa3drDnBqahF4o0vgf8KDii8pA
Xzce2IQnqGNnSbpYlClRyAVokIZ+nwng/OMKdmFNkoU7RpvmP/ijE/vpUzhwpEtw
oBiHnxZJ0tXrL8ElYT4gT8cL83Kpm1AJRnY5WKKg7JBDi2XUrr117fPzO38AKoP9
H+iRK2pmAX0Ch3s54K7BquZHy2nV0U7477HbV4rYI7KiRPOVpjphVc0i/5H9I4xQ
ie0M6wZmfsxN6UF8/rLPGiC5eU/aod1bf6vOaUrSoJAQyrUgerCnLcV3MvxJXuwG
Q27wnTpZX6xgj5Cv2vzPsvZMCqgxV/mPQtB5Di8AvaZP7oA2BFVoo4FRcS0YUk/e
4g4r1nLOk51dkJh1/YvRSVXYU/WbbQRbHGBFZaQOM70Uqe9nEgClIRQiKtvoZBwi
XNG5/HZIg+gqhSoBWwjbWUYg90spFZiZmRrKo0I8FguM7VdhzYPFq4iu3R1g6GUa
rDgSY0DGD2+Ju8wao8q4cUJyPIyahA2XcDUz/z6ypme00pQru4GTcKCYUSIOy6Y9
yUg0ct1yDuDL9P/xARQlW9bo9vC0yXmeRhqPzv3FHQMuntMSEDP4Z6OiaG5YEeJI
Ixp9fcY9ynxepuw0zrxcdX/XgBhwrn6OfEBLfEwBwfF9jPPBFJIbKUHryFGJ3F5o
Gbxm+QfSfmOpJL0gMufXiLHPj6eg5nbRJpiRs75X2t7sK7g3RT4/Pkx3/TfzMJoG
2jYjQeAMjXc6l2gq+987NAQ90p9PjlE8QGvhpdRfABmqaczzFLR3C7TpedE6DEOi
WNC3+Lii8z+FYHk76hnZzERslwoHNDVvenbKZNOc2HJl8Zv5BYyijkQSWwOjkUaV
HQKVQSDIK+ymEoR5IsJYnSFO6Fl3UvA/VI0Ar72q5IFc6+2xOR9XfzQTazwUcNaB
L3vim/X3mB2u/MgVkNKaR5hbl86C+i4gEgRpI0MBy25ZOtLRFAuDVczy30Yw8W+b
bcfN0cQ/ChdWrFRxkL1WOHXuw8EZ5VxaKY+RGOQngb4PyXKua2vKlzG5LdgIzLry
OzU9+81eyf4+vbJRRE/JeWYtfW2Ea+zeuDkzPo0Glec53akHSSdLyPsg871pFUyS
0vWl+LXS9s2iA+8Tg8mowwK8Qf0aqhd1C0qhYMnalcOXD6LgggzD0KT+eWiSchNW
7nOtAIUH7qBv3+OPOAOVOggu5CNz0qFeI/lGkxerAe35SXoaY5/7az5nExIcfAm2
KAcJ7vK3ErCEbbbwuZUNCPtV4k2MtYXf86Hew+X+QS1EMdo3/oaHEfjnD9MSkK7r
WWruiX616qyk0BAJDs9ZaoGpTpSJQd0DyUAQ3AgFGIBT7YgnB5hROwFrIcnaXQ0X
LgA2TXXD2wgpJLMRYI/GrGy0EvP31wE1tHC8iwYLrwdmjuDvbbT4YKyLlFEYe6aU
Z75/RgrSxCK6XwuPWqGEyHFh1EeVWYjNGCiXDBdNp5lrRO3MbKKUjtm7rlPtb6bj
CpJMonU/N5Bnfr3tCev8k4miq3NrF/lsdAVwU1dJxK4FOz3sNqwnorXDT5G8S0G7
yc4XoOCxnXzyw+I1+LfasvUSUY6p5kn7Cg0je8jrmDWwm/GZQvKypnRvYDEybaT5
aV9goXr1085aRk1Lh+7Q6mUFIf46zweS84dcDXU8uuEjhGSfzuP9/AjVlRFIxHxa
i1jwCHprbMi7dYoTcvAXQ2awPP/+F1Qum9dtxwS+3qrxdxWbUsgb7YhTCNOQtwpi
XOr4c9QrYHNRcFxd+oQh8SC4PXuW4LeGHc6wdI03PpY7Y8E0iyZzHkQCTgl9xp5Y
hnMmqoExCIrYiqQ6GnsFjrBSoc36DX/wzoroTMIYOv35KMlo8u/7DIin+I/GL+6k
rZcilt3KlQ6Qy+Dm7fmI/fKtZ6Kyv39aGDZHJr5gziADFY/3ndpBia79PUCAdgQE
I3dEzfjpBIOj1OOFfxVdkI1J4BtJHXIWQoIIUgxwWxmfwLwZmjTbiuiEv4kiwwoh
fd+Szzww8sJ9otv0cwHqS/Q2MbuIAxCrQGhUJedbWR8JNfj3w0SyUOUtvp2gDH1r
KqMoM7Elb0FLW+p77xqs9rhweQ0MOcdBsTMVsYH0I324sFBz/lraq7AYXNE7sNTx
aG8tlXyZ0J/ZRXhojNN5xP00J86Xf0QDS0rUjMV4q10pjOreNO4dMVtx19riEBpq
GhTGNjk0hy3ctOHAUZ7pLekp6cEJ2YLlPTePbvRQyI+ZtjUOfIEvUr2evlP7es8G
jfFtdw31+lYATXHa0Iqyi7U3UKXJF6voy5GQ05TvRu+n9Y2lMQBYWbzBHq0zclKl
eQKbfdzYIo4HxuOQ5vY091hEfuLduA+HWmbsU8KtVF+pbyAYIyKYUqFBrh4qBJVn
55gScDxOQ0OM+EJ+vXXmIgGsn7uIv1e+yUFMWS5ZGJjRhIk+m2ca5Jge7yKBSlvg
T+Gu8LXIUFPjQEAHmh8PjM2VxiaodHQJQFJuoghvX16PfqPVOqAc/AxiOt+CQpKQ
immRYgmULfOa2KkLQkvMe0LjOplaNLT98tiC00b+MbGGDNQCNWKOyGA/PUCAlryP
5z6scvIv8eX7uJUcwwPOch2i+bnqlbtEm7D8l3aFJ8an5l93efa3Di60FLO4reSx
iynu+d4MRlveNWfZ8IGyAHhywEyVJJKpW36GOv0F20TOiokP3sbIo9zAn3JalVwM
3BoJlssu3lcX/wfo0Aho+sZJRYmk6C0/PppZdEr1pxmVqrG97e+tSc2NOGFSjNNj
ON9bOCIVsSoHQeQhsWs53DKtMnEZJ4hirVlYodc0kXRIefIZemsXF64QDBRoDPTe
F58BJDXmN6CAqFKAgS2p/gCf2wad8dxxILUfkG1i3EJsNshDMAyoDaquMxw1QpOI
yVFHRzXz5rUn9nPiQSegxX51NvKCChsI1/QyMU8JVjcnf6HlEyRBsD/+EeVyhoMt
CAsoX++TxKhpn9TZIngwRVp3t9BZ7UcXMfMYFO5SuxzHeF9y3q8IqADJk7R6g71Y
BnZMpCC1MFn6styLXTaZ7hI+6ONcZ71fAM9Mc4SN6uRBfw8IxyQfE7T3TfLyCess
ieQ1Vn1wyn7dzOPoDE+NBKHHX2MxuljyUFPHbCr5xGQK19fBmwB5mTLefn71z6YW
wNOA7Mmc+uHQqo3kFiffLtu5RYBYpzJMiVKd04wQied4nnctabct14ZlLHIIWhPN
Y8LsC2smgLe+0D2v3X5M1pTU1n/5hw4gK8gE0KT81pOAaQ3P64X3BCgnWREQsS2d
ZrRvIL5jdZx3k/JY+htbQ9Q+mjRByJZDg8OHxeMJZwHomS0xcIaQOP8laVNzDGsZ
S8b/W8gWZv1vYKO6141mV0P3aCcV9R82HEPUzNQZd+xi9We6qk+3bqIhAVLbYQhq
OVLCXS7xWvrH779/En9JPp5VFZjbHfwSUxJf0HLdDLUQkyRiXWBNsSZCxLYoZunQ
ExXXpFwU9p9sWqVlDEyNpmpeuteOIfY0YZrbNDT7UsiXQ0z1o2PhjxtfSxwu0uIv
DmjT0Ekf0GwS+iw2rqqhzbPoAqNYlljXJOxZ0eBal9PEYA5PH28EHW/O3VVz6FvH
V4V82dfP9yOR5W3hJJ/xXiDeTTqWxypITb/8C62kR+IfsyT/LtNTM4Oaf4Uvix9q
nyaKQQctLGMyTGXjE3LWhf+6y1hMNk7WkvgNFXktIYO/sPuf5W3dLH3qyn2Kh4+3
lgOaR14Na9S5Co7wLWgkR9HcGoAFOAAI13k/7ph2z4QzrJKNHdMd6ujAs6yvU5rW
IkhEoa0OeniexuoAgasFHCZ2n9/bivnTPYAL6BztkaP6skf2Thh2ZeKdrovjnoHa
Hjq6ks+YZUnYGQqSfCaVlHanaF/m8f0KQMB6fp6bmAXleYGjN17UOcswO6j/CIan
WZ08cpsIJdbO4XuiWGXQSnIOaSOtrxjvo2FS4Bi91SEJTKBMfbTMzpXyEJTS4ESz
kTu0AHu5GBt+3YA5WzrUFNNsZ+iJWc0yyDL2ujn4e+u0686TJ16uzZ13ZTvO8niK
q38sTZI6+OTgLE40AKfmdPQCRfuioOhdVQtXpkdesRo+RZAZEV888fyvEEfNtRhi
MkmvdrbQSA3L69Ia45Imn92mdKUwq6mqwnFTp6KBBGelJu4yFNY+FRDUp/IJHmZu
WZyt0svoX78SYEg4WlX0lZDYa5aMtFlcYKN1hI68Oisoe7SgFoIbHxFXUUnPUqdt
skwtUCG5LwO3gYISy6+1SpbEvN6Lct6LFCKJgFK/OLWI7SKknliXKsBSEk4gwd7Y
qyRuV/43dehmNv5no+k6/SLcv5OPuyfJfrVt9m0nWrYCysRewvH9CEG8OaOIS8Tu
Lo9yP9BmEOYwu8jwyJNLrbyYaom46rso72RhhWMUcYvalapMfrmi5xSDCBKv8ehS
8v4RTAzn73gz3zcHkodG34MY/iTlwfLomQ6Lxm3NCM5BxeuVTaxotR3wTo/06V+H
jarRtSjE/Xvdf0mJmaVgkGB/0TXbU4ahUIrvZ0nOtArl26Bk1hCGmlwHpCVPHyKX
nr7yx/7Lyjgsy9OIHzN64oDjQd6a2YCKXRzU5kURoPPsGBp22M8AWthhXM4J1p4s
RiNfIermMVYsg8XyO84SCRKubun4Jb9I4RcpOV15lyXADgBC8W9qV2KNw9Sa6l7z
jD5plMOlvLu9jS4lLO9u3wl4F+sDN6BttIIQwFhfAEvmibtP6/O3l0sP3bGs6IIM
ta+ikMza6orYN81OZo5+4oYWlYzY2en3AGcuyJiDc3d79yttH5K9/d3p/+vnUuBu
9deYtMpU7ILPkan0F7ayBn7v825u3zCRdTQ7tK0ldmgO2hjjFdLzwX3nwHWQVwdA
ZIqUjGnzOHMqXxIlqOYJY0yEcZDMMkchhxJnydbezKwT/hwhJX813xe1SwCcxdVx
yNzWvZupLszzLvtlphmRh9WSqdf7yKq+qu4igiqs/BGthCt6pVWDGwN58dxwUU6I
Uo08ubYkbU14AkAMtuWIgsksp3SE0Q39cMk0IpynhxrPGB99YflxMt5Q9ULz5pcA
PqAd1P3JpuWpg97QUYYKdbEZaiSvRrXIMkxoA8pmg5fv2P+0CIQey/+OWQKGHp3H
MYDKqBahlkUpWwnvUk/kVxMLbBDIWZyaHDrO/zMWRaBjcvhzq10F0eN7eBGcvYIY
APykrBTVe0euFTdCtJ8d99glRdgKionRIZnKOEQU7mQBB/bgsfISVFkmx5N6ggZB
XyXYBoCdv1D3vLeYxy3VZRroUjYyAM3PSrXToeYK2rWb8o6q5hC8+ytqcEa9eSat
1zlApGP/bLZiF6HzzRXdf4pM1LZIMJlXGCJtGvRe2wXoOdY3wQJxPGzR43quITOb
PsaSzmMT6TpquhAnsosPCwlZyfr6todop8zx3ENTgJGK7B1Jb7GEn2LSgJAwE7LF
i0Wll5M2VLa8c90f86H2/mWVZB1L5y81j8SAwec2MVGpfwTDsXncDMAzbIDWoBVn
QzVqJYQR8wBXCpzajTKiLMuzB/BBuH2pLbEf1yyOyGvC7f/dhIB7KBUqZJ+oRsLN
p22sRBxha8kYk8htnbd8QxbhT6fUB7yRwD/f4aQCvTsKKxSrpju0WYrPJ9tRwbe7
5ExIxSgPlUXTnY+H+sVY4Axv9d7zXPnuj+s2OgTQr/BPW5rOC/wqqxaBk6ge/2Sx
lF+QH9eVTIRNHeBzQ/V6xrOUA3P1Ulw2FLW/0YEzBLfjOHlYopyQ0aF/zLX1ifa1
RH1D51R6FHRCvbQ3OZ5GRwGdpS4Z4REZ3ztVa6hMEJlOIRPNnmFJyHAKe9HOyo/8
lzWNPlW97TJ9NFhSM3RonfcuxJHXE8/IlRcLnC/ln5JuTV7D5fDu/buXrnIm3mxJ
x6DAFlEWJbngEazK6Z2pzOueUduZ/9yOI4CzsKT6TfeG5NS/tUaoqB6Yj22p0FyP
TUDVkzxL6Tol2hqZdZsxJzm8N39n3r8/to6wi0zacYDq/cKvbJCyRAHHio6WeYI9
sP9xjbMmqrrjgeCbPtzOV7imD2TCw2XXalIC25CKX7s7jq9QibVnEH31Y3nUJwyC
EYpwAdkLSRB4safaJL80NdQq0ZuTZMOLWgs49djIIR6Pd20SBxrN02kM7LOSGNM6
dNvtVSgl3htSKPPSptqx8XvbmwEqiqjchkcO1i7wlElqQw2rG2PHVuLvtfXCuaTK
dKkCwKu1AEOjlVg63gBqrXqPIRieNXDkAaqEJdXc5kYntvkXv+E4CjaTA2ZRD54B
IWMCMy5R8xwgXSgHv9akQKRNkgF9YoPippudRld6DaYJWAvmXB4hxNSBZpCnFxpw
wgQCY+e5G216Q6fNqEvWOcDXW3TkPD7/1jtwOPKLLojRoHQGKt2WXqY58IO+8C5R
ivYPgax1ejeiM12zMGhfuziESrAPnpo/2JDjsPBkrdXZ+aMvSGgY0SkqQAk0PqUX
+7HptfR5QJ8vM6vQZQAKGA6TokLls7A2jhn0L5ulvN9Ir8Otnoh1Sumqz/hlkdvX
nQtYekECH2I6TQgPJvsihKdJo38FXLl653ZbKQNe495qGnpnPjP8N+3pWc5bjxop
EthwMuQjJd4mWXMv29JA7LSxXu1iF+3TXI4YPqd4kU/0DW2D/ihtij/KFiOQ2Oy8
qyqX0gOBa0mVy/gjPRMT6JqtIxTr8xoA0NjLIyoJzXOrwzuFLmG6L8HkG8BnRUkV
+Joq7Iyu7pfORUk/ds8VkOGlGx+c53g2f8Bf7XhCkpo0z4sIvbSeTq5mTuOiK5iB
DvTQ6zNVRVx9uKEzzg4NFnkV8RoEgQMbC+FIDoJeYPUA6NmsRUZAzD5VluUmN+Hg
ujR/60FS6LiuJqcSC46tID29kHc/+ZSQj47pUodEYCynzEGMsU2g/atCrs1lAt/4
2DGjVrAY6+wS9Al29SR/gjccgWlc6liG83pl1GUw1oEoju1V9iPOahzutpsCZRT9
Dip841WrTrDQhVdhR4U/vBYOeOmld1HFfN7uGoy06SeSDali7KCzmKyMErg32i8p
aqkm2WujiE0wdg4gQzW2FAG9A914/52eAVzL+hGNCYMt7JJAK0aTh1M8/v6UFJeK
I+5mJXw1Dl5fkjf8bBs/Ju2d9WZptk6nnwDCw4R9HzklHsSk+WluY6MfYljlZJ4U
eANoH5qzKGYe7+jZKKciOLoLbji5usnV/mAVTrtNtOo41d1EzrliDfjP6SR2ZN2l
OUAZXACo/RaQBkJw4uMScaATI2LqU6ywaMS8+EDL3+HxJt/awjjaL7Jx5SbeJC1v
Qm96+TsReN8tznSi/ZfFFcOuZeIhj9tvv/vN2PFy/OYx+88ScVzI2BqyXjRkhUeH
CSMRfpB0ytX4db2UrXhXzDUb+LlhcxnuLTc8J/vKQoYfKET5dP45PEvKJ6IXaGN0
8MbtT0RuP/YaaHZu+HvIrL2pbZDlmmGoQVXwAZtURzVJeuVeLLzKRpMcFXHDz/vz
40p4ARucxnu+5fTIXnb9QsIjnKKdfhVEdNl73jVXLZ6OqLm3vCowtDhLpxUHWeWl
AEqsdKskHeC81liUwibx/kGHkXcNLmEo2CP/IB+c/aLtfOvMYOTdOya9k3kTboGP
+S2ZoYQ/i2dhJwQUPgVhTpsnJO0eKWXMn1D1tQYVLqxn/rdRZvEI6uo1MeRPuXyL
x35XJ4g/TILKDsExglaE7LJJbW/cqKtgDa/XG6sJW4RFFLia4zM8wACLK7TdbJM7
ihr09/WB5e2U4dpmaeaAfU6678nNsLMFi9h9StYH3b9ES52gTTDWmeSY0Top7H93
NGankW86ijnhcLsTzVTOWx/kY3LAbcxlIeeLapPqEcdLAkBW1hy6n1Xdp6Mrvj8j
8FOZ+ZrJChbXS91xAM2hdu1tgFNK9uxq+BbdinYJe0499TCHA40JmwmDTfx2rNzS
WqA+WQ3QW4MPtzLm4oaDE5PrgENkh45Q5DpQ5qfGVRALfGdHg0e8ZNb0G24wyFMD
i+YNAGXtaWRbEXngSaEQFFBD/hgMB3VgtiRrBtkRAmHU+SrJuQO7Z0Of6a25OQAG
/c8uD980j5hlGGchAlssNJlDV7WZQsckx4c1Sg4fe312KI/QDy2FnD5oKD/dPd4e
glJuEh6pxNg2uPoLkAZPD8feKUaxh+CwMzvrboBJigsqYh2HJGK9WZvHpLLs0OnJ
F+hzmfFdxB/LW/D3LNZ9BhQuJmcocLcDBU0c6kjJK9aTBm32YZ+ehx3Y+pDskR1m
hXmD97VhMHfbQNu7bb8UhyKqr94BZS8IVwO3o8HePz9uP2pCAqAWgTNL/CaB4K5p
7T3TZU5xptJQQRwaW4S2ghXdGpe8VO0NxC2PsmV2vCLrFgDdW+tb/vHx/8JqAgxI
zJp/f49eYUtB6vwGoeQNczDTlo+5zwa8QCFbSqDFqTNKLiIm1R7XFpz+cyqvZrBd
eWeIMBpnnn/z+P9feTxROaKNTwgeNhgczB1yj0/9oOrfTLgEbfecrcBK00406sQA
CV0LkuxLGo8N3fnp4WYKj4cHGxFO77WAcvzgVzyRgGNVQ3WFdD6MuwmNNoDVo0ES
L2KTq5cj8r02ww8hFir4Ogi4IRj9IuWU3rc26U9Z0afkROgmVrEGYfjrHbM+ZLWR
2V+UFFfANpz1RyyeZCe1gepJ26cft6Wyz3NhNQQ4sQqeqrycxWrTOr6urJ4mUg9c
iJJD2IRSb02lmx+UNClVALlaYlcU+Bhntovclb1HnjbwPRItrJoJf0eFT+u+xETr
H4QZqWwjq0sTQi2S3mr9278CoUBD/RFxFknE5j8IVZP1ZZzNpo7dy61Y0c0hpycK
8Ayz+4hYx7uiFdsed2NgpTvU5krM10Ne1WKhLf8a4NGQs300rxf3RjMV73DYlgHo
c//kjOjzAFqSC69W3/zHvBhJf8kutqZUgjaf1O3QI0tz3QUd4TxbcMcteFv4HxWg
nv3Sd04pqwIc9G78tpafJWWDRhboPr3xgwvcFbEKi1pWpDkZt4h5ttHgkHmyZ4Yq
Q0w92uOlqjpv21WdfMbfjkhYM3DW9IP253OxOxB5aXA6evrlIudqqG0GqiLQFJeN
zxOhVqkCqAAGrCbidclnsNcI5RTSO/LV23m/uijqnMfU7WAAYQoJ+0zwoeMocBQq
ZEfANvKpzIGzSSvzbEsSP3k1q6s9yWK0bdt504HIZicrQYSnYsoWnSUU76r84BMh
O6tJPQYU96oPXNoIRxcfVT8eVLZnF4SuOzu4dnSWwWxMoPk+s8IEeQvAa7JisfpF
WP9UimcDRfhslUKPZ8hWlgQMrsJ96eLU2ZN1AoZmfQ5sJPeAqmMRDF4VrBD3exGo
D4DDqHhGj6XWszedes841nVgYboAAgTniZ5OuVZogPwAgfp2E4RaZUGHE7LgdOCM
IEHrljdcApDMv5LR/Obvjo63J1zpi/znQ+7VdPI8irCwHPmfqgTCZD/9zE/DanM9
RDheC0l3DttW2P5iHMZbcjAPO3k+l9foupAAzIuSzN5KWP/GbDdU7KmA0nt+Ml7k
AEJ7WOWK+tUh5TaxBzq2LVSBWVMYuR5d9uMJEY+kM5EUXMfNXG7E8OQFCxcCOOek
yAT10J11OJr/xC1DtzsPr+gQwA58BhUCKqtPd5Vn9n7TCnaIX0F8lbygpP8yA+vz
BCiuh/IuQijAv/zD7bIKAKP1hfDP26uXnEJcVJdInLRjbefL0KenoVMWoKCU6VkH
bSJ7z+FeeYYK6RDQoSRlIAWI6HIx6c7sF+i8dPdOhE22hQuMQXtZrjt1OT3BsqbD
dLa7DexjiXNHA9bqfJC/DlhA6U91Q2moExM05yWdJPh8h8x8kfS7vr4KTTxv4npZ
TCQjYMXiCedyso+Fj8Ohd8NXdqpbxyjxsyhpNuaattO2v7e71fkG4C98W8f8qE+z
NRW63NaRcRzCz5seyyspuLYqbu2h0Eitl12jBlVYStm2SZdVlzmdvWeu2xupZnry
fPlfNB/937ZLRg1rA42lV4AlsP/uuqLAhNUsALK2aE0X9Im89ekI5DofpPmcRP5L
sDDcatGnYDguTv5HhK1lpjNX1cnrnqy7HqrBUUE5rshlUaTCpcnF/k0YIrMJcqV/
eoOwULPpYA3Ai18JH1BByNlVjcRLcEp0sO8ZNuqs4E3gi8fIZ8uEJ02A+YjNQEzc
3ZDYuxXkBeBNQsy969do/SqWiogjLryHnT2dCRLnMoaATlN3FWfvQ6JZX0vcuwMN
2yj61PRgqtzk1/wJl2/CzBc78v+V/07uPrRqibrEUaGNWXo4hlFeyZtYKsVF8p/v
FWpUPf8PrZ5U8KJWtGI7z9XKNH3BkUbVIGDN/hKNjKDQDpBGFKDsJWgdT0HLypbn
03ktUfQ1fW16Pz5mgOmzFl1RIJ9L2m6/zFFmFByqhRTLxytEC+cuyKs9Urj2/Xjx
lbW2bP4N7nPT8VuwRXpUfwUksgNVnmOsZJyzcaC3tSkYd+FKPpX9SoNF23N2GjdF
SFZWdWNGVI5n+qgk1H+heSxnvd2O9KAqOSW8O7WC9rbTw0nxhRjskoa9A0CO+993
Is8hg8Tu79iB4/Oelyklhueo9v8gLhVQA+FPwcskqlER5DBapvDCP336mBrDXk98
deoPVxHmdNNAibUJ9f6krH0hPEy1hhMTH52IShrFmEveyDq4GznZrmILga38sLG4
nGSVDhbZIq+vEsGQ6JMAwkMYygyaloFbE9McXt6LcsJxCY4r8a6ND3m98uK00inb
bzZjB/hWgiUEvhcU/A+7QaAzlHKSxIRdiG55Fvt/FmpT7OZFzjTn1A/7XX0mRxTL
IMxmIJOi05VVxYr8JvQhS/ViJs/Wf1cfoTm/uN5vCw33jdENipK0iOvnhcBFy3Dj
VPcO8uxux+7UpMlsokoX6Z+dBwp94NpZTNNPRJ/AfQO+UKxMv8exNtVrnkm9G+bb
ygxN7BUrXgDGEi40cPSJgPN4GYBMbVVpY3UDEoyLkgkuZopHLBtkZ3FyvYMKQZGv
h1vBAJKRxiuVdUfsweo4Xa35NspWxePc+pz5FGdQkjSrPSrjOjbXCNGVBeMmFLSd
UIhca9SG1P/L0Q9cuZ+UKEfIlR0IARLBa92k+Egu388cFPUB9vd2h2K3SLN1JOsM
j+aYOyL+50VHFI7MqOHHPEz18IHjMZd7aV0v/Zv2Ayws7K22UjCIX2PC9S2muf+M
FTuXImpDUm9RmGukXH9Nj2TJic+Nqg5+gs3UjR1boqpzlhqn+mnCO+D0yHfX/CXC
Avxvc+4q+62Vf+o+6xaPZvcyFE8YVhKfz0SoCiVLR7rxLWJmAxYoKBmByrQYY7ca
MZpxkJJva+wsTb326xXMnvn+5HqcTK0uV+G74aXcl3R8f0iuWzJ8fk+nqcdRsh8S
UozAh8TelEGlJSVgw/vMTvQSLvW9eE1GCnxhrCLCHGQFTf8szfkiVE3SxETkBSDP
Po5XENupYZUK3AvlKcw4+aJULZyhkZrcBWCIj6wV5IUuM74tSwwpjMA3mLeQKM+5
Ech2iLtG9A/yO98pjJp392e3Zqk0lE7jTDu9ZNyCTpXtwkUTeXPjNGeFDI0JQ35M
J2Ktm6qihASQ1iYnsi4qZA6wGgKZjShlthXVdQgs2IARGDTVyoU3iCpcK2zvm1/b
7NEU7IuMVvSBvI8Xat/6tSueNuRu6Q0vx8km6WXUku1V9yBb3JqV4txmGJ2HLv/7
B0yFifn5JNqsdnda2yNLye+V4Q3sB97ucc/cy9krs3bfMPFcPynCCaWf3V53tNdl
OhbYyKPLarj//hmE330qskI1GESGPDAhJMrZWs2xedFCp7ZH77Fq/1AP/M21VERz
QN4DVLS61AOyjMhdNuLF4r3MkzoBr7Bv4UUeBeLFSCsv14spnCMf4neSkbZefG/1
lxdq983ajkC0pJFpUWhBn4qIZvuUiqAJOxZUsMkW5yovkScBx/sv34Ppphh10HcF
eC976hl4/227pYdAPYioH3k9FyVHUpMn4Oupy7vCATPFVDTGTbo36x1LVLgnZIEA
2nig7ZmVB+hOgH7afSJreWQbGJ4PhjLJo/Ak9MSbfWpVJo6gP+/sHISyZn1D44H0
x9c4cW1JpVhXvHkjr1vrrtOMjxSqqp/alDj0YnQnzFPZGrt3HTeB3aXXMt+rCWk8
uMKcrTqP1vQII3A899PgQhBJeh8XxBxfBUySKIt2hwhbm2zYfBjSTW/rt9mpp/J5
XR2DiSeUu7gVtxyuRuyIwVOZ/i7fsE/0k40UFHSutIZL/uiy0bLhoJ7p9I9EWBWZ
b49I3FgffoimU6WXXpjQtYzxeFNpKaM8rm8Tq7y4KQi16Wb2384mf2wzrzB3ymvJ
ybCUasyhgA7xmnKR2LJorgwtnF4i9oA0qdNfWfnF7YYLscA4vsOmsHkpLFihSV5u
rw+Mhg+LgZ/KLV6Q+/4c9ehst8aDvcmvbxJCFZ8zqBGdpLHaYEOkpPWpaapRJL3q
flA0iaat0OwLTs1Im2iZxt0j7lVy8VIJ78JpulErG0ONA/NW8a6zMG9eYocnAfpa
7OMUd8QqMizb1/FYGyg2xQDTQdL+B6noeiT4xqurr8R8Dxw2T8oDIuPhTBe7IYop
rRp8QI8ioNSorACUY62q/1bh/AVekIMZNieD9SdoSyqWGwLgA1zok/b7VAsXqs4T
I6YRbgbRZHs8DOdcWCMlB1VQ6FQ6BCXfBxFLnd+LhclqXJ73IZ+dv8DLiDA80r+d
O7Ch5Af4fkTA+2Y2Xsb8j2JkzgrVbu2yBZg8jvESB4yIZitTLmy+ZIucFDv8U1Ql

`pragma protect end_protected
