module altecc_enc_latency0 (
		input  wire [63:0] data, // data.data
		output wire [71:0] q     //    q.q
	);
endmodule

