// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
Re9yV94LevLlR934P0Uv3vKb4uqLB6wC079JvhIDTUGwCzP+51fuZ3l7TVdpkBvT
rqrc1DkFraGQIrspZAzH8HCwcS3xOfb+GlMJbKGZTq3Udh4G5Y+HhxYMnIuTJRVG
MXVBqNks+uZiL4x7LOh/pbYWf2bO8DrOr9/ZVpyzpjnp1BZpVlqOvA==
//pragma protect end_key_block
//pragma protect digest_block
6DrEwxSlQYQtsnb6dE1XUHxV3fU=
//pragma protect end_digest_block
//pragma protect data_block
5kxpnUhrOUgsabrGYMiAdFFT8f6uj7hokevP9RTYRUdFf/vEgbm7LJfuuNlAf+hw
V0kooTf9WLuLxXQ8i6aqEHjdFfpKknakpHAau4pgO2B27hfX+V6li/OjVYcDZ/2X
LZJiTg3cFCdwj+ynvjzk4h/aQBX9BxVYnK6pcnHp/isCFpLrYWRdxPv/WqiYfp5/
dHzNrQmaQlcp7c4wj3QhEvPQ7pLSYkCVCDgj16m4sLtEgF4+z3PjZgI5wpdGJwII
n8r7e31G/NhvSyw02kqhLuRVPRcw6xDHkF7buFciNSmZeL9phSrrzKr8Nsk/h4h8
1AbVOvBLECZ7wlva9c+eq4xwaiDAr3DQ7dp+MaR88FUP5U5q0fGmMeT6COap3EGM
mj/3GGm+rw6wdIGp8PsLs8U50NWZw7ogZrx+PbWwYiR++/tCy8pGdRNxLgzrv/3v
WU/8ufxLl2Psnm0FPlcNrSYwfIKGYMH4hywqmMRso8FJ+ujvY9/cKfyne6sE8OlK
l/Zl/8J4yQZQCUFOeMoZqkw7dsyAR8R+GkHpaIfgHTr4b0ujIIR6op6QFYrAEQK8
7nuDbl6L2e/3ufFIXNFfGYCQTn77CH2jFJKj72VVKfWmGfnXEarX17J80bDlBXuf
bsKFG9ZJaQ3kVfOvgmBX/bhmNY7exZqVtmbOskm23Cta0QMt7c6ov6SasAHW3dax
NqggkizarsLauF1lu/HEkBZwkxGdDvQT8Bny7cTc62n5JfxAffMIP5eqXxryUmlN
rEt0/uRhN1Zz1oujNfZDH57Wi4P8ytUnrnZCm2lMs6l6EeWt0SlXy657+kH5M8QK
44WlqylJYgkSdy9znBv5wgrgDQKAmcssU8vcE1WBajODcygdBDtShvhuy5F3H5Jy
SUjwU3Js1uPC9k+F96fl0K2bnj1qky6c39gv0dTYM5lf3XST2gmZ3w4R8zV/TYPs
deU2Np023ayFwW1ueSM2TTfOV2n0XjJYvt6BTRUSvmmoj8Az1VfOoOtrqYgI3iFp
B6I5YBEXrH5OFGuEqbh8KpXI5Q6dsySzbTJSU+b+aVVpkJ6f0bG+aTv6nxxWhkmw
HLgZC+VWMLLPcqqgdZFi4tZXsbtRFI7OG/576UCy+liSMMvdG5k9PNJJcPuCwWDb
ngfXPSb4vfMkuwBO1grw3JIK2wdcEKMW3ZnClbowSGppnVyZjdkrR1SNpkWFVA3d
ybFcMneY4ds3pp7UbHCOoiiQSePRuHR7p6AOwkJiqsV5ys4f6lYdotXqJVrBPZQv
2T2W1mL6KiHvuZVqgHjTXAXk04V6iAGHhT7TzsTR8UVsH8aiD4cm0Ze6WtFrFczb
JygwiFRa1Tc9RBxQdgAC++4vuICzK887kE8pg/WJtj7oMsMJhWAggZ8x7j4/o/PI
VuQU6k3ZIhLBPu3bfnZk+K8wuUcRoGXO25xVWpZnPugvRAx96E9msCm81e6lNo6y
z8Uhc9XditkyQddH3ji62Ke1dKe4ehGC2EQcz1P4W73xmnyy/HkNmIIORF2+zfIv
hRHwvsO5aUW4WfxD4vHe5/FcES6LRzpVMbpXza7DIi6Uh9VrrZCaFh3HBrsATPB1
0aV4dGxLSrq7J3aOi3fCLAVge5US/U8A4HVHAuEcI/WdUXS5dkVMEnvcf5Jb8Rk4
6q7O8XybEriEWnY2+0bg3hhv0buBdVoeVPHwcSrtHLnsfYZDMmQoYRQMa2X7kZP3
+S6b4Ltb6+v+djnoluwaWmaoWV3ZP2PDuz/dVb7UaEJNi7cOoveOxPWghpqrbq2q
671D8b2fzaIk6Fc/27fxPY601UZOVEnPMuyBPclr2CMDsnb6dLwpGFWBHq5VBaEa
oap993hZZbsIICLhz70gNrtN9RyoS+jUrIvM/3mPWKjRdiL8hheVbfGRqZ6KYtJE
h32kaFjqjfYc4g2SAiaPeGQWNJPII4vGsikJkN0P6SpaHnLJmn1x65FAQlxgpfBF
n1Pnd+W+dxlOZrAmO20JINYCsYw3uEJONdnCDc1or8GhEx71YRtYthj85vnaVjO6
nX7zMXym0PAOsu2vS4svTbHsvCec5tlx64Qb0ZycpjqxLvgxT3PQKPG6LoNwRlYf
NnAkF8BpljVDGPJ/9TBQkYzUzga118GA3L8na9Oa0BFprB4s6t52jrw2c6NrNswV
m1pACFVhVPsSEzbq7sIkzTrTyJRacCxE6tu0oYk+k1QlA/X2QkgIn2pH9vs69sRW
ewpQoLCMEVMh3/a3/ZORD/uyOEOioIXsFOJLNSQMzDka6Ulh9YeHETduZIaFlhjp
Md/tEkAQJ3RvT5IBZn82Zmm7zovZWs7RaflGzlOiMDFmuKKxjgvEWexldAeQe6Zv
Wm3yjkcr0gXwYiYYp6TbjDBAVO7pM7Wxhri+5uzm29nH2hbS9/IHXdsHsrqqMqhZ
P6C7ZyXKxNVKgr3C+2aRRzfkUbhQrkH6MAeQ2R2aCQNYGJ5L/vhcPXE/8dtFhszW
300SnX7zzTJd4nXat3iOrwiMFFi1yHn9H4xpjuXi+0J8ma1qqaqIhnMp7hB8Zz2v
pkv6PWZLSpu+EB9dmLObZTY8iMS8qAVwh035QeDFtvPumDhPJuUExldXvc50U+/h
41b3mQk4cIqbmfSuU3QIkDqCjPOQx6e1Ztlx2LD2CZWtvCaQwC66IrLqQzO+HsE9
88bW+275ua57OPTwRltVov/2xATyYIBGcPqFU42FflU7BHaSOjavU635iGekgTRH
2pvLO7RnXcvmMyvTgE9vZH+otQ8aSyEx2HIlJ4RtlPG2T0hj0bJ/95jVT/AzuOlL
l40AROHXUzMndwcqmxNAfsJr+kHF/Lwio+2DZoRgShfHfuVkB/QNsuWwNde3L7zo
+i96qOpy5NdaQLJZeMN1bSdhu6qMluhwqqHKH4mP0cwOPDVU5+ygDGcRAnfQ9wmH
QLDauk+h/mzN5kwmO36GiHbAZTRlZX/NJFPWcTIfiYuB0c3e0x5sieaQavvuoQFW
6d+BvtGAb0UZPhL8Klw2/gWqThc0CrIOSmdVb4gPhRIADtljW2STJWhCWMkFCsPo
VIQE68/5ItHOcU1s3Eyw13el25KRNYNh0eMpG+qYM7K00q8fSvm4W3G0ebuGx4ku
lQhJq+v7a62StTGfVRjxSia0hEsUGdvKBSG6tMH103BNYHrGHEiK80wc3af/jJ15
/XNHQ9Mt9V6ESCj5KGAoeGsm+PzbpCH7vUjOgL0C6xj1YPn24KL3bbq6eCmV3PGZ
wsatJo1NRRXJeiy61UZikynmD8Oux+HhUzGTGcAlYnH4czNZPjxT1UfleV0RzxhN
kNJ7bmycFFmnnYNlvLUwRep97v+RdaB1zGQoAcA0vVLsTO5qea+d9SD6PXFTyeKm
U4e2tFWchJortOUnSC2zzAEOez3MWw/nH21Va1TSjvrF3VutsH31QJJmD+YdOxpU
Myj+5M0USNfTAF9hMgYq0Ws1xv8zjCnaEZc+YVf90isQncYAB5bltizOHyfbyXZL
+ozPK4/Xtrz4waGm4K97/4rWoXQXU5mwDL5Lv7uYz0ac9JAPAXeqdaNjuJx0bzcg
XIrLIrdFZk4q2hlrlRVJax3W6Z8tJFfNmFahub5CWgpFEFo3AQZOpznZHSFSysRb
4t8nIf8rZ/a+YB7PYKDMNZ301dmcqiI4DV/WK3Obct1EUflqh22+FqxZ+2rkKF75
E60AsF+MamO4Wgq64dklfMWFmOQhTGf/CExD4kvLAUoPilbm94CqqzWCReQgKmUE
LX2ygsQrpAe6/P9yq1uS7eYj1+TQCNEQpUTgr+daHIXUpx4HBbA842MZuqyNj/sj
yU0WZ5w/UuMQImKSsIaVX5UT4yvPaIt5FGDDVAw1z4LUG9Zs46g6jqUVkwna8hOp
TXCxM/tqWNJsyB5wua0f5boxT6Tq/wk8M12KBNTSlnU1e9vRx8/AykZafe6R6tGY
C6xDG6CIZOXowsrasPFDU7uXGov0YuCqJ4FMLUKTvaaqvVuIhTBCL50urOLhQyk2
5qi1/hHRC4RUqrsVaPzhIPxJ/SbMnc0Y0ultiI/lr49Gsf+t2yRofZ6ySDDirHCZ
0x0/QWRf0uPZOQnhVRujuBt7hb0x2gT60cdej/Bm/Dd+eXsIMzx3Ze8+wtbEll3f
yHRtYTNQDVkJIT91apZ0uEkghJ1pw2RtfPqm2ItsqCiOWQ46LoQT2zY8SVG8WF52
HlfSNeEjZVuM65NvSHsC8HkXNMpTDgwG698/jR70KW/3oIZSVK8OmeMg0bDKzCB7
WT9xjVD64EcqQ4tJSpNI6kSYPJyVvIpks2/tQsETZnPv3XEEVSBfHexOTgs8II3/
JchsS4W+sWVUXxxK0ncdCY60oupqXkUPRQKyOd4uP7bxh7Tu478njxCQZ+wRwH13
Nihx1S0z6LlKcCkaPaeHAogfcLTVVrAUIH/71walk3IbbudcV32ldeJx3TQzKfif
UshWXwDyLNt2oi6IcBR+Lk352eEpWTSnooDjhXqlMQoq252gqjvGNxYrigd3m5Uj
wF95fVZYykOeuLJevaFVZOtgbs7KQibjd/nZP7FogspWVetOxdovINZA4U6CJTRP
0NUGNxcoyaVliQBum6BNUCjdypGvXRByA+Auj1gyL+SMQN7Mfy7BAbqDY38xuPS4
a5NCQ97Q5u8dGPldFfgm+4GXhZDrL6KC7vykD3RRACKBbuJYFGRadCOSHZTPTN0k
Y9aG4FklY5fSGJlNH+SZ8SSoVAijnx5l4EcFlqcunw1wbDD8wqw4EGjJVxU5qxEm
r8KULGLjTEVbY7l1Mt4ut5RpNTpTmmwjXSvaT/915zOKPWq/iZGjy8s+zw85n8Dy
tpFlIBAClvToIKOw8EkQAXyv7ryycr557v4Q3AkkEv3qQyUy3lMhznMGnWMT6CF/
kskCf54lozUqu/f/gK8bR+0sJBWkWViU/FCfznVmt1VZa0/Sb/XZO1crrNtdT/jc
M2mftvLFffmuavBk4PL6vx2TdAvMvpHwSRGFBIEBeTVTLztksW8VqGf880wBhatY
6ZFw7BXg4i6DKWxOlOZZUxC+CGE8xfCB2QDipX895FZa6qy7PRga5hYoUGqfoJAv
oOSqdasg+vZu/j35ed9d4H33i7M7DXJO/XMGwPP99M9BcuTCXWMfBTGBWFs6fuG7
CAQV4felonuAMjbu5f0a1G8fAL34EBI7qkP/7Xc8rSJBXHVVWNkePryyxwKihfoG
vcuqSADP7Fa7bkIo69VkIvqXupcXWujMHCTsGlTbZP0NPAGyMZSC36uQ05+7/TLq
uOb5QN1WRFDDM6NkgukeeR7Uuc51sJ8U/jFJ+MfjLwm5yRT3XDtExwSzWjiAdAdy
CjlHt3IEn0pab+R2umNyHONHpPx2O9ZuXHfbq+8Jb7q8sB0sfs5HVg7vdZqmxAM6
A1Fml6fZwxQ1Kp1acJDGrztUX4xs5vg0QjeiLMd/xvzb1Cpm6uD5hzISEdcX1nWn
vliSaE0EAX+fgCKeKgEDAYyUEkccdqMYc7f370ADFKZk9U1/IfzYcVznPhxocZ8s
s42muEvkYZgfc/Yg7It4MSvYQYMWsnzMh6iRY5NthOT7bp4aojK1Bo92GMYFN6pA
RT2NhNBcU/rM37lpDWppEi6Ri4fb59riD2T4fBEU/LA86rQ0wSqPoqNQ8wTdHylW
btQVwJryfMeJsHimNtTBaz8jcKtaQQ9hVdQsmKSRbDrQyJsDbfXQ/xlXGO0jUApA
kDfSvi27OEodN1H/IfY5lNfe/294l0jsfkUAcxIHeWFoS4pETkrelW/qefnYzgIP
eZesjIl6eWwZdD6iMBj3XtWfmoNfSxXUQPODDl30YzhLjeMYoJ9n3r6qZAQhs82D
icCBYlvRWwgUIQ2a1VerSFaJkF1KiKJ6tQuI1WCFd2NzvXzTentl2m3bkCdJeuh4
d+8uz6tCTjfmXplVKT2OOhrCtmRUdEGQsVssJVAiENpWdbAnBsK83B3MXVvyOs9T
H14VCNSIaSt0110GA6ntRTYBMxZVMKHpwCzIX2dYFJwk92TqJ0UzudqYOJ6So2Fb
1hIwLcZj49CZSIq4jEUZODl3sNBA2+QHSOfrF8JpV8s2vWIDMBiLMD6kHW3ifBo5
MKIZPCJFdhoyBAVmlB7s0+TRcuh9gRnlEi0GJx9BCAgUu3LiW/NPhcJJlHgD79Os
OQ7Dho48MKpSVWUXWbub8AHQmex8oucuSr5tFnU2KYadmyn2A1S2rUgJh2jPYtwm
uNsAtnRgs7kjFlTErHA7zKTgaUUd+Qoac8oNcpOPI8TaWyOBjTdB6QkjXc+QjlI8
cdbRqVnp+NKSQu2HAnLpemSyHuqsYEamxrJjGeMuWzC3+zSZX2DICE5wJVvyxLEv
af/aN/42DE9QcszIdj0O/GvoVowL/qYel1/h5kuXzW2YBfVdJ0LEhORuS3tXP8R/
5SzQqP854UgZZWOgDixRlifc+vv2MsRyIhmiDRGTGisvvMKAr9vgNwoRWifG8RCj
0OS8XBlrkg+aGsA/yIdjcv3PCMwyfzefOwWu+0n5d7yfhBsSQlJ2xvaxoP5a/pZ+
unhwD1/R6v0VkM556ymwBwV9CXRP5Y0NcVeZguLYFkenS0XAL2FHjd4uIhNo7I+4
2G78kZUIs+3FA52uHxmhRkTNcispTqJd0QZeHvMbo3EMwX8SZ1O3rplfMKco318R
m3ugr0wU2OTq9E4RIqmX87BxUT/PIKD647pHq9Dj+aDvBWIrs5U2piAZTwmrBzb0
0MVVZrOPaQ9ZA51cR5y8mu5pZfbdTppRtm530sUz0d/DYlnxtbG0Z6nv1oa0GXqP
cAG6oSU9WpQcm+IX9dqUirQ7P+fd9b/kUos0sLPkMAzjzo88rv1lY/TEaxBgu+QJ
rn8xKrc8hfsQz+djkCYowGPwRCyKmjYb4EEkUKqUB/P2ajd1ya8r9wYaj+d+pM2W
xTnwIJCtRDopj0XlaDkbd92LjkLRWb0Z9KE5OWERUMgWu2RAqLm5PA8zlovqxVrG
D+wTmFhMWMi0ZLRgmkuuwxsLH/Xxll1/g3kyWaXoWxrW11l/9Tfhlo144J8TTtuC
Iye1+lYFk2oc36qnGe4tlWXLJ9Y9Qd6d+sASGtq4Mp+TQTya/5DepoyX6AIV5Bsd
lVPcs9qacSzUUhGvsvKvy1g1Pjj/2Acj2NYAH9LSe9eus9vrhK0B1j8/I1bABm44
lr84PFTs/E3pS2r2ACZrIX3THz2G2UwCSqn8LFAtRTzcaeidGKCyx7C3CeCuFx3J
W894z+vwTubV1LiVNrU5XFEGGaey1XaArw56TU2AjIsrm3AFFGl6gPrsQ7O1ddAc
ZePOYLufY/pLgglqAdBYQQyj28FL+Y4N9LgdypQ/hNbq72OPF7lg8G0KBIf7EB1r
CMAXzqg1vqS487GOEVY7uIykv7Woh4uwsBrRfRjZVQ23PWcK9nqxomnD4c8UOlrV
ZKJzt2RMzxRKz5QPjCahoNjB6GfsqjWEK0iC9WJ0xkjcYFwheGNSOyehPbbAHJZB
ISygwBmxz/oWW/fMhStcPaTanfZGPxwWy/SHIIxl0uqQOhh3r88C5ARfvdyxBPw7
hUNXuaaL2SKvvqF66DZg/mAxvYywqn5wYcwvKCsFu8A17ft8hSb5pny8Y+AsQZD/
HbTIYMImNZZNC601Chc2+Mm4pIKCNed+ynI5Pvdxg9eOCB7uUxaG3e/Gx8FeGqrN
YyoMCpfs0LwkbtrgkVOzkVeIwz1A07rbncxzGwjuQFLnx0OPQiezbDuR6+6l/g/9
YbrDqdPQ0HBo7zTz7FgBgRDXEs9JRZkuxwgHt6TOtS9EkY6qkr6bHF9XuaGi51p/
gSb3LO985vFWOaRlhqj8sAX2SwaMgGPlrJBcI3dRXT3QXtM3fXE5Jf9QpiIINRFp
gqfpOlB4Jt9B0pQs/FPpY+MXg0zGBIJg6PKs7p7tsaVcZNCIa7s2ndgCCShtwUzN
WANglzmKHHBzWlm/3LBGg5ajT4p5Y+zPqt3YYWaWmB3w5rnCdtc1GWWISGqUwANI
UrASYRcj9RyNBI2GHTLVflvUPOp8X/QQeQDlr8jLHCQed0v5gnz3+JVPaiEdXuaE
hnPyyEhqPN1UX4CWmRShm9lBEM6ApY/ibG/fsnL9HyEH1JBy5+xee5ZosNvZghqk
LZl9FG0qeylVsEHEBbKBq5dpV/gbb8YBw3OxQaWxkF7sFuP5tynPPjswtxUA5G6O
T055TCEbmkdxGNkzU891jPnP2umBC7uA868Eh7V3sQap3I31i2jl6iHYoLTLoJYs
fodZCM7k/9sdTqIR6EmFlB0eBesvCDsB+Q0zgZAjHjgzoueOe5inDDmwdLPfCxj7
c5chwf+CIErupaL04MmWs3+/Hq/QOvGzHLFVXNt3g8dScmhRpx5XZ/Jp2CbUg8xi
O3IDZZyfnNE/Ja+4Z8RmapozmCOC89pLEp9bWU1XkiQ32hrPy2NwHCRl2h5giiPf
mW0F+5gvFKNAfeJ8ZaB4u93Mf0HtVTrFjFHH+5ZDUeyp82uutqQImyvegxtWcmCu
T4m01kvexLEHpqGqoEgCoIY7VJXKuICxerCCoRWrwO9IvP5cAyJgw1F+RJETZq2c
sSdPe3sJv987sOUXG4atR8OdN/LmgTqBCe5iqTutetVDqwYZ2DDlysl0dY6hYliF
gJN24GNccsIP88dcU2dc2BKmgcIMJCusvdK/Z6JAvlSla0sJvikGZy06gAzEBLaE
c7BPC1NyvYOdfKwzLrToidieqszLrGQz6jvAYL4iEbONnLIWBj+CSh29tteiLWiD
LKvY4JjbfTwmN5I8QLDBBJ5uFx4+YSkwXcfA+R+AJRwI0+eZP9AJOOChA+Qwwzna
od8RdCzx804cbROChnNDOJVuY5nk7jjWZUlZbO8u9+J3NJLDjVS/IItn0vNKd3wS
x6E8GHLjdL4eYyREttpQgVl8w/P0sXJjk3IizRZZU2Nv+fFrFmZw5lTKiLCJrUO+
QKu6dA7E1UP7H1C8bkethq8dEfLdaA2Y9+QVGNVmFuj97GNVDRrEvmzq0cnTVTOK
BvDIIn8bGC+OyTDviNLiuTLn5KDbiyip43s0ikXWH54b05y6CKM0SlzIvVnlNQvr
DUEQMMiOotRaLuvKJb7/34oHM/GtMozkMZiAcaHykASNaCW6wdEmfsmeCfUOYPaA
7oIY9OqBVX4ybpbKSLoS29MeLiFrkRqQyoopYKR7ficLcifh66M6nGGIbX+ELtD7
SwF6RgBf9Zpu1aqkU4mFhhEbABTAcj0uUZTUvsijOF87k/nN1Yf/JfzAH2wZ+y6z
Gl3s/gMLCU7oFNeOYEiHQrqHJSoQd2n2bvqPNvxF5bXEa5SpRk0qCkla1DnM7LmB
Xk1JuT7HGOihLbRgUu9fwEG8XkZi1h7SMQz5Unq4tCdRQ7Vo0EqNWvYsPeziialW
tLnGpyWe4jF/c6LhY2KDu3ccoxkevc1ggOhvvSl0Cp9iLMTJXKvOHa4BaK117RsP
9Zr/TlEXtiTDWczVTdZpKS7Kmk34NYJh6CePImYW1X/J5ZsQpZdJ/yf0Pu15YuTn
lqrNz4dUgAv324QAqvxlMlD/MYpNZRoae/MF4pFbu3tyjz8NnXTZeNjQF1UuLhKc
dMmq5bmUWDVBjGecz+uHSGoIfamKARTNzTVnmz+FVzoEOekKva/eDHcS0bMQLsD2
YnAtY0+zUK5DIEQEbIIb7yIy4/AM5VozEbwvK3CQQQRE+gW1NHitZpPmGfKAUAR5
zpP+jmcIt25VMN18IchAX5sWDeQ8FJWe3grRrjbegFjwluXTdoF/sWEoWpmcqzv8
b4grbCcb64ZxV4/+6Hjz5E4u9h+k0klcTaBOEwG+D4OYDBluYn4BqARKILYkmKaz
vjDll4Igt0gg0gSSHyNVNnCfVJvpLXo7x0rAUbsIo0xk+ZBSmx6n6t03FviLcP1t
TsD8mXz06ui6L43ecHHDZbXceCzTBc+eRJwbQYnaSMSqVrVDV3GOBWhwlblNKibW
LivLnJScxkCSsoT07Vmri2EfRpVEY7XelixXPFQGG9IQiHYrhgH6dmRIlQQwzEuQ
eUv6vmcyGtE5sqs9oMjJjxtKpw0FtFURNT2P2EaHyRWYebhw+uQPAXvxAxdl5AxB
mecRvFwJ4KQDyBoqiMr+U4x7HkG6qhW+/wIOdflsLXXSJF3ynKCPioK0H4LmUzrY
W/s42EH95sFybvOUq6GzifuhjRzg8jpgshsZjWExBjfee3VURyJiOKl2JOEdjegz
CF4JhnHm6YG7+hVbSUROuQFLcXWKTFId4ojkTGw1CZBeoMZYjnPwP/QiyiIRvKtw
AVYBX+Atlddo822UX+/pa1Hld5lfBdMT7+YzVPFYe/CzRVDhApnpsh5Bup6ObIdD
SXNIA+EfSt4lZ9lS/9A+3ck9DxQgV1kfwH5lEQZP9VERdX1YtQQBe0u1jCWeLl6I
NYFyunjHrNZVGakKuaN+JD9ct6L4hrPcrROZpbVAJSBjRdzzO51H5IhjshECKAtq
xZ+IGpo6t4d4TBmBqMIEs2/GtljIVEPNMsZ8n24tr/1zzTm6KIs7GfjRx6V36Ams
O4c5e2WCCZRc7iXC2FVAyAomDYGBFBC+BkM+WTF8UZlogrcUDVwtwDZw9+4iVkEN
cnWRTL4stwxx3hgC90pFzF6TRe76HkXP5//okWew9mzVebVBDrOlrlntDvJ8TQV9
gDG6WBnopKn1Typwitw3qXsefCL9kgk5iT8+6+7B7ji1ffmyqSCJYD/bX4mM/opY
YNO7jGy/WJVNB8XDrNDdj4ovsLkNKlvGIbYu+W8i1H4usfHaJ0k9LTssdrr3gK3j
a87HOVexoJ0pSxIcREKxhIKIiHrDLXidN+SRz4OjT+iVON3wsdewb26mTrYGTVHF
Qk5SLItkwSD7vdzcRkZGmqVGaN9nIgtwLH/cmm5Dcb6M0+YeaI+8x8Dk/YsU8A+7
Y7j2DHxeP9WjlQNyaGQZBT+KXEleoKqHbbJEVr0AxmzOJsVldtjg6jUlPWC+rmUG
ESuj06E65o0MfGQRMiRft+ZlOPUhNqQgnbmdePIzuMIhp71K5xn1CqJLUWboeatA
5litq8eaQQPw2zGbhblnOcEdWSGWo+p5DZVjM+KK8VDV+pnXVe4IrZhvWtHVRc3q
hGZvcysUF+Ms2i+cZP3jBvyTvwFmd7Ta1npgCJcrVCrma5xyLhtaWHdkXygY+T0Q
oEh9CNJEqPb4SMyaDZftDjcjzIOHkGBHDuvQIShzxnXcYahHFXJHLHpZIUm5ovtn
vJ9Yumv3aKyxt7z+K4usRl+KbxuoLPRhE4TdTcRFVQ/yzK9kydiJLdsQl8EG6NDS
kM2oct+qN+xyOVq6/1nKisW0mmaq8d61XuNB7SVVfdT8GIzqBnUy5FoNGM54fKFt
c6WMrX5KB9z6KDxM5Os+PnOsvxMpVxIeWZuf2MaHgZUEXQsWu0btn+idDkjvtsYa
oRd+38sER0p1PWKw63JfNW1dgw3qP7YgVuO4+1TCKGN1XmHoUL2Hca/vsOtztVL7
4EwVrPjTr0EsmutT+C4ftRfGFAbRT2noJJjs+kok7Bn2mZWvz+kwMR2JQ+1sg7t0
dkOtxeAZAqsc5hlHzbUNBmBji+B1ry2nYu9Z7gCkU391W9lOnrkqCmkpb8W5mYRX
l1u9eNwDIDCQc8RKrWBvf5iwue1JWfS0JYU8LXXi7o4ZDG/rxdVowSifDbzPAAlx
DuMqrH/1TuJTsmceTUbJnP0u83CxuCzkwqhPFaUY8x40L01UQoKBXuQRgcCufgF+
LAWduXI1Q28k93CixhbYrdCvHneMHnueOVecc8miI8CiOMiTFVkzIF6A+ShWV19+
XdN4Gx5N22xaDBh9W+AoAwBUpQhp9xX7rVNA3NdJpDhN/YmQL2pRuI1Czb+DSFi1
+Z0XM/XYLvd9EqcoD0vEspCNeRRGXmM6L9o5c2CzQKxVwE6lc2/klBWOOgYA4TAI
ClcL0DOAtvjjW+Sz0BifwFu53DSR97xdG/86ojF8ZT8nnTwfrSQR4wTV4XMehz6P
+ZMiiIYlxkPLqGz9eDc3TeDWNQtJcBrMREiePfC3mc1508gqpH21ebV4rlhIRU2y
FOv/oTdWkQvY95GfKCtYHuKoMb0fmEaTiMJmxPpCMJ0JxNG0QqK2BOROwFazmamr
jnO/qTOEmbn9jBAAINaWm8bYdMUkmEy9sjOsbv7Cw/HGl59mFz1y6WEMhClGV+J7
6QMA+pYDkloTwvM6BTt022QXewtR0nEujP5PCrCrmAuV9XmWeYZHxI25dUYGTUo5
oZTqBNM1EH8Fxbhb6yGONmUlcs5hXcF90/rokRxMIRzTHTrK88PVqpRy5B7s/anS
m1am2tE0etjMSVs8nUuI5iidnzGufdvxyvnFvf/ZV3xN3/bxNVZKDaW1dL0UI4mE
qJfcFNDAUhBUkYZ9TRPOyBcFAefrdXh6ptCFPZO+mmuhj/2z5P1VylyVRAxbwdf9
7G7aexQOpCUpHqzPxxGGni4tzXYegYos/R02jhqKzTs+Z0sjoxkDWJSf49ANzC/O
u39H7BY831BljWZJSZWU1BeduWmshoXsLo8zYhgfqhElzvK1Mid5pzVbFHnGnetu
67biv07zO1ghQp0KyLF0f6uF+fRKn3hltHDeRnVWLN435eQBbz7JfWjHhssfvlR9
4KNys+JyWmXL0mS6NVCEXnrTehMJtkToL/e6iU1PNUdmAnwpojWj097rqG+C9PF8
+qOjfOJps5tAdLJJTdckAV9crDltrfQT1eUxP49Ur/uJA1ka/A/fLwcRQf9ErN5M
iReCTCHH9Tqz3B7sh9shVkFJWD5hEHEa9GJGhtM1K5T1RDM+aDOqi8jL+jXS0L/e
Wmz+YP4Z9iHi3OG2mlIl8hdqiYAk8aCpRjrAOYbQeCxmT6dBhNetDy9R/306riXW
XZIi4lOgFYRaRtdZvC6Ja9yjdwaDhxyC3mpbw0Gn+lwRsnrE/3E/06rDQlFgxcXf
z9V+U9mdeCuuBzrqEaGC8mp1EZk6JMZyJaSbjY+sKZgJUfD64ukUWPfTJfkkinyE
NTE/NzA6OXJjdAFJi1gvsrcFk7Iuv5Qp/XOqrwDg5jge5uPSjvXOiKZcbrK4zxxw
AIa4dK+ti9uBm/cdbQNS8lxgYd571K3RIdjz9OUs1JYfK4ZfXmYC/Y50sQhV057L
T4+msiazRk6kSDMEvpl9PC/60G7RY5792cxS/IrXddDX8BfO3oLPKLH2ad1YF9Ej
lM+EwuNlw2pF+VtdWjYVAIj6upo7MCcacANh0FK4g7ZUUSbdU6qrvxQqmleocP2K
fFp/b1QpwGQkdftLCPXYp1+s1Kx+7mSf2EFsgnfXjh+IPH05gtSsCi4n7PMDTAld
4nofWnz817eAbWftUMdThIjt+Kc0Ypu8tur0EcIkbZBUZbetohRYtPt+7CB1eLDI
k6XikKY7Q+eqhNkO3rhFs1AYaGBFuFaChjAeLBwDwFo8ffw6U0zrqWaOXvzclR8p
sKp1jShDb1ym+WatMDL4j0sF3v7mZBGiDaFITI7muERcb+XOyPYmIRDKneMrmU93
VmHl6KMNpqpofelwMmqXplGpuJByNnn0JXrdZYyRNL+iL9tsFKisjz9QO71oe4//
jOM6ZvxQlmuwMrXeRJjDUnbrScck6mGUXduxuEE/BbsstBjwzLqIUG6WeA5Uc0a3
J4hiywuad+OgFfgVwB7ZWtre7A4p+y0AXGYTWvthZX67RAxYTJacIqVURWD4RmML
p7JQyn22clsz/txIiHbrxyxq0lUr+/hM6N1bWFFmC+Q5aGWNAvGwBd8MK+iBoYBN
DPUGE7Gr3BCP18jQClWjynRlx/1uzcm4PDcrLqY3tCJk8E1679Lgq8+llkzZm8Id
mDjw9IE8lDIdWLfyPu4GLDa0X3joYAxbLJUmpnLRGNmBh8xk6Dw3SHM2K+qtcfdG
NEVQ1gQYIwUnsanzosli9T93Cf6hgXo8Y53/U2NNxHDt2Ca1Ji7/BtTNQZQWNSi7
4kuBPKy1o2DMwlk0qgQJpHwoWimTyKwlJ8ie0rmWiFVfxYIJ97p4gZTD9PN+qK9h
4hp/8Shw0U2XVfybf96/Rr+guXYsNk+cAamsOCV5dy1kw4MWUGFSoC/AV8+f57Fa
fbogTBRv8mSQFRs5LCYk2npviu2kobSP1U4dcvad/rlBjVswLFw0q01O+HrnmoFL
DoHhwQnxfKhkupBRvXoZSCkjNFA9/uUWaycimNLm81ej/PjTR5y34T+miNKaBh/0
b/yuXbJMpesWh8lrFE/mDjdsANMUe0GP+6nPoVhz+tHTDx22uIjlebiw8W9iUjsu
7tRnty7AWycj0RRDR+w4g3SsOpHWBv4JKU4DPt70vtHtacz2bp6GmwaP+n4T/7Ny
BOlnPCN7oNH7mwk8jv/fUACcv0EBO/0vWow8OeF/4Ea7NuAFnDaI+ReMaCCzb7i5
LC/mRGNN2VS9/2hbh7pNfqnpc4Otgz5GGCl+CDSM7maVn+P1dfzzI6Ji/PF96bmP
PqiilMT74sOWn8convXPuleun/oyyrvspGgDpQKus/GYVxx9vPpDnQmUlhKuI82c
SO9RzUkVyIN9n9cMmA3Wu4o+d9dw+Smxre3xWRgQ1vjfoyy6EUYWVIn71L62jI8Q
oYpOybbgqEP7KxFWe+wqrWzblWmGRQFbUqJ91ul8nZ0ccq0H6ZPXOOavEbNJpQUp
CsytKEY45O3sQVI4pBs5ewS70IAz/HSorMVAJd20R+abvCq8QJ9ZVYVhRSoDbasH
irHhG2OTfHtV8t4j4l7JNU2MGVaihgUWU6yQ5ORG/Nd9szCXHvvzDdvAC5MCobrW
8t/H1KFGhQPTCFDxbvJ4U6jWFEhLChDU9snpL7uQh8+hDNwVo1fR2syCboWfnhg8
fUAUJfyVLczTkJhaFWlQFq8UJ9LuR1kRbvC3OT5YsDoEbk40wCqVju0IiAeiSzgW
n0SeNsPg8e6pciwPDeCWbL6bb8KfB4KB+nlC+688w+xCWVxlQRBg5OuO0oP7p0RN
l0+0sYFTE6uZxlY+swi5mjv1za+HATLKN0r6cFFfsrjgBRt4RVVWd125+H4ZLcps
+mk8yIvQah08zoAc5OqO9CnVmccTMsZ0kTGNIElybsYLaHEUCWJew7iKB3FO27DJ
Nwuo/A8u5SSQOhNGzFjCx/WRoyzgUpXfQsHuBVhZVsaOkwbC88Id9snd2zWxwoQJ
Y31GVE4c092d4MmmyTch3qmcStUKG5SyYvki2OE9q0QLOSsEgf1A16eReWYszucR
KXGZFRw72XHp4wOnCVIZUgIFtPJVWyLYrjRq5wqF0Ju4RG6xXvX+vHdJKywuM1bB
VIrlYa7isa6n9hR66NZ3z/w/j4TLNHX5bo374bYGnFI+6d7NJrLHgVW2ggXnFPiO
c/JdSNBvPDgx+LyBLjphkM+OI6MMtcEa5IIKApczt6L+/sMp1GAiXL2bppuSIQUu
/m8Y4epI5xrn5JNj1wWpNCUoO997NEsd9ndz0kPBe1sXhAx0/s+4nv2nVYnK+dYc
P5hPeKO6VRMNY7H96j5gQnqTSlPpBy3JdiTBTRSO8dA69W196gJsljDCLqC2BK8w
/QM8uv2DZMlauICSxmyuiijO/gR41JalEsVvYHrmR6UMABuhx+WhWVSTZbTyciWF
jC0YvjDXIzTrQEwn9mC8rnADe3FaSJROfaKwSUCNu+n7CMvkP+xCg+fKaJSOgyrP
3m4GyX5AyG5noads2TOkJxuMwIBVc72nDdVKmNocTiBpbYKkvS5EPNT7nCGSsRIk
2xjKiEwT/2aF6mPaEzViuI+vjD/9h9ZtN/A53Cwm3S7nGeuRbvA6WeqEH9UivDwR
nw6P/cQlPlxYv77KPVMauHLQY69kIFN0UtxMbCTbebijufdZ+aZQIkYHquDoz1MP
U/q81v7cGmgkNM5NWCBO7PBwdNguQkknkb9J3d/KYU/Qvc7nvPp6ymVsh3ZXZQuz
STYiNx86IArVjTsU3mjdLUipEY6r+xQeCOxJRM7WfizpEYHxjQQBp21hulXGvmuq
qobpghiX5snWwWpytisWXTQlzdr9ASXldEystFlaVULzMpqsb4PAbl147CojNNAk
ujmmnKk8oB38kjGrVceeLLd3Q6Qa6qrZRewUQ1Ti46V/5SyJg5//HF3lb/47wnvT
CLTLvlYPs2vIkp+pBLGjRWwpXlNzFFfssXw1bF2b3w8lmfKBMB3zfxmk8PDevChk
QFkAFhN5uDYALzKrypYz+UCmgzbafYrFbfbirscPend+p80YLqUBXzmDo3vxMqJn
E9+Ku0ajq0OgOIU4ieaN2Fu8YM8Tx86ro0FE9ZZzegtXsKnXbCNZtYCL3RKVvAjC
DlGV6GZh6PWMd2VX6NWv0huTq5T5aODYbQpUXNE5l6I6zBeecx4OWZHXRi3NvX8G
0UkbYFgBn+70tpxqQct183rBWd+CtMC7lNOmooQHDrotljSiiz8YHtiUQn8pnlgy
VoNKU9QcEqxT/AqNn9gOJEAQZec1dapmCW3eARCKRtJvNgkUYRgrPKZttqsQtaTB
WF6z4PKGoSwxr2YFxhARVwB+nqgmViFgZSD1SpKzFIT47wFjXAzmuUKdW58qNNVM
PFa+Ws/utndgOEKTA5YHxWB6pBd5/WEvN7Fv9tZ8xRroq3rMUJCWPCgcFK8fVSHw
zlZfMC0XdRPEbqfDjNEMhxsbvybUs3aUBYyDg8si9fHEwy5ZKH6eK6bfy2ZTuSQ6
46HOh2WMZjf9IB0BSb66FDs+lHTU6T9GDi1gT+5XgpUP4o6o1tuM/TbqwWtNIVZy
O2SQLhoZvu89Fw5ZXFxOxtANVRwNaHe0DeAvZKe4aP87hNP7ssQio+9sm3z+rtlj
IrsTRdOMEXn9h86f7pvspDvOsg/x7+x8qdouuh4q0aznibbyKhIPSiEP/8rZOGOo
J1k+fwuyYbyDVNF5Nm/3BMpBQCPI/S/fv3up1DOsB9UdejFS7wdh4LkVM/Q3Kye7
wlycnVXcItvZ1dWy4cepa5U9pwkWPJCyrTVIFbn1mQ8feRYbt+mQJqWfweJvJmUW
Z22dl2a0gAp6tny317dZwDEv40olTmfbNRy52sUidqkjCGpkKaj1bXS4ENHDMXAr
7d6GvHQlny7n7PKihemLftxJI5tBfWBIHCR7pfItd4OETjJKvstHZNYBwI6053/9
RXBXRu+F7N1UzFNXJUeutjWYqGgeROWEzjCQKYMyqh+y4I2r9QfZmzfRsf0g3zFM
S7O2Hn3GsBFFe0yOFVvL+0U8XKOfQ94c98wZWqBxsr7y9VsuyDQj4QMKHw/OTrm5
PEBIMAay5+ACaDEcvxFZX6KCM5MP0JuSsl+FTmUj8plTR8XMjl0L4aXMQpJbIEIn
hep8f4GiEkiRZ6WW7eXbbRc3rGljtmTefI84KiB19IkCxMkJ4oSLNlZz2KnnffCE
mhRubJDXzD6oHxGvbo9f+kfddFQ5Exqmif17nlGBIwJgvEV39KUeZWGMiKGuErdo
vta6uXY1XV7UFiahHRcuBoVJi5huxgQP6qWwVIXaEqY1Fk18c0GmC60Lp7IWY/R/
zvVGCr0R4Q3S31D9JejTNAZHXRC82d3Fq9bxSc07sAMa0UVKS2UzV3/A6UdvOQV+
PLiWvTIozrjaQC2ZlBv3RT8+9bjRV0W48akQI5bPloLndufIvbCk5apK5T3ZBaAl
/SDoG2iJk1w7TNpvJ8H/WAm93/F8HscpldjAkWkHX7vDXSh/BzfmDblzcZMtWtWl
LWfbzQuTlxuZPuQC7LZ7R84uZ/opmg2Rl/BG+SUC6MvXS50OcQDvFhMcjzGs4Pfc
W+c2Olldvts40ynih/OgviqMF3q9LzxiQny0zigClkm3w4kWrd3BlQksdgEBgTP3
ZpAIAI9Z/tx5Rh/D21j6d9ybQcDR6fSYXwQbH92RVEsnNvKceRFVa+2uQR5ks86M
qoAsD6X4AACPAcHnnmhPOh4cyq0VL43ZbSITv8ewXk5q3/Q52FN0/0fSoVVCBk9s
aLSbJTbgbxvmgVaKJC3bgSFna1F0vcGZq6FDqVdPT8WlKjwbAUPqaeJDmCz494X9
FFCf4suc7TtIA2zbwb+0pYDOE8MMI5p/qgJgPh2kjfZstAS/gYzV4LwM9QWP635t
IKWDBasg8ENN6Ypt8YLu0IpDkpcCpwFw+QJ0nF2BbdaqduLzLLQ5t7sTOaLX/YuA
gDQ1gOVD0nD48O/f7lWQsoOdJD7emROX8ab92E0pS39yWX91NKvUKUfC7FpO5wRo
bEkhK+JqLTH5HRrn1lCvtaS8C6AbVSu8q31dRiW/KFcPuqwmARA2HtRULkkJ1xGP
vkM9BNhM0e09sQelXzaKBV9x8QB3yjy8uUIZAXi7FZ2gbAxgVaFbu5tNjLhvIHF8
FtTaB/JVDaQPxvF1Q0gJ2IdmwSR75qKDsUbYvK3kzMMy1RaUpPgtThzH88RmCAA0
g6vQby0XAps+R3g4cTq9iZQ4VWSV9eLiqgfF0TVngrMJW+CPtXuSf8G3YMkD5eau
0wMfNRBTiRqzfKvgopR91yW5YcjxYWUOjeFr91YoF5ldRnW9nRkNo46DSWadbKsl
ut3KqqYvDzubAUUuIkBaN7GpItQAZa9o9ChRmjQPGPnJ4U2mwhbr0NAgxm1JEBiE
lLVDG/k20eBq0vuHuUVJcV7QIXcp1L0HfjHQ26EirqVUoM+dL9bAB+jGZKFGgtNV
KPf3S3/h4KjjXcsCcs1UIDeHKrwdYvx3Q8Vow8eBUBlI1sWqMbIajngmtxR9BDX4
D+CJT4XpfN8u7HIbzXcYtVECQjOgeWdtCPnqfqKbz5OKXdFLEGpGNBcwDm23dCEi
uqJqG4Ym0pjZX/V0JTYySlWt6CE6+6oxsWfRKLT8e+vebToT0JlhQv3aIdNulTNv
W6Lzd9uyplZzVz25X8S6v2wgDx+ebhQvphl+TONbxQpfA+xaefT+k1bDNdY5qF+b
lT6GDEFLtJrFHms/rGSWpENSPIJ+4RfCywkRrCrOv0sWoF3vq8yl9+dySexU4ePG
MK0VASCpe9TabL2bChJx1p7ngOnSJyx2x0HjcrY7yx9UJzXXVQSw8KlRjpgB/DMz
MSngLgUWlgoeLTcQY9X5Qzkr9Rhn0c6KqrnyvYuKd1zQ0aJ1pYcS4QXl7BHeWnlo
mNYV/36fmw/mlkWEHtWPnMkpfEPCeFFqrbsEcna0LVIZkTvdxms+4XCDbBxhOXKt
YBFfVejizXBi+GLI81pt4ah+zrpyQT21gP0I+E+D8a/hSN9iTNHOTw635FDtRWok
d8X9CNsLAgbc0xOF3m+TDjBEi+76/2w318VYzSr+n9A2zdzo8l5wRTmd2b/Tlura
3dfWm1O3BxVk2K2I+2pfg+Ssabes7zAc9XdDIE2de3I3nvslo2uhgfxE9xvslHj2
HZ6R5EmBIhkEr2riixE6ehFLWAfWqWu9KFLdxDIqJJCHfoArgMUoGWC/8BSdrhVO
1JydYstoDppcrzsjUjf7n1WhE7afw43DzMvWnlR7V3x+i90zs1Tp8FERv+Ijy32a
icjLE7cr5BnJV+R9rbpcRNldhVOSAPwgnIyGLVTMzKss/qNk9kGxg2pCR2RtGrWJ
ZaCHOH8YnIsNQVTyeoJ1ijuJtWqZ5Et2ie2xBo8surbtd2MCcbmnzplWDPIRiDjs
fQRL6yIhW2OHuujHPaONKEDQ6TipOrDfRr7BSXaNGBXoFnHw3VTVTdy5ss4NCC6q
EOy/dQnon3+h+KIrTwmcX1TmRT+zY01zyFDG4L9FUrb690sS1NBVk5NiA54Q4sFd
TUSJI7gFUblOVRT3mlEK4RQVy0L+r9YXMXWrC7yX0r/npmb2HgD4YTLu4/Nu0U1N
R9KeuFPB5uBYqCl0SiGp5R1+/eJuZ/vFMZxl0KycF4EFFcK8YNbMu8rYKMI8dGr4
57kSqgDyO9vu1YzJqhy1dStSC8ojiS8Vjyg6K7ijynE45z99TLEzFyGSt0OfFEa1
go/unBfqDbgSkdp41qfoRY1LIdXhjNnw0eix7p9NXnocdktkKeT8UKUiQ//1o+tO
1HPmpO4g3SuaXVjQbZkIQJy6z+0rgfQrqKzibOGwUKHPSeuu04uUPzWi0YuPab3S
1bIo/lh4GBkbDXTYofLNADBG8fPyKBth5yl/gH1HHM0eZB8QY6iAmLSv80uYOVpM
ev8+YG6MxE5aeF5T5VE1EQ6dxFEFAKab8/qxz94L3y/QcgywcyuAgJhtAjaKS3ix
o3DoSb5VsW2ycDDb2/1/xEPIL/1M/Gop/dMEduESqIk84HBSDT1vrAujUkRZIWCa
TBVh0V8WP8vuwt/McQ5AW756mmizqSbByQOr1XWlQq/s9yYwDmn0d4c9ZRe9BxlW
axZg0vNhoB4bMRr12jWI5WkChOd0CpzNm/g1QZwzj0EOKlgJsNewL1ozC5hkA+tP
zxLGgCwUOkRaHR4rkWuCPrqp/VSmZTadoPFA+hhULGLTrU43h7wIb/zX2bsEQF5m
pPtIL/HJGLjAe7PpfS6Rl4f3VO3RZmXGkoBxtRCIlbAlWqsc6LcABaeYCuGGbn++
umDnimSNV7dbmjreZefBhNj51sDDFulflzkMtdp4jXJCYy+BbKFLXi/nqU3TCX0F
3T+QGx1RuzqLhhBhVQes4Goue2F8HJvhAQQXGucY+LyBRdqO/7A0v6GNtF6czVqA
urS2R/zs22QVaI50rZT5FvUF2proFQMzxgEonE1h1lGLYhjHkEIyswP7n+RqbwzA
bJBE4tWTBiJS3HV+wJnFow0IFlAW4PoSUfIgtFEcCWQ0BxsrItZ3k6RRf19q1Bq+
kDC/FV+lpnexCXgN4Rrd9LqP5Shiivs//OAeONkrdXlqmmZXMNdltRlp9RTlxejp
iUA4PuJmUknK4vVpEswzSp5Z25+nTeeRARezlDpahld0TikY546dB+4AdZ7GUksE
Uiyps1HjMIhrzJ7bQumf4ZRuuN0uA7IwsWT55uEC+lH3mqG1/90oSr9eZ44XaWts
Kgq1S5R8vuErK92pqW2p4XbX3md9Y2VdaD/Fwve+Ho0tTdAF1dFcUBKlSgetRj49
UyYmMnt6GV/ImtU3apgoDSLtPhloEUDT/F7tPwllk7XwAzSACJdZReCZrOwMB1LP
h9lfbf3VbE7HcS3mQ3AxSSIHTSyAX7pkaWvHq/HrqN9Oj8iNj045fQe+SDSwLxcy
VCuaoV8MFJUQQsOQABh8j6/65CpszHkitc2lgiwFcJuRsE23O/FYXZgiT19RGjqs
TJahdtz28LSEluP67v7ar1Qw9ueMyF3vg5lDnwGH75ib+JMjeF7AV4UuOde+Mbkw
s6dJTzv6rd7YEDFpdPO/9H+T32e45UdFJz/kyR2DIvYbBYNIFOfdaupmNfa1DPHD
ANqUK/+41ounIRQZTLNzohBteoeQoTAAHGtsH1qVE6h5qoQXQQeS4urk8JkUOtgH
j3CTmjSSJ0lJyMnTeIfuSbD6wFDWDPBsvhOMVpdnyE55f+Psjl8WOaRTxjt0S85F
otzXx+Dk1LN9+jrBGdBGI2v/iC1ohFUImxB62O8qVmSOxOJLaKlRZW7fwVneSq9N
5uVf9C0S4JpxOmufvQe1OdKztbe+gw9BztaYNkypqMgJS7brdUIdQdPuxGO72WR/
iiUMktFO4Pp62LSq3WJxF259VqqIDGI5thWRcTGEbP4N3Ai/oQDVqRBqVcWPOIRD
7gQf5ditUA59A5TxitFCE9C04gz5X4KrlQ98y3x/vStCeuC/gJbzL3Nk5fXqnKSD
Qq3C+Lqsl2rUF3dPFi8XnJ/rLBEeScWBFR3Dvry2JpQG2S3dbFjwZahEtldN+6eX
jFQTkXNkyKCUH03DvTLX4n2XSeUpHC2p0xmklU24IhNvalhOvQ7J6Q/1dnz1qUcl
GdZiETsLehXtkatdl0mh3RLDwN70kfAbnzmhnWTr00NzADGeg8wlyZo2Ojj19saC
Bis48g//CvN9OlXh7s34fsljeFmjdiKqurWQyY5FQyYmmgopwxvAFl2O/K+IbcD+
sPq9AYsL7JL80VLLQdXt/Pner5py+0qIucGxws4473buXo2zoPezzKGO+Ba5j/Qg
fM8L1vK6egSis5f2JowA1rqvlWRZtVryMZWfoI7KeE3+m1p7jFblZHYlYuo+BfA4
6RER4A397YQhjzc4YP5NuMTPM2YGWZ77W/lfgymT+kAe0LKgDLzEcdDFsjGKrmnF
dX+QD80qeDWNWV1EZXRfj3dFyenlpIw9iHSUXU2CYYSSJBG4GUS1e/zd3+YawSde
gNrKxur66ibUJk6cqRSMruPcAL0L9yod1FWxzPIkaVvfLEgIJnZDl07TBXo6NFNi
RYRitSQZW2m+t2woJZQRkg2g9GsykwyoTcm9n9KllTxTOYjk74nwpTgmlYT3Bnpn
rPecrgenMt99rEWFKr9WcJdS9V/K1CU14aLxOBfNx433AG4lWpwCoMBCRijFwDpf
RX3f1FFDV1+KiF7y19k5rOGTeKEPkOaQFkOderGAIcZrldwfbAcDpKtagbVrinNh
ZLHywckQyI+BRS2hxPG+nl93+mxE8rhP43ZYFrVLwTr6FT5DEnwR0rWyaSHovoSA
Jksv5VvpP8HJxSnW/h8RJ1jaF2ExQ+A9fw7Jg3ebrB1pfDP3Duk4VbJSGXxsNWA3
ZteSaXuy5DAhvei5MM1OIi9cUMUU9MnK+mM2BJamG0wehGmzUQlQQWwGDoJzuB6M
RKVxAZKq8FD+QLf0cYYj4P0KkPoyXpZmyo5YLbtgPHGBub9LBLf2rwCjer/o41xy
+klobsUXs2rOaQpPTrBJON0a99gGsS8x/pTsqTV/TCOvSYw5hLsOIpjJUbRzF6Xc
/Bkx1xLSrx33/KglU1Dt0TcG/WKXmn7GAaY+vA/51bya97YqsX74OU4LmNKBkC4K
bEHX8OZWWmNOso7sRAikuvRFRNBoWOqrP18kSQ/gl6y5o112yoeYsUYQBT43nG0B
Oj5jJ9/YMfwEkemQMBdwT6ii4nBhvN1UgPDiP3nHwnXIRIrpo42EPhA+HYy0Pz/Z
SQmb/Rq8EVUm1t34KxB8RmcYP+09I8nSz10wXmtGh/x5XIYRRPAnFkQZ0EhPzqIt
Oq1U/Z4lBWnJmyZTSN9mCoXjg3gFrPChnWZtZyLFm2yUCyIZUuX1FIUhNz3pNY8r
gqmDjsyVCiGQTmHiHnetzgBWHCuocVaEuU7f5F9zY950w4chREiyfEhsOvpJVytg
kr81Uxl6OsSt+LgIBejnx+wZDPhPEYnHjPq7znUbdi3odpGXGQoUeT48S7C5C6Aa
FZe7TTFr6IZtUn+C95Jnu2kgY3n9a9ZyVks42cl8LhJ4rKZqzE6KebaR0+Q1XG5c
GsyoheLsQ1ngVYjk9B6O3sbfjQyyE6Mvh4KA14VvBrabekMCXgNGkYC3K9e88CWu
WejqMeGnX+eMOhy0Bpvwi96lDsgOwgT3Cts2Pj2ITSyFtt+jfH+uPFFoYyjunDdu
WgT4+kiktrk+YnSxAlZtNgi4HIapdRGQbAgjNF9Plkb/Vgzu4p46pzXY3lR02oZP
qjJ1LishuG5VmiK0L53O8ho29k9mAg9Yz7KiNUAd7MSfe2wAhyBwehQ31IqOWLeS
PvY2DNjF4i/sgusjpIJrbXaGzkoA7b/vq+YprCJRG4Mi8qNidsyxSJ7k4biqhijV
zZmtPsl9BSRboQumdpfGtBEWlYo0bj6W7Nchy+bTVRsPiYzR62CG33bZE7P4RX9W
ZMeCxAnDmhe9RcSJzIKFY5+Eri9UJ8+QrbhhVl+UtCZSt5D+4LsTmz7c8jiqRGYG
eHdTGI+5HAu8tlI4CNPeHEzfZXKwpbwQCbv8TIZ+X63CMLa1oVGDCCbvTaLZW/5O
InATQzyBbkyPFGIsEmGxSz06ObFLKcl9BTkbktFTukZ475k6Ec3uxDVdKvHA72gx
MhGyM+4/1qACTc7v9s1x/rY5qJo85MoyhHWE3eMiGt9ws9Mzb5e8VSY05wxjLzYN
BKNqkji22Das6QmGXxMUBCQL5m6iKOiE8JoN9sx8EOgXtFLKnwKvvfpP0XDwxkg5
60Mj+MRPv+FNG8gjiUz1LXghg9CDc/qxJXntkF5yZj0fRHCkFOVTOccfHUE/BGIH
SwYygXOhXy8oErWT+upW0JM77pw+lkqlsXLfDKhCekbSSeWR4vZ5fCVdHlI4h//R
l81e7vzBmhv/LL3ZniSiQOz8dFJ4CVSywCisCJUVdtxgena7saS9Op6axsgyJB3n
weKRQz1/G0C8nABmSkcDm0Vmmg4P5K5ft4p1TdebnNvqsk8IJO70V/p7cGj/uwTd
pFWLQFWNqNhBeu6StNq0vAHKyaT9YK2PgXw+UjnqVC4pPbUCjw6zwBfQI9AUib1K
SVzIxInUz1UdSXYc5Sw1JmAknDwU8EaW3VSY0U+VL1mlMUMp2dTNlxqGCsn0vVwL
+y/msvA9ztGsOghHU7ChJdDryw4NVdU8rKOqi4nFPeZIiBiW373MnbCy3vJSxKyd
7qg5cJ3RJ1khfajsajHHrDdKb9r7ccyCcRnX2Kj3kcxgLMzxtjS4zbF7DECbZMJN
VT5501nq31bKyjyUy8c4kF2EDSZMjde4SLsWlPjWP+lD8aGw5eDyMXFIl7lxh3Fs
XT08sjf5tIlwwZRjHPqNDoXnXpUEzylh879kQ7b30aHcaTUBCTqH1yjV3dWg0Cs5
bR7jAJqy27vzhHAZS9RvUdYxwNi1qpJFAIQ/hlM1PMhSCKfYzhNbv9jyLuhB7sXd
6sVGzNMPIKWM6UlUJVRNHVEtybFVM/fFESFIrTOU8fCF++RygN06M7HdwXtjC/Ej
OmY1D3U2KdVgy4NBI4kU0YYH+QJycxvymGJdSX8ZEuYDpxi8O1yohVd5sjwwBMmO
u5BcwzKHMNPM+3vCK0J0oh402odhpNx0SqBu9lTvPOuHqbctMIsdhEocwKQp+bCL
eo60FzmrU+W/5WPdBEKaVH3ugzv3wchHZecfGURXETbh8rroQExVrnrSTzcNHOLj
v1CGFBTGRAf4W/rTtvBqoQq/G4ShaYKlccgxFl4BUkd/07eswrzHZkiPfGa6ZodJ
1I10w1fVRpkrLPTbruuGsBdTu9OnRqh4aJo1dkgctI1nz2bPvWkV52o2EA9iphIN
KaMu0C485tIqIIURN7QEKvr8ZX8tCXjiIQ0KDOiXNL57bePHfLyB5o6THSlUGZaP
4htPQ4p0TsKYcQhOk5uzrH1ViK1WWMICFgB0835oTvKnxxEMqc9GV+X90/2rHsw3
BOjHivmN7eyWz7Q4sdZ85leH+yR6AUGb2aLH9EBMF5iyPDhcY9hThM8sgStUVe1X
MFY9fppcmKay/hY0CzFfONK9UFhkFYrwgYXF1TzOHjPzQqvE3MaARQ4Mm4713XsQ
/95yuDrDlT8MV9VsTdJWmQiPp6+OK4qKd088lyqzuX5nrssNNI6G9QKhLk+PDymE
jyv9HAJ5sv+1JPJalYGy7WaaMAAtdWSULfwnZUEjHB9pCQs7UxelVBVOPEgJ1BqA
SMUAQYvefRol+a59hhIz+Lr8xv0OYTP9DWqxUmkv3StNSa7fQR2OCUUelTFuF6g3
eJSYXPQT/S3nnnJnAlY3h32AWW8OMBfixHfaV/hwQ/lQy/3FEHEE6VU6P8U6c3dN
WTAcDktohOwL1cZ/abPDCf06S07/uuiobwspx5ikirvoXAxb6N7hpFw9lgZlFqn5
tvX+wS52tIoOz3qfcJ5oSPOQqPnzIgQm2KMreBTLlze+rP4KUL5N611q3CyUogr7
QySVgMoQPR7FtgNp66q9HsKmTkRqYhv10IpJEQqu45Oo4qke7rd3lGfa3SF3B6+u
utHsGjp6xC8XZ3yXQ9UeWZgCVkJgpZPjl2r0kZ/k3enp6Wjfwuow0TEk6iosC2H+
Ir5JsDzEq6JXr80JHI6XaoSa25OUo4EaRJuqp8qSY9OS3+XiUEGEcu4SMfox9T/g
gFMtUR4WJztejAZEoCrQWpRtUYxC+bx75KX/qY0BH/glBT4Mpnk1EHJ+0DTF5Nsi
mZRV+d/1gGrbgioSHOmS6NJu8KJPUKyFc/2jfpRxV9QNfZrR45oqkHAXi+oen/q4
lZEfmez5N7hi0Kn695sI083IvzR2pDj5euClE4j0EWxa9XwAoj2jlLEx9bK4yaLU
lKD0b23M6uZuo/nwXbKwr0HT/fOZFaXLo2WZutG5XyU+Hqm0zfSJBEDGcGpT9/iz
1YT+ZNAE90g02mAaOakGsLg34gSX5AyGG7nUTVwCJloCyd33lFImNfdl/gN7KPx+
Dsfdyvy5eGcB+8+HSQns3ovPTl2D2CFASx9TARi3Vj4lLSP9Gp0NQad32QTJrY7H
96fTiJC8lpu0bElYl3RUGVu17XdcGreZAw6PAeMCsuBTQvxIcw0AgLAqh4BOefNm
wTpx0Dv/OXrYPb2A1WpP75Sx/A/nIHsVlbt060QlbLi7D0bzu03k2CZ6bv3s513+
OGNV3wAB+eHtswr/DPf+y5SJCeP7dx93X66DmPPMX+eEf5HcVM3xvT66cvW/4gBw
Mz/pnxxuxICPJ7xcHDC3SUXqWrMkhBOI0iijqlx/XG5j7ihd6AkxMb8+5OPrt3Dm
ssmV2TxDrgJYB0o/WbdM1hRCFu5Q0XUrRlQfF9CNlH2Vw6HXmUDDRa/5otC0sLmX
MTn+QnXxs+CHsmYPOact5Mjqk1AdzkGiB6Q3fTvBX2VAvvvDWWqj9DgndJRDh58D
nWS5HwdWas6mt6NgJLceRffZFd6RwQNdNlYzm+bl615IX2gY3rim536b/EqXn1Rx
m+LytEcTPHCFhFAsqyux1M4seMUIo30YRPkztIGXE67jYL+4uLDQ3tHaOxZMpsMa
SpEJx0X1TuJbc21Hr8KzD4eMkMiJGA7InNsol1idrXHnq9ycJsd1yW5N9jHTudGf
O1r4sQoYl6c49xw0G/qs287azEoeT4VxS7tVj//P4HV10vSxS/s7MudHOsl69Xzw
eqwjj/Z6OyA+hXCfDdrnkTvV34BV5BFLcqxqFwO2tZQqqjaVhloKvrKobD63X/on
RGh+OEJiY8rAw180Sbz7YDnJmuvkOHOxx97CUOyb9mikzNwfxXCxH5Ttg+dvDOXV
Tb4Np/52/MSN+rLyZq3tPemLfB3rH2LFOFpYZ9jY779DP+Y6VDlCjDtBBDrO/b9o
7T2w9frlvOHJl1/6twopj1u3vl8TQSYQP8RiwvXJOTz4vHu8M0zMCVUlKADexSsV
pt5VgTnuOizQRaCTOT0q+WkRBiIJnjAX2SQZI9lSb7dm3zH8yvN2VUnRgp4z364M
gtsRYDQxWE9dFsLQlNEE1lw7NztnIEot6kkOzVJPRuz04dOd6tSoVg5cYI6FgOC1
L+YSiTOio75n8+v76D4qNiMt3QLbxTfdg748+KWx2OUbcBOjUDDONTAehWRTx1kx
2/kxZRXORdFj0WXB/b0tJB2E6S/i73dn3ayW60MD60DHVbqVsA8YGpLC1RRGBQOM
xNmVPRDj81BIQNevVdu4ZtTIpF9uFrQkc/yqnx2n27zJNnsJPbJXyy3QfK+UiVRf
YQ5EVkz8LYlljMD8Quwt7Q+lZteWYSkPezdhTUePmRH/02C9QY0qwHJQkThL8Lr3
COxPiplNoQs8MMymeuV4YvaANkmrMDU3rwuteu5xDhFmDWnH4FOtwyyzfCgHnxQM
lzT/loxu0idcFangzJ7ce2mz/CoMwyHdD30ZZCtwu8oPRjvpPd2TNQPlQ2D27JgP
RZ4+XuX/xZgxLD33KT2D4tpRcPUkrFKScdX5QpLKOurzP7BogIxJ5fXLwz+ZcvQE
mVbP/yhyu8fiMPAZS7joWWvlfnPKLrNLc3dM7s1VlAkaQzHQaqaQJ8DvLfQR4+nJ
ON/p5OhNViuHfkbso+qjggWHLJitoaNiayw+9xcyaQiw3x+TBSfm1XJ6Wt6podcU
0FJBXHuaWeSYTMJESY9bYZf+sefxCpNldCDyLFLV5KvuMh1xDTKdmtRaDJqE58JU
M5SNNxKFpA5WwdzeGWOl2Gdya7G7bSyYYXALD7ONaRTpFkrkhJTqemoIh40k9ynt
4nbXQWnPmxf8Ua14XA9YegHG1mi1gVkSRVLLI9elR52NBahrg5jgw7OQ3+UZasDu
vZbZtWfnKPBshTIRx9kk/jM1pyBFR2TRu72r0TKUzAjbg1Dbt81JDlBCJS9SdV+q
2hJOCviZzrwDtLueE45QaKl+Lm/S8WJ8mKhfxTHpCCPBh+/TQ85FxOozW07Ky0UE
SkzxMd+H2I6GkF18WlPKk36tUvWiMwGSCTfQqK7/+/kqN1KlPuMskDr0hcS+9McO
HAJzEwskltHQv2l8fU2f5izQbIDC4NDqVjBZkOFEpzBh+rcNBDzmA7yRmPyIOqYU
po/vyrmqx1FHIOrzh+mIN7THTVrZ6u4FsYp7PdAHmb/ku93O1RquKjyH7gnFdexa
2BCWwQ3/yvAzwxXx4S5sOTSHjAX47vvCA0RuV3Lh94WPplmcVslyaM5MEtIIx466
y5C0lk8U2JXT9GUR2Du/mEnERkzmQK5z7EOY8faYii8eVRLV0xBKGt6MNmc6CtL6
49N3qMf2ysjOdxgo6lMrzYtpycCHwld4mST32e8aZAUZTrJhWAglRis7QS/sPR33
YYmMum7JNPsaLKtJ1URM/iEuaKlww1ESwtwloW/ziqP3GApCJ1FPuj+9/ga3a3zN
VnBHYdU7Jk/ORMC/Ux4DJua56o0AQgRQRAGfRN9SQdlkD9rNvGu+FLP1q8GYjruO
cRpEpq4G15Qp8vxsCKgxZmaRAtESzcCldcwyT5G8Ic0SyJhq2PtpYQwQoieP2XUp
UB1sRQ+G2EVACAdtkNrt57VFLpdGQU4IfAUffmUVbWZ1nxiBB+iKRUp3w+iqDJza
RcrYcDIq7NtCkm8lx+OHok1mqoPp7qmMGb8UvTBweTpXEE+1TOsn3Fw+qB3k5PdU
uNlySNrdCjetNt/QY7VLEnuO7+PN3ihawFsb6GeJA3MXxukETxcHkFy2Qqbqj3kF
sccVDkfQd8OCJJJ7HRO+glxK6B0r6pcWL7Mbpy6N/WC6EL1gp6P5EAQjQc1Gt55N
KToB+W1HT32lOoqCYts9r5+Nasv4jW/o5uIrPy06PMYyjlC3V0GpvZIF5Flvg/Vp
AulmFb9QoQbw20/cD6aktbdwTYaLxREknCtggsFHrk3E6+iU/PMfILCLSB/F1wNd
Zud7rOy4MkzhC9XqAggnlcmd10HGUclKykS8qNdjA0H//qC4+tnYqNqFlnVTr9kg
WqbbvSFdgpMn6Xg4iWDBAJpNUQaL+dmTeCq+A9MBwJxRwIeZRHR3OE984S67PuAh
NCYSfziQiFINIKBVF46YSzeb2D7WdccpQajPucf2J1eUldR/M9Ej1dnivCiNWiwS
sVm8sRKrZVcHkd14WNYey4nAsn53rpPi6iNmBEk2gDo8GT0nwsKHX8f+oWQpmxtj
i1L+BjqRJ27LXJUHkf+Wl4qU7ipHxO+sbk0+CiQJEGiOctz9FJWLwxIuqhbjefD4
uGKZ651NunOi5Uanjid3QxsV+fN1Qez/N1U93ceCZpv5L8wXC/IXx2u2lkcVsXN6
xFZnFhiOwLAzVrt526flk6doUbEb37Ktq5f+WkzmSfn7JwSjzDZduUtVOLUXS1Bu
5jkVY3bzEQYrYLGAo6p8AlAjuJGg0lOVJykSeXC9Luvrts7hjIFfSCiguA8pZ6D/
6HV+qsjJinWOLkmDipA96tP0qNxX7pRdDV5eVI7oDmOXxfLjnrNbaLZbXpQG8bEU
gu3/g+cM0c8/xvPvtdx4f+SPH/57jFchjORHVOQ5EmAj4wyUyLJZTExAoMIIp/za
4PccyWdwyYNE302XOfMRY9aocohIvc1UPsF23ydAeSZgBD0DQE8ufWXzsonshtSG
1mkFLmcypJrDpikZoUmXZuMjvWj5xi89xuUYRB+AhUQAUHeJM9P/90T5pzYdn0rH
G1xytmDN8ZiJEYCbt3g30y4PwASjn8XAMdNZhjEddHQ7zJ6OcftFcXyC2lBXG56X
SF5INTx7e7NvP+fjHDbOKjvuUCweDJUleHPEJkrDUZxKSukRXu5uHwInT0sVffGs
FwTzKFUmumiw6jXRrKrqqKoyMS2Z+H2x9Ll2QP0seFVC9XodeaYKon5Jg44pjF9c
Z23H6rC+L2k05TFtzPG71u6vDlOYoQRADvkAGpUZBP+lGSEKo9Co/KY96vWG4tOb
+zEr0k/ij7QsRdBdXEsWi38uYQUB4z1UCQzx5KPsuaCmPxFbRhxkVh9HhuM5xVTS
nRLxI5zg+JNUA6h8l59RnPZDC+gE0xZaodbZFwshJXKMRWi95+UlyQPLv3jE4Xo6
UE/GAttpQDswuv8rgo8Xvq9lV+NlBDrWr4Vvck2/fLa1Vnrrj67J9b7n0D4xv9+c
YA6yo12FHewhGw0kmGuu+GxsVG8JptqU0DrFp5Xja/c=
//pragma protect end_data_block
//pragma protect digest_block
aC1htZpt/jwYGvjZoyFp+CwWxKE=
//pragma protect end_digest_block
//pragma protect end_protected
