// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
+yIeUZ1P4MYePLdeYi/rJN2o3AQw0Z/VxwMP3MnY2yEt7gtmbyeRB1DT/0gtQUuF
f9iNOpjtU5JSXI4+UHEKPG7o6KvnNvtAQDOcT38SZBttINVNMdqZ70PoKXPf47UV
Mg5kNqN9gRbn5Yj5+PxVXjrYXjc2Zhp1AvD2qqOQsWKhExhf3QVaCA==
//pragma protect end_key_block
//pragma protect digest_block
JJA1gdPBM4tEL689ZRBYxwxSWRo=
//pragma protect end_digest_block
//pragma protect data_block
pbaTlOo9naWh2w0ulZLtdE+7YHro26HOlsh1I/vj7EOncZq16yM8ptuSthz/lXpC
rAUSYZrEORm8SFu5ZJYAO80Iscq9H66h4cyjEpYp+yKOYaa/Cd1yyZW6FLTosDpf
gOCcFouZl/cUTtlCIz4efWnEjG6ExCXDlydxqWWAGbVoHl6a2yelCFgCcovyUwdS
DFod45d8U+QwDsjFzn+aOJDhnxCr+4CJ25EJcP5wfSKbeN7u96tkxebSzdyxcERp
ckWE4cpJWbUiVI1cwHfS+Hho+JWU6umaArLCdRoNYAnrrRiZ1cDSF3NZatFLJ/9M
FyyEnf7rE8NfEB9XNXHkw+Wb4XCEbJO5xNy01jMOqwOFt48pPDV7ef81Qjhh9gqb
8fSkz5A0/6hwQBtH5jzEiwFsvm/SYLfe55TXMpRokuTlXY90/HSqmedkaMkbCykn
7XzUYwqiF2LhJHrs0dS4PxlJc+lEz0i+r+Fep3Iv9KRqWlBDbRCykvv+VdO0KBkV
D3oN0cMGPIXlIset7CuwX0Oeoxp+OvkmZw61/ZrhYX42f8GRMeUiv2/bAi8geePY
kM9281KFg8I+MWw/5qcLtCreTR8D17iGR1oyz0a//9q4dZgp9iMCy71eAV4mm/no
zbavjnGZtEi2S3gvn3pYfGg3cnPBpQLXYxoZS4Zac6oKDoVUMJGsfXyglU/0IDRS
GmNyXOa7YWaGC0/phs+LJljmtExJKvPMKBdyhRhCKuG9Eyyo80wmPQ2uhghsnVzB
J51GgWt6kAzZbHqNPZ/BuknCNmygLcbrHxOm4C4itKwr8hkNbQM3bLPxrLhVolQu
ucaQx1BEvpjX7At8Q2PU1Q01RrXkbQEZq8uFwsMuzKCzx3YOmwza++x3QQZW6sPY
eh/TZs+UEJbEv6h4PvAenDiH3/OVAXXPwyQf7JcTd0nJHAZh1lj6ZZqg+WBKPfq3
vTI+thdyhL6XyERjqCX4yvzns/2A8f93R3QMSohn4X1IDto6/R0uto2m6rfdtZj3
wL9WZyYDIIYVtNYf+4YBW2UOGS1ZtDqLXzDOIYwEuDtxyTwSfHBrnlmz+1yxn4/y
XfwbjtCdJysSPnWfryGiRZlMPe2tUnpULg9S4ajI4LpfNeBRupOfHHeF4Ss2q8rl
xtNj5B3xqRKC62q1flBsP4Qh/3+hn9s4OM+REg+8z6Fp9+9o0+Raq+Aykg5rD3/M
P3j9dvV7vbj2Uk0wSVW/mcqddjn0FvG9Ah4PNdKn3gnY2+YV1p51XB02kCeuWRsE
QN0mc2BnSUTnSw9X4doTvli/IvfEdMKZlBLyJHlYkIxtIJlxFD8bHyPakn4Lm4Z4
S89gfSHLLAWydqtOlKWjFF3S/85ExArfYA3s7jO4uXrodogZSLSLS8F9rfdC3+9k
jnIkSscp23HHrhiT5MjNTWuMYLZxi1pMbkG6QcsrQ5gD0U7Nroaska6R001QO1ZN
9GCkNsQu4EI7oDXgCJAZa2uE73S1Fw6qpRXV9DK+X6VHfKmp9cXx1kwnK7Jrttc4
irN6vuuCFLQF09vwZ3gtGFFG+LlKAHbY76Tem7ocEwZ7QrOcFo+JlLGeGF8IqGca
VU9EioOpvPsahp7MAsmWvQMnOI/iI45lcYIrLlxtGNyCClBR9aLgEa/kB6jKjKd8
L4MhUDG4fIaq/slbTbAXi2lPf9YNCl5IeuZ6fQpddZ74zAVyRrjAe3oNS+Q5X5nO
ZCAdOGCTKR+m5Is7NHreYYIJIPI+Yby3rT0EtmEEe+Y5qItyhozLSCRnGnoKZSyD
Oo6ORo2FbVnEy3MJhATfX4gbpKU2E7o2r4/bjuTCkAv/sdBiEuN8kGn5nI2Z1tgC
r/yVV/sa1Pts10CG/3uaujRWYX0o2uQcLwlkWwuLsckQ2V6o4T6WfUpD+LcZV5qF
qKcAcTutCNKlg5O/MaHOWdyUJRr/t4D61lUVS1Vmo2hhgq7W0GW2K9LgRRNwhcEJ
XK7YWY3vkbw9QYwWALN24NB0jfep7ijMfgq/y1/9zMcUd3jlG9Fn5exPMmdj+sdP
w7tg3nx824/fVr0t7/CUaanX3NtmQsm5kT9nC9QW8vrvDe+VJfTTODAS/8p3YJ8d
FBUmIPaoXninvM6vYIr0hs0a8Gjj1ocMWcYHtKGMZmO+RD8495Bun8fZco0dhi8d
HiFdQ9cf9NPJs/t2VHpgd2hwQDLdGOMdnzM+9WIrJ9vchrnkkW5AwI42M9GUI46p
awDlqPDspXNfW2KYh32FjEMXlwmtQIKdEkiI4qvrUAImtciaxSIFSdBYscCgIvVq
JhbuJPVMNUqXY02YlKmzfo5o78r+x4pZJWPVx+O9RNcC0wV1cDvfFUZxnVGQ+XrJ
v68lAg8Lkox44sOkS5Ba31sKfZgN3Vp5FDfDf/E1KN2VgsfMFzuzOVGCWNJ5zdaF
ZdcjzcsJHdS/ieKN6sixO2WYDVHZMaMo1MnR6xUelcNFZ2jg3YtPn+J5O9UZwWEn
HushoQUgM7aU4N229y6AEwfTjxjfpwYycmqgBrEB3ij28nlziFw4gLtcd0LnTJVU
ecby3UUwExz476dYspuOwoTNYYCISU5wz5gR+4BUBY5TcocFdP0JjjhZ4Y9amna0
5q76TlpCMFNf8u0xnOwhU5jFlqOx10ZoOrk8/MCfSTLec/DHRHKMUqnal5h8cMn1
swCOAWT01q/1MkhvDe//ps7OxunMJeW17ZbVYSGa6OLUXB+kxoMcKi/TqzHQLjdT
EMRjeYvKiT0RoWFZs3qVOyk7vybW1aya7YhLTeg3kPeYuYbV6UqyQC0IGeq6zwjw
NONTDb7ULcA1c52pgrv6dJ58qxa6zvkuy6HWt0IwZ4fLrdI9fSgfWh5f3hlMAZDO
FeQSBEOtzsCJ8Wv5/+0Kl+sHgAmuVM2CIEQbVoeHa7e+Ahje4L7mpUabqWU33xr4
SJw7xZEsn7SZcBARTBJiLb3Iohkah45hLl6ps4XhFY1tD/SKCK3PETjkkXN17ZbN
oir2s7CZ9ovTImoRRDMPSD6rGvOw5ZXNKdAvSXoBpAergJssxlmiFFHK1gDBATZA
gV4s0dlnceuhtiA8DfjjXL6H5SEllGxagAdUx1EAlsRXRu31XPdADj516U6Aqfwr
T6AMiShWdLPrZ9ahrC/70m7ZAu63tvg1RyPmE6flqU1zWmG5Z5oYKyCW6ETop0wG
BsupeXmIm9omqFAah8jgLrSgpwwE6aytokxzfUKs4kTLMlBxY/DdlBM+VasYG291
k4vkH3B8k/jO3s3xCHui+buMLwxpMZV/ikuIcEf6TqJre0Sgv5o4ICslvsVFiRAc
sjW4ud1FcYrV+VvxyGRzR2wbhIkcnZi7FAmBmP/3v5rqKVOBeKb3dvKZJtJ/nwKn
q/GqeHoqaQ6iLD3K4rOTteiRfmsxqcAl4Nq4yY3yADT1unwNonElueZ3LAfhkUkj
5DWELkAqnieBonRBMTe0jn/vkWhyIOLSdEdrgUrDgBeJj915FhgXlXP3w9NuoDPd
U+1kZqIGXFWn3fd2zcAboOjUEAiIrauVEwErS8kwdRPQJCIGpNlcuKpP2u8R7MLY
446GmInl7NyqFIXxEjpNb8V2nkzHsFP49+AnM/ukIrgMRCfkK88h/tGd0ER8+RD+
yeDp6mVf8nhqHqJm69ETu22cGMl7Wi9IcuFO9OQz9y4lJIHgwsnYZA296/dl/XtX
CqMzWHPuAMV+zXrJNok3c3sGMazpTz9aWlpuqkW46EX3gv5v4m7aZwESpNhhR8EL
7A8yjjlUwZ+QZySOeScxJjMhRNHxdR6dPhH5gm8O0/sk+HJk3O/owPH7/9HE+BMs
Usny8qqstunsei92Z2+NXx01GNXe3Urj+7n9sKgU6D4JVGsqvmVF3TpAwxNQ4AiF
ycRk2zgcQBY6/JtdBGxzgE3ddrcogJ37Vfnb6NcsgLFLWlk3kFWIhMxy+mwhPXDb
qfcPcBeo4wtJBbWCOI0WSDOycq7utxtS0n3/nrWEAm1S7Oty2LSOsneNmLB3wUv8
Lp6Zt2zxsMGRCgips+aXdKU+1T0KKc43M5ruTMEJ2dxnpW6fUiuCEi1xp557kZP8
DUniCakTmnsrNDw+wRruDEZeMTWi3oFkaeWLCooog8Ky/pNl5oKFRZzwrPC5rd+d
LKUDAp4Izb2W1FKhsmULto9GVvQ1EjkCElEOwpsjJitOGsavVgKXn1SD7L7i7gd0
VgR/hXUHh/FZq/SDXjOx9Cv29xY88lJNNrRwsvlLjqkPOvwdVm4NbbwwhD9tgiUS
VdC2oDjNw4rN/6fBZJUVEgL3W6J07IU/fbLEibUr0Ley4Qsr0V8pqK7gylVb9Trs
RLNzGvvKrh6OtjyQi+rAp0RwvgZUpVtRgdB+dkTQKFFxdIziMoY/tz0KFgW6mJwk
OXLsIUB89R8D0du68D3DhMXc32oyha38SGeRvGAiJoiI2ayvgk6AS4z0nXPnealZ
puCwOnXzVv9CRqzfQWoGrJ+a7USQZiBuCpuJUtrRFt3rphUenDr7Sand4C8EOrUl
e0uDUtF4UMCPrmNskdaVt66AgHf9zP7DBOiqZIsqoENbYRM2lTu788e98dQyT43b
+YQ9KVPcElw37RDGHK+BK92OlUG4LVMYhRFvqWP72jSwPntm4ysA0PTP7ZSTThWn
qBYcxUBqE0LuFgLhoEukkZ3fVVls/kfVLvkKS46D9j1oEqdjo0PPg+b6QYVgPzfH
6SoV9v74aRHa3RQo5HDuqdJADjkJk9tm8jTxsdYhmr+RchkB6ZJFHdN3egpfQoij
bfICy3fAGsVA4S0m7aE4Kl/m4QbKsnEa44zzn3OfWHhPqgv/lRV1PK0VWZVD3wSy
k45lsWAx4gby0JuCZ4K6+n2xlTJmHwHYpT9v7dfcoNQmm/6Jiz3pwPZqQ5RE38hk
TMCl1cDlikTIiq2Gf5ehiAfYBXOTLO3933hMr3BRpKKv5hiWPlB4izxnGeTcIm0g
EcfbpK7Uk2qy9/5ZPlEuYXiA77c6D2Lc+y+J+p6amQwWK9ASA53adsYNK3q05v8K
QsR08OLkFsK4zWkz2RrBgxzcUwhok+BZAYDra8+LDsi6iEtPQvuxkslUuG4A7oKB
T4O8teRq5dFkaOWaQm5Y4fyfX7W+bQtQJiO2R9iw+GQ6s4grQTbNSDlRYPp7ElzI
Nrt/FoP9CGlaxLq8KmUKup1CCLAeiZySUPs3at0/ZjF3+iOO87Tjf4RP8obFUs2f
mr3UIcr1JkiDSg2OayMzQ41w/ZZ6FLaLgedHWBEjvQKYQIsZXlfTXzORyxo6zae6
BVpUK+mFMXBQf/t1B+UeyQ71Pmgp5xweQKiKjWZH2BvzVJZu+Vp8CT8+m3hu2pdy
MYW6sw+ptOPt2hnZRZ2KeVRz004OBPzf9dGi7RQdxfXwLKOv59QxIskUUdzwFgoj
IJU9nnCIYywLG0/uWaw+DisU61pCX8KVgRFmkXzCMuOh18lL98ASHKIq5W3o45mX
bxisr44wgZRh0jH0swOts3TRp5539PapKWJ8Qz3g/DWG0fVns6FTyyrnlcqKrifA
7ak6h1B4BU0kI21QnvQkcPgmEq33ypeFNkUmXK2ZzZPM51+Tkl3q8V7U9F3b9c1u
/O7bEQas12K29duXxT1tmvb+PZzFsGJcT8vlKWHtF8bvyJrYMD93rqS6EDHD1fzK
V1tYpwegfjlNrOIDSbN565tzXctjT6hTtn7+0EP5atxm9W5T1BwjyXzuC0wh7Bkd
U61+81GAP4tTZ9y3v8UrIFTgC1hhbi56bwZcG+9p5VPDTZOznlw3U434yWPa03Rw
1e6Th0LCJJZTiPkQeLOrC21129jWBmUc8zEfWs0qkWhlUbQFzXx84tY2dQjjXYCP
1kXX7qmbgFubImklbRt+a/+lmXlbePRdUTo4effSsXpcfloj1ocsZ6x/HMKXsh8E
x/ryG62ToIHmiXBDeoZcVYTeW7BBN2h/mmccJlV4LEBmkb3/7de9Rqo3+Xx7TFHH
7mI8B7Dmsf2I39azn8kWbQqllLdJauDFrphAlr3qrMnIBgJ9BawljbGn3DsfC2/u
MtmFhDQ4NtwSa5LPohCNLnhWxoBQEqqNBRzPaV9OnitDJW6hSTeYxZrqr87vSV81
qK2hj+yuHQJ+lXPLqpl4BkHUrYKGbDBSl6HXCvF/oKyfZe27lwvYCBfKylIF3x83
Q4MfIsoQdyCPQEPvGVF+aKDRpmIjeaIH4jrbcJBkfqU6HHIXohd3scFZ3Nmt7v8E
MKxyacFPBm6Zw3dSp6ADi7iZmEUkYxwaKH3DQakG92BJT8CJlIl/QJz52Z8py3H+
CVlXLlUuz2bafs2M64Cc2Fw60J11ia0O/U08WbWbRYQkrh3fasLAWW1ToSgs/s6/
GNBSO2u7xNgeCOLq9E/X7phzCruyWZZzm3LjTvArf5qAzlx/KnRyCcRZn6egGFcc
NH++oeUiONy5ExeZ5We4L+1CwnydrzTHLdMbzC23bSCjviu6OJgcrhHsdbWBkLta
e6ONq832u7zdHLyVEeDU5pFkrI5u/VL/1FDej3GEhZ/RbUaJJi9DK8pzl/6CJ8El
V/OyhmG3EyqRph8IqeDlIw/hAcm+hbSzxzjKDmjF9RiDoCer/s24FIHwiWhbLQg8
alenHOEN/dlEOTmy/Soen31KgS8Sq92GzZ6bJ6OXj0Xech9ogzQSCL5R9BDJi8by
6sjgenfH9K4R+54OsUlFvzHrVqxu308D9zphpcKf1fafiFh2ckxFfpXa/3/2KoNq
ISCwqChVrF2uj4BCmHzli3BPFkIhTNuN86uaVDsSMpC6UjaA397bLcEWEE9Tt5Xu
JK4HYbsKSv4wnTNy8syubqFpJhXbUUA/WYp6oPAZCv/aw5xC1DI/t1h1JviKUy3j
WuNaPuJJZMQy+o1mZl6sULPyopPQkn0oSuYxymR+Y4AFMyPxHQH7zEwtZRAapE9f
W13vck8yWAw9HbPf65DRPArTtxxcEPyGwIDNEE1nhvDcnJJSu1qOYqhl3J64hUQO
tG9HsJoCa+Pdspoqt9hkyaKLa+HjdVWRikDZM2Fpm9sfFPrHmbPRuq2pCdKF8W8o
V2mXFw44/tW5wny//kAK1F+A/wCfao50JD2vVvpC17TrhB9yEJSBdbj50YejFCC1
clmaIVKsnybtq6U0Zxjfo8zonj/ePdjD1suMvMxq2BAvoiOjIc7uLOfanqVBvcic
lBAg3dAUZP1pCie1w96OilJMtoKpaJrjdAut4sWtAKi1gPTZ38TIs6CEHKGH2B+j
jB3ZuIarhpwgiQppVu6Cxe3dwPYOdSBgwGkz3leVJS8y5pQsVGsU7BJJrL6apdTy
kk4hNLj2PYTDmzPlfJHrKNcp7Fk0fI4vrSIKQjIETkeFiunKuSOtuk4jecpjJ70X
+wXAac6wapUbL+lXZ5IZ4Fa06uUM6O6b4Fa6uKIzQimZw/TZt/5EpGhG40LTZtzM
yVAZmaghNg8AnDPAl/Vm3brDUjRz+tGm+Z4/JgHpIUhBPaeVRepwkSz/KSBZqFkP
GBKFe8TbkSvNmCrf/Rbx+bdnDl1EXftDaYTi8deHwwmukPZ82hXkYGgLQdciswse
ZnshhAUOMX1DIAwFd401bXpc0BFir3G5KHEW6jfNvGxFn3lNFaAgi4KmFg2QxQDC
CbZylJTVUvIylOAVhydGAkkMH8wUmjhB7O1PGY+cGfiUy1I5rF8LvVgMYEZ9QRRn
xuem7DNZAZneoSi1X+O7uwyjXfHAwDrYXne/wmSHsPMdO+QowXPiHscmB9GK+65w
3F+SU9PA9mmaEhfkggvW79wKYJl604raTw5YCx3jxmJzYgoN6wC2UHsixPwfe+cG
kNTM8LVvt1C8vzSXhoiYwdvJ6p1FMKGnvZ6djlbrto+cWxyjRQdjrlzFjtxIFnM6
FJtYS10Xq7cuUif/CHPefQh6ceD/sSaPXSTWIOWAzsqxkVVV8AkJCoC0AOZ9f/Bi
OaXPZBIN9V+xVY7SzKfemN0k/I5y/8m8mzr6/QnE5+3GUvvFvyYh6LkX/Bd7AcE0
o6rDBlDJPy+WsN0Pe6g0k7mdoQSmkIx/17dzy/3cG9t7lB9o8cfVobcLHiEwJdgj
fx48bOax5fpugkD6s9X1xd9NnSWiKleYaQH1kbH1+kcz4wlX8cBZ3Tb5f7jc3mD1
hj0XA0Ye+gU9jQyubD2zUxDutR7YeldPhKNhPhs60qwGF7Z1jb6bvuIQ/Wgh995b
g2RJpgntFb2qz7n8xPGNCWCOpfdv19jFziMISQAeouYO5NImXH4tAi+BeELSQO10
nlSTagkA4Sy8mfc8W6TMgVnyE2nJ4IvRc5rDoSJok0LrPi81BUdLRcDPOBccNW74
uFLU7NYwXeBMqkli+zmAbp9eAXMvxBURCvv0FVHfP3xKZigJsCRY0lZOapyAX6Mu
yKbn08T74/oQcdh/Ak2bKkyaqohgc8tcm9jGY2cPgjVym1GKNcRUONoSu7Jz2+2e
fydv2hvF277Ws6t8PjqyPyqPDc0hFQO6fov54qvjlTI+jfybPYB/jj1qwDm26oYr
RRao5mQvPUagXF2J/zRBql45z+wddDTExmxwNm87ujIbuXJtZxGyb8Y0oJayJmXY
UWTFr6oqm7HumUaqiTzum/0I/tsLRyBvxmaGEQW1ecMRufXmkJJSNCGMtkIscZqx
sT5Do/OGKHBvEb1lm9+ZYbc3baheV+TWCInh4M9SUsfYLqDu1avZaiySyCglITZW
bmnIXjlGKXN0rgknwzU6M2vg7o+IoPrCx6LD2CuyWkN8nNGhuAyiNv0d0Ri9n7Qu
TBE39vNUzv/E+bfZ7WYmbhKRlF6X0QFAjWFnadsU084Pz6bDRapY3dxc/WWZybZB
M+MfjJf3McQNJLCXE9eR8X9+qIRmzErS1W1NHu89l23oHmlaeiQovd2l0uxWfvnY
5m2g417xpUfJcvhRW5b08/9l2xMDOG+x7H8y4trZbHBGOVQhjiEU6kGM1yHCacg8
ezOUfI/vlPPan4s7RmPD/MuBtI/3FWlW52w5A/OemvZ5cnjwl+Y7ULoEtGJ82IyD
C1kLu+qSfEzLQa9rn8s5PinFvFmTgpeDo6tDyrn99jLOmGawyzMr3Jdn3AH+miz9
F8AVuQI2WWYPXeg4pHitwQvMpYAO3kuBT7jjEEIyICl7kZsQvR12QK6fw+Yg8oLJ
jN1kUEqtTps9Wn55q1NFpdMExAdi8g897Vb7DSmymP2HLWR4bUUyD3GHFQ9c5cPJ
Z17l/IknVEGYsU2qUfMSX/z44Z+xTu9mAeQn/zoR+50k0a40W7wT5BDM7swIucsc
gNjULfdHgJaba3QKFhwynoz/OD/Ohz5QImeFh8knTZWD8G/9mpNP58L6mCZL0NbX
S4TI2cRDCHSO/0vyPnw+6BwZC5cm7Kb4+Bpj1QtTlG2da44tq8M6/lbJorhnxHP7
bo418paXJXlvgPaAh4jRCExALxBuE+gy7u6eT7JS/WqVO0u+VPt5lwPvGjjdmjZS
vPv/CWI89Z0YyZ7lTbvy5Y2ctOaZ8Rv/k3Nel3prWkzqf1l+/fpPpB+tJS+O2v+J
bWQ7Be2plNHFtYrGzjmGGAEGuqa+gvl/2TT2NJkH2uwsaE8MXQL5sRq61yMvxSme
7mWJjbt4+V+Ew1flo9AMk+ZVVZ6afJVAIiZfqMUliwdut6wSInnhZG5aB3mnyiJ7
7di/R30YIC4ogkC635Aowf2AZJPJZS1STknmOWVkj/NMGOLW0JAgClzeIrrslUin
GYDLkypXw+XO3b6Edftoq1nIgsLlp0PvZwFa8Ly79lSi0rj6IfUY5AtA38L65HOI
L3vv0Zk4F87/0WJraXrWS3jvdIWYrDhVnju8slx+heB0HprhldAzv60lEBSj4Ehi
NYR468REgL8KaoK3xm0fO1wMoDTewDUTGdXtx0+2VR8uvOcPRl1tKzN9jelyB7kl
kCSow9ykBQH1r2iHv3cX0hUIQVEaVetsuq/j1nrsbfI0nRjWArCvWIX5TieW+9s8
V8jVtVPHchHbtj5+Ifl+fhyjwXFkdgUlHJqHiKG4jXDT1+PTmwsGTg92i6EUesvI
3vjIf944BduI8GGpot8gU3MHnGaeKIvUnZc/w8fY2zQigE9hw3ccx2OR6T+MXZ8r
NVbA2NlNru1elL1FKH/kWcX+4Hqzx9Ct0ftN8sksRlKLIWdymbkoYGhmdUMAjvut
ipm2Oll15pmlE36wd2TGADDX0Jnw7OhbppC5iogWtGZWIyyCDd4jxP5c4jlVJqiR
bqGqXRiAZHP5xuAO37U4zcAh2nOwGEkOGggpE2KFiauv3FGsEE4fOz8+Qv+tpwEd
6Os4XyAHuP9j2q22yzRYv5cZo0QJPOAO8YUMAkf72lcBdRsz/RSvEhyrTlVNakaE
c16GwIMmjffX+c+UgkPUtiu8dqXaOlGbThEOIBNCeFARnWpjqyiWOjfTWT++rbCM
owSalu2Gm0AMOiPVXJg0T0zloKlL7Jy4B/1kTPtX4IUDw3Vt+kLVVEmiC/u7zJlH
v0jqQeqwCNt9V8bQ83gNr/LTJkgz2AhkWVZUEdcyHl0vrlY18yTcae/hStf2gaWd
OmHIBNPey14/w0x5AJ5osm8f/R7q+wKu45K5KaYMBFfJPuBzblMrWAEcjEoL59eF
gBPMDJrRoaQzYP6BGf+awtEbRf16XzMGuTTZ9zp1blAMOFk2TN1guxYJNqnIMdKQ
n6npsAEZyeTuDcKoLwzI0ohVioXGy9V3ob2cNCC3vT533xsjF36NQT67Qa9h+i2I
nnc2kl87O2CTg7leBUpOQndOP6P+H+XSa9jgRlVE4Y/jPvwxhNZ8KkP7SMdiSQHS
hf7zMWpA+ji4TwhuTb0kgam05Q8Ull6u21E3uv0bvQB1Q7g9BNkEOhLmx90gm51e
ZXk9WfN5VR0IUMSsqSo3k8gO0gI48kT6gtr6xv7PHgsdDCyk8KdzX2j6vtwOkYdN
KchqLYM6WBWHeY2e0KIC2s6jrs7VNX52tyiO9GYovuGuwpgHPfshO/AM92Omn6br
7e02JPpFK4+6LPcZC3WxLdpyAeHUB+2pMm9siPaXrJHc0SlBh/ua8AzUp0B+fbtj
mypXnW81NXFcq2dghi5ujKp7A+JavWPGEtw17LU+PZ296/5K+q6DZXrU01xKCKpR
jbmsx/vGOzGAp6J6YYrf4DlvF62AV65803sbOvw8x2F3BopTM8Ig+F+2BLqkyq19
A1uwxoR6KTedJ0xpq6GdngEEXUGiD01NZ6UuaTzOA4LB0hVd6FWqyTFhQDN1dNTE
0vUpm41PiGvNdaFMY7hkJ5s/lWOhUouHRaN0+OTEC2UbuGoUSE0ygn6S/T8HOPer
brFgSztYdxnSgpaTjUlXfiCM1mZrfWYTO4tyZXTMp80Xny6Ixc2Ml08aOBaJoVi2
xVzKGNNWXSkTdxfhi5DIWdF5NIJENyDSXSxnNylEiyzq5fV2H7lbFh6boPCZb6x6
mnVEeZB7vF2BKQj3TI3pmKnJxarD/yO5R4hiiF2nEstfxIUSuubKZE/31MXPUDh3
Wq1lBbJvr2vkZt1A+ALINNneQdte7W/LEx99IPOm4wjiJXWDUpYiwvNpc0X5i4n8
NOqiJSLmO/jXbA6jhWuBqsmh5hNTI0eyxJoRyk3VEXVCu3CZV/wL0Ea6sQOeAZ5E
CC9O91PQCbMg3nMVptDrWxKkp7A/V9wNqU/dcaBJSV9B752AYlIeFbPmTiXt+RKA
z0ta4rY4q62C2K69sPh+4sPuGkCfRIjnugCmzJwwALtLf/TqLS5JEC0XxD/sT1t6
3QkDufI/IPkYGU1qwryu2Ns0JNnPw0i9qK91fspY7L/xbgMN6g7XW5oHKyVCha3M
rlYrbutYvpT2m6ZsAhdOSpreiBN0b/I3tJWhESYMDBIVV8JIxRt3UEilzOceiJve
ucHdm8DjIYdUsOVjFJ48GP+8VSEpGgcVfTsbm2ebxnRs9WhdRmhX0cw0wMkF1v2I
rdKVYu6okJJ1qbNztllb8oDLjFK/15L3thwT01HhzGOIM7cKBlvGq5CsStF0+tJz
icq2ZkNkaXb0PTNe3MkF/G7OW/Rnu+OsTT7hIT6OVsGJo3DRHPp1qqae4BIFwBe7
m/yPDjybiee8bIlGTaguLPxcxKREqzaQFDBv4Zj4BtGd/uRKBq8m+eGfMPcUjojg
vfr2B8Oek5Zpu/N+v518YedL0G5m20LlEGIxafA5AuRd43qIDnwodArKKTPpMXPN
36hC0EdZXDxgyFGSNZcANzanlB1XsZyL9aUBN4ZSEHz1mLfNFnQzXDboRwTIVto8
o0hJmjQQj5URtfJcqtEtRE6VpI8sUh9IYZUXI23llXVR9Pdua5tGeT9JpWcivHLo
rVOufK0YmzdkXBDf/0DTttFjiSEANH/mhjpYo1GDNcTHE3k/CbCOS458ApBaJlYs
V1KWQMCz2OGRQd/hII3GBPSHX0+W1nUXBFT2WZ1WctyNqTQ541cyfHkTcZVBAsvd
un8IdXPv2B1lXrji9s55C9Nx5IXbndxYWykZgvtZFYa5GhOQH44R9Sd/z5LTLkJ6
Qpag2V0qpNzZvJyleksc5URlLokEaJskKZMICTtFoXu85AJFExiAUkndI+NMk8le
D/Lnu4aJKG6nt8tq1+7ZJoyTK39bU+2Bv6NPWZ0w0UY3QBgMJgFkpsGDasznmh48
va/T8HnRK8Ok00LY0p3ww6Y+5rZnO4OOovX4sDDkWnWiYgaX/+IE89JV84Lt5/0S
mbTYVTHZZMOpNApNsGEdHt2oEt4zRn9UHzBFGFTh0sh5gOCNmBQNPj2Z9VNXs5ue
S6k7t2rjaUABB0sMAznHArieJ24en3tuqT9BTZHCfVvhLRkdpjZVVRdupjxa1/4O
2ChHCDOcfhkeTq8rRKnqn3z3gtcgrwLOSGSl2gHQFjqaT/oKriPdzyEjXDRZI192
uCKbCjNPwTA7FH3GIxpFjcVyzZXV44EnrnBjRGlq/HFpWIzXR2oluRQEW9DBJhiD
2sZzSy8rbTUNrqIuKjts3PnnmwjsmLyZShwNdCymynOF+ZE4U7Kfe24cbthnLme+
vebAuuAMFBcGqP9QF7w8CC6qvovqSjsH3wzuIkgV8MyI379C0Emb779dNyZqtAv1
N0FtmtDHlhmuAiNbfWMC3YHG2EbMAGfG/BoK2Nv4gXLi5RianNrsj5+4iId3KoEJ
cbzPTa2HynON47oqn+EorxHoAX08sJhV2eX2BeA7PtjkGC3kILQvFxuifrrAU+eS
tqnwmxyeC8sKT5q82e+Q/2qgs3ipMzsRRyqhruNSfarhdve29TdKywl+rDGkVlOJ
d1BDNHM1g2VzOhit8XhykpzpCy0viHEr7KXxGhdaTwJekXMxyOwNkWYr3q7ZwB2R
86Et3C31rFkF2IkTbxHFu+3BgDmBDYXr6zX8IA7Dzn1wMo4XSrNeUu7T2O4Er6r3
dYW6TMtG6fmDsjH4AURg+A9hxlUTyGh341dyGp5J6tZ//SrV3ugWBuPX1b7SnsUw
dTJz2YWbUJHwG74ifR2/3atwgmr2lPH3eeE0wtUWhgaiNvgM9dMIvJHqIihdyuCf
RHFKgJO6TFKNdawLTOnrgp7jWp3kLEeDXne+Suqrr8a18H/fkxcvDe/tc5oFSvRy
xH9TMmv3tLNn2xCwXf0VtuTGs0uqqgCrPtawEv/zqJhlF7jmT3nHnvc40d0I4aab
O/fADOTTc3aljjX5/IpIRR9KGFldW6gRF1SV8+ERnnhN+YnD6VVs/+rtk9GrhK5J
qzMFtKfrcgpimxlxruSeTE7PKjbTVFwQO27ECtIo94Up3K6n94GUF44yuPDhBdD6
QvQAWAd29J6k1IpMBJ4sR8+ryFKxXB1gxtEFd4Y3/D9VWbocaQMUMhA3CmlNYxHt
EZiksVH1I3I0VkTLjoB+7OMnRDmu+kxv4qRrGQ7fFLKdim+cXoP0WAB3SlwnGrsZ
emwS+4UpkB8NDsB7amoTJkAwaGdV6jORxkBgsUdHxttpGIsWLHlDU2+zK7uxU116
2LAJl4EX3nm65RUDDgGrHBINpaIon7k5gWVpnHwnsTjrI5IlK1lmBb2O5AF6CUpq
RfImJQUTK43yPnEtzCcsI4m4cP2Kyq2+Fyh1sUacneq1BnwfEw2VM4x9Wemv2ycl
NGZlL0PnjspeAZkdzTMdguXbf0/TNoChufqisxL8XxnW5ClyymcH1kaFwEuOM9SF
xTUsp93dwBwzaaQlMlUmlthpLTMVL1V5dhwOkTC8XN0InaW/O7vcDtIm9AI6/7dO
nKKGkCu9pN3xuHJD3GOTS8YEBxN8MNElqF7klrzmDPyGM9i2JCysfxjkWaokWsYc

//pragma protect end_data_block
//pragma protect digest_block
AmqIONOxWuljE2J0+hC64KOVM4g=
//pragma protect end_digest_block
//pragma protect end_protected
