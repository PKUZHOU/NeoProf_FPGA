// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
mB2zoKgEwJEgYsCHUkAcCjqEOLJpJRrqEYnjE6QSGVf6PWvsxDd1GjtAPzCn4h8AseEW9+VPkCcC
+vSWQnDSYlt+u4df/Y2KegJChpnlTdDGQ+IQ0j2Vlo7yXqG9L2eeX9V3m+W+P2pzsm1PxS32hfvJ
isiIxguEOSPumM6si5x/AP2OUabvPH3v6jyJtyjppg0+Gtdi0kgnnp5zv2pBsVUECuJS+/tljDyx
5U2yY6dMgWIB9ZLyoFPdHR5m15rVkgOlq7xDti5OLhvfd3YPnRRpf9dZ8le3hgKWsG7CZTGejCcE
jOjfgCSM8MpFoDBNLhMgg7694UDtIAB8yfadCA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 76880)
07zsyvgIUViUyuG13XMLpnTyJZ9ptoPwLZLqvwl2Jocmi49nRQbfoX3/r8WVAY8za27SbKSNJMxk
84x+/WJqGSnjyVDo25ujz1XsYlGMoSVQ0ikLW6DtZ8QJ/62JfygUXO5ZAyPdR+LPWIV0AMNm/oPB
7EkLpWgqbA3KTNkTdu9e8fHnM2OeTyEp0s32EYerdxSVNPh85XchzX0xoiHPkKeihRwYdYFPEj/m
I68eUY4SaRIm98sPIBc6E1ZWr85RRf0j3oD6d0AGPoKnsDeWxY6pNPrglJEIckqpf2q5bNGFjSNu
QsfcjtIjmB4tHHaR338Fkwi2eLnJiN/30geDJ2p/uBjkD9q8vQ8QoLnKshI0xJE1rGAUlF22hfus
y0laaUw7MTTG33ht9WoCctBVHQDsHKrhIq8oWhGlwdLcy6gWMxYhF6zxibUI14LgW/WL5DJUviOm
Y/EQ1DG5CcmvEQrOwK9EN554dO8zrF/CGmuxSVhhhNr1DNtg3tuwxtuMwuBx3WkqErNFRnEDwoqN
vQTWXXKnhSZUVc3D00l1NnSjXG9Kj5MIXQ5mA3A6W4FVLBejAzwhR9cyCC7LZP1TljFcJ9q+gSO2
fS9BprlgErQLJsIVTjg01AzO5s7QA7t3bh5DllV8QD7fyacUTkH3c+2p3V0fmn6wMWb4owoiwm85
wU3LSDYUYWWmaSwO2ZNZ5A18NFBHz7hf35IIYIbbOG1zFPz1q1Xixsgoxu6xTKa3QIGxPjRuAaiV
XlpkNr7Bz0qtJlGYyBW3k7W83ToMAJmrgDUYwBYLKGqOWDvJvBj65CvvqIBTW/lh9D9Xe94H0k34
7P2ggpvwwX5Z/monqNVQXRy0qegXANsSmQVuNLJAAo4SyyKVr9FxwNyvrcCVnDgDLjN4yn2xfvSe
BstTjXPywpEyHWnoMQGfQ6ZOEEvf6A7Kh90HFkcztepfa0DVk7Bpih6vvdeeriBHWSWPF2EZahST
UVFJrfL13InuCssUK6sSWdhzK0hvD2U0PoyyHbd9BdpHN4IDGsarMbWqbMp0v1xJx+p9RMaNjNYS
01FBGUjhhT+miMpYK1p9CSwMuRCPo1ZrRys2D6yokVHo+5h42+K9Xz5fLPLLckaN5f+sRASS779d
02PPKlEnqvvU9Tzbcjem1O4Uubl1qGe1SvJs/GxvMXNavuSag6pwH3UhGOpbMhuKADA+jaxrpMvc
2nFpxxbg2s/tdwrzFpXYmN5dHAuWQ9D17m9C6RZUdhuIC0U11ILj3W+9T+T98fX11KbBg/cZYXMm
6UWp1H+YRaxu2SSx238By4pAJs0XCtItszNGUzkHLfbos0Nu31EHwMk8YJQ0DfkF8GOzT8gNfBtk
A/QTOeNFs9HQzoRk1cEfQB26w9AzSBqPaFh4WQW81Y9ea7YQOc2BWwrMa9Ia6Q0uO7KmTs3EUmUE
wmPEYSfMHnzpx9Hu9wv9UcgIGsfdEf8DPmZgeoE6P9ayVhO6grM+WSL+8kOQnA0pQKFGiQCst3Wx
ZPrbWvaGmSbc9V6CTOzN6YQbI/OfQs3WXinHQOUWpRrgr+r7p8ZYIeHJeCJeZLgOPX1cFnbwHb5s
PJ7JsXyddJ+OtHqe7rPM0YXMx+NFh90GJj7LJAnJHVcFLV8RLaN13ER6AyXdkZrIcdiX91dO3hR8
My8pZE3mS7fwvSmTNqCoJU3mg49I7lvZy8p1XPWdugN6NkKXX4CQMn3ey5lavioxycmtOHGP++Lj
iVa20lmbvOIZAopgmfTZTOG0sPmew2aZpXyxKPRO/RIc1Qo7eTg5MRSGc9TSf27VYpNfy0Ymq9j/
z5wKcqPazlyjkagOLy6p/HVcwnFCjH73BB+0Ly5NNM9/u1GwniMAudpmJPw+G1MLAYPZQBa6eOjG
k32PXv4MPd8gfmA/YbQFfATYecx7h0JGy1XT0ZWkpwpu9cDxx3nG4w9Obr8FoAw8JFbg4jWc24AC
MYUfa0M+1nMU7QqbFHlOXR4NFDGHQinuVewNbDM3BiHpNitSAxlsf5m5QmJ9BJx6FrxJDhEXD3qT
chF4tFgc7n7DQS4rsjSwzUruzVgtvR7WmITo+K+gPWd+a8DVcnOcpPtQsNBZLqqdYi7LC5KaJRRz
3oIZ7Xc4qGkfyXkBotQSCmSUtJwq6bxhan2MfBgiQKI7rA8IEtIiaEw8L8UQMIKwhxOeCWgx+Il/
AhMnS+Armke9x4/CQ1rv259e9tlk2GpDIKwUhFoY0Hq80qsOzqKWJZHTouamVkLKIZsCrcEm1BVz
bt3dBcO6Cwt4ozcG1n9mfSvqQyXJPQ6yDsmOvAQJ0E4gCOICNs3kkpdv5eSphBpObnzZa4i679A/
0OgitOPoXSNtvuGr7ZeiXvYRquRzuYeV9dcIh61QcxJlaAkiEQy4Bm3o//EjwTFeeo9MVmkbhqb3
t8xxAX5MhZVvtqNM7RrtbyZWnY0DwYF+jtEAWafv+TAjZfeuuWRvWVRTM/TuhFOy+deXhSzwx5ng
M1qCUZSxUtbxtnRArfRo0V54RyE4mob/qfnDaB1Hdf86IPwsRUQklr1fUGqqcCFZSZWECFiu2OTV
mcl5TmmEiDwZiVoshfOJyenn1CON3UwotyqIzZ+mPCMXA6e7xAcpI5UIGDRd0rzsoBvlgi2P2mW7
/4M2YIHIikj1uNyUovPALDy7jknbqHyvulFfUCXXg4tf/sxx/U3ULjLz0ucxht6BJmzPbMOcUgei
YmqhMcghDv5IJLSVJoo4AtAauXZ1ZNQRRF2qi7A/gUvd/UV6sM+h+Ls/Hql7SLgxl6+jrwIm7/rG
Dzb6bDvADufJVzmlZgUMUHACnUScX7SzNUT1yTaQo6CBezN3aywRk++x9mh98PBsncEmzDY8ozTt
B17cCXvbC/xGoDP2gdjQxYgUgGjEV1p+Jj6U4XB2d7ZvbzT/Ybdf9kJWXFoLDWg1Wv+PT/BeB5Ex
TyVHs4LYH2hdAHJSmHQ+48HvnzjURNL+Vq0iUUA9q0bXtbMMFm1CEbNc/Fj7YHLUtvF09FGCshAf
fHM44nrCW1MftEVgHak16eIDCf5ZK3lGn33Hs7FB7gg+RTW1ZqU8dOt1Nwfi8q6PE0XhAx8wxEXJ
bBbAccHxIf967w+3+EzEm1uN83FH9MSUW6nR+iZ6sppBUpuT2GGtzGiBRqrGKaI0zy5ERYZ5e3FJ
otVj3gYnyC5uPpGUNqu4V8n0LGIe0WKq5FD88LeEHoi+0SohihwWwAEK2D5+umi0mAmHvWjuEs9n
6hn1h/JYfJijYku0/9KSUeBe8cT3UqNUEHxw7ESl2g+I3TJ9eQh21QCnKS1cd8h5FDnoG4QCmsi+
JSL51IKe7SnggtoXAT7QCDYo7OGR+eTZTfar0LhUwMphleqqPUjkoyXPk/LK7O33rlP5W65rw2Vp
fxz9mq+Iyt6namNwRWe8j4JckLDfD5/fxOGVZvGuNOr0I87Y1SPI7tDy6nRatlgVhsLppWNy/saE
SIoMozOMnsJmtJ7aOiLqYzxAO39nlkPWVTrD5oIdaBqo/l3Z8zY77e1AlwIjSnaAzTWqU0iSQrxI
GaSsJMBLOGiqfqXDsgbwhB8mWeOxTPKj9MAN9uX/npnC3zP6j3zp8U2w1ZkO/mOKwdL7GBYxrrsy
KeFKjSXwQ6hWM7U2Pk1vsBjOqD+RSr0VXx8/JgLKZhxj2cGdYAUXwQq0EQhNJHUR32zLlPN+2JCm
/08Ju+S9x5oEeA4dO9DFldD0eYtKxGjQcFuMR/HO6bJhwqNEzUHxyoddkwQQvtEinwd4T1Koe9Ea
Tx9pV0F0LWXlRTKaGa7TkAjYE/xXmg4kSpYxJxQf+p2sAz/B08n0Uxte5FIVovC0rheNWJ/Fm0ji
qxXmldWpNVC2u47UmtSl5OTL3Uh0qZx9ZuEnLCZ5iD0X0ZP/0mjirMZA3mQHoMPgoT3dVwSqhxll
pR+3HCl8brq0KDcJ52Zk+NOhiJ+DxyrZAEel1xxk7Lkz5Cg/X5WemwApuXVeOdtN9IW5l/aPedB2
7Ucco41rjJ3RWAlyjFRILF3CNXAm6bVjseGLBR+buHuG5SzAYO8qKbvUJNBcRslViqolgMjrZOuO
lKQuXseVCuTpp7r1VNS+3a9hrrJaovTbnFBWuxMedbAHpRjvAIsmO2lQY1/EfjfxjTCE/pDoAd2x
LpUiyVMLEfu4bIfblXea264cngrvgBtQamJq594eS4pbqKZ92f1a0U78FUTFIogwlKWcWDkJyff1
xAtVBO2u0m4k3VhB18Vv6YM0YCbpgVszV19pPqxyqZf9jf+rwF3VyTeaJQd7GQlz42JKX3HhPEpZ
WaHIziYrNH5uRbh1PWQYKMUasuwyYgdHXI9o+vc/xoS0NlX4mCOYsMJ4rO3gr0aQ69TwMqCZXXfs
U56UZzd2zO+agoeOzUzACL2eok+nkNdRvWA2wA/2molDZvHm6vGotTIc062s7hXtsisIxdo4wRag
7bY8+P2qCpUqgo08iAm/AY2Llce5R2Iu9AkpiT82T20Rx0yxFoVrxG2NT55caoBCnffuUHkeuHhC
JhJFkhHsijLW9segxWmRGXIOXap5qmoF6+h/gwD7vBAgLyeJMS9ByuAGla6/nam869LzVB3SghiA
XEMqbxIDcDPOO/ut8dhnOomV0dCIUhXYvTS++45ASKrcAhH5KDBEYRF5YmdCJVnkKXjLJg3t4H3l
DK4l+oet1KtJJIAon+PIi1S+Zq3F95YpUV5plfVw9rmZgmZ3GN5XmZrpI5duj1gYUbizr5lZAftw
wncR+152MWZXSy9kdbqCNj/bmETwpcNTXtrNWyFudNTh7ABZ24VWYL9z95F4J4gYiDHrLR7oIhcc
WFozAMwd8ChHE8sEow+gUzboYru4YZ6cLHaoBGHcfTAEfUOoilkBYNCNrj3IPWlDDd9wKGEB7lwk
zVz1327P1klin+Ano1Ice/NSOiFeuPhA+kJsujHmawioNSB8mkfOWvgforrdwla1p716aDT6zF+K
JqnOp6pCRDILqbegRHLPLDrfj3KVzmn+3+WLKuNTah8Fu5LuUewh1t/BY0h/1IX1ksdG4ae0t67N
GBT6wQjSlNCfiD65K/5P2T+MWU+IACnHDCNK5wKNImwtaAeOmc+AfE7lPwpfc+R4DLBaRDvueHPB
iAarqaDaSOqDoEP/v/bIb5vhT8AqZCX9sH54GSrWoBxqe5d72Kl6X5pl17XnXubq1edv2jPFdwwE
HrQt71hYHxbmOEddGQKFyzoltjRS4Xjvg388hJU5smcmBPTA+MWCZvtTbMyQEqPGuQljPbRX9w3F
K1hiF1V8p6ycPxus+DIZcpeen/lUMyVWduRB9wFWi/9iABSwzqQ+wn/s4z7VBeBfLEf9jp9Fu5Fv
9Bi27RJIvowcKt/d8x79V9LdvJpxkCYjqxs87Zf+3buM24Gh+BHNTyOFGrpCFoRj/Rlbo85ts3DM
CbNyUE+gFZBhhGtZkQ8ku0JcNSM/llIwQLwD6GkKzSIQdC227ZTvxVeqnd+BLZl06EmIeyz744TJ
26OKG/oDopUUK0+LnMeiWVPrThuwuMvRxfpEM4xZqHZPUB5mh2q+Md85t8dYC6GSdhra+xV+lJ6t
XrKWG1JnVek9Ideq6oStt4cqqoKLs87qUJmGjpg/OLhNizZREAORlMCwL0OjjLn5Gk0daQE45eLF
X+jsKAdTlCzboBOHdyKtucI3aYOcSIWlzEKR7EJytWGUTd+pAzx04sUa1A6+dc1kU9ZKYz/8mTPO
BZYM3a4Xut+tC0E/kr5PSMrT7kyH+GMdJK1NtM09+ojYiPJf2zmJTcbzltnvw9h2AS0QJVBvKLUY
DcnDkYaUMccEgyNdtLsIwZbMne67IXGpr38Mo/CQUNgrR6PS4/qxtS74ZylR66rQ6GrjAOya4p34
fOrwBpof4It2I+41UAI1GOnvq0qUVZwt5FJPqYMhJj2mT2b27YqwUe8kDjNAvbzQZWXXToYPxSyt
Fkw9TPAOaVIKgrT/4udr1OYIrkCMd/d2sR/jZyOlh7+UoQC0fUNMU5gwfS1UkLdmbUhzmD80XTmX
wb3zFoJrEin2Fn5Y78SwIAxrAQPwDg8NHTlh5WAc39pimWLEEo0zE9BqToCDLE3cJDzvSA9IfT/D
MNqQIsCmiZFh9JkhyDDLI68nyp8qvuxQbvfRa9/Y7QPkcJ5ToVWerSpYvLLw1mxPf6qyBi5JNccT
NgH4hocTBdOtuW9e6QCoBCGofB7SPtAzjz61UgkPyN+L1oAouV0ttvU4vJnkhKfCcaHULBXsC2RH
LLen+PztJPTWeOJsO7GNOISzcawpD+nvCTRuIKg/kEgcKR46rwQIpjgvc8YHIXE9EMdAFzB6rols
tWQoe1GWU9AXnv3bZS/qyeezYF2f8WOEATGHHuYh/DVSGckOpVpuki2AhjKZwZvw99z5IBGu8iGa
iULPx0tH1fvPoIIiVIB1pkSEr4bChfxF8p4If9D3EPT9To/kW6iVGSq8tC7M/XPV28yhMixKFEIS
uizBkZROALVUdVSnnYJRru/b/soJFrWiZnhQnlvVHiDUu6OFfow06Ojme9sRjrgPhj5cndgWzU9D
Sk25AjrVbeDX3entrhq1YfTBLHI055Xugno5Yz6AaJx56VHtQYwD92SW/gUO0qrNx2K5eKHYF2VH
PtHTtJUT87K9+H4JzXJ7LMAit6Cu4HdoOMku8jbHQwSMFwWHkLAetYRBPnR36yEakjVtfCqRMict
HGBPpbX7cetPB37Sy10/b13on5u+3K+f84r8HTq0Qlu8epA/BApMhqi487SPTFvSjgcOZabMe52f
YbEs/3bVV8i8Z7CFpfUyM/mYs4MwGIgQ+nnc80VI2jCAi/PR8g1KsCMcVS3W7ZeXiYgZSWqhhFuP
enNjF94WG2iEH174Qh5UI3rl7sdyapgsojNr4LQWxkpLmhPKMJl/4F5Kxny38E3erx57Cb2d58Ru
f9oR00AvG7Xg4dVOlo2Za0gxqAA/Lp23BOnMAUyTTV6YQYVdESy97dWOksdMLqxG0KWoT+6oERI5
VgPLBMzvd93SssTMyjSi/vTHyaIUvPiVwnEO80YWkyry/AWTIOCcjHJ+NRzRHBhrfE8lxAjjyIBl
VHTa1eQnwV9FRrG8DvbJd3g4iRRixVr40ANyZm+7dpWuCrKdWAqOigLanPV39A9LZSFt8vMiIxRY
YRqGhKpHKkujudu8QH8yTLkHeWSBdKJ3roSzG6PeKNz1HMHtp3TYiFcrMDMx3LdW4XNRQhxpvQq4
tI+oYORc6z0RscbiGm0+2r5NluHdgCRdJTpia4PoMQRhQZZpBALQ3hgzWHD/mh/s9xZC/ZfJWr2j
Y+pjakfUSmyGvbkP+64ijYP0iSMcwxxWcv7RPoFgSqN7uGyrR8VU26Hu5NDdL/TXMrQgJQk7biM9
xstMiBZL1NLZuAP7zpC0lE1rm4XnepwApFU5nLE53M5JHplfSKlHX+yOEpXnROqUMPF3/lTh1hBP
QHRNA7GQzM3Uki5P87C4//Me14R12WX156AOYenoSz06ErwpEWexB7Z6pmpur4avOa49J3ImPbpl
twCOy+6HtWePCMeyVwB/oDNeDBzjpR/KzPmxlX/PjgRJWtt1MT8i9o1ArLIh+rDCId8fBCMpVJea
lWIroNjtASUXFBuiAJ2nTT3QUDDZP69lVHAfiP7SL/kieSZqCJ0ByhEJw+ImwT2ZYJ/7dco43tkp
zl4/6ZiIAfgdB9I8OXVKkYe4IwUGmcwTOA69xS387Ai36EST4uKheVxQOfTk+O4qSy6ey9an7otj
5hHpqvwrHjHYT2M2lzRhwOPYhvDHhc0862h0+7OgcjSRzmUPKnBcA8WcG383hvPEGfecYWw6WuNE
umgCpfjIHpXpNX3UD4xvyHBzXOmDSieJ0hH9DXAy8Bm3HKg5e4enbd1iZC2mvMBO3qePJUpTTJkB
W0KXNxxt9gPJNN2HZODpXNgMtPM58hLJQk0H+AJTjjY1tPyB0IGL72rVzCpxOFyElfL7yImECpBK
XUDqOPopHnABxNwGF5CFDzaF04GQg5c/YlBl+vkwuqNQ4L+R1SJpS7Y8x3DvOk4zYfw9Tdlx1JCJ
idFw8hKRPDqGCkD4qTu06xBwZwns8nyEmFTnMDVCXTlaaZjv9J156nm/Zx0OICadh6qVFB8hDz0x
nFFvSJ3Hg98X9xTu3CaysHYkJCipgPwb1DoqCCH2CxtnlVtzYXrQoQrSyygqPf4Hbm+UMkihe4zJ
JDv2dZ4dZ9cXPhqB3hO1NwJHOGy6st6EJc3QfROjHKqox9au4q3X1O1uSvhi9ZW5nO22uk7+ibIX
P+qddJ2KQPVsG4QcALBwzr0nUMNR0t+npmqFruul1epHaEEzZrrYIA0whY5gV5/dfpjn/CpThN0H
muCjlGw0fQ4SX0siXi6t1KpmwHLFyez1cQdEGdHzw9dqTBKhRi+1zTc0Cm4WTY4+/aQ55OlQEMuQ
ibD8E1uxGchxgAw81WW+9B986oNmF1o3xuEAZgZFpgulvW5dPcaOoH9M44lHtJfz4vuq7JcFIA8T
tKlGF7W9lXTY/TvDbxCCmzwTnK/l8tMJB/JzlPYggfO6L4RJzdFB/38Z54n1PdrGyXpWh8R5Vc3s
RdJ+CBiEa4UxorG3kTL5EJQEjTyGTqB+5Gvx7UNBnmDehwJyYw3izdkwkHHXRaeBRvlnnzfZ1rHF
H17Z07ICTVzee3u9szMrolsJsnFgKOyHk/toCrjk4wbt6WeHKCSQoVoGbYqClf/hRaoEjDTQ4m99
GovVf7/WUTlVGxs7A5r6XYRDHhQhGJEjZ5v0NnXjDmrmA6gMNF//SmT0LHPAR1uDcPQOcpvMTFSy
EhZwNJgxzG5/apxnF+L+KzOum/cnL6wWX5Y/RIY22kIUlHMRs3/iERADM0uiCa+1EpgEyOrVAdhV
HHt5BIziAEreL4pL7fvmhN34J3or/DQSBkP+CRT6igl1rkEJmjyR/75j9rTLAbfbGzQP/C72ub5/
I+969sQBRAwI/A4NgkVRy0VKtbTyDVsyvXcHp/0F5y2c/lcxyQxwSE4/6GlXszCDYafZVD70Ll3k
GzD3+xPlTq+0O9HcJBBCy6w5CzwtQnqSB2rUansOQOc3sASm6v6EMiWr5pX7axEVwj6MM5dhalXJ
Ew6JzxCZ4/1K3gmU7qrdQjQYKcw4Mxe55sAuUhsDEhF7ZuVlfrgP/kqkwWL/VQAFRNCLx6hGgsNF
DGfWejG8eqDdaG5GDe1DGRK81d2kca/MYECxmD9+VqWfeHUJB145f/mvS0gGgO8V3BVDZOgFiJIS
VwffUvjk+i91ZkuBq6bdixMSSPfrIDnYwGpkPfapv6p1pN4E8ofNVxA86M0jK3EDik13ZW1YxKBf
bk7qsYdhTjlmex6tQYzDtCG2AuYe4O8T2cZ0UqdNogn7aW8HzTj4h+2jWxX0rIHJ/TR71Cr3hPTi
2l3IoZrdko2YF3vyBINpD2EmnC4I44PcZ66BEBCyEbNuo8YGbl0aPAWE4eC3cL5vouiUif9MfWMI
7SbPQRLhfAKCP+n6s4MkZdioeGMuqR1E7Z4KGDNNY+8WbifDyc2QzbJswQkZ71uE5C5fFiuyaZ6n
wvpK1/9IpNALVTfF50eV+ks/uA1QMQSDFo1fvfiephd2gTTRlmFPBUYgoV1idLxlaum8eniJKBaL
KTMYdyhWjAvw6VvFzXvcqROet4FNqge6RxL1l/CmAzkG1vHZKy2izjMiJ1lV0q73aszt4A6oCKGq
JEDCbncJmye2j0XqY26j8krQF8TRJUBeODKPuTSBWyfL/7goRX91yXZBvdk7QEaGzIYX6lrd39Qh
1qaUnijtj04uOpV8TBy6Z2y10WNdlHrlaNDgXApE3RaUCrUh1tellKHTc6BM6mxiY+2OyjlO/odk
nuJkdv8fpzFHFGRXnD9mMAUwwuTRr5agV3ff5tK15GcCpvo9z1tBXb3aqHmhYyFU1pL1ajDKgrXw
ug3kQjz0QVnB4JTJC1XNGugNUZivg2yZbAXhDLUO9u+qi5a7Zv3y6s1k7c9JxJohFUKrWMsr4dQ6
pJi9C7HokAvbb3qE4s/wU8q5gUL5Bcd9ZzAJB+VZL97NSBIRh9lD0AEyzdM0k9P1iXux2lKslqfC
7BYfoNuSRVBFtdb5OI4Ic8+C8ZIZAJlA2B/7WYH+D+RWWPTiZadcj4cbQeHUZEYK4QzqJEOXXoBa
EQkocHTAkmE/CkpLbA0AIrCo8TGmR8zwb4etT6NpxcJk2X3kAa9jvwk52XdILFzMZY57QJLUcZLe
E8PPGXmDxrCfY+z+ZYu3HqgIDNrm4ngrb/6mdpajmIf3xvGOOWcLsxBL78Q83KUAfxr4BkIz4XjQ
FFo8lE0Tt5C2wELYc1FnCoCV1/MyN9G4QnV4kLZuX0St1FkwDMLGYJdxUlDyxFXA++s9R+uK9wRg
y2uzqkagO3953vZ632J0h6ztq27AV3mIArVd9up+D7nusmgR8UzYQR3k7K0JMb28V9podJrfPSMW
n6Ysw344Qn2VcUI7VjRxpdmQBln4AcjVCM8nwCud9yNkzlqTwfjJ9O7N52VB1LrPTmgc6qICSGFF
2XWWcIHYScYFO7bCB1ziqAsjWI8K0OtxhvtdH24MjEK3vJDeI+6hCACalFSZEqm9WCKiy0Hz+Unv
dpBSe9lk5CBzR+bzSQ2PAB5JC5lWBu4abHYCAnlKg1DxIGA8SrfAmSR44DaEJUDhsBge9znbj8Hr
Sl6og1XoDHYSQytjgqsXR5gFjjDZRUqfq5wgFk9kIJMok24GoTfgwFouyeXpNkuGSJq8/NOFpFig
YU6V1/hE+A3r14welAJI/MkKN+apeflO9iajirDl/Zz/PprssVZ+Crg6rtOxWPlJqx18/WU2egJ8
xQgsdLVQJeb/T822ieX3COmQYJ7DNFzFB4IPguSaW9eqtuXyi/1S5HPw8YHgMvA3nWOSahHTxEsu
WiPeXmpomkmcMv/Mb8xwujQqkpfDE3Ql39cEGkFYwjw4qxe6dI38fbMT32VL0wLGbjPJNVfX2k2N
spO4ab9nUzSX3USsSq4aEvJZ+U2wiLZTl4CF/KS5u+Wg+A2SeYvsvsqurKAa5g+EIlJDkfY05B1I
3DjAACTT0ucNTpFADCVsoIS3VDz+TY2UXLWKeyep02gaaBZLra86zW7WADAySrSTtxIcd0eBDs6G
Y9lJokzSfy5+Y3aBrs+2Hzy9CYGSxegwCCfbFuRwvglbSKajveH/UQDw2r8i9f+OvT4e/GeKCxYc
xdD/gkhvYGs7G/0XH0t90a5EGK3okuCeAmQs4YZdqCN7iLuAmnVCf4N4fktbBVxgkaviuAUAgYo+
kVrpA9AZuF5j5+72l76gxN/H4zly0G71qU+ZhcGnmLUiONoCJT++CVXvfiTndl2+LMr9Ml/CyaOf
q6+bC5uJrc6C2tu69PfwWtHNXrQiWMtPHI7XY7ZjIvtQO1/GTnpGBQULcRQI8UKld2wrwyo69kbG
eppmZnoDZ0V+lsJisOnB4IyEhApraQ11RGRGv/HRdkmzsuTUB0VY1/E7XkskNZhCRF1c9xkTpL0b
2ijw4nFqTf2YG4KHIVOLJGY/vPYqfabpeDx5sST/1theFpYObkJlbispy8X2fCHov03abvB9ckP4
t8ymwZtCln4/kGWd5z1Z/DrttCq24i8y35W6D+lS2CjJIXxuySixujH7oYIDKZzw4bHDkxkRMfGZ
c0NObSlcHa3cndaLYkCohx2ahrQxaER/xZtzheO/oH25BaLrBUDMoxPMu15nCTNiu1AhMUJ89DAE
8c/BhcXAiSN1GYKz236DN7dlF+gHusclrnjxwM2IK6eqOe2hHhrvMaSsACzV2s5MRCc+UwGK8rEB
maw8PgT/glr0STdxNh5QpNLeXbPu1r/kAuuGuUT31gNRTqsDeVgSaAZTcbm1xEbhf7ySzuZpxMVH
kF/Bx/roPKxOnYMMp4kisNGeBVNOoEkdLq2RGtkzkht1MbHr14AyAqsqGr1+Dj/pkPSgB4FEU7Ak
F7CvKGf18XbyGQhO9boFCjU8b6lqv7yvdPXXUuELY30TwwzIH2RZ0yIxZ2Wl0fK8T07kng8SVJtf
Nw9QfJQmtp5eEjtlP9w1ocaMJ/FiOh/l60V87kAy9H9laIDVO8o3g3dU5SvD1dk1vQQQ6RD5JB26
MF9F3mPulgF9aI6UT6qY3cX/KzWhM8JuakRB4QG7bPK0iDrCjbwjEPZHMFZ+1wPL2ljODbFnd5TL
bhNldmDYzbaLFrnTgum4QLWb/ppmacoaCrqfC1N0P1VjuvzX8wwChKUVA6r5z2d+txNEkzUgDqfN
dzmn0EAYFlG3dHyJPn758Y0EBqYKAJ5rkR4ySwypZV38z5TvLz1lEDMZuHCG0JAPO2tP3+n9dL0r
qF/E5GcO9MZPVsdyERFqjBv8Pd2gXIahBN4QUms4y9YBULFNT9jp8LGHjrQ6h6UNShviDxPU8JnK
fiUbE1ykS06Zo6GOY9fRgLjBbZjG7rGF1sHnXHmTlmRgedztds9W0wRgsNRVzP6E8WdzBzKd6Jto
zg9B7qGKMhnf4eL7BOVVWhRpeAxTQy+gh5NSEDbw9M42XFatFdaOt/M2oYXP+zntWQfg7LnfUtz7
pLQ1ZF8NZit/wSOA3NyC7HJwM8LucZnu1Kv7O5i2v/Am8jUHImz0o8Cs/B2t1OvJD2f9BX36O5Tv
lhP7YaiN1MI54GTz4yv01Ld3WFsWxT+KfA1xdQSxphXAInAl1O6SVtuR5CVSkwPPfKOoYCzJ6Lae
sdEOMBjtHCPtO4a/d9NNa2SNl9ltq4c/UlNVe+SjM/wSvvaW4kSmkkYcyey37RkdTbiC0MCSBw3y
pqbMAbcNnX+KZYAzcXJfm7IGhGhhJF4ex+fsZ1I1M+z1ZCCr/Szt5Qn6cEXleKxkroTWNzXolxg9
oTe/ixutrHeIDFbc1r3c7ZqcgqkPMfC6rNxv9GaVCVeskIer1dg+ubbKMssFPapt55/DpGr1gsnS
WyZ3oLmAehMz5HfU73UilhwvbPFbjPxFLC2/r7gTM/+6AcvWDTSMK3Z4bNHUK9DzA+jMF6xwvoh0
Ky8oDWTGOSwSBYX+ayCzDMgn7sORD1K7LqJ+o2NDX3N7TPpqUnXflO3mGgB0G3a1QyI1VKSoJ1xk
HLV+lPxpZnGgYTvWPOfnTKUBiElqYNmv39kykjcbOWJ3zVN2spGh/eIqK3vbxOzheEVH12UfpWB6
k5lxlAiti2QSR4E/MOVEpqiD9L6FBTDexNMoLPtSeBWqXVMaD4yBE/c8v3KrDan+GGJC3UA0X7tX
3isH4Fbzl1o44tHvMSpD+aKLL+osJoDtJNVfFxYaBdU1zbTrdRl3fRFJNoIPQ7Eoy+tJB7U3w35Z
4hkiSNchjljOf9Sew9veEAFaXyHjpfGokn5qSr4sb0RuhiqgjYYzxYIhLOgR4dHKkRPnqFgnXtVH
Kbku95WqFYWJayy8RTHftnSaaYWFyj9adfsHoX9My6yW+65i04HOUQeckHAc68CJPVpuiiUsXjJr
RqUMNunEsfSk7wbmHWeFel7iUyC8uaKFFZmmLBD7XydlE0oWunVUifX6vpVXcJRDvHpb/UtGn2Ob
dKITAprRulx/ToREnfKpDI7AInQ1XRPE1gyygqR3LTSynlT4NyTChTkGf+KEbzF6HpqGm6zP92BV
4lPQr7AZmGCgR+kJlSo3OEvA36DWwS3jrc96wYtvF6p/YR8zYOEUAapRu+8OD6JiXcCfTGxIDmLb
rs6dQTBNAZwC7yu40GVZsjY/+DCILxtD1Bu7NFcQ5b0nXfjJdVvxY1K/80uhwXzaZDzRnJVGP1UT
LwhA1gibXwfGrfB2vCfi89UGktU/C23jgLq2oAv5I0dw6gAZ/1xQD/hk/V39hHlROs5fIcSVkZ2o
KvZUxDaeZ1UKpNgI28D+pJck7W8+odm3GtOBKseQO9mHgpuUMlcwO+KJpgSs4FvMRguvayBtvWu6
itfkYM9Mp90KaKYQA12mlIdELETa4e1cVxKMXmtCCodSlrsjR9I+/GIj3UBasvw6MeIYTMKGBW+J
I1f3aPJTCrSL8BNnWro/kDkHn6uAV4YhfITT02/VmIT7rH6zHTOkQuPFR/lHmq59W1wsF974exGK
sCm7in0mdfuggktr149D5Zaq/m/3/Rm6vbdDtxAR9r0J6Iw8B8SonBuJLPl7A9wG6uodZSilWoWs
0KWHeorqvroKuSYR0L/QAJrBFnmkmRCntifi/Q2xTR+9oneasgHJrUPWTUCVhzLvjpA/EFUc0Bix
/uTUqc/9LY0r2Wn9HDXVkllYhyFUoaSMzm8oLGI0pF0PvKC2hasTlafgxR0p8I7Y0mk7KLDMvWJY
PxgjWrh5SGFeUa0mCSTufxVL93aaSqyCduwuQhEgaeKHCP6rVRc0Xfb9kbclpe6lQHXLEI7vDkV+
Se7dBRsaAkVqL9PSzvevhUPNjdYnZtO7BG+n5draIc3GewdtB1l53pOVsZxirW0GuEcG+6ej8/Mn
7KjDXxOPmcVziE+Th8efUTyAx9oCe6iDJVyNl2Uo8g5vFyNuh0YYNwqCKjA8zQxOC1+7OWqCvTvk
mxcZuRywlc0Zl4dTblYK7HlRgvi6rdaAe9M7W2YdCSNH+MB3lWeNKHnldDlFcxUhnMCDDw2J+OcR
VPMFr1F+G11GiPmxglqY+PeJWi2e//0loFFBKJjPYrm88G+paj8rnFQFkNEtIZUAfAsH9IFXsINY
uDq+a7rOiKxbLNaVScVBc1UbhGWj8u9bdXT9vNa6WD/fKl9ddTr0RMXE8jGkNLBWbsJix/AzQrzr
e3iADGqAZe3nFSojpQow1aoa6+G26Yaj23hI66ZPP738BjF2FaJtsICQ2VukYVouGADSlPMgfPDs
pvUZPV7dwtUvjAeOpNDh5JP0ZmObyu0HGBDtkpANCsn1nxpEIjgHVRJSWLk5y0Y2xEAEKT+APsqo
vFm1mI+dbHpOybDVJvMxe5lXY0h5ne8gqEKx8srL0rIBvF/sgCyIL3a4UCTY6GsJK+tsAIpao5qZ
QUQmq7+laiOwcGgTF6Oo14fUDkepdiGz/rbyeRJssKvVTxkgBe5J+bpsKVxlA7NIlrPj7Pcjz6DM
IA8k+5ml10ZmF/n8DF9JMPD9xPdad8xrDw7ifU+gGUhqvMQU+hlZMuVvJIDXxgoT6pY6AFmmEpu6
Og3f6shSTNdGKuJk8A1Frca1pUzGRUegX/mW0eiIuHvNDD07afUthd5UO3h8oz3WuK9+MhRonExf
LNjMghygoKFJl9d8x1ZV4aG71fYy0ykhnD3/gH5BraQVRrzpBhdG0QoNcRlMiRJ7CKvYN/2GnR0s
8pqUkQXpj+mpiV1ETpxVuKZ544pNDFYQ5E4DO/gOAaou9LHZC/SxoObxFulJuuj/jVpxFLCCMg4v
rlznp2bz0hT2C1x1eYlfDyEgZqP/YBIs8JNnDx2dMVKAuMyI76LeFlWOu9zpQueOulrs6kM5K2LL
QrHXdSIzYIbF7VSY1FN0UI3hU05Co27uzZgU2MONeddrU5/kPv1Y2N6gl/PTFtpqSrAhr96lh1aV
2G9UAtZWB8XmZFKxWCuJptDw+kFap/Dc8zgrlZgVOURV8dWWfOtp/MS7tRS4RV+iAasme7B6eHwe
cjBuH5PLeCvg6b7iq+jzuz3YlRpyY4jyt3hSb1cb1gvzSu5IAawJSQqZddTDKnd3RARNBzIngksN
E+m9ouD2A2RhXuxvLrNYhzKYgkIxGLbmnf8Q+7iUueynhoZA3ySiopNi4SDqkk0ZI4wR7AoZT7rz
BruLdinL91jqG5SkOGqjFLrJNr9dXcY6HZYI9SvKx7C3HQfV12m4zeHTVRiewm4vFJTnXxBqU/ku
ptU8c1L1sqfTyf9Pjkzp2WaRXB7lTGa4l+u5MLG3WaH4o6ZxICUqdymDmlJcpYlOup/trTgGc7wa
aFNjz+JvGDAeaTXGNnf/+AzfA38aesLwKRcgFFlzmcyWJd9KyWuVHoyJeMOhjSN9B6fVzZDfFCKL
BDCoE/ugReJ3VNEkYUaxjl7D0N+TIVX8vqEuuIIAIwsLW3QB+68BS9aDm70oXqiLM6aTwrPRfxeE
Wu+h2iOZ2UvtuMieNjUHds2OVnBKI0mtD/bXTz5UwLVbRRQcvyL/en2oMr7mNFdJhmgG1B086Wlo
VPgyISHZQl4LOUfih2nqc4S+OCG/1tT79Wb5I/iHMcZwCYsw80RYO/XplHiRt+MujupOY2uEcKMl
Qhx2XI1+kREVhl6mGOl6Dpt1Drqiz1pEWDxzVQNGkXnrDj4e7mcD0m5mXTDj687i7AMz2nxuf7Nq
8rHXpzNC3MpmaIsboRxt8QkU7qQRxjyOnxrsJ2Mt1LasuUd4kRqkQdk69/a5d+4rfEGBQDZtqeEA
90tJb2VHcmc9mUaZw/ZFLCgRpI1FWrMu+LwOslQcS88SO0xdOvYtRDrtif23lzv0Av2cqiQP+/Ea
4brdUP2PHF2idO64U6+6WTBfMNkk6XQsVGhRd7R5cL+VUwVk5xIQDtjjjMEEwC1O+H8APZt1oLGR
u7X/Yd8RDcRFpV5HJ4w30Xgjgbzm4MULUU6SUVTaoCDwpiiBBz43D6JOu8ybT2W2U3pBsB5K0pVQ
rIH5mlsOS0d8JDiOQqQIDQdVrx6L+hM56d44fMYIh76SQA6t4aMi0vggskxNT4jlXbxQg2DUF1v9
cdZjSg1pZD8vbSiUMZiClFLqQV5xCDNKpg/x/O9gg9sILIUDb3IGWpjGuCcPpJ2O2UlBhe6MBIuY
ZbAQWjcHlM6q+xGT/RPcLknQ9y+Xsv/CwtNmuesOpyUJkY3tGybCVnyqfIQD6jXfqL27oFceqDzM
HLg9hVHTpmXJxj89cg8gC8+7+wejOllD541MDPyakh4430cAAM7qGvXEo1ZJREJyn/lgw7yN2cis
cYFWrQweYwxgRM1JD02BnfuMYnq/+Jhy+Pfn4xLDXdHCu/J4SiGrClg2AygZNK+CNB3D+9HhFOc6
cfusWSA5YYIoPbgXsdc+y0nd7aUjaq34cil6xWn8JCDoddMdkutk2Xz4da74ZETU6VoRJDKpCwnD
NJtXTYEOTELiNOUnhksQ3F7NTn7Ks00ytxsNTAWqv9dm2kMsXtebMXhLjvPzkXjotwrvHfx8X9tZ
yhUIro0eUY5LmwBDI6YTDQB3riUtuViQM7EfJ4N5pM1sLBHxWN4pVUm0SD64TtiVpucjYYN8AmPm
PhdgON38FpLTpnJ2cpL7s+NhrMyEmW0UcwPN57Sy0+XiRONZ0/RocWwSfy8XcFURiMGBbwo+xwkQ
FQXLI5g0qfGnxqEQY629I9dXcoG3uIlO19QK+EoDfJDWx8xtiVBaoMVIq6S/OSKDRezTHuJAHdPR
X8yglPgbctatUTDDO8P019SRSmbstcBNij3PucucxCjAnPmtKzmjO0aUOPoXw6giY7Fmz9xLJnkE
JMo6nyovMeZIblSNAkfiQBljFfrOAAqoPDi/jg/h8dxfpGDhmkEJTnFBBS/9dQe80ED5pI3epAYO
UcY3aKYi85scwVNNOJI/SOzcVbptfrXvmrx3PWMXKy+LqlCP1lU7oF80olkJsUSjqtJNkGQedMeQ
DiibT1c5o1m3wdGU3ALXcO0J3wajBEQHo1UI1VEa7eZrGBeoIG8Zn63EFxYjHUhnBVeP8hZP5L2T
JNSHGLihODDQXhDxY7QA94ZKyk/LRl7TgymIFxnWmntXsRJJkBiqDbBpxsBHc2qZJhsBpUYFSvaQ
KaSTCNQhSpVSGCjrjJiWE1v1dUqIjl4iWdV0DmitS8OJk8njV7N2wj25jKsp4qBX7wrWZwCah/Qr
SabQ1wHxEOsB/B3puBwdB806yjEglzwc0mqA0KT/sE1DX6Pis95jSVPoxOh2nbBLo4jmpzlQqpxZ
Wu3J+6YAaUTJG4BAKqGfYBQ7EIAa56lLDpDXjMlcrsluwZJPf1+Llb9TCRr1ttVOCUXnhKR9pVCe
1Cfmse4yUOsh+DB0ICD0n2Ol5kPxOyFL9yF/Ad1vB9GMJj9BqMVKf6YqwEdgPEqxtrAi1fd1WgfF
iqRMqUJeIcwuv+dqaHn5BVboX9eR8Rm9AdpecNNBufsTuYKBeBF6agGNn6E794PUs9C5AyK7U9Bu
td2PfaO0X7jO4zV7BCCI/x93VTHhmHPbEnMiytJ5F8bpmpYESwY5mCaDhFkiBvXqN0id6xEC917v
/yJ8Mxtk/h05kNau8ebyKiEbwpTDEwpP2pCC23uQpLTQC5SPBrXcp/vJYBhfHbiKMFYHV4L/5gr+
FGnBnShGIlOblqdoKF1ZqgC3aPuGh4vzWseRfVcpXGmL4nt8qw7fPer2twcfiY4wVq3rlZkmUQdb
twOSOZ+ok2PZDcc+d39GxeBV7+3CEk/ZMWI0rDbqL5jsKm38/htWjVWbcLmxP8ETp0u4M+PC3keZ
gJBEcv8p/HMm2adjUrYgK6Ho4Ifn/bSW+Dvw5z9sizKZTRuvaLsJ9x2q2mvnPWTfrajD6+tAQw5u
83wDeOuyDQCzaMBlW0G11H7yMLUpNjPv3bmC3cQKj8nfrTDFXyjjhL3ol9vrnVVAOZmRPXPgZLaN
LANAYdyC5L8qjS3q2Xp9v0VuI844euC3nxIhJyF9e0zZcwSRIb4i/Wiue8hqRRtB7AX3JfMPms+l
+W5TvSez0vAX35h3a2JRVFyV1oKPQELiP4LGONpMOTI4h99sYvaTmoeVuAYFPSGNVzkmPGZ92vww
/AjvU9ySDmVcnMkEJx+J7aZk3+QfoHhAMEy28moGEnARBf3wyd6ypTpBgJ4vL1d6nkTaFmpKv38X
x1Wlv7689+HVLtRLvTS+0pmP8XY0IHBH0SQSrFVXUTFvoxe1LHLSLdU3JcvoMnP922eJZl5R4TML
oa2EWpVyXd/9AtGbmeD5+9/0PsAlzhiBrXdbVvf+BNKDiZCLALWI3axIy9BGgVojPdix1JwkwEe5
x5GA8Ri80Eb/9AeQlCVe99c38FWPIHSvBXPfpiZ29XqNpk+kfsyenVXa0ZgTywwhsaiZ8Y+aUOF0
XX0ycgupXcmxNnKOTdY94pKDFCeLT2HMsR7hBiJoRbooJu3+EeCYpPMe5Elz6WF/Uy4nrJhq62zQ
rwB/T0SMKSaxrI5XHxfe9xKmLWUbPUKTqL7N422ofsbxoD2nC03rsvh0hPk/mVdeF2UdWUZbdvzH
kMVeQ/jkIrp1p+XaEQrGhf8j4cWujP+S3zGccOWWLHGmTf5v6Y/0xrVlopMeN1SkY6rN/j0TpoU8
Pl53sz/gjlSicA4q9V8MtoZ22O0UpKU5vXQcbOdXnrNRkfkmG4QGPpBSR6/9/0UQ5FiDCkQcrQMk
5nhwZNXULlLlclMJcD0xq9RX93oCQEa6/O3tyOLG12/73Pk0k2gRXik43WjZlQzhZnASFi3uBFaL
375Z+7ps/7wBFh9R3IJ6OG4bVRvo8tEx5p4TwE8BhQrJOOSjoLmqhppjuT59Ogw9oqZV4ecq160Q
gMNAtRv//9PkyPYHpatHJC8Paed3rpQfoGUEsg8xHSxh9b6tCbjxBRwRBW7xHjbVx5LLwAcqButD
yec0dbChXHkJYkI4zVoSlP+QUOVxGwxR7p6XlJbxEoPDNS3KjjPYh0HabdY+Om0eoSsq5TAowK5e
bfUjHBOucgmllc6nYdGJOVdzCWa3ogsPLsePp33x4DxUHCG7C6O95nsajJGQ6pu7+ZSQAq0AFEuk
v4YjROCa/P2bl8zRK9wx3HqxlMmu1EJPx/tZrAcU+7FMocgrcG57l58UCueY1G8UxNZJYnHL2xjS
/4RC7X7qQ/TLy+vXvzavxsV1lP+oG669JFxr4pnfnhRmv0Zegc5HDTDSUFWeQoKs3/QvY47Jrvqx
D5BYVez6rcmY+PcF3xn3Ic7hIIaKqc79y+IzQy1c9jLGcs6RJXkoql6wBOcfM3sAWMGxK58h/YmC
SOw0UW4Kd4BggpAirAOBrQtlAG34/P5p2tvZXKgqxR825MwAZGhvQ4QIEvCxQSOtlO0r8sJbyGSs
aaqbXENiXzMDGISRsF0FM+e25ldd7ixm0c80sBmQZgRjO4QELVKv4Gqra06hMIZMu4ZgbUAcbH+7
kWneq6fe5nRuaLyO3978g7N+IXlpVYOqpOveBAj6RK435PML2+JZzqffWWzxDVwmd87fP/O7PlEg
28XkL3/D8dVwaspb6PrvC0M+ROVG1ylgPQOLXnxcPtgAndYaNXgizOGtB7pMtckCfnKW0EmKehqi
duqDy+g68JU/iHo+VNAz5jbsv6BO5EXgA5XPHfdWjwiplOzAlvlHE/SjwT1JpibgF2iP5ekGUNJB
yqcpabHKuJGjq0XoxMM2oLVspWPkt2h5IvDarbZ0YGd0gLyF++BQu6qk6eIhgOxpUx1M0Z7znzi9
TphDCZGzbe4iqwbpHJsO/d/uaJ/Rb51zpa/MVqrQ4xUUTHG3iC/R26o/w/dZbpR3nSzp7tJTqE/1
Lu3/RPvu1JUBbMWUvxVE0Rr0l9w/snUB5en384RldHDIkSJ1UotPunohtatChJiVBF0A4X8ZY+O4
tw5DxJAcJdkQ3UfqmyjUuzORGw+85l1odNFLJxGGJA4S/4Wm69+LF+Us74KLxQX/+4030UqLAYC1
8SPGuGwewelKlizUVueyf4QHFXNnNSAfoGUvZLd06kJaHCpeXo4wLOztCEUAS3i4lH5fYazhtupU
XaRzl4uoLtF6NBmfK1vI2PXQ0urjX0k1wUp7lh4GrpzSgVMejM3RA4S+Ij5Y/xuqhg5KmLkpLcDq
MGo67KDyAwTDHsTWX8bdnTAA9rnnW63jzh5Q1z37NUyFPchmFZo0sLKDsPzJdCXfcph/kyxH1fv9
W0L1sQydxNs5sEwryEhxVIfSvW4xeHD79XMQEf0nnuKeVRMUscrBcWEye4JUPD7ZYrEj583bcFYx
Uak12xYoHXCfUR+IAL4U/VwTNHz+mZtUaZ+9OfM/2wRE3wGofdYDRmSOt4T/wjaw9sqhlMDc6ger
EwLluO51QPbetQTQeK/hbLhMoT1xShJ06mD5FKfaMdt+FeaUCBFLR0rz66q1U9QYv387ThHyqJqy
VUgocFAq6AVbp+gUJj8OcfPE20b98PD8YaLQWB7CHoREI8wTK4y5hC4L0g1brkfU/edrdVIQW3zA
/hM9cEniV/aL7gFW5XJdvt3d78UNCBJle2aGSpJ71rpTMVT+sMYitJgr8UZn10GFf7dZmwQXLX4d
/qPeKQ13DNGflveszfILsrsMC8FrFmZVxdY7tVLwydz/CVW2J4NeW+Xmxr8vfZxpHoiEBdVDUCnb
QrayAdpHEYRxtjbST7n2DdoPlbIn7Q48RlN3852uRDXMYdwQL4OXtfmEwnCvByM0bCai9QWuuH+n
XCDpRrj8XIM6Ij5uDXcz/G2yRbli4ChXPUKUQHUKxb9SjeB+LS56OuwW2fFe+xn6nUYJWj7aEfO2
psdsn9+3a+Pin+iuX26Ogbc1cCagt4tCtHrLmgwm3LiAUV87xgpkKdsE6SmkYQeI/q4nuM3OZVgp
cEtR57ApKNT4r5RpriW8JNu4GW1esEUwYmHAHemlsCnFNieJgDReKB2fPI8wV56+PAwYnCXEu+nA
P7knR6+wv/Gzb7hPtARPBKrh/QttlrCE/VdbRYu7AWBO4ZkZztRhtVvvkBKicekX0S3znWLgNQPB
zio7DiaUwmlzvS7HsY5KtbB8NdVGOGGb2OFeaS90iQQn4z6bYgCggROfIRQCulbOlOziLCQjdfna
3i2aSZI0vXjxZK6ArBr4jFWl75Xm/ei9AgQ+6DttIoo1pj4uDY7WiZi8a+IFpj6+V8a/kx7wXSDa
JScZiDYmyWeMffoecXFCI3wz1bjFV+SZqWgyn1bSz/mybDwz4p4NjtuJ9ioe8vsqfQtaiWF4AJ0u
1mFCo8E+MYLUo5BvkbofNhIOm3+IFUtssbNLpvlFRw1Fd64I3rFUkRfnjGV82VoIJ3ph5FTa1Pm+
B6Bz+Qin6gUF73LS7z2nYN8QRT+o5uNbxI/JZc+CuA7kIPflDVOqgZn7JUzcyq7SkFqPGf8qeas1
KiNH/jmYzJiRFsC9qZgjZCsNkcrA6bJXPLGrEAp7eL6rvqWZwvMFvbKOk/I5J0QmCqRUMxYE3wbi
3TANBatjy3puhby3oP7K7Pv5AHFkMyBnq4+ExZ32TkOd73DP8rSxlkk8Df4SqwORv8IRUc6YAJvf
zUhL5L4JZ1s2su8z9AGXaAAj9yLoPj9D/R+yxtLMm7UXjf0Tn02lWKGhP5lvM8A8B6EOAAWE0ZGL
Lt46gWVfBCTkT7556xDAOPrCQFtXE1uopRBYsF1PWn70dsn9tUrc52aPBa7HDIXx0iG1HpVHzp0S
IwpNgmh5oUoIYMgQFaoGcE9tmoH1xLTkjvkT6oItmxw2c4qQTNmK1tOLc2GMdAH0q5j7TpCdktHL
JU9ObN0egsf63On3FTkYZ/VnwZqbNeo+dnAOGLlPejh+BjAfUiGOo4AR91G9uOdi/+28/WWMsVUG
5Cq7w+Mo9FiaYcT379LSTJxbiysvSnriPplr438po+IznozJnEb7JwT1azcpWNZ9fvhtf96Bqmg3
cWza30H6zNyTCKPg8xgkmMshw+3sVVAD2Smh/ImFlTy7Z4++CWv840BAr+tCXNighbHXhhDusW3x
f9Szrd5LRiFKC0/gvFEQRXDgjqYTTmvEBrv1aSWGrCaS0OV9RjK2kdS/1lX/zYc46uZpja7mlZxp
JRDbI/NzgArATxwClavYxddfV7ioJ0GYt9kl96d6uCElDqTlxKmd5xqxPKTQE8qL0kLVskBQ0ZSK
zKbgsr40qd8ivwobQAUztqIM/4n5R2ehu1UddAW1sBxoiBY1ByvRuhNTaANok6iRevm1bygp2Poe
UvMvr+HNEhdOSe+wKiAbZIT9+HW6TWcSfEUe565Z2wNsfwvjrCqZ7B/ztB8CWga0HJt2H8Rq4Zov
gwJRRk6w9s9mXXRI23a38D0fYNamM4PWGEGgjcx/XStshmc9YmNJ2Clmm0xqqeVQuvj7wVesQ85X
qZ08cs+ADqZHIBuDWEC0Pk7V0ycXgirodHIZvFMI3NNqUZq9HRoOd15jO05fsy4hxT78/Qp6KySt
5uGrVEYOUVIUOKGO1Z8jHFeOx2T/AnsN0B/A5YG6LzdU7/QkkYBAHDgmMl0pD4TduRqPVunJ5Hqa
DTk4uqgUIPuZz5iRET6/tmUnIsiLJooJDFQq7nCmUkWLsgKW5OtI+GHo6HbDu0hhshJbX7K6fnlZ
wdZwyo7UHzswqHpyRxF/DWVCe7Eiuygo8U7Q2C2OrOMsZ/EQqZSns+LFrlww1elGgIVcfuhebqGd
qyjcMj3iwzVAJDL6Jq4S+GZChDetARzSker8klk+/D4QQEPD/HEXkGY7Ka0P5EbHyDHH1BLPbVI/
sv0Yr1c/5tVQmFrzXhAsr+TS9BxvkKNNZLjsvJ7Oe2bAMVzbjzbFCanuCq9KHvK0kzKcJAh94i3F
sko3qli9+RX1kp8h5CyERkQ6xTScmPTUq7BY2M99vM8xQnGGh07ufdtgTw5YLw5td21JbRsL513m
GHkk5mV6TKslmcLUMdsBiQISb0rLhTa4//PyOjvdPqcCcDgBix4uh3KEPb5XNcBox4wVlO2IRh7S
m+Ap7QvJJVXe8oczu88KMJ4ljMrWszMxmThBIlLfj3y690m3cKCEQ1ad0MxH9DkQLAn4s0nezN6J
DH61yufw2N53BXvg4WU0vB9zMXB1uranq00JpZiaPZgZRzJzUwb4BPR0siY6cwOtXDjCkdY14Lx/
p7bmZY3CqfMgvMcFAWewZO1SmaPC0D0vybKb3Q1E/tMWp6a1qT8cCD8dXV/vaZSdP+mI+1igYY0+
c5Vdrny1aFI6+8fYreGFAbPtibWfhnTI28lQJ/+9bWIOHo17Ub04rQubZ/3zExtJ411S+UbbzLRG
hsstxmfyWZ+Nyd3wmd3lFHSrnuu3xyxy3C+jEIh4UQxwlr1wpwSfCs2uJ74oMqGH0yM/bdRU0l6v
uI4u40ZQufGbBNn3z0Q+0g8oAVPlHkkqtLItBe7hNYlFuVpUxp5aHnxZEUn61C/Nxr9q1RCD/yZE
kChEo8OMUAD6h/Cb1nlAh2L0T9xkraIAYhewiEY8aROVrnXxa769MNvAXSIW16vELRWkbJ7+GqnY
pYXuhVJB4Bn85PXU9j9+9iouyxbbx11TksWB4cagAqRJibnVQGu1SrXyKMsobIaXjTyO+0le2E/Q
xpFv9rOdWKf0InQ9GYVO3y0ETAUVgdnDgILt+1d2RsdMXTtprOeDCajTjQMsWwEpzB0vDCkszRb+
xrthyopd25Jx+vEbX6A3kjrsUz6UBrUynJL5+nr9oFzSiGaZIuT/zy7kxXGMB/fbSIPIqyv4lP8t
CQ3UM0RTiHgL+4V2P4RxpZeiA2PJxFmYY2yStXP/So9B/NyBEbotVfhjJfaRBD6EWzKotOh5Tkm+
U70OQu1GZLdUs0OKzTNZ8yQ39Av95dQ7vACFxgE4G2WQkf9EWN0Vi1kyZaisut22HF3eVn0CfOs+
xvgD85EKYPm3CfJwnuMX4YZuLKN9ULHIARG8lGX3pOAzqWHOVxPPiuDoHo4+Wnop+u9dD7y68OMF
YE8wMiiy8FgxJLuCDQNkNyAwHA2FgEIrsEqJB42f00gEErT16X0ni0ZVQ6qF/Vd4A/zKJB3AtdvN
cw4U3X7FKvYrrBtaDdy9PVmBaSP4ihWAAkV+jsJHc/nHjRdhU9wSYTm8XvlfkYuBPA/guBM27iy9
lk5WLHBmL0Q6YbsowqjXnFaIarMptG8ru9VyJk4rqR/oZaomnoB8PYUpMu0+H9v1CALHFFsC32hc
XYvvc3vIcYh6kR3x9z45iC/8dMayXjaaMi4b3zVl/PlnKzx/bMM8oRrDAoBVycgswbeGnYK8TrU7
dUilTp4pjT1y7RNDGrCaKUIlgEa4WWjcqYHlHQtmEmH4XFTVaLMV6CWRjAzsMbEYJnrVdAa321KX
I7UG4MFKajIujs3SLdIHdt/oPTaA2J3OXkbtkoohkoeRKISh2Hu+t2oT2U7uP2UXgAGcLJTopy/6
nbkdhvi6Z4Fmb7+6/mQUv12cvOKDfeXyNtEJ/Q8jjGn5PtgU2WsRyK2Pu0a/qIYCPiETX+eflS5m
oN3JYIAJdgNy9Xmgz1knfz9sCTAOrZLdMSOs2Xij7Dg+2aeGzrjU3oB3Bi+2Y/Q9yJ9/M5hfffI8
mLQD7AiCh2W2fdI/Zmtu2et5yindIu4lRbS63oheEhQh06PHFKTiQJo9W6dYddT3wZQjwy2JgVBU
QkctrxcZJnYBCn6Rv75BxLHxn226YmNKCJG/lJfBSS8iwRXbY9Jv3GwiyrnCFjeEbi70jwjIxTMH
pFlypa3kAovYgJT/CV3gXq2Vj8/IAXvwOO5kUXs4qmReVLXw2WUQ1fy7CaYTBDt0qihsx4+E0zh4
9A1qf6174MkAN8w859/2hwrlLNAjmyCr+8CKQDucfS6hdyljrxEp2JK20u6kD/Yq04hvVuBQCHGF
yc0nIJ/mr21Cll8uOqrBHfTW+AYk7l9Cwh3SsTjdqIYIEoNcDLjRLoWzaP19YLWbV9fembeaQ0GL
9iLRSiIYNPzfPDDhXIiGrCSf/MdxJdexW4bghdp3sOpoGux1xUpS03oqz6j3y9ESq7aslQA0Ln7T
e5Lc8wxryIo8stnFQNfar0mpRrfpyZe5Q/Yfl/773pUjszUr+dCyiHFjqiJjR2FdL9aYPED1h2sI
dmo4WDRFJejk3/iJyCKjbjAMiPnq6nIO0FYBU2e97FH10icusDn5Yp2+87CQcFNCKjYRNuSQjxqu
nxptYqLOq6jPPEwoSeeDevao0olKPDF6k8O4F/q2hZ9q55a8AaDvigpexsVt4if7/KmDRGmWxARY
0qxhbL82ZfGXE23Qkr6Jr+yYN1iEikjTcFsq5rw/gXbmcNjlZBNO3pQrVaAV/dARA8q++Sz3lr4L
y2BgO+PzbZIiKDi7VZffRT9UTDBEZYvkID+B9ua3kjNWGFLa/+bx6kDZ4s5Tv42oi+kDZv0XNqZq
RyT6i7PYJq2SFmGKpXwiPxI2rh2jIPWMdIAnBlK6FpdZwfzWDBz5aL3NriXPwRhSWH0SdGDBkxKc
32ZhVapawntR1ZzF6+mIacHz33QB3iRvcj9TFtb6oFcs9OcD+6EOAjJ8mbOx101cEEgjiqbGSukB
TxlpNYwmPeSZnak0ObZJ8W3pu7Fz/K3N5lQL6CmQowEmxw+VTg/i4N0hdpIaUoZdErAFyAkqLDqe
PTka0bOBTeX6Ma2+dxPCuBQJY4snn4VMI8DcTnRm1gzMMKKUZ9XYPBbxcw5QyQn4HmQSQylSDSS+
dD5S4Ji9t/7K9Ip4lhRPuECK/rjmjjRDAHxfII18gE+C9Fv/TjieamYHZkRcxxP8IZem4oBCBKFx
zvae4j0S/RhAP/x/dN3trjZJkYaWL0Hd9b8lCt8C9G1WsTL2uEFALfuONL0idUb4Zim1TTKqOUPG
s2Di7tC98bX9D2l95fOQ6T+aAJySHgws0d9GOpwXlCFs3NUsj6XplRAvD0EYziiDqYdZciiZ2b7w
vS7nrVH9wORt9U6UD+aM2na2Q7UWDGJ1zM76lRea1R02J6uI6YpWbwySUN3xKlsbJkgBXP0R1iQE
HNLEYG47GjYW+TNfKM8tpeZ7izt8johup6Kr9EaqVDmiVD0t1kQ2hRhV6RJVuLl8Qb8sP7OCDTdD
kPxgHtzRapid2KvDNah+IjIVdVfbUbIUDKTYcCauZiW8eTxaPTXPOouqKIPseHZ/VCQV0Szp5WTd
ayYzo8oo3QJKMZ/g++0YYAMhYQSu66RN1/YIvxtA/eijMq4XidovzgJbOUkcGiT1naz/+F0GwQ7z
5GICsfCcME9iKjBfJzryJFUwij7OAjHTAQQh6iNs1OP+ky8+quV82OISQkqSMZ7gSIJ2OEcCBIwh
UuXUzvzCliJUU4fHwexCbF84JihrFT1ORWprZ8js3lE0yUQuP2w6lytcO/iKOG7g6loabZ0xt4I9
GTukNikxD5ymHsTfUFJgLAFyGXkieYdetrfRa9e6yx5pmv22tPr1g4WTKbJ/O5dY02V8++NK4Gfe
93MUXuD0dNax4Oj87qjk5AFIDffF3hIiS2xeIVGj2gnamQfL9anUebjOXo5UOVSloUDg1RF6vuMK
RiL4D3RthWsGZraosEkjf5wpw0AjbVyLJdL6+3VGX55D8UfmaOpoMcGJ2XEjrvytbKwVcqesL+rT
wgmwTN2luft+N5QSZDK6DGm6JiDriLnNCeuhEaEgrBz4967uVYTtPM9vagtY923m9v7nZpQiivsw
SwX30z3OK7oPuXrED0IAbQjFFO9nAW7m4k97HEi/i4OIpdNFtaczKKB+06DCeYA5H4dFgmpBKrnW
Q8m5o2WNWmxnll80IVJCPNsVRkYOG1oSUJMQ5jJ71wEh7Hn5sPNtl6rpDoGHC1tDByYlhcj9FCOP
NjqgB3le2RRBi8x2QkYHCNPIy/oS5h+Kc7Wssf29Va9zUygkNMBFRC/1ywdyp/oQiPxvxv+H5ldx
mDytxu4Gv64pJhmXsvIGHH4SASOeoJpmpxfUeaPz6272fAdxjlPmOcSuj/WZHwjGs/lp0Zn8uWkd
dJMfbVYOc0BE+wVppfrgVNdbHgnnBJ50baqshbaXJ6SE3WbKzbR99Xwp7S0Wx7BaUhW9AkAw8DLJ
sPjLhxv8+FkmSbdOX60nnhcD6XSHdkyoE+xkeou2NFwX2vZAnTmVaoZPxmUw2ifwaGTAE+DwCABl
KuxEUEOALFi3klUdgvujGF5ESBrfjRUwXomLiJBGTDhJuHyYrzeLfoqTojPw0c5PYvTU7HPi2mqF
oVLICrgn1Qw9AOJv5VA4AQJ/HvE/eOmyaxvZ5kAurrFQByPjrLgTp+GJsx3RoEJCtwHACLOoejig
57EFCHoeFkSxN2edoybFMIKzOu/hSuhEplZfNezFjZsf2pZ9kUZ0hu7HsQOeDb8ntpvRZdInNxrO
anSA1bPcPe/Vh6JWZ6R1g9e01O0DXMcocsEuwaTbgbef8VMhsCMg2mImewTnzumirpXY93OuSJne
ECH99LjkJhdj9v6rHAcegVbphr3md5cKZI5+PbcP0FFldUtyraZn2j5YqQzLEv3opbGQ2hKVv2OH
MAlSeXmKOv6Dj5yGMhnEKAaxHXmlpZHMfXInT5eow6YVkLvoBtgOL8D1ZA0AelA9kC3rq5RnjNrr
ogA3xEvzHA2DHXkO6x9uD/RVuy+TDrbEozQF/rHon2ZmCypyThFZ7gva890ycD4g4sFnZjgWq9Y1
CTboREpi/ARWDSzfgy6LJjjadkRAsu5A4dsfCWTT2SA+y+d7f3x3ENAIE3K0/+JTe8RsWJU995Dy
GnTjF+C6GgnCz+e0+uSAny91rPPA1U2st0cD32tGfu0NDO6A0V3FAvKHzBCUB4QpV7BpaFVlJuJ4
9gC6vr6PxQnQVg1iFttX66pVwVT50L3Qg5RbINneieTodpY3o1IpXBT6t7ZZAhqDKj/4btUwN+jB
hV7ha6dTBUnmtQMdS/8tk8V92es8pMpozSfd6x+517iryhWUDGgOiCc7NJC7JXYo8vqi5mKDnQbd
b2ZSj1e1dm9o9yoKSWVwUfqNmGlmoL3VMrIcxGTCY7XDEVv0xAQYCtv+d6K/kosdCepmWP/kmRS7
PSF91Z0WJnnM3k9H6NNkX3jqy9b+p/8JbwygzmknrXlZzLQGGiYilbVmfzd8LWMt33PrVPTm09g8
vBq5NgvFgnKqKtiKbwOBnvLy2sd8Zx4BDz0McS5Qi93X9TwzZhZC8/NRy92GNyUUqlSCUmNRPLEH
b5rQnav0KBa+h1gA/oSc4lbvw6lwshm2OpjC0JoyHenKl4L3AFN7Pj+rLUxvNvY4QjmBXbiYYSN8
1y2+LKKvh3SCr5zh55i6UJrbuZSyGrNPKrSdJgFoDhVxKgeDSZ3rmwixbOkeeF/OvIWoton8yklo
rPo7Z4bAcn4K3nhPK7rlJGV4hIAcNWW5NdZAxicZse4cwLbBII4cobX0b0qM5h9KkinSBeHNKVKF
SF2qSPmOZ7ZkIjusKUO3nyh5dAZ0KoyC6U2yEX4pOvIaU9UIB4N2OD9atuWePLugsCUMW0yS5D37
kSHniX/OSSc5cR+S5khGJBnlKHbOq92TjbXEljMud74CKPisvAa1psvy8QBm7zaGzRIbFbg23J0n
cy4vOSoQNo75+weoIT2L8Wxi78ts3Phnh9ltfhhLFaMVbxc7/Nl33DMGHoubHLCY70T/1F8dWYOR
qfSyMJqwiQ/65iwAvB7YXEpGOOy6AysnnE0vyeiX6S1pGWFlqNwj8mRXWqB4XN/ZPSfK3EaFbtWm
xJeQtFAzNnmIEZhqFgEDgkXjnUBQbk24sFShupXaECND2PE//oG0KuowENMDBY4W7dqBOPpC5q2u
FlL57tvknuu0PCCA+IGzu2EBTmkbDxsLIr0uhzmBLIcg/upbRJj+HkFg03hp4HTFJgjJVfB/qUqV
BXJyDuMfrp5T7bvrohD1xpvRG2iecq8iQ1MiSQTMvd9lhJR/xfsMoVV/b0PEVCOTsYTSHEJw4vP8
fmSr8PHw/woOw7jFFpz3GXTd/Ylgh2e+YbC+CQP3ewWHt6nHdtASXJw6f23ck1ebNrqKJ1MeSIR5
yXOYC//Ey9wABLblTCP7RfntI/Szb99wuxW+PFTVrtUEw87lcA72BAPzMQa/de03ILOuo5EuA2WZ
qjA3Bf6qaLqaOVW07Zj73WnyaioXgDftLlH3C82ASBW8yJBLl5ynhwP7xfZQg1TbDEyBCjLqoCWW
ZqTqK/5DTrvnDk1HCNZIz+Lg2GyMJtI+/on/2LK3Y4BzMgzwS70dxTQd6E69sbG/6ci4hwSBwPqI
rmTAtGzjA6EqXxVMwH9/aarWMrj9wJXW1H86KSYc6E5gbvLGk6CweKSPBxNmhry3EcFG+WKWEnK4
dnytQbNfauzpB0oZ6CGl6Hqzm0qz/djYhU5Tm0Skws6EcMo5UjhdvgkJgYBJ337uTUltjYYMaGYn
qpvPFDqQF7f7rI77NEUkFNpXrg7X9wAxna7HGoJBc84SXP8ujnW036trtujDJhyN/t/0rmoNcOyq
I7riIVUlOUsuOdy3B5JKn/4eTD/H7gcEfrgJFPTsLD8VUXjAO5gQfEHJlSpuD8R6o6X1rzFbZxAH
SUZZGV5ACtqXN2dj6c68fMEAvvQ/bjB5waNjXqzPcCyo/K1f9j4QzN8Zl+emry9ykV+KxdBUqAhg
bAjXv3Gbv+QLR3lD3z0+cdVjb3Vc0vJmUjj8yOw27EkSRRr9XDY4NZ4IeMI+sI7w3p21svFp3+l7
Hdg50o2XYh4M5e6wTc5jd0LvBpzUwlbYwWEEHih4dDMlh0Zd+mKWgE+jLtxQ5op0ZPZIzr4jD4tC
Jei5eIyOHlMgdHWgn5KUTL8/lWgxpTZzk6CIJZe3+3S40kQGhqmuXkchxqGeKoJM1BYbBVP+LJcL
+tVv1miioM9yHyU8wTl6yfexOsWcO6pQAYwYTUXUPhtQPI4a58yaQGTn9A87kDpiRfbqHM3BqkDh
MweWmTBNjK9QWbI8E3VP+Bc3VxLjSUzBTeV/reGKaMhePiChQlgCF20KNXTX/olr9M6fqw+oTZzg
NF9HjiLbo3++yXsN+JyvxTck3zrZVwx3/LWqb11Y8Rb/YyM7+IpzNWSwxHzIGKpr+zOsPobO6u+k
FytdrILceKzpJbql4HcsGp5QgeHDTlmBsGOfi2TTU8H/9Lvk/BfJ58imbBSSOg40pw11Npq8uD79
eyVwujz4Qz5B6MabN+dS3ahWGGBN9hTWwqwWB3JK2xpz+Mi+J/6vLkMrLSnqx2agRyM0YaTQd62R
VoYKuufz+m4CviHNICsYgXANg2ewgcLoCTnvecf0+gnSHDJwy7mjUiu/RxdBXapmEo/1HkUpr5Yx
nfgaxzywWEHqrbhSPleiA3DXLDVLUZBezNe80T7Dn43wKRDZUoYBqG3wXxvpVTwNjbQeLZhgV3Gg
otP9TcA6NSjTb7+IkoeAjFy8vNprXjQ2UaWfGoQ34NdXdCXUE8XScCE8aGf1DYfN4PIbqOmVR7E5
U+IUdD9QByFRx5tMArkH+0H1/J/4fo5IOQMuQPJHlpGvhD5i0n0oBM5t9wWzZfDwj1nh1WKd+0/d
mmiBGK6rqePBEugj5QaYEjQ186mWYRtMztU9S39Vbm9i0m7RpIv2evGg5pkdj4GTHlNoEsCH55lG
Jvrf1tmtRPyrtgGY95jUAdLfkdqrFjqUyt541KY8oYHBU9hzJ4vnrj2k4SVBHPkj9ba9V0d0Exhh
s6iKc14s9LsB5/IHBkhMgQr55zsJGo3xRQX2hd+4njSueW6XCwSs1KoGmusBo1Wj7YdZbWoKTt8x
VEsSwNE0gyAL8fzmjunclER5YAjE75/jyx1+e0C8eV8bs1dpCK7nDi3dXOpU6MlFw44tBlqd0fPV
pWSebt85urfFrCBmtUr6JmHdEuy21ZKTku9Znlno2wj1WdYpI97yagbEtr/wwEoiPyvF+JZ7/kZd
hcyQREna5bwhCAkt1jDUgUJFY9E+iiwNm7zXEZ3kVmmhX/rq5Ruuuvdt76pPutS+2pJo+MAl6C/R
J8X7g/k8LmXr2bdep0JBPKHP9EqRK9K/okjUf3Brs12xpLplsuVlnbVHCjdbEcPJO1Lhw0Fu/BX9
3Kfc/CV+ZuDH56ORgHR+mrRWNOzCaXIevJbffM/b8k7D5HenXwpmTXtnQFU6e49O9L1J7Yy6iwR0
otKkkQnD5zhs/jCpFH9Nc0iaBwFvnxxKarB9KmULYR5C5bmYIWn2knYclORNDDD0o84z2KIEvG0A
gbAhEgHh/hY+1GnoPO6zEOJeZatKSglbPJRYoWkArv41xfqeqf49ZfB39V+BFXfkzrhv1W5cJINM
AZoGHF6DqnJ3RfyA8RPwngx9+hSKqGWACpKq6n2dsSHEbfsaNte5F84rmkX8bN76wYVQ6rCzxRau
O0ohlhnnG52jXlAUmDHZl8dGfojrZK38ldVhKoNxSftaQdpCnZWMrh4ikhUV+72cvNoWZh2HHyFt
j/oz2t1s0vvrMum1kt9z0/DsFhLFnL3MW2fGPTFeRxNOA00yfYgZ33K0HP4ObHacZV77/xEA2BrL
ocSvBzXAdot4C8RwXo8yUP1+QDPBQum3tVStoOzUjQVUtT/daslL6EnHjrHqKZuIRifejVyG73Pd
naua5+mIFfw9Ujn5naJF2MCASDia54Gt4hzQDyF4o2/KyHKca3HECmQIrnZ85QDYI2C5S3dTV2YD
70VFKW5UyM09IrY7s6/DcsUOnryMFCwhV0JJ19cYFXntZ4mux6pp9q2Vwe1F95C+dahO9pGxm+x9
B/O8lgQDcXnSTguk6Mgi48248fXnlPhdtnXUv9vmQVybJVfW9rtr7wIaiS+KRlFm0109RONeRQoX
5zpmm7l907hznSud6Tg+2ihh/zXPOBw5UimwDmcjcjZJReUzdDvJbh16XZKco4InVphRV4oo7DXS
3zQ0+6nIs1wQ0AWmiibunK/d3Qb80agVNhac+mjy2VWcwY7bkuVuGnnhHjk9LUQ9lzChhk7d3nJt
l0U7mA7iTlm3fpjLWZjt7pfcaHZCrwI9KeDJL8ihKuvVk5Quq0g4Z8KjLZ1WzqLB/T/qWot9EvKq
wIgIuh7jaULcvdUg88m0sWCFHX4Pk7QM8Z+YRfzy1FS7yMnVR0KZ9UAD3aA34RW94pCipjPDgYlN
HTXqI+M2ieAwumSphJ/Lq74GHv2lF9rxlAuwKHwEYz3XN/6NgvBBKUJJniIUo1RfH3RR2aEAjymH
GTeI+utL/p6eJKlTY0F8H6vZpuKriWSJmnq0teFfiTCLkd7puHW5LGYFFUQbfr9Br4AWsO8lO1mL
uFzwwWXRbdDeGfUmF94yK+wvZLhhRXNc7sqhqqjLCOdlq8QZxdX4hhOHufVpOOz3ARA/avPM2ejl
SNd+hAvvAcCffRGenKDV6H/7UB5kPtSLw4VUNDja6GuhlrzVtKfxIEoThIw8q7R8A3vK1gHzIFOY
+x4Qy5oL4OsCxe6gdGAFGRuJkELA6AkuQcD3415sEXO3cJYGyoyb5WuqGAaCvsbWBCPCQYQIBYXk
aI7DFdI9wsUBAUIf2ijzRkXyaIP0VRQuH9bsOyDUxMLTmonfQDIWTv6u5p5RLfIqEazdLxQdpvEA
XXftbYTQIYfg8N1ykRgpGrc3yzAbYh4yeROpSonGddMA5LM2jS6je+SvOjjtydoT7C7ic7trTOzK
IuemC4r2N4WFr4bkDV+x18sKi3a2Ce8lyq5gTmTRWUvIvpvmwiKBxZDWzLojBNBh5siAoVtbhj1a
vn+7orybHc44a007ZgRRV2UNTih4j/PcmpcbxvDmbwksgQ/SivIoIelMNxXhtIqqC5u9oL18PJ+d
UvPY9B2whn9ngEXG+oXnXGxZIHuV3VmONR7M+2p5Ng5BxNZ6PEpc1d7pC4QhA1233BPv72L95YU6
+IMUPxtGoBCqZVutqgOggPcd44SNawtFlUYFfOiWIb7rZAex+e+OyK4E/SYAirfuiw6avMBR/7vD
yCyIPauGd0fX33to6zLLRj+eEqtswBcL/OOC1MFjqPLbX6mQc0RYTv5J58GyPBrEs6d0vxAa/+zP
sZTXJXcMwVFxjGOIpEaT9lLvqSFmugHr+Kko9vOpuTGMm81TB1riPZAjO4rahege3blrCcmPQASL
uxAzfTsn24+iTnF9Lg2EaLQbQ9uU76Y3foIK3GtmtvZvfEaZI6BhbfTYNjDD+Yfu2TuxsOwXexmj
20Odqx7L0aTs6EBaiFl1x6b83Xyj7lLOzxF0+GgyvruWc/jT3owOmU/hG61b/8gsGLbfRgNvJ1xi
nL9OogLAd5Qe+iV+C8vsZsQYVyWXz1mdy5ZytgOb8zrNdwqFT4/GzAgrYYttiI2yKZ+ASfEoH5I4
CRWJUY4VCaWSAbJHYUXYwCtRQoSfJI5Yb3XPcDrJJVlyyrjsQ4/TjFLhJPr20gkOzPsok4EVClEU
XannZxJBxEJeTAzpy3MK2QFtlYB1B9f4zYZ43Z6Qf76XqGcp3FYEJnidGjX4TyFGm5V2GkMoFMfv
LcJ3vSOVkFciFoZiq0xeH+QhC9d+Ez5cWja5JHmn7OIiDuYxRLUA0+v9Ci6gLjuvBo3eWSntyd4w
POkF69EltQ8/2vk+hZup84rXBQ7W6qa7msKEz6rlCp0lBeZA897ceVoYPt6NgZzQEqCw80TYucx5
gcz0Mif7J2tTvzw/TMijX6n/Ttrjk3EgKV1a+FiNT5yY/qJgcKltzu0XX+ExTBi6Ra/90B/DuaWd
4JiLoWfYGfMsUgcdh0vok1mdTcHuRsxIWy9vNyxoPGKXToQlqNmT1AHHAFCYB19dncqWeN6nJ5wY
gjaoNTCjPRf50ODqAbR6/rLOMTq99Ofw0p3gVkEvP2LBID29bOzvNvfjsqIi/hXlSJmYIVtJRX4R
e9ExzkucPUc/ehCKSgYW5y1XZ4Dl/xX7Dcsai9FndSubTXlzZqNauVUTGkwszF0T+8s3pwiYSyPP
IN4eJu6cSwuvJ4O2V0C8B76rp3yUyy/6K31Sd+J54Ff4fhmgl3/9D1Hs8aAozq393bDzoWIBO0Jq
duunR8ZTT5CWcJ7BKEAqSuSmORDw5kAxdK8Aa0JaO3Rl5oZ7FLoB7TpSrExCazDGwUJ3HGcD6RZw
w7Iw40e/fJbVOmr0LKBvPMVTTMzorORUtcKYw6ZG+L/p1BYImpq3sXBn7gdAbN7dz+BLOXo3sajP
o62u0PgJpjNK5fdBiW/eNR0hDuWdfRThw+oGaM1ew89nJ9zQPc3Cl35Ba2eLcNmov8Zax02yeP4m
lMbPVuYWVf5A+Kl8CpFEP6L4jYJuVSRd38ZkSOHOWjzqinPV6y+KBq+l+lv3lBxPoFkHxbo1SPhG
o0RONSQc6paaSlJBglN4huYjNp+kyV0slWa31Z6y2+s8qhmMf78wb0J9MXgRRLjIAJnbjEPxbVUw
iAuWlPdBJDq3QuBskVt2LjoQjKFhJrHR2U+WOvpzGE0bWObsY8FO76VGkFINLqvLRY4sjFLyL/4S
LVO9EOgSRwBPN+O7qxz0EiXEp4d8UOEkFyQUJwm8q0vATdM5Pi0DVVGc9Ii4xy3NRTfck46mYtk3
VnKhfjFFrjtN216eJ0sfxXQbnFM4YCoiWrfbic7O0sp3wehGLlH5uHr+RCHpqcOcvNcZSKrlahNf
XpLIpGv6wX3iRakOLYKcTU73Xwf+xcrJkKxgh2xeu66rFj2NAPXa7YmMBzybzWbXshzFDaJPUeVO
qvAE8JdWJ2vvH4MLPNtxNioBDx4bAj32EpkAbb3Tw0KQ9hNn7D+lbltlepDdRPAZcDod/LpRH4d9
PczoVrOlMhLVrvQerczJflZrPkKyBCeO6xi3a4rVyZhkHK2U1E2miSTbiGU5AlVxmBdkh44u+lQP
DCeD3zjhELAeyMqdmATZqTlRqonrNHZB7MO5XGETQ5RDWJb4AsO8JeZK2Bng0HE8/JK2o2rmeUeW
6oGob1VQ5NGHCaTfcfnJGIgRUleI5K0Ov4eP8yeDb7ZitiwN/pLdiyP8XX1JQXEXcDpg19X/LsJu
rQXPMZKDTW6AL+KKHlsn4RUzh0TlQ1UxbXtt/wT7AV6yRES93WFUCTYIQv6OdPDUGO8BYIoVZAAP
nZ1c8ln28ByHj84IsDupyEuav88U89gs9lepdJRpdkw6Kkg1vxatXMl/73QsKYtI7AYMagqdKxII
yq5fWPcHRN/iQsLsYKGTlV7mxeoHSlrU7WNBeTlK1PwMFWuZNAKbXBI8q/pGtuQ9HX6mKCe9zBRZ
1ajC2bB+4a0j0pBiRjaFFkfqY6xYfmuUnh3PHAMSIoP/8aOiZ9hJFZDl2cV4bk1Rok0ZLb+KN/Go
2yuntnWuAhn/Akz8glI0RnpmLr/EK3gTBPPc0vEgQAwFvLtRMzDwUzYq8DAgK0cHucEDEKLQiDbp
LEj0+u1LyOGzvlpPa7atyy9mEey6r2U7zd9gnNKPJJEgyRIyNXdZIoFt/xLNKOS4Qv92idDn9PL/
hbZqDOhyrwgY560okEfj0NoXrkpGcpY7SMQWgcr88xosD5JlkG+tUTwaFaaQcjyZCw5QyzEBgyrm
/iHgPn+0ZjrbD4FTx238dWhAfUUvNJz1CviglSzRALEURqeouF09pj83xLYcwyD5HMO5x2AbN1Kw
kzbg4RTmeEdEXHaezW2xHTSiWXBxAeMJl+P/WhfoYs5qSVouJYJiM78puiZeBzDDdqMxsgLYZlMf
+aGIdEQqEgo4PavqmaDIKgaRA4/ZSK1njGYS8B98z+CTr7pIXNAKHIF6ptrrPxl9uKA8vjGvCf1x
K3qTquPu4hs2E9PX8V3xebVScUCbmwYErcGZJuIenDQCQZAPgvpjYiis95eFMb43Hd3v3Kst3PM+
hLNXKVSIeD3oimiihUxDrRMHhSme3Q/H+Q73+Rm+RZUQ2aRDioqvIQeugCG1tP+OXgeVQo44j/jp
i7K9MzcRsHI5umwZiz61U68MwJcGdNWDSp0ae/XvuzJjkkxGxe01zaYgINnNwhxsLWFSwNRNe5Ce
+1WnVr/mCC5e/T3uAbiGS4/d/awa2AsKeZkvU4iMffAuabPUtpVUPEpnnprCjM/n9n+kqzJNjpOI
vHekTRoyDK6QEvXd+h1aJoI9/2aghYLG8LjcnKGmWQ++dMKFKWAIi+G2sQEx2gE1PFxIYIXcHod6
BGlPJDdaeHAlXBKd0GthnUqPFJ43PKjTuLSQdP0aAkdIc3yjvq1lFEPLZr6gxa9NRNZAZpKf2xVl
4mPVdoXl7tz5wkaqmgtDGEf5HM+ZfIF3ur4zMH4J22cIKo5a2KK4r+EN1dZIpbBrnS0e8CAyAijh
uxLDtXh+KTZNkbRyjcsWi2k4kAxuomepNcQIEkWBTLVrOEYoQal2a6cvFDXYDWTn5aj/P4wFPzel
IP4E6+loGF0cnOJn6Nz3JmyPMy2GBms5dkm+oDsoC7nNMLTd5G2tPP5Vm4hJFWkEHaXraZkYgZNx
mAXAlnGFOhLvCns3oypAH11RgSwEjzmBH6vQoVMdwBoRrqmJGvaLpVxJ6x9AnWsyzL8V6L99Li2F
xKGilLimoWAQACciI/9okunvz2u+bGMP+kADRqYq1y4YJsFbhWLSnG4lf1rktvfJch3elLcE2Me7
zl3DkADEwGz5JjjuCNj739dBDI4vWlHukuOTJy5bmu+00UbNiznsDjgQvddFOe3OjDWox1ADweSf
t4Q6dYgclBIYZMWKfwrKi7lZqQs4XZeR/wYuRdNXLYqKbNa19LEGsMFB+PW0mHIAtmrckuop8ESn
1egNFPak/x+ypaGVm4CHSInzGl8lZvIszA+2UBcoW49C5pKEbo/2ErVUknsacUtFTN1+mFbpPOVu
hZEwYhNbbxXxnLdNZycZV9mW1akYN12HF/3cnO96eoawp9aJ7/45xQ8BVwAspOGQS8qucv66LmBS
QCqj2zAitAAqupv9z7oL6HRB/b0MaGT9RZGrujz6HNkcWOU0RPn8jSXFoGl3kpYKXLPbQ4EdEvba
uqCtFVUS/27FLOadwTTdy1KCc71LxCdG0kwplro3bMJ387bvtRGt+CbzYOL83SJVg02+eSa4KKvs
OLewbFTSX5mnycY0KyKbgXwwbSDHXRMnC5QuWKAMb0RQ42plCIxCj0iIepKF2D09J1esz79+JBZK
DIWvC6pE1rN34HPG8s6QkKkJamDOlv6mcQaDVnGck1L5etcWnlWWMmcjKBr/ibzu0d2mTyJas39z
CYt3/vvRcj8GvuqsMjUuK0h0f07KsuF1z0OGT3+Tln01lNTRrmu9z3m33nflALsXu72aTL9K5ToZ
i3rIhJPVtO3EMqXRxAQZlYq/RNjW1mZEzM+JWcmE/p4PckLmzlm576AsgGvnIHwKunggiAQzFzoz
B7DqGKCzso3i1L5Kq81foryYkuTVJidVMZ5UjdRFda8mTA/Z+o2tyZRjTU6etzcoesHB73xo/1O1
ufiQypxOTxJJTtTb5oRxSqMwniGATsW8JBaQMFi6ap1pEHRnPTfEx9WaBWxnGkFHFVrAmbQhuBCJ
UP6/pWU+WvbsXVFafX+hDEGw/ON7qcLRZuqKlDWgraLlE9UDHE3dkV2FNf/3dDMLwC/2lpccy2F+
y4JTgEK/qezOTQL9rB1dEo4588a/Cc/aaByXKKvyMLzCgL8cjdlc6/lUtPrS4JPjliMIYQmxdL8W
f3puy/ryYFhM6+5ax1tCYeUha5d/5rfYNfsAAVSKVGA0yhnkc6N+zY5xUqaTLlQgS5fphbDkPTue
1VvIRFWdlYw4De2GcqcvJiHNcvDdB+pPtG2pc37ITdQrbH+qiZZ8JvXxYOMkpgKG7xYqWkjwYKZO
IWEOFapmdh8Y3odn6/2CRZpUIoHFLIlPbiHOl0SyYmpYmFOLwgryyiNCUgLqu34Yh/fsCCN1qM3J
bHAoKAJVi+nbH4Ky+RF+mbVHe/Dp6ZDrXEsem6ekf4PSgnihO0WQ0l67ix+p4o/gSkDfBW7osvRs
P6dXzaTr0JCWw2DRgZ5fV5sX09bCKw68ux0yu13TKS41u82pcQoMcIE5nBc4j2+QlGXDIxUJESmF
Gyn9sAjp99N9JFwmg59AG0aLMMHq4JjhxjLT1ZyUOE/6cmEKZFyBBbOPDnaTfUk9HTWyrovxUOYQ
cOQuLbQ0LxpB9zq5/QYXXtvTxMU59UzVGQI2sSmhnqP35df0SnAYctun5SG+NWko1N5Nl2YyK6lA
59+CPQDzH6z8gU8c42xGd+iO/qhvUEJ/vVxsBZy+Yk5yc1hHLIs8bXchoaVayjX8hhaf/7xwL3qs
eZ+L8yffZmqgAPrJztWUvvqKXMmO2mWjyT5mU4vcJy1FGq8mBs4faV3Y4olgUGk7RFjSs1ve1reT
i8mcwczqI4Hc/9Wv+h3nQfWoaFXMm/xhFIjkKw5vCeCP8lV0ydCXBOVNPJ2JTBCDgWDUSqCsH57J
rmZyu3tvp7c0nJ9nsS85X0yZfHz6VpZ2tZJ/gFx0L0AG6IoB/tsx3vyiHKWJvXE36zOAGxfK+TvY
fQz+vGox260wiK0BRJ07+s4J/twKh1soGq1ADYPwklIFTtp2Gp62j84VYJR2rt3WC4UcbF3E1o4k
LYyt9WWxPRDWOTLTkKCz6iwXAuM0yLRnRcMzlFeef+CO5CccJqIG7ffgBNTPvyi++VQWuT6FJQH9
D4vCSkUtg7DAVQQkPoPWovdhT8zxrEaqjmCXpUF981u6WJuFFFyFChUlibfc+HG5FcMHrdSbtJOJ
VXHTbDGssxFA+EuBqz6/UDPVLHWMbyKayVwKueJT6eYWQXoDskDOb5na7u+t4qbssRQ5aJuhOpDL
75J240zSAuB+fOAL71AG7oas6IhShvhQ+GE4Bd5YI4yUJzRErmXcp8DOL2wvcQnKZQpAmRL4n7dM
a2z5+tXGnAyCPLWUQFj9wtPtoiABcI4k92D/RAJfReU/ThqBXQIz8vpqPm1EX5oUwwzl1yIJQ78+
NgaHPETEH+bFBAYQ/SPbAHFQjA//t+ceewmnymo2N9tSd73Hof8lQ9Ctgd/yk25mPPLR93Q5j/K5
zKft0wj0inCZNXuIb9rK0p/Dz6IjlixgKRH6Bs9tk31HHkBCKjZdgMisAeSawTxd8nzOjcVwEfPi
6ZKue8qUa7Ve+NzcHFfnv3PjnnxTZIbTkKhEJU68ukWgnvB0X/Z1LtmmEvqFX3BBP5zjtUZ+npGc
/wVHILn8+j1Bkv5IsgJHREXOVzgwB1HLTUTn6/iicC+Qt+uC5tken4p49jrLphbRieAkgW8Cdi3Q
6RUuUeVGydTk7tKTfPpFP93MMLl8OW3VEYi4w/zu0Ao7eX9Z/H7a1HxG82NS5+fHyDpETng+tAeG
uEyj8ce2lL579aTQXvtPgdYaRHKq4qctuiNtEBkRuWoj8Z95PRYPVOYlWuuvsnvD+/mXok6N0iZJ
XSIBUB02FPy3BlwmO3MNK7cfYA7FBWKEGOmSfgLKmgmzhIy+7k6XWBcRdhOYkxmsH7fqyrXDlFrz
tmiQAXGVDJ0t09Mo6IiNVOySNvZE5d9uDKYvBJy/9vxQ7aa4Q7EtHq1YfUuNrIOASsv6+YccPGMc
IAuIy/C2W/49H4Wxdp9duKTKItmFFX16vS1ndPYGRxKS7gZoKHHcMuDMuRwECi4mlKWKsa0IErGH
lAchRf0xYVQafsY2R2N+AcTZUy0Q1OQ10AB+A3rbJCVBhy3ylXxJqncy6ZQxP4OKr4ty/HpeuD9j
96O9xNta1MsPxKms97cAIzmPQRI/Zgrpj/Ux5JD6usoFzH9LYLHyisOexh0srf2GvzBTqDjO25DT
Gtp1s+dcytJsqGAD5FIeCSg//ZoiLqOORDj1MCSEIHOOzrshTJunLI4vBUoOij+Kd1+QqHPQ/fTB
J8ojwyIC7B0HSeSE5yHluB6TAmXE0c91zGC3sPkdCztCOEmkOiw+lQMbT1A5o5hAfhxH8U0bV/iI
s6Di1cINxohp6Jk0lP+PcHUYQwx9ANdoaFzzouIQkyF1xCsy3jQEB2fxEdgd86rM2wkXwNvKYtNS
bw74qNa/7Ygygz7C3Y/vZMRKRKWOBpz9VpK2+70gSXnhfYIdUz1V58S58wJlkKYG1vwNLWeb67We
KHIdh/coKKQ5U8WQDs8grWG46MfLPjtOt6zU/KF1qAPVw5PojBJ8sla7eqR3BepTMx9ZLVEUIg0U
BIp5dZ39LaHuGLT5CCvjmexLFHqF8Q4V9ZOX99qp8H/Ik4qQ76YiUzVJG8IBdUrTPFtzJs2GcQg2
q7UVHnzLOfeQ22l88Oy4K5+LKJINOy7d5FD9QSwA948g1/c7AekaYPwX0Ou5tUw6a1SF/nx2FcA5
iYxhJgU39FltCtIYCg7r4I8XSNOA83XtmjGeIVGqLyNUEBzUCEr37vknyiMl5brsSLLqAvDzBH6b
AM30JAuQYYIpFq2tXHvdDt9Z8hxx2SEfGov6Xfdu4SRUVqgNg+eg7axHevVICKIPWK5mjk0gT7bZ
r7RZXg/GjildBXnuYtnDgRDphsTJ4eCvt4IZ3B/EyHBWDR+RW+hKaO76gAORZJ9rGIWxSm65tRww
bO1SkSGBmNzEyI2EdXK9DtRxcL6X2btqk23jhjJhoSU+1nlk6dphXy2E8TwsM61jbpzuR5mUT1mF
LexVM5LFJjuTzWeku720y4Vjtq2fznCsVY/IB0QSnpUGbbTofofSDkOvDmla894MZl1jUVp0g2Q3
jAw3bbxk5L5uTRga9eaqYVZ3Jggc2FF+gxAgpGfuh7B0IrfUGR+YTUb6gHdLxj1f8Tjg4aMnN6+U
UKbD8gC8dvih2SMpK+N3Wh7DhOBmFlkeyxd1xvmvDQed3ohWWpA3pfGot8klFYe0wyqTI5syg1gl
eFzDv67aT5AZRRThc1+5M1XcYzwKqjAE6gArAZDxFHY0HFOCI8qPL8yKglZ8Aez2FD7UPWfwnVxF
yXzcuFgwsJ43i+ZZ4VunyJ+5TDBsDp0arc9AUJMVJkj5sc6BaWeoGthYpcIU8Qn8NVVe+lOEMMaZ
f+bMKW8OV76WyHyEdBOIcoghSLa+9RLViWhI+MgVNK/Wn/j2wx7NNuE8NI4jdg2xIChSPX1SNg2d
pCH5/ql4wnIF/cm7WSVZNVEaybaOfmrjNF/GMemKcKgNweVTbZA7h81+ey60o0KTKsnnr5+EAhUC
UK8fyXM2Ki/oyd8QQsO5L2aJgwulhPbFm/KUxFP4E2MrAUyeeQOUSL+jl/lmWwg8e7S9cLPuVk9g
DjAwi50/4Xnj9HPifgu5Kx34CI8lvpNkonNJgrpY6qKEJ0ZJW6k8VbmrB8i5OiVs8cvIxCVRj7PI
rMIZZtRQ6Dj3X7WvV7gGTZHlQuSLkP3uxE3EF8QUtjUfFd/SGWIFzbugZVos+DcEyOmZvCd5nJit
leA8O5/1DoZkk6rFNhetn0ZoDse7uHlVZMTrQ51ONo+RWTE/6SDSlv1onKZ97xYuPsNPRszei42U
eVX9ACHo6PrEUMm4l+AQGRzbNiopAQ8DgBRUfOKqF+HzgacSJKC3D1aOWUzwhxhxog6hXjDcEekb
eMwgcgRt352ADzrSqlsnRevKtBqJ4icU0aAMp5EWV/KIPMyhmPkDmICe5ItXtRjjNP1syFurcJYY
3fCms6tDyhcOfLr5Q8KTV9EwR14W6ZpC1qMa9U8JgceGtvPN1bYYgOyjQDxzHuEgXPYGK8HX6Sio
KgyVKl3GKm/QaejEvzE20THxrlXKCj9FN42sbG+/oKaqWD6CMgj18jRLwMw4/ud43J3FAqoRChgL
Kdz+7Gjm+DYeVucxiry2sQobWtL0KmcRKFqCtCT02uHbIZ+ZTlUOCSCj4OMkFKa2Ju6YEO7UWlsp
+JBnbI+7aFKi4Rh01VLt2m1weCBjf4nR8l7NuMLhL5pE+qUyldTrCDuFRqIxdWmEr1W0s1dmsMpw
X0YwuQwvDO3u44ZY1bT56ixmACl/Xxiy4rrkbJk+KZ9a7SHCOOj1udUau+hjDcIAqW4/q9WI3KHW
1lp86JytZ+yohtDOg0vOim06kjX0t1DpqMu8xAGDoTFzW+jbms5pTE6XlDXsKgsuoGNUBn325X4F
1hLAVi5QaLO85TIcuNaT7f104aYWCvl1cA8TQduWk7UyWjjl883QXHyjJAuj7k+xuXyjchAV39Kv
Mdzy7mt/EniHFQSHg0jBp0ygLA+on1+hTt01EUk0KXPGZQ4VPFHghyIpevAU96e5P/CN5sQIkbtG
NVM35T6mhE8XcnmLefcFE0VaWp4ZCNTNcpcM1/QFlSEIL1lHTqSYSQbsInBRXJjVP5CcGQGau+xG
V3eGrdVyWa+gYoY/MGQboFLqYM368qxYZqw/jMXqGYlx8dIEUISH5DvaRTQMk7jvX/3WYNhwMH1D
i4o6IV8Fzu2UximUr7aQYG+/hwXoCrIDm7nAtMteFayvo/07/ykmu5ZwLUb9lgAXNj9E2Ny2bK1p
+VRfjmvoDV+/NTYXbua0+5+r/f/i9fmWpthA5yw6QMkQHfR4J2gHPaH5pfu0tjyaDsBot/9iDdT+
Y7tiooq4Ihr3Ie7vWGJ2zNygfYBVNz1+iRhVeXmbo0KUarVWz3qFND+Y5iccddlBYhT0sbOYksL+
ho7D2qbZ4WLGQgs7k2VRpEGKkkxucdxZmIColed8WFCMNZ8ql6MTCLFa50fB0ODVcEoWk+kvLx+l
u8RWHyHRat0OiuyrKiFKM8Iuwv9QdLSdSfuK+lAICTzTBV436QJYqmKrnktBq7Y0DOpEPfesPgAu
RIT8Ix/ROfjL5Vaw2UP1oRwZV5uRRYzg2qRmar57yOF5+gbZ0iTrI8mPuC0NVbMIpgxjyQYVlYoH
2PqHJ1hiNbLXjTlHdxMVE91g9yrJFdQf/wPVR5tIrssx+HZRjM1sXcQq4Pgoj+w4PgF9lW65G8F9
gnPEO7O6o8Cf3JSIViEfI0uj912d42pYVeduGvqaagoizWpjYSzQfLt7G9bmQ6BS+yBcK8VaheQK
cVFhj3Iej1ZjttFz17Lf1g/vhee5ZrbCMIfoIHB7H1Co67kVL8ED3uGzlAIXm5v6bWH2YqLaXtCi
ZnvRnKeEKAijOfA7u2GH8KMhFqNsRVPEZFdqCpWHx8opSbfNYx3Hb7M805AZk08ZqQKetvOjRdm/
5KZWOUGaSYqZRRFeCyOCi+y6fhlEV3EPx/rjT60EG5CFwib9xxK6UGLh3T4GLDqvlIvVk/bXzG9s
dYBMTkKMlCfsXC3aUOxiybX23ayI6bjl2FvOxHRTj+/zA7mWzxCByCo3jaxCYZT6MeBaViKrpWwl
xJuL1tMOc4eWXF+HW7v5wFsl+zL/aVjyRdouW8FYWQNZCXsxJmMC3Ofba1Mlw05ZsP222NKId8bD
TdZEOxKd/uywtiVGqY+OdXLXZJYrl8VMHj1CjatFEv7QVQFmd0tx23l0bn+OP23zRVlZ0+rh4XK5
yFfOvtgFoFChL7mYKh4hWyrINbYYRc29JHfdff0d/7PeZSGlsq1IgnY7cFD125kuJrgKk1pDS9H/
R/NsRdeUvP2IApOE7m5R8B+VM65IaUCgj/Yi92OXLYUdPFaKsDXNIOVDv2ULlaKQ7wn7Ny5cZZEV
rizHkU5ajkqg5PC953FDWmKHEUB63vPpHcBpYYCj2hVbuIbYc3NKkKoXKlitC94aVLKAkoFaBOcS
oolDoTXH7XPs9euMOsX66frCb9GNdwdjQG2RU1LSLrBP50Y1ANDMHmmU6V2A6bYAzMm6QElGpb2V
ClaTPzzqIa0ur77PmVqUgqNhZJZeg79FKcVZOOsVYDOvDACxti94SdGpJgQwLPLCqSVI94XCEW9r
786SXzzkgVdn0HBHsr0XO1WeXvhn/OOm/TGn7CELyfogrk3UC9OWL+Ij2KPc0QBbK1xLHqMEAymq
1f310o91ysoxHhq2vbicFiO15Yq1Xhu+Fd0o8Oy3JMhyI8n+tLRz3dOZbMn0T9obdH2sGWZEe6i/
ulFi7xcLhblporjPld65LQ8m0vTycFwyEac32eUt6AIrvX2XyrTTui1jEArC3bjdbHGk+VZcw2cv
nXLODf/t4OQnlGoDt4uU8YXykRMZwNTGiaC0EHdcelFjWxXa+W4Y5a0C7LOX2JSftWZyCnVE4Qfe
MHf//BK/V+WFvAP4PI3AEekYwmK10+UANPdqmwLpHPBxgCKDkaeZuF14Kp++beUz1h4i1o3ZFbZs
ME5V6gWgOjfnKrVFHX4iJ68ARUt2QcxnBCGWoVLAtvp2uX14I29cHxleEI0i1mZ2ZdssxAbmdhta
MhD1+Y14oQLK8YbA1GqXObOkMPZYFgOZBkybSRPbZXnM6e5KIyUgxITKhcpSgWlknycNdEVghwPY
IJ1ojfFUkIhYYjFrdL5u0V7cyQLtnyuZW1tWdEppgMqHBjpP+gnUPdpo3li2sXIzNOVKJDn8Fc/m
aJHJvhOupvx66Cc9eC8uqrQpbaSptmEwP0lhD+RUDo4Z+xfGCwDwa9dophq6kZ6UjW6GUKZ9b5zJ
ujLPEzcUUlKHHa9uya6md54jR+D2lSSH8YnmDFqwt9QT5grH4rSquvjxMZgPMh+Z6w9d30bNW2r7
QusG62D9quCG+OjRuAP7mhbeLMqSEcqe7yc9qXcx+ynRv6/cEajXK6f4dsgd8/fUP9bX2XY8Rwj6
TwICifQ3t+zJFCa192hvNqBGrJN63kLv58TPHZFgU6SaDzLIbMaofbpREH6Uv0GrQ+BiUz2SiXuv
4za4uLrksV09tcW8KnV6o0g4yOGTvEhWplgurgrzmxeYfshwppwrPdmYI8dRz+47s1k8y0firZii
Fs7R/Ihz2KNP7wxsu/MfKFtKTAe4uHjX/nw+szogexTrLooW+hca2tZ4h/vrpXEC0sMM0VVjQUWp
hUu9jbT/nKHr2EGP9BwJTSTBFTWbI1L5/iOUldbPDC4PurYaxHT5V2F8z8J3dzFIIFtiOy73Po4G
1vlMMjQYEca/wu7tce75qiOA2Vc2YihW87jSYDFGFGPyr0SzKH68qXPO5P8Fd7rnzTROQEvrSNKg
TVdcKgt6iP2BbeeZSjcyAucYvodM1U9IN7TWO0tsDLoqEW4DY9bXeHnXllZVDfoaoyLAVyPRVxSV
qmxBCkNpS4CIM4hz0iVhM5bIs5WUEibB3C8VsETGO4W+GGxgVrPl9ZQXWzm8dbqfKHWWsvLMdTd3
SLRBGAHW5ZW5fcAoXsoljUlBkbDDc4tN0TASOGRvrKV0C8v5b44IogTpo1K6T6OHLmnkhmx1sC/F
ldVwe1u7nby4fzXYJp5LXxMPOfMT3tq4i7l2HqNuQFqLL3WgcfyZ8JYoHuTpAOil1jfgVXYf38ca
rEbbjRAqiHn5B3UAKOuDuPBcSnNeJgvo3NWOBe4Fvk98Dwo/GmUzbrkpkkc8o2HR1suXOp1+BJDU
L2r6AundQrtWk7kyJ0jCrbOhNycps7QTmdex/QBnB4zsGglu4hJpYtFPqs+78dZSURWequONgDA9
d8K0NmZprvSluQh7dcCca6lv5rReTw44Ya5OzfrnUawoyRRkTbhay1lNoi4zvqCeB9puSaNjf+lw
unEZtEPG1OFswru0pnKNNXpAwttuqV97Te6kfQg4MqXOlT2EvVk39KirQ5CTdd67iZceVUoILckN
NDwHMOOQAa7xWGigce9+XX42yNH/S+Htnm0jL91Iq60/3utDDa++lq2qc9Zno237sDXpFF/tM6lm
5idxmqUmEsML5H1T+PeQVsVuGGzC0Swo5SpTJ+fp9riYSfhp1YOdKs1wYdMsADQjlXIlGWhZB8Lq
pYH45ZnSj/MgcIqNpDLeRGtIUMH/bWl8xXFPQGOTn7FsXahVUtK9KBdCev6wmfOTBQYg+5kDOhhN
70LcGDdc+b0uIH7CgGtEugS2BXFVsfSO8jn7v3ST8JVBaJh05ewBMxYw7i17lZ8Rq4pcaJb78gKl
L2zL/XpyTV0RC5A5MkzqtkR2BkA7/Fkdrd/dDkUtVQQA+n4boBL4agoTrIPJBn+D4kbCxkIHO13Z
bg/Ydxylhq08Ah8vMN82tawVUmhe15nKi8KMa9qgQww7+dm2toqBG1vw9GlCh+L29slrBpjDe2r0
0Zxhs1cDess88q7tUzCMslePnnh7pHPIewtFDUVMkRs6o82VQjOsjz6vzisKzTUfiYAaSmQI7T4D
cioHnnAnYAr+OUrj2NV3FbZsZ/5wU4iCWqOJB3zzATibEIqrS5v7FeExF5MD0MHPrWeCjh9PrY2j
py85i6grqkh80wvMdNLOZjfNlroAcaxjilrDRpJ0YuhskEz/J+J2pIZsQlms/XHdg7+dWy1Lvbso
GaXgdKqZKue27manF9chjfickwaIJXBg35zo2CUoUzvImwEtCoS7bRysApBNJ/I2x7iWDkJIVM7O
YHrEMeAQIQk4BvJMmlGyC2rzFRR5te1Od8X8gljh/PSTNZy+R8P3usjGsMY9XgNKJNibHsPwlIhf
xryInEPaEtq7waUOIFMcOI/8R75HthyeVMmOh6yiDumqbTusyVU1HVpcQo6fSv3LfSxCjYFa83oO
d6twHmdbRx9LY5IYPGshlFvPpPvkMrGnAd5KcD0z/durCAG+lP6vP+tdqgFrY8Sdtg/PTgSrlENT
mq1TCO+kRlaxjPXDY5haeGoOEdyHMQUP7UUQd5jDj37n9dv+ZJHdrLhvXaPIVoYxwQFGItDDQqfz
iXeihoFaGI/cvc7p1VmH7sMPlrjmIYdJMVuTZSy53p0m7qdE/6YJPfbmddSEUD9NMtKala2uCUHx
LPZ/fP5tqB4tNYreT8To2NK54dWyHnOiTqT6S3JXXC1Jq1XFqFZBOvpvljD8KxCCy0Wkpxo0mCVg
DAj+vfhOgijpjU3pxDhvGqUTPlP+jPhNYgxiByeOm6gt31Kzh8/0TKDoS27iffycOwS9pgBaZZ2q
Sqf9yCb9UjvdVDR8kHt4w+IQcWEWHqM65vUem00zXD1r1fsDa/MNl70gF/3sy8ENVAVKukRo9p4v
gXR1xWDfs4l5HcP2aBT8pT2DVWiBmm8Y26AoV5TYnPyoCP87FuQtfwHeSWyriXi3KN5EZ5zwqHtJ
3yEbPSuchxK9LLV5eCzGkGl8Io2o55v/0fTP228Wp42Yt1L5AAMRFdmT0CfTfvKs0Zap1hg8VIdC
pgJbff6j8g5wGVAubI6/R/Tyhq3BMO6Fes5qPOYH6srJ+SylD5PTxzZyADmZKvRmPy9Sf1Lewh7R
Qprvz984FbeKUtWD1PCSuRMA8g14rz1XbTeLqpOmcjSAO+WkawIppzJi+/UOGffHBz/WEPXaS7fN
yDcw1GPeBtLEe0my0z5CQknhih6IIAhX0Vom/VKJ80NwVfIy0xFUQNO4oNN1GTFzNVL7EPiCLUV4
dHUJVLV3VrneBAsdRAA786gwrCoEABDWNSaIl6LYU/hO3AFWqDQpztgWwo6qG0z/JNCIo7pmJdKK
aARV9pbA4aF+eH4jQMQYOPlE+Co9M4riUx10q1K6Q6c3zbNvegh+j89Qtqjx51sln5sMgb7xb17H
GilXqwZ7p0VBNEkZ9SD2fM1o6otht/kvYfesOCsF2z9M1gwFwSL7gVQkftpv5ER6s6Gu9UZcfYgL
HZBIAE28VDMrcwuzG3SGc5kAKRu8deT5hcAv0r7rWX+Xky8oIdVBfXEzTOGtHDrL/IlZdlAF2QUK
uQd0p/+Lh3eYG2W0zrnd+lizV/p8QZWw7Z0KM2WfWX5z8ameB5g68Pi3E9jDieY4Q0MDLQGGHpvC
mwe2Y/x22M1fkh9RpkikQDKT7ku85wlBon7D17MjQWk6+hVOPUCrxUmGvV1AO065T86UDu3oi/j8
d1Zgp0NmSTD/2E/SFnDxbZQ0j1IkM64HRxOXBlOqrRPlXPnWo9uFpxoerfAxpQ00cJ6T/EP7SCvV
yWIsEhkp8ksSL9CNYAAiAq7/8R9RykcwwmsNKhUUeLflL9paSIno6BFs+V2kVBU3iFh97/z1kBOf
ss9FAc9gDHlHx3tiuYm5Tby3kStk8yWyPLQ2/eFfhDyLmOaJoiKnKN5FpC6wdyU8R2vsffG01qJ8
8NbfyHV/nv0IZSz2uIjNHq0T6dzRiIjAtAYYwul9PoQMf8Ij6FPcA8KQVFc+d3NTbcTnmb9AmXYo
FLEEk8BfObX2GHKaNZEq3kmAVHGNLinacB3S3JDCqjzPzgQsUCQ84BATNbKS3a/L01I9sRTEYszi
lgdJok57wz9ljxjTzkLxRNjVddvd6VD5taC34lVSRobYnciYZWtq5EgBgJflY6GCuI6QWXhyOIS2
8sn/vpTGoBRSFdcsJO2DB1AgarqgTl2XcBRBAlelXnYpy9rrgJbO6cq9HNZs/EEMpzMmhbqUatn1
wAme0fTEFBwkmIa2GxoZkMPNJaMawVFEqBG8wi4dIYZpnI7hSfbkHFwItJuNJPYaOroO/d1SHTGD
QkxRJ7RrXSD446KXGchQfhbGVlK2KBy5euOiZo7q1SwQeqXtvstF9OlxHUpzZENsZYBeM9o0oIJM
RVYcmMy/z+89de1YoUtxFACgaO1wYmg6+XeQo1TZazdt43gW++Or8CI/ViaXO41xBCniz8tVuvL2
va9Yudul7DrIZxQssABqN83R4Y/kc5w0z8lQoL5bJFxRA6sZ+C0PHsCCPkwPl0/m771c6qcKAAVY
ZjJphKjNVgUuc6JrqUiPExXObtn4Av6epyZ05iXLbAGDivVrY+Ru02jp94WRbnxDBsLRTmJlRZ/4
r+mxVEb1NM56Qyj8dHDoQAH1db7wKMAEJ1zGPYQer+AWFyWIwhX1jco0kO8clvgqrFIBPr8arkH3
6SWSfIr2TjrEgBwWeWhGfVoW5R4XObyb4kzh2Wl8IJs0hfd6ifHzhBPvy9sV7q1/g6Co9zn2XpLy
TEnmByhgmoaZuOF3BrdHhAN5/Nzyumn/0ZOiWKeehJ/OPmm1focim0+zkh6T/x+UVT83kY7d6SDg
5f7iJoI8H96f8HQz0vxVtNmXGe8eytyvzd1yysZT9lk5Jz/5M4P4/WpDFaHXwqgetmsU0mhAsTgN
Fm0vIMTOsbfK9RjtNd03oxk8WTd3vPLEyRGzz+m8imQbPh6dLCUcTiRdsWwfKzE0+BKzhLg6npU2
dUGFrvF85tlrqXFENmCBk03sj1LRJjjgdYTVc2SNnZpszX4HNyBzPj9dB70hE2a5IBuWoe0GzAsS
Ndu7RCL31j9YQPPr7/HFRaxMk99rSr1JjxwYg4PZaNDiVGhz0/xHNdifug/VK6Z6jtMbC1YGG4Y4
loCUeqOton7Tk4eabCS3C8w7UBDzyR2J42/jtWkvFCTKcHDP4Cx9stKfAsQ1CXjd24SK/Ik3askb
/paDsQwjbwz0oeq9ZlRwAe0MyEWwRAwegeNeslnYsasz8ZDYIneufQZadyOivjv1qUpT+KKWWK2I
L7b+3pDc6q7GLMs99DrNEZ/AFfPYDp4H7g58/u3HZ+jlIYkiuHhIPs5m/SHETsP/5zlFjgkbtsqK
rOG6p/ExywwFUs+tK/YNQKXQ0098ih8pbBC184LnNjcevsTsgTWTF8BmbqAPoaFOYKWMSpug9tAI
fViH1OBsimKhH/pvvKXC8dj/3Suxo84ujzyQ66eVkn017yBC/7qIt7CeRFtoT6Or5nYLeZIiBWj3
afoaJdxGhOscOvvYiy7T6gIQ3ToasGmSDo+GDLTvcR9prootQwKFU0wClsP4JX3DaqXJfjNS+5xL
HiG3EOs83STvvcDA7VCcThM/PpIGsrw7oFa9oyKySVECbMXN6Bps8yppVgZYM/xHnplQ8RdOUu6Y
oWyNANwVCSKCnTOMaEWTKZwHF5x91rvFRioUx0sSGuJlTuCRdLfmul5p8koOTQErLNOeS9LLSGki
8fJn5bS2dSuzEGlgYaVyGl+RVfEW2xR9gIyX1gg1n17jtXOqzF1EjXbCxme4shZ7ceWzaa3r7mgp
GysNIuNmGa0JMhGBnYWortu9GRFtOaudxBzhBKdhLldPStq270odHRiSRAYGQ+lbeOSD4971Szm7
VwWnhT98sZzs9NL+vEO+qGXwpSZB/VKKCaOnAEJm/LFWlmFt4gU/LB2yLCK9x6M2pwQg+xUhIdaJ
SiPDQorBXwI/t/XNlZudbEv3oeoAxDl0bo3b1EnRhj86PBQcOZxTjCtMe/CwZpRE0QqW2UCYbKzy
1Xfn2daJII0183tIojdoj1+ILVxqjJqmiBsWbsAKxdL+QD6COsBxU0j89buDnZ4i323sv5U1yGqC
VSxouAAZySBeBqKJy3fghmBc08DVWBGuIW5T5c1a3AfoPUeK45FSKvaUNEqi2weMn9qojUwO62aX
dqLnKOQtV1WfQS4KtuaotWCBXDMcxr8i/zRHca/XVLw0hiynlcaPpF4OfAowOoK+7NMPYJ+skhOX
GMowq8qBpeum6DFEuqrZLSSWNIEmB1xD+k2kwWTaC7J7RVZI6c55xcam/fnstwPOR4zqOQ0RBw8r
g4VYNZ4opQT7U1ahvNbgqLsFtmRC3QG9MCWDw1ByFu/gh+EnILRNB6unP1AK2MNYXutX8NyvK1Rl
t9ACaT7xASJq86mf56yfHx79RBaisJGf9buT6CqV32BCoE9kEW6of0hKbYpcRO9/KnMUPDn3cfvB
6JYNLR6hJCsjLyZhIsGlYaSPZgvORW6oEAB6gDLjQq6BMtWjpVP23+1uoiQZMePFdNPvYOGoF2Mh
e9rZlD/uOrMl/cX6WCuUZkSMTRl61bWcxq7aWMgK8xkWJIWwy3JgKE0uKjdFaOgW+jFAr6G7NBGs
YQKCXBYwzCvMom66sNJl5J5FbwpymrVr8RTNCDzrNAKh2mHx8PV2A17dsVDwc+33eaqinHkJzahV
tFV2thI4WMEJk6la8OTgRYhXeqLetQrMRX1GMgXaLNYCF3wFG02JejUjzz0+l6AoQ5FbZISIkrB7
x7orsW4VhuQpbq4P/tw7jH2dcp6xC/1MpqrViSL/s/AZDV9rbPGwcKVTfqvqHfPcbSoljyyx82X5
/6EfgKAQjZfZtzfMQ9vB2458DJh1yWu6LYpOW7tHt0tIlJ5dFj2XHr7g1pon+EDdCdTy9pUni89j
LuQiU8rN5FPLh/UQsPIUM6IK1LzhcFi4Ixm7mAUAOxEN/eUQiW5YthIFWDNeqzC8Qg8bqLZs9mhX
Kz9WifAqClMho0mpS6AU+n73xuBRMBbWdvNVmkblkYBbsrpcMCgAP/pufqcA0xumPyvc/LU3ZEx5
Evzfb2Fv/ONnaX2GYdPFzsAY1wso1soqbXBET/29cNx5TT9fgSojUnXGqZFbN0K1idWZ/aBVxGij
EPwBxeeJSXnH5+osUkXvJ9ag5W9Zf7JFZVZRwkvN+7xIch/DQnyGEqI3UQ25r3PF4jB2ynaFm9hq
VrYPan1sa+pUsSAnPi8Q/Kz40W5z38YUIY2/70Ae5s0Z7tUIWKnboFg4uQzXA96xD8CF26o3MTMy
WlB5M24ajHppugI7+rkzfF3rEUypaoIzd1mdOfp56l+RLB0Tw5ma2MfC1SLE+iANEKFZtECuknrK
Iy/93BCY8yUpY0hpg/l+PADU7axpZBe6UF2PvwsSb8ouxomqWi9qIOOOpOuaOjGEzK1k4qaqkiBI
PTfVTycvjfnGcsdmHNwYvP/IEdsHlxi3Z+DnEvC1nFT1wXbmuq4hweTHJf7/EBGhFmeiUb/lEIpK
3+8DTbkXwrjHB+7wpSeUsyh+cJm3NnQJ109lBQUVn27Xsr9Mu5W7fNnsIf5v0VKUj24SIaqN+mao
nX52Ej/S+5Q+904Mvizm5wUnYi3hgEdgASp+iLiMFVktTKbGPwfj+FV5F62Rf2NCLVa4qEcVzAtt
UkmxkZuUjmYI8hBX6ZKHuyk7Ji2bIKd/uWDy/YUCowzr0lCvZVhQWiuHpTSUgn2ARWJk6oRSioSV
+DluZxTtrl+R8dU1+yq0u/HrAUhS6hNK6ntqj37+CiJTpjHxr5sP3hhhb5DhUtgrff2PPwShWGDw
w9SOzZofB3aR7JBDK1WvBb7vlpu+5Z5OWtQ69qTGcCF9WGjuVRYdriVGJ8bYbeGqBsWQVM/R7TeQ
2xwA/xSmsv/XuWNE3nYcZRwzHOjBw6O2U80ExN41xttG2MpS0rvcAEZ1S8zAGR3cnpXatB54f5eE
YfRK+ah40dofZCqECP8jWsFO/4qrqm7kqNmEWaNu/LwLp6VmqLUnShBJEjLkB3TCyHkNGmTM8rwh
JbKnmwPJ4bTTVtaFveAKwQaQfiC1/LX8bs0HlC0eXmBA8bat/b+zliIaD82H0Ai+AKJlOcOl+eqN
cIGj4cbfaZwB7hCG4nY/P/mAd+CfcrTPcftzhthySLSqAB5smTXSVcLh6qrnbVdd9LjnlcVisHly
h0hIv/7J4HGFz4+O/6oa2wA2/y3q39Dylk2Az+d1BHbrBbX4Yn0Mx233JupzkD+iX3XN+t/YBTcj
0LeG2yjfCcCK0s3phSsN9vpbIhrpj5KaSkdxeij1SEFQ3OujZ8kj9I7XFiDHtyOKUC7eHGkiJSO5
9oRfSZZB9HH1bWa1uDzZLFZ4ioXw804p87j7vDOlrxxg8iHimuDanj1HblZiUByKXQy9xD9RqPnx
FL2HFrCKHOeYDeSqQ1OTAeJEf5xWf0IdL/554bGkFYMCV7gKosVFHhWpPGRnxdtQbF76cdiTWg1W
xQH8U2mzsGueLZh3bkSEOfflJVTA1To01DGgPMw8kt9PLHq0hg64NL6bdyN+i0UNIkwdr9+PiKGB
XyqnzwfZRgCiUgzoCpV0zO5mjwUFlffys2lbJbPQxX2wnVrIpd7kn+ysZ2KQPvB1RKq9vuQT6G8P
NTONG5an7CmIgejxbQRfiakwWYhJT8X42gIJJaunEjy2wpDVf6B/9ZafkoUX9AGmr/K5PCodqcBk
PnTnFLqmeMGpzBzDca9eZwk2DzHSNLEGay7FB4xw9DTQoCwkfgRT45j8gDBsh7c3Iqbz85B5bOoR
5zuHQzrQ7PSePjaz0UjN2IpGqFiFc9eW0HobBBi8/vyzLiuNR4Bz/rQdDfI9SBCpuCFgBUwnkQ4o
7Z23dUTb3J5QhJxT0ex1i3zezttMlLScDCYUaYq7WlSgkIGlX/aJ0+monBBs+Vy1eLB0QXImXij8
NU1t42xW50gz2FfnXNZcl4Bvl5F8Se4WPReb7Osw72QEDoo1qqsBcmuOmOTjUEplc/69NYsZAehz
EXFcxmAx4SCnv88K5l/QxVe5tjwLpkWeeWUpRBk4IgYc6M9CIbMNB2MZVBzb84DdMrEteG6PrkjU
u7+FyjY1dpbDTWhHhbvh/F5suMls/WJbU8XhUTCqEyLY8s1rNaoAvNgwEflh6mnsvJtX3TWQn7lH
c1ORXp7wdDThFOSDZ37/cG4y1eui4np1HJiOg2xmKZZhJzEQl5GSTSWi1quFv7n4gWdRur4vhKNS
VX/Lu2SRxNvY7OF9axo9m4OOCQF8x/9X6H0YuFE0MiiC6Z2g5X9R8d3RDkczqkTkopnHcKJwBOHa
BlfZIseHWS21u7P+Ivq5GaTHb8TS1plazK3yC8AOs6mtrgysFt1PAeufuwawdR9oQ4Wutk3I3HmW
DtvraOx2LA9fDH9DBkKyrKW3YYxIQ0wW2o64wdWHuVcbwLkXDvtLyqAVY3Fy0txF0HHPyYC4inbc
N5KPlO13UtbC4YApog08G1iZGoYporF25TYMe0l8YlOaWTsinEuYYG/qVNweaWIt/OOfhjfYbT3M
7BC986TtTE+a46Bi1Hwgmi+ZdwXR5KOLtfSoL/XnDmanaBZ3AO9DdR9SmPWovZXiqoBjFpc1ZaZb
TxCFI/RObKx4vzOurG7DUXVd/6U/ZB71OzkTaJqztsE1h1QYHVLntQ2Fv28p5HGVinhzwDJh0t6M
fJANCb1XB/YDKejvG7G8bHVjaV3EHb6iynrBzpau3kZbzX0WmBr+Fbg0MwmyfciXEQx7C4hIOPcU
Tqt+nZjhDG2OapZaxzSyuZznOXb6NqlbJiV+a+dN5Ut+loOb1vP8akhhTLoF9aEo79vsu4/p4BjB
CT2QrC8/4awxxg9MHksZhnRNJG1wpxjDWIYU6uPmP6AeCncCDyjXckAc5aSZA+a4a73NyxKE9vY+
x/CPv2sXzzb4fAtL3d/gKuqO1ZDYMAMPatWDNPc/3TjMDoKs8clSGEGmpb7jjVJbyYGUJne5+cyH
gdQz5Rm2WCGg8kqp7A4FJX8sdvhaLmXmm5T7DhOfT7sAaxb702FWTGFlNumxJ/3ydlaRX5wuwvpe
9PZyInLyMecako5Z2bPR3JMdV7UfgJoAZu+iOyIj7rxjwpwJ/4MUvyxY5A4fFfl1vh7PtQ0tltyg
9/hV1EBQAfOcPLnZAz7/hmyDM7ep0A80HXDe1WdM7FA575tUt+RtfyUJ19mK4NJwCi1Ooq2z+aw1
cblgwJIWMkuS7xAA2/00Ml3L4obsL6vl1ZxCbwxkPN06ogVgg48PljuXwdVO1qJX7c2pcx/hds3a
DC0qih/9Ak7N2q6L/Ay/GiKb4fYhlcQTc6wz6KZdiSMCSF9ZPqZgwhvqkn4HzRY7eJzTT3/R4d5m
DrPw2raHvZeUbyhRCbRTrIvnIlS2WY0kg2okEiBC9MeBBwciyjE+w2ia83jP88wj36PlHMsPhq8I
3Cp3chMo0K3VGhEM4qebjA3ixrHXHgZvyJgSCpu8A5usuIwe1yhSeag3rtIij9hagIkXcH/KLwsZ
6HSbEfYzPGlVhrrXcKc2uPHtEw52iZra2jBUIn7fzxZFYIyJ31hMzXZ8OFEg9oIh/T6eB5pXNJ4C
353TnL7M67aZS63AwJ0s8uyrkhg3tHhxz9OM3p4A154174pT9MxlqRF0gT+IIolvSa0IZSDih6pB
Fmnne5+BdRI1Ksva35NR2gWhXF/xUbBBC659vaoWuWoIghp5qRqAL5+V2svRLTka9nSb6KlOhui6
9Y7OVCGStIKKBl5g810yPH/OgANKCKfyIF70nBWceooItgaI444W8iPbo8fpaQMSCyfpY4Hy0h9k
HaV+O9Y3tvLATpk+R5nk1YhhQTxMVd96uyGMCJcprD9LUKQSr8YiThqOgS/R8cZLCuYS/oz7WZi2
M73k7JGnBXG4SOUgRDs6vc+1NPOwwtU66zDXgHCOrqj0KdNnna4PQkDoK2NfbOtSiO+0WsIMN2SY
ll43C4TJ7ih/Xr7c78YeIHCzcD0g3yWzH2qZyQnrtzFf4CqxH1WLtw4gOQeUDggoz02k2b7aY1EG
UD2trh9kXGj4DWP929efN4Lwf8vYIu5hGf0iy+mIhdZxwF7mDe9KMNqck5bShUH585PvezxS4Pgk
2sexh75JphQGVIfQT3famn01AftN3P4chIhh7tM0yCn4AcpSg8z2Mrb86BTE5sszQf777VahAsDb
D4bPxDBTe7KHdLVeS1li/13WUuvVCIKqzzlMW4xrHPScZo5CFNnVQJXCzPjB9Vbxk9LrxLURDXsP
9AKGDQtkUmDLuY6urX2Nko3EsAcpSq66Tph/od4BoNIqdcM0KBWdb9hdQQD23HaINW29aK1RDeIJ
6jsc57XiG7wqkbpERutDkRxMZvXVIZgNR5toiwcvBlliCnAsJzuwcm9OGydvQCAnLSs1Wngf0smQ
ejVZKb0kyIoZWYoKjrPVWeR4+RJHx6nPbTO/YddKjI6ymGmUKEPtQ7ggEU5w0Rdx2Gr+PIRQlXlt
ElsEWu9NkkRwvGKvQR4RB/D7diwAczKX9kYHZO0kPtp0GxMYDTcMUFiWYBbsCLYWFzu82MFOeyIf
YywBR/nqMtlnPE7ssJWEtuL4lmowPE0R0l4NT25lyfKdds7v8CdRGBdES5Lw1SDJ5ijMZfcTH5/u
GUrVi6NBwIvdcttbBnA7F19VrHkEuZFhmbUM72EHOTdLOMfC+AZZU0sZBH8gVQ8BzQ5GeWX40k26
QmDJS8lEhlUuIS0DLK+MvhSucm0+qYkuOPHyU4ETKI2sb/2z4/M1/qMBZG758KfFp6MUyw5Vn4no
TBvWJFcVMNp6cVURipC9JnX6vGdFYoIZi4gSvrfVEOK6ZaAdCNkT74Y8a8Hj3ZlZiuDExn/UrrVK
yPUPbzGXHJoutoUBelYrTiM5ntf5s4Ugozy3fqA8t9KNvqkxh4QXKCjdFOPfluUf9d4nHa7smyux
ozZcI3/cHKEK1vaMm0x0iSzImsgK/YffP2lAuNBeTVifHmjebQw3x9oN6Olu4lmVmk4rTs1bQK1l
o4aneiwU9qGtBoTbVzzi5ihCYEBS7Md6ic7ol0VjGJyiF8CjOWl1Br8qjTb/Wpv8pOOzEn2b6LZP
RJJbS+smmbGdndU8s5UQ2VPTU/7YpMU/AnoKC7PvG/cQtchhuOXSK6nONb4b/BLtnWt/fE9RKaOb
gG496XhmMRVSdTbc8roLwDMw1gfTOHdd/oWVNi9NYZ7g+N3aZZl8bXSJt35H0XXOjuSx0ZSCKDhG
B3CcjJZt6tduLH+S7Sn+np3ddAXZYW85M6DR+ggX0XMR2oHPruQ5evLQyIzMkUaNLG1Qj5raDfZc
56XObhIgO9J/2zDg0VkH8MkJF7oVgMr/zRh9vHIueRq9SF1IlwAC1rxEtAbZ9QJmSQGNrULrRxBx
jAkNd2f6Yivfq4Jy4hsxsWUKC7zNIaX8/lUI2gv1ta+bpQLKU1G75zuRcp/fVcF9wKeAud2G2Alm
htVTD4GxRBBMzuue1CLbp6Bs4lR1kCYkNFarXlDQTNLTuHOhbN978gh7eWzRbZhikJIk0S3y7VL3
Oo/fNfldvct+L+5hNa3WzM9PzwihCe42lukEV+Om6gsqk8TKte8MmHbnnjFYvWRX+wECZCSA/e8z
9ATFkJdzsjnmiHjD+ExC+Igq3NijO+AlnKduWXyNzOdLi8r8EP2zn/FaSoU6h3N9f/2SR3ie41En
MHHfyaq1rVm95c5tadKxHQtmjPNTlDuCH8QoCXv2ZGtttZ3LoSJqM4m4w/C+2jL6BGdM2P8RJNlG
rAsXQpl6YwA/x+fOLfgAYpa1nAix30DWWVW+DzoalRshxd/tHlvqSfTZpQwfggRL0Q1v0pHBFb3I
Ak2RQHkwaxuH/GU1PJlPfvYV54ZoZz+w6VwTXYYdm/jeEsHBLsf4N+LFY0FNleIZNoiksoaLABnk
1q2iYl2l9UmxmMRkgKLUm7ZuO5miL5ExK6dooexnaA+1gkogYMnSMWVnPk/YWh2ZHxlOlaErUwWQ
PaPrJszOX5lAVR7pNMKifkLj3EwOvv5bulUhPgJGW04qs02bj4RxN2O7xRwJwVqJeXOb2nFO4t6e
6OQgz8xIdvl5UI+P44ciS7QZmBMP9SeHGzahKShaiOqDRpycnLCkgjq+u1KOPYH4oeOjCNV4ZMLl
bTOvEpMJr9rF6yMRKCwzFIMIPo2vOJALOQWvpyu+ug/CEmQH5f3ikKfKY9r5nzVWYVbo1bM7q1IL
URHOgAHPJ2cZ3wXN/v3ydTyhF//BfUIiU6vFqvQBy4mu0oHgU+B81qR0FlV8lIoKStEbFBqrGOca
q5+U/NZjm/sjdpY4mhVSmnfYOQpYC0+FAQoyZdHYtus2sKw5s9MmdcrRQClb32D8KQTcW1tRA9aM
NNQ4YcboSCH7DMhQdcur/COfjazTxJ+UIM3igi4F3/lOtxSsNA4jC79DZxm0Olalv8xNt+yZGJv+
0ER+Obi3B8mNnBiFCjLcqG8JgULyNdEZcI1NLKJ8Opeq/UsP0JxkBtEEyr+Z0ocgX9kbtAwe2w4g
zLCbIhyqfesVBUNpV/8VeBn5uArenowh2Gg3AyPOprtUflZ1ksbUZgnQM2pOyl+Dw7hwHKEts+Co
+6n9WoyeSZzdAYF9BjdV0oX2KIKxqY58s4mvSPjfIvZowQlf0r2WeLFoM5VQDUH6m0kV/APJGFeK
/cWyWWPG+rOMWW/N7Da+wWkj6W0shu4wSj2eSi4fkHPIDcIMZjzAdlbudGKtJRa/VY/rORK+UImI
RkEfWS6ZL+h7OMsHm+dMGU/5nCc5g38TtYUCr2Q+TdVap/1Xcayf5fbWZND2WYBJlX2/ojBdNMj1
yyLrXz36UcLek/h+d4kxufXEDX+febj2RUFfaf0zKkgHwGDEgDSxvhtXi1IwQAbDgaIrulz5vvVU
c2ISS352ILlXWc5/pn2DbaXhP1KTOmm+H4tBKBW9noYI2jaWtGJIiPIt5ie7FvyNpULaPNONLwOX
SNUQhjYaKpRgwVQWx2xaaqRM6a0YtmVbN9rLHmoDiFFF8Io3imiCIYAp/MubVzTw8UumNvyjSbJg
AKIz+HsNut3T7E2+7gtW8xL2Qu2VZMPA/adWS0L3zyVD7UGDFLcXvj3OKwvqd1qglw4oslOPKvHJ
zfhHUdXTnD4d7zxzdk/3pDa7mCzPE8EUwtYR9UBFGcteaVMErXTk4n8ZHdpqJZS+bTpEw8M6LzmA
9lqxfNEiTvlH9sOzGJamAtyQatyeEGjpLDexZF6N67aZacH4z1YU+RRRvubI2Z2x6ZvMH1gNZBMk
hCkCOn3qb+iGp+Npt3aY6z+LNbDUlTGIX1QFeI4tvmxnxNOqcu/94C5C935eiI4ofNrwwKYe9Z4m
CMl/C4IeRZWDMav3mA/CNa60cM8gYRvV3Dp4HFJtr0DzuOpq8WJVzD8gtJnxqHNtBPo7/+gTQoYW
XrUnUuLXlSjo4jMiqMdDZysb1DNYlUnnvTldgFZaw0LA3uys+fRYvy9JvF8FfVqf2wzCOvkEF1GC
IxQZ9hD2N7hWbjaIIEFrlXqRpcZ17/2i9Tjhja/8w3zq4ttowj/6EcvsHrWDo/MFITDfJ6Dy50ZU
egaVZVeDd3iL5EJ+OfzfZIC9+g0HugzMZWKNIO0PHAtXZeYb70sc0hfB4ciPsGxF3m2SDbVkQ3an
eex7frjuoicJv9KVhkVxvHhI86KH6u+mu4cswKzbRsVKWYP8f4TVnrcGPUR9WEJzQN9fAB4NFQFX
5kUgc1lQ5XEQQ4afOC/AIXbfQlv5WX2caZbatXf5SkPEmPj5aqhxawyeZ9y9s9F2oJRlLBuFtxcI
pdSFCTRsm5gh8swILIOMw8XBhAD/5KrO4wjJn8rPrI4sGXndqozASBuRB8cs8DdpuMrIg36y2xI7
FUdkbgQnZHz0wta+ehuE2TymlBrdF8v5VOCXqk5kgdWlE/tGenp22UkU1casIPKa0kIbd1O4+Y2V
AgLFWCWZo/gpoF0+R5gaCBIIExhcnUYYvHL99v5qftEF3ig3hV94vvJQhNdcqqNF/iiLl0oUI5v8
v+ee3PbCOCGctlxBPwKDjqc8V9aM50shxEDhH+Eox7hWa5x6RW8zH3VZmEEvuimVmxlRSw/LMHXn
NwAwVagVAFahZOghyVhYZUdb1fcBVoaaSJceg8BDcubZOacUcZDk4olS/iqPUItFwWhZYSzdcj7N
hiAi8EaSaIFakZA+ENGZOJn82rBL61lJz6AM9vgfXQ4NTcLmGRwgrVuOlQsyOe4/D+jdVlhKCZOs
jM6qiBoQSdrW2aSTGwHJNh6c9fMOe1J8vIABB0vPp1iGVyZDf1d6CJqVMCYTy/xgjZ9Q9cCQq+6M
m/xmAVtnZqDjeH97l+5LW/T9rBQNCURI6caw0OSrIpxTGC0nMwvRe6wXYkYgamUvA1mYyq2p83zD
AhKsKQnZMrRJjQJ8+UqN+CD7lWuF4ikh/BEvrMrfL2U/QlbVwbKqDJYbwor3fw+eR0ZcKJHg4ING
plM1FIOhyJMR8Tv2c09dIwJ9V/mwKg8/4tz6CSax/SCtkjzs2zoUy3GbYbsg6VmeewtfB0k+sPcj
vVUwuxZhEw5nzVKQFTeBnvXMtcSLkiwBg6d94ZJ4RAe/FtQSoBndYJt/2ZjM2uwX+UZ3hq14UrJp
UeeXpqZD9YCx92A3NgYKJTmoVjYl8BLJJaUDJWPmogBs5lzMrRPUZ98my2rCiizZzrunz6M10wHz
yXsXI6/cHCgml/a1EqKmC0qW5sYxcbBqXeergOO2rbNAclNwOE2tsU12+iM9Hlk0h3UF/2Ai7Nzx
/vAKmMC96skSp4eHA3WyeQQZIIczjp9Vl2Yg3eZu6ugaCVnPESFTAror+so1K+Cfs1acT3hQqhfj
tc/6iqDg/hozpGpt1zFgUyd0GO+RFhu7H0hbOQxAb8ImDVFET/lkf0KZrP3LZyHRdGbLcgpgeJ/P
etSRuFjSO96NDcZZi1mvvUqd6R12yXqW8Z/qDaMFzDuTrXNGmWgNTvcIYu2/TjnbM7fmHhiegN8V
+LB/H7NQdU88PiXFTT7IBeqaPkqhQb0ZiLuAfGeQyBn6SzcKa0j0NBW2NyKIq2ED468yvzzBt2sL
az7SpYK0XTlXNvOHHUrIeZX3vd83wZ/zqxZCAk7hZ6mQeNQ6NYz4VUdNUvSx7UAs1/pUFu5yj07p
Ux2YT4GfJaRDz3ufc7flPYJ2BTZTpGCcqyVKlcINX0QJlpkPc9budrBXOjJg2E2zCnqQ5SdtgveV
DNbW45ouOy8+To1sj3qkrZ1OlWGZhPP8jvVFmh/P7wgt/TlHzFxsTVW3Cg/G0ZBu91K5h/pwEUlD
/R0Gnwh3MI6zTW0CwXKiODzIa9jgeREbqmjmR3K9jckAS30QKZdHXbjdpkj922Q9QzE1+Hy7lIT8
rqPnEw+bYwPQYw3cAoEhapuHyhxq+o/bkMG4ijcSYFiwG7Ymfl6d4P/yFpNXeLaQjFd1miUrovWT
8OVRcMIRB6HR4iLQknDKx6dWFqjEEqbO8NrTIvRrXcZp6m251GZzI4eIKdd2BLPq9jFGkIo6/Qsj
qetfrb0tn5FS+mvwaBSE4EcXyyFHgdpyEA06AZozzVYAvLoBf9NVwimshKz+LSg8f7uPhUnIrD/K
R6n5TDpTyQPRIh4HojOSulJYGCO0r3AOxcBKM4Czq+T7J/GVLFkNQjG1130BKJv6xnWNydsys5CI
f2gyIOtFGwcQRaGJpMHa4GK6SFqSk7BuSmiLMHRbzqdoqsPqUU27Mt3Vano/KiN2FD0HFvKDunK7
xgzVPkdYRL908wghUhBCNk7BFjJfGduMlM6UnpVHdFnhcPu10/BOVtdTSwSq3VCjlpIUZ+bxfor1
EVjTZSj3x17aid0rQLBI/aCHkCuVzjKKI+tDD+UWtDamYS1Jyxx1PNB4d2vp/PSs9ds8cqnqZPDp
yZzpofyxySdHkKXmzXUbC9SFerLK5/u4OLw+rEDQjkDWaNIhMskWNW86Ee97eKJrb5ezMGutbe8f
cxkZbDE8XVyZaXkeQmeV2ZDEcndC1b9liWJPB97wJgZSNnZ4GXpVT6j7+nu+D/AIf2cCFgA4q/2/
8ChfkSKRgAx88wOMs/joQVMaY1KsFvkQpDfCOQR5KqPCv4iJmv3q/BjFdCwso7vj/cOhL2nu5Ypq
8Y208WWbFAzH40zD+UAArQHhQ0Cmwj55e7IOHTwEqdd+kOg1ysM9T6TzGoTlNDZ/cvYI9uLmH08o
x7Ip0/7mKsAo1jyCsV3MLAMprtOS6h1Jc5eMhdbiSQGFeagcjxJUJQstmAsYkMVl/RrN0ZD7M9yu
3mLOtqlnnL9m7pvkCO9mco8F1wTtPjinl95GjYY99fkuxkXDOP9fjk5TkFyJnqOqoUIxCad7BwNm
28iJon5huC6W48zlWnmRLXAU/NFiD8r3MoMZpa5+IjLDNnxP+PVHeVRkJG9C8Is/7dRqVTo/fW3J
0dqEfsj7IDf/JQpMvavJES5BrBPoMve4RaYIHNparWpfGItkaUmmpyMh3yoweJdIkcpqhlge1e/W
iVfaSaWlgWiB+EU5elK3HLPsw8RR58jOXz//6+/29ZMWMzI+J2DmEyN4qotc5qkBliFSkL7P0kAc
DAAexS6iZ/fwSaj9/JnBb2jD/snuicqc5OTBLA9y9nPzF6V5vjS2pnWOkcXL/g8wbISU8rnPnvQV
b1dKLlsp3U8YQRU/AlOgbJywXMDvUCoTZlT1nS46o6LoxaDTb2oqCdxWmEyElYJiTLKnTvIFYvn4
Dlzkgtc9Zdvhy+1osA/58T7Lgh7E4gCMS/j/NiQC0gYYYuaz4KVcR5zNjtQHJ9mbYfhomwaRgkXh
CKvAb7x8igCp3dw1no9EYFmzEiy8NtUIAgXPrcZDghwo+FmjdKc/K7AnRY46Uf23vh9WBwELAlqV
uo//fkFYFDNmOXYNlAOOzJS1WYlqecC5wRQvjRce2ObgD2cEypR52tLGXcqpKTYyyoiAq4V7kxJN
qOIhBHE1oflykWLWTvEfes36LtwjCThs+8KP2tp/DJ9AHjGtDHFV4Xj1axVB7OOrA6Hkd7LJtIF0
evqE9ZyWYZs3wD62HskwXysAsMaDQWt9dfv8+p2rt6yGYQ03qBihCcdTWDmycesBS0qrCV0Z96mC
FkFBxlKIbtHx5V9I8deHBvZSZj7GQTOfPAfeO3hWZZwmxXBqeDhW31LFELt222Ia+ZNx1aJHz+Td
CvgklZcEhi6ubgDhgVdbP3Uw2sI89J+ylzbVQMIzmgj4jpGbDvTJyX7RmP0UgOZcgMpPahWrdb2u
bkDI+yb2JnK+c3fyHhio84OH9hKoIBZ5XsufjsVhmMzsGK8amXpjoa5V7bEYQB4Ug8ph+XtdiNWk
pFDo0B+1roEgZUqI0lHpfLSH+s5FyikYg0Ul7MIbQtG3h2DA54yaj1GIHppv69DbftzMQli0gEC2
rA/R9lFXuALA+7tfhnFhe7WLEAlw2Q7IPeMZOrQUlcvzMa21U8Ix3vaGc2enmYtaPsEhABT0ExmG
VwG4ZOlvJnO5qI8BZtW/5MiXNms2gKaU/tB24tjK+wxyOABYosugcpNLI1BareaKfzX/aa1zFZaA
/mG7zVvx5qNUFflLmqN3Q+IPll61ajw8xCxquIVAy3u2fESGq3MaIEqyJyf5PgfA4d+8l4p018iN
+E5ucRzFSk9ThPXcFl1et8+Yg5Tc3PjYp9IHb5Zm6hs4HvWEpxGtgUjQk7+EgQXux8lNOxmPP6+M
abdN8x3AVWW+zNDkCebwN9e7/ooKPlBf+QTlTVzbaKj4U0LAiwEav6As9sWOv3PHEBv3dE6S1E0T
z6onSkmG3aQpsvbOXBB4aJZddYATMzBSc00sBGpxv+Ih0x37zSPraF3kdir9d7bcqc3pL1OS3oTv
6sd2yfriB7zuBQqNlia1dHCigJSS/uXJMKKY3+IhNXacQil1hdwCf3GSf+v+67PT08rHmpcfwtA4
5frgwk1X8POnFjpCiNW5S0vaRrrVxir5X9mscgeNjzjHBZxQXUdhN4cfmTIo+GKn6pqTKolvj1Y/
rtLp8zh32PylB2FhvVaFPmg79bLq/WUdEdlLDOo0AC4cYkYMuZcuB4e6WFXoPVX4CJY+sK6lNhIY
7HlE8DoTmkMASSQfXAwXt4OYk4/bRFv6jtQpE6KTarPCz00yLvTvvxQV1Rl4ovpA9mwHvbpMv2Ip
RQn3wWJXQEBy2u0nrGntbWtfltQPLSQ6MksyitRYeJVqY01G/I4prh3LE87+bZHvTJEVwQN9oLiP
Reb1ntG0Wu6H7VRxE9YJWgt56pQtkoSIWi3Ye5yHrvSOZj3cQFLmoiGqfQshgcyuvMYNgSw9t11/
1sffdJw3oyNGMpLX0EvEK+nsjQZQ2aztgbxotm7v6UkpKonbnlnJA/8AV3VPSkP7c15f9TTgMk9/
qLBuoQn5beXRg9VneAxhVd7PUSi50qp5RBgL+oar+Un56Bl4fzoxtCA+714ZNto7jPkyXw7wVr6r
sJCbDYez2MLcws5gJLbA2+bEqwKmyVa1HlTIo/x5hDGkvq7pXoGjUONvEyqubIc/oMfq/05P1MAf
gAs6xQ8n3JPbkevg/fwh+sKvXQIRdMJdaALDVsVjZ4Up7e8wLxc0N99jEY/2/KxsMiXosGRxAkfc
NJqibgYpGHXdlM++mlcumDgnP/Ircp/o/CdH64oG5dyHGSngJ4lIcprOPqxq38vZgBkDLVQ/nUaO
WDUerNBO2G5f63hXZ7DZGT/5nE/X/W/ZiZII+MpXcS4zHt+3aKpFzw3I3YwGNmfYe4KpmQ4kIcSp
+F170AUtHvWYMCTIVqsSgDtVV2zff2UQYBP+4lnVFUYjreGgJZdq0+ebAVhlG7m2vyUnaaemkK8L
gyTY0GPkACmGjxPmsLkhf+dqDVMs7bZfAvxx5UDPLhT4/+Xoh9A/ss4uPsxAFFZl958ASXr2SW6O
rcOWRBl2X5o79PyYzKtESyC6pPeytKaxhqVSV1lRzlb86AbYEBxLlaHZTXKb2Nrj6r4SwMTXI8GR
tZhXkEXcfBqPsaKsxRwQSIuMr2L8uXEGQDcjwlbn5JZ8AqjbY6T1JQy4YpEWydszZrICrP2NtEw6
fBXTBzdhQMS5e6tDY9WkMDYWs27gXqofY4vTpjjFhkEcjFBZ8MTt7oATJ40lK9tcLajW5c2OtyBj
AjHQcTtIMedG9X+gyasAK2uAYtJM5OcJjRhx5bQCmcB+ix0lr+NspTwM/qt2wOcJFTwS2TKdUBpc
+yOMfRT/HV2GFRR2bMc4iiw2VcJB2HorDWMXQu8psh/Oktb2yD8UchSHIi4yX4kZAytkgGv3iRwi
7yYyXbAP7101M705y4CkgMBgYB4zFob7G+YItiNBRjjgdDNIHYYFRLh060ijN1gGoJL6ZW9kKWgM
yYmpvdQMJycbZvFJG8Zrw/I/kW5NoWup+HZOHxsLIT/PRx7j/8FtG1lPJ6eGkmqDDAT2wN1RReO4
Y4C+OdBUvgpmYCyInSpTRU4L3rQg7ab+lU+F5LtnSZmd9BwbaB7GMG4nHv1jlTWv9aXGWE52lD13
dasX4PpTKMfqK0siE9Kkz3cuM3AMMirrrlKi5UeePi1SzovR1oBEhMKpe2DFzU1O6XvmqcL0kCPt
KTXye7B2+2qLEeABUHkzQNMCKg2gEgsh0xicgdr8ssVG2Fc0obaB0Xus+j7DxkWTduqlTPtpGm67
5p499ir7XBexfAkdjyFr9upXeDk1jbe7ICQPmvxEpcIio8CnFm+sNKYPoyc333kaAuLjhnOQLxMe
/MMylULZyqugLRcfVkXyOYVHx9v6IPEzG4J8m2T1psqtFEk/39xxaYPfpGv5QezuqHvxuIvVYCaX
SMmqBTqzrdybJvcMLNue6lC1XBXwFmxGl7ULs4MhByuXJCO4CADlkLxiXMnrM9G20q2hkrj0afGB
yBkG1HxzSrh2JeETkbD7usFdw5CW3uzaNPxVccRfSvGlKqf7/SbHYXwURaUo04IjBkh7YTxTMARW
pet8tPg9ybE+7GjE3gps2+rRU7FZJund4Y3GNomcui0enimmaWr8DiKZ7s/CGXaXR274NrlA6OgN
coS8AUcEl34wAWLWs1so45wKSgFMtiOTn2Nxdlea3Yx522MmfPfTtpx35Bwo4aAj2IJHygst0eZu
p2uw8Y2gpC/T3oNX8LI9RLCibQIm9uChOtYe8ptr6Xn85z6hE6C5dP+hURU3CrohT6BEvD6IoHMr
SdS6bQjHmX5b5II5VsgjSrYFv+m4uS9vdcLj/GJGffScCOv5KDLwWD2OVEkbPjohOuwOVYoPy8rn
C9KQ8/sRBc5SO9qbWYW4CgqxK7XjEs6r2xkroZo+8FKa1m/Ohke3SeCBNB3QaQa58vg8Wx6zEbME
4DD9tgPtbmSQ30Rn3rATCFCBDKooj6IsSH+UVhH7OIhJKHgYjERxTXGCQhOk4RBWnNSXHk8NPXcC
wO3PlTOlPIbgXI4m+4jDGHVE7jQvWCN0Qz2XULVldc4qkO7diE3IQWOcMVlyg7n/km7uT8sCRdxq
KaFAZ2qRWrEExrC1RDzmtZkx9ol+g7u0EkNPilrI+oJ3mhlijc2LtDuYdJJKGAEh1PeHjAlpIJe9
nxpa6BGiIDDMAT/ahy0k6A1ZvKkbjnjNiziKywJ7nz2qEfBx9RCcIt727AWe1odRGm4MsiDO0mSl
lQd+wQxox/o8UQ6V9LHXAKLUgg8wvOjq/bvc+9WzLvZLkCwWnYOmfawKrFBmxQJSqyWymrEw2B72
aUbx6kU/QyceMwEs4fKm+8DieELSJHPzb3T9GsSNuljADP5hMt8PDR+1vJmY9RxgDRIyBaH02RFR
Mfxhwlgk6NpF6rX8W5nUr/dRUhgsVAote3o6Jk4x6lB5JQn8Y7BWmTyGtp6C7HRHqlkW6tPgibbn
ByO07QjkF1y/C8qa+RAXZfiWcj5baFh6EB0ECsikNUZCoYAIJhbe7eCKzqQqD3NSM631JY9wpo5t
UstmJLTrg5S7z0uw0M5yJqnNDqatILrQgPS9b3W7ihyPnz6cO2VrloMw55BhW5LifvgF/c5hRihC
uP18l+f3z6HLwQPOtVM911WsudR1y1l8pA7TtXBZeEVIAX2L/IVTjuCSThQroAtcLO8h6qMfCzC3
bdJXSNEtXFrX7MIxVJL+8dJACg1iHYFsAsIHYMt0siqthtU8/W1kliwQHFB7bvT34DvlEwKzjB8Z
6qhu75NLc7+Kc4meU+VwK4/anuVf+CjG/V7PY2GzhrAYptcItdfUUu564udqSmjE4GVwEa3El/Cx
nkjk4JSoFrW0m+WFcWeJU0XAezpH8vXZtxMI4+DXxOfJ145X4jkkDTMT2TyucLIM0Dt7qE+X9ku1
TkNxnN9Sa1/XFCDCEBGHD3gG6/U9o2oTfuZtPY/dfaF7S77p20P7y4gpfvqwe91hNxcdpYeuCD4/
1NkPscZcfrMHYS3wVhL33R0z+ljt9lqF1NtBbVBgv49wG/U1lnKTmOWEj9ThxHUPPbvHycfsY9hE
E+hJgajVT14aLGAbzUw/BfqERpDLgrOMwGuSEB3tYXr8/Vx/ECL2/39jKqhWNkfGJjr+hFxtly95
05A1sT27xI6WBX0DAINiXztPJu0Hmo2KDQWEnF19T9PVkEK3nJS4G0z5BUpNa5wxlfLHAVUc1E9I
GixSCBN0wx1ycgtet7JuaFOW5z4ESFFXNRvA+OcymxMfzACFRfkmqOZ3F0wZBPyXzYew6si8r/O/
txeQb4Wf2s9KZUrJ533gQtTcoLh9NibB1QXyQkDgkAP0GorgTPQhKOTxfEAHXcLbK+eXLsbLNoVK
22EFBNktg5bYDUXTUduTdyYG2pkCg86+RfOWchBESmuiIB3fGCPvbN7HkF6bKC2qoTx5NCxTkKD7
l/o6BLqTwawpBNIJPG4HXIo5JmfphXiZyOsKDF3AgfHqTXeTD86sv4sA1V8b/ETKrS7Jlc1HHxik
ci4sBScs/6b/g20KOGLB54N5ZEoKCfjw3cNAV7QY2hzq+klCeUxrmE8R93Xet0hxrcDrulxjqV4V
ZDSOfBMTJEHPKapkaUm4ElFXtcgHHntpM2PrSxDefYCzKz689e84U4VqZbrhAFdpzwM92ArAv04f
vjNTeu9lDz4tWF5Rd9kQAR5xscRfijycXikQPGlbRBx9JDiJldD5UoUQLCKzQ6nb8jQV0xPYnyXk
Y5+fJkkiKCvr+UxevpQ+S1RpHe+6i6E5sTWsthMOb15aVprvR5h/IJvvZCU/GHc6IN2miECT2Tjm
baajlz2zml7ZB8YxGwYr3w1sleJSKRXnxGi5bLRAF4j1Gyl9GiOpm6Natbj5tqUt9Van/KGXA7S+
6ZBinujpAvCoAVE/kOC20PNDSwM0XyhwAJKOxaWWdijOo06Eb4/vKIYl0TGWKkcaFRUq/p/nJ5pD
7z2rwXXHfkyV+jYkbvZi+IN+FLX+j0yGU03lt6xniY/lAu1EzTaHDCOvz/XcVKTLKshhLap+IsSF
TX7ctcFq/HprdVgwTviCdo6L8J6O2zaPv3NpjVc/yDcEoQYYEiKV7bNWY168T/Eu0gNcDNtD/CV3
BBqookkmHS8634unoqfE2qaFTSZTkN7vA/VOeoYCxZtXnWnH1+50YYT6GtL5c2By84Ds4OZKhLpk
CuLdLejQ5ymRTP1eVKc464/unT211aEdiVeQ1FXWgT2/0sO0Om5K2b/kOTzR2GWtEL2k7AioYckn
cngMLAGkr4cXTO965siGUgV33cM56/skCF+rfe00Dg2sAKoCJlNqYfIIw/LHG4NK/4uKXVQgkSdr
MO3FwKYJPvIH0wI1BU2oS4rohzmwr2gGvynCOVpn6xChLTTXDCMXUs8XUnW88F14qK6dlIYcTVO2
JiP2YOZxhpMy/HONrxaV/pDiSswTUOrxZFQfRTX6lFsu8c/HpcZmQwF0gdmNctVvSoyLMhTO1Uho
obUC2hHHcMdzuKtxpqfPFPyuyrwadeGeYme22rtOKNb6PP7g0UN0cc6gIo3gvHTkUfF8GnVMoNeJ
Am5cn2XfHeOwAE8+NUTpz8tLuzsDW/jW/fN5skACYhuoWvmgG7MVFcODd8Ji7T234rDbzhEuAOjP
LGZIyB4fm9FAOCGyrU6g8gDwZdWh2CziNWlZUbS6neV6VxVs4TCp8k0pZK9WTkI4GRRfoGBl4wks
HjtDyvGtYBf23RgVCiPqK5jU0xJr6ypKDDTE7XeOExdjfCKsAecjZYqLlEvPx/mcctNp37SzYDSv
Usrfi5nz95liatVa/AbXp2hG0DWmrSfMOEDeUeYQYW2BqreGdro8J9YoZBM8GVcYjS/bdtol/EpY
dP8YV3dhGoYlAHW94Z8b1Aa4ndh7MPyzDzevPB+tDjaj8WnYnopscpaSF7ZZK2PmO8cytZeyR4pu
Zu7jdXo2BKF7iMzUDs8We2iLnq8LEZBFyWCq8XOKUoKzZWI2R/4OnonUls3wv97qJZfvR47MnGsY
mvkM9i1QkGaRpoT/Us4GnYTHFJQGmzTW/NePV/Wg2jZRNc1GlRWA0Ty+TUs1FjFQtDA1q9+1ToD0
qqWH4/Fx6WuDUPNZVnOUffbXu8pt3kXe1RzLBKhGk1dWa9gow6jIPw13ugYkqPJ+c2D2g6MJ6GvB
GIWuWLglT0Ik7d+2BSzC9HSEfE0DC5KWV/dTbCpDx3bG4aCFZWjto5i0/KV7oRfffA7iptkvzbmu
o9eDIL/FJF06ij1oLAMf6RB9PfY8egPDQYIGG6sOFIUEAnCx/uUGQy5hhK1kKO7tw2BMCdmfTRGq
1CjEruIk0lpsgzoHqKpiqbrAs2HFwNFS1RUaH2Af6/t572HPyS7pp+QcKzRYnRQ7bKsl7eNtWGR9
mm3/YSE4qqPpNrRdNfzMdTJGMNw5k+Rm+T3BUTTQQYDfA79JZr/rrUwwmraKB/5ilEeUb5iIzXvH
o2GYy/y3bbbP/x6t/trkkpWSN2S1Zv6bPgh5HiZfZg6GLCPSqNgrKTxsHyFungDYaHDnopzIpirF
E9+RO4k9d7j1gY7QK/aslR83oa9WA0l6o7eElYStuAaH7Y/UDML5RAUuKb+O9EJsg/jk/Ydqsigs
pwJki3OOPwFPE1+M3e2Z01QXgFHEfniRrNYrMpyd3xnwb//515bJuc+T3UVdBt0X2q/RwpI1BbZW
Up0oyVy1y8E/wmLPv4D60/tXEAByZFkWva5lWfKVdmCsDUN8bu3VfPLvbcNvin3/jb7BTMonjIx3
T8tZGVLEl0jxSk6nARRYIJdBdSyCmlrpFFPI1ukhYZEm+zPwKT3huvDuK2zSKGk0EEex5WHx/fW9
I+l/+YikHhkEb5bAzI+fLmYFUO8AEsdTjsW/13An4wSSNdOE0raT5Y7t0/pAs37UJt8X9zrmyGH+
4KAGq8JNmPD6xJrHEYKmF7M08bAbknQvghK1QQw6kYKcMR8TCpuQBKzsZeRS6bZZyvuPQwBS0bNo
w2Sr3h7sJMxIcF1Yo1DiQ6qb7GjeZ00tIw5Uk5Z6eWjQEvSMcaP3G9N6dGrnpIUvOzni3wdpV8K/
SfCV5iHj4svFgGmSom3bLaW96KcrBLH5AGnX9/Aksb9YBOHzVDJiSDv5Fmyrhqt5g/RHX3EpU85Y
tjjshUosNkW55FuNvTqxhO/DLnKJjuBgIh58DDM4piUya8oRnSl1iSM3h08Y6v9Da49zifnRz8XJ
YWZr1QDfRQ9BewLqKI1VnyHL23I5VYcCDvvxyTVsVtElKlGvd6WU8sL6Lg1sYEpl0/eWSo5Nai1B
FGzwXmDjJzRJq8lhI2u8mOFo5s/mOnm2zNlg8t+Zx7jASrYrax8bYg2KoADuZLaL22G9K7BUXCwa
gKjFcKZgAfRbHXeTpSdZqaTz7M1ViiuFtLk8Uza/uUahXDaXN42cnK+TYcsQbibpHHBb8OyBfHqy
RbGqQR9lDasrObgGyEoXfq/dqlmVhdKhwEoFjXFrJWAaVjIqhbTl4XdiQ5O0W6afcyzxpOfwtp5u
S2gnkBDBGGvsun0P6pWDXj0PzacRUvpERV8Nt325Jns0lPc5Lym/+OYMXbuEn/akpQDsBj1A40+R
1yR4yS2aajSPEQZaqYw66c88by5NVMQIceyY97sEtjQl1kXoatiOrQPLIHDL+tRYdw7uNIV8eesi
l7ktNG0o5ne9Ibh75KUG1vPtKBG7P0I2o4FjtNAyc1fNMNAY4a1KNqIpXGroBO758tm94iDj3UYB
c5I29I56q81+/mkG1u7DPlzVd7RpzOdl/MHU8gzB5Kk+3r/Oez42/1qF+6RldUVbNhoNeh4+pnx4
ilQGC10y3TrwHoK+LxtRXMhZhsXaAnnSaUl2aIdplk8G8CtoSwoCq3RhHn2gd6/uET6hRFS5q767
0vSw1QINgTtTIBiU9UWpx8HvBoTFVacR/g+3F+kfqzkV8Ie1Ex0dBAnZ2TdRgS5V05DP4tQPExYx
VgMguVnQdOG7RL9/4MC9tQl5c3X8pEDLJusQS5bJDTWG669D5AoFj5qX2q4jns9+p+0IlQiv8VLY
nOAR1ARUrTwigO8uaWBsC5uzaPIHgliEvNbxKJuevjiT5/iLhht7AzhIDEBs62+LBI3UYJ3am/9L
5zpCViQmLPRO0Zqe8qPVtILZhNVbA2KraA0aOCFh0otSGu/0GT56KeYidnXh4vzhYeKmij0Hq74q
oSFqmk0blNSKN5vVuBhRkakCXYQpYr0iOJ2J2+Rbtz0ds+Ew5JlMlKcXwbjcwgCcX3wFhZZc7mIV
17NDSw9q8YqSgJ1ZlGvqU2GTMLsv1fbkgsHFuld0ivaRBRu/yVA63U0OhZNl2QlqmYKS/XxkKh3s
iVibPxPb0ybPBMnc+lODsTQxwj39Mu/GY+L6BgIyN48QBqRXWBUCabHwuDXaVVndSbvM4b05YJNA
LJ7Hby7S/lseYSP5GQzdiGyg9bHdI7HNTpkp26PHq+CNkBiiJhpAI5wh0SLQwtHyZokvhk4h+RTZ
Pm0u4fUTRnjfBZb7VCq0gIg04MrobXuhsnP1wlkiyO2CCrtvYQUpe8POutVI76ozQcko/peQMVq/
/Zt5m0pyiAPKDH1PbwmpgEG0u7e2crdUgptO7a3mzk0QBtjchiNsi4sFw+dE3mqtKbV2Wznkim1K
Gko8njEUDZTy8oNA6LI6HuWn3LzXj0OYilzix0hvOeGrbznISzVUwtpSUst6EQUoLUEWO36zrq+A
2wdX5/jMKPYKY/fiAC4BLDtJr4xWqaUHZUSRgLonBNkJ7qX7lqwetqXob5mfa5wEeKYfd440xjwe
UwF8JERbGPqYovbl20GoclizIn91At/NTHg2Z2o8d5UEii6xQorIWk4721kEUNzaJrUJTGYYPMEF
2x0ZxIJEeV5LCqS1YWh5M/Kly5mABmYEcYyT6iD2Q4jECi3kYKgLAz3C5Yen8ZelhmEocsosrllW
+PREza2wyAHchBO68gc4OBBiqbO3b7W/pm3E9azLMdt3wZYuTon/4XbNPCbeSX72HRGi3NYASPp1
oBhW6qsnLaoxVn47COiOMIdXMWVgjuxOm85e1uGog1zrshwn/P9gRfNKadMCaekk6CYwSgjaleOP
cDfPxAo871eIZoO0fLmT7y/pY1aMWVbrX7orXoz6eIljboLMdbXbHuBd5F46PGqYr8rr5klAu+eb
X/Wm9Gzbf3Jc7vRS/tEs7DHlLcILAouR72Od8tFf9ogFxiKRya5rGibGLuBSl5+fJzcCRiSTivvN
tz5j0pGUCBkHqrDTlXmsj+LwINVe7gjk6rLGF/lhx3qDir4PLYh0xbItce/09Ha7i8QGwq8jEcU5
BPf6RQsl2vazS5Ch9jvqBmHe8SxpwmL/qaDv+MAWC8mttmPYYakaOl7sAFQslz/rlkEdITZBTL9/
xKCpPd14YpjWdqERpmYg+yvngkjdhlboE4InRdX9afFwTP5rO58UtEyUC5wbOrqDRM/ADO72Xrnp
K88DE1i8HgreTeEy/qvVm++KEOs+75RpeZzPugqINaPOccmrNTAtBN8VST7qQqeG1xCYWzul0Ez0
qnWXY3Tqku1lZxezcLOEgoF3TELfzq1sFfkyOLm08gaSH2Tk1evSYaevam+xz9b7pz4bUZlQsGds
TnuFRNitVbUshgLOKqme6HD1NvzQeUXxqASGXLtyufo0xsWztHvXzz0kXiKGpgqdwFQZxTCU9AHa
qQE48645i3U6Qm3IE6XZBpYDbR5vsg+eJ2QuONiW5sPg8FP+tgbEHt4rWwCVKXv5roSlnRKf6XBv
HBe7T8KN4tBKetzUMCZmgHTSeFMRZqe0Esla1ijexPFSYZSHokW0I5qcE2W3UdgfTRtd2bbwWoVJ
k09GlQp/1tOp4HbV1sKpsEWwmieWnBonkC535cFaLXuRr0L3lmTKmQRU54lHWfXvq26xHngeBJjb
liR/IcxyyfQInfaXShxzYRkk2uEdyfUFdI+Jko+twou26FPIypzrh/ic7LwkaWe1zWIDltIAMi0O
4NJl7u4GwngknOa6ZUSWx9Rh4cQOOwITFlooyEkSYvp0LsJEPSkCGHv+6YgwwH63ZMyYU/fuKvGw
dXVjtSG3ur/adly+Raof7jeWR4UvrvIPWLjRrHvoQkFNz060fI10pQtXZSmz5G8A4NbJVi9CB/tr
70YSaT/Wpnoqi+frgliJsN6eHd4LFWTvIRiFHsORqna6CUxS7z2Q3VkmgxtQPgu4DEbeqBpx5x5E
NbRYjw9mrpX0hxxfXX7QVspA+fgxHzjiY99RqYIovyW9i3s3pf0uuRjIHxqwHV1rWdnLXzC2EsLK
3iBfOvJ9zQeHlwPJ2HghxphDzVVx6xj5l9PnTA0wWdxad1C430RkyX/UhLlambr4qGSMXDpF8oEI
JMLs+LbzGbEryQVQeuT6cw3K1yRvEPdhY//uDuCNuZP6gcoILXszyJqrFY900PR1UapQ6jcC3/re
Sw+dNcaDk0aX/ORhKGkYfkLj3BYhdbLGBDD2ow6eYgMHaNEp8MTvSGZZaIWwoXwIbw9V+UC6EkFr
JCppBAo+G+nvtaZ7X2aD4RnJPfr6JKfkmbkvhb42LBf6ofboTI2X19aVwbKiSKiWsbB9lIppmsbE
HS52uraSecen/RJTDBt41P6rKkJWey/rOTvvFMPC0Q461F9e1qGWz92gqI5NfuZgIQakmCFyoW0s
bihFQ/Jchf7UHhFmlvl8/RAigH2J6wZdHKRkc5gwLQaryO0KrEw3r3Dg66o2d+LN8wfG8r3bI/DA
VstbU4c7S+fHQhWk7Ajn6jOBtVHv22xaDpIsrOvrbezgV4jomUTeh3IypGbLj4LfI2+9vwFAk4xX
U69NDtuGRSmMhATMrksncZv0kkZ8khwJDj69uTfkiwWBmfKcsi3+LqyCB6Q8P1TBsZejXpxZG70b
V6VyfS9P1FUZpC5erAj7dlLkFpY8IDzyLzjfBIS9x1vxbUb1+NoiJv2LSoPAniJib3k/RPvTKqYr
WxHi9GWFwHp00VdgUlbprFDvqaDmNAj50LPu+G9YcnNbu9wHAxt7JAHlwM/mf67FOryiWAWQziW7
kgaSG823bVe41o9HsAle0fX5NpVMuOGn0bLabywocfj94rU3pLupzkG87Y0hYxLH73p/ls8C3+yq
cLbTkpnfNCxbvK8sb7ghHobtMpop6g0q3iFfMx+teeyj2QP38PUSYQZE51BgOcndVE95tpnK31GT
mXN0tCC6GDRiPvc5zhO3m7vFR4nkaHYm/JHPkxD7xPVb/pdWgTlzNsHYBEWCkJwy/U3ASRcuTHNl
gmv01Q3yL60HqiwVmF5dxvUgII9OHe+jf79b+KZMD1WXBbi+dHcO118YMyVIwu/dUebgX0GEZCsu
AcuR9Ka04G7Ob7sDBqByqrHIUJeZDt2alwCek1JDrQf8SsPED6Jyy6Ml8J1cCd+6VeSziumpy6ww
U6gFeO3tH9FpCKzXSYww3ODRs5zhJWP1VA7m6gQ50SCxrPvqnOvjpmI8XBKc7PQwXnpsZDQaG0d9
i0EEXRBvmne/fX9obSUlhiTtyYVrWSWm+NZoez5BMlXVPs0nEcJ6itkL7XMWidkgilxmkIEAWhOj
xbbiLKV0kVe8ItxzoE0D2pf15V67ROeVNE8YEbmcAYEnRCZwJF5GbBdwyJufcQA8/RrS6qx1/fs6
2KJaAHN4JWD0nHtdc+xGnsmR0jyL9MyYZgKc9OnbNVKUoSOPfJAdoAL0SKfmwnuUKA/T1OrI9NH1
uw0wa7+ZaF82qQPk0D8kRD1RmKGBAAE+h3L819DOOA8Bv+4CC0O6qLyTAVifbUixFASTXNBu+Y3T
iyMEWiCQBjVgoyUazmG6lF6AmhFasQb/6Mj4g7cEcvinHkllMM0EzyCc13x7Z+cDxVK5CTTyAFiE
ascCCI2FgG22Pi/13lghNx+/Xv4pVTNdXvUlTIEh/E0qDRyjicRZIT+Zq0NMkmqxdrJBAucXroA4
45QKda6m5etnagrWmGMWsgeyshDayLBWtL75h1iHt95qwMKw7ocfClVhtOhBUq+6KN6TGaSBQGkk
CWw1di1ZLrt917Org37CIhlhA5RsjtDpObjIbhnEfgfJeqHcgsNurQNK0U9fWuwGPYkpEgjDHJDP
QtvV9YPS4CGClY2UAAdrDYDbb8CWLR8kUuydfWrS2dwMLICSan3OsV5tI15xNA2TqTw/XggfA7b6
IVhGv20Cr8R9HI+/ZOJ1H1laFZTA2tVvMLY8A8fw5oECjqNBJXDVF4q0jyV3H7Y1Dhl/Dxdf3ZUO
tDq1OXcUJCz4aPvpOE5G8wKSAyCmgRYtk1XedEIHeE4vklWWVmVDRiO2JLhHuW8RELL3aY7H/IsU
cMJgrcdtJqkHcM6AjvSkeN5RLt8ttg5fxIp9HmW/qbJaAeDgKNDxIXtzVX0BC5SfnFxtDMvXL549
f/z/MVlbFE85JRXP0os15obpD5D3F27yfZZXmy6QpLz6Qt8hySf/sgwumezFia62GeB/Lq5Foe2v
3klqSG/hdwbPMrYv2LezXvmsAEzA+ItXdiVY2cI0IU32oe007l6ZqUcEAllkIL8SnimFyG8KXZaB
nz5Mh9mJiKH793RXuiqSFonWXG7EPm1JOJeZEyr0p5ezIQ0rYRme5ZllXEmHmfISLogIZXZWQV8d
cttNxRTcBN7fI6naxy+N2PQmxqpHKVg7mmMfNxSO4fo+VmNn3gYWdZvXZbMhZTPJcwyEyRYsnfUh
qgxgBABJe+HEuwxXGXePMFF0c1pZ8GuPsh1seizQKXRraTnEdJ9AmgC9kTyueKJyhsdsVvLu6CD7
bvcHq63sJA+YRxZ6f1oQpI+FeHe8CA6c2+FWe1RGNmBUUXXenJ10GFYqtxm3fMvsCpMEP/4LKDNA
+yBR960tUt+tWQxJJFPSH5d6+QkCcnJPb2P9YaJxoLmSgjH5xBD8d4GtUu2pVg0Ve3871O082ywW
o7IkPHxV+hVTpyJHtbsVvvXkLl/X2lWWVq8fj8jYVWUKXIwS57w3KyZu5EbdQwvQD/tmeWHEp9ad
M/Eu8jTFzAe9ZP5uOr6CanhTU81XwtHKW2+B3sRSlriESCPc+GFAzKRJ8bXEZL9RTQM4QMmZUyMc
1r8tEUX1KxGR0qAnn8t+39Yw9OvH+hEpq9XKddQBjIetRR25i5/o/066YGYgcH9Z6d/6pOLTbiao
d4gzh0oTcY3qVa63uIL91Q3udOaxGLdX4jexyJzHue6LKzUHiDm5G4G3ODGgstZ1L0MENS6aEmrU
E/80QNzxTz15pxW+5FPlp1uZ7jYN+qGYVb8gRUmBQg6bIKGJf4/dN2IBe3VGmxQTRK9+e0Y5bZ5g
AR+Cf5V3261Zp1xqhgmeDAusdi3CkJ6M0OAPJbP4yHpHM1gP7TrS1dXgPdL6rqKAdK3Iho/WRTT5
XbWLJV/CwcbVBniluz8GLVvIOPCcQG2SnPwzKiqWdcJ/lSP8XJAVWA1HYAwZuxlxnw3YpL4xGn/8
c/7E/tDLgX1RQXS8WGHhlyRyUThv2fQXRVa9FCIk6wxn7dcSJUpTS9R/38991BtjSkapzPYGNXey
AEKuMv42TAR85DqRLDkf5Sfn0+WPvMzfIkAigopYKnYKEUBvby5SQgzEy6WVt/pKYq3MhhuEsVdw
CteWglYJIY3ejYtNcGlQ8zH5+8Y2nBYLWDpqln/BT91H7oWipG4jOcrUa1RCLQBalswIrIjke2nP
OLm5Tbd2x2I5dSzHoaL/6SVObSp3txoLEMGR6gtgS7gJ4rJn8ehaiZoiKfgVueY53+T9l75BespI
Xbgkbur6kzbQuDiW9E0D0lsY1YjgLmhFxBbWCfGgDYstPpdPd+9bktUNSSNy8TzXyzZG3b76OBeM
JUe7EaCrJWX5Ng54HRakso+aGWG+lLO+cao33fVs+uloRmuolXOykMYZyCutjkKOloE+bnqi0SoD
Zk7E2bl1+a1XsQtNbQGStNilOTn/dSgwH7EnY9DKP/UqEkpGXHgAJWQOHykPNVkBdTZwECg64czG
TjwYGAv5bhgM5YoiPiFFVXxlbzpjbuVydBDfEDkTlmrzzXpDNie0qt8RokSeYzcj1BWuMQD3n9Ai
QhUVRH1K33KV9NR7/GNQyLDF7uBBd+IGLiGctF42JSJ59EbUxY+IMcKPPBCHrA2DvF/rrHMAWbNG
JGyiLMjwUeEVK159nwDRzy4gFpQFYL2ghBSpfWxU2HjPw9XqF378G9HAzZp5ynto+2KLfTYGvyOV
yaRg69fz5QsTa3zMgn//RgRymW8radze6GuOwNtirIIFbeX0lBiFspX2VNiju6HLdW0Glj4cYx6l
9sbjkIVJ2pAdidKknVkgWp5hsKx4cUtlQII07g99ZCRVmBawcmWqYn9YFudrsZ9VGLl37f0nVl+H
LSB5OaIz90F4DsdC39o9tOeoTvhp52oj3ET9C9viPBM5GMHZZJ72ZgcbOIr6s7l/XeXppLjLELVJ
hy8L506o/+/oP95B1j5ThMrcvBsw9Urc2Mwmt2/WBLSROaktvie1isWo+9nQvhmc3is39wfAqFAJ
lQnKwKzdV1hZ620f8oJR94ffUtA+KgYSKqOucZ2hBTq1P9dNBbcBROUqlRKXSOvFLavrgH4L4utH
+xDaWtwyOEZrqvIP05sFiF0TcgW4ugYyhbzjlANRB+nHQcNI5wTu1FlVzj4sS1BJ6pHBHlt9Dnt6
qVAynUhYbYR68d+xWo5F2huBwhoKLBIfafz7QHW+rG08KHtuRR+pQ9GpImxfUrZtZUy5JZor7kGw
TYHFXw1crln8YxAMXQxGpNP86QmPHBDyH8He6asWc2Z8lWbvYfNST9Yr808IZtAWhrHOhfuPgsIf
Bd0Omgef+GH+wtBwxAln5QRy+8d5tT2ZBP55szBPln9Vimph6GbXKl+LyGIkT7Ze4DuzdLTqDAaC
0dMi3R3MWOS36A5C5zRzgYZNK9Yb+qtVrLZAFMnIKIikg6X6uEIovoYfH539md02ghD+twedToKB
xkzvZ2CkqBST+EGALFCwtcrhvgvrLbK8OwEyeGtsizXLZk8QR5IqKlfJOd/ARjdowL/7C6iOhM1U
va6OLZZpUp11b/rWX7PY8YjMCWPNhRc0DoF0EJ1a9dsHMPZzBotwsxEk59/QC7261lB+ChjWilKH
2dHukyu5RkVmQ8WWI6LM3YT6LVNzo9KU9HaD7R2OMwwNm0qMaReZt01jpdClL24KmmK873Q7l+Xo
k58g9x7RbCHHR4wLS9w5Rq/sgaw5sYzoIUwtG0vT4ean0LIO0zwwa9OXRLiPPuRal9eVGKSvI281
b38CAjTO1btFU0CDUqb4zfQ5dkmvHnqRGnswx9O9E/TEeE0/bagQpcVLyBR09YB0KtZaHtwO23zz
KkjVJ1EWYAqvHa7zNRcj4vxHuFn+2q2Y0VlVgI6fBRVw94+qqHkTXlrzhMXUOn5VMWpraUOzs4Dc
l4m0JgpSGEk83i79kkSbO3Wpp60ClcVKRsrodQZLbCSMNhSQkK05WGuOkOqCY+MKUi6g93cFajiv
B4HNHIbdydcWAcDTIO4mOKRq8olKfKEnYqUrSOQgQ/mKoHzWqEIDiGAIReBULkOxlamO7UyiKctL
Jus6HHn2+iako58Staie7FAFdaVxG7aJep1fw+q9j/tD7MG2S+lJOKz3gbOm0RQ6RVU+4UADlFuN
mlT7YV5+uAi//8Nxw4Z28nAMKaq7mPPHen/bB+KBAmecnr9F+FS1hZ6O2VJkzFyGvgSe4Cn57a8i
XzK46+cHwHfbR1EREmrzaZA/IKwu174Jo3M9rm7PlC62uL7oG/vpHtqmDuASUu5c1/Mb8cRvIaxA
XeHdEyeP+49nxFGpW4KjBImFNTioQh3i/UUsCKaMauhJ+D6hnPiXwhSfVpax4u2iz46XyN2qtfFo
VNlPUQhKTNtuxpo9vqoLGgKh9s8UWtGUeDf7YKcIUvD1rd1KBUIwYb+v4K4DYpoK4rprgXELRKeF
MqIMGQy+teSeQsz7s6l2Tbr8Y0mF0nc3dNw8A72V2f1i0h41xasoUtm6MIO2jblmj5EHnG6N2neG
UHZ1KPnK46eEKUNMYmmZ/PKAF4+AaTlJ7jIPrTz6aX2cT4FlIrBOFWzEy7VKUWHhao70Kcvnu2If
iUK1PaMaQtJypuvKTgY7e76zWabN1ac4q9A+HqXI47PohwGHsCvjYOtw8TuKVZYDo/Zi9Zcg7P6G
WH0QI6HeiV1VRPcj1cFd1GSC8JBL50kraLa9uSgFjJwwmYAtKGqPq6ZfNxicjPgbtDAm03vEe04h
dgwQYMtnDvTLr/TQ1aiKBpPXyzbfy2gP/dbuKsGgyP8XwtBB+B/l7sk6LTVKfW6fovndXAxdd5y+
9XZejKQK4FkeU7Th6CIW9t5Y3oTGSPyOxRqEAJ6/o3gA+AYQJrlCU8c43qWsRqcTrfM/Gf+ZO2zk
wn6WzvD279V3eQ1Eg0a5Trgd5i4PW7zAk2rArgpofyaCi27Gnjibu5z2xgeg0RDkYdiAnRaD/k6X
DjHaqUVDSSUPSCi6SaXYY69ZnCG+U8pilc8anvc8biIWdhtLC3fOajPFaTE9y1AQDLh498kz9duI
EmVT/yr/paOOpGiZn7G01/jDP79XIQiRfJ1Xb0b42LO0/Z67bKxQb/v2bTnKCpldqV/4R0aiJTW9
vQ0FANQC5lbfasKcqTX3eci4gKj9YK/1JnfUrnLyH1qyZQZdLmY5xjNFzM7y3zJx61Pjzk6w+KgS
GlWQc1VMbpA2xLLTspU6E0fZCuJNN+R2EqNZiUjBXuzIOnhU6pYzxgSavMz+Szs2NJaqmV6bZ+I1
KTncZ3ZOVDvLDehpA/slCKjmUNmN92G7yOz75sGV8qEsimRnXMfMDqU0eOx9nNxFGT8+hiadnPML
MlXXUKsvypPr75GGsmQ4mLEZAHHjXYeQn0L2/bRvFRXjT0zblVOeF8Odr1vr64V5ty4XzZDEUATi
vQRI3InKIKN0y6T7Zj18m2OUNZgWC1Y69JSxNLbA/s8piAuuZudg4J/bcki2bSB4duqJgRoFbukN
PPsJKccHgED2tOu6s5Nggrd4BgQId4AiYWP7IJNkNUgFeERwNTd1u3pn7qsbAfvUyizRbdxUQI/b
8I1r9peodoSz1/oE7qWuPiofxiSZra/7TpM50dDlMMyrUlaIWeSMFwzREtt1LneUwbYkk2Xdw1e6
T3zszcNzR97gwcoZ5L4O3dfLg+W5HWm9oONc698P5p6BIS9eND1Pjg7i+9zp2/ZXB+Esr9yw2ekD
5cwafea57o6h9N54hk2VqZWc7klm8LKtq5ENU8aeQtYMApMg2R+0g47wM0A5ht+tIhF9+yPiGzlG
jM7UFpGH0AV1ufUEuCDf0WJJXJJgCINP6foYPdRDqaivz/kcCENUrUcTPts2qsNxMjp5a3Q+EN1s
j3pi7SfMHhbQmEau2jsUM/UNjq0KXdjdUaUPYqG/1SMSLr60ZuewlUsGpQ7/zPpSwLcJA+AiGnqU
6yMEPMtF5UAxdvCsIH0SkGJ8hhsa8jiS4bojO3VU5hPrRrP7z3+f3KfxD/0J1jtpA/mi8ePKbyhs
Xeq2J/gXV/u+kKO2pJjJuP26ucEwGah7GiyeOkgErj0k3zVxaRj50CuvkZcEzBERmY0ZE9zLFLQl
j2Zwpzc6r+cl2RoiP2ouVGbbmCc1DRZg15o0tbZKbcRupQ3SKH+Rs601WtNct8+FmHFZP5eyevtd
XKFw37TZGP5+EWwG33ZJIl5D5gKjRSf9tJviIypsos+GpGhQDFEWESU9CBC/d9DoqbsshR4dNUqS
iCBHFaZSD+TNmjUdwErUsphgAYW9xGXMg/ix5RS2lLZOkv4opRC4Q54/TiCHUWkPye82SW0TlT20
c3z2VwxT971mC3Nd4yubHbkUWxFzYkuGvs7/MLFOV3yoANQBJA3uJPaYR6ZLPkc+5Fgo1q+E1XNg
1ilbHzwAyDGuH3M6yNAJGz/++C6ZtueF+bZbufuc16VnVbB4Y7YI6aSCDfmTF9+iMg18v2qnZBGA
ZkZ2ALGegefh+hI9UVjfobBR5uo3T3hyv2T7zicozt4P978S4JVJRKnZmxDlWIflJ6khWlnF1xV5
frrfWM153KbYklNGrIZgtx9qIInMWU3krXfdRhrWjcW4RhNHqqJeo7Gd1rCOZpeiky0/wrIut2ET
XLUovGHyanLND0tN+mrtLYOk7e1sXyTNEsrVXvVpon2tsfp7lnl4XsIEmTJ1DiXzhC2+/irnv8u2
+QYPiNzEGderU2cfKMf/iJRqo9QHsvKxnkdpE7Zc0igpXySBwcDjs14N25q0x8cmJNCmZ4Q0stUW
9U50ZwnUXvrdQp8wIAduBwI6mQFm57iMnr6a8rHlfyJMuFo3xYycUHq1wJZ4DGz/35HGKxMXv4Pv
h4XDGq/ye5fmk765yDzgHKMJRakIctxYYHIqCsP6UFwKmiqQoTm1MSg9raXr9czYAFTHPLoskVjv
NoupQr+HUXzEUI1f8z2DIsh6e9Ey+tcvL7D8UVkao8fBuVhwwJ0YZTWpVQDWe5m7gMCAUorhmdz1
P4k1MDWUI8Tj8wd6ad0s3CHuON33qM2oziPcLPBYwrtJgCAi2aHPrLAexmIsZp4XpGaWMjcfEJi/
rS6OEXmmvte11nPaXjqkgLVX8Ue7X753c9GTY2o7Ot5nH0g9Ewjq4tLMJxMeTuvgWOjdD+d8dKt9
qlD+KvRcQPC8YYadxmz/uyh13F6hmAqmYXZ5FLj74Cow7Erg06DnPQN2cKtKHiFQbZFMKzfpuOQf
70z/uJNLDI0SWbptExxlt50ZaXXzr5kIK4dbLtTuCBTcVujljQ6eoJe9iSlfK064jX9LOMxJPz7H
kndfYEMpXsf1SSbCoZ9yLEHpxsoBCFx9Gn9CBxjDVVGWLVHfNYJbjYtVbJUxu+bmz06+UTaA1yrG
Q1fJDYwKlHr6R0lr90sihjTB5EuFQv91dLFCVRB5mg4DKNcNuoFYpoPVctoP/4u9hXrAPjYDz2Ur
MWPHsGTPZ1sypbu5FQFgqrX5pIdpGyj0RgcQAgeOpnP05/9acyAFX9B56BiVjsTrvdZExps4NLtX
7TGJr7M3FRuf5yichBsOIdnctFJYk4HfrXuD8QFhLkIDYNA/cXh0NcLc3x0glHy/SnfZZHJE7/g4
dTin20FrJJw8wHkJXpKdsTGNfuV2xn91nEcw1099XM/tFEuweVuE4BTVnljQOa5nahtQT0dfTXr8
fycG8y/rEwjr+pH249UgCfRL3u1z/zPfYqh75T5IbKCX4pqwXrjoDXkM/0Aqpi++eS9Cwd39/P06
C4GEKVVyKPrZvI2YTjSvy9ncty42oCfZLHYTOQIDwq9DJwkRExUWP51p0TP52X+GcUP63GWRjjQq
O7jUpv2x/P7ozQySjHtFmNeDrGKaMMxNI3uTgQnHKuTBkSNJAwurw2siBJrAEiYEvnpbSrkk0VG5
xoQVsPpWsyzP8GrWHnwhlSm+O/jEpMOCTVLFRbQX7AvFe5L73vP6vHIuLZ7NkwBnLrSIIZLE+sle
0av/PGXIIIyG1dYkZuoShUOBX3Rcok6c2yv+1YSI0M7pQ3N3EsabfkeZIrdRlqM0h4+ap6sNqesb
yk3aEWqer7F6mnle0nhC3HOSu/xxksv79EYAIl2ZieLxCpkXHtyFc7NdZ+MFJH74LZe7dnIRtc+q
PvcWFbd5F9mC0TzTXjGrG8o0kp/VWp+xnJihgyvRCObM3mT1PdQg67GE9Aj+C2GUnGtYRxQy0mIo
5HCQEg+u+qMbkUah3WQf3fEHC+hElBYk41Bk7ShnyCT2g++52ew7pz7DdQ4YcdQvWirGgYBsP7gt
1Z9Avcvm3V0oDUuuYn1PiDzLP+IV57bxcPhtpksTMkQPukgnuErOri9bV2nc72YhvSosjUwQ+oVN
HCBo5dWyB+oQ12jGuJLjwCqLZwrKuUcMaamlIoNCz1KBPlB3iF3Tsp7C24z5qj7nyxQFBv7edN15
ztO6yJ2/vx4EMRvEhhaenQRE0mFjKGsmMv0rlR36SMXTkvZQw6lyEcmQ9DaYpuvnxYV62v21Qkv+
Vf4sfyCdvCQC2jbLzupxf5ND4AWRUj0qm0Ml+NE/iFyw3+Fh4WdxWfZDodspqGpOwynzZDhVQ82M
iCOEJk/XgxOODZVGCD02zK3PLKG/PfxWULNXYoZO7chzmbFMbhHeiJSybJbFNB7kQbkKauODg/T8
lmMo/uYcxAlL39Z+d1Q2BOibvk3SF+99aJoADvYcF7NhqWSZsjWlMHVA6f8ll8QH6jHCeKnmPXIU
QP4L9h4a1dkvB84ws4YqLiijgLl8UpynMcnHTtDhKAcAPQanQShUY2T8Ybuk6IWKsIG7Y2aYKDMA
O2gdTSw+PvifbICagdRzWIWOvpjfTtRUf4/RnFVAhpHpsuxDYjhi3M8HvJyN+Jy1/mQg7fGmiX3d
E2VFClEic8La5Sk6p613gm2Da1CrK0qSvDOEzGtolUNKB58blozmdMdG1AZqX2fp5Sc0+TnBF9ro
91zb3aIdQE1d1KQo9Z3oGxw6fkZ1lVGq4eAwcl2PZ5ZfUwqy6JEa7oMu0TF3dgdnepUqWNmeJ6EY
vuszTSuGyFXHeMThwQU+qlU09Ilu2+pxKUzWLAPuRmEUT6G/EHIjcSWxoJTK2hLyBk7BsATTUUMA
u39WuvjEeKOumBoT7O96ktXn0ksXlUCfE2tM26TWAjMm1Iud+NAdshGWih4QFFTVIHeadnO9UwIb
TpMe4mFFM1QPQc92eq6KdkkhbT4ZrqcCsvAkn3IuvSsMgRYSDxHKKeA2PCazzxx6hSBPXF2CUXQ8
iEsgk1pLHwuutY1S2btk2WDF3+eQlyn1Y/5SIxefnacNZiTRs+OCRl711ttHfwgsyVoynsyGe1p+
BRtJDjUG5O1zCPj6fEJ9GFbpoaIcYhcX2AVYhzdtvrH97vuu9F65qiMDEUIGvzoid70FMhMa9NhE
1jwqdzkYo+jVa48nyiCH5sp34jxnRBvSnsvVCDGQgv5rlH35L/9i4JPgnH9HTbo2lOhGWtOpO7UP
MFEZg3lXuLeW9tvZ4sFz2PFgPcUnm1yCR9xUwtogg0FiHC5N7JZl/mNttTwIUi20bUU/f1EnqWtu
r/cCXfGALZgQWRVasme6Kktm/l+Qc72hTXnvTkpBmbWhTMnObOMn59q2idNUn1wcK4Gr74ZUx2lY
QjxAhzeVj+/FNn9DrPZdJVC/4y0aJCSywuaT4IiNAQmn8BGieWmAKte5a2BajyFVH9SGTDiUrCeV
rfY0VksNyuEF9VCkSwocIgLBzh7KlY0fzenBvDqMFdWs0A8ZYBjQLS4UdleuPctD0cuZLH/rJ4ej
MR/ddIN5snwcOb7uRTTlefFK3cBRnEI4phdEQZq+A+nv0q97GKzhl/30/E1U9d54CfOOpnaH1aJd
0n5jb/FK4ijGMZd8JDgYg+ogDVCtMFvK6o+dXNeaAkqbMWGQJsOGmgF7CfLMffsGFGqYdgR6WVJm
+FpPfKKITx67VRieygy0G95uNhCQ0EeylzbDPkKrCLaGpaYTWpjPbCZ9Rwf6B8QjTzWsr9HPR3/r
At20HRQu/p/UW9Cnl2HhYZicwz2lNIOq9cicpuj94QjmkmcaceAKBZDAXeQr13D2fD6iAUSi5yb2
LbX7mRaytkU+ufwU/6fy1N60gq2ZQPv2fQFu1MTtvZ4LeXFgQHU2qvUN8y7Sbl8ZlI23vQou9g/l
7A0DBbYROiBk7vnsXZAUt/NmYjkfx/OV/O3kAIF2i6tvucYXiJEtNzKRw0h2V8jaKKeszq9B1io3
LGofdm0lUuuRZMyphOjNcyFuU4h+m3f0kGTIKO2gZ/bxv5MAO2/Zo9I21rKsl0iRcv6IFy1s8Ihd
d6Ozn2PnzzeN4p/83kL1uYduJ+o4ZSh/oU7qvAG0JsrdMgarhhTxrL5Jpk+YYc5VbvKyfQbP+ig8
m/Oci45po/dZhDpI2TqMArOPG9PE8mS/BEtAM30Z7/cbvg50B0a+Zm9pOAZNvYiJpR2UWekd3I6/
2RnuC2lkI9u4WpWFWkQx00QOkHqaWIxdcn1r/CrxhnNfRa8kQ1NoB9lBc2NFF9a8cTakAUKm8hW1
RGaHyblvdsNLR3SYXHf0IQ1XQSg24mkb7EzFLzYAskKCwQ2Ko8sR6h22D3nMPTYzBIw+MbzG++ky
nehpzIKZmKxkuVrNOintwXaVTO7CJJ065pWqa/AW2fsfhQLD1YHAt6sV3E52OrQmIH4EGoMYyXpX
0i+2bqqJhYB6Q+TSFyNmSM3TfLE+pmEQHrlvNmV8YxHquk2CNlFn3gxme1BqpR84bOzE11gNki7w
zXFJuj6igQjiDsk0xExGw1KRbMjEIE94YGNbtPKqWhehFwwH1gnX2QG98rAl3/Qajr8qBy/j6MD6
34uYnKbHPSmwTm3Mvp/9bFxPu75SLCuvaOx1X0q6j1WdK/k0qUs7a3f/xuDn3YnzpuJwBmxtjwPf
n9XtUybG3e1lK2FkCNjvJW2VcS33qY4K/ibmcEVOdW2tLjKywfAmisdMgdrKer/5L7RIS/TRpeY3
1Xnfzvm+3jUqosrTOacWyfjNMB7WjxY12O6L7OSoU7d5Y2M6NXVZtMsYZ3W8L1qzfqQm7GSnf28V
8AXFb/NGqL/DoMZ7j5CVp3YpnNtrcQhJ4EOB9oCzgltA/pLe9/5deMx/BekmWlVYAMiGAsKVXJMg
HnegmepRFBazKosDzV07XnV1YoN/+MuAuGSFD4mTWtjjzddG/louL9VBmusiKwwThX05wmcaLdhT
35BL4mZz7qqyohA26Qd2LB/2IFA925+qQHHT5+yZyLnJT2ATAkrLhjclntN4YLswsHtoU2JKgu5n
8HNEM0loGnk3r9FWRQISOcSz2Z2t+L6wbZ7ndjmlsFSWn7YlNSqun8kU+Ot3q/URwFkFCGyRz9Zj
aXnynnbR4Cyj9CdltMX2F9NHZOl/LCwYngI2Y3fw67YSZC5dqNVyCD18OOgNxqmH0liSLewImhEE
tTthNCIhuFiolfpduiutbpckuYDt8gNI8YMZ6ruv8iTXdfXfZd+0BlBGxkn9SbFgi1L61d1hrxfi
w/+sQcEQ4HnZuAoDw8H71jXiY1oiewpnFPmJq/2qkjm26Nu6q8C6HQjzP7iDUQZoaFXzWpWy1x5O
tWhj0v1oNnBGSV/RNY95Xel6OIZ1lSZRW83CeJ9z0K/5x29lu0hC9YJ6MqKwvXTbXCKs5MCOGfSJ
8OFSLp3V+wHBP0YO+5gC1ruBHOXibAV1s6q4Fsot0Lbi03DkkDsxpvzrGoYquW+g9m5MuVyMH5pE
jaVDYDvU1taHjF+pmOo4eEC9nJE6zLPDbDCThwYWYrrdsuzTR31GN5GKnZ7xqTp0lRth7SgTwvHe
u5EYq2q0RkRJ05B6ZBsFSwvcg0vfJr6wGJ1B6ybjrb2EJmj7dhA8JdAvMDZQK7wvv0aqtakMRT5a
d8QFFZz3R16y9NTZZVWLmzD0OF28tNYHSIEZwxI900YqKfV9crqLhpeppvLXqW9HskHrMKejyrxJ
A/hr0PVYKJprUqLX8E0gzceio2F/V4oJRFrSKNNQ9t4oonjJba17/nX5MjOMHWkk1piR6s9BE+pk
tlY/9RVrU2jLBxxLGQcRRD1njrUaojJCcrjS4/4akzZhjPfkbWG90+KXU8VQsYFs3/sDRe3oUwDu
7cpBD2Y0IRkGK9MSEyfVPBVog2TyXroNf5kYp1MCaCovqjBRi8EtgFXk7Sk+wE4A63dnRS1R1KLO
K1/BrljPtIPEIGOxGdQcShtgv8hBuCMG78lIK5YBejCYPK3pOqZR+OjS4WExkcgBiaCCWrJRK3pP
jkjLCNRoUIp9u/chRqq8q4XK3sP+TXEdd0x8s/Snot4CKpKA27zf6/wD7hA7NGaM1isteIY0prNg
BKf1a7TwJnAaVqqcDVvRK8q8RsiZcPdKjYCaobmxHHzLFG6tNCKzUuJmJt9/+c417KOxRjZZKnhG
jBAhCwTk2k0OOn+/49WOkMsfIp8xjWd7yMpjHzuTwTq+zi9EHDhsqpFlkHjIzstZmXTho/JvCiLd
gX9M6pUlDlZye/tqRYbJ1uengs7WCcrgvYxFELf2vp1A+vZWmZSIjsLjXoFn4OEru9AhpzUixzcx
yPnadVA09wWyKsFq9tm44mK+b1SrBS5TRBte9CSBZT2hN+fv6h2Y3pPEewd8PqWB9P30uZs38FdY
oGoD5vZRsokG63+vEWg6ywnu+xCJBDuvRYEvIzjsgtTsmaEObfR7WrVxhTRBeBhYc9+JMh94kg60
dQddBNENSOSw4VFmEfgLA6iaiS2gnORqHCnzKBwq3sx10kUQwfMspHEX9uLj4eVqsS86e0P7R4rw
bZZ8cFZbdoQoAHKMX4Wpvq6AqjpXA+KMFamGgIwYb573+iS0oztxCs+Q5mL++hEgEtUL24rtYPWk
XPw0/d2pSag5m8XkK7T8FYavTFS2OTqvVKGAAIZTL6+0PidubObG6lMkrS4raZKKh5kc57CHaWf6
pUU/WrgEEV2je3UdFtpkgNkqEfCVW5ngodnEhz/nLmeqXx0XMpQ64LN8VQU0hBueV/TKa3YpHE0P
x1bGByjy1osBZgpfFDsWsFhsUfaXjCNa73uBiJOJOwclB2ljBJdjfxwHz4zVtIjdXdwy6xdVxEHi
x49F5qH96gEzOGybyS2toISlHPwMGmWrVhGo5UODZi3UYSQlwVGIheF9+IkA7Jgwp7rITEK7JebK
rAI9leF7KpfRjaxt4VcXVhwPp0YgPpQY9kwgwWCU5fh55U2dJ30A/n4SJ6zf4apbTTmiWZ7sg8i+
2ZAcBMNXJVB6YkSDw1UTrFX9huRZj6K7TG9Joxjo7aA6qRXM+rslBFovgchgFkDj+zjmTtQ9owCC
xiP1IDU6ZKhKbuKCuez1ojYxbncPWwlBcocvcic0bWXmhFtdKOYzDXd8EgAmxWXeRgNiD9WbraLd
KenxYcm/3i8Rw6GtgdJ/pkdHioxGl0hXUQ5yYBOzAIY011+ZCfDuJv3m3q65a73REXTVXF+umVcU
A5/L1QCrnPL/IgEmPUgoY6oPGu/0GH3QGd0s1vfNBB1uhwjFrY1a7whGNkswvlDjwoF4g2iXRuzn
YUsO8/mPmqummHCx0lFyL6SIasQe5jMMhOmRgCPEn+d9xz4FVtVtJUuBrob+WLvdyNhjWkL8ltk9
Id82oYVRAYSLheDAs/jyoJoLCekFFbDBr1LJyvvsSyYDcUAWjmxtAWwIJZIt57HM12T9ONJCQN5A
wdlwS2oU7FOEC2Wb7RC9K7H6Nk9OLa2HWZZ8bCn78k9ymEP6FB9y3CvyETLo9qhY3cTtLGqLFKy/
+xp8X69iNU1jYLdIFusge3qjbSxvTPIb70SPvyqqHhrBz8yUe3DgrbO75dOYr91bLpTaLZVN8iSK
c2LS9IhnDkS90xxo7p2PVYw7AM/w7gNYXvKvP+hasrR8NcrGcpgrS64P3u/azBxYlluIYwmBj2U5
XxCVWnY0w8TU6+pOeS/ewZRhPk69semfdyrek6ym24AS4l81SXBu2QpAhJrnn32g5aNj+vuefmlP
HLg0riU6wMgt5jLZ+9kDVpzVC1Oc64SMctt7j19ZD3N1GHnUMeq4mY721HvEzSYD1QoM/M6wYOJX
2RQfVxyl6dNGoaPkcp5bISIcj/g82pxUW/hUjXnY5LfL09+Kl2ynYanhHlreHd/5hVnmAdZTcrdA
hJMss6+2Os7Q0wZ6LqF/k1hFYzGrPg07ia9mCU4kLUspETYtaa47yW6VUDD3tyBR7RX2J1k6jaie
wI8tGz7y3iAug4oTtgIEHE85Og6pxIRo5pavYwQFL6O2G/RHvK5+AbDe3jaVLi4BlJmmY+fSB1Qd
dRa7kep/CX0EAUcfzUA/QkBNo0kHHOpCNWA4Pis+PHAnXpULkVT2Z0YZq8XOcTIj7FrD/OhaViso
uYkk5gvI+sox7fsy2/vs9ScGPZiBAW+8RCcyPxZZZFcu/W+yFvAs77TIQ9E/8qm2Wzb7F/cvI7KU
ZvoGj8zLT+FsOje4V85fVOQ+3q5eeXw0leWQWqagWqJ3ml8l7wQBnpd3sO9ZOIHssWVGBNfeL8US
T6Lj2R+e07/rjmHB5pX/A/+X4yeaGg185KCi8cnf4sZ9A+6nZ7IZ36R5NuA8zbu0GMr8aIQNsWYN
1s+Ec5qPtm35RZLCJHofZv8UZlb4ETiQg4AzitejdbqBLpksYqqRPwl4R45OEaa4FBXKGugKgbhJ
TDcTfhW+3kicM0gUFVB4o14JnwT9XV1TdQsmigAnUwoTPy8AEd1LoKhbsAtBydcg+QaPmLhYK/+D
F5Z5tJl9MuqRoF7rh+hJWeRrHBgwt3qOF1QpjdkpQ3fpDiQVVk97GEk04IJaQzXU/JJ7U32GBYdh
CfZSeAEtsRLpVXRCXAcXMZqO4eLeQfA0wb7P5K1A7NQAo8cJHZISpyn3pEVOEzSegnOCyQiaKpZ1
B/IX1eCbIFNIrjAXGWGf4BUnCbzSqvaRY8jbgR0viat6+hBrOKa64QmpIugyh1yQxCmCpuIpEPqX
ZmqPJDTDEqPc/Q9rK3A7kwzrwXw8Ha2gnRWldyemlGTeS9xsSx3Sl9HUNOFXzwr5zP/kRmbFamnw
JZ7DHnMT6vC8qaRR70IjFcaHuPPX9pc9fYyeGduEofldZotKcIBbtHOAT9gVfFUU8056M/vqBJg0
PAQjHVdFCsZBTDr5FYM7LleS2IbNsf9rjPPAXgCv0+vymxC6/mLOzI7OV5QbuxFyprU8ZfyRUoxO
560zsQosmZSRS/ecuVgWVKnlx8HDNUpVZaXuz0hqfjLBGr7mfg39l1pwegk3lUGDNVuNDgHTeCqH
AXAz6UTXpMJiVZ/grnNbO5UjFnw2sS61dBbT2coDDqBZgk+O4AzKCP4EW+rWU6fuE18E5k/vzozh
lun+HoCMcf0KtDaTl/CRqaLr2kjSiWRQkU7BXsByjotZ5aoac2fPzHTBBJM0TBsDctiRbq/d+ore
3gwW+cq0g6Smq9QVx4FelocbIBz/Ws+xJdznqPdpG1yxNGf5X1QIJ4OW6uE1xnvPEsyszZqs+t9b
yglZLkcrwxzEIQIxLTw8yXva/5D9tgiIRvzwvRrqCzfPrPT6LP2eSAez7QotxrG2e10K/N957qMS
utJXV1Wt+rYIyr/w3xXVN1JpoRU0Z8SE52pTtUGaoCUehw+eLexCK0zoxs79tMWpO5iz7ngC/k2E
OLJPE/yVaxyQzhfchfPWdDmhhsv7DsDx4Pz/XlJSTYbBpS7OaBG2Gi38G+qiPixJqXfA3bYzwTJv
HdKAF9XbecvtjRMre15q8OrG2PKWcF0tqI7dfBnqUzoOa2s2R+pMQW1FJ6z8D9+7+Q1sGrKuqAwX
4IkUhL5Uf2JAN0UFxGX8yMs2YesMxIY/KFSZ4/zFTi2mma4VAlDkLvHgdJziWdsI2MqR1VLoPj6+
MNwbwXx3Vc5uG+NfkkqItBtHreGGlc4kbMJSblG4L5arfDzMA7S32Pa9P97zf39efPwcDuyhyG7d
qz7k2Lhgwt8AQRigQJxP2Ta+GlRGGOfmPyWw9MSG8M8wcrj5gUQ0/t0fvjM9H65IFP87d57NNdsP
KX5j1Yt1KGDFNEWO3PSBiWFPklL4LFSyWkrTimYmK2H+LUmVocoa/eYfkNdQ8eoySwLbk54B/L3g
9rMcAykk2eaGNfIhRfnDc4ukDJSCpVzjy53HjZj76o/hRCCFBifV7uvOWFP8OyMABLAuV9qXAv3k
oWpLm7agXb5tvtmgVyf77WdIYOt0jIRs7oMrrun8le3Ng3hGg7GBudooSkMkgp7sEeN5zfdyfFWI
3q/VHTa0mUD3mfo6S/DYTpzjWMp5HN17ioNjTN8OEoZFzpuFNXkTGK5cRzcJH7mxpfMStGhg5hNS
GciC3UV+r+GSvpV44rEXlkzzZPnzmyZ5+ZaCsGGE2PORVMbNCC5bP76Gn3oD1jTGDkcu2h08mZ9p
pG2+klR6CLCtXHcRkYEKqBu168w4Yz1wrP3GGKgdp360HhDPj3FXIwsbQEWTZsY7WpPakimevfS9
OcpdiHUyeukydOsOzfDPYnLYklR3fABn1pUE3q/aclp/lYM2EqVTUV/Ewe/bPC4JjtZjFtN8mWPu
qj+CgI05OQFR54Wkp/ShpZfS54XOVlW6k1qdUqyOGXuCoZQdnODsqxtd4O0cSBsIIOD0i1KMZfvE
lx2liRxyEIBb+aRG3Jw/Q1kvt/IXqAqPCz3UEQbEqbcHxVhIAEf3uERFCX895OIVD20qkpMOxdHL
BjXvDjnHTYhPbrcxuAt6lMb0vRyZ55qXTiCBbjQzL4A4+bsxbAaY19b5ag1pV0kxUiJgGLPgRyJo
7LaO+fQ47b37SOnyBOMvoR8+F+SkYufUP5g7Fcml1+v9s4cMMlMvv+M87ZC+N2CkIXc0QSddxM0O
jDkVTApxCiN0bGgWYDIVbwBtESl6yF4/kCEJ154OUusRSbA8tD4vYGXEniV8nGIrVwDTvfLwrTTd
IwO6Z7aF+cg++8LWg5IMK/5K1D94W9FCLRGyrjBhk47eJ7NW8jyFkwSRCWPPvSU/hZD1HheLyhIP
2P/5GiubWhOC8RO8mwhlAHH9cujaLo2Rlyj6pdipuF51kRK45qJMsfzglnWDt6hnzbJOVtds2mZc
t+7Fs2KFbv6QIhhArBFgmxSv4O1MMXCePpAQ5dYknBWrGxYIP3zUBoRjxSAP3t93KCzodDEX5BmN
zohnisE1DynrR4x1CL/tnPbHTGTuxdbcOA63AZs3/M4zF3V187W1j2h6KhuV8R0QYv14RtqgxZT5
jv75jlGPCPiNKYamrTaPrAQvqbuopcgI784DO4Zk+m9BSpiZeE3kKn8A+y/EstB35q5JfUNwJVPt
KvbbXQH+LJ0e+oBmXd8GQywDKZJJZNA6qUgo1IAAnrBi3//lbdnHTQe7FZxpcgXQnjcISooAOHSk
jUEFm1B2wHTAZtQtvG7+2e+nv7ksITfbSWvqF01wuZHZ/+wTXOTVeKVkIcJTHTderor4iJVLX11A
IcCqb7GfGKxTDkiC5Y4Z4lEnt/xiXHk17nGo7wiFRJ1vbStdu54r8jTVUuO3xpKSfviRM8CWK0yy
MSPRR8Pzy3XZd4yn5pM31LIqttGxK/FE68aGNRp4sTi8lh/sIJNrLFyQwIKc/SAu5iwvAXoYcxBs
CvQEyMjhiXCQmBI5dL0Tft930cDkKYtksKJT8eHikjtBOiKCVP2HNhbjmWbDd1pGkt5VPWGzGdKD
0T5RrzJEtVO6ew3/VWzBGu+7dho3xVI6csp3QbvUqwsGrhCy8apeMc8oJjed20HrVIN8LX8GpKGk
HdoQsT5iepB58zt6pTYeaAjmLbkKZGd8H2fpRAgw70M7jH/mR1yr8Q1BgEwr6tjwv8jYxNkEvCkH
SVoEACNcSgybWwGk44v8+lGrIVEIsghIo1eruMyEBDrJNFUKe+0CEqIhBZzjdq3BM+opDKTXDN34
hBpKICCBIHhSGYMgvOMaK0XmF5DoUaXo2Q7YhUIu/MFIC/6mH8zGA5aGzbWR5wYh1NiomFaCICBI
zSMikFHRHey6ggL7tCQ1cjOnIlTTUVZbDWFTj7q+55RaWKxV1ShYrL6Ddw8msx/rdM3iWLnjHAin
bJrOSZVFNqkkZ2VYWQ4gBnN4uSXrq3ayCr63PXLnKbnhcuThLyc4hif0zJ8PW6KvG8WEMOqPrBd5
o3bLdcTYew1x6G/k4RV/y430I2clNhc/gTCD+gKiTAquY9Aqk1PGN6w7xHZoTPogUWDoRiEsWq8x
ToG0tHLgOLM8rnhJJsX/cIvaBGIIuHh+5nxCJp5bqIAdb1GKcqViUxSl5DLNnD0dItQCoejdrTYS
5lJDKhJ0aaI4Hgh9Df270ZLSpdgpSXy9/ud9gDv5z1N2fyXbaIqIcPyzkuClmGO4+Y09sgV9dKnl
TM8u0GiX610lb1HfNQ/RXhX390mrPre4Ty4t4gnCva0Yn3QTJ9kKQX1zgFTH2+Ak4VmY8DWHol7/
uuyYpNuyoc9JtxAMDl4MmrNB/yrRyKUd2ghAt6m+u48tN8CN+IE6Rv7m0hSIpoc6eFBOi+KFjT5Z
w03BZA3XMMFjkI9URho+4bDUn7Dsc6TmunAsx9GAFPJf5kcTmOjC39OFFeS4btX19LI7AoR2BJLT
wSBQqYMHeAJ/l7yLg5MMtKhmoBDNUMJiSJmxnE/bwL5TpFM0uPS3xk6FI9nI1SY6xSNPbm46dqFz
SuK6bLXJmfrDPME3UAyGcLf2P3hvjcYLrNzQICby2DcVKVjcEH6Vsz9GPhkQSblUN3rGqI44aGfJ
Mz4CrHLj4STuoocqpfanTCE/JQILAYR5PwEeQ1HQnjpOsJUG95hCjqnN2QgcRx2fJ2yB2E6BYeSn
FEHBPmJVyJRNba3gQVFidzSL5P2yrD2DfAiMYIqe8Gb0oRay118IUQDyawYKN2N9yiAWwJOGe2Q+
F8cYBFZ1M4ktJDrEgcz3J2ZXYXxdLGgJgPaNQ7+BP57rgU62K8eMHcZCSti6Zrk9z+PJslUsXM9D
2YGhj3z8LLlQygda8M7TXJ+RVFJEgeVYdGtbuF0QqtaTE3EbruIsUT+i8aXoL9UcpSjO1FKDB5O3
Fn+2umJnaZ8ZRh8gOgR16VHdaEI13CB/thRAkMQAkmfDPEVvlRi84MXBBCrzIyeKUB02gxm4fnBM
MIebtB4yOd1MR9HMHxZx+dPTGoZUHupR8s3cmIGQ3ZDT+pNQojuflWXkTfllSiGwHRxcA3MxFx+A
GPzkJ6jJ2/17e1iw4wz8GDWVxZajmvQII82RtDX5sKF5xK4JrmZWbXw1YPy2MAvJKpMIQ9epq3K3
t3ISnU+NoPaEcSyeRWT5SpAhCgtuboV0y3+OQu4sCZp9SOZumg/jQFuIJP/VlAahP6yHEKCESDPy
DtTzV2QZ3q+NgiBVTvESNB29Aj6h7EDMeWQ0Pg7Sxupvhhe39zv+4CcKTIf3eiwW2iBfK7Osufbv
xPubahhabUBxD9IJeoT2kQKJ2wJET0TmuIlFnKYVTsJmsEpfvPsUsJzVIbuoiQRY6Bhmbx2noTtc
5l3+6gccPbnQGcbD9azn4E55qNQupev+eGJB19vJsZGf3TrWY8xkRwin8ZvTHTAVYmRVzkF4klJw
qOARlzAfFM1JcnkixJZ5xHfJrdaMNEbeAxNftfpyPe9dTvk5VqXXZezJW086y4EoY5qn4le+mzFr
jPSDEa/CWJAm24HVKBmk1Noqmk6C+WzRfJeMacF5v3fZ71MuEZGM8OxWjgjKcUZgU0351+jhT9KP
bRwheslbHRZALROs7X7o4pZzFJttacvvvEabt14mbBZoDowm3U6stgzSUfc6m0VPNKb0B6cdvAn7
PXBELWmEqU0ii8LwAoDkQ7adShWqKabmKUzHBKv+5Ee1LBhp3K695DW6IQL0l9O7rU734MY26nE9
hVNj2hnqxvkKmFkcqFKDUJLcOqVlE1dXnghA5UMRmY6vKysLj2X81053nDWwpVThbrx1AIKktWl4
jB+Ou1OzkyAJkJSnqxyt4tFc+DAHyzFH2Y9k72UEckQQgojv54gBBoHdvR43rJHUYhEWCnQH8CUk
sgj49YhgXWoiG1oIHf4l3n6NYL4V5rDrWflLg0xEZx2cY7VziukwuMwIKxXUjh/0GEIaIB8E6jG7
phNahhZWHVeFgRkWYxIgzKP+iFecSrki3JHUhZ++Qz1LWMMuGHA9KXpWA1604u4MsSBEs1zfXtDh
pwD/Nhf/7q+RJ34wrbFkWUy+qLOzr9S5IPzjMrgvvI4n/kZ1RSqDJyiR6sAoQuICBdHbpIVUsxC2
oJRjkMe+wRRWQE/TndnTdFR7Bm3ei1IYj1PYNB8/e5Jnkgqp0oTJWufp+cwDnV8T1JtVrI9puFbu
LFOSjlyfzvw8jV3Yxr8zpx24IydWOJNtmP0DkRzkQQ8NX6MfVv0RvoUJWyaEumqLP3sksapwd4qD
KU84j2TANoFdLScDq556vdVdXqM3JwozdSHxY1UK1EEKlKuPBt/5ABOAc++hIlpWzOPQNo+y/zpJ
qB5pJY7kAUsVuoT6808OG1zaV/2ErxaHk/XJJfH8k0JlyxzQJiak01uyaQRpoZODhySY3IhmJ8pg
oYh9SfDonObTarCNu3m5xLm2j5zkHqqOv/F901VFJ7Bs8cNy13+xWRZzNXd8ZcwFj3fFHdnXXbUW
mfnpAlr2eed1K8btEkoQCPZwI8UR0b/9urZjjQOmLTiTHgV4sBHaYvmTl/bRBp9OW17JwNFHqQ6B
JZ8TKDBg12+jvSpI2zNmkSWmoV6I5Z0N1+ajr8fu4fwZ8/nOkv5mCB6YqlsaXNQ7zSb2dyi9swOZ
WpC4HMC5uLLze9iplY+pGeqk486SLUycbn1rGcZ2QGF9saOzs17iEpcwmgD1b045DBjLN4eNZl8Q
Vb64QO1gznsSGu4d8rYDCe5kmKGeuv0IEXPjfmC/JkIdufB4x3FIoDeMzXUxY/LInwOnIFl6PxIR
9Xi4RAG5hHLW3XI6c1yotdAFEXoRPQFEtbDXO+oTfKUP6fRG/C48pP7EhczpaWRPQ57Yo1gg0dWG
307fg7RAZhAcnKp06tX/w6c7Jlm/lFAUiKSSTvBhOnQU/NgCWkhLVTCXdb/S9twYGWzSj5nACVzi
d6fC1BL+EzueiGaTvBKqVXYuMyyhdxOd5DKoWWBTGh75B+EyBbknDqXXEKTZ2WYUXMBtm1AAX7u+
jUwbl6+qHtoGQlQVWEqXPDkFZIBr2pa0lJHkluw3knHTB+rmfx6j0rOMIjDBpJQJFuMEhUiquu5w
S533lB2ayQYRZxYqtA3G3KJ13Ndfj+XJJM46bbwg1xOzNQwIhIzG7FdohRkI4nLyyECan9SktXOw
YHz8PIT8OXdQ5akYNK0tyGv6e5EF+RWQXxtLUkEziEAHnfpfvbiajI0TPniGgGF2GrcGp6nFB67u
dY/r+uANBm+KN1D5ZmgNTjMqyW9f0YRjv4XQ0mAOSxFGBU1W+hXfsGhFgQ4rwf/ZNckEVuhRNOiB
K+QlgVU25axZP6PtgxcMUD1yLMZDS40IDqqWY58Yn8RTVt32WN8ynMBjMWR/1pEukgS1Nu/jIZDI
iMPiE1p97GCwNsr1dPhwCsOTMTsM2e/PRIwriigWRXmCCjXz4rroEVhhdDwudkEMIEIHBoV1ZQca
j5mKsPHiNK4hi5bxn7gy9xJnA8YLZOST0ba/56dbWQyluNHX2zMaPiCaE2L33Ykqsnv2FIVdeFP5
beJUzbUaddJC0SfBHDnRtSVwGsY3OY7WKak4yU4QNvqwmma6f+tsEpjirLXcJHIgqX46gaX0i6wE
L2+v45LLoV88oBGIZbK5Sgw+7tW3IN9jfnjc8Xx4R7YoSiP/QxjuVgovNZm/ZJ+yqJZwpUnqH1KH
cLR7+QrKu5Z4Ddpmsl6OXV8uh7sapbvdDQ/D0MOzJ5KTB+OPaU5w/gA63XcA6+k3FLPbiLbmW5Rx
No377NWhtGP3sseg7VSQz16Jpf43A4RDTagwsWBgEfXPAKxYaWQCsOAwyRbL/3hH3QrJvDdxGAjF
miB59CGCCHJgvfqP3bOYxMVLO21wkXiIVZ7R3dnyzFrFmUT5xGpyOdlB8U+byQrBe5g02zT2YVVq
2fN5XKArsuaQYGZksj5XKKfLh7MlZxxdt8SpbdC8X8zjeeEN29NYxv3hL6WSX/fZEu1i1h/4rKig
G2KZnpBCsOQXRnfRcy9wsVHBtiIda1ez1dTN0zyNfQawkgDDDyQfuOAJfZAAwdujqgU9/xURtoLw
70nJet4XgZDt8NZAVqSvgYxnhnWcekjz1DkabPZxt6IytxEBKYNtEX9MkKxvBYiRn7ktlaMiBCFV
gHpi/Bvjg+jBeGdVDfvtOB/Xbq0vpvxqc0DPOcVe+7nx6n5H8TtaW63BCqEKBz0w6M5a8jaL1owV
ogNT9wB15vEfpOAeIQUehuylpWFZYlW4aatrTfXFdC9D9E/55kBMzx5mev7ZY5vyFmRHuxaliy9w
KBOYe3ah3HxZvjUxh9pXWLSbFL6GkSGOFfeFejbQS9cBnAhS/8I3LWHwXSVHJtRojohT1t4KPLCH
/Q5OVgm3TSkN0x/rXX+++YC0nl/Jx+g1SemZZuFcBvEyGDqNWcqHfuWvzmR1PS/g8/wZTwrpyycQ
LNvsKT56wdKpPVgvgznLkLSSe3nwYVdFp/G7fgwhcoiErjaC1bg9+KqIkazNxsY5J3Jxxj4UzGtP
8Gdxqho3aD9KUmHUFuEqMcywiiizHL4aNP6QYWzd2i6DXk2PiUIoIFwkghSEictTgOzzTBx4CfBr
OdBNMBUDGFhQ9nSIEbkoL2A5cqvVRg6tCeBMbLlQbGTmcILzYh7/xGKEKVLq1EH3O00kLY1X//mT
RDbMJGIlzgFY11G/hpvToKO9Ic++3n3NvVx0Vwc4BJSptTwkDGHzAsAPN4ZuMWD2hFJK0JsvWPQ4
Ml29MxjrJxDqxoB+o6VSTQzfLVPAAe+aoNGpxEd7FrO9UzyKNnqEPhnfdOgcWoITetRlMzJR8Wc5
/rVYKs3Sx6goNMTD0MeBYEouuFBoJPhJOWMXAT0IemxkHE0/PGB4kiqmsVKLS5S7W52rFdJE1Tw0
9rp9bQadrzwfM1QlXgH7rGE+hcqKM1iFJekQGQSXo9V+5gjVfM05bQAH2CUoD+KHaXM/5yA9Ka2j
qMHhKDiXoLNt4LJFV1lGNn2LOjOMwMhPH3QiMgqumY4sIcQIKd1Aut2aTrP+v9xv6HJQmEKiOS31
5DPjAxWix8KVhv3mWuIFouBK4XD2nQpApr/Mj0Q9Ul5GHZhdH3bOtSSaHtxuXVFpgPaiDc3Tqq6h
T1EjevnQBPYEMJq+7J0dgc6m03pbY46gVrieOwpmqOu7lKh/P9XiWbx85jxvbNg3st/xD/evhU/m
t/hL/Uemm2rkVTqEN11UUPaRRq5Gbik1wlEG3QOX3Xy/nOF+3peXToHlXknVhZtBA9u15SFBYEFj
Aruaoa4C1p8wymr/IxwdIs9xEwJ6qSeEK8IIPvV5Q3+73BFWQHeNLRwr6W2XFEV0FuaRL6m6zIO0
tKwDaoNqZZKSxoLZDZ1amtY48TRS0U4fqaH/03KFc3K4KkFJjunjdJXwwR7T5nktA47yiUKOgnWu
9KuAXnREgovKPL5Ih7QH0IMqtMxJK7jXHlsSRrfPv17QvKdmOz/thg8gcy5JkdxV9kJOsWxICCCK
13JZGXiflIPrpMPV1PWk/a4GDgiwE0jiF+hN0G2VKFLSscQVyUf2O8bU+BqOw1rDG9xvUJHQrKF6
4KlOYmG6GKvu1HDSnU5fmy0crvIOHD7Rm6kCVGnv+3B5wH6aixbho+z10Y/38Tp7dwg+tsmSh2io
xwyk1q594t6zluymTBlWkkAkTY6xSOT4ihXn2aCmsdDKpuGeVLhG8IXXU+/Iwk+dAoRQFSy/LlJO
xXQQYPEQG2KXTH1UWiN2HxV31aodW/kMiBeQv98dsyuhF/ST/mC/s9DfCGN+hPs2VU8tGWjAaQv7
PBdtk5NekcV65Ty5i+usKzRiYuqrRN+fNw7fSO8vSxS+QuduGUx9hBKZ36XKbhhtAEpsN7VOATAE
744OmEvohP4bwBdo+u4WLL3TZeP0o9hJ8QuGUdBQfs8UkIzQSUVvir1VeSQ4GC3j3SkQ9mCmBso9
w1vT7pJb5ASxwTWmq/EVEStLTvdxot403Sdv+Zno99DNzlGoMI4joZOgJN0ASdSL3IP49htvRWOM
NNwB664+FWisQSYWj/6sjRrUc2Oe4dFzGniugFtKt9CkQnu1Jj91MnYsjrC9zU/+e9cQUhfjdb34
oBEDbtN7Vk65er/s80G12q1n0aOK8047eIwOwedyn1n2sJwIDsuIBtJtc2PQmer07hsSKsMl0cQJ
Autt6Dxluuy/6uAHEEINTOTHKZ7TTM/d3lyjxUkOalFo8QHlpWDjEEo8Q+HSGbiZ8D+3aaVllpGn
l8FP2BANe7nFwafocRC8dTDPey3FqAy948ZE7Yf18tgJqnwTUPyWKSl44eO56TEeUixY7ixzFgAh
4FqFx4WrhOfJGJw0uSrt6gpNuWk3vvLUQxr5LuLphqb1e7VLCPh9TxXtTbL54qBvkr4KqELZU4BD
pBYZ16yOXb0zz90/7rYnFOQThPmlZt3ehY2a6XbvsPbVGZSE0jpMB1ZXyCa1kPArWlf30kPOgw2L
hx2C5EbRlsOrJKjx/oQxen56VzdXh9TFBDcVUa02mw6c2KTC8UIA6av5PCH5qgmhVLDyDigm8oK1
XC1TBoq0E4QteksAk2QN+H17mMlwA0MWEwZlnyCwXHLFY0VA5c/bJpWUc8RlC0juUYmBc/0/zT57
Aiz08RBhDW79VMLDe8Aih7fqyPA/M+g1rEfVhYTHKGVxBk4Ekf0vbQvFKvMcIKQqmZPyAkh739mJ
vX7FFq9Qr2N31XIbgaZ9GANJoJ88fTJ5lyqzma1Dh4dV8PR/Ac8u2DXs9MRQwdrfPWMghQNuPwUZ
OaM9HVXQ6jZyMGRlvNcOfJA8rS7C9zt5nqPBZLBktP2R9U9ac7mqkBqC+dbt6j6yxE1NML04Ptke
9KoPfrVZsgN/kcn7WEBRjEF0HK5d1M5f35d0zCkHhLhZeTexzZkrznpgRnMSMKqP4CfYyq86vj+9
LBS2og5G5uqsz20Aa8+JP0Kt/3uXRuIP8v/Q9MF3dQVEQG0v8JtKmSselUYugcc3FNbzCdJA0pVl
IMETCa6ohoozJOpPP17pc1SHl+iwW06mReUaB62TTtMyp/bIjMJFirUAPe2w24CQVczGdhg0KPF7
lp326WdtjPQgIkqxWbspGnni7xkzgBth7fuP5KWE3SvQ5/M8FV5wD8nxR6wZ8Q9cuOs/rZyfvGUZ
QMRYOOfOIqh0ToA/FfdGyTczHVbXDiofAn07OaHhpXqfmA5fP+E8Q95aOyEQrllC60Ql1XCp27Du
xm13MkGbdsbamNe8Ulv2XJeYtg4roXDNSq8DM8e24c1fpTkZPv2HLaQ5Y0nG2WqqzCmDLlLYwsOm
SXzv/bWVGr6bWIu1paUwBBQGlF12w9+lMZhj7g21k+fwFZJ5yidu5Uoa72D4kKG06oinKmRfRumd
0vZJ0pFamGkUiOj1D9DyCE5U6OmSrV57rCA2C+386zuIB/Y6jjJNlLXJ4gjSxUx28hXUN+mornMI
lDmiWj8qqxmF21XWVOeGVJXWsbo8caIqGJvzyQWVq7GPCzfBzayubrUALiKwbWOkOQL55NCM73uq
/6876idBuGnwwvcQjRfMkJi92EfMYfBUrvC3RkX3nDFSWRdQB4thv+rxM7YG2Q81x2pr+IgA6glD
+GROaQ54pug3E3ODa06Jhh7z4qX6thimr4E/Oou6Vrea7eLLOxx1tAeiT7XjR3C6ed+Y6adbqoK7
22JRfFTjdeMytutGIFviSXTzcFoJVgPIizo3J0oem88UbVL9hlNGFkKVqghkaObr7rG1n4soeW8Y
+/lX9RyY9H5l3HfEHOGsoJ78ztfRrdnd81U473i3dWgPimOLbNt8LStHeO+aHDs7RGItJ7p2HFqB
VK3yhQ7Djs9MtsUKOPWCrEOVceyC3prkUsOywTzr7NbnfrfiY8hi/p3XGhcuVZ5bCmFxbHNo/ShW
paX4Lh+vKnoepheHIyoMFnQs+mv3xLPJtk572Ie+VJimRdgfEQPfhrXozlG+YG29gtAsiwjU930e
iG4HmKC+kUEP4WBbP+1GYHj3de3lAgrcF54fpx8lY8GinIZ71gP8vHfRjA2sIuxq09+sYAu3qXrC
DDGIVOKyXAJUcuc97WI6/To3B7UPCSDRwOVYdnVacLJZB1fXSIXtCYubrZYz2LSoQPp1eA4Dv7G7
7uIEi7BmXZmWLXarc/UJdxL51rXSloIlG0x7MxmDeuZ7HWDXaUYbUdls6xhGYgB3Ydg4vJEhTQLw
jqIo+F6hnQVn1k+JsouRYTaNfKwcSPmbMwbfssK8hFJsFD6NAwmk9eXkHf62uG29G6wnrtnRQSak
i8eMsaTDFuM4BXTSEuew11YHZGKskdUuPSfYHUf/nv3Mmi4dd8FiCiTq/sZRGZ13OA5/PCtfvIGd
45Lh2fyu/4suT3O3uIXbPkvJcUCrt1P2WKtypFw48BhCs335fFj4AUjwQw2FdDd0Xkb/612siWbg
cBFu68Nf7btYXmpD5+g8opRe9eZm8TA5F20yITMPZAMQktNYaPZcR29CWBumXQMod4wiDGFdHioY
uf85KSdUEbYGB1jnv18wovfbVLGjxzphkygwJ5IVXrixZGKo3X5+1ea3sCdZoMKHSrdXFTr673on
t5DTuJt/iwwg2g9zXQUiigkz8oiq5ZyHt0lnKM11ViNvzogDq8i+yUS75UrOzzu7LxhiJ7oVm25n
RUgjTqAkMkLDAlsbnjWsUAziPuerwQjzHVWUJSAEqjMgw/9eFZmwV2vRwoUNklAxrFelrZ6NSiJH
PniyWS3G9kQ0isYQ7s+am3TlrEhC+d5agh96bWuzvmcL6g/n+8uxTfiN2+sxbRhubBigZAaSDr1v
Shl6FLLzGnw2QTbFanXHFWQqC7WkNDbmsYNdr3OoMVie5LVCHyjfRMcmLck=
`pragma protect end_protected
