// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
jgLg8u5lcdZqOClczw/v+wPCM8a/A2HzFDTNMLHfc10QwCllmAUWZg0KXDw0
uYgD+3Zok6Q9teaXiktiXkhLQmSYyB7SbGcl9g8wWp/h1xJlfYj2/VtY4saR
bbPqRxTfzRmauqu9Y6FvwDSQ0Os/+3DQ1cnjDuJbZXRViQaFC/ReXmC0Bxd3
P0DK9IwwMfNxsyZMxueakQagY96VUdfSeDa635i8Y3/W22GIZZShzTU11T7p
zllXkJdjY5H7M/bm0F7e7jZdEDBBPUS4iIxppul6tqKAUTYjdAaapMHIU9ve
260LQaLiNtqIxlWFAlgp1eHzuJnnONRVBTst+uaYsw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
nE9qP5Q2nFEplH/IUCkhnHOz3egmNXPUpRRwVHGBYWGgrLUVbad6FvvOj9iW
hrcZnpckBZ0iwrU1pmBbyChY71UcoAZC6MDmzA+i4tTww+8i6MdGbl7ucQwZ
Dl0m/4hQnlGR3g/AxTD5xn31h3wkLyN+/k3s2z1bXWNEaAtoXEKjSD++mrIX
/Z1TpmWBzvNeDijXZE1JAFYY250HRoiyMLbROuGae3aF0eJVwcvC9p80ob2m
4Vx7/g/oVo7e9DZL9wRbU6/0d0RuDZeJvu8yLmkDHMZ7y3H3c7adx51W/Umb
QpDWhhSRKLJYlDGbGMyQzF9jk0AjQsgBXGtKF2d/7Q==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
d4iw9XjLxs3tzt4sbhZGWVOPOAvUQSJSSppf2pQvtv0TNjMCYan8wxkxMkkj
t2j9StD0a3mwEg1C1Rrs2FYwd7wNZ6g2xzeZ0YudmbjMVC2OZ7G8hsbrExTQ
TTLtXEWc0cSo9/FlDnRO6Mg60saja7fZI+ZvMcKpgS0FZEcnHI5+sgx4Oqav
y0CVHgUNz5FonlVMvmH34FTV7hhK6BGn9RDZ8RPPwtGSt8Rcc4NECgMasMJL
zcnVsUaPKowLNruqzmB1EAvMoAiIuBDzSw9JWDuK7hYKYxuY0yai8SYfOZ27
kIM4mcNS72kjNPJh/71ap/VutO6Eqe59kXfBP2RDJg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
XYN3QRe8/bEw4P4H21l0+R3YLJqSuULMcsB3ObDMmzoJ95HLTQ295cyXvluN
viNN11EYlQBLjYh+SWPAEc0XYk0Pbx0AXOUzJL6505s4W1TrY0YSZ8llurXS
jF45kBF5IESbt0vEWI6tvbQHvMOaXgYb2dhzmZVfNZaaCG52ESM=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Jg4y5r/ml4az8GPksqpNIn+P3feCL1HK4rZJwSR7GY6RBjtA6/pqqOpDES2P
IqklwikQsszygcEDlhQ7cF2Xo0trNMInW5zRgt+JkIzkDpINbujQr2zn48eJ
r8JIopvT1QNYNu0Xhc5y8jkUpoWSzslSRuhI2QuhKTE/05DW8Q6c5YJz0smA
ZwzWpyVA8LApIit3KvZwPrj3JYgk93vLq6MvXP/gyfyaqsJOu9erErnRe81+
KTIRxWsdT/0ld49QeR3wYnNB9a/KOi7inJdIpz94zANKNAs1FRj7XMF8OETA
FnHgey8ykP/uUd9oCnaDEnr7os2G7kxH8L76JWasONixN6d07o5r7OlsEVws
5nCVbyu8m3w+OnAP5kZjOK8qUXvc32eOGCBXtRviHS3tDokwFyNE67C1iE6c
ANeBHun5yFHx0qb3CoRuJdnyagr0cUNd+OounrrEJr+YxqBw/2di9Ig+2GZn
uf9NiBG/lFwkUUqG3tKa/tgH0SNZuI/8


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
pklIuopqHVBFqM3fTq0yn3cuvldEshImfLjDxPOxRoaopMtAQJs0pd2qjUVk
EaYzKq46iN6Vu5y9GJEMCV7V23fvF5YFzFk3AYGNrdN5HIxoQtjdkkBoDMLP
oPpXKgj7l1NCePicdNFypjMdVnguIU708QiP5z0ikPREazrMwAU=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
p/mMHknVaPQ5UA41wf9nitUoD79g4rmxlqewkipLzgdQa2eCvDhSkNVQARfC
G1yZ5WIkNJ/e+b6Z6gkRFT5TJHVHGFEsCpkZi/FtYw9HltNNzj/NiHKucoph
dGx5r5NdE7MFNBpULAIHLXLSJwGBlYyhqlM0sXfYpqCGVT/Zpdg=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 10656)
`pragma protect data_block
Zr8NZH5DGSvy1jSia5SZIsZsN8b0iHHl99pGdmjVgZpTntZEbTKxTGTZKU9/
lRrE+5imv4r5nWRCtOMjv2CT3tM+r+NidNxCEFyBfs0/onspUKE9WgHnEKQS
yxL385ovS0k+3BidKvp+CKAxXhJpUGNA463w0FiJToKH2QykL3Y0ZepSUrHF
LKbMHKaXm7PuxRiba4Mpr8cqWbj2VwBHjTglcNhVL/iBqcoBcMa1aU4+A3D3
GGOhccuY77vMvFM3gVwX3mFsunLAEtZnDMILmgV6PMn+cEwJan5e7qPrOexx
o0cgo8StuzkuP4pDTyWLK83+zp1QA5TUh8k0CQYhBWxm4wez1L6iHOiBrUON
KXVpsR3jsqlsL0xIHa51fPQx3aYqYG7JlByJiokr9y0lPjBVPDHjDT17zjxD
34nlpNpjpcYS6IjB2NRlC6jsiwpAvAhJN6rGuS1L+Lz28MoC2/QNuZcMJLRH
AdcZ3514mHHcLPEAJO4wx4o2vyGq7pqHZtn6AWihWaLSvJuo+e7N9eo835VH
H48Ci+Tv6g9A7FtExnLmE3BR7LAarY0vThJmshZW/zP7fOmrrrZ7s9Yml2Ox
3vFj9C3MhgfpWwRZT1EqEDJdgzHaz2aVFx/ORO2IEOthXNBt8d83EQTBY4Y2
NFwtf3wnSH7kNuBTXuv1sCqlcVmqaaGBzRWvSVUe+DK7H89UFI+RCZkxT2/f
T7EZllyY915zHAVbLozoGLbfCqW/VN30UxyiSwcWXHxl9rrpDEdTWg9dJdKD
jDtOjVpM+UlYMEsmCo7/ghl+kWsdfRsefY1c+LIyZnhRpeY+3OIhzsL1Mba9
m818myJaENLEZUrnXKTfQNKD35Ze5ZoXaxTg7/+rKSBX/qljf+EpKUcBfnYU
oCY2+C4d6qqEabeJwUJGqPpxJe9V3cKS98TgeaX7uu69zPE1CmimsitL/WID
TR6oKiWkiT2qiUaBprcuaPlKa99JemgK08rcijhomlsrPzwfx2js8xaMv4dj
QR7M3UMldc+rvtG1gBky6IUUgEwXS04uGLpbSRvNOjN7LUfadp+rzZEhnqCh
0xuWcr75QcG23u557h/vDLvtduLfSBEKTYnBQzyXWAH2KQEBHP+aYrkP/PxT
OaqZaMMVsFlxoL78Fc5vfkpa9wFbYPXZnhBUAXoqBrQNoRV/iz24l+v9SeOZ
i1sBwFs4U6n7en1gDdf/ocV36k0zWGsz8IXyMh8/1j8gz6ymzDlXQfzChvYu
vEXkZ03AZZbWRJfPLbS8OTCY8bxOREQfiPVNOs9wIOc44LKp52EXqOhnQVD5
2DAwRvxjAVxw6rIFjMO0pwroja9TXApjmTJtn41v15ldQ3waP9NYR2lx5zNy
OLrKJUKPiCTxpTGsQKq5o5B9RolDxm8trioEjvXfUDlMZxUa2w5HK1dWxvMd
elfXjgDPdFuvahTLBVZjWdX+FjHBmXeDJ0fXoEDtodu7twZHkbmKb/Y7dWks
k1d+4eEdcwubPkLdlyeFx1R0XKH1bA24A8LMBcmdWUi19Ge/L6yrcCbs6K2e
SuLre6P5TtFvPx8sF9lYxO5dqGUsoLLnmgadcp7iMg8Ptfnprvr2aihuHxDu
hNbyMjv6gD0Isca/1IrvxqrOImnSSdmq2az9/C7NbgZc182E1h87PspjDtt7
JO5/4LQpzsFQ/2PibyP93xaJnBDGpwcgOd/iVbKQ9qGMOkLFkUKZR0ln44GW
IFD8RRhYBKxvTeF8uAdQ5vcyKLIvmWyzB2qoDMPZbRCy5fbG1B7PKFFAsMT/
YtczFkft87EDutH3B3mJTfq+Edfje+XAeZcZm36/omAto/IQ7n3QgwkuA6oc
QA0Bo0FJ55uNYjSa4y0oyr6NN13oZmi0lfj5rZ1mS3PADpQu8odRmP7IZK1q
PTJT1pM+3FfncejMu4jP9234oilGzI8nv3uoIGBuXabg5Ry3wJx7K5BVcAxb
W64yN/3jPVGzaAMMaA93ZMCnxD+Bz79ct+jSSQtFaQI6o369J2yZczqvxf5e
52dVr7g5aYGdg9Ap5dsZlpuQrMWfgnaZ8Q8C9D0QEAhQiuCKPqj73HVsMDOZ
Y+yZxf4BXzrzBQkmPxxSGYf/Oq3ypD/21hJ4dglGrhzJ+M3W2Wq0cIg5ARRL
PGlV4dOesl9AOjH0NFSDtg7zmcRuX2Ttl0GdcMSImvcviEPdY3gW7ViRS/Is
W5cEq67ZEshsIRpwizP4E5ffDTjcbDZhvSuTe4fNbq9nCic3g2rAElR8Sk5i
4iV3rG55V1KAXhd8EULN8OdNSXi7YAp/6KAejZImy4kGxzb4p+qZ43EB78vF
rkbCqwE/0qFsXA6S6MLnEvvskAD4dk/urc0xrgAAHdZkqXhEY7QfDlwfNc9h
oXlff9g389DDHaHINw7R3Cmzd7bk4EqUhR+vqRyqVaCc0rwDxlcDFeWGqoR5
qYSf/XM8eg/XZuldeQNZKU46cFJTIZXZC3QmYH5PyH+iiTCCvOarTGOZyUl0
ZXSV9iA49hrdpSTUS+Q/XVC+sAPreQqte68f8knXOPrMp5Qzv+Qjmw2AP3eh
N/p2Y8teFQIEQ675IPAf6NhS5LcfrCIwS5dZkDjNFr3zzakokzGhZ0eLn7Sk
Yho3+VC3VtHPVOBzm/PsifcRFrB1QfJmYs3vMogHoeXIZlTraR6D9EPyxvm0
ewszkPf9Hm5gNJpQRtCq3bKqbTYEIk4irOo97qPXjUGnQwsiAALGDAZJo0Rt
M8BugL4+qbRa+ST8tqK5drE8VGoF0qOfYksAylDELN3ic6WWWbHPYNKW20kt
XCC9rC+5A9oSRK/vbzGL90oEMCv75DJcvM+HKdVwm88/hve1HeV9FESZL8wa
X5zQBiun+cZ92nz27JXhBoWF77j4bsYikiB6x0oH0xqDFDU2Pajz/CPIx8bQ
plQzFyGMtcLu3oe2yyMrwHqZ4d0U+npqphXZfo7cHER2TNDeD8gTSR4kvAoF
RamE5wKALdNbNk+ENfCc8azzfq/wqZj9UTj67/lcHAR23TvwfOrqjpJ7YOBo
go4M5ixTjlSbZEfxo+gSgpd/7/69SavdNcMhxxbUNLyoq9RYNDBoIxXR1zZp
eO2Emq0qMCZB3Wxo909D+oGRPoYgu6Sb1VPbEoa8CFss3jY+3GivjCuJVxLp
59LZ44vTGckEfgdypoEdkZFoDdS46t45a0h0pjz4GImBykAz4uPmm5u8KEjh
wCh2q+SUNMbtdVG8+yLfBC/PTwziE+jSQMnEBO0CU1S33f0T0kIrt5ts2DlC
SvQB0ena8wc2gAEROdkaGhg2CVJs39kXpxLExFbkSN/VUknkd5u6Js6gdxk9
t+qW21QMuFYL4jLMCD8Xm/CrKyAyE/V/+hk1oyX7YrlT0GS5yUE/PK/mxdNf
CXGcpxZw0M9WyOR5l1nyHzYfvGHt7E2dVv7E7DpAm4bD4xEjLh3y5SPMsIVw
XV/5X5p9hltIH85DjcBiW6vVfA0s6whrqSBzogbwn00H2S+KeT1eDGLalggx
YFSucRiK/HTLGR0SCoT8fmGabT09fOgnsBXyhD6IdOp9PyILbtrmSelmbVhp
45rkjLHQ2HM+0VNBeCSIcCn22GBYO0uD2yRtwmOwcG5huJxe/KhEZpeRb0FU
Zsnj3iAEKyC+Peh2dliUmAPQTEKs1fJyQrGg0sqXzvhLIj7958zGL4OAiOmN
WthdBCIPNmZ/fhLfjUseC+0MzF6Elxt8/2VHS90+t2svw7V/km+wA/p1HReg
j7EQP9bufnUx8yLI67Ff9eg9yz4GjXMhtIBoaHh0x86TLczhKDdOpBFQHL1c
OmU1ZCHVbk720gEaRWsayjwhpSTELYxixhC9f3+VIzOgZMC9C2uisPrOcqtK
QURKkqAbmY2IH7SN+OU1uwl8oetHNp1xWnYGUKWdaPacyQBYYBHoH9CuByxl
Ai4Qy/T7136ryaU9fRiYLFLl89707lJsbSbyzSDVPL8vLeX/rjDsWIBMC1v8
2Gzm18iK1BN3NHfvnngoyRX+dczI5WKOBCbet8kgjHKCwHlCuMAQvUg4FRJ4
e21fpty3K2ytGauiKK4FwBOLn+5NlvVD+1YOfR/PVNOxHJURSY95vngi4Dba
/aBadwXpjbj4ivEeeq3us6goWxfwx5QDicwyzcBKu8iSFqgSHMIbWekqF68H
RUOm9V3sDV5M5bZ7kUR6HUus3Iq0zIf0nmOuDaLC7BX68M1DT86oq/3vf91G
h26Z+q8n05d1rOtmVugXCJkEcVmh0eXqKpTzrQ0LM08YyDsPqvKDwsMAE3kM
yPxmHE4FTXSIotPsxLM2OaZW45sqFd1eBBeFiuNYtUitq+DLDkn+LNeNnWwb
NyBrqyJ/TxcGPGIDolVhOFK3+gcTlrzhju+FVBsMgpyZj/Bpm6WWNIjOnzFL
dhn/FxB28aoejZ8Z311O4AF37oYVJGvMeeHSDbguknXyQyu89pdJ2ahMcP8o
7tGafMPU3d7WjwkPMmFuK13rv/vp+tzc7zDrJLBdZhQ2abyRpqjjHlMfS55u
dSH85iqLFFxYRQEIINdRtVpaIOwUdlRzSirlH0yB8X5V1/D1lIDwXa47y9G/
WkIj4Gz8Re2TAT1AhXhF7kBJ88wD1ioZTpslWUpMlWWe0HFdis1iOpKfN2yo
/ya8i7Z2FP9sKs7ZUSnF6WVdOPJCe+J6I0w4I5p0Ot7oVUbgrDEWDaLlmlfC
nS9tZ3RthKiJETpTtVEujHocYxBdtHv18qR6BH/90SoI5fM+SSFrELFBu1cN
VC47xXkCy0/DcujzYPcNai1M7sA5UKJbDDukPFf9PmX5V9x9oZVAq7LEUX3U
jd7n53lqmJC4Pqz2IP+znAs3ijSdvovLKDlDZM+8I5owWDzMZMa7a4tt/9jW
exZrjH5SIK7WLQ6E6BOVXGnSWBBSVj7/o/Ia827s/I8xF/sdiGor0A1vHOMN
bFQMD4Wxd0N0oBZVMwwG/RrBdPXscrcfAYIIkDyTT31+Z0uDxnhMwrbOAf+8
qcI9fzAXvfs4MS/5Eol4BaXOKidyuUzJrfFRqY3oYK6CpMosB0SB/ypicxjK
hIAr3cbRaNfzD3VQTEbNfHL1g/jQ2oTTxY3S1sB5fNYKu3x+74mON3DyLdrf
U6mexwzQ4mD/Cn1wnuHqGDJU+OAACUWj5Pt+SWf45Aq2el+ZCSAbqPqG5kCg
V7k2sGexh0XXIRt3tKDpHvqhXo+nKmMIFUVtn8LUlDq3eMiWKFSxnbiykguo
GobEWxVstzlsaTWYFA2p0z5XAnG5Olr0SKVo7JC8UxQ63qaKuqz3zCFixqEE
CoHNb1pyFuenegNghmTbjAkicD93YZIAHg/hF19UHjL1YxcOCrw3+b1o0oGq
dvtZU7mTLYxqKBIaNuXgsE4WLOiIu1Ekn1fzHlqmGXgY5VDQhU+9m6iz59BI
djEwH48JtD+ekAe1eEcxA7IsF9ZFsfSsXEF20O+bN7UaSibCcvOL9XQUTZmz
PJ0oBrWKLeSBw9TrJs4YdVMT1qPssoiu3Dw2LtgQUNo6gBrbuQs54wsVPdWW
wNtKun1JTALKdFsVbWsac0AOYzC927L0ql9nDt76r6WCy1CYQgbcC0AIONG8
jKJrb9wkWlJPc1ijxkfNa0mwdvkNpYepm3BiVWmwPARk/CXMBnvvoRk6EokH
3Hl5V7ih2QQdvenKJwgEn7wYHyjAUYJLZ6BaRChnEUMsjFQxpCcESI3+i7Eu
aPVFikTNhX2T4M+sK2C50UiETJQ2C/XDz+zc41P6kELBbvjUwLIzg1Zq9wKM
Szd8KMNJrLPtFoq4OIkw7VSI2ovTj9MmHVm53BFtoVGygacZMji/GPePO++Z
tZq5zfDSCfUxSK618Wo0tNvfejoOHP92e6cBaQ0PwJdDFWA4yGAYs3yHk0S7
GXJbX1IjoVmVaYNSfNAcnKS+GAQw3wtrPc67GcbohRErqiyupSw4IakzFhS2
C/hkJeYui1ohxLkTw1Hdhoz2VZNef5CaHOpZ9YfUKkWTmmJ3EUZRtDSFbjcR
K6nPCq/ftrLQUIuihSUvTyAov8qTHyNMnHillH9Fnb+gH5nxn9x1hi+8pR0Y
tZOeMHWYnLwerZpcAswlD6SsTwBabR72uQBUbfQQv/95fdXNEWL5JQ3F8Zyj
6dH/bLIXXDRslK/vAhBFO/UYElpYn/+9jzL0x72hmlVYqkVEkZb11X0Ho9oL
Y6DJMzHD2/0wmaYZhRCJV/Hqyfu5MYROpOgvaHfhTkX8JTgK/Ws47kNvyHck
FdfHSF6XUEqq50tZdqaFn3sU7O1h5PJOmrb0PJWozPYqOC/wtBz91BRTFWai
t5Vg/yrI30JVALuUGAqXJgmj72993ojLUEo/QYn5WZzOvjiI7HO6mZOwLgVa
1M447eKKOM+FVnagAn81OtvXKwTeAyub7kDs+9OtrDJoZgHUYrbJlIuQxruM
Kxtm9UHIO3vHjASilUsakqSu+UCvGtVCd0Fg++/g/JaVo1ja5TzDr8vPk+Bg
IMDmVdARhCGersdjlsvsoNgDovswP7j82wcewBr/iPgOIk86VreLKqnCJQiR
VbWke+VGrWPZPpSX7D734r+Y3mFtosChtyLfmWnnY/OwY4ObX8EwNEhl/2cG
HbyTN2JF/xwduxIjf/u858iWSISktWsPmW2kj30smRkC2IviRHwKs5Nq5QBr
4shrOfJFmV/311sQJetndQ3iNil+6ig3keF4CVBngafbsts/Khkt9IGiio54
FzC1NBkLtiRduOBz7v+0nvS7r7sjuuIlioUz2XxxKphxuMF/+JzPdtcJZNAX
seWcsZbyJlmYSMZj+bEaDD3yBcF9y1HsudgoWeYEOogfEkQPQutEpbqRbKnI
DYAfbVY1UcUbjliS9EtPh1dNt7nq+7RXiwuy+xS1BCxfLIgsdZgrSRnCk0Vo
sI8uOGd4l6Io9xJuHP94lRbwYo5Dd0NjGXviIKatjJd/3zv+H/9ldrFT+faI
GBWdTv4G807dIi2+/RTeyflBT4LFDkMrUPAh4ih/IHKyMXV2/YbnGbfb8x/v
SFDwCgleiDGgrwqVPMQQCi+ZaoZ8eXpK4sD0bZBXmg0KdKhYQFlxhKnigB8E
ztcISoramlje/MudgM7ubuMWUPxvGCQbP+FnW3lfWFI0yn+bV/V3TPyiJegz
k8D5XpRYNgUzEY3bpbA9N5+34xId7iUa4cUzq5b2s1PcRDKWKzoMR2Ym5vPf
tuSEeHHabG+9QCatq5lW5BUHMiKKBXbIfUS5oR+sGT5Vowgl5V+iPSSCQWUz
KQKjhdOlhCD7OXd3i7OV9zvh+6YWYS4draU3y9e7cLlY7gPiZko3ThSM9MP6
wugTGKvozOGWFA9xTfTbswyR9rWmM0pXa/br7xfpkakSj0HZhprnszQYlzyo
+cS4x8KIo2XLCboCyAS7O+eq0QpYUysqL8MjRvZ+J2NnyL+qJS+ODonlug6Q
2Ww9UTNk9Ssb3RTZuX4qLKL0Iyt4fpCevIZm1z0QR/eomSL4+oixkRda3IxG
4/ndsWLjlUu3fFoJBiZq1FfWD2KJLXRDPXZoyiMuv5u3Uufuy+hvNCFoVWuL
wvYJM6Kgq5oKObfnFCijFpgs5pdfHFg7A1RvnTXmoUQJEJSEmJ7fU46yo0rB
drOEyUwNf9Duu9LSMOUMzwvxMZxBeDSwutuRUIJCbIqSPXm0rUEg9RXC3jaK
96Ym2hdCRGHa83NNtWW3pKnt0ugL5wQ28s6eC5gizj3zRBgGO0bMof2X0E1S
v9YXvPYC1Mg1aEQNnvIhxKMYDLG8uCWO6cwHjc0DeYfXseFYDc+GHn4uuSfP
FPFg6HupOoQykKKBPjfceXJILMeZbYLNPXz89ZCiZMbRPfc1u4bSvyztDrcX
MTGOp6HwlQVGQRCEqxD+PbkchKeHM85wQKoGWMCwgsUF2SYTnTUugLhON5tE
UxH2hoP+5RjxvC8kErs43GsIY69cdfDSog8B9aY0JeEHHnyY24mTLO5rEzrJ
R05tQBTPqi8a5dqm9dZyLOw2Uc0rTjxYBZk0s48hXucLcRnyUQq4uFtfZS6n
HnjxeVb20trshlkX2Au8M5qybuvW1Z1ggIj1zII6h34AQdisR6Ul6BVAhOY0
zRrxXaw61cJlqRy90VYrmHZGwKPv+0KWGyzmT3U7EPSygqDbNJ/1U0PInevX
B2wBW5j3bg1X+LFuvfeJOlhBjbQy23Ye9lEaAcL+ySF0q8m+s/8S+Zclmr2F
2VrsZg29NWcUug+72M1w9v3zC+ip5nwNAO1ZeEp4K8t26V6Rx5X7g4sCD+R9
Z5/09y6McBLhP7EHeMiHgKS2Y0Eid85e4jqO3PUdytzY031p+X2Yl3vL2T2v
R4357b2F1D1sq4JZAv/5cZV5+l3R4PEUifkc4pJvu7QZy47fLWabO384p5tO
Jqup5XtlUI6TgCmT6RAO9bRLMSTGyxs/vGVUH4EVlXds36BTo5a6a8B6PdZR
ag7ZLf7QtIXdN48ztAPP4WCCoJFSHn1489DaPH61m/HYeTJAkoJRDiYklyac
xeikarg6Kwv1KDUX/sLw3FOVteOHinxu5qaBFRFbhSxJaee+LG/Q4j7hrBnf
YHP9amUqqF+we0FdpuZZTHy8xystGJXKjE9EXN+oBGttTKlMQ23L5/bleapv
Fiu8nqqm6PVmqdSkRS1jhkRh9s3c9xP13V/bcp3iSnmQsK7B1ye7P8ul9H3y
IJGpo+OQ9D1rd4bpdM1/8dWe57BucMiykKHBBmf1cnqxTiCM/q+xO+HCd4Qn
MJ+m5Tp8D3rlZ1W5SVgDEooNh2aKhiGtmjnpbplrLF35C8eWViI9KCXLs14I
RP0CuNnpjNr0yGGYxxbDkThHphct69HsOIi7B1ueCNuBaohS6Ht2qoXM7XtY
aADFoYfcDmkmrp2GAJfVS+VMjAQhDp0bma8ZdnkPLDMonkDs1i6B6qNUd+Ww
RDlCmIumcMTU0uUwU3Art/rrRsgfWINLrB3Evqc1vXhiduZfBSdROye2P65X
s6+iU9ZMJlAuXqPkHVKLgmDdiePug9iNDr58b70rQ5Gv5EIU42QX5sp3s3Kx
+Ew9IRv/cL1zpDSyLhj7LNOk73GzvH2wSQlv6GyKE4uh+EKOPhX8dv0Lai6b
txH3F+KRsTnJ9r5QY9Zfm1E6Pi1Ul6ugVUvK3OAktGAofyxu2rb2FoWiVcPN
iQTgG6ubZqM4wAxxUc+i/r+pvyt/lh2jhgjXg96FrlhxCRW1cWeit7AGv183
pQGIpzRMq5DzUPK2iGRD9bQVb5DAIOIjI8jejnIxOQ61xH3OhyL3YQBGeicq
9oJMg/EcbobBXazel2EU/X77j3HCKhGUpmG6juPVypS2gKyxSh3p1iqSS7y+
8xJqE+4/xL0Z/L4R3jyI89AwhydA367453D4SgbBVVj9qSoDYDjCE7gcRXzA
loYMm1PFjQAwsXyUX6s3ZI7ElZEmdt+je0iIXQX5uZv274gbwt+Kxal7HJXS
nofBtqGYVp+lUWVIpTI76enPmwowXG48QTS0Xo9D/lUAgKx7qHeRdRWMWf8Y
oSjwigbcX3/HZEh0NDPo37pyoFBO9x5A+0zOEAZicoYaiZuQ6eY6BC8CZOH+
OBjKnfvhclgqTqSQ59/uK2yPn1FsfuL+ONQQQEzDHmoCeYCPd0iCe534Ujq2
jco1RTPyqhoCnSMfonuxzBWvSczx0Ue/R/KkwpzuhSWf4utVmZbkmGnSdpYD
213bkK+BRNYD7NfzSRbLQqv5y+VEGeq3DV2vJDMyarvPQpprI+xlzAxOMG/7
IgQlekT/8f6ISOcfX4gumgbAn3cv3xM/SMgtF8PyvBC22l5XaJDAmiLJorrW
DFZ6kDrMtgRR6xYI492fcyl8ma+lPmUnaPOfEI5wP9WpQpG+oqCzyyOhJbi1
8eCK8gXAz9cNO7kWWEtRUogerMu6yoM70oU/7x1NnIXVEjD9zAbkDpxEJ7IS
m4JQcZL4DuiPo55yZgIJT3A7pvdkfMYOTTw7yKgnqdenHk7P3XpibNVtOTYI
6ZkhFn274Rhe+dDtaeyxDvXOo0hbGR3OchuxOSA+kneOeAktmY48XFl+6+X+
KL3aFioBTN7V9LLFuazVh8E3TgEdIqUtd1hY6QCtuZeDEnPkDlDNbDHS4W/X
USgDumkZfnBTWXamaXW+mRo/EysRgjH2BDjE8k5yBwAABl6qsjP3Sjb9BMD3
NpSvtKMrJmjvvwRFwgOoTeXT+WDebx/LkHRXmkw6tfIevDGSixloEzRMS5Cs
heNLmXaZ7IzlX6J95fLwEJxMVyX5X7o+BCmT0kP314zBAhLrnBOTv3zzoxGY
pUPi78aUA+0T67yeVUdrjl4ry5AWw/VrppbVIDO6Je+01lY1xaZq6pW32k8/
P6NJ05aqkczx3PLiGbz5O33bZvgdCwirYFjxfk8e5zqhO+mz8fIBWk4pP18N
b6ro4Cwngh0EmpAg1lhqezhys/C//dMILfXUw0RXyn3efeY0OQhPHI7H7omK
P2RwRGcyn4TCmf9IOhdCJeOGCI9N+FBeTDN6pBy9jPmPnX6+IL+S3D5bL/xE
V8UXVG1SIPhSOMTkrOanZYukVleHsSJV9M/XjKbaNo8vtLSxv7L+6klUQYaH
IvaNozjp2o6+OwGBV7RfqDL1uqEpVz4BCUiuWvtb5tgiDA5Jxr+L48bfcTw0
+70f7BtC+l9BmO3HroLijuHmAVYrSnSoEjeShDdDIzLNv041WVGNeooa7wac
QpMvqsM95e/92G3lnxOctqMn7hAawBkch3pSXoOO2Wjc4ZPXDlP3HaKhaHvj
n4y2f/nxHViu69oDGpBa5ZHBka4R4BrOKXKzcua0tWvY2AGMeg+0LGrr0zfC
zdpIPnOV+deAcFOjQ9rClmca+qw5NNiO0Rk+MZt+elM2208TqMv4daf26icO
lsT7pUsis0HOA6lYyqv9rm7O2VLQl4lG2ryFrwhgixm0Q6B/qx6XBKnfgBvD
vv7TuliWLGu5Hh0Fx/z+OY2DHcB/y6AcTrH2/VxRS78cq0lYjzX8mGKS5lSC
fxVMQPQaxRuA7w8WGzAsOQUbNKc5/kKYt/hkzABgndwC39RA06iCatDavNRJ
Wb0qDZE38ZyVObuRaWOtSw31NbSknZvtzswx6m5QnM5+iOiP2E+cWdbT1lS9
sRyeuloMhyFG9rpb74qDIlOMiPyzEDrp1KGd87ab3o9JThppaONJKniIujEn
tYKYR/Ju7TG4rYgjSTtvOTrUL0i1YyAcocWQNlCNOSoM8hC+12AzUgYJuFGj
GGmGWU5fsMSehJtxY7BuhGxd0H9oB7Qk3c4n6IGRAgkw9NxSC6ECIUVwxABa
SvePEi7HBd/3IMP0cHQMZjaoRvWBqLNUNZSkMk/4lzqGr58h6pgRrQ5yYmt6
x8QxTdBiVt2qI0GAqD8NNvDjfTMZtszZ//di9LNvf1uHo15R769xIRRy9Hmx
FxBr1VrqfFeFpwonfV4CN6EZrAnGDCSKXWp6sLiKo5zqTMb+J4lnp109+eBY
UsiWb/Kz44X7wApi+ijGHd4b4sIiJOClVZOMAhohPIJSAgi0GZqFfDbvTMa7
ezLC7SyGsWLwHbcCgdjBnbaF/nRcRBuYL3kcPNkI9u1qYOZivseKUXIGmYaz
HE/ncamZdoQyUKJE3KC9OSns6VXBG9lzOkYooSiZpX92lUU0xB5IE7KnRh+C
vYUGrr2aDh7xG6vPFcu/xGqwe5Lx3aoyr7QwgiLU8FVRC+tARZ9I8Vmh6C7H
kMu45ue5F3diDe+B/hXcWOnKH0rcDNKU6IJug5/OFLKIOIBexxiX57sNOu9J
RIYu9Ku6nDpHcBUI0wB/s2KRz13LrLUiPIhgwbPZuEkSfygRpRZ2QGQQcpSg
+82HHyKg2bx+q2GLd/xA2fpODRDa47qOX7G6PRp2aVjbENSb0fGvc8Erel+0
x8CVbEOVO18HwhFLnG/1hXhk3TeyAIW/mbb+Xn8ITGwfa574HnlWiig59Vj8
MRtlGvze3LKUmukJyC9q8dEHZhci5G0uXE61EBLn3xWRn1RkQ0xkQZNgm4zK
kxjMyl574a45C6IboorGAaOAEJGN5fxghS5aUIwCLEQ1e/knWRLzZipRGTVo
d2BS4w/OeW36Z7OgjDlnHMoraHf7WU7qqjo/Fhu/WsxsbeK2CilGo/SLQIt1
5+fJy+KKWgfMB1RxQhXR3UaCtmRhPbiwTqDJHVNPUCktUQ9yr+6K841FlaOI
8vvMKEDz+fg/LNneyN2RJYeECeYs75NnjCFZPrJQCXc00usNe+FD5JXCONTT
Im8k693Pfnb6IUclNt3n9uduZ3L3LSZnWyFC8guoJlC2TJ2omwUWg2HIUWUP
8OKX4aY5s/kW+ZqcVxfp1bxhKPW6j27lLdH/LtSD6FaUMvHNvcWn26hHlhiJ
j9CCJSjTPKV8aZscImioLE+aPQSKsTzdNarImkaSRq/v12fZokEIfbPmiwJ0
sYYR7ojWBbMsp4zftImhGyhzt4sP7kgSn3+PaDUsJEB1vIw9YlX31LUIe6bV
XINDFtjFBodFs6R49H4lEpBDYXre7YUkxfdM6HOJJytoGpnnbXTArXG1L874
rhhnWEPP029SnCA1ga4llAcxXXyhoGwmPgde9kBQiM5kQWBWoocyiLshf+Ah
GWqjIIklDNux4/zFb0Vdh0aAc3Ixd7hzGWdLnzYXscyT9w0DaXedRxdaeJ0Z
rMmAeyARSOXj1UMhKgyH4+XJENXBfhDsEhjXDPJW9nfyAh5pJgFr8LgfV8fL
ewsm6egNw7ygbqbGyKrMb/L/hwaBOCmZVaxgq+WRUBjCYYPkj/Y9MUzR+j86
fPxrkLdII3XMvcFDtnPDlwIuujRQZVD2hP9WfNpYaHy4bXM0MeSHk78JY0FQ
L68mk9ksN+az/y8K0PoGzI4xTVyHriTFk+oH+w+krTvIh9GPA7RDlpef24yT
30zx+Ao/aBwPDw56+IgjlkkhF7F+eENDmPh9dYNLstKOd2D2ki1iP21DaSN4
WAgQcyasiO3sHUxOLOk/FoHvKonT8pv1StcoIqraabED/JsaPFQ4CSeto0VJ
S6W/XJNZEjj497fe+Yxx2Rhv53/sw1qZR5Co5eA+1xmI/3nk7G9iSlwNoDv/
ThpNtc5o+i5ADuVFrj5LkTP6m4tUwel5Pts5wi/3fXrOGGpoVQiMgXx+8PCO
vflGXIAGAQ4c7tt+H4xDmw6i2jHDMIGUThVdaB+cboULS/4+fOddk9IQU++y
WaZHIeWYtTTvvCokLPBTJorfeVL553QaZGSLBKZ2we03a3VuJrqrn6ElOaUQ
JfmdFUBAUqeP4g6LdkJZvwZrUMajX2xOINDNRxCyzQyT3qcCyfSWw9dhvhFo
NP4x+jBc0qvxA9V4PXheH4qz+BmBbtXKSrzCHi6U3idTcQGxLX/UtXkP4XzQ
BDz7APrLYKYFup8tiKqnFZLDcMDTSy9ZGk2L1do3yjKsEJ7vRtz/MoLWbzBR
SbUIrESvoyB3QflbLNAsWUSPmyUROSb3HLqLRKhs4tHb1CYyIbkEXBiTpCwH
NpSXTT8YCi4hIyMY6/oOUvoTOYRTiS7aBua4luBCuQjOm3n7uDAJjcWgCNvL
ZmdcTJqMUOqOneAmqnpPoVNtvfgQbpQv1SsEM0nmsqW6FK9qDoOJzyo9qJAX
gPnm3stx8nVT2u6LN4jQongP4mYC/M+ysEEQtjkjm9KPltVn5euzozatActr
tkan3nNMBvOvlRpAsK0t6+wl+Ag+nxr3FuL0bAME07+No1QO9WpoXatDHyuf
0m/bIX/NbE0JUCVAd3INovIXDQQjb4dgScz2uo1vW05iH5K2VbPd7JbL7vDV
8g0rLm85jdOXx8R+AJc0D0v8Clfx4/WX42OFmiEUPP7XBdWl3WaRySJ8ljDS
/Wd4y7TzHc1JUzHICJgYBS1Ne6ce10YWrP9ZCMv7PfVfGREJvLGmVVxO1dWu
eSq22La2XMTAungDUz76DQA6gk/3SGnTH+q+wJngZvtwIWLOqvEQ6Hd+HGON
BOF1T+LN9CAHQHp6NLZiEB3cn8LZRobBzqI30SO5h3Cr4mn3igQ95pxd1EBe
bUKX5+RBYsFG9k4fQn0xizO/LMFbTZWWeZeWQGKcsK0+uXJC

`pragma protect end_protected
