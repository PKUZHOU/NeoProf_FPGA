// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ovCaYQ8JaQKyP9dKNV3eQkZv6+boc5bBfcTwchVN/Z+nLd7CBrVKmS8YI4Wy
cz2K3LA4zVT+vr+SoeUlfm+EQ30aR/RX2hgrTixBaYK5612mQ2r0N35McTe/
eOyr0jVKIfXFEcig19X3BOY1KSbSzZAztwzW+Buf/GQi3WOfBNQ2jkNEes8u
r5AgwQDcSUhM7MTU4vtEwG2By5K32GWQaVRDxrVdLUXo3644ERBvSLVmnabT
mCZ8R9tXy4bKxPPhIDI3rqqrENqHaWbWLfxrwYrXZPeI6QLrEvy9hR6Lbezx
FP8ESYqvMFNcZjOF2Kzed7tjS1+450wheCtPRWIsVQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
cLJnbbfgxPSZ/6Xetw81Jo3IC0QpIaLe+FfNFnTf6jo9CYyL4tSIc7zRAH8Y
7hsDZX/8I0l4xT1pa1Ujbprkj3+gLz3tii0sDkkwI/o4slDBC6EpV/cOutoO
FkcIAYOc7Szf7DJD1BFnzGmsYysdHLQfrsmbL6AxdY5/FeIO15gfzcttw/v+
0ZQhQk6nj7mCJIIQv3eZ8est5pw6LauRRN66feVlTtkZkAXXG+fZ2jwFanf2
pKZ8ojV4aC9FHVN+5Y6VtQNNOqmjCa4A/Peb4u4ift5PPSCjbgA7Nm9Q2SGf
KXze6ku41X69DV28GIO0yeB+IZV0+wemJ1PfIRa9XA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
rUq0MD9z6GGWSvbRjXMFNZh9aEAN15VV/w1JUYuUUOnzQHOJPWaP2Lp1KYIV
PfJKB2Oqzr38K39wtd7Thi9vtIFrB97QVx6m6W0bZc5mSGVbmFxojxt5vDFM
CXU1GIOu1GAtIbnv7ky8xMwS0KJqGHMVf/fs0DAE14HybXRtMkUH9ICa774v
CTFu0E88wAGllT4YZbnvl6T86BTNi9xZjpw+b2gEUhDMicftDGKNinSyDHJU
mnZSYr0XNqTop8GkWXJDevGDYq/JmpTEzNB5FNDP3Eco+vgcm9Ns2rzfEiay
3h/4QJgb/Z9Jo7tQLyzQx6YwkiLdubvsq9ogLDSNUA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
MC4k5AQinPZNLoUIgqM3C+pSzaYjwfrRbPccoKp5uH6tWgruWK9bJJte0JoG
/jxMvC4Ui2QzDMFTRDm1U6aNICXtAzR1pMmP8AvA/FairuQ/TYqgryR4dwme
8Nztr2kGMc20KcnoL8J8GF4BvUaWauzDgePVkKzfAlvmK1wCsUs=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
aliFGUlPHcyq1k2yKEXr8XyqlQHfmBDwItQrjt6zqkosRkUzh7E5Y+JpdLO7
bQD19HImB9Dbn+K0/uOsWarpBMwXFVtuLZJcp38SZvRIh35/q475Ynp1xfaR
1yK62UH2IsjrX2mFR+DA8ED+4bjfM/5/HFO6yQT0pyyjUsFChTIgwISNYbk5
LpMTj612xjnMXfN9fJ9s7IHcZWVcncd+QyI263fBzz0T9hBk2o19YJA2mxC9
mcWJefQNDRsn4GSmOL8UUce7IVuPVB4tcZ6bTdkl+djgk3c6b5bgQfaoaFD/
VeecuWsy40V/SOWh7oIKwVEEOdpL4T7b7sjriS4MbR5mBjSm8MMjO58C3J/N
oVsu0F+2cLRD8vd3ofLtbflYIto1846Gw1uj2L6E2ohKKAnTnSMxlZit2XEE
Qt65hD8pw8N3OVvRpr/UmD1kzl0/iITEVIebN9Fj0CXr67OkHqPmrWFNzYca
RmkfnPKlu/QylTds6i0Fdb0XT1XQr8oV


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
cuHIMA7Vs8wpS8mGzW2TQ9o6uUCD7jxEYKvaNjs0ctVecjERxgT/6k5k5bwy
LnAc9WUGvp0zrMQTHtPqbUIPVQyQRxjjW9EnkeIwMPBbt5U2alOvNZu90lpo
NCdpMRyRQYwKfqLn3xO6zKwPdA8LYi23U6Ldq+amws3EFBsk+VU=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ZO0DXefPfrOdZK+1AQorJ+hAEaEBq3ZBnwFxvf/7hgoakLcvq37lk9iMQOAA
6hs21jMzcY7dOw3JeyxLiSvMMx3/30AG180L/NL2nkwwAVSlp5OttO63btMl
sPodc/SeIG93/BX2rK2Jh+t0LocD9m548228o2SIpi3/+yXEn9M=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 48784)
`pragma protect data_block
VYfrGFEh0xa2Z+45NqthSWc3qR+jfD1LE05HmDY8F9cboYPpUk0EErddRcVz
Z5k8TiP8hLJcRoJn495ZDGWUzuLx1ZxDvsO33ML62D9bdOjFIhDbrYxWv54g
hqNBmLXjj45pYq1QDGJz7od1wqo6JeOa3J3GsHQqBZivaefcHqi20dUyH473
MxTlmVQMJnImYWyLmGi/7Tdk1SABYAPvEOBMtUYQBLaZ/eHksGRqCFJCYg7Z
ml5pv7vydzh2/U/W8/LmhfxHe9j4E3tjHOVO6SzuAHjSWlqf8hcY+j2I97wL
3GYxed43W4OSdVVV6i2fL9AMvVAMJkUXrZ9FgS0RMa51Fi3BOZPU87evXB1z
j4h+ohWA4Bmz045kV2Y1iWwojh9/nTCPER+VK2z7vfmwEZFPO5K+0baOa+ra
2nIheBjuSYipB/x0ZZJKLUezgH+wcYNTe9j5db7sSIzDekMjrzUmNdJSWycx
rT/WfsDhRVHA1tszWAPpPydT14extanIzDg/TlSVESCESV1zuuR8R515y77m
0wHC7iEVRkoFN/bH5KZANMLDI4OQDeMuHgMf5Vh9zvvHjzmMOYXV9bbnVsQv
ZAbnFmfTE2FgEAy8nkH9GIoxUuzif6Y57AItiF7eZDj/8dlgvd47iwPgKSQw
cjw2wFoLb7bqlRwk8puk2odZDB3zqz8Sle09DwcSB00dq5pRkoG9aKqu6YRO
cbyKGW6ww7tM0c8L9m26CvrTzru8yB9KMoeAt61sXsUB3Kc/WLH3E2JZHAp5
oSBJHuf8XxCawigw/fR2WMqkcOvjKa5nzAfZmfwImoESD0Pk/X1ggLneEtrL
tjQrmAsNYDPpJ1jm4Vy7WliEswIAtI1MUMY7YKHEwUkNVXlKVrBpGiCRWTmh
AS2TwDH6iiR8gwgCctBxRN1pKmIwK5+YMF1NwVnS604NWrQ7wZk3SILHlFnV
OpxXdCHCp5GsGp4WCbAWNRpLQmuwzjnnlrG7WRR+rixtt53TcUr1MBvxcr/Q
CF8LUMH5rbNeSElg7Kp8aYxLQuuU04U5E0TOB2V6kgkPv1KShvCQmIwH7MjW
v155tSNceinc3Nwbebbu3s4aUys8mt2fUc2gg+McfZoXXGqWfs5RgggiFbU6
qttswtC9+uDveeszCJftznwOcLMW7pb19e/fMhWAazNCw/mXG5e2ZCCpGyjc
6nET2Icly9f+2fqbkJ2WNlh07/pFhEUN+vnKyu1PKea7z8rizAUaZXIH9owK
xcZroIzzipB9C2xNp5U5FSFfojndWiSiZsgalhrXaCuCTiEy5nBGbk5whKCo
1pWET7j/LIB64FpJlHmX1E/iSxDEliKBA57MwWtkW6EmFniFWottexJC8gOl
bPFVUN/tXTaJfXWcKlqwXBvuD0y21rvJRWBLRhLEutUDx0tjp5aASdsiuJd+
T/hpA3dnzYjJApxquX4FEoMPgqUSlZR59d0t4rW57/LDXIU+MAK6/83dqily
wElf5Li3hC2Hqn9W5NZZs0hHCudxzpeVGbIKn/GIx+oIV0BMFthnfvpieXBo
VogfqaOQcwBjFhaamEOGiCs0g3gl6P5gOIvumzlLoki0434wlVRFDUBhgLZJ
vEsHqaCH6+NbzA1E4Ih8ytdJn1RxHe3tSz+IJJ0+7N8RdS1B3jlgf5uAO1+E
ZipgKYNbNjS2fYOqUrcJ0virnX1wocmBH0xHgI0gpNqT21hOfqqE7TK8+fV2
7WT4tsLTXwdm+SOZeroHOPjrx7PTb4+A5KflpIZoryPVotnSdeiSD4LRQFCH
Eq24YLdipKL9U0qZFg85Rx7is9cPZGMSZKYkmhIXIUSlJNSVeJDEcDTEbZT+
HRVtWXIQBtkJ8EZSOx8+00UfsS1Qy86DIRMO9KUeWyeQJNGCU4ZxJayNUBpV
xpvhthoMPJ0c8kBCQHhBuQvjbEn+2sV2ZVrI64C3UtXFzLUCciYSPfYAoK0m
2mtfRDpp3hLTU250YYGLmnKc5qxUiNND/4BkY6J6uVBQ9mu5d6NZ7kqXLUkc
5hR0NaMtCJlS4dEP4duDZcLdcvNf8vktENFoTjYnueslAXkoJcSvIU81G1uZ
Q1NChAnfqcUqLs+aBZkE3C62SjknE342h4OsVS6TgiFgzIAAlVtJ3G4KoDeH
venViOBrZq9ZoBM+pKEdYbMwCMTVXAl5i+JtsHNFJx2xi6FL5c8VskaxV52G
BpQ2xbsX4FRXopwsoPX/j/wZQ1cEnZW8Y7gwBc+CBDAPqbtzHH8T30RcRjMm
goRP91Cbs2jEvV4Ode8cxLszc3AVjWjpat8nTqnvdtdXACc74r1Mlqv4suLk
54cda4jC6HZzXXv4EyX6KtopMRMXFCdRXAlmfL13QbSa8nicOJDjp7ouerMY
XoEG+NJBXzi6z49CooQb2nqpn0Qcumi86cky728wQWKAFmH8X+MngpPMbZHl
CqEBhMUB1EeNXg+HhEcVumjv5Fzqc+YLsw1jJiDK9NkW3GRbouFI1Pj8LQaK
gGDAOHHwB3n+RMtvIAjGOlGT1+kkvL9h9aKP4wxjWD1f7jLBMO2sc+Ds81Ai
Q4umwFksAqLUsvpvW6TdPXnI+uanbguVzwyHmaG91z5DK8HeEH5TBS/9fKXl
/rGaP296OKUx+QPqdbEBXNK9xzRHgCejWuHE07t2HE5qKvO7QuK6JcqVSztX
pEi4as/a1l+CECaAKXUZfa3o1/S3zBOy5R4tTMskjeV6F5ZCsqm25kiIQXlv
67SM9injuvFr1+mNm8IAgEGaHQTssjRsxnE1tzVV3h75vhvyS6VP5z62+3mU
tmLMJwwwzoJ7YGgHBhEzVGlHifHzyXtn4SQXMv5JTVIAGNbO17a8P+aSTU1z
EhEymZ60xOGJtw73J7fn8aPBSyTJi9sXUFtn/HopGXxWgKg0s101na0CEL6c
e0G0O5hmHhv9MpU5gLU6V8V0wE8V1K+B82oz0ywZvebWQ12Gs08OteIv3Bd0
yKBjvgObezKkauAeIA30FXvHlsunL9OE997WjzK4PQRgMsqoNKB7rfjrWYvx
yjW+/y1cpPlnTtHBiPhZ/DuagiZe/MxNoRv/jbpdy3NSHy39erQHHVHAlbud
mqiJqsp3SIb4b4FiVFGCfHkq0y6MTVKpWeCLby7TTiI0w9PMOhuisdiDrSqI
EcRO6FVX/+r6Nxqi90kqJsAiPJ1RfqdECksHPPucy0teHFVeSHdYFyNBM3jo
e6UGiZv8U73115cPSh5X5hLgx2Pm0zQoImivylHp4iVzcsXkV8m6ceTdfnVF
NRj6J2AwnChCkhEtY2HWPwqhw4qQ2Bwt6php8QEIQwejM9uHGvxw4Ze/L2tv
3OJiH7i4Et3XEWIxNQ7p481GERfHJYgDfoXSZQOoe1fWUPIfbAmX8tHvwpFQ
2fp/+S+YYPVqwkltirYS6QPkCe8gAKqsUnoibN047293Ph2q4ayTr4Um2puk
YVuDQm6b+6uU2C8w1u5U1qNd61GnCrOb9COdkASkOt2yonPTUF8gFdNXuVSR
iHW5ZQm4A/WauF0W0IAmJSV5Ea4YexHX01y8FElQEDYZb/w3SCJipvFDOOMH
s/3rSyfFaGfHoKbg1kob8Iat7C3iXvbwkZKrDNRjLPys/5DUixzBr2Sdsj+l
OJD0HTohsqa/Z6ZVh9wTMt6O30Wscx7aNcF0exyww4tw7Cn+mpdR7lhyWD17
t/fG8ibSPgpLCIYJMqtVIAP3eoHLJ4LbyMVZBBYT6aApzwZwAJjZF9r9myXb
EVV424Zh8Q1h7c+XRpvK5NLG84eYHhxAhdOZWFy34TJHl77VTkKAos4x3sAy
rGYP+3LAvGywO0ZTzh6B3kTNAuQ8zHWYxb/fRkRzBUkXysVGpN6oQilWwIBi
pVvbBur8cpJSBljISkN9EGZF92PCdQEgY5y7498nYFCmIBNpuulCwJ/oAKrP
Bz9T4D3fu/bsxp/hU21/M0ZDt0z/05vGxWj1yKAERHjNof5A4xfUBbW5fsXl
EuLHwbiYJ5S0BeFuO+yuDbYZ8il9M4cU81fiWNTS97z/UT5zpbJGOJx3AsQQ
6yz8K1aenHuuxOauw9eh/2h/+8pEeWgMwALLD4xSVVX88L2GpRyriOj8NI0d
s5lnw/dWJUYJ+dHQ8JK68+A+HIs4K/WQIlMrMJptw36SjjwsvxzlJn4xk4TV
prb51m8Bwrs0QmtMVDHnDAwkMNnC+rDuC3Cum/0ip9Ea2WVSAuAyMrbTX8xc
VDLV2ClzAqWkaoYWyzpE12NH1wxzQ60iYZap08g1CUTYjJz6DrjAJzOoernl
GAV+taWDWbMqRphbOteKXJ+UtU4ZUcQz0xWaZwtaVuwhqeiibZDnRATE22kQ
KsXJS7I9yqwEzp/CBGMgsSGVzQKbpPnnloXuF3V/l8+tWNAQApNdRsuTTHEP
NGVvSFCOzSQ4fHxLgtvESH81zxQtjd0r8VCQOZX8o9zoOXPyMJpBd5Qa+9Tb
LCZgnTqSEauD8/YweNPW01eHtOesmQdqG/jFtc+cYKWQK3s2mmgqbeHqsduk
64RtB42yu2xRTbOFk3vglDM+zmrjkGswKJi1YyI06X78xB1Foev87mCuEAWU
d3RmpG+y5WF7JGFMJchVFXNouUjPs/PUG9qijpmpSfr8+kse2kYUPOQaM131
YLgVvtz9J8tscYk81xyVOHYSVzCFdSuu0nQWNuUk2fhmA2Tdyxjs0fCtIc2u
o5gDrgbygFcpxxxgqhwZfeZ3rTLnx2rb6tynMtOJVBM0G7LuxDBAUE4rIGyF
u/8dDc/MOL/dHazHDidol7MDsO5L+ZKVZv1haVm11Ug5FPpG70T9w5di6uoq
x6bWUT9Gn8phhClcxulnMvzBcTEoDl8aS6HZWjKwt9Uwq1wt2Q8bAk/+wfJV
hE6OLvHWibD/DBWqjbcsSwvCD9QbVoxEdo57ab/KTwLBwsbYvD92C5k8H6g/
sM4GlS1X8LdJ97+Ulk09yTzGKGXaIFm0gaBbHVRI+BcCK1qDMVYzFJBQhTB+
bVqhrP4LRDLiZNv44meb+usIIcfJdU8jZ6fZu1IDHmAtppAneIlwdBkkZgan
k1GQCrI5Au8vCW6cgMZ1j7DQu9+BxCZ9rz+Mn/rA7EJkDMoIycQASiI8KXgs
o59028+VymyvRtlfWpDzVj2LkPDaIVZwVJ9LFdQQ2RIGfeoA3h1TZL+RvONT
THsTwta3/cp7kjrBFwK1WHgxXqhfTnlmKIqFR5eWJH2fnUhT8Gpv9AE9pAez
ztK4Nhudeu72MU7n/pXQt5t8gWm6g2fb4OrH9bHRru/Wfp4o7yUftt0mzqGq
EYdXzabaGNRNsNpGGXKnvvoU2ydVBApeaIgdZMHgKgttPfkSeGxA+9stNUq9
DumALrQk13bpjittrstFKScIw6lPXtQtAjn8AdHpygWAu2w5l2hRWUKmKXTj
j4/CPJUmvdZAcvJakP6wSc85f0dDajQkygH1uryKAcWLS/LMNzeslssUrmr5
+g9oThxyvXaxB7Kh2pI7Q4Oz47r9mMW9mXzXrDpDG1mT2wAeqZB84iE5el1M
D+KLh1UsT/tVpLObSbWOxiSKB+fnWnw/p8JcLCGsCghZerLAvohgCKWaXCPO
STtwdHut5Sxb5s8M15LV+hX+Z4l+d/mArQ6pST2tQyS3n1ekP7cQUfQI6a8d
5QtcAkVFZw8Mfwbxej0PDh1MWQ/cF9FKgDEuEYMcwSSwLF5qlqUoyvZZB2eX
W2KQe1pI3AAJyjUO9D0NUC5bFxxngAS4bdnvQ98igTRSiFw3Kz50nuafiH+/
q/6k/lx/byEfypHGEDK44X/rU0He4iY4t+nvsYkWGQtUbv5lBCVxlM18Vvwr
OstTGp8duERUSYfAPdL3H8C9FUMi6qVfi2XZfT1R9irXHNOkUDNtZsnT6FXM
EKi5vK6KUUPI9bgppWRuZ+ke/zfYa8arkOwalvc+Rh5uMU2slROOGUHmRTbV
vLSPKmUe9X7+Z+GkuKf2nlDHd1NkMgPZggbKSf5h3tdjso0K1CCKcn+SD4k8
M5Wc3hNzt+tBP/1qBWGyqtk+nX986a8AKm8YiBw4/LPZ1H6ex3kMRBM+cBNf
c6yYj0O08dB1WAeXlK7M9VnbWqQFKGKHUqKEp9Y3gzvbnCn/JFeGhpNiCTjR
iE8NH1g0hGeGrBnmS/DJz72LswBtQIMWrdpP8XtKhJJh/sFdY3GeCubgW8rg
NCIU/x21kGVppPH6jbJL3GK2n/yk2nils068Mi0SD0I/UkgGzjQpX1icnEA7
Rz7E9ZtjkjOZR/rwk2GJzmjKiGZCw7YiHyfvmjvHhp2WTb2fkkKs5Y7dG7Xy
Rzf9TNuZ6dYJciT6yZhg+1EevpZM1FFwR2hwzbtmhbacPodi6+zfEOhih/qO
OFAk2dDhCfWuxF0vzKVQP4PkIJuKcOu70Zb6gVznzIe9sh1C+pUiV1N9uG5m
dYH4mNKnzE0i57Atx7JFUC0tkoivjb1tYtkwR96ro+lbGw6+q2qkkRWf/U+l
2OZN/sluszk/vWJXs4B+fVYuz+WPdKKCCZAgDWRm674eOvNMqDOcnJnGmHRU
erMT27aShrA2WJFguytKAq+whsMyhrUVP4c1+OZf4FoYPkIVYkmaBbn9rK0R
kGW1AW09D/CSY3xS6S6h0ZyXqwn2w6QOHNeg/mefijox9f0r5uFnSsIDzH0o
K3i3w2y/DdIGJrfXPc+WLHfWdCNqtrcMt4PFdIz1unaV+14UJFvpJt2SofnH
RkuzPZG6M4rm4Oo3xpCq7Y0kUKrBq6CsWTNywPwG5fymfYtHS4tIgH+IVKkl
M0cH8RZbrI46LFWFHBb9WvXWyNMUxptmGAJnHuQxK3weMB7dCsHSeAx8mKh7
Nc1PcTVgIfR0EdSBeIvQWTkH9ZICvn9I0+fdv34BsbTPi/dNcx2NIsf0RXsD
yQEgx249i7YvYuTF3EDkX8vKWgP8M/Re/YdtIxmSo3M6AyyUHIeCQeLL6KQo
sxCYYoqBjz6Ro1XTqzmMznvO6QBcZiRFix0AxdqOo1ImOwEyRXwi4IgdwQsk
/oJmv65pPdNxW13d3usqxwqLFRz2J19GsQcIoWlAcqMpQbYZqzcrvhMZ/HZW
gj5AkruYYbhv2y/JB4Cxqd0QYkLDmXdWCJWOwgkg2gyL6Bjq4k5FKqJ3EaQn
rRtEP9E/ZUcfK3cziwmSK2xoTLQn6vasrDwFzrlg/kY/7QB5dpkQiFFVo+4A
QQFAmvZxXVXCT+Rl9+f3u4wlu9EeAOW8jhnKN5Jh9N6uzs/k+x0Zyd/9d0Dy
EdikQJyJKzZ2TYRCsgKDQ44wpEf4EBvd0E7j5eIfkzeYcLHQycU0BQlkpsN1
CoRXvpqEgywsfK3e9q+XcaXBRpJ4qwrRMovOvQy3ionKo0a94q9nv54+70oB
4o+26WnIXOjnXyuePJI2S/817jA1JGjKY0Gk4pEEfeVZaL9OthHhWQiLnJJB
bYZgWDkHReoI4Dh94tCnnMaL6pXsNddcMdQA1MRU2hasuSeppWjddhlZtj8F
DzFCcx5krVBjK4u+OlW7XtsmEGv9msCgM4GSJnsXFlK5JBGi18b/wDYkvsbv
zCtXGCrrTcGXjc7X2id5m17pPZRgoogQO/QWobMv9iYGttxhPR6EY0n8LwOW
xNTkfn82mNmMANt8S6+oVY//mFe4VEV5JX/gyamIPvQKdVCxiDRePAlwHwkd
pzxvc8EOoaTN2i6bfZ3Jtx+ewWCNgnBFxmNubffLK/GyOHP3TPNnsMapsh8G
8qMFasJYdQwsuuOL/vXn94SyIveWKA/jFKxhqb5Nu4mcwT+zQTiJv9GU2a87
T7MX4tjuiC6B4SEhFVkWZemzIfm+VV83LS/+SOW9bSji4JB7YXcFBwMk0iw9
AdlM/DTfVMdRf5VT4qdlUQFizB1f/XbGpMi/rr147yVt0NvEcMG3ysx9wrr/
by0QJSX/oCY39tLzp/FW9XeBgroer7gjpY5ENwFCUAvafowLuXmLmt7GgUdD
4qq15LyCIgsGMn+6d2AKGYK8D9TyMMszAmpxAGUKGpfbSlFntYKylynHWnM9
l42LTbtji254gkFrxWXhuhOgjDug+YBqKMDblpw40IXqyFXNbuN51fDTcTDF
wcqjR9jLFAZQlZkVq2I3Tt/7DJ9VCbvgrF9I308YoKD9Y2II0lDFOS2rY/P0
HI1reQ5nrqUN7Wu3/cXezm5j+Uk6XvS0mtxRGksVNLbmT3Je7Aoci7NoRdPO
fGyXpJkcvpI55xpnIyR6Z6G7Un29fpG0H5jyjUXoWhz7EmL0Q0v/6XSz5Lwa
E1CQZLIDAtQMFQ0RLeo9kxqFG/1aurzkEk2yNXCjRsdS+Zhhg2lvKQXBt033
sISlJFNQtA7u0hRuE8mibHeKCaT5X7NZzojvkNXWKpVbi42iF4nOr+WE+iRc
mJgOep+8yWnwYBHz1Fl0odZQE/IfAEdtwQKstG/9FEVPP8eUr+oxOq/BqHhv
kS/8pUHKXzuNObyV8UNy1qrDV3peygch+qS2y/Sov5yyRZd3Gv/IFHgPjVdE
I4h3SP4uCHLOyQHZKeustRISaE+dgvqN1uUBSOmZqYCFcnmNlyHxF5YlLNmC
rKrgjc3EqvlfXUPaj6TfRCJL1sXuQj1zvNEhTUdNArWLJMhGw56RXTqNp33X
l2m62Pomwmp5eS7SGublXoEwp4lzI8SxXTCpu19vpksEyf1nz9DI+WM4MGIJ
UHA0FRiBrM2rnRS/YAFlVBEZQM/fmcSuLe4pI7V+M2XEU7MSG+nJ4YaS4cRL
ltXaWc0xOmHPdZMIqpXZCP3y509frlTiGYD9YTmyCoaHWvaH6BlSJEJdCLhc
UM04g9eJ7YsD73/1LdtEFgEvH40QNIK2liUaPOR9c8z5ZGbn6/NaclcBiOYi
FsMBkQ7qM9NgmeK7X5S6Ts09NH/ucHY5H8IwWjK4OmXNEM9mklQWwsbnP1CD
QlXXQRjtD1rGFHyoiGpGoxVIUbwghUkHLiZUPhwt+RuheomAIgOnedhzwKqR
DhEheLC40WYhG8Sh+PbA/lZbOBLhQYXdQ7EhVvBtMnrEBgorlh2FfNkMKdfc
TMjx/WkvWZ7HFupur5lUg50/bweIlOp4uhLhi2IpM9WC0R4iarGF6sf1wZc9
XE+h0riMmb1NQ7VYE0HE+40yAFeCvyNSmoyurCQtZsQOQNfVFCmo0k9hYDDq
iwdVfF7wXrIT9DGBFmfj1XDPWq5Ov91J9GEEqmaWiZ0Kvp9KAWvw3k13AVIr
BjhqfCSFqWfowkTRreWUNPzxMlZs/kii68L1rUFq+pQXtH6o8ANsNaCb8aV8
vFeDbqhl9iMg7/vbWUz/Il0LslQgeH+LS3tDv29Iwkhops+Qz1yYXpDYA3A0
Ib0Ay2dbupV25EueXJnlsJz90fNidy3WfOhT7wqNQtg/zgvk1FsK/3hmUpHo
lsvUKPXPe/F9zGalJKBoZFWYXs8LLORUitC7nV9j1dZgYhf5aelPtIf68+JN
dKCVCBP6XiwPNdUJLBW1CQiZf0haFubAIhIe27p8VOA/Vk+//Ml9+lX/Mspl
LXrjBqy70nRgv46AwhYil7AS4Y/U9aziLSIqDKHBYOMO36Fouy/Xevrv4hHq
U0t6Cokky3B4k36Cg0SPn05fH98e8scKHX8hpbi5nTnoh+LfaHGvBpkfklGc
EQ3EDMaGMlqwM4gWHrUVKPY0lIkxKbx1+No7E0vHTqaUtKfOo3TMrBMawBW1
nyQZ3Q6tCEQbhDPf7RvZ35z5ph5dlNwHss8JDXtlEGjYmyrE5RSh2Vw99ipf
nkhvDLIX2PleQgNYmR1cwmVsJZisq0tiAs2Rr8r8s8sSQ2FaIlDLxZKn3GeI
+oRngg7ZkmxqdgVgbAVZL+WO34lIS9iq9tR7MKVqJGIaYRRKueTl6IfPjJFn
bSEwOK2K05w2nagG0NGOu8Ee449JthTI6ds6gNEI8yrEP6GpjqXBQWLEzlrs
a7whG2CM1MXPJKLgYUVgHMKxayl2ufWRzSuBjx0+yUZ6vkkMnbyDOdnEsg2v
08X/MP3E2yejK1hNUkXpQORV7Bf1KgWiXfdcMC9WbTfABk2HWsHam9Nd87I+
I4fbfjTXTsrxblwKWsPSqUu973IOWEa5EW2J38dns0VgMPPSfuNWo0xc4zi/
3TGC7Hjz2a18mCnWdJQL5dONd1V7RfNolCRlQUtvoKP7XSHfyehjVV2SFCel
YqsQ8pGLVp9+73cYtn8WzFMCD9QGwMXTSxXtKh97L2yUgYurAQpYGnHbKzjS
tQFwzh99hQ38TFuzwDHwdms5OcFFd652h0+/IRq6eT6EGZMgzH+l7RmggQfI
Ha/i9yQgvq+Xy654uovew/EeV8ZfmmwXhrd7PeReylB7XdvIbRGcQgpd2B7I
5P+Rw6kdzIXwJwKjx4wfez80rSKo/rB059+zf3lgmkrPlTSctuE8sQbVVf1L
fb5vwcYsloE/+4K71AnXwgQ6EVhl2ihVHybEI2UBQ1J1A0eXZd5GIG6EqhYT
0OCgOOTv5cPF/VNa/17p71/ANGlEZKB2GoUVJRwFbiWAAHvRthQzOjkPmttQ
kksSUbwfm9JpxXHYG8afUaQl5rUYW5HE/pY3YTC8Xwnw1T9JDQ4bEOPw3V/1
Ina4KrxhDOJt4PQFRbZWm9VxnFMm18BovIV3BuoWQybEuaBZLrxUrn03MW3H
UgLzT/sxzsICaRD9uucacUPE4JgjECAz2izcSfajfNKqc3aSXUG/GMxwJkec
dPjp52eNNsLShhOH8+hsh/YZLzzBeVYUhUjPjuGVvp6IPuGSzvZJAuWZz72O
wx6vA9qFgXj5CI+vfTuRKq+X40oz53Cx+9jFQpy1YhQq2mzHfENFv7Ko4++H
S5F4YrhmchIanj0fIJTsux7/Td/+QsFk2HioWnRTjSWuVY31+TSxjZW0I9sE
wn05AXoFWIzVmQoT7hDeMD8vVFRcJisjTzVk5AYR5El3iXVz5bZGqyr2gK3T
LgLQfEu2hX4PGYOE3sejSgSD2KZDdOeYC4UDNWD2HJZYapu4N3UEsSLp+p5i
j/M5/riNAAweOgW7u7e53YIUSaeC8dcZz7x3rQkJI0fYN2zScVTw4+eHs4PI
rvYjw9Jp4037rG7Q+t3vFQ51tW501mg41Obd4RP5Yd6wqQYdFx5jXP8RrMj6
+63+if99ut9r7i8N+4NyJNVCLcoLsbVfzLSKJpWGxiBkLwMgTvncDFs6DqhI
E6Zvbau+uqJ4XZGV/TCJ+gwHXA+uK8re73uKTeGKz9pBEyVUzwnavSYW47sb
bArpsSIQz4DsvXvlmWX18kQluVNGBWCkhUsjduyvxxB/Vi+Q4iUMRGh6Hsh8
ApzW11wrKvuqQ4sJYfWffuw21NrK8PIjoyK/sY8XgZnufr2wsIUEb8xO9RSJ
+8h2oBzw5A04FQxI2LB2VYYWAzdv8P6sO/HeyjE27UiG8pORUk96ZfOi8UfU
gzELYR562Tg8eqzreH50Y2aIyTPh2rtNh9akR2Bi8aYjrWhE3CICd5xJE1uL
mQQHzqacULv1JDIBPQFSth6GOkXRqJlg/y/YixDYeNLWscUPPQAK0vSVyZzc
gHEHLdndqZDFK4fou7VF9t/HUxxr4PDAXpikQGxAWECFoq6inMY7tt9EoJUt
HjYiBYCPCgXb1jqGREkuBrfXFGbtgH3A1ZjAlSwktulO/KQUcXVYqJ6gvEMG
2BVQ8ak9NqbH3/yMlBOJD9YNegR0wAB8q0bNzJ611Wfc3Mz94OnC5Pbwu8YT
hK38jP6jal3YSAmQAfIEl2GTFMHfCL8WC1uszEg7O24vvD6Dt/4Ac1dMGBOb
p7B54YdoJZs3QG4bi1DxGdO24JuY81WmddMnwSwpjoaqrCjz6X0G664Vogs1
k1Qx2uOckLml3Wf35r6b64e9OFgOdYUtC2IqEWUu+XFM8ngsNjMm5WFR7Nq7
gCogf53EDhx4GJ75gsFWX8MQ9bqzXG4UzerVP1Nd0u6m7UXvS1ooRibdZ4zf
1v/VVXwR86sqLy42gXX346YfiOuv13bTOj0btgdEF1nfJa0W53myNC8gUJhu
UylzA0MWK4hj0f6HvwtobGZOpjxipshxo5IrnU4UzgTyhyLpDvvAsoUhQr0G
hxU2RX64zWOGrkv8RNtDNpDY+HwjreelRNuo8N3eOH/bnmJHlifBCKZ1JrhZ
zT/m/lO4Q+ZmkItVQXXbB8Fc9SvVZ0yf3Ca6lTAs0pU/FbNcns0n1EYzbvBu
lXgYDSWl5Slc/MBCpop2dLeck2uRIEB+x/0F12M8B2URRtV/yzVLE2Y6y3KW
73RTdYYlSpJLth1BadRflaSZH8JRuHPILtGyasHwSOI3fbH0aC9HwV0+jdEo
eMpVaLcXvmhKjuDHNlBFpXWfYpY0fLRhPoMJrfVxTsAur/2naF5vCJ20iNTI
Y69Uqow9MP+1qc5UHqXAF+aizFeBG+NESjDpTPUCisKa1yEsm/xZcn2wf0vi
xGkWvJtq3r80HoFTv+Mcv5jpcgDRUIRgXEH/whZ2sZO8pjSs8TRY3eQdjWdx
rcGjfe2i43e2hkTdh6ptNFjNDLCetSHvWVSjKzniQeiBocVeQMLzLDaOwIY/
q+NnZ9BZIwYLto9TDJuYrPL8pZTCk5vTKvJ023bC5s7DOsi72OYZ+QYEhKWR
LmrUe7npqcMrakuWvSytR7vPTfEw4FS1HVb+AvE9liATFDWFY+zpjE3YgBBl
Djja5dMcVFgSIa08vo/lJtFRyOSOyD4bxL2AuTmk5aCxufwtwSQsb1J30kh1
V3r5gFhFN/Nrj6ojil66rbvbRdCwzZy+qedkceftFXTP4M/64OaKmDmuio3Y
plW/TTll8r9P0+svgyL0cnrCcV2bTP4RFWBwpCa08aGpVVTjGDZIRRZSiXpw
pO19opvFBTWNj5JFJmZHCuHtlc0idD31v7MaorDK8+cQKBgW6Ng+pkzwK5lo
d6Lu1PvHIbCC8taQKQ8F1WlXcKe3oyTD/Ffv/o9FB3hiKAM5v0TapIZM7IkC
8U2FF2z+3zv7BAbepUf90kazj3Ioh/P+elkmpjw+NnBN1wPazB+vokc31Dr5
FNjBF/oY0r8wS8jXb3M+udUm89T+WhxJkZ6DlB9rsSbvxtlPMupj7jkeR5NC
OQkksdLMTjp84ECCx+Oa6eMwiSEQJwXHUyWKgLKAvw8LzPs9VmjF5CGA7aXA
vw3A7+1qug39XlP/RlaVFoUgIphH7bN/fv/el+7qDSryQAC4uCC1VGwq2o3n
snxHjtiG1qT1udH9vjeGGpOIRJp2Ut8nFWHRJ5tk727WsR2GTWJgQt4qzmi/
9TwG7uHIq3lnhcSbX1i2491KOXIWg8ZfY1/GBkG7IkjFQdRx2K5f4lk4Zko7
klp6dPr/lHzjdQUqRk7AnzZP7jgT8dYS70CQKwaHUpQT1IvUoMGruKvXryOw
9f3l5Dkg5gEs+1MLQF8KmHpcl9U58uNLfmo9c+1NmHMPxTGfh+LC8HD4NI0h
Jc1EifcBqRDjGbFpVOBjnCp0FoABbOQSpHx25C2v36ICIuTsT1MRLClW6LIJ
X8pnB94X6v032HS05hx/K+xR30gkxyBjZgOlgttIJh8k4WN+RKeJo24Lulup
7eZCK4Zfg11olP183rZtN9FZb4WAesYroGQ+aOEMinUFEESkA0h1IEsSi0S7
rh0yCIEMXAPa9THXEDVo8azcJLzv5LGo2Bn2TdaorX7kxY006LVH9V8DRyej
OF+YR5ZQgHJ/a4Un3lg3+OQnF9mwtbEtUrqQRNCpvDRORT4CrlNT5ZdqxgIe
mOnbLStFLVE6C9lADr+u+Uz2dJ7/G2D836bYRrpveQaAh5QzWwPWHOVsHFrV
Fh6sc6aSfxhNesLYnxqE4ZQkwIOUSxx/+RLzUOFJvPzELr/OidOEMvNtNl1E
Z+X0AmDG3b0tct4Ld2WlVatMjQ9ngKQc9yOSxRNq8jDWmuSgqfpsNHUfk8Az
hTLJX2yQjrTOIRCf4gaRq7UxmAt389G2KiECD51ydpVYuuU/AZVDfs5Z/tyk
VzkxPDZB7AgrTf84Ykbkz0iCXPSBZc0h3xywic82BdgBNDGj70jkZ0WoGnJ0
Gd5un//Pmz8vg4Sy2t1JW5eBxlRG5shsQ+O9KE2AlyoAr9y5fCHHb92lG2ez
4OXSa3O2OzS7drresnMfv7Qxh8yQ4WisPe8UvgRRvmI5OTsA2vNGZ75XfVTt
SdgIS3/ugj+/DbLF1XgmbyjwZWgsrBLTyXF8NM0GT4dGZc7K2rpna6RJD+50
bod3xv/M1qTql0TXdQCXZRwztSry5zXPDl/GFOrErzcM/fJMZd5+GjPmGBtU
T9r6aiPzjuk/aWcWYnhbUG5fZHDw/w3MlWTHQvj+MOAcqaVXEafP/VaFwIk+
5QZg38wEdifIokNPu1PLY2JVAmrUit1jGQA+eHlM2FwjVZi9DKKydH0XY7TE
gUXFSlgCFZBaj7Uc16ttF7ZNv3QinqSJyJasCs4o0oNQTvcBzxUVhC8w11a2
5/WZesHNTyov4FU/v1bON67zaHZC+/fPCNZoy5qphkMwFeRq58IUW/QztK1V
iJCYXBpOei3P3k8RN6WSJo3NyVUHDIA53EnvbKvbKUGqGBW9C2sRCJYFlY9h
A58dA+7QkjnmnM/MEQHHEHLARhK++/3YZODpGdLh259cZlb6JyNK9vwr+yxt
RUvCKmG3nUnV2CUg8MMPdY8cyugpwGHzPC2a+X40iOSQEi6rUfXzwW/eSfJs
Rb/UBEjlj1UC6dds9E4IHs3AUSPOQUY3ZDk8seMd+2GOC5oIRAFrN3iQQ212
uJNjP7uULpBgqEoZH8lgDbJRAyAuebNduRTfdEXCAVpVvogg1b2pGJrX1/Ws
2XKleyrqIT4svwfyOat4hovBaeFhPSgNCijnwxf3Z2h0JsxdD0fEHlA8DEri
ntt7c4DkZlZs3BOGRwgcoebdj56QHY8D0g1BEDUuNaD8J/xjC95UpYFld6is
wCnyuc8eiF2mO6orlbKMGOTFsEWlk62kffmfQGae45727/2YQM7FjuUrq+eu
xD8y6kShxB7GPQXXTQrUKfOdYAYg3/ys7D7sYo7Ttef2osfmIwORejGCxwWN
qLWNY9XRTvdC1ycCrC46Sq8+ekWBFfKhs1+mcSKKmZcv4qvPurCkcxKd2Lfu
2T+J6oh9gBDGhNsjjSPVwlbo9M4hyKjx8gDD5rZ/nWo4BbjJkD0eTwbxk/O/
iqIGkpO1+KiJ2hcrgVIG8hM+jQ+iBKjrunHiX6xd3tNykWSoesHvY/vrvn2Q
pfeC41F4FYia3KMiVipERFn5nFtpkdZI4VgozHmTbYsF3uCALfmRNajLsC5u
AKj0ige50cjON553RacxhM7HdW7xyOuOZQ4r8DSe/aarnacCYmWZRMusTtZv
Nrmw/dhWrelHMXPhoSfnUIzZvIY4s19I88dsSOv8+IJcBNRynQxFOORw5EtT
Bgwop02VhuPlsorgSCsJBSH6Xydf3Ld6kboyEWGVPiCYNsyzpfLBZjsnEKXd
Bt8ya5Mtdh2kVCmqe53UXalZTQ9xtncmfYQ4I5jLP0OmTjWTCbKZqwoJaIjz
qWvoDPfHUJsEPHhXMbNfyisVtWrKA88Io/uwNuItNzwxw9yT1JpIo0FZ9y5r
gKt5iqriNvwU8CN/lDfcXbL6Iap1u5UvGzTAJS4IIOvKBs5xC7yMYh4P9CoX
EwqyyGyxl5ov8ORz/S5AFoXE8COecLmR7px4+hvROT4YFWm3pQoj/+BJEZDk
JsnhSPwwmWCZSn8KqEz7WH28ibRkawD6etq3l4nsyQPyHIBLpRRquSm29HLr
elAcHr2YpPdw2vCvs1Jb42g2D/+rw081XEkaFb6kaO/ajJeDCr3wlQnsA3Wy
ZMam2NJ+1n3uzA5EpL11G74mMBVTkkZGiN5T9Gg9+dfpv36/RPXfcsJLpuqp
QGvWuD0yam8VDEboAewBAKSheHeHqrfIXOZW5M6SsUTrlKNii1hinrvx1d1w
WoAt6+EP1crOzDAqMqReTHclNsYXDvwC1w1osPEKD60yUmCvc1EsBCubQvwG
WJxhAgqXK2b74H+m0uvHpqjGl2ZL6oOUMhazGdhoruGtoQ9VOt8CW2aSz/vP
meig72ziYN+LZfmcG7qQMnrnJ21Nl6wxPfEuBRiSvvP2dBCOBZfO585wxyN9
Xpr9cERasAC9mAp5g+akZHDlUBaJ2kRpMu67PZKr5dHnwW3BocpInczxWdla
ILpNZ7WStodkfsn7jB6tWD1RpMM5yiFKlY4w49kDT4FxuI0m29fnloc86XTe
QoWjTECPvfxYo3zdN222njgrm0HPGeXfa+OPoEAvGtnjgUk8nSIP7/KBwAl3
4cL/uw1difgZXuDDI2e1wd11qpBH7tfDaZ6+L36CJ25bqbpCy1VlXcxDLq5I
6EEGmpKk9KP71Xwv1fQYXewOVgEHEpzvWe3yAPR1tkaHOYFhQgNUuqXJIAf2
tORKD7zOgLr303o11CLuHc1fn1U8iinN/LEAbFRoMLb9IBEKMD3Iuenhk4vl
wown3npRQlsmvcJv2zvTGtuUQuur5iV9T+FIJmSna3T5gBo9uyNG5NJ7W4WD
g1wko83gxBsi88/h424E2m+qnAtwnscWPSF4lllLmj9NKrPrUxTAGkZRfZMr
F2WR8ZnuZhJX61QOLlEQjDa9ZJrzkOseQ5yxtZsxa0Px2scnFMRAi4+4IQk6
IACgVZijh9AFvYrY0W/w5Rxnx3L25SPJW28Wm4AN3iv1mVV33gtOI8+E1zEs
YdC5Irg4NxECHNfIqe0k2IEkIlLiIgNTV9ReG0DefJ2BDHNHjSQWJJpOLfAn
kEH3B7oJA2bSboG8tbUnGYsvonTnEdZti4VQsukAPq+AzweZMIlkTqAIxwQV
cioCviT3PY67ayPuV55kEoAf05Uw79baO5U62dNvJ7RRZmd0s9jzPeGOwGPF
jbLbo/YcrUUQ5myUyLZTtJazWSo9OOeG7mVDN/uYGu5e4dSK8+9wCtlqVxnJ
DLkB6SJg1KhcSTH31CV/WKTQNXBAZC4OeAkcpA9j5EC/kVT2gxHqasEDOsoK
FOv3UuWqPpXWNaPNtl04+6IPnSTtGN2arItTMVqwEAgU4Y1SkTd//GwsycN6
3h7b6gAcT5HQAc6u9NU9aX4gQoFehMsjmyFu4nc0HoTyx3LcVn5sGAmm1dLC
GuPlMscPVkeT5AnlWXmlD5Fp4+iHQco92LJ6SVl5LSJ3fP8b0RmwR6FP23YO
uQzhiY805wBP/jPCbaR3wxDzgWVxdoQsDjKRRbvwqbcSk0xO98rtlqNCGeGg
K2h0jobb55DLdUHX06wjcOCQcF9wBH1/CXePo511nX+U2wC9ul2l6y3QXh+M
OogRBrSUj7oXz0QobQ3ul+2TCDBcQ57V4rakNVa9rlt8KR82nrzHpoUnaU0A
ZIhIAGr9OHkP+sBj1HpfBOVxYkGBMchgA0RB+a1f23Rkc5fo0Qu5v6dto8sY
jimQd9MkFynM7sHmPquVnuRwUGk0Q7zsHja3Lwk5vzMuJ9WG9AZKF3kuu8iA
jE9srpv8wnIJwDYiwf40M39zk0bhGPTV8vcAijzWAyGKryYqS6xF1RDDEK7H
P3FSDGo4dPzB/v0ifz4+4sKRSAycz+0zd3Y5WmdbqUUMA5mk3imu/cSWx29b
gZw7uaI9WdUNeqFrUKq/JPAByf5Sh4cdPuB6gfGskLvFOC/o7K9cNB6iOWYB
AWO1CKCgVOEIly0XI8jIa2UdYV6jUTIe3ywaDmupgrk0RwnGcqqJmMs3/TgU
K3VbUjosjyOwMKCZfa22Zj+Iwm3Nin/xw2nEektpCo3GRCW4vEhOAJZ9bHUU
+8VuzoUCY+g1V3gm7hE2ux8+AXAsByNMhUZpEeYDqmzwRbRrldC3QUrsgr7p
7vKmQXKgQzNPKZIxxHQnolH2tAs2NbEI1CYT0f0deGS2jkdjRLupJ+OkrkTX
6vwY3iWarMuDdXXwsm9c6fUlNrEs8UnqddoeIeQYov7sOMbiDjpSnkDzFt+6
4H53Z/YNW0QbR2pjdNuhwUovsHtOmSn7//CFZG6iY+nuw/t36rHjee7m3+Vg
fGQujTJrEdVRssA6Sh3D5UuflaON3WUFGMyPK3hnPhcwhYAL3bj2804M21U5
YypXXFNPOSamWENQ6UlYtgy89l8aYtSUWqZENV7b2eHt7dmQ6tUVzje7x0py
T1CCY1BaBs1Fme88Vo5RxRYGknJAsIX0XTBTJc1v5gxtUEHBNj/t3X9nmKou
lGzmNXRPZhyAml58x3Hc46RZn9vezGuxZj6Dj18iP4WwgRPq2+11FIXKl27F
KmhrnP/NOrZMDBDms+H+Kfq50ryyfkHWY4Jk1NptCIS2sqwZBLuK1lFbp5Ha
Fi5wQaSlNVWqxqYA5moUvEPSJBYoscO1KmHaAkkzttTemmyj+fhuidxWJgTZ
qP0drSlvVqmiTIAozRMn1Glb2kk8x5nq7pAo6TVfLieh6IpTwbMeZM0DPWf3
Mhn1Jw0l/V6QBDya2XJBNTlZHOCT77STXTde3DDEwPrRnQFq0G8kAl8CgZAC
8txHXy/v89BRhXORvkEvRI4Pt9epVj48PbaCIW82mWUXsHCRriHZ8OQ+Yk+I
anaQPBrBouAL3aUPu7iW+zKbLy57LiCPaV5L+JsFHYD+3ez5P+/1Gnc6HKeu
HZfR7Z4YDa/Nt9XgZ/yaEmvX0c3kuqOOYU5WnLmLbzVHEi5cBS7dj53SlSEu
/RV3bPlUGEkqbZ6m6AKARGjaQTZGgSLS0FaBjfqHj87vRRYeqNzWOaRcFZYU
Txqdie1TyUEo8HJ17aEc9/lb8eWPRMkwrV/td+0ox5olnUcTP9q2BXbkmBW+
h6j5XtxaaonXYs0niBJ06kE2Na6iIySD2x+6X7pxofYJ7LXS2Ij98+VuRwOK
d0JF2AATd4L6FSFQp/T/JYMZy5W4yWdC94J3sQVXrI42/1LqGqimxnWZPqbN
bLqz5HdB4KiXGrRfdCllpfj3Ro8NLeGbMAOL6qTClmr4hfjWlLjF9V0y2Ww4
Ly/O+hGqlJMCjYE3uKp3VmVDe0zTYJcpUA8bHIFNvB8lDOa1moVy5F9vqWCO
B2Opn9GZqXPBqf/WMAWLKg1+Cr+mFRRTpr+dZIl+ORJfVkmSn/izYN71lkdX
0u5WzdMyyRv83r1S+34tpa2sjmvP0bvKXgGP78obaJMQYrSyclwX94HKFSI+
vyzdx2R79Bi7lyySwVgTnemYo055UwQfqfM8FP12yf/vPSpzfCY0+XG1JPQ1
obfemoVm7kL6V000nVyUAFieLAq9TaWzTiGWbOSSAON69hckq8CLJVNyNyXb
WZuixHq1Z9Y1csMePLzVNu+sbuOBIbzwATAEacYny88uU+OAqs6xCw22fhk+
aZO3M8suCCEOPfk9D5aZiOPrpIa8Doe+VkKJk5o4A/CFSY4ecDm3Phiqnzyl
gHyXYk159vpC/I421/nvaNMDVdCC6k/2rOK6aVp9yyQBKFbajMIiKaOODzID
uboksfe1VkND4M6zBf6lBueP0jmYu5H8aq/oIu/SQ/hVnT5kTq/v/1Lk3BBE
sB7aW8c6uaAHE0DKE1j0CXO05VC1qGA4vM6LQOyBR8Wj3g9TB/yVZSI48jPK
BDpygyH5kXSkFVQod3YxGH29ti5rSZyj8UW28Jckuynjn6bQRMKXqA0nkrss
u93ZDvAuvpReIIHzKtxegRqAfp9+JO7EtGeUekHe8WQrGk5xALMBRyCobgfL
os4UonEOi5CbLbAQftgfTPDwSCPKUgRfuqCDifEI3A+OldTirNipaU1nfc2a
RXsi688spUlYL78xSVZLzusmzh0txClPfSM3wFyX2xn5Hu6RsO1IV/AINmHW
WAuh5va0pErzAz4PZrMcThwaxnGP2rW0Yc8oMFAcKJFeLIsgjIr6DgUF6sCf
Lszhf8BQqFjdKucFNs4i+LPj0kYlACbCZ0C7+FQPz6LfJmOsK8vjSlFrvxdp
NeHNzkf2W9Upup8z89yLNexz92ahujHhR8Bn1X7LxI64WdqXHnW3Ft77uNdB
V8llnJnw5O7dRwhya/DvQzC/1siagdxv+14o6cHruhrHh0hzkdHr/VghrbX+
eoqxZzYh4cG0/35x57Omvke+PZYm/zHDzeUy/BTGcxzYDSu6Z/R1G6nldqwL
8kzVM0UpSGjhOCBhoVSO0JxFe/YNR9S/V9gFuQZPlOMkGeRgXDSMXpRnq5iN
FzwiIpKt+blQwgnhWo1yotb27jFaGazGlNVQY7fWTcTt0XwiUR98em2dD+3J
cAdkMzkLixBtm4x9kKgbmWd7e0XCShstWwwuNXgMZA8sIJ9Ms2EsyzEl9hkM
+HCMBRQqSXXnw6A0ki6UHEczsn52EoIYRjtRu8QqMwo9hgFe2UqU2+p3xxJz
ilGACZt6LqFmOhYIvkXXdreL06K3U18S2zXxJFn9tfqjmltyyIWxgBCg4Q84
ncM2DLS4rMKEJbrnm7GP7yO8dWN5I6Wlo0q40nALS2QwhTXRdqydqHfdDCRN
EKpvdG4ZkkRGuwrOyTuZNv2JMXC18YgXU4y+lqQCz4W9dNzTTYQlYuTxIBch
lzrfRrzNv785oyuvHSSlu9YiUicZXQf+629FMuSJUDzN87bMeBSrYi1lrBj1
GWG2FuDWBeb78zBXedd8lY67evriPuHT0NtxvzWtWgam+PdmBd0WflFl0xG/
xIWE1w8lsUWL+VaLmVl7MK0iDVp82OkQF4pKEYfhUmdIvo5IumqjmiAVlH9U
WmRUCS2QVcf6Xk7aJPfdJvnZRnFxZA+DWc7TOxCZ0pt8XuIwHZpdEVx/Lcjx
Wq+s510ofEVAXbz/Pa5wcNOlzs5uXMX16hYGydoaaKKQtIruj/GAud1p0ni1
eWMCsb06chHRNFmVA4b9C856gwVroguLgHMtv83oV4hwllKu4TGJNTuPpXld
E32thJbOscCV1qkJA30UCHwnGNNl5cQBSawJGX0fOWB2Gqdaba1q0iaWh5jO
hkVMf3fryymGdpPsuIyps0RS7P8mbb88dMtamJPsL8HWA1G8s5ZffiLAzcGw
ahSg/mVTRABqvDDilz1X19ZppP5cd4iRHBs1pGmpyyUCSPhVgFJmSIcP26Sl
3RMt3kFG5+88IiLRGiMd/DjnQsEEL1qUIcTEMVgvAZvJEvzYyuknjFHZrb1h
Rh71qGwGwI5ryU8U7TwmSJfY+PXQ8dMA2hhkuSUGkAW72dz85cdnHu8urYkF
lXby+XEH5sYh84/dtlha6lvqFZJsoV1UVfdkA5CWGCcAkU9AJPDK8JDvdOfX
CLV4E51BPOIxYpnc7EJ3LsCeIcfehn9T0TVabGUzu5GWzvYOZ9u2lch4YJma
gSNyl+AdVfCKfrNP+6JIpXCAR5mEV9gc5tdmCuWOiX0JpMwkhYPyVJokRILH
BgtRwUcc9xHNVIQVut7WQ4Hc8fz65sWWf/c6sGTvniXyNSR9NKup6qBEDcD7
8DfBjTmi3/D1lD0mTtZd1yJVo/bFBU+E/NQ8srr2SLMxlauZQme0dwTJsGvc
udXaJuRrvIdxR34sEt2IkOGtr3UU3uqzvxPH1BRHOH6VYhgoEXgku4+hqsBv
/geEGruCqYMu6GyxAOQ4Fuy6K+t2VdDDcFicDh6p59EqK2ihozzNtw0xHKOM
mQplwlQZnBq7Wbj9fZbmXKsQRKeKwPWyR484KiJnM3Ty1zElrJp3wO3Eqa0O
orKlbB6/igdpeR+6twf+IpMEwQR3aDugoIa47Rh4764v5eDqNfCE9N3FZB2e
M8dGlDaZQh2zT4904kAekHHdQ1Oi2BBBsJXnUjrtRWYUsNlN3p6oDUBbmy/+
LB04v6EqnxdzpRP01oINt2LGl75mlRenQAKXM8mJwyriVMaXHUSnP9Wv5+c0
vLX/D5aqb1OUxUB0/eN6TzXOg4IgeK6fGRaMyEnFVQ1LwrEGuwXwH3g9Icfp
87MV8I/QO+YmqFdVEUVVfhLkVxjhsk+k5TzanbhqPLWnAfPtI62YDwIbbref
KbmOboZ9xNW1r3gzANhLXnteVxOZKBT2pbVPcrNiDsg6PfFSg3jTrNAtzOk9
oXqHs6sIXp6ynd6dj/9JGDFQo732P7F+ZvW3R4qT8U9bMrdYX+y/Tc5wIKkV
NBb9gxe3RzwQAykA4k3obfHLnFKGBW3cLKhJ1pzxZuP1Ys9VL5lLzbwWy3dc
NzVIeqskFdV9L5RYOTVlbzISsn8iwECCZ9z+rac+3CitttR1kztKziDJmbhV
bCbzzzBpvILJI+E3oLS156WL2UDZGDRI8tMDFTW2PPNL2+icAA/zLtsBVwTq
Bt9XsntIZFgvbKAtU/Z8eAzxWajbhGOnQMasX6T97teSB/+JflqJyOvQrbl7
0PJ7YsP72mzcPoGiiUib/p5U5W3V80lHvpVQ/bhGjqzIEeykMrS9LE1qjDXr
8FrVNC9BXmqHE6qZaUJcTHpIrUOMBJbqc5LMvQrMJv5izFbKHYKEfcy/6Qmu
OHpYOpMQnyGLzZTZNGfSvE1NUjZ6XW7YetRPxNXqNXV0WjUQVqFLvKIH11KX
79HZyTRtn2x+WU8pHDekNGhouW5+RV1IYxgaU3m6KIVksKAxlaowQWtlP32k
lA90/hT3d1HD1yBIyVvh7fR7Yb4C/MFyMTmxNAYKulCHOaQvE1qSrUusigWN
AP1zyvgPFoNKCwz80bQE0+5RCVCOFFm9osU7KavoP6pp/cpcMwnWYUMXDSJL
N2tcF0iwHXnhjnVvXrjI6ZYMSVsrXkY5fGXCXTb2H/I2nIY+Tv6dSiikIeqc
i8m3MGLyT4SzCy27ZC/JiAvACcxVCY9I/3nZKTMfsmzshbKfnc4J+JQNpSLg
r72sRqNKnTlHpQD4HQxsa9qvoqhKtW7ONd9fDeQwbvzEnOH0Qq62FmaTrXrA
YowBNcPxTbQwi2Hz+2OZP9s8lpYSKpO1HH4M+lI+KVnNtzMYH8GscwdGu/4C
JsKrOtrrZ6lVmpfAZvSYkJFxzLNLcx3re8IXicciTi3xSE6vqAGzuLcZ6cMz
MwUa0d0BMLvPwE8DZknywXiKP1u8qK16e6FBkLAIvU6erWZ9vpaQBWzzWKID
Jk2BypXLr8ggnISUt3L3vl1z8dpyBZp96Lk0nv444R3lf1dh2GO3uNx56C5Z
UzlRwsSH5dr8iZVegWQlDCfZKwEcgArWRMqF3Uhr1SQKdUWiM7/vVmcGER1J
9EoYX1ID7mFAndEYl/F1zq1tMS+giaEOueVJNa9edJVdt6jF4jMs9dd2Lx1C
Gu+9iyBPhqSUjCBZ0zvMyQZLw16RNE79tjqLpidDzSQA7JLP3PjNsc3C8JbY
S4jX57ZeBn89dsSIjAKb3Yy8kw+n8x7AFbFDkOwnkBHUWA70geWIJxp/uKdt
w1cZ99q8C9iWw9iv2SmrntrKmF162xHvEJeDGzpqK3fNGyYXpvmEr59oVCec
o6AnpGjOtuCwP+kM+FDcjhY7thgbJ3VpxYvC//8p5EdIngKiibKg37cf7KKM
e73JO/91MKrJEWns5c84N0MGK5bEp9h1kADd9w4uewqdXRPijqJsWpXL71Yt
kC5oKwIHz1Y8rlGkjZl+Ag+L9SDSab3kfBBmSpoo4A0PTwHnn0ElyDY31zb5
2GWrVLTVTufjM/2YzhjtSsnCuED6/z5SfHFq6E219OD76oNlfQHIV5we/cG/
tkVMb2E25baUTBH7ngqbCtR1mh+9e0LDoOkCwvYlyxxi84VYNpNfugtR5xYv
3I+B+ugZYuJy6hf0SyGlpKov7AQoUErt7N8ZCLv2UzxYR6JhYIa7NryQrzQl
sbCgc5X9wQq/oUVQQ+Zz3fHlDRi45BdwI4MUPOS3rG0Mqr0BDIXPMV2tux+A
PydQfxAKJ+MKokLVZ2yyR6nODeDEAmNIZ/msHAnjlWiqQ6JhWb79zXT50+mP
pPuiuOW2GMakqpaczIfuJricnRG/z4GY8oXu+vy/Gjv5VR74E2Q7877BjRVU
jO2oOBrKejkhFmDUuvQYNErn//g7CBswMHoGFyHtfYBWyI5DcQY418QKqMA9
HM6YZBc/yd1Gzk33kurzG5yC9mDxus+0NxloFBy5F/7roOsJFhiHtP2QMHP3
nBOuYLgfCG9TfmylcrYscHyHI2DOqLRFX/L/xV9Ph76L/ddFuFmrnv3eI4Bp
EYVDoy87wc4FyFKiuGFuEuS9ECAcbFFzmloAbFLK3KlYIKg5zJD5K3qguxAN
Hy/sfaS2psftiAYi/xyxp5z3gLDCxIsNthYhd235VSljT6ksezWS2HRFEka4
WNXpQrLmhSHPXF6K6iNUDxSXezSntCrGDh07WKvKJOja0fRnwoSYVbdUcLMu
ZjEkR4PtxeNNGN8lriOtNd2r/tWYz3eo6z08iWoINrT9JJ4q94H5jKA06yF+
mcPfUNRYwnERfzChE+yQgCWUs+55Ss0YQKy/Q6WOaX0UTrf1PseiqB7fxzGR
SvCFFqnUI9xwJP5+l9R69DfpPKqThyKIHCp3kvuGRW65El8XTv6KRbKymSZ4
A9NAHaARctVhqK6+bykhkKi3b85k/xlSAuMaAiYgsCMiRcAFTluvKcmZsNZX
Yh5DlNOhpNWY/SqEE3JDhyE0WrL8H8JSRXEb5wrUv5SeqbkLLBpfL3/EHOUt
NKPpPZ4rrpilyDal5j7De2cy5sB9amobOxGAiyHHDuLss8pov5+uuq+woeAv
35IChAh+uTbS0lhFtyd6qB6ssJT20zDzs3AevWefuUfZ1h6keAxlzz/P7RVz
sy3ADnj6PVC4RKOjQQ5CK6TvBycW4ISQ041CTd/gBJPajmseOwG0W7gqE1vf
mrPWrcRdSx/tE1zP7Bqna+vtjs62+OGSmdHrsTR4LIqMAkA+4tKTsrZFIu4F
x08Oj3rSr/vAXuWTqGt7Apj5Lv96/xFWrtVJu2Uf09/8i/ll+bo4mEpEKQDe
FK5t4ym+0E+RLIbk6U18DhdkrlCSrN3/boGYV9U9AgevYWaqAsX7FdV/5bh2
R/kGjxgHlaEeYQDWmU/wgvI2/yvhDtw6enxqN1u7pTj/j2WLBsu5HyAuzNEC
NNTAqMana2TojKrfHqUoK12HrAv4N9BkiNdQK/1QqRQBlMaiIvWKsWrq4old
3Tbaa/Au0wxTuSGL7qwfaWxS/iJOouYLTG4D+ZKfaXGlyUd9PWh5Ojrek9M5
yrfkhzyCHQpSCXfgTLnFx4zLfTTrCgvBwPoyfJVQAm8ehhJChrPkBIoNoNA4
VqTO9qHER//UKRLKt9td3XWCHgvBiowPRkmlsuFcPlPAAN+s2fA6UH0FmgHy
X7H9SvXUSSCHrY1fTpcB7YwXimWh8H6gzfhosogaVD8zAvZjM20eymuNtJlv
sWex8UFDLCS+ZpkTgmHE3jqHmZlvT+/LrwFbmZwMouq6Q9MhIt4M+buh4KCe
uipdi2wjGaGeUG+eU45Fuh9EiKLgcKTYqqHHMMfBjgElUAz+O5xMuaBKFEFx
HQzAu37LOWcjRLYT83wkm8v4w2s1A1aB6j1F7u+HKr3Ild0zTnnhDGUOhkfk
PYyqoBZ+yyhSz/x0PVZYSjxpF7ATeV/Nl5aRp1WUlyMnCW8LmXRUuP7AoNK1
MPBkLbsk10UxZHlJAFdxKwVUJzHkOFKbQEtX0dehjeI4MhXVRfDPDrqUgeov
KdOgmS4er56d4XSCYisByWbt2STW6/Oga1/kwo5PK2TBwlQ3kxQqTE7pBxof
6kLlf4sUCn3W0Rrrny5MagHpI8Ol0tVlv5W+/mUAQ9EXpJXHqOg0vvyAKtLo
bpTc27GnIQxekl+mIVLM2IiaAvgzQo6GpsqtFUf5wmPAD008gzDyk/5sXDTY
TyTM6Y/DvLnlxW5HRp/OT3fYqFhyDhisKT3gqhGHogXvFbElbzV+3ByaKRhe
M4LBngPG9lgD4nkcydJwJ/rNts25D5U1Oovdra44NZFWRtgz9dDqIS/jwqji
bq91KiohLza+fj1tmbZ9jdjLp9iNiY2LshysSDK41nW//mnxt1WaMPYTD2/U
pkHFpWKRTTt/bas4MNhRcqLKYq5/75c1khqX2mOjqclBxhj0jXJaXmPv2vil
dgbTXZP691TpcPHEXOANFp/nsX9UKUgXsZUNaPkYdkDEu4W9RHyOoFXwrQle
NAUObhpxYVCJTXezOycGzUiRcaognTs6m+H7HWxJh49uJlSUqrA+Yca1IzGg
YyeaKltrVTPf0CaXOiNIxbHbi+brZy/aKpENb4AzGcO5l61MOBRtcy3KqSxM
6j5QhyHu45fkwMK8L6c0mFpROyGQJVaKaE2Ce1PxsmTFeDZT0hGpZCf0WrO+
5h/stJiKMELj/1BWqlQ73/l7SVlaf6Omc4pKgVuv8s+jQDzaYvwjrXeM32gH
arTp8SP2VCWwr5sE4UHV6OLfcL8Y0Up3xNySIaKCMZ3bTearY88LUDtFch85
lrLt5fuoAu4jDnVu20DBPk0xbNNpCGlcU/HH5FPm0AuaeLfB/S12q5xuVIB4
hQIg/hfHziC9y6nmyzXNx/O51XFYWk/V0FPQRFNV69pu7nM+8A8NxXKq1bRT
/6LVuGQD3+Qnbc9UpwhaShiDOY85xIZYLSZntO1TtweGSfIIlMu1rUJ5R+kV
lpwHOo3DEznsoV8pIll7NQ52Ec1GQWmEf1X7rwmMLxylBQhwOoipN2Q89JgL
9u6IE/9pFVq6RAPnr42Y2pMNL1xQjG5uwleH01jIz2Ybc4zCBSu317ZwH+i+
wGsbULDKLru2vMj493L30idbL/mAbHUCzHS2AoFiPIu9IOa9trZKXjJnT4vr
ttzRVMaGhCuUGvDOsjyBUrxrRiNX96zb09hbUN9IptAzUtsLd83KcHO4i8PT
YP5eyxQ046qId61pnMkG0brp5pT1gLauDtfUSUq0lBwq2ejUw010hAUTrzfA
2pYxkmKE4krLLe0q1SKo2hBA+M0ybEBv+AmSm/I2TPfgm6EXNl23GK3RO+kY
0QUDnJ6TeQzxxpgfnMH5ITzcUY55hqpnYVEri2tRwytw2AVILao54nwpL0LU
IbHNvzeRaDmIIJwT3Ng89AvkpdkCbXHgPJ0snTaeAR+oSYmlOMCA1NmaK0ai
adRvz6hlTK0Wy0OL6E15oVSRXSDwVGuvGSAb+/CK5TvYl79+UwDBp6/8oFLp
d+/SQiMJZdK3ptI0w2aMv97dKT7d/yZZEMNdM2EFKps2hBls4B0NusRohORV
EeTfrTQboszVbW1wfngPSIrVk5K+00vL7veEBnkRPug6dWoPUH/RkXPR6JBr
VoA1ICpii+MHU5xn+HeeZ3hOhD0NSvM1wxGDSR89tbv+GQeGh5ZJpwXDRO0Z
juAxYlL/hr2ERF7HX9HO9nPe8yddykyqYNBYyUM9AMSwF6DCyflRY9MtxNzL
s3tXYhecHsLwu+EVZpkdzt2ErG8QeIlMaOAj7vXjwwhQWcW2OGZ//9aFzn+2
Ez/L32m6znHxkzrkFbezRXmWZVMQAOCXQvwYBFL/dHU0TxCrAiqFgiC4mCxJ
lw2s/SP+DlM0xPVjeJpTOwvj/AC0TdfkX4r7oZaSwcUCh4jQMpSdukuMu20T
2uSwODr+wt21O0X46QjmhN215LTRrAyRv1ki/glv7RPMQSAlQf5YzD/yXYGx
RMpkJeVCSF1DiblU2FyIQcRXY2JGtjCO0nxOpid+uAhikRPHcYtGyozOrpdR
a58t3kggEB+GLIKDbFo2PIQpBThrBhFs0mRRQUk5gxpV8b+wgn7CpxlHSb1e
9L64DpdfhH8llFjz5Ks2v1jpfukFj0xpAPI5HyQE2zLLdFvbiCc743eZt4YB
5N5EYirWN2yrbMEptTbBNn5GWLepgbluV+QpJObna6CJL3pmPTWx5jsj3uqs
YanTB+uDrg17Ac9WiiO1CGs0Ug/xYvUYak4wTb8pc1w08k1ktd/KH2lOWdyv
UB9Ezv6T5HfMB8q7WU0SM3QEKnVTqoncNAdB4Iwd1cLOofiIaW4jEoK+zFz+
tbfylTKEuW8tK+BoGZTucjj/On9zREWTGFCq/EzTB4BgwuO5uirk6fuNATcM
QH5WYrQYvbI7Bab4y4U4kFzf7VBC9+Pw4H7tk74OFbVxF0aEV2HvGkSc3T7p
l93RdGoG80mPCTg3IGo1UGwRJxb4BjH49Wv8kblx1PjBH7Gl7eSXtN8yRT5L
RfsDOCPbs7vyBCNpx8ukWTKqHAngCbhYND5/cOK/jPwXPkG2Y5I36X96/TKk
iE2B3sRqRJAIsFKxNVlDZYtRVjdVM/c9zRhYQ1ZpiO9IXqphAtAri94P2UIh
iFqkQRNDIo6DMIrZ9dAuAUkOguBLEZJkL0El9FD8NM0MYGzNuL8ZUpEQBm5D
e9kEmkoJwopjYTqhCzVrIyKGJFU/mQ0deSx/MQmoOw18emmzq1gO5YWmun2Y
FlNsbLLzykv6rCLDS1OqxfTBrbRl0PcjG+7SacuFtzx9wcWstRJrjA9E9X6a
y5Wa6lqSJbB5i6oiVG9zK+k4E1zTECQljPx5z/5V7C4aEtlbW8S8BqaRB1R3
W1jcfA64r3ZO15JR50UpL4+g4U3GDFrIZXGs5Nf0rA9dG567R+W/WQqql/2b
turVTi8N1HmXNQiipucFFnu7IAKrPmwXh1luoL6t7QV4NIHo900iORanxA7T
/xUW3HNmX6j3CICtsrW0CHKHeK0HqAh4sbc8moj+aDKrH5Ezhsilh4nnPshD
IVPGbMi3i+cVQVaRFE0wdC9uCFioKkgfoZ/K1SYI1gLwPSgXaBcUMXilSDj4
iafO3+U//a+mwNoE8KtZkvhFebyJAxnQ1nq6ZjixwvnXK2586DZpEkqjfChn
A/aKGhx8IroRYeO6rftjU76LFPnydlcKYiEZyYAl7MlYT7Bmb9tG8oa9Vbvd
sIo8LjSeHMjF0OffUOASd6RYY+T0D78y51NeFeOKgY+VFkdrzJN2Ko/ZH3s6
T6TuOZ+2hVaPE9p7zGj5YFP4inczdZHZaaSU2BnSDolZcBsZyypDfjN0ao/z
/CTcC3L/0Mk72ThVHQRbX/JT4O22Vev61C9OmTYouR7F4oW875HOSYbmYyHY
eOY5IVFkUaZUyVlX33LosmAx7dxOt2kqs5UN2DAanvdWXoV4hYo/2LdPcf7M
ZTw0Bzt69PDtcY+egFqPZd3AAtCGMGnjc5aPRcAjVcdrGq7rcM6xcbg/YJiH
QZTZhx+F0mZHtkeHS05jr84/KS6KjGHuzSdGKObBI5RXNdM/fk9QwqJOlwSN
1V8GCGMYTqOLfaO/8vkTR7P38ez+RbeIonzD/LEG8qzQYm+im/LZOl0W2syu
jD8HMDRnPZU4zACUiIZPFf5yNjaQ/wjg0tzQ9Hx4LRdQPd7/MANFY2vwj6qz
qhM/z2pw84y6F1jfi4NNqVm8U9iyt/pRJ3gouYNqMaEiNeL2OfuMWVPP6lZZ
IMuObCV6w4smqJ64y5Q8L5P52OW9dd4HCuCIvjGpHhgYiSPpWJ2X1SWaCVDn
YX4zaFjejaeLH7XOu/+iyN0Vu+cAhlYEI8HpifGGpxkTonhgBzlusiOAcb5v
Skxs/WUK2SWDU90ToYA6yQDMlr8X+Ad9t4tgmDBU9Wcr/2zRIIl3CXqXgH8b
aY6fzcTVgI5VAqQqYoynBvKgmlIisUgBQuC6bNLuqkAiz/+ftMFTQmBeEplJ
crxTWEo1rNzTc3kxCBBRED4BH/pllYUkMz/LvvOMy5+Jjs/XaiC19T8K7mqv
bKH+l1nmAZbI1OIOkQfqWNG42Kem0KluXWJGEqMjtNkT0bkugMaxELl8i15g
3lL4F7pzvihrwZWbsuZOsMfYA82xqIbjxHAIlRgYbT970vHt7RBHVC95G/2j
GtQzUrTKnFn/tQuLZNCfIe5SwqQXFHancZDGCPss+Rm30dp86hdivknvGzQH
D3qiaI4Krpsj36LTbg8XW5zMNgNwVCscmCRKBDNgUWf0koGx+fAJyULuJBlo
PI9BVDuibmjztw7l1O1Jt7CTeE3nn3rthQp5FzxUEaG92IYYj8mzUSqmO2pD
lHjRsiWWQdNw9vuCyqd8hbyn7fLLCwkeR9r4i8riEYUWz8VFQdtVdlsebZs4
upvY4HLI/b3eHgAQcEt6J0+fuOnFkJ0KCkqC5/4Fla3sWE7Xy2FqSgsd3zWe
V6PzKHdPhNG/CY7Yfg2qYPmDwUpAp+GW6EAapoRn+wWtm5EP1i9glk76tZ4l
h6Zw0wBBTOnqMDurDXoQDBDBjQcQ3uXaGOTzP81a0IRHUnqcQyuJsle1SwCl
pwcRTzDYHdfifu6vrVTfmq4QhXPDBQ4/spKuY8a/D/FxTPLfz0K0BmclkR41
tmqaofhcCZTkJlD8IOQ72sYVcN0xkHUgJSy/a+hvMLyOMFF7GD99uW4eNcbF
7JXZvP4MVhbGpBKEC6C3Rr6GaOAYHwNpoTo8WeRO5YzIuriS5/N13ZOeUDav
kzz0pCdXqOvnEm86SgkNJv7X1r/y/a53Q9CQKVPGv9gpwAkfTY2AU/ee+Ahg
tMmSA5G+CzfH2QGwlTR7TUjozxGEsOY/BwzSmwV4Le1iBA8flp28ffsMsRu3
Y288qsND9DSnvfRd0+FCyA4YqJpN0bNF3QyVZ2uLc3mh+A81Aku0ThvdA6ZT
loGHQWN+QuC3ySoJo2QIJXQe8YLyY0dCiduNnnw98PbkkgGDDMwPCFClDwzO
dWPDBCSR6J1qqKAC9Dxl/GD1RzY//Won4r3782zrlV1JWCqPQdPe6ab6CrMd
SD5MaLmR5SapRp4UtOgqu+kuAqy49HzrYXvcKNXTFNC+MBeKeAT33ex+JTdB
fJEqiadZE/nJlsiSifuPAcUUxxOXNY1Ih84E7tDqEbMYkEUlJupo3/PMtu5r
KpnKC03/Q/P29oTUb5wrQizT+S6Gqr7njOo85xLOrK2btXLlV1PN8inT4Tec
L2+JRjSe4DhINc1tqwUmxmBBuW2xkmpRgmkJw6977ANHQX7VrcA7yPTup8gp
2WhwTV1BJLbxZZw52sSCUEONOtguqD3CDRA6yd/PDLuUZjF9QufpCnojMWHE
5H7b9rX+cFni+zlm6ip3OT2zTpmOZilzQbxN4wZOO/4hbsrZRBB9Pu9kkJuA
tv3K+M3oa7csTybVUeGlhSR1EkKortU+L4S3pk6BTJeIBJ7f9LuST2b0BmXC
VTGMAv8NzH3II7s8WzMixZbDRefSA1bBM04v2vcuwrLORfQ3RBFNOjVytjlZ
uJZqjXE/B9R4/7cBHUumL2WzLIo8s24qPbtRUcbRt2Ri5ROOAvZrUkwkZOsv
k385LSJKSzcSezPmQXpIVNDFRabutcChVMVmq9/eOIsSZ8e8LYM29PQ4ftKQ
TeKsu8hEnHI8Dg9ZI2cyFPGbjNRdixPH3++MipMb/WOCs6UrS/bF1SkCAh7h
sDmj8+VctJcdrbSS53WJhcHpsCElqD+pyRIKEi46Uvd6mnlxSmCJuwE2+fp7
kAeEdfcqRYM6WGYWGvvcJ4kd0rywXWo+UhrU9AqQBps+ZlUo8KsTtTrOjF+q
/RaVxtwfJAyl8KRoivuCvySGRaTBPorvhZKddTart7XusMdx5+EEkkEHgElH
+Id3e8gm4/cSJkuiWjs8AP4PJlnvm6Qewx3zKLa9Mjge7ajqY2UjR3KW9cAn
Ws1AsUuocGirwZvEr6o3DoEiC0cMKYCbZhi+RbVCp4gCJo4tauUJHonMHNB+
5R9xAbBCO93vIR6pGpMRKISUKsCfy3p4R6mNHhs8NVmwexQRZc3RUvQqjxu1
8CGNP0UKyou2b6fHg0MyhmV7GPp3Yhwa8jt4uHS6vjbwGfw4gJ4DZbSig4Ux
Gou5y0taQ0+uucYRm6UmoThI7MaoQr9LxAH31Qd3fqhVZ/XToDPsj80jk7Ci
Kp3BaO3yGBk75ZM8y6WxPX++04cXPwpr8YwEU1VGYyc657s+80LUsjy+4Uvf
NGeg3JxUPCa6+v+6Vzt7MXFaJac7f4sWAuwFfzsHEeNUzaP2E/FJlgqJrghS
+dwJIKUU511YXNJ5lZHDmWZpNAl5IR+iem3hd8FNxA3TwVxW0F3EXv9YxMDj
+bQ7APQyddaFQvphd6Uzuyn9E8cpWA8eCLq9E/d/998iDGUw5aR1mPHJ9JBE
AUzQEdGlNJFgpE1p9bhYu2JCpgj0zKUQDzEJB3WAoiZRbJS6fh46x9pIT7il
4babJ7r8HfWqnl1vY4KnCUO3Dt4ukoUYTJmEFB2DdMewQ3yztseMEE4+ZAaN
O4fpYYlqp/QO51deNPK/qgXrxyRAWf5amr+bsAqhfLibiCPJE5iR3v6FIHq1
EkTSHzGnkCb+CQ8+Vb908P3osZOqFIpuSoWtaF4oyxC3Q6OcpwJUoczKXudO
YJL3r2iApsBRqdVd892RQml+YAQrEZWBNTBW7PxFuMlGzHY/BrlAKNrY7V4+
0CiAgD1KvFx1Qu8MFngcYw+n9Ox/9F6TawKOvbgIVb5ASC4ry2GOqLiOnRvp
pSgATxS5fArKaJIc7xSwujfl0PDzOeBh51/NtGVbgfCdztt3Z25e9y/9izpE
Q0bbfv7mrVcJt5+1xvEro8FRe+SH7kGyg3hEswJnsrRDgbDdlEpcTK52EVGg
GqlW4WMETWiojypEdKfEiItXmdsB9jUWjfkf2kZLK7+wbZZUG06ysUhVF+/p
zKwWgj1VUXkI8MAIDwl8zA/WNym16I5wnF1Yz1bYbTFsN3u482ifvO95l2Co
jzE/W/PpSdwjUQoSrUQ33YhVRRO62blItDNY+jyC/hs6SljztCKVLnjjsNVm
45pxEuD8f4ZhIM4G/lA/1JkBric9RIvjG6w8+r5E1o8ezhiddiwXBulg2CAn
0paW+ZpqmNM9CEsFJZCxmDOwVx03k2qVu2/e/fz9RGZU1keEqp5upD21ZQvI
c9+nDqClPMZ7BlEDRn0EZYtp+Raincveywa953sEtRQXe5Tyk4QX631Hg1Fu
o1RO8KvFG6/EA/Qd9evjbAGeL2qZkIb55+iyi/QXkcST6BfzRz3cFmBeZ7+N
RPQb+7iqyxDdspZ4gpZKFUYGxVUEIuvOj6NvwXDQHKTZxdOtDj4N9rAAbC+J
cBjACSP39x+yirUPYpTfZOhSoaguOJFKz91ivakQ4s355u+NFmwAj8VGqFm1
hQGLDsxukHQ899iQqN1jAHHC2Rlcrd5juWrADlZO6t0iY6rQbjfdHX0qIEDV
6Yx7+7+JwRKjXQWfpxN1aNlByZZcxFjrI0EwQ6us5xyCFVhu/JXL2R25s12J
RX7VETvkffxkUuk/rct+kDLtnXGXcoCC1oGx3JVB/mkzCudv7e/mgQAAT1Pw
eNuEIjei45THgA7aDL3tgnzEYu3jUyzS1qV+QGtS1ChgfF0CXaphCQdX1r3A
X1UqmrJ8MZpScDaXc8WJHPuRMgIwkN2Theetz8QxEwwYjWwVtLwzTZXt/7/Q
urJmkZSqzp1kt5JHnaF+52JjZlu1EdTQdwlOgNl75kKRZjRMThf+ZGejjvP6
XeAINo5SSFW5id7JUMCCkSiMG/zlwlm4ZSJP6PDR3eU6GGBA1163OgFfL567
/buulqaadAl0G4XvH2OI2MPl5wehRJctv/1uqI5riGiG2YOIAAiMmNJ73tLv
qWainfIEWYo+wTDkupWfGRw+RMJKieLAqgmPQH5gkknxs/HqpfqvJx9vMhCG
Y0n1gW451dKmXOBtg6SBxbjU7jqKItXur63H1XVBsnWUdmUZVByQkSYD0YFc
ID5OQMCIitLhfwSApRtgccoZyrm/ET7+W2LIQ4tJE3aEhgl6TaK+/xxdE1Fh
3zXg/L6adsT9yqqQWZpvKznDEIoHKPbNGT3hh6SFVUawXSw35vgK/eU6ZC6u
QHonLRij41eZsyV6oeATmQOEsQWkiJj3nv5ZD/pSv6ERXy/s/CxPoXs2n2+G
XaESp6GQroQ5DT93T0952HvdrF3MsOcw9eH/x0iL0xdPVCiUh1G7qMGG8zeo
BdGXT/7u1hAbqSycFaYyIxRMnzfJK6f7JToP+y50KBoEwt+lzhaWA5quY0qc
uAg1FbIQxjUIOoumaxff/XNlm957Y1jk6/tu9Z+WI3/7gDokecIxkBldNIwS
ergRQVHaMfeEk/Sv+ZfP/OXSshKMIksedA/pizr+P76hGKnxJm0wGdTu+YuW
+ZvpF7fk6/Sbf5fc2ApbqXbCyNkXPvjLEvb+dCq17RqadrVoypbkGODpGuDa
UbAy7deZ1dwuskenb1zOmBts0NbmF4SSwKqfPdNYuajcC1mTpegDtWOEfLHl
HQ2yWRIKetyu48YTMuIxdrd+AdYf+HXqlMTwewlQcAKYYgCKZaTUKNdWt5uW
zjEbG/OB59+FxDbvSwpKOeqAgT2PgCYDZ3Zfjl4RjjIhnaU6uxMGZ8aj/sr/
G/qnQXwnairBcdQ7CtwjLMK7K+XOLjKs1Kyw4e8CTSFVYkffQ64ihOnIgY1h
jH5NV/g9hZbIrkjGsjtThcxpRkFaNyxCz6hNATWjfH+J+hKX0289wGo7t9u8
uML3xv+LCUrAl2kHxmPIpVi2dtSItV5ZreMWgMZIUlBq/S2EOsqyGMxwmVRm
wkvnJ+Oj+T2E1WRIorr7j3frQbJWr4FXJWC0/oGEFXdDTbrIiDhDfQBteHg7
whz2vtgQYimOvTF6aTWxpOrpiwb8o1jSE6p5Ntm6APC6iGjDskSOvrGHNNVZ
s+rBmQ0KDaWsuODv70tuFyKl5jPNJpSEqEswXVrWUjYYXe0K8NHk+KPIYU6+
zQ9B5gH59DG0WqFdXxbTVAjSN5Mu9XV9FSQn0JgqtJzpg2cNkrgKpVWlF8oq
Yvo8ErXYGcCjYnanA5Kxh4Wv5Vez7779RmuoNvkG6yAdfvpmrgxSWcaggNpK
ahAHo+bQEo2QwUzg//QlprV6Cq1wcQFIrFjnU9/SHjD/O3OJPTTxSPkX0Ona
PQvwtHL4AOy1wMD8SdfqebytsEpGJrqEpUmKgVKwjT/M6DiFCndNmv2R7q/Q
RkdtBr3Xyk845ZWXr6JERoU6t4cLJ3X8sXYuoXbfMNRUR13sF/vjVoZUNZtr
9wqsH9fPxYo/T6cd7lWq0WTng0BqDNTYnjJPeNwd8SqQf5ZFuQVtPz9Vo3Yx
cjBzfxPNE3gc4FcZZG5mQS3eY/A4lQLjeKjUt/EdlUmwYRvYKyYilZ9rI9HT
1u/YmM6AnO++gFDjsq1QGWZmgP2Rwr3WcZ9rW9gND9t+QCDC2TJmQxdE6nbX
KY4uOomuUsNuL95ROv5rqxG1zeGSTZJIx+AfeLMc3uSB2UL36HYEjet8KK+E
wGSnlOFRwDE/xE6X+cEydTcUqmDwBIIKHuRHeCNodoyas1XHe+gTVn/p+RZ3
3tuJ8BifRCI8qtlIuMzwExhABoTIjRytcvSFGnF/IEmUln2XBQVqIOANGpDj
fBYjOEhbaXFU9yJjA8u6fafJzLqA6xWGNuDNWPNGXVYfEgd5F7rJySqO9nG0
ZWqjOGHs48d7QiYx//7zLqzSMZY1myQaEdtwU8cqAb9upJZLiUCL4lXvf4la
Vpxh571s+7RAq8/F80ukgDGkLbgVZRGBSfO4lyoZtavYcao4RZsnlLZEACSx
00EQ3RVRWLXUQmV4bCketgBkv4nzGvdJgKKVK9cRGdavrQsVaiD8GmYugGpe
WebwED74OS/WA045GyQpcpFSztSBdDdylZCgywE/4CJuWg5xCBZq/UcLTIvF
DmXCjHcuF2CZmLiQ0nrHdXbQObMPhOm69OhnDhGZQW+50xpjCR5r0uMkFmvi
llXnafY+ZcT6vdzUhMbtHeUuulQUSSUn5lZ+126VrCTAtrB/UVks8i3M3Qok
6dNhqjEJfrPJa1irNfrxd5p5BPeRGEru5kWx9wDTwFvOoB4ixZbaYfH5OALz
m64byf0qR0o2jdFE7YPiQs4vGAxxQKXO+oY5Ep+JqynDuDxrf/9uCjp39naE
Cre5p3bBlEl6TJVbc3mQubCanKk+AQOtVxGv1Nb4ZrMCGLD3ruQ4mpftO8CS
QjDa28LAkWOIcIn72vEk2vAHSnoD4f8T1fqdGULqO6kC0pbCXnrhjlgV7mHu
vWkGdqdESOwWLonNbjYeIaXQgVbfBKFGiUUYlLbmHzyp6HD55DqlsrjYKYwr
bQGB1sqmqRuINTaQZan59AN1qSOZ+gMr90EGLrLmYh2C7aoJwqPQn211h6pV
jqi/j4nxh0pcbJwPM57WdKYR+nKIiMCoHBtjjtd9PM7d+Q279GrVp3DYF02i
wte/mte6GimWMiYmR46sr2R5fw2guOnZ8/7lHPkOUA05ORGPwhoBEceXcj4N
1A8Qf9NNV1LWWGBdesTdOdIA4ll2itzGPf4A2RdT3LqRmFS1H9937mewquUj
MyDqpyVq55lIMtQaRPZKJSZBkK/F1o6fEICA2HNU1bUcokaWoYjqV+hwfArO
phDIPNOhn84zqdGSzt/JJNNuKOMt0Lmm8qtGAsGJsgQJT3ZxnmhHAUhkJPy3
CcIkA3YIHf2NXVISrNacw4yhpnPSdarZ7eg1nMeDGYKhO9ziP8M1CQyRf3Pj
D/FORnXe0gweS2WSBAogOeKE6djvNYHApKlbPbYxtfpfJhATtOfqjkTMXJEQ
jOFr8MjYVxlsAUxdsNqq3oTJ1a+BUnCJaI4sKDdQqzbmIaCYklHyWEQEMIuW
Q3HLT8gYtyKP1BvTFVBRKJMQlcpVsiA+AIEHXDvodMMzxTmMIuN7uSbWoH/B
wiG2HMpOljw/Xkaq/F7aijWj7WGhJtpQ3PbhZl7ltj06uSo+2uZxD4heX3Cq
f6EH3S1ulw8GveGvP2VQdf5KdzVma/SISw9hoxX1HX14BkCb4crlDYkABpRh
YxaASIFTjodASELHWX924NyI1wP30WJ4MxJch0JkLixYqKXmR9YIOBLnO3LM
Ec6V6mUwqNSuvavSYNTqkPFQb2cAzg93Wu57fZ4kfkK+wa1h7hSj9VJiiimd
u4BO+0NHPkKWSIIY1VauegiyDLRVK/18K6nV2A195gkiOvggdOSCOPJlToOZ
OImz31K1X6poZedufjd1rRpk5agYE5f3G/YsGjgOJr7JuJ5jeo+Y4e/daezh
/j6r+fee0/WHusOnDXUgx9jqSRo9K+BKvryEgh/IjTHqX2ATOzYWPDs3JPdI
d2yZIma+CjFinlLfr4cbKUjVcqU7Qjx8xVA1UwTKZke5sdXTzB4AkWiZR6vk
ZBusLVEqCZr9K8qsE9KU9uMJqTu+MyzTSepSLX7rtjMYLOmumgOrvK/3YtD9
P7+K913fir6mAsEPWtguHx47EgIjt2QtKcmGh/zyRZdz1RDrPuI6KQz/RWls
MH1MLPCLwRolejdN2EhG+8Yi1jj248YcEkRjHy+P9ty5uM79SgV6/hGCF6Cq
J7qtq7hHcnynI0y29YKRBWPus3V9OAvgVyvWGJIEFamioIWW5tDeP6+uGec5
n2jz3ZFWARCyqFbdi252uNE9jWROn+GPpsOvNhsDXHNyEOLnm4kQQ3cP+oet
gYWxxXdiQZTh/1Sc0aNXxtlHK5CIoGEaeK8l7fsotjKrsaxMHQ0lBuRh3X69
vYJLx+XOZVsePpcXhlBc6rbGAUlWIoLCWFa1NfxL67+7TwzBfqBSozB0FX6w
38fmqjxza5GJMd451IGiXH6XwGZncKg6jKD+qo+dEkMFgQUaDwULnWhOyNw1
eoKPZqqKf2ivhpsGDaUyKFPr4tjl9PVFA6+b4hqnd3b1o7YSf1K8EoIvC6hS
yoZ+OSZzSOepJSmYW3qatTCtRGrhZ8CQJ009w4OWc16+YLTKf26Phpgy+Mvo
dOdqL3Bk3pVUozOf4Y4i2yo6gcdBqndxhsgLCXaf7m3e0oXO7bFUYQkv6BMR
c32hyrlF/Uf9bAArGlCjy6R5H8pxtBrpKH1QvpJU1Yl95rWl454ozPQ2YfdK
cXe1GsCrMYwxGu6E9ViBCxmQ1/AlR3SNnE3Hqi1f7w1eXht+PYI9gPbDOwJl
CdBlKDASJLaBIVVrpvY8gDuoSMjcpKiWHMyhrUuKqMz4qgXo44/81CWN2OJf
vefQgmv6ijuhwlKJu+ktxrIm71pXj35Gg1kOomnoM0iL37u5Rmw/Tt+081GS
iN+X+SG8Kt+32pqoPtTQyNW6DTqIJoWGxGWhu2e7EzEbGnBinJuzbpBOfVuS
aD/OLAdrkDVI0wSUFyNBhkjDLZNubC2fsIVniwgCDQbmGBppvuMWSdWMNTtd
DogQpiGVLiF7cnk1hioTD67mJrKnPwHg3sAhNw8lkfBTmbB9lITk0MjYYl1A
00A3qNrAvglof0GXxlT0ny5fzBUVtYxwyFSWIMl0xpirqeyroGTAI3SYuFCu
eza9R2vgJR1AvjoY4puqVb2FmFbhaCdWmKhUCE89uPiJmuMvR11U7MY0dQ5V
mhWjEZnUgsJPQiaeVC3E03d1BGu5/qcz097Zzx4DCq0cumQ7F/QEcTdxa00z
FVUExsbuvYVUj4dZGfH5p07WrVBJ9wnEo4E+Pc+toV1s2qYfIYYwpNQtq9wq
jCeJoa/J9RoeHgBwB9XIU80vDr3R/rLpZ7Mvobj5L3k4gHmR+hCoYgXzfKhW
bKRMFVYfwRuSlsBMb70UsvHKCBb9PJrmzmCqUXaGzZXPbTx2rR1cymcCCKOs
c4r1NmdUHRUOc5SUVQq4YncAbaIfO6gzVmFBqyx28NLyKt9yGOOLOx8G5hro
zLW54BG9fi59lX9fDkTHHbjEVkVpgz9Ow+Xzqk/ezMoukOAs9LU4VKbKPgId
WNGl0HOW2neMqCIMeBC1YajfFOYIVFH0nZ4PMRb/wDPwBPR5belXmgsdtm8X
lvvW6979bfJAZoyQnaLfAY1lx/ZFbDSL9r7PIGUwGxzEM3PcdhSVBo+qbs83
bEO0vXsMiCLHApampFxLnBM8pQhuHnyjyITpZ04I/FEVoPObrAdzHMkKOYr9
hz+rL/1LgxuxJiMkQsOXRUyX5DbfKSMO6+v4iVGzWd04A29wU9/8Il9ceYBP
zf2W58W/y+gRx0b41SBl+d7w/b2fwgYHxNI9RWijFWzhyvBqfezqxQQStQP3
o2QR5MeqP2mfAmx9BzZBWSoO01zWR0X7zk7wLiOPYvLKq0dnVh0ev3siwxyC
dXxm/wDWlrGSnAHnObyt9HY+WQKFr6LxR765+X62ghx9ogL4eWHE7Zu/xlEu
vamp9DRRYoMjAip9KPcU7l4J8I2OqZXWSl3E0nnf5Oez2O48wF/piN90X7C4
yRyGEgiO+77NuEs7/ycOrnAGSSujpY54xvEgFXiU2/7p065kkpxoi0Z46gev
YvoUZhK0i04iLJYT5QmmPc5m1KEZMq+kRb7FkPA5uabQjYJYw1u20bXhNvx5
//I9tFLpjiCw+AF6m4m9ny/bQbrbFBBbH4F6wnr2kmEH9Jyq4UYUOgFO1Nj/
B6H+rXQGfw20UGcD60eN9Y4TiQxQpv/96gs37tTgq3juStdMCpqC0AmYN80E
MXolx3Fo5B70VTNmrLz8EjgPYOXJ93CMZ6ZV6PjYLbdhRiUPM/TrFa4wQC13
kQ9sSXQif8xSAsBm3kNNwz/9rfJCJ/+CjElf6RuT7qJodM86m6D0po7fbGsE
s43N/aDv5GLPBc/EJ3dH5ydMhn2vsWJknU7IDV8jx6NB2Qz2bPGezugX5MMq
znLQzUU1O4cbz6Sy1lv4RitAZDH825J1g7YAiX+FYduu6yguJT14KYLqFB20
o6cdAKGABX50UBSpUS3iVtceMHEiPATtXOkxu61p86vj6XN8zXgbB0EHNjZX
OVEFWbWWmoVXwiIogNCYJfFxcfu9IJJpniPfyY5OcUSl9VvR4bKDVAVl4JGh
E10szURmF6XiejABULo06L+6qyrwFpj2uPZtG/8Fv8qBnOShJ3s0jUeqLUxS
iWqbzQR8T9TxzP2bGbizxumY/wRLhCUierCkpVqQ3y82Xxb8atrgEfIYqVBb
eXFauI65us/vYH7mK7Gh+M7ruV8dphW2Fc5DG/I7TMC0Y5khSONWvXW/XifI
lTyxnZf6n9bugr7AWqQRzggPJjj92HGw8bG1waYnOx9itbZe+2Znw0/G9Mr/
Hcf/2T7tSxmRtfQhshWS7ZnIS2nLUoPfzv59dRBSI8jAtd4RBRcmHV2/BOzH
kzUEg30gerqXoi51pEenGKbhx8k0VTXOzioqXfVJ+BADh6OBUzj0MFMW7wQZ
CQbgizTeJbQfdKHQgLWm+g389HO7DC/f65tRR1lENWr5KY4ZHHpWFth/ss/b
S2YTJzog76iMgkzEPXdabKS1sYqJvlSrmypeoitstJ4TETmDBOk7JS2f9dVI
E4g5g0ZCjaEO0uEo4O1/GYtiqrQ4wcX7x4oNG+bBA7t84B3133RNa2snvxlc
tkFmTxUGvEr+PTziu5TTrMl7xdH0xtcsdVJ8VoVqV6PN7EYfE92Ma8RFsIYM
YMQrBpdPJ0el0tP0ONkjkC3k3JRSkJa/cCdganLIKvwgwUGmr48PGnXIno7a
AiaxCnREMHeMyulPnv3U4ceypzPBBCTJOBpZxuMllllFKw//oyUiCPu4lQRK
+LJsP8IQb4FHjuv8bIMEwfd9vKMnFcOFLYQ3YdePK1eKNj3pNhkm7tqeeBww
AyX920bAmugveUUrORI5Fi9jNtMUGoHUF6PyE7JJc6E62E+/p0SMqhetI8V4
9jy4ub8GSBy0i6Dunft6hSSXCVf9HFUh+bDXsFtopc3CFKnMoqNuXIRHIEUU
GVceOKWXUWZJNdardKjSJHdH8g/OpbCf77+w0BzbS+i3Prhdj+g3karcQ3cC
2JmvQpP0CV9JltgkWDxem9rvHxf/RAfsJKXtABFlSdf5OgJ+08fyLo+e3shM
RVuL8vpG9OPWxBnsripqLOSEJGGfj1zWS7Z21HCg+P1fO6lKttTT9wRW9flB
zkUJUMN0kdYoBIfz7YyXLVG5v4LGXkJ6JFrFjHns1XkQW0c0YeQE13KSCD5j
Z49QMn1hn4xSkDd3P5EOChTr+WBvBjXclYwfzJqyvL9xxlDB3gLpZrjTonvC
Ug2lA3Z21fgIQk8UNDdx6wfrQXLw4AEHXu+F0QbzzjbFi/JbCh5jU5ADcMdU
CygWZ4AHbp2U4H9w7SoXA8cxSy0UpHDITJdB+qKeOCG8MX/Gv0a+Coz2o7Wr
Rj7sPMk5YIBg5gN8dqmtHYYwthGuFlqM2v9W9HcTEhYrl3FXgKk9taeSSE2Z
NnSZu4EeqodXj0ss3bL9RHdvAXZcV9kwtgA9RB82xvn+qsYsXsID/VP25yu7
SoxdvybyF+65zLtHlR46NDOqyTZQvVOmgstHNLDk/I2ce1aDgFjrIBwUgqGM
h6Y0VhFJrIC8QSI1ZZQXe6ivnh1GV6gYLI1yOTFEYNaqQ75rnZGozEzXYkmf
eME7x+PN8qYNaJzpvUGaPnwD6ZUHvMjvV9kU5/gqx+ac9QxdNETUKRAfymrT
8898IITK8318qJmBoOzTWgqHGmGKlkZiYsr/ifWdDeVq7gezllLov1i3QlP/
H/d7nizLPhjfwp04VxnLUde4LlBl8jp+IdoEvOUnBWX8QaccS4Ll8YPCzIOJ
rKOMHUwpgz+bXmOtsHa4S/OdqSwJts2sqPnp0SB7fZiPz5I0Op0J0q7BRN/Y
1PUGXmhA35+jgrSD+ZpuvpayNseXd9i95okLNupozN3E5Hf6ArEisRAJ/Dq7
/ZZV+B4b7YeO86wl4NRBc0Y/DtgnTqxX4qbADVZ35Rlao3rZon5gOKN49zoh
2q58fNEQL5ewhCUEu8Ai9PBmYmuNwAI3rEaOcIFh5kaETGC5zmlzRNKwl5Cg
lBCoKvIv0e9KimBQYAYTA1tI0NR0bYFTB4vvMFLqG7GECfGILAGXGrbyjKE8
sIADD+mEmURkj3T6BlJ+wnBSqeTLaA4P+SU6uIeTs5cwGp4URFM+N/s5+Swr
cJpgXHDWZn7w9DcHENrL0I5ptJceGnVAeEltfqRTi0/9GYqs4x4QKtA28Tim
8/+44d+kTvhaSloSqqD05siOXvVJoZDZUFXjT5/qqM+8sY+Y5HhcW88UQwLQ
DnwHrf8QBNKSU1j0cX4eQmrknL3Qd4VhSfDnx/XAUa27idmVSq4xFMz+ql3C
Dy8IbkV+c1L8tvCGUmgWFBgNmHPrpzjU1UiErQWqAFnT2JY08yjJMF/xKAOn
7z3Z8BUdzIUIthuLZDeJwzV5lxqPEG5Z1VHvZ9AxX/8DbW4ZSN/dxXsU+NUL
jQBwMyqcUGve55nf7zW/WOIVRoJsXC3CVp0PNqh0WzL75p38kth6Zr/MKCs/
tXEnmTsAktAas1EYiX00YUOsQ6tPJppFPmKJwbW/ImbBiPjxGqueNQhWt7c7
o4on3yZK6cfgPCF4LoBpiacQ1+aHO7beAIG/mMDdQsHZM2FC60DmUD/ik2Rf
HPqfP1HoK/ZHDgC7iRuR2qXJRK+WBSAvZtzpDZ52/5VH/yAJlG0libbjpQbl
B8/AcsZ8z9/qxnUinhfMXGbhu/AEM8Xi03Ege7oeyCIH3l4Lo8Xck8oR8wuZ
mvb0Ozbp3p5CxWzZNcjYzB0BAdKk37jbd5TJoNKnq5bS40ewp867y8Ovmxnm
yBT2v/g7mSVEhFAxUjh9YNnml4ybwltwfhW/klkaKZm9BSfuwWu+qNgNwqFv
Rp5Dpz0Kq5o7ueJ3AEgMwsPfhIxCNDzKlWODbseHxrGA38ZPhn5VgxedDXGn
DlyTLWAncIfbe9Avlk3P+TavFMI858oyeLGtOY4DMVqbZ3ysAZ/kCJAYUsnB
TQZgajC+PKPym4e5nzaX07u3bsDh78UrAAqmLGMrbLQ1vplfOQ5By8l9/CCZ
Ap6OwsbZoF30T02QJsVg3hXoSRsfNoefA0tySXBVwlSETmpVbQLqYbreJTGx
pfLX9Gab2XEDLdi8H7a6qaEle1tOe5mxaIdCgupp69UWGplpfQoVf1lrbDAn
rOrw8lYu9A4EqNAGb+N9FebkuP790RcrJyw334LspinZJa2m7xS5lFksmGEk
1b2RWWBLl7jmNFq5FwvT770Funk61xI/jthUDWBmr0CPdONKPv/+IrlB+Wow
/5cvaaLW/CAj7mONZnLtg0y9W5NDqVJKj46sbfliP/Pce2+NvpbRGwJ5UigM
zgaULiK5QSZ4VTV2z5S5UwsaiGTHL0qSgKBnz3syH9orqsOOP3qf8G2YRgc4
HHvineoQjccL3xUcVQZ09dbf+hSM0LoSRnGd2OpDp+J+O/5XnUsDNAxDe+b0
hM53alK/MU5UFs3f4xjxA8PeTsrO4V9r711R7LjZ+NqaNSww7MK/+UOlbdfF
o/iQtXxsHb4riX7Rpfy3J4KayNMlmxkSes5Q2iplh5d3wqqyqQVwv7Wjec4f
nG9Cao4p1sWC52a7DG8IXJePwpsMgrVMB/Z9NNpAntVlZiuMq5k/APRBwucF
zx8ILveMyvcwcJ0i2wH1vEFed5g2KbsdfJjZEcDVmn4rSA4o6cCJeHRFe2vh
50mBIDlimP8CbiHc43mTUD6tSrKWQ6qucee5fVcEluW4mjS5krkT2ZDaxp3X
AfYKBaLJVkAWe6eWxT67PUhsqUS9o9ezeXMuN1TepL6fNYEHHdx0kCDn2ULw
C/Qc6KlLaXQHsj+Xp3iepoK/YTbrggIFiXESJawa2WRPbulKJCrXfeAqeaal
Q2LjqIeN7dcDhzuJs8BPW2d6d9RAeVMIqBbbjD/1wXMr5W6rzq+CDqhfxink
M3CvQiD45+CfMwbvJ8K4JWxjKdXny06aHVVByfXJbKvaChcxXcCDqEW3GqU2
SPq/y5qiMSpjvzleJLG7EJoBO75+DEQ0sNtUjprrB8KCV6Z2DHMAVx7TIBTk
mCvDW4tpgcIyiCVF/qiaw7P1Q4HXvgPlzduq/GtL90vBhm4VMJveMvt3cKME
QhMEvT/qxcIjViKmFzH+QJzbY5G7cncS5CMeP6VToX1BIbVCnatUKmhh1PbM
GgRHaLA6Es22wvwjpdXGljm4BZ4PwlvSi0uf1jNjSbhRIscA6hy93JkFK+3y
tG4csSRCTX1aAuweF1fkd2whoZ9b2KxuvMAs8sZgj5GMlt08p41pChgtrOPF
ASbLFBF68Kl37AsTety9TngQETPimBxv+KtiPgOVAEfQHZ3e023U4xehHGhb
G8vzOSP9VT40FQFOLFh8ccRsHv8skziHhc8JhGcSerOYgoHrnlM+AF1f7GiH
wA55B4jzvRjHhhUjqLZNDmlu7hGBhndWET/buIwj0Y+2yp0jaIjAfYrzSH5l
CmYRUzaElF35ws0McTUzz80Xne4XTm7pRq2LhG0LLNiU9qe2Xx+2ImpZezJq
eZKdg7FzPucJM610IOvxESMloJoTu2E0sHeP4VfVGz8OYKsgWR9F8UH/DYfu
HE3j864XUDtFQUGQV+67/KR7QOoqTMEY+Ac4q7e3kQWSjqxBOLuoX5Gatfw7
LGRUmC37YAX6LtefV9wKuWEn1/zWas1+9eJzy0234fJhpsQqVzHS8LZ5mF72
gnoL2wuvD98aFt+OET3MgU1CQfgcJe1AQ6oraT2q6KvqaS6AIbW0LW+AiY0X
Mk+4zxMgm9CN5hGhUGH1AUHH86EmSBmyLJ1QNwk8mnpq2c5Yy5xKlRJYvkUY
Gtkkae9kx9YSSmGR50zPzUdWIosQrvtTFFKua2O0quxTNYqbAUbxX9OMPMZN
TYt/SJOMmguvXRk04CXHWX+nz2ovpoGJmkQwoMFy2zYv1oiRWAawvGoou4Ja
UoZctPpa7kmt3E8hGK9yDybDiqiHXpv6J9XUHNHBiSiLT1A+EfyAtjWuWcvA
ehtjmW7O+7nke3GdcF0yaTC8VaNW+lgGO+UsasO4EB48ZCYhi9zW3J0NUnEo
12BRA0/O6R8p2+BVRtY9wOeuUwE1BXh349O9XBD58EXY78xMEIhykn5Y2cOt
CSNd/PcltLiGQOZNnGb7It9swAecJ3J0fpn5AOTQpBxVWy4FkdOftNj4FKMZ
5bg7pUX2NV+Cc4Y9GphaZAB2xITekVCguZyebYA1IuXGCM2UrRb1UXG0SuZX
/1p51dGjLIFUSHkMJyu9lwLyz6h4dO2xhENPlChVtgnEZYElv3m5GtOlqkrO
CPNkWjCltNvuKH7pD6ItAABER7lgdwHgWGTzetpu8tfbrZTjYDcpGw8dy7Jo
rCvmrRceU36WmKng0Z9CWuo3N9ffbN63pPc+t/luoUCx7XLIsm9rSsPZhukf
1PIOzWQRJ5jrlt4Agkl/URRYjjnBIjwKjoyQeaHr0kNmpRkf8NTLelMjfjQS
N0MnfN8XNcGmJ5awmBaISGV1vOOPiIO9/i/Hh/xu+hKU/fgjFZG5VDejUCl9
hFSLIDASDt/MsnpfSLR2FkKzKT9TJVqoa+ciEqd6A3z6nEl460uF4n+w0mXq
OkfFOmyEjPztsw985hO62wBN36xFyHLyzLUp/mCiFPz1VHogOl8dOeDipB/T
ZNtu8ighSEgEIIunSiqqTD2ZUnwpUmiO/r3ue7cyxN6o0LlSLK10vXP+UCUe
jFH3ZDfhhvX2hAsfjXHwR9cldiskq7Q6b0vItjTbkpPOi9GJ93eHZlWiHIqN
NCGuF/elD3K5fZAS4BwRY3p0p+sSLhK+A8R5ghr6opFdoIyHQk9kluF3ALoi
wgiSQoAf4GrqcCHeFbv8EUyFNvZmZX2mJa0/KqjPil9kLI8VfTTUIpxaBlIq
q5FSE6tmt2eDsHc97+TXAOa/uRKpLsjLtzdlckVEt8KfdO5eWJ5/26yNx0nc
U3VY4EUlLNIGkj145gzEmI0j2LFUCSaIjOXmE7MT42UNzfE6qhFxAU5m7Muz
Ey5aJD6glnx5gzirhvZePMOLF06oQtG3SlnIOvD8CoOmdNaVfbuBVVcLgtsU
S86nlBE4bRBTJDCJ1XlrFculGxHX8eUaQlRHeIeVnzu/NLKvveauC6lZWDh6
ixClaVPffWFzfE+soVwpQbTbVFRXWfP0gpIPz0TfGX5pvVM3ceayAMg0cKLH
TtTPaiimp+gIJv7Bg3NUQ0qa4jlTqlXWCvL0fgJB7jEoVdModV/Ulo/73v84
cK7aJ3vIrRmqBSkZAYZNR5cuEB+sAiAahYXKQJ3fIRMQiRp0YvFnAvsjk9By
hUJjXlgBD3L83ZYxOs/jRTsEqE/x0N8C1PPzDfOvZ6Md8et5Sv2fBFWR2r98
J2zHjYARZxhTe94iZep+V2ms3kkM4ThV4Kccgd0sE80IU4sBfwQmgxLppnCT
YONxHCHUTxMNtSjPFy7jzbbW306HZjO9sPob6zYN9KTnxG4/fR/QXhV/QpzG
/CQLZ6144ya7TLJp8mRFUF3gkwpMUJVOhPsA8HQyHyjavuhrMD6cJYqJtX00
VlNh5kzmnknn7LAiOXkQSlgBcpIFgQf4NynbhrWMIqT8SWzjKMrFwrvaRZo5
k1h9tiX+vy2s13WvgXJ9H/5arIAshK50jf2712pZOWIUxQB5XMDYW+ce4ejZ
fgPFHkZw/66xNQaFiB/ThoFO2oBwz1hjjwS9ksrqeKFumI3K5c5VpSnz7PdC
ebdiJyzrj7wFKZpfh4VZjJrjXLqE/qQdRM3zHw2y2yP1ed8NrHVKNFZglytk
HC4MCXokoI/OJXXVDcd4BQfSvZveruu5Fj8cuRCUr8bvOerVMP7LCh7+ravA
KPA5HgvxhhJyGa2IUAdH80I8YZy587sd5oqeoYcAFdm3/rFveOosa4Wfmk2n
b9AkMItsl1hEUU61u6qShlAMtINU6KFz5dDT5l4fXz8tpjLTeWZIYcOTOGQy
4geGj1GMKKbpal0SK/P3BztAlye0nM30r1+adZLSex8wS+6gXuncRe/Uq9Wd
HodM1xwZnDD74cLLjrRd5NcVuCEU7bnmGFhTn9y5pwer2Py8gZwnEEcCSsRF
fe1ZUyEq2lAjRxPOaOLIYu7gMpLJbeqE2qRvISyngNm1I0anj8AHloE0NWG4
xigH8+i4wLMjx+GHskSzpOYYAHauVQasGZm37DiiEKW1hDzjHSb0R9MHgLin
gAgfphMFeoehZqELG597O0mZhu0LdnfzrqTfqRg2DJZdIsFTJd0bygLsaA2A
4Gejidyeb48iCY1Pj32sXtA4MxpWwdhJsjzm46lo8UE3JTkxaf/BXcRBQkq8
SnArUibMllEqRFq24mfAnJxLWGq4OBvugbFL3we09S2xtD8/KGGnkGg21h3k
XIHFX/eZmP09NWob+6ENNgGkPOcLixI3qB/qbP6YKBasvmgRpa/Hbzpr9Rdv
WeFZZI50bJ3BK+1gYX6Ye/rzbIAST3CJ4twYZdQPyEZdpKgOXKracHEkJEke
dVh3MEMnfEqNOCUS/iya9MtgOdOcC6gDpxbpmsHT0uZBi3FOPDhCRAErFW3C
KhYilJD0f6mVpR+znHlE8yv9TiGCs4P4hPM97+IfOwq84J1LcqOlU266qCaF
omYqUNEftwxSZV1ixfSxoomIQBKugm3LZeR8C3GGL+zYa9ULJf5fw3IsNbE9
+H33LGoqrs+bbDUdC9i8ehFjp+rxYfvfdJdS3VqneZbz5wC1X0ymXgbhzv0l
1D51cSx56IgvJQWuUTftI8fnty8uolzmwaWqVhg/ML/KImm6eQz6vBem0BJV
+cKxX4ywUAHY+7//OduuZUQ1TqBcUizwq52Yg3v1G7pE36+d5aK69xHPwT4C
kYUFMZW1cfRGgxj7qbSLMG/4NCjPnNjgYBZfh3xeqm0c50ALtmO5to+VdTbD
/Jr+EZT7xsEC79BmRCebFRoSuqB1df6ygouBhIGkPIdlCIndGIB2Mnl478BN
YX5x8rbOvx0F5Dug1TFRHAfUezEQ9xfkW2IiV34WcgR92QfEMhpLqoHDuNXK
2pJE2M0GWwhjOgIMe9Nr1W7xny4CC0TSz/tnXBc44pi3b+OLXybk/Gsy/DXH
FZ1h0HQ6e2DzUkjZyfdlsGS7Rr+vBGMwh2vJxCaPlhU5IXkqQTraaBpANuM5
sSUuYVmvU5t7YdRzpn13aHF0wgvAsKivlYvTUPCY2VujzANcdCDU4wH6GAPB
fYf6nsDwsrrXuzIoCw8GEjEFiIulCb6YJhy6sIIRK8Ny0nYGJZJ+974NIjdC
59PuWhSIzgD1aa/SorhKqYDPzhqcJxRJ7hdZMSifEYD138ehpcZNugjhfxtN
UfcEkuh0mpimvemjh+1j9ZaFetGJBIawsDYZJzvitqwtbDJ5uNvVjlNxCi88
+oWI2Wg5FGjHskMV1TTC6MHZiLf7XMKPtzzAXdZGyCUOBNS6qlTVYk6U8hVf
XHpHzbUPRW729KRy4tJvMrWsckioXJqPKabnNVqRn/WF9IK3e4BhwqpXW/78
kVOyEt8o1ZpgvbHCa3RB90HkpSd3on/cTGLuSJR4B8evRrMn2hPm6tP9xAka
oeEbrmUNLas+j9Ho+8RRdKvJxn0GVTEpiK5z3wYfpnDG/e9znBs/23JKdZSZ
/p3AG0jZtsPCQOIJfcZcRiHWpDVWcEYaPkfnqKeoWGOX5njudzJQwsOVbWgo
yfjtSWCtSFJ7yVSeKyaqI8M1Nd7kkTQQsU5lqizyuF3TGApDGgXruUlehJT/
1oBviSkDsa92OtPs/lIUT9knCj6zl2XXlTSb02M55aiXP5E7YRQDxxAmNWFU
F8gWYhfPPE7gOxihajh0AxenGP9X04KFqIEJADEq4joo5YYI7tJZJIERW9SD
0GVGotUGSqRhmwH9xRaBn0EoZlCwP6tqKrqFWevzQxPsEi9OWZFUdHtajm1A
HWxYoerb7ftQokvMUCxYIkFFSukrqvHg6v9ZKGRDWU7ui5OVjACPy3XRRvXM
OIwtn7tlv+X8qD6jaLpDxJYLzZAr2RI8D7Kgpy53Rt26KnwvWjBcsV064lnY
j+gjcoBbpFxnIiJkMHAqxvuQaHYRpB1GRPsncO0FUWpwqvyAvngM0tOsc2dM
tuLGr36SdjKD8T3bBpJYUjTOFQOpmhTh9wgAwL8HNkIJEu5FrWY0N1QqArCH
a8u/hWB/erEBFui2HNtz2lg6eUAgElJxWoJhcECGnGpwIEzYip11hsfNx5wr
Jvw/3uoV2Blkdo6HYIWDw5716SAeW+7oSz1Fpl6AZsSEqBAA8uL2HOCoxd8s
fyzeUx1ZDr+/f6oMj5WlxQ23e6WftE1kMtqHHWxS9i4NyIHxNq8MoF4X+q6D
GW/vN7Ra4N+uTIxEIhvV6YjEBAX9yImvQ+h1IyBGrNAFS4cIzPtYyEtZaT8F
U2OpiE3C9I1FBpG/7Z49QXAsfHqNmQ/cgJM0YhCBqF7bZIITqPB+krBAjKTd
6cQL49GK+dqIKwsy2nh8dA5RYmnz9e9prF0JQZcpGq5oJM4vFNUxBYui1hvp
pLvpnQ38oO5OHrOyi0FYwDvgc0FmijFBkJ6gRS8dPf4cirOV04FJ8Rm/AFjr
xEjOByVQcPIB0Cmo0r3GW00pALLy+HWl8OsTQ4iTbbeSQLhYShO6u4DkXUGE
YDKcbIl7bJPWy0gJUgVHveTHMpB0RXw7SNdDLIXlVZLYlLx4bsycEogbruhg
f1tqmLMfY5bIaplIbgA0kfWjNPRSd0QoxRORHDJ5n5y/vXoQjC9S+MxHoBHV
QrJEMtlRjvO1HdWHmbUQalZ7Gd214xN9YyJzgZLfNLQMfQL1ErS04WGdw1vE
rmIiqcv0+jKVbWVeO4bxOs3aFMzr0sRrbtAqR/2CeEbAibLFEAILdzVOarut
mxSCATsqnguMIiUqRcqRdoqiBzsaQwP/Sz+8ebOowhFCJj3pqFdiPWZ00Yo7
IqthV5NmftGufDs2QFf+o0csQnWf5L87/VoSPxcBNMXTmfXQzFd4BPpgc9We
0G3gDkuMmrrD6AYZyU7Aj2xNZlmUUj8BS3x6DpJmrGhtVqwJCsS7O5897Hk4
iCJr+UHHpXpGZWA9eIXu1iQzcQKaVg40EByiHgdIwgR0wNQaVDt2kgUK+hA/
4pp6vy656UgbhDhvw/vXfTrFGjLLUd66KK1M8HMflFhL8bQVrlOGAFMbicQ3
KI04fmD8QcPUCkFtkNPBV2EfRLWoGYn4w9oXRGcqRInBlXvNJNuTydaOcEhf
nfb1+dQi7tj3lbIZUZOrIh1FjRpO9Cv+fzDHOn25MEgrR3tukaMLWmk7S1/u
9xuxOkgCVb3OSXYmd+X5FJ/mFhgNzBz18qJF2LlGi7LnYejIETVf5s10cPVP
9U4M7zkbORGeDYNA13fhe9AljqjlXS/RI5MSF4cAxDv+7QnaNnv16Z4qUH52
6O7WIGvfEQWifLn//c2QdgOxrXETNpxeefktIpXUtEUgiL7TXck/b/NlCm6l
sL2DfWfcw5k98r6keolu+SzzpYNgWPaCTtC9npiNmJZ6VGn2nw4ronhdOSG4
L2aBJ7+CUUvxjtKjA+XeAACtAIOLG4kcigpT5L7mQ2daWdbZ9mlWRq4FMjlZ
w1WyypqVIUf78h/fKHxbudZvelB3bkIfVHTsIlbGw8Bo+XKa5ekDyyDHd9J0
Cz+eDmIsA23uaOIjcWS26mGFLN46Dn6TZV6uBEp4uqkf9FHxmyQCsR6dp4rH
6qbZALGRkqSPce15BsHJi7o0e6YGsBtK1iaQwSJPnhclIXvUjAkYIu3rIBTB
6LtxC3gWlK5JMP7+h1PQcJ7RyZaH2NYIG7o3sGhX/fWshV4z5pwRsN9EGh23
pMlgs/JrwKtPY6IJEILMgKELdtf9aCY7ZLPyaUSmLogrKPiC5HoNbbvgnzHe
zpWXumoBwGriMoAagf+4d/ybXC519WVDWw3+KR56Rhxl42E4g1+d8Rby/Aev
zR48I4kOrYg+HqlzA1/nN47vZxr9KceArg29PYJPwDpCa7wEaoh5IxEetJ4P
QmBl3iikZid6k84EWRbsYK6OUBoSgOVYhuwH64wY3fLwV5bPRz9idWGiYlFt
BKbSZoseaMcjzz550LZmjt5qkAyxV2UoMyThA3HeyrgHFRId5AuLu5GreF4V
Bmlw2C6dw8n6Kp9wkszY6S17cxrN7qSH/U0DwjfVWPMjNV7xdAyH8hiT1Z2Z
ySZQQQduoxL1IQZlUFUB/ZgNzOR0qn7sTfHJ6RKauNZlfpWKfku6VJJeLGXu
VfcdHZ2IUfXtIjLVaUB68UttAcr51730vZkGcsQfo0K5oROTDvj7HoC2/yt8
/tgHk7FcpLBF5ifHJEZBRaULCyXmJuqVvUGNBcc0+SF7o79oX5/K4VFV4OEW
kBu6GDTHkRGThG1heiRccIjhWvDKxby4JnoLK/zWo58w8nAiHcCFqJMsDxS6
aSW9JfD1u+ER2v7hCwG7tmnpBUKR/1+MEvN+WTygP/s4v0lITHtaHT8McCdc
cYXtU6tjUrTBy+I3khR+7kaWLNm3e2qf/p1EMH6xDIWjyKcvIWl2xb8FvutW
fLXJrgJbsAle/ZPT/Fo5LYwmjx52TOzee3cSMpvJcF5NlQJPX+LxkoSyyMoj
giTvKkRE9hC4Vl7FoAbTcsCA5es6SRvFf55XVDbZaBbpYtfQHsVraL2sFkNP
sh9FNKPArR8ePGJ6/pURs/H0U/l9s+VnjPbeFN5kcXHnFZccCGLFNASOrUKk
qs037n+SOTCJ80fvcDAoxiiviVQj4blCKJ7EFhDlQ1Raz8nTMQnFpTRK/oZl
ycjvLUadQRVunpX6TsxaBOqpgFzQDM4ZdvEGmXiW5ErT4YZSYjuwjlb1Dtfp
2lvhS/jfhSz5EIbNboZE8au4Y/JI9FiBg6mPgb5UrUnlIDeiSBeyCXUBGzPv
BPdfanZbZd1j/pwsmWPJ2nT6JyEEpwGeJx7hPuqDNh+2eqitcUA57FTpMuI+
jiGEhbpN4J5noa53k1NZjfUpSOX4hoeNPDKWVs+YfudPnUr03dWaG0bpJmX4
WeU1cDTcxalYHqnhC1AaxIIDIDtFTOHUS/AkhEREStJ4JICla9lBe1gBTcmg
66ScX5T2Vr3lvKYGaR6hsO0zC9+bf+G7iGU5Ddg5XWC3TPvzo9Qc7mMFDue0
wIjAYdvAoU58yjkoIHy7sEmF1UZUX5KIka5mGydDfCNkQ4RBjH0v3j1QmBem
RD2sbGuddTNQR0pD97PWxkh8BYPNphNHmG+ecSpQ8dFaJGnPqqP3qj7PntES
hGbmDdMlPos37yWkFkNwuKXju2ku1OF2Bm6qrEHnje6BAl2VMlt3MlqaNMoA
uexFduC6A21z5cyWaumwavPUfiftvMQg43bJ7vPNLFKkYt43WDFzdwo2LHhv
32zW0jYON5EIhQZhzzGnuFqnFWWtxehvP+KecsFN3aihQO8CWbph5rSrSGGg
YuwIyeB5WlsyL+634H0pWueBIvqS5d11BN2l9urTV+OZqcCa4I4fctQfGCkK
FHvoyWP1SME3pWJTUvaKFvAGvYwVP3mQpDHZUXudmYuF1gSd8TBj2EBnI72X
QB05ZEjss1jvXGNWopNwWzt5Q1gdLf4gfJ4bW7/dcQgGttR2a/Mty4Z8dpS3
3uEWO2wECSZFgD6E9TVDJEvHbGbwZ7bJt9JZvN9wzTknN8a/IQzhDWPdANle
gy4hWRS4pBl3LuMW/d3WkkS4OsNLjI9iUkOv3ysOaFl8TBMoHfLHjTZFzilv
qzFLeE9tspWm+NlQ9l/W5WkdbChEE8iDsDuSfqzFQGlJr8E8IsWe0D3mytMP
qR86+xb6gOYjHsEiDa6b+4erqyt66FwP5Z2p9m6YaCRsUWN+4DoAi9KYdbK9
QU1XY+T5sC/k1drL6jCck20Z/ojqq66XwQP8OW6UvKJJzIm8mSNQNqWQxQCs
MPr9q9qQM4FYBjON1mzNOMq9GEpMrA2jNZW2quB1N2BzcTh0YK5gFo0zQaTa
jgVTBJ0BXOgs4IBRlF11697ousixJP2ag4dusCLDfn+EwhUnc6gYfp4ffF+w
IIT7It4mjVb8ywHQbCSE4pk1jgGPV4biYriD1bz62O4pqpNVyqiB0QboacZ8
c7n+ybbVkTQpsbZBK2X31MKH8Nu9NBZW1sY5iLU/3sdm2M3o+GyydvhNEa54
B8B7Ws29psfR8f3KRCsmAu+bRurM25tZa5ARoc0IH2y2gZ3QmmJ4HO+Xf1KT
2GMH/svWxn4jnuw1mMyMdiVboJ2OtCD4HSQT4dJjJadYbpgH3agO1imKA9hC
OIbem5wyxaXv15NyeQCPpE2xChHSWuAwQuXKaAtoSyBwN3JKtCguD4MgpUzr
Rc1A08ElOyJ6wJSTRclw0CvvUQy7PlDIDVnZ0dvs+hXlHySOYv9PTGt6pvzK
Nb8tW2ICXTOq2sAM1PEyaYrSMCMk+IYHGMSuynNseqZa5HAKH3LtUBSV9LC6
Ca1DRKNIM4rPOpgei6AP3/ep995bV66cI9b6tynX3d57KHBAXfpvQOz3usa0
Sg8xVmoT7M65K0YMZRnObB/bXEU+NZ5aCrfNJXMvTkA3OgeD01j/9EVGNjPI
u5N2kV7k4ncm2te6kx/vyLIUOKauUdPVgad0QIfazw9GaKcgaLCW87x2+pP9
lrvP+fo+2Ph6OkVwbXFFDuwk9sW1jMdf6LDNNxac6WVbCpOlu2UB8S19BgDw
ecvQPvbeXu5z/HbiXhYto0mRw6F7jGWB5FnK+JYTiTIQnCBMK+WjRZCAXF6S
aNEHLQ1amCLZKNFyu70n58+s/9EsK//WLtGE4SlumGDphJKBDKuNufO4uCEg
jigiXeL3t78jtt6YaPr9FZ9GcqITvEqiJIOnd9n7oOANrZZObV0CXs8t/hbu
rxpxTIZ1JU6A7jRkUd0gawvjqr/J8v/nuGF9gTu13zvJwLLrCCW6RPc17GdV
+I5b1RwIn1p4cPlLzXv5FG+tX/ug8rspsRj7gj+BQTrc8eiGOvS4lDswYj7R
a4bhcLrJtIVxeHokpUmme8yUuLW5M9wsGgM9eoLqPPpeYEya94MtNKL0qnEn
Hwr6kNoWrs3G2v6OETEb2TBOKG04ppmqglcsnZZHpjuGG9K4nrMBBxSKcVBx
wUDCWsNWiuahbQYhBMs4CUrZSNweQM6xDGIK15tBYShMVI+y03sVKxIi9XLG
0JujgMLrl3g559AFfpocgYBIeDHbwNk6Ay1gs2zv9wJ93v4HbwXCgkOFRPof
XqRUa+c5WFYQjWoCZOdUgqyQTDeRzRY683tILpQG21ShooWbEH1RIFeO+Jmm
tzcYsv2XPioTPuZwnbkv8cIGGebpzxPhh3Kwi+YLeU5aG9GOSopnTLZTR9Oq
8zmQJ1CXkJEcdMgzW2BN2JCUHaO9UpTvvohW9GB23ieCz3B+TX54BbPhxWaJ
tj6esBdaKmNd/1rXpAochnHYCTbL7hM1tiwEsZaN9UVOXvQlj2sEX0FHQciV
Ofl552B7dazcwkav812VATeRk5Yt0WyDtqdzbbh4OfyXWGE6P/YW4k33Tns5
hzUuLXj1RS7fdkG6Ekmx4MYCDx9J6PZ8hct66h1dTxcHJholBOD6phhyWRp+
xgWsKpiUxPUVG+rI6RnL2WEBWemL/3IZT2gZJAGujdBTxjTVS36bodayrJR6
Skc77rNdXPJ7CAaBWLc1xv2R8n1WOmhWWRxcceFm+o6G9/lObNTpewNsP53l
Ygg6ghGDUUEcVENG4BninzjGC0NN1b4zno8zaikkGQC4Y0MOOkwpjFFpX9Ja
28KD40oevzNlid1ank64iB9QkO002CkWvteP4Frc3N/TUVfYZaYaBorJlagm
Omwr8qFoOkV8za+pkququal4af7120DWe4Yu6VcmpJONMJVrsialpgfTAjOh
s+LiDq1zFBrar5zjMwWHAI/XxltUEc/Sss/clbfFyxU+LIu/40gEq/L6gA65
2lMy8mae+GxN02C2y0TX8hxbpUwQsNVEvdjKERhOnZpvin+XP1n5+DiNMwZi
4JjEe8Nx5TMOs0aN2tPqBG2VqhD+6PjtwxGHAmzp2AS6M6Hkol943rLo30Ys
W/3JevqVPsRZs6S3HDzqxHkDDWIOBv67yVxPNf+RyyufQn8c+zPkZJux8Zwh
M/YkEHhYW606n8fh0+/oV5SA02QAdcHrEdGGX8oRxm5iEq+VgCHo9UvVJoFg
cWhBHvUFLHwwhmjVrySaqhvWrslEiuhZX1D3apirky1CjZSikW3PnbGanbld
9b5rylS7i6M2yTW13Yc/YfgwlKIER3ib2tlyuKI9Wdft+k1eJEXIuYjF2PuR
HRamXmbuGbQw9DXfI3Xlm9L2RuUqzQsZ7O2O2v42wCHxlKAoI9g/JAysUOlY
/0zlEF/pTp4ZnD7C/C/IRbjLCotYRDQiCsKHvIVZTmxBnIlZt+Xfx/5xZlwl
vRz98GAEJVzk4VhaZtoBryNTViNhLPH5KL9MG0t/6ucHXsbO/J8VXWQiX45N
XG6DWjDSytAjQwySqKrMR2GYdAf5SZMS3KUPAun4uy5WZL7Rx85uFZ/rJddW
xNFwvLkGM8Z5F1+8P58s2VH5JQEJcRmKX7Q6RjW8n42RUu5cr7z8pTNjB+Ns
q6jDtOX1eoih6JmmZ3W4RtmXNGctpE60ClENgZ5HSHhyt2UwJq+H58s7GhnG
hrbxITVNqGrleE2pt9vv7RU21UE4t4sA199Ia8tNq1P5l6D1o+VjjNMeA8GQ
yMEK5MdkdsfFUebqDXTupGz76ffWOGPy3IXJ8/rQcc3wZX6NfG+PtDdM/iXl
2f9F/wWXVXKlCaHGqwsP6gaKPEBFYV/Jh9aamtFRJxq/1qsLl0mC8rVcdb9o
XtirHDocdN5X9KJdyCYPNbiH2VZaVw+LvzFvwhzkNeLl+EhGiLiEL9/eAQ4R
v1TH1BDVXhoNGp5FkCpoyUo1THBZMmZwVFN/eTLR57dTP4gn/kzihd9E28pt
u0/tPrd/i9vrHoLBQIPdleRjiE8MDsWF1nZqg0jLqY7/hUIZM5b2PwJw+CI3
cUq8eOL+1pz4yQN5GMC4AjOQEu59/cYpqg9MoNgcm4bJfpoQovXinXzLJ9wh
jsuY+5UBvEn8jUCfe7xKRQobYLCJ6pBJQxoXm1SdoUEXH50DQhptH4yHPo5M
DVRQERNxsiy4p8yZAUkTjQP1oZ2qSLPPwj8FshjfN3UqK0f+Ldi5jm42WI7e
VwIl0LTvZtZViRYxICOd9Aq09TMNI9GugrUVwy+gzO1TpUB9c7KuwJ3DMfi2
6alv4XY5pur2pIYksAzTt70noSc8ZWaESdavFZ4EWdlCkoHeSgkisq5I02IP
VwYTRFZ5SDcN0gTjIs4V0T4LhAUFrz0c1xAa2CE//ZWQz36eUJzKzZ1kcvgA
eD92yxyJXhtd80gndpNEszciliAA/Fyo1Z5YfHzqVB9Lwh4y7FTircMdH+hN
Er/19B7DVRxqfpIJ3rBQcZJasKiPQuGSpvYnfpeIFBM4O6qhizGo0KKGl9Wh
AVcb9SsmKoLHDMa9oWkKdnFeZk48ZmvFpL/cfacGRfHBp+nnTW195nVKhxqy
j+0sSU7P7zjHoxKuZBnkEl9mH1Qr9OTbZL6UnLN41oZPDMdZWiors5jY3rCF
mZIiNyo8sHhntCY/y91Cu9YFmkRfg8suVLEW8s3idfCLe3l6BgHz7w8gRMuz
YpAwSScQeE/2SMIKHLl0ynmfsK9bwu34xAM8N/6thha8K1LQ85qL+UzrjNby
3m/vBSyZdeoTCFynWjg/qes1dZ2RFwWOIzrHRz9grLvMmHnoag1k6msLcUBq
V82LprjGjIcyjBkQI+EnDMtT9tlZ/15KYphBhoqv1TYSZhcyB8n9YPH8VGNp
S2C86QUW1HfU5ccYWfDO0AZGNJgXBBQMSEI7Kf5/QonwbSFULhjtFI4k4NIL
ZWOfDhBe9rBV01LngfnK9bmqJJ/hmUFRN1gcZExDBNaUa9S43TLa7gmyAgcK
6zswEeqIro2PMcV9QK7e74G3AF/L5KIalvf6fzRav6k8FBo6y/1wKeFiA5+m
CQIwM1gW3vw4I2uzB08uT1BQpzvb3wBfwV59PnFog/P6swwkQT4mw44zWqwu
82zaBuYa4b21qAGiMqd3xC8HCJmhmlt5IRsGK6DFq5Su4yYimh29mShmGk89
1bOradmULSXjKmtOwGz+gnSB9HpYFtx57XFU3d5ioCHNo6mh++cKNTk0e5rd
Vk0rwJrX0106bH2pc2lMz1wJ6uoY8dFT/4rEq2MyrI+chh5hZnMPVZAETUkd
aGnonbWLw7zgXhjM9/M+/CWlqMk65jk0JvNDHdFq+esszBMz5sqT7UmwSnQI
zVh5u6dAcVZ9YH4rpitHs+808kgz5fJZZ9kIGyR++kayG2+Gwe4NfzjBDhx7
rmBkn11ui+ZpjtgOQuREK29OB6RmBYIxTteUFXBHddh617iAcqVduiYhtsGM
JbB0QvyZp09bQoDdJt3SBZMTdW1D8VgEvC1uqvQCYt0gbAEt5nh505vQGtXy
a6ajUuYHmpQDR8cVVRRejHdwFDEx8DaQOR06mlwGM9WpBzNNj85b+tx7c1+H
8JuR12tln9RSri6stqD9eHYRayhkULBx7Fnv/iYeMGDzQxXHkYWdvYNEQ8Oi
SqMK0pY1kzUlS/seB1yJV1MgjxhFXvE6XYKWcbfeBtUvlGrotIFdFOj3I13J
/fKYttTDszlntUVAwSeC/RcKM1o91S7rppyb4FzdaDocLkjqtk3Pj72gIzUR
jfIm/GTloNi8aXy/9X/duB2eIcsJn8yQtHOnTZ7nOEGpzcRYARL3CXq71jjU
BIWaVYlEGrMh+OlQ5OGnNvBazjeveNVl0DTBbcmrjGqPDu6GUAvQm5GrQKkc
vqkZ3kVCSFFoQ57PSPc7FLLwCEFxPievYQttvEAosmdLcC2B4qFiUai/3CLS
6oWanrSNLpqLYIaKzkRmsLSrrTqGPTd0ztAMT9od9j/bbTat9rvV8TlsPPbH
5dar9v1+7eGrB57h3PMKVPDBaPSp6cGuXJBBprFmpooIl21fvzBXQ8d2JpCZ
NiYjGL0QKGpz/0wKXX/M4aWOo81ftV+lYKY+3JUUqiFJ0rVWKEeYrg2vGcEv
MqH6Lk86IZCWqM0LZHhLK1BZBdorn6QZ5ERLNRyBRn9cHbfebbQzTXuaRYT0
ktbR/c0RSBXYT2bRiHxC8hrtUFGAIW08HePS8RAr8fBmcJXxliaTaj3XHTy9
FQudpnpBST2vYqGY2n/j52lVlOymjn6UaILm1hUwAXKjnVHEQbWcnSYJP4Lp
OI6fbS0IUX7czGNkIHXL/WSyO1KKAT9NZ/c7r0DNdaLcdSwsgteffAwrqCmR
vEDukgGlKtLau503zFIHX2BZlPET1DyRb3QBDUnJs6xxcNE0SzqLiA6vEBzJ
cFgpfGoabCzY7r5LdOqUah8H2y7Cr/jmgxCfY/yfX8CRxA0I51puRcRpb8Ut
56bOUwdbmX/djlTiocmPaM0znJxdJ0q0iIQxSkBlUSLpsRJQyGo3nA7H+PpN
aUx4LPa9fqMtArG9ZWJs6bhw3gF9rsy9t1FsyUrmY1r+GMMrjAdjGs3I9Wgf
0uT1+KYo5mg8hZ6KnCP37ka0KhWPvyOO86CL30FnciZ/BuxjKZ+fYvU/OdjP
FT3Aa1fq5bc5Oy0yZv5vstRD9bkVXajuQ4IJiGLVUHU23eTqIAAo8i8ZJ6Hx
jDuyv1EuyN44EXM/BeAczKgpP3r7LiBB6/ticzFNMesfpdtZ5mOEfvY/8/Pj
p88yyC7f50EayhAwL74Qs9QfwolFJIAzRkV8+MKSgKSkRKpRMW+6ZJrdJlj8
h9VAhcsqk5amu8kxcEDmg7BBRGnwkMYulH719XuoWaHnpLDDmj6WXwdrRI5m
z0G06/0zige8vEqqzX6pHs33z1HpiVoOheUm45iHq41fWol0wMNQ8unwUxG8
AP8cE+URdiM5dTz55zwCUWB7mzYiPTrKpvB9KekVBYf+eFsAj+PVm240+7kt
Y7YhSszEQJ0lAfYOseHKDCQNNvtTCsLKqJNRsxmsUoXzh7J0uH2hFEgDiTl1
ut9UPHb2H9i5Y9wWgk+u4cfYABkIs13QXCThfObp9V93lXV3KIK4zYI27/Jj
AhU5AKiC3G4OQFeRRXCJ0VPQQCN0cSSSdBXNRNHhOc7/tfaovGHA7BD87pGL
A7T7kBd9CMIcShl1QQK17N9iCYMlEvXvaoRh/Jjeyq7NeaAEZlGhMrWbnJ8m
5ATkp6gdHgQ2KT3niHH3WWU42mrds1y9uWFh6WQSFm4ia13mvEjVQsuK2kjc
1wTbvmJeEGKZzmTya/7wNSNfyGjXpFg5FheVamc+esYsZ6mk4nQw0b/zzmey
4oZWIGJGod61BD8d3S/oqwYpwfrifWaC72EnLUFyuQPqhRH3uwjkvdB1/Crx
TiWGIxGxBrCcWNVvIBTLj3YAgNqxf1dAt3Xo37uxu6h+tcmmSZP6OToxZUDd
uyPvbpoQoaD64DcjcVYbg5uHfuA0QLrK0/TYjX/NJUEhRqsVBvfm2qaAhJDg
YH2ON19JEqfDVo5Y5Vatv0RMj6vUbvvZ+cBjBIVsFCkp1oYmyTmlfvGGpEuK
PGJi+UVbNKAAECFu1oDIVQYFq05LPSTfN2bNVqhCbm8IUUyHMKuUgdVkMJHp
XY/jQhu4lVPFqrYl8AiyvaFGsAhQh23gqTX3ORR14YKwfHRWS6DZp3RO2lkz
kk4Fay46SeZMOy6x+9XSDowYGug4paZ973oyA44eBQtLJdNYOKGq5DcarV9i
DrhmSdoB4fQopmv9S4cYSHGUDcS/+fc17dGRGV1iGouJlsrSbpBKtq0PUc/M
3pBsUAezvEW0fMcXFg/lNSEbhAH+yfo/13k9lgpkVUkULcKswds6VAPbi16t
9R8sM9se1jOAVStmMadZ1DryyTXH2CSOQBdZRcirbCuNOwsZvpFK1/3xepDD
eaH5+4faZIXt8fMygGGsmFppRirXDcNupfG+2xgYbPaKlkanBKzX704l2WQ9
PfgZLWDcX1XiDGvf5ym2JM75CTxh5MMCp6ymDVCGY1sTajCD0dNGWUeqV4RL
bgBWaJZc+cqBMw4c6XcTMNrmLbsfghUxAuKLGLO31UF1TBp05gJWkAl+Gqin
PIIMB4SoRAEUvdZlVxqbXlgPWl5cM8mU0XmQRZfCcJSem2zICOipUmimFifw
P5foGOQP6pWaWpuzfPTSDWeZUqHCcTYGEnNgir+GKQvJwSLiE97MKQuiFUKZ
IUt847Z1MHM3ZHtrshgpDc627inuYYwFZR6hTYepldeM0nC9mHD+kd2Le6m7
rN2+ZIB9goTFTX+GltgWSZEJN+EUPw6ohYEQcc6NmKeiH14ShMflBVbHjyoL
zOZK0XvkuGqswepUI/iMwvGY/pg3UXwLRAM53bU8VqWff3UyNiw7Ryz0Ynnb
h61NV2UxRgZiUoBZHeZ9Vnb4r4S8AQjvM/EQtUm+QdtJmgykPy0fOSKZ7kb/
iBtPvPxOym/EVqZZcl4DejBY6/f9kg2IgPdecG00aDwxzaXEWj5fxD2NMbOS
hc7wjd0TMxUKpU3N9pxf8eTFe+0e3MroGJKcNpPMUbqmh9C/HF5BhpcZlrHf
ad/kt5tpqwMnmJQhbXc9TGi8DRQ9oOwn13pVQzunuABsYb9vkxy24rw1JfCW
2KjgKPTdjy67GODDL40ZSxYqx89x0jcqUoKp628EmVpxEVBoSZbbZwxcd3VF
VIA1GWS16MQk1xWSknGP6XMs6gCirnPfpUv4yY3HZf+FN/pJT0e0OySFkTaS
Ge570PXL4osDSgMzFGhk4z5Elvj5uLvr4PH4XrKV7UbQwYg+pA3REpq/qFW5
Qr97UIsygkftyB3Mz9NX78aO7QuR9ri4kzfgZpTrkWMCJCjGfzSjnteq5xCL
5mYK1qIUtcGpH1cdgAfxHTWjIumZQQBSbMmnO9jw6XlQDIr4IuCD4GM7423W
mX4xiXSzYlTHPhYINnMWsMYZWImPJsL39xWnnzSvrPiXvoDjhpySJ0ZslwX2
nknL9twzcJByHCzUaNvOi3wkTfa2A2I6Qh3sbKpNNowROnI2F/oxebE1prXx
CWjGY4/BFBV8Z0s1+/UaJD4wwo602iivMOuFnJeBAANpRP//XhD0klXsKBrT
SIbY5sSxo7BfVHcIFKbRNhezNHLIL46Q1AwR86FQDKv91iv1fvGOtaLiMpgi
su6UcwI0CkfB0a4yYyxgpZJQm2pAupgxGX5xfcKKRyfpNDvhRcgBbSs3tQVm
vkudgK0a/rQp4YAwDRYLhZErGaZGfQjbSrXIoRkqhGUVq3fQUArXrO4MhJxS
aSJg6RtbknQp3bXBnhslyoNZGd8zNoV1uSCE33a4T/f/zBGGQHEEFbbm3PX+
8DVbGWoIL4xpexzDkVlwbJRrtjCZRDYCQI9IxOf8boI7tA56LPinWH2vGEyU
6D/j5BDFZ5ISVhGgeOwQBgUCQvaRO5Zv2bZlAOyEcs95R8PQUCGLl2Z1WA2x
2tLwSZb09WXfstQA07DZUFWbKvILtDkzuMZTyCr/h0Nk9tz2h7qtUsfX/ypq
HXsBi3X0oMGkSZbXuHfYRWlkAAFkVm6ENxqojV/9WAwJ7VZ1xTawbjVzUjCG
Goma5rlkTl10ylUCaLfE6kKsMBz0IEdqOWDTcYSLgxCNWqhwEmYwJErMsqSP
q5KvUr4+1gIE4WJvM8nZ5z/9DrfyLPRwga1sf9fjMrzy+9zYCPGsTxmOMCd5
umonLiOxfVbpKTfepQv02IHpMxMHgC95Mn9V08ku+B9a3w8745s9EHAfJUd4
z6TLegvz6klSnzKBXAHgX1qrBAS7u+bRbEa43naTCHVWGiS8IM+pgoM1QsR6
K5xWOBjP34011VDWpUYwQ09XLXTxseoK61Jdf8ZUiDbU5gzBL12EtDjfolFe
DUO7OzgSGI5QDYj0VHuFXIdGsv5cEUY7KXLZUffcWsx1PxOyceqrWMYpJ/jW
L3RPAsw48kbLf/H2aUcMJxaehrhO7G7eEAIgQPNfjY+LOl6JRrbWXRz6XguY
r27HCyhuOJjArexjegZmZ9i8RiHQlUQy1sPnj8/chBZFiAf5hv0uHRcPjPlQ
JMN63iqVAB3ccOtydSaWyuMm7ZxyTxyayxf8+YZR/tbDY7nK7I30vrG1laps
Lu5MOvnNsMJ0xiYCWqxxHkqFFfsq1WATcgRs/gSfbl3cVLFtpxYdkedPT48M
A1ZfmkBjsXmZBVrWvEeHaeGkJPpUOJ3WoaodLGHrKpLVXzsRINdPRVDPlOwB
cWL+myIxBpX1vgaOlHFacaD/cTc1bkMxdAZC/nnlrpc3oNgLk5DUIzbXDuwZ
8RJCKFos4sequg8oDH4oMdjXZVT1DGHT4dU3al7QqHtOqnG3YrBjEER4zYfF
ZsPEbFLsG/jlB8H5b4fDj+1CQ7rr8fTSCKLg04TLP6QFpYl0SfgOYiXj6FXC
6C0W6oNrqo+sCSicXE4u24yC8jb6mOQ4EJ9NBGqZw2gm1+mvea8o2so5sGgG
wPgFXEpzPjVdOPhgGceTaksML+eOeJRUtsonFg57gBMxEFnR5MMT0MktcSLE
KpX+JWU0eJE+c5AF7RrahTZZ6hThJvaS+dlFcJnSg3dzLBmK/PjLg69MimO3
FFog+/2JjFaOSlOdyTCXibEeeWASe3ZOCStU0J8wM1Otr/rCq2tybRUkzNIQ
NPESvwHV0rsKMuVozAk/Bufc+jczFVCLhKfvaL4dWcgQ+KXDwhmlxMWDFqPa
vWCgjykuMaRNq/EHNFUVxS7CCaPXx0vzjsBwKJzvtMGiuSjjAs2dHwxBpDRP
Li6a0O3c6zI7Lz21aeBESPpG2J7XmblBZ8g0F4RGbdjGOYqoolnBUkejSbh9
8Rryl2UbjH8JHPkYB1/dIk7UUhAKMnhFl6KMqw9QbTD01/EtoUlZ8vJy/Ic/
wJNeOgZvYeaN7K5Ps8zWQ0xiL3e6aD965aYVARaxos3PXCRLeD5rq6llmU14
4MbWmoyg2Sbm8uoP+SpQpVuLTikOQgW9CCZfmoEJW8UR5cPN2KLyp5msdWW3
soNX4njPzBaEFC2IVl8aYhRHiMHeTh+LMvTC11qgz1ZIWTAE0WAgC41Le4uo
jZHxi2Wy2Wuq5VYnUn8vdp7Nf9cfj0FWuhOQVpMBylq/qGDxNvCAgNhEKKpD
KrR2wRMkJP0qDnlsi1zX0REgrLDVup3NnIDsCx3OIh/2pZlNzko7XA2m6Ak2
SFTzSotN9BQAo8yGUuke2Wn0Y4stSoULSAIr9uu/ywL1NqAX81VH5rG6IotT
BjUqRBcR2OecNJGn6V0+Ih2xQLWsQkwxOVk0m2rD42STGT92dHpZC5S8G7Us
9wFRUsZY8O8yGOJ8hvhAv503sC0zhZPVZYEF9YjJdV7uWep0FXdHQUphtJ4w
WUSbTGkLRdUI9/30RAkWcJ1ChTdj2pjlzk6h45hyeKrg8rMXVPLKHlgsJRbV
Ht/q8LBRQUANuTI9EFHzqV1r8ElpB6GYv+fK1XoX+3MDXstBj/neg7ffjCWv
6tbdZb1jOijbjPiNiCphHqOg8XJkCt/2WBQCQYbAGt1Lp1yF9VUtpicqmzHt
qXEIwZmQ8KUwTxj+U7kq7Nku9EUSVu8YCKZm7RpGSP6r+l8wB+QKkiNwEvpU
tE8+z3ZFCaK6EjMUzFf85Vacn2N9y7h+dgSF3YixSZnPMllPN9grk4dOmow+
ApODZYPmJWH+W397bBeReSwQkh1Ybq2wVvybJxXNREo+/kGKQtsCPUFO5qvo
7mvNJIopMoHKf6fjz3XReNmRTnYpYqnM+4qaFN6hMG9DkezvRDshpHjwQapd
BsPIyOcww3OB/yE8GaxwcE1IJGf9gGVpIfuC/tpEymGxhcd9wf20+8IK0tWh
YY27NGMdx7BPVbFaiyLNG8LBidoh6oMvTV07/tynO3w7Ym7e2lC/dQLVg5yR
xwMNE3SnJLfH/ZRUb9VTwXiem2VW9/q/YzKbEn+8ZgFOel1pe7TUj91/o3qJ
ekdG5B9cuOX7M26GAx0MSRMGyu+OBoOI662N7WaZFz7R9KSVsvBUEzTplcR9
T+lc0dVodcy44XKWRUQ6K8WBChWwzrsU5b+ENn3oPC2fQN1Yo56jKPRR+tre
Lu2pmxvb1NOfhk4IuvStSgQ/uygvJXkUN2L6rTPFLQwwFDHCud02uIdGdHMz
d1rAG3R4DtxgyZaTM9Nh95Q4r7pheeZdZHoLtJRoL6ehC4B2EdANhse4erUK
inFGz5qwsXGeC3GCWuImSmXfAlMc9fqtUw2PH7NrJhiQ3wSUJNRULb0W+3jz
gytdgYN+jy7yXCpwFPkdzjIEnHx/dwpSg7/lJKrRpgLfqr8RzjgydRxfpIaZ
S/fas+8EPbqAhtpMI4V9m4XXFUmZKFrq+w/oAplV/q7unpHhEw3lK0NWBpVi
zqqeps+3sE9p5af3+3zkRAMw2gWagI3BqAs1FkLCCtFGOyLUyNewoW93S8ik
watmyzH0mV6aKqCkmPKhU+A5eTF+Yu2Jr6x+RJHGS75rqcg8yEVIAKw0xYxK
1nCKzvWQIF+zemJ+Ev/cv6ou1sb7W7T6xJjkvbN3adQMBTpY1yONLRkAtifG
Y85yBf8YC602y7IywU/P45qBAW184o6dcKCJuZZXnRiGEWNEo+XwLFb/XNys
KXQD9g4mzClDiFCKBS2j982nr9Gbt/v4RkFWpIsBSLg7IyButfxIp42vdC58
Y++LS+M0WuzPzO0MO5SXpB8HC1iOeP61AAL+kwxJvj+xGPaYXDjk81c0iTMT
ycSxx769E/6hU8vaedkKYVf8s77wjMs6c0tC/mLB+t1L5DBJwX1e23D4pOXn
nXxNNsA2oX2B2SvXsPynlpwh1wtclhUMTjPMZ7YDTIxS17fG7EQY1KbKqW05
F/srNw==

`pragma protect end_protected
