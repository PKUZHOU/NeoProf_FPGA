`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
aYX4fa0tZtvHprU7Fjvmv4c6c5wnefahOJt7QVYx6FPSPiNPpJAdsKp+AD5V8kcC
sWRtdkW0LWTqLzi0g50KOxoS4tyR6OO8hTzGRQ+DoECiIharOcj9STZ/E+DST2is
fxW95cL+8rT2rSNCPcz8SoEV5SvnGBG6u0CD1pvtrT4=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 11216), data_block
lRo8Ofy0D1iDSIzgBvkdoi/s9M44NkotY/++2N2wiNoFm8hJFzBgC04gxJgS770C
ZJPI9Hj0PoaP7rUPIMxLmdWZ9cwYbqICuSDph99DApWEPgqEAVAP9E/nHubMrQ5b
VtOR/4w15tpOLwnKgnm7vI3i3/zdXO3imXLb7gvHMNeFQyip6JlGlEDMT++yGZ0M
eIr//URCIAO0eoD+LsJLXv/qQY35nXYDbyv+1l2obpkiHFJmC6fvOpMK+ANICtsN
rosCudSZXX6ZCxLEpm3fECiwF5VymWyh6VSeIrBNw7vD0wMKtWRJXbTkX8GG2y20
19CJM/jkk5S9rwx6Kuhy4oUwjpztIW5ZRsHzG+K3s5BxoC27niJ+YvN8JQaHUD/o
RmTiE3EXgpD8NBIn9QiptlxqPJuEiUTMxMCcualyV+Gef5GjNhU7R8wrl/NcISNC
qIuZPr01frmUa0l43yYx7xogvZKRDzh1wZg1GHQ9+yFOORVKNXcOri6ni93Fl2qF
JXpYjdy50Adb9HonsvlONN4qvSQDxJTUhPs5Vny13pFdi2LQHKM3ScfmFKyqgX4p
tzoI8ydcz4gXz2vegOIoyarqVlLMs9okYcTAwqx6LYWz7/n3baTQabPG42qQEfu0
Nbi/YhvF0IyulL86SlsK+PODAVYvw6oipW1ltUCevHRtzI6QapCZQCez7ySY+07+
0tX2jNfIpeiRHok2QsLjnYMycKqRXP0XQGGO4gmFqTUJJ6qwm9sozv06IPDpFUyE
lKYlw/n8nb1LSm/kUg7hvKCV4Tky/nILW/8SjGXZyB5MVYGFrgSy+aG06fDjXLRj
j8QrcgB9fsZzNmJpiBclZwkBYpc2OrCiIZr3kuNrh3IbzIL8FzIhD1SOt20xN/pI
ml+duQudejVewI50ngsO+zyH5zpyWHpuTsKcyXeeYbiofWO7xtrD38tllNe2R8Bx
Hij7Cxgl0E0XXFmr++IoZQPGKFbdDG5/nKNOFe4I2jMWoAK0CrkUix48fONk7FZN
5NwmrKL5IzcLKj2bNAwJZVNJxMPQWeHvqn8IEImP0dn4rAeiuGAxruOO08erZo3J
rQcTOEI3NbYbqwqfiB50bLLd844JU/IvyfK80Ruf8aF9uhqqhtnqi/RKO7r/99SB
jTFIqPR+Kh0RedXcJ85VLihAHIaEl83+Uabm7lGQ8luDuy2MO+LmGO1yS7zfjOeV
wKKn6/TZ6yC4jn6q7nxvE3U8d1a5HQySnrQCLlyVObyHsYEEdwzzi7c9spRkVxG1
h6fNc2aH0tXUvePrZWLhl/J5d/TZLgJ6I/Pebo439M5JhgGU/rKM34AACim9zvW+
bMNMmqhq77WvotNKKJx+kwVaSYfjgL562SAgicEnVTjbhJtwglpdLV0xejSatPNA
F5r4aZyN4cX5+HZNb/geh4pKm1ADW9fU5ChfuVrBkFS++dvKyLI+5SXs9vdmKwiC
VbnJm4hWYVp06BgSUAkSDKz0+UFyItDKzl0gq+14ubUCgvBTQWtk5i+8FfvglYEO
drR+eMMQVahe7njP5yMw0UsZ2DXrKREo8fdY6Nv728C5WZWYowz/OhCjgSm7ppYy
JkO9z8ppPeUrWh4LmeNqS4ZiBCQFjgqiBYagNLpW45afSlLqMTlZyTImGrsXDl33
td1q+cHVMStWkhME3ro22aC3+uEGJtdp4Cty+Dh8cdOHhO27GcCMDjtF6T1vUAf0
pOpqcfAfdvLQv768eeZd4fS6LVYZ1Y6wCRIi9bNXvdODVPKCUM64K9hFUXCiKeTu
fbu/JQIrNytsiftUwBwbj75g8o1r1X5n/z1TPduM85jP+4valcTvz4Eh7gfA5RBY
KS3lA1WTj/fWzgn86FtDYx2gPNnvoY6J9UqkMtuwEghMnnhz+2NvoRGYAuOAVrwI
zFgtiY2oS1z1dx7CW6owAJef8JA3I13zi2iUSMu3NX/bJ+HX9VFg9QbMkQPY3rV9
ryraTMW844IgogIlSe3Zzls6vrt+wBF+xZBmGaBnR58qTWhEPCQ8cHEC2ibrZfV8
N8R6G99bZ0vhMU9k6sWKEMXUtk4UD5IfNs7qo72ErPi3hVmcvHe/LxOxwvWIdByh
VTrTNphNtvzGBVrU8+8Pv+2WgR2i3j4axf3/xVXpQCJr6VGibdYRjaDTFZjnlYIC
/lCkwWxiKhFGjPdGX5D6MjsMfsKSPR/gdohAAsbT5CFmRPCI/qnIRPIVyPweMw/Q
lPs1YibZSOAiTiIJChveIroKedk8eJYJcFEYbXVHrmuxW4UFqZygZEG2aIaXdBxS
9kyfMEiS7jFY3NUBCzR99Pkg84tFOowH4IgvIZAp7DAqrqzaN5ynCZxT7oALbDS0
Sr6DKaX9EeEdrCqjgvBvt1PMKdLyVA6WrzW+ah0lMDmSAYd7XlnAdt/QictmLrtk
KY3t7gamk8mQBOpj2Vwdgvx8YCoc0e6vFMAR9S9mbwGX2OUTPcOjl1K5Bh8/Rf+5
2GbpgKfVcRidAkMAiDjEw09pFjUWqB9OsIB5hUI6KPESZ1ibdeUXIFWRyvt4kVAq
iHMy8fJiO9c57t4p12NCYxfKBjRkm/8rgLIQ5rwdXZXGeCXtpnWciLaXlQu+FTFl
mywcIHWPweN1ocIMrSLOkjbGFqOEiactj1/qdKlORLT9iHg0HwQoHlYJvZydCAnH
cBmW8ky/P4WrllTZbshz3eCfDNE9gbMNLBdcNwNnL9QWqRBGGZ0dXmOGF5wcIVf/
KLI16RdBCZjPfTO84GDnwXWVRPBZ/b3OxX8Kehx525lwV/pFbYk3yHUmbjrNxZlF
uzmcHGM9nmxKmdycSkXj0/OevjTBc1or5n55AFgs0IBEpURqUebc4sKg2TsNqmPW
lqglbph/CpvHYJzWXK/6fFQH8i+MxdPV+pulmqMyXHd9JUfe4rEkA3nNwb+DLeVt
zdSOPAfdd2UEOxDJ4BnR5Ugf5daz2RfZ38g7Lz/WddglG9Z4MtqJOscOX8iGTOaU
1ze+jWGDtKHn0lwB7i7d6ASNjeGftOfRFM+BBnT+5M+r81QkLiSTVl4/wIRf9GPN
7Pd8I/cvtwx6L9NHyJCa9Vd105F1Nfw66jAU/LXjgA88BckOzbNlpEeNKG7+NRaa
BMsX14lSBskPlwIErRGhDLt/7CyMMlxnpGk0BQp0D6rrHFCpbDImmWOUH9Mz0NCa
hRcvCXaAJ1JFpyM+NHqidh4q4EqU+q1MYKWRAQsAsEh19rwPBxYgtVhtuaH8Ynff
pMaP5lToKgmOpVdZ8IGfvapjveKU6ggLgC8w+da7OX/7Ywkf60cZ/32dqBWIeL9j
O6yfb7gLHCWvuAbLgt+PwrVdEIvqEtipXSgV5yzJwsT1tAPEVwuzaAbwDZtxh+Eu
LvogfJnnFhYXBUpm4ybnsVCITIa6WNUBizXTqEPWvmEfNQyOHySUqm1zdLa/Nsaq
VqeKLKfsp1V8x1+TCBKGahTHki3aByp/17SHvBBYNCTLuT70dTZPWAeWomaNwK8v
QNbhcROmkOJbFjuPdqmXGX01Ty0oEJ79RkPm78h8BBUdDdGFtF0NzDt/vYtnjujE
Lb7DTtldZtlelexDHLqLRoEGiCvJJVNjco7yLJS1Lf0/4PwvXjSWHsRwHsDYVlen
THNiB4T8vzyhgBlqRWB51Hbf9hCRJEx4Q/Db8S6yZzMFZxYKItqrZcnJO7u8SnCL
mRvwiMTGv6q4kqfcVVN5o6jOeQrGMffcxspxYh4z1HKeoNKwv/bqSu1ITxMuvOmh
7whaoc/zDGLK2unXLYIXfzrYbB+StnLTjSeNXNcHjEMhrJc82hur7zVft6+RzlTC
PJ4JG2etOot6oZzWMFssVuySZ8wduuiA8dN94OuX0mI9GpYuvOn5goeva9zC71Bf
4pDBSDPVVQJuciauLAlUDRQwRrWDMMbKgnL7wn+Ad4Vqbd7A+nrszIGt0ykCRVZ+
tUw7wZDbF1tlyG4DH4GQ0w06BZKMVrQAl9hYsQzInHLa01S0NiBwqX7lXv3nJZkH
l4/+u88ephkku8bBFbMTPtbmuvE7xFZVGb2/uvbaQzb6Rgbr2I/YYQaccq5dzhwz
XNtLZFvd/StqA/uHbOPf9mgjhlYzGNsCxsh5/k9InpLJd4ZSdgjDBTXFJv56HpL1
VWynsrmyNrtxyFAHo3SQNqo2KRpIrQ1OyqdyOGxk7Wq1L1BHDrXb8dVmvsyDfOUl
Ozt73D187ZAc/kZ5Hb8RI8V5efXikSe8GkQJHuvwNcJKtYWRbr1unbQdC3qCdKp2
rKvqDwHqzGWwrf2su4cJhiE435jhT0QbgQXra9fQLh3WoO+qdgvESYThUC6cOez4
Kd9kP5QriCYz/kOYmwJa5JM46wVCJdO05gru3jnVt2B+IQsE0a8RHwO7WQZkTUd2
nU8tLQwjrxymp/NDV1/6EcnV6347Ht+hpmnw6x22KI7RoQIkHWG7R2Kzr45hKBr+
wJyT1L4WvXhlrECiOImBEGJXtI0zG7iLO3vbgUMi4fnwpZHzU6kMD6EIPhl/rw/I
w9uNNzuy0e4uiLUeBpdnFXXDsplOi05mssynEqPfnzxh7tBDFDdQRwyoc8S5sTqj
apPqUdl5a4dL1ZhB4QeNobhgTgXxJmk5hIheydYNbA1sxqpTNewnv/Le82DrPLZH
8gxjHdYdOvFsAX3v2cUzB/bHxyICBZ5M7s1wZg5lGEFHC35LojdykI8ngWCLkjKO
7fGxqe9vMF8xK6JgJrEU2qNv+FL8xcnc994GkSMLJGrgMnSlIQ4PveMRQO1A/aXq
qnAlLdPN/yeoYPpCRle7vrUVv3L0TsDbHjnAZvztXjmoMaBwomZjBuF0FsRm3CNt
tVcsnweSOfuB0DwXemkiDjlTUYZ/jpczxSNv3w1l/hcXZk1zKM80QURx5I+/4WIF
tBy77vSirr1+NqlO+EJ/e0zE6Fc8FGnf4JfbKscX8b/beCUEqshBPnCxt7Y1pzMj
z4EyVWkJ/49pcwm9h3eqhjyJbc6bQ1fOBYh66jJBui5FQUIf0C172RjV0nZYFHNQ
tgY8Z906Sfr1n+jnp6Vub6PvwEGrLXYAL9ZxYXY8NEcRQd0LlbuHJ9BizlCr6jB1
HlQOBWauJWFIfgHE0ylJJZ0tte6rOD126GFCFgCUx2vSvuSnMS2Q1N259Cs366kB
Z6LHyv1xspCfNOifKM65kJDz8D2bM1/jkMaiRcTe8xA3ScI+o+dY8RT2inT6aDkN
RW+TAXQgwoVCFJE4DhYGaE02zz6LJ/61t1Ew0DM0x973sLtkrth4l1K2h3HZ6617
7QfJadeZrQEWhRsuGK82v7WRUfMjEzwfNFh+3WpoanHXTQJt9ijwxcI2c+wkChyJ
N+rxRmS6wB9mjqiFnQPJ9Tfnt9a7k/GUogNneHALxh7BRzLh3K1hWfZ4Gus18RIq
gSvBzNF9isqMQnD9xkA31VIwFtZGtBrn2X3ZUxKjFFuUli0Au9CRdAUNz3Nz7Z/8
Ta7QSqqFUdYJKRugLo2mAA7bXj/0pLYDSKsDA2ghORhXUl3sNuVxZ05VlMN2a9pE
sn8dFxC4AnkwlQIDNFgxNduApwp/+Puv0WpXoZ9Td1aQVSYl6r0rhIEU69mNAJHd
rJx1YXGAek16CSVrGJ3N4L2y7cJqnfssg0Dp2HuT4hB3RopmprLi1Flw+Ny9mP69
HAidJrnDSO+XKJ/htukJRu59IV+Rvjaa7y57zwcjBZcerXUVqu2sN9I7aMHd4XVV
8SlfPaoKmT45kperqXRlUDJ7fjLLc7MouFvFka3DOnktACi7zCeq413QF0JlDfr4
oQ0LoN4VV63lGkXnIa5GBiM9FbOKp3dwXSrLdHJRI7k77XAEBmFYC399FiG75oKn
9zUTUZ0MF/qqct3ih8VCMIaM6yYD3omvLYUnWkY++Mwmr5HXLgfTzc8vn0kVwDaF
JswgpLedreNhYrgQYDcrDd+jAgA3CjwuWKa8nAwaPW6yrOcoIt7GIBKKhhpA85OR
L3iAmSuCl+krr3ACdq9JLWvfyRkshLFsHUb8IavtD0YNX9VY8hCqHaVLtRBxpzzG
ZrhXd6EKbLYOByYR+gZEtjtCwtzRauWX+E8bzrCYo0a6uWknbEeYBSvuRF/uYOLP
VV4JV/ctVXq73/L5k1uAoUI0fj9OKihksE00/p2UvMB0GADoTmZAINybwvap3czo
flFuIUZjMbox4iZAaRN1TxGVJZ+Z8RCzMSoeasbOoYA9qbt0YLr9nGkAwTbYz8RO
Byr49NCo+FL9r/MJz/eqA2BMSjHxVqWyUugcVhvULKBUQU6UgmJUlByumwYUYwdQ
wFyW70u1COb2C3CLqXAJ/xODIOV5CxsVCLECBAIA3JL7/k5hW0Qf5r/950pzgDZg
zs3wXQf3YBJKs8Z92ngauaj4+ND9zH/fSMfE3dCoqgL9zP4qb5jdgbHeQEz1mm3B
LXTg7NrDVmR0IPzVLaw2asEXeOaAdlg7y97rodzkvq/Sr5gdzXgA/8ldhYIGFSqQ
u4Z1fbl3QsqF8co7bTr2w0A9RsePyP+P6K2jNV3MAunlFiimhuKVZikmXAdUctcd
Hpuwe3sBNp6prNVVTR1zm6EezHyOmdQZPW9u9qoYN3CwsQdkVEogH7aTc1IeLo+w
JkLBvzRy+CtvXI7Xx09fvH6x6655M5jdbLZa/gy1doOsyrTgbtkgFF3G4wK/jFfQ
WhXTqJrpLC9LMEXcthkmuSQCi/fJrCG7aWTTbQGQFPYP7Vujg522FCy6ziXxDf1P
F6M+KA8IwBaDXCm3lpq8MGGmB8ufcVPej0kdbwmO+tjkU2Qj5m+L4assQhHhWknl
VZzCp983Q64OJ7lCA8LCisWaXxqf+gS5dVqsGaglOlsz442GRSUdY7h/veXiGLAX
poK35B7tpbvNJeUq/1VZPYPscYqupxAS0eGS5pAD6b0HvmWl/kwRXXe/Ytxbe1fU
vpoFklVddnKvpd+jyxVIte0nUItiBJvld0OonzlrNfJgg3l5euHLUaO0sMcpkfv0
xf+5EVSyInzCSgB/zR65UYuragqmlWNOc/HQeTwAjwg+a+CHzy5NEtsUi8bTLjOT
qECTseenARQDJs4YzXpbXWvOnBmFjAwCnl3UN2vpnonOOJLBPLonCtjJz7D9Mqh5
7QMRqEidnO8upEWStx7q4oNf46AY27XYiyFYzYT5mrkodox+y/RCHl5jEeeytbtj
zdzRBPDCsOVDMneM0/4B/Fjhr9u6pnxSBaKDLdIQgdJHqrDSjOxQWavSAj22P3m7
Bg5BToJCPMD2xYE7L/crCyxj5tY8X0rluY5iRoXVTv3a4JBNZnZB1xulwwAB01qw
B7dWRS6TqIUxLONgoM+ORx2mc0nybuhZEVjQHi/jTmTYNA6Cw5E2tBcx6lqoFYcQ
J1k5BZSkY7yEHae7srSIEsnYqrf38KSFsWYBWT743/xqMGxM53lWFxVE+rYnPWYp
NGkOsBecRlKV3vvy8k8qJfIcxpwLLa3+5Serupi3vR5UD09GfRK4zfwol1RFqo8U
WmpZgbbM2kD0ZZp68K6XKKNLgNDh1Gnve3rvPvODYJjijr5rzxgOGu2zx3YBbQdF
+/VYrbenWTh63QN6RLErRsN57OLOYKozRAJ9qlfMbsbNqYwrcS9C/7aj4piAWScK
pRbiDmHb9niAdbRqCR17Sr/gjIllSM6ltk51Cv+GHOK5JEDceCErAaWP7H0KaIXd
zmxn1LtZwX6jlz0KPnWPd7zhipqYCOFRvEvDgQXGulqq17g1sZnZXVYJPEaof2GQ
UTkIqIUoZpjclvpOEt7pTzMpv44wRjvRJHaoqoIoQrek0vO4sriXn9IUxiYhbU8d
6Q29xBvkLGsmi0BNqonb0+dy416V+E/FbL1ZPWAT2E9774NEHNytEGNSGoxxm66j
Bx7w2+txV2UH7e/1jNE3QLCfB7ilnzQgLgl2Ofu+UWrlEbS0H2UVHa4ACJKxNaN3
DWmkgfmOsFD7kweHx0O+CE+rLtB+ZYaKeFhjiaIV4psH19Pj5clValqA+1mokQR0
91f7xrtG+F7bC/qdrANWGve7TFLjZGgAXQrw5VPgkwbP5CaKHVIDZzjLbIc2lCfc
REYx4ddtTu0HufPyxP9Lk8MjQAzYOLcWX5m+oKDJbQ9wsifCjpjqpAQ2TafFcMgx
CjsV2CgA2ae9H6I4TFw2aYirfw+W0udbQWtuBqZLm55IT5eOcWiOG058gjjJ4BKf
1vwbjelaa6wGPXJmpjGm4S+bt4+qoFlNqTz7kYvkooYLAO2T/gc6OCxcVvZ/1HkQ
0G4b/dzisnWy4oqzdbkMbc4MQeYovLNzbpCxo3V4iKAP2lZ+VT49wWLwaP/HoNm4
esvUUbrkz+6p3h/oDvfNP9Pp8qdc/qhpKNhAVHlf55REfV4SLWloRWyxnKLOnN4t
wjwi8rYPBjErPlr4sRwHrQfE/vehe+OVx4C2YILRjwGlGQUfaY42pi5pDxTdEhbw
Rt7ehAB3hAVdlP9f+igkEvHOhb5zVcZWcHeFaTuN4LDzBBhMaxVX6rG/CWBBRcsR
jTm0vGvPJUIsmc1716LQkiHzrxWlh/VIIHy6+NCR2rKEZgAlZLEOvZaUmiRCCGZI
caMlH95bCY9qKVgH+rUveAt+r0l8DtKUXSuaI5F4QKPVtYj8ECJXkvJqQn5R0TJ3
1nrxE9IEs7xmsbXGkV3EMSZCE0Q8g7OhQTkdA5U289E5ATK05PcllWKcQbf55xN2
t4HO6L59kS8L0kiLlVNOj3cMm1s5dhHEMYbsgT8iPG0ZUgo+aK2jSw4NCUIru21y
vPLrp+vbr+dYJykVu2tdhygI56Ozg4XHjPW9WSkf6afOgTAJKjjZYHeej9Unp0B2
m7qEoBEtsy5vLNpREzkEFiP4ap+0ExvSjMFp1lSEjceYw0KpW5o/j/mYA7xh3Dz3
rqDxf1s9PPMdj/TF7YgDVVcs3ZTr5kRxkBgh5CB60n10bhDLlGPJutIJUCvMHTHG
xuLF+P3fUH7vEW+HuNym8L4pP/FIDpM5GrW7b/eVs114X9205baNJGMYauY7hQfC
MIbmgea6sGMJVw/Y1d/XCwF5Lmqv1RxW2UpLbWt6faoKOAYil/X6Qt4WmmuFLKRc
NEBoHAobHAU6m4xq1oJKdItRqMtyNMnHYJRx5Es+pK3ZgNhbNVkyEOq8J+EG76Ba
ZrN9l6MZFmtHDyV6x/uQCfge+yDsmu+kUh9FYB0ptsUCEXQwzfeJpwDhIP2tuiDD
qINBAV1NmwJp9vHLzv3K9+vu9V6RS0TAzm3Trt3921yLIVSyaCbNOnD679GFXyUQ
Uj8Oq345u4P+sRTlRCbrdd5hyGdWtVUzBMW7yP9tLalHP1DA2euSFmAsFsRhv5Bc
dUhPlJz58o8lkbSbdhNZQ4fBO0xMdKYtrvrKMl8oXsJxMEu6fZQyx/N3yrQyJWP/
dZKIRNWsOHW32CvHq8i9L8E4wbaAJuTcQWdeDHeK4eKzlLHck/dpgfknNVqo9w4X
bU3XXYUR1DDiMA+gj9Aty8uR0f8re9A1Fd6YTss5QW09tevj9LYWBB/RfCtG4g7/
7r3kqBugpv/jJFG6sM/Ia1IRf5r+d33aFyuttYvodicCw5H5QLJYsETRFkywGzxi
o/aZqnowiy9VNI0NtyYMHG74l/Btw3txHDdwHR6g7z9tAdnySHSgOh3tP/fWdiAd
YKmhzHqSe63DRDEu9lPofbkuWn9BJi4Ie5PTOkuVVXrs8t7O9M6zk3002WEekOeU
9akQywSvw6LZVogZ/qeC3AtXd5XyAEuUfY8YDCmcGlQqIt/Gw3OngTO5RrF9c0Gy
+Pw5xgYpKMgCFL8wNk4Ngk7f62QgY87r3xJteRUJXk9sTgNlb4x6IA2RaNYQ1T49
Zdwbl8NBei2e3+JYFZ7x/8dhNxinhWsJU1L5EsXlfczrKuGlVJ4FKOV3DREEKe1X
LBj4j0SkF40pX+tVPNsl50VsWlzG0b001slX98T4ymewEs/y3ey5POmNsE9U2jwZ
wBmuEWJ926vzeVKw66YtmnVlfzF1wfArKO2vJ5tyjACvgWOxvt4bRzO/pG+5iqMu
ADZidjppnMxxPO7xZMU5RQwvh7eN3zqhf5n8sh4f/lbiGtdjFOt01826ixYrTik7
ut0MG5FuW3sFDqbyIozpz5UZOrkIlHtc7StiUH4X28VJzXNWMmsWWBHNFFuBdUvd
a9XkZ7NMvmj4qgi1A88KxjWTJvTgGwsL7DrnuBFUu8MzJSUu1jw3O0GyeXHByUx0
ysapM3fxYqkvtatExCHWUFgkC2AkB4ipNwQpPlv6v173I9ylVH9fBcVUuT4XKDpK
UgK88G00mkL9UCqWeAxaLWVUpMkq2r/H4B5PSNHeJD23eAV/i380jwI86fN9vP0c
i8edEUqSaFjnIeh21bkDjjQWWBJc0RHmuHiTUa8nt6id6/UJqwUm8qePawe6vgiT
agZwxBev7w/uQthQLJPyJb4BcacTnRU/6+WY/g6Y/fkoibjBhVLI0E/kDerkh6UU
0JF5J4RNTOVPYAW3S/43R/lfpX6FJRDSqQnxNTXbpIiMoOY7myYhOijZeADSm5Ku
vvLhnkmoyzRq3dzG2MiK2f+mu16+7bBbWUVR/w7YKR48GV3UQayubsm8lI2vavX3
x2PbLwYv58iQcCqGuXgAkWbxPb39HwShiIrumBaphWsKpgaUhITpxIKaQ5ud/5Yt
UzlQmOXtSCfQ5ye83U0ZuzQFFLG0SVL/RwHNRer1soTRCmf8SiEyTVG+8PQDvbFD
jsZZGxFsQyYpIzyTQvkzSY4HBQkxVOgEZ8reBI94Eo6admMa1IAPlAVALIRXiMe+
bEkxkUTswZJx11d8QJ3rX3GR6cym4d2Yi7wri5OK3k3A3s9IzGjIqCThxOlKOB0G
dxZNkDMUCDC0RXVafHdQBrErsabFLfuEQfv+TRuvrLs45X0hs89Sl7inZaRne6BA
wZ5grUe8hXG9HIPMk+t94m3NYTw7rrkTJHxpi12SvC9KdugMogCgR67jae753SYi
vOeaOuxpSlWhgZXlw0O45HLibQLtB24eOxOHBqb2ICE9uXi9UJIa/IP225E9Y8O7
hQOHWAmfhTMw6F37y+iTioAVc45eXGj6Ci8EuE4UFATfPJ3rwcWz4yclGndlAF3x
PsgObYnTEO4OgU21BSpZSYP5S26YWuet4Ik9V/sOFBUgr6YgTLDHD3M3h8kkTbSf
FdEfBf4RnpKtIKSHHt5L7umKYQYuNJ/i9RSHFDQUbUq6VrXN5VLpEwPcYovQOzyZ
YrsyFIun6cOKUE6BAhv28hWu2283U8lDoBi1LzjDAD/55i4cuK6k5sxBBXMRE/s0
kOLPzwY9WCMBDd+GYfO1oPkz7ORLD7x8hrhOBM0M1kKGeklheIBslnbQZoK2SBR6
dBdYZpNTSqUW9iLdVW8TX1XLzgTX1ssW+GHhFv9mhtAu2MGbMBYpBiCalohQ4Niw
ip2fDbn+8uuylz+IEzpFHmq/bSITO9cHcxh+A+6tV4eghimJt1y/L9wsmUgXqo0o
vQWbwoLrlJriFKH34BZ59nRZVCiU1LrfjdLr3HmFbEa9jnysA4mAVBfi+l93Pgl7
cz5FZ1N2VUbU3P7Pd0o6tYNUr+R8fVEqRPq+eMtfvYwAmmlPDoV5ujm/se3lRb7E
hp2KDcXx1q4xsCHKNMXIh6e7rhCgFmMY9AyqA9g9aVWF4lpxZBYN02gDNMk1BEzl
MAkqeKlDuu5fRMMycHmqj04ez0wMD24VEZuEcpkPQaB+9U8ZsoELjWTZsXyslSqb
qYyBs+N+04pZv4/E/M+qkEOaCaJy4Acu3gwueQlYSU8rvM8/N+GDTQY+tCJNzbqO
ZeGshKOg0QevC4OgabnP5bcHFSc4RLuwZdjpj2CgzbgPu7V/8AI+skPvWJT9IWma
q9Limv0gb89e5fIgHtw2x5r88CfnPluY3U3d+L9F331z/KztykZQuuIfLzQAEZ3Z
K0dYzLXrZPRgnyHD3UlhrfqkrJQkzjDBhwOL1YqpoNBRFJ0enqaAaiLUUEqtzII7
I7zukFQe9FGYDeZB/zOOfNklRL/uoQ8CSRlgItLqogaCb03WhTudtS5eSg3QXWoM
S9s0CU/+SgZDqYOUg+nxQpxXGhotrs6/WI1Bi+bC72Qt3nTub+KPcshuBKErgXxp
tgPrHxi4s/2+Bq5uCd2lJqKZzuPpLxlxko8uk9xABPyDKZqInBqmudEraRxhwQpI
d1FY52Z57asguJfaR5GKPIwAA0ndmPXPVCjV23ySS5jltEhflEKk8LpOWLGuZ+bQ
gJxRZDCjI9ytx2OzYn/RNuBLg+80ZIs3wpzOI7jbfOQppZNPDZ3ZZlT1KfAd24Sg
5xcvT59zZKctf0dgUg8RZ4QJBrhHxbwhCyGIJCo5Y9SvsSersVfGZ2vGJqyCx80H
CY2u2Jz8fZN2oYmzsb5dGTF4ijtxvR3XURzbBKGKca4Zq4zHUUidy3YuuC4rNvWE
x/r6M8YUkbYc4QF4TpA60v6pUWBOU2Eqq2bmsBfrqyFAw/Toitu8h927B0Hu2BP5
JlZB+vJQizeN86PIsndesKcVR5Q2DKH53424SL+TbwO5Z43Io307cciuZojrT3GG
sGFJzS7jj/9NKF4rEZIdtUzYFX2Ljh6lp9tLjsUnzdR4IyTe86t3bHrFMPeyg6MU
r5hkgG4/9Dkg+aSD6BeXx+4NuIWHviqznosK+dqWJhhztLpw4TsiLO1Qi0/nGnCF
UtnOx/C0lkj6o9wr9cCRvsBrwlgdzcyPhZ5VKfC/a7K/7ga94rhi38l0Zli8pwiU
LKUj/oYxX+z9bPrKM5hPM44xiXeedLJH7PG17iygTuStP8u6/ia/jrI82TqUyPlm
TIvfwmFl2PZL27dlsMIPbMRvpJ0J1rfqB+sQcB2OIGiqFAmRyCt/7YzFzSMrsMKI
z8kCUmPJMYI1ZpW8lcy4pjcDaErja8Xjv2oE/loLZ560J3XAHzWovf/PDVo08kDm
lJD3amPs6p2rJNyFWu2U1lOoxtCVwq7p20j5kn5WJ3Z2Bkqmacr4Qh9DnXjmXKJI
hJ79WhqY2QAALHglyGLVpuss0g+Ce2f6GZHO+Fo6ocJ5yo/1eKwqrdv3JyHv8Sxk
THMygiUnOM+4XCIxWVhacHyNFhkp+MypaXHzYmjMf0i9bUp63Y6i7D1KQBzgPRPz
LAvkgHTNDKULNYzmwAsbEiPb8kVHxW0NP05cPMQvl8wFBOU0eq2fWVHdwYoXh+nM
RfQ2GCUGPC1w2K6SItvCDqNu5o1+Ge/J4cH4qGcqPuqpmGbpeeNBosO6p8H8z4Gj
lIjHHT5A8BX/rHf6Uw3hk4W3iC9WB0J/ivgSUmNzJjfL4W+zufNoDa50VaNM3QTt
uztKFzJu4yRv0dfyfKcf3p+1TX3WiCLUdiFDjQNykxKYy9JpxoyuOAxtD9SJNQ19
/AUMUR2Doy9X2+1spBkLWek7oi2WH0BRn+TNUxajSDQDYLdL4gJyFyWQ0a8bD6lq
UZHvqNIzj4g+tk28DjeUGNNTha13+I+UxRlHquYKgZ8uCSnsEc+9an2IKoT+m0+0
qrNRASLerTnULOa1R+psSgr41PZyo9ARNyDFoSQmNSUdMAQXzYyD4ZSZDFazNvJ/
DqnIGr/tdmHtz0KP4Jsno/OxwMZWSdBTJEgEZO2K+pEwnClA11zt/wGi2086DzZQ
KxVrlDn0XLKPWVyNAlRiEmYAR6fImOPAXnwIpTEf/5NJiE7i+N5l3uCyPMjRqCSz
zO+Xwv6b+VosIS1ClV2Plasqoie2w3uEOySgtYeS+epUNBEzifKZOdSLXcxv6grt
AX/q2B5lNYkvlYx2VcANFhyG4jSaQhzzAJCGOwwzecgXhyDYwZdvb6jWFwq/fy9M
PfdIJfU74vVGVW1Wjrpn91UwFecsD0PMzHgMPUZRXmD31xnSwxA8IIpkYfBNhwP9
1VG++WJzDP3IAWYNmXzuJtGAlTCm0/v+vKtz2g7DNAb9LGgJXIUtiAdb7IvwS3EO
Na3fPII/icCirkdZAZM4w33XTWM2khQ63JlXUtXeXfOcb+fs9x/yi0aKXz+KzfRM
AoX6vIKlFVzqevhyCp84hBN7lfRKSWx626kx2DhtqFVugjkcD5YnghE0ra/tiKXe
4CFVbCPlg1LYNcUMumrLAaX2YhD9+QBLF4noVLheupbzGRhI2GD0fIWs9nRpgDs0
/jrubnmodE/9hsIXvPfFcJ6fzbwWI0FAyz+5mghSMfPtd+C5/4XNkqNV8jATh+u5
cbEhaix1bIXytPzqSJVbTRmnhAnK0IPpgLxiYhKhIK/S9KqUTv+GkGCqkoCta/Us
OITJFlMnXejDzf39MvVS2lcTnjPSZvPaqbeTh1iXDwlr3KdktaZOJmwiIC0t26Fm
Zyj4YnDmL1msaZc/ehVj1FdByIXWwCyeOqfmn29kJ0tXJu/1Gyllz3M34eqLCjsc
fjyjQNWO9zICcmx6W6+c60AkYsigjgz8jFECTs+XqebZOh/QBGXg1HHi+udzhH/x
pdbK6Hw52O0DT3OX/TnzkdF++JnZK73rseUyquJexy32YhsxOC5NGzcIFgJJJpbi
S/XpK7VH2k4Mtl7m1/hZDQLmF/cerqPHDrcn5VwUvEwC/70ZvqGcEveLCuYZHvOP
s72wHR2Y4J5UntwgT8TiXlPLPutw048/C4iUTNKgqaICuDYpTrQ3U6uzhbwGphDv
srZFu1YKf64DUVYco8twGm7xKbIJ4PFsobQyJAbblKJS2QfHaAW5TCisO9tejJDk
jSE9qDFU4C7IvdhFdfHoPMmiNE2cK/JvgRu1jAY2yn+my8KYdlBVqnpVBNtG578P
OAmeYW8Rtw8zjRHiLvxDJdlTmPHn9A0Z1GdbWSMcyYQ=
`pragma protect end_protected
