`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
i9nfEBx0vilYzWnuTxUrUQ56xL3Nkh7M3eW75150fKEO9ERnJyGYoSNZZsoDMqXn
I/EcLMkBhAouQsTRHka39xxzRi6zGUEZmpThhd1SrCBFfJy/bZryLmsgm0kIs90K
fGtf+U5e8uVz819LACkakCYpSndmZwc63IMbxPWCwwE=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 44944), data_block
7txxRhyIWF5CoQgNZTD7Q6nYJ5xYYQXK8nkeHS8exUpwG6GixE5Kd1yAY7YUetGJ
AnGFu9OFAEUg4r5ZeEHiDvLeoAGLJoGY2xgadBwfU/5Kwv7bMPttVwAP9tR/3yzj
XZ7Z4q5N7qWYzCeBa5e05sCYtURZ/8PDXRNNBDoTDU/fKjvpCryf1K5tzydE8/i/
ARG+2utqvN5eQgGn/psqGkNGaBobWR+w0eBjw3j7QVysdruK/SNpz6cW34FiB0DE
U8GjqJ7RvrHdwJXBjGxxv5GdXOzQ0fPNqovwLhbvAdiC89pA4zlcE3Un5u1s3GQL
eIdPmFxtonDZLFsAxfzEfeuRdiCKZYyiJU3IjMCVE0xIwaFfaw5nQuhR0dVk/oqN
/N1W/kBzhr+NAHQIqayVIVPtFsSZzRodZbYPwEBepprzJMSYwnrj80KT2KRvlTKb
mOFfn/emKkk1qU5MyvFoxSUzfMrQr/8yYH3khwqOUzbLPWL8xFymbc0+pG3Y5sd2
+Jial/p8xTwYjDiQKDiotuH1iW8FnZspbGO4ItvTucQUeZCoKb47z+vjFvHs9h0O
BGeQvd9rHb/PjtPBw7NMH1NXUCT5YkqNpqJz846cXU8yimIXKGrOUIDH+fTp8gXO
xTpNHxGYh6fEXPk4nwtr7aDqESliq8l/Wt2T972HdKldB2w3x4jQwbWSTYwqN4wB
Xww46Vzc5AtUUa8aT+cmytr+EAIOomERJdAmG+3mcz8+yHchOl4oDJf09Rxsid0i
6BT3lZItUxmZAfSDv/0GsS6WSRud+Sb9P2vpXDXkCXEXXecj9Tpm5V7PUxryStYB
ds5yBWhTw2B7PMg8/AVTYwOGUzLCvysDGQ1fmJvdAEt7OJje0IxvaTQaqZEuZaum
I2tD4UjFxEKf9SiWg8Y3SaKDVqJB3TjPAiE+N8PguUiHVL9XbVfUHvxAZxl/OiL7
XwvuPe5gh3B0PAS6+VK6SKvNtATwlm7j6VQRxjvi32Pifx/JgIw6fRwsfu9OrPCN
ArFNrfcZHr6P7WLblAVxGPiZ+JVg/3sHZXE7CTtkVVPyc8pKrA16AWgUySz90si5
YknDFrlb4xEX2XXJ5sm4l6YY9v0WaPL8Oweb2F+pmg2dMoNO+w/66VxQ4IrRfhF9
kD5dvN9ERb44oXCMl4+5dEGrhnFcrRf6IhDO+zUw24K1gQyd2XWz3MTDtDrX5Kxu
xeNS54ymV4snHqNvzcONfsFpts/JELJBixzhTTGGuHVkx1YWTrHfHVbk17ZkeFe6
0m27PCu415vjawoSRbYSHept9uSYWnUiR2h0VdzLU6HJmHs7t+eqdVYt0zwBePW7
KiZKoiSSdYhpe7DTzPre8MatvAxtBqG7liQHyg4WyOOJF28qjaj8VgrEF6iyE8sr
5kpKgbLo5xM9qS6p+UO3BGODWyJVD3gdzCL3ORDvQNanKn86+XsG2FWB2f97+bBi
k2NzK3PiS/oq/j9Gd6yKq41Q72vyMyTc0MMiU5A7OWMFCzZ/aXRSmA0mPYa9FNtn
tXLHhKRmLTd7wBch+umlT0CfJHx7ujzRSeSA1KGavFpY8Vdn5AlqvCcW7QJSemZm
C8pNpZ5gMVgtBG8QqnF68igEBsZlXS1VaXWqcJGrbKIAtE0+a/d6umHX0GM3/Nwj
pE1jGCzz0PKqUtYAv2xO0kIwvfZoSUUSkpjWYEAUk1KK89eGIaCU0tDrE7wAgcnR
D2xP8Ers0qdsjC1wLgOIjcgf3EVxYlrHL02hUdH6r2igacoiIYmD540heNBIkts6
3pcEX2UeS6qBGhT/CpWOPwoatnS7FzP9mfstkfZ6fcUJdscPEoDS0cxhdQomuM/y
v2hEbz6PuJyzmnCVSFvN7JBz2kRn29hP97EAFEFDf7aTrHSrmmpXMzQEHaU03HYE
3CsJkwU1whjDgjH1MLG1mMopqGPP4MK5ClPjfoleHS8713dfWAE5FjIKO8Gves4u
LCTX9KNvFjMnM0tWSTTGXsnaOezEjWjFnCAdJKOpptf+RuTMbaPN93YQhR6dq7bO
vcHCwCA7Cr3stUfWyfH2nSEAQ77Azwmy8T66UkulGCWo3ijbsUNeQdbXFyh6RmSM
0D/2tFEiPMm160hG9udS8lGEj0J1yw3HwbcWpTxd8FqEwX4f7HQTGjjp4BQvXxiV
ZY49fOtsiXetsNwoamFWuiqm7ngKoXsw5R2e9JLvViy3NDL9azV5Ds8W4ggLKz7U
wj3O/1C3sUvJETVoKYC8GnbPOWNFTi7ykjvAiAiz453rRyxcukKnDEwoboBTqxVo
E/KEVTOMjon1O3sfCfSm9Hfijh6SUiYFT0r9i1VfNAW/WXWHv6paW4NMVX5T9QSS
kd6fexalGOkPgzeaWEPkW4TVxzlxDK1hRHwXrnksXJsAX95T+CmHyupxwW5zCoUQ
hzKuGaAm9uW2UTVVgUIUDzAvd5AQsjMKpVjvfGeh16IfH1P+jq67UQydkSp3Fjgb
IgQoi1gfdtjPHWXM6WVjbFnU74XNwIlwmaxeT/uYASxmQqe6FCTaEVWRJm0j3ZXV
6q5o7KSejv9tFwr6+mCSPQ66xQIRndfZkizns4PAn+Xu3YMXSlukyvsgWMM+uabc
yn3sMRaOYpDcgGvsVuOKur4BsVmPcou6xgp07u76p1Q2rwod0cRS+qlNX9GUfRkd
NaaSBZpg5I5DUPpJdRtagsv7H0R+SyQRYcNjwQ28OV3s/9ZbtUh95mkBdbHZhyeZ
xxiRpgz/B7eQS2REL3NH2Zah7ivmNeP1uDjjDN28O4OeQxp4mtai4WveidX5HmNv
b7fEbHsJ2fVPr0xv+O7HE7lCwf5NE8p+Wlip3NhpOUThheJjB08dCst0ACT45jbk
+FWBwjCxjEB6FAwkF5zL+/RKIMOsvqnZlD7FNefGoWQjQs3GAuZfPcoloy8POhsX
87+8Fhjcm/PgsNREO/IZ2jBKqnUQYf091A2Jgy/9ZSl3lPwCrbHProDDTCKyHqcS
jtEV4PcVYz4jMVGEjWTxIqyGHDgT2/fwlRcRbh6bX9JVPTYxXzTmh8n2C5Wz/Y9c
h3XfwzeLqj94s4/kIOjPV7UrF+L28ZS3IGD5eLwHLwmEoPPrFx2BjZ8utgPM1/jj
w6ohj2MscI7nvIzRs3OFQhwNXJbxCQRcFnq9Tz2sn8fCELaDpwOJfh+EicHhUEQT
0FkgeyztOfr+ehN/T4IjD7sUvmeBauj+Z7XWfK+c/DySlCiuEe+oqADoh9KmI3iR
KCz/38h6kxydplYPOmN6lFmCJN2nzLX+L8ZE/f4sScEhUtMvX2qZtsfmhTiTNb15
n72mknpyuR2Nnet7hezIOPuRxmvc3ecEi6+6uIn5797zonMHhUajkXCp5m1B3Yun
L2wn6deLYTq+k23ebd2d7frGstC9cyY0hFBxSljLkZ68/Fubw0P/ILuuHNjYXtQW
/vGJYbA7xb6T2IHFaZsNfhxCsbBan/4j4XC6KNtgpCyQ4L4XP7tOkPi9iok78Lky
xkwgScmk9WGraUpvQnIYkpU1PCS6tpVpEPlyDl3M4hAk4HZssaYPanRlw4qKGFC0
i2voj1GE49ikkfzGNmEV42qVRDLXby5aJ7mydOwXmJkkWPnQLD8pVuGM4ZMb0NJ5
i4ELeymWvMHUyzHWl0CAqhGYduL52VQqXYikJNGyF+A6bXwvmRdLBp3ifby5l/8J
N5AhCkUOGCQXn5jWXeSwE90Zp6ltzn1mYVTCMALLtW6RZ1kQbVFbZRkmOmu1GD5w
O3D20DFRE0z7hJZV35ET0UckMIW2EvcAe9qcTN232DnJwPoCHmimAZvThwl1tSOJ
OoJhOUSOgZLSJCBrWpw1Nyi7GRavxCxOYocxsl5RLDe7H1zNbeR2wFQdRlDsuLo6
+sIWUYgfvfbxaCOnss1/Dbe74619r+3X5b8rv88aUaHI1vC8J0eF2s9cWb9yx7AI
6OqU9/hWWspw6ovcJAX31wj9yAKRNYvBbqBcxV6FO3owWotIN7kX42BzC1NJsx1G
uldPLMHZWKhC0BVZlJ1jaZv8b+pgnrlY9Z4/SkA6WOHkkdf7qKhHmYQC6QnkKgOx
KY9YXhq4d+QGHCEzwbYxprTIs0VG5D+5FdOfU3Ks3PckbumUo6D4rHm9DlZ3FXBw
L48eEM8CEGfiGiE/hKpOoB2STb94ktkbX2HQGFGaqqSVTSAreX+9BuEq0FGnPfmE
Qg83XmwbXpcidQycZt3CY5N288EuTJaHX6bOqFSarFJ5a5UpQJA9efg9dsYKNAOV
Bn2HkiL7WsMkljVB8vEbfdavmgbmfqZytr7wGXizP0XOlGRMOLyB2obdZtV07/7A
bfVSbP7JeUr2v3mNVdXd7VKlQsyNOQijTzm6rJ3Ruuij5spjTgV0+YEh1vpmuLo+
Yav0lb4UL5FzYx+NJHO5NwEwznnhAjphLx3oVpDGgmdDNLO9OjMCLciczbidL88a
NiHHiFGsRJn2YOvLTZQDkLBEsnaloqC8bL7PcLlUlyaBGP+FcnmSYpNtBK+RY7l+
IwZ8BBAWhd7Mmt9xj4Q1SypcNdgotuIScAUQpmTzFxb7pZuxOCvJnyuzHaDZOXTE
9mO9TC7UIfAy6qZRFsjWe0idS/mPRPcORL6J0EwPK8h9aAL2ixPrWd9YraJkg9r0
l4rrM3D0ZWPQ1a9MhbQdeetwl1BhD/dTOGzVV7igq/ufIoVqv1j9hDbFShLSrwhe
n1suG4dNRj69PQuzA1LvTxAdii3jXyBjTBUe9iadOi0ovvkuzt6IX8qGg+R0M7mz
drGUI3UVFUv0rqFJC4O8mBzpYYmyleP+Q1WyOC+bpUpZKpcjl+3rtcDrUPmSz0sy
klj4UC2dv8/tl72z5o8i1iny6XYEMcWMwvwjP1d0TkeJMp658NqrY6EOn4f3Rdzk
3TxP6962xpabYriwuQkf9oShGG0ntEQFhFOXWVOjSGitcv4ZCPNtp6aO5t8LWyiU
0f/2kktUvZLtHtUXzEAiLc50k45uuLZjEuSwAtyIC4qF+iJRItVWBgq7CWs93MvA
JNk/S59p415m6gVEdh5b2TnpWJ17aaFNSFbj45mImyRIzF47jMO/pTBetP+tI5n/
WSPyLlewmZdrFOy3Nwk4Rfy38FDf6Czak2PJimmHVsFHQRYLtFezo2VJ2/4n9DQp
zWkhP/9O7X2btu7FVwfbqRO2eJo5gglo64bFu2ZkSc8adU2HgSPfJZjqzS/6CqOc
T3PQSYUyjHHX9XDhvF/+Z0hFfsrk+mT6/Wrj4Q5lXKhv2orjBrjL92AXFEyJHTlZ
Z6saDr0QdCSiuKjhjKaJ0nBHvGmpGCNisq6wf4X95TWnRzSU7RFxGMu6f6JmyRM1
0eBA916x/YwwW7uyIpHc0KCm4m3+kMtqUYe3O53rjh5QtBt4IScQM8nKJWNS02Nz
egaxIWsZ84005jd2ACpQHpFNLR+cikL4E6jRns9uvEdarcSz8pUOfi8+QGa/9me2
QJAthEmUypCJmU0z0KPPXlJkb2EDc0F8HKLlB7g2mxCvBMpaNqxO6g14mElAdjNJ
MFopKUHHF/jsqFmVINPuX6u4aHoixn+SEE9zQVxNmRiKLlEBxK2h0ut1fQo/xqk0
sIUvNRWx1tfrF0pj5Sw8G5FLdC+PNAZ2gW/TzuLm+u9GY3D5VTT+iuAsvX2IbZRW
bptWB6sPiapVcZTYV6/As4qbPOxupZWBTWdu8GjO32dJq6Ys/SIPbwByzmP5t1E2
rZIchk8d1lYCkiEVUuyce4gqMmLgZnEeJqic5EL7N7bvkXmBTyh2UiWyGDHv5gw6
KyJsFnwh5BWkjaI87vCqkXmWI5TVw6vGY+/Xc9BPFmXuL6d33EqsRvXMrciV+lff
ITJMWbCCBuOoV1bCPsKo6NqDx4YYTSoAnFk8K4jk4BzvFmPDYc2501G+AYj4Lo6J
nLZYNYMu54FKghW7KB7RbgGTTDBCN/puYSOYByvk188zyaBO3WWGkwQJebxX4kDX
fAXlYDHlZcxN7UUzDIh5+Sr/ucBUz7XVlI0ZqsLf1J82zdwMn/XIR7YriuttXDNH
wz8Zgz6nkUIt5XdEL0ezAhYdEG/AfOLgJd6cSnf/79SzHGwis4mJb+JPS2RLDJPG
ocyKdeR0Cvn3VQSn3AhaZlfZSQicDeJRetviq5x4PixK1yDl0c/axVXrHquRAETN
BCgY/Wf3yfks5IX9/ZY3nPn8HUQW6QrmtCjZk+E5AN7htG8AK1dSkC77vAHw5I5M
dhYAIErTeo0W/M+jRervmXuRyHFAhptZ8ZSAG23dF3FapynpUwH9JOGK4ZE37Tcw
rT8QmFD+DEK0IhDt1/o/jnHF8oPgQqmQi2k87GqLkwJbSCwgVmpnKorZtapnJ/Mn
j3oVwT5dGL1pUUkuq9ZIX3ZGfSfd5V7+XTyMkerdYUk/WxmyvCOUdmawrZjhMPZ2
RujRJNk4ugu96XKyNgSOpU2+luqo1P5w/3ro2iufRZzsRXXfCARa1vJ9phpjtDyo
5E9vYEvMWUQADVzbp6GlJ69qTVB/pf0ef3EzOHmljONPL4Qgv753WV5cDOs9WZiG
42LhDBd1cy+5nA2OjB5aLYfrsCwzvWNdI8voECwVjKCve3w8u2GxEKbdxqvt2v6n
hXY2uv0AQUcLDAPcCYWNXqw43S/WIMs95brZuKbUqvsV1g8EJFI/yo9y8VwMc8ky
AEEhNBkNrp1b66/wDZkLQnqYp16ivsi9fNXAww82driAkQ0iPpGlNHGwOPNz886I
k2iaU8KsCyCMJLkyjv3DHDJepmBY7Sek9Qsb32UOzYf/VEuXCyMk7ak4cAfvuf46
cBBDsTjTrzTr/DLy7vgx1XFTQgo2DS/SKQFXYvZ/+OCjF/s+VMNRljyXMGyPy3qG
RiZaZQW57x7itbmnvxeZdwrqnI0zecuSkEI64TRnYsLBmgUETXUJgljGf5zmPVyL
fa3hlVVEF5VpFHothBrlRoVpZedpfafBn8h4pjqAAuagQ7/6YB1IysDpK2DJupfC
n4ui8eIupnNoHgs325gPV5Pq0wS1/hl13uK3QjqqlDeWERHhDmjhruV7sl1j3J1N
p57SjaV0c/Q9/lWLsPvkDVOsabR70u/p9dEaoYB74VDaR1AqB/cxzQjKUrjmo72i
ueQqDz8htUw4mKWwkwagPisa2tkQJntSsM02Q89cg10SANVFyUZA6OTh6KR9ExXv
HbmyMmR+/RV/5wnM3UJTWAAhpvBrIIuWvU7JKR/pw+6Sow4x+lA9gUX3N3jCNFWp
EygqK2rP7sSSBWCIPgH1Rvwz/UXWIIFje3js8xxtqjLGSEEqXf++NwO9haKVUBst
tgoTsGuwAJwdzQlIScqlKKpD/CgQz1KB2XzNJazaWPOnUsVsIKCYNVPTFvisWrqJ
v13+H9BzGVR58x6vqJDhhhMJfHMgWvNpejih/HLgygtVd3PAB5fex+5OH+mx8Ljm
uTBY0J0hj4FMcXvEs25AVaeM5+zJ8xZAPogpedb81L4hmogQJoSffnSc3lKiFmh7
Agk2B/qLE/2gVoP1kx1b4y9V+QpSmo960Kv0z17+zQOzpZbAAAJgn+LDlQfoWsRp
DFo65qRek75VFYHEmraCvxnqGZhGQBTYOgNsFQH1FSn+FnMRgOBEvxBxtKslpmDQ
114EKMSzqsumNLFTQ2ART/Sz5/Q7KhzzMKwJDQclIJ7uOiyv7h6LYrEtDdEEWBIs
oz60bs7d0OHcxY3STtIdg5EQ/wmIPnNf0RhKSL/mJD4vpW5TkK/Am1R0FkvI9lJ6
PkdzD6gmTjCIBRAgOzZhYZgvW7Slw6xNFiiAOPIDQPZu0tB9vmqMW3MexRIeC5l5
tcryzAi3yaLASidx4a3ZEP8N4/Fxiq5GbzKG0L5MYQhU1frRztJVPxoZdOqbJOSP
3GExIAMAqIK1y41BzPKPBNwKJoXkCKNOSxIZQBVFuH2WuN8KazftYeh8lD8Iz5lq
j+h8xtkOeyu0x6ySAbkUBTD/OAT8Lz6AdsFpJLNy75zt70VbGiSOCe/Dq5vd0zI8
2976r2lxI4PsqK38OsG5fauNpVaKYOcOHpfxn+rN7rKLoPiXhdP1Vsl2VmL/AJXE
g8k8wUk/iTogBwVVMnhSJxOKgENEsE1mT3hC965g+kS5VelzkDPFW3ZQkvFtZtb+
W+HLbqNdi5cMBg+cTXrh87XlltEhr2AaWjaUaCeWt+jICWpp5J5ylnMVnFqP+Mdw
XRwwcCXBCsh5PdJl0jdTeYW5dLvl+NyBk+hyPMqWWaDrsWHx/4PUm92i8/IO7wot
hY1EU1JtiTziUGf4tgCUMXmTfIYVCnrcrdO071DQ8WRKQOe1cVUz96oWptoZ/Hfr
v3ZOwgwn8qLfSHe9yYAuCROeMUnYmuyuny6wBghf55Yvms7ywedixVKkokL4ae4I
Aj8ev+P8/GsWcOAUbhdpAFhtI1W5tuVSMLLuEJ5lqG8V92EY0XbcMiWAXsxqnnzt
pskLvLOcHCFZEesQzStB7f9KVU3vh3XaRllyDRff6+PG+1NFvi2djiIIJRyR448U
0EQP4st8uJ4sy0VwnI4YyNoIm7GMLGmPpfknv7nCreSB9yEZ/IYyoShpSJUzF587
6Hwcb/ZN/0+PaFWFmYVnkIsVa49K1GI+RXmNpB7AQbxq72+RMs9MguBBkCNomfyB
PlkNp3pOf9VeKYlPWOCixsap6uN4WALE/pO7iuKUTLEjJNy1b0jL6Q7zm9VHPyhW
n83wrodKKxmLyh+bZkatyCuvsnP8Mw3VvmNYosoChzTCFoyCatJByKyyNiCSq0ub
wWLFg9o8euPtswKAwVBUpZ7W/jW+373cEBWSwpSDb0fkM4NO1ZfmlWlbq2vSnRa2
jMBoZAIi9gNSSZe7tnTIRt9TEp9A5l6gJl4SThCP35EAxE7K8BRV2Her2SNvy2zy
LWV2j5NgV/K+iyHrcB5ghcIVOF7wsHQT8nwYZTTDWCzgdphyTXlbr2l0KDNvk88O
nx8F6PsQjQEN40GivWbi9NUpI8iGh0JLsr7JlSXpzCyYy4WhLQtglfcJCKK4PBb0
rHvIsNMjvHBtxiprrJJsyjGr72RPO8lh2yvRS3pn4ridu0L6HGUFl9I1ToSQbE4w
f1AlU4rAO+Xsdk8j7sK1p7WllfjkDoiPQB6HTQRORlQ0MSK8QilXch3LKnKgiGEB
BDS/Bfltv37MMXv2f2f9+4rpeDU7o7MlGjqfoDezao3F0wz/fzJtIAknk8Ih+gnA
Cnx24S2O8jAqnD6yaPG3oP8tr3w5iCTwsCwJpM1nemPoZ8X7GWVw7ZhjuX064J4d
01bz006Sn6TIi0NiP3H4mdsweJtV7TV8lxwJdx/Ncr3oGEuOdvLwy1/dalSYex0e
GgDA1VKsrEFBLMwpaHlhyojA4zLeL1viGQJlQ3AzlLJHtOX/6yJYnf0Y1Y+olTpD
+mO3P19lZNbFPk9WovjaMgGQkt3FSINbzsNrQOkiS23kWN9nIkXBj9apjy/5GJvq
42Aq1zX2iqKUDoj5xpCavz6A+hhUA+ex3nG8pRW8/miypnzFlHFEIZHEpQtnkOU2
nJQd5sjwfNVgjpL4t6GLCYxuupfqFyuqFnzVUo/mDRV8xPO0O6PchKjqhPA7cn6i
NtmVcYlCKMG2SKQPbjzLjMnCKNk0BUCpWNSK5NsPeEAmg0O3V9uuEiNiQeunIDgf
AOdESHlwOfgCFrWlrTDES+K6g0Nb2sKOauRqV1eh+exKAZNvn6jlB3VIFUmcViaL
QoRFCjCC8ZVR49zmShq7pc3gyFzh3tpJslhxXXmzPs6MFjWooUAaVSD0Z0I8VnTH
XP33VFH1uyvTJxOSRyUtT+NqHDBPp+Gth7/oirw7cIWEkmi+dj2CBxUW2OhjONVT
dwSyzpclGEi19PlXxbh/hGyeOzsNFXrAcPllucz4kh0sz56N3kZu9PNs/G9dMWnq
fnJHiTjGVJKD+TH0r6SbZ1vtVvlV9VBJLpC9qit57EuSagLi0+t/OcYocLr8/70y
qY/9zV0qsXEHPxXcju7DT2mY8hI7e09ylVhZBbetpEXL2v979bTp/qop9w7Tgo/W
bTIlUHN4LZMvqjwY6+US9ywPwIS2s1tDfoar43rvbcyjs+FjSyxyVBPDBclvgZQP
T/3lCmY6YYk33qmNVeAoEs/LtAddVYIzhr4FNnPhiT1zq2KKgQ6CzoV7igv+J/Mb
xiY5qdcHfiVNrse5tYKljZIF6aPf97x7kCrNLxqCXzNVZ91yLiipHiiiJJsyLeoy
RsVl0lU2MUQT+m3F+rpXiH5YE7vP1ilj0I3VlbHTqnLacTFWBtzuRrlVDmPVj9/X
ZZq8szf8KFAtRQSFr6eFWabISAikHbqc3/sFoo37QEMast4lHXDBYR1qqcgXzzjS
qb1B6iZmN8Z5qcuGD37V6oAytSSn1qLeKAhuapBUuGsTEFyDqPtX0ztZERb3rkvH
tA+T8gInvThL9GVGPgCwGwOV1XHnqUhLlzWVfYq91bvPLTIFcD804PrRPTof3Uzc
FqJKJXGNkLALVswW0ZD8zaLaDdSHqsJC0dk0ro2/Jm02bA6haQon2WUF7J9q74P6
DdTV9FP5keFWPyIR90aQCaot5hikWJSVepoZvH8JWaoVR6U54BgJG9ftI+N6+pd4
qa9BLxN4yFB+HrUfAjBFmgxr4qOpCK8+dVAYCmlg7284l4IIG64tN/wElDSjf50x
XTkBJYnUPNeCWzW0sXN2CHVYdRsW+BHgJNY8wbNzCgmxf3yVcT1aWl+whrRtEJcV
6zSWcOZQH2jDLhPROsBwvroUgrYYugEq87cUL1sXz9+FgOi6XHfl9FD/ZqxndARh
zHXFSrTsKsSIflevSeyVpYijIIoW3TEOIEN+ZTakr90vZhuhk0WNV0u6XR5j8Nbz
2RfcxPmxV1MTmpkqnyUkfHcfS89laMA54s06Q6MP4YBTqVL2EqPBU5MZffxm4ssS
D10BCfNpZhWwwGhlIZUnJTnfjoKQ4gVntP0xIwD9NeFIPzcusH8tFONDf1L8H6eu
WwfVAGaXv7gZHj0to8tW5dRsPpBpTtu4fzr2kO1CaGFh8vTzKj+7ctX4cdUELyj2
T4pGE5dO4VUW/V8vF1WHVQOH2eWc0KGKD0UWBCzfDbOMLgK/28BzYqclj0x3ytt2
407rK7fPO3gpBUR2DUcewvi4MIgAYpYOLfP448TRgTdDt35oRORuKsI0ApGxPFSS
B5i0MHIkNKA9cBn5X8y5AJLoVSZ1r/9Kj3Og1kJ3kYXbPpAF37Sb171SWF3B5vlv
1p5oiG8i+v630pwvVd+NUUfKBp6aWtArKhPyjyC1XWyCepJlY3uBty+pueeRwEJ8
fgsfsfo2JW8VOz3uPzhRZILk/bGlzPPAZvst8aFe2GMellOWaASNzVZbvfPZkRV6
fKLSeBT9ZCdCvSvaJ1vbUjCvg8qAyJ8CFdkiPVYyWKSO19xdl7WzPefdEYxkiDFU
2dbtuDdcnJ2hIoeLfdl1M8ryLYGNwBvA83gjm+B/rP+0xoL1ijximKz3x30CRNtx
b7cvGMkxui4tD6df/F4wjgI/Pp/xpmNwaK3Guq2yZaCu1tLvctcc4DpVe6UGm0oW
1I5s+qm7DyYYuPwzt7f23dZC1ssjrqDqbJcLajS7c8dkiCY05URHwzCPy8tMXco6
6kdPeYkcDXL2CDN6W6de1XIBYJDRObrSD/DJ19rXvaC//pVuCVf09AvVhr+RvfEh
SdEx8VikmtR7s40qZLMFPxSji+XhwpldBghsHVPIC3ywYLvHTeZCtzJOP9ZRDqS7
JC5c+AQpYOYKZ9kOVA9Hf9yflZO59d9xfjUQItV8T7o9WQ+d0Oi7VqDPukmcjIhF
NpLEu//ItTlgmocVVZyE1p/SBcU6ahhXV4KIzk0Ni4Dnm/SIgTL/MSafp7K80002
l1fgHeT/GZpr+tm2d/7frXedG9R7aX0Wg2gJtio838HWfjjYVMtyn1lupZQPyinx
g811d/ga7OkrDI5F3SPwhHufqmSaSl2u5nLB6cQ5vG3D0hms3SOY/c44Xo6/Gvr2
tZ4NuYJCjWFXeQnFz2RdxF09yGNnB9Y6H3Qk3ZBx9IsqAoIvcKRnxi07hSXrEp46
NVX1HnZNlN9Wcpd5o1XWFWoRpKLAJHJHRk6TwouODanJp8tuBp8ksfV0RWV2yJWQ
/994rT8kCNwll39DUMocTboApqXU2qz2lZsED7q6MuhDc547p9nRH+T1KR1Yt/Fy
f083K05/HkreCuVQ9qk54rqFdfCGt5DJzvOmWOVZ6J3+6XNm1G7nSKfsFt5C3q9C
fJxfQ6dV483GPfL7fYY4kccaQwcfOBAzuUKQutiYDZiVgXHPBfLbLB/pT1hURtuP
Kv97WhTfrs0Tby/BFUFwmgXiVJRUfnzGwyj7fNjdRFWCFovjOgbmj5iLr31Pz4uc
64My0x0xkO4Fy+OQfDv5/6DYkcat5aTja3kl4z6nBuzquTJmXyrmGxpoql24hqyP
6JF/qU8FHcAKJBjFOw61qIVoPFnJxsxaBFyLSoiO/APZIaXETz0u1sG2PWpSWmS2
U/n0mnsWcjt5YLfGqXSxMAhMH5MPfK35XWxcLV46oHWHxAniohQNfORMTsUWjcC5
8TJvphQ4KVrrylZTBu0eyaUR8I4PjTPaAnfS/oHD26gvSafszjJS/ocNhCUzXYqz
sZF4hR93/7cBaWASUzDb7bSP57tYNtT7RLkHh99g93mcNNGk4HgNPWcOnDQdwMaw
eUYDCZzKcfEm7+DkB8RzbnbUMOZXt+zNQ+VF9sVjc1hC8dvVRiAAEz640klsN+Nb
O3rr7dF9KtTwhaz9MHorUxcxIN+s1P/vdcJQce/qgdle4F1oLNTQ1yZ5i0Iu3MN9
5wb3zk1BapTTqJWcXCI9gLB1RAOaOSz1+pH0VpY8INvDqIPG0vhu3oR7n4OnDJ8F
zaxNxYLs2vQbzGRke99jPTpB0QP6vYyNeZDkHU0M/eRX8c2eAWEavJtALH2OJkqH
2bzMvVMXNaaWLK9ktuDMRZuYG+YKdeu4pm/pJ3djRy+REaSW7seINfvCAZCMOHKF
90CXSviEGIUnKKO5FQ57ieIaYhTt+Ke0Oew9/mWopMFgVUbqgkBZGry7Rj+A3kku
DOZZ8Wl+INnIWi6rKgQdUEXlZh26DsfZF9IUHnUb3pPJadmq7qGM7SySJHqmKB2Y
TwM77yCvh0i/oslHPBoeVKqxB5jMjFPAMxBX4aGFhgnpD/iGMdVeOAT/ECitPbMM
JLPFs4cvv+fsl7EmyCmPVmxjV18q3QIA6yC6DgFyIQ4eZTzkmPCGHsPKP0kwmCmy
sTV/1qrPsMZHS0KgPsQRJbonEJ7jSQebZeZW7txJeSLRo4YHRh0NQAGbv1vOOtE+
GOIh2aSiSvjP/7t7q1hbzdZxVMseEksumRtL+zyAXzlOLAhJzk3ohRbqP/BeYeGU
rQG4dIdGwT4pGjxji15xu1ha/PxSKfeEQF2LOJOH5FpMLitfRHhkNGIKu9JLSAMs
WkUAZa6nVaS5Rtd21/f1052ejCHNXzLQVqclKug4ya8ppnLHqmANRLhcdydtz1CJ
igGYQDD0Uql15++lbnuuuz+9IV4Qfk4L0x0LRm0PvaskTtrmfwuaPMUlx9esFRh6
wmuNn7r9H+/SmZMg22XqlUqjkqpzFwol8x/EBfPDeion6S2FGrK8G4fu3RVp/SQS
sU3gOHVTxNGukjHpLMbReSIzLfF0AB8wJB4ZZDr6P//2gKKobV/Wih9+b23268TX
m1siU0s4P3StTJ6SdQkJnJnJs464KTyxVH/sUcUp9Dbwt5n+HaZA9pzZ/8bsBXrU
x4Jam0hsHXEO6nQakUYQUQB4JuvqN37kVO9iQHbnO3MsWl/lIbrdUvT3x+CKOK0T
In+BLEzvE5enQLcAvUVFthfQECPWqCI8fKUPA4eL6NHCRklJvlR8DtIXWwwfh9zP
g8paUFpmrjJADuSSKq+hBDSZqCNK5cPBVbJh0bjFw+20hUq5Pu9JEG+PsvxaUZ3E
homgKI7YzS3UJURk4D9+MW/wPvcifHapThOphre4NA7gQAGOSrUWHxv7IYrjCs6y
aG3oYzihgityZafooXZ0epgHLAhuh8KhKXLaWT3s/s7LmSWpoCqX/qo+3+z0+jTd
dWSrrWlQCzm/ZwBgMewOz1FN7iApnQrr1q1C6PukLP7H7PxjOCbqfVBW5xpja7Nk
iPZE8SX6wcsQSRuUlMrYdqXd4Bx45KymCONvgQLVaDi2qSoKv4SRGOWkVL0RP8pz
vbbe52Owv6gHZYk/FYtjovXOxnPqHoDOIqC5dNssrkHn1WdiB9blhLejbw4IYCBb
34Lxl8hTihRRZbakCXpY0y1JgLf/WoB5IdSrrO7L4yHExl9DCJ85aUBRMRqTt1Ua
hMY73F8y5Zk9zgDjN6uZzspAx7KatYBMDFeuZwbMsO8EPyo5ewqGFaXgaKExFop4
kalLZwPHts+FpLmgh+Q13LZjvXEXTbo6fptRh7aTfcc4HbEqVesoZtYZRRkRHtLc
RWYPnGqrmQMQeXZKmrciluqD2NEP7vwNg+QsstBT76GGR6yWlC9nfiV0fWUr6hgc
KXJuWgD3Yf+ubH3a9qXyEYWlOct5C+OocowU2hyncCT9sxuFraRICMLp8153F3tw
HavQkMj8XsYHGhoxmghK6ygkf35MyjBQ4AUOeE199N25wVXUAClGMFiX8wGjSbBG
OGe85bw7NKr09sBF+FYVvh0y9u6IUL3VJQh5QmbhBVi6Pk5C85/pHAtTcePNaoHm
hxWoS/TBvW4pZXouA8GJ8vuRToPD1yDn/4N8Okw2aUeZQI9uvH3cyfRXDDNAASFT
AEKbCm5ptGA1i+pF9thp/D+i8nOXFCl2zXWfXR9zAa9cpyV2uRUsYK2h1no4pMR2
B9+cH9LT0TWcK6amhzTlBd13sxaiGJJV90T94n/vX1cqA6Y/uVo0dMFPecTESTPi
3ZgQ5RwT1T5NpAxpc/dvSednL+3mUzGGWVghjEwbdXg4PdxB17zsAQevXVtPP8eF
q3M6SY2ZE+UuIa3XsjNUthN/JgIB+v9SLxfj5FoxfFFZJ1ulROiPq4ZXNKrDgPWE
2QPeWbb6/UEudk0N1rHnlTax1dhjvirrtNtI5JeEVqk4JTVIZoxRNNhxITEBD85e
dsXxKcBmI+uJOBQUrKKHNY3MHCGr7ELgMC5Ilh1LQ6aCnnzjptfZ0puooHHUPb8E
YYIqmR5tQkDw2EIEj82XottNv4+8jO4ZIljiYl/3LAXf77pgRaKMeSXG0IK/WaEI
/ZAKRv6OKZamRqvD+mEhhNjAD+TT7HP/348qzYOMt7bG7NDhTmBD0fvurZMV4Hur
tcvjF+wB0Y+bdIvWKxDTnty0Z7vPN9kGP9G5skBovSjgGr6r4heTL9Y49LapQmzM
pCjjgvPhKUxrRPTXqhrcr/GXRS1pDZJeoLO2dAstn9x1DHFLoZrOJ6rTiWDb4ZU8
RRKQCbWkCo19qJOd3O1713SrlJ2ZdfERSur/uzQq9WUPghWjaNr6/mCHaU/Kw9tJ
1dQEuGd27wX65KVCyLrf0NpUBWMggzO8MyU4QjsGnZm5nVHQwHPbXDFCGpxhV/xF
DWYAwjdiwcZAKtpcO+s7JtL1o19vCzyYBpmu0ZokpiOyBN62vxejxy6A/DZXioY2
mM3nXDLjx3yAsAMr9CcvTaLOrLkAiJ63i21j0D6BXoxfiO4vuqUCUwQkimAEJqaV
HUzU3tBLHpv9Wqc1qlyRM6cm4YyQlUIu66t2GQUdvIzgF7V4lFp77g8iQtCkIcWE
jDgkfM8qjv918U6YOjQD4KykZ7GYyiVq3/eAyGwFzs9tdX/h/m34Wj67IgCaZymo
1QJwkGBCtKlVR0mrI53Wl4RV+IK/GCMRuWY7IOdljBXjgOJyLtrjQIkoECp3JPPN
wd3g7PlrS8vPZgyWmQcIguWvCfvEL6tpQdDiT2QSucjgPI+o7xA4apCK+lbnYTxN
M89BZfJofYqHrd7doO/IoCgp65UlWgXJCTgXYmlXiK2UedmrM2g9MvYgbKIWYQkr
yjCBuBVDI5f00cLnhm8LhHOGPTcMPuUTAmf7UekeAFerOI5OtdgRqvpoaZ5MJrPc
bU/uff/TkUvBw66jpnOj6fCCf3glSxlymTy9k9GI9Q0veDw0fWmsafAzdxiIw1nE
phh1cd4KNMSGIRZI/e2++97E82VVWUn+5LjOVQNgPutiM7WIMjIa7mJPM5C/hT5O
A0pjefk9YNoXJqf4LaEA9TlKIIhEnZXHd76figrgg1nsEWvnGzbYPTpMjPWI6rq4
Z0p++441y898/yLL3/a6hJOqHgWDi6K3wnjv4Pxmz28x4vzqAJU/oEHpGt0MNZQU
GN1ofczss4PxXIbbwcaRDu1ZYkfV16rRvajz8JIrOxOuj60zQTICH+oyEp5HvBJV
62/dpwV7CCEr/cO61LWw/ZHxN5HmEg9nYAmQCDXnJggkrENJLck4kkW0yY56rx6t
WN/VL9moTE2YlSDN3NpgYmgdl9Daw8yyq5hG7CBfrE4ov8XZlbWNynY8fWspAX6T
xN3vmWSz5KHPbn7rc8jXKpyVdihriK0sc9No9NGtKj493v23IhvWWqwLBhlS8Rbx
pIMyXCh/IEcNtSSggAKBPUMxHwdOI8VG+LPhuzBKTYZN0IJA6Q3eE+Mgkom8CqUI
bz8u/Xy7ScsN4+0jedSxpWcg1N/OS2IVv6yOc9ObQgPL7dluiHZKxQ5n7ibvOT02
MFd7hNltDCabvFjBykf4U0qxdjbsmKYe2VdH6eszLcH815SUDQ+rgdqSgzEPkOL9
RGB9Pr0PMwWIzhLATpiQ/8gQfRWCoXnKKkXMBLrHEGoieZeRxfIPNQMAStp61JY3
sF9STIGlUNKJdRY27UfYRqmmVByeMtPz1MPiC2ie52nrcSwK1I1+WaGRyrKJuN0N
ZUvvzut9IlvXT9fvtetbVLJP0m5nzaFc/7M9iE5FDhEbwK1O9tRTEZ0ojBssP5oG
4sQS/Jpg4fmuxSJXH9ipGms+oz1dBGizwiwhwW6hsws8+Ejg39mYkYewCJFMz7bV
ABLQ6P+0uBfuYhPWBiRHPpedmBXZY4qw50WUhYzPY5086U85uAP5YE6sdaNy7MBh
EPaWlcd1mk6Aa1YxndMqIq5ICQzefxt1Yx06NLbO81n7ofqkyDK32MkljqCNyQK2
y9niSMGIiGSro+gVDshbAzb2X+460lkzEvPLfTwPe+bPW0xp6/ecTCIx8CsMMMs7
rYUx7Gw53bAkaEFl8RcUQPR5bZryQEXT5c2Y516oFkE5mlsassY9lX4Hc8VcM82L
aePcZ9tcouBhcHUg75SXBbVo27EZG4I/9IBEgMQEpHCg6mR9PPSfUn8Hc7mBFpZV
nPQ6uZkR5DSJfWgia2VCjXAFuWImAiZOzcuZYCrgostt/CaSn+pkkX292NLUVQEB
lh8ShMvlwmCDFC9CBybGYUKIA8U3Hak58Fal8n43iV2RloLAcETAAa3gy0jJhtyP
Lkh6RJyPvTaJnxehiP3rQA+SDlaCmqMIt0J7QLuDd0lwjMUvF0OnkC8QjChrX1I2
LgSeOQ3Jr4qlvkgrUH0QQ8ehvFD6A+LkpY3ntLYuKe7tPnoQtGQuk4r9DPfD6CUg
K7xgOtdR69Gx/sD+xxOMRuutY2FNhW0dtcg1AW+GNqAsrz67748ILjz1ibrwfADn
MokF0iUtNsNSw8M3VYaUIt6n+reDP0oAayfHer5p/HI9R6vYHY25AaqtjGnhySg1
JdJ7Ad3O2nENIuOl924teSAIuZ4VuWfZ1B3/y8kuyBRfigf0/pUIpDhhxnRB1jST
HzGKCBVWQflHq+5O37484hDa6ocGLsWRjd/dgXNjwATSUDqsQwJ5Nz/WZlI26d2T
3lu/8Ih17CgKIfBRptW6bD9zfII6a0V5Ahiw/vFaf2xAmtTbng8M2iJXOW7M9tiz
bqqydQG9206hejlTQERvC3tEhDAjiAAup1/qNXC5QONKAzQrbobeWYFOf0Ghacll
dYn/hQGpd1yru8TPWj14O2OEuw+z1AH++ENEMF4wYilyNdh/8JPDp/icppy1q81m
P0UtFO5PhcOBw5rv064dUdkc4o/cfBIFiyF2Q8ARVzT+JntquY3+3oA7SYtIJw3/
4/UEBgp2/wz0o342dEeBg8TZoZ5Xt+b8nSO7bHVfAei4CS2BshIFFyBFYMqLZJud
qJzu0fQor5vqij7IUlekwNOUEsKQ+LfbKMVQs2FneYGyi2JM+mawYE31JxUxqitT
asoiiOI2yBqGA2iPG1A/rMlk7oYFn0oNpc5rz6dJeIRwYSgub2zbva9D4ExlsRjt
H11qcAbxR9xsTncwBBIwTwTmulb+jghjFF5lq1Iwzg28L5dmYYELSGIG5q4K1Bq3
KTdOB7FJd2LSAu2uAnZIRcRXdUmrWYJAHs+O04pYfqutw6B+tZDnSKDTMFatHAHO
qUhrbHIhVfnh0GkH8x0QkAI5Ie+yB7roh70pOoK6+9L0nlJ6bQX8eDq9G4+lLxpy
NurOkeszGCW7wgcWqNTJ0uQU4YkDmpJFJ18EIr90bZu2lulb9CiCecCpyUG0fAYw
Cla5+Q3nS45suvYa717mSPT+wi4dKoAQStPG5I1l8RJtfvOmGgozh0CXGq6BatII
niYuCgqMcCMokBPjFqUCOUtftdOq4JrVEtjF9+pTaCn1pttFf7mPrlMgNfbeUkp4
g5cb83GkWOOSL8BsDSA1GYppXTrrsIfGepHlmWgmxGyq9pGJrzIh3/eKanYKzaaL
3HJV0xvv/FM2V6PYvJbsaFq/fdiAd2e4LEQ/VqeO0i5++WmczbMZqlATMquxYTKw
U1Vr504tEMPQ72RNb0i96+EIefRrPMlCNY4peZ6xDzSMMUOsm7cVDAia/sHZe4jv
dTUtQASFGFdUxm+izEetxU1z1xPcwOpNZnHkGeMhNMOAMvEey7bKTltlyalLG9Ry
D0mM5BWcDgDFm71VWXC5oQ3iJ27+XNyyWYIKzwrPuMAkPzDcGZVJJ48qxo6zEcxW
13HADhpz3FtUtCOIKW43ezVfWle7sO/6ni8Y2zI1U1SpCO9Ue8iOAkInA2M+LKKe
JHSzpzKl5/RFNOxOZPX4bh2R9KDCZH092IG6lLshssR+pZP1Y1OqYzNa4O5aq8ok
eewlSJj6VgxZo/z2pNUqNSto2IjNtCk70Bsh/Ta6WORGTmtTfmJCiQvvXXD3Vldr
G/P3fUFJA3Ou3gvF2HLpwu5AHOEcDNGmNuVbUPsADlq4cU6TCnG1F/sUYLttDNut
0nhqzMfn3iyO9+Jk8bPyMtu92As39muVp5GMpTyUZlDFHT+Kfe1Aj2aUeotWs9oA
6sYupy6EoQUoW+y3z1p2JOqMWtoPEuk+yAtvamhBaGnJLPweWag9yfwnLM90N1vD
sTOVNJ+AV0P3oVf43Pa9LdNu0xhOTrg7bIBs47FHyV2dWVxL5a+74kok59XUgafL
DiUvQE39WEf422/Ud3y05JbFT6WYS7hWOHEra1h+HTRQ6eeEMZOAAPR+rDT/Oa3c
+H4DNir0RuOj8VxaVrSZpI9XabxfI7s0mAalXX9V58lhKEyDUD5irPC1luZ+0RNf
L9aXFnW4g4d5NsQv2zsjIa6yJobDJ6/3bPKlU6P+yz/gudKPMMbmLo2xCkcWgE3D
WO3ji2fnQKrZKa38ckV9PYLBnhIbYxYv5bN69hzQ/yZwCqpGbs0uScGUjbPjZvd4
G/IyExPod11W6eILd4PdlD34pMp8XvYM4d2EPRfkT0F4xcR0aZKrVsZVzbODPra1
NQJse14qVfjRHkW44obnT2xU2AVPqCbWrwKXGUe406mArroKaXMORNt4PpgR7wp5
K9QWNuA2kUp5ofzSDPY05pYXd2xR3Dvqtms0syRTcxKn3QbY7PiCdTXqE1bKG2fp
johDti6bzUyqG30aaHHpXP1rY1picM/RtGGt2gO3fbIWDmS6IU4EPqqnY3xnWZw+
W9uEttvTHxH9TPEqaI6AcR9RjsUBPyZlTYj5xaNheM3ByB10MZvC3CiaUXWk2UZK
G+Y6BPsCy+SElLYqHE90ioteB7T77l+4lR8twFNFua90XpMDDquEmxeAEKFVNsGl
sts3wbnWfoV0X7eckuh9I+Y4r1Q0iubXW9gfyT7mznm58ZldgRd3YG8l6PiyXnor
ojU5DTIZmBRj0Vaszd9Z2yWpT2ToOMdkCvTZ9qOwOsg7uq6Yj/ROsz+YWHRegICx
iujXKz3liErI58DQdA4DnXKdkVPA6xxHow/MeFeaqDKzmM8st62GxPGasFBuGtyk
mvtMSSRMCwFnVYW4L9AgDILD5h2XDABkUyiIL7rANxspz3RkISON83rfb5dR0274
zDVYGVGBbS+iSAjiB3C2N2g/e0fUap0xBqMH86qocomkS+433dc5KJOgPIk4Xszj
G2qRs+YhCdImH1K7+hTeBIGghZa03Hweieu2F4EdJgyu+j11giJaFVOYeaVPnCxJ
wGdbxZJSeJxBWR/eVD5/PETBAf3LdGIJUd72DZn+yxdhWG1tFKMy/cH/y4Nk6stD
VUh5hzOBR5UAPi+38osYzokMj1U/wT5HFZt3wQm+UpEl8MjVGa/Q0Rf9CYj05hUw
Gce6HACMs3PhHclMxd/XVZJFK2cphHgfCsezqMbB37DTEwYQfyXZnm/+rpEKdFtl
sl8CascpFntlZyhqJsm1s0vE5lkcNey6YAKeTLr3ni/CuRZLHzoPCfQ8LjOaV2za
4YvBNmyp7nZk8im2hKULAm9JzilAjFeCqsdNjQsrIpV5yJ3tJjlY6e45tGKuqt+C
36CnK+TJVoalmzkzKT0JKhJ+cL74+FvU+uueKpZyS047rrrXCHyP05ZEM7BxILHp
TBu/3TWtXVk3W+T9PBVdNvpzwB+Bf1uFeUyCz/DICz5cFWeVqO3gzsqZfI8KlAUH
wx4Y7I45OHibPYDGWv055JvPknXXqdHdV8U9ncuyTBZEyea3A91fVJ6hWk17xOVg
3Wq0K+Y2Ud+vy8FI1XPbJq50QB8ldmu1Cquz/KMWAJOTOA/WGPL8C+R/EXAyNXky
+T7u5AP0rDrQM7j7z5/z3g6jONCUV5Tt1056dvYfltZvXV3EuyDULYcZoVcXywIt
oWR6tcOMRgrKfi86j44gx/ks0RD8C4tMiiWLZ/kJAF2yyEef9y+FrSfGYX/79IMW
sthu8YAJW+RNeQKrhaBY3Dmne17B2dmQhpzjjn2K0vQqfLpUGVfosVIb81OBIGJs
bijT5mIbHop01VFdiYgHm2oDNSRx8+ghQ3PaMkRT9QGz+NM8VJ3fD+9r7YUsvvuK
MeFxOqZHaZxJKpeGdNKeWkPh/dIrotn1puYopxQe897KXLMb691BV1ooCAEDupA4
Fb3xXIgsalrMNxRKf6QNw8itzr9SaD5ATPoIGZlbsfdy3p7hsew/WNiz5My4qPiI
RugBLjqUzKqG9+ORzUJKxt8JZyK9qt4BU7CN38Wzuao367om4XLwCnl7TbSgEwr5
7HnAZ4PI6wzvE3+xIJKgiiiwQeqR+0hfk4/C7dv9JfuQqjSpGKMl50H+GRZqeN1h
OoTGCfC2Gk+8wy/XJaMqyPMTXW8cTeDd+g0jryaSOGmBVXmrZf+Rbuc8jA1QMnS3
kaKSqr0yhCgdOB2Imqen+ZKwcnxeYZrfiYfQMZJf86m/11CqO84v6Gu0cdEBeNS9
ONoNKUq4AbCAd7A++FCGPBXaWF+w2VrG/KMXO2cxWtG6MnSeKyL0uro+TC51a1qj
UJ4VJ3oaOA6R1ou7skethr76JSYuNO0LT+2yIeoelZlJfrATP9WACZNuhdUPQoL5
tKKqBqxDB5xrMPQmou4sTWppGLGjadm+fbk50NZF2OX9icJr6mUgH/W0L+mFmUl/
S0kXkP7cyqc/WtRRADlI+E8aYjFMGTjivGCSYgYE7RZuTKRG31RtEHHsfJqsGqym
VejqIUWs7MFCPfn062/pGg0o+3bNx0zFgjmIaWVRMZdgYs2Ts+2txQwFER31TiSM
FNJ4UsdRnrEjlDqz8reBBjaGIcBrnIX1/U9z8SC5sP3TIcNFBv0e5SfJToCAGJjp
h5m/dT0Z+ZwvGnzUu5Qm6qqFcu3BiNCQmdE1goAEUsQW0BzoohsWaGKBhTf0GnPB
Kp6/D/d7r/ayKuHVgP70YayTZVyERyRXE5ERUTnd6aSsjTowAj1Uhs2CA5RFZXCs
wiGGN5/GcuT1c9s93MDXupAdLBe5tuF66Zj/1z4M+b1D+d33M/kZVVz38XMWqnbF
TGrSaCd8dj9jWyknurzslTxRQwbhHXurES6GFkAIzV5TkliZCxgoqjDsFl5UWuBb
E/hdz0BNN8QSIS7NG1TB+ViOqh5kAZ+WYu+OwlmxyrCdXGQUxCdd/6+5IAVzRrgT
GCy3QESHS8L6QBYJliRdCZc3fbToAiz/RfMqecX4aFqJf62xKwYAnKt9f16Cw1KV
CdcNOphZDcNjKh70NTfjhxcA4dT4Y9vD/YLr1jI8ceS//uEI5OZuSskXr1p5/umq
HQMQjWr+wKUwA68D5K/jUXqIdPhmq/4ppB8YmKogQtKmqapSbs4QBcpdGP8+ZcU2
Tq8nRbLC7BFbfDgFwvAnlSDR+7qyLt7O55BbcA+nqB8ZGwdSA28mRsalMBFdXkob
I2wuYCBu+HYF//BkQ7hBddeA4oIk8msdoZ9zom08LdHuNx1VsVciZ8Dcd2Qgzp7G
yveiJwVday1xZxOlNkMzOz13ZIWVKzqjr7M8i8BR9cGrvC0NCT6UeDH4FO5unJYx
DJ8uRL+PjT9R4AWPz4JVNLuKtBseoTbWLkhVweAIKhi2TcP5xympWK77JoDFbZOC
uRVn9FpbbVkTvHrvet4Za/c7AfVMX5Fv9b5bdyG8GKHSP4TEGlYMBgGj9IOr18BG
neqfzsMQkfsqigrMsrpQHfhBxWaVFw3Df9ZIAtVR1PpwEB7Y2vQ+GZoJyWbEuVXL
uo9FfVrXxqX8QForf9Vr38PkvHCFAK9PVnQFTOu6iQIZ8nWcS6p6NrIOT+RNSe4e
yKRrikpFNuUC5woonQ37EnOMPjXgqNhEAxvtZ0gnY1N0//o86JEv0zf/U/yjtYsf
+NLwEpQS1RznoPvg6haQ8X4D1UqfF5MKcNf9BIXFaklSCnxOpGwSM9ylCO5vwWSu
SQjRhHc86+fDquaiKGN3T6s9EEfGRzjhx8M+1O8teGYpx2DCDkZXeDGn0t7OrW9w
jMGxfLZ7zHYbQ0RIvmLLXMO/t2XjXncy56rUySjeel2U5utf8VdUj9jpUywT944I
mrQ/FNmYaZzbYAKD7np2Z774U82CijI81vVRMvKFz7v62kepzWafHEzdVnPKmyCt
yCdro4K9cD5zwr0Xc2dfqQET+4+dr5bj+H/s7799FB8FiPF7706n1/aroHiQFggG
CIvLIhQs39dAEOPYM5zhkzJZdZvnf8R6+gmpCIYtk3b1OqqVjdVL77QIN4kRE5Nk
oyaDqa6+a7AhTVeuSVC6O5lyfJk1s0wxzYP6cAlI0xfZLE8Cg4u8RSdcofWnSJsk
Et8bvUwdWm5obYvxGOG2m267g+kAGgQrHhMcYeBpIj1YgRmTTy5C6vncJutXtsGR
jSUAL2fYDxV/joNkP87/89pI3PfUS1+0zoMHJnNsjEQ8YcR7pLM0AAHjR83X3xRA
xymfoxloTaT1u+5vbL5yDFlGBltnBG4Pjhmpvjs0IPdvmBNjHnbs21IBgMptC8jq
OITj7/gpUy7qrDKtEVKNDlqROgEXrmkUAr8OOxs7L4aNJDli71YxHFg+OqJrqZd+
VE7bAtWAO/JiE4p74bkLOKHZJJz7TfbGcSq4DNGsSlIW6q1ZdDp1J/+TlOgmCn1/
34OeGddnijczqxPrY5UOjkVVZ7ntCIizxE36bZrIvlh+OF3F18x+v9hp6kmvBfhM
0c/Q1m0dN3pebShD9fN6CcFnt9QGCtYPLDssTBzzA4Z3h59s3HDsAwlHfSSrk85a
rP5BavuF9U18Hzw1KSKW39Tzyc7/pIfzn5EJGFc/luAx1n2xagD030Orw9LV7CJD
TtesvTW5YygHb+mcE5KF8zDo+ukVsGRWFS2D7WkKiRWUOWah94HDTCm8F1aavbGl
AcNyfB36Ixbi4b+ngRVBKo944O9ogi0jxyDVA8bbiT64luydGdEv4IZJlbAnADLk
7/lT45mxGrZ3W79kVoAxciNGbPePgXEWVIlXfhfU3LCNql/1UA8V4/fdRyXtgR9P
M3Zo4YoWjzpvIvdmUgzy+dYNXPJPqT8HTBwAltSdp5yHfIOxDInzPKRMNvsdt3De
UvqVwitS+kIGkq+6r+HnlTr/JDjh/qJvxJynwntCDKcB5QQsc4eMP4kCXmgOMemZ
smsd2UY2q95ch0PrUoum4jVoFxF1iMXrJZJcqJmgXE7zp29CLxerLsRUHPNFK8Ph
Hy6NNmISKpnqUNMxw3esW1tSP8SswVh22VMOKosn8Xqi+6cM5/QqUjQTZ4znUR9i
8S8764iNimemGnwIN+67HlXYN3A5bwGgme6xIMSYkcz4faXLL+6Gw0i3yQAXNdwo
MM/vfVOVOTKMJg0zGcrHlYNzcidGt7qY1IyTPzS/ERuv+wj3R6VVzgDJRnidtiiM
XsKKOa7IGaRbK+Nl2aB4w2IF1kiSn2RtYKMMGjQT1acBkMTdu/G6MxXJe3oghQNi
mSdIkMM0Yujw3rFmJ1iZpF2PBUacTPWnStXvKPjz2c1Mx6qb1aD6emjGTGurDl1Z
xr6hoXpqZ3KTPyKLAy6EuERe79wipZlagoVchE19xW6UnZ6PWG330bpNyjX36eqH
97Mjjs1CzbGFWnfiAz76LRRpf4PGs1/cGBmPxCvuWs2uxl02yLK+MWVgXqEwC/pd
7A+tMQ4INDqcTnIYplJ9uQX6RXmiBdJjzsHvmlpUAHqhL3SFFkeVox6MuJKSiXoU
Hbi3gFuQNARITqgVByfpW/E8H0uqHS0BymbMFVY5T0aKkKULOaGYFQ320w+UWFR7
U2EUcteozHZe6sqGy5hYnXeK3SDnzqKAstmnEM5vZ5e9LhuzpvJXZ5mjNWSGv3OI
5sm1o/iwcQ/17LON9gdA9mdrwxIoncqncOOedP9Gzi+183Bj5caFZtOX/OeE+KKm
n9HahbQ1FOEPTStl6x3VA8fqDi2hnrt+g/pnjoPCzbicxxd6/bS7SwGC036NZgBu
s1Y3sN6n/XeC2GMqCoehwtOasI7OrP4RM0Cc+Ic3LFlCQp+be08riafQcK2Aq3dE
CHCTqd34xriX6FoLupVdDUz3SsqfZW6vwMEiRA9u7ix88ML9NeFnfwxI0RDSjapc
zshT5w2IxpZYsM5BDnf/1tc7jeeoIZ0mARYanRFmx/vxXKK9PY1/wadTUVisOKzr
pQrt5tQkPMdCOOPB+Y/uS/7T03uqQCdnRPu2cWQlwYEDqOs/ltDXlAfVA3BH6Zyp
8qsRnJIopZGuEHKzUG1T9TRwfn+VLjPTaRQiX0aL+xk0vrf9nO3hJX6vUX6uI0ye
5rXQZ4EUWdI1RjoARUWzVeisN9qpYZtiC8YcthYCmwMx8GIF5yBzEUoSs1PqtWNS
fWHLCDen7M7fFEt3B6KU8KCmgIQK/dKElZ5cO6dPJSykhe5NW/NyRkzwzdLdU32q
LXY4mdg11ZvkSNt2cotQhnZlwE/hbPeJSFZ+PVu8xsWAz+qaw5gxGEjyscAX5+Gr
ZoRRRCBGok2sNa89AbiUQNuuTNVLqWUWcEIUi1XFrmocPE54QdCNY0RUYGSdPaKB
lA+R4zxfiGeGGP03Vt5/ig+Fd06D3tY2lZMFmEUn6JBI+Apsa2teU+6NBWoZB5cc
B5PR3j1Lc/G7wNGee9iPtK8JgFggroqe05AGgaF+zMfPiWcqOSOPVbwPnAQupN5h
8XDOiPt4syifU3zD7sXHFk4utDPc4NbsAD2mbCypPobLj8c8hXRCug4bmtnggyFK
sa1867/FCvxiXGqdXn8gjIrmJsjpSzPI/Ble/9fmXNMwUj8zmCsRduSWVO19BcWl
GG9osWUybQMEPAo55MbmZW9JHHp6PM2+r6ToNNwGuDU1I1ZVUJMNeKeX4XDWcmOz
JqDjGYC62u05UHGI2WYWwDd4vQfh1LOQOFtkdMC0UcQTUxIUMrxLtKVVl5sK/bgb
f2LWGZpeN9XY6NaOPNVMvhcXV5HRZFiWppuBWfr4R12gtwyhmPCOVcpt6E/sc6I6
GRM0GrXRcCwmH9SVD8PN6sDw/BlJHjPsftjnKum3cHUXdkTDammD7DTmdWXjYCIa
1r4iYPvFfuNRwjUAv2tIAqyDP+wsh0beYfTcRnonCMboJxxgETbw8FPdwRHL9MFY
rALEcLxQRuDjndwYwAbPkTfX3fMtvxb+irvCaFQB/hmWexMk/gc/j7r+FGh5Np1A
bFbwbSV6sLLfNrD6ZTppm2X7h4xTI4HOW8lfxTllq2MGz7Tqx+jsnW336KYA8DqB
NzEWUTP8K2PWg1mvSzVMzPaNmLGWD53yqQfVpG1nrVmvAWNulM/Ne22Z4pEXV6c/
pvf4NROREUlNrSREEdVEwY5q0qw51tdNRBHfLrD2Gs7XW3EPVNwXQa/xdggiqr6W
nxsAG8CU1G8VjKHmsDR4Y0Dv0353VAK1PPdMoYxOLhUbFjRVmCrLKQIeJbzgKmhu
xNN1l47BpIp/CXnC5aQKDLL+3WYJBR2sB/KxKSq7ew4QaojpxapjWZsqqX6StB8i
tFDAYWPFzD/EyonO6K6iQ34bPfQpScE54WnlDKxnZoe20Ar1KsT4vCuZbpzo0dlZ
1spSw1Hr6eKt9kjAkHXYRESfvaxg+9yjGv4RioNXEON/D3Is+AwTu3ZUcjKHsO6n
1KVaSqNdv8NDrSH7RCd4NH7U9OXAOgVEqS35rOB9pX52fHOfurlNBK8xpAaQpcVB
MvsQwmSV1CH17zAL8yDq70Dmti4FIxCM3tJkPstJu5EA0p50utOMDUhctSp6rxEu
/paWWwNBEvUh1I1ykuUK9RUStsBfgBk6GOkHa/AOnHKtb1CvmWIKzfDO2wXJxR1G
6v2a6GRWPS2sGYHYnNwgL6RFVXkMimzyhtx7pOb7syex5Hrv85fnnOA+0kWlSX7n
ca/eQFO/kmy6A5K6lrrBhH3CR9opZ/0blmitxveyP+PkFSOlgM9IsnYtXS+JqoaA
4WVKbubt+EztP6nwYw+V0Fxo+M/7IFCqtk9REeY1RyL4RUgB8/7bkmXmZyxsExhi
VO6EzC4D2lDrC2y3+/tAMI1/9LK3UAevYE1MOA6OD6fQ4/ynSV8gUHK1AUJYJCpc
5X+tB+doIKEZAXaz/kqkxHMpoxCcDxTVw0bxnM3E+efGQZmZHoC+71IOwet/Bmw/
Fr0qwKSkokgoPeHjMHtPRNVdwtN1NRVX75z7KXo48zTi0I27nT5gkhSMNhASxQRk
NfM5Wn2yB3rrgSHDItFAJ19MPlKcK3YRrRhBHg4sBPr5biShkbbxvOtWjPuuLS11
pxR0OSr7Jt7NWRs4P0lLZQdR1n+IMXM9cEAXnExUjbur37A0LBeJZzV1QKaW9Akp
j0Ix3yKiHE7nxnb1U5hpHTdYJyyAUg8N77NPLFb9fX6p0ib2ECLbfkj4JpnCBKSL
xGSoi8FfGWAQTOBm2h5wql3PSymaDcUpG5G/AMmXRmdqDCZ9gpk+Jf0eM7NV3qhl
xiMQpZa3Cf/OxjWzU9+wbwRHpGW/rCPEXDnoUVNN4+HUK9JYgK/F//sDIEUPoete
cfdM8HqcqyRt6fQEC48PVa0PRdOhQvOwN84hNIMjmVCbGfd7m6VCKsIBxt+C57rO
tWRJTiWQ8fmX8vGZdQwtItU7U/qSGEdNUpTCrn6I5N9DKohsoZzE0G8+XVlcdWL3
CW+skJYme/xPvKCd4ycElukAsZSMk49AoP3KmJH9tuKYUOVo7ebvXTjUI3UJWZPL
20YgKYP/0NbEcZEspDZofSeU2H+Dq7Bhr4sQS6RLaP9Abvifd6ePZqWF58In7AO+
T8nE2Po4yM5riIHi/LFlFYid+op6PNwkGsEeJ90Dt6byWzr6nvwwpEyKzC738EL2
OHJtx2YDGLXoO1fzuXyqgK7crDaL79nThwQZdMKOWQSJWtVmORPL1mUJkcof6egZ
QhqNRx2pnqnsaYwjn7UulqGCzE/N7W9qv2ZzrhcRLSxplzTD4jfkphc/N1ISoSjd
/p9x3YZ7fLz4sxuI7k0AHqj6jh6AHR0yd7n9t9KtvpSs7mGGEEDxa7BbmwoBP/Ux
ZhLnMoBl5Z3tVsyXCVfasOAv/xEu51LMpAImzJNhjLlV6aAI+L6UzRF5tdgjWrSb
0XusjUHjearFDuvBSPS6rWlUqEzFHK6hOsGkhqUmqeg2T+q8o/R0Mm9iMpBy/NeH
ZUO6/jI3ksnjF650mRx/qFnnCgwvMuNF/1zVShLk1z6xBKU934hir9P7xrW1XQm4
sjXuhamBLArMPsUImc835xum9ZhMvm3+DBCHOJupsDOT0hgiwXHZi/3S5txtNuR4
ZRxsPA50iL6MK3XSsp46K4V+lDySgYYQ31z36otqgqJ2NyQelNv4OSgDXV2Vv5kl
4iQpJRD/eBUd+BbUl4URs+AwdqKoy9l/tHRitDlrZGoErVoGs0aFCs5nJrn2zyhT
9dxbgBl1ogy/hEGf3Ean6vRMYfgi10YIapkDk9TAqbuivcSEyB2UzNaC7te1hChL
LoNS2IuwnpJKRSU+wjp9VCLVAewsJvEgUfvq1+qSVXpQTCllYlsIgrIXd2ZHadOG
Vdt1oq/86n+h/DAzTmeXwmskoGL7Cf9rsXafXHiaQ9G139YJOs3t8VTQ0pkuaEag
3RRYuu1VNVh8uRAlOUnaSi3atnB2CTyEe0pSEJ29nIWmjMZRHjzbuhXWrN0RGXJa
azN3wk/NtG5rpK1sgWdV4e9DxjayHoEt+LIuTbRzMsW22aDAiiBtmqRszT7+kdQ+
W49192IH37MMS5RCxcRBe7l9GotMVdbO62AaMPJfLJZ6qzxNG0IWntYdPBdJBoZ8
vGBV96PozMJPzhRshwfzuLEYWzjjt0dFIL3j7kJnf9ys3lZWY2O6I0o9CKIIqa67
Vqc5FPsEz3WMYFmeZTXdDyf1t2Is7r/2ynMIiKK1c0pn0YU4DIl6TBQLJ1FGAtgF
H9Rz/cVsG9TkVgwlJ5s55/lNOB5q6+oh9nrudviqLQYxkYudUXmichIr0Tph66fp
ddAaupsnYWrFg+N2w3mbQtxOeqFNwTJxCalcNBomTe2GPwBRbTUX33owuiWCpSsK
VgCQmxh3J57XmI/E1YvrR/jK5DiURVBGme/3M2mbVk2Xh4VZDWmNvAPLoRSLmgUp
MWmWnwhH6rLH7PLIQE1kO1zdCYqFNR5PzdNI0dh0PvVAggkWpp1+/YztLZP3AXRH
ZjmPPfW4Wqq+ju3YvyseOUFnbJ0DEoN8+Nz05r9dBDU4n65yKQvR17hTVItseMwl
+RT014tM/1D7nIFUgHM1RuJLT/eWLmxIN5lT21fnFLEhtiw2yyLcWf5s7wIg/fhX
aRAawq453NGOr6bZdd0zMZn3lTqWK37rcowyMlIL2ag/AkjKCRJyVuBuE/IW9035
OM+BKUjk5rXnn96gpJ8tGmQzyHsZajGvG5nwcIpqmFhFKpwG+gG9oYIhZLJRZe1+
zNprPefYEoehqgPGGj7zqgs4/q++BMeAZzMM+BjKOU8SC9uJkUW4p33rxbqq5byA
qyukysI32Ubtusw17oFQrgbL4177xcT67TqKe4fTNRdBZDHsZs/OvMuzKBVTP1/X
S22GEq5PoBgr5MKX+KdI/mqztmLq49aIYo9aTqMzY78narAd6/TCvvCIOVk15lEz
IUTCcdJHyjW9KGfizEEn6oZi3WdedmYGKnEtsxO8TgylPcn0OnII0P/x7w+5s7QO
a10xAGdsODnWkyDyld5+Eq4Ta8jl/p/9Rd84QpWhuOxxHr6pFGd3m7oa/Kh203CE
0p/+nJdDBp8/JC2RbZiAquVk+USHN3xpsbt/d7Ru+7KznfRioNuY2ABPQ3Z6tKwA
njWRQjIzt2JFzf4vyArdoajVr44PJHcpi2XrLpa0c1KrRVu1DXlA156J9eHOyY9s
0fAY3ZA21jF+hUnrC0JdaBJe5efVwZzP4IzdbT3Adn74L/B1ZFT9Dkcr3/lFBHKo
BvXbGccLRToRSrWUlOI94powL5SVNe0o6ffO1Tm0/ZoMZLexmhZ3YAM2wjVPhK9Y
EixmjdM2KyXu68YojbdhL8JxpYrMvcfLhiao9T8MhL8Ah9zeZRbB3WPTwnAkL/Q2
R6xzThLE9Oct9nQumzHcP9kEb0TU+k+09grumAjmAMxaCNEjzOeBgRpYyXF2xQHx
YF+23aKLgetk/+1RpAccSiShgMVAocNgt884+RZavY5gdkdm4PKL92oJPgK7vk69
FaDUeeB5sCzCZ5+hYulYwvd37DLDIRYgJ/4IDhZt3EM5rABeHa90vKkm5o0vSNMr
O7xxpvrI/acWw030T9ZwKoVKPHO6XgnJ3xG1UVC3yDJiwo0FbOHFy7XpCmNJZGml
zJVMqfDwmCNVZI0040Y/k+4J/FzIHniWKKDgtgbdFA2WZBb2dmPq6TkrmOtahptw
FajNdBu2xAoXxinhVh+4qIvlB5Wfg3Tlo4TGgu0s1dXqsb/+yKH+iIP6YjKKcqYo
hUeKn7G8crBaVMytdCCxp4fAVH2dGrcPSbxT68sqowULB7WVSN7JIIlwammhSP1w
ogt5aC9uFrmkB/2HqmhgROhISiZiBo6lsPrFrz15RZVHJbyBy+L7GFFmlfN+qaiZ
cTbVRRZywqHNCn4lAVRM9Xqf+FXsXVGf2DDs2ArCdq8OJ/i1ZCfiz0bNbvzMGr9k
SPHaj3nUrVFtI+Ketzpqxc8npN9qhw2eXIf2N382vgGpfD2z+avAbZdX4Ekkni5r
0BzG0UwB2LmqyT5kCimwKKz9HsG3wAw/iEvE3F/dIGpWc34Z+Wm0s2HEE/njV5qS
R4qZPIbW9bilgjnPJxXkUdq/NiK1G++GxXcJHc9pqxcp9h7kRMThNlfS45W3btMq
G0Lr6sWoewf7YIxd4+GnZtQqGwGs5i3P3dAd7yGoWLDxsb+gDwVkEZPa+Jixk3lH
bvHPn6ahDLQ7WZ4CdvKlnAzHSMs0fUHnh7IOtxMdE3BguxSpYVTGVDz4+6IGjYvm
4Lz5uQ47PaWYYyltks2sFBQzKyXfCIe51neNYc4TpBzmFfJ/c9j2ZWMdCE230zHE
FcANCDuWgl351+LR1oqQQhO3eVbpnNFkAW6vXhyQ2sydizptZ/eQNsMBdFSufo6h
+4UaAaG3qS8cd4bG3Z0/fZFfw2i/rjviLHtLYAPhmTLtQxgjKTtWSUAB2tskYWxv
O2cjZH5tB1vmpJ2+jNFCeNClQ0muxRUeDkfGvRBAH0bBD2erk8zjRKeRLQ8vz02F
jDjbEaLVytTMfddueCF01SASgSnpgx7hvzwGbyCH1uSRDg8cJ2H47Q2TlUwxYZNI
6R48qGEAygHjWFiQgCnNh8rjJS0MWYvhrgEC1509gVmvatRHgebJp9E+3dNOOgJK
msuW5e0bDnIkVOO21XcfPd5FzNZi8mUeK3L4+3lZ2nA7H6NJIuPbIjEQhK65FdPG
3wqILZDFB+C3QxOnsXv37lPCtyteyJ1LAHamT93PqTTO8RDn0c0sVrTFtZcHs/4e
zDnbxWlQumdjQvnnU1FGAdw7RZOLHa0GMZpiKKorlEtRHGHOlg5AL/Iuiayg76Aa
8rbAMvJeN5+QzCxvcV96VL6mBUedJq1g0HA9kRI8zZJ6FM5nN+UiEAiZSDQcJ/hW
gva1w9KmZaMjypM+dxm5/4bnCjTKqe60kRtvRUtCEZXrQScxfnvHvuaJoBW4PPzb
koSI5Yn9ZFcZKCn7bsHLHK8daDBcbbGabS5LLzC9mQT8Dpx1zmYWghY239Qei+7C
rytxEH6oomS40gNNqsAKe4wKPmFvhWhMFL7BSccSeWX6WckUrNVAPioiJtcqWfYV
qySFw3tcdARjBOEj5EY6po/8UtY316kdLYXyxbDS7Z+eUDXHpltk2d7nDtnLWfsv
YpUXY+9l3TRw63vHsq6LKI5CPDJvjccfOKsWWwBiU6ePwbljavtVW5Axj6fXblcC
0meZhtKCxxu9kBL0OhScvV0LjXkKBfmrC2d9a2iOOWHu1c5PmeOilOTgsGMYSqlg
2izW7j6tkF2uUH3gbcwnz6Y+CwoFn4dDPn3X6uV+P5paYoUvW+7A6HIfRshuYt9j
bbaWWpmCeZvCihwj+8nBXzQr9wN0ju6Pg+njDX4YIqCkkACIBb1uPUQwmbrtv+Ni
teA9f2vANXVSBIQw/gtHB74KaXNzpIW2J98k2AS/2VBnOypgEnjY+xHEPePhRccZ
2QvFE/79eIc2FvggNdtSkBrsXH1bUYAqJEnhuP7qdKHW54+6LAOyQZihobCfuEeQ
ethdW2LZDgrs2l+vgZaTM9LOfUFI9qqXIElqXuxmqQojepTP0ypOA6grq9gfO8kX
ll8nkM7jYlWr709lxRHhNII14NlYlclesub1wlgmgtfh97uwbIcPCW6u+lmupV4d
NZL4Hwd7Z32guOsr1IFtM+/DxbBwmxd0Zthihe9tf4QrWgTqLF6BTKiOzIkJZ3+l
A4WsbVbLbGPCaLaftT88WhIboZySbVQUQU/Tl8x0SM3yrSb8MGFczPBcyRgrf/ol
WqCwFjBHfGC0Fo7o+ZiZEHK37tzmu/zunjJ5qxi32Z6bol9gqW3KP/6c+nthw6e4
4EEbYLTUXPLkRUMAYz338E5HOoR80zcutjc1w/gpDazJ10nE4TUAuFsEq737sjTF
1Hgm8bl0zBTCzQzla4+DSl9eoQl+6fbWyLCk3WhM7I9k52iAQKwYnb5FIczkSBYA
25UPyNxLvr7yD3fNU0PPYBpE23A7atAdebPdiI4XxW4Rdg1GlnoBrIAkkSe/h11J
gCCrHMGfCgd07Y/Vk88PqqGKo8pwo4ProB1yQBmKYx7P/YG3wIqE1GsBJBOuNXDM
5esXQNfHknCtFyfER7DhAKM+ucdpBalX0bKSPfBSdR/sGcBVgeEfHN6Oem8fhGz0
JPFneU3vc18vua8ZHVwH27ybegTSuPlUfehsyUvM+q47+m+P3pgjV3HeThEByh2T
6Ecnw/teBlKNwfa6KtKKTuHHk0yZ/l05Hj11XGckJVGV7a1Iv/7L84pmsDYz93gp
OpVZ4lM3mWXlvMgBkAB/sBrT93iC6yYGaooez4geEgSihbFjoofnp7SIH6PhT/oY
b3hMnHXc8VKyncX9jEr47H0e5Do3nIMYyljnnyHdnSqSrJxUy1LCETMebMT4Oc5g
NsXEbK+P+tK5otF7k3xMc6bHMMZLKIcajTl7jOOPeouGK2BRqBun01EGuSwUI+1a
1ybBwPFnkoistY8dqM2JsBW9vDsozLuFesOs3jyP3IQqaj7NsGxGyRhfJrZZ4Mmv
2OzafPnJv+EVpZ8TX52glSRPjJtEcl1+/gl0U0KcAod2u/7jr/1pSpJHJnAY8OYt
1AVjAlSAVWHcNV2e5s2nSq1BP7SikCvlisk7B8uC9Y7QpPVZNw2L/YmMQ5mju5Lp
QR97AyCud/cKs4t3OOgePahcKhaVbJM7f7WCDWxRULIlVduaK+ng8yJtD+VzMBdo
PusW9GAvBqjC771AmAs9A8dRmGkLcIURmb+w9Nxy65yulW6+xNRYRbZtN6r0db/a
2Ix6JfI7qiIyOV1VRKtp49hpM1oQ0bcgwy0RRLMp6fFeYncL8C36r4gPlhKTn1i7
/grZUBib7CaPvpsgUN2XRHLKni3f0AtopoHzRvts514TH9BLKt2pjfIbu38ffeyU
3fVTb2QbgTq0A/M24Su0NnfNAg7r3x1LU1H/2tkBpUZlD9duixcfVdpY0xejS843
LVNmxQls2rlWE/lW11/Me1aZOY6NUAyEWV6/feYAZ6j/sxLsJKQbvBSs0YJXuL0F
zkywYuENQtgt/KDyhyT5RDlhN8eYXYvACcg5XuQ2mV8YhlXo4LHhmHpgq6AcI44C
fByqgZnhJHyjuUAS8MICcI4xuyJTA5EfBx1VdaFgrCwtuoSGcxaKhGpBnptsBYdz
gQO0wsr23REiz84M/qnOeQO19rLu6VfQedayIq59aJo9cJ5jIZSkABuYfuk4owE7
kt5nyK/+/8nHK71h1w73T1jmYnSwfpFfcwe6l0570uJUW6vDYN0WOCTLJYvpNkpO
oYzQH8MVEAIP/7OJt2AL0+oeTYRuXAcCcHxfRI9I5PTGjkgiqhhL595LX7yBvorV
ucfc3FBcuZs6wEWcXYsruRo5vFhhLJ60hB8BRNptg1W8Zq05V41i14TedwHKY/mD
KXzynr8jr4guzRM73qrjMiAD36a/thwtjAm0mkAc6W6pCVbgE2LOjjQ7mIiL1jcB
HF0/l1q1Vo5nNWG1T6w3tTCGbDcuZwanQZ2Il5C+xsdXg1UAKoTdzq4GxTSLvcPN
yTQtYWU5q8KQ+NklqRk5bPUm1F7uScbHHO0XocYuK4YprTNgygin98bSlXLcz2g8
UiBUb8LTxzz0I7iqFA65VXpPloIPbKl/2IQUyZ+EnsRLSc/ee0SrOyo5F1fZQ+83
m65gMiOFy9I2w0BSLCCEBbIhkc+9HJ6wTmuDSdjQx3qa0ykb2RnRrMfevWf+BCk4
52m2P8FN7WV2h6QNZax8slxmW15vdkE50C7YTbPci8AynLnujsBt2DZFL4lcMKdy
GMR8Oq74O+dLzF4wid1cwJzcAo+jvn6vajz72bcjf2JYFvzLxqhJdoXTrj/M5TqQ
ARm4obUGZFHZmo8Go4Og5+JHz+Re7SpoZu1UOYXFB2lYnolm9qkPw/+RTGwMKP8+
lgQQu/mdrm7OvKIEfZJI0N4xWpFlAjbwYcZpFSAoy6hqPfI/Dal27U0AWONtHde/
6Fx9RKsSehvxiCzGAHopGlSCMiIQrSLbbc7CZ8MwH7TDHoBwV2KL0y5q+hxo9UWo
i562e2BBRpfOrh9kR0HT5+9JCJaGnf+N9gY4DyafWDFpAYzQ6+NL5S+wg773lxm9
Mm7b+/GRqabx/vYmpWflvNJhLJmZ9P1hDAE/hsowtjyHrZPCOF5uxbUXjhGppP48
0hgODo0YlSSBCbo24b2H2O0LiZPLwypNx5MN/BnABztmOyCnCZZObnjGjYhWNa0n
cMxjXw0Kb0WKOmdDp+D5K2JnQFi000ksL1dWGHlAp1CbN3deRIcuK7kP6v7cYtmm
dKxsEIvq+kEsCurlbVfRx4B3yXQ7SvdWV72XNOIAxo8vRHAdChIc4x9nd3A6DxrJ
WYU8sOURI8cKhg/uUnsihmE2oswkylXPtmPk1xo88sFeOO6ILEglCBBorWwjerMf
kIPkeyMNlEx8lSqd9yHXPfgX45l03BqrP+adyLglZ6Mk1EcLcu47rGtlmlP5Sp5E
b0GVnkFy6B5jCJ7TPH0LRQfSONrZGHMv22R9Sq4/MCKc/tOGeZeiI4WWkvwXcJrZ
XmCFJwLT/+FbaLuQ4dW1eDtrt2ihfqcVQObf/WOhOupZsjKmX7dScEY6x+5sdzJj
QKddWpHEwEFgG708zL1/qGi2CDpHbFrRy3weRwZ5lLZd7d0TfknrEpglCSTrnaqP
agoOQp+yKEGHFuuibcFz/7+ZHeAIsZI37bnUwyeLIBmRXGnS4QsY59ufZ+MgPYwN
3413WhQVlAB0T+uEZO4uiuFVVu3KgrSU5sjoeKwpRvfasL5R7TqG8aJCYAOGtLhd
6OP9huOv2qwQpUBGSSrXUs8W9wZzcu7Z0eULws3yNFlYSkfC/Vm+jZrMmT9/MSte
BX3VByAF7d3e67Bt4+Yv29suzr46HNWxEZaD9axC6WZcK6WRBFkHHR6sgqpp1iyF
tSGLKpF7pO6XnEMiMH2uSE/8SeOpA207PxyIMscxmcecjlV17gm6+IAMEaD01Wic
ZdCNLu8ZYeCOshWWoN+BUWCB/YLvDHFmC+ASUuQP5HqOMJNVH5O3cqS2PLfcXMwK
FvaZJipGHP2ga7L5Nn4I/QvdG0sm2e/GReZrlZsGXkFIo+OLN/k+yFGGJMM5xHdo
GYtdKggqVtZi/ji8HCXofjwYnlu4HiUlRZ4agH+TYF8dR3ewBx+WSy1qpnboA1Ia
HrsjYxwIl55FoWtqQmsIa4ubgdGD+XBHDYYsEH2n0fQg/DCS3YHlZPYs63LW7KGi
9LYlKdeQF6P1czmZlHi4b+IOsR5uAJ4xU/wO8hKhuAE/5mRRxrjnCN/RmOyieBLl
iw4IdwDyeqECfg9nTrprFmH0QwF3fTIOKP/pmZKmiHeQILU2SB7E5q2R+iRw0UWs
eAIjjRFhjTUC2B1XxcAxx/YTRK1RCfbHObaoG+Huv4NdUMeCIk/fNeEuvMiA3Nex
T4nSfPe6ZKlxTnLGdvPjDYG/mpJhVEyEU/X25ZVFAnH3Y7a59m58nj4rlOQ/sW94
U14XwMF8szED6rIYD762PSh4Jm2M73C21B3pt9r3QNYi1RTCC2meM36yPFn/7MD9
/eG8OXVHM8ZZ4yD0Nv7fL+ZOZ24Z60vGfOwWTgx6ib/lejNI4LDnaZNRy5AieInZ
iey6B/dxjDoP0gyrQ4qNPLSNaLHGiI43QLwpUNsXleLAhwGzxz8bWUTr7aqJdPtC
nOBFHLUqL0l6pR+JaVV3wqwGVz5y5J5yA0yHQYVabDMI1fwBN9+VeOCWHuR8pCpl
dmT5M/qPWby8wDlrlXXx33gbxSS3vQ1X+2l2/tlXwh9I0eK0yfoAPSdQoWkWvqpr
U2A4Ihhw9VXu+YXMep0krYW1DzIagtcp16yrR2bJFcb2H3svImr6bXzbtHc0Twey
wT+6ujAAHV8Y/Np8mGyqWwCINFgPZVNlnqNkxKfIkfaNCxHSHLjwFAU457OatTZY
JbtNaJeMM+deG2KwvOcXyqv0dAaUMbt+3CyGjGBxXOIXWCQXCK6tELmjAxnLujxd
G0Mv4Bxhd+l+xUe0xuDYnYUCK6eCqhKSyz7JoT+KAC15Jtj3AA76Wi5WuSAVmBLZ
yYnKBqGM2f8cdAO6wjtleO9aEnqRFchM3Yz2L744h0c98lz1Mpw78DomF9btFyEv
XqmISg0cunv3oNXLWCycLLL58k8pF1kdHnQ2ApD/W9oUo0ke7+prVxAwDVRVsImM
lyn/TGTC2zM5U/wkM35hucO7NOsUxE2w0Skr/hAGBLPRsDTtvaJe6TubVLpW9Xhk
MkT/oD5D3Pi/wWcy5x5FIKkB2uWrW+zxqx8SW8BBJ9tTIg5dA/6NQMyV+K7cpq74
/4R20l0hFAB4gh8dvpBI96+/GqCfRsnkgTvg2NZ3Ata9u9/kNhG3yF6aiaXvydsr
Ju0GjRsFe4kqxhKjaq3t88o5oz1l+vpO3ltTQj2eTC/cvM94xAMNUdUES/LZF7OP
63X1SO+MNy2UhLf/1QkKG/RwtezSvCkv7dr8UIuI+3cO1aMiBbaHdDGLGd6Ebwpd
VRzPaCrxxJYAY91wgYt1juPBxq7QyRibzWtyrM0GtoDSNV7SjyTUWMf2WtIJV+4W
yQ/MoxYeG5ibQrb3eVyasHFQ7WFshw7WKb7KcaRP/A965ztUw/DA5GwV6Bvb4oRs
Jb46UWIdRIfQJuMGC+LnPa1/IBgHym4SqWlBx8TXDgkoRU+CmqKHswOYSsZUX2OE
A2KOWlCH7U6NUfCDadqHE/yYwuTpoYrVzUbXouve63fWnKX5cFQv2x41NycjZn/g
vftx7tvrcAFri5L1yPVEn0vtjHq5ICU+fVAoicLiwQHHLKku6WNKVNQPRXTQS5pE
hnHPORUNvxuxdqaRgLoc2t4M6+1/fnc6S95A3tfQ8NatP+/Ayp+HB5yIoELsFE/E
iL4XMUWvBBot9lB5mcHnudWDEAjxae340KHYg59FfpfXzs0Vbsf4mFJMd4tpi6J5
VIyVMtcu7TjvKrSf6gNgNZEee8l8P+u2H2FdzXMGrGzw1cRTgdRnJEZyewDghmmJ
q12oAAdEO1ww/ruQNGz9hSVIncBLEJlB0WCUX2H3744O06ri0tKaEWexnIPnhbf+
nmjbonmxCF86cHPvpNX62zQVKwMpRzhdDKl097Tgq7dQLWVWH9wzL8frVr2iOmS0
UmuNyf5KosNdRwyiByJdBC60Id6qWOBM45k52ijE+Lh+kf+BvslBGo4tKUCfVMQs
x52273fBerYscrlySXBGli4wtNHCxQG0gLg62xbbJVxxxgPrcYVWAqUgP5XL5RCq
CempH3IkfBBUWJKLmnMc4x6q/iv/J/G7SwAJyeiMlTqMQlpP5HH/uAJhSbjj4jOy
LzxG15kLHjkS2p1GjsDOUK+IEVI6lk8x2y9URAzm7Nq7a8+XvwPUL+llM5BE1JCY
xA6T2x4vj+A5eqeSo9stE/ycgi1ySVkA8RQJH937iZ3z9wj0wP/Oj0n2NgW6t9oR
eOSAaasSTksOM6PTXQh6Em8pcMXyN1aAsFzA8qLr2jKu6rc3lM/ukYFCnJD7it5D
O2j+uTUWNJNhdma/NYJJEtfxmvDAq27PsN17BAXIh5Ot2HaZBhENXho68fdUiExa
1MhZSn8w3Z2eOY+WrOrnCKHfM9wx7miDPQsymt2+GnCH5jZjX2gRwkxzhKqSd7Yq
0akJUQQLkQR7kTjeJAwGJANeXGkoGHJykRNq2JQdbFX2bgpS6qiL6NKw+MIQVB9W
T0TXXawj1qhOgn5ZgkHA8xF1lJxlWqPzhIHgJLycEjse20GIKlTA5RDA2IHlYwnD
mdMomnV+n+Nek8TbEPnFy6jaLct6AJfM2krhaK/aT8SX1VY4vNnlMNfEG6Kxyw+t
tf83bs8XomZOfs3nBVvrl1B5MyuKdMj+FiiUX6yNOk4r9evm2wsi0JOGIzAVHWEj
7nuuiQFm8FNXLEk35LxzQ+0K4CN2HyZpmShLQIWxvBjHBOqBvXHAcK/lEVmbEfMS
/oV5dZ0zzzTNmoRE1rytJJxG98hRsWDWzH081qCyyBiihbCT67PKJeFSkTC6+6eW
vdOPv5S1zrlSZChaaxwN3vNld+zraoUiC3RATDY7JEzhCS/hXaA7MEqP21g8hiU0
mXV4I4lfBMZPTVn6IClTmvdV55GF7Vf83p4GcEgNFV/Xxh8r5u3QqbSjvIRbBnhk
DZlNDXdIYtn0KDBEhCcbSMLsCOipIOT7n9y3XiE+hISUlvuX+R2JUR8RilbVtC5P
4Mm/Tvuq40oD3bvyZHKJOdr/bILkCvMd4DjUkwas4ilPkwecruKrAbtYS83VFynk
wgd4ckqoLStY2O8Czd+db4zxQ25OJagrV9GicXKhg/q8Vl2hl+yEjUNkpEpf/B8m
V7ysc2z3xXoH3Juzh58NgYP9VDVgV9El56VkLutYdEHGiUe/ISareaURFq98EUEw
tL896XsJOBiz715ND9ICOAvF9yuzzVLiLuKF+guE+Rh6uWFNLH1JBjPx8/qSyiQx
BAFhYuvWQNMcUc/2jkEJM+d0k8lGOtwRpnIldSNa8JHquwLJ2slBrdr9USTj7H4H
MkE2eq6qHgdZW7lYUj4/q5GDCmTEy72G7oomB3jWT5lwuolzbsa8QUZ3o+qlmQIx
uWKvJUA3uj00/sWXmdprUzX8zbY74FNEHCIvN5AIxPu7SQsfWk5DnrRDTpqkLjjM
QXooTXx11vMeitVyy8Q0oR178DtcvyJEBqbZO2qdpQMDobZGEYhWANTWh+ZtBOpt
HqZ0BM3odMmESy9iR0c3wYG+R54vfELueJMyjenf1VvIwMt7AvStnQUzaEht2REd
12GsEkRm+1r7mGNuX+RcMnFmudKLCenawCUVNsfH++Jii71PEUL63GnnipN/eUll
Jt53zFh/F9jSelo3/gM5vhJBsiIHWmZxaJCtTbBq4O6EIWv5xnI8EUc/B+EG27U7
0TYF1EMc2cYqbYIa8Pers9O7qNCEHmZFN12+4FO8MFE+RSejAauChtANRu3AwRwF
FJSWRvKOIVe5BcavX/lQcEe0L84U+3JMN6kZMHS4P6Y+cowGghSXgMooG1NXNebu
RGpkDPwoyBoNeTbJZNyU9nw5vpqjcYumz2wMQAUHiaFHkEFdNPTrZ16Mmzv7dGhF
Uxu/eudcG95ndwoVrHBh4MlbGx9b1AF5gs88xIXHf+PWe3VkeylHhImnbgBHxeiP
fRo26Q783sip/hFoR0qHWVStItNYfNkcbn7oAS9VDszhTyKd+ElJ2Dba5SYpTG+Y
EFe43ttTat0XVpjv9spwklNZqPVo2TBfB2gNmvsJrx/DqUJZthLTcuFP4dEGryYp
9n/WjCYAGDbH6cdMA2IKKC4iFQUt0i+9TwCG/IkFqlzW5YE+iHpK77/f4Kk1fQkH
BKVhuD1j9b2h1OXgv1agf6c9dNYQMfmro1lFkNXOadT0oxF4MagI1hK8LyYgwe9y
vVvNA7jc1IrNNFePdlHwbFRm/fiTneQn5XweWKkWsjciJLpo2gq7I/zcJb9OVqwj
SNrnlmVadaNsTHiBKSF4b593wuu9mjat3yxXZQ8t578U4Q0ypfz8b4TzJmsDHMPG
NDCRyE0UqBt61xXUVuD/AaZ2wRaewSfH6K2mKwk7SC2+p4ojWfIagq+E1KwwysCm
aCFzCp4tnQz07lVDKt19iAUdty60RpUEf8DDoCvf+XipwT8xd6x7nRJUH9rAUKok
3uYsFQNjto2X6Rh5pmCIV+mDG/roWektdl0GVYg9DRpvkpiohK/TGq/BMFqCC91m
daUBX/mHmnGQ6NgkMFD1URYBrPqSUSOsoEFbt7Gnee7jWUDC3eEMGpAaYY482TIq
0+xmBeDpGpBzNikYQI0AI5CjsvwGvegAV42tKDJFCFu1PMrgLJuHEdFaILlAZLZz
jjoEYefrM2rGqAmOVfAfBOud0vqFv2abyJAwnrdiNcEls5fc24xMFupuDfE/wK3S
7js0DHu0flaasoa2/jjDoR0acAWog2R2nyvxZi5p4dqcsjYEvj6x35Q2iq0udFk+
eM3BBSVa4HgBEyqxVGTnCisS84RViBwKxcehTw+JVZUIyPlldnLxyNSGLO+6UWjv
i7eFpiRy42/PVf0wrRS9LdHp/PBoYSICsd0miP5LNttwMKf6YNzWzvTof2LwzXno
uWWAf9b67xUwZTU9uKibhatN5LPatWeQrrbO8bVV6CixDp4Al/9nK5QACZ4OyESB
5QAOXXChRW9JdhPfQHQ2/KDVaqBkpdYkktGpGUFnqbvnRlTQdV1dVq1E+sPo/Cny
7zMlDol9LuqmNP09cGx6q+XM7nHXA682A4/irGJ1Tso1PjSNImI+sy/bA6tRpUwK
EuPpnw46D5RKvNlbWJaDZR1VP47IShhzVgJcq3FHicUnLSimyk9jmWYGHFWXqZXk
WZaXNe96hbbAEux27ZZaT3dfM9Z7QPHh10e3LMXY8iZyEMwJHqSfjQFxn/ox6qy/
xXTJ4L+3yn+VYHvJ+kPJpg+oBDpbrRN0FM7346bmvpbTLGl+OQiTYaMivVdbb/Ur
zm2RcwKcjt3b4D+69nR0sq1TfQDsTpb/rECiEvMPyL27xgkN0sEV7JeT00RXoJRq
41QsXLbVPqezJo5J5wMLTkOvwfQfu5WODOi9lELoKV4wFBZVo3sQzGEJ/92WbVxa
88QPmRYfoZhqmnhwhyNr1nJtNPYmp5kzG9tMIetFccH0B6CNQvmGu9j+5f+wMgGJ
PAPFldUQl2U1xnDZmY8t78FWKWB/0iy3zePKO/LIONnR81/3shBQ5HLujMuWcJS+
luTxogerUVz0l3hixLjEVkps3x9SKC/iUp7Yyf/XWVjT1BmSygJaPFdP5d/3bnho
ttGFu8kysmhyzkx/YvuJC1Ew3oxtZxbxozj40+dcTAlKCPgXT8pRDpIIexjWIDCS
mQ0v4FQHLFLEvfGDs+fW47L3vpglLhln4hz/RXBnZamzkvcFykLXaAn9g+LhOglk
LN9hk90nDhykifGGryCv4pLRDvvAU8W1BOWdLQEIn+RVjrHaD5z371tbQhfgRJvu
CVmNxQMnU2Utnes24hzdfhYKWmlkPPFU7hDwgzSmBBdez8YL9NQ/pwHWlS/YEdQS
h3+7Nj2l/PgMw34SE+4vrKndgEgNh+S1NrkTHRO6psjlqDkS7+UUIIQKfBfY3hA3
fCViUwjBLHratMmhY7oRC0rhHaWKKyn48n8ALIpFVJOwgmt7bdbFpqGMs3hka3j+
2GksNgg/xh7xcQFtUACW4g+buDcSDV19b0uvGawbFAvsUqETywlc+v6T5QQW/bli
05d+OLmgGM4zTMR/cE0qW1qW75zUkBiwG8/wWxc32mdxPifyctpVAJE1f9oOD+mi
zGPjvdfXJfpf9XDoZzsh/ZxvtieOCs9Rn0369cBd42BaD6rEEKlK3Mbx9ZQ9orHz
zBaf/QEpmM1cGXYqHfXkSEnMPhA63ctwjlXDcUIV79mIDghWFWCvBDB5vSe3nueg
q7xpSt4/UYH/attap3TEVqY7gVBDcJQaE9YsM4a5EnuH/Ee38UZgsqgY7Gi2jNcb
3vILbfK3kMr7gXUX6U07rrHLrVwLA9YgNSFCF3ySozogarYMe316hGd8zMaTyAQb
Ts/FwWE5V7VLlnQ5yc2LWR1rQopWo9NGWeEGCJRUNW7vVlmAFi77Prw44Ho+IRJA
RtSw1oQTiYwy7RKSvvV2ym+IgoCtUaHd97ZM4eRSzUdVAubWPv/J62+VsEtejxpV
fE8sXWkp9/zdL8uHU2Bh0HBWASr+HP7ad16tF85MGMFNhbqPgJYjZ441DYnXiknY
cw3tSF7U91eptzRd7TF7HWYc8r2ncLEPjCOVZyMmv3Gw1W7hKgr6zNwdYzmyzGwW
mSt7r1d+sNz9bwdoBZwViIAVDU/JQSLVtZrTK57CNFS6ZfqXccTSbeDgJyxM8BTF
6hY2WMnGSTO2rTz8fJ0NcjtFCCP+GZ8jgBHkHRomn4W4eYhK26jYQpnauhfu2OK+
uLqyFzXdfhw8eMIyKoURJAZyU56j/pKS3uzPbVLQjQkg0G7bU3rY6tHu+kquFsJl
mgqMPJxj45WTB5nuWmqTrLF1Kg+PHHKy/M1tEm7iUmkY7lNaAFl/9ci0Yne8NyA5
FdOUs5kpb2P6n7hbvLHNyrjsxAG7/e/pOHqdDcBE/sW7hneHJ/jU2ujeTNBJbtNo
EOgyMv70KEfngGV+w8qFuM7NLBc/EsmuTKKXfhVo2xvt+xZaN/L4PQgu9mF6hJa6
D9iJW4uGFVy9ThuIVQsjXwdMwfAD93gbyNRda+n59nqMWBvZZ+JC71WTHGfXzjx1
BUsCvI8TAueQXqgT+7dxAwcE89NvWlI/UwaBH7NkT95XeMdV13Lz5uqgwT7ds/Q1
8BP/eEPLGJSLuhB74mX2HjhVylL6D51qTwoUx/nDfx/+BIWXd87+Pp+hu7IuGXwA
3jEgbfWIdHBvjiiE3gg2eZkVl8aizCL8riOaUm65TsVPfiNhvPJjQDzZ+o2l5lPV
C7L8qIY9x1Ei1hpkBvDMOeB1c4M+uv4KXuKFWbFmDHIuprIxtwjlj+4tjOA1KQme
RdM3uiuVtLyIardH9MbDVRj/2UAZSIpg6vWxO7UoKJ5egkxUQi0i65xuSlVKHEVx
UIVRXGehadiQDCXF+aGZOyGDU4J+DRNEaTxFYtLetVUEY/ARAEQj+j09IXX9kQLf
uRT+WR2yGTcl+o8O/REnRZN4CFp2OnL86om0MmZNUdcq8a2ns3pJ2P++wQNc3JQ1
7/vufV/KitStBY4nmkB5NuqvKBG4FRF0KiJ4UO7RAmLsWId2zLMYqpnD/xw7F+59
DyJnmro897bODrG6zsooNGu7ljLM/0CeZkHd+hO2GtUh96BgLZ/ffPsFHMz0DOhq
2n834vw/n/hhnn5WrWP6zk44ASCN1DHo0/NJubmwnJEC2mCaVpo9oZVqrOHQnwng
MsPDRj/vbcCmYPnX+z+fYsrzetiBl1AWr03Pzy/gD6CcBzJNJ/RyArf4158XFJnd
i7QhiFAoAoPg02lrpNQ3pCNI4tmPnQXim3PXCCqPuwGonl7ngkTTf2mK7ql2GG8u
3nVykPY4b3HRDBBDOeEH66Z1Sr8GLHzgd2e51dn+5g95mj8qKHLXiNnjXYrQLEhT
tUuy0EOQ50eQR12pcZ7/P2Aq0Q/Ggf051xMHv8pcrbobMPBhhxAUkq0LP3zNDZfi
Fsc5XH7pRQuHVqs5SE6TiyI7wM78FpNFpABaNUa4PoXfY4A7qf+0hYpa+pgZshlS
KECufkU9E8uz3FI5Dgzsr/9u3mvfrmksjqEZNcRgH5meIZwVxib/ZninjzfLEFja
Lq6JvdIxnlNmv0Bwl+8808Yi1mMJ3WrYCF/11yuTFy/I8fMBbDIovHUSxc7BXSpR
SoSTP6cpHh4XAKstAQansBOYRnJguO7hjWdniEFc5dhihsM5pP/FGEJa34EXpMPK
UV30+q66qAMYv+Y4tYXRuqOWRPyZ7TPOSK3uxcJMeospqnxkdEdzJU/6sSI43RaG
TKaZciF62lEOUQlZtQT/KP8NWM5l2DX5YyGL2hjCt2Oy4mswVChDaEOIp1t7+OfU
UtWoZ5T60iS2C26+JSwAFZ1KV0Y+u78r4ozsyDVvLJRmc+hNcQBawcjpSOZ+G3JQ
Ely8/HjSj7HF+JBMLoT9xNICred3qsGwS7P5xEt7Zu/Xs0RvBhL3hhvxTApNv30N
j0EE9AITozDHx+1LsrAXvuKYawra+sfD+MKaW3Dk4gV7S0DbOPFhKchf1Sx0ddkV
YYcjWCcC+DLNSTr3aq+TU2/Rh94cCahDczonoedH+pygZimQjFVB+Awqs5goC+Z6
7zliFxzF6YnOzc9SuJk8yKf2LtGVPNOCTFljOVhjBltCDbE31bmSe2XXX0zfv593
3ThlP6X1s7fVKRcbTQ8q4QG2qqLaT+lR7BPaNhuTEtPAqftR/89SYjKYV/z3M0td
Rf659aRM24Kp41owXLf3ECslxCA592Pzzbmouoh6boYK8pfm1l8AJhknTBz1tjsp
dU2hTNZ+rdACMy2iV4hU3lEFXGWsbbmCOQRQI0VaJYSpT/McsJLpnlrPomM6Hl86
1Blv+Qo2UxDPbI7Wz8hkxDVjn+DQo7qh2kyLS+uNKOB58AMM9RnxHkpon2885LAz
R7vDga5zkQnW8bOIrTpyC1mkF2SvAfwMP+gyVV6M6q8OZ0W5EnzRCRh8Rlo/ipmH
noYL1IKksNJQRuO9fdJp5Brp5EUgfBu+3WAwgURaoLgYODau6Kin7DnurScJ+IRn
52HibEAXYgThD9x2to9y37zgq4NkO6tptxJ+jngkDXVBBeNXHQWevJNmYPAv5mbx
e3k3ai3ZaCW9Jcolucoq6/6UMgToma0xVlLzRn0oLkdgoy6RQgher34Wewiycxmh
mO8ZdC9+tqWK8sqP9fGqGhJaecJ/rW7LgaXNNxrBpNu1EwNIC2ZaH1bvgdOQVIm+
vQR0yiLiSJCfl1pZr7fBgT3H+6fqQ3l+55H2x0k8/aa5bjzfaaWd0l3W9FG6gQgP
LweSOqYhE2K23Erm0nTKaP4L/2UMj3cbEOcuR/c6TWuzzPRN/dtou3FeUGBNIrvs
0M8H2pzC7KElOAAJMzKpRHCMsdovPKu7L46p98Mei0Qt9tg24TpXUcNcplHI9H6y
2ADhFMBKgzhcJBMkHSBjt6/jsV1HkyM0GDXl0AzBo8wwGZS0YGri8ig/J/wlmio3
ELsGH022lM8TdP2SEL2M0S+3pyPjwTjhF0RKE2e8+ynip3i1GvlCTV412xpsTwki
rPFU8CHs5UPailR24Lh4Z8f6dnQ2pYNva3HVXqY8VkW5NjDRSdp5yxoJ8LDsROlJ
yVGjQNvTwJoFMDEaiXV0RSzD/J/UVIMiG2f84h3qDpmNRsRiCKULjIwky09MffHJ
g21l+WSUjd30VWly9DdgDtaqomAwGsC02giB44Hz6QSTNgovT1wxz69ojz2oSpY7
FN1CLtYphapoqLyZNr3JjzA/a7YjTOX5PFlUYByxwlD49Z5lnxkXupF+pV4p1rIZ
/gYb95VuY5CZvZZhHGH0xe+7jRBOvSW2wM6MhJzZ3tq5NZCS4imsbqMptHf5JvqC
yDlKzULESfNcrStl1s1dJ6DoSHd/6/I1Ax0mh7aLTWbvHFjsriWnet1S7lhbWlfm
bYjvI0aAcpE084EfjuZS6EG8fWF9UeDww6xtJ5sm0lOTxamRLPZJukptKwhkJHKF
FLyv3i3zthZftUUUIQNpAwH16VTgF48qnFwMG5m+cWEbqRU5W7D/1L5iFvy6A1nm
u/LrCgZMEH7N5t5aDZ7lShIPKS2mDjvhdOYc2dWA/JaHXY6zu+eaz/hEbVddBntn
B36tJpEUBdesj7G9nBSZsODNeTNCS9h/RD6iuzou+LT+au/aLHuDil5+2TmkCFbx
41bgFedxScytSX/OxjeyBROc4kt72nIFEqOW1HSvBdKfZxMTOxgoZAiooFAbOipG
5QgKJSX/aJAMBr8OrOqwQ1OENwBwHGIKlEIzVmSia1qveI27qB+TwCVpGb+tXuzR
l2GJWuu8wOz5C9WaNnZCLVu2F5rImOh3dCSuVct07YifcCPrUxw0q3by7ApoWg93
SMnpDow/xSa8E4Gh1CnNzUMtu5JHHtKOceWX4Jld/1vyLTRtShAuiwDD1Lg+GQ6S
GYh37HWFLHLKfuwDdZt0zSpsLetxcCVQwQ2FVGchYGVqYnHFx0UGe4IBgVuJUYwI
rjSpiM8YNJkQdhHWNWQSXchVb6wtHvHoJAmB5UL4PfsNrDWRlzmeFj9OPMGj2zaU
RWxsVdmO53ERCUEP4HqWKJdHn6xkI6nWgiVTOoguJ0G8EXXLoLGMUtW1R2ztprcn
y326iXMx1I2tQfRHcY+uxHTW2lhsF+W6SVndACju5o50rDyy0CHaHxXLrofslfUu
xdIycgrvU23ca5IoeblyXya6uMYERp5T5UDh4HoyWPPpSyhCTAiixUakwYoFZHxn
e/vFBjayo9hYwyJ4Ohm1mw3aFow8FATNC/dM8lgoki5gIS4ldXltH2ZN3Xx4+fb5
WkSlFTA8b7/OwHbnL/8dfBzgRygTMrTtPM3WUNKDzNXOsXTsMZuybstWr3cZO3pN
ZHvObvjbl0kHyR4yJ6cVwUG1PYcMaERbeOjsxSVBdbPGiRcgUFmB9NwryhOdfwAf
jJZWx+M1FanK8R7koExEB2NzHdsQ737T/bEnVyBkOJcjvLg54ZfRUID7dKu2tGzz
OmNg3CQYYl/QQ67zPL8ghRYpDhgA9VDYZmBqPW0Wr7O00MD1EV7bPGxzvmT8lzIV
T0l+VqfN4jBBqZBZmhpGDCh9svGdhA46+4zYdpqynAfvvRSvBmjdiQhtArcjTS8p
b3Ws+8IORcvnvVtnLOiySxNR0p7z9yvd93kr7ZXY54oDJrv1CkRpVg9Ejwuw1RTX
zoxO/XbQpIcOF6ytPVTFPfh6Un/wAv+EREOcQKcRHYnFH3rI97k1TCVYIQnBeL48
e6Fmpc0PPl0zgRQphTYyFbhG1rdsGRDLmgChPmzKLFQqa43HqC0xweN6lpHzg0ss
C2JrMj4kf9ty3/NuFZ8M4S4YssACPVnS/oZpyLlXS4qkcNSq5elvMLObuxZPGMlG
hwmRA7pagaCDe+chgbUHl6vI0FklySywUbMNitMddwZdKlFqZEeuCs2xrAXIkGVM
QzvNCcPMWnEaiOsKfibmOanYK8FpdkHUfRjZDiHMTRfAJyPm2ZVGNnYzS9sibYNM
erqhXTJ/HKik/6szugt2cIJ1r7lvg1wPyIz/XtoQNGs9fdCXay36V3jZo4velOQZ
iONLqkuWbv91oKSefELPUDApPRov2ZXngNqAEHTLu25XbA7XlUlcooElhmtIiMBV
xfJII5b0S53Zvk+v6/1Blioitxmsg25OU55SVYDWxYLwBlwvzTCV/VfqNLEiXu1d
E47zwGcxn4IgOQO9kySbDOKMzFW+yFmag16H0LMBTFEK5yTm88hmXxzRyP77TK/G
/Zr33Ye7APlwF1sv/gQ4nXaeYjGhqtITkqX67/slUeEjsVf0DiRo4uDNYVwERHL+
Eonjr9ytC8q1ZWMVFTe2F6nKjOarfJEkWlUbGwmUUTk8y+f4d8R/wooO3WomNp8g
/qFlcD764ongaG5L7nNT0IR8DeqLgdCEt/ks5jYGu8FREmASTME8bpvUeyQd1WUc
W/g+TztIm/nJ6kxms3qRh3r0M8aslTn2wziOPzHuK47ITP4BWRkWF3WurGIpowIx
pogO7xd4cuwzAOpnfkoZIPW200o3X1cm5Arf7U9JJq7lIK7YJH0rPDb81GFUvj7/
FDKuGE1IZISsX0djFpEaeThAEkTtdP65bZzLlBp9OFmdLix8/znO17wPvkrNFB7F
V9YoN44L+4HKU9jsDtMHPfyxuVOO/WXdfVOMTSjjZCCyJ75EFFykqxToJ/bg4khL
HqauzT0YeRf2j172z/00O5raDzZfCDktyV4izyBZUNF+VV8aSYfxbxm49KrK9bsw
YaKefHbuuvq4IPcAtS70AGVkqPG7VeB/1raxPeYmqUa9Qtqk1JYbwo3Yc5HYS+fA
AgaJNM22hmoldrm6aVEznSLzGK2HXZ6wWfZNRUN0mw+b64SPgmXo13rISBrHggKl
ESBaAweK7iD4M/VqMWeOYj70dUt4SvBPQVUhqT0AUcDIpZFN6gDIp2mHQaQkr5+q
TF7Z8VAbspIJGbJHkBr41HFquBr5t7J/Pe0lSuzBccOcEZRsgUfqbfX8KVHzmCU7
aD5B+Uvz4cdnDFvhp7Dihhi0LLAd4Mg+GF+soxuotqkxLQkudSv6LNwEM3vTbub1
dyfJ8Vlpcrrr+usXH7harAwtUGZESkZho1lICWbo0HA/HN8nA7Fg1sELl6MT2ceW
FvtVxZCM5BHykzRypVaqhxxQws/gc4Arjx9b/RNNb2kjughjo+KLatpXuREWZ/fq
MtBmq6eNlYeCINfQNAis+VuxO6MdNNj4eFS8l5YdzkVf0CtnujmlLFbSzPUxaAVT
2rSqnzpJbOIoPY9OLP/OI/PxdG+vxmCtCzL3joT6TIztBsgLIkBXoDH0VlJhFsDN
Wj36vUXk6TILt+tYx8PThtSpSWK2qUtGlYgCQ1BkMPn83z0U/g7TXWbDYqfiMwoo
f9EyLga9gnjetO2+KqZYV4jrqRZW1EjM/Ams4TLx/lHUuSXjncGETPKFptnxF8py
E0A9iRdir5XeCqLPEBjZl5oTzzQ5Qbmwn9FWPhwSnk31o39ts/RKxCXLNoX57TFF
0mz29fZZuu/ECmUS6MfF1wpcDgQS0U9lg0zgFFcFs1uQ81ZrVpk2eHChIwW82f9b
BkTm1nC7s8RBAmVqyALDczwszsK/h1bFeoJ/HNkeF2g0sM6N3oJYr1dayOc6fAui
dmuuIXMYAzbSejiTP/lKJS2oMFe1sKyAHCEQriP01mqiPECo+tWHRDdfPxpmlkSx
ur1Uke/OQiaa/B4H4OV0MaRN8VNUn1+n5qjOWWYSPbXWHPPeYTyjBolVGFyo1qU2
HeWDo5SZtk059/MNKv32PKzPmKtMK5kOOMhXIzRbCq5mLYtyMP/nbTz5ygRsjXhZ
9osDy93K1SRinsqgJeyypwcSW6nid3RWUFpvWvNhG1IOGx1sAEJREPCQFbpOdm+X
GIGtXLSvD3lK0TNvZhg3KuU4b22w6tCsflT7vLmLsgPpWi/wuU9p+m5SjeLXSrTZ
SCrTj/BctjjjC4dGIP2Ml0lGg8viXmQRtyweKmsVs5mgpE80gpoi9ofbnMAh93P4
TUc1A9q67abpWfMHOMG/gOqjkDVW5p0Dq7kGHyV1uWXBu/yafe6elY0z5UTpP2SU
bUSPWCOb6P0NSm3gstKf9RLchtw9B9dFsldwTVADLLMbNgH9J4w6ukaNs8XjQF4+
t9Av95+NSTL4yolaCw/2AJsvcRv4PA1PvNO5hxqXInmXVAa6GXbMEBcV7YXFV8A7
swf0J2CfmtoB/5xMXBZXHjTwEhJovSSrp/p4vlFd+MrDEYQ+G5KAbBWs1uJFlZjW
o8DWftWSBtremZ+w41WYEZ6gMZW7200/h4Ob2GkxKn0jzGVZZecxaEfvyaLtl7Mu
Xm0Y/QCXZZCNiKbqqjM6t3BUAnAt9i0lAp5ro6wd3sYEEFzWtviX2qlwN372Zxai
IevcXkLNGCqm6BKgM3/30uZ1F0tiTpyybuZvOs5gNX2M58rC/BDIHpQA0rm9rvEU
AB8EumQBbrxwnTuqeBPf01DWeKqVDSFG4lyGggxuLmQXLTxZszh+l/eg8BUvHoBT
Ml3us2HTGAW2jsRkElbQXmakgXnGYGuBS6Wph+AeAiHWKZMPKx6LoiuwwcqQTkYc
e09/RX0fZ75H0zA4oMnO0oBwgRAPwNuXW1ZfgQXkSMnd7/zNMP9vy65zinaZ7/6F
OJLXfpkcG5OxtyE9Kx0jjEK4RQIEg8Zmyjel489gKoaYgs9fK/pu419Es2EbPRTn
tVKKETBOAizi6/DDejPERC2ZvKbsBpFl6pVfj3j9bEVLcKpeYkFAp3N4TtK+jK+u
NJgZfsTYFCe0a+sEegE4L/YtvGVf8E/Hm3/fJmHj1T7IUHi8I7ANCXcpBlPlRIaz
JS5E3S5AEJsEhJb2BPxTvj3IM1kZ2WhUgq13Wn6fTck3ziHf98lDV3L+iW8d7ggB
t1/qEA4gwu+X/QdO0U4u9RaCUoKiM+gMQzFnAiJ6rVtE3fXzY3m/+8q2oH9tnYgO
B+YGF/n+Tad4bbDoz3snZg0P+bTnXVL+3xKPTUHFHMWP7IPNyeR2FMm+SUYeqgns
uuJZvPBFsEsvh2Ek0wgHEze1CegxrwFQe4xoczVHjKt/SU5c77xE0qXWVa2wUrE4
de4iLaz3/8+ZBDhjA2qURdNprjdmEtfOAKQ3Ud/43aG0c5XjVbptXbixxjrgV18T
Fa/yR8zrdDaNea8IlkBU25wotxGCJq7CnWMYui1F89GyIb7zZ8CCrTQ6Y6BV8Pi+
FAF4oArXIFxbL6URVhGPqxjBT/zQbKjYVfhNgE/WmtrZVpvNajTfJUmZltUweO9k
v+AlsnepryzIBt18QKiZ/ham5eUFB9UcGQu8PqgP8EkKt+esL28eoe/SwEQfMi1E
X7S/7QTnbCYUJJiiMtASgnZNxVRBcyUUSPdxiEuwnLNlLCELXK3FI+mT3vdns6HA
O39vQLnqdsrRkdCn02uJA3l179hUhMxXBi+HvezWKxYuzaWZJwy6feWqx6rjjFZs
xv+E8vq54ibuFcQoZ+7IVJHouaoomaG3usr0ySCSoFW6lWhunDUEo2LAij2hQptn
DFmk6oW2Skn501Kea3A9x6Lwy9fNtKgrge7otxJLXwRLcaEo7cxUMoG2Qtajp140
5KtvzI62wNozBQkZmhWL4jEZADOeXPSZgIbIUsFVe9ZbB1v4lG7bY+2gVc3gV+Pi
BqabKKYuwlXmLF+fFZazjjuBaYGX83yPdsLjfcYCEEMGZJpjJbCad96enU6SylnQ
PpTGsuiBjR+EWD8MjLkGCYl2AVH7mqS4swQlNn4ee/73O7lVkOw2keIMXDKozeLP
hAtsVQC2b2DUkW+3Imi89tRkzL2jcaAzQ9pFAdiPmg3juaVP9YTP/ZWU19vESrZH
tc0Sy76H9t3bQ3mKjyc0LY/GfEicmt6bIQJK/py5mJ2NRl7t1mxj03MobutV4Zt4
cAHeB12wXi4SAgGwt2K3+Igq+/hZm3sgSjtN5PEdQUt1dFeq2QhP+U/T/IlE9WJZ
TOa+OZDXEGmc9dd3a4AF2xD4t72d364s5wcm2o2Gy/MnSstVbawq+NfGRV6V5qWi
qQS/giP2cJ//9KsDKqEc36R9z6kZe1Y2GkVCm/Dt7Cv4i3Lx8KE38WB9NsC0gc2F
RWyrholuj/xIwlH5l+R+MuunkNf+gvXKFEpfeH10hkeREj9OL4YLP9mtH/PXXCjs
9L1B2giijKUALFrFXo9mtuDVOjqGqRvX4UC3/oBMch1w3HhWzug1P5RU2F30dN8C
+lQu0zrP8VtxQkek6FwbdsIbW9iZYGBXl7qJ/E9y5i7+GFNmF2STDyiqoRCnwsgV
jCarAAEoabjDonLvxhLOgvp8tHaGNUAOb6GjrH8o95DfzfHti9x4Q/IAq4LyRafz
PsYzy03yWkwvXwjLze4N4MNZLHjQtCza4HLyD6uqkIp/3MREiIzSKb8Xcr0uHMUk
3ZGYkScQLiL5+1ho2KxfeN0dOPOKGcoGcEHKXlnlgBJILn5uZ9qpbGpE2+YKhtv7
qV/tFnR0bT7zE1NtMvbHGcqwe6vNgXxVwX82o79/e96qXI1X4mn5PDLx7k/dUObR
u5rJvN6Bfwz5E6ndsU4Oj/t4iEZZKTIVmA2PF2IHnyrY2N3LK9wA4FtKKp+PVgNs
QXrb5V6KLDvrtTkVlZmcNG/0hmuWU9993hY2Zyy1H0tzDeEL6VLPJwjCr8dn3jwc
OmFKIEXC8pF1SS9bd6rGhnm94STlvYaAEtv9mhaS0g+hZTtqtAZ6bZOJ/LDuabbv
GNG34J/vQTEsPlAeUTQpTdLe/moBU8UTtl+qKX0dt6/XUROPD6SgrmoktiHA7rQQ
iudXgQaF91IlxJqQF+i5upy33b6wbQY7UNqMVl9hucHGcXmteo7PDY2Py7wsr+Tf
Vsu1DRH7yIKSvwEzGwsJFmuhnyXUViXJetZnmnQgIGhu5egPTGuJ7TdlgQBxzgsK
W9ntDIorpQTjTotV8HzW+msTDNTs4Rb0gG24eTXj838rj/WoFbAuDmvkRXzHNsHu
d0+3xst+DO/uF+oyta1CozYAhu7I8nQ8yyh+e1JA4qoBOiNCFIfuDjGRrVBJh9KU
ojGQYAESpa6P8OsixRfkI5dFP/lUR0XIJei7xuqrmD25e3cU6cGucZSmqYqzBAkt
zoGw9gXew7tbfC1GVr6AD4LjmZYs96aiNm2+ZZ/XTUAg8o8jXCJmhZp6/Ec+kdwi
n8skI9afjC5jWOGC1Jx1SOHk/KjHDpZERYwAPzNvILqgce0PBSbrUOB/syeF1r1X
0bBHg1YRqa4/KSEjeXqGZzOLJk9ui4UcAvFPujLClk+oKL/1Tu7UtJZXQjUQFTzC
p+fZGVldtNnqZ7mTj2L0yz+8GoAmQj+n3x1/HGGQHQueXPDFazfoawXJuXEQbQ9X
dFWJFEa2njCo1bkxrZBB8qnV9+mAqyDuehK2hcEbY46l3UG3Z4bT0IkSUy5lH8bJ
hkf62zIBXUpOPOzLAyA1DPZW9k6fsSfCzWg0r/PrtEpCGUqOh1jNlTUwx9Qoo80K
U/yf7ulNpOX2aB1XXnH1wAr2ZBBSuv9VSHIZDEPfv5AHtK1YRov9qTT+vIJ2vk9j
brzZWeWUFDSZ/Jy4WIhSfZkBwcwMcGxlTmsxU6tLE31d/CTmxbEgTDJaxN0VAOT1
kDjR5NpNaviDTt3OBfVhrDMjQ+ObhcWwBqVXpnWh+tgL6O+/Xs6XZDZ1jjF6RDbU
0m9oufZh9NreJffVrY4ijhGOJD6LepwcnYH6jQ42VwbSn/5TEUgN4eyoZzi9Uy04
0nK7dtSS27Ha/noskLxRTQKoqu/cfcjhFZ5xFbYZCPkWJDr+dnj/GuFw5uzi2M9i
HdaUMLSSEV4pR5W9G78MGBZAwDf3GeRwtmuETteNUphUHgwSXJusdHYjbaAOm7g8
X8vfK8RmzOndlGkMFdGYnG79zdunFlk1KqJPlnaiFQqzLWfORR/ye5Da5M77Cbfw
m1+SWpA8ntEJEDJP7wphs8K8rsbk7tu1UFvXiZHxGY8GzovXFNWxycGuDDWorX4I
H9vsYf/Gfpei7LwtzyIEpBPjGA56dyfN1wmP0usif17Yzoar4kau/vKDZOoIjMgY
4K8nHtEoXnCfJMapw5LSNxf3aMWRvXdmQfhJKAkHzqlK/NNYB9PqFL8EWDFspGeP
yH2yO3tFoLxDSuiMluxcUW1AcRgXQitTN1SXeZhNfw1lF+Bq9UWJV53mjl4Bwmwx
zKQTfzEOo4NsKyEobxv017Fzz6yXMxNjytA9GdxhXPeG3XkygFw2R8NgR/XYHF7k
RvNSbIB+q2+KhSHlhIGaEE3ke6LwIXa66uUjSwc/LHtHVRtKh1egbnWMbnKGWQAZ
NM25rwVwALlApT1VkEM2ESIxrcrFp7OzEgJDRtApjGXFExN/FWr6kURKC8MWS93A
Z8J/KEDpT1FiNPOUS61zyM9maodKFx/ygzjTJSQirbG4McecjQwMOe0FlSEvkIt0
v+oZIk8uO+6UsslYOa1L0VyvdKTMNKUkMIS5w8+NMJ8QnqvFMgUJFC6sNdD+1B94
enLeGq1Y3NDp8muablzGfvKP+RCo7dCgk9C0Hm0fezg2FYTQYj8JT2eINIHgEMAw
HkPVTk/Ck9d9imfBHSXdMwm7W8XQIhZKDozrMjE2ShgICNQLAW8t+Ber27A5zwRG
ALml/LUWwC8c0Pqmf8mYnxSf5M/S/sxEiiAEqdQolHRQCltvlxnlNoiEWG7RuzQQ
ow9ZmmveWxUeoqMgOeYoembXyyoHzLuxDYSRTB6TTa6aqK4ejXqci6vGTNTGnu0y
KLDn2nXS4LdOquXX8w0xYnlMGjNfozYgy9Av2AZ2BS+f4xoM+gWU4c3IOLp8+x5P
eqp/GlK5wBFmxDjfOK36E2/hLcJ3iMg3PGGNUFp0ZLM2PVxx85RkEZIITJhAJnPa
/KhCNqTTsD5rK8cLyQa9sQX+3K17YYhBx1Dv/hsjdzO1imLvNymxIhy+5iNptgqF
xFeu3tX+jH6vpmpb6Y93LG8R8deyN7PaNqFLdp3f4jQVJ5B6wBWcMWAyK3MMdhTm
T7Oiotk218DTN8m0wewRAeMnWr8t5+vP3C41ZFMlry+zAGGvwonovW9RNG0usaoY
Hh6PxdUger0i2taRWSt7MHeP9Y+fvHtr01B9wjOpXUr/zBKcFbs0g4mhSyzfHSaa
EziQ/SvlR+3nWjX4OiTyYgvsp9S3Kt/YVA+titoQzb7wsvxprljZr/bWbXpFiVG1
9FFCjiczFBx5yEZ95DmCoZBN7eXY3hP/oYq009fBE7E42aGv8KLKW8PfoSnnDRC9
DZwpXdVR8kWjXi4i4RFiZ6RJ8YSRSLnNrtqbHULIKW+sjBXy6Ltxue4vbS8UgSes
MMHlaKDcrGvHSsJyEvv4KZTUVvLONwrxs616SEqbQ65oJRvHiUEX3AMqD4VU9V57
kShEbDroF2Yvdj8z7SMPkfoKPZte4Q18pvdNiCkFPXewUFwA1Ds02iylUqsYz5II
Al1ldMjfOgWBhjtdLaz9m8beQuO/kbW2ZB9EEMwa/MQ+4gj0VV/kb0totxUMxod/
yAtsWyuyYbkUgCuX4ljN6NfucEVkxM+3m2xEGXZPrVNu0spo+lbbv1N/rDWiuSEt
Jkb1fi5g6Db+hYMEVc3J6/5GxRVhxKGTKg6x4U+AqXmzzhp608s8qjA34d63QTKk
RrsHzVXhnFNPHzo3aCINDfFlTmT0FjfXud1LSEb3eqq+iLZ7wmCpN+bPOu8gKXpw
n1HL5e/vnSzQOeq9QH9AmYZkUDIBDyvPlEb/2Tiz9XXqv+W0mp6Vo/oWtw3R8/mX
mEf/M9v5r3iP56a3avBlnaxjoNqeFukfocAXU8uSMN4lGIqtjkV3D6c26/YxgrV4
1aUaT1IcyKnV/41U1bP/OC8sl36ETuNqNALeNqCpEBxa6v84HPDLgJLBmWjW93az
w83JO9vH5C/88KjFBaP5ezHzn4FJlVH7oS8fGIzcJkOFjM2ccAcC9SQ7b94H93Tz
GLPHkRgKg1R8c8XHWmVDmPLohq8J7fceVywcjjKetWiVL+m3yO8QZsGA1CVs2ftb
JvvgN0SxBn3nprLZE1sCcrz02yn1qkBxcIhny4DnauYJcJEZQupDvfGjuJtHRpGB
V3cXuE7DlHjXsVRI75/loII1piEIYngRakp8K3TK2qdUjDIG3ITZMT7gACdykF4O
qnBZTWcQuCtR0ppSqMrY+hNKpYiagcnHrY9IZpUMcQL0HEMyF1zcVaA5ba3HxGTA
3ljuTvkmd5pun/DirYrFM3UIskPvWPiMZP10crnRiiiJybv/oVi9GtW/Z1W57Liz
k03Un8BfGy19ln81aA7s9oA8UeCrA7l1DPJ2KG3OAUHlMIzSzpUgWipzM3qNfLdt
9HaxmMrpORMhBeahVABTDIatPP+eC0PLny9zNqArkvXXM58wBJ2R6p6dktEf/cgJ
OZaYUCbUvCC4IwCtzJ5ouemRg+HrK1VZQAZCr+oijVsa8Eq/su/v+Ol1QqUz2P+a
NiqRUSAOWi89BZtfqp0fkovt3L169doSGltCdN8heYV8iHeQWkNfg/guBUvbRjbW
LbUw7ee4fcl1iG3ctMw8LN449gCdTOtljTyKFh7pQKjVD0Fu6n8322KcXozgu1ut
jSWy2o7N5EToelEZfVZP6nAI/fKlevxpQr40v/L9PhpKqDaRZzGAFR2OzFTFWuQV
j6pjWsPVpF9kiMOKqqDMgPTUIPZL2/rqQmRYZv40JBZqu3Ivim+Ho3Oq6QxWpVbo
CoirNq91MRjxav9G9QfHd8iMDey0+8GAVI9OfSWQq4jDXJfhV/vfl43cYh7wrIbq
7/ViEBLii0r2NhoB6N/K63/Vwp2/hLHtAnN1699xGxk0gFl5B3H6DB2AKw2PCIzQ
2sSxwrkC56z1HWdoWIgmF6B1HUk7CNY31Pur5UdooeX0U6tCMy/wSBrVMz6gI7mk
cWHGbH7c9tIU2HdKW7DvjTRsvGRPDERBg9xpnhY3laI7jf/y2xTZr836qig9TvFn
kwqKuTDN9bauVOjcP8fmSawuwFDpAIDgA+D4c0DHxD6ss6GQ00qPdmn9QJvFgnUo
7i86HbRGl+Q0Xi0uP6FXU0kX/DlBxb9sEbvWxpdXAxo3S0ThXXd8UmjqzzXWsuoE
oF703mzgO40yuCCyHCIcETCKw8LvhCjpeEaTVdgBm5RVJ1EIjh5xVY+n7e/ecmer
mi2hfOefzf1Z/1j73DDIWxAU5Hs7SEPJ9xnQ9X4+/IPcmFzqQCPZ6TtODdnw5moT
LitVk9bFTZWFKKMs0HDLfna3i38GAcQELi/xLokiCuA2/YHPwmKGebGju2Ulqa4L
L4Be//lEq0N0Rm2yVckwimFHZSzF2Uau1yOn0HcX7K1U70z0iAtar3MYgwmOkaXK
vDdRJrj82+HmKpHwGkISiCrG7HtaZ06eW1pfrVePaoJtkBOyfmu5oUdEjFfoV/Ed
8NRxNSQhA6jkzRFv0vPdK4j54Nse8OatRKdYk7T7TVzLCR+PbGwbcja4Rig+vksP
9RD6mVMMSEZ7O5L4+CXWkXVRLfGXnxsku5f1PCI936biWYWedxvVKNq1lh7EA7bp
TYz8WtVho7HV3k8hzfsxkXw2kEyMYDpLselMotQTtkGO/Plkb6Nfx/We3rnZ41ro
BqVx95HuqjXes6qfHiTkz5/ELO540KjqrUgjvrykDBlRib6MkTdmNGtM/dq/IGfy
bVQu5Vwonq27eHUzmloAsvx0Z3dsnSrkKl/53C7yFYrEYeymscgl1mLsKVjRG620
v2Z1Ldm9bPy7VJD99SQYV6YzcCCvCBlhfNpO1hXdqqa8cVrOUjQ95RroFxhOTrZ2
L83eFEOfFLKqgIY7Bj5nPR46Htd3NimcAeZ6NWd8FP3Ie716rGpeHOVTNVqJMsTI
Kzi20/9nlXOr1CY079viaKM3hdbaa5ZrnLBDvdD3RgJAeOHuYw6HFvIK9h+rIPHj
ixWL6lNdhgFtjcUdOtacT9JP6l+npO8HUfEKouCCRxYjfzrfyppaj5RtsGz3HJHb
teManMEi9fTNFprKX3x147NYUE45nklhRDPG3FLS8fyulTnnPAH8Pdgr/kWt+v86
tk1RUi8cAFx/CZU6zvAIFTEDZisM038ZUjzonUB3Wtr+QEFgYRimMuezGATB5ynq
zTmUhD6Np+i/9XNEsS9yahuBMYTRElV5El6f6N1hpjAUjZULtCrFAaKaLtrNXWVx
ZvV8WAtA0CrgszOAF2gD9zGPj6iRd780mp28cQFAfLXjxO52etZrrHc4EXq7XDN4
UlfcOj4fx16uTxKl5hzixQ6/XGF57830fpOXPTPHf1lQJLoIOhDT/tbZ7C/PKlwz
P5iDIHGoExN5SdnuNQVcydWTSEcOK1DKipZppUfB1DD72byc+BprPyF+kDb9Bezo
OWDb9y88xC7LTgeo+U5Cb86yzaWU5658iyGwBpmu7Mf2EXrknmEslFT/9L9+xx3P
JPsBJCrQB86FyGl98BRnmamZOaxiXiw7a7YuaPtrsMqqZa6J8Way7QVll3EtKSS2
llHiVhjblivLIAoN3QJqU5es/SEa9PWyf+EHKZOavB5i4WCZmSLfIhNAD3ifQ1Xg
yT21hFUCz8bMfAEOMOaiSa9qHNVcArEgm0Xsd+a34Zsmcg7VCVuNd54ZRamn93dg
MzIz1uysKQ/6fMpq5UI9JKRBaIgsFaJneIvwuQ+yEolOG8McL+Rc0d6JRgANOI0D
do7OY4NkkZ6M5CNrUyTmc3Q8BmDj6TDVV1qg4BG71WkD4ZszDERPS9oqhKARJcYT
JT8QY2GhIfq7Vp2z7S8stWcOQBrLkHOvZl2Qdwo9ZLBBV6m9+8/l5C4Rfdg+roDM
wFDVIsck2P/s1XBugRKOON0eV4/1Zc3j5c6HsuuDcB4MT0HSs8xS95bCk09dlBSR
X8fDo+IwuM9ful47yWT18Grk/cp++vYbrhEJDZEpuTNwcQGWZObNQioV8zkF2+PY
Kfz5AUNmcKbo1/4n0Wk7s1s+vU9VSC0dwQOG53oW0V3WPzfB7c7BQcBCCYTAc8E8
qdZCM1PYsvRe9FTRf8UvNqtp470ywDdvb20wHeKFQaNL//5m5Z9pEd6HxZKLwFIL
1OqgbAJjzXFlbkhobDb+kH4TRYr5TiQF5OKKxqMrdLflJfYgWDrmb5bRqaz1cONO
pNUMIqGDCMfRdgIx+IX6mnU48JMe424CLc2eQLMlUIiqJC60q1TiBaCFukRNtM0H
AbNJa0bgdDpfTe+R2lorzdXPlP2+zoCWVK+X+oP0KU4h4XOemObpdXlxrAcfUMu9
+xu7bbWQW99gnO9GnvDWoyD2Pd5TsOAld4WKkP4IekWK24u3x6nfUBD8lTyn4r+U
+UEcit/WGcq0jDRUkrsNCmxH62Y7ZZaRrZariv5aX403nO3fd5BPHbpc6bqx0ORI
CEJk7iJYMIlpiDKUbtdF8NDL7JNBi6mT0v3QRcxBQnhgx/qDfC8setRUXtF63Yul
wQ96VZ+9aWws4iFPDlNpzgViPBXRSUrJa0Y6+EktCSxuUBNyGWebmxTjqOYqUKpc
CI8u9kA6YdHpjH3HkPYyxWNCOYkDbO+la0MSv2K1UcdFOKfJEH1KjH+G4K8KN/rT
vlm2gqEaLaes+LUOOUWBxilqC9/sp9MSIQvWAL7t3FxnP/uFjwtd+WltDd8Mlkdq
v9WOwXNwinM/IMqXCAHsoV58j1S3mc2aT+Io+Cl96bamvySRK6Otp4HbyTTEluLg
zqhzwZjGBqyCCVQ7VJvdjWOFlnY2CoUBrznCexV5Ii6w2tbcQMOaCLcoko1+w2s+
z7C+4OVAv73qLRhU8qLy2Q==
`pragma protect end_protected
