// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
B0hFEozGHoC7/XNmNe9asND4gznntShav5Zqyi0K1bc8EgUUluzMNMTltQIXdyu7
qcb6b+5lc+2uYP2gxW4Zhh4RrY0jVwEYE1aT0+TlxknAMIsscot/U7YCLjG8yKrc
runSJ63Lg3/9NjwgTGiled4wh4yvqS0mBv8sqRSkBDYOjCfMKv1gIg==
//pragma protect end_key_block
//pragma protect digest_block
sBH9m53FCv2Wf8mQRF7kKWYCIQE=
//pragma protect end_digest_block
//pragma protect data_block
bWo5GP7qtUGE+rybiwBb1Fv1iFqj3LJZRJFK4HllFVyOPnhLZiVg7neBpCq8nuWG
ID0mnKdHWpLH+WeMY5mYu0UbWt92qzjk9drRiB/9gY+xil44fpgu7PxBYDyaEMJb
Fv1smgQIITsBgQkZ/BeNr6IF0LhJ59jMukfetbi7fmijYgbL5ZZvjv9LR/3iGNcx
HgzcBYYZzKtxSxbzX0cKhC11wgoEEovElv5gS7SI9lR2zYvNQtO6KuPHtH2Alqpn
VmvQ346EHdA8721oYMlsxjQ6p46tbRf8LTBWIg0j8bNlKMKrY4jeaFyLI+TN6My4
n5+TnzLvTqfwMsgzUWB+qvku1sh2t9hhxeJcqlyrXzFwgQ8xh3Nnm8ZgZqiXEnxK
P/5ZxHtAScymN+j/5bGGo2OsqsDPOnUUtK3mVQlVWvHaLdADpzTeVvGN17TrsHnz
qmZZoUkRMInKuCgk87IRW60TABA7EXmziQUTXjE+EouOzc+RB+xIazaVbCUTBB7i
zPJEFqN7ZGPdw8xYSuTkeu3VYlXwcUHe/YJu7bI01weU75SK9rmqMs89RP0DkyBN
ZPB4T9LAUkvfwnIFhAt+PMsrfgBEvwt6oHeW4xdOR53bqjzoQ+KxkBpOJeEF7lEM
VAAF4jmQG5DivpZRl0gz9KwA9LbfClGUOt/tD9GV3uqQ/JLkjqJNwAxruZ4kkaKx
MYAuey91nvi0cXjN01genxNQ9dKcAmQ823AVDqBGgRAP+TPPKZ47Y4CzEBPjDCqI
wAUZyNsmaQzcOkOOfiXQQsWGSSdkcaVCrB65piPthbvxv8XA5NkLpqAajFHIFBZ5
YjQewV+x5JN6qDMr6PtELzU2S7p19vRTLs0Y7JS5j9hbuh9mjjgTxs0e1j1lqrJl
JuV79UGvR1HX2RUh/z/Gc6FD4hTIEGXvwCsmN/JTO45wAlQittnSCbJeryZBxssS
H/7wLO7MimtDc/vPwSGoO8XT31W0DQ2oBCyfxQGiW/01stilcGJcKYo2L96zu5zx
0SVr8vqK1VpNwngFrSU3E9ir8OuBFSLNLnAaQBQPOvy2WHysdLNS8VD5PqOTEMpN
J2TKj9kAx+69HfSNPQTak8Inb0OL2NhapCFUdYTGjjLoDrD0v5uA5y6NvQ4BBpiZ
8R9RZBTbgzAh4InccxJmAH04ujl9RF1biBS4YD6bWDzztF0hOdlRPsPA/2QU5sp4
sqQczlcdw4Srnp8ht5bK3EUcZk2H/3LM3JyiQdpdTviq2fsBVG+ziL07kQQCKzgm
YY8/RuYB1mOpwHcPDV5XOkLJ03RoHU09XrsLZN9qgUv+SIsjFOBw82hsx0fje5/W
AmoxmcULPOhaR0d30Wr7ePYgL542NQEk7Ju/cIiltJHcV7SHA4gGYsG6AZr5JUnK
auXJFxJozV4+rpZy1QRjY4yy9c8XfY+v5QQ57hze8qEBYivHRkS9zg38DEj5JcQz
Go+Vy4vBewEydQA8fGfFXOip0+RGZT+oB+YOhXXu3MpRQ0yBh93MviK4hM2JK8Bz
qKdbIGyXfwMo+b9vX3FLNbD74kDJ1vUiisWzc44dE6lkdh3Mp6Sqszar/Ah5PMoQ
Nct3vnr/7BZ0hWWxSEsflJzyHwz8YdRix24Q5H8UNbzgDZCtYRd88aQHR2/+10PL
tWiDdHRzkohmcpNEq3qgG0wwvrwfLfONuRAkY3MJnbxt4TBy6F7wEeKfye5fTUI0
S8ZE73mXyHl3MFtSAH1y70hlFDOVQelfBq4SQHbkA/myc9aIIyBJ3OhnsoWifIPf
3M5xiPGkOsADtbKX5dANadWMm7u1zBHAQUT7COx0AGw0icLgPuiSm28x1PYEkn0m
u1zGjdnkKRghFJxRXD3TG8n9syCK7fFmqgxDYzsworYyUVbvTfA7KZSWyVT/jlf0
/M6wKgEJImVJrd90jr+VqjavF64z7rznyEoW83AEQWjfrnQrzo6ak9Kjulr6VebR
swHoo583vr1Cjo3UYwb19i4HKc9srYKIIren2es7rkQcENwT0VxUoza4CkNrO8xV
HdN7hsK2yJd01i3X6c5lPe+JkDX18C0EDuECfAD8TIjjpVv+UF2OP/HZesuG8ROt
9Ph3qGQ1ltsx6nlX/i2Utn+URyJqzc+rDUrSCxhaTiN3d5hRIjbF8bdjriq/iEJ3
3szFo7w9Tuxh9mG4xXy8JYRv4bWO9DUPwGFK3DoTWEzYHjMNSX7oobtst80c0z/H
s3iQhVH0SLhad7lMfJ1DlXh0hOWC1gwdLB9yZhOBMB1H+37SLI6pEJ4woUn+XKiN
MyZz6yezxhuhbvF6q8GHn+x41s0jObSzgcy/+hqSW6/5XHE0MpJ3XoUU/YSi0vW6
yp6S9ibxfo4M8K/wlikg5XphEsBIAYZJ+QOlBmASH7UKme4JTqekr3PU3DeTYsxe
b5ML8JVQOdaMwy6LeGMgqS2J0Ak/b7ALfVzMULMlaGnqbNg3t2Nm65onJ+XKr1uN
/Mt3PEdHl59vG5gE2F8JS+K0Bbd8Ev9HadggiedliiOF4C5OjasQ9whIVWWqBCMY
tsiyiNj6be+9Ca0t7femaSUNt7ibBuP3oTx1iphlKkJ3nHLWIGP3BHwUuYSR4mde
XapDiDh0RsWBvB+6yGNolfJUWSsnWOLA8XLJBUvNuqwq1cFFAAdggbQ75MvJGgoo
EDJ7WuZlFJOKQ/x6vHjETtEbqg3E8QvSbF0/yK+IhLYX4IXpVWCowzxzKn5TiBtC
gMjZwxFb6nb3qGvWyKVMIIMHgDc1GyuCnSvYCVYo2ytD8aEw9uFGYnsQkVoG1b/Z
9kCcX1187Yp8z04kHirdO1XgYCC9Fw1fuXqGlvzRGheiVVRnOWGLbj1TfyrqQDQg
8yrHNCOEO94e9QF31lsqetHbJZObrxobR7ODmvixCLpRBgsmisZjvAlDg/grtO9T
pOFeRtunv+NGicJx7wgXZGKGu1H+r/5kQHfJ3mJXAEyQJbKhHoT6eEUQLK9r3g5B
xTdouJ5D52zjnRupvGM5M1BtgnFEelGxtY83OfSrJ4KynFe8WlX3agXfDwocK0Id
zwULa1Yp+ldxiW/NyHKG85FHAE0s8ODoS5WYpTrX1qRyxQ/ZqoI/zxDYuPrJVNj4
8wJKvMQJKRQDbN4XNACnMDzRBMzOw8HMoX9nGkgX/qjRVWG0x4kzXDJklDLAz1TC
9ktjcP0g9i8/KphSlGjP9dETt1IPwuBpiXvt/pzYhQNYxXy2WGoCj8qMPi013vYS
76C2Echwr4pjg41OsqQ2Jerr9U7x/V8E/Z7KO7h6rbzHJlEy3RahTdp4J3W4WLgv
QG7MabDUCf11JYwdTKWV3POPi1WET1EenjbT0MCIh9cWaPrKZVYMbisuJO50+KIK
1qGdCCe6Y+IT8QSnSexQuL5fAnWMDBHenOWrTpxH8HxTZKUyN7rjUdFXldpcqjJy
lkq/OKLYLZR26UmHlPi9QwFAdCNdqPvMSL6+felg9wM//1m+uXrmvOt/gu6in5Jw
fZDCNz/iB/0oR+cBxNjHqUGQMkb5chiecliEoL9n1UYgdluRM2lxzsvtcxdf8BHd
tOVb0hiafeiGht9rVHAFCVLFR7Nawn43HrRLsjyoPXNl48MSXutUXGveaoREDXpM
5OvMwQemaEVIvyXY84/rSU/Wj2RHe1nHI0qojFtP1OQA/QiANwXdCx36l66lF5VZ
Q5cD8sU97Lrx8EYDQHDY5NrzPxeefgpbuBv7wL1OgK0flqVV+jwL61EzFF+NaYMU
7G/uHqQWYA7xA+uZZK4ud9zD9R6HC51OpgLVkD1OTwzc/wi9Rlg8piHNoZA6VEm5
aada4L6O490R9N7iEAZ+lqgzPkRGBFUXb9etuz43gcx0VguaFFEjWmswHrx1/sRI
WDimBS9KTFAe6fOkKuQBggd9Uy5S+SR+YlPncl+sj1fHC2uvtjkcS5aKhoDLmRPm
khkrKAZUeOcE2T97jiyv1b1JOoeP+9iDg+9wdKwMD07vj4DtD5Wnjkv5I9occSNV
rPiRvhoTYLWoUqzRbkvwKHVhi7uqTMTRESeUlaSPA28g34zR85fqtq/3jbpzDqsj
Y++1qWj6FB9a+ecTw5lV6tYfNUTwSNU/YIHJrOJz2NZ6+2Hd3irtGK3h3Qxgt+wF
bIx10dcN2m7GS++VTXQ7sJO4K+9NtLI7JFHvRaCbyAEXrIKdjvZ6kgvw/9WmN0os
0D/Rgb0vIS/GaQ0bmuADMEhuY54XaGTJUiYMitJRtA10NId/mj1It/pCD0Gwxw2J
02rjCTXj+wEfssCmyENHnUL5BIF7V0xfVWRY7j0kDRZz8BEYYpVp5bcmHVW1Ty3Q
t9KwUVxqK0qJ/Ofv+XVgoD2kbmA+lR5+dFqo3/GUHtNm24Yp2G5K2wXNT0zGOfoz
dmpep5qQYxctTFdCRZdRvfKewofqUJ33VM3Ou2RqCCy13KcddjXwlNUlDBu5vTfL
KSqHFQ9O3u7kkYfLgH+veWQEIO/WVa4KVodtv0MMSI7sNJ7sX/9tkJQI9NRQIVpC
6RlQzzsWtwdJns88TNzAcoct/uLHfpRgwrDocWdkRyrDrEfGOtBDMWwyfbwGtM2Y
/pmgcwL6nVxbNKGWurFurzvhWo5TfyQO9Pygulb+/s5n5ZJSnSzXf9iReFGcD34O
tRyU6VllRxsqRB2JciJCuVyOLVmgGNvcLjYFV4+5g1cavANU463iz8QWpFmCN660
QYz4IasA495jAxvismBkDZ3aYam94+LJiTqUDbr1NwV/OA3WlPw1qYlKkcJEZcGk
yOjeVtEqK6qcITnTT1ZxhoSVxdbcvToet44OQ5N2K0UTQNkhR1WSZMF9ZbGinmvW
T5Mov5fFDdMjoHrgBnAKXQ1fvbdqoBqlwI3rPVqofHVwR5eRxEYPTY7aVCmsSKij
aN9MOUYt0XC8hhOGiKC9xQBWlTb8S9NKzygKNAipsYmiKUlGHi8mfJhq0ymGU1DA
paQY3Yt+ZoXSiinLAlyCG2HQIZJ8QzyBgrqHuujQrSInnjkS+R/h31hl2baOEGUw
LambRjN8R6yvpgo8EBBfUl31TBP6HvlAa0i58JYHAtUedorTXoEk501WtwUaQ85/
2axM+pY4OaXyR1UCLKy/Fd30y5D2WEaHrh9NhKvCpX6IJStuVZqdcOpR0V/wbfGM
nAaJSqf9jsAqunF2LrtVa+iY9KprCYCT1/onUz0cyG07VNv66aKoVdzhq601L9aL
GkizVR5QWGb031JyKURzx70p8SyYI2BIRO6FP4bKP4/QPAFLhf0nC9LGAICrucVg
MzCJWZu7lf6t08scQ8TBQYC5mrkp17veu6r5X/Z0r1gKeIxtbiKDy+DFjtGps9Up
zI1pCerHSwndAoaiUzZw3X8JVVFjF7ffF0lJhd//ANhGE6eM6HJjEws8aobPxmSS
kKezrhX9nxQKIpc2lL3toh2WofA3hFVEcnGoB8bPIBcxtxb9SvqbrZjTwxSvKQok
NoMtk0YloxdmJoo7e2gCuX3FhMkgntJK+FULMjGtOPYRRD4t/qiRKuwJI8FHOMRJ
hNV4uUHLjjkt3apfcUCi+1qgK0SDOercW2QNXQZHnHDbcnz1omOfK9xNCEQDS2sX
gd/SKV9GBnp65KZv0JDghEzp1Hmu2ooc2JKSVwbqKf4aD33QcxjmoiOKVHwME11z
XkJFugDQCeah7Wvqy24B2jsuBlLs/de09OvylelNTgkjnpZLHjncAFmmYiWdeMiy
X01PYpxsaJ7XMFDoRM8kPyhfsF4OB0m/dqiLqvgJuDIfQ+M0G2o49oGF7mubYdpi
0kYJ9y5j0gkP3LNNcGjC+ZOPR4fo8UAT1jsKBrhhM94qlMK2CJDP+m65EPRprIAP
6pHQvu1IPG00EdnuMAYu/6QKM5+BN+8VinsbWWhmXNuSEk73vWDSvCSaHtMIsNIs
bN0LCx071aeOo6xVcFk5gNcWG4/Kh7dH0BFbNHOsI71C7UwieArIGJUIj7eOgnEb
vUSZi7xI2z2cIXOCNgwCQj3Sog6UTEvAbu3DXakR/vmZLBZDvkc53HRz9QbTqUsM
/6OQUViD/JI5xYo6dqmxcrwuYqutskeI5YW3xPDDl4FzH4n7eeV2LWDHvOcu1kbP
OiV/ORLQWdWQo2AGxDJcWd8VhK2uIH/NyRpLJNAOPzOY8S/COfsdy3iiwIGxv4TX
ctCkwVWmYwmRcpLzMGbRcQ+phP17ZSdJlHyhaImamJaqOnJqLBiOzXJYohGsBViP
OOmHdwOl6+8oHpIff3ve8YD0QCZDfy6xU0GvoWdP71RrwyEAZGSKCRy3Mcw3i7BN
kiFxZyfj3Qm9pSt8gFJd6OFRSi3xxp5wAreORaKDs66Nfh6sKQ5cPG93IFpgZGGd
qH9sPiZQpED7ucTGU+yVCZNoHJzt3oJizDlEMNsYZBfFNVkc3JXBrlQA/SBamw4J
kZciTC664bO2PQtFsv3Xz14lXx237Qan00nx2+v97AQoKm4c9ujAZzx8bOQNYztl
ZIbK60xHUbfO5gra5P0KjHrqAwAhbSX3hpST9p2/uW+lJuu2PEkavzur5I5SZwTR
N+DgXpSvgO87p16wN2yxKuFDLJGsEOyAjp9wicybAxy4jYw+Z42skP1EtllojBb5
I2N3bkW2KnZqzWZzNLIkg7lBaqi0pWj3/OWkZjINd4AA3cpaoFW03HVboxPN2WWH
h8o9U79E4dO1M4lBOKcT+V8HHhoI9a7BKCj3zavHMB94OoPeNFygg6cUf7SQRK8H
QaBiZCwsQUCNL43+Y67GU1+TpJ80AXcPT9JVfOA0oFZjtIXrZFnj0nWHleasiq/n
+S9jsP+LQSQVr7IDHCWtIcEGU0txHHLatKy4o62Q5JuUejEkPeNS30R3rfTWMcp8
3LStow843j0mnJv028+RYuG0PQpgGuRfEIVn0bHR2EtUEErKOvX1mIFNCtK9iuWg
NvKcuc4lVnHIJWdLV7xso3uh/A5W+BwEU6pMxTUJ8QhRUNjVb9IuZW8cs6kxX/1P
tMcxl8neqZ+T8fVE9LMFJB6Pju/dz317qhVtPFxFkF58+QA4sU+V3OAJACpVkLpN
jHIuQWEx+OQzkK1pS7PuaB/XM1VTnEsFm5bgBItTGA42yIvIXqOo2+Q90RMrxuL9
QSQZJ5khNvhfUdWMcCjJoB7SkJmUu6Nqy4AranqoeW8f5sbAge8Mhodj7AyLl+6z
GmqY5s2OPZghNwkIBqUnQBrYGik+LnNEZQDHbH+K5r6chuohNRrFSA/m2ZgvUgMA
z46b3KejVT9O/ziitse83ToL8vERnSyCPziIwDy9ZnSSAZ2Ps6BqnHZtpCex0ouV
5vLlm0HszZ1+yFp9m51wZLs1lLVTPpVmzp1QmaFPUPQmuVS+mdzcAVZql7hcH3vS
WOuEpIk8F5rmTe7AyCW4hWCgG7TjzJAHGHKX6MAs5Y2EYxn0hpAY/ja4e/I8eRs4
lBlIW1dTdUXfGMlnf/hIUnjDqDUAsJSIzp3a/IoEQD5QWFVwfJKFWDjrEaFyPMdG
Xmqfr2wgRyV5RJKPvU22WIdhahjE/2Zgc5hXRRn1Varv5TmEnSut+Wwnmpj7pRwl
A/sbXMahY5pK1tOaolx6nBTg7ozoFut54hP3pEz7I90rl3tt0+d45Mo616sg5pjW
rA9El5/h23m48hETOrA6xjBl+cY30DEleEYFz3P6jC9l4pAC8ORBb0kmFsH36JPH
OVRA0+kJoaRakqsAaEK8XRFC8pIyWSH6uS8USQ0A6/7wyw1uEiuesS/hbLhRfiXm
D8rtiKFHs/Pd+cXEHPbpPF5zeojDDsWojgBsAthAyejW7jimEkaNUsR8+2Z4R06z
8000vZXxBTLE8zJDqpT2bAtol0XOU+KeIrYD3QLOMOZz78P4fhm94J8Z1crpOzI3
lsGDcXfAz5rMk4LVQfN9xHg19HV+i5UrYvJ6mq652clRt+5zDqHYh+Ry/xEkdNLZ
BVT6vGy2MrkSGLl0UfIWk5c0/pSevVaRNB2LDKG5N/9rssI0fJXnAfxARUp4bP1+
bl3obSc5p7c1GP8xe58BiYIDk8HMXs2jQAD5QGQd4bfTmCiija0kUihHDrXGnwpp
SBVDR3ISgCLG5f+WYndfiq85eTpndN4Ym55D+X5tDT8arEv2ToNtj7joCZqxtgP9
yqNDfsQFj8uYsu3EmWi+rnJxNe2JgIm2WerMTyLhTuyI3PmZRxBIQjmVhEDhk0xU
0FXha/yd1OnJQ4ormxsSqrZpl2bsSDvJ6LiSst9P7ds3CclmhNEUsFkl4rr6Lpl5
3BX5yriEWUxqVNJ1PD3tsxoDS1HK9pBbusmJiUAXUwQE4qjdpbIMsaHyDG/eL6G9
QP4Ss8pk406cl2+77aSqPQP4fX0v+vjaVRhxbwZ9RV1CwOEAfwjUbYJY4lqsv4MO
rU7IP3RvWeQNjxR6POoXHYUzHKMT0e3pHPdyEmPJumuGuZD9+6PQAOE2FBx91JEp
68ntUuz/NbHyhJEicma2Eg+oze4+SokFVsggmTj3jyfeiQ87mfAr+HWCcg3Wsmd3
QZJY6RYOwUiNUJW0fafZgr2EQnbobHCHifrf8iJkfKEeD625B1QhvXlwlwzj74zd
gsMI3D+Su59DbQAr7C6CLxDRKzo4ufGdgHj40XBEkPK8fL6cFdz52S1hXTSGSttN
NkEB5HYtlAWn5A9xvtIaeNVqAl5dmw7Da5/WOT65dlFVtaPJSca8rkQBFGVJ8Vep
vm461mGZV7EwhsIkJAZWdftZ3uvTCQ3NYUC55BUL5k/4u/I/ZIbPq11DPRsCdTGX
3JegBK5fQiccauVVGthGV1EX1MrJ5A0XuV9M+PCgZABzdyYuTTvK1HDFFT0rWan0
WYUPuUZLnzQWgauWwf50AeCypjAISTPAr7t6URv5lcas6MVKPSq0YsB5ltlH+luH
fVG2UpOhyqyDrQ7xmvhJYg/w5VRknRo5UDxCR7QwtRbLj5oERH1Jxlq/vQWPEhaA
9YlJwEAmZa5tzJCEcr0eoVDM7zOtW9PGVkcVc5bH9NTRd+zoORi39eadpum1qiHu
E47gmNvez9fkEt+NMdOtLr3poVIMu6qF11LN1EVavUVarY+a9zDwncQad2IuJJxC
0CCwP7pLNt5aMSz3qI4ycrBraoPpwbVEdTY0ioZqTi7LqBz8mRvZTN+ykzGmARKw
hGMPcrAe5fhDyF7CDQoIcpISHuuvVUvoa2m+Z640G5nXIp+43ikIJiJRHmbhRYpk
3vewHr6NBuDr6+g9UC+wt5Kuwica7J/xiGx/GPMYkKJ4qlapNYZSb64I47ot9JSL
UbIy6juwQZjjPHt+SOAjY68r7JRnd/OGyPV8w26+GvP4aIX31GENsANI9UCdEcqt
sfKjShs50KdXTJIR5K0lsk2M7SoZW9PIdYhyEXc71cfAdOXpFgEh4AR+OERGIh4v
dTkni6RP0WIDZP984FDIMIcREy62907APTyOpxtg6AWGEhIFtTNfSxnmrFVU80HP
+QcEth6vV917qVfJk3BQs9YUIbOgMTXExLULtzfCwx1Wk+h92X5pyqwT98nml3O0
Rx4F3uticKErTcVvOXqkPspph7F/XIl+/syw6SfXSFc02+sSWWvCjphFFiFHpiVu
KllspAGodzM870X65UqOCCA4Zt6ulBTaZ7Blqrti6a8rdC8IXgQGd2Lx93mYjrix
2j/QZ96wusKJXiSBTTN4LFPegjATR8UkHFSpCWZZHPO6ktnE9enjWbhM/0fp4kNc
1kJC6RccIjZ+vgTvVngcIoTRoMQK5vAxne/6/kCvQKAILq30A+ELrCae16gvULGd
TmECYgTV8hbVFnourE6S4egyFjMnkc76c4ixkLYgshMQo1V7bSIEl9J7qTOvXwIn
Tj4WoWo6cKZex11A+/zqXz4JVbIiO2OWbcZlb7htHYT568Vi0KOW2DgxyoXJijb9
BJwNhDh4KImEy1gtPIoAO3wyHIRXfvkBLsoyWdfYl18unpClYOS5L7U5XR/Z2xDm
eZHGByvpHw4BPd1CHaEPSfhmHaAErJRNA8dOVTw4NPX/6dTAElGhs6E8J2Og7kVZ
K1Lw2Nrcud6qqwNd6Af0GhHd5JnY9QYp9humFAzv3dQKiKRfROoieMI+8d05AA6B
JA88wN4gFi5WeQ9YGMrFqFc4obf/nTT7zYtDmxDNDRlrYUvv0sGHwPHjZrq7qPkG
U7xk9jTac4hWL2RMnZ/ZDfuYcggpijb/FYaX1vqAhTAUzAghS4WCuj8ARX35g34b
Wp0GEtUzZczD/xcIpsZmydzirt7LUIvt//KEmma1GiMvBQoUtAsNBnkC/Z97WNqe
cQUiYeTahcsXmQxCBQpdAOEMwydQfeH2GFle94Y9AxXK+o0ssIXhyKX/+Lqod6B/
s9Ltm1f3pH3TeZaXufwmWDnUJcZoxiJtg/SRNSKlBmT/Eo9C1ZV9AHaE/MFvMCX/
oltCMQBMHCPaKlufF2I/mcOaxUnN/ahiLJAcDTNjKOq9EmIflXqme0TooTRqdyqr
ssDbpNAfnbtHqU+E6ebaNhYkp/Y/PKarIl89+cBhf573pS+JZ/rBmoWMMeEwpZIE
56K3JE1MTA6SnSGxv3P12SUfIPKFknV4oyHqe19gavLeXpyxhApI9vYMV47mvi8P
YiNkG+gqRp3/NlegySsU/rCNGEV5xu2XCIbOaeA1u6KAnS7ulKM9pOMvH7jr1KdB
U4xt5+2LxqZIqvcntwRpEc/TNSezDiufu3CIUlfxiXhGD2BpeF4ppc59XLWxFskc
L9mf1eqXKL7pGLq8SvAOpc59nMbuPbB3IuxmXrj52gKCxCVqw9Njbu8JFCAXKyf/
D+uicT5PKN4fJi6lglfrfq0N4UsI3YTdxC82YpJKcOjLIqDmWTjC0uiOY+60g92P
zCy2XseZstttiPwoGd+owqqqC9xiV7Ktga6szBIFT7HSgUCNc0+o6b0/pCNuJCna
MjnzCU8iefcDyDi9cb4E09fLpcL5htKnWITBHtVyeA1xdn8h4zzwPG7Z00vf9jxA
CbjWT4ozGC7PTSEb+kAR6temqevh5o/HUlBWDAJCdwoN2Iz6vBe143lv1ZMQf22R
efwHt0mBGrIDiTxeqqMdq9p5940NL4z/honluFX6zxjntSnCjVAZgbcYL30Z9Hp6
/XxYDEbe7PKI8yhXXGOWqPrvzQnpkKKwJQvhP8isuVZm9rcIzESJL9QdKSXUhEGw
oqUYG7BRVGYyKl0FeRDZSGGihPOpnGFVp3B5M8GPYvv42n6vsXv/wN9Ki6okafie
3UEjtQ0qEgc7A8irkCrb61E2totFdpabCCLYDwD0x0aJqck7qA3g+KSN6LBkcIbt
m4KDiFOZuEC4T49afZdSFNE73NmWYFhgGptsEzyaZokaoJJpfZtbSWuDdHLDsypu
EuKwzckmhaK8ZszNwdQxe/rPli91GCEgfrQBA2UA07bSr/KY2rlW9sq4SfdeScM3
JxRTONEucDBexXENB7zGcVevf+MhoPzbUpoQbIFNVEpxarbAxoXfrolowYZfdDw6
xkwM20pYgK84zjJWSoPVXoWHwydyHGdHV6PXbnxNwpUfqhjFFnt8IcTBNSXTeb0i
xPLoo3ZlwlmJM1dCKYvaK5v0Spvh0JqnkcZyy1ZWFRk1E0ygzxWNxHWDpS8Uw8WW
45FlPcyyveaMvtcETOb5kLK2S0mru1KxaHLGaMEy5We4Ngpb1jEBuisEQDhdwoCA
RmdTaqhM1n/btI5qevbN9GO7sJNzVAAX5P3IIHhig9VKZCKd5zczSlAkDJU1m8kW
+iWqdLIpd4pXW7Af0VVQox/4+UyVcYtPB0IPvrEohbIK2C1ekMLNvOSf3DWzQ2kw
/sNhTgpADYuyiMFytKQoPQ7jM+VJcGFPv21n1YGz/HEvVUyCHvEnOgy216YtY7AL
5OQF9yAk6V2SoiLSYxE+p4DO7dgiYjnjCUJBkCUmqrSNIz84/hluq/nBQe6uLiVL
nQnAHFo80IPbk03MZ6a88mlyvhi9Jvyw2UULQmQh4M+0RSE5noNc08XcL8EXmZxx
4SNxaxK5mB767GCtGwetWHr8IeT3NVgCkr4d+YTqhankFtNZVjZzJILWvpoAOKiT
qu323rf0NctCTVhTsS3VPEgRmuHj9wG1YyW7ol49FMBo/rCqAVZKQ2UW7qmltoEi
Kzxr1K7ZIKJ0wEbUtLsv1cgfa7Q6wWiVPFc4l9/vG5wyEwLJUD5C5WwNeXbWsdQj
DpKSNTd3Q5HV4YA7N/7qDQQRqKRyDuIVa0omF0N9ayGx/fwVcoiOdVjtOxBW5/rB
PHDKMbtfaKUgs+pNNb8EDcMeJYB1zeg7PCE2fCFM264IjqNt2Hf5T20Q/H48ih/S
MLilO99RNeTfQskBACSgEN8/P8LElkSwc9R68Fb2+mBOg415BcvdIx3j6ktrIkUh
TJDLRLydV1USK0IqacdVv2mebUPHnGUisQWmv4QrvSXyIKwFMNAk/sdcIwpABSwm
bl7nqfAMatOWQbgolIaiqB3HLz8uXD8xfA/nHOniHY5EzQWs72JlqwAOgeTP7rn4
+mm/QStP2OcHFtKHc3THz6qxXgTvsYIvfjrZvCvkV3hOSwwygGgj4H7PsbViEBKD
K8wx0wTy+rcjYYADsreJbuk+z4Ctc5Ca3hCrYdsMzP/ARsqU+V0YVzbTmvwp+e9q
RkLhUKwNCuuogz1O5HfxGK7zADc6Pz16DPCx3JRshcGb96mVeELptgYNP7+DP0SO
OMlOGrLPyfTMy87mxOTwKjDl5a1l6lnLWmZdfyTFDtSOFKXSTyqJxDnv0RRmD1FD
+KgMPnFze4woFSrjmV5eELZVuu1fgDghurYVpDeXK5Pn3ORpCsJEwmBWk1Nx8Lmq
/Flmn1j8ymBdjygjz8zU7H8L8jJFg1P7DWKha9RCG7cT10xkVerPyCYbcHR7JU8B
e8uunz1M7TcsPWYB6+a+5fJ76vcUyrasZ+PoTnn4XiTR3TvJ5hc9N/WC4zzqZyX2
4UwY5HwW0Rm8YQUTr/nGKouVGmk5iQ5fG1JLOJ3MYwpBFJEHiv4SDWE1yNZSlyBj
Yw4TrxIXxl9RbNLJQ8FA1TTIrc9FdMZt49FWjSTX6ufu4La0XXkThAkhN2ZD9FZk
cU9d2tKJqA2leG0ajOXLVZB9/crGIdMrbZIkxS907o1GOkiJIpn/bSdC3Gaji1Ab
sxpDffluzgDYLBk7qekNO9mOZA7dpA4NZi+eHpb/h3NqX4sXwdicC5rPa1AtVaRY
K6w/UPrkgFGPlfD2La0SrhSHZOCo/y4YRgT/l6p5VQEgh6n4nOGAJ35fUuTzR/aP
54oGgUzx/OjDBZo/Y62YuIUiTVMUxmQrL7XYs4VLChUtH0ygG3dR93z72iK+wPQv
DHhH+h1VshnN4pitsed7Oe8EKvWL9Su2Bmtba8auD798jxcZsmFQ87tbLLWCLSZg
k3uMN0Y9n1nLU2dpzjVgS8MNcMiOo4fzWRU9O5lWQA8vezvzYlQKxXNgZy+jUNJ8
qQwesHji6ruh26Ko2usw49xzzHhob5hO7Aawbs5XRLbZdbFsVLm7/HiA250DjtZo
J9eSEqWtO2AEjQRSiSQjmFaL/Fdhd9WaRAxD/VhGdUtHRmFrd94idMBMmbYW81gC
yxzgpK9vGvdvl9ZIxmbUhfnzPX+kI42H1xRIAYr1NapdKdSUSDWlhYqa+19x3pvZ
hvYduhKRycb7Q8LpVt5DJ4lgcA4Z55RJ9CTDlVbF5ZF3JKt0hPuorqEjEqWy7Yw7
8/3fybHP8gJwC1qoDJ2KyYevYuEEHQUlXTtcUeZb0YBimnzscv9+gquG8+Nh+PR+
e0MuMctsZ+aqn9J4H2LJRpzmSQr+9lzXojWU1H+npc9Av708+bzUgZAv9jTmeHPG
DNgb2DYr/ngJSLenoiFPReZ9DM2XX5WHHEIZtZ085BQOPaajqGcYuT/O+s3xYIvk
h80rlUhJdUGFs2/Yt/LpzwE7h6EvLfhgzZeVZxMOmUXaGj+6vgoGsl1wBysxBao/
VmO6ZkWHLIEeqbku3qxC17PAio/8YU67lhE0uCQYDydZrNoQI/IyE5Hb0xpUw6lr
Y6R9tL5YwJOzsOskeVjvDqORFUm/tfrz1LvA068duUFYlYNDXCK+MFQL+9e63hdF
VlCt/Pazh4ugFPWTdb1ifhsPyKRng8xYr2F4RO57sPNczhFZOkf1y9/bOzRXnuUd
93NDq7RwU5oRTjcpvtlD5F8oKcWBOVaMAsxXm27AUAtJpxIfJBm6iDnhO2B97uJB
EboLiIRgKDsH9vtp7wn4NWJZMFlxlV80Yifs9NNmImuzsxnEtoSUvBIgOfB6I5xq
j2N2XfkNp+wXlhhoMorMsOOO5JxreHh+3kWgCX54HWREcnSQi2BLSlTyuLUw1WuU
lXDbDF7lhlT0FMY/oXhd2lV3lu51QOleWJ2fyFm9NtmYbznraqhZoJk6FwAoqdW+
Qy6/0ilz4d+PoBeYokLrclrevY1jle7h3aI9qL4I+zA97aJJVVsEca8Bl+KDFbsr
59ntIC/Nn3AS/x0sib+DHkCmkke14qSQ8G8c0LAlRbXJqcDNs4DBpD4wVawE43uK
DbE4PwQJSJVfBb093Ux3tXLeW5GDaIMbK2Wb320XdStc342tM+/zkJ45gxUGr6Cd
EyU4vuHO8oTY5OjKuejpmyvJE/mnzDICaZG1QPeizYQ002laeSh8B953msrUo3Uu
8c+AlnKwYx+3028a5PyUUksEVAo1JtASMmib8K54cTXNZwirNtZ62Yug0aRbry3v
UdvyD+MgJcnnb3DaIJTZIFKt3oogxW5F1HZ6iMqU7M08Xfwewd+coEaRu8rUwZSw
WCAtmoGfQkdXm1bRDnt/yQLGXjft5d54On4LM6Cj2SWYeDkT4yn/65XEzKEmnKYX
KjBT9qQbmHnThstlFf9Ui5SVlMwWgqKUE6m5Rni1UkCT9FcESI/JZWGIy4Un0mNQ
uJ5FNAIn92pcPneX6Ux6Lpn0poC5YtWe//+qhHXq75ZvWsnyYShxrAUZLAAULnjq
m0LA2ULkiEHwnfCiKR2UCXBQDfx1uSjOZDiimQCqSdDCaeDsV6xp7KljRHpEQNMk
IWnN8MkdxLUEQKZRO8zn4scSTByOaYTLYdvyw2kLHZvEXCSdSIHcYHuj3G8AK4pe
1/t1/qjW8abPvmd/UXhn5z8eFYaCAXRzJ3eGApCAqU7kI5Ouxp8TneGLyYndSMZU
pl8ouvKe5c++XzJ+7fMNmXBggsx7dtaQvwKmafVUtuf70HvaT6zsRhESo2LMJSFA
JTpbMsXEzY4TRSSS2YZlPyFfOJp12UvPoy320jW9Cy56LR/xxVC2xGtRtBHyDuDd
NNScYGz42IqWdB6xn6HiX5CongKFnWPp2OjUDHbX/fPBCIb6L+xcLZ7doFYsnJ3+
2hD8ACCZF/A/ab9ijwHMVA2PQDiymo9elZKGwed2k5aILluuCGVFcKZ6eBVBhRpr
jhH4BBaZUajH7xNEQcLTHixRiGYfgyqKNiUrWSZ4j7NAO3uINZqSZD0GI/hbISLB
nDycovwXV8Mwt2g475GDFHslchTyGGVTE7gTSFr7lCKix/Q+U6yyC5I5gG1CNrY+
Za4UnHte0B/lBF3CRQlMCVY5o9N5X7NRqq+beupzEd97Y4UvQZZ8MjBG4Tf+DjvN
vThDlKO1BYpPXypghguwDoLGSYTS6eo+Eiy1z99SePluJF5OSXKJ8p1HJl+4JTHo
XVUsnDBe1HiViPCkkiq74VIHec0RzxZAGpEsjXWuCoEechzn63Bg8aOoY8je4fDg
LbJaX41CwQlYG/FWh7NXvB1PzaDMiVTXzNK5w4Bb3oX0zZ4X1Q6ca0wDRSoTcRT9
jsqYVaxQPS5GilSrZMVCSOPYZALnK2OS5Si8M9Y+Olq76/Jon8H5YBY58zEvymLw
cRXkfdTDgltkbpNQC2HxrjGb7iaP4ZZaQcmEtKe03OTttO/ueLWp96l4RVc3nyTu
P0ft8eUTQljbzyKg0QT3KGx85I1I2dCPBD181808ava9/dPaOLw1gHlkH6FiTgWr
3g0iQWkOuvrKs9rwYeNehfAUYRe4/RdC64jjNTKXz1aoTqhjo7lmIrXoZQ3yoc7Q
SP8xXiEZSHk9yHzmdsBIpJLkI6RVynDnqk8SCJjaf63Qw9eLm9gctGTRd8wEV4EX
vwxJ7rs0zqb6XAd5Sf537LmHDuoZDgZHyAZobgSuwciSAXsOkhb6Fa+CzllKn7oP
NVZwhtxOnx97oCxK/JyVRxpmiAJ9O4w3ZShDiwQGztSjDqATwjvOt2vi44qyZyiQ
8SM8yK6Ql4FVOkDfIOAVC5GDCItTrx16CFXtvULNSnRU9HJdOUawpZmX3YMY3/Z4
IkoJDQBUxI/wWWzvHUB+3epEpRheWP6pfPEYRJoJ+zO2kFRfkSspkcavvRzMf2ig
KBW3lG6aomKN1MZuSkHnsSeIih4hdzoYWWyb8fcWHM/KP98U5wXNwGqLG5Lrlejp
1s2UEmBVV7Yp5FJ9OXpAc91l4ZwYS9e0HQ/AOHlne28q+FQSZp61/w+DR/YQuNT1
spTF1VgE7InZFSoUgxBKdL9lmE2gtHWqOAexq7bJjaSzZ3VGEIX0EfhgzReWH8pG
2vy9+Dr9ByGFj47NkVDq/r03MA/n/hMoWH1SzdpW6JC6BI0IRtMKVw3LRz3I6z3W
r+WAvXoslxI5vUJFTdweBJn8ijNSMLw/IsK8VoO7D2EqxD7ikp979VLbRtXQP3/D
uJYjlxGCgJ5nNBZJY/7v7Cg/zBdyX4DXB4gYb64KpVKHq5xQuh/txQ++L3goQpfw
xjz6kQmZ4kiCDngreQO3b4yuG2ei/hkcRpt4LqFFP7wwmRGO6IHO4hXhXBQh82Kz
x3ca2/i/t85mqH9aOatX/ddL7elDx0r60GYCK6+FK5PyJps3u72t2R+iEyYMDLXt
OBSiSHOG+TtvAMDqKroqUpG4dV8SzVQE7tF7fyGBDF71V8BUkwNfOPUb3Xzr2WbO
cD0+jl7ofT/tzsCgMTdSAFfU6v9EMZQb77Hm3+9KDUYeHxyUro1ajuhMCC4Y4brR
d8eN8XzfB8XGVC5JRIjuun77yM4Ps5TosLaq96HSigwqN5YcO/++yJvznd5C+mAD
xt2mTFVPPtCjMu/riHXcf7xIOta6QlupqvbvtOEWhoIvW/xIK2F6fn1vcQFiRu1w
slxD8vk8Aje8fdovSFp2ccHORS/tlK8M1dbuza1OC0SaEcHPeQLxBP9SUZigF/Od
YQxzdFgdVBRq/AM8S30Uls0buKv9q5tM7dEmKUdV5br8hj31iGhmiZyDkV22Yjk/
AR5T5+aicx33ser7XhNCaEWj2sRlGC6QmXQDubWBBnwIRyVeRGFEpTVPl2szxCU+
/KdiFsny1wFDJpiv27xpRcoakwCXar1ASI24SxaqOPXJ7E1tzRY5mIOzdznvoqK2
WONqjA9xvZQJymXLJ6BH7DgbFQuhTKSrxjhhQJ4C3yhWVYnVTQVOsrkezY//Eg6A
qS16TaJknIGFMSnntX4JwNCHL/kxYVOmJZcFfQf9HDj6xOw7oN3X9p32oNHLQo5R
kQT8urDLQIiycZSViSexgAMjiDR/DP/0regjnpDKaTfadhkC7gUPX3VE+8FpqDxS
UE+haUJjLJgKU2PxD1yknCDhcxSO+D4bBCixJs1+RSNxyrdgSxYhOkTa1GugXxpA
kkBXX3fs1pqe0nvg8fmyL299ljVWQoCrqtRNTps2oCZgFKwxUOXNXGG3PkXCut8s
vmvbi1Crc1Ilq5vsPLDHMnY3jVnJ7Hama2X7ETlmytITxIWaISRma8xKfcuxDqq4
hb0rJ+u8IOFcmZc3BquAUgQ3Zs5NH54RqW+b4MiqjFepuW9sCxI3VLAwda9HaU6c
yIAYsOUmwba8MozcibtHEDMtT/l5tnaCoEJDdLEWh9zsTldTYQNRO+0ws8J7Tgl8
efxfa0l47oVdElULu9vl+YmW74PgTqyracDDgsfWU6Exq4OO3L9oaYnfPJjkPUY9
wquu+9AqRW9Frxw+E9jMeNU8q+Iyug8Bqv8vh6eIwKdSQaZwM+niF2qt/0UTfgPD
vv874jLyKWNAc423QdFhhEQA3AW1eBSHOKjZwmSwXrJf5IWRNfC5f5ojuAauurTc
eS3FSMk/yY+S0MyrVzG3O75HjN8+bLBQYG70br0RbGbe6RstixEGO0kjFUyQPE8L
3S7YJWG0epZ54TxZ5s6nHGMfYXRazX21e8wp7AkTDmZNuQ5iWAY4/ZlHiMjd8SRG
5g9O0C+fb0Bsd35tPBjyO+6aGrc1rIdZpLxm3hXrXqomLrLmWyUzYyNKxv3MeXRg
UGDCBabayiG/tQbYwn+Q9yovx9ODVxB3Ca49tOSP5hW8qYNgUbpLHRj8467ON3c4
T+Sbg92M6e8QZQl9edHrmkt74H9zlPxI6J7Ig6jIkGxpPXKgll7dy/DbmOmYhIJK
o39UiJVy0QKIVNmhFTE0E7ylgLXc0qiBQBpLGK/NgbXuuL7ZsUSGEShQBwD0REoA
GSnN8nCNljPE6bNeTMHecxVsLbY3XsuQH+LYmX5YGBBIvhW/QUaZnEaxQv0dr6+5
lS1qGkav1Kor7NN+Szf/F+727EjJburbTnmXdCeMjabpQhwDKoWugnBTYXisBoo3
i0DcIrRz4SSaXYjiCsy9I2aEGoFa9pX28Vw+pzPvKfvVl/MMeHrW2SgsPU6gxcGn
bel5hYhtBLS7g/4MewRlCFs5cyYPu857lRhKplGQZn+Pnfckj1rNx6sNXfHOxPN+
UwzDLpRQalpyQYBnkT/HC8GzZTc0uwbYWQponYI2/XY2Gayxpkxy/4iTBDoXZTpH
GSL13IlwdbKxQ9Na7FcmduyszD7WlC3glKw0cFQj9TentfW0W5KiVZp222cQBYO4
jIagJoyzL4z2olH6s2sB+WXkSrhtTpkB+tt6YWleMtwhFHS2JH9Je7a6abDZ4vxc
kpiLzFp7T0IopTyBvksH3X5rB7Tm5T2ehgMYbEv25xCIsOnUr/00AEnERvxGZ+Wl
y24zbNoOxD6qYbLWJVwhNNoJf4eb0/dzqD5uoqwmK1bflD8TilD0ia8oPHg4FwhX
aBCE9rkPpFqKJaEe7XmxlIuPPYleU11/067t85+vhzCSAnpxbqCUFFrP05Ah6vvF
XnjrkdFogaklw1xpA6FrLLoZzE+BFhrb0U37C5ExDOGJmtp+gYTVJCNf4iQWw5Mp
VT/RmZA7IgqhPM5m+81uZoId4NPmVV0N1/ZvFbCApmLTm/YSQXtKGiS1ucqv2XBA
2+1fbXLprMybSfYLWgf2BquzDvJJpdnRJaTnxYjlessOXXDMk8EexC2WgVBA12S3
bMwxW/rZp3I2WTxkmNOr2BTnWsVnm+1cVq8faxaCgrF2IBHSrEXNPTDTP1xBncgE
F4VQzm18d1TBwBLIWxSB16IGBbfLt7+6vawB+YgA47aj/PFmjyvGm9KtyBpQDGGj
gVqF+IowItP4VInzT5uMl2yD+xfv3/+RX1xEvaMML/iFGVbwvkVPSF/V2pzcugz2
skfACHjuUbaQVu4e0gFy0BjkY6NOwsoa+5WdLXAgwaugmSLr8UItHehdftcQuILV
k5HfIg+zfy0LkMnIRRXn/9pQs03+947QBAjchYYNz76wya3tQ2lGTek6IOZ3x+RX
ijeEEatXIvR9O0+gQboZZ/8eX0rUgBrzGJUpyZnWlk85Y9vrcojJq9X8A7E45hub
ImJC7z/Gi5dOZZyWtpht+N4zDlXThqbEFat9i7j8Sf3l/pYuRgnN/irS7+uvnmI8
k3P9+C93nZIx3kaEdiBbzW2c8x0MGMidlv8PivwCF1Qw8Zulc053hduPYV7NmMpE
PWENBEGb/ZsTTBa67t2b1L5nSOtjASTHLigyrplsvfIrJGRM0FpyALSa0Q16ScBJ
BuqEj3YDoBl73ZqRdJ4oAJhIPUGO3Ue4+PgaiWIWd2JoWUEK+ygaAJ/0y2FxL9iD
Tt2FTQgEWVFk9AtvtpuL+hxQi6j9ksf80Vet+j/qAZNUTvmgaxIVfryqG4HATArt
CjAo6WAbfxMpJMI29K9h/c58o+rIim3I0JIjyE5tvWFJDTAh4+0W/2YFlPehIltk
1CelhM9Z482wpxXw8YI7TquHmR0c5WzlcOq81qA2GlefEAME+S3OmVcTZZ/PucZH
V+ZMFtofZi+FtDFGKFI1497zX/kC+W0OA2In9A2oal/TAzX6eJY9nGexWNLr+YKt
/UB2VUfRIZjExAEDKsQ9F3qZXnyRSP3Czt0Fpp0T2IK36G+IsAieBQULpQgfGGrJ
Yf2NwNyHtcIaREL5ukMvs5Nu+fklUyacZePnljn8x52i6BEXHHp+3EJaxPpYfYMn
19LtMWKw90EbNohxYlEoNliKah8vQvp5i2T4vZR3RyrUGndSlqKYKaYagv+CriFs
Kn2yGj60Nr4aVCHUVLP7gvAXAt4mnDtBHTzoUztNzg0t8JgyuAAv6gfN/6bAL5Xz
JuDBUfPs3qWX5cH6z6QuWRniFxgIrytfqMij6BkxgAV12N+AaD313c4OdN7XO8wm
qPu5gYLfMeno8cvpE7PazPQAkoVVgJjwJc4qD9/wKy9a+OqPwF+gTgVDksOdXcAC
KJPbDBIXpmIZmQxNKx2xlvuwN705NfREsIRm7vQwjWCBk7GGqAh52JfBl2hATkjb
ejIErDDa+HpDaHPdpObgIOUzMSQmgMGFHqcoC4uPUmstZBnwwk1TSKBGUnp9X5iO
FKt+aRFMVqyEozncsSLsXlkwRfQydFrU+k3ClbBUhg960yQ8uaHjZHM3+yHwSxMK
LmP173yGT9tnJ5Bj0OC1abmonE3qbca0T3wWs2A+4w3u49xz1ikbIBgn7qjWjgOz
QZLZl/z1CIONv8VTy8NPyKmy0fSyj9tfSgs4TQ2a3Tl6IbS7gg8MOH7/qZ29+2Vd
/wqTy8W/SZtRW4/kXDlu1ptX32mPNydBg+VSPWxt3tnJ0utUXfed5bbwcdlD2U81
/CVefuHnnUvZNE8KpWAOFG3dSqWzAZJCsmcb5fRNq8dpEFORnuNdcWE+/6WoF4+6
Xqz3RwG8/xy4VSV5pWCVPqldLlyiSrZ38JUWQUFS/9Zgt3rlXP7KRS59PNCDuvu+
0WBlmF4u+bocYwt+tUQ3adtw+bmxhYEhlPIn2MXoyTDbZKTGfvwJ4L+Dllqh4gBp
Dw8TZn2uA/WXGuCHgktZvSkAvrq2E3K1PUx1uS/auL6LhIB2Gv9S15yT/6ShGl6J
2Z6qMPnovpmjDJP4PjFi5L7t7E1IiFcpsQTxCjApacl0QYByK2a9/G5LA94GaUng
1DPJfD1M0gNyJg+76GQtRPj5oMjqZHiph1SqJwUG5E82qhgVlb7Nf6DQNHdQmaii
beZcoI01La9ErMinISQDla1mgGtkAGv0G62e1hDxjzuPsVv77c4gmwuk5Tr7u3HX
obmWDBL+UgOyYhOPg7f02iuZqiPctezkAgCR4iYMGxb4VF23//cTDEHKjUkE+vY6
gjAlludjT7uQ8KpPUkeURwREmctOmlX73f5IAfD2ujONoEkfAV7TzcS1pA01cinK
7Jl+yTNjoza9DVJ1mdCPRclyDFn9GCYxqhx8Opwde4Qu7T/lpRb1hTbSLk6mUxdY
GXyvsoEsDtB7QOjm8WFwYGVjtyZvLGyJX904KtlGB1D4r5/viwvfAklJ+GGoKYA+
W3Z1rFp2QRRRw6fv1pMPbH2mR/mzbIVFt9mnYlvJed0MWF+reOPOTUHHSe/cpxEl
pT5/GWqCTTuoD7kI+irl818IUEwizGk0BSJJW44/K3CSPF0nda9TTFTsaDluNkcz
LalU9tfuOA5Djwy5YX3Qw/DsAbhke7tnww+aXu6ZxUPN54d0c3NX5WOZK5vqQRA0
6YFR58RTq4Cyz3hBjLrD37ajzYd5wy/6oIeTMrnt4bO5xbdxRyye4aS12wub/PhL
W10ZSnSXQk9dlKYC2sm/FOXWvYVO71YdNWkA59OSqD5kebHvd0JztBLIPdGwaExL
rVio3HAxb9uiXhPofk7ZeRq3NScwl+FLJvochdwuMYppYRFn1JVWoZ00dY21phTU
VR9BlI1+ylMwTEeShPd2GZ0+wcehF/IovUjZ7soPKfu77rZhx66KX/+ZyFCWY68I
E6lA7ibDcPH8ZWXV/4X0vTeEGvGLiKvOmi+fSp74k8U31tVqojLdp+aoOyG4i5Tc
JBP1ADT7ZZxlhno59sfKl46+oJ7c2dvq/+7uD2aHZUQYeEbuRvxTb2Afs4DO9J0u
7g+kBYmzPQIOIIMQlOQ7BermwkohDNbZaIiRhWeNDC5g5NlZBTHW1r0DNW3P7NQO
01kkXqnLr54yufwDQVKvNaLTfPYThkBOwJuIjufk8aRxs9fAH1ir6X6ms8bAelEj
DKf7GxXjwwOvGxeCr3ddc8iuC+4nE+EJLzqfBrHAoHMPixDlyWXh2W3foCrDMv19
E616ZDXbzU4m1axwFj/nKukRQV/oLSF9w3S8tPRZ6vyZALMlzUJRztgYywI4C2t+
yB9AwEdCMZUM1971PZA1TguxydP6JQ48aDxtoh9vYKTKWX1dho6HgXeceTZU1t6M
op5hoKwhdJdlubEoaGCUc+LAI0fsfoopv782nBvvsZ+2dt4yV2oX0yvkvQIXVLup
2xeI4/AobYxKn/IGvKN5W9V0ELvf/OThcqlhc08iz0CGOeLY/IadXTBomGfcRMmu
TBwa6IhCHJH6AQwIUJCyb3ZRcL1TOSAtCEcleeKvGfG9gOnWBH/pruQDl8Tulhnl
+1UmLx+05QII0UmMNZZMwwP3nGSaev1sVhwZbjbksPCgHTjTZ1w++RmiciOP6A6M
WYMIcMdpQoE1lsScFbKeQ2Q2YC7HcjuGilHdkaFWNK0D2qiVsq6DNdfa5HKVRzCe
+NUQsAKjbRhrDmUYqkbJ4ApRFMN3x7korKMvx9xlIE2a+FJMokU2ywCVfvfyG8yH
+1swebpo1/Xo7iweopIiCXuEthzbJytH0M5p8GV9Q+zOufjJLAG3lmOa40KiaGwT
VAXGHGLluyVzdrIit6Y/rj4HXhZP7YvXBiBU0XJfuKVi6rSeAeIzDlZfIIC23Frz
MBe/mDuWI9LHkMLoBl4N6vaWFnopWwy3BvIxNs18KLKQer8OKFyRv8D1Jleocnem
xLzqLyGbUch5yhw5cu/5BuVajmyUV1v/AWKR4BbYRVFeSmzBmymgQ5jCifNEsV4M
u2W3iwF4WOId55cz04WdNbYyTEISuUL4FUe4NCAaZEPxteFD7EMrxZMxAnK+374X
oAgqEXlMJ4kts4omLsOzqy9KIeZSv6VvWsVcTOo4jKuodjVxqurfGKa6qYAQjMPk
sOA00dFJwWmCGfkBVEhbo9rcgvOBOqr45loa37yNvfH0umvopwI+cXhybKc2t2lo
y/oJbKYS5zFOVitRD63ORekBPN9jcCsf3pldwaUhO3dxfsQQ26pfMMsN7/3IdTLS
8L9SRW33Ngh1giJyfJgq57ehWYv369uZ3sK/I095s8XsYE0qig6kYGwZo+s8FRTY
c4wHNn/yY7g0JWG42uLJz05dj8sjcBd+0tabU4HnCqdQ0EhdFbnvd0WGGL01YuQt
Yp03lqTDSXyUeSrGvFCEky37Vol5BcOpxWQ2vosvNK+Fmk6CcTp/7ASdk16n5k81
0JM9Ctsg2IYXB6pAOCRpZX5BVkWOZcXzDmWkVVWPQYDEaNAoos9bLjaicWyMi2zm
kDJLcWiyULXSRi+934MQjvoh4OJDsMQrqxqajLPjoObwMAMpHMUDrTFZ7AswnUhZ
8tloeqmBsLTQMW7acPaTvAXNent5gJ38yxD9/FoMKMQZg68tfHV67aGielL9WoXw
MrLer8yI4muyuvKk9CLbJCaUwZUWuufF9UAMfyemx8RiBeB0WjfHa/Zo7TuILkjV
eceok3dwguIJxYeb6iamDTBVMbZmyOYvB7EADsVIpkKRqDr7adFBjx/mnBxv/42R
htx7D3oUaOj0jLyM6ZbEnGWAhcqIwq1ru9ucsHwY9lmtlykAjLEkPmDFN6tPHMer
EovdplnQVG0k2eozuEShQwWCdSmYWxolHwaIcKr5YFmEPWpxFAs0F4hq0h8jjYwA
2b55ugDOgyeymtNQ66FMDf8kRz87R2h/Z5cFW6oDL80uwy2Q2wytvO9xSAOqv2py
NTzTN4h14sb1HHn1n/f3GTsM33zbgAYb/2qFQKtCI5qjw0RUQSJ1A9MxdCH0KAVj
ex6GNfda1zEgqPBiFaJ15cTTZqykU1PjImv+QhpTvtY3J/vjYORoXW3Z/iDXzCq8
86cv/h2jANzfvN+KR1rHeGRMFCltSbbcuzobmLipUUNmHhZD80EeuPcmNwqAd7I9
V+pmcDvzu2l/elu2v/7Y3SwyYdCofbU/pn4t+7r+t1c/+AXer8GvQg1XrnUq+Xl1
Xy0eNHUDWQYO7VenzByh47vgJon3tRVz1dGNuRF9UaUCr5Y7Nv49O8P3LdHBhK2K
V4oajlAoNxwrWzqVpUlERx8fruNtH+zGEmouAiZSp25NuS85GvHMiqwBAkhT6Dfz
jjmF/8R/odC5Wvn67Y8LJS4M6roHhlppGNO/Y2xrJqrtppxiPVgwUkZX21mKwban
gfdcI5NMSAPnSteN8oxgz7aTXu771OEZlSIvf6L63dU8WDHz2e/O/mjssv7Ncixd
ogKW4yTSSNof2gvTX5Z05Tmfdi1bm+U6U3PgxCVvzV+X5Tg5uZG1JCzImHoUAvv2
+7VcqVka1EAn/zEc0It95wF0VdlKRODI10GrXu4475cH3KRzqa+5WztN7O6dh5ua
q9PNOCYOEW2QrmtsszAxqGxELS85GLxMR8kUwNGBybvZseD7ZLv04IznSSjHHKoO
f+cuYqXDDp79trpYWnSCb2t6xgdGXceW+8TzbA9fNmYymTsy4waNG6ZXylQcUAqs
L/mfuMnuU2LCk7ozXFwrFBmQbMyv8ue1vvlopNCdL4wyLMwER+fbhBuTTKQahcXJ
F6BGvA+07DQb/69S87atW7SS/nQ/GlrgVCX1W2IspfQRW7r/DD6lihOYneu540DP
rnbTEpEfc3sZCX6GGRz3jPTwtQK7qaQU4oWG8xRVMJCym4n8hEIermlYCt844rTu
Uzp+AYXetQ0NvR+wZ74+WnkqsD7zmwJntVqeY3aseGaKizzawoDUsf0gXeAtLdpG
b+JjNoIXtHP894ZMMEG5iwhikE/QZma8TPQPt65KWFhHaVMKKgtp4LJhRrs3A/Vw
43Zx/01ArQ0LwE5HAlDSpnIGbg4sz9GE5ywGbUPQN4b+0ePca8/FhKdYfw9W24pR
D67bn0gw+HhQVO/95Axk+9ajzrsm95W2zvT6XTb66RfZGMQXuAp9tCGujfb9u5Mw
7r4AJrsa9Y4fmRJlSDNAEltFXovskxtJzQu7etc52Q9l3DUfjC0hC7Byz87fophK
Mr+Nj2E+ahhb9FJBYpp+R7cGp8BlwvUMLClEkVcHz37oF3f3jI+/su8iO21RO/dl
D4cmM3SzxWV369keK2RtjV/3zDagpR7Ao2VZmdkDhJAFdWtzLs4ZAJTLS3GwfZ5G
NvuMxlGQ4ofp1TZa5HcpedTODlg7d1c/PtpgLjQ/9PKAj7CEsTuxJIVVrlSUpD7l
lMIDcZhIPhLRfh9Hc3UQwkUWMec0v0UVAt22FZCJdFQtAKCx/iXD9LpobFOBpyKl
+OwR2/drBd8GvT13izqvu0OqOJTSRlBBRSdNJlbdmKDPYMpaKKvUXMa/NnAJcNEQ
TGlECa5f6jYOvh4fNrbPbOX5NQXwRXcIk88pXxhVSwpn7Z3ri23ZLzmYdOvVoR1o
P2yuLp18j2ue8+7ItlF5e3hsWV9bCNDRYOWN80CyeBfsyLjoQ9XP2Y/RqyY/d5Kp
7n7ZC3UfY/v+cthL/jQym4fks55K+iYAEhc4Qc9F9vZtNl88i1DiNCXC0tbUmBQ9
OBt3aPYLRjC9nxHyW5RZjMsznrHFmHMTlqKaZZcg1vE+Zva5CnT0Gv5B40UEPP6o
3+S/LBJR5IebEMxSIPp4fStw+KEe5O7J5uuGcG26RTxVpL8HRwuioDKOguV4qAW4
WpY9zsyZzYKJv8xqFDTUEI2aVi0isIRN7Jp0JzcBV9INZQ4pozDM7qYiW5Lr7HD1
Qe1jcfekb3Djm+WyG44f0XkA8tQCOdSY0Bxb93W8aaNRdJB/MN9H2Y2OX2U0/9i9
B7USA4HtosLRHJYG++ziOVoWjFRwPKUZICHPGtwIZ3njcuh0MR6uhxMFA8n3CQ0M
SSIsG/5KwZmbTShSR0PPLzPZMCwYmkjB7DtqZ/UgMkpB/1qbWL7brGbUJmtLR7Er
3T7QZL1cxKPRtjK26UMz7QzMg6RdQ8Yn1JrljayCHXyeNjc0honQRrwj/gY1GIKJ
lRux9bwIEuVN6k9w7qUeM5cCz/I34fVbfY9kNf1Vq+qfMa7cYgP7HeR73oZ149lw
hJ+Hb6fRm04tlHVVK/4a4THlK7kCXzC7bEez7xLenuXcCjiY+QQxNkMCilPbmJgU
qcI+aALCvcnXY6Zx036zmo2fIiU2bvnIgsX0uB+Dcv2D3Ybb+Gq3EdINUV01mllR
LOmin+aI0jr0lnqKzKwMGxDBPSuGjKMNEQr52eYcjgu4Kv5T90fPLQdskxsXtMEZ
QKF0iW7USJNNLC8jD5S/dJQMuhFOWP5wNpIKMSbkSE4RqRfIRWCD01aDtgl9g1lL
G4YKiZLdo94nwxNSEWQ7vc6nwT12M+j04Xo5zhnDoYVvMqqVy4xq/RjeILIMfV70
nwZOvKJfCCtwAewC7ta+kLsUkkMp6ZroLHTP7H3d9rymbylHCpdKyV6BkZzvpJn1
YtmPJ8sPZbOwwo+8w1gmgyPCNzxk3YSZMBGMeFfZj998Ll1zdx0Kh7b66SoJ8WQ/
uZaLL4ErbFfxs7APh48PU9koRbGTfBReNGY0xYytww+oQ0BV3m3+hvdaXBnBfzyi
iQozh6Btla/+c3lklkVz5AnZrf2RaNBX+G4sY7d4+JnUQQsLKrw2nD/ALIRJGSZO
f8n7iBzM++1Gi9ZGChe5GGq4aPB3zGh6uWB+0fZOQcM3F345JCwRXGjI3s5j8hF3
KsUY187jiJAqYtmwXMPqc+UXiZpoSyTlC+XRdxG94H9sDpmDZxdtIDoXXe8i7Um5
i3K8hLTU5yAizQCzxsIU8vAeNaEsPSDJ74cGzJekqLBZ2k73XxiohwtYhwJqoshp
DnODzq3f7pzF99qr73InMyxB5p0SOheldSgY7KFE2C9GK4VQgQm1sjHDkQPzhL3q
DIA8OfHam1J570x9mUtuac3UOVNTsWMYWV836vqEx3CmCVhXN45g9IN8Em44C3Lh
FvMwtoEl9DrniNMEks7CeDcyadOtfiUpy6zBKQ/xP393j93LnI6x+3Dbrv04Qb/d
sRyJh9v4fSUkTJzJslpkkiDhygwlGWsTFEu+Wf3SYsGMxnQWM7K6Kw8xATBC/x0N
Jnepl9dYvzBTN40wl3CRHCZffWuU8q6NJqCMD6oLpsneq8ViYZHbogk/WWnHHfnm
wijlPbQ8mdC50qtPpjYxhRsJWvG9ebisOiWRtPGbamjvx6IbB2Wlb8HcWKJuGdnO
0pehT4wheWAfrxkwG8ine/ys6KLz7wympUUlIi2xddj9cxVUUGVB1P0dUN0UYWz2
3Bz7kUCM9bY2TkYPxzbSwDQxiqORrU/foDLgvEkD4nQtnRVQ/b1B0WpxXr5YyvAz
NDEFOUbAkHCeDpX8JomQzKq17YPqSYG3QSzwkpspdz0nsGlqlQxBEdGhUpQ5Ry6q
tBM8W2Tw7g7u1MmGmtY9O49kt53V1pisppAWomPl87PhjmN8bhRQfxKfJDedZioz
1Qo3s+5Q1gqxgjGAfBci6kN56rmWui2WUqgQ3/+ri2U5Tf9D+aih8EoEZ8P7YL3e
aIXtk/EEhHl2ZQJRBsSsP1OoPO+QTniDP8T4rDf21EMkTTflDFzb4f1J3BhJclfP
OUoP9nH6BWrAwZ+ufbfCPgoqQ3s/95Fq9YCBnhbhbMLZm5dsnJwFdt7dkiTcF0Pr
ruHLHpzp3ctf35C8idCP10oBBql0girRD9R01K8PSqi0q/oEFnAVi6tlbzZZHwZv
QaEMtBocyXoSpyHCLy4NDcJJc63ADNcc8DALfQEoyo+J4w65m6SQ47LCnfvpKpOb
HSLPdwCCVOeJYeUa6fGxT4SZ9YZkmUk37JYimvp7sTVd8pHKPeNNevQdZLQ3a+GX
JKtPYYQGjQEnOcPWNxnYt3/4CbxD06bUBr5dKzs60Ql5gtTjEfY0iBE9WilxBI05
D5PtrwQ2PQeJpQfMtJlf3d3muPo/utEV42I73or0VgsBN8wnuttprAaQAKSCqea1
EW0mIahoTFlGmSU8CkZ5TGQGrjNJqh/Zq/6pmh/pAT8YmPLpth8OdRzW5kgALHyn
rHNp9Rt1+rIvUm++Us1SwDpxWbL/UAjPSD5aPRec+soUGjsIVS60LczEf4LC4uMB
FCb0VYnuKdAi/xNTIA37r4Om9hGY/lkfdZmgy+iN4sqyeQJILaIS4rfsU46+6Zxg
6DCmPSAWHWUKq7qPeg9O+S8dxFLyfpnuBvWwwU4caNNDp/m7ddpa5xPYsY/0Exe6
HemcPVagyqXeVs1/RU4TG+yryz5cZ2lmRuOGXcBjlLYk7EKFzaAL7cEVtR3427ph
Lg3PwjqU14K9DTJD8wppBAFlLEw8axvNi8MCxk172/LagFAKCfJWvwXsXVLlw/0O
diwIev0RaIus/B86UmaG5y+2aXXcCGdBRYm5VRGQ65cvJhw9MBawZ85PmbkGs678
msdvPyb42/bfH0VLLfxcIxBLPeqq8PGQ6N0Ddg2TY+9RGPpUTYqLSa/PEHKLgU+d
X2lAj686QE8vsrHBVi8x41P8X8faxvK8/DaDdp0mZYwKxaKtCTuFtpopNunuzNYl
guTgxUcBV+tBu84XyPNPNAn1BwL4nz1A2sxotmXujnVlQfy7Y920xqpkNBhEnxOz
iGztt8m3vcphS/muTeOnSb0/9R6MRj1YSEJmaigWlTtlQcj0G4ty340SmdNj15sE
pQJvccdUylfJ0JXJ9UZj5OCU+DHjjXnbduZ41/3WZ2T8vQl5W+t33oXs9D2aMMc9
KlAIQVjZQQvqnpbNpUhh+s9s7Il9TKVNNfW1CrzvtXXtYeqPA0ohfh8xrDKPga0F
jrXYjn4dumC1dV/R3p8PFSsHVkS8vmn+XkfQI8u+CI00aKe6NbRLl4BtVPCkpaPp
GntN2XU6I7rQlohb7ruEUgd08+4iJGKMxiD90MQJcxR5uznphsL/31xfsODx1dwa
nYPbCLrqmiJjkyMIj+QM8FV0/QgD0j4M+4omhlH8WYwUmYRliLswcJhk7pRkc+zG
YVNuMeWhcUvOve4X4D+SXbmIOkABUkAQiV7Njs2BY6KtEJKB/VZ6HkbrwC81pTLH
bmMhtCv/jJbB6VYmPlvd8k5+z1SrwxbPRpHKlaSTIZSA1LVcU8xAMsZdg4OYIkhZ
FQBqFAkuNP5MqKCokO3HhfusqpJ/+Dtzne+mx9SBmgeH4uC3z2vqlIjd9V1y2fGR
2kCJOm8sMsX/6KNum/p9VBdVUrw/6cW4+hPowPvd5C9funwIZtqb5VT/a+8DZY5B
RIPFQC6Zfx29LleSaKHMY4ghqyO03zkwQ3eVUoFeni5UxKxtHR2Uo4iQry25hzI8
oINF8lj5KHqTWpbnb49uxqI5JEo6yU2n8g4nwMgbAzta3dtkCjvgPYcu8+FkNKQI
QtLhhTHpyY589o0NnDR5dGnhCc3RU4X1sKUJ6pwQQk7xkm4rVqRWMxW3fH4hPChv
zTfbREw9qjia6sLLyKKnp0nhCw7MIORZ6A0Sba7xeKfplYauL0TVA4u0g7UbwYuh
9gjSgHUB6vbmnTnAOlklmMAxlL9XVKXEI9SxIRHPtXf3VHLRqHA1jcQyn16follV
Oj86ASRGI/EcLTmjJXWJPkOltJ3zoBTs4J/oAwSo3fdzTCn61unSZSj2xeI/ZU4C
usQ1mqDtp3HLyECS2hFiFHOrK7jE3uFUABC7+M+j6mO7Zd9yalPWGMRHxE03VABx
yYTWgFV+U17qGJ1yTdt++Z7VNZADagE+dpstpDAmOL4gQRGIaPzSYbKxkjGiKrV8
CupbeRQcdFcSjX79Uluym+meo5qzXUPozLoQE+kT2vuxnpr8D4uKUjeDdDp4efQJ
6WX0fJsWtIN9/SbdwHKNNDPE03GDFT/LXKOnrHyO8Bx9/oXqk139Da9jc8Vum1DX
BP4P9HvD9cJIjTwI/k0nktJ1DmYGHCyPMq9HwxhVxX9B5PYYNJgiN54+1xn7H6Jw
eKFM4hgCJ20msKnMHnhm3fZfzMVqtLyrANC4TsuEsiCFG7oC4gehF3eD0hoxgHoN
xKS+cBNllBUTuimlia9QJyNSmi7TfnmmvXU3y7LkdwCLptWxwj/hwpTslpSJJzbO
IRwex29eJ1GtaDWxK60fHO+KrOAd3cxI4q9lhinf3VYHkCsYkizyaozGYoIA6mzI
a7/Oto0b1nKUH7JcHzBh7+ADGnitcjnGXeX/E+J+6BV1KD30L2iRPvrDAQGSMXgM
s4IESnp8x8JZAlQ0nIUp9+RAxRE212bSQtupE0YYhjY44v4CFsHQ2fVC9e4ScD+w
dppj58Zj9Vs7HjdP2ZUIxQRNuNV83ajSBZqkwQTXVD/oTSiz1cOFNckvErelF075
TiqXDgMRZTy31IPS/KKxbWMPOef1wQ1fvTNsngONeWEFUUdwq85qI4T2wghY8kPH
hdaWP2dHDlHiC7jul/OYjzdKqfrZmA2j3ND5V00QiVxBErOGxg23EpCOe3p9UuLW
CPEumsaVCTi/N6j4RfIycblA0l9Sq2/lqgaggmmgYTh7UzJjjScGZSXKJNBisyrs
Nmjm24FLmuuc3cZZjlS0qn5istheKPseLjOSdJZlMGjF8L1kAZvIXgi4rU8mzuTG
P5ilC4XjkwTJnxOqQMMb6CwfsbKdk2sEboD6gsXOBsONvTk7oDao4av0vbJ28eU/
DZ+ZkXRVl/ZGwxqJNtqLjPoOT9vza2cBALUmW5OdyM3epseTyRxIYJVfx7js0whv
6aXulOtCtFUcikA7K0zaTXocnZ2e6dLAIu3P0ZoxsnFyhJQQjVd//O7Y3Z1dfZ3D
dmf9L5JHGGvmgBP9cMUxyulDFdplQHtEUZjzrxGG0ztGgbHVUgcyJZP9IB5W18Jt
MfDvDyXCwTbnE3XhRmLJv956hOYAPB9pcdxjIVIwUBCP/A77EVdgsViQfME+ew7q
2ECC16JYL9nL3ja0YZk4uQtTVpcuun4BUI8vY3rTUca8QGrQrE54uKZz1gCA0I2b
hQb/wksp04jVQofF6zBiw/EflG65f/sPCwbEd9jA6ETCLhP+xskRjqEvRFAaL/P7
Hl08mKFADNyD94ypQ7aPY18PLCE/wQJc0vlJNjrn59L1n2aFluhmaHaHAOhhXpGP
o6m1b9qxlw1+cHcbFrzIEpWB12giKNT28ClNox7F25sQtCwDbrltVJSpCbNXQ9VE
eaU+xTDDXGW+4hjlS0869nBEOlmQ6puP2Gj7I3pRhte1v1tNLZEROerhN+/fPuy1
LM7XjbHy0tHqHTTCfENqfJPysu9+nEgs8ICWE3czXq3Wudp/bH6TPVND5Nuz0Zuu
SReHXoSZo49Fl2sfcA2dh/STV9c35CVim9cYG4k/qwdi9MHRWhczdDjxi3fOyUff
YDIAodXA2J9hD1AwV2q6i96jPv3Ti44aURZ8qhZK7HqXUvRMPdFfgpmuCCL2jX+5
x4ed6iAOMlfYva8McyfuuYZJKRLOAh8ZkgnYTzRCbotldZyFVzKb+3eI7b0wGbtp
qjlQvRgwzTahgJWshQAUtuAAw7UHftBC4eLG9Be/E/OHlq95eOZu6qgdy/+dLXpi
zo1N7O5/u5l4xt0r2UITln6cjQ+53C2i6mekzJ09L1RF0FqZFZgVc52vJeUl47tg
aGD/IOXr4iAdD6so0hthrolYsu2MudDLqU4EY5tq0XivJJ257R2mrGEeYCkhpbEb
btzqfIO0NZL/o8WA7ruI/G4EoumUSEY7wCKvnHT1/ytAAudq9HfkI/YZDDidJrii
KjmIPTrEePEZdSmwzOvRv1jDPX8Rf62pcBseJranTo0ik71g+7F8Wqd4JqY2dHTA
tIOUNFLHtIu1G+Qzr2CP8x0/WkECpv9elJGpmgxZIMbQMszwe9Jl75cdMd09GOVZ
mOYC7tBnlt7ncjZesuA8a2ZFDSRA/Fi2Eo/45++RH3DJQ6k37BoQVlpeb+CY4xGL
ZOa/qzYl6MkHOHVEADvlCes+m6FeaOoXttlZgRjaWktGCFHGNPKRehUCkhR4n2dV
amXFy/YFuTR0V0cWVtl97nkgJxWXeTeA2Jg9A2v5YI+2YkqCpuPSc7LT3r7pRWE0
NYosJqJV6K4QRRygW+iEto4nlZTvmLPdXj3ZU3JwBAfKbYDDP/dNU4wzVJhTW4ru
ZH8Jkti8siaVklSGco//TdcsqAiJoT1+cxOBKkYo/GC8HLoJa6lzersMpwP9rZtP
4KGUnRAKC8fw/7VaBaj3DP+LACp6KNcaLTkZKK3hq1Iwou2fQjXyOKjGmKjPEn3N
lIlsbS70qJD6735x+n6B7gwOfeP5+5H+7I4lC3Q7EtMNZf8IHIXFPoLCin0MsdwV
5s0l1QBx5k1oRXLhn4kMBiq+QNxzEWZtToLoeaJRkPNv1uyqVDd9qUi5K+svAnhE
Q14SIqRl6g0mz8GMow5jQip0DrlALs7VxMvPwpsQd6jpDGGZ4uKm8Oy6erCwKTrK
rAQGwQO6ZjCckA9iBN0T7boRRFCIcMPKjlW0RNBzkfoz7HqSFyYOw0W2tn6Ki0sf
obCx27rFqohVzJTMc7NbvsEgUtXmxmxQnEKZL5jriqDPKw/MpUEV31YoKCywj4tv
/+Bo7fHzLm0rCBCs7hqI0ViYgq/md9DHy9Jpc1O8H0vYVEHTHLqNGTfblK+db8vi
biQyAvlj7WJT7qOyNeAF731H64ln37RPdjNscvn7NHaKZH/qOZQf4qrdolrDvne8
TdQ2ubcgNTX0i4dJvbdmN4QigIPjXF6J6xwSaJFEyNHlJ37idtJhBknZLxdTQ/tb
wnBT20P0mYdRxQnCA5GOe1hJlYXLkU0tpX27fXjJpuSEDxWn+EpEbTre3FJpKaKj
WpdNUaoo4dXw85MsaYx8Xo2tKJkkB/C6bYFX1Vjg4JKkWRp2GdYqo2BVmcqsEM07
yXPRlUbQKtIcO3GQ4Fv56dleNbm6NSX7kx/Ae3H5ErzrRmHmLfGWlpzoq6zRTSEL
8Arm35zRHh2wuMKrC4u0Yr0ilsDrAw7PZOs7T1uLD885OxO7Tb4Wyv+HqrkHtIFd
XCBEOVyZYSacARgEDSfFaUosoAr6cfFUTH06VG3AbKiNEOx1cg+vo8Jv0nsq51aT
3RG117L92k14cS+Q4bfAMkuSIK3IknU5uw/SBR5CqyjyruUMVqYDlHaCBWq1r4Zp
PoPCrmpK5i5hPdXMfYRobZFOYSjAi16LPdVOLXbY/eJNclD4AfD6vU5IqmEw7o6e
+iB/chEtQ5UMnrxJFiWPvszqoe7frk78lnVFGPGkO8hWQLoAxRHwzizJ1bk50RQc
TGY85ni+nBYWJ4HCsyzvhRsC8Q1m5RDF1MQFqHZXQ/ppePdkuFw3NbfflKNPIp/I
aIX1EP4GsK80RPe7FlCvRkPvnmRbedNq1uXXYQknHaImzwwepJty0XmPboBUT77M
+16x20iJk7ZsbaOTp0DZX8GAVdl51bUGHNs3IgVESAmekdHH51l/Gw2RYKfmG1WJ
qLK9kzRH/sgiNhif2zvr/1Xf/RF1RG2spRBbREvFrM5QL03Ae66XFoGiQGcd/g4p
qM3Q7uhuP/00TYmgV/NDQ0gwiVnlYkG51O2984XpJUVONKuUE9T9Z3BXTJA1b2a+
uJdm+3JCkfzGr8vT6hCMiPsXzW34d9EZImaYX1jGelAC1kV5sEml6NJ/+0cYqyBh
oL74A5A8gBx8Hd6YPZxxKraDeAWZhqABqDNPFOakQHQ5iS9axGD1QPrzbKWR2fqj
L9/RgPpmUyd6AEfVV3EcGQLlMJwtvN1EQTNi4eD2l63/13jkmZ/5omSlNQNNatm4
Xq7jOeJcaODpNwoYo7B2AbYZ1JFovuedLJ+ZydXknHWDwcUSLipNZB16O34K0Pdr
pjidLcd/NnbVh4iOGhQfeR91XhNcsKcvmmiBmvJG6M4xB0vDOIbjpabzT4gP3EbX
57ot7rBCigVOXc55G3esdEir792xRociGelntxqoUKWKyYbiKul9GDNEwE3u00X4
9uoU8SdbS4OI2iYX1q1mxvOTR9+PnODj2A3vRVP5AnQ9WyRWroPgHpjL5tUoTGY6
abyJnjSQQb3GDrVrbkn8oM2FEpyU8Eo6qypHVhbl5OfjDOkRXK30xCE2WcGiqi95
dUvLlRmrnpsGssCXJQciDynEE1VUP4k3zxUNycUKjJLMQUfNAEyNmfj4A0FrlJ7F
oO0YhMvEYPbbCW60zCkUIauXFXN+niR8upzXiyAkiASbAij8R4MpADKg8eIFpsG4
21wODoZ68aQRstNQzHOTkEvwE5HkP4h/MeCep4SzYQYFuf01gDgjgkHORYpwWcOi
kZCECHyQaB0lAPRoaqZMv/jYHvDo8AODynzYzTRBO2PO8vhOZRIOMLKkEm34UISF
+MAZaBML1uvAYHNiYC1aqMvhDkEW6gVnti0v89HeaTOo20wATnrsw/dTd9w4j8H3
XtwcXnHyqPRBMLcBfWmpMojpqGgQJQwykTaNCgbMn/yVPV6fxi+mrBZE33vuzYFr
lsDQeBEDvws5Hb8ZsSBLELXjD1Dl6WCC2QgH0g8IJ+oiwTdTJOFhVkMMsu+sd1GD
c4y0wf4IfCVPfR4sPMfYvVArbjuXrIn+FMlk8AMh3SP6a3vkHBMvb+10zP/vIWqZ
7381W2mRfLUWxU1LxOqDtVvFeYcCh+TI5CzXRYX9ha/X0CXCuYfeAduNY5XWXZ6i
kCGMJrTzVWpNnTeog/mChRkjkU/lgQG2pv3KLuIfi3cOXW5tMccm+TXU2DtEMvyl
GoUCmb8Z4ejvtrsQPZDNMF+YFC0h3jMkvtfTQGrujlhMQkvRUMvdBtuAKBVqE77r
fEXHKlKrPY5G/HiLbAkOFh87BfD8+Vfd3q/jBUCekqPduBXCQAaTQ41iKmwGodz3
G/pGPAju1HQ8s37d48bYHI+GhoKTKpvOxwrysY9qYezNLnY8pYJAVIIBbvjCJdBg
Kj9o3WHDtkq6Xg0pKuoFGzbWBT1v/mt8RKkW/uPjAL8otV/z/P34E2FtdpGgG84S
H3OpKHsS9bLKrUIDbWzF1lmC2aJt2KMRtFE/GnJmrDhzOY+GYRmCPAQaACdCrF46
hAEb2rZOiNKD9yv1O87V8/4dZQBPKz/zsahQOyg2SQBABHKDJGVogpIaf9YtUq45
txCZgnos6Nl13kVPIfXNAOgDkB/Va/Xh3HN+TJL6QupNJPz8PLavBg5eIOWvqGJ9
EjvnmM2NHr7C8XIUjAYLD/NK+pebf3Nf5eTrgBqrB2fLoYNmpRppEtpLN4HLe2gH
Z6IckuMFtZQpJljK4S9DjMayqHMdSAMNuM1KIg+gPu0YDvau7I0xVYvfXisM5pF7
zIPtgeYuZe9tFeAAEPSNiOMNkC5RRZgMpF3dQERBKzdSGltdhtCOBlupB9lt9i1e
tQFDm1SXpeoI8f0TO39ZZI+zR2ufXsi/CgB+P/pf98736Dfru+EqoOkERD7QgMF0
s9vHePvQO5dMb/guz57PNEMQQi0EhIaxPImDd0UHtyOUanJRNddaC/LBOl48dXHh
vFYjj4usTp5Ra72ZF4GAdg0Ee3gqA1G6xIm+wDGTbTwoARv//5qKeDogkGZpYB05
xwQfxsuUnZtSfFtvNjS8V3UiceEHWbxStgFxIXPvtJUVPLJdI1d9hEn2tQVVCHMm
90fHGNj/7chQ6WFSIvMEKFghZiKti21bjVC7nLrrMiDMyPc+XwK+PZ/7f+MkFbJo
KQVQsFN+TyyJc4vmYWccvP2hI2peHbVyQTQT6WaQMgh45fTofdPjSsaO2KIrVKNH
AuYow9R7iJiFmiucY0pfB3PupO7HIp65LRZtbDNmWeHpmc234H82NGt82CnXBkN/
NcsfwqpVhTRrpUAScx5z2cJmWTK8d22cJ6dCrQFRBQcmKyzR3/wHy/hR/1PvglY0
Ltx+dJzv4Tc4SsTpCUL35rVlqcGotzeEGOyP/ObyTNtYmB5G7wbKYx+5rLbyohI4
3p3//VaEQECwi0nu9B56izMBIwmfzp+2MnQR8dEZ+Ki02u5c+HLaqnycKyU5F9wW
y21LxXW3zAGUuxrDk5iRTrKP+0wZEwyvR1e1htrTrecvyOhmeVW1Ko79hWrXR1ne
8xqVJwbgeiN81G+dGL/b09IysKfilIH1PbHvn9biJXftM3ZXqn/won8kN6dUSIci
7VEbq5OK9cEyUgC2PxqALLET04VfOpTBeU/lW+AFZePBuQv2MzyjjQdADRZSc8Tb
9Psa7mjyMn/xEHbA98R18z1wVk8VsDXFtbZgRJNAIuFFtz3fpL6gYTglEqYTkYkU
KLduxnkg8lzXDFhgnRfr8nAG6F0S4dsgV79CzxjDjG6lTR393RLHq0QQKljIGFkM
5EWufezNAjzFjKgagF7Tg6JN1PJXfUrm8JH4X0hP/UgUhQiSWx64+LslJ4FvEKTZ
SDIKPjbxXVj9iQyj7o7MQBuPrTcn1ZwPAW7M45vKerLAmTTYpyXc2tcXD0XOX5Ps
Hdf835/CVkkTILAakiy+uwElirWVnSoUKLqBj0DI3dv33/RSLtouNO8ax8YzVt+H
rd5VQmMANcPkW1MjkZisN+HvqUU+B3HupK/9T3LQE8iNHDYjK7SHyrYcjTlaoyXc
fed1w2Ob3MTZg+STcgBfzrBqYCc7OXKpmmio6M/Y0Wy1Mvmhuwkqwd9Clw+HL4sX
HNAZh+oE7V/yGxcnQmH6FF7AqLmSvnCTXp/eCl+YE22PTvuEtUUjWOB50ZXMqWgb
UQPODDqY1H+5z2p3pffq7ZKtd3RKfKx9PSHsfk8u7NpFwq2ycYWpvxbvv0wYtaQI
2JrF0PjmzFF29GqS1UpzXIoQIic5wHa7jahQI8fDC3/F88hKP0N8UobK92I0/Mor
Y6mahiz8IxB2pzC2GNzPzbL1WKqe0CpOwTrZ+FQkKNZeZocmfdx/hNWW0UiVxSqT
shMyS0n1iuW/05bkSYAu9uoLhCCnJowmfY1GyZJg55c3eIsOevmPrBd0HAItVRP7
KyZVriYO2hHMgz77EMqzuNFAgg9my5G5tN6y85Tbyw8dQZRtw/m0LyGn2Mk6FUUl
UXNcJDDofBKeFVM0oRMNsM4Ofhh1ZBtW+0KyXy2R8gsQWcMbRasJNcvRcd0POwZC
7lIy3WN7WzRPcvlUxgkfHBjl0O0T1UTg9aKItKVrCC4oGYuTdpimHrULI61XrzGs
O7Pif8NXAmk2DP5Si8O0gNheACriSKFjUHYCy6xeNLxztATmJMRsyLLqLHdRSZJH
hFFDSLgcr5DvCHQ5AbeIb2tAXksVfVzYHBpoAapmbJHhWDIh3rqqh2X9q5yBuYQ4
IxvOOD5sgFiQ96eTWpeqwg55pogvCwn8iOWmeCdqSgU+CYAOEu0aI/CBd0pXs+VZ
cRPHWxDypk8C2lMuZ+su3pQ5o4C3eMjJ4KBfyV9Nqef38k7Q7LEIZo3a3xBxGF3R
eOaIwdJ5o0mCIQgGrDpPmzW2BmMpxkBBuMTPqn+NOJoWDRP9M1ByQtZj5bQlz4qa
+Ed232QndrbtYb0xc6bvXaNX0nbwJ1KHBZO+bFQQzOk95aHnDP8JWZJ13Z06rjhY
psk3IUPE5QuIJpeS1fF3DawfsTarjF2QZC5D5nk0LDRPcLgEK1iTcBfes7UKJBRX
5vguC6b8Ghk9gz4vMfznk2cLBJ6q6+4aOuhJJa2Dsp1RkIuE3encOBbOCsBjUvpk
T+xcS6jIuWx/skdioGnSgutHI4cFIXFdVh38T20j7I6Er6821ba//mVP6KzXqbCT
ZVHmFnQcLt5bHb/fhI6OaFHB1owvkzwoIwqJwpawHtIOZDXPib+iKcEI0pKJLQVn
j7/xRafU6RjCe9o8O7pjbyNd6oeEUFIKz9aw/DBJ+sqeJLSCTeHf4qAvysdw0Trh
MzWZEN4uDCxEtUq2EYWArs6g9p3STYc+zj1G6xlVb3SwynITX5INEK9cQ/iqWa5X
HfDvF0LP/ONMVB6zrCOtpVktPccFfrO9dVA/4smyb1VetdsmFDt4ZcmiGB6pSH6G
0J5LVFAPymqkn66gJYLTwPBtM7fO9ikgEO6qpjEz1RJBYpOJr5ys8PE0oKshKFWO
/760VaCRtGYmEWF0WnArkfbstujpooK/oueD+hlKnPWfhIyu+KZsuBxmc6FGmWI+
uJqGhstcpAk3r4fYFFPhRutZOxSLP2yXyeufMlOl8/UfTLQBj5ExaWFyKXQS/fJB
5/9xiok5lEO/g9aZ4FSjyNLMLJAOJBhYccvWBkgdh2FxHBkPs7lzgLkvo9UO20Ne
P+kHxWi80bYUTZD4IMaUO5w6RDR7Qn2DOyDHUOKCFXsDa9qtjc9AH66Or1iqyEFk
ZBGtfssiXmDb8b7UYhXBdOGiCFLQLBkKg8a0KTffSBMbjfDMhUUL+ooygIBKzx7Q
gRbfx3NTKO5ZJ8Q/doD23vV5nzKWGnK5viWR/JBcQb4IPGb0h++/A5JvAMPttlB8
xVJfKTpGVVJaa9t/to5SB1OCXJMLf9Ps1vvYS9r9jSeehmRE/EYw8ibEUcrCs/Od
ImQjPqw6anIpa+ZA3ukBU06+GqyejZp4Pf8w/j4wvXgoZ+sgGe36pSG4cLElk1HS
jwgXXahhk01zYvqsDOl7w3ygrtfK8OR61/5nKtQ6doyz6di01WbnOaxBLrfuUiDQ
vVdHg1xCB1BzmXlDqRM/zEJa+F5w+fnKNWu/fZaWUHX/GCOI+U0pBsX4LfhUs/6j
P5cE9bhmoZxK1kSSrq8MTVA2GJkP+x7FjMrPAvxsWu72Jr6dgwpe11LWrwglziHQ
d3fW7um2FYtJPpltxA1KUlGPQ2neZoDW7YvUfCzv+lt7Hya1awLel8Uf6/JT6+bV
txGqP9Q8l8i+V8rRQxFF25JJ89Z/JsTOfPNhh43KT8MEZBCKMRmFD+szEFa//1Bk
Zg0BejwvJOL7eVuW+lVlMrK5yWMFhCr5uHzRWO5cbaDkDCcglAtw1yEazfAKoC/U
bE7WjQ9Ok33WfdzvyZOBhbfWzTvoRGvR8YS0JlmM4+gFXeFofroU7aMnz45U16lv
/d+9BkEeJGbZrqDsMr2NNv9Iawq9hMkFXrViR6/tfheArzG9ZZYc3zwYCC0ypnZD
xJQBE9rFz4EnZuln09od4MaeG4c6rTvzTnXyVMRmat9DFRESdAdGSok4FG95OpVR
WkAcIjK/jAhJ7ud3Ys99WFg32DOY3EHdarS9ow5zKvTJPAhPpgrxi0kjrjrBgWIk
GDgPeE877VDYJ7etC9pa7lMUKlKfiZ8prFbbDOM7aJgS8c93YqNyYYRVpr+hcu4G
BDEhuS+2kZt+5H11rWsVDpVeX75Iq1VUy017ndrOQtKDL6aoMI1xZitnK1NXxoUY
J0Jgye7uFgMrT6QpM7SXXHAJddQGC/OmsO6NyCz8lxOhUFQdrDSa4NumuIt9FLy+
fr9a5WqAYD36OwJgWD9UzmVh0VnH6FWJYVyDyOcZMWJs8Pxi0b85RqiFZ013Sikc
PbQB0F65IKiTWpE80lsOSn7+TlBwfsSay+VM5sG7Qon3LfnVYqGNGjIem5WCTgri
ssK2m7nLjsJMAdo1ysPAKiFsga5kDncnGwr0XTobZg+M/3pKODT06vt16U2gTGbi
HUxSka6zNllXRgWxYGYPgnVK4E8NF+GUF7OUUTBe/DHvAevKsFC8da8cKysZJ/Iz
xlQwBdD+XU5eOcO2n78+g1qXT3dKdn7acNdOdMvGL6fJmy9zg1xaReiNbtyRM7zG
wnosVoypXC3X9yJhmxZC2G+Nig+t+VDkc/AG65RBuR+sfufdpG0+MdWdmOpvxfnl
kUQ3cEuVpK9Y8J3yFDZ0qM242Kau8/R91K82491JBzhu2L3LqzlneDm/qPoyNz6P
VmFxjFSdN/NWSKWsaVcklpXNbjKvVuDv0nZFVEeMoR/5VToeVohWSBH7H5FeAk3b
fMt++B25L+V4TqkbXl9bmdfLuZDURT9BjzQdfeI3IOiAXled1ET/nUh6Kfa7JYVW
ItxlgIrUz+2qpc3MRN20JIOiL7kAfzy5Qn/evTLwNkZLDeuEja+BEt8D3YQCD9mM
5uEiYTgYmnyG5YkDQVGzg0JBFCYldtZnK8FgkErnSvMDtmAil2c8BvEF6wNiJG1/
BrAdqX55EUirx6I1Yy/+dip3dtixc5WdTgXdTiYo7ZlRSF/W+bvxI1sFBIrekuWl
JhYPS6aSqLkYntR8YX28W3gDcVX9qm+mG1Btg+0McFmqk0h9QP+Amq70Iy+htcLq
GuxEiRKLOGdDMyXwPbHKJDo530cceCrwN2ZpOxDsA7MLi05iXrN8IWXRwfpHT0SI
EA//8N6g9TNyDv1m1MGq/ZN2iSDDRY8MYaYfFPAtgAFF7slbWR9LjwFBFNFBv70J
jVLo1409S9brOQdQI+IJZD7cgD98e7dABEw9rilFHMrsiUI7BZxGQmB/fs+LuwSw
q7BrdelIG6OiReCffl9GDm9dIFbCOeeTExRUoAdKlEBW2Dbgn1wx1BPjlsFfqIlE
Ee4LrNRwe6P8nHj/C/U5EJBJhCxkxFOeeT6io8x8eZXgiVDyOHdbF0i1WMs4n+Ra
R1z1gtp8uoZKeqQLASQdtiUcU/93qoWS5bTL/e/89lBHbKaFmFLlUV45DzUAoTv4
JZoZWLVMiQYfZ5mON5eEEpws6CO7AL6EpvB/prJJTFFs1EHJ5j+RLKiAVWsIGGeE
oy189i2R4AWjGSP2cN5hH4sapwOdWI64vDb9sGz3Bps+rAUQXFDA3JuLdTmzYX++
lbxdPrS7j4xiHQcOCL6+MKA7ARtA7mv84kwIASLPjm3upLeCdgBAf8jxtWTd5y+b
qaIRCZOJljr/bMHAcbZlSVVeYCd1IH2UQSR0WnpdlL0rfbw9epAllb6zXOj4hav6
vflWqqOwTy41YZ7fydxOik4CI+p6qBxJcnY1x69g/wezQKv4xT4oq4qpZizs69Jh
KMrqR6Y/9/mxWl3adEUpcLlkhdKUvi1XzzRUcxNY6Og=
//pragma protect end_data_block
//pragma protect digest_block
OfxS9pN2ClnDa7/EXOhpEST7Waw=
//pragma protect end_digest_block
//pragma protect end_protected
