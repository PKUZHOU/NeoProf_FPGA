`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
gAnAAytuloywJoyFDQh8wKF9lNMF63R9mKdDNMB5XQq+4+F1cROAQFZPY0Gepktz
Jhj0aTukNX56VQBTGVNBAX29fg2DP0ZSu/uQOXKXiISzoAg8PL8K5YA4rARqwPC+
HwyuzD4sJUquYi4TNcRN8uR81bcmcOnLaqkUepGB84s=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 8576), data_block
1aukxEW8xk6CMawis9Sa4LTbyz1baDa48oqy4ANUfLTJ81WI/9/LPQfoD63+sXqR
jPTqVVdmgScBPF58LEwacvAxYHHtDwxX8gFMD6SNrjwR04zYkMNmtqqWsGpJpBiY
nd6Eulfwuuc3AEE14kVjokOcXfiaAezniFfPSCZ/34FPuObjl4WASPywx3PsALdf
kL6DKxaUDddyZh0W0jx1DSXragpx0g0LMnswObBOGODlImeS3MntKkOBWYFkM+/c
TtN0zGmpl/4+VfiRaodi8/zqhvpz7U02YU/iL0K1QqpiCfIaaXWZGY6eyTMecP3V
fHJzF9KxwiX8qY4/Iu+wkOA47oEkKzxrT2NLAWcoNW0uTzJUjtg4VwtA7ZdAqrp5
MJWW2FiqlcBA+zvjey4E77F88lhmpv8VmcbaS/RSWKWV4klF2C5gADUZr6iFqTQZ
+2Pmf7ey8ukMdu6ti51qOIYHGFca8Khs1JKiPuPQq72x9s4QjFAJZ4Ntmv2+FE9W
jWTNe9vVuCcRJtE6qkQOZEoPSSwkYgkalTBn/CwCFEh0NigSy+md1TDPgyYLMYGy
+GYQFyozTZVJytSL5wJdwrKGw+UfjjJhrpuHalBMB+qzDBZuvS3SkYKQ5XsyYJW3
iVF/+NHqmFs54wngSQgT/syZBTewDsweWa8J+i9KCZ+KWt81yXOoJ4CVkLn8aPsN
uuW8z/3E93HY6Kk5U059OM126G7GRORE9QcyqMM4PI0qk4LPliRSa9sotyJHt8H+
FWtjFQBEA//4/4/28ByfchciUWht3lgWz3LXWa7TsXbE3DO6McftOijmNTqIKjDp
COkODFXhyAUgylgaMaqhhycCboGEOgQYuJpP8YYwMQd2c1XxScLgIBbZyhw565Ky
4NFHK58p9V9Tzffj/xWgCajkZaHk0L5BFrAjRvZ9Uv3eqtFVTY4ZK+g3TAX6dt82
gzwVeEIRkSpT9MqJaL2J6UuLj8EjofXr+EViwNfoMYnvbbYKMxalxSuOBxzIQ4x6
WxhhbIy/ejEj5QO6vQzw1a5jKT1MOlKGhKf9fVL1w9YCQAqVSV+ATc6GfH8BxP0V
V4KOgPu+1uuDvbAkAjGLwfBY1nSvHn3c/xliquOF9QAMHP7LPNqrwNiLyhpUnJPZ
jjdjRb+pxBt03TLUG7ZI5gBnYmjzw6hUDrcTByjgBWuOgARcuWfs28mhRRCENfXd
tc6Zy3+D2q6SbVB+s6FP0b7gyjn/SDYOV7YX3eSMLjLRS8Cvy6Tq92DDw2lQhjQL
K27KDL5fXxcJboEJDsNNan42+Q+DhYFVv4QPMsL+Mr8etdN6Mt0m7+5DfAAn9cHN
V+1AizI32AgbKpqTrJoK9euFCH3G352rGvfFT3Egf1a6LfEYfcf18WsF9//C+wss
e8tsrwTwivINr3VeXrK4a3pMQ6pzaUl/r3J9ND9OVB+9NeiMKDvqXgOZr+oVYPK9
JRJgU3MhB7doQXubtqT/fATXP+Z7dQ3SjL9Jf2eKstGDUZS/ZScSBNjVus4l/UFD
3duA+IUCJs5EgXbXTmC+SIaNfjBnDIy0X8Efhc5f8d6GcrSLgteGto+X1itiNbWv
qjfiKcJA6PXrn1N6ZFbNuKkTkNGaxuwvdNOfSrP6XinCUDM8pwplDQZO3vL+9cWK
lDQbmpa8J32Poap4K/DD7+8C8z8RqOYE+TAwDY/qdXfNrLhib3B/At0P9p/NFAST
xqEubyNKGWC9xU/wHCK47G2Iu20+2nAgXv5yKrTmektUi6/+vS/lPjugP2x4LgSs
Qj8M8MhIunou3tJ5Ql9AS23W32cKy0WYwFqJqOolWllwo6hDSk8Yaa25fAI2Gg0Y
hHEWbFDHg2Nb5yLv+VGq0yqq9VB3b+6Di5Qjxf/zCMizOoOGrYXMfjQaFvlBG5Cg
teXJSzRM/Oipwn85DrQgbATuveHdnsA7QjCPiodzzU40OZ8Z0RHWfUIa/06573U9
8b0TZO3VBtyN+BSXujYFCR8o7XyXm+WGbjd0mAOQdKuILMrVFbCv2lxmAK+FZUaY
FO6+oRaxuvU4dqoFStXezudBecjyn5ov1TYVJFeliZ06LdUb1EndxQsCJv02waob
MQp2WfUfQPHdkiVNUfaqBPHMZ6Jy4tPpoqrhI07Y6M8WCC1G5EFi6Dp/j5CXdFzv
SFjEHqyhS4IWTyMgDzaMIApPxmpV5Mfk5g3NvvJU+DT+7IBtkZMTdEeVKtH/+Wu+
Y9Kzz9irfJI1s2YD7s4qgOItMi37x/TroEfQGIZBmdCYWP8Bckub9aJfFeTE4TJ2
LvSTHLQ5DBSde8OM9QEaZAofllTafAiBodX48BFmUHVuPQj7k9cD4toNWpRRjDpW
gGSq450ruh0fQIK7Q8/41icL1HWjIdtyjCGCUJeb3if0bDC28CgutH8k3564uXag
MBS4ByZNHHy44PhU1em9civLP7t0z0qfvnqvsTxkqT2qJYwvWhUzmAGaUNmo9PNv
s0GBhCAIlVYYpMBRpXMPk8wilzhjsFD12oORSpzDSWolrg1V6t94u4ZmV4DQpDlb
IdSgYInA9HS9iUAMywAxXgvOkiqLTolurMbTwlA/wJDHrEhShXdGF/uSjpnVudvZ
WbHZ9y1Q5m/I9b91OTmszpb1wnIuM9IFKvtYHI8U07TStWpS9TMDiPpvkZkjukJr
m5mQczv+3sFooOQX/8sCPdifeYxG1ee+WQnXyI70fVVRWxJ9Z5Nhafv2O2X2Z8rr
hRsFjBb6xZoo7Y2V2Ktk8Ou4UzG82IikzUuuAoofzbgdzNYISPlmtkoMAqiEN9gL
u0TCo3ip63g12zerVehrodm5P6ZXNPcQdrD3W7LpQVvjCSfCqApr2ubCoiLzk8xr
Ly4XfIW546B9bACAK5w6TvfGBVfyaeqSnHl7BYbWZy3hid3Mnd1sPlqY9R6adUGE
0OGE5VvkUrNdMBPAvyI4zGsJa6323hquxWY/uORtnOOd9ZOhPaN3t+ak5OgGuD2t
Xi0dGMQ4ZByuKeZNNLA1W3qcpNw8vOPTLzs5kKEgYQPEDTLh1AYdEZoQGspTTeSf
wqzj7e61bx/rN9tjlDuw+2kJgAlRmgfu49m2LeKfHHy3vENPvnMO9a+nta43xKIP
y1fs4AJPxxf4+r17BmTV94H7JFY3DJPdM8BmHj4KkgWT0caBP7UAdnApRO3tJ1Qu
OS9KhcX0nhpapouoXhurobdOhzUBPO4FWbDFDUx9vndvaS/NAjy2SGcy8n1+EXo9
gqMR60UEKeSB5o8W5yrRpDlRzKsmHLaGoDAQafJexhCaJu9y4XHDleqQ5MtRLmni
wpROqHQlTHaPVZ3Es9zRTXFzL1dBZ1l0v5xIa/cH3ZvqJGzPpdjJ0MHbnVKFUtqD
CLoQHHvav3OAY0W+gyHixYkxRad+27mKgGDkw68IbbTS4eOv4mfKdCn3p9EPVLXH
dFFWb1dXnVJ7s5cWDfeCogMAs4Sxao2BpMiIlUec4LK1wbmBN7D/mjxTmBX5Cmcf
Ik14PEaIbYXeQfsToF2AUCSClKWBgMbljkpi3d+/g6P819y7AYQDJwN7hnr8Irko
ZKIJ+Yje9yonWXtZdzNw5V+4mJlJ9ATqQU+76HSmMbFF1dRnSz8RjYjAlMZgeagl
yPTU4Bj2VfpAA1dKCZMTsBCe0iAoLndFuEyJf22m6z7N9q5G9Og8xeN8y9D2g9Y1
UBtOIahx7wiz/Xv1s4oTh27KFJU1Y+i+Ex8LUfvSYKn+Gjy3C0escH//F97FHO1+
atQP8K2WdVyt0/jBZBPuucmJul/cnRHmbLhrWSnNkwKVg2U2jPPUN4nE06B4LQoh
ylia9lzZImhlau6JSUgRC+L0MU+ANRwMSbtP7U9V0xxheZF1aw6T7Y5Z3gorfIDo
9qsCTYAcTVLoQjoXWthiTBXLUBk49C+Zwki8FdKHzPwB1NJ6IkppPmRqrKPNU/UG
XDkgjARku69xyMqgrhbkBix8ay17oHjUPtSbLqtgBFgOmuVWD7AOyd/AZSS/hUHZ
4yE66LZdfwGKtYcWYnvbnfmK/Ib+clX5CqA/W2gXnND6v6MwHD+n9XLcUf5Rcg1Q
ma8GoMUsLg04PFv94sRyD9vB5pamqndSy8qLc3DmpyKCx5TqnZCuVB4zP6HRJVLe
z7gO6TgezMqjrNUELfMQKYnynITMHKo15x90jlVpJejrjaIr1P8Q/IIsGVEbvtXU
KjHamR6eIdmQ+wwugvINoB3YrInL3WOpmKcr0YaXWgsHt8XbZoiKKjkPJKFSAb4D
UvLHGRD+vOsyPRAsBognBAXHFgA+IEivX5YbadscitBy6McP5ekR7oQhCCjYQ8Gv
5pqhYTYfOqj6liPm5K/wiuVXIZhtjzCF9+BwbCIC81vXWqy7laMTCeQ4RLt2Ahyg
lMIR62AwKxL31gI2kAHbNSmR+LAxrvT7TqZB/hdbrq0AcyNrZ/NlFM8kstgZOS/A
kAQ/PfKvDpHPJ2BL2EyXrnDH5eE8Gd/z0VUIuk3cwr6x3/8Z+hyFDqUTwqnKx5v+
IZ2oQ0CWXjooH6WtyZ/kxs1J5PI8IkiiZf9IvSe4a6oiO0bKmxkIv8a2qS6Sqtd5
82UIR5dOWrjZ3CFm9iBEFRE7rPWvBr/237Lu7gZkxs1TJzR1zMs44UqYqmZuusZy
beMg8v1aVoGTNnE+ZFNFEqtONEJZPGsrTe25+XeCzThjOvvNanNBK8b1L5eE9pd9
JM6tTQd+nv4AhOGgo5Okz8TILpk6WBh8Wx6jn3Ber492mhf8d3OpEmc+DF998mnq
f0ToT3+/oN+OtGi0ahA1JMebEuC1h3U4WiWmiQ1m0bJGNByro3PaVnzBhfpdedxU
YKvEMkDZSnJkH4ukpzj7tALzL6vQq2U7NqzTX4cupivzFk1f2jHradX9XtjF1F1x
nuzfSgO+MUi9Up+/O2jOvh4XNx9cidsGpEzX5tnYCCoWf4PeUoBGmL52SzBgJTVR
T7dwjeB/7QvOicwy3OM1uERVIOzVvsyIFIqOd7n5i99ltVjHqblWX4Y6Tl7BUoBI
gxgSg8cRFhZdsN6g9p9JufmM2DGqVBabd84u37lAvJ5ThZkfh/XXyyBMTxNH/c3D
XLhHFBKFGYzdb+4RpM2ATri34s4WvJY8vSOLsFgbsP9O+kf3GwLlKBmyq04M9hwO
6U7U3rPVkm4PqpkD+Ki0SMlVJEe1OW5SjFYLUHEgyAIUJCwGN2jKm/0ILqgMWvBz
je3ECvcIIG3EfMB+whzErQvbFLeRsnGPbwB/CkU9n8n97ME3AyaWjcX7Yayw3fwZ
pN207Ne84qwrixd0f3mTxlcuWmryoppnUi1G1p55lQYFdw+HJyBBYUJUnXU0tDhy
mz4sKOxQ1MzgphiWNKqDz3b3YJCKhUxBN6Cnq/vwLK3zIFPP/aHv0kK71CS6QsE4
CFL1Tsl6nhQBMfvX4UejtdsvOaIRx08fRMMqW+vy644JO+hrzwI5KR+t6/3eKVTs
cDZKVfdepvo3ZSFlBQEFOZavqpCuPJT35+P3kEI2cuT9oojUMXqMnc0WnOsMFMp7
x/WggUizYqMwmAvtXuluvtpfEYhIW/ez8FNC3dOf1pBtH/Q2YlBbkHcLvYAukPg/
YwMQWVOOwzyNkmirfVzGsv37P8aSU2iGjuj7B46m3R2TiharsZCaSiLC/Ic5Yiti
784CACKzwgrbrU5/WvA0voROXsXNKVj1lYDFyH1bnXTv+dwpOACfRXiQYiizmQ2L
+hEn5HDZQyjjfWEjB29bPKKsnRjzJUV9SYJpcQL8PnnlqQUThHIdHGbEOCtXMwIv
DKaPdbuzNL0Y3mwwSpHDJOU6HmQoTtN5GDvaiMdcYIeP4fVmqn9SVSXcdspG15UQ
2X8zHwZ/tlopIzkH+X1/r+etKT/7wIXcHNuNgegiq7dBeUPL6oxueZNqiRAim1pt
EcntsZsoLAx4f2e3/nicHiUU1rEb2Yk3ziYjVoEgT6JTlN0EZFtwhWNdQyHBocNn
ZGGntOMDeik2Q1RyPslk1MwgS2+d6AiSdUoxXkj17PpCbEGFxtBTUss7HDHSlKgz
KncU2hy15e8Nng017LoS66jLgbdfNetxyrx82w9Hma4PNe0xhCeaQMRScC+wRPot
4LHTNxdINEpxHNAUN52z9zCjWR+OTws7h5XYTZn/J/+abtff1Hhq5bB6F/AGKkSN
3c+QfGThgdHAKyFAu2Xgd8tW9B147Sm/vr/fPu8OftdJFmnob/2hUAiEAWWOfrGS
Qxp5hlR+ZiqNwa8cHaHjCsw2tE79MpvDqop+iQyvRo2yyf/jpnIfkzfBzAapxh9A
ADC2NFfoRAoGMW0nC4jZJpZbaGSf/x9Ox68bsHm3d4Xnm5oPecF2lDrZfeYDVvn7
L4vsgI/qLpszdCipIhIOOA5srtULlohBgsUqJS970e2CFamMxx/MzDYT1/nO7W5M
qpMJGwZqI2PWqhx34rXj8KldFm460A9JZgW3YFObOD31YeXoEsJPXoM/4YRiWnlN
2zr7webEfOlE25hmhb6kB5t77YqVFc3k+/AnEhjBckxC3CWr2IpNrXVXFnQsgF82
4iB1Uks1JdGzIUzT0dTO8bbyu2T7xfJSQGlpz1QauVq94nQJowNNKqNuzADfUxsV
1ApB9hyukWQmg8LDu/m4m3NH/TqeDO1fyJF2rPe/gpbcnAwPko4kRzLtlff5/Va3
dSLqDULjbqyC0u2OEvZETW6n3nm30OUNCZnEz0t3Uv8x5+a8ek0ib0st3RHuF4N7
7BVb/hlI2zNHQdkKBD6+yADnAsPuiG3FqsrU1iKPpYRN1Qi/poIP+eyVeodmz32f
q7A3DtRorA0Jf2S7URbemoTznfboLvSIUDBSKpmasTkMx1egMHJ9s1kzZTr0aFzm
VAmZHIY7MZvjvFib+biWWCocVo4Tk6FD7dS/OX9hWLf4k0uSn1mDLv5jTr2KAHin
pcIgXoVypeFHldLM9G2kr9DpnS1dZV3SMs88Hv1ersyEbP4zF/nL38tIPhhCFFq2
MQT2IZWqQLB85LqmJAqqb9v4QWYfkKb9KpyQJ4VgzlUHjqgMZ31Mh/l7uzW/8BRj
UvLQV5FAeGJJqqxRB4nt2zGPQOYWMnf4fDQ7j2lf677SLAbu54UokXuVmsUbxvwv
niYMzvLdQ31dGu9JnorD99jrMOuxDmna1NvUuV5Cj4WI2XrQ0g65bd602P78wp1Z
7L/0CaMrpxLqdkr3DRdsFxWy8OapKab+3E0ZP5kDvfAPm5J4992SkiUf6UasSXnL
MZoP/YIcX3k8hoH7C47JARUjyvI4RRNHcPsft04oHOVi5nP2q0AXEH5f7UxEtIJn
PaN2aFCdhoc+dOZuouOmkHkJE+D7X3/bWTFoPl8QqP4yvsDNCll79BM1u+RcAH1Y
z8yY2FAqybolerpka1R2/+B1Pez/GjXmTkbZtdVEFFsNMWAAAh7WMLeBwVPnkqcj
zGoyW94k+qHYAmB1JBlFlwHJI6Z3NNr6w7B3lgnCZ1AIzCbBRdCbvqg6aivvw4cP
BX86Lp63nGJ2itpbXQXSHArfxB6bmNIA2GELpWn9f+6nyqMBptYk+YNxijh/N9dF
MN4rQQf33iO2KhnCkW+Z+TukzGlqVGsNUBH0boGZ+oSitOzNxKSOLL4BTZdlLppE
f1+6ApEVgwbSJ+WUeCgyAM2u5jRC6gjOZvf5lr+rKzzJ5Ors6IMqTTtc47yO+P1Q
eFLhAiLQ5IZa2OFEvFlFBCwcyQjckwtUJfQWVyp9mNLVXDom0PCiEVZvQnUZ7nOT
i33I2m4aQoftv6ZaoGwrDpjx2FlsqxcgYeTBzyihWCtGtTiSQ7eqsfLZACaf0SO8
ohG2ek6UaB2Rr7sNk+ZuWDTc8NduaHOKSWB/2HUiTjHSpM0PGL/GWdPFaKFNCr4H
DzN+xMG5Y0hLZN4H9m0FvWbqoWcgKGV5u7B2iMCk09G/RGxMrZmVcaZGO3/PdtvY
JCbn1g+NiB0iJhXJv6lgZm9PnXH+IkPTApaNSFkVuKO+ppMbk3KAKaHaE/RaAhZ/
yjI7z7CJGdnVQxl34kcYr4g61C3C5zXW85zqXZk/X9nI/ahMince2YeWkpqjsJD7
8/cjdRmSmKg8bw3SVtCkPG73vD2T5aHQ8qQn2oC6OCHyAPHUqrnQxWd/JgxRndrr
JOiwG39zqW9y0ly2dpyLuFCzJGM377jxdq3FwY6bDxtmY2fKPn930AMUhfmIlQMA
Fp57D3awJo+WrRP3C2JZ+Uz6FXDHwXvRUlbSAynjuYdDoqK8FERn9yUF+PJhzwY8
ytvD0Wfvdv/1p0nWPjO0Ky9FOy2n7MIhzMI7Wh2e8s895HcVm628fhTawSw//++d
WNqZ81seb3Q508tED3RvT4YF4s95Imd//Xfq4CvP+8PfpGQz+zSjhs9Lm7YF4bsm
gHz06UEdpP93FCglYqmMSbrEsjWE3XEIaYJ7Fme8jNfet18+zodTsIBe0H+ulVdX
Nos0BuHH96rYShIl1GxXMW2kaPmhW+OOB/Heg1LAuSpX68w+skk3ze6Pw6muwZBA
WHMDkbjIzN1CIt9xrwYOdlwnc0LijqFvoAdMIKfCZvZvKkOEtB1sl9SlS1/T5KvI
G4257QVsFRGTl6nD1SaryYL81xWIZ/pFqpbw293aCtAcoS2nbRBdb2JsNie6x7Cb
Y4gCuVWy4VB5aKX5um6S+bctnmhLFFK/KT1IaNMEFvNhGNDqauVGnleo05qW/Dbc
3Cf2b8fVIdFmZjA2p+qoOPh/E9v9/Zn00AzEGxNv8KrZ8HuoZI8Y+DavhOlLj2im
2WprtsFRrVvw5eeclnmEvuDhZPQNZtLE2hU7JNpzGbfy+W9YQVyAYe2U+1vY7Z+h
+fW22sWVSYjb022ZHrzEDXcv/zZU61yElcPSfMwECmBSysxavY0sAwqKY6murxVm
dF8X1gIS7mT5EOlu6X6qtfgp+HGNxjL3Rq/CAqMNTmyjrsGxsoU9DIqcgmVCeLYt
J777qT8CYa8XTaJsg2YRKgVG4fNJrgHqV8Jq7cZaim1kN6LQBHVK22IiS77tHTxk
i+sG5MIDlla6k+NqhMsoMen8U45QuSW19AopEAWhmLyLi5knVStGCsUaIgQityMS
fanjCqK6ToxPiNxQE6AQISoFB7X2osP3Q/S2Pl2ttzykEUgV6YVe642oW4EqSsNi
qepdoYwbzMEYCB+KFUu4SUHZxEkRvUd+jHlBJH83ZKKWEtgjldv7PUKS5Jvyp/wu
XRvHnUChOtlvQdNwOhBkDh7sot04OKreroyUPZE2394caQRcXZ3MFuFE6OvYGsZ6
k9jjCjlQYw8LFsDmVjr/hu6+SdsIz8IE7nR7rVBQnMJoLAM3wk+kW7asy6y6mTAm
ySIvQ31gtQB1u7NUTJEZb6Dl89JzXaFoNix20xoNGnsjp7Jp82S5Jrj1nuRqqeOg
YL1gTYsf6C8Oe7PUUNRbrY6z02HJswORAbFeeECChd52h4JEARaEEVw5I7hi/eOS
ptyNvV0BBL+FWNzgeZWc1krbBMTtvUWDUEJtoNvJrkv6XBVnr6wLKVJI+/dZPmdT
AlYsiw+tx7WT4Zp5bB82EVCvEltTx+XWO28ZbFojSjshFRzGPKACPKCDv34KWHFQ
GkE79IXDp1E+D/SINaXVqi0ku/S1gXeYRyK0HJ7C4VWL1NUwSHoXPuZtoa1kLj0x
OTkn1ryF7gehJB1r9vHW4GjNfSws9NN+zPRN4pAUBmfq2NKJYRspOHuXyZZ8rOaC
q1xEoMhSmyN2Mi9TPKmXijEY2I1Q66aV8qanP9KsT+35zvAxOoGTizHlI5m6qCEQ
qCqbcAtLZlCxY8Y6lEKDj1hK5F3nSjnj4DKfrOQAp1xsfGEOLZ53SRlvG2gJ00ix
Ml1Ub73LZn+BH9NefBNmZsRLM8GxKfvvsBFHN3BHftfOTIM3wXumu9GP3GpQvZUa
vF7lBTMCc6paOgs3+1Xr3hbmUSK3fJzO0wygpYWC6F6VnNB6S8NV+44aPngkrZKP
AuHcGnQZxmnf6Mf62taztDhkrYF3xIaKnmY46Bz9lkYLXFJdOSF/D2IxlRIbZX1g
76sM2yo2Yv6d6mzQg2X/rc1sxlgYiBPPN1kxQoY3r8KCDmsBiP0QxdWGWP9r7KkW
hK9DU05xeD6RpBZ5x6/RGI2DH/SeOs5rB6BGjuSgUkiJlhPQIl0MHTDvrKKpWwaq
pgKbGd4hnnbaZhmPoy7QrS19FNzcTLlQBzHqfxei9QzhbsXnBt7vLU2649Pl68ny
up9OInXVtm/y510wuhVlrCWhzn+dXgG4K0y9Q/pIIAVLtFNOi7Pr8g03labIXMVZ
38wwhP69mNtwaXgGkDPkA0y2j32LfkkCeJiNT2O7dXgxKBwPnu5VBH3T38/p9YzP
43LrpFjx5lrQssctVFn4lT6Yb+Rm71nmF7VqMG1s2ZlIZJU307O0gH2Hs9gTKf+a
HX7OG1TIL4BqgHeMUhyhams+G0EVFQ/YY+g4GE6HB8vA/3/khxhV4lcPW6IDzwkg
kB7oLEb4QIOWt8ZL1hqgLsQxidN8eKUY9rKUxI8gAhb97asqF41/KN2wZ4BynkGo
hs5WBG2xpkJuKLkusv3bsN/Ak/skMRXfKK++hIDsC9Nv75WturTN6Cqw0AwXSR1E
5mx9JbCRWoFmq6xyf/uozrfWL5g1SsqeODaCEuWnDOLLGSPOYEy+J9egkn7wwMS/
c689kchTwhMhyITEtNVJcKTmEVkm3gcR3EA4Y7gAPgB7uUONyLoZOSQEG2VqZ+vO
gOmfZsr4Aq+RA7JTnEuCp9TNb2gerY8wUzWUWnXukZoJKj3j69gzVcuDCd9+d+Lb
6/20JnGddBim0hSZKHDnQ7UT7hbkyMjNQV/iimPXzh/PVmXbXoMrT9p3oLMjiV2Q
QXlM6ax6Lwl2Z6UTmH7AP2e5BMS1V3B1r1TBGEzX5DCtyQfrwP/0ZjX13FO39x1U
hE2RwPDLGAr3s4fhQdu1v81Tw07DUvqB5ibLjRpYDeF5Uv6T6TanlUDJqeNnlROE
AV5D3iEK3UugPvVE5mwBTQMMjPyIecpuGjx+Kl90Vv6lpaZVaMzZRwXSadJB6Zwq
lAXqcImldde0RtfAb74jWbdffzptVtAhws2yvKolJMaM8jhxP8yXFv56ACgtoX77
Luhnlv+QfSfPTsogmC2z1YSdvqXEP5gtELvWLhvn7I7izQH3hxXEWX1eLMyoI/0Z
I+eSqyEpUtElkLGvlaNNJ3T+8WZHokveRYQT9zZxHQpmMcBPKjYIjtUQdd1c0ckv
S57fL3hmaCmF1xtUMLaPS3Cn1cAQLPeQxCT9jUrFC3BF9AzcL1UTnWad0KejTOJ0
HLJ4qLyxkfeiTzBZxo5egwr+mt6ac6aQ8PI9QYSCYnU=
`pragma protect end_protected
