// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
qnvKrxCJBfe8jrcZoI0q3z1MsDdDQ9JhpPzprIUfA7F39mJmXNhat7u+XKPIBXCr
e4C8Q6zPVNRra/w6Y5xmFhVs4jNvYFUh4n13Td2Ox3bBEcmhwBSDr1lQFbxTW0H/
q8mUZwL6WB48WmXEpiXeQY9CaKS729iKEsby4Lcr4nw=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 1520 )
`pragma protect data_block
+h1r36oQyIYiH7w0IjV8+IiZHpYwbPcCeOA9e9DsCVXdcG4dUvCibK5V83tvYRpF
rh27NI5AvhuTTc9GE+d12pZs+N7Gx6iV5Vcadw/cbaD3ZcBef5Fd0Wn2/xr2bPaX
hR4Um4WN9lOkgzw6Aa7vx9GAa8R3/IFvj2KNqQHvrbvS29P2ti2cJV2yICPYZEWE
hk6YIiBlxG7Ftlw7uzV4PUISb8Xfq2IbuPwq6r4cZ1ALtXKMWMxLSkSg+fU4ma+L
DcclKBsl2I00UOYDKKRKE/8OAnxfrymDkRPWk3YFgAonSGJB/KTLmnK2loA8GvE9
L8aaTLLzS/9k1saXw4zq2yG5iBEge6NWO692e6ZSI08VgNlETaKXCYxksrqDIoPv
djhZf/IrynzhrEbAW6xBPePWXalHeErGGu9q5Mwhh5JRA0SAm6C5bSk1U/DDml8K
6C9tm18jHJjN+B2qlV9aiTynbHoGrmUi7zFYY08VjzIFy4LZEl+UpSuA8KMpq2WU
m3gaWMWMcPJzu20SCXa0qq94kgBJi3oLrZjL5QXpY7GGhxlRyDJv67BYMzPLYbP0
GCsWNLPXFt+JFFmoxejh5j53OEBccPdwE7QS/jSVMQUWs+uniif2Gt/VyOd1nSzD
W/5mhaOXzCN+RO4NujSRGV378xMtV6XgV2+ZeXzrsGvGU3WzxjssLeU3cOfu6tmK
CJr3jlIsJqXm0kiUv8vj8Adlogw2hVAKo+e7PVDI3THduBvxFy2H4cIoWoTA3qVm
PCl3RtWTQlb+Q6YK9UEvFYOC/SIGsLht87FhmEgahO+LMwTVGhhOEhm5uvI3tjKB
mo5ANZ5zwyV7fa/lymxCgjCbAtt2GCagHqtwlwGd18j9IYp5siURRmeYpCyT2xo+
QXyWr5weXxOUXgxfZheET+6cc8I1rLO3oFO+m0lMEypcZe75ziRWA6ltDT+TQlS1
aYu+nQpVpEK7UANgDjGwkbVlRWIsbFndNV7FhMBmHR/H/rhjleCCBG5zDCTRT18I
kjYr6L/FSdLKsN6SLQiQhA07neR87lUco2s8rCoceMqCTTs3Sb06LhXkiyKPgSXZ
9iCqk4sgBm4A/sm7zFv2n5AacIMbIqSodha4d10Bn3ec/36WS2C4ofwMCFr1sJOq
/IOjrYPVxK/TWPjSgeAMmZoUpwX/Df6APQJC1T8lQOLVhtP9m7xcufsXldyRFpgR
fXnQIC6ZTYmc6PDbx7ID4RlK4ErCMRiVnbPCGF4M04HkTJPvDP/uuRVUKE2rBP+8
oZplYf5S18Lvuhw5zPFBYxlMhspfJk3Zb97ifvYLb35LLvmMzxnZvWdgLATJSurP
FLeAtKAbLqJArsmr1PYJY5N17UdFj0tDfxMHTon07lPvZ17/busopbrjFgVRdsJn
KND6eaR0FJOrmwwD4b9ye/uxcTtzZrHvDiSpO4Uli2tyQAlMrmZZThoxjYKK3GZd
TKgPUcmn217LGpOHD6qhz8jL1OnTfpzD0I9vCyiQFXVxL0VEP8avpVvw0LMn1mCS
6vzf0lLN99tB4y62yWts4+XiCxY9tuDNpy2/7JT0N0rcA9HJMOcOllpcxSq1jPU2
q6qMVnvuYk4cgMLmAN4fcZQVNeRrklvc/Oi/0jzewW4Vy2Xm3MwHuoYbgwcTpBj1
vayp7+8XWDB2h8eltJzYmshImXHMZBXZnSFJ/SmxemGeFLbg9FizeKWm2WBZy6Vx
3oNJkvB552QY+OucsRJHa3N4wpAiSMFQfaRrv9zGJ/JLHruv4QQrOGFB5Q5Xb2kc
rpY+NlfukSCwRxzy9JiG0JnmT81MQ9Sn7iT/ABShJ70/9qZmpA89PHjHpzn4Qi8S
0UOkzHnLEeBsv3OPGmVsynqEKdVGLO6l3QSd/C0ay7j9mtcWtUMOUwucXu+QbUs4
y5GOwplzX73Y7VjyTwEocXfwuLtTOr6CH1xbzuGlb6ydY6pIuHRG2wPoMDraRviM
6YyHDZvG4Pd9kAHJAOUPp0+3MHEaMLscf0k0cFa3cus=

`pragma protect end_protected
