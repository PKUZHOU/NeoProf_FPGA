// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
1rULuUEh0CqsrXADN+j41t+zbV+zthdtUTeSFSP2kZ/LIfTAAC6aUeMyTt5H9Mle
DR5PvnfOzR9AnKFOSZoR26rJOFXN+nKf59L0jAD73VBiRWlALCYhnyneJDfVaOQS
LAUy0BAjOIIoXq34MoWC7hhxi32C0gECahiAgsO1WxE=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 10000 )
`pragma protect data_block
bGJDldglpeIKY5qhAITmwZw8ZB1oQcLtmeGONIaz2JL7nlJycJAVjCYeo0+/uLO1
6JHxC5P8+6MhP1byyU1coIpsZRkjXhHXZqX9F/+v7kvFBwTkX5nUBCGtQinSsEFg
wS+dGfowBXc5cr/4PY9FyBbuf2B/Vo/haHViOBjQpAHQL+XdYOCCd3PacXiX1RwK
JmfE4Q0XCe+n/TCjqVNZXGc2gYJUNvOPRcRQBRKYlO0gf+CA/cEUdYrtkH1T2vaq
Tv9I0xZSy/U/XT+ke1axqujyBtK5KW/dIQOEflX7IMsEFr1I7SF6Q4WQ+caMMuMg
u7o3Q79qZG2nT2Aa5TU5VDOLjR+zNPv8COxBOzbkXktuW1yhFBYmrm5zAVuxdJnV
OZqQQQVKylseainyLQ9V6JJTio+NI4qk2XdkQAjQCwZgwlEkbHRHKTp00oK6v1yG
elcN+sjGAOVjRuVUYzwiPBsMy4Lvc5IgTPsxx2FIVrZUtj2Io7aCy6s8l42xg2LS
yPdnPi7oLh8HF1oqd8VwE2Y5MP9P7yUWGzWL5aFSjrPDC30kF/yX+Jwh5HLIH1qT
sQpuWlpNSdMA6AeaEYd/NcYrTBuCApQio1ljp+U25n1coGcy5BDZY7caFLCiyYMv
mThYMQgjlzgm6Y1VrHf1ZH4c+r+aBEV2zn5AoIquNqSQSAwbmXQFIx+lNF5vet2c
4eXta1U5C9r3Cb12ZlLt1RiunrBEoqS37ZkOFVg9mz3sHki5v+HLz0bzrrCxKDb+
UrhNUzvGTUip4/6Jr0LA1486ymJqUYAb17hMCvRLpEV4zyN7GbqPSs9DPRLSNOBX
QdFIECPXINodxhKVlJ4Zvtz2PmPCtS8Sj1TGw1PqB38JkyAdvhAqnkcUsYSZY44d
boNlFpjscOtdHA98/YCvDGPlksOnZ0SvHId/hFvj1A0IeXptpQIu8DFrD5HXi2tp
9+2DrEMijBSd7V5AXX2+jUxqgouCj/bIJRfY3rXWczT2/06eSZRDOBsUc2KPJsuw
3JOep7m2HhHLEZXS2VPHVjpA4n6as/1VKxhOqkxiSVex2FXbbG3bYsLF7NOfdMOm
ohUL1ER+UQNVqhoIs/VdKpFUdTDIdYhiOWxcsr9XAuvp4thiPWSH3ryrMjq45A9C
tQll70a8cpJrlh8Gv+5ELQVYMc8iCo4+q4V4m8KaGGAm4Gt5x6D9WFoewxv1jgIg
FD5sQvAen8IfmkW0oMsXyYx/3yZu3uAvwRtdqXALpXkP6+aD7GeeWjxOVGDQlvdd
rt1HF3CwcAweagLlbIXy+tYuvlG0lFe322XZtr5FEo4GpcGZiCoEF4iKrPT6d4gf
RaWVh9TAhK3BDHQT2HnRbApuxjggIuo8b4xKsZMHsbXC9UxEQNNl5gorerIEguOC
hQStOKY+wMyML0tGr1AEfpS3fOtR9xyV4MyVCavt+YvdLmzaCo2Ig6MPamr5UBml
YHg1riaeKga5zKP3om6aG1XoxJ6kmU2vQEuvx7og25tEQcb+08HZHyPIcl/JASy3
v7o4pfBmu+Vz2lyvYHYZxigDOyIYPiAJ25pqGKYL74nT+o+KTZGMSZs1Oxet60t6
/RsEZ6eHueEc5hrjhXNRoBjT/t4T+6aUCwkKKf5NPJKM6O9bGRSJTcbEa4pMOSML
kdkFUoXyCv1wicqstqphyd8pV+tgw9nX61WWajE4Q/5d7IBXkzJ7dKp/MGFCR1o9
E6yQKpDusBE4PvAnxG24lOeok7W2suWGvHb9itHv1PVj4USG7UgBWydsve5th5I6
P5v/eA6h1ityvasKgMEoOhgsQ9bl9YaZ3Xlz/qgS33dIM0a8bZdegsjOtKOA8D2p
xT0VM9mVJbsYILLLBh3T6bUwrtsi2RiKf2OY2gjnBMQEo4l4Gnou5CWflEQ4W+2x
QpG2D/1O2XYM2u9apGq3I4AG+zhkWNXrkF7rgU9yIOHsvTR8lMV/4MA/4bSq8wcm
YEskcVSJvzLwvb+LLt73W3wTjNiqzSlbHvNbQG2x8jXtnSvFBvAaI3mVnHdQ+WeA
xHExpta7yT7ptBWaPXUAfImYjvcllLhwosJHJ++UXSOA9MLTauUjFDRU6v/53eYn
dPAFyFGMmPVLylJTw3PKashIXJxflQVoCcK/HGnEyoylYGcY2TlZtDzdK3M5Sx5H
mcQAGOq3NKHw5Kh5omDEuZaPrLSTIAohR/iMSQmyaahSJPBm/1bdx0hJDb+paF+z
zCdoOkFHtZdwffGdtChOb+JsCLERm8478+DbLknn4y6yUerK1vET3pQPmpxZMQMV
aHopr+MV3E02AHmpp6XNn/7jaE5XuaILLJTPwZnserDf+cFnVajnApQx9Oq6kdHU
WMyyNTSUwx4KI25Su+6G13RH/VvaHEIyPU11H/zXWiAsRAB6J7rBJ4B9DHTBmHqm
exf02MIQzarckS/T2hMvh4i4x2KIDnKp5GfsqcRNdop6i6Dj+On6Hd4gMgx2Loyp
QdRnxF8KQMWUgyi0yDQzuYabDZ9pzCT+Ibd4JHkma3WY96mYS5jlMlrCBbvhqjPv
Cjzc/uJGTz+nFnnBQ3FGR5LQFp9p5V1oDZUSPq22m2cHdp27ZA/OIrl7W2k8aa9s
dHjUAt6Bb3j3jWHFcu3bjhYj0Y3Wo6yPRKm3QRHpy6iU7Xa23MqRs9FjqjLhDVeI
306aTmzZCxqsQ1RsBFPExu3MrsQq9vmFZsJgMG13vO405mEKhS+IOA6c0FTBsBwG
l2F7g9wKTVFEBBZpWIUerK57jbkCh/JkI6eiV4FzkfDeKocMYkNG6hPFPD3+doHK
kWyfPso9DlW63UcNreHpegmMhCKYd+wRZmO/AIObV52XHOrrOkmDm4HTkYaTytvE
FjhK19+12/kBot0oqeqOzp3r7eR60Ae+aJ5SmSF86QE94qIEvAPhVZ36kZiAtHqk
yGpfhlZiAsrBw4Yr+gJj/royz8Xtq1/3She6VDjQQKS4t0E0JYP31F1J7/ytUY0p
iPWZINSfS4g6mSFZK5Cz9en2G5k89BSf/qDeChW/tZyUK5P2EMWV4lzsS063a0lN
Kq6E/xYjO3Dn24iWgHbwcxoSb9Grf8GKO+sKqLstGXmJUEXOxjSIiiCC+ZorludI
mBUpPyUwLCaD1Vt4lGpmQHP443GJgyQ21SENYwu222jyUEb3GfIGLAMEzlcKCyWz
FEK4Q0brL/eplD+bo868F5xJbpgYyq/kX1Fi+BJd03cL78blDKLu+uPZ9M7nHEWE
AlABVFknYWsndqxjIMY4VonSL+bquRpKLuQ4sHc+q0+D3ayRBty0G/wTzGSt+JYl
cHFZ4jo86MG4LPUlS8CDzROdEQwl63FbvcTJsL0XYH7u81bFPbd6D6IVdoNImcaM
h9Lk4kPeRRvZzyniJ85E8tcHY6hi7IDc2e1zmI4BYeiozwm56bsBQX3b1LQ9s0rV
gYB9QZXkKGCDWZ9L4LagtzChRpe7gz9DFVn3p2wqowQa82rtTI3I8deBONmvgOm5
udT+xhz5VValpkpo8xdnpnAvJ9nQIfeSP2Rzypon3wfMQQV9h2S0I7uOSm5pmIez
JlVELrpv2ayMgxbPeZxy1tP+UY0NmgFxpFjmPy3aT1k/zuyAj7rgzUhHhdMoOLE8
twaH7TNq13axgQYxkndB4EvqqRjqu/IfmogRi4yU0u97TDQ0Tq1W2W1qCqjUzSXs
OhfiLh1l3TzUwnK6+rHHIRSZOR/RCy+9/Q4t6QxWAUI8Jjnf4J8VRgvqD7wG2h2D
4e6KI7ax9qDrVGGI+YMQyCkcLTMszlEbeo2RjZLUoJyD79V8lOljBe0EjgC7l1N8
wftuFQ+0WpGU9LYIUg5WwHqShKpeqtAfvxTgInhtLUkxLJdHHZcfl64dYIeUVfUi
+FbrkC3PN2Ix3i6Rz78yMLHnkpYLXHUmXDGhDNMLwasWycamYTEszJ1bJHzS1j7u
z8bY2mU3tsXqcK2Eu4tQQHhyJpMX3xxtVPkMIcgH/pfUAsgEJdSwa30seUnSRC5S
RFb+fu+lLHP8sXfIykomgnUOnbCX2pibwOrWUTQV3CEqjPWPWRB4AQOu2Fm1t4Sr
sqqB73sLPmryR3MAOZNXkLWkDhS93RZoZNC8+c/EL9+r1RI31wK3a2e/eyeCrdKG
kkPAUQENuePZCzO3wV/VeX/BPgjo1o+E4DbjeGqJFtf/Bt6Sawt1w6bMhfuBMOwn
aiayH7Nu3loJIrakYhsgq9cOqNDihUgxochRU8Y7gGOyrpCbyhRG/Ii75C2AZ/ON
ebiQ4Z+V/XvCwkSKPOvMY/Xq0RKEIZANJYCiDnKmZ8lrGz0AfbGBtdgNIBazHG06
DQQ6Kbwl2sN7hEhbmMcgkudZoXxzGpMxNXa6EdUUDY78WiyCzxWU8dvlLVYwtT/z
P66W2U2M6YTjY17sgGLrd4WLoyXVD4x8U3TuGF688mktbirS1WCzujAZz0UGIa9i
mxU8ultntW9IaTiNaQjojgt6IYfV5+JzHiO98/G9yTjuLi5traLwBEt2QUmmjAZb
CvLlVeT5CF3WocU2iax30iI6XL1ccav0xwLeu1I8pSxuWHMiahhlOO85jgvASv+l
cU0P7c63oXlh7akqxR8PMNacUJh1apNznvPyiKRCxcUWow/j+qZ+EZ8txr/0qid8
xGylfPhCBQIH8+mvowbD/pPhAkta+Qb+fIWvZOl96PbD5LlT52fsaqkObHDQlFgH
BDyXZ+Sr+JkzsR8oB2sLgqEBJ7Jyfi+ejHkVj8s6KuzA+WKzcejcizbPT1GYK+4O
b4nU4TFfaIq+9MRpjTyfaJR6DoHGwtjJeRUwTrVWlWN33NoZpmgvAT/IoVXHYk9M
xCtZyRrtUpP48U117sd4DqZkoeWyR2Y6sZtiEpgNY6kA7Vh0iMnOdDgpnooLAT6i
jmYPoH/bMjsOcsQRS5fDEssiTMbAQNQ4oNEWBCqTnpOSk9P57JYbtpZTgb3FIs0r
Q/nYhrRMqMmBJEdiTlmQVoWMpqWXKfZajL4OdxdmFtWAQUAumVk9Vxai2VUoDC3K
2+GMdM3Mz70FcuQ8+rtiAEmQYVO86pe7Ho4HTW97kstjea2AIjZXmAdHJNZRVBBI
l9LJf491kqFAc5vdcWkOHEJSdZeHdLFCORNgHVZAk5ZCwIKtODkbwyxdvX0IytHk
DnyYI6jnl3TWFHytPieu7Bb3+p3YnJlUIghBV9Eyg1WwEPROUwkoVFPejxlrDUz6
E8q9nWek9DGTGoHRqZUq2fnzAPSOxjyaTgXMfLy9JlS1B+kuFQzv+iIMj6Za6wLg
xjca4GBDI4RvlfGYbBqV2z7g/0bwJyzVCTUra/avBzDUXYF7z1xNFRnoMhZJCtgn
GPdGFXW3+iKH/hDmsyN39+LNCQV5tFbjXcwts8oO3WamrPK9OOhEQHzwMQ1DwejB
udsP4PYTqLHvrDmgBMj/WDmuD4VJVPk/Kt94YTvGThnTwZrFSzHM/TyT3pPZEnWx
+/HHHhkpn8fwzoWHYGE5Z5b0edIwNjkxYR6YNDdgVxpa4eFzw1MohYU5sRsocB9L
wGRmRQGPmGWL2oj3oXgwYMkAOB9GOk2p2wq5OnC5CRhGpX9ZdFYFkHaihSclafMJ
FYkw+9ci/1g2Wdy6HteINupgd3Mr0RrocrUnHcQdg8JNnnC6VyE1usuuTLFO+toF
beu9jwFjKJ+BxR0lgm6AuMLoEapq4yZHmjb07cewrgYOhiqBXXB/pzE4pm3TSIGr
FTlx1o0ReVaIlgSvKgqs9K9O2jFhacC2z3O2D/UKXn2bc/dSOo5EgExm5uT8WYIe
9OmvZKZN9+2oeaGM9mgWd5Y/2eUA7ISsLDGjofrHNOOVvmjsWu1K5Ur8jhx+AX7x
qqwmBCC/ykhkZxYYvmE01/WEpLFJE4nZtvlD64jaugeW1ADCMvGJpngHhwsxWIFg
dtepQ2g4GgwEBGXEY4MrbfD06BbvgYOfnnAQ8mkJH3QfpL5WS08zHCygEbSIxIt9
sSCYWCg3RNy3mKluAB0T6wa2KWIml2RTHhDDu3b8KvX2C2qWDgC5J5fSH+opcd5w
apHHM60j7zyfDKZ33huS4pdGCqSp+xCd5voZmqvu7NAgE3WIC5RXo1JCZ/UrP1cW
6rmr3a9kkqgx8gRcgPszvLPw8K4fqjMjz7RwpfmYXH8bThHqXZRgwAhppCfdoJJW
VftW4ULw3PRABBiBSV6GWLvPTw3OylBCHkqTJ9p55oXS1nQvyV7VCmbmB8bzYnY+
LMw5fjmrC+zSAD6fuo4wUpHv1wEaTY05sozIlQOxcJuFmGPhzv3IHhXqBwdDyEAb
Z9U9l0mhxSunVLxz+LBoZBHVhLXZNTHCmKWVOTHpL3KPPeDV3tifmeb4JU/lACtq
Vg00nREdoY4o3fFGV53w63JeJdOJ+1AdECmS1NkE5obKYcuERKaw0nAJKiRKHQSE
zNT0us8Pn/YVxG5BhoP3RX9wMgTOMgLphwy2PJJ10qjZrZLSrJG9NMj+R1Wtq5cA
PrbvXdAJfc6ur2b8rTDRV+mQ0gflNxvTTrH970QJPpE4EtFt8PeCtOIkm799SrA8
heJfzkgiqIPtgcjJelZAB4ztj2X7a1pBJAy+/ujTwIV+i5k/TcbqkY2Zgl7fgEGf
xNJv+SunGpw5zQ+fg2QeY90RjvgA8+Sv3HZCj4aISbHYh/HD6SvDIqX9w17gktIT
AMzXQRLFs5Zr1eZre53Fr6rsLJpL/CVai0u+1z3DJQJCWLSzGor1zSgHehv1KeXf
lyXaNbn8OikPvw6nXk3s36gK1CUikBM0uVw74wkz0JUchLeiC4cwvT0g6W4Hgqn1
jaKeDpUTTh4G86p9ugTcUMeb+KIkDAoNFlzww02wDs+7SQbSQXU2QQQVlAQGglDw
YAIjxAHoYDmIenOSkFTUy+d8XQSw/4Fg6AHxGMI3SbgHWj1fYhPwb21LMd/Y4AbL
Ot1j8ckCGK81QphTLgCTl0xCxY5Ndy/CcO8/68rODZ2VIgJkYdJ3SUDNDMuQ/bIe
Hig5UmvukoGze/MeN3bEkZDGS2aX+TpXnXtS+58voR6XdiBDNtx81O+caoymiB/c
k0AGOl93WMN1y48Lf5rlfaR0LCgHb1IC1usbyoo3smRdP805SeVQlqGZ2EryF0Rx
1BXPpeMgUX0Za5w3kqbNoeOb8tng+OUbqNdYP7sBvvuRTDBslXvd/FnUZz3oKTed
Tez6Be78h60hJNkOjCflLdF6qvFuqu5YioIPzDYauZFAvVRTv5ptOA4N4c9805kB
RaVONALdPr9qYWcX/kOOglAaLiMxiMV8xmfS1cqixGJyq+95qI6z0+OXgs+cl5eC
kJ7JVo4dOTNuR/fr6q4GtPiNn9nzkjr7r74S1AlB9c2BkFYgTlIuxvW++TUtB7ve
mbDtYe2UP121+LAlJyOEIjDnCUXMi3UBgWeA++oReX7uuI5XPpKSR5wU2tJYvs/P
tY3EjqD39RUUArMTRPtQji7Z7nS19wTwjHvI1OkNcvNBTKlTv5PvZRUPaKT49O02
9mR2/QJsr5npPzQI0jhjEPLmap7Lx/ZoC9zYChmgNgoMbdseiISmyWawswMUUaVb
7SXVeD+XXP7kdynjZFe5NqvUojDUqf/6P8PeG5HhLPAHWUdnpS8/e8csrQRrZDfc
7Q4xVR5jybwhd+02vVRQfuNnc597iP1HSohI4en8lNmM47wYwxrd+l0vtQajsz8P
zc6p2a3Y0+aFW6Gc+le6qiO7v8vQJX2RHQ+4hhJU1I0/tmq4lZZy6c3jAqyLeMMM
tQ6rswsFaU7CWMVZMPy5layn9bG50S4B6ZPt/QoeVtn2NnP/5xwiBMuvBbbPZcQH
nlqWqZMTusfbP1urT8sz6DtbBzp4A1iJzdDxxTS0IG5GrcIc2RKnsSsMms8W7UvW
jnf0b21reHfTw2vU/zAxvwrw2dO04I+kzheVNtkMpehGqdTlhRJSO21XnoIJo8oN
EdzDl7k2/oY/g2TuC/emDcHKSijcYqFpjqlxAcRb4wXaHLm5tTkN2mINSa1puHaQ
Ckip3D/55qjrOFCMdcVcIf1tCbRDAb/e1/1aYsg7rMYJSXLqtrX/j2bBqkxJyav0
Kv4OdHcp3TxcK6L3Pi7DMgDNlsg1Wu4M/kN7IPCPmkoBDof2Y2IhxVFpp+a1gT/k
qsEI4CG2vn61rJGn7skHumOABt/lNkoUbO8n3ZiD+p7LebA7btM54aknD81vEuAD
D8VVZvmFp2MDqajo1LCYExwNwUjV0tcBoKNCVHNUtDa7nEzVKb1uAVOYfxz/iMGt
wfKyzlYrPd6ObrYylRZqdf02vrY6Ye51HCXZ6E+5USfIP1g1t5XJilDswSa5c0gj
c34JJSGxjD4oyGERrVkTIFWDraYuF+RGu0MwekQfatJUfTGsQSQQuknvTOqvDEco
XE9sOaggIMG4iGOtcGfINZSZgdtthLyOnIzCZ+ScWORC9ytTxHeG/f4cNR6BbUao
6qytkNw6UOauvQ/wDA2bax/gaBkWYsROh7yaNzHkODwMhRJ4AN7cvjsyp5B2HcvW
f055M8qKJfI5eAAyF+42g8PzK+QbtslEjCNze6jS0PL3f13o2GgiJSb7mqrsWkUy
cm96vdLKRtcECHOudakcRxaywffACMNUZGl9rG/WjVryh/bGQ3ChtuArm4EqoTjW
kgnQlH2BAmsalOmOxdTsnxk9AGnyaMLbvdI54mdyl0d3KFHsVkf2T5lTA+cqMjCh
PTs7Qdn2ht/cZvDRlUBOI9pmJaGzbJgvnueTcQZqsoy0PfTyk9eh7GwzZSrwhzOl
ipw/xXGzVXkWPuoUp+HPbpQlIupTAqfsJbyVhcZkK+KnS/kUo3wPWqSacQfo0Nvi
f6TfIfnMWepRNkWScwM5UAiyUXFbaJQEjNO4ydI2jN+VJWXucwNiWn2nTgrl8tAq
8sv/zo8bZz6kpvA8dI9lvzdKEVM/Qm8xf60/uOwIXiYGuGK4QC4ZYbzGYdTGJvhP
Q8ksdsG197CYLHm7SMc8jRXZK4dK8XN2ozf31v6D1AcC2DxM1FHuJ0uGtYrCGGkb
yCVF7jeh1bPl7RwoNfzrixuMF5YGJLHUoXpTOzvfxsl0d7PC3X+Bw+Si+n10MZSY
eHrwm0DygrUvXzOHUnb/KcUwrOj2oeXOnUJgpqNpJtlB6NO4z029+OKgjMz0TUAl
HrF5ndE+0D4KqC71AEDk3BCTJHclEc5hWBLJt9uBs242jyn0Exoxhebc+vrrVs3n
MVrGX9BJa7o7/06v0Ln/Gdvx8DQuOgRnx+q4DtEDJtu7LhSotkG7nGvUuZD3pPEu
ZUCdjVt6Fk4M1xpVQWo6HbPd8n2NveMys/9pb/Dw01xRDRwZg3WkS/sxcP9rGGgi
CTAR19cCJ3mXN3BghVlH26x8hAQnk/rixXoEDBZLTfXVEmmXYc+fsS0iI4uLQ9Md
lMLt2PmM7TioXuy9U4EJcXxnbTs0OiYLyEdXA/xSKNFCIPyGK7Xv0GCfFr7DI1U+
n5klL8T7r7Ndm/Y8qBoC0D974faNiNqLFCKlMGpjsFqocDQhqkl4ZQ8ll5EXzix6
eJhckkbED5D+1bqrhBZrxtZ4YfzCI/x5sacK5mtDCJXbZOwGo86kkQRjvUHsXfn3
sr2iEM7pBFxP9ECsKfZyEsEyk9BrKjtZchSzzWvkVAlo6Ha/rBMlY14sU159pe/x
2OwrxwbmyU2qO4NzlP459jgteGyRSszjrd3xJwzHmxBjw3iVrHFnkv2+tCRppH7F
jDQIjMdH/JLAGNlks27fmqmM/N3YKZC69lir1fegr/2K4i2ixGp6jxf9yr7D3AB2
ad2iWcuw+DvpbuHwvNPURqVCWbbOwATQemMv3qnzIcnd7FebpiSvP73+KwxqF7Nw
+WqThRjAvNiB1PNMAi6cP8C3GEwL5T3wos49U0SzIUwoEoKhcfdytrbJ6USTfmcJ
kC2ZoiG4j1DjpUuvWtgMynfeXNoJbqU0PMYup+4O7H/SWQXfyhuqgtOqw3KeYTog
/I00ypoDYcr3FaD9j0Gvkd7FoAG4PdvlD8nMp9xFwqYxlmgU6xagQxCuQJZT8SSd
Ene8rqskK6nDbJYEDYtpDrCy4PgEVccuTo0CZu+Sc2LMUiux5KN5UEPfum7rSyaw
TsTKk2AUPW0SSxjxaL162xG8noMaMTrqVWprPOJIzNXscIVTCcmWwUGYiB1/+YlR
1NXes/txKJGYQ5Wcg7TlH79CE9rhEAfJZ5WmfjDFMzRQtjGfRPE8pFLOjL7whUB+
sQW+k7hc/qn2v/CR6Z+OTufkq+luFPeBbBKe/2g4EQ19KX1+hjR1Nz4Vu76ERQm3
O3WeevTu8BLAkHnFpDjv7pm7SVpsgVU1xSNgWbYUIpP6tkOI7tilF/f75Zk3BdNP
rGzMVZBLy0P/UL/DqBEge0fR+jk8GRioIwUmUrjK6XQRRL9ciljvfiLR+ZotcNTp
uVrxS6h84v/hv4JLfT1xJ1GdMJE/A+68YYaSqHjIaBbSxGKvqYnlucPljdok+1jc
xYHQSyXZOwGrc2p/NmHbtOkqpACCJH32m3ZenMMMpltmgOzZEY3fYopdEWhwAdNR
85ql3jAjREFNXihdYaxAPZsq1dh3E54uIy0DA3zjOBjBvmP5pJJj1ThzibX1ngD3
Y3Z3LWHPo4vamnSGBDAVPtlNRuvi7j6g14tJxYqj/bUqPfFis3LhaiSX1k2Oz8AW
wmq4Wm9B1T0SZJG8i5CyoAFxVh+/gpZJWmuzwAXt3p43RGZ4DHfjIPBSMeY5402Y
s/IUGqXKxJBkfp81GjzPrj3ZvBvbQHQr7iCGRnqglzrCu9uhmy19dbXpGVQJx+CN
7GMNRUUIK/1dFfrmKLA4GpmMfF11IiGyjesycGvQQgmDIdKqdXgtQpxG/MdQvh1y
xquVJTO8Czt62+V2BG2vV3JVnCo0aaUy0Kdl1yekCwVCVvU38wuj09F85O0cHf7H
B0a9hyEeFpLien34T9Kq0cdURXltvz7lRopNkKY98NFLlyuIgwOf53SkDYLXE2s2
hRiKc0FvJIQ6dwszA7qcwcZPDhQKU8UJNq1F1FprzVYF7INp+96ph/QkPsCeYjLF
EIRabVTaNk/flhawuvVkE6+h0z1u18VdsZ32pxuXjVkjqMVD1ZNpsD1S32sC0rSz
RbJr7ncf0iYdiqUUmZfuToEpvkvJK2qNMkzwlm0PfYui/GSGxDWlcCSpAi87dBin
7iGN0Dso0n1khnHaA3R68AYfb9TIfcq8pyG0xbzD9zvFDoK67aScb6zHuXUF4Cw/
091OlcIJJhEpCwaHQ3bajx2o0eXRfLAQ+hyY1lWUgl2AoSXP/GSznY8Keg18/tO+
7Muig5N/cICIV4JqQ8yyDcu3pnU3WFgfq2yciaMzKXdyV7XW+Xw5KXCEaFJoJN5/
HN2yCBDPxqDnQTmN7vM6MKCf3TqP2nhfr/hQNdgaEXZuk94AhTUvYFzlcHl0EMgV
0b1N62onaoOh/rzy4H8wr8CfXI45JnG7QgbbPABzayV1FRXt9TE2Ht0J0E3GbDnd
STXLUwd9lMJXK0vNmG5FBNV/z+naBBfpVFAb9orDN1F/Vq0Pp66yKZHFKI9gbUQw
MF6+K5BIeKAJVn6I6tau0JJi/IHx1iWQvFyJbczmW3IpZdLpOb7sBv5pdHH6z+fQ
72eODSSGD67iG0f7598BVo0bsx8R+s/A9tA1xyXq97E57AL73z4iWDERKqjtWjse
usZM2XZkUQAdJ3osXUBY9uTQaeZAOdVVWxbc7OK3FGO+oMcZtiEa+U8OLHIYtAE1
HDq6DxIl5FYYYs3NUPZvu1B/z898PCMde7Uaz51ItL7cJYkqr7G+5kLVd6Auitll
Eobr3JEmPwsHLp6pYyMvUl9rxFzLxEHp1UFEy+b1XyhV4YN3vawp0U2n3/RposAi
thZTcXmla/c8flQ5Am7ULz3s0djkAtUKyqROxiOzZUUeIUaYRiI8FGuk18D0PFhr
4+9UZhH2kZc3MWrlMcIIJVIAEx0X4Fj96utcNc89Dyzdjq6XR2sUs1E6WQfHarzj
iDmUegciCtxrNGmaOL62d0Aytg/McTb0lqc+Mq22z3KhkFwRuSH9jfiNuL/HNn5j
sIqkmGJasyEmQ6cH28onKj4E4pAfILZzFIeTTf6+jHgzgyvMawSNfk5d1hqfmzyS
28UoPkyuf3WsfdksCqpJcDiCh+K84nioEXYA8bNQhYU/Dy1VyH+D9Q1d2YqHTNN9
rbsRtYYl76P76z5mKOSEbja9wt1dx3d65Pfhqv8RT4lQmpM8lMfti099Men4yD16
s04EqYj7ltqAr7Tn+6JjX5t4CXxK6/5VGInbSoAHwNO1wy1eIwEmaeoOJj/jojj5
8RyEVzoENzfnSKlhmFz82mIVfky24w6NUsFU1oN0sB4sNj+UYqIaw1W3Bq4dfcP1
7hxK65tg/2mD4CntKKFMSkT2v4zqhiPz+4mjVsOwgAcS/7csrIZNK1LD59J5QgLY
TaIsB4v+rmhbJbnHEQ1D39DsJEuK4/p4luG5Rd810SqDCGrdLiniXp2v1M1AY9XL
q6AB8D4zfvA0oG40haBtlcV+KggEWmBumggs9hqtPAY1/fEhsRdBuKobfMnM8tXE
dRM2/5JExs9xRDDO+QGjtsnFSwXosH8JlS7iN/euEcelnrHqt26V3DRljbU51oFo
woQGszRnWVzxJQ2DLw93c6jkRYYU+DWxA2qSfycXKRJTBubT10wFnHJSuxJU6w3w
89+XJ4eX2/g1xJ251+FoS6THFBBMuMdj/C4/w8plPGyi3VcoF1nUKmIip4tw3pD8
p/NOZ8/bxkMUM6tEEvefZlMYFtVz7NOVHiSrqrXcIRCEdkwUkBwMtRqKZpuIsau7
/GM0QP6SL72fGsETDSXfriI4PPHgU5YmavYExHs2hCPHT6qlzYwbMusqQ59OOMJ5
gqWMw1vUOwizjxFuCLQX7MvZUAODeeJsqgkK5TJJkN2BZXhdu7FRx6TEtW5BIdRN
ffjXj8uPqFkCM4teXX0/Rl1r4C7RMgE0qmWcUvHvmQpmZU25NKge1Srb/85gFtCr
8Dm1ruxnqSsobCU7I3oCVE5F13OWWIvqwSmCFZBv/M9Iq/O5NKmUIV+cvzMkF8XU
k1tdjd1Uy5ky2U9CdhOAjbSIlhZhypv/I7+vwf8K+nAh8bO4pTL4Fus8ya4QNKIY
JYXlrV7xIWRqY9sR/iN2YBv99DfaO6t6UF0a9CBPVaAhjzdCgDo9SE27iuOFJ8x/
m6nwiWPfsTor6jAMQo1Q7Q==

`pragma protect end_protected
