// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
oosMvudzWQ3sLB9QqCcs78ZEjjpH+7sYIZlPjaqtODEOJ1JefcrtB9XXTZCb
4nYIPXzNmqTrfDR1GrN5RyduJ+eQ3wwb+07WT/3l1Q8+7GDje/70kMQsAI2n
tBT91BlpPK5Z2tmcALyY1xN1MCpHScHDZ3n6p+Lo8KOctqjXGwLH8l96aGE1
In6NeEurHFWHSeBvgFxi1WTOeLWTvwU5HpiI+fEShro+7pa1lNWnJ6DdpQTe
XLSZoyftunUfxpIeC5518uk108L1LfSjG4uORRS1oYLGJdKRKvz4xShEgD35
DFxgSncYRkfnYGLr4abatBZ8jaGstPm7LzvX+fNupA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
AZvddnrxPDbLp757eqrgxu9Dic2aIsvEjVaAV1hF/0ZRfUoTDXfVTfP65kMw
mPILI8978+/gVbK0qQ+Yu/JV1BFGIPy/xwhdzgTxSIBI+WZA0wUW+xq3hSFC
NNtROrUkstCZOukqzHjWVYrlibOta6Xs6UbbxNEM5626eXwlDv1JinS97FZc
i1Q9ZNUrVAjshYSdtoEnqTom41swArRZS3ClehqgRyZnKQsy0TT4u6E8TEzb
A5o09hWw3k659V5u2EeT0jc2FxkxrUWLayhJgqyLi4BkFFyNBFGsdto02Nj8
YMHzNa3KEblB80PhTgSnBBKLDcRXEnRwD3UFnAsf3g==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
chBu6OsfbixAHzJ11obrG1NnwjpRd9wzHKj4fkWCWfeDasxvWWIacMxO+PYN
lZvYvoUculFFBrF3hTZoR3q14Hmu/m0UEycm+VVTdNJu934f4jNpUKpMhAJ8
Qh8/zKgrinVZUDbvgVWgecM/vvWwULfar+LD7bEnxAb4xHlibMLFQCcSsN98
8hbX5ctuF/nE5bF0A7WmD6n+w5JK/XRCTQNUOJVH7TJ/yRql2zmn5xvWDKEw
ez8+SN1uuX8G+m/UfQxPDoNAGa35NNxaWf0R1NJSwxtRbEZfH2YFcx8xcVnm
oGC6CMR2/ynbcXhouQoKKVx+nvt7pM6Lj444Rd4pfg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
pB1vSxtonrpOfQLKck1ftnKVj8BNlIMn1gZ/lXujpwk/eXLIJgi1oLCv+bzx
Ulu4c4mHldJ4BJJXFrsGE2G0ubibVm8ATYjsIgv93tenzbiJ6LCy6gnBphKE
skl9bUNdh6Fm+jOFeLw9CK44324U13LeIIy2DgQvfKQOU4NNzCQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
XI+8NuRktM3QeLdH+p2CcA6v1rDNUQOxdH3H/DgMzgvTTitSleODplAzHXvE
uM3y0zxpGBGF5qOqx0GAAecaJJLjKvwb0EIKcZcmIXUw5NdIn1nmhqpJOrtG
9/9/Oyf9aV36BKQkyMXM08TS3+wLP5fLPfTp7BTARjYdyZz/AcyZIPOAjw4w
M69voURFdrSZumXH9NT2Z3KQQX2F7ccTIpJsm2qoGKpBOq5B1ez2y38KV9B0
mmy77XR+BZZlk10qp6pEfOzQ/iGpVn1gOrV51vaOQVqpWt3tkt/7lrDigFYY
J2DWAmTgGMfERO4K5If2GDZryclDwjhSxTHFLu8O1fkAEJ+RRDxNKkto1jbF
xQnQBcKmmITOgxphciGULGc06RukRn+qXob1xfPAgkOtgHo9vsvjXb57ymQd
ew3WGrAkAiRLoYBwyDQwKiJgFLphJdGLTsLm2KzzHtwc09BFbfdoFQkfInBS
bo7SbHX5a4dRIuGDHjukNQy2UCcJdNXG


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
LmcynO1PTCVYFwS/0mkpDSowrpkEp4T/TU7IuEJVvbbK65Zt8Pcui0o4qKli
yPNhMmnXyncI2PCiu4WQoNdSYnF6gwiQ2p7OmHAbGL0h+rOMSfBG4Cxj3k8F
cSWfh6AM4W5I7E1HJsnUw9mkdZkKA2b93YegXuWQMSXsokk+odk=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
tEKBE1Xz71u/i2IACU1Nx4xkc6HC4+X/avqkwmRnubkkbzcYhUWTiwuwppb8
Cg2EZbiesihMiYjDQ4AuVneifc+pOLCm8OfjwTcOpTiL7dhM+u+ILhRow9nT
GxXoaJG56TPb0U4WN5WTIBAEOQWkG8jxsRtiKavtXANTvr90Rxo=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1968)
`pragma protect data_block
6B/42xBdt6p5s6rDCRzomg6LxIHzRgLL4uhnDz/A1lJsLwfwqCzdaIFIBMR1
+Y254RqWEm7YMpX12U9KNGU5o0y2bU9boix0swo3u55UiBplCLIP1W/qUwRJ
kS/n22n8a7xPbH/tELIJxv7ZpSHHQ80dOCxKzB1iWtIm2nI2VTXrzXytDRCc
S+qrc7dZ8ZQ5lVZGKi6vxeKb9M8tUTG1NlSk/hQBxyhI7mLqzspNndtX08H7
LkOdgZZEUufPHrJ/O/nrprTzzBqOHwiUIluuBzdLHBZICUVWncP11B0f/kAw
92AtM6+U7SitjRJuNdZy4Lxrp4Dd4KI7jfioMCjZ4xWQjbfbHllzfxpdqSdF
A0jjjnivbK9z7aBz1ECCtgpqUBT631/nsrm21jLLUHhACfuLHSl3jYEPP7h/
1ZNbCAKP9HT7CpkPyl8/wMU3pPJxQg9O0aCQDITfspJsanW+TCt9lV5jHvQk
i7hLy6Xut25nUDtpBTRY6j7oUem5FPP3SLxLfEoW1Y1NX6u3K7ojAi0Nm4w7
pPKQq6imyVL4Dog4rH5+eWDVIdR3Jdtx73WSwPx094MmhtHiu6te4KFIm5Iq
z3OOuEQndYgTL0COu+5ykZWiRX4656NtNwFAAIElSn/WOs/ywJ2iKhA42GJK
LZFXF1faWDmedpfx444F50Ht2m1YISbzOEI+MQ4bR4XkQu7gdXuwjTPyLwQ5
inFgZun5OZ16oWrQruWmHMuAPp0CKBFoS4DovRqYIduHoJay1LH9AV+kRjVq
B8e8DXlNnIa1y9KbbIa2qMJNXSvlhhF85R07adVut6mqrzsvxPRfEKhbpUg7
jctqYwHhXfBg1x3+HR8O7sOpFE2CNpNFJvrH5RRZ/gig5xtcKYybMiT5mEh1
E3dicAVoiNrpy/I6/y0TlhzQTxXRw8W/JcJO9MYEEbf4IVKTJ6yEsMt3HtXN
TNKoZZKdfIK3HY5ygI+VDe4WY7JzAyh/584l4uqc5nsNX5ydlgCQeALPpi/p
8fxuNsGvVkOzzukng/SaLfOGM90GGHq0IMHjI0g5HRw7ojklmFONIp7ZvxS4
vsIhfhKsTNKmBbD4wiaAiYOKqT/XeCRF1JGmxG9GNKUSHIaROPXq7bt2UoKi
K93huVHLkyiKARvxoH9O+e8SldsWXRfLgQVZVQ949mWLeJ/tHiKpy8nRwT3T
uuZXxL+lKOozrKdcaNzbwIehQ5DSCdzXiDTSl+s6NA6nGEj/LdWzbdgDtBhH
C5SjY+kybPDuvIVY0CwPSUO9P16jTINXwIAJOsegbfAqP7V0/y3LKZpaqlqC
PAfQrw27NANhUz6TufBL2UQ33nWPuTQ8tBYHsQtojwcENJ7Ksd4UPCKsbeg4
lqjzAKeYyWTocKdMiqiZznt4zMrjnJhFzx6O1JKT+GPmLzy39926zoBehFhi
TkcayE5rXpTrWTfAJBW+fDEVYF+XT1ZZhQim+j+2hchRIx80O8oJEvpE3tNs
IHsFr+VXOUnAZWIc1TrUkAWg5zNEGv7YGWqsxszrsmo1nBSZG4ifE3vo2hT2
Qd4adcYWkQDEU13mR+YBul2fzPKfTDlTEefqdw7ia+3djcqoEQLGXgJS6Hqk
Y5LrxQ6DonLXsRn1SKq+KQT9xpxf41jTEb+IzLBNNPSWfM481wfZ7l6kWcfj
lhVas8NYKr1Jnh2o73DxsYRy9N6lwBfh8DHiq8MO6jqLiJOZYFahfdlsNknJ
Tcf7nmskA7Xa1KttVvUNEKUOhB5CObuz9KiPtHZhXfiYX2K+3qI/7j8ReK6Z
MStZeufDbYZqrb/m4zn7ryXOmzCkmWJvnSpKgWr5RR87N70/4GJrVbOTP/7l
oBoEP0tS2q4j/4baNeoHDmtY3Z8VxGB5LIkwwMzIfMdsKEjECLlZ8+91c+jo
Y4IuG/hzKeBTeAnt6RGOQchexCJkTfn40wFB5GcD55dKXp5yH8UpS8/vZNDJ
eyKPNzntPPZbTr5sOjiSYUvCp6/VnWwnRCosRG6hYcVo8TgBLgo9kKSjkeRb
GS+47zXe/YjOMN9AQJefXGTRoXWzit3sSCLes9wIrDL82BbAzlyP0sBqDrB+
RmdRv/wk+rO6prdd2VDPZ2DXskJPXleVr63aw1W64g3bqBpoHxtl2Wh4mOz+
bkGp6SON8Ap0gg2ydYPnbBXujNgEJVPRL0x4a/OXO6vFkPokk/k0prr5yeiD
iTsLzM9/eB5wZDJkcy2qo3LQF0JtWmqpoj2l1XoZvCGZrCmY7QKyjzbKIqTt
L7EnSZjmebomfPxKKxWHY5LHvcQyASnD9tyF0Dwxf62lsaYiYb8/YYIkK7du
8e6EzvG6YeGd6/OoUjpfpgIIOk/PBOykuxYAQuzLhNqyzCO9FnxID4yy8+Vr
Z52I6Ryj0r/ighLwl+QtFgOZ1/QrtHTYHbcpDwqOdE00Z7bw3tlsT25K+UBe
dVx/WVG+ZikYEMhhKDBp4nY411OPD+BIwurDx+9CuTzkn7xgwTbcb22LZELG
SAgRMXQk6A4SF1ebeWYrOCnd3ANM/9fI0uV0t4RagLGr4eWi9Yj3RGEmBINt
o/Uvk8nwuYa8dr/quFJwrymhNLeMdnVzrG3goJ64/YWG

`pragma protect end_protected
