// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Um3nI4gRbk0hjLHCeNRRznAPRDp48UkhfrSp6yudNicnljKpttNMiB57trBG
3CP2YD/5BPgu1WeeObOJMpRGV87NiSFGkM4VrLd1ypSDmX8AoDsbfNbRlzsr
j9bpLs2hbIiHsCjgKzOEIowcpQsCIwfj/krbAUtoI08IcORSiii9VYR0FG8g
UW1m0YwjmAbFJIbrODRxfwgkrS4OXa6EqITWpigBdS2RZg4IteFNOTk7joj9
0NcNdvfC2aNzRoLxxt5rb5OQ8wgkisL4IZr2Hq24oAHB6xvSZSsjTRGQOHXi
Y6JPfaSTkuzt4vbeol+mAv+acxXqTNibJUNDC2OCog==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
GJ9Q/xPDilTiJmUUINKrRmnj9AwADuwDdGNXM04qCgwcIvRIvqKXO7M8bxc5
ZJtzMiK+MJhnmNXbr2beD66tO/ftBmCRERO/1bmgNpAHCOQIVbzKwHewLy8X
lgi4B/eSc1M+tpu/x6WnulPSW7rnHTzUNgaAXYGbpHbhYDttVNGQvevI1Waa
sKfwYyA0EF07bow4zlGBiSOJT55B5rbfikgauVDwhldp59zNlsXVrl0L1hNp
t7mO2d9JtSQAWykZasZxWjwicpwhon97NNdjrKr4TSmEtEcOuqV8TP5oPkQw
dKXrRG2OuCMmTvlyoXWIfXVu0I1oWa2d63fEKZ6bhQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
cGaOXfH1omQ/AvP4fQanFVFEZDyxDK/GxuJUMk5td+qWPH7dgGSPJIponk+a
PLvxdu+e7oHijFcN6qYD12S63W3DUuUVQcfvLeY1fyw59LOqI0DfuCgFXv+p
l9Bjp2GZ5A0QXdhx78Bkr68FR3ZEjqTnQ2t8GR4yZu2QTdu2xWvFpdX+wMaD
dIaHVrAVV/sseO9PMKZY1eakwRuvmYWlZe+P5owaQ6TKjfhSHAvESkZTEnq0
3VYnWpNTRJxi2jjzDYNWcOwF+GlYQND5W4UHZAKLZezdCxvAJC5nWMuVXvHf
6RF5VqqXqyblRDjktfILjhRwIKz47ukKYET5aFM0Sw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ShgGS4isEM/IvTi6PHXdBorwo9uzFs6V1CRzkiM0A6dhZkbnQiQeTNR8egmM
RBu6IpGGcHVbq2RF6mL/lOY/1L8p49DehgSOVKRNlzQM8mUDrWjhsh/WEOU1
Z2RMZOPa/5ji/MmwM2wTjBo/+wEUiXAAbIJP1SCBRUgoRLx20eg=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
YLidw6FBGAlzfAcAKG3hd3/FFfkDiyvnS45jYF1QDZqf2hfo85u63JByNWJ8
ewKJPaFHMELIZKofF6WZBLCcOItWGaBibV9vhtQmJb+6++U0FYsA7SeAePG4
wqDe8eXpGOQ8cQIe0oU0ESwfC/fcgemBdJCEX8XmU8C2PWUtHz94IBmbwimk
jaljN63PKaoUYCuRwv05CwnrO9uQ9dKEqOfWXPeYpJIoLGYyP7Tj3oiyPT6l
ihE3B5TaAX5loFaBTySodmQ8gEOl/OJUvEki70jpVoddPmA9NGzlB+VV0dMB
KL9+imkokJzaNxxiRj2hWFlAPLypb0NlEWJMwwa4mk5Qoqi+gLcxinpewCTD
wzersFUPjkWc2k7k9gCG5fHgxJlpiNBRCL2LH/aXDAvnMBDZXLolBux3zcny
YctZfRto5nG5nmwMMUeIE2g4dpY/5mHZdjTPRYAWAXuIGhnPmMfxoKHT8Gyw
xYUlwkxI96c1X5obqA1REAVUqp8lYmJw


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
GPVJtP0G+OxPztrLmdpB6M6pnm685o2ePYBho2qH+DBrqJQKn++t5UMe4rYM
medAXNmdeS0+76e+sTfxJ2KesSs1wH6esKqRaN/T9BIwd6xRrdEZH6KHHy/X
WuKfTg/Svuj7pzHJwl4XVZOhD9Fy2fsfj0hExhYa8fdSXPSrR70=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ar99FQ2z94594u1l1HF42VoJosqS4Eu/NSsoCrFsOP2WPET44TjXRAoh0+xp
751M1cTfCfY2tZ2+ngS2EQpaoTUyyLrcC2pSpmqMVdb1b7TFMAAA9cUldElO
Q3dBqZABTg3SDfxXjJVen4U6rbFJ+OcL224Xs9Zwc0w+pnAeVCw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 13040)
`pragma protect data_block
AJfXpsRrF4VkX3P/YgrJy5GodZLVdkujqDVsYW9Nn+KiGEkbyHzdZZFCGKdk
0DaTKbE4Vi2wcBuidjxP8iofiawSdrVO65c0WNkApSrgjb842XKkAH+vTkLI
pUSF1aYcyCU6nwa302w2lpjKjIaTjtx5npso1B+cijoHOiuciY5DjgJRkxMI
xWA8lJEbZ+vn0WchF6OIulv99/vF66soWyHMx7wIYTPOnKQilajBLYWIsFLa
XjXM46y4t1yba5hfipOwZIkCez0RIVRWyCWVsL63pW2SqBVfbE/apqEv3Vkw
/1MEs6IdQpfnPD0sEmvaP6yAmLL6uRtDzMgtO33y3kSSMtvXhLzNhAk2sq9y
Xfw4/HL3tFH1Yui4pLKyiB3Z6clJTi8RXQDvkJWV44rEjPhyRLPFpLe+tPSA
MevnpL3AP4SQx+xARxTfJxNEfGU2+auNffxhYLbddg92bvBayRC8pONheWTb
yPnKDrIGrED9apzc7LmvjtD7gYj5yH0MhcTTp8k+USy4OU16l9H2O6oo0KL+
eKd37ArVDakfz1RVrMrIiXCyz+Pqio0lGPvnVZdXoE6yvsKlUDR1OQd5G5TO
5QmtboxR9cLZx3kcI7P8URB+pmwRBdciDJTaMWZQYikxq3PXSgohJawWQzzb
ZIe1eKto6+ReXnsK8Wajg4RO9zSGYx2kLK+LaptWjP5NetgqXs1ex0aXQmak
6hQ/tO9UtmHgBhrLf1bw+2xgdq8mHnF6sY9xEc+a6KPTgKwMqYyPBUvFb9Bb
PqWOGohUdH29IEXMZJsOw0VWzQgaDEf7GHho4opo428XGrfXBoOje49uICcQ
UaygdNvGvYE7DQbKsHX1oIR5QTpIQvc24JODNiiTF7omi18iOLeCSw5X8bj1
R4AlK6A6/4K02UzE/Qk9J5M3EuPwfFsXJG73A5Ea/IoNgyGM1+cZkPX2+S5N
QYfR6wyBQTN6uKDtqXVsqcpo7IAvrZSrpLVMN6lpJbL9WPj9VfVpan5e0/EN
IDw/h08j1cNLgrfyGTjx+q7QrS7hU2rbXMFTEY3YkjEp4STkXNsbLWc4Ym3M
eKnHrd/nHaJgrEK/63uvoMjLfdI7ipOlBgOd/uPqWV4SGBcA5jzQEvPdz1ix
oi+x76i/NE2qJyWy/POnoexcnzRxCLDhf7QNBE9Bq0qlLF0swQuk/7KSOOuh
xF3rkQIB7bZLY4fzcYLqwDE3roodKo9Jesx7kmyBDVePCKZ1cPt5Lrl1qSBs
Wwhe9QSzu8ERPCUOAXLY5c7SPXoeymwecmhGAJ0a0ZUXMDVW1ECpq6eo9sUD
3v0Vmee2joRE1EKb1XbZormeubt+s6PETIz/TxGAuXPjDx9p0TEcQhX5RXYO
FGFYKgZ+zaQ8sCLbYwto4u3knajbfDPMlymmFozq7bASSgzVmSaLsi+Xhlvm
KP0sjvxEz0JZuwXtXS3OFGj55ZI2gSOfqOFB1WPUzKaUh4kD9X18WOSzLoYw
7PJAdwwyEuqkRq2jCyI1Kq2tuVm3FRq9kQOHbqSI8t7vcVKuCK6ofSbwKbau
LVKzRylcr6kZAQhtFd/SBnZYfnjOLezwrfy8Yu+kO1WOuQQIXABoMttLbZEP
OePjJW0kwtol7tG7VIqbpQYKUdS3KNAD406jOPKBY+PM6i7Ll4CKQlGo8u8C
8cl6a1n76j+U8HaIAcEbrNIbpXuto3Jtcs4rBBV1J8TDrDk5QbxLOHKLzH9O
+LMTPOMuG99jHeMzrqelB9DBwQhaL84UkTHaiCEl1IWKn17BtqiN6Chw9vzk
HsIb2fopIKbR0GRkHu/42qKXuB6iwoM4lPMSEncXaYvU8TvASpwUAQJcbMDj
CwXDIoJjAX7th2XEFJvJw+rF809MDP5WszIw9MgPBBJu+5nH04OX5/0ZYnuv
Bj60SOyVB2p5uWLR3WREtkNVMns6ZTDSco2oWudBFIck0C6d+/e6JdyicMXl
4DwwHCwPPg9OErYZNIUCsE/ZEqs7dNle1PqBsp/6Z/CJuVvx1r/rW7TSAg8z
+eOChh9gL/LhxGkO/4HkJbwpyFaX+JWoCqVFgvmvgaIBxiALtvm04/bTQgV+
KTh8riLds0I/yoolWGcwjr5Af7jYj3u+WZtk4JEv8KnsIS22lqP4zpRZbNg9
pWHbpVLCq5l7IRETS+CJBamrJSQD22jSWUQCo2dp09DwPKTi9HjXYP/lFSCc
YhnjgPz1pdKxix5XzIYI+XWNn8D8l8nwxLfCBc1RN8l6wa/KjqQu95PdGHRG
cJY6QND6jHvBozeostJhzsaQYlQcqtCpBpaiLLys3oj7pWwlAHCBStquVRWG
vpAjUgHTJOAm01t3fcsZxNEypSuA6qEFWMxH5oUOHdlZOukdu8AtuhUNkufo
Pv9FZ6F43VF1dnqdwUwzosTfTs0TEI3QG9RuwZYJ/LiduT+WfIvZunDPKMHf
2dfqDHk/bM8jx4P/3qmVApHz6WHaZ6rW1HJOYxdHewBhgxFiKI4uSx/OVFko
jxNxgnRTQgNfl1U7qO2H0Vtf8yyGU3t000p3WynIBchBTtHX3RPGs43V/t/M
r3kuLTrhtGsz63f9ZcMKAOeH6GEmhUZLUqsrYXw92zge+tWmzaH9sGj+/JWP
kJvUY62+U8cc993yBLleFTZzegXjnmcgivB3G+oEAs0ryNN9LAorAQuVqyK2
Fn+YW6c08YcEhezbl9b2iF85lW2jd2HzXdik/InRtlHQadYxKy60ZLYc1bJu
CoTA2L0nqg4ymsU4I5KThbVcdMKDGm+2VO2zjVDaTLUmz7v2rLzIS+xZ3fQF
g9Scu7uLxNn4Hy588YjXyyIGWOJaSZp7amIosMQvW9/dpA6u/zPfEXapRxyZ
tYRATCcP5qBXGItjWdT8uYmSBSCNFBe0zicSiXQVU6LW7i49dM8jdH2RqRv2
4GTVZwNCwbuyeBzVuLoyNbmx1aAJb7O/r+1xqfAVBede/5MwgkaSuakJQBpu
Rv+lEXp47Hf4GyCCsA56aMG9FFrxloeL5OFDECwdv7Afz/qtBiRSuvoVbgyX
t2Xi3A8qb7JNPrCUxcca//n1LCfsZZZcfMp0PkK0XP7b3OBDOsjmKuuXzAdq
WS43XxF8UTyhLmn2APLIAytl38uRIM3O7OMqZlwX2P3kyIPi7SWL9ebJOpVy
8iVbzo2wlDvtfUn09TG2SxsEe5yjNpOYcHyiGnHb7fvFySR2OIzWA4IJ74ke
nclXww2gNBS2uwStaFTnhAxRogd9PAisxA5773A0TkkuILxlwOMM4f8SfkOt
Ei9TiM/yRMv91Cl4mkrWTAoLmpgEOQeg+6Y6iQjY9+6VpGUlcuEQJYaET8ue
dzgG8zY5ioAydSAotiey36raNXOE19mpCNTygSu2RuuGXFPNpuYk5YSAbIVV
rVhs82nOxpq85TicVXTgD3S09JJ+s49iYnw2ywDkcW5Fqw0vrBbtoOhwfiva
5mcN/NF1gaSYScS8fu/rncgEkdDf7WfOtzr0bO3vrkVzAjfmo9R77b8jd2UM
rt4EO2a+1Qpzm4f2vJnb/T4b6tC7KVmo00cYMR4hpqoc387v47tj0jTwHtna
uoyCW4XzHoGDYQtq2Rtq6Sq1gYm7MDt9xU8/pgPoOaR+ZQNj4Ri+H77p2TS6
jqSQyo+z9fJmn5VOL1ELXwF4lIWZqgh+B0ifaiQqhoWxL8cBR7AIK64f+hNP
FckG/IWcbImyRRZ/uPL9+m+hXHpARgsHUnHsRJ9rROcSyz0KJHJiccgk0T2T
UqcExN+iQ/h/VXZfJSm8wkbu1CQk8/Oc3n0FVyjiXjgP0e6kyxe5dZBIHCde
uDhtUJmpP0FDHABCNUOqyuZIpakqs7wnU+kBuieYXXDFJlImbLhI6rFp6eEI
uPIPdFS8npyH/jTd6D1uZQcmXnveY8mVBkZTqb0PU/KWfTX/bZxevN++8dg3
Iwh6CIlENkCeqfJ8yLYsHAxhj/Vazq9PymvSvNSzWxN/7+rI5zTQcQXDn4jh
1XZ1jsg04MlmLJY7IX4ljOMP5Qaj4JVOBIvvKdhm8f/XUNdROTBBXbUmj3I/
F+nWki7u10GsOWqw9O1wexhgQd5hIWEgdeXBCcDUAAlgvE4HF9a4nWMNjm1b
LcKbU83daOxKPeswl7KSyHBtl5leNMlBzwy/XCWEfrX/oZZl8qD3j5FxM1q2
zsBoZYhRzi7MyPcEiUeWma4Ub5tMxKbWIraQZ64bjjQBOShJdvpjHk9LEgGW
+EdrzHeAXONtO3jGEbe7PxZxxvBFFUuTilEz7qvoZxvabjn8KEVwUZt0QU0O
SLxFGvW/3SUTtZPiZxSnsgWfJVXVAONhWQMBTwOiXAjTq47/u0zu3q8UlIGJ
3sNElxjUTVY+UTr6DrMDhClXoRBTZnsOW2GQ8RMjL2ns2++6vfro5UxeCEl8
4y29+JvpY3UpFbc9D8RIToVEN7uAIozoEdjmLJRbM6mJohmrZwA1kjbzl8d4
DNVrYdxs5bJcPA+f3haOSVqjC2q3E4Gw9+u1oH4U9dLC0LXd4+9t0WwawzaJ
Jw8QcvOxzM4+mp8E6yX87s8y85DpBFhiXho2fp9qY/aAQ7KpQq9XbptuPFo8
LPf0ElFotXeX93vjErwSQCfGP+cjtkoKjZZLh3NBsJ4tJnWWNT+/apnRnAaf
2E6IpS8rCDYQzQjGGhfQx70XXJK5vTizvuBopfxGBFhmsrREDpJY9XZKaHuN
hTTXU8ubeKti+2ohVnlauJuIsTdZNHpO+VAIopM2Xb1NGPtZmxmPQqOy6/Aq
l3fkGGze5YZ7vKpDFyqYAnfTNONTWtFeTBBatknL9VXBks+DvEGKNKKEsKq4
U/HberOCQHDevqxkgyMldDIq3AwoWTcNWbx30fJGY1VyI3J2+rG1hmFCBl2v
A2Qi85zCl29PcjWxtDPLWR2IX6kQ2D3GWZpp8yelrJ7hWUDIyZq51jSt+MAn
95gx3exS58tGi/uLyZaONC6TKtsMwXKI6PJuVfkquTzXoorLfNk07KcGCiHv
e5po889OABDcgGImKlEHTLHAJuB4TayRqQl/to5MCWFKg/U85E0MANA2421c
8EAmlVVZh6BkXH6Y+B7NR7XIcJqYiOKu+Bs6aJX391MWKRw5+kdMUfaWvZXb
bd7nKAakOjt8Q/yT4KJk+DuQYjFsbklbVkAs6P6JPUaHbzJN62XjzXs4mM34
0/gKFyEL7mF92Ed22wgXdhKH8duQCSeNAD2ybWCPxojORNcNAZ2fGGQVdLgn
PLHq1CbWCJ+q+8R+m8IT76Urn2r+GO7FNVpCHCsxxDIw+KAYkhb3Vqo7aVjW
65DI21wxYVFm1GdTchAapoMYPrW3DJhU4ZzZD6aQcs2aqErsZzpI9W4dbaXk
r2TS1m4/y0+aGCzGTTTjaUPy9lA6Pk/7G8g+mW1gK/9dvDnfjar4kugrXUfG
ekJ7bX1cz9miXeHfqHT8TDcjUC4fN493mOXKxWRCKQxJ0h3Nlza4927ksk0u
m08QJ0t2ChhvzqeDHzRYaKdxiQxOw6jYa0F6eJUbmto8n/Mz5HZALE3ESoVZ
1d1DYSv8f4U6geY+vMEsYOCa68mu20yuxjb1spYqR+HTOwgiH+yNQSMbu6cU
JBD8kxUJHyfxGDoxiDEm0r9st08JxXf/1BA57PF63sRhQyJsb6KgdBZrPS3t
K7s5nwWTTgUBfO84WuiYhTDbzMByrFGHupWg/FjT8IvGpyyCXww2X/pW4aG+
F3a8NZ0fX0h/jqOeMrXfH6TP/eHVY05GgKpj3UV93kivpkmKJnQ3KTarhIvI
N8fnTYSuAcuWQaKSW24/H4P9Hfe4ox5XriU9KEwuza8kAAey7F8YOTAZf2IE
qve+aLkEYuU9SbXJWnZANtv9jBcZgE2s4mWWZmfJ/jcsaodhuQFyvhlE7D+1
eXST6C/UM5yLveKkuR9n/LggP/J3lTRcfB36q7GcXE/ox0aIWskfoR+PjGUN
OSkmIlXCaWXIlZyH6GmA3FAHrQHyFQQ7d5B8oNh2P5Gtnlwsp8d25cg+JXvS
tNkKXImi5A7CHFXnk0ym+Pj0R52Exrjk//nnqGwSLcrj2+7ocKP4bSUdWlFL
4LLkAojhlBT9G3/kvVegJ7iiBxYxgJfpbDE3H1XCe7L9mmyN8pUaEFuja5AA
id3G7HnGuFiYjP5ULuIVdYMLfqzQpW2KXYF/1SHzB7ajduho2CUylYaGJ7fi
F3kEFmDaETBHsgfz3avpQDWgagGXHaYRi/BNygWwAEdSj2+Q2zjEwM5etkMT
BZltAowvIJH091NmglS3sZJZmFM/Vq6JwD5N7onIdtwEnSLVZ7616CAfGTM4
WjbbJWMtwNbHRrZ7N3LfeP6yjAg/3APTbHDaWoxPFuRhcpS3IZbdHnK0U7SK
M+img780dH/PFLgCET3xiNHyjR42LCh8CB7hDDCx3pbZXJkzp5ZE83biURh+
iBT2QDK5J+hItSzAysGxvdQ7m7ZAee5Wg3STi+x0rHnMNJlrSQz+RwuFFdUW
+76CC85Only3myxMMIdGZ5BY3BLwqlUT8yDsX9v0GsnfQNYcU/6YDmeyQA1w
lq22theQT9wQHbecA9/1hkVzaHoXiuvnlwdZsl7DAOU9D+VJSvigE+HxYIjI
uCIAZP61ajMXBtT3o4rKtphuOKWS7LGZ8DlkjxyBmH7yQNA8BspLH1rk17q4
d9VPQMmbb7mq8sLsC2F9YOWFnd4EXn+onmQnAyoLulnwzpTv/LS7+zODZMLH
L10bsUULJMKEnyyiV4RhNr5tDx0ITYNvNyfU360GwJopgazE/eDQ7YHpYQWD
laIMXwXHk1arNJ0pRbih7QYhsVcWRLzZnVWjA73xOaMVE9WUMviUT/0HfREI
hHinVLtDr/zCXmk/MxddHMUQ25h5exuinILAcHN/NIx1CWsGvMX5bMFuowh7
8UpRYSVLycx3HUgaND6oXERXD3izyk6MtIu0QXqpKXVH5ulXQfzMnVxoSj1P
qea8PwWNYaGBJeielB64aI0xlkZvZFk238CSVdn91xItXIym2E0pwdRq6Bem
0ekz39XHZ/rp0X0g1XUELTLOS4BuQVx/7P1pBkeB4r/HL0AbTOVdZExHplV2
QGIQJnY5BC6iqcbEzebDIJqDDpkv6bluDpgujxUbHdVmDKmDaoiiz2YfslVY
2Q21uX6jyVVTKpZqpRh1DwKlSLfNyXcy5IMtgp2Tjd8hWhhUI3c/jyookUcj
dp7bfU6cL3RUQhzg2V7F7em+lIdbld7D4Sj/kDGv4JZawKOsLHXkFtFpeVJL
x2NDk4jRbWDmxyrYT0TJmPSWF4/RwpPM6nRnUryRFEPGelP61fB8kNiNOBQC
vwJeLQ3vTaXeKcgm55P/voMKePFPYJxRo7/8gq7rb88julPIqfQ0/cdJ1fqd
Gbh2mQWJlwsIJ2LvpSxYIzwD+kdeomiod9/W/5/28nHfcgqpuh9Y0gInr9XM
jvGETJkvqI7AhSMpxfWoCrX/YS16cJnl1KvbknmTHH1ONyQcgYdu47ZgTEon
YZdf4fPghHFHMw6v6GM3c4kGQPiM3N6RvzjoXxhi7ZP86KtS1tDN82iswofz
aRzpbZm2szPqIms1ZlcFZnuLv1fap7YPhXX7a/SjM9WS5QjHnBVUWAUS/MLK
hPu7p5de1TSVpIAJfRNnN/gZ1XNd/a/glU793TULcFrOlhwv3/bOkj8ab1/2
fIfZlrlN9armGK2Ku62rqES5n63JMEN6F3dKuefixzZDpJbpIrPYqC+a+ONU
h1Ppvq+XnLRJyppYesSpmvZXlFZ8fZlA5qwkht/wVuRQapSbBojU3WmU3drO
uHL+8hT8UT8sWwVuL4T4HM9+q+jF5Hph/R9gb8IaYCtI4R7tN2A7IA5Qc1zd
vbxun8sXYC43u3JieWp9J6jJFqQoJyhRda7vxXlYFd1BGimOGsai/6lHFLlV
vW44CQZpnBDJefpANlSAlMPefJfvhWEDFjeEtMA/EfP4V4tz5QqacwmDheQi
z+b2V+Y5Vgu02qXN8LQwV+yaR6O/+iE90Ipmf6eMY7Ig5l+MnQX8mTUwRgUu
a5DuddLxIP+4iAgyrmaFUpWPNq3rayd57oyDjFMEvY7nsIa3UIOM/fZXeS4Q
lezhkw8IBNnZ/+RzUw0l09hg9sle82uFJ/UH0p51f9/C2iXetbbY6o55HT83
M7nnWCvgv/F1tDm3aUZCrfSFhb3xD0jCYWmxBjDIU1+lrIwbGXIrXWBm5lyd
IZpknYaUexWk24VlUikwrHH3dmO/hamh3v85sIK1tUdIFXgTb1BDhLG/w/zg
/FwzWETTWaAKfaKzkRnx7nFthUGoftB2jwZTYre5MyweXmD1EfwdOD4emwkf
HV/8ku2CEnpgYsIv695eTw45sohTklj8FM3cDZPsmPAVh5KK9LuktsrjEppo
9GzduuAapcc9KW03zTWSbe689szl2tV/B9vIlnFtLRkEGjA66PqwbB7MpaZs
Xubv2IcElPNC9+Cn9Towjm3g+4Id19GAgH9MIKRhJeeRzesPasoWNP0YiYAg
TOJia4IRjvmFTxouZ+JzrBT+eYaozcqrPEzwB3t2BKvMyVpChtTIPkGSXleP
Lhf80uH+etvTGK1Xg/MzfR9cBbAoFNsBSP72LvrgqMDL1ugXeUftFx723tdC
TiMgZxevlCSGl9v4WBapm8rXN93MFM/nIgKRZnB74xMqGUT3EJhRt+/oBdcF
osNyjlxi5l/VBhIhs5R36sOuWuzve7WAOQ+YGqYdRafy0SOG6PKRMDfK3jeH
hmheChi6xYO17eaz61E9NkdfmajY5MSSfxBMQdgCtLeX9dGhgjbNLhzqbF1F
ZNuVcv17+Rhnp11ZICEvF13w7SpWmU2SXa67vXgdrk4FxJ9hv2Y+8a82p+g4
+XZI94rhAootGtQ/efyhbiZHPwAqjBId+eW0MAvEy24OMe9NEHSphZ4qKedK
wLxir3oNc44PxmAmYVY2UH0qSsXPPHXztFk6Nrb/qWxEVSnmMZU0FgDG8XW2
I0VzEhPsKHXIO7YPlhZFjcB5lD6CtLwT0Mmuf75OZmkloVjZQg/63qllJfpS
xJvusoTN1VsEwno+wW7Oghhfn8Yq/mGXTFsxsMwpTjZordp4OrVW0eiJkPs8
W9/gm+yCuknFbqHKmyne9tmL/8biGpd/a5d/hlALEFkqIkAXADnvc5k2NBKa
vbI2JBA2RRL92wVkKUd5j/b2Y9rNjbjw4+eyZSjJnK/TNh7f7tfD//aM4txN
tgUgb7bTwwrCMTHiL9xA7V9HIuaJ8Wmva4wiuFjLjajNkGr07D0zpigPK88v
a5Lc6gbVBzPRGzPP7azc+PWb+ywWE3KcAHNPrwQmRRQPMldS4Q2Yu3YaFh2V
+lbiglP8YfoecwC9qTTwqoZTtFNK/dMAkCBDDq9FOxMVaXs0nB79ibDSfXH4
N5gYQobIgPPI1WWL5Wf6XLRKQHJqKFUZATr5j5BmmlJ6mhMsxhYPPZ5lREEN
cOxbSB4XsFU+jRF9JoMjlEsfSJy7EhaBr3/4wTL+fVSrfnC6MGfXOwSZwA2s
y8WW+u+SIfO9pD4vk7h5QpFtMol4n1jvYvIrhHT08na6qPZEU3nE+A/ToFT6
pQwk99v4cMCwnqJupO8u9ZK///Eom9Nq01eqZUqz5i1PI2EpAxyITOek8G4T
oRFlkTP5INKZJcMBjz5QSeBibdxW6pApSNePc0sM9oJR6K5tc2IWKKp8CdlR
fh267Vri/OicKhu915KlogSQRRVUP/TXo1MnDcAXR8wZpSMyVEKArc9Zreyd
WuqDgympW1u1y4ugl24BqwlFIx8Ws1q2JS7fKnyBDvfhiIy5D2KdtuMVWYzC
eY8UDRrcUcE2pLh19f8ekKpYq3lHkcB+fK9F0z1+pYi0RR0VTMZ7Gone2fme
y7kRbpEJH/NhwKxMmz56Lnka4z3gdXIB345jKdcQZPr5TagXswKYIOV2YV0j
pjJmYVjf3ozPg2ZVL9jCui3qJrIAKKisqseo/RKTxmU4Ya/UZtAcobGuuc1g
N0RQNxgc2PnOw4ckuVBR7w39P44dpO2h5r/70cD+K3ldIa6+WL6V+vDj6bMC
yspZTIfbay6pgn5ilPJwG/bTZgmjOHmKIFHpVrHpFhLv2qV0BuKS0WIqRATg
7bTqxNM78VUZ7DS7g9ayiQtt6lgTX0YGVNG4Ww4D9gQkgMlJVDUvZwGnU9Pq
MzhERxfjaUF/PPnDMJbub399tMnJxP0ilH5drqyqDQkJ3AZO30FYpyU01zhA
irAW2k49cJ4/Mik/D9VDu2mBU4GlCpwEA6ZpQce1QKuuRynToCaCMOqkV71m
SFayUGifxy4dyNUCfoR1BrzDikafVowreuO+JAxIDZFjSdd6mba/CdSMOkaU
VshCbm/HdWGMqwJOqjCIyGqU6qY3oLv3latjnyHwPNfm8HEpKL+iHB6yFXev
E32cFH1D9imSvPiYkNp7hfdfzHr/LKLaeTFIJD+0+U4hKfV9E4q80DJTpOo4
lT/dP4NX9rz0flhsnweEcB8U4iyR3kYejz4/gGKPqoWgAS6aQtylgaJERsff
fyDP2X+lX54udXYOd61NWPh+zI0xGgxkAoKghQ+8EkVUIq48khxlK56LYPzz
ERS1pViaX5Y9UsHjIniklSM1VL4OEIoOxWg1DwpmaSCIXK6c8yQcxU9q1ZO0
ZG+DFUyp6jj80uq/Edchkp/Wn9cjg3/Hm9rf/QauhG67E+CGIZRTv8/lnEjv
ccJ6zVKmou2A9OH4SDJW0U9wRxuXO0bXFvPSzeKjWfFZLKNEzqbCZ0+5p1GM
WMi/uGXdQXsltilkhNCbLzAN5el8M+f50QMo3FOnF5YbKepfSoHwDwNemr4q
LRedj3x5kh6pvkRR0u3bcoTlQHaDdi8FAsxpTjMCUlPQFHjZ/dytzBBaP2Lk
VubxyFTUHc2Ahyo9qZgZCiVVl808cTFaG9MPsjl3W1mhzfXxN8LSA/egLjTy
2H+vcPm+uKwoOeUW6L3e7hKa6PhNjazcpEVMvX2wb3c7bpA3XtKyZ8JbuXRC
IjpacOa3a11xhc3Fxl45L8QY/8IHJwMEo5T5zjeh2+vZhoQF7zt/kgczM7fF
45x6ZIEMsZzASPvzROixY82P21GcBvSPyNg4Glnzpwawxn/2HJmp2F8gsisf
QPU2uIupLBBuJTeFu7udkwPkXpZIuzkzGPvciL7QV6jnmxdysONE9iWLflK8
oxzkXSydnmkz3VZLsrXkPV3oWRetuLUWwpdajj8ifs7aObv08jZe0NN5p8On
vg4vU7rnlHv1mOADax697EDSqhTKMVYOY/IBvM11q/dGb7rHaZaNG7HougoV
qSs2RIBYrVC24eHcToU2YNcwcAZx47UL9l2WbxUIEeqkJ87G+/zzHxdq9o7D
UhIWonqYPlBP5c0CmTluKZ//rlSvRyDaJlrf5U17EU6GnQjCSvme8+OeVxqh
pU/IZbgzcRRzuIt+LTlB3UfO/b09IHsRFlwF2zn4mPIKT72tFshTgHtgVAub
mmWRsBlNXwF1HqtT6jWJg0Qmfkgujk9OEctNLGAADnwkBQOp9AgaIIQUhniY
dL7k1UjrmHY75oTiqHkHDA9NBHcYOc8Guk9sKVMZggM1oVoIyffQqo8r+6S1
/mVGLo+M2gaNOdSukhvgBjYe1eSLQtXYJcvtiTHa2ZvMRzcu3bfe+HebI9Eu
QecynGjVTgYSYt1ruHIBuQ8BLlPy8EpNQRDWUUklTMP44eo058Ihfok+UHfx
jbeHybNS5s9eE6R0JEowZ8vk/cPB9ZCb/e5pJdmrqBP1lMa07/0P7P8cLnZU
d91wA5l1918Bf0yve0F7+ZNo45iRYuJwrdgG8ADO17p8CznNChiMmVL1itLC
QoHtZRRlIdENYD0O5oaLDZcN3zs/1Jq0Je56HXoIudnBPxZOteKfBdKjd2m4
p2j/Na1a7aGCfPEmJg8CG6fx0ddtCoDNf01bfNw6m95P6FjHcrqnFBltteIG
IevKZfsJToxis0oLtg4cVEbXrAKDiEj2ob45pF+pa0RX852v3bzlaAlNUmJB
rWLTpLHE9nwa/GpQ2vwhwETPfmG8zFmHxznayCTJEj0yKEPdXFYRV96WZKhP
XDJ5tSnbqcWDgmCkrHiFN6yogkZLUvmdxSQjMTvT2oj47MuUAMkT8iad22QZ
r7/gR/u29yjrvRT2ThlhTz+AwDsTDlnpFVMMG5Ty1WbBD4W+4asw0LtohhSL
f3bHmki0pHDPxZFAhI/irJqkZRqg1y0CF1H8vWnOklvlloiIsAqWlKV/sLbe
gRbB+Fd1Anm8OQTOEcicZo6EYwo5BT7GCst/sxgWBWcHNP04PoK23OPqLgW4
0geYhwxZEc1hV81n6wmkiuwf6CKikq2yBJis2+Bu5Dvsz8dyK25j2hWaPNIN
hUkAgtGLa5VWYHUbZAHeN9k5jDgppTrUyZTlLgNGLzgiU65u1d0hIv/4lNmG
j1oreN8m9Vk/aKXypdjV6FdGghZzlJ0alkhzhbr87bWXjmwNCDYtnIBSbtGt
kYbkiOL09sINo0G3Obc+2Lqq5uwwfkBDNeI3hcQD/oyjaOgzWNQGzSXM793+
OfmUOel6ONv+1fR8C0ouztwy7ZYqjG4u8Z6ayhf1kUEPrS5Ej9gDMqalWoHS
LcWbW55goNUO7pxwQ1Uw22naFuGM/HmlsOia53CX96LzDaPQTUSEOFoiMJAZ
sULpc1Qtb5SzlN7FD/3R+ZPCVA0oCy9zgxieJX2xdufQns9GR/VQCf4tfGJ4
4ZS0FVcUNtmbrPab0BjHfknC1d/SzR4Bp89cAKvMqwemZyOBpTXMXFHXGH5v
PGLvBBmKW6E/G6vDMfzexHWVfmeAQBsU07UuJmhnA/yRi/7duS6zeo2GpbxL
Pq+H/+zQ0+X1hbcvV0UVOGeZEwoZm02bmyvrYMyaQM/xIwAbnEvxrxGZB2Id
j4+KYc6dNRSoDPC5iziMNzO6VQgEnJjt9ZfSc+O/6xUNBLUP+5zrVd5jQILw
QYBwzzNA80B5gvwW/ka7r51rktFVjRxhNOEd5QI8oxKE65xDFagbkhRZms9R
srnOxs4UhKg5/nDFpDEap3eseSIIdTZjLmUacj7tJrMdY3lNEQfY/w3cwFyr
RBxLJw8kRb5u0Axz6A1cgxYWawM/aTfiwZVXSQlz3Nd+pk0hGlvMfi8GSLGC
LxAjTp8AMnA3PfICh2qet2rcdWy9h2BmN84yaox8pPxZcWjHMtCeMIhSeQyS
NwrAgM7GTCfOSWlunHGbEICGM9stg30fwDiW7krjjZVdX1Yf8WM87viUSC1w
GulpKp1lzFkfManisf+2K8Pf873IiPZvsej7aij0je9CmzB0VqVf69xrvSd7
2tNm4gO4Sr9GBuSV3HtpX3FFUaphVmVSQlm0NrnFnRo4XXVLExISrqsUghHA
AYFT8MgODtAjJY/+FYr5HifQKDTMKdAb9BmVn4qBSmGyZoUQo07rk1QMOkO+
2x7/UvPAz0mCx+EdFyoF8g5XEuNn0wR2v54+aegBYsO00FAHOWGvfRFbJbsV
czgAGkw95ME5yMjyfD5rXYoqJjHjfG0RDNdNN3RidszIhgtOiaELmhFMLnh3
L2DUz/DAPyEl4FfuvfLmtDj/krNtyFhFyK1gi520dISLl9bWFcY9zmhweTvE
1X3o3s5pT3T82CP4OZemGMUY4gZom2cL0C9YdstOi02Ss5NDWBd80F4jfOw3
oQPMZ4KZu47aW6ULRszNDlwD6aAqroIGKYgM+zyhAUtMuw5zENVTwQgpCV0Y
fIjZwshsjdaPuz23T7hxL/Hh2KbBQI6bsKHT6pN8t6491+phMMhNnoUdt2k+
tygqacj7/LQyCNLLWRbGcmMKfMtjYoV+GZC8ZP+bQUcMZymvokbqvRQS8ic9
Su4Wy4NmReVd+7uJSp5tetkaMYq6+RBg9ikWL/b3cbRWTsG8bkfh/TDWXD8c
lEyzC7Cjsm9UNDKi5vRDkXTdDlYvCaYd2LeJX367iQLrS44UG4TGXIQ90+KJ
+XFlEkl5sU58wYD7zGQxiMribqzzgyLTCSjIDdtlN7qu1uzCm9NjvCtTjrW1
VIYhohOAeKUBpD9OFro2uCzD4dUSXrAfrTPEKN1A71yxE6IHZDP6sCPs0ion
EUoeTngGdfHVJbile4Ic4FX0y3Zdk4lxM78Nqf4U3hO8e8ZlSp41jDCSf0Cf
VaKeeTe/WhAnbs/P/+PWrDEpsyuZ1TqJHV76kzO1yPc2cOqUKcHuUtoHVCxy
MSQOe6mcjVv9uArc2uJMz+6lJm/imBGEVsIWGnd+JogHdk9hm9AfucQn5sLo
ZJvx0OGxXHdh2SrcKWadhUiaHg4eOrgW5sLlXSr09Cp5XbNR/MGAAvIa/EiQ
wPOeRzYzbORCr6O0zWYDYYRxi7fEUWmvApIsugKtB+7pQm5O7n7rbgi0QQ8U
s5kiE+8dMDaR8O+IV/Ek78nIj1nrgRRnKRro79TaNlw6ccqEu0SH5p4cTddc
V2qO3/V5R3WcchTcBt/fRQ7zitK9J2gcenMrfSaVOhuy6lRubtqXsiQINN6m
p5oDXHecCtNLeW+kKnEpaR3dwo3r25REeToviwAHfLCdOOATH67ObQIc7xcJ
exoPtoQXMy5t9lFBZIC7rpPAUs6Ajp/4gKQDW/gZOHkkUGIpWR4/5yBBeHcU
TvqTCvKb/ogp5fYNE9SujIb0zPO17VUbJEx2gUrgDFvBVuns4x9NAT1DM/2k
CJyohKClVkemh9FMYgndFWzP2UuEBWmtvNamOfIYrxasCwoecPbNFTvUv1hO
i6p5Hjl8xqi3r0E8AIha8YtZJbvx8JwcOPETL72KbMinve9l+ax15+jAMHR8
Ikgi/ujgf7YUgrTd05/KQSyi1xk83ECPgWUCBV7/VU3aFd0xGtdzLyUjRIuK
ftPUlOqf2gm4erXQV2Ram8PQPbSWpA7Y5mRNUeYWW/ewCJTunveCK8U7qSip
PPn+biBX+vVi0vVsbBNZf1yU5FHpSktxInuC7HAv2Rm6hOjTX2bhq6Tq542f
Hp9egK6IBSi2SXFGblyh7eR+oXY3jcZHrE9a/2YizyxgkiYiMEudc2rgVO+e
b8PM0kzEet3kOKHetD1QR0rsSNvmzfx39sRegTEl0yMvmcUNBhOPNV98yObQ
DUDK56rs4+8VSFn1/+cQkIo6QBvrAus6pXSf07uEdFGU9Nj7A3P+4Xp/P4qP
8tBNmuvg7F5icT4owEedmTMPapqBlGu7EiTRtACyM5fJCzXRiiMquteTCHy3
9fJ/dKdn+oIEVWFrzctDaxJ/qBNhKEFPiqXbcFMuMCGdfCu5tlpKZDBe1ZQP
rLosxwcvgXkRbgYtyR/loa/+8eCmJYqzNuItsMdQnEyT8YlD9WVbwqXki4Bd
mbYPKfuTO1K39oecVHwDi5ISgfrCI5NflpI5FZ7wnyaUeB2J9X3F4fSIVfMo
vj7y/410iQq+cLdOy6xKsgPopyWiAfxGmWnWO2o+HFTklOJExyYkkfXknt8r
2rJBDxxWFFWC/Y8/lyMGzjnvEzFnoWU9kuKwJtdIux+sCy0WVWM5cbyrMhh7
SZiCsis9xk5p+jiE8cG5SMo9/6g/LCEOm51YiOknaAmnQlBPxCwBGCIwx4/b
qDnyAmQIlfXbhBwI5Kxe8cxO0KMwNWQkVa4ojdmvxx+jTTeD+K0WC9cu+cL6
5wLhxHgviku5ysAj1B7uMGZ6XjBdxznm1UR/aFBltbiPPMyuyxnoYHmfW/L3
cOxd8Fm9wMf13nUePdPD8iFtroYhpDpxKCnipxoEUP912W402RIQ6s5+1RNr
8bGkJcseT8Og2D7tRxFp1Mm5qtUAYNihCeWsSNJI2k7W8/9ho68tv+peWSER
XbLgvz25T+ZWhurbR7r5e1XnCcGi9JQArXrug7wgvZCtdIwdLQEOsFY6A+OG
QLv1IG02QfbTGI6oUWslGINv0siGofCTSJwOHm4+Kydd7fszgWKHF/cAhTki
MGeaMFKG0JQ9ft7TYPJUjhCgfelaynz/Cbb9RzwdrGFc8uZ7/ePoHIdApxnl
dqdJRlPW0BlAyhffnmubZ9OREDSVXSvI6VM/t7qWt2DZSSV/HLuom6+MN8I3
AGAD6VuJzGFTIY3k75qje1cZvjgB5gdoXLskCK8sKt/xf3ql+Gew10gnIIkc
hopK4wI0A1U3X7M0IV1P/AYIP30E0WzPB2Q7EHRquBGBkRRQBYMMrNlgvYp1
sJmwsp9clR7ZIdoE7Dudu40FEbNq41Jadh5WHUv3j7mC6/BDy1zctjKx3Cn3
7cQoUywduS6gNjPOtlEwuTurGYcnsJL6LKjE6e0ng719xJQcjUCsR30U/FYX
N+7p3uyMqtJ9d3yZhDBSfCnfFI1QcE8L5P8uGDd9JgqWcg8b/T7WL2OSR9xE
/pEiEgl140hLb2tyv/nbLBExDwOKtF1OR/xcKkWRerdtgRIYvSBsu0iRMAEQ
lG63sNK/2AfAYjSVQIcxR6PiwGU0xqp1I+PZFdmQLGDIC0WkdhTFG/V0XUi8
09x6SG1Sk4sEvHfN9i25LagPwIR7Mj6S/zcWradkizbf+AMOBmsrHMkzuDBM
jar/370JYM2I9szpGhBtaVPTBwodT5AJN8Yr/tbQ4CzByMXOvE9fvyUXzndP
njzOL3ao9EZ6mHrMkvk2OySCesDvE+OppQbeTA/aNoBuU7L3+yhyevFS6g+i
/tvsYfwIMUr/jqzffoyN+OTMin6dKHgWV1AZ8IVAbhVnVzDpM4/5e6om9GvY
mfku0lPDeP3tLzRXBUHoQlNKuppwiZfOshWAnn9ToIh2yaqQZsLTClIr3nMp
2K3iJRtqMymy8ecORLRGfzXd+cBr1MZ310ejGxziWW/DamL74PBPx7/mST0U
AqXQta8/igppfQPjvbf5+MDuad7j5J2Qqu7+XIXe0QL8FzWTJsAs7J818FvF
9BkEitY9wb33Wrlfkr3DnFTLUAYCuRozh0Q3G/gPw5xmZ9oHtGMk8TC6j6bk
UwT7txeHPZrovM/GVi8hxoO7LEGafrcZo2Nxhez2bSn5+xs4XSyTbb4CG8l1
cJcFPu1rNQLSA1Ub73+De7vjdviFw14bjtzLGpJ+qRkbttk0qAYGT16KQHyu
zL62UwAvqCxToyLMmtaJ+5l6Tn/9T0ksnd2kIxszW/LVoqZBgR9J9HVjLFLW
8PBrjw7gKWluBQERZU41D0kUCU9iTbwmRtN9z4tRvX3J/lsQk3j/2tO5Dcxa
MMQjbhiWpmEntPHl8XweC1LXldJtxgWiDLZqPAbwtcw5Q+c=

`pragma protect end_protected
