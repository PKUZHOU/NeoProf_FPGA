// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
KshNC8iin7l+VlUV4BtWcauBMrWPsQkC8aIXhUlNrvSUYl/k4dS3e2cDTNLEgipV
Oyx0aMpIBnW92y0LZ95ZKOmAEi3Am+y+VkhILcnjfGJRmOnOOMUsinK6bwPIzn7O
+bsipleh/t8SQm/mGy1VPGDp3oXvlVGuordAY8tJPpyqhUNvZY1GNA==
//pragma protect end_key_block
//pragma protect digest_block
kSeI6SYP2VKaJ/16e8bgPqXcb90=
//pragma protect end_digest_block
//pragma protect data_block
n1YpB5CGF7ig/1ZC65dWRgJ4ZiJTiR5xA3A1vu+J0bxRbmy65yvw3YLtNmZ+q6gW
IlzVP/cx9TBHZGrFNusrp1tV/tJlhOz+9ZJd2wSZvhquR4/9oWDi5F70xqlDMg/J
oxs5Ou0rcnTHfcBaC9mgorpwTlajo8q9ACbbScrl7lBSAcIlB2L3CmpuB0SnBN5B
GSnwhgBDDIaEgyo4ydKiR+cw2ElVV1pzaowIz9SI/HHjo8wD1rCIAN9rEkdVCxsV
5Bc5ZZ7qJTOUcghZH6PzcsBEGUw/2hCAG1sA0AOUSlgtA06Dxxny+WrFsvV2gwqj
5dzbespNI9ds636rYweC5SOJjUUB4Aw8/EmdeR7r8YAo37wQrcd+QIPRpJX+7I1t
juUmDF+z2fhGBrqEyW8RayRzWN6tsAbOOfkdLH5vDJK262aof8/1pNTjlmnWPMvf
EIccCSRw2hCPMh6YjERcqSoYQBWgyTh0k+owcZ+ZRSfL309Cb8Exg9oNhwDTHERC
oScsvp/qsdCxmAXNGphRd21weA3dcv+9tU34Y7A+TuvJf8pXXTE9L6GpUxHnQqpu
FM8eA5TL1dZ3n8ry+c8osZHPazFocL8K/qH9QWBi/pqSkdcgjMoy1djCQT1evq9z
OvQ1mb7BJVnQvcrYXvWkXQaoiXg+snUEz12yITpGBgcRmgF9Bk2PYtLQMBcLOjMO
cYOOcEq6t3v1T+wVpg0Bp3FFb2CjnKEg8DCLHCVoTG6xRarY9TNZYPChmCV7rhv1
MsfW3TWsEKipjECRyugmbQ6bVbtc/g0GLlrig6sGI7bCiSdQbi1JpDYkBZirXLru
nuzwOSTMu7OL61rj0halvSvnFGZgqeStEWTtRz4ZvpAWtuOfuXk2r+e55F3m5oym
B/dqHIrbsFBO5dDxEKuW9d83UZyx4DZCa5eqPPJvNnvUYFUQlyrXhRcWa2Wi+nxV
nJ/5BaOAH1BOzs2COdO7/oG6v0Q/yTe6lXlmV50VYZzxW7bk8W1s4w/ylOCGhMVc
QzLYpgDYUJO8n4yU1dr32i2RjUrgTsEXxDyKD1nkpggUIwEz+4ddiDRZa9X2VSzG
4TdvjXuPGpRiJfQruHXTcOKzAmHrW8vjjnmZzlK+7NgnWNHQ2So9ic9HlUIeDD8m
1TGUiXIra0smiFcoZQMeSwOgHYCIJQ87nJ2uZC8xAXk+FOmFmIR71tuJJb0uBgVf
zy0LnvQWf8VULQ0G2iOHC7Qxj8om/f2k0WMkKCF0EUuTJVMNQBAOy2pZyGLd3lML
vbjZNNl6DBrWertpj6tfRns4EdLKG/S8WzKCSci9winNedKsgfRrF1cp+ggb6gsV
HMz4oRep9m1wxQrLRyFfyFUVHq6mcRiH+p5SHXAfCrMzVKAhgMDbRY3eBU+zPKxz
pHROjWFTAftFG72kCUuNd4lLS1qCNqbx84oRCDKhw902Z4jx3mPpZRxqVQsgrzDO
OD1/PyrLNcifsysdce+nMWuThhLnUflckb0bEBUnyRC3qj/5ihkIUFoO9kkDArLf
efbDu3BQr8JgjmBDs5Kzq5GzppGCUH2eC2FbRi+3ZgmhBf4ttueXVQZZ6MBFEL1p
xLJfrspAeA+4SAuGfpH4L4YTNKxCWPVTmDcTbIEFI8P7IDPdVGmZS9zkD1Pk9KIk
5Q7rgEe6Wo54S80kwzhC8pM9g1dCx/mlyDOO3bGhH4HY0d2m+EWuayxr1u9J446W
17z3zFY4JE0UduySRvrPJfkSyAZu0zwB1kG5g1n7pOdMJRc09TvJU/LsDTdhmTvW
W9Am8JY/bcvh8O73ytg/SXmXVuE/KAteP4beddLc+ZeD1UflPf7YId7pSXvv7CW8
OsJWl1BKioGA123ROESmDAyxvxA1x9FRHtQbkqC5CVFasF9uWDlgTat/pD5X/LB4
a0HgvK/gt+ahJSWFisJmczWFOfPLvhWlskjYRfneaPFbWuATncxZ0EGBe+S2vImY
puy0vht29+/ligiRv7wpiwtzk5s/meLMN7iRRuS5+E1jMtZlvenYguRfBu1uh5lO
5J0kmvD1+1eyVdsdIiXHqFw0CbCKA9TeWLzN0gPYgDR5r4DCAoNc8myu/nsgPqvu
FtX/uaBz7HtzOCT5FDQAG+CRTLQfBfSvLPP1HdVx5hIWqx82zLq42WiIPS7qu9IY
SMKgWYpgG9RG+hsDTAyYDjYo1nbcCOQdJhswOJ/cSJrQ6ngEHK4EGxSgSwOcVcTr
mxwB1r1s9aeRbiah983K+ctSh1IEYA/JMPHCYcbR1g9pehGXUgAqbJncPJ7Oe6K3
SZS5Xbc8S+Up/aEvAoO4XxlIkvQJpQv+OuqXFAhLbtNR2uwwWKBP1WSga62HCdGY
n2KsWHUOzHVcvLI2TDM87ocfnu2NwX8lU7dM5hdv6baibYz37F3hEi93IkguaiCa
MxV4Dw6m6O7caHmLKOy6ZzwwJN/I+RPfVA7UkMTP3ZtT/bkvb9+xssOn3l6akv2G
oaTUSmHLiHWGHgcbBMOxuUsXm90rSb7GOs5+d9sGJVO1qGLnTIaPHiPp6glqYnBL
2NEBsHiEcL41FnsH3Y7WMR9/7tT8Q6ZDg4CaoEtOtS5v03fmJoVwow1m+9HkJhNr
9uAyK8fj3RRte1gdtrKN2t08QJSaahD6V2Yhp+dRfkX2+6UzDnr68+V0FJz7YTlH
08RN/b0FKWz0Muh7BNrtx9SuJNccEfN75ylBe5qfSQ3vEjJPeeZLAePWIBbLONwd
Ra3gYksmRY/Jmbt03+kkYDY1m1fUrXox2ZO9k4sifT14kWy3DV6ifH1uzOFJ08/s
bHHZA84p9EEX57pMZ8DDjsvt+nIWGht5YQE848r1SURjRyV43EyLpnKbr7l9X+99
Kf2lRa0FdqvdF8fuebj2wO9n8v9cafW63BhHEfXmDv1Gsb/QnD5Cs2JTHM8rpyYc
wb5sDSWKBMCXn/VbBrO/QE/7rQ4kQc6ttqfNp6MB2VDeMvC9/gj2TGeVa7obbYip
3dAHiL4G5mWvkUG0HbZrWnHmSS+dxTIZPCbAgafMcmNy/W0ZIheHyM/AmpyrVrwu
RMQLXVT9diyXLb120HCffXpTcDvFZWXpqz5G5IHogGK4GMHlmmUc+v1q0JW7Asao
whePUC3tneFIHhJhJ1+tdlI+NVinMXP6tnmzVi8MeWsvwBujgGjHQZj1Eh9p9KvL
DRFrwZMpn8v1pGNtBmrPiKBBs+wsPNfmOLWoMN2zWrZqmonYTRJUY1HeEepf/jOw
2fvgXjCqq/zIasFL4sfKZbiDOitngGZLsJaZ9b9gxpFTSO7FLM1cKt6TYjj5hUih
4YOy9CEodHbapWIAlmy3EvuV+dQgqY8sbT2bh/GG6HYWB2dh0+zvUBvtuigPbC9M
fUu2HhhlCqVg6nvVNwujpu882nTnusAF/J+PFUZYdHe9cpKsFm52PeuUgOTKtSAq
gwCU2P8QpvA2ZQ8hb1XxYybzSq7vSR/qIPze7cyiPBUUAxMjOX+Xrbc55iclGmkl
Q2SDnm8AbH7A7dlo+76pNgEcIUpBubXzoaVYOl+ZbNomHkQzdkkwKQfuydvsjSzl
+z7VLFA460PhZiBVjgJrHZbI/v+aAAQniZFVSuQ1MbCalxmOR158QB0dRtTI0PLv
76y7iraQ6KXpwTUQ97/sKd9xWmEZIZ2l46RGhNDS7V3ayUHr3L/iWjRPp5zVUVgM
OI3cTeVlXok7yR8y8Eotd5pRnB3AznJdrobOs4a8JgV7BVl/c60wE9u8UonAT/q6
OnVqGA93Jv69WosHYl7X9FhHAgFfAG8J9h8DaG1vEAiIiCvIjA5PmrY2ixNRIgW8
aigE7NKlxqFZZwNFeZ1sSb0m3toN9NT/9re9V+xFuTBvttS1oXSysArmmFcw+XjG
IFZGP1yul0xL0X5TEnnJPOguMjvh0Mv31QZeVoujQJvGW21djH6cXtwLGGJMqZ1w
DTBBLGJM4MvNAeygAGilQpbAJJSTjorC2235S8lTgPyvSJ+PDGXOjbo5cud2jxMR
z5cv4plhqCb+JCD9lAc9A+S8HheEHAozERs7Oarmc14HSx4m5hN6+T5eaZ6Qa8hS
XqvFDo8CJy71DqcZ9AtXIyr0xnPPw1h9bmHYjep9Pe3pYStU7jCrOjdYwQOJdFun
DG7Xn0+NmnqUB/udlEwImRW7XnExFd6uRSU6x8K2kLrQSnSZpNVWU2Ah/nGaPA1Q
ryunc1a/0zhhdpskXZLEPZ+EE9U/wrPpjtP3BmHwfwux1KBlAcI7s7hxW3nMWA7z
uuNKYFJ1DE2Spoc7SgX8jWv8icLEdREr+jMl2CrBWGdJ5bsuowuOY3p9UfEm13KI
2qteH2aN11JZdfW12Oq0FIfH+fea8XIA+3oU6wSOLHvmJwi+UBkJjKNPTnycKe/W
Zmf/X/Wh+6dmvhy6iTQrbucTdtoMQL5tVruG51LZBvMHRcaDoYJKuW5u0anNB2eu
r5rL/v8TMDfKfnWZfuJd/kqM8DibIMEpmfjKb2jcjNVQPTb2wZW2s+3zg27uoWAw
gH9wACUmPr5qKD3ZSIw1DtnQzedtxa5OOZ3IjSK7QmFWsyuyaV8xuw1BjBJNRe9B
wNlpb+MC9Tzvpj0fgfV4fd83havhDe1vTF/VbHVFYq7BoH9LfGHrLP7CrzrnpjC2
MVaN9qZn5DjY3zHVPlYNGLn3bEm9rX2scI+7bQJ9PL8sxPnhWfnSaashwC4bxsxy
p4bnADNS0KUHkBE/6bzuzDqFsF2JEdahtAC4uSGa1nyoD7cu9QzjamD+n3j92Ylc
8k0Mj3s43s9vi77NRNxYfFpJRfZiz2SQyu4c6veoMe/MPJawV/P1/L4sUKcfPhBo
6wLsrqdhPiWvvmEd37okzXXRSMJ995pubaDodpTapNMiHqcjMS+vNi5cON8UhMdq
wLlvY2/Qbx2NXjPnLjEjBuhBhDvsSVEdjCib1ompOt4OizD6CiZVGT/bbK+8g2rD
wuzCw45v1D5DeuXO6J2C7KjjKVtsEvYplervktw3aSMMBf/6ne9fLmlB6ANVSQKx
chEzcWvCql5tsfNQiZTVqjRKRWn6cyswH6KisMC9oKdTbJqakPJyZ4jDqkTD/J92
TVw1xA+hbN6depniqJ7dRjEgLnuMEoYTeIFIr9dohDOmL1j+EvflhLmxGt5R0qkx
mJYR5FU/trNylWBKG1htjeyFR0uHmMiuXPyXjUNIAj0Tb3eNyX8D0sj9tN3YMytm
/Z3gJBbhPQXVQUwLlUBPPjyTqCZRpk753lp6ZsiE4ld28LezwB+XyQ+B9IHIlJy7
yB+MS27P6uMHipjs2aoJ6cNy/Wu8OiVjO92avSubMGBHX8XnVvCrVwonHcfDVM/U
pujnvqpEM7bjbfkryy9MeJ6a4dGyXqm0pSrCpWj/7FHY6h7zF0rH3EgVhFLKm/Uh
aL7JKthKk0CjCP9IZ6xayZb6tTFSlULkpyHO2LZ94qDF9wbUCLRhswb9sMPU9JsZ
3F84vaI9xGr30x8rm6KOyzbvorzojkDdW+unExUCi2HUGEFRUxW6bupX5cD2dVIv
jVs7DyCWCeCA97SVvXB0jIQ70eop0IJ7DOrB3c8nMwqDKpgHtcM411qM8MjUenS7
FVxWWniQcsSDjrPMTQsq1mSvQPF5NjKwAxBmO//6u0kiroOro0yCMfXthI/CG+5o

//pragma protect end_data_block
//pragma protect digest_block
csZtP/TtplwDYxguuLsoKT9V7n0=
//pragma protect end_digest_block
//pragma protect end_protected
