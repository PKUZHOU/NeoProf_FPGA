`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
hHhWjuaR9z6SRS1sUwzHsWiN0LCBTIYGG5i7xhxKFYqbUwGL0kCYz+uWCEdvrZTx
11mmAr6W8Trmbb42h1qPqDcooCuq0mI3J/ksGtr4Bx7shTPLXFEgZ5W899GAxci0
f/fN9GKCwgr4CrFKIpZy85A25yrxv7jlWKAPSqtZyN4=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 2240), data_block
1B6bAfPTTR+PZFj6XZciRY73aAqcDabSfZbXJSGgf4nL+kqmYhPLPPibiJHn/B/m
8zNU4Hm+6QXOCQYUC1Ko8/EFgY9brB7mRrRELYu+nVH3qV5qrA0VfLKotj30Ttpt
qYNjYWSnt80htP/MlRgvpE5y9amp3Gf0D5WFY+o53XnzPxhUCHVaO5ksm6TrbLjc
Nt3caAx/Sz/Lgrf5KXDHKUw7QvYBmfmLpUEh+2yUAVCjcOTPpLLBew54YbDFx3Nw
DOF2R2BPpvdW8J7wSKhQc8SOwokAiTN3vFYxDgO4/e7r11BZriUryekQ20A8zPLo
uMB8QQb1/zMNO/ztbYP5UYRcDxH1dFNIZKhtwvx8DasfI6aTApcGnpxvsQAsC1Fo
JEFscWCmzPSD8QedL/m7eZcPNtM17yltRdV+hpvNojcq+61By1PUEJF0k5L9mPVG
f57EMOGw4OwR1JZffSrYGExBK7lDPFtiRn8QvfXrLWYSjsqAxpdAgNr775ha0tA3
DxHhiurd1AoxuEmPbPQvYf1MzY5KyuU3m9HHwoxnwkLkURhMLlJMXCAc7M3AEgCf
qxrtqFOdb8Q+BVGU1OQTxsi8VyHXg5rNP9Fx/mIkydN1V3WGUSzAFpW8xtoPvIB/
Qwxo+4/DYsL/dR5jqcSFJ6kRsyOLFODTmLyAvjPwrfSQuBrBj1q6ZVvqPOfFR3PM
bEaKfeGu6Ax2y02Sz8uXAMLPCn8cATjQzS4TAgnYxpomGEsdKXSDT1/fHzfrPDlK
XNXsp2KtXdX7ITG1RTKZfZ91efusSesgM0ohwvrxY1SLb7jMXXtkCXkGczSJgfdW
R9JoDEvr1ia58Q0bitiGyosKU1w436cy0t2LElUhKx+nuNns1xkQTjreA0gYCjdD
QY1RLuHsb3S+F4xLnWPBZwWKFjJ8FGPh8XJ3Vm/0XxsRUHI+HOHJECWcGILMiRpA
yikfUp9UqnldTBxCowrG/kP4Z+YqLZtl8pqfrCSXLLJ80KjFAfJbBx8ePbQfa/j7
wfkgO3cEAvD6kPNQgxO8FuUA85lCNOy4UrUYMoR9iR5ZIaYsKz0lNi5XmZqB8peT
yKjjAUs6FMPbRcHY3vz6wet3ciYyLI4bATd7hSEyCOB6AQeGMZcsnMMUdWXPTUlY
1MAIJO2uRO7Q8B5lVR808jUzgogVlaDvoNBRXpk0FDgubQyh/9aJQrn6Wm1UHMRH
uY4KM52lJp9ieVgGqgWBkTCzcCYFofU6nd/NHJR5SALjXfBAgAHMFR9sSCJ3vfHw
APgJg/1XYjYtyDV/qYJWMYHK7GgjePmL9A1gyRnfDu7wohEq7RFleSZwZIHwfbqN
Ju8AQKAdVRs+jJhNR5/YUDcBHwJAHvNSjo3hzveaKudyq3UG8vh7qwW+tP8cEdmO
ip3Tmfo4z06Z1H2S9qKLfMi2kTDd0tJf0byiSHWfTS8JgrjU9QThkWROZQhZk+Ft
Q00/kS+3/yLu5rq2rNe086ykypbcSm3Wo2lzbKhvoqU1WQCGbiWCqO9wIR9W49Z2
f7su1ByGyuOZ406X/o8RAEsC5J6Ziu4yc+oJGEOaTrgaMYtazMoSDZmDTNcHEfwB
10IBJ7h48/6ElJK2x4js5xMd3POkteu8oqLCIM3T9JGNANRD9iKgna3kmwE9CXHJ
5GBZ2q6fVSUrMwEIxLjrC6Chk5mvGw3DeYBhpRds9pAjzH/2Ja0yl7fFpLswuLFF
L6dklu8iejA+79BDWJLAV37mD7M67D2VLRtpjZXxruPD3NvuUjXn9gJXOIoiDssz
RQ8KsBExio+8jumX1JOwC8AI7yEYtRGPPm8sIzbIxX/jUxWLsGd01ORToEWrA0KP
NuDfQkz8ac1ABvn8J2pPeWL+F9Jdnv0drL5i80jG3ohdifEhHiC1qFNVZS4wJMS+
65lMU0ozYhNVW3BgoVhSw8Z7/gCIUNKK5SRLiUlSwljLDX2MyLujihi5sKu/26tP
94cSkjjZRTt6CKDk2F4zxAyol7L4b6NKO+JTmqesprKLlne3zmruDjjBlDi+EtXk
st3NyI+UpNYozQWrRV4BMjzTBGP8jE7j3AXdbuVlvqLBvLskIgzV2LjimBFgNoKH
gdUOm9yd+mRI+EeuJRUVTNmfzVrGjidHEdUNTK0sE4YKQGdg5lCZ3y48Pv8ml5Hh
c+t9kUKNo05wZjPMhtjkFmu3Mvsf4K4DovSXZJre2cyTKDzrxbHg0lT19rJmOQjI
Yf7zrXeKzEN12ZZRIgnvWc5aL9wsa7Q0Z6OEFdnu+2Ir+3NBwWTjX18DkKHpXB//
FcKfxKSnmShs7T3+kEqGzeh2m+zDL+DNipOIkF6y0IDa/pDNT2S10y3Me0lYepR0
wXDQBlXudeqOVLhdg/sGoKR/moJCyXXL9a37Dl8oXyBpq0gzj7HTnO/pxSci0kXk
A1lTuM7xouXx/6Ip4m4eS+SwJNrcQDGO8sNXTLVULE25rkh3AR6U1CnpzE9ISvHW
HMKdwqIVxJ7U/BFH3yNNrTiCr7xcnUIdbopG60BfVPYl9PJxPxgBhMgxQop0ERYa
YBKE6P26Ggtmov2prHk3QGk+rHLd7KIH3r9saMyw+ggVLlXuyI5NTMfk2o+R8xRj
Oq1hRc+XLZsuKtYMw2qGefXPWB0kiuz5CI6AWVq/GfH3fwyZ3FyjMVj+7bttXVhU
XvymULHrt7t/huTRJqCztj65ztcQuP8hpHHx+RmqmFfXArXWz9C86hcXDUbB5M2m
pr4sggZq0mpFad6HdiwrDXb0DoKFvyNFpxS67hyaH7VoNV37/dicIMpolpZc7vOW
xuZi5wGW/SuY7CcaTBmVFO/M2HndgGViS4/J2qVj8d8ZRaLcI1LSewObR8wjLSkR
iB6SZNzxmw42u57gmOUsMy6q+xw+ittmOJnp2Qs87JOcMDR0lYiqIC9tCqJwIHZC
m+UkGWJV1M0WCK1r8cC4oukhdie05RO4a1uNvQcUA0s=
`pragma protect end_protected
