// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
JQhuVQV/mR0W5hqufpvdpXvj2DEwVz6AV9UksYnzndW3F+YliSPZXDRmGM8C
IGMwNIkUXQiBR8qWf62iPSheWXIS38nr8UNY1DhJjUpVmiv/uM/gx7FLuNtT
CNvQyORuYSWvrEnOhlWpy4Fc4GLjLPqJoVAHmEp8c3vKAHvHcliJRVScJBm6
VaxPlUeBpVi0kFVLNplGAr9Gt9LSFJ6vEzdWgKcecMf4TI/gS106oo6TTZjm
uwERnYaQCQnnJVHZa1E6lsDktFSpBvGEt/C4zvjVeTQu3VvpTEQQY/FCBMO4
CBA5ephXd0VLcg0MYC3JTPFyf8qINFTjiILe65laFg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
X7TCCUNuXGn7ogm6sFvOjfz+Jx2Oc7jgbNHBDxpCiNavnv07QVFvm6wGy8dA
OQCVMlUOHQ+wMQaQV4VAKNqqcumFYpucg1FGfiWYnFOokbwtSCBeXSo4eWVr
row7Ys+NycF23IkbAVD3ads0lNnd0d2p1BWuinyLIDH5U+vlKfl2GZqRkxPE
MndvWOwRfeeGZdhQHea6LtpEisx7IccGhI4AriDgBuZWCGkfo0er+3hWAnJc
wN8qHCRbWihMshHm4ZeFHey9iyNrc0pXp4lxkZ10Koic/0gEcZSv2eGXJtz+
DBqm2+sSOKB5mabqrMi08vtznFhiiL3jgime6ruFyw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
rYMEa4pT43D6JpxzNxhtCjl8Is3T0G+9jZRMTld0a/83G0CKbRzbJ5cQYJih
Ra5FDBGt45hQP6Z9k5k2cE2GogsV20SKTXJmqaWHeC6/yb68nxTNIJUGq2vc
jAXT1uqq0FgbQogM2TwR8x+GTNPcMdrKxO/T9BbrMPg2x0EFJxDyoSwOzXi6
b3P6VxJCHt8nRG7ng6nizvNKJyHTOtkmmVzw+ltx5fM/VavtDvXQgdcCaim1
8L4RqANb0jnnmMb9QGZs6w0NA0381oXlyH95M46j75Kiy1SvpRRLxFD5deg2
Tskzu9uMgVeMC87CqwOl2tT2fQZsz/xdMmvwzpnvvg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
DaItZb+edp7r/H8iyLKaPkh/PsqrB1vhAYtdJRHuD0Z2dPU6XADiRTUDjBuG
xQmQvmFXfq2/ixA3aCI5ftTgrG75OrgnZagGeR1M/7+Djm8c7DVazy6ZoucC
A66pTM44xeRaKwxGg0fz9bYic3wwOl60dn2A0Af7vOY5t4IvxJM=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
VA8uc2wXUPvt6StjaCRhmexV1t1ETSzSwJzSU8ggZy0jf+h+f2D6YvsMstUA
2GIv6tHjzFFsL6bXkGxTkUWo4brmnY+E5Zh5aZueNpk9yRDq/aXthKl1uqYx
3JHQp7oqvDCefNOYWsuiZxNb/hncC82x00kXvUh4LVvWc50+oewRul0ODQ4N
PZi213NteBe5XkngPxOj++ykj2jT7+zq157G5/HfFJbA6DVNF08vd/du4aIT
nrd+BcCuxVMx/Z/T5+DphhTIN+zRmZivkO4ozd4/TH5oX1kyt6o2p2cHlCtg
k6qySbnYZr5IejDFLRzCXJJlfbBof1/jr21nXhgNh74LkhY4098DwP+uRALX
BUnPY73omVcMlj47qWCdxLUk7xzA1/sbPIFg1yhCEfcM0aZ2FftJ1Q6S34OP
sE9vAzu70N6IMKPAF9UDMDNfCYZcV3YzWDGlHUuBCV1T7MiLluwmVyRFy9Xq
u+rbQrI4y4r4Twg5atU3rjbS/iUuYOFv


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
BzsaiWwJog9WlxUyvzgns8IID3eyn1YoxruytsaaJ9STnP2mw+y6Ydz4/euC
vTFvxqju6Ko2orOqKiuE12xVV6YXlVGTsyexeSLrXbt3TxEvUFaAO35aNiR+
kIAirmwkAxbPh5hkN44S+Xgstn7ERdLJmkmRqz4SnZaGtyzUGhU=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
O+xlS+aRLVhzDHdG16gjbwRORtXnlPOlDKxsErmiViBAE4wo6w/bLWRv/QVb
8ydtI30bFSoJnO/H+qK2q+NYmwrE0Nnr6JO2Ice4PzzMcjiA9cr0sCxQnOsf
RCkQdhtd3BLO5GG1+OM3n+mkb28mgnzEDlLtCVY6lkygMMUjaWo=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 35184)
`pragma protect data_block
mcp2ZL/W3uUJuOfJZpi9KsmSnAAA1xpjliIpqwgivUxjbCU8EmE/CUIK+1rG
AqVW2cBnJyYaAOOgrmUpn8JXuAroggIXnM6lwynEHtpOei/lzQ7sU1HnjEmz
HIXLQ5+xxNMH6Xao1133wwlM8fjEMqMvo3aSadn0UgtZYwI7lpFzaqLt5Wph
+dBaVz2ocpSqs1D0cwE5jn3ppjp+92v88ccoQ0enMjRqTo2lpe8JCyAKxOlO
FWjU/aV6ji1ooV1aNt7vtJB4RnNmufl/pOkmZ5qqA3CZbwD7nVFn+BQLgAz2
kD8IWAjWbTYpCfHPSCD47AI0U9wvmziTUFpy/VqfHT8hF7ilnH+NAib6aqd8
MebDUVRqUiQobR9iYT29hlvrqpyY90J02EfrEf7DrF5bIJjoACvMis+XhW2Q
HGR4fA5e+eCSyG5t+f+L18UioOalC8MWBjo3qB3cAT+JbZJbhWW0jd+n+hcj
MBItJrTnxSZ9FZyNGN6Hj9wf+NPDNCfgSwUeicUeUn/p9qJACDlvqPZDxW8R
LTXPznhtr6Q03J5CWQxhm0Xxyn/RKwvbOucnkNfxvwqa94Qp036UkyAqDwYi
Qp6SYxWN2+rvwG5j/Qw2OO9cFN8SAHBDVi6bsWLWOEAxWJLdPF0fY2huHmew
Jflbep+dLpZr6Jzc0xQsr82/O1W01RjtTd2SSS/mNhv2GdWxcc/ZFwxIbpHo
KphNgSkFM8B8mj+dSiMyWwmvi6yVuhjVXccKG0gyQodOFJZoCKe/uI7jP7Ph
gKNMO9LwL8BXE0zrZk8y93nlUYklw/gshGUF5Op5c4KgsVyDJ+CyLeXxhJMl
O0YT397HlFEprpVuQROAz1nQxbQ1dMvpZ+mbrNbqGLZw5uIPYqRTcFANKrAU
O3W/wNTornf8JrwQWPFBAKwJ8J4yYTbAXzsNojAldUrAaJxqsEBBAdzVB0kz
yMQ4HE8ozmn3S4LQIhu5HeAWQDiFCk3aOCy13s7k3rQyjt4cn3Bc16Uf1Zow
h06zcWAv3+cY/h1i+lcb4VvRVYejZPCDT8DITDpSCIjTscVh3nIU3PU0bqmx
B2VtF6aAnpzaZxMgZfYWk+zMW17l3Yqes927HOlNbhxMYNi2jSwYYl4zapB2
hgnSlWIC/bNW9Oj8KP5cOjM8xaC8DDc2jN3czov/ZFSdfGvr7d8VEFco9T7N
ukQ8m9xkYwWG/NalJB6as1AzXY+zfHgT4sEqdkXKQ3OZWD3f+UGDBdw4l0Uo
x/7xMkqvxuWdC6/qijHx73Kvv8b9obCUrh/Zm4YqKMdod5g6DH3/2wOH5I+j
laR4pfRtoaPbuKZuQFJkePvT2R8KM3SZLELI9zpJCE5OlrdebwCuVyuuR2BG
zbt9dDwasv9h4ltqWXklyAFcxJLBc+Qurd/ILuBQ0noLlneAMnAQVfmlv1ow
jdhvAN/snkcXPT7RnPTfx4hbDY1Mmh7d4dsUob67x8fnDy/2z0b6RiDpQnks
ETZWHFJuFRjSInD/nA3xQrKYCaXgW4ZAs/o0xx75IiXf0NxPUWCtX+3I0zWD
t1QC30UgmaXe/ZQJPgFzOY25xM/nnPmAdDb+YMo5mGpINsDs1WyLR7WAZvtf
6Xdc/+zkYrMffgaPV6IumyOuUvAVHP9n9rtilfGjDrNcABnrgCdgSMI6eShc
JRWLo9TEWfgdocB4I/ZdaFeuz/xnNZytbEdy/tiCSpgU17wJp8u+qG9JJhCW
7n89iLWjmCGlDfZ8VZ4kTBRYFeAM5ncErRTgeHM8hV8rLnjhHgO6AQh92ZrH
avqLNdudTX52zYomBH3WoxX0twk/XSqXL6Tn8y3GGVO4fcSWmTtXmrfeVPS4
hlxlm7lv02tOE+NntZXf3e8Py8XougguQQcq3mMgYk9upydQQmOnxxB7/lOE
Pce9wliHU6wgkvnvARPKjL6+9Wpj0TfxF4MCZKmL56kjAlg9XhhMvwWnrTtK
a2ApsVJofJ/03SOy/qeFopztsnWM8fG9q2PUgk9BnNeT1dKZWESVkRzxcaW2
z4xJ/ImwOMqsiQDOMeIMuWdeZ121R2Tuun5sZeCp43G7sEi52p/2me54LR2y
Sy9ZbQtE7RsI4tlKJWJ0YS7zgnLoMO0hi8OswXoFOwa0fK5JMmIKFKAPUlqZ
VrDWyWbwcn/UloPIhuZXACKn0CCecyCxPHJSCJU66qEfb3IYpzoqzNaeie9G
qcDul+bsFHiTiAGULgls/oSsojgp4aatcYASzeQXFOklI+82yf18O5Xe3RK+
yT//0WxsJsVoRQ4w/280r7zd9uBgshYLkotD2+hyvqAVO/hNVn/raEIPLhyv
aSRN/ocV3/5h5qoNRKPLVi8T7bYJdnMO1MPKgg9+29bh508zFy47F42w4N5U
MeZkndqWY+dCudoKXaelbIN8GypgMF7xuEJnRd3rKkgP9H249jenVhi/k2o8
1DcyEnSwS7JKPlu+IXKwUX13v3wgNAij6G2CsVZLXK0eIB/EpeDtRZ7Pt3YK
awJjAhoBTscwcaAfDphvxQmndo9KyeCYZQeIrb5fuW8fHHH/X60zwWqI7dHb
W1pa0YDBIOoxkFJrJmD3f/pQCR/VIx4VCxGdLMHsVkMvHC1ueMIEGZlRFemr
NhUbtspNaLl3Q0uWxS6Dz/zHHeNPhLoChSi4ACmLf284QMQfhdhMxpgm+RjP
42ptKPZj/7hx7hXA0Zsblgrz7isdOTmdniU/EvToUrV6Gl22NPHYpc3nWGGp
Vs8oLCkt3u9PW+8qigOmyBQwY4M5JDcHbO5o0e/Ig557i8h/W1AjJt8xqojc
k5/qyIPh6OaqoMqhrC6+5loPp6O4H37OBK93VgETF3wMiqrSGukm+gbwoqJT
RUdL9H8S62llcm8ZPhaRBwa87pYCHZoSX/K2UYmZXBLl7hWaxTGkxd07dZfo
F+EgqpblCS7YreT67/jJGGPO6k3Kv527AIeMB+VblRXdPdOXCPT8hFjlEB6f
WPfsVNDChtRl7z9FhRblQakvqj8x2Q5Q0NACOtUG4aNK96dtMA+GPtNvmZq4
V6KvNC5bOEj2Jk3V/5a7SOxcAfYNblX45GoyNlG4leJlzqgpSgscV6ddtfMm
BHYq7VTpEhXmm1YNv2C1NrR3aaZgZtAUXujWTLrZbYiHdr4yAe+CaffiREvm
ZpruHitIN8htmPc3ODhTPh15ezsVLUBOhML53HmPV5NHNDGfoJKKVQCtPT2t
3a7vlbSG5PLYGBfvrxkieOi9mlFs8RX9iGPiZv1Vlm8W44UH7xJteNyTEy4u
cxoPioRScLLxLxk51XDlWkb4BH4T5vgNFuyVYI+rwyUCuqIfvI4KhVRfjIL4
pkbPCy2ZpQo3oYMbILnmCTES17963igRJfZttlpELXdHTWikgMvKcXzh5Tyv
Yecd//SLI2poLHYnCvmIG8J5YLXCWrXNRqTSdXZ6sDtvHbne7OfTB61OTU2M
JkM0nXQnWO7ELUQLwlpOHx5CJNWSXRnZaBRU5gg5brEJG/2myaTmm5K6ttsi
WYjtrbrCcnH26lGloUKOGABfKoVuAfYb620Kv6DpnfveL4gwrzDFajcV+VSP
u+QDx6SnMGjiAKZqEQLAUTKXQVfTJzL6uC4Dwljem3WMbIzvj4er66nDuMO9
cbfbuouECCXsVlywWLGcPGfCJ+ZrOceq9YC707ebYGVFZumIiTXvTk4GqPeh
g+fETikCTASBn7HguNZlMdQQ9W+d6ivu8euOp7oOPJxR6GZt+G+CMUT4PiSu
aSC9GvJSsOC2waC4psrKNDbahuplOlZZAJweP3bBp7dLNqa+Tcm8ogo1YPek
4LlkPez+EyOPmUnwZp+0Iu9xBj0AMrvjl27PAcbLGzx5KW7ANdBYzBzDlYRj
738Yq6Ek/BLRrBnBYbttjxDLAbHFMH0H6rwT/AD//C7xAiaar6izjDvQNHJ5
8Z2SXB5Wu+b4JfrG8sYs8+rtGF5bYU3gschSwz+68OW7HbirjoZPLrQUovx+
YDpvyRlIttfJyXp36DLyVZALGSzV9xJSYF7LXxixJkDXuhxV6sor3IqGG0KH
OgoA3g0NIOlnaYHM6WCEe8C6D4HnwvvuoauEpVI/6Y8SFJ8Ltqqmii8K5hVG
O44hlK91xctI/QyFU6fGLUbaCKHkUx/l8Los4kY9ZfvKRStt4ofQAC7yUyYa
FTNoO59IrR3oQjBzDv8SmQQh3YNsLqAwR0nX5RtGK0dWzfR5QKV6UkM3hBx6
X287L+9WD8P6MD1d94HRoqHt8V4aic4ltIcW5L0fkd6zVcjSvtSx/DHxP2WW
TuTukdNAUD14CrrWnZS4MHKOH93GstkVvGGJEKILGSr/ibSSpYtRhfd0mKt7
e1x2abLXyhBwWyqK3Z0kd0EnjoaW+og8BRSvu+7q4c27ipjwxdHyUoE0o9TH
Xuo389p40qkmqfC5m0UhlhMJhkpq6Uh+Lc9/Rsuy3QPrsKWzoaPRiltroF3t
K2MU8u6POIiSiYtaajHGeQULbFgoOR8wtrtzXaqQw8elegSudZn1vJU14Ch/
FaP/0DSH454BjNwLCXwQi614cl26u9dQz6zzTL5jiUwjHum8omjUCozU6uJr
BL2WXxx/DqWgaUhD14/QuTWq+IkAvhjCXcThQwRrs1H+veUG7KwU17NPe+8B
gAtXeCusOv3nXp7+a/SUP5lONVjxVwBepIzmXstx8T5TIUA2s5V0iuZRJ2CQ
JLuzNu6QELBwbTdbVs9/MgjcYtTznUkbB4HmmlWS6REPAS0Iklf4PYOep/Vb
+656sXfj6sy81QnpLzLDz6JYnCuWZzM83/v5hv4ydMlWijCrDw+llcfBlbM1
+J1qVobRg1WHSgrSDNHuWZ8pkW6gT82EwmVqVLrZmDQoi5LOLUmjlNhCp3Zu
GCNSBHryq82MuFi/YGOzWY6LVJKnU6AhdiMedFHiTUOFoXaXzKuXKPIjWs2U
qQSPt79a0UNXP8YZmY5XrkvQuYSEPq8tbIHKPMEecF7TPZwhheaOl3Ui4yEi
UUu7TvuOd3Wrd26BJJnwoWjJESWdzAhzyUIdqql5lewt3ZX9VEot1pQ/96vE
nP8iqn9SevjVJN3jCsHkEebHny1vF3Zl4iID4p+6B4i4HNa3xoUfigCDeC49
hZhvpU98vejotD7IPPUjqGcPwEGAajM1C7jMgsO3zKwoVzolcT3qaMwNj7HA
XbJf9vuw0PDhkiJIJKaYPksugRxOo3H+Rg+qkS1nftDBmmTBNsq/D0p7IlzR
wHvMW9LAuUxYiHi92XsVv/kcMG7O6b0bYz62J8N9FYcm/ituh6pQB0ztVPq/
WlXeza36pVVpm7M1YJtaZhb1UhanPbUA3mYC3YUvHagWk+LG3mje9MGdEvq3
pWXQCshKX2tpkdJR3UtFQV+j5lCyAaArktBTADTy5uOBm3JUqYTGJKbQiuVN
8PsOvj2gL3J4XRLny+2UTre/6Ba+yQqsPHFFxGXqnZO+Nl/cEXXpP6WbTIGD
28dIRDkUfoITQaqpOmYZBe2kc73lq7aua/g9wyVCMu/KnP0UnsgwvotnEUAj
3YVtGAjBM4yeg1Xy7mv1uJK48VgSjzjMUANo7XKucSMqJ8jDswM+yb9XCimc
SC2uab3P5FuDeMWxR/iSUEDYjbkUzVsQXNac5Q0+AsP1clOrQhVisKcyNrjB
fkgx0sMgzwMlJ+vp7lVIVVRiag1sWFlHO8MdH3+ETxyHLwCpa1Ls9y1xCbQZ
qLN0Nru0mvxVRWpMs/uFGPhMVTvKCWYJD8JhH0ajeVvviPHpMAMTJC93wstI
3pf0e+tG2AGOt8I0Q72AUxEW2gRrm8Z7Bs3LrHbShJsJLYZkPDvF31AAJSO7
rQjZX4nOrZud1f10L1nLeS82M8dNpg5Qer6ApZIEAKU/Btq/aaXM72ef1lm4
S5f89MMmfVyiG+1oNhJfLYvsXZ0AyK4u5Gf/+o8lcToAbEt/9orxLku31tss
eFgTaev1Yro2EwqoxOQ0ext/x1YAQzhFPZBtrFQcZEc6r1Wr6wQETLCvCUck
bkKB7Ox0S4Lnf2TI+Z+XwDG1qJmtZC6z1HBu/mDLs6tODHObtYKNpos5Zbm5
rSxoNRWCOxFPPkdkNZXwv/uMbWBuxQWpZ2YbHURCM0aRm5ymb3tQHVr66IbI
LHYGg5IRwKYmMz2Ek2vy2CAAaeY54ev2A1gee9aPaGw90VFlRMkGVwtSXT4s
iiwPntybYlsRX47U9MjENTJdVymrCww9ujaByYK69mNeWDWAwe/DONSGU7em
W1mdD3GH3BP0yWwTUasZzfPBd9tWZq0e0qQ6b67xzvLiCqP56LPQBIstsLO+
Z+LavY7b7dzBZk39ZQ50nfQfZ1otV6Y6CApGSqHX4oQzX5qa1IGyzg+GDA9d
shuIszSuXdl0Rb0sNebn3XAdbWc+eWgdT8b+Aq289UH3jOLQ9bmRsvS1TytE
SRttPZ9gzTsrK3HxceCFNREshKcvzwl03n62DrPWcbmG/xJagirbioszo8i0
CJuqS/NWJRZEK0rMsSQCA4trAeLFWlUAS3YQIvUGWu5ixGwyZM6lPqbcJ8un
Dm8ch3aDlEure0lhOi46GwxY2OmDMVnfvHH1h7RN3Rd72P3uCsAIZzilmYcP
24Qe/6rlzusRsvLjauDadPQlXsSFlYivF6T3iW7W3ySvBOGGE/W3SIu0iztI
PjSTDZgjgL/Bj2gTyZoOVpo6EvZe50rEvX0ZIFla78GusHS+J/IVrzVCuyp4
edKafMmbetueuZoBNp+7JYXhWXrHM5QdkkaJ5o8xDU5oPFd6JXm+BBPu/LA5
fT478wtJTiFY2qPklAZsVkKMoEDTMCr74lmVBs7skF2VUgN0A9sm+M85WauK
4yVIFGUMk8L+0DfefK1wmhKjEc3GPQ442WbhunzWPNmygWxTtePxPUF3bFjQ
WBT9JUkLsMFP/9PJ61BEaoORSlCsdpTQSUVayme5Y4b4851dZVGxgohNZF3T
BhxR6/uVEr7RBjqy/wnDGF6zusQgoBQTXgroKpuGz+R0Q/YZnD3rvQcU+Rvf
Jrm6ruvyKCkeXl8IDWdW+LQtNyGLxB36EgX1EJB2wJs3MvOIjgcIYTh9uyyc
5aT+dA+m7gtMzsqwmxTUvEvlJC+WArMgCOFH9VrJncl1M4YDii4iQJgUZu5Z
o9NF2CfTbx0MFuEQV8eraTlU0ivMbeXRF1U6tI8Hesh5HUEuwEOi3ZMsaC6Y
Jofz47AjJmMkQEyeEVhaX5cWmTumZ3vyMsT+vyhT673LtPmoEnm7CEd4paUh
qg1EOI2DCnZh99ehWWLaVAL8njGx5FqdqmOr1DPsft0sAD94BXwkST3nuy/Q
hINnwLSiG5jiTQcittt4VfFf60faF5vQGNbpZ+mWWjCzsXFb4DW1rHz+3JLH
ei6pliwPHbWdKsdVfelKeaaklob1/aYxBIq4Ekjp4FiakLRkdaJ0NBMFQZ65
98EEy8DzYL+pBqPcE+IMSxQoAJIpVtuGDz2M/fyEkSEG8rMMjz0qSXXhY0L3
PGnxuIiZxTXDbfG9QjhBHFOXqgI1KcGxw3yIxySFc/Tf5Cx5byjGpts0lgU2
TOfnRvf9whh31QDld8NRkcyB8Ei6NfXr0p+8GihGjj+DwXPE1O0+TogyTNXk
/R5wcuTXUjReCTgSmrRq7bocmKR/AqeUWtQd7oWyTRyxxkTZZcF/gqfRnyTT
QP0zWwzQMv6iQFdNWEsDMkl7KR6GHbXXELi+sUNL29A9JmjlfERuCS3nPNPd
dodL4s8LAilfNCCydFCdtnEBbAU262y7t8PXPRMp6XJDPWN2wvosibUiVmIE
zCUwy84b+HfNDkbupD3FEiTwPvl8FGwWIVgZJ5WwyqxT+uIkLdQUyefH3fjH
tl8MXVWpgND4u2y/lTbq+eE4F5NL1pvwOh0QOZPkLVBXxyYVhpADi9MkCj3N
oTCbYRr0pQXYQHJSv1q1hC+kmJNVOwIbfmYxGqStk+UlvwTKG5sCleui+vmL
CBHqFZ9LiGZN5F9lp+SH4Qnn5ia9UEI9iv7PKekzQqHBjjbpjJswP5LJWGa2
HyQQzQJJNM1FlEveTl4dbWb1Pi6M+Jyz+NFxB69bX0Fzj/8Hhw1kapiksWjd
X0/cPW/rxbDJEv4FT/lAHlM6sCn5cDLNlblLPlr74KJjBFmwUKONnILooXzy
unmKKogiheDFiFU4DCAybhK9RslAiIRA2RH6k42YRzcuyyY9RtLdDi3MUPeQ
HxiJGk2P9j1QZJiCahPthb8Spo1Y+8yF65yixqSx/5VMSS7EyRYieT6GY9X+
w9I8hnUeYj8wGQJfXFGtfE6LiTI0ClW2kO+A5HyW5L27xqp/bIMCeeDXBPXo
NjvFzYssB9zIQhDVO1lZ1ujy3fRS+tyIkdjIrbgkLaDGpu5QRtUZRstgPmVo
9WVAqBXwBygUhuZ9UVYaVYFfQf0FvwX6WwryEb2KmKck+NY5TJZONuGcVYSa
fQUjy6iThM76D3NDf2BCjlvvHyiYvKkKOG6sd0pLmwbDTA4kaR+X9MjYTP1j
kq8mFbUY2nxtHMstgNa6gLRAkNtuqR+zDtsEO9CtCU+reOnb2p9WufwxkIpA
r9rJcMVe45rxpLDIvvbcsYobbVio88MQyH0W/+Ez4WLH61uaX+22MDD7hvrE
9oZVNR2GZdj7AaD32WTJpkW/a60xP8ijHJRK2epPJ7X1ylyHuQOagy0MYoKF
UsxGByVX90OgmEGsDt06IPFtBA6mMoxB53qPLCIMQXs7atCQIs35K9Of6pB3
ocm7ShC+/3EtsZI9q66GJo1ZoNBJ/K9xpsg6o3NYm9o+taQxCZKLw9e/e6Qu
WYhDdC9doKJYdgtjOopKwjNy5EzAImfS4iX5TWXt/eYGkhTXsIp/tw+HX603
y0PK7a7/tAEgP0wZKzr4dFRLvGhauEDabbdBqIfSJrp+MMjqS/4tjPQYL5Cx
G4OCbA2yfbGX3+YJwusAea1v40ek/SjzqxSxa+jsj3C3miA8R62Y6hkDx4aK
4gJnaBqTGOB0gFQgbkAVWORoalHYKfljyMgIleJajObY27zmu6n9fW0y3xLH
UYKCvoH1fI7oN/lUKtaErN8LL9AWCraY61M5TWfQRpmvmsHleAlqzhbIbuZE
n5H+WPYIqqixeqqXNLVuydU7tmFp43VpK21cQWSVDr/uJbLIAnqdYfHV1Jbz
5F+49GDdzSoOR3xoV6xrUKg5xgiDEZfN+PG5cBv3vjS2BZL5Xg0JYXOr22r7
h3yq9GXcvHuLp0sR0k8At4TNLkHrAHFJVoStSyt9iAmt8JJRUOHwIrha5q/R
qtg14WNHPkql6z3tgHi4+sVasyRuZFvBO4ncZBxSEwr7BNFhEHusIj+2xr/z
VwgDeg/H+XZRWOwkh7Ubice+JjjJDrTQhPHTwf2J+5z6yc8Hnx7PSWpbTlIJ
jYta29BLn4eP8Qm09fRYUeKz5ibO2RFNjLq6cHhWuPC20RZ4QRP5lPgis9pw
K94UJinKxoIFmcKXKcGqBSUhI7UlWX5YYySAMo1uc50cd+Xoqx0F2jwnjlhn
20pmum6R+2akQXHM5/DG316r2jPms8G7FEwk/VxWdQ7BseUHzRPRfiXBL9wz
jUy44zpgYhJ7IvrmX0ySKYxQ2lPOUfQly6kv4Dd6UA+ThzCM5Je+99DIejHm
nzu4aZbeaUzlBjLkNJ13GJeHEbwI1SdLsy/bQUTnlE/fqTTp5Am2k2S6M+R0
xYuIzRSys4dsXzif5TEa0pSmhnIZ+Orqd4lm+Qq2cE0mTT895V83rlAoL/4r
8l+92thp/6J1s5OWTsvMey2Fo33cajZlsjLh0yRDO+xxmBwFBptX2UbfZub4
Pd0pedbNFhcPHSLIc2+OApAzHlGCuyHMwNBHWSdt/vxz3omKiWMBNLOYI1Zj
LMcSKlxzNo9Ygog29U2BCcOyqsGUgWGP6mWPnqOS8YO80OUrUK84348db1kR
w0G+DV5o6nx64MmY1PE2hvw5Ni2R0Zeg1rb+9cgntDzla1YmlrXEochFkzfk
Z7++1OmXIItbuB5hojOTbi0mfjyxqJg+xXXN1EFRjdg6a4P2YWWVm1AORxMz
J+zSoK0oU1a4h1y2h7eIaBTffLDQY9SDLFwhZgz6RcvuY3n9LlcE3vHWGBnj
LqP07hUpCYPhqRBDeGsQtTLNYeyD195pEOaVbz/gMforCKJK/uv7LV8oWAPu
59zbXcwMxRW99XqxbKp22lx1gcWMiNPzp5OQCsjli2DoHYXxI+php85T+jze
wjeuw9ossBSQwoh+MWjj0VLwTnWgzf3hI/EeRhtKCiYUuf6V+fMnyTM92dI5
eiiZJvo/Te99nULOZfVYLgvDRs6LX7YL/P8yujSnGhmoH3eZFWJAFn7qwIbw
6dXaqG6j46rXHRYmDDyrD9U/qXUv2xR8rj+fHecxEEYquQt9KRV6gdMuTCAv
H2VpiEAzLban6awCyFiZIxeSZZlArfqWfn1UpJ14HudImAStuHCw/kZcniDv
DLVIEMUbw17sP1F7TYMa9CkbykE1GKqMwelNDrWcUheZ2VeVl+m1Ip18U9a0
m2kMF2B1D3k2e/StCIFYGwP62t52g/K/jx7HaxN3yKpG2Qg5kh4p9jBQrhTR
OvGuIzK60M7WUpIHOEPdjRxCrfbcH4qhyB12AjitOX/z2Yp9CY6Gr26hdiwT
ia2M3HsdSlb0dzhN2moyQWfcWFt6cqp+XjUknSqWqmSNHR7wBBxtb0pYAShy
C19+sQIQE2K5sh02baw5ebgJv3u0Sv9OY2GDCMlnSQsqOB4cUTBIFAy+CwfC
tTmJX8KKajt/ShwHJBMUIM7WgZ0tctjKq5TnPQV06WNGyETWcd4giBc8MaPZ
0fb2yY0BvGJ2BiO2fIkKd6rugragWTCUfuydaOzR3Y2ozwiEKCQjSHSycc5j
QCyLWVUctAFHuo0JBjosNPMKtPws3fNHZyhzQRysl9zAia83OJFi3DqmQq+k
2UveA0Rgr+Pa39aEUApu3VCLAQd3XzkAdkKK7YDIpjishWooys+JzAkSlQrz
ER4LI9MRjVMm+Hp5XnIr3oD6DvAxcTf+SF395SWrVdtiI84fWzcCxIuwfbwK
0+xpE50mSNM4YGjVS+2V3217jfxxO1DShFs/2oDGzNOhZ7LLBLm9ZJhxSkON
NxnihtjCqk2JSNHIP7GZ+6qWJ4lCdAvo8OEYIlsdNR+dtt0KOW9xT0Y7kNBP
2Z2MAwmeGmz5sKTYlIMZs/3XcBQeLhHFTEd8QIzJ5c3+RK+aS4JECpNZ2leN
v63vUQmFA48V9QTobvDFpUkiQKBw50vbUroIc9VBCl4hkyD5vrzbA3Lfcd78
wgAWZcgZ2xIYqYOpdgWR9TD5Djxinjxr0EJuuf4Qsljrq9wm5dlwakcZfULv
hMkmpynDn9EyCUM2J1WpB+KTF3dRDP4O0XynwNHSDGwgZzcvUPVjdgpy5EBr
DeuWHvhOPrM0L8IaMl3J2ueK9iJhqObSgx0NSQZWgnQ8+nrlwzmD3hxDLgib
yFnPovqfBT/PiVKUSdimphmjLJf8oyEivAiJi3nmPIVw1J4HYupMrKwOXw7r
bNYsRVc/xaIzAAdh/KcDDjNV1oQ3RNxSbokNtLqR9HO0tzXmCVaP7Bc9w5UL
V/hzPxcwg6Oau/k31GSRBp62tsKhUVdPq1A1rZuGQzGZbO0YLVvzPv+AarVn
3LzRrg0eZiJghrnLa4tVOvrH4FZCrXfZHx2B2K1X4hBMkewGpvLZuQZA8XdU
tF+BQvdKk2SPLq2W38BfIBrjzvksQ/LvyM8Rk4gZuhtnGGUCKBmHYmRrr+Qu
jeMGX913m7TI8DqSaQCZOEHQFMu3LokLNgLKtVCKROUj97E/EUKwk+vriiFm
cnAiO2LLlrb3EOJCYtLrZnoD5DydZSi63dvci+xIqkmgjWhpzW+MAwasXTz/
36rUlPxeYNes+HOThSVYcBXQWURgCuTd/dII9fhj8maVHd9++Ka846ultYGY
DJgWuF465kbpSG11TWsaDFqB+BqmlfTpKwDkXBx3vsIc8AFobpH5kaxULMmr
iuSY9PbxHtN/OlHO0BPN1nF9l0FBoaMf2QDQ2GSYvU/eN1k9ONj7WfdAHpGX
y/zwA+IogTcV6A05EobfJuMsYOeFVpHycSxz7LfKgUysGlZMTRZErQe9E2IQ
0mq8D7FTd8a0mOn/BfZUPsxaPucPX1sGgzGsfp39fh/B4okpMH+vqRRcECY2
OLQrDwY6gKfCML5qWZ6usUjJWpoA9VzyXLmNaIdjSBdXvzd4pFT1o2FN2l31
/cdM7XjIJfgZ+y0U8GPrxvFsUQqJOW+0wOft7oUxJVkoxjJM7tFNT4BPMJuY
oxS02lEbFIYgiImxVZc4Fc69/kCok1Iuf0qePftZmIrGacEcyCdXCvphQslr
+b5tzT4p0CNuNK9AFl0npPBX3UQ22kozwiPQ+0KnrHvdqI/XbUNpGgp7wfaX
dWmWfnUnuisxeMuoIifWbMDsQRimRoem2HxI9JOaqWpmiMb1Xno8ShRf2X9A
HMqc+PvzOC0hF6XChtb7Qokit796KoTvuq5Na8LfdAJ/h+A6bMGIijtlSJVZ
nhryWRcSCuIigqyXFzkp4sX9SyCHypz18LriVSxymxiincSQF/Vvi4vSUEvj
tebSNK6H8eX57woecwsYehtoSoS4yEgp3BU5SmmABp3Tq4FFecS6tRJqwrLf
ul61hgLfVO8bRLiUwPM4v47lIkdxliXzIg6ZeLCM/3x3rGgPyidCmNfKjWLp
qxVA78ab3INJ/sjjun/2cz5pQ1fTXpVMd0IP5cUKMlXKkIX8EYHYYJZzXOVj
JSarFecMQ7DdLdsFn17ZOj85Q0QHxS88aFxrU+SWsSh6UEHtdNE0fjUyyq2z
kJwG2O8futIH7r7Lqtsv4MAWcnjoxPy6o67vqG+U5AOsN30nkMsp0byxcEkw
lYmMRE9gCKj4ICb10eBe+BEG/iMTuP+Ozb6275PzUTTiH6C7NIKXj++uGR3r
2/A+frTBRkhsOSWpISeXTmeltq8JWt66lapvhcIYzUA0D3Yf6XHu95qaKGUI
CdyPWJyeDcUmIuLwQ1Gfd4hCOejUqpz0TCf8EuEtkkOQfKKtk1pKG6IXE/uU
JAP5upo7lbfWxZFxiTuXFqehtH7xLjdqbx1y3d17jRiOzXoEsJW+OMMbJlTg
DwfXJshcyg5DXf0PhM7zVyuIfby56pDTGpACVf6orpms5VLFpiQsw4yvrNAw
lppo3//ZsI25Y+65/rNdbU9EH5GEh7GYeSlFnaNMRB1pBwAFMUQbvcz2vsP9
1jhiVDw0O79D2+NEqd6Wnn+KivBuf6c8xvk/wncaWu/5gTeNdy/iR7g/trTT
GwkEk0xNBqWGoev6xacs6b5xbY0L7qHuqHP5lZwIqlSsbS68tVTulbE+NcrP
8eElPMQxsPHVvoqPaUigtxVUrx0DGVnwXR6EtC7ka5zLAm7kWmHJFqe+xwbt
oWTYXksAAtJt2BhPTvY/JVB1Gxp8jKgjpq0gc5aDGEx3eVzCia6p3BmwpSqc
rsFsr30RG/idAdw6Npd1gs3iI576DKs4UpPektBJoFTQ/6AniF3/q1zJXdwy
d8kEPVB5z66bW+nrQlomL/h7BD7+f7LycdHo3927xXsUuV4BKJOAHdsUnyhz
y0MEMoqcdQ15cmjAWqYltMEdTrnwTY3QrsosapPiLv7ukUoQ3Khekbv4FCyn
LIcSx3/BOwOyLaeMojIOmsizety4D1zag90Y6O5kUCAGhQ6Kqagx1cEMklJ1
a63r3afnhEZZjLJiLHeDogu1uVn9j4DpmtG36L+mVzdWLJhsgEmf64S/Mo2Z
A+w/nPsqiOXzXGREwRg9Jj73tuHBotmoyvdSUOK/uz6erPmwjdideZ3HJKZ+
vkPlzocwjNqtf0WexI9a0PJSyx4PnBqQ7CApsY2FFbLZigaeca04XcyATqWR
fyLLSmWsoy5GTnqOFsOsdV8k2cpEQ1xXlI1m8Ovz/UotrwQFid6CExcMuChh
CXMbJ7xanz6RH2dSmISoMsrYJSOh7PZ3UTeY+TYXM8EWzgv0QeVT9XLM9lzH
wgBnTR6e057zMzm4l0/NC2rdBD7MUyp/YUn1MVGkqmnT8JrIWX/J7nY61EEg
98ownt6aaFl61lckH11ST5hlFoYi1sZcUUNOyY59Ez+hnp7DUvGSgACEHKOV
+lYYeu69rNb+MeModt0BpnPHLuynohMbcisWMy0zaxRHld8Qpv2IodoQzflD
s0w9qZZwodKSSZ2FiVW0ALED3Hdo39fdCrOAGpkgRRg8sPg99wMO/aiImq/O
wmb0is5d8/wOvluj8hdss+pRtZwMchV0f9JzD3r1Vf720sczYGBgy20x9orv
RRSvm5cmGe/+yfjJ2X8BY1hDpuP9nK8AqgrF633XTun6Cp5Bjx811Dxi1C8B
BJju5xP6+IZOpt5dYjereIGO0W8z2Jfewg9vOq64EMmYA6iIUJShAyRE4+tN
pRxQYFJd9cwIgNI3JjFVMDDVZ3dUlIGWZs8UiZcrGValFBJ/wKbsH8b9BQf5
yatclHJo/68raXWXq+/buvDfwGIsbLIJyGLLVx5v6bRcSc6hpPHF7CDsFgV4
DJjWK+YNxSqkxjUaCW8HZLUmtm+aDU9i7RNbOqu9WGoS3unKDRspXLrDswfj
tpRDqYjuO4gaCM7i34Tiw/fLHI0ohtY2L8cYAB+m+IVVbVlSLDq9S9kUphLy
dryFOcF74o9cVljY+FhOMZnk5LSXes6J6LrkHHVZ1htaS7Q4CPSB5TQXXF0K
beDeNJskbVtDPXBkJrW3tAaoXojv9l5RMOnSyTEldgLaIm20c2lmGSuCoDqY
m5Fe6QraVA0uTYZaJbah8/iOE3PklAnINZHE+PlcssBm98KsFIpODiAr/+1G
qcDPRbNcVHTpaN6E6A1/TaazbBSJEVd8i5mb2nj8uEyMA9U49hhbLer5Ighf
1J5beuAWgpY4oZoZc2+3WCKr/Vta8QF2fmtzRJiO//3Unbxe4joJV2lYO2TN
NNHMrMC0rAYiZsGY/udVE62Rjmrpv6Y68tvnEkYlzZnYEMtUO8lM/ASVlhFe
92x9wnX+gM8hNJjxnj860WbANiYKA+3OfqZJrplUCpNRFIyuGizQOHZa7mVf
LXtxMCJsMpjpU9FyCcauGYFPbTgbly0/OEYN9Mw8jG3Jk0pgtXW+wujoxd/w
Jsf2GvaYi32vghet5GrUPVUf2R9fUkojYLQqr3bqGzQoBMzSha3c0sxeP3X/
Tm+oIZYQhkiLk9DhyXIa6suXX/9x5eSPBvpaRpW7J1/5cZizbni+0gzHUHsF
7/3NDb8U3AIW5euAy/LGsVv/yzvmJcBIQmU7hw8enqEdKryml/hM60BO3fvt
Suo2qZAAI5DayMW9S7PMCtGBgug2/dMznCd7N7miGnObY2jE15/em7IngfCo
vfz5mdk80bzrpUMMi+MhUGv2/93n0ihwBKKjXxrUod51iQ1P6DufLXG6HDvY
LSoHk/P6qSR9vTnqkbSu1vR5v6CL30WO0KP6CNR6BkuC1vIeV8n8Xqocckr6
PvQiXSR3kLQn/ZSSF9kMPcxCEbmDLLA9HaqYz4TJQ4n6AKSdp2JhCCevpSPU
rP6w31R5ibRiNwn2V7rcOz9W2mFummItfCGq0zrXrx0YbUf1YStsId3vw/PP
vcIUPK6bvlamq67V3p0uilu+sXV0FVbm+sisJxbHEKUECMM5PqZ0XmFQfofz
xMD5P+/LwemedqBr9vxTBlUdACG905C6gyIQER4oAGKr7zgzBpwswCZ4FKPk
DgHJ8Pin9Uu6nRECze7yHf1x4FHWAWooh4JpblnujhNZYlyQFYEeVg5ELuul
WTrs2656CZ3o2wvjz4z0jr6MWKZ+I2QQzBUQG50XwwirIq7ecRmoUFFZ432I
i6Zuj1CaxnFXA6SYkX3G7twtziWsgvX1zs5U885N+JQk5XGBBV+hCSL2mAEp
AfKNLqg4zRmAOghxbsY/7kUWF/pkMhFdcowT9UWEx+vpit8hntDP67iQuhao
Jjg30Ua2YtY5qGn5wQcHSbH4eEucL/yAC+mIYetxVzQmI96iXA1ERWzaGWoz
gR9HykmTYJ8pK1mUhDt2N/vPNOfd5zYAD/vIu/Q4m4JfOZNt9SsOzPbdLQcu
78bdmoXMUxHgeCxQL+VuySDIlf2NK12/qTmRPFAyKEK7LMcIhupC5GBt3fjT
+cyS9KUdQ8zT0d7XkejatGSZI2AIh9iSn7JS6xURucvKyTYGSUQLvSxP3eo+
pzQo5A4mq/jZJVAFA1jmRLTLl9QhXV7eSwhZljQ9CDDtPt8C8XZFvaExb+hi
unOIBPMZMY028/4XkkEre7s6HIiPetmwBtdNfEJHW1qvEE52JANHqDByaW1w
/I+X2ox93FFGhT/gqV2aVjjvJP/IhqABnpOY5zkystYQLTL3mklVm9gx/UEg
CcyRhQTlYowxJ3onjQ74qseofRzFvBL2auqENPh2mCEu013IIjAK3o//8Y3i
28qAbe1gPHY0Qrzdtgel2nObf1wl0aVqz/zAIqVmh+UBbVZC+AdrQ+lGAB4z
96u4ufnwUDw4fwKSDHFLEXLy28QHlcRpYHxIHctmo11cqijJdLC571wzsA8Z
weT6/U16WPvkkOOVZxpRsm3YANdVXZp/Bf1ZPnUOMntWAlpHXOYqsBrCOYWZ
mfTetZNmyCDc+Qs8Va07DClghV2pwAcus47yg7SPKLTY1qRwGVDvF7Om35Ha
8ielVSt0OJNQnvmmhBncrcFS9+4aRhdJOVqiMxQLlxA3VCyh/aQ3EL6uygaL
AlWe3aK8v04WUIMpoH5rUnB0iNYulc+na7KmhcLO7lcV4AC9eOKDTYBnTd7S
XVGhJliy6KUH9e4AKoDojLaRRj5wVqsLORENwi9wYIhKlPA0chVOq1lEP0fd
QiHshXYqhsVz4JEuusiL1ToOEwvutnVFWylwGRFRIrSxz0c0L8Wxfo9cDdKV
EX1nr78XK5c5Css7610m4jZlIAAdBoRs6VM5CIZmRR8ZppJrMvEzuOXTqpRv
YypplYrR2vzrMSVNOSYtAyBFlmmlyB8EOCFHvf81yx3VcMAYjQvrdnmdJjCc
e7xgOXBSv2bzydX0begitC9pFHnJuhGmzz4R98QX+PIqR48jiDIEKU1na6EK
0U7OUNGuTmJEGmwMWdbBz/YTQDQf8Yb7R6McasN17wwjeDqFS1143ynQ2lKS
doNmdD60RdCicqbZWqDPsE7Of/S90NlFQjCmMhl8Oei9m2wwDGfbjqCr4bVV
y1SgVnv+fDQ2MpQd1Y6+Sp01RZqZBVBLP7d2uuk3hdg+vAkJ6Ts7DWRiQUE+
2Y5H6P7ivSP+S8UelJn7woKlT7w1Jo2ElYzyEDeMuLqXasSmg0ORZiUgNQkZ
58099wQYpD2tlPRdJFz5nGQYfE8u6XhGRicCduuGJ+S0y8L7hZHQ8RHdHRXV
hvMOZpX6CY/RQXxZLio1qs3VGweQZhwwx8chqwRE03iCOp5Xx8qFvjCi/Op2
v7YsIeKQcOfSZ6prwHgY1HnpQx7gggw226i7Zj9yWtUhBrYHma+xozya6OnA
9vv+9ExMDGXuGeh/fJDE0dOr3pXm+9HJdOZGwT2RQFC4GPkVuQ8YApoNYfXI
y03iOKlCuSwiZGLGZdIj9tHpmN85XwpTkBZ8N/ymHvPkjlnWmnOPEb/7++UQ
dW9HDeXyY+kNxXmhYNYCTf1Tm9kpFIZ+FpncFW1wdaOVibTxDPWRoLXCQvJ9
uNydaAKunwx9oosYvkpX59YDWIhx4Qyc4TX+5y8mEnmUB8nJXNhY0FQ5NhGj
bkweE+JIFsGAYu/U1Ghstgv2N7PlOxUHfEUz6KsN7nokwqaI6PFzprrMctqL
6IdXW7sJZSBI2IUAfcWdScqzMHewexxyLGgB2w9HT1VJFBzrxxxGOvH2iiC6
incNF836x52vRtlu+3/5Xxl6NmulLnr6DZ1zIDwWBmekPCxvTWXMcvPp2I/k
pUx7K/bKJ5MNJZRBia2PLdMbKMzp+AaFsnnOf+L9thwbVJEMdI+eH5vapMEw
fPTNibPX5gGJlpxzkk/zR7tRqS3aYtyYoU2kfiYj+E37ha/cpGtQ7aFGSwP1
DFskF+dizeaH/ezslQYHFW5qZzeOVAm01LfdVw8Tc0ZCws3RP0Ne/92L9T4f
VZDzzynRgl/l1B835ytPu0natFZwl1BdZIZVnzSQMwOnimNtj7OfKptglqB2
EkNtWiqvF3uoJ3xhIeSiOfrtl7iQ2eJP3hzaOxJSeow5OL6LpOup7kLAtqMW
XZy0wEkaGcoj8EbVavu2rvdgp+084gXtRUt+bxB546h3yMcvzskPVaxE7d/g
oNqLrfKWQ8QC0W+zakni8Zm+afGPd9aXWaNFMmtAn8TEbOjOWOPrVFis1j6/
T4Sq2Y14oH3u6CmNolE46aRfPxUYmDybQzrbQXr0rCMxTkuk/kRlfvi/TqJz
9VWLy3qjBT0irdvwXmmSaYffnTc5FhAcRVK4xFyCChmhaynLO1aMoT/1KTDK
w2Uol0N3gm6YLYYTw69qsA0uGsUQR63x/KoH3FQyEgyg+0CMoIWMgxBtXggB
buLgBj/WqUUVOQyiUZJbNxFKRgnWg6UJ4a5WObA3CM17/YEiWdFw5z6Zg7Lp
tZv4LpNTHQ7l4YXTSI9h1nfdcTgIEcUKBkgmkBYyABnEEZ1z0XEq09JXtTee
OtgNPBtKuDsucwCx9CoktNoqZwNY/mqod6ofK1VsduNn0KLK5FsgdjVIaPi1
Kh36d3vG3/wMTVLGNWCIOylbx1JmtGU7ZEe8POH0S5D+15ESkMMRirQHtR98
euUpwnbQjWeUro1C5t3Kz//FfmAFZot7f1boFeXgIqWBnFEWxVl6SexBb/fm
Xzuc4JKtKccOKwfi9IQjARF9J/vYv/fRGuuJWqxR2EN8dZFu5cjHJjmelrbb
Ydu4O99RZ/qq4B47fbuTGJ35JYK0h6iQDO+8VBuKYDwguEZ5EQKy5RSrrcpy
kxzlPysN/KfIsZP5SQS/L8H3fq824UJ42z3YUQvnhZKyWYjXnWHDU6XIQj8b
gOU4q3j/ryoNq1IhaeTS7CofZA0YuKRCl0lG6wjpSYIFVvj7ifB7+mAtpvqN
MVSwfF5jRQnJx+zW6KJClVvV5GpdNtTs1R/j8e6M1CpdYfxL3uTjCDCP+4lO
o+YQk+WP3EOPBzeKquU2DXb2ZSh2SzkqluvcAYEuZavmt9e5cXmeFY5wIWeQ
ObOmBZdu5v/YLUoSkYCz35Sd4Eg9WnmaRyzQFiAGrYJ34/ZZ6homl+fhGjVh
jiYtiyMZnFnEYQ2IsImb+E5n7sZ2L+BzuEVbUfvllLnpkGsksTvuZPEkO2FI
VcYBc4aRksBqC5gkMkiOLitaRHOAAep3F+uPmy8mmSr8vOakWFuQG8PdNtIK
PCC76fq0uVLos/1yVHukYmaI7tjK1wWfojY+jb+wo11CmFYNQ65xOO2LsVXW
pHTx0dk9tfuLLpKWLG8JwR2HzKQcBsJyUPVKIK0fOpYusflIfQRKKbDUfpb0
tjXtCwGVb3QUHwsUpJ1pcW4DX9fdVBPSdsn5yLThd2ci4alFIbEIlbXgpWTK
goHLkDIl+ElH6eQkJjL5bTh0NMbV8myibtF7n1vRNRdHjVDBxJB8C7JtvqO4
qcmLH7akfMuvygcYbb+80K/H9jfZM7cgI4LVamLVKjTjB1R3ELipjAKDNvlb
4b9ePEDfORaNPP/FAeaACqgZ3VdqJWPyW3sajXahqZ4vpqKi+kl8x+10SFlt
63A5xCEKBCGDgNMvx7z+ciP2kw1CAYqWNgsZ+9UAdEuOqe/n2Oy5jy1Pc1Wr
NNzG8HJbn/uoOGO+mktUsQ59R0TDqWn7w0yqQN/eE31vVgfKVK6AfE6QpyNG
bP/ED0KS6XyU9PTJU0z0wLYZftx/vXlmic18qVHG1KcmDYrm+DW8uFjNouBn
QPglpbzCqYjSOTr7nfyxk1D9/oGn3e6UAJIqx7HwC0tS5phUB4um3Ad4jpLY
pc1+9iA7xEJ/ejsvSFj2/wkA6QLyzJSNwxz2zEgjITyTj78bdIYFh700vsz6
GuZeolmJ8B+shsOESWp9MtL9aQIYtVPrJklgjZlJNaonVtIoZuOQoKm1F0Te
5k9TDSCGTbhqoPLojS+iptvF9rVIcROTfEbtjxs9X2QNq6CXegOnhsELnpR4
urTBB67Zmxvg4U0j1AWhPMImJMovRz7l+s4Bvy6+HCv/AGaYGoCFC/vY6H3c
LmLnet+QRV5jb4S16kVT5dOKc+siICzte7hu30Wj7eX9JA4yAgOnVKy4Onjf
nyvRvxGAocL2bWBoDm5orJ3uQ3S2UF+C4afRgTNWBzbE4FXepKLW+/HhZkyU
4XRMP3LE5OhaMvcxZE0IXs3BB/TD+4iCjwNxOiSptKng1q4lD0C5MhkkWNIQ
UgPF6eSpyJbi5bTvBxywmc8GluwnvjYr85Y1J/fdE23/i9Lc6Y2ZoD1uI7Yj
jkOcgI//MIq45GY59M7KuDO4gCpRyc/afum8LNJ8SbqXJPBzoVGLDRDMujvE
V45SrwPD/lFyvHvNOkGDADfyQAebng9FiwHU/UjuwU8C6B7snkxlf/kG8Iad
JbkX+BTzzgx0BD9BqnW/htamTyAAR1mJYp4ABeVzcUPhHTX6O3Z4Erj0SIFo
z//9DbNjeC3wK+tLGQW4m03rzSSydOUa49/tNJ29lTTurOPvsJ4gEhAF7/CY
GzkQ3pHtzoAg/86hRzZxdNzb70MMrvZ1V4L9/heIOHxhu3HKA8NW+0I0hA4f
ToVFsR2XBrqgntMSB9CbZ2u4XA+IQnkjN4lft0rf9CPZxOXf8lHGYSgk96+d
r4R2phBahNXKiwMwPEFOM3pA2npahUqHGpkGSHan/9PN7YFlpm58zGNU3BE9
0oEc6EYw0YPiZyel0wUguLWiRz3eFU51auXt5BjksZuorA+Q1PolfqhGJx1/
iX7EdZC8GrfziJnYov4vXFd4gxklNgePneFrrI57wHoC/rB9dcxSF0TEuQYi
sMVUi5r7yliJ2Z78Yj2ywwS5JB8f0VlWoiWNY8sr7z83A8ZfYJkFDjSnzdG0
YfF4/cpxkY9m1LR9oYqIN1VvneU53R1sDf/OZWbHKkSoxDK4J4lMMtCdx5mZ
ysIQYsKlVG5iUCtEQKWJ7w+MM6EP4mIt1tVSEkVTQUjBiBmKTfQjBTdrCP9I
+f1LVHiE14qQm+X0UPkbAK9YpNqvHOEarXzfgpu1GuBfA93aBg++l9z46XBb
EzZu05IcRphjppFv7uD6pgSCus35+w9oL2QI+CFcwSQXrjfFayNh9DNlU0HS
fq1y6iH6U1p2/alFMhA8v5qyac0oR2Z4DQ40dmI/Y0+3XRIKytgHEB30dUS0
Q7h6DR/CyLS2ktTHMuTwJvrr8KR6zcwAyANrx2oBgbvfDtMI/1bVA7bFMJg+
Pk87VvPIyptgFSG5r3vPgITG+gbvOtGyNYgaH3KvSjix0SV9HaPGjp3cBGU9
2AUkcUO+p50aGuUG8wrLJvnQSFIVBW9YUJgmWF9UOuJoYxKfx4QBh1/j2YhY
2PFCpUbfagnQRJKZ+Up5tikNTv6ja0+Y+dxBlMHJCmC5kcB62s6sJWmyTfHY
b3Pk8vy2WmVKy0esx58ej9a3MqKyaONTJhe/kWxZieEeAvOQGzAVTW/ObIq6
lg8+vUJB2qZzwjCPf4JZy4b3JmnxHvLaYv96N1w30Am6eGA5lUgk7hDWOTGu
KGj298xNAtVQbgXSW9MaB/pWauv8D1hdvmicT0Vly7gNalY8RetNJm7EOGcb
wjN9jVuo9mCIZwLIr/+qJhkvp9zUpdtfqH66WXosgSwHwwjC4vnc1VfhPnR5
aVCURR2WbcQKu9CFawEbubTZiNqO6Y8yi1UKGB3Hd1oMmeEcGab54RX0seLk
BNHFpHFMJ35QhrFABjY/aGH+cMCsZQEKjpW4CKJfNHKnVTiIybKDDZhJvKBs
386zSIvccI9zo/h+YonCwYa9B5fgX9dm5VOjujcEONv9kaUCdNIBewWNT9Se
n4aypj9vCoyhpcuBIzlzURq62L16e99FOohiAnqvBOqWUAQMOXBTIb8qlgk3
pn2QSXUxFBycWcPXGg6v88wdUKLHbBuiyxav5FaUibXMFRzafCIoy4DFCvZJ
VWSQZDsIQDLgMVQU/0o3etWTNfWAmLuDm3x6lABRrJjZ7Ph/SJiaIVr3BADF
UzejODZ5xXQiyZSmLqJO8eVEOCu+3C94wA/hM8WdvYEKtT79GrptbswK+nT0
Yqf063NrH9kFzXJRnVvDGlEsSeErHjjgBZeyvSuG2DMNLkinmbl/ElNuY8g7
aAmZ30BmWGSBmxA3pgcdpA0b+D95lVn6vIyPaBjWV/t57ExOvug9M2qdVGVh
udMyg1YbVIZ3V2bgTIl1Jn6LKbiTxG7mAXe3fzAO84Qz7CHYhbXmysHk3g0J
tb5rylccpCgXpBPPSeQ+av6qWLOM8fslYZ0axG0Z5gjrJ87aKBhRAe1TW5+/
NBfNYcrlTyMHJq2nZrk2+AJmH9jKTCcXZpD921pudK9unN4KUOdJerGe1+te
/2nG9eGNmMvkwTkPihu/3tNrXqle2X22n4LrHXWNloN3CfzeNG2A0eV1VIIz
IFt3nGciRywCzXXNZAzl4NnFT0P/j73YhSlPu4zJUodZvRa8/9nZ3WMapJPP
hP35b167viBtwtVX45wI2nvf6AKUhEQxd24F01Vzv51PO7DEqSiUIlrn+g2F
8ERbOLhGePwwCKZK4CLmd1kA/Q1ccH4Yw4OmBosfEQeU+LSQ7gp0ID4j21dj
ulvAgByBkINCKWbQ9GMRtcc3hE23dk4isP6RdfxK+C9xlA8PF67zBJbAV0yL
Y3PkIKet5t6PnQgg8aQ3jMkKAZN66QN6kqrv8YgfLes4DnLjgbsjSSh1AXZY
zdZF6cEkfuE8i2LXKPg54dC/IhUU7qncnCgz6qXCTnwwEtkpjOYM2Wptavmn
sSk3duZoLEusy3CuWfRunRQbhddLDhqMroNAfVciW779WHENDyujZtldDcXQ
Aq6vCZUU1BPpwQkcwQ34rThX0CAC///wQViyqj1gB05c1Pr7DhVV2jpGBaS9
ULzvEAu52B+xmpcS6l+shgB560Nm4HS7ylr5hKuzAsEsLwfcPw7XzK0NnzJu
FBGH+cfxzBmpO/478y8lIiXMVf248rPohA0nSoCFGOdC7XL0vJ9a+35qXneQ
fCWafUmplabXg9rMPm8GNIE4VI9o3RRLBFF5fBODylJ6AFnpHxVSh+Pieso/
3LgfZ327ss0slrHkZhoeulOp7ozh1EpjNzvil4Rlq7Hct0EtzYH7YjqY32SV
X5sqLJJ7Hc8GpRtaP27Oazb3+x296JMo5YObBgD2tvUb440e3R/Kop4Avhdw
fq4jItyP/5zNyoZIAYAQVMyPkqa/HoIPzeXKSV0dzMjcFF0gQsL84my9iy/g
Dt85F08miDruumJyXvQ55hhy4Rx+J9yR1GRgMlOSnV58vBrk9FhnLKr+GNjv
33+bfXxw3yiGnS777gMuiYQ1eRj0UIo0VCPdv252xJKedJtkkhZAa0Gmq16Z
0gF5wZvy1b296BSC8Ofec0MCaFgStONgD4tt9ySQVZ13vakWfpamMjJcYKqk
NUeFze71nDEgM4t1jtwK/1BQJ4lnPaywZvAFghHyKjh3hAfiNM0DEsV97W65
8NBKkC5Vdbtt2CQTW9vRm8fH8glM678SgIWXoZjoYnCGJzRCYcqOj5F6/FXp
fJRza84JefAGYKPBFq5zuPMStuAiiQ9xNpkc2liS78qY0UisDRymF8O4++WH
13M1drTi9ZHSISsObgG20CBL6M4uga5kn+VQnOdTMnQs0zZcP+D6Ti7+z3A/
bzRDIlTGNnvJGwXAn4Pb7mg/MUIASIHw/KXKrw3z89Cwx/L8tzpD0YGNDc6N
HnOs8z/b61kce7LKFT/uraqlkeJtEaJQgzgHwOz5Q/hA34deSCI7UR5zfLUz
JmkrfpMRP0S2j8598pJdwlHHjEEFWmUTOBhpv1lzrkNy2LxpPZbs1AfNm6Ta
UdS8htDs4D29YiyF7b0xDgO/w/0NOQEfLHaYShdcrXfDw9MDACv2Hmtl97ZK
2neYRX1VRCjau1MasQsLy+DPbvbUagJ2lgVU5KfOmogecUoWV3Vp4rsLLOPH
mpCNiG2MMyF5+TG+wyBBxZ0joCHsyGKcjgYp89QruKkDnROE+lL4tuvjW7pD
VC84ZXd4gbUqlpkxEBuXc1QzRvVWqRUAyfFgyv9YDwjkq6SkXVWnF6xrXmEB
NA9Kjs0+bQMgs6DTJXy8birvX17ogBxdwjHa9MDhgbVSGRTEjlNyZXWsUdjO
30niweCD+KBEcjdxBufsQT87JbhUanEzG/f3iPKxVG1r0/T174OyoTPVOzty
WwZfV/X4XWGJzeN5Y55zHSQqrthlPIPOCspPJve53o9TXbKOSIojoBz+ZfDv
Z5NN2YH7cVTspjINCJrdCjqxuGqxsfeTwPLgBPasdIF/PJdBHvRh7cdK8bM6
Z1xaA4JfyS4aPBXOdGtIgFAv94PkZVovkZinlt9GDMVWKl4gTCxmWdjmzOk3
W4F3SvypQ2xvokDzl1Y4VA0pYLoeiGDJ3CKMjjARUiTR2sG4T4nUKYw+38p5
i0bjTZo/rEKUg3HHwKBLvgZzaoUi5JrnASKXsuC/kDBIiAeVmUk7HcvzU5vP
rPTXb8uYEBkLFw42yMPD1B/StFwW0kKB6Rrbk43nQ76pB38ajkUGVYzZQ4Gc
rVDGjTRPn2bf+BN5RKoEGTswXpzSI7Lja55kBJvaw4DDsNiP0JG6kjMRyOk4
wT/Sa04+lok1R+8dd5Z6feSO5zl4iwHdU69sdaHAN8MaUV4fs/GiaKWB8nLV
YCMyve1tyZu4D+wID40/5lj2U7TvVaUU3PFrBuLaPB4fufwoF/sosFrO67cj
0HMONeFfp7tMKoIojoN/oa/YNtyNGG7KD1aTQtV0Uq9nYzvcWBHQ1d8s1fDn
p1iNQcpEpv+Zr9tnUzZOVIJhmnmCHNG7Egs7WQLFmpyYfDI9knlzEPXBSLvT
Cu3mviC0hZJfl/m0Ipn+4XqZ+28Zmq3oblgTTCK3TDPIwKP5ZRcJHjR5kgCU
Mp2bzLXT6fnEyYjhIgT810L5/zNV+1VOdJ/exB8j1kaUbOfJ+MznEhNny3xN
MFwpHaG8QXdMerjv+TPOAbX7oqh9Wkr+1c2+uRWeixJhu0T+1A+wmpDS1aBj
2g0OVDrOqSzk/L2SoJ8i1w+K89DO33m8huknKL/UbRnD1p+2B4q8lSn+1s3R
wCRfLNmqCa31jfr7jvt/2Xp3ldspZ+VcfxKpuFMu4VvUpB7bPXD3iNjXhY5W
yZxHPvwLOk+bP75nydzfeJGSFSPeZz2qvimmVcq7jMZmvO5x9O7LHHJ+eIb+
aS919tjd8ZtjxtbMdOaZZHM/kQOmQlpYInrr7tSKu2Nb/Hf0kg2793J6PHih
Vq/K1bmdR3L9dgITeYir9b2vOOv0T913lZb+D+AZgNCnDxGFXfng52nqNcDh
/GMO0sb1o3RlFcKCRUheIILKaAOCVSC8zz/4iKjoNb2B2Ld1FdWZ3ZAt6AXs
31xPaFtEdQEEquL9SKmfAmw5qpqxOkoJTmAhYgwxZ3NrUVnko/NNnczoPC9T
fhaYJaSWq+qhwTaeWEKYqIQ+XCjVWMmZ1ttuSIEpiuMuYRVdOX+66N65oa+7
BGHVpooEeoJ5eJ3R2eRiyndPtvf4Ss+HulDsILun12djf2ms1xCYHkCuQSqR
ggFkQuAkqk16Xd6A+EKe2mo48VvhMs8tyzFokeLKE3JungkBlvtIF2frCz5W
DmDlOT3y4BfSb/du7VlyLP6L7dF9l+zGx6HYNmxuVBxxpXbxVNJdAFM1xYrC
Li9kNF/uVTRop0dLa2PAk8j2w7LMJ0XznXoupzjntSrB8rsHhvmiobw17wc7
bKWRx/WUbrGLZD4m7CbS0Qc9kI619hAgK/XMg/dXMg29Oegcga24BWHS8MfE
5+ZqZ1kmeLZ7+Enhqh2hz60/alHzZp/CXJSHXOoRZGOl05yFLeAT0dme3s4w
hqnkPWVrvNSbiFI+KAyygMccp+TnY1NnND63X8yHpENU+8xGerp4hloBcVy6
EJnmzbk/essfaSj16hcuWVkbz8svDozbinSEcOBcNfXSdUjwkO2MCZtuVpkR
lMNcoWs1YkdLL3NppENGdLmuEZueJxzsXXgDnUzR5EU0/gvR7v0slrsYRUjE
yMdmMJA08AZbVRDw6FBEOarw8vibQPj7CD7P0kURJpGzL7zBC5NOz8zy0hEt
qsn0QaPM82r/SSbMWK1vznHRrp3kvlrv8OZ44l1VjQOSDsSxI/pew2YuNQNf
PFDzNhYMt34AdfwnL/JVjGhlacZzG6mb+NYhuvfTZ/BMfMXmoLhJ3nlzOnoE
8s3LCL5/pkk7/hDYygr4cVJt1ZyWvFPRtQboxcx6qrp3Qx/20VH0vCPiWbtA
a6Iyh4rhKMPmqEym4dH8sLTTNvLUxCe3cJJFYYYhNHXuKpy/DZQTBPCscvIT
KhU6+8KJ0OAQF4UpWwy4+6is5/sjdS8znqyS/6+qJahDlvgHWaQezCB6r4+w
+XldNharPdQYkIkQ1/Ot5z0TZQ26JyT5Xi1Oc+ioRWrs8UFCfiB2R4/nxhku
6wYqvbn0rQjk2tV06m3dmEA0DjRZ9fqvg+HgN8yXJ8sUHsaGsl9nFOf4788e
Vekt6xjESDZ/VYVKkt50D280FPgrru8o/q31eO9rbB94DL/4RZrVhVJYH+5f
9YBBWu1h1IziVlvCCFOLRydyfb3+LynJ0vUl8UybccNjBK8a/Bi2iKYlr+Vk
t/44qnklwIaxrD+cTYb3L2+rVMqxztWMUZKAMjTxjau358Zfex7YxIOGkV8d
z7Eqrwi7CjB1/S/U8sAGiIKca1BvSoCDrHeZSwqMKIg4LcypQgyB563TWFwd
/YNvhyORfqPkVM53/lPANAZWOAeXnCBAltRAEuxCxxEhkogHNxtsGspeIj9f
4HXDfUEK9oBg7KO2CghLV6NPsnC6bj/G/DRFeEf1somL9ZDX+FFvgcMszWVK
JJMDVzLSgl7ACv9FhZKEsWgdJaMQDS5pGakeyfJ5morjUwWcG3I1Sr/+9bKQ
f9FyXlLZYZuUsguuQ8rF/fqzWlmsxQf1n7EydfrXWrvYhFnp0QK72Zr8cG3U
vL3i3YVWgGCUC1gUEUvMNp0rkxWiez33ajedfmdAwcU6K/k8hnr9lp/lsBcM
SrVrkPBGP2kbavcMMlzdj9Aq6XffwytLHt7MQjKpiQCHF48M+g3MdZkmfl2C
EIdT9NavfZ5Eb5qFoKOeRXmYhOFwgp2EEKq3/vTF3bB7wQf3zxkcFXymFB9F
td+ofI+yT0ADaSEdXAZEXfQ/IvHY1a4TlE7qyhkt1Jlwj/vvPyLvDF6UxpVl
5RciQYhQV81hBRC2SGwf5E9qj/jWJ4hshn/aaLz3E8cSZuwoJgsjdz48JYxX
VjpSmUKTsrYDODRtfbFn/oXcA0XefLiugBKG6zgbArPl5eS1p8JyBDW1bUui
9ay1Lc42mcv2ugj2xolQAA4LjZU5Mg0VrQk12u5yKcyEoAUjWITUCF5HH9pV
XQFj9zl4QpnNG6sE+dNxW/ao84H8y2PEUzsbJlmeBcvTnZpbdoHn+5tAfdMq
1jsixEgkl+B7pdazOCXoRGPuGj9A7XoP51onhXGqJMQcfMWVen/s9cWwNpZX
lJCtWnF1hhZWhKU9K6nEuI6Qzp8VU9FIlY3y+LWZTn1DOhY98tE3m2h5ZKhP
CYtPEsIFZih4KMJTP/9iQi8yGeW7eIpPxk5qJpOiOsViC0rTvOsruivbd6EL
rBvLj5fB5y4a3MXBgKbtAmZFN0omILpZWY1MsGhu+jEqKq1YmpfEmmzUvWny
nLfJKjpZGaCBTy71zjrwbQOoT3GA3UHoTQXZGS+cxdpVn3jHGL1/sPYPUq4s
kKW0Ip6Y/C/jKcpxAZ5G3LfdDyt/h9DfrkywFwqKXwsTRMIuybcUABRpK+ZF
cZlaSnOYqUR7/yIgvwv5tDfm+jtROkYtamJFwEXZOq07bycahs5pJ8obFW3v
HZoHD3RsRiKJsCIF8VyMhS2xjH9urzX9mwzpiHAg8VzQs/aBS2TUUyqjtb/k
9LaEwfOOqvoebcFYvqc5oeNFlQlHbueh27BuzyssDPNFetlksLiYMeNKfbzT
uj/HbB5np++CEFR6PUa/6HRcDz9iSfUehz1SpoN4gCEPXRxpXGeAFhtCJBiS
QZ5Iv4y116H6M4uth7BkunMdofzWfyKBoDBWSZqj28EdTk5zijbC89ppNIFZ
1oga5tE0+Wl88EwnJF92UHOF52092fJhtpUJDPgbECxf1YaUjmp/T7/g4DHF
kxWMJE8I3lcABeTfp6VaoIymqI79LWlZukorjJkMYvfVhm66NIpZS3y+Jcrn
LCxacnabMFBpi4SUK7i98ThYmcg2artse3e5zBtK+pClalfbkf2VrIejnVWK
8IESQ3CCSV+WX6eymNHiwsHrkpn0sXemSzDFvZncoi92zYXrjH0bb243KlS+
9w5tUOEeieLJ/9iMRxrmwOmxlkZgVk8g7AAhd/61uePjWpRb6i/Rj7hOslFA
H+Cf2XUKUJ1/CqrEQ+4BI5veA+0YHAQoGPa1rIKK3+LSYXMj0/Ajdvw++Bzn
aIlAaVGPEfUudZXIBgVKZqk7dGOwrKVqhCh1PSISTS2txDJtjohENTT64LzJ
aFoO2iwbMsBxCXa73oOVM141+kLRrPlgMT/FBjxs9+Anw6oCLoriQ5EB30XJ
PCOSVONkf1CF5grOaeIdkOw+tF0auDltVJeRTTwM3m/uWe8BSBFanetMQ1fX
RAuQ0poK/e7I7TYkc6BkMniQMw7TqMzMnupOa5EXGGLO5osM2do4Sedmgral
lGahh45gHDY3dSJBRnEnmhhxESD61LAtDN11/TIE0I/Ts4c2XHaH27WKpYfb
wvXq/Sbd6AUkx7RoPYndYKIXWOdQHjZEY3OkL/wGdhC6ZnjcsFneqKSAZDUT
YV5L2IFIUp1fLQ6XS1uBX8nqTw8O3P+SsgAz8+3bffXELddvKoxsHZZTtKVb
G33RTAaSmsD4XZJI1xzpvCxUC6zepxSPw+ikmZgphtpq1GTCLR4hnmkGev7U
cKVWXFFWl2eJdR21hPqVCpG6lKyarcol/3vW++YPwGdZBYM8FaRg+w/wbUGc
JNm4dYsCHCq8/Ox13GFnupdHloW86QFWwZ74bLWNQSjZAd9Ici9MJWI1ip+4
DvNpYIOF7biMztsx/E9KLZJDMNQnB4n/uOp6C9BY2nsPC9G2Pb2fgDK5trZo
opYmdPBBBA5qq7868lW7I9BH/+4AfBi4vfGmV+XuF+f88smaMti3rMrK4Wmy
+nCTcqbkTf1UW4Be/MeuobYPeNiyeMLUG74j8XAurgYmHSZ/6hHlFXsz+TL4
5msk5zdGfY0FguOYUHYVxQIKs/kR8A9WQP6po8XVrYKh96CK09jl8h4v2Rgn
Nr4bLWWHWb4CRO9vFsttTMu7JDAfJd/MeqOF/ysDsKgXCCq9jR2chN/Dig1x
p35hrLii3h3vMYrl7nanlY2k1Op0AYmslrcb4/iTp3GWJPdX7f03yDkeR5im
cvK2dcr5PtOREwDhulKbjaWSX1aNRz3MWrmoCVV5l7HXxysSIfzXqjGhiZ7q
X5EwZ9WJwkvwEUJhev6MB+TZ2KlNNKVPEpx5mTuyLl0yCqGw1u3leo0CRWVH
yKhymfos80j0pJ8icyLlACSproT1hi9pnJvoTsZaTyA6WCSlAhCRbf7y8G72
ajJklHCTdGcHno0jiKvjjBf5YeX/B4Ky4ZTjbY8NKIbcCWwC8ZnlDVHM/gic
198rAbpMS1Q5D5Szb285Nz/Lqd9ejOwmLpRpV9Yslj6+u5MgjWjMNkOTYVdn
YFkQKER/TwB4u5UohpvHC0XAK8odYMZYglvpjaMXic0PiDL0lU1o7FwW95s4
1pcB0GOLHS90T79nlFDtjCvVFXY7GLLV+rK1x3xNA7N9+n2BUGf+pId31kTg
n1ZT84wATrLM33/RSE6ro7o3Y4SYqvjW1JgOdRsoboDVXu1tgXrCfMlMx63W
3/Ms4Zaokx9/FT4REnsYiWwIhwtMsAjyZ28jgLTiwP/zDRi4a9Zrp+xqZK5F
fcCtWlveWXtzhbO1o/ol+El0mpkpIdZdbii8lPP54eeFOXvNk9NvVAcat7y5
/oboDiC9ws5zic+cc3YU+FORe5dDrhBqWJAe1RVmpYn6pJSevwC4epdieDCU
ZRf4j9x5wPQaoVYFqa0qNdt6U282oyQytoeBgZE1dJzNpIoCf96s+8vuKIHr
r+pGVUM4hwV07SMoxNuotGReX+qbkyufT1n2fWifcGIHeHlIls4gnu0xtaCU
notB8mNItEUcrmjuqa6uB54paUkS55cduO0/ldTnjfY4ygPCd6sYTafKafoB
/b6nYxRlOzdNSBbaw3N0BbjZii2YNWefcRbP0P4zbEufzI61H/bSKIJl58nK
y71vcc45q6YDl3D8X4ps0Rk+8K5lETa8aTa+HAUch40K4Gb/Y4MvNGxf2gj6
b5wd14OYio5COFzqtTYotp7r4HsduGkDNF2H9MalNcoW8KtALiWfNMP3F4Bp
DiXdXybw4mSwzTA1s0rCk6awR+EvUfepiPwlwAd7nO+2aYNvbBs1Iv22qkop
GlRFfXuY9igAPSesvgvO2/GHtiEo3P0A2w2GnGM0nl2Us0n0v4p5qSHq9vRU
Crwkz5pEkSVjMiDM/qEUWZ4sQT60FVD1FBLj7kfezjr7yMSdwq0607rXHGsR
YciZSyR2z7fj3Mpr8DvdF1XFykGz+HFex5e6ndep/T+b4zdZksfqJdPJmsj5
3+9zy1FrOwFv2OyS//5ve+KNXKRXKuZ9uoThhV9X/2OgAJeq5GfbQkXodxbY
7QmMpXqftT0mdodcd7iE9NRDl7GE0ZDKSOd1rzyszKyjVOwRV5QH42RnwbjS
PYkLZeK4d/g8aYcwy/H9jSGHefADv1+ohfIlVVEKaedq1JvyzWTMjHJVrDiS
6QRbRQ48z7CE+fROyLB9a2AOiarcD9GUlJ06l5oXcQF3XOhIqv4GFxwY3FbR
fBmCUvaQTyDmT3kcO9/BZ+HIdjDAjNBQyyp3cktfRVjSWF+IQnyfhOqWRyuo
gjja1yCqXZQlPsBSGoe4gIb69M92fw+lUHaDCp8XwioOCE7TiidkA5hbds7z
qV9gElweil9SKAPVR1g5UEJEAoszDmAeeffkX1tSFFRkm8a4eQ5p0AH9Ottg
mjWdVc1ewax3JJzCmp7B1fNEHjPe8w5xG7tbVuH6Y8OI+2Ftm0tbKhaHe5AA
1pwudH/DJvy8iOcy1YvGCGKh2VC2+pE6DyUZQ7AA6X5KcWhsTC/d1aV+m2+j
x8uw9cxU2G+Q1/KL9Zd/vb8MAzXxJMu3sOYOwLRlge+r3qy/QB6mdmk9x/O1
Z8Y9cFddQij04vYkvkaYQruzcjycHwm6xMeVoHAkFyv9CGPcRTlFHiHoW5fU
f+Rll8is4Hvv2cRT3WuKBSuS9/kOCnL45XXZgg7+MvB/NL+YTtraWeiYxdNr
7SpJaFjddndXl7zcVNVfqNWzJs2m4gLmlWaRQg/dQWmQC2XnwaMIKO1Ug+35
CHoiHQ98gJwET77FDiCm6dOfr1Slze6UTEF/0ZaBwJ6BeegGBCqimzrxZev+
e9X5WvWM1Rs3Zzcpq8U2z2xgRxANwjzQfKe/K96tlCHLH3EX2GxoGrYvhB4s
1bms8ZgeINw8CVYgQQdTv1DlqzGQmU6EmjZ3lpQgPwLXXqnQR4dtoF7QOWgD
3GkFKKAekZXdr9TVjrQVrcG0vbDA8gWG+1F1ZxDy8cXoSvwbSbTQ9gQNkbyG
pvd+azUAVuPJqszM1cWT5RieHyoJXNNXof2BbNg2NJ7Ot+p9+ITAy88sR89x
cbqYc92X+4eX57kO6n0nD7DzBIFfIurJMf+1kPaEqCxxYDPVGkcmK35lk03m
Tew/C7s3FpbWurnv7Z3wLz8pqb4uCGl0IKWz/FmVw+bfQ2riXEvhxvvKCp4F
45YAFfOFapen6oGzeqdmVRcwJ4fBEwKCapi+TWIBNvTlExCVJfHmzYYwy/Ut
Nfh0ZF2BObG8imtNmxfCQf+zIJIf7nL2L2UUZ/wu0+zBOIP+/GYGv7of49ms
zwdEGvZOcSKMiizQ87SVWU4ny5uFNMUF6n04iyh+jehyBkuJYF7NNHzNcRZw
vD7H/pTAXu7lckqfZp5xiSfaxKiQ+fDjY947O1Y90VSQHk4WOdrPVLZ2ojLt
oRu7eOExOuvyUUaMldEczQyE4jCNrTLMH6UKW2SD4HZCFlvLU4uD1QplwWbl
iup3Gxxq4LME/T1lGxmE5MdNqiHf2TIf/ZwNIPuwYnNr0A3tv5uDdFz/JaJY
z1gSzCNw8urmnUxbWbPODdmCGjpQp860Ko/qaD6pwoU6AKAQt29i924QI6cT
W44EjngFnc+92Cpg2Ff0r9Tr3L9/SiJbUl9wDma6HujzGsePd6Fjjm4umnLr
3K3fNjA9uI8mpVXnpNKbDNX8pkxEkW6bW4WVKaDn0tLyCQme0gHKYYNw9FYl
kVML2yHHVJFlzN4cuXaciABRPbA027P0Srb3JyDoXfui1CE8SQYFPDI/rgYm
NwyG5phfkWeP32OLHK0QdehQdSff+hoZrBhb1yRZcwcwoL3gbXge+GxNdylN
lBIl7yBAoCvRhvfkmjDtzR4HJMicYNAqOzjT67J8S3AbEuK9jwgwC76tGf5A
8OdlolYTfu/skc8lDranvW3SbxoT7WZUiCq8g4r0ShQEWMIxU4ZTG/e34X+I
MLm7vFhu/tyq8ZJJY+vZKLI1mRo6WLASPYAAj/4Jlf06tp2WR4hZEo9JcNXy
h7VuWSxetlyNbNkAnI1j4O0jeoxeHOR2prF9TQSCD2fRPFqeEjWnOaY7KJKp
fj8idAPKJ35qB6pOCrdK2uuodzR0vUjRoFCMQ4B7afvYO/e75ErwadIAKNYQ
h8PsOcwiShZP6oPXYVcAyvSnz8i6LtAACu//uusnXbJMhsfuFLjqJFlrUypi
oZa0AE5K2oODdcgclLnE4A1HfZtbUvZ0mFUiHZJs8JbL/xCP4c3NfqW5XnDq
/kj+J+n4gIdniJ+fwijFCeF8QK1ar2Vu+jrjzFEtEhh+A8kd0HjpYFSnvAP0
J1/8vUo2WCyyzTf2kbHGq6qPaH+v97GceP+k//GpGoSIuD2CCKhjUG354ZAW
+KSOq1/0bI0MgwuMw9MuKNtuhbTCvvEtLJqXcghtr6xJEualxHlgtPD+zj6T
fmuCnfhN/qCsQiRwGO83ee5n/4wtZ06xAwu/9kiJNMlpAkLeKRXuXILct7DN
H/OzSyT43FscfkmUFqTMiB0bt4SOBC7s4i2G/yisiNueD4+RgS0BRJOGUOn2
sBsyUQOmK1fqQdVOuuF1SSW+pTn+gFu4xCQBWPOBibSbfliaaOUsGky+vvmY
3LgJ2GlQ5p5WamdOgOyJ84bLS/4ejQpI/t9IigXSK7naTNXZzYJYvv4COWHN
WRYhHQqmcs90XxL28KBkW+2dQ0QDKAL2kemzKlQQmP148ukGDflvcRPRlNCX
4cvoxn4Fs/dmIY1i44fDua7HdbXsbze105gR8+VoY9Nqo+siu291Mg+GXX1l
eHrHkVqi4dIDDfId0p+l6S1Ll2qNbSySfHXkRQVx4CtyOajf1BxO/D+wM2uR
LJHzMH8FNkW0AMl+11xWyPAWodbDzajFsK5YfCX29S/w0p7EpMq/pIUvzus3
w6HdPUQE9QTnvhGJiPOZw8Eg5Rb6I8u4usFHjHG7yMtnQ2JoN5TPIx9iTG8/
7eTq3jahby7yIa9vRepYjpncGNX7jQJ5oPpIELybJiUwSiaB8lWXBTaXuvBs
JPGyi80a/jpBeJ+tksBpd8mt/aijNThHbOs6O3z88FvCY/hFluYs5EJan2xT
cJ4kk3H0V2gnaugAhGk+2EX1WtFBc2z8gKYpmdimApQ7Q9wEXAUWj4MU2qbd
iSZeY9eHIYOQ743hcDJAHSjUhYgf9ZGUaoI1By994xzixve2MLlMADnMlhEW
d5O6k5fnMygmJv5Q7hVD09OxFvTTSBX5pnz6RGxUWtuLEVkxPZla6oB8EuL6
d2uHgayFrSeFrTioy5EPP/5hSzTzUa8aFdrz0IVlIzA23dY0Rtja0h3dDd8T
P63naToHynrDR1oDzwgiAp8tmG/Y3bOUq7uj1PQ3SQ8fiTH6uZabqQPlPqEF
uZzggI+gcHdI2g676r0xoOLbUzmcUhjg2823J2cjTriD4qUaZEqwh4Vmt7fW
IKxJ5TofcvS32kKKZPbs/jY9cObV40joLfPHcX/5TpQyGB9EA5bju0X54fLk
SSnSsUi9EmCZq46aBtJk+2B6mFFPQBTuvSiQDj44nPnICmeIYYeGVZr2yk22
OMFVrf1LhBtv+5/soX2yNebLNxc/6ZahoZv7aMsR8dHQ4cADlLBJTZ5XA+jl
zCzDvJyPsumi/cSP6Pq+KcVSiL5shkHmAHALjnayjup9BVdwBiExfIvC+OIU
2mFQOKZqZImAxfT8iyo3EotNOJwQGCyJ+BDhgbGOht3RudvohXM6BuRKn7rz
kwLbpyPHUqhHh+y2yMg1wioyP2RzCrOoFvQHHVWFJtDTNspzSchZP5VjkHUV
4GGoieU1IFyUeSsvPcg/i0Iqi/gAi/i3HzgZfgGdgg4lnXn6nPIfhnrEk92C
O7FIuXpChSFykJDji9+v5Ngy5tq5qUYMQEvAgQAFsKj+M3Mb6IktDaJVn1bq
eckovkBrZpDp5rDbVY64LzfRGw3RZbIT9UF2r1SwL3pc3t0fN2mG9jTFsaCh
54OQ0Lm8heHeOHEbDWMCugzfKhO0Myvky2YOSh4H4s3ezDTlTIz7qeYxMEBI
55DgGFFShzXh8UVvNrA9dka0uKrbVevVPr9T4lGvfnvTCsHHho1NtBUWURS8
hzsK4sBW/qCu58Wr9twEeGVR5h97NJNFpCnQayy7qELM5Oc83N9sq7OXonF7
68Za9TwZdgaw7vQOuzelIZ+UJRcQf+hNxanDMhS0RsqkXUc6p2qb95yPWarS
cTg0+Pf1NWTaNU5oMgaJIZH6HcSEnc33yuyaU8P6Snfzv2mBve4PUSAUYY0s
2T8mBoECGPJlNR4PK7KrgvLS6ZqYYVt7NTOJDGMc75KuptEyrnbvAAtwU6ad
BDctM7JAeHfewZ1lzidp+Q8ky/YnyTyXfGr1LzCIkmw48NkOOZ33Ca142j/N
Ifrbyp+dOZGd9E5dm0s7uXUPsJaY3sJGnD6lLQ3Wb5IPukJioZn6JDnSUQ91
kakMy5Js0OJAnwdDYL7r1BNlMPR0nMdHxsOOljSU3Gozk+VsWOg88Tp8sQLm
MNv0WFRU+XxV+VNI65zG90gfZN8PZQOrVxLyDc3aC5pqja6TUUwSaOUNcTzf
Z1+VKUxNA+gBXzW1BvqC/c/TZ4yEZclc4+UjiEzEtIkoflC2BPVvo1CICTsm
0Q5msKQQ3/P+Ov3mPrr9MY3mh1gP1Qcb0vz+GL5KkJc9juV3i1mjqwxxlWPx
SQ+t+/mnH3C3LC/ACapdL9vN4ptg8fxbmqRZ3ituLhkVngCHp6umYsjcLGWg
3v7lAmLmwSKXD57qk9QiwbK6joC6Xtq8KxY2vpDhfoJb4ahPZpONoKIuSKhq
8zA9C7FNvwtxehwn6LPo8rKpyYicXpU8a7fSR5IfMRKPzyjB6TKtkGvDoGFG
dbXtgaKw7aM1DhrW5cKgodT/L3ptwVLoYY6NsmB4QKtGAIWE6+raYNQ0Jt9P
3y2l6rdSQe13PfThHNw9+pKWRXQd5peMTtaaFIVD/gJ1kZYqpNLvCNXBFJNo
8KUWgzJe3XPsed4B/vwpMfKQqcJuySgE8J10fUZkRE+S1/NU7gNSNlS0n979
SC0/XFr/gP9sXF7ZeBlG4Cnv9zuh8F6QsbIIK78ADM73yQ/rZ2zOSgeO5ONy
+h+U2Ij04l47Tc4y/JOn+ioYvssyrxb3RiF4vmH8qSXHjuBbyI/d8QciCGdK
3vjVQGUSM4U+CBGzNglPfiMVps1kV7awKcAPRhFpfCI38N5r160lp6vM/RR2
v4CZXlLQ1pXb3fW9Apre5RIyO/V3K2T/wug/u5Szq8mevQnc3G6rBKtUAgAW
nAZbSfIeNvQSzRCxJ1Io9H6hHZKB4J9ywG5X5Yl1hSR1uwsTE6twPI7mirwd
IiX1JzkfMBF6WWAAkXCX4WfLH0lwLVXeVO5O6E+DnR0Kt1+KUFxvm6j/oJ7x
pW25OLOBLhHYRQwyFlwVGGth1qWZj0Hray31kADu196UUDFbfj0ubUYWb9+V
LAkua6JEIBYmjLb450M5dGhmDZPCeSFH9pVocb/J+h/jbeo3a03f/Is/Z9bY
oVG5QJuwMCfdMNKWaCv/HIGC3uyowE9qow/bQo51q74ILnzpY9XLKE7Twku2
sI2Q3ae+KfrpLDlybV5gF97bXA1J0t5kqGDGNFSCtb1Brhb6KR1TyYdj8WXB
C4kgiXoWmu1nOZ145ru2v/Ed0LTAIIe67S8sgsN7QdvrH+c12e8opZz5yGBg
QJPvPAoSKAlBJsPnHSVRKYDm9u2QiGHaATHU6LSe9e6iNjC3oPUrR34Q2SEf
j/NFVBY9TI5JfanPsk9T8d9BJCVZmMV2LMLh2VSQg09OmKjY4McBass3Ykh+
N5G5CWXuOetuJfMK1ElF/81U8kMnX3MfzupO8xNrU6mrDU85nPGWb8cpRX02
wn4am2KOqpzFtZ/nidkDPLUKbx9XGJ0j6YIZ8HFCPq6mNvIxwW91D/o47G+r
9OUYZa8xBclO6fTn+KqIYGlky8KTOcpOvaEjV8BuA4tcvjHahBT7ycvGLCe7
wkg6O0KycTpvHfiyuZMxD/h1R5rv6WloHSCA6R6ZE2LxJZrhodIQBc4lMCYS
iubGDsc473WPyvHXuj6y8eaFeugGr/QtMb7IgJE30buDWX8sHEWGJCJt7WVl
AGuK+z+q9t9zusKhl+SGYN2wZekU7bu/KA1kOVqtmbuofP7xoxcHoZMJFsDv
Ji7MtD3kiM5kvFeHILFH/A9cNzvwnZUoAALRJ3dSCrzLOznCb9snCfp3xcGp
I5tsUZu16ECusaMhExRXOs5r7GZZfK+jVdsWXnSQ+loZ/afC7tyLNWhEi5rA
AxSxRlWusnNBH/+aiksVTLVmgGUuPTkDMPJAhpyytwxJ8QlPuvnhNdWufBee
JPqDANoqf7rjN/NuJR1odSLnaY/IuQh10lceW6M9rDGi1aCIrz3D+5gHnHhS
YZDxc3rWs4Op6s/wVUo92bGbcR5VKyu0HhSrrkzfy/Gs27AcsZssVXRffAMs
KBsOsNw5JqayqrB98R5EVmdgFD9kR5Kf9XDcacIHqqHWPSvrOqSzVlgWB8PB
ktI/fWt9gX7tU+CyKUGlYnNgpsV/BfoOw4KkjfELuxSPwWHfS7fkIJNyCn6d
sfTWVgKnbv9i7yFfNwTRQbKZ1oWogqbaZMx1PNLH6q9WsXdcslRaUmD4+34E
2kPocSWy3bPF8NpJXrpZW9ZHNvhrTgsqBOUpqccpM+vFPVU6/+O430trjGCp
Wv0OcRN3xPUgoqb35eY3IXd9gwpUqycaFtiUKx4VQUuEBQw5VCGUQ74L1K0s
83HCyMKzHOLhuAFcqSyEVh83OiiPCK0vN5w0Zv73bItuDB89DT3GNMXLLzSM
OxdUeZMorTALs5XNPI/Bti5ncduIGJms4qbBMhMWEzWagfuFVuTjA22Ie4xc
YL+Keep31VCI3kLDCeO2OyGteYNJ5tcBi7oTEGs30qaP1V5ryNzzVuDNRW6K
vqN1FfLIBJNKDbOntInHWFa2R8K1k2cICk+wDNQ0gq6dPMcXsTnkqhdYEebD
9QywDR/I2AqLVgwel8MoCkUWyRCVd5VS8Z7A3KYjJ3P5bEwoalxKa8GYvO+G
sJyHNSp+8zj1/U/J3d4ro98NzjNCiUJasPZI/TGrIc9OFbWEgQwMw3ajConf
zDvWC/HuwRS5HVEFI8iC9Y2TkAyRKS11TdHCEWo+di5Q4UV5w7mReGAwL7N4
hNqxUOFYfsy/elfv2Mmnyxa3xGzKV5DDF/+ZWZ9lec56eb9+lYrHYIFPGlcF
/FYOSZJFmxbv8CjExVq7zX98LYGoD9SOAQuEV5ZOUdK3Ej1993h7ZHNzTMUf
hr2fcO+Xw4Xkd+SwsXqs6jL/pQCkx8p+h7j6zdbnvhxOMVjHZTd7SCYQUYBD
n/wPqr1Qz0+XtIFOxgx2CjK9SvVnUtobV9d2v7AedArr1Tih17+Oa7dVDYzs
d3ZyVgJeHQZgkmw3glsqmN6ma/nvCexpa4yzLVAu7ErrjBhLPAJ3bTcitrvg
ID1G2TsFIpuusPskgMeruq9A6mPZgBchYAhB6Ne4XxzUSz7BZd5IHPS0lLYW
jyN69Se0nAvgk3VHfgBn3yYR/TXae2KxgxuolyRZ6IOic2fgvM+/2DvBK3BS
gFTQHgMzYtQ0JulaG6mN3oq4JesWzjHU1pUeM2Rw19To5jAAuoip52Y2uJIW
tNp1aDU0gl9D18eN3G64mpXgGfWQREuTcSFoNt9w3fNkEZ+J9LIrzMib6Umt
m1NNP9NospWx/QwspzxOOT7OTHiVdeilW0Lvm6rkGnbXMZxNg8C8lOPKCQzN
3IFCGFTdtbcbASiBxpAp/n7LgB29KXCJo7ZG822VRbkhG+fCdub1h+n8w3lO
nC6keWfe0vS0rv8U2aiJBDtRiAcN559klnlmTe5YwSfgT51DKezZTcGDmsa4
vIA+FaS4DOMBZznitt1ggzrAwf3rrL4cmmnHovqz4+h6eBKi2zvKADZX6Ydi
ZlwoBUmmwXKPez1BbeLgaryML74INd6DwCnD8xS/u5J5bORqE9FrMltOnyZu
0UrJOkhXStfqRN6nVmtPFb/jPpLeWILhyJeF+fW1Y3f6+PJc5UGTN5MJIjOz
RF9eob+Dw5s73JyOaN7SVP/ciTnr2gSQFSnsjv+hdoz2yc9ohAHWiuqOONJB
Vub3quY4t3PY+BtIvuVGsogDAVxcBb6eKG9YZ6QWwmf3RxRt9HJF1eFYgsnO
sA0w5+xEwPNzvzXbCTl0gEYtE1zrmoqtGlStjJ1wlrbW45Er03ccrS1QLPzG
23qW8lGpv4w1xddBMeGl/b2Jq2CFqNLGIfOLh9wv+yyukfMS7eHQ9zXeYnOb
8nJ3FcEqmoZnNxVOfWFoF89MBIhBxqz4FS2UiSHr1ev5U019Xgl+gMNYroHZ
NGO2kxUX+qKxC2IuAg9jK2N5V9s2gQYWgyyoNZkA1FNcPszeqebk4+k+6zLN
pqNhES1qQbHtTQT3uWjhjAC2aegZJVKJlJnnydGXD6uLtmDU+HFqZpteZoYG
7F56guL0N7o3gm6YMPEmU4LVOOqVbTF63y8YuJPWOTuW4iW+q1UNFBQFvAHr
OQJvO2i4sDirY9kdweh3ok4to3eVS/FSbElY7sIAEbYcoHGNuY1C8u8Kzxxo
amkGeVv2BbVEhl20mj7pyM0VhyGlaPRNs09d1mRU04cHyEsXq9iNDkatcCAp
gAi+cKzzhzVLhdL2cuI30wNJ64Uk/hOH03HIN6f6xEMxegHaqO0Dx/CwlxGl
Zpjz+QJlzyDC5og6vmnbzF91KHKoa+lQY/L51IzUFNQi9kbcpbH4H0J8WX8r
jxarmY9/GPfLDpLHzINUJCOVCXgt0nUWNm1IhW/aeMr2GGxK5c4mPeedcthf
fAy49B4k0OqWyBARGvY/3l82XjrUitsLnG9PzVrIdSctWeW5lDZEDDPGhz3Q
KcK+39TvaDgCk9iF+ztZadlIbagOoF960cUvjd2T01kVFTXZrh8V02RoWWJc
7dW6yKchhJ0Fp1kIwc71X7NKgPqLRpn9TmzIsEktVOjGN+44wjJfaO9cZ9W+
e5mtkjW3Lb9Ild5rhfBs66Bc5Eh9Vhb54KDV/wNFFOJIjIbjLYL2hKPNvCIh
4T/W/kPE5iGM1Ad4jE0EvygmCy3/HIFWV1vVaDPRwO/8mqPr8W9BTbwP/txM
kZHcXekasYIwQEHPrZ+MqoDDDgiT0QXDA85g/FBUIXWvEVLnHDbWGqiRB9vn
a2sA8wp/1cxyHPeGNVQMwtf+YDD398j0NHmfpgxM239C6T35jGZrjtg85pvc
H4Vf4WOFDeT00X4hcB6iVYalX9DXryyGug8UZa5VdWNcfym9W/eTXkah+Xkd
uvASDsKHsHlYaiUfehsCE9lqML4Q28PTr3cu1+ONkSMQzYEnk18TiljKATXZ
rSHdUxz9Vha4lHbOtz0LfEO9CH++LPngf9A3u5FblNeRFDWDlf55JQJLR0Iu
XTzvmM7r0E+m8VpQK7DKf3q91jvrxVurO2n5UZTcixnWrSEZfqKGs1dqBfmb
Tt6wXzmDJBUzWQCGjXi2U5FtWGj6CBXk+boH1gYuGoUQRFCu4GzP6n9bdW22
10ovycazCjaYP/l3S3QFWA3btIf4gVK4XtSOkYbh8XQivICI+OwUiTAfSTxC
400Qy6KRODmi6r9cXevikt5GWaP+5t14Rhw7P+M7X+NNvXkFE8UXcsXxSknS
oQi3AwmDU+E9obsgFrfJYzxM0mu8dlDyNE5HYfgmZCHqwB4W/Ybq/7BDS88w
kc9Ami9P+7ENeQF/yTAlLJoxRyrlR8bhIbw3DyTyUrTQk9XymYPyLHF3qaD6
yxJz3B7kNHtpB5jdnIJkM2rBWS7xSgrBXuia+FQwSbD6xA3Sg4kX+55/AHFh
zE3KBYDOQzKcaPhqyfdL8hATRVx+9uJrhOUH4ZGhYYjX0ZM5lVFqXbBbuo93
3c9SyPYOFJUIw1Orw2ZDAgEe8+A/vn8XfqrD4a85TeagJ/xS7Ef1dOXNV6f1
URNKvLoVFOiwVgXuj/ipHR6D4ilhO6TZqt53fgYVcGEkMOTmEcPfedVjthrO
dglt4f2OQZ/AvivIoqXyK+lufMKr2tIRjLTgnjkgkpIMz3BgLspERdPbo1oV
Gn6GtCxuOQcdTxEWR2uyTOor11tMoGODgxX2tfpud7G8FlRAU/ohTdRBFLjh
6eYf5IH2MiQTCGvbMc25Hl4F5GUviAwc2TWBGoGhmauxABo1VC97zGJT7gSq
SW12TErSyoDUu0U0fUZdukw3MDm9fwRoa/lBfjoF1DX3+N5hv0LoPpgNSERD
zSabSONpmGQwj8PBUXZfv3Ug9u6VNPVq+m06zOqT81GjzLG5Bvr/neKyi6fj
Zyr741/WEfTRrLlxlkwWrJWMy2LUm5DUE2qA0jw06rkcSmqVvS4IVfkZdbSk
kF0cfP7f8dL0EVQnMtLk2IXoGuywa3D/Y4Rbs52wowIjJgEvkDB0V+DL1R2M
gkoSoqOJSA2mJRBLNYDn0pCgr1uoZG7E5Ka1qhpTWYYGKVfnReSNJ/ulDNrW
AGu+/qLyMwdUSX494fXljFlX6UpR5Ir3hPyHtO463MEiEhE4p9df7wdXN1mC
LOv4HCPOHQGEoyCfHIW+cO/vq83cq402D4YJfmPBKhUiNitESxLmPvF8HHAz
cpw+m0p5ynOrL2TzoaqqM55+X09huBmBmEV+2qmVtGO1iIOSYoq8byHkazz6
Y1DPjZvYdh2hPfR+GgKZCA6h6+fuEIiV/pjNbxRlaMOLpOb6fncc4eogfWSR
JJ16i/wAiCYJ5NIWbPk126cvnwcZ0l/ZQe0KwvOCvoVUqAipw+27Lhz6OUJj
MjdRGdvJ52/mJC6ALRPWPCLlsFeaTHOVNHFB4gx6lXkt6dNJOlHF5l5jhfTw
MA2sz2djzoNUka2cQWLIOsIY5G8NuvlWIjznnKgITv1hVtX+ubM8cgNpMs1I
tWAP/YFjyBDPQJo5HbfZ9xLmOtrn2LumVFPBPlF8D+FnmHXQkJvndZ75XnWz
33VNyscIqlVRBNg5A007R3Oi66XJz6ln8iErfQL7afqclH5BSFikBjEueM4H
9/iYwnKDNn7UvsMrYJo56+ocHzeISn8TLPqAU87fWYMW7mrgdQuck3/aNuSQ
FsSwglaaIgygWQ9rYJUbt7jx/e/8TVyOOQTia+5QIvJwJkkvxwgJ80HYP01F
bvHAob45TgW2eNvhuEWQomODuEmKYG9AKw8YlfkEeVYAGot5HSYtHR0x628j
4PQHe5Isn5ZNarym6fYgZgD+Jc0nWsiTD+59tjdNNgL4GnfmSZElnfLjaO46
WrrsHG/+cs8hY9qeiWyB1SStQ4ivz+neF8w06hy56HrquKfJdUvbi5+nT6tw
yFCmWfgStZsZj7kAUA3aQXICco48wqTJBTH1KqvrLt0mS7tgdGmBBfxJ18hg
eb5TVqezZECI6B6YMne+FJuyNuYjx2MMicUM4EPFqB9F+naifpWJmK8Ptn7F
AV+JFsaeU+BUxolXKudcqBHyJsfyTgCXVshW3I9ouaJ09T4Lt/HVRPphuYwf
xw361gcmmSS0Dm+VYSm64nAnDalKayxxeF1ZpOVWuudjs9BxhlZ3NPKP55pm
u4RO8QluqBtmjMRunjDrgQmQEFThXcdukppAs6nk0CoDiAUUIUw+6kRLupnU
Q9cp0XqJUm2XWMKfh0+W2P1Iesg0u7Dzg0wszvRRwXLG6wZXitVIeD4w+tIn
/J5WNvHP1Kois3J//ZLSll4egekzXHQMQt+/wIaReUUrVjvlwg8LxTE9PtBa
5SUXSe7HCU/J4HS650htZMJXK+r4KCC7Q3oPgjPg50N/bd/pkrc/zsw1YvWL
TWn1wuWh9O1ZWuqphs+m43fcmKqfyoQNFLSU6VB+pGJl+8jPfG0CM3fgV9lx
ElOoSRExfU8rbdy7O+EJFRmGEr7iQiWr+Wjb+ahblt/3OCKCsEerZDLk/Y41
T0joP83U2/OpKcmhIsCmydWEzNgdLaAhaoTPFIBdkeYC/OngdqDl5cIKHeJC
G88DKw1wxiINyJdgl87URhsQmms6d2EfjHHAu9cXQAhLSY3Rojpt4Pm7NE8g
ot61Vsa6PtxiBJB0nWZQVYtc4mb3TLoazNYkShj0J3RuxWUVgAWiaaqUDucg
Byc4NVcsiOvnYuVpl1AxKjAvaKCgoI1Krc2tNxCkKzGnJ6aswumfA47IcewT
85jauFc95edtgLuJojXmkx1j8FkFV/AYeLHgZLhGh/tNvAK8NJ0WWfAATzFP
20fXo55LS3XcKhTWPnzK73nTwO/dO3qsQ1DdvrdfDjp4/ZfNuBCPwFL/aOVF
DStwY8ymCunRCvOQAPYYNIRXh7+spTxPYVvi6aKAMAFIf3Y0oBwDzvtxIwMF
2kxU3++vJu5ohuQcEVyftLwgfimRzUiCkIBKZxPFWByFtT4epTbDTIvsY4uc
Ln4f9SiZOqPE9yL1rFs8oM04PtheA8O7XqJSNPNiPmWN7k8u3cetb3YTQRBY
QsKXUi96LSaT0N4WLrivM6DbaBu7qUDRUWpOsZ45M9eSS1Nnw/h0uTUPd2a8
XpjcDJTR0gC9FlkCJm0i1TiiF9hd9K92mGqvYZdsjTciVZr/gpEaJ4Xt9JkR
wnRvyG/T09UY5Q5xztSeT9wnnl4VoKxrU36WFiTKi/5uHC6FyINOq4DuVNCx
iy/UqCvVbSlCrqeYy5gIkWBTNLXD/Fx6GpAuzIcEod6UL4IUrDNN53hPFWP9
8aH3QpDaGwAAPK0iKNkvLzz9J+sh6EpiM6WXaz60boG0QC2BbGp8bbPTv5yK
XWUdbY5trjZJrYeSIAgwVQJdfLeBczGv492VxNG+RvsJ2blzhE/qzsLDeqPE
SU31HwRXIMdHu05lfnvW0Rd7n7Srx9yviX0/yk2jRyzEG+YqKZyCbNfGO+GQ
5ji0APRkVaI2yoXDyXS4tt+RoUrEuEdmMH1mUr8sJOxbCNW4UlWl7B9YEa0p
9hzwWYbts4C8WfyVeaIfVD2HlJb49VtOhPRtbuQWlcYhbJhbIci6bmggvt98
lLg5WtkxQ3/owkiMJ1NfWL+isAzTM0j2DUuwxwu4EY1PYi+iotBMyeN5BOfO
wGWH2ZGLTyFLUq9gjlVtxpQmegxRl2dEXLE5Z0B9ETMXMzIdJDaqgUMy1cew
dwmlTe3NxA549oSpOVA8b/O9unkogZ2djO9jTVk6pmB7OZudN+yQTfod+RwL
tl4cGQADrvgxKKs7UX/THYC1uqd3Q76hKo0GNbp4AMa0X5NzK1Rg2CR+u8OO
mXMsnMm0oyEfIJcAzJpnAj+Atc1mer9dGXwRMV8lexwAXBHWQ+DPzV8YyIWA
gR/9RU3bABxLFrjXWOdCAoeXJj8ZALCBpp65JCTItx5peRLsZ9dPK8EttXpl
CphRV8HAKb6y10QNRRuxC6MFpvpfb4dgUewgXgUX6pfrwjm/nco8tb4Qf1Pb
B97cphi8d75daxbL8IS/7BUZeWKanHxqNVyRE9qlbuxHAWdQQYyj5G6qO5gz
XEi5yfMouFZe5dclOcEhKle0rQML7+DgQqVnpdceqEfeLZ1NQ6fosTAHzRPP
MchjMu9oSfNosgzSfrjgb/ZFQOekKlrOhEX6fbAqlgJglge0bGNsv2R5vpmb
fOGBAGKZx5o3Ej01YtQS55EnLJdhNprqsX7AyIY3PYtKY0UQb8DzLYmU8FwL
S35W4/8/T+qeRxFn2xxOnBJT4elDLH7B/gTmd8tHUC7eLQ6Trku+aB5nLZ5m
AcKa947uwsksx41qM6Mum5yM8pUyORbzGvabzTKNGW878ZPgM8UXN6bFdKH+
buaHK5+RLe4cRtIsZp6id3aHyomLZgCJK1qmGNWukH9u/ot6k2iwuFCV6Wkj
X9h9OdMYmKhdwKTsW8a9VAJGh8xr7Wj0Vhha7qfFR1WuefYLDN9BukshNZat
R2UXbBm7ksFJZmBhegoZ0EOAi5c/km9PMRmXPZzM4FgDaQjhPg8Wjn5I+PcF
HPFDQIsHizfZP7b6uEC2S3ZMtvV8jOrJhJUswG5UkPKPCaAtk3vw2iF/AcGt
PXtC4MXiOPckfbdANWDl5irYTqmJkY5gBBp/+RIMH0oahORm3VRJY0fmSURa
/qdOKijaN/ACE9rj84xa08V0ca/F02FZ5yP+Rivr6puRi6xM3XX2aT/v1pjX
OmP6rTQQ5wHzDUgoZRhUuI0Bx3MUH6Pd75K718hfDCyS8mc62LC3Y8YPP7z6
AaQDRbT1XJSrPVOqXFzHR/bl7HQ0pInEwxW8a8T7FFl36+r65uivKl0BxDSK
lLNs5O8jFh+HdvZhNjCn/eUqsAzIDTxzy2TVPzTYbYEUaB1JpHt62cptW2Nv
T1RZVSagecq2E8QbkduMn4E42oN/Kq9ZRCUsAxHIzU0Ii7yZX1bPYsTYPLjI
XXrz62gqHP11YEk1A2GJ1bYA/OfUkVudQKQ+MEV9cKTifqezIO9CA3gxjcA9
WavRB6pTZDB3CINj6Nacv1a+GwLtH0Edd5oUTElHkOAe+AthOdMRLiw7BvxG
u2QPkDcA5cEAmLuxIh6bJ2JX1F7Ja8NZnVbXsWogLMBufBYxvW2IlfHqYLj2
Fyvlh9akXRmpmUA3lU/s9Mpt4sNojo1iTTR4wwxUWkBbT1tIiUQM29HNYD89
EH1rW7/kqIctcWvB8gE2XktbuA4dom6McrUUIhOFnc+0vxr5xv+GDoDYL698
jV+wk00oICdmXNuN7kkohLW8rFFRoN67rrInlgwp1Hv6C5jhPnVxwSWT99Yx
ZDaQBr/1SE7Sp1v4ih7jIhDyIwI4LPPR/6GDXoEo38SZqdfPYxaNuAOMbuut
MCAu5SN23TL03SiiVvcZkPlPgC767uUT+A/2hkcOMZnLg5taGFG7oMo3fwRb
BD+rN/0JArVnBlkbI2yUMJcP1tGjywLYiHgHajCa+51ZOIfnW3YsF9ozavJM
rJ60jPoLAo5lYhJUqAXRMWsR2dck4BSrV5bPpx9k6UQ54nhgWOC2IeI3fWpw
qbxhyzk6WFvFXHFnhamSOKcZnTF9x39ad+31QOk+CYJyPGbExI1ItalCuqwP
9gI/txX627UvKI+RUU1yHx/oWR1GNMGtdjIR1CKnQBiQmpUv+qm2JKFJozj8
STacy5dy3TeK25XA4LjC5lk7X4gcPKvlQzmDZpe4HZvpCzxIchBd/G9xHjop
WTHEcwY/3kjRpMpITuUPcSk70Ca80k+p8IHr/rJRuGVhyzBj083CeeEWGbCH
gRi8zWUUrJSOYQ/NlqTCXJcZfZCl1e9dWHflW4KTyLV4csANey852l18bsq7
rQRPc2Yu1xZ/ZNqhFIli0JjVOwmM/55xiYB8bv5Cjy0rjJhHXsjs2nFboawM
WhFfoRMkdnQ/DQ4M+OTLoGknlHeKFvyN4cyFsg+eI63YYwLHW12x0Fnvng3p
iI38uNnU/+eW8+ecqy6RbKntpdrcq03M8/e4Q94HlmKctYA8OHMqvJ7bp3wK
5Y0AewMVvkFAiAvhguK7pg9BtsjviKUfEfHWuJhQcDNGWUZuOPVnGUaVmr3G
S/bBVAt2iLEOUzB5MPTzD+UIlmyrYu7mDmq6nnB5t+AHnD5nbp+AR6OmDVNs
SqnzA1xXX9dnL7E/I20cTDq7dhQx+yMv/tevVzZ+pDNp7ftb5NBn

`pragma protect end_protected
