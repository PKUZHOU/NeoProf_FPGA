// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
RQGM7NUOFfwq7MDWRwDTERAorTyzzNjRivqdkZ3lH4yku/YH3g0EtYu9Wows
zVioAjvfP526pwGV1JeSmT8ppo3a8kCVrf2ZIwVtULKsePos/722E627+jCQ
KBZiVMAvUq/M/cb3DoWFeGShad4hEcOtpiwwiG3E9dGVvZLcYwmEcDpnuBlk
Nraf0GvDyKP9/7F7bf457zxKAhn7PwM1dmkTtpt/IKstMG9qCxMJDKjpO84Y
WUnKt/T54ZepOCU4uIFTqXpiKtOoOnQROL6XqP5z3jHN2O/OoXIO40+83dN+
8m1XCcvOh+ey5D7DlS5ZIhawQBJgmRx6nNMFTTu9zg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
RDeRbGZU2P/pBKKMMv2cAjevR2jlyBhlcsLZonwDZLxAShe2CCfEmxEzKcOL
KyEvC8jpJ9Hiw1mUAQHNx7HD7XQSEd27NwSWHWSFj8IWSHrqLm+yH48ACP7c
JVEu4uBR1sHWw+/lEI2sJ35k+XGShji7CJuimk7HckauhcC0srUovZiZCd8G
feQrCLCaJw2GLnvqQXaZF+RKGbyy1Rh7gwRLdJqBx2ZaaZWFql324ad6dRXO
syB2OI8OELWLLEIlxNEeCZETg7dg3DDW2ygjoyrwRf8uhG5SY3cPr+0PsWqB
Pwdukw2BjsXWvpkHePMpE73HgN1v+NprxTZTYEFwTg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
azoecsLsEyaMGXEWYescmUTZmfwgocK+ciGi4TYEL51ddptQbMZ141bVaull
QmFjFLkY/piMCqB5kFaeAHP7GpZ8C4lQlG1o8nUIu74IhWtyZVLUGy8V+g+Y
4Jd148qINY2V7pdZMgUre1DAnFAoT3ukJ7BUkt343E2bg7pINA9jObVAayI9
UdN9nyLhn9S0YIOJ2mn0ofyni0i3y18uFr9jLHBokW/lxb7JIxAVI3hKW+W0
jwS9WgYJ1VrAXJGSyrmZc2h7odjbmy3xBCjvHPf8NsmddqN5uZEbJHoATmTH
ymp1zyFVe1eUoNnxK654yULegk0oX4h8tMD8LwL6lQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
II2C9eawAYjp6tXAduJnE+eylzShBdqrYD2LplUNAQuOs6o2xHaF7OctN9Rw
AQ+IOa+mrGf1lf3qJRE8w4JFOWgGhcWh7yMpryjN5e8HWZVPf5taCTQ8d77a
oL2SMy9ou45U3Fl/jedybMgZGmMb8obcJoPoAhwG05D9SHyFyaM=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Z3SQxtfiUZobUSf+91nw7eNyoc7JErYkryThS1dXryVL0dYTa8/b4LJ8C+kK
uactLnfz8qR+BhFsntBn//z6SIBH6fsclQHz9bfZc7q4ZcpCL6gi1dNPbUJR
cJxalEy1hS0t6aC9NIfaTCgKYLWVQQ4X2ZG5DlIAJQ5OfzHYj17Qb4fL9na3
EmrpbZC6lQpjK9gVB89uITtctb3rxKf1EzufwC+lKAYBcP2X+bPQ9k+R1LMV
uuiSkfGQ5pLitrXwlbVJsP6sAHBx/BuZVv+G4WyjZjcQqnOSkA0XeMhgVGSW
xoRN/JgnT+bfJH5w0ogQFjPVs9ao5ks9VNFb0oSYiJSq2Ezsj9tRH5gxmsg9
Y63fAkAZ8rYfT8HmAAaZH8O90uVODr3vsETqoQCkP0o1B4OTqkATMj39p/fj
JJen/K/txqwIO7oeR1tvHNoysqByC7nJ2P5ov1oyT7/ZVzwzRoHXG/0XcrxE
6cBNPgktg8ogm1juQL9b4DurR/Blul11


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
SpukWQxgAAVa/lQU7117dLQFvJ6j3Dt+8avzgBPZjMoYrm+b9J6AWPgplnhl
/gI948k9/I4O6hps5r7Lz162eAclundaA+8I+lRa7OFvzeJJLZ+GENNw5JzR
8p5GotX6WlyrDe91QQh/NRDLm8dg43AOHf7ni9+4WJtrjR6coK4=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
QWWloMoWjn+Bu+KITW3bY00vftW9/DB7//yPEkyelEck5FnEoWC8VRl/NBaa
unffORxU4zdU2gGwCz1Fg+ObPU41mWNUpCca+mrNfDDlFZdXtRvOFKbYpNoQ
jTYAaiupXIYaYCKKftaKB60cxVdrf9eUOFMl8NTyZG1KOcw8gAw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 91936)
`pragma protect data_block
Fus4wmueNqsucGQw7UHKOHxUmXdx00kmWf15Em26jr2YYNO7bVqal+gLrAIJ
tFdYSo3ZJN+M+5bSjr2ULdQWEoL4votrlBiUMqcE20hwKcgjj/91GSH1mEmk
FS9WQaFzek3jia6Y4GR/wxvL/V1qmlumcO/+J81ol8zzlD2GlCpNwGFacaWI
rPj4fNjC44IkHsYu+noFv7PokwwVMkxO8kKtB9/AKzQsh4lLU4Jn+oM3KF3U
71vV3rQugEImfpaq+VIpNAn28Dq+CLGylayq8nHFZf1tr2Bqq+xv6l8I1bQE
Hwqz4WZEgHh/a0ptPiKTYcuVBUMR2qMebMdJJ5O7FeVOLtwoIDJE7CDqKKl3
0877xMLdrr582tsPUiuuiuWBIhcsGWvhZCavW+jsuRzORb95v4pbsu6kJVdr
l+H2cHdqLgFcU+c0Mk6pwfMmbDxxFNzlWWMXyV3Yjmj3gg9qHcdASX8bWDN3
+K7RhxknA2aK6F+TJj/7LjvptdudCPJS1kD1DHCunkPXgcDKNcdtduWxr7/y
1373baEeri5PwyWO4YOOPmdMlTS3IbQQtUI098tlFe8QtXjo9PMf6UtVl17H
nfma0zu7hvMp0suC4yFouLyw9OtbPXdF6refCwocUdA1+C5FX/Cf/DyqG6M3
gpX70YIfKIhukNF846PBW1kVuPykDPm6EiByFbkY7E07+jtvxDm+xOGV6kXp
gJ/NlzkvN/18Weki5yvW8eiCa0mboMVMLyt808+cpN+wjxXTfGDGibhol82f
0hVlbVBGjtg1xTyZWV50xD01s5rO1WL4+Wa1zBP3Gsho/yR8V8fK45pY0j32
7zM2iVKc6EoYlLJ4Rm0UDF9YBBRXChfyitqu0lzlw8XoA93rVlAes6DOM8vw
yVhYewaiuiv21DuxBrjrVEPEam8NECkdbzolGYVj9x4BqiwfBW2bQ/kQxDUy
DLXlULPxodC/ljF+mGnixkqXKMpjlRudoWqnE08+AN84ssv0tDXG2nfFLmoh
CL9kJWj6d9PN0GZEGTeDVhX5yZWSxNfix6pl/Z/w5Xk1cIkyq7/yI5g+qzmx
KZp92NJgVAXTiqcYJMjznqrO04AO2Ct9AY8pFdZ49eqJuFQTfMXLbTtJXFaW
5rHPPwnG4196ZEL5DLMgE31pVnBN24kj2sc9unEUnR2lZDeq2giS6Sm//VA9
PU2QgVaGN/500leYtsHys+LQWv2yk78cUxkkv80BD0UUtpmLH8txScuqKjER
6oRjT9op+uAWe/iJIl5FKYxgERMqIeUi+8VEUou0YbgB87IalmCpGsswXkA/
4r/86UeGTH7rzYZLnaQBY/lcQOljn2qFp4rmcuYF+Yt7KvLl0lVWyhmVk7tA
h9wCqfWEQpMs7FlDfeHHUv+ORWbjL4RDx0KFzUWDG05rc16vcoDaauDdw9CA
kEXtB1U6IGpvKK6tuiirfafn83pj6oE2cmMrJ+xywUzXWnLEWW341qGGqma+
xng5gvS7nmhuYg3go1NUQqjn7UO8XFzfUB7vP25j5xt8JckCMn+sCsAALvGZ
dOfT2izTSCSmS+sjWtLKM4/VAxVHcolmNQjMkT/iCaewNqZffxJhb1SIkLIG
aqZ0LzZ/A7mltHjYlACAlDYsb2jUH4N9xfgCszwRIrLTpxrZuzlEzMUFMVLb
8mWdrpf8A7gbKcpKvHe3TVXt7nx/DP/+zYaqVovvzIP7dyN0SIDmxfVbEhY0
oDrqyYmYMqSy5PO30z00gKZqMbSBZZgk6lyxoZgCD/r7Le2wVScMuS7kqdfU
df5+jjx8v39CdwA+SaFsiadBxCykXsVvfbpAC068i1oEdCgDILmkfs7jGqE/
ayQXFHWOC5PbdVZHje7M9MuX0QVFHU6Su3QWqXNDS5J8YSLMt5MGPYPj55ho
bjt5Jk0ls4OzvAsVhPTVyE0U/1SCWSfq1gk6Hn9RLBdQxn6ebt67UmwTTSYi
cMCRof+hO4NQKYIgeNXOXFxpkJl59nVxlf54jMSjcc7+QCssWgvc08/uvoBf
xTSitJpcV+gIxQXzC2ceR8xVSvJibGcNOBRD1J84lkfEPbmjOTRotg4gTe06
zW7kT3a9JygaI2LsSFSK5sqaiw+mkM4yNy7OYMBIIiH+1bfsIvSeJxrKr8kJ
AjixW1o46LWtcC/yBWLuJ2PEs1nLRQHlsdxhyTnEcrtidDQjj2hoEzmKpoxl
F24E/qv/vfGfk7tai43FKvGQay2Q5iCL8F6Awu5/POWu4FmLZToh2fHyALg/
LWtBbE7aqlOADe4WDC7cqgq9WEErOQi5EzSolGR8SbZRsO1q3qjn2NEt8Rk5
wgI8r5f2+Cxa7UfdpARMuiNVfKQkzUxITmRSSMOV8BofjfUF532c3icAm5wd
PfNQTqwlGmTjugUUnLtf5VCsz/IcypHEO/4zhXCEIit7yr5jMrLxjRU4Gw9n
2cc6ajGL0+qljnfakBzUOoisrQMvUM92ZPbWLkKiJGgZCc/haaBD94Ikki6q
JHRGZiXVFVKTsY1udWQYshbpamPp2G6sZmkmGGgc9/oT2yU1loPBqoCjHUK1
FTHreHluR6L2v0khbfeph7Fs1X1ZMGGFTy0dnOKhr5Oat81WiXeXalaSnu6i
LBGwJED8y8lTNJsQ+pg5g1RRna+Q3FF7bqOoKs4Zc5T+1AyX3z8TA+r5nOt+
AmN6VFHeUfP7DdgIHNcAArwlAC2d9v1wdGYf7urE7TWFuJrXrFEQmKY8VKl3
haA/Sx7Qmyhge7VrIeXHxLFMVZr2VtGNxO0naYde/gRa0b2Zmo1pux1R759e
77e9cc1cISLqFEXqTvT4+XIMLI9vtNlIbKX39PLgrxgDODzHzV8RcThSrM6K
ErLe0+93Oh3Rcwb5aYsfjadXM52uGIH/KEN9Fq7bGvbC2bJUoAd8v1udztn0
P3iaDDcrZaqjAaZ8XxiJ1WO/G83lJS583x9E286VEYABgG6xFzBXT2CjDhaf
1jz1JKRPluNiG5f8dfS8Rc4Z2IzrszN1bmxE+SIDnP12964wBBj2mIBzDG9a
S2On1jI0Ccp671Mlr/CkI7MD3OSeqNfNCbS5M59im2irKhqD8sy28614VnGb
7H2ikZzik/FG6nIOHDOvunuGoh+R9UaEVqF0Lj5pt1KJpJ0t7eeLMT0CcbQG
cPdUdrTNSK3K55fpAhjfnYKIY2MpET5Ka3qwvBilVPcjYD66xDjqmI+Sbx3H
Lf2A31563jKjoGWlbtpRkFV8Agv4j7xMFkCWu94osFkTDn50w5FQzvCF+T+K
vGMZkByJcEgwT72Ve/UYvz6AVRtHUZfBJog4OzRTG/+16uJw7OXRDawrnx8A
fpHBTgJeu2nNrkiIokw8EFYvTleQVMMmTxYLKwvsENFZ1E/EU/T8dVifH9de
cSuW/UhHxO03xzGtESC0pZHdfAFye2D5EbAc+iSKWzxqzy93jOEzrmQNWm3E
3Jwg0/+YXtAtbqX+2vVVcqA8w/ii3Yp7eRvnfLAazR+4e7BP7qB5S4uy/EVt
GLmvTqV99LQAs2vTP9yckX/AdugdAQzWRpU20N8Dy1vgLAawQpk5egO3POcX
Z+CGUcQ8k5UAAWBFhDpe00ueEaRzsOY7aRLR0H7OC8D7/M0x434HsW5ZkGHW
7Guu6HTCnH0B2AyEDwmU0O/tztyqUSJoaJfs7hhSYjO97JTABQ3fTj3VFwSM
SbQMctpFp+VqDimtbZifWGeB6BEIQMUwKv4jlAd2lRWsaOGwYqs6TfO86F6Y
tcEFPzQZTZNIehQIACgKLHTVUt753WmkC6yqPXlV482vVQRe+uIRtwoeVbaF
lxaJfX9cPM8+TdIbCBDoH0me10pho5nqVJ3mCK5kyhOmD1Tkx4ihtLGsduX/
95CCKGiRXROQ4z5XH+sZto4lHcy8qFWlruE5NO3sEfKW84CLVWnQv2D+D6MI
VrVyIDsDs5My4sEdxWQNqTtJ77Ksp7Mf8EZXx0dGHiOEcmZUWenvP6wsZG6F
bgNiiuO/lRT3Qymwgl+341w5uMznXwnIB62L2aBj2EWAMKX7h8nroC1teF2B
TEPJi7X6XpioIyI9pxR27MKYri7LU9WZxYgLcdWFQUFS2q9MKHmI36zkaUN5
YC4K4zTokEcFZRWJ0yhbDDdVcJn604xx0PFcNtzN0wpWrAR5zKA+sT71PweQ
EA7We+Cb52lhgnMRLemW9wWf5qYudHNjdqV8EOtGyXS6S4ECVSurwrEavVqk
yqz+fXM0AJa9uQgQfW4lAvMkc23CqsxBofD52cWyO1yZotaZuj+IvF+gThbF
De3gCwcOiaD8Adzgs2FD9tFhvhun2dC37UaeQ5/WmzEBjI1kOrst1snxX/Mc
2jWPivblKlS/TdQ8WSPcuhFN3dLDvPgY5cGFO/pD15LQ0f/kt2tlYBZykghd
9fYF2GuJ97ZlKcAZ8l8jioTG0+lZTBcg1yx63c2Epy3M98RfQrch/Rj7s+du
UhMHADcHZ1kApR+xkcAdet4Hi4N0zueX8HjJZPqTK0WCgQRePVxWQIEGLusj
LF/lRdRi+0vdGAvXBypeA0EbSEVipnoR3eXoGF01HZzNuGi5D/pu1MGP6v9M
WwLoZ6+qcUPf5yePPzjqFrToLDpRSMtQwrt0/cbpPmxED5h/4XeTmMGMgENy
Gx7OTuAHdU6s0rkDeOjDtndF2imwZRJYFUuhxfiZqkGx/2mqcXvAelub1j6g
XlEu5e1oNPw2lAhNY4NXC1r0/T2eYqCfo3ATTV/ZTh18zlOqXjPTQ6yBMxyV
y2/HGtiuA5+Cgs4IgBBJiELUHM4N0g7uwpLcacS/b+KUsA6uzzNkUlK1P4JA
tHeaux3M7UHu/FO8aXoLMbWU++8XXezwJOaCnS2GiHGdRMsW7I3ub06gK58K
RBL7tzBnKJFz6D+J3tkR0+qmMILKcQRAMmqEnyzy3o9esj0oHpc/sSXz5Qhk
THdqQrhX7KYdppULrL3mcUAJz0bEFjxVJYF7lNUOO4cx2wGaRtyE1B0/wx//
GdUjQreT20kUtBxM0j9dkVDhKXB0qVYX0uYRv5pfWNi2xztxBCZ5cr2bMRbX
VFbMLg3e7MukAi/YKY5oG2lN4w3Ys+G2I9KtpnLurNzSCRZIpP9FYmpy/wCs
n47Ab5/czUNlHfcqvopwiDWA4V/Ty0kLRPYIcVf8Lt4MuFe9C2VvNtwQhTuC
3C37rrIiJf3CQWRWuyF4dIolCvLUIltsNC096hHruX2esLM8lDkeqxrkYSko
1pM3xMK8Bqp/p6xHWeUA5PdJW1ykkySV70R6qMnjPnwtfh/8MS/7DyoYGH3d
mmMzwuhINs+jIgVtff3oNeTVB+vjri5nlIAu/+Ydw/GqYCJjMM/MTU+xchpC
FvDN6O10Icg2DfO83m1Ay/kPNNVlrWEi+90WWtq8Am1V1Akf21vJuUlLiFR5
PDzAtwA1a1SIqbzHQBX6HkLHJ3RBWlU3F/QCfPxaDdE2R8mR/yfgZlEO5lbu
WB1+6rsMWz483k1mkLx9GVpo9iNzQrkELeZinX0vd+GdeDJ5UjRWshx5fQxh
MD1ztFwsANLNa4YXLZ4O05gI7rLhC5m6fONixeLLpqmefQ0euz4xhi74HSOb
5vAavnChhQWf00x8oOZBsZk2/3NI6DQOt/M2DhSzOKuWhevYLpm9eBGzz905
fIu4c1lMSlSSoz/gVzlj848/W9ccgDZj99tcqAWmNQ8J312YaJXcmifurEJv
6pHvFDoUceyLGkFEFqLlTPOVRAN+lCxBgIw1Y86KEZRwhTJKVP66iTpEASSx
ckQvQr3t1uDKvCw6sOCehBC/gHeYEnuTdYfe5gvWiLqFQvcagZ8FrLuTK7f+
ukp/eq7wUM2B9ShKB8E8bOZj8Qh4hVl6XXT9vP5FaMvukFcEDyqB5oah6PjV
qbJtkvoglZKdjDlzAZPpkIUQl7s572H7D2G9gTdsrj2gWWMCx48AB+lHeYp5
/qVTEY7612Tv6KWTkGzUiNFGdxo4benz0tGOiRWlCy/JwEy9KAQZJvUJtmHf
OAUicc3f+sTCdbLdEqX15/phJLgt/AJx+/mWXhCn5BOhxE64KuOD0eKgVLLz
JoC0DGGQawOH5mNofEKV2NIE5lKvx7xPKmyamYosHFhkO29A+jXqQfhI8fgQ
PW7NesGyGnwwNWMxCXcvbU4OVLABYMrjl6sAb1lbiD2e9x6z5Q6o92NcfUXB
gAcy1pH1O2s1yAgpFGmUvZG40tuN1cfNRpq7kJ4JkMyDER4jlmC8pKN/0D/c
jHFO0BOs+BO5G6BS+Uv6kuw1gA3B3JHDu1l+078wH5Ut8jrmZI+5AYrY500j
yPSrYlwvBxUKSxF5oFPINL41/9soqAW2aTZDVEVce/ANSOVnuWtQSAaPXSER
cUbd2eK/wYevrS7ZsOyAkgUcdXc2i6ZGuCf8y9Uvro+O1dMZq2gLWToCUgpw
fvDasgfk2HvE2bfGiHXqSu7VzEqwcF97QT5LxFwRsAt0uGMflSuSglp9rdet
5u5iZbUPLUSEDT4dar05411XaHlU8m/UPIqRU5OE+znL7JPNSF+7zBKCQjWJ
ERABc0b4xanjHt8tO8mtiOZ/DfY/QI5+3lBS7UI+TgXTpZf//dRqcHGo2PBw
ATzSbMYSdm0XxNwtvb9OBbuXTFYNSWyUZCZm90OE3tLTAFDtUNCXL7S6twcF
R7d1fgzets17ZqCv7oTKo/0gFxxp/X1K47sl6By4vUUFhuxaY/uUSPC45ZD4
5UxSKem8d4zf1RukxlSomcafAs2okB8WfcYfw/IJD3TjKWL7vV2qMLpzB1RQ
b9w6phCZ0OHSMRLaXuD1e/wpxwLTpnlIRkvyXI+ihxBvf7JghjOcWtDkBFap
Iq6f48+UNQ3XZcyeptDBkjSbu0YbkohrFv7+KUZl5X2vIIt7C/26PzMJFR+7
9f6BpCDf4b0X8RUmzRY8eBF84MV9OYRGnROZWe4Qh/rUDmO+BiP7xeFcf3Pz
8SCznPmcgaoKDtAujxn1ADAM0UPfwqrvspr0YnD8Hp9eWW88Kp71egB/4NGA
WxcfB0ZpZRuJgvEAjja79Q2iGlmT8dCbWCUUx21o50fEeglKDFkCi+psqUQx
JsnD7xCENicRNaT/QRYvuk3s0PYSEP//DD/Ak/HeQZuYO05fVT73UN7Xpyqi
J6bibwXND9PWebukTQBz2wf2PS34QyIl9Y5q7HAbUKKPXlJK+7muaG/ZRIse
9Zt7LOFfMgu550Q0qSvniE2Q97L7jyPY08s+QwmrQm/XF5NxLJTHaxmhQuk3
Nw2UrF5MwOJEtk25AoF7S3pgTOTc5kfWc+cEYZOfIGFwC8xfaIbrerIZKwUj
9rY6r2m2NmMp3yWaLyCg9KuyrkbqXJ4lpAyaqYOmeFau3TuH+KgD7wMbTwmk
5nMrWnJk5Jn3H5zhqnGFZnkIU5q5i0BfNzOMaGEM2/Y+CV0EjCFfsEorQb1Y
DMscWhbCE3TwnRtePY83jSzdBtlHmAc7rKPo+q0uQKp3k9GRzOYYZeeEiaTg
iHdxJLILvQ4i01NJjgMBlbq89uI2JuuAHWlllA9Dr8erVRJx3nICYNe894Ea
TAHhb18LMND6+GBdyNi12nDzlFmz1JCfC2ojMnOuVsDsaCURZ2r/KJ6sAPf9
Ofv4ag6sMUgINkH9ZONZVs1eRIJojR1yprd/MMS+nMv2yy7HyP1mfiFr+w6/
lyOiwM4SM3jUoE3uEtSp04Ys50o3ALMsEidMgSXHlK/nHRtCxSuiR6gqO7Ab
n+jxC5AoTpIyDEp00RQeG2X2eoJ7HGcfNovO2n5T4HJNKJYbPMbBulvdtguM
MSDXsEnO4HpXrixiX6Jiaw0tlyYVobnkrkuu4VaNPKGpG2Rdn+kzT2ttGE17
O8guH6uZ6EcpheD4I3WQSha1piSTMCDuvZ5jIeXPLwHHqTHajzUnzzs/DEDr
ORXp1brHcldbAUJzLYrd4B4u2Ww6mAXJzKdFIIgyVRH/J0EkQRPHjmX5Pctf
aTAvRWaMMgR8qokbELU6M4IpahvWJCGzvia+7mZFb7dEwjxviAxHBPItNpgJ
4tZ5WBtdurjtysaT6PAATSo42pX4iSp8OnisHFp5b4MMjz5qYJ0oacapqpzj
0uLTMRjn7vhXImDfjNo4xeDnuOKVw9Z3RKFBUoTxsooxZO9Zv0O1JtrgdBOw
cYuY9/uP+NosBa+wEj1XvTCQ3wQaSDr1xzVFrIfuI7uCLK2etgNfvpyarQbm
tVdzInxxU301vaWKlZU+Po2MvSVR+bAL3AnRweeQ37BQNF+AsujfiP2+HGfA
zK/x7xlvwZLPuH0P+sIrGm82If6xvYg1pM53fT+QOUdFtxz7Vxm1l5DmKUlH
gScqqvgo8yRimiEdauRh65Lqudgmmit8iSHWtq5JUxIiQJVGrU8uWGo2Qke1
gfMReW284z3d9HVw2M/vezNY0CIdNW2S5pWC634qvxTIwrhiQ5PgTLeEuVaI
CwG9uB4PIjgZ9cIZU7Odv/uEsy082oHmKTEX9cJpNsxeECnHyboyEdvp1kFT
pvq5YtaxcYuVKUfIjWCLGH3xFeL8FZulMWNLXoyGzXEze3QFySIrg5vn/xE7
PpGkxLeuH3j+NiHqemhxKNkFb3ligh1zYvQSXcksLNxJFd/doxRU/nITgVXE
fhVv4Awp+CvQyci64UtLTMzQ59ir0Lg3dfEjkt2uxpr5OUfEL84BAu6FOaPF
qXORizbXhlGRZqyiqe4c1GKLDWCFgT8Yv3pvNnB101IEZHKnMvmEPFDCVjCu
vhp9K8UX9cEuEDRAG8vThsNGaVeeap33DD7yb35tL1BjC85EDi2cCXRLczeK
GEejoQx0GEf75l6xGv1132csFjTdX6fwnUA84w1WqANZOw/kvoWZXh0MgDPU
0m4/SpKhBgWTMgNHmBTT+enhSdkyLuyZdPsGInYz7515b/yYwqcB6jfVWC09
3KnqkDvmjOU7Ldh6e2jlwskvoIJkif4ZanWMBv+P9ivxfMNSE+JOTmrUj1tX
t9WDPgIkjbi+nKFszG+dqZkMfN3VN0nV/JQO1+Vj0WoixG/iwV+p8H4Voxf8
X7Fh+JAzhs72x4cRSJPVBKxBYFIl4yp9AnD0jEJucBsNlpnrYowyX+lpUJBM
kIf4AGHtjj2hyYKMXxniwddZRX6L6DMSm/fAx9i+3yuRaImvesJ04CQDR7ip
JYkjx/SKDcKRxWoNCWe07TOZ14W1AycOK5bBpoqzrRpX/ienfDJGhrptx2FH
4YEJeCA3oAL0Z//+KU3uXg4GiqD4/HX3tdvOW7GcTLd9RzcqUFWk4P2mBEXk
CtpnroIQfGX2ype6j/gqRSxTtwiVnaf2zyKfrAgb3mrJxQ7uNx+j3PCxldcf
UQS2rAuDyAFsxPuCOj0h/r6pMaMuanVRuS81QQLVSzH1u+FwxQnKobr1i3uq
glp9i8w+2jRCwQOZQUlmY6jopA9mLJEH9Wt3r++PppY1rgjc29SpMwDzJ753
s8tjxqClaSwZMuvB0TxgRPwrHJyPneL64GtVGpTrr8viSwL7kHrV6Wntmx8Q
PCFHziWyfO0aaXhH7FH43iM+9OHy2Fd+fL5iOjpBjSFkGitFlZPXn294QkVy
yBCFJqsXXgdN0h0Z+rrAWF9TjA/0Wk+14jFVH1Fm9NbPu4EecJiBXV4KVg1l
gYi6d5E+QEKJApVOnlcGeVOe4jPBcprQW9p/T0lmUempZyW+kF04wCD6Btnf
fMGvFuzjIwoj5VpU7V7ef/J07ogNBWK16A50+Rz/mA9oNh3+TPZA3C++zKIO
v+bpQUpcrcQHkR6be0YpRHfGaKELY1FDpUc/ZlyxKtc0/dEb/fOd5eJd/b6w
uMd9wIQabz7sN49tFk5VzGlnx1e3q0skmyVlgXofn92nKRGXZBDRslA2LieE
K48rOctXzd69odRAzFI0+SmTMTPk8K+EhEdWLqw8fs+Tyn2NN2ZcrbTBdm51
XOsWpazR4BS81gV273Rwi9OQPVdUFH3EFC3/25Uk1j0s5UHOGC/30LFkrSNZ
JcWetIAvUwKJSGmyP/aQL8hC+8yquyCMxDVPkBazMydqLvil5cXcLjYTqj51
ipa/zmvJ0wNeFMt8jkFHfONtEFqerGIgOTqudW9FsA3cPdCkmdRdKv7Y9ULD
L2tMnTTk8FY/MBI0BNivSNA+AKeqHwhbw9ExPUtPl+aqgipy+qwz4OndT2E9
NOs2eR+C/Toj3JuM5IYdjC8cRiHEZ6HdXknwvSKfYLqZxAS7dyp5xFGhBM+6
lNb+R10BBT4gF1aJHPjQpT/VPL1S6KBJD7aMcX0Kq2dsMx5Ixu2udXO4jGyG
AoTGUlkI9sdubtH1NJABI30imyQ8ZjdrY+u+W4saY8ZdbwTZkZA2Nn11O19a
saIGHXIGcYbsCOb0f2nWM3PoxpFCAAouDPM0ZiOgua4tm5OcZsfgFR8RnsN5
5cnlhrOwJs13vgStv+6tJdg/UzJfjXDTte43EfXg+DWkYsT6BFgKalImF5gJ
w/dQHpSwRo2DnksMc7utKIK1FVeIMEJfWbihJgJnryGPDNQ9q5wnPcpONjQ1
JCn3Zz1OdEdLBNwOOMrmVipn+uZvivRsl7RIP2BvTyLZSi314ieJvfMnDSh+
KKYdVwZYq+bfaBmVPBl0+Rg3ASYL0Ctesp425/Jz0lh7VUgDAwKCwX5KocIg
YoC4Zh1/570X1ToHg/FVvJpJ8qm3plBddpxodRr80JYUCCo5/lPiuH36Y9+2
p+FJRP3dI3dqVTatL5gkRXYezJYAmw9SVMVl9lmo6S/4bWLw6uufP6c0vpZT
SESfiXYlzfV5Q7HpiTfQJSwRaJNpIlPSCSTTIAPL9wyCF+xjf062SV5VIlip
Rwb2hwYgA1Rf1C630KZ51xFCIpE0TvtASnU2d2TnRWHqmgGW1HJtk7zJdWV9
csWRwrSG8hFmxyBK0vWehu8c1aKcqcHRAkL47+RKO0D5SsZYBdGaLPma1HKX
VQDnlBcSq+O14AoQHMfzpEv8fi8aNNxdbc3D6X7wXX4XkbdITas2kgRKbcy+
K3eaDs579ZYhxjpiDxvvp8fUhDVLWmf8HHBnb/LBi3SntqFyqTB5pTzlTa3G
PjYvFTxzOb4Ml4/hCKZgyOBfD92vCQkYjhDctpt6uURZo/xfTuCUJNU2e6t2
Xp0yqF6vPbalWc14e5Cat5+rpd4xtxCly+aNz2yAC/y7HLtggOPOW+GKxvNw
k0mK/HL6LjnWH1zcUt+v3cBXV4r1wBvg27eemnITXO+WQW3EpMlZXJVBTXD2
ffsHElpCNuL7dr8hR6jnLuxjb1hJhapna7rXNu+mIITbwTOpp9iFPSe7cUEA
eh+Z0fuld2wIz2XSadXVE8mXsIdlyt7ItUwdDYtwNNe8U3uaOYKo5Kz6Ryft
Hn2xbuOb7fhpRNqvRDHWlYaGD/7v25kTwSACq3rv17oUOOzAf9ggJeyradtZ
TeVtP+87JO1t5vXvp46NRd762uTMABirJn/D8fB8dfJ+paILHBTZev0U0z+9
UHH4z9robkGzOyXcQg6nWy+eh1tcw/qY8jQMuMh1068xvPdAS94lBfLswoTG
tDGvask5p6YqgDYmKo4U5T+jiIUkqq28FKCokx7SGVVZlmA97S5vjkw3Lt5Y
DL5b/mDWDMdpchMr382x00lZ6G86DkENlpTxjcR+8XUR20XOE6r0rUKLCaNm
UyDCwiWDMjJLIN9er105sF2RLrVRY0BXmc/+ruAyPg+mdpUw+08VT3N5EA+e
O+XHLi/oBV3DtS6XskeyK7HiXWKohr3Iqhp6+t3F9hCaqzy7BWY3x6vyZP5i
Hn5rJy6SVPjeAkKVvM2JPiSw+YApUBLkoqMdwDM437JgkBmg6ERKdhGKZXqo
AMtn8byZaa23AG1cYonnJGgLotHggOCn05x3+SPKgt/wtDz4Za+LaRYqc4uC
yJ8+G4P1gPFiJPtWF8LqiCKqBZvu9lwfHdlYy4AbrZy7PWmmh1kLFX5M2XJZ
5nJAbLqWzoTOnmuzIbMi/yi94LgxOLI/6q0cksR4jdd3GlmfUFDbVPWpZhe1
ihDE5kf2R19NqwrMl7081aJ2i8sgrInebQtzpeIQIRisgJLcXb967t2FY3yT
iOGl/Sd5aR3CIAni0geIm+kFsAggued2vGPmjTTLRbwsX0sHCLR7SjoGyZlS
Hze+xY+pdio85L9cgj9FQsQlLeNGy6O5khH7fhfuqtKbE/r0ehj/1WAM3x5p
axnDurDQ+1GyfubUlYGh9VvQ/ffqc1hXuvC2Csj7AOoq/Sg0SXoUbcW6bd20
QInrWogRa2CkiiR5zyBe57qPW+VmTnJEfowWW1ezdmYgVpGmFewsIQWmfkL8
eZlDofPxDX1/e/jqodNnLElx8ny+svYMKUISN+9Q+suL1Gr57WZwJ2KusnNI
NxHIG1wkNMbYJSIpsueB0NtooBN6CV08JiPqcDFwoAM6P/1BrH5yyErVBoat
Bqp1sq2vJofsIkiqY2NI6Dk68siJnoxN9WHMKC3Dm7LNKysSFgMZmHPwYio+
k4i8nFb2j7upRkeORThagypIHmyPnjYlBb8yV51K4Pl7MvxxNM7TIJ8y46oB
LlBXGbB9wGMni0A0T2MS9qHbYVuQ93GSwGH8SSMtR8kz9tnZphvmcwhKku5P
AhjpYvvnI09RGQYFqxNaviWrXgxafeml4lkukihdWcaSRLtyJWEQ4GFuJ/ve
XkkXy/HrtAXCe34BDp1ifrqnHFnVuH3kvivuLW/R2CE4ZOHpoJWQfZC9rZ06
Xfxz4rh4Ck16OmC2Cg0VcoISmpihs6UH2AO3XAKN1VrN+Ugr699IZtpcgfk9
FnvcDuSnQMs7PmjgBb+R2ykpQD7qASN9XGbS2gR2Z7u8U3rs4cZIjI22+XeE
cFDe0QtO3IM8t0ydcSAK9XQ2ypvhT0aeGBLrrVnFmXA1yw2fIYzXb61KXq+m
4orFycWdqCy4/kkiN/703S7bfN/XbWe7+EkGbEAxClhjjXtCofv4x7kVtobr
SdqSMhO3XNj/FtYNEXAEOB8P7feFMgMk4R5+5YvdnGAvRpllnYQJWD06k5RY
9dg5SimcA8JVgzXGt14HS1bjXQfgS4PbH3/I0+R+LnT+TmQP5eGH53cPSFjQ
CdWIVbThW2LhnNdEMvusLEQkfS7K8KEh/4Yis+TV2jm0AQXqcF7o/CT93R1G
WPLYzqedKQrmJZwwN50ZwHuP3B5JgApAE3ZWx2Gtcc281kCRlv5KVMfYArQ0
841Pud8Ri0vPpRWcvSGj+EMHmAFCVnQi/ajkE41cFntHXBJ2KY54hzF5E+z4
XHr9JrCFJ8LDnsEYt5vCHR+hAPY3BnrsipzPtN1X9Tg7Ki0/Y+8s7CyLgK82
wp/aBq0jT1J7mHWepC7v88Pk5o+D+/mpjPH5lpp7WXTsTWRmy7QjVFwEUtbA
RYKOhS3mzmy2ZHv6jDGa2GNT3Xse1jBzJ9DWKk1Nqc/R04MtB7KlP0cmJyrN
d01UlvMrQ9LT0Aljh/N2uy0sAJfJhMT4TqTynKx2jEivgKBEaLLxz/SV8Y2Z
AdACjHYLMhMXElHskYnovq3Gk5exPvpFNTL+9He7zq207NlxryNDHlJuN6OT
aZ+KD0o0dngz/3oiBlVXN2p1hqzNC8n7V2Lo0OEzu1z+o8cK1NqVoeFXvI/J
3XBvjHa3DumHtveqHlZYILm2jgRMufjzrgMCITKGkM1Y+5NRoWQ0jGvtOvGN
vPkUNEA3JQAzuf8jdTCdVQY7+UxFj8Hn330G50wUO4czKCFcAO8umYbOyRJt
9EMNLsTXAgwQH1it/sZEXMUWcGNMjB+bfP08ewEcIPgJ2sSHcpJWNv/xiPaQ
6UHQnsYvRPnMy1Gf345yz0D9yMV6BuGq6eHUsRMHx9iPmNfGAf09n5v63im1
DnGTeeffui7kj5iwIAb5qVdUajFihJvZZnExpwG/URgTxOOOjl+P7pvk59j/
zU5sWkSqGepYuSLjUN3ruVpAdzdKlPx3T4v6WDFhqrUhhtmN+88HxFkQC406
O8LUQUJqUZSyQLtVT1KsR+KItkmvba5A3nYKpDngO8MYP8fRb20GQ3+RcTfz
6oAAHdCDt3voO/WKGMZ1yBpsqTb3yVcUOCl3+TIzLlt2HfGzSTaIVHoZlGGG
BY9AV2aCocuAvZx8qvwuK+MqOVobOP2v+Wr4Uo4Y7KmAxnfx3/NOOGPo8wpM
te/huTXRSLgGKSjkeP/vxk9SZPx6+zQ1NwDLSbwrt2rh1pToN/J+c+eBW3rJ
gumBOVONb8UbR/A/B8BwtoLN3ClMg8JbspAQxGSc2bnNT/stju9ghxfGfANW
5MGoGtiZoWTclWE8KmEBbcXMZv7MiV5+CwklI9oQBsq79DWC1lgzQxvGXypN
oAY/KJ8FqqYKeZY4YiNAXY14DAppQ31SJs8iKauSRYA4r4FuQaPn3nEJeQQk
+TK2YbMxCOYLlLoiiEvyu1uNCDg54ps+Gp47iL3yc7+h2ul0YKt9soAFVvUG
ovCpeyh/dEWSN/qTTbTwwV0jpaTe5au2poVMVLgmHf/Ac9kEVV89CDGIUSaH
mlE+ZsI2E3juaJPmjVA7qxud7DyFY13lveMTs+F1qxLwjQ6uF9DtdWh76JSd
kQUvLkoTV/pfi4NH7BiSqs0NVtjdaXFXbloEiH3e/la7+CDmrGw8j47BdvH5
m52l0ddBtbD1sSqwsX9/3v1X1DgPqy0PYcq/P40tEkSWkj+EeqCFKty/+q3G
bz/f5s/ja7yEGdA4gUxHGSKlyQuVEXo6vV8J1WIEo4TTAfdtr3oWJrltEuel
sBQfz/YhpJJiAwqdbccyR0NNf7U1g9BLVa2y/daqIe4K5MweMbqJ4O2o1YS3
8n982n5hfFO2hCZ4OVdeRqB+1Q3P3rgz0ipnS0FrwhDjmXL3kmkH0q42B3BD
AKdTfisl54Rz3wOO9npjpti0TDU4+bg3sgwex1qJ3lG3hNbb5U/bqLRRsKYh
5MK6QFpzWtICcNpMyFjlxDGpVmTm4MWLSLvLmTAGKcTZIKpyrgp8xJBf6k5/
2nmP7waMBY2+QB6yh4qtXuL8/LIlrLr09jxImbyVVNuNSmnj7I5xqjvaduX3
LJVBp/RwHiqWgUgNfwA4haMByfPPlBhALwoAaEzePIn1mv05BREB+lNGTsVH
/R6Qic+EaM/I6FFAq9l5884B3fvNlzv3/QeTbkpfUhGJvU21ZPE/CXWrP7ef
ALmyYCiPqDKYb9mOZS0Hj6d51Nfj6A2J210CZdVZUPYHcxkLb6Qc+GGpgX68
UdQ9Ssg7fqfwRJdIQnkOztQmAIu5IQnM9YRCkKPwJi1QZKSp0nxJIAnQtA7M
tQ3+htVQ+2UVVrzVZdXe89m7kzCTpgcIpsIoS28zp51jSb+H5QjlzX6fIFPt
0BNNXtq1yKYBMB1pLoDONhBV7x++eI8ERMNjOEBIYy35G644zA0q0/Jrv0+f
QK4VTDUUdz2bQ9mTm8Jb1AWjAPv03ht0eQ+IoacBUMrGCoJukq0U7c/zIs6e
8pI3s9C9q39k2wbal+FGBIeVD+Z2m5vd0Vh9HAK/cG9y6GDpu+wQCmp1fXCW
kzMPhwo+ul6njeEfQImMWsEjeHTOtAvBh8GbPETE/ksSmeifgWPUQPlaYrCO
M6ON1fqjRQk4DRCpRwMRZJxGsCDeZw9/w01pQn2VPywghkH0hBfBaTeNu2Ax
PWlB9OCNwBFI1cxXUAL8SAAxvqSXHPeXAqFxgHvTWXWRzPeXKlr8awte1E+M
CuImJnpvj1HiK83jnkwYPeN0fbgmEO2sFhGWurZm9jSZSZfbGWswRnO8a0SD
6voG+EoMwoRrB3WTNWr+FYuZBt4m/LizNRq1CetfSKHV3PtN1nMoxm6TZaSr
Td+0m4nwXYFkawjKmfC6T/QAJAVa99tSzELA5XJEZ5mwH9y2MJMnSG7RvQp1
+So2iLn0YSzbGBMDfQGdFhSwY6lSj/jucGkQFOiWMsB/HqEX/V2Hb/eZvCCy
9r56QMG+576ZtfbBabYeYjzsOLjGA1FBESDX9qXsmHi37FzhnBlsm7puhsm7
dhBZLr2qNpWTnrTz0JZVaDQWr8t0aCHYOBxPQqIhnIYJ7nFg7/62M/04+f7n
CtyZ8nOdMRUAl/sSmGeBLJyuYDs2DVus7tI2M3+1XLOM5NaVuJuZU6tCPTm8
5pwpmREFD7jXA/5YttP+7LcGXiji9+76q1y97zGM5Na6eOwd3zGLnKK+ho8o
yV4YFrwwy7ms2hDXXfdtJcWT/Q5roYkUQKxiwieW77V08Uwfguvdw66xYGWn
PoDyEz0CD38QZdb4UOqUdHrbFP7aKvwJFhU0cwl+wF98Zk7RXYUAt6QS4BY9
MCPD3tgLzmpcisCqOWUx592njFEseiE/78JeBLmsCgRv0GfXgjslzn91VAEj
cenhbQKGq/10Zple2keA1nmlO4ma6PEib2eHCvb6FYCoUFcqx1q7KnjJ8ilF
BwWd6lB6HwkZW0nuQMQG4iUDlgZsXi55YTuxSOnxzS1E3qWNivO88EOgD0TO
rJrZIUknDR18/5I384UCS8y9toqGGx/ZqplKaR1BJrE8rErc4W2h/sszo8TB
1aZoeM4aCOMHeVfs8H/r330OtEuBefbXV6Bp2EYLrl5FgIWX+VZyskQyoDHe
Bes6e+Nuz30HkhWy+d70Uw0dudaW0n9ebPavQmoZnktOedwBiLdbdvrnZ/oP
0WSDlv/r5E1GNlePlzKuPf0ijKUHgInROCKRqvjp49AKhqXxjxawWpkIQ9vZ
3SwKU7Jrk0Yh8ldIjA2Fg5z0it61S4yOAO3/EqzkBos8kqUVG5EhE+RR2Tuz
UZZnp8UjaIRN1TW307xfsMtbq3nJv+AcSMNwOokDpAy30apdeJSgl6uKJYiB
pCBWiwqnjGoQgV7tL2wEuK0p6yaOa7JTegyxuvG3t/8XxFLPEA1RyXH+ym1j
RQFoaZLAfsi2L4s4A5KjoPR39eCdilMG5newNxc+imjM1wlqPmej5zlUcqPx
H7kBEPovE4a+wwNkHFaVV1iDnnyJuUD0p2Q91kLPDVkC+b0VDR5OrBwn6FPG
kJGuClvPKzUGG7f3laSYsfdqeF9zp5c5+UyCkN05caCIKliPUyMl+h1C8bUL
7lM5gKNyVuSDjJHTfApl1YeYZS25EVxVgq4P8wutmUsoud6TF0y0zP9dygVb
EKt9DTRwQJTM8H5ldw2cKpmwI/MEAeM+rK6Pk9TjpD6qbH5up9g0byMYFkVC
r54PakLey20upNgY11a15OAtqB90UHRLwoRfUiOLw1sF9xVelhLEkj7bta9s
8HuW3lH44qrnXbwj69Kui8ZQRBUGEibsOVhBcVvWYXOrV4urabpNecNpZbsK
NBse1Rysg6V7oTGD8CmToaX4OknGiYLqF0px9zrwGmyr91AVuY8g8JPQecNA
ngQiLyqN+Mf3PeQ3Q392KC2zIvoBOuQWUsjXPOWqOYjaYOWF7KAmjVRrQyxm
lgtd1riBeS7AtuAVib4gS8L7MnhhPKCgviFlRQIz/+rutmnxcAD9QVX7PKad
2DabHj5rll1SAbqU82kipwRTOnFQ+iRPV17DVe1lcLAyn6wlSKWRK9vgE2M4
sjrdkwIgQV/47/2X8u/yCLFlU+uGIMyT2y81YGeg/LS69gIHEHpfGk/g04h/
+AmYrqZLbgwOdJI/YLGMMCVUdp9yOrjryqsdRRYmXCa7dE8pUqoah4RH0eJs
0DNntUNA/qDzIRHIXb8Ckow27vEy0L8EAy3ZKTZWbyyM7yzVyRiV41dhbznk
4EVIewGFbEETdsOPKE7kn6HslNHswnCGQqR5A0K9r2qvMRFfA0gLF0AtMb6/
x88YsgPID7xViJszj7wk6RxMu0aQNAOHns0GOSX3tC/ucuLeizYz+E0woyCk
E2VTV5B39p4tOgD7ML19iCi5VZwjE2p3R/rDGUEv21R6XFl9ZNjBCff00N6I
XlmXmCmL2Jw1Q0H1i+AlwFwkUqLUFTWqk9yqAaQVHA/8nLtiA4shB+gYA3yc
VJ/oLrSh02YDAOwNArDpaNnBxMZ9fqy88FwYE9Pa3+l1THhy1d1ozIHiYvsP
E5r34SSdXqJCqF7MR9sGSVjP121w1NbrIZvKXs+mU0gMcViAfJWlJziw1N/y
0cilgoIDC08qafw7CIt6T+Ysmmu8IrvG8htWxQMRh9qm8qh//+mjemfMSMpP
Raz+NK4XfKKPUpytJ3iGLcT8S4EdkTQg4mkpr0MWOmX3ZXPSYkg+GCzRecYf
IiHYGSx+9UuHLeJXNOaBfKi7LMkViW/kXWSWuvcNtNNIi8EohHDCVAJeG66v
A7qBYYpbsb65eARlw8mKRFpiSvzxjlm/xb595uRvVupL+Jq1I+HMZNWwMVZC
6CJ1Trtc9LxTfE7V76NgakZqn+gNn1y4mlij0qPkOko8ZT05uXj8+hkZ6NpK
hyPFjWceTsiCz66+ZdS+dYj4RewSV2murIkysxYEGf/rzeIbKHtFb4bME8M1
EXRZ2cKoutSxNTq4mdxKfe/pGWiydPS8SVWEuNSLZI3sEeIC1t62qZyYogtp
ZuZmiUcyuzoTHyiwHCHxoy4X6mRmKeFWt+Gp7wKE/MWklID+yP96Bh7Yd4aX
29dc6T9wA3Hmvy3YwI4B5ADDQojkkhQd/+DSOKLBBxUIYTJz0Hp5nUZE2C5D
tt9g/ECxzHobs+ViT589PqifPcqRn+yEYgDeLT7ThCSEfXnUJ85HM+Bj+wpM
miy8JuiEU7LZH69itdaI2FPSHz+/SZ3tUtqQ+Z3K8ZKrOc3pRwDkligXaPIr
+erV5iDiXzyFDGfkX0c/O2cO+i0133H/zSTkfU/6+Rd81YO5mo6kd5QWI6A7
X+RTvQ4W9vFOS8Jarue6lzFNj8/8kOe3PkosY8H4eQgZQeXwh+j7aIgYSDh5
mHhZDnhLs1hyGt1ve9IR+VToIrMUFQQbzmhV6AF1NQp6eEkkuC3jUYW6iqfI
J01k1hvVcJJ0dwRj1ABcvMpFMdKioFOoPsrvcaA94nsJyZz2S6XIbzfQ15Vd
sj8wX/iC6k8UNYD8/MfMJy9YY1diyHGrbiXaZ0LCfMdQMQQnQcdwDmDgPvw1
ze1PS/eAlv6oqJ+TID/hnD1byfGcVZYnA/8nFREuLq8Onnnpi2jzYCsIlZoJ
tZUULG3WHseBd1MhYprUubsXb3IEjt83bWbQ/e40s3GF0cw1KO2m6M1Rtxna
U/KQ0vM9mKN+v4CG2aL+l+lHW2OZ3x+a/ycwss4I4MBddtWFdwfvaHJ4g5AI
Sd5nQsVnNDJAbPSFYD9B+lxnc18FYxqp1ETxmp17SBWfxAAtcPl+BSyQbDS8
jVfveQheE2FcMH/kl7MBWniYkTfa8SIydlbJ0/IIxKWR+uLgUHG+4Tun0w2E
IjnbAKpaUDzP9jzqGuilwm0Puk1ZmZAEedRsyk4cksux97oke6lbjFDwyhDw
NE59OEbn8Fd9x+EOtIjXCSFHQ8zTVsyM3fhNu+PMVblyIz5LmU19p6E69fjF
ub+mUavPTytK7APog/ty7ceIJCGsgocoVAxfnCzx2jTRi1ba7rppNBHdc7G1
52zt4aTH7ni4mmETZvWoGrDN2THyQd61yDWnHNSzgtxNgpCZ1PvnSM/p69Pb
07Cfz7N01I/aqmX9atVwawtceGGIFVZyjKR7cC54MonVy3VBPWkw2XENUjLP
V5Op4VwbBMUzOFgR4caufbe/nzsqNBeQElPFI1BkM2wqvw0QndSc3U6DI4rV
7qrr4NKNKji+2kMPKxdhI/pBXTjUdWs+TPSeFv5mywbEE/NDG4P7F4eGvmdf
gvSLXPDO+mJnLJwAp6wdokMIgGpIaJawGpV6PgyWWpzcXwP5hJQVtM+sPvaL
l7bCaqUfqHC3XFktdincX+T8VrvrgsFMgCOrQwnFAnVjNhgeynr6bMDzSzio
oYWi/01ImnxdpOdTXjzl5iiJImU65KLvjhrnHih8fTLOYqrsZXLII7pRG5RY
CWCIfzvutcZDJJgJQNMoM/Jc1MaU2ekaEgrQbWIeiohkY//ly3myp+Om/ig2
ANsTwZL6UzOcy50acd0QC8R3qGhYjYCfAL1e/ACMHtUr5seZFtkNmdrzeRAh
rGb1xBGl5V5luviLuT8mcGjKSp5KYRGeuuWvGsy1WP24aWjsqWE+C8WRrQsH
vOJgLFPbZVG/bFGSbOxM3tOZa1FfBwKhjt5Ifmgwhc8zjzYRLLR+HK7o3YEv
Y950fo4A2h3ysuTQ8hfSFox5ArObrGM3lOtMdMQENlP3S/CM8xKfM6TOWzRQ
7Nc9z1Sfb3HFS7aYpxFh+BQI6MPk/oIiGsuPmCdNSZF2Ton0m9VxSwWXS6P0
lgV++LCmWy+Q4/VQP2SRwX6UpbXaJMZlb10vdiNln2z0/4X7gdN2CqLnj2yA
S/PHzeKx1NwQr1wB4jDwVNYtfDg1KZbg9yikN2HlEY2SYKAfKE1dRpUKo90a
s2pBO4G0oefwNM0CW4pPkUj5zJ4Ab6lA7YAE7ZJ2DePuglwg37yFVhvZPDDj
av/apeVK2vXb3gHc2lHumDYOdNLkVZKoCXQw1L40yIg+C7Py+f6ZzOcDqDnl
wAW+gQ+fJbr2vXMX+fjrN6kmiHPU9vaW+PQSG5gUd0Ono6m8kqJgasUuCGaG
zMUulzgaij2D50P/8WlbL3n7tJAyA+03HshBIO2k+z3tajiOPkmpL6F9VMWU
bkpR5KmdleSLVd8gUCgUbNCDpanCa0zu0EOREYfEkS8xYpL2hewEIPbszAT0
uX0XAaEgvQyjyYkyY3L5X6e2yku9qE41qrA/lekdtRgCQajNCVBdlQQwbeB5
UnkOX9aBTx7FHihrCva/7sUNAm9S43ZQ4ihT6pI4fjIM5YV1tbnxQ47LXR52
rI/KEmPMQMJH9Tr6124+N6QIHSdRBLCF1HemeI+P9w+xvnuJCcXmf0ZMWliR
SNCWnuoyMwp2uuVOE/Y6OkxT7TD3BWQ4iRo6T62Q/fWseo/BcWlJ0KNYXZJu
MpIm/Um0+WLZIWFQDrP3CJod8HxQbeNLJaYOPqw6cGZl+mM9ZyT6l1VYprWB
D9nDCcUYFckl8Kn6RpkYlNbf/5VP8+hf5uWxUvujmD/S0Df3TtNNVxedprAq
N1a+EPtw38aORr7Vp+Fo2RhuQdoDtWHgf8ZALxkAeV7rBlUFCOLJCjUnjAZ2
i2siaypi6GE2O9NXD3cL/3lga3DkFdA6M2n3E8QT+ZCOkmZwZKfNZcUnqdFP
wLz2KL3hc9QZSXuE1rDjqEEo55h51t3ipMzPKyffBEPj/OihsnQm48cLGMMz
YQW6b9kFf9fEnxBUizuxb8YZsQks0jPt6OMFPmo6fLD0HjOWfhHGFL0FRngv
npgV9Ex0yfUHze9fFEVYNlo4NeiNNt9VwQulRvSxUWXRxKGwuutKG7GsIzfb
dERGtvgIvEQcpy/R5h0AUQcdlIHctUh4kZTosgfYRNPu9LztoJao46Dh2CMs
hNuFJDinES1D/SmmDruiKPYwjmViwLTQRXzBzDFDovZNsw/6V/dCtbqVLUpZ
CrxN6ig08htdiWlf4fQKiXg3qfzcDdQYESElDgOL/UjUDM6PDcbdiMCQKMt9
xtJlIDI2Q6u1tLXigrdiVObWk/fNGhv/SW8LQ2Tnv97Pl4Y2S1A9gWjvCDCR
GNXZeWR+n/kpUJMBPU8vysMAz3w8rei5y8AYiEpDSbXkV6cHX19nS2OXLgtu
+od9Ks4XG1WaxzkCWIDcTxFaa4tkUcfNrOmlyZ22j+sWnrlgWltkdGO9pTIu
XTr5eD3iKSaEOrF560+rxaac7kWXplLdvUCo3uSc3Y3TM5/oJirEsWHg1Wfe
bliZR6g1sBYfMzcO72cBpYxZlucgWHazSO/KTDT9C9Y58vcLeBjfDyyObNDU
UKgN/UXhQdOt9dqnu6567lQBbKJjpMepszM50lOlY8Ay7R8oa2VHWP9aDLYT
+lGVK2QIRMdlWmtL2mEmPIiKF1UkCo5GzZF4mXpLEsi95vRZ+8KH1kmQGewt
ZXVJSXcg3UpmTW20qbWiNMzPgE964pmGsfsTUzzJ5cgisSE0CpK0Xk75hEzO
0haY0Z9/evMJzHsWIbNPbMp7G27XkNvlsUvAUKIdRvNzBO4Mf/fCs2x337zk
tYzF/je7RDZgt8F2xDlrWvpzcyfysEAbAQNwgr/vrkojFLJWY+dS7gBbeova
5EGSJMr5+WWvx++6+GbiTpMOV/39uzOKZyUPJ5E0EWLgEo76xXvGnKuLJes2
5TcGmFEeyIc6/mTu6IRGboKmAserk3BHKUeKkTiy1fsuS2dKgiUT3wFqsA3R
/X6phGOpgGN1XKqWmAjiwZmQuxfaCU+hpHkDms3dxJuCq/OqGZlukMzMFyLZ
+9k0JJHLcXF3A+jiYXydbfFnGvA2q1eAcEeip00734yzwQExmfcBi8t/Bk9/
xlpbgkX1XjrgP9Vxq+6qwiuSm5VdfS6gEk8WiM3BVazkEJ86SwF51NtZEi20
6qDXGFEIJrDwLPbmNy8N51W7jpKjTF9HGZKoi+fcOlNPBMBWsKFrcbFFeflN
nmGLlkpjzEfSq41p+YhBEzkX13rtrsBfIENBfDNML3W3J7hNXXZ89H8Napla
3WyjCBS9HNMdY/zkWTwsAlaxDnQDiUthv2Hy+q0kf4bQHhJdkRghVxL/d/AT
llIm9t7hoYcsZB8GfZDqr4TsKvAZjAqNVLGHTzAeZNP7x/lkz20yF8WD4YR/
rdcFBI1OIM82BRGJO4BsATtpCcUlaBjFyjfX62rPsj0+Gc00RI+vVrkIoRfZ
H4YLvzd2QSWhoWFbiIOF7gGBB7ybSASFCEOgq+6uhTlumNW0/u2f5KWOBg/o
+UDmxi7gB3k6njMJA7bEKC/+ClRtO/ckQcyxvqo868x9WZxyYo1SyHXdCulU
NGLALw16z9Z9HrSL5m1q+Jd0OuaygiT0v83paKmqKF1fRcKZpWTW3uabBD4F
idG8FjfIy6LADU8INb+lCBd5D5AkPbAnNomJkWeajMDlZBruJvppCH9S+OHM
cZDelC58ax86QSL7s47C0aLn24XffCN2etlq/kpmo8O7hy6bCTK+LlIvtCA8
4vTLhf4VaZ3YluGoy4EpufZoWDkCjCOVnbMvNbklv8jk3kUdMMntqGfVMs9Q
A4G9kilBrUOOGCEctJADCfI56L8VFVcZ5+wIwkhvSf/sVPs4swYO8XLO/5tr
3vEWpibtnuafsYl2gL74zPPM9bpkIUbUSfSf4+k7y+DL8rzGeuOiNFYrSnl8
i5dg599UZnIsqiqIQSLROzaOg/3nVJ7/9f5jQvrkFm5KdlpMesqo1U0XXu0e
p97mnOVJt9X+FVQ3bE8lhUQgtyx+PsOlKAmVUvhQ98xDzuhohr9W4tE+LkuW
1PaSGwMXnT+WwqGtCZV23SY6hKHuee2T1SL0Op+OzPRoUKNHb3rKCpWEeo0S
FksZ61kKW0Q0VpfLO2zz6C5yFDKicLVz25HsfKVrRvKMCe89YURhlDoX9rHi
+5VCWsV9BVHex28QIOMgO+noIHkluX+HxA+oGwyAG5yFx0Nt6acM53x6IB/T
kqqDZNzFA1WQBdUz44l0VT7ZMR21AeDa5aGhUWF2t5nzySTZloXOrUZSNcEX
IPFqt5UqXr1DwE5d1f5MK9mhJdDx13iStAKz9sCLgkE5o51e5nAk3mHjzZV5
sXVQ8Gt7z5gbhbg9KPZEkKsTP6h5BS8EVbuqFNz6OzN/Px5xK+kwquym7XUr
JkbMcB8vnimtGqOPYnVvD5+LEoalnmnBVb8EI0rdZbZwodcJO9IxdbA1wzRY
MUUuiQ3XA5rfeLG6i2J5L5Hk1d6q/yV7sfULoyj+FQQDlBEw36OLNvH89rdd
Wh4hCgAYl4WC4DdRZULLrWa4eEGMCHY0f2/Fwuoe183bANC/vcHtr4OmkXgF
IOeo8Nr8mGIPMebYK9KcdCGlws+3e+dnOVj2dANx2OvHroI+jXegHuOITpFi
Y41i2Xvfa4BJcRNVDl4R4SSWmj6LMYQmpXxxnjDC/HguKhIDuHWP8ish4AMF
C5YUdE+ZfkMn1EJxfTC8jgso5yRvJR9W7FAZVh/AExdLM78xMpZnMd0FVEcx
F5WUZug6mlNUqTGdXD+0gYLW7/+LXLEsvCTmnIKIJwnewWvpS0QvQI8lqBYF
scgSK23cZWqrPF2jCYOcPQey1GU59eQgRgTMVsdyQKN3y+Up1qxrvXytJxRn
IwyDwDo13/yN/hWTP3PanKhiAGMH/ZCcMuKWAHa5kQRR5sagJNeVRXG+CZMm
YOi4FeHo0jjeaY+AvQkxKGQHj2beOD7LFsgMeLH6b7NXQW4UpHkNDkg4uWF3
GLUujWWyHk5URhXrzUw9D/NU1S2OnRmBz95aSfWuyGR/e6OWUhfCE5rXEwv3
KBgQUkmyqa48CRojJlDjicqFBhf4wiqjU3iSKxrmE+bz1XXc0k0qlYUPqTNt
GFAfRx8LY90ii3KjXuy+aHnGsPo/pMcPWFgR0MfzfP0juMy2ixaOuudm4TOJ
KaDIrtsykQlHrPVSIa81lrwuEubRsgSn7ARVvBCA4TQmQd4TMQTf9rY3DYi1
uexoTZNR/NU3FVkQeEl3EhbMlgs4GtegwQR6prdgxHEMwsqEgzmNgySfqeUu
OLfU4p0ChYRV+jyyR1KEzhLrVNZIpx7MdXvwVbYb+tmO9mq4NURoOZQphdWi
0PFtmS6/EG7dR5IsxlWWLQIVXlYnOmnW5oR0VelYH0DEdWYTEtZpi7qyDiLf
7ldt0bjvnYmSX+IiKMAwwWy1uFrqWIOhY+C80BO4PR7XzlFxGTsOoO5QdZiO
5bd8BHI0XChd+wJSgW/L4JIALjFVaTcb6kI0uM8ND5q27f5tgJak3GLhPVFK
YCmgLgmwXDohCWrp+wr9Y9ey8ZVEo+OQEuS2g328sGJqwHV9aiPhC0R4m2Fd
xJPge6/a3iR0zU05tWXUjfQ+Mlvnf/fCz8piFwzBVlQ9wPaDS05AbSPa1CSx
Z6wVM1KGHjqkPOcbJq3yybfEnlQom3Ns5aGstogINA0mfR8GqbTPvJI+TK45
3o3Cm1OKKOU1gGBUslRTATrHJCqvE79C0jq0ndhxF1E1Tx6TsFPE1p08KECG
fvYCXCf+1wrGhduuPa2v2N5fHYE8ONB8Y/DAgRzwwdKJ9/InXLYxZlpxbv6F
B6G0ERMX66tx79KOqHMtuhHn0GlTPUHNbzDHyNzCljHKXpPz1EC5A3bMiJNq
wcuDsMw6YeBS8pfk4N1rzwSVYmCyrJ+3hsO5eel/3jVQmCVMDaDg7DYwkePH
aJrmK8pM/fOI2JvLEQV2UisVLFFNLFch/oYYuLQi5tVlOkJB2I2tI111hfpy
khab6jVYy2GqmJ+2XY73EWW3JYL80r6yZzoB8p5JcSZozPnZBOoP8Sii13kT
C+2yvWutNJqKm3D5szqjgfPtXa6ZwhT0aciRiEHVfhay0fBVhFkPZRzDHCGw
8//Kk9pgUDeMF0TC0V3TOk3HIUY0RMZA24cgvTGOaluX4LuLhXiJoxoBbCSI
28NmRJK3rUq584zCrfNUou3uhNGQERP35UfUaACHrZSY9Wu7Mrr34iMR4gUr
TWbpBZ3yYwbX9zLnvyHcRKASFam7wVKT1IHkw2cPa9ZB82kq0M/1GtnyrEBl
5efZtUriHxOu3AG8U9TVR54iDCzYOneRH6COLrjlHgm09euQHxG0KJAB6Edw
awKV0laqmFjfte8Xv7P4JFGuOgU97W5ji0qdt0MhN4d2lee2LCoz8dUPWx5u
yOwj8y8kYpw4EkvcgNqP+928tY4FlKCwLFh5lpvCC1uQ8KkxPolUmbtlafVn
DLWf44VF0kpAo1d/EuND8ab6Dt1+szY6Zrm1JFkmH5KWHR/1ZiaGbCykZcRg
zsfPOkcO3WUKrL5BCj+xV/fHme/XKHTbzwVmkyyfVGmt5Ht/SIUMxd/vHTZr
gT+eJLecMmSbEnJWQ97dbSM2qcrRm7yobJc1fUDdEy5lnzNF3s+6gdrhvU4l
bY5dtTqbo4GzX8k/mTg7K4CDKhZd0fIZdjovg3iMD8SGtUHOcdhbdlpHBZhw
3mKm3l8qn3suKyYvC+ez1v7Oy4LzIFJh1a2jZS3KSU8CI/XQ3XYuxXxJbwOs
jXw6sEbqHHeZgmBxW009q29unhrkTaVv600bDptaAwbMSBvJqRwR2iOK8MA/
sOgsG/Nokac1598c7X6n87fSVim4ZDQYARbjri9sJsLizOVCWUOzcqK5nkhd
DjNmUZ+yLL7IIGiCYWzX/WNLVsnK32lSF0hHD25K57ORW4s4012mt/UKF14g
cjWXtY734tzLDwPjaVsvENsFVvBuJwxLCRH8PRASiOyUApwAyXgjyfSare0E
Jwp9QbTiV+keIJTi8h1DxUhxpW02jWW9tLyhxd/8wsUkxGO2u4Kl2rjjacb3
3kwQYv6Sb/+ZI4ii3hN+iseQ0LXUuTOx5HO5wz8gElWTFSUDXh+sOUVWaNDk
dZRbTolCzCgWotFZBLLXTKmOHffooTmBCJ7WpuAML7koNKSlaFjzYT6kMUOV
Hp4Vu4sk0LBYIj+HEsXEqICt4QEAhPdr9mXoFRdEXd5UeFJPUkPsGA7twmBk
2NI701eEx7w6Vr8P00d1wPbN4w7S/EIEWRxuj+s2HwE6LQqcFpeJHnIa5ehD
j6rj8ePUQOkNgjKmXvrPTSW3yu34CRu6vpPUo9xDdQBSYgxZnCvFpEuNMW7G
KnnvHM8CWdsjZYqXpvorlGK3Sedm6dQz75kDIrGZAs1uAyfdIBxSTiqDkpeY
J7cM65gIWcKHSxpajCDKVIWtVkfkyHXipwqUBMYJzmkH00v1KBP1Jf+++b/z
SDVubQazSCGmB64+4EmWqX3zVGfhW0wmSk43BXsyqgYLHrV6KIbMGn90sLS9
CnPlCpyT1+JzO4B0cFajZf2CSW3clnTOi2qsCfC6SaFfMRp4sD/xZ3QJxpcn
WHOl7kt+937UBZ1WwwCubLEMH3YosnT1j77fquVZDif0khk06P/M8SwNiuuQ
mwnVLAHUg0MkikADHShl1UdPjBRRr9aEBG+yOtwlNjwPb2OOTO+naKeSxNdp
Fv33Y+WX28nLJez+iYoTI3Y8ovEccRqaMDN0+WYPM8o6ZuJ7eoFZTYU4tiIg
3+dkysY4QiC4gQ0jb0fuPm0Dax4Kwz2qE6ARRGVOdeHDHJFZ1b3Dbgzr1cL9
s7tcpQ1EnWAwV/+H0tYVlMw0Q2/KxgqKCqN31m7J8I1ve+OIfs5auMl3ugPx
tTAGVfUkbfGdhH1jWWPR6uYqmCm9TIZpQj62e8U11u1veE8OJB1toYZ5O3vJ
Mq5iGH9EZKMY2pOYUw6dXL8UeDJWAmMsEsf+E96LpIfzk1zxKg5umvFeWFbi
aStCGk3EMtbS8per7BM1+PvAr2MOSKcZUlRdnGi5df81mgIrtqvIz7Uyi0NX
5BeojhQLIPTHQuMduutXYeR1YSFNevPHSfIqnxtezy6AzIYBCR+jnFsCfUUe
sAkhb2AGb44g6h16mig7BVWDIeT3pdNwE3UP+TgdM4WIMo5AiEilcgO1Sf1h
616omXIksfyL+0H6CEHVOKU2HdNAZqiDMSJBoKizJeUKEYz7ajHnZHDoahJL
eODSA6Su0ZIj0IB5CvuEnyZS5ZpWWOVtHYWqbKpDrhxn8HFys0nSEO1m8j2G
jMfBJYFGyf2dy826Y6/lhpvTahBj3Pnu2DoxgChMi3bVvlg5IMEZTskjw/o4
+s6zY7eBjMB/5UxfciuOKbNJAkIG+E5e+lB7KV5/6utQxhloMxMME+04NGHn
G818nL/IBf54o2PDAI3oeC10k+/C0RNUHI+ph6qFVTvAC2xAYEBvt7hq37Zn
zU0eZiTXiGEN63/qTFA1c9QSPe16c8lhWBP+tgKG2dzvtsfQdTtn3rzBcXtA
YFxpUes8lrbXPWZoNQ75PZbY1XxbYuiiN/ZyiZpyGhh7LqgVX3n4TyrwJ2iK
lpMJHb5HXR/IejC3G3d9E80YYnMksjM4k+BpmQx1AEN0DfY3D0IADkB/AJAe
7ec003xDSeTdzEFwUhyaf31sBRupR4zrvIcAuaQdNl2FGFG17UKe02nowWkn
MYGvhd4pkc1ary05No2/vqUj/3qUNWW49efMnxzEtjy6NAgA9Nk46eoQfO7y
GjjKdj8mdV67UsGDkjyA1zWA0xcs5zFbLO//OHLRwI8RJ6Za177BkKBAyv+0
w7qLpXpnHCH7WxeN30/dwI5e3fALNzumuemfQVMgPwffsS1J4/X5xQgkOEVk
DfMiiaR497/HlcKMrTw+bE+mCZjUh+ICuYkyZUErwr5X9yKUxChQoVu9vW/C
xUeOqI6M+yAwDl+kJ08E8b6N/088NWj2fly3rWWsUncOmnePV/MWSpM2/FkG
dKBy1jviS2lZ/NV8pIeDiV1aHkQWdVP5hT4tkCbJ70W2FpUoV5FPxMx9hNZ9
vNvLYNzzaE4VJ4JFpglvxUzdnS+97PkbZRifS+8luoS8gjFBzM6adyAGK+08
jiiQPPf9H/aSlSFjF7eDAPPW3QoOMkd/tEZkKozW46YYBtOmzCeS7Qm/ULAg
qVqH0x63hbmSTgHksPvQnlXleDvc+y+82gYNVG4djPy285AXYarWMaNQG/0v
H7MlqCTluRvYG+m7ri86od59H++v299P5s/b66YNsxgpynfJqEEFcsE3cFsL
ftNlvJQq5/r7+XAOhL8gRlGsDB/yccwrWispyTpZb09n6+eObnDFA2QYneOZ
p/9lGhpiShilTmWbpXo1spKCQTZAefpuDcwDRpAUDNNrKjK3TiIazlJSFeSt
Q+9VSel2Ol85EEs9hIjgd54KoS/jHmKVh5SMdvs2dX1Ty+Q15rC/QXacnf1y
66S+BAxC8TYp2NAB6WueQ8hBN8aNf2Tw5KfaG6c1SqB3Gkgr2dFb5vzPGvfD
3p/jOq7ohlVyNz/ni2o0wobMtMmhPDaKRbgTMbVGcqrbbDdTvYzX1MosLpIx
NuyqAj+VVmWkBOlwf1+i/7OlMEQINcpvtMacZuvSI19rvAzkhmz9rGu8ok53
nXDnAlt1L1s80+WIlJwWjHSFK9J8UBD4FtAnVtLofMTo8MCvfexPfS5XcPtW
Ld1yvwZwj8SLoMyHokp0N8G+4B2Qw/x0WWJuubVz7g2g26ZkNL/RDC8V5D3N
WUGh2EPVOkD76gG7daPjiCE8XfRZQSFZf7StuKK+np4E70Yi4kHWJWKRQiRB
QaQprLN7tlVi+D9XiatfHOS84rmYwR8r8KcxiPeSRc07dSGr3z5GVJOS3uOj
obVpc5JyNgMyR5rmqUFLD3Oov+KrgEp1uizT6+BJZbwNOG6HXTeKqAqXEJfX
KymGGyDgDG0duX2N8ELyosJ+GN3xn99/RVp2dIC6rAYYBNuIL6AuuR0VgE+1
f58PMYQhwrKZsctJObza6KT7dLs0bPabdGq7kryB4LKSkeXo3jGsHdBLjPYj
bDeLhIPTklv0BuI22PUH0fQI12djPCI5oSJibTDG09pM5nnypn4G7AG0+xlp
hllVsDc9b4Bl2tS99pdNQD2QIzpWUQs03VHDcQ3kA40MLW7mc/O6hhXYcTxO
ipKn97TikbvSUvnkJq1CBl0mCWJcPNQ2T/KGGuNuOBIGzqWI6sEN/jqcUZis
peC4/wI/MMBP8RH5dZOQL3n31is6nLKIcLpnPPoiwMwU11FcU/oipqeHJnno
ncv3cu5mD00OTBhvsU0eD5KvEkwOPE6920cwmIGzOGB4wDygc4I/sz7gIGAD
1HDaFZvOeW5zrZweGfFyyil45BnURBCcLlf6wt0EI+/wZER+MJ5+vj08HUoy
FLG8VRCyYlONWQ2gCqEbiLSDgEuDIhOxsG9zfIYV858sp6YwPtcoHbdOJ2ST
xSNv395lBX3fRa/032yHkWUFjQACyg5Fdi5asmOiXaUZAlcPQQ5/i9uAEzRL
6pdOtUgKVoXFkrjkX7X+nPymuuMCjiKLmIUIESYDEnvTMsPad6jG+eygUhsp
whrUkIkh4Vumti6J6FPU2LVAOlCcw3IRdKr7OEztGKIcZ9UZmqHeJhIfJbXO
w+MV8eM5rEjUdA22fwTmJfSxt06od3wrrKrPRpzBrledHN866oECA0CfmzPw
kXHATZ1KJxVSbaXyJWdCMe60mDAJtMg6aWOLybC90iZhehq6ny4n94wPqCW1
MO3W+4B5QXtHgQeJyte7Oy9cDEJAlgcW17HZd245jO0wdbh6X8rRUMqh0Tgw
UtYGgve+1h3YBdlBHOoV+Fzq5gU2+g79oPEmCXDAsUtOPFS08gDnVRPN9af6
9OusIPQIHhSt8AluB9/IPjCB66Vby6Trpg3rrHuHrP5Uz9xgFMden4lP0A/0
PnDQmyNKZTCPaPjyDkSf/7e5B6Tif0cFUfs9TzB/X4Y2U1PRPCxZ8MZu5P/R
ETrp5IYpPC7AisXI1cDfjua1CjnJUwgwC1RGDqDngJgzsZWdjrHugruu4vP2
HTqg59JsNiGOpaRdb9vd8mAzuoJM1rVAX2bNPvc8x9mfuBCh5OwXoWEEM0Kr
LHyjt5spf5hWWFPQneyp7lpEffmyZQjXtwGi8StU5p4rO8hbau6FmZ3Y4UHL
mn/HAF1u9jRZ+xvDCE/jBxsgS4YQ6xyxLUbHq1EJba4WWfbLxn/SlFcsFQwI
3u9xvo7cFvXFC4eBKO1KeFO6EAI1St9WUzE8n20nHcCMjRONgH6S3YEEmUSk
2ObP+63Js+tU8mEaEkWFTDC1bniWOqV6fEZahUzaa+0lRNIZs/uiB/02VaiU
mx7ucdpuacsJvrx6jxEQjpU+2eoey3/biEHnJWLB6uo4UwU9LR4UqBRLN+T7
NzXAmSyMWc29fUHWd/Q7vFmPhgk8p5QzMzMjsilL+FyqUvA7RejQ6k1faoGT
9EJns0Kh3MkMCciTZ1VHI26/5kYQd0zRaLs8bSroYfQbh+Vl80ANoKP26PqI
DQDXGK+/aJzU4YulvHv1JqeYyYT3roofBk7ibol2+XwP3whJdOBehEP4MZPV
Q6YAwJpKcqwZEfl4Yg9FoT8gWBUFfOO9gTqtOCZtHO2Hw1U1j/ZFfIP8o/wS
zjNukShPmon5I9GKh9VzIFQhAOCZyeZcXXvIwF+JO93ARhB8Zjf4Q/XyUKrE
nGW7eKJbhpn++R2qh+DuVv3ARlLnI5wFm3w2Jm3g6qewa2hcVxHlcOVHj/Wm
7ino03Zz6HiAK9ZnNIo8jf+0EbL3jE8FFFyrqXTmo1ie5+VBK5LCyiT+SnQ9
T1wz5UV5uMyMR/qsyd7vTiS3eiAAFHmZavahe3ZCwgq29uSefnNdkcAObaW3
aGyhrbNnboNw/63W5fJ8YTpYNWgC1s/rdetXjwrOFNWqqF++7G3ys7zdZocj
tZ6OqRjbLrvbe840kGvt9023Jjm09Zhmex6bWaYIZ4+lzzsvRq9noCVWiVlq
Mg38BOQgtNuKfHmUg9UDTnw5XUvedLwRUnfunmZQdTxFK4bGzGkKfR7FW6Ox
NeXIT1bmFZ6++plgnHRVCxeGci/lu7h+VparYwxqP7Hfkh06+IwJgoESDOe3
48kqnwHV46LRdP5zPDQi4JS9LuLF7o77w6u7Vo63i8ibUFkztV+VmjTv+j/W
otcSNRu0OGWtLn61u0Z0NhmVj5fu4xfyZ5CfkLTy/ULWMZORgQ0dcMbNg9p/
qOehqesmgZOVR+9oLIJqOkWeJBg58IYDauo9Fpx5i5Prpym0w+6D775/qUX+
m6uOPTGbmr8AWg8UxTAxmlf1E88haKV60YnoYBa6vUaXsmfi87UfIp8CQUgL
RJvlV/Y/hEblMeeFTGFfXHJHt8E+m6i791zjuuw96A+B2p0jrbu0IGQTs6rF
teiRu1niPTGjWgum4MYBDgfrYpcntGiEs+OuqFhUtv4SvliYwkcRPj5IrZxQ
Q0HNvUAAvpVriyiisJHr6TzgskzUMyjJXagJ70uABdp8IOkGpB+z3qRCw8Z4
4Vd8X/GfL+lSUwQJRntcuyzVThpjHLXAaqF1ms4bnLdhkzECy+09W8ibOlZS
6TAulatcNYogaR2jfSoOVAKVRaftkVggCyXy9BlWKbA2WDPvIQVy0cILzNUw
0oQ9QVJL529R5OV/iu9XILVXnXWlzFP1hJAZ4NAF5Ah50KOk3ukOSfaiD/2C
Nl0P+MD78CN9RhkjNo2mfDl2R9SZ62rndBKPCOMbpQdOLrTsbbojG83uAhcZ
0Xzi5yl6q5qTls0/2BXVeNu7GfgOjHwLHHULpGr+NoU+JquZ8AWiZdHkgxH5
8DqxIIJ1CdN99CKgVR5+C+qn1K3DVGYoEjK+gixHqxxPIjg9CeVrQc1cp2Me
Vn7H7Gg3gI3ZGYTfqFavweFvf7NIMqd0aVkvo46PXm/wFF6b8+wj0FGDXgnm
Q00TcAv9119XKVGMLd1UhLWZGLQdWeQltPNJ/MxxxPJeb+9oJas0+sN5Xund
5HFiTo+fRPMXX9EaaLayvgBScej0LucgkaEsQ4UjfzX3Gujhnsy8TH59FidY
tCYtGyfFzOu5lN6sbb96aSIfpCd1Nh+KPTKiQyeZrmChs7DtYXMSBhBSGCQQ
+SHh7sxJLimRa2VP1lGePxoDDT7c4Np2gW0aIimA/0YVFkqpCh7Rnqk0SbcI
uZPclU1HWzqJPWAQ0iSIQ/N2NZvnS7mN6WeTiEjXopDWW59qL2tJmA4ODro5
HPnoL8gPgGxqCchjl7pTaz3YMKaDzl6CVZJhSmKOoGiEacJjpfYQNX6/W5fK
6xol+gOXKSBF9Ee6KB+bFqMpZSBOjmvOOjlr82NcywB2niWowC+LkKoptNUy
z/eegjAIJRSSNeQHafgBbSaqcLtTlawwe9DZP5PQkWC06CCUwTOPX3BF7bI6
BazGu1piW1iXvR8HbtrmZ364yLoquvs1kuMVt8TqPqgqFd1qzGf6/8541HbU
FOD7tFVqPLamg2NhzWXEPPGL1gga/KjI3AICNcvgrpKWECOyECShhy3X3bnI
hnC9auHA63F61Ipu2iXRElZlpd07+Q9cx2spXcxjvht039IyvfTBeISrRgHM
QxW8CwJCjfIu1qSkhaAxItSoFyndQlc92KQGlZjTEjoqgQILEP0CCjwSickR
/aMQTtfTbADW7vejvr7VIWrqHFC/CMcr91REYxLwxLUOD3Ft5EcJ8WHOIg6s
85KLmuXVNyadJrH8pBdpfzeDeo10Bb7/Mz25WJEvkH+mesGBA5op7Q+zmSIJ
bqrXRFSwf3qA2iB3zw2+UgHeN0tPhH5eUKeqlyyBt0P9y2n+19Ir7dYEtnvr
0q83NmWzztWLeAE1NzYQyHOCy+y1qdmGW1wq9r7W49gqLrCO9w/vKtTMe1TO
OYeNi01UNt3LhiQt6uISYN9tJS0djWdbTzKw964QX3c5e2vkfvoXDDlAl0rC
0Oob4wW+ep4Yo94SiJlmpVuk9Wqi1AAgBwPxnwskjXqtxgUBjgB1OWT6UFo/
R2AlvAB0VFcJoU+PfPD2qFELP5oa9EeKcHM0vrpgbibAUV+SJyN2guhEVfog
XsTUSfbvd6E6IELpqbmAIRfj9f0AlNGPMn41QigXgWUdGjY0syruK976d6n9
BYEaoC3NXFJapim2rbFyF4BvVyk79sPRcwC1/9P/l3D5ggTIM59oHPelmMb3
v98eGaNJYP0CzqcHio+Zntp30aH2X2trgjsRBTFUzx1tD1YB97HLudGhY/hE
HXSgLr3IOs5M/9PBOKid1Gtvp9B3eDuv/BuWUvyk9AGu6NdzfXjkRjsUrgUg
rOB2fjqL17wN+BPBW1vwGl9aZ/KhHSDyvtRYjT1FbXbO1WR/ki7Z/9K77cQF
NP2xWXt5G5/bYxGd88ggpT/7TUSbps1r+EuzQNvIrgrqug8crHzcWhvZSb2q
lphK4o7zXfNFT1ZFFH9g/+G/50d8WnfYF60F4WplDGy6nmkVqZCzjp8szKPO
rCzLvH3gmc+OdvVF5tNgkJuTje7Xq2T8OchVuaHAMlKvpy61Ve4UjUZOWFrt
cY7CtLQYEVsTWHwMbZ177Y6wXJkT2FEaolAc2UgztqEABb0iBkZjjcFKeX0w
VIkKRwu08Mh8INaEKoUa9rXOIneRhULXayODj+7gQkQzmSI+zRxnw5t2iZJQ
qnaOnnf9kqmP4/jGI0bSBcUR9WwpNnWiS6HjsN2rm6lP8qiGH/xu3WpQAWN4
LUaS+0Yd3oDy2hW5qp3zkilAwKJk2jhgrEGeBnJV0iqdBQyFPugqPknJ97c8
rLZUUiNM9CDATVCfnG3le3s/kQfXUXZXls4+NpA3GQo1iyfdGhzLJq9Pkbd7
9P7iMdPstDjeShlGN4X26RMv7zychySqFNcuachROXmSMPo1AkB883g4ta8B
JaHqQJ7DgdUlJA6MHeM2yxP9+R56w1VtfrQYFi5Tf+PmPH7yKG0hTFgq/lCX
zsz58iN1mo+gduToUHgk4SPJINtzpGDInPY8FM4tee+f0M/1TZs8++nEPxrO
BPvX1+I+yrrjIMPcSVUrdMufFB/32aDmYTw5VuvyD30ON+V/py2LU+ufYJbV
5cE03z26FNMQx6Q8uxd2xPwoygQk8txqIakqzwTk+msIZvyNFpv8LGJIyCSQ
J3L9S5H41Rx17Q1lHJhVfXUjGbBGOquFmfudoPj8tzs/2aC7d0KvMJnDdTRl
xqK5J51Lh9az5Tjxpbj30EWa++HNZRFZqqCh9iohY453Q4zWWBnCZzamUzid
fg9R6H+ogRNxNDo9WkiQ7LdK3qgdASw8C4XsNv7DsnHFOnJiiHYBBYKI7e3Z
ms8PA2CsgT4AiWKmAz1LEqW9UDH7vMg36ZCu5w0c8eTEDiV8o27H61N/YRmS
In7FFDk5mGjsgsGOp9noBv1fhByLQHbffOyaptET2fN9J3R0Dbp3E6hkud5x
GiamMDbX1/vEo5jR4PP16InDCKFvDLzmlo/Wf6TxST2HR1LeNVpEBrEDZ034
yc5ubnCAEZPfRPeAVWXQ29qVoY4wTP0uQyfBJiVyHB6kqD2bpYeYrjN8yFg8
idfbKwxooMNC3xd+3+NpD/yCTu5cxcILDc3B8ZF3qNlDF5tI8QZSDAh53oaO
UyMMVj6K9nRSMvOE7BEwGmjFI8xP8vkWEZA9WNcc7IR8XWl6iaZorwnWLMSx
GQz6i1rH/WSA/PI1/E8jpcGnwInl2QGil5fjzlP80FfMPUZOBFAwTcrOKsLl
DYvNMHRTmmyBDq8KuS/VghnCK+9+fSb7l7OsFx0QDFCbusuu7/2Va69tkaSi
fFQtZyfSI6PQSI3O5blT+EYQTO4G+dXXSpEs/nAEbNNaxMOAbnOGG1PduKFS
+atPSc/gXG7YB3hV+z5aCLrk0MCWVxg7RTpBetkehylq+PtRR7r2kewNsgVW
94ppo2WR9oUbOCqIAXBviWdyRa0BihvNveazcbDOlVHLQPgRua3mm7AWNjFF
pzyXREx6HUkIwGL8MEjEuCQA7/U9chIifZZSx08D5us24+akZ7uRcG+U8G/6
5G/G5BtgNvpHYLMpg7UfX+yHB6Y8dgOw9kl3x4IkUjje7yV6sEg3Ub2ditLp
fqsHtd0CXbINS4P1r7CDqV0o4g7JozUuDdfo0LSWpxPEqJLibyWUohNZhgon
GQ1YFACZOcBaxpR7wf6jjxZNfwZDiCi1k9VFtHsWFs4Z2EPnT8CcqXH/zu0G
oobqN/SrxjiFBisxW75TXY+ymQ20fVy2RmvK7o5RNMDB7FEhsF5Bq7jDpdfn
VS4odMpQeN6DM4LQf2u5MDOjmzwESCTANpouBO9WxvhHFFNQvU81/tneznTj
dCkIXLWgu4YSVZCBQTiO+ztJhCq2LPm/YRO4tYDaNKHcfnjG/soRkFgvVEWM
qwGkFHdQHZHDvp/oTBi2DahgEkrzfkrE5I9rdasQmcDwpym+Lcy6scAjpzLf
rlZw/rrPOpCuCNP8cHsN6Ljh4uTmksFkl6X5RiTBNs5faROyBcvRWh+dxFtj
e+/jm603etfGYRj4UU6v8GgxXfa8bA3wwApTeKX1VT2FxFqsvuKH3ymW3fp1
XPQs8ti0Z83nNAVWqULyBnwRwkvM3ps58E5nXmPXBklnPsj81JNaRNLhJlk1
Ey9bnXxswkzuGTwvoKJkrGBKmr2QxLe9wiNgOS/kOFwsfI5VFs6ZYlkmvpGc
v931aGT18MqhuVpGk05Z3om6h1sLsWelvqWzMiLAfMu8pbxoY5lIZIDcr17Q
VsKpb1vcVzcfaAbqzBkvjjdV4U7oJ6GQFssmibFKTZ8HZCZ7C94ORAT3tLnn
BqdSlJ1HG6XaSp8rHjZLRxvFBGIh6PzCMoHPewIIF/PcvbXBXqAM+dDONHeM
dk9pN0W9pIjxlmpRg5fo58iOZrTVHPH1jfU6nx0t2UPP+zmShB5/kJIMWgnb
OmRfWtmNvjm75u/cL4/jGOINleDOAcZRfMXdjoYlsJaXUKOzY1EnvtW1cBZv
nPFdekAt/xSoVdWVnXdz2v+U5PdgOZTbfvcvD9ynTwiFKKgmg/h4+0HVIDPm
PpnwUZmDOn6bAy5MV1Ccg+lNUHProIc+jDbnWAi0Et5e67Dh7A/j9Y/IcnoQ
u346kUx+nfhRfk6GcXJGzgHe6p/QxnOeVQBpVmGYcQZAAqD0Kx9MzKZ/Gv4W
pfSXP7irgNaIJnnLfvPUo9ywddPDtt1NFj9lQPxZgJvIb3duCMCEcYGDvCfx
mmoVmyLCf8jzgtovPDsi3fTxqHT9KhXaVUCpnK5dnBtEV9Mr8fCU1zMc/lEX
CthKdbopYNE7L4nSqdyW8LqkXwShoxGjdpJzBMiCkDBW5O5eEV39qH08xAmy
FIWW1B0qQPEr8OCKZ/0wF5oKqfXTmK8XJYqw0XY4wKMTb7YwpMQuEy6xZMj6
GWCI+cInA2bnU1UPx4oYTqAV47AqGrbhQqbaVod1lVkamAzhQCQvZhn381Qw
lakVJtdFxIsdV2eNEgnWv6PREqW5JgNBRhR+aRhfk3TcrjKhhypsaliaQ4N4
zDBewV7nN0JwEpbbH7r9RdmVnggip1J5KE9yihGDmtclomK/ccvcrFSgVFML
o1fpEfj9dX5mxxbvTJwZPURE8A15EeouHZWyWdF/mHLGCLPnRreCyEfSTcT0
04IC4f0sMbBntELyHYpqjR+6+jaPjZDSMVYzTBwxQXeZ3SAeV9YE6QOSvGL5
Gl+W5ZUDpPjJtC1Y7DS4kJBPW3DmTqEZ8+dddQnS6hYNwXW3p5uTbq0N5+OE
kHcg6nXPH4wr5d09g5M21KCc2XnawXehRCQCVQ1d8SgNVTjbFXAZRNqqdlTn
Lq0aY2HwM79i/Vif/57LSM77ynkJeiPl6RtSJOF8ap2X1woszPkXP4c8Giv7
Wi5NwkMXLS00bpFTcWj5K6PuwY3TWiTJEHmdqTjNzfTE3mka8qP30iutljMG
o8OvK71FYtt1lHhWELcn0XmUUNOS5RL9Tts5enm8jx0ezY9nXZNVa+OevzGO
Lt7bIqyzkmN9DLDjGymOwkIlUURZbKgFrU3XDSX4g5Q0Ww/2IYvjwt/ayb0q
Ok6VqYvzmLaYR5OCXMxKuCPdfU+GFLOO6MlEf22rEuILDAUQBoM0ofd2eoxA
aZylV95fZedBeY6iYxuI76xxBz1PUbURYX2qfv9ggTXXu5/yfGh+jdvX36S+
/wN0Fnr7Kbth3eqtLSJP06IgUxk5pSvuKBHZ9OaHd+5MHdjsnRD/MKpWSVhs
xbExdjOvlWqfYSvM2Y3ySZqbFb38MQGfXDQtC4NGQt1Po5/llJ9DFM+hhZ+7
ZwTRNT6L5NxGJVjLJJSludLshWenqQAXJpJjpegM00wMlfpFueovTt6cIpuW
Sjiz3RC680co5sb8/Au8RigXzoxnnvHkJvhGkPI99y2WRYBJ081p4p+NaOn4
DY6QpstKxgITZHPHUkS2vC3Uye6JXeHtHDXL3bxE1NyGA+WBsHSKySzvj8a8
iVxK/ARE0YLmgwwJhqQsR8V8VvzQNhH8pk+EW3Oz8UlYbNxr4peH0URwRZRo
GqDKyo8YKuVT3E1aZX1e8/QWJ+xTPyx6MZjUnIUYuXGMWjwP98rah7C90l09
3aRlqhHM83XFojGZ7iMin5iU43OpO3rnNqKX5fQE82aScFx+Bbw8a2LkYU9n
m+izAJVOOtlWPtSSNgGM6QVLqVmYvvWfRemCPLUxgeX1j6ntgVDJrEaSJdjO
b22gt/oLU2EF/Ev5y9LjV2P9Og7ROjHbM2wfui5Yt+sE5zT8L7aqYNqzNxHF
svf5ZKzy1LTrLtFq4jGJSVtcn+C6AgZLVk9LigaiMIMGkO+U4TyBF7vGmeeT
079gIU+y1aH/TsOVy/KAoNvtQ+6cy5m6+eB1PrBAKJD+0bcvNB4+UbueBA9S
awUJiVwf7mJrhM515HDVS1ZwzGkOyXfD024Ahp+U74+hnZeqvto53SpExlnq
/nTFB3AuNFYlKjFi8H4rP9ssGjrN8YpJpsIUkv4d3upNL69bP/RWNksLzql2
acpWwbSuhq9QlpORRqtIC6sSbKcYB6BGeiJM1j41vRy60e5/JeV5Qd1IDD0C
tnPg61ZHs3lOYvOIjX91mI4vmeFfKMQXPkVnL2PFRxN6fF7OLdtS6iHWP3fn
ljoE998YqdNzlgVma513iA29b7HwmX/bHaU1ogz8oK0DgXe61ZZZxTgPftCZ
RF/pI6p5Hc+KDquce2KS9dBjFZkCxIwehZo6/jSET5hexWJLV6BuM6x36EkO
5WR+jXcHYsQYFyceKnOG66yQzft3FL6a+CP1ekCbqWTiYJkwCkcsLTgmwohX
JkccAGgtA2iVAXQ70nD1DSwVR07hgC3PVpcVGF277noOed7WZ1bWDC96/MDq
vjpWFuZJI4dONdthAuNti6u3qYJb66E/VErGlqEjP0UnRZ/JqopvdZolCE7E
6vihTywDAUeToMUAmD5f8bykpLxCNELKbECia17Sem6kNOrY+8jU5FTZz+ZO
zlNa572HAcavnbyIAMWWhJ2deRhMbXDnlh6Tp5PTwcjuDlj/qO/TDZybgbUY
fzJ2gthV25uv11oiBgC//XIMGw2jVD/n43yyn9OR6bsKSpLeZw7667QZLiHV
pwrpuR9ZB+Mc31iXA7544BkeDIPWKfA6nR/r3irhODpx+ep7Z1kYp1B1po+B
vzJurEqdbaRZn268KGqG6xI4O3BREIF9cVbXjqdfXsRbCXAWaBZvMQMrvQZU
b2yjvUj5YhWXqLKD4Vh1Y+DA1hKhBsj7yRReJk/XJQVL+ROUjEpuDEB32IfP
FZdvwACMHiLhHBYIY6VmhHjnZQhKiuM+GjG7yIvkDfYxW95rkiL3E9E2TQVz
AdcuVM8QfewavKFqqbMKlIFs1NK66gsnwa9INYO2m/DH7byDmzmuif3eI8mX
aprorZPG0ALlzP4LYL80ype6UXYl+NZUoAUsIiS8XGynh9hOgMCDbZ8DSkKz
K5I1smSUm8ziIrUPugJTxeH3Kcp+LuUlGbqjLMJx0JPn/L8gWF/8cSEdnlUX
2VmpG1mzJZ9nh1DgiaHBKnUAnMJBeIvnXLY+yFzrXkjn9ekETpcCYYr/iW3L
niSAoPwgPsMelv2EqitQp9gJnt+EYB8kswshQGcGIkpROALfN9bJB6SOnWiy
lus15HcKCB5k2OefYc8bhmjTTOdK6dUWtbPMdZx7fHxBjV7h3JKqfFxX3ZIk
NNOxZ+TfvFqRKyOxw+jxQy+2jniPi25bE29oJP/DVWMSgd/+KC04uoP3+/Yl
pzF6aOuyMiEbH4zdKaNEqyacOX9LIeVs8qibfQ9YSGsz7MS2LxzCFr1t+4NU
xCd3+igU0PKXv6Aip/eU+PytwpYZ09PEZn5j8zcT3RFyAZkY2WJta8VeJoYa
CH5TksfI8UgiYryZfq3+pAR+fJ71gqo94bI38umTwTVcbgunmjHcpx0sgbNo
45Y2xsXSSih/JDPrepHWZmU1/tAnJXkGm2/JCYfm/JBLotnFKiT1N2yaLplx
tir9ev75zhvKKdilgpRy98IpkhwNJDcWMeNhJN0vD53RcRaFPh3HM2kz2NZ0
aW8+s+x6hkHWD6ObdNCk9l12N5L8XuQ4z9GgJY0h8iWpimBJi1LM7Oz+6iNT
PbW/avuw1tIY3zJWmFmBRFpp3hhExYJSd1uhDsomWWg4kViDhV3dsLG/MVJc
mKEyrpxoIPd61B8QN9CaHtdCYeRUfgkZCQhQws0i8h1zi8nC6ZCESGXa1ftN
AFcL4cWGA/3izJebBM0M2H3ezGuInFTtoCMJtZk+cAFU/cpZtPjH8axbDMmo
WrtENPdYiuNI3uAbYtsn57NrMV+sdPUzz55ZsGpoUzxOovJI8GspD25EPZ4g
e+9TvDsDtkOQuCG1iateyPujASyueItelApUAEmMmreITRHOaJHMUcdUcyDX
SfvjAEBXsH7ORFoBY4u1BGabd6UUE7Y4Sd9fHGhVKvMLEO6gP5fBn7Cglwm3
3gZu9slCDuO8m6ICuYUmSG0NsyFptkHgvnJYXs8ZyAaHc8TFsBS+slLGipHs
kDNmn5kXaS8S6xA8y2DJIOfa4HOt9DUvbEfAFL8WZTi8UwfZMBPX7dbxXg4V
GhdmqRLyFLzdatPG2L6sDaJXG8o6rEknzu9c82ag7yCRvkMhK2JqhuhJC0o+
ODOa2Fns3+1zuCQKNqg2aRGVgW7TPtR9Oq8j2cPhPmXXrgvLlR4kJrO9mRjS
dnsQidmEGyQePIN6h4qOR7QhCM9vSpmoCpC1MQ1yOKUEQDxnhaafoX8tZQXR
28K03ckgD2axJjq3j3wppp5DpX0nNLVXF42mc5QHko2RDMMdefC5UkVwJvWZ
vP2EXDq7TRfy0ftFWyFaWAlHpoFPuW6ZCtxPst1+Z0GessWirUNgPov0OBlI
0R9FfSsWs2XlsZ2WqfKl6uAEzvzvB38uX5fuEn1UG+7c7lZGazWW8lcIeE4q
1hpQwpFHc4QHrGjNj/Hal7BzmOdKl9P9QBrO6jsKi0A+695dwxVJ2+qb/NmM
4x9ZmPtpVuTUB0T2sfgiXzNVyELJfYUREfefnjcgcQ7KLgInqsAQYWizCLqH
Oebx9rvsf2NDegiqEPYUS8fNzbrx7K6IX0kzGjaCEN3Htq4IZpaVguk+mXYi
AvuWdlPzA0j9SSvPDJ8asaxtm3n7Jc2a1aft8Wvx+eOGm6t90lNhklY3kN4x
KSATQNQ0e/E1sAuUUHScndPEfWFjT3E01+Acva/L5qaK5Ku9vEHOMHSaQ8va
Ryl3BvL/BrYj8fLXv3kI2Hb0QJXWIXdSGrPObQo3wr9kGVIsrJo/u7MbE0NN
ysSgUo/Q3moWih9a7t2mOGOjIoPOaD2SsXbvLp8AQnVxQLGUw+Aa2e5mst1t
tfirSnjYlqanoT5hHNmwVcaJEGXwgw/xhB73X1jMgn2gAhLTc1AyGJT6FhEW
sirD2MzglN360C5+1cIsoVbvb1kFWPsok2f16fhG4ccKoBoFKDDdH99UabZ1
pmwUmMLZZnND2wd3SfnJkpMbT/zWFvFPHSwx8NvkmdYdXJYL5/jsSb+1XSte
cIlizGnhPwXc2O1c/svQ+OOlZjSih8FloSwtApeUwVd/NkDrdVX+krzwpHjL
FSSRKab/Z6CAYFFwObJ85b2YW36xmcMJROzbAGo4xXV6PV0sBR9kboIIyMzJ
Ftt2sOrFNWPoCgh9XIXZmamOteLJCH+YnHKot9GyoRSpw9Fhq8ULSwWpY7vy
Dx2NTbBgd73/oNzNl7xe2NchPUSw98Uw+bscS6sSfWqhcScNFcrzzZb0v3Yz
dZENUJNcPwkPZ+KQVbiI0Ngw8U/Aq2wjM2r6mdB5JS6G8O7s8xMgToOqmAn7
jyH1/tzlENtpX0SNegcOQ9vEe6D9vQOkbHTGnK6VD6Mf4rMCX3nQ24dksCEp
ruavj/ikVBdQVG2KuRDzNkduqiazwzRqnGWrxPJmSfI2hN0goJ81iCStzmaU
xJ5ovB2EApOuRKSoYLgIOJBcMoAlQekZ6PB9NKVtTS8rkadR9tMOkOorNfG9
PMNThWGZCdR3VCT8ZF+qqt12AaQHsYpRtNNLOzd7hCEb8gvsxIpf3DkkryUi
1A9z+lOuzoZNixFPr6L/UsMl5H3uXUxOEH5vsfNVfmJuL0i1khQb1dmGiFdB
VcuNdJ+5Nqu8RtNe4ypRSO80WUtc4IJFKo9pvN4XGgvxOyHB/qd0jp2Ita+D
nnKlaa5HlkBneJZ3vl7r8VvXbeI6weopZJieUOa2FweFvK3BvVCpeGhPEnJU
qRavBcywDbYUX9rnY1uZhhRIRpyoBpLo02TCJftZc3sukH64fJLfDxGn8ih3
4xxESuOrCtUfBXr3U5RIDdXvIeFNAAIiJv3Nl7f7HmZ8yZN+sLVhXLGD6VSb
EhsPjBW8stop/zydjSoaNE+CiCP3LfIxkN3ZdQ3YdcH9gtk7CuXtwdDW1xOX
N7MN45LQEWWgxplmje/8WEKeVEaLsxdcZ5f4WCKT3uh1XcmHZvx2mEX74oI3
7GFJQEEz4gPfWUkBh/NQhhkYSYZCqhbkP+d7llPPXgBskTkogdP9wxbUNvLS
WXG3zd1XLDPzG3T5B9CWJ35rHUx8IYvf1J5yQPywRwLs4pFWQBhuINA3KOyd
BnVWYGO7tSSEwWqGz5CWrk7mX3GZW5ovIkKThNx6qT3mHM0fT5Glra/zIAXC
0owl9breqa3nGARGR5H4urqBfdcYNwy21BQf5Jn89TcOShNSDejspZCTxtIB
3RmUorSrb6aEKyM+T2UHFVcDXMpUVR4cvvSMrgwPfT+lywW4piZHOUlLRPPT
TO5H5YFJaKIVhgaXQhOvyPrGvRgzKhyCokz5mk101X6/QF6qY4W1dr+jRRnE
kV2sk8+rXalx6vjCJf2A3NjIKCz/1uqvUrfartW41f5/1CdQzrojBhJUFVUq
pjnTn0yo0SDAKS7uQrhd3IRxX/erSlKyVSZgn3dS1/ySZdhr1BOA46i1QEB+
xqZ/pXFkTpam6bTiP3hS+m7cA3VBiz9FHNvdcSCxjM1/1u9IK1pR9aq5Qcr2
Lvd4d15FrwpNLZgM8IgEF6Mq4MmOL7x4b7EyEUTKwOX/WFmJijYwuFU7lbNV
Pf2Zp6iGjLLMXNaW6HWQVcoA23sv5mEspKZhsFwY1yjQ3+LBcHe/Cj+vc/AY
F8meTjvC9s269X7mXiBakFYIlmllRuvqbXhj/Bzx1x0KKiI5fJiCyT4CZeeH
1pK1pYDF2N5zeWHLcJQMiqYs0coWltSvKWAAgxUGdnkey+gcXki6CaD5cMai
YWwc9AXqo7ZYfm50l9cucbtYKQS2v4VsmhfyCkTZIrDTxMkdWevr2nMvMHos
9C3rOhBHXoIAbn2+dLovayZnkcK8Wi6g6nVTTOX3xzcUH20TFB7mNip/FYFV
xZaencA8ywKiATLvmUqwL7Fogb8+dYIKkLGL3ibTI2y6Aq7/OYqUjEJ6a5ei
Kf7rpZiYD8HX6Z5+HRUUqGKtegvs8fP/+m4IaeyBPYfhnMLNJNHjL+3JlMtA
qH+/KVJREV24YUw9xzhHxoGI73EkmmRDG2DdyZ0Mi+1QGZL53koyWR4N5yJx
VMCqwLoN0kqytD5wXTEWSpaXlyp+97WKDR0ghSuZnF3BU3asmIN8OEdcfhAK
N5Hv5Jf1cplDhdYfc1s8savb/6f9rsP85OLLHQ8xMzjL96ww/cPERCEn4Qwb
XJPolGAzZ6AQ+K8W8lNMZ0/sqlYiZ9rqp/m5cz8eg13sv+kKJw7itZVTKarl
dGJGYGw8vURewX66ag+u9q4nZNoQleQZtC73vDrbhyI/9bRoXzYTT1U/++Ta
Q45/nDbPBbJqfMODdf01tEngjKM1iFLweyB0R4qX4jNW6hfu7aeU0x8df5vP
h/ZCzGsxpniYNObkfHxtMt1cR3j8zZHo3mdeWXyz4cefTShtsWkjproI70YX
+SZIJZCCszgkCa56ilp1PfjWJZDpTXKk/xaVMaIDTfWxdERYSPzuSAZQG7Ph
f0J94VvpXzzwyB1w/+HP6oBKBUCC2Xa13cT0lsxKRvtK5rqv9Q6+cE61V2Q8
Jp4IeNvnmBpm+PVy4qsLiCTlJNKahRrzd5rnIM48OxMrZDMAJLsf6gnlEQc8
YgXkZBkg9w19vqaq/nO2NYyTixFqqRSBqlR6Rsr56b9jY1FH+TyLc07l7oXh
K6N/3c9ZgqR8JlmgF1oiTvOdoz5dQ2FuKDpIbXze9Ova24vfBWAqBDYi8aer
LSSuw7xQmN5N+/OImwIOa4d5uUWjEG+Wt5dB1/H+XCmnFqsfCKr5qo64s2JY
XxlNaV1MLvqZ0f3QOfIxz65IvcuTzogRO4mQWGcxsCpxEpgPD1CB6Fg49Ygu
BTHfc7ftGEqv4FDXY8cBzqmsPAUzrvDES3De1SH4rVIedeqNrCGGHECTg+4c
aKxpbyfttkJY0SdHoINjYaJ8pXHNtZVOGSjJEPP3h+DLz1jrWR/YlBQ2hmh4
yzySn4bgQTjIq1v/urEZmzaTXFapDG3bj5uHTeumDaIcHdyVbe5RmT0Cga36
r2XcOCSPX9sgKlj9wr8xES5JQNRYxisDvxL1eB2iwbaILKzabezSbCziH5Kg
U70S+mompsOrSZHs2Pq1rpKxPNwFfdiU6gES3698ce2/uLLAJmSdFEbNvgNa
+sIFmZaliuDEca8EvG0y7kIDDkv9fqXgLXJdyGxc2NWNW7RZMwEh/MFkS5hD
TyUFrevRnMCQVjxh3UkWIByt0ME735QeAAXTvS8MU9Kih+QCkyuoKdDkUs5p
Xl8L++HbdjXOefUAXOGmfFZAvnZHihY7eGGwRJlV5OFSK8ykAuz85pdnk81g
q3L3e1/DdZe0eLtMDHHRD1khyAT6h1pRJta5SkO2+JqTFisIejr8G5+I8St5
UsK1E4vtnLAuIhje3G9kFMU+ipJu1/dbeHeX2toDJUzcFz7/fXpQamFRMGI0
DJi0gJf/4jZn4bO5SfnFyX7ItmDrSnGERUWhcTc7SO5PJHz5f4rydZwfZmWB
DSbXQk3xXV77MzM+EI0l+AceQIy+dsW5ocqvbE86EjztDw6tCvK5nR57GiCP
t011VJr/60oS6+yPkGogzziRO3N8YsahBv6SodSUv9TuadrMtQcZuWZYn/KP
vqoiKkVRhUh7cFNI6TXlIJKiO0aPXHrQw7XTur2Jb98dF/q5amPCGc40w27P
Y+dvw6NV67+/d6jQ0EGrxU1gLfZURligb5tr+wVxshelsWMcpvEB3Ndmt11K
yScQT2hvBhFMbeh49kM8dSdRzJ6AqRLMW+og9yUcafHCSMYH7fvf77b7UBff
raR1pXYYOEWMXpBw0+qypkONN39wwXaJIYy6cU90R3Lt34pXfLUnKBU0fqHh
Y3qz/KukhyVnW/P0m6XG6o1JHybjnTfift41WtidCo8bnbw6gGuTEQru2iEJ
TlObQk3TIe4qXpecV67k/5ovsIrJlm0mSI/qukrQhSs9cs3Bv2EB399hdq2E
8a1WkfD+8D0UYl43jIbB3Aclm4/uzztCrLj1FTQFjIGg12N+dxGiv7Hf5uRY
jRJRNA6S4cOcZAroxFuMrWVFDo57ZmdN9/s3NSc0wz8hQzAj5ITeVlcwcHYW
ampyllTKP8/wC0s0VXYc0mjIrNFhn9om1Gjr85wZPtqmR+a/m7k0Cz/g3rj3
S+oATXg4KIzRU1v3hlBEFetYF7lvndQ+ZrImOybOiSRSQ4492zH3UcluCHlp
8FqU1icN1LL189J2IUFFzdZgbvuCim3VUPPmAL0BDpqwGQQ5WBkg03NGaGD2
0E+XSbgVnYWgXn7ycfb91nB/orcQIVm4BXtLI7c4majejHb3wWz9T1j4DfHU
u1Xx+OeLIaVCrBzegKtFO3+BNT50E8z/UQaDTKbXcRcjtAonBlk+KhnyRmnO
3Q2EuBa63MZZ9v+mhMh8vh8wZAKeYxAUUdWARzfZ/BIL/1vpaFHuseSycmh4
oTjpyICmqf21cPKBhN/oeqTh8EiqHH2PRnm2bVsjBCaFUPPXTtWF7RWfQkpc
i9oAC+4tfM5UdAEurzHNXUWqqdJVdmvzDMm38cQT+nhQb1XNfCK0ijkliPLg
3xs0FPMJiLkT/6oOFFisOs1Le4ez90lDQxPPkicjgwhC7HOBPDJ8bPHiFGCS
7sJLMtwAgDPdKssVFBHymLHUIV+Ko6fLUlOJ8FX9Cq6/F7AALWaVi+M/G2ba
q3EDVC8Obtnn7z+0BX+Ly0O5YGuULkMMQos7IbGpIYEA0yPBwcNbIm3qOAFc
ihtzUgMKKEfd8HLlcoXFLb6WrI2nzOn71NicLJJSmeLmjuenBmhzQnfVCxX1
22oZs+gOfmaDxeNdugoA6eL724aBFLofrvANMEAblYKwGS4mz1iiK9eDHrks
AhJyBtpYCLnUVs/WAKXWhy7g6hcFCGjBv+6oqOzHQONUPEwN7J/Gbi4m07Op
JAjRc1+obwBzPL4j3iq4Mu4Xk94KCMol5H0mnjOMZuxfMTm7fksGrxk38mG+
lxBiD33Q1Qml12Wwt2NYv5EjG8YLtvgV5mELgZqsSxYd4PSu2jXj4g6OxSUq
M0o8/4gWcLfnzveXlI3XPwU0nzs2Hmy/prJ/1raA69nAT7dRgm9DaIUmwrDb
BPCAC5kP/U8etaWBQ/t+IHz+PaZTRWDibm8lJPopUquLwFkhPh4GwnEcGHIH
xvbyL5ahk9QquCA5SyaJYrOoalqavGfhcE+XNjA+n6uK76fS1LMIV/ZQcYuz
/7Ony/AoG8WZMxrwxRSZPDcKGgvVuRlIvc7WZXuj610bxA0wghKIgV3HfFUl
uhSugZRwP1WJBoAPclD2NQ4ki5J0RSw7wrDQX6AlUmXBRBLdk0GwVdubu6/c
tOhwuSuvofl+Eb9AtjT+F646m2LUUGpRJuvRvRSYDdfVACCF6O+gUqESkGqD
ci4szGYUGnDR/jZ9xTvOrPAQLvnsO1kASQxm/Z2YfLNtmYFzm/2P0BTH2zoC
1MEdinvV4gLuohtZvsrhpTtBFc9VUoaX24RB5lhBUGv7+P5q5lXKvtGpwqV6
+O86T1Dawabz8fcldyIr1Xjgz2v6kDb1A7ZmkgFfMq0GoQXma48xg7it6baU
G2n8rVUhUfLKUoDO9tu7MQELSyCIfVEBjuwUJk5/7vUjdnnFbv7BgBnb/JHs
buKGnJd3y10c1k56eLp7WPibHBtoiI7TGEq2siqqcObnwaglBN4HAwsMi5xC
Zl5k7BJ97wKvZLTCmalM7qnIjxu2Zp540DpuaPf6WqCF+YbhBxL7DbM2KvFV
Y2pxxVFciV9kG23UQx9EaGVT2+YRh47HZOmr7gcd8zSKCtizC/3qgz7HukOg
nYhfsyRHbGunMxj2zP5rc7E5S3L0FfGPTYzC8y2OKSJO0JKSC6RAwyk8tND9
hUcK036yqvehDQZwMKTT7nXwlfFMie13R1rfyB0tS3oziJGAfREYO+KTDWPp
U+x9PgfV/B/WdSYj3wdx4O7xOjrdTelibIu0FMwAb3sBHLJf1WIaSLdA/Akh
BqZD1+pAu4//DKcvCz2QGtTEj6waF8aRZ3c+o48aarIWkWyQ7oE9qBH4/PRo
InNqGjQzBusd86n+QDj0NxAuoAOqIchbL8m7FiMQplQkdr5/DwH7jHCFnbEi
iIumuSeC/Nf1/RllAiwwaIqeCxcuVOT/FODJxrHch+cO+OdD38EkjyZw1Ycv
MazBiiBGexfsFHs31JZWJlGgJ/6hT0w32snFSwfEOg6406dVmX8taZLiX+B6
aNL3y64LeCJ2TNj4Lu6puzi9AcCMsHLk+uV2HNrX8FFCeTVg2+9uZBQ5qCQg
oYODuM8btwkAzYdCn88YZqsOtHhZtFz3DQ9y2zRYwpd+rTGG6jec0q1VEFCV
tSENge+i/r+9NQB5V9NFaXAkc/wayCisflvz0clufLR0Ph0PvjzIKV2QRBPq
Ok+XSAvhUpgpjUcyUhNxKx1tdPDCTpXyxWK1x0k0LpiUikf0qKDfvZiokrSI
842AO3dkGGvCal8Q3oN+LxMnso4VlY7JMMfcLbuUT+iSuWisH239nooQleDP
y9CnvuT2yOkiAItfddhgdwoHWSZouE3ttQ8uU6Xk/OqKo9vRSi4szychkUzG
QVEgJZ9WyPi/C5kPEpq2acODnTXE1JVYvZeoV9WAGV8H9XHNTVeF7CEih8EQ
arjbPzJ3QuQ1eQ4dgHZeHCrQVFMRziulZmxk802zkAnO/RslSNXBoLFNi9jx
sSAVZBdufxlWWJDW/bhqb2Gh1LHDZmAxdTkgoEZJRBsuJhRo5sAsswwxPjIS
AgokI2kD854Hu8qKVNA60GXt+pO6/o6IldOYzIpU3gG+JmWC+RKenrTCK3f7
s9wryq9lu//J0dJxLziK0ZyBKUe1an9ZHEXQCLXgCZuNb9cD/SJlIZORbF6/
qmg+sXZq3avLhA6egqUDrzild0wxN+is2cQt63WPTRY5FNO9S3LfKCk8PtEl
T7kJ35Fk3fyhbLctnZTIUKhQusIZBKR8wWF791ZEh91k12L92vsUOON+tIv0
FA77CVl65ux1xCI/OvU4CB2RWlDAi6O6AcXCUw7GMeZ8AwVWidkJGZBnkAQg
W/PqGRiJRAmIJImDXPY5DA3RwIrmZK9ffWKm/7PsOwwXllkXlGkKE93/yg/o
8oH64hNgcon92CjHo9XlFCkNj0WhVSyP9km8HucoK6Phs6kWhUyhCYNUiSt/
g30cvfZ23o1PT1tT0s/hfcJ6hWIuTM8WjzSO+NC2huQe0q+LP6+MVRX4C6oB
rrPKZdOy+Ts2MwyldebpB6tRBqOE0QLv1TMpz4D4FlaG6pKj2DLmGDCtzlPC
SV7OcerHZwvB0/8LTEdbfsFkitadFDdDc79BBvpgQD+tlebywdWWcaLJJARL
FCiqx3xHRnNnpiWlbGwG/LMvzXsffeNfGoicYoKpcimYff4+INbp7wnuLF+j
LAip0V14HJF8FbNPZ9xZT7lVDj9W3lrLvgVim50yXisVgOoxMHUCVisveanY
0dqDBhWA5LTQEJSTNYVc5AcrN/lhOGJuoIp0Z0tkFzZ+Mqafb/I4RPrIXcHE
nA2kwLTdiruKs0HPvucaPYOsNc3txUbA51GP2vrNktsVhgh3ZpHX4lWNN3Ns
kiJTSDWOaUeurc8CdKhFb2P/UjpJxlgWnTSnKUarwxO2PApYv8qI5FCG3efv
yB4cwZ+Hp4dg+3kzq2lf64wWzeb272QxQ9uJzxsr5k7mVGmOlQkIIkpSOjY3
0hVZV6V8Tsvmac0bD/y2qyam7Mx5KcLXFBpF4520sxevAP0paSwPP+oF9Tui
SHlJAW60aGW/gr4kGfCFO4eZp/ZDEueJTcOVkriMEF0ilKXht7t2EGx4tB1k
kVJP9bXlPYOUMhyqYNXIL8Qxr3npkq1TTNjf9d2QLNCPLyBt/PREaEaWnQED
xR9D5T1HfPCcFTWfI0RcuDnD8soS4YBbu+GQgVd7z7jTAteSygn6xymIqfJz
MzPkCdTXNk1Dt3mVSvNzRmB0CImFqWsgMAPbrTEgLtAnkvljIHbrvZmZteTk
17yK2Y50biwO/8K3J6YXbkAFeM//jwkd17GRgJa6XPoudWcKHc8fr1mn9BGK
XCXMfriM2coGPX0cFMtbeitxyBKRnmA2cIbVDLfbp+NOekSGRVdn6ZIVvtf1
bL8MJnpODRUR6nAB0mhR8F7vEb4plxu0hS3JUgTF6di1CQoe39tyEhN5gdlL
rUDmOCBf1a9blDXF4rTwy5x/sCa4BRfye+cSNCQvkJJDoShA6ju7pztdwJqe
RMpFnx2bss4Fz6/CV82WSHEmYFC+feGnfU0djwjHSsiTMchPDzEspXuIeMa1
Bn0qZT6YpmLojPvVrL+XXBwkyUIUklleaERp2RHRzRyO87llBjKR95TtktVb
DsVu92IZDOt8j0TEuf1/i9JTZNCH0kdoAPG4iquhG1Z6DhivBhZzpUKTnX+3
pktfYZHw6cL1UP7FzXkjKc1i/PjPfBaNSJ4FbUNoudVGHK1+wHhEuy2WTE5Z
tFDEdmKQDsiaPIy9JNW4W401LX9NEzQL0dBJjC7IcoGTQSiUgV2XZyJrJC1v
3y1m2+TCems9F1uiHoCFYjEqlSUhrBsaQ4WA1HxRdx591tQ8VMKmh+nuD566
X3DCcLBRSEAsXCO6BFFNsECvdr6V3mToo478urLsk9X6ommATtjzDSX3k8Y3
zH8bqXyM3L5fIxsxLgT4pZkWPFCWKWGqIGZU8lKyLh0zByipYcc5AHr9pOch
HhUX+Y6fjfd7SEYhnpuK5iOrmXNRb2NmkJOaBObjYPsbB0pub4MtUIqlIXRy
qmEeji14C6TW6/HHpmcQSPQXnZMrdy+jk//EPe22UVuttGt0SSkV7ZcGmbIb
e2nH47ZdPJe+Ao2C8FEnHIbrgivWQxzK2i8yC2Sj4odSju4xu2z0FbvtfEYw
PLbCag8sEysKhwD4pDN4d4etqvILr3Y/sE7e4rMzCQ0HvZMhs97517SGtm1E
npFkLiWFIbYGG7b0hehWnWTtKuzneQ3WT2Zb1j2ACW8q/iBtBNZeeof5+MKn
BY9zx8d3IbMLmTsmw1vMz4RMjh8JZXqW4UnZxFFuPZIH9HgpmbCCrsXjXks/
zHtChnoxfJ3SEzlRohZjlXI4EO4dHB1Mr4yAJ2m+o0ee1vlRZV2XKB13NP6K
43Amksbk2zHhpUCx+qnluaCp5CS6EZw4PGDol220+tCEJATPe+Mb2bYBHB0X
nzrsX9mFRyLVqGhOyxa6mfKj7OVgmzzlLqcCDzRReLZEdm7ydjoQ0hi1gGMD
fn66C6ZNuWTQEyeP3K7tOGL2Vr1wFzontmxxyEB2Z4FE59Rlx5eDilv/yvnD
PTsLrN03n/BWxoIk14ja4RFg6HaDBeeuBhuNHA6mqZjmFziZsFL5hz7h5Apa
2nhlcFlwhbAd44Qzv8iP57abpv7Rb1gRKr9LvONx++nGFqxU5Y5jBY7GjJuB
Q2uEhr0jdqpUbp0qTwTQF0YmpGWaUdoahuG9EUCFiWK4QXfIZE3ytupGBa2W
XBc54Ucw6rj+ubaxM5pTTrdr5mZWtSyqgVIPuNpKMfwQKTBLyAYxs5dSf52c
A7Zw0/ZsvdZb7+1piIXt0aLQv598d8RN8jgxxjf1yTcn0L+VXSG36IAiRNzd
el5F0mGL25f4YgbtztMscNoFHYPqRpMhaI42dqlb9lR3kViNCYpWkq6RonVz
0jRjgFKmZwZ9XVpkFb+tCJNrof9oriM6sSu0Djj8IQKDOlgvuYAwg0tumlB3
araeG+CymIMNUa6LgzJKfclGaDV9isN2HNCwlrmDGeRnd/EvbUbsEooDNsjs
aZT1Wmll462HZ+6bDCD7qKJjWka2i2CFAx/oeLigmnGcIUyBUiecmXXTkQ6w
8PywZqu15QSv81yLFPdauRcUXRbzU+V+fAOp7nTGSvFV2e2fl7cleYNux0Hl
RzOlTm/CLTbPp/iCR9ZghGs6gIuFJjrGhSv46HtJEhNaChznaxYVka5aPgM+
Kj70OvhUQpGBkE1vJNuJmOWYDYpCVJBCNM00yHqH2wTaSv0iuknUGdf+p/UV
wsBFavbTcTfw+D9LpylQJiJ4jrQNZ1IBtKqFVxn1lsAu82Q3qamwlfN+Mtay
cGthOp9y4U1Z088sNKyClpIKxh2U7m2/gsYXDI+sOqBPDoHcbvb/5L36VPEN
pRsZ2y9+Fwbz4FR20zvhHzYwR1DqBOUDZ7unYTgNr5G9/OjIpS4o8Vmt5FFi
19kKVRLyaNeYubjSBx1ky32ITkCP5FCer2EVipAkqd2iSiPXk/Td7u8o/9Sr
jTUaeXqrsnMv9nLT+EtAFVTk7n6umZKRo5nfWcwInC1De+tu5GKM3cmbxRzG
Jb8tzB0M8KixzBaehlMw4/duSHW0X6mGpR1Yg3ZdckO0aavrUuxQu7hTyBSc
WPNMo9wbnO3kP82hfNzG5CRNl9BKPnY9innySwsfBNpbjPSpEpvJMZn5dzwy
OatU06iCoX8ScvQHQmXifbDyIn7AwN57re9fF4oA0qa6Bvtk3pW90CnG1swT
RYTldJm/uhWrjrFBl73p1UJWko5iFIp8OyHCDXKw9FF/kht+vf2hhSe3/Ylb
Z4I3e59GrBm3tk7hPkDyzkydciPyPAx7DrYMnQJ9vBfDNhb1BF/vcFklqLPY
s78hCiBG/Vjqupkg/eCZVmhBUnqRGLH5iwmBkYJKQVC7FyOhK/nNqxP+91xw
hoiUlLcrZDgPEj6dDehWOKtjGm8YkvuYmwihWYG6dktyEs+tVlUajfUk21TI
MTMjKXFFVJbyYQTCUITwrtNN9QtapXYoPRkVhD15jd+CfML83aWmu9ReMZLj
ct+Z5XER7+Xw7SyqDIba/Os8n/ep2hTJhBWRR84g6by+ywFFo+ufXWyXbeuL
fMp3DO79FSEJTBuVy2eRt6jEQQDRYI/qkMRY9vQa1gMJxLHfOIfeQCm2F6Th
AwY4SSdM9UDQms71GS2kqZD+8eyGDIy7FHhXEC2MICXA0TYkc2pcl2dMZ6Ui
vdw832mwJuKDID98jU86exTOENFh5q5IE8opX7Mk4xqXwS8IgrjAiaJtrffr
sX5phNntzGklR+EkwsjpckudS+Mep1kuL+1CRDpz+sd9VlnysQGMmUWDslZx
NNasLMu69ZASApJO1kdc3Y7zLPCD1y1J7ZIDb9aKvcqmOzZsyeHXgTgvnatp
VROwT2xhxurD3SA3X9Oy3dwG5Wn8JuqgOkvYl3K2czw+13y7FFDt+2wyfr37
c2MT+IxNwYnUNacf479wzRCWYLRM/ciM+AryXEh3tjhdxge+VvELlcq/2Zey
tFr/r33st4aIUAAewXvlWuX9DiDqG/r6G0LRnsBX7R0hqCNAqy73cKsalkX9
JifQD5nOscWsuqH0qVaWhRoIIi2bymVv5Fqpu6NhTpPbLrOXcJRX2RVeTCyk
6Rik61wmldplblGCag5naCYLocO/fvPfYqOMxlYqmPp0d7MMBKnOMDY6EJg2
Bj5+r5jTTF/BqvuAd7t7WmF721EJvovuJ1IQh8RzJltPwKbXczRDiCf/F3Ei
0DA1vfT27KS+KSzobV3Tm2DahAUCJ6EzcatRMf+VDjZyoDxAnFaHtDBycAzJ
ha9zgsYg2S/fCrCohXpic+BmUlAVq02fPFwWmFtJ1BITUJ8eXCnlblHXzbJs
Cm3v0nF5FKyjwgfJ1oOmyAOX2gbj0xVpbVWbGYB+KwrjznTdN57YjwT1bvNW
deH2woocj4boZeovrXxkJVOV7QuLVnUY0FD4TivyAgvTjdfyuS4pa2P6uCRF
F02IhYxyvkC0ENRbvWjfFLQLBfP3wzympQiGl/3g18/7Dki93hl4QDL4aQ5X
7ATfKaVHviVlnUNEq9ncMIRSpidBrZAyCM0gHvJ0P9OwK0W8qfT2CK0gc6Wu
tpXJcGZf9mCMBiHJ3lj8VILTS766Wdme9D1pGLYGt9m8tj7LGmoGgDLEzSLW
gk9dLf9qy34Rf8t1JSUkCNGJqzoixRewFgbEkyt1XWI3P9mZDti3Y6aX+vzh
utqFXO1M1AT8pg3IK/z/meh9KSbfUTRbuZ6ujmdvr7QhzhLHJy5SCNJVG3TS
jMzgAWbC2pElfMbrybhqtn+ylsR/dTTZrOyVXqFa4ILu5t2RCyCYjgXYnjUc
E+G6T4V0zPa7cHVg+d8RRusOQAL7rSqtXhBOxXt9Jw9CKXV/PbZ8AF9IH1yj
xxrasH96B2WAOYvdGF73wkZljqil2etwmrJAdtv4UeICPbSWEkKAO6siZufx
ZWBvFQ/1F7lc2QPv4Kunb5VWXwHVtlLekFrB1T39pvVNXmMBiqGStia6t7GU
u2J8I4srL7j+1XAea3wq4ZRZPADndOlfI9QedRaWR1/WB97BDBD8woq6sgez
IUywA8axm6iahiLlneGUOMWlgdv/v2vpCwDD4yfIqlGtzxCiEoHZMoZKCZBt
fGJDLMa+/qHuIWcnGG6EqxGjzVfKI2NCYXS0UVx28LkRo9s9xbA/yFreuKWS
rKrwzU9WawJBiF0FwJXCv5VMc+UZ9cR19mAhrFyERINKreWupMKPGT9xG4wr
aFSiwwZFjsT01QXzrbBNPbbw1pUm9Gga5fVydb5VnZ5mSzR8QmXxvx1d4bVY
rdo0uB27d+H79Lb3ujnsbAC2zjj3CIK4MKGFdgiWYm9TM0mkdTHeY7w6woff
Cg8jD0Z6VoiI2Dy3gVNIQALfPMBAk+BocrZQgN1qrCPlm+D2l6msv4Wm+PX5
Jr8br75ItY3h2mw/3H78q7f5eadz9+F4c5OERI7+h5XU6/FC1sC0bNOZ1NQu
yfc5/ZWfWVIjxtOzaI2vLnZXLSSfwWkEoqxozngQJ/IHfyEdxNIp5yakUfm1
Rr0Vjq7vXszMXCaQ1BZycM2WwiQemJ4oYJBlhiPFlKAwxAAyn61CgKZjDqlr
5z9jBJjoMaWoKao7iMIuT0nUfB4B86tjR2iY02+tOwIg5/HlLV28+ShJe9z7
+3Py2d4cVp/oESwsNWQfGgbV9eYwIdcWsY+bhjKOg7hSBW5PpnGJs5i2LQuL
LbvPfN6DbA1x75r8hIEMO0kcOqjHe8Ni2nWKhP1nJ3FW7XVcJw05D3xregnH
zG0TOJ3nSW4BNgtTlglov6oXpeuTU27SGSLs5juBj0oE0JS60577TgnxxptG
m2GW1wXmm2+C/h35HkEHB+Bbe22xAOtd8Am6yGyCfezPA1JI6gju2dxhnv4F
yy/9Y330cbnTANOmDsTxeDpG5+V7dUiWMUCdhFMxVsIxVUiJlJq4Fyo8SeyK
B0aIRdiZbLLG80Nc00VhVrVMs87h6QSd/Ab8/8QkjWM0stoQPI394KUhS5sm
9UM8htMme57dG/TfwNrxkPSpKP3/LIpajDLNmGuy14ap7epCLSxJ2Li3NghV
QQZgZ5pHXRSj8436vMeC1c/H9giFUkoZ6WJzAcq1AV9ZHLfJYxo8IzzM7pYS
e1RmkgqwcbsoSh+4e9EYl+yksVk9UjX3t+DJuqdKpB3TCUJCWJJw9M/pGb/5
VA4A/b/cJ6OlbMfYvqDSvN4OLM/TzbKwMZ+wuf94kzP+Vpz9XG9GNkYG4W6P
j4utxodifOWdmDZerRg1mpbmJME8/cYg+eyjhC2HxJozPU5HAshMggEPe0Cs
YKp2AnV2cuIe4jksqJM+H05XpfYxxFYVSyi38YCpfBkLe7CEGm9Kx2PpMlxC
aSNnx5fLLNj2ILRQGZB3Ey+2gztD7YRaY3/WAUauQ+cD3hPCl30FBzAALbhS
3HV0YCezxaspiTA6Q1nK3q7aBBIgA4ixQ8DXlg/0XiCaOL7rNxGGuVov26br
K3+v/trRhS2Np7LsYfQumWmnY4JDIkCXDBEusrdNdgWYYUWanflZej7G0oTL
8oQzyvRCA67rNSLpIgJA1WKSTls11ux/Zb+0ZemFhCmXC33FYR+9eoLOuZfB
B0suYNgRbKHqPvkDYGUo+zVOj5c7pm4FyRhKgZDvcouT2n8ODLrq+CO0cDZq
ld7R3m/9+//zatEVvayA615WbdR97843VA/VxOjDUk+j8wER1O4hkhiI6u1W
YVbW3VtCanuPlZrl/G/AejOtE3VHxogMa8aWqyDYyznPVqnzv641+OdAMhK1
Gh73NvI8r8Db5HJo3hp1KbheWTkO3cK7s2UcKRECMSRpJfbVykIOkHZt3Xts
aXw5+Dk25iKZ5HdqK4gD/snqUY6LVhnjXir3EZ9fSKTN7SyJqcsCPPR16rvt
mkL3xwFmRVoShmdeRpvmQoYBhIBCk3goMcGVHK0hg4DseTriE6MoBZ7mWgmh
XfMADpGGH71hp5xJ5yHmGytBA6DCYQ57J0uAXpo3CAaEV8r2uxvxqM6XLsC5
nMpeWQDqDEHeQc3vHbkChqLBRsMdjetxnk1215D//fITlmwz8s6nE5V4xmh4
mbSDZkbzbx9qIfFd1Ardkng499GMQzLpUYbjO70Y51Ndz6gal4RlzkFeECdF
N7HIdYqjP/P/XmOWwzbBvYXceDs3Tfws6OoQGGSdqAl74bM9BiGKBRD2odE6
wdLJ+3q00DNfZj7wqtSs99Qpgr9DYT7PhsurILeCBtFivoAldyuqlOWC6b29
8Jbll04Ywu2J6LP1OAbuOB3yh21VLG4HgxAleS6lnnmc6c0z7ZaAYyCR+74D
ci/GcCXgPP2L4gvGH9WTDsKQjASToERc1kNbG2ehNGKJM4i/kFEbst8FjnP3
BHKz44RaDJFLqd4hzu2oaTi14Ez/ahg9mXSLyqymb3dlWxLjYQ8hBAmFexNd
5rYVtKHJ+zRtH5rRguz6H7/2NSHwl08cj5Kqbv5gF51HlraRsFz6GN77rYZy
HZ6eL8D4Lplx5EOc9tgzQfHAgZzxRBrcc2N8hThLcykVMNn21vQXemSIsTSJ
557uYvB78EmBYUKRTsWcT1QytGMBXjvhHoZHXfHcZmlePi0paPoAGNLum/Dh
XG8Ig00NnNCpb0drZm++IhFg57emWSvqQmxSSZLCA+jGoOhw7sxA8gYY2qhR
8P7rSoP+hElnbb+mQgekVfx/RV2cT951sIGiqQ6oD0/qGAcV7c/eeJ/+QmOM
M81QrM1jLyALIOOwu+FOZKIlCDASfqyWtsOFxptaOx+eOnwMCzsEAXYqrDFJ
cilXDgNqMUr0LSEB67bMcEs9ftxr8qA+vPLvv7O8DvzuLdqOJpsjQjEbbA9R
r8xb/xPjZyx0/SDxUmSa5BqSB20RhqVHA0RBniIS8IQqdFMa6zx/+NIE8Txy
0VS8fdHoa82QSgxGWksdWfcxbklVenUMt3ikNOMYJWm2jc3ctN0uMsR8RFLK
Dfz7u8N9mzMxUNJntM8+fNcgiC55DQrM4N94OduUUjJzlOnF40S+sT0eTB+A
SIqzTVa+aPRbcxyBLTU0cjGcGHDlLu6hTTnYMUmHXXB7t0y7OeQpVaqpmYMj
zl3rtCvou+qROLvY7B/Tx7NIv9afqAJPV2UCsMWJe+taoJLOqMoTc5v0s6wl
QUfn/KdTg8q7oRXQfqvOMpuw8zE/e00o4C3iK/xMIny8RsdUNXbHlJ6oSwaS
CkfCCzGLEf6nuXAAc8SFyo7NoHqjyWUftt01+ySuA3/nAopou0xg5rQ7vYj+
25qU2Fem4Q7NvGEfecu4m4+ua7DgfQrQRudZolwd03Brx07xahyXMJTawGBT
tPczDv9ytZ11OuF0RFEMsCe8fdMa4DPc250SfvFtr6YCxdFftZ2CpZgdNOVE
gryuFs+j+9s4BzE05AoKEZfrDUymbPKZxEiX/UGnGlI9/vjB92pkI5uKtmbz
IUPTVLu0Hus2biwZqVuB36tTNpMnXZuiyLmCFzj8ABwwC8KjiSGSx+TD7jgD
OYlIFFF77Z4Gil8ctt1ckkkeCiw7VrQJqtFFAdQb2xCEz0vrmouaOq8+xc2j
GkUnKsPXuE5kdjI1UVTFUdyyFuVj7rjQYbRVC4CP+XLt6CVVJPZJZQMK9Pcv
hYV4xQ2zHmfJraTq34q+hEimgvMzjQgY6VemOWXymGzxsnFJE4qA4sau01TB
H8aNi3qTKPM+DBF2UMcw0ZWqKoifv4etPOGQYUFQjtRwI6dTCMh19LMC2iiX
LZfB9jJ1NZpjARXUUMjQpeL4YAIUma85aLxh+Zg/n3RFUGa0+Cexrm3f6uDn
6kExnsR9xELzT2IOGY6MJeLLB4Yc1Eu34CEJvqiIlUujl8GFxbWat5dPWs05
gjNtE6cQlyDByYH2ovTeiUjLg7tPwvYGo2czNq8aQQHQ7tWnlAsC3fR/6VCq
v2pDuLvR0nn65+18D7V0gbNDMHjUbK92NWUGP6cPgTTi5EA8CXRpcGdrmqIC
l8qaneiwkvn4QjXYc5kRcHqqldu1I7s6BdBIFgADN6lpj0QFmju4wPp5Hro+
ORskCF2zuU2FlU6clRVULznBQyW0aG59NfocK6XQ/8HJXRZeY8BgFWDu3As7
bw3zXvP3YQpap9xN8sbJnlFxFJ9nLwIEgjsgVI4P8xY2QoBpWydlxmp8dl1x
okPLupfqYTuMzDVlVvOm6/iQiwmixahAl6+a9ua/pZKEjd3Cr1O95GTI5xYT
ItXbYGa72FIve6anFoukDdBL3XZJc0E1QfiaaFrFgoR3EVSTuYnVGpcgh1GC
TCskKDbz2Qt3S4J9q8Yya/k3WJt9E6juFp4ijSPxn6efQ021CpXHdOgpC9Qi
Cmfi/V+il6evVFLZGIdyMntXufBAGZiFm1RyKGjEyX4RKgR37QvLPfShXDOP
hnzkEV5np1EPucv0s9RjmoITSHdrAeUp4Tv+c5vxlVgB3Y8sIA8HCuPx/Cgh
Z2zuYSZQQjkcQg5CwxzHZQgIIstUqyEWiCnpJ6X2ulHGx5FxjsKHGWMnHLO5
j+cajCmaTaFEdXx7VcWGQzNhflxPyA1VdzCjL4vA/NiKroMJtAdyiTpUO+iu
KI+qzljJsnu3joQ8SuqElrEJgYmKMp7em5x2sy6eCt4GARY+4Lb6VXmhoFVO
su6MJwaXPxcUVjUmVEKJpcTWhNHsnGxdVEdU/641r24W+CpfstvobBQ0Jwjh
7DA6vq3WaPIrPnYrLPNBGlrz6BIfSMgZn2a5vv1H9RvsV5kRXmpcftvJWOS/
Nc/DMuHldXVSJO8P11za2TS8JOCkbhMPHT4JlEAnvDjn1/AaG5z6GmB9vQmh
XsfAoAtOgBMBPxLeNEA+z6sSHmbnq6fBVWhbzfesCQhWndDFFt1sETBRlImG
PgEyO27UKFXtioDdCy1qSL9Jr1BiEt0jVyDDV2USz5+jxgHdylATS+jSQI+U
K9aHSPG7Okyi4vthkkiYlvUCJknwRRbKXYPl1o2XMr9go5tv4mLrTv9QIkNW
sragvoSOcjNu7DkNRd09+NJjbp5aglTLG6NRKmkWUdTs4ap/pFZMK3aRWNl7
XfHTr7fkiEpurRhoI451DCG8DJCgwjzy//fPbEjxwMnBVelDBQikeZbrlg5m
VVPIePtNytXZ9xRune+iVZxMmbWhT/d3dCnv60dPFh/uvYtkmpSPAaWOkwa5
WU2P66bjA3JUDcbc3FYeLDGqspAiObQJOzg9MgDyiU3UVEt9Mjl9yvBeYu5n
UDCVr1x3uI3b2R5vZz/lmuTn02au/L+fe7vbg6bbttvUvG+mgBpA4zwY2ir0
Ith7b1BoMR11ZO8enrxaVyDpHHIwdQ9ETZNI0n7q3RUFObI63sebgT0vcbXR
ZS4+8O3Sj+VnSif4kz+H6/S6mzUDRIxWcFXWL/jT3GGZ0Xx+vrbTDmaA+JLU
bvDlh8Oyqfao5TV5MFDW4PSIJ1IU4BHRk6LD/tcZrXypHjn6Vdw4FLb+7ub+
CEHlKXVHUxEcsIt87cHkB65yfVkH4xRc979Bsr5WNMsvcb831cID+CByS0pK
zmENXbSzRxycZE2j+uK3e+Nd3Ep6kHIpacJj1kiC1/RnU7kP+qcfTuZjcSR2
FtjRIdCFBhGpG8V3jtR8RjT5RAZYmKKDlACafRzG3Ddrn/ZcABlT3aT/aFWV
Enrnvpvi0+Pbj7uz8eDmMAD95xH7/pT6fm/ARx8HKlgA0cClZQg/tS/OZBcm
Xn3N+CioMoNNJsUKRRDBnzBdRqYE27sKL29x23/ETBp1wE0s4qCcjIOmAVSZ
CgIQwL4X9GcHK8QHIYtwxrkoL9JBM6x3HhL8a7R58VsSfmaJu1O5VhmiiAD3
IlY4fcmlD/V02lk1ShgsYokvjwuSAaNYu4DaTm0P4i/IIw+brEwx+wXXaIZF
Oru4xm7iHvuf9a/aKgAvAMa3502pOrAy8DkCGULCmLypXN9J2fc84NNDVNYf
Xjsq0PubjwX2cJbtWEkmzSEkU9TMNhtjv1zb0+xNaiMlNYsrh8i9bQq+cKka
D/eRfI3oYZ6f2CJ5rkrEnPoxZwgS2XFWhw2mu1uXN0j573OCmfYYoVYNqozl
Gi1ZlvKHqeGI9VPGvpnPDWcfMMJyVx7Gwm8EDl3xpwlUJjg8yUbAlbojcSve
FZ4K58nQ3UGPa+5RzKyd1H/XWLeHqHUH5EM0pr+AnNdl9wbTsNmW8VBQjclE
ZM9Ott6BxjwZuWBN/Y5OWaHgUkphQMtj8pHg+XxG/cLTMiLKqnPUno97eqfK
nXmEAL9k3xIygv5tdegdf6YIMZpfEA0vayi4Yny3waqCHf5wASno4Zv4GORM
QK6kXOyzgpnBx3YhthuTewTDyw1r2oCGmQCvUrrM6e2yd1KfQx7a/a7Dv720
jI8r3iWamNZgnSFZaX2OGd6O7JCCxiqJ9ml3wD7sPx0BidASAIMt3HojyYgo
ULcYcbPNllpNccRhQtZgJ+qodOUR+XR3e1SL17su/NYvY1yMTowL2B5xwiTa
C0ic+BYZx58WDU2F6HAmmd8fToPrwj/OloTJumt5xpjATUXcbrimunFMnXlw
fYv/NSxgPTy33xrLs5SRBbIdsxwWfN3cqMo8aNV857jz97Ni1Cj/PL+84Ibx
AX6aqCZpLv+sNskwJFt1sACH+rmsRq2CfmYEaEsTTkrGaUbHOQQWnShyqRca
M5rkH7X+Z9Dmf3VdrVLzIe4sVONVzo/wcwrRjWc5yXPicmCcQIbP2bT+NTq/
deq0z+WLA3N03/gPmz39XpsoZqCpZr4SwVRZMr0nrZoVFwwEOUz8x+UlIYLD
aEfKsHl4bx1OzS3P9rlLpbvEe75VfEd3LEDhfyRmKlKNQodvZWMqhG6pM+A1
wABZOZPy+l9KRmcO3eFYyuJAKluJjOOqfO2JskJWrmSnKoXRNy1mz4eYjdeG
GTJEzFVEnbQ37dE9Ow6UjtBDMKk/YfFo4u56AUqayPQBF6hAHFE7ec7G6JcF
C3fvFv4X8yZ6sas+EoC/O75irBrqza+C1E3373/ZszmrCZHJelwsBUS9N4Bx
yjp6EBO43iPtaci02mpMC0Vc8nwJy2TObCgJAxKNnsZPGLD9gkkoORWyeCbO
UbCr1vU7x99pLb7F/3cPCGFklXC9ddcPNXenCdLOtcsutvWhl1Etf9mCGjqc
TUwouS5coBBkYGKf5nLLA9OtXJapNgjn8lIx1inxSaUIBawAgTcy5mIE+1tz
0/8igjecNMjdWGUJCRgQpET3IyRZImeusc1v9p1phYk98jadNUZLKp9U+5hX
QtaNe43wNwzbTLEMAg38QLX4SZwaV+w601vF5eP7I1Ds6FGHx/FrdCB9xEbj
EN1SfGYrOgi5a962dqqQ95CvWrrJmuz6NYZwJQoc6Cgk6ET/cahXTNUa59Hw
joOpZQK0iAD8cyK4pzjRZhKXiZHbdGy0UDm2iXCr+Emc+ZZ6UQSvcvigHJYE
+DPskDrTcMptK1/23usogAs4pTEoWg6TYx2U6W4kTKoCfIT1rh8VMBQA4EXg
Qp1h0pgac0qMnTSeMYXVt+6iaK5L/cNb0j82nvO7wPnrU8AMcI+7esRpp6wT
CD530dRc8yMQFtnsFRUD4og2BRyFY7D21cARLFUjNO0idpqj9ixzb8NRWsxM
pJVXQ6/OPcGyA6P24lLItzGbDVxqyuVmrlaj6wnVkJ5Q+RL9N+tomPKnm85S
JDvOKNfOPF4L8Mgx+nVXb3W4+r5vbWK3hQK+cgz5nyjFLincyNCQLGdEfJJQ
vn2/g3QbLYldxoQjKpKw0nytkzTD1X37lecuWkEQgh2PjK3ItHiEUdZe3YFl
umr1jXwfo1RvWTfos0lkaVdRdYzhLgWakG9ZaiC3l9E7JRJL2b2VmyridzdI
7oD5NBNXlKo9VyU3XO+fDvS/GsJs9Vy5yhLMM6V+zmsuZIl+bv6WxGif9N/j
ERSxClcG9G1EonJV/rOm/WBu9JC4okX7usd8SpSmbi7FR7suZaqcOQRY2Fpg
7uQtILYbsjxhCUROgLkra6ThcAPYBux0gojpnbhW+JSklnLx9KvLdIV9EZzY
2dswigK77r3PxOb2IJ0v4zzkOlG94tQ7fZJQI53z5CkvPw/vKruYlkK/BCmv
NRgdzGTC4dhQsfpEaoU7oFDMfw+MZv1dfKu2lmElMwO9YbESfs6O0Za0dr2b
S0r5YP1AGTUi/LCV6y17Q9r8OS0cyJV2f1B5jzC8kyW745S3k+w10WmiiUFu
9TS3SKSoG8K48gXBvw9mkEbzHe13sF3DPIcC8X7PvPyPX5eLIk3aMGGvuowT
JopQliCSNPaCudtILnHARd75EWX/e04ZZQwo4gCT2DPEMnLIqtc+hYVEZP4Y
CrGnHtnyY0bAl73Cc2A4Mr//c36snn63JMO7M8NgzMY+1CeHujxQCbBXOAXp
uSI/heABmVCNeTNEkHFIsebh9OQJraMirWFmCMBeYI1Oxo2JdK9hGqPwIomS
ZawYf8detlN9oj5biAuaV8Xbo4CZ6gz1CKNnQHkT/5QMfu8QBmRKcc4ctp6R
j3agl2/YTw9ZIGOY3T8McM+7t2m5jJ4bQTWZEkceeMzHI+wjDe14uW3+eYA1
upaxU2bIW/8PngzSOtb15B26L6SMb4Vj5BxlaXWq5Qd53qW5e6tY4qKpKGCh
jIwh+c8tF5wuC7PEvNk+HXTBG9qpbi023ocDQkq3FRkj9Z5T7E8DsW1fAihZ
2VLZHa5mKAZ6OtSYdIrxV3wcQwM1+OBEOBeP1JPn1wGOWbgrsBJ5NfQebvC9
AqUrOdCfh0Dr+e3bfKGJmrdvbw5y98oszOvNUMfNhTZQkkVJVFpZR61xng31
sSlXMJg0+fOdIvBhzaqXcfO3Sm+fDjwfsFuXKWlHYkd8TfTX3etORNMBiN3u
zqwcFsCr9Gu/qB+g1hPqLvrCE+NEfd7TvM5yNFSLuOySSXhsDM7oef6pP2yv
gVF1+nBrfVv6g2Etul1hMSvWvx1reW3DHqc++EzC5XSHkkBzoGZepBLflqGp
ZSTqFckTquPLnupA9fUUV9Iw3tyc5MV2DhDCpaTLaFY5m95xTVl+MiYcng7S
+NrguxV5Yt7ck9KuQR1wk7HLqwXdqOiDa/eLeyZfi+O+FN5YXmJ+Po330z9B
qxBX6OV29PmETxBp9wEYc7/zmbKl7hGnBIwiY1YFuE841627FOOqUJKTm6t+
lw3WRmk1QsPuD8i/MQChjwdnQ5hZf8ZLK8iv1/xgaxcwACD6YCAOyNpDfSoV
5Mdawd1fU7sk8zateXDIX5k0Mn7BzVJ5FXv94/xBO4jKn0YYmXIL7IIGfTWj
PX1u9rQEOKhXByPJcBW6zGeIKmr88buzNTXSy/HHDZ0ehwtwCK669ZfvXb59
EY9h4sN0TZrMf4FFa3XZFRB1Ww2uTa54HDnMlNjCanCtRxIqmuOdqCKWLzIw
73CQpxZqqHdFSB69IuQWm1JPP6FvwpaZmxYkaXipA4ZV4sZB45t6u8X/s5Ze
W6IKRDbTsH8GyExi0yIdTUOlUVwbFuyH09nyY5jL2mrj5Rbd0qt2jM5/zp9o
qp/vt8zmQGQj8vd8pzr8gBEGr7H+ofIjHqwWkYnkOVnPRuOmMK7S+90DoBVs
qR6EdH/jrjFvciPAJ95rneXmhaxERjsKeyFIGwo/bF3iX8TcCWloY9+vDwNh
UAq4SvzH5c+CMwBVbE3uMtk9+VH3nn3v5Ceb+Z0G+JmUehIDU2zDG10Lp9cT
BSO+yMnWU0c2fowAA/L6kL1eYzrqbnkf9vX1/B7yBMy6+/5MjILwjDlunvcQ
WOCuPs5Uli/h1MjM3oKIaLPC+g4Fczk496+rwlhCqhdjkD10YRtiIR2yusE0
D1CdDWlKpSNk/DZN+CB/Ww9vASJBUNKfrr645xFEIU6Fmsl2T07Aji2H1NK4
Ll9cizcULzt20yOrOwASPQx7o8PPsZbl5YmZe4Pihv6Smhsv6WkYT2eiqUma
LQoNisV/KDhogJItSK+hyELEJ4JQLFFZpi/K3n8wVxmaZaGlom6OxblgeFYm
zE+qMm2WgZwaDm82wtwDbTJutWvtZdDyrZuMCSCmSoJ1pvXcb+X1yOvIJvC0
hKGXc3SDL5PrAsl2C3Sa53lKjByQ/eNFOusDIq5TMKyoLbnjhOon/5vE3cgg
BnXnRxuawoSRVCgALQs71YLteHcrkVUJKF1nzLGQuoeKpBE2koNx/WdVGqF+
ieIrOo8SkVK7198kisTcICKBUaHxTlnt9LJgEWsvYcyySuwplF/J0GnRvv5Q
1Os2B2K+YVJlC0hIt+C1WVQgYx+PwC7XTdGCkzuj94sOAMCpiC4s78UgXfFN
o8EQTkgKEUYhHlWwwatiI2lMCm7g4yydIcDB+Xm0C6lHjVvp5EKisoYKDZ5b
JbWqal9KM2MJ3z+YnF7avsv6f0WFQjJrrlm12DY9GsRnVznlIDGw0//CAaUb
3cCsHB7eTnn81Y+uMjVY/VXMEm4nuC2/edWUpxf09sB6JufMW6jRB/x6uIoU
NN5zEgnp8UuGVW8sci/a2GdzJ1m7onWbfnO0XqQ0+nf/XOXGSVWWY/cbZAHy
Lm4GLII93XIwjHTjnk2dHYKYtrYWf+t8fqeY6igMFmA88NxfsUqfpYh9xdkU
1+kaWsDTEwFrZRQ9HtEK7txq+KWJueGkQYEcE2h0jRdNcHas5jfmY0A4dJN4
iinJyBwlvRFosoeWV9ipNjp2I8uYlyOAk30VfQeeAyib1LzVppqyHInpdzG6
I1j1g/paXhwV9Tg1gBVj3Abf8P6rN9fKzLyhJt2kqv6LdErhHz0HZwQAGFM7
tf0wKtrN1gSG2mqqPe1AE787/56dnqZ8lxwZy15yNs8fCkxbOlwHGxrrUpSi
ZOIc97u0hA0NonymsCvQX0pYaCYBrzamL+NczV80aECAr8Z1Dpt88B5mWOI5
6DQC6tTSP0BVqcW/xB2vUTwnDF6r4CRGRnZby5e199w0hTwukeVSAPd+0qTe
j7Iue/06RHxg0m5JHs8udDS+090KF96JN5yHmBwvflun/KLSFrXaa415XkhO
zS6xMpCfJsEyuH+pPZFEphwE1G5yNnyX93DBL0sMqWolKQzG4l9inPE0n0TZ
teuC4UhIEn/W904dsU9OojzAv56G+Cs+9yvyChuf4OevP7iLLH5302otxaJ1
4tsSUZG+Y68q0jZ7p0Y/GgAjIrGLPrg0R/LShFjRJLnq8XQmNSjl3fODyuDC
RcjAP9aissjobzUInlTo1iruWfCQeQbSVHyEUcKMUcV/Bhef9L2r44B515Tv
TN2IecVvBvV6zAmZMIPHLwyR78nl8QbN48kWj1AFtWFuQzKgYgKOgr/kyYDV
eMvQXC4wVxwoxAllRls/eGhy+hGmUdzX+N7bEUGKpGCAb6Zyd63PboB20EPE
0nLNv/0Vp/fR8Udc2C93sw0UWBBBrv4oI7bwcSB9+Fz9rhQ5D4AYEMvy8Aaq
XC0HsQPWGtXYDqvZQZO2lKz5fCoTyYzx1YP/ex6eyIpU51X5j/YSmWpGTINS
4quZiW3UpFVMSQyb7Wax+W3TGmBclQ1ePb3Rt9Y51dBkXuaNJxFuvMXDrC3A
dPrUQ0UCKh8GohvspXsUOxkhU7fy8nYv5GPSGRsseYeDDqAjV+bDU+UmkjYw
azmGy7GnGoMovLst6KDsxJ0t/bgRvEt85+NRZ4XVzlQLO6gWCSLzHbvw6qqK
jV9udlhpPWcHIe4o3YpedVVhtBdWMwIMaepfZkRoabqGEpcANQhqf81Y4tF3
OLiYDhglHDgZKqUvMdH/YWFc3HJWpGSxYS6m7VW3ENQTpaNn4cEZZGGfwPVN
tPgEfjgxCXhGbsQXSbf6aq8g/+XfJJXT0eTRKEedWK5NeB2a0b5/zhzMjYRw
8dAO/ph177hP9EN2FIPKxDMI/u0XGHmedLF3wmrj5uqwZS2IKZJMGdn1aXQe
rdCKWM0ZH4tij3gLNlDf20doG4/NilkPZWbHyM0nvu+3blAmDMxVJCHrfDRI
YGrBZcqbcQCjJRn7EltuphKVrPnztcwwVKgSjXIRZlyQwTW7fkyZNp8Vs0dh
B4biAjevfY/FVvjWXUrKnUsP/hOqJwHkxm/eY6BzNUEyO5sIlgCY+GPg/xOB
dsXP6XfDED1Wtvu9SkGNlLUmkr5Ghys2+AFm64+HoD+ktJcKPK+el3XKS38y
wIS3jZJbHiE91gmaFuw0pPIg0JyzJXsj4jmycPauqIsym5KUsxGIc74EoHRl
XQFovh88r/yRLfJ+M6y5jzdso7jrijtV+k0Dpyf0X/NnrkuCWHiG/39zguGb
dtYJwem/21wcXpj+skYAe8ZpscPvoIpNoE+aLkWfqiEuBInuuoMptGqTTCr7
EJO7TB5ZWZkulDgHHUUjfjjn3RCPmMOSfsF91d0ItTsEHCkNcQ8roxsjX4AL
k74HpaW16d7ddcZ1VHnUvyUglKmwIOXA8B5DauiS10c0+buY2qJhMofrCp65
ioUSUTkvpBFRX5XyTAlw2Dw7bDlT48X6eQ3o9H1KvyFiZXOzDN5M5F2BH0JB
dC+dJZ5iDxyCS/WO/sgvZDkpbZ9Vd5DDIB3eM1lP+K4tPaA2vieP/HiFFxrh
Isd0ntPFEpHLiQUryk5B/nG7H2EmpahULTwpxBZej/B9mlYuskQ2WoNomp7s
lPWtKEjHaeOtOpzeA/VLRJipJxLfnPO7V7W2w9+4vt93cZDPk/wmVd3YAqjN
gIulAkJmQovaN9yB+1EWFbBL0o63Ba1jOoWCJwlalbTlBjLm89wXZ5cMdt2Y
ux6wWAOCdkIsltHBbminRP031B/yCBjaTC3RDlYmyxEg6xIxjox+PNXOtbcd
dnxa7tOwOWfmSTLuJTQQ3VvttAHqU6QoGcgPFBxLRBt7kdKO5JnmTeo6B1n5
yG6r7MG+VzsFKqPlrKJd9Hp0bwXsj1nqRfs0tiliD7+BC8YdSSqO1XSGPCDJ
uIc1/HUYp2dpeTg5FShtWrik4S92Np8wl2Kl0k8zzCXD6Iow4ke/Zq7eOu/A
aObO7H1gen0kqaEz+Vrd4PK1Up0A1xGHdHTuMQaBl4yOtI4RS2IQXdClV3QO
UGdXMqMBTEaWPj53y7lg7XfKBYUHP2oG4S4uN/yili0hZ7Q7fR5AvJuZlFQO
YAedmfrbvoeu87oJgva9Vnsx/XCjLLBaxLYDt8dl2HPSLQcuH3wW9wYKWzEF
dPgBFSK56Zu5fI5v2Iw9PgY9Dv9oT71LIIbBpThw+SiV3xW252/pX+KM8VRJ
69lPc0oOezmjdwM78lRBwTv0YcpSm4Yv//rCzc50VNsIi5poULEm4d0Ux56b
J7I7HVcpC965LrxH6JGDcxQp3OvluKNKtn3ckDqWVN/k7IM0/k9iEVdY56TP
zxz+LygaAQghepGU5kS/n4n7rpVgOrKaJoVxbksGkfDFyWFrL9+dYAttfs5v
ZnJZflBxWgT3wPmiURSfPjxPkRX8kNkEdngr6mmDoeXUVLb3ZoOG99R0Dq6C
Ynv1r1iijPoTMwRZl/LQ0tAdrBsurejsDC063fXfot1bWHhs5JOhh13eZpwd
GT6z+s+t2ciWOkp6wk7QUpLMQMVyy20MhpO94fgcvCPEzahSmuoaYkf0BpcW
L9Nt8q8F1h9DfDcRvnASgHCIVJvE1zSbdP7lPDmaz0bFMuH5JBRyzs9KAKGD
2Ced3uajfVhPjgQ5OMv9Tg7vmske1wpeB3MUlaP8wf1I9il5MgniVtKWuWSu
jH5YGpEhsaUycxwmCuJ3IBeHHhZ7RlwJvKfw8D04ZNLrsEo1D2p9bUDQ7eNG
qA023xcHV+uA1gorvzdnPZSYz7jy8BFSThLhcX+1Il3OxDqPgyUsymqp7cQm
TkuAQjVCNeKz9dA8T96HF1Ew0qjChdTN6Y/vZBnXd9wZRgN8MQxi0QBCi6ZQ
p8mpVk2obKj8NMYkDEBue+lxrdvtUJVanR1Bo4SNZfaQpjJSsvA47RO1QQ1a
p2tV+aDsdNcNH5brS1B/4HfFy9Q+tp1l4/nQXEOXwhWsrUcArq9GCFRdIrsk
qkZrJkmCrCFtZ0cpl+ksR/j/QFhPNrVszprqCjKuFek3/illq3PzfD5ytdv2
yEarPlJbNJ6R21CDbLD8avd7ixyLb5VGYrcV/QGLLxEd2BjSR80SBOxJTOW3
jA4n09sJZaQVMLI+bhIRzfNOCRxxJJ8zNh8h02nAkaCUU96OuWiVPakell0f
zIrwN/Aq2eCz81D+ptamwUQuEEGXTQt5xNSekAvfmHHob0PqlWonKDkCEyJm
3Z17kTNZQ43FEPQHAdDEsatoz/YIDeOfS0ugJWWt+KSl/lqCenn4FWFDp6Cg
dmzXSi//Nn/d7dsQzC13RVye5rZslPuAwEHCIqXvm/HCuhAe7Dt958IQwkff
XKMR7WtVJDxSL0smXHrnZUG2/HDVG8jRem93tgJWbCJocog3NGPiKCzaQKpn
DrD9A9FMiYbz1FyFm/6eZ2H/ZB/DczLgPyJSSnkKloReSsJblIdfHbVN9aYR
uqxfIyA8B7lQwFJ/VzLvoZBTo3l784J42f9bM60KUP6LyJQMGsiPjei5JMeN
mbE4YKAJ6SNOQOM5FV4xnq8g9BkGFvo8vGGWTcGoPoXzgvNR6fzvHQLMarbu
ExBghjVy48L6jp2zoE/j9QyMQa3CA8dXsstQ38R5IZ9gsqd7Bz6M1gm9V4Fp
73gzLpPeCYrV2lBu13p5hemp6WPVNsA7yuS9w9XpUWPRuFMKvoaxZ6xXOYI5
p5OdFj+oQqQG+WCt1m/lOnBuIX/AyJYbZ/KBxbynaBgZf4uUkjjOFpWj1bi5
0xd1tqebMJ5gt3+iN09iuFS0g2JL1pk4MrZvZt6jzDl3f7FUGVDE9+3htbXz
5migfpeUffwyvt5CJBQIh4o/hX1ps7htWWg+IlXI0wmN1tLWsm40HZjzrpX/
LBxRrdgpj8+ACtjgaNuXUGBwusS+SIfo1tg35cAgDX5wwMfdYI59exF4azFi
8MDCZ4X2NXh0DMeyRMe8wYrh1ASgd3nXFvOcYT2L8URIujtFur4ECJDY9hha
5xBx8Woq5WBDenCZYfxD9Ozso1DjqPpH7vL2BjWW7iQ9XvZQtFO0l5jWswc6
YQM9qJxLAjsOpxB8oEwbZDVRle6iquSl3WpLWhmm1Fw5NZYIs3iR0AFtWvWj
mgtAjB8kCzvgSb4Mi1fxxNdTJ8n3zHipnyci37nCPKWoc5hVIh1flh12hZA5
4f3mVDUGDaiCBAhQTYDLSkXhF2doMy3bKUtf1rmufi/ZNDVRVhcP/xg8D58+
D3vDFPZLmaqGRVhz6VNGqMsFYoUfUpN0cIxIwa44kGZpcEYQm6S+kiSH6QpY
d4vOi7atAMXO5LZkWDhitp9VEbZsUDl5tSDACFtKP5MCyM9OfuIXEpaY0i9e
PRVRFdN3GqgZFIX7bx/aJtKRzm8ZwSQQ0y8AVvse2wLsJv/c+gfuQzvJF+uu
lkNmJIusb2RDYmVhNCFuvB2dbz2tkiU0mp/SLGDDXvZzXOqOy9PqueAxDGAY
gicOdjguRl08L2zVVVfqLbo9rziaaIU6bJIIhsTBgMye8p4yCwZB7mc3MUN3
v6AMDyogUECOmVE+0N/yKfT3lp5+SW0VvSA+XtupEK7lzG99ogz+jAPr/jU8
5cI9RV7bR5NtwCJ3rAMdKWmCRS52IbMNi9sacUXTFrNi8AQKU5ZJtzi8qzsp
But9epehfvtzGurxFGsWEZsbEZFunpMbsO3y1WuuVUAnet2f6YH2x23FL9yp
7qYtWkWGpXqjYOp16+MVDJB06RJTA7SnQPqLAMi0t+OurcQuI+U56f1pdfn0
6+DbPsGB3bO8GTIzWztAmOUofPz9uXjDYuo24PjbLYXxPJe/3cYcA7CStdij
+H7Fab4PvdFUp7TyXXo5T/seQknITq8WlKk1NsSNCKO8ac3gQtQ8ANfzPpCS
RAr2Ath3slGFTJkJvK3xG6uJmZBmVo+GyWQeVFy2mkP0s6hnTWukdo3MuhRP
g2Hn4NC1fPrbNSNb6HVpUARwR0sIB3HyqET6QnknfDlHNBnAi8S5BnVL8zoJ
RYlOGvc7Us620Mt6bk/26rcBaRsanc/NrXidWzB8E7hf3QYNm3Tmti3fjfh2
4Y7JoweTVRvNBVIR942PPaCsYIsBMhzeLaFxhc7tlLKlAKRATVgPhv+fhrid
RCI46f7B/M5TpQl8PChXE0FhAEUHNdVXt9gqY06VxeuJMQ5Ads/g2Mxkp3d+
7ZVcePYco+FiJ1mKJbR93B+eRV0kwbw/M0jYWz7JzUqJC8EyaUopeNKLgWTt
IqjFnlhlB2DerZqCyW4GuZm1Hvo014jAAOmwK3E47jxw76OSZ+Dh3A8NBqG7
9KSQa/AS0V8uTpYLMsvVCpyXAPjrXm3n7zMqiyVK580ykJ8D7H3IZipG41kL
mm2yl8Y72hec4I40ErkwBLAHhm71fZC2zz7AbJebcZR959LUlaGvKTxJ3PKn
BQ78SjGQjuKLXayxzItBOgsEcN5d+TstzsJmINtC81NYjaYoq0kupG8ylH5V
lklqdsNIStJlWU2ennYdEsPWdiDP+cupjdlBTErmno6rqjLFnta1TO8tvyeZ
cBoOSByv0mH7H2qIblJ/+E2wgbJFzTBEilZoQIgKTDB+skzTKo3nqAsZ9vza
1li2tZRcPT81hFXCAYEXxcbVGzySccBq4ktQp6uNAze62uVqjQy5bzEnIVe+
huRKZbRH0OOLT56L7ntcnxWGRT06L1vrV7MdPkgAjEVCSiOacpwzJdtAAnpX
WXDkYxNgfBgN8Pl0D3hdvtipxN7lJkDy22HtMLREim2lemUmt5Fjg/XGH2SP
q+gMycd4FZelLABmH/XYLT2jcUmyq++YMlKfhvBd/OFsUTamOWkXDuQYntHF
EZtKGUIGbr9vLzaBJxQM65ug6XsXvMfvxCx6qxX0E1RVGHItVROItkmbEzyU
rgBg5cSWyyRIy/p9+aVEuX1mBdVnV0a2ES7moR2uqgPn73ha4nqaTGsatlJZ
F/EAa6Asi0BSuCFEzvLhp9sBWYxJ6jfFZdsTxY9hcsxt0mKd4wjvItQ9qE6+
WwesN7ewK22wSRKKzFFhmbC7agGB8ZaZL0zutWaNiC6sUvqOvxzAdCRIQrbX
xRFy/RBdq8E7t6SYpOy9mTAOY9Kt5BsBA+6qvACtQ11p77TUjeLintl4qZXi
Qtp84u2GrvtEyDLWVtoaCmtbIrlMTzTkDwG6vcCgphuK587G0M8O7MBq6x/l
9l27JC6rOMa0ARkr5uOYM6Q8Xuw4oUEdfiy5qYX5MN7WyEPnLfsNwfWoTp60
jIl+i+t1YCtNYyIj7IL1dKyuENWN3bt4vfrWclq+QhBGxRCZcHmRBL2ircf9
ISY/Furt0CN4mz9mV1ZmeQkie2r3ym65bUv/GO5gyYOD87iboS+rAop6zAXO
L/xBOaTjUrfnA361sRpuISZ/X4Px0ttiIKEYvqvq2VHEF1jUHbNvQGGlVYHz
12EVJ/Pr5/n93v2LkmziPLSRsvQQaNcss/sjGnS5nWf1qCXFvuqhRCSTe0j2
1BvoUCyib7zb2YyHn4qs5ceiZFcpXBvSk/Vqu6gaLOZ2ic+QemheakD9ZEhx
Gtc7LTjmtS9ZhNZ54vXDQ0baX/rKik3lbHS7qtz/0NGpU96D60OKZwHzDKVP
KolYjFDFEPMnyX8A3FPRK4vuiwlnsGqmDRDomDOEwZP5cTP6W8S5ZRcEZzIE
ZpJNmqJ0Cr33EA6ZXUMkXsHP56Aqz9RDFGRp1uO/scVxiPtSALTHMGz+0aX1
6D5JMf9Hn8dppOPQpu7ZA7hWu4AD6W4wdJih2NCGxgt00RjizqNCT7R1xGXP
tYyAS8WzauRo8UbNQKn0MqzeUb5VxqAfF2c0pOxZJHL2Dv2log9DcD9LEfVo
b69Q3fD/xqgwAcFoDO/qCud3MwZb15vqZvYjhG+mgOtbnO9dTKY1IfapHlNy
rnOybmlnxSN0Lc46veQig3tg4xsnXTSic2lxcZrvn2ekTTYOs37Lv1RreUYv
M1brgdntzyqxtpnIlQTmrYJf288ZUMw9lnCz+a62PppqztzBQAt7lUUI8raF
e7+HVJtsxYJFMT2pFh84EW3f+6Z4rCsN5eN/0f84ANBpKaw5Y2HLp6UdHAT1
e3CE7qMOI3Q90ANa638lHn+QoFkujcwvehtTEu/EX7cWxwZfgpgoilQQQ3/B
hTw3/ptgTYAK9eqEMLyTkjRjGr3rI3wH4JfWOleE0OSCwn5CFXSMNMF3o7NR
YPcJDn2RDq4VbbkugpRbKzn1aj+IAmnAJhvmrmGP3CqX+HMoH7fZ9TcW40B8
DAFQlX9IWClRouwVQwm9yOk38N/6e3Og1uQLvolGjNdyyBqJwJFHryXiUA6g
xbHpWlS89+poUvx+XLbIiJ6Z4rRvX2Z3uCYPBJMNhC4JtF9MkhSaeEWcjuuu
glZ4IFzh9vGq7TSNPggQRa/sQIg/uf4AKvjecRSpM/hdGEo3jubbkR/OBaHM
kOne43P77qhdBm0G7y3aM9/FpjKlMCPBXFeOa0S0V6fZzpvCEn3xrCGYYkgf
T9DL9B6ejTXuIrnPCdBfO+ekQGYHnx7IB7BQmguIwoBJeCPToEW2sipZJZOg
xd4WPkTmGdfKmakblO3cn+8RnMoQVE3tDseOGVD2jcDJlRWKYE5CoX7Du7Jt
SoTYB68MGv+j7WnP5tSv/CSNiFa28yuXwmDcLNj24G3+V0EUSRjAAMsAlxTL
Wg9VuiXJfi4RHfUfnNosSTdZqUWloZKZJLx+QI3xva0q5pM8eJkxREQKnsG8
Ie9YCb2HCihzTdUyxiniyMC21T3GqHukKqfgDb9dhzRaZMNhme/UJO/X+wjT
lepbmCukHsa33Vtn4hOY/TitF8X9d2uDJiqw9HC/r9p8m+1sR6k4p+eEfxUm
0US8uCfJv63RoNOFftJj15qS/Tm2wPy144RWr8qT76leQ0sRcx8eT4Pxm88Z
rg7ie19c0vtnTs+5jJCw1eGUhWJq61xNp74s3RDhhtf95hx7+jZMQsl9OF7r
2uPAl6FurZcSohrAGBIrb8KWL6B5qnwdW3gFD+etzCowJuN0U5HXn1fEVAZI
S5y1gSW2xTFoA6Grpd4hm0qVZdUacKO1wqSQJqMHju7JPqhcYm2Q4v6jz1PY
WBAjT5eo6sBWMz5T8gK4GFwfy91PcYa5WR3V+WRWHGYJBW/aGaYUDaptDzuD
rRLRLa86lrChNJqNbMTPghb5DwYjE+kK/DbaMZYTPqvR0WbBpM3xJr/NpMzl
42vjHBgUPIV8FW2yymdGOs4EkolcKWYwiGd7pnm79TtymowioItCkv+UfS70
Bs059cFVG9c6cEwjfhiuXqiZXc8VKyUsIAvZXYwJKj8+yFgVHLm+2ZOs/I1C
uMvjf3nOCSM1FMq6wYBao8BzKE1SKnsjAlVfNtm7udXiNyQCt+I/85DJSU65
KCZE6Ac2AQNyjQ0DaMKg9eQc+cUG+mrpYGfYmr95HNTgUHYLVS/2Xieqvg+9
+NaXH0b7W7yQ+NTlVYV/78mws9bCZGt8s08bYfqUXy63SLNrfeNsxHIrxqnH
W1f548pJz5aB1SwXUlZbAsReCF+UVBN4dR1zqzLbWXV8l7UTNIfl6zq/65Ig
N3QndUAAvMcc3BaNnM8gr4Ylv0wkHxhAeGLGh8iguN7ORZirl9+P4CtoVLqi
rPJo1ynVCvQ8Nc1sD3D2yjskX8GaN262LgHQd6j8krIaWksgQFMU7XaeeRm4
LaSU1gvioHYCpLf7CJ0BzGBwGXly57ku69PeoarBVpS4ngBeoOGx903eqK3/
HNt0G8NHwmGO87DilBp6Ks9B4EdosKbXDIOaUrwz6RsOVZX1WQjKaW6/+p1k
VkXeCcKjeemWziM7VjeXde39P7R8mYGxawNhA1VmaceMy8aKZMC2NzZjQoPg
HOJ4oTJyePFX89OLo7phAJTWxFUnVkMqKVL3vNxBMx4pXJHsYfoBnxhbXcak
WK2RqY2Em09g+q7Cbf41+ypEJuo0pMKu2TqwNx0+Ukd45wMh8aFFaav5q1cO
CZTSe8aK5/XFBGabkD5XD0z54liLWBWc+uB5Q8AV8BtZVCYzqdcU10VkOu78
Pyxljm4JALvCFBhAOZZc2P511+FbLMsprasJbccHu448a7T/CleAN6+/YIik
0TwAvJjSjLDCIfxo0nQNwlfNgQwyxJjnbo5KUranvD2EFPxF1faAK+OjBNoi
Hj9QEMlvVHugrSC/KxhGUZUkCetq190/tHnEiJA6IdRjSg7LeTbyDNod6bbI
Ur/sCMNgZmeG3rm/d/gDm9HhxG/fde6hHeEMa/EpZOGHLFZTRAzoddIHKZXr
BwjiFwyl3OVCY65ithBk4dpvUrj50CmB3qPR/FW4WWLCTLJzyMqNDZ9E5u8c
AA8gBNIy2s/P3sKdCUvRxzH2vhLrIqhWqzcyfzbhZoISV+DGVeWxMtz2QzHk
BgdFhZseb8ZjMaWgNq210uh28p+iQSTqF+u96GEtXjlN6BsCmcGJajC07pdJ
qXzZc4G3tmGqT1nEkzBxH+8eqmxS9h1gMpN7hWRU18KlxD96vWdbgKCkuVUh
J3CRn45XLkNJCL1DgYgUovluLQwSXJXhFcWJSorpOO+M3C+FjN+Uwa4GFVGh
tGQHePhfCh9COLMkK2ztcmKCPjjIYVuRnY4XXHiDBIGOOIwS4i8SUk9SeGvP
UEZvrhz0TFQ1t91llEFUfsqbKyteSy7drx+zhpma9I5TakAPeu5AyUJlDYCr
gVMVm1T2vEdT1V5VoPE591ebG9JJmMCxAWWNqxa9/L89yPJmumy4RLhfYdk0
dyT5/zeQURX0tJQhhGFHtolF5UVz2bzJr6g0LfDCJwUJBAQ2kPoAevjgPu/k
dP8FuGlr+U1clkHm6d6QlGCaqz6hKcneHQEhebtuD2vNLvZQsr0ppaucbJX6
RGtZPLDgfhmCW4aJhMmevcNQUyXm477zbcbOWHTz6HrZoeuClBLinNqAjQqr
uIFOlYBDghuNiOkVsLRrci4aiOIDfNa/O8FkO+ZvQdAlwER5Jx3OZZP8P3zV
/56NLMKnDH2/qJenzL7iPwyT4uvJxbaiaW6V8tsJ+SNGk25nXkZi2IGtHOD+
UF75dJDUlvBhtY0RHWdUY4YU7vNb5K1+FKtRoeAA5NR/aOaYIUMYrVaEmecb
/wf9tqkWQXatN+owAD25n4xXMSSOTYbbj2iKUiJv88szGDzyc2dYV6fciWmJ
GsfElx2PzNha3DbJPfQnyo9HtECLAcMhxqOLvxCBQ4TcPMI9XRCXjpMT6a6R
x5n1LZo/Mau8PnjVsB2QZkUi8sgSiEKJ59gCC+Hki43YA5t/+ZOOoKgIt8vp
SR2czJKdUe74GFqYVDB5nyWIA9WAiGhdNu2+DXS5q0bAfQAvlCkO+T4TDKbu
+cS1Y0aSIifXKYpQr4ExJTIlvaSrmkHPMt8aOOO3WACgAL4m9Sjh+yyLOfyt
B5ZLHodCm/Tay4I0cJ4Oj7kxBNISODo+Fl2eeXDLoESYuMMFBrQG0UZn49wV
Af7nyq8WmdtP0uqRhTp8h0qQCOob5yKF2EVkzrgytmK2e3KowGEsVbAHCPRH
tZbUKfXXdbQ5ZqdSzuRx0Eb0xQILqNSldjbfYUqASl1J1tBc0+IBo9f7CZFb
U41NRzdtcQWrwW/M537C4AETNeNVtXa9hm9EOTyQ2h28KZfXJD3SUZeYM03J
eTD/7K2TZIpG8FhUFaGfj2Ep6Q8+gLSYhxvE3DsllrJbXISCivvmLZHrPopa
0bwN4M4+F1hdVVBdYanlOuQt+DeKDkKQQDPemCxUfRaFX9F6/nZbgMEEoE8E
QpNJIQ7HrXxvo15KYstwoTE5hHoTHn0oXOtDKpvhIwKNGbBzRvwY3gxFKD1H
p2uxZjdCDS24B5ozO1cMdnAhzpsdDdc7Z4FQ3QeQR52r1ngC9UWPhgZYyFx/
ol3EeQGkyVKXld+wyF7CL/nzDncMMvGRIFaSEQSKn5gNOqjzTD+SwoZBcj3o
6z6HF9QSZLIwN7TMYdcFMhW6fxMWzbV45q5g57eOnjs6Z799PSAaItn1+mxS
V0ZPtbo9F4L8ngn0sXBb6LysJtobdD1GiCbkcF04zrrr7uYrKfugOBsdzDkc
gI9NQO0gJoV293cYFXHO+rwf0chwusJtwJk2t/GPpVmc9d7xEdDak4PmEgWT
4o6pcsxqucKBCGwkTDD5+dr2vpPKzKZLO4lIx+d4hUEJtJF0zOx44boYeY4W
e6LKcL2BKnXyhw42klOC046SJSiGMGjKAJh1Z1C1rwQWC9zphURTd/JBVe+M
b+yK+kRW66vRjAdPDPxwFRAIZc8zTjB7q5zkm+Pg6aEsgrtAdfF7DX7+d3dh
9K8F5GxOYj8XWWOj5k/aV0bU0xoIbHsVNhyiCKQ5VePjlDq2bvr7xEk/wb54
Bc4hJp9zHG0r/olZPaIvu69GerRrfkLHVx+73A403HMb3boRfH2+wwOB9TUy
Xu1tN8vJ9XMojCqrwHEg1p9yJnBMP7pSe2yJePeuyxobN9i1JTWjA7vGlGeB
a++g6KBvy7P9ZX35F/qqrJOq34XvOngYchfIBmUQidtxSJ88apeXSwbyxnLa
KUDZgUDG2FwS8ngfbFztSs4irK97pXbTL+r+vwhk+2eX2w8MKE7Pta3vKB90
epZnD4ybH8bPn5YDooHWV4EDnXq5UlwZsWuNHRP3zFkVoIulH30BemfZolPc
t+au1BPUuN4uZeFpvzEriVLwrPaFuVMX7buc/MKrSDgQ8cGPTVFxUiCoEEw2
HDZDhGS8Ohxo/4geMHRTjf51qI0jQEn4B0sxYB8K+69SSuvNrLWekvi9K5Nv
TLN8wJUrz7fR/tjabotCQITkodjeB4JpfRCTUfWn4RtXCrCkFU+heyknAU4e
FKsWQ4jxAhq3QkBxcfBlT6+fpHNRu4T4+OGwvXio45j+WkSlE/pRq1WmGMpO
6KIg4wp1qD75QPQNqvsgeWRRWDoehwCSlEWFDvzwluy4H1J/9d5SED2zh9Fe
OpZwSBmIzJawApelABGaQZ8Yn777x7VGmmuOWGVQppvQ7WZFKasKW4FkcooT
o30am3XOPPxMS0jnPnH4d9mLg4Go9aPTPsWBr/hUdUPP07xj4+gMuVBDSjSe
gQVgsvXwuPg3cnfXXQso8hIn7xjPJIqszN8Wcx36rW0jkxBPe5jREYYpXzTQ
ak4F0y3uB+8f/XeRY5CMU6ls1vgV15yEdazo/4Eob0Ld2j8f6PzpkyAVzr04
Jl+P6QezeUiyRrh8nDGiQZb0V3USqcVOW/I/s2rQtIA6igjoZhHRnl25JzKs
X643yyWLnCrEHP5JTZ02Tvuz7h3sox/jfHzuERZVRTb+mczDMaV3x4Ms96N4
T2PHYExHC2ABb4ox+AEgVdUm4bIdjjYoLK272y2WVBHnO+rEVdKzR0eo8/0a
uTm8vCYMIcxk/nI/UvOwZVe68f30cwoUlXdexqG5iDm8qTgF+Es1EYfya0Wg
tObUQkthsnH08D9ww2846iYjtmYxOnHf+Dst9UpW3gDtmbMAORaIstX2WWtK
pKN298mUU6Hpyz2BioSK43whgXY3PfWb2Bb16CbAimSp14YgtuBBWxXezXAZ
73hyghjQd9U8VNgFdZniLpahTgfTa9CX/vwAI13dnACw7OR8tZ2wqzvLkaXE
vml4F1HTweSijOjFRiLgJVGeA0H0KpMKi3atRwyezCPpu3NbLA7TKdDUZFJz
X5thFRk4DWftNf0/+7hFD3SGCKcscgsntzrHt7PdDXzmOdTJa+Mj1ADOawba
f7qYTPrFufcU7/HHn1TnfnFgM4BCPOyrFnHT61M1J33FsxzqH+W+65gbEgH5
K98Z/oFEWX8S9NnyQKFINsP1+UuciV+Mie36TFRk8GJc9Q/u05f7t3tAfMKu
Zl2YDP6r5aCvfpWplCkRrhB3Q/pqFCbJCj4qMAZNu2qMbl5OCaoKoQeBNvqS
iigh9Jf6mVFyuIZzRTn/DqpER8xpbLW71ImSZsuhrImXfEWUVVUBd7EVAzjR
dJHfu5V5zIZERbinWsBl+8oal4snC4M6nyPAu9KcF0NZFBiGk0t7svBr78a8
GLMbyVXsc3EFtLUG+PpIGgVgypWxFudHDdNu0+8jcjZlpKJQubBmQjqJ7Ttu
w6JmwX4OhfCDCOs1nsKM3XfqcL7j6zn+XKBzgLMH9y8iOmi5VaREKo9DBiwq
oMxsHD8EWHOjvYfWWVa6rv3rJqfoou+GR1qYlYWM1wHC5JeYyQC2ZcCS54wx
1zl6EOx3zgM/9gJGFoZ3P8cgsuJjHuSeZGR/BJ/UC4mXYoUJ8cNrdw8ZQnHI
A3YsUJ1jglBu/3smANzfTZPkO5tYODBC0SYVHQKlEKj9kARA+Xzz3AJd926v
psov+d4okU85ogpMWuX/L86jFJPTXkr+RqYfd2xSFaZ+ie+3nV/Zn2WVqq0y
5/Ewl4PiTkTCslPS7+saVMu1sCK2STC7boaEga8D33KYtkflQDin87yzjVSG
c1gIDso/KiCxh4GDQulmwPSi2QyCmE2V/m8lwyI4bcW0hGfmMYETYPXFhf0S
xXZpgeOqoNZvO1+4AoWjr4OzS8efL4PtAmBKRqcSTgkQNa/O7u8toq3cOFyC
9Wc+ddCegXAOmyAozjvamV9BCFchG3SHYNK1vaJgTXnbFcaIjRHXObcSHbl7
j9s2cuteHfywRlj1f7TGAo4YAZGTtI/Roq2UzWVM+wcr+9G54hMIl/JKAPml
x1wcSuHtEOp0m4aPbDysORi5l76p0h9eTxERk70eSfCbVLakdCAV5TBMeZ11
CdnSU9Vqc5F63o0QYd/DpKUEwtM3Eyl174Xc/O8YRof6gjz8LcKlOtJgncq1
5VhXH+y5OuQ+KqegOuOsKemQcAM3wwfSWK29/rzmOkcacE1IeBWROMfws8xi
utNMpgj5SI80zdinyVqnltlWzLRbt+MpeHDdbJfClpSSpBVbTZLynsnEJegA
3SS4kBeBWbo/Z7YGI8FybDeA8l2oeStAwgk1R4zIRq62A+fmcI8HRC6rzVBz
/Gb/+2AWAGlSZWD2WoN4YX6WleAciT5fMhuNtTdo7GSfZp9lwaB4rFfmyr+r
2o5u2MZPWpi2sk173cUzPGPgjFQfKGif/yZP840SiyiQA7A2obeO1zVTjQm6
8aIz/aTKAKRXqIJYlfATmh1PvXGhrDSRXX8BTIp/qaHNcn90qISIEALYP6FV
Nc6nXd8ewpkaRJzfQpZisbjK2EJHbDUWKgjW6WTrAsiF7W7bC9NC5hup1BJ7
SaQGT4RVPcWpkkUiIknFi1cpNlQ8fjL3MHV6kHW0Lhpow7H4p1rEWzxpaXqD
uth55mYvqZmD7mzDV3CF/kSnV4MvRikn+asoD5AiHaOjQROEuzPKhWSd4DCj
3bE+Qpy15dGXRdVzIfcMRqXJiTE4fWGDMGyRyll62bvcBc1atjM6pz2MNcxl
vp0d0RBisFomkmYrdtBv81P0R4WPbjoUtfo1QFKb2dCXwQ5WQwypyAsNAON4
y21BT9NdaCEOQFxkHt/KK0s+D23M6IzctaIZSCnfuiyV0YjnnXY5G5JuA+wA
ArUw+MSzMw0EmHXNZADk0naMhtpo0lYilLVvLKPHS8KiTgxJOe+U+WNugOPh
X7x2dITkGzx0WJthedrWYNG685tV/eXhOmF4dTdAPbRsJIc4x2HV6Rq1gHy4
rpjwBvTDQnfSRaYhfTqEga73+KnxoiCLAs+B4QXA9XwcXEavaOLbBuzZ6Asy
cz1V63Wt9PbLlqGPHFCv6yRWRt9O7150uDV1IYcGZE86p3jgyAPBjSSnnG3M
uaXZhhnpfier+yU3Nxq8jJTqTSxsJO74gvP4a9P+4aKYb9aIs5El6QZWVTrT
PPBsw9kYDSbXfU8S8fn13xgcWBnkfynDxMFt+RnPJN1TyHlHLpB28jB/719S
J0nr5nHJb2xeT+uX1qjR8LPgxUaJ53icVf2fN4tstxuXp6YGKu0/k+fk34oy
Byzxjtq3tMBhPIyx2IQTxAzPLIEHL/6oHU+Ahv0rol/F2xpxTo7BWDDzHwSu
M/Q6UcFNIuUwja9qarS+KjX8ywFQ3NOunNUiAy2VrzqSgReG/WuJx1es77NG
pg96sUyDU3vXlVLmsnDJlIRT+mmVZ1Ucldi7tuYhe+dR3JkLbir+Vv2gsxc+
uzju1G7SY/Xc/oL7Xxh4lBh6z06xpCpeXYwiDP1Kpfbr8kFsDvESZ5hyy/mh
4T5iXMyiwp60zru1ya9nLv8zRQ2REMA4/pVvQpyWtrGjUlj3QeMRWvSooqgz
aq9+L7us+mVHDUUaURxQDbWC29+2pcSmCXyuWnMh1MRFJFcTgJ+U5v1Dd7Dt
1Qd/WtjPz7LxA4lVkS4lfDVuoeY3l6zj7ySdGMlH5ZmVP1i4bE83Sb8zT9xO
KOaAK8fHJ/iXKksUuHzkgKtgfxjxQ84cUcFPaSfpltPdyJjqnCtnsGEqFL58
TZP95mALv96eg1QPD5uhxNMPct5b4yp/TA9tcWfklLof/TUPFtQ9xMQ5ZPum
gLnpaV+nCXRLWjSLASwWsjK0PfLOqb7s+S9bZBtQAmyGLF2NH97ewVM1LYe1
EL7Xemf1aFktfJBeamnjoug4YtRQhrQuSyrPTRZFgj25mdOWClRsSPqNdEqm
8H6Mb80E4SROwH58yRHaJt1LaAcEmQlr70Uo+gHlymvD0u5mkYcqt5/z5heJ
C/AQ8cVIBLuDG9aGzV/eAHrnMLkb6vNQLCg9G6YGCXSvEVoMgim0SlcIVA7a
D6haS3XdKPyYJpRcxxzfzcy8BSey4oKJ1IDuSCZii9J0S38PJ2P8YICrTNX7
HU1nj1HfcBcMTujoj6Di2S+JPnbMPO7g0BbZ2YbGBlGBwaDWncGRGB8d+5M7
jOWmq9ndu84loXk9en4SR08enI6E94OJyLM7vTz/R8NtLC4dmZWwX3bFvATf
J4pAwmYpS3DzDnnCPT9djIcjJ3YxiCyIuT8T/zCLQiMkl68dXff2zc6DKGiy
8vQLBCd+RMEzUygEPLlQxuD3H1Cb3zAJqQWClVeYlCl3HN/wHQYstrvjIwUU
0k7AoKKH/gXFK8CjG7faXUu2FrhfmWiz+gZ8WAvE5PgkQRql6vCBhiCzJgB8
mXFCTQAVis1jj9PDQgLy8VP/hSuaBT+r8UXsihISThIfJf1RSYYzAioSjDjb
t+0jvCcRq1MmbAuZ1QfVyZApGIN2Iz4OMOuLd9jhvlLA9DWlov8DNA35J/TS
FZkO4hYcWDMaZa6JlDsdyY5BwO7Fsnnb/ruEEyJsq2/Pav7m+29Z7MTfT/gh
7HiwPLEaimWt48jJSKcRdYKAm+0MBr9fNcv7yM3KOdrxkJ2smcjxRdfZWTzo
ak2mFhxwiDquE1ozIutpYRxMM8rSEHFA4Fk3GZn28fNl8MPS4PAYXzhaWl7n
r8b8nVESdeH6rwtWOJ6zv7wY02UFGEZ7mxvjIlX6vofiDbCOlQ/LfT/k4pIT
O7JH/5KTZQp+p95CWL8r24HoC7nDvy/WbtgLtVjBHEBnKot4q5MUjOnziMTW
0acrbDWVb7M99XWk5Z52zNlB59QkQykZw5y0UzFz9KjZCjjk9kSOCWfPj2NP
/SHKFv3C1VSPiUaW3btW2Lwjs3hHmQbBqe/1ws+CtPiFGGwP2WZcNgmZ1TMz
6VpeLmGumrr15W9fCz6YCqUQLVh4RK1Zl4QoXBCopULCRC2Zzg13DCrW9z/l
O3TGljV92Ob39Th9SUrtUx6MtogbgtWkacsRjtua61YD4EzXKo14J6px0yxz
6mBb+zM+LIm0WjaUr4fbfAjkhi8coFZ86MPENUj20Vnr4zmpG2b9hViBnHPq
WAjgYUNQDqVyvQXtfkF6Xm5hAMGzQ6slVf0J51J1XY6vN9Jigvjq56u6opnp
wZwyUL27lqDVzXp7/LIijDz+yi47Lx8TFsdwxu7dMwq/rCpa755LjKc9HDFo
LMskuhSLAB21YEwUmLjxWHpslzZfMDWMcA2murt3QESWvnGtt+5W3rFu+4ZL
+ViFoU3N3nf2/kolXQEgtRUTKYCpe6OLxELbBpppNXCEFb3SZKZ+BKEvE26E
BFDGyodbhokunyMpm+zrSfO3BUTEgCwF2SyDoFfqNYKrGajBW/lLbsS32CoL
H2YagIHyBcqe7roCYZIMvsBvRpYTmiDbS74EqC7cD4Sv65qOdo3ZO1dFnEgc
AmDKbhjTUarYYNmfTZR78e8yGhzSGxhFZwFni6JY4S9F9giQKF5XyZ0/2CW5
Wmk37f7rwN1VDnntFoYAQU8bvee56drbYVkGBz6kQy/KSX075JBdEsd3hr29
CdXnW8uTj2M09v57Vt3OJ8L6E5i3iAqDEp2Qm/LK8brZ7N9WC6WDHn1u+40J
0Ra5cIc3ynMoW8jDTNld2Tum07M4G13SSYssaIMEHqNOLGOurFVt4NR+yXVG
dyYx0ogq+Y6tfZoigTZOG8Q63p80gyAJc8xNU98yprQEwR0CTLrChkpefbe8
qIUZkxBZjOVFlkqp3Ara+oDZEXq9VO48QA376s2+O10vsnRHrOXl819zyJB9
bth55m+l+OPaIrWw0sjs5LOczQ0Xtk2iSxc+bGFQiuQJSolWbSaGtz97pdUG
KN2H3N4znhFJQuGr2VRboKJyR3c1RaJm1Pw520v8IHbkTZoaA6Xb0BUqq9pv
q/bkuRRT+GhUEB+5rqBymzZFYqbFOGULzhhYCnhXQfVO5J76jMetlb8u8DUq
iHuKrMxvwvZjLQFjglIkAbLdWC88oPqgGZ8WLIi7Nxx0hSYZPkZryKNM1pfU
K0M9Fg3mT6geddiHg0TRLe8EmjZkfrkmd3V9KvRT+xYdZjgfg2S016AXOUCi
XP9DHD2cDuw0+UOJm9YYogGqSpTOh48mJGtbWrOmHWBUQ9xidOb3mRDiqjDx
aZd5UYYQwkGoyOBxXAKUW3cDpRRfQnhz2DAjuqc2esfI8rVr1lqs5T6mXdqm
5zMbclnqTCseqhX1xWzmpVVxfumEvV3/usBNy10mpIz8z9LITfjtTJ2rFSda
8h8zGxljm5F/jTwAlAol4u7GQ+4lYePAF7WNmW9snnWOnHo/R1ApswboCWdK
fGmwHMACI6vgr2SakNZP3Q6YOb+ewnAxQsFfL3Y8JHN01BUrpn30ETJtQOv+
IufbxaZbjQw1CnXrPDJ6dWnki3Yhj3bPRpukkhWCWVqaMvkt/pS8iH7dK8Xu
tJ86U5HnItQLjUiNK+hcunaFVAqO2Nv0U1quERbR6GUnF1RHsW9zstlUwx3t
c0AXbnMCYPio6u+oUumEgHP+5TpvQfi4MOPNKdaOU1SLrj0XMnHHV0mtIeZX
2uanAgCpqtDVYlcaZNhYc2l0zJ8QE8XaEMZ9AD1YcjPEy7pvCPt5rapFjPDT
X3ePjfu79awRPr1nxrA9uyRrL+3T7htPamGDGCwjPPPvDqIoWs1+XM/7/UzO
yWUt7o1ZGbwtZ3zUqa5znyIDICjg5IvpyTvCv8mUHdBjlaoAfN1BVmx85nic
nI9X9IKP/zFG6sAurY9bZLzz4Xse3qmNr6D7FrkM1Uypi4t+g21apTsjxIXV
5tvhVetj/KipkB8Bq+mBWvYJZEfaVD0vHhwaF20HzCHcdFT8zAgGmY1eOWuW
b/Cl9BMkxYZALZL1Dkfby9jA1qNjkBsVFH3LeTEnY1bWdyTu9kJLGx87klf1
uy95MB1oevBRXj6f5kXiqBMwKLhqdoYgUdlQqUk1lXb6m0vmh4obCVaLWHeL
bGnHS/7liO9ePbs6Ov6Gaz0GCNDXzJVtEb6CCZf56GYFveLskLKPPE50BlGO
eL71IvFap+gU1T49seLLhcsRkrp46Zzo/KOXB1RImNsBwm8reKIJszs48oBv
K5Va6+zg1GPayKiXlB+c65vT2+IPSfZhSa3wJwzNZeFHs6q6X6YAvL2ZSMj7
T5rNjiV1lIiUndW/kgFzDdDafTsy6aI8bSCWPsdm0NHXLzxkzYm4lAo0tZ1H
2MBnO9m0apPFHOzex3FAlQh372PwbDlnHooQvIag1ofwnBTt+7ZpTvrsHMCZ
O5cpNRwVQCGAVtVS/kL4n6h2ZugnywvaoVCxM/VTkodUJ+7EUyZCXngctYNs
29IFw/u1lVE24X/pf/iySe5EgZHUKnRtg3/z71fitkeKIWnEi+CRPXymjMz0
tB1+lBfxNZUmYBEHY7ByR6YRplQLKyYnQOTKnpbSurLLPQ8DrQqqvx1cLacX
DzD8Oi1BUGAt1mqhK1oeND8whh7gGmNarH94LhwdjmvpRYxjzo6HurnZc5LC
Y7Cg+PgEvAjIUDVFUKFJ+10LGgTvR0HQt0gyXDvWm2es8+EdP4FWt59mE2yF
8CcdSlI1l/UPVxdtr1ydTLiOYuUztQYgp8GhMx3heEbGgfnYmJmQR3eFMoah
qpZWS6BoZx00rvdEsGsPOOYOymIBqChuMroYh0PKCLQ+h94OBPPbpmD7c486
k+dx+lSeZbR/hjfD8uzxjSTk0eD67BtCGZL1R+tn8RATZQicUwW/UO6aTss+
T153mtG6B2JLtEGkU3DNCO24RPckMlgvjfssBrqg557AOXBrBCTbwko20KF8
oS16AXHA/rLEWNvOUZC1sep+xS4bImaR7yNzmzvFW3aMva+940AcATY2+F/H
nMGQWdXrbQypXC+uAuIX39hniY3Exdh/3ygXrhLMAEIzlGsPjojqN8I8T5No
AVh6lrHTNmE25iI0k1jsBnvQ6krM16fhI0CWQAojMRXGbzgYt9gxafL67jGq
YBVMivGoGXFoaMMTd/3c49B5f9ryHonNaIjS2v9U9s/zAaV9y+iUz15ZGHyd
B2za8BJ5wJHYKVPDak4CuVNXV4+M2LMxaV+e1w0CfYpD/h7TZ3cIZRJatd1I
DoWFUKrJJipcEQdItFPL4WRixWnbElni6WG/UMqb4+P9IKpHCz7DIfcBsuCJ
hbWy71UqFTSrWqMwnR5Pcon2YBAGOi1iA+xqVo15L1z/4uOdFED/Gm3p8lRG
qmy1ID1JdpVtqOxztaqx3ZOi2tFlAqgUFbb/GoVTbi4kGVmnzJIv2YkSdwVB
yILcMxnxDY2NCVe5n7wxLA9EYOksMWDndiGSyQVQ20kQK65o9oAbl1QoAXCK
E8kmZDDx6EXvVSNqqyBBOrW7Yik6PciUu58WpTnl6t6d99MFlhO5fEWSuGKF
cVb0y36/HI3jJofRLyBIKsZKspNLtt3JhkzND6IuYnLAkh6ZS+j4V3kti7Nn
Uov2QQ5kNWb1IKEDmUbERttm2TxjDJvpQBzJLtk0eMrMcfQ4yZAfk6Of22HG
obKfOiZtTkLkMnfanIKtX6pv40omHQTxg5Q+Onmbv/Z4/dg6ifLBc7+Ukcww
hiunl+kJaZMeMR8uKYSfnumAExypYvnI8kFjVWaKurhY7ueFqc83Vuwr/jZe
LEz7Nk6hoyQxTHsPXWMIgXOAGv0qNPqe3rADzDdBGLxGN+TwfpalyExOxHyp
ZBX03NhUsTGffQXgEIof22zt+ljWqNOkMfZ3FrrA6y9AVoilWJ2jhhdo21Gu
MEy5NP7hDtn6KDWsrc+vy9VHgYhhqEfbMDsWjnYd5WBYTUETaotN6p/Rng0Z
u/qVB81py8ZC5EoZ1qrEHL/yTr/K2EMKk6stBQcULMCVMgUfuyW9gnzWRlY4
S3gq16gC5fwp7UAk1Jx/JfVxBC8wetUBLHj9d29r23/bmMccpaH0NvQP3Bsa
T7TvI7qCFtdvpaU8cIDI+Ko+6/PLoHA4NrP8W7Emo9HuA/tugkX8j/hEulHz
HrsbGFqQeUT/1Z+v8vaQyG/H6J3vkZ2e3ZQ41Y01SbgJ09DRdAQY+6ja9kQB
8gdgGgLOD3ePoh4NnxUgAPWtoJw8EeJGH/JDq724MdzfF/a8Oieb1SDd/SR0
e45hkBjRHufn03K0iZGhdUJSl2IWcTUYxL+THJJ8oQRSHW/HWH1wu8ZT9bb5
p6mpQBlw92LhK8qQ3cG7x4Vyzc6JtvajbAdCa1vLzn4emv9V3Cx+IVGkORNQ
vVjRmCbZNrvZddYgij6JQmfMYXAwYdUTBrpS3H4H+I8BlsV1Id/x9xP1dewk
o7zGBrhivsIUe0pzwDqtouXOX1XsVAqf0BX6zUAh51y76HkC6cOSwTmTh99k
X6ZMj02ZMPOPP1CghhaCaoAMEA+2j63z+v8JIzJsdOI4lC5RTEtwl/vAUQ+m
06KLQXTHs/j7AcLNhv42gKWzCpEXV4b2bSZ1SmweyWGmCoZWcWUK4h2afVoJ
v6XqG/4ZD+C/RMZIAP6VDwmwgB3st2qAXfk8/4e0GfyxzeNSFrZyoOdwYFOY
zWtCremWNRX9uIrseV679EWwEs8yXGP8MUrC9rkfECN13n1cZXVAd13wacYl
1hm8Ejn0JRosIWn4TkqLUlX8S1pmxdz8rKIk6Kr11iUC5uJGFKQsdQ5TdAib
X2BuHaD1vLzb2VrHZfJdocqJ7sHoIVZmE56nq93NNxO9LPm2S3l/p2RpCKxB
rXmCKS8jgdR9jFjsXb5EmLv4MsrNXSFa+DIYI7mgnmKURIjiobVG7yXMVEsx
Ke2u/wcFmfselSIy8xp9y6z/gae+v6qwSjsN4D4bii7YoOvV4RQYljIBgH3E
P/4yuZcEuInusAcu3IzIwBRKOtrO0C7z+8wuZNAteLu+/cSC/Dxh8m/++nbc
sky5t8atyq59JtxPxOkRiGKmNbgWTosj80mpWGjCwxhgMoxGRDitNoSWNQle
JFaHYp/0K2prtBFO+c/cfkhh96NHQNgBFA7SqATtYAfBVSmddxRdezeUIloZ
TmRjEaCy12lkjcLq+XQkX5JjwOIK9gY0ZBnabJryPPas9oCub+cupoJDIX/V
Cwulb9aCSfhVgq7EdbLnfnhJmXlADL2YB4GZfc3y/tPmq7V6LEDN45S9a923
1dtpZ+HLKpGN4NR+UBSsbYHKov4YzkyuFUqgT+GpU+I2vQrxFEY7FRWxRgr/
wrHdYuaqguC7v0878nUxmTKE1HVyPws2TV4NSdgGVMpXApMPbSZcLsdN7ys9
Zx5eu/L7bJ+nme+I/TJRhodY7wP9lnffp+2L4QER14f+bcEkeCC+FoMbX11A
fplq1MqOuPUEklLTlUpwCzuEQFkcoMZ9MrFBiyNo5GL2DPvJCW1Q62fcsXgA
vfhRGJioTpSs2PDuWirTO7MvBV+rEtT1wF38SM4BEuGuDjs5p/dDIBbaCFqf
THkcRJMClEnQzms7BTuNXcXGEvfW3M2EcP9mT+IjJwtdoiXG/UJvWW4VuhOJ
rVb5hJBGWmHe+QWh8pBXEW5jZadA/C7YQe79a5w1Ia5Qq2NYMF4Sbl2v8oGg
t8EIxmsVDM1YiKM9wbESvcG3KhhCF66kJO5a0/+joseS6hw2q6/UAdfFntf3
nqWshCbWjkXapZuoPfNHs/0TX/mtsJMbQiqqcXOtZqrdfx84zH7mS53HBpoI
clMquBEZZW2Zs772CbTJ9F0zORTfxX2fmbmk5YwPbOTUDzl6/mbcDRVU7oF2
4BFmSWb3YDD5tagzcf3hidW1V9naIrhwqFB0Ok2SqMjHpRZUtRV67oMUt+oC
tyArDJGWZ/2m4cjlbvmr+1ib6euKoTFLWAZPfv6phGUcqkqzrOuKLk5e9jfY
X21P5nRPbZH8/LVBkk0jNY5mieiHLmFQylGshax4zDG4tVDR/6cMZ/9XoWS0
EttVvpys163xk0mKP8cH5v47WhAlksjL8KPYgOKVD58CqOwTQeu2w8/R30kg
Pe3UoQ3tfkJ6YS8JXAzdqhWY5c6Nc2ZOJwkfBDWnAfUD/hmRklDG7OLt8OBI
DvZyUlnxL0mK4riN8A8f+JsDlPi+l0K6xBZQCNx1DLMTvxbCQ7fVssorCmtJ
Zc+ninps2kS0BM73v3nbMzjwJQxtK5ao7WpPimBltVe0ghZPCWuLRYmugYxV
3AMPJMaLIRYyeqKl/VLjPQxXkYo9z0yrCk9uXVbH3AoJm+otwMSvzHI05hQ8
f4e1FobMSsSjWyN7TuUUBRS9+oluRjGlMLr+HG1J64CfV4UxUgkHX9gCqFWd
y/qB8z3W8kNA/1h2C3RraJ08YlcxTFuMuYKzOdR0k74K8O3UdqknDL8WUgLt
mE2Tf0NGSb8HtwCi9f1p9HPhlYVPqQetzca0q6Ac9jkO8t3fqFtjyiLQ+Jtb
8ipg3ahFdCEWY26bedwXjLbEk3lKtWc/BLl+ts/TT+Y8194A2MDZTWI+dWhA
kC0dfDDwZcX3r11OxoEG/8eYwDhqIF0MrGzkTJndxIRMl5DXEgZ3SacGJvOJ
8rMYEI/PYjmDeKRNeKKZXv8I73BXOlY1mKdIANGfx9vuFzjhCNNtbVYCY2Ek
LQa02GIA18UJHejhrEoUglcQLGIv6pizWPYAsZV7GmjK3EEQ09B83g1l5Y0Z
tDhDflPPwdhUaHtcDWVMkYtyMp3yjRTjYIWaB3wfXkZDvtpm++hrzkiY4jM0
irPBdcK3H59yo0Y7B8Ry4MzMQth87RTd+noUq0V7Q4ZQeBGISTSWorOFvYxp
YC8ECuxs+hxd8BM+T9JbM78w09Qs08g9OkZROopPoXuU4bvyTY8sdef84xBg
SeqM512edpPVUREE5N+o1lXu+cvN84ropgUF1289QOQEfwRuPRP2eWJkM1SN
v7l2XIWnGnfF2kWHBzB/KzT/pm/vYkNnVYQC6dKh8xhfl4PUoSGckQcw3QiM
FkJQYnih3ZCXtVm7qhfN1yKGMaIeVNV0/XPgsATSrLDejSyff64CuTJa2l1j
wm0KddV+9ZyVsxO4+zGIMeS0kdCoTwzHoKs3w1iwEu8DU/Le/RcLphtvjNRi
IRqarj6BEAj28baSwbT6FRjOriwH8wM+QLNc0iEbQMvn9vHcYMEFZcse3Z69
Ri/zjyGyDnBizvXN6zyqcovS8tJrPgeiczqyCr+zkwKcnrTGMNJB6N/zHFGF
yUXPTDDRy3p9VYLsXVkI/93Hz+aJOIFqO7PEC4tfOW0RXVmzwIqVbqUTg5Hf
4DMN6eBRWxPFCNln+b34fNZHJI4OB41jx0ZFhPR2tGpW4FD/SNYDmqJyILhP
+zAEhBdxHIG8m89Yijn/AjyfcCFOBzFn7P3qnK7eX4fwEY0EvdEty0QOliok
/W7+49YxHAwmtzChvqRtU3qHmjuJ/g+GcNpTwB077C8q4Yzfgp+qKIEF3eaN
RljU/7egA7LQhL6+rmfllZgcDxxdEW25Hb8Xrkw8Ow7BfzvLgeSeOd+gxsde
0IhXpN5UZODhQVpOdEnGYWTorWXltiZ0XfM6ZU9tR0TUKXdva4l/L5pV3vNK
y9aKdJt9mOaZZI337NjbBGFS+jgHt/gqwp5cngQjxpoQSxMQrF4wgsH/luZJ
gNTgT4XzY97fkpHuwXAL+l+TOWtgicVWTOOszCYoVB7xNIjmXp247dUTcQAB
GkIu+gh7ht0oSwnZ3sMwObXSqI04qSIemYKakKgEwxOXttZeKshOyo8iT7Ma
UxxVpWC25gfqLBXcPZPnIB/aw+fS+KPBWF/wbLv3Ew7xH03Bhmjz1ZySFE+1
dVK4Y6LWeoJ1pQEqY95iMET9r43sAHqTR6aSCmWZHfZlyIeqwJZX2Yjy4CEQ
WAhgOEjSKOqCFEC5RZAt+kXHXJuvKcsDCSpRosVW9QA/QRNvTumpZqOirrxO
qKs23lJNitHP5ePbhW51D8PjJjkmPcNRZgzj0b/8GgC9L992CGt2yrORd6vr
n65JDEB2UECpCHywbPNrPwkRFnlT+doNOJijtfqeMc7gO+2J5d46hsVMxik+
+JBWEi6ctwhvvpWOqhxtlcTaufgiWqLBVUNc6F6i7sd3QBcY+cJaWpcQ+WRs
DaTmUy65FftS+WWRXlW9S3I1KgQRnvZjrZw3vI9CWbameCOs++DQtNZPVW3C
K6WcBA4quKpUEk9TwwFauQmkgnW4CTQIlKTyRqs686wFJbxbgtBVka0hJWOR
Bz2LNsafY7ehrlmzP2VXggR5pqZSMMrzX2HBjqFAeguNcwGxHpyGaXbN+bvM
cGhz6+Zu+JLJ/6zIj9QSgj4nQ2VGc9+MMTXBvzikPjLUk66W5v321c7/zoxu
FmwVBWQ3UcCBB6bZoppmWX3EX3gSQfYhE5m4zU8G8+aXe9s9FgdJqB2YCNym
yNv8XlXUMraCDqj0w4a10EhEpKfaG43Uu9SbKU/C4T6VU2sTOK/1glY3edIE
rH0eOurX+ur3MZ682HTALfjI6buntIushByO6dBqCe7dGGl7QrGtry0zTi/6
iFZopGNKYJ7mukMK+3UOlP4KyV8rFIObt+N68D4h6IBBt1btkrNPUiTpxVT3
6k/jTPCHdvoNa3gum8BZcT2MShKw84m5GlivT6S1/8jHibP6heWCSZm6CAjv
NBr0LvneAOaKu8kRU9mnIliu/M+BUhMqkngtbZZdpdCz86SNvsmD4Rf5zt32
NbLXTyhrvFIbUbB5Ec7KCvd7BztQhn77v9+QPBx+DsPSAtSLuOGzOqinjYuL
gkOp0g4IHDmafjUkyOY54Nk4K0xBa35CCYwXHgr+EpfE66+wuUeKwKMgQcYE
Pwyv+PqpjTYBLIEg5yZAac1jDfZZGzylEcGeWlBDmQrrnDH4fvQSAo3YT46y
5SQSF3jBGh7IG7NOgwaw3R5wWqCi7y9WZrQlifFZzUc+B2wzL8RVhhpNX3Oq
8bzbRQP1UWusOBCPy906OMEv8buKNBBIqK4wwT+fHng9JFdOIflL/AmarchJ
sP9PDTwui5YnWjzyc7svD0XrdFq3m2EaIkopHqENhhlZ/oFEYUTq96VWfHOj
EjxvX68k858Ppzzqhg0jxeQcqgSx84kd+qskHFlzF3mt7ONUUnjA3OjKOLQr
oE/VRAWgJEISKl8nrao0QYS/dXtvX8meHVGIyNySJnv7BUxXr7BTmXeEX4Aq
mFSqdc/8ti3J/f/0RGUVhkfPt4OgeLjwB7ahJFs8Guhm2hF1qKIDpfbprahq
e8BUubaYbIvdmDtM+zml0yvIYrzjpg1DGX4UuZE2vinMt2xbeRR8wfuILBr5
TSwc5G/GRNT2MWr2No9IlQGOSEv8G80hXcABlKBO+RBMSHstuyf2gxLY1Jn7
c6Xau7ixhMVJs8JOxXiRCK4l3zl3eVwvfWUkQHEZ8LgKbwerbbJ1/RxOb9bQ
KKm5tAx1SsaEoIcnsVUXOtYMpUdx0VxLHlfF+DfpEL36VT4iGWj61TQsPYp0
XlNK/dF51Rwv40GbUP+2W+r5dLtW2JEmOlLkbRPBkoqTinx9QzXutm+HI0E0
y0Q8FlLbwM04GATunWgIgJ6Twy0YWKW7X6lrSggYMCOAirBG2rkv6VR5H+tM
DdOiKAQgRR5Py/VXDFxcmFGL0XBozBnDX0b1iG/8+z/o71dPPn6lluV9u5K0
+zf7Iq4SQtdDzKmfyqq5O4yk5kHltWdh146UH0sg4KtYrEVGctNSnriRb+KQ
wNW0mSi4NOt/3i5drDG6AUfp548orLqRY3qT5K/U7eUjyE/rO3aZSW6jESA2
/wBNvQvUHfPKl9VdM57XAN4irS23Gv7lU8pQEc99GnyJl48yseyMPEfpFDHl
5wjbRDt1vavoKPxXeiXcugWQvfdp9StrVYb+46cyimny3A8R6hj37LbJAxBF
5M9bmRpyAa+uWdAs/4ivDWjbXAE2r3PU+Qhuk1QDLweX+BiAHi9u76pysGDU
nfeu8JtFk3CeVemdDVikrcVGuYgsyJgS6eY/s2Y6S4912mNMLsaT//nSUp1K
fwKoyWSUwYDnXeniNaDOVr1PlelgqwWagXjrMRl4bsNQk9ou0oPjqoonHSxo
wO77k7y9uwlxNneBC+9vgFtPAfAKM+vk1XgOg/DdoyIMzKdsuVlhOKlfNNt/
rmAuCxamSuGUMvjORdZ3yKh+wrlTc9HpP6WCFjonrKN0J72NYsRNS/IUlHXJ
fJhWkJt49BypZhfe/MV3FdEdzbF6B+pnI8bYa8jQjqOEFxNLut5kV7WoVdWV
FV/85uIJsEEjVioWV8d0MI4Gg0bmLT0qKJ6Il3DWl+2gm+5X3a4V95X1QyYK
YXlWYM6E0XzJclgkURjUGjQxKYUppfsgBd49C1ZwTC/gD/5/uISXTEPW5WxE
rm8AKkBcbKJ43v/rWLA2CQxKv08SQoafogvOPczRC1GwqKBNdWvsSsGYNeUd
erJqN3xdcwvqb1lefjsKam43071g9u8eLaU38s+BxpB82O9w7y9tYGYIhzre
KbNSadMJKj4WLYVOxRI2VS535vMlJ7TSLCEWdXPbX2jo1qj1ZZbpUFdfiACh
4TqRsSINp99pNEgfvcO2ayn8ALcZ22tb/escFvX6W7okeYJz2B8vsCofGgl4
L84heBjuuBJ6kihuO64zlnjzUVpaEghhN9VzJA+pXoc0QbJILRszUEMt4RMf
yCVk9jBbOqAWQ4N5GgaB75tJsy02fuX2FZqB0VRRovleSXE4ky9y3/2gCSVx
lTuBS4suBIzRYY3EX5mEm25cqhNrKMUgdY8t0abja+o73SmV0JhBbJwSYESn
JP3ZcLzsVPP3gIFXHmlOd5F4oCaNNCZSybax70arqOII8nEnswWWrmWIjmvz
3Ly7y2Vvo0P4H+7lML4YxR5iWnKEYSwWZ5X5ODuOSkxe5oWa/saz4M1ooH9C
71xHknYbDRvGFlWiSpYEzIelS5g0OPguYvIkxoK2ibX8BSv32+fWayzghL1m
EtuWFAzF1D+sAUDxkQZ5qJnbXyWKPeWgLT3augzKlrLfvsVJod2hFsgQWS1q
2/TwE4I6rM7RBQZkKMuAqe7fVUa7jhbBSrf+1YyXL/G3XzsoR8Aev0BZ/zaF
CyeWa5/gGqNEi1Xg928xzHc0WcFNdp8p0mwv1z/FXdfz6lum9u0xm+Hu+0de
eSLSK2Br5xKVr4vDO2IVOTCzYOkz1xP2x1jegP/J0Kv6dgwGASuxV2Jo4MEr
s/wkYS54V/2BqqOE+yGwgT6Uqp5ua6sufTbOGDYhkvIUy77F5EsHVjD+uyPc
SCYmUvO5rF4H3VJ7EYmpfHGogax8sFE6h/8o0UEbTLDCOO+pVZVcbO9/2/Y2
RdPHxRQJ7Hp+Ic4TJ16ia/rMfJkfbhL1Qi/IOwVkxh+YkS8cJvXzS8pb/qgu
ho8u8ZGhgBAl8TDh0bFCNaCYc9DgpXU+gPBWgxJNjNvr9XVEGNTUYRNEfMpQ
l+LzurPyoBuyqrpbnqBPyjjwTuq4ROiwJtBsLWBr+k8RXhwOAuL9zY2jcYTE
vdaZqn2iqYGgQVcsnoAeJPsRnG+wYEnUk1nPl+t5aVENhVKsNccyARHolNRY
43DhlZQyr815PcKFdMNR97x7O2hVkI22gShK7yiOOA1gjqo0AXVzG5s+zozI
EzPbqIOS0pT6eNAikdT0O2IeySuHBH8IB9IiAlClt2nw8ZQTjiIYX8czaL2X
ZlSOxkM3plDXh0DkpSk7ppnwdVpxmhbMjzoIK0dy8cn1ZQwiv08kcNVZUH4S
EhOfDQZj2G76qNcnUfHULAfChGlEoDDiNozSu5ZkSvpyToqzZuT0G9zSwnxS
RgLg9K5BslMXsdvUpcP2uJ7MS+KgMdfavsGJGuvu8/hBXtKl6rxyJE8qMQ3R
PQ8qKuIZoDR8M1L2orOUYNrwEKX6JBtM7yrdttdoW/qP33zjDDx5utijJBcl
PFwQfUj7IOWV0J6FOvxISRYAqtj0SVjLKSiKSp7I0ranx3ZMcZqb/lU+tjkE
bhxOHg5VI+SWzybaqMyexU1zDMuLHVSL61hc7kHx+qKf3T52q0kf1BKt5sFz
G7C0bce47Zmf/awBO2iAO4mk7fxEgDSAZFweT9/8JzC4CbLLE1da1lrLknUz
b6pOVbmlNznAXbSpCfzX3UeXGjSb3BlW9SPTbqZRxQrKzYPkoe5kbKOy6t81
gTNUOi21g5IUY9s3mCBwjZR9XBSh/BTPPSr+pVEs2rilS2rl3Qpnd7fo2p6X
F2znROJ1SRfHyALQPmRTRfuOh43jbKRf+wBZebJJVF6dBnU2klIwmf+M5ykt
j4AJawbIALjgWcCeo+R6DLb1eDH//tXCHjrtL8bpo4ce5kB6Tn27qvx+q9tH
ihMIoVYpvDzo36de4tna6Hjh39mJY5luWAklh9h6QePBGl6QjRpAfxsj3MvB
Kh0Jcpovbj3mxZApSbVENuVmmTJtN7HOm/kDiGNVCY94Yv/I7MFQbLsn6GqW
Po8ZrEqbnOJRHr073P0T/eamVm9ditXsKpAhfEqXZ/NeunhHoWs/3q9Xmjo1
IZVf4MHlamn2SOsLqIwgLrwnn4LcEMxUARiDHxW91yK/acFmd85hNLekTKtN
LCj+iWc5Sixxurt6jimxb82Zt/+7Tze1JIIupmZ5CennUXc6v+3I1fBRZXhl
DgcsQdWT13DuiKGsDMko96kVdwhw6xxz7igXXsuv9cnME6zOuyMAF1DfIJGi
ycW1PLsBLr7J7Q7yoRwL6XIO2Jcrv4GrJt13h9hpX/TLXTjtlOKXbY0Plmg+
H0zAZGWp5+FiIq7GO+ZcdFycW93aZXYXM+C/JJSDpV9T2opKIVMsXqEDoZ6D
UaRW4rOfPVLSSNn4aGUfNFoDCU4we0dGjj2sVfHsSGpb4O6JQs/fc//WEDQz
68w8/QRLETMCDqgER2yMn2INLqEkD/CLc0OG3MGDjRP23y/j6cmdUhyATAzI
Cp6l/6BVwoLlabQVrqe6gEk81gMovE8BOEXhwJZYp0V77tSthzSjEqcQPLqY
lS1XsPLnexQxf1/rRKmGOnlZcHVnhYcKGyWvOLUk0GMOwzGI7bOg3aRNMenf
kzsbVG0K3u+/wWwZ8Yen0ZBfv0WX8icBLMk4xDrtBP/AYBYX8iHLdn+NnTdw
QG2gYXR/dASL0yDCP2ZKZ4pALCbBVuGIRWl9gCHFZtGMAz+lMtU4dIhVl3X3
9XMTH0hurNGbifN7DmxvvKKuOKNS6F2pXCJDQTaEwzZ3JuQPh92ACylg3mJs
DWxz8gSOD373pXhpFCMcC4+4T0YF4Wi0TPh0kZW6DJUYzR716mRpaaZxQeOR
yt/o9adJdilWG+YK0MIwOmnD9Hn9q10bGj34sFKcOf0sCsXuhK/t+5qdZCfl
orgRZyiKTtHwvXm7Y+DaN1GuKCsudQ0hLrFArDNXpXpkYekUKioBmoqoa60b
i1kp9eJJTFb7yskvy7SO7VvumkVJaAeEzJ+Q72JP3NdI/omJCevb7c82UROF
E3brotBZDcF0sm2gVwk3gVv2q3w4y5xvA11bXcVXIFLaKGWazkgkrPX3c7Dw
MXv6T9PnpLD0Qoot2Z+lB3/HPaCZjb208yqoE/uDg3K0cB4Bt73LPzzhXW1k
qZlorm1f30z7rndoDgoRVrYQug4xXaserSGkP58AcCXtTWrSfDzBQGtM+arp
vKFlrEQhedOGyW0a+SRr2Gw+xkNaI2aQ+s9baTDHNlzfvHW0ZlGe/OpgWhgW
DQ7dCNiK4KeGMa04yS1QUuJElSNzNTKud4uu+OrE7A8rTFlZZ7n7uLILtVkO
PknPwIV9CXawIE9MOLvCACicEgz9iUjgo4EmINHkQ+JbQD8m3RpY8aglvZmI
RiyEifz/MrDbgyCOUA5KHUfbDEwt9aba+qFza24rNPayE8x/fD3QUFRQnSou
CLqKEAwGQXBTzpFhgFdQ/V9NKmTZrR0+zw6dwQr8H+MMU604ixZ3skdC4jUE
7uR7rFApG7Aa05RRPAmGxrT2okUFvwi9aIOaAdNjX1nb1SfgwsbZ26OhyKhg
KOhSei5F5noaWUjtaEJQIiQhXdhPLkKf6qoTgQlcefVjHFKOglrvrFpqT7ZS
SCHYJ0uPXUzaoLPbxgPjjZ/dgdqe1y9zuVvb2mxz+sYWtriJcx5VRK6XujRn
eVt8yAH4x+upAag/y9FZpkim3NNFFUXmWANfHl00YJg6ZXL0roH5z+swfKqt
Euh15K7HHzXSMO6/tF3anvvSxtOIttPnIL9j9mGoYKffzNm2hwbQQGVCs7dy
Z22mB/RAmcXWW09VJxEWPjh7NkzEJ9Y2hLhBbyqjozg6keOxi8x3nxBGqA6q
v0UXTw5h6yjka2Jhoisu5D+j48MCcH2Fl0zaeJmfPtsIcUnWGh/u3Irnie+E
Rd0MjN/FrYmYFu3xg1oHqOFA03EX27dOlIpuKGCvVHQHC6z4nx8Gcq9Yihc7
9iEl+dK0D1zkONfAWzj7oY+btGEmfs7w5Hd68ZyvuLXuK2IAAuKiYumpNmxv
NgJv32JWQKMZm6XV4S3USrEN3dmaNRAi1bajH5j04s5xXCpOVpAE47N5VBnv
dMfRLT7Rvs7HkUKCbB1n7TFvYnE9gTt777yTFdFf6hbJF/eeGmlb9MdYzcAn
ZZmbCnMn/D4hMMlrw92Dqw+Vie9y/bqe7BtPi3VAx8xNeCqSd4vTmMiKtWMX
1k01FIOBk8Hu3UAuoDF/psOO/UwC1tuS/lIvcuhyb2gNR1KY8LRfqOpYk7xK
661Gp91Ka3mR6ydVSoWjfiAHRusO0Xmno7532G0P9ejGJFa5lNAsLF9p1kWf
ED0LZSRoBQgQe6VOEoKLIFyTI41SK3pyrFu6sGSjTiZhRrmvyO9o5mR98JtK
Xe+pqF96lvlAD0U04KcW2EyXp1dhQkFOfNGZ9fil8qhEanjpMG/lpBkXWcU1
CeOZARd565BxvyenHDpQ1lrddUDOyeuc1dUvIRT26BRrG4htGJVyXnxNEH/a
JpodEJbyr8U9STK7OY+PJ4G5e/CT/sUF+HNEuI0c7I2iskIUl3iw4hVWjDCe
ddWE+JpLsCXUs0nj/DL4i5mb6IDLgtzbC+aHMSJF6m2BZBo54QxnxmWcoFmd
H93mkgPXUaPv+k4B+eObcuJWoJbyKoAc1LK73aLZVuQCfydKBp1I8xhymlPg
8oOwR2nizSmep6O8SZ3RWhrNfl8pXd3HelxmMmB8H2vlm6L/KsolTJbf3UqP
csEQcvgyoMVw/DLC+l/mfDtXzttfeeQmUO9vFFHN4eggWcYUjt59FHdZQ6Aa
n13mcnLBkPnx/ote5uXwi6gIeyD87A+lMmMo7ADSv/B59mDikz3c70xIKKOT
X7AdooZJtMcfpdSQGXKanU6HI3Tcb46b8rjj6j7vZXBz+J+TYZKY24884wLA
COaBMEV1qZbw/1CTupYPd4lVwcgkKbJ7ziYTQvwLzQd3PQ0POpJyg5NUZ4sH
pKPqlkySnnQwVmc/TxAGIulxi3tIR1DS+eWwAg2+D39uuJpyInL0J7xwjImj
arIxeZ0XMQOWKSPEUMYxuVxhdbgtTRd9sPzSWMy81olfQVI8LPIKVUJ+Qb9z
k+8Nc+bpaHUWfuqcnkVAbUbi/v88ucQz3Rcvgq3nTZhBS/W1EQK/vcnkZVRI
JJj+RyKNcx0SVqWb0KVv5I/TkOH4dPK9BZCzSF5apUmzYTcpq2exCHpplDOP
k/VKQPKTB+8l1XsRuMTyuoGkA0sD/UOq7l0Z6beXpUNun1zremt+bZR//1ZJ
EM31ODasVbdBsNNEeXhTAqKO6fr/iU8A6oIqjIsaEXcjbftoagKSxU3JPS/o
kFG0J97NYqbfuIJ8a7l9lv/syYmDI7ADqH1U4NZFTkFY5UoeLAKVOYpFqiUz
uchCmToY2ehVixA5g4yyZoc8kqTXzn0zbMpxIVIJd5GxD+BCCMybeBvohuGs
Fk+N3hKOQhMDozBPRuNIO7m810fbbuoSj13h3GJIwYAUdcJMP0kGWwcEG7jx
O9IgXU434bK2wKatagzcp33rgB9MZS8gJrbZownJX/k7LdcoR1BUrQ3nL5P4
Hoye/lmFHXOS94JtShc7451Oav//lJKOqns5KSuPkvMJuMHS9jchSiY9+i0Y
9ESjHioDflA9FjXYZTeq6/JY0mFO+yJMSNpaz7n5dyhITq94rsk+BrAtwOxU
fx96KWFp4SaDbCS/fJHnejPHNzn5vaGuDiVKoFMftgaHGdO5plzEY8GA4OhQ
YS6uUozHm1FANde1V/+jWj3TFNAT3uEk17SR0MHYcatUZXPp24rb7kz1Teea
M5xQapPdbB8AuU0wwXrauoJlT8+5lXAVmOJk/XpZ5fE75Aqlbd2v0w+Hmp61
bR/2bLUtClKAgk8EdTtkZXFLTWGACvNpGMWROCyaQ2ZTGy0KDhreg6tjojJV
44tFckrYPcl4jJELVO1F6Z6DJ12J/puED88KOLVyMi2v5Y/EHe82xxyqISNl
y6O5S/s/jPsXQAewWnD9wjtMJL0xVdZOH6d09Uix6AyFGPmdWSjRxLd12U9K
ZxUO68Mh1FlOBYILz/tB9je7Vo9Hk+QhEiyuLASQDXEo35E3Wqf/gCgY5KcV
5EMcuZ9ByI6LYXIxs6r6KUfOFm6luTqAw4QcmIMCSzPbkWOLznq4V5UXgY+F
8GDZ9TE6CKCeheEeMonWVN1mP4GdN9jC2HqAfNUKJxSeuzve0+nmGY/Z1v0M
60tTltyNotOTPSi8myWxCUSgL2bJcNsqohOScSEXDb5aqlomgy5iCvDx+YnK
TdwWhWWLbGtrhTN7FPS8fMbom6/ng0WXu5VRXNLACWAcxOlefmbLAmQ9F0qp
T/oltjOt7u0tSNWmBEUBXXBiUVXBwWXSkvXT0AQSsB5qY9+KZ+vfTyGoU1s/
x+Z5UdLixHQt8WUC+yS/jSuw+2cnZiQHbzPD42qzkWMgxkPAJx5AsX2jo8s5
2HR906nrxQgjfXjOGKWDBeQG7bavV5WLwBpI0EsmZ42t4drgge9EHlSKnyUG
MLH0gqbzWe1VXAlCxivU9LYbMh6ziqwnaF+uSWICvZkobAfReO4LIfP35Fd7
XfSf1ix100q9WeWrUWJD5ajSDqBTXuycS7v7dt6yCva55jgz5wA6kRilfXsI
V2LYO5mWIz+xBMRvSOHO14gqsclRZHswpMtyAYcwltpsIni9P2DcHIXd1O+D
ehjXPt+B/uUI3fumD6KPo6THsZmLitZ95XoHz9mxHqb4IV1vV7rWtbtJ1FO/
UQeqh67BNzmJN9dN6furvPgU6JpYJ7pHi7wtIPExV3Eg3dKtOq7YfwlQw61V
ZtDOG7P5M9jYFvQ2iJQimJ5RbuxIFll1GMlcSGbLicpny3ldmrroQR8yJ6mn
B7j1bSlfgk6FfWfxhY12do2WN4gppykpx6M6kxgKaKXjb2xzDVPLKPL/z5hM
+yquWX+eqguOtAaHAOmdNXE1Ws51j2jdPKr/zHMYOBLOmoTGCWVjMQocJkZs
HxOg34qxfYH9JdhTegOBX5XnnEaF2m0jPCPowzkNy11h7gvJG8BeLC/2TKjx
UiXQh3DvzlKFhux+aRSCmDsvAr6UQICOT2gd50lm5vbUUzFJqJokAVW9dws6
YouFU5P/6PRy2bJ53/ApRUsWgbP295IWLX76yM4VYL6DOTPi4VKkwzkDcFBM
p7v1+r1/zWxRRhLkvCYGCuucBEILKDZRJM1tO6o6JF/2mXvLUWX/gGS/9czs
ojRpfBoO2CLLE6iQNjIJMcULyZB8QbZzrUg9RmyNv1pcP4iWCOBQ3ou8cgmA
Vq9gPSzaIAfDyD8jbWx3ikYw0aqk3Dpjl0Pq8b1w7hnk8+ZX+h3TkgEkaGLI
oOGAJJ9SXcSoli7q7tSg3Lcp+Udtnz55GO+3iGmTi415Aio7qT7/J9//n7rE
rPPXjd3GkZIxIgkIy/eiaJQoe9tIC3vcT3dShWs1ZccQXbRquweX4p+ZYmC4
RUzDMAaYTXPKql5ZuYbgkFQM4QNzMxqYhxj017eIo8RydfPTPr1Xz/VwN417
uxReIDGffr8EEdZCq2y01nxT8zAtlzaUbspEuFaj/vawzPwvS/16yuzkgQa9
sepbrag+ZKb2LqT1YJiELDrV2WOKW+8uDt1pJlEICxmL/gqzvdpxOs/FM43c
02cW1bOVpoUZrCWvOyAHhFqGrVGCgzLkXLIuM3p1ScEe1NmugQ3/Tj63UiNg
cA3oL7HYWOUk7CA5Kc0kWVuC3yXEWlOlS3vjz4qbxPB5zZAYaUtxyMa94xVC
k1/3VoL3GSrc36P2nJ04nHp1GFBQ9j9yTzfCLDHhFELfD42Z8hdPjYf3Lua4
Qm3MesIZaPA05P/JkWEtlR3skQQ681wH8el5l4cWxGIKWxvlZBj5fpCg9wYJ
TNp9SmscNd6rd6oSSQ5aga/Oi/SwNWaQZYxHpS+lCiaWxst+vv3dbLOq5HHJ
0IaF7BiKPaDSoLd6pGe+YWy4EkCGnPujbjfRNfbEmvysDfUqgteCNndWKJSK
mIih8cjuwZbasnKzjXZRHvlittD/2YL4CU+breZ+FvTT3Q7QLO+Kw5UIA5ZX
uxSPEawk4ajfalAW4a+9m/xB+4N1a2/yF16pY6Qqmvu7GkctCUgE6LG89IuP
a5rROLX11kixXVOvhiunbBxQCf7AFRSLs1ZUJdOP9CiTpZt5sKP2ahpkEJtv
977pv+H9IPjHhkLbhx4KL6loZmGE5f1e5BV9G2CN0lwvybg2o2C7mkLudtNW
9PV03WFTq/Ydu4S9FTuylQiC0O7miKee9GDNuT5lizIlZ4x6db6ryS5R83Ea
K3GH7sUvVk0dkcekT1qK9anupdg8chktyQn+HcvnMZv22S9s9aAn1evjdAtf
IQHJviixGkbeOJturVi6NiO4Xwlx57jRSI1pt+I+jfnXOJF0hbfHN16cNsex
EmOughl6NBeGTJQ+U9WyVqQkdbl5VGz4sSrM4oEO+ULGIuF+3qSelIojTmwd
pHCL2eJhyD54RKFSkU/MobpalbdBAgELgqU3JWksLjoE7UothFzBLkcQTVnX
S09qxXeuQwxJOFaLwAhJ2A85FjXxqgm8u0cCMDrYXnfzzwHptmKm58Ah+PdF
E/mEY976q2eaKNCWA4ddzhQXsgEGR+DiUHC9D1hGkAsy8zqfSniz95xL7Kyb
33xeb8qo12gA3G5Trloq1tFPpQmOJKSMvnP7Dts2LiZO9jxOO9xN7kAkT5Ir
iFG+5CENZjK6KRunE3UqdyAh6t4y6wPDAgtPhlnyJNAP+Mvt5lhN8MLlgPac
mUSWyelik8CPrwynDL2uahT5dPBnC+bH7ri1I1VfCEvEXM7RkOUX++gDgygw
IT0UVOMilCwy61j8t3FfZZpTvTSBmkotggxn6exTNVdVckMDaHXOD/FUsA+c
O2VKPn8lXrtMQthL7My6WRRXKzD3a54pGIqZTJwhp+Tqhks+6QC5sNcjD3X9
E0BbQ3NUN9lHjM4s8fuXxm7Uvn+extfFbUFkVkadkDM6Gk4UhBSNBN40TDjM
TloTteMEzV1deg9UidTVT5vurhs4W+u2h1HoSyj6Qpew2yuDolzR8FM08bT+
Lu+uoqxmOHWfdXjuqyfy90L4uf0jdGvwmdoMb7mx4AOJ31r2fzL/5pdg2Is/
0gAci9KYo/m8LNn67rsKXYaHQv8MLIkjBs3KYcHyoqtUkc+JWio5n+cTCCAg
wWhixgquL9Jq20fNfO5YZxohl9UY1uf2ngfOev1pJoAbB2EzcHEaGvGwYnBu
Ok6yrprh3iOmYTafU/iFxabPGkurpeAVXSCVRbmheOV4MlZVjfN2xi25HLEq
Jdt3st/PsCRBq2PXvzKBWxV/k76U57rvD9o016Gs7U6CmitWUVAVyi/mrAOo
ym5rxq3Da7oD3yBnMU0qpsl4CpMz/S5b0MjRc1RyieSEMxCpIlbX4pNAhgj0
etifT9j4wJjXLZJ+k7TXyHBcysdpaWbIVWTjG6yriDJh35COir8W+6iOU+8E
1l/V8quXiErvbZ9EfwjxvxIbkVwd4bdVaItA9xG7LeNRa7+KA+CD6gOtZ0Ji
cJsu7G9Uab+4GNbql3iLlpbwc/VjL753S1OpDFHg+iTIA/KyY8C6vq+bBWzF
mF3h4awEshtnoYxQZwzVHfpS5C1CrE0LKfr8uqJKu8XYhLjDYq4IYu8IVcbx
hkOokQM4ZhnLMVxnYe/RiYlkqJyKWOZ/QkCBY3vfXBYiHca+IR87BMAtWUKL
P/bDEhGTUL9LNEe4KueV/N0cuZi/D49Br7p5MDZIPE7uPvRB9vTxdheYXKoV
R+L6/sJYwi/ywbQfwYCtPSxKCBE2ik7lB5VVWdRDNRozRRiilFA9jPa/+J09
hzI+RQD9n/F/vW1X776Dw308yD/OnsQGLcfCkQusXQp6hgWZD+DyzvE/Smd7
iBPlbe4UGBTPJt6bkBHrQvwNmKz3IssIwmCe+jJvZibmNyfw3AlG7nAh53dE
DlGY8bw3p3WEe18owUjoExpq3cPuzxQYXsUDNgxLlPvctTla6cus2LHX4TA8
sXCdLcSMqOH4H+eHrMnJzFRCkl0RACC9FoQfRo7ch3OLwVLEa+rSQl19tyXj
7SqjxTAf+P/2h2wVAz422BHluII1c2JaFBTpDMfspLBdhnGfQitbMUz3SC3F
B5XEEx+n7xQKaExVpUAmj4030L+Bn/QOwfBoYzhDHvXQmwyvK6s0zOeSSQNw
Ylpu1ufBmkRjwYMBJunyrcECjsN5Dl0k9ziiyBkqQvBRbGPsCDCQqMA04NX1
Wit6MlEyOmq1KhESnwQl9RM2VAT9JMbaGZqzac/XZOxNWdenkxC89UWy4zLF
udQiXc5s+cQK8vbnDVMC+BypdotVW/eApOg5c8scGiDF5dvzmG6V6OWJvq5F
YnKQCJx0tzY9nQcsnNKA2kJSIKKNJ2l39YnZJ5++hYONBOkUjtL57eIxtgzn
4tK1SXswLNQtZk02b0J9WRCxF5nowC+50INRosrVswJjYWwDNlytGAdmEJtl
hnTGsonN1UVp8E+9HKFlkxp4TWgJq0yqC4Vmsd8GwTIpwiuI11CR/T9ApFeR
Th+gf7BjHb5NaqNBV10TS6sENyHgI4C0H5cHDDtluDt60LUtsyNnLLV7vMQI
xZ8/SpRsgNYdehLzHgLlCcTYBH9gAB9hxwUNKPO1xwH7ufmJRlFVEym2Poi7
ao48pe+11YA14rRYJu3qvdDBHDUAGU/tcHP/u2d2sL9NNRKeLZRXictCTfpz
Lt6/vP4+c2iBU+EAt0XkVQc+6DhSz42bcmZdVoZzAMurast7zom928ZNM+Dw
0sATdxIEeyBt7s9LgJtzYbxlTFFZkP6SAJjy9yfmVffvDXo41+VKu8uZMZj3
dWmvKOC/spB4FJCX0KQyZft0cCxvU2DyUBRhzwoiz07kTeYcxYyiuC5BnhUj
kwuQMrE5UNnZOAUMPGy8m7V9Oahsk/hmBkfmkNYZDYAZcOnZX4x1JIHaodix
hnJqeeshNJNNEXmIdXBqqjSdZIf3knvkX5TawFM0DwZneLBvbJf+SIRtsvBq
6i6shIXIj2OO7O6I7xj779ik4wiIlEtLCo7y4HXtsJXMOm0FUeVWeRLFz59E
+cEA79BdIRuAmJe08sY2u2skf7tKiHcXW/rgCjXNG+4ezxcbbd+pMI9lnxhw
Zm3fO1EHMZHitB0owIXQS2JHYF+eAQpTtTM67uDAvy6uI8kxMkBpP8H2WIXx
HhjznJGAy3gNBLYuDdyTREbPFEkWz6d5eiOll9gFGLI2j2W/daJHx5BjYUTa
RR0uWLYCk+9xvDF/cnMzmThJMgiRHkxLLw+PVAyC+/D61beo4TtBfZHwas+9
GvJohiFZ6UMW+YgEHvm9la29uTS8ZHbyXHfnCtFNat+qYMlguTZUqMDEZc2s
9+vLJ8GpzSFa2Az8+k5ajiRVZgPDQm0MiEr+7oWbSYiIJY6Bd/JprkhgYOCP
/wME7NjQCKtz2244SUV/Nyhp8pMk+wtyZToQyOWFgcLBmH9fwprEyT59g8gz
phokPLK2LrgGzbqwizxac6bngOY6JrUYXHD9cP+Os5w8xjAe1e9q9h2vQrzz
3/FUZsg075rPEeg27lAd9xFv6htGNR86To8TLeACa8xwYw3SGry4ksyTGb15
+K2AHA74jxth7FALo9DTq4TYpLLADLZF+A62Orw2Zv2GbIjdiE+Ckrhl6r54
7byen+lM2GYbK3kKvoYsn1viam5NVu8aMVGixTDKaROqvgs1kee6P1HxFuG1
dgtkoYzdfoqaiqpENdKHGTsPaUxUwOoehgpvgcQ3IsmSpqwBNhFi8tpq0Fgc
tgv4ltY1ukmmkRRM++DgzXmHogTE6Iemlyc4HiHQIqzzG6wm6X8WLHUc1I54
3JIJBtrPNnXF0/KG2dYPARIMOnQVtQwEAtrbmZIo2ZzE8bW0wfK/824WCENe
Z4cNIwaoLHBfAH0OIQBXC/zCrHtGl0W3QrHQX2ktTlOoHBP3fCEo5fCs8P00
ixxyQ3Kqhq4H5zFx4e5gM9BH/gAsUBosfLUTfLkkvAbUwqaO/ulrAjmO8B+C
fH1fb/t/nxqZPF02ryBHsCClHtYlCMgEaKrBhiRT7L4sp4XnvmQZYnyU1+ib
MJPetWd33gEES5yxsUgDoBQFxQIvTwO5aikBCboNfP5KZQbZxHYAOmiytZ8F
Q3e9UTzeyZFHrgWBZnct6YX4FtAjAEozvIF9WqfDDso/28R8kqfWUerD+iyl
gNNWUHnDiXvFpHIL6KJT+3GuKznl3U0iEIZLwQO+s9yyMAxstJKxoMhrVXmv
lE0dvVjIt9f+mvN/vS1P+qeRDtupQM6Zr43HOIZiZAJE8noxrYRw34+XtgYA
OwMCzTWjv4uU0uyU977xgpWG0+W5WTSWg5OdQEKuQtdMktM/4n9VHk8yH4TT
4Jf/Mm6oRGvPNfr8mcsXqalJLi+tIN/ed+hyvXbWrnGiPqAqCwsIIUuokESE
ODSyICGcES9w4YnIqGLVfX7R6T7RJ4qqThEtTr+/bM0Jpj+JyVEjpyJ8IUc+
09R18vs40oWtRSFywGJDAhewvjjliivVLbxzyzcXHsLvft37YQ7Ja+HHwA9q
R/wHi8FYLbd95r26zIEEGxDFGnvQbDi/S44EDTzmYjtQZGWv6+Dz68c5UT6D
yQOAQ1q+Ixo6RE2l/NPqk0NxvKQs7SfK1k1o5xvflw4N3ALYcYAMHTDqwK/Q
RFvSjer44Tuec5Cu0rjHDaaVfdOcMYHyDSN/CnZMK0ww1LTxE30j2hRRLe3W
qIIYoqk0FawveJvUynGPH13Jl6orKBvkK1RJZBdRJcHc+s8qLWF4eM2mWb5V
ixcFGyeo3d8KzPKw1AAYC/9XdMSP5sU/xIGg0uJCZm7ppPaAmb8QnaF3B5ed
9qs50+CK4Vcck0P3rNX4SExRGWKt2pZ1bW2z6MKKfVTmmetxMRWAUbUJPvmE
t6P0Q37ZYuawkesph+RgJCOX2aQYAJEmdMuFFtR51Fx8fQqXuBEHMVsOq4u/
pLDSx+3hHBNW80ubKqJg3+qYR/RH+pp19FBtto4s/hYQkxAiZaqA4THAxTta
x/1bgU3dMg9JMS4oD6RHJbUJly73GBBK8qGNYXGHQJyRdWoflq9xpwqcz62X
sT4Via2L2N85XN/SQBsBTSAL+Vti1oCKTDHEvqPmmURKMctatjqmLEUx2Fsd
EoFglnK43TH9P1hheIC7FCGaEkpXEsrngmefViWtYXK7VfyZIWMSYdEkJ+pT
bavmfRE/BYX7YfYNjCmkcaZlfUZ4haGF6XLRRis4w1hRDQLJY0uCZTgsLR1P
bfEeQ+DdzzUdISeys8/59TRx9mEB08MQ+94zMOhuZDLlIVXk53/hqDSQURnm
dXwHIQhhNnL6bGbl8E37SeElDGaOb/Uusy85kLdfYP3ytrGFS56cYg3DCBUc
NzeYvcv7m15yvVpGAvFSscbjbxkBNttY0fUNTqXmvC7ldbdlfjHspeg4fOfd
XdMWP59mpM7rwoLnNvoVKxAKL8I1tXV+cP3QYyeJcyhGqxXh1dsJkAOz7pFQ
am9REq53q/bjmGXrshyNFkdjbm+0oc7JFLunfqd2Nm+BaSlzn0guKL3PCnNr
fddwgADHOUKWXApnbZ1l1NG5pKev82zKG+B5mmsazygx401AxkhXQQ15DhVD
lm2+wLGdJ+cvX1z1i88KFJavOn7IJghNCKG9Jc/vVXNR9qS5rrWstHMbX55z
CGT/X5RmL9zpRXGtV+tLKe7g+Qz+sOzvxTu7b+yFax+aF1CrsB0ns+YMOapJ
DQtQraHaSJmO52TzlyAhNWVbczY+LRMpruAPxF01wCZGfzhw+4sOR3keTunk
M2AXgDjAasXf4jlwhGY75X9kNOWLxnBmDAB9Uo70HiDjp8qyZbtQtjLDCN8T
QDaEvJDBT2IqmN2RFDUGcdK7oASSbCgA2H3p98iEnLizhVYwDUdn2NOcxIgs
lxrK3LGT7OtrCyohDa1oXEFZgK9j72RyXRwDpNQpfPtj3u4Js1iBxcMdFiTn
UivlwdHjyGv96Q3V+NOTkwyZoX3TkytY748wvU24JC1STqaFV5DX4cvALKUP
tIl1O03ySVFJZf1u7D2UptxRnCRbMQIen90xHaDBxloaCIph9VZyjJwgBt4V
H+IZvhmavfkhPOWCVQ5iduvVtUObixqs6l9hEeNoESFYIICW/PxBy9Lbf0sl
DuBxwrQ66dYhaVCwOpxgobervasVyz/hEAltUbGbB1EXvsVzeVYfO8+P1CoU
PmwWnZbO/2P9yx57iS+78RyPPW1VEfm6iN74sPV3qziTSU051MrFHYvBOZtm
Emq9kn1Y3YHltubjWNRQI0NNRX0yzCRag5AqoNWFxUVGIWyTe6OVfrB2tdTD
Z7mMP0d3Ii3CG1ntSCjEtBikY8lIPKIWRddkA2tXcVu3bsFUhM7QI0YYptx+
Lwe5EtM6ANYnlRQJCqWkerdKrUbgTT6A9YKtkj2Do8xLhs7kXcFwApxsoCGk
rn2EjZkZJEfQ5MK71KCevKqLl+z0+ZDBQNMWsAGq+hnEPOLo/trI/YjvY/ua
KtP+MTY5fWd5bT/+W17NfNLC465P7CI5K1bOkgsOLHmVN/j1yA/5NKoQazyL
JPjknIfHmVT5l+oqKloWcLvboZPlHquPH2mWZG2X1URqAiQnV1Yw/tDZM688
e0mipR9GLM5/5BrNpc16hrKEssz75P2eTlf0BEN/DVnyHYk2G+mCmc6gzPPW
ti89z2cYWS1gzkqiei4ep2CApxxU6gkzvLu7Ac/JknAn436iJj5NtsxjUW/4
Tdon1QdUtRRXkk/B38kxU4jlfUM05F6PR/9BKR7NnqdtEgLIwMt73vA1Q2ks
XI9EVFVcZmuOqBHLkyDNimo0N2l10bjNSQyfa76WJcTfgIndT546nVJiDfNj
CeAGTWBAo8dRF0yCIaMRpzieEnSEY8Sp1f1ND4QbAVWwW3T61jD+fykACYNa
H9DUHBRpALp9oC96A18M6csncdk6tWqDSOPbwJoBIdiUtU1DM6lKnbVBeFXV
SP1wZrzNNafheI2mdGBiTFy2gP9K4xT348p9u3yb18EzL8HVA1+oiGESfE6E
rrhx0xsmr/pG8qdN8dTU720Lod2s3+C6lnaJmLD7nyaH0GXHOEbJZZinQbZx
vLDXZlhiN/oIkgU41RdKFDrs/X27MDDqoNsjO5WuNIryYA1YNo9HMkrtgpgD
j+XuJln/Rb2HH1weCtQ3rWDpW9Do1+P8i/KSwWMZiCoUsaDl8uCg0u4q8MKj
+xhBaAqGIRZBBg69uHmFewNkXR0v73t6tZC3SacfSqq2MwpMthykxH/hqx+G
xLPsORKCx+DkOwSeibAIY/DAcTdts9dVSyH4eMuDIenJaYAHhiXLgAfa1EHo
xj1kHCRLe1x1lhwvQDuY7ANvlNBXFaR9EKNDZzlRaO+HZJj2R4wH4Y6KeD/H
/jkn0IZ0IywQ5pTngVdfSNe4Q8inbYOJnIAC/Qm/QyJGGLa4hjDR4zHbJfZT
31Hm3ZJcAShrS1qL5lD7CyRW2Wuh28bZyQY+v5Tf3Hjztm/Kpk84ywigGiTN
pSVpscigiMG/yTHwrtdERooUZbDbiULiR77nfI4RAtohCp/5sBHbzuL+YqqZ
Bgc2ZLuMbt+1iw8kSBPGXZXFxcfMTvg19uXHo7VSROVFj0UoHVrabpOud3Xr
p4sUk3UzvMa1DMX7p5J1vCeGnbZOAzhOSZH2FO4DUP2PyAGBVGL/zKTvVzsS
d1U3o+m6ZHdBHb4Za2CFtPZt43wA4baRBL35prUueHaVG1bcMoNWqVrWMY+q
2lPozZKpTxWsfc0F1VpqioVnIxLR8xJUs9JVpS1GHe07npvOtsQjxH/RECz2
EI08rl0coLpL6E8NrHPMnq51wPOlw/2ZqtOqp7SC/94E+k1fGTu4ZYb/tZ/u
ZDaZVvEU+Qg/LD2dNfWMSMSR6qF0WG9gBJQDEk1SQRa6zFIY0pmNSqsPq+nQ
XwFKlatXbV9VkozkHZcDs//O9aZo/+7T51NzCjpipBPHDam3F1pYYCF2Yvww
OLGYcSteJHKTaPV9/EvyPPS+e4wdESNiPQ1OxGz8caKtdvtqmefS62NZKa6w
sppQAcaCUNuJvbIBgoovJG7oiwc/qH+nvm2b4lQKwLoJm1zo3DLlNia0Jy/7
X06vlST1i08jd8DqvzNwwH7PCvTiLCxQ0B8SAY3exvxHEe7XyJozfE61sYXG
vH6LLu7Ejx4h0oukKH4l5863fyPXYCQKZAs6NxIVfWfd6pkArNM6DXkER1rl
ycMxjf5ipvBFxQmybBcKWiuV78HAEO7EsNGFZqJ8XzxjljdCYbb1Ymt3nmD8
aInLkcSY+2/BXY1RE5tHekxFTqsq0KhSRL1v8AVSPyHB/VyItexl/e1xwoZ8
6mbzeQR34UeY8nXqeo3LziOgbGP82udQahHm3AhZBxU0Emh0pFOw9EI49td3
WPH01DkwCfHC9g4yEJh12meFCdgeWK7ZpATKJf/JNRX3937EC07wzbIa2Et+
zQGxRJ5c+tjtu9j3xBfP3ykXjFko68AMvymtcW3v1V5g3HXPzqJtiQNGe0XI
fp5TbbpPjgjA8zrto1ObpYFrpgdbwh5i/Ci/za0XMWdAUQAd9IwesGkzb0J2
S0enl9oEVcHjDjRwOqTZN3vE7CaWe2A9Y8F7vag2MOQko9QcuqEZ6ZmxGZdn
eXTYUGr68/keYRbaJaTx6G+nGp0rWoIT0eS0/GtIH9/FE9U9cU6nRafrq3/p
/i6555bmYraiXmjue72aSAVlD0rwaXxywyKn4vX+uWnC1fjv1EUmnXzCraYh
Ec5uRXMgQZSV3qbM19R7OT2F5aJyslz/lxNbw3cmiVtLxhYUw9wLNrKrDCox
OCjL8obZXjqs8fVxSncYAc6KZZtQQ6Ep15lcnUxdQ4vsFKY7GFpF9qQXWfYF
SufTzIcEz80kMO5ouZ7MVavR97Mc8mkw+tz7P1M4h2P6IpRf47qRjPPHQSVB
R9jDuPSRP8/nVTba3shEYDrMBNY/JZokFqWeOIFnlKDcRffv2ywubUAZdjkF
iDIDWg83qK7FT7Wwle6c3EN8IfoeesZVUefKTZKMlJXzu9gXI+UDHEQ0/Yc7
m6FILNcF45piMWRK1mSUHJnvEl+riAGaFlINcfpPKA4bQS5zkq/Bfv5cb05i
MxOR7XhRmarQQPIMDy4lQP4JbeZr83iQMSJVhnBqKKPl1zknTLxwx1eSv0jP
9Wpt4MzJVAmW3kbtwuoV2cw2ahePxS0EWzr3aZJehhdepQOCyni8lASEA+CF
tduYtYcLYgycXbvvRclXzfhVvey/d0hYDT34ryH6AnY04oz6Nn1X5OXJIgEW
0Y9g/EJ0C+gE0YwRJpXGbwTPdNhnboPL2SYzGNjXIlZdSka66ylO3oUgzgrU
OVUr3MY61tODhsudLtAWOOFOPX0JQLy9cTUgMaezsFYr22OolTWVznytigG0
hShu1twJ3yU0jOyLAo/OiGdoZv6f/4sf3+8PPh4ECNMFczRJKwPrQ//pjrGm
rzpCSwp0dnGikoDDg2H/pWO2jgO92nxRybb4adR4YE460lw8lR3iKv9V9YOE
9Ta8zGoqCL4m6AsKRkfhfoRh7kvcLtno1se4sc4VyLIsjezZ75y9X5CoVNrj
xYz3MHhuiDBaBNkmk5FcEzYU0xo1l0AsELlDK3UPfG8uYh6V3mUn2JFEKXjX
SYtpp4Y2QJYbWQWwJHZHwFWgP4h/ysAuQgArr7NvAucWd7GcVGhB74dYJezm
YA5I8vdcnglOBwu4TkSIdN5eqt4PFF7k3gIcQQpJ6rzc1+D8brbtsP3Neqc+
v/2s2m7lVflvpU0Wd9pETkfXPgPeNEXnRRROvCvcf0d9B02/IMSt7Ix5WWu5
VN0Ep1GsmtTCQpP7SL9x/Q3qdU9Gs1hFCYlS4W+DGqznHugm/x4Uab/5GkjR
s2kBM37jDDeEM0WbpNY2mi1CS6i6czfwj5i/LBlIJ50FJCEk4r70uaXU2uMw
OiFy32+1Bm1rSOVu+4mRtz+0HM8xLVQKnUodrR0ogMsTwKSXpNyrUA+ro9Xs
nfbjDy9g2QBzjRXgEpGnLQWx2vJHlq9Xs214+8gvvXn9XrIwQPPZwTMTgvS8
wjOTJ6rnSeL5P29/HFnD0OceZjenWFuyl2JX0NEyd5VeWmnsmPZXxaq5GEWI
SWrFr6+e343aQ2ZkzJ9r/BUypNDCJSycR4d5JrFRp+k6lHtkcn0fl44aSfgz
7MOVlRsnaUHjvInfVTDTU+Ywfcxx6yreeD1WreAK1kQt0UoOAPIh9OYIPtX8
E82s2ccH63BXohfV+hTja4WocXIGZEpOhBeExVwvb/1uohPlwfEe9WXzjgLW
bZg4OHSDsqt247/Jinem9GpkXavslHEc2Cm7P6YNs9O+uAmTEgBPDVBrOMN2
VsCkEn92bpRYXIZG6UVupKpa52mkOLC5PA/BpxklZmZI+m08g7nsCWZrEAK9
tCXMwEPa15YhRzmoKldwbYf2CVPVcPTt5DmSGMVHGdcfsFpM5Saie15sxEzv
409lj/4pgmReNQgSKbmcnXHzLwGM5/xfDYHRMI90ab5OhBH2tNdNGLxsAIla
xBep+2tdT9mNjBwU612Z2BoIEHioxzg2gEV9aMAPZT0MGA2iWkr5mW3IwFFE
wt/xl+Md+eBS4RIBBlD7sgzJBGkpmSraVWibRPKkyYFz5/QgSQw3BDEQzzxZ
hnVUA3oGp/+oultIvZmGbDCc1QKFcYKnqAbq3vARJ1FlOJM6lhDJZp1kEsRe
6KaySLCzTyy0ZVAXlkVVmjBtSKHPGL3W9ZVfeCn+oreuSCJ0VxsNy1vZnVHt
QmmP/HE1yxs5rILzSRFMFD5BqeKQG3RX8Q9L+opG7BUCHZvq9GfYp5GGwwIX
iWF/BwGfZiVxFLdZYXthgRww+0OO4XWtW1oxfLz4bpdwxa2nK8XWbbtX2aIJ
V6yeK06xw5oHe+r0DbsJp32rmwMdQ0iTdCjUEIxzJYKayBUaR1/ct2Cv7A6D
121I+aEWmIiSJSkFRR9oQtFG0JNAkar772B8GvRoGJqWM/2on40nrDuzTO9i
UHhbDvgP7Ytz+pom1tdfGowvOa/vNeE07nQ2cHGH9yc+5FJXRvG2ZTkJ766O
K+qLV+6/dcHxVrVPFLSQfSmLqAj+6a5tg//DF8Rg8zrp64w0f2O3VUkWzHcb
0GjqJDzqfAWNxQlB9bfCbkZUCDgccUw4sD7R2b8aP5gCADhMyt1tmblWv0bV
l7Fm3rtEyEGO/nIhs/X6w6bcevpiqo8DwI6d9Gd8+9W1NzvYvZwW2JCs6+XS
fb2tfBdyZDcpkvQ9G9+JvO2qsvm9tWypz2lGx0q7UeL6ZHT46EvOrLJ9KxIV
rgn7+EyTc4NQllUJMfnJYYQ65kblFsTXsKowarYmd0lHaJX0WIgM3rUFZk0F
wiWpte5u4rHMrUTtsI2xhRhymQBvglRwnwyQmIu5ykwwgibactLH3bMPZZ4Y
pnkg09m0qagrFs6+Jh7Xf+HFwMAj6lih7auoG7alJ4c7ttB8yUZSuV/ExH+t
sSMxkudV2HHKoLfn/5gP1kCwi/CtJy4fCoVU4dVBJlG/9OZi5t22Y8+oKcS6
UQZxkI43CS7rv7v04hyXrlRl1nkoVG8I2xMVHNo/DGk3GYUugIja/b9hjDlY
K9cZdZSC8Vdj17vtV2OLNbmR+GQId4lQfqV//whvxs5mVwpaaCcY1Ht7LQKn
OWFR4ItOtFJX693bYGrDLYuW/XxUcbw9yuWYHPoo1IS9UYBiwBvhbpl70qv5
x0UvukPkAxqGL4+sTwfQAz9h8QHJpuGDfl2Epe6kGYUvQ9JwlCylUfmNVMdb
KcsipTek34oFgJnUvHq4lVuGS6JwhzghOOz2JIgG7jwU8uEkKOH3/RE9yGJA
YEQ3wl9dIPxXv2HODbxOwI+nt2L8leIfGnh0GH4VVP1Cz7CpDqSXgmheuuD/
i0tNKmJNd1X5qo0Hx70AhM9MIzS8OuxOjYa4CSqix0c4BJlcV0wga3R32IIJ
HyAMjDqkQ/D6hIlp7Uiw6hRjwdiDUANC43X0MbhGgmS55vqlOxFgDbMvJYyD
9GThoRbS4EDcqOnmYt4BpHVhs29rFE/eJcbaElRTk0Drl9MthoysTeQmmQHu
2bLXeXWBBfWf/O54maJmA9JXXEW1W0wRajjthRftc8oSJffdTcy2udru3QpM
hlHRZ4eQKTB+wd7DXkxXfWnmIOlRoz7iphJhEl4t5nzPtWBnj/tMqClVsH2u
iwuBYJ5glOVhnu6wIoj0tzb+iuwSe1L6fZ3szK9Gwu3eGVHpb2PkytBzsqKI
r077PQCYEkQDgBwsa+ct/KvdDk5dtX2pZoFAbyVS4LMp/6PL/0i2hYGxMgbg
NpsTS9jNMPUcHElU83VZAcdZOiQRo7s6hrwmLaJDm/0ILN2EHShxz0AYgFje
fum6hSX4vVKUgaAbWH2zGclJTSgiaRDcv2m8lRnTy3fZdea6MEM5F55/v9VX
msD6Hd6qGZdNu60TkzKdZ9G3gDf5f4QOsnzwRzPomSatLJ8ClYEkqky6YHVm
xvuw+Pt5yKrWCU6wzw3dNA5/QtS5SkUQH1+kq2SnUqQ3CcVlQ0D4eZ7ZVC4j
gK3BMYLRN+TNjYPyq2/oZiNSr/GBTVMKO5FTQw6THYPynJCDK3JaS5/Eul/P
xY3FDQGrdoTpydM54S6dwjgh0Eox2+juD4DH0qSo/BxdBIPfNX8qRkT7zFuB
rFrlxTJbOPOa2EwkFJHHMZ7KBkGzZ+DSku6QTkwVB7tMxNaJF704lLnCMvlJ
ivsCrq6OZierHJZ4VXyHuW7ZADAaD8hBKYDxom0+d7nIaLQhHYXwexjF5SHZ
T0OZViR+3VFcTO5Zz6/zQyN9p9ojXNk1721ldTps8GgTEGZNpSafNJocasH3
NQ8RqUfwoPeN1jYX5HLTKf+O9Z3f944WFHO/gMD/bkI3Ur/57tPADFqkHStS
P3QEcn8EO2/KrUe9XIVTf1CR5/PUdPGbjaaHOIyEwFJIr9qPthpTtrtx+Iis
/5bmz+XtqRUuNOIkcit+i+ZVgWEDpJbPlw040133B4g+o3DiZuAshFltBNbc
nDSsaYs0XbgD2z8DcT8ZpNe7HelCebusaxKN1KVx7edR830Oc5I+5RwMdV2H
1hUo+uC+xjRFEjF5ihIKoHH1RDVNCw9X9e1zW0ogaJgNUGHr/uiUHxIkZZ5o
33r4ZciHOyTUzVmATKfZoPXfpgIhm5RtxnohP+KT/me9E/kjquWXeDSqULWl
+ASS85WOrBEEQ0ei+OZDgFP/Ab5ux8TeilM2G7wPS7fLKIag/0REdr2AN6ce
mNW7sY5qXMvhHQQdHtEkyJBDGaFOCBtvo1RLwTntD025bvYdmITbSQZbko7Y
bd/2mT4KvSf6J2FpVhnnGWfixktO4LGEHwHHa9rACX5k1JONVhZf4428tMyJ
TFaWzuWiBlsJKyBpo9Vqyne43DTSYNWmrJoHBtkgaR4R17dG5BcQQPyQD5so
eEEKXeGm7ndLhDBClLNZkCiyT0Li4ot/gqY7siVb7vdYFmzQ1UgLdwnFqW6C
rV6WBQ2360FJ7DmLvTRlIvM+zA0MN0tsgyB+XFzjDSrwNEmbdSemZVW8T4SW
uCxxDBfGFqwFSbCYV7VfSVt3NkzMEC6ti/8wqNPTFqdi6f8/nCz4fLzTCiVh
pMUjkGVDJT9BOXfafggThH/AypwxOWFXNqimZhKr3hwMEi5+bbmgUggw/Jyr
UEo1Rk2wmwyFpandxHlkbTcutsxG3gT8qApLnFdioNVPiRQTuIFp3+5O4HK2
UrG5tpCDcVYscXZiHIPNBGyzoQH+TH75e/UQvT39wAZ6LxbQA54R4lCO0JiD
o/mfL+Hphb8IZCVNsbF97uF6R3UBgANYR5UhuB3otkncFb/aoCOxXe00S2Jt
ul3a0Yh/VKhV1BDx6VwS7AkZ/J8VJGSCjwmCQDJh2MtByVzwalVkZ794cD+N
/rkgSKVSI6nQ/nxvTbdRCuyGVJ9mJ9vYG/V8J5qhi8xdLPFk/BMDF/j/bv6P
k4v/TFEIAjtiOD4CMXDF4azpT4zXI6yxu9BoE5WMaskBxMqAtIjWzTuTVory
DQ7clfqx8r+NLO9U2P00Jq+uKwaAkBH0J3fnXlVLnRJvwSmvgB8blOvcVWq2
44tgWt94yk/VYsGETIYWoFw1otiHARsaKE9WcjYB4LEji6xwWAPMU2tFKsaG
JGQNaQZ+CPPJVQJAChNcMP7fL4PKaiky8cniPRVAoHRo7a6jV59U5J7yUWLh
1cSvrT94m9DltmPqRH7/SbBBCjKVzXQpjfHbOL3WWAOPIv2tOjqbXZMjmytc
VJmw1AZiBXszEzqPhV0nGbetuPh9TsR8kOY748NqbUTnQYrm5iSSUMVSVG/w
tTlqH1AiAyhCmSim7hCLuAK53tGmKdyFd4RCYy83bEsaUUa2gWAISo613rGT
1zDGfY2Dn7lvHjxcMLv46jh/uEtxJOM+ypReAk8eF4aHbf6nQKO/rvvJVjKg
TOWyu0GPwfkiEFWks80A5BaUQU4L2Cr9vlLFxixezLQlVGPawigg8xShx5ex
ibQKLwrlnEgnGLpx5GFs2HVZrNkZOfQVaAY7ZSzof3NbA0B15nmTT5TRQPu8
/8tG6TXjrZ8BDBRr+Lb8QnHt9dS5uRPO7+P01/9aymSzS1XOqHzUg3M391KW
TV0Tq6In9MikzMFgmYrHTnUSqaqMiE8OY08GLCwb7656EOID1+uP0hu2nUm7
6Ga8NRtZnSrHO/peU2szqWFYcVq+ILZtlTfPPE0Qrh2R2RQpNV0Q8ZfrZc5n
Hh09wdEgcJNgcLxdkDNAAQvXu7QpEVuOhrWulbVhuKSFWFiz8DPiAjInRHW1
y7HZTP/tNigSYpod4bp96AVxO6ivibMadNOozzuPp25mpCjSIzVUhxjE7EKu
QApNAEMS2zeZnkWDk9gCD0UuP+pUiD4BXyY23ckswJ2kXM10zBAmzNHAYGrE
Hpllqh7HQOG5U+9Tqcv8HzGq2xgkh/+y0yAZOPMNuxRgkiU9fnYtCN1eoLeO
TQ1GVQlhmi1HBmjqLLL8Xp0YFGHH8TNpmKS0Z2VBoNtVlXSrIS5ruDEH/K+O
dcDxQ4sezbPW8weKXFhB6j0Jmv7lOnnsRpXqvXNZCWoaejMriAqNZJLDMzBw
wGrusYYtUK1zTM6tGS1CWGQ8sg7Uj42RRLhUQtjWLsZgLqPoc6NfPJ6sWXtO
IBasr1+c+RLU5SIB3/rVmJmVCA6dGxpa7AUeYr+/b2MZR1j4vSFkKmRDd1Z0
hFwWv9p8GUV4W1cqm41nHIsZxSg1+cU9NGEIS09JoWwxCo8P/cHZ0vJIB142
reeW+Mx8I42F4e/njZZ6bfzq9khFIrDmZKjY6uhgYDEKcbIrrYbdOvZjOnyK
QW7X2lZOdR4x/pv7FqUrCPIJAKetLEshqm0eND/7MhMyFSGmCD61v8q9nsmX
gYVqK/wbjSvd8gRevXCh7IgXztOwbAGNcy9OUz7iFGsl36yAWVjaN5lTJmbk
+bH5ywB5gcBkw4ZNNBffFw5NZPXx4vUXf5YDNZ8BIKDAXL9BYduTB0gfX3x8
K/mLxYtjkEKgDqWvBXwoc1xCDn7JSakCyOo1WKn0kONr9cQkykZZ8Ba7fBCQ
NZNnpUDpf41n9hBvMW9WsuR8TOhVYsoG8D+aBMvgQ2htPx+8r+jJLM4mUMXy
1XpQjQl/CCmiu4Fjx9KMxkgFsS6Az+/jDwXQh5mMvGHccWSVgJBpDXtTVD8Z
M7QsE/mJgVdoUD2hollU4qneG0wDCBI9gGUoQUnmLIZJ07JYA4eufYhDsKqH
CMrTSTD/QbELIoSaMZ2b7orj0wBVPiVGdGgvBTTRldqqQZUNM+LuapazhhZm
2sNaELwCorK0On5WkssLyzxRVj52usPGnDL5H6C+Qcs2Rvvbj/AmbjwFJzZg
rSIHl0FeNm3BqdAVVkO8i/f11RCvXYL6SKmtq+/Y5lx4MSl4K9qlUptbuPiC
dXOOMFq+r3TMHapuZr09Mqpiv/d2y8x1GnhVaFhxhdi5EiSu1mCPhM/0rng9
eEXtL18rS9ZLd5QHCYXD8LQmEwVdNGE1xNbJLP0QudKPx52J3wCaWxNOoRfF
KIfq3jzOuO4JEIIVwE6LnpwtbvXFNemC74kApBdJ+bxuq9f8n1+Ch0pXG/EK
tZvj5NbGP+JfSpXsHSUmWzGaKcmlh4Z4MGN2j1d11A6cNhM4fg14m0FDEE0K
CkaFZxAlbn72OIKMwAzeWFCfgT4tasecIPTIJ2SKZoPEhUrHMK/QtzLirFwu
920fwHFhzZZVaa6fqcoZTDLJFZWd5hsAa6LW1tfpmu5Y5jpPNrYNg7zVsNLx
kt6V5oFcX+eYwi0GFAmgANEdgestgBJdNV7tazN98BgjpugS3fOauYguU+D6
a+NfQzysTG28Na7hqHTnrxxnx9OjG3SbmKZFyxsFO1SDHD6CjYklTrEn2u+C
11xt0KyELBki6iRqnztYfJf+qK/6YV2OwrLONezpu5Q6kguyvmE6jDfro6Iv
iNkGqrcj0zzSVaZXLb1SJzX0aVCfvlAspzjqf6tCYHm+I3071o7h7odMexwt
VhSqer8wWAIpxS6WzlK7Bq6yxiVHEwEnIyZ2ZbRAq9KMhZ0ZEbx7Qd0qKCCy
fZIVJWgFEq6sSbvvkymDcCFINg4BB+LekW5eVBoI+g9SIbTUkAGR9BaiivoY
WLb/3cSaW0NjvkFZRTKR8cg+p2sOwjlTI9Mn4WnioBQJGy4mS6h43P8DmKaA
ud/EFFfcaNONG7yYgFMSnWveV/B19fnWuDLQGLXfSa+d9Q68coCOKEY1g6+k
/p1gh6E/S6SSELgTJ8TefqfBiDoPCxOsJXxYTQW14OjBEJOL8cHEpm+6MLjH
VEymhx7MJq7w0MJSReIAy6CBsfdDTbV/kHq3kClrPRZ2TVXNH+40WG2ogsNz
Ns/HwitLl9WN9cdcpjwLgf6AADq/XWjSbp7uwrsDooUrXUDrSOR9FAi3kXdX
h+vn1LgZE1LQHGee9qH7rV1AUwH7rGn3PVKBbwLWocPXPKoi/1d5M7rZT5YR
NMLaoORuYa6Fztyj56Rybq6o5n7CLqj/X03EoagJIvgcNlofmWuVTKoOYHHo
9q+nabu6Y7cKOr3pyd2S/BsW8TlxCsA3XeHnaaRYB6/w2OJmIcCtZvqWo4wn
pryELBHTO6E3twbDnZl+XCdqveJj0I693sEvtkTY1VGmcZM2Cw0+yeepKyNV
1DwvI1PTwXdgPmDxwfkFnCz30CrTC5Pnf9XoaXUcV6tF2w1iYs+Xh5wJai21
nm0iMHn8Cmh1Oiyvx3f2n/xMVKQ8LdwclaizM7wZBF8MCrXHtq872K45lwN/
nF0Ep0UcaApW3yQ2a4LLLc04+nytq5EqDpSWCjIP9m8d9yJ3D2JjeB9+z5PA
zoHY/t0skAr3loNONvYEccI48Gg+qYaDuVruMEv+qiogAjtkkjNeRKn6ZsAu
atXo3bh8Vd7pc3PAmhvDjgRx8H58ZFndrHKSBpw+FguL/K+y+1O8PjxOHvJr
8OjqdkqbuhW1i3VYs8mdsblZrC413ZsuZSk5rhVKSFzfsI+zHX9sW+jg282Y
YQ7mUn7cgtdIXyF0aMo0HH5D9VHx1GOOb+0Nsn7PlANAv+Lx3ah5Tt6Qrcja
R0b+/6E47ydGnLhd5tlCfM+VIRg8iHEGGEdUIlA0dLV7bIL4bV6WXUk+G7uu
zuSLUEQoKtvLPWrVtcKRLacamAUloJSlEM/K0hwg1cWu5R89XMQCw9PHtGCV
nYeEWfBenE9kvLRwTuSTYTE5/ecV1nd+RKZBPBMC01zNs5r6cyiupBccvUCn
woQDGT1ovdvJelnvYPfE3FcvuyoOnKQe4dbO/th5Nd3u/NmZmHQtsj8rfis/
XdisJ0VLqzi5ZzYCKEwS+6IUbDeh+3r4xKnXyCQhvZuysdaRYyI5j5DGp3xq
ua0Pi8YDw8OuRcyYxZfTMwxS3okcyFmqIAfQ3Wo8LQW3nSwHW9yVLxR8CPBQ
ZjMcsZSNcOv44V5hYoAP/5RQriQze+AFgSG5+uqple6Fg3iR+Z3UCYyjqEq2
suxo5gl9/CqSh4fjUr450LCFjKqnBeKfz9Y+QdtekEVjWo5dWUw+5AXsadJz
+TyM7b2qV9WUlHJJjWJpNpQqZTKLgTIC3NwWPSJwvgEu9+5mQvZG4UHFAC+r
YmXRESs1Fln/1GT35w5xpzWbm7SUxKzfxN9ONJ59u/kZIol1kYtJtacSkCR5
SSAABix18++vyzxzgMcEk7yPSXgEIx5EP9MnyivDB1QuQLPKnFJSLzOyVXw7
bafYnOKgxQEiFcUAWzsn8UqvUtp/b9BOfm5Gf2s6G6mrrYIxmpEZgHycz7wx
QDnghQTKKLan5Zc4Fw1BXj8owMfeRDqB433KVkg2tXBi4pCj2f15E1zmE76m
TtlyQ/srhtzi2l6xgxfH2OBmNWrnmGXbjqHi5BpZfbL6/tx+jNeSjnbCc3uk
gjF3RUJxqC3J1lkLCaHc/UYaGvx3eNlcK3hFj27CyjqdeLBeOgSt8ym6BfOu
D5f2vbcHAMRwJKGXGQeg1gBLfhHno/eCzNjenyT/p3BS7SbFSLVaAbnCFwP9
XpZisaikTqRFNII9Wni0/5N/qtCu6YRoKYe7+0vw6yLrG3Vd6EV+ctWu51NQ
Gchoiz8OTLHF1sPLjmSorDFhdGe9npw45a9iLLNPybAU71fMiET0RDQp1+p2
bD6R1D6ln3Rx3t8yUHmqA6YmLivgFpPO14yCr536seF3VExK2uYqq77zeM0u
l2gg7EP5mx4T5steAwQ9czrzUBnj0/0I1IrevfsxDPD1anPneJu6TGCNs/Wm
30RxZsUwBWGcXil5q9CFxu0HaoP5CyvXKbqe2/qyR1D7W6OfWStK2kNGU2MV
PT5oIeLJAwUiT1M8p0WKcxYdJ5nYJUx7+y8v/GDCNE0t7mdjxmJrJpW7/ze2
zJ7OepfoAGUnyYwtIsDF7idEe6OqGVx+5XGIYrxP2MKTK04peBT2pFGQdAlN
0sWcdH4Sdfp9/Rbo99k+5ZHgsb4fB9GnHkz9bNnDLa967kIUuuifa2JCOd4+
aKeAQWIc0Af6ZMhdm4VsWKaD3S1rpMl8YoJcfYl5FQbdu0T3R7YdqARmBXjr
KvhWBBcEELSe0W/FZ6W2PpUrzssHhjuHWGD2liJPSpdjY7LrEOQKLOBERM7B
vZegyjz9+WK2LiI2Gugsw/6yTUaU76L+0JDNXRIXeA4VdUVeGU68M+DJWwbI
6UXa6gQ5JIB9bePPFtCobCuAlr02lo34Q2dzVuQGp0J6y53Esg4f6wKcAjfI
bUEBwTTJJq7dSCHZ7plL7eSM3I27lRzzlhm1FB4enZi9ewEI9dwrBWx5Lydt
b7GDqG59dBBLbvkW1YWxcRTidmJD0c1sUAQ9nSSPlF+hZ1UBeYXK+NJZIjXu
Sf7hc1cFG0jTMZkP+ZMOJvTZR5EKgZGUxQxv8LJN7SKfyD/7wwYvAYBJTX4+
UaSjniRQX8CQfnVbd1YFW/FoOVtuCXOlsaM3Oc8gQCIHNpHf7GiTNlDHxDCe
J2IsmSZFbOIFzzbciD4LMhFKkG689OtpHjyUPPacL1N333aEJl4WgvW5Tt4d
dIx5TcZmjmslF7l+J34z1WMghT9bmYZfaTn0nIbwyladllLhhDB3tpNtlLd0
zpP7rF0ajqf0ytn9lFUJYYh9S9Ls3fH7xrxxnzBaP/ZLD46ES1mZ9KTdX2tS
8vsKxUtUHApcaUGlmT67RfeCGKV7AFXY98CNDh1s/wV84YBEa1lXkqunW1FI
U23jprT+vfaCYFtpXf7Nl2G4DwbefJ9tqy3sSMe5zAqNGGwJdBmuHz/zlb7S
8RcdZgLXHGzN8QBNQpeEp0yyoZ+NUhaN5+cjnJjw6fPngalBVgwZMeovEEEL
Onjzbp6fHPCGEzpleYbpGFWCIAdsuDxfVXpKH5y3sb+DZowJtmmcJbLjYASZ
J0llkkcD22x2APydAX8UR1xxstGnqxAb3i1o/4bdoTsiRtCSbELs38HHEoHi
hVok9CBH7y6oA5mRef7rPvhW4rT/pNTyhS5h8lKfX82J1ug6mLVJ53OF2fr8
eXrwfN5a56+cLzKkbx+b9mdDUzOy2mlrUkw2SyPMBbB7CDyBPEuLh8PMQsNo
VcEX1mPl/+/oezGI9xaZXxnTEJQyKsRnKDTe0qoTcli9yxebntO5hoTgstWo
XptjfW0kF/OrHipb089KdLxucecQBNSy+8b0OpKMiW3gU25cjGzzUmVWcebn
5gJa7Xe5PR6nD8sOc/6AxALrNQOIshm5yrZIJG7hB5Slf398S4SU9P7DBVa7
rCqA7ZVvHcoPThgJEd0lYjmeKcUcCgroEISEX13uio99BlGIwarpoIy7QgE8
hpA2bncwmO7AQdljmEESEXdImxduXh+6ubD76SGZGAgUPje4k6b9okmMK0S1
H/rZ+WaOkARiT/z+VwGYl06tUm6UVTpwka09vuVWx6T9ewD8Wrl42x1sRzkP
+6y52n6oQIkavp3n4RIq7uFEWF2SFLPOMrwJfJciI+4YgLHgjjsw+9bEAqyq
u4/6xxdEXBp+o0sEYiOysdh2kX/sgNXV07sSm5hfxglV03g2iQrm5DvAIElk
nl42KRvfWW/+WJ+hoRBPMlBSmQ6BjDJAe/rPen+h/yFSH3gbNqYtvtUprCwu
dQOqBgdqBtwIQzGtcN3KEBuBOH0nuPygIkn4sqzjeWnqG9KnpD5EjsODyfZJ
31rk5I8DNPbEWN7fxNdf4VF6HPezvKXBgi00mzX/3hamqWp6qYfI/6/9ju/b
6+rb4+k/Ij7rP3KBm9g22p/dtTCdXZp7bar1rR+bX0PV9cxnhd15rx0jMm86
gTuxSb7H7HS/tKvdLe+erbwSo+LVXYNySd6mHnTs2HqkJ7gQgy+PwsySpeZq
OoGlir6AoRRUXw2F4XqEwsK5DpRhezrF2TI4WnqCFiW4kgpBAgcc2ugRAgwN
j7Dkrutm77Obh5cbI49l9BaQ/Yrz6BPK0O2+dVD0wRcbidnf4cSpUoSZ5F4A
fi4ye1SeMK/7yX4j2fhZP5sU4dXhkJIatki9/yNpd7WR994gTl/ZIG8rHpWC
/x0MXcW1DjxPgMKz/7iT/y3pkKmFbyJq03LOXVeVvhqO0KUKqlIMJwI1yJHj
pEnTbRszFa+R/T4cc/5NL73XwRgcMOS/6h2h2hsSxbwEjh29nZdHDae0vBLa
V8FpQk9WQO9WgZA4f8EyUZIA/SErsi90hR2SVRhC+3FK/aB2xzYIhrCAyA2s
I2MmOSTM5PRSI+6ZrhmsiMtj+tl4aUxLHl/pkZRHmuHK/55wzRllq1uAfprM
rTye1bY/I7S6G33PTcy7gMldcsgsJkg7m5gPvPDLDioPL7K9fRU4o67H/3sI
t2k8jtYE5wJ/BX0/STAv7Uoy94Kh67/OyQigzKVnw62bfENFn6qoGtIgKFNx
jEKHiGNct6TOOBHgsGrsTFobz+qfcywgpIIU3wU6iNExeJeKU2fhEymKp91/
pxUHjmx9dNAKsZ2WFaoHF6pZZdj0OFJ23BtnCDWukPlrgKcSq0cdxDa15NJY
pgUm+6wTdBPngAzKia5IAvYgCkcGE7Db40s5wVWJM0LkWZ/ygWDAYRkUc5dj
HKBaP2BDg8n78qfsvhPUd3k0k23ZH+Z5RCCcBe1UMdxrqGFZzGIb2aU1CscD
jAwjxiAZ0/ZlIyFyB4HXNTP0e+6L1LS4w39EWUaB2QIqUW7mMZauG6914NDf
Hw==

`pragma protect end_protected
