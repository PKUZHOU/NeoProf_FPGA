`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
S3zXcMTYVa5QOlT+BY9Pf+siTzQGbgNwjVu2uvfY6N9GZQe5u6Z87z+ryDWbmjik
niJ+GFvDuwRzYV09otdO1G6RxjdQTsYxfWkTdK84lh0CGLVIb964vPtZfub1MDPR
NHOfctHH3lC3KT9NepCVXEBj38u3k66yvwTYdDLmZWY=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 31488), data_block
Jk7Pd2gzXJ66QowXqRhhrTxeBxRWaNIjgtf2+1/TI40b+eFeyTvX8dw2FlTZK7Wp
pwkrW+ycIaPftOQPZtdvDYHNdKHhpv4L8ceOG1LHFoKaQ4Hpf9LRMhIT9S0L/xB+
a+QpEGRII0vs/PIiz7vRHBdDfAovlAIwPD1NhjzVo7usQ8SfmRVWKDKwCgX80Ayx
0nuX9plvE/DNUDKJuyA2Q1KmfvcAWFbMFMmsbCsu2LjuSDe3GDPoCVMThYOA61S9
KMkBJ0OqMiGyqMXyvAR1kd4oA/gTQPxSdkDl+zcr1JpMyY1wM/1vQevQZyMJ+PtE
dIJtMeGzbzCY8BjKFKLWg8uwfH89c/BbK5A7E9NQWJbOSp7KbnMYo2P76cKlyp+M
Rs0UcPS/qWf2AAKoWiikiuU04vcANSgskJffJtWIhepN2NR3T5LMET0ptfD55QHC
65gPv/nSo0qnpIt1f9lOnsBkqCVwJiI2X8qbI7Nhx+gCvZKNSSShjX/eja6pKUnE
3Xpd8Za6TZxVFV+jIXgPmpEsSSzzOL939w/3bEdQUVgi0k9nlLzy5nBd4S0wA3jr
nIFJrnQqhvnIjVSyhxdVGNwLw9xgs1krtVuaTt+1J2R/mG3wVcnE1wGBrRpAcuji
tyY+n6XPNrZ7R+iTRpjSlICptGX7VfYgWAOMz9Enlerpcb0gicmGS/7TZPwqftF5
mRE1Z/EgxE+ieab2SmjjWlOFn9nvfrTNByKb/jiT/lwsyCIUh9W7ANzGVsgB8qON
JbtkUOwx4QY3q6foVzYQeQ5xQgqq4hr/bpagRNPzDWZheFUKqffKAR4tJP6SLBFp
MfBFgL/WFhAllaHaRU9MqOLUid5NMCon55qwn3j6gNwmzvLkJwN8U6cq7CkT9GvJ
o1KhGUf2Toc4WE02F5uyaOcxsJrRY1TmE8RiQFOX+uK84TK26tKMnpuqyHMr7DVO
nL0C48fpcSSW+J4BjrwAmadI/s+P3C2gRV115o+MRMPLcr6b/taU//7Eh9+IXemE
WWrIC7mxbiWyuP2DTuCkgIgk17G/2NFI6UgSqXqKleW2ofB8jZ0tKSJ5KAkUTWcB
aUoxakw3Op73sewMVvK2F6g+9E+K2gWY2OsMuFiA7u2F7yukJWPX47HoG2fZDNCd
xOV+h7l3dft79J8kgDzHtZRB5n1Wi/+QWIihgf3YCYBq3k2AEulgr1YUnEAEgJz+
rtKww8fIaBQJGXMqFQkO9BEMm6Pwd+5UODfby3kv5QMXqlbob9seuHgvh9+8ujti
MOPm99Q1XAHdpI+y8wVLjW+ah9lCo6DtQoSZcfTch4c/xD6h7nt6Y6GFZ8eeCOLA
g3z63Bj92HS24Hij1IeDQ3fIqRBZZlEGEJDVDcjGNNnwbzZp0UGslvpQv07nVDef
KunBwTOrgxz1MsHFswdmFXuSbM71l71OqILVsjE696RTTx2x9vjG4WcNbnibnam9
crxvKK11Olhag4OGDI2xhz8vsuZTeWlifJbkwawvtsew7TsOAP+2cgJwzali02Rz
n1n4+S+qCBUZyIRg1w4S4rmYPotmUuJpeE989aOjq8GesCTSRipK6KpjRme2yq18
FF0yPwUkRu0+CNwI1Db+e51Jeo1gEBo2Hf5AML6cpJAET0/FY3qdFI9L+sJ+0L/l
OS2M3PxgfHkeNLBdFa2Kc2mK+aJpTikoMIHbZ9dU9B1qTg6deKxAPxRFFWSGOGFr
BYDbVQDdiY5sNQGzs4uyNrMifG5Tx8dn3vT6gjAga3iSjLs7LHxbFLPc+bzvTWVo
YFm4QEu/MQ78KeklH3jUtqlo09eAnnlCQs1XY6Ch6mOxefo0lm2r7YWE88c2UTDU
ZHS2Vuep7v95CPTNU0mTQpXl+a/F4yA4R/VFb/QbsmeyVFiiKWf4MDFSa4m857h4
zfvanKAojgVFy5n2l3izQhBDgmepmJKlmwKsf5nHlR2SBUyQmc/XHe1TdtFSABkS
0uGoRXPnVSrtTTFEZUpF3nyJvYLgnBIkWn++f/dT8tTeRDl+uochKr7VHu3J79jR
xhAh/X9M0QjjvHEEEClZNxqfnI6MznPlmGv02Lin4Oy5MWUumUu+qn2p4SzTCZGt
yUgexT7ZjlDv9M58/5fz+XelLXPLEU+ZERM43L/N+7t95Dx3tPgR5T0uEKhh4+1A
H/OezHY4HW2wE2dVDDcyDp8FRsXDqZVbPw5GziIpNIxw+73pgW3GNwkaH6LobrpD
DZS3PJ+duwcAkuks5gAfLBLAuK27zTIoix6YddE6UQ8ELjKeFISCr80BfT0vLCj0
1YgOYfgx+P74ZorG0dxVW4vmbTHeXXM7I29fs7JJh7oPOHd6KlLvOWb7vY1m6tSR
wD4t4jYbYTv5FV/GbdIY0bK/J97gUlCmO1xBELj1fF0CK4Q8Py9rarzl8tYUveRj
WqPX/Y4TVTTTUCD2ela1OhM+b8c/x1ZrENig8KTVEs/IDGNUmXbQki4IAhrdTv2s
2eyqvnSgaGKp2FgwcRq1vNKKNE6Aua2IwPCvDXWA0AzqIbA81KEMo3X+MFW+gmQQ
TlDkeGi6I54xELP9Py8ONemVYELU9chCdyKRDUyNPGnY96UB3PkXIPFnqjAerCNR
k11Ug5hcLSqlGago8KaC66nXqIErmZ7BKbKmN5ne6WTLhGIk5KHqA5odUdDxDvEu
UcFgc9rM+aK1hOre0Auis+a65ND/WoJXghbwW2XAwrZbAxHPB47RZehYUzuNDMWK
aBna2H2l666nveBv5Ye9+EA7nZbXYgnDTmUygRU+CYVYvKRKtTUQSAedyF1uT/t0
aEHDb/QI2HGXB4QfgZdQL9Lgp7YpTZXAdUIXrWPy63hR4HZ4jgg7+osYsu7BxCma
LseCMTew5+Rj1q5/jszZg9QFvlpYQ9jzkBPgVbl+Rfq6JWpydPZZnycc8hpeo7ye
755QJjVu3fQ3cKXVrvuYlv75zjx3uu0pz2tdpSjU1Sb5FINmqrIxtZAeTUfEJRDZ
wnLLF6G1MrP3Ub8DTmAz+DydsK6HQ5chrY+PYRieCdMtlkupwkDyr9ScP4XRIHzF
Nwo4d7ftI2EIjg9pFqQlUCzl0u6l16ULIv/FX3qkJq2TBNQjpWb7rL1oOIe97NOC
jRXpRqiyZZaXyAECAANIc8v/f5we8Dli2K81YiwGcYn6S9xrdkuEA7tq2MCik8co
HNXX4u0aSDjiYd+NoZcVqkxGLagYQQP5TVDDMBF3SB/ZxeZ88BmFmKpZc5zhhL0T
ShbtGjUzaQ2r+JCoRJ5ztrEWpbsQm648IVgMDqnw2hq/SkTdbT6MFnbXXHA9DqqA
ec6DCIdxLzZ3QgtZaIGDGIlb+9djBSgmQlDGweGmu8oLSOk4ZCXxrQr7YNxymeU2
X3JgDQJIzWjlYEZaiBha5wdOEXF0BLzm+XsTn4btmUKwB/8VZ4mdd7WQwU4GQS1x
0fEY5ovIMm1fJ156LXBXjxdm4qoMEluJlExzDBSm52a4rBiUwdE5LVF1cNDl0vp2
BNsyt00GnNXZPXv22vUXLCp7Z/fBi8sjVStk/YwuksOBo15rSImVybaWxtjNCZB3
Hrz7kukG/vYvcNnWzdXGM6JXydG6EyEdyhCUByl4Sc8IH8YXs+IOaV4TJhWbtb1X
GEfrka+seBdcOc6Kv9svweGHX+Qn1X2ZGxBp45XQX3LUQwZqGmZChKBl4G6NviqN
KjuNQ20lvIzxNFa446cUovqEZbTC7gJZHuM1vGgr7KHxvLTQVVUESgxiMP1ERR6A
uATQ2+fYjcx9Hz9srt5kAvfN6QK+dMfXL0YoY+KFFwIJT8y77oeswysGmiPNLUYN
swNDt4MnVpWCxT20gXuSVY8DCaQ7oLMYdOyUbc2pEO8y8zR8ey1JbkFdN/Nel9pn
VGXC0oELnjLgcB4u0CZeliTIdAznLVJq+qj4A3KfNA2GvmjbbPQAfL0J/eZWjeGn
3BcxFT7Li3T3NFWW8o3lBMb6LYAUv7hIgoHAMjvopMTz3HJsyz5FPKhBf8wJZePI
b+2YBFH8p2scQOr25zHehbq5QL910xgpsKuYXKAYvY5LGZqezULST2Oy5uXuMUEp
6Iv+sNPQjgUmpnclkhvCkfBNnMkxRiLyqyhMcaAokxYmQ2hKeLvwprsAS/Nzn4gA
ReRAFesjoPyUFE0aa/yF2DUht9SKrZdTqsHuJvLi7cpl089jPcishoR3XgKy5/5t
Nl23W/595sI3gFCkx/q5dvBvWkHKVk6pdB70rkc0KVGCP9sXVjN0e5IX2xb/ZZTa
7SP+cWU8zgwUu91zlDh/Oi/OJSR+opRK/TmutK2r3cygWZAEzAxTW2yo4P3F/yTb
473CaQf3KrlKdCvL7TktBs/4EguJ7H6AiZTAATCGX/MBKRg5exJWZ8Gu+M0cAbbl
DmJ+W2b2Gt90G03Qyw364U/NHEDn3+xznR3MAlaFobtzpPHFdAH0dyd21c0AWyQc
QqDvNg5CsyX0/PrnTRVQ59OTHJ0135jIfr87cdFpIeQdeYTOcmetgipbYUGZ9xsF
lhhonCkPMQy5thTd4ZFVEJ6XYA0foU0qEELHnBfv4/h7R6MHqXmYou2OvE6fK3l/
q4/OJnhNTCwLeY6Qg4XyLyyheSKCCNR0u6RwTaVGm3drEGDzdeTySBiqBB1tdYkY
4NvHcL6jq4n4tt5wrxIvZk38m9tnbnDdZo/x40p75IcP3iBnFYdYsXGjtSj6UCtS
TfUNPf/RsXseTSBIbnCvn3KoM1W0fYuMDhHwBw9oEBwCXI93rnM9MYmDHLHLXr3n
czWKabUOduIpjtIPNTonjJn8MhIhiU90WIE/TNv3d6M5n2UUtEwmo6TVt1TZJx5C
m/pHcCCb/aIaj2Bq6pYKEOKSJpxQwn6iYHfhBHhGfyV1VKeEtiJ7x8nsXSYsZUGN
h0U/lNOFm7Mgd4p1Ev/B9Vy+aaFvlB31aBsqQRM94oRrfLgJvA9AYP3/jBl7aQjv
Ze8ik8iz8MvS0faULuAjl64VHBd6PdjWTx/9P0mkNizGulVZn6C/Z7QwRKTgJq3a
c5I73aAeMoFF0k5ZZ0cEuK+RTdzy18QRICC5PV/IXbumNFkNqH14Viyb/j20ujvd
DtLmRsnNevZuhPq73sTkiw2X7OeUvSQY33dBStv7At5HdjpcoDy3kGJM2CoRE0Zq
3krUfI2unTpea0pFQwnKeZCrc0uNh6Xctv3rg1jGOlX6jmAt4bqffyu89wZ2MDl/
BgnpOs7Sfi57SKchaxHxk9yGLQMiLtu8VnnQXA9FL5KQKRZN9uO2xxe4wst/tvyJ
4eiB/mXrReJ8rwRdg7bNxZ05VpmsIbb6pN4syu9sMA5WIeO4RFtIrEp9se6w3orQ
rJ+zsyaEDf/W3kOckp6D/lEt16kdNEr2kYEzVgPakVLBrOJxuUlyP2kY+PFxT9mz
OioQDtgCvzQHJpW2k0iQCFQFfdUdTW20sbw9cIX5KCuT9oRk4Tj0FsbB2LG47cua
nwpKro3rYn1FfimYKfKRozAbH8EmqZge7IYiBRYNPx0wawbqdZWKnqpe4wruyQJP
gvCRBLUFKCBHcGHiTCmYgfMGeoSRyKLwjGi8W6EI99gGKazJdQq+WDkak24rjHYe
MJ2MVHh7jknOOyNlD00KB8rBOBGF8mpjl8Y3n93h5sDkKtbbjkeg11g9HhsRCPjN
Hf5U+4EWWlLfguuQ8L1H/1W5V1V6zSy5oUQjmyM9mLgnvHpRPvLfDwRHNPE5NVtk
029hsjDfsuMv38bg5CkeDMnnu0yLqVgS6iE2XyHJU7/ibL1+ybN3SSmN9S2sqhN2
cYAkJjDO3TWRyx4htkj3UDtY8smuzlxXQ7rsPEDuN5lucD0L9aT2xI7PeHPMh4yn
u6JE3wEBaWIJ+yJNisMl2NvuGk3F6TxGn9pkKNx+PVIrZGZsepnzI6tukTXiewGL
LoHBW5V/Ay6wAFATsw1iPcTDCDK3/KC1yV4/n6MUm/LOWYM1coPwuGc+EYQuAbeC
1hkY6aQHtdW4kSn5Hk+AB+Szulk/LHEa6+i9dKbywlYoql0biC46nS+81gPEF3ns
UkyGaWXucYOfzm8XyyzhM3n39EDdJ1M+6Ww4wl/O5mdQZ52TeUAD9AeOLpBtuUM9
FeeNOikaIKdNRP5NxKpSKyOogyVJ+VEjHGqA5nyJ8dlhPjYD9REechkJppuuzqxn
vw+YpAasbzbBBXl5yi3xaj5xLJ2QEP9hNdJ3nqCSTFgbWMloelixUcGW0V+06Nik
1jalfaST9oIVXq+tySBS1cuZYIPHbEhoSchSTfgMqVfbvWXxYDJQM52yn0OTE693
uB3dOHnVMshbrV73n02CYQZ+C8j3Ko6Cmr8EogZlGEPL3z7pgJYIr+KYw6WVLgTs
xlXbJ7wLtbmPUYmN1bB7lWk3VFrahswq27+IV4ysy1luj2JimIR5F5VpnviKDyUN
nW/duGIN83BgjzbTvTX2KwNu0p+3E9d/hSye8fHy97aZsY8RI60bLHo5m+FpK3Cp
OwlmI1blSwU6UZOTea9x99W+N6j0GxqdAh0BrbdhfWhtAXwCZzweqs2Kep0k9z2L
6m70BnW51b0lZhRWxsnmU9AUhmXEDmuyq6pJpPcb/F8sGDUINf3XYpAGiIxU+I4+
MvXAwj3eB69egqf076kp9vWBqrjQHIW7g05x29B02Wir7rworh0AaLd5SOm4okrG
5Kpacf801AIZ82/DUeF+uAxUMKORm8jWRvsYznnerRuySU+PFd7xmOy+iu1U9RFd
UI3i2E0iNEz2Dsbvleyom1zPS5VHdT87AGd0qNSuVKoDhieXUNJJC4IX1q35J8wB
s7ciL/m1/frlVFhy4RYa2KQ/8JHescSdm1Pkojwm1VSc8JZ1ZhUFZU5dp5uzV1lF
MEaYiL0YktE5HQNk55EVjal1E633Hq4I34IDmWbiYTVXtXgs8yoJQyCekxh2QGe3
Eua/C493LCcqGu+Q2D2UDjdbBCB8MkJccEKgyaEOGxELviW1k9mgaC4uV07U/7kV
eUl3EPEDK4P97fI6zktHnbC7vU6RQduncHafY79Agjnc5sc7POQ3AGKO6SLrAsQk
rA4CmROipMKc8qtyuaeh/qyHXe92ErDCHwb7Bkno0PN05mqvV8009pHxQsEpoiqY
ivnW/whas63xcFbyta57m5fsLjXlw2zfslxNfICvC2/y2Tc9c+pf4rRbWMJ8R2pq
4acBMque2cyexOGBNdfRRfwDrgrRZU6NfOf2p5xIa2T7rN9syX7qf95VXzOS94an
5qO+56iUYKZh+pW+zKZvGatQ4Ujw7BTgSsMrVGJKBSRH2sQhP0TWiUyOf6Zw2qj9
kSNV3g1oL02RXlFJSyCm1y+Q3CSwjFtmzkCuapiFGODlmiWq68UK9gYPBQ4BbLiD
dNJ7k0M86UdZXUzr9AZ2eXUEdy4bxQu67my+WhE37KeSvwk0TLAYMSJchRcwIcoH
8y+KMzBV7fTWoRBBCfdJc2StppDz/ZimQPi7+wVBJ2j6RiULuTf/3tKnnSTO7PuW
s1WCTeAsLHVdtTrilgXJ2ggplKhMStS0oK+ZpR5lbb+jK6QhpPR9cUu8Wj0xFUri
+u8HW4vmrOiO8yvY9Xbkx102Yi3XHYxh1v7zRPJ2I6qF7FtpZ2ZDVnXKvKhK6Bp2
4mGqSpxoKC1YfZhz4G0pgKyj2f6PiOZ/KxCcC+l+I4y207EMENSUHVA9RvRnOpGe
+4ekPkQKVr/BL/bsdSdd7Yczo928WgXyh/vvNXgVprRzo58ao1Qt1aov8t+bq8d/
NV4nUOW8szst6gxBgEFOXeTQ3/Y1l/5hwFBl4v23C9gCiDeB51hfE5ZKhqLs78Un
I1lqA68w1FAaObJk45MFohSoN+i0ggyjAjJy4zv6G+N69suW2UJFqsysNXEFaSO3
I69mR0sZNaXK9EUX1XF13isyWvOXQLaTYviLYPwmzDYUvJLkfUC/0VSzF+WYFoTX
BGWig8bfGG187A9B8BYm9YfbZPAx3MA7iJc1i9B45dDzy4EJ1iHA5SPIwZ8y0kUs
k+sEW0Ivk7vXVTV2EnOLPTlmurSmk237rUNdy2aSypWql4+cPXarGUh2B/We2506
ndJ+p80t4VIAbn5zgkfhqi5RiAbN4jpvunKxxV/vq/jeWLZE4kWZxdOuarW1wLCG
mt24GTkkZR02Di/kaEwT8HVt93HY86LsOZzTsG9KMMY12eRIqri0w3UBMfZsWzVz
qQQvLfrFyEii3ImXYCOh9fMsSYg39s5G/A9EwyBeSelVAJtC9XNGB/SMipXKC2tg
8lOl9QyXwRfOZZvAbYa8FgTwoekG2ueE/nJayFe+0706LBi/U65HoWN3/F0MZ1Tp
8Ok6u/CBzePuHMU1lNBqfLeCZzC3AtoRtw0FDnKB8y2NSJpkp/3wuku8XlH7Ga1O
RDHKj+wq/ngmynFxsZc2mO3MmM+4zcw+LBGPJVjccnL/De2eVc9QPtgicxJ3xTib
HBrs3tn/Mpc0ViUJI2FeS8PFm9c9tNSWVYRSidtCZ0w1vX2IuDA2XemiCJ6NyPQP
NPCSIXdb3whionK4tROKcOSSDNIaVJ0CCcHIW9X7VMt4FHzcAj8hekkqDwRWm0KR
g2motqbSGnYsXC9nDIpxZwqIn2F6cHgUHz7P/F1dEJll7WRR6OQHZzYWduvFY6F1
xYF7phVMUCKXPXN6RHoRhDW1OVxVeD+eWmC2sINPGXha6fA9GbyWnMT8tijHHmuI
lUUy6AlMYpNywDHqmfMSsszKGp50R+9eAsb4KZciuWH/8iYs89G6yQj877e+hm3p
+dfTUWATbiqw1EvKtFQ6gyT/KZYiIMvMJnEia8MeEqrUXys5BcXualoaR4F5h0iv
c8+0fdAXjXSd1mbTE2G2EEOM3cFYm69Lf44JbDgWn3Y0VfruSnXQgyDPAU7XSbG9
XzNRBaJeR6OLlVgHVeIU/OE3X3MbgNVGfDdN8ha1FbuAL+saA9DMURjNXRh5v1Hq
NHxvPuRl+kRfRXNS+5UHzU5vwhtjJ4ruBS4YawViDEYJKAr0Cl3p5inSJbhSxOBO
DKy6rw4Soh7NmlVhVtvbV7siHQyV9xuFTVNgs9geEk8iFskm7OOEWKVQTHMsym2J
Go1XvY1zCdYK0il0m/fQrSMu3nxIIPVqlxY39r2/BlcY9GQ14ekcx+a0DPkc19uU
bKe/v3Kdyo9y1sHe7m2R0aKUIN1R5bGEsJmUFpqOVv7A0bPkJoXPLXIRs15582FE
nLWx6pi9g/JWSpjBh7PXW19KUIvRWtS8njHWCqBwsptNB1gfnRBEQu8AX6mlS+NY
n0fzgGtrvR6JdrUvtdBcfZsWYpZgtIQ2oKkr1A3X+OAH9R3VQAMKyL3ZeXTDS2kT
H2sQXsdPCIeMkPhSpvf4tv+i0rwLFgo9vuaZLmgJOiqLVvY2HXRAiuQhZyyK4/tv
erPdfHl1a0zR6Yc5HZa7/7eF6n0pYocI12NP0zoGfA38MlBNijSs+VdYPcKrOq8W
GXWTGyajBRR+K0A7a6ZoN/Q5qSoccCWSrzwzN1j3tPQz9d55ES16jKk3qt4K1Xx6
hK4ILMl6CzaN4PD7IFeKxJn0vLmhpUuJWVAQAdMAwmspndB0NLqYesbDYYuQhwVT
qhw3dS/eo1/8NVg6LYZu1B1QwlZiziOKr2DhmXnfDdR5TBfGyRICb17yTCK6fv9g
4+k0VPdQJ0Cax7z5EKaW9up+2tbJ3KcbBxRnWwGc6r83eRbukhu37Z2j5DzaR9E8
X1bE8kOL7VSTokBaHy4u/UNqCgkWMdqb61HEKC/liXLSbuWSUk774AKO2AORCBB5
Ph4B2tk8BcEEeSCT3UwltdxGpH9wtHdevxcaoeSHyFkaiSCXZjYaIfYExjD3weNk
LPxUvPnCp3ZecBVrMJYuPNVFvHOy8ZThpAB01yVItR9OPNbNkVMIMDv0L0cOVyTQ
uEdgv2MNZkl7NxRUVEXkH6KGxs54r/UCwnSiC78e3vpn8J2ptdCGzHDO71ztXynC
z4Q7+1csu+rHuuQn05y5ByeNDdbKMxJgiLmS1vtxINQ8yTmNuGrQauwzcuHyJ1/2
88wBXa47Mu8QWsAC++B7G6vb+ERH7G++W9mD1nc9KVjsOgUssXqZ6s0xlMdu8Vkk
Ctjz4fal7TcsTpjk9dQ+SO2qXcUBXFPOv9ETaDs9G8n0j+wodQbISiZZyJ2SolsN
PHafCkXoOyCnb7dXnnO2E8MYDrpw3Ek5jmYEyOUw5vyZ8WqXIybqRR0ImeYnt3Ok
qdLPA4MvZ2SDXSLeXI2mDf/S2MmgDsEZ07nRfRjk6KFPTg+Pi7IUQHLb6RvsW5SU
/eSS/V03SbsuKjYJFn6qI5RUUqSjhi3QbPLqVt5wUHDO6dnUX5ohwTobWWDpTEjv
x1bymKDKJqA66tuDXjPMg65Ze+b2PQ5ZWIJlJm9oS5+Qv5BAiXSV1codmF0H6/jO
qAmh2GaMuyoao419xtr0iMzEJjLG1MVhzmw8NyrIMq16SJgOC9K+BN9Qk3l6lUI3
2Fbe2F30miEpRw1vDfdYwRweCrta2wUrGzsC/GZcAqSqE+MeZvFuI4dEt1qKme9B
jxoD2M7RQHNvMxaa3XrudYL8mhDA202OnLcNw/5mVYsPU7BYuBI7uQXNM0/9Xo+Q
JkEdEXvDLVgyVNu3k8MGAIiP8Nl6CAzRvfgjjrQhJB9m1AFTH3ruErJ6cRlSU2LU
NRvsgiL75ZO1CJPUnWJcu7TLODQJ2/veK7gx8pXB9VB6PRs3iz2GJ1525foNu2vP
vgqzTvy6+GA1Wem7cZlLkhhyu1itO+8TKpt42IqJDqRqSO2fhkWntYnj7ON3nbec
EdwPyxkVeZUbBuxHad3m2eyfg8M+lgJKIwNW8M3lg8IMsA/RcmqbQ+U3a+P5RIT2
j3aI5iXvLu/66GBHWIkJzMIlYgCN8I7XzFKkh9JxwIF4K5RodaW/jdeFhCa01+Sn
Bj45WluDWeLh503jRT1G9OaDRh2lsJUciGqxK9S1DfuDLBYyNSD4S6oYW7UEV44D
ORkiBlVRnQ2u9RcKayvEVZoTg7r2cPmGKxMkHti3YwjI+UWNuxvJjAEPCryxBhYr
YxSSdu7/6NY/FnJ5BpYWmEFjQsmxIP9KobmCT8q/YK4dcl0CPXVjP+sEok288Qo+
kJNwiZsajFj7/EweswfJHSXgYzM/1JQ2hcBVQcwNQNFpeLXlZWvLwlDkCzLVQvwk
UZacLRpHiuws5tuH82rmxDIVxp1Lq8Wn9LZawqJFAWZnYPJJc3py/lYV6pL5K12U
4Bk8dVuWfoFF61yrFETmid59YF/o+0BYAfGEq/1Jl9t+X0TLGrXA59eN42xV6SyH
Ek7UnuI06yuQJ4sD8iWg6/nqVGLj4NSk0Szvn+luEfBFGx2Myi0HSq6re8XInTU1
H5MOKzGkKfmPCiEeTsm59kojCfdyl9v6I2ph5SkiATr4ailjXBS0GEaZ1QDaHgG9
HxugtcSaxg0026liC3r5zDdB02Seadg6iHnbGNKOxTmcwrMldE1odJwJNFWalqb/
EY7I0sFK97u7yB1AkYvkOXyFXh3Tag40ru2snHGsZD2sehfGwfpCkzGupsw9QnQ2
3OvjOM++Q3wLh41tfMxJQaNxoCf6EN7X7TE1Xw/ELCOYMS8GHPUoVvnl5uIbVWha
+u+i3IRBRMBCtrnfKF8EfFRe334Cn4AAQrOrM8xo6Ay1mkr2F/kKYz4VDUM/0XoT
U0RnUfkChVKohx1mN8ecJBZ6TDZ4Ogt2q0DiDqAFE0KiCl67rCV/6fDwLGZ4d7ub
F76JLZoUH77UUUp02O1PS+3iAwWeBRH0zqa1MYgKYhMi0YqoQXSlQJSAZJQg/SSb
OR7osswwBTf6GMcJJPXePz8VbHo7iTAVoyKF4qw1dhnLBIuNkoZFshQ7gPbyMn2p
oWP9xPq7Vm/2Zqd9w1xB+IOoSI5o306FVK4OFqNaumSrzjNSoqdOOLFIEb72fZMZ
tXSufFNZWavC46j88Y0uZdUN3vWtiH7hKbetm7q2B6NBuxuIyuIzoTzvB5aDKGzU
L3VV8Ld9F94lycoVKwe/WW+CVE8ODYHH39S75w+79Qm15T5PH1H7D/vhkw+bkiXl
eQ2JOzUcREEsKJBqmFiN9Y/dMc2WUyD9Hx+XQm5fXJZLJeQxV53NDPDAgCgQQoGs
U6EwNQ1bP6T4eepXukVTtqdevCEDuxy27gkeqeU4NgvCly6c64fBJAfTz7oC2Lm7
rxatyqlSYWNWi6aas7Ti+9I48y6cR2exShOINkbGHKc07y0zXnctkTIrwiq/+6lu
r1wwAlUkI2L6FgKQqZ2d1Pz2c5mpIDHJdqgXFsHoGqtqy3Ur7mP6owx3ZBtEccVr
Z0vBZnCHGEm81apxYjTn5LO7X4qr2Xld9XC7RMCV5GqDW3Wr+/FoZGp4jwH7KePd
Zgxr/+/CZqJrnlrPyGaNpukZql7y/7rwjSukEIFBu+U1MJ4LOIh4J7d8p/3j4Gfo
IB52/GdEH4mpSDr+H6IVJYirc9duwa1BUpWFtqQyBa9wxjs3Ebaeq8+W3zlk25RM
yyUacsB2P29PpQgzSKwbii/7mkQ4srw3qZ3Hpp2ffuqUTNPhcIhhpYj1RVNXG2z5
lvPY3Qjp3qvctuTyg5hr/E+O1AwLvEMeZd7OQGoXEpC0Q1qPZxZz8fzRAT1qdpVc
v8tef/D6KJBcv91dsrgd3g6CE9Y1hb/VA0LR0YOw5/zHrqyQkZoPrmb/UzXACMBM
x59XWl+lsjd1VQWQg4JkTudjLmw9LmKEXVIDqNIV0h+hHJU8UofWps0oLQfITRpp
GCb6kdCt+HjObZ4OGlr1L/rIYmStP2P6O7FIwduCvPhp8bMlbB3r01K+YVJHjABp
L2KD8c/SCbNVY2ErudlohbAPpl8BPd+iBE4ZuOGSAoVjRQnRPNh5TNvh9I3UdsK+
HRblNAXSgW6TN42WjS0w7cyUweEmoIIwZviY5Q0d67W4ewn433wUm+1aO+fMdIY1
kb1yC72ngokf0+wf+QFpQJjshMBs8EA2x0au3J0dPfdrXmSlnnp496jUJ6Koxyjk
3RUwge+tyY9EcnboJDzVH4tvFtliGRlY3FHJRgD/hiTiPvRVSHPct59erPB5+9FD
6ywoChNed8o1bAoRXKB5R2YU8kZMNJEgRU7jLJaKh4HTqEaJk/UywMI1hd9cek4S
B7sA0PsOzrPIurJ6zBLgm6fgjZo8kiVIhK7/MVXvr8ZvS4TsTfPGemnJGaktPvI9
pVkq+1UwUjBRbbDifuieYKv7XUJXcarZWVEZgRBlcsM7wQ7d1IUM9ihybHm+WzFG
Fm7tVLSjlq2OYLSLTQOhE4HqPT6UouOZitwhi09QH8J/0FdksyFcOTwgCZymfP14
HA2rWgTB6UGfzQAr3JcHi8ayI9XJkl3ABtAgvMc5J0FkoBWocJRkZTRj3RK4uq2P
crzkEQoTZHJhc5Kw0M+gBOrPlOUYkRCbRQ2D2CeN7XWxeYVVsClBX5fctBWlEHlU
SBHLMqQF7O0WbDeoL6oQbi6rAGPvRHbc819USvzG3V2VlXzDxsp5IRIaq2rBIY1/
Ug0FyFjzFQ3eeB25UfGoXLMkyySgwlx3+UB6uC279IOI4q5IWjZu7C2tdQxLW6Kz
cvhSMwK39Bppst06rCsONDxGd6eozqpHMPUhUa4SNU3bpIz39PCbQitqdnWrPW8M
/4fwi0y4QjOLzFANunGzpqbqHOKAuOAAzw+mCejkdKfZwc7LhPdLMw+kk5uriTCN
KRrHrLrJmwz6fxqZrOdg1AsqPt3QfZOP6cToSMjBErPKrEUUICsnfZGWwKyJMks7
cumJcy7CfMwdxW6H8WoY3hrJZ8KnfZau1VrwTeEEGsOxUlISb4zpmuj1c4B40wNJ
fce7Ey2DsLez9AcivxQwFvnUvu/HQ45idrskN88zgSn28BauTrKB9QwWCMnqWpTy
mrbrke8nDsiyKWVOFW+Yojg7jBPaU2R1VuYZK4/gECothWpxHZNE1+Xpw41bUQyu
auQxeVcdLOZAJqu7x23Lzg/Tbxy4KQLfOzy8u2zuNQwCL90Yl4C9XXf9YGlf4+Av
03zrw+OC2XaIkn2Zxhmq253BwDYLSOsQwjmP4igynO44R+CV36qioP9g5PszjiiF
xgt4fOAp9lgA1FlLaAL4BPat3LVSa3R//75uGtP8V5NbQUOdNHRgO4u2ZBRIUj0R
9KFr5jJAg1W8fqzG2G+F13FwYD2mGGoXIL4XxkZEhbIZIWuPnWNbX9r89W+TolCx
AiP97qz3c8FKHcYOW1Qtk93xs2K8mX5EHOIGU36fy+3p76u2aUnjKnXWxYO1JHcz
5DmZLuBdq9rn+PZgehcrPRK4xzVkxGSAdkuq9vsD/zS9K73lxTgrDazMqIk8HjwI
yjxSIQSjzPqwCXuV4ekpjv7T9JGMLKprPYFJ+sLWZlOpaeXG1ODRap6skTAf7p3g
THkVZFR0HDZRuQYZYZHVv05MbVmjQLhru95ZYvwgcd/qbz4nndT1VxjPJhMW9EVB
WW+6HAXY7BjTDyXsQY88l2mEaokOnXdUqS8IeUii+LRZ7hNBLkEVZ/Gg9BnrzMtk
br1DV795JjyiTiAPtjVzqlov5jYoVlafNYICn9hT47S1+veffC8feNqgDf02Bgv3
D2Tmlb7mv/cQQBc25sW6eTb9iOXKwy7C4WHnxukD8zpSlhtmpLf8OZR2kpt3GyDE
thcDQVraBzD53JiluXB6SSe77CaxWx1lLl/OM+SynMuep1CoR4m376W1eC+Wtdm0
z5ycYjpziFwqXwqIxsqo+Kt4cwsWGVsuylzJtC3X2nvRjT6Q9xafEGSYuH4tEwl2
0amTohV9f/+SQJHGiUzIFI7cugnJoLiyzQJ+AX345jVwN0/NXeh25YeDBaihuQIC
4879h4ATQDzG/gDGHkTtcdcMiDPIexf8Ms3mdXhAs5RnI+/d7yNCsZSMIB+JHXsV
uN3Al8LGFjK2b8DV2LZQzPJ4CgDx8fBZqZ+I7CsjWdiyBM4Elk/5EckKlvTV1+W9
kloFqEsTH5avH4ajM21SVT4qAUYNstLDeokf795DmL4nOBxcUQry3NKmbGoCXpXL
SfXRb5NEeDrAdYR/i+C4WCGES5CsbxZfUkctLv6urcD0Yr7zFTu0wdFTKJy30QH6
M8sLWnCaqndBHvcJPQobTuO71sF9w/82bLSlnE7S6u7wu3VUIRZZSidW0tfAw2Pq
PnqPisvQqkRU/JwUzuJc2ADCsTFaFxhz3egh3tILNABNIY5kfFCzc/WsVBzU6PDk
+TBbqHNF+zXH5HT5UFEK1x39T3trwOLKXBHFgr7bhIh/5cUJqoZVXytsp+SWzTtU
smHtFonN5fTXGtMv1F+bjXjn9qwoCpDguWYIyGg95L/LtnefYftcRcF1K/7gE66P
VMbN4/9JtmoizGJ5arcOpm2MY/VQR9/+GQ/V5Ga23vzFshMJCR7mADjch22B1eWj
GHn2j+7MTOapZtpyOGm2qAsCy9g5/JKge3AxIQgTtSVfbaDjwnMvx1FbTYQL1qIO
aeg1n3SCiwt2XWjx/bgLKoH6lJB953KfrD4hHDLIxPmM4iqvbRSwFjVWTRxn7vb7
FyFw6GSM4yAKzg9pYj+SHukxGOf9F+KluoGUIkV1Y5xIjZMOQmBkXT+dW9tBfweS
DYOIKpiHkCkARpOrZbDisT4J8whLLG74pR6WPHvfB9uRhDJekpTiX0p2zgTdTn1r
fNomSgslQtEcmZeZE4sldSgoRYdEUBOXIVCALHBISkAktFpcxWcAFxfRHtygo7gp
45d9wncWbY4sS4TdEdfXvM1zf69OVMtt/ANaeVO0D4134xIVv7RCfab7qP1zH2SN
REyv2yLQXcZV5iS0mOGhelToys3mDUVhMLoiSz9WgzNp303ZQx805xJIwc57P2Yf
cTW2Mxxf0IhQdrW40AoFEFMRQzQpf6tSKnVxI0M4wIy1OgJavRw8KwJIaW88ktRT
lEqm06ZaKT5wK2Q6fI3uIRIeFPjfohMj6ijBsciz4FmYdmTSkFLhOUjEYJ0xjPJn
ZD0t08qZi4rbcCkbqGKVhKqXcZnwjPEpPvbH1Epuznkp5O3Bo3VR4+DiAArtSqZP
n/9/cCZds6/OW54qj00byPHp7TIlbHlxBcQnUuHKJqqH6qXMGGX0fQvFOvMEyNpe
88YXUZrZpLyzVLkqBDwAjCGGpS5xdpqaLjRpsbJHRJ1CqL4pXZtNiQiNYt7FJBCW
SyKZnGLqoBg6HDHcnr6ZVCJlia3mGW45tCWS4iHinT9PGdhMYGX6jawtmFKEfVgQ
dw5LwIuWBiGT2ozoPnNYEaDGxGmqj83481sIMJei3aedc/wnVuoRvomT7YBg8v8w
ZZrmEBOWCC5mmDz2I28++XE8IZMVE6rDUlLRW5R/zMn8m94fzYovSOsMhLA+IUbw
aY7C/8aG8Cw8YQlF2GCsetSNm3eBoUktgYTwaerRkvW1THwxP/jFvvmB/2eFf30i
SuG44P9GgYfMEXpFpUrAjWjjBRXEdiUTjKYClDH8dCTqu4UdfuPJGvi1zAuv9l/V
M/vB/kZ8VAytYBm0eNXb7RYlwKqvlV5Ap+fNsXJ0hN3ZrG+T9D26iwUBHGvAj3hk
JmGGUBvy8VBVN333sPwhzmlWPXgxfmS0wVGSKil+nVkgOxaeJVPdat+nPeeQYzWR
tH04uFeCiQJW9qGc6v8pqTL3/5R/PpvtPO7xU0dtmaDOnO/MkNBB5bpNTV09cuIp
V6C0BwcCnkVfPFdNmUjVC7htoGZ5gXqPnpE1BBKgBO35s+wuZzd8xspKt63zKklz
yYaG8vdtj1fsI5H91QAcJbcnAB8PdEnyW2y7G393/23jQdTIWmxZQOdBl3B8VvwU
yLR1USOn8a1fWRQIr2d6gTrNSaUCTkgXfji99AizeOwAYtkGrcrfpFZlW+BZKn+i
BOe/tVun9uqcvQQ8ZIZgTHvzJ3K5QcwvLzyZF1xuJRoFrjqKoKIcRmvksbumB0wA
ZQtV+FL87L/nNB2yVgwSZZ3xEVC8a55EJFRQtM06Gfwh/8XNAwxLReuBfMtV7Tic
JoSQoefwiywVIiuEixHmd4X8B3khyci5cRGGfEcV0lAGUrq+yP1Qnxz7hY/mmsZl
KjOPbSsHeRId2V90dGfiAQmNMDU7N1JuQq0ez7lWRVOexTdc2kMjVInaG5TeS5OW
GwSxylUAhtPDVl4uoqQmTA/0VmVDAw9OZbAS6XflC7IcS6/w99RCcRJnPZyXLo3B
6YW6zWzmgKYTXsO1FZb5J0cMcZyC4bppuxQK1PrLLOU051wHZdlSK9zlxTnc72A3
9kIqtTLlyD4TLSB3MyY2o7I62OO0HEoDDNJptxiZqWRNQqbbrj8VjiL9mNrT2/K1
9SDkEUos4CSOh1BYrIMxdkUr17usH9mAN4NDtBUxLPrt+59uqDwtzrzTXWfsoi9f
aIHOzptnzuqMF1TTV8pKMUS10WtvutCKTZnTK5bD0hvdcrk6UGjOtKIkNwIy6Zuq
+FHDzlDw16qbisWQjFqV16P3/zQawVddxYlIKnhKS2n+wTBzLf0zyaXKncHPkKUF
rK6F82hr3Eghb+kXRff3fnmvQeiQqYcbCQbswtwYa8BWsRFvFmghS1vv8oQaidXW
QYKvjL1cR4B9k19MHFBZglJ82uUAegWacvqcjnusKbv3fQhSWpkHWbutEVdD/kgl
y/bgqEgzuomv+kZc8uH18tbsMX0VXUZr9R52Habb5YtSeBcTmMQuDmZYG4Y+G8Pj
pKPRo1B1qkFuxzN4AzwxsumoLXeQgvKUMwKMF7DfnT3Q/HymKypyCWmyC4blLxub
YqLAfd0u8yPsobF/fg4/0JzVGK8jxK2zO0ctH8Nmqg7nj6ehIoFbpkxXXGNkLFW8
NgtxMvNUVTTaq9V4lqGt2hFSGrbw412t0mYflXrmz1WddDkWxTABF0/7VItioTr6
N9A0zHUZW/fvDjlNJh+POwGLd1Q4oEPgCvPXc3b0kEu8L1yrhinI67/3ua0uCix/
WOY6RO12g50lyJXv3L+DBN5rydKPSzrp9gpo6ptbUkijhB0/SJL8FWWLD0dbgRzE
MUHhGn/uZLU7KT1y+EsuBxsnKcMZ3N1DsPxE/UXgzI8BxJ3KrKuK9TxSFpiLX+ed
V7ewtJkBaFmCOEQ51S9aBoo51rLY4NuVBhGR7yW6HR0PgsVTa8DF+H/5AHvJLZfF
vjY5xvnAO/Z+4viAV1NdRmA2LiRJ/ghPwd6cvH31M9v8x/A6BVNbS35yMrA0grPD
chVuwdjwM3UgJK8Qn6qY4yCiCT5X0/6BAC8T57+z7ogoHwpuXg6nu8JmDy5KcquB
gw5MEwSxcHqkOe+I1jz8caZnwwe4VytFTy26ZDpt0P/XluU3UfPd+cW5CKXm9yLu
zPlpYjS3i2kquxfqTYjxJy6Cy0h30Hpp0gw3WUkBG5JH4Q4gErzXPQ/IpO7K/1VJ
MWGhgjB+uM7ahkF3h8JS11TMmc8EvnGeTkeVgTCc2clDffXVf26yjz393qmJSRm3
Jf+QBCLcoMi4EREQIC974rffQJ5jTVEiX0RGKvLvyuy/U9w8M5RItzllIgLd//85
1Y9fgmhHvLD+RqJvTYg44usXtR/9C0ixer1oTht0AJCJQHEjLnaSF3pYLudMkz2/
Sm8a7sUbpaROTLwkYNc6VMnUWfHJZXPTaHuvuHs3zW/7/R9tgbl0EYb4Q5CBaoeI
f0fWZZnxUNO5M/AkN7e1HeszOWmUO4SXcWUlkZWQJvVqgs4zdtctJfB4OoYm0yfs
CnSjIjbfMUYxErjkqr0+yvQAiMZ+p2QG3mlDNM1pw1Dwwu39M+f9vOD2jcuGFNXs
bSUhgmNAV0qIqIoVrZ0XK/l5yCi8m6SekQjuvo4NFx/4PEipRwml6Xn9b3WU+kpd
EzVhACkpNIFxtStiXsELOKohcWbhJGnfj81QCfz9JICat53nkgpHUcq/dyY8TVYh
kw4tj00KxJoYTgK2q3LgN306fgMzeA3T/lbQ/qAFdYaLNutws/ia2zP0t5EBIdTq
YwGjuJuFdOQ/gyX2YVG87OyKeQdqYNghucmDY9eZ4177WocJC7V7iNZMQeQbhckB
bj3EA7uzmESaMp7I3eXjLghEDmjNq2czJSMG+qvMnQKI5dkOI+MZq+uAKRSxi54K
zjQRbbUA4tsU+yaNWXuQ6WUP8lIYp5pOUH7guQs3PncvZfISOZFJeKMByAWYw15s
Oq+YGOFi5ug5NF2O6GG5Zih3uwNULY8Mlmx6fOEOZNRQQ0JK/90gWtR/p66VylhT
OduKpvdSUlkp4jpVhQusJ1CXWULqjzK2yOBBu9OWHaYQdrUJYZnqJyjS0BNf+EvY
x58gIJGHW6THiAuOpu+h15L76WVjcnlueLlMhZLRJnn6l0bQW6Da4Pg0FjrIvFwb
QlKEyXmyErsS4GfDgUYJR9lQPd0utyUvEJPuqSIGRkJWNwmbWPmNWEQtGNpSfpZ0
vXi6XM+k8xE6wioBdrmHtboWPVB/IOJkdeNQkdQBVhqv3qFeWwU9bFA+0nwjlz4/
ewGM2vU8Dz2uodCsvbFw9Cjch7vOn/37wwzMil0Wh0Vac5GT//4HtSRlOczHr2yu
wRSkA9NM8Vag+9WuviSZw4aqk2VFo36nglrSLT3yWF0SJd05Y3hhQfUeAibC0Trx
CH7VhjV3BDNk5kKTWKkxtgLGB50TPwy77FfaDB90vmFADL+z4iIJbfRMF0NXJ36H
aEI2NFuGSpR3txX220KYub3nSnfeDidJlyGG8zHWIr+Dg+kcNLELNkdEk8kyxzPQ
1md2ULnNaLuCGMuV2yVk7TRqj8djn5r5foVGh/HHKQBTdY0jR+aO6vPqGnaQbyhR
llkjF0ElyQARac6iWgcKOOykyU6x95bpUtvAazLNyJRV1lk7FX7SyjSI5Hz6RVxR
WLUWx9Rgat8xb5Yf/44yrvD1HHt2ALStHteGMCC3OX3aN8kxmLb0F/UDzJrN5/S8
/uqnBvn7JBnFFVJu7+2ctKxGgcsD2iHK0zXMPYDNCykXjBt/7fvIhF623NXHomkP
xCxo4uO9K6uecqra0LFo/hi6iBXgMNt6j+6ez7Fqd0s7KPMxKWSlZqPokaVqFiGP
Dmrl0H3SU9pz1ArluRNO4XSELbMmnIRAI7rEecZt1PPzBDaODu5jDPXczXhasCvl
Htnac1WZem7qaSr6/jYCcADhHViaSOEpz+dC0rjaGZG2Ior4FmGRTvhZ/8Bt/jcx
JWkZRfjj5gR3vZw32nihKjaOqzx3j6HhIZFr/aujk6Oxa/06/Ym43t1ZlqWnnfUA
ujccVlaYRK2ULHp3kQDDmWZwRwMNzl0yAOnBExwvpH93Vj2bBB7UOF7N18LsLEDq
SRiyNQCoY6OlL2jiFFaogh766RJS4nZpeZH5m7Nib0XGvc7sx2EZ7D4lGXP92I7h
YFnnYXs1q8vqKiLEuamIFZvbphgyfyriZagKKE2qmNNjSRLdOHnkhxUnJi/y/FAY
lgRYVo3xFEIhY+cbwI4LBNjVGyFgvmS3/hRaFASQ2c1Nz6PJDTg+BIxU7Y9Z5yiy
xcwvcYaHBzyfJqDxMUA2RUKEcPndKTYyE58yTAf8pXudCB/6DrsRq/6waCch8m/T
uKSUrlvYB3mcV+XKoT/cVcDh3QBcuNlooGrFb3PQt8Wz2HMvfz0Dt+3chJIGCwHc
L7JfomB5tomGKDKOzq45jhaU35XoO98th+jo8KMXpqv6NPg7hVWseem4EUbklDx8
893lAoQsErJCmTPBMGhURaKyioIzTTv2uOW/FzmFO3MYiNqilldQtIFuGFRJyXZR
hxOHXi6ZPFtHQ/rzP/E7bHMGbyJvhdo/3c4YoJDjsTpAXubkWkAriipGl3jXxWTa
P5sHNtNx+WF44Al4Jd2XRLT45K7b1fawOQEAaBgGoz3XimTIxbnXRejBUKOxiJyf
KUhnno5XwCRwFrO8beCTGcWo7JaUjwufcKfMbk2IkaWsumozOMbFkCbRXnk6vyl1
FOG1Vf9OalYYPjy5AeO6sulKCtOeEDJCTOWu2U0Y8na6Elu5Jj3VU3iT+FpfKgtv
vo0mjUK1V9l8k6PTZOybfmI0/JFaxgdkGKiI5CkxpJnVtYDY87eAc2YdN/+9qd4L
9OJBS+ytkI8pF4nsHWcTdvgUl2bliPO/R2xSXdgv1hxwNbrrKqCUbWfwbFEhVO26
n9A27P5DM6JBC34opSNo+MAn0k5mke1p+hAzk1B6U9n6ELDFNmm8uRJo3jrXUopc
0O4XGcp56oQOu9TltipxKsbBlHu88OARld4SrcvHzWk6c2nJxDIuslT9TFWuqi7Y
e09jsXC6ng1xnVNWXdzRdD33PaZqvDLKi5o3iV5g++eN+8VuRB++tczKTk538J+N
kC9wvWtCc+Z8NtcngHyJArZ5U6fcgLFmRGne8GaWDwguG+vG3g1UBK65LnuOIGnc
yZBaRcM+epdL29JJh2AF9VQPvXuvrQv1c6Nf4RjHO+Vk1iZ0/xyvNnibn7qd6iT+
YPZywLcaI+jl9PHnrcCpiRZDGznQc3qI+8Ca9OA/ReYqleaJkoyWU1G1brZ1Fo01
UjV9ClATRP/GBQNjJ2J8cUKqsArBEQujl7i8QRq+Kih0jTNKU9li0WpveJYmLTas
0XwW3rFVbLz6vrGFzWW9R7dDonfX+DHrRE6Z8QKu+7RnIc/B4Lf5DMoWkf/M7iG8
2H8JGF2MYi1hNd3bR9dQ42gIeLt/cL8dV8sKbyUIc2i1Bo3EgetaE7ML76GSIZVS
JynAVNcW0Bp2t+RpUo+saLvnzHnEBfn3IEkxlz7p9iiHxP2Pkl/M5GCUO3mPdMv2
71ys6JaMSaJgmhN7EgVqzHPii0mlxALLG6BjZ1yJgR30A82aEeq10EwkYwj2+Dh7
gsvDKYmg8TJ5Fm51LtoaiMV2AzO8GtV+OLUPgB7UaSM7x0dXjspfwEnhnfWXgMTy
LMhEYNO+D0nNx+bPg9Bg/PjoGW1foUnMcC5Vz2EUFQXFbtA/YndRqYGDIgjJ/tpo
EqnQ6MKv8o+VTKppzKYEXogd/4hp1fUiAHSehnsfGHqrEhQ2dlDf7wz+nnkxRsG5
Ysgtw6SXNdr1ON0tmekoHuqUf301lR1FQYV89+YC0DL6iZ8oTyzuVPOGKoPeofFk
FHJs57arnH0FnEqnRaB/XlEJKl3tVNnVqGr30hbCQElFhrr1WwXXCckQOoHeNlIV
jbPwfp77cafaUo1S/y4u9NYuovZn5FuIVMgyLLruKKaBhfmFYzX6eQpP/BXLT7y6
9zxQ8TcMxNnlcOJs8o3KnBVfM5Vq02FCkzshGNDh4K/gAlRM3PMQS7f6YrpQhaxa
mR0EAWDHtAELzZuHLY8kJ1csbyuAjzX25/9wJM+eMJKfOZXfU81YzXuvpKaDRg2B
apIVIKvWLPnmd26xJOWhOGsxF9aXgmffvpZYBny1tArI/kWVU2XSCseRBoZOLx6y
pc+aBcFe9shD4APi6zcoMTMvPsSEkFByGykXsRi+yryTZu6M8awbF5vXRQayzCw7
D/CrbAOfoMHaWkZiDB3o+HgnfVb+5w/PSKZeCROFgcL4yO61rPbQZ5u0M+kilnr2
G4d/fvEqMg1jOmwy7bT+WHBj8JVJ7+l5TYOuz1yQbne8FtVQSXMWvAAqkpfFii2L
Qbxbbl/iWs9lm+FIlUwAErU/n048GTfniX1KJFldm5Mqx+TEssvzFhPx8imdpMKW
O4vyBg3tCEIDnITFKUc2sJ5YgSpdU607q7ru90hX2q0TeDdFFAuznzsD54ofpDfe
4pl6nG0nYsHtXsQ/MTDr3mu0NnSzeDMIUUFLLnpBocLbqVhv5MGo9Jcs++XHExmw
PxRO/7fsPEem2E4o3Jn7D7NXo2Ymu3UUeXtst1aMFHx3WgQakCf6bcodBjXOPf0k
J/WejUpr841oFFLf4whPb6fT+/QNQCxE5rPctA54Zfsp9QZ8qU8Wc22YOmpDf2/t
uvYZ+t6aNcYRIH2q6JhHW4DdUjFutusIrZ+F9F0kEPKsUIsqmf+9exxLXdUBB4Tg
5g13w7vvDI32eLl3txDvlli4bkaAprYCEmsbtvWSQVnWDbLH0rrJnQ9jbdFdBOfA
fxxpEFmiGQ4L2hbL+lUoQl6Z8KN4Dp9D/VZ7cfyz/92hvDF+Zw33hbux77KCdBOX
pZpZTiir8so+WOL9T9a7dD0ftGEkYn6lxPD7T+wjvYkqTl7vytCo0rDH8P9+AyLL
RYWtBtiX/6A1P+MZBhqNfvyTbtfviJ7Kihn5rhUEClGlHNhLiF+8vZj54Nbf1dBc
TqlUa9HLzhh5GEmOeXVNylKOZeo1shRdWH2YiI0f6ei9skNrh6R14KAQdYUA+E8+
srLbmLBPAidIIkPIbjAc261HWxRq7nuYyucujx3IaCqBeOUnVy5pZuFOC8nSPh4M
VHHWQFecqg2x3fSeqOpw9A2WpzwOk1+FHGonRSr0VD0tgFu5OwYFVODrSb+WCQ+G
huvThPc51MLGaATNmW+SrPv7dJICNpReb21VnJJrVa4d0bjb0joeY1UQMIUZsUGm
IKe3zn0n6CBbBxZ3aGwOHtS+mzOsOvN4SEPp0pE8CBztQg6z02yLt0GIHcr8fyea
BeydXM5w/c4yCtSPqzCGnVlcKi2obozAHn4TUW/9bU/CS9Urx3medqkJLJA+aF+D
TCKAFcu6x+O4vlhColFXhmm5rxagUf23+FFO51NKzPppu1fDACvb/DpcY6atPhZN
fqVEKJHhtZY2AGR+NBs4xIxrCIgmAhL6R6TYGmbZC2w8OHZW9ij7POceDz2EsS/a
vDPCAnyCWP9EOf4pFskcbmwZ+haom+ZtrNZ0CQVTLk64XQxpcODfY0VNxxC23Y2K
6ssArMzUx5SFtiq8XiP3TSbqoCR5MVPWJJDtRiq75xNQPXTT2xAd0SP+Q9EEIM5R
4MucdsC5Bau9VWNe+jxo/aw66SbaNDg1tAzm/sZBsPpntByVXJ2C3iGRQgvhJb2U
JknULyEFbbPs0fpCeiDHNn47WomB04OEuisQdtusMMQogcWNXKs5ZGNMxWd9ryZX
GXmwfyHRjRctGTAQzO+lUJy4TD2CAiit8uW810GkBVjkyi1/itMjAmHh5ZdSXhMM
oS9QCx+P8QjFRUyCbSCc/CjarZn33ovZMcKhp+Ubv2K7PTLGmjBgQwNeoXOmViuz
5g0pJY3e1305vNrhCrXCdfseYescnRjlUa6yMYvLAYx6yEj23GXEFXdEYher+ynK
Jb+YGSD9ZKXlkXtVz8D9z01udko5yotIIWvbi2RW4l4aUPe6i2F+jcSSvx8uGWqi
R5pfCshaw8ajmQD3Ri281B+mHHkQIXbRdlP6Syhc5mGcCF57HZO1r3bU2n5P8RGi
9pnuWhhCSzBumw0GkICbLgAIW98Pui0u1UA6tKJ75OaGnuRKe9UE2tkUhxCgqwla
GIB+OiByRsoeJ5CBpEilme+jZnGLfJoQS3mt0tnusO5kMTD1EC5mL2RwoiIAYljH
ABKO4BZadMs5fpCVXJxoF50KCfAfKJwucbXbc87lVT956BNAwu82P9pROfEsDUZX
80F2gQ3crD0hRY/YYzfyXLMdu35CNHDTbjYYKleHRYK8uIgHLEHwTu3l6uzWXzLr
pZ9mYilkZO/Jt0EnXMb6pVbkZJtfAOHjIiHwaC58avldhl4e8cDNmiQdJZ7zDyit
x/nqXcTPw1CaR3iPSE/GNBTnm/yUjyWkSPa6V3Ei7iapWH1VteqfXi+cjklGqf+e
h1nO+kR2Dn7Ea/Yr+STH5FfNZlx9O0rWFq5Wm4xtzDVBOddtlqHy8Qlum+lrfcAv
x9wLDvrmUlrhanYxBrX18pbi4q/EPaFi4OeiwpYfA0GUuxmBsOIaVAsrIuvrpRkN
a4hlpAOgc+6m5H8MESJrb8i+AkUBH2jNKbLkQ4yylhPVe9oo+lwHk2PdqjWAGz2S
+7mLcoP2DnpwoAQyQhHZBSZVlRLoxU4/qWKdVCaT3sFNC5v4+wYUAvDKNA/7v5vK
H4xcKQ05tIwEkq3cMP1MCQepfX93JpiFZQIYw1GfyqxvQWpz0jFuBgCL7j8bDwdI
ov2IMFej8Tz1SUX6bGd2HtbCB7lAR5iADdiYMzZbpZi2m0cmUqUWoOl+4cu+GaQA
0hwUYSSxLDkBVxuVKAmNplaIwRDPAYmfi4FADwpoSVBZRqPJduN5kb3dAMYd269D
CmU9MLCkpp8BGoqvlK7sAbXetxUj5alnBmDEzuUX3v1whtGP98V+giAL/3MX9SUC
FXCFn93RW8ZlrexVZyX5URWkz1lrGxkxA6fZpmdaHuEQGoVUm45DydJfYEA8Fjku
wllVoHUTgOekFF57EdRTBusNGG3l3kHbZxoEDQyoBSDuvpqLZtxjR+JbPXwTV7Mm
CaLLBYG81X/2Re+Tnq9KCkgjzvOUPaMTGx/8GWsvZWDTalxvIIUdQ4ev5/5ccGVu
viuwpF4JzKl0Utm+odbcVQbaTD5oCF7ZCZ+E2tpdExHel1sEc504JOowwj0+xQ74
DLr0If09qxhowvNhFtWjuwq75zAWJU1wWGoCl2fetfcEbfRrsyIbD2RRRYbH9lwA
ArKCvU9+0uQusOICO29D3Frn7Vh1WhCGTFbeKRpzf9helk+Y2iwj2DF9Jzbr4Kes
X+GPxJJdHeFRSA2KYK58LxDMACazFIS6GiOpBHVIrlotnTM+h2dVZiTUCYrY9YyJ
7lQzymJxsrgci3RE+K5GjvINuZeTyDbvq0TXx6tRZHq8YNnPUscmEncBQ0//fkyt
HOPWdoEYo4tA7DQTbehhU/ciaAQDAq4kJhIpxx01zWFhKYDpVMFLkJ93J/aqm/kh
VPPp2DBbJSj0LHgxTbZMr+IwGBAflHk1I9B7rVc6lrFrAm+QQv2r5LnH98hIzbil
CW4px8R87Tb53dxkOiDN7a6HLV0rHT/KTfXR36a3a6qq5ST5MU9T5rOtqOHsWY5f
djHkKteic4Ia5j7OAlmDC3ieGlO4HwpyPuAVgKiTaUZC89gW6kfsIOZmJCdz0CIx
tTN49KlcgRbgzpPvCTme7XCSTZuIYo2yhqSZHGYAigh/jAEhDYYC3tSqvvWS8zYx
HFR39jcVqOBMDitHBIayhUjKHu/odZXz+mxGfCLorcaTElMMxvJqQoTg5jUIPZ6q
hBYnlE+6kj1pq8Bs6C2kJmWr/0jFNQs51gnkL3ym1fjLsYNKwmlhVD+V1mbT6W63
aGA4nv0e3q5gCm/gJgb15WKUVrt8K9AlP96PxizHFTVRq9EzUi3TYdG0Kh42GXpr
bGDFtiEwCd2pNwA5kqMvF3qFoCqdwntjTxf47MTUEuuuuEvofH9CY9ijeo53uRsO
u1fXEJQwvP6kKmuOx3Yj8kWOt6bmUo2PQByiT8y9uDIzrEeS8Po659kEjS1afIRS
JXq/KXFw3bdieU4jEYkkmMSVhloHfSy9kDZevO4uQeh9aUfIcNnPALmBtdKjQoex
1iqTkTzWGcaj0M7CvrAcSEXnY3OMquvFHtA4gi9eouJYDGn0+4FQGk9vnj99fK9S
PRWpWit0ScQyfahbyIm0OG52G9XzYfoVGj6vLKQQ3jeUB6BQjMQqVZuTN+mVuLE2
SmerZeE+Zmqxxmw+l8j3FX1gX8jvaIr33hSyEJU8ZD9TcMKiZaySH5loL7IV2WgT
Zau43PdrnlSYK0dpuJnq8HM21ZTuPLEDRL5UB+q0hTCSB32VbDJWx7+jlKGDd+te
z8LkN+v3FRncVoYOAxvpIvim/ACv1uKW965O4a4tdsFAwzpAxePMvspBNW/2kM3/
R4ExC7gIUqHmio43jvvSpMEoL35cykUCpSlhlDUJjPA9Mo3XFS/G/5bwYbb0qz81
IJNsBXBclLAhwh7u5F7Ngux2yBr93uGnYeJMOK7JDNjQIatK9apc+/pYoK9e6b+3
lSmW22gh5ee2wsLj8262vKo1JM6/HUebuAP4d7b0HyYBy9qVEIZU8uX0mbb3WNSS
rDvj/MxuUvL+QDsM3bLHTXSPLLBH4XRD41aKulQS4tldfJsAyUFk68hkVRrHG0gR
khXfyh7hTE/rgS8APIvv0Ap2gjXGbrhQjhGq83/0IO0m250csH4LKRMPA6tkVdhq
Y6yC45kmY4hvij1sD13Xb6dXzWD8jWDMMpBKJbi7g72NrwVInXtfeEFgha2SCzol
8L9Jq+X8UsjHrnUcS7GJxSlhRtos7tLY9bGv//DDLLOcc9Mq930o8a+3n/bzK6Vi
pvZ3LOEmppnLz0op19CO7QetEIrgwf8fWbiPnckrIx77WXnOsxq5DtFvTYHe/jJH
4TG6+tbSFwp0KFu0oH0KwgDwN/IECQ7A8Ug+Ut6U+MRZy3VGiiUP4fKf5uiU37BN
/q8D7aRtN0doNYJ5S9btUKZIGrAtH2XhSvQFWcJhRxKQ9P903MWDyxIE2ZOllgC3
0la/EEwlQgFoFUY6h2+bXH3PH/dLMWMYAzUBbwAURbgAPyxQ1WqO/WZGaLtcCS/w
aCrxpiiS502Xjom0I65SbWRTeYUPnzrDRS8uMdAzBeA80gHVdN8SG5qJOg0k/hAe
3Gma5q76ICysUvLvxMhOOlt4KpbNX3vFSSdmkK2O2gi21Q2n3bXlK5OJjllXD8+6
7xRgi9TkeM1mwptBXoTP6aQv463Em8TUevfqXY6vKaX/s5j+JSaCverL5jar8UKb
DGXzTuYwzKmKWcPkBaYFH7j5T/5wEVyENq+I2Nf0YSZX3ecBl+e+56SsvxjvrRXZ
UBDeXRpY2kBKgG7W1SZ0v+y1eSDDVKsiSANENKhtBYqn80Dw7gemcQmtJ5OpGJK3
l9S0S3ogDjWgSX0vh+g9EWnHqjbvajC6aU76HM+hNaKmqcHg5pII2PZqhG1OQmIm
Qw3accP3B+iwMjwV7zuJslXz+B4MAHuLTLLITmk5rl62ARestIZdFTny71zowpVC
HygTw9Kv3itvxRcg7Cf3lLimZMee2Elj1RCGtwI5KYSSgf6Hjew6uffOnTMB/Em9
OBnSGF45G/eTcsDND2U/y5Pa/+bVJpq9HCOW/FTVUQC6ZsFOV8o5sozYr2kXW1YN
AXXgy62byManWYV0mzbwCu1QGrb1KByezMbwfdZJE+VBa2xmzOI1Tmvp9qQCvcZY
191VWbBmnV0AGRwMofR0jinHijKgCdRmWyQX1fNrYEkd54dGvWNQuDC9gE5UHpkR
jV5MRFpCca7bZInW6YohY/2ycz3VB35bBZ7DOMQTYh+i16uxhJ509QvMbR/I/pBx
S4qNgQ3wkAVXufo+HKpNvxO05/xFcOYPnE0+j18FRlqAE+nXjTfaB3GcYXboZYR/
OvyrpmqS6BeM5ySDnhyN6lYBzgAtcPcq5JO+Q//efNW/ayCY/UJRA/6Ua5VT5LDI
YL3Y/L2oAJPop0raQksqTkkvD5acOQDN881Psxe6mKRW77IVvnl1ikhQ4AwPPxtk
AJGNVYjCpim1qL41fkA1X5vcT/ro6DVT5NlmA2IkNNVocYtkOcU5Tx/RpF9hZbhj
k3q2b7S1wENF75xKRUWVfKwfBeASOXtg+Yq8VxxS2AlTcVssv9kvyl1ootSg3GpX
WaYc+B64M6q1bVJ0X7tMsbGw2ERLJvSJ9oBOlSuvht+S4AAc3jHb5PR/aQUZTfu0
1xQA9LRhPNklbZsrIvbYKQF09ywc4tP0y/2zHz6oH517XYkNDQhoPxuy9XSrud/q
Np+1bhYC0l0cXgPqOqWTLorlKgo65/hAxEi29Aqit8/hGEmoNokHDFTg6q2Zv22q
l1Yg1THFwfYBAs5f3Xu958Cz/0GIr2W9qlPMwffclYC4lR/OZUrJs/mHdswmjpPI
1UR6OsMVmdN+QqPH8/PBcn0MaMWRC+g4+ZMMr7yJAN/UOmW/YYbfYcAiK4cCeFnx
w/Z4P4sd1UOADRQkMy3EpxgB4x4VIzHvm5I0Bz2DaqysT1zKQnwoHQ1NHtPPn1eK
lBw3vpWhCgohdL0Ty0kCHXvybpc1d/t18nS+7etwyRIJYa1E+yKm8MUe8xVa4WRe
dj892aDrHjexeHWQhqkRvMFIZrH62rd+nk64pg+zyRpLTj6YARqBG1aRIz2FX5CT
SuFGHP5Oa7LqZeARLTzh3jcKCSORLUdbC9pRthlFhgAat5NwkOz99VEcsn4kHHb9
xkosG7BwsTUWn5fRLPb9Ai1XE1JX2mUMqGHjy6RlW7Z8UGgfgSyxLfAbk5EJoVR0
+Lp18xHJt1HOIF61gjg7Tn60QjxlcHreH9RgdyjYeD2gWV4jo0WE0O/F2bR8JbL0
xlALvpyRwEDUeppQueg7YXYRvVl9VUDIs+VOd+n+RS6KrK44wGEbEPrefUh0n6LX
TqdwgeQCv5aW/vWgVFvnMwrlF2s2x4mIVPuCn/43iZmiuJ4M5YRvBudMpqsNYMIn
If5W9myx1s0Wbd7ZaoFm4V8roJ3kZcW+7qzc5PAZkVNVY3f1oOXU5FuUSI1MBbTl
wYgTi8fGL+MIXiliQKjyE19XsRdcxFliBFudXb6bPVLiwkPB71M6j83LvW0djdfL
WXVyRjvFdldZsI6vwTrUOxUkFtBRSyOz+naS3sFqIghxXOCBcNMo12PBdDfVpA+3
08JGva8WGQ6Ld+LLCtZPmN+d+ChMEYaiSmMRW4CQ3CQIx7Yqi7ZUV3ny6DGZ5Na3
8/3X2ekq5/Tp6Z+IYrqRYbFaJPsPSQHTaa14fsqtjvreN0O+PDiqSo/8NRlwGrU0
a30imFXKJs50cMhT9ZFWqcL59bSpYQhmPfJ1lHjPLFGRJ+f9JqzZ/j2+LPX8P4Dw
pRQoCOF9b1JenpkBSwBnwYNQJh2BWZzb1mE1hNyfHKkC6oUioWNhtxI+XAm7iync
1bjGXi6d7cejI41PiTPDniaALNY7bmYeYXSJ6M7Hue/Xlc1bs6kSr2GN0iVfoC58
DvwQeurJZ7XtRtVH8iaMwPihnHWjOm593Y9ZgwYIp/I5sy7d1mSsF/SZ/+KORiem
p+5AUJV6FoWi5fMvl2pJclVLxNWugaqmQ6X/y7GSypYYHHya4hCshoJ5vNnp5ifI
E1PE3BdyZzPX9GEY81Ax5LjMKWdCaZYhrlB2DYEO+1mQC3a6MMsvH4+O7qf/MDZi
oYPytWLqn5h5PwfYrU+vgNVJKi1Ydvb/6wAFU+7P1ITrDfl0VqsgLXcqUB9yKgT0
gpRiPCOqnE4DDYhIr5Mv12l26VxCdQvEqY1sT0/NS3KCMTL4t6ecc/hT7bdp1Io7
9JEr7S7fzigasHQQ/AL4DiD4yJeoVpqecUmebuOlYb9w0eepg9dFCf7is87j2vzg
Isl4i9co3GoQPh7C3JHtpoth/c586hp7O0yurRV0E9dc0Z2iyuQw3PDfIQP42Lz5
ihnOzNkWvVbKPSkoA1NmaMDTu8C80YVEhkmGFPHvrLZfFaY5RsVDGv1aKtLnoZJ6
GLa5aanKwmRgPoHM42ooxJizmftYl1K3YI8j0XnLnqdUY3L0zdU8ELUKlhyj/3Hc
NXTpertnukNkRReeFCMgPhDztikelTOyc7k0/rswsu7+h0eDAKfBw4/N/8RbRVJ7
xHH8guXWVN/ShVOQZl6ddJS9tvBGnF756y2u/8kxnaNqb6IMJw9DdTVwU2JNcCwG
XyQegtBvOd7jdlkH26qmO09ltPn7JgGG3yEJrrL96uhWEKuPEeGWqKlJrd7FGYBf
JzLUoXp+umb7WzExx47bFRuwUBQpExJ3ttmju7ErgHHvUdu24UHR2XjlYzP5FyWf
qmrd18Ny5nXSkAYeb8cOCf6iPNlRn7NQwKa54vlp/uXDAJarBpZLUJGzWS+V4U80
GO7cHJQA1WVJCsGXABOyQ53PsQN35hGdm597FWjabuCzkEzZJtpkG9EVhEzwpAjc
UMwVEvaCuvkIBMKzsX5v85ti32qeTs199a2/4s9cjI6a0KuucRF/utgT4ff6GzLf
LFVxtS1qgYpYxCGPG+YhVdeGIZhheIzwnKJDO8gZjgGmqyYorzPiijqmlQI1lnnt
0IKlcnyRk2gSINuqGsTnx2BTBco+hzBbgyi8eza66wU6Anm1r2TdJuTMoOXUSWFS
vA+O5T87y9/Rc0IMbRMO76bhECm+rHM5Pm31iNjCsepwRkplepcF17Yxe3rVGasO
YOXRMLF8D08DOHdLZcwbLZ/mGnmFVpBjzk9C0s3pmWla2p/rbEvBRpNhSuDVsUhN
bA5eI5tJd5ezH7gdY4/BasgbMySor0pdbb0jspS1xd1UQZ+PVdKOEIXflTVVt9Jx
Q5O3T71SOnh0S1fjNj5jeAmTBYuifUwP3Y7VNNoyg7mEzgpBxbbqLnO6mhfh3IX6
OI7nCEc+PSYiLVi3CCZgIhc+q6fZ4Lax7yX4MMuv1i0JHNyP0vvxi0AoxvkgsEpq
ACS6/uOkcw20qQRYENqaPuCcD41iqmv7RtaxqAy0JfFWNCm4vLErD3m0TpKz5SNa
1lK3O7O04xLlHn0/obKApKCNqR0c4uGJTjMdy21QLaTF1+irFecGfRJcTir26KMc
VPSBjmDaFtF+nYiYxlWrxVTnrWhVb8XNn4kiLYI6oRqs51MYSZI5OjXn/NKLVXJR
u11a/76cy5CZGrLchgbFrZyCHw9bJO79Vc1s02hwnTx9Cfu5D1rYQZ8iL3dEo+Gc
ZeOivm1faLovW0PmLeiE3jD9hVipnN5Ct4whc9tUzHkhUIQfTVXay7zlWEeZZj4Q
t3O51BAXb4nk4fOBf0Zn7HOwWU128yAE08qEY6Og2XiBBe68DIlWu17i+CuEXTdi
w+m5rrKhThIVOZJupCei/MyT/AMqSTe7Ta62TA/wKlA7SCCEwsrKY0SnTSqiVX93
jyD1SOZjJB7bALFiLQi/aPM/gg6FVqqxBtkdDECLMXIDTsjjWlSHsLZoou03+1jY
2ZKqmwEP57uHyjBEeWkzxcXVPh5o0Oz5owrovyc8XmToxVrhQRGjv5DkbfxJd2B9
I2dDtvdddmrH7m85CVjfa0+JPLosYHTaM9FEXQ5Wo2mzBufwrYwdKHFYJ6n574sw
9OtgRq2cVYbktZfoS5oNAux2lJK8L4V1j+P/1cMsjMzCA3HDNmetXN67HmCuxi0T
5s8e2mKHfTVCFBxjDbCoERC1N5fOmiW2BFejff1iZ/vMsoBIUHnA8pdZJNn1hXa4
Z4M0lasjRffhm6DVc2lgiKC+06btY1Ip8RUq5emQSowOjKxJes6ll67q8KlVrx1o
A/s1+uEVRVz3/pMmB68mYQ3ZoWpj1aCEXC6odexdQokxX4C+Ff0hmLkmOH6RQtm8
RLgS6kW7hjGIbzT4om0Cqfi2lO9E9grY8qfZKY1IM8IrCqpqPRCJnnCdH93yYVTT
kcDH47ULnA/h2WVgSMSLionzoHEM7PZqTu9p91vuEAAjsBBrKcTJ2/2cp0Qs0WNc
X+EpsSPne4UM+UIJP14T9ScM8dFHpN6V/naizz7y/BfXbpHqt9bLatTXGMkCh+BP
Tn//q/Mn1O6cwesK/1vlCEDANHR4/MT5EATa8qGUuIExTjDWoqCY0/k3i9hlzmW/
865SiwIB/LCq+KYLgDZJFed8273AgvryzLkWSAMbQbhBH32u2hlRkEvtR13sJqBh
lf7vGrs2XhMqNgASrI5X/h9YH4orZOj2jSWfmVlQO3+TBxFFF49D5K5oVpekEQoL
TX8QWWhXHqIODT7bx3pHlELlnLaRotpWHP4dSxVJueMFXPUYk0Khrx+PZ1lcJd77
JuJQcFKp25UOn+NxgnpJiEXOI4VX+Po/jHfelXhPfl50Pc6iM92cvsy+J3+8aPYV
eFcVUK74I4qIM4Tlx4TsPVkuHCMEFne9bPSbJJl9BdpQAM/EVwgtJyRfROykcJND
jZv++1psCJCDQoKjlD6gLNB6F2Wt5sa9oRn+uTEBsQgswxGXnbRlsQq25DjStaHB
iclkM7OniKlk/FE30exJ67+m12ToigpB3dnOp0QQY9B/b4tebfFPhrjP0gCge0lF
ZZWonRStolmIHhD8oMPAu4bFcjkWhTpj7SZTuOhGXEg55ccEKfv3WTs3EACaAchW
UtAMXj7LOzfbc6kMIRUtOZ/OOqCyLC1nTH+6C9vxK5Uxno4ITU+KwOZFOzslHh2U
+L3pT68JaV1IuIWZeB9snoSASK2VDno+beXNtDClLYo6fmtNImV4xbYhzAV60k+K
mYc/Lt1DNlIDn4WWBgg4IKmhP5ofLO3dPZLnrpPTcyfeXGv+xRysyl3Uh7mrID3C
85iPOWYYTm0bFeHi0MHZQWuKzrt1BbABC9n9dnn1A32IqSyHv/iCz/qodpv9AMnV
l8sJCQmV3ZPvzyCUQcc+iwXMNPPHF2tzy4PRV61hZb5HpQbMtjsmxXbfYVDD/lX7
iMbgFuOmSbPDhoBhiakgdqp3riFb/S3o7qlw8f2AfMBbt+lTkZ+CgQK+rCIBJbKq
AG+RPHkqcAMPnGZmv3rJTLWxmGyt8cG7GlvfNmUPvIPTBVDkWcKMcLhFaOy96c4S
3IXj2+kkdu93n44JP/P3okXW4nRhBr5R58TISX9Mk9IoReo4UGj/qE1dXm0PqaAN
h2cFwmhZcir0h4+9RfRPR+E5lXpiFePGB5ho++tqxGuyR+tZvOBdxcbmYKI0Qcky
5VogqZlHgib+3xfBdoDr5G8fZZ1DIhd6WeQjOMfhzp634FRuQizs6ipMYjraOLQj
ZbUjXslLBUDkhMdCQ2vdnMe9A6zjK5rLMCi8llO4oKA99UeomkFnUVq7jfkFIl01
EdGJBOrP/LRUuzm5Xkcds0zJUNclYwU1XOIBX2OZEBNxPZZoNYJqEo16xQXSubze
z1ZOf0MNeeZCR9AjfVBZuQjKyWd6gpjvbZlJ397V4fZzhkSh/4Oe2+MHFdMB5Fjh
GbLk2uBk1I+gr7SbShARJyShdGEqutiFMV9AUxMIqks/V/EJ9o8v5sF1WHSgpXMl
eEFLyurW7cMZ0vXUNd9wVkvM6dl6z4EcpHOf7sHoT4h2gA7pIYRCJS7dv7VyRcpJ
smsnvg2p1nMJUOH3QMw1XMcYK7YvlPu3HOWWUk2Lz5i6zvrJ9qTW2jg1wpwHoM1M
Tnk+xPN3TqqJP5PDxSkdUB9IetMNzaYfC7XbLT8/4oHgezdLBL+wGAtbdtTu1J90
mZlfBKg1C6rsviFTKhkLaHhvpGrW7g7jJgbL2yoOOxR5/dg1e1n7hyL4g0h0DgjO
FXu7Mj4SCU3jJwLqE7iZ/A5bbFjYCkNk3NlTWbOyPRiizkNzusO6M/7GfsDn/KAC
zPpc1Kw/IU3/goy3XCcbJS0p8JhdYS2kttmRitK44TYoJzBmuvoh6KwmFc8IudA2
ZJD/QN7z7oLPtFNDddYTEeuxicMvgKEq3lGUo4h90Hb7hF95n2tZ/oxJKgDlj/OT
MCkQ45mRgkEdwKMAZ+mMOb9J9OgJ/XHZiHP1kNKbJIrp9O8XaaLhhl2EDiHnyQ9p
fKk2mzVzu0nod0S/IBTOCKU/9zOw8mO4J3u/Xx1tSqLtSHkYhFP2+an4JWen/kk6
H+d4/WfwGwi0lBEpPPNOJWszqnhlWPK3Kt+PZRfFXbo3EMj2dhUSBGTGkOidT9Jy
9h8XAOLHpTE6piDcJSVpV5M8kz3AXHN94p+kkvETyIaTeQAEYUHZiihbhAOZIhZj
SFuiD8cy9GcYuf47eW9SFOJVYA7Hfs2LgsaycZ9dxk5C1ElaJKpb5y3NL/MAq0g7
Ld7vC+4NiQfwShVvoYiA0BkfmP3zE9r+e9fjrgHzDBV0Ni+sECY5WNln0Vg+yrs/
un+69W7suo+9ta+KAXaXW4K8xKvDWrYQU0ueXPvT76idSrriJ+4DFASSUCs/KWLZ
BJ6+KV3dX20CqSpIWBBjwTlBTCGXzXgkt6uyxSMme2O7gJq17peUuNNuFif+yxfS
2Jvb/UlxtCM81RB9znUMUr/H/kzhru1MVGsAI4V+93Z2Wj5B/821r05RBc/ddsPT
YxKG1xN1CTX3jUSWcAeN5RZsQ/kOcDOidCb0Jl8lMrF0McXlZMD/7x4M+/Qm+2fj
hDuKf2LJGN/5B0FsAC0zgjluxkjZb0mOhtjLjnfCA1UWap2PBI4WY36hJPoKJhfD
dbW7jz3/qvaRuSrQy+tra1SuGi15rmTB3FIWdQmKpWR7wVrA+uwVaiEHomKILitb
e7MGz3XpIuqoS3ZTS7fRVOqyJbpmZvsiB0bX0m46I/P3Rxl8COOLszGZwLRN4bCU
JUNNEfgzcR/j1zhuel5VETCtw6Ivwarg6aZE0KtzOgFGtvQNvz/wJsF9nDC220t7
EL3sCYordrjS0F4iKjsxcYslUEtvnWzWtmmoWLQ6YTarnYnUHptNaLvs8BHvYv8d
pw0tSKkOcg1q3oDYTAZMM+1e2e3TL/RYOMo2GEpIxwz+v7ymLs1IPlvcBttFPGLr
271h1uGzbiw+My9sKYyjWvazMxqdoMmvL3KYUMXQFmswbSY3sa5B9jZz+qb/9bCx
xQv/mnWaFqmSh8gv6bWeQEuTdAEKX/d9W4t84qs1cTa3imowF9stMHICTmgJI+6w
eC+6t/r9wYIyP12PaaOAY5LblQqnaoiaWGo6GzzaTgiAWi70J0qcaeTXHj89Bsnm
fSa59hacySDebJmnU2QXESD8l3QE0m8nMoUCgLDlhmlmzbAu7Vjx+IFsHN28JE8t
l6XLig8CQSYrqspEaNaRQWrgPA+DYCHGS1FLgvXt+XAZY9y4CaGxH0vUMPf9ufa8
TVlUlkColO4PGpgnuGHFsuMYOOck9PobcF/wnmw8ctDtltSz+h1H2W0S2IIY7z1O
lleB8lZcSbjH1CNxuViYb5D+S/Mg82q5dE2XxYKjc9VclE0Yd6gYi2RlqymzYdKx
e2fl2l06lVh1wj+T/lgAwdlgsTz1EDp4MzV2GSyHZMf97ECjHnisnOONO+yWb+Va
4ur7xlcft1vEQo0cz+7d1tO9m+wh96bTrEFOukNvAVitHsTUBL/+kHZHVw458voO
L58MUwx0tFRWifHpxIGjcalXiUGSnBW0SSOk606Ub8ywS0W5kwbLQUCYC84yvGW0
PJycZis+axzRfXIZAjM0mIVJlPU0D/vN64IAikXCpJLKdKqOuyQ+0Qo/3u/6Kuqo
3RogeQQJ/JQcYh4p3jVK0YycOg1wKzrcexBR5YS+ZOqsXwn8OGVDsBPwNo+BeiN9
4r7lzCHkh5IM6/pOz447kg2s31oH43x8oUyyJqw/Wge8/1hUD+0wcmdb+BLdwzJk
5p9G7bZKIIa+khtH0kt+T2a8XJLoTw924IGXvQuC8HbmMJa5/XPB1eZpvZAUIhJ8
SNIgefqXiG8bBxfMFMmMAaVosVUwBTszYsjta6Hx2QbHqzuG28bCBeL27H1MQwCi
ls5XfJh5YkLkvJc2/+fc+cya0EDlDh8n0C8xZmk/wMPu0NET8gqU4JaGsKG/LlLe
QpTpstx8nFct7DrTptbxTLsFZaSh+5WIBvVjn8K6EbXm0FPpwQc6ios1dfaS6ele
NnG/weoJYuUApnD4xKWsnk005Kr3iLoglPUZL+gWvcG3LeDzfKM/3cOsneOKfA2l
zQhtLlzZ1wsVavnOHIJd499jJS/SQ2jahIRebjY1C8Jdu8hJK3jCRwkUyLfLFE7W
12PXRdjNff0gFoe+91VIjfm95MFGLIHqwYx+rz/a3by+kHij2w9qqyVcqGaVcYxM
tFzm/33t1jjowjvdTGpOVTNLtw1XxIf+kshRgqiIJvu3QE59VsymxezfISeS1+IM
XH63A9nFZv3Ab+vnbv8IwFGKSEtwzp6oA5b3LY48eGFMHAOUYKXT30hb6shktq1k
ztHqjanbenn6C6ounY5m3Rw9TQP1kCSQKAvce9pkNowHfg/nFRajmZPxKubCxHKT
Ph/JEc6937EGRI/FsNZfOtsXYtsAogh4+vg6en59DbPUXgSl/7yHzMcCkw7HT7sh
kXqYYVfQ5bETrXoRKEN02qbb91IDQGdSbPaDMFskgFmTFYqNQ67T1pdChisVRcDA
DScmfCgI2Y6emHYSQfu5EjqXCEMXouK2wcqZV0e2tBbMZMV5rPDDshgdq7aVPuDD
QGl/pRs8fyL21mlHQThSA5jOPFGn3Z/VM3mR5liZJ6ZalEmsxar3JO9/KSkiElTj
EcOJU8HQDd0F7z+edLErqVIG9WY8MGkV8NuN3mYLVGrltSQrJvxQltyKN3v2gFdq
lpiL1WRxJhQuh8sn7EUvp47oIdc5Aw1zoSElvbIE0LOg8e+XQaquONS8Y271qld2
Zk8fYsOyCMACWG5pVf8RRMIOhkhZhcOH4/PdxRQOcrqCEyX22Hrbf5dH4jQP+bV6
UlbaLdicOhPZxgqGEzqAqNedH8xUR9ASm+V/YOKToP1K5lD+tMbB8VqxOhh66AdV
avRUnd3Mt3BcdUyP6lshwS+5n0Gt53vOo8Ig2VkAi6BPZEyH0pti3vQfy1dv9t1/
6lRQvE/GwjWUHrUGTlnBJZPbKQB5W+MbabaHs46t8y6MV6JHnLsL9UJLXnT5xZvI
yYV3M8JtEkJxbRL4f7x17Y2eTQeGycSa9mRfHtbXEhuxRFCYF6PzhoFXKuuSc7EJ
NrLkUjQcsizm6YacQsQm7imIynw6izE0QjmvLwy/ks6xI2g/2oLzqz14AA9sVvuu
kt1JSGwZSWpuwZGbrvC2H2bPuLUksRSynGhoPojGSnPlZ9qkKOYcTeOToOFstR6z
eNcHd2nsoyE2mTu9F9DPVnzqnIQ0dJO52PMweiVEBm4uqpmmAgxDkfwvor024cI/
XoUGG7KR600BaZEx4ZiC7lTXiRSpMGg2aNtxP4o1uSgnB2lr741Tk88d/9H9LTD9
St2PchGK1Y7TZmFZrynDev26npgckYncULwtYfBKd6lw9P14lIuCwCngaNl2g2UD
AYKcoloQojgSzJmriSyrBvbo+domMRVpJPxzVvKehZr+jPWuVzvsk3d2UX9yW6M6
BBtx+osRhWRn4L6dUf3cGYnL/tDnB90egliYN7xkyG3uJey2yVqcG+HDUjDioc20
133kaVH84LeT2HG2N9gMlCy0W8r1zjW+rGHxhCO0DBz3V1if9KZY95GuQeppwtIf
jgiaqYJnWIgZ9hGALsFhusjy3G0YiaIJZsHs6z+OUOrW//7ZUYct9OGXrO7Wi/x7
F2ZLgFclM6MIIdSjR3u9mtmCih1foSzVUqLb9i5IcInympknLTFHmPCdQoT3yv30
QMGZDK2GW8+wQ4o8UmOFkgtPCe0hDzs8S+DYtcB1dM9ec+/IPKN/GG8/xN+96EAI
HuXnfVtHCGXKEuFHHgyHLaKTm11010GNPQd/LjZtpL4hGDOg1hROUBzQ3Erq3Bjt
K5hx26Mwwy7BVnyKChnHpfHL7dDKyRx0/8ywBfjzJNRz/VhSmkr4hhhaT2C/pO+s
lP1Kz/2zcPZIY9NiyUujG8Vu2u9keCmUD7Epe+po74e7+C27fq3GHzxQ3qe528WU
bHMtcOo0NP1AMGBn8hHB31Kbv4lEterDu49Ahw0JL+RLA1KSX2KkQdo0Wz874imd
iTAtG67U1N4iYcBVTn1DUDyp3jaPHqad2CpAfhTYzOL81bsw8mARW1eM4ntTC1us
SQyB92rv3hNJMQsUF+XqBWjS1Vb5zVERZxSmszcL5S6WAt8OxOcnnHBEQWuXkiqe
sU2ltKZtbooStpPKAluiyKCiTJ2YBTRoD7nGt1pKne6Gnp9ifjL77EVOlPpsJHIl
Y30SHR1See16GDhUqaRp5to9gQBMtBzTnG03iM8OGd8wMEIs1Zyf8N1a3/fVE5U9
2Cr6flJ0CS1BVj24fxThNSenWW35BGhG/5JRHu6UQ5sQ9SVQLndBuarV1GnheVPa
oFa7Uohisk4rodmxh2sfXyuSEpRh3WJQJiYaeKG0IcZfe7E/7iLlmj+Iaa9F2KQj
bF/pRHcnMYQuKqN1tuRuaP1PZAUg9nKLdw3hCQp1K1wAUajkqAuIDPY6j8Z72haq
g+NFiefmS9rTcXfPGZ6NVxto6cWRsIH7HTLGh2diqOmknQ4LZDbnlB+ZlGr214Xn
4Q2/7adR7c+jyRu+aQEURdXnSZK0o7PafPaYGfmAw1FK9ecnbDm7BHkOIv+SMkSr
VPf4qYNnT/cunZs5vF3afqeqo7PVBGTbAfQxhWflDZa4D6cpQRU5SRZ82DRVwyGg
tgaqqAVP1BETSVOrp124/P2NsmuPmb7UvtWCifUGqidmFfLg8XX2V5ewks9lWa3b
ufAPEah7kE/Xexb9IorERjTCR62efj9gQAl3Q7fp35T0iKde/3JBxBlMwHYu0o4L
wa1MTXjBxNFvgqiuASK05JmAIRj55cXSGFJzK19vhvVGsbHqn742XTqm5AH/KdVd
hW/E/c8JANfPOOlTaLwqDKpV31r6aiVYzd1nfjauhnhUsRjz+iEEYGNDfBgPOQAI
lRwZtLkK8dSrlrbpDnsteWpyay7UqMiKNdb+/RMIcQr1bNCtL2lSd25ywJJm4hHv
e149z0M1QqMVWlO4OQNM/14hzk5kIpp/CW3I2PUkPZWh3yPptusb0xEpRKghgA6y
i3K4l/X0RQZJDHitRJIzVupwrvombAYQccSZsDtPJ1MT40yhPOFbq/4MoHckn81A
E/LuqXqFAPm5JAOkKyzjjwGicgS+4HNCYHLMJ4S4dfEyzFvivo8+7ryeKUaIHasN
UWel/CdUoyD4B5aNQniLEUq7Gcvwoc6MyM7YYkIIALyz+YiPxcCICcsQoiAH3dXb
WTilKHB6/4bGQhQCESsJXYoomSJy75+VWUrII99KlK4pyFxt98adM3XpxOghzS7b
tl6Hl0Qabn8DVMV9cvZ9MpWUUZJBktb5pX1QBZU5a7fIaymBEusDnQRww7Ra7xWB
jJ+DFgGATAZjnEIyDcqzFfGq75sdiUROqH3iVlkXPd4rChPzmsmrdbNocP8EoGIM
+tJy6ZX374s0K5lfz+3ZWvd6ngVKmGUDMHx1a/AnNE9zaGdu/Vdn4GRci2ChMUxO
D5Jwvcg2YVwrZBPDpPerR6dZOd1vZD8zKer3mNSX1ItQZCdWK+5fZschno09hSW8
VhZU5veEx/ymLlhoc/PVUjBFeNXDCbfJb0AqmWOXRNFYZKIM6x+Ym9Ur5FgVyExy
1GkW9A6zA5PfdZWv/YQVrFsCaAiJ1Q7Pb6ZFE9e7zNWYAaBDY30Bmrr7CKOIUSFP
aCkXo3R8Qs+R0qQP+bdIOL9atcdawleKN92Rdz9ratEI6ybQESyMG/5asxFD/RpJ
hcT3Hs9rqVV4STqytyZ2kjjvbxKJmsH2+cZ01V466k1TnFk4XVTvx6At6XZbwf7B
9vVZvU6CzxC57qDU6VvIIVpNIqKejRknd/trbNWlaoW8VxH0LjKb3rS38SFjOb5s
5z1sQZ0JtucO08OKtdXGhDxnfS4Suvq/vEbzQhlDncO7IGRmG0hfy0yucjGsyEkr
S4QWVvC6+8KRTTMz/scCcnA6NKA8jMvdSYMMQiVv11EOyZ4DkIZB7Z6JQKYkRNHU
KIP1Ytzg1uNX/Gjds13FXaizNzO+BPOMXFHAr6VkFKbb8YtQvd8KxvDwoH5O3jmI
SHI1P+KlhKtQbPRjRd1j8QTOPbOJtkS6XxAzfODmXjcyAFXOIgz32f9EKKbFKowJ
Q3dIuKfyH02TPKpoB75NRqHOSZEDFJZTmEjfDfJYplfUrMzS+A+bby27EsrCzQLB
G1K94YfF4DZAKg9y9UxOLXWYzau82ZvaWMeF6icSnoWylq6G5ILIfQNBKT6rbwxm
ZfN8bfdmni/8ckyA8ipAjtGiiUo9M9QnloNE2fhyrZUSDkkzZEPRxoEPsMZpbBnR
nuZaydnqQy/XWVwjmeP3LMyIO6LvW/d+3iE8wBqvAZIqt1uTy6xvUtcRvmnjzw9D
+0qvzzGUPkhYJsTUwGg27CxSENL/aqT30dNkDq7OImIH0ugNPlSZp8KnF6XPs40D
mL6jnC0kOuQklwriJ7OBbj5sISZqVBzB8YmuRQwwVGnGl5TrDfoA4hrtwDfJ1dFQ
+PxumkCwStrAWHbWoT1HqTkztS/L1r4+HKpxpWzqz0IXq/sUgWhc8wuq8p4GdCij
UOXmgjpSWXvYGRZJ+5MVa595kt75YsLWDqjwkMGDn1M0re0LqB3k1RjxyfksDxlk
OC+nExv/u7WxigmJFL+Nc4A9JsDvd6KGFhedIEAe7/wM1Z7NHpdUv5NHLNmwBLMJ
xk8INjcon9fwdXWcTOt43avMZp3xoXkAZPRuo3G6akcKgKcNpwWgOdbI2g2Lv1jN
QuJgs6Pi9cqNjjO2tS7P5sjpgehQ3w1bO/1+LmLjynhOZCFLxvv6uvZlTtv99ScA
5rtjUZfcXJZLNMvlJmGPq79zpj3HEiLxqY9H4taHMDr5L+NuEkR4b88/h2UT+SeG
KMslYH0CsEOCXW9lD0jai+b8BxFyAUjLtPLWWcpssK8fmtnMMHdPW8ygcrQ3wj0O
4+FvyMUwtl2OhnRtv5OK8JIqShJU4twlwA3sNUDJsTWO3ESzSgRInR9iu3D7nFgM
mIkis3B39EQb06SgDNct1PzaueHQoChwv2KFkoRE/i0GpA5lBLi0y+UqILx6I7ea
9tTwlZKx1zYgz/7NhDLwe1q0t4F1MHWUlbz9O6Yf4UM8taxofnGiiK9DMTlqne1W
4eo9VVyiYMja9/ALiWM+i3VqajH2S5T2kn2FKKzMTG3rPqxugDttuh7sRz+KQ3hL
hLmVO9/ARDBlCzujzRgrRxVNcVjmhAzmXEmmLKMJwEZCcyrTI6eeVZsmAB+B15dO
`pragma protect end_protected
