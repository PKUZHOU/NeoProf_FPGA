// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
BidGahDQY+Ni83BEi8Xi8Z/4NZd9cnDiZmeKZlYN5ptcFEiy9wm85k7P7qdxnQBkz8aKwiosJehf
uxcx/Ifj2rbe7tHfC2Gbzcg32ABcJV0vKP16P+n6rohyZ2BsuX3qC6iC3vjWlLD2opWZnhmCDnBI
yFIzHZGy89deZlNJwtNLNjTFLNfIHryzn/a7WviH55vRWL32OsKWaIQTtIUBm+D8dIv4wjsfUH7y
2l6Mq3Q2/zZ37mYuroPyBTSsA7opjNwcKJLyOQX7pEl4PeW0/ryacABL+3zlYpT+ylV1N8dpi/sH
4pTsNdTvaG9R5JcUdfZX8kcW22d7ZBSUjswclw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 28640)
jI4BUYgNByZKHiYik8n0CGq6hR6Yj8AoOC2UTuT2qZt7/twXBA7u5s+x6OMRZHnpaHYHLZla0z3o
UTdVYVrs9RTYyVPiIPUeFWXN+D0hFVqnXImNgb8wZKDZkgmdO36GMznVj+mjJr24gJcycWtJDVWI
Y+Wgy7eoXAkYRHAHYS4p1GiNPekRU9Nc2+l6mcSyNVgyLTxYBvvSfET+shNqrdw7mICe4nJ8xUqo
kt60caJkB5rAFSvdVxd7mesgcQ2pmN0UNyv6T03Y1jKMW3dRAQQdxWMj1k/aaXsVuP7EEDAbxj5c
GEARX8nyGY+ydnf2NFoduPMQHXEVHzt31GSz0WIy7RET/nvthuhRrmjL2Z0CYzbKfskPrmzAt8ev
uri3fSF+S26xcisyEEFM82aLxKQrntV8VZokisbnjEyNhrqOqgRGZoKbkSopUMPTYOGNDHiZ5CD5
1Y+qYLq15CkT6Kvie6oxIJkbhOJ45+ex71XRk/br91V6sge5gS8E87eyrSjgLE0exz1MNKswqXRA
qW+oI96TGndMY5PsfDR/TXD4qL8jyzS57drptTCBxFONojlSV0AdEv2lCM3xs7fsvJUd8nHS+wEz
BS9lMmqtqXtOLUAhPWLylfuSylzD6sm6oPZ/Z33JezZRyIspBuZtQEI1KVAGIqHFa5+TJWC524xL
+L3/3pvHtFBSG59iUhaqW7DjK+eot2k6VlfPpY8a0FulvPPeaV2ErGXP1XkNIadd65MFaURDzsZE
oUazUdMc1Q2ms64PI5xEJGZRjGlyHO02XtgZ8Bz0xZoaj2mUHX5TIRgbfxVJA/o9rbYkh29+aDN0
24I7PiXxmhsoYAgYd2Tu7fLQDqgQSCM3G+W/DTiW06rucFoTPJxvJ77v5jdjRJxDefNhjZ4FKIkB
5R9g7BhH+6wWQplYyCZ87O8zI/CamWFqkcSxM8o0MEYiD8QioKjTAZjwLKoqe3Rm5T0Xyv7fAHzi
YEaD0i/OXh8Q0Xo7hYB3xJK15/3v3FWlpk6wK93pNKjVSU1ThxJ83NfOKrlpbVrEbF9ys52Adw+/
mR7LkhDM2lNycy74WZVOgpoglDS+9NRavEFDjcvTxHYs/mRx3YMEPQlrIZM+/IxXPudrn7YLGC0r
RAkqkilrDnUbJLl7ih0X9i7/zbqQgKvKQqIjEAYyQCRTiqRxDhRdRqaqCc2DIv8LSEYQC2vgWlPa
EwVwSD0ZRLB7889Al2dQy5RG25em4QAKUIeRsLknNz1tTnPoh2EQOTQB3Z/Wyf9TuY7ypWhz9pux
d3HvInhL+ctvuNhZ5cIdIX4YoHZhJ/B0Fbg/DmSFmtkaUpJQ8DjdUnNZQiH3H7b2zGsAsQ1vUIys
3I3dSM44xdkly9EOlE/A5V/2SnjIhjbJ10+p9+K7HTBRFRiyRJd8VkzMqsanbE3s49ZGdFBmLV9U
EG6SFn0aW6FLpmeDuSZTXMYE0aLhznr8/QLk7IhEwwnIZbOavJxqZj2dNwxJUUpgFEC5YS+oQV9J
2KeeFvcK51yc20ZtJ3D16KSiTFolWnmLQ5qH513lmTFTLOudhGJP53pKgdlXb55KSZjRGvN23aZ6
E5CvKtrqv03goJioOMkvwjRrj/2slkWQ8235Ik4voTIsQNwvYaWOZvgUIv+1qJKi5kEeI/xQ5efU
YeyXSPI1XUMA+mJhcl4tokZH7XTE6OcgxDwa6kQ9Okp/oZ8alo3HufRtW2rt12WOcM/xhCnq3o8d
iaCLm531HrwGQr2TdBEgcaQ8tFdlh9+qnqb49o6e1D7Yrwhnvo7Yt9WrrfsJBEgCWA/QDwbrIefu
w5DQktpFE6TINJ+M3NJ6jELpScWrj0uaRkiTzdixAjBX7ulxgObcYVzNaAn4K79NK/uCb+taCrY8
XrgX1mKA07MDQmu4jUvfOxD/+UpCHHZDr3HkOjbO/J85JA/LAojSjnvKfmiOSqryVddlGOR3uT3C
I1tXqRRVDPHmm0k24/zbh0dqXbMuRfOg5RDQVmqxr0f5HNrIy7e0jWcBC6wZWNU8TiQe28tbszgk
5HJEtO3xMSEwsFe/qzMM4fYjrtHX1IuzCeeRYh6p1dAOuXWbqeYEp3kuWsQGptfQDbDjONMrb+KR
e60Sl77nx9tpA1R7sMB93UL0205Uv2tsGJ6O61DGl7H1gzSBvMJ2uBdOpArwbvKi3Fq57ch6mUw2
BQ//w1+1bPNXlDDF7ctESmAxgLicjTs/oxN778Nbo0soNYIxbxX6vLc5ob7CN5dPBGs376/keE1b
oUZEfMGT7WM7lmd7tBTNYpQWOCIHc+iQJGbtcL4NJ6b23Q6mAASqeDaXaC8l+OZj/ryO0k9MDypL
hT2MHMdXSOxc1Y4UzhAlFdr0azAjl5dNhWNt1E/sq54ZycDYnOXytDHATP+5o4RA2XO4VIGUMLvt
eivi1dJ09PB+dgyRn4UhBMKjcDt+SzmzbRx8MSMdC9wPBsOrw29tXHSpZzhDki+WjMd59wDQ7qzS
wW0maVdyVwpUlNuTSQWfNXwGnXjJLRT0Yo/0dp2/gYf5OG0e9S+zyQIlA2yraSmZM7M6gop7uWXI
26ocWUpZ68N9d2pVfda1pq8cj/3tMwY1DnaV0m6NDYvadGKFey2I1sVk+8FGoQ12vGpLS2ObGpnK
qSRN/82zUtF4IpuPP1wNs4bb0V4/2bSu6lUjvGPtgU9CvUvBq7YfQi7Wnh6r7CAJgDJ9l0sB2R8e
aX6J6FWspuSrkFYNTJ+T+1vVO+Gpb7MEiYNV8lc9GHJFQDUkJsvdAYxiv6uPCmEGxOxQP7rNNrcJ
DY7KnOPWkWwxsTpJhoruBdvSAXrBgtoMtKtrkOplf+hw2EXa6oZshJppjRwN3LFXUrM9CXs+Bk9U
R3CezE23kP/NA3FlL5EMWZzbMVv/qEbmg5EBXo8Q8VwBoPsoixvpi6LU+QcPl/5Q/ln6k8lQN+iU
g7ws7DUxywQlnZ48OUEu+6fkvOCyZEBtxJnIf2eGXOzPrWYYJ7OQcWY65HkidoZGwmq9L8iQ+g5k
WLASOPuwzrpEXDFK3MI4zK3dMIw4qY6+sX0NfoYQ3Qwz9mh7xgb/t2nlx9LXOxxOcfE+JNzDiSnr
nyLx7E8+zqrVf/gIhwi+Swe/V5wJY2r5gZLYXbGPEku1UWewTsxW2eX2TLz2nSnl/5LM9w2vzCdc
LIMGJn1J6q0Zt26R2rudWDpQ3aIYs1qxIra5rFFjIzEq2FM++pKDhmQTdqHEC8bsyZ1lJ7LFhYdY
20auW4bfY0Ahw6qOAxqqAOHye2QsDYiLjRJm36sQ9Rww/onIsytDy8ryNTNw+jIMhUhErSmK6MLN
kEqi60FzUj24nKwY/nMM21I2qc8Lv+CMUKAt/DUnuGYglZwo3cSXKhGy5wWKVUo5DsEsR+Ck4b66
JrR9nmKzDiTDzINj0r8kwJFZm4SfcL3FM1l0puKJ61iPdofD6oliBpSS6RBpTnOoFbF37CXYA3EO
3FOJIYo7kvo3/xkSW2eO+LkMiNCWWyJqDTnJYHaux8gLAD3PNfnTKoh4TxN0puC+A/1XoXKVq0k3
KWdCX4Hc2cTrCG1d4CVxr9x6mPI6ZmO8KDIecRTSEndLR+1L27DuGHPE7vk7Wjya9o7ikQ1RrxNu
WVduR0SIQYpiRdVSxJwfX6Yxpe4bJ+nRlT3GHxUPBR24wXRmX+bdnHhq69hFAAf57nYbtPx37IPC
v/oTXFo/sst/lUPDDwcw4SPBVN4Yg+drMh5Dd0UDM1wzSYvkYcP/nmNi4vi2L4/f5SgwUcwudTNJ
icVPPZY305lBhRHg7yaqMnYhsPIni16WOilIHgiStGXhvoDDkrURD+9DyCCimxs7I5Bv6vR56a2Y
VehN/9helGcnrSEIX9e/T8xFB3f3H1YmSUXvlNTPi9erdweHjIy2pdo4gV74vO6fr9Qm2ch5w/cC
coiGMDsDk7ej00r7Se3bUMVTiHdvyuASGYciFUPnC3KfA7V/Azw4thXqFL2HWoj+nMmShBdeWxq1
u7OjvIcnkO4DdFXuUjC6ymbis0VWo7yKZYCHsMQQs6enmSpp3K/1j/Llemyiw9J3hG4djvq8owNZ
TKK3n9VLzz6VDCxvtb80G080IJ1b4VjgBC9OxlnIbHX34qeR7KWN2l0KWgYdbG/1kWG41X1+ZgkV
4N5raVjzon0snzPT+PLcwnDwqnpzEuxtpDnSp95nERA1bBilEHyu6Y7eiwhU+IXqxeyuKL6dtoq1
vSb7IUOd3kYBqqfzK03P/FaiBKtoiNBDu5aRpDSkfn1tgPJ8iq533CCh2aSJYUeYVTE9xnLfsCso
4ZHDywJEz3Mhpl+cfinMclUv8+B2ScwD7idGHaVi5g5mfqkiLVkAPsO7vdEyaH/NeIhRARy3QnbX
Ij4PqCq6bW47F/rNSKRM7ZXlm7AWj9/DbJZXpEZrGKQAbjuIv3ZZUY17ZSn1sWrcLzKdAdI4L0NO
1G0gxuSDi/TImOfoCU/EFu3ZYYt+nEzUz5Cz2W/TeCVz1AMxDu3xVNl0SaKZ9ZajAtOOyIPwOEcG
6035aA6ioVyfVxFKbcUgfFiE4CjDGkePENSvf1mIY+v0R4avsx5S85XW2q6zXecGhCQbSLsMS6f0
VioOt1OYl6IjfmHsVwK5CMyERPOewRRW8aG4YxTm7+HA/v3jTFadfkjOdXQ8A44C1PW32HVyfqFB
+8o3xcQN4SeMECECcndYitnm1NDtuqJ5W8E3zeB5nB6PiTyfHlKmtZz9LUewfP1yzMitQUy/Lup2
5FaZ7hyR0nBAqPHRb703pnCgpN51+oivpoIBBghXdlJVcPc5nEhGrCqlN2TyqGvE3cMm+nY5+omo
DiBEJ0FHQbdxwR/epwCC3O5aviLX7iCVoDIP189HKfZJW6vUyPTmG5dhiBgG9Ur61qk/UV33uX/8
+sosNlGt/E5qGgPBl2GWbgXAMTWpjH45j4tg75Krrt/uaAu7rdHrOfDa9piVCTNknCigNpwv3AAk
iRBOTEGW4IkHcIvAA7Oby8L2yV6OgPhXco5rHY6LXME/IRAVO9FSqHRKtTGGydk/Oc0iQsSsFkKc
mROPHKBRpKs/mvD3vH4MxHZeRW1mJsRegJXQ2Gs5lKmAiKTLSGsF33FQrsUeWvmBfJx0pK70p4Ga
/svak6vlcGBnMfy49+SVBEPbGq76WamjADpqhRzf/CEX9EYA7r14xbCv9YJbNjfA6PME3TnuSc7V
RC3oHFbLu+lPcC5DZEZF9YpC7Yb7NBcl9YMBArTejgTVpJ+Fxnp+bRxwCajLppUcacJwBVurjgFN
J6mrntsSFqFqb3VkJ42uId/xJmeXSjvv2qBGkJRyAu+vSRF4dvm6bMr/ezw0VLfaI7sNUIUm/Jz4
GU+6iiUDG2oj1uG5ObQNp9/HYwl2F9OdTx3H2Gusny7ZLW2UJ3kikBT6q6k4N9sKooh87YHpQZdh
XTUcsaoSm2xJFu8lzXw20Rl92kbvLJ1jagg9FMWsPwqql0YePr+KVcoNOOO2S1lRvXMIuxtAcoI1
NuSkJiMpPTt2Jj5n9O6UWp6EsXNGrOBvVGOmqVa/WMRtRCL9EDAs5L3R7nvTs30eIsoEg4pVTGsD
lwpDJChLutS2ktisvWuQB5oyFcpTaK0rlmMOCOAGyWcSiMANqVfQiCch7ECunesVFWtmXLyj2oI8
3woNZUBXRc5iXuXdXA715PkS0Ea+/KkiMsRsQVbTY34AhSd4zYu7SrFf84iC13WK3NiVzqDUDdV1
wI7z+3MD1DrWJMUdHT9Ngz/WguRK8i04Vr4TSIUp3b7+FOgJH2UprttqifJuyUrKQhjB2IN+fHAZ
3Q6Lb6hjSFvgzPoGdH4D/QuUlv1+vYfR1OFhuJwNyjdBtHls18VmhBynkY1H/M8wRSHnpfKmviFH
YZs9ckq+aH7q2U6fKRwGuMt2zAByCQD+47FYdUF6YnCnIInTG+NNtiHJvr+Z2728DXvpzxFdsCkx
AxIwcG6TlGnPHIdwCKMRtNOySig52rR7b7g/47CcfMBVN0zMilpZCwngls7gKyWSuxXT6lmGQpwm
bNijjk/tFhFRisfjo3h0eiJupxyCenCTHdrrG3U30wv2+NIe6PvU4hQVP8jzVCQCttl6DNIgmths
/MnvT2d58eYohxfxrByC9kgdTmaWVps23GB9uhBDpmlwOnAbDjPxETl/z/xmL9tGf4GIIdsJDVjg
Ceb1vxOUSeCbIoc3/pnPZ6iLqOl/hj+QOB8ib8Ndoix70HImLyDFyiH6g2cw0PPCJKloHX2pWqrw
VlzE4bJ8pLIErP3gY+WwV2PnynXqAyYhMzJ/QcFyLHWZpVaQuGsb6OOns1/5ES30LVEmnMpLxbb9
BpCuRZ97Qd1QMwN/irFAT5KqswzXSOcQ6al4BMIAIIJxtCPIEvUZtS/tkMOvVUkFOzky/mBIisRt
suPN9Xu9GPdrdIMsK4v9asdnL+MVxvRrkojDoro+WKT4BI8LqyGcrIFXYSeVHcXWDU79EgpXIvuQ
tnq/fywHvY0NuHjHS/WkArH1H3GrmueVhB7LMl0JBR/qqtDBbkWe0gQef9q1o32RtatNLqTbw9V9
bvr1J4ED1hT5YZHesdc65OhnevYlj2yR0R1xtxGro2XbxJ3jvGm3RhjoaEF9h5NlyYIHzcutc65m
m1C+Kg60vtPryGk7y4y8xqd/KBv2vCsxgWYaATyggLsLmHlchRMVCzyx4SVSaiFZCEd7v4dJpITr
85Xn7f05RMfgGMX8DHUxc9jQ9Em+8T2xl9TlZgoBSU6rhWDkgT29Y943umpRw/n7g5Za2MfbWWDI
6f9mMBwkG9ZAZOxG7yLDXKuxuxLz+ib47pXWCRFQnMQivTHind3874Iy16rnq9e+pYDSllZsAfdq
IEzencfT7CIFM0NPQAl5pvGPkEq0oFDhRclE8cp/ZLLEjtlkp+6Gim8b4Cjdf64K8XjLKcU2PBm9
y0+11HQHiKXbfj8h8LZDWNZjxA+UtOxQRJ2sqOrNkKKob77uibWsNls9fnVW91itYHELnHPSBXBy
Oa8/0cGnzHwoEhpwG3LHXTIwsEiRyK1WrSsXk8WJzpJ4OdRYGY59C/ToCnS/LiEzb9X/42Cec1vk
Mngyjo5kmosVATzREFaD6Aai07kicWFe40PRjB4x/TSD9BcsYjqTAXlMQx94vw4bm8K+14zaSMBI
oT3A6an60n25q5Pbi81TMQ0mlU2+ahzsmfWe2gGY3jr8NY6i2TCa2nMEXL5S2+qjoRk6bk8+UzJ1
+3qMlFj+ZfsROxIDrCIK5SZpwoCFT/jyVsJBfETd+Fv5UxhSyqtJzfpbI1RtS9paXDzNT24gG+wc
fF9la7ItlMVnudNFS8VbRVxLklU+UKE158SrxF2JdAI5zAuojbumPionFai+hW0IZWr2KT81Gq+r
2uBQt+70eHJVGSG2gLJIUXPjQnapVzvP843ap/Y6C1MyRhHn4TsM082KkrbTWLsJwAXXvZIyj7vP
34IdDI0PEVVSTvrr1fsWrWDkLmNfVQct6g+UcvzYqvUZDQLgeaAjQcdNRqqY4mjV3mCIx0stoPi2
HLz321sGnzAZEpm88mbkySL4omaWTNKqey05gmv7uSdmArLl1inBAKp1Ji3HgDHNTka0BRjwN62w
Oj7UiP1dfjPOZuWM+t3wmZ30QIPkYA0/0dd95SC3DzGmj36Ol1aCSpc1otNzA85NFtV5RJm8q6MM
r8N9dcI46hrp+/IqCwX1agdDpRHxrkGax1Xg+eEUDVBhklJ3XzNhRuUFGR+GLHKYPJrzcs/Rd3yr
+A7mUlR4SX4x/w25CZ+DxV71ZBsfhRvSnD5yctIVMUGyyQFx3BSCHcPWamqKfIcC4uNe3dwRlGvu
Guev8kHNr+5gxJCfi7A/SCjz+hi+zsbplmDOTv3uV0+GGs9VSn8PBqQ7BPkRABh+4N06ymFceHkH
d0TAgQMVbZFEPM5BqR6nlamG40zm/mnghxjmBbS++A/JGv4EDj8Bav5RPY6W2SPYwghSNmb7W2WC
uXZ7ofQ9gcQJGYxuguXhm4SZEksEcGrRGMBd7kEPgEBLrui8gpGSsdt4dCACc5WSfW0PY1lBVeHJ
4VAJ80oS+jvKfiQ9NXLBkTjNVOw+WWzSfNu7SnCvfPrDZoGzcWOLDpK5Kou/w0+TNme4XyIHZVXm
EFsLo/nBL3EKTGr+xLlxnyfn6NKocI3ogh9aDah1DTKBwuLmoFDeQmv8rT5JlPlJSXzTpbX1iQcw
ArL/EtlVglHA13aCIUrJX4SfCe4cWjEAgyImGPyaO36kOW820hrIfrC0TXLfESxS48d3zf0aBwfB
+KxHGzX/nCl3z/1vWss8Py+hOkE93mXnZk8Zrq1E9vgLvsXlgAbnwcSRMV2ahf68SNbv0Y2l7xNR
tFEDQZMYWtGrZXfn7GzFHw7udiUDUAcdbXMIx5vigbQPhSGTn2zpAIpYKXZyyrPj2VbNK2Lft188
ffyV3ZYOUDnZExTegMxk87fszcWTUMuGhBl63AmkhBDEoWljOt4K1OfOmxgyCU46yfXxR/ODRCNI
eJP2IV1V0YTbGNxnZgpgsQ/XRckRIQn0u6af2SZB5/ful68iK1bJLfacozFFKgsTDKJf0hstne7Z
lk2qep4Wfdkl7GkO22ChHEE14FLELEziFlkv9g9gDerACSSwDqZNSqJnrfIQi0db7btbOxZYbXbQ
8y9uMIDDrrpNYt/AE57QWHuFKVjItk5s7uL1bXrWqlvr+3UnjPrqGtoWwgGxLb/grzrbo/SLM62S
taJquUQtazNxlcqo0/fyKzANNYwUmpreo/DF8DDnLhwVisyRxClROcwwGROXZQKhDu/0bXuQ42vz
n78sKDvpMetHvBb+SBQ4qfzdZiMT1vWh8QBSQHLgDKwieISp+y8VfGGcKvUeQLe7hsReZBPihcOY
IHTeA8dycu2rueG6SpcJEkI8DX0xJBuvDspBhidrmxc356FDUYOuQ5BtnTZyQ6P6Q6EV9rHIGN8x
yxu5/Xq3kwogOr8n3unooXuenzYhe7glYxp+0LWKrYGH9gJosJNVYiXmJIYz6Jf2Ihf4a181jPri
czJEPaCkr/F6SJ9tlSGDxaw9H/p8Ieoo/KLgJgxhj8j/lRhT8rewkMx4ETzWXFZW77SaJlhvXTlt
syr9MHdxc1QeSMm0wQAR2Pi6j8xuc1gL1uKQnG24uTCsACI4yN5O/skt09K2D2BRVOzAngYKXuHy
Z0sUEyMiegrpYjf0ykUV5GiZKu1LmJ2JsxOXwyYmxgU7RkV0FmBR5JkycEIJypT16IwriJunDD1x
3ckij1gZ3XU1g4obO/7bg0nSsw1JIXlyUUtTnz2TPfCCDf3l9Mxq7tLCnZHR0a5CUpcuLty4Qbv6
N8BmFlydNCq23n3yUN6PoeVSOVQSUJhpAWcVQJt83NtJRiVTCvIf2s9MfMKWAoGzEwxVWcRnG8jV
4W30FFN2Q9l/VTFRUYZIg//1330tVxov6gJkE25VSYsAKIO8ql6uKC2n/91V1fSCVUR0te7Qz5yc
9JSFU5R/X56tffBGNhTYMIEBE57D/jdFJ4gkqcutmvq230jZzkBc+z25RelVhLTUXITPSjwTOoZi
FkFlLXrBK5rnSBuSPLuW3dMv/wI3zAT2WXo3w46tA4yiNRmoYP/4S9lMDc77aatJuNSswgIhdn4h
v4SVwFW6HQ6yiF5dUKUnHjz/qZVobbAhf9b/k3aDK1CvaeMZqx1WB1Od2+haLQge+OxQJYrAdG7N
iXRtUgYWpPfKXw++L3m9+rhvZbfAsGxkaAlX+ndMk0stjfoVV4whFRhTpR7RVyOZ+o1Ly6KkNc/T
2usA3BRQBqCpyf3T8Md6VR76RJCy/eMLiWuY2dgYPLKwOSRIItshqaf3r0kFc7JoiUJLMtwuDxqT
D2dh1ocUMZjKpx5dAe2Tr7qmXwsXGXL2WoohvUXpGhiSRWeT3SZpeDNEPvdae+RSNKNdrLtgf0yl
tuUTpyMsg6t3m8E6dIJYGbTAu184dOLvG6h3Rc6fbJVvEPTLdk5ZBEK5Jo02ChQsKXoR2OHBtRfa
p18MuNfJDAlETDink51LS60LL6R7oV5CU3l4VCliMy98hPrd4nr0kZ+Y/ExO2RPXqO3o/obkK2Iv
VT1FzOX8hBCVxjzgQRpvq8lA9jqSltpv7vZLSF8TY8QkXBv+ZNLuCvmEYwQaLGs0MNrxOP1BAlT+
A6xbGLhbZRoINtPxAKXwmFenGicml29NFKICteMKdS3p3p2bduqGyFMYCEbrND6ZsxbTpX1Z9cdc
INBqfrbNOUWWZWMfsl2p6RWy1oB0TVettw35sJ5Qev3mLrTY0YwQxRlKeLGtDM1LH05QwLuqh1n5
mq4wvj+D1b+Ie90uTxTeVyltXaT4VghpG4J2JQygbDeF1HH//ChEEA/mfgg2RURfo/OBh8Wt46DC
fE12A+PIQbEEoJZAwOnBhcMChR9DDtSat4MKb5nqudn3zXcWoscujx8Bib206YdFCjBXSb3XgQr3
mD1vAHZUZi2YqaqDHC/nfxTvloMTa0MOT6kKd5CxdY+AAtGrlLyJWOLAorqQHi0LZ/TiiSwC3PrO
13+nipp5Wkpd9iZ82MgyXve33ZqDoPtTrahzJ9lftitcYMlaZjz9DOQgymlgnepeLPkUXf7iQh3Q
qjZoAbj6CgpI0+Tw3nq6W8vOoAAG8l/ZvBNsx9usle2YVWus8Nl8HJrUqkmLvu1KDXB+CEay+xHp
gGFB+9NNEQ800VJirL3vaO+PL5uQ6fY8y1v2zrBw+uIhMNnZcB6O8VJ0XyAMtDHcDPMwNgOhErVR
kjB7E90wncbI/lN0wX9QWOc2ZCaSQDVWtqKM/EnD3C0SBfM2kxiCtHO++84HnsJnRLsmeQ4dPOxp
qAk+H4N+ZREaneTeVS25EzsSjhnDq8FHrgltPpjBYI7x3W2Z3sXCcXfhmAjcbB3K+nYsMdQ4JVtY
QnUOJBQb0x4ydbCj+DylUMLx95gf8FuW0dNawInt8L20sC2hSyhYk1cQI/zJ8s8nIpu5vI85zfnc
ncGL8MFUvxeJnKB9DGmjcZ/pO2d3gKrq9c6HVXRBgPREMFgIIihO7AEOb7kZY7RtbVOzPDWEfoMF
vlNvMh7zkpqKxeXSrYaD79VuNePvG/a6NZSs3R7Buq4W+H9i1Fi80to7VObXesWwc2eMTh44OfZ3
OheCtIP3jW/3plETC/fks0ZHKYuuBZuYry2nWWZDOqgwDKbfLGkImPWPPPY7kt4gmIuJdCECPEg4
cRbhXeuc5fDYX797BK5E6+5xQ7nqJXXl/9qrS9i6jzvdDwNqHWeokM4kE1XgRdKNaa2ivni5KuB0
e1apdU3dJPwncK1zbg484fkUzKh/iqykvEJg9h9ULnEm5G/glnaWFhOM0LXoVoG+KVey9NpfvjXp
sRPOn8sxlW1RQBga7GePDLlzcPVNwNFjGjQlDwFgjtIPvtoYkJ4qmaIEt+A3oUyUgjza6OZv6zfS
OmBpWC6s/9OflyHw3mmPYa7LVRENKTNJhMNWChf0Lv2SmZS4cqiLv6JBQ47VipHdMJXLTEeBCGYz
/Xea1XneAYNYqjV1xeoxmlaYQh8C8pltSD8ws+RlG76QeMlYXsGyZLhhf9XmYdJtIp2YGZo76Nqo
K59fA8Wu1YEA3B8iZK0OZOXRBq5QtZs/3mpm7G07CO/OoZFRCqBf6s+VuWKZT9xoCrOF4+sA0gzB
xPfUqaP81SiETXPZmvNJMO9R6Uy4JrhwGB/6qWlPlUx1v2RqBlfWbz9Zbrd5rDPSNpRqzMMVWb+Y
WSFypU6ocQoAqNhe0l0MOxLTLoN1CCm4OwlRZh3tl08fgqBRoEza+DPIjkh+IAbcIixWSW5wL5ZB
SpI+GD2yzbkoso3tQSpQnI2BIBL5q7gw5zPq/zl8IdM8++wWcYjsel/Pv5Ljwe8dp2AzWiA96Rrf
gPn5Qh/zk2ZCTgJyF5kCv+toz3mBomheBt8zcVCxdicoHmFt8yKbL/61V5v+6ImqLRIj+QbmVFD0
tCxUiUg15lACSGiVSAu4/WIiD9je/8cATnYpkXQwiIelzVwMkHIIacimEc6YqlUndxbvK3bWZrp9
6nGTUKu+4GBrA3ycGcBt/FIdKl71NvIVDt0VklYQsokc5uvSqgQQxFI92d/QVn86QhzbrSRQ7L9g
fC0bKSp5PE9oniqxuaTtbgjwtRMHEyjud4YiLmQ4iwi/lWiibDhuV4q73r0nqGxMUykfpZoGToar
zh92WrHJ0fqbeLrbswM6a6AwLnEPbRvTPenlEiJ5/wLJgdRi0xgQc14J2pVNsbN3n05mTnVWuhEf
ecddnjo72x0npXwgK+QXnMhyrdylesWRJhkjk/zca3NX3UWvDWhW5DoHH84ZMuEAOzgvFcRvdhzQ
idqC0qSgQAr13g550CgdCgHRcpb16I5GZsfrvTtu79p10BZuczYjeXcZqgDqqSxM04ppw/UvfiYb
J/JlebZfeTFw0TTT5T9oIINKNWLHDb52csUhYCo5kG6LJodRvhULmkfLEPdVsGgLNKi8Ya+UsrWo
ohmC30a9QAbKwV++8HL37PE7jtlSbo+tspzCU4AIJJHmAXR8ncaraRMpYemDwe1hDjs0jMWibiuu
WR9EoJMlxtRl4Og8VzLhDXI8LZN0DUl+2BM3gzXcJt4fWQ8s9xK13yHuBdbyHR0cLLkNkNfJwd1Q
TTvTaJOPecGPEWP+HgSHTaPHASznY2Bsej0cSsmHiIkFu0nG+ToQLQCf9ye6JITf6prRUHmQcCCd
rDJA/WQkWN3YuymFBzL27fsr+WanpQI28GEzF3ZTombz5NlPKJdHXP/E4MJqTV45HaqqREJZsHWQ
E20qbfBKryMuAfVtaPakzoI7S1Ex7MECgJ+JQLcxPinTCSeJQs85+jP/cJ5dbSzoKkQHsrbpFB0D
q6SO9PWhC7rZ/m2QJBR06QCfS2TPCNAgF2Yi00oU+FwgE0aAoQ3WOaro0Bze7HlIwvUj03ueE88m
Qyo/7avuSdG1drcnvf5FgtQcgsPy1kf0QKRK89VHzM61TEexri8HUJZPT3SmhnxoBOdtc4koLvts
T3m08EUZfhDHLq6IPJdNTAxh+3+k70XKvp+ewKU2Vd3NamNRMzTkseXAReFCFO0CyITJtj7GXAW1
l5BMRXc45hYA0fSqCX0smoqYh8f467ROvu3TxvhQvSvhCNxhttsZHCrHXZ/P1vgBMX2ibFZjZXyD
Xdg+mbIj923wQ7CNCj8n53PKGhDAbjKgZIpIWgLtpQyhwINumG/WuhM07vW3hPdd0UkVdz76qttq
ODSsYv8GQI3BPsUXwn5C6cIrsDABRPGjpgTO8pF1HN6hcFx/J/alfu/2QeXrXb2rTWJbUKyjrl6z
lnhoRvhDTWxPZJf0QLD6tzLVuqZmDM32BDg8rAsHEuBRvzlpoZzDmQKSQ5/QxBsgnka5tED8xTcQ
mNH4WOkg533Az6oDwlZO6YaELxuiZghGlU4m8VwKfou6gW4KlSP6eYe5u0xerI9A1qghgFDTwB6n
dJDndDQuOvxowmNkTHrpxp3947V8N9vcB52Com021MwM24JMgUCyOrb8lYlUAfhRTZOU8W3nq18N
nBsIzJfvrbk8cBGwyVIB+qGcME1BjSlo+NgYLFsXNnehiC8LR+wfok4Uua1RDC8PlHjBslguGNov
0XlltSKVgUM+GzhLpN31go4vowD+VMF8CXzaqghu2+B/aiTBPUvGm84q9OKRH3uqLIAjMQdxCZki
AYIKTWV/ATYLnRDivCiOf3vHGK1SHl2NICBK4BXgbc89PwoW7uuXF196A8j4/HqhuLBiKOwolzd1
6C3UIzY9k+/Wxeq7ehd2bH4ZLFgxnLpb0gxC3Zg8EzW7xUZ6j6HeXE1jpdEYl/6mKeO+6LaaTX/8
l9glA6p/ta8uDcQxmLS/9WBXUiP1burummZH4Y9S1kpGAZsHkUi+Cl9ypqwwiSSqIyXoZblxlxoV
r6er4Z9JOw7QpTtTO2eOZgRGixscjSrjQrbKeZK4wSo7FMmMTi+lyUhnbfp/clsSdREY/2Wxck+h
U/96Ea1qW8QvhR55wEs+mC2xEp1qIghlP3PW/ImLCDggHFSaJXHgEA2Nlr2QhAbZbwZAZ9ddGVrR
IYYJTI/BFzmUONHz9CTQmInS33EdbM6wZPNDZKFkCazRLVYWqx83QpR/nsv5vtLet6CnMbFCT5Yi
3o0arfJxh1UiylQxja9uCZCA1gmqc/DiKIRxyRmkWlLxDqDrK7RYUS6GECPI++5CxZCTdeHIZo34
n3IGDRmIyKkOcJAU5xPsjhAU6mDGLAdP9sFKTJ8xBq1HzORxMjBVtbdJVaOaOYQTHJenUzTDGZjY
NQHhdI3pQktl2WgtXcZSpWpHZmevQSL8srqnHSV2zKzak5b5vkfUIRruAb6ValoJAUkl9xZbzcI8
1e/SQ33rrhKz4lclbtqLshwWZPvJQ4DSIFAEwsfZzNpy8bxTSQsMRtNgoxlfpTde/r4o6YOKw2Vt
qhMHM2J8PKVERAGS8XtJFopTuE+/BzJSL5iQpb5bWA/flAdfWDpayzy5/BE04UZR/evdv8Dvz641
B8Sse8Vwv/5IHR0WL2IjYl7EBV/CXFDzvxFHUrMQGeJNGcbsnnjuIeBPWbBe5TB9/gjW8xOdOyw/
fVInwqhVbWwpweEGrGtLsR/HxxMHL6KG4PhFvq8b9zEwV3OG4UHkW4s978yCGW+6W4qv9DN0B8zO
+K42kZMgwEFD7RUjj6m3UCWt2n+dqv/mV6SDKurawrwVnaRAB4bTAd+KkxLxZ43RoWkv73WmcF5Y
wCbw1zbxpau9nw3l+YJb7yU8BdyhgrhEB7KkVrqG1UqbF9Wp9w64ngCAQYlHD0kCHXpExwnYcyGL
8SxYqHtl17gv0IArs2y2GesoUBKrcLnojMP1+kJXWDZSPKqjgs533Y4gXN8op1/3WoPJe+qh2zmh
udC5sHGi+fd90LBVHPg+GDgbxcKFYiCKBrrIdb1D/9NcqbSZFJGyZjhkS9OPP6JURoTkFYH0OWVl
JLuQiVavc71fzKUoxFs3kyLLMTzHWuMmd8q3emIPxJPOE5iovzCPTr/bQNsYnj1bBkmOYCozTVtR
/Fwmc0Q160ts/p0hCRWh6Xp7o5N5ys8BzqgJrL3KRGLlZjxFXQAFAAxExmfWmz8xrFUz4JwoOm5M
2z+sQ6i9IDgdv+lKQMMFDDn47+rDxhfmvAm57RhlR2J3pJnpE66H8anPfxj12kWxsdflsbwdTLYZ
slD9eA3cenMIBLEVOGt7fqC8vSSa4stqPkeJBA6wiJKPuPGLRLX65ybYWluXsr25ObLUlOcBzeqO
qZGZkjTgujz93xp6Ma/VK4cnu2XJpVhl+IbZD1U8I7v+tRBXkB1pFlESEWvbJDcD/207NdQ+dXrr
qB6N2hFMVVVf/lHjBtjQFTxoFyqYx7C6C7TrJMSLSdIkO2PkES0GC1sPp3R+OaBT4ABXgi56PkF4
VeXLe/0KfxKejd0TFuEjZR707ZvU99O98U22fIAq58fSbHRCQxoHp3of/HVY7PIc3RapGXj9rePI
vAkuItexrrA5YLcMY4YkBkJO0EtBAaESSUPjDzQe3dTJvG5J/MoDBs3SL0VW6CwSyAjyqkt9HXkV
bPlvjq6tlAZLaci9Kxj04SgM33RpeFAk8qpDDav/3orbsWdIzFIcR92U6lJawSJkAo/d63Z4Ey2A
MS8ncu92XZ0CXHvEaVeqH7ZBVvLTlEKBn9gZM80zYc0wmOnptXme+xkract3vEXrYKXQqqG0X7o8
f137dfIwV8G/rn8B/n5d5lNpTr2xRt2ZWa/3qjqWHQHexHvJSNvxJr85/dr3+ta6nfn0B0kcn4Ss
+cPZJ1v9C3+iTACwc/fnzMjeAoKVZoMW3yeHkmxah6zL8/ung0FyUX0mhkaYJsOoJ/cjZwSOWnnq
yGy7wj5/LueG2mY9vSPWmf9RduYznLw/FeorWMb7L2hD2KzW9wbyWrZh6YsHrpI6wV2n8BMxup2Q
u/7CV7ZRNlhYWwHN5X1ycLGDV57VXbKtMOSvFKgbe93lubjJvGACc9SBYIjF+LT6hkfelRnKVlc4
UL+eGaWVXIhH5lZBumqzd23Pn/mxlz5jrrI8hsU/eh9Ghy9tEabGfHvMbNDLRtNhHBq7bFRkq3Rv
bTIdpek9gNwJchrExh5pU+0ZxNyPedtpEJMG1p4wYZ4BJge2EuzEroKvTkL5MydGnok0VxPgEfnn
I4OUxAsLpuJAJ0udC3QXWkmw9ovGrn+SPOSWfgEsttQrlbAoPPfJBeiU406VRTPKoxVZkz2w2acu
w/RwJuwZGbuWLfvB8uk6MwAtIXS72ytxA/LxsX/ttX5HLJSZwY1Jo9AnhRUPv/cUdfKfVoT/voyN
ebOhA3Mu28uatC/+QzWwwWCmoUcsrFvzfPmIe2uOSt5fPw2V11qoVkmFOU5fSMSCox31InGnXPWd
LwCOm43v6ekxdsS0ZgrgOf3yS7dEylw14uYPHgx2HYQXH8WExKDs3h+TOe2+vNQIEp58LDAj1hFV
DT8LV8rbIeP8p5SfaSnyEwKoqnxfPU6O6yNoU+CaBqNOTo8L+6w1ArKqrwYvXCDwEbGwjQIRDa+3
r0z6tP78Ih2QEWCAilcElP7tiXJ1cQ9HieQc+TxnAI7qxjtQ6DmYNG9K1zpXEdcUrpXOr8Ug/Olx
3E9c+7mEVVyHyTn9sajshvdp5mlPTOkiakkT8N8lMVgEXnLanJGf4M/uAIyNRBUyyFV/tF0YYjYm
1e5Rh7RFPqNgK6Z8qbbvQOL8vK7SckP9GDYhjoOs76AGl4E6rRudOW5d2/1Y3EEGNqIf+KhsTCbw
68NWOZlXPtjQKiaAlqK68zA954q48o8lBer1tu+OoT+Wql5uTpq89YeQmz2ZcIdhfvCtd3c35dTv
/px0Y9rfqTS9fQHApS+IQtqkypTJ+QGbOwgrZyg4aUkTWCqXeIHjpLW+5ahBKLj4GoQw+nUz6GFu
9K9WU6TcYZikNVuo+oMvg7ouzQCN+42mM4EpAHuNyjcYX2vZ6EvPotZopgYrGo5nazoLH+YLK1eo
pIla5GSfkQybVgDnqU+xlinc8JJmdN4JrGYnNB0HqDiEKmIaxAhJpT8Ts1pB+Wj83/VEZSDXGaPG
eYCc7qOf50AZOmIbBIEM/qTfe5WT5xAHNAzoyp3PvBMeOHwzRwjOuT/eAlAwqXGWSxrCNKOYKakz
eddwTEmMdJ14OCPkxu3foLSKXW7Gm/3Lu3bmPOS3PYgyENC8o2RXz5kLSygLplC0f1CNuLjGkjBs
UMh9c2OTlRJqTrB/RgrhD2PRu1fJqzSosTsqEpiSabid/5mcsIHnBaEuLLEOizUgDi3CWxIRwRt4
GSZybJyCayLLNeUdRmRD3b+jmhCy07I5BzICuiz7upqg5g02VTwMkW0jnD1r02qGwjSMuLWmwXZS
DSshVUJljRBYWoQokmbb3S1DtRycQuEdMY9RrrCJTYvrWvML6M0aXg4C/Ofui0wamYySKAvYcnKD
AdEa5oZzRSFTsG2GJ/qkiWVTRMRxqVDzBHy1Ld1e7GTS6jVDakz2xsFCSXzsEeUGH5Ee7G9567B5
2ySwXAuME/JCUHsz5ysiZC9YFazufxcglx4/VuSS+jjv63lVNzh6rOUNCgU8BAqh90xaB5d0xgY9
hf86CZczBfLiI5L2d4PYozOXl5vSi8pwUcEpVFGd29SzmreNAXknACsc+5266Ss7aFKbYrm4RpOP
k8nsifWGjRgvxhbyx1jNkTllV7rIVaO3IYBqCR0QwkYpznYEVP9RTnZ8vdr7Zt+gW5YepuCwmQlT
+S//Un0Y3DFb5KfyQ81av34Vee+SYxEan5mUm/xqMPVb4sclGxF7lfHkOuZAl+YYH6HWOwI1lURh
z5GqgXZ+uz3pPpWu6Bqnwzy5CK8u0W7YAGGCU5KvdiZt8FZWE/J/yfubSfhX8RlZjJ+KpHmlCAZ6
VdLR9pa2c8iUFdFP3HaQ/J/ygiTNM93jpo0dfZ6jEfCePNxwgRh2H16QMoNOhgip6GmjcfqapdT4
u20ylMn+7jU+06kPhmjniVVxRIKsHCqrWYJHthDcC1zG/nyqyDm6Ino5J2BbAAvaNtw51A6cVnlx
2wiWWJTTwNXSZg6/RtR5/ckLYK+6PyfpLStlNGWy5VX12rRc4eULSyMDzkIjmZT/Z3+XJLkzeUwL
Qi3sz9QcubdeIO2bmzhA9ys7tzaswhSg/CwMa5Txnc52nkeBfIgviFZ4uXQxLNJk2gYDksC4kNZL
t4M8aj9r7nqutNHlhBxFwngZCUJs342OmuIH48DVJnYGbpIUnvFcp17CyXrDAK1slnEJ9hrYT4kj
M5dLbCIRJ/Id9ov9Ws8SNQ2+eb2f+Toq4hgMjyOWsySjBAtcwosqazVLOJzyupX82b2tda+LXKMZ
S2Ndk6zTno0I6CWNQrndBu0gfVYKxE5g328NJdep5B7hiHpf7m5AkqngK5joia5KCO1T25VfPw10
x+cVgKh+NZMhZ6H4KYztZeqqYZv+ct4IIUkijoCICFjOgPIVu1cwcGGodH8BePXQ/h/thZT0tTOg
8X0p7fYISeeGn3pUVgKtAWTuOXxQoHPFdrDohvEM7W5cGZbKjYlgicGCQuTihkgPpY/6OuM+60ea
XT80RS+MAUepZ0ucoCWb8N1kdZWke1B30cCDQ41d69Ze9NnfvpCyG6x/lRAZFCGlKo7uSB11GyP3
UXmg48PD4RLkdKtVWROGR3Lqk2mmgnKZ8cdYFEXZpaRI4dPJ6+FmZnAdH5W72knqEmZim4U+rZkL
fe4CGwur4Livw4gpXQEFxhB8PfllnXlkD9lddey+ylHbD4wMjAesmfo/+TNeHjnK7bZFLIHYjg6r
9XoGtqydbaM0kd9RY1E1TJsNfwe1bynOe4CIFYtdIr+d7GMTHpxvGIfvkNqoM4dLWQdJL/N6J0Rp
RTQVQ95nkL8a+tUn6c25lq6BB+Mb3cCsVZuudv63h/SCDP/zZGI1RbkZzFcBD/5MRw6/K8KEJUVv
hVhHtKxyRENqeC5dab6qzuRvi7xFXAtlow//vPM+edgS2PgFmIPnOXKO0SPhJD3jIzRmaDEMnNRB
aFzMdtwshS/wUoLbPT906QGIJHxODjg/4fk5WjLiPIYNR/YBQ7QpgHdCOA8KkSqZsuSXuoG0iwgX
+LWhXSmVl/Rf9VxhT8ZfUCYMD8CDgHnMiWBlOKfRt2TqAt0Pay6xXa7hjtFRN60sxt16TruQGCF4
17WBmuVI5v3F6EvbBAXufNRaxLYFwEQzuNCupwAv+8EpAsbLw/AXBHCzs5eCwEBcgNfmYE6+Tia0
bKzhZnrcguz1ukA+1uxXqanx5gHeuFCiiwSK4mPdHXF02Ax65DYkEfa0DVEQG3Kyp82IYFsa7tW0
20akFQ9YngoTp/iEClAvbcG10w+/74WcvjlHb47OerTDa1Bc4TUmcMWD7TmTmki4q89zc9uB1Rac
iqvZGd44UbWCdaNYSDwzn3cIbu0mheJkMw1p1etgT8llMTyj0YgSbAJV46G8ZkNneciapwW3AUHz
Mf7WoxEU+e9feMfBWmtiqVKv59cClTWhsMZTkfnGRm3rkDWDSCjqem3hK2GwTDzI1rkeuXW6Rfpo
CW6RZ7DWf/uLvpJMtVs+5qANNV852pH/SeBahYREkGmihzlD9mhHCZHmbwaL/DuvlJWsAMPNY5CF
un/Cfw/fWfc+gBZpZrIXq/mKB7S3h7ESI9yX2EOwdM5Wf5cdhkRl8VLhTPsnbsDd4J5M6I0zu3Ts
8Ct9uVrgvXYdu6ZPIOkNoWBpvXLlMI+iYGd23t4YTAm58/t+QZu5Vm/hiKTMBROsA0lZHJlGtgcG
bwpYqUnc4xNDxCiE1spZJHAMW4jbrWcbqxKqiQhNqaTXCQlsSNMbzVBCKYmT1ORmZd3RZVgB5taO
W0d/kqcSAGBLcKSq0p7PDtyisi5Cu/YtBObLfg8WOVLT0JYwSvVs6BrpAx/TIYHnuTJATdSNbiDn
e9IWr9r5TX++T+QF+Lmc5mynzrXV1x4W5C6KbRPWyglm7/PBcEW9zPHY8UYiJTt6GijXdDg6ZelQ
MmZk8O6XkjYTyB3Q2s6Z0Q4ts8Azl/0c0LcjMt56pe4aDwSnMba9eSncWZlloQDn4O3IViBYDeXs
5v4LxjZsTJO64L2y6phKULqWo+pWxA/nxfYOLZOcRXNMd6Jz0DPlHUZN3Z4jI3cC6f0c49yjqvNY
/dC1m4J7dH0UZejwZAHiFHtANQVw99ESwDsc2J1VHH9HG+Gz8R8XLWozftAgriogW4iQZqnI2YjV
euvZq4SCnx0a6IgqrI3QnQbJFdEJSLD3dNgscET5hDll28gLw3zXWA1jPSZyha831SRHh5qm11/h
JmFwdvQBSbqfV+32MbOSvsksh5H4XRc6Ocy3zAolzTdtifQpQ3M4d00h0A2trDw7Ic6jkvTY9Tw6
HOOKRgQxPSOc74t1iWY65jnMG5qMDzU4odG+8BfD73aTwhkNOCJUTiCbnYs7Mhpkszw6qtZQPzI8
iFohYr/7UnW2SNYRA/jETW+U8/c0l7zy0g47XAdORugr35Keo0jooavcNgQPgigRb/lkcrT5HU5a
iPLOi6xDOuqFggK1Tlx5fI2HXbsqHJPCWzqPmD+tj9jujrNAEQLPRt5S5Fv491MZEBKbYntz4lJx
MbBjO9h8qpKTbO37TV3wJrAld28B5cLfZVuVvB6xJldE1Md35a3dL8eR8Vmcx99cp7wdGRJtFqFY
XoEEdpM3HfRDx7nEFHaFJ7phf8kkiWZQi4dfljQe5cA/y05jCI86mH9N7jXIEYkys+Qj7y/qGr9t
GwxSMbY2yEx6UtZcEncR9nHeE9JQvouD365Bz2dbj2TGYqsGasUiZYRzih64nzpgO/a99gmfsknE
U91jDH/ZM/N3DusOoKcoiEiVvUBLJA60kI2bC2dYTnFL8/t2GAIq+f4kkH6IUCm+dvuCF5lIA1K5
wzV8oRCE45LhEZx/4fCKdLpXtEPjil3osq1yHh0DP7FcOkjOYCqnmGMS5lrA4G4dSCx+OmGtEZWC
cdq17rhs3VnFQb786NKIjoxuiVPztdq8J4bdYQhZ6rBYMOLASVfzHsySG5hqFhDUtkO1Mo9xgx/z
T4a19AggqYegzKh3EoRiqEU+ycV6sMQY00H1ZOabWbCnm3iUrwfNMb3nP2Z9DbG0DnXQ6pSZYZEu
LMS8cI1sIutyBZ1SCk0X/DRGdp50QsRAafiDGlQkJ6ftB/yAeHK73MR8pPW5p5pmkvvX2hdFDBI9
PXoRChhIs4C7vXpWwpIiZcBlAawUeJWhl6k6nxDjQQKyCMyW49FZRWoFfCer3e6979tIy16U7ns6
571HxvJ2ptQ6EmoP4BiEZygkjBRkTpBjc1BeDUUh3TqvOz4JP3uC5Xsbb/SSHwMHiWMSxbuT8pd9
44QygeO5/Thh2P4+PkAP/gQZNEsg+gU3YMP59aiYAr1EcOZ9+T8lL7dDPnDb1Stz6rXh+BcI5w+4
8qXFTJRwi4qQTqge356PGEudAbIQ0lnbVHMXnMFHH8ivKTWWUNgve4UwxyLrqtUX2WgPa/glhJo4
vcanHHngqBYFIftKTps7FrfQWI3GTRm2onh528hOvrZYRttp7dPkc16qgwTLFvgsQQm55e497nbB
ZSZZo21JqTADdzk4WnGwYgJPUcovo4FfUk2W9msaa2fMNCTz8Z+Sytrnah2O5+OSpw55CugPn2ZB
Pvf8ErC5H6AdGV539DgbdYYkuucBNZA+Lq+iobVHz3c97q4yaF3WhK0Ad7de2oNGYdF4d5BQOJsJ
fk2t0ReBPBKH5AiU5ATIr/pIF2l/lVpXKe86GLsZGNiDQwCYdyQkplxXX9xF1KptIsLMLegEvexI
mYOCKMINOXbPObuvQnpWstcKe3azvTqO8uz1KcisGUJ9zxI8UGh6xNM3Ez4ZihnvmJqVZ9tK9s7v
i/RYcuUWQnfoS24Nz6maU76IUeT+qxGgqYSDUV6oPa5RZuk9FhC5UThcEMYJsNSHDape6St8H3L5
l7wnQz3iRYjQeaRCrJIFuPA3fdAjWZ8ExJJiPVMyp2EIJn6wbhRvCDVlrMtAhDDZdPXCllM3l/M1
/dcj01UL49tg/U96fmEffNnV7MEkj1sMgFzWH4Gacn3NpR4LELgVNMZC2TQmwJHKFVdz31Vt0Vol
tYowlTh+OXoSXe2JKs/MCOHGvdA6+OUzDxqSAEqmedhDZtDCvgYFYtSjPRCEDWrPhbM//BaKXRdv
TZvCe9lREkpMu/sBRVdQy3pUKPf1KWNjFq1bhqu61CkBguUkqnYEmCWmJNyPCNVzx24knIarscIu
XEewR7s47Odu3ddUGlD2lIQzPpZFsgU4/BuiI2VxgDEiG4JBq9Qza1N7Aj6nhwugd3uSH0vPQQQg
gbfg/5FxwbbdHu5oX/3nzZLl2A5WxKIkFyQvaHJhWF/H1guTpT06R7ZQdprTXjfmXMBqlWuoVpiJ
euSTQ/BiDKHY3KH4u/5xU8KC3YWodHbTjs2wwY2ksQSqIuCECK0qU6K0WFbDF9MlvWi6SfwBYSLi
YoSJImvXxF6eEbr6kuXtORGVR1Zt7NMhK4+4TCaCUI7Ou/8y2QGuSZH9gChaiXa+TeJSm1gjqoYw
bTKnK5JxRN5OzproBfPdkS/+JcoO3bw1Jd4se18o2NTkFdEEjXO7+PODpmOz4vNh7whcZcwrLG57
3lcD2j0rtHveh1eSwjjGRXhRD15teaPuSEPLIP772yGhNL/dzoHoEWrmWBesgmk1CvJh/ZJtuTm+
GeERn2x/ENgzWXJnwahxnKZlajoTs3dT5m0U9YInh/h5HS2tfqtGsHs8cTVNtoMGUk5D2qznu2lp
H6kbM50fUAvPa3+DA98jX6cfBr3Lltc9J9n/AUfcA7jWUmT6wOzSR9DAopCFkS18EymlhmBwc1N2
vzFpKZtGOo2o0hif2tIMAxack1rmfqg7xlkGpxtGgKHFDUALXrvTf+Wyxn/nkVQVZLYyt1xQTHsw
8DB5zcok7sLVOWGENX7jmr1P3ryiMaMEhUMlTXMQykE+Cj6GxcoqB+nFxuqxkiM0zjzjp8lTeogt
EmielbVoig28xpw+DNcD+MID6YO/UhfJlGXYqqhkGTJAG8CGTSUqCKrtpyYsJWIdUbpzwTYAYelk
Nb8k9XzEU4825G4cqRqfsxYCyZV6vM120tSz+L7frRvaqq+V/9pCy/dJzYbvRH2h9Ws6YU5GOFMs
NcwgUFuz/TR+ySqNTs703L8DTEUoNP90afvmXo3d+oX3MqV9Nc3KHWdgJp8tj10S9Q2k8CenSgDP
hCVRk3n539cIMmaMBIezYtba7g/3K4hthqGEoBwNcZDnZLu5wfaXHLoQCA1k5M1b2c2Yc44k+pV1
7OkroQ/HQr+D7QrOBcnQCHa0aJx4uMDeraUx6T6K3mLQIhEU32xoclqplJEmS1Z/L4tg9S+3U+r2
j08tABLPs6JHYNWAEzhyNgBMSmcQWouekOAN2F6grNkNZI6xv/v9xNaNGVmLhQJM8VWcImCx08Uc
1zHo6UbzZ7eEJyyz0biYfb/ImtlyS2qvXRQSQnqlYOMUB4FkHjjbqzp1TOFz1UM97HeLTgREAeNy
szSA2AZQVi2ykOP1QoASgbIZC3ogT32Xc2IKrJcb7rhyTvNgIlMK3VMg6JpCdZY9irvqVoycugyB
oEr/eamvYzoAl7K/zOtaa/cgwyqVbIUNGsRAU1q5vJtXuXb+srY0jaq6bXoKcygVJHmRn1/zimob
fs9vjdZzS/LV0Cr9WEasaj/57FtZZMOmU2qcdxmGNzclugMDRbCzGjNif6pXQKAsj8Ck/DdSGUFT
JPHsEO2saK8Sy+n6VmQnixP5Mi1Ctt7XzSWiyxVqILrlr/ABhdYU+73KZ2bqDGzxpBGMOQPl6Jl2
CeI5Q773FdsIaNwgQL0M/th41gx4Vkt4DRC3kEdJiQWrE+i2SJ/VbpYVOnRA1qtgcqtAUx233pup
LmBTlV9E955OJ+7iU9EMwHnExWiSP97ESNNFE+LHImVq/RcmIerKJgIHd1KbkbERdnhwef2IrtS1
rEI5SFYSHJ7FjPAN5F79KsyvLSTzAf6pB46TKLWmaT6kMJuWf0RS2eiMAiyZeUgp8VamMKDsMgy8
JnDemrPVQOLomf2EyfgJUDIoKftegeT8kkJa17mEko5+P3iPS/w3D3TulaljQMr1uemKFvtTKtBH
MlAHlrE/uSH16fEBLvhhN0WZwEAsbzg/FPrOPXzwlUPrq7e5uMNNF0PQefU7lAZIzPf7wiLA3wpZ
3GlQ6gS1zzCh3rX+hev0FopbsVwXUwGjJRH1CDu/jgdPGhz/I61PasFX0w36/TbxsAXKCaV5hdAY
GYS3PSEOg8c+8zx19BLZZfjO+q8fB/+LEiF38MGHG7tx1+B18RhoGJPSPpUhhwD7BsopjPXkeqWC
5D6YOJGUbPCVhYp+L/7Qp2owkEi4qZwjoVTxybFKxg6YVp2pF9u6+fAzC9akOHmQRj9jGof3OGcw
Ks2BzasI7BxtALtD/rKEbz8IMdOkZMe2I204uyeBVU8jDZn8O87ygIkOq1FNMk3n92QiTDGOyJ2P
B2DaS0FpD8hjOTuMahQzxgiXCWVP5QK0p8f9tENl0w29j2iKlq+I0KCFYY6Rqe6e5b1q12BlXUr9
zPDxDpIn7E4b9Ey2qPUeFrOWUOuI7O+xHR38clnzQfNYKJJ2MqWhnWR0AZL9FIrSTD71+faC+qzz
5jr/6U8DmCZqmInFn7zAKzO18g4DCVe2i8gyDdMBo22gqL4rO+nv13xbr9vw/A5sFzIL31wYIE79
jWG/dKGFeWaFJTqgh/k0S/lr1R5Ypoj8Y5shk+bYpYdtcsPvSE54Vj8O0mDandl7sinsYAfX5Y+m
RgvNj9icvQ16PdmfyCHUr4HSJkgkKaWsM3Y8PMWwNppnZ98+L7U6kt0l4e9dhyqOLRRdX5GnZARW
Z73yIIdZU7kBp6+m4baP7ZQ8nAyf+hbxR/l3EkaDNNPVP4sMrF4fZ2OFG3UlXroc8fvmVvoCfiV9
gghDJzuCe6cbFKSqJ7oOxPbrY/2wmwCbbS6FNAaqLGfLFHvZC5iSDjv4lYv90R8YDAexU25e6iSD
OfsOzEMe1DgLPLwU0hCusczlsJkg5VAyqBSRPqnxN1nWDmelaKcPWmDM+kYVc6eo8Tej+meqf59y
f5Eb9W2wLoAooUIZp0xOKO6HgwCgFUuj3k5NLopHQ+dU6grZmUbYKodwBqUZSc+xhxekzF9i8kVA
mzLDvZ9Wpr/1KEPW7Q2noeO78m1o5CZ3OnFL5YxL28A8GOmRt9VdbwXETpQ2D7huoLqNS10pkqYi
KrVPZIW3ZFJqx68yxewCMAeF+Io7FKWks4KGX3WdT2uBeILDBzxs/z9cHRjO/TUxsJoMojy4uFfv
+iRGeCthJ1lVQH4Sph/5/Uhx1EbxO4u0NO8AZ5mruh8ZbjW74mSAVLK9Rv70EUoYmIJ0nO7BYQ2t
py+iYSYKsgVaFbWZBF32BBfFnqxi9C9bmsGMXDAq/7XlN/F5tP6W+OAGgI0sOOza9jjS8ppMKczx
lZYXmO4YytKEqd8ciAzotDL2TsYiX7Ig1OPgwUnnzWxeECNg1Zqm2VX0NN1ejrxoMTRmbgWrYX1x
Sfol7HS1fIBkBq19SKs//RWXjwAJgF4GovzB4BBzod9Ftl33qAMgmrOFNDwD+8SLVOo2A3XVkiPD
4FP3JCvZH7uNUGZFnJJmOCMvLeVzHfTljLgwQTMY6b2VzkPzxL13OHfCwTMhyfS6DO2gt9hJX3by
hP+m6z3OrgRUQkWvoV43HNa66R56JDHgTyDgJ9MJE4tinwTmDGbPNwuVWN7vZDqCyXjsnx+XzctE
UpTyoaB4M/L3B3I9LXve+IOQ0WLWhGOCj86zZrwS1uWLfxIkqk3Kd/7ZfrILathsDe9SHJDFuzxA
PWLIrL03Sx0rIepUpeySCVpatYJ+/ypATgltPiMUuf16RPTF/3e9pL5MJDV73Ql1SsJ0v2CUfvo7
Mv1rhNd7kZsvgoV27BWi5uML2SXx/BNFW+XvuiKm+D3OpQSvIT/H6NAG8yjEWtEqxC2HNDOl06oY
8mAihtMz1GT99prTrGkgwCY+xJyvTqdf7x3KNI3xkrksQO/gIYRS7AFah6EoFEm6Sgmr//wTNCrk
OvReYkT1V4FW0CzvE1rSz0JdN/NNFFL8FxBZufdJaYa9ZNrLWPdVpp4yDLS7x8tfwQn4kBr8gBFj
JGaWAPZiDD1IThpubqK2V5NXz8xuCke1Ds3bPZu2I0HHsBJl0Xjfls8FexCfdrJbeEvB4xpHq76d
aw+iQY6qati8+gWgmDBJey2h7m3khcsHAaodNelGI+5HaERNqLwEJeNhEjptPAGXsaV/vW4qqu3i
4siJPpv6FWKcIfYBuaynvcwzoJE6gbdorlOWOeZ8job/1SgLt1W/xpdQ70k0aZQgLW+YlOt5Y41o
ocUYvAGDMsqIVGbrdnot5cZp/I3eMBRY281DEHbKIJZsK7FdEGzR5i+QmWfgwzOccG1MyzCj8D4h
7AXWcS/qYXJCKfnSf1MxhXXTMRpnSmRMWILMFK79VySpXfTv/9mfZ7w0s0lWHsDjsHVp50w1hP2g
VkCIhscsXDhflpIbAlRnSc05gyIpgMdKrPyqFSzS5oFWo0vucQ0WNHP9tp9+gZm+5M5uUtR0uj1N
o3G8HaHZwk0JaYGq4fHl/0TUJ24Ahq42ZR88F5K/V310GzcW91s/Bb7p5WxgrAJQGrpruSkpj6Uy
tEG67EQllbCKX5ijKnVWnWjIEutO9LLCyZ6dJGGEzkFaaYtsReD2z0ujzipgjiZ5baiY+casMfte
ZbDNBGx1VYzSVLiObe+rv79BYVRnCZ5hMbT+55q5ov1Y0ADnM+z8Gg1zne2045kOMIvjY1AjA6s/
LLjyx+Oin+PcOPeIBGwXw/L0ywMuUd/Vtx8u1J+4yJWulNdXiG4QUJnJ0EU3TAdBIHad7sTtKBI1
tUCgR6ljiRj7aso8+BpDATlC3glHs+j1gAFZsBaKkeaQNaBbD9LCxe82vPBCSmaLylEr7eFXCHys
VySW6716F9j9300RBX/nScmbcr/ID7xN8y4i7k4NowWfTYdnOJLp7pCFO5DYmzq/x7O6Ep8qPY4p
q2MWG4UTM1KU5yY8vkrATexW5YmCVCphbXKCFPC3v/78ba20liZnYU4ZoNBsXNhGD0DV/JSDAILL
bsVHhy6WDplmXl2Wb412m6GjALvlPsccLn6RybILa6RzmZAwEx1EAnnGfjYsdwqQet9VBMzScRCU
pxAjS80muUqUv94Mb9WBzfdx7vzR4ncXz3DgJY4Xk7Clpnb+jmDvN8vMDrM86RilWntAgUfQ+dvJ
ZIc+y5iSUB/vNN54TIt5gUkp63PrknbiOjzhbDecc0TcKtNpHk6xLSKBXH1Ly0DAA3UYIjBCMwLN
o3q60KgiQC0KMRzUc2jropLVlP55u5gHeRdlx8gDjnAr/7LQxpiQEK2xsMVvITtD1hHWefZg6fyu
FHhqq14wiI3qVDAm/O8iwi4gWH4A+TXCrMWtjHrqGxqFygY6uShkcgMIFsuAZ1SZIb7zH+ho/rou
ciQxfXGaai1JYR+1oUA0cA4P8mfqMtZhGmWHBZtPE06HyD4xmySX2Qih8WnI4wvpmVUUEk8GQUzp
2YX+APf2Aw6t106kzsGk8MQD7SUF4g27byxIfrvEyBhAZMdiDZa8QWBn5CiRB4mq+mribQP5D3zV
76/yaEkYUs7P/9d+QSe1ElzgK9491o9HozJK+DY4/wFiRWKKGJDgGVOvHzoU2vY+1gVg6MqVVz2w
2oDgDlwbKWWWHzPpejaj/FwVA3UghwDkziS3dCZVv8uYtBuVGk+ErJ9k+bZmbt+PKVbfum4danGs
k47EAXmVkq/Qu7SW58DauH9SxP69F8XULd38hBpEeyQ3bWlB6CVBuyxaK9AQyvTRaFpmvaMTGgiB
IUbEBue1Pr4TwG9bipQV023yh3eSz2V5bqiDqcu0MH5tffGThQj7tS/HZmKEP3kSunoIkbEmVnQA
asd+AgQWLRa5f+safL2S/Y3RO4mg/kxdhg/pxk+D1E3pWIzJlUyVKSOBbKGPii7q8GgC7Y4o+vOL
W26FItgLZ2SCupyi2TvzXvALfKJMYuo9qGr3gJFv0jz4aHr9V7B7tG8DXwz9mhLjitzAyOE5fUXS
MqV371hEEPKfXjMpnlynvIJnA6uONs8RdbhvhDHqVr8gL/YrCt8Gf8f3DmYj/PEKdkCYEh196DpM
FcBT3p+pOox33Wv4DOOqYNE8Dea5Ob+lVpZvUAtSORuF280B0NelqyONoTQbp//R72qOCwH75VqB
msNAZ2GUXR3ro0xmjqSfWY5iVtlfz1+0Z6h5spEU8HUJ5TXi+d9e/X+fvOLTvTG1DTVgtRB4G1t6
45T1/qnEX+v228MyGzOv09mBVD82yohM0Mn8IVXxHluHzG8U1K3qzJQrNRZWNuItqdCXj3IrlIu/
lGaPIVKuH8zmtZUKPvO9GcfT/OVgpVy/yp9/wt8VvR0a0emZaQSgA6OmWOr3zYH1wbmH7pJTXDxj
ME9oONS1AXO9sBFFmIKBAhGW3dOVn3IPlkiiGFUXSaGwFiserFxzFv/YGTG9Yzd1X3d5D+1iQEhq
9Gz1P0JqkvN9vDZBxAEfp6uPquh/YxOsQOICuzntI311tZ2TZdWX7blZ3qZGVDLGjqTaCnW2RQgv
mEKrGWv7v2bwLP24K6WHl0ZRgFQ2+jpgd/B9YDtsyq0f4bRRChCp/yCGSRRedDVI7OcrFvqYH07V
zyPop2Y8pQf2rLPIyAlrncsdd3BQ0yG2l91JEOf8x39eDubC57jFeEeTU8ztCKf+cCBjBXqfG1Fr
Qh4eq8FGpmc+5QNYOlzgdAvQCDA3Q4d7zMcsP/TU1gNT1Pu4folC+Uy4AJYP9s76Q0UnkzrqMKbz
ZU1f2DZ1rTWc0GujwUqQnrvP+Mb0VQ1CAecmlw/6wbmPqoDRzhc1PgI6sXM1bSapoN+wpiFvEDup
WoXDEnpqTDb2Y9DyvCth9YEHLAAPHGCmE1T2R1sBXMgW96udI/JFDtMGnRRF2gBPbxx5uJUDdRGU
J3QEZOKlX7t2IPc9vPnKfyKhu2pxQPPgsq/pUmUcxclci/Tuv666no77kS9hX2GWIW9CfbJbgHEj
Lxvmq1P1/89HDA8yBARGdi5bZpmAILq56BOzt5opTAMiCgAruROaJLzd5gBuOeq17xbOnHuH1jns
J8CDYrSTF2GBmJFOnqhP3greWmBvuiN7LX2Gtm7GbYa5ZTMVzgqbVxmA5+ggd8n6iz4O3MbZ66yE
nSY1N7AWCqKIXtoEc1eLiPyKNOoCwuSeYYnjoN9AftW57EKFFPIi8KdupBtljxVUxw2htbKZ6KkK
SKOnAlZpShRfRXR6s4z8lVq4KiY9a8fxwsB61A5B5wypRnP0dGhzLitUQLicpjl2fAIHxNJFl43c
eV65vyi7FIvAxwbHfWSRDEtqXptZKT8ltFdOL04c4SXl9O7ETdkqOqGDZyTAS82Mf+sZv4PrSHFK
N9Dvn1Gs0FOl+NwoPfl79n+bgghMmO/lANEbeT9JOXqJ/r2fqM8jhsvUY6vCcMj8ox8nX0j6A9EM
bzEPn7j6zUSbOkJLm3nLs7A9H5FUHkZAQ9j/1kj2raQe3vzts9BvtQf0TNaxJV90nH5zSVlJLQPq
O618uqiOAxHft1Zr2GO0K0nX42azJ2K0dZl+6svWj+CZq6ImB8KkcF3gawz9Ts2CkPE7PsD7hbjJ
HoX/o/f0lEdnfjKhUSPQMVOHQloFpMQimVLBK13OxVhkxKhYDh55EiEXuNyZgHaXgq3LFjEDvM58
hkPdVc5R3PzP73itoGQ8WOOGo0jqxKlOAPUtAt0/vX0IinV0e3iypCDNz2hfXtCScKN+qn6kCVA/
48Bp8kXAukxU7xxTXbA202RhYHyq+6QUCIZKpcTXutsSN2VBpycCREXDBP63ZdyR0jZoDfinzJ4d
+eXZA6hUfxRHptmOVGOYYUe81GpmtjHI5vfVf2apbq/FLW9FKkzBOX43N0tcLJ5Kf03Orew4pDmM
/ryJtq/dg32/K/tOV82Yu4isCt/2T5ssz3gZAV943MeUFLsJJ1L2TdMVPd6X5uraD5RUt2j/9n24
Xnah7CwCLncb80+0zxVb55RW5iRJmGfF7HFKw5I1XHC8E0tdRtyuGUaTDemFrf66Hdn6VmOfN+DG
ZcBx8RqnLESxJ+BlPtiXyx+ch8tFqEDkIiDJDxD/UEoIrq+ulgokJftYnlrUUUUqEqYmJm51nIlP
D7m/asxN9gN7e/Ku5nE1oYD7FVeznDGkq4bHG8KfyNgQfmflQfHKBjGlacZTew6e3YMCvu2gkaLK
N7Ugvf71MofKAMUTrATXSc8zzwMMOH3uAxdzvyqMHadvHWs5vN4OFvXeadnCRDBTeHEVH63wdM7z
fML8qiWbf1YFRckazeVEWmG+8tO5xvBjQZNyNHn5v7yYJS8WICml2xjj8S1x4PkAl3CtkC+OlZXK
Icq+WcqfnV2aCRZxo4K6OOAQJWdOPwx0ZIVc58ivm8aGaXw699W/d3tHrEPVEf+AbEcHVWjf6wHv
IYvRJiZQ6zMf9PYdC/PPcn8aXWF1Tjptlnx/LMOP5Nlxk8Bwm4709VcXgkIIs4XA7sQwhskKsWuA
eDaXaDHcWTtPtIz97LL1mcyNpPFlNsrm9vhSBtJfvn0D8US5t8YdXSTAHu0Qv2v9h7rleRmo5NRN
G49XwBPDpsIK36YTAMnaMQWqfMeelaJpBNJchp0vWp/0aQupxZFXeH3k3CYk5QJq0nhCg0EGHPF/
ltJKpY5DzFZ0rpe5Tb0etJxhP4h8I4G/YuDcVMF5UKvNB9H2/JXlLVN5CSNrh8lPbUJB51xDTsaN
Xrcqa11uHzlhE7zFBzkm94C8pQ3dGvwbDKWQkSk9MWtHMY9kowi5YtcOEWpmgInLrJyh/Zw6FxVU
tr+XkQbTPwo0xKxKkofAdC4heOFnXCRt2t9LwP2YPdyAqkMKmfUXJSQmy/wUNz0zE8+ifHgPZ+Pg
iPuxz+34VFUDlOOey3siLVn6tbqdJAN/LViqQNqbFeekaYUuKWj0NPErNR+uqq8+y5LOnrgAe683
A7TnDxy9oXjiHnR69bhtn6IETOcuZtewBxpCvI0Lcy+T0i9r0z8yjq7WQuTlOopLGVWspk+UXWdu
1Dz51my4YrbLfcYEbXkFPK/vLxk1/d5FK63iyi9bbFJd1twFsohF8JMxXsspOA3GGhluPYMpXwt1
jsuHkdfLb2n5GiyfWRlppwxDSXDW1b7mjh540CZNTain8bMymGlCjaFTfJy7UODU5yQPzpRB1UQc
GYFfgwwBQDBUBpLNz27cjbCKr5McrY7dkaRauDs3iVjUuwUYlM0VChULqHY68AMiZbGluC21MJW4
G/Kh+ZcXswYKsBOmFioOytzkN/rjkTiUF7uMht+XPJnHF27UjfHVjjFf5CYybn53el70I1+05fCV
avjTTjGKEIyjZrttS4dIs3tyWVhuNrRof9PF32EFVr57OyB9zaAhSTX9how82Yk9J+mSHiF92I1a
HZ0NSw4/tdCbkJla3bV5SmfPsJxjb74g9Ob3SG08NoNRMBCidr0m8B4QV69VpY8d/U7Xyi22gHaS
TEbxw8X3YWyv57FV3erESMV0tmc3/m5BfOIIoErzLeV5AZd9H0Kas/0gI3YB1M1zesN5sNofqVkR
NPIQ2xn5AfsEdlyH5oGaj9mVE4An55BhaydwYG+uHMw+a6zaXuJcZReFaa4Bv9zz8kTnKLvZaSAF
l2C2Ymx4M8pI7SPwBUZkR9Aak9gqdW4czA/dK6BNb+m/ZH3tEkd0Buzm/CEYjhTU9YXZXGKK7gug
NoyvLTBwDkF0sJUprWtz/P8cNxDqA1UUqPlp82Hgxz5qL6j4iIUgBSj2UBX2wHOMHtK/vXa1K9e1
0Z7dpwPV6YIKymR0XflkVs04ZY6aoKm36Heu/GAIWwuX74QV5R6FhPfhhtI2vOZ2L6krOIADF2RU
Zb/wofFp9Mwmna6rQDF+qR71RdowZoTc+S7VC9gVEnLUseVxDEcOx8Sjk/3k+6dTpIkWZ5QPJ8Sp
C+aJAKjActoJY3A8wgLwZozuSVRcanvvVNFGSZVkoMAjlP0S+H3BO/uFoIuZ5pbE038Jh3px5ZQ5
hZo3qarKvYqGW75JQH52RcPuzQCDucc8nBVOBpIgJ/7Bc/fI+XohpkdA63jHnFZKHOg9/2g4smQk
RchL3hJABiGbs23HHnsRkyIsd/7eSXuS2P4eOURVPtcLPJPtxntEOb6ZL7SSy0VQ4zcYbUUITiuh
7r65MmtaK4IJGupxw3EAyilRxjPSsFGVoBXXU8Wa0DBNWi8Kp1SDMtgmiyc7CIP/tLYEf+66PtHd
QREmm7eFacvkBa13W1BB5apmDAIE1swTkMqf8wEE/vaEaP2wcmD/WyJbOoxriT2rjaeT9JW8eCYj
Uc8obCUik+hbj1Puo2wFasOdCDvHyw8YXLC7+bmFdPOmcVfx7n9bNrZIP3MFINumlKNxu8PK6K7f
ruRfA7B+15dqVj9a4HZNn2Tw+VCvUbo3CJynY3vP/g21Ny7MxphxMtPOYuvLf9BDvuql94vsJ1JC
QX8dcfH3ZISvxp7j/6pCqhFL0huxJ260O3G185QngnltBZseVechHtDFm+YxCSa9u0jCaI6l5tkf
Xmg1VePOAxYdtlMgY0r08B2KINBOxyT15pbRwNq690o2udXPFx1OSAaqeb5FdELE4BM1vGE/zqQR
bglt66Hfa5ZBOr3Aep0uhUIst9+Ia6ba0bte7Z8GUO2fNd14XSsehiJ1aExs57mLEZ0AUHTGAOJN
0Oql0RimPpAPBo+3jQU2M+MOmp6sDkOlQcaESQgbMOGefKfz7gVEK4QE5SOToBJj07SB0OUeJhV7
PGlStYtTMdqUqbuNVJwzO9nLcy795eMPYPI1922HuiyYUoVvPev3v/J8yr5/ICnfHaupZD1Gapik
d2KbxjL7K+Wk65QvzC82utmQCq83RHgXy2qIo5b49U8RcuOlyt5fpkTh4o25/1Ct0kbT+3xYBn5U
G32mICJMTHIEIz5z4hJT4ZfrX6A2UTpZT9IIB65Mrl+HsC7P2p3tE/7wAHiZASz0krwyTTvhbDmh
nPWAxZAgURgLtzlmbHTY6zeiy6mti5cgDIOjNFdQj0iGyrVhTsYq8Vy3pr1/rMOPDIb/u0ItKVp3
gEMvqeTc7z0M/Xu2oHGtnyenV+CffLe26axaRIODmpK9sp3kz5I/QrzpNF8EFKcaCP5Jf0Tq8AHU
3ujkhikIxJSFMVOQ3mwipXQT51jepQNaRm3VdHtsdXNmvjCtINni+bmjeL7cZeUnT/JHkRJProR6
evoKqQxyAq0F2/JAiZnXRBqDGYEBIz3WNEPf/RsUfNAFEFl4EwVsFupDbQSeJvIuiCI46j1aDV/L
nH9TjUjqCqGiUSslE+b6GsGXtLO6Q2m8Ckn04QNNe8302hl1i6zkTS4bhMpEVcC8o4xOBlSN7Wmk
vHMCwgwI/wohxSwBfFbTmorOr6zGmzGs+TPt+dCZ8XAYJLBZPw90kfvC4wVuLLXPWEUtlowSovGQ
cP++qupOzz6Slu+q+lWtAIxDmnD8Qez91FT6cYR+kH+HJSkhTFp4XuJ5QVkWrhiNDh1OJruq/1C+
CuPDGgu5e3SAeu2z/W+xF7Ucy/oGRuFUg8uNYm4fF8y37IDZ2jn81b2azl86sP9O2zwoVncT9Ns8
gLkw7e4pw1MEMCIC8JsTo1lI4ByL5ZoFtdDz61w2OlGjlwXNLzQ4xsYPRwE1Av5Kbm5lXGsWj1no
HpfZTGby0iCezo86NWlJxfG+8DtpXeEOKo2z2iFlfkReoJXwpQE5y106qIXFHoUfOLVbco/o+Suu
/pCPzQxYXvgAzMdPTsTAEMicUfolj6OY4hulohsNw8ouA3fQBtLF2qzRcvc1xsFUOD78saKxisV3
9sjqrOkbbd6CsTN/mdkdW5JWKbABioMn7ZJEy/qvyo9D/QLbTTGyfW4TxaSrjngm9FGnO3aQzoiv
ktPSy44QAqYWHLgCAWLppltQx16ev32FIhE8N0dcXGQyad4vRqKSo1rWfFatxvVrecE+ZAUa+ni/
V/TYjK9BamJ4l/F2/ovd0bOQC+zced55Y3Ww7HJ48FJ+lzQbL6pZNGzBF2LmHBm5OA/BfC+kQVeE
lvo7Wyl7VmRZczIRtLPEA/heA4+7xdnluulPp59s7/qAjGS/XZCvDnjJ41y8+XXwTLP029myWI4z
lAHns/48DuC1mSCkyNHVZycw9VnnyKyRM6Lw4LeET30UJW1dFp6yHvr4HP6hSms9T4D7d7rnhrB7
r5yb/dY10dVPnqhkK/Dmd6bKPlXWrpJY2g+OkytxrViMvBBzJuKeGFke5tinRXCHOLUTnidpuTg3
sWaFO4F+/JANZM450W7iCJPNVAN1eeaY0kBQbGwoJguycGxrAsWaxfFkR8WCn2Rdc7VsGbvfPnPJ
+mMQWTOCpgyWTXivFwTHh1O9ekZdP0MiWzPOtfbUNOtSjuwgBdd7gCIa+jzxPLRPSBED5WWAtZEH
VUUiaPBOLy5XCzRi3eJCkEmTdUvczMg5kH6y6DEnXbUdOGU2DsKk4429zHC2by2SUnMXHccbZv1X
c40DiLedF4Do4LoBexYvr5LqPc//HlWxvT6bSFf624skRESixc7+TR3apBuNT7fE7iHLFWiQ1sS7
OGpzuqbddUjQd6jHPyreHtdxx3YBJHYkvTF/1GvDdyt7UpyhEFgyYeIQ39g2deyLScyorjybeFgm
hexDVZzaOFjxdNa5kV6dLyWjhm9qZ9A3JwXgFcbM41+ORlfWth/Sr+zH6rTof1karihCC6fSXtak
L10bnonlVKETiLLIUNba+ilxnwDMUQhrUF2afYF4skN4ABk7JbtpUR1a0i+07pyYOCX4W9IDpGyH
TtH8HuvBpno0PZG3aTExq6I/howaSxURLV00CQZLjGWpjk/PJ5V+dS4afXXKbwi99xiVso+EcE7p
tDAMJupgrSGOMNVpUL829RSYmAmq1YYDraSxLaYq2apwj+C5caTotVrIFHRsb6XdXfLMErBMDIGL
UV9kOMqw8JHcCnALvn2F/1c6Hbt0UlhKkOYBSk4lAto6ShHfWxfuyfGXvPc9zQ44rzkmF1IrPSQL
FfilRLjp68Vn8BCTkRvnVZvWBDnJbseZL15FL08Z87hzSkoDwBG+9hPR7Z2wozAjYb3x+B/SXsS9
WGwHQ7GUPU+TfIp0dTrh6T7vOge/anzzCmqStHLfDaHVQNj0VjC7GYoVINgL+YfvhDYQsjtGRi/1
AoldP5UtqCmHQHSPvlb9OZH9RoGGE+gPhAwKMOGkCAPHO/FMxi8qjj4p4UR13x5/DkgwcsaQsPBJ
WNeDYG045qKPx/lGsf5yUA/a1R6DWicG8LPgDs91yWP/6LJMQCCCLPS8u93gvoV29XHLaB1H/mT4
+4Vy58UQaxXUEeD9JnagNHs76qAtQqe3iUGmOfJDRctgVeuwM0AKRzS4NT7SfF2jqI9QOPTPZtSD
pG66GKDl6RKF6lZvV4q2jKinu5MwRFiEfQ8WWnc2IbJqw89QKrVWzmcWHHpgMFSGYgNRrV3Hv6mg
Du/ttbFW4V7P8HtJPyIcfox/sa6JFnjeFZXElozHxgdZLOLFFJ3//0bANldqt9MaBxc4/KRDBo4Q
wpi4nkMiTNKPy/wmH+BRDG1vPHJV2eSWej0DwTjTgLExW4N5rZsgHIr/XuuUqXUI8cvcAcpJkCMp
DCrYCsNwWFtNQNPk0L3UbRRSew2KgVvVY+qqfiPsuz+CX7acEJurx/Gsz/Zo9GzeFMvKguoUfeek
ALFw/YueQkxD0m5yfkBj8zIGIDswwuGO6okIsOOGsTbm2hbrHLA7z+hD++xHg/OLtiscijq/E1ix
EUoaE3bKO5LZ+/OoAEru9UPU0cwUTqEW47AgeuSEC9HLvVsciFqtFRv1TZIueLCelciCKaFfOW7U
29pK/1vdnqWJi6+6mYlrgjcOnt+5G1M7mQJAijCYCQWA2lnUTNFgv5plJjzSf+65ekpRR9ckpaiz
I1K90Lfc6AKhjVHtIKkGOLqR8d4W29Oj1aa8/kAnJpSB5WXOUID7daCeLPA0Gc/QmnMM4LM5SrsM
J9brQJNs8mcKcJSMkWX4ZlBUoGIjCy5nszsd+425OWob5+WyPjBy4ua1OXBRAGOBuI8Chg94k6XO
4adOVT5VOYvDvR4lwvdCedgZjEIO1S0PpCYHj/aYxoOZN3C1OqBGxIC4CFAtKnBB04P8VCZSx4HB
5hZ/F7wJraPo8Lx33k8toidnUx5bHUaiuOG2c9c0Y/iX6/2d/P6U4KQ2SjeBorbEeHMIZzcVF6IB
CF+41+VRfnK4lrlHRHQlOtr/BovIjk5LPcM68MaJsaHmirUfgpKFpobx5HTMwz5bqNgRwciBsvl8
rmRhYcwI92cII/ZgVXL45a/jACnFqYqJbYUuWiBS16YnLVQVpaVacMKsGNbGbARglL3U/NTuNC4w
I/nQV8cW1ftLcWybbAboKV4FKoB8kZmdBwltFLxqA5+IIXkUpXkC2TZ2+sL74xlBPv71C217qoot
tccMWttFykLFHK9eE4Qia8NbTC1clOTfxFm1z5WLFWeUB49OBhPCkaE+ay4nIMRJn4GcQfjdmHzm
GoC25sCFWUalurU7fIOqr5vT7A7sCkU9P4BphuUt77E4UGronzLrFm+1lIRebw3N8hdkBjUmwDRC
K6kc96GzQ7L6gk6rApRmUzVv7IcCtkuWpWnL0HrUs3XVtLzlJfOqxOosmdwqKZ1MUL7cGUolLaNT
avCnPjaZeIE1M/KIqhzEstOcN6GvAmXRcN4p1AjnDD9/uw85KFVErk7Npw4S5IpImHEMoOPoDTET
a6XI9owD3ifTdXurOWvft7+Ulsg0tWh/L/P9vs8j8JhavCkqpcSsTCf9vAwZx7AEEepjaQwrsnbo
3k9mV4v5aUwXuDYuOTP+3CpLlsT9UAWdh2d9KuvgADe8aKnFuAmGzAyOCZT5/qvTyf+yew6Mf+aj
tkUUhV+1E1AOAWe9GtC4lvX3bBjj1VUkPw0uQsFiLi/O61svsT6e6nqG0kGsHhQbYL+cnIK3938J
X4HDk5yZYYygIHu2vOgIhIYg/LQZFrGTT2o6yKnX5JgKN66dmam9FSCzxrzARTKG5YL3L3EKuZaB
hRw2V2OZiuUnUV1IAXUnDOTbhJWqYmCf2clcPAAELvVzKDhkBu1+xVPLUjBERtoU+pJDH6YkYu0E
ggxuOStd2wikIjKLi6z/aApv8V7ZlB7gM7C4DPAZBLLfDpODTjq8iV9mHUBc8dOh3vl9dlAx+nps
qrGievxE8SFX3tPk5Q+mblCyTuhQgvdEAHnD+wWrugWzXVJRofzOCaZCSm6nvJxVuSnFx6MLCmbC
iJcBxzf7R/uD4Xs/MQ4wk8+/+JrnBr5HWElgawUbg4pzw5OhzwkCmfFlLEbhQ+DIWiu3WRD+0Nkl
uvnbnwd2rEOIVvd8xbxUZTm/DcwjW5lPLJbe2lyLKjKhTgCWORQWtKKkbEBRmEE3vsHGTdBaaMEs
Jnq1sraO6TA1MlaMLkOIGfZt16uO6qVk/UnpCBRiX5BbMxuBd9Wqe+B86lqhBM8jR8HXsVMAMV/c
6TuSM4OFquo5D706+td39wMjZ3aLzTN/+qEtA8+lssTd7FDxsy6uWKBmNZoIxtipgqZxmpbqUex9
5KMPZRfJGDhO2YgBkX/nZvb9J5O2RGJ9N6rj4dc4Habb4IcfaI9RESlg4iUuCV5rKG8zIyHgHNbJ
7VqgnFIsz30uQhzMkAmBnvhW8teJeOdrBN8=
`pragma protect end_protected
