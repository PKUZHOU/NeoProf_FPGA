// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
uBWvYeszgMEmDQcTbZ+Otvuy3x8UjtLMT8+uAQCEnRzUQa4qXHiiLCygrL9Epw0XJ4WzEXmwSicU
7OcviTzTptes43sUfgLuIWzfVlT2AX+hDHmRrQolNtv3/cMeGaxpoywfb438+crFhg2FVuz0sQ1h
Vb6+NxTGm2fdZG8p6O5fRMsl1rvwUjRRd3bBrvOcg8+2mOiBqU4BemqBn4HL3LCjxKJnUk8sRWJN
5svs8FZ6B9wqkvGaPY7RFgmYlD8ht93XhMvFYC4RTqlOCaV+Uod5dmcmE2ma42j/0/JKq+KwCy9l
zm2XhfIlUrj4NKkWjFd8v5yEnubMK8aOuPDfMg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 7040)
mzRguyqoy4qKKQ8t7O1GEbCRpeEPlPuUCC2qojFdH090JhP3rIuRtd1w1xwMsdQi4u9JUx2ALzOO
wHrwRfeNoGcbGR4Ro5XH5FgpPdIQ8OvyGYfhhXfujYnyZuR53euVnJYXAvyu7JoFp0thL2xrIj1t
D5XrVG820E/x3tT1B4N4reYS+lDs2IyXfISu9b+Etn6BF74fdUunhBQ0v1xX3ywgl9+Z+0xQAzW3
tYpO7tI4D06KRfRKfWPIfIrmByBfhOja/5ukjkuycwtn/alMHZOK3JE9dh+V3kcCLdc+AtIxAOtK
dBkcGrK4iXY0jhbrnqMwr3ZL8d8YmInbDBY8xton5TUAnFAFgxf0unU+ngXUF8KCF0m3VFpD8FTC
NN/XjTExGC/oHzRTCAvTQViLjhova3vz7RJ20JvCoTQF9bK4B8VfC07Sdn6HOyEjM1JivGUtYHQ1
8ZRlMMOFpw1Fu5M6SyAZZUzUrE11g4qiAQazRFOe6fBl7W0X7V2S5oNqgC8u5R31P+P4XfgVS+J7
eY/VtwLPRHFS50uyyLT/o4b8zxHCptq0Ok3kDidX3omxAeKyMaQ3gKLJSbWE3Ke50CQsnFNyWLzY
PB/iXOXz/sZYFv4lQIeK+I5WUcJfxhveSi/SvV3YBzf1FUFa5F/lpqZI20RM5iUXHvnme9IrOPe8
zztlF3QfZnuP1/8HrJfK9SPRNhiq3VFPEt7IQDspYyxa5BCzZQJGujG//bZxb1ElCbV3SiRptN8P
cDE0X72FjPom1uJLEHcnbeGG2AqclQALNwASdGI2rswNusGNa7GOgbeJIaalRCG3Be5wD2QCBuNl
nepbBdejwDe15GF59qU3GqKSErf6eMa0CbKWFzpxFOG7ycP99odPt3CL6artpo1qAmkhzcSa/Pdn
X+IvHwwSid5a5Qn8gpPtYr9OdfsNIb3Lf8ZY13/VYi32Wepv7Ww4LLJcqacD06TqYPjoY3CucIQZ
J3f0dVnxCDfITCkv5nR+GYZ6Tbrk/mAr+C6cXw/PCg6xx2R6bnlfWXQQ6l7fc7wRDu+MuCyGwJIB
iRVnPQKsrl7VYFOlHoPmJjtktxaDQHmpkWteylDH1Yi1QbmgARtcCLd3hf/LlQMI3LnMb8o42prl
QDIWlWV7IepBugathaq+lf03s8HrSlFo1s1/PDjfGRVE/i02opBgcK5ILwYp+KcHmPUWgWfSBtr3
b+nuWp+cK5+dG345d9bzjTu7USbkhg7bkAA/YnqPrEVuNjPGYruH77LX+EBH9cq3KJABAL0VhHzT
gse5Bn1hotgr+8EVSFnK4yggyrZmphg9aSz+g9+kR7C0ud6vRZrdCGnnmZZLySs6XxfwdZhiBZpj
DzX0/ZRPK7aqtvGm0tEk0h98+ngbGvtF9jptCZ7ef2EC9IaafiByQKMQK6VsNOYB6NRrR2gQURBq
IYrXA3VYK/k+rihsmkcbci3w64kGwOEYeAR1nYPx+UIZs2+uUsyoZuvteHHiK0Se9y8w6nSsi5KM
eytFYgdr5oWMcaXhJ8X8YT64ht/55R0GHtI9PIvzB5DYyLuHAld4iKRvP+qa9dcR5Dm1dwbScxzl
QMPsLkDBAu2nWvISk8zL0hhvq/S6aerIZ1UsTL9sZrm7CtddwDCvT9sCQfTXxd9aFIhCaOU+OcxY
59y9sFGZQW8au9+93t0oVcOY4xWlf+j9dAMZNc0eBq47pE6PksVtkQBS0HFZg8GRCeIX0/tVXIh8
kLrMl3kyF3Bf37dhundyg+JHTKfuMGS1gIzKsWe8m7goDNrvXvY7T/AEfQ7XkYVXAICIhmjEhC3s
XeM12eEDo3ql+SWSkhw+7qzMGZKep9ljHYlit8E2QWL6sDK8VuuUIk/KwyMGhXm5JrjZHTkVPKbo
1/AUC8izBol25dcCgl5JAtK8cat62K9R/DyxuRRk01ZpCSfh0kjQxYZOoMiWnxO1Uxd5EOtO9rOd
9IVvYDpHnh5RlfuFVBCJ0jaT0gq0NIDcKcPYHytYUcEYVEjF6VtNJjfQp4vE8QkuJm0Dsf+yAZUW
uyZDEBUHAHitjyknovpTAkwTeALt7TLCbHOakBH/c/TTpQfTJtjtMWwVlbvlDkwuyFnI/3waccFw
YGvu+WtCq4OkFZ5AtBzn44TUgj6+0xYw7UhbYs/serOPTyZAQbVea6qA25MzBBJ2xM8KQcokKy5Q
SqvIphAj843+gK4cW92WtFBbfGZSorTL54lfIDmxyU40+xjaGeYSZjzhYd7hEG+aezh8oGKOTWqg
qYx2jhMKPBBdgJebCt0ludWcrg63/OgkcnLv24p7ppEGztHTQ7aXGtOnQyO9vUPv0IZPBn9gDKr4
5nYA8UGjh7YlHzvc9UH3wimmDfNxPavQ4dx5loYmt+0i2zzNqHFZvG5uR1DkWUbCYDzqdzWGaV8M
FpNzVWAJJyylHsZEFGiuD3k4VNVVyV/w+34hqchc1S+uXM5/hQSxCn5Ugw5yRAgQSPz+vahRWDuD
k+yBTBzSori1glCSMJ/6Tsh3WYBf6apPDYB75efOqP8OmfszrboxM+pE9Wcm1m9WByeH2Fb7TylZ
Z/aFDXPEZxka3+LjWY1VpGUDLlJTKC3/aKnQQhhfqZYzV2GEUnwY3sBY3am5NhUQxgKfTGKhRqgd
QGcQxPDFauo2jYtkJ6XBFoJsxaUcAmfVbrX3xaSjiIbsJzlSJlJ71n6+xYgPAHWcXety6+3SOz+N
11Q6TF/mmcnA7eGSSQbzqovIuD5s/1685PXItrnnEXvm31Q7AVbJy44rO44brexF0lFZL2S55HmF
yG7DSK0xs1G09No2VixLcO4KUeGh8clkBA9TfY0y+ubBo06hVICEj0XZgD6CgrsNk89SOujY9rfz
6/1zmEKK4W6RrN3a9myOPoRFk+yqVeq3C14+vRthOKiaF/642TPX7T47bL42oNZ3mVe7bxlZJURy
fQIi3Wf3RpuQgANFBu8/4TbziJb0q56N49OApjRdfwJgfSGFrqaN+vDfU4oDDywaH/1wx20zCmY6
CC7VeJK1D6y27Qq95eRl8nWlgU2tM9xu2Xlsl4WkyQQP/cXXzbTW83PVjW/k73j+0WaEZL3XCx54
lEelkNXx1NoDBcyUk0J0Tx2HkaIjAyaAaks062eCikvB6ti2YJhqUIyupdub6y59Etkd7yULKD3A
pbN7bZsEW+2+/1pa8zkHtKKayxmIfn8QpVjWwdAX3k0zfip3QaRXVA21JayKEYSIuOenP5aKeieJ
Orsa6Jn41ninHIB6LuAPT+ImfiLfLmXGgA4HDVlA6ijH5oGEMiXuIS9yGzaBjWWvPP9EG1qyY9zg
VX/4QvZpZDebfk5lHK0EPto3UMajeY9oTQB4QocQtAbPPSSaQzmPAxmPYt0sVduD9Mkag12uVKuI
E/Kj4dektIP9RRa/wyN04BxtE3YGqkE7dx6YmYJy3Ud9DRgRif0HNTx8u1kGBuQh21y1WPn74k9o
8DRLKP4yUhR8v0tLIr2oWXRza8t7myD+rXA5ZoCSO9192Dxaa6Z9abbrsXXQ3wV7ATOIrQPsLOhJ
EJojvHlkdHSk1nnD2sFXqCrTER7Z5N2xhar1XqqGoa3Fz83/i2zM3aPnCfpSdMDQQsuJmQQF7RMh
SDc0icDooitTVUfPROj683h/alo9EUNVSrtTvsSqDJiIFqg2E7kniNPfH6ZpArJr7rRkI+dygrzk
Yq6aY8keoVjrsigUjtrWqyTa/h82rak2sHQops08SV2F+3BrZm/SwI96xWSlnbrV0D0C6iGtXyli
oKmxnQdHRN+GNK9FlJzwKiXYct5dAafsVhtaIA8W2z2Q9XKenQ8/WwhSh8UpCN7540k+dK51OTCt
ixuXtynyYCaqqdk4pwhWz9v8KmsVl4Z4D9vtvfkEkqQdnbmJNJ6vi30zZo5ADBYgT7HkW9Ft4+NX
NMXiEp/+MPMoXlySRrx6R/6uxAkTbnaSFgRHiD0aCEAZZRGlN21qUNRmQTHbo60J6t1PE5QMoPOl
eHp4c1W7xL+oKlE5JrhTnOfBLYvy5aehc7AYOTjR7voQoZoT+LtTxBCUazVLTP40iWH2Hjim6ize
HYuwyWJfzvqgwfkqstjhbiBWAbi69Z94v5Er7AFe1EBrCZNJPpVPKnvpZVDTv8A1B1JKQKrkJpHo
tyMTcaeAi3i38tGj4x0eRl70KN/PHZJIjVS1U9rqTNPTChPrGER0OS2jZ56FH5CM/NPSnlLT4zDu
ReO7qcuJrLHwzSRG/kOROSxdWHsAIdZNvZ2hwPi7SJdHnkQQYDk19oQlS92Wh+rWbDFxe3mX/2r+
BZppJn2SvXcxCEjLgX+PAD93BWWVaRbm6fYb1ha+IeyBpdm/0DjlOsy0R+UcZwss8UZfRQQplNXV
Pm5TGfS3dscCawsNr3L+Br97kCL6ALFQ311DS9ZO5IqwkvWaLwfmyLTVvO0hxPg/NskyurucH7Q2
ps+zrOvpLWyzQj4c4MZDhZRoNocX6GEB1F6Qk4e/obpawLuOV9Bp1fN5upKPakdDfIZLBRybjFpR
D0gSEyc9cdIzxhYR8RkOBiHg97lSL3SA1Ndp8hTAp3C0CHPLsY0NZFpjN7MrZoD/ik7WY0vk7PAk
3BE/ecyXTXEj4ol/cEUQNrTcvzcGBfvTfAPZ07LlVgaDeeyWCaNw0DZlUu1qus5y7l+//XOQRutb
A9TL0uwgzNQt11hmSpKMQPReVhdsSJj7QZTV9AjKnmuwl0KNMWXxx6IrCSqOOL+6/RVLYwKx3Oke
03WNdX8An6Q7u5WUXF1l9KnBjyqyLuts3rkDXQkMqfYzeVPiMPJl7r0qM1IW3PblBrupG+Bk2OlH
DupjWcr2bgGfUl2eI/tpsOzFV6EBVGF0jp1WdrHvQREIpBwk3D33SKSw+BA1OZasik3FDVE6nrgy
lQADytYVy4CtqM2J8eWswKEhQV5I9+NxNyz8ZnacofVd4rSTOsZuYqaEICyp+JFncxxErmvs4S2e
WzxKnoS0l65vZhZZ2jWk38Ktc8kofWVuTYJse9+c3zmNnJxS81jHJaODPnHw/WXTm2UX4Luzi2GL
KZPIX48aLPxWOSkU6asSJbdRQOXHzjjG642MQ/wuZnQ/htI7F6cVYwIumrGDZTOdWy8WTjacYnu+
O+ub8AFBRgWiAN9s9w7NYYpjOc4VaDtQkZOyylJi8LLbi17sjuQ5ew4/XaBjhi/6KMKle/XaTTCq
N8bOSAXhmDJAW/stKPw6jOnb9xJFBQqGzgSjk4xruet1X+UUUJKPc+WYy6l14XhI3BeXQpQkeDI3
gvXb7rUKjdZ59FgoS/yjGBEMw1gY0I+RlEuzvtpFVZ8AI+pY1tPWXQimb3g4G6zSid1e7dzT4JAm
1nzL2M5gjcZDCCbeimsm2Avr3FYq8YXGVZmcdxc4Qe+iJTiWRcl8akpX+O1QM/B3Rf2POKJDdHOd
/S2/nxfAKgzFvz5iMrVsEnUpRPFpQs1/L3cVjvDpplTBET3b7ctzJ31DNupDys/No8K2HTLed7+M
lUBBFvk4YLbHF1MilORMDpXcP0tHZxDctyBBr3NI2t1NnoMkBqgJsqId4vY+MYjU6+cZUpBucQlf
m9ida04rVssXCFAErWUYYBAmRjSDV1WRj0y4PhxmnyIMkshQwmHMocHfJwp/DsbZqhuLDcTzTC/K
AgVZgw9rMi2bvmy9Cl3ukYycuZii5UXQbSPqqGVyjAhNvPfP4yFFDDaFEuoVouCU6eU8izdyNQWc
VLTTfb5u3bFSTFcauwcvVRY/zlLsvwIQ/Bi7DU9TACBITB1PNLneEwaVnLhdNqLT9gHM+cZQVcfB
hgXhNXsZBRew0GwsMkwn0ZBXKu5mo5U009BGY5cq9AHFsFGT7e6gHT8PJtNIhWxAnb0F59XWJHC0
IKny8txVxQDGhwCxa3pOoypjETlNagBEOMTG/Ub3S46K8KAgpjq+K5AK4GEioU4pnJEMuQEpGXou
TVEN4rugR329v3OMqXuf2OFycUufgEli4XMoN4iaboY8v+ChO/m8+Xn0Dy6SlqFXegtn6DkWoT0Q
xia4YwG17aiFFZ7+bLXk7qqQViIT6q3tXvCJoqP81k0UA/Nxg64BEV5hUod4nx9mOaB1KW01tGBb
d7ESv8cpWe2bbUVcvlGxgrrQFOpcXuJCUjO7Gjiq49iVK/5bbLKaYsemARRiXirqXb3jyBUxtlxg
Pfx5W391J5JxyNNQMEfX91l/Qn0X8gwYDLYXj5HOWKgaDiFKlA3cz3FrjHwOJl4KWRoJiOuachbh
hVywMXfCVySjW61wyFiJRsa1jBX3ZB3uG2aH0//hOrDrkdhqCoiaJQjbFC0FW9PAF9VCOiv83+e/
iO74cdUmjZotbVVplNCpghnhTDSc9KZ8DQ1EaguWbYcE6Z6IaOEew7rwFHGarmPdTovpGx+7TIAx
wXSZQHv7Iy6kOL3ACj4HsbsXrFxMvC4v+9Ozrapqf5P/ZE7uwChj9/Gx/lB0k93W/Qkx4g+zqyHH
+nuDAgdc5sTr9urLnI9LI9h8nB04lBm3pepbU4sE60hBW5BGtAGKuODw1Dc3bMfb5GhEZYzL5CpE
aEiXF5mlBC4H6dyR4NNSco41cTaYIkhYtIhy54TVE2Nc5QN0mb10e0VRdk2/oV+N87t2xZqtS6lr
VLCPkdvXX84dN/rLUvT9CjWAzvNDPvqaR6LDOyscuu/3qZc1dyPxae4Uam4l7R3w/lsAodVY7/1B
i5njLE/QdLhg6tVXjJ+RzCytRP5J7BHWXgkdAMVMcrVRZHuotLlr+ClDbzobjN3gJdwhrj7Ba2Nv
TF63crWfQdBWuix/tnSILWfiVOJPq1CaBtAv5uAYx7qaKAClPyZNMFnOSBvdswKaqk2NFmR2Gilx
U2I4cGFrTpBuf9V9q7oXffwIqJ/PE2zpTTEiFgTlOIZsZ93JnOkVajhimOfWqhKlzAs6+kZKqg5Z
X2wPe19Dntq0IE+MAw9nKbRSSzQUJ3/pAavhuLHWZqQ5D19fpb3OL1ApbFT8ObKMlKAmKn0fYAr1
S9+lxMy4VDa44THuwD5sRVDVZ8ruRhA6graXjMOhiRFQnUKQKb3/xEw/8kYYj7eQz2Q42y2tHug/
a4gkmLX9LsbhMHesQ2bf+Pnuzw3z5OroD9lsUmHRPLA9fvCmAlcCu1zIP33WlCaWOU+e42nTBoby
VznRPCK+bo5gC2+veajJI9/+RhHm4wQr/aA5AYN3LIUWUFp1dMHHrpWOts+0cqavGujEp2KQ3xi6
UqmY1T00Au11pJXpmXU5pAHYAdanz8eom5Ou6VH8z1H+Aldqj8pEOpTxOkb+qLPAD5YHoe12Mctc
ZXY8Ye8Hrc3wsCrxdXxbqUs7SDXvCD9NMh+v03HltaDKt3pmZs4JA0GfTN5Zd08id45cHIXinj0S
6itHvGT2jZxJyONzE1J81iXQuqKE04OR3tJbMoIHaHisOZpmZDUs2iBe9ekKu5sjrLVDGyuDK3IK
AsPVOgSgFUH/9nrcfujX0EcWcJAVBbzIwPcrEIq76HiznvItpE5A4CbE5gjXYk+7G9jPbrL/0DVB
WykZZiiLiD1fL5MC9OlPmwFBC/ivCguGbJ5ykaTBHVs3DNG0RH3c5mP22NPs3uMp4RaWJIOkCNY9
B97f6dW7r2jPGnOt/2TEakivelYLTrXdfbMqvoPibkfXap3wY5rSnKHK2lXkG1RDwkI1A9wLT9cB
hqJ/wesNGl9CuZpfE1CLAgG4GoTX0Feav5lBOKTFT4GkKukvAkB0ieRKGGJXsO5gevsMAD2UZWu/
ud3msy+dlE8ARvv+BuexMrSNPh4kcxafuM96LBUxViOUnfifp1GDau4XWrkfSRUNCa1h2lhJhFMe
3z/z8E4krfACGm7y6wj2Nfw9z1cEVQuviUKOAIfY4Zr8ygz1yt6BY7L2eikG4tJzc7YaQYm/ElyH
f16eKbqngNzvcfk5jC1uhGFVXKkkEluZ6+LGEyNQ3vmYznyxoa5mHoQYPMRdlpCYgyfS4QVmsygj
z3v8pe6ihsm36Cw9yDiMXU9Ji3HmP6fU6u8LkTH3Ng+8G9GZqwTXydjn/ZR5rTjbZjYjUpvyE4nQ
v54pCHr2PBCoa3KCVyHUqe9vbEPv2KQklm6u+wu9urVmWfWvlK1aRoUgHwnGWoTlUUAUY8WbSq3k
GGULEqYo7R62ctlTpFpJaMGEgv0cXTqncubK7liH1XZB4GW6nlHOu8wIZegT9TyGoDaSXPJDwqdP
HQ5XrPkfkfrX0JbYjeFvA/eTj4ko6EF+SlF7eWY1Gz01EVADb3LHhKGzpri5VYsw3yjOh3pS19/P
4pHyMwkXVD3e17GlWiuXWujR4SeI5N91qe4+fd/bOrKMx3JMzW0FsFKksFbb0gRaHy0J6yzyU4J2
ZLZdrtPnUU1mKBI3yA6TL8ZuswwDFOzaR3oEr2lVbLMaG9DXmPahFPSKNLd/9aO7WxazhunjZQFZ
VU3kBDL039Pe+sA5U5YYoaYaedBNvbZaR08kYKR3SD0gVTRGrapW8hyhXDuuCIrw4fZ6uGGcSy98
nFt8fBpldHjUN0f0hqItrTftlbL8PE4f6RUd4OsfPV57XEIZ6hbtTYMpMn7HpoUFBw+QT/UJ6IyM
vEDFfjvCRqEAqHapBdThHlCNhLIoh7q8TdNOHBH8fLXLieXIFA8abgEKh5YocXYur5qICTyvoest
FcVaO285Q8LB01zD+Z8HeSWhMdC6RdXovm5ebcetdWF8ES0SSEVTwmZA0twCkiVoxgRcJZUTYDRt
LnF7RPrvdmDYW45XV/1fPl9Ghs0pLeEXce2hZz8GvvInLagABAVRZAxUtcSRMhTpa4GD4zqwNfGG
XbnaFHpVPhkI8XlgeRb9MkuLXeXCUGVMjGAHKGgQBsmpiVAXTanfnD9kR5RyrifRGn65Uu5uUYH8
71C8QkeHI5aSdX9THwP25epO/ptMqpy06zv1kG1vrB+dgl55zeKBFdNsTryCsDrUAO+YFZVLdTrD
i6uKHGgVKZLB8RoYDbLdA8czUzhKKphoBi1SUH8UdE075f4NsuFrPiCJwrY++sn6HrHLZjj5OwOW
3frPJqAjfJqbdG4vddVwchftJrbHD9YtE4lbe+LhOxahvEGuJpOeFG2ZtdOKohX9OgEt75qbIaKn
Y+rLYM6Fr02XmQGFo04qBAGlfdiqwjeCMgW6jRq3ncd/sozHjUPGPd9bUaxAo2srBIHdt9zpLhPa
V47BksqVilkb5bAAuvFaH4GZVmTjXEUyW1/B/TmNiD3v/FcL7RCMNIskrHc4Zf4Ygfy0AxaFJ3IP
LNyQd75wVEBsdwGPzI8+n3ElPv3T1hXn930v9PA=
`pragma protect end_protected
