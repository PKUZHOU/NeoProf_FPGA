// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
XeptZcDLn+jQ8d9BTKb8FHOykO9A8WJRG/U51mLLwup68PxAKjrAZVX05zq1
pmaTD5du3LTJZ1LMgF+VcWDYz0LvKjidvXcK9M+qJ1JoLhjkOeTGbwc2Er4f
kexPyOUzw8m735FW0tr92QLM7ezbjnjtzHOyS3Tbw17f7m0Z1NeZPj1vqavV
Q02GcX3XaWTyGFcoTJIWIy1jyzXqFFsmFXZykcqr95HKkZCtex0NaPoOkdqy
VI+cWxddEB8jRHuy/uqCd25KuWgCgMVcs28MkY8UytQns7M60Je70Ir6Svtd
vX8zrRThynwddHFP+vXDkzkGdlWxBLan31hEHYA79Q==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
axKdn84/7jXmipSjvS82LvirPqxXilzUP8iJttMP87+DxTqiA/WDlMCwcljj
nhJ0E/KUl9GRAK2UBWMY6lgi3uPbjrjeOZh8Y+CF4pm5SC3VxWLl/wL0gH+e
DZTeIBm1QiLtL0Qy/8mQBWkF1UWQGhaIkTV/O0rhg4Cmi59J/Jj+X5PrxJR0
5WUMy+Iq9Jg4lCzvJhprw8ShbOkEtmG+/hfh11emPgnNWbIVuS31ZEusOb2u
UgHjvP6HJma0QIFqQdxVcqUXzK6gBW88Wzdx+lSHgejPyxhjKrF/OdmvYwql
d7B7ex0ORSe7sBZvZ3ihstoGWCWRhOtF0R2TdW0LaA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Gaf/NlRT3zezDyy7Q/G7V1WYdTbQUiIbzGtA/8Osgnx2NpMs7XuSCRw21tvb
Vt47y9J4UVUH5BH7ULcVCOaU+oc72kng3s7b/LMfQFyPnTtFi/DTksEUou1o
aVALLJyqfgLkiKgwJRtAKX3oKpd955CGnn1IR3FiL37dU8s99PnlPep1PTnO
ZOnZkugalfHIv9TBVQ6uT6IwhYIxlEjFACBrpjMIFNTZGoShpVUgUw9+vOfX
6AerRgEvmwy9JIVJ/Mp/DyLYRr68C0fumnofFvA4vEUYChByvgMwJaF3ykiw
MSPWeDvfA3wvYazqe+9P5HgZcxdkm8RZRTmoVyJFLg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
IsUuRWzcsHJHZ16AcFXwfenmAdggIUqtaVCMO1Ne1oYr+IbPf3nZbf8wgGgr
QjnlfDYyoHdoyfhs0vDVEfoLzAxi12ri4i38js4Vk6bkrePz3woIdLsrwSSL
P5Qf0IHL2hIWO79VlYHIQQjVZkUYyKJALO7TbPvWSQ/mSU/sTuI=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
OeOSqQEQzS7A6RLhh6zms9XBLd9ROtoWYb3Ub7KZHTIoyKZtG2IsmH9lh2Cy
rMq8HPCqkn5A/fcNLZwxyqHHoPvr8spsIJTxGXLjSrfecXpHdvz6M8UuU2/L
/4DM2B6dRetQ1dH8hgvBMYbEoUMWRrc/ZZPq/ug5SA2BLMf6r2pS2GiZGOba
jHJC5kCM7gtiu7DS6oBP4JwZ/nExtXCEKbeg6UsHb97if8NPZTaDXKIFmAu2
nhtEXhc/EX+V92Bv+GLITViL4FnQOKNZtbakbg2lCwXc+dCqT1GofGcdFtTv
fBrdb8LV4q8Uk04h3x+3dieyMwvSKgBS9NtKzV4l+Ucmscbt8mOeNQLLH3vw
7l0kDmbLXRrLjoAbNfGQZAjmDJIZYUBP6FJ7F6GQIS6dof+xSxIMeNWaSqXV
cMun91MutTTxksPrHXG9hzDHYTQpuZUbH4OyZ6N6eecTusNLPs8XhDXfp+xk
6r5Jx4mioPli7FFr+xircQaZ3MpszDlo


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
JuRkmGlaWzjmeP5/YOP9JSePq+eYpEqgOCOX0TSM9D7/E+XQ6ZVkXq19qKbP
TBRpsriVS2qWx4/azX7QFL+k6dsmynNXUZ0t6iZXgjYWtmaKMSOGqAT2268i
JgEFMXE4bzuoMAXdg/8Bujv0ARIrAiSBZxt+Yhr3w29445Kd82o=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
YxFKtwyvNRRnXTxUxQ1iTU6Bn1/zPBgaFlEMM7qNycwA8BeRQTwhS0YcNEqm
WMyhp76Q0vADx8yv4y0cl550n8X6X/zTJ5MDB1aF94dUMOBKdGko3KB4HZat
anbwPuOfeUm+Dmy/3pYz/VtWKcjivNAFHVHTaJYDzCDvJiDQXms=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 14752)
`pragma protect data_block
q2dvRdqmiGjuwSbHGbKDxcmgznxxkZEV5laHlW5fuDgp4d81q1oRspoftNnj
RjtkqVKKYcF8WF9IcEuuSHegePwVSKyFJF9Hw1wgUQhoPYeUrv0l1wte6cQN
YAKjEuFsYtjWq/dUNniRhoba9Cpl+WF4O5XNF361CzKYiJ/uLeocW0p4E5/J
shoNu/hsO0xbS6UVdX133elARnmzIfvkxwUVT6ntgw4D+k6S+YQxfiaqEyag
tesDA81IOHlCBBIWRFQVWa+aqApTh8yxryL1ajh2TQu8qVOAab+sx7mJ5XlN
gD938zADNsyRmEu1MNEWnBQK8HzdQn/vCuDhpXAnT4j9t0ziGylBuuXNni/N
NKPixbrh/9IFwgbyAhH72H5zPAhZ29FxN2hzIsCM2JTQ6/cnf9n1fXeBD67b
f7jjJI24Myf5+9yZgUDQR8IIjJfsukPU2k+p7I9BXIpirsr0wmVOxOxeToxQ
sYsKzxN1ySyFEVoT2PTJcASI2PfxwqGz9xL7hi2DUQGCYQTKrA28eGk6r9eC
AaqTYMofsgb0YcRc3d4//wWdifz7PUN0pmHcVxW9YM3xFQBy7WhhF/pxUMvK
dRz4IIqGKVBQpKWYgOtET3m15FwUsM2IdiGT4y0Ml9Kp/DLYOZVLbQR60T1i
Wh7bZJ4lvhlXr3ygD3FBQDo0c0AE8mAInJ9MeO9PyEFcTlC9gZf/mqYbpxw+
BBJaXq4Vn8U2Q5yVZKrZpNbjBE1jmBgbsUjzlb3NSPeUlCmcXEpZHPUe5Z0P
RdpPaqNtRko8YmFyelN4IExQ+acw4ECO+IQ8F3cFGuJMgmRyp8yHU1TpKSpu
qplDC5uexa1lf+zkJkAQrTaWrCjXG3PeEZHT4qSl+34zA3FCofuJ0wCcy49f
AF27xoNjeYqQElCmxkX1KAsZHNYoBboIVwmt00IX5a6juyyXkn7g3+geF5tW
GkDBjBCXUDTfCg6TsDeywcwpHsl6A/bQVc4hkRONRfcuSzNLvDf4KDEclvfD
us2MiKWRmqhor41VPhi4s8AfRmKQwrXfYFbGBOK4Eg/PvbqxSJXwwqzix2iw
2BXHAvCOZkIDQcMKKCpGVMNlQKjZAvgzvhNH2JpFoRBBo8aU9al1PUnPX2rt
18fpl3MZbhnZ+krQ6Y1lqBtueEpSntKvMrkE8NesZzM8esWEhaRMVjh7FbG/
p58LG8CA269mKEF7GObq1Ik0/honHsvyKjT5rjNqXwtYhG34iFZJQyvdqnGR
uHpKs4e2IYvOaUmeJ8o4IQTKELqi968+XHEJ7I5Lllr2WPKQKFn2tKlNZ6wR
IAl7V/yNh+U6/J2J9HfEn9zdOS0cYfwm7i0dTJ2HWaEGeMJbhduOKxJ35rl9
QYw7DC0tw/HvgNYtUdXrR5jIDyzHjRRZu7/rwgtn+KVNT1Ng7jcDvgEny72Z
RhRQSC04CPgq35+dLSqs86v9kyPCsxHxEnwll4Hu/lBRkdxfnoKcK0VwoQ+a
BxmowdIpf3HdvKfvZ7CvEaQylXQ44Bpph3lk9u3twPSLUQxuv26Po2e2iJaY
P1+k3WEXwQ16BB/Fmoh+wwDmVwNB1gmGMqxDqMKlZj532hQQGyuIe+HSUrtL
Iax/+xZLDLk8UhJX28nHanN1Jp2QF/oz+IUrgb7bhiMfN4++1VwO27pWjG7I
NIwE4ZgzJ8mvc16hBzgXU6nedL45B/n3PZRjcbgfovB2QrAG5Z7vRMtYkhNU
CepXiELjjBWoeg6/abTQUjdIQUqsuI5wcY1EnoqbiYpkmgFAj/Wu3NKoKWYI
2M4JcNgyoLfvokj01cLmI4D7ysnKn1Tbt4eIkIgjw3wMOZlZhKAwV50mcp7z
AHdv3PUzmhkDLFYN14/UxU8dTfMOynCers2zTPlwOK5NgK8wbBZL13/zxiJD
2Q18EV5gcROkEFceUJghHClDxI4JWrc1TxdiEiGFXAOzHnNgj99XpuxfpS3W
gQPPK2cKa3hxCYAoWUdAzM4NKe2IzI2rO+e/H5AsoAAXxWvYfVyZ9y+sNuHB
kbokR50R0+iwqWqcGNhz9dS52tRqNb5Mbq4hjzy8EejQRJJBTGNvL/BJXfRl
jb8/11qc5V8wKFjBjuP+KMPWcfGZ1fBzVpQpLYQRlb+GR7yIvHJAp9jU18G2
4+OB3xmI4eKq0ZS08xXIAv+Dmzog8PdXRfLrwe6xDrKlgIkbIii75rc2IYeo
xqzOyW+MCKQwC7szul7yNP2c8U1Qqc6zh3tvFm/KHnSdOdAz4vlEm7nKf+BV
WqZbyA2oZJ6MbvWST7epUmNdLnA297VmuSzWlXvix6AyXq3t2M5/p0adMxh0
HVAq7B+Oveg8/JjXEfKjkpDIFoTb/rrPmzzhgunUTbgCyZ0AYg0WntvFM2uw
h7RiXlbuSDRDon6+z+AdWF5QXrjS4G6WnLC3PG/gFjMz41me2j5inzp9ylF/
usAKR38p29AhIDYD1xleba1rpS6/67ZreItBY9iuRvRSzRfLkmbJxWdSO99M
4bvqHev7g829Smc7V2ODhVIsQvxmUMKwEFJj6XsILEeHVea2H7v67kW7a53F
XH2AWdKv04MKbxxJ+qXEIQvWslNU3TpdmThE/ldv7hFY8i4w/Qwch9my7kPg
lZWSxP9k6n/zZhTMd+mMTKuXqQ6d4fuWAJFwimYgRzjovgmOQFc+r8ApuU1K
ARrTY2hryBwLjDQ2aARf3ceWQAhYiRzO5tHokjmUMTCsk4bM/IEzvj6+6sv9
aN3NQ2SDYdSUDZJruTJg2XOFUMoY5lWlWrajFWTRqIwlCV3GeHaXcPDBfpMV
4bZt8m7+01dteu8iFP4mgr8bk7ZuSFkDSrkrFyyTu51WjmKNssaQ/AAaUM4k
UCxksk16DkFN/7SQ3qAODZD93b7j1QsOCRqEKg7XAdlqm3WbISBt3GbRNIu5
1d9v0uDnY4rYqy6sJn5u6omvTYTujPXfjW9WesT7/S1Nke+4YVT7SPrbZI6/
C7s5Ha6qdfIAGf859NHSK5/Bh3X8ObTY8RYbGv/WiYYTcF2G9VTTNupkmg4M
g1yiF5js1qE/txKNRIiiuMGrhWSsj7iL2GHjIhv/qYeuP4GLZFf0Fqb5MT/U
v0FAYWCf4MZZGTmiZ4WwfPqnkcP8AbU2Bl6VcO0Lhdi+KP3xvL17H7TkxNkG
kEGo+cpfLlXfugYny6VNUrwFMGfs76gIX9UKu/+wS/CM5DZAGkJ06pfzoZv7
oiMA1GJ47QK6vBEBqfMzcUMaIGAv2/h1H1ibbtXuAyFBfaM2uWvJ6zVfjvAA
6arpN4tM/picJRKGrCczhCG7DluvvIl1kEgxBUrB8UxJ9NehS4vDdTGvp6rw
QQr/RPO0uh8amfDxgzVPaCsRaejzVag4mNH0tlrJ3nwI7IuSAhJ4LqEZz6Qv
PjH6FZQVH4hxT9i32SK7zQ0DSh2V47q5u1uSJDjJUdTngvcdDFlazlzmU1Il
2+GKGLqFd5kvRNO1gv/w7dLILCqpr2qhnbAOBD+i8VR4ebsHD8HW4Jr3ReKb
5iV/Idn/ahVZTXtRATRinB+RPV4nHcSALGncfs4SoxSduB51llW3XtUNvB3D
Qmm4C45LXdFz1v1trwPbM7JotAa9lMp8OjI+GdJOyGNHWabypbfdSEfoFkaB
f5CAiBq140bcY4qUYSFwM0w+eLU0AH3I9Gf/j4r3B45qgjj+e/OD9uJEwlSf
CWVohe9DBOsgShhUP81wkx1gqlRjjpxJSAlw4QbhHxMDhLe0f80yTp75ZTim
JEri9SwfG5rA/Sjy1tFVJr+H27NrV36io8QG1SMrEH0jgJaRvRw/IwHcnrCW
D8gvulq5B5uLMxn/ANIshDMdd5fcUuJn/Lt1Oh2VwYIDDjNCcIgMJDUbPxXZ
GB9hgseRb5pFNvnWPfZ7XPecNhC98I4tGzE4fjcwWHZPbxRAS4NKupnAxj9J
63BEX3GdFv6hntuQbTWimZKpXsqdZn5j7KF2E5DgnWlRUIaX9wWtwHVd/DpF
TLdorTj9yTiXo37eeXKciokaOlqFofIFm9QhkMZAFftAxXV1j37cRDCISHEH
vPGEHwgzNCIGVJI7bdTr5PaLziF0cNdqq6spN+NiS4aZK80zjY/zwJfNO2Y8
IYYjJZnC/jobS6KhHQVu8AEbqvMjUsdl4y0vYmN9CxBhJozJXJXGOwtNIEDb
EKKyoASAc3bpkdYNRKWmtVJKgCWehAUWhGyjIwIQRPdG7hHbbMDeuCradkKP
S0VV+VT5fxnMuyNEeXLznV0AslgFJl/VEQRXCkh/PfmfkJm8B6ee2OkFubW1
sw6nU1vrEvLIne1BGh0VBTY8BCC4exzGZnm2j3ilrKjbugxWuE0VOR+f2rc8
C3xcJ9PP8ZwdgeQMGW41RBhgUsbdejg7AchvR9hVVhjXcydxMQkhhXLFCxe8
rVfcnEJNV2O0TC7F8vatA9bpKWOmyPnrSv8aGoD25GsXKAmsXZFGjxRMzzjv
YU88bWHUJDl1GZV6Yo4ljvzRKvIVarfPJYjolxOcqwR1wVELjLcghkM0hE4d
kZEMw+7XCG+RQwb3NRe2rJnRDSMlrOQORkb9NtuH46lReFTUAvOAj/LkIttg
nmwjrmJUr+/bFAcLF2iICHl/0ZXz0n5Jk6Cwws9ULDoTdT7Cqc0tFjJnUnFk
l+YR0LO+cTpAuU7/y0j4b3m+v01BKmufFaeQeFzEW+eFriICXPe1UzfS8DVu
9VXllVlKE4HG5BqN91GbwnUKRnwc7GiZ9SibDacdYvhUyhjcuLJIdwzVGH5g
f2FietcKJsy4mI1CAkOGc8/ss4XW5cFQKdx8lvjjIpfVX56NWeSs0nGwSzh4
WPwC+uPRsp4zusM3eDAjlbhEKXoyPBIbTItwWbOD6aLZNZoCeAdFvvTPysHR
Ylvcjft5ESlNOQXgM5hXb9b03buXpHOY8KGa66iRecc7aPVbxSyesHeLo7yL
o2PPm+p5WLz70JLgr/BOTtLTz8FphgBoaMzjGImNDuDkA4ACvo/YAVu1eYRm
GrYs/GdEIW/fcAiOVAKqsg6RUqlTENi0x220vcW8Gscp7yOcrmfohwhmBKKJ
DU6aT1VtJwdG5q+ZuKTlegDBRrqGgS7vk174Nfd3gbonwjDXodQfQtvNWgCv
ltMlnh1HaTA7d9HTIYc30HXITGwdFj/uzyJHMxzFoJGqhyW+lBN2CaRLFqyl
ix4WjZ2rLxTQ5+0jSTK2+hAVcBP52phllFQ1X0YnwyyprKxKIMZXPo52pE0/
GiBc0C1cpdXl9jY7DXbU/c4kyxg6r8UK6ZUFtWmUKcIPuVd6MYi4FRkFtrY+
XqMhRoPILxEqkQnbhH7H8+ZHRKUOZj88QUoLomru1dtM5zhjHin73wmi8MS1
Gipn74l9WimfTbmmcjisoHVOLahu54p1/UkfYkVh0CVZJySyWSXiqBVul4qQ
0z7LyGO3KeiHW8tkNDVCxH5OJOWHIcrNAMv/iUez+nhTttPn1w+CRSoX+qVm
rsVsH+6OYRJ8LVsU/Ei8/GlTDbYIUMvRCro5IjpHvGDvmcetFSIBW+IkBbg0
699gVju5ShFfYV0sJ28JR1MYMpNZ+doKmChNVevXldQUuBeXo9oJwNsY8N6U
T8AkQYLJkgigN+e8IgpJgWXj9wFh17su1MPaSaIHTDpuRVeJd9mPMB5wuRtz
Gz+0EJk7IYxs1q3u/enYIjQ3HOvws6fF2IkEXDfRzmk9BtfLVOhmDh3o3sgz
Kb8OMN21mdrvjo426vExM1TrTsDx9Ozmx9GL4TLJRrPV8l9J54jFoTz7Wqhy
eLnV/r3hi4Xr1bCVqVRlEQuJrxDyrEQal74nRMxqXHAct2UVMxzHspDb2ZZL
yniW8v2TaRoNK15ZyzwURswKph5QYLtQSopVGTNwDBHZZaxfse4Ey3C/ZBqN
3Kb5PHFxx3nJETo49g+UrAgtBBkRu+cDCNSKTz15c7bBF/ctNSATkSdD+qcl
JBGFVHoPCNFQGv+6tbPkHt5KyMwtReqiDF9u4PLcx0paeIOc8rkaAU4E942f
brNDQeMRl0cH5GkSmTMFRCM0VHDFYjXAS4aXTxIkLWe9NIBQ5giQxLT+qToQ
Ksk+40/B1wFPxdK1w89qwM3YJYa7hsRlhNl6Nbk5sFuqdwb57VY12moG4miP
KjwwqBz2sdema7NYNJaEkEwe2CiAEl3QU+/h7rqUJtt0WjkdwI4qUz3YY6Mw
syKuOxEa09QySeBinM7Q8rJVz+6XO1jFyBijPCBr/la4WsIv5P3yVCL+vaUV
ckDZmRoLXCNhsDb2IEJFk4BRr8dUCn5TlGmlmPObywhGqlWTkI0gJuBAfr7Q
c/6dGU2RnVWyhbpS55PhKAwHmJ+pJB3WlNHYmj40+NXD47bKDUUjD+UgVkrt
uTA1kS3PGJlSXrXZLRWPt00TvY2m73/IG6X7h9kjyLQFbQIb+SLY+5Px924V
bSz9fbJVvGHsZzhtPoj5Xm9hBPiOdkqFNRiNxydeXavLPpb+qbwts5LGKFa0
QcysVFMATxhmvPXOWIxK2UP7JBBk/6YB4w0hVKznVWLNFhJH5Z9sldmW1naN
zKcmPiTMuJ1Lv4K18mhS/Jtgv6zsZt/y7CLw5OOZeUS3y2nWGqXbDxRfqISx
0jS6VZdaDgV58LE4oM1A2HxMiPGWLMrgSHkU3PrL+0IQJSOx1hk2WX0nwQwY
HO20+LGVJeVkr3a8KGPi3aOPuHaKNXvuTWhReLADGICpTs3/YdtTzttqQSle
37MSMkMiE3h5b7nRV+K+iyM5PUtdaxvXf4POoByCTN8tHQWn+IqrLLq3W9Ke
m9XRSRDivysTrcbxbBfj0MPqLzek1r7TaRjVbVFvOV1NrYNa/pyw657kHnwh
NCXVj4owAdjdWAQMcVBMkapvL6K2r4lp2K2PVBNEdykAdGWyEfabAkM5s1pE
IU7Y1cFAA3BroBmSGcftPx3xVo0rTnVLfphgO4OEfU/dybuoTDoLB4rYYVPN
FxwhBxT5aYaYKs/U711vOerOOvOpI3Lv+dsBkOMv3PM5FIQHF0b8l8q6sR9U
VuSFSz//mbuf7ZAuHLcHD9c34cpp6C/nyJ0ae1t7MdH19V5cy40ivoHE3Elx
9fShcuQk9q5ICAZguwj4BDSAf8U9l/Wnlszr7wINv5Q5XKKdvnajPH73vptZ
870M27aFzxiHBU4/Jz6hXgE6cfQk/3fWD2c3S+3ENgEd1CRhS39oKYQWNNdP
XZZZFS8QFVkoBr526d7GFf7nNbKnDV8EmSZ8esvZ5oLi3weT/n1d7eqMdu0X
LyMc6kCaxz9RC7QBh89Z7aBsT7Sdb9Hf1JkNsfUGZFKCS58O1d5YpcerrD3l
iecwB2CoEQJnppLGIBeunAnAFGfJfLEKszb29ZU28ObLZ0bMMQXILBscX3dH
OgRQahAYKbZNTvZXGRFyxaqVbMjzEO2Zo3t3a1Sdsp4xIHEZIw0jzw+ux9GO
faPb/LCrKVn5AbD/cJKkorddP4MD9l13Q88Qo8MsRBXNGd0zgkKIMoE9pW/K
daqMvkvLuP4iypMcXIoPC/6l8CeiBc8lyvm2pd8gGk7ydHMTdAPIQtdOxsl0
sHUZgijhnMJaRC33xxUT+qfh3uZ9TyVbQAF0UsnnrkkhWV5KlBVbk0MZ+AMh
uucZO4g4xdaz9ohzKnIqFKE+lC//yqVKaQfsxED7W1C/8nKrWFlDHUgg2Mtp
5pxg/Fx4UcJ33FrCAF3N8Hdvs9MQrhVL9/KLjYhwSJC/AbHTM0okPcIQ/+tD
Fp5bSFsu2COSMrDOphYJj4N/02iHVH98JffUJQh2wdZJCgNqRj/7IUqLdlRC
A4geGI6A89p3ugqDO0ixoa6EcKsLAfWbKfjefIR40QYNiFnlMJzEAhgbdRzK
xDVPMCtkS5/w7GQHjfhkImtU+xhOajLz69Nhi/rQhVCniC+sS4AsLYECUGNH
DU1zYg9qAEfmwPlV+u6JuigKn8+bDGCYW0+UPcParTHam6qFozBItEf/1Oxz
fW1/ieAGzsFPfnVm/ODOJAPHlI9NKPJYABbF9XuMUGzucYOiBOZkMQfmpyiB
X+l9RfGl8F/1qO06TDSN1GdxV9OJbZhsBBOeRGu9J58h/G1mKohK9u8B+RPR
KTZ59PcDNCFtNF1tJW1bhwdygvJCyTRv6YzeacY5DVsmJiVErHYYRhNFPfGJ
N0+azyvwTTvvjuDhHw/VCc2kw6HjyQUepbZIAL4bFWPPOx4tqzEk5YcwnHDq
SSBbY73hKvRRRiRy/rDdXkYe7u+jI3votRSL2bx1hDMU4pALiCeQFT1IbuQR
eVyehcq46eHTZCH5S2O3h9bJk/Ir5rXhe4ulDet5CF9mX/zH3/oas4K/85um
bCBlBHZsuT1+4AP2V0zblETUU3GcagwUeYSrgQwQDf2eH4Xa3CpSGon2XKw5
KtA1lwkgRgB5X9b05xaUJe4n5MTSuEVAxBpBw9zbVDUbyuIrYLE9D/ckJALr
bX4HTAMR4NnCYa+Wlrzc/DLm/sYdkYnV5bZ/5GQDeSXmammoJTHdywX8rxd4
rahLyE8a8mEvWhXpnjAPXNP5Yki1c1rRuFMuRVHup7Us3JjCZXKNfQZvb4+3
1KmKO4KH9kVWmC7mLTFk4Ms4uCa0yXYJpUMzcHftTMSWsxC0ysJC1x5djJxK
MlOA56MBa3sGUvVOkVh5yV4P0hGVlHGpZm/AvwhI+RhNoAi7UTZQPSZ8CkTu
Dl/8pFZpkQUxTI/EEbOcrjCU7S0njK92PnB0nVCB7a1svtyKIcyiRQLCGxoM
qbgrO3Rg8Ta3uuvOaWk1dyiHbmR89VmYyAvazoVwXZwes8BuWCsCf87emTkZ
O7mYW7C36sIMy1u5G09F0FkhcmfsN2iDD5UHs9O272HS2pY7uljDrrJu+wP7
z/QPlxysn/lyDzYKDOePJTlfOEjGMH9VetjeOnr+H48dfXnA9tb4K6uXEEbP
9OZL9RzyOexdm6lPJdZauhH2JEJBuDJtVY0Hd2siVD6aroJd6BOHgru7aNYW
L+cAtnMU/ytBhQPOCZrjbdUOLICI64ELzChnbqyZuOS/qOcJnnzErl8SGDFf
ASYwcSkoADnFRb33CrAcP5fMjkguQ3rkZmWS6uDL5oeeF/F7P4mq1kSEc7ls
xduGQpVfNjNpy9K7PyPtpSWH9p4RB491nB+mMxQ/usChTscDoH89BceNMNT9
rDvN1Vt47evy914YR67HgZAYrvyO9KpHEEuP9okVurnxwIUt6OEhKFcgVibr
ltmelFeD+H2tHEpXYuqE0ewwk4TyQM92V9Bflv0ksauXQu9+FugP0XMEFva7
i4TpCrmeAxf3UUR1l9+IIm7pJqYm2KZpjaE0YUJRkeXjzLa/yJ91kCN/MN68
N0DE2kbB2saHJQpuHyvgpxOc+QHaHKIymsNZN0Jf+J6wll5x7ZGSpfs02B9p
cdZRPHK6bd2sOWFeU7pHQJaPHBrVewlOiuSR4VRpD27H+ImbkfeSPFYtKp53
5InVT8V7DHj2DnY9vrDrBTp3YJcre0CzNO+fWS0icT14HEHagDYJGDVv15bM
JPp63z7jXd/KgtCxitt4FwWtSiuSHYtPUQ7G94mQkREb1Hm1zu/dCQqRHXgo
JnGYSYU3cqAQ7nA1co2+4a6gTBPua/eYHcjDinmP6BUIxm4a6Q0/Lgcy6NEk
P1R9fuem9t3M3DEa1P+7249xxOfxAssFPCI1ZJ5C18fk/Vkjo8I2MmWfA2qM
KbOmoLRjMT6TwiMj72mEUbQH4FxQEwDrL3mlMArv2XjHz7IU46YWv4vfQKo2
9Y/181yOT7hSfgu71uGKLbBN+1OLFOAamHncvYQB9KrlUGiCSzPuZwFMu0AT
65hSoZMOmMA2F+cGZy7Pop8dqPhYjROg1qbyozhyXvX20ty0l6zIc3uM/vjc
ujIhE5M8fBPC3SyYbixLWG18HwJiA2BKYUhQX7K3VkMUbwSX2JidiCCwUPf1
LxbFPMmtTFGr0gWuJfnO4M0K5htzN45NuueU/izmd7KKHmPHn4ADK64GBv5K
AX65HgrDc5Qgs/Zj9XKFlePFjb+aTizFBjwn9A7+j92PXUjufbZEMHWaRXVz
Jcz5X7Fa8RCzxu6PO/RQZc/2Rh78sJFLVOpjj9mlcrMbDNU+P+C13rRCw40I
JQXwVEGxXj5oRjLEDMiNT5FelNYzEFsjG2tHkv2UPS/8ov1fkWQuUsMGzdJW
fam11WtxpRwV6JejjIs+D9zrCJE07HsLsVLbj4wxYJkHG7dGMtAcCNsoecER
tZ8QkJFKJRMe344UcpkvZ9rpZ2BT9sfeFs486jxbaEzjYPqoQGMgnpdJEY8L
PqDKhT6cNETDPcGNhpPR5FRa8JhFCaDHanweaK63Na6N3GMtEhaEJPbHjRKJ
9a75gsocZ1JJtEScBWN3ioGg+oZxvzoHWlVGtyyNUlHh4lqwS7YamFDYqM+6
jXgG72GdqUCjlRXt1t5JXQCZb74CKGzZdkGFqGqjzuA6XMqlIRCSyB8maiMS
lO1pajmU0B1jCwpCyzsu6ke5sksd0ZqSG34tbkGQN3uqqLhDwM6/+uIIZXuf
FaABvyr/mQHjhyxRxXhz/dlq5vTfuZaawwA7c6lDjc3DeSmizrMxZ5BfUh06
Zl542oIfTZxeV/myuz6yZVSCZu27R7hEEttxM3iSbDBsMiR8uIvbIb1hFSEh
GccV8UMDsJKQnCCCE1KdIyRQPfYsOj/V+7AtUCGGkQT4s3sYs4GgF6JtBOOv
cR4fH8z/XJTu7DXJDfzb92aJLlwzONcWWER0Wclp025ztjwkxh/xDm5MT0qC
xxgxLBK3GirI8GNLQXCcY6ywAW+qf+gIDjE7TBrN+daVPT8TTA/0DpJW7F++
C3sPM+5BqxCrTjYypx5U0IU0NObnqwJfPHAPd4gG5TuhJnyMaSsvS8OYxvTW
OSO/JvAfdq5J6SQkvHAMN66qzhvsIq1r4bcg4wasIJc0gHrpHrrqGp3kk8TP
Q+9QgjE/Cv8zfndl6SGOG7FGS/CPOGNjpm1uH4+syOxeLaRr2D4SCcujhncc
oAofEbBQmcuomLDYVV9aHhelUinSz+XxYxZS1biMX6LWJ1/DHvkJIbhbsuqb
GuVY94zyHUWtVuw5PikpFjkPIk1zhm+py/Cmz4PRgPaH2kThGh4oEBDLjEGF
HQ6Jcm5wvY+pnFwW8a+DbSh9MpTnY5voYWpVPeZpAP1Ipa3Vor8Apw4nkkuq
lKqyS5gTHeWeJMjWWAD/tvN6nH9vTcHTdY4JPKoo9TdqXWFcDNKcVtvOvIq7
OUPCkZ89CdfENWOzhKoq7ileSXiimEq2SFgdH8pQbVl3/QMLqZjyY2+GGswv
FGx7IMyWlgjggU3rjs5Aq6CCg3ZnCm39NJeA3xLKcXxeDQ9Ci5fhZjEPTxoa
w7hdvLXGgl4cqGRjxr7JsePo2jQQ+lagxh/HelUp8n0R46Eg8VoGqzoCpS8Z
998HPuh5U5SccLGt6nSPP6yNn38gMDX5RcLcDr6/snerR5Y99tCGDOd6W3SO
1qz34AetB67nb1qeMWv2aBaezhjz+tlx7/xebe8cWHQBC+BEM6FhdyNOQF8j
WFq8YX1clQBVyetf/ZMRD/E1MlF2Y7eKctwRxWgr94if2/bdqwP58D0uzWb/
XwVhd6+BGIwdUYL+LbaQS3JDnOUrTIl8XRmMuz5wllSY4ay/Hg5armavZZWL
UgQ7yjQOUVFytBiCyH2l2XKpiqJMD8MwAuPfVYUfEVIJ/x/Nr9Iy+3h4Ih60
3aq2uCH2pncJKF1SxSyk0Yt7JnWsDi2mnWz8BbsdTEfHGhXSzqXHLFaiTMnK
ckQyB4ZM4epBUodHuQ7VwQIjuEpWqyr5I0QA6kbfNGnBuY6KJ2DglMvdpWqt
oIWPrpJZ77FyZISZqBHNvvFoMrpZqYQvZx4ZSRLFwDJVEmI0QUc6t4tR0QM+
x/sTwJfD8gbtKbhRN3vaLp9rHRIH81C39pS9nb/e49x0xvasDCBoTDWLG7Ls
nNJ4cySKyma0p3DC4jErF/+yC3OshaP2UTeiBQ2xY+oiYN+YFfJwOLoua2AZ
kym+Umu3DU7J0qeGxlo83SujzUa+3W8QH3ndl2WjZ/x2rC04zVqdfLfbVeP+
YSei7rvjEp1IP5OSuCzeGUvftPADirRBV4r92SbwAE7xwQAPmAPulAbZHhzu
pufUtMzOqzCILUV4xVJT8FMVTfDc+PXw87k4m+LjLFYfT10w5KwGiepi0X5c
aqZEzIVVYh9C8X1Uq4sZuna69PL/W5enJ4B49uOkqtVMWj9WsuSuagUs/AuG
+4B0Dw1Hz36GKYU1xtI9kI1bZpefXycLJvaJLmExCAxwUZwht266aOBFNDbu
9zUPhTwzR41hKsJeLzXSHAAZaYJGqEdlaTBxaJK27fsc/XQz2vMubyjOLlqy
X3xWmda9KkjPoHMDUg5Z4K3jTQuEvsSWq3ULHdQuLwXVqq/1rNCld1jvnoWY
4G+AUlcpUY0XHCKkTC7c1XpkCs54txz0qoILOXwjMLLUtDSUGlbRINzZHKjw
mCuyCnFRbtIIJd54XE4rWP/aXikuPBObwbGEX93JEpOX0ugauBUDETuh5+SY
OCSQLDnLnFfJ0O8gxUrlXqRVE1dqClutLPuvxDVzax4jC7UxfOCDp7Cqyp7I
ss7f8qkakV7v/pG9DhOAx01cSdU7rQ0ra/dDZo7tbyt24quNCoGmW5ZCWqLn
gPlWsvQL86ymZZKpUL1ZUy9Ec8JdAZoBNfwkK7VaNOyEI/UZgoSUG/VMsI2L
RpPNyy1Fy3PUo7Jb4cFUBVAk7yfsieQfcLv2OyI+wwN9pLgiiR+YajN+oEJK
wzpPNf9xhDBztICDtQ5mcrll6ewYx5Cnt6dPaT1+sci6i8kNGDYP0YEBvXwN
jVxNAJSwtY6ff744inmYtMyZLdtK0sur6/GvG6j8k3Fk+cjRb/Xc+6fqqjU+
bHOOOI/ag9yr8mLzYxBzWBHwCo9UmHtjur/D+G9cHl1LCHXZjQQNm/+1284x
Sn7akym90u9e627mVljuRPR7901hNLFMnlCoQ3p903muRr/dKQq2zWPqv1TC
A9CEiTPcWk4eMYil0ACVQcPbsRTvU7b9/+Cq8VlTdKlOETo23si7c6IFxYDO
O5fkDVMVdNSRa6/c1ATWIsfTXgnhJ8k0kFr341Lo0sPyQetBY7KwAeGrMqYN
RLJTSwOKrb4x2Kvt256RbGHIZ/YbIax7SDRt0D26YulHYTP0BHXyHw9E7//p
OpECAmErb8oXfTfL42VRj2AKMvXuWj3rI/1tvypmDQt3Ckcy/cIXDZgoZIBY
7iVed9JF81wEDWYFEeT7GmqeX+blJYsw5gftbH0wMz8MvrFu11ICNcarHf8Q
skK7qECUDPfoUtajsK1zO0kGp0yeWoid6l0QgULGaJbFm5EmNPJ4mH64qTCv
Q1qgWPQGRFYFOd+Ldgmt7wTZMQD1kKnjeo8udaNoCrezfSRk3sDkwiHgcLSc
7tlscYE9L6eamJZG7twEZ+H655SRJFcjJTdUxu2vfe9v3AeeB68yeQ+8hzcf
IM41JfZbNBLlZQJjdmRKY9P628iUkzQ+aVyr6W4TLnx4eww0eSLN8zlWSuUb
pMSpdFrjlZwUJOAO8DAtDIM4y3d/wrJetkF4593q6pDLv25PPAIRxXabDsMN
Tnm9sJHSB18CGqLQGKRek8EXcR2Tb1MjkSR98yu5QRlGA/HFWN/W1SfY9CHN
crcGTpn/UbwYqCI1Q3VHoDzDhrfEp4TJjhLe8OSArDViGgc8PAaldIIlXhLM
Pm7VUrdBQ/8pyE1bHV3Mcax3voPuO/j9xGf5DjlFoMTy6B33W9uDc58kVaQH
QP01EV+L9jF7q+Z2oLWtQlSAf+35BwX4UNuvC/pNrZPTyVJpUvc9phtUKU1A
9hXXGVd39AQ+tUQMi5FecuSsF56T+PnyavEuown5nGTSZogZFA+7Q14upXJg
8Sdkzjl3BiVhiZTzAaoxRwfzioujkhy3e63ZCRXa976m5cjikEJwbeQTcgrv
WRCgUkrmz/oic2BR0F9lByERyX2zsBU0CJQQYhf1Kos6oPJpqRzoBgr6e4JL
xGlemubMWqDmB1WwbCDNRHamm1laeTffab387JDC5YlRtMMPR9wbU4ywt+J2
t1NPHKILrOgOtJy8kA1xaTzx1ZhAyP3FKv6RojFm9szXizx/oVqStCc1AnP9
2RSaimo6W94a3BUsoXclY+bPqxkkT/09yu5EMCklKJYkePdTCuWb2O+cmlRw
ykzVti7Kut5byTL3xLLdHnRnExBvw90S1nY5vsyaLgTZpQJ9PrERQbH8bhGc
M3UYWEqnRzz5FRcRwaULFovGtXGWbNMX9/FwyvmRVIJJmYQQr6xB2Q6hJ0x9
gvGlIP6ovqGJfdQwOHor2ZYt0Muu4FbAV342TuGKxw7FQhJ9xB3w+7Z3+FLc
igfmpT2M1U3awmRN6npJ8+NCIceAeeOKCU+b21yvMjpl8ksevSHDyoQT7rZX
jRCj78b5PyDAi4DtkwwuXaidBMZRGBFJ4lcaCgfqvwKrx7fFWk0si8kiHNk0
qHr7hjKClXxYXLojqe3UcEaMhCaCFT2jiGJBamooKRaRsU2KM5RXDK9Iv2qm
hG2PX45HjsEK1lMooZ7+8N7noYDvtmg75JMxmtwXHKHjZz16erFktdvNplph
k1pPC2v98RHPGB5Zd/uHPHK5ml4SmaCGosKeARJ71kbbX2jyGnFDXiA7dhap
X/BTq3AQE0Og1XDq320UhlSXI6DA6r7vboUGTd4bNziOJDtvSZBcTD/szkV+
wEDJVDrREFc4aXL7zhC28pWKEC+FVIqVSJtawZYizO47v4ye2JIUVmMLujmd
OXzHXhrtrEFxNWfA/u329Pe6W5QfaVivBl8WM4R5YLzDO6EsZTz4e8o/zyQ0
zyHNBP9AdTu7qOIdY6AhC+vliuqRx5HH2iKnq1lEqHdwqWy14pnjNUl0LC5g
et3OQiBGRCeu7umu8wwAQ2NbF8nxRA2ZQesAR7G5W0VA31D6zj0urfJLbKtx
upS9C45xmN+ml+jp6TvlcQkdjYEwcktNgvDLx41dvjwtkABkGUAHH9KV/IwI
ojAKFTshC8+NTZKk94VLuHNA3s8JXeJIKbFlXZ2bNcT8UzhdRvof/X/J+w4g
x8aSfCPfU+MegJEUO0FzkTFXtsMTqTfVD9/TkBPkfjsq+bgjxKxSdn5gnTxg
3P1TopeHzSNCMLvSYQBc7PwnKRRhyY7OYabpmbP4tiOyFO3lC21s+sa7oNJX
F6d5jHpQIyAaVaQTjd9fsSYOhxk+bqqgg0/i5g1mpEz0Kl5gyRtWBKL5LKp3
7WeLA1YPUrjlzz+tmQwkuKaR/39+L6oR96jI7qyrOyGeEXPwDpg84yIa9y7a
zTQVZmLwLhhs4U5lgIDtI9nkRw2x2XR7jRmohXDIXytvXQcAcKrOf7VcdcQn
sd+IZcBfy40fKtcGruaW1DCT0ZbarA1YjoocA4rr56xDcPUL7miUH6rmhfGX
/0NZLp9q/yPYbVobRJn/o9kD+f5LlrHY+aHkzJIcp6CXCsItcLk/Lup8GkHP
ApCkbxvWNdqWGgFJGBYzBx0fXew5CkXchjA3L8yBw/a3/fpZi/FmHRxq/YrE
NobZGsZiBm8j+p5HgOT9aaNJ00pq89TZa9wj7775ecwF0KZPkwYH/bj3zWz9
qSya3FqBH4ttxgac051RzWA6ibkDPmgLVVJ6EWLx0mukLUX8pYXFXAl6S+be
O+j5V0zclRYUC3eeSdkQtzzUdzFsNjhdfjZ6UFXbijqr3QGh7Nbdbcpl5OVl
5Da9aXTEBPEbpu7pc2iAB4fhg7UBdH7L2rYsMUesDzSfVPEoUAlh9bLAdoGc
XE3UAhzwWaBbN5mtMPc38NHk4Du95q6QDerrktSHnqbd+3Jacaw1vx+XcrXb
Ne4pBBCisHj4ImPnhCYREIhSfhy1iTj3k3gywvujYjIL31wwlGHpzEWT4X3t
+iKvFAy24HgBFBvahBje9auDzKKlgirZpNixbImQ85SMnq4xuQg2s3WNRfnj
wWhMCmZGNTCVYkXMiFR8kAam7vSKAhDSltYUP+zQeWToRlVecsQ2IU5d5F53
aN/lpMJ8pkCGyfkAP5ua3l1dd5eZd0RGAW86lbJtWOuTHP9aabWDKJ7MUFd7
+W1VL9fiVBHE3SSrT98FLxqrUBMGGtKC0iCPR5zSJy+qQfXLKspFtp07CoSd
F9CSjv9lJYFsHovu4MRZj0czYRHbxZQWeG+RmJcQLtx1p+cBvyiT/2AEoddj
u0ZCcCOEWynqrla3i1INacx+7hskCBsuNBSjbXLu7FTcSHUacIgOx4Pb9gaV
Ex/PTWjiKfCObSNDsmplCorpRP0xZV2zetMOXk+JCGTGs4W+mCxbnmEVqsZc
WcpHS9U+C+XzWtJ8WP5C4ntPHHqtbOdENz+iyj/y0L30kwrYNH1kPjBg12oh
je9+JfpP6T4LryjstgdT/XxwXeW6rDamEOrSjDTyhfUMQdaR+uo3e2uejjOA
5RBbmVkULSnilo5MkZsj+cj6KEnn2/5XgITbptq2qBMZjNxjOyyFm1g6r+Mz
gJkMYOH+BQeXQnIjXfs4YaOoZwDRkUeSu2vWQYr8JyXpnljPVJWJw4I/e6fZ
ccF9bz17flMQE+Cyf+Ra926OUh4QYHkHc9bY39Tj09SJdXyp9dc5gDXZ2VOK
vD3bTLZ23uiqTvUnCFKUEagd4y6wjjmMOv/BjJqsMB6JJvF4EoQ0JT2XfDke
zo8ILolJRvpmRYm/TEWq2ScAfdabw/OJHHZtpeZXRPiAcTb+SgdkruHqqKA1
nq3hWYP4njw6B1M4mm9ixLlqzGHdhdy0tlxsTy50yb7KmwjW9Y5kq8FWn3vL
rJDpjshF5ys8RJRdakNMr/gqajXeTxevg21VxtsZgpwd4CPTjqyEaIk+DJ9J
zVs25CPN+ll/NRvrN6D41iEWc9YnQoLpFXl/TfULkvNq0OCPwv76k7A7on+I
rMivHumevXQ54AKsIodeajYlX3TazZr/Su7na71g2YPNguz/uP6KtWXabnVq
HBgRxs/kceztrrCaZti0q9URguUs+sZGgNUvGaPuxIzmm/Ggs2BfvKdfkijC
1+Je48rc0Tb8UAXCiKlTqfFeaG55wUBGQ3kftTxj8mAgh0dQVDzhqFGAdo1R
hrcXwmkAytG2VhZLnGQUFnktvpxH1hOvBPOCe5GVwXqq+sGMX6dw9a2X8AYg
mppvbuSg6x30X+bFToo6foDo8PpQM+pzBT9z/CNsHcuxSvLZsKDk+mPFHPJg
+HIB9FTAf8x/taaivg2SWlnVf6KPIzc+9LaZ70nUk2GSEsHXpzpFPXrjhbIE
ov0Mreymp2c+uAxjL40NUAgDdTzA1XevRupbWbL+dHc4ITwkwz5MoLmm9bMZ
Ud1XcYXSM0kahDvWqOAj8Xmm66iuDXG+Avg7Ez8GkoSoOIRv6Aw+tuV9Ind4
+6VBa4Qd4D5Ss+e9+EiUCkkIFZOFqc2ppaEVmc3zhk0MVvRlR/WmobA4jdKH
Hpds72ocv9UopcElOEpPBX/6d2ZSEXD36RJGVWbwYM+4fin0sTTWwKvEpn+u
5UMO+71fPYfULa/o/QejXdbPQQQs+dkQAz0aN2BSSoni7LXahRucNhlf0hZA
cNbm4eJ09/oczz/xYnHSGgW2mgz62wFY4jTXzNuZJ5jJihwk2gq8HF8hFtmq
8IiIS/0Azye4NurwgLqMczCoXGD2155AQdexj4n0HlT5SWuh2P9hMbPbr0Tj
vAhIAZEVNnHDgmlrMPHODaRmANiMxUjl87ONnHtc3cE7xTM7tbOWmlOzvs0g
4mKXrKpu0PZCMthYMg1dRWIrsX2hSaojZ+xycEl2L1dy7AI0omcm9k1GSsCf
/XnjgJsHTB7POUGqGSf5ojW6ha1PQow54oJIuAUIVmtTdv0Gu5uRaj9KF5jP
W+uMyJELIG2IqZSh+/bYbeHsOTAG1VHE1shkeN8NU0s0qxGg10+ihgyRkx67
BD3GoApWqLvFnXktgcP6P+eMP5QIMFMQpjRA8Y42Bifl15vW8l8BSfwTT/FE
IAao7bNSQy5AKR+WKzXjO/wItB7GtLo8zyUvVk60op5Wp1+3YmW77ZuK9Hag
sYk1cu0lJ+JGZ2iDJtA2Ihkgspas8Cfk7Q4OvHKqyk/gR8z5NCNxswp30OMw
z2paL35ssf4doH5nrPavhBBaP+vbV77ONdkj8qOi+2wmO020U5LZSJCSY9Ce
H+CLrjbbD5fdKEprDxxC8Po1F5IpGJgHjAEA2myahUxU01qL21lPB6U0GAZN
v/3vAiESkym8WfUWaRGO0nHs2fD3knK3bkY8Xs1rrfsa/nlDKcmAhoSWdin5
Slqbaqw2OersUXSwEnFc0QG/PhX+s1SCEAi62SkXnyUh9fSO50HLIstD8vFX
xbhBllUWY3pkacM8AaD+ZBkz60NKiqwWnS9xYQWJyVLipK4V1SypHwd18S5Q
rD/MpPAFFLniu/9ffRDGcdiZzySo89U35LQ+h4F6LHeYNZslT77S4yrAEDx7
8QlT71DmC83CSrmMo80CSSgN+inQBvg7kw1tsryisuDnqHhBffahMIx+WXEI
OUCgT44M/AHUklal9OZYnCNI/62UyrlDQkY7Sob+i/WmNOIxyc68S+etmkTF
8T+f6SNtAV2u1yNbe5LiNWBGSmuHA5uGocaXZYq3J1L3GoeOKjwQrzPQ3t2T
J4H55y+SXFSQqkMjSCwQPBJNrMb6VIg0avhMfYjviNMCFeYqE8Q0tYd0rygd
ASGQn0P0bd9PWkD8xsyamt0O4r9kzEFndE8nUoo/di2+XhRCT5kwTzjB17Vz
8k6fC7PAyNPNx2JLcr3OEyDVtg/IZU/LivKSs4a6IpLLnrD/a79DIZ+73Y+t
4NUdpUZpuIS708mn2aXPXFJ1Po1FujaVhJA05U3B05dLPSWz6mSTInKhLdY+
nt0j4cZSJb8hwpQsSHlWV6nbie36SdVksNTZ6WSeHA4LVrwmJvkvPu9S4d8u
X+MpEGzLN4v6wbqw7oAXsuf+meQM30l2QLs20UJ2zWXvqYvlX/AmZL1dJrfK
sP3hstXhPSYJT51jTc1SFh691VHveAXBILIn6x9A+01h1xrz/1+bliEecUDi
Lto7VVTBLXNR7qmde54ySdfmBaKCoCXIa8VJ5lJtGdrK0ZIftjXZtwnx0TyR
2euknVZbZs6ytOHdgUWdNw8BjG3QgB6uYK65wX148nB7LbqT7941da/gGUo2
8F8t56M+momT9bTLUZjELx3g0R3KIYgckhRS/liyJjuArEzYv+lVwmOwdw2r
f5jMhU2b3+Z+8VVxvCQEpgWb3ypGmXmC7H512oo59mxMsZVq/wsHH6Ix+6UJ
LB7S1dQ8KBSK6hKnAw0HC8UIRhzTv+IA2IB0iwIf0v/tCvab4yjZ5lvgfYvq
5di+6C7gaQ2AYMJgAQQoKkzQy+hMXt4lvL29ap/S4RjvU5aXNnbXdtKxwcPs
kjd70CMaVyk/BeTYv8A+4sX1rqsUeSf3w0+cEJ3rWRmvVt373A==

`pragma protect end_protected
