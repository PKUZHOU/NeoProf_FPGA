// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
z4mxGE4UfTzr/y/BTzg92FjY3UtaXW078YKOyIlnTqdodtpEXNevEvzxKl9glvdT
ngjDwWEAqP/EuiGoRTCaSMWt97fOmXgQz/nO9RQxmUT+9NZSuMgUM9boozbXrPap
UHxc5HdtGj1A+d/vJsrOQ4Alz+28fzjk+Rytje1i0d4=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 8464 )
`pragma protect data_block
bxYwS7xEMiDOHb4dXWmPZv2jDhVzIB9UHpZTYXtw4vmk9HRUxZ/sqweX98WZAdIo
L1tQGlzG2dzDpMfgT5RxPgiUkmcshZvyWtsiD0LKwuSWlPFYnnD6usSWFrvxvaMw
EgSM0ZfNbn0mLwaYgVVkUTltZERp9Zqj47dPyFAOBRP2AkXFlGie1FDEgeswSL04
PIv4t3n3J2a2KG7qhRRoel35ZrUdrrfMPPXQjsbMHt5sBnO3JjKIBV4w/NZ/bzUp
fNWHiDCJ/0xYHzii52GR/YPrNxW6nbc6Hp1Cn+m5xcT2fMLeo+C/kXV+UUAwAW4e
2m12R/9bdHe2SAnY+j8da3Yuq8exdtO7H4fIDRPBHjpeFdINkS7supAxe1xjW1Ga
laTRfZqeVMRNyU7bwY9DM0plwUjDxI9DYcr/kIjQmlW0V6Cn3IpQYzyD58htClWb
+J6OnHUQdkZGH8BWEls/OjVfy2DSfTUrCGH9ZNmQo33HZa0Im7SQ8KG+ft00Meov
KJZt3rOqZW1e+O/bRSIJ56HOQ6st9J6vt84OmE0RcCsf+xO5evneSBKgyN4ATTF5
EQt5xkAG1WXMZNxWnXsbA+AN3i5nTXsMjhDvu2nuicvCXdyhebxgZAQRANRUGwv6
s8X0VH8z8n47HX6deQ6g1Sz7FAn3OBlvmbRjT7wbAiXJcS7LOX12QHs2oLTs73io
mpDgCkuanDjPLDjfuTptF6wgxlafglniy8VXm4kNX/qT34REc2GS4EpWZT8tGrTd
qRBqpliqntvebw4QAwz8e8QLpUgVot2hSHkeiV0hbrAo3zD8RjlUksEOBPWn6nq1
8X0CKLiy2EnIrWtzVIKlL0ywLFZk7cwIHXGkXoqxhUHhlDJeQBa3eid2d+6Ywesi
wFF7BDHYj6T9YTpDqlwvy5xPTMNRrF+cI+cCXEo7262F/B66fmeWygD0t1tkR0Hk
J93G4rDcUOSeuI2ELlOFE3IO1014URKn37gvCohEbCW3lzOgRVj1PpI8dhH72spR
5Gg74SIhEAbWW8p+YPIRzTjeKvPkCYeItlZYxDoWfYQaIgdQ+6+F/vbelMnzrA9Y
1TLnJKLj1JxhEH6PihW9aLPoqbQkw2WH+K7t85Kq3/XbXWvB7s8s2mvzHtGkvRv4
UGAVwkabR4Os8V7Q8K+XrJnDVO2HIN22UVYB5DstP2JEIVxgnR3ki3ydFdVRrUDt
GbMKXPAV9TrZSIAv6dCbt9rTF6MDB6AyGbfm0mvNhYelxobKsaHiMcr6f38/ZJYr
pYfhU7GdkezIyrg9MFUQZ1zgv1q5zkWvjOMp+l/lromFw2YGBpS48yhcebMRVNXa
i9fALIjd4wJWlGF/YeAuEcYi18CGsxR/J3a/G0n3j6k2WMlGe3vh0MPL6MQqR4+H
AS5ihSNEnBZPLZyfNa1wp9GdWOUqiTCPvANdgT29hdpWVcKpeB29Bi6NY7/3KWtX
eerw7jFZhmPZDl2hKg73yLgAlum+m8aoJrg/xTUiO/WljXmYvwoQBhAIVqqHSRA9
4uh5mWR+j8L5kgOUPmcK7eJTnR+E7AbJF9AkaLB3ScHWJNSwiBxk6OP+jwds0nFj
rgPMpOFV7cMFRig+lzxzR8vLXmCVpeROm4AAJQbPD3mhEOLaPE1wqvroYaCfhnBc
yC1hlCnV5DVQL/vZhL0pMQij+Z4J+zGRTu9t9Mfnm1m0CIGxHGIWIebnb/8Hh2Oo
K7fJWBqTTW6ss0B3OZKum6xI9Nl6WrJGCAvk5jfculyaC4v68RY1XMUu3Z8u/7a8
mY6ZMX105S2x3OHmFYqVN2GzygiLQhkmGhKYZT/BKwUGPUo7/H9QQwKtJJUc/FSv
Ry/v6+GFVPxMxwU+zv4c9x7JT8js//Gji651jcKZIvDhk2ccpj0xzAdTJT/+lZXW
O24MnYE7qAaE3ZLpJ3uR3ukTsagk69EX+KfCfNDNB7tlXc872ogFuTZeFc8fY/R6
7ZaOBk9zkjshKJskVKjvIaDv65/oeQipBRRBS8w/Yw3ec3JcOcro/ifvq8tQRE7n
qXb/H9PuGLg1AkSruF7WJbWa/3h4TX3HlGLpSbHnN1t1ixJv26B3PwYHXPkypB+R
uzDK8UyD20n39iY+bsCTinZapytmE7Dyj1jQyPxrfDzL3xQHZvjxLSwxXxbT3t4J
96u/8PpIlSJEbrXTomaKZAe2IqJjfkiq2XMKdHC6AHyAqUtQnur+nb+zvLf6b8bh
Lg0FmnN1F0dZACgx2BSLhOJbKAQwozYTtAEgwoTQkbvL1qFgDKJRxBYihb9nbr7V
k+jT7qJKaSr+OdyTUXRIrOg829QlHUgfmDv5B3oGle7hfJDN7qcIDpTJnaiWZjv+
eJ0GPpuxdGP56vZF3HTqZEgR143+50Dpjx5uEA6rd/eZAX8QuJnRRV+UPiGSd64l
C8D+5b9edxCA15M0CFgl+UThZTtik7ph+qA+NT7Lfsr4ixek4cmcOlR6Ppmyhxvf
dNjLP9W2DIw/nUNHziWs46Oc95AEKiuf5Wy1Leor/MCr18pYv2mmI0f6UTli9hHs
Fm+50BfpikmidzFCZ/xIyNkV+QEWLW0QluzpkRZkCEcI6dh2exbNaXE0faJVk5Hr
vpnOuLyhqexiJksKGQHs6+ixK7suic2I9a00ImF1IPeZQvQv0PNX4Ru7QWXB6ylJ
1Mzh8+vzxTykCOyGZ45ZjcXHAooC7JU5BOn7lZ2WsIcaFTS5coy473I8vebPE8OB
GIdQGO9mxGCfpk8u7CbBWzbq2LttbgyBKrLyRXEOc9a0TCKZEWdi3uR8M+ohCDDi
Cg/c3j+182/UTpzhSgBPPyE1hbxi3vhNTbQIj5W//aWWy7RPO2MgXjMzmWjAs/xE
tSeP+Jl24WLU7Of+YycL97p56XkP3mOG1LSZ0HWuXgTH8i1NIVaG+mr/VQn7ZQuX
0fs+rofaRlQCMtd1vJ+QDsQyec/jjvKxNqPNTW6dLTFetlXvacPPdHpTrwlWmOps
RLOxi7LCjzCsJBPrx4cSsLsnOfz+vj1xR8w5VZrXMX77mnIbLdaocBbkEBOY7oy4
1vi7W6E6lIVhvhvSOnqY9G8cdYl22pRYmscR6QI5wVRZTDbJgO38whnTlGw1f/LT
z0KR92/pACyFBhDKVb5EzCJY9f06wL+I2aOt+3s+i/gXXgKYVQIyptikwTpBz+WX
KMJicGgp9MnqlIuCy19mvYC/owfplMNDtT8XjWT7LAtr9eP9jKC6p3ubjh95+nXX
x6wfWvLw8wakoOhHAUZ+cAvj1ENPntyDOYnnp5XLS8C5RmZhkQX+vhqCBMtGL3SX
cho3/VkX6OoxpCdxFJyysYXXqTqw3O7gqGYGes0rpWPOlbQreToVQUIDvxvQL9+c
KZTHNrSasSY9CfdQOmaKizTK5h8Y1IX4u+obTmMeqo8taxVdvB8P8c6oHObfY6Z4
uHnudd9l5ZixqEMzO/7ont1kvRs4oDxomIdcGxjb1VxmhPJ07gwydLD3LMEWoBR/
zzT6S548qwk6H6pBD/RBmni2kjGUYD8JAEnFVLoeERXT2+oPB82Qw8DQoMpLxMw5
2fTxTAPHgWClC/MfrxdYQ0U1rR2V4mYbW1T3c8K5JkO3AQy7LArqEyZ/c/TMug7b
s5gbhy+Lbh0u5EZKn7VotpC+dVBjgI1lEOfFOU3haoxgnVwD/mQI7EVmLfac8GTl
+bfrXSufHEUFQE1duFbnLnEaToivO9rmx8/iseqGNGtSbsZtjyEuqEVlFOIQhieP
1vOS+iV6HubHNaJJ0FD9DseDQN1ZUifHXvfZNziFs+wQK1/VC1/+bgA2XjcZ5ed7
LSW++wIcdYa69JOpXaRKVrDiz41NzGWg6+FL9+iLJj+17c2p3Xo2yGEWDPk/mty1
/YqayogsmjlPvtOt1D1y/Ixx/i/mjAL/P/H3oecFWZTYt18mIshrpMv+ymrxb6CR
CsW8zBu9mW411n3oKbijghpiAdEhVNFld/Bo0be0Sx2vBE+9AuYRhFrnEb/07yGY
l3iB9gAS9ra+S75I96KHkcb34mBZcdqEMyk0owN4SNl/s/x2HDFfIsI0IBxFcecf
wsU/xI8NJ8LovgXGhGo4cIERFWi65YBy3OkHMX436KTy37Bt72oWMr++flNohbsD
xjLo2ZlzqQw9SYBFJrxONdvFYWeRitVpi+xcJxyu+xxCWPs2U/t4ggytkTez8Wq2
9GCLP6Gz8FiqigjGLaQ2P8lPbuocQoqLrIDu2HJqLhLrfRVQid4YjJNRCPyBi92r
pQkw+UHXOByeIf78dcbDGd9dkOvfJSS1vkNBekpRN1yEdFby+1cvp81OtM+bxuha
VQ0LILf+UXduHdTSStgCA5qB7uLEe+bSIOZheFTufYXDG1DttxkBgpLslyy8NEp+
aCJgJyq25i02R7lWIiMfCdyT4AWCbsM1cyg3zefcedk9aGCVFcc8+4UiA+djfTsz
hNvXvitSxj5NsemUsNxj8jt7FP1cF82nZa3aEKAFdSsAso7Myq4Y4O03xegazL/N
GW3JGWwau1AnYmuwmKXPGZ/WUHnyP+f7klUxwp5lMFK00+TU4aNnwxOSbOQRh1pr
ZCQALPTdsjIXGJj9Oh5HxEOIAf0hJG+O/8m9qlk4WkIKxrJN3HHV+2fhdYHrX98f
uPE86HRIO1pTSJCBxQ/S1L2ZInKNXLY0oNkngWHrtfKPx8RHLhqPT4vllUR5o6ML
1XWM3CCQnJgfaNFUowoZuEKzHEnmvB6h5ljvz6TDNnniaThgK20RWaE4gw2diovQ
d6hkmeNcWJdNtBP0PfW4Rg0LqSRY0O0aAkDEJXrCmDMxLp0EZLjPlv8CkTK4Fde0
hay9EtmJnhI3cgB+j90TeN9r+5pSmgW1VZfMC3K7HfbwjfhtZxvlnVNk0jbqu7lr
EWysa7AJJ0TFc9T6HjQvWARPzzVFzt7sEAEiZqdLfYxrQpVPDB08K/gOQmX1RwQd
Uwz8kSXLAfkXZwlyKd55S28y70jEpQ6SvrnmVs1wEGQgBApYh1GUnxIg5RceUC4+
wsihpuiLr35pvocrtvHyZJvd5XqcuKxOTcCak9iB2/3YTDBCLJ82IYRuUJ73LjoB
SCPHqXMWPo1ss5QkGH9xMZYOFp7Nd6q0FF2GgO+kKcCt+KIUOmxoB0Xe2ErDICs/
++yxy4yOwltDCPus3wZ5gkfw4XzrSWOn6efE/9g+iBx1GHOxAkSohfpcWwwH5W3/
y4S1Fl8ywyk7PDLqXWmyAH4EFWwbpXpYP2tUvqJorqSwWIBqTEC2mMCnXjQHePEE
j7+0DuqVtVkEAoNHCon6772bWOxzF6tnkhA6EYpkfCraO17LxrVP3t8v1KfP6CKv
DLk22Nd46dhH6sjZImymnh/wfqmK36Vk6W9nrvFRkkLeJCGWCdkOtrPbo+jKEnLJ
uLPPeabqF4ONvIXi4VxNs9ghATK4yBzQa5INlp/5+mETfb28WGw72tdrMaqH9zih
1+uRRszYY4CyDNAWJAwGq4c3MgcKkJ/CVkywHI5MiN3QJ55SfXUG5wdRA8aqrrRV
DDkvyLsxewEx55HJeXZ0twXVw9v/IOgRHEagXqpGON0MZa5h4jgxYY83I/dKSEow
Gn8BQPle3JqSwnAEzdptCXv4/nk1aVtKfYyLScLr+0bA5fCMjXGg9NMn6t728MLy
DaydvNq7A3HMx0cwH5XaYEsX9T1lpRRaBERb5EmB3dO5zDQespcUHq6Qzco4WPHv
VpuAheX2d200t7Be5AEwt7kQli8ntykjyjRQYjm1Y2xyihttlCkuqo3VGqNmNyW7
qC7sH6DEpp8PDy+v/sFOSvABc+IdLQWg61vVT+01XdH0723K0DwJZrlBrp1mcTkF
w1MhtMz8uNS5VpaZguioYirShhOO+8NB6Fytzqa6N4QvYwNtRcY0QsAA6pms6Fof
S3YvRnQnJEJQrw29Sp7gNWad92SFZarlHOapRvkECY6n4tHC2bDVQZQNY8KAXa6a
BYqoQGcYJAuleTjaZNNHWiQsC/WeuIUnGqTL6bhC2bCnYDcVEe6uQOljR6zadNr6
mQJrks/f91AwlG6dySZ5VYyWtqz+94kq73Q2VxdAKuFcsJYZqPZlVhL4aMXc5IsF
+hcso01AuTkr60blZhIvKW25tVr825HjI4l4sx32eQAsLPq6mtW54mi8DfpqMdcq
EqIJeETzTQ+3y6hZpJVXczLWRI86MN9cdbNYytVDhMVqHM+lIDO1gbch5tYwvZxk
luwtw4fFUBNGyyKzTWWoVWZTsbB9YwdC+gNaNhm0JNm1juQd76lecuwmkHloAFcu
wbZyrfYqkCtWPbA/7paD4k7mbVOUKBBlpYh+Pu+QYQ4mjp+ypLQeabp7QXWm2NHm
Ds5KsqMiYcafA9h1d57AWkW9X10X+cXmy9G7w1467sxYRf3j388RwFti6wM8/5Fz
mkWRIBrt1FO7zwgHj/APXcCQCw1XGlGsdzVcmMrw3GQMCDoeoMDdzP4DzSDpGM3Q
YzTGX1/h9H39HT8s6AHwwtUkKCmCjqqaDsqXrMF+tekWWFXJQ7jGz+liYEUQxHdL
3uH1yk3BGWqKgQMSGoaemV28udPJeQ6QvGzRz5dLVvwW9QpRlvVCcxj11beY00+R
gBCilTPRE9K+lJCfEU2uu2u+19/TjMkgt/ZJ80WAHnRc5xf1LkP69gK6KZDM4IuI
pTnGFgHhk0Dh53bbNmr1q3wOnQyAjHIkJYvjKEAFvHacsIDinuI8xXTX8XTKFlor
Ul5rvXvN2enet3drUUoN8isO8VoawxF3gaVGw4FxWAP0L9LlbzJSCnET2ZczrEDP
GoVj79ndoEWgEL8eEIXqxo5S1EZk8GN5zw3Y4UMUMz7l8+RORSVYVR+uUVcJiAw9
OuitBFwAC+UOyaLOcUtXnwkGytYw4+2Dg0WfUatNjXrwJunnqCIyeqopyMT/fhzO
Ebc2pOnSfRGDJg9+qPVjJ9+73suq/an+WTFm4W+fbKLMY5joHDxybKcnEwvLgWCP
VK9cfoIUPd3mW5ZdEgD3/WMcU6QklvOeutGkhiDHoyTn8y1ugRruDDhQlr6zkmMs
mDxI8p9nbWL7U1yPiDYYZJBtwJSqMUHlQb0njItND5KTxTkPAQaXQQOTyw4S61Xt
caA7yP921Xwb9FpBtoscWZxEia/bCAOjhD8TyuB2xu5WxxdNXoqU2I4C6b7PRYjg
D/f7VyhUkkcnmYD4N6LhuUnNAQuH+YOxMZsH5Hvi8ZCjSF/UgbnyPvjAZuvS1I8x
uyTnCoPAKjcXBDZG4pjgoUtSydZgmwbJU0wWSGa8gSUeSZlZDg1BrwQVhWjzrIq/
DV+dRqfei2VcSq0FXDwl4euXCtLuS7rCZ+61MEpNlccCDenMcSwtwT3d4zurZoOx
aNXPYHoC6jcLL6+xgzbseDXJ1GLaFtciPDJCnHvpBed2lC3GYPnnjkCaUPsX3rVj
kw5WVIM6aTwKJzwBPmd13WDbqKHgWj2pz/8Rns4VCS2pxPf5lals0AaNE3/N4EBg
Anh8gwlQadOInxhIGPu370nUWHwHtD5eXdDmRFJcfEXw1QCgkKRFzhwC5zIIC2dp
zJouyt0Lt0LtHxAsVVV37sDlUWL8RcorlNgmLmA0St/LoHiMdP+Q/xcFCISAuckq
0svCZbIpqJ7u/TGUVxLe6BGTGocDoTDZCcLKk0HDZ/10VIyu1/+PDWyXYZuSScnl
TTk4b1k1gkob5LZ5/aDeteT/UTqTi/9YhujDimhCgr5oUjSHH9jY5O6cD+qVOpaa
HXOFiAfF4JKYcmurDPOV3k1aAZNVLaJE2DZRuSE81HUrhSEudscOAiAHuAaOL9Go
FEQmHEOEXM51cQ3Xb5MmBcTh3cO7qsdw+An2VvefXz4/NHSL4MX5h14BKaXN2VXi
4KG7BNG8p7fSPLyr/DLMqzPe3PnpsNUL1yszNLEtKGahLO9SH3EOBpn1d4dCF3Bj
Etv+wiOZ1oRrxnfNytNfsowXcXWTKHI7BnZyjMHzAaKfnJrMumcxjGdPcO0AwArt
OPcnqDtT+PxK00w9TEBaLRL62cHN/UNNC0Ma7lp4KbdpwRsAplVz/fOzrjihXomZ
IbenCUlJI/oipHjLnLf3/5UQgTpTJVoHlwDXyMbdjGrDs+6woryqirpaLWweKOyz
3J8lPE2G2Xk+GoUtOsfmIohX9Up/Jys3Uozf1EXWgyM95bOueYVaXP9clbg7o78J
eXN4maemxMRTf4+6AroQo1dmYF8rLOdID3zfKe+c0yLw9MFEuocZS29k/7BYxkIY
ne1H/s3RLJ1GIAhsdVU0gwrIdvIZOeb8fl+U84Ndw4k1lV8CiagzJwCjCnxka9ll
0FZFyS1cmONZbZxOYRYApwij0tQIzl470NXGqSvpTIJJ3VmM4tyfcOCb19mqla8z
lTFjzgkewM8wAR3hUGB2QfjAHVxB4qMwzhUyQq/Q3TXfTS1uB8/e3xcm4eOZQhfk
03RbLnewqrJAltAVNwAfiTU9c1T5CAca4yG6nH5FfAScVqRuRs66dTF8cLMOrEBC
6f0ekRMnXf58Un/QwMLmKhMG0KCm7360525Td48Dd9L8cZ/OO8fzMPrUyddHAKfJ
/vPlQhMLrkmGYVWUBps0Pfi3pnhB087HM8cHMcg2xRIUMjPN5zXEyWJFv+YZ9/3D
SF7EgIuwraiKsMSyQMVwG93txcB5WKZL0w6w1VCsJ6wsT5OZPID+pxwptNtZtZzE
RQy2qggH7WYHlr474sEQyKnFjbfNAz2aY1ImEWlnf7ObK3E75IVwm+IpHOmt/QeT
RS0ncUuSsSerpUEOsW1JtVzEXoyqmdIY2dVrjJXN6Q5c9+KnHxdC/zZ1xeu/1iWp
b/eXdNEupr1C8KbPuQhcUJffBn5m5zzceM/6KE3ecKDwEBgV74A5KxBmsVsuIRF8
PnV5fMPi5x9pl9O4KKqz07fmoT7AvStj0jTGue6FBHikDllinrQjmehNbMfyl8ej
7ARbWq2BlN8zlE8SCrqorHmiCOE0/jcu2YiZJIQ3Vk0lFlJtjObwK4kdrpIBJGwQ
Xgahwy7IJUXPlsyAuBHdWBPJ4SKVeJN7lDwCZszzRPXVDORef1dgRRf8PQXKC4p/
LwabyMVfGdv/AYrlCMEP7yK2rUeO2i7vwwsQSNY9b+3LCfQC5fon6Bfahomb/lmK
yymBWBJ5B3JjszM7gmNiuxpYt26izMDbHCMuYULJvYjfZZOtzWnB9VTesALtYfU9
uT2PKqXtCqrV7e5gi8lpcZVptLLzuI7hQukjjcA49G4jQGhfzZkrr0y/IdOB0w9v
Vh73Jw+Rz1Qmj2BKiC4y7FycxwYJjQ1ULNWZoUEzcUBYuBOH8S7XUsFyYnRHyXlM
AyF/HZYm5OaLpksw0cgjFrBPFT+y1OM5rEmPn0WwvEeuscPojMvITplR9kvQ8ABC
zZ+n9nSqzkkKv/MUBx75csSDT/DFneFQL6L+n8Q/+CLPCl7Bfc0HihHw3pZhRtGS
Fr3l5gu+WFzu26nE8CQqtU0nsjHHLcQ2of1sZZQeUzoa/9Lo3umqp7vyIeTnXvT3
V5q90bDnf3+bKQQ5EPn0lCi7VZZAxyBI1+Q+igYmgcdhxF2CT41+ZCNZwWTztOJZ
4CKWFy387rR5R3PIUdQG4S2gf7web52VAFssIyJ2eR5XeA5Lrw0XJwr3XurqvxRP
2p0TnKNNt5a8tdT7QBJ1ZBNUHklbQxW3y676zsUJsGhEocJ81+6EQ6/vB5g7v8dQ
TVwQM/4YjRBVhlIOYOu1dPXMHlw26b1AxuOdOgrFG04wC0hQ+r7pDoQF/jJvkyEg
9SLWUGdYTAcwqIoauV7BkHSW90fytCdwvRfrD5XjivA1hvL3tIu+W/f8yL+sbiXf
izV0sVFXdEHWxcavgC1rdRwW8UfNh6PmjnKjiWdx2uXbThKscwXLFsriMBO61rjz
3A27K1EF57R70ynRlhyX/tgTQ7h+miThuyp1S3c3FQw35jYYKcoEGzjz7SgmTJEc
BCPY8xCfrdeLrjOZvw7oeVFQl4fEFif+fcA6SvU6nFSRZ4V6+07Inw5fFjGr+qIk
sJjk5oj++eme7BHKPfujN0T0SxE37U1f9xUCcGnc2ENLbq98TafT5qBC+SIs4cUH
A6X47lQNGAKtass+IPMqSj2rgqE/NPH6+2uxoMChH+on6LdfCOteabIvHBjqUmOo
zb3hqRexkruDDCjQglXVLLrRapbxuWrlAZBdh7rgTJ586CIfJjZrccpfHeV+jm+K
Z+ibwv+PeeA6dQraXE662A4qjMk1GqMqooDPnxCxWnsHJP3vFfvkzucipav72zXe
OLVmNBzjkPH0Ok1KKrOzYh/3MiOlolwMYXI9vH3a+WXtskM2Yy/KuBi6XCKZgL4S
m2CvLDAc0Isal3vAwi7r20EpxCx/1bmDYjiERKwG2wtgjUYGXsFR3sKiHRPO9+Xo
a/FLcVVtGDg8xEAzC2fwH0tYJs/KKXIM9veUfdeRMdPRbfJHJFQaNlX1p6eODV9y
2kVae8B01WsgvzGT0818SFyy25W91kv2Nd16OvaEOW1GUAHZFuA/+spksaBGspFe
l3bVsx5EoPWekkW/YMmT0vADq+BhDZ5UuhdbQYl9jm/JOdwhpAXeAbm1Sod+Kiw8
aP6xqJN2ivdd0qlL7kmpbW1ihApVElnfL2aSg+rWl00CKuTSDIKAXQ/36XiR1UHX
H6HbWjMLRfOkjdCLOIsQePq4cnqqRbr1bfxdq0GIF692fErCBY3Lo0iJDZofQiGE
kQR2JyhjPbdVA+KK7Aywv318cKJr6d9mCf9SaT+jVnLYHuExfQ/erE6TuqlL4ugd
SbrG2+QgKmmUnYVM1zUmiVtZgYYrA4rGnGQQBrmN2wRt0ZKVm44GTteSosEqRGte
85XUIGUYqX7jrY0tXaq5txA7REaU/L0oZ7Xnv/BSP7eTQ1MNVEWkOQScP5cP23JV
Hh664+6/EUmlQFCXz5yjNWVzP10yxiiyiIZQUMReA8rJbc9a1Texn3P1o9yuLSfl
wniMXmHrt2tbMyqmKnt4JRqnUmDWsbZbsiJe/HDryjxQzPyBUyyqCPUR8dcomTt1
a1XXYE9/A0VsCrrvJc82/NGQRVNuVH0WFqEzjGXCg6GUNLy+dejhv5HbodEZ0c4A
TuONbOQaYlQiupQmeuimCZVwxnhsw7Gjc8KxYQ7SBZCpbuzgKeuKnA3h2w9YcvdQ
KTv+o8LVbLQivvBvq9kyfQ==

`pragma protect end_protected
