// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KZeV5GSkVtFvyaRacTkjLwlioz+7Ezp57MNZp35yGy9u2I2UMIn4XEd1rKMr
gxRIK8FWZrKrw1YZp7v2/+hG+/o70ct6MgCmtOZqNLn67geSBX711E2Mex87
CAtZbsoFpbejap9abFB02iB9kD95j6oF2TXy94qjh4ZSjQdJlFcY3mn8LeAO
bhxkLc48RxqgeciF8NT2cy/Rvk4ylAT5u3r/7kTi6VDDrnBaFXxie/Vh5NA2
pGLb0HGFFMTDPQUX7sC+y/pnJt8KNgmXk8TJk0VcDwRYV1O4MEzDAFhtS8qT
rKP3ynFOeUjYbsj9Msjo35by/OId+qUsl9TFy8/BCA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
hizCxvoiTPvD6lTHCXb7n83hnfMfL4FIqJX7ynpbuGICi9h6GjE0iS03WkhD
eQbVCMu4b0Fv5FbJITOmPiXvHX7B2Umf1Tzn963TBAfIekNyfaOhozjfDEhh
tzzU2TdM/bRRwAMS+/A7XzeLPf2cEeRQSFpFk4Q5X4NNF2D4iATtEwpBtt7M
t9XGk0+SrGep21lU5665Q8aIV4YxeaqCCmYfaCY93y/n1G5d5WxgnYGMYG3V
KepIQDZPoBF9kISz50uD6zsI1SzRjRyMgEI6iqu6nTon8kI87vrMwNMaz/tN
8uPJOFwjwz9H9hIi/4gLD2Z0e7NQpdZeEm9QATVF0A==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
MuK93Eg6iJVxRBC6NyhctEs/mhBBwb3q2ObUGaCbWnldWEyjgUW0phbLQRWs
lbHOe6DeGq4HIj8YTyr808h89mvdZnzYvm7dDY8fPV5xXayh6OE/96/7NaV6
FZABo06bO9ZKL5Cv5diynx/WMrQ+0BOqKD3NZVr6v5UE7a3x7uYqFQmas9J8
NBXcrdpqJAEgp9hz158qbxwhw8wfDPuGJNOjEPuIFWOR6k/dxNWNoBsaroIf
gvuYg++LmgUAfpiSeRcRQuzs5tU/+WOXfgPI7/zm1qe0spBKXqHSXbqssvqq
Ye7/Vxg8kfni7XP1WWIAsbpByDTFy8r/Ikus9rQOwQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
DckOXcW0Tsk8MgYCRbyHgWdgyc8gkKiMF5I6Fa2R657jlSDd/EtRbeQ/Ho5g
EEGSTGD3QMx1wKH7QjEeqHd4ZGB2uWN+IianZ7h8Wf1S49bcCG1QkbpzTbxz
ii6+6nj/gFMgqY/9h311CdR5w51ymjDTuKuj2AZB2npWAmVxp8U=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
WQgZQ2qs/yPIyMH2KgwB0mFXg4A1CrK91tCeUbWjWzL9HYCeiGOiZIDRrG9D
6QbLebiNaTMqVv0ZUy/HH7T25Lw6U8cFiM93Y2/J4dpTZ1yiCcFnMGOBDyTl
FnIMgz2bWGpgSaPdM42tVIwGnputUAP+HogqAJEz+hBocxHyuX22H9DYg3fz
5o+VnYqYQ8DAZLj8g1EgX2ViU2lYCg7FPBghwiqP1MH792NgMRdEcdTXHtyf
AqsCBLIc1Qwd2AfMjJYIMbX6hKF86ysa7VsDB2XkcopL66nOyi/htToOhYTx
nEUy6HJWIpLF2sXkdb8v5RXVVCHOIwwOqMhJ1Erua++P3pZRrMRi42iyg3cY
D5WLb9NfIdzDsHQLzrX5TiPHCXElQOJuzAQBXDBr7iHbNVqeQbyJa18wr4aU
hqwfa1PkgUrUeKYjMHJJRtasPB4PjKdEuQmjycYrpLd+k6BmjJGDrryaWG3h
8DUjWAAwps4TA5xOfk7sLXJDZbo1aidu


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
lt4UN0hMGd0lLJEP2ubNK46SKHX8Jx2pkTo+pOMTfQ1Z5Df5i1dTcT58Fzf7
YrntZcKUbdz11cHimWsRbf98Dr6ycHeyda/0z11+9nw/X/yOY8RDJJhbQoBg
4iRfkVjFZbAGNBTTxt5xUCxwkfuAfmPGx3KDiranA3qStH2jURA=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
uaZT00Gw3NqhwtKRsFHmFWQJc3p4GkUMG0AzxYToobW10qtCAwVL0U4S6J1m
TyRd+syhCmuigJGQAtpQOP8nPmJh2Gawz9tdMg7dqraE95RR5vNa7RBagc8J
gpby/TOoUZVawrNVpEIC1CIpzeV8UT5c4KGGsQIjuUY5DuIgl84=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 28656)
`pragma protect data_block
FP4kKmRQTMaYBsUOFLlokFebLPFdTu6j68RTYejJCt1c8M8lkc/0fJBB3nRq
zqKguqPmWdE7DQDcvNU5J8UIW3Q57SBvfjyu/t2OEi4xZETLqHibZejWQhP/
f7cdTBY4VDP0QJsFnJmn1e61EHBFsRCjBPNTx08evHhJYhGUKX3z1nfzz+eg
UOxhMWHH//XWv0qjYEJyUY2JbZCcjj9IB+xRFLC2Ocre5dz2ek7sYR70zjyg
v6zrpc+Q082Sza6LF3DD6MdksUzlF4nMS6wLzc3fKlPRUWjTkpp7/ZFhfAoQ
kDI/+AGLxSupaU6j0dt//VAKALbJXdmFbwhukBELral6At7Fe83OIf86MCNb
cKBDq65vdHmutXL/vWfFNt98IAImXp+90zHmKZi9BMqCXHWWQjW8mxXgzSFi
LalqsKPwvs8VJYPlhF5awxKUkneqROit+IZhMZPm1N2eJ1DXDuzGLWpCFabP
1VUhZztjPS5yClzrALrrXtr1fsZl462Cc+D8kbqDtSb8EkdWv2g2H4IfTqr8
Pghm0g4KHM6K49oY/Y2YIkM46ulZCLwYHV9RgplTYcUALYPGNWpLKfU8t7Ic
ostHxKHJRxMY60kVL5tP2VeCJMzFUSuh5F1PguQwW50pjHfMmQ66Zp/KLhr5
U0iHuYcg07U8mV9dvfWiEehQ7k8AH2o2vIJG/tpehk9ottLe6c6L9yRCBMzq
6BaPoQwBJRAB2jErTr/FLbALaMTMbF2qOMRYaq9FBth9uRVu+aBh0tzNqDHj
8WtQDyd/EKHSiMF2I7MlILxfwtqBiRlkb2i+rSHhJmt24no9yYn7O0eS9QCQ
5bNFzlw8mWExArgF2AX/tj3uQtU9nrRu6QfcqsKud8Gl5TAfRYWWpmTKCZfa
CyHGwr7xZFtsffquv8IiTkP4alTFmmyiJ7/6YuFEt+izW18syIKIjw5QlJ3C
Upx3Xf6V16tk33EWTBHhVF5tH1YzY0PlkAJ313qHX253+XSBWoRYMQQuA26l
/ULpeqpU+r3wqJpPFsqjugwSniXz1OdQyRSDC+HiCOFGGqDa7Vgdnqp0R3lh
geCVH4G5JfnAwy0BRfiM1y9/COcvocsg5CUvqA8Wl6oTG8O8cQmdRrGytxLu
X5Ww0uKCAKPH14o9JRRuVisYFOc1yy7b2wryrySUs9FxDcE/iWnhCOgyEWwp
+0wJwbq/lDp7H6avn8cQWzQfCRhu8dmjKlKA8jD2z4Y25KuYhZsDqTkQC5th
bLARO+ZXjX1DgCsh4ibC1S/SPipOJt48inA/DRBN/GOsVcDuh/bUsNu2GkUX
vpA7R7tOPtqRuKmZtuX+79fT6lr6fAXUhLHtk38Mh/EbU5i9o61UAj2FxojR
2gWsloxLPPjUTKpmopNwKqcK1cL1qFvljJz4AtZ9se03z3uwMWjshZca497N
jugfE0gPGUBe/zGswSiNMvMxKno/eqpyKIBzafiTiNLFGzm8+CP5EwF4aF3m
GdbFdjJN9tsHB+NuQL28H7xTDr4tZjRJCjnVBNCTeZm3SXZD/UPvskkKQNc9
DDpdLbNmx+4Usmy5wkSdcnU+gnK91kIPbYUpxffyXpYbfRDzutptm+saiy2a
BwhYdc763mlFwl78pcN+B8o2uRbU4gg8zHTaZg0y4RMR64C9zcDcy8dcBL9S
Gerx3mDOZw0V/XjfMH0Qq3d1OXazvAtrIqCT65ooJkG25H0h+I9316OAR8vl
06+Csxa5wc95yWggBCGpHYGm2Znl6Ro/jY7rdhjoa1q6J/EiteZgUVia4Rmd
EOtBqgp6qpjBuyISQPqBllRTqSgZrqi2DQJ2whCtXXy7VpUf0/q38/mT2Ru1
OtfRTrOAJT4ieZRB9R5yen24CKFoJ91AvnKYxyz/yiudtATw21KEtEYjviSA
5uPj6cLuHHjUHKz3MYhUK71CAc+VtNUYEwKge9fovEUgMqJ9x1YffbpVglYe
RlBMdfrTnBJsS6IFhPIDwlABE2KE58jjvIWmlbAgjfLPGbQz2pFQSfa0Y4uZ
VQIMI9H1qFZRzLJfqUAOSqWYcU9ayafgSKqGEbT1Awn16RGy8TSURHC15i6w
vDXwGb/eFgzfQNLcqHkGSdIqQfh2i8aOEXn5taNd6E03kUEaUx+iLW1JhPZP
0UarSubl/L677xk3AxVdBvRjsXu4ISE7pnsLK1YHk+Vu722XYMfftl4w7dIF
t0m2fB82V4uuCY4YtcU6JEt24Hy5bmVgIeaBOveRhmOd/Jrp3TMEaUDW+IKK
tiB1k+PlYisTyyfiCNElD9AtgsPgLONNXpX1UnULCEmwBr+qL+y18XbsJ/83
4831tzU9OtWgl/bW8p27qFh3xaZFFyYBhVXPfiJQJ61SXzZevot6Uan0+WCI
HjTaz5GeOlkEKyBRBSFaeA+556uhjku4Jk16mp0El1FILDnlCmh/DUPh/b19
HXg85X8St6dgX/AIAvWwCNrkhuEGeswA5s47AKa0/sJu27O8wKWnF4OW/WdF
t/le8UOH5d1SNxVcq34GVKNQwP2FADu1hwzqyslK3CFagpEnk1GrHMy4vnzW
e0luMr2C85OTqZgMtrBdxupav7FwfyiYCmugjjW3vZwWuIC4M3dN8fGd5//j
jGlqUs+uv26jXsqm76vzAwYTXJeNij5rLtp6Lu7Uaz5Syh9/JadJ/2xR4Swp
5Oyh+D4Vzp8Z8qlK7VteIEfDU2fUs6vnHr9E/HyOxQfeWx6cNO5iTDb9mlV+
yvHl5dECtohGgYC10KYNVFOE4K4vGa9a3erfbWID0YlAH/nYE1AHd+8dytYD
0R1JdfKO8U1zsuYGrxgtH9iHhGBCRU0DhAoH6cR5drhC6p4KZWUQGDrFekQi
7AlMGr0BLFWWz8yk55Egst5ZdCi6ox3zZEfTBygtCEDAo+f35StrKyXSWZYC
B6mB12yQt552CE3BehIOy/0Orf2Kb2YfkME0A//W7SpmgWZMzTSorWkLn27d
ZH6AnuK4V5deptT64a98oLoGF3TrHBI4JG3gPIOygQvNCj73ekqCPLOWxiTb
PHnOolfBwoRCJczByNTjZCnSUiGY9TcQiwAI3zDHfqubEhxP3xhjpsOewlW+
lNzs8Zrzy0hZJ8Uofdyjc/AtnjFVPGQ4tgLiXKVOK9/huzzo9+ChfiDDTesM
Xc7MnKa+ulLmFscrXdhYqlWpxUayPmba2pLle8ubawVTvlbNwdju+d30sEQr
cOs0IbHl6gY9hamd5bRq0JF9BVrXG1tRH39oQmhxcosGbWFt38jrQdyksgmD
BbeVMjXJ24leX/GPYi4hqytgFMcP/fUQaVgIP01BLHGLYgI+I7tVHujKlrSx
9W+5FYAY749X0eL+OPT5q+BItZK6hy95RQklp8G4RvVBSa75b9WeegZNPR/V
HHUoMxbDcsyPskdjL/10EkW6fN14uy4kIj3XrO1OnrOeCtuTvLGfL4FWE8Pk
1FF+Hn2njMih6V+upIOL+f3W7R+Xz/d3FykTRBZR91wq/2yCG1D7O3wjL51h
+M/al8yvx8FcaMG+E9ZKJDWg1k79B8z9uRuPPmOZSJr3ImNIv+x9w0aYV7Xw
yka2I/60T80FOQBC/K+WKCDuDuFjgo012jsig9CQVO4nyBG9ihJMJoz2PZ+s
VvvFiAdSuG5hsU3VoYKS/19e6GyAptfkFHvyNZmD2yvKd7KrlaM2XRuNpLC/
wQ1jnbqTeFeZJq8WLvrkrpzOYc8+QJVFCXzkQBnXTTkMX/7g7/cV11Us7TQy
hU8+QSTuEwWjmJFuAmjpeDzgiznIBYFbmi8eY+bROClJ8F4UXEIN8m1XnLjQ
QkkvfrJnDgVAXZrZBu4JjRIiYQPz7XqzLDQpD0FM4r8VY79R7SwRtj5bhmRg
IxIsiiNzH46+P/g3yFQdPJCQH0Mg0f7zoTfMhjjhH7BRZyZOIl+pge+zUUDT
Nstb4bVYmRJlSrOwYaMXDzzx5dMu+PqJLu4WRJeFwukDobU0oFZHmvpKZm1P
vFoauWYUZnD1xhJ1x7710xUwxJvMQcqetfvfsqPZ3dyVjJuJQiaL4cN68shI
emqvBtZ9GZdAQqaF6243Elli4PH6Zn/gK7LOFPpntCAacFKmdz5pfSNoTFXz
lmUgb0JFNifzR5c1OKbf4Z3+xv0FABD8sfTm47FTQwuDLnVISsQ8dbsaPmAr
vfI3R5HdYD6IdHEYGPoVaDR3n0Mdu1CAjs67MTTT3G18diq4uV3Ez948WJOi
LsbWfpCMlNeWDN3+DL/xZmx9g2pm1R94doHcXmJa3puZHlPS4EUYcFsJwVP6
0uZ+rPD4evDT8ODcFJ0SuKzdajZM4anAr5HJHz2WUGcrjlZImOCwJZgt2868
Bfi8pFBhfIwXuTe2I51SxHovvkwbBb2TrNLhKHdE9BvWMRJbBuCQRGr6T2YA
JhFePktFBW48kuNOUeUrjgY7DBcNYis4/BH+zoPwMV+tVETcoJjFYONivk+i
VlzvqbgMYcPGDeWbmlZd+anvJ+yiaHqijVWdm4wr8ZbAB0YhGYEEfPNKJ0m6
Os9vbgk+tE0kRaiNllrEGvFxHqmwz7F4KTkGqQqsVF+o3Yq7pFNBODOLE+QF
nU5e0KeNcqYNERsGQmb2YWYJR+STyFGbhzNq9p9zNHwb5qGOsyayUHScMYec
Y0MEUJMkH9AiH7jsF31+5O8ZzFA4UICx6KuEDR1OwVfBlAston02t/yHr0EX
pCRtNY+tibrQJHBWvp17DtTMh60BMeJ+8yBes38OYcX5KLPJt3HhELU4RHyr
JxNT+S//6RG5ovRpoTy5A+zL/PiKBUA/pz6Eq7XRBG3vMJfj1NIxO+sGyAJ8
KiVANBcZ2y796NelqA8ecL0Eg3szCCIeX5C7A5yj811KFckVAUSPSwIu9spB
Ab9BXb/Ncoh68Cb6/MKul9unCTGZIJGwPXN7X4xbE5n1obfydtNIyDTC1DGc
KcD2mNfshX0jNpHPu51pyEQ4FAzPYUi+WmOSlH0HD1R8ZuS2+LffzZWl+YTB
hrqAJsWfBug577+T+Vunuh9V6/A8arK8j1/Xgk0DMARE9Y3b+CZYYQyTd0Cw
LJTWA95+ZRBxNwDCVoLwmWVeGUAi+93+0K/FLU/MsQmtEUXuTub1E1YvG3Pw
NKMb1qA2ADVnbIT06T1SLAvvHHSx6fT40ZWRHg+wmsuirRzZbR/4/gvHJp67
QHOw/LcdyCKuSSSv1+XNo4D8jsfyLzfZ0ysb52sEBLA20sSXh6st2IFgJmBz
yh2FiumyoNlrmXPHhuxNMgjrjcwHkGZQRWNF6bMWOa6ldWCrxN4ZoBBAdR2/
Asw9FHvIBj99vBhJ8IDBfcEU9I3oRcRYnNB9Oud7+w37ARnANrRQ8terkin+
HfIcekafSZX6h1zGFn+km/NpVEE2EkgJ504ePU0KN2yhyq9utftHOPA8sLC2
ma8SgpGf/9iouAQW7ble9rxiovusJpZG2zUwUIZC05lf+MLjwXkdTIHYMlee
vj/7NkuNEmWtMTP3ovD8Ws+9Wc1+gCcsE1DRS30tHYy21dieqgiRRJI7B6we
SHlM290k/8AbJaeKCF8knhzGjlmEA++vO/iUEgVsl4RIxl+Y5CwlRe0xDj5Z
IHHE4u9+8xQrXysJjvOLpxrSeamoKq3e5p14uTsziHAjki1yGjRtQYyIJFMn
7ZscPo3UOecrquMS6Nr68aRExJpScEi7mRIG0i5MhGT1T8OXMtzq+nS3frj3
LMu8qMKa2TMLfRsx5QyLMe60K5MxoYmd6Pj5n33bfeA5ahZZp0ryYN9i4ZxM
6aegNtLUrOSeMHzVkKUivxCeolCKlXZoIc+mxTDKLy9S5G1YHEqxxMdJ20yT
RRpOA/72PICo/p9LGS7G4VLjhcU6q/dZuUWNDTWcLhz/bz5Sz1Buo+9dCpJQ
2AFYJDemmEjlIMqpkC00VnoxYn/ZQ+dQcBvmobGInqMbFA/HdZkJ66rJ/gWb
yJOOEzyUvZZuwpEYkD+cFbKV8l/lPQ8aPsEIsvgCoOJDe7u1fcmZgb20Soe+
L9pCWVxaSPsckjRJG6JPTmeExMjUqp/Y8dJ8Hgg8I5BNJnCKrmsCsRU3zHeI
C884tHwSz+satm83yutZe1biYZiN5j/jCTAR48BSaDgSRpQAkPVfcj5stEh3
Y/vmRvJH3liCoh4Q70VlUqcnn0kc28RXpvZiWfrVGK3lHnahHA/afijj/HgV
xZ4fpy26Oy4WcDjWFe6z6vWmVNMH+kji+ZTcWa9RqzJ0CwY8/9YNeDmnS6oo
3KSP+6YU92iTwWQtbeRHQdtyo7W3+Kp+uyXY8osMe+adzNW/3YqitynEl09f
68ScrOc2friyUm85CvTdLBl57KxCNSoC/vbo2bPob2DYLrxOpwy1vr5CukSt
3Dri9jtAjgfmS/8wBuweG8TITohXMIAYz78Tfz1I4ciRITe4UY9J0XgZjhQH
V+QugllNuAcxoyVgmgXeFwcAOCt/cRxantEDNfbf89eTdLZPPRY3DLlhYYiF
wGDA47JoqQhWJ+bZh8LtyabMmyqYRkuLovRiyPqbz3AtPaj9supgMa/bE+il
D82Mo/6qDyf8/lWvLwmu5HszX8dnzOiwglO6sL7pYsyqHJjROljTYfOVgxrG
CgTtElFtsAdq8vvTdQX4N5J1hqkywo0qle9/kgH/qmvEENmjsCpvyZ5nGyxH
ixO6k4Q4eqJMu6+je56W1dkLvQmmLlkjnLrS/IHTE2MrNW1P5RdTJqk+DEl4
cKyqChxuqxa4F7fNh1wsnKD+uxM31ljYFFBlXcm2+SVETS8Ms2XXVmQFeDyC
ruGLL9ThPIPdORDXPBuRMXk0KRBbvq89k4ClVjXed/NCAalxEd+G3iP1mVw1
Zl9mvt7C/j0GAsS/uYd5tD4cDHroqgCzG6+ZgDKUTjxCqvwUJhKXquHwipww
Pdj7LXJ4X4zhIBROF6dto2Y8EysCVhL0xh3D/qqicUMisd7aP3l7QtF0w1CT
y8VOGfLzzrKFpUV2DAO2iD0ObajyK1Bo+ZswYT/n/diet/Gi3HBCuDQu4+Jf
glICI71VllJAjbDVYqKle7268DWDar16t1rbhHtLHpa92vXGW/xIfwpfdYFn
VRtZpGK0cisg5BiB+YfwCsyWCIxdBY95Q5jyZv3KSGYbdwY4FyKV5DvdsrzT
04QFNED4cJeUQlRphUMvE8i1ilrR1zaMIACtuOPFxKzImnX+SQljWj/Uf8vx
GBf9rAqRzmWjgBFBSkllpPEKbunbrLch3Z7q6npcv1eUh1Xdwk0EUGMGAMgz
o8uzjmxlBzVh3h2z7Fb8B5Y6rDvgA+k6VtsgRRKDcIZDHBhmiK3HfpL7Gkve
qM6uB74Jkib/tHr9/TJbPiUlu5WryZNoShHvgWSFYG5HNdxXJB3H8vZStXph
7G7SDd6QMVpRw2VNJInEftNwVxkKmnrx0uX3xXS9m8E/QaiQbzOPj7VFDV3a
bl+ak5Vrujx8uePGeRGQYVzMISDWQRtxf5yX2hAEdt+bm6REB9sFG/Yz+3T7
By5edcRzhmpeIZfaKd5lpfFRMIyVjjFBg4XoJAdSXyACwZiFyjbyE5B0QSaE
/y1msB3NGp9fMX8tM45B4X5AwP64nAbTcRZGDZH4eLeIMsmVtOrfl7/CwUgz
wNL6wsKF0A1piIKabldpjIqLlJPZyIIOU/jEzMxjd8bHv0Ty1SOIkd865H/t
FFfCLYLcXueeEveVQJC2nl/EOIHQ7vL66kffiEc15OH3D2ykd3DLAp9DB2bw
mm7uDQn7+K+PLdhS9ZrxjgE1yvp2a7Dw7EEprlgpj96Y4GvocTmXNmgdPlwi
UuvRukMCpQY4gFfwvkxB9aKAjlBuhiPauETqpOPmMARMq38nKxtnwtJSERku
O8bxKrmS2xPfXqJMPc3ZZG30Su5SZfB7BKIs1tc67/0qvms/wrFmnOSREBO8
x4vIB5R0pj6tvAUVgQfhUtKQBasZr9hfTDFO8tr07Wg6nk5LwxdplZ2v6Tmc
NsqEr/I7HEi3A1WG7d1Bj+6bCnxFUcsEDWkrtpGBSIukl91DpY2NGchFvGjk
0F7ZVOzGgYKwyGHP41IG7iKQwkpOzzCKya2Fig9MtWa67djjzFnOGM0Ndego
EDYRpUDXMdAMmVcLlPTYIqr/XYVAiOPtjjF+r5uI//1ul200aNIItqeVgCRr
2yCIEXXta60XUTuAdh2Bs4TVQpdXHIvrTx8tYzGBfe8UzJKwOcLQgUUhWkAH
gDmHEmY/zabtm0CSWzwBYErcPhRvTCG6OQgd4E8Rv6HAr6XzlC+RS0hG0buU
mJ2zqV4So0geIeN/kHPHqLy72Rr4wnN3Htom5w2Tkz22Zk/8wWsOSNQP5dzC
tf4ZQNrD2WHUXzSoRX6TubwtGFaHbb8VjeMv8ce8grjP6zzyO2410m77U1mp
ISzn4Vm0M9NIW20O88r5NWAjywFeg6CypD8Q+mapUZpoEy7gZYFOIp4+5bSC
9w0x1ijixMVwqyMFihQUI7VxD/IQSsGG4AuP4tbiu6HjqhHbd64NTwlgqMCC
nF1eR05MncjiyqyrVgM2WigfV3q1CNtyn7Nkt7UmpDNlBJru4O/HW+11V280
1nHca5g1Y/ZAOztjxP0Y+UvXZvTUtRIMnp0n+/OuWH0biwVtPmZ+xB/Bo7B4
81GPFyD7IWnwuRTj09hAvM1eBbFv0rSQxDrcDvp9iBjDxpkm9wDxgk05bt5U
WQdy+NIoO4//06yToHDCR00Y2nlAVuuXmIt9Q3cGDRuQmLpeWa4dMTGF4i6u
wRGnNbbhW+oVHyn8azlWu1IehFqXA4DKhB0PVodMYjF0834opl8c276Ringu
RAySDEa22nOVysNaffyk5h60AhW0f45W0kNFsweK+GMZfL7AUfjqRlwKjRB9
b/R4Gde9u0BznTk+Cap3RQrT/bo1i0KC/RZis5G9wZOYWG5LhcupHG4IWq1K
fpFcvJr9LBLD8QzUSI2BBZIARSmDasxQv8cRFaEkEuBfjmr0aaoKHzda1Cb9
MJGw2TknvHrxjEbBT6+B8oXc1U8Ts+DQmyq0K/R/8872uY+oRbY3dUfZ2kPM
vWe4ERnz0op2MxqITtHQew26Cx+jTGwIEJTOh+OVpTaiT6aJdIwbtzop20f1
WbTJpvRrmg8oJtVhBY5Oef6reUSTacaY/cgD9K/G4A7w8ETHVWRapyQUrsrs
cPHN2fC/eLW0cmK54LC6lBtW/gdyezDvoouiRIA3vbBEbAHGQ0YXVCf1M+D3
bKSnjhjzQu+5fAZz5WFlQJXrAjj8VJfk9MW12W/NW7wxDp9t0PjOY+9J8af6
dQnK6ZmGa5TV/OacvWBKCw9rCDsetQnt4Tq7oL/yqOQtwCjJ9yydYlvGfR/O
CdB5snCdqqF7wi6Ft6i41iatgsJFltAEW5HWZJ3dm9wNDf87aogTs9VToz9w
hms6mD7Ci9heH6dj0wP/TSPe7gq856B/KmHe6ZifaSi9PMtHypHUetLGuGnO
NCnfwbtz1VongMuE2BekNlqzLEsAr+OTzVMmyypui3UUxZP/esbz3tN87ZZ5
8LLaVQhFB5UJbGohQEerXIzd3aq4ANCWXZc+m6jF/7ITgDjRTwT9w1okw3TB
HzXbQjef/GmFvtbh9bTB5Nrz5A6w62UY7n7JKYVOZMXhTjUnMZhY4/igjRGQ
g2DDgGNWts250FVrZbX0jOd3V6h/pYD+rdg3HpRx1TT3Ci78WBa/xy1op+Xs
IqP2UEYTAsEwLf20xHz6eLegWKQUWW9zusQAdqURRpJuh8o6JEE+nqjIeSH8
XM1m+kCaYXESN6DKkf3U0ZcdjjivBFASFnxYSrh8fw17WPkqhxbtLJJgXuTZ
9Zvrb/8r9EiSqx+46MxmpKbRYkDNLMwK5a2R0x34vSAecc1bB7f0nNfiDYC/
ceYllPJw9MS6J7JL8JYPSOAmhvVQuHfWBFyoEesmhVz9/9UrAEo5q2pnRXcv
VUwXdU1ArjGijYUzGCojAN/wKibY/d5m8NxbU0NdL6wL1RNlgfiyr9QLOaJK
Ok1Urnn0dePgX+Af3vF15jUD27WqvRDqdf+K9/Ns4khmFyW6wXEfyC9LNvAn
tlngBamVa3mzTSz4/9rQhgW0RJuLvoYgVDMbLxRwJXVNBmMzDfnu6Y6Qbx0F
+NPKVnXLvgAstIncjeiQVaNFEBPz7vPMAClYa80pKwaY423JVnY/IVuUBg5l
/gkx9oEVC4wtux2BzDw0UoRi5aKaX5+p1BRaX0bsSaFJeUrq8lfzpkbQgbYU
6EWpz8SPu+/9qH5JQnpliyLxYVqC0AjPgYo+JzbN8kP0RouterfgcvxEb9IX
M75zQepFwIBfiURpUJJbhGHfzZEspacwBwtOglK1f9ZiVv4b7G6cUVvFEkV7
OXiTjYU9DqErZTyFq9x6XyFPSNWaz08GwB3oZzLNL+Xt0kq3BBUMn4Tp4c+Y
SXzIZ3fkhCuz38dOI7Bv4KaKGKwU9C2vse7iU4QODdEUMcKm7pKjoO6CeIY7
uaMxsmVZprGSgaz5acnB02XBwwHrr/9C4qmy2m0NvWBB+XEsimEcj8SXbsU2
jnDeMa0ezIuM+hipURSoO0e+lluuQiyt7iJwqGJOzwk7EMobW9IgYNVswxBm
lIhWt9b/Z4adGb1ZVLf+y03/eiSNaKy6wfJluD8DPeHonyaeuNqz3IWqorKj
r6sUXZov3wIbRu44LwUEUOrnXjF87NO5y5PG/UghNwt0ZgUK7TjXkgjWzMGm
C9xEG1YiLD2yFkF52Z7J0HKXXe4SenmL/27MGCMNQiWbNRuPjv2rh7VOvmk+
pWk6ICGiaid53NHWuR00JA+a7pZagEd/X3Qrf11uDOW+CYP5KOkHh2+H9rMA
t8AzASq3fygW5hLRNeBthQk0pCC2wBKEp9NIuqaJMXOosvbgmmspQdZfygc4
QqGIRR8MudXXzGdNYZIFzxq8stAvhyo1MfNT8V6zbQ/eNOX7wzs6KKum4tms
CVSrOZQ/+thox/gsvw411reAoupsH+1Npv0ZFyrgX3UYTDr5x9QpcHcb+lm0
3E47udxeHrLAlJ+Hyv59ZbW6Tj7eOMOyx38PdVEMA5uX6VeWoq7MGsgLN74V
aquHaucb1tnMHnGE8/XlYpELO/xuObZoVMmb++LE0t339YcbAKJJ0ERF9ZTE
VX8vKfgXK+18ukYUnyK7Djmq7g/0e35dDxO4MHIIt1Pa1JB7MgxeEK2nORop
v6QkzwFCc6mXEsT3Jxq31u/8/IzeGzOzatfo9sMxoih2Rav7S6Iv34ypVBDR
+cEL8fdcaFXlIfTXeTAow5y/d7TNeBJT4VtCNLjHAHvT66CSne3susdx1kx5
ZFH19rhEibvovOVK92zce9i0NtuKs1gFFPirAcWUlqkAkMbHR3cJYw9eQw8Q
6gOxR2zGwiSVSXgqBN5KStksPlLaLZN843nd15cSX2+jzbrUQF44aLyo6aXv
I5mRqMgI4LR0Xo8zWKXUOdNTI7GjB80WLbbHf8dRlLCEvQO3OM8IjfG3OsQj
dofG2mbKUr4KDTUvPSSX/crULAEcDAkzYa61W3R04n7fxBOiJ74qFUpOOGyk
D5/NVXr6czcwZvabUeB5X8Cp7xpGjvXnxve44mIw9V5XNiECzYYJ0b35n75Q
Fki43qC31QOAmC/5e15TYTrI1mJ8OpYYpGnhIZKaGRy/WECM5WXJD0Z+GH+X
CTHOGO0qzVWAaaWI5JmRRMIH0yIehFtYA/EwfzmX8hesTpBWRvzBEvinahcA
EmwOjd4yuYfmIGJWiECBK1lNlnb55VWKL0n1kwLsvV/AEPJ06zzt5XwDtqTy
yr0m9OPybyKraeBlitJeficSjf6CDqBzLclTxgowmgkAbhCO0/coValVk7YX
WlaASplvCE4dSYTgIvVCna/bB+mfOf4GpcV7eSfPHYgiGk0nz2ml+ib7bzAS
cyx0TZjUa7jBMu/r61L8rtf7FnQlKyWF9lW8LjSn+1THF2YZE70jxz4vlay/
xTXbiLUMTzxeUTKEFGu65d8T3SQhJQ5CXr5FYLv7d1gKU/LOT/zN7MCVdagT
Is3yrUMfjXvFI+QYCB5sKvFI8kL4zuNMMYVIFP75SQMNnkovtiHmTZpzzhcI
4f0Nos6OYic0+dzGWQT9k4mhhQdKy0K5PX0zOo8REjmw0wplGJlJDrbm4HFK
RxGR5OxOGo6JnN/PQ8frBIjb4IowQEfbudQSZOH8jJxHxd27AaQYq+VlHVv3
cAXFE93p4FALBjMESXrxlSvxD+E4/eU6SgaPTLRq/itX7CiwE+LpP9TjG2TJ
TUsJMKPBSZELjGo21FP2vDYapG1AyGUgT9YrjDVqgjtEJFP3as7c4oMg0+b/
aSGFoyoDGr7du6BtILkG4f+uw0llj1lMesex2WaoqQ/R/MAUd6U6LcGPRRIx
yvYxoW3GzqZXVmRDj5A0cXzo+j87W5tVJGrjn0oBc7UEwuBtTxCIh6WXRA5J
fG3ByUMz63AfdN9i1GC6wVh1k5m0hlC7dOAFhjpemq+0olZIf+j+zVNNyyRw
SidyesmCjlOwMHb9aUn5gGiw06z204J/CAinzYOfWCQBQ6ktUMYaEdkaBU4u
Qa6nU3E/MG3NNlgldRhYDssCEmlz0xLnJ/fL/OWGsbHLm6tlub6j6J7Kf+hu
2LPJz8CBljImIlpfZX84hFqXRKmYBDH1p8fOgK/4kVNDjTFFrE9onNpAcfbR
MzN9lfE4q+sRZGUU5rLmZ9LsY7Z6Qj9AISPGigDwX155VSfjke9JUCDTZZY6
dsBbw5GgRdzxScou6VcaaBatKItqB+iNoSwNbzwXAQPxiX6Y3DljtVVUborA
CqgGxI3Q9QEG3SwebgVs5nm9aEmtf6f9KnbExf37/vzU3e1LKFrNVNxpg+js
MAktelL9B0EevsI1FKer44XIEE9v7UpIzkfC6L3veB2ETekZDgaROmGl3SOb
BEF1HXuUtjYMignrQrTcLcHc5ii/hvBR9MXZvQcU7gq0Jddctxa79B2Raqke
fBzh2mM+ZlTpL3q8/cFBg7iK3ZICpBQcTsEVn2/m1sImdKShGIsSDIiwO4B4
jkinfYHNxB1vK8N2WRDsgkaoPf9KUWh+AxynzZSjb8b0QPOJpw6b7ozeib+U
ZvEEALWlbbdzRNJllJpwmVh6xpb6dwgln4jQ/0sYmJPvoJn7+uHAas/wLeKS
DSfzFMR1j2fls6RoG/2LjqqHH18Mp/dF//wpmUGu+YYqzpWrBNR/0Nnq364B
LfISxc3KtN28ELep1r52qOwD23dwpcSjpKwMatyxqma4yyIIuobE3D+WvU+w
4D9Z9l1ecisoQj9tWrH82GUnWIO9Q3KHxhzAbBMI9zoBYERfS6a0tqMkezDk
MZGjFOCsksAbKJqMtNf6F2bW9AJxXDzp9wMmfx9IDonKMX4sLaApPk2FyO30
DAdbms7yxBU4kUaasXZhtPNwmRX7S91ZPqNAp1nYNWKU2BXpA124Mxq5Y8r1
CMifwN+KhjUZTp8zVScvWbmrN9MECGW7TjCiHhGcegiw7IrF33VABHLvy26C
HMdJTMOGmwaI+2PnUj/y2//BKBuo4Ah45RuKChEu2pdY0cBDYkGRUtLtQMxP
k25U3d0Sga1LR/I6i8gukqep2ASceW3nQTY3MSlJ5/dgDDz7dSpGHI4yx8hS
gfZ+2RmdtV6n7heMcXP8D9tKhfF1xG20YY36feGvWJvpIE7JTvgqF3PqcprX
zwCY6eJn5JTJ3H9p7h99upjAvcw8eg0kCVPRuDhHqdaGjwr2ghqoamBNUO7k
NhYlQjzjYlbIlUFUhq01Jp9P+pXLHzmSyZaqKTS/UC3mGVXGN7pmcglru4sK
E8BURYLxTlwNfZtfEC2MrfQXp5mgstzlY/DyR9Gs7WVpv8WteeWzHzoGQOiD
RauoOzrMPvS2jdG1lssp07fYIi989L0UpJIG6fQbmmtnuS2iMruiA0EQvpFq
JfdyVcdtiLwW790OSwUte3TvEuBztyrfq+rFcoiiMw6MsWzli2pqOdQZv0Ze
UA4QcW+HcJDkGoMuv2WMBxQZ34embizVz0Vrh8wNCyVolr+9CBWhemCJYKIH
hS+Ow4R7kwYzjB6VViMQ//c6z85/FHbKZ1JH+DZfaOesErbONEThp/GSKE8l
l1FeIGkjRZ3jbv29s0eZMT+ZTXVdyNVX0WBVCGKWZqtMIJHmn1cITLoOtLLr
2MJisCsgmddfewXYTC7w3M3wzLiVTvsNFcpaZwiMNbR9RGc4mOngqqRZaMIt
ts8x7v2l/AYNQGqh+FH4oqa3e+4JS5HAciWqD2F0M88Qc6zES2H/AJ1hJ3wT
uS4kRYR+aNBVp/hB05Oj5RDi177JBl3M0uG+9tfeEWzhArk6Uh8MifwfDpSa
wCbjdlJlxJ24W6kIkztjrfZW8NNFv9AdK6kBMT9qBMrnNjjCiKlmMdpKABZv
M5BNhfb3MVH0QfGz9JJqNR+nPs4duAz/hTiLRJDGsK7fMhrcNTDGo9CnJ2ib
jBNaB/BEqb6T2fNJK4ue9icZidjvEekNsYdI6qz0TzuejxqtvwHIw6nNfZ2Y
+wHtDzsHB3koKEXuQlyVtUIim9/WAJc6SRdtTHtFWvM+86+ZHCUM7YERTbLE
F8lfMlM6UqgtiLpEXhCmBIrZXuanF5cXq2JDnZVJC8bgCMcpQgzytiTCzlE3
L2gehqNXDuYYmgx9Jt4T2/dEk3vo2wHUR5Bw3XRJmpMk8biGf00Ic9f/gXQy
aWamx2LNZTji0oqfIkPfKI+KkoYf6stZsMvTk9o3t3Vj3tHK6eZYSnYWquw2
/3A7Ge48xwwQMViG7zea5NnfYEOxrXWdxrnQP1xa4OP2yh34SrT4mBrOIvGJ
oKQYPAMjNJUPd+jSDkLRlgZWyjdxdnIBq6w+PCM7ZSIcd019M6F0RckwRVoc
xI1Qs2/OxpUBWkqKBHK8SxqJG/9Yn2R+YqA2JizdEOyF5/ZgSyLXJb/zMkV8
D48jGheqUvWlFQ/xFSxEld58rin4Gw2XMgIenBCrQkElArhsWHcvTJTexdVs
Mzfcyu9ZYzvSqgQark6Cy52kxSAm5BhtHECCP7OprE8RAk1fyYdNjysoz6yL
L3YWJGxoqPYgpZodu7VNSUACJ1anzu/vhz+X+7ueU/djU7duoyoCG/qmWU/3
TMljLfku0LxuXM2SiEP8xaH7gaoH2qrcBhGwPCHj/oMZhkon6qnf80VJ4/m6
Gcou/6wTQS62AHgxXZrVKKAekpVjecq0plqFAnMr6n3r6wgEFoESh0XYaL4f
4rWAZBh/DFv2qD/pRhyR8QWK4NoksvgaeMA/x5WY7YQoKAofCLdCNtSLs+o4
KsNF0+XbqFzPjmE+kL8iDR7dFWvtrqoiRNS0xxox+ITkWOAp0huOra4xS/GA
Lnw4wZFQ2/Wbja1VWp/F3wwnQma2zLQlIHbj9VXMUutls6Jc9qdElXpM/RJp
CYH2Ld8eS3XkuGQB410EQSISgK2cdgET5UOl4FXhhXkYBmV/ucY4Fhbaob6p
Jt2nNpLJSAsYLEVC86hgoOsl7yujYTFfWnl0G51xBrXMeoejC8y4Scpd/4zi
TSv6qRQkjnbRKgk1UbvDkkBfEKjkMpUFO5Gy14/C9bCDb2jcb18bx839wOs3
HGdUoHqe8j8a4TVU0qaIsrNFM46wWcaHcPbheuWeK48k78mWaNv/4wnlNVM0
EjjnrTnJlSFej/e48cTExkb/zmlf532O/XWu3CcbebOlY41M72Xn6OwV91Ft
1rrMjo2rWODJavN5+XWyvgUP/d022tzdR+xdY0FuxUpLkR/EJaq+51H+Fbz+
7WZgnwrMr7kAcuIjJqwar8uKrH0UZntHkIrPo5Eg8Imrz0EOemv06IKDcJ+5
TcxeQgUg+1kuA+f3dAQGjmO1IhZKWrLJFRX0bokPmniguh5sRGkc3hOgOnux
65uLPLQ650P/hTVrEuHq8CvXPt1eVYgi/raMhrQ1Lvl3wScLGTFXSqswnwqA
snmsHF/5PvRjkhen5JyKYUa3ltdfBG49wtV8JA9xCj+cJKpYXXF1yx77ez27
aSpWNzUt6YN7sNuq1ywlbtqM2lNliUQcWmqM+ysL13EupbvTwIxEeR3Z4w7h
jT7S8NErfgSWrLkchCQS9ie7rn75j2+i29pa3K+2ziNAF0jWISuA3fJVEg2x
O6+x8lB9AfVrck3m7qzvdsZ5164vnqH8Aarx9tbUVamMRKfwq97XvX1aDb3O
RmAFkYDNS25KWyRc9q5sF2eoadDz1WYvD/2ahGWgyaYZZr5TlnaziBkVHSgU
BwKUyRgRwYYv8zzF4j/4Yh9QMYlbrnTCrNGINgh03H73r5GUk6VS4xwnn2Yn
1nf3XtRv+o7f3s2Mb1BktJV8DNoWQckQlpIt1knRkiWhpLRp0dNgxt0JqQR7
k7FeN2wRwThelWquLF6mOEG5X2oZLSStSNiXGBdECqpi5Ja1jTjykgPr8Q8f
Xwkyeyou7rQJuici1DA4LpLioITnOLeRXneLWIudtaO0cd+V0ksfu5o/ccRH
uMBU9rx2DfuS5wRPT9QXziualAlv5zliDPpsv8eyIwk4TyfWJva+tI8lmbfI
uFltxvgwSLT660RYsWAZwPQgsHBVgEmrFkNt1+LXWIUfqMI5PX1SPkf/8Lci
TKlcMacdHX2akfhEB9eST/LKltlD5Dn1Oc6JZZP/328RAUfVTUrL1/rTvuqX
BnBvMdHAnsQkj9bZO8anIVz7xpjRLEA/mM1jes9+SMwbtDdOuCXiHOYLUHAu
p9W1hCrnEx07VL5w8nkOUv9qp7kvwKvaCgA8pHo7Gp6pk7WUx9TD1G1GbkM+
gXnkrwucUxQQUU8tjjMp9+xqDWxFSZjQyJv7UQesTv35k1fWz/9uJ5K1mrlq
trmtVXeFbCEgORSLtJVzXpIIlJoRHFnzUpSpxe7cb2tj5ocU5EFLoBXTbldk
P4gR24JSMKP5Wj1nRzJQDSD/rdyXGmXSGtEH/ibRk95EUN6tVX0hger1igT+
EwU+dAwe3PJYnQrUxyzUTtJoiqcapkkwHL84wi74F9d/7OZjywB2j7dzL7Tl
FnOt8vyKC2K8+CbchzDpAoAUZkIYlS3+YKL1HpUD4860TtvhP2iksmcn4hjk
rYOfPylA2JFSJ8x61byIBuyW2rjiNA0Vo3Yt/Eupj6B4QhWzAX8nfAYsbdWH
cmUNdinhBgEZsDy6Nn1RprFo+5S1cRhyahXDcLPEFYEFJLqJ3EFruHIJzHBI
Yrtxtk8qBnI+Enab2nzxQQe6IokRJXAUyCcLM0H00cOFnGVQN5sPnQjO5bEy
ztk/nvx+rRapvHNzBe8bTguF4cXKa8Li1ofQnRzwDf4fPhgd+0kYJzdhF74v
wsLTpyylS91Gehb2JqHxlMpjidntLEzDfCg74JRqqrorxYpyVonvPZK+k3lv
h2NwBntCLRhNg9ycPFbgwrgGEVflvVF+9Y/aHufUOuhuLoa37NAxduXnVqUc
2o8df3j3sULiek0UOJsHATs5vGjxdusr4qIJPeoMZdsbD5cDpow6Rq05cC9o
sz7ilC7ITvvCfwHirSW6DAZxr1BoUUzKQT9mNEtuTP1k/h9ksdzeKCThAgtc
m5IQWj3aeOej1vyogpwZeT2Bu1OKRMrcb24FNhPApCfsDPTePWOwjPh+qbP1
8r0rq4RF9imFj9z6olbgx+XjA0TpowC0Gmgdmt1lz6FJ1rjSDuXu8y8fWK0S
yQAme+s67yBgny5pQyiNCBbKulpt7b2y3hgI3wcPegt5gzVoEHfmDLT5ZBZB
heCnE9OYaf7d9yglJ+XRt8ZM8JekOYiqlS0J/btxLhEqKiBRdG+6YkWpRSbQ
XsfjjL7FL2y1PVZtZrVTSDpng1PdihUZ8T4JYo1nNSlqoGx5HtxfbHlVD+oF
MJ8/y86GI+rPzHaSY2/u9shr1sDE7hyVTBpuvYNDN+AEXwe1dfH5VImffOOl
MOpSaiDi4cycHEc6/wd73nzyHv/xQq9y852xOXTL5WeEQE5xALz+p17F1aKh
ue/BGKh5xD+kIfl5f8uyPfNXAMp/pWVA0dgl+xtT1o7CYTpZzD9xQqiOelcr
cHykES7inbgQ5yqLoQJgdxzeDlCFOaDq293AY+pH1S27JoBwU0fGDIAdhJRf
xpY28uhDLr2RDlkz5saJorb6KPULtJaUasU1b7TNz0yl9n69I15r++xvUlMI
iEZABAEWJ3fFqGerVjUcrrS6+YwUmjlYtfk4mDW5zwhKF0YSqPFjwi7p2pAF
IZDuIik0GU3W9Ch0qcME662apCCsQhcvIjLsi8z+PsRdCQeOKjLRS4fiSkJa
zdSJlAjAtZ2S4lZQEXm0OUhRO2knWRO+aSGyeMTO+46s7Zb+/iS7HqNMRY86
0w+YoGl1OKlTtbhu0NxoZsgpTJz19EdmRcVs2wW4q08NVU1KEW0qMkBUjntm
mWI9RZGUloLfx8cxJlwGcUPSrAcjcApDlmpchWL2Fh6kA5DtkrJfmxg6ucxl
Y5HbS+esVOXMMIUcyFUeAk67sEGd3k/h2kCIz0OsB1i1cDkiD1Q6mSE3cKmS
V5JpHpyPuXBeirYGBCKW2IlddRuMasDgswgKbz/5bO2Oz5Y0gZIwioJGmdpa
w1mWAbzvmF6E4lUr6GurIbgNGWNptwwcUolGnPQrucLaed3XIKwJSYxht+gF
Z+GbdfnEMSOYjB5rr03A8UTb/kuxYj4SRxwdRpTlTDRv3FcAI5KayHdnSVdj
B/ImBk14zWlMFAMmO9Lpmvfo4Nw4O9o+4Aie/Ot3gxEqrx8dSpLo2rhEgHU8
DymSAGMEhaVgVmmPqhEl1Uhv2jbwz6QxcRMFo4XQai8yenzQchcm4kHklwcy
gvvjshXnkrNA/VLlZtEo2712vgubZSdB/ger6A1uicKylmdWuHkGwhKz8y9L
eZq3HtzgENAYVewobST4KR7WDyyY3Xrr1hksb+pWIxjpUDMSeteqJxbr+qzy
Vag3UEcPNAvNePKFBOZGp97fdv6krcxtr+oXVALPbyQ3z7/iq27ZxjYTaJOY
vvHR3LJDV3FXPxjIRBi2pwsE5fQAPZgRO8PuEzweoB60XDvkGW8KoJIc9rwh
w78z4uy60OXuXJV/82NRm96/uCYiNk9iZ9WKoRzHiSzcfzXGwTT079G3ZCWB
uV0776Bi7957Q99KXpK8XF3qTnOz7gcaQcFt3f4kYM9ydlEuRXV6NUFWrs4A
U0QtY4fy3HSRSwzpq/t1DOeeR8OXEjdqF3FP/i9tr5s4+hGJ+/ECVLfI91Xq
jB3cw4f9XUvB2PDxsZr3tEYEHGzQVfCk8FY1jsinIcdl3rBSG24xHpw9dy4S
BcQwGEoCfWpF7OShtCTHwk/HNSCfpWt2ptP7hh0MsMj0yXoczyusyZdfMaNG
GU5jRMEx9qSDNpy3hCfii7UEzRXMrHQOQDce20KpmV/EHhSA94SRdizukaPY
4ZwzXm3ncYNF5JSwyRc3mY0U7TGJXm3ko7jX8sHjM4CbVcZ/rLbYKatWPAJW
VPXXBUGGLsvCubOujwnyLNxFqyC+/iDIte0fWiIbSzOdma6eNpTQK/WM+qcy
ncd1aexTs/xr6cIOrTNI8jug4Epqp6MdQ7Cb+W9g/HCrs2JSY06gVQ1CbFfc
Jigcz1yNo/yW2XK5hEiNipd9Fs2xUAxA+TLcMUzPDcfsyvX04pB58/ls7M1w
3M7GTITJWc+PxkIlzlK/+yWB9i0hYwRUx1jiuT4QMKOrpDpDweZflFdyv05X
EKoEYyaM16j2eU/reBpEFS4kxANojiRHTlcHOx6FLwrB/DanGrBNtKLIBMSx
c9hCD/kDDZ9bZJNPhcTpbhMUqJH/lSCqfl5Eb04jBZbys8IJg6gWGgK38eW8
Xcej9W8b8CXMiLObT/jCdsL8lcbfUPPh7qMRvnDsVet/FUMr2JwMCMWDT4Dd
5rKJBA+0lGFML6lbubd95z5BCNpk1F0h8fdWZeo9Ynb8iyxf0VYaHgAFeL0Z
250GW3FGHmkuONS7Vb9W0/rPw8bJcFATwVmDn/1pELYRyyn8TE92GS7aie5T
hRrm22MpPax1Dt0TWpqLwOrnRa3nxEdgS1kKW3ZArsCrAwrM693Aqrqk2ss8
j7jT+yhthfSSJ3ZoP7eVtbRER74K90QV8t7sV92rB/7KoTeP7Gl7h4jrLz02
4aSWyGPw6ri8Mxl+RdnbquIkpAc8ZRTs7EigG38w424oQDDcpj3zyakpX7VB
5FXFQ2zWAoMfXNPofqX7rBgfRPCWWYXXJbSv7Jn+BRJvToNvssdwA/X19r40
t/whrqV+bLpnP5zie4pI3v304zPkUHYsEDkksrfPATI3q1oRbSbKJQxnpRED
XgX5i/sR0mDEDLdiohJMui+yXC32BSo8qXsDugY3YE7g5/zgMXR23z+qyzBU
H1l4tfxYxcJ4WT3y073oJn2FShdG6Gj/hAS5Bc3tys+Vw9lnrADS+cuJ8rqp
jnkGhXHbRQofysSa7Gek3g1NgtC5lb6aKV7YHgHbsCMwLn1cQ9no7PRsdpTZ
QhjOhoGC6GBrJcb/CHJZBpFt6lcoQeZVnDwUIDuw/x1LnKMYtME8o2uKVMJl
66tqY6apZ4wv9G3C7gCrjADPPppJEp2/YOmb8+EVkdDyei5/DexcNh3T9o5u
iikz38NmGZPUjXJjiK4lRzFXqaQkIOV0Ew8UCkP05IOCsEEDPpjBKLqvijnC
hLo1Iu4YTzkoXUy+Nu6EkbubNdZdZFSTtj0YY57BattCEr9KarLJWQCtUPSY
Cn8RE/5wtQHZH/lher0v1LdHlsyzMs7lMfHyV8pKqIdIv7EW2cLsyCJCTSQf
9EMtTp19EAea+BJpwzW5yXPM6ZOVBKWZ5x11GQzFjknKF67bnpZfcUkjnKAW
BloVoZjDm9xMJqU98yii4sfg6pD5n0gszCArJ5Y1NHSoKRZ1O0zjmyzFQmr1
W/KR0+D2d490clehkcxeTtskfSBzMzoC9KSfB4PsEnI6iKSHmh0kxq805jqj
gbFGw3636RyOtT9N/meSOEYcmwqmRApQytWUVnv5rCMnul8DEQiGxgmcquV8
e5ysGhzfl1FZcv5ep6GTOO36BVo0huAFSssQPbkSssVJx7Rtg658xWeqIpBZ
ha9A3/NtJBffztE18/9Zolu7entKnFUStqCeD2LFC1AWV0CdfFKPAp7C7IGd
ZntVytdwzV3U3qnRRCRiOXXLOclog3wnlmNdcYfW/wA1j9l5+Kg1ymEhJFjC
Hl/2k+2HLHOUvT7uZn2988I4ul1JcsPQvA03CsVyEKnUtPsohLuIdGVtPIOM
TXuDjUfBO/+jpW/hfa/LeknxyVlsNn8OyHgPWb0T3Mf8nn6ZqChTo7KAJ9dL
q/Vp8avGWqh/x4oDK5tLCInYB/FUIMtRBRvc4sAvlNIOjafhd1F4IB6zrCyg
/hkBKiP+OUVzIAWpE5iD0Rfp18uX1vrxDzi1fYiNGiTsvBshLBASsrWwE4vB
SCawckCR89Whs3tOmybd+LWMZe3IHqWrJTG5U/iLc0HR6RjaLu7ab/Oj90tw
4kx5/nCJ5F/4rxBUJmeWObvrQ1PRwPcfSJBbZ6PfwP8cq6031Wrhp65etjHN
4KHzQOC5Y7k2h07RwnZYi3IZtNzWjzPGelwOMJasZ/Os05sipuoVyu5M4o4h
0VAA9AGyuJ1F10TKKJbOXqmTacqZuCa/YNdxhs86lbCcIri3jT1XpsG5dbVr
JZUWlYiTIjZZQeWD+btfgUDYt84x98c/HXqHuI9YheOiHv6zPOrOe+ezv6Wf
aJVwo1Ae25hjd0ecKF8Y+97LTJGPyaNpC0PIPe+bQJQg0iNwpqGqkxdwyySl
4VmFZss9TASq9PtpQasQFaD9wI2SZfqzR4zZQEl7Aesr/erVVamFN6DNk9MC
RjEv/mo9nOxTvgmCwSgV0MJjZisi3Yp1mwUdkkzvLJT0gh3soXYS+Bm0ee/E
76JwP9OT/eBIoasHk47s5kyEVA4wVnD8RjT5aG/uYow/udXDAWFbAlqSP9nb
OPPjqFcdeINhDPn+EFyh6G7WUmTcIY6sVN6fIlvTs/OB7sK2wWGNYma5xPId
fwC9YbK9mIPx6JwKNYaqkB0+Mhkzf6Bp8HCofqDl6J+QDh/KwGGyd9uSz/Pk
T14nr+e9MT3anFUsDNPPdIHjDIerXPqptUm4nI22dKLOqulpD1Ng48HSAUyA
cS/XHuH/yZX+CGd+K4RIU5wF4t2A4TlKSjLRZMj+OL0Bya6j1eZ5FpFo8fob
gZOc+qVjdi07RSmFpXDD0m4d8lQ1CM15Bjns6X2VVrXTC/mNQqflp9e/GTVH
4mOO2dvPvYENcdCifng+GHAEgppVL5y6Y3CZhCyiwj0HOVKIO6rLIfSyQdkw
kIr+T1dOJHBZhgfbcR9O603PqcZLkSJaPZy1KWdbheC+WVlMHgsF8a4AOG74
sYJ4q1sByfITNsyLhvygF21CsmMy+CXWocNZXS6BC7OQ3BB67N59X+3OGKdv
oXgp9Lbq/Nh4ZhBtxu7f2AvN9+dsz1qaKBJFsCbEdz72t5lM7JOo65Pib7Sx
jeqZ/w4PbiFjxeUWwBwjxhx8AO+ycbq7VHWwfhRtQ/LwfR86+ki6o3O4WPIZ
TQrisaVVXGUItHYjzv6QZJUlt1tSGCZfzqPOUC0rUDbc47qkXURFqdCISdhX
BYk07uq7tsTYvq29825IjHUaI5i1PTjQHkl2Nmyw7y+dyXHt95Avww+ETtVP
i1DDTRES4+2KdmK0eM/D4dMMMW4Ijtvh0B//EHgS46n8qZo8M6BI5mVnp4k/
sOcW42HSNZQWiSSFD16VEy5mKxXbvkPni51AB4FeIx/OIg7EeLc2w07wJt1q
m5tBk8IW0aXAGH7Bvwu8Z4qfJbcJtllBFG1RcwEJwA54C/UmKOWPN3MQhhZu
i/AxSQEsMZGHLe5TXI05SnxyPwgOEUDy1t+L9nDBjlGFYgSVlkm7+A+N+KLE
3t79N+TXEIqteCuWauQ5sYT374cGjE5gfM/UthOSnBTLClWgVdZsJyep7Mpw
pYsMHgwPWp3zxLSrbJPq7wIhqETmddz9o6C+XUUdY/RVw/pmt4zqD2MiUn4t
Qg/mjUsOfyj1G2ZtQ34AhAHFBMI0GUdgE0jcx3HP30mraW/6ciZCk76oSUrx
OwW8pqWTs23hGTkjtOHck94TO/dMYg4A6HY1TFVCwUwERXl5QgXOh2oEqHGG
6pefdYSd8RZCLSylLBR1gyN3uo3j8/h019PPEGQDxJX4rU0gb/u22aknEtpj
KAYhvf5S9hO6CMF4hQAIvVsswhQXMFqTAGfi3ZsQM00xvW0xOOyBTon5R8jX
AzZMfkHVNK9ilK5xxTaoBVOvavFEMF4wRZipZi8HQxGFuRLt3idffT8fzjQY
pM9gl98wXuS8imlA4ygjhg1yjdgdJcoKxKGFsfRDDanVt3LkpmhOHaOu0Ave
6dWUpyCm385Kp0Fk4dyw/hjAmUbdyRYZjmW9j6LTZVO9uWxQVCmrWiywpgkE
NSrxmE1u0VU3OdV4HOrxt5Wksfv8IGLy3Qp1TQhKX2bQVGHYXuPFSVWoOU5/
XYGyauFeFSrjtLjRIHlWpCA2YL7S80PuWqL5ckUE08uX+tzB+Q/K+nVQyVPO
xbAGhrARIsvITS4NIx0xkvMuLqIeMZbO5cqmfzN3tJykzU3zmGy00aIIdVyq
AUS8qk7Ob76DQ7iT4C1Hv+jx1VfIptdPZSc7VCQhCd26tKIuRFm2oO8RcG1f
uwO8DopeLgrW0Z+hTneFL1+4lfSpXlonbEr1c8/mAISegrmJlbMelNTecETE
zRVGzpW74jk2FicSzAgfFj/ICDPS/HMkjmrlB5JRAQ5/xS3AFPMnA3EFLlz0
GgKFE+DAmSbkDoVcj6e181w/ZySCVIK74GkD0x2NtXJs8BfJ7wIuHT36FePd
SFzqzl20LqZPSxA9ttifKknuvX808l7oltVRqqoyD4we9QtENn2kv0n0ewH+
GTNX788z9W5ZlFaaaBVlt/KKusyI+52Jqlt4/s5t1gFht5AvVEpw9L6po38B
7sbHhcSEi0tvuX5msXw4+ODHh6aZywAdsc+3ZsBnzBo5zU53KTza8nxxEuAv
7Fs9blQDgjz5asn/EZYoHhK+zsLwSe9Tq6yCQqa8weHialBCTq79c67++Cqp
C8s4DZvOpJ9479erl9SnFT1yWYpm0kWaSYvNV+Bt3t2ySxjOaB8a507zBKgn
HhiF38dJbsj5sk89HNDvqnmOX7C9L+pxc8aOit7pEx7Jff5agJH/kJ77nJYr
M6t5mQ/pM/gT2pAh3maO4SYtbsKb9w3xXxrtANCfQ1jWOZ8Woy8FFocLJ6qt
+CgMQNM6X3JOV4S7NNNENALnxFBeaHoNNUf+iiW824+G7qJIbSmpbMKPTdWX
rpYXIUYworpzAyxhwU/+rx4Gp7ILMKKrf/rS7fVHv0W4zfxnWvsCCOUfeicg
jDlFJrD6Ghn0VD399p3Y9G2DRcWk0aIn228DlnV/z7k5hIcpw/3DC8FCno+e
hONm004iT+t/dnygVRV+TZq8tGAaxFBeJWoBKeC+OR9uI9K0h9tkfMqmXSoR
L5vXvNrYSkb/V/iP/eNC9skbSau5anG+v6crf7U9jH5Qpqr7rqmNeE3tT5im
ktPI7oL9BfyZUNfbVjt7IgZiJ7BchNLOKYWk3o5Kn7MRuFHF0z8b8zWSZfzx
QeVjv2tTkac/QgsrQQglbDltNoZjWw5ZNnbpT0iLB+cgW1s2VkTRAbygfFTs
8/q7YyhQdQlPnF4dDzSoEWBDiFqdMNfivpZo2Vx/N9+DVsJRggt3c/qhPj2C
i2S+6tkCruTfeDZc4t+G+oHVUMCn1fuNuKHyci04Uw/wtN56eZFics/pDpXB
+SrFVsdxYyCVIgMC8y13i/SqExwZbJpXYCnEh3hTDt2KFNvSOP/A8Uf5DKTw
6NSV/Daz2DhBYYWeOCl4PpmDDTQqrl/rQjJNOB3w9Lc2zZhWf797iCY+6/3h
6793Kvru1Xe14nwYZB5OGb8M8w8LXmZdXA/YvwUdwAzRI6icheBFy+aTo35d
te6KXCy8y92at1or76+IHgOpgqi7ZluTpCuEx6GELB8/14TTUoBzslnCIot3
zLAoAr7/TcBDxqvhS/9a9D/4Wj7U7OwXcciFknQXC7NloHB0dOGOKK/+Y04J
N8yvJRDBrE1nPcFhIV9g3TY8L4i7GFHAnl8jPvhzf7eoP9iCniHnD/Wpt4sk
RX31sKK/8A783x9egELJIDcDx43qXr0rbF57ugJo1xYY8fskig9toRjrrf1X
yFyOMUBkqzozayu7L6nU9mvGfqbcUscUQxLO5MdaZmle6B1fG1sLctbFiIsa
J/AgyIlABZXhwwZ9DWpeYS7cfW0gGIBq/2ZWkuvtFajt/zgOr5z86PuTwmTe
Cr3hkGuw6MwpIGoSZCaEn9exVB9H2ogswclH5a9GxeVaF0MIRid4toQK9I8o
nAyYyQprd8a5O7y3MFdUAoQlYNgMCa9Osj6oAbJVkKIPzQ+h8qDXWE2u1pqx
pjVE6kL/aHYcfEIf1jO4GH80oCamj59DN69MPkTIJRxZA+sS3/HBSJ7GYGFP
kOL4VInLtHT5zPcmpv/YviIue9Gse8o4Q/pO+w7Ew5F+ptFTROvV2Iss1vHO
Zt68OQQ9ivjpdOCVJZCBedNVM4O+gE3uUZD+Gh6ByNUuDNWKli3L4SKQxN7n
g+HmmFby820cr2Hzff+cqrYD8pZlmvor9Ld2yxfRc//RXeur2EcZlAs3SNqN
9axqpob0ACkPc/JmmCOSi3Z23oHPho3YnByL8KXXwznfRM3J8qWy0StBZOwd
I0luyO54FviTLkUKkVhVMQv6lVeFKqV48LgLy51Df8DhSRk9DAf8nilvq4Xb
7J8m+mHSfGBk2Ls3E2iPvPZCkiJX2yQWKvIF1pIsxFCMvpkJlX59XBa6cFZQ
0OMxajaPlmUivOMNQ0DRzBa1v3Gs+6WYfdsm3Qs4pYFmfOYRRefjalzvcZ+A
mWIJW2swi2CmTqB4ak17cT3I1l/xDlTSiBFZ1NuDs9z5ObAAom1fWkS3h2fc
erLh91IVI1MGV8fovQyf2KX8APsfCCwbzRgG6tWEQk6bU1hfvmbZgxpWb1nk
HaTk7JblY/841GNWU8t+wd8GBNOdT6VpluFo4Bnj6e6V1yap0D0dNvH/jsfG
qY9zDVc7MO30aA9/0Pxktre5sfef0B4jb7iovThO/c4buBdGFJCwUUkJi7m/
aY4MlyLpqSLD3iQFbTyzigRW72lTylippYnPy2+xl4RinHV53RdnrB4UHogO
Z3O8oD5YG05aKsojreiKlZ2s/ITmlk/jRoU60iqyUf9le4B9ZHYCWlSP301H
w4nTsXBBrQy4kheT4nh5RzyFGoQu+S0wqUWcYqi53qNLzycu9gGhz0Vz3WHW
wq06IPgWf9MMBPLCsgGER1+L955h7MPe17TS72NW7Jh5PqbETJtmHLnBaa7A
aePOoKrMyyKz8loknzhZsKxH5mwrfxcZewujKzlZNlsCZrBs80Dx51DxsQgU
xi+NGd7OtLZYDG5V1/LP57Nnybd3fbTS8DqpvbzywGISMNH7Zd/8KcM3LY6C
FrpP4DpQBaKU2cJwAKdES1pdR1LMF7G8paJedh8dGf/Y9qx4ircIqcAKDdcE
QD9g0DfB9jwklYLUa3NLMJYMD3cavctYE33BKl5IXjs302p1pvX6/yFlBpAw
IvigIORdHwc0UdYBkdzrcEw+e1x4xU8769N/A7dBqpwrPuJWO6kS2EYr9bmY
FiWnH/z+bsRcwvSWIh8tQVnoz01fGLga6mSQQGMDtRc3X2APGU+Yl9/Jy6Oo
qlaNmSE3uYtdV91d7eWRIHigV2Qc86FJhCTgCJkTj2txX7gmuMDoLD/c/7Mq
x1hGIvUbe5mgSlPvMkQlXXtTeoEjlPZGNY/PPnsbq9ylU0jBr6zPi0HCPfOl
e3NGumU2QHGBiT6yAnnrBlri9ay7VCojDx4FIVjvSmEkZO/JksMTI8K8CApa
Yd7T0aNX5o7g7sX/qzdp4AHZGd2jN48I8WG9tiMC6FxxQS+OmuyfTEPThjxx
qpAVOSFfduX+M3N/lUhtpl9+mae8IeIiYxWUlGryhp7lPKD/vmFTZXHk/RG4
hgsYa1B/qdjBK9Evgw2VcX679G8rcClhIqYzKOQCeUJj7GxYZ7tHkYYm/cJq
lo8scOZ0b4Fd5cn+O9HEbpKJzTbnKiJONbERhX6JbgeO5Pgtxilc79GexBj1
L1V4HXRJ24oEzGrcFHOfRBlAuPAFrB4abApAbGxEqRzzKHqbk9z8dCUyyznS
kHNQHQ/r92nJC902UnJl5vGIi2vLgDMSzqv2vmc7d3rbg+PXEirNpCNDfWFC
KWy+FHW6Ky4CzHhqsEubWOwOeqTsrR8uAlPuR9NMCI3CmcKKHqxYn2ikPnut
MD6WDQX0gXObQojolrlCl6wKLB/rB54D9WUF1syD9J/eh1KQIxmHfiu4u/3S
dHW1Qh82kFW+zO62Caz/gjS4a0How8SMQfa7TFaR7UbuFZPtkGNZBfDto2NU
YoUmY1xLZM1M8tlbLOJYwZ6KV/bfw6YRuTr1Q/A8f10VCZBWeFRymkGskWv5
6dekuJ1omN9cpqVuN9l4fo8zPGJQxqqC/W4SbsI66nbf3IB89z/4Zrl7KC6+
3ZMeyrODjbUBxAbzKf0jBVnT41MGltC18fJDPzkL3yyG1OAxU5DBYbLGMB77
vKOxF33dKIPnPbHPqy8Nv7sGmwijX0KX4fsl5H6sWPmvwmt9NfVjwKwsZAxK
++Kj//dI6Dx2mez6k3Ft5KUT84G52ZLTmPEBVYHPZH+f6IK4P2iJXU4YWJmY
bsVkRHfqAX3v0ptIgcHeB6SFnJkXHD6YAVwzTp00bAA2XsO7ELRTQgI8PtR1
mbFppX0h0AKtfVNPnqD3BBW5wpSKgnMq6dm6sCo4LcDFX102QiMRPt5bd9VM
k2EZaRcjHXdYWMm2Brut0puFUAj7xhWlF6svNWUA8QrQsA8YV+6f8S9Eev3q
0TeQ3BiTnmyyprLmhOsgHcJacOkL+FfBnP/SXj75WoCaHXsvcqBlj7qgJy+i
lqxNz9VZUrFEt0HlwCnLLQ5TfDfmZW7PByf99H75MpV/PpzHHYhZMdGKBsdY
dD/Q7R8IKc88lRdt++J2lwijhdt2Uou+U1ojt4M7l2kUELdJbMlt0fq8D1eN
0clQaw91dZa6b5GLK1fgDV57UJfSsn+ok6Fs1Vra1oMh7FW6xrXymQic5TLR
V7kZ+t/SVLBjZFgwPOStDnb0TYPkxwb3Q9yo89yYVUHx/I9zfkGtzPIBDzKG
SLF+SKPudyYuie4Wtbq/M97Szpq7xwuJpkcIMkfL6IpGW9WVYBH/ZMfXwfqD
d5BuRxxuZQ2oedpoKPU26gbGvGS5W8QXSDvBM69FoO/TISYeuvxnE+g5Tlo2
oXbZO0we2Aqrr2rgYnN6qUuM/7ODppvHppTPAHg47QzHe+EaOzLD5/xU4LaK
qS8bnS6lVMArZeZLt3jXjAMb8Y8741DFFdk+WCImc/0ull8GsUnVLjiHgnc1
bnlV3VULrvuID4R9yba4r6SPJMw7OsunGGlY4GO4FUQGNq83/vFIp1a2/uKg
RubnAIeUErebLF8AvlE4fWyTLkSnfc3StAgbUh5IWq1Mneh2+YhIJW/qEuTv
SIe3oM9dHgDIh7G3vFsK1hVsEAnXeAxnggsY/Q3ajlr1rqbzgRMClAJFprvT
oluaZg+4uXbCQDHHVl4Xu5QS+QqDirfZA/rkaI6eYdy7PiuijANouXmu6Al3
8IbPDXHXkVei65dvxPSoSImGcTWNA+staaLiRTYzqBdnS3jqmc4LNT1ELtEf
XNe90NDdR9FaM2wIV1uNVHOT8r4sAqs40fGyheNV9v4NDIuu+0TblCbLWKXK
lg0MCcg+ynLha4BdMF4xr4+XDaSBnqrf6L2OQ90ihuLJHMWoflZtSig/GGps
E470Lxi2gqnyS77Q6VXi7MkO3P50hDBZ/r+W+82FDo+5I8ltnIF7L5ssFsNU
f9/dB9UXEDKaIGAqDyl8uNDRyyyKk046QtdN2NABmqq6MNH7z0Vs/LNFagmf
diqrwREZ8QZkVoz+Cd6fPONS1khPcInCsfZzge/BM0MxuzHnyRtRewzu/1qx
N1TQxsI5OPeI7+VRl3EV/C8wHDO1lBRVunejrIbtCb6nlmbcWOQGYwt6gGFZ
01x8c01Ean0rNtvhdXG0nUp4iklE3uBWjnZSp3GsroBWdTaDR3uM2BH9XgPt
ht2PJdtIBlb+zp8cr7zkEoy5qFbUxXe9442jZKjClvkn/z4QUX3b1+jNHIPu
kgr23i8qgmrLGNz992wylM4LOSdc5t3cJX7jj6P58y+eZ0+DNfd+tQD7I/ZT
I0dPzmW0yeVk2YHoQ7JRU9NwvB/B1ch+ecIuE0kSo56zumXNjZnVI+kw+rZn
4qLE+18/Rr0o6/1m8OjnXe1GCCFRr/di+i+C3iO77iiW7/seIcPFRflaMBpR
NISyBo847thPX1hNZfRccijC9P9Ixm8YGcyku8G/ESWxzx6In+CHmIBAY2rt
305z6MJTPNJjY/hHrAcYttZ5zYxHX8GV6SeWH0oL1jQN7Wsd5qLxg0ypx9tW
A03q2eVnWq92yT7V6YGfBkoAlS9XlyPhq41lfCk7rDwPdHKWp8WFkGhnUx4u
XbEG/WlHI5P5YLUgb9mOEzu8nmwi73kA++GaK1MTVFO39QJhZd11oss57oSA
jLtr9H49Gwl6Aw6wJcQxoq8Ui/Ckr7v15e1brD6szyKxJtv+kHCfAgek0/R6
Cghb4DkcCAqyCS08PJkgS+C87l0Id/cNVzmjxb1Ld+tKftkkBAndQRS4W4QF
kJOxGWO+98QNYfWfzuJ2aqD2p2VYkV+bbFfboHbYuaRkXkeoW9OeJtuW0vP3
h15cBIPiIMByXoEP4NukhaQSFmOqA7CdKJj1jxDXbUfXucKB8yGYT4B+BZsu
VwOp8ACY+ercekXL/qa2DlZJn8hatldlCHZWj3FaYK3YpHvX9C90UMyXIVN6
TQFlD9QIw10/yJlRuLpgMrHXBj6HgZxopb1DjixEvUhi/CD+Qn4jtHXIuERo
/VjIn6UsrgHgBIzsk0wiQ0hKKI13GOWLsbhNd2JitlmehIV6AVVan/kmBW1E
rDe5KQ3XBqOCuP6QQArFSd28JL/KjdWCSc2ruSo6uXjoEXzbi41ki9YAgtAC
Z/CQtKi/Fyq4RX1676zaDoW181ciLXf9YQghe3i6yEpdwKB2t3ypa4e/VT4o
mg9FYITLV8fqpa+rY9AZXh4hsERUWUvrM2NmZnRWjZI/oPVMMLgeKeIT+z1f
YvasFFcuCzk76GVeDZAAbX0j77js4gfAP948cLXFA5xnsfkIBplPD31LD6Ll
31eaabJ7qJpo3HQDlgjGxRsgfuNn5m63ekvBMFmnf1ruz+nwDm9F/5MpVEex
LXqR/F7eTB3eWTrL5+thtr2AeIMjySRnA+ofiAk7lEztdug5u72aApqeo5Ea
3a0ZuSn9Gu4bn07X1u0Etu7yMQk83347T41M59Cr6m+ak+tsHftM2XymUSgU
Q5v3g7q4Hj5oueq9B+O03u+ToGryqNmNgXy87p/AjdffPMT3mpyJENkdxP/s
GkDhk3kw+lEKvz2szVqcrjlT99ZHyCirshZfzbG0BBQPpAEmVNT9lvyZDRcf
tUm6VVemFltwmxO1YWI6Lof1NtpyTQUM5prXUNCtm8ZeB3D5ffMHG2eZfxve
5627BuLFi5Ug0Ok1i6Y0GPBGKw8v39pT2oOlpmFFkUIex4onpGe1fZc5sFoI
QvmaPZkrEw06BYlX7Dr456X6Ab4rxH6lZ7hSn0iJ8F/c2owOMpCt5bYDIH3y
lT42RzV4ajOav6IAN9YgZIk7yxJE87grtS9RETpDxaovmrLJkm1/cQKejo6b
91u+ZOxK51vwxRIED0wxf18VITZ6DC3HyqEcq11h5qaxT6ozRvDhoz+ngMkU
tZEv8ZwR3Fj/zwdzTjj8JErD5KgwqzI1/AbtDDUXCqD9QXq/mUF1+dC0tpjM
B+Jvgqg27GySBZ4dnnKd6vbqtrF12qPRjYion8GJPHtA0SUCg4eAgt7PIHzO
YVemKY+9Nkz2zl6bQ2vrG/l4aoLzCmTbOjGtMifCbSaBP83Z7fvq4dQCVWSR
Nk0kaGW+rWwZBO4cdeTVTX9ut5mx+66qSqLGiofIRE9pNcWD2hawdpdP+mmS
EPsD7IxexBg8SoBpMWpjr1/9kNAITdVDoRDK0tSIaQIHP0eVgCIq+yxnTGXH
BqsjhKM/kR1/CvaTvsYA8X2Z90MXouI02S/47iHleE2VOji9rsXSigvyrbfb
qMGzclylDBjoT2hXCD89MB6sYAF/7dpc258HOzvptS0UtF5PiIKsi1N1lhYX
TPp+OIDXKE/ekVtfdjfMCuiwBUeoZZZt+DSVg4qZc5LGhS4mF7KeuMAAxfj9
XhZBTwrTgxIIqDQCVGVzq5YX13rx9t/9z+AQcX6DDLTFlV48M09UwBuAM1wf
UPrO1otUClmZHMb6KiIBTIZUZNKYXQ3j0DSDGEuF2MgI/ZmRGLnljaIAVU9N
wx57DmUFDgr8sd86yiiqfb3278GzDkq9giJSRMIe92f6OvIFgrqFve4qBdM/
K81z7MsSYfSILiBBbbHOxLNR4ADVsXrBibmLEhow21cm3BtGkAdrsc4N38gF
vPZ9AuSFteHfGatmKEHD0Qi3govXUaZ4oTgj+dDbruze5eMPMLWA5Wm5K+t7
9fd/UECo70uIhRRvPkk12TbmeervX3A2rMXsNXwZIjGZXJpZMd7DLyt9pRsS
HYRzfwX2yqQ4gzNQ9yEh3Cv5Vea55eh0BSABLYXHEBCB+KJ39lZYJizMnBas
IYNZCs5ePcUydxtPiEivdEcel2zvUQzFKUxytr6a/nH4x2ktseEWOX91BYnY
Xyu1OioUbky1FCPJIoNu+Ob0K21RD3rx0moaq37ommPka8l9u5MJdBGR6oER
R5m8pPcvngahJCV+ATpBqD49D6Gvuq05C1IpnNX28PFCyNz0ItJZd1ecU22E
pLAnqX8xJuaX85dX8ZlIL3sZtRGVcKAkg0DGtdcl0vs2z3igmF37gP4JMV2p
c7sOyDzF9q/ctATmjcQIXVKoUYH0AMPBeEBFnF7v9MM9yWUxwX5pNGAb2e07
N1KWkIHUFwm2V3aJWtcsnqOQ0Iruh0wYHcL4KeRK/sGprn6CpY9TPM4k/KLk
ubnVgD0DB1CU4h/xMapRtsbRK38kokKbdrirSg0MEI8nXZOkoC5/Itc8Rxrr
C+6Z9hdl4XsbJ0U7rymlA08rLqDw1q47icoA614CAkOlYa0ZfHBVM3PP1HoY
hATr5qkRKCP7k/E6MP4J6TyKWOhVeoSwdIlTiIBysHfJUt0k2V0BVC0VQ8hf
NtIBPQP0tk6pyj6xkTUo1Y4wseOOIeMip3LalS5xgZQoG9DkuC6Y0C4PbOWo
p60gbsPMklB5HzAEoYAQn+3v3lrdPg+U8EdJABJQO79MDqS6rrAHKQvD3FTN
wFrn3Y1uOe3BCnS94xTC24XhAEi4BJ3wBjofcNiier0Q7czRdV0MXmkmQWfs
ILwj2bAtnKK5R9mQWE/FuO5bBvW2F1wzTzFWH2vXGo9eRY8tmNzsYvfO0RO3
0a87wi3KzkUIGGWly+xxzV4msql2MAvfYcyShcbh6Ay6wT/g6trZIZeOr9g0
K9sPYQvRK6TOikWTCqWIP/c1gFdQbb3nsMu4PYdQqDuNzjMlwHN9GokDrf6y
UlGgfWz8OyQydYffXvvuh1+myvodY4uKo4/8VNnB0Z3vJYoATUOLYweYMpT3
7FIxMLcsgzNRKdbuR/Sor+BOWyFtN+y7V/MHh4/zQaZ7uR0sxZyCPK3fgwdQ
I/uPzqOQi5cLq7xH1mW/vT0pzERjyGy0Ic2/HMaN1u9j9Ub/kaoO2SZMIk6X
pWzEtJ0YRzBizLEfORN5plBA3DMCwEjF9wrvBu0TF1c/xTJIDRmKtPrWN3WA
JLkAFeqea4taAdH8qlzztZuEqoUeF7V91n+6tmvsYolHf1Ttfky/ONC/ynYB
vY8q8jF4PWieg3jcWiSlCmhFrMNRpeSOIO11uHmwH0P9AByPaKNCw3tUP548
SGO0CfZor4+Nb66PbBfw28I/pKLxlJfoSbtO0oo5jnCy6mOeNBNjd307J2n4
mxfjI1fTkoRpHASfMnmhJfZK+Ewy48uibaTt44HG1AlgnDoRLVodGws5lssk
HRf6Xl5rXv01CX0G5j1I3QExI4AiAeyqLmQT1skGk3tUrnauGVDqZnfinY2n
rpoDfUQZ7WpK8j9pDM+EA3bMQX7vv7se6+UHMICjjudbSA9GQPVvJNBKOnuu
Wm6KVb3X2RMx7FK+z0f+59GqklZkAyzz03lpvIJZKU8wpsxEJgiItYhsklWu
FmcTRPJDRWcp+5kj+yHO/559uUHipUEUn5sOko+4kKZGWte45CBmcfLaO23b
SDAePDfDa58O6umHLZigGbMnsWB8A7xCtLqCOwEasJ5LdjND3+pklRp42Rij
/YcUw2BLNPh5tC68NWEIUB/bILhTWYUw/8IMhyFR2qmEVDjje/jTzhY+4UZI
YFD4zjbUR62EcmyuIb8qaKZscm0yHEXGn+0BOe1ka0gRPsMBvKWZeHuuQO5P
nkAAIAlUtMpiWLgStBg0U4rhM0dwo+U+yTLXMdVeA9OFVivegDqsjddgf8QH
Y2gAk1KjReFq6ISKznDHRcvW88D7+dqfAu0rgtwuycYgP51VlEz8zmwD0JWv
nrDSr5wJ3kfYIrW1TV9DpgXlVV3i8FqqIlk5Y1S9EHT8zgxT3vASLenTajcG
dBDt2k7uH5lRhK6JSBHPXofrDKlMv1+ovQuITrv69iQBnRv3PuI+owirT5qc
gg5okkMuJc43a5n4KpgGorhhUUTqgE8qTjmGtDo8Nb+uA75GZuRz0hfDwPcY
kwWgdswtG5Kg4KYBKS0npP9KkYF5g6QAHwqYwC7IZgTnNk2L5eSuizniZnVi
Ns8A6h1ZdaUM7xhuQeubih9TESPa360ev766cOI15iKlLJe0cr9Btx5nUvEX
jnebQZnovB8NBGbNAZDo1E93XAPwndw/MBDeq1EH7UPzOxbFR92WW1QYWzAN
ajg2fxkyNAoxNcfqgsrYhbWehPKGYgwwA1kHrf2zM1wXqscO0QuFDTm6uLgG
ceEkZpUMS2FG+CIgCaP5MHmzy4lWrApSIYVYKxId3dZ0VIrpzUJ7PqsguL3h
J4dWgjnBAt3Yzs/Oew975vTxhMHXn551Pz/4nL10YDKj6O7GXfi5htRLeklP
mrkTTARhQ6vOwYJU7B4Nq79y6DKPWiSWIcH5EedpNQmQ33DqMMr+bE2Du+ui
bwBh0OzojGLzraw46r+u2sZZkfn9la6oE3wLfEB0io4s6uFjYqjz7CxSTjjL
SJOPCkxQMKUuyP63VQXo/SF4Np5+wtWkpGy4g3e9FgLQP/fogiQqmtd10w7R
jNoWdc/DX1/IprxO9ToL7WCgNRV8iLNsU0hYk+3IxTShYDNcr06s+lsTvPBd
R5PeNe0EUg0wLz7rMPmV68hhsGiXICGMtD6ZMgvuwwlfi8ESYJL06jcHjnBx
r6zKngKGlBWGo3uGccg1xjSm8GrvTPitLMHpe1KNw9bkCr4faOJsBFW9Ijri
P/Evbf+n5iR4Gbx+00o0Nwa+I8PtFXKcXRKwzIg7r/tvLhyup66Sc5h7Xybt
bNl8cssbIN7A5c07sL4vvCcSStv7fFy8E2CcGVScuv/eurX1JPDZEhu+D5aa
HnmySpU0sBXnv1WI3Hb1JifjVDdWc4qdQjci3abu61O6woLA3bIuIBMZNcAQ
wX5NXGf7uqTSkz2DtXw/fgeYCCcdJOVpz+1WJ3xNtc6lSVQqyJWO+FTHeFa1
1rWGLvc9tMkRe5CTJWX2fJsmU4jEGUccQkv5jsC5jx56KM3JBAK71VrxdE44
pqe/M042OEiKKahwW5bZHad9LWH4Hl1L5G1jF5QGsgei7K7VT/pHKqtI4Mu6
OqUOrsi6yN37ybaZFcDbRn++Bg1EVsYdoueZ8B2F4MslgxaNDU7WN5d/5JF7
mw7XjnUgbiqsbyYggTdgsqOV9K7JLGRw9yZ3npmGsbh/50UVImZvNE8JPpaI
TmB6EoAGrKDQEUL4Iai/D7VyrqgpK4n0/xSqkk7vfn8X5MiQqDy5nVi5EtTK
MaN33L4iNff9qnfGDzPIBLuUO/v4RlfyD8S6m3pomA+d1XGzVF60Q8B4g5KN
ZRUefPhTKbigf303pyD+Aq4FXEbwpNt048yCEHCK+9zK+l8lpkD0n9RxcJSL
RwDBst8Rv3vEHyNRdNXnYQCIll7GaZNNmQyNbwYiBEVIV5uRjtB+1CiVms3H
1xN7v4C06cvDTdRCLCVTxsO5c/dnaSYFG15majyyrdj1uHJxuvZrZftWq7xd
QdU8H/Vn/pRdpSHZX8Tn2nNVUWCWYjRjBBzfEqzzGFEGcKSVhJ3rh5/RSBcf
3e6arNsI++/ku2WOKSLPxXIoBH+YQAtDiTx0wMrk3IbGDhveK5L9fp3ikK00
dCEyNvUAjA+xXiPvCSpZHXwyrpemIyLYlSSjNoqtTknC3LBKRbdinQ9JDrAT
ikz392hekoZTzGnY7eCMBK3YUY0s8XuDzSkyIFPMSasR4roOtkCUYuZSnjCM
wsYmC7PZDAd6NBQiurJfOV/auUHvMANrn8kP6pGESJqiogvVuSaw/1hLZIf5
BO1qDhwfXuDXQ8rU5ejzkujgeahJnnOfOzCahGygWVOawTuyKTzbVkXX2dhi
dvvzcjavsKJ/B5a/EiJ+a83+IS29rtTNdw+LhmGpA/oHzf+AKKCbtzCfgvag
/AhSfp1ay4v+PJkasXcbHlucvzF6ASEDlwj3PQtWY5OjTN4WZve2ilJgfqyb
a0ldsKDAaACAzh3Iq38vQurZPNvY96V3ACO9NvWbM+Z6KXuxBWYozytwenQd
4Yt1sW+39IXtYy/ZVBCOYiQtnr+Jj8S6/ocahwD0Cyx+PWNEV/Pg1ee2mqBL
7HB55ZQnzPsrFZK/6HPzRighhUDYg1L969xqop4AYxfGFWWsGjmH4Ga4XNMa
V3WRhF693jkb+XZzK/lNgh5Spd83vQXQ9tDPifrY6pdyPtd7JwheZzqO5lsn
Z3eOYb/RwUC4AGqonn9sLbKZgWLzfG1atkZZnJZgql2lhb76batd9RUk8DyK
PX4AXM/5DqpE9L52mardTpCOuEWNFl365vSLi+KUIl3N361vTtLMd9fJQNM9
+SX9e6KL6w0V66OjNrD00/J2q8HgtoWU3UBg85TqzKeGpLkCYO329VZafYxd
n0C3MB2Bj/JC56QrZp/2WsJ84hK2/kE5J0qFShgBLkUq/uhCrds8TOMuNb8I
1R1vcNLFSUKKkBFoylX8Oe8s3o2In75agvhZX4PypF/+9/XLUpngNoQNns8R
mDHC/yN5vOBfBWysz3Knb/r5u5fVb9iN/6hLr76+AJAnif6xMRl/Q4KP+CPk
v3e9pHvzEdZMKw577fvsEEpE86oJrnzNwmYzQn9fRM2qisaLEJTguyJSUnbZ
4JgXkWF/MxgR2dw+ozLgzY/BmUOeHZOFcGwFg+562nn2yAoRXQGmezrZUDdw
IFjVEvrDllqzZorINhql1jN+noXvyFlQ72xDVD/viNFt+FuVNPuQMFgL1aGE
aiOwrNDJE+l11M3jvzZ5Agc2A5S6R5Tqd6goI3cSIA03hw08tU/joTx2/Gc7
TnqdzL4881vK9FXfSj+IntMqP1IbUSkShl9PhsNkUMJqVbFx0fVX8fl0HoWX
rJ/rmsl1iS+mtLhUh5l54Hm9R+Tg8nnZyAbD464lu7KPLMsCmxqOmmnFeoQD
2zDohOZHCKg/NYwkC9dfKctFxblrrj54vTh0qzJVJh8UfYzSHvVwHunCbcyG
smgEhvE8jQXpzFhfEKGyvAvz6ljmUsE8Bf6Ycy2f72HrKl1cHroqOA0UBR5M
5kFSsh+0O/V3rIEOjJ1ljS3o0ZHetDGUCN9DikEdUUqUaTs1YTMkH7ZKAI90
v1SwUMh4xEmfjO4cEj0xt/6ZR5RBjoSjnnNgHfCgxPqq2NJLD2WPJRUDO9Es
dlpaHBjb5YzOL7y+0l1LHrmQ4jXrkCG4mnzEm8bNMmjBgGrOWLFiRm9zfyp9
Bvv/BbEpeH8IiBnTNl8gra2yBEI8gYKYhqvbpyq/KaDeMpPrRkGWtMZuGzjA
s2OE4v7uU1y5gEdc+5gdnW/QSaN4K4QD/Ebu+v9HfpRGwrOeEVg3e+hijsOP
Ed6baiIqI4nM84/yZlqxmM5rHXuZJ6AewQE4PpAQc4Oth/53TuPJnRwIE8Da
7qQgeGUh9iR2lhdF2iaPx6MwYLPETvre/0+G/U6xcRxqm/GEI7xC1YcoQhTI
L2F+mHFO1dcac+XUTy0CCG9l2dfQFbM/PDf/bM/RhI9baW8T18Da3bQ0dyzu
wIjkI2q/QTUoU3j82x8SELj69x+LZkz7InSWiLKoNyxXL1thn8VwvemZAYZe
drKCPkFv8BDctXXuvDBlUPoXv7ctMe2PVQaU6F6vD3B22ERQEi9U8I0OCFsY
Cb+rTzuPWybO5z3WMvAJqeU1gUdBPITY8MLRa+hSI0bHAfgJX8No444llRXF
Aw4HcTNVFYp0tKJhEXeCA++f0ug/XLyKFaQPADqu17jONOfue7SzVAH0NpwI
JmHOxjE9z7pIdy83Nu+MK6blwTU2V79S6pS/JZTYBqLR2x88RLjmHvPw8jrw
6f0Ewz9TQ15x2MLCZoB8n4HVUzx/ZpdCG4gFs/n0enwjyFk242fqukfQQoEW
uy6Eord6jFrZR8tUdCbhrnxYKh/c8gE++kfYYkuSsTC318XAIdubSdm1bIPF
PDn9xiQ4VuzwdTK92kYZjjQQAtE1cbAkBhfxCfiae7VVURV6

`pragma protect end_protected
