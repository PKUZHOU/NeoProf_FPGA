// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
AazHe0QteMouIA5Xsj8jwI/CTeHTA3KQs99s0VxBPVKWJ0qyQakddPe5C70BAGv+
vCJ3rsE86yURfv1k7aTtfBVnbrxrK55xO7iVlUpZKJzNNCj7VJItawYdNAKz1YeD
SAAPqOfJZ6aZXdEvBb/O25+onAEPiv/8MPeAzQ8KH/An5/pALhD0Ww==
//pragma protect end_key_block
//pragma protect digest_block
WP2ARKVXfrmxWMaWR4JiyJNXOiA=
//pragma protect end_digest_block
//pragma protect data_block
h9dVDNS0R2UK4Oux5WgPl1g7MgjK/IKvIeUl1Pp0f4TtX2B9UGaUSQDNxxq0AnBt
OnEZJuyjI8xoWbjdOvtxn4GLujZ+kQ2cDh3x/GE8C2fDGtKja9DylAtCr13b9svH
El/e8GJMqmzV5X8DlkZy6Bq2QvXQvhIpjIm3lwyBCCSoFWxZGYB0iKKDDqB7c9RE
90NJmLCpRrnhfb67qjqLjKP6VPOuaSW4hiavVKaAMS2CSHXq9wCHis2L2lntKkwj
W4+KrymPJvtaTadKNm7OJLNBxnKWSM1ZaxO+K8oYnFWtR0uq0hefI3n+Jbla/baX
UInKPnhl+LJ/BCUuPoFKrVEDmcr++AKZ7rJR7zWYwgJf/RMLi/xZrEBq+jwzpEdc
xFSPS9xo3kQ8qUcV+EhxpJltUzi9+n2uUmr2hv8x11bGa+cJVz8/pR/7Ns5BGZdY
DSM0Ekn4HSAZYSSymzvjUbwibVak3fVgPqujVgg1rOLxw9c1r33EuOcO+1Wba+ku
lfjCgi7Y8Unn0pme61WG1GyOQm7vkIxNavEyaAehG7rFVVk+XDs1QsEk+qZrUELG
JsFoocErU0VsJfHoCnl6AATdF1tTYvyVTUNRucX10EZ4QlJcM7tYmvuHh2vuuYdW
eI8q1XRBbOK4BfDVvuGclZBuGhDRPjz9Ipqs0SCf1lJ2g5wyBjsYLqohofk6VkNh
Qw+9Yu89ik8crYvm6xxLFid9zNL54SyoRBlBL6w9P8vsCNzCOaH2yxMyWV4uv3uZ
XbZB6wYz0Dt9GkI/f3sGAFsYhgt5EcZWnCl6InRP+yZLiMJErEjZ9p+432/EGycN
yHxWqLLI/tm+H7ZyxX2CfTnck+Bg4gagsmhpCM96S3uTdIWGphsA8MqaegFkiEZ0
Qg8yjdvs3vBL/ox0TeI+UzbZhxACUms4Su1V2q3Dq9dI45Ep5DKxAGhGllp57AMS
Rv+V9laSW6T0HHPvGpifnTi+f5s3nGHKrbl0JF0nlsMLJwkIe9CCsojB0jBMi7Wj
PH2cEsoa0QpN2JLndAG/5XcOBosJ3uY2hd7DGMo4+iJLwn97eSDnVop0doCX2i8a
8IU+dM3YT74ZFv6jbFGX+cumIN+rEnyC+ziTgtO2OghiKjuM9mL1fozmlGjBZboG
1l3fV/btkZLLuy7RsUPVwcD4lHWEOOkyUb196CG+6mZM6T4jDZzNB1dcKGLgSeLc
2gExl44HFCxVV3bA+/Vt7azVYz3i6sKXbg+a5EnMka/pWLkyw4kOM4vNzrIZ+MTZ
iARPofDkY38dbTRL+s6796ZJYWtmpRZIp3D9Z2ifUBpx1tv6iSPYzZq28FL+E/QB
Xx0LLEFBiuhER6Kqdf+0ozURCAJ3C/h2jlelTs0N3GHNx85rSNanRwtu0LUKjNKN
cN24JE8+mKTKfKfLcNewTWwwti4+OYUXQdblVUvbZu9OLj6QKM44YFQULdz7r6Dj
VpTCOEh21yg4Z7BDjCIGqiiBbr8kEyaE/adhJ2y9JSX8icW2jKh6zbQ4B0Com5Xs
ob7rBFFkAvTTJZnRomYFHvMkYTveErZ62VZ1lxO/Y1ApgWtC/a5oRDab1z6jTftM
eE2MuXn8P+NmuEwKzgpl8/+hU69JUdXX5te7huq7Z4xrIqOAkrQ0yhzf7OqD7R8x
n6YBME9Sz6jOqPe1Up0ZlELSrv1b1GSkqdWKXvg9s4GasJ6a7bcqIlgdg4ATzOab
zmow7apuqQz7B25NE3ZtP8xcAtcOfSihy7feUYv6VCiNDuIbCWIokAFraGhYgSmQ
HDKPeRnWYmwBHKjrhXkB3r7ca0zULdmrKEFt96IcSxTkrQuu4uSTaeq1l4w1Emq5
ai+cY9HzZf8cm+epYVJobOSWKbXUWY/kFb7t64TpoOmJ23ukyHIShl7vq9BDluik
jg1B5WaTkQgQUF6UC+ZsyUSGkHPLQeWAhfTzGecESKAQcA4MuSk2Iv1hIyb14BiD
nyjg2vuyZWJeBKVCrb6lOE4aEByQ6BpoRdnfOXx/+Ht4WOeY632+8B4gL7dt/VHT
C4ek7jravXgC5ao9pMeEGxyS/xhq4TqHA5ARezEve8dv3HG1QmS62OR8l9y+E9DI
qdhnqmny8Uion7Q70gIvzPlQT8Thx2mNGhQR6c2hSjZHnHd2IaQXqew8u2h8XxqK
E7mf//I+JnX7kfvyfG3ye28PrAI4+BxEFDrb38sjuaIZSwF6NiITPeUw7IMBOwqV
0Ktsmbo241cFJ9ApR5xTXSN1X3S9yxsIwR0XIsOrCinb4/i2Bn7D13N3wbKixdRn
U880OralBJfLgZcoeKaFV/EuzoyWLET1QSFq7WsvcXqaZZU+WLh8sZSYfRbTiQ79
ZlUIaDVx4jTlD+A6QlVzWpe/BcxnUC1WkBDTeu2XoXXrD/ZWXt616rlnx700XWmp
dUJOwLg+SYgmyhQoJYMfnlBCwfyTjATP6M68RfXa45OuLnYVTqPM5PV2DQAD4N6i
l71HeIQCCPMkqJQFRi6/HU91e67dA3JJN7lH35B/pWom3XVWKAswMkezYid5/kKE
4sJQnzZFSFaZyFbEjxcE+mpOaTf5TZG5EevZbJneGf93bFHowtpNYsHnmKd+ZyI8
F6M3+0I8Y0Yh9PaoYSY4uwpkb6FuiVSUNhuUEu+gDg977tPF1+EQpoVTgT1TUXJt
Y7596EAts0xeXNjpMJF24MASxz23elxDLfndeL8qGyRhruzUcVzVFejaFjoUmIjh
mc+VKf4O0m5iccrACFRvD1FJyX7Pb0Sh1vOo/hdOXiOE5fAINMARt7FcKVVvxfZt
Dz1072WjtCist3zjWqyL74xAKJTE8EUdhqfPGTm/zKSoG1Igvbf8ir2yZuypFB2K
hI0qh7d5CreD27Xr22ijpk89gGhU/EUm+j90eCA5KSD/qZmpS4QoXrj6WpJZ/Ce+
c7tvUO4waSAMLz1iw8H5ehigs2YV15fdDaH8LcRg69hX7V6idYHcsyxAdr+/9EUE
RFE6rCN3fHQedWDzk/0WYX/iqXQfyoNERyjMUxzlmNLIfXduBAbLQcd1cF3Sne+r
eDOhIf7+I+M7kWzLSFD16S+fzjP+sxjBig4WKekMm2w/qRdGkje9BMdjqtzH/hJl
OAB27cu16jwEssKl8MJwZE3YuHtWcUOAQdPjd6z+RIisFL3mqbJhG2jaGi/L8KLf
inr/OxVv1KTSfkr2gZWMpIFdEP2jBKPtwA2zppcFrWpknYuR16KiGb1+YuiL+ksf
I8QhjgM49XEvHSuv2UNCj+Yop6Tcsdot2NND2pHAfmBJlUwzCrDOgbXAtNYufT5i
3SHId+AN2MIhMXr5gMN/+Wu6FFa+zckAYx2HqiF5Lpu0/SY/W01MtPp7qh4Idi6K
zB/qbkj8ur6eVZtTQ60toSOx7a69ieowM1oPt2AzgrBQEHqPW6psoBkLQC+hh65L
QjxI1KLMQVzhf5gZTna7jBU+IHun/gBqUkX6P9K7PUX6uo7SPdmJwiv8iWkSBP5e
iPhXnu5l+skv2SvuyIGtEPW0qgC0Z1Yal/3aghK0CiF3G1XJr6uOyvT670CXs7Oc
cildq45DlNGnHU2Z9MVHMRpCrQ6IZ90QpLFF9AvyboTZST7Gi8NRvmz5UcmzwkBm
eQosJMW4BKcO5VhAnbM3aU+cxCycb9mTTWXjcJkz7EPWXO5qZHiplRc6V/bX2qGA
uxsYaW1BMSS6dkW7DR4nOAXzKY1j1rRkA00DPlNZQgmHjeti3Zz4DjF03r8j8dvI
yivaqpJITQ9UwjXRZTX/gQm8+9iLrI4wI7Q1QpCxZzZ2UW98oLQpJ5oZq61KmfIi
cwVNDBRtjj6+AnM5/lQfqb0n2X34Yq5NlT4U8rmxaas39ZOSTQ1JMcUwc559pL27
IiqL3zNBUwuaxpkGiMp88TaNdzrAtpzG4jrfiQ/W+oOOTzkhPGPdtlvSgJa9TdfR
54N5oCh8KQSyw3IArZvJmWXF1T9heWahy0v+PwcFioaEv9XegD/b5VjuwIPuOdVa
P9P4XkgSvH9EN3Zcvz4ir0iEiY7iSGeXi2bftsn99qhx13kH/0xiIJDu6QeXoxAu
h6dkWtvKSBhkoMTARJ4CgX0Gtv73kqgjPsf6Pafbv0d4d4jgO+w3nKyohyedkT10
47/lk/rxSJhOjbdsLw8P2ui6Wv9K7LMWtsZB8wnyeiEig661OFf/LeUXJymCbgvp
98P9GhP2wO7T81zp2XsA0VLmJRgfddTlRkhMbQ8oxlOgKCO0IpPK3dc/76x2dh7a
/Js9xsbRHS0Q6/SB6MbISlS/drh4StF15lVEaj0OTOxu7gvDz9nT8nP2fnra5fiz
zZSGHbPXwZVcGWR2iTnbF/jV/LBCSmsGcmsheonxj8yLdHNYBHO/o6yRXz3eiBZu
p7epcBKLdTf3qDRfKgzSXDnvfys045FpbYCh1dCYZsurd45LFM7blRNWO8WjV7rP
cjGgNzHOj8DNGgci1haj9TP1ISqjCroKnPjD9yEKSvv3ZtSZ+fs2YrkpVaPPH04N
46z3iY8sZ9qOAX51oWkuFrMRAQvKoTTSHHrhxn5+dESISHN7FmToCbb1gbtCLGmJ
NOjpsUCCOIfc11tpNnO9RpVicrIRw0eY4Ov7oeejBn/DZWhI6YaiVBZgvZIvh7us
TKnhlMiP/5LvCO2Z0iPe6lFerdvQGDlAM4ZwB1hP6o717N4kps/MtAbA9GFpeLe9
YeJPz/l5RTuETvJEERj/G6XncxrjH0Vx5RcXiFxocsFrqadBE9Vfuy7fBCYWFN6h
gtAYGpg2UaezWHn/cjHWIjovHQ05tueKV1eshoiKcNzF77HBVwjs36xTfEel+NLH
J4T5PHctLjW9z3SRNWnjdHmyEa6O0QQYu4V/m2o/jm6z5eOFlYXE93UiCUNF/yPL
KwqFv7S2jYVrGWbdsZx0lHfMHvMmY2BsnVscuqyQ7QmXz7B6wuczkjHCeq+bIFzi
Ul/pMgRlBTumW7QlZKXY4ZZTJ8zQWVLvYzG+6+aOYu3B4WfYAnPXmg1HtBjUSx9m
VWYofe3JWdGu0AqgSVOQA13owZVAWDGfI/yMk55l+gKX0vWUliVevgiDsZlff2YD
m1rQ1CdH3WMmgcX+kdsQ86FimpNjL0hPUp8NkzyCeQAKn9Dmk2Z7lP2GB9BFbAcr
R8IaRUlxaQySHWRVU/xIQWWB2UMMJe7ue9YGV/QhFG60kU/g8C6e10q1WfaFfrYf
Aif1PEMEALDkZrjFRJV1hfiMmV/gFN66UZ3gclJ6hHtUl3TJC01JJ7wI42OtEmS0
m8wpFmyWbMadb8nwTiS5RT5PJgWU55smh3ai4v6ZIUFWymF7nb36+OsCCFEUa83+
oZgpU50DbKzsaBxdpwjizfhyIILCPULmiaQ6nnZxBQUN+2meMkN0DXRjc8wDVXwJ
UCk5Y7+T1QMzf4Xg+papiP+G7xDysGk1YNR0mz2h1/VXrnB1PY4Kuk2W0nOyKq7q
EwD4gk8DhUD+jxpOfpSNDo+Tzeh11uLf6YL/OBMMGA5yepeswm9btXQxjyTxCP9p
Z1QN8BE774qDSqE+pcjSXNAR9M8d+qpAb64JV0aw847yjfPc8AlEN32ZaKf4k2EA
uxrvotbGQhWVoc7aygEniz6mS/8WbsYhs6QEeL0rwSGtV872+RNcDdmuGV8Moukm
A39HFCBInVxKgs82RRJFXxOeNppxyo7KNmCh3QY17wmUy1YA8ixt7gQ1E28bCk0r
yXN1aXMDh6W9N9OHZ4x2L9NlaSa10MYBxfLvYA5XchbRhATVEBrc1ZyAfc+UnHm9
40ZlMnd+WNgtIHueQ5dDclT+T8Z0ktIx86C36137dgCazdWcbCTS5te7kMUObc0E
jfqPLeMLWB6JOebRqEgRkiwThgQrEVp1u2WyHtmiDJVFhm3nDLjWic732Y+NJI8m
x6JUT7038/VxbrXLt19z/oUpNU45I0BizIsdJxryYgEB29kjJob2Z7chBZlp2J+d
uyBbcX3PB8lUgZA/zfxxYi1+yRNqILf/DsoHqJx1uIOhqeru2Z18oF9Bs1zsZ30/
lvUp7rhz35OS9xN9oHiXg6V7sQ9RA9YjR4uRJ7ulV049wl8SoLIqaG3V5130vwQa
BPV4RwWD76cxBNs40CmsEZhu+trOfBKZFqrB0ZMB1TYrPhNyNJypQKVFwGyKOToA
JyL4/e7JSOmR6KY7xr7YO7/m2sylxHNVA5XvbZ4NRrB2D/0RiRV6dN8Je1pyh2Vj
er1fonpH7qbX25iyqV9ibCkYHKVmG/PdK3mNyYIoJ9KoXXnzdeuqjVqXTEEFJ80i
TzMnrXzNU4pPv+a6tOjmi4OLlxB847IHl62l3/bQ/7eLmW46tKIksFtDENoNbU7u
vbchlTcGhYZ9cGubVtI+PlcaX/Gt9eDyK3cw/oY69oXYU3Zzpk1equc8LH4umOsb
zOKGYubWSgVw5gh9CbroThp60cZrixp+oAro22t9uZYSYgtG6mN1ceruMpx9ozG1
eiPCSX11xHdUQEaUv/ns7yQ+LPMu16EJlfF5wowJo+/ZnhS0Gkx0726uoNqtN7Sa
fWu1haxyB2jWBpC2fjSrGnBl3b9eAoCB598YAyJPLSt6RKhZ38g8g8JRx/1pgGO8
eX5I0O38P7hiJNfucDsA24ah74Qdr7wrTYU4S7EdJReBJHdMjoCcb6hV+dBw6S5J
Wdib63D21/HISlRUnb5RGBJDAXif7uVv5XHDNS78wucYdiG+/kMBWRT5SP6h3NWo
BVxIXWIpV72UECK2bdEv0CLTKecA6NrER5sjR3zF+9g1jXUEpS7VgbXapODJvv84
LIfJ54m876F/KagTLAkjPtWEFgJdy+2jAO73CntKj0vpvOObOBQ/6vplFToYyukL
uxJoPxy0vUmEQUt3W/9TzaQ55iIcNlX4leLwnTDAoBZqCRxcjqdZw8MnM9Ee+fkA
Xx/cNwGZMhw+coPUhAA6uIh9S6MugTn4hX38h+IzhIDzjqPWrFRLWat9Xg1MH5Sm
6+io0/dQcvn5CsmTkL6h0suKsWDUdFIKK0iRe7I2ZePsOkPpDWGChaOyStOYPS7b
49t9M1apw2zCUZO9qWVUq0z4+PbnAr22hzVrknsGZaOjiCsyU0FPtJN9yIosyDUP
yDZYqBruwztkrmSZxks4/cudRlJF11bXrdSRlZlOVph6Ak4TGR9ky2WZAKPwqwfs
8NliFZ1M8GYzO959KT7+BGxBN03N0xQGsHz/JU3kbbqn0i6JoXGdDtbyhMLruXSn
e2nSFAk01xu6X4ga9vy6YX3xtgvS2lZv5ll90ZGVdaUv7ulTj9K8GTPNjQkPxyUR
B5LL9RZ+I38nt4J0dmFjnubtIYC47JLn07n6h+t9pJSGOtA646Zo7TWqXClpmK69
1t6NoiusxL+p/tD0iREpb0kagkUZU9XJedO2+ZNzN+ZYJsrv/0OjPgI69//wMaq6
3JPOZyI5yRz36TPM+bNO1jcd6GU+5DRT3sN6U+kkhFit8PHGnpiIKkY2S2oH7+uT
eckPy8I8wUX5MStilB8Kn4BiPV5gI6Xre21hF+Y+DdRj4uw6FpYJBVhCjtwzQA+Q
08l3O0H0ZOHxMvdRBK6611JvK/fDCECeiQfbcIdO0S8q7pmntnqzPqGkt8JnC+aY
jD/S+OkRDz8MOPxMTUfYB8CTVa0tr7hQgxX2n3TmKEl+CTAHCM4FSqebGRXM1kWI
JoE9MOz+c/FV06ns5MqDQoEX+4IwD1MsVnBJUfuhklCrgoHBfYUu48dXon32Q9SE
5phEugSeyqUhahht1ReOk/mWzC9MHMh23N8E13e+VMjQ5Bj9yGV4wDtKh+odIH7p
Ecc9sQtnm9BspiWXg15Z5FVpye42uKYDpxnSmCNdgM8gWiXcfG3QKPa2gKJ9RTMj
Mqdeqijw5XFYCw50bpJFLGtQSpNZmQlFbbf+gPHrUkYYKKm+0ZdnJC0g+1a9f6py
aMCx4bdDy61h9qyTOgfzii3e3qWl9Tt8dwuhMcBYP8zuWvTUELZ4ssZlJejuf0Ov
zxrnaa+xiFx8ZpONcCNu5kVp8KUoOHf4hNzMyvdhm3UimdsEffNm02fVGP+ysLMb
oTRXrmeQeuz+MSsY6c8ubpt1vXlyyEYUFtgAK21ZvOMKZ/azd5SDb3ML+7goSYMp
OFhclNSEHEYhMFFdIBnB9HsSk4GuGxBIxnpokC91qmRm0afnNyq3qY4cSzynyaN/
jHKDEu1mS1ULcBG9uNuV+7rWdbP92AF8ddIayMGRAMInvu6GnhYZlEtT7W258+2l
oAGHOcbeK4P5aV0Ygx1EYJhxH6bX/GksTxOrhH5Q/TAGl43OCsOZ7ztXTN7jLU2a
o/W6Ir/JJtIzi2QOPq1PLXQVE8p3FEDzbv1KxjyYaLYg4KvetmSyupsilpibzOA4
t+eaglzOpBJK/+YisFCIXH+Nr027QotO8SsQbEomZm5SVyE6rXWuxP38pAwYL2PM
EIgeTpSc7JHEduzG9/qg8CtTNFFz6+QIs8uHLeAVCfsx10yEW82BSqRQrm2r9zmw
9h8BFHbAfRUemkDbTObCU7GePPRoD0sWxIQgomKCWrm8BEh47y9e6Dbo+WvTnSkV
A9kwoTKFeRfd5arjY/Pvpu+fHWtdQ++PFQcFL4K8Xi4nPaA9NVw95HSqk00+sxYs
ks9i0KCBdpzM/uV+LgOpphOPP/5FGKKIWW1fJXcsGaK5sy0Umw9E30GhdLT1VSmD
hzV+XCDngKDTzrsFT/MVKGl5woWBdH2OFmmvj+CX9IvcXBuZti0agKaujzcKddTI
QVkH346qtajdrJ1kJzudjirI2101qvsdlNrs8YDqMCqIAqo9z+yMiFHpfC8eqAOn
7/CsaggM4z/scdXTYgyUeutKJPVSJ5JkYC7nXwjps+CV7qGulrLIu9x6ffYhSDGi
XTALCo2JP8ch2WYoHXAqRLStblFemPf1vxfby61WUdgaSb7CgdwtuZOaco0B4UMq
a/z/n52lJPNNMt8qFgLkC6GSJG7SKEpEG+ngXmBx1onIhQjR2t+BWuuwks2PAfDo
nT77tEjkF4+mzonavBfNEdYdgDySLZcLHTO8A6mfelY97sPtNqZKUgJfx6Mo+WFE
XDAgubn73K9RZUGEoRuY1sbBCXlnbJVhXh/9JWK+eikSzVUE3T9v9LiCeV9ond6F
EgIGtrNU9dAplxgreJyilZVkinRU9ulm3UnpJ/oztgIRh0zIxmFvQ8FXNOlwgFWR
sQpmfGeMjDPQHomhd7d/MTO1ZPiL9tWY4x21Jmd7WQLDENehcs4NpYLhHUo60Rs5
10F8RbqrfyLSCBJkBMDq/eUVlKecw4WrwHizK5D1OXVOcnrV549QZ0Xe9lAV81dq
dMxIu3wa6cAtDA8c3oZssDbc4sivsRZY7wA9HsEPxv+Ka6okdOLXkBKBF342SsMM
LbSUkEaCN15YLC6M74tYOah2xChDx0+BApsqHPJzzjsYZMD0KZbbDqAHr2//7Mv4
u5QBTTz9noVr1A2LX5RHLK0/kZf7kwYddadu6h/8AnStJkBdM+5qR7WbGY8YUEr9
5/SzGLTVRUVEl2OGstzwzXnegbB5BWksoNBEpbQ46HDvmhrSVW8SvPz/Jq+EBCv3
mvQsQtaHYnwIdbqjh1WH7h1ZNBhih4Nr9Cs5+Tmh+mmjSbvWMK+mLV6JsMwiRF7E
NozFk7XIlYc+/HvWI2+U2U8fURX6a9/usKCjaroxBkHPEzOsFEzZSjKeq8SdX0Lu
X5Fv6MrH2w0U48PUonlOTMTpFvFFhc6UGifCE4R7Pi2rDV8cykNcpwM/TK+P4AfI
pmqwE5Ul991+MrvGlcAdyFrNj6r6tAugLHTUFrQc0tq9/t2kPQsxNUFqJoRlVryX
XFfFecjg5sa831QSUNPlqSIYIqekCBNLqfAzDeaMzHyzdomoQ1CRPOff60aedcmO
KBjje1OUVH76N4H/cFRBQ6gklu+zW6dRqRhfjstFnXVrblXQ3UBHEfE8NtYxtDvK
Emcl5qKo2nBCM7Xf0l+z57/6uuEDHA63vUPfzxy6I1sOnMPZorDTb2SOGsCtjhgo
05CVpOaAQ63HXJrUc6XbXdTiAVSqLS/pf05ZaBvfqdUQdqxg7m/lX9VzBmX7YUh1
W3r3A+82Ys+brc03oHx3L214QD8MH4RDGhCAdWZTQYbfUzcWHfY/sdnhYmJNv1cO
2e2b8HZRFZ+EdOFG436AP5IeWcTY7fYyfoLgbb/IRGLP1ZhUSp10RgS0GUXqqOmF
85fQJ7WL6YDbby4NZZ18FhoWMsHLcWf26/VIoNIORo6Y4BXC9zTn6kAP8V9UxLAs
LquJ9WxboagSkSFVCNIAllMZWOHXBiBlWskwescBjJGuHaZxT8VueQDxjzZzZX/3
J0PdBlaWyPwfi+6izjY3VReravb4y/21udnjAbZEDoHrUPAtMEV3KPGfBihBVCSR
DBOtbZTuDkNYhJqRzIjcIDyP5B7aBApwvDmkZ+ocRb7bZR3IBmIf/Vb/YLBOLl0j
vHego47OBwbFytdMfiY6aYnvdZ5Z905yjIB+dqFo+/LGs66o0cK2QnzFcwNSWuOe
ZqeF6lBXRvT8pOZKaDUwLbZCDZz+BxPGLcCn8wo71nFag615fySQau+j4MkFcCmV
JaQ42/GiduxlJ2LxlUFHdyNU5oGSo9kizOUEaCMeMpfW8MSNHyvxkz1D19gaofnP
X0pS4PX8+vltca2LP6wqlW5m8lTHPbAj8YhBOxxGdOIiRxka4ruUOUZNnF6qLmKY
NW3jYa9N2bvxNWjl3deITiuVfk7TshUyK9yg6xNna2PZ99dXKzHjyR3EBT3SR3it
UjaGVqQX1UyrqiDGz38r9i7aKOzcVqj0T0p+H4yMMG1HnXUM0LaBMlxvRfGQBGPc
FjkGt9t+AIINS8Fd/LZ9fQ0W9gkhesZ3g9bxrfiSCxqgypc4MZ9xyl0Sl03CvTCL
NGS8iMxCafdSKAAG8HAysarplPXubrd6+q0RUppey2uGpizcKvh28FN6ESWBheo9
7RhhvptUtPOk5DsrDTpnKmePSDQgP9QqO2N6hzXjPD/eYb0Xq19Jhn7b+XMvTCEI
PLBxB97wyFg4q6c3BEZCrtbjLVzRUkIt7qPZ+H+ozZCrzjxBYSZwmVDZINW+TYzL
ZDqJhjnLLDzMAq9H1uS661bNXZNhOJVuFRKL9+II9PlMyPZc6m4RnIMhtdKL8p+a
gw+v2+8LSW7VOV87RxvQJdnQnkppi/F2bS3gLyemxOU+AoyxDNgntx2STmnyqtz5
JHyHjpBv/QACLwxUjSus37J5B520X9q5YOSUDo9o7UQfemaQHmsKfq0VH3zz9Mme
VIiHQYTXecbzxTG48ClTLKY9vXyGlvN8AS04uRsaiqnagOZZLXOONt9GnN3wkxwx
P0SpCDQw18oFlSizVT9oFgOgd8SUpvolow//sgfJUDxb8cgbVsHEU4VZszoING++
5dbHDSfHbC2/2LfsuZcyFnL6zHOQ++3562qsN5fE7MP8iGpGxRl1Vwk0/s99Mvsf
NcIqvZ0GFmtvgcNBzcL12Pr6h/W/maCIgADHiBZ3lR4ZsXFr9hsuZkq32ivcq6PN
NiL+dmruA9lyMtmaYa8kSgMcYSBPof4+Iw1JCdHeBJFAveemhJa7CzYftBQr45eP
967jLF5+ArmB+uz0Q4Z9hAKbM0Pqf/2DpxuYcLxFwDktNqHuD4jy7bD+S0HUXCRl
Vy2V0CkB3kAOOhg0U6PghZUoE33SV87HFa6pZnaVLJzoK0KUMozn1vmwPf0b/5cj
DMNlmf1e3lT8jeE0+J706ORXXNc5BLuGwNkmt/vY4S3hNzIebOWbryahFPnkG9+4
MtzY7jvLfLyFTQsKTw9uHyLi1nuQDlNXYDHmKj+RcZoQk7HiJWkHXAO3xNVcCrJQ
XAOdXDp0Fp62h9YDPM8MoKXWbwDk9iRb4WU1si34JirUoXOzy5CUGXmu2OcgY4Px
A88w07s7XYZszagZCyh1H/ziDUBtsT1kXDzsXf9iFkrRFn414IAdy0tHsIM807wU
o5k9cN/IErxcuveK0wiP42Dg+YqbXgh91HDvHYcuMAYgLEQ7Jy2lnorq0l+YVNLh
eCGoILetz0hXFyn4OsnSj1bbnfXnzzCUPN7ag9L6zmKOcIQkJ0jv3vXjasYSZCzZ
awceESge5j4gsadkXz8LYZ7fy61mqRkEcB0XK1357XKUrbuWdb6ZXtEKeT0wwTFy
r0m/Rec90byWsNydy1XDTP4v0Y0CVfOpLM0Akk1J7kGM6iJJEXQND7KgXXH0aKEj
5wnsBEHI+su//iPe7bsmlSts5XdgGF4Qb1q7cnSPoKghw8nJhDFSwcG/GXdYYkY0
o99l/XCkenuGZPhGvF/XKU7ltLP2fyyTLUFBWsrsU5y3upam2F1oFQWHiPd9OTF2
FLGcn0vKzdCS7J0HIjqa3dJ98e1EQrdc4xwtEBrsdQDAEbOjJhRrAjoLVo77bICY
KNhsD8UVAgGX3wdnUFQnKHMb5n4TlZJU8fNesFP0pMTj0j2yqnyXk1HyTEPwPF3B
fvnjlYaIEyt6QRyYjxFWWkp22t7KbyyGxPL498lLgzFdKKkuOyLm0skA8O9vIkrA
6rh4u78IBX3kRnMHatI7ZN7Qr0CnIhN2DWXOZmgPoMpg+jMhznGV/vR2zhCauSW1
7xnrcjj1XvjChBBNLEhVdLHB2SZAnaDm3owwU50ZB32jzlZsh3pytCiII/Xgk3Kj
FeqxV91f8f3gUUMrj9qAdOWQwms7CiAVCKnL9TLiiCf4PWONMsJ3myIhaX8850vR
DgvdL9Buj4DuTqAbvbwMfXXKw/EkSEELhOCpC8q+LbUQH1QlFF0DanDTWHyTAcOw
NoIAknd3WxhXC4Ql0bzcK5eqznk8mxpTNRPGHLCiMaF+0/gBdlbfAKYIPROE/Jrw
RnB44V3wmNWqhRrDg0HyTllNljKORz3cuGat8qIYeyAVkfnZy/qZFW7ox3B961ip
S0HuhW1RCKRwWDLMGA976Wu1g7Z9wZiJ9F6xJITNNt+9OHG2l7+sbdpoPnPtjQ50
u9eEtkFFtwtIbS3z+W1T/v1nz4f5TDoq+HlcwZxJDtf0m/a53M6C0txc4dvObKV3
W49PUFQSE9GG1raYlWXfq2jHfBqNjhMxMV6uFWVja8nR+CIubLawBsl3MuPhIq81
09xcLJv7SjE3lW/V7xqG//bFlsh+r1dBhDbgQOkMpIEBO8pra2A1OpID2K0+5Mf3
4IXuTvRRd1EuQz8hgXzRB+OI5H/dPj+s58YsXwVCdT/uvyfaROPcLVuUkaatU7k5
Bzh9Yvw79N1ExTgHbDN+Dzyw8vvkfU73zQyOF/Z7vn1w/3dSaJ1v5A9ZcLAE3Uut
UF2wrISOcxSencHKwiIKEfcdtqphneu685Ek6kA3TSb56EOw1+4cgwWkEj3wygvx
n+ED/EqxlXi91OmoU8cJqtC3qs6oh/l3rTDCGZEtCyc7GJxQGfg0CkIu5FAhpUFi
nyrJjfysMRsZY1bXlYffVj/ofqiVu8bPp3gZpuzo6aUVSHvYGCuGOfM1jIDzvKAr
cCewuoIghJi4p1zTKTb4+dtgDxc9cYtHrF9MsAVGY0OIF1RSYBu2dAaMp7MG6f+j
eLh4X7RrulLkm014y78PuaSmMBUNjJJo0l5sz/x74cA1mjpyLSNytLDHSRxObS6y
UFk+CDzy3hCxTBxi3TAtyMPjY8fzIRTIo/WgEtgJ8zm5bztx8c53U0/26QgSV8Zu
1PZ2S/yJvbW6x1ytnKV/tL0AhazWRvQBTlnzVhu5V1iDJdgtRpDjL3bDEHEuESLD
hh7+sJ5VDwfXVNxMAEVYl2ClXNnJ4VXgL3UG85u4KmNZ79xYWbaA+XDJXqiuCM3b
kPVOUZ1xqU4+UrF/D2ZY4Tic2vvfKjHCBmC4gSZZj7eux/w7SpvBEOrrnnEBjZyj
mRBpLjDK77MkGzIdL1qYj3oDU+928tz0wcH3cPx3pADjeDl14LEGQ+nZjNIZmhcy
2adrzD9nJrYXOaIRXsSL3Qo6njvfik2/nFTUr5DVhDGC3KXR3IP5fUCQiiyao6U+
gIYIwDIMzvtFsO5rim6Xgq7fHzXIWo0Iz5CHzrWHYXhcDNL1OvUu1BdHXrNCeqXp
4bZR7uAoA/+3Al6v/2upMUqTcVI4unOQexrlM6AQ0MuZ7hY2yfNOHfXcPrk6nvgJ
nHYRi7549xoOL6+FUTlG/kumY1GTM/xOLldPuiq5M8HzX9FfQdmeIPoC8Bmx+Ic/
jcaXNs/IFLtpDPP3r9kEnDFQoUc7OUwfuBTVzhWTM9eqcf7fPp6RsQUi+58hS7SN
FtK4fpdlbHKMBZ+yz9VC+BEGe2zCuhs4b1gkxHgrr3P8LBXg7RGhE25M5p+YH3n7
KmvdFI222HnkgiylXT20tbjvCXfMEJ4Y1vdAvApSTQUGH70T2UvLqTEuujS09bq+
rs7WYGY1vslu/Y00L9LnRNEb+SVsEAHm6nLGFlR2J8FB9Skx1rdwTxTNCFgTmGFW
l2Jh9RUy5t/A3GqNv9LQOx0tWpSske09+JyagxCEf8mzymVJg3PakNcFVS5F5rBj
ZYpcHUPvkEuE0vJFTXffNr45G9rcByBbD1ufupmsjPlVlkyQATdQvSg6mevEKdKN
lYOSJ9stHEd3+Kf/V2Gv2ORi0fFFOyZfr91Ia7sMGOZeLqUQ0yVd670iETmv2QOI
d6FC1u46LxC3QlQOaVrdSbwl5TQAfzOY7kjkm7Q7gcCVq0faz3GynptCiYwItobO
T+B7LA5ROPtTur0EuQM/4w0/UARn2yFOzgswI+QE2dS8+ZgxajUqNC5/yoiU/BG3
m3r+89k5Xuz3mpCO2v8lwqecH57+1SaZ90y+D7cfDXG8fx5gBzXM8Bjv5X/ov69n
EgvE0RZ6HcwcQ9czxye9EcOczm+e838EiPAi6m+yiFg4nwxVr95ruMNV9cl9ww73
dRY3fPxpeq1IAKdEXxCJgjMXGgWSJuQ9ViWsX/EfKo43k0y4h5AF2RG0Me6ua2pD
j4pkY43E+jeHwl+IHNmevTqtCMwaSmWSMY+P9JuHsXS2kc/QPxcH7NVXmR8MlhsW
ysr3uu/Tyt0HKYcbAs2NcIYu5YdNjryCLc2SGHqSje50FtTWjHzWIfI0eMCiGP6e
vN6HcQeNYF4ju0PerodEaL4FYciMYhIQJJLLAYg/wO2dRXbP7XGr0OVD4PWnyEnm
6KLjEy9GvuyyyVu/qdl30968NXAKGCn+ZBZceH8Tvn8f6aRlfAEfOiTso4EPMA/e
kaYgn0Hv18K7j2htHQN1DmDzflxiSTEbcuSJqnISxSWtj68kINNj42o+jLJVHZU3
dmhHrCac7+Hu7Tx7rTtMkg1lD1x7J8tbnlQKwB9E8IyTFfWmHXWoCyfHG1upgbED
236+T1rE/1ZgRp7dL3R5kepvMVdWUM9/l9qC4Z4IPPeiy7qmlxq9xaATdQ+yR1QY
fe5c6ELEhLmdPvlvBOviUXD91KCCpUEWL5MIMLbfIgxutjlsznFMsaPYhJFIpAGU
BQOFD2T37NVZMwZzu4WHoy3vmqW8cm69xqQsvXkbrABubwKGpMR8DP9zEUZ8PrHK
rVfRKEHS2s8E/BATdXsy6aqL0Z1LC0t8HsEu1fYTm+91hdfgdtmGcY69Xp+xr8oR
94yfixWCZS7pYHY7QkmaGN6iPr8+VizEwGjP/4WyVLL1Wo59Z3eVKg7FgbD5gxvF
6uiF5e8l+TelqCWDQZa58mb5s7SXF2ki16Ud3k3POGDG+0rwmHutKkZXL7TK+UVI
ualu32xCS8PUPgwVHbiShx9DY4ZUuAWZKve+DQM7eILEp5TVF+MvhAy+VM1m1kaJ
GYC08ODfBTqU+VS3E4HYJut+159j2FME+OBErZdTDBsalQ6t+2zS6EnEA551w5To
BSSvTPuDNzr1Lq7dp/nxU/XfVuolI0kXc+TL5nuISA8RTyQ+7UBOvjU3ruuAEVY0
CfRw2ntxqyK6vSb1GtOOg57BrjYbena2Ho6THHXsw/gbBQSIH9aPfpmhrqxpcW4f
9Zr5gT8Z6UAqgS/8pXVlIKSAzVr7ruIBpneHoRLypXe36uuCyT9It0VIykwepyAd
fo33eTc7TkDpNZr5mpJlL+4EvdUG/fD2rpJD40/C08eWkzVT11+hA6AZWkEzUtxW
nTPbNmxv7ArZIb0/3mm74Ef/SJLf+ZAv173N2K3V11o37+D+RwWTHKZziirZF/JK
JnNbR1L8o5EurILxztsxRTaiTYCo7sHJ7+OcmAhry7HMLGmkXR5aXgRPyqLX+6UF
8HKeIYxd8yZJt5nFw1uGryGyb8AazPHb/mqmz1u5BfnClO7GLRS21r3DhCILrMt7
Pvu/yo8iuzw2VMjUSJD47k4pfbLLRuPETBzbv9Ta2FmsdrIzVFXNRz28MbKm/iBu
ui9bNgPJ0JqQ3os7pvX5jerT7b7fcqGT1NkZSgoCFhFMJjVT4/ikDqY2czCIwCO7
grkfsL9lC5WZd8pewS7f82vExer3DWXQJaWqlih2qHypbXuKVjY5+bHwn9CfSibF
W64R3sWXFSZ3f8h974l6Ju690oxDcZ0E/qaEhrId5Xtc/jDmSzm2GJ4Bnt5tvR4b
KGsbqDcNuSjC0j/nxzrVMS0osWHkrR3TxW21zhJYR//7a9RsJw1lI+L93i23TJ4k
vEApb/fKbZuQF0gSsWVP+k0Q1KdhXg3d3BJaJeAP5bYV1MeEzX0xPTy+oWBWcqE/
/RkCbCPPLAYBuyNEjpZAlap7Jj0bjdmksfTENGvwyymyyMkCOV3n266yi5NTQe7+
+diiIEDF2MnfWyY/5bJ5R0gD24TkGPNlDKjIgA/rXy2c5v0/NZ+ct1m6J4JYHEBI
sunqRXebhjQL4OHWtJNC78vzKv3Ft9B1nQDk2L5oHnYOSipE1MomMwdv+yCqC77s
ajtnaM8nZQvGD4z7l3kKkHO4jBaVpMSryeqzzK8QrPbdnjk+n3XOT6jwkG6drMGb
erglHsrcwThQ5XSQakUbo6LGI0D+yYYZ/NdkfXVmZ9heh3NT1i+BR5aywjHdUvBc
91pTCiaGHKfixvW3QfeyDEuZVxFlasUsHCBk05/yMs50AIoOxxEu1RIqhRyUqyWl
T4hysgV8cEZxALO4CsqnMKIbl5UuicH4jjF/Q/zCq0he5XtUg0YuWGfC6vNNBlUZ
0rNZ3jyuroiB3DWUuKCF07wilTq/g+uiFm8LoFr0AB36Etd61UNtbJkH533uyXyl
u3TWynKTn4eM+OIYnQzTJMd9hJp8YAzHfvrvu8yFM7n7agk1KZ3W/5v+lan6ZAKo
8cs+tjd5lGatZmjGrddpLjGotkW0kULt5jEu/pPDAFp/DpdDIpZwKenBfDaqjW+G
Etkd+7qgbgrSdxK5O+WTjt7jBcLGU+XVhLXALFl5wUw0UUphhc6y+VSv2pa6NjV9
8zDujHCdEslaHYPZJohjKdS4otgWZyCNTGHZG3+cZRnxxnVSRp38YNiQjPJ4/rjP
RjtfblF+B2EdaTr+rQeTyXMxU+Ih5Pu2VbNuhC7vN6euIhTf/HLK/IKGjtFY+Aec
mRPylwFKl4Uyrcj2itYyJj4RtIC3djfmhv83zbAbVXdEmJHUk+0s10Gv9CocUwsG
G6gBruJ/So/4L+GY9BLP8dndWk4+hAqL9dvI+ePj0yFL2/SwSTWn+dYVS45TTBkc
TA2x71tQzKj5aaVrwH7AZHsopJhuMZ2WryL/FVjKuFxYDWIOpQLeOEcwBMAymq8u
epKH1Bgl1XNrebNWcjOIAMz7Kbt01PQJjR7DtGH2Zkact/Tgwo3dC7YaWuqh1R+F
atTKg/NUdlDxAgrtl/4b/9lTdMgcrI1MD1UqZSOQuUnI6D4gevV8QwuLZg6G6FeG
AA1ZcVGBi/AFIDyzkADR83YSxY5ZDFWQkckpll8jZpcnEkv3vHbw1z3QKeiQK65e
ah7YUN5PdpYLMN6i/1h6IWDzn4f0eO0fmeSvt/Qln+SJhCq21ykKP1pe6T+GKGT1
ZRXtY4FvPPoCWoC3bDzKTQyiSM/+3j0Wwj51ao+JxDOKw0Gz4xC2jNM3YUZ1jAeI
SvGb/jjgM15qe3D913V4pQJx0k+9MSz8WM6jiUNPMuRLEYPlRCxAhtS2FV40M5E1
bh+NLWqUWKQZ5x+u8y8ZA0Oa1ZWW2oXgGF0AoFVlm4x9pqr0yKyYl0ctc9DwATP7
DQ426zIVZlECAK483l2/9M1wiNTfTbemDvr/Wg8v0nVHTPMFygLM0rPIIxoTlXaP
Hcknb4i/yLbAfqhb+oDzwnRiWiB2vAl1ids2sf62k4hT28RF9d1XS9TABbCowED6
TKH6hDb43UZhgiDV5dHNQDIF+ekgxxMrxJNyG59yxZl73rjS6cMZVAhr0L7Ui8+C
6PfRojbTzNutrM2C+Y3Wu+9USSbvNdXQEFGTdD2gjjBrb6cyYUM7rL+kQKOulRVD
W08fpXaSvzchAeT0kxgnyLag5jJu3AH7nP3OqjusF9sxHsJsYYNaGvD8lZGSQJaj
QzVwvLNqX8aW6KS3/g0UhoDE3g0rR5CplK+pK/DA1gBiAb7GrLMCrPJks+90ojjv
LVJP0pyu586jX7AhxkMPZq2QhEdLDB/pfuQ9ddTRcDBE4PR9+Ld+ISuNsAXWO7cY
qmTEVk2aBtKruovdciWl8pzK6knOC9avE/jewez+/4JqLBTEez0LsY6DPqDk3GhZ
ORzawRYNQK9CV+XeFbPs4ErvwbSvo/GZrSFHqktfRL7cvsArkQbqSrXygcV5zU/V
vdMcYddWa9vDsEzI4lJhjT/bn3KE/MtZS2WmxKqYsiG0Vd1Cdrqr19od2bTxEOTz
2+0jH81PgH+2uBfo5BevjMgj+Y5atYu+SFJJw7Ay7RD6O74JHWhdk8OoKKyoYf7Q
mJ3wmlM7Boxp/jGChhElriwTgZTFiQkMMh4QN43FyWXxOGZEnjKXCO+l6LNKaIzW
z9XlMDV+JGq8fa9+KQPjsirYnQVC/6kIHys23AsRRUdJY/skGV6m+vZV2LE/R9yh
WuwAXUraRCnlIQySosiGx1AeGOFA3YrXyKbf2KxLpB8CbZzZf91XCs3FAtx8eYtT
oO5YhcVCUr6/wmXaugSuWSfPkfCNZQZV6MSPml+vzFKUlKYR9oXLl/hLM+7t23vA
jpCFqDvomUrU5ze4AKb29xjff5tZbfkL2ucEgVD2PGCXOcbHVgd/seqCS46u3vFx
7Liduf5Fc9++TV+2fTL4+eGBnUqt/x6PHBelWzR6hIXX26AoZsYe/tWJDdLBqWJQ
lH8Biq3s8KgaU9gzPD9J2a/ZR0RdZrB1418OEMuNXZbcc9zLita/9VjAQCD8bd78
VZzJ1GYN/kMnDsjIhFCdos6A4GB1dRflY3KZBgfrzS4wofCSNpLZhjxPB4U6jUzc
ZI+987IXAXaCz5cXsDIFRyaQpEfNuCc6RL2nLux1GlyELag7oLORvEOJtdk+vOVl
GvdRIR+KBozD5VKEzLCatfz11POfvAS7EVb/4Tl1rHTsv+coL9Lm78Rul7SbOFdn
RGl5Sibdsv0W5+p+LLg9gmDskK3Uea4V7SAdYQW06pcZwUzqsVENblHTo5SgwzPl
5H45bHp8oR+mjNI0055Xzc+MGfEH35MNq1bInlJ9AKi+DV6xxzsa6rI41VzJ9aTv
iZW7ruljOx3wrcZQHVOJS2Tm8mZGN8Jhg6GeM2oH6Eav8gqeJeNUuyt37j3AikyA
zGt++FxWhFfH+nrPooJ+oLFo/u32jPzsUbhogrD3gcnS8xRfMKZJcBjS7/ZLpNFH
5Hbm5vR6hGQLQ34+OY32ohrbA32Jq+wXpaFKap6wNTlsgnIexdpOr+5l1imPrroY
gkPW+7ZD067lnrTNmtu1SXypudKh81pTBizu/KuCYpTGqEYesc8eHYZG/5JKNOBI
4DMfzm6qctWTq14LldN/p5UcN+H9Ffa2GAL7CoxIFg6o/3eeLETavnwmw5FUvB7j
Oo415sQBa6WKejWAJdyBGvUY6hD6vSoH3QoYA4JQwDGlUBnqzYEnY1IaD8Z4rOxd
PZDhmtgyBywq9L4QRbyhwP5iInfOEBWmBbnfD2SFGU1g8EqLxguSccKKV212PMvD
SBpAC7fqjKyCghTGQLsYhLsr46yTSovj6UkXFd7nEwixRp31EbhstAbZCk9Wt1Ty
1/HRz43uiBjVI5tMd5ij3hz2UqtQsksZT+Q2RuYyIbzDjcnkrWKFRjGcsYuLAeGZ
DMGOJnTIYH7w2YzMPyHSNtU38fHJAWC8iPz9oUHEf4Cirp5w1dbWB+iZ9yib3jGe
Qir/U6tGuO+uz05nUAEyl7hifed/C22pdhlp1tHFwYiwzfgvFVOXyudqPyB/FZP1
51iGysYhwLJhG5xXDhOH40+502A6JbAKyxoS95iaxZD5IU+xhoOsuYmwP3cmjGol
T3jbbNB18xikS3WcHaNx/a2pa0em6raT8W7/yqI6M5fkKC3uUJ81KxsJA4mPVXOY
ZE21soSHad+oO6MImywcaVRhjyUF2wL5jLvFCndHul07xuapCb/pBhqoEogcy1Sj
A8J74p11ega0+Cm6LppEcW9oacIygqg3VaiKLRr6+patW5IujVwwVA09Vvihyg5z
kYyVMoVTYN6skoQFUqncDsUyPIDlUY5fgihmhqd87i8t10yLsvqC+HFtLdEpMJe2
r51UR6YUmUbvGYTWTIT0yFddD+SzhS4v9iAfzgsqBbVPXuNdNh0CUl4E2dx0qCfT
iBwm2CAOdoUZ+uiCxAGtAhHaa4OnX33stlG1ux1PGIvmMumM2qwDDikeb7YvYwIY
MuuwMLRd6UPWOgcGZ4ljYKKpayDhIARlpcSfn0XNSVvHByM9CL8g6Gq8Jp9+rSTX
uk8n32Q1EPXYVwFaKLspGWcyTO1f5raiLkpzUQwKChJwd3osOT6e1tbpGOB8vD+y
FOjN4le1UnPYBEniFjYX8MmvCXyfS0R1XDyg2NCEUy9QgamuF1LVoVE+BOCgOt3v
cLr1P8XVpY2H1t/igN4A7RMpm4qFic8F1NQbeArzlwZSQq2aWM5cTsV2ViLtktiT
eso5AehNYYVz67u3bZBWsGqXyM+oG/nekhBgmXoLY18TvJIZzTeRbzJh2wRHVXcu
kVzPx2ZpU7nZZqjdlY1jdWjSEtxCzs2sD9kWOIRJ2Z9zx+QtXHkSaayY7rgksTJH
qhpegR3FYNjLUMgjtTP8fk9QUUsuBpdpaEj25Ueasm9O4+O1zIZCyrdO6hlaEJ5f
xeOJKt7X2mXGRKsh7GMsK7BN45qmh3GtCDUt3BKkUGSOAkcE0KktQPuWu8QMvxzP
EFDgHwmV4GzzxW9JV4IFvkfmCGlrgDsTrNM/yXNy6VhdFsIPGSP/bvS2BgRe1+kB
jZKndUJxCbubjVjV3ShuLCJx4x5bC43nqehOAHPGn0Ns0o/Yi7AqUhKU646+9cyy
ORHAJ+g83ybxX4MBO/4Hz5P8Rakud9fNPOqOOtC6pkJTMIxDRqrRTp4SWoAyZ5+J
zZMIbUmWo/wXUDx0vXreLMTSaGXcrlOS43NqLHyjijwkm8IZOieqiXZ3pj2H7grH
jbl4BVqqzEa2zKTnpBRcNBB6x8SHVLl6oFoD7Qyt07iNBa4McGJWdr8u0nzwb0Kj
J0iUai5sNnZK9LFgvJYIKwyobehh3ORhe4wLmtsnRLEXXBCXe1vJ7dEqhLykBzHq
PqyGf8yBbnXQayF9FoVMVnt+OUF4ajZzSKJfHETZgP2DC75lNpRH6WRsI3nugeim
w9LaB/1HKOBtzljlaDtaK0e0xTN+XnsjXjGs05l5V75nxEDL0qsOGvmuAvKWR/sZ
9NeVmKxjayVWOvTU8+C4KFDHXLha/eMiRDcwRcvOCgyOgBbHlOVqtbtS01sKcpGi
ezNjVkphe+qrbRGDa8fuv4iIUtyNeC4oGjULtjaIP9WXdYUl7p0fDNif+ncINkm1
RnFJifaD9w56JieSEKiGjJlc+PKfQHSJcXHJX0Zz/cF1JMWJ192wrb0+TKZUOiWz
y0e8Un0zyZOXgzT0nKII6wCCRgVGOF+jUIJ1DdZ2+xDHZmCqS1cR7LjWGl4Z+6lL
SiE0yBzZLn9vEA5oQ8xbcBmfysPMbkFwZsrbUJQ2J69ITS3ZvfuHiVbIbyIMLdTw
tpuuvs1duMCzdZxzPymdQRKQGAJbJHnYjeFe1fVie1/f5luEvlgyqfMQOT/FvSFW
59CXlTqmoiiA3ZZyrj9GOI9FPiywLzgtjhQ+sChHfyqF83DE3QGAbVR8N9x7iZEN
ruDO72VDlkCamqHmiqMmi/5wO8npZu6Kt/D+n657OcRp9wS07crjDRpAqABkRIcz
Dx5X4fW9kdz4QlNhUrLr69A/wZvcNDPjYdPr7AmVBmrDJFvnEnm9wM8u45Rztp4G
g7BMULcMov/KOUAmmDST35K8+TflxF/XVzrv14Ul+D3i4IKwdrDuEX3YpFBY+WWG
dNFiphfy+syAM1U+Ijk6icYbQka+MwbTd6oz9QFr4Y35+kt4k+HUnw2xw/YSl9M7
mTh++YRlAh3Ojv1Nafzrb4P3KqsARPcUkBDsNR2UTag7vuTcZe2ymJMxUP5A+ZOS
0ZoY0KMgQuqrqdAF6iqj0PJfsimKD/fSGMtWWqoE75zFKXQck0J1xoJhgywvddS2
gBWwg1L0qwGrar5bYPpvTC2DAsStUuUcZqvbsbxeNbCqJ0MYDa7dCRgH8yl8fHgs
/fYudYp9aMzSPRNt1y7FmSX1cO+qcjso9IPJDm1nLaBsl4Py7sUrdOd8E1hRuYf7
HMNFkJoL600feZigdAQvsye/uWnIl+H16qXE3X8hyC/s17ZR/b67yWeHKiI4K6HA
hVCx98cXsHlu6EdMLbmFCiJMUn8TQZuraiPkzyfY2yJ+wZk3kG2079saUZHmWwEa
W7yo6GMYWr+Vw7uRrN8KXxic2IpPD0zxkXIFweKDxioa47ZdjQy7RJzPjYAy5HnJ
zWiH7hj4WAbLxQOneYg7gU8PmSmzzRk8clGNFBzIbANdxsAkYj4SKiGWQ1hAytKn
XhlRDte15nBiIOenql83IpAg6K0j98rUCx9JsDWR17YX/gTzrYI/rmK0j274NiR0
3867GoqOcHBJh9iDOt70D23DeRaWUaK+WpdUY5Ozo+CoBw+Dpllfj7Thizj6bC2P
dG2/9iMHl00UXLIaCzBb1fgTV31Mxnbp6A83FdInSCC9ODwa5iLJX6XUeJjqp8dF
SKgp0F6e/TBr4umglxdTv+cyfTre/21eW68Rc3ayJZnHbdp+BKw3XDOh+gGxAtud
6ZvBYub8IUCL9a8WnLadIefgTaLFc0+KIt7OMhLWuAiAAP5YHqJMQVRUaKbD10pi
O7gJPR6cyoyV77c0HzsBQkYf9tCQ2Df21nabeXAVZj4ml1FrZify4WNENvDiuV1A
Dt7vScMsJ0zDe95q5JfD4/uwa2K+IdskGyZXf9vM8lkTl0xHZ62u84S2k4eopu7U
rw8COiiRFRWR7G0oY9Mo9DSbXjyDhZX7iGRb4syULWRGahFgu9jzNHPp+xpPmbiy
XXy/Gbemu7pjKygZ5N9U8V5r7ItVwzhv6k/fGEyyP7DmIFSLhZgtImlNxeIV63zu
XDs2I+8xJcS+my+KQnHE8UCTDnFRsL5ucVpnXP6nvmyEatUPj2ap5SlxW4YbOSEQ
uQ365X31rjDGFOm1UFZIlUJ3UOJdIlS7Gr/z/FsDNNkEIkMFFfi7W9a8ui/HuQBu
MPKhxdHTcJVc6+bgzVaFgpayinbgah4Nk5hCMEUb//8cCNWhNd9Xhj3TIN81ScvP
zp+LW0hj/aVM13vAgdxama+IQACWuI2Mh5WFKSHgwy9J7fpC/Org0PGaseR8KhZh
KMuv/5k44kO5WZjVso2bEZkQ8cG/SEUhHeFVDmS5iHMymx63HZX7RLqP2EoSfxV3
s+BpE3LS6qbqh24SrKvp1hbyQm1zhsZX9zmh4BjejtsVbZYfNLP3q/NU69dghtAh
TR2e/aTD5BL0tVag8D3bT480KBagpY8YlYz4DvKf4/5qS04e/r27PI8Bs1H5I1xE
GoMiGgr0pvTYl45R0iuDZuc/IkBh07B1n/SG7NWAMPdTMJzjs7z1rQHVnSo+cK/1
J3Tkf0S354p2QPMBongwa5M8dw5FiGQrRIDXAeKnqqbauLfJcEph35mVETE8AIC8
jmEWEoyN3Js3n/HF43Cc/IDaKAU4mbSsf2XMHKwit7hQOW0HD0QmHEEXMJmEgNeX
Re8L8NMOnJDJVke407MSzI8vCvrcS18FyQXWC4JQZLjJMbdKDe5WpfWB++CmWFKS
+Sy8UU/2PsSWyzaOFVy1s8gV4PEMBlbqLTGl30ay8w7MAHT0v8sL7pQfkCRaza1u
quKxVyp2g9VeLBrYJoIzehm3DAF0SmWG6mqXXAn4gURTap4oyTLcVrJ8dThXFigS
GBW5EMfDv5n8vCUduV2016+R2BR+AET56bDJJaUVpjy+bDMJlQPK1HQ5U3UjUQIT
DcgQ24SCXNKIOut0lxFMqG9oGGTnj4cIIRlem9eudU0UNQ8L1xubow32p6o4G3UX
a8BjUqVKT0dp9RMTaPFPmZ6xsRTSo1a4czTJtAkPjeJhK741exgJ2/qFqJf39THz
k7xXt0w0gdZVY25ZDquwl7mQC5KRH6oslqHbXrOk8aOgKNGF9rJuQ9bEGNjnaI0N
DpOGS8MvLVk6JYwjQ9aPACF81u3DaNH+Z1LloZcciWE+HUmBmvg6ubTOoJEw1dam
W/W3SmXc6L1by9d68cdWDv+U3vZ0HjXRJd/rb4SHWNdPGWTnd9scwQFUYJb5EyuI
EXJkYYh7PqIfDpCXj8x3p1tiHEWIoO2C0jbDZjDDEORhX7W/hEUIs0rRfm8+m7oD
yT9Ycipdx+vwBhQrsQRB5HhC38R77DQM2L5k9PhTXdpO+hQyjzKxmVYU/TIdKeqF
jXKKKCm7/skptb0ctcRDb9nC411JX3bBhlsrrtTibUwy3O40pLku4tjkm/c6NFzj
/Fgekh/VQL0Y3Ns9Fx2wDRS83AECq3SeA0OONuNm4uUQyRsbMohuB8OX4nknJJ0j
xVnyL2mOddX+xveIU/YN+oqqMdDl0BWbsNZJehjdqgiKXvUZx3fFMLQqSDuUYwPU
LILuwrrOfOJuXPHMNZWznOM5+m5hBrgJdZde5FT80wouCPl3ahQHZcDhGbNEVkVY
dgIkvV1jPMg0n+cdI/oKlcggN7O9KC9aoEzQSxmwR2cMNPMyenfgjWBpb6OAWOjJ
TjNSTTuhmiKyhnItlikkOMU/50zTC8d/YlupQyhggoJC8Q3kiBg+iHOynU3NqZ1w
t83t/+0unRaJzyYaIJtrNIFAq+CeJHeq0/cUemO3/Murk1wQAgVsQj27U1/Y0EI2
6KsSP/PMtKxtuEoY3lxAdKPf22wSQ0HMHdsjs57GY2NIsepVOFYQtahPrJH7M4u2
Nm1F+dXF3iXPWvWYILjhldmS9Ix7AztwOxNI9D8xMZ/cbX969V6oFGuyjG1Psvma
+VNaMf/MX51/V/OMMhT2zdmhRMleOE+4l064+M5laejG3uN09jmcC/3f5C1VMAJ8
stpZHEVrBQU5/G+YQ+FsUFPgxcZ1h6RvaEFe1d2iquVgBjUIiZVotrs6E0Z/hUGy
/acHB3IQZjF9EbpfwZYhb5fkYEDpwz0eZ/QTkFRxCanfJpwOvqoRSXjfBrHzh3LH
ZAaENOiYVOOPOiXShN4DrAS1Vucz2E4puYrT+ucmz/9s5vbkM9JTaZvWLLTBOmnx
JmkoJ/RUHTFD7Iql0Cfnyxbal5T1TzAwZIX2pNINntAqkWlSiX7lGbROFGR56o3x
36dSIMsxH21+UZazysMwZAmJWe1CLfFd/rjb2H+wEP3Gk11DicfUDNVU2XscsDOc
5h4wSD7lWkUgkR5BlhYixGdAOjNcUFBZ7EmyTtpudg69FDGbNdEOME0us+58p5O6
17CUZLmfEPk1gVNexHsIlaok5AWzJbj34fdgQZLzInmDFGNvfMkRjR8mDRVsiaaT
03O6tv/d+dmkAPPBBOjXyNWtMmIo+ycuFPN4omQZo/Y6Fgna2qykXnSbA0Kq3czt
H3SgZ7Y/B/tgxJ6QiSnr3qgKjnxZ+RMGnR34wEZunr0Re4BgOexnvQMrBzhMaONK
iLOxB0q2FXivpTIzf0mFpnvhEDXF0mEZ2KKm1jthBR9BYLIXanu642DrGpf0Z2FX
So2MOPLd6XG3LoBkD4xpjRsAGuVfK1MzK6h2waBpadsWhC4oje5Zi3uUYB4FhvtJ
p4PXEEPfdMzpsOl4BJ+P2LqhzA4kRqjNXGwX4o6RXV9YrSefPgiHKrwWeM+Jl8c9
VaTt+KdeLlAQoVqwrAWAs0uaDDoDsekUtJkGgGigazliaACpW4NyJalyDH+JPZHw
1CS6o4r1AaezRZ3iXqzw049wyPgvnruVz73PT695RlzB5LRTIir3LFHm9JpCnLx7
Yo0mD4NFkAgtcN0LVkO0bTn2n6m6qDMKzWdJg+/2cW0/9+2UhbBzsgqvHd9V6L1e
29SKWo8z3HasU+g5j8hMolT431vE5ZFnUgt2A3HxI/WTkg8+TClJgozMdkrKmEW8
UC/Ss5W0zJd8AdO02vzbAH+a32OashQ4m4Gu3BtER88526JCmcEK/bBzkmKY85fa
EN+a6HmXR2V5LZX1SALsEmUesSw9id3XCzj2GS6bBBzTz+OO0xyYufDPWcY1yLvs
2GW5iOq+pADvBzy9sFaVMnXCtfjvEmntK1bRWsjAVhAUtUFGIS8PP7C7jz3dGWjb
ciiWtpGH3W1PBZF7S51ISRa8Wh9OV197NiFE4rKpg20DJFh3j/8gFIR1Fzasn89i
oIdmUjqJZToLHQv8GToSOQdj80I1pBG1i8PPpOiQGo+DtFsHDmA7hj3KejEb8hzQ
drwJmDrWVfOOmgkA/CoeY43n7R07dtmVdxTlR+ggFe4xfaVc+oP+x8+KcdTt2hhJ
7m9q9zED6kj6T/hVD+XXI1+X+ZuW90ZNBXdBojmvrvl3lgwpBAo+eTr4DrCB5nHT
BHQdM+cBQaI6v8EZL2x42T23uSd11+XXGi9Tf2u0HL5+5ZsV7W8mISRBb1IL9VyY
JOmlqfyM2cEC4dRgNTvGYx3Vt7k5iksSAepsUM672ihU47WYCwbwRNqM31qSpaqb
Im3OucLj4j+3W8mCmfOvWvrTtMJvicKcdlZErFUxp6z01KrYPaM7S1U2rUsoRW3y
pFFM/ALZya7ABM5BHBUm3QYF2l/CHIWWbmHcKiYRqQHd4DfPZNko9rvR9+nAta3z
ujN0kqafwiSdHolManWq30rdsEaImm/inoNutVnThsps20F2ixGoYUqfIDh6yS9+
yc3hc9l4+kPWcIHIdFeOnankfsE5SyqlgJDMPbKrhxi183QSCo3yHwJnO6FdiugY
/kQWDo3iI3NGjQ2UdLE7DAsTBVrgomvcmWgKVHC4vUFV6WDyObVzR14/PqdHykkA
bOjnOf53nIRMLmRFuq4LkGLgisYi80XBKfGByGk3DRcB+iraBu0+yZ1WViKlcJDc
TMeQJRuAs7/zo1zxygd/vbsiVFpKYK6bzErtVKLbi+Qshusms8WCymMjF90BKWPI
WAU66oq0vg9ZwPRHfgbSApMSel0g54l862vrKzOw5Q6sJpcM7jFJ7J08hDLfHRLO
IYfwZTYVyf8AMs2DiCU9IQQRCpoJ+jl1CIDo6qWlzegrIZVAbXddgo9Tfx1Zj24P
5xKGBHv3nWKoDYAqaBLyMkoKpo3OdwwdSEdraUhjVYjfBFlzPsvzjG4N0yrj9Xz/
24+fynRLK9DE/YeTSJuK50EdYq+iXja9D2Jcqqg1HG1nTtAooFi9L/gFZuXn0Svf
Y/rwu+dbtE8UtJAVSTu9dHmw8jUDbC767ygyNKelw+rLaCgg33avNdk2/SZ8EurA
L2SAcbZJReYyqTmHFRHygC5SHftY13iQuTfNrIX9VEZrKZ7b0v7a1TEigtuPkW0b
qsE/Q07Ra8/Mjh8j/czWe6k1h01NuOpQSRP2JdCJBAmyhzWlidZ8KeMqssJU1lRD
3KhIPoGnabHhrv3QkNWRos0GxYxHtvHVOWGPFxBAa9xlHzEglMSuIDdb0QALFrO2
IUjMAiEF/tkqKd56FSNZrM4fhbWcgs3AiaSdJkGIAQzYw4c4ReqoHshSK4pPhykI
ZPh2OKWfJJKHFIth7NaDPbikknm6MYITwd6JEh2wOsrVd2oV/dnty00m2lHiWhSA
9aJEsqC54IxT0dznRbwYdnngM8itRwNjRRU9yAFSDrEICmnzEAwaukSqscCu4bk2
VRIFeda2u4pkb/apdsZcLGnugB1rZ237l0FM2YjDylf1ezzTJRJ1z6OwZC+2ey1T
GinWimBExtZQxwkomIjDQKOWBLaXS5JmWVlX1Qtr2mWzu7YEBpqNWujtfE2tqG37
oUh8A0fyypzvMvNuyhIVJOaAou+qOkW0A3EbXcDvYxQwlEtjHGfa9jtbLyDvqSBN
LM/lEnjAPV5WEcnauxhNgVkqKoc4oQGG2NkbC07UJzxjKCbM9kO7R/131EyFAHWT
HN9eT3meakJRsZmKsnGVVRH8Gv+NO7jjSKSM8alLzpH1LBDpqUwVa6o3nBIk4AzP
9Edbb4nvb2z2HL6FU7r3Ttjb69tzo81VCX21P1oPH/+UZxs8f2zCVRmTDvR14FP/
fI6FgLnBVrwCQWcFk8NHWrAnRcxI8I3fFhcBO7Jwc1lbp1VCpnAwAt/7GZ4ZQ8/g
nirFKmdmVO8lSC+FpVf590fQI6nx3htZ9JPGVE9wgxGYOqItZZc+DSFK93r9ZOUQ
LNCjTK8WMAmZ4qUzv92xg9kmv/h/IQJmS8XkpxtHobA1U/Qmpz3uEvOvbp4ltv7z
3Ya2NASUdCJHuKnHitwjflHhdlYmeoPjuSyq1s9W5GoOz9C/RdvwKApODO7+lwqS
wl/u/7eCE5Zjr6MgYUlDTw7SD81vVXJucTikGP4Z34wIcP9Hr2jjQgEQgtIeXN7g
C0ffTBto4UYq6cOzmjo+heNm1b6n2OL5EIWIIgwz+i/MNyeW+fmcGdiWWeQvOR3x
kKUjo5lzwBD1NwF+SlzFQc5s0mShD1UU2qZfpbdhlEwsq31UandZdSvMjQlVay4p
hOqszrOvifaRBuV3UkUE/ztWOkJsucaE9HmeVtm2mmGMAzJmwiZDZBnjOdBr9Rgb
uI8VsxrVXuBhtKVtRF+Y7ocuxG9xvbyD2MFjxPGJ/8BQ2Ses9KDJJRsGyBVjGVsl
GjvytGVKZqtDvAxZtCP/CrpBsYJ0xA1mp6vEGvnsGmnGMju6Yz9+XR8B9Aef14j2
dFTHchDcCZti7q5vW/mdZV1D9DwyvXMUmPdU8KVVaG20pEBFZAltEunv9oVH470H
DIHtLeS9zDaB+GGI1OTBRiLqlkNUkonrOnlwlEMG7eYifA2eaVZkawmk6N2yJF+9
MAg7aeZhNrDYuNsM63iibTqcZT3f6tM6QxvR7JG4/esR2auY/pne5PB+Tyq5f59G
Q7Mg/T+kfOF8j1gyGyM8KWpBkhKbP2X2kvLoXTOkm2ykdy+aflidNFy2swhuNAlO
SXJ21iOHK7Knv+PhXcpAiZwwxfqY+6cgj+a/3d6sbIhkKrHmQHeQGUNvHXH0tK56
ShKUEcszYTRZrIcm4WAc+fXwI8SG3yWcqc7omzD3AZY=
//pragma protect end_data_block
//pragma protect digest_block
GCLAdisbshQVG8Zg9wdMWwGFp/w=
//pragma protect end_digest_block
//pragma protect end_protected
