// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
DP8RPv0u7sdDclYCTivglr4pRfvuLCML5Z8yxVIuYufKW9Vjd6x/3FFLI9Tfgmkv/HhYcZMZBBer
epD3C045Ijb/Kzja2CkNP6hBNSymFnoQvVZiTa7txaV08anBq2lMGdbc/YsmZfJj33h1ZEzWUHSZ
wYs3redZmJk/Co/CBphJhSjpdhNycfzziIjDLj5IHqgPtNoeZPKj69NemzSpjigY0O82VaHnw7On
+nqYKPsUlkmifB/q7v+rhywPKpgGMvJ5Efs8u5YPDPO1unsortQoFbGcGE+Oe1VjTXdc0NKUS5lM
P2ut3m7/MOVmvGnUO3kG7UQOm4bD4cbsOJQ1LA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 8496)
zYkcBTpuIOFyuL5Qzb+zzWmLu8Tg3d+hUBBe845kb1FNRQLCjwIkqO2dyt0qj8Upl1XYs1yRo4LV
Xu7hJuHNSds40KL7s5Od6JCv2ibJXG/h8rSy/xu1+ECJAwSHCmi3HLKTknR62O3VSkQ7hp55Cr/h
1c4G47O1z467WDdGulqR4aw4IxesXXX3BnepTpRYoiTwB10DCFa2D2NkmP1aNBmqFvcp/lNStKvL
NiXJTZKqyhcM9pQ67bjXHlOKGBQbk7uJJPSXaYzFUe2d2Zf6Y1Wcqc+3aGRJWFfsGEChm+Mm5Nnf
yQlEoBtcqojeJv2McTtefTN17bJPdWRLSJN8Ag2InTKoiOrnMQSZmbQ79nhxzSp/VwXxakezRbZa
1NnX20sfyC/MHz7kswP6Cafc6LlfNWUaEcMtbst69e8KhLY7e9o2zewSKhTw6490OR5QvKBulGDv
+NBNSBgJaeARJ3x5E6uzdy1JqpoNNhkcOewbhuca1qNUfYfLdP3ir2rOCiAxgIminL2wDyVqPllQ
QH7UmICl3RBfnB722aQrbr3+xwQy8NALTrXggLkzuHB+JygQvbynMBTgTiZO5xQ8DqohpbM5ib8V
XnreDzIe0YS6X0LFEmuO9RIPEK1JzGcba91NQoUTO+ehEubvwTq5TyARJ8O7BnAHIDq9x0KYz/yN
abomVbUaKgQCdIOIuPed3sBEXz/utYJg56ez9wLZMGAnaYdEZtmOhx4qX+zS6pYlQKlnMC24xUla
4uS4Lkm7yyFyESWPxVaTLEdN/LZPzlZBZHQbq+yU/Fb4Vr3SjeNrdbzQwygRZllV1XSqJ6bfBcCK
GmZQiXLDzISWU0XZE/6tAK+YKsioCwrRj+rQioO7/8NE2WOIAVaKhS4V3jQTmplEi3XB4LOsZi8u
6Fr8g/tF6GZSVfWtCGB7kaIw27dLh3k8bLv5XZSN7Fqm+jiMCjyL0VGxvNBNZoXssr2Q6WCJy7gN
T3W8Rm4RQOcHyJid2kSx58Kw1k7o6kxaDq5/krS8IWMIDBeOC1jCZlCa1NdqfgfsuCAyvp8yLRBT
yq/mZxD00kRlExsaPHiQoy2CVInrs81aoAxAempr+/MYOZdkKgxwLohwN4emA0I/gBXJa5AwW+BK
guydcmmlrGuLv2i4vChqgJTDDq2/jzuGQGvNoW8b5ooKK5g009YD2/Y6u5UV9kEwXUsjaUXFq0GP
8zil6hVQrmtVzDAAUr49wytOsrixgODTEswjQx4ZX1Oq/XiWXHTtvduNPpBYW/uG18p/F9p3NIr0
0hFA+wiF4/DcMWcPMW+mAGFs//Y6mwEyFzoVWSWfnqauqppsjbuXvufo3t/FXynOPM5qqRGdf+c2
DUmgMOgjdvZ+J+1aq+mBqfvhhGMPHsubRmhez3lCjdoW2OS+tI2IGf5ccGIWzkm8uuYAgybRW2HD
acNaOrWo174QjYF4vth79cXXJSMMYAZoMZHCa+GHVtmDY+POYJmASIFN8/44JkmJnF5K5MasOBEp
TUOwk8UZav3ic/8OAi79fxcNDr+nP3PNLvcbFmtWxmZP165oOJBbCKeitPyglBu9V97wRz302iza
eX0AfL0JEoXrqcCTHF8RdyWSWpNWNcTte6uf4oZfHcCMhWIyrJEq5hqtqVTgDPBuGImKU8Oh2NKs
IukuKbod/RJRtJrkDmVInOVzLW8rb634iAO+Xb7k7eyJEX6haMaKipKvvaOvOJk5mbpEzQXmkrgi
fR/ALMoYADCjyqmbNNewTlPKNejUf8WCyd1HpAr7CIEbRzmjR7YfkiyYsGHMZFOiIyx1EcuxKuLu
T4/Zvqy3jnVQZxFFeCsvANyLhv54IxbGqEDDss05cdIi0ppa7Hu0EZM3b1dvtPrRTT+xAoDZPTgd
Nbo7CFMIRVj76sIEiwYwwkU7QAQl41KCSyuEiqVeH+TdMbAo9W9aq0FX8MCcIF6CO3EVTkDtK2DX
ZnjUyp2HAZkbSjvOH8XGUY+jYZhvIi2Y5ehBGjZx5fHj6hWUONYn18nLM5DsR/vPCmOfrNj5UU4s
0Z8uNRk4QANVOUttj4JjLJTZaULrDMKafOQblUOH3dJONfOQsi7Iry97OnfxEdesgOiuNBZiS5PK
elwiWPEdUq4CW1fPTEn6yE3wWDjn1lzJztOjRXeydoXeFxy+ufwyuVG+yRCzKvhRiwHp7br0ARe/
oVp6iBh/JOBhafwRlwNXN4jev8MFKxSpC332IOZ/ADrTpxsUAgJ/sYcufXMpUWN5PEj429Fg8+o+
fMdxMiTYD8I8J3e1EKezbvTJ8jUTjuuV/KL9vhTc5FRyyn/zv7UOiUaBZKztPotuyCsUfOMDIKER
YW3GG6UCT3BAoB+2nfVrMSeG9cX5qkndyEtXMwbyZ1rBfgD3fp7JcoP/EGVoTIV6Et7rQLPCzvcg
wZh5wXQ+D87WGGMhA6sVIN65VAr4awz8eoExVJCKHq4IX1Lg1Plht+GDI6FNVxvap0OEBuBJYFaY
7oOm+hVZOWvI8qnqclYaN+1pkMN5ruF2KIDaqIHPBrlGjmgzPXv4UIp/CXx+DpKBKTukPg0oQjeU
fiKznTk+PCqY1esu4liyu16FaN0YUxy8dzriT7En7q8EbanzmH7r8y9gGqz0DBbrZo/0htyFgq2h
6rZ/2EpIGQ9lIilkUuE5iNxWG7NIt9Hh7E1QVw1hC/I5a89kiLQ4mu1Rg5w3XNzKrn0KhAK1xu35
qgcn/3h7ZJrkn6aOCmBELEjyf3qGse2g9Z1mPgvBwlsr4r8ol7ThRg4qhiCJ13A2neEpQ/DixoDP
MkDs4E/DUY6cQmjsH3plzmoPN97tk24FOYITTTX0TgOdAO+j2VFIN2vVSMMaaWxj4PlYb5DAAZaI
v9OX066pN40Y7Sc4bk7I2gnk6o0AYzWywADoPgk3wPpbNuRbLTAx9K8irTaIMRi1vmmleq2VXL9W
oWvQr92Oc74WTLbhyDyrxvu1fHWArpvrUvq3B7VTh8OKAjk2L8XCDSu1YkojJEiaTYk9/0phkUHI
hzC8nld0ETi6doLIl9drMwTntFULipDlTzKDMWNaDFFnttWSYPlNUkiJP58FcZyqUeULNQK8Q0s/
ayJx1nr39+Z1TT+wERSFK4dJ24mDOJ1HHKavOmFAZFtk/5rhTcVnXQBcYCq+8ehtwMHWQ4DZ8e2f
2kqJTSeS6fr69SpkKakYKn+UpKElwnG2nL3pKI1ndmYzDAOBqsVzVekjdYYDcN+4kGPR/ETWhg5x
SqmDLEZjKVkm2vRCnrlcAj5R+RDiU/dxk9Jilz/qWKYGoaKRwW+BaQvAO+RqilJ/CDStaQD6mgyk
ZOvnoj6VvPxr5MWB8NgVr3o1S62rheW2A+qAD2A2U8W12wc0vxi7z/ylt8QShIxAqBrVY7u1mzl4
hrzJDXkF8kKQORJB1q0SE88l+68+M1y6w14shjK2kOUIPl5KBo+aIWSsYl8L1Kp+44l8vQ6sJxux
Zv4WHmyH/f8AUg8EB/HA72OPqLXMWYoqHVCtTGFvlZkLjGFaiRdJ60DW6svm/N05S6IL0Fx+5XO1
eM8b/e7BxKaRVFtcFB8kazVP14LTEEwHbyhFOgPtnMWUs+AXBwLBNIf35q/GSd0p/JR9dLWPp2fL
nfuLPxqeX3pvx9cBvlcwhuCbgeCju6TxCoIxdRadOWg2qxtvlDBoyOZaK97a7xz73pSsI3+d8yr0
Wzj/XSthZGEyb2OYLLsrKe73k8WGrgRKluxMHpOhlaQ+gKU0ahjdBA7hkFZzoJiU2L4NfvrFhX7q
+7uFWqMfhjCe3Sphatc+UU3pWhqVfWdpFgQYpPUGDmmjDoU7PHU7sGJ2RBcOuvLnnBxyIHYHhsIK
yMIvIqNuYsaUb67d+8PjNTor1SGO6Y2WTFxk+zrsKDiVl78SlUi9IySnlnvqf85idr14vPLqOVYz
KqjAPLI8j7DYn9B/66+Ok4BVegVsMJHd+wuHyop6ivkFWjelwk4283+r2/vS9hJYPUvLoF3cGf7b
/5fnyEJnWGmhp72yU3qBb/llhTCVKGuf5N/6bsZbOpcIYBycNDadbONobxlyhI9rlg4pUbjaFOTN
SQxE1ty9PhUdLk5F/zw2Y9Ke2fYp9KMloquTG++Bd+GqKvQFip97MgOvDAwqfIak5z5eHbhwG6tV
moozDqpnyn6B+3+j0qQkjzeNWafStfXZSwD2+tlPdVPLXFTms6U+zB+Droj6gRfD6IquD/Asjiom
4Dl8QSrwBkr7Gl0IwnfzeyhyitzsDfRoO6JGsjPWOSIgFyFH1NLJ1R+ozHdE90jpls/+S1wUY3w1
FlEkIuV9dbv6pnnUgdrg6VHvKC02coSWsR7MVUeugR5nXY38XDAvNUqxluETERBMzFvPrZ00PjSr
98HZYLyUeEAbqRlFP6XkE1nYvl+fbydO4QPc6MGgUQxlCeFEkLkD8X5pqpZcxqpqnEJ/IYxaoZv2
sRiI1ySY/9IkXkXMyRRHs5sAMHhyIES9DgbUwN7DeuFx9ycxWTV6vGUuOYSWNP2vPuARK+nKDSC2
WHgckOpBSuCiolN5XQoNsJHoC6IEGL5ON3Tj3IQlgqPbqsiaSh5lcYu0QzxddBQJpHCTVqoRlKh/
VIQ8pTGmRRzXzjeuBogFIU6a/gBm0oVVChfY2CWdUvD26/DU50qBxOK0fUjVp4y8cxJ/Mm3GVye7
95vOEkx4PLr3yImU4xKh1APl2yeXcA49B3ibSuY3E+Nc/0D2RbTfopUi/peF7jLDJE4EW/XiT/mG
kdYpT2jXy6gjqPKg9iIoh2U4e+heHMwDSisA8tzMZPerShup31B8GmjxeWq2SZi+9Fa9NmiUA8vv
t00FuNCiKg2Hy4dXqT3UYk1GY84Vh4LHGsOmuKdFxSoh9rX9wVvg5a/VDR+RKPwcFaVEoLqxhQ8/
N4NAJ/ZJrVyou+7t7YTmLI3//HLxOog6fWO0FDWxFu8TLDvpCzbnznIx7tBUcroTz1PGpwVK6+Ry
hLnxJFQL0vWpUqmvaMeF/ZMB9BTsT8gkNR7L5qp9IkOKCCM0iZPLtZCSI84GEkAAmwhVUFRVnKdr
KC9xyJLSbFysVlJ6GJcS7KPLVA8VpqOZgo3fwBhVg/SMNG2dfq0Soka3y3S1s6/mcP4BuaHOgmGQ
kT+cAH2jTjO5kJDUW6kBkOE01cLVj1BwhGWaNCvKpLSk+bWUji5+umaNekIpsk3s1A6ULRcsR1Ht
YQqQOjGLjrSCt4yYpYdDJhSx0BnKrBzsmRGyWPJKaFZja7CSrWFg9PTwkqYKvsloLUEFY8lPsM7K
uTqlOalJmm2wTgjmJHkjJhGTzgRpYg703lZ2/PLbD+jF4dRtlrIhh+66zjodkbffvzzZsum5OVqs
JXCCcPkupnbU3U8WUKpG0rS0wCVUdGCtpfVJwjvZ5WXpFy9q4YmLKbHLHsNfBLiWvOhk4tUiAbin
yXLaZJ+ghrA7la8648tmjJpTyXFxulpGTvMPogTbEMKH5nRsUat4k73Ajj9XyjBwkUB8Qn60LOHl
2sqgXsdITuQ13/flSW7M3NdnrCpi2eA7+1JBJnBqqz3dHSKA/2eW9cIvbPLlIuC1C9VWuilI+dpZ
8O9YpIz98599F1xSEUrzbStrzLADevpXS/kC+ZJfK2bc4MsSJ8aslWkva/svTt8q4j/atDXb5PUF
TVwBEUUxISz5qyWANcA4fvS/vnzSPvWDSUejNBdlaEJB9f+Jo5Mxz2CWWSA9ZiZJi/5jfL9wc39z
mQaMYIdVoyk6Yk6igodLaDuCW3LTghMmjoueqP4syx2HbEAmOBtwHntIt57f1sVn8tXLiQcWjGfu
FRy2tvPHadmJ0uYSFoPEkLk9EX1FWRvQW6E0TVdvI9KaU1ZXA6pfvajbLQguHs3wAj6chK5+o7n4
LoS4cj0o+tJKj87r9mGzN0DxsuygK4FQQJPLpKR17l9EnJcM+q3BUMVWW8v1B4Dw9tCDAR/bJMgz
x2aV6rIOG5dpVtd6wsN+mnws1wJx9IEiV/MyBufBjomU2XY5iwekDUHuFik2+pPJ6HRvWApgEB6M
G2kbfT4MQOO5/4eDLpSveHpxvpgfLEOfmF2/0ShQ/K4fM2TG7aOWBJr2KQf7IX7dI83m++HoohEL
+n5IIRqkEQlHOjUp/+Atxw7TFZIPUXv8lqzImlnAbrGYHvRUiHtxDRv9Dx3fVpKtF1XCUGrgfoDt
BoN1FFTXK/6Xc1bHipn5Qa4uiBycsdwmng1MNfETIRHdo73IduLbqNJnJR0g7q9iYrVdTxxB2/+O
KOq2CqO8xHw2B6/yVnkZqtMSv+9mPk+QWNsnMoHnfkZ6qooWVfLof2D5H85VebKv1YgrT60Azt8N
AR4cms8Wdjoq5R5ZbBvLj6ebjsxwD7eFSfLDW4y5FpYJdMF8CuXfrujF4ounkAaIQ2Ls35G+lZgL
3txaPxqoOusYgb9kM4GZag8MemYYem8iE5VBJGJraIGQCH3zmsO9DVMni11o1EV5bgWkBwws9lAY
+vKDqF0L0CiYG3sAmmESsrEH2lMdal9ct49xaAHhNw1Ziekr3uYAge6LDCJehJNxAmCAzDiTLJM5
sw7DPzvmWqvI9yGXMTPfWkUXOjvnmb0uUTFoEaL9irN6xQVa3+ayDXU8cigTseMT8P94uVWahIf3
Yoo0Dg8E669ea+eAbFivqTOhurRdmGX0VfE0ZI7dpk2LSQypVhfmfSDrqzwVFmlQ8QKpVsq1SIWX
/7AqG3Scni3uqiCImy2SMXcGZqYGHR4scNBDN8h6ZHtx1JG+LYD2czBNZgxyFAbpGulVKX3H8uwz
lExe+91rO6wf3oA3kVb5hFq0amaOcKW36F6fiJY06ll2ctwoIx8z8KXso/keexusveKaqlKazFf3
84KlC6EZlOFWWi3HpHCQi93FlZdgi76x6MhqKZ46+XxQqtzzh7rrZxbDhXa53gVZTOrDGabfTAE+
TagX4VrJmRhl/SEuWJKPSy9bx13cJrc3EpdwVEBgYjUhi0XKOG4YMnAGEhC9arI0hZCyoOyuWWLB
U6V+f+g2zX1O9riOyZwK0/xNKlUMMFL4ca0dFITID9f26MAlhXiOaAa38jzbzVZbP8D32D/2FR4R
eAfMjU01UJF0EyuQGySJD1Oo5O3t8RE9M7CCuyyJ4pHLVwrOliTt9eFE7BdsivF8Uc068lz7uA5d
ECKvmFPKVTy1tsJy+wQY7fljZhR5PFGig/5XgDNVi5lOouFaeIgZOoheX/whJ0uHY/62TsLzpYdg
SqwgpekOpNTcBODlJc2X0ONfe8UUzy7p9j30LgZQjkZg1kQM+8mkcjHzOxMkf57UeiFwJ6w/vfwq
1AZnu0ZNytoFSEt5nB/CR+t1EtEuauGvdQMCyalmNS3D6nJe91VYSu2SkGFzpl7/U1w6RdrI3cJn
WYO7qLVo0K5ik0hazUaKZycL4HfDtTTxnydvLYuTHg07KD8WAuwIO402ynwD/9w3XiO835iuH5Ny
8oGwemK6jbVE5+XWD6Z+/isVqGokXGqZcxf6m680hiOwF4qOYPviY1NaSlr/aoD193ne2UsNl+sO
hR90P8uWMMEr+fxz9VnRWql/0F0oPj7jeDOMM6UyVAjFHcLQ0hnyKUtIVMChoKbhZCr0/9g91kR0
4c6+M/Kx/H81t6iPidl3dWqDENf+56zMHnYqeESDYx/wzXxd1IFdPkENpHRY6+lLru+h2YIfy/YV
D3cFgEneZyWrKRJvvvIxbHH/9hTccPKrSkUmaSfLeA0We1C4JIEuf/N3s+j/hOvcx0hcfd7SbmRu
FF4XMcGmfEnrx+0z8AutYW5U3NsqKgCF8H6bTTzO5fpcfOoUX0/1m5GFo5GreelnARoz/tOB9+Zh
349o9nRegdqaqR1dq9W16ZfuwbCBXrOUtpioEL5pFCrDa1SuxpxmJx2H8ZdYF6kIz1ZlQSHSBd87
A2Nce2d+8nbl8ak2CFOOItRBTrcKUM9lStTceAchXuO6TxP/rY+as4aC2PDR6IsUAvn7NseBlXao
XBla7Z3iW52ebHS89ZMrjSngY90PfOF5/NtvtcvFTAV8dE0BUO1bEUN8HJiwpjvruL+C36wMHpj+
pgGfCF6BBhhHWYFFbS9WWpOKFu/crCGhOMq9L/SZNkeYQ1hsxrgjF+iKvhD04G9j41Lmu0KhYfDD
KvctC3XoPNhIt9xtZg22RLdvC/Kej2DJybWCnQ03haeMxZjzsam1lUx/ohaipQDeXzW0y2hpMfxI
HZ3D7uBfxJ177UnDI66JTHOv6Z2awBebwIQjVCyrAsvOylrb+lT72eE4ryiXYuJWCKqhJUAUVpwa
Wyex1O4rJtnWtD4EwPlIErUuK/LpfqkQBEu/OzP/YABaZ+R/1iPgok3Ge95a908ufn2vki+tPVu7
mSbZNH8dNnAb4JJAA6UJ7NdJPWr3e4WItEswsnZScYYLk3/tzt8ox+gf4kEGkmxoIJwLVk/c3BBv
otUHiP6NUu43AOKD4uru3dTd16LUwL4YcHOZcPcL64VpjM2tWu8e9Byn6aOaukyjCRNBi3Kxla6X
o/IjxyWGTYe6f2UbFOaGab7zkm99vyZ4raUxXSOVJjgTW2cBK8JktuPclgYmwLIM6lbCMcqltxvR
w+8m1WHxQMit1EqJIau/ShYeuHanDL9ylHLrFMEUtFgqkIjEtMsEYTOu2TnfRL4ZJTcfpwQsXi0i
T3zr69tytgf0EidXKvvHds0gXXieH9Zpg1krdQ5BHBIXVc11t9zDtI+xwfKGGQrp8EVKDXeD+5Tw
MgmAdFmt9lpN/utJXaqAkMJlkAyHbnrfTSpzl0Rt2+UkUdeW5CxytZyjhocMhGzHwmFRPQ4/QSz5
t7l1uW0A7u9pwaTzNfcJkdcIn8tQ9NvSW9h98QXERTtOb9xr4NVh8dPhVMaJQZbXirbdCGpmrPYt
mdujLHwDFC12v729EaX8ZkcwxlPh19yuXrS7XLmNAtju3US8vcuE0UI7atSw/XOWAA05azGjKL2a
DoSaqXJO89CSp2rCjuwbqV3+44Z8buwJqInmHOnmbzWgmTL2/4sNluXbtlRz6fgsQCwQGV5fDl+Q
ZChNtUsflJXm418IUDN/nCNFE3w83L1mwgseDmyFSYickYyIajQORm4WCVq7Je6ow9uXfKu1SqBT
GkRPvCYVbDziwPXErnX6sAjh+0GwukeM3BqgtVRMl7NMWHcn4w7L0hqfbOzITn1aj7oQCJJS+Ovb
18gHit53voUHPNpD5OOWtq49roBrIS6J1jjhFvuKh9anPeXcwrTEg3UVnoICP8iAz8gvI9502Vhc
MF2A38Wx1EGD3uhY3KWmqiyb0QEZ9wj45h9SVgCLXfAJqmBj6fH7Vx9tvGf6b5S7mQZbzRJs1t0J
y9t6ZNDmVEn/MB97DtTgjAOImMOgA96UKAQAPVU9fae9e6ifau0K+wDXHfEpTYzMcUmJlQ+TMymy
IcQW6MhEY1LjytvhTY1lMcCD3bOtLxCQTDNihRt7PL9imdtdfV0r0jdRNwcc48uN/GTk0gjj6p8U
6EzHZXmFDIxXewCYT2nhR0R+LXpC7uA72uJ5/zCuvc67n9H5BXsiaWaFz4d8C2mgQxg/kT7CyGJY
bBrnhc5agl5E4pjc2Uh6ZSFXLjm5+CKFdQJFgLjyLfTCCsV/P1IKrWXqiuwKTnCFFy03gV3ag264
1ZG8BB6i36BO10nIoP6VAHal8lZc67n9oy5KkMEvlQsMohsNKEzi5cqwvCUaOZISWpTriv3hx2/T
ftfY1savdTU7WzZkiAcTvktp9XE246N/IXtq2MaoFyr7VcPP0jcbrZDxeoJtpgO2mYZBXcW9lw+o
ux4gLQvqFsCM69jkN7SeOcrPJKqoTUqhKeyiV8/5a7G/8+jVCf4tYwv54hvgXWqZwW/RU9IQWWnQ
wTtHB3SgAVfga4RBJfQrTqzk6a89ig9M6Ll4dptxiXKmY/QvAOfDWKSzVNFW5mGQlK8T3no6C/1/
zTuZsC4jSU+4p0jJUkYS/gfUD6fhbHvsdoEi2+1DS831VMNx/F2MUrRb7p4MOHseJWGSDwsTxHvm
NRUBw/5ZydezKSlzXEmxYwZCeaoBkD2ubrZVxh/bsUbnOkCf+4JAlTmNSqwzMPk5Zq6m/XBX1z1S
mXDMjZFmZuGIqP/XCuPzn74dprBTEDBrVWI6Lz02U1ci1X3fKxtqTjYgOMr+Flh7By+SX8iB/PPb
SOPS4vbgoT6tM0PxRO7yP8sN4Au7om/nPVgfVGgDaanTYY+rnkczVDbKgRiBdl8L4e3uvBsh8+7J
6nq5UO8CUcO37j3QBfbewBBOiyigB3yNX5rdT8ohz4OAUa3xKCTcUK/R3RG1Sk0ZrjmmDugZRDl7
XTAyEmfbMU8CFwublaYeMTbSN82iKPgyKiOWQPIDOzGZ/+azKEkiDprldcBcW0YY9P7JAFSVft4u
J+u8Khh4vsJLw918eiCy6CX8BbDXwszkFjhpJKVRWHVngOc8JJxv0lIRjuugXeTrG7BOXYXZap1s
hIIuoq1esf1apZylwDij5MFVNNdqBPiJVUxyONcQ+9tZzYCmsFV+7BZRnSyiYihfOMZBJDp/gw0f
EqR7qDbmvzbynp0tCFrW+QOjywxNeQdqclSet/BEwWhHgUBFtWT3KneU9x284HtQpfSYW6sD+M4e
rr/hWHJZ0FzPsps++j6nYuUalHMxIf8YUaBUtnEZv2I9qPSr6FHGgg1EFecXeORkyBC4yABy8PFW
xyC2NO6N0W9bZ65sB8W2OGtTA+wXaK1C5PN8mfGZeOc4w6TI9AgOlfXUwe0TSCNhm2ko1Cf3/nbC
EyxD90mayhG73Nfzmpzo2yzRjeV1JQty+EaTcRT8C9LKYtr70Gttob0EGixDBw3VnowSOfzNRwRs
4Q9GlmIpb61UKPXwUFSRA2b7CVfNCoH4MJMR0ONJzWHTRtqGli5IXBImLNQ0aF1XI6ZLBKiqPt30
b9HIfa5L1/+tHgr4rPEM3UyfExyZ9caZXbhCazF2A+H+jyWe/H2sEmwBJKQdJ3jNkg+yABnX9iHO
jWmitQEXm3DD6NAxpyRfGxSTndlrz6h8zIOwqTTK76maUS4PAUW5epddYJ87UF+40feahkuY9TIe
R1R/KGsvZleKn8ckemjccUF1tpDJc36Pddnxu0hhs/di+JYQqQsEhRI4MlXH5U+c0dr2ARPp9H+Z
B3EdoIB2orN4azg3G41RWnPp+ORAZTiSeWf/1t7Im+BwLsa7IiCNO5lij7gc4VeGApZk67q7+KDt
12y1
`pragma protect end_protected
