// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
XMaxAkaNyetfXu9gx+F+K1XsiMxXmqEcv2qubiW5xBE63ZNGKM7OiLOncrQod1ZN
PwraBo0x9GHMHjjIAaw5F7ddwjxEP5ZBJM4I09v6kOniq6s56HEQRKC8hCH14cZV
gLHZpCYqsc6H2Fy9kAHJEtDEcObgDIuaHKxJ6yY7FPE=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 11280 )
`pragma protect data_block
RMla86Q5XQZz1I0nUyLx0EzrPoVCsFKQ7ZUlHtdYVQZy8lu8MTnTiTvhLPynNODV
mS6qo0FoUJg5QO+hxkOsVpN6XkvIw5eK4Jc0R7JnlNcj4CAm+R07g32YWzUnersn
Nr/O7zqzYte0QJq4rduJcFK5oOGKECwwDhNMLLLhPGZZzsgMbO6ihwhePYFk2Hmk
yhDTFfA49k+ZsER4Qio3EFbQTxD+Rd02XX6NSCwKhscvzh7/lLGFxLnRK+No/kgA
8DEYnWcis9bcB4/RDUS2NBrnHeZfW+SqVQqQ7bT/oAX3v113qMhkEAwerhJy1uU2
1M541J0CM1XtOBWDcrAKc15wQfgGZhlLfhysmZwS6ZGBdu7AOVUrLMdK5eyyIjoo
56CGHZtpeqoQD0ZS3i0VzVQ1gBghudd9Wv/h7tq0ITpL0/w5lboDj/HM6kHA4X8o
lVwuYyzlX6iq5AC8Lzlm68TTgE5ulXqSlzVY+mM+KwPbCbH6ZuAnjr/RMX+Ey2zK
UBhiLqABZdrcEIG8IlmixcBsq6Na7L/6c4c160ELgPsRgWzMO4HK+Q2+vWNG+Zcy
HpEBTEY/Z5i0HrV1mCWVJLniWysmQ/OiBq6k2b10C+/SAFIRq5lPLvHoF5UCoz6S
FMmOyqcvX3DpKDL3yUql/5b7ne900o8uBvl5rQ1fTfX6hDPi1zRj8lGi/NQ14BkR
+aL6rBtG37N3tFyjzihSdCe0SEEZJSCgVmlZI+VY70siladhvr242NN5lTTXXxiq
MI/p1BC/79yfPPEpdZoymCDP8M6N06OusAlk6mSxyH3KNcHpV+XWGyvLaKFtamHf
i/tBOW2TeWE7ANnBJ4imszWk45vnzq95Ja7TuxHhzinlAjn89eQMLNUQjItiCJOu
SbSpHCV3bjaRK/ZnJIsttGbvctOrQiZUX0qyxFfsS815j99NDxnWSPSk5/7H1rnm
fM3M4M8/ln6oRZjr5BckFv0AMkNi9eDbQ9vfn8yGqnCwDWD/9pP44JBa9flY92LG
lck+xfBB+fEiByFqB5eIvy+AbhXAOibcDSAZZz38yupIf2pqoHG/e5tfTpaolQAE
eZIlq7vNpdbflCJKBVl+yaCsrM3gyJsRPl+/CazSEPl9byOypt097HB1bQdBCIEI
4cjm8ktrr/BztO3Lm/H+4kSCIbFcGeVzjUddGNMXhxc8K9OokjDFOWhPVd8pNOv+
e4vXJYCOCVxd8B96UdvHbkkYBJyCVkeh2rRJrVsoVExhGATBdI5QWUzJanGFJzJc
SB0BaHbjEMej2fK6ROWTNuggEvt6IxxOTZe+5eICtZWA49yPjoG/VkBqbvILi8YV
u38acDPmhO1kaMisjej7qZ+Rk8/xqK27+NfABeWYymjuKIuFR20QxeJ8C8qWBT+u
a8MC12ZMwwEqW4DJSunLcgnF4h4UVA9IVtqXW57tT9ZSLpvnZpIwbmdGq7ti+abD
4Fnx4Jmgu9u5E8CRzooDRythNyRY6y4FMQHVScQsD26HFjJTSi6hiBBDHKOyXTVQ
KpaS43nT6imObodYQQzzwrzMk6IOsXRoPAveKJDJz14JQV2sOAvgP3NlTEGU3p68
S5soGuIyr6h3jAr6BkzkHhayWDtFRF8JCAqskNtBBrPiZaNQaN9UkDzDjhC9ztSN
cWqp0YuvsaMrZuhpO0bya0D5ak0zq/f4bIAymmINa5dYmxzQKdQomYbkf9/6L54l
V6Sl+C+Hkay98tYELD5C3Xc9K6xgINpT9x7mIboBYd98yldvwdr/l6auL5yNfoNS
G68kv2wWLwuYrWgGyZq5TsQzlYQ9lTrvugXFOv5Y1r0YLzsf6lRh6qQivFziBSVq
XeYaoOdNVznCJsX1fX7PgBta6wJtZ/5+7eaPZPAlhdH/B6YkiIUjhfY0mym0ol+c
GVd04JBFdNEMZqn7/Jtf6TvWYQxU1Ggn/2p1pYnD+FMQIPJTcWUrfHS+YMcsRfvb
DfSRxWWTpLXKTVd2BYRTshE6WNpnj2HcNKLsgm7lejlpba2OHKwEHMSkMSLW52v2
9PRCZQ2FluBCw+WtbWjW/A70xkWtD/WMcJShiowu0CW1/PRU2KzzOFMC0BBnctUi
uaNxKofznvXyTAemembSCKZKD55AEmRRoZtLnPlcAwf5ghlh+OfiGuqib3etOWtN
npbsO+au5PF+8hQD3sOx3M0io4CHJUwj8ObVaBpOd29aKMgkoAWUTxRQx5riQibd
cFLM0dBkJGC0rSHNczAiXW9eoFqR9Lrc3VQOJVm2OJpl0C5m9T/6xAiBMtz/nxuF
m/FNhzt+2dzfYfKT1dG8VuvV139w9CmqmbS0THB+nR/N43I1eGU7NB5lYOWCdNFU
niZrZVVprXGgQy/ZPNwE9YvN8J70f7TtAHyKkeL9XDR0yU9DMnCKPXVECvqZafLj
ngilzh6DWP1418kn33SjZPe1GS3twTtHJ2rK1ps9YS4hQHbstVhfnudUUvghBSaz
9nyaXENsLns5twB/bZastRnfts8dGVIzi6scYO4IVgRC6HyeKsDHA3zxWBlX1Uil
TleAAYiJdiEyxvWBfyiVL0EvQ+0On9h9/IMMK4VAdDzdNoqeA+8Ca8JL0cvk2+nf
ATWLl1QrkwqhDkwVJasQdwrodKf95gP2fZV3QsKXUTYGu1US8Er4FpM2FwJshM6J
wgrNkcSH+PJN1qOhHNjVR8XFzzuXJzzeOhxi0Cb2RnIQ0slSOKOZuo+78xjMKTx8
1o4q2SJI/kI1/E//eUfv0zjqcyEJ2v1sY4IruzXNCf1a9JwNwEifR0VsdBSzLVi5
kjibyUC747+RNfiRbwYVbbkJD5jqYS3bA+jj0y78cgIZNIl4W/tCzzejsoWl+7sH
TObPNlrK70U7/3EQC+8uzinJ6+qNcdJ8ADtRC+JLFOfUrVAxBfPJxJPpUlYi9Fio
JZ5AvwZ1Igjau01n5+HmvfC7jZckRsIYoe8/sVpRJHQB7y1RosHpyrpEwb8ykgfw
x29wrubd/1Ra6Rz+Nt06WW4qRppZFrAYCeAIuNfVLe19qtIBPObBNu+yE2+j3uhh
xHVMEYntWBNTQeHDaY1BBibP+P9yrHBbcrv0OrAVWcVqPPjTDjMimlOU5xFbPLTX
aDyt3dzqowokmBKRmpk2ezGJx25xjRCW7/23Sle8Sez+vdNTeE3PNwwFTiur7VQU
e/L1rRxVtCzv2UEXdo80Un5j4UNmHIuw4x81RGEaV4LYv+GDUhhn2u5GSQcPE2tK
pRFpzxXvmCXQxxHdmFq7FZbkdCouhRCQY0PmbTI99W91+wFiwno6gQXNLAifRYVd
9+4R4mxll8q3KO5TJ2BgKIt0ZvTuPSQFUXdDv92d6Lhpb9Vl0Q0gq3gSy0m6BnJ1
H8VONhQ94E2mMhIPMBk6mV8jWCu35YEhVe+cXB12aH5OkPP0PCg161kVY03PPJid
ua0z/fCOMkURxD1korUG41HJo2jX9K7171bBas0UnWUChIicn+2q1KdTFZsxehnz
C6QtyjQo3t1KlesgafEP2xd3h3uVEt/2K4uXaaSMenxjdoOPb0VnURzkzYIHsS7Z
Q7xp0wDbpUxHx7W45JdRc1N9OZhszRZDjtrD+Z8x1Q5JnKEuFC57kTrL1YS1UYcx
pUB8To8La0wQLpuomGD6UMb3lEYx/ivDXSAb5hQ3ef8omfcSZIuEcKkZOSb90/86
L+uulzbWV0G0Z/lutoCpv2q4tSFaOache/b2t/p2Hyfjv7TWdSEYWKHv0XK8x6Sj
nN1kgyBilBjSP+P/ISo/+pCafosPDilzNNA/cyoMPBag65PUQaPkSK+nJxgjU9V1
jYecJ3DkAwsr3O99qzLqkziwKLO3axoVqjOKmqgLTc9xCx4997MHEFP6oWK2We4T
YcrDTIYX+uvqvAP5bweleg67qRZXsN/80P+M6z4ApoiEcaiigbUhxPy609ba8VB4
OejrQeR2jYhErlaos6EpLPt9LAX3fBWw5pOlZy+2XmKRitGqNWyLiabUYHl2utr6
78NLm6amJkOL/7HbK2c2xVHJz8XKgmOn5IuZQB7qDyuq9+//0E2lMPifZPneycyX
Lrbgtu9DNuv1g8++RNiOuSyilpDIYS0kM7XlQWID/7rexqUHjKbbC1j+WX5Ieguf
Fnury0A+tA9rrxMkeoDzzIHBIaDyNejzOrozLRnYXo6eUKpwV8LayKlCDVHCbo7k
6jFWaKVPTF6L/LafISHgrPJM4EzRNpgO3WgX41rO3UOIuM+6d7XRa6kZc7yw13Go
XTo8GXYb0GQyoHfTCBrl98S+3Wr6BhRpfZIN8Eds3qZoM3qu3NyCQgMjXM8BaXnA
6wai4Zw7K9h/Jh/BySwl7WHQU6fMfXGXSZV/T3+Qw2WScDL7e7bvD6o64fx9KNqB
SJ7sG78kzR1q8JJcQBWwDqJ1cCZcPvUnPQzPj5UcYrjcngcHdMF879jMG4VZ5xF8
7cAUIWMML26RJl4R8cL9yID83HXyzKJUBLgkepGTcK7FUnYtNN0Ono9Jmc2xO482
1QSVatZqoVNiVtXBFOzuBdd2RMgFvcVAZYCZtqI/12Zr953w3+0UUmM8m+MKsV0c
IHR3215RT7Ig7W/46f47yMeUOR6BON18Br7r7y4JW3TiDZsG+AIVJUOxcPY7GD8Y
0ldLow/cKvmgAiw7Wd3loLaAkfEYDaQcgp8AxMHsaMvtfpQ4RbxuI3N8dgPeCCt1
4fPnaI9hmgvYxGEyDXfwvV/8CiDi25OT5DQ8iIR3Dzbc70EX1BviHtk7wlcxsWzw
X8/wzPfsbI+GYiz+MuJ4ozGYNnKEkvgm+5xUpm5ynqfzVfrADZ/NC4+93+Zl+htN
2HMDDotgST3sC53cqolwYS3C0Eal5ac2W7rPZ1AUWefQFadDm/zRCBIS8E6nuqtg
FH9ZLGBlQ/RwCBySUO+d1uka3o46EgjlTfrNS8IwAI95BZkR+/17cbJcpMXc/lFo
X45RAet3Gxy5GNVdqhc2PPKXLlBB3vAbqm66QKiCQ+mFMQtMo6WhT9COjYcKSRBA
ZhBT1O9/uhhd9nMz9SaUtWZibcBiiXdqyANY0zUPXsKdOzGmTn+HchuMwU2jW4iw
f5pSjWlin5S9f3vtVPKPLKvhIs4vVwGqPpKBoBS9e1i81y0NVX9SUqMd0WlQR2gq
VOjCF3RewS/RdMrzMVicm1bq2kz5CFjFVndLce1bQ6cGCv7p2iVH3nV35qnX1N4y
XZjct8egyqW/FAaWtCi/PY1lG6mBn1dxORzDu4qAXtR5MiCiuIqnHAorOt9f6Gl9
Wmhs/mFtIwYA7iHK3NXemAG/w5aQnuNxSlT1wlwRT3HvUTVG5dOldisX2S8jE/wy
WG1FSW5u5cpYnOVN/LmloV+YTS3Al89APe4ktDEY1ZjRHZLeqamZX6R2gK5eFXlC
ShRnNl7nKCoMrtdtZlAJjM7lLQvRvYekY3sXlgc/VQKeDSYHxN6jBSMp0OZ+O/VZ
Hl758OadfwVxRcrsD2wjsD2Y3n5gedQYNLvoLqx6qtZBo7uVm2A0cpsSpUMz/Zsl
0f5tE8zMhapgpIsGTdlFVlPoab6H4W5J/C/kCKG01ycBdlITTpifwUatLDzE/EKA
kpiGAvfxxiuIpAEnziNgYSNpNHsHf/ETDTzUQl4ctnSJEas6x9RozsFAKexj8/a2
6CR7fHB6SeZne5K4GoV3cREim/2EewyHTVGyZ+Q9bGnmitq1ls+XUJ4AmMyvU8+k
UjtUjKv1X6yBAKc/RjMs/dYax2T88oj66H2iL87YmHgDv6G19EAc/Kfnot1jStot
cKKJHIYdy7k1PEJ5HJ5qs366DyAdDNlvz8r9D6zJ2PMGsCeqSEo+xbM0ZPXSd/LY
ddYXzVh2ZiODW9MM/sI8PeW8HA+dFOakKENgV1E486MmYxB8eqkEKMXReEb5rS0/
vEzcsruDGzj/82GPk+rVGz3oluXlqUUxNgP+5883QDlnOLf1Zo8O4ej7tC1xqhyR
TbfH73dpWHhlSRUtulRT8RmnxnqNmqpkBOEk/27yZVLpqvDleKJse6XDS7s6myua
epkepOkrB3lVRgRCSDn2YymWfLCUfkGreAhvJ0fSh8NZITaxsatEGqYgyGfsGTiH
T5Kezp9bcSSYFHznhln+pLhHZwXKqYSnBzi5y8kneqokVznMUOTgqKPGEcn+2DZ7
w+kpKCIk8ppuvd/HV7n01og91O8Ut4+kHtm3/2KgjzP6WxInLKOUCBN2s/fHf0IT
gVxyzxgwg7gtudAkefjZ0ijiabYtjNV1pvSoL3GoBdJc5epuH7y+F14Tlk93Vyb9
JhBA/9gs8fN6zeE9x7dulBewyH61HDor7Oh0PTrtpMytaH1XJMpoCKYM7+VAjj5D
VybcKmIssQ9GYb+KlUCs3vlGJmXK7KUaaYj35sA0+ry0Qo7V39Q/NBOJ+zQpll/8
KdSyjocfHdiDq+JRyjszH+j791k4FmHYX6MtSOJ6Y6Gh0bSPXFt0qB/Z2YCVebpS
d7iXW4EjqbozfuaqPs5J6WGkrNUpqUlAlqfGTSKxEJNd04myK2JPZG9ccJwzE1sA
GBxkGpQ5Y7pTGBbNPSB5E0r46VnRin4bOEwKesvnpTgefusbwZMob5ZRHTyxmot/
iQSUAJSJGHETIdRRtUtoDjs7Tpcti7bwWxVz0/mHprS2rWChmXIwvHXUhNA8XnQt
bcrQ6nSpAPqnBZ7vnLAipoFPAmwIITnhlFX9FmmyytMqug/sQJyu1QvlownMtuBN
gKr0mE+eLkHBsFywMfUAgti5IyPhPC7Y9/xn3DvVIDbcAYjk+2Yx8NC3hTbrA5Jl
hAVam+XTPIlYU510Pf3GVddvX37sgW7SuturnnVLwPsOaBPwqJSZxDoWJzK2fCvx
XuAe1NZYqbXnGk9gBudZBLdGZNOyHkVR99DgZa7MGPdaL4W5bhbVn3O8MdiOCImq
rPXZjULYS7wUJB+wXqPQJAfi1bOpZd0xjlAcFXDGFlxcDiS3vTzBwEiHhkHT+3tF
2L0lvHmyaCm0wJlPB5C823uB9ul2gp2XFZKSHlaQAZng1bozAZOs0UGi3Y/LTmHV
+26v1ZJisJXCE4Lbben5Dwj5ehvYJWP1uarmbHEhNCRGUyt5CqpvbwecH5nGk+L/
UbJHvn/nd3p6/ifr11HIX3VHOApc9IJF+BvmpEd1gyW6h67/m9L7OGZtSt1z7aiS
6jt+SCuqRG+UdE2Em+UM2f8U/le59mCfXkrOqt2ivyaODyOPDpmE9I4Do2IzCy48
Tu3bpkThD/IewtNT7vPXojA20Jp6u3r5CgPLbGO5wpPi/eVk6ubrt3WDnABoSsAP
AIAIotvk7RW4L98gorLUWnju2Datk7qoUPD6JejZYxnndiNC7ezyx8xaZlgThD5A
UVqPb4KAbZf74jlQ/FcOCCDPulniImVaShpiKRnoMfA/rBqXbyuojbsxjm4Az6HO
INoWlk7UVDGXTIH/ijTXGzZAv8LrRyGYdhlcEbaBSmqLwx9Otdp2NLsyEjgD0Bqy
1UplH13aXwGK2LX++MPmV71amXeOql9AdvksoYNeboG/hWfk9ltTqu4VPtqa+CuC
JMO7juns4oxzRk0JDjs/WCDPeqRUxZqVj9YhyKRy3FaW877h1YHoC7x8IS9BxGt+
6WAvhkH9rWxePwXUXlBHy8L5hLV5CkmAxYbLh1BV/gdJIB0LFTRhStR5ObnP6RQ4
1bcDQb3lWncqCasILDmJ/Z+BR2FCL0pgEtAxoX4TiHWjS5O8sqT5wjlZcibOrJWV
ypHqDtEVuWxCp7Rs2lRPiPUH1/dX+6nawkt2IJfzlYz/bAtumqM0jXcTopeZvuZh
TilnG3/lO010ZpSwlqv4jLS/C1YT9umhTWCxF2BpTA9KGWmf2oCsO9U0jyrBCKNV
J2Dzn6zRvLq2bkjcSUwt9I0QNb7xNX6qgmR1ShQnJ6Ij2m8hrEx3Bu6U/gFmoWZE
Loaeci0lC/gyhPMjSaVl0Bu4UscWVGXfTAzk0YkXf2Vbl31gTLavnCCSX4ogaTn6
nC/NSgPkR5HZShpjpW/Innal9zorZ58uMcvKG7/QvX97ZiNLosmWlIBrK67VkI2F
3M4x3XOzxLvRy/3DkTSDWLJ1Y8NEyYDuSsTCMAGA53b6RfVL2J0svtclzjNrtjGz
DqENd8bCdd519tfUqXBKbz6W0kAcGgvA04m5eYPZHfkUct/gT6yXn3Ng3L/2z7Dm
btqlcLJphV5DKc7YQ6bdUojlUXNs5OtOhb8F8ZVr7tBSwu+bonWdYfl8XE/eUdFf
WdVHiiQMwvpUqPeOKw+CrmOyw+KUj3BAkjowvy1ogZSET9Sb3XuKN0vyGiW6Gjfk
LbkNQyV3mvZxuERf4QJlW37pLCoLDYiEbxqXWsdSixO2lbl7MG1raaFSsaFbnsdz
DhMgzZsOlw6JFRHwcFpruDFVYLLpL3topPGxtT72jkCQxdP+VjrQ8o6oLY0bHvtu
RevXUo5/hb/qTHmARZyd0c/w12tS6Y0zVbIALgalyUrdCTV0GV3ad2XyX6csderM
1Uf28sOSXwn8v2LMcjd5jeJul5mDKwKpOZGwopCcKPcdqggzChqmm/2tSvK1GYz9
WyBc3uQ0WTjtKZ/pi7QAat/DLphNR7265bQpLxAFKhWY/+ofunc6gMcgdwvyqy6f
0ckku/JjzZsL2ZVEz2dWHAHLWX32EoI4a9vQxAktrXzK1lTx92eqaD7DrKl4bc/Q
qOZF8I8SP98CqnJFUXZQCvSdZYugiq0HESXTNs45F3lATpypW8qn3/2cwyUzeCYO
kHZRaBEyk9zJvrWQ0ASEBj9tHX8wBtDb9xKGCkTJvqISBe75HtB37iHSxopefmuI
VeJ/wfrWNxWl1rY2XEYWV4aeZqv4tiRea2OY5dxXlQwiDdl5cgcg7wc3ORG02FAZ
Mgbgba72iR8VoZdOIceCA4HSAOafonrWnQPW8z+rjd4bFpHWgqIaL+UGHzTvTEAO
a43R4fGO9njNXmB+Q8wR+/YLkmx+4A4FAkhmbRc+4YuAXKei78lYSU8azGnO0JQt
lzzC025PNDYSSTSrtEh6jhsowHQG6PPoOlo4qqtd75K3bBgbtmx+OKNIQpZU/u7k
M0oNVrU8v1dYxZk5m09LlROafwB67bgogZgiUUcJBPGNBplfrC2PpwPAv3qfaWtN
mhHk54487mNHDL5+jX5h2xJwe7G6Xk5rq1vSaTKLG++1ctsm70gk6OGSqOcBvgE0
dPrDfwUO2Br55uySahNk1e6QSzuYJ13jYYd0tU5lmEPMK2cIT1gTngxXonaXBgZR
Hv2lvt5sf8az29FDLl4ZxbA/bArVaa/haM7LLs8J1EyNOQ+SgWNMT5Klb8eHdBpK
hn1BM0zLLqWpL5DOIYGE/tcBvJVWcOLGiYR8fE9uAZ2Q7lsLcjdRYXz84cy0IyFN
5FXqYB5sFKhZn46if08IjXmk/DxQceVJAJ4T8c22zUpVJy4mAczrqO/XoiFHtsq6
/OMq5gZpDcGxXNgLGCPi4FMscfcxB1RZW2Lo1pXr13NQoXgxFmEKzC1mh9JpJu1y
57qjTllE9LeTzJ0oUEQAuU7fIaHOypMhgdfB39epjPTvPZApcBfZW0BllQmUMaiR
qtng7UDVjs2e60ZKqJqikpDJUo6yvr2vGb/gMa1MAcNXewROgqXLKiU0FPiE//8x
9n0QayXRw7ibB1z6IRweZHt+8sd7eQJ+tAK/ASop8U5qbpgb9Seq+nnOE1ZO2Yh/
FptvHE4/rhUo9Ryd/n8cByWUk7fvqgXwpdjP93zQ4zl5aDrvp1f458srtupXFtwY
4da+1iM+WiTJ4s9aqX1VC6ABJNmTGoi3Hzu9tMzcl7BGnqUv7Gr1Bh5PSHnZq4hE
c+vT0aDJG89beOfpXTikFrNFrL4cOxu44+URWFCFII6tabHfPqrecCMh58OoFEQi
YcRgQrBaYDrj18G7lPGEeAeCBTgaOqBP6F/wJJ5HIPfyrTI381sqyon6Gg7Yrj/F
176dTczYJDKv1YtYmoQTb69uz38ixfLdCSshNON7YIGrZcFuOhe8s/zPHHRRdQ6z
yvxy94Y1Msoj5m7YTgnjZfuf4ZSTwDRbP1CZ6/rjAOGzoSdgE+42rU3Jr/MKPLQw
UG+eEHyabL5KexkFZnFk0d2xXWg5lfkRoVdPlPdb5GmEvYiQPplQx9fVw7oxNKgW
csdSBZRl9yF2WSIY0edplgzw6On8KiGroLF6/HIGCGpVC6rj4JdGK+sJmx+yxR16
0zUvMLPAs+5wEOyXWU9AqGnrIsFLFQa3XZvFsiS41H5/B1clejzy1auAIaiOeVSk
IvAebUfET+1gZTm/x+9x7CbuJ0Nmu6bTJd/joemFRT/u52TFDf73iumiT9cEdsuE
MObUMVRMNmTrIRbnPO7Nkqz/gyFhpxmhGhSaQ/14KEZUKdhZMJG+93POv1iTkoj2
GP9M+gKArjlbdJ1yYCzqaJP9CtzJjlSzNlO/MkJ6S1e2KKmWMuOFVV/FE7jmdb3D
wcjtOgtuEu0o1RGrt26djNZI/aRu3UIFj3hB7bchE2PK/bQ2JjVHyII2Ev4dhkuI
RZfPqB+eaTNi3X9FrKV4hKBB+XcUoPM/z84oIlgsV3opBujW8ZEPMu92+ieqReFf
xmimqfgms2F32EI37FYZ24LsK5oyEKXjHzhya5CZgZCFsRWN3u1PQw6dty/fgkjR
l0iHJI3eXld9JXB5U42dmmMidh4hZ59bweMu0vCndL3/HMqlAn38v/+RXPgmRoMW
DnFGsS3YPheeaBG0wR7NeusdMyyY+aLehVoe82Ri9udz7QXKrHfDLh4ajx/7chXc
ONzD09oBhlZK4/YOHJquIdstOp/CAQey1yawlt6IdKBi0dbLIsBGv+4P3HkHrCy0
rnKqE/khQ9lZzmfyh4blzTNbKCdL6/2R1Fy6iGhO1qqwYBOTs6dnxOzXNBqoI2A7
XlRVsLy8TSQgHIGN5Kqd2Ujmg5covlGopBbZP8YYB1dfrC7l59Hbvuastu9hURy5
A7Emp8Jd24WsaFMBVwaAxhu1ZBIRdyJW6c5NKLdW3Fs3pyRuMOxDaJ5Z7P4zA6OG
mIIqzipP0oY2ZSQTQV/IsFvZOtfSwc2mZ/KY7IDHJPW0GdKqdr+A21fQXWLVkkm0
OO34J0DL0RgBM4jg2qeGkLRvnBKSy6Vr9zbUnTQZZT7awcdS2t088B9ykFA4C6Tw
C4I8qkDrjdpDxnIS8C+KdJR2P33qgXEHDfYQuMSC8x8iabRIsX1aIde9D5Bq/vxt
5YG2Ydh9orrNnsYBDSBRwfdT4hWVKlLQrEogUeeX5T1rzkjAZhwnWbJVN2cSbYLd
6/RTkWYbsUjoQsy4mXXasewB/fJn/RQ0jjYnTEWpCpKM7ZuH+WmgPImwJf5PXOni
jwv4C927Zwl6srE0mLjw/P0xStEoJ1Beu3qVvBJhwNzBphosk0a3p140F9pwKsMV
MS7Mm4H7z0jzLBUaOP7qMmy3PwaIn2pOpg/0C/yyxgbR06u7ChLzTxf/UgJLe+4V
PGUYER35FCdyuxEnov7TWv179ZzgnIcX+Lio4J7/yetc2iKcIWd7gQTzvTFNOY8x
W11tMCTZA1ZrB/0UTMY8H+NWs4HQr56dBDVGYZucddA0wACOpHJmH74ymP6P+NPv
L48Ht2yROPeJm6ExMYLspyOSAfoKCD8YleNrysZ9l2a06f2GJXRcKsUvG0jywNX6
KZ04Yr0P6UcGUY4vo6jdVMpHGTdAmc2azu6GV0fN25VeeZUZN5gIXjBhZaatc0Xg
jgktKQxuEvTjcfqZdY/uHt+QlSqOsrS2oNBouzo6+sdy7w47l8OX/tluGMwWSr33
zjW38sIEPB1lite1mqOALfycc5Zkp78ZcVZ2QDa6Yl6ZtvXYorK2NwDpDRUNMQJF
5/0ookvnotU54I6j/yVklyvxD4YugpJXQ0Mqfzvs4MZZ3Kc6eIO/b5q913OPDDV4
tlgQkSNajUfhgV7G1JOgWj+MD6vyJBg6nJJzBv/RGoCcg++bPm8Gm2MKg24Fwhy5
DjnTPM+F1yyR3QjfCalREGrDaCleCx6wxrN+xFeLe5a9Fz96KO9rTUZXRSlMDi2b
Fy/Jcrk1l+iF75V6upcitJVwjGoKtPjPa4nBPq5D0+mvMtOBuu48uXLCEK1dc0Qz
8wXgzhkSC/UmmB92sCNKVhBCLPDtGucaj7h5ziSiHCJyyc9KNC6U6orgEedHrY4z
LBpu8d69WiCc1kQuwimRsFp0ekcCGl/QvP/GIo8pm+pbqLOgI/8JBFQyZsKR0a1K
EStvtKoSYgtG2k4X1qWw+mNDUFLa8pWKLLR0Bqpl+npo5UNO3mNpds2W/GfIunbC
LbVQbAX1VFEKBKlt+zahn5xXLn1bZ3EN+7VBIMLX8QQ4gtZcFU9cWqMNULqJAU32
EFfL035Uqztw/xkTfaaL8lARQ5/p6YANL+6bUiOh/mIQASkxRel0z/VwNB41Uzmi
/XE5X8y7qufJL2Y7fivQ2GJxbAy3ReBQg8IWReiWqliEfn8b1w9hG00uLl6rnUjh
K+wdYY3ZZGnqK8upR59pfhqO76L4QVl2fWGxFEIbJKGWMWg4BofkqjOIQicZdN7l
b6x/YaxRh+NIJSCUP9wwxHGGU7Vza7/g0+owGf4lOFJNAkD1vcVuL9QO8id4xGQ9
bg+CZFsPnWohaqFFEmts7DNmNMetCvnaBCmzXuPEpmcVg7ZF5I4HzflVQs7b7vbA
q6/nL5YvE4SHdzKQy1Ou4CCPw6mbghqA/DKwiGv3VB8RTG//X6bPlQ9fWPIDYybs
CWBW4zSXpJrAU94gL2waLTMUCfh+yyzYge1mhCTjh9ltlEJPQ/l66UYByjBR9kxU
Cbx7s7qFiHrIvUNcJz0lHzClH5InTwEY22RD4ucDs04yK4vcfPUSWV+GbkJ1+WtZ
ahsa8/sCPOttLZNRYB4XmYkqcxbtcC/b3rGLn9eEYQxW3z/QlCeTB1HP6oRlrVE5
z5P2Q8ahYh/E+ewASTo7CDUaBAAvRFNqUG/9lQMNmVjHCsUt3hVRmf5mKtye318u
k93Gn7hfpMzRFWM0nhhQxofNwdl3H/eYOPU1REB7DGKxy2B3/1XJ2CF/AW0Gm606
SETRJJxPHpmo+SIThZtGb2oxk1b6969slJBUbOxEm2Raa4w96cENy4YU2SMXep9y
Y1V+e6SCbkg/oB09Mu5juaPoVdJMq5OvYCPVs+7rIZVIk9YfdRtaqqx8wz5FXZkj
d0cQ+U7pYt4Xv0RsZr1TgPsY8XxzkSnB7MOz0HGUQR4m5rkb/TQKonGL8ZNQ5qef
xP7kULgpDObhTAz7gDXSzvjjMYq/Sc5hggwD1axBvvmDQZa8vEr9a4O4CvkCLQFM
w1zzbb1ydngr19Fd16dZyaGzuLsmdMEjNWYKYgoO4VkdEdRr7Brn3WaGAW03SxrK
mZStt8ohlHjwBI6CqRlzXBpTOOBXNu8gndVSEhgwqB7cCzsX339wmJr2CfVtTBy+
9UkCD67oDN7OyS7RE6cXSfKnUbyr8Agp93/IjFUgXes0on3tCeofV4qsgIHJx87n
+IYlaE3yuMo1CeVjJDEZpFFvj6ejtprBjQklvUZoUxy4Qphaw/xkgM1d14TZU8XC
e6U3jGdFvlXkU+oJafqDR8ZoQ3NOwH3X7Us8Ignr2H1205Qk6fQVO+cMtziA8Uur
ZSEQGfSn6K73pB1gqKi+CMdf0EmVQyF1Zu4mv/rPHlGVSCfFcAbT73XVRPZ9vcpv
kT3AVOaHfvH5Jg5778Bqt13/Mq67Wr4gQcLmkrWhElbLu+hk515ezpoDdQ/zGvWC
06YWne/zIUttrNlryFYQ+cVmeBQk2kExtTP1QdQzBPwFir/mZ3ToTiKkVT+4qVQT
TF8tFCWhMHKSXma98goMnmmYyPHxQ7qoxD3rkIX3Zkk/FLsG0BWDDViou8cXszb8
aYcN/4t1jzfo5HG2Rj4XKwP4joPh28MR5o4AD+IDVdn41kEJUdZnZ+zMaJPD9tfy
hu/GPaxgGqC+GmmdU63OsuSw61Rgq7+nv12Sdj259EdM1Q66gtWAwqR79YyKrqVA
qkr5BWd+9PLUtjhR2roDWy1Qkc4CF1G1T++Z0ACBuNOIH8TI7PwL2oYJhSxFSYBW
XpjlVS2Hj9SuDQBwtVYH2Rs1C7fMxujRwS78sVbYC4fbTHYj+NYlAV4c6xicNkEM
OW/HlYCQf0zJrzL7dh+HB24QA8sgY2snan+0cMYu3hqw+em2dk6Hf4g7erVYJvxI
dDAwXp8yWc6V7ze/hgbzDMy6Gd4h2QNfiExofc0VkAnFmyjZ76oFeYzkEGBBVhSa
Kl7rGG9NjTKNC+ZDIJUttYgKeBDHtAf2aOSilsNw1pNWFgUo/GL5C5ZcVpHlfb3k
TIPmI/rgJfpScSHNuc9NYdrhkjZXgAQrUZPRP+FOunRJWqIKCocumaFtkH9B5p66
iw3+9scW7+0IUjf++xoMQO1ASDWWavzaMgFeobDVEd7Qn+4P76cJ+9GN2dqUB5Xy
jjJrkfmasFeCFNe6Q5mfv9QgLAzTsfC661MUO/Zq6o48iAIwCAiio+qs+TK6xQL8
MswkoxeEcbWKl66qzElmQV3mATCMfCJxOP7q7Kf2WBQCoZ6US/LYkt0YiSlDt2vk
UZPYcCqpJyj3A+Z7oDzIupD5tm9y56DlG1kXUWbj9tpPuUE+Z6l9KALSHEQ1YSHZ
V5OT2psBUL4UKNTrQUNdtk6ew0k0QlCJdUoWFj0tSaJP4a8Wof/IX0Nn3uk3auun
D/Mj13dk0mkl45U0ggJsGirjAsVzVhAJnlKXBhcptlWG6zuRDQeqfWcFVpP1tL9e
OIztOGGsOx5sVq4IywiFHE6+Slre/P/mYWogst4kRNVcF0+joOyb2/O56xKZFWXK
xKbzOAxG+5cxZXim4z22neI5onvUerWyDsRaG1nVxyqgPKvyKxw3AgOnpcLwnRbE

`pragma protect end_protected
