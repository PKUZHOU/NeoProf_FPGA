// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
XXi2Jnq9X2KgPl62LAacmS/hw3eBb+g3BNOjqj4EnNRrgqTJ8bBRPtGKO4qVcmaS
3rCxLJYxvkpteokyut/l/foUFPXwu/w2MeZb22aCrnN6XCb5nRoqxcr45obn7kiO
JEv49MiQrBb9u2+YtFBZt2GIfU5g4LhHDqO1V+T2r2g=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 24128 )
`pragma protect data_block
amhyylCehXhL1oAXJy2sRq7R7xoTHw2I97bwEdwnNT1xpE9pmJB/rlpl7lOStrqG
popqTGPjSZCsUOOIH95uojHp2ujsfBPFm1U/d8NtE2/ZLGXZkgIuGDcfLsNv9gQG
CgiJe064SeriGMMoszhuMi1P1e010hgZ2iiD7N5cWqu6+D0Ua6Zc5WI1njEyVto5
KFsGKSbDh3jyc1yNpbbBi2aL1e+MscRi71a6hzrM9gFTQtkDfhCKFnkR1qgUYZSs
3tKZi8xAqWgA2NBKu6tYTbsQrl80yy3O6PgngXHTWM+HFqZW/aVjTh5Nfj4K4lAD
LRMszoDzUdRBcqiqPBXI68kdYgTP3emThtPz0zu17QGVkCV2ijqGoD6SNVp4aUlf
yJKXoZowDKpIHX+jhsKv6nV3uk+hk0PMsuLzWctB+lIEDW2v/2pVQ74tD/1h6QI8
LHhBlD1lv7BAA6AlGq3UhJsQyRUlv9u8pbE/U7TSWjmgYJhXko2MJK0dtwofZwA8
mygERpZSJU777urJJBNsh/m6e3DvlLYw3cJbHyB1Xv9Cqn4BodbVz7ZXUldrHhqD
xz+gOFZjQ8P8eBNSk7LVIY2KBkW28EyOsuo62NWuEs+dI5KDRdK9m4GkNoyg/GwE
gF1QM6FG9ec4I8PH/vJXbGVkWBlhxg0wC1QnreuuGihFz4dXt6TFM9fkzr9kM/V8
rQTrn1fct99fOmvV3tPS96PdIgaCXsxDbR1Y3tLwX3XfvpdxbxdJ40Ua6QUT1+T4
nHjcXBPh4mDrUkZDHm2Lki5VKfcPYoLN+dbZvsvtM/+2DU7cPxZEEcBrJOMFdOK0
0nt85dTbWf8tqnjTP4W8pbH2iE+KK1Ar2Z7LSTskxdpQ8UjXv1TMslY2Kpx/w6CC
reXxzpObPZYsqHMlzt+ycnJhJBD4EXquJGssX9wVHkb2/T0pUex/qErMsb00EnhS
wXpJDwIo9+owdAXSTOFqpfzODD5AgnN11VjYenqGz1beQo0d5ub9JSzGB9lqxrYj
urngr7zP3+4+T8MUNiax481/aHo3x3Xke1cVGBYwbgLcQ1OUNayhTV60tXfM5gIT
CfJkYGD3RIMSseJtC65xlHTBYhlurHAePB+c4yt+L9BeQGPqBwLYSgXx2ogFAwdx
n8jlyBhXYgQZI5CGyMUnxMX66uNrnuKgIotCDQJp0iRF5dEWQ4Saiwfzy9upSLjs
MP3AQoenlidajeEW7aHAmXa3VEqKjRl+sIGsFrxzjqHxJL3b1YNboOeiN+QOkBQV
ek4hgbUknrvh4bMLUltPiWqgCSVM8Gr0b/VYLQKI/gykwmMjooCV7PQi+SBfhBCM
vCpaZrpN47sIVNFDcoXZsgpm+7cxdm7ajwwzmmkVUcEVIy/C6mdkjm52icUyk/qf
bI33EBZtgKW+vgcoo3rTXMl7NFZD1BNsyMcALg8lzb+peQY3+5v4UZH56tsxynls
l+a107PiirC7ts2UKt1NpeDWJoEPs9CoQXIhIA++rhB63+X1WSUSg5Nr+RW073KU
sqTz+f/I0M4hrU/XgnkMtirty5US6IUO7aFUjjE8YKk4W+SEDOs9D5ib+xHpkDWo
mZgE1XABpFVLySqSmDCylHpT0lzDdzDDR4qqewHfwU8uCxnQg5MMQq4Cre1s69/m
sUJyyK1FoeG8y1/XIKu/aH1GoRMh6d+C+mdnTht7vMkUEAvZOGT82T8YcvtFgZsq
kOm2YbCWXzcptnQMJElGmRKn6hEWKO24cpR3qAUdP1M0ihgwgD2kUIZw99Mimkvi
KQ6GJ0oV5gchStlZAzBkOClAPnEvSsp8yfmVBNEloMpvXw3JY+nT76sjoVpiFzMC
7Y+GxxyzdpwLFfVe31OhUchr/myQ8YovgY6gQcpDj8YQ5hHtpBCTa+RhQEwPvQRU
26x0hCwKcXXGqSXL1fY6cXnOfVqWg1E1WSFT/91HgQTs2WChiLvdfaH5+NoPNo54
A9/fW6Hhc5sPh7KMTk4ZHkxC2aouqI2T9K7STfrGigZenrpP/16d191zcA8DKRsX
Zrn/rnK/muoT/W9HW2m9QLHk/8mM9iMKvXvOghu1+/nkGZ6IYsdnJ6j6gxVqOQfT
WP6o7Husz7UwBCX0NDTDkqzZZHdUbNU/l3Coony9Jxq8pDkRuuoppUI3CfGRXYT5
JAUm19mAzkv41btJGInK74Pfpw379sjFNjQ/Y1lJWz9uueTMTIzjyZt/eHjelHRr
YZQVw4E38S5xXMjHkM0p4iCz72Klbp8SPyvY4DkxBK/THsVojUcjBg+dPEJZemLg
siqxTQqMCHqtH8W7EaB1n4DujDZX1AHTaDa6zWc7hS1WS8Pg7cjUANL7lyez2q7j
/oXgKwpVqyIgT2bAks3pQLz8g1jRhk5oyUvHRWyQVQpT8EG6nnqyeVGcmQn1ctA9
bD1A/sz8RbxOdZS5ISecmjoJAE5DW5en863G96ELb+Eq8lghLigcd6aSL4Uz73FM
RtvJ3xIpzUy2jY4wlMglrH4bys9GBKJvBChtLesn5ky9P47lJf+hN5Lp+er0i/MJ
swpmVfVMMGvkzibIbX2g0hRDjRGA4AlnzCTeYtkIJjvkgu6Adm5hXcHoxZh3Q4k3
bzrapyC0J146OBEI/QlZlMHTXVf51aDPmkD6v5laIHG/gZ1c5LQySsysdfq/ihvR
Z8sg5vbeYtlrtb7fXu4i2Pa/bkm3NtR1wZr7UmhJ0K4XnEHABzmDnyV7X6TSAkiW
O/BZPAcMsO01hCaSUk5DooonRh7+St9Dzm2+PSyKZGD0t+CIJjz+m2t+mLchqJGv
DDh256Vo5pFQW3lW48jLcnC7LtrLe2q8u3LlBrB60gquSUtS9xYUlg24MTYi8JKj
XWnJoWRXjHq4z8cAy7pPzltrHwFT/nyL0JtVvf+KL11MBLoln0lq/IyMv2UyQ9pa
Xoqa5PGqb14+SxcxzVA9excdaNxSaStmqYHfZ/Zw3WGYj0b5nIA4fD7xjNm9b4Tz
YwlNwL37zQ2YT2djm27BEco/8k3imLLjCLGIzoBw+MwF6LiLrGpCLgP0SCwfor7x
4H2YlSWmQIwJuz6HSNWACV2Jo5rX+711ifoPCpoSioJmIsj3IJXflLlc45P+twtX
vdKPxRtXRr5yQ1qVLIe2GfdC5JVMIF9yy43PttZ9cjoaO9xAvDGbtIPpAQo/8JQQ
ZxPka+W1Ja/Tp5t14CAo9M8P7GKtB98j41w8OuDrQlcgmb3lN8Nj+6N/qp44soIO
gwrGoo2JXTW51ZUTaSqgOpi7HCxL3i00ZrNR2Vz+CI0vbcQ5Z4yQnw8OnPHjLpKN
vC3cSocu14MkK0/hzxM1BVZdcC5VluSt81kgQEieqUWg879O3J3b1FgR6yVNiLRE
KwRvwxO2M9b0AccibZ1kblJ4UW7xctPaCA85l89WXr1A5FnPT/b097bYzSl3ucbV
cKo5yylBj4xzMKrrerqL9wi9vioXcVnX9tl6Ys7sUe6nXzM32cmeofRGy6uiXjv0
YqxHQtvHQaKTgiNF6106uYdXCCmiM1TobVtLgHhwGkqYQtwytu67vFV+XP3130h9
+qqcaqUgs/7oV/HxTJX/BaemAzeD5eKY9K/2Xwa8/SjMy72Q/1gl7D+Hy6Q1snqc
T/KTjWboLDDqM85FmeM+W4NPuJb2JC1qxJcxc/PLRYyorq7EwVPL+BeIK/7efOtM
abgaDEa0xlCeBaP9ymPtdKbe6NWC4SQ3Mu1FDt0dr3Ue4jd61IYkhwtH0DRqDrZf
QjD59MuoTMWuajG6Df3BqBO+Jui0vDE/Cg2H4OFzSU9f8igAwcZEETcBrbqNbTW5
yReD/ZhctKZMkOdKe9b8Bb36cIq5YF0rMMFMG7AEEHdMEej7XphD1UexSurLspn8
jxIvXXF2OyqgkDqmzrZK3l0zLCj4js7wzJWRq7N+471eB01VmGRcCNadOxicy/Q+
sx69ScEtqam33M9Bvyapt6okWeqRgiTUM2ZcImP3q6iS98mdwvZP9iuzoqjO8Z35
kewfa0wAfDC80k3/TN5eIy3YEKeC2r1+QonTI1+wBXzdr1/n/swJfPB2vrVbZWvh
O1ua/QTh2L8v27LMmCe8R50vOLcGgOGK9T1u8Tjj7QVy0yLNjWlyAD4TxviS92bS
uhuytTuGq+HosWPj6uJgvzvZ00KaUrfb7sCIhjuUWJI3rt/PaFAvXP+kTS/xyz47
vYz6wTmM82ig0RwFppYKq2LmN63vgN1cHFO8OU/zatRkbgxOU0kwakUQfApSbLvg
6NMXrBnYvh302L4Mlv0n1BARymbTwQW3V6BhRtsASDQPAFpYiJmUZ75tapVU9PQ+
0QNVl1rd1ELmnk/ybLeK0sUyeMW1upONkaWBcPiG7UsD/3E7AIuAE03+DM++N0Y4
p8Vh6ESogpDlTL1oeCNkHXQfBwcj7AnBNJhEjOmYRXvk2MUNsvMZhHKeC3XDLyFe
eBOCTOKcvEGCtXrp8jLZ0722kTt1Hi50ra5XWle5u3TtnPwGf1N4KmPm52lO8W5h
tvp0NYjp71SYYOnWis7NHNytrWH9j1F0K8OOg6ETDtbZWdwvS+fXa9y8xHmnXIAA
v/yWuYOFY+xzRTfTGoyeKAYPY6T7PTSzgupR04bZ6raSBXNfVNbkYKNTiT+8jTCF
fHjLh/l2BlSABO/0Sjc90a6iGCywcTeoKQ364QqSJQuo1kQVickz3WEC/CqClgXn
/QgUqpTlnTRXEkzy+y1OWW44QhA/UJ4lQIbXROSay75tpfhQ86zeKaLFgiLIXab7
CF3YVAnrihwluaIK+16eDAyMGVeaZv8829be7TiLpDiEvF67yjjp9O57Imu4Q/eB
lt5/gT84i3YE0+kw2H1kzYid3b4Xb0Gkb55ehGQhnrmeRtuKQEhTnGXH/b8q1JAI
25le1MAUOjLtN6ITp7yulyZXQuBEkjD3qlHiDafcfISJR2Hkj4zTjp9ETK2ImoKD
KvgRpOr6EpzQl4EejvtOkuW+v9R2L34KRPSnlHZqzzAeDVL0FrBvEqW/DawTUEfN
zpp+U6pcTHXM09Knh4kX+eriU3tfcApR6kYSvJ1MuGZauFzBbmEC32IAhkdIJ8vC
yaLVptMxwFWC5nFAbzqpYL3WMRlgwQl+xnUBy6/Rtx5Tn61BJO0MqVWgT8RgqZpq
qySOy/5BI42UHK6t4M/XVMLvClPdvFArN9W6voJGNUB/gKbUudxLjs/NRGNhJ/4x
Z05cVGh81QW/AyStQJIVdoFW7OxF79KGZ3/+bo7VHkpPGjTgs43uFYIfzagezSTe
+rvF4DdUirV8jCaECtr0/+eP8UMmFPo/V8IRqqv1HimfS8seSAiUgIHDxpW66ory
p32xRt3dGiETRh6PMdRu9yurFGY/0LHuk/Ss4dsMWaW1Fof+TL3MSgLB4B6Cxvfy
Bj+XEed8ioaV4ARq9Fppfdj8enGLH9T1fEMfvPrqg+pJ9JygH3H4Tr6cQx86me7A
SiowMIMx8lQrkaBhkhQ1L+0JF/z/SKj+FXQCe6VLHSjbTVOHDHtgVnr4C7E+HQwq
tkqDxTbWNXpuYhOYqb64p1Pmv6neBpGqhEMp1cTn4Sxjad9o/F0S5aTWrm14ORWO
bS4reWqem0oKp9a8+SPRjW1gGOyM1ezuwywr93Yc05X2aO+ip7cXgR3mlrQL9C6b
wRs29SDEl3+rhKy6RLSL7Y605iWth/4uKAFV2cQMJiy7m2oK6hq1JuFymxXJvsjm
sCETvfs4SKa2tQQ0SBvzOISQjXFuYYOsse/F12wIdxa6yhfBW4jwL2t2FGQev+dn
eUj32a147d5eU1rjCjU4ARDwNlZ6dcsGMSWTrX0uDFxuQcygF6GoiKqDqRnsFGZY
4ck5qaR20sraTn0ZXDY4JQnpZ9VJSnQgSLpOWTCZLQa8bxsNOw7PV04Jo1RK6ORp
Kb/aO3zwvl0MDdh5hFALMzUu8q6Z3wv3jhxe/JthCuD7L/8fba4q7gPVw9I3MDYZ
3tQxVjunBphtIWvZ5qFnG/FJPyke3Ye2HIYcGuKLYJKhw8rOIcsgdDulHIXk6kaD
kuDoI082wVT4r+uPcBmeHd/Uc3RA08ANMi4wg1dRWOUroHmjq26QNQa4Zwv8N5dO
DERQgwO6/ABgMsRU95udLhRYOeELmIls3KkxJOwee0fGFqO5/tc/oFq8WnaLGoud
RQ31NWVjdk2gZzs14PJ2tywcxpCIdGva+gXiUnWC42Mtg2DjdOQUjxWhCzfeiGAX
w3wcUvlgHwk7tf1f/bMo5MABr5CTC0FY+CrW4WnzcThzZXck/aOkf/V26wXFigL1
esHY6fCCJ49OmHCaTQZtcQ+34IZsKvIjyjZ8LyWtwyPy9dzCWplwiDBOvEK7Bkyv
1UYeA37kbPAmEtwSkatJvjeT27LR7lcGRR7vYtKX6kvwM9TXms5+P1mAH/BF5dt9
BBhmpQmZzjK/EgvCSLcdk58kaakn+MY4SFSX19NZwXlARsxqUMZlj6/lemFDEHOA
QmgT2zWgYwjZBCk9xzxz6IluEMoWlDsnFrPH9hUuALAYq6j0pfEHAKoorNx9eDwV
AuDV+DQ1PB4CUjy35KbUquQqmPjfWhcf7chSuhRE3pxNKNsBRKbBfzptMEh4dFH8
s3GVjz1PjPlrSCyKo7LNqMGoZ6HSHVgzz7E4RPUeGufNbJ297N+aOifhhnr2cKf+
NAUindN0+2cXYSr/IwQqkSKBWjwa4VV2P7/wMQn1fIsLZdbduKUPEJS2V+N71fSu
dRW2MkO6nm85E0ddYxRJ/Md4ASwer+lhgslZqsdwpWuhut631dY97o3g3j7NpMLC
sYcNNol0e7zKOOrzeKq6MnuwXX85xovgK9MhBWkZPygMXTExkVdNQMYavRFj5hsC
jdq71vSiVNpPADp6Xb2brwKwgZrE50HIFdsx5Sr9ABa6Ns0+non/b8mOf4vcHxL6
P/AR0Jb+dZn1ZQaQIehvLlIB+7I6F/h2s+vIwJwCGsVXOCC3j67l9Q0sThcyI8dy
1IE2upvv3+SW4uPCmWoydZ8fW8IvIMaHtr9LBtzaaOQ7LCkko2R65C0Sa9uO3n0i
UGhrVObbiQcb1zIgM/yNv39hu+Dfh2NESCmd1s8CddQsMcqLtbWRnUyQL3TfPw3j
xdCeswHb/ykWnfEm+rG/jDZvP43VCJ+azWXbu8IwegaXcKYQ+Qdu8ys1VsxZCgq3
VdJMlw3OUhfkAfcLL74o4fO5YCp1AbMJ3YHnB8w4Sozo0138X14HrNf6HLDZBkr1
xzxRN0G5LkLPXIjplkF/YRnzP8paSXGK2K8DavwOYYxjbtqLjxfP1w5v6dq/m/sO
SkNNMx2/zltUPG2C3gb7VAOFBmLV6ymrJ9qvqNz2pdM6/beD8q0ugjhrqcFLio0V
EDu3XDNAoHgUI+WKkhBwNOXEYXZkpEsgmusuEH1ZDaWXAOya6wm/MYA6L0lfUm5a
Zr7YIakJr0XDVyYMIWRyzDVdrgNeyPC2y8HEd8oebOSU4NNAxawdJlE3ZP3PGYAV
8NTxndvpgkrpO1dgh4bJH0jdetB0GSBHB4wIgbwNVH7791u+luChy0v1E/Evs57J
/QxRa9SVT/MYEH1fREMFoPVYUUN5ApOy7KTvmyyn0upfQckkrYS1R0bgymJ2V3oO
I+58kc7QASv0XQKBdVdLeFaVY9j2gG5EzvstPJHQd7cJGXaENiitIi1HV2MGSIOH
qgmVQDd26DaK9ItDtLIvGlJsp2blFaKgQ8n0OkUB8y3Mtm5v06HJ19qqGzZira+W
QWUFSaAYPM0h870nzYOHoM0nIBAhiYN0KGVrZa9E2hechSTbwzg8h2qW72nAIPhU
aQHWaVZirylvfF6/rC6vcA0GB95fdaLAdSjYRIpW9mPsGcv+NUmNVjb97etLFMzF
pqKIJrx7R2V2ZrIZLXb6PKJ6f/cwSfrgUo+Q2rbi2D9UeW2nxjomeNEPee7GONqC
tcJGxfQI0WpwJKT1ppGmlfA0kB78DNyP5Ts0uMBWbbMQLJmBOeoOBymxKea6ZJmN
FoIBIzY9DSJpVjPogvCsdpFReKv1td/PHbZDJ2f3VMUnANgHTd/NIpbJ7FPzSTQY
g6/SEh4coRxxq+HZ7p2spcLmAonlJ6uny6GylcuSYWByu70T3ncrThS1RsjSCdKM
oY2cpxRh+uGRuWhR2FWr2n3cQxuCEYTxWHfzyOKFFPZiKXyEoIcVT7Ru6bDVDfWM
qaAyKf6J5/u5qCURiTCAHu+vxD1zk6JrfhkXJFXrnDpBo9YiANGdkYOPR0sEfb4C
rjI9DuQEex2FSwdVCvr5lr3vIzPCCP0jtWIuz1tBWz/ICN5mGWH84GUTm5VZFcfB
N2dZIhS3WB4Q0a4kltTfZ3FkcIGYHZi/fvD1UHZycPxVpBxldDSZ6HYT67GZLr52
sAmHTNFSKl4HeIHCRn5Cp3ZkPYQ7ydtX2hqa3Join71ziDf8ma20vgX85Gh7vyVC
AIjZxDAtDqJrimYZUOZCSMNPHaMurBpxc39SzH9ciwHlXZ773MTqbV/JjbDom+rr
t7xOh78Hq6nxgeDhkw4wuNE7yNlTMY16vo6Xtj+XQ/7JmH9YA4ZxZfKmC5b33ON+
Das3fglYjisNDhZ7a0lGlqwaAuUe1cFkLclkoPKR5TYkgCs1T0R0o3clRU3OHam5
KaLr3mvXijpA8stEObc3SgAO5XD3bdd09Mm8yJ1zdZD2kWmsrtGraQg9u6MMcex8
peGzIyoGhJmK9s79ldX0KXOC+HgZePkPrAVNc8LrKQ+H2nf8G+b1gYA5/DWdctoK
3RQrdYuTZrFiFbrswLqlK3ZZQX6m8O29ljHMTgoPyMh4k/p20VghSfRnUw3rFf71
/V7+wtP7/wh81R3/kcyaO3E0SdKfG3CrPbKzTBC/fjEoECxIUb6Kn8EFEkJu7zUA
r95KCEWngwSsuEWShN5LN88bg8v4H76RDzOa6LhF87TjRWQhwZa24Y+BfICwDNtK
SZd4MrRuWgzOdakvE1+lI6tccSTyF01+DaKU2yTbn5xnt0LCq++IapbO5tO7giBD
cgAdQN0xoSn5uddCgTHepFDFjdpXrfZJkU/mRjQHBIxBjN+WafmHYVP4+3AO1hTL
OZuEqvXh6jy59GrvqbZ5Il1oF/b3L3P/yj5p8cSk44mFvAuiS9sddpnZF0eXAeFb
4jupckvARynemaEHHUbSkUXswJVftoKj4Qe/8RZvXcjzyrWze8Yrkjkd6sqnPhAL
Y+sF5IdIEsZYiP7Z7AVJ+Rs3e6qv4cdh372FbKVWaRbpmBHFMVlHnqAI8Sh/6m71
+vyym03wjSzj4K7JOp7z9iBU6dnQsnDoGh8UkLVwEhUhNJOPCmhceuGMwjouhzgB
NdicyhiwLkoHnOpa40wWQf+NIXpPChvBBwNe2hBDI/MwP8BLpmFLTM3KIODp+z7c
Zyf9q8vMULPxKBmNssiUcjP/uCSrddPxVGJpXIp8vB+0T+i/Iofr2JM/RxzLlkla
iG9AtclTlisSsIIvE4UIelTs2qtVBf0maAIPph7ncdyU/yHEOEwVaC+jeIUIfEqb
H/1wTLWAzwkVMdwbRx29Jox1HWSatDljb5vcRq2MM1tfeEHnL29QG3ErtoVbCjFT
ZAtc4ZoLKbjpwqg0ounktfkbEXaudu7qG7VH+3gqZ7UcqNQp34hJtyebsNvMiV3E
a5cbDC2bppsFVy7XEkWLfLClor8G/oZ1M/54ixDLsmNrWuybVTXU35iLJk/r11qH
3e6FImJf1ViYqxTYoe0AOp/lnvvQrUWvlSgFCX4L+g+4ETEqq6FneZMesW9E1Txq
dzIcOBcFNiJBqR+nOGawJaNoNimj6jNWCYdmflOzOQW0T6I/pndiBDcl9vsm0C/C
8PZwLAlC9QzNgURKjJqt7C0wslv6ZrUL8DZJbThZKJU+UgpKrhUe/be170kazfdE
5CpYTru4LGA7B3D264KKC0PIzEfFhOHAM+mH5snNh2i8MjbeWujOGSTxuqKXBfNh
8nSF7zDz0BHO+pzFM1kligIZjsmMCC8rLDsASeXholsixeaMxGXvB/cUawW5zfIw
sHOIQPOYU/zgkzFSSZWfKVaizlzTZtm5ejX2T9aeoD2ktCQDKZouhLgf9ZECJB93
ef6ctzrxS1UH32X4iInFNuBb998KL2Swyfb4gl8VZjmnpTaaGlfjOdOuTiDZYRZz
5QXvkpIEpE+Yup3seJovLfWnzunWbFHnuHZfSj+FguzC0Pr6vZTWV4li576ariWa
7mlQLFv4ix6M/DOUbiIxqqb4s63xzq7ndQmb1+0oQijUiuDT9WfZXBf7kvGXj1tC
ziIS871istMpvXOs1KHFWxO8ZvN0SfTW/G1leypEfDAWJ/EyzcnvFKv+N/fctziB
siJJn6bY4BTehGr8Yqh8XnzNyYfst0SbaU1nyqjcF1+apwzxT+vtLW7C0o+30Fka
5MGhumlNABgPX4OvZ46GNelK8CLvumjEn9OJJFb1VX0kLR2m5xpJdQBt38YF+jyX
Q9wYH+WfA8zjMW8uadS7ETK5yNnGKP3nvH9raaqZ3eE/Vp2k91z2XFpBJy7owf1I
gpB+k43JRNeEPV8XXxRUgbM2SQnooBaogeTxhmpwfttT/zUSo8mOSvZjDU7iHkEY
yxkbQmAj8dyxsqPXZkcCkZ19QCy6c5H22QoElncFNUpTJWU7RCIvVZ1F/KU5h6yB
aAZSaQnlDDWbH5drOaBVFocCjHhtTEiG8xRoUwqjSEba0VbWIr3DPTQoeT+dKZUX
FgcgCHAUuW2q/J04CsjVtJC7Z5uUBoDn1DXCq3lo5DzC/R7t3vaOLPkSunwkNIY1
AZRF0N6z2qxFDFr6AhV4kfeU7kFDbon6o76RIO/mCubc28x7SjN5a4iS2BTXEnDr
DcRKNFdFWfonywq3tgZpHZDOXr5zA9mdczqHM7Hyq4L6vCWJBnDTpcZ/7o+S5nZC
3cvEqD9tAmbpusfd+c0pOzmzjr7qDEZN3+Oks6D7dLf/DcHxq/7UN3wJKuI0fQux
g1Q/YNCR2UirpJX1E3Vy1Gi2aSRQRfaWdTweiIz4XDKXSIrs6tXw/fYfp1iUO0Ix
sBqNw5XJfThyJd9ID+pLUeN4bzOUm+vaVl/1rZm7wIr3AkoSCMLwY2/cWccntIhs
uIToMv3IX7hfUAhNI+y0PkB/blNnlz029MrMjb1BHvQXcxp7Ml3q2tW02YZj3zvz
l0e1/ubW+DBSpWjh2gYAU5w2xpuaUklYjHp8hcXGjn3mc3lEtVEo4jzKmgn+9P53
jewxvgekdiPaysdfxaLQhMakN+LT1mVxMNmvSSE6iZ3nQet4xWqCuzKp+E8tSvdJ
9gYRD4pdxd5Rm9S9iv8YzS58gHjelmp9VRrm2Pw7cf8ZmhpyJ1ZvIB7TfLbupAOa
n3r9XI4sjFXc2fQ6Q3OF1XSFd9gh0wMvA+9ANtQAUx3oXUSuCa5wfshUldfiv14y
baqkqlPgcsgJQv0MazVwzIPYn797RYqEHYJeU1AvDHyK+ArzBYK2FAlzbyFH8ePq
9C3aWyIsjhG3hw/Lsc1fony/CHf2scZHkdrNIv9oypZYkTrGB/xQ+i+ySzO+oKXf
8YT9bAdn9Szy5PepzwqhBXa2kH03Cta61WvoWWFpqJAld+zbTceRXhN6JaXJS3i2
i4O5I+kAFk3nOIxxfchaCEg8ly7KgSiXBAH/TpsTKkv7bO66DW6QCDzPe89/WfP/
i8PurDrXpshh+NoFyOblhoPGh04co7HxZGDmzgETvNwbIxcx5Yo3MaW/I4CMJBxo
9qS8BEt7GOyegCv+fbzVcq7gLkQJGsQJ2naVj6Gxn9+Jt8hoOYDiVB9ENAyNpHF+
2sLJhtS4OaYtW2pW1/5+PaH7D7VyiHaZXvME0FbRPOj7AfiCI4k+loFHZVFcUef9
iLFV5OXt+hniJYe2ldZSDoXbbGU8jrhzIWKD+SZgh85NGjJFcxD5peb7eOPsLPt0
DGd6QFP2bTXw/T+cyutZ6yKQlgDlSm+co9zwguAlfEvpzsTqHnJphtlpmuzYNkzz
1QE9TuVHd8bcac9m156gKj6NrZvjAQA6OY1Efu7VYGNgwtKZqbFKhF8qPx39ZzhJ
NvcyrklqSURHU9aYaJodNxJ/ckmfMBmsWp+4iMDB6fszWtWf5ouwLrQFkDCE5MJx
0BzndOeDoyC3WO45s5aEkYKBPa7zzDxtrzYX3Y32QFLzms4g1dAGlxVV18zCoRfN
APx9YFXWkUVg6Ud9l+Hx7GOGBtg0rFsq26PeiJe0BdqW5lTi0TD7lQmyNBgsbdVH
dLtpwX3F9/sQQIVjE8NOZoI9MWoz8WoQR73Jci0LD9ixsHR12F4qB6O2cmpfwTpS
1V9zNm/u7JvAdpXWbU5gfmaqfllKMOFVBWgPY68QdYALuIAbIIVvVeZm3q/cltdZ
rk1g/BGfKUgRex6UQmJEvtgQ89Y/eWwwQpsBbOvPDr/G/n8SEc+7Ezijz0q5ISHg
5fsRjZLEOl2EWmdD3G1iD7P9V+6C9zJSuiLZClDOjwnlOYhh0j1ciQk0mrK0oauV
FLaL34MSMFkgl6BnQfYy8IrsG47e5uDR/+iSvYmuuSF25/ACEfK+kWSx8xMUE2Yv
qh+DR7Il1IgnDDKQJPiVhqO1WuWAqAFJOXUAbXgj57sBLVVLbODKersancyWJ9CB
bMmkR8iI5CwzgQau6YqfkzcuYV57oV1V57ig3uukmVj15qSrj5mZOLj2Q5yY683I
e5/0jFfjBi+JUno7ePpARm4RA6+0jGtL4ESFRff1o1I3pLC1imO9ZfipFCCdsHgB
81zgbflrAAI4Z0AOfIf7ymD8qd5Q+D5So9INDA983ACiCPprPY6IiXSQcHW5cw+C
UiH6svu1pWxrC1tf5dH4JYcXv9P47s/UjQUBCPMqmlsO3ucO/JbmQHSkB72m2oV8
ba4nNPea1GCFM6YLUI3jPQNjAk1lu93IQ8UylaXLslaoL3X88lq4U5BYDSt4uh/r
elsGzc37jz4e8Wff4wo2RqAtUegeBvvXUA60KXe4GaLACxvxQpw512MSn3RdrMuE
Q4RLiUtIK8qLYtaY4KqHolXuzJMC7DoyWjPv1iSQxAem/5d/OI5XXFSy+4NCuPyc
pS4ZrJwRJKcPzO265uS9iNC0nQ7w1TksB487j/Jc5xaFZ6g1dF76MqbbUuNEOfV2
6FJ8dvFvyUq5z0y6VZweSxkzuRjsHUWiUYqGOoVO9K7C15ctxt1eAvahJvmhEWjN
1jAP+rx3QUGJ2WjN9qtGJTLkyp39yXCqM/ED2q3aHl6Jcl0QPHsgFMb/7/fq4scR
zWuHc5rhBEYE2G7nXRrbpVxSIAk46Nq0jRLa0zAungCbE89mhurx3CHofvMCKQpf
jd5yK+xL4D/PCtFu9JIcSzY9s1PGkWlSYk0/btMrr8Iwg9DeMdX/IHyqSz/d01JH
zO84aIzTJG/5nOxhg5tw4s2GEwuUXtblXEO/sdyzqToQyeuQc4sRfxq++FNISK2O
2WGIOK62z5cU3Dv0N6zdt0RZbXxTC8TYvI6l4VWrYc5wT/TkPPrXjgd0Xz6H9/sE
44ZuUigJPqbwHBJxkGOZm102T1OPvmp5RPzkOM4x+82dNs2DgVXypwIlBZb8cyUB
ly42tI6a+sMlQ1yZCx/YlCJZNl+L+4mAkTsU1A3KgkAPtjjmQfeRPfmPCjOSxVkz
r7e31dGOJyjlk/nkjLbCR07xJodXvgE7Q+Lr7HneQeFZ9Esy6fbnY89nFVzHUk88
7kCXFiJPLHNwz3YUgtPrg7c2MxKO/nOnsDjFcPfrCNA65rnBVv9VB6fT/sllYpMv
wlX/YfzHdh0d/46D36D6ETuYxjFxMO+F5jKqfcC4zeu7czj+8WtLOXyrUZHy/aUf
XoDhVqM9pwXDbCAbVL4OgrFkOsljvqoGTqGfJwzqZAgwtAoQL6mv7BcwA1Qriy9I
KYjgLjz4zN6VK0rJWs+NOsuM9az+AiwjQ7H/UggrgI+FFMX4VMDKE/Cq+I0Oh2eJ
AjGw3lELalOqIA+mE3accTUISk/7zKcxZyBOmfhrg7+5o9Fb1bXQc6szK+BqQVHI
8ZH+mbV5F3Z6WNJLH+raNqm7hnjdrqHlfWmYAIYTh5LgiCAUMSlnCJcmvEhhQprh
NNCTydM0lDWloLXSFUZzFKg9pwUnG/KBvRDhmaKuOohpsFIftqgcbp1xIlMOms73
cKJMBTFaYWCDpAHGgR1xZaTobiunGzzigbGB+HVGzTB4G/JbBcpz4rQ9j7tj74oe
USQsIKzEIMacgcitIhCsNkmHB/F5kMvAuX8ChpdTkThH/CBF/G5beSvS2NA/QZL/
v/7NqQO0cKagFMet2E1a8YXfV7u6Vf6hHhAB/dhIFr5KMFL03KnHu9WPp80a1vOo
pEHXiUo34Atz8qe72JQGN9udVcmo78e7VNUxBo9QSIH43+Cmf0vqv+SrodicSbJs
iGvOMAsMfo2xaxtDfoWPyZHq9XOPsAcINhiUsEejuMImbfAcmVmLGanBP2RDAmBt
WLpxyZwxZSbQ5PZuulw86ADaF6zDRRe9jAzv1aea1RKRJjpXXfN72+wEgY+hh3vA
j7ZI4iLjaZmvYOHokl/37JSioixbwqsqkE4HKuMM4ucPEg6TUKRcqGYxrk6RxkJM
wY8ccSkyoX/JeTguiZC6m/uyOsVDxoMzp1flxUg0G+7fXhewrFmbiQeVpPSdRtIb
8LnHN9lZM72Vj+Wd+olhIPi5pUuFAB1IDCQ3GB/TgyikDgS8xibdzYFZ2yXoY1vd
2HY3jYtyw2GYubrKK/2ogc9pjulJtxXl0DHQi5JqtgYPlC4FMPsSf3rndUJoW547
UbzdoPy/q4Da2Ebyrr5oulq0bqmwaxYeRIUwYMERJTTwxoxpZpfKQNS6TG8EWwFP
/ozeTohgNDxfuIw7E7uww4SN8omgNZIKZr26NZxujgnMIULsB/y2I6MRbdhKHE1M
PunN2fnJKjbrkhvO/F3olKa6YyKtsYx+xhDExANsZ1Sih9iiPPmqIG0oGQqZQ523
TPSVl4lWYYRU1yh3IMeQAetiqOi8RtLaF3bvle2Iw+aD11DyRd8v4JkMbMN0CIOy
e5gRmuU3Ho9TfmCZrf+2LFIgte38jgeHnmn3ayxwWH4ZxmfR2s9gIYivpBrLy3RF
Ve4222h7bXxea5Kd8IBgpEZwMHCngkksDoqnGTI1SgQfSjJQKY09sFkVKRUnFOuL
TOSQrem1/1WB0GhtyQua4DCEtbqn+8lnhmejV6MTHbugussKdasn8O5+n18C09sw
c/4spNF2f9SZevfZcKgIUagPElv7k3NpnEFCdxtiFQsyT0hImPdgjLaSHhy9FDIH
4S0lzAWA4ub1wuypl79/X05YnC0eZ89ezo5Km2p/09bNlNRzHAXC+XVZxzFz2eLv
tEH7KyWJBEKq8WAaa1uUObReu7C4sV4hNArzm17+xGMiKc3b+t12+oYawkHYE2io
GIyWjjIEkRiDVvX4P3nldeR52lumOSap/20Mz/SnPwFHk9LM6Nfg9L2KV+hu9htN
JGG36+tAN1d+mXDwSOVb++ZoYU3qxroDNLUQETNVAilZ+YtgpXBj/PNDL+OXOazJ
AppC7RJJ8JmGt+juRKPppTLuhS+Owfzf0LKLzv+s/mdXkGEVuu2L2MCfuUQsWGgM
TTSs5HIbPq0XXKkX7NoldYcjGGczbtiLZkt3deUo1jJZ/I4GAbqNUr9ZmLkMWLkd
ef0wuCILDe5YVGwIakUiIgj3jGDs/iHGGm8hXEDL4IvkYPjL6XM3DY6r7uBR6m+Z
LhXFmZ17T7p0I6mASLT6Vc67+kFYbE9ATxZZV9Q2Wjl6JUlVMAJTqZuSLepoh7Yy
4WT4N7y4D7A76rWPFuXS0Ny0j19N5R38MCtAR3XhCdjSTqLTauoaLpZShhD4duPI
OMvHhDqo5w+Il5kAyfp/uawk9IQ6LVBkVF+9VhIhdahb6LUBAr0VAE/t26hUTfi9
yEzzO7RxAHVJNEtGUe8BviJ39xhlxz4Vhst3nS4TIDJJ/AOFX22R91G5cNKShthK
NCn1nakbhRRVsf9fBcpnkLJiTVNmb8zozEm1mHgJOplXQpYO+JWIJwQbZQdkD5hB
Ibmo/0Cm0t0jRqOL8ya4h8f+T5Y25k4jZs4xKnTyk7tqWshM/lQvfOQU3Z7ZCkxV
C4tlQG4hpsJnw/Z9J7s2tge3Wp25h35HlcMZBtpGMOItHRv/cppWo+WgJzbWeaRr
zsvR6memcDbcIyHlEqArW/UsQCRQOBUSvEMQ4EnOjYD/x8szGM2/yHw1pDNOChdx
pdK6kmJob95AMchvm9MT0HbmjqRzPUNkuDCKZ2UROjzUDWQFMoiI4nppd1XjY9qz
H5MsD2WhFBVLS0ivSLnrlZgjgcdf+/Z/yB/vcUjLah/+JdjsrxFBGw50BnegH+Pb
Xc+wqA9QcG3odCxibN/RHJdksn9AtME6vZB+cafazJrhKi0sAc9xBMPKzMtHmBDs
TZCKKeaGFWezgbBJdkR1aAlwY0voCTEHv4uxxFU22xuht4Iv7pvdcOsy9mTIGfGh
QlnejLvcIvOIWtUAKd5P23MZZmZsmM7prI/jHoO9CwTyVEDxNotvJDaYMvPl+G3b
CI8XPrqRQ5KW1ZzOybRRqpfXpYeN3LVdi7e4hrnRZpAASNQkPcXTw67vBzXYvlhj
OB7UIZ2zv8yN0/iSvGF/BXIyT1dernoeLfl1lh9Utf5sqD/6gbwDU4Vt38EltCrK
yV//pIrU4jAHp8+I7KXKF87v/ZfSopVNXGbQvoo5fWwztl8WiG0ERFpJGNGyNkd4
MGyxDs2+a66Rn5YWnBo72bi90rE3Ru49IHlx2WJPiA4UcIoqZpkyrLa0NczC050X
nYiaX/BGXwYsvTDHsjBO6pbXq+SHfPrkt17BeftI7Y2a3/RaBmq6SjS/ra84wvHN
gU/Dg/Xj9iVDFBqlx4HdMiLbQD0XSBX/Ge1GAcFjzcvR8oATL/2VJXth8yiQcfiX
Pa9hmVj/JSVjGb9KUJcjv04eZR4jOzPQm6pHrGDDvYHi6FY7767UcO/uzOHaCRua
r4L0hDpcf/3jYXm5UkNVubmr03+LXwLLaF3gsXkP6Xi5l/OnY6icp+3sOu7L+VZa
nxQaDMEGUsIdJZ0fLjRkFQpLmf/yRiiK9dlYdYk+y1fINcdoddRoyM2CfMELfnlj
3LRfErWZXjcnzZ9eQiYUfmod8yvxwnLl7+taNOiK7YNWTGBL10nyJuLRpI/vQ/sp
VcaaCKSIEvaw8s4HQGwG4hM7fLKnkaAuEWXNrwvu4kzGoiH38C1jyB3D2xQIYDOB
yMSLdesf+BbHKKcV3nXjYe8Xwxlw9tMtqYI4jRr3QWGtMGzCCUdC/P/lTSadk++8
fnES6Eu/2d8s19HPmTHKhwDKTgLkcdhRYAT2G/md+32Cjca2VloWV5G7TOZ+tPkE
nhcxHQxiOEQhSq1z6gpQ3G62h4/xqfvf5g/BS/r3c80L5bMubcHQGUURoHRWhIM4
d5iRuAZxWKZdrJn9Y7MdtGTJ1b2t7bIcamsI7irNEEKWMiWrkTtqN9OJQQ3nKdJr
iaACY47gNcxErzXiC7JK8eS3LwZkEoBoPZJDhkucnsLKooVoDfLZCPAVJd3hEwKC
/mkx3BJ810feEQxRxyV1nBSmsK93LdfNm8oFGXgfJZgjJ0969QzQHjYPZ8B+oqf4
6eJzlJ3WiAxTbBRMEbjkmUnHLeC06VDNKx7gRkuGoaveWkP/fdVtj8mlOJdTKzvz
HB/8Y+PeyuYImM+pkBZkGPrHM1+jaZybCjxxRu8ofUyotBNZY/deFTucRbuWA8ui
dTd0mpAVYHLPIpGQiFcXojIu1+FFZNrZaVHKw+7fNV6lqB7fhi316oqh4n1CX3Ap
sFbx8eRqaqYDzZqMSirHwD3cYFgRLcRZh5EBZsylGpKcbKoFRIMy2NBaJ5KPdbS9
sFqvIUfn80z9daSywAKbnoUa9PTxro56BZPeCk6GiglrHfvZbS7zOHz2FLAL283o
/j18MrJg8aEN0ZGzwCFzT5p1XnPt8h6Pmlg89XQAsV9ow/UCKc8bXxJCGc+c9LGy
E8iMRe/Fx0gPwlE/yN7ujJjnEwUIBrMhG8SGHsrXRcc9gHc4FFZT8P/O/Dtjg0i1
0//b2v5hvABTLQ2ghboh2OtR8vJC7xbwevp1sW8KwK37u+Cx0/HJNnM78vdNHDL+
8MbCCY2F4MXfVcm2rMIg5py/3B3CQEMc4OYn3CTGKOzOno2FSe8cAFbc+vgWV2WL
jWFGJ5dSocKEAix2Tt2ir2hy/ikCLBG0hD6fuF6hO73U7MifuY8W7vqAu6pHQg4P
H+6KYqcEvTe4YfX8Sd5ZgmHRIRH0S6ue+bTTKV/OAhc1a/SXGvT/viN/Iku4jKp/
PTxJbdB2W09SueiAwQ+31RgR1pI5DTvINhcjRO00lsZe9RvA69UrM3LYL3TEzy8o
6aaM47E4rkT/QnQCC3n8K+4YWUvJX5ZD5B5Ryj4CggnZzVSRr1/W2lqWHXtyoAdj
fN1KNtZpom4vu0PCHtAh8TYqMnWDmuAYFyY4+Vp9DnrXkc5TQeQHUlLhqTziOO22
XguDV9Z5wzqJmhw11FGT6VO+szuBY71BfmemFCNdmQ6213iEos9qkudRLusLYEqU
cKRz0h6eKqiKcVTR5/Rx5RVZx0NgRz7rJMnU3nnTSajRUEga2VycnOM6SMhYxEoG
YotaFTX8gjJIzLjTmD8xvyRQgwOOaTiKUZKW8xHTg6pHgrYIWe/fuH2E8DGoYUcZ
D6Si5T3rmNnZha0IRp2ZX2TUDrkKTombJdvK5AYpqCZfffWLjhSR9wDxcak2U7yk
gOHOy7Q/6BNfqVSBRpbC0DsQzj06O3szY+e0oFp+6I4iZ3wxWWDmY6pPJPO2nds8
12ATY1Cg7vx/oMusTKrcll++JqYTecfTYrYu2iHqdaZyYjNWeaiNx4Z1XoQLnpNq
j8zzPCnIdFsCqrBdCBpg+7E1/Tw/CFvlPq2CqYYfrEulVx0Vwv9U/eRUuCzLaXPy
VxIwno+d1ArNEVKBBezOQlevj1WSacmXZH05Cr3yeYLbf6CIqJo0BjkDIFTwY4BT
Xkuhv7qef/+ChZWYrU3YF4FjUerqq4JSvD8Q0TOxredKed1u0KRWF/Yh9gKKRCJF
5MZjr7qKphdxDA5HApdIaKeE//bj7+IEr7Ri1+d3YraYjZ6EIpaUgkK1jPiOPMnO
Q3OAnyXyRelZn9QibqQyWEEzFck2/6eep5FKzNEwz3iOAxCFRPPSFE2ZgmJijbTH
mKgQYcnD1SvCUBF++wCPUCMrj5N94/eywoV9o3o+/wUu5qxGNopoMfCXq8mWFbSL
itqO1m0vkgTUr4K6uK9cPWSH6NCHyjHsULrtOoAShxgJG+7NQex8ek91v+OT2nUv
ny913OjhbD+YfHsiNfpm8N46v6PieRvhWn/ssa29K+iPs8c/vG4lW2YgVLh0527x
IOyZFPkNxHOgQj7rcTNV8tJ72uohunfDD6GB7OaRk28LdVz+d0b8yNRaJoldz97y
AjnqrHLn1YXTh0OfHLzIwigS8Sd0Rx00fdVzhCHCxt5gsprygrXrlqahCamLOI9X
KtpQVjghHjd1JEehVeribdN/aIQgN0clcxsr+z/0ozmSgJZzp3uWwhJg9pbgEJTV
I+fXIKl+qI2z1zSxLpRYoRb9Qgvi3ShMA3pURwwl09k/sQ3gDz9OJypxA8CsiqWk
oA298J/7qtjwJHLpEBIZUIgGyLdLsZZ9lC2JE8Ci0w4C/KVeaMZCXpR0cZcTjPPH
ol2PLJe6Fwd8qwAfUWA1sB4Jp79qMROjwfnXJvGCJR4gWFP8yWyxthPKCp5TPCAI
tiPE1HyCbTKjbN1b5HFfiS6fgmvHkODrXZQnXLkAHTsgSq6+wGbylmLyY4t/buWs
MSIOXao3ShhtTaqTd9Qe3w7pa1S/DnpzCKAgc6gvs7QgpvXfcwrCm+rtwRYEQdlr
5l6/sbOxalPXt/z8T13KvUU4Q3nHWHMLM/bdd8efe9gc76gVbUi9ZCzruIeCJODM
eCfYh9zBHnKZJHXdiBXbIN4Tvo2rW8zCzEmhGTvpSUVxz8K6IVZVIKAPN3m6jIfc
MH1Nth2V+SOM1xhBsNg7ia6oRtpXi5q8jAqRhpeRcfnXKKboGoxDC6mOsDH+10mM
z7NvsDlDGHdYJshTtvAb92f+yPlBnUpqxFmhWWo6uRo4ubmr85AqGWLqC1X7Pm6S
vqSlVt3UXM061B+0HuZURlYARhBDTrG24bWTB0TYJYk2CJitZHtun1C+mD+q2TQu
pUS8QAoXida9elPFwBl7AXX3Frb0Mht2vAciVpWMylfK1wLFtpS900g8JSEgmyRg
hhpwVsYnDS18GAd8E9nNC2zHIEbf+bkcQ2bT4sPojEO7+cJsdASqDljqFCSeMW6v
LJ3ktpWYN6iEzwrIxKdAE7K1TwzioB4aq4ZaWCV63pWXizvgK/ZbKi7Xixklij5M
XOGn8RorLbb8vrRzPtdgbWQQYe+EitHpaqfI+MjOc5il3aG+cubXW+w1HFhgBVgJ
3u4wKTALt+NwI4yc6/hsXQ63soNfTLYxvTX+VKzWN5+BfF0xtsdWI3i67Dg+yUi4
nohJOJMH5zC3r7nwfhQ7Ba+DG5moJ6zoTDeGtwzzm7G3QlsMbMShJtWEtf3T+jor
vvgk0AjwIFe5egJlrB8rxFbLaTwtZbcdjId7JReBGD6oXeCRP6pydlfcUcgIF1if
5RcDRhVQq5bljSchU4mAcrKqbzLi0pMyLIecftNPfYyFU+45uBfPee1bvA+qfKCH
1P1ER80Esx1KxfMKMxJmgnLuGmDjZ69Os0GdJJHmyxgtTFpdkAXxS5D1APqAZJy3
e7OyOCXLEvzjd49mSn62mRE3eFua4QBurH42nqukr0G/J/ciCdsvLf5Yul25XJsH
6E4LWd8Xh3P0bFFGDcDXNJt6tmFAfXTIPy4Q8/EU3zghNreKzRnuI1e7acO4+2fB
JtH93tYWvMKpLz+L/xtov1IANqzYwe3u8NZ5FLD6rO7veUshulS1GDWBlq/j7DOp
i8Tiuzn7QjPVhR/Yr5JbzhcsGifqFrVwpppBkyd8E9dycYeB5j8+nkK6fHgnvZko
CITSiUzLOjP+aB4iDtK3kv3J/3bIhO4CmEpjcBBFPbBRagfjIT2t9Rv+x8sCoG9Y
ARIFXcdYvl1NNQHya7U95OFhDytCBrs8TRcJQBjiy5O7QDW1ywBAtYi97opwsEhE
b3toI+bj+sKFImC637gwPmM9u5eeCyeB2yIGcb1j+BEfAkvietezku6xZAIdq+YU
3x6uf0Ib1xx3qhtugfogpol9pUwhPU6PYb6k1RiZVeyUn+G4FeaThZ9K0d8gfrk2
wQxHraB+Ao7Bv0I1rrgIGwc0cbyEsbTuQ8dm3wbV6diU/ZYVuI62hF3u8NUs22nl
mkLYMLbcclwvmFudzNVigDdTxHgDfM+O0gdpZ0VWHzk+6NmZzNIcsSlUujaNevWC
Py55IXgKJlt6V8b2f5kwmo0Ylo/0uP46bm2fQ8xPzUguYhGnmB1fxaDGLOiFL79r
/yncRg89v2AAA+RxUNC/CB0tUdi7krKXeXHcBtmphzTnfMwV7I/hsqBjnYUO/0KE
0oA/jZdpXfBNqQs88isGZ6YrmsJhpc4699lV9nW98xXgDrGasLEB9731Y+6sRoLx
H2YNLb3bp4vZFHjrmcQFEh/pGEIKPqBB8+87K2JaY+Htmt+wXsjGufXRgDjoIn9+
1CgVbXAamKIzFo5shcBruOtG8UMJ8Gn61/4JANHGZOKzh0DEFVfQfg4dYwJWru4k
EqQSPbQ/DMSdl8OB3ViMukxuzOH9btzDzJV9LFdmBAHUlYIq6y1kyNTE7d9S8gft
g3xbXYWMEvz3rCS5QUWi8l2OwWBV6N3nKBLWxDYuGsT4+R9zYN+S4WFpg1X97/xo
kDwNrDBI/e4hrlykfjXwOYU47fQLAP+tvgzcuM8nLWjJOgalf92cQ5ikDV/p87wD
wyXZKcuVCrtFi4tNqmpyDVtmkfsSZDMqIxBuG+gR4n+PD0MTnixZJ73qTadZW9lM
bTz12sKjRLtwyMXDAcQXftReezE1TvnJ/czd7r3oSlx1E2JzRZqk+WKM9fOw//2W
qKS4vRNee6ksiUKnbRCanw5pvjVv7YSWXm+3CZT0Chh4BetCgUSENxJWyM6ea2Vz
rjmRxcyZyUbX48p9qlq6rYEzdoHPrvnnL82y+sd1HrG0t2puLD252NLB7H6CXeWX
LZSk2Vgo4iUhA9V7m7A/aElUfC6PwkRpJfz3T8Ytn9SJiSaDNAKbyvNY9+VQzZDz
C2IBq501Ar/ApNq5fl2E43we6WK+E742vNgtlQSjIBkC93n1vfbdFcIRNIkwgyP8
ulTd/d8kYmevaPd/D/cT5qFNTw4kXmlEqhwf5Q82WAaHMpkXU8jojd38dg8nLTEw
bGlianFGEqEGuoG5GO4PpPCLnvLb59ROxSkdGwf+wVviGk69BEszS20IHGswbsCn
RJJHH6UC7XfglkVAETncmM4P4gaXT21vOtmAdYaOKUz9QzNDSyLayMIpz7PiYJ/L
FoA6CNXSQViMuRK3sud7PEgEsV8DEaw0mfGA0gdjbMTuYlBhQ0/8+7HZGAcY/CXt
FfCnoxQIhOnYhFZeAH0xqx7B7Bu73Qa+VY08YCF6HNHbW9o45MPTCzjiGmZ9ob6o
Ce/OXyVYKFK2w9kWMAVCb23xxPFPF2TRWcL6CbFnH4rV7TigtCu6xWyXWsh4GhV2
CU9jOQre09ClQiD/g2TpXTT17ZmAG59sgaULZbRHk7B1y0typ8B1xo+4BGB2a5zn
iBs80U3WoO++YfVt9Q07xMdOSTkb3XaZOwIoPCc3v/F4nqvuA30v2Er4Ndd2ezp2
sN94dAwBJYbtBos6/Qi8tSXhXafkGcuOj2xUBI6OJstc2RtxinxLqfjz/4EoCgLv
q5mLXCrDcprUC89VzwSJcvP5fP5kMKuUCRtEiSTbC5OQe7rF+LC21gsPjIndbsx7
6C2CH79E+TYTTuPr/4+o/8ksiMECaSZ3dr/dbm6meS9+6nEBoktg4Q5M8Kd1kFYn
O2d3NikdOMnrzCTydrYCvTG7hrNqrdeBwyMEG8LgrkbyDmoQL/pO7N9Y5l8Usm6T
ag4cSKWKJ9z4UBFQxcJI814tYWISVMi4LezXQGelzzQ+yLtJ7hWgzS+bWYkD3+85
nHmnuJRHqVZF7iPZ/hHV10iSWGnYuOda6NssemIP1T8/frKoPayTEfnUnGU9cqhv
bhnDw45PnF2TMX05G8DLe5pY1a2I6qw9gOUpKtuFKMZLaMQMcDCweJuFFcEORVXV
i+Xb3LybA3vBojqeYB3c8eVprloanypRhjTSTWk/DZnRDU8+nbURRgo2SIH2hC2F
yuR6v64eG20iqRph0icHf+LQkS8bIGYkOun4cR1KqrRp78tiKuH2THd2S6GxfnWK
2FWH7S1NIpKcGuSOEmipN1Hawhd2Q2Dm6TRF8JKEJ+MALCU+8vD+BNIVIaYw9vB1
nMB7O1cih5S6eMDuwC1IUEgv5uRN+FyqOg708xNlg8ynM/Yl2dTbty3lvX+822rz
ESS4mxiTZtBqKJo2zPvxqidO4g2GhOUEddheBeRqnWpLvGggbPSlOlGxOCPHwt7L
sPJyq3/QqPp2ee2uBmFCfso23xbng7NDKlGJUqTTy6k7qZMfRjEqnVE/XUFRF/qX
/vR8tKyXVSP2hgp453Z9YzyJxFi9OYpSXgV51Zp4TsiELMjYJS37XxSxdbDXezGD
jEeqgyiAdj5GpIWqiTH18lU0VGKcBcs2+HBk6mM/0TNsXS15Vv/YGZZ0mOuRhfh5
VX7B2aSKLls3BelCxVwoveE0UQLuNUx1HczsfX9kB6G/Sp3EMR6VQziJXACBB87a
hDh8Ihufi/f1KGnNccNfVJsvO6urMepm1I3pemRms++xhTTsNcszBt0auKPwMZjZ
YkjSI9WC9tw7KlbGYkerrmuAS8Ju3Sbewp6Tnu3kwPqM99Sc4UiTeSP/ZLXW+A0M
Dhd0eXrlsz6xelpZWb88MWAuXcu9WTMW0Ejkpq5SoacFnUEv/U58caaxfmDnSB8L
NSWEUTTYNh4sh/Dc8uAi5LveGgu68ynBQ2ust8QAhJlq+1yVlzxFSwoXCIuVROmM
u029kpNEa+bx/vp6d0y1z8x3xz7UqaUs0mo56FIS9CD51beQ09yKYtYywyaRsus0
hf5JQSZhJAaJDwb69xMSez/v0P9AtQ0IFgCkVpJVJ/zr+Da+5Uez8e2vPDdW1Rbz
BL5c9TFn7vpnyCeDGAyZ651hl525cyqERv42w4EbXsPGmc45GlC8OzF3VNOg4C9S
d9IWoFHAwDFmtU4+70NUJIVnY7iZHrqfB+ZLBogFXLp61r4bP7i2AmbGz9M3V538
eMgJHYxTqV4bwGRhm+Vxp70vezF2cpAXs9j5/2WXGssUQkZG6cafTk+uI20IyEBm
dVqTdSNpC5p+cmL0DVSTxxcq0D+uEHBGM6XnO+CKPhqEWa7slnnv1FbkFXasHlUq
A7cqzvg9SfJeUTadyGN/ofgsQPaCo84jVKL51++6+ANAqO2ifvHxeSh05BesawAx
DyM0wKDGM+jomtTo+mNR5lKCqIXW37WC8yQ65S6zUcVI8aT1j43yTq3/wRcj7JJR
w8McYCDQC7oBOlYGhVsB+uU+42JgYCtU5osJ0AEaslMEJ3iacP7bp2mSsKSioiqU
PXiB9hu/poR2swtoTCeovacndcccPpt76chXLIydF5O3aEEnCzxWpJN9MYeuADQM
kuolqz2fo+MvBXAhoqQst2SYkBCVKFdB6wMqgoJ7eKkMM8rwafJZdkQU3RBHfEn8
9kSUHR220U6oaubpUyMpWOLfE7/laS9RX0mt8abzV0wG1EwBLiZgcdKWVPWKVqUH
c800x08qFJRkMTY63nZ3jtjgXZxEp2u+AKB5pQupnW8doL7ys+fiOan3/qCpHOua
U893QEDGlOB5mC7cNuvLWWmADRxxF+wzx0aGM04LikCbCX2GbJsahRdVPAMJSLBK
8UpHCUzRHcAYiY0DpDqD8wEXFYBtVb4XpYHW5YTXior/A83LvQjMlfK2oWSN+tfa
WsHKvPhOd1mGMyNR5GbbG1Fq9iQ6udpBSdPVHzmpWQ2qtUNdZA8pLRq8jalwvpW4
Ao5GUH/lVy2GDOjaQeX8E7dzU+XFcRO/rt9ab0KlNFrQI5D0OxXpcHDHyLceERUe
XLPc0VnkajKoHBWzcki4QAYDOtNQ94JC9Zjl13B928sGtEjWYy7Bb1qDWbePzNMt
JhHc3cvcjcaq8cjjXZd/K6/kqI/6aHPooxya7oZMShlkO8qRyfjiuGh6zAFW6WLU
hpcl68LiXcbp7DRs8Of912K7gyMe2Je9xfpuwuZaRRLIkIK9dcGW7nlgxjRaJ3An
RoPJ+Nxqz3MK6KDYRaxj9fIYyhCTXrVzHLDaVefg64rC9G/OLhXdWZ4yfiGYBpML
9yHfjQNM17FSNWqe2CjJ8OQ2tNXf+FjXQKQHurvcgd71xeBNQhGnYFIZvR5NpMqd
I6xH8bFSIB1hY3/v7bcdFQyhtvG3fwHNXJw9DpHCtpR1zJhxYGJAlolPOJBuCVpe
jwVyTujTtUNv1NrMPyMqOv7R48XUC9Z8qK4MpMmnyln0WqI3k/9YNVJ3l0nclWKI
MElXDXPVDGlSsuOnLOfXT+ctoAKy222H1Vw+EORAp8//96PRO7vEib9zqbPPs7zl
c6p3+Un0ldAjL7nXG0M8cZPNHdrPxIxbpir4CyVzZL3lBr2V6K9NR8RNAiyVE8bv
/akHdo1gad/R1/y3m2X5Tz7PWDNsuPajjNwVcHAaqfv8vCYIloqe5FR6fFyUyDAz
cIe13eTnsVBpFRnxgkx6QTsExeiYZIAcATqQHM7Xt7KPT8E1ZyaQrfdPwcIR/Y9a
JCVuZ8gQj37xM+pAFrQfPIYW2ZIz6nb4qEDzOdfI9Gaq5wBJe9XQxlbNUhm/x0/i
d+5DCahom0yCSzM3A7qdGCbw3qSht13S/toPGIRtzA3jgupBvOWI2DwG/DL0aD8Y
cUQda4AGk6Ldr5idxXlua08FOSt5SDAwGZZyweOTkBwKf7DX4Ns2kHAgZr7y5nde
Iaf5NSGlTqsaj+AX1kQUSDQtotLWiXihoPq7eANTU9ZGPBFSYhtbbPRSq2i7hVR5
BHwcz0TGh1Gs7B6urPG+jK1Bd1Z8THta14jDZUfs1/G8CqBceMvmbgmC94O9K9f8
k0LR+Z1TwbFHp1B2Vc1OFlorW6tkMOQ04KWjNm89udNMnt+Ua85vPglE3kf3FqCS
SLnzFC/Ki9aUuQaFM//+16vWKD62SOrzwg/qjPkEZ/v1NSGci+eI11OD0gK6nMaA
LDJOBEWl68dngA2JZ0PUbOJFyqFYDzukoS+Rvf6HhS4E4oiC3pOaUNT4zYZ0sJyD
L0bs7cUYLwTbVX/bAgWsiXqewg6ws+4vNkkbdAgVhjL7mjjzH1F7KKI3KRvixdnk
rkrOqcSoXZmepmZLcymkIRruCGeBP1okWUfMxv3ULF6iOSZfC7UOiqcuA4IjCVUD
squgmfTNAf7Ozp/Xj5nOhBhPJ1nNlRIw1PPjVWF9ZNwPo9+9LCKgt4x0B9ETYiPg
fAdJhBiZTr7ZD6KzSrCwzEMLF/1ycVIs3n3LNvtRgJWQIwJRUOyNh3BBklJfzUqA
c8wilGdznvEzCh04LRLN2d+vrmGh24wLyZmJCtf4EOpS2Wu0t2isgYP3AqjnJvnb
TmzJIQ63mwjY37r9HakSjOJH4CivxPKyatYpMRF+I66JUdsAEel5rBwhuW06HofF
IwCw38uedUfya8J1TuXgPB6aFm8rqwF5OQ5PSbLm9MWZplMuX1k+jPIVsk76Vvg8
+UZyVMIXS7bfwd+H9yyK+YiMDaAX3F71PpMci6E6ntKyauzEZNE0s15bMfwge3Gu
0uqOezrGB52CZGty/C3dVTcJbadK5KB214kkzFWMRXbhA8p7fc7NsEGE9OqszP/Q
p4TkuKnQntduL1peJC8S1Eah1XUVVWBTKWyaWqVxqSmBdU1o3I0fdCq1RV180k2Z
dweKLy5xIrmTEytuDusgkJnOMe8GCz44yiRpFc0uBuion9uCEeMQggPTvDTXqbu2
suNrbjCyLnF1RVyRgx2x8bl1ivTpbgJWxgE45dJVVW+dZDEyOCgYHtfp5e4sJHF4
Fu1KuoZCSmv9Z0luZTOrGf9Y/xBeZ44uXtSB8ddcedYIDn84f2myFWrhFTOZfEUV
uXamLI6PHRxT16S7MynyzCTJcf0Le+OUvwqQEJQ4+Bm2DfdmKg5B9+4efJ33M6YN
6G4VGVmKtHKNIfXcmVOwgszNfUbvp6Xemr/MduMrcCIXH2xbCnJYMmmOO2RTWe3c
oZ+6Iw2G+3vm2BLpUbDH7EFySUCFBweUMV3Dm6Qvcg3EsHf4DBRBb3Yi4OV1/qBg
X1tvrkD3eUYQahjlaZFfx34xF24fLrDCrVf+fxDrHYppaJlooQZUkAnww+vZAKl8
GkzIGCrp9yYOexDuBgKtBPTWfpERs+bOiUHBVlj3lESQZYgPaRPcD197gKY10fXm
zAWWZXHA3ydD1AI/d6Txp7UcamJpfpd2BjjUdwfZj1sNfW90rm2ql0Rx5caAxJTn
kAt8RrzEnwgMlaCyfuOjwJBgf8IhyEeDO+vY6JNv8R/QMEKhpJNd/oZNIYOvju2n
to3hfeC/80NgcQhHUWcN44m4i5YmRGUKxIwZgnMJmYh8ioiwHowVjIQ69cgcaQGQ
KPkIQHtN8TqgYgR4qSk4UltnIlgPeAxO5hIo1+hbI0/IGzAqK91Kw48v76JdjIlK
YcF4jR2569D3XS7YSzrw/znW+A0sv8mzYNbPxFp+fm4qw4+7bCB3IGErPcFF1UAr
r7P4Lch8mVZzD5G8VYa3R7mDS+KuSm50+z0M3lYoDTkz3dPSWZImimtFRP5tuVyU
6GCydTDpjDlZaVGUBc0eSEc0Hh/F3gBEYaQUgIyIZKGjh69et8Zk+wUIqlLd0MUs
1nalvBJdGstRVhGU7K3o+yTG/DiV6U9a0EOkFUncDTRrIihmPur0UVHxkVfZW1Yh
qf3Ft/GSGrsa8XsJy0Q3bmAyxtlNWNx9hR5UsfNei/WFZacxzcuX8OZge0vhcBaK
9feQfm7iQoEPVnyAJYk+c2jLY+78U6ivvRtHjm3vFHfu19lxxFvu/6TCoPV/oNVT
kHb0ebSO5y8k9D+KaF0CkkFbHqA5kU0DCaBYuUqgfgcvDNLlvKzCJ8TAz0YgoRr3
QZK3hgu4VIAmbrGprPXvNZhk7X11uG0GFrxFBMERIi2M1PcULeYhqR3hxZV9HJ6o
QyzUgeKp9vsQPPaEqa8UfT8pkaazpaSOtwZ94kXHNI82pnum8Af1cyc4nGQBwB7m
kprzWpdnBMKC0ymU/fLJILcknZnDWAstCM9mKoj9/DPYONkV+hVog27xtROATsPU
0Cm8u6Rr+bvSuSPZxvdbmyPi296Pe/k7CJ/Xf1xg9GGIix2Q0YE8YM3QfXzLpXgE
1GzW6t/rCm9CO+DmkwKw8Lpo5/yXWofrLIH98rNAkEd/o5+h4d5stDwE2vH4rNQL
n32zM3rOReqnvQxwvja4PwMt1ESMbircNAhhjKFMxtI0qV6Qk7+r7MPTfm8+ossl
WXR8cMINs8b8GcXP99bChBYZmisfjfmqaK/b2kQcGB9D+GpFVQ0rKJMhetdNGVQI
scQdeXAz13jvpljlDlLAPr3LB6LvGEfQfWEp8heQdUvF8CvjcXTmQ8ISQCxyomtn
hfisD4AD0I9sf15tcdj1LhI2jmyxjtNTf36IjxMgPVQnbsjnXfWFf5a8ZKFXwAhI
8cTAQl6I+eW4+q6fNTEJtxj/j6zGZfiBX3JaILpR4Gva1McHpD7YHGg7TyxotMnT
Js7ic+dMDJaO6Y4D99+2UjtBCYZh3kmXSzUwXK1Dgq6q+k0XTgMyP0DIrzN0Wccg
8ceRNQWIwCvEbYNyHtgZooq7tdphmbkBOzUv6rJQYdWNa9dO5JsqpfQ+lHkan+di
KdJZG7sKK76VGa7X6eV4dTKSHSFza8SNUGFpFFzfF/+SX1OMo+EjM2l3JFQ+tsY0
cT9YShmH/aOfYWKEYqsByQ8L8LSDkgRxoi0SUoNwTftqvUQ6GDwDEaJYBFHDEUbN
TX6L5DB5a27ODNd4GRSqAXTOZ/wKhHbH8nz8xIz7QzuyE1jCFPLuuZb0x91FiqFK
T33iJEpYRhfIZHqp7+kt07Hivtbk4p825rzFvSlsV7CsOj0Vpv1qup2iM5yQ8Ng8
FB621mHrS0y4yBR43bKH7rHa+53pigqlpLvuE/m5OHWsuFxDR04FwDz6j3Ala+YM
VsbEBBw3eo/ma7tQutaDjcjFuV8mfX/Uivp9lNYakXNabTbiU4JlE1PODrDse4OC
/j0hoOkTUKfsUyR5d49EpAoc4PPX285zqkPYwwgqeiH5ACe9lnQx280i+hZcAajI
SNEu0BxTGpgqxYaRsZbuqO3LKrxv2LBrb+pn9i6Yo2iDrwoy7pjyEHxm3IPW6Ho0
on55NKq5wzo9sTvU0RLnYUwGUFQmBIH7P3GzjrfX07jPHeU3VE3Xc0nKqQ3zmOTx
mvqQuh0+igFk/PtoQVMRMV6U7R+/cUJGeP5NPgP26olr915gkrggUyydyuVnm0AI
hqoKqyEuc1tzM+H6VwEXGE5e4+ug4Shhv4v7XaiYpQJYqMjblWdQaXvJKafYhrkS
uWo/6aHyru4u37kJxJrCG8kaZmVEwNGHe+rEmxrlOaUHzczA/jOdP+iB6IBPCrkl
ZmPTEccKIt3MPMceb1HTHSuIy7iw+wYGEuqH3yw/zHZ/lLLmGKAqSQ2IQ6siGSPr
QLQ98wVbmCKbuHag3N9+hGAIVIquNRCOwg7vZhrOBc/1kg1zPzw4NVnAp9lkeRGA
mzN5HZ3xQBem+2YtXRrLZ113JjdUL80FqZ6j+poxzKrFjjTsj2rqATx/aiPeFgjc
cWcNPwpSu7Q8T9rD1EyitFvyLlfAnn2EDVHmJ8Cl0zUhrvzZJRWtTt+Fba3ss+BJ
ykIhQaqWze0mCWlLPeHcW4Dtjnm8OC9grv7sLMrUjkc+NpVin6FrRsnXuaGuPrWB
2AFgxv4jzSYzZAOimX9fhI2Yu2tY1+9eUOVuu/DP8L+igHWxB1mKG3borHFLajXb
xemtL0Id05Pnd/IowyPsdc6wEt2L1SkpdF9Je1OzMnSgElV6udvMys6GlhA6WMP5
luc25JvX3V19tKReoPERt7qlHycVDlk5Crf9dYCLMrpSHjizEvMIB455PNJRxFl7
S9wVULSTmijO0JKj6BgJSdX4vT5bo+MrJAxvZi1DOFheIqemLWd0aw5dTpmMbE9L
46RK0hqggNp6iSypVBrtNFYBtpWJBx4Gt+THkYdpddfsGwiCNHDhpqR3Gd+Wv8+b
ZdRGu/ph+ZBGWwRNpxu73hDSrHHrMadbM5rCnHL5ERtF29LdJITqjmKUZ/mVfcVY
CXJmpRaY0n1mJ3Rt7T9fHyePv/rFUJCq1ggUAYNAoiZQypxY4M2Zv0qIuuvzmvRi
TcE10q2H37EXAd3CNkonPL4KiQn2zN4eufo3z7u1ZgX+W78a+9Y4+7zPYulJtfYp
SPgHy8pZEPhTY5XAycPPaTJQhwhaUzLHfzmSPih2rYY1vcK94PhjZtUFkOSqb++j
ofKldP/aqjo1e0GLLwh6cgWtqfa5niJy4Jhm2PSP7Bmrc8L0qvCXkru4RJo9bGhT
gtRHCb4p9ICnsZ/8bhY+g1tURPQ0F7lmcQZAhxEZOe5/m7ih/J34nwaTpuLaFiTF
DfXC2+TvBX83V775CUBOSuD0VsXHggbyYjpWgeFOYpZNzZmra87C1eNuDZsPKHX8
IBicqUsAzfz1SDu3SfEG7PKU2IF3vyxEafTsqj5nuVJ3q3wSwY/CQN4lj6mSs2YB
+HwtI4npRhKdONtAKz8atGWSBZoTyiloLbqEWMzhwIHqzLMtuEC0EjNi3x/PwaZy
xbCKlSYjj3Y6xtoZzq/vYtIImWSsuX1sOP9zZsvwDX7/x2evvWTJnRkdElTANzUv
ny5YJN8RGPeFWH9NRa8sNscqV66Ym8strhBXC09IOtxL6vEN++uLYu0raALLPien
FQI8pomHHIP9VMmcJxmNHI/o/PkY9qQ/2MMdvq2IRhoCesn4e/ADq0+xyQkQDxLi
x6OoYpwOi6K3ZTfq1mEsX+obC09jYzllE+s7zTYN+v2DzVMQIg9cvnyKq3lDb1SQ
08nXeR09NwkZVwsapGgU0cHBUNYI3/Qx/JueX+aRhxkdYPeQOQ7iU+8FM/P9StV9
4R8abn4KT6GsULWcmmtZRw9UvgaH13c537dCEJmBArzsmNTW07lhYLJ0GOaOBIX9
//7bevWKQHCB4ywo030VmdApD8zs4eHUGV2KDDt/5SwakvuJmg3bdCAJ8A+ah81u
xsHeChw7FZfyiVAy+nEqOwZyBSKeiwSO8KRJrEtOZ3gtGDflAyLc12rhZJDxl5uS
qd3qdLQ2MG+uf5sXopzoh92UBSMIQLzqdPN78Alpj6fQ1Pu5AsNHzampdgPJD/wE
kG6BGszAt/0aMR2G3B53uSGXBna576+G+MBhnj3roy68q4TNWeVRNn0pr0pCJDhI
utFxzUmfrUKgC0NJogybLFZDQ7VCRVMbs+TZfGACARzMO902WzKBsbSXlqZttkJh
mK7GVRjFuWqYiw2FCl3eP/TnLPA6EgTyXhYOjD1osg282QYK3EpmlAbnmxevOz4n
XW4FQTop4nQFC5TrtByp/tDdH3jLS7OQD1QlqcqEr3Nx9PL9aRqxPV3YNlz4I4xh
YvVcB0/40qFaMZg96VtboxqON3tWw1/2uJLzyeKwlQppi8uXdNCPWqs+Lgw7W1Jp
jjH7ASCCDCh9Tg0o5+AZGz20f03Iv7/87xnE4/VvVTE=

`pragma protect end_protected
