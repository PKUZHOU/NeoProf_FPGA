`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
DCoPYLxZUA3H2jttPRuRbjx1hUizi/RN9KEq57z9hm0IhR8QJufNkCN/JpHthunO
i5gLINfgkzn4oeNoVwIsnNriXaZJCFGPmChxmbgUCfBWZyrBP33VGBbrpB6m0bLW
xjg/aIMCZh/jLaXHBUc7fHQxPYPBejIzTy4yn1XBUMo=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 8576), data_block
Hsr4Bo0C4bkCvvDSg1KodEZuCK6uePtxBydXtew7g4AB4GO4ENukBwyrV9+30YrZ
7afH2hQ81DOWXQer7+MK6kNkqy3JezvagYnoL2EwwwHZNNLjk1WGBZSVTDAvH2eX
B/Pj7g4Hib6kjyNujD/hMESlvMBU7To4Ey937PbWGGuiu05zzmKMT/yhYqwajsU2
7QmcgVeAbKbnTDkpYih5WPXbj6/C2s1k8m7r08h2KfP17C55AOIRtp7xPrgYBwlA
1QZ/KZke2gD5cJAZyvRJWOOCf7+C9LYas7GQmnWW0j+5Eip15dfpd9Xn/ZV1aWht
OyXpcR6hnIQ9Lj8JlQ/AurkeesMzbvFqfhXVsQOLRpDT1gzCOO7f985SWE2tXIqO
zwIo/ksBUOy1Zxuvp+LGL8T+yb1a9DGa9/VQzbRGGp8Cyo1JW9Fl6hdpWwtw+D8J
KIZiqM4oK6dTrN7K59uwgCy2MJr4wwdsG2sxXs81nL65MTdX9gAbtKa1lsMTZ8BU
7/mNpB4Dk7edTSIH7Ro+g38FSsoLGQG2PKh9EEC/wm4WspCw311HFwn3Mx1nO2QJ
aR+Fwhh5yFZpkjA6NMZkkvg/LVp1/HUjGSEqhCNvMSxQcRjOIC3Zz0sgxeuscfpY
CO4+/II3HVlddvM3m/FJWMnjVortwgu7WpEPTfk2/deECOz8qvnhIS9sb4Iyyzhc
RztMEMBxMgoW2/Jlk4vi9j/M4AAa4VNeknRKF9D/MsznEu3bE8IxvpQxOv2V/9kR
LfQfJAvUSSrbkhBDV7TLF0lVweWA3eehpB8dAbAkdDBN4a3ksUJlvxxHkrYZgSnk
YIlxhfvPMlVb+OEk4YjZjjWKmDagYlJ4m4to2lNGmgE2EHpzu1GgDRBPE6YGimfV
3DFP9y3OuBpVXvY2hudlyfcbWbeyFVJyswutYg/gL18DcwL/MKQWEZ3Z90hkgf58
4PweoTBsyyD/08sCMQeuLhwCo1d9OYRWlYEaCuM+EGHupKdLkJSvy1fTyMUmdQsD
tX4H1FrivxTzT+YlNW8IcyfjnBoYnJ0BckdZMYHj7QOg+XMTJsMgOxYT8GB4hhhI
v/4V3JIBXwDgVCbobjAvGCsNL2FUYi4FOK6+N+miZhzmXCwPF8q/c18VArGuIDuq
OVWYRp5ZNSgcgBhsSjAT5U/1kTxTk0F+5NsN65z5t55pdVitYOrSzPhmH815wOp+
KaFtAY+iCKQMehhASG7vaBlePiDr3tXQ9nRar2IUZ1v4roW7J/8RDm+C3yszP6I2
BoKjt+tsPJJFK4TsXKoxeAJmmvgNU8AXHuJj/MbF1ZutwXrPO4d5s4X3gecaDjeV
TQJmq9cTpjVdVEPQdStcbO+fLsPPa5V9/oxajfEf9OVmteP+/2tHAz/J/iiHHs82
H1zZfvBJmo77axOEGyVDy+Mh5skYM5/RxaWRMUN8jKA+yw0FJth0sB8XJQIi2Y4q
MzU+iOn9Yd6JOlyJoSFH2wkm2fv3DIlNLpxrVTmFYx8+GB0WsskU1kA83HXjpl5f
ARDretQZtD+n3ILfcP5SPxhJmb5DiEWLrY2VMlXcbhdCiYFT0hKTSiUx0jXooUWM
/SPet/wmOk4K2qqTsHTNVjS8O2hsEGwRESd+ehPuWTwa3lx7v7fkYUmgBAPdJENQ
e2neeGAhQQnkp07nM4vYpc2YFIERhxY1Sedu1A9Rtw373MtoXX5oRDyGPYB/lFbZ
ZGl4G3NDFKenXrU7yF+WCmZS0dGmyUC08p+PpkP23U50C0HeexGPN1SRuLXjOfW3
5zAqqjfUdmKyhdh8SumKcgFOqonTQzLxJWIkzIN56P4NGYNDojTqFhlT7tpVuPwE
2dpmOGekREwsJz4wp9kt/vh46ps4YQN/dVgKjOAPoDG+mJe3r55m2ID85WwEyjET
FxVE2ZLg9OzShwO9J1BzqyXBSzOj5UbOkjym4eRnMzRkdnKWYofTsq26TKVnLOTg
e4CIvNwn8jq1/KB0Rc2aewzKl0oFe4uFT7OAAvxCd/OgWft2sRjmJ/4G8GSaCpkc
ILzPyAtxcPyULd2DRrc3SChQ/UPA4bKwvOu/oUM4V4rAZyWUHQmhnGzLdCwf7TLp
6a4hICXaSqX/c2WKjmcbKjOiZHreIMoPIxy/zTFXbZ9TMHpKra0M6BVxsK+L96Fy
qo4Am7JuPyxRmbY852OVgRcXOOEdH6Dr5FvhnP6YsT6mwq41XV9OacZXli/Zqrnu
mtIdQ8Ft/n6OEU+T4a92R6pNZI4h1UHEF8pB78NfQtIRILdexuiemBV/KdCFJ9cP
ifWBxOWwuIDs81ZIR4D3I6B0IKD/ab7Prymu0I0VpgOAZPGez/r2+OO4rfew2HDh
vzYnjsm0SjIk+NGKehlSJWffn4TR2UhADM+vP9jX/GDYSOHcgt1OmZjasNmgdMIB
j48WSlFYDMihwl+IMi0w+yfMP+iGQPZshN3I5Af0ztfxewJRTWrbwthrm0gN7G/3
ucIqeHMFt/NMHn7Iv/d/L/RZTxPgPcwwaeSKo1v6uJeL1ewM3suJ3TrMgD6M0Cop
IbhUYQtFUf8bRjnHpbciVHYjXmcfO9DWKAibwi/mavig1q9ScLbtINh6Y3XpAWWV
SCuEtH+adURB6V0/GrTRGw8JvcdbN3CQSGBUzj6waG1Ru0QppLjWq08p+XZBcKf1
VHlJBsWRF2y7Zy/tDulZmR4BVggG7q/0j6GKgrz/OUezTWRLlIT9cwEr4RKjKYSg
3+Fw5ythkXTEqDm+tsPmTZ47BxpPWw9Cqx4YznFdKH8LXAGn90C9aN0wgvpR4VT5
knqNrsDsk2+dA1gMWcz4zmD25vuEfsnAH2TyZlmJ1MpLvNRTAnZl2HSADfK/tZ3E
X20Fcs02oqZCkE/AmVU0qZ2R1zbWT5KaL7p+d+xNvRioIy/h9DqrfVcWHF0gMUSW
cwCUTVjQxHnrKqI9q9X5UJrihyXxWTTeHjM29l3lVEp4z9l3x11DVhOf18mwlCOd
sU+9lyicWbPuK083wpejnkvKn0YLUmbj49dmYdc+9YowK4zSiWefnh1pjzCPBBFz
0fJLWJSSi/WIuQtjNe4+EU6PDNUKXKCzGmLBuVL1loLq5iYJLgOGQfWZAQKSbuP0
np5e/+R6KvPmnW+OE0iPvPMGuKfVAbgkIykBV/XHFaIkSyHd0RLrlT747RnaxZX6
BvaKzc6pKEhPEnco32l0EdlZvUSsmKZuPCf55MjoH7hZIdG7jbPtuGk9WpbObES0
gZZrtpiP+UYaht3iPMxmWnhOVzDGRN829+oqLtVYvVC9FQTer3kwDmMyEOhMXKbm
Q3zxF7GOlac6SV0Xz8amvigI2kPqxrcRccys3wM2BFSI9zwFiheIRFEcEG/Yl020
kkYAk8AYOTGipa2zZDzI3n1pawkXiulr+vPW3Oy3Y0kkYXzZQSKUFCWWqayHtNbx
PNhtTU8XqPZw4Hf6fKOMBN03fcCi9yOrYd0AMKk3PQQDSGz1xZLIOMWwYQGWlLEn
FyXl9KqSn0xyW1qlexYFrhec/OGqg2u+O7vKnzK53+wAHZNdCJsz6JRuyEQbIM+7
/m3HeiAg5nia9ynSndS8QvM/DCJpuc1bisCwankt7sCMf1PEm1zOb/pWE5VkG/xU
nIQWvGTn/WdvZ6ihsufiiQGMq1DQ4C91z08iNCuozQjDWSpYUGzKBjHLvSXOvXvy
NpSvYPbsSBzqpvyPZw691XZI53UTaaHJvvwbLDSlHMGCJdMphspOG+r1aRMsBwDc
DjfAeraI5XEdzGsgtq0hrQNVvRQvOqFkbgFo6ZAsnKdHtmFJmTSCPjf/h1sBltxa
c6Izmx84BaircqXRm1aDqvMC41kAKDSLWILFn+TsJxMLNJFiga8OxLMpCSVlSpF+
lNURZPDCSCZ1TXstBx/O1J7qnn0MZCBQemci40AN5RijDbYrw0pcqPbGz3x6U7QE
PuBLJzhVENxG9AefpqTC8ejUNa5tI5IGqC0l1yHE6TRm7nAhE/7HsjbAjXfqS+Ja
wEvWsRYFsvRGwLC/Ilte7388VQlP7j47g+ep+2hGqsJj49hi5oV1fJnAF1+NjTzf
TEu4fLcTcpEmxibW0ZyV67UNHQoIs8rBIh6RSVjvWQNu/ekpZgtMRfLq8wIGWShI
OR3CiptOHfHDvat4Cuzl7KVdv5eRXgO+xThUZuUfd4E8NY+cHdSX2upJi0G5J2++
Isk/ZmmnXkvjLGfJ1H6bqQOywEmcRWdlyKeh/St65FxbniIxLa1t4T9F65xNXCi1
dLF2fpPcMY9fOybnCgm2FVGJ4Z/35ioiWYsBFPxHoJPSFJo/kUJECiCrJTKXHtBy
oGvatv0m5WjUhPCjG9q00ODrmtZ4qJIBaDrt1+j9+89/j1NtPME/buDlRJmMZJzr
EqOnkJUp5jpWgMKhnRWJbCez+ou3SdrXAYa0Y/1P4fLut0ej+w4irRV6ErFhP36B
UwQImUC1h+5nEFDpSARY0XfGD2mbOqyG9c19mQkkAF7sWOQfUd33ffl+O74LsAJY
IH08vLxTx/6qmmxaVnsbaN41aZhJCnsL98p2rbqmvJh8HQ9S/QpWDFz9ykaGLSd4
Ch/kehQ2BOVqg0e9q0LMkE+AJoHB4M1tK2ptIyiSVuzue1yGSmofJekdMqP2L/8m
52Al+uiaITDghdLp6I23j6SgwEiroH7FuqK7zun3uIcsSK8TIyV+SvpFQV/+wGB1
nhuvx7bpOMB72wK5nYUDxVTm2vzXj0mottYKsVj/nKIlCiPJnWNcig1DbKDFhn67
3XBnGlo/VnxRf0i20W+anJMS4a5M4Aaq3sSiyRN+XLeCanKQkF3U5+R5S4EsFGrg
D9sM2I0fh+DQZN3U+8wB0KQ9dHr19fWgdIsJXMFF+bA8T/Ks7Dcy/yBEqRjwsk51
+ce0V4OUx4qNfv8EGkfFB2YOIz19hlnTwKX40tc95ZzsoFMvfWKblg0XHH1oqUOK
dPuDfqd/+wftWzBQCtdFA8k++vhVLtYiSxlAtCk3UDgLbu5sV4YAfLcZPiqPdFNh
PzC9WXdRPoMhw0BxdhWPvGDi/+JXW345JfV/EyqEurn1xscfqkeGAvnljDH+9rGL
yy0KUht6nJq+PnqR/B9ExwBCYv8tBooTnE0qXor+V3h3CA89OHzbHniz+Sc5+MkO
RifEv3TVLPTB3w/PnLrInHeQSDeAVgktDWx15WH/FBoNem4lDTV02pA1A9iqIbxX
0EhDi9j026CJD8GXCGccPW+g5FES4dyzGN5pClEt/zjAc/lhQZDidtJGhl2ndf/j
VqBPRgRs7/2BLqcSNLRUMWzWlcxCY4Kz4PNM+lVnqH6p+Eo8OO1Z2C93ohB6rn+h
sme9rkXVAtxrjdbhJxXBSpoMquT8rY5ikAoxWqKuOCWrSVq2m5uAOIbXtQJPOt/p
QDkX9nVCDZdR5Zt5Y790mVzW54uOccuZ2XuLMp5L3dS1QAD7FIdpxSUYsrNmpa3F
jUCgDuND4rdufj6LvcT6PlC+Fn0hktKFhA1U/T2aKaD5HVATSSOPjSUDBj25+AkJ
VVbe8UhSc+U2DYLv5rw6PzvDBDVs0e3Ghbjq4Dm1Nvib/w82lKvAhlN5T6sHS0qS
CsZCW3t5AXp8/w9vfY+jpqCCBvMeOUr93ou2p2bNdVppT2S7B7oi0xKdo6iWPPk+
XL0WWA82iAiqBke0bR270vYCD1sRYrBdxU3CO/BI32irJpTDu8jSXxJ1lmode0G3
kLDdvLItrkabET9mW+JcVufHqf4iRrcE8d5FrwINA23rwrVhwqRAsMCLToXLVHpk
UJhypDC4fBwxnyLxLY4rW3akm8sO/CjlXzT9mQ1y0y0J9ZIiOjoATEQIfwTPneRJ
S/LQJfeh0+IdxhX61GH2gb+f+l9TnQ6osanIHrXe2Zxh7ZGHtJGAMhj/MR0vay3x
0NtSXOfiNpkWxbXV8jyMCY8zODtJXsHEV77yF98r7bdLJlNBOOW8AmhvM82iXMLS
tBJZFp4X3BaoVEarUhaZIPE5Zu7eKFg9DjkoBjVXktHzWBpPfC6OV/buOu7aOHjS
mbpR1CGfUEPgqZW0BskMLvdHMJpSuE7s4hhTV4sRnYWjY9AwsqJaP92QP24gKTFU
uTH+JEsnsZZ9SnA+aJaRx24+9Va1P5wkPPjtdTYtnj0xOYxh6NuclItuKRBZTuPD
cRCM6sB3BBaC3El8bV2yPVZcTYSJg/Pxp4PyHwqLx5gjRytBCnortk1DPfDcgQD7
+10bQyo3HCWsorCMZO6X/sioEDj2jzWMyLhaU5Eff/OWv2UERAhkGlKG2VRdS37S
Z9/b9nLXBkOfN8CermQSjAn6dL8GqXhiYrd8NpAqx1CgrTqSs3w6fmcGkv7wXnto
RSlbDkYX3EaGGhYAbqS//yGFYg+LAXtzxcsrRMuR8DQczh9yQaDYEgaDf8SLbnIy
KgQ6CSbs8CC68j9u32OyC/wv0LMMJPq+K8QJbf0wYul3IQQ81rbxDO223mZgF+W2
RVd5Rf1JMy+CRGN7l6F1Kl2PBKK3zp9oyYM2CJ8+53x1vO9JSHRyGQew3wTyibR9
l1lKLMnIqcan6zzYBHs8b1hWwTvnTgE+Cr3fvGNBQq5mqxRoXxR3qVEMpceO5ryl
BmgEtJXKgd1ekDgQIYuDoGA3sXsv/fS9DY7ctiR9Lz4IA1LBINOeySsYwHMIJbGn
G3KrqvLUD++MiPujegEZ3VvIwU63Fzw/WTRioTuTlheVQh10Z3TGWGYc0GxiU4Mw
xKErL49lbv3OG7g/ZPy/inoGuhiosZqDsjHdE9mQ3zmhulzXtiYO9uNZs+lQxztk
DF7gtOUQj9Q4BBM5FLZEAN8J4b6P3PXblmuuRnHjksjC2ERjGb10tmMeTKQyChJx
w+GBecZtvLvTh1Jm5CVXXLebCExWU7vs5jBvD52jBC6A2R6pbjFAGAoL0VMPd+vZ
/bRK62nyMIAjYaT1kZ7/m/y5ZDMY/U1MIcNRVt12a56Vb1ji04Oh3lGZM890yXed
t1RrWQftYTKGQGfY4ACFXvFTZLJ8KD3a6gg6mPIEZoSQ2CVWuSNqD+LERygeVleZ
kGruw6VFSkdU6tB6jk8xIfW+XOL9oCXE320v6dJeBnnYZicJO3UgPaRnVpw+Cg1p
F8R2hOjH2Lm/cVXPDALv94HYHJznXzj9wOBw3jrGHHYLDBF5zBhlsN3iaC+BEsnO
9Vpt/qtvQeTphoW4WLZ6zpAyOeHN1hHlDALs7htO0rD2H3KE8Uin764BR/TuxcyE
710QHHwGJ6C5UCk81lvF1BuPWXmZCG8zV8wjv3IdK01fdcg97cwJiPItbEZp4j3C
Wj/6PuxfP9Znt9/P03QdXdqSxI2fdbXtOkkZhrpQ45FZMdShAppwFApWFJ4sWKfq
ygQR+ck4aVngxJOUO8ksfAefEqMPqXnlk+PErzUov7j/IaoFqWHFOMcl1GIdskEd
dTpPLkoB1g49HF09FJ0kOCcs7V24joN0wf10GtAIucj0btDgac2kWUG63PATnOz3
/9L9RB7l9vQNxU6XF3nzDFwMrfN8f2VFjUYrIcL6RbvYOrV8ibAA2SQ/HTbilfMO
NMOQzySC0q6f/AoLQHboWCKnGypq2ivDE0qe5RKXc1BYmpHflgnsvkDtdVsdU6VE
qeu5mmN9gkS1VeqO1MYlfOwiBk10VO/WAIsDhH61RIYCCyW4ulmmcPyS/1y4GQVy
Odkc5qrZyr/FjpTfY5KXVTnFpR2VV64+0D5uUmokgh6hXvneuiCPLm7hlsfhHGT4
wY7VDL4vH4bBClZuZNYf9aO6VKBVEFTfb14SRfWESpXbVNgdce4ezFLoH7NukpN0
186OgkDFRDXuoOTHjELaF7fJCEmiisYn/NxFOo2/JJckJ3oeF5xWepfLgZ04cXpi
2azpGLB26X2K7GsPU4Y4Xm8JktTYjrsvHXdkft9XCS2aLCqKwWyZjfKaa5kAAENd
pcjJfBDbWiwzK/bOHlMBYNQCdJ9D8FPERhf6rBI+uhy2/2KpZwUdLSO6V8rMJwlL
U6v0RiIoyEmRJ5eeIL5IXp25iSGs3w2/kIGarctWcApW176ihOasA54S8BppH5J+
2121rZx85Grzv0bR8P8w7sl5hE8H+/lGdPVOhCBL96A/Sg2dHv8P6WxoIJau+lkE
ji71+nqLwfVPzXR01O3U/lXWAKcf3I7EXj3el+fnkrzudusbFuk1fGYSEByRb5k3
p1itQ/CV8g45uhe1A/4jru5DSvem08qpZBXFg302ZvkJ+dGe2cy/P7YbZitJ9kYF
fwNeSUzdIvbDVHHr5sIiXozUTPGfMGQ2TOSUR13Rl7erR8txhItuYgY/kmTM2K2P
T5M9zUhdqP7oHvT1zS6mbtSLVzmu0szMkxSYS8tM0JgskWV56qHjHQqkmTUmlTtP
9jXL90EuzCEGIBdUokHFlJujjwSflU3ze8nrVEvaWi5TIs9hMxt6zmXStfb19JnV
WfuBwIXESiYDsweMaAnWPBXSWhBrQGrnUlR7a6PDXcWHNENKGxTLV8V4lg4oWw+1
9xoNoUCE42KVap0znCmwofNcfeiDuE05MkE6Mk1QmVZgk0h7x8LWx7AbLezg3Tb7
u20uTr57A6CqkvBu3rf9ATTIefpzPTHfkbbJNfi0s4rUFtjyalH4wNsdw5c3kuui
7yAY9GXoo0KvgoE3BCZFe4jn7qolTpPsyqGu84yQS8m8lMqmY//9/n9qzt8N2Smd
1oarzXxE0YHc1HXY72wvEe/1rFjhqrn9dBiZSJCedN8bTra1Tplq7UEpt9CzK3GQ
zxlNyR4JSYhT5igBvKVXwAZu+rfv0ejkJzoJxrO9VxQI2G2f8rFdl8+JjMQ5EEIG
m4DzLCA8FAfI1pzCotUhK6m1nyhhAhXTVaf4swwIpuXYA8LOKSTw+Y8FtrVmSBPU
0dOhLNzDdUdOM7MmQzypOXL5IoCuQkArlVerrTk1bgcfoLMnHElxVMH+jpUiRH6s
VFrDoLncmXLJzi4NqWcRjpZig+AE5CaKKIUAGf9cAXI2rJc24NSTWhxhod4xrJL0
sV43A7US7Kl3HSqz5AItAVn7UqzSy0ymh/eaHol/6CDQKoT7/eN28PpQiJdg3iL8
tNwUOabv+LXm4J1EVDpRKNSzMoGeVZ1Hx9PrXXYEtSY578EDlJiG+5z1RGTeST80
ecn7qEBvnf14FmKwP7GEQAThXTAlh9qWFqt9eUd1eFSgCIpJl4cfoMp2dMjixuRm
c0do65UyqN8nJI7QESjVWdapns/UO1BmgLYsCaD6QGG3kgfcmutJtTme8HMWix0o
BIl+PXt0fV7JAOiTBUlY/6Ki9KaGsNHIPDagZJ9fy+laIrGSJyHAOCLbguAUAmJ4
uAsHjB8eaX6qEXQr+zMzSWlgb1WayH0rE2wLAwNbU9jrtzsWJlP4mqV7WlhaufoS
hn/ZDZ0ghnx4PeuBblsRpR3bvgLCeu85YULxlaCx5m6dpN0jhCuWDs9sSIXwC6Fw
aXyo0LMItEoD+zf7cP15xqvMDfNkx92+x5Z2XSXCLvzBk7thqLNBEiG20yJOzfzY
tS8ZibwU5Qt4x2KBReqe7ZYWUlCV/OcJ781VmIm6/QDrpLGsLhObAn6NZjck1TZE
qUSjftaYLh4Fz3PdO/5bmtHOsiWQLcdd23TfyRjwCd8eTeLUR+f5hmTihl4mfC7l
WmBt2okIO/33kcYas1rPEGmwAK0vyU1qsfbQj+2h0DaKLc8kULk+jZiCA3+i9jDs
vjEZagRsVLaUw/16Tcp3mSAc3qwl3SmuEmtiMCgHpxjtfu0xw6LzqXbdiZd5ErWG
egH7CgP+qx+HIkdd9mpdXzJwWwnaGwj7F3Qah2/KFTiWH5xmXU9NthZuo0LnqUZ+
UJJ2EgiknsrGL4wQ/M+K54dHITkmXVBJzVnHYrcauXNLlD8x3AfIWf14v4gYAI7h
/56z43HnzSHJN1mLtxdvNr9YzpMW8MIeCRzl0w5WxieFmTelptcUghwUup7deqUf
ZtWFJbk2YCemjqBujJ/lDTv07310inHwTaGA9eLifN5zmaUGWb++yNWakhlTeb/R
24LFaDPEatyn6GOROgQ7NG6cjqbGEPAtE/fVwRIKaTiAFLbnfYAhTHM51AZa2ASA
+JfP+yeT/x11MniEpCB0oz/l3uiYKMJhchgD8Cl3L2U0dawKqUouMQBRxVACy43C
8ZBYqcpveYWv4fBtqcyq/+timIYYRSJWR6gIY8kAajJ/G8VdBN+OHaEov4VvmizV
QT1l5+PsDhST+dvNU0HNCRkRiJpcxJpGdgUJLFNQ8t8mmOJG/L9UqlCwOtgplIxG
bFGI53T53RotNdp4x8VVYKnTaAw7NIGfm3lC1hioZkZ3bIb0c/zCpj6f7UzZx7V/
QbhQpBdBFd5KFvqcRB4p+xOlhavxo9QWXKgCpJCFmBBEZaY9xPDCzTxMoXCZ3Xc+
IyiKmux6yWkYYGuT4TbvrGCyrE1oQczubnvxUx7nqHe5wgIaERX9fJIP8ihkF4CC
EFLIO1yX94zFpbxePEII0lHatjw0eqUMhvCg2E8Y5iHhlSxjWCkQd8FGJGXEjxYJ
3oBh9yQofgbRS9ps7ymJ0zHs2D/MGS3JbZs7/1RPK+KNGE/0b/1ZCUjXu+QvfBoA
AUZia0d55zkFpQUMCXQCAYG79BPAwE8m4Ay245Pdsjp+Ri3E6LOA9Jo6gXY7luLI
5/fYp9IXRIEcB5qINoMX7uwigQJb+o9Js+ZjHRx34brwfXRFLM7uN+XNevA7gfP9
fiuo1fmOVoU31s0vw5/boUhx/XtQM69BTGjeHxNEQ79Rx2qKb68CyzC0VpYG17Uq
9DTHwmfZ+OLPW3BepKTIjs0ubv69XE1jjVXRkiZUzhWcj0c5VrKD9aeTmw572Geb
2N4eK7eqIXbsvgY/GiOX1ikHKBfODniG0JqTY3AfM8AU4Np6/K4oBfIGl2G/x1ki
/B0gi0ZNdsj/67lejbwCW+PTjtXlY3+7YaAP1mAygdVQ/W2riQEGWLb9EjPFu5yZ
MHcHw5w8nD+uzBC9jIF+uOGY6zEPDIda4dvUNEm4ChyQvv9/q/TiJWEqtCs7xpf9
Wm2wX7ZDNg+x5n7MsivPvzN9KikIdXjCpx65vF6/Qk81mPo0EM0jSslPe3c62lRp
lMpp0xItlSiMuK8Bzd+cBrh3sKr1pXbRwTaoDiA9iRDyWEP1GjNkZZhbp04f8Hxr
Bnn7MAUZRnpP4OIfP+RLJZZi0juDuzbUdXYNGzA/yPCJU4f8RaMWajb0r83HaJyY
3zbARP7pN54lTFzMf3Zwhlc5KepMugI9NC+G57adNugkEtauUNWvAxxq8Ivu/vTc
Hrr6nugNY+OYuo6jKwZZHWaUZwnRk7RPTweZXY5ORDQ=
`pragma protect end_protected
