`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
IThk5GeuYD9ROL84KxS84j1YO2q/cQkHwGqw9DnB7fvrStKcpYhLKo1hnDzBjCOl
crPLXhqXNbax2AiuOHNumsV3Q2JyLa1axL5BL5EHVx70JTBuyYbpKkiOT0wfn1ac
FD0Q+UXQsuRoolo3Z/eb5YTyGejbleRJG3pqZwd/hV0=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 22256), data_block
tzaIr/9uvaslJQHwWj/FJCnimXZ6GBIPLqbxyca86eAK6YRRmYJA1NE/Yo/XUiEo
7MjEtihxbn/LQg4bnjbNdpr5RjmrLBlMe4oW6/aGoGAQCwmg1gRsIiMC3AEGwXOU
KEKx4Z+9q5k/wGOXqwJ4hnudw9q7VUbnEueT0kRRgbaPCBRMvbvSErFLx+HYNnjr
AQ2iNNEJbBbCeOJlZwvgkrF7DEdSxWQ+erdPmQcnAKj3yxzQyc203pW+H0MRcAH1
DWy8axOb2LnB2XKTK9OeQJXPZy8YIMVSEOTfkhXDKr+1GU+dwnxv7WFY6TsvzHWx
qOFbtFgV94kUTfU7Xp04lhFQgJF4zDgQbegv4mDkw4E4hqnQBlJwMFCgmzACtDcU
Q6y0nFtYyHwulhawdAD0At4pJvbXN5cZ+pOacddgSnZtRYIxkrwVxm5kzv1Tg5tv
2x9U1v619CJ+t4N1KZLOKZBrKxMkDT2ALvX2hHT1X7A8pffaYp1eXKlQZCyrairN
SR57LmTzULtO3sEqfamkmUNiqB/qb3qGc3vnvYkMISl9BJIPw5imQNtoU66DfMpG
Rdp0xK7TP1AooAdpv16h2hyUY90krODIX1s/p235MfUdzfzlar2j9ssuswp0IqGI
jRxOtCteNnOVoLYJE7ZFwpfEJyF20Xn3l04pxhJB6iQHtr0rBhk9CvJW1rX0gXCj
QBkVXcIv/U6I9kvXHPaBquMM6D0MjX1YkbaBsUfY+VlrU/zf+LnQkdjdvERfhHRh
9m62Y+5U1z7wNfOhyzyPy/Xnd+5m7oBUMnU9zhmJgb8S1+GieofXas7V/15zDK5A
Bk1g2xg7GBYnXRPNhI+qMjZTOE0vfzfoTcf8B9ILInzPCMrsHW0cezpKBGCBIZ30
mOsbqb7bkrOj7hN1Ck5tdy8c1mANQ2uASO8NLUP2dvaJZrMU3PyjHScaK8D2VwtF
aUYLDoLdGtuSC62xG3aEY5fvuFyOFODuq9pq+CPuw1yyLQrMFV279am2pRzeLvzh
qEuhNINvR5ufaZQBKUAuVWBCYJL9e589NuFBsFVRG6i/+KpL9RXxesJ7Uq8kbcjU
XnvX+TpSj022wM0tSlaNXXjRFh21EgLzZqCvb2xFosxW5UrZ9FPhWtRa8sxv5M73
TqK6jscCJgr95FXfhSBByt1SVyEg/u704q5+dGkQwmi0Ga+Sdc/yAVk7wb/HGbjm
JABqDxGX3zO+fwKqBThJM2fpKZQdQsQaWhdrKEPIc/wN18DouxMBIpgqPr0FUdsV
7i6ickV1axnzxLerQNwV5YpTye1N0u2McR3qOZLcG7aLArYOXtQ2xfLGr/ovBZeW
7E3e/RaA8vVV/GplSaoq5BlRF7c1K3MZkMNSCSIGAJ7TvJgiyAXravizX0UNsLRi
g9P/m2Grq00DWtT324Y4UCYeOaMJGTyS347s0IV0mnZyLWNAFqcUDXFQxMbAiVbF
nlfWT4+iphCdXAMAtPuFUtHmRaZ3/BE7X7EDV2kiEpnMr4sS+UcyA3etSoIPG0DC
Ytqhrm/cARJ00rD/+MAZF50zTnAkr4/Nt8bu0GFlKb+gs+oTn1xRtuFIQSZYahwZ
SUi5fcqP4ZVZXvk3HP8vx8oAuM3lgqfXLMphA8np32FiV9REP308SwxfRdjDSj3x
ksL65U/PdWeHLHkJk2mF1VLZEXzHrHRspO/skx+LBevLBl5J7w5Rhf0QMPO9gU+x
dNDYOJMkZuroJv65JK4Lh7mVdawWJ4kwM1Id2Lqe5rf/j8xu7D8GMQscRz3OmR+Q
KYIP6mbzdTVkTlYNvJqM5g7gCP2Xf4zswJdm4iPtHFTnaI3apJ9Mz/j8z2uurxoA
5E1J4fW7K0YO54seLVLcIcFZKSdLcTqKCkOdv5hW+Rag3eTNVXMDnCZBXizhPngg
LlLuuBogsxMxfOMbnpJpVYpFUCHNKNUvKO+unqoU4coAk8TRERFjuiVb6IixJuRB
0oKfhB0GyoDbZPSEjvqOgzAfTMqsWbfiv/neMld5DImV7tSlZnSnlim33bVXHz1J
ehVtmcnt6CjzRgQ/Ppo4T6ihiXPlUCU08ItR+B/h3rsoqf1u6uUVznFdOVH05Yd+
2MYEq/cCcFY4OFOeKBoUEoAznulBxBuhKOLrt6+SCOKd/ZKjfaMpxs/2kYlV5Iyn
RTXUzt3tFFxC1UEzQz+mhPQlislqhMr6HMW6Oj73tBJqa2qgr39jKwqQUSWgzpcl
+/7ZetB/PEllxL2Azk8AeejOWFI+wWX2UAJD1HCFqaCqEbpD/r8/0Y/BRbMKJkxo
G8/vnLpaxP//+s9+Z6KkSYdQvUD6YjSuU32Elr9TjQS9m7kKqMYWB4xSvXMrv3xj
cTci/Ho8Gr0AgC1dLawo/Z2kg1roHXl/KzU4iZx65Je2yj/70KBLh+uCdt1Fn5tE
0F3s6hBmKQbbOKlftBTmt3MeWXnssLAYPekaCqAHtDZjOkXu+qpWDCDkEvxlg65e
Ph64gLbGR5CzkbmxPK5U3SkfkqtOgWmP0EtvqJqNdpK0ci5RHOrjsOOwM3Ld3ezl
wD91R4BSgeNwbPmkIyE0Df+E9OdgOTb14QKMxXso415M9Ys68dHdobxQ6yuzpJNO
Ie9eSqeYS4u7N1JuaqEVvxtt3PGSJmqAAZq1DYUuAQu4gP7S5orO5a/PTcyr0byK
MXnx+xd5WEZjmUSe/g0IQqZoPAn6rd00x6TjjYaY6oy6QERxjKuhTqRN969tLIgH
UVXsOarCkRpite9yMF3L5OLtHGDl24Xgvy0nr5GSOfVD7Yix/FGkQI9vv0pEdZb9
Vk9sH84k7v3JF1UJFNCCFHKQD7t2YK3v0FiG61tQB9Ln1GmEqetnkQgob2OAaN4c
nIC+W9PHKXVAl3I14b2yYOM/75Atq4P5I1p55eC41bXtSKkVKOMQOah5hjYvSYlB
geXiIi7aANLTXxZM3N5kUEqmHPbUl+Cvxe15eeTUuNcxHeARWlFkDY/R+bEhXjAo
66bzUus9Rioyi0NzWV+OMZkBAs2US+ExXx9w60QNwDaNWFr12xy+cQ42mFGKk28U
HD/xRDC19MC857dhoOjkDwQVWYBwFzLjRIVG2y5xRxYgjtZ3J4Hdi4jiGA2NI9sz
MdfJnBJQyDJSa/ZYiCy1zVGQKCWdsfxPclIegsAkl5Qpo4kYhpq6+ESXh4J/gJFr
ES2Gm+fYyrpYtygxdf9oyQGiVKEjkzAPNJ4bZcrM/kXNkCpZ2K9rLR0s9M+H5jaA
mO/26I69CG0Mg/WVAHfPrhKGGiJrBnLoCWUIyzyqT1ycVuejmKmnjVia+tMQnkmU
x2AqpkfGloZOfX7uJqJEp/Ryfe/iix5KffSODHNNRSgmBNKsIFxJQ7R875NKaQzG
TmaWA9HZchod0mrwVCPNXBlvQ8jm4LhkPWQB8K3QkgungG8mTs8wSAEPfrAjWl63
pQTybW7jEqyuFwuNjVL5TimwaxowfVQN2didvVhjuw/acWtVfsm4ScVqKlKyVoEj
04jiERJ6sYXPYcxQB6na3VTJmz8KsFNsXv57VU7qVtWhq3veVoAkF8yABboXlsv3
fusARbDPwwbPKGOor0iIVSyDQddGHSeaAlUSVtxW2nqD0F3pzYwZQ2XIVNLLl5PM
pd8sGTUrtOFTcSLfW67yAK2OP4rtN4LuuyIWAKAHKkqpqdXdbrwCzKXerQvsNE/A
takH57XMH7NjkCye0psysb2dDO4h/4DvZgCcN/T98kAttsMaXpEZegenpv5gcGWb
8xY1VJzr1o+mytxwX6mYYLgeCuCor2GijO2TFCHdzC0QirPHdaHKQHKNhF5Naovz
ovr8gKREYmHmbGyyZ0Fqg83ZvkmyecMslYE5jT9frIKraarchX2i6dAB3GpPAFZ0
SVgAhUWXiJ6So6Vhr0saCq2yVM2QWyFqPhBDz6XtVyS6+mQhGY7GdH/lm7zX1DN4
LtGCHC5etHHdVK0GkIbP4S+5dwHrosohsy0DBwLf7Q1wv60n98mw48XOER766+OU
3djKpChuI5TfGV0EAlzpvXVPZkoqSQaR0y10i9NZ0Yoc+2Auali1kXa4edtlgkIA
ZBpZeSzXiMIrhoRqS6lArvJ8Ypg5434nWncDvsMFj5P1ANN22YrHJkW8Aa3eYUg/
CJO/ymzirg+jNnTB0ufM3PY4lwMol8TbNYuqqjN/IQFOM8v22hZsWls3VsiVprm/
UGrtZw2ZFoJWZWanlOGPo9SLEoXNmvo21YsW5syb3Bkt3Ifp8hTmqHdeA5qGbpWn
znAmozQIoGCRgAM2pmSWTuJcO6tqOSLPXFgiP8x6+dwn4otK+8LyzlA/IxVQ4MM/
tnewKJVoh6AUO7NEkLKoDxohv2E6AVwxKtMLaLCCdgfhy/Jbjh+7driYIvBQgJZG
7AVtZTVPbQbW3vYHGpXcBkaxqimaAK+Mau6LwjHv4MvVaRlAai4ER/oIt35cBhVb
sZc1inWcgY6gI8fY3Oesg0SD2LpcxXYH6EVxh/6rIinIKWEHav07dujy3LblCtIf
BJIVTRIFVud0cQm/9yQQA2wmWpUqJvR4hRxBi72594N3BEi1pb4baZ6g5yZGmi+T
VQD+p47loXVyqdLn8eRhglN3AmmP9C22bLLHEJvBY/c5m8F2p5cJw3FmYmkMThiM
sLFtyrsf6CNn2USiXzpq9NEVbfVkWhBdn/E+/Z74kFocu65PfLRZZ5NJk/7fknPP
MhhWPk9X7tamoAEkhJcU1SkpLeP5ZNNirFzgn5Wj1KkD1Lsf8lKEL2/tm7IAWdZt
X6bCZM4YpYhW1DTvdrJQZrMuTRYNGiP57CtegBI95s7twDnuQeAuL2S7/eNBtwqZ
l51JlrmxYK/iJ1XHUHMk6WQ/pDkYi/W3vXnVv8c6GTI5TUA6DQkSvuFCPd5T+3pD
giNlEvDtR430Rjac9Mu2shOKvUjGpFd7EZ5uSIKSt9KJAOpRot82kO8bEt3GEUls
3Kk7INtrcIRjQ0HhNVEkJEe1Y+JI4cSreF8rdVppoCgX5fqYKiE8JdlAmYklC23t
7QO3/Fwngj7bgaRDTWK8j2kUa8NwZDSnbEpuTk9o3oglrNI8OBr2rsA8iBlEOAYi
91dFrUs6toMF3V5xPdqRO5JPVHaWJamWHhDMUA6xQt9iKjeKXsEfOq+va5IdMNIy
fgQj+bVsTmokdiXIpfkB/r36eHKDOOVyWooQo0xrSA7YxFkLREzmMKb9nL6TguxW
Cme60yq7i+rK7pllYUlv8OgejJv5ePJj1BV0wuD32Y3aohWXZu8jA7kfa5i/GPzR
Nyd1ZZnTjazJ33F8iZNnjCL3WRiR3ICxQVKPTggRklLu6vIICpnltNnCFQkrQXo0
wfILSCHYogJ0uETGAiU40oGwi0hPetg60m+Sg0LeK1t2cpZcgL/V/csa9oou+IC1
2jSzdisxQtlEPViVcAzi1RO9xGDPJZ8a30bHZwGrXB2SxEGgitowg70BbHFw3r8N
5de1YX8gJKDKA3gV/TYYQwx6nhJEsF+AFdLD0/XPcboNmDfeiBA39fHkBV+NYscb
AEr2Z+qAuW/0IHIsUwWPQ4df/OKuV1/xik1FVYutF1XcE55k5Zemn3CzpTHtp02h
xdU37IP1jW2uIu9AiQhHij0mx1gMOX3Ra2wYHxP2sp4D4kBEzyIZR6AuqRDZpkxp
R5YD+kPonT1UE+3CElcX11izzi/xKBZK/MlVQwOLmm89rNGnNRMlV4i6q7T5UvF9
2nx0ijAcTeYd1X3krflOFUkiylQQbbKCMOeYgipU9Pw/r6MTtfYLRRIPucKBBSLf
msAWwQDgg9kEpsW+xC77Wpkn8Nu5lRy4qEw+GcAo3CeIQXQniRTNoV/e7eoEyZR5
hUAsCJmmjOsdIqyD817geKcaTjIantNOkCRx/gh+1a22v2M378iVVyj8og4Sf0A0
Yi/4sIquXftyv6phDhDBfEX1FcZ/BXp8Yr2blbK1n1yAqnaZM/zy6eh1me7D8WKQ
2ptZcOAl22VXcE+nI9bzSKK9yoxhhekIW+EwstkJ3zFOuwRF+3d3sCptI4Utvc6K
/6DC+QZAzVTTOnv7EP+pNIqF3y4NQXoL/X6syigfelioCOqidiGZkK0tUK9ejQUs
5XhkZbDlOy9WENzFHQ1URS8IxB1aE8UEUEB28byGyNQ19V2LI5fynKVDOJQb4hCM
YAaLdE2aNcUrPUT4yh4IMeeheWmr24AiIUrvIUZiMTObJysSwSy87Uwri+b+t4l9
2rR+lpk6+9ib63xPNg//MQXzeJ0udTPffNjIRCGfb1OqYANwXFu1+P3kBhemCmj9
g146VINPfrinfIj816I3aJ81PHe6q3ui+ky5kseERosYq6+jck+e/w6u5jQ/L36x
fS85gysnDq6rWkLLbefYR7ujBAzq4eNYBdAYYMmjl9aAshfEMzbBSKG8P4Gs736c
m5EAASHVQ5CvBV3wax1qajSoIVc5mnHxtt+gdrofH1/MMWyxrTPGH78i6x5wc0EI
hz8yKaOf8OTRgFRvuCPI1Vmc01g0IhlxCPtxqDC/lrCKchBdigfjRslgvT51xZk3
TdDBNWkhWYN/2BInZ7Y2y6hgbcghgJpRkyrCFu4dGJZC+112X+Fj3DTs3UC1cHRz
jB/n0VHDE/Cw0yX667HbH8Nw8qEnxPsL+P7lOcO8JBYotxYYsCWs3Cht8YvQRmDJ
2D9Zrva6KamSpwQ7YkzLkPc54x0V9dtWATlTvcLLK2WHABDxTHHOvRQ5wAOhZLLJ
Si0jDCUbpruWgIwBLIEyitVbpRXJ2LwON0ScEKU+qM2Kh+XUyLY2Z4ReE8KUBwyv
P2u1x5y3/YTnRMDoc7ErR0FfZAH+r57a7gWVBoK3nNDUsk5kGZOUT7mwCSAmlcdx
1X/eo/rYws1LplNCiOSWA+kR+lM6BP2hDJNjnbYcz8vPZM1uffYWLQgCW3vpmmJG
madsy9zi31f7CvXaVOgOxRmayTRyJyK1V6+iG42wzKRfNAvdc4/7qJR/GL3w8KkO
OmBW7UCUEV1XbGKmsZjTvpvWojG2y4rBZaly+kO7z1/dfSNFOFfBgAJ6EzTDCwJI
RUFyt5S2OI8zc3jaSEj6nilbJnPHRkhTvkZdrRY/i9zFmaLYwqdUY0MfJjK6UQF+
O6A0OHe5z83zZWqIm9xQAMY1qrxahGiRznuRef3QdXtCuJQO6al8In7i+f8HJtCI
jK8W5Dnh4DjZXgRN6yJLGK6KcSZvpg6yLz2By2094iWeJteupCGauP30JOAyl88q
+RioKwp6zSs1HTeX6xSNCj/WFCm9v2OpYwlLNLWn9e/+8tSXUxalY1Arw5qwgXak
9XcRGN3/6UiRZKNEPR6yv/iU8QtFlMeSutWQ5bxVvjVIOw9w4AF8tBnrvOCwD7u0
nzJOcpAKReNPxQIRkE+qSoBT4NOUD+uvYmB0HubkiHefSQsa3qS3PQDCvCklkhTq
+4H2vbU9mMM6pU7lkIusLg44yPQcjoFUDRGEAJ5HKGdv+05p5jMLTzCAI8sTwI4x
qWuy8dELadDhV+lD4J0NuzT72m5lqYRqGYLA9sWI9Se3ICSKyzA1+FqUiEoWYwh9
ey/4KMnG25EjHpNgOQsKvB+BoyvHbFSxlAXhqtLxK6WPADYOXhVfeglvm7qC5GnY
4f1hdeYz7HkqLM64N9znrph8HKULyO9aidGhy7XkZk9bOaPQ9JlM8FplB7Tlcm/P
Wct9/HwpQn6Yq+oWDwMzhcGI7iJo9+RVmM5WSzeBd9P0+HNT4ZdDALcV3BANgh/w
d4H0jaA6LrZceSBGtFfo33gGMvFA+QjHo9PkQOXOOEmRisRv3O06taPo7+YHObC2
WXxoMpQ78YDSipjZdhSHFLNFHYoXtblNb3R+oS5g0JiaKLV6L8WwGea9bkv3aCgY
iDsjQfQUhLkAKnDw8dJiRijcvxRy7rF82lrmXG7sMjRdkuhSWzhu3ehgCVrGE/aT
8tbxhA8/Oo+2STwY6TGHbOEOtM0who5OknSmBjLEqsPI3+ECg5iSOYAHxHKHDyTI
GyyUe+dwAHU3j+Y98eUMSScPlDvFlFQ1QhjfWlLWiEDWeS2P2/odNjNVwN8U8HcP
pvqyBo56o3XJA7QCWiM0B3rVK5Avt0gk9KnGHzBPpSoFthY4JElIqYBkqbbPrkCM
YwmWpxaHha2weN9O7U2udETcDT+J60CEAYUrI/jLc6cNgl0iSVcqGnHkmG5YKuE7
dmCSKdOy4nIK/WqGCGFBm2kaokFLuZrbDjmpx+glB1dyEeSrrrMeMTKRGbSbiACG
8uOD1c5hdsiFafvCeKD3IjeR08unUwoA/oR6P+oqHhNwzX23ytpNVL9b/mJbxk/k
EY2Hmhxn9EJbBAvlC7kwdLCeHtgwv8MM/WHZc7zTFEMqfjWoawSy6n4UOa5P8SK/
1imCccumUect0I6M1gjyg5/BpVUrAXl8xiTfopk3k/ujAeHAU1BcXGmYDgdFlLpD
tKPrgwZropbapktGLZ1wY2ar9bdy2kr3Oci/sb574uu0riWXtZejf9JV7/qDsrEu
oX5pswVYuQBsfrBuLJNn8wu8/BmKp79fpsOeCmRBP1qfc1A/dmuDVQctWEdIm4yX
/vGo1TSz6/piItvNpiX15vSkstt3TllsawrU7DM8onsJn0FGEZ3TVgTprV4jiwLm
tL5ECGJgeupX/biu8hPTuvy9crqcKGth/nh/oL1ZIx7tV3Ob9+iT+QbEBoArrBTS
TVy5sfS7unof9cdpl839wBSR/pwNAR4PMqlSSE8Dc0Hm2r6xSvsWo10D5EzYzdyE
RLntb9tewi9ZOPwwuX8U0Po53n+Rn16fqIkCID9hnr0Pg+2U7ynUX4eZ5rt4bptA
oPgQvA5j10Qu5/pZ+hIqImn6pIRL8kKq87l4MKs5mws2oBfAxc0/3HQ9ccbD6RLS
i4K3UCyIvtNbZUiaNndxDiBED8F4KMQfte/A/ybZIFEPgOGEi6l0/NHFC/UAAWBP
9LD3uXhIEgW3i9oFTx3G+IcZAzWehcDFDy+M5901ur2Klb+UKPi27AIXPE/XYWaH
48LFJfuWgSnzezR5SzWOT+BcH+ggmL2XSBaACOiDIIB3eWKn5+CJ8HyWsq6ju5tU
pJmb0VzH401XXp8GzpqjYjNWuDL1mZF3mjbP2PqOqMV5Tny4FExjY4+Oxmg+a/gY
eQyKiBQ6L5nAzMHGxDqwAoiEAs8rsuaPVO3N2GxsekEhAqDgGyKE6llcVMQe+oqQ
lfx58fa8XLdDsVeuy8JIv8OdzzY5qhCuEhJ+rlxT733hgg2eskN6sRg9Vhbt/TXg
WCBWsVHGFX+dzoNlLsp3ImqKqcLOcR3SCZlIrCD2t27geh9ckzpRCpuU6Sid2Csh
awNpldXtueLS9jihhF1YFMPqbZBsY2RcWMXd2XeSsGsUnoHJkv/+d3L7DkpqB8KT
xkgdQXnImvZVIsZKPfKwpiBMnDqgQErO8IZAWwIsisM4VWGkRddZvxb/xd5bhoA3
2pFS36H0B3sIzqcWuqSsRIcvzFD9XHJA4/Svu9Lf72JBQKeioy1V1GDeDK1rh4Co
zuBxLn98zDVXmkZwSzWG41l7pgd//aKcXxROC+97UEbPX66oaMB0p/BTMGeWUR9u
zdTMXfNk9Hz4d8AiE7D1bWnbGGaOWNPolwAV28Y174L8zbfza6BisdJsLYBojyje
2FbxPDHF9Xc8Uvw7Z28kiu8PZtE5NsQp/9Duw/s7OB8zyTMfRp7MVp3zoLMlEUEf
jR2dYQv75PH01g2KFjw5K1JsjFcbvzMvNSP/zrhmiYtlPzYH4KSUehoI2JHvN6sM
/bXp2AdAyA06FRZmCh0T8hBMxw5hRmDA2i2cXe7cTZFvLWDSys/yZ4qayrlLcJsk
UFSbvI0iUxt07HIp9Vc9hWM7fvAhfogwYh14A5a7xlKdr55zruDNKZeGZJlo3X8Q
h5JGHCLpHpyLf3aVIcAQqYF8XmOM73gFHs8P+q1n34TUFllNgOiBgjEwFPACB9OI
xCV9xh0CeLolM5l3/uUmV5fjN1FrGLd0YaZHkLENCpQ0fawuUaFYP1eAKD0xCsRn
YqgSLSQ/CoSVZAZ2s4LwdVB1ivTQMVvWeTC3LH4GlGRWyO13Ps7okr/V2tNmbzTn
Lyx56smI+w2l9OkhD07nC5ajRpddByr57z6PlptAD9PgpuVYzo5EV/3yqgaJWW19
xiOyOR6JMrz64Wt9JjtUs6lLj434uLIiNQoenesWHPyNCz2D0JMYu+M4sWT8aMSP
SnFIWukc0QPNu8pxZdB1DjirTS3gaFaHsAgVaglFVJ54Zplv9mYwjMPA4LITmbQZ
BxZ84tfUuoUxTtvaL2fw8nFDp0AyXddqYzjkR7LfMBGgdMTmKIllniEIJwm3wM1/
XrW5iyJoetPlhptJp5Z1LppDnd+UznbzeF//6lqIbs99oB5jREGsoxynR4reKGVn
x8sHgG8V2I4EDaKn2U0t14wwNN4KaTzgyruEcueIaBNPwszvmI8SCBTD0NdiZL7M
3JY3WwuqnRl7ADaoFA9iBXLVa8y5Xf0fo1cOQZ56cC1VPs+b6Lj+3acLv7JuI3Z/
NssT8z6fox1kalAeMS1Z48OzFICxr6CB7bN7i9VH1qAxhvCT5GGGODKaDMke00f6
ew96RCJhLOaDEytgkIHQfFZNEXNSogb1IzkolQDaivUOiYMed3Up21/lhfPQdy+P
UN304ZU6lMx75Plxp57atPxuHzeF52Xc/WQzDFBKh+qkAuRuvbmELZ7TOBUtGnIV
dQXpBikla8LQoxYd6LwFIghSy/aidW5byBxdL5YaCe7tpe87N7oKL5/4YgHICF0p
NAwJerUN7+GxEFu43+R2moGyz7+fZ0kfA3FpkM7Ius538t5kteRO1pCtBWrzTeLt
JSxLw/V12jtIuXINbK4w6nJmxNj6gMOqmaOwVvAYoy/Sx0rfJxioWFQU6nh0Iivi
P0ces5hAJspDxwRyj/kwDS7L5H6i8POXgndczj0aIsPiO4vlljC9hGeIAqkBZK4M
YGhXbgNBPeDXDF72C3GgTQd7ESQQC2U+QTogtNAnwZFtp9MYCsX0tl0klVd0aDCq
8MNOAHX01FBse5o5Vc6fXd36DCJrG9Y+rDIdhOemmcPb0X+D8TpEVUrg+YJDE3Wi
dre4UQXU3q9JGgQ8TUDCh0i10SbNylWwtjwi4LD9KWXkve6sLftHZ6N3kOrT3EWB
s/Cp/MvdLr4UJMH8H1MMjklgUutttEW3St2OMi+LScd2LOz2aW+ufsHiu5zj1kc/
KgJfeNIL10gXgt0Kf7IO+wUaNH/9LRK5II0OZ1236NyAmRPLXZscHElpKG7lCAm0
OtlAxIjIPxI838qzB6iU7Fdijba433Cp6qo74irYuUsf/srhZdV2P16gcTsnMof5
jCWE0zgjccU9lu14ka7W9u/iYYZ3FDxnxPmQA8WP7Bnjl7ZwLd2UvvYjmsF+Fs4E
ayUgU6Ic3pszKq6KPyRMpqlzwGb+CI87CAalWpAnYyfr8IR7lD2XNh0SjwgAtO96
VNtmkR2rTQw1aF3oVpEzDTiHrhFGAB1WbZqRnBC+d0/r8K5sMuhPL0RI5/5R45l6
rOKisXSsi1TSWw5UQOtaspFIH7HKnX5gIEl8pT+kR7eh8d6eM7BvUZnirKDLddtN
dWSAC9gxBaFFf0wKx3bbKbPctM3Cx3Hra8mBIS8XetOR1O8dg6zFLQelOpF4E5E4
Bv5d5yvrfLKJhs5xXS5lUi5pTGDVv/4eWL9Y/xVSrTwfUxebNB2PT+CsaTE920vG
vD3O3xG68mRyUborYjCiPmTVfWqt0EsLuJ/tgwgBd5QxrMFQhfrIzF2yhLVboYjA
UraCsrMIMkSOcMx2RRL1C8Wivb3qnVCPeyNc/nkX/X0dKc0nhhTVD1rYNNihwwDr
45aM7gAoREHGKk6hgsFDG6yLTbSgh1jA72yfG64oJJtxsjCAJ8iyaTYa0h6kOo0G
999QUQIHzkRtGNe+3wSIfwPvJWMLIAtHvi0IA7zDTOGma89LuhWQH3iGZrL5oRgP
oMdr/j8g6x22n0QNFlzaLgGWGYVbWvyqQeP/bys3aY1DrCa8UJku4b9+7w0s4VXq
eFMSRNMfmqKpnTIRGYa2xzdyzSJEKX3RBkXdXe0rFQWTdhrn5p05vrMYBB+OLN3I
WUCGkiisnuHqRgu+2mqN5v3iOWjXjUQbA04T4OHld2l9+2+lja5wGlrsIX61O5Gi
3+Fpqs1Kf2RpFrxkERGrg5p7mPBMtgdPaAJEyxNCGpi4j+qLRH7UMjNzhyrdCf4s
9btxegS7QUhe0h6mKqT0i2yBnOe4kpos5KTH1deKhnRYy/8BbL00VjybhD7NuSOy
LpXG8vjDpLpZdS7/HAFdiDHjhu9/wIkofihPFbJ9fcntzQTqcKmlB73tNrxvVaxC
CKqU34hEmzvgyK4iH96dm5YbuWNodjhSlrT/KDnAy+1fnA4Bd3KuRc2z3Xy0IcbE
fsSuDzVGZ9HLPysTyinoKCHIlU1fPJkDXyfx+noeDbE1bSqoaylfDbAzwEAvfSE8
v34x57EA3dZTBdowPXkzYTPDPhR4DwlurysDSZF5O59vMrxUmhrICsIzY6oR1zYd
dfE+oDQVEysnOuV384heMIC38z+RgnZxBmRRetexJNrpdPNgE0qzjEPn1XxtJ/KD
74fTGBdlwkVuAwlsBK91ACnn2XgQCCTD4eznwN/FVtXSI+rJ4rWOHQLk851L4+e8
xeQ2Ozj3rzOuBxvQjrjE+sDCLqWXV5SzAXkrmUkt8qrcpuuFQ9R+vxF3UT/ffhBk
sss1MjL9Tw6arxU2OLT1GFqIYdfWy0C6/CjaHMrPpm/GRR5TqR+xasg5TMNL0Ic2
bC4RXyU/m+6Iy1v+wwkMp/yVlIE2YB+6sUjOoIlIGakl+pTBHYPvdoCns8L5J51Z
PAne7M4HYhmXbuSVveprRlALwEU4pGtdVCQXJw8WgdY5Tc5lTnV7BY9RLR80l3uJ
l0lhQCR2Bp+bdddvNtpGJq/JTvo6TJcdOP7JRqOa/CbHAf8hcncIaTnRhlanjZZe
nt172IgS4TTqD3oOqQHWk6PdyfqeioYaNrzEc87H9oEZlT8/XG9TTOYPB7XUGZ0j
QUSmQvmgbXtfB8qPWMvoFoYB03ksXMPM7u+aqOc06K4X8/m1pC8CiUIptBlk7Cd6
YO7Uj02LS1q638aVKOtaJ00Ig49kYq+J+rhvzL/LIvmigSmYW89HxA3cziSAXTNz
FrIQdbots7yL8Flwpx569je69+eBfPCKGOMsgHiIIVTRs4uqSCkGhyPewr/RJ+CY
BtV/fXYboIC0qsLI2K2025WnvDb7/Avy13Lep+6/kybo/rMvn137dfxq5zN+OLUw
0+4hvJGHmXA16/4B0mbsSLoEjNk06lJl1gCnZfXCKjMjZiVaY4wmUPG7BZ0UYI0r
7+XnAKbB8okMRtmn0bItpLWk0djfSc+sSZNADLGx1lopQL5c3n3oaBdVOb2Rkcrs
3ZJksjQA/MOJWYqqGy06gMpsOmSjbRGInUFiXsbQ9/5U1P2YJQCBwYRzpSJh/naJ
qwiX35/FwQ4EbVII+EDxHhWh+KJ36yqMa57MGKJ+vQ7uAo2LebuXkuGCqTGQHhGZ
W1UeQKmQbMO4zqjHZ+w1WYUeRuSTZ3nlRcwGRv4CBbg/sV6Lfig2PDeeT3O2PHQT
QZzJ2m+ODX+yv79+0nLIdZ+i7WP134yEF4j2XC/UJpBcne+8BYxUBROUTIDP9v2p
F/fXOvtkn8wtsQU9dOclCTe1OYpRTNW3UvtsGMOtnxrydX4ziZj/w5bvApjzqEMb
8eJi32YDkZ+LWThwNQF6vmP8TRZpBxWRUpfUKNLJr1mES3yJYbO5wx4qymV4OL3P
ETuTMsxV+D0B0Ms+Jso2626aAObWSryE5ZPYg1BVFx5aTJDWrMJBEj8TsYkKVgeQ
7mbbKI2kKz3Fof9WnPv9AYCG1tF9XhrIYJXt2dXPTsuFNQrii/0C4ZKNGJWnO3c+
rgFT3YbkgsHF13X6RCqZuDlqz3TGUnCJmOyYN2RKl+4L0Cg7c6rXBdMXOJO0Pm3M
/dbyjDHFzP529KCOZoVOxsD+pI0sMuFOf12TpmRD9dChpPI1EHVau4wSqEswRHLa
HddElKX18nj8u+xQ/ZWk76UDvboirU3ScmNCQlaFIMgKifB8qJ6K/KgEBQov5y/V
uLniTTAF+epbrAIF1mxJS/kJ4dBmuotb187j2um9Zv5CdKA3xlwir/xDkGU7qs02
N+sdVCIb1PbZ0c+qlbbQBhx49NqiC/gC5O1M56shjQEADrztVygDHgIYVREiHWLC
tFlPPlkP7LoW+Sfu59+t7G8gZ2QbWpkOSAOQiaVff17QR/eZtmW1aMkC0+lTESLa
0BZh5KFqwizow1q2IWHTVgAd6KchiRhyBSzhsHSeB0W318n6nK1XAwtF/HlWiQtD
vEFDd1+LxaXjtS3bIaj+mqc5xa96/r28V7s36BLrX+mqs3RisH3uyl8CD5dQZdh4
Jv2CWaEW01MqFHKW77HS3fVWp2f0JCgWpBc25gwH1MR3/RpswPeL3hAOCnJp1sAY
NE/fa7pqm3QSxmokKidwZBr9tPikkCfBEd59+fQgrPy/hvIDW5lMpkpEZ2R+AcIs
tJ0cIRHV/6yf+Iz6uA77rsMagKfMzCwZHRiacrGb3pfRBkmG0hDHvlw/+xWp5jXf
L6BxhX2am/U2TThhdJkdmw/LV42Vh22/0GeimGCzBNBthkgoDLvIEjsoZb0SGRvo
8f0CojIgJJYHHDTyK+y23KzBUWqos8oyfWmjC3Wi0VqMlBfBuyIxluuug9TISIty
SmzMcr10VmSCB01IfKFsG6Rgn+qtbw4+l4vXQXb+XW3f65egNqn4z8NQVD5gAJx5
p3R9HUFABLm0mUiwiaDTSdQ6Uxjq1DKIjN4qfsE3P9v3KC3RtXaxg/NW21DMn8zE
QutW5FxbcOrB7YqP/8+yn1rOHUPxBm3wG2ru2QzEuw1UQ5iz/J0KA79TnjAWZ6Js
cK6efzcfALzs+OTeJkOoTxzIggN8g6bi5j7XBXXz5qEPwfsxVYbNNppzz7ac1fw5
5ggX5VlJWGNQhPQR0kLe+KJG+pCVjBcDtUen+Cb0eMnE5ATUUYkAUbySJBNLSoNJ
fOLN7YDV5ClhYX+9EO9eEcwiFDFM4vN5U5YmA3Vbvg3+GPU4qg++PgndQYjTbgqT
pefREtnEV85ONR0JuJFxd4hvgUglwzj7rAcSQF86wrlkH06o8R9Nc5dgi0XWtbA6
qA0Uns+KvRB5caMJGeW01cpm4KBrNIhDKvJULj7GE+Bey59PfXz1GofAleoKeCfU
8RSfz1kVPxMSSApeTPvWkQ6b+m/tE9BVdRgY0bNJbtMsdmVM9qotKnuvHd0n4O77
Zv1gQy0KrBog367gkQUJYpnx253Dj+3evr2DbO2Qcs5j9CCIHTm1x+Bvyw6rBOeq
fLyrrmIeMhbpLtzJ8/wu8+1xGnqELwT/fnUCe1zpleaRZT/VbN4VuE/KyyZdBHLD
4n0maEQ2H+qJdSHhWTdXK1slFDqCjMQCJNBsogh6cOkqCwGHmN04QNdrHY6dsFsy
h+6mulLfwmzVS0HhWAQKy86GgwzR54QCxO7O4Y7L5yNWg6+4RqMHMMe+/0TwpeAF
wEA7522b1QhkzC+/3Iz2YogqlfQbItBbcuuHU5F/cCYAy9xH/OHdg1eSUNQ3c75z
e/HkjO8oSNgJKOLhZxUFgnSSx5Jie5htR8dofB2bZZOby8q1L21iLiUmwNKcBTrb
gsMlssOhtad9IOlnBMEqD5qIp0fzgSqLi3wZYdWc288gCtSX1bkQgdORWJBNO/nC
8FmJ0jvpF5P8MC1KP/8ycs3ffvA9LfUcqbMUCzDsu3AXlf3bxYvY2OWVvIC8wjkK
ppJvZfQXqPTqMFZIyPe6tn9PImmVeuh0MMW8ZH0kNAZhWXe0VrutPt7U+l5Sim+y
yRYMT/Pb4kg6SBEM00IEsgfYw8cbFg8d50O0xXV0zEPhTbu1MxKB1QAAMrN/m7bB
E5n1aU4djodDRUG1gOUcFGe4s+Vgt8sv7d5skE8QKjk4zbMtPAXX3ByaIsgUmP3F
3Y/ivKzmTgtU/WPWuxFIXTDZupE0TSGXWfhwb56czwGwrIsjowmiGWxiJsh1RdbF
sfedSS4UQN7r8zvL0hhnPpeinkvLjyPvvg+Z8+qjI8VcjEXD/+ksKNlr2GsB+A9a
mpZMJk4b9OKbcuPkiPfspl6jYNQwH4e7wrhJ6G5bkoWEts2fDF0EfZ5p8x3Utms1
JgbXzYy9sZYtrnbg/l8cZux5cPdnnv1u0+wBcGWCLiTls2SGcs2XthAnab4eD/PR
F/ZJ2dMelfexY/5nlSq6vIvWvCA0CHsJ9YmmsSNKRDzA4hsqOJHkrENkL/nnB3nR
9j6/VgttGCMA8G0K5zM+IVitqVQybjHlKtrij0NIT0bOQ8gyOD1LOWi2qKuwjCIx
mxLqsvdlYJko945ZTmqGlh8LxFgzrp1uJZ1wBYLVBP6olNWB8SPCY9bDuVl0dis+
Hr+Dj0UMigiY/z8cmcpnjdI2+1/fAH4hvk4XfPmvuUfYIfGxuAmZ4frlMsqn8ULE
t2o0+Rf8dQNr+s+6pKlIqwHweh2X6q0Ey1FXatidK18ijpzvdf1GmQPHNGsJI+qQ
sbgSbC0PG1W5CLkvyeInUF2AnkIkwjhTMWaOyiGZLVeQVouZbSgSatN0mCK1LfD/
aK0U2zMY8ZTI2qrDpaoRyKfkZ3AZlyug9OrKgdE3y+t2bABgLcF4hTaZAA582vYu
hZ/ZTXohOVe/bsmCZm6+gF+zhn2fiA44alBG3HKqlNPTFcj/tvt3MXtrkHstz4IY
RsT/pg/oezzPu7fwVXEejrQEOHJ0y26r6FlmqCNmZcJySBBF4g6HKvLOxKUjbD7g
TDTfZrbFP4s56XhNRTYWLczIOSE/1PcPllZ7jYBX3wXTEK87FcPDZNQbOHof+lJP
m7M/tK2RfyKj4iwDKzhkewaObhwKsr9mFBds8GNUYOhsNxA0HbYrwybVYpIOsnO0
Sl+RcFOwJUPYbDHzVK7F2eqvjzWK5QscEY0cS+ClxEcSTnU6mrFcrGl38W96zKvw
84cavumK00n4wqmM8nb+zzUkcpLQP55yhkwrOwtCr60lufz9ph9ZhXi/KOuQOtgl
W76HrdGBxX+nYsvR2cN0iLjn7DcIhJH4L56jynRATtedeFpxdf+7ehgdEGDZYlzH
g/mDjLWZO03bgGXAwsrZPoJ8eCRJBJTcr4a40e9ExRHMqVDmFIJ4hY7I5xv0828R
vcpaPZeGn0GQ0VWYemaDkydMb3Q4xsTIrzgMj1w5oq3dks40E5IgVL1KSUL8+2TC
uBFqXJU94JLmthiGWRRMNAWamnhlFukVGoHPPI1ggccbaGgbVvZGzkX2IoyT7ug4
8qIrxUcGFLdnA5vPmjYXkfwd7uFPWShdDmophL+D12JE9HB/xEfJJf4CshGyWNnH
j9P4u/8iDQqOpk4L4/LTW6hIhkm1qOaTDf+9OQRLtF9OrKu7CEHQTmRb66FV9cfx
IKhUOve1RYCCuFg17eJ9QMVH1pIxDwbznSjckFBlImAPBqmU/RZ22+93TRMoRrl7
4FmmkKOxMz6bvs1zGAkNAnvHPCjXH8xavH4iKsXHm204ByWGMx0vpem61BDvFzOd
th0CnfdHev/0F/XT3aNi7nAlY+hyT2JVio4hGbK3SO2IKHeNlkd0Xd0qkg3moPXP
aArH5TeyqwKMpAF6N6/uZ8AkXqgWr3GueU8rWPKcPx+3IqkJWLQpBP0f2SP4OcaW
64/nCW9reKsbZ/VhD6hVn6nlSvUSgAhcwSuYcqmwN6lHtiy8wBtDi35mNzBuQ/sk
v0qyl0ZQL9aYotD4RccUmo/ZSxC5nqQOQAWw6F0azjqPwNNbZXdwUhL+XugPIC8k
TTXA6yGE51j6j04Ts0MEEtcfSWqQO90y+PjLEpH3k9bpKJur7qNlryypcUya3v9Z
M8sc0qLfOc6K3KJL7cp4rUCP1mCzVKB7tUAt8nu8tyDxHSu6l9QWjvEu6HIDBT9U
rG/sa2TGLnHVbeVPoTpPjdC0O3K/IyjAJ05t8aqJSqXMmg0/3chmcd4TrlycXWwd
6syML1s+eeCSSNQTZjTamaWFlMVzL+TAYfOkx3AE/M98GQl0+b/DqdABQN1ySIiR
3NpjzkDhTR44Mswm/ON0DMmv7a2b/DYglArPDYXVLArUzMLSQuOMjauFab+oPIxr
g9UF/CkSb+/+5pjgcm+pLXbHXFCNFllJGgTqkMvlhgRUnzcGZQarzK3rVwKiMPFC
J2sxOrrUZyQWE1RE28iMzpP8AUMcs8Xole20iyiORYDhbKvs5N9Vr9Zsb5KlfD6t
A4/5ekFXrruKjffUIeW4fQMZx1VwQU+orrgonvF9R4V4t/oHMvse8hjZ3ECXndoR
s0V2wqp+Jo3ibatYMiWqYlRTUP8Cr7yxhQj/q3Dcm0tnnQ5OOHvVFDA97TIhBcy3
Zd/otu8PH+29KB32bTbEsC/MbZXDN6sFqz13jeg747fThcfgEShPinmcnMbu8ZeP
7QT+JSLWaZBZ4I+dqzxw90RlgGLog29JOpTVxxHtX6eQ+VcEsVf89hb5jOoKUZD1
RElxH7z33IcEk3fDFv5+PJXRnq3LZ9q3LHCp4E3Dflm1FBgoZVCkXYkhgInnd2JS
wTFzUDTV8nXYkdeO2B5UWa3hwoCi93SfPdfacZejyy7bdqBVMt1Zca+OJH68yAWP
LrPea6NEMoaHJRO4rwHuqs3pabbICVnu+0yUCsoqAl6w9m2uTqHDagVmH9wx/lFh
uh2Rg7fK8/vnk7vXfMwenyAV2/evK8RdpK6bYpvlkc/2Q3RHw6UQRt02RkhTivbg
mFalZfbuy91F9Hw+MscbiStsAbLUUNy8YNTdoNnY8mnsIkkg13fHeuxfZW30hC60
GNr/A5lQZp80oN7qYQcM3c5IGD1I83OCFPi5JPexAr1Dw1zBa2oxB5xyVderGtjJ
MVdI5bhS+5Qt3m65z8LzcSAmKq+J8DyzVudQdGWxGpQJbn/qiL1Gi3EtIUx47jV8
MfA/uf4K+wjiZUxHn62GemORUAdGaZPXxrSdmFPsfL/0+wcFusvJhXBdpA5EnPWe
qSr2eg7Y+5D8PoTMFuVNRuc4RCw7Y3kkHzy6uQzKGLucvcT9NpfWKz/3F7FnqHvK
Jq4XDfhUTNC0KArHvEQUiQl3Hujch6CFjJmxgLOiHma/j1ez1S5nlHoRy7OJmsbV
zZsR0Xuivds6vao6RULPfEh77wcxfj24+cVwO2Yyz59Op0TjKte6SEwpv9ReAfxR
xr0CVMfUmLouIUhXW1ZtNYASV7U/uZduttJPHJ4QrUM6lSNd3wW8/KE2WHDdN6zJ
WNb+J5tK+2fAShSepN+JS2FoFVHN4MzdYipc/n1EFPms4bFmHuivl9svq0/eoEUU
J5it8gE1eNW/AAJHuuKhXvyGkyzw2R/p+qP5fgmtTnpOEvcM5xIcOzscUrMjOb9V
XhOho69pXW//tITpqTGWTAY9cR5aSiCXwLcddidhsi4+oeImzYROl0tQewtHmrPx
f/16xGIDo+O8J+1YzT00PT/HlCArYjHA+6BmCqzAwddYg5bq/zZcBT/AYExILLty
z4qOPto9FceDHmXtuJOIDSiyQl4WxLDCcXCSsr20pZMWCzut47jlK/O18YIKhNpl
l0s2nGYbOSl52kErVERqzFNZ//MJ9mVJm7MCNgEVWv351zRicedALEXnBCIvMCOk
qKHB8Ivel76O9v64Gc6Uc6be67CZX5bRmYi3KUNQD7w+U9CxUKnnVNIVIzwWkmrS
Uavt0C/7OxJ1dBKbW8mS9CpKMc+v7P9t5zX/LyztaanZUmol1CJpnK+MxjQH722k
SsI6H8BAO2bY9eqW6pqHEkZ+Vq62Tv7jdZ+njwhJgsaOCIIrPLDWi/OArnLPZt9S
83Qbu4EV+aw8GTzh9pD47FY6gpKuIxln4rgr5gBRb3xjcXBZVimjBFnKESJUWSNk
NT0U8/+UtO528+SgIvit6jTLyNJpKmi/5yDrpKT+Yx1oygs6xnvqVpM+c9m7I5M0
UZmFX8ucrEVBgB1RSGZx+krNWbEVhnGqhAL7dO+Ew1ntBUUxbOw/CAE90juSK6Lw
aTphMgmunZVnOPmi02MMrMLLwtxHXtwgCt9zMxKcp0pwX0MLEqZpugWJ5P93p+dh
XrLWx/AFKzJNUHvv0CNtw+o5Ni/QaBuw14j+LzF7fDp5cAX8MBqKRst1oG2/f9Y0
/qS4dkrxyDMzD6esQt4sqZwbWjFK6wiyW5pe/RhnZ0mRhvI6c0roRt5JM7KkCQR3
jFmt+1VlzT66dmFB6aXsTr64/AiV3kkL1t1c4Y01fFaZOK6p0MeMT2gKqG+BTS6c
RVZS0CX3cNRnEm30IxWEOchEioRgYFuLTaBjEeLZsiO75T7SqoUJpSsboRV4FSqs
UxZks2iLZ2mYm+Ur41JdZ5Jn4UCQ3IH1KwC4KmvtEZ7GmKpRQimjI4D77R3T/q70
Qx0aFzKtcN4YXTEEN82z5m04Toe2VWru76c+/0fJ9Zsb5XFTGBEX5irhnVf5BItJ
B7XlNIMmfkqLJzJmBjT1gGobACSWp9Ya8lTlO0Rq+EgK5z9U8KXw4moA1MaufAyh
3cwMhtlBAWxiWB145LMwPrFviNnZcdZCqnDc9Li1m26qWZUuqAiOFHUhF/xEg4yd
8JFuRIqMP+bsfF+/U3RC4rVMeumZD7j9qPPgN3k5DSE/9ct4FJbhBo7FBH+Iqk9L
zjT5bC8+nV4bQJ4i4hqAWKz76aunCLxFXrTQr5ln7KrFI48Mz+xdcxZYdnjtT3eZ
UxYDCjX1mITChxg/XG6B5p5TLFGgwpaoWanZ0B/fwMg3skCkIWf9LUId3kcsiZ8+
8eMnHemLL6xJbsZ0lw9ZJDVsdFxZ7l9v5ZRteD1tgDGY17rA5+AByja5f1F8mNGX
BdmxwPehL2hduI1QNSVCFczlucdwnG7P+Ua5kyV3clrSDZS84VgYmIh0oYTSpHDI
IyuiugwTFgXKQrh1QX/KbfCA5mlGiIcMgEfhnVYzj/+9SWTl0oBaDEJ5DZYXULVg
Gm4bm/l/Bl+8jRoAPo/F7xbe6XPhdXRoxqw2GHwejz3MgvXDYf/0ffjH5Wyq8dUy
3uQ/LLhQXW8+sr8KRHWzbkfzxE9s+L1G9VuUL8Ok519TsNY/9lQYAPDqneFo40Yv
IphG6XFliJ1CZ3QhTKfBWitHIPbofE/go9znqHt71k4ZTcNoiXQog7ZICCaNMx71
7+WBDbHotvKk4gd3XipY9IyUbsyTnKV4vZW4PZdI0E+rd8yF+cUa5vt0wYaaID2Y
Xq2LJ8HVo+0A/sTtY7kBgzPj/5qC86yHGc3ZTjgm8r0voGCXe0iAkFzanLZ2/jks
7/Q9zTMvjkOr+lW5zeiC8TOMrYtMZLTfO8bZ+e/SFHfnIOPk+Y6mAguIZC3KIBGt
u5WOzBNp8MHm12Odcs0RIYdLbjFbJ3xoqWyZ0UlDMG6en/Lm2+p11cNKDUlCw+Cl
26RyD6enncAxEF7ALXzAUr2PiUej0kI/I7Y3k4EaxoRbyklIJjGzUOBF8D3DfEam
0i9f7N8KLC9IWd7fQ90rXKKYTy2tikgwvAvPvOtzaO2DVF44mVQOw1+2sDCQtsxo
6ULutUYYr9nTnwclB8MrFnooTM0oJ/4oZU3E9OhqcM4y+uQuiy6rNWQAA9UftBtG
JRvRXorbkHtMEY95FI+ZdSh33j3t97juObzDdL5DhazD0BiLmWZSrOOoA33T9qqC
YUe+x6RfoVMjE/MpFDLrEG/+Z9++rUELrVR2M/fYT2TrZe5zLfuyLSfLQAZ5DJkL
2e1O3ybNcI22eTZw2QqlLdhg4+jGOZ8nh9w0+7/ahunUq+xzJT1Uwt+nh0EhAC+j
5/sLYm6wl/ss2cuy0f3e6I6BaWISnSRFniScu6y9m1QCFNQAcWq62EPmG1PHmaMW
9bmBO6Gdd8oInVPVlLf2nUIkvb0Tn97JnNzvDbCP8WSGfCJe9Gl0koj6dCGfZllo
ydTMPFWV4a9a/0yJLCaFXTFRMr4qJjNoSYagNpzC8RlQmkRTelTXPD68aqTLSwJn
6Sk40jOXOxVimQx4lgyx/dX3rxBgDurkFU1hB9TCiJi/GENLVLlkRYbe58nx+fNE
xnz9jHodJWzrsoe1mKHVL5Cx53xjGtO+kwB0gmtuVzxhCWDF1yuG3qz0GgOzDX4Z
tk6XRCkZBfZJ15a++xEJbVDdsqaG9SmTw5d58aq3JtOdR6/axi7fHlpMffM1UKfs
Fqk8cPvWIqFVS2I/y0k+pIgkxm2k62M9AtyWjHaqfj3n/ykgQSVH/IYhpaGQFByl
7Tsrh5asYGVXQz3KWBjp0BNaOdePx06SCxsDQ+QFtwjSnvV/MdCG04GA7hHssnN3
nku/pTllGgSwQCaWXdXIe7EAM3rOH/f0TlC7ASHPPQdCT2AGHi7PeQAooSRIW05x
1EAoaQpQ+IUeMupIQt9/oSrLaO3ajfpbGkRkofxTBeM0NdyCf2VU1BiRs5E+0q4x
T6yfB2dlXgmWo8YhmFAaDBoyl+56MSGEET5/aF9c7tkwainGZ+7CX69Q97BejyU0
nfx4vTzo0XxIqvpo+LWbdMl9C8eRni9sVGhubvuNZ7G2s/m891mrYPunJyzENSWK
rJSFilhtL9/xwLZF5388zehDJmy/01adWKhrZ6wNYfYzwuDMeu+FmUapUK5PMcKL
Jgfb+wsvi8qSiNbHHvXV2g1MW3vMZmj0SYZl7npr3La8vrYa8rUwcUvG/H+B/SD5
FHWBEG6SJaLNYQ7KhzsBb196TeeXsHuDiecQ+tF37RJPfng7w1H2U1h0daIHP5Sg
Rqssto2f0V1MmEMM9pLj9QVZn71POaZjCGQWfPz/vHlV/SKrIvmE5efxegTPoUoB
E3Bfo9U7GHP+9zPESGUn15eAxEQ8a+HK4H/ydXglzpvHP34ugkVetInCE+zbhnrX
ZH4DOHnv/BX+ElKDHtmYk/t2ECcA1sYrf51u7rT8D6L02i0wSCP1oKF3jiAGvm5m
TaOJm7vfLZtLbc1fjnWlP/SzJkc8W8O0nMaGiH5VcmcEAksJ0iGlSyTRdH8cJZB5
TSD3x0lkjrYIaOdLt6GdxS8qwTsMlTFeq+7PM9s6hI2UTIrGrVe7GtJQl6zNtOCO
lCsb7K4D9wM6JGdr14qdPJBNRjGHrYhlxAmfvNa9TzZOd+SpG9tpzvsuZIV4dhHG
DJKJNEH2Wpw9Xd8nRiqLylui9QybNP7qz3Mcm8zdOsib6tjwYjoExvJxHnwGxPMx
ewiov8wBaZHEwqNFcD9QFpWCKNM1YxAtoFYr5TkBFLEVIgF48jApuW/thIAojROp
XCV2wE3Zx0GKNzfapjxJXymU3Cxc1CtNYPnqKnKSIVHsc8WJikrP5B8tz5RrCv9E
5D7RYX5Qa3z/1WHygkSsA1a7hzMMWU4T35/vGezJGwBiGWr3fzPECCYlgrXJPtnX
qbCOFW975sxlM7janKTIgZN3aw9+WjPwC7oqb2nL4ksNhc7f6thyloRQtqs1EX3Q
PkB26AWelts83VLeFbr15DwNujvgmR/Gydfwx3e2x6ENn/n3sJo9sthlCgfxB1v2
tOUGyC8/22JQBxGcFI39jVrUxtwUmZlO2cHPILpXcPCTVzjjwtH56S2vvHZKFlDL
3SEYhOohUWAs6aKVzwvYCK74Ltn/slvLDiWtLpI6ssiXjRh0YuZy6PPJiSsMls/q
g3xmlH26P8hm5h4hF06N15/bdPpWQg6OQRpPzSy2EGucRYD+p9bRZ+dKBXrx/v6j
7SJTYufs5u8k8ZTupkNlSo6MaXuiAqrODRTb3mlpybNVu01yACQoGSmMPgTJCdrI
B6RbNxDzLuXnwmGEqw0X0899lHIqIiju33FBKmRBZ8CmSnVqhgkB9mB3aP7PA/V1
FQf8vM7h5fYcoR7QQ4klMJwGYUGREO+b+etuwDYBYfvrYq4EJojJ1VlngCrZ0Unu
8RIqZlSnQkG3yuMrSiEIywUFpw5IPRfaAGEXg1dVcETR/3q0p+G5naTy0CZpWW0v
YAwHKj1tUcf8zkH2aTKFwmNA3lqqdwPod3TziikHLa84Mp5HLggezvdDpkjluc9N
VDHfAAoPHOYFuJ2WsWmoN9ozdxE8RHBZY5YrQ4de3S6k5z0KA20bgM8nCy+g4gAP
u0AOzafpW/Yjn2dlB85xBey+XtfTWYSK54FkYyBa3GDwgnKs1cA5v7AKtiLvaGP/
9UeijhIp16pq45ITRw3wqeYjslXOYEZU2Cf2dKKoPDKFeE83+flIFCJBSP+O1rGm
y8hojsmHKqpu6TVQkKy7VpY2oFBh6rtD0ecdNZTsurm4cwKGpduTU5p4uFw3vTkl
GygfWCatcBfNgwyCWDVmjjKs2kKzkdJRoj59hOXA1TQMy65ue3GQ+Tg45iyyxfGF
Ikn5gMU+mjLRQUaervqB2KrUAk4Z1+7Q1b19zMD58KgnPuV1yH5KAIOWkvRO3vXi
pD4hG/B+InNtRC76URklgtF4fwLdXZNr1jdbp7/Iz4jJMCqZc/VeOrwbnmE2i8tj
Ckyzjf9RcOwIfGARQ26+xca9Qb5cy5pdg6xwBfhAVcMar1PXQnrdmZnahselsjHB
R64DyHmnzp0aWZT45i17zxXuK3ygSmrG1Ltxv1RK2EQ8G1/YSw8Q3rj3MlaJvShV
ecXwZAyd1mPZmDutT+pp3BI1x20854eUO+Yo9Dcbs7s2Q0kNE8GuiRNs68CYRhyg
KB4C5gezZSaQDFHi4h6mEvaoUVa/qi3KdXY8bhkKpAH16hUIVrq+rrrBkl+tvA8A
YUiSd0K51ETuq5B5QArslUVwBxuZADxDEANcdDzKMdnsVqIa8q3psSA1+kDgVY0B
rY719OKyJ7lE7N0oypHDsQEKhApHXpBpBOXbD9KA2lpsgzYKqfAVW3LAztu6EDFM
gi4iRMmBCIZcsnBwiPXMnwdb59ow3ZQVGH1OcuJtha2ENIk1oudaFBiB62YQrAP0
wExoJPnxVpxmDJSMo0vCA9yQtftZNKDZMMTC3q5aUEydsqUngiIEswxcxoOYE1os
UJ3uKNIraKW0YoBA0Z9T25+2+rot+1nzci6e+DrZ/Up1IjghTDKGWtih7aj+4OWi
nP9FB3ne+ptARqADO11YySVCKMm6IzPTiw9LMYc78nkF1ibSSmTAGKtq+Udqw7fA
hgWJyWtL6V87e8dLoUHtavfqFYinwV4U/5SWS1aGiC+Siv90/wasEFQxV9hxhK5b
G2xZSsFJwtpHm2bRkWJ5ICwQRd8TZePQ/2Vv7HQLsX1gYcelEDz49ArNGInp1Cbr
LYJnVQ9dqYASbW4fJRJf7VUW7zT7uieQ1n/3OSrH1SsA1C0qGB70q6L6UExKcLfq
DC/N90WvAMxWBlR1WpeFbn2rZAeQkvsHr9oAPqv9j+WYu/ZXtnlFObMlcwBfX2lm
HtZ1DkF7GFGVaqmtEjpZNbiqzUgbp022KYtFH97uHKSz8FFm+tj20zK7KV6jGJNu
eXoYHaS/+oxT6FH/qMDddYjFY0QELOyVegbkh7lgVv6NaE9zTEf44n1BTKJslGo9
5JaN7NWT8hSLPCYw7bZubUJA8FSodfcj2XmS9kzBdBZZpiNHe3LRolZrC2r5hwsI
A+UZ8KbFS9ndtISsbJE4tB9gUZqBdorTKzkk9j6QievPpLzOiVSYX6rS1E7au+PA
uDQJXFJ4CCjDg6Ke7KwM4uM0RZE5OnFxswSQU9mNGDPXDbfjmH9lxD5j1YhpRK/W
jHtkt1YYXUqIlbbmCF9zOuFvAIzAAgcvPIAfxxzB9jjlOjny96D5yUlz+zuh6FQA
dW04e43QgOiPrK4+qonC1jiKAszFkxMgcXWMblw1PDhf47gxRZEdXFdQhdyPyJu+
XIalijfmYJaosBicvkn5z2vnwI9vzNRCLBGjq+7qRnnA1s91c6wkPhPlWhrv2ioo
UCSo+o+1XPHLO7rI0ErRTCssp2Sau6f0vFKXR66h7ThRc3K9WRgBfRSoSL5iEgsg
b/+QkA3oADl9HtLGhTEceE8h/bgqShNix2EEZJngsa98+AG3TexcnYcKI6Bp9i5t
vYWdaCTpu0QBCcOLcgA2rj9jvc7KcPPu1ZNetKU6Sg3CwwwU8hSSLqr/PjFdCb8p
KfJDi/Km0JqWfv4BzD630VO9lxEOrwduzhQc0elnYA9118is0dDZ0ZPsqbWn25K5
F+vpZg5emXf3oW96+FEmewnWuRh5K6xLwMmzIYv6DPaNgIjv5XoM6TzHJDwt/eni
RlnMwWaXUqUqHY8zjpCGbMAZaghbrSlrzsxMWI5SPZz4uh2G9lT41nMpWyPFjFpD
n6Q3acimA3o9VZXZK+LdC/jOEelXgZOPPJaxJSzgcwIHl3LJCbzkTk/+FTZfFI2A
uk3vYDz8ReZSXvbS06ZNkjGuKu+wQJGhAPVb0dk3gmm9/Owc8u4uT9HVC9loRyaO
lfpU43RthfJzm6eWST9PkDtepwUMbPRnLjCsEUtt+FNTeSedFQ7962xJEsY99aFy
XdfpcIQT1MhBFKZAVyGEDx4Wif4FV6zjKYJiqeD6XFGJT/3iYPL58iCBbmCm9hVp
WcvLGuBte6JTsgpwiwWAhuaAfDOa2p9JTvBxJd5LhN+iz5uiATXb4rBntf3F230r
DDK+kdYlvvqbZbu6jvjS+CtS/HL2hVO8MhW+FwS+z+gW9knA8IX2HcKqwg+Ruwvt
PfHnK5Dbxr6KuOj7MV4nct31dPOT2H7zqRXsPF1XHdI+Ewlp9OHsscAeYQ47s5BO
qsgvtW9mkrD/H75lfXLd+RNe9M3kWf7sXx04SIidO3SL7T61OHKNey8qnFcDTZnO
xkBqY/d7W5+XmpDDm9z/4u/trNNDr6ZdClm1r8iW1c6COq/wPoIBqoLkdOqbR8ik
pd5D8MFacKVHqA/uv2Ks5nW3K4v5QcnaX+3f7bmjLEyRTEbv5gSwbc868+fk0U0+
8hoSBFq4Q5G2hGG2o1C741nf4tVeQKzbqX7+R9Z+KG0Gl6dDIcSiavpzC5+p6XJN
Lu+uTy9eEtFQWL4n6w6GUYKlG8VN6P0NQXmp539p3YEMb3+iWwI4osJbzpKg9OUu
o4Ic9heSaXvPuxIEtTslmD9UCqwmWR1Dju6LFokmX9NJuhGU4Riuqm1gBV5BhhZ6
mSfGRT1aQxsiXzL+JYKp0zzbnoq7eQEztEccseNnmapdFPojHXxcL7/KGVr08IJ6
jzMlMik7/Pt2Zs3j+9ivugz2ctn9C74FyXTatM6YKneXwAUBwNQeMiaIbyXyKq40
iBdLaBJcBDKK/pLWKj3CXcSltyJomeT/Btb2/WEqjD+YBI8B0RMpKSHc80s5z4u8
wVCBIuzTHOPxnca0Knfx5NBhuPRKSw+iek+Yoyhv0gQ5KXUHi9LdnQKPRlo3F3Vo
64vkIPmNWe+uUObdychNgyMsl+DnrFN1l6+rVfuCQeJP/V70CYzHxlF/oiUUljn0
HaUFetorrcpb+XaVTjbp9S564FLgQA4y/ywk9saCIsimBQzUKGw+g1lkSkOP5ZcB
fyqJ9oNDy5i3rC+MtipKSqni/CxdiwVpufiNNfWVsgHULMt2gXenVnhnwJyVtD0P
D1BGf8/wZHI9+O2+k+4C5n2PQ3+leqiihdIhjdQuKeIMldLvlXjt0Xvjc1jthJjK
u66DWF+eB2bm1An76myEtyAK2T5UFuEQlZ04y8D2Vng3YuxTo2Kt+THP7NK+BeK0
CtZTuPFPWuZ/8yKNNLB++JQkZRsNVc7vK5rk2ANIFRjL/2rSkAbh1QG/O+ZuHwt8
sZlSMEdzyjKH+5yG5XAhjn0QJBZEcp68706eRMN5OhaHq3y2ktq7kCickhyCirfl
T/fJt2QqMKpZWdWQY5vtyPhFB5Cmld/TAVD9Y5p4DEBzoUmOeppG9bogirs7Rprf
kI6X9adoVy7onGtE1uPzbPpJ5ww8yESnccWi4rRi5BkgqtiM9ffx++Zn5AFKA0U6
dApTjqfq2Dkhp9aKbigdB+pp1Ete/g1wTZrI2ojkAP03Q60KIGYapHDevdmpSLb/
YE1mSBPLBRt2OUof5CgDrNjsDPJN/xoDaCTebLefsg/2IHGxAo9bOmTvM/0bKcHR
kKoWMNHkCtSVy/wSy9M/WuXCFFbspQsfZBC3BtV5ZrZRJhbXDqGA/iEjM5jmKJye
FZ0AgA2/k6fvwYcP60S/AgpYeAn7ZjRooHG6lFDOOQr4y7ekVR/V4q/aSay/+0ka
yKiXxAnWZjFFSKNIstsRBG2rdiLxtFERC+acyXNZxuC9LTC/G+Av8hqT9Qg7ndgd
SeticCFpWo+iGQYE1R67U0fhE2CrliiWnjWYLY0vSQ+LZmu0i9TkDokfqT0LsT5r
na8yanArvl5qno/ZDgpyw+klOsYBhDw7gP3oDjmQ4WpwTUGI4sKHoCFAMBb2AnQc
DhAtUk3rc8QkxvFePb5aALHCkX+1QzDJJOgFnvq3Y4ma62xXfjPqRXb395c75faJ
XIWkkckCA5+3209NdR+Gam3WqqJhgYc4wdPeJkpBObZmWHYCZQemr/qT3ZBpKzQt
BU8X7kBYw5f40gZ+TuCs+p96W4hQUE1LMMexfBxNRT1rSYDIMpL7YQD4VvCXMY9z
LEbh1Sm581N3eHPoRN85OWgoCzkhSHXOG6s9+P/4PvIY6afeTSVLYkhHJPi39LNJ
QJ26LUurGpTGTVoULtQrLFThzfrbfLoDIFc7upeCQ7+0XGIGNUz2JT9bEYT1qO+3
q8YO7BQtIMgAkGC99Y6h2vAJ5G0+JeKOpvX2add5OAS6/vNOzHkjLnHy2E/UPb8U
kU3K77QE4Q5ifYZq/wcfoXEfAquOhNUUdaJcrY1X/IrfrNRrAfblAP2xkWyzmS42
N11r6zS1+ryN0nQ/reiiwE63ZY9Hu/2iaZzFxVrr8yvWDzhoNBCiudafSdJIpK/O
iKfk7cd4D50rMHppcYxR9inbIURJAJTjf49uzoybcveG+ecND0sfw4inYGknxfVP
cl+YwzBe42xNKuli/OhiuXUSfwC/lC2ZROC45J+bdc5+PkYPoIFS/Otv47BVkHcg
PhbPaJ9zHPJXaphbq4qEokAl7atGVsQIZd9BGci02QJ7ALHPdXhtbN/0jEtSjSut
qFB2V3UXGtadi1u8+IkWYXJc04eGsKIxEXhNlnx2AIjTe56hKfYPHV8tQ4Um74fV
xMzdxIEBQILEaua+C1hS5O9WoyBSvJaFA86iI1k11+g5K2WJqXyICTizq79/KdT0
lkix+ogPhs3I7wyGmhmWDwWP9n+J71aqq7OCwXvXlq9x00hnuOVgDpbB2BJ8GNDP
SlO78dDxpx/ZK9P3fHHXB5uy3IMmuEREaSatOVtrI0IXup0m7MAddg/6Jh1tdNzR
gCmv7RLEPSiEp91B6LCQsVJPrChW6csmsWSpJT2mMuU=
`pragma protect end_protected
