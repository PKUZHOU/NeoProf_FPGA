// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
3pJcEeAwGG/44TK6FSsTMniPIpyKLSQv9omcKIUeQeBg0zsuxOROGng8o0RrvaBm
rrSGgoeahwSEZk/N5EeK5RV++e8yUxzaBdFjYSh9x4xJhPFJ2aQDhq+OrBppEqLp
ynOlCm/LNgn7aad287uliNtc+WPOdXfXVZajhgKiCXA=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 31632 )
`pragma protect data_block
vQ7UkrS0mJa1qtoFY1PvCE9uvmMqoE1hX2ut34K3RgwjbtAFuve8HYhk/ZPB6aU3
WIrAYyXvAUP9G1RrdhrMLHrwJ3ozvoiUNJzsUZKvFyC7iDG2Z1LG9SeKsmeGV2jS
O2a+VuFj3QJDD4z8kDLFKerXDrNYYtyNzf+HB9djhVnR62rdWKdUXylbUdhTe4mN
N1UzFHvfwvjQKKsR8fe7lYlfV4Ah7zauMvVzbn3C7PrA+lKHCUl/DW9DjoCpS0RA
SDF2656VGLTLBBOlXx1xn8FUodlJTeIAZAIB+dbA3xLfIPjrEtgsbF5iNoh+zXQ4
S6KyB30VlsW+iWmBdFhnlFt1Cj6NzCaw6jRqOY5XK6GvKQ1C2pqmW8YJpwK/L+kM
OvPwn175Pvp9ivgJ6Dw8VVtf8mNWTVc5GMKyLE2gtPYGQyQnRbq1jybCzCV2DOPT
5eeOeK/Iy09bvJ9O6NQABrc17JpyefXbHOjIG9Bm9cK98jnYSwT6NQX4VGbdMfWj
o6gygjsmvBPKHP01HY6W84I/w6mTovScl62Kl3D+GISR4ZutfAYsBiESMRMaXYyT
9Y8CErNVK/OrlzeRNd/jrfB2TEgZ4+PFpW9WRmuL0XhIUmNLTs0C+ToA8ghM06xR
lDf9bWR7hSc6j4B5RFuLm8mRuEoDyLNv5I3uMgex5pQaksaI5xkOKJhXi+tVUzwQ
vwkDeZvzUPw25KedgpSsc8ByYGpV5dhKrkPqSqT2P0qbx/o4YGzF4pxAYN4ixzHy
NT9RD0ZKNzNW524Cdp9UWzO03OsJEImGUJeaRwJ1afIxm4pSaZ3N95WJgWiySQ+J
T9xfqs6HxVWZFPn71DjmPtQcwwFogMpcNayRlZJbZZ2gYBNLjRJSaCxwFGLdguDd
1Bjqb3jgjUqTlORO6VWyRlooZ6vv+P0SNeGJpOaHNl6jyhAyM6cXAAWR52voQlBz
EHmVF1ktPFMAHBdbDGKh08kE/MUbWzp+bXGGH274boewIr+leQO6GlOyCam5IwSh
OIDwFBiHgN2jn2TqGqA4WoCtegg5/5jM0hsi7QXc+PPJrKi/E+E7gOuTJlw1KgDM
7gv/kSPqaGt6ZHzeO0SzBGPUAqQcIX65JLwHNYOAYOOojFc/j3/ttCQ7ZlTMyM/E
6tEHy3wbpJwHP/9JrZZLjD9bbYVlfr2FDJ0VuecQpJz1KqR5DTPw3gBcFoFTaaDB
2+SAlcIZsWNE9zEKSnEogRksTS/LOKVtnE6eIjLl5dEs3hwWEF6GRctzcCxRJaEU
xO2u1Yr6o776D5YhTOoIuRZzJGaeARYK88URTenhWZkK++W/Z/s2nkji4TFtw4cA
aVMNQcIjeuzvUHwfnIsqQhxCpVs3OZInT/JHjtTf9wobgMNeq2AJ1aywjn3akDW1
iAW406EBYvi6k35mfR3LuExwVnnyv11+7DDn8ZQJgwXSNtpGvR36wC7r3f1U1lYf
yYAVCm04V0He1c4OGQjskjFcVYGfjaDuF3A/0WbloKhVQ8uKvoqW28KxOhj3wQZI
5w6R/U8pIPtxMXJH7xItxBFeV8LgyjmsXymCfOagNOq+oFrcgc/N2wKTEbWXB/st
0z/ckEBKRo45ypxNEkoWMzCjuq6T+ozWKx6C/FGZSLzp5q5YVCwWZo9yY9yxk0BC
iEj8ku8vjP7czQL05th564G7riZKDDIA5UK3WDmCM3vXxb40BCc5A9DU5mtuf0q1
7JYp+OcjgldNSTQ/gi6u88miNqdB45ZrqoQT1DehdQyLecnpcUONpubo31vRkNof
htqS1Rh4P+RerNGkRmq1f82OKM7dt4byTyA5zHEacfL4DdzG3Y2sV85Oa4bneYD5
JcMSItZL47YAskLB7F9JFD0lUvgdWrUB2Z2ynpUgP8odBzwY25mey3imqPUyt8WK
b11Me7Ivo5fu9H8Ov/FhKB90ol0oXzulAemvtrjwMRtUJO2T70AldWZPMb3Pt6Tj
MQpItLrR/1IFtV1vRPdPSwPTQdpJYVHjPnF21R3fPeOjcbRX/sNCbspS6w5CRpvZ
vD2RMuBNnZ4ArYNGlVbMPPLt/jGc5s8twP0Rc2SZaVIK6pQR+VhEHJfag21pqvDW
PkwM2dpukw8X5hDBj3inUDj9pVLHoYfSvT3Oa/uH3waG40hYBSMnvMLOLU4z5OrA
Nm7UR0f4SQz5/8d6hDUACXT5cyJ0+peGM/yBdWr8/NaCh+88DV727WSQriSj3LUv
GkdieQsQzKSjHp6sB20woQP95Jb4AgJ7nB7k7ZroO257KCQoAubTJL2YStwU7p9N
+et6JfRjRpU7bzNzaAl9uzfSnhK8hYxmzb/pKKInArKOJC6IC8KjQcc2Ls/nWPOm
XL5vLEctWbQyv39XNyQXgp3wGi/Y5iUrglY0wcSVlgsKT4RGZfByvNazA6qxhD4X
QkPGfvqzFRp3bUr4/b9V8CqJ0Vc4QK6at/SLjdHOis99AjmbBzXoGdGuXyT4TFMe
pBhpqnDe42E87XdQaJ/kW6HzkF89cPRndHo3Vo8jPhO5AcRKO5X2K9U8PnB3LPfw
YZrR+9w23yNr1kwRER058wN42BTt6lu2hAh0w5o7VrcgkipPYeXQZ2py60X9wPHL
JOeaZv5h7E7oV5sT+/nBxI2y386p6e+N0Ry4bktIZPO8kr6JC7ULNJ2AqfdUQ2Ll
DSOofoB2wsIDsGu1e53dxY2nL7X3bkw+Iu3iY5+aLHjkcL17vdk6Q2KndL7QLwne
a0vavJnJ0aSLsFUYfRetgEG8dir7p1maF/fjg8l9/Sn40iSfE8H7D0wuHDHkfK/r
cPYr/ea/JJ8e8qXnvsv9KM5LhI9I0rZcYSY1B8HNqxHyLh5I/SlhX3vAinBj7CRf
zVObWXlE5UWIik0zVggIUuK0Cur93ZiMyo0hK2g5GqCbG99AM/8ezNwWwnOMSOrz
ypWWEOokOwjFVW7tjF3aQN5Z/MMigZVA6TDtm4Cy2d8eMBHbOJkesJLVHAvVuEwS
gBCXgBbq93hS9lTEuIysVPzO83jzgBirKEnAQEPex/bOY1nN92Olizhv/qz/zVDt
eOWJ5yUevmqBvhl1Y8n3z8RKoqK+LcyMMFyXUFpPmdPqu8p+uc1PYHFWh+MUOOFA
rlFqjfZIxwIgARjZtpoEq7TjzB2vHCtRrUCauNUZsfWPbTw40rYmbtk0aZwIyZCc
LT14Yz27FJG7Usj0NFYRkjuthi07NUf1N+aXr7C50RAZDJCxMCWKmM62Qq4iRMt4
F8/jFwNxRUK6z2RRvOJqQswbRelTAYzn1kkmmDOBX2qD/7fd0p5aDBCJy8hXzHV3
c7qJ9G3Y0UIHeQawVJVC6r61U9ZVXm61ZZ7zFtwSXJpeWQlSTmb/16NrMWFizVWI
CSbygeAL83ErAIlJG2gR7NLwPO/zKEHRpChtAWVCMRP4ljJkzmLAHUt29NIHysN2
PW5M3Wxt3JDoqU6+7EqQqSyDp9ItKxyECWjBAV+cI+s60AjXbqnwwTYpAwGiMDLr
AZwMAAUjCFnQAkLWgW+2+sQ48uEUQD5HDnawUgTcRwFOGqU1dT9bITh8V52n7Het
P3MTzvLBziia4susJpvqaUHxt9JauENZL3dCrXIkyOkvs+rAHOwqHqiYFYdUINbA
X3qMpnA5SurEIcVSJzcBjGskZxULOufnqE238alg5Vo8jUq7zBCiyeF9hsR37U7c
CzT3Rjta3HnrxPER14M61pw+gWfvF3pJS4BnJbTEmb1j/NWjyjQeUg6WU1EajdyW
v8VwgwXeTs846CA/IuYCw2bJAsi9RDTFS8N+bl25YRfVVZGR2ZoVTLCpYYE7zeun
cfiF311zk+mv2/aPZZofUAo5ZUWesj8uq4wYi8U4l1RzNJYFrVxtwiHeq9WnyhuR
2xWzxoU/tUI6olOgCBxp2DhkB6A9jzW9LbRic065o1Qp5NznarH4eqlFQBf+j7cu
L5lH5GNKUrP+/X27xqfmI/flbVGvBmVV+lnk1xettuZ18XuhXIU7bV9NSmCa8cGL
7Q/i2kDqpFu6hhcEAJW5x6hX8sTJshp4cQPtYpY+OJGdzz9zY5TaD1scsUEfkMe7
lrs2XHLQwx5k+GVJ5nun5ykhOR9Ui8ouqucSK1v5O7zjO0TBrPzoWSYdWrIXindQ
itBP23eGgLXmh05jIyqgoORqY8SO/7FzqNptFEZJFP63QZGibvljhVvaa45ssHMB
y6DVS7Vg71bhnZIcrmegcfR8Uf/xVC58bgNG0U+IYOH7dlOIAR9v4XAwWZ7yP6e+
nPvRK4luoZ1w3neD539tScH3kgEKxCWOhU7Q01Q2PZzwDOKcNYFHUjimAy6VmpMR
Tt/H+cX14wD5A1LUyeNkFvVxYUZN10A6R1NTDdp3A1LAzwmHQtUMOi3JBMwqpNyd
WtWxtOe1ySSMVzmIPvgSHmcK35MZ6KKoFK3SbevLd5YrzPyZIMCDi9oraDRTWcJW
IPKFXL5wci5e5xIwuYwvSJ1OtPtr1Z8iSz9kwD4dvRiqh+D+eI1jZSSQNR86rwMB
cGIdl42OPLkfN6zBFVJitVG2DFL7CcPrPB4Y1tBAE71CgYkT2OjlDFL52DX9HtYI
U4OwThL0c5wJk/IArqbgamCKza4cD3CQGxEYTDhC2uiuiH99xF/2B7MKDTP/b34e
ocG+n7tM4t4aYDBo+YrDFYHAM8aCD93qAQPh0dBPPVZ6Z92/WKWdrdKtIRGEtHOL
id3v2FLRrbJzBlVt4B3KsHldpMGtHIE13SodbXCuExbPn15cPDiQcikm9k7NlD9D
W/YbywFiCPmg7s+LRKEMCOHo4Cj0C0Xl1oyn0/eXWsQC/27eDpB7L/cmcw5+hB9i
o400NzZ6cviTbaosrodHJO7tGFbo3jtJ+D0AMye+506wrDqoQIoBvB1UVbhebdQK
2BHLlnNtcVmPvzgOAqqYSh2Lmg706+hQ1GiK0McI0e4oCcNGvQLxpzoQC3oViB9B
bX1burQPBGoaIq4vbdQBKRdnmHNQX50tR3NkgChsXng4V5txIIGVApgh1UrAw9C8
cRRUnlcSlaB8g1q7lQKewOCq4PLKw/mJd8S6XEljXorCMhWOykBO+DUZPzsjXuEC
culEaAMoOLjakw/+GjmUCQYFX5NHwCZfyjDWENny+qdNh5PeQuOK41+xEgOCYlJ8
DDfg5UsBR0ovR3Ms7m9MVfqoORMOoMTgd9dnVKMAQ8YCOeBS1VDcWY49LUt6uq0h
Sn3rJP2Bh++U9/8/8sPZvJ2cy33DzvgmNEbAi3jyIrR1o47khIKYTzj7hG9aRTgT
yCGVM8iXmxcZF15OAUtZ97ooduBVdagm1p2d3zlH8iVWbFg5TFIu4O6OjypfeSVv
1NfE7NRgPvKnZ6Rv8j+VfFC7iHH3Rdtj828iXfjnef1OuwoGIa9yes01G+t0vioa
9/vwi5td5ds6adDWxIIdVTyKBJWBJlRpObUyaTpFg9A6IteK43Gqr/jEmp0wGhMh
fYkFo1oS0P8Fn5IBWG4T4gZSnWqYqNo3+FsaQRXclB6jjbStJbo9vJRJYmobSZoe
eTyTz/OQD4XHz4CMbxsjTYMaR/TFnYJBF0EonzhAcx3CF3AHvExmRhbAY1j18gYp
AHewPmvtvWamD600xqzKsWtSjhNt4+5TMq/wcrL+JZuJh/PgbWOk0FMPgSDwNYiy
62/+Yr8ed7ILI7Dl8YZi+iTbXT+oQ/uHkOwYVwe6G3q7Qj/J9mFhxbP8PxNM9jgO
rNtD4lk7yScudSU88SItJBZy6z8UdOpQsTIYqIeXbTfG3nMk7e6zOVYEp86EdF8/
is/9EaiW2FP3wJ+afFdS2HpNdtS1yzqjxEccSIIc9S2Levl1C4QJV0P+vF80I0lw
LNYlDaGB/K14QeyT9ojotD43CayV8bDqBs5zjlmYPPHB6OqmyMzA3HeUr0gADIkH
EXGYN7pIDzyMQeRxHqv1ok0BvY1oG4GjrONzVLNTzHGhetLcEjUY5XkFTl7ZRvcR
de3vpVCo/onhXhUDbhH0HHDDSGLi2vqbyk5+LJjR46ytjygfkD8SdxWGaBfGPFuu
gNp/66PdcsGnCFV3xoQdMYx20w6gJjiD0fG+N7GfoLTXQ7u9PWFdRLD4ZjJtIA5s
3hdmtwpdRC1CGm2dQgJF2qTr9ir34DkY/oCYaA2cQ+4Xq2gL4iyVthkHzAmZWjmX
L0rCT6RcjSGE0JbAXYWG8m6sAV+6sgQDN4Y47gvF7wgKq8nfZggCFbtYRcqm0m30
OpGb+x5zXtHQTi341u1LcTs/2WtYCBxo/zJ91HflIN/ufcA4tQnT7MF6hEWp/kbN
fKNJIyY3OZjsed68rGpzBXjbgMxUkUYS5YDLyZ7w8lJBZ6Jwo8uQrli2aurOThEk
R7yNt4QF9m7TXznPrEhl3AfK2Gf8JXt2AS2+aXF70gp6czG/ZJKTYJWI9cIem2+R
PD9veK0hjqe1f45tQGcHV9uTAZc0c/HQeXiowsGM72HheWyj+me5gg0FrryG8WSu
mxNbOlO6/pNkyli0GHSRPkNuWRorGTRhIklCf/sVtIDzOtPmGzIeM243fx5LuFtS
8O/3fGX6AUGRouripeqi4vIZeyqlmk5JPCaK/6d85bh0yoR6SwO+L9qO7fFdMRwV
va/Lo1qn9SpdVtzyfPYQ4Y5ZmziAF3ImmchfHLUtEUdV5J4Dzrd2WbsJv2uGVgdG
ifQiYkRLQsXXyT7AoEyaSlxfD8xuOeuKRQdK7Qs8hs9ehCJgiNSfkNXd48GVdblm
7eBpuHv9PQD2mQg/mN2h/KrDZopsG51SR3v+ExBvSHH4++/GM1KUmjo+fjOpGxa/
MCmzWIDapePqM4J9SwNyBc8qFnoIxT6sB07tbD6clOroNQWQv0/0ISwtnvDys28v
G0pKhH9Z5chvlDHJOfX3RGw2EnTTjMzgMNdFuypJXLmCe1DnxqRZIoRbg1RnJFLb
59YinLvDmHCbf3SUj96tmRnNmwWdjL+vy/UWs0jB4eZBiVvRCKc5lP52naRjhLFD
Gv3BNGTC9ck9EjoWQDkggoZvvbk4MhNU6avbp44JzMhLwEnQc155reCDLTItTkVP
ORKKyJZQZUFbQbJXYQSqAgkAQbJbu0Xg23NhypgJLZm/hbbIZZj3xYUwd+SdWrhO
y901EXz5xVYoEQ35ukLmJznUJcazF5uzWId2zjcSvAVaKYTSyWg+LNshewg5nk3G
Ebqqyq6BtlMfSkstZAYTbzsMhSkUoBJsL2YhTCzmJBKwcrsDqYeCZeZ9O0LFOZE/
5Ln+4dOkvjCAtXO71ACJsGhsv7Erhe37lhRLcOLP3le0Bx5muvulauxfqwE9skac
YpFgoZ7aDUW1GAC8EtHEFJHIYqkaiqU/oTKLDTt1GOb487FoeYZAEHpseLGgPfY8
1015QvVTkfoCMPft+Q3fYYA1FZIKxZNlTU9NM61AwQZ5M0MQttZPbE7BgaS5qm1A
dCI8kCAZJc7wrJ8/2Ckgivu6EHv5coLauLSSsBbaH5cyKxXxL7Awrpzogu8IUSLZ
WWVNRpXd8DxqizZIZ2NOcuc5A9GxgI7U0/CR2MlpWen/gkF5ISu3TuRHzJ6JwmN5
rRG3WwEOzBrxbZ/q7pA/106XTK8dGlgmFtVma7DnjNCs4pZvRMn3GOkwvqD+SPhJ
achiUhmPI3/Q1jCi2UfhKynF9M4s+bhi9kBZs1XeuXv7PeVmqTGn0HAuYW9u3QxD
+B9LPK0Rd4R9q9bJ8lTM8y/CEUn7PHyqd4vrM5WOSOJeLZuQvT5L6MRG1ZzfVkj6
2Q05BlD1f+Ds9IsyPT5mTHk4LSOniZPaW2EIbX2xIZd/JLqRc/pS2LvNQCTBHQXj
w4m60f4LW71ZDS9+plRcf7LcYPflVeDSJ7KhZIODnRutxZ0FF53Cj939hC55Cy9q
ZDiQ2jYvo/tKumjO8R+Na2GvHReP9wii8fupJ/6rg0IYxw4DeUpWbL9+d+CnzimN
JGPdHAyhrW3cPhkQdWXQwy70OLVL1pMeJeIvDqEKtioqf+uAAQ2jd6c+BXGlTFCQ
Hvl7LpwHJpKFcChm1hqakjGH+Ch96ezguaj7u9K3wxZpoZHiEDp3bQYSIqPPnCwb
pqNtYmqUbY2ItMLmTYimEdY1JZGaOS+SNoOvfXtSBEanIvPW6HGMeE4ll4LKnVpO
+YzpjOVq/lnW45f7wFEKSZ/oom3XzeO1UFi9y6Ngde99jzEywc0Uo1VXdB1DtWfp
QhC62XQyIPdWYTkH28dPNdR5HbZ6z8GWcx7bxiIQq+tdZ92nsroLpk6GHcoiFYLG
/SIZC+CfcvE3w4hIJVK100sJ0QJ5OpGM7l+ZDny8D90QpV1cfIZFjR8aqLcJ6rdM
OMEPjKLNlPQ5L6/pdO6oy0NKNlc3zDoprS/1ybpvVUfprYS1eaPXD/ScnwTI9oHT
8nelOH7BbY5G8iUoZJztg9NmDP8J+eBkr1WNV0oEl2/CjStWs2Gc/taIjW4TSSsQ
A2YcQ0FB+USFD2MTmrXy3F2Gbnw9sU64HdggNiFpiNAMiIwCZ5njJRW/8luQa16S
JNBvVjkbfGaCTUV+iu9awBl6kI4eR2kORg+lEJoG1bdehVvk5RI6ke4LJN2OFfMe
znpsBcFdKggOc4rmqTPBqRkIVmhq2n4suSvEkntnbIkLTGKEsPyN7HE6iaXIq9QZ
1dmoRrpL8iO6JUpxhNWxoKMUj3K55t2Bs6VWI1+rnCgzVEI1oN9IqNnCPKBZmzAH
HCqi9+DO6vbi4hMbV+qnxfHYfCKKQbEvyZ53MtYnhZlTNv1IlHOj9178ngzEkXww
iUzg0IRqqatAuFh0CpLML6m7wy0WJmecg0X9VMOA2/mG2umnraqyOcovuIaOpIdg
o+zKQJLFH87jyPMlZT9HHRVHqF+X3Q6j8orJXswQ7hf6bLwOtGxNTspL79B+9Yq0
gIMuxLtAmYxnaQryeIZNOHaKC0yDooLEdSloRwkmDzGLwtsm1LUvSdR0kMzsgzVg
hXV7h+oEhf3tHib741U2M0CY9FXrnFAO18PplbJh8gvPd8NYwGwWOyDAdV8r85YO
d6R/KGu9zqXOPAMgVlukOEZqQQthvEzWX6wexJA9HP+bk4bC7sU3AJ/kNkki24KJ
/hfPEIlVSEk9XC9hzL0g5/+Z6CzaYEBj5PcmpAOasgxuySj9yhjq9PQrnX8JWzD6
VFrpERrCjbiWovnrL0bOQUM2toQvQFJ350+Ej03184Ej2YPX0jpxzTKuPPJIZ8n9
bdnOuMoX4CerJRH3DnItP2QFuRjt7nzxrgXjB8qJ0GHW4W7Vd+kMdsaKK9C4LO6t
buNpy8H+dBACqH1vzNK5J7p8TZvLjoAZxQqYQdJ0qpdiU6H/BjmTSmW9KCFZis3a
ml8t2ZHVnT2sGnR7dRPvYGmxYUEBcy95J8Edpqhj14jzeTSPDiMIys2H22f4zVzG
scC2BB7KGGObaEF7OPaz6I1tDgz0fyR2bJqVuZWC7ZZgZpJWk9BEu6lMM2WyW1am
sz6LnD0aM5fluv0l4zRhnDkPvAVJbModTevfYzdjjtcA42JgJpjvHbOhDXKn/oWB
DsHoPyv9RCqwcrpJVPII2Ccs7ep5+y1lUzXUrbrnjRsdsd0J3hJOTtYSfEAmv4qS
D1Apaw04FxD9sUFrY0QYJPz6dX/JzuuKn1cOnM7aem1kgqgQjPNAgNs7FeHx+CFg
7f0O+f/wLgUf+HE5BaFjTSBe/RwXdAAViSD4pVA/9iV5Acw5lU99ruLx86IW3d+z
xqTAq091Biss1Xz3Jpwntd4aByepWEsBHEZHwCX8N/U/fYiuZEMbZhIynPV/6nMB
O7STIEhtvELh+WMXGAI907zp/Rio2yWuWLgHzfPx9I5vtLt9PfRU2FwVwk0RCCi6
enSd4KZ6kkrCZnxCEYoEu3R+a9qQ7dbeG7iwtxWIfR5fg+3Y/Uqe90OX7FKjbY10
SnIW+5xyatQr9vHhRrxvh1yrBKJpFCZ6OiJPJnRzruUNBpYZJnKE8f3MKpGZ9odU
CtUKK9Kzf1nOtUBGGdJApvCCBuuhfPdpwMribov8yU/Wuzyz9GTtkFoOng9G/eG7
epHw2zvp9iLqbQFYM61yRc4QNScp6kR5nWTbGFKxDeNejsknua3Di1zlWko79Wi7
skQbUCGpY+cfZLpk5vQMhGB0AmPFj2t/aF+cuSf0HW21ZBeavMzrkkIuq8fpy2YV
zTd6cfLv7hHmFHL2A9tWqaHQqXkuKrjaDMbaRZQcqahM/YF5WDkmRWAn+VAetYk/
Yi3/s5qafT/rMt9L3QxliqB3b6f8T9D6Gav3Yk+VjAAZDngCA9uh/zlVQsDwwqIY
3hDyxb93ScNiY/xeaD2kZ9tj9zwbJ+xuFANwD0bAGjC09k5EBLmPzdZZz8x739AN
FaNo1zjxOIiPjhz+BojlBX4PT9lj04PXBCmEb7WN0NzBtcO9+So68XrpreKA+hKw
RUYeB55lHj9pH6uJQmOY9hff6NW5lkjhLYVw1HvdnAa9a/uzeaB5ayhvYTSPu3mA
0RBJnlpL+RR017HDTbzcVioMb4SfAVrvMpyyt7q0TakyQLNsHSShKSqBYkfkgzBN
EFihFiyGmadJRecg7wVH7IXPxrxQh/ExB+QX16OcVj9dKo9hlmkLg3rx4G1j/+8m
2/unW5SDkMwbSUYVYvIjCCpOSAO/QJ/kKoiNBF8GM0wAFd5VUiABEFCcTktqUkae
76hzil0+PFohOBX317QdI0Tku2MaROCm/TiH6YQBIAid3cm1DIGAKnjQ3fGwlOY/
te8uRgYxZHP3Bgrjoqgk4bDAzV1NOix2xCB00Qr1bdrUBjsXg9beRnB+Uj/comUJ
11MVu6on+6JG8pGOZ9WvGxib9RlUxmhtc7gTs5S5GjOA1cFJvrnDRmDdSpQAWt92
EPWbFsi59T2jl1qOl4/ZEr3e9TcOuDzudk/9e6+cITL64I9bk5NZ7y4XW91Ed9Sc
b23GPpBwQONdHrzp+olxoT4DZaStPE+kypHRLC87HzcZxt9eL924G4Eu1dr2/Tk+
4QWWHqXNcWqpto9QWO+zARHrh5X330Y8vy8lgCbC7MZSQsC6s6Txh2C6LPmWnlcd
zEI0TkGDBNalFjIFjgxhvZ3Pb0Zeug3j8c7atSBwgOsgmn9hJf7vCToEKo2hFYGN
gLYlX/stWs84gFpiOhBKBmEspVNVs6Z6rjKkmPaeO9YW5jhgb5AVogq9UEwQkNpD
T2kQLPWx71JK30UuJ+fOb0rPmRKnUrkM13MbajdT44fghKSTM2Z+KQ7r9991BK1a
C2NUTb428cl30CuqbOv0IYFkulnDEwXUHX0yAfrS8WcHttPmgSDOXs/Cbb/b9MST
1Vcel5+l9A/e7b6fq8CzoFRG7XXg+pfVYvJdM1oqKxRoGjL+YTyCGbvCS3O1lsW2
LKoCeVGftIMCYtkE/YPdvGhyTZj9t8CZzZ7BUwV6Psf9kW79VhoK+wUQv6ULJoeB
vKPl5yzBdjfnZYyHVpfRKM6c7Ttsmb46LVMY6BeX1K9oSiFwhf0JucxNkEMf9BBQ
3cMlpOfrE6vPlqL5XJknWwKrEt8Rzbti9cWXdIjyGLetZQJi7Dds/lRDjbq+Z8T+
I3JVRsE5cwUtcsKLGRsYqz+LGviZcIJzqVqBtmt7xxZ/HudgbFHvPMHv9FDslR5E
ubgxupBBeaX5MzPyClbjjYZgQpOo5L4ul00GlM40otOCrMMzBOQRpOrMsLchDrrd
1cB6CbVUVsZx27ifs75LYdsHczKujvnb00IZQWzKOTdmqx3vXf9a6SZu/VFLsdAn
3BxgwjLeNLLphwrKPLC+3/t9204CoBEzBz1vQ93PyJLQm4qt9J0L0FX7RPrTHLDz
6yFtK2LjHmlYdDcftg+jEL8TT4SGIEqHBJbRB3SYI5I7uyF16ct8PCvhltHfp6ZA
iVNZ2aK+i2HtM2pStWOqWd88omSGqclgU19+A6Z5bL1X49K31AfthshrkUHQpS7O
04+t5wvt41LMK9+Bct5qAmnG5ijOXSP/pSz0P0Y97jmogU19ex52gskkT01yvLrA
SoZI8VlwmLxrTQVOJH+zettAIjZFJ75gi7okRM7wOBbFCelyu8n+r2sIOIWpD1t1
QdFTu8xcaLcSmmm9wHBbicEhgYAyC9zM9Jy0M8kL9s8Z0HnN2bPZAl5Kz1cNy4C+
B6oM/EKd2wsRJVoY0Gf3027cecWxd1HVSZK6WDcYkhzFxmRS3RBL+iywINkmbNp7
wbq9jcaDRNev0tmXzBrzIzRzwbsS4aG5Dku7ssAuGSzOuAMU3VxJFYbPxWFRgpMO
g6ALYqJ5FRyaV6x6cNz5mkLy/Yx4E2fBh/BYy68AiIENuhjjhaeUBlC9WMZZuTRm
UYDk+uxC5Id37Koe+e6LBmk88SQP6sv+XsU0PdoSlvUXB7JX1cqIaIpuBuHLDuF4
BSLAryz9jfyP6pyVCCKdDI85YdlUFP+XaelWNijyuCOzThUzeCDKtXTksqZbCgtx
8WHE2vv0HzjfyEVGFlxjNa+Qr3KKYKDqMgJUAjb/od5FkJtqt9DVkUI91pV6BI0y
YX/T+DZv2qcFEd8ZSCo5uy2X3VEn/xLiuAiK+HS21trcnv6ewh7Ui7hQBOQMpszy
44mjZGSiXKMfJSYYaZu/rmbS36SwQ8tIS3i+a6Fhl1JKjxAufTtkBEgEpM7EXdUG
Rzbd+2+Qy10Dffadbnsc0iaJ/rPXZXG+FlfiaLCC2Qpib3rJGK7P434C/ezsiHFm
gQbH8RoLp3oON3N/Sffhb62CQEcTgoeGmNEwDhFagnIaXsXTxbhu3RehmrMCp8LM
A0/TmTK/n4wDbSQ8GVA5h4tnYIxmUrH2egQFeQxWJAMatTlHt/d6uDUe1hH9uePA
cSFgyzif1oXELFlj9YsDQRVNuLmPAYgu+Y5mAMSl2t2jiRUYPAeIit2uhEwZyWat
DOe/2VzhmfZNXJTGF4/JIONhjXXaA+vgsmtJ/yNs8pP7Lp+GHDgMIXXsqxS5ZqrF
FWzzjMv8B4tWc/ZxTMB7Q3HM+Nyy8loK83CSX8omxKbNbeGhIn/lXUHpgcfz1rx5
Lj8oEseWHO7hUuo2LhD+1HQn76cZOR0gtfrRDY2j+5xu+wYX0/jIWtLs9pzNk5kk
7/3JxbIR0ehE+yGTg7DTJS+b876F6IGK80G0ZLj/x3kHDFrkRO1IWgWloq0t5+GB
Vj1GB9eiMJVYoU7SUKzzB7yeVt+RaOI3ZQIzzSiyTd/r57+4Px57+AYiozkjLV2e
csgGPwM7+Liu9AApgUfEVNbh/Q4ATmRdUos6k++F7SeEOqHBdNbRit3uG1ipVM8H
1mzfCc3QGqqLK5hqIcCfXcEKzYqj9cjrXfwfXy+HAdmkOza+I9qgdEibYM/y3G3Q
mYQmEIZ2K7TZV5+6rIRo1JtQMsLEpx1DtE6naigS0h0RrDsSfximoc6N7TsQv6ys
2NwEL87EiyxFQcbpXhwvPvgOOQk2z4E+7/K3dF4UAqDa2bCqu5pAeBKyA0QxBUgo
QiOjHXRFwAuk1iW+GdaK8kkHgJpWR/qRs22F+crJ6VwNYS1iIy+qgwQQlNh6WiMH
u1UD2svTPbQgBgQH1VPmlIoxGDzYdkz22+gpes0t9T9OHGdnvaAcjrhEaFyWQl16
ERZEzcHVMv1sgi1oDuMD6KjFUs3KSqxfTm6Z0RHSr6c+sdc1UqJTIvruR0dldnnO
SbxdJO1+hyM+X8mEptZOpJl05UcEg9Y5/7MQJL60cp/+DNrMvMouInEzhzd9NmC/
obnVppT9aFYxh42x3NbvE/QGLLm82nQd1nCD/3sslJ/jV/nkZ22tFVDhrTMvc6Cb
Y1F6wmrivU3G3TEmHtzae0SK0r7s7Br3NkzJ2f2tQKJ9+zMcgXFsQ6s3Od+UP3bO
AObdXC6dKtkWaUldzoZlQ9Gq9s3xWlM3Hd3PA+fq2FfqxXC9SSgwyguxZ+6PmUli
bMXoyXuSgoUSju7z8vjuL0vlQ+DK4QnXZjJW2VhBdPwIKr+80kVQfhWlVZUX4Ivn
zAIZdzSb5ZOuclFgam6xQqY/sDq2TBN2EkJKrvJhy2Y1nroWhy5TL8KE5uUu53VY
7BklKlgML5xIVFSkCAvEJs6eozDtqrqS2ar2N4vWhY1pmR1V9fdyBM7ZhKj2UcAg
XYNYr/9u+a4Zl2v54c7t9baneaBTJ8UTSE376ereyXabbso97QzBXbwwRHguRMBd
6bnJVp0jQMzrdc2Ocgx0N4OEPFvLQYZksh/qVZ4AHCB4DnCmSY0tochcmjVoVm3b
GkRO2dkeh0cpWYHrO+iAgu8USsdONmijDRZv8xLFcJOZIU5XMwsnhHBkjunwB3cz
tHQl4TqryZNQFEyzxobyggjJI4EHiptTaU7rof29FFsAOb/kU5Fz3BgJhTqBnrVT
oRPeOih5n5DZVUmP6/w2JinnOk6TeSwb7T10U8WRLm4s0XPwZO1GZHOx4HpVyD0Q
yVvyD1VSJu8y1t8c3KkXQuazoNZePZkNg51YevCJS2xuzwMZBxWf5fQAKscJzNVF
IZ/ZfsWxNqCsOaXc3x1DTKw0hexfVKdMfIUDTj4fSxxrqDsAqfbn3fJCavzr5XiJ
es3cNHrVqeDUNV22+G9jwyfXeCWXbxHAFYWOmBf8KNA+b/XoNi9jupjX0BLQ/KmG
FA98u+8seAfaScvRns+Ts6ILxZH4aXC793pDyWN592XYwwaE/4sDPuaEo1sgG+mn
xbLdxDNGgcwqfHg3M9RzXgVfCv49FiC2jAnWBMelD4GvrkOZU5DUq+4IHG0iYHWy
LWon8ZiU0ao0qvsGvvO5rH2k0b0+R6VPXBfWSbY6ikpOUZCudLXy2t9b/szJqokN
DEaaHFIEySsD9q8YzqeUVYTx85uqcp8pVMArEIll/Miev6n9JJHQcEwEFcjHMiOY
BWHODqLfI85cllet3octw/SfrNAK/9tgUCaumY6h+bv0F3zjob5ImVKUDQVxNlSQ
NInRPYkpAg4KuYR93xwpYxULIih9yrdiS7BPKak2jOrjiEAWZfREG6choFSL8+Gs
JewsWU54iMpGC66A1Q66XtVyVT1B+VRlF0ow9z2wKzdxeEtIAVUAtVkDBs3JhyDh
E1fgKeM7rMT981w3Vb8s9kR8/DFHV1AXs8iQUEPn+IE+9gUSeWWWKJmIsCvETDYY
fLPQYrLIm9vSIoSld0CPZMQKRUsGzIfgeNMe9p+1ehATSjlsmi+4vupA8foA01qK
5EimOPTfISCeXHUmUUxh/YHsz2UW3v42BQCtA2n9YBLmUZ7ZlNA9iGaNu29W/Iec
vfeHFJuE0pcJyOzcuXCWhmknL2tKeMnAj+E8GPJaE+SKVmyPEsEOB2QagGcH6Gky
gZj6+iJHw4ciyxT1xY/ZcnniBI/3UBYzxGEdiJ2crfYHADwSq6NnQG2uJNbFVgO7
sYnzF7c6mXn8CkoFIk4voqtE7PK0eat/4aG7ag0T4kDLEvzryyjjI9+aA8VX0jbG
2Vk56Ldc00xzoQqIdBj5IXwjisVYug39bA6GkbG9kvDnHL/pp37EVUxv9ocN6Lvk
JfEuedKX1dmonOC4mBOfVBUopchFShLy6qmrqe3AVLQUgKOb1uZaTx9yDnPqCH53
9evlAUhgFFh6kwZtAxWZzVgDA82Vc8uTrt9zyPMFeGnUpeUTlUwl89Y6kBxvz9/f
CYXimNEYiIIfCxKd+V1Ah8nBpUYi9Y0V/maTp9OoQmEwiTDhvSAeIQedA2Nl1hJc
5uKkojze9KzPvJFohrtPwuKZeBvIf7eGJjwbc8XdfmSRrVMCgVvP7q4QH1/mwVxd
qkh9aDqClu9DLGc01I37gcBtV3Cq1zgoFwCSd8t9gkg8QrvMlzpR3mTimYIFhm3M
KezKq72ePjXkaNP1UxSlgEWplcAU8F5v0hgUyfjuVt86xata37wVkyAwPsCqX8/g
isv/8bJgrLnfIxYtP20IzVIr7ZNI+8D8v7N2F6TUyZ066LJW9yw3BUHHhlLsSS7l
UgyNOqQPtn/uDjz195xPvyKu9SVA1ggt7t2nRZsNEn4ARpwc7oH1LSXH4nxDTiag
D+ePaIZvFXu+bXnvG4MRRIDIAEEngGcPfE+ZM+DXYvdTF512yecwN4Ani0vhZSIb
1cdm4DDo/muQlSFA7egK07IH8jSmqprpMdYzBlPq9VfNntcpYydnXDYgiI2vI717
B8OhFzG+ozlPX+TxL1P72oFqV1WKNbDnmGN/zW6lhRU0KNPJVbNqArMvoOPHCxpZ
wW/amzdmg6+0KitUx6ZYu0x5N9Gjd2S9tzFxuSYIuj2IL1r8F5/73SJkHD2dbxst
3XlVoBF8aVbybYM8pIOyFCSQaCSiSnPr63ugjlOY9IQLIwRyYWnDokmkBDneihc/
sW1wJEU8RbWdCzOyvzodhosBoiezJolEf6tvYGs7xRjaqIB7uyCMvh6WWmM/LAvr
TD+sgB1lJWIovQYu8z4IIOsJVQTV4amoP/dXeo/hJlROWI1erG3I8fJgwkksCSN/
BtFstTcsChi4nt2y3Mj7gSPAyYNA4QQ+3XDbycD3BW0cGPtJTNUNMOAlzD9vrQA8
S7Clf8g9AHjjrr/BWNc0Xkd12SnreuTlUhcIV+/xnixijbIWqCW11MGEvmfwRQHA
9GGVe6lI44b20vzAmDbVMKTISrZvAkAjsmvxv/VTjcwSvKvtIHgrIGtSj+CcM/6P
gvtnC8zFLG4wLdYIkBer7NtQxpyWfFE0b55eBxLZkBkuwfJQrBg7bRmIyruGCbz5
90eLfYOj++S4SmV+cbTqveEZa0P6HAz89F9ZnaesnJvN7BEWUoCPG8EbvaBAt2uh
xoKXrBr2RIwwK3Fjb79hCG6JYIZ99JdwI5moWhYgCK4mYN4pLHqgUKQ4in8+ipFi
wMgAuSF7gB0kT+4NxkGKpZWy12illLp1LlK1L0LzJc1wy8iW0Vz5nMXVm23r51PU
afiIgJBf1/x8QEAtoSn6fgDuay9e+qAOCNmdTwK8j3+/x/12G+BOhjtcKPfSdhgJ
/k1H3+cZvarpHNqHL6asDPT8JprQ+506cKiHUevXG0Pxspw4GcBa0F4irebr8uYg
TxsKIGt46syW3ez0EzNwKwDELixpkiaqE0zcAkzD8fhCpSCeekRCyOz/OGzDDpQd
Kbf7iM/hI/7hK4HEAUk5VlJuvRAlgJfv8YUnZDhmNcU5JC/q0p1by7m02O6M8gRt
ZWuPOPNtWcUV9my9Bm51byLpjw2Mpp+GyfrsRZU1j62OweqZmZSUsdg6CRor4tCy
veypD9r7Y21Z3f1cLGXfKkmBhmYznXSyDiFt2G5XKNxR0ioQQsoxN9ifoeaIuwFF
8imgGQYLKFGQjVo5frxzYYYPAwJM6h0v8S2RcxTsQK/8dISFC1s25/gqqRpZaZEz
zxjdrHHhmXbaw7g8WJvgxUvIipzcUoBDQMyT9FaAAckvtWHKFFuzkIbXls/JhII6
gIyNaMFY2oHr1BSdMlIG9SvXIbW7+wEqRo8ZSZZXg1YgXPejdfFFbqOTkYUQJ2Ux
8KrYEcFuyBFCXQHYs6yPrboiMtSDPQx1u90ygN7pymMIg93UGPmzdpvj1kgzyfIY
uCCr3fJXqgckRoajJCa+OJQS9jLN7E9JAsfSXAzpGyp0yf+g65JmAwc6Io4bWe7n
tJuAbSSTlD96RbmcEhiC4v0jVRFz+9+HZLSHgqyR7qBJW6JYJdK+J+/qXIuJJSf+
7pjyjixg/a8ueRxidk/aRRAy5tC3MmbbMwDZx9UpDI944j+T75CiPDXxM0MULbVq
QxJxxdfP7+Rpx88XE82BwAC+baUiCkjeF4xWwVuXDg6qv6aGFdEQkC972UuyND+6
BtpreKow2hrwD8Z43ytES8UjIx97FcZ3G1YJPhnCFzWIU50ThYUUlfvIs0yXxeai
CDmomlUf9FrxHvcmka3qyy9zLLJzpZ9jiu8sQ6hd/nd2Yfg0kqjzLz5lqoXjocmd
p+IadKrlZtuix2dK/cEL38BrtCsiwqmVD8pwldlAssEkGH65m06rcEC5tp3rFPSR
U7sg+iegDNtlnHBrnwsbJVDjNmkKp2HSyMJ27PSykQmbZzHTayJvjBdk/6/QCgCQ
bC5qCM+KhVZmR9hppNHYF6/MDA0Ds2RYuBZkZXAMCcJdc1lunbXfJ0giV7rlvK2M
TtwkBapOVunww7IiDnI6vKv0YW2g6F4swGpcecHskNTXrGeg4BIILNLHdQOjZd9g
Sh/gWUuxD/X2ofxyM6kFyigTsmHueHRcugtw3ry7awAXHikuH3YtG0T2EbkFqD5t
L+bdBtFOJtM1NLKqAwlytQr0rVbl4XnPrQMB5PZrrIwtAsqKEGgSH+1MPT0RqUXx
eVF0Bf1CenCn0z4PpfjdnWDS9JDxOagGIUIqHjUwhvXgou/Y6EZWTKQUw5uv2pXx
ALQ+xtalCp4DLe3btynjQX/5aetNh45ToKrHJ09M+tk++fTUag6ScN7+zq+Ym/GO
AnLZt7Bs1cr7VRVADFJeZk10DHwkTG8uN92Xekqw4zzB1hjAPE9twj8k6WpO5h15
UoFOTy7+Cl1WathWzqC2VhfCVS7J5I02sS6KC+kqFIRkWh8zjIo0Be/x/gBSUBT1
i/JjJaDWp6yV7ujEaJWSolSTasLCrGO6hSY/9JSkY8aPOYsLbt2kLwsBlWoLz20+
3E1z0k5/gozy3oBxemIoEnNETF6mBpLuxH/zY59bxHLztqoKQQVIGDcy9fYrFPyC
peCJnpmO49/OS6YKbd77rykr81i2DU3+rXlTMMxot9ztaLhZv6p9pe4Md+PGWXQo
1LVRE00CdkayeEtw0c+vwCTd9tzwQ7DmJmSqbKTvHbucymoC2pZoYpIwh5PiJslr
CT8a0ObSRp6wxeGZR5LbS253YaF0A2xG44h3OWGGLiJuJWhULv3VabKKmbW3rYMI
lImDyp/GlqqwOy2P4ZmwnPH5Glboscq6OYnKZq2WSnXmfwtzGLmAaeXh+MW1NWpF
nlNGnoM58YKLsGtbh7F2So3aw7UujsnfbLltVh86QUmG4BWoel1ok8WVvoh1bQBd
HkfotA9MQYX9taw1AuxG/bp8+gRRZCykw5Ns2D2DNm1ydBGOUOBbLprWSHmQ4G6y
SVg24emIh3BPomJD33lQmNDZYlQ8ZDTJ1TqhrlvbXuLjYHUaFWX0l5AUmZaEle9U
EAFQvBpXrTFlhvakwocn+4nV7K/Sgz0IUJUJT/MjtQfD9f5XQttgJVYR7CJv2oCI
yae7Q+8b47VCkr8GOxH2DSlNwQvu2Un2cmw6vyP2gbaDVD1jueKhjWU2fIOIjckb
Akuc8E/3FWxeaLA7+z1SDZZiJYa6HQqxYmgSiVEp9o/aWL1dYnGuKQ+bEPqKFXv7
jmOP9PGMR0itboKhC5yMY9ct92YisFLnsQ9a0Lf8v+ImBrXC3GMOiAXE/noNNqet
IgcgXyjFz0HrZcK78+GR+JdfFOTHxZKvczh8T+Bnx5p/4eY7nnkPf3qBXcX73cLQ
sv1D1EdK0TayhgQlafnt4/VjlKfTAtQWTFJ0ty5srOb+ph6oajYGoLsQtQlTmP62
y+soGoUwA1m/9cqjdWdTiDiejgoKH4eVdiLzG4ZzEpvMW6E6zOaPfDvDLGR7BTQD
x4vGK/2neh4mnkUXcUJdNr6WnWgLRHp+cp8PcDY0LoXHNXuxP7XCAuCznBD24r+B
6uRtLesNJaQqHa7XrcQJjElQKdpl/150YPx399R/CWqQL9/RI8Jw88AJRdem617+
nl9EXnF+wn37nOK4WMyZ0ueWQrTQp8lXWQrBHu94TIfsrb/LwiQqMLNAbe06sJ2T
+A7DjdOQJTXscxyCWRtxjRH988ddp8Kfzbrd/U5cWMBlPPUMR3saVXn41igQY5BX
JtpJSdjXWs7H0xDX3vativg9PNE7LiWb0xnGDFlKiMzekS9zr4lYCsiNGpJZP/M0
XXqBUQN/6Uvi/5yn9AkBs7q4CNdqVSjkH3MRj08MLSXbBQuGKxnGG2qx0zeMNJ5H
+FgVQldkZWAh95PPLiuQ4/jQ3mVVFGHJ9dkFDxHjo2HesfsP4x5yZPoU7IkO48nc
iLBh52vhsWZIZP80+js6nLdKPqUy/HfO6sgYk5UA2dMOAdoQqC5WPD3jYH6FufWS
6ARqxK20AUum1pVK6EwqFdM6qTSMT/POayH9R/xyB7dvnpN0hR9aWg5L9YIdohzM
U6g5wszyquXYKcHbJuBmS3S5/sQ4uHO5ykXd0+tfmF5xJmCZ0BMU+LHgJtX3KGJg
7fSeD3c8ZDY0rapoBtq5IkmAsCDXJvyI10+07FZ/ANVKDzcN4R8oD3zS7ZjUxc13
wB4YdlO0cXB9Gv6FMB8sVTjiACg+Djp+u6l5c3z1g+m5IViQkz53q3jQy0wqeK2Z
kWoXqDLl6L2tYmavx/nsC9IQBMkEHUzW8D+7aTiKyjuhgEBo3afCS7YZI5lEo2wl
LgLn6XfHAoA8Ac4v6uh5N+MkcwQErohH6qga2ltR+Foz91Wo9wA24YOyjgGaPle4
CeX+7JXFd4CyIF3T+FCYeBZEA6gftSWKeigu4irkGcmpqTt3ii4DKg2WsiDoKEtY
/Q0rBi50bj0vEGPeEz0Xv3kw0gWGiIgSD8IVcU6V8poFrKfscDJFJKp0nU9Bdq2J
Q25SP1FDmQstK6P3zGXLz3tXExcpHy1wTuPQjyuJoY6g5ed6qrNzgVmmfz1RiNxO
8pZT/SUTDDo9i3vl6iXP/NHKeAz5nO0cL5Q7qy/eMt54YKfc857aUvlRH89HSmX5
889fCggWP9/+84JtiiZHASy8m6gpJAa9TUnQ7G0ov+ZiGY8KUiCrOauAZQ53gTOl
ahY4A/lbZolIlLLko1cDTkUtRTpoeMZSEF7j2oHpUYSX6PnbGhTTxjkJvyMXAgy5
wYCYo/IJzGvE5zh8cYeVPTTwuJtVWr/ruCarUyBxXQBPsYIFfLl6kb68wjcJ7Lse
sfr3PIJ8dUsVaYWfnvgrgv8ihj6yXVNzNWgDE2JJHdCaW+N99D/QrFh8A4ha0wku
s3PNdwOSrpbUcvbMGmwznQbbRZ5gAwSd9gEcNX9LX1XP7MJfoB7FdcUsw5C2wwaq
55K5o1LD/y+cnFeA9rRFZxAFu6UBrIcr3ZPm6N01cNemvrnmqrmwe+xDpRjQqSWv
6WGDwoKKJf5GxO6lQTjAZ6HAdMXWOIt7ePTrUiooxyi0f5oZEWAIJR0lSmnr2P2i
NsKNOltI4rpO0BObh6thnt1068zldmsWr3FBzspdAaYrbuzyJZ4w1eiCROKP01ho
GXOqbK0AXbqxmIV2bSEU8VWxlsKOiEI2kGX2hWsXAbTjPzn2cQHqA6DSVJal+pyd
pbg+4Oh2pX/R3/aB/TDyTNR6Vq8ISPB3KI4CCKQfuIolsh4KvVEj1FQVaZudOPt8
tVdPKi69QzaCsuIUlDLi+jbepDifN/oQxi3823KprntwDyUtx9oOJ/E4xwPAavQa
mkZnT4TN3onyfhvTpFsNLGgUXXmccRwjzxNPcYr59Km8G+wVBusLrdHDs4RcH7BE
+69k4TeLtRKsHQzgsv+w41gxMR0nnjYCEd+i6K7O2QNzUrz+0+HTS6DaplnECQyx
c89fEjk+yR9mtoNuuYOudtvijkq4ATFN8WPwxdom72z5uXQcgyv1vvEb9FIkjP20
WLh8NPhzqELxeb0wcFDykshPgqqUca3NstcF/Kqpk0TEYZaQhhzcrXGCJSqZQtVr
4nLpRrEyTcDMj7IEomfRlAyN1T5+e9Qv/ipsVGlqgodyzShuWAMvoxzWL6a2przN
s6vHEG1+XGOtNOAFNHppTQaI4myQYtNRHXpWvhES6+pJmIEd3YCLqe9LVrccH98F
y44I+jrdSukluISd/QdT3D2iy9G7XF5BoSSXQYWUnXd2W4reTYg+gp8hyDvye6tM
k2Mx9V3IzoBDEh0urAxb4bF142uTOX8xnBwSYko7s0d40ykEkJAajMfZomZ6jE55
K9FvN09dUJ1SRrDWBfIq94wLAhO6lCHmLCPfAy4JRb7kuoTUjPZfUbOHIZBik4Ea
THaassW9+UB0dkDK3EY/cq//phE8j8mTNOug19tuAm7HCCLEbe0eE2l3HuEmU/r6
xHigJoASVNbzJ3FVmJlh+YPepJQTtG0FkhvC4xvknvlUJrzkerCV/BdX9/lo/t+z
l48kDK2FrUCPhq8WNHsnGcs3KfIcsHQ3FmgT2CVeDN91nGj5VW1xMfnxTfBBHhFt
U+S3/moTZrlQA5ET1/2Q4EoXlE1m1I65uDuyHNl1CdZEpBHSk9Ozbv5zckaz9Iq+
29Sp+FXW7lcoOEQbJ/B4eLk332ZqiOYFhwE8TFvpRdwkCuhK6rRzt5P/QA9FyeRV
bwdVCuwZ+RyHSuWn193HghCgsho38JeWMwHzdZ0FB/Ic9L6JLOn2ZUgucRhYmqK1
WCZez6yXpQn0Y2JYzgFbF62ruIfmmzXdyO5PQKnvWQF6Su5z3LlrE4Pwklqh6xfP
mid+5KFRf7Ct/FK/VoktIHLNj8E1kh6KXSpJz7XqXC1+ql3FNJnV4Z9G/WcJw6TP
aEUiL+ngyMky4sA1TRfCpq5MNvU0yhG4Ud/InEeDjqBQTmS6l5LyGSVx+f4luEh1
V96XlgNrsSdZ8M+BJrZL0T6g6u6rhT3BA7kttZMH61JulQPtXAA7B0KpQJhwDJB9
YFEz5P8C8QWAzYa3A7Zc6W6XmzPm5I6236ESi4zjnQmCPfw53jm4LfeI01Oo3MoH
4HXDZ0FPGpT82T0LhkjeIezC6wDlQT9wxRy/cybvAWwt7REik+5vzPSh9jqhuCVh
egh+C15PrTrDuwzPZfyDg1OCecD5/LRBlt9FohyzxhcSQNoYMs6y4C1i8Sawny5+
cP7h3noqz0naKsyIU5cX1XuPsIEf/JXQTCusbrTnxvmh6L5+QJBArLNYb5O96nUL
k5Lk2bVdSO6eGZhho7v8AzUmp4S80xeUfIW+GGIoH5La3xIu1IrNFhipOsJNBSqz
iVVVkk5cO8hqru4NkmEZ36djOUkaR6dVb4ZHIbhEjjWK3KBQ1B+dWVld2usovrMl
FudJcD5rTizNnXTfT9Dy+fj3+Dwm6Xdn4xXOGW/yRyf0TqmzXcOP3BVsQuWCOnEn
KUMefKpIMH9NjW5QlpA82MsUDVQbJ4LRSx0Pt5wm2ZYNuqPXirfa3UUSV0LQpTtj
S9ybjX8ifT+6J9arqMd4Nu8NY0ioqBA1g4GLcNShNAw9rc6mLQByT6qqC2vRAYZj
bDUxp+L+o2Ekph1UgB5k5tVqNfSSqmguxjgjCSqYPuG1VGAqYN15WyPRzPOZoZFm
gE/spazfNg22sjQOxGfJmN7LixsmpHJLbfo/tkHWQd6RO/lobVkFz5EXFvhTMP+T
7MtxPtK8ksWxYO8y4dg6dXon/6kSANOsG5/dRhuq44hS519BbP8PA9rUgweSaH95
q5HIVMverN9+jzGuVy4GY1eJezJtSM/0gfqat7XfA/vzYG1DxjhJBHmrB49GoC3U
sVVsd6aanglVRsD7P3eIr9HTq8HLtpyt5cIukFXZnPYrOCVw6OULohfSa+Ke1Rye
VtWEEKtUH8uK8R7NUEqnh4/va7o2KLEz05jgjZ9CcrmETxuhBH2tKN7ql4xVwoG+
Na4knoPs9U+DiWJ4YTSfwhJG3EMReJdGXKjiwooCXiuCNNNM28/s3dlrl3+L6iPr
yoZ9y3eMDWCht9Veg57eBl/PFwxP4QgWR2+jgSsHmJMKEr+R63yWNuLtTakUD6fB
gAps2LkWzdBTV/R0WZP+G+agObRJVfD9EGfC6NITPa7v2sbKIQNEi4RWELPHPY/I
jioYhepP5/zua6k8XfL+R8gvBHktiZkUxkKyNLgSfozQfL6Oknr6BpaqsDW/7VDz
emBEpVT/x4v3Zk9I9+FhBT+V2+Cqc7NSvoOG8s0313pSKQlVMcDffKBzbJkBZ18U
ABg12dKFwh+G3RHl2+PkTKhQsSyjCTFgg400ae3tBzW6FD14kXipRSzudqYwdeza
HQGCHtWowJ9Vwk5mPMPvnYd/AJQEp4PT8orHPiZIrAv8mmmh4Wa+FyRkdF6OVmw1
6kJva8grYQy0qNLNrXMnweSqmWFuPvcO7zZ5MIQjNAYL1dikRJdrkCNTMSmkrj6F
1RNQIG+VV1BnYho7y8dBp1ueXxtq9gFku7gxHnCqTkoOTKuzAnphcOJolGVH9lqW
96ksD74bP0zBike9GhyOk8MxG16mLDPwoPOHSCRMy4yD21WgtZzgsyte3U+4LnR7
XDFvAKQJQNcTyTL25JsoKxWiS5YdfGI/IRouBzuQB6UzbvwoIWjg17OtdgUg6y9x
oyi+Cwo2+g7RafaKQieGrFeBNf4Tle6kCYWxrH2EbpbppfflK8wXJDVhodrW/MTn
xhOeax6OV+2Y6QJkIRsW5iqXpHMYbHjhpwdqX+pwUmlvRoVurTJ3yVvH5+viHDz8
ss6EeeqxD26gN1QgvR1K++iJU6y29b6Bjl54Bu4rUHn7cLB3VMXpGfiGtrXCVFSX
wP5+WcDwrbER5/s0mUTt9gxBPkr3tia0wFduxdhVrAdIqjMBaMeerg2Xs/X0De/i
rWEHcmYr0tEonioKMcdK4NxTmdEXdhCYqpzSzghKhK2GKvbNa5vzSwyf80qyRp2O
+lddBHsfP5C1+/i9AubQPlkc0WVaoyRwoPCeZ8ZlpwuX4JSuk3zhU+fS5FhgiOLv
y2NYfzsX5P3s3p2+rypNaVt3UB4aGpeNpoFG6EywROdIDVOxzfJXUXGVjdIEJ6nS
VnTl5NTHpXAbKnZCRaQfUMwBzcarVrcQSowtGl0XwDiATBYd1tBUJyhF9nJhYpog
rvfQFFSZglWNlPcIjEKOjXqMF3JqnHs+LcYrQXHtgf4f7/l4Ch8qNJbgy+LNtnYh
v6nKY0NFfJiBNAVk/cHLHLKVQd9fY0lwBYW6cuh3b27V/ypspN6MAJNRbuOpAcjm
hZ0zWcv7Rk584JmCm0Tsz3AufJ4j/75r8PoyNaqbcSb3r5QZYkyng9IYskQ826XR
Wa6BtPxrblsGl0PMf9gkkVeiQBekptYpFhfL0RMZ0bseZWGNQmW2Scqa8NFbyZu6
gXTX/EK5qXuZoMkVbSk+rSyujbgv3u5flVCyAroMwIwDzxJQcj0uQsjk1CL2dJ5k
o/q9z4em2CQ7dQzLiX0ukiWXAY69ACExizqhLFOcl2ypoj5HbW46wcmAHV/Fu/Vm
AnURt2orh72lbUHiyYhWOviTMINu4OPGaqulKNurnBJXSH5QSaylpilMC+YS3ny/
xHKRkd6F+7IHRPO8mAO1hekrNjjIbHT41wlZI6ezNmuEq6+HYIvF4/GJE5l3sSi8
G6MWb/H6tx8T5zwi5Pf8+3Y+kID4ZqHAphxHbzPG1JWqC6aaQQqH2FVFnepApiJx
b4dyRXASosVYhvIJ+xoBLdUs58KHZJFKJ68O7Olyz2F3ykUqedKJFQN9dmRVXB5X
mADvtuysxlofH58WTMPmOKcIJzjy/Uqv0lRxRkThEHVOOcx0+jTIlpzZ93xZdQ7r
0axcRtJbrwpEoRMM1InTFMG9o94xw1QhIo0F8IbO7yMlkPng8NUgID6uR39/Dc5J
2Ob9NIs84w8mq/RVeUYndiHj58e/CQDq7vQepIAKcr1B7Ys1JTdK8E6onzw6D/q0
ZmMzfwMBzvkuPPniuCmzq1nxmva3jAP+mtEwJMKreut66Twt9YV2O+PodztwxEhQ
5WqxTxqy1cr+An9jdQuUStCDLGNP67ylmmoxN/eIScHWY4/K3daGJJVUFiGt1NLl
e6BXy0pJLgVRBVIKjN3LVpdq+13unWyeI9FxlZxSPfUldY0KRPDCucUYBETxtU+j
0VFrwkOHKgS7y5wUixzEMoArXVmI/04M9WXM0QlTMef70JO2J6bTMoODiJau+hOc
E17NnOIXVr9QjOb6jYPTotBfF15YkC8bmBqziJOM4XNdCGM/72NXBfSLOVvf+wsv
zyO+oZcNQdxYOyzOhANokJC5+JELMwl0KqVjKAAhwMlyw/5TlJtijvex8VRyO+K+
/yGaz94anyeD0EhPGzR2+TXMD6sSTzbSgzA96gYFMFQGoF4pCv4vXqrqUmSZkAPP
4XWVsT0CvlwyhIVXOcB37a9y9tznyF0BsB4/GuATnbg1YlC8eVuzaSW1ds07V76a
pZe6EcojFlMgfv5o6dsr4y7z6j01B2v/w8r98nKjml+KrdASvQa6sZAecapV+7+M
xWaCTSbu6ErG7Z/sEZMnd2+L4oLDrFWYPnl7VEaBHHyuGQ4FJ1lo1WgyoSwqpACv
gPTx09STWPikuyAdb6NZ8LcTPDT4WkTtQhzaNgpG/lTjEFiuqEp5pZs+AhmBdOc2
YTXqzhzb39d+nYzJeXaXGjjT0+qNOHwJlZlbNA1luBTtftxiYTGTAWAq1LOzFKkO
TXUNef4DLRwoP6m7BY1yUPPgQvuEZ0aBJyleWu43jbZi1VPLG8e5cKocY0Jubh6j
j6ER9/eGhqagfC05j+bcNaRQR4wdGjWGFR7DgDvhDEDJ0Ii4pFmSpINThIACJ1hs
jSbxGhmLzgdGRxTnTlzxQDVNUossYLqnYMrRCuL9JDVs/3tAZm80j0wvrBBYbxdU
7brV1SUkgvKFaD8lhq4Tm3xSSWxNcXNq8iMYfbHBGqJMdr6n2eE5DRDJ0DNoy66u
4Bj0dFNsmZF/6grZbg/vagjjqW+7kyMMH35pxTEbYxvgX2zABOgShwzjTMIvIiZN
yPekeDqDiYD4UMnEfbr5gBBW5hg9Z7lykLGYyTSyp8A3Fvss6wDnSGW9gNVhqX1n
ua91d41H0yvqG3FG89Esbadngu5MfCbBUN8c7s6K5XaYKV9UGtebdcNcUn4ugiex
yXi/ZMMgC89Q8W7n58WEMg3NsfwmbtqvskbNZKlVL6dj3tzjWJ1q/LgTQRuKmr97
sx2fcZXq1WY62p6qjF81rsk1qUILaQrNgB/AoaRUDggjGjhDOLs+f3gZ1TPInyV0
2EDu53XArt1qCZniA16I3WI5aRbmUi/5XLZWhKAaoSmd5KGL5ODAu3dCo04F1VwK
Kfx2MtNLZYqz5E472QazqUP9TJxLwyl9OIxakUNmDCIO/0WSOt7OCJN9jjEMEuI3
uilByw6MFq+NClvm6OzrBDkugU7HWW9MTjaAGB79rT6HawBH3x9af0cwqOcaSUOn
ygc6k3cEA/lw4rmZiOmkjpzCXckm0S0TDQHFPKpog0lXZzI/bTNlWOw4n7SafIZW
a0DWfyPO0TX7wCBBAtI5OrdEoOuFPiBtgvIwAqCsjDHC/MjLeKzGn2AXFh4cwlwP
wpUORTijo/sFYheQ0Y8AABdrtqiP4+v+lbRIkv9sFmc7b2JVBVz8yu80UK6f1J59
CFktLnjiggMr8QXwLkoDp1W/qXTNaJvcPfK+xzwo5etewRdwTVcIuDeSMQPskf2S
zLzYzdqcgUZrPcQgcG2kqjT1EBx6ZGbKJhFWdyhXOfw3hX4EDsQcLIeLP6QdYqZB
JyLXVUuU8+e6WDFWGtKwQJdQPdx7ceOapqHdnOvTJsZhFi4JmY4gJ+6KQnSo5z3h
c6gvdXwng6lV90YXEt3f2W5WeO4daWUyu/g33xhDCdkIo7L8U9p0ysje+8nR0CNu
02AXxglrRqAafOtuqLJqeY+QgDPXIhNJu25DZ0/XhcyDgOTDIUoXiG98DItRuQ+8
K0h2ApIqigepJGtBCBPPkWbhgKpTQbzci3Zm6cZaGfLd8VwCUInf4PpBsFlZMYPn
NWAGstbqUNQ4B2p6EywkNyVKL/2wo+K1VPc5/L54PBOhjt3MktU3wsT1aAYwUQii
FvZkiW2QTJzA9VtYRCh4mCiapM5sqETpxGQlmi7y9uLpeo5/wePhEOVsK0nCNfFM
BwAgXRM47cw3a2mjbCanAFKTod9tFiRbXE4NeTSeLgCZRcBVTu7bnpgQoa8OXGWf
TFDUxktKhQdqWugq99dkv+5xJ1aEyxfD62rOW6JheI85MuqbD2IzXmYvQHsiq8Z/
T9dtDpqoM9HpGa1RngGa0g002dRZigDay1fHIQLcIxZZD7cRc7cdXDYlqD8I+K7T
NoTB/2fpqrQXRkcDNd8UiVRfKUAf3sPzNMNKv71ujt0JJu9Y5sSYbRlne+X/sAMk
58u3w22hE6nk11zjKnIB3vyzCsUcrYkRKtUbIGk716LYqSi3cnU5BBh7bJpgRDcK
amjTpUKdT5nzAvp8aY825ZoipTXvofQfhmB1gB8XZIBedsvIpEFS7kp5RUeKFHjx
cT1TXeB2l7/7IghqUn4PUWx0WcRvK7tAMh/qq7kYoJJrljAYYDL8fCd9pLKULhnQ
ZQm1RnXYr6WU5VO8eet7lQ5PtnD2iOKvZlMKpTpfskmvALX+Vf2eTkgQSx5M5h+P
6iuWafr1z2rD4h/LCDmha5+wSZtZAS/SZrc1xf+10TxdcGegByLQMu/iTNvHbhQf
6JIjYCJ4RvKb6AHHRDGiwQVmdRKRlQgYl5OKNCnb4oUJzPeDFuXj0vn+1YyCVkDr
l3Df9J06AfST7l91oNlAfkvrs60kpSvIIGpMAO4fpn15a5TyhAMt1twPtstQ5j1d
5IJBf4C7E0Y0X7GVYh3zhuz1tS76iDk2NBSJ733yn63W0Qq934jrOz/GkaZMrjwE
xASnKAJxwZRzaMyqve8/83xVlC44IXJ20EhaRzY46Tlu802sjuCEYpVSraXlgvqm
3fjnKdGy4jxpYqclXitqYrzum4exd9zwfnyH0xD6++MrDh6sgwR9CKtuXgx+xTvh
z+uTc400P6+AjL0DhAOYnIAI5Yl6zjLnDsDxzgh4Z0BQSumf+x8zvCK+0bljGH4y
IXZ/DvmR8Ei+cEfYK+Y9G0acjCHAIhojo2nXaaipVwx/bWSz1Dd4v8DFemLib0wf
6CR7nM0igeb9POUcSubrzk90uUUt/JRFib5Be5nqwLg8Z21/9DPYWey1RyDJGfr4
vXB6elF+0U8GjsSKvjXC4HG9zdtXyVOOoTvBxnFFtkzwQNWr5d9Ac1VGRijbnsCh
eFSHoIr13yExMZ+ZRkw3TQU7QPcL0VQKpag5ZidsxEBEcmsnjW+srf/H7zKj4yr/
33hjZL+MsHFLLGF3zSIGVpiMBG812lUwreyEch797mXuHO5qTtNVk7nQ61eJS12g
iS74NwFrA6xeXkFL6i6epvKpr0rVnnqMcRF6iJogzHaJTTRgYXdS3HSHrpXJvRgD
PQlczyOc5C4/IAbWHF9L4/COVvZXORIj2x/b/HEA2bxSQxx/ScAXYuGfwrtlEzhF
2hLL76Y3FZkRFXiEupgnBpX7EW5H8aZ2OCf5cIJR+AQFWr+WimCDd9SYk0Sev4vA
OuPkhc0khfho8mBWHMkMhPVvd43csMhMc9tNYdtYpIRilsk5vxqbgaC4qDh7pv/B
wbe/R7JL92IYVlKArmJ0pG/6/DbIlNsIlBa177OCtoB4lnn9dP5swe52EjuGJwoR
pfr0mD3iBit49PUeGZMew69KUclBy9lHnzsnnutWxLzRjzb0IOjdVRRZ4Z0ds99C
2azdAmsifMXA3n9i0jVG1VdjjRe4DKDDmLrGV17tlRXpFcMCudLndtqYPu5Eth6E
b8utpXkZJOyjBrwpnbp+0xeWCsGxflQM8Sr0d2zQqVjLRJDIonn0PlR020rtwMiv
91wL9ZYBIl7QHb1Pk9wOOcwy7rRcTWyYPqOT10nPrpQYFKCWH7BOvlYsTzdXXjO9
jMTNg1/jbTUuqdfXUx9UE/wJ9DvJe8lFg5ncps05tXW3DUyYkW3E9rAcc8q0Rwv1
4behvbWCGOQXwMg7UNAhfIfq5gVRFn17pvdSQ/wL9yp5sLycgGz24c4WHpdeSZwY
zuqaRc5KPEeMhOffEFb+t8FDN6QJk8SMEoRCVXkW9+PjSCUmz+QgI1lvXwRgwRPQ
vKKGAHPsRQzHZhFGjkBoZzPv8P3VeMm5P7Frdnnb6KEH7mAsxR5+5n6pKBZ1eckr
rpgL3WKdpXD+zbQCMVmQ2IGs+bw7pGo7c/9YrlgIFZG0e3TmcOp8I84GWQ7CXXPL
+A44ps1rpR2eeCqjC7RaghXoqagBS93ywu13VdxISwQAZZPlnPkLwKbL/nmbofJM
qM+lo0q1Qy/XxiaYxHAXJ69aHP3eJH9ypuNnxkzpnDP2AR61c5DNAwXzVp9Srxpq
3FRrcIY3vTTEUYEDFuLIbBzUrZKuT2LQD1xDYhT7qf/5tBKG5mpZjnZye0helyPv
9hp9SEBiB6NzOjd4UTvxGtAQ7Dbx8K+6NSnC5aZbxO3+GAvQm1+u0tEYSHtjP08/
Hl4Xo8EmyMvZKsaaHaaxrhsDnlBFkY+GDR6VlxSPe4T3Nufvb/KxrXxGkfmiEQXp
fzTTn+7G18aw+/CESg7CjKI1ScjJ2WH6d89dT+ufLdE12JSC0uCey6QAFkzcwqvH
IkqmDmAmDQ9L2FihohSrrbyUy+sDlGmBI/HrLNE3AKdcE6dUhpmw8QLNvdDcEUBv
EeHA1tMXvKR6g5tx3nRhuEmZdEyHbX8HwWIcD6GgoM3WKo40QZlpjdJwWwHAmcQJ
rp9f4oW0DoTFZwYyy1v3LZJ+Vo7FYeXCz5ymYLe3YKPUVn1opf4TaiNoY70IAaYF
ehLCgPEBHUlpt2G2UycdbYPIQx/czbz0BJHjuhlPyTZlNeOh2bRyBkiJ+POEY0QQ
OJSj1iakQzrxZUby53LRbmpp6hBVwucXto+DT6/qF+D3wN0CB2Rd4qlcMVzXyeV7
DY0b+YhdpQ3FtGLaiKULZPL/ym5XVXXsdSYW0TesuuF2Il1m+BXsGASDy324g9uh
LYpntf+vXTgw8eRlq9VlYPYPvbHC4wBJEFZr4w8Hwd66NsCJGnAWbal4WMxpddUK
gBZWRXXBL7HjHSRBNzWNPEfNsvKCjCMNDBEK2KKWWGkPaOddEKy3u9UaCaUfm1kQ
M19zfhKFdBTTmLE8qFMrwQkAp6m8pHnp9pGYM3foP49PgrqEmJdgISa2ITlEyZMO
UBKdcWqiOhQmrtwpVmuj1pzTLMb2iK5iwWkhvw+CvOf14M5mLy5zXLtJtOEhB1UT
6qA2at6YXCXFxZRgNG2Foe5jxOFS7MLtWwwHqfs8wU+bz4birBc4gL4Z16FpAyZZ
Huhbeo4vp4Y4j8b6QvcJfcr5Nr9t3iJ9utHv7Vtwl6uoqDxKTjCZs9bMvi41+Q1t
dUq1IDqIR+FgJEV0nZAxuzjOckr0JkaUFNeiB7WDoaAvk4cnniXpu+D//JQZ/o4g
luwHQ/kGs3TMZoX55ZP/JwZckDo25AIhTWELXOsfPS6V45DqYZXgKmFd/sjy4xP2
zv6VT8mxHJBK/QycMqO9iSLqRMw0dTSHiwAHHpjKFvUXt+B0gZ3G96gedCl+AT79
BJb9woPtm0LfQgUHU7z6NvwjUkzB9hg7ohoKA1Ta7eEkCf6LSzI9ZGMtxUPYwjJy
HWhe3QHoOqV8DxbswuWvV3tpJTYDTqcmHfqXZRnkl/uSiZNTc5k/Vq0VsQrZrQKO
/4RvA3NVah6yZ2CcUBc8FB60awoSeIXhRzpCE2DdqC8OxV6ZqK1QF7Wjkd0rpQre
B+Ao/5P0nFCrjMoZXUCtvIkXFRoILyNw2tZrBNRwtz5A0pXUnLJNS7xjrWTA1kS/
h5myQLbDXeOszGTZhisZCoh560OV7BLhoug8+ohg+HMGqZ3Rnh/wy7DjB0rhSpCh
SO8XBQZOFqWSALksoeKoQqHF9KUiNYiunSJU1WbJASp8IoFjOchI3MWnE/aAmtTK
Tje59Tba1RtJuucjRNqVM9TWxv5tgTB5g3l8o8iArld38OIqRc3R+/K6Y95I0zOq
jQrPY2tuj8ePRph/YHTATDyNB19dXkKnX4bwxsiBqTf33Jf1CPY4Gl3XFKlFjAdp
1/nMyJGJl2V7kpp3d54tXjFDUpJJO7DGzsHw0zl4Qux9uszShfLxoKdPNzqxVUgI
EhD5NPJLQnzLXn7XuJls7O8M0IamW0dGIkE+BMwPQJb//c95fUlxSx0862GbhtvW
NbJY68BdLJLfIF+LZa6zXq6JGTxgJbjmdeFuyiCAjEWysOnNvoomu+oT3uoXVtRV
XQp6Hlfs6tpigLDcw7+vPKFW9ZPudolL7aV+7bnAkzBdg8L2UNHsEXVcjkNNTLjq
ZFLmxzetO6YQZGhnJEmNkVtbWyMBa3w6y26Mphxftuuig4xc9lxiegGjRxvxFOxr
mMMtl0WRjP+hl18RfvpyzL0Bi4AktAhj4M3KBhCB3DFS3NIS81pnvX0sxEYko3b+
bOzaOkR8A1v9OVdI+SwgnAtqeMM4CSf1wHRMjnjNvxuIqGysDGNznXGhwZArmk22
lMc0hf1FVkhiS+8W1BeQ4fWbgX809KkkFuXg39hKPagLjyQTf2ftWVcZi+UdllaW
dX31KCQsR9aH7Y0epY2YpDuAr3yxuS84t3Sxc1gtkJojLxXkwv64LGf5nppoihDP
xnfl0oIJrtPNo4ocK7PbX104689hdKAE4RUzuAJyGHmneQ3A8uN26XUyckbQX1vC
g/hhZ8Pqsas8s968ylQyxaSf7rl3Sn7X9zotEzgCT3DoXcizupjq+rYnyqwUWF/I
JCW2/DztiWZd1bbiGxX+JhiTRxQY/Ajq5qttfBNrs3BvN7ZaXtQ+y/XyOJliWxA6
8j3gA4BHplyTBkhJ84pBsyykuUa6K7k8XO1hoF05XCrTkW1gEZWP88dRDKpP2H4P
dJh5NwNhILLSLw4ekOlpMx2eVBcvWVNENjkg6SIIWcpq4CzuKdCQPVOZW56vP8rg
MHO0FP+DcHsAK/g0xQGkeUXS/9SmVvGrfDmfdwcXCOIbS6bZlYudQ7hse3zH14gW
8b+KGYLCd69gz5qRR1FmIBveYMcIGsGh7xaGZzHuBzxDYGs+5E6hetI/Eb9oWUFX
mNh/VeAYbdc6mvhb6THWAmISU1UksfiqWmOUkMOXFMIZ0vPh88sHTtaXBlZQLk11
krtleGLQ1m6BmGAKcyxG3Yo50O6lgXexpeRnEaxbFwPs6tf5AsdJ9ItRgHGqW4kR
oqbCGVLJmpWg9u1k6VE5TevkYWwSmgHA3nwtOHsXbr0NzyN8RrDudCkI1PIo2q9/
TPyBsDGX03AipUbme5Gq/bOKKU1U5UxypwF2G0RuCVLCHM1P4V03KwjWWFHg8e0w
FXbbMTYdvk/RcZDD3w0OjY5It+Oy0huUdvBJDJ29fGGZT1biyX1lsTetXZSDtecf
boaFdzh8lkLNqjkEc/ShW6+dT+TSH5/bsJ98cFZhaRc9NQt6JWmzRHFGeeiDCBnO
e6D6ec9y9KRsNhrfpTlTP4Zvvtnb1JRLVz2eo3IAilNnit8vgryoMiZBGgZinmhw
WkgFVr5XA9/GlsxzgqyyD2ccjzgv1XaCN83JQ3YkqbY/ZRWQJ6miYWa8/a7zkdz9
SZ6vRortwBR652usrvhxnduk5HYUn9+vdubXyNOf4oINRplOQRwe5rnmV6+Rh3UM
IcRGGgFkwi40/SkV9+0lC+wrCrBx7C5Y+8HoJ+sj2qlSTEkdRCI3JjG/GTRqbu3Z
OPLvRQETDP82J1jylcRgsD8gqXQffVpSfvmKE7Ogs9+SDlEPLQvmrqLl+mNoYwvG
mn56XAbvCLtlt0d/g/ODHWOcHFCYuUYsR2uv0CW0Sv0C6efK/SqIMhyymMTvgE0d
v2lqcQRMYcgUL0Vv34TBLX8CVStjt6RzXY2fheXMzrkURjNK0YzZl3vd6WL9yh1+
Th35aCbgfk2PURyaN1cQQupelWSToMkOEgoO/ktibne7dxT2dTch36lxlXj+qCqv
CpgaBw7ijBHKnaeYKszAPei+RluNpdcDECPTcrFx010Plel85RdvhBkUUnn6ri40
GRfIjYxeAkvRrevbNFtFTYEIhWUBxplnL8jM4G6pap8wTnZbLUcLyN7F+OxO0A8v
YF5ixKiAgLCyfCv7y8wO/s7lniBjFmjfNqna6yBGMzuyOnSM6qRv/VMPRoZaJrAX
znelGwjTl6izLGPU33MtQULhJg92TKKz9PMqDQnlJsvIjcScw5r502LXJ3wq9WQc
M86P/HZkXTY7EB+8CIPKfT1bwLrQqp2tsLaHqqf8aLIYgJ1SByEXLb1HOp4KYsIi
j8IziEW9/17HIIu/yBAITIBmIeofLqWz8nptSKo6UGpx9BJHBi+hPaXtpdvf+5kX
IUqxOAlZdm3YskTCN9GsgIhjbE//T6E7ZIjmwMbohqOd8SM2t9d5l0GD6en6b4oi
d6Gp0/yNxiLderf9uq2BVFTwsMgF3NNB9CKY4ELpttCQxsHrKYoPf6My//0DUode
ls2bzfNb7Y1RODYDO6aDRJE9JsyCCe8+ppwUadi+XtIL6yShRwXj0AZewGaCdpgU
HiOCJsTR+Gu/4rFDR344UEZQKV5qPKwEnOFzjDk0phpX4EMT2RydOw/Eqco8N6N8
c2tskUyYl5k4zKdgiZflzoYxYxwXHoLP++FOCI6h4XQmx6TKnOqNjrihwq0jaDUY
3/79oQ2Iux5RW72oXug9Fsbt+wPmEgjsTADrm2VMa/no8m1TLOQnMCsxJ3l42d6V
98qyUH4KELBLPP5HRA+FTNW6d/S5uEA8O5C5bOKS5MnRTs9IRhT3rvjPmMjr9Tw0
zb9WeGwZb5lpWfUPOrzNDqlSVNyvIVl90Qx1B5tSIj/agNfG4bG1dEXsjJS9p2bw
tow8QiUCVabTUY0NpWeVSxTDz/3UjjUimd3tGWIfLmmiBRzMQTsOkvDjRQf95frB
8K+4f2+uuMt9fg2jo9voLLZhxiAh/QBGk+z8rBeXz+mEO5r73cD3F1LOqDYHlESd
212Pu47tCoDCcs6fbVQMSLOw+PndRi2Ma4gJ3/9N//hVHyJng++rLMEZAcqZRAsn
FIny9SZtfefiemhqXc0Aa1jKRv8RzJoZNCIdJLXmduGkvCgwjfRd7fQFKursLLv7
nPLA3lg3Ylp6dibPN3MJ4VC4H95fe0HYgEmQP0YqVY5XFSm9PFGycVWxisu6J6i0
70TFAUKVIorLtgsPXU2GG5jLLsPwqFoj8gIa4j1JmERvhPNrv5PCKfHGtjJqk7A2
QUTS+lleDyjoZPvs5JgxinNpQ1vyOOh5YkucZsCnZ29vQxVAXM802xyxKhnOCHaa
CN6tOWMxLKqf/YjbZ9xK2IAOSK1idaUDTnUWNoZFpoD1EVgb5s0senyqqSxVlsE2
3ptQE83hORnyeyw/nnPl+hfDL4mYfzdouY1AwkeUGU0xmEl2GIL6OSkaVYWMfU6i
ACMoMPSmW+1x0dYtwXMYemQZUdxqrbUOuLgICUDeOU3KHMtPowUtVZT3hzxQnJt8
CNFbbFVclFZEb6S3pvp/lHx+QwQJskNCpxgKrQIj0GhheBle1U9xR3EAysmUtKJT
yBW085Vi+GrUEblIo9qkWd3UePz5DFI98hDohZ7s/0/vZw1EpWqeT7StXuIfqGj6
0+LHVCPgd2DSkz1DYYzI7OQQk/D7ikLjfYWamth8yRKcSlwEPrGF/8fcaIvBz8sf
ouYYznxBjBweS2CHOhSELCqVIero83BlTcLgh+NdsV5SiaBKuPQdeVy+DPOHkB5e
v3mnLngIC71guUh7J0ci8kLea6HTi7JzjioZsVIMeG8a+R8GVt126hlm5/GAeaLs
UoaSoQHCVvdB/G5dudFGmlarGRtMuupbNKT2jmdt+ntU5PFqEgAwK8bTJO67CF+i
4ZUZ492LEAIwNoQ+8aqfdKDIAeitaEFsGoixShXuSAZuN5TReF+V0vIZYHQP70Ad
9M5MUgtZWTwkeF8v+tHUw3YwAEW6VMdTJ7v87kILR7Y3Yq7nvxG9912j1NXfIWkz
9jL8Rc7tPocuuII7HBgEMGww4KFx78LeKn3zqmwbJi8xuExS4TG03704soEm5lai
NigmiXlSSv+zy9Axq4YT/VRt3Ul2IGHxPCuJ9993nMNfITYJ7ic0jb12fffmwJk6
3NR+/sXdYIX38/ENbpfMS/2xNgzrgeIymTlfmMhzxEZxBzIkszJuc/Lynaj5Kj9q
AK7dNaZnNC2YJ+N5F6Z8J/DvPFofEKf4gjUAMDCFuiqSKXb0SEe7KlHggSP2CLXU
SGARz2DMMnsFJXXslVhK9LfeRN2c5eC0kX0iKAPcmIcitPEv7riLwow1BGZ5rzL3
iu/iMldkREY3wpjDYJxiqlMoMaXB1CGfKtZwWvOjU6phznWUY5QlUeD51s5d+j6L
1QTHQQ4SAcwvyVbAqwk2ltLdrPe29ZC8oCBOM9rolOlFDhcMjuZ8Wxjsz+g9iLza
6bWn5yQC/ebOYjrzxsmZzUEVcGTip8LtMM2SWzTPHpmrBUST1j87Ahs2beAZ7rvM
ss8JQ7oBKfBM7j35rxKp1+689F8xp9HliA5binOvCoZ2IrhERnriiogptP3Rrxoh
CNOfzpvyF1XzEr1S2XFsEKTuBp8f/3GJefDuq2CYU+Yx7G8GnBxikjXBsbexying
awEId5VXUPMvlPN2M8zC5/R+YQJ4zzuHPMKEYarHpJEPfhIry+TKHrGdjc23eC7e
0MQGsTWICKjP+7UsWM95w7b847L6nQO1uQVb3hf0VqvK0XR9bt1BAGTxB2jY+Dc1
Le37dvb7ysQ9fhHIo/6/56Cu/NQpw+Is5cxLBNWKmmQ8sUvSMf4OElOPt2igYa0C
F8OahhnxCl4vF2gFcedavEntM1KQZctZ+E5utrJQrZfWdfqOuMeVhAWQrT+bPH3n
cyJs73P7wcXHELOUrxETkDO1T9UTgsBNRKLsHrC06muHru7r1nCZISUUtkZaFC/P
cAseD/iAozmrkbNj2vKs0Ez//6fhKWSRQBn40ELNs2DNlAoaPxay8wHljKTgO3Ot
8V7rFmg336MA9YzVU9i1mWWol6V4T1pYwvrQhIlgtpV0DO6kT6YGzVC6CSGVQ6v0
ocEZmbjPuU+jKisrQ0G2V7516eaXGcxLY3F6FD3izzzZlGJgthOJzcvrEhmNj+0T
4goN6hy2XpjgB0P2aNG27QEShq/oS1sae9aMFTg349P0yVVgB3iZzyltU26e6wEM
UTQ5SYk22VLG3sICl2+b06UgdoW+e9AZRRaoon095jhHovIQd2et4gBCB+wmWFjW
HUUq4lEDqivg+/OVJYTUFivnNEgZXnFGfG1jLM9Uz5Bh5NHR+13BLFEVoRFvs8Mw
tHBBXJfRaV+Yz8DXH+Rt9ECzIsVGTUajGnO3YreX5k98e2BRMw4tYQ1qWJNwWMyy
s6bfGIB7JkciZ0ot6o0lgJB1itUjDzWtLLVBM4sJQI8poOS+eaAg9aYZZO4MxdK+
/3x7k8MQOAyu2E2URfBfdvSGxBnzcwk5TVL69uC38xm15EFe45rfVPC+oIE+Au+9
fVx8QgpBZxMszWUT3yI8dgWDlHiYUL1ME6n8voCN07SFMGzT3N+YO/aOGfHjOnQi
Zqhk4SrYILyBjVLPahIoxtT6vAK4eXnoVPjh+AC0kFf6L17Z1sa3ew940Mgsmgyk
NQ0G4tUjHXs8i8JRkH1TcXRxosSl6MjovHeJQ0MhWHTJgh+pMeB4z4bcTpoJPz6y
pviVyCKCyBZ2w9IXA1nPv9MybuNaHOZbHWOw8EZNobIkdgVpPSWZDuQ9ES5ZibMp
KppImkj9zY62Ip4urBMwjHUQfJnkJ3igJpsrQArO+P8t8spRrlqWvLPRiNdrG5Fn
x+YkFjzryapyreBlkyUekKWo3aMVPHV5vzrTiZ50vsvOHD6UQ9uKLmyX/K+F8Gm6
qyBzNj7L238dpnQN+65aFqbuitYO7VIT7WyR7MYIBzEw5PKC/ZdQ7+OKmZFrfVXb
AvBdSJvjLLsuYEnNFoFSB3zWSEav/o5C9LYVTOY4Fp19DYlR2QjlEKTPkRTGlO7/
ReO3LLTyR7Ezld1vTvOx16AfaKbfRgJAAX9f8DeNMXwZfR+Kpwkk03wSFHskBpdX
FZRzKf+gf3Chx87ynMMMHZovii9x+mn4CLjMRjJ/XP3Q15X9MWShbEFTP9nRLGgi
jWbNVEJdX3q0Z3PMLibyqsoZyjmZbD6Cmb0vML16GvL11/WuNVdTaWkNfMXxfLHC
KSF0iY3ttH/pZS4h/+ptuEwBRU4KWavQ19NkqsIxeKlPO2cu1lxGQsLxAyj3hoVJ
k4ECcTTyK2Sl+uEJjaH5QlT3lw1DLOAg/yhW734hjBlNc1K+xby1EJQOuFj3SXUC
jZLrzP0Xh/cUCYQ4QaYoKAVQr9DPhMXo9jlsLeNyYm9om0acbfHx5GDmx9vS0WyX
ADwcsBEzAZvDkKYY6Wsm49J+9eudfamMRdMWlNJpraUX4dn1sRHIaqqAupr5Gbzc
AwEDjWu7tp/dNvmDvjQvjqRNstWSu8VaO67oBw2OQkX1jf0eePPfllnmch7QVsIO
EsxoZp7RF4otGDidcblzKDBknTxiXEvhKuNmeEhnug/0ff4ppvwuVjWkLLVsLbTC
gvzB6wnAdiywzDZkfuuvJIEu/M2JphvkSKWF8/TY/88SKG5tFvPR+ElLFzmI6Qg4
tp+Ms0IY4Yp6eT3y33KDEcbE3CKRRHm4yj5JdiFBRwuIWLiEukzJicSviCDGq2LD
9+Ok2NOESEDyMkwMD3J9RaOezwnDnp5KV/Zvs3SbpYJX6iIMpXOvs9GvKj0CQLXY
BQ8PepAoCFSIvu7RIkHzKExy7itYizQR1oJQABsQTVRuallfxDh2Wqok/hc9sORX
i1QTjSFOL5NH334iqcs8eeykcP4bddoU9HdQTm5rOiYwawyhzOOKg8gEveWAgkxC
kGqjTBhdMpNcccfpupzrKyGgTYGnGnImEnizcDE5wt2I1fwqPSGmILCBzP+N9PL5
rpNvWznPaT7VWTWbfwkKEqdd96F/Mc3OqmA+STwVFYmFlLHAq/KPy75UOvg8qm2H
GuheLHD2Nq/gDrCjam01FA0T/IxA16IJy6UdMN/hqq2XHPCTw0+CxcunpvpZRhPV
OYTylSlgtLtKt9+5GRVVjtZKokkq2cILlX/5zgSTNIAoTllYZc/Agc+5nw9oupU5
Kmnwl9NCy0QKYWkMiVTTfTTA4uot7qNSsWxTLb9wWmfoxUsSMhNtGNQFpcMsbA/2
B7w2XF8gzyBf0CFrf2uwy17u16lLyOwHSDlg5zcMblSIg5wdDTAtPDPX5w9p20B+
r0JsrRdDG7n9p7GINJBNCDCzQaJz042cuAxiuG2RMfvwoYnYCJPMPhh7mW2Up+o9
004JUFP1/k8vCtBeDJs3rPe1lP6RDD/K9fyYoq6SSdbhj2UbcZiWqUZEFGCYWAGB
qal87rk+AX4yMEIgncSfqAyttaqVKxWiiK6wphHi9BXNKqOM/yFX8+KWNI1o1y/s
Td7Df/iYwaY8G7QX6OXcF26HW/z23ECC0+GvahLdnH7X8F4YWcJ6PGM+800ZRgdR
pRK80G035SRAfj3aqeIj/QRnomac6xsR1zK/8NQXLZfxMwaQQtDVeWZEFGLV/FBM
vFs+R+NMXrbrLK3/LndySsPT9EnLWAZMPpPLJPHCXHlQGTLDAlDjnpCmWUJuDYWF
SL4MeLqrUxZNxbDP1uDs47nSsDmP2qNxpG4Upcotd9HtuXhbtyiiyLEpik1lAPsO
ZQcS0bNP9KNeAmNVeJOcJxBh2UJ5w3NamAR4eYVs/g4yAxgR0yeOXquJNYLGW4yY
XeWSorpqSfYF59YbjKF3t5HKpvG2x9Mk3q8kiUeXMRuEY4GhMg4CE2gMcqRyVfE6
itoQrRRpwX1xXJP542bECeSOR5VvsjM9exL0dlYLzpnN8llvwgci8QYluyJlXfa6
zcjuZkS8dCEmALcT8oc6nvUovW9CkZafOV6ggjWme3T4a0feVYk9O8fX5CuudBek
TH2rbMdWJ2QL52EqvjGLY0s4TyOjw5ahW29hMktqQzY/wUcQ0POqHUa8947WI7WI
d88wVQGdQFs+TTrsKzXhNFaaNJ2kljkOC2gIUjjNr7SnT/MrSSaR2A57ykAS4OCq
V4zGR5TstH7v2+s/Kbaj/G9hoPP/b/eVItnciWk5REJv/zIXufqhsOmWGAIseKhH
CuC2PYcsBgBip7Cqr4Kr7UojxqdUQeH5QvuBBx7uojjWGgwVkXz4NxMXhW+u/v8o
zqEYgh4Z9AUR5RUK1ASrIeXcEEjJoG1nupaZnSdqUxPaz1cslBAsMuqA0A3/wLvU
L0SBcnAy7N8TY06FJJC83Dzb8jt6kQh6jBejC2pghAuhNUVvaWmp6HmfFlFJYBMp
mbqMlCrwMR4JGHWVaN1Hdzo0TpBoVWbO6nFs1xHHUQ/rrws1U3U7ocFq57JVzy+K
Ocif0vF/X7jF2QRhCQlxQHpJPs+ga8IJq7LxC31DKuer7XAQhho9hO8PHxCRxQpC
61h3kEWjPdw3y53Tzo3ZnYWV3ngH/aAOKJezuCBLGmIZvwSGlPrqryFEfeIbDJRs
b1Xp/FyWW0ZTcH8AJSMjAFkhW1+rZ+rr1DKkNBzUN82M4lETlxDVLI+M83vATCJv
6rXsljxOrhcmZrrcMpEZJPKbMREgT+cNqK0kcFSI9lnMr6ayiGNJf7qEBNSCyBfM
HJ/qTX/m+MnwXH9zUSuj78OdrRmtjUQsprkJ26bE7KEN0yH+/dnzEgfaXqr5+kes
N3/0Aj80mWYE7k6Af5LYKNovwOC0oLsayc51SUUyEQ1YVfZ4IO4ntAo2zTPuC3k5
cM2aSdubI1XEPe/xZv81hb5zprP2xut0Ji22XB5Use3NeMVpI20Fp/PQvey/RjBl
H77KhPvtzx/5gXxkpInzkQuYeeZGZ+W55VhHAumBFyFQJJGAMQQY4xgunaP7Mx95
T1HjxxIdg2YmrtMXbI+/KJR/53IOlvstMwgKoIVwIsojsasDxNoUcrDmZum1sfbz
36atwGmWR7qZBaVQq9TJsx6j4AMAj6RnyXWBt+H8gWBs0Mrrx1inYFqKDImmKi+u
oW4sVdP7zGE981MpkPPEMKfsraMmP5XX81A2xnJfDBTul9E76pTC7fzvwReqOAds
DOs1t6Xtbg2fJnOeMYqQRQcf0i0c/c+vJqjyEyujKebqUZWmbPRo4BnQBLQ4mWId
l5fwEYoiBb78pFBuoGdiN+d3yovIAq82AYSQp2//IPXzhi5sDcOpL15JsRPy/DP9
NlquImjiiQ1UExel3ShOr+jChc3xmld74kEmtnUCZESjGfo3K0pNxLGeajzd+sbW
VBnnVJ7RFozxnd/XXn3X+lWx8j+IfVsn6PK/AzciNJMufxcJZnIzFp67GPRQK4BU
4U045ksADoQjPBwIzsvUgHtHc7qIZqZU5V8k/O0vPe02XiJs7cGYg6L0f6bLB8n3
BF88DwCQyN55aiQOC7gDpq8LQqrZm/eooYGgXhOpnu4uB4DB4PKEsQosk05tRtOb
z20T59YAIKToyHpOMq7v96xTu4z6qkMObHpPaV+ijL5mpuifpWxOsuYbQaWp2Rsu
ucjJZzl6BZGY0d8SST7abIwhw2vvx4bKw36T9edyNNFQdMwfmSlvCwGkWYPLuVmv
ZWiF0G3A53dYG4BfwofGaPBtw6qhLGS4MyYhNUZrGTC94rfqpub5pBgNEeZAAjHA
puBRmPQsv8myv1jjPd/yY+gH+IDtHO9Cnd80ezOoqYJ3032u2kjDLFGjWy+vHiY5
lWcxDaHIVdv0x6fX4aU/xce8r6ROYSpctmBkboft5N4HXWN7W4LJmFFE43EI+/no
IExtl+V8FG3D4pNr9SJPmJG/Rd821kCfVnD7vY26V+Zv2AK6E/eJKCvB6XxvZ187
O4K2UCR50SAXdVVf9/1BPRbJSE7iCeLf41h/qob8+GPVWlUDyguEmOx2jZ21E9VQ
jS21Bzi15GHeyULbV99VkQjGejJEOPugR+ieRYJ4ISxhl/pshRSalE7EaYRwUv+7
U3pZSoZuWF2ct43oCv4Nz/h8x1uHafPAjRXOgiiXNEaiNhiAf24kOGq0ZUN4pfXX

`pragma protect end_protected
