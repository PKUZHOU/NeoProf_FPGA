// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
MdWq0payBn0Rmhad8kPEa7ndbD9RS4k4Zzq/u/qHyuLpzLH9rrnbjdRgvJwr
nl9fifuKy7yaF4cHlsILlaZwBsNnHWAvU85GgIz8dAlOgKwKYsQIvCcKIse5
nl1iXIo7F0VxLAm6AUQ218t14fyxLwyb+oPm+O5oMFKsnC1llIQBAVS4QRCv
LVT7gUCVZEoNLcrYh4TFNojZrBvrJs5AiXn0MUdb0KWt4+yEw2v5oyRYmsE/
fuaCKga91KIRaOPoA6sUtlTcRQejartIIM+gUXB3SoqAiADnsZ3h5h6FKkf+
XJRhP5IZ0EgjcIlE38XbNygmqnuJ4un3QoCEqNFJZQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bROGWCBQC1T2955W2HgzyzlK6VfXEKyWTBB/VNbpHy4Ew8GsOqPXvCw03WHd
8k70k/Xaht9+/1aS0gaDyci9BU0vNbcKrfcPdJoctuciYIt2HmRUnYeg5Qnv
wD85pgDjlENXr7/1xyeSdzEWWYHkWi4CUOJjgpi/hKYreTtsaTcIFsRDJxh8
47OKnt6RoyWbsMp2/5GW5APEuIcuUfxynfqJkrl3MQFFVwEOEO67VA6TOhsZ
3uZU6jHIVeiJIfX+Fa0UfO75RLiDlPv9DE2rDR45bx59TKbbtKpv20cMQ9/a
IViDZ3/LOAQmAYJpQlL1TWwDE6SM2jnlMZp80M0DPQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
CKzLj4cQrw5NdGzyIKvx2zqPCvgfT7SMZM6AbAB+Q3I6rV2qM3NpRw34L8tJ
H+rEKvPukePLihqmBAiWLwjiRTRP8DfoUFr9+oAVzKrCCghDhpZs3Go8i+Qu
sWCPVV2zmDhID6ztX6OVXrbWACd3EC0j7/zMnghxoioASAhCPBrn1yJIXWOj
9W2MY9QECRHVgCNJlR6rueMudwx9YOCAE8wEb7h/sZjtJy/lclSrfoqAEEdY
eqwC6Q3ncF87ByoU8eVRlywa96R4I83TCRdGIt694uo+UTqwU6MWKbXDFuxv
0zISUszhDiggQaiFvmWCnZK4Etdd1iDA60i6SdVypQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
BfgL1NU57BiQrky0ka+cThvykXojCRo5vYhh8rzplihR8huSo50DFzvPj48J
u7LizGdDeG8XW5x2GpxY+YwM8HQyeMOSxBg/LEn5q5WA/FcWQ4lV3g0ziT9I
grxqv6RDmowg/xhbwEL+yCOWsR1lSQDRdh+RsumNzb5XcQxNUAA=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
ELpPOTunsC/6kCEghkx9KrfTMjrOfJhk/YB5mgWqhlloaHlCIT+iVfe5qe1J
pMEi6EQS0Fb7+LreEzr3I/93HuVIhV5pk2a6B8MGJ5jKEPYDvjCyjFcXP/hI
4JhRIIzVOGZRzLEFeCqy7ESbd5foMBwEsl2TXI0HHeqrNPqXIuKHMwF83r+X
hhqxAsC/NqKCGZqSg7E9ivoeDmG/D8PSOwZ2rgzm+ldaJxOk0LxFk9TVq59U
PtDMwRrcjospQNX+i9iIxxiRqCyqP4WjXnXj6QDcdg12/KzKnQONYMgd2BD7
3HPM+zt3lUhOXqhCCiLb9+nkje7/rX2XJzqdOFnn/fDzFWPk/HrpfnNpzdRG
mX2tUuKYsMg94pmzYyC3zwWX5k7cFLUNmYU1FfHlA0RtlTOetPZ+vnrbREz/
z8UgkMOkGSML9VLVqWOJslF9Gl1W/ZBfrtgeL2OQXjA4Tt1g173JbaPo3mE4
b72HMcyq07HB1CWPyAwe4iAUfq8Og04G


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
HmTIVtdlYNtHRVyCegCCp3MR1qo0zTaL+/eqUI8wcdczhdqL+Hbs9freXBP1
IPFY8AdADGcEigKDfmoDftEfqsnvzV+j7pyOpMgsY/AXX/sVuiE47VDK4bxZ
ucy4Hg6ZUWI5AUBI/eM9oyZlv593+O37IPRFW7xcI6UjTlAKoPk=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ONwCNa7UI2PJbF2e8tjPmQaHtO7ljgCNJ10dDpp2XvT1xUvPahxEDeroHuPh
QWgqACrsFqrs+A+8WsEYzftLuVViVrXTINVuXbEo1+0iawbjVXq1GEXUjh6T
bxBEjVMOGWl+X2A+OIeTVOVSPIiK5q1IU40MMp/94Xkp5irfkGc=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 10608)
`pragma protect data_block
RHIxu4y1JmWLaQKw05C2KSCvju1UQhFTNCGmdqI29DtSJ78qUNg1o8hmChP1
lDk2dAUqI8aJUa/fSx70vZ94n5ILsfiSKSP+pPfh8PTttKPEImGFf3hegjjx
A1c3Azde6THDb45BogcAz8dVYBWfw97bBK327Zm0q108R6ju1xJqR8CwZCLK
F8x3QkgrNnc3VU3N3IvRhSMPcpMYKU9MIhC1wGUwqPDo4IQS+tHd6WPRQe/o
7ea/F1jQwK+4m0Vu2jZEi6kOU+IGHF5b4IIGZVR2iMkKzGxe7jq6UgGS1vS0
LsY2IA1GrcbvWTYJorkiS97AeIW2Czut/OD02FM7rGSOvbKE9NkYGqsP0wMY
RnhYXq3T4NHfLaOQqhhus46ufr6T5a6Uf5kRNZmliCpYycO8VFKEgl9ByxxK
8pi+RoWiV0/OC2p+b9UKKVko1kvV+Ioh7xQtScO6u2b7JOILXtVq28tBj/gX
W0vqoriL7euqFBQYXeUQkiDS0DFIODNeeAFDOtT9KRMzkvgfpIJwJq4g1JZF
ifwjAR5Dp84bB2fhpFCuevCWlSHxwXnargjoPUslGV6iHeZhSbdJVxqt1lQv
Ivscf85DAQhC+ml1WQ+ZbRiqxt/XSW+wQ8nxCSrFiHU5rprWB12rZmGCJlj+
VW+MSg4k0RZ5XjyBW0jkCY+L5QmUaj+m67aVe8by3B88lrolRD74i8+ld/Di
U7YhQK2IXMbmKz7z83q67kGnq7HngFsoC2fXQq3ZTgqjeJ6S08FMUcLJvrGH
udM1mlnfZ2yE7iE0OtmzOI53lykJOek04A6ozl6H2gdOLAZuk378IsQFdghj
NO4F91VxuY0EN95J6D6yq2MDEMNKL5W0JFnHcwgvB0wuynKd8S2wHhDlUmJW
cA25aXEcBVulWsPjNlDW229yVWO5KEtRUhtmsvyFHez/q1Bmth6mmMVhKOhN
w+n4jreYA2vU+w+DPW67RhtU8pdh5e/yReMpgKg5OjBXttTTrvBGepJ9BksF
Gb2crtTWYsGEsDxjcYTOh9KhBuquxwrqlfZg1OnyH+xdD5hZ4traPzWtOBdi
6GeSctxAS0A4auLSxYWb1e2FaHyzkiXtoX5qw9IxxLRx//I4rsQtRUbdAHyF
p+Gp+EDhYLhD3Hqua4wZju8i9b+SalLNX6/B+rzOYxbRIEcR2p/MJAFE4cu/
JBc/JOuILa1ZjNToVj9uFiI8SZekF62dxO77nh9RoQbnMqhI7ZkGIop1inyV
TbRfmYvbQz+UlkBcfA64nwhe9odcSaVLzD/fKFEmPVvC34DLJvsfP0TTFf7d
+75m1YU5craRqhQD/GkKkQjYIJ7YVcWqw2XUFiqptGxLhy/Zd9BbOur17KhK
N9EzdLRRgIAdis/ydtncQ43wTYk+tETq+NFLvmbbCuZvyXSCRhCAthRcwxOJ
lGVJj4fHfxLRjmljqJhI+TdYyKIB0F+ik4+Mmp6avlpYZKOK9gtIOt/OJ9pZ
rvQuezXKi2Mpe6rKUuA1zNNaPiW1JKmbhhQecwDmX33dswYUx636bWHaxDB7
NiY+4nw86wDXmfjFd/ko/3H+65ecuBDCzSawk6MLb0Duo5yLU9xV5pr3aYx5
MF4N8QCwQYd0i1M0dulX3SRpKWpDTWK83YVdDJAcbiO+cSBzT6HWNIUDFOJd
J2kWruYMrhSVFZBnhJ3gOg/h01mCi74c3AEcBJSCdJoKE66oDQ3bgK+2fzBn
0hhTP/yMv40vJPPUjaK0dQKF5bcMN7cByqfbpkUJxpbk2lfImELE0CcdRlQO
ibN23wQ1+bc9G9hA2ik02oGd8BHkwWxr7zB1+uBKGjqillmPrDL9kTWCDLnb
2biR+JZTKEYMqTAWDxi1wFP1VaDf6wfCcNT8TbQvRi9y4s6OVkdK9A2nqf8g
5Rco00al7Y6m0J7XTpWyRaPVAwZIwyq3ffUplwTmcP4XFPUSIRecR9I1j0Sz
dYO6apTxKUcNAPGuKwzdp1xPRh/IvorrvZlaoX/tqrjExrQ6WTD8G/OtJZDO
XpvNXO+BfwVX57VCZycZEGTco/UszXam1U8nr2RArGQftty+XEjkiimOpsk/
nPPTMXwc4T8ieI5Eyw12u1Ah4iea5LTF26FnqLsU/xcJvjV3s8BFBabTmxi+
Uqx2I/+kAIiKFTMppKtEtRz8PfJvJpRSl3Gi9rKlWsMLWWige1hxO3HXjjjn
WNg2809TQxdmPuSw6R5iAeOidZObgAeuMncSBlag8Tqoi+NW0jboBuZXhpQN
llWXJt9JvH02RqsFupYUD3SuqpQflFlSTDs1+OVKgGH+j2nD2BOnyeBFNaUO
TeqAl1gTYtXb9HbhaQ/ttEkIOQHahVGDfvnVsPLUxT5liMsZhmCWUt7sxHnH
HYCcgRgi6XMpixIrOHF17YXZ5HPfGfkPqOl6iaKXphTD/v6+wFeatuC8GTH5
k2e8JatZXNBV2acYKrA/J7jhj7MhtglWcjeDnOV08jGFLMm1cw1SZAjNLkHO
yDDKXLoMOLFI+WhY2pMPsNLWLGUaFNlLSHF1ermYhGr7hUtQX7hnhRWlEmFH
7IgAXDXeUedB9sych3I9EO2AFeZVLDheV5E2145B61vJbryW2qc6+9gs6fVC
RU+jU2QONFEKmAZTa9IZQ++ZGW7F2eETPQs/sB3bM/0NlwoBALiimt5PiZMC
oI0zQ7+u3l7PPhYKhb0p830dWf+AwOKa4Pf1WObGAweg6MkHfAKmpzzKLCYb
uS3hgfbd3nnxtyrMJuDqWh7dErulfWDaaeqSEB3aPTCeiaDbwT1C1i3gU6YG
uelk2Z9OiTeF/6EmZs+6vQNC/XUAt/pK7290D+GhrqEdkCNon5GzjttriBDP
gIrnMygYwkCnSN/a2VHfl0chC/Bb2jrNyp5IWsN7g0/B6Pv0VeA3W2hD9Ano
uWbUBkzuBIXkaV8IsAgz+WWaOcZnslvvnLfMLUeFnsRLnHsMGaOmGY9EJZMc
3NZqAMunfpYJ1hUPwDr33BeIBrhxPPJK5vKmqO6RRhBYuHHFyzLyn6VypzGX
QH6WArhadCjpobXa1t+h4UhCksQF1TZeWioKargM1oqV1DFTBhWuSPmLWBOH
qbqfAvSJPLwrVReQqjD14c2VI5ico1uHV39TNUlnN1h5DRuaEcEffoyT7XIS
+gWroz2DJF6Af841iVveMldbRlzp+dyd5eE4ZO7erDSv/o2kTiwZr5pCNKFf
u7ef8Z0PuZ7ZTE+OkIePGroZLl2wZgNG4kOKH6AfiHjjXWbnfsXxDWk8hWQP
JqF2bl2tWKf9CKBajrEuq4Ki0YejkfO9/lbxBmEan4T35zSVlVY41cDfCEWa
9vZosL51TL/k1M+Va6QApglZGYlkFxhhloo/clX9vj4QZ0yH3SpTgzoJcgSd
sgW4OOETLXiNxeU6lobGQWoFVehms19i/J1xOmVp1VuH9t8RNfv6zTPqJUsW
gC6p07/wPVNoQxw6QAqLoE/OanOqVcYdFtfS07ixNlTioA47zVCSKNTVhw2h
Xlp3PT8m3wUntISEZpnF+pE3AV1Mp0XOwOT0RsZ+n+z+5pZYKmKYDTckRrQF
zXVJZHEVWL8vxxeY4UlFTjeRUAipQxbpmLdsPt5+8tdybRMVtM5MDlQvPV1c
mU8DkVLjHo6H5u/vAFXZOzuaeiSCMNNWDPcpLwJEikV2vcx4T6bmhNh/Om+I
x3z7VNcDr6/giwGg/gCkwQYgHuuZjepZNoy9x0DTaHT2qcLeOLaqqtJqFGpI
bCSzwJ0VIcjsGnbNdNiJ14v1jZ8G7b4Oq8A+TG3fP6+Nd9QpgOjN62PpBBVn
3sZw+cWFGCaoxD/ac05vCXQcMGG8yFYluE8gmMSSXESNsCWjZg1A/5M1B23X
24faF/LVdMNSKmYkoQZWnSmJNGIBa18Y+qUTPD9uIDl4yloS1hDtuLiD9KtK
/vNHhitRVK0DRT5coDPdc4zRobx0rjs3lByQHC81vYhtFZ2TaqLKwrO70S5y
QPmkM6/zCSd88Cxbekx0LyKQI3QuPhSZXttOkvbkivyuHUXbkzVw6VmJIT8K
5fyIBxkRDQf/VEm9jGyO+MMpJCc8X0ZRyGWF3PIYV9k92gPn+EBo+Jjyn5Sh
Fi22VgV/zzhkr6ycowLCxsEubGEL1oW2Ccvv4vHnd+kQJ1//cDUrUePMIUQx
3LchGfte77ZIuM/9bZa19eFrhN+xlWSzfDODrlXt6yChUyZtrwHsA/pD3LBJ
cXB+pSZ6fndqZniag467I9eyYi//VTQpViAEsTPBp0TnbHi+NIfkF91gjHPk
FkxNS8e0qxQaZ/TL6cd5tYqOj2BwTUmAAFL9t3rinVctqjzqVi1+62AhaRqM
I/3lIEPTgvZRV127GzX9M41USY/dILezbxZmVpVzaQt42q8O49lXx0uOqCzX
OhOhcDXgpZybcovrtLJEQp4Cz7I0FxkHg5HrWAlKvVFlNBM2TaqcOG2NkNQa
H28ABg2NlKFh+uAsYidnP5jh1/KiTt1T1gX4Map7+NVBO/ZTIYnX12ifNuWy
lCr7sRexgQJ8Bq/Y4ptsF3g/H0VkcK7mP1OAtACTw/ypOHldmlUPglCd2ssR
GCDUhUMLDJcI6HJF+c8696quA6Y0TkjSJT1B/8hJHx0Hf66dMqYzyFPUTBNk
g76yiQgtnNF/CD7k/KtfJQd7tNE9PIF+pxaxLXiWEnaTijYvFbCP9gcTPTK5
vrDXIL2Qv8uU8kEYXDK7GVR6QcVbLv+MmvpQhZWB+rudciOHTkD0tA0dHrkZ
Q0NzBVQis6aOPvKLVu9Qwqf0xYdgests4N8dHB1m397S2BJCJTb/0ybO6oqZ
g5vy0M6ksjyJQk9JjjEPpnOFbW3NYPwSLLhIRrXUbK3eDAOTIZTsJyJ29IWg
EWbMlFBSlzOUSwsgJZJLMqG7rebPYnzyFm+sCRSydUNmyWfk5Xf8UfidyR1e
1K5a8pPSc+XCxBwRgKjE8Vmkbq4iX6axBYbwvUjF6DWZclVdnz9vbU+7NjOF
YNLN4I8Ru5yQJk5ABBbDZ2k25gMU3AkmZt1c6LUt4EUixLDR1sPCbyhGeS37
aygmlVkV5gLy1mRqENUVqktprNA+MloMuX9zB0wKWjPlS4VR2TbcW+L/cIer
ciH5cyvP8bT07JCUZXoBzJyBn1v3xJsuZKZCdITEop1fDgqTTbuLJGQ3BjZg
HmDwiByFZPbfgfWQxDsgDSQsvnQg+iBSxQ0ouN08UftGbOdIjUgTQEYZ4ZXe
KRpm1/fi4plO2JBTptyA7CTwExBO+DElerhWHvAnkLo9AQcxpJXSx+JZqLyF
+apqe9e0cYi5ykNVUUYEvr9jAh8Q/nH4WJslkPXJmEmTTpdvYfU0wtx7OZUz
S31lORpctS6vnWxnYA4wy4x7HnOqMFc+53VadeLKdm1skvHKb10kSTzgE8Y0
apd6nc9IBxg9ZCwnOdc02PKsUcfh4PE5PgfY/njWPkJsH53YhlEAaaG4ws3F
jLT8CNbXKBiImpPxKUoTnxMQlgJBBKZKKcrVsghXNT5Xr8DUBp4HZrxmqLJk
Wly+Ua9luQNRI5XghMe0qICmFHr92M9apE8gEEF/PiwGvpzQMxl2KlRgdMti
Y0T5U99UN9m6l2V4dn0StBu2J+RKPMo3MowHH3NnyCSr5Wo8TarHsICArQcT
/JUAVYXh9IZCs/dIsg6W7VSy7EiBC3KP9Ufuxt4dMZDG3aRA2XxOYaGbR/x+
4jD5maJYz6ppyEhdyFPSBwKxeHeoPMvR9aCG5ATmm2F4Kl6/cLXY6Ht7GhRA
rFhh3mEfFCxScxz6MYYgBpSzWC8O7DMwI++cwWpQojlZJK3R9aSk2Tfs6Fy/
Y0tkO79L+hIXCZkHZGRODsTv3zQzWroIWCZTY2gPHDfM5IPgHGL5MUscKXTz
QP7tn+IYWRq0Ee6dH5fwtYAuAPSj/pSrbVguG+lzCUyWnnAk+03i/+GHVrcP
7jrXxQXy8/sZLumeCzIdTJm6t411LYaSZM8T0VFkmJAQAJO3dOxdN77hOjHU
tIOdfKR+SP0nT4RRhe32qIHLrsLUBuMCB3dQ8m/KCIMCT1c1w+bXFJzzwODe
c/mP4nr1cpkW/ZLpopjeEj2L1W4G7hgOsfGXoK/QB28ZX+/yugq0v8+e+T3k
QtiKWp0KTvvpBkF7kYMVrANqJ3nVkCT7E/myROasnq3Iv8S/iJTveMAHw4IQ
7EZYXvjiDRLNoyvOjt2z3lxwHX0+fqtGGsMCAkRtjfv7E7VUAQg8uixQar4B
IlkbI4h9JMRrR/4m4j9/7wzFeQWCpEur37w+bjr1qpe8p4zDhm+7OUPM+hGh
7MALJ3d4c/Imk+dsrjsljL+UhSjx6BYqZCVOFS8y3+Fzq50X7DE1FfBO0Vwk
uzubjRYqoEp+dNWI0blSbaetW3CLCOEPTR0cgN8xFmE0LEaTPil5vZFdFjXg
0+T2Ke7/V2dOjeLy3GB0g+hh6/p4GTDxs/3nKVhEBCY1l2aSqkzdI10EMBUq
C5n6LEh7j1wSRwKgnY8iQppX+YF866hZM4nsA5Lf6lTQS18rOx80aACezJmN
/lLUZzqHj3z3sIk7o/y73bg3l0dFI8QYnX3Pykcc5RSWVqs2+NMaxU/EzluQ
nYQL4YKnfX7B8XACA6X4hglJXqn4LTYIxpXtKVJ04UPkx1nBhH1TXpQnnjs/
RCtJ1eErmYYzuj3bDMkWd+Smf0T/wWhwZ9YuVNafHZX1Ohg/Q8UJjUFGDSSd
e4+CA6IZaqnXdDtu6E02KHYDE7Nkc6oidZKs3E9+raXwh28NYBrXNWDuY8pg
gxoD8gfWHV2sTXIbIt1FvNPnSgV+2npSAcgBqE4vi5VGCE+f60oguDOPXtC8
u6FJ1xHgQrOaun0wct6O7mgldC4JFR15BMHAQxRK0Uc0ijRifd97R+zuHsMf
IV6zwxbWBh6PHm4mvABAmJFVCWWhGmZ8bu3PL9vY1ur2J06lRCUf5aHwqI4r
qnm3kGrrwldXJXCJySt9bhwWLodxZN12KUP8J5Tmyo39HLAMn0HL9u0kaHoy
fK1kzcuKoICOaDWKGsmI/y4qkq8XkMwyMuUEhkafIn9/q1M/4VO3ZexLmHSE
wV+ieCTOZp5SSOG2+JWUiaXabYVoXIctaS0zO51WKZLcQ2eCqD1wP4LxTr1T
Xipgm/vjWBi2s8tZmQYg01sFD/h6gg0nQpLzSXfUuoWMP1uBb2ik33bfu0o2
8pxaPuKATlCjSX6j0AFEFNmV+gRglFGNFBEaqUs+XIq0NudOaoKQS7IugQjH
qU8ABfoumj0f9rJvY9vkbFOYQLTiWywWPqib1IvhEAGSvhcbt7NIbgOYOY0G
QG/NE0aMq9e8quGS68KOdLQWgkJh/nhMm60FM5s/8K8HHTiqyijLxKSaEF23
HR5N4VPF9qnPR3Zpb/QT1XOBNEvVQcauUIX+Gp7bpGQE5EWbw5FH6SGJWfPj
nzSc8WuF4foP9gflHzsXXOs6nm+eVQ4mXSCQf8wjJehaO7cwWvkKBNYsFH8c
yLFdafuZvmJUV1DirO5XjFKgSE/G8Jt2DgjX2PWR6bl80Rt+asFI6QOhDU20
N4e3DQNxJUk6fOV8I05vL4/eP0Xs1Qgtfbq3lKYHjxwJkdIWAiH3hseC9pob
qRnN9bjuioxxM1GZNsKejuLhkZeEYqB4q9XkkQWa4LaFSHfeRZtuz51v4C2u
EXeApWFvYOg4wuMQj3R3MF7ITAnBL2YXoawNWW58E2sOcCZSfNQO5tToUvB0
1NUEXS63dI0KVV9qxMd5t+vKsdnEVE11JoFwhd/tQG0gsyFSZ6BV4m+LwpsA
6uVHc/OtarSDrublVHZmuQtzPkpXjrFHp3DUi6kgGIqJChukzqJcDEtF+33q
0guapS4eHVIRng1uFLCxzwRnwFHjpV8fqv3oIyxJlBJKQNnaWPscdk7jPuCc
wXBqRBlCcnxc+vFASf4Njd11+tI2ZzpKByeGSxnlmkKdHe/pQE7EUewAO1ZE
PqndBnIu6sT9P7gEmWZXrBXNBx0VJU40GaTXC9WHmyk1COuMNEbPEmedXgXd
4wWHZBgSbmdIfZoHKWfSR5O9PH8C824FKxtaCtV6vPoiWUavGk0FS4XIZt88
xzd6xdBmcIzJtJM0DS/MA2Wl46Fa/4aKqFnf3vZB5kC8qzQDhqzJNpMX/C7n
ZyVo72yLfUp/vg5kb58ebIfTbdxf+vEExgXt/8FBvKB4Ai/peQgVK0VLoW25
RdwFeq7DqCJ51a1Z/Uj7IOUPcBH0mUS61kRIx3Mrw3rqC6RHPZ1jZvzlOS2s
DPTBWRRCWCWJQW6X86dEQ2W99oKo9BoxD+EKcSNE9XGTIuRW6kSGuNl1iOAo
3TCLQCGlZWwnjvSYJrJ522YjHB4rLpslVDDCVqioP66yUMzwE3zILRi5Ijy6
/8lUKdQr0uaUGUtGnpJjj6xLn0Z89hc3voY1zi6do+RHBn0eXma4+APIqscN
i3l8I6WmAoPnNoOJBbQuxfd2dsLmScWNb/6lCmyxB+DLJjiNw4W8X4h82Rsz
t0TQJcR9Yjmovu/piWtZleqSkYjE29gnYywpVp/t6O0Ep8v5JMd/TMl4hMvO
UR38VZIkbSXOuA5jm1FTHxKVFhsN30d8tLaCZOfHV2gGjkkXoWCWflHogoPZ
ViUF9u82VL3KT4BLcw8eO4kTmeKj7G9fT90zPeffipyf+9KMra0+5P1fmDEY
u2hDwi8anFT5nCflcOvGwKGGTSzwlXAn2X0f669uSTYdxMxvxBumgZDfh1Ua
fzqPgKy4l5LCsAWmcvlKTzH2BX1otaEk2tEmd0XtvxQv/e2Wuo1PE1bGP+R0
YkZaPew7ieoAyYIxjnu/nCgo9JudPQGGoZ0AfeG53ZDFhAg3AnwcFRlmSyPm
feqsXfXVRa4UkIfCIxpZMmbPKuyBU/ZqPeqcSzh9QS0EkJ5wlLb60DwmetcX
zRlDt77v9u/qi7y0I+7XrdJiux8/U2ZdEhtJE3tA9ogfJM/qszbpwRPGnvAA
N7TmzUINsmksrrqhE818vtnFo22kLNcrsMRB3E+F5/GwoKpz7bKHkz5fFvg0
y8oOvGs7CadgmDV/riYZivzwh9c8qQhAa3Gy3Wd1nfWHnc22UBxPKY50QKen
5YFkxMjpGU+Kmp8LI27N4xg30nMqjWBkxGyQFMvCV0gDCMHnuR/hxepS1Fgc
j6hudMyNPpYvKQzrRD+69X2b6rnyCBOC7FAEbAYxKVbmealMMi64DJMrjHGC
XDgG6p96R9Zvfs+/VLe8WQXADDY1vJVVPasy+cLWsgqDV7r4ullTco3k2xnW
8ddQaGbGHdIq5Wf+Jr4tseWswyhD6qvnvHDe3eF/3RsyU3xviIyOX2MZPsF3
+1WIqeGG3WQoCb1mn8nG4PTC9zMF1OLmYtvxO8Y8LIjprUxxitBoIqH+qdNS
KtjuR4UsZvV5ebG21JJ7dFkbm0noUFojKG1QdkqPyE9JlzFadKXR0wTW9udZ
srDPQ5yVIBeiCywzik0DaztkBbCvIQR7i/uSd9ChFSKnTXgRzZfGYZ6EZ6eY
Us1M+1E7TACIYSm5I0qIa/H2+hk4ArbAJpxQ3/Az6N4+pUSkXuM0GrmUilf/
PTgG/1EjgFxLdeWjRNasL9OdSQjrEigK8/Eb05JB5pLvPYPeMfBaf9OHXkjT
D5U1uczDzikcbgxG7yXeePfDvSQ3HRrMC4+7D3++0Xylh5uSv31W/ERfxgDg
JChumeh2C5NL/ouX148qZmjG+XnqYN6ggt96enV3+WA4tMmFf1rhhx3xFh/e
m7ufHEHTtGKzUCkLmK6JhZcXTVz+dIWIs6CVBUBWQEeJAAMgelxtM893ElkT
c2aqoleP1/1HO7e56IkV46SWcYhsx0lQ4i0WLzX94/SnYseBbXLfblx8BoSo
VjLTTQpR/HeGOadok1K0xDm35sEdLSAux4kninefdlueI8up9SAH0F+zbo21
dbvRKFcldbfIMT0I2uJyaR3ixTnH9Fkne77pIjWlAHBPXY4eJ/uhF6kruO30
DVxAAiump4x/AB6mCAQnrXPxOiHBhdai6RD78NhPhFq+dHwHU6m8UKhLmgGu
NzfGjl8IXnWBrUhpm+oOf/lVWBBBacVDD3Jy6GfqC6ifKxZ0r+BShIaDdenR
qwYQMGUFXVtcslhD5+VW5VtGlWMsoKQjzpKcMl31ewVOnpmrq8+ti2nqvobR
s477MhAUaC4WAtfBNvIKAg5s7usty0TuzdWfRQG/8WG51NP1JM0C1X8LT7NS
QgcUlIrOyRgbPKxIsz+PH0ap9qWT7QXbehPY2pBRNtOKhSkW0VwS+GyBcPlV
ln4cmXE5XaPLfcw/mWJwD2fq74Mwt55RY2GKQFYR1plifcsk8df/0AIuoMZ9
v1YWa6+g9cQX1neBhKCSY8qIufkM0WFBWVqa0UaABzvHXAHlqypz5UPoZWsp
Yin220l/+q/ZzbEWoHqN71JLNhbVFyfyd7Fwn1P+4JQSFOIowbk7BrmMINej
6/L1CV51OLyojzKkeEthc1m3+CwTYCosj3mq1mwXdLVd7QfbQNVQSOFIbuCW
O4v6yB0wLyPbg5cx/St4AbSOgRwcSFoPl4c6EWaIP0HOd3+oaNaL+og0DoE8
avm0QxEnKaW/O3fX+OOU+rXGlctQOg223vFsee0+znBrmVaNKUG3pVGDwuLw
unO2RUjetohD7i6H6Wgk1CpC9jzL5J2IGEajgG64OtoRmyLF+feYlXl2y3Ua
N3FcnEGNn3TTfzpUwBkWyaxM4FHESylxp6dpPSDH0vGwlD7ZcRTt3UIxg2xR
jVHiQJWamufpjNvVz9zdrG0U6U7/kOFDnDDMThDr8PZUnMNFgL8hNg9GcD6s
KOs9Q0L2I8Nt/e63wxr4/IMYLBQ8yzhSxExB8gBswVlz8jB2y/ZDoxPInTp2
s0fXSgJ6iv10QGEHISqN4gHpUcQrJU8/2yQZy1trV7sz5VL83/vgz0T+Qe0D
Pmq8mM76elvtBnsSu1RonCPptx7YBtvehbeRTetRqagNRu+PkRLYBn0wov28
SnQoJdIElY4ULiHj+Dby25SszjKwyfOx5zJH0zmo5dCiYVkDCnzIC2xJuh7h
DMpMuqaaGS/I4TfYYqlNENND1Gb+Gv2/jr+Rav/0vpv6DMKtWs8XyxppJU/F
ObRwGq+6lH3lBswGvwDL5WFTNs0mnUVyhEW5Sz4WChMEHWtCAyXlQUgddqMT
UuVE2fF4yrPBcoycCJEJG8ztUAeBIvPbNZJ8tn0ePppS2ocX5AIA2Mi61Gmg
E4hYDcBikM5zVMjM9shgsYEYcVOz8ZE/v91H12j8f/fY4XT0Rd5eZ8iipMxZ
NGB7RX8g4uExZ85F6F6nM3IlR7QJXVwaxDnJWkhfOI7OyRNp1+KA5aRL6K2o
rfsqPYd2vLIZacvCQaOGMrOecqqtJiWEawgK3SZsCvUfZkccanz/5+9C+dbM
VyYMDKmuaFrwEayAvn5FVlI7GGusem5wA7WhRHIQ9YcQVhj54VZDlXJJNKLE
c3AzvwixKTD+CjT5vCTflJkkf/E1jgZvKtdF7d/uYupkKXfZPR8oFdMdjG69
AaDO1jGgbBLqORGCtpGmGpoEcfbEOqcTUzjgazpxjkscl2MrhnsZstm89Dw9
Rz9i3QadfrvwEscYr0u0hwi4R7646ACfZjZlrJx0NLTJSkcADXMj15HCh+c7
LPqzEVJrROsJeSZhjmSMNYLB9rS+TFaIp3cfmkTkxBdvk5aYsTOTtkvT3SaD
nDFbfkDSZppTKsXVoNg/uBrogTrLSbgAX4bVKH1+xUL6JMawGvx3hwtLmmoI
+riyHeLZBMuG1XOGbFAy73BS3ac/pz+MSVVggkTXi6cJD+6/zTIs1ymDC2wR
Z/OJWhPWeQTiURff2ysWOmqOXTaTGjYZcHwYlSYQMYBu4XpUjevChfv1b74q
cKqR0FmvvWwq/QLvex/DxgRRCL/ceHK5ql6x8P1FdD68MdatHjtYrdXSlTrt
D3yVHFHtqgs7wafMzY690A0ZQcFFlDde+AnaCc6Zss7+0UpyYfgbYcZuJFTU
G8zJ8xCusPVE/mU19jB1Qieg9b6J0nskGGghXgfBmmPqy3MqoKtoL+Mis9ip
fweAtQs1BX8POqUNxhyNJJNQ4bP8LPkVhM72cAUuP9HWmZpeUZl8XAr5MmKk
LgBCTvc58s9Mws0ZIJksenoVQY2JgWWQQXUyt+5nY0BD/gQzI9q0QGSAQ2iv
yNaSbVZGOH6cnj9y2LS9czcnE57KO/n/Qx59rUmySxE6CTOSCeiqjYDaalTo
y38rJx4g0ovxku3YQpBHc/DpttmxF8FTpXKkgThXi93w2B7kM9f1Jwb7gYrm
83+AkIbXnZjIjF8rTo24QRjMXqE/xR7cj3O9G3YbhtAoFQtLy+bTgOWRsmtB
394gnQJBMGqLd+OoAp3Ojl5vrfDSxRx08L0RMioaMu4JUDbT8W9DxXged5Wr
JCbxBJTgVAUrwGf6ogWmsomMnvXFURKa+MssZ4AvIQglDOx8GHmWyOI1md7r
Buetv4da78v53u7fbI67Vqs9+9A/cwtpdxfRGDPU1x+P2GSSDt8EvB4xEj+X
PEQeif8nHh8SZkvo1p5U4HzIJ/1NvsVqIGDUKn/BD/8tmMvBZ1dxs9Ron/So
ATY1Mihz/OKbJ9bebDqp7KjS/CP2r+luFegM71dG+aAD1VMyYTm3ky+hf5cC
CAaRbM9Dnoj0Ssw8CoJPcfP263RUT0Q5f5iLLlqJrtw5xkslHFY1Ddyre2z1
Vnm650TBLn/24Fxp6fcb1hIZMzTlIt/2TUB4VMQXP7in+PhhAUJdPAuHKTux
xV7jrCd6wthmKU/FrFR3IDIbVYBEEe26GYsYwJ8sq/mi74/tNH0v/7EM8Ar+
WSFLzf8gWpa8J0/cFgMvffF3Od4moLvT8xpkHojdQ94Fx9YiugMKYfZJBhG/
0mbs3IShcaNV6QgNX0AKLD7bADhzlxAbXf/3cQj7NuMOiWG4a5OKm6SfXvrx
Wa5t8aU5I7Yo6XgWO+NgQag6tUARJ5XhD9fL23IC63IZebfhtO6mp7Ob0si9
CJcPLYUV1Q6H7PRY6EvXWgcDJOyEnJpJbOaqEJWyeaSavXeGMbmFGJMnCXAI
Xzc1HeZiyU+qe0O1kTktOljHQCJERPPbCmU/wTyPB8WuNRsINlzjrVSv2gbp
yti/TBPiU2Mxc/Jaon9pp7pXbSnhHdc/bnBwttPJo0PCaG6+pNkZSw1mRz9i
QuFPRB40va73xgn5KF5L9bcL8l9PtpenpPh0seA5d5OpN3eyE20I2uvUxbaF
g2kfIi0/GAOZTxxB8kWV+nSNaMcrJgVK2x7YRu2yEWDB/jG8mKeT02R1/lXH
/IuX/gqRsFRXyFUkNCoqa5rtTtYHpfeEXCc8fKKrya2ueWChV9C7TzyiaaAA
VeOLkV9vZwVNdrYgQriWb+G+LioMJGVwWKQKHOH3n/qw8s5ugNXxlz2HzdMD
rxKNyc1uFxW97PjR1qQe56h7FsQqxxPfVSar7r/6EtILK+RZxBeMUQN1fDC3
XabNSSV22c0aXosV9169v2jyq3NQ7izjRUl1yqXViNgdZe5ygkFYX+SW2PIr
BzHGViPMjjUzMF6WEasOazFSEQ/UInCj66A0ZAjqXfJP6EBtiN590z5slKvI
N8SKLUK5kIPBTV3j3B+D5uVDN3XQ7jtZ8cKu0/wDak0Z4/7KQa62fnwX6tCI
S7mTV1HTQrG/bMHcBw26lWy2cM+ui55GysLBC00Rf1Xnz+gNlpfvGWqliGK3
BD5kdOl8LvYDYEYZ2527b2w9bL/kpj1/qXvghasrG2m0SWA8OOwHv9h7psQ4
1jsDwrs8pcQKLljjO/5QkTZPmQEp04OfSCo8LlX4Meawm/ZO8N6qWv7xENiI
v4SQcr8z3BA6J+weNPjV4fCH4QBJQNv/Br7/md1I4exJjxpErxPebzSOCKbU
rDBvGMdcmEWULOwDV9PRE+hwOK2mt3s59OakoqYgospIqAx5IT0ncKmyH9iM
LuLWWw8aHbIb139wbEZm1lizGGLF5lIxqXeoUL+B7liC

`pragma protect end_protected
