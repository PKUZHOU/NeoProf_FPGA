// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
0uRzxKC+XTCknga8eJ8CR6EYu5hZZ+b7N5t6aoiAoyrpAlBX+055X/hTjsn4
NP8HqYoj20iM5bkoyw6S4ZJL7TUqY0fKFU0sdyJnSqI6ZW8/IwFYc3NxvrEx
lH9Xr6w9MQq8pCezpXglMd8eMx/WCZ0cFfT8EmB4Wml/vyiXWRAqe/aB2Hjc
mIgTcdk+mx6tbwSnanu566Ah58lA2OxJ+H86drFqLoxaWyyqknGwXYb1pulS
/b4baSWbNCNFiPwQxFR4tCwskrPGBR7KJ7Y/TKqVyhYIUKi1KyH9qNucsQFr
3/d7lrKNwZ6WnLB4NTptHTca/jHXwrMLATet9y05EA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VGXoS2862HbF96nNYj7kah8F/FMN9f7Lyz+UNw1dFE2qwIB5Ln9zwNPFDysn
/KHWlh8CoCRmMxuTsg/JBt58rI/alMRxMf+e++UhQJwd3dJ2A+jW2owjCu+i
MItUaLRACH7rnawzx0w6GcEXvI/IinLiFMV8ns5ZDo02o4kHqUYFCZQUlrpJ
CdFqncI+zaTCelvFwE5HRc2RrX7Io/fLFNK2XADrk0iga/xlL/gGk8IVutdS
bOstxCjFv2/RzgJe2uRofpVqV9zRqXrnH1nqh+grCTD6kimkow+6WwjDQKgS
HcHj8T+masO9OegS1w/W6ou7DKLHhldHlnLz8gnggw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Q7gDFsQkPqx31oqIl2YJnaynSRzGfpb/SqRSdDcstwoQkEB/be5pTD7dy5/L
YH83JDhvGM4WuE3eDnYW3zU2F6mpxct0FmcM6gAuv875RJAg0C4DEGwATvW2
TZKVy0UZyNuWoAG77uBPMMD7HO/CXvKr8qKTfNVyrwecfW8qDjN9bFnxjzIk
rY5qOLu8F1RtH18MOWd44bdPH0CeqpORGh4lRTMthIqyNhKijA20deeKj2nE
1iwZrhebNw3VowBV3UYoHOT7tmtlAY+7EajYlVjixvewClT6nkSRlq7eFRGx
y9u/D2m0bshb79vy6dflMIKLDaH4N6aR6m0pPtMn1w==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
iV/bRyRGI3qJiCkk37D6bU1NuW0r8a6B/VUmMts5UrpKUDeFZhB2r3Baqb4I
lYv+Wi0XXmjUpenfeSQnQXrxiaCsB55R9MleZEtAX8Ic/4/B0IiCPhzJmSSs
qFhI6kPpJ2yHIWIfyjS9umUNnUnRTdiMjdlnB+MDO6vTnR2WD88=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
N5vQoMkQybnJnaTuk80ZLyLEnGF4x6Axg7KpovODOLl3kvLHLJ36iLZmt9TV
W4vtzcTsj5wwYTQogFtWlUfcnuC+dazXjA0bNV8fggxRUu8cZU/6jZoJ1n2z
hUQlp9vjrzLHlCBTB6K/ybxptf7VhrWjK7UvQu0hnRc8Vc1ZXMcUAzhpWnx0
nfZnAGeXcNEGow2vezQdC7HDrKVPj03DDuR3jjQ+gFPz5xkr1Adl+sneXbRE
IGQPSprKzS7BqJ1yguimaM2ZZL+pfAvBwPLzHFfTDET7Uml57NDWGzzXwPy9
+/P5ITzXIUgtiyM0CxXOinLHbOhCQI7JkJ+8EC43Eo/BDLoMdc+0UH9GPaIw
C/1ZweRfPUztWcDosrCVtPHn1TX7AY1HiwX7Q4PFCd5viJDjVusrBBNQ7Ff4
X2hXn/9RNSa9WS0Dvz9KiXH2KoIAk58Wkaj4dBNRohNrM+TaK2E5/4Uqib5p
TcfR+eYacv1NF0/7gEpvhyuFSsNKcaJ/


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
B4TqJWmH6AK4cWtGQpZ6K/RCFqPEmz1SOddI4BiQDD9M4durxA9Y0IuzreYa
lLRrH7dWQ4yfO9DVTX93ui0dIIH5EyxTJnJoYdAUYjBe1oSuVrXI1QfZwi3C
BBoVw2TpdQhsXJ5QA/FqtXYbTn7AhPNCKzzMi3IEBFf6DRo9Dlc=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
oyVbM5Hr4EqTc3+HOeJAnydvW3A9jiKpukrPRkelNzbaih2MXuH1b9Pr5YNQ
Dj9c5cmifcYCnHpF85IESeq15w3HLZv0ru6EMe6+YQfDmfHldn6mqSs/oxzL
Lu6NlXtPsjTPhEg9iqEs15Tzi8CWsaWdTzLXZKIU+8PRMwPLs5A=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 31120)
`pragma protect data_block
4GW7feBQ8yweIgTong1O0v+7cZexQRZXyW9xwbhQ0uk1P3dzLsAsr6XxL7D/
l+YlfuWXLm5A/wXX9IrRcF4PguS+TmqkSYpF2zJSDR0eIyoUHeOJnKXQfZ8J
WyUp+wfODckNiRFL+yiNOL9Yh1w+bb+d2rB6ALN6gmCGqn1rDv/Cznjv5aSV
/5XCOJJWMW2a9YU02XcqFrrEPIyoQqygBrb0LcvXYvCG2vOVyp92ISb+RkFz
PBbPpBXiAPhfXOnz7upYg+zCJ5YoXYNi+RJpIU45k/UCcmkap/MbPAvkK0gP
CcNIvrC95/4IGhHdyuHZowBZteByOHN+7HoPOlXesurKL11DSQXuEs+kTXif
nw8cT8gFHCIBLn4xKhpKZsT8MJmgZ/gbjybhLiJC7nkmPDyes9T1WMykA0NX
tTBSsznUmW5wo/SdxZgEnE99qINQb1MAbws3KKHB2t50wSrDvNtSRZ+PzItC
bVPrPSPm0rd0G//PfuZ3SbEfx/yNsAG4BCxqQ20rE4iESIaPBRen+ABJh85E
6FghC7F/iKiQrsQIsw2t4ZdnwZJKqUEDuBiqpF9xNRCC4YpdY5z+ZYbcfUoi
MFJHxegXqJRjBJ/Ec5DPcYmJsPa6PZ5M3JYUhZwtlvHFhuVD2gts5/+aFLOg
UU2Ph0OImzkr8Jwa0O9+gFxowmT5K4fJdtiqosCKLlVBZnwvTxk9fNN33vlG
57rmIQnk6Adz7hDBCJrqhygAA7sJJp8+s5pDCyI/vqXElXN5FsxHzDynnRd9
sKW9B2knUQxMbtUu5CSpHBbuI3+sGz3r2AIki3EHorH35Omp/fo8MNBFdplW
TSJKALHxrfbOkqrzjpgPMIvCs6K3nLDG5ip1WNGAsXxhXXwIn8F1rH7WnRwY
wqQlvU9hI4OhQIbTt53+vZk6cMvbupIL/Rac4yWX/6vMMV3SbkuQXKnZwvlF
cYO29WV7DqF1Dg0qOHHrxvDZPBeWGVquBEP/coZgY+L17sni5e3KR36q7lTc
nu5AJtY8cr1RUu+Egomvc649QI8Vgefsg8h8KI2wEVHbynw345heDrxO5Agx
moADKfBg2mJC4X8CgRFa1pYqtrdA810bbGQTrIqgw1ScWFJTNMJKuTbueE/r
13YA8hJiyvAU29NpvMuC/MSs3fastaTWmGuNmjvJ9rKIxmHdV+73fXh9B0SN
Wa4xLABgg5l0hNlDvcGFqu45E9L7OpIxA2MgfAwq0hNUOI4BYILhrwAImHKJ
iANTTyZ1HSpJdkQunpljWd2C0vbemzM+F+VafpjVaRNBazkJsSSwbZPNAd/P
4dUs7JbRyKo43ws82PLj9yFOe5qInlrk9egPdbgk2Fi0uGBKVpMWtHB53dAa
f88Xqj2UUn2081cDOwsRlVx6h0u+ui6Cq9zVxFUkKbA5iuf+me1i4V/lbRcG
+IP91zNEDlLEQ1esGCuWEdfvLiR1CcmmUB9IMSNiFH9cgOglqsaQKFDEQEw2
T2P90NJqZoFm3Vw+gNWhWHgHXV8iKteiaCk7hn2mGw5D3VILQ0nz1AwuVkkr
5lKiHXoMIlv/sHVF2MaYmebElJHyIpbismt87aow1lCga9N0c/A1QeTyrGCu
0sRzZ2BfHE9bfjAnw4nX+V3D4Z+T7/L3+j3LmK5BOH/5JVMTtarv1o0MQKsX
qqoZAL1Q5yUCDveWkBZzHetF0wmeyjjJYR8vYuBKU8YcvFdzSsmnvLRn+Xwo
wqOqHGGJWe9DxG6JbeIIWAMqX5bzoNrzzGsa7dmK6kOsjMy/dUszvjxC5Edd
M2fj/oTdql+OaPLQSQUmzOOZeZHNXCCQGWUih+qZSY1t/cZI8miM/vcXECVW
wAbZKnocT69ZN5FHuHWn+kfsWzCtPnU1nceupNwDDJUKlkeM3kJwZCO04FSJ
YeXCPAHXIzNvvpoZ8Si2e79rxCNRto9bqyb4Dmsw5hnlDUlPfb9naP/x+TtO
6DDBgdhuv64UDmJOsepBoRI11VODCGf7BUBybnpeQo+zFtXdvipj6SdMDGcX
uxqglHmUUkCTwhQOy+LP+4GbuOgMgwhWOekC3h9aYE6Gvs5cEWIwdGAzpjsm
xpB25hAfLbvpOvdsL8d4jJ7rHDaa75De9DBqiK4YNyVzkBnq+xJ9KhRVfX2X
dUOSiaYWjUGejsYZzqoEbfKzRxvYIcWk5Dhlv49w9g+YHSdbJUaojsgYnx1m
H0iHw2MMBwygMxxTe3Hd58KiE0bkmXhkI/3yOfwU7s4ZHFfKrxrjFzu3S/rE
S+HzEDTkTF6h2ynjm23oa/HP84jOr/lOIfZ5ohH9+ge+ZiNuStykDL83SKhd
F9Jq+HmTeUkd+IwDabD6o/xxO/gYnTVSQ1AbWqbW+D5OxIw/amfdCIcKC/dV
LzEoWSsgQYRj8/iD/tJMkEdUkJhFOfP7OS8fU4aG+wWCRRXL2MbUVvPqk6My
Zs/is6joJf9Z8ArnGJMTRwUnBgw39fnA+kaLEGjU/FYRTgzaXA7WiEtXE4bz
jecdEgVnX9FiOkEsO++8uhVCGLjfe6uvE4PJKjnNmaupKkgY1X/RFlQr09Tr
t0EBBartbd8MFr0/TVpHAqFxTw31WQLDXWy/xHiAMO3MGxkpNKVIWeY2ECkm
ivwYPAQqJ2g0DRMSaWtMI95BAh29LKE3aL95zvEALaoDo305ghC1KZcaRNEM
5BCjuiQ3ZD4lCHiIC2FgAzdFXaHIVPmyQDEKtr80KRndCMpTNVup6IXrUQXw
8s56XVqqJ1GA0mZxn7frS3kaMqKASLiBZRfS6AgNEp4iFaBVToa0Rx2bVd/w
RKFFbtBBMQFHI5XE2fY36wB4Mma16CrekDOX2zDFe8C+7I7tvGVTFwgf58jG
mdIVKhKTCXshPH/c3RoUHPzl1Jfls2/lPNb8Ceg6WiIrxNEqWlx+7nEfVHiU
6I95R/JrC5qusw66Ro8L8kninV30KIX3Dj8UHwRGflNd5GiEdQX502tKUIIb
lbTXt4NTX5LrIV4yD2iMds7d7ClZYiFkeGGN6oL8fEYcg43aCUfwxjcc+jHR
iLwI5Jo4GGreV0lgNfk6TYypG4ovkzqg3TTwzZF7wEl45o7CKpXpDHYlozoy
i6pWfgCuL1yC7kdjDF010G+Wu7TSvgyeN7S4WrAv8j5P6K+UVoWmxqoovfdN
3rWNi/uHL2pKeDVOjqte/oFO9++k/VyrQ79C86mh0gB9M+VOCoc5IHGfyeoI
pDaqv9X52i26qqWRUJmI/PLDd3hlsg0Asj45UBLbzOuhEgfTV4O3JHJa5Thf
3MzCRiFWnTRqx+9yNOLmr6DnPJ9/IAaXG5vA37tFaFCGVPgCLDr2ynTRUF8L
vRPCIHq3cgFoTQj0sEoju8eQEi9Lgvx00U1tW5BROw1yy64htdylxIzGntN7
bvu+jjcJXEU0UqQ4k+JCf5fixujAtgdyNy+inAGg83xiwrj9xG6k7zKtN7wh
+zCZr+pf5xj8NK5sSgjozSoLFGA2CN4rfkYq22UPRoB2qCs/ol8n8DR7WUxY
8CNwBJU5earWJEXsKAiwlN2/FaHgu2983l8PxCI9gDc883hynjspBex1JIG3
79h/FMtoMtwQo1AAuwKXm5laDcxXdfNc1MvopEXWcwiu9S7UCwzXXN4EJ27M
YNtzjSAzGLE+xcVtuY/HA7/aUAu4NgfDtbD0emVNyJJgW8k7vb3t9DmWAGaM
Txsdw4ZmDbBVG2rD/5Qyd6XFxfvZIhqgE4E4PKO8988GLPo9I+icO+KoB0qF
sO6AiIleC8U1lx6DTfiI2TRLEnkxYOj4FEW1+w260G71S6IKIRTZLfPy0l4g
Wi3LNTfRbnhMoNLroFvflsUh7vAwZCJYsalYEwfmvmxt2OvyWJ+HKM2B9H39
kjEJjEjaszos43riAoPZNjKb0gyrltmvWEc7LzxRSCCzRxKeKMcDQrYrkEqS
UG66k49cEgVpxiSmMi3jH2k9jWcjGThJlbDUiz3Yqz3ptJqKyo4YBIG2sXoo
soldq6qF3uD8L44T7gdJdx5hMvRrOe/HxO5p8N16fbYDgOzFXw8ERpFnziy/
9NyMBpXJDJ9qRbAJlpIF+F15j2YJue0VtMgWP/fQ+ZKCXKzQDPLatlvzYOn3
8iLOASMJLoA5SpdRAJcsXqUjz4nl4sp4VOeCE9lEFl7h0tqz/jnvykNPrEV0
4xoGedyGeE7CvE/uLOecS8szUdn0yumSJAaUFjB6DVPJkCAjLtnWYz0lM1CQ
UZnUgbU+QuYRm/PJiVmqDR8FUSZ3BXtMNm30elBjWv6sICdhIJTjGGOCK1mA
Npj1zhoS0lnbARAVYRCyvAtgJXSzIVrWy/Mv7SkWQXVTobkzLevOVXPwF2jm
zqywKsjFntad3Pa0QW6YpnVwCdoia7P9Zb5ypy2mvA+EsfHCCTnTigZzOYRw
3RFL0SgKVqSa6Dy18yxNyOx62RA0bWOHyt/FClFXoyg9fgJTlSijr4CgM6HQ
6iD1ZTOkrbour8wW7pLrXdhqnbfqNFN3yqY0tyHekdygBeVSNEKlvmC+Nv5s
CFxSSsjAG0RJ0Qth1c9mra3NPCMnWLhVCuYwbpOKMoMXKTx3HVFSJEnqErLg
mu35nMU5qX/FECimXRxu3Q6ndjYWMQ8uHauNomgtIldmwKZf7OJx5lEjculc
62Ip4R94Tpm3JV2nqVytO40Kdlfl/uuK3v2uIQUokOMncQd/DOCaLofVgNBV
iqvIlJ+3RwnjQOqQHLyp3a0mwF+WptThX7fBFcBaETeRQJgaoATP1U1EBG47
gq30lWwE2sIqgzRrUDDJegxLWxriBb4DJ3ZHgpR1KWxxoYVDIcriHxBqFdT2
rfQqubnurOi+PTkck4TNMmAStWDwRoKFuMzpT07cZfvx8xpoe6AEbadFZzy3
w9n0TgGdLt8TaFIsdj2G9pPkTbMqs5QDjJO0bqQk7btmJhxCQrlZlCWyVIjd
mXlmEIw98TUVRp97d2TBdX/mzxVeLRJyeW/F9OdwIHVi8wjx2Xa058tg1j7E
ANgYIyOXnltDALg4zoCv7thYhpmdV3Bgp8zk0DDxslFb4arw87XXycOtl3RO
n3pGisNVZGfGqoV4PBWHbiZUEa/A1A99b5BxaaF/6A56YcaZ/luIQ49zEipn
Yw0JmDHsG1mattPJwLeJYQOwLMa5pKfP7jUbSGMXqe3m2kjniTuagWROVNzA
zI2ees1H0cGZukvsab4hg/QVGC+APWGium4Sl5dQOJAjY+kGlZfsA1H7YoME
gBFqn+t9kfnYhf3x0CQ8eLVt9pqT3WMpw9oMrvzpYWjljUYVNixKeNDbWpNt
nUswb/PmJvjxXYp4J5fNDKVoo9gX+zyucuWlyweStTaR2xMepQIHqgvDjHAx
lUkclVK7hmhVZj+UJkxWJWo6pAMK1BPoOoz0n//H8XNK3wP9EcZSkbCxJvWN
X6QmSyUCGHVihZBrjkOGufbnJSSB7seFcqy/AS0a1XOi4jVUgyAeT7GJB9oP
C5E7T4oL/RhvyDQHfN4dMr2RPjlMT4LJ66oTz2mdFc2aIVuW/f7UZnGK2rlo
XGen0oB67/NwAypdDrn5TdcdQ/WPetZFVArRl7Jxq7NdjDberKDzDHLRCmAo
rxualM0KvfqNCKb7aYTwTd4ayssEvH6CNb6STTs8vlNdEkqlaGk/V3J4L7Lt
RZXJYun8NsigPlTUqeZ0dT08yUFDAUwdW0ibbRiUiGcGe+0uW4uC5aALC8Jk
3mUXITF/NpOJYX4otXX4aP/obH+vchcaj2OOYiB1nYVO88KQAlVDswAoZYQF
XJJm+f2zhO74g/mTO7VB88/7l1Ow7TuIJt1J02XyHOUqDnSiGJ78ENutVJuT
VcDu5Xbu8+WlQFJv/FHerYT0K4j1aQ5KeKpfZAPepsqU11odsfgfmKvlEaeh
uMBAKKQsovsEVjIGtuqH5klSZNUV5UX6Bo3YOWzrijUgK1/o8SquJkCDN9hH
w5/WNgGxWoNIdZMYwdhO9qlcnQtvedOetTmL2BxXQq7vN2Na7CqSx3YjT/SB
M4Apvm6itX4jaeVASOWn4Pser1cK2MySjrSayRLqacsG0KxJdSN2JchjEU6p
xveBiGj0cU+gb4/cPUaZilMV2MUT4xIw3kzBGvCm46XjwR85k4Zf4gy9U1yn
Q3SfgmGFx79T6pEcyt/jcx0eKhRFj0hst3Ky/oQtVgD6atHMoauKskq3QEJT
o1wneFuIGY1PgKR6qCrbEzT5cJlXVuAaJ0FLKr720E53x9frycYe6H3nNSkT
7+3UDAAnQjypHmf5tcXJC+/kmp3oCffOJco6FFb8SAFp6GRiL2DH7LahDpLr
T1uGefEWG8wm05An4rJGDIzqJyzErE5pRnXEzHHHGPhdVYvatTDtG5S6qhgs
oQFr5F+K+P9jhzSleuM9wMiVD4FvyKqCVNDj60jh5dAEU7k+U6UMyrHLRYz0
FKWfrCesfvatosRABtnmct5UYz8PtYD5ACJQXZlT6YJ2SQWEBHWO1ljT7Ife
HxRT2TtSs6y/j6T/ZoC6Gf4q1LuOHIq6XJAkL71JIPdqZRvDbLouzsr/NrQ3
Ay3bxZYA2f7I0dcrFIdLfW4NS3CwK5Dn0LsXMvCN9YDmjr2QwftsY+ImcTeH
hOiXL2+dDGq63VSUic1LPve+b9dogQs3NZRCQGIlCxasWmg5UkOdBndY0xjX
5PHzh9nFxIz9nw/801lNof2kWLMrVtm+TLM1qexj4UEo9wID+83XfFquW2Zc
8ddv/2qsNEyw0ZT3F25aYBxVXFlg02rgvr1YJxrh7ppPsWLsS4FPPZ+Ru1UW
/7UjTsO6C+k0nYzA1hE5MhB/ipjAXjOieZVqAz/x5HyK5NAJpPQLMYWYJlXJ
v2c9fjabHlqqMvQLxdcXlqEmXmT7we31yA9xtxvUJIz/vOrZS97GzIN461dG
iUC/OEinDBnyHxMocbBqGq9HR8+wcrimwUf+urq2/rML3VVl/kzKHUj4DR8o
XW455XAaWwF5nkrmDrN8KXm9LhetJxPgjrH2JkJeQ83dYo2zkKv14/BH3XO4
QbZdZ7dCq+WN4Ri0aJlt3W57yLmhxU6imjfWU/hTcNvRHq5QBwr8/PbUteD1
yCvNH2HLYsZnr75nQ+chCoe9ApwQWWsuqUU0hZ8TKdykIl9zpgqadLEEDOjG
47GaGEKqHbVJ+rXIELxAzdAQBDLlGcGqjIO++kcC4ZeOELa4Zc42RCVIHKE/
s/XQFEKVmI/EL6tuL+isRSj8tKpb2ocC5dIDO9BU8tjRZsVk4QjaFetZs8Qa
F4vCIMsfMf2KLvO+Ck9qDiz0PmVGBcmUvORpn47ARIyATjcZ12zioWN9TzCe
oZiq0mNTI2Fij5maJJ6MHmMrG3kRTVphTT1BiZMGK51ZVNGxE5i3cfijcjS+
K7mGltEHjRQEvaA49LhXM8qAnUMq9UGsM8MALCUR1lDq//jSHlvQ4o1ULH3V
VJsZdHicOORa4l/FGmBVsCdFLLEBF8BsQSUfAcymhyUmWQD0218aPXqvE2Bq
Rq0Tbfq1kgNRU1RgondM03RzccIb3SG7UanMbBQjMla+DV5fQolC4JfIpg8C
dJPPrdTVqG47yDquE4GwT60fUjiUiO2iK/LERVkqsVfhIXGqwvTC26WkeTUH
TA6m6eDZ+Yeoltm4Wf3jvzyR/iiJjO8YhyLgVmKdCVZC5A7zVG/aAcGMVpyF
Y6QpM/l/Hf6+4FwOfa0Rk8smzLE5ihcyjs8CmE4a636wr/Ze0kaqN9eF2+9n
ommhOt7UAWXU47h1RjXmslMfpmt6bjU6lq6Gp6rQ5obwuGdQhP/wsOBMDtMM
UR4nQkXtBOxvoUrNut0HKbe0fJo/374h9QU5uh+hlbzU9cf9eW+7LMS7vdMM
oW0DfzJnUwAZqfXJyAsj8GZnpswpJE0jSdCTSeZX6a8ILdh/WmAa5N0PpWAz
eq6t5+ZAiMpPpOk3VQyy+jknHEYKUDVfycS7sqzu68mjZ2EbDGKZ4v8tYjfC
JHKxmlncMOO33kg6AWfntgtGd4yWDqNcjQLSw1nkX8kfd3KneJG9uZ1lYY4/
MeGD1nVivxFdnw4wwQtcDvfieIOdJKOWYPz6IwuuBxjJjlMI11lCwa6LcXDt
QKLoKNgBIIO6qDUWMVPD7D9FAXDAUrTf0p8yw+x4uScValI2xlGSMJOfDpMC
QG0HBWCK+FiZ2P2tWEWINeNCNv/rG1tzeZ8PaHvlxW9m8/uEzfwRwbcm8KtL
16X6rOkFGLlDsG5XtiezYST31CdEKKbwg++tuVsdaAgVoH1YbxI8f30Sm+q/
BBn901gNWVtXtv+jzc2Wx3qe4CKu2t3tJ28uLHG7cc354gBy/PrwAhZ3uKZO
oVxvPMTB5yfoB7TDJjb2174wPYIcwR/qkunlWv//08difPwpwa44vBuF6/oH
lYGoo3Z5sD42slABWH9cPayMOMLj+w45YFi63yez+yuRkScKhje4Q6EdHC9K
hboVDEFOr4vprCZI7KSHigHkjWdTtW0tC4iSHW3wFQHVzoWU4jY5rvVnINcG
DfA4S0y7FE+Dz1NgoRT1ZftQTUAKjWwK3cRqV1OH19I2C4EnDjmauBaEbjz9
PK9njew/bt7SqAIxkTaYGF5T7p2hinlfu4hVKM+UT6pBTgrnTNFojJkzoslY
YuiR3pEmI4Ff/sb23pZV/y9sSH6nBqp95gJC3k3K1Yho9QhhSSN7dwMQsnjD
ON+pgfGNn/ZryRC8g9Slvbg0p8OsJoxy+on9S3rchmSiL1pKLVAViAsqgr/9
AtMvrHj6Y0JIj04U5fRt2KGVx8U0rrUGjg5u6TekW8ZdDK8KnYnRG9I4bBkg
fuQ2ARcqz+sN3vmLkWTrZNvPdvkaNB/op7GL826K2gMhtMcb0DlaRdUTlvuX
ECZ4ubpicnv3YTKJMPbN+MmnQu1JB/lLIS0CF6SBV12XJzcK4R0DuH0Iea6e
voArmIWYZods79krDNdJLzFavFHqj+Qk1TWfs+XOGEQvX3iY24+01SaBFPMz
VYr0Y96s+y3MN2tOSVRECxpde34ZqV31cMp5m0Num4qh68ZW8m3lCWj35gLo
+GRnIMnclnV6ZlFKFLXkhGacSy99XSss/W+kKZqugkbuD6SWgCfHa8CPrmxz
wHy8udGoUpPVKAWapadepeK293xoOvGQKVt2eU1vOqdqWvvJ3a+ZlBUTohRJ
yGZEM/KrL7Rlvd713JHctbEXAx8wC8jgm7WiW0evW11+MJEYmMpfxz6z07Sq
jXi3i9ND5RwsCaTGxuVVwT9vJ4+izeV6jCcoNIvPioLbNBPbdXoLTNMltjeD
rniA3O8noRh+jRqe6c12cMPhY6XWJaWPo5w9Uwou32QvDb/mLCTZK1yolB/5
RMME/7b3WyUNeMXLMDpBA/+JreOb6bSC9sxmUfu2rYpLAMhOUCjJkn+XhcJr
zGpPhuO/FpvnATIPJUsnRP9aL60kTIvzh/HMbVmO9xErcG+4L+2pRJAGUllD
qrC7ruuyXQ2B1va9gZ1ZJckjt3WCWYzgtOsnetOStf2fA+9nOkSd3Qqi8w5N
UmZJzvTtiLBDu8XDwfJ1oY3JSiZntibjCV0ozYd1M1rxmp5ODG1yACZSvELa
h0rtgvl72qD5rGKuIGvscmfo+a7f2ftPrOwpk9DxweoxpXxHFUEKPB0RwDNO
HBHHrXqozlTcP/MR4xpo0Au20XdvGs9weRu6JBrPMnkBMAsugn0WoIfgeIWI
i7KFF0rLnWKfRVmL8vW1mHSKg7NKqk4lhUBF3yjwkIsQXLWixW/HdXlsbyo/
098qY3opEXNGhnj70LJPuS5e8/3mlFBzrcb8rjjUwjxCgLEYVRAsUWkCCjBf
TfwYmx0YQvsLYixBagtadP5DsyojRICfgZxi1IAFgUJ45k/3jPJ3wwrUa2J7
bSfmWV4giF/ZLQZ3ZlECkc7Q5w+Y5w6shHzhnLqfqCCqhyZfsAZhAD7WyzD4
tyoHql0aD58qerdbVjvW1ZPiCGerbwwg2eOR/u+QwSzeWjDX0lJriLtHk4I8
lXLSA/5m/8b+JOjVTmc13zennMpS1TqOxYlE4vupWvL1TDinDfQqQbfrSBbm
uBWdmqKbZ02L4TI+keTXIyx7OjMLeu/fNSi21de/TxOS2smM0CrrE4sCEDTf
d/H83Ly/5Pw0slPbImj4MDQg3l9yKOuZBP9yc8KSyhp1Lpqq+/fJowP43VAM
ygWqLqaBCaMFtOLHEt1Rdx3QCZ2sbmBTfM+7eQvZiapskTGhYGEizoQaejTe
MRT1vozVIYrT5ffQEAdU73UIq4GeK6cpRiVEPTv+//iGL0uLlPO4q4j4Cplj
kcaUL30C/dUkgQoqtdKZxiPEvXrhrh2BHOCtIduZ6N8NyqPzH0w2WCE9Z0FU
ZbhHcZuqRnTPoJB59mGV2CyCyEBwYkRiEEfc3sHJOneli4wislIydzAnzSwg
gSvfkXCy8+/P7mPhXNVwGigjc59+cCVOhuEtprBB8Zd7xqsCYdX960fc2WaT
q2uXFjaDOJYkht6kBqQJPCor/jtezmyCnAQ7duqDrIvy9uWbJ6rdhIYvMyu/
N01hlbtmxQ5UpUisZxDaTRyhlmWBWtS24+ld3iCnru+HqkBmTDEc3PWxoLzr
nJARAIdbJcprGeKsq6a5uIIQpT097wSJEEfShNZbmJjjAnr8LUG51k0Rj8f4
KhS5AJG5vFy0bG2gTunHhiC9kBJg8l2jdPDIA4tG22aEQtqxOrhrgyStfuQW
pFarKQfE+1qCUCEv/kEXZPQ6zVuDwcg+bdyNQVFaMCYDU5c+bOduLTf+iW5p
sfpH8HYSONkFCSU6EferbU5l2DxBZ8TJSgcfDgirDdqGC6plNfoMApnNwmxv
5ZkicPyzMTYWW78yvSZ10aek4JE0wUDLo+CzxO/vH3W1Pv2qPKGP1ugflk1l
tmVddYnBiZMNwyYlzdXNQYamuPOPCDiK5DVn1cXyj6H6we3FHh27jSG5LKeX
yTFTKGXe/PylYAWVnPttvg9290CHzL4xAjMQmVzqgbDZ4QUvdir00YExQ1IR
Tnp5vdaMkG2n4+kBGglpIWFtFrprChERnmEY2Jb/nsVAMbpse5CYdgy15qxN
/ixhEILN/F0YFmcV0beBxVJsWJ/0iVskCIL962UCRvUHxmrYsv+QzRveFn79
UIxQDOyFms+FE+tcQ2bKaq2rXQpTJBh5mwaGo9iqx9H8ye2EINlZku0HfPVD
zOvlkXcp2FLYqp+03qei4yptqg9IM5B2Emg86M7yijfmqycvRZVBedZrcfFR
uXtpWKl2duhR+5IpNNjX4Rpfl/xWmby4nbr7iHyIRQbBYZ19thA4VPpTVRYh
b9bBjpg8I42TdRIjNlPC0njBOPr+VMEgeu3FpKJjog6ki+vHPuLO679vGpHn
EDYdEFm82IV1QMznLzWuIULRseciQdRXPtfG2uUGSPqjJIQspM95OypEmO4O
pkGVxumy4/ih17uQs2ab1Rpt9nGeKWR3rUkw0Ez8YXAHbMZtRxgPQRe2wlnl
IWoXDzs2wakSQVNjvPbYZtNIXHpskDpJ7LXAs7u4mOtBiG3LkbX9/9gq/iKq
dK7fjkY4KeH89EkpP8mAcSdY/IsSijtVovnRA/HmHNpjIeHE8ASjgsVe77Gr
W7TNHD21dfEi8sX8UIUufJ1HnFHmUbuxio1aUE4AoVJEQdTr1r0yeIAf/v+E
hvszZfEMDsxFqWDCKLwWEPl/CQPztK6ZHLQvkVMlKVivLzC0gZaHeiVJoQG3
wcsULaWvCKSAj8AHNWE8yWPFwQThx9riZtSqI9qIGYxvq3tHFOn4NthpUp+p
MtKJ6uWkx91lgsI74YO9avJpF/eQY5L4gShim1lGbQ5kNsOjsahr4gxUOazf
oLfo9h37bNjHuml2pPHXyZarOSPda+yaIKEpF8fiUz9jBNwqY4sQm5o+SVW7
SP5yOjP3cCBCRUqTGzhmlMLG9vvkoNqtBElKF1oWPxm/ET8r4CYxZifXLqUO
+tNBlH7RUk/vvopMJrGNoE2s+o4nfDMLDekWmueN7UMl1Umkosd8j49vfa9y
7i0YTP4vHH/YTInbFYHY5TPxAUguHNXBuFGjmKFArYc7oX1egR5EnwW4yd5B
ExYngMc2p335b4DvV1iRDKeo4fLVEyFHyVGoj3Vm9rUoeVXdO5FLHiJHCzwq
TIjBWjs0HGNDZto0x8YobAv59i/Co+dLowiJMfX8FpCNsoJlSpeDIcDhtteH
rqqkzHQjFqS+3N55qOMb8Wx+S8KJu510G0XbJ80/xkXHibNG7egXGkNmgsN/
S726m39K8BAaMJ1eQ+RFk55sFuiBSw4Epbyi2lUcL5cLXsA7/726sxR+Vrww
HSogQqiG20STWhfN5gbcjgNENbPUzsnqod4I/OD5o6Km0fS3l/7bQar7xpEU
lkwSMOyV188F32DsxMmCiT+JQdmEw3sfklEKFl9ilGWakImqOGl64pE8yWgG
XwOln/8CJrI5HFvSdl3QQbNR3D7Kd2ktzW5W+u7GwCHyIWLci438xrICDCln
r9vBjbonkyq/u8hguLZThlIFrpwRHmeVGki0bHmedKnjFIDrbJZhmBasm7G0
SQwKEch9UjKSxvfzvOsF1eTiN0u4LIny0us+v7gX2gd7bbEStO4/aK4jC8VX
tKHaBlJ0WshC3fG+ejqbgO44Akwq+hJ79LVg3f6uVm1Y+Tl9DHMjiCCHghin
KVzCmQZMhE2SN+tUeMvrVX8a/WhtprcmL86BZAHsBz9HEPUdHWqSP58QOdg+
i3hIkOXtD8NOkVrq0ziLg6jXnVgzM8dNH2RlLmCs4R1QAtuzmgfzdzaqO5Ch
AuJDMS7JEMrpvIicAGrg+PWsASeW3r5yeHIWhbHnYFcgIO+zV419AYyWR9y7
Sn14M1rrt5hLEqPeaVrR5UiqeUbXyaGFqUMmRN3Z3TCGpaF8gwj2s4Z5agEP
AXbZeaYuSSwIO8qSd8wjJyxpv66/EEUUrlVn00AD1CwRc02IJu1r+Pr7DwDX
K7AfcgIYRVTKnr57REN8mKHVyGbCY2zxvr2sZ9OrOQ4lYaCjTTWjozQiqDZI
YSCe3vArxCYy8q9hcYGdbeYxojJPB36IW5/jTBtBtH5Lby/yL+6a8IrjfKQ4
u99B4153SRHcY8cVtX7+KdqvSqDQ1/UMNuxel33lBG6C2IfvB5vmRWt8qvsn
4j0GogW/kBhomqXvKylCqBZmR5OtzxenSsstQ+8XliwKtJSyAcjB/tngnsWo
wNySGvFyYsd5FEvqkrdwbU5wQtg2FJyk2JWRFKTGpoxDrGh3gi6L/UHszGgB
xI7VbVyIsBEwJf5Wj+SFdN0mt9AdzI18MrLY0SW0YJhGdWFYMDSES/4ShkgH
ylDdVW3jMw+OJyMuar5CB3UBjO2AXuRLsg4UbxIEMWOWVEXXMlTrzkxTIYjr
HrLOcMDihGQnSOyZXkk7vs6orqjVBTks+96vEqxwrRtC5KCybtvS+UltXfFy
4IbTxLfc+HstDzg59D0w4qNJ40c6LiusU/ZEhrXjPS+oRDurxzcBu79SZElP
CNrkdHOTJb7Mb6H1ALXrxRW263biGyV+1Tly9QiaAyi1bCA+dKlZvN3eMju/
EdIfd24PPLvH2EMzpG0BJ764/lowXvCZMUnDAEv06RB69F42uA9+blr8zASw
guTEJct1Q5kSciDh02fzsFcQLRXMHJMWwJwdnlHQR8w1xYgp37O1H+LhNKMI
30DW1eL7YLZssuiVhkCe2EtxeEHb7qQNxahAfVDbFd5OOyTQPvbGzCywFanM
/zMz6Lnu+h0BylHSige1q1uvuvVQW34KjYTpaSK4Fvdeui0Be+DBqO88BLTS
3PXlSFUbnP/v1DFT5YMn7KyXwTIYu9gCA1FVn21tmac+yfMrGIzKyWC5RYLV
Gb4YNHnLp3Ylkp9iRWYDFcl358I7NLYGX2HECQlRMpyD2aw6udMYz8Rmnh8w
l3X5KvrTbqjFaMwprQtlpVK6YNpliHhnhB6Y1fs6B0517uW/2Rz3PZ97clBe
BVM5qC/Tc8JXidVCB3SE4NS3RS9sB8qEqG9lI2L+jDRMEfAycJITu+xNhupQ
5Iv0lzS0k45DLDfapAvfvpwyaaAfW59EH428DtEp/WFMA76fj0Sj+11m8aK8
rk4Qi29A6CGbu9dblDPVRnuiQUvAtLwQgpvQPrcsv5MSRuaKcEfv2BO4WD/v
nYtNYGfmCYkhMegZAT6o9Kz6AKVuKhymj71bAB5+o+ra47lWOQrXwd2V//KK
e5/1o5fkV/dfXqE65+KdPPDQRZEF6c9ktdB7tm2bH/JmNGl5CA+zZw2Mbl2J
7MQknS2jyytXuOftqc3rCOG2DqFojSaceDVeGRTXimb6Auxv8bIHPncwq5wr
zMDb2+puu8IQQ65vYdfQ50tAIB7q/9Yoq2mV5cnvQlPSdl/UmFN/iJgzdn2u
r/+zRkpWAcHyKOnVM6qyu+n4yahCp8bzb2GwsyX8yIXdJ9OGYNy2+p2TRQiE
tkyf550nlDXVjTIP+7Uh169BPFA0y5kKVD90JhWfATvpCCra7MggnyCrhCSj
cPpdE59gTV3qS2fNjitic9UTiH9FQAtK8T81J/rd/lxXxBijq5b+B4kr0lLG
zC0kywfSYzkWCmiJz2LejhmBmV9yO4edVGukOkmIq8BDx0GCidvGNKA8bmfq
4qJ8tG7twYnGjs8Wgm5eNkDOS+lm8MTkVVn2EWHgYvApJN685q3XD0fg6aIy
KvhwREqhFLVoDiZXSDVW7cAS4Cu4QGrVEIPsASGeu2gyQxLj0Iv903sg4jsb
Rt3GYOpO5/Yp8jEZDiJOrranB62dV95gBmR7d78y/jCzrAUDD0bTlhOc9SeJ
rPDKF55Kkdb8slkiQvZDGXuJueG0NL/8kEoOIGp/4tYzKXp5QwR1hqBNciYC
IvGvahMaHG9QNUjYSyYj722V2ztlP54sETEipqyOQCSuUPPBp2QQr/dzeSZh
nUjy361CHsKLqwKZM43hBF6A6vz2M2WwapGSwJyn5JAL84UZgcMXcCcS/L2A
kfuv/mdkPG1T/lgkOaBx+c5yrcNkT/FqdJz502ztc/C6/OfN6HIv+Ne6uLri
4Zf+ZA8r1UfoByn44YHL5n9UCFfpSGGbAfhk7bwiPyV48o0PaQn+v8bNiAQS
TEAmzEDUU4NNLLc7R8n3xWePqkBI8BCx5hYvlHZzMTRbzg6sQzLabUGamizn
GdeImNht+jCAWp+7MqHn74iFUJ32Fra6XMd9mnc8fHLsYJYwoqKnCpk5MOof
29oLOJGsfK5zoxAJMKwU7BoZtt8N8/p2hfaK7eiFyDlgu9TN0UQD/dBU6kZp
/UyHnj0venC8e5Fg4IWXqIxBhRIjltnqanUOQzJDOo8b6H8CDhGLKQPBF7lS
CcHshuUmLeqtd83ElWAdS6uEh7bv5wBLLih4vR03CEy+WpGdKK+UAEY4gNQj
sH0hRsi/S5t1IpXsid13QkEpdfRLeeoqek0gV3HipIMxQkXAXu69Oa/OY38h
0MZ8+u5nozQPrj4XHfa+N9+ijzn/3Tjtk+dTrDWr9sHw/8242LL7KYvck8RA
oqyAAQzRsABpHtL01am8pplmYWPmL6EwfmAwTqC/xLq2H8SkZV9pbMcgpZVa
O1cyFPUA7G/MsEfH98//CAAozBhSzoIAzinW1cSt39CQjgKgyYaDciAmPOVS
gyizHOMYREpXXsfzBYziGQjvSOhVmlLdbyBQH0LoCBhPFHP/XnzBXtE7BfND
mRATNj/fPrwBRGTExKHvXbRAr7DHy5l6wBxwiyWaanpzqI4sGrt7MtT3A2C4
dQh5oFS+aKBLHOxuPsLoJEPX6e0YAtu92WaXOhBP+dpc4aoWSU0VCwo2EjRK
ZvXrJH8Z9tbXNkcp8qIA3XmykIJHB8as2gICVghmob3Gu+Xxe1oLO+bSts26
uTdq9iewakbSusVaiviADf64govvubZyFa/dEm5fEU4lVjUrKXGHO+5OcS7y
3fsnCX13rEeOFErtuRSbPpAL4GG9b9ftSZA7rGxntNAgbDjWU7zBjDQpv3yc
yIkrO01oic7a8G+SUK5FiMaBxjeHG/9OVqUXPcNyvVUSc2bnCt5W4GSeVY7r
0tbrpJdC5ZE1zyroOM0aY9fCcnj71SVBtlkzXjWkZvv8jGzmXUYV5OKMC+ki
TPm5khqyerzuedYdO97Qwu6Xy6WTMUczLaHWgpF9agbiR5P3AbqCdGWmUTkm
otbphfgK5U0j1BYW7DQnaFT03UU+baf0kKFkF2i3nvwBwttEy8sFHUPK+kDI
NJoLSjg1qfHUnrwLF2nKGFTct9sOuI+fPXkGR+HvcBhE8W8UE7tAEh4Mt7Yi
oAjDx7Zvew0vbhcLXWjX/4OBtwE48ijaFAsYmZ9I9c284AeQLXx5+jcnTX3o
FHLWSSMrH7TyFMUO+lf67IoxekgljMxztUjV2pV2D6CyYOiXbsT8Y5moQabt
+cZ6HEdBH4V/p1QszohbSXpU90sWzTdPT9O0spwYYwiwSoFRdB3EnAiuoAsx
Iwugpj/Bbw5Y6FnPEyLvImpxpj5UKxjbzM2wCfVVDjRGh9BGV1krRwLA7Kap
CdrGcA1UVfPtI0H+ODnySt7HtjLBD6t1TMLIgOl1GdSSysypS3c+XFKa2x+9
4SO5v5hT7RKENm1AWrrVjPYXFQIZh80AcfAYrYAJK4OBbHsmXVELalYjMKUm
1rOrcapSl8hEShxYVgAZtUGCM3GWH7kdFlynVQNfN3gd4/ROONxvhzHj9j1m
Pj3kel9tGqOTe/5gymeH21XvP6WzfDDElNQY6tE1z0h1I/8QI/BnLMv+SV6s
p5P/vu/La6sBxkPKvrCDrjUJgdYlfAnDKGIzXxXZ7nhWM/mbgK66s7zp/Qm8
fy9j95XFrTSM0dxBhNf8aYTVYMpbxJmqU+EKENnqC9DNfyrY9qd6avhw5XHw
Jzjbn9NRL8a+paauTcUWKkLB8Dj6ykZcCiL4Z3exHuFSZfZbeqBiTyGC18Z1
418ePUyRfnW4tuCVtt/71Z5Zuf2LylCz9qnzD4BlHPPfKGpWP7QNR5mCHhEx
UgxFRWhrbIFjEyWujlLHMzcXl0139gpYy8yiaDf3uyQ9y+OP4IWw3tX2QOQY
rtnOJU2SQAmAZb+1ifXZH9HvbtgpGwMJfICpEayFnS1eaUSZ5WmXWWUClEeG
FIkusLR8af/lgRD/hFnXi5/UuOZ1OlRiHE4uqyYiNIANl1gpYogU86NGMawf
VnyCeZGwIp6YnQ9rsJf5D2L9+KR8qnPtHMUjIylFsIqZSKT/OeAZauipMycq
iz39/AHsFEQgDd6aUI8M4reVFR5/jqc+ytNI7H0n0Uf0ejQ+CFY6zzJ3Fc0Z
qhQcrI/z1kUqJ5le90ELTECo6LRRYCEtkSucRGYdZkBVCSm/Ug4L8mvK7RP1
7TpGkV8NTr7XpMYUJbYo7Cj7Esv6Zx/9esC0H1Zb+R1/g3yJuMHouARHt/fZ
HQ3aY2STDip8W3QEh3/SBnStddCZwG+HNxuXMMYnSweqAN5XKEO9SSXit1/3
HfUzSOITNSdyFR2byusVWItB1H9W0KLO/0Ccj/zq3KX4O5kRcHh0BZfTofNb
JusXkbi5g5kxT8MUUK/hRlcMKLy/JSC/fcSG5MBlnW/a9SvrKI8JP72MKS03
Vukz+OE9UqGuFYg1hYrlx2liC8rTJJ9ekb8uJ1reQ5D7ab1TrCkAovpggXcS
acVSvmrGnGsPH2qfGfBK5irbPGPk++N9ePNyhXtMBsLc8KJW30+2eWiJyNad
Wye3yYLqIhD6JnLMODZXbk8NxO9CHRACiMsxunwD383DL8ig4HghPId7FxWs
TErn+qkHnAhJ6K696bzJfHrrppr3fWcTjuMbn1us23gDSDlX36TUwKfc+oMC
ZKqHxO1CHm3lBY1MDH8dNOC5GBntPXrPSIhvq3IGXoD9NNbajtke5Hr8IrcM
Oe1wWEMFTkDX1j+zZQzkL3SfYODqfFWuZpzsY4efnKDb5r8DrK7UITG+mvD/
ZFwvgKaHlfO9ToZdvBuYYSmIFpgXg1pKdShaKY57wQ12foKxnVzgFusVlGw2
J3ffj2+y6fq6YuC+CsZqT6BHXOUPItw1Q05kQGadJ5RbyZIOZIF2px3cgiDY
d3DZHKGZrLY97wZ8BW8WBYAriQq//b+8NI9iwiLexB7yEn7nz2dbnsMnE59J
/ByQweK9yNcnYBApMorkIDn3ba1czVbABKANB+k8VJH60+qazQ78WCiHP+wf
/IVzuIjMWVcbT5PgGAeZqbSEbEdt93xqoCSSUpmU5A2lu5I+aTzPryYhbIni
WGsiXFPyqAiLAXEg7PYN/2AC9KwD17DZQ1Jt8jgfSDnBZvEExO9WO+40pDq0
cS7G1mW5/vaKsCTqWGPyFHHlWOxDVoHxBFPIY0sPzWTp+9dP9C9Fqo20RSTm
9ZR/BNt3MjjphJEVNLp//ORVt2DvWT3UV5Oc6jbQR+1q4CFeD4T7L5wnRZ2/
06HMU6zIgxK8IRABH1fY1WSDrM5cyYh5cUMwZnjfXQOgdIyfXoFyYxF1YlC5
gLCs/H6zB00Al5LJBPGkDAzUsmFf777I1uNwMqb81283zm3qj1+lBzI9ahph
Y8dVVL4Beej3FQFfAINjbOaIPMEdyZYR2OwgXzp5+YflvMKRM1eAKvJ0575U
IMhgRXmWjoTYySSFTz6DiN/f7o3b/sI5Bc+BYVQ95v3g24eU/DOGsuUWwm/w
rICihep9NqZu1MaACKLPxRK0trQaxiOURiP+6s1fopRc+xxAoYzogEYZUvGz
yQLqqiaKxH3fAW8BYGN9d/Y7s3fyzcNaEH0o5aR/j3Kzl8Tqf3qOpJ14JCnb
BfKSD5AIZjSj9k+5hqGtLGkg+h871HbfsHMjJWAlAOjBRdz8KitZjRw8s0HR
xS4HJE2pImnf0SfJ6AIQCBWSPofeFpLecX60DgMx1cgqGAAJxw4GxUHHiPwU
VPiQdLgMN4GphtX4kTmK/f99z6cx7/hNZjWB5sE/rCeN4I1JEVQEe1QkPRM/
GfawC+6Fn44oSXP5TrS14C900jIflbxhbL1KA9WDqFmn3U23O8GoihZIGgEc
IvSZkyQaXQ2VttXhDK02R7uIy4qyl0H5QEl+xw2Z82EYCeie9GxmIcaH6111
Ibmk2jIFCxV7R7LRjsLpgM+LozNe68p8ol4Iqum+7iE4gCWa/MMTz3Pzi+JU
POn+yzw1ZTCHG3wJht9eB+pyU6Rx2RdeupU/mxS6EeGSufzDCr94oj5M02Uz
IXvbtPhvVALO1F1uxp8uUUH2dZyxBMdUBNBITZGm4XYcL7lZEgA3nflWD3vP
5AQ9xmeWSXwb20VnNFjowWDFGYkZL0Dq49GlyjA2C5PwSi9qchQ2qUXe7Icn
Uuu5NDdDNf6Fm/5IL4F5dVPw9c7Cc0CTNa88iZXzzSnyiJHe5CaQaLJREFYX
CvrGURGFUrJzCJ2HBCre4S3PcJeubKvfkOwXj3q4U8wGlHnfkaO4OAN62jC+
oBA9sm654D4/wwYZxvKbsbrMpQ2tCoKEitwuifeNfvNWfR9K5z3ct918PB5n
A/XZTzFoTfQvegZk8dNjVR8X+ZdtJQMg4cRgfOZ8yc5aoW++0wDy9d9usdfQ
0sLaKMRFnyxRXjEDAWsDXAWeTONNQznZifRp6muOl7cBCoACqQ5l0Gp5O4wP
Gz91Cy4gThCQzdxuRRV45p1WTofcZC3tHR2elfrvCwRWZGmgCu6IcnJSrq+h
/Xqgqtc9xsAYRs4JXvHLyIT11C0WWWIs1Rof5Ts+So8GrdtssDdfE4HqQQhd
FzXCj1KA0t31cPqqQXxc9k6sT9ve3turqBhfO1pgsBmfBNU49xPZnVHTjSjD
EgjfurF8TXHk6vdMQwpLRNCchs1zm37BQwk9//cTgIhfq8x6639En9KytYVQ
+lMGt0/ooXHPwt5vlIg8DTXbaDjobORD9IYNelfV4IqYPzc253O3lH63u+Uf
ar0IDdIUSc6y68hak66+XNvfIRShvVVFevXvw7fn9pCC7BK5eOSo4W75FVs1
7yegWFdzvm7+xlWG4U6VtpzauoTmZ8FTOtFXqCE3ZXOKadXHxGGH08nYWtCp
LkAYh8habMMdDyNv+OCnS2hgaIeLA71VBfxgXbGJCnKOfUUE4mYppn8Trgc2
WddYFUtiRFsFJsPVprsu77e14la8EVTvJ0cdExP0WVoWnEBkpnt0dd3E7xbt
lWjE0nLKxYNGlVK/YUMhh9YCSSaXZvyeVm8XwaQJunR0RwtJVIpJiDW59r9a
HaVxIsXRPIenFYUIG3z38twlwxXE330m9EDnLBr9/eBp0GaFD/7FHpKm10xW
3gyc4IYY4eA2peek+hj5o+NQmwVJFyAUo8Oo5uEgtfMx3N8s1RyVLXX5fOF9
S59+xk0a4tFI4oZM22xFBISdjqk/m2gc46OmN3DYQMrdBZplnZgyJ04volgm
hHwtwBgoM5bMmVt12f5PMYRTg1+tw09nft7Z78+M0oQjBQIDxVycAHH6fF7s
H/G5TsuNQh0ZG6ZMNjlKTRH0mkwPYMkr64NsFo6ndOz0jzefn8xeeM3UO3JG
zq2741L5gMQeD+FEOUNtGHl8bhgzKfjl7ezMWAk5u+tuX+bDHm4Vxlmd4U4k
EVlnA+paGdFyIKWgyFQKVliSRLpNiATapZt997dhA1TkVpfxZOEadcZnEneh
4Qs+W/86vfCxc8+s5DXKkUDyeAG+bCdR7bvglMi7Ki98JU73+Q4ROiFciOz4
3ZhGaciBdTPxDEkdmfDiCvhhEIoqNYzEx1JhlRWlvTUK9fYEvO97VT73IuCu
7pod4ZRHWgisB5TZUoNUa6BzLotcIs3of9WJKGFSfAtaAnuE5jYAR9iEVt/9
WJ8xI6THzOGbv0AUj8GbpEpatUFRHhR9552u/yNidyOnqQamh3uIlQ9ORKzV
QSO/Fc4gu62gcN2zrqvF+4jydD0RbfK2C13mFkViIvKMtLeSptaMZbH5MC1J
nDcht4vYBAd7WkRHjOoTRjVXlJeDhCEUxHfX/WNetO/ZbKYf174TQAkCg09F
UySKdP2k/9eyClmsKF4y9c6ZoQmlYbk7v+EhK6WCK6FRU4o9CD3b65vd11Lt
gFun7O53+kiQjNEK7hXM2RbxXWPJF3nKNPJJHgVFdCdUmq+767yBXCKFRR9U
2I7/M7Y4fHwAZpKyHpgGDwox3uXklBWwH8VWk4jrN7PeEV6aF0onILgTlkcU
ETAdema1i4vNVAvgAT3vOiz8IROENt7sCQuuSzhGkZu5jZHCiBvWP/clKYo7
YAleWBAc5Uw1YFQnhizxJJpLZkaNZJfKbg7jSoyYN8d+RTpYG3DwTzDUFqyX
Mp0uNrh10fxj8lAsOn1h/lBMmtJHw9K9IjaywUFltiUr6zV4NJArt7t+5Wi0
I+YA4ZHoMEyKdpTsX//NOxRx76AoH/ep28X2DgeYkR1/AX2XRFzt/gRgIJJS
wNe/TgG+9iETYu3lFUy03jibq05botzgJEFwSjylI73IOTONUZP/O5JdfdN+
4UyeEKIB3DHI8F7tJQdP8hrGHwL+dpbqlxjJtVJNCOp5TjZppRJYEMWhiQS0
i/chhONNuIzkaH/vjFFfrLGhB73bbf1lsMParaNOX6rKBcRGmiiDjTnqNVwk
O4WakVY2daR9+fwp2mxGzJGJARfTwhv0AeWo0dfjw4v+0CHOIQmUfDaszuF6
55NbmvXhAE07tuMRtqnAwvw7v2wuXY4xXN6BY4p4IOrSszJXwgx6N5d6mJhS
xayHemRo7EOvueOS3SWpN25rC0lJodmesWYIzx8SQtlI7WpS/MNRwgPWQefA
f8PhJZcf5Qcyh5zuKZRgyEDeBk0CUqf4v1AvjvqmExzlVMOMqKE6eam89sX9
3r+706yXjCkwe0rVzGjLlTZA2g8QKAK35+XzTkZIKAJm8C6tGPMHNn0A5PQ4
AWZmErx/lhnnRs01WTA9DemyyrHGQXs6G1BKErESkujCng+yoLnpRPJ0V0Xc
Txe/12cogFRxtCAdcq6KWrVyYSq/uqie42oJ9fe3QX1WlFh9JvMpbUlBwyCw
HAEqdgCkUVbwcEE68nymJoqtKhFKka8KXCheVs1VHBp5wiYI+GsGXD5LwBHQ
xO/BTV4+ufj9EqZVh468i/v00MmFrUbkZ8upW/aLqQdLvfdP2bhUZkSUb8yK
y6p/tnsLHPT9tpyzvfEON35Thr/JF6JeNlCgqR+PTXVjVZXQl1/THXmkoeqQ
nKH72mLV0rK93gcWuUtJmGOcrv3Qz54mFHVwdQs/u55i9grAhTkagkjYubhK
CIX05riMzTpjc8ZPHErjbshMmBMlrcwsBeiqpyBrnRG+I4W0T3xhCmS1iGDy
7EM3xw/yj/bISbNMiu1GttkP/SmWFQVgbmpMbgjR5yoCQXqmcs/nDGH1hcZ1
owREC3bSeoXS+K8M+fQ//DQs5vU7Ao95/f2eKoGR5Dq9lOXoHOW+BC1oVj7k
SyUkgl3gD+phNmemIrZt5SYEClZWTyoPEHEXTKYLu4XbLHLkAa8IK05rTln1
oNBSwA7dyUwMTUURRJ151kcaCm0TudOA4AiOwlRstxdbpTUMLR5MSbCKMhbY
SgFIuxyDjUIkItQga2p60Sx4aB0BfDLkBvrApQPYY/wJCpDuWG4GnRBjtzaB
RLI/KVmB1Z5xUJRu0tiEeOwdkOXkm37u5OlpkEzMLaQ/I4R8x3rktYz0T8EQ
t8k7M8mR0SECFalcnSrBDO/XALjCI82EDpapGTUTj5Oz2DgqrhKfAQdz3+hy
eFkCkgjW9PTTtjB2uJvSfnSP31l34MkdmhoWuOYFJHc6Etg/CkQJYfsfwwXu
6XvgAF36izgyIE8kSTVkKgq/TfbuDmAwL/lmhGu4meluQUnPVJ2sgG/VcRq8
YYQhaqdwbr4maSgjvAN3eeDDrUL+t+z/2yZA1887kOpJZtVoZiiDmdLHsJKt
vHpIRNl/4cyRTDZQ61eWsvdOQ+xgPTu74t0ZxVgWDTDSEbf3eNKngsTbeLmL
Vpn9kqQC179UdtIsS5r8A1zGMw+drLRs05L/DHzpJ2gRjXWVzBd5iV2Xkkgl
SmT91Tve7lvj2uSz3CELShTH6EpzASALMUVCUrtAzYk5D6MqNoMSqgePl52F
uOOblhzuONNwPa/iAevegiyfW+M64PBKk4VeBkkNezGhO006UzciNkhzOnek
UHb2NuaxM5p1YVN9EqmC6FQUUZCaFr7LJ4GI5g0+pZbr57CPj5VhDsN5CB2x
sYEbfq0BukrBF6+j16NULyGeuQ6vnskw+nC96w0KDVF2Gr3vbRClsR1d80eE
Xp7c003X0JI4n+t7gbWJtRVJVEHjUKZHJLPnzsq2Gac0cTiQQBxzgiEAliUW
TDh1gmq+9NHDzfDWcHZDjIkWjQo5Gh+MYefKEPxNUHOVA4byo2MrIL24KFgd
OyukBmgP+SDYBiWjh0rjIVWFI9PZGfdpAvLtOsp83EEjhI7e7cFigckCkvIV
6wgCjEHtxLMe5DZZ58k8qCGR1KrZ1npR1m/HjVuE0DrGH43AXRkHSrY7zvqv
adTcXXAFAHDfxA25fQ1I+jjom/Xhro3zolhaGG8VDOh5CDc8vaA2/KsAZ5fQ
wjwYVw3WuZq8XEzcZ8Sq7mfAipUSnjZzEeHHzNjDohtsrAqxFHABQr3PA4bK
URaVWmu62SjlgY2jU5u+RezLN8b5d5mS2hzdiuT8NCp2/WYOURuiAD174/RD
W6sEMoXWYQSYB8oRiTQNbvIg4H9pWiDt/8JssMRZPNIyOSyuB2sN/BLZ+gkm
D8QELjjpssUZhuE8ixek9XNQ5bRPvoj7JsRC9iEYX/wRUos2mAhMrUSHEZtw
eA1lEpWLSWG6JjXCfDpHO938XIObYx2VxwEWbwcIkNST2LjbWJ4wyLTYdweE
Kp+Ii96l51s7QS/ZnE+A7Xiaqho1enAcAd37fRDrvBshtI7c4JqKDagkp+i0
dsheM4juA66J6ZtKIG7n1PdK00oqWoVwuuBCatnlluyHjzQdRlf+NFPPCRlx
CXdRbFpIPOy2mQEZJIWGF3LY89lIdR170xlIG2+28irW33YPrwBpgqrGRCiv
by4Yy2ETI4Jarp+wfpVJv1otmwuQMtdjMXUXnlGHDXyxeaNa+tWk9M4U+wEk
oz6vTULDfJzLAIrNjJ9+6WPiBNw7IJ9tTIxH8uxqeNQZkP7k9Xb+Mg/xiRe7
3n2z7rp3m1DLHD3MpLX2lvJXly/UQ3zFRHSauARo+OyM6ZqH/9GJ4R1MqWtb
4D40bOK+ReTjfnZPXYxSoDVETmu/iP2am9presR3YgDd2FHBhI7dZQWxss7a
PiuZYjqIODOPuBKfQ4xVJBYMhOs7qrdXzRwULlIQRBWthPl9XVTtk3yzucIc
ovCyuSwWtN7GcaupcLbeJCpttfFgAhwz+pslk8dQmTdoNi8Uu9xauF/g1W3o
BJczIPTIIrcveQD1SCPpw/jBSqidLnbk+rThVg7G5CZ7uCXK0PvhbCelTE9/
7QniP9rgc6NHRwEv79jeuGyUqjq5W4+Fk5y0c/MH3F06Ga2H+RO+t5EzBmST
SrZ3Fp+TyOJt3msJVBFWO/lTrMSm1UJt+DzJv46+BaTuBkCfL6Uwde2L84/y
V+rZ6KcMuby9lgtmKsKI5MU972XKdtXSp5prSHscCU0v9kjfuSarTNWqy7z1
gDF9nXRIypIWhvARH1ZUR1kdboqCMw1pGwWR/MSyT9gWC5lLlfjGzDIxvSHR
Vwe9Hj0Z2GXW6Ldb8Qce/8D4oIt791sLE7CJQ9RG5/DxzeBVJOWK5KB5BBaW
RzMJGu/euJjrK0zSKMB2x9oIysb71IceX4zk1c+oQbM+zSIl9gVNg/78JNWy
1A+eFiIOo4hlnyDeNI7VwkTpwxnPS3VSSoGPX/8sjeRTxRz671jorqOBZJUH
B2bgdvf/HOK3CDZL48c6FM/RQaoqpTpNLavS/y16QDtaYNJ8LRn62UXsaYPr
e7rRUPR+qP817Xym+5iPJBj5Oq7IKjkwQnbzEO4Pw4H1/JVzaoNdgpy2fAfa
Hpq3tfRrJJkz1MUnqyiUV33bK7B8UTJXcnpMKKS9uGn/k68Wqveq+5uG9eNn
B0hZFCLvv0zpxU6P5wWSlsIB4EaLwpih3zXSCcaphcwSkIxRIXg2mdGgey1F
fU67CxaD0bszMpyO5F756rzXV6QjKMkNyq1ZV3CIe6WOaSbFpmvkkmp7e1Eg
r3icE3p6I7OtfrVS1RIp3+utIlAU80tw5FvqF4KaryclupjQ4fh8kKcyZCTp
35JAUMVE9ss5IGiXB5XyjfoiA6tU3vwTErnmpy3bYjJtrrhFvnlt9JBeKQBD
MHHdmBvrKOsg8XA86Eu1f37axNvrsmsgus1+DoK6w/8YNFRpn8k7NEfoErSO
9MEPoCZzaAP0i1fpgRYFLsIaXqawUcXp/dmnm2/8uovPeApb0evqOMrgeSiT
kbKUSB9/38Si4U1I0NYSc1uoqS+6XvhBjBpi2KpXLjWir2qhvDD6qDFaNQP+
KxsDsAXFrWtnl3TmeClHK/UZMJQnzF54/c3dBrtVWbmMshiVQKSzbCGWv8f7
4Syd27VQCwY/6s6mExuMbjUH3+KCmTe1/yZeDJfRYjIl8cFVTvytvvPeoomp
bjHEGN9KWl7kTKpXYl3w8h3ztkXvfZk/pUWsvf3+y8ndoS1jp71E2jM0HcV8
cca60uZ4APTcQQzpPgiGF7zfmip0/BhRf/z+TusKAMMC1rwsCerjvpWJezV3
bYv5wkn98TKubhi1wnAthxuwzLbUNg9pfbWcIldW31E7eJcREa/KW5j4kMuf
7W2SXAVeUNQg6PUaNkty1k0K4KQOHmmYls32QC+wbQWOOR1KxYcpRbV4wKdk
K1txrY9AQtNAIq/uE466yaexJUwe1fT8tyqjKfGU8S793e+ybtWDTRTx7AFG
A97Rp5qFcozP2zzdgrIubYI3pE3vHQAIjCA8VjFcop7/lmges/zW6WaoBtu0
er3AALNpSKqXHZvj9xYEel+vByV1uM1zPEFc1hr+PEy5erQCf+uBRSXO88Ay
RmRQwL0vPsHP8w+rHNiDX7qdHh1A8Sk2/o+RF8KZ2icveNDdthjXeRfxw9MW
WPTRTkDiQT66zwKRRt0+iwXGj/YifPV+WINspRomGzs8/QWyVRxT3SK4iJpO
0rdHqnm6Pw/AtpjUOhbGexuJq94ON85XGD8Z//Cz59yVOl4C56goWbAxitqj
Tfesy0GCXYIdo0QN00oU0ICbf8Bv8DWWhNF18rexAOKcXlL+amki8/rIHQjl
sXM8gWmOvnVkYjHHTZx0KEvmbcBKeWt4jIrHAPXkWLGTDZU32BXBdmB9xI5a
UbWi3DKyTrW2nh5u6Vfzu/ce9Tsd5edzHHXTPGA8cOAhQF7B5ilUmmztgm1s
L89K2r8TRYrzn+R3qe3mtn25Nf25sFlucsDyOKgGbzNpbyupEtBm4CBm5YZk
a24rAPNt3AXwOro0ErTYZfdh8hSbaQX0rkJnI1Au6eInrYilr+eEMrFHj76D
hULIDeI74cp5W9HK9fmNVOfbmi7P+CzX5H0xCktmRhIRS736u1H6gtLopyI2
MfjmJcfIfa4cNPA+oehLl3eTVYCIjgipvsBdm9LKAFYsCKDSa6gtLlMRrP0K
9ZkePxqVr1olFKpfqO2zK+tnvgBKXXd4Ou+1j7eNwYK6GvI9Z+lVvqm8wjoo
w8j1Hy8wPDdZK3trmx69lCvg+mf7XK48QZJUg/5xvEFCyz9ITUuw+/AD69fC
y6i3K1A0aK69oSqHiSGQ8sHl1pDf0GZuRfeGsfBpkpiSYnanvUWPoef5ptt4
2AMUMktOPwaZDCNYdp/NH4YwVM8fIGpahM12jvtTBnQvsCtqxX2+DcTFqG5X
ICmCsNKYt4/GIpMOr6+5aXjwh6OxMmhRmefRKB97Llp7prJl4ZwJP6b8ukcm
g5iPcxyC4dh+OIguTnS4ai7Wx0fvHoHuI7gm4hKOT02QnqDKQDnA8PZ3rFEF
tK8NnHX7WerDwLDROfyrfFO/PhW5U8wBlgQNolqLZFYzgB0xFK+UkdYHx2nb
v2B/SWK23NDlvMdWchGmNU3bluuo2FtuWlw+RsQwhtp/IhdXrQA5VBuwBrWe
Jjck7jfL/mIh2u8DepEmcrcjxOxNvbkcCTyL4ZcadncZSJ9S/VKW5bPFNec4
Wiy08tGIUaFjymD6F0pA/dDpXklMvrUSE8FVeDxfqEBoqMfKl7mCkPD7sV+7
9fFbp7zcPwQJx3lYIsbUWJDsMALCKCX1qWaGYs9LWfahGc4cU2u3cwbzlVTv
Eg53PnXWpvtfoZkvAmHepGP19H2RsYLCEfdXZhEeN+NQbCic4oSuLoRwIc/f
VYVJciM26911xjGehrhneDWenH2AVhtsrGtzheEONYRYOHn6fyTJPnQYCzxY
zO9aAjUAgqwimIt2ctJUhLqldLcHAVf3p9SRWjasdoWjwE5otL7m1QLlYKUZ
a7PjELi3rEbEzxrZgxVtuTL0FaFpaRfUnVdwbgP6/gQM1f5wAWDT5ahUpOJS
iqoGfRv+XxFH/Btlb4j05W0+ufEPHC00lWMYwnBXOTyK7JJFSLRen2S0qlgJ
V+AwCW6HK//yLQiuFYZyVQeCUwRzQC6CPpsCfmI9RuGqKZDYFc9f0DifBzox
OJE/MGsPkuyQwXYPzIeUG5rO3tCUBFDCRYFJjDAMwOldRqL+taNX8r0o1FE8
SmD+q2ZKzYOnRyNHBqQfisOu+GefZw1h08fb0Ica2ZWGHExmECkUXSVAdFgR
hh+ugs43Ds9QPHHDzrA+g17SvWWacSXTBocmzyI5BDZm3A9GBxh54xZfzip/
dz3BtBOZRHwmv3dPBnZma+wpPdXO1k5hDR+G+9TXLggkp9pFzfBrRtK1yJS1
aULW9+QubXrA9vvQTJZ6uRHRTcikqRCINDqSyzvPGQTGzmQnoY+pB0yQyXup
VRvsPZyhgeylEErJopy/qugSgpms2Q7Wg3MeLkzs1L/mThYVOMVrZZWUtpFU
997CuyahHNTrPOfxjnrZ0NyLwCsMH5oe84px4BY2ObzNrpH3E/S5upoqheAi
0ASkC8Zj9st591b3mxsmIfzFby4pHrj1g2KgLA/uPno7KN3vVaojTaKrtChi
e32w7t8b5sJR6EumQod8M9thZyi3SD+lyhiFjjIlvM1sPiw2j2gm7s2QRLhJ
IKdcyGiZ2nUdNtCzZLF+t89qqk7SzjBeO9NWIPXZ7uBsxWnET7ZNlmNdWMCe
jVh399Low3Cq+ftlzla5S9OFRu53ewEbHzH3SmK2Iil5/kB0S5luzijjTr5V
gCz+sIYLnha4bf8uewEeuUNaId3VKYsTQvMSfM0lZ7tZM4LuZqfyLKnKUpUW
wge0drbw3oQ07pFKbw7j4cS+zSTDrWBGcfDupetaG3QraieI8vokLQoraOd+
FUPvCgZHw29FSxSS1LcEy42+c5iMaNB2td3DN3Yp157lOAfHQT8Sg1m7cO/l
YCML/cd4hzVYKSA2HEZwrf4oKKgaEktHAORxD7nnwMK4oqaqnhWsIqgeI5eF
cTTZ8ZCU+ymUueLuFk63YFpuOp50fs/eMDcuI+8wOm1CPeTEjrtlSg+ifT+7
29Y4t8oizg+krNIbWl7beCZpXdqOSNIJD7AFyftsnlRJ7mSHrlAj/Zd0ouHx
aZCWxWz8tuMnSrAryv2sn31OMHwAKFm0CgOWIoVXFJ38R992Z+jTQODNeK0z
Mhu3D+2AFZXi7tXDr3mFEqgCsWcgGm/mCloxF8b9qBMtfcarDOThsTUPmq+2
wOhX+Gl1DtVFKZaKJz4AEQo+K5irKSiriDJEOkiRxRV9Z0osTQHIVa3/WSIU
0fCHvKCBa10x/WUg2X5NqxPWHWFfEbJq1NgfeMpdr/qXWkE1tb/THbYtLuui
taEz4nTjLAaM9rUOPgbXXO7CLWRZwcC7MqFiTOmv4FtpZKxNWl+lNs9ClEYi
ObeSnoY3oUjWuOoxTJ7IidOYbtr8kK/twULJnKGzHzvVOqE0NV8XElLxMUye
+5j1+Lxap+T3ewrPEJaizxFQYGJXi993nX7Rt/0QTcUGpxspWVoCYoUfcCy/
VPnU4Rq/M0M0WdGCvge4s5srZu2TuZDEaoNFDgUVyTrNw1wcIOzzDbxuaqH5
0eEgzjgLlc5ZWCn8u9+/AQ4YKMuseZxGfYSwBmhQC63AZRRyF9s0HN+YrTkJ
ohv5d55bi8gfS4KgxmBvHTyUS4XLYK9tZRR1O7nADJoHSju7OsqFS0HbXJsp
orbwLujVgwUoQ4VUv9SzigT/w1M/taKd7wzGMhRhWKlmPKq30DmSgQovI4x8
tOz2TfrBf2xzTh7RsD71prlGfCdqUvnaDObaRWlyi/oWBJIjOxextRAGw0dX
Xj4k3T9Hx6giL8XwtRPTpCUeTlcLWOMwQ5ZijxxFVremjWmlg2cOfPFHlcAM
ipu7ID1d94CVyWdIrqIS2wQ2tAC8DNa8730XLWhNy870SHiRkQRqkFSmk4ou
/xEBRgc1RY8pwBUn4aLEj+L4ETXGdK8YYeWFL9zc6U5vQppFmR4lH0eLk4bh
g2Fo0ckwCGLKEySkWrDiq36KCN5t9fZgB6WIcjuLr/qEbo9nK2TX5fhKwi/m
VbOCI9/pqkWQ/GOwWApzG7WHH+luKhBGKE6prv3ltpNF4vUZYYwG2HtzHbtp
8jRcO6nmmnqL03Az/ut/sXCoqzCW3Iw88IjrENMreOVRRcWTn8pGH1s564Fx
GXQDpI3t9rockKSxil3UJTjxZKeTNUvG4/ZVjmW1wE4z6NXgnPX4Nh8Eg9Do
Ylv9wAsUbH8CWGT+0RBw529Ljcr+9EOYvQCouNqvtJRx2iSjtqtSoNiE969x
1rw2AoxWrz9m5UX6VHTSQVzzsQM475rZmKx8dzfUBs2E8/67Aey6nOgUl0Sz
s0nS/HrJe3XUErYHkJqnoAbKO63YxlO9XXp/1a21+C9boPJdF8Ffy1lWyMq8
Wh29BDJnG6CJt36BoNJxepaPMNP8goM6g0qijBf9QG8ASTCVE1OkZZbQpM4/
3OSGsBkXrNuc/rHsdMAHcANhYsqI59lOBrhkxQIW1ekf3W5cJfqF97tGzei5
68DTeH+F58wdjiP+Z4jVF31aW1bU25i07MAwe7QdKiBa37AtmgIxs4gBSINz
56V2DGDKijjDF5D6OUysCJ1d/XFOOLKt5hGybR5AWhbDRDb49eGmwxFmja2X
roil2x+XB8JLCmVGhvh5snXbUzOMbkwQgV5zLO1bxIHifFEme2ho5O4IBzYl
tt6X5LJsGlvf4JhAlw4lauRSpFfiUsRoiQG9u3EMg5aw8ICbjb2rvcXswYe5
eSJg1NK9JHZa2UKHeotarmGV/10nWKjB/ZLHlIGwuyH7Lx43nVZEr5Qu8fYp
uc7E9gkYkr08mPQLl59kDBQBbTLYm+in24oXdILXr13Wm4ouOT0t+HpG4u/X
guwiQdYXZsmZqCsqkeAvR4P5jno/asYEOS5EX3KdMb2o47Yhxd6KTYKIdpV8
9fF+rC1H0JcCPBWzK7WFHiW2B/CmOKn/NeWUZ4HNrOO0YjbswWN3a1/nVEdA
A1g4qmUBlHv8POAmTUSsbOWkCdYLacaVDWkjoNuUfYu/Yz5eN5x8WVX2/i+T
+vbGxKf5REZWeVRjVoL9XbMVBGRZH58jERgV8YVHKLz9Q1MYfLuSUIYF8IyH
Hc6LFnW9hcRUxfh5XoyusDEdDV4237T57eG936A8QXMzEBtXVaTpde25OYaG
t2WEbirAqxq2Wga40PJaj5IsSusffuduJu5OeiARxGSDyvgkwh6BIVqbrlaw
ep0UuxKsWb3R4D75CAV99hcy7DhCQvHncUPj6IUi3MV3PruoUOvOLd3zkFN2
zRzHaQ4pLVrUpOfEh1ZyeWaXTsMOJ6YIqiuD1zT4EjH2rLGmQsl5sgZzJ+ll
zmkoXT78gdf4hUm3/eEj8JGMNGk6PcaAi3n92p+gbxZQ8JhH0Z/qFqaGcJR4
OwjIy2xG67v1daOhZENNq8hj4gHw059e0w0Oc4XjrW+dynp7J4/Q5f6knngo
49EQqXC2C3l9BmIRG2ia5fI66Ev3aac2+gBNzslviQ8QPwv/uIWPUAxOcWnA
wZcprNy+w9sn1tn6gRdHqCxGI+Nlmrin1Owh60J3aEku4UJg9xH2kXyluTcG
D3BJmYxi9vUd61MuuBdm/9Bu1wuGXv+tA4oTQ17o/C1GHwv2u4yzu2m7Dilw
73uPxeDVEChAYfNdyH6KNLFXZMyX1UYYOjsr9ofk0KIfi9sOn5FiUiZPET/e
4HY9/rx3ZLQMEQWjlwZ3z0+LtxzMK93Mj08KSDbaPn/ud9jfZZEb4km9lUoi
ZkoBdyEW4nzVaLyNir9XDmZE3fAk/k5LAGcQlf9NkJHJP9s+hG2b3gsjPlgV
BPiXUjEs4YJ2ou2GZxkJ2IpaUjKWvOX655V4OQKUtURw2TYDTm+juK3NQNCN
Fq7T3YByiJZ0CMT/5jBOkvqF/IBSk9EnIs0I5+kvjndeNiBA4oSLzCzky2zu
lACOvkMiAMz5lN9jMMYIury9R7CZCX0Q5ZK5SprSliXWmKyTxjq9TmaV97BX
dDMbB3z0HmQc9tKUE3Yq0i19tReN8pIBrEqeysQiThDwOPD5dEmsf/WtpzlJ
pTaQwW1PTkngGPMo2aUhbL5zxZJo6VtdCCJdUolDtP2+dg/4KAzz8HPU3SUg
a9WZpWDfaSCg1WyNxvDqTtppCY9LALdROlyGiDGR+pW22RRmMi7e/Hqhe5en
eIr6pNKbOBTqzJwFiVGGAuMN7dIX+Tct4OeIbm8W2o7ghxCk7ZQSJw9MvDBv
wlyQlXRrfjzu82l38gHH+7FvAZtNniOuXxQNSe2Q1ZnWh4g+N6t4+nFXrare
5W3p/mkVAWL4S/HOr2bSeWJLHpy2G7ox6DyWe8uArevkiVnSyI0TFRjDLa1F
qnbMMJaEZo7y4CkjIoVymWJvpHvPDxG7+629hoKzEJIAcoshhosONR1+6sly
srIqmgJIMiNPrZNnGzFIcj6wdxuid33whdIha7rzQS12+yz3VV2qPLiWMxbl
C2P5AvYitPDokbCcllp3H0amw/81FfuRuKUN8wopb+6XqBCe+RF3WzFDuhED
dNFTsyHhuebmKebqz+u/b0so2NqDY8GwwujSJXvqBJf3j5GVtifepi0MtUQ/
T9b2jhnGoJIFT43G+yh7bMClZ+dx3AThbBvf+39Iq4ArBcgP2WcsL1PFNP0/
cBBuH9uvxAI+r+aYk/5AM1cUEjXHHu/A5t+Q55PAtVbcZtbUchx1YOFi2VBA
9c/PgNwqORYBn8jDZXS0+nyMesnEXSDunpgVI+PlhARTJt4nBjLEar9rSppN
6IGhqk4QKjkHTQmSnGDlwMrQelBQX17TEbxLjE2I2Tk3gA8DCYr3aLEHV7H/
ug0CaSYXmTzmYnEawt0B59e563DXOBJaRAEmRug70dst0jLqkk9mysVEnP1n
6o001yIsfReuXj/zXnIrfLSUWqSXrCQnPi7fbOWGjZ/1EjW2TYpVp7NoEdnl
n9aicSlL1As2GcdVpE81WWyLiFBbcfLFED7P4ShGbQIKuKFNx8X7Mdz8OVRL
t5uBeIV+ShyMLFq0iYqkKWqil1+E2+09aqD9aC04bTmZO/SLTpn3EGtok3jM
mAmlIoIL/xkvtJCPwyAbRrq+TAb/k4J2AM97aginhAzToTfU2grmm9vCyuVc
z+hziR83pMEnXuDzqNQHMzIIPE2YKyaMnI6ji9Pfv9Cw9DZNajtkSp2vRdsB
WVVlMDGr3hu9sJUR7uDYL27hQVGQ30fh0fQcCk08z0fSbWLBNXM1OHLBvkV7
eTwGEnZNSsv8HR+H1H6UnytFOBMDBJ9DAF9Rhe+kwKCLLxetkhTfqWy3Kz8u
kBVOq3+lm+MTdcsIPIF1E7xSkfLHYmyQjzBCdqWVZVqtyrXWDNziGG/bBLTG
FNcEBVBKzL48/AhMJz/2LkSXm9S+KaOiejNK4jJe7jKQ/3JnuH39aOcnMZcv
arMGnUfk3EIjoWlThfUjHnXxK568CozvxjJ/gkOOPxferXr8ttlBNQJa5lvN
GKWSobp2SmQ8+hETIJpH068PlfVSWCscsxexuX1qkdGuCI1RLtXROWvUhX5j
+8kLlDv1C4EFz9l8m9R7IbL2IAW87vbZB1ZotIrfZD7ndnUXjqjDYFJh2jcU
9fQo4oVrVnAhMLlP9l/U/g/77I04e2rFLI5fFWTpujSRnHvRAC1e5zVRT9Q0
gned1q7CLW6B1D3tAvGxoV9lvUYMRLHCv+uXaYgtKDn/f4bBjFBzv/XKRTIE
Zoar+C3RV+e7VTm5T3xw/MaEtMXW/etzMNUe7Qrsshwc7L0np8oB8WDtDlsU
B0I5EjloeiZR9PFH1jtUxx0fQqvRmBuPSLsFPV3QnIHivH8/apQPoPZZhPNW
4WV+uhAuEgQrdrdu2u+OAb4bFvJKsjC/lP+jajekK/A+VAlAMHV/sep05wpT
Ng7TRTLbGNQ4wldJgzDsYONRdrYIj7o2yteozeje9bkdKbDKKKeDNc5fZY3r
NPyPKXhzI0hktgWcLFc4nWZCJwCk/itKzklJRZvepEYPR6EYcycUEPSD7+Di
PP+PC2qxvyIjRH0p2dY0nvWiVQNgyxEiSKzG+ECD949JwOJiId1ZcYrxKbjA
8eXDKYDzhdvH9ck4eUs7jGdyLnJlE2uTpSuFAeJTQnfAttNO4cH20F+aHSHN
HQiHYkrarXZqnQkdZjz+Lc+I/UjYuELQTkDxzt63Ptr5OTTNnNThFXOjolWz
V1GD+toCygsaH9L21w2xir+JQn+P6crbKVtjI1t5XTCL4ECZd88Ya5skiajR
jvl1i2s/i4CyLfJXdLZ2tR5KrLWmzBAGK5wop5U7b2qU8snyPMx63+aeYwpP
mix9290o9SDJ2ZgFi09BaZZGgOEPviCWhiq7Nm30pDb+30GZ+t7mg1TF4Ofo
c7oKVH8h9KSxoI3SGQl/OB/cMPbsDIwBySQslXV4H0gkYN9rmIjYAlNVGUYc
N18NRrZwETp7e9CQHL2+lihNjFWHlVXWx+Y8lx2Y+SS5K9OlD78BrT4VkUr0
9L6oqw3OSTJWD9FqHUxB7yAa2bSwmj60SP1QhWxeZOGRbHawDdLCgz9Vy/l1
x+ra8P5tITuSlZopYfc17tmvtJpRyYc8LgKEKSwvjTGpHaVcNiimURJ/vKty
zahDU+puBjlyF6pwSuqI/1BYT2jtE9u1iSA5FKYqn+a1gP542Gb9pLs88Lrb
NgDRxMBckCvP8w9EUj7Zi/V8qQF8noJMQ9a+GKq3O2RrAHgsno1aoLWne/gz
T/BvHZcjNC7myf8GsBfwWY8XvuQk1mycivhL5jtiLetahW7dytK36R+ZhOoo
+X4bC6eZfsAf/qq+6VSxtg75fV+69wdmAge+id+kaSLYSr89iPtcbpRwN6fT
wXt4ZcsJFrpXxWPfA4TYUsXwRcg9IhKOJh34s81X9VVMlmZEasYfMAtg6iah
YQzeWvaK2NdMfvqwbnPzLbsuJbcpVlDiISSObdJ42467r9NFVJLo9L6vOlEC
DoiOYQhPm0M+m3qjv+Ujtpgv9tSuCxHHFRgmS8E8jwcE/iqpRiT7a3inDyo9
xqpBHn0G/F3h0rpqrpc6y2uvU+NAjeDyXzNRdqe9AHylacdf91Nu8CejduC1
wqdOksffZBNQB1BYQOTzCgpbsqgMxpqfDl8s+r72tYT0HAJTDj9wApY4vJg1
drd+Ow3QeQolzedq7KgOlWRL/3cVhYlw2jJ9YxoGI8CzKx3LK46jKfVF/Fkx
tH5rQIFDWOO35fh+MKQ5T7mKuhQreGbxihB7lcwEXZHSPC+XJV+LvMIDxseI
anAqpRYXFf81pn8Cgt031B2yPKBMo55Et9dPj+z8OKL11kxEjmY5OH7QSdTP
GXNybjyUuqFs0fvxbQcEeYMZOcdGWbY9JiybrOX5xUY19/8GUYGCWJe/HMlv
F12FB77MZuX7t6+hkGevz+u9qLBtFvukdxzMVRz3/yMgRRuJy9wjHXJT4C5m
ejdizEyVF2168LUmEMzTzSsqEVfmooJFaxF96kIyw1dbgR8Izw5P35GCD5fe
VPg00DmPpv52mPsV+xmsm9ngY/Hu+n9PTkYDwn2huTo3GSwgWdQPsTva8sYK
2lL8GiXXw+GXXujdn9wyPYNJK4yPmnNsHH0xHBxXCgs/a13FMIahx7tXfyET
uoyv0lopOb7GcsGCFo0lUoGsKehp/uPZx9Mg5YQUl1psihaP5LwKn4zDMCaA
7dvaYECZTBUpvn26DZ1D0w5OiJe8JNqXG7H5b0WCrZqQvHMKphzytPSgioJM
6kaKn6zIYv8So3kdFgWwAv84RpeIGcqoXRQdIY7WQ+EC2E95ZbTAMRslmpch
Kem9y77Jk/NbnPz0fcrdUrYGAklgW22S+DT0h57x7Y2QlE92U8bhFJh7QnzV
7DX+5fcqQPj2dvty/yANghamHGYCx3sQ3pDIq4johaQatGyq13Trdn0YgUVa
OGv1zu96USZn90cdGvXdWRG6J5d+EEv0UBKsS9U5NTVKpyPfXoDee7QAzzHy
9m5MTh06xCKGSZv+PfLK2TVwQcp5676RZuD4k5rWEOaE5xYEuzrxKH40ziUa
fxDCaT1vh6KDlAtdxpcE9/koyrN265wgVIWb7ss3nF0h0DK8iNghoFYIHTg6
DA5p1YZ7fk3Wr9Kpr2RWiQ4wTlTNFEPorusvvAkdFPNROhmjM9ddgpWWU5wF
09C7BMx39MO45TS75zsJim4emR2oAUbd3kCUIYj6S4G5Sp5J6W300pnJlv7Z
ITV7Exx0BMYg6k0/gvRFSQka8LztJcHCq6ttZwJtLreaBCvhbqSk6BZdmICP
RTs86OHu96rquIUfBGSS0yEXkPpeCm3WYxo9MgWLPSI0Cq0rTneCpujbfLzP
PGtC4ok36kLY5B/g2J+pCFszJt3C79wFYscyZYakmP5bUMp5ZvA1hZDePMvl
0eUFtu2ZUsGYuTwSCFdoDbv/S0KjA/apT0bSS4SKU8fFKpIhL4yxwrvOzs+p
IJMSfYi6O34f+9L/xrHw09/WeyA9S9Aqf51LCSoTd2ruKCTvms6IWRJQOanu
guYVFTISi3B5kCVM66CnuNuXX/jWc5tj2K4yxEcU9LJ8ydqLBq9kEbrkk58S
oB0WtgQeyTctTYCCbdYjTIXqJJrnYvUGKrhcXLOKFUpvyB5RfUJPYMzkHok9
xLSmfa+euB5D1XBEa1/YucnT7Q36JQVMcG/zeCRPVUEFBPefE5/2S4I+OQAs
SvD58F2OKUbhzniavpWstmwgk+vQEdSRBbGqhfz/aLnQnmSIt9JtbgQt+zLo
pokT/XpXQJT22/bFxy7678oqlpqBwJy97w+Y/OJPS+Kva+bRxF4VQW5Xf8yg
S9dMWd8qrA5NgmpbM79xyEtWDtBnAlkAh2wcXW4xrpOBia+Ysehx9WpGkQV2
BhxDvCkZ8F3KsRwIVyoQSxUjZL4sfcXAzbfh1gbBOhgqJKgsMiHlrPf1buk8
SjfXjPDW1Z2sZHS5wqCNofe8Ums538bqE7h2EuCHilEwv16DzF32ZgAobWzK
Bhd1wpKw06B7Oql0y1uYP/33R5PeDzrrhn7Q/kADpWHiwhFA0RSRvsw7JhWY
w/uCucGG13bebUv+AlOrhYZsqx2wkgsc74KvkRSLvZcZLSiEcbehBVW4YEjo
08VBrvhsXkAUiKh7lMXhkwvcANi9vYqOs4Hhy7ZVORnF8AsVEuwFk96o9gjh
+JOu9QvWSMwWE98hZk4uADv1M4fEKHvns6Kr1Me5Bjhy03uvbycAzZ11Ukyf
741W20hPTHb97M9E/QASTKeu0A1zUxXI7POl4ckPArQvi45I4G4u/4O60Bf1
N+5ppOkziYp7SgFw6bid0MZgjiz+jRahAGUOXgBKp2uxxidY58vux0ksBZ6u
BZv1kZWynr0MdaokN17wgA0dyipNTp8kqKUWbQI6nkoOUCfBHTs2WY20TYvA
g6SocaW+/YthACMK4gYyoqmScFXEwWLFWrF3U2WkFj/TeQV0lu2MHzINpZjX
mkcKHDlrv6l20jGf25Lx1R67lV12lnE4I6M134l8vO0FIwEi4RMHURTpVPIJ
+C6oqMxaCq4W30IUAKGcts14L+zvdXKPqUyzzbk5zCgRxp1eNqqOqc5fHMzs
nQNuCs2c9nTHjK2LkOQ69jrN34bL+QkNv7mA7zGMSLH+jUdgJ5pibNpOcVBe
vjUZmuA1Gzu7CVoJKF6JL04aNkjDC5CSYalOouyRR7Y9q6fxcy3DoYHMdWLz
ETIyj7rHZRkJS286fBxnR3S5jswTLfV48R7iExHBwpucdaZAijOC32KumxBi
hsS8gyOXiHGV1kAmVr2520vjkbxRhyXryuBef/4PRIj/VDHWr767zskxPAAT
Uzh2THS6PJ8ebKeNRVjKG95eKMuE+yXrgvpDuC63eF9ILJPNp//bLQn+Iow4
QB1hhpnGTs5XIY6cR9yWVvBDZvcNdnk9jP4ntGWZOmfY6FDh+7Zay6uYuzRG
DthaaJWI6PsN0xXQ93OcKLQx0yNqyWV5dIqnpmu0xzUmIx50BmLEsn2gpZcd
Q7kH51q1x/fp837Mws/yKlTZUrNcaOsXvTM4qcrHGy2P8R+IWSFRGDW6BbqM
cTvFNEs3bruOYcSv/va3KqvMNTSVgOCrhwAfpSszGNa/GyeVnDXtk6j/6O7j
3AAllYbkCXehye6jHsLcdafo9NKafugsCbPiGJAWWRLtIDQt/4/mP3BrwVLt
eRx6vFj3yx26GF0rq91iVX4TSqhINn+jM/VbIxNOfP/BIlNXdwrcupS8PKtZ
eCv/tGqCRwZSnfVG5Eh/rUO4PzdrFNHGeGjP/DEYFDTtyhYzrV7LjlLoePOB
GNxiY3UlDdCBeoaxYnXsWlylhq+vlam2u5CsElPXhtUBP++N+Lp757/n+Et2
1H8bbVPaIUP6xQS0DljKUKjfD3N/VZiddCfQVg4kvWob4LkOUOMWB2A4I7Km
s7DRuDv01jeL2yYlc+/aY+UPKbNqVEP86jlkGbfVMjTOXkExFzoanjiQO8TH
U6OA7HnQ6Y5Hcd5kSo3b39g8wwXvGUKRReUOyRa9kUWBRPOd3lsoUbgL/V/H
6sHTQMRUGWPY50icP5xc2/5QDlumCEKuja+Z8nwQbHwV8V6tD2j+bhsLmqge
PANJfoirZ+mY2gFZho88HJeu4OEsWw5OuSvbiwYfNx8lUVZwl5jRkBX5GBnJ
2bsezHFbwbwskSrC3XZHWfqjZo+8KY0OWHtNTHx6K1Bu1KKd8TyXYM8ydPnE
TK89V1QZG+z1j3y3Bhp1T0d99tJeRGMBBChtDXdat/IfMckYGAtdYtzsAWuS
11WMPPDdbaOZ99axpPFVD9ZXFzOF8YOrQebYOcyE6jheclju81MCsgB0HkbX
/4hGECILBWnprCccpBSSQj/qIAivnZIVPW3PFx7K8g3WXoKfxqd7fBZuMMPB
TFe9tModDURSE+wFBcFPgJh69PkABHspyoJLS9Pr/W2A7QdiM3uFXTA9sfsf
f38Rvd5LRaE3ZEiqzyVOUQHruiC0zv6z2+kBm9Sj3EB+nc6dusjqmLjjukrt
wwG6hRsubNyjkdUmleZ7yapf/yA/Xr1b+3ydmg418/oUVn7An82Btxt8HeBA
T0JHZtIlA6DHFIqfg79DYUJ4Lmuk+yfeaA+Xb3M4xoGDrEpbeVumWhNEWk2D
xG4PQwdq+m5XVVprBHlJalZztq1g5QVea8gs+ZtqUj/pCzMv/+NfGV63aE78
Wj8x4W6aRBMbnzk92xCy6gMe+ZJc0xM3Hm1YOhvHH4F5nnnU8VDcnz7cLt7A
8yb1sDghOk7erj3ePcm+TQTQHQ1tk1nw8AS1lx3beKjzRJAms6UxJRGWjtKS
hQUw2W+vTyrYCkqkqnOFW7crb60gIP5OwZTXsmmDvYcu6tXuhoTtahZq4wpm
sTur4dpU00UW7weUsr/vdRMhz5cB0rxvZO9c+Atm3S2JiPZJKHgofvoYCTbx
rKQpa+GKYCY0Fw8aKneb6MiWEaNQKtZ0iOqxSazljbRfhQLTAZfIr8KIz8e6
ChQb6dVankLbVmAa6ZoRrxIwYfSrbzNrFqiNE2+8a1Mo8+xAOE16PPvaAsk6
5PpWPdkKp9brAidv4ziDNjzxnNa1KMsNRaRGpbXx8watrbOINPBoDL0dDxxy
1eKDw1HbG7kxz4OQjCA9KRbNu6gVEF60LkXhSr8iUxh5tRFxKl1jmMFGAEE/
Ny6JA79mxxCjWPWFrWHRu5a36bCpAzT6anfcvPAa8H4w3H7R5qDnV/UsWog9
qHA0UUlKC9fvaL6uO/q9Yqx7s06gEeWLjvbu2Wj0bf1q49cHNd+CWQBec6/V
d1hcmMm3UM/elG0HylGCMBMlYQL+70zJALe+cD39Fy3kLFh3RalxiyxShdRB
3HsKElu7PMh19Yyca8Yym1BkphhTDNryQ2FuM4vpnXIMOlz7O66gOWYbf8ro
6YOblTKD8p2akyiPLLGkfoA0MZHL3F1vBxp8PJ8pi2zmLjInSXxSqxBeTRR5
tkfc7al723Y07HAko/xQJzP5bujUljBgqNF3VsB81/2fkWJIFiI4e6TLT+xg
4oJwCtPnNcH6HMQTLsizgoEt18Br+J5skfCheGj75myAhnOCrTwO7/OschXw
1nctz2akLcmNUs72IrKkwvaG4zZnWB89Q0eY8aU3B872M4dL5QwmneeUCR4M
KccU8gdnwkBNOo+zC0iNvJiHBodraBbTGQuNm0/tDGYfsy5uDObkVQP4faaf
h9H5+Ub8jMQiTvhdDNiG72YtXMAKohR/YIcOwIe/wPbcFtovJxQzU77GbOmX
6c93QTwSyUOPmLYAlJLZ34kq7d8KJVq6JOtGW5VwlIyq9xjRN0mK5byf6tVA
E+HPTEMqIjunlm8+NYn352mnnEfG7SKaVAYO+iIu+d/spone43gIAVyMv40X
pQDp8mJFWOnV0Z4AcfURkqyX89XlVuioSCQSJ2i8UET0BI+zjS0hWeqo3+qP
sqWRGfRIW62ZkKbyN8zAA0nNdCBK7JBDRQsY6TV0V3xgMGxHKNsplZcXYkpA
95w71hydvOpgJA393hyNHMH3JaAl4EpDGlzWXcXvt0BXgNbRXlKBp7Qj7djP
S0/IyLjlK9hxWNr0NGmxwhL7T0yyQkzuSBptKw0srYe2a0Qlujg4sZHo8I8w
dMkpMVMJu83b4dFEl5xlmicHVFySNuU9KarzPo0KbuWSPeEaI3NbSxatIGiP
rl9+pbmvKKDnmMpjFTsNpZ+A+8MYQgW/e5Ucjsmee5h8hjUDfanCHV6W0ly4
q7x0jCajP1q9nOHShnu+FrEVK0nWcEBQsie+SG2EWW2BIxTISPjC/vYVVF9+
lymDTtmQvuddJFE8drh5GMRyrQJGXu6mmvXw1eVq74p5kFvG4oW7yxxAAq3m
szOWpZLZ9KyrB87PVdyqRLmcehpMhlOh+t5ME58aihaYRGla9+BrK50J0B5i
o+E/shZyRe29S50OPf87IDKw30k5eLrzvpQMaeh1yzFaFv3mbrkC0ejfLN0b
tVF7S7hbaJXqzxEu/B9HUvk2IcNhviSVv10SVcB+qeTm5+3etGJnSnLJjn5H
ydK4uX2C9ZBDvWUbFGXJ75WYmBZyDh/mpnGNlt87Z6Cp8gBz7YEsEjy3F4yp
+WT5/KE6+V+tajgymWoj3PxiyARorinel14RPqlyY7hcERAL1pAraEoQ/apv
ulDNdOFKdbz1/lLaS1XFPw4PFLar00nj+1g/7f13tryJNwECTN3osq4jNe5M
8NsWru1z1BDTiAib54ww3m+n43uPvrS9+QWBbbozrTrjUY/mddDRfh703a5p
pIztfAIg2tfHCju7tOPOkAmHX1RYhZoi9mAtjhKmxu719kozdQcklsdHwUua
Zj1FWLO+2MDIYMJpAHTxYAItgF+DgAwA8IKZMicbu3JdgjGWbJDQvHDHXmu4
4Ttzr7yW+r+dKm3RrXKfvPBn2i4/ghoTnT9UG5bFmwS6CPnK0wlk5Yenq8ml
z0WBNd83W4vIfhQ4b7xrXKggJjA31n4gtDsXiKop7IS9nHIKh2dhWhWi1F2S
VtGkpNetHLrELffv6msAWlLKn6WQ28EIr87FqHAZ4/rPpHGQmKelmMy+aLvw
4scBtZERLwdB+5OSx0YzT9lgErITL+snqA==

`pragma protect end_protected
