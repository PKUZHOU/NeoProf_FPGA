// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
V0jffOOMtz2IJ7Bla2z/sIIs/DbINFv8EEIq0NtSSLGe89vKMkXHg6FRb7R9
R2QV6hPM3D9HPfNjJsCaL7RI0m+ugiGNtJTzpo1RJ4YBH6CLP7TSBnahseOf
i//oY3psp7xbKUsyKOHkVqS0Ea/fIatIQWL7oddqCGm2ApfD9cjpgw2M4HhN
zrg1xnNxZjlfiK3epJXh9uHe220ivNJRN5zouaPdZImA8LHJLvzt+CNoskW9
1hX55jMsjhJnseeleoe/jvGKvSDrDumgL2emHZBlEnMSEMYPlmKUT1Z3UBqW
Wy9DuoQ3D9CW0SeNTKxf2mg3i+oqdn/PbnPbc0D0Jw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bxrHRZLZupuZgelkd7qzEifMHx8E2cBpRvF8e8DIlhXR0ktcxw90t3Nl+j5T
djAQ6xMQ+s5lxXCAaPvu/CFF8G0GiqGBAdFLIX7fJSqbTvqX3Xqe5gACCMyh
lijMO1m6t7RviQ7uaHwkhODEhnGK5rmw4wHa2gI5LBgp1dm6Z9rAQQf9xAFK
h+PLqw5qBCk0km9m4XmgHbSHh7px1Ca07L86huKDfcYA3de+Kz3EhNz0y4ds
vzkVVx7RCls9gxebRS/LYVCgldxcoaeXtDgvTtuuEWveQtTmLwl0zlVZlu3a
XjAiQhxWmaCOZJGT5FYvHgjW9DLMxexWkrjQtES96A==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mdju6Zi7DJUMzxdSoSAHiX1XWIl3t8rbLi0i8joTUyrLENvfDn2Tz5qiwX2f
OXIbM3G1lsUAZg2hj8A2UMpyC03Dz0Fqeq6XQe2O+1uaK0SlUvslBVUnpt7y
5xii9uVJhSKQSF3Zj60ob/43OMHq156GaGjrtn2D89dSOLVqnrpuYdveCE9p
qlyqm4LdPLa0V34iE+EclppMr8VQvV1oifyr2FO92eYzM0qchrvTc+PSJGIC
e7xx/agoUGfQ+ofTdSTHzt3p5dCNfzPpUtpCC2HRJ7Bi4FjnQkN7UZieXiG9
C9XYpYOctW3swc0/4agyq3Hn4KrSkKrq7RQYeT1jjw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Yk8meQtS5BXP0vVg/pxRkqQTTjcHkpOGOI11+CSR6gIvEfSBD7Sn/YavF3s6
AXjYlsSgqGdt/XyWy9Bb7VPmw2M8Akr+yN/wWFex9u4xE4ybC4ceoUxFNd72
yDFTQndUevkSyAxfecypsjirl9RR7KA0ZWnGa0m0zPW8ghr0mwE=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
wHgCphZv932kpiIvDEpo1BEcqaXlHVsRpWhL7cZXN3ezTUP61Jpr+2B8vi5e
r61RkKuyDgYYUxjqg+wjtYyyoOYnQZLmzF72F6THfOAaEvsnj8ft9+b9MAs5
DOqIxHep+JiaLtCdpQ5e1vTnohBQsUJXPg+PA/KE5B59jgYFIbqmigUTwhqM
GG1kkorXch3KI2R8S/X2YhUfF1PcbFJm/Rs7qJ1hs0EJ40GTDX+oe0Bpae9x
3w8137i81M1tpaaJEnFBaqZH3Zs/Fg/H+CACnCx7rHODXojYlCM7xhoGEhtL
8NwNqtb5BigDXAU+s91BHRPGRLgm+KOYhCTXY04ubSWElDydPPANpvyUOdj7
2iXCoEumpwsjGqTG517PFBQJ6WUc2XU4FWVvoIXd1Ts0X0GL2wtj1zUMTnpx
KUtTYvT4kvkRdvA/9xoSiM61pjfS5RGVAT9WYs5p9DNdVHHFKUX5PFnzAlYL
KYTJc+YbNjueTW0gdqlBxB9jVdwW31RB


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
BJ47ij4QL3Tq3yjzTrQyNuSiW2EqfvXxEIu5Br8hu9BXC6q0p7KEYcDG5Ukm
DgCUYwL8+eXAekBHDSSb5KQH6IstQLO0HlGAQ0VefRskTIfxLKDJp8u/WmAv
/pFQFWwbT/NMnq+ps8d8MjGec+979Re7fOS4QnbO5VwwIZgbwck=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
G2sNY+5sUuW7YWbDlK8+/nX1OWxJtBqYrTSjGJeyUoZgu4ZOi5KqqQS07iuw
oYdr7gluWzustNQvsaLAJn/ZfO6kmpBrtuiCk/rZia4saD+v7z0c/h6MXomZ
MsEaw+rvGOXyDKkCS7p9NkqPE0w87rgU3J6liINDEpllJI5KaFs=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 104096)
`pragma protect data_block
O9WBdQVIfY3H+ujXumKgrkwubWDDv2+pCq83SIu1ChVW9VrCXuLGMWk687B+
Uxs6phNm7KQN+7Dddctd5Ffo5w3TcgNCkiw/rpK6UYaoWBSOOBQY6fy2XAdU
Kgi7yN4XKZQeLNtYKUA0zBLCF14Dc3W56j9VMzRohrbnX+fb0MrvbVRF40wC
ykVPfWl25mPqws5Pt0c3sLElknGJ2ES2+TJrfFR8iXjfql8tGUoF99bTyUwL
mAcOVH9p3HazSnVzxXhNz7cn5HByZ4YBUsdL12dlSzeqI0UD97Ftts4bS/G9
LfQV0A5f9/TdxLrQWUnDpr3VdrBaiwMvX23IGRCaHV5ls4bZGLP7h3+UgBdI
+tCqtRVlmSOjQUAxWEQ6lKJFdFb3/ZWn0vhO7wHHeyYPurATi34R9T3+abWc
1QXGotPTERUzeYgtWABn3ipSth5DsADRB3npoLy6K201OzdPI7Gtf04KVmEB
OI2muQX9KtZ9uzetwHiqoxZAopLHmCscGzvaeNloGB/G3oUSAka3RtG5nDw0
1/DT19d6i6Kz6Qj1k09fq3xdDkVxM4th4Q1xENH5gkz65y00axM51WWY6H72
1TN0fjnGyFoDyfIji3cbRaWSKj1D5MmKtoZu3pcAd3aAPweXVTdtTDZ5jiHv
/YYhKdHE2ZkZYmerPaSpr8mKFcW+1FyT4TxtNiReqShDaSAeu7vbb0yLhZyA
30jikidtBTJUHXx0dtzHcjqnmtvYhdlKUcqxvAQIHKa2pBFJYa0qAgZAg1Fa
SfuExZiL512tqJPZEDNYh48bwXQ358ICWcd9kFozyyEoAhQgkAJCeAemUOHB
K6VpaQoXNrVchs4I6zz6tmfdPyvT3bTOPNr51CQuJi2Za+suzO1nD1xbzSmv
bDK3BSRLfeiCjyLnWKNEI0ErzIs7Rat447e+h+0zW1Aw4v+lFfErxGGcQdr5
pTmxDBVPAnhrk4h92mQEFeE5e/wbcdvQdRJR4vi1w9/2BxKXU+saida/DVZQ
sMdhh4gIHi3REM1OS/pK3bV9zYI3BvW0XXRTp1S2m7bLR3EEexyoP+Ff8CSZ
pZK8PA/l2HvZZZoY0GcOe1lnhNYZTBnB61JtHpD1ah2yNX5O23gcN9xraT0C
uXcOdPetK6Bo4i82hrhw8j8fGTH5gv2zMk/NfomFYKURmN5Yli8qfwch9WfX
GXuvrnbHp2ke+gd12gP29FAWtsB5jb9r1deSUqjQ+/xS6oQ4evQe2dnS2Z9F
YxtYaq4frU9WijJfDnHXGsloYmmIf+jWCGjAAgMgCSv52N9t/00khPhzz8ih
+ZAZpWIxxDkiSxs2bZL/5iOYJNisqARqknw47opMY2X7Ab4Rf/lw9Q7U5RKP
aNSst0TW6RLrODYbRFkh4X08y4X7gEZoTSzurw/tJ8+e71LAjQugiUf0vGZf
g0d6EuznjINXwwWcMF5hF7ukGd2JZ/isO7pD/rHu+mVi4PDyq3NyRiBirMpt
69twirXC7M/ku+mIgOdAl9kPl221swqZrLDJamWk78BBUpJMpqw5GrJ65CpZ
oiMz5TMVxMIbw55SA61qmEUGnuWSX/cWyEIgfRlOKOwBr9NMxU6rLEiSa1eJ
8xYbgwX5bpoKT2beXzSYp9Y0lD1jFzNND3zdnyQCGPPKLNazqmi5Lw7y4g8m
CQxiIZIiTCo78KzoLSeqnHxEyLsGv3m+33DdNDVg/r7P/ThVfkF0/aqBIrr3
jXmxYBaD0aJVH9sn6RLoUpRU7zq7Q8Ow0fXE5eJStlMSO96B+SMRT/hGGWaO
vi5PWM8Po39wC2hgycbs/blFrTiaFLGw9vAnJlxyeyiPJuWqFej+fAAEYWC9
xJztdfm9V8s12feXWnTG/rQY1ue9Q9eyP39i9hLHBIt01Awxccd5jZfPxN7r
4b4tq5eTYYkExxC1kB3igEPzxgwtjV3gH1AwUKq70H+S7qEmZmLzZzAnUON3
V8ZdBi1KDK3jfOUf1xSOED7H2th+8gbN5VgzsZNfrd/ZfqLFKpjbFNRRrXde
S2NA5CAm2FOkw0QHn10SXOTkuSHlmySFf3SalqVOR8kx7DlVzxhmhZs+wn/L
oOi2ED35qn/o/xW2KG+kW+gccZER9mycn6To67s47/lB1rILIcGMwrJNnl6Z
5qsbwf4T+LB9dc6RjR+xayssqAPuX+BfyGH7tn6hHunsW20ZQBNsiqlcPIF6
nPvD7hexaAjrhxctSxuqCvNUnWiS7hP2CYcL9Vw/H7AsrK9rz6YOAlO5CNhM
N9pzhM+cjps5M6cum9jwRFTJbuszz6nQHnDOdNbnSCPkxUBHiR5770dIuMG6
9fijVNUmrtxhONwKoi9JG7Cub8w9i+Kjqe5wwvWT/BmP5sw0sktBMpvOQ0ti
nyR92cY2BSyviHR1rVc3Wg6cBSyjQCxPtlzIBeQn9+kQOivET5YTMSEGBF8F
H1uSOyHQk3T90QfONLMUb9jlsPVdw+QCn7yxae3BUVt/LPuwTMpU6WP0Eqh3
OfeUteOKbQXsCDIaIUf0cF1Jpw9TBF2FgQth3xKRwv2EP031HP61GIrElrYe
brJqvUwFLnHblJ7Dl0ywTXOr3s0jicPx4l+BtbaeAvOkj336oqdhjJIp9o2P
8IQZfcO/ZUDnK2/nYwPwXRbX7imwBp5UnxtLsu5virXPagROTGqZnncBsoD7
dbWZDY7guZd/j4fqYZqIBUHLAerz08fzjGfWAFagH9oLYhplt6NsDCvo73/a
4hizhZ1VYxPFZnx2l5yfmEFl5pF5eUFDlSlFkWVApoBPuJv2O3AEC/ZgggPG
FrKhM/vzl3EE8CvRfqOoSA+hIGiGCijJ+iIj4nUsmr4pXpHJypxL/3xTWt7s
KJ8aozLXSeLY8n9yiUegqob3FrXfIpOUq5nwqQs8bAQc+sgcribU3E5PytsY
ZNYLBN/5szlDXhvaXMDp/Qlg7R3T0K3ANoxgxnyxB9HRKjgVdU3ZxglbsNxP
tlYAJ0PUotWP7uRXzMML93xbxBOULhZo6NUVaAdmrt0AWqRD0wBVddtKv9hV
Ypvepjd35cT4dLuav7yt6QgS4agNdWa7uWAYkASfuXtHJZOAeh6UcTMJc0dy
CYYEH//ix+JyqZgbGJ4sJoQ1Ms5HoSilhY+g6bSMCQ6Rt7DOhlyb5RodK2YB
lPHjFZwYvjSxZwxAinGTyOVsJdg3y8Nn3ESEJevyUyCeuVQiuuryRy3cheqa
oBm8aL1FPpTjzW8m17AA86DdMf9oT7beOQWPrDG8GSXyBbpaMSW6xzhxS9En
IdZxk5Bt4AsidlfEXYJ7jkHXDlJSBgkR3RV7oIlpIR6SbW5TYQiiQEp3MASL
11QrfCXQvmgGAUleI2NV5+H3yS0HXqfeTkRmDLNWXzLGmPYEVxeIejluKP/n
0R5oV18S0ONWfZNt5FzCMOfwAGRGr8ZUZmv++xXDbrwbgMxiOK+CQDeulDG6
IvSjAohlXdHUax3Bbsvd+qsaaKR2XPQZgZcF3Uj1FtTYoRDE6NdBwNkYKZGm
QfB8N2E8j+UMtbhTybE/E8DRxPQ4HWTUgI/GA50YGbvURUZ6XoG6TvYeIJkB
JDRaiSjvE6p1MCAvqL+gdNZ0+/JtHOFyURxJLELjGoxBDJua1Eth4lp2isR0
0bqtEKJZYRTRr4Lvekjh163fV1Qp8KbIKAo8JC74JMYww9pdt+PTgZ0w+zJ8
KAdGi1AHxVxKI9hNopv8/6wm172l5kZQ1N2HPlhASaLsGoL54sO1dRiByl1a
WUZkLHvtPTQPqJewWPGUeWb4Ua1V5kdbKBw7wRVFGVTWhVnPBr9hTGfml5Pm
ml64pngbIlIpZa0pGzrqCJ3veHC32reozT29doZ25tYUtUaiPFcw86trWyhN
ObxZ4AT/cKuS1+aRm6uAA5Dk/SC6/jFx9GPMnmr2kbq7PsiZT3oMb+oySBPv
n6jvWyx5tOa/eeFyZOBF3GOkrL9T7s/I1oyonjnrg13AlLCxa29+QMdPTO6P
blCoHQXXczjLUWMeJpujSAPoXxsnYtudcRNaoGq56vDe1++HSrI+yi1BVtkL
FeVfQ+g3bYEy/bqsCdHPVBSyiMMV0ew2YRFH8ijDfG0pVrXZ8Okl/4i7QElO
Z/MKIDIWEYhej1qR7QlOXWlpe67tptgcVUxg4Nu7lWkLYfpAAJN7Et4HN15L
aGt4DxxXLbk9hwI+ovPe9mJTD2tH9E1MNxhwhZINgiL12ki+rTCgJRWEzFcb
QtIa4rnnXu4Hxhg6YHMFa1u60V52J/MFnQ1qCdqc888ygXnsKDwKXIh1QjjX
OzF/pgunPBHKpI/fGf+8VDvn934PFGS+fLCBQZkhqURfeHBloHA3qxfrlDXC
5uzIx8bRmFyZWNsG8ra1kC1yWC/DMqcN8ahO4RQloAqucVZNFiiVtRLKpJLC
5QHz2YsLScAgGjpN2jwzpIMAFysHKvxdQ+dqdbLzdbwkuw2ESTGxvRIrSZgU
Ajx4DE4KeqhbIeW4gJN64DXqBN7giNBuz6+0WEFc4cHuvFLWEFTf5YjhoHPQ
Cq6fHFQ8gTJ4lOEZOr7cB3qW39i49gZQBvS1SGFnmWCh0DicUwp/lrV8rMR+
xDqqSDnCzFbLgJ4YWlmKO+BNU1ggniwdcdlxEzpplGFwbpVdO67r1Rrlzph3
/vXllO+4gukB2+UIM2P5P+2f9COfh9ackThqyls/bP+bXtXnWW2nhs3q+FX9
bUogZN68kR+tWZxGyeTpnak63R5gcoFYqK8J9JKQ1XxC8EZaCpdwDeYNwVaK
5u7NI4R+Jn8494cS9CzVJWscMVpCR5VH5A6SAPUvs4i1ifCmiykTo004K04i
R/drLkLgKt0+QVLikukkt3Ju1o8ymKo+7tyUMw7tYw4UebhslKZ8PhoJtefP
DFG7uT17XcDJC8warhi3IvfQieWNPVlEuE3Fx6TxTmJY9uLPdk4hIPGy2BFH
cDx9LDT3Iw2WOQzSUzwAu+cMRL1iN7Vp3LaWPrHSj9ztvafmu33YJt04LdbN
qIoF6VxaJTQfExxVu2guE7KCqzwxKKBrPBzccsMWUpiWWEvAEoRd/IqhDZlI
gapmftaLFE+XFMEzsFPlP8dpKDXuGPaLssIVN6nmtiwLUG7JyS+vTEmJeoIo
7GRJK15zlS6nnlBxRphpr9b3Iq9EPjY2xc1B3rsqI9BkpghcUcLRhRNiFbbF
KPgo9atbWjs8fU/DK0BW1PzQLn140gT6BUHGkoUF07C74+kWdqf+uuvOG6i+
Th0KUe4esp78dEWSMi4fveqy8+9u6geVNWkdw5BQ5BoRe/kKS8RgyXM+a6CH
IUAwXSxnml8yHwQxVADzFvNk7q2zviXQDsWWhDydzFsoINq/GWn5gLsFXk9w
EPOLsM1Lahgzn5NCFWl2X9zfciBdAbCAgOli7IOqVxy1PoZSlsyhlszIDXn6
eX8KV1w8+mbHt7fMG10akuEuMcz9dzBj/lXO42eEeqweyp7joCVWNx9Ra+E7
5Hk3jYaX8H08I8zBjjJlTj7GSNK5kT1wS6PS+C3iKE/xxgvjaB8Aq9BkpSMj
bmitOiLOIhW/PU7vC+REGZaFF4SMS68OKVPmpZnkr5W1BMXfrcxqqrrj6/T7
1CH43xjB4TAJcjG5s4T76DfzVZZx8zfXDXsRf34tiH0l3kMdCTX10A0uwcNp
VCX5G4DJngkoDUmHahQm9qqbM4HecUev6b5aagGKNtjB4ag98oih4x5ARi+S
NPgeDPdY9cSfq3EziOmAHBGUOsFEG0tsCbZ7qVlnvrQnlPouZPEo9yZCVltq
0wGgMDzeUY9b73HqUGHKChiT11mL5m4h5hkibhoC53FC2qWMB9ShI5Kq49Hv
C3TTdw6GRBltQVAWGrwRrKutxB7uNGo8Cj/m6C1PB29kjF9N+KIxih/xAWEE
BDMS2hh5qq240m16DVz1CRu8xdL7TSemcgHjyA0kD+crf53Z7HjzoacxjHsj
gk5OTxvbp0HRD2HJhBkeKXMWBmbAM+RjFMcTQb92bnEMhb6yq4B88FZZNGIY
Gz7ksMFX8L4dZflrQvjXUXhB+qKePEfaH6J+cyI4XUq1Ll/w7KgcT9RrHDuY
E6T7G+qN+Dzw92SkrrnxbUvXydHD9iU+hQcSQpJB1st08qNP+yR3p8Y3KQtK
37O72NdI3QOOfezfpsLcYo03dLoLzxIo+oB01hbiEEq+7pv4VGWlqUKtVjlH
Y3wPv8/+bNEcQr/8mpD8VtGQNNJI6p/a356cYU/sfpiMdJ+BLJM3Mx2fD1xm
TSUqMHUWhdhZrGVqEjmB/NJ7AqJiWb2atadqePeLd+Mfvn+a96ICmDTHR8lF
LM3m/zbx6A+0XXFVLQVBiNKmtiWijvYJn0AlqlP5bjPlatiFF2rf+QNqRf+d
f6wo9VP034EmeFGVyuw4l05Zf+2M7xP/sDl7+5gtglkyiSN2qhCjtTcExC0b
ELRtNUMxcZDowfgB9rj3qRR/66G8RHBptQLebs4d4SgAt9mSTnyeoH45GW5p
lT/WRJ+ockBtAKOH59Fxd9XcIMwOlNUnCKu0p18Rzsv3TZuGk10k0qINr0B3
gVxRJ+AbpvzIgYKfD+UVF+X2Ce2+c2NHwddSK/rkJd2puzEI3EeWgvX2YyD5
WN9FWljYRngPSi17VFGmuTUC8wLwYAJd3VJitE3OHDNcrQ/7wmDRGOyYY8o6
WzeO+FMv+fcgU8hXQRCG1nueaxguxXmjGvG3VAP8yQLXVNRx0Ox8nQgJI9KX
syEvc6SnhRzkIoGZDYJ/qQFXUbXu+STsEQABViN8tUQEiNUtmOrvL/E/4k/I
p+3pXfa+k9P3ZPt/vgjtJwHzCPXoEC8+0fChThS2ve2+SbQIAWinlH43+fQN
+TBMUVicOwINCbtNbVFhtlXGqDSZcpJyxvpc4RKojAIjQ6gzVDEmUZi5imX3
W9pxE752YDvLniwNOJFaDGgCD8hgDW7a+TrqmvsL2nbObEb+JK/ANeoyXnnT
QCWqNF9ghtSbQFFw0wi5t1AvoVb/2Zgm7lS8xc0TsIVru8ehhG4CxEmE++ls
tfw6cjB3uLIoBpBTba4m+r9e94/vxHNCGJa1nRSY5n5l7LRSCKDwczkwTLVM
8wYjBed/e51dtxFnaLc+Hjwywxvr/ifYiqnumpCtGzBG+cc/HC0Tqm+eO79o
2uhkJGdtvullyqwGj3r3FFzHNR1aicTlyE4n/RqaPokimxMEZBqFdQuTKylV
Vw5KCoEv1bgMW0bS63gttNh0aOmhh0ihY3HhhKOac07vcmONqeG8ApoYw+BO
YOEDkDM1iiqWr6mlv0ZtZEAz42tiJMcAlBrOhF1AlkU9Zj6TIEod5DSV5mIW
kabwLjQyMpbxyyYgcY7dAK6yaMRYHkHR16NTcySegJIz6bI1PZMslD7wn9Or
W2ivk9/WdVwhyZaC688+gGtxfJXH0+q1/lmBY+/QNf5sctjn2wJ9nbJx55zZ
O4sla7V6LjdgYlbT7VS3XoFVacKTnm7UXBftWsKz9PZcOgbtJvisfEES8T5F
g7sCjYZD04LncZbzw4yrZ5hVwn3NAH60aJInUIeJAhhaWn2aeFsthVehjGlB
1mc8JGYlb9eqP1BXKgmc9n/M+/iV68BmgC40KHEftSPlvdgQW4y/tbEspquy
xViwlvHiD98OvRNAVds1Rf+R4srI1R6tQ5ZkuIbpgKEzjQQf7RLkWYcn13rO
8LT4TQ4XRSRwuTSLv/kWfiYZvs9D3BG1AFED2wtoTxo1VYieCrmTonKWZkYA
SvzJErLGL/ojHvGEM/jE/+xs8B36pz6TDm2i7rC7B8Gwl+QKP6eJl7R/SGYw
+VxTjmRhjn4PfHl0XbRy+6P1FAbEzadw6SsNcIYUq75VwCkHa02iCXEvjKO6
U+ZAqxKihKcByLubhNCYh53T7Cm1B19vOMhEUVajJBgMBJvMY3yf+TZ7kIKS
RuUpV+p2Tj66cCoIc6zFQ/oHBNps4CEQh+pLPBVBBy5j4XXA8ktBBfVUv8sO
9pu4ZyLfHYjNEHbEGGda7F2Zrdc/r1MsaSXYC4Iptk2RfS+QNGcMC+/sI2i7
OKqKcYVn2WX2dU/PmK8qvjVWSfnSL1X2s2asRVw1WsC8xP4uZUN64he7Smkk
LQ5mzLiFwAXZIOt4QwHCSa1CXNa4JHDq23tZoFgl23NglOJLIsXjWahjdgRr
iag4JXuKkiTH2uNvWH6NXAfNU9OmjKfKf8Sbyd+JGd1yCl9GsU5iCcqAX7bk
jyRnFdHzJgp8mc4FD5qsf+sLd63kcxstgKCtRvBc/uTVUIOFNZCF68Ovyx4J
ARoRERw/wRIlGqstaFTq57h7kaPfMhELICoA2foYwtLuCZMndzOyCrR1I8ig
PGZBHOSWpneTADa4Pb1si7V2Uo//EcGTWLvPzgTdp7CLZGkS3xCxx+411pSB
x1ToU9EQHM3CYMxyH2tBFiLjhqEZhWR/OZ6ESsXJiAIHcFujMCTSM4jmLfu2
D5kH+YUFWn4/LR1irQspyT0ioDSU1225/KFGzncVV7HXKh7+d9FJrrcrGgvt
K/Q33iwAD5zGONAzjy8HAAAjPSoAnGQJT+bCz/C4EbXapVNi5a32T0AzE/sn
nPWTZVCMngvXODU7Kqd4ajxlW5cYYxaUvxOz9fuyJHuLbv/EbuG0qY1SvsNs
FumK1EfIlzljoFVE/2AyNOfTyHj2Xk/7ufSAkiamY8LkZjz/GhAzX5ucgKv8
vNxiTxwT7zmxl0+Jy3Ulg7fZN9nz0GGFbui9VftkWascZ/+GEYktvNo3R79S
oYdkvU3LdSuAQ8D3C1iU29ffEyRG9vvGxWOwIoQ32S5anEBCIv0TyHg+BQAa
TtmCyvRq0CeMDeQqgpqPNmqtsDCJulXoH9bwvsY0r19oTMz0cPDByu+M54FJ
an0t5lFfiFmNYf7iMsWTO1iX2w0kZpSlDgP/MXfR7EwzihDTWPOzAlQYcqC5
2uzqh8ED96ADqFHUFDcrBe6XyE6O7QV/3hVf6uY60Y8fIq4GkGRlSvQP2O+w
NrxN+4+YAkCWYq3J4qG/BnDwuV0xTGSqD/QA5TsU7LwJyCsGvn/qt0vE2eXQ
GbhLcW73vpoG53R3cygEwOyATrqoK2tUasCflRIYW06Il5Kty+N6r/BxNYzp
0VV/AyMdktLXXl/zq0rGVqu5/MZ3cBpaxsyNi1bl274NKMNSBVv06B012EOS
rG4TyHfgPE3nV0hJYyZhL4oTo9aBQOcJlX3ZXk24ik3IAoC9XNJbDEQiYOkT
0epHpf6c7EWjaYcIBcXeEEa2n7zMmVuyXzYj5YxcG4DcawGBodcqZuNTTWV9
tYhs7uvhjvpX+Cw5sKA8QpgypsvhD1lBWeI98FkNOcaeIJBovmNzkWxUDukN
VVIOzgX1ZDmHNbdXUKf/ooy2+CQYRMthOdSxNKb1VrCPV0m0qPfeRaWCc6V6
gyYA9O2wdpEiWv6H2B7W88pO72ktnmtbLpSB/dCZ76jAxQ9d2SuGrTQVImqv
2WHeDI0+wC0YZFDMNLYFueic6u8zLnPxi7nTfMNA41TkxOyXH3Fd1A4knE5X
ZZS7WpRCwLWHQmYyTPsjIccerUj+ltcVbH5e+IRnJ1uw8yEx8rzU+YDJ6YWM
GYQ/sAshG6OJZHUhdA1bcNEYrL7SfeJGDKvLD87uszQX894bN4bz4m3z3zsW
A820yg7TeA4Zc9EBe5QUbbXqpsV/8u34eepspENrh+ykQky7o99TZAfv1kol
A4/OoG0zwrHwgfdh695RdM8CfxoBl0jdHaHqWR0YZqwnS69ZX4Acz7Btro/F
jy3CvELbfCE1vbR7WwSsZ861p866hasYjFoZQw9lEQBqoi2TCqwFtN/Zoh7v
ZwvD0clRYZTQubY3rs4t6sGZSR8GAfG9AAAoJhyp8ECh4TGdrwk6kccYgNUK
k8A68Pu/qzXtQSTs4wxPy4tRropyM98gLlNYln3FnaApFJO3+Cg/2lJS30Fy
6CkT6asKFocbsDMYmuU/4sfypg/XkmuBYlvEOq2Iymf5ePjQVfCx3OtKck54
/JTbpOM9DF6qZ+zS8EYMLOQGdCjVuZJsWRAaFxZ2ejqLqARWLhCzffzgnlHU
V3zD/jiulqEZWPjyXmCqU3k4XlqG22HVwuneJlbLPhAkn2Yh1FC9IMYZ46Bb
TE8Xm/f8xHaEMRl2AieGH4lW4PiuBJNCxae83XblFx0eEfciMSkVv4E7KGlj
Mn2L80uFevQXFF1xAqnVKBR5qdpaf/g8guF1sXlxjkwXRTkPpFzw9N23qXsw
Uf+Yh4uDDX4Ddzqj60WlNP8vaRDCtOsBRIgQKoqHahzH/tbKETP1s3aRiya/
27EXX7mLQdf5SwprLE+nKSc7WXoWfSFcwBV/aWtP3MzHOvhW/YhJ4FKhscuG
u24ZWd31TBVUr64ABiT10ebwGJDerSIgu81nizped6S+nPV28sqqpNZn7zZ4
TFv+COPSip6J/so+5ejWW6xs0ug/PLCyRoRgXGi0dd9W6YlviQR2nCpp/2Ua
sGygthPN1fDdBTJPYThzhqP9ZOFrMxE1MwczzG4TkYXvMAF03s7+DMqURAW+
P3gdRriE9kW2DnzwSmpJ5WtoT728G1az9y91KZOYX9dB4vKF7bZdFDT9z0Mg
c73MAu13FFuoIkSU4f1SEcFXQSTyOBwdGf7LFrNSSZFpIrs9/We80nPhPmRo
A2aLc3wJxaXbrg3L4BjANCHZK+E2fnAJdBLc3K6PvBDOxdiLYg1mqnfQIKiv
i24HuQx3/9u+MGnkUltS5qiGmHdGFRlbKHdQXWExhEgFOkosmQjk+81ajjeY
QIvqCMV7+pP44OtCdGJCH3KJxPd5pXr7ne5QLYowWDWdC3PWHxQlAu/hxf2s
x9O1xkdb5EnMQl92tkCrk32ycbA0h9CmZz39AfKbbw49+lMXk+DhfG63k6UJ
hQIwaaaStofkCucj6tHx45xcXVGUmI2vWHsJAtIFUWZFhxw+OdoT3tIIUfk9
MPN+Y41TognlWFn3fQ3DI29kdKpSZMce5Pl+4o4ZD8F7z69DIiVDhSQ/PsR8
2sQpxsc8snbJs+z1LgwJVlK1IL4ZRCkf74xzYKiAg3+4bBPJAVEny9cAmgPP
lU3LKGCQAIKikkdE4kRmjdtz+0o4OU7FTMKDgGyI/vCd5xomp4GGZaVJnx9s
t2Lr3cvr4y+6G3CrwqvaIsohntmvib7Fi8yi6aYzuGYTvacKUA18aJ+AZ628
m9sFu3bjlA9Xc4Qt3d86exvnvtKtww75W60XPU0YpWAAtwqRmB9iveHKxGU6
mD9vR91EX7Cr4szZpYWpHUeCxD9SU6x4CriCikg5Thh/qnqXSntQqCn9pqGF
u4bUvMp2CiBwiV/YOq3FkWgEW6nl/W2ULce9gICSOO776aHgZMez62x646iF
G/XVXMxDPe9e5jTTR/S4wMHFKFieiIB+FmhihdPpA/sKN2Tlvfqr6Fj+NIBh
6q8gv+bbmza2og3oXYhKLl6ivpXzoIZZJ8Faow6Ve05joXBjPf4Ql+ZTVKgo
5yWR026H9ZAS/y/LDOd9QjWJUHtrBGPwQS0QJz0kUQAfVG2vrp+o4VVwArHt
4tXJour0mgRe/UGHRO2L2HGFvYLTQp2pYb+reZuHfLBph0W7iozxi0Qa80sF
8fdYR3zT9jHbpOVEyeW82N6dcTdpipk6kZJdMperN3NPeAmTPpuLec0EkORr
JABR6SweyMlQqXkVFffQYZbfa+gpflnayeaZNXlQZUI0RTZoSaSFRd4JxzX4
mzUDLHt3XzMjRfOkiFt/epUKV1YNIIqqR/CVRmEwuNrCahy7VFaT6T87OU4B
1LIZsRzN6+thP6Ef6XcIGD6VCSaCYv6PWY0dkGka9qyj7lPOf4OJzwSKlNkD
NQsijruW/51BCkBqWahEZyBtTLRP4Nx4bRu7cghloMFRWJ4l/wS8kvjEVwif
4ba4Q1ZDkIQ8vFaODuBojjWs5ILQh7OnYtIxQAJqDR2fL5zmrzoWUGgS7bdB
cBraM48KckfCD5EDLuMfXcZYX4MGWR4LwrjzvNm6kmniT2uY2cLi2c3/4dL+
+XRFNglT5TFhislk514B753/lV44MeEvDry6JNTt4YtOiuafajV4EdNWaq3L
45/04USqUtk7V4wjDgbNTbK1TeCJSKNggYVJVFOB2cYCoopyDmnNyEmnUYUu
7wjnU+zdrhy9RLBuMRgNHJ5nbzd3BKfglFeYk3Liz7lRVfIu0NnV0Iaq3+cS
TaTLZGYDKhAQV1IduiaVgO2A41Dw+P9lZT4OJT9ci3XUlsYWnU36SFDxIPvD
08GeucoiIgWo+re22K2bZQsg00JBy9M2WUVMCM+lhieUDBxhJEnfEmJMRtfG
DtTGDIBMNRWVcRx00u7ii6V9Wiz5wlIpcK2Ws6/vPDqYaVoYdR9ZiBNaK1ha
Dw5fkNTdDynv7kj7iEG+xCTgsqHcitSaI/BQU2V3wevOPXY0Vf0L9jO/mRqT
ZwUj+JQaePbNMnBxKjxUeD+WAt1dFCafbwnmFg6vBYnFT91KR4Hxesw2jXgm
nWCGB9T1cROkv08gB5vL1cA2LQpi8Oa4ms1ROQDZZTeq+pdyzUIr5W6K1yb8
DiLUAM9sNrtRi1VAk+5Wr3al+z2lwt6ysE+XlyaqD4UvIsSWp1LwAG/jZKGC
IQNCUW4SOBb2nRZJsLLPbKvfey80K++sNsIhg6vm4XKr4dIlUbg0nqhlzxjC
uyx88qkONiPyXZxnFPHIzqHTaS/K2LEh/RvJQ3abNmn5VwL+pL3xzfTmsCua
1CgqaO7NM9MBpbkRASL209xEbAcKJqKepb3ZhYYxg3qgUmNpkREjOsdd6Lpd
MLwBpw2Dr0dDgAa1kYXjeu+En/L1yYRnl7qx0rF0jJktGoSkg7Rac/4UtIUp
Hbk9K4jqWgza02QcNepKmf9UpXO4i6LcUWYGzeE0VCHdgfWCi1wUTVjgXQbq
IJewKQbfZuYh8/n92cc0YKy8GJMufa0zIngi7rVLPn4k/WIX6r2IudwSqjr8
iECTbt+l5Wn4lAok0cbr96zAObhrQtYxzruNGOSkcTai17/VviicuUM0ug1R
VJMDyDDg+7eYJY7jSDdkHgZLTxlWMm8Xf1iTp4v8tKBviK0JjOE6PE3/N9Sm
K5aHSIPoI9yD0xhxQzR2q2d0H6RdabSy1Aj7cCre8c6OgoBEHVPxJ5y54n4B
De4Jczn0Czym7mtJF36xbNL7LaxqNfjA99hIMiT/wPcwj03lzhhaOur3EYHr
B7KtAx64q85nOBP3jeJyJPo9uRN3h7/kyZMnSMviDOqbH6/tgxrp1blBE0rB
/uCgstQ4yzpGgQAedGNticIRG2P1XNuM4FNaAa22mvSj2bS6hOBtHp8+qaI9
QGvB+FWW9qPshUOxDIw5T6pjg/nkpHBQO0HJ93A7o+wC8gIhMdzEhEKae0d2
QJw/6co2+ito98kjyEz6lBd0K/v7jBNd2pkxL7Gf+1A+0ecq74ghtgd5ZNdN
Bb321eAQ6MoYA6Yg9Dlowq1jC/5z/jd5Q4TC9j7GibgkX5eCmSiH2caKDsF/
CDvnxxf7fGsWoZr4YJhmaci8jdxE6Slr6rZpK0P/BE4e9Q7JzVy2Of8KNJIf
V5Fwu4oOX1/HfU6NnlssvaCPnzGN56jHP63aan+gPVouEUOJ+ZbXcS0u9kUz
NmJhvunjKNSCFLbeE4Jfy5AXrXF/csf+asgEkUNGFDdpSKuMtLVkXw3u4PEY
szPNdQK/fGbQ/9Hmn/ZmgzwjeBK6KAb0aVnJ3AEwaCzWsH+CIhlnPOx6NmcE
TQEuRqLCbbpvyVCQ0v9yD51Ifqmg7AoFYMdlkgbx1cJLbBKjIDZSzgy2ji5O
wIEC4VmwHrC8LmTQfkzf5FInGjMzyaxZBt73I8h75PSgPGeZE6CF+39KIiCX
nh5mOEWEfLzqnzExeROmdkAeiZaiCjTrniZMDNFFJyAhckvWu0G3ZE/tIzNG
4RmOXCQNluE/MJnlzFoa0LN4/FYaz3t3p9ts5f71/w5vqgvTmFLJ+VqpcYs3
aIwSQmGKUESco8B7Rr4/sLqxg8pjLX41Cm+62yve3KZb3IoyJb1vGB8CzBZJ
xMJ7imVh7/TgmN17RPzM22QIlIylwjh8u08u6xQ2+85N4dznkkTUMZF7lo5p
sRzdGLrfn9a69qzesVYh59sz7J0zq/grnKGHNiEgcypWlb2HoEnKUupkz0RF
8AYqCb4GsAv7Hgl45+j7bw98Eyz3qsIoBCFtiX6/J/s1Mi0IZlK5v54TdskS
c/U9oP7LBZmvHBgEB7T6aGkQj7EMXW9/qImkRSIwK2snhk2N9cjdQ2zN/1n3
bhmZaCqX4tr4zc1xp/U4qltuged3dhJsKYODSU3J5f/oSWyfFIFXjrNS0taG
Bbk0IuWJ3jpqPU/ptek2ndirw8fSlBMHbZ1DGxofV6EXuM3Vwv4WABEHnAVQ
638us8O1RgeHzhY1No/5bBocJ2bKJIN9EZMxqe0qMPp+otnNNirV0qYhaaxv
engR/ruDq1uYgglHGobAXzlC48XNPcq0305A/BbjN7o/g3stOGL6HfbfOttC
BCVkNJV5qyzOSFwplpUn4/94YlQ+rD+DZIIR7aB3QXMs98cUZ6Wrxtiks6kW
qaKHOB3AqzZAOc1EBEgRzP/oQ6o8yTk5mBL8rxuDlusGfYf0wWefh70BCPtt
3rPRAbzrPzdhhhabiPQz/piLHBYJoTDb2cNUPkDe6DwQbMQurnWhIGyCXU3E
YM5zstNuZz+mJ+VjLPjQ9F9OA3EJ8jCUtrMO3biLK8WSE+08CXAH7rqKJHtt
4mR0MCcGj4Ur2eqICZ1/Q9yDhwCpBT3VxaGUjoDoETp8IrVjLa157+yp1e+y
mQh+2q09stQNHMSjhIrgk9kTfu6dzZsZkaLVn/26AqXXLBWXWLnWde02Yl1+
dmybuYf9t7KKDsovb+L156Jp2Dhzt17D5y66Oyx8BdCTw088BZ1c0zI2iyhO
sVqNYqSdmEvg2BInCT/pkGwCmAQN0rXjS53jOg3JwJWk13/i3zmU8wRhFCDa
n/B+sQOOWGn2qUXWt5TeRh/dpZ7lHsYRT9mwvCeHqQ6Zd4/Y2S7QNbAO64AE
s/cnMA3krXnTqMwQjylroOs7Y78/V/gZDIeV7lgg2ucfkk/xiddxqAr4DADk
Fb4iEEdo4BRVRRCT/ClnR3jS7t0PDRDnF9leLpNpOagqMT9c0QzXpxdGQTzj
aE8Zbf1JqExA7UlnTMVoZ3FdNl6aGFpG4815rHfmeyCpzJ2k+xciOS7v1V9D
mEIicthOBJ8jTC7IpxRKj5dDLvlThChHgpb63WR82TB+IgG9TCCWaQsDlLRJ
cwETmCVByVAWrgWBpCFPzA9O3GTmFwV//xSiSWsuaQ+pGZK+blo1FRH700pL
zhYy5ZeaG66q2pM40i0Mjq0mEaV9fn4TgoAwFuyOuAydwusMXgY5jpZfqGPa
ordZosMCVZFIHIxPGSvx4JYV3/DBHh6RNgY9G5aTikNzSz3U87sf8vwCER1a
5LLoxJsnJBbKGXsbTEtkv4G9EJcJuhfDxtozKRMMKJaSo6Rvfje4pBvr1Kt9
ZPX67g6FS4f2lq2CdI3pnD3wGRmWnZd0OBjlvXx+LGia/MERNI8bB0wxL5Sk
5jroIqC4ANPhd5phMFpSLKYCuOdRvBXVvUc5w+Yr2OtJxVpMCJS9503Yyyk/
5Pt1zp7efUAIGU6Mq/6NbMLpe6+791y7lX9528xCQx1MfP/TUJciLdmuGNiM
ufkwTeKRNnTwhJ3fIk59fK5cYn6nadLBlZCe3V3vShmo2QBAkhyLjmsvwrMp
8Q9pZLVoA5IU9Bc4kujDeGMaYbV1R7GazX8PabQRL5hptQuMo9pqgF91ShSd
/q/B7C2hP52zTQ2QXMPXxXjsrep9Dg1X1bM3nne7+fcEbsRkdFg/bebpuqPl
9KjCGC+bLRan7iDAMC5EwN3IJ3QENBmiBxna0AH4gLGEDf9nBBbYN/sKEep1
EKRaeUJLlrx5S/vHuQHX1+OB/59yl7IhzVnRzCQbf14YkvpAuE2Pj3l+Ruvz
FyhnaN55J1B31/AO12Y4+80Vvpg8yINOKSZr1qmhxGMD5E4b2fhP2B8FG7HF
R2K5II3bnSJwWhp8VYYxuRDu/FZbviBEQ+xrexORJz8TiaRKIcBfWYckBt2q
C2LLY909j3sNYzX2AbzELvN2aK7dHNlIUB17y7oONeJxqKRV6w4kwYpM6FtK
LMYDB7S7tHva3PwpxH3xB+1SYjbt17jGs6YXz/VMghwXeiymPDfjS26zfsB5
TZHDuCrkzm16BPP67Ip2mq3J8rv3l6A2Qduz0/N14wH3lmCB0CiQFzGkJ8xs
x+cNyj2qDZqNbe6TqKjtL1fUy+JQgFAZtTwDDnM7jAEMHUh+epUj4B5QnIxk
HFbpfgnKkHfi/g1FdFkzcVB4qWFOGOfxLuwJc85HtsGISf+yfQ1yHvMjUG8o
lJumY8RtmBqIfZiG78KgVKO8q+QRMt6sGMUDs6npWK+WseF4dTORETIPpnIi
sG3T3t/YxBZ+e5RLA159Swy8MrPjy2XgIbcRBdopjnrTQctFTx50umEegUUy
tggn2Z8lDhoLMqngabqI94yDh1nHk0EeHW3MUyMR9nVw8e8WQdRwSB5kln97
YXgSxUSd+seoqLFQ5VF2wnbVNvvYTG0psnKuFdIR/BkcUP/p+9nzurnzSoz/
vr+TZtqe4QcWvehkKN0hOCJj2B902F5sVimM8/clZQdzoBDma8O78AnrQKmo
vkbuEqUhfp7zJlSkjJKZCbBAMoX6Lo0YdpeJ+cfxit3xgALAGyNhOO/MDepf
UQFstqCbVgZ515nWQSJxdSHaAIKUyoMcoCFavmBCt/r8M5C4bzT16DyZ95dY
9f9OJ9BhYdsQi3x+GsZCjCkqaw5JxhQJXJc6ZD042FUgM5ZJoybxwhYQhcVm
AOmINfc8oaSeheqhcyzo7FwPl9kEE+ky3/NKd02nmiUHeVrwWeVQJuFtjZfa
C+zOfU91RMqDbqEFnlTZV/6OrRgMxvvqjnLzVLPoL+bBSBcqY+TJZvfyi0Co
u4znUxxsGdd5xejf4wrn7qsatOrXQZgwKcuGV9Jy6yVdvBEwJCevEBe7p6Pw
ZGe2mmfIqRL6oPzuNuGWw59Y2NqQzB5JmQUrKqYgAEUF0HGJmY3vldQgfe8+
yGZSR7o8we7bLAOZhBrX/2tC9Y+BDcrAmniaPR0P9h0FZcV6/q0XXpaKdOjx
HbGO3v0MtBBz5sdFtv+TeOjK8zbhZXyDS08+nqlJ2ugoAS5hCNn8XTGPftFQ
gVTB7IOfTpONG0jEAJkkG4s4bnM545ntkCj3voJq2+beluPcFwdNGh92BW4B
yPc8J3pTj/9x/KYg/WikTp6tdn4gNab796wOSiaOaIxeh1/LWazccZljdEFF
K5ph/gxfMDXsBjC1ScClzbbX54Hg0UbQCbDTnsTAj0jL8C3RHvF/FxUgAn5l
OyXyIyZ/4y6Ky7PM8T9muE87sahjBg7AmX8loRZSYaY0k6akxuXAl4K/nDmA
enkIPMc7axlmUyuZLLXl/fkRitZMkKY2v0fK8Bygq+jzbqQYUtO+poie4tAQ
1FwshgYUHcnA0M5J0l7l/MNC1mYvK0kCYL7U3RBcdynSwyJ0BQAJ/2ObBTTY
piufdMSui9gh96N5+e+s6s6h4ShAPxdtJw2Hdxy4gOYdGqAEwpPhSqu3xNkC
yb7C1BraaxYQBujc9eztXtRCOftMxjRmPw9UNZWznGG2wI4LOWbzRZM1/k48
VdBuf1aDD1s1JqemeHFSw3w9O5lfFDvKZFnQ5GEsapJlQ845kXvXDo4FV2lD
GBSRxvIT9NYokWgC5YlPi07DAwA5/DykbmnJCdOaPgNxgu8U187P2VvRpRLe
1ho2XmK3GHJN8TbxVDgAKXBNZRvZIHGhFtuKJ2m4rjuyL5cUG8ZJu0/zzhVx
jqOkv1sURaILhr+HZ7wooxpSKbhHxicZMN6RA3GK06GzGRMBS+62hXc7I248
bdJRRd3t7dpPurUKIHJEU7GHCpxDADZYVCgFz9EuhIdKu04MFqvMkHvUXOBG
Fdj8HtuH15ZM8Lr3eYaXbEjrMWbUxlKSPeEy//fF6xQgpFGbx2GPPhyOCY2k
tRW8Y+EaIYljMyA/+OO5QOUXmyFNS9acbl31ReMkufcO7cGTFPiwpkc4TwtT
CjlIpdutgxBOVVSy4WIY1DcANl5OlwUNXqFxB10HoEp90ykdJfRNA4HZIBmu
CklqChtgOG5/a5t2UEsV4UB7G2Abe1ghqvTx3TivbKEuEMlJFIbIlsjXKqdF
N63ggMtNNp+XI0hUeiTt54MEL9KDszDuKeLWrcrBmhgV4qKN2zfGlK/ThbJj
pcJmntk+nEngPQnkUxs1/cq59uEhzTHZGh4wf7P/hL6ZrJb9lftMKTCuTsHG
MI1FZavgJQVMQFJVsOn4lWEIGads0Cnju03mQFwvlu4UbQ2Hn4p9Gs1lhHYj
R87nL3siY5jaqPiUh58GdqMCFZEAxpKmD168cJD2sntZiG2gqvO46Lk8BL3P
aQyIGgb33366U/3I99/5ELBrvpYCQuWsjwnxqKkbCLMfR5AStusGgQIGEchU
GIvVf+AUqDSCC8uBAZnVv9T3tvIfLuAHINr51Wx0bWkYXmwRHcd2EDcxqtqr
OeDbj5Ht1o0rP9f/DfVlRpJ3cWnlUN+Tpqrgw5hE7NoJXCQP+uyx/nmp+k+w
x9Ni+dihIN8LpgEx5F3Z5POuXGeqdvoUb5ypBRlrvtunobNuH4UXs7Xj9liv
LrRmBDFeGjM+JXWt6xZeSs5giPALdC1xar5dt6S9ykKpiD1gb9GYJ02aZmNn
WRS0yCihsh7wcxBkMDfp3Pxo8gaHEw9JpIppK98+V33CDBoogY+C/zcz8WS7
L3SPHFXu1Ds0XYmn9716pfY4VldKGMmf9ghZHtLrBBmTGEz251ZKQaiYdORu
UJGGjjPpZTDFr3G2HY/Pe3HiRxLYsujRXTTzlsMuk1VXSALuXZsuTLLbNPLC
M2huI4OtTLQv9QpRELwBaINuATx5dF+7a1YLyynH7H8/AbpMApEa1HWQiT5Z
K0tOOMf8/3ehIub4GtAoeqgLIIMaNCPORMD+amvyh2xCLtfcWXL0tQOo7NY7
1oOQu7PVf4HtHfB0Docea6HkyiHnn7BVxAs189dlrq5mKsEr24hce8p3O5xn
pCmMMvKZO0mrRuWtLusuWExwOjZiOxs1xpmqf1Pd1aiN5SR/BGc+ONygQd9L
GR3YUYSLekIssTntukXk0zxHLgZvNqnYx6z0ow1iqMPK5OA8SIdjXY9rnxLI
ksshQNI1Ati65xhOO+oJiRIYNFDUjRZvf3U7StyIzX9jTtj4/SIa2WiSgfJE
l5V83PIiYH4tfuu9hRfs3/HKcqVEEQLJL5R/wucc+iX+GnSblK3l76ItrTUH
t6zwTJ0Y9aMBvtXCpzRQOofaMJ9WWVLL8qzcM7JRzSQ3YCqYWHShmQ+lkQ+d
z7JdXjznYkYLybKY5Obl2OL6agyEMKJICDNTqXNm1rRSA8hakOvhMUc43D9u
4qDnPIGJ1LXesUpH5dg1Z/4v/BcFlW160EXrtA3FeJMprnmdAjcv5z11NxGA
ArYOmVRL+Jf/lKLQ1sTppQVtNmBHQq/x57YlNrQ6Xqb1OfZOlYzv2oHse3Mb
1KfkHFILujAfbxZizuO+MpGDu4GIzKm8FWmwf8jx78x5R1mXVfYiW7WYjFqd
jM2ce1MyWYPo0rTJE2zYSJ8IBttW7XBnms+/7BkZb/9khHR1OMPcQoonms7e
tzMfz2oxow2qji/GuiJQDruxEPSvFM/drCs3tdQG9DkFxyaYClp8/iiEiUxa
qUpyIwqJeDKcNoOXBNL7km1MRQMGECvmaIiycaj7IHjr2PGTugVAe1gfT/tf
bn0g0BWHRaaivTeBAeCw6y8C/6TbUUQE9V5cuM1trjgMOZuowfjTO90PnpC/
WkG3fx8H6tPwIlNuSGvlg2cZsuqZozdU1ACIveWRxp9EIjaCHka69dI0ZMUu
wtq9V4M33/N4ovbeXrH3lAK+ZxOAlKTNjTQA0pA59aDfnXpoH55YmQEK1PyD
G53vaPiLEX4dpWW8d9kIYduAfMJ4FVeKI39fqiB/i52gVIqgJZqxO0GVl28v
lg8m8PXLUorqpTONGn+/lhgFkPONIBu24WR84inVBuPlrMHhSy5/3atdQyaf
CWu8pbqoOOgxR/vrX7dNBNG9Bx9Okm8dhhT0Ia2h5najmAzbo4tJlpf1cU6+
SAkw2dP4eAbP/jl57jx5uTh2F/jALIMgbI1fIS8ru2RP762StGFYdNcNqDpC
A/iilZvad5QXSkmlhsoJf4ZbwqZAj2DwZY/zsRlfZsfFB26A7S5yI6lK1AvM
2d+tlwxjVBuQuPChobaS1wfXnFrqctpP3iyIh8JeVDaYzYReop3YwvUUp7t2
QcsmfwkalST25bz2hm99Ftm7efal5JDedojHAE9V4h6xmztJaMb/kY7+Qtej
r0wCI6BOU1Gw1UkxJ4XJGk1Yn7NAqIwKm5JsHXg4V9bxdAKrOaAn1F9qpEX+
RoI2ToYlDIFhNNNDrtvyKzlZe8uTX+2ZJfW788AMN8LV5Ne5jocfj+WhpqYE
/0EO47hEt/2L9DdLVodv/3REAzlhIXOmkiqvIII+Rowmfs9QZqnGms6oqggg
yYhvMwxISG5r64EzO1lnssW0VfFdkLvjeY2UGVFlJEf9nqG3a8HablEueVg+
D1d9334Xs08rpdHgD16mhNXhMhp0MRFLNl56hVQs1ZhmBWBSInrxe/RaJBd0
MVT3hsFnJlQezdF67hB+XrhrUThfljwSAw1u8FgniDXDFW9mAf+yU5Si1x54
pk0ugtyVP7kjlGe8i5gEO1hN8b7FEiOJfdPY8GukNT/OYKxvpagarWw7lrJD
SWvgLNNh3X1IHFjh6i2B82zX0dVlA27wsacteeojnkj+9CPaCDj6O0OvuIoW
eTyHGw4ZtH3tzM/s5QIIUlQujjAVdgbFNWekJVIIwp6RYK2IZvZA8Av3CYAQ
PkL9/zqJ7dkDd0Z9kq1MHocn1H8OOjiCKf5rAOGNr2QybtNntpPaii2cvYcu
r+YPscNrknTsJGU7fbpQ82HpsniJ+Pt8+oL7Zc9R5QFkS0RVUwSYvHPI9oZf
oH0f3NH41v78FXczkqMS+AD8uvrEfC7goXqI74phyuml0jhMAbxYH2/hS+a1
Ccrs6K7Pzugr7ByC2FwwqMFhZyM5hiMMWULQ3/NhR91gGAnfW0OYlAHqEzPR
gAt2de6mhw8TqhI4g6kQDd7nBsgCv+/57bQ8RzS+AX6SFzzffrUzBZBMeGd+
QwrFxyps869o1m4bkHshmA7in/XX9eAPBTO2OMKOVaHFwQSFYo9kuAJ/NjhC
fKK7L9PxzLuogaH9F+IEC6fnzxUB/sC6Za/LjJEdQh4ydhwUbbev8MnooIWn
twTrZRLDlwrenW28Qibz3Y4g4vqeN7LIVBOxnJRxyL2E28ts0wqGbrJJVLgC
cgETfpNXUv2C+SzTYXcnp/kmVZllpnhXpU1MVSXESJol+6zmGx6KG2Dngmfi
6dbQRZCBEQekP49mf3J1r2PCpUMJZf60V+9mpX1xjTt9FnlRfhX5xcub11rN
jjIpuk6XIeowNLpU41i0F+5yY8WThBc5cl2nxiCLeKxzotXWDP1crNclUw6R
2TdwN2wjJ1IQHi9myD9bTmQl6dm08oH5ePfGq1RfWHLG7+uo0Monq3zORUe+
i1lmgVGI7hLoSR8R36Wpu13eZWaLU2wPrLVGhe4MXkGVlq1Z11jYiR/7uwwW
pkVOLNvQUtjVYdKcaDZnivfsVH+XKKPVrLvekuezrMH9GgTori55EbsCxmNM
Jy5JUzcByyJbtqyUg6JYaE7PCltTd4tHAZZoHCuY96+dscgfrsD0R7P+/Ec7
y8gCy1jMZ+pP4gF/L3F2KNQLdLY4DLlO+Z2B6SZc6X7jkjbeMxJGK5qTGqHd
4N8Kh1+gc9rXRUMr4cr8ptF37wGgUXR+/HDmmXgsWngIe60XC9TPyJQWC08a
EBudw2YPqiBzWzu98gf3jmySKMejVmnMElrSn3DW668kxnSKs5HHV2tK2xo6
DEadciLLF6J36Cp9Y74gP4HCuE9fXqlQPhLdgBKW9ot+p8yOYSPpOPtBEICQ
XnPZWXS5X9NO9qbSU8kZ5O+vjLVUBMOzCZwvKUS+2VGAm0L5U4KOUhYuYY6s
woL4kI/nDVXn/1TRjsLWs6UVvD4RftxKEg4l1QcJq73SKkvfNzuaXu81e/F9
GR+Z2f2maS6IG+1O3elLf5QSZZPECsBa/tw/9KDEsA6l2SL0RHoKpRYf7sBq
ywJJRZiKsRFLCtfUoRKGFqvbAZj/76Em3xqwDHiSZCRguy3opPxreE9eSu4r
9sgI3BfLmQETVpNo8tIPff0L5FivJxzc/ohadTm1Q8H4DWD0l/UNjqKsx5l/
/a6goumnpyDPOKKSRVA6NSBYTV7JoxEbN764WlQLWAI/XBIhhk0Z3vtslKBW
lvUOO9LECrVNtKg1tR5/X62Brd8WP5VAF7/Qes7im2Zr5M7RZEZOBycHg0KX
Dsw6OYY8i9H7YUKy011uXXA1xURB6nGPKp1Y/t2Gkoe7Ciaoo7hmGmhaNSTq
gwtruV958VzfCpfTMqNIfOBt/EH9Uckc3uAZ2APaeVCGQ3xdoZrj13HxTEVx
68Xo/1rZxHmOBt1mknRk9sdlAbDl88xG4RjthNdDmih5hSj3JxMlVzBzWaWZ
JGPVDnQThUCxxhRFujqYEagWE1I2J+edRhL8skuM43BI8T4hTp17rsrc745E
i0VTD5Z5DaMoH2atnH89yf3wg8tlUwENAQoduZpN/6klSrsrMB31HRt1mRhY
rIdCMrDT04gwVT/6Dx/8wCRPQ+kkzxy5BnfAqGz/jUoq3wduNm3kQZeB6ymm
sYQrw1h44TrdMhEm/dpSbCLiGLJxB+q/iCmnh1WbeGvII1wr1sg7mLgmLql7
DsU4IjW82XS/BO0X5QBDMr88ks5TZ1u8lss75a/w8ybRVc/sqCeVOnFqFsa4
k+f/BXq/N0q/e/Bs3WRf7mPO3R7rSlwkGS/oCo0FHAcpTTP2H1eWiqAcYNfw
VO4h10lfEQ/ntICS6rMLOwE4+3PQBjebRaX1tpMaMJsrIbyvxL0ZDJYcVE72
O9ZFjQrSR0i4RM1b/OxObr/N2ri47g1Y4ZG8dRyNkdgQkwNPQ3DL/zNlq2n6
75FjnBHEbL3yGQmKqiRNAZFc96gQyNqKUl4ZVP6kaB1OgVKibu3k892gVMra
VcryjXfVmrrzQo1xYMAKOWkLlrPTsiZD23kM+Cxlw282psEN5kH8yMAkFqGi
mvGs525DtlnUpMueti6Vie1BahMejFqQz4iWFNK/ZS9dKBX0776vZJm7adPN
SCA0iIHKw7YnRF2op2OH65xCSkxiEm1WRw+eidc/Ck9imW2J/3ktpXHochrM
R10rsOH4cGyQvcvZAEW1E1IFq+EqcCUsLLTFYH9Wwo5F5p/7GAjfo7ve05iH
IcSpsiTAlQZp668p1HdgjTm7FoYV7E7Ng9Lrq4GGPxA6ZMoB7qWmk4014ZJJ
762BMLQWRvH9n6BMhHxTeXUZn7J2H6/PmEZdl+bqXhCA70dLMIQ4udjlR9bf
CKq0ZOb4MkBWrt/DBvhNhwk/XM3USlMle3QrpK/+zowHgZSedyPS5qq2pMkl
CGAK58Gs169MRM1IdWnCdxYr8GkjtkFbGXH0TtRVNPIECZ9FnozXcu040Oav
UYZ/XOEYgB38O3hTxFuqK7ozCDPGXNbSgW030+RJbw/7YyBIBzhMOdK5sGmQ
0eCkB93lOTJhwiv1CktcC089tJJIVsv0V9wQof1TGpWYbrU1z4w4ALZW312r
L8Z03dUVwnRdDdiUf4klYdFQz2jjAEKmR3mWk/fRwMLpTJbTfgZcKsSMAqii
sdmSvJc6P/IsJ0tTCEKrsn8T4GvoyB+Y/w95FzO6dcbcbT89WlfSSpJMA2zg
pnSvuQQadZvQzBbIoDQaNxBZwbd+NlUf/GsO2Z2MRUlEEel97b6LFCwESt2G
kncSpaqZjreaR0zUTOPbUvLPWTBs1do8qwSNCwMEI8Ag/i2UFz/uZhW9wyCj
zYe53mK1U8UP2XiJffGrZUt7BFYt+30IH4+2PnkMJS77yhQw1BtgcAYpSBxO
E7E8c4Fsa9b48FhmfQEjceprLe+lDrSihKejxCWdMT5tAB2HpkrB6Nyw3F0e
d8Mlmi3SeOv7t5wkE0CC6ZqBOgrIqzn9DujhBK2R9LOOpeA7WjyKPqBat/cB
Q9g9Z+QEwHz/yn9dwIyWCfjpmwC6pcLmvM4lSyW7HQb1hTCvoTpkzRZt4OL2
EJ8aSz4Gq0sHbX1G69QTHFjxDPiC7qhpfS0txIKMU07W7rxBN9Ud7LymTI1H
WxwlyXkUgk/rIeABqIGcVBx/46bls9Zfy26GfcfXO2xpJZn3j/pmGLspGgV+
0kIenFzioL9Fm1CY0r4KOkIEb2BzaSjWv+vsmqOhcCrEOEGHFgwFT7N7s0ya
V7irkoXajHi/FaakoySpvbpKcScl5JkBZYyzhImjDaA1lHGcyuskNug3Zj/8
PNZwuSTYH7zib+OiRtNdmqxAO6z4fWLsImOWEmcOBteKjRNDXWm2J1fbpzev
Tpz02gN986unKdrbICdslSOEHRI9LB6e1Cr24XZE+euk793OYBmZqZYksSzz
1NtDcSJetKff1P1l/gFIJayrzzPmVpruQeW9DEQZtVMlLdYPRqOa47kpqvM9
9ecpB5rd4Rv7ABQac6rcUToIYUMuI7wyrCgGnDS6o7exLjz71AmnAwHW7k64
1keIL92FVR2te3ACy7jFIguRnJYCBiSvaCy0jGj2OntC9yPZF/tALsA9OQhs
cDDpz0O25j6mJuwNUEtYXv/5Z8BmLguUGSh/eimVYYZxhejmWWdDQYubCmg6
xln4Tfx8JBJd27eL53LXC7IENNwFIsRSULE0/Yv8AwvrPtcoVF2JQlkMAeck
FqX0E76iKrneli034KH3L6fnHBKdXvbe/CerB0frNIXvzQcdeB/U9T/Ve7WL
IU0ovsURHCmZKlF8vlGo9UJHgGcuSnvntDSj34l5+buymDKok+yTF5l950P4
8ZyzY6LfdmAKbLCK9vkhpOnazJNafdCE500Je28nImh1jUvJludT8EKETWxn
WuFDtX6Qbszt9JeUTUJGknXUSGjLCfnssq2iKEI7+v3EGzFwxXoBObG1QX8W
USO3Nt7zB17Z4d5QgDkxXN6eBLKAstbA4IfdSeSQIshQlDIE/AOW7WQ3VvJo
GnDEp/fD2Z8itATLqb41YbCGrPi1N8y2/OdofW6K3euVPXPbEn5tF37hT7SS
I4ERswZFF/+Z1qjC/9kTepbNax/v39SEQxl2sUkChT4CnViNKtVoSwhv22Tu
kw5FQb7lNx7GnJ/nj4s1ChxN/PPZrnZzZhw9q7PEXJ4+DW3ey8lAvFQCgA9F
blg16mpg7zl50JyLyWu3o04a8nVkcK7YBeyDkLK642a7i5NrGkyTsaZv7QJx
FoidohcscvHLiAYSOLL9OrgYgCQ8BKkRKtLNn+YsrP5AxgK8PkrqILumbU1r
xiHTB7QzxqhC/+1WssIQ5RqrGxUbY1REfn8fH2K8QU5p6Mkz1WcGwiaRI1Ka
s5uTk4xGTa7TkBR39YrYIH0ae/Lv3sgf5Qz2DDh09x59iMcfYxe4QEnoy+ZB
KIV3smYuvlHDBPwh7vpKnDKz3TRReAGhzN+0cj/V8Cti5f2FgrgZXvou+1o9
5geYO2jO4ZGvkeOi0zCQ0TLopvy0tNX3Mpb4I+3jiyuWDGVy6J2whdHcL/k3
vC5Sr0GDVFiMjYyDgVOEloG6NiC0Sr1fS7lWsx8WIL+b2X8NLZLa2YGmnchw
GEWd3moZ+0gjsDu8xw7ghw9rPnazmkUyHaFJJps/ZhGqDJuyspQ57V98fYKR
ArmcMM3r0ByrZ6wkLQUSN2756+FWauMn/kcZ53etenjPD21K1OGGBCdiuw1l
0DhUnkLtQj95HJflD76u9U4a93LfeJhWbhGj8kPu9zpIx96YrEO2ZCBp3L6P
G+svecJX6+3h/I9e8U5G2/scjQ7XQtlz49cWMg9FS5jHa+uB9Bn6X2hJpAx/
hfAeCPySJywaSrggCPHAfBwEk1USgp681M5JgntSHnLnzUpSewTdMoWM7s8G
La8+UgPIq1bLK0F070Pjs9c8g/9d8hwnS6aYcwdsQ3DULX6IzJRQ0o61xlXG
bEoJs2MEByi7wdjS8EK9hPahDq/4Hq56zgiYcV0YebjLkfqWbxmfFyryffH2
GASOaCi/fOtgmSayhokxPRMmkSA9GmZrkqZxw9Uzk+Oeboc2vEHJ+YY5qaTj
xFAtyRDEztGHl6LhgBooO8WlGL9VQIf614cGDTTlaixXIqFfx+lb5dOKCdtu
blro4sE8xGi6KwiK03wnDkAcWJ4BA8TxTtwEJ74dsE+ozIyAp/eV/fYYlj+W
Wq6WEOvEJ2b0M7R4Q77j4PZo6HLWQ3gRbviWyJerwnkTZmzW9BI/UnMmad39
Saiu7xkShA/f9eDoI+Q3f0G+HKnmvXWRYqFEg+Qb3j0ixkFte2PvqDbAkFAe
GeLn/zU/SEHIuRscuFtY/kk4/VyG+C+2gp1azppUNChMD6pBmD6O74TaH1nI
qh3hUpQ8C4B+5NK2eNTXPaEofWADqa/9pMhKb/l/LBvzP2mYHnczd0E+sqxC
ikcyUxspoXyGGAWdV0lo3lYkO/3GddKe3kE4h7Cfi9Xp98YFIjm/SnQeHNvn
fMwwUSCsPz2YZBDSgdLEbH3ALpeLkTU4i8E83+yvQMbRRRgG+MPtY+8qpTyK
9pS2KfTcx/uSCBJCJ2A92HinSU1tbzZcp/cDDeCrC5ARhsd2jXhXHyllXhSS
msM5tLTW9F03Us1d0/zMBUowJfAcGNRGoMZ9/8T8lRUqdi17XHAk2DPl+AQO
Hb9HN8ZpeInH3WHkL9Bfg5W3dIEZqZ+FEl2ZNZOB4K0z/VrKNK1GYEsUIdhj
zhfl+YJqDDzmhj8GjGOZhXD+Ukq7BzRVOjZAQZqvh7pZj0TO3h71N/tMi4bo
aF3XRHJR7MUBeJFO275zBybtFEosDRfaNe4UE8IXGCDNQ82hCZcPBOEd3GQj
OZKCyarV3NaiiQkuQdOPDYjTCN2Mx9DxwiFF0VmU5XD4tgWWMuuA+INJgxE7
Oq9HMCnokMmq9H88P0mprwmhyEyHRf8OWKXkW1KXSu1u+pbO+gv9+bCvK5Y2
lZgSqXjIQsyLMquNj4DEyCDVLM1Yw+P/65jwqmHfLofAO5nLOThjuScewwWw
64FTeBxc4np/UZhsDv9VHBSE63sw5D+qTkmJVXDv7KHHhkTIsdaNubpVSeFK
CdAQHbzfRMv5J+grRT5lIWc4giteTnNwa4D21Jzw4snFo1V9cxVXqVu3hmLY
K0F0xdIR2FHusT3FZMpqmwgiaD+048/sjLCb19HOpDBn/ZQEFyaOGnRBV73m
N/8o/sLx3SUHctr7Ir4hfQxHIN0LU+4lEYrnTcvi+tjIXActz7imkYBDDbIG
vwJNDadz7ptPDnbYeaP6YWlb5gCs7iQXCcKECPWErdTGB+zG3bJ0A94OKZ/4
Ef4Zc8W5p9eaTmUVUHC28+j/Yj2UnYlmNNCGZ/tpyMijVk6IZYiC7HelAHGa
X01xMBqV1mFgOyye4maJ2ytb3Zj+J5Ody54xoAj/vpXdJLMQbz6gStXBPmw9
png1LhGxtnkMTKqZu6YOfdwYtzbfTJeMAMWlR8oMFMgKXxkqg1TZRk5nsehd
Bh5DbAX8pQh44o+ywQDXlTiJRdnk09IVWviICKCoAMFGgr9m+jSDoOlDkAG2
ORt5bsVAesW3XiYQwnJgdMYBRBTdlN9y6CXGyPqjF4bXrsRZU6icAkgzbcxG
bq51ycbkyKPFEeFqvCssgX4O90pcERXLSE9eEG94cD10FdU+fK/67wWKsgkY
7n3fFcbIoritJDNUEm1xdv6iDxI1aBiLFII49rTQ5VmYUVYrFM829D7oUpfX
cWiZSQYXm4/+GDXyCAK5zAVKMbJxOrhnhgZroZwh2eJLFE2bXe+nAZoEfoGI
phwBWtY7KQHjYq0TLLOQM/16xW++mEBPkNQL2/pKhm9sBU/KQ86uCvr1Uot2
jkTugmUxrmiigXKzmKnBZ1hHw1YtpWKur9m8evTBoyK4VJWe/4Le5D+b7rBm
mrddLn76LFn23gan+u09ARX0wVpgBDTeam3BYOX5YBgsCprmVSUYLO7ffXye
orllMZ7/NkL+0eOeR+eM0FcKZeDo8LvhJ4t+CfNcqg2cddwCKtKW3RN68uWk
wSi8o/0ipsRN0O4KwbGQYGg+MEbk/a9QrJAq85Y1WUHWy8SJKah8+EAJZETR
gY8HUW65xKby4EA1Q/tiJk43dyRqqN2+jOnKiesU36HEMRvs6Mt03oaZz3bE
0Tx04dhmReMUqkhxtAc+BMdZxtomaKMVQYx0peptI612TWLqVpMYBCWGXj3G
fgBx9lZrc1o1YawkgnKRR6fUfrgxdAyhwT5/Aq/geJf8IZhDoLsA1EHj0Kw5
q0WyNu/ZQrYOTC1Wxc7dUAKgH7YOyWPZwp4GHVxxGUwHgwzCIgsnkBiarDCm
PtYfvD933/XYlwQXyzPF/7uXXuwi+aSckpfKVfHNdalpBhOlHG357wx6JeDL
/RGlCXz/T5J2hFH17w/eP39GxqBDTybCdwCY6ZggnD9tNTkEcXmMZIO0OGX2
Qq0lEDe7DmFKh6i5TV0SR7VRpfpFKeMaQ4T60kN2KEObteN6xgwlDGRZHZIn
Ue6LvCjyEisYLcm3D9CmfdgCAxVxedjs2u2N9dOraUPLMXXZD0zmXHWOqrRM
nVFbQjCZ/12uC4B8pBAdHvZ3aYtp9EgfoZR9wqFhi+yW9dLuv4u8WubcPor7
gqkH8sLLd8jNcnVNW4JQn1x3x9zzCFeeW66+p2rd9+N+JCCopjEIkzgmqV+N
iGXeiuEvC+RKjJs7pokmH1cmyuX3NRXrDWMzbpfOYXdveQ6MCLUBIfAO8Y3X
va9Xebpp8TLtiId6HpFy5zyhsXZl9VE69GKsOv/R9kTW1dJrnGOtcDR/p/XL
5pIHfwtOdyTd1Mo2mRq1kzFKXJZ2dMsgTVM4fNgn2z1uJG5/mE6skZyQm9ux
3BHa2RjumrmeZR2hmOMaGMCdaIta3jkS0ZNpeYxsRQ6/hV8aR0Jmel6ldY5v
uSgz19UkY4Kdp+xeyD3WHsGHDxIoHT7xvdAqq7EFf9RaHlpaE5vwdcpadBRP
Bc8rMfEJx0i1urqVu+3Td4rT0itov2Ziz7n8TS2v5g4dPiwEzvY97MFkST/y
nZDjbKVfV+KVwKUKT+RqvR6u/FVnIrC8dmSQAidPE5f9sW5IdpFwxh8HI6Ot
H7TYT5zWLJhpMnTY1YSXFL0aLwp6p8EriHMAWBq3uJjRU6sLEgaUQrJey9Oh
M3RUxs9McNT9nx3QgBOmqyRiy/c9x+8pR+QvkGugyFXWMqPWXtnrkd7RbWov
TRvE9Eo32mDb/UitPmSxcNCVa122h8Q1oIngyEuhiXgO/Iye/HMIrpdSWxu9
ZBgXV/Njj/rZUzcd1WquSdspcKdO759BUpMysBSq/JrR/aUmxA6veGoPAh3g
hd6bnSb92JpqLD8kMAqd129ku2Vr+wGIEPBeWZsSNYgKr6F1YCZyXQMXgaVU
HbJcYB2RqjOdOMUJ+ShchjOv/kTF8fgEHcoYWa2WcIT8BpbBI55+MG9erKlT
/dgcnGseTRy0W5hQufwBTpbeWmLhOS8xz/n9y2jENmryOSiYaDENw3clAUhF
dX63kUb8ABMHJwhzURQztNh3S+mVCPnz7DkusRIHkd1Lqo4O5lPxLssaltAG
Ts5OZimn2rs/6J70pTivg7ISUA6msY5hrGrai4w0BPSLkUqslvehLsqZLk9Z
TDpRmTgXoeMQ9/Ov1s8t4KSTKmewdH3b8eRiqN/xq3n3MRQDRWoi1MXVTwQX
9N+f92OEJ0laDqIyihuOawAndC96KicWDcTHZP005iCRJ/CaoKPjmu6eTvdt
bfuNOmley7APPZHd04PFQv9CQUdhEgXBP8//5sHn+nyIM5M0NlB+F8xgMySO
2/+f6Z0l8VPXzxM21YVUbkqaW8ShKSnSuB6cNivs38Bzc63c1Lp7zegUDX6J
bUSFv0rVyYgAKjCOIjU3nEsFg1IKJk83GKxKZPbEdn7wmmDM1eA6bixcAwZQ
M7NYvKjG4eBJ9syen0+i0/4mzz8ApH9zs4kfWcAdYGxXBvNDviNY3XG3hr1a
FzhqJJXOXRn/P7rjaYJ9I1eS0hL8gEQKspFU5ZAE+TXXcIThHMrzkFFe96ql
5IemgQMirr8zY/oF7dzFPCLd/48vosVplCCXQtxiil+YrYDBpvGtWhC3twoQ
vKwbHvIZ1HYCm0FbFEopHNHiQJm64Jpj5QUFLr1nYXbGCtsTJ1/S8wHpUGsa
7g0n79eoaf5i5WKVNuDw1utejQflvI3qD/JM84zFr1nCCW60zOpQ84d6sVhz
nXzq7c3GkvdZr0cnU+bTZz/OVQdnwccmix+4YLnK1zjaYbEFBWAJPpWnr4Lt
26m6EWA+6PrlsWjCWN80jzdjuX28oxGZ2FaLFYxvNrJTye4ATTDmViaUsGKk
Hy9dtqS15Ew/RdmLSf7d66otn3Bqa1YHOZfPeSk6X6pB4wC/0cex1VLLpFRZ
L1Y64/XKQe1UP7tTP4uIsr8isLTOdYn7IWR8YiPkftYuzijw0X9xbhDNMZ3R
wFDkK7oMryznaqs3V5ZhvN+1Ezy+3qO5masxWPCONp+TSN4357KJz4XptPbR
YfBZvYCf9edkzwyTbnD4XeYoYQHXY8SHI8c/LpLJyRcyljTqinE9Yn4xxhMa
vqWE22B/jdc3EQ7JkMlt7c9oPAuHXg7elD2isGsKJEFWINTSXBgkekGHB1fG
4fvHiWjdrf/U+gLacX1Wl9mt/kP8VCcctPyRcf251HmDkjEDuXpIVCNz859m
rWscSovtBF53yJgvw0wdJTODDigZxKhQgOrkwyarlkvvKdO1LVMX44BeRGJO
wCBl6aK8H1T6oU/LDmcTCKtDEUEt3R8iFG8k9C+1EDvgVUaUYgcOxeOg6qB/
Aax1vmCowU+T52pqwd33GzIqk47SxV6m3EExuOAd/mB35SQRXmVWmSa/iLGY
uQkpCqjK90anRiYdLVvlS57kxgmrIvCErOVZDKpv82iT3CD0Zi9WJvEwvSjE
DmJkH7PHUhmbBqkZglnvM1HuPpf/yAJHZArVYtPoV5it4voaRiU3gm5wVR0h
W7Uo6O8a6rL2704mv/ErQwL4oPHlnBONtA/WmiR2mWgwPx4a9gXjLJtvGuhD
bn7mKHUabPGFfrlQxHWhvj/HDwT2lLVxc0nFgx4caJOqMayoWV7C7xH/TUH7
BgSX4gxBuJmHitYFgJVigJXjBhEbjoNzKxaHZFDGnWcmQk7wHkmQvKkTObZa
Kk4olP77BCo1yJ6cnsnHJrcK5TI/W81O71HxApqwNYXdxnXqd0btWuUnzes5
9l+qrsEnN1V4zsxmQbtetP5UrxZ7ahYYUDIY1iSMVqwPbXsIJr50Vqi+Rc1X
L4lJKUC3DnPmMSzbSzf5UB9U7IA1yujjFDC7J1Q5bq1hHwgP//HFiS5EuMRZ
ipPhgZapQw+YNOoVbnByZk055d7d4XO2mncKypq0yMPYsJ9ifZDP+F5mFaKa
/9WQqvyZPJDl+q9FdZPlEat90XIeQ2YcGaXruPBOtha/HIBYFpwN1wBAJ/Vn
XNA9Phov58lh+c0yyHwtIp24OT7mcZg5g1Z6cNgUyKXKRX7aC9pDu9dy9pYe
ErXroywX1tY23ldv6MGRRdl/+n7e/CtY6tyZSniwam2YuelOr2U3fUl8quCz
+KtV0hyxtzJmnr9QeusryzfUxlUZO2iXPmxtSWcHMJqT+kxtV5s/kg7s9/fo
XC8+GtUb5O05mBefFpRgJqjUYnpidcd++6qz1GSlFP3ANNdeYYRAOYLQVcWl
gILd6s/9S7koMqPTHZSWUPYPyILwLHkpnu4PsbBtvEGCP5UMmgCWofUrjZ3Y
ywf/4vXnQHYfamrLQhI9wP71DyaeVrVbJruVPG7L7K87YH/uKPpm8dxgDkRE
DabCD+iaTjp/ChqZYzzfm7mXimZYXb+PINiVP9qIGWn6PTyMruQTMHRGnl5I
Ou4PXn/dj33En2KPuGlcvx1Zhpdc8wx+nMAr5+mbFuVB2YSMmkVo+Kw+MTls
oakJu8pr9JMOmW8KWL6otNrTu27wNlJYQ+bLAK35mQCpjr7xxGWc4o2bfDS3
6RNHOqnB3uPCHi3ur8pZHNhMiSyJDVEZRXuUzNPZPQdQXSABxZHx5mRYhsdQ
f/0/Uhyi6zef1q7SH0XzUPRO/23BLdQ7XCAAliMg82iLsWFGaYiI/92R7y3n
upW8JFeKdGSQdJ1xpVfA5FCqgIq7OUcdiP6BqrNcuhdaoTNObP7UfUw5rx9D
EMUDRFjMA950nuQQuftgOWeRqDqlgpT3iSoPhpOySXryRIwp9PrUfLW/XW9t
/jLA1OYR2ZNPV56XKZjeKQV9x880AvJRIqfKzMuoN1KSgXOTz924qJ6RD6XB
GM+xa02n35TcOYSYL5Gtxm594AYdXiP7HQbHeDB83by53LOsEHLuUBkWOKdy
yJ0FGeFCX2hn/IpVxtHWvl+XkD7sxWU91YUZa5VGx8URBBHzLw5sUSetZ1Kx
9fGPp4VL9j6qMt7vzInh5PvQhzvqFWq63soDR0Fe/roaEFqS5WB+KldbE3A8
mV0ehVY5iDLfH5O0Sws+d1QFh1jaMHD6Z/a07GnpEo51sZC2YbfWnJ0v941r
VVbbchAuZKwivWeCrlbRbw3bFE88MWShpr+fGX0VwwZwhLtcD8CBKuwLw4LO
XQoV/vVMEm6Zx6rClF0vYzLFpKe9MCxdbgFKwLtdLAQB6FDBQWhNQDa+KHni
hzp8ucZL4PshtgakZ5TgWbZ6Rm5YDJrII6RpfCzGnZFfsHQU6jt6HuY2WB/F
XZobzb6kNsUYxSZ8RZO97VhXngZULMSytG/5z2vM+QY6keT5/2jsb2gO+QiA
L75kLkZzsAC8ZNT9XZ77RoeIdn8Vt1icj9JzPc+6L7TB1HI60ZtDICqSjVc+
Sw3FT1yZf1Dqihq6rIifaRBPqs+/flw8H3x51yETyXEfxFQpBL9swJWmom7j
gC/7nZrAtSEKdntqGc9CwHoNk/J+bxy8IU3aXfwXR6l40Ew8kL4ROkgLMkpP
SG60V8jrYUOBhcyU6mhB81hUSWnagKtDwHofswU0eB6VALmDOb6joncrrDyZ
c294u/itkqj7lu/lwRqFJrVrKD+l4L3IFASlxu0Yhw+IwBk6BDKtjlFwbbcj
TUweEWYXB0AYC0uAKi9UtprArm/xKKMkIyp2kEejsWoR/se9YyH/WkEg4UuI
hWgswQhBodA0Xl921CElRx3GvYMio1GuQ+z3leqOKkrF24fy7u0FriMeLe5z
LsKASVBsmOU76YiEAouvL9z5Wl3C8FGoc1Fp3jyiTlMAasg20omkseS75lJN
UP/jJol4/KdnBCG0Jbnmkdm5yb1eUnABeYle3k5XcgjDrvBjWeewC3V/o/Bm
+72PLPAotv3uflnkvsGlbk2ytbxFcoiUHgAW45xxb+smsJrRdf5h+8j9tcY4
o+zuuDiva380UCCBxKg3xafv+DnZsBew1krtM7J5FSoTpbuuO+VeNJHrYz5l
RXFAL2+BTK+k65Y25vcyCxC8jtTTofBkenun/EXNGgIHnHEMNTuVUOqQZ+7/
TLK+RQZv9Ra+aoE22kdleRWuZ2U2xFoNXNFhdsnUjK8qct8UvRgCoNtLSMYi
EhbRQjtxnA/Or6/yHu245BFYvXWbP/ae3+2hrZwjmvDOS/AS76CUSuHH4hp9
45vwD8YjVtzRWNtyk4B/9cFrhlFLnLXeM9XOm+V0/sUWrQqmpX3J6Jzvt2Dg
8wIUrTyt7LkyNkngxtTeFJoJ1u51Fc+jo6HP6L27CivISgsaGzhdYCOoV7YV
vuTn43duupL3yXJF29eJh/PalCxqwtKEqzhlQty6drx6sX4vjbNfQGbMGmyL
5R1oyRptTgJdr97U7Rw9Etlu4fzAbnjIkJDHp8S234W2BDeI/Z3eti+xw49U
EUHAUP4iohirQs1HFxPqB4Mltvf6ciypJXF/pTTGzIeE5LsgjDP0aPTRfnFL
5IS3jH295+8qV6/TiDQOVERsXA4zSOBZxGuOrqlFMoU10SPZpHAdoxzOhdzw
Iq4ObtLqAW999S4BRCs9FNk809COMPScKxZGabXjiGVhdGbAcWN9SPTspWpA
BLxTnOT4wOWW57IfySo5thDNzcF6yI2z6ipQsySb7Vk1D7GiGOMvrv9OmpKc
SKe9VuiwIBNyYyY8pc7SDlq5wdi0lR9exwYO8qDEHLhfe4D+209AIHNFGpZ7
29irbKHfUzQnfrAcMPFHlIxFb3KZMkUx+t6IvsMLY1FwT+B+0Iqo+DGaK+1J
Yjrds4AwLbUntlYLdMLi0i5Wh+rA3hzLebsveY+/J84e/5wfFRqerMfKHzOy
Ud9OwBZx7Xdtr2XWrUghJtTNpEPqI69tLaPYfcm0BsebBszjT/kYcIbslu1G
nnk/vyzWdrgJQxMZj9rmVqbppWoHezPfjO35KhoN+2zF14MLARB6CaCK/qlz
lEeghquasnz3S75PMr3jn1vYkOoiabkRnfCxoPazVehQzSkcUdE7dg2nWIUW
Ku/lw15Bs8NQF7+/yQ+1DJc5YUsXWYqECLv81AJKd3/GVQT7SfZz3npkNs1X
HhuPq7eNmfWIqLXuzHPuYaC9arJk3FABsjje4fiGBvoNxZWno+VN4lswQl3T
K0lUyI9dnyEdAbEXIWTgKEKwic4tFl20vdRy2RG41Iqqt2jdz9hdTcsir5Au
2gkMQK2mP4k1B0fzQxQp+tn5CmfRF/+yKjMdbuAY/McW41dB/4EVAVJe1zMn
060bz8SmtIzkZJoPnZJ//DJQ+fp9VL44zhE1nHvbgKwpDhoM8uKiQQdrxcmB
uYtiVTYW/UM14ApriFFaBtJJl9Jctl00PlqBw15JjoqOJxLxqyblJuMzuEn+
dWV05oVkd4Qji5MHkt0WQEFS5s5eCWa309lQIBFE/JlWNLAWZqLV/QOQRzHs
l0i0g8760GGdKdn5AUOvVM/z7hdiRi7k6cs90dyWZiO8jOP8zsqcWdsl1UuX
FKfXGgW6CCRZKzdoNMcGrSsM/vkuPh4jyqbK6VNntJskiyfbznA6OKG++w99
lskkSb8W4XjJopRBz9mPfbT+g6ORC0CMX8gIfaXpfXKdA8KtfOBZkxforQpv
4ay9vY7Nra25f217rPkd/CitO8GhtNT0V8NzyjglfVY8VFhlDABkyOcjM/uz
Q+EVoThlZrbpGWdgKZ3m9oLnP7iBQ5DIf5brB3Kh00F/xnsUpG1JkumKrg0U
3RM0nfLcZWdKoXLwT9dV+seBS9O3SFiaPdtny2I/IwU6aaGGKUHwVgL4goiM
ZyBOxdulSoUWMmHqlGFJkJedFORSjr2uKd5IB4taqGLZkf4qSCJeU8CFJIr+
tbouV6Brf6u/Q8sKyDfZDkbJtUm997QgnApwoMQTkCEi01OFDocehsh0WlOX
yUSiD4H593Q8rQE9NGUgxpfJ+vyNNgCqsT++/+bSYYfA3DZctc32mDVcOsKW
rddjh49+5R570LE55l6Yf9lTS0b0lS4a9ARghqhjPIFwzwCXoyVENl1hYsTs
V/auWhoHG3JLw1ZmcXjkm9M//pxx1MLzbQBjkwFRvVndS0mALQLmkYoyAcM/
JXlTbtQgCInUFHU1Co0IkMq0cz9YGGg/vgk2vJKJ1XEVQOPZwL3BJ8x7VVwt
buNGGbr4m72wW3OY1UzJitsW58ewYs8TpPukS+eYQ2Ip7q7jS9tHEeBidVzw
b41TTO1qFLyp28ptVPFmcxUJjWU4WVc9P+2V+lS6UnoDJCiJLgqbiafGnrfZ
EPh8R7F5nM6SMeDixfd+p08qWYzOk7V2Cfl+HFatJcGjfGiT/saqbGqGvYzR
wi89M+ihYycegXPSSiJu1pO7qPinbJdigk2VhV4lByjbvaB7UoHK2v2JezvG
9pGU+AqniPneSJeYQdLGaBYi0wXh13kBqxgL/LGM4+zOGUJD29d8GRqg2Pwz
ULk1Fonfy1fUyvOqYpgZ40qITlYZwox7ZINPO1eSnNCYl1TXXa7I6fMU42rY
ZopmgZpBz9TMz7QY3K4UKKT/bqgwJeTyWTxXzhwybfIYdr/tJTAiARhRBBei
xQNP9xiJLFd6/mgTOvnIrJhh2d0Ujbbnh4pqPjWCAn56ZsqDVFgX8U0kKbre
629ufh2AuwQi0swrOezmA2K68bJ62xy8L8wvBRu2Z/S0wjEX/pXgUFdZf1mB
2ttcTn18Y1AGyFPMzUiC/dkMegAcDAcNC8WqH8FC1s13vRt7KAloobae+R1h
dZEQf6hg9kV0junQ2LIy2svOBQn12pjdvdBB0aWQPKcnYznXGcxTah0z5Gt9
5NgUlfQLu76oP9Omf8jS2O1p3y+ql9c0EL4bky9NDDX/cFISu19LeMuYvHD+
XN38Zsy5mQ3CvZIc1LMiMQby06vh6zCPboF4oGtDNLANjg3OsYBxccWG5l2d
hbQATax5a8gVXnPhY5m+g7oKv4HvdNb+PKcnWeW9E/okxTUApas5OGQ1g+v4
KcRHFxGB13ZfTFDrT/e6eZDnh4WOWx1kCVR69qd6l93R3ZN6FLvATE36Daad
xYZAUdQahNJ9waKPmauPG7HVaCJPylT+lXquzFX2rrsbcR8uQQVsy1zUgHME
jeusL/Q+9xTR56nEFvO++IITgvQiNk+FbYWIX2/p0RvQA1v3huKGod7RftaL
5UHE76vqCljOfe4rrvdGkYt5dLF/wsf/hqR0xIbnWetwk2OQCZN65gm3XqbX
lXJOIsBTCS4cCSJLiczhS2DNSbu60Kx6vfRlb6k5NC0zCKoO70nlOH2HbLaP
ARkKHXjrikWIn2jv9QwUgqHFbhMIVLdk4jUB4Qud6DMKokHkI2wmoibMjltT
i6w03KcmjGPRWKQ8YL1xu31CpGXTjH3Kr5hczq7Ww1SrtsVajmhYLqHCgjZc
IHEVnafIZ3ouS6d95oOBxQNdVkLCbOwcmreuwXutNF2ubKXZxQ58JN1mrDR7
wzQVZvwkBwpacYDX1cXtVBdf0aRtZfFR9/iDKwqmnYq8IAGbORPGWzYBetnM
3gkuSoaf4hN9wM1eDqvl5vSqIP2P6/Z2vkLPLjvCv7PAO83VSJxRR4PTqBe4
NnvIByMQQhbJXFHqcPArJAv2so2LAmvkhSiTNzVe614tvhnHA3MqSkONWQ9Q
PODlwdra5HoE/ptt92Cmrh6OQ58jApvS8R/kFq6l07pmmb0eDaUcfw3jFy8L
cxlNQDTU4TuRXadgkWypJfyFhCDxp6V+ierY6in2TH+qkJIPUh7Alh/QObct
h1FH9H8dUMhSGkJ3yVbXieC4LiNlAKhvT80Qte2+rcY39l9DpfMoLjA1f1f0
2AM2dMFNSQcMdeOxWMo1AHTLr6H/PiL1DZHFYSzlSEyVpGNQdK/LhzHCZGdf
gcx1yOr5aO5dSJaE5i7SxwuVMSFQb6QPqETm0LcntgXn974qfLHj7KpnZjPo
qEoKMFRN0+Or4zMLewc4xlc95xftir98OmvaZ8yxES62+UeTrwfuWTe1y/em
OfEIrbIFKjHfQT0WWLzUWisAmJ1wHB2d0zIlb0QVB6/sG9npIIiUAkwWcPX6
tWL6rjD6rp0iDvwQNODt/nMtB6CRqwUBNneLDwEOyRnnxHi/uYgtOp7hxfO+
HoGt2w6Q887Y+WsHStKcHXWsRE4gldtdxRRbk9NzOdv3pdKmHirCBVq9+Gtg
kk5vOQ83QLPtZcQXWlP3eXwMAH9RGjqOXPZGd+ypW1vWvhH6mRV8IcLGjls0
FcZsyIgaBWRakEFQuFl7ZVUYCfGclYV60SIVBuhlCR8LrpQbqddSYD8o0ss4
meRozE1mxPqlNQP53vfHtIFchLDbepr99wZlYo9kKFoE6SAqEIWu8rv1Ni0C
Mozs1BMe7w2ForgeWp+J8vcgPJnKKqI+21zPKq0ApubIIoSE55vE6Z56KZwZ
t67NHSVdjIFrQiLo1vDn2cvrmiCq4Qe18dYNb1RwsCsvvtT5JNuo+e5Ng/y3
UbG+P2OujizXiqgejxw22qNZ10VvZyrUtMUpHGM5a8/RCXvFhY107QE62UZU
gDs9+dfly10eFBxhGS0S1Q9qWeOxQicRjrA5w70ayowQa5/HE70lhjXj3ifs
xLCI4p/vc/KvClUdEZxWyp60yyhVuCi/u5fDFJalTND9Ti5RqPyDeeAzAARz
8nYlc77zEr0ojMvuktpplM8HP1cMdQnokhilGCl4WIOTgAVZSAVenKmjPwDg
9mNH40lEEQhMALXMswohf/WQv14EbrU2TttRib0wOmXd7vfYQSEzm8X65/GY
UphhA1JFRIcJ/1RnZTxoAVszWeoaAckoRKlb44fwroQKdIZnBp2Fr4V9Ios4
Q+DUJUKYAPKY7T1BGIA92bRE9iq30xmZao0M5Oh2mPqhjB/KQ0QZrrJhZ7zo
exdiBlcHfRX8ARoTKhn+qlJIN7TtKiwovEHUOJ3tWbY7KFUJCjQ9qkLjoLse
xOapqLa4pQ7LYDNgzEeN073b/zn51mDVRuJit+vu7BHwExILHNEB1xqgPB7h
oq+ZzwR2CbftHsmQBcQ4IEq7qmMyz5mxLwPzFe/1yjVZ+xDdyRaAJreoE7nZ
+eWM/WgIQ8pTB7KcI+fg7X9Pwax6bXmr9tg0qMfK+IYalwDImNcc+5C7TwXt
CKIBTOHJy1JrijtBuylP/P7WgEDV4SrYcFVjE5jHLfQAgV2w7rf08DjFm2iz
DKmST5M3N3dMNc2Lub3BLdE/7AwiCdtRmg9MVHkgjGx1KUtDbLmDplDFJ8MG
jRxyp6uKaFA9tnaxidyOAPDFWcJZkiqzZWU1kj4wfqXtMpw1wrBsIED5YpBn
k7cxujk+NEIA9FQlcs9ddCcQmSjzIUium4fmIw7I+0Gjosd3LK3VDT95Rzv/
WIX9ubM1WlryD5QE3W0mRvpAeobLgRp5IxUAPu5kXqDgX7LCpcZwAmnvvFul
i8dSqqUMZb6LfHHn1gwYh3E/tTkEBdicj1Hu4mf9U34RIZ1/StsATXVZWoEm
f0vVD5rhUSbsGUuOrL+AlilZO+nbqvV3OfJ7Q11i2XlAQYGIhBMQVTemCFhs
TaGofVDwRSGFU5geIIKU5LATOWgysXa12E2nomhYyuNJY4Qt7GjYO+AE1V6/
sB+tocfkA9j1Sht5XWs41nen45fr7jbs9OXTB6/RVy4gyCtWNCkP9quQgaBB
KW/LNWgJ9Lcb2cQpqYRvrsgExbS11BvRG+o0pOw/LOvbgVkwoAVl4Tej4F2u
fciR29ISzltrs7OQN2NUTAgdWFtsCLozidLGZTeHUDlJwqq8pcu7uhw4nFQi
2H+iJRzvn0qhTUNM54UkaL+700KvCR5qHD1nycTiN0T+jSxScvtK203vSIJE
xcUpvIww9c5Fzv4Jgo2gRNFt2N8X0S82Bc/crGhhIYRVsMAv+FGMdpzmT6Dy
H54il9oIhchDWacv9ukPIgG341436aU86yzNZm+93BB0oo8Dpz0mel3YQrmW
ulGpauYyv5dQmFEdAh8WJ0YlimTcBb5BfwyTWiwSAxQ0Ixf1+sKLZxKwX2I7
wos2yqwJBH5NpEccgPTx7L6xezrx64r01zrw6bMe4FkDqAzfUDcWjyj4tTrV
OMZdmbDSUTxzu71vndH5q7XKfc6EJxDx27CHYQGHjnnTty7X4HhqI0tzb1XU
VzmfvSvhimuL/X5z3or/QbVrgoaYzRNqGPvmmkKc6K8ulZArR7tpzHuigRGo
YI7/XyZ54ea/blDnbzcpFeIb5tp+65NYFjFgXbIk2fIRrZRMabIdjI5GP+s8
6k+HSiTenAhZMAHpQNbqqNAta1/tFwes91wnp+Zr5CZmDC7JVwSpmAxXw13Q
ZxZp7vc0QF71JaRUADOMKotFMyL8bpDLX4P3qXdHSFt+3j8s8dnOqGh972uB
aq8Y+YyHSaNSByTdiucDCmTQVvqUO5NYL97oo6FW7ZhI9cCz/1F2o1mkntr9
+Y3TD3tLxgknLSLEll+CNJuhXdzDHYE3hskkulrHYL0XWKebeE487YxmywZx
bgUOSB2CXiawV78yl1k777NcQghMEg7hapAQMUlVZ4RGx6kqe1HV7eGQy/rv
+bnOkDCvJ0ljmmHNMwXuRgTC5H8Tl+VmJJFzXob9otsqX/bOXd6OaScS/SeT
ohHUXAIr0bRot1Rmxqc6YwYJEsGocSPnOcn6CBE6AizEMR2m+ZNTi9cMHfNc
Yk4GlMQuGhHehowNe5Xo8SKuSAQr8TX4oyMMh3zx/sMZygQcxqGVwKgyd3CY
PoP4T/TlmLiIsZeqRLM3zrm96E0rep2vvGA5YAxx4H4oFyOkF3g9qUt214FJ
S4aCFNndSMAkWBs+zeuzM/+dVg4lwh7Ww5iw+ydmVsF+KbvH1vZd1M5W4jDq
l30JXGOFfVNP1Z4bgxD6qbqiyuEarrlD4hcBpNyz89EIR/zvSrMJm66y9SGB
xOMEyAmPvBcRSRxlDeZaV5lGMBaU0LAiwm1vEGMgAyWb0IlKFN9v09oAnv6M
xPb9Uw6AapOgUhP2b267UBjfhgLnTVa8DSiVRiR7eVdIqBpsfV9Uu1D6w0fq
4WKaCYHAzVnWJziMQGGwahmBZHjU7FF6FdYOTnGhVMR5WAs+zhsKTsCKZSfA
QsWUTV/LIR16SrUp9LRVXTaAzl+1HNdM1PuCqfCD6AIKFkv06ILIlnSXrzWS
Q/KobqN0V7+AhYHExzRt9f5Pl5TK03v+QZ1SGw4cjrLqBXdZm/w2rzLscrRf
lISCHfyLRRs2UClFGJrnC/UUWFiUx/pYyYRF/LNqRahRLzxuZUphVRdWxPoW
GUVothEeLeTQsWJ55bQlM4CfcdhjnsLS6LETNTAkdxyMl11SeLMLIxQ/Iax7
++piR9Qi0efQUzixfRWzvd5Taj828OPZLn01AKzj9XD8cFPsvV9zjaNuL09x
KvERyNHpSUjdLGmDHv4HZlCe+9ioZ6VynGMYAN+hH6bHmqGBYknDYQRb0BA0
S7Uypmt6faUxt96XYdi5LwgJYJ2oCY7SbUCM8fFSkQ++j8NDt+05BOcIu4pt
e94OO8r9uk5Be5AAXNMzNoVpMtoApp246P+/p6bCp4RYhZO1elh+2uLZvd8k
UeDvOdR3U5wUdtkSCA2i8TCwLA5fJmlbdfkvvaSYq+PL4OodysnCZbps6KtN
eQS8qzx3dlqlLHLiKU/XJFsMd72J6kKEJBpsmXQrRTEk62WvsxKs6vhehjN5
LI9p/AZqeeAnXZdtE3HCqPDIwrX4Cb+N+C/sHSMhm0rxp8mcT3mBkWjzVDZ+
9F8r7QRbC0zb6kvZxyvf/avM4Zhv7otk2tGDlVYGeCVRuNlm3Z9+SWX0erGR
Ms2U1pEVW9rFbs2+wxj9e8I7pxFrhmDcG2qdTda3W4kqRUv4nodhCBuRdhPw
QkULTaBi0ES5IMMcsEUBB0asMPm1463XJPTXdmqOQukk8rLJxcmyPHOaduDm
aKGgJnrPoycG3KhcWY9Aurj3nTPzGVTvDJ2J68Nfo2v6mcm0LB3vOiYL4pwK
+DlOdCpQgBKqe8MjDQoqh/KJF21g7N36epQSOPogpQy4tMPCqhIKEdgc65db
HJneqwMVtiIVN2nggx0OtlW6gUfzEcn7UXSId4hzAqieXwUMdYUIUyuUYaCE
bU2QR1dBN8xmchC4yUJdpj4Wm/dVBmQaGA2jHBmB4f9me+wraUCwpWnhv9O5
flauFaQaaZu/XO2MHog+aCkeXOy+NKS4JqN808STNp6N/MUr0kCfkJ5gPzU5
NuUywxTA0I0Mb7gVyOj72++QVuILeCsVRYenAdZirj/TGY8FLuK2vKfNV+YZ
z747RXgqoecB//W0UcSEyWaihJbBfFqouH6bGXQT79hQLewPZhKM6yCR0vE8
DuM9GEQPWp/NjzBo2g/lCUAOA9oHmlgWtiJw9Mcxixrx2Ej1N/zG6UvW/vY8
ZamaS3LJWyc5/2TjxkUJO8UthzaNqHHbr2/IYdUv8yGHuEfTfOcq5BABIraP
BXgHR21UW8UrLRLM9rejPK2Fq6CIj1jyUFink/0zSjvhNmigzD2ZyGK41FU1
MmGWo6bE+dTkH9hP1T0w+LMn3PmtYtNrz4pt3oG4/zV8oanpH3vTd3Pu+xXb
Ssogf/x66mQ/4mxFR24U1q6Oi6Is/YJQ67LDhvYHF/v06EvCr2NtRfA3LNOX
8877JW7oNrkTJQsr5Mb1WHES4F8wTi1iWQh+J9IGZspRxUXDotId7KBeFF3t
UeDvBhlPV1axNFz9KKMYFl1fhrbSnlC0bePzKh75CWmmuGIGZWUG9gwO4neB
v+WNjZCyWVjshdAAMtIc5eyhQy6u+trj0HLdjJ0lfB12Fk5HHKwQul2g0Lhz
PbpBKXFehXHfRcG8G0UMfmHDeQDaGBFe/gP0HWenCknY3aSuf7BA6OH9yyFV
e7nihCceKL1T/i8WKCoWGR7ws0Nlipk6mE2KHmORAYFCtA6OMTG9jFuSXYY1
XbJ1v93nr8XNnUSN3bU5ArjpgBcwMQrMjY7QDYKQVb6zIDhjTJrKjs833xPW
1EHZKooytrJ/30eVYCD5VZk/qqe9FIkQeNAAg0TGPcl2CB61Z6i9kfTRxFgO
vg1afQOnyqh4781/GAoqDXltn0vCfitgpDGhaufvbrkXqaz9WQZsZuUniMzW
6RC3ACy090ie26HlytMwPBVG9K9C4g0mY/gYVhw1x+MKPSk+FNR9bhuoHUXI
y7UJbq70U25MAAVugCifflnsH9Le5xgFoYhCUnI9kS7XG6efbuXHd6E8fy5R
2TR8WysC221GyjUWdzcrFCsuZGS09YKCCDyYJvXA21YsBneqFfrG0vvt5FQq
ockmGAC8jcQf+4798845Plh2vYd2/N93BX1hB2FMnKfgGcyLhj2HXLzXIQvR
dHrjSex5Uuu0pcJpy1kP3iCQcln7jDKZnyqTzFzrekZJJZZbd6EocXGCkawo
ylnJyOH2ByblW4fRXjoOlT4ACsZ6bZi3umRLueXsbIGisk/PeSMWinBcwVUa
q/q6zfas0/q1f1OyoXAgUs0gNkesMoetPCIHq40YyxW9pXT33M7DmIbctyR1
J830GcmRnzVeRUqem9l0sINCqpDifKW2yygJW4gG0oC1r6JnVLZcMLgbxArs
i3WLlwyrwtqUzIjIY6IhAYTRkANEmH8Hl2hk+H5h+hsAsRa2D6ISDtLaSuub
nmXjP8kM36sUZ1KpzFpSKqWZc64uSm5z21OfcbnkdxT+1pSoH+0guhuLztAt
90PiUYThC1FyZX+Df9rLg0qbsHAEDLqWzhJjUNo61kI99QyfBscWrh2+OdTO
B8c7F2zuQzUnYhHDjf/ewVJoP58L6qXZn5Uf6U/rfUSKn4sKacSjuEBm4W8D
mbetIkeZCFaxJ1B/a154H2/WSkZ2v7nDgk6E2wf5uQ8YVFrfzokqqQWxlcW8
+2EUJWLxAW88nAApFjrlMx2E93qO+hex4aaRE+S5Bb0vD6dgiYvJHcoyth8H
enF9CA/CDGycY7I/JrEQ5AZTTAg31IOKpJoVoFLFN2w4ro3LPLiPsNo3lucZ
gKRzG3iRF2G3zrxBgmKeVv4KnMO16RPjs0iVgYYWhak0pe18TKJnVZlFSBFJ
bNsY9JiGpFpZRfFPaJ0tcq+j2HNd5zvUD2Uvb60uXgJDFZTefna3dmxjBUg2
Ul2GWb7wBHmxwzHy8oWb5hO7G3PMvSOyBwaDPbYt7zbgSl3JrF9SoeDajdVs
S5q2CpTHUWXmoGPWe9RUTY7LxM1sBojLRjJl9gsZA3hW4YylW9G2qXm2/oyI
mk4ARiQVQVxA4gu3LVeC3/LP90YFrCYDCkj+zsZNGC9FwaW1n7A1RyRhl3Cl
JEKW1/u+lgFj+poPtis923vTGUObbg20RuFvipiCcBI7Blh8RIKdZdlbxd7s
fi3Nt/nxmDgGKxxn3gFJ2k0SZtzJE0ZNCSXQMZdy2yyKp7DlZ7KyomBgjmRx
lOKPjTy4b9lHTcQvIZFWwsXa/bZRU2CNadnZViS8hoUZnF2MawklvFxd+KI5
qtqxSQBGlQW2234TaXSzBOoLQjyuhSfY7k/hlL6iAkHNn6LOiBMJHy61Oaae
3Zt8e0nLynByGxhJX8FB1lkKnHNP5HviEf9uO2Jts9zKVOoY/4+cKsX5pbX3
V3oWdIqg4YmOEHBE6E9PdtITxbV9WlLiIVf8GORWgC7eqUhJmPWGVMXKY5cx
jVqe79lGlB/zuV9GOVQ8fV76zCNqyt6inxOiW1yo3nRXkJ8r5YvJbdlNE2pF
UuDI67Z67tBKjZmF9PRIxQ8MhG0aPXavkIQTAkEWDOJfRffaKXGZd0HcoBIW
72/xcusjEtKPd66EkV47rPbgXDO1cOTsClqHkiYtPGzSr4WH1GgyEF0nNgJc
szVILbO6JahvKFKZPL7MYWPQlaqlhHR0U4UzEnYk9WFWkEBOaoezuzKjqr2I
Ipq2C2DCXDraqsWbdV8CmTE0udHPIvGLch4D1NwP1yHq54CTuOpBcg4m9N0u
F9oO7/jJyoWGolcOh8sMQMy4yQ9laqvTtwYDvBAww+HhBMJ88Z81wYhI3Y8a
p9cb76s9BQ62jlp6pG9nKut7ffWBpXRaJBiSYB1fdSjlAy1RmOAfJtY6iEir
nBmjg/TyuIx5iumfTsXVOekxVLNb0rauKZR9Vk583RsYoqL/+8+WeolBfPqx
ke1m2907R7hzeybpgF3f4KnHPHHf5hT5WVxxG/KHWafi+I2+iEhaXS2ll3y9
473XFID/fP48XBrAW2syARlWL8lJ1MzPoX37RNQ4oI2JWPJHGAFUphvh6Acc
pJ9Gv7/32p8EG+vWHIm4+BYeXLYKC/EiPsJhZ8RKQvJQSAqf0riE3fyuSy7T
uGI16vjRPhdpfJKeooAzYXgKDmfi37Hj14hxb01s4v/gogF+Vx7uAfQZv5nn
GAWHWJlH81c5kw6HwGSUEGSRhupmjSClR65Wt/eny5V+MqcGr/51wc114A+v
OYYCXc4lEc47zrJ4Od474fiI0Ul19VE/84SpnWhy8O4TjMDYDUP1R5kZ+VlO
7QGhzDiyfdZFtxws8g3+qQzx3JxDOcAtLh/mMXAFO+m31yU3zwUAFI0It8w8
Pt2EMok5x7NxusUYDUWn6AMgUvtwRo1YhSZtSoRmvmr1tMDw0KX9j2ceuixD
V4tnO652edJ/Gf6+9auoCzke3E1Zo3GfsJU8jiCkG/0jeC6RU6qZqDMQX1zR
FtnSs+33plUeurDgoYo5g9Yn71Wn2/ReK5+sv1Rl4dfv31HBojdQYl/XKo6p
7sQYrVyQkB/C3MxbCvE4qeBA0A95ZaFPs/aXsAz6SMC2VjZDd65c3koCWiE/
SCu5RziYwtIg+EyLE4i/oS/jUGGBVLfgUmVGxLS2fZMlmDaJWt0UnxaZld7C
naIp0QHjl1FamFsDRvLqR12YGo7rOVsyN4axig7b5P9JDW/OELJDS/Beyl3D
sqWopZSIt4blgtL+wNY8UjGDne5cA6idsNap5boG18VBPNvVWggcooAi257r
c4rRfApSOmu2llvhgqSnWJmNK6VwLJvHc2W2wBNjSgD12tPHB2Ekwci1R3J9
lGIY+giloUIHj14XWusq0TunMaieXnkNnGYZ+R9uwcTmj0kNq6tQGEYYS1Fn
DYInuDNLTXRFmbWiZQG/i54F6SWOEyXw+kMUkIYwJzLOUkuN+PrJcs51hZaV
SWIV50rbycXAypjbSGXwqyoVfnugivNZElbjrwNdOJ+L2GZZMxB/MGw7XVUV
ZPcigsefmHDN4qPVLGfsjkSge7hB16si2nIzNJSQDy7QFoc70rGtrPqxgtro
zgw1Q7wuWO3WA3KuUfz7d1sqkEj8QUIPTByZOlBX8RRYxL9MY15+80+A5Ylm
IE3x8Kw3+j7xsY+fOe45VBMTwCPg/QC6LZcUK8ZbIxRLLmgx+KK8SdG4h5Dl
6pLfBNDXACXdoDZDSv6fNsF6iAvY9wdBsCkw4ZKmPZ//4tEzYsuA2WdpA475
TssDL7AFCwmeobaOW9//RdaXaXo0HorV0wkplNpkA/mpTSsxm0iHK+kBDikA
xAHQpRlKifqNBjz/tYB1jE/6RKRIjIqnNRYe0HOAffkKWfTb8jM0gbseKHHo
XAsxNW1HBYeOdXrx550KKmaNIzywlvP2N4RGtZRW1QasBlFuieO/E/ooTn0Q
ujAldd+B4OvIHKrzqcoJTPX43yFWaH8DVkU4m3DhUKbGojuGpMTcFbUC4HmQ
CJ0qJ8y1mAy1AFbSXY+pFy25DjG1JTEvUeEu0y2ntVfVUB7Nb+V50hhTxWZL
a+ynx0byQ4p/06hpJUzUEuusfHU821ZySEQQ42mwt2SgUZ3+PmeV8iwvMOEq
bwOeC9H3tDMjRNbuSLq3yfgEdz0pvUYRBoMT3iyayZ05UDQEPGv+airDyPZv
Z/F5o7I+4eS8LKT2qIj1hfPwdASzyk4G14R3AyBE1/A/18YMxdQZ7RDLuo4q
OMnyHIswIz0KtJGVh2H67DaFB9pIFHLxmNdTJJCFQhKzKSSPvR8c92Ehkz4U
zGyCJaw/iLyFRpSfOZX9QcbTA3IQkrBsc0HTlUz4tLyR084LvCWHW1KrRPL2
iUqzpaX1Pk2bxYOnZvwpuTiM1ebw23HXvmnklJLc/+E1G2uHgyjgKnHEu/9g
7yNC/ngEUZOjmf+zYYPFKxMWeP5BGB3hKnZETUjps1V1Fhn+p8qWI9J8Bo46
PqHgF0J1ZYT80miH7QfFQ7pVIpqXf5kYC8+uS/1nIr4MXVuMlRTxbVFYjE6o
KckKsku+GgBzIjPKQ8B1f7BHyiY8mgr4fOPJwI6tqf87i4fsNhKuQpUpSMjf
hWBme5bjgaAdlCxdaFIKTby6QDrJ1hQaGy++j6iHz4MSIJfSTue/fw5PRLEB
PZ4R4qPfKfC7A163pGUwbf/94hABpegiFYNnGL9F4Q/NZ9PnTF7TkhHeJuIj
NiAXL3ww7MnKROPcY577DBXj+IOyVTqKcwWqSTUzDuLmo/M+KwJf98o9gzV2
Sih0sK0jX4dlfUpTpAlxBnXpt/EtUrUHjjraOYIMTJxHqk/8ALpkuianudyk
G8cIjQIqAxVdc5FKqRYRJCM33avIa7SGGl0JeuO6++uJh2GWVVCrSAGVKhQR
+hwi/rAecY0tXflRWE2JP7gNDXacUvVGw+cJP/KGHLzSOD/IBvXSAxPgt4le
1iYJxirozVhd4wgzHNLVbNPrJp+XWfIqUZG+ffN0xmRPNgArbjjIK73V0uv8
FDlgU6INQxbRTWSyCrkuFlWKMsdtXkJl4WhtcHPZDh8Vz3sfeOYQQpaIYPQk
7kyp5Pw2mRptp7b2kSdu41sMbk369Ku7eTDzW5cUOMa18JRvOjTRROadlqbm
II612wj4Ne6ONkJ+JNxPqSHPZ1X1sGEn1CuWvtVAwHXVd48Hq27RcDxqx70x
WxHE2ZlWav7d89f+taIAB12PAyZwOrQ7U1r5HXuWZg8P9NOk85vE+WEsjs7Z
hiusA03/y6vEItKFVMCJZoD2O0rnSnHqLI+W5CVUBMUS28rRSUnCBu8MFfR6
mySg6S3utMgsYnLrresEPJKON+dd0yNOtkfCB2rnI9m2Uu1qQhJ2KNUf+INe
pNaPznQ8evImBKrSSjR8jamu1YrXIIxx9JrAibiVKFq0cpFUdI4GB78bp5Lu
qzuqhf20HPnTJqNOM+JUg8T3ZzsHF/B7LFfKJ2Oak5sCJmnZrMQNxQ3kR2q+
tGoEbLxT/i+p3goBOw5iwVlK2DpF+YFBo6LJ2DiNeHvgU6nI9RnaUp9DWo0t
1aYM+D9YHpahF/lqWB9nacagyAE1DQOVLdyqkZ9EwR04EueWNFM5gaG2CKAX
829dRX9colZvYX8Yx1k6ZS3DrMMxGhcJl+/uLOzETwD6OIsXdc7WbPiJkESg
UolVh3sgU8s9nBk1upgoXfUJB9IMcA7Y0Pp8I2oT79BYxyY0gSQ3g3uknvtJ
s3dDsYyL+3NXb9ye+TOggJYiinGH54cXJpSUp5XPbfDqE/mg06EGf6JIOeEK
WKhln22uADrvvrEiqjaBS+AZkWqh0uRadh2n3wFC49eyMONXZO8FyvQ1da6P
TCeqHzGO4yu2dBOaUNqHxewvte44knMoCD+6Hhr/kJCgMPd01TVJmeGKiRkx
gsUIFJVRJjPPw4wc2iT2LzCXHUEWXUgghAEj4jhcW1781lZwpUT02bELXhqn
xxjBtbCRlEJpy7Q7lQtZ6UHU6Hpz/QNrslxRWr9EXRaJPZ/rw1DLCFsjhPc6
+PjODOwg01uhQfPQLa9uzz9V/MJ1yrd96nHE1Jo2Md/US41QX6Z/hRHeEwWT
cMsZxCd7K3VRIi02e4IZF/HtD3XS4t6N6dhCqOfyAtPNIfJv83bmdDJ1atui
u0iRdN7gNCY5EcZmt36b34oKnRilCaied4MKeWKY7lg2ADC3btk+GtdQkxVY
D9ZiyHBnC8UYp4aPpsJ6Kv/fEwV/Qy+yvP/LCHbfPyEzgi6XDYFHFv3z3qCE
dvwJyedzOcdnoBgRVs/y519EtvAgmQBJPN3ny6XjC6bwSKU0eupPqs/R24u2
1w1e2Jm1Sl7tzAfyQn0gufT5Ig6DftYKHi0Gbz8VpFs3uWUTgU+ARKp5LhWm
yajeSWm3EXH9uAHXubBfibXqydTfVW2wi2L9i9VFN9sJSWedYiSXBW5Rr+iT
PGr8oXl89XPHMMGvSC3+ueNJogrFgkg+1uyJLCwnofDZbwd7KBw8bL5I5MU2
ZmEhVYPFfbkUG8KH3+YQYVL6TYljYoyjxzjRxd42Wdxofq+RlJheXCYaCBTX
RKEnUt48XY5/ccRt00tOU9k/1kr4qWOUnG0Ucrdkm9MwNkoYNyGzjB8OhXV2
r2qbBvrdXHYMtmZd8WZrvQk6/OdtSuTaOFOo+GlIdloCVz+fGMJAkB7o25bE
ZoyYQ+cwsb36T1voXdm7gPCO2vpbCW4Dy2TXN6gBkOAg3DX7fFzLSoFBPUnK
KqjdoupFG3MsqCFwv1ksS3eI6rT30261ERu5Xfql95vKhYBeIM7Ou1mJ1C/H
viwSAY7pZQt1b32V5VzGfV+Bs3F/+7o3umN7xoD85/gcd7SzNza70jpjvJpQ
c0GRxO8Btj06ClAe6jQDMmscvHLJyyzSLe82mYW8avrpjyJABClaoDsAbKOY
EQejM6Jp+mcCh5KXrH9T/eCR212DdE3bX0p/siqokLjZVKEvf04ygeQX5B7k
uK+6QkYalVL0aXrJVao/JX2ToZzYo3RaAyPSeKpZtADLSD8mQ/uNwxWfse8o
x/MxfMMx3d7toZ/XePJ7P+pg8hydsmTihL9mxRJ/2aUWtZWnAT37UkPRnTdO
cFW56CrSJ8zVavqL1fqQVZf0SwjLhlWGZ48+3yGDOJ4OofxOhlsFioHegkLe
taf0984xNUj1APCqgLlLzaFMkbwfuxn9v+TfW/T9Ye/fweK36OmGLER265W/
OPNDZG2lgaCZxihJwneXY0nNTcfzjC1NuahJWwWg2cfpHQiU/1B3svijoFoR
e5VNrOpSELu9UZRx9c2XryH5cXW8Zg5QBUCHGOFWNcsjNPETN9TiE0a2ruH2
rQC/CyUYpSEoFeC4Gwqasu5fsPEqZbS/ktTzKKpGNAJCEj+ZWhIVQPpTMkZe
reZvz7EnL48xbD+Uz+FZlFgxO1S1LA5mX3YZF2Hxqa+p0AgyErlu5WHZGXvB
yX4ZSIb+z53SBFTs3qQ3ShQe+L2mvew4LhWuDJ5CoDlh/i09Hbz2l7I02g+z
M5FLHTK5O5mekWJ+Ef7sNgDDqye+uy/SD+qx0Qze21B+nD0M+pPnwSznT/Iu
jdiF5xtGZqSjT9eXwaBXCjsMKYoTXKuBKKsjUSnr2QNIC+xF4G/Jnyr5rg3n
tMAda9V0xcB5Uxph1idzZv/K8gkDbF47IF2RgZuULSFKWTl9qGdz0RF3GEDE
qhxDA/Ia1nxQM2JjDyjoXHBa6dIHYX3Aw/ODWLPv8HKDB+zRIKHPmd5+dTgr
NNB9t3wqhtm0b+913rq3+fDZrIAECUZ37nN9lggN5hwfahzZ5PtV04CQSGvw
IIXMAt352tWUqVCBg3eWIASYKvajCrLZ9RSZV9XkcCA3HS9tLox+W7xkxLQt
gdUmfoKlTwp6D0LraMpe4pqTOhEo73bIiZXdG+5NzemVSrDC/mQ8YNW4QIgo
KSgdFbyb9SoLpuWSZ+SuCRbY2Z0J4e6GvMZMy2v6NAACBIjSYR4jZs1WXTDZ
hiMk+TqLkkKqyhjeZvoqYh7VpklRIksAMHBKAyUw8/oV5/66QgMnIjFqMwR6
PSmdFb6uBO5oRLLJj9PIJqgQG81nAAHlWU/KTG9YkAiy+faDlKVweKZXLsRN
dvNpUPRdEEifvv7NyxBY9W40k3IQHq/E1900M6+6mFDnkvlHNTynJGepgZsu
rWBrQtsPt/2ogIaMDJmKy5i2EUfhzSZzOicKxt0AES3ZeiPpSp5xCWfhCi80
8P+xK2NLEnx+yBNC/zdQGK9E8rLsGpNe8MiEpP3FN4Euk/iEJLef2Ggfxeta
d6/ZhsTI8GW33kqEhgZD8/PgI39fM+3idGW+7ifBV8NpAUm4TXF1MCFrGn+M
PH5HIR0RiiwnA502E+cfWYIsKhF0XxmhCkrg/BTc0vx/SEh+bGN6EA+006J7
BkXxVD7qjV1D3O1HG1q9VuX6XBWBQku0ipCcKGtZ2p+vOYuH9F7+kmY1q4qQ
ZArDCXQi5QALuq3lP6rNuGlVyt+jfQVSuKpMKW/Xh+A2ii2/oT6zezWn/q0k
ARdg5YlFH/1Rz1fft6qbNJWWy+UGwecC1gpzih+VmuZEMUIbR0dP1+1/luJm
boz3RSToTaewx9CKagiHGKzu6vKiCvOI6U7WO2bzRRGOUBrxPVEYtMNc+LG4
+YGOy7YSOwq7YOW5D4OiB7XSv85V+5tpE8y80/jhpyMrBhY45+CMK+Vkr95e
MVKS2vVsm48vVrlbGaDqe+lMNHt/5DQM7wnaqNfOqM+UiJB2Ns1GCKX9tHc0
Z/kZQN31bRxQW4SG4RAq4Ie+RJPc2R4ARpru5Q7ulppQ+ufWXiab0r1iHD2N
I0f9Yro6SrfSBA+r2R4z0HPhRixXxdS8lqtj76yZokdd8mHeWJv/i9AKWDNH
O8FFUPNm829/QNarQW//27L6EsOSZvxHeRtjuIt4OYqmKw3jWLONmiM5CIj1
Yb9IJtyC9KwFObixL5Veewy6DwG2iWkhfNZH4dHYxj9NowTyXD+XyWHc+vku
HzHVcFs7O8DlZybGyEbmE+9Y/KBgXG46AXv8KvYnMmSEz/p/Kjay+pj28TF4
Xboi7mELQAANVOujiuWmgdkoBwy7BqeXcbrzobSsU9l3RW7D145MNJNWb3H0
1JCzKWVSlyXMYiYihHmkycaY30pOrQJoJbJpSULjsCw2XpPjNaN/aFaKmmIw
8oXLQDgu/+mIMB1gsW2eur3iJ5Nep8uej+Sh6bEvjU2Pfs5Ts4DCJ1fADWq/
A0o03sua/4BMITNCznTEeh6NVFqAgjrBWreZ3jVANkFdj0y6VRAmrNEHto/P
caxE5/GrUDwrQ9BvEL28LnhE0Rckb7uQqYfVZ3+qK66nj72GZi3DnTkTxcO7
JE2S3ZyJuZQuYUndrHq+qZvkjVIPlY9EDRwkxnn4m641Ea3GFUswBr4QGG6n
nLoIaqbfYoHGyf0D9GDe4TXDQXY2kb3AhgRQprrhzrwrBAaIrrIQFr3PQHZu
c7Sy6XmpO8IBEAp/p3rQNJdBQW1T9xKBUxJ+x/WEE4ssuCvFOJdSEJkjl18R
jSziaTqb8WJzOJSaNTgrsvrxenNaWBBuJFqfGxmBwTHAd0GB4jwi1TNbWIh7
VAJIV4+4gXn0ON9AyyF3P8H/pvKfulHIdTxRcazrV5E5uoCNWupMoTij4VfO
LBmnlUcUQJmf+//yXwLzndowd1ZJ+WQJ1QRh7EmC+Qc0WZXd5JLAMHveRvqa
xbyFYO+PrsiTICk6+wGLha1vN7kV+SHh9EpTHASUQsvrP+mE08FQqQbG2mr4
sHGQrSUW8VpcO9+ddTYteBxmehXIYFNbMZpxGAJTSQsZNowmhw7fvn3QmC1r
xyLmlRBT0biee5lnbGAaF65Ix41CNm7obu5yaDoa9BiArzEcXolHwfm6yzY7
CiZZkXuoLKmtAUp5dY+fYV0cmS3u5EsXGIpcKjpV3R3CAiB9StZYe1XpTEue
ioi7gNppYMdVsqNFWt8gx7BdP0jB3DpdzeOScD8SiZwVjxW8rLTqNBphsbbH
HJt9L36okr/Ay9EGVLZZ3cQ5+gVbY2PN0831DUI5f/Q8Zu2LAKUbzRmm0TpY
YvtURzARdd9iULBmGajbRnygjpexvUvpDp4OKr9zHl7adNcTaIpZ/BGX7Ft+
ZYgfJeJslwFwnJHpwD4+TWOzvb5d9eLkdzcqGZ0sjsjeEHHm/IZtkHP+d8HP
vH7pl1uZ5y/YGSij9knAw/Xu6HcfEfldQs3WXZUERPHXyCcuEKE17lgmi0UW
myDIOYujun2leCMxkM0E/u7fkVB4B5cifpYrYB7RRj9eJZuYsc1LFPTMOkOk
wEoKddJbba5cJLPK7bx6UsEEr1AUmiTMSARWyxMRhfXVPXjZKFIzDeJyzGxB
QzuXw2anMoTcLAZmklaIcWTdFj3+ADBLhJQCZKA29Zm08PE2c/a1WqxMmt6r
TsLLiBSE36ResdmB63ElQHVoeooLK0MIPFGUIvTr4GeCBJ9u5UxyqpTH9pKj
f9qWEEmB+k/c2kqPRL8Qj5BQzVUfJ+Pdb1hHYEVRTlufPwHR3EhN7RxJTfM8
y3NJ9PsjEUtAGAIq9738Muc2MdBtOMN4UFTB80sButjFfknvzrXqvHHqJMCX
pyrs3AltuqOljVmTa3+GlAXCoQL5BCa8/hfsXZQFg/xfkhJjp/OOHs0QZOoM
n2HMtMEqTt0GGXJqoXie18GJWyPRqri0QIxADhMGoY3CtlHSnXjTBYKgRqCG
26mhIDd1JfxEoHPEARlafSRzu/OfG8Lkuk8yGd8pToN9L/NfIdRYvp8OhYAQ
JQASGHaE9emXdzfy1PRBe4c7D9mOHoMvwsE+mvWRZjGwtOQjWWuNt0sFEG6J
/iNvEGUzHJkaOcF2oAor8IsWSns+AO5KKtqCYYbdva+M7JhEIuvYXwZdPaA3
/B/EkYMIInGFq+fwShm50WY0kvA3xVGjpE0NEolFAIj00lxHxreaPz/0qepY
voIdijcpHNVPs6dJah5ffSLg/OWjZW1rbmMIUcTdAs0NqDSzc8loQloyPLPP
HUgwGR9SWeX9Cl4nvxmipU2Iuc2SkGAtvbYetlHVPitiVXMkv6mGxtlki/g7
Y3EUm2X+b1qLLz2G8+5WudP8RbDStpBOoj7JLr7V0GNgzIoMnQfILh75bkHr
A3H1dmgDRElWkwHwqOmEaqFrnsliLdcxKqP2JYLh+oxpA5SNk5OrcEJTfoGt
2YkSclxdqHWbfkUbESU73gJtU6EdM7ejwZP+feIkZslKG/aYM4o3PBX15nL5
A0vdfcefDNSMYNoMLdVbpw2ZzKzhk+9PCf0QOU6PZXptWCYtpu/LSzmsJcXc
yaRbfEFganELtHp1ft9TXGf9NtkP6HP4upPZOHXm61hz4/1xJ0tK/DonDy2g
tDFsctoZfDUFnaH6sJAGXhbiHkrZPvtMN8WyhCCcjH8ayVShE0hRIBosjEQ3
/el915WnwCsVbVge61S9RAE6GNWhGVetSNSgyjgslqA60BlBErs5XG2y4Ulz
311JaNQAz14xQREYNeJ1gYVN01IRD361NJLKAGAiQwgugQeJpnb7IC61+3F1
6RibXZV0eXHv5AyiGRUjJatRkNEaILPwzXZ8rgprTGQ6iQytsbsB7OCEgFi7
nKb0kMYhtGPtZ48/H2ATigBW2uibceePb8RhRtfV8BHyzuflh7k8Qape1B1v
8lFLwfLLYKRRMedPx3MMOBYLX0nEwCNI1IDDMUwqubCxZP4S+BLELAtGIRLD
OrUaRN3HSj866sjF0xhBSz6IgXA1aiO93Px2HwSkZr8x3oyUHJA2I2aA/ZDd
WrHcymon39THMs6j26ws7QSrZe7I9tZ1hGW84//OcPPxrqlb4GLeAFlz9JC5
7rgp0hpEESdbiqAhOcFX8k2ckRkxanBJ82MmBoamhkSAOLEl+L8Mihhf0PQr
fgiDcUfL/malY/WPODiQ6mYIE/SqAQZm057fihze/chOEklZPaKmZ6HUYQ9A
GgMcYphAE8PEdfMKEH7VOrzTWd+N/zuDY4/hcgiD9xoUynNGO/z9DMtIT6g8
bv6yBuQZy6F+MTxTPBTGl9J7ChE8mS5//tcxOeMiKeuLPu0Gs5NuoqQqjvN1
p9PKeSwxMua37wL0eB9rzQcz72b3stp6i+LajoYMEkKkYzvBAIk2ANNYNiFd
9FphsZGvKu2uzRrPcss1LoY0U+UjhXcW+9dHBW07yJYz6hHq4TApHaZ66JhF
7xjGXC+xognzBp/ko0LYTOa8Nr4tbcRzBbB1I6AT7Uq4lI90L7vXdfw6IxVI
fqtJCR/kOoSPjufLN1pwO7363dSWbj/Z1rC5p++h+pQzmobZ+n+YdpO024zm
D9y00KLH45xg3OyEk+gJTCOMvK06OWp24GY6AsaKKhsCvRxkWMz/plWUOUDF
FGqOoZlxs9n1T1tJhZNhg/lPV8KXIhjygSTrmKunUv0EhdbEFrgtiuxyDJr0
Hg9vlt8u7thwFYUImcw1zkqxiy6VytCu9oQSqwXNGi1FHxrjzTC2GpXRj/5w
ib2P3e+np6lNG44TCRPNqIIKTYsipvSls5U73vOJEc6F759FTbG9V/+gywfd
Aio38793Q5DkbVPIAbTPD0vYaL8xvb0tTqQNsb3ebhq3xqO0EtZ5s54orUvV
lyskJaNaoIkxZBbtZLoFMLlvuW1pMZwQQMTllJE4Nv0NWayPlIn9nhEvajQF
ZVilzCaECFSi3v0Lebx67PnXv3K8RnFtVkPvzWY2TsexxrIRPRhI+WJbavUS
wiRzD0R7/t8P/eXvwSgULO6cKuT6KEMMjIVDmCGDthl5PlFfjWAL61GOSUS4
VABPjPAw4l+tVQjUAqK6Z47REOitLrwhzqxIKG01I6Ky7Zz5gHCdKGAGeM2e
YQyTwK0IE6JwkMygK5BII9OC0DBZXoVLT7vWV6gSL0jMlo4tkOwZ/C1Vukbq
lrkV2lML098Xdk8TCc2uA33qVRNiw5A7B11rfSmje+lHF8b6RUOS6NLe3j1u
q9ZiUVABbDp9na36bjMETN8ewLtE1gbv0jJRDruoC/DoZtNBi/NqQLljU1rY
FOWUH3zEpTlAUXHaWSkToj/cz4iu/HUFAUmAMG75o1UtUBeyCdXqcaVeactD
utUEFTjryZPLAfXJtimO0ERHqpvudj3/z4XCbd0BNyl6KyGl0kM552X6WXoL
J7BHayWqQfbb6amV3DoaQoAMn0XHJK2LMqVDiWYoQII03i2UyhUqwhc8ICHK
jqN5cHeZk1cFztYFlcH0omsmuq5KPWF5Uqbp8dHlaTCOIr03fezLfDfR0csU
rCETW7Eq+LCDst6yfEzEDoyVnLO6OpuR53HJ/WwH/IVnq5mjmd9JQpdUITc9
/nuxjcYYYoKSbi/ElpHiJu1Lnwk0s4J0qTqQ94/BIE9z8opk+BR9UkBh33Hi
JZudHdLBfGTtwNE6awN9vDZCO/MMeXSSd34u9rLO82AoHaAeGc22y3X44gxs
w4i53/IcL3fAfyPiSUkUUSt7UG+vaF4xS7gOr/nze8+hOCt3volmGYkkARcp
HB3HxK7pHJerDUxDfMEmwvLfzq9KnFQFVE21XFZRq76D/79p1fsiMTlntfac
mh+L2QHTNwcMnvCAMGaVnkyhtWQ9CMutTfdJKr1pt+Lr3d7CFgJc/PxyH08W
0WqXyQuVlRsJYAmxMDxeZytRAPa0NENY8Npuan/9CY7t5ruBMty60gstrCFG
+JG2qFUfHUeuE9ydDwblLFt5HLCcMeQvoLX2wx/0EYieGyK6RK2HKV6H544j
rtbHqWsS6w0izs4fz/ONvelZ2KBE7dYhtlwbYCb0JbNS+sGexUXebyWDHnCr
3l3H/VlnMv93P7aATKs6lP2gorHGWtNsWqAppXrT8vTY4hP5teRoq957soSj
5qu67HVYAM8VLLc4J0Jygnxol1HKGnrJjULgebyIRI5JhTE6o/wegFE9jo8I
3Ei+pNLxGtslKAUk4pFxltVj5C6gin6PCR7QTX4DVExPcd2/yIFmmijpAnaK
kma8HMb3ysGn+lBV79YBEcWGEIWC414W8iLHJt2jjG9iJWj5ACPxxk1391Mm
auYKZpNet2DTC/htbjK6FNXDPVyKJbDquR4yGIkpNmH/pa9+lNQg20gpCxcA
PbxbqmKXyhdAmD0H/UQLmzWENhQh7p1jqksk72CxvumvNkPZfp98ply3p0ra
GOAKaToTe9GcWCay1xX4I2ulxkoxt4ONCnkMRJh6YeQFZ3iYL4bsPbgUbx4J
EKN81YCe8qxeB8rtINU2CEhOyGK1qxWZRZ6YgqSReSITj2kZHzkF0CsiELPL
kwWAESxYS0tdVQ9uxP4kzad86pvhXKS53IloPaMkgf87Y9+qFmK/6alLYYy5
mmkAY/9Ls/iIojipb8lFJUyNfWpahHr2F0ZGpXWfKXPMHfEOUCHxec98yBIl
UYM4us33o4SRgNYRqk3YsKlenH7aaSD4JUU+UixFvFlYNKpvw8lovPwfhDCw
J91UucPgh5ocAfvhcxGZOSOJgvjsczOkdXgyFhkwWxNrQNjHuWB0fYpMZQHB
Co4qMvC7JUdPmHZFpBa9ONvF6P+RvCCvcN0OdW8Pes827V4KrtUgyZzRg/T5
zzNKt6O6rmIEi5aLh9Lly/vSGNyb52kxjxcNMODz7HRJbcpeiXIlcKG6nQlr
+un3PJmMt6tEwWX3Jo6/3EeIfwDBOOYhK3/Nz9UKeNalWwqV2q3WV5pTTXsi
BzB5IyrxhtUhprtE+RLL3ZOT8OAq9ERU5g1sGIyJiPkZQFKw5HrDwIIORses
dv+SQv3cMhTpi4/11r9I71ezdRiPnpAZcw2Me2CT40myxKdGLCkKwlDZBr2s
LgNpgxrzB6x6pEPz9MaRM690B3MfYKwNKtsMBGQMQYldCSbjwapfjTvXnrdN
3brt29H4XLU4CMuYd/kPzJQ8gJ7ZbTjy3q3kIO70RHZlBSHmhlAG2BFyeKeX
N8+3IBtBZf902aJ4auucNgHEJCxwC92lVn5FZU4Du3tTF1e4eEeAqhKW+vTV
8wM5jPtkbqmrRp9P7y4WgJm2Uca9m+Qtdio8PSOTyRmd9/JHYabsATJfkI7x
wND7XBCJLySuAi1HbfkLfrv8BqlLkQhlccfMFFNcIiPQK5oOvIpNYa7BkLMy
9AROu8cwIWQsB3ouz+eSUOZohYhE82hIrGR7v5dSv2iqbg1PqjswKt9vZ8F2
zj+sg0PFXdFgT1fy3rJkwOSAiCiv5VJsJUII43q5zfp0bco0pX64ZOWWKnMX
mRdDlg3sNXMomOJKWRffEYD1HKiWFJKlEKkkWlWUOVJNR1+rEj0sYg9X0uZT
f4JBZvIVV9SXTDgOrHfz/GdxCeCv3RQBN6PoB21aQpv2mAIdQ61AwS7KnfYu
fwIlciaTDvLBegPW7PoF9eV9Pu3m3bxnIthBECfqAtmWPQDjDWMAfSROTYbj
4TmZAAHUP7GO78g7keziE2C1gQ+E9nARfLD67qDKjJQ9rUbP95TqEzRYP5Xy
nSP/9JwzMFQKMrSEFuWYHXtssYq4TpcP4sqExFdC+v78qS51o08WbbGwzsbo
LVYSPb2mv91h80xBvoCOWi3AVu/U5EaMOGipbpB5ddBUQiHgpQ/mi+6TTwvi
yTmCSUXESa4mWZUWrspBpEdhKZRenrw6a9+o6CZmtQ0yVc3+xkzDm5DfJTN7
xLz+p3cs8TFkUbpIgczANKjFE6gTQPIp8BWTLqc92lUEmht0iGBrSCaa4A6k
UQiKpqC+XEJiM0xTeaClly8vtZnkOb1yS5n21wd6j3yGqWdVhY31vS/eXcyt
lxLb+MRODBwKpbr+zYpwzcOr2WmqIPq5WoqoPa6TCLK9AsRWswHVpWccBYn1
X4Y/exh+2uD167UshYvrVeRC7xgM4yMx+v3RaqAlZi6hfH15Fg+FOupFn/wC
qNM1kXdNhcuXMtEMjs5uKJ7FnP0tzYjYnMrujNDj1FZ+GPEholxmLR9XZ63B
vIyP77BevsXAkCBlZ9RSy/sDixfgVwCSR7aw/4Lv91GQZzi0kaJd4uhxgn0c
Ou+f/5Y90xQ5UQVwL5yhTB7kTtKGKRJZQMtdn4EnBgeGRnYXRLJ+7X7Y51Uv
sX38CL7QPSGsUPRuBV7uhc19IhcNhCmmeeHZIpLHzJ0llWPVNIarRQOnjhQe
c3ZjT4UtacBWK+XifaeeSQYnTrdCRU0O3jhXT5vfuABAJtVKTaXaN6NReRP9
0XMhgi0as8qfie0otZ3wXWJmTzKbWD89lRgGwEoW6jJgV3DYf2dPOEDjImsY
5kqHn7ADzb9cfZfXWtAo1ifLm5AfaAWawW2fS+rdcVmWtvv8qmzUfwionbRE
DDuae92S7Uh27WCr9CLq0zkgLuqNiMXm6xrVVEx2q26l2St8g43GlUuo12QZ
GzmYuSIPzNvchse1XwjIaRffPONn4tf6lKDhbnRw7MSDSUyZQFWw277Lhx9W
gB9mBmyAUl/L6BCFS4hmezy67UnkxlGnDKDxXfoxXldPzg1SndI+UQLPNqGm
+D6zvXeAvTbzfTzZKSgZubiIiUPu69BZzQkediPMRapk5clAaV5u+4uyyLY3
wapc4jBdE3WyJ01BKpP5F4BcnmWrNZAn8eTDIDIPzn9DtRC2IjC5+mdYgnW4
d2ZDtSd6m5fTDorGJRGUFDniTHHYO01OJfasuv2v2QVSFJ0Xf7WKteabz5HY
gIvJ95pR5Uhki3PLuViXomRSNmeks22kqDcZw7mOm8zqampWTeVj64syqUhF
CXunEJ5xGnKAOcBauJPzHCLnykg7s4zY8Td1gyP2jc1zpDKEN7PCfTHiW6pd
wvWEoQHShTEA8MGK+T1vZ23VEs00ylKZNLOf6YzAbNoeYUaeKXb5eYgMIsrz
BLUdUrxDbF1gFhgaLJaKa7B76mT8vdB5Ph63uX8fJWrHwYSvhgoP0Yqgh6YT
9aqmloBlWavlLzGnS9UgyBXEr4g4mvBaEcTPwpwVFTxTV6MpqrdZVhIp0ICU
iQ3Gv8H3G4l6k2OGqodmUFZfUaoysVylYzi7fSzqx2GEdZp7E5SC/enj66C8
Te/PncyCJMzlrH2DXCWnheJl6r4WWIl/nFF3YvCLKCAL/Kr4ZMjISGG+i83B
x+W+qu+qUZwL4LK7mU/7q6wiXRidz7Xla8vr7nNwExxrwb2RiGqxfTLIvQZb
c8Mzrpc8Od2NcLJjyqbGzwFbrwy6bDuPVODPK21eot6ShLSehCAdiw0ruejJ
7eDXyD2TG93jb1sBAkThzlw7FdmXX0kT5/vYgLhsT/2hjBHUxYU+moE0rYJM
YOGiSAZ4Jzezg8pU7C3zwbPtuQ6SCDsM5nG1AT9ZZWwx+rDnShzh+DJkhqbf
lzl5vRfqbsAEcLofqC6gT214N8MR2ZK7TkwjlsLpjl5BfFTLjGRZOizhBFzp
Piq6uSfTXJxrTeZijr86+/n1t7+dJQPeaJChsXUdtGfEx9YIrtbzTh+POu+R
hOI9n1nnHIzxCEzZlMDP7wPEZW4uJPpA6M0mz4I9KwntkV7jxdlfmZD7/WAT
5nd4VLWuu9GMOo4na3EcwMzTY4J6WX5pM4CugS4t79WEX6lobZmnA7cWyyET
1jj0v613PIlAju3jXpkxaegsy4Ceq/nxjfN5NrNsdotTq6ZryyrHrxbJ6zmp
O3soP+2ThfMh32CjTXJScxGdP50XKl9CsgG+og/xnK0v/uRlsSF3p6iv4JAk
QeLsDfgQ1yCkm7iWN1XHQniSNqyGnWLzeedpnqm8BG67Mhp8tPCXT3BDjgpM
swnB9zkj3JpB/U/ZSTML4nItrvIxcVEVgqQXGB8W2vDFYw5a7PxmtBYjIbVs
/96VjCBUPf5q9qS+BQp5ezbtO4YkY/P6yTM5XsFKq783MX4sTEoo147u8a+b
RoaGLNILwrxviu8wqyjp2rSKAP5MpTYN1d71aKhkLF0NIIMYi0zCr+1ILdFT
g0cVJE6QHt1IBb9uSXoRpPJOXOAqwrvrkTNGTD3TWLrNGRxfnMl9ExDr5XcS
d5fQuE5Nuz65dxNnbe6ZQ4+tERrWc3aYv2Hey3khKhVUoS1WR0NkLClxp1v0
6cK1qLnC6T4BWIWvw7/G2z+4GrxaONkNV2WISI+RsddvEvE24KMLBAs2Q6o/
fAYVB+p0a6QB/mS4Lx8PcvWzu+kQtAHvPG8fbx+Co9Q4U7fSgJdKsguoxt2B
CvYpPo9wOQmb8/HPtoj13mWldsnZvt6FZwLR6Jlds3luqHgziQDFXw2k3u5K
0BTGS2cjV6+ipYdni7YdWQ0wEy+RwGZexf0imdDa9CetXnDnAHkHJFiq4Hkn
kN0ajnvEv6qyOu5m8YPc24hLq4WnrHqFQAdKPNOQh7I1tnqC8o/Wkpqw/tIq
suOHeDy51v7Ftu2ksq/kpvgwhvOvyjoIOquFuw3mXgcigILlL+6ECEXHNTEM
ATuzK6n3PvfhWDubR1PYuL74Cbx2CDzrRrs+VFwraqVEePJlkjC1C5h8O7AD
1Uma9rWWImMh1cD9D7OfHZHzXk/SkucCp5c9lEEIzvVEU3J3CGur0Uzk+47O
KYFZM575ldKMEO0SliBdmGmCmgYOS6iPNrg9cUdsksoznqgYIYFi5HtDCMeR
UG+HNPxepNC7y/pum2xQPfzXWRnhBWAum6kSfSJIQLB9G3zI5pzFICaTzd96
/DfjUuEOtfMlXTTHTChF9FEcug/v3eHeEssvmkipeDmXmq+vf0vjhsn6ubj1
euzM8bD4QL9QUxFI5Z9pxqCsGig64pWCRwziK18E2IijLoIC8N3JslyDNyeN
gS96Q0CZY5+RSVCY0dViynALIUisQyOBXicRrrtQTPgH5jTo8x0ovpjrEH3M
77pRmN5FGt5qi77SR5Br5g2JAVoQAgS8vYMDbAetnfhY/LiuBeYAN52W+dgy
sUD3iYUdtqKdQQqedm8amLTgZBtgvaxG9YpHKv8YMOEuVdS1fcRqW82Sam3i
kDvIhSw+B1KWBa/ZEki92JWYxQIRzWFYMI1rmUA2Vl+BdGrn/01qMFrWfkkr
f7DXenXFn2UtaYQ+dkQfs0AvK/8Bkf+KDYYscsaNHgs5abI8TW/Y6QG96XRv
8Ba+XrB6ckaeUB8nZEHNgZDcF5t+WXFQfuYYE0GbS3IJVMGfxgtruK4xCU8q
10QKZQsa7QQpPNFh/gLu6dysMxRvpfX86teQHdFOw/3GbqNEwlfXW1rtlxUC
i9t73PGwTyV9oG2vxWm61ykgF1wJMSEepqm/s6yukTFy3Z+yMNMkOMHQST4E
UCSC5ZRpfTE/To5P6YgBU9BZxSS7sGUFjUsLa3+PWjqtHeellVCmfIDo5tlP
nC8Rip03l5ySUFmc1WnvV2zyKyaTfOntxR2rlS1EdXck25ortj2exHCRmHSs
kTNIjqQjluJX7Gdag0vZg7BSs1zDaQpwlyW7g6oSP8AWzTe0TON4ZF1DQ/8E
N3mx3CKcJ7ppUh3Asv2QBI7Qu7AOZJn8Ta2u2a9Lkw1LXyNyEB13WHIbtkmG
iH7AXjDv+ZCt59NKCVHt+dxbJ85mrdweziEPy6FvWs/Z7y/o3oIBmWFje4xQ
Dqax+XBIB1yYVQFe4jBGPfNDrm8ZkFLFnaUiTT5UZINA6L9Ahb7h7bgRcbNr
fdOdYnJaHYHzfexJKiXmbK9QxrRFu8xUf28J3kxLDY0sqWSEX958npQ7zCv2
P7a25ECHlkyRpFRAomdUq1BK0nTH904wqHDLjLfS4BA8im+ggoIMx0JycY2p
e1njj2fmakQwRiFxinCDaCuGTuw1sZ7CYwqBnfO3EccHhv//5Sjh/uBpiNAl
a82gOiBIawTbP5RCuzuA1RHbt/fcgi5BfJT4s9rZr/Uij3EmB6QNeNbV3gnO
T9w7EozhFCM+jnKppXIqmVMWqZWUfRK2Mcs5N/0jkjbobmoy2ppFVz6b1MeL
mt1LwybNgqauGoN5hUv5xbFZlZhAzDsaLafYSoQ7/P9MbxLiF6equwa/jcw6
lU3+seAoXZ111PiqfKzBK28imwo3+E24Yw7qKDRUbYXsnosr7weSX4qXe8pB
ZH07axtZPm5N62/pp/EPxHmHaGXgUK97qI7Ko1O0bAF/FDupEfa6M1ZQ1l1v
CdLeiz0lpb83Fs+9QdOClwrS5qy3xm1Kh1qLhvmRDtZUg4dbLunGCWgNGsSl
xczgim8ufYzhM7i6FNqr0S3Hc+XyXlxYzu3QGjSur5JLu94/PxWLJEZUF5Qp
a2WCjbXGZg9JKtDKByYHvMggNdrCrXk4VmPWldPq46e49LJm3MGYhdkLOwF8
AsvtvC0SLbpu9CD5/AJuDCPLyqOMkMJfVMg5HQO9Y84SfSEr3hvy//COZsuo
BdwsaBwYvWEfb8hmMfFs0aCQfcQ9ldBkJ89/UqVJ6OIwHEui/CiDgiLC4Kxy
IuSyfouyAqJClb0WcVL+CjjHR1HtPt2hw7vY5ZvVJBdWrWCKF2s79UkTeE5Y
lCYcsZP0j8fSoIGlg7p+AZwYCmAQm7xNwaH08odfeaNfco1WycG+0jCImOVs
VgzmOtd2YKI/RpAmezFj7e5G/vrMreeVUzR7I/w3BQbvJuej4Ey5XhajhEZm
OjwZjfM2pkISdXYcjf12R50+D7wP9w4Y7FL3Wir5xs2hCyHuWQICIaL02zAH
Y3P3S9e8URL56rYjGmQwy+5ZBfjJPDCBsVbZGZ3F7u3RteSU5VMoTLCGISl/
rEjNS8Gj+sCvRRxRjw1lqiUZgHzf1mQkCU/XIT0KWQ8manix2SnJFG3Zn15N
MN3rwg5j1S4rVcJdU55oboF/mnefdd/RmX54fvTyhRFAMcFz5C6Gyt9Q/oMc
e+IvR2bFe7sLnwkqeOhgoJ9mhY9AhRK46iOqCLf+AlE67LFz5sOIxzmOmzkz
VMzvUIUSTnq0nYjY1VzGOJQmBFvzWsKz2EzUnPeLIe90jvW8qhKB6vLpHGjD
3d/tHlXr3ugDnoSSXZq8d9ZjAxf4Sz3ejZc+AP10iiJXEueRMnx8fZPTu+vj
5sIl9890P1hanjOer+uv4ADPnU2XFUNVh2uw5cYJyYDaWTJjg25t+bulHPzb
g2hjZx5WwPItKVD87sWlk7A/GDM2es6LVo2cGyUwBj/T5E40yIULVbHK/wiK
RYXl9psP+sVCHMe/QiBXUIL2OGunf/KHxpfDqS6TNI2mmj9uZKI9uX+MDTv5
yopk4ZMnMxuk4dJr1v/2HdqS57voRSrQwuZgu3nfty/J+4SnkH8AW4s6v+Nb
cNMCgIKFPmm5VHyf4NjEtXoQ/2QXLrY0lpBQc92PIgRH08Reu8L47MXQA3BY
CVEr6haKL+vYP+shwCHsjjhW/RAuSK/v/R2alNrW7E7fbqkAT7jpqsQIJz/u
pxGlyzyfb7y3qe3BZz+hPHe6hxiG7r4ikYHOKJpbHpxMnRD7AeZnJbNZcXx6
mG2C+6VKDH+6+mIW2wUUEWJqI8AUV7urQ6volNyWSzfAVLSXZVDMWO1Ftv/d
+GPxhH2rJMoMy6z3u1TfnVUZD70pagxatis1X1eL1JA1MYcheAe9y4FXxLiZ
xsITEclrtzDpNAcJAdWc0SlVqTLikbbbk7llKzCZULfApYlxc8vQA3P1LCmZ
3W9+HtPcsB8WVV3iD/hyWuOmbgFpgy5THLDjSDghmZVBlNZv/cl8zTV49PBn
yMbReB0PpaeG5RjkCbWxlDArpelAn0EPvVsy+fL8y1ieZtQQmL4GWq7hYFJw
QpWcHUQ9ew1swSQD3g0xfypo6fZFjytRTkrl0j0ndHDBmvrYGQZg04fa9f+6
5mJnKLC6ZwD7pA32YmQ84eNSUztSeBo83pedEel4hYsfQuA6IF4DnTMwZu3v
GHlUgH6iEGxpX3SERgdnb2tDy0YAYxSJj+ImSXTZto1CImS50viMBNQM2ZRv
4AWqKm357j8JHSqeufb9x8ENLqggCD1o8SABgmn+IgJalXi31Lcr0hs07pPG
nHjAP6ZjyRktHnxxipDNEjoLmDdLMDf5e50RK0Ol2ZUr6nmnKZpq/dChjxQH
xGMheYvGDqLuRwjSvFWEQdjWt8sq5xPFWjyPrXRPAqF7GYrR3cg3iu0GOIPz
pbLBrqRzO5pX0687xSOID34UekwCSfIBfcmhuirhq5+8cXA5daGyadcV8jcS
7opQLX/T70htFMkoMz6WiodNIX41WDcBhYzBiTO5GK6K7zi3SxKtgFzoH2D3
lUg8VTgosEMH41tJNGi+iLY5X38IT6G/QR24hUGZbSaiu6VQ/k82qwZEaIKf
U0TKmhHA5NJxUM6sH+FpE2FVSZ/6fqdu+5Ym3hmFHsjiyY0LCNHKKkmB4NQ5
UIuuiTW9zVLr8iotPAWYie1qn9q75L6kWDnZq2PgV0JlWy1fnKL18WbdG0cM
03txvdTEJhwQopRcFks0vi9/Wkn76mw6XPt6EZgRI2TG5fZe7ksn7jhwO7fD
+OziGjgorqz9ONnrhjxQFBeueu/H1cJcykw3pfgdfM/DhJRmw2hCEhneKya6
2YiNiCk9AHzhHnypo5nLSXv6JFZP05Q72TUjsMxVJGzpP0ITX2p1P7cjGuNM
IhkAUdJAH6VevWNZWJVJtrhgnNOsoXVG7Gz6jXVOHIwuZnz6x+Y0pm8FleAj
K8a3mhZ9POZOm5YzbmYcKc2ueRI1yF5jlOsXsEKPBgTsgHJB0aiNuyYXN6vs
/+WilGgDbezJlnP85hjDfmoPvRqkI51Lqj3yzzGGXeRP/2R4VCnF242LoxZ+
1vC9DXiFjkZuIL34iHbL0UfKmgFdvfMUPDTGGEXNztAW87kJWPfSjVNvOsv4
z8f5N/E/Hn5hwp42h8J7adWNmmjMyIqOuCqxZJkHO+L3IypzxYxAc2Yudh3h
5lMRUknPiYv4ncqI/PDKCiEIRuvNcZ+7dd1dJ+3tfgryxbDvjLjBFTk/zZZ1
B9UmfaPJvcnWo5nTyR1t9ITF8b3I7BiJF/l1RBksmbvTAXr/NFWDzn2nYB0d
12SlYIZpGqAOUhcZD2v2lIN00+A4pE7q6CccFuLbZX9GkKSPCH0CJqovBVar
a1hpK6uVd13fXgroIXg9GDDExI3KzLrq1yaCstzw4q1c4fcJpMYmsINN7M9l
zD+aCg2MIGpaDsi0PZnHZo9sTHaTdDnjdorbyiha5oiMXMiKuHN++d7+j4JO
j0iCda1LocPDWRC+6qTUu07w9vdhNaa46NdZcmGEqE79euqkotSgL/Nims/D
NVTpEL93Pi1bcoHw5lEm9Dfj3AJeQMGVrM6bJl3siqlznCAruiffZ4KDEDSp
E90G8Xamv+dRAOVcAL1IHG72GJo+Ws3c7DNODdYDqmL3to+ihJEgw88RHJUZ
t6w/cpA5pMdIJHSTZi/ix3fRU24aX+IH0yVkv6E1geCcpVh0xe+SN58wSTrL
JSWubiNlzjpmMm6WjYOHTje1RBgZmdXwFUEyzVp+zZy2YiVHk0HM3bFNw09T
W2gIvy8ZoodOl1aE3EMdmG6Zn6gYte19BpJ18je2/W6SzGDKvBu2Rcw/EDdr
kppOqXR9xuwdKaPjQ+iIq6sNE52+YEGQAqZ4VPUJNjmWy4IkyNmpGV5ad5NX
8bbbp2E4KMW2PxIiX824GE8kIHPDNuocnwNQQx0kkzreVnccZYjQlc0Pwl2H
nV0d+rvll3lQGPazn7G2+J+INlCE2Lrnzayp+Ptwr3APOorgP0tQJaxHFuWS
ismCktMAc3LAzMmfpiVIsddNPFIlR6sA2FqvBG1wc/9Mdh9YSZ1sIYiqmfhJ
Pqu50njYblgQHA7vVIwtoH3PPJxGaQY5LHbf2r+/Gy5kKg4B9zuNvKFlh0AZ
BIUXILyCadZnbWXlFMkDakGvYT3ODB+PQpUOcYMKqlqLsTYKEI1M2Keuq3gw
zXpqSZCVkcOJUzZbO5Aa1l1WexKAeW78NVYe8Sm0YyhqHIOWbY76UjpXSZ+O
jrEZpesWkGXUtDSRjmJ5zzYPA1mmDIkei8mx3iSKXH7kvVufj/yffhvkmVJN
jQTMyD2ccPpL1OmMHVW4fruaGWxRfGAAcrq5pFeAVmx4flYvTH6BqN+v9uco
tdVhg9YvrD20GQfVy1+pc3xybGZsoB1yS1JDtPVKBlx5hnk8sWBO1LMWQDJ4
zdlEaZcrQJVT6PsCnzT5ShnxcF79pegJuTeKLjVfSCIljRVGjI1F8ju41iNE
bH3/6PHanuQ5m+spv5uhEC3FyMqJiaio3LtkZ32pEkiwgp0aW9RTuyzNsurj
RIQV7GUjCya+HfNxA91gJSLjNa5EWOhLnTkKkiQOItBmEG85Z3schAmcpAwE
fsLU0+o7jk916XbKke0mH/MU5F9X7FIBh/BIINL1fYOspQ7Km3c0XHy+41cg
T2Vx8C4YF3a5i2hjeAvUC8i9OyWX1meLrsD/06w5eEuFylCMsD+hkdTgd5PN
NJcR2KTV97h4RRQNzkPYz90FtHAPkd46AIwJVJlD9CsOrncvCKRjGcT7hY17
2EcjTYTeZXeGS4U9LKb9h6YOaRNCvZC/2jjpWeDdVgmiwxVtI6o3D/91pJIY
XqA2bAQoudqbjFeklukCCG8Pu9Dah+ahW+B6QQVzP1LN1K+reBZJNXXGl4/f
3XJmfrIuQzA0Vfen6utBEeucv+mOLWe41H8CkhTPxBCAIjkpY1Q1TpjKZMaz
i09r2+nLXP0Fu24LZrYrnfvOoPPHk/NvheBHZZHQPWVD9Qh9+lmo7MVyG3QX
46T5eCj73pCNrwElgWYg+xtIfZD3XpNbnXtZzaENinsVF0bD3A9agirP1sBn
Evlq5TrJPnacH1YFnHuExsNIiEqXEyaAsENeCltYSeVotVfooL1jLmvwS/1A
JhEcQKBVhC3wpJUIF5IXHgGjBD242tKczd/lQjojt36QRjyjxQ8nMCkr9UID
jqQJpuJTYA8itlUVm2lBHIvaiQViE0q3w2KtYRmyP7c7xNZGeJ8iqHyixlG5
b3NrLLIMCCquhzQRg+2aSSBv33Troaz5vOkLSqVqzMvnYPoRy2JTp8bc+NeE
1+A0j0aiboT0VGEksTQmGHq2PcIPmxa0vT6Yp9ILYW3VVAIWvy7Wm/3E/Eec
oaVSwCvyZiIXS2HxoJaqXjbj8tYlKIqt5GR6d0DThQWOEBlSDv/oJv3dHBvz
DpibQ9FE1EW7g/R6wsQQXP8TU+ZiERzN8HdiBEj/4ZnxJj2In9FMfuKOWzKG
L7lbDS9J0jlhuxSsYnfHxDXu+ed5MdlEuP4wmVLfy9legPNN/1liR1GsYi99
iQAnk1omaioKgwf8wUPf23A/CSP2L6WhdM0Mjx0CtzS0DGcKUxzVxXQyl4Vb
aGvB8SFeeVnrLXlKdIfhdCB8Q4PemT8q1EjqaxdwpVTmdxAEAS33iKClk417
CiISkDLiuF7pmCZzmfpwatb8lLre09HMTz8SWDK63Ke2Cf/Ty/birE4JnWcr
P2ZWVKrLcCgBDzLBiXCNkJbxVFSIz8GbzbTjs9WoONeo59iOBrFCqv5VRSAJ
40sHxkYAtj+/TPUnpoQz9wBANxb6g47HWsj/XshPnSxybpzKIm1/HLpc6YQD
IsxYX78R0wxfrCeK5C5vE3nWdvPgCfGtdBqkzuIOi/bG4yLQPG7AaJOyi0GY
Rw8l/pVCwL3Upheo7FckkAEcb5rf/1pU14U/FDGPWYhJ6zDL3KIXd0NwCNVR
cRye06KTAl6YuGavKssGrxgwEFpguK9KHQ/W3HfLpY0+frpx+gpPRWPt27zV
tgF0DTfzhacH2o5DjOxjg137v1FJ3YrQ/E1vbLg7OZD/tjMyKNdJ3GVKO/7b
/zoQS768NOyFjWDSdQm0jZjxN1q9TlAzYJTkNHBgG+mIKXMCuQYNqW1q4Kaq
N1CKUtiVwToUP/rRriioZXnzsi6SqrJ2t/3rD3bm5jpHDPM5Tdqk+lvozc6Y
Prxgipa3iTHnKlLNafFgujHd0mV8iUHg/h3gzljbpWPfyhBwfgMmHvX9fTlc
Y5k0VSmiU4018BpuejXL5ImRrLJsmA1lH8a1NvyeNigIWFd+xX3rzwxbn/pn
NJAG4eMx7gYpfjc3TH8AKRvhuJIiQ+jRnUHgVKz7jnS4c7lnESY+AxeY52L3
BcZZu+L52BjS7bKLLQv/qtZcr6uOrR9W/xETzEqTGciiI8xraIQaw60hAmat
y6XmQ8wEAbm5jicnMwpulU5hT+oLAvre8rllVyM0Hx48VZA99W99ZBt+ueQB
PZQwRy3S1Y6Wg/FzgCFAYECJmUr73DlrDU2fZFDbE3bh8tryOnzBKsBqKCHm
VNpNK2WwStcg1T5ImapGX4vOWtjm0E2epQyBO76yG7yCKuQSXthvYDB8eO8A
aXoXMLAgHgZHj+JnAPphJG54CMuckApVFThKu0DqXTY4xYwppvxe8o6TgKty
9VYGrKhcRRGm0A6xVPtV448dGPe3k77PXn1rQeB99v0uOPPAt3UJX2eroSwP
N+IpCJ4anVNJHi6JcuyL7I2epguUWRtqV9Pz05HNkRKXicyaqqE4rWUg3Zvi
02bSSYUQ2gOjwRIMg3ITCCpA0NQQg7+bYgj1DIAWFqr8+oXc+r84/4gUSkSf
xpLkEk6aGoubC3wE6G8nMYMm0QlRfdALaUPYHMQ9wg2luV2XkJPo10aP7NzJ
+HiDVNItiEcEXdbhaaOcc7oM4HouQwGOSAPAcCVaVjiDmO9+3x2WDjuDWKIW
9A7f2Ir6irZ5boVpDMnpJR4i5EOVCKb+PNEVy7SSBcz1VcaoT7L48YSdrllp
ZwSz0PMGmM+gej9LF/QrQNSjeH/TpxqYif+YJXBcOIJx84zPNlk8rOJyUNh1
2Q4qdzsWcARoEq8JN+ygZVGvy4afAJMC4aBbJtc/64rz4w8cX3ihhtS5aVOh
zORNDXUJw4v+QZKKNGq/aQ4BfLIl+bu/FWwpkNEWVnIxo5XCRjZMEL2rLMo4
XbOk3XrQ6usSnddFTJPmJL/J6XxR5gT3dYQL6tdECeSupzms/g477gaT4wrQ
WcbWHkWSz3j83jG6UAWxSnlVhnlpoq/VrrVCjYMISykn1IMQ1SfavfbS7RFP
mbH5ruQyZyBve53GrHua7Xqgkzcsg4n9fCXbQr7vPuh+fjfW/HHMn7Xlk0Vj
ORNwGV9G0ta2Elsxbr9JEAnZLtMVF+eOyuuiqPgtWor3Hs3QCNrRuya2nuQx
LOLlwWDzbpwNLn778oTBUO5sVoP5exGL0FnHDNBvymSayoeeOGGFC6st1Rca
skIvK+5ca8Jmq/K7JdDn67ohnWp7p+iM5KTdBRnO4l9nBXC1lQLNL6HAMbVf
5Yk3QgOE/AjAg5xZg5tkTiTnZlJdfAthFKLXbFgCy//WUx6HXbhJ0gfDEuuu
yv+075vS1oPnUFJPhiq94HE9JTTyKUzeM8INii7pKeUJciiRicTb5tf76okW
KU3U7J4UOF/GZQpCLG28QiXmQHSG3sYrRR6A+VO5bTCheGV43N0PuLuUSdts
1OnZcuxfdaSMMKiWWA4EwqdjjmSUYxgOUWdDbQIrR9dBi8dJLvAD7r4BXVK5
bwqZA+bwowb5q4wAMNjZ11WGDK7Qbqu9RCZJWivwmvVfzEgUd5G1YQInh/9n
9qEqf21jO3uyKivtTCN0FC5rfzFQ9nIpm4JOCmdruNP9tyQYPaWBaMr+7m70
uAAV8giWvF3Lk6dcDzJPSV+ro0buYw7vHMHtr3LWnQJk3KoLrnxdjj7Xbl8G
uoZbDGRGV4+l8GUjqZcC2N/A1/7S2n2co6jkijdOkky0zR5kxVYYgeipF2Xw
m99IY47FmycMK5zqK98F4kheueuMYGIMGKjkpfXmaE85yaUkO/EHAOlVpW32
jBMjab1bswZphBOGpkpyYHaJOMDkcmpHmCXIjulHCQ8g8VrgI+sAdT0KybKH
o/Bx9PbHCci0XyAzloK53lTdizsoBjv3kAnfA1G18wFJ4ZEwLrwWXjfVbsMB
/jGVvlr6w5MoEO2J2c1o5ZBAe3or5z78bbayR0ewmwl1SrtysETBDdn/NAmh
o1RI6GEveJQb6H44GhzUVzTTJXPW3r9cLW8U+6Mt9BPrh+9UhZKrM7xkks3l
2CvaPiyp66uj/VLDJhHW6kPIHu/zdQJs0XiarnUqVKqR1DP1jmYZaZSKh/UO
ln2Td9d1j/86Jka6iMlg83jUCm3Bpl/lYElzM5CJKr0+BcuhkdDTb4muPWd3
Y/+4zkBdUIZ4KRPb7HnPbQ+FSJUaUR5S39st/8PTMidrYrrHTwKTfY/i3uDq
r3uTZDUGqgf1Nc+tD9Dojzml+P6fFkTcC0Z4a4TMKGIY18DHRsWD6EH2I407
iinBFhlJo2gg6NgHsdJ6zG4f1oRQhpz/neGfGaAEFODh7Vu3C9LAZFdiJmOb
Mo/6msV/QQdyZzYMmSmDyTgI7/8MfslFRvn3AkctlCbb6kf8p6S1yfSyA0Df
7BPVe9OL3ik9bCaAvQUMh2vAd5H6xIf7y8OJn7FgexeaHmI3rLjc3UkS8i0y
KWv/UCuXokEYCwOXrb6hpWQ7ikiIXlEohmjo6oMbHuenuftBI7jrqsnMY3Yh
zYVVyjvbhFoJBXnSQ9OJW5UQOobrA/1wNey9I76XhewrKKgUYVx+Pv1LWo7E
YyhvJGstkbvEHV1MW+f+3AMJpIKRrbJZ1JZbjVAlAUnJgpfXj97XVaf4TJW7
rtWN5OY0+A8L1SLtWeDJsUWwK6bl38bzETSU8tgELMgY1Lo7lfhorb31SUHW
bws0fe3JJk1G/+lYYaanhXEkG4omMvN4Nm/v8ycrVTC0Q38lGfjdmNHwW79e
RpfZXfhn9PUqWrKMpSCplfRDMi6xyJWhXc5aiTdYvXQ6f2K2Zp4V9pHI1Nsz
fWj11EfaKq04zYIxUQzOxp0uqJa1QvGm0SvGxAERI6+5iVM2zUtbosuhNAip
Zuw+QN7Rj1HbEY1c3230LUhom3JrD1CsKjrTQ+aUL8TDV8gJ2JHgKVvgCcOC
AAZxDygzCHhQ4MFfB0OKWtLEzHfvSVdPL2/A+yE0y0wxISr/x8/fE4hvxGkX
Toiw+V8M/U6HuYYfUrAcl1cwoc7G4/nlkPO7FS2m9USIcmSvKBj7Fi0MkyAW
Rj+G1erPJA5N/cpUplE70qbWmWzu1lCuoLEjMdOdsZ+WWzfaj8mn9cuxnEUx
rPaNDlFCQ21NvhggA+X9CI/CFtxrjUY83xJxcSw58LJNlQbSNCUmsCvdFgA/
pKy4THZ0P4KSAVX+UwEchKAHo3Gl1vTo92OLQH7f7XqFVlKeCu7cE6Epftcg
lZnRl8NorzhRtnx7dyFD4hkSDRl2wXrT+5ehvODlERatVutmAkLMGk2SKOI3
T7KZpvYi+GrXOTsKjUFxCJ/6WljzQDscGRuiroUXImBIQ1ED+JUNEjiG+Sxh
SgWsYbT0PgF3JDzd9NHqPpDAi9yhuBGqYxrqMCM4PyvgWkMIRS8qodlY6J37
fIs+c+RBNRX1uKPNIY9+YEzPcnt4BJg/LPmnAGOsXnfQLym3t+KkMqHqxlnO
/YPI3m22j4+yu5AujzKehh2Gemcj7DPGWcPqzOCOaj0oKP/P1158a0OlDgVo
yXk79fJYcvQHRq0oQarYJK2xNAjQaJWFcavrhUMd5mQ8Tnr7ZQtJBL05rUfX
UU0v2O6+KdeCVtNDhOlag8vmBG9B0WA9f4IRl62uQ00B1FgKfzdVpD8k+0ZM
sYPhJl+i7QWJX/6F4qGQTeCgUoN0vFQLcAGRHYT1FDtqE7DHUTjYKPpyJX0P
W/Q3BKAiYeEwjeMjA5PW/UNMNw4D7ht2Y/e9HC3Ob4QcNgZDPY9ho1xrtyML
GFmJxwTK8Sd0mpmKdvukeNp+/f9iYl2qBjzF+37BESgH7hKw+1t9mMBlW6X4
5ObbR/Iro3jVLa1RGPtTRn0fJSYb6XlFEtaXJHXa7oeR7i3dN2NU1kw9pfMb
KMP6TGAasx0wYIBClzhoyaJTD7K9tXUd7O4k69amdd21HapQ8wZld94uZ8bp
vZSYFZwACvow40YFLg0zD+EwO/nwErchSslRqxYS5yJnScs93YxmO4RkVgSb
osjBo0NE7743a04qxfeIZNkt/jyTqor90uMVdh4mbdR1Pmw9Ym8zi1GL8x0W
tB8Qi3ccwg9y9z6vmkG9BlyK4Cecd9z37Stf2Uz1nTTq7OHPDcuqfX+ac7fA
fhf6FCFzyeqnDvNRziOkIEF/PBUYVWFgGslhjhHBNISIHYRmvUPlUprmxuNE
x5derdWu/b7bZTbyoiioWDNxVRp3QFdxcf0ZPkwrUycmDM9kzj+Q+HdTt0UA
uV2RneussLeRa8UUNnhwwo77eMHqfv78sijD8Wtc9aVdgrtZZfrxTCOJ0aJe
J8pCk2iDil6Yxseo3qdPOaFkIBpyUudbyqD+ZLZ4YlbwBSLjf8MY6niurs8x
RGUsc2YVMArn5b9sbb3C+DbYFK3BC6OerLo4wBJFzF/V2Lyl1hQemFAdoBqJ
zm/BOkg9tZGNeg0ksArgQvni57QlZnqwEogCz/k8C/SNmoZhoMorT7Eu7urd
3RzNDIYIj+wxgPbNXLq3jUFEpH+e1WEuF29j70kALNG0otipk6P22uXKmOwd
j3IMtMZk2adhaQiuPBXE5Ip2412Nd3Ry4qXgZOly3BgocojpubDKvd7uWKP4
mrGhA4j+EzolcU6jVGizo5sx/ZvK8MR+zCqhSubs/nCjntbFxJOw14VcVBl2
3dkFHj/0WzCy1gBbt+hE2NgDr6wBJkgOkl1OhzMRyWjRrgX/7DN/51dOONCa
SZ3y/Mcz0f/Pg8y9T5Fk6W/r2Qp1fuhtZj76W7l7c+L+JgOfBHpnrsNUT/8A
AZ4eMwVx1qo5Og43frKcnfcDtQY07JK/1cQGPtGomcTIvnXGuMY5NuNBZU8b
7+/VXinIgiZJhcjEAGQ8jrWH56gWSTrYtmKd+O9k6KHqTHxwS9W8QSLEvVML
NM3XS8nB/CwGxyjoEslLUD91Xd+1pwWvyEHlj6YKO1etTQOcJsjf8Hs2GOV7
3B/pZ98KQnsK7uEspf/L+q26hyCT2E0Vgu+hnwceQiUeSDl/tS1nk92EtJRu
GqDtO2IpA0d2tj0cQ5tju0GVt4JS4sj3KRaPCJna9z5n6OiKrrLfo6xH6dmS
b6JsNHe/moIpDdeGGUHQkJJ0dM+YNK73reBZ/UI1vaYcQQlINbGVBu02pbHx
YLiviVSPsSqlFedcDkRKBP0kjOO3zHtwO0Syp/FQfpjfVk/wk4pjwOvmyL4Z
DSAgZAT/s8V+o9GvWZ1JwNAe9Cq4K9kgdZcjZ9HBgHDCje3LznL6DVauepyX
/e6vF/kvawWiXcdr6AIqbeK1zCnQjA4FJrYLalnlBqOzAU/sQzFdgzBMlrIJ
BnY6ExxIL3/RWwTlfCLobYDSgmsF7zARWzBFmOBJU+DDbV1wvmkcNecMmmev
IDOIqzIAfHJaSOjvqvR7nRltUCMZzdWNQFepwtNeEk3V6wnxJnfMIqadSKC7
b+wCg5ARQVQsyPEmo+XoYWLuVefqaNBq8/OvLNaoVKMzHIhByv2XFoxRHEnV
QurCjprf9p4sd1RVYCOrDNqw8OXw7Fr+y6Cr2aXqDOzVNI9BGIzENDPpigQE
kwg9O0saJhrZ1ztBBqhtdL+sO7Et/oL+BD8wVl+T/TY0KW/hhA4YTAv6Hvbu
8dMQELLhIwJlK8TduECL5bMFliSEHehEfal0pc82uHktFyEV9jUqAtBqyznq
mkIYqptmZCMhqpDqNf16y8a+O3CyhPsvOCWjs1HILkWB5fbc+BhrNu+K4S+n
LN/IP/wfR0mdHuXdiwcxpE5H+9adoo1ndEzVOE0SycZYyiFLvZmzU7hd06CB
g48nY974tvsPkj7/MehHwvNPrMatDXasJFabFYOj+uzRU7d9exdx9UQo0nyE
zXwA3nQnxgAp7DHvAJuiDKIZ09qi+FPOJkcKcuqQU/sQX1rUTBGwyhtmyxDQ
Q6TW/MVO0fX4OkUE9t16QZa9QNVseXEK0bcT0e8So+lHrOy4sPVx2AQbAgOE
m8KNuXK53CN2JpjKMhsJSqd7lO6i7h4pKTAlBZJ7ISCkrH28hrchA3BY9cwh
8I+IbRwEBSrfTpUd8MCPlL5loDrWjfDntrzw55ZxKc4SxC8wW0jnv9t4MNTt
ZmircpBRhvf91fkPNuBh18TxzIJL/+6qFu6mkNNKogAoJ56oi5AO+I8iHu5t
M9sqqeGhlaagEa3335O3mXntyA9Ejfz8/v/csXRWISu2GNGfcERAYZq8ramw
1ccTaKZpttsNH9Da4blcY4x6NpqC9BRVTkOrFojVReAMmpcj56wD5EatxMka
Jzjy778cATnpeJ6b/SV3iH3oKm3r0jiX6T51/3YqFVl3qBJY47DTQfnok/sP
X2eePQI8pE35BmQTuhciP0ov9rHYwdgHvO9cdtBnSLWCjhSIyTyRl+qwSP1j
jR69it9N0m2/Q6lDSCoqepGIB7qpXUXH9Aon/5XAeaWO2+BpX+Qy7TGshKY8
gfdlufR1gFHuBNsYEMOONb0NF7t6n6/kVrghxsnoRaMwYFQe0CqMbh7nJZM3
buOobSuwFNOSMMpsP7DvWiCqoeOvsSQi33CgYMYoYVTBiGVZyxI50nH6ZUEt
HYr55Or81DjuefSM7z0lmwWyNJDfeMUwhfez9AN0xJhTlMtTpVKUJtjegf29
o90VeFOXSSS479DSdxUmQDk2oFH82t9IBY+kVIdS/2O8BWIb5giZzrBrMe8M
5Lg1H4JYVU/yMaBvUb6PA/Qs4857EP9perf3Vftx+BIg3crjbgvela+XAWkQ
l4+nogW/GhCdWgAjJvEaYucSUTwLp/zWY/JSG90UUD9Ykoh2DqgQJeOFkBqQ
Xb5ikOAD6GbWYRNb+8EWUplPGjeP2fk09lT8iR3bG5E4b9lGujRh0R+CDoOR
AXT1kFxzCfL2hMn4WkP9U/2ip1nABxKHjSnwrMU19/UdCg5/bgBPco6znMqZ
YKkLZGXBhCn+dre27oP5S/y0KeBFmMEOCjUjfguI9ez96jqq9oI816NsPJqf
isnRUv/OAjUTFCoUC03nAW6TZa1PSyrNtS8cJkTdQzd6DulYUP1Yh5cm0Xue
1vVPVLWtfouNXoIIN8c1zyYSZYLX+Vp9Wgv/fblBMKTpCGh2gRp8qBYu62Qv
+3do6pBc0tSS1vmCsMGt41d8O5WN0bp7pmM4gG+XbnbIKu7d690Pu2Onyx1/
hfpjDs7wGTq+ADLfX3bX3E4s7XTQkpWmhTepBwiKaH8jfyqL07wRNKG0Djyv
0ZYWjwAjsSbnEVCSsvsjpKg6lgQJBlX95nHEieI+5enqpuhXwwdH3NayeSZ3
IEbG9RkA0VikKp4G4l4zFNiMSWO8ElMI3BmdFrVftZtv4N4gJW/ms3/a3eR+
+QKT5+Y+NjpDihwaEtlhCmlNLyZLjMABXK1BPSm607An/wjf3UZfylbkHt8/
p8imJVaCVMzuELY4XHIss46hbvLvr4y1iBVnoNjiXTP1kBIWS6AwZcYDJ5z7
s6ZfwOWG+W6Mv0pHqADQsFjyh3gtGWZ46PPFZrtEG9rFLuqh7ZuEsp5qZ5Ay
IqZ/sEyBiGcC3+GNBsJOlFOgxUa9KCnEF4GOeNkRdzhEE9B/33qOxYmANDxB
1VIVDJCC5CX7tKh+YIFb82vpXdln9VAjxAgoNy7cVspH8HJkvPSTYt6ak+tM
Tn3dqr4sQDtl0bQzUhzg0DCvuu2/zAeUwJ4gZOo/nUBG2h9Nx2halSQjPPD1
mxOxIFG58oSoLXPw3Sv9E6tv+eCdgR9Gq4cLVhPENKKZpCB/SoATtOQqDo/m
NyEJb2veOW5mE5N5+Oc3S408OOAS4R43texM93yKVTEqUFqPPLxPHofYI7e0
qtBOxN2krYQRPta3cHQnMgEWy0DXsnSgyT8EKOL/AahMfQKKJNp6f+KBl4Vb
pH+YOUnzZ3J7yMNJyf+6n2LMt5KWVSwSlGvqL9tg9GaFAT/PP8JAVbvil1AD
Fz3bPIT/1by3yn1Zv7Md6mDJ791my6jTvKmMB83DSUs7v5U/XqzcSucOS7M/
JxdN8vxAvP2+rSX/4sSSpeF04V+P3dNogUqoQRtUk3IULLbqqfMDWrrJy7xf
hnt2E7KzsXteShoDe7V/xRncwJJg+zj8uHy6mKsbTxikC8AjjEH5br2+s2Qq
0G8W0/GlZSJ8/WFPhnYp1LeXve8ZEUDM5Wb9wzNgJn7d9i+ZCZqwexRPM2E8
ve3t+ppm/sgaP2MtMZ87m5yos4jv5KLiFYpEF7q97HWoxez6zRphd73QwNKo
usZKrvMV0xikfgyjxdtRO9GzEAfHVySOBblEDJnGvii8t/+2ITI3D7h/jltq
fRyTV3ZlOvFxIgZdkEwA5mU6TyninExy0OT6h+2vYGn6sMUsyAYIYOJ0koQh
7yl2D5jEtw2Tu7B/memA3MWxzzqdLbpKG2o3wfx85rlVolOF1TCZEn4tNcFb
Drme9xVaHNtdFUAjOV3jc/9drSFLRbpy01HAV2aAmRyl0I59t3k94h0Bmgss
+u7+N2Nu4GvvRf/3BR+DgMyGgBXHk3SDMoh2DZRIHeUvrj84mBtCWj3C1Lfm
rnUbIyK6KXfp6NC/tc3lYMtViKeZNw4H0ZN8pADZWh0iDbUK5hkLOArQxSRH
3dIIsbUhZWz/wC7pLe9uDLr1G06jBJ0siRvkb9lHqzatTj8VYS9bS11APVdU
RqoLGm8Iz+RDhjHkfTuGdqdWOVFTmOrSWeRvzle+6R6uK7PvWrGTA1/1St/Z
zUp8S4a4N4G8svZnkGzbsl8C1+3vDM4bVZmGeYcBv/G2MQQVW5MwwRw9/N44
mCYgDf80pUG0rIwAzRgskAK5t5/DOmWEVjl5cE3+NqyQEIOwBhVS1kpFS6/D
rw6Gt0hiweMxKpAWVkHGV92gGrTkOi+WtjSMle1J9mBR4A7FNzYfiT8I5gPg
ubKq/4pltG1igl959zvA6C+hnxMzDmzd8C17XDbTx8NCXayj1EGs2lxHPH1y
euKsxdGzq+fDZXB6n14bjFK8suUkmCExzy7b5VMhE8ZntNorZAbWR2kOgJf0
t7MnAY9vQh+gW89hqg4n97KmU9+5RS8u4x6foMSOsnopgTd8008+TcLLejY9
aHrJ+O11gY5ECZWWrvMIFexByrj0dQjjRECyY7GZ0df8JD5Su+bt33ZAj3lI
txXdqn6/1S5gET1LMj7ndjX/5B7Iq3uHlTUoGTkFfCNn9N2STgoVBT8XcGSc
kDshqgRfM9WWBx4/Nm5OUjs8oR2D0hJLX2XrRhL9P3Wv7oZY84vXonpxwbwU
X4uQTlSWfodpXN/k5U66zaZeKCru2zAMUjtw5F3+mVQAc+zXcOU6+OQhv9FZ
7hUr0QmUHJlhvr8oqsXL0v33IK1JNrlq7ev59Bs7yDMq2x2L5V0zpF4ynGYT
7yG5qqb7cZGs0VWRnJLlZURdoXjGopimf7dI4+tFU8tyBnsA3M9dXM6xF1Qf
PDk2ejQlpreJdzx4JoJC6+FJKzzZ2nUU6APPkFHt/R1dOU1VvDxEB14MNckH
gbd8PsT8MkCiBpd+v9bUU8RR6j4YuJGTUbfMwCawCpM4hm278JLfZLz8YVow
P2Wtpl4KdR5DsEsud1RCDzvk+r/pmst6M8OgOnJMpr1HZptaX8rcZe8Hq3b6
K66nZNNkgKrBB3LmrsDkBbzHLWlUZwAhyW2BZGxooNzhU27lLw7A+E7p71pK
U41h6u8MgYdl8witdRyjUoVvVzky8rgMDj5cq5/S33x4Wlfy3NpRNth0zt+k
B7u5rH5r/lN3a3dOd8j9s1KkANF+bjv6k/0mKtSuI2XXqwsJUmdkg9pW2Mcx
Dv5ePPbPDRkib96DGZ4OyaaAPk+szYrHWSpyLcMmpZAffqM5+NwLn9Ax2RsA
HXSwU/YtOH54HyIcSADZnl+w1s7pMyqhO2d/8ggGMZ0PVzFW6NVlFa/BgSOk
2I47TZM+o7yp4yTe7ez6t/p2fMiw1lXCT1OVxG7VQWTjxuSMICfgf2lHKJgd
phwGuS+TJtPDaGkAs/nrVOdP3df0DRGt2zysM00bhtJ9QbL0csdeRyfwILRQ
UOXtt4aHPziLfHni38eblEVP/+UEz9wsWbydxhm/RsZUDe3LV7TPBA0tjABI
qpdavjQL2EeaJDf53kYQFJ/7CRtyaS+ZHpT8Xt4qaet3vrw3zkwBP6cZ5HIp
kXJytUJ872fgKuDCG41NbxRYyxQKFsJADYkb5M7Wsxa7smlZ4Rz4V8MDyk1C
CrnGSU/yTMjqb7z0fdxRGAPxi1pAiM2v9zhmcyHk0IM94oKuvqntHyhwfMCl
c9fiB6DRRuEKPRBW+78pI6e5LCOp1ceaJVbdigkAHTwZcqqWeBC60k6UsZMx
O/RWuAlTcvsZL3GaFdO1YGzuuiabvX8DyeyuOLJs3XkNA5V+lljv6zPwVKOE
UhmIIEvqLjyTPEsmZ60ZVVsNv8U8ilSi1SMuEopinuMo6YiOg6w8fFNsztGg
073SE/W9/b6hIORArIzG80O/KKArFXS9atzbRfFAaDBPDtMi0WlOrUJuWQXR
2cTasO8cBh80FA2+ytgEtI2NGNwpVIDk8gDbz/+yJK4NIDv4eChjbXKaVa/A
ckAf7DZbWZlddq8/oM6ndxkRieK/wVP1gpeY7j5C2TeBNz5R5LswpDbJYMHU
iYLLIAq5sdji65wgC5NLK7kCQJ1vGgEFIt8KHrvDFMrs5zGXrPpNcW/JayCN
0FDegA1P8JCGJ4oLNf+GhxqbkLAIGerhSsjJKcxFCLI6Xv7uF2u98PTz30e9
yafFMXBAZFPJCjQIJ7EdzI1gWmWrZSGT1EEajw7fpENa+WbF0Di/B1CEsdaV
/HBuKq0zrsKZ/cNaOK5JfAkByWy4KNhkqoVeCgA5D6aHo6Ya23lTOI5vVSJT
zr+aIYBFDUTqSoRH9w/b+C6M3XioZAObui5d7PisfAeLP2rBlTPxeTl4NXxL
VZ4bTvseEjGEpsSXF9zVzWNYdhwEK6DWJ1jgVQpmlUcm3L/GpNjUd+mTpaqs
FcE4xsPlPR8oOydCQGxy77Moz5nujSQ1zmSFIxT0gH/PDNDuQqVuMaLZO7Wl
hGnZYFLgBGgxZFTlDLhKok+47Y1LE0zPVkubFKw6He8COSUK3SdDQTItf7wO
PcK2iGhnpxxHwuNtC29g5qu752USagbiqL/6BjwLuNQU5Kc7zPnb+RBYZqAZ
xotuhe8sWVcS4Fbl71tN6/4ARsiOc9VxqM9YVO/LEIVWCmZ2732TgYEHdNJC
yQnoZNCmDCWtFZjNqRGKM1iuAMAAzqfwoHkUYg5h6xLTw8qmKeBFW1o4OksK
XrG/kd052wr3G+iyCwEB72UaKZ1U8zSaQK2JbwRu6vd1k9K+i97m6SoXA1k1
GrxA9jkUNMMdzgvQdns0qqYt1uQcuOJfB0VAjD51RKTqub9mKuc4aAkHq60l
oViM9NJ3E4FVGyYPFWaup6BcIR2t/iaJD1ELxFcKUHSpEB7TVViw8psqG+qf
oaGflzdThF7tF+XfuU3XsVCoEGRhe2ejazu2HSMJMSjxnp4Kke1azl+V0gV5
GN1o3dbIrR5q740SP44wEFdSz9GtLVmgeuIOohZSi/LBKuozzgqVzM1PTus0
79WgqEQVK+q/qE7HS645rOjXWWCtkB2C3JQK5t8VlQeeApThQJfqfT8UdSfs
M4i54f+R4NqqgIARlT2VHh++3QKtN8IiluIPSPEugzvZiLH5dCnF7eL1tgPb
e0HWjW+nfxKcipnNXcwgfZriHwP0H61DlRp8CIkaufZOwhMu2oWx+g9vp4I5
NAkxD7n496D55ANEK50DfHpf1DPnJCK6geHMvHij0HKd4n/0r/WODQhrvOWq
NBgJdGu8s9hg0dVV1usXwcgpUALuT7vQGfrFQ3qnLHTdhKDZ1PG8qM4aO18t
zqH9696uajkoLfBcIOnDEh+0eVbaOK4lgM0kvWZxWiZJTFVERoNUgxKmsWht
zzQwfwIUDsS3uSvkne8SU34LKfrcF8QM5lFPe0s6q/ocXMMXmagEuG3V4Bco
7lSDJGzLSDF/He4bCw7V+yDvcsAcPLCJc/PPAhGLJVozHqWFzLw0zLfImbAu
SmcuB1cfGGOxxuwQR111SIdYjyB65VOt2UBedBjgYLsoIPTf+Isa4+D8Mqs6
eH8VYcuIs2qsBFRJcJ2xKqM0YYBk23wGSZFpNTBovWOyv46mNx4V+9yq5DKI
btedZS8va0JiBr+LQ+NwjQpdrkdFb6lqRIgbcRv1pPAX389DM5/DtPrzae1z
72pr/+mPqdf52UM9h+6yxWF//pSDJHvcUKv88sgbboxk6QzssB+vInV/SUa9
QfADHZ0gnVH8CbfwlrmBYf5g3bFFifc0em/qUyyolgDAHV3su9yArENfBXnT
SF+kM3p2QAMTzxEY9LcQgfaqxURrBVFOJ+kII8/aKQHQQn8eJpXj8IDzkdIY
ETbr6NlHMWPCeSNGOx2HwrFrFxsXenI02uovfb/3loY+MHPHwqVdaiSgjSXO
TxNK7N8ZpHrEZolsNKkl79Nu4WK/RThNGuYL70bdSELB5ISmvtGiLvcTZE4k
BBddJgrA6WVq7p8wuk3T3vhGESgBa5G92BNzZgc40mYZLAzgS8yj5h2VUQft
LiZjZlZkXWYT+qKgONYGZRUfmKOLG9dixeBMTgrp4ik7/AEwsVufZHQwbe6u
UAc12vIdWRH9KRTUauH1UGXMtic5njsDD9b4vAuJFMxxKkGUGZ+aBbcl9S/L
GFDpg6PiHsvPKHB1GlTpXP2oymCp7N6R6ZOaIZTckiHj2VWYA5ghgobNXwN5
7cVLr85wsyjTYof8l0jBoSOdAIIFevo2b5mQcRDOexyig09pWxF8usANaEll
N5cjqDvLQr2TiXlzbj8SYfqj+gGt2HTA+4mb9eUVthUc6CYiWaziVPLl4hLk
Xz6jCynVfw33YnnnEohAX29Q7DrxrdQgWkEHraVjnlu6u6CIAaUdSnvi/HKu
h8pfLck+JGSrNSqDYXeQH1h3QsxnXkLazc1SIslK7kKD1HGRAsSvrJOQ4sBX
FdQ/M7qi/RiBjsV512gNVVj1LMgx/k48yne2pm3KghHW+MP7XrQ4hnAZ7EIx
u1sH7wOMD829WMxYg8OOffB5f7NnJ+aV7+OX8H5s4L2XmJ09tKrUqGPSbTcv
iwbb/SnWjEyrmCOVGWViSZAiRPZRDdFcQ6VYbXF6eL3yfbVjrfKW468A2CWV
y7kTpTXGGLI5jqvnkBGgByJ06WtgUgC5m91AadJAbz+phrP/6BLq2bDQ2M6W
MUfaPj1sINF90Q85+0bZIT3D1ukcBgfNTXuStPE8J8kvWma8AaULsiEt09sd
ZMo9YcEo85alq/YGRTqylnoM+I1E6QiirPMhuAXVPv0yswTehNHysccA67z/
iwKp9CnAyf7Oa2wqtnVA8dVOrOXQqAIbDQv0dSlF7kGNzUfvTOxS+9ida2q5
YXthK1xJi0cwKUYu3tIshJIDEAibgLzI04eK57MonoQH5UJPKMjH1PuYtgLT
mdDWUf3KHED3ONBpwkeiWa6uBe8IHXB10ZQSTSHLpUuv4s152PoZD4z1Labw
wD0ANllgMjXbimc+Ox0Zula8yg1zxIq//wBkUWl6hMlk9et2m58hWyVua59R
cY4neuhBAaShciR+dBQ+Mwmmnv/b3+/nYtmBPH+DHmLkjr0eYv7nBl2ewUfE
dm0SmgAGCPdB/DrSPI4/sudgU2ArucbMWhD5CN32cwxIT5qHGa/SihzwugM/
Th1ElE5sOBalOSnTzSvalRf4YXAV1zUs3Tu8du831B44UbOg+H8atlJ3BVL+
VwkX8yLylYrKQ/S4ZUdDqOBiYS/BQliMnoMzYd7KPAYd46frCfyhNgj/IzKa
iMpqOAdLaIq7OfuOaS9DTsvuxelBYefXyd+FC6MS+j9SDIwCM9eCOw9Cbi6C
Dr5T8T08CoOvPRrVjCEtbHsAUM8sC7CdtrF8y6C4mcgTfS50nyLCyRdl67ON
cTebu+F8bPkr4IXGJhsHzBYLXogTR+0F2EQah90KQbLXkFWIG4UrDUykx+6B
veWzlIZROrn7BynBs86cjDGDS2X16gWh75qlEBYfSAGJ5bkNng04KpKr46ew
zKKFbF3mf56d8WuLPECgaxuk2ok9Tp+ibZ7xV8Nzn/I3FP3RBA84FgIofJVd
XHAH9hSN1++br4UukrA/iuTByfYb73qvsy3hdCpTTBax3DF0biMEfd+1D0by
uWrYkd7KPOmg2nEQAYH+XH5sh51Vt1YO4xCsF2BWxUial14QibsU2/pVvUGl
VGgcjnkkcESlbd72d5By5H3Ls59g6EQKBHMF8OLBgDtBsDCRfEtcnnce9gG5
3Hq1s/uPdFJ8IeTaNFEkEcBrgYs8OPr6asqbdg6SBcSvzUWzLjvNIVCiKZSv
uJrHRmtoYP01xGQfvcB8ocQT7Ie8J2WhYeuvLfX5f0kwJO8dac5PcGwSef2S
fqevoFKSgkUcfmoOG57eMzxNDYRz1ijg3kmdIb04zXbqZMeTjM+jEski4iIW
MZGzm+w2c47s3gQEi/lfLVUzbFc85i62aSC/d+H4co++VmQUj7/zw3vjCdc3
22SNJLQszBCWKYh32lrlsA9QqpI/dngKALKhuryzR5ONB5HIUsrK+Kq/BuBI
mfIEDisKt4CYxk7AWChvlSDqqB63/NeX3W/as1nExuVHptMyXFI7RnW+qBMf
x5ucnXLsqZl+xSeAFyt1GfGMmC6jZjrlLfc9y88P07kjLlyKDXkdsa62tr2M
aClYHR3qNtABvITk7ZDAzSxERn6XjrSJlbuIJjwQ8Nf2RlkENnisX8gBAdpC
RBDEUQsUqnxyElHs3vTZXJa0BDhmbZT6FcfADf+fYZJdvWGeA9+az8GyMcdW
W6oatpHG8A+SkSaJ3C6SuUxBH4ptHiqbcJA+BgE4IrKNyw7k5cRVKSfiFImO
7Xl2ugwUvxoNvakA81hQDxz8NCb7/dYJe1Vfm5mQIJDj6bBWybM/29A5dwHw
DoESLxTI5Z3marI8aHHsAwJFAMlvlUCW3c3IsU6VFM6O2FPri7p5voJ3qxTd
pc5kAZ3SZXK0lqqmJd8SkCivpzz8mlm7lL00FOS93j7FNj6MhfYRzPCk+CzE
XDE1BZNobRKbJFaSqSQ6bzCGykk9jbeMQuh5a6FoFCXkE8M+BUzxx8fsXsTA
cuCmIsgr/sJhjn1xHMBOVUVPFvT3ZTcSP6Cg8r8HUmL5L8gohYo1ZhhwQGdS
xmPUEcsNLRjZ30RPi4N/JTk3YFt1wfafHra8iLz3xHz2D8NqxnR55nE0U+8b
CRXP4wk8lHb/NPlMq2dFS7qGm5G3euDJJcSB7UfuEE+U2Qpp1HZNfFF/0bzd
bUkkhkEGF+/anlLoCtpZ0+5ZUxRn3p5T5SQf41y4RMaT68qc802o+r00sxaq
qMO0bjtG9Eo/cdZ5lkq/0LyEDZOQBJhlNV0Qku2FMtYseIuembf7XXbgjo2W
BlXkdh2wG41HJi4+vafoFfQAHjdwGGS0KTFIvCpdShCSx9tg/MvV1s0Pj1Uf
0ftPb2p9wd4vA9vQdCqFdUmGwDuZqdDAofaay4T/1ho+649s2R9193OnIrOR
37t58UpHbgOqHmEHxRxDI7x02wGwyVreF0OzhPKPS/MswUsdrf4uoMKRsD4M
PQiBeOwwIwQ8pUZyXLHbSYeVgtSP/F8gYK7tYvbJPc6YcHpY9JiS+tSC6q2Z
5E0FgnEBgNIP18ZR4D9FMXtNzb+5Jm6HRRBmlWbVLNtoPwlSUhYi5Zchqs1c
A92m8AljLAdCswwExLLy7e4vCPg4lkLBJJTaejzmwIPWzvCWUounOuS+fXia
eTf6/iciE6OPFsWJ20opxYsnoBRJWyV8tlsPD2KrYyW/IXhStwU9EhlKiNZ0
d8T6AtSvqy0YjvToqh905uhzOAUpfjT21Y1d4uD3V+wsMtmVPRvcDBVtitJ4
+72Pf92tUeBtX6+6agZZFDOQmpCei5/15y2mimgtFtc+5L8HoI6hGYvJyl6z
AieOUU97UXm69kMXVReKTSamtD+prKFOJ48PolSICQfEENwPNi/ZRfPmwTwZ
ke1NlMuX2pIZ/8z3qgtCaNLpM8X70r9MhifA1AE6kogfJGPTKD5hx3J9ZL7F
HZW0jWt5dmIwtnTCxcEg4T1qXQ+270WPxpOKG9UWSoGCEbkhyiolewAmODZH
X8cvAGzB79h1h3T2RqmhE/aknzS4s8Jj0ib+FOdbc/ry0oPB0CsI/RwGscxw
Q/STJ/FmHjKtUr1Q3PvEhRSZEl2GRWLfR/ZMtCT+0VvGafv1oBaW3hRMmwDW
Z8/v+qXJFDpJpJXP7vmwgxkuXamon3YfdjOteaADeExyqpqV1nfz2E2o9dxM
qGDExafFmzwcx5hjbS6qMuR4oogR6AH5gGDqqcWjCh+rS0K4YJy7QfNy1xMa
7gu4fhwJXmc9RoqCcWA5FYmhR3R7yOvqA/TY5Ml25pSEU5HNr2etdFaP0+CQ
/3j2rpdakpkegrjyS64IvP3pZoz9+6FMHDMeEpnbwyJfPMg7s1ZX8gd9WYPi
vr75nzJKmxnp3M6oa84rnBKBBmp2wIwuNY5L7dXoQCJ9UtDz0NxXq0iNk1Kn
PhY+EI8oseZy2TkSn0vu2s2/CUYW2ZIB8wrY1WTQqpqMpXo6iL94TP1xJHQY
N7UqPzli99DdCQN8GuU/42UT2YBB5bo0CooAkQhzreAFo7E/cZxaefE94g97
uhXzEJ8lapAnTVfe8B5MKzLCYSgBA65Tcpt+uboRduIlVzctsGwdze6uMTbB
ocaUIwZOAt95Whs4xhkHu/u0E4yinfNQoXyksb3Bo4Wstwgk8UGNgFdv1Nn0
3M2WD+XZnFpXL4nYmg9+X8U33Y+WDHUIyc4NHqq8f0EM8rrom/o83R235OVs
ivVIvYVlJbe4I4CfqNGQyiPG2353G1CNm84klZd61CEGlWngz1+LGjgowaSc
GJf2xJUNmWxcV8u5aYuFFbTCujMKKhM1YlHPOHGI4hDh0wCQxPUuRB4U8IyW
fY95JrraDL7odz4P4H9QjVeVhcW3yn2qY1rwU+Jn0RuHupszauBnQpLNQ0ev
LKCac7h+aWKR+zbO3UkUFV29WaDcTTvPuG7oX+aA8bIDUalDU/Y2ACO4gxnv
4Wh5fOCyIBJPI9wwUyxA8gkHLcYJ5w1D6wIWm+iwU6YQJ22VhG4xAZ7+Q1WS
CqX2DLaIhe9b4fFrch4X2VgvmOzJ7CeQ0iubRNeZ1scdL+EbsuRsbQmKTPj3
12uLki4+NrABtK2RjoupQHJCSpDVGuyDQonr65MhXv4p0I1YgWoMn65y2R3/
x5iDqF9Fssy1ejqrx2VesCtFY7YPB2KGeRENy7uVqNHha4XQuiEL0t15/HSm
Ib15367pJpCHYl2IkILMGqRGCqVrKVw8xqU0Uz53p4to2YiUk3EBkxlNvhB8
AX5y/Dk/0x5O/fp+WkGG5E+c1uV24B1GIp97dTFyLkcrMNIKMvGuWwOddJyo
5OPTRrySRcF60wX7SYdx3UguxW3s3ml5gjr/pJ3nDyJetKFf2VhmR6mdH0/v
EbO+Jp9qU/qLmoM/jTqZ4SgHlH/jegllcp2ZSUr7puJ+Y3xS23J+bhkrK58t
HHRNc+Q1BnrY+OcGtnPPPRDpootttiSIwf0Ffgn+DF8G1QhGZ6TKDmMLUyyY
TDtr/TLM0FDXyz4N6uV6ONtiw+3/3CA94CU+qP4tNGY4yEiG2ngvgjE+WMuJ
svxRVYFhBxo9xf+NAtzDWtjDikuNwHUMCG6iOQ1yNiESDbw6CBEjJJNAqXAV
kRPknv+J6ngEym3/GxxDYbm+f4f32doD8jrpoKKK//7FESCW4jVacPuj15QQ
uTo6x4ppSL/vlcSxAMzrTkWqQhaN9o+mg3oZ18552x7YHfPVCAlrm8LYueyk
t7G+kspiBtxxD4QxP+NzK3tEwRI3tf1mUoZIEANk2AU1CNLG8ee86QaTbuTL
SXjNQ1O6eyLXjmIAEy3Ngjp7ArKCWTeAuwgahm6i0D47agFEfvnWPwh6d9q3
XWWp0voxkXmRrCe+70lmOb9WEsz0/CuEDs33tt6NUmutq4+qTUXPY5uX51FN
2su80yqF8XnezmsKHYT3iZol+dGcQ7vRfLqjZY9DhwKPvGWXn0gIGdZho7tG
kvpRF7/hkFRbWZNnSbD7mU+T1jmJUjrIJilFW8Oz9WmYXSU+UCDjYp/uUbSK
TydHjO+z9oMg26CyEMVlMxAW14WH4LOfjFM+SZjvTT69RwE+3PPuI5I+Xhu1
7QOtg+0YJYfHLRJcjJN5DOK3S6yY6Cj8pEwqUP+KhZrzeu4fs7/Ld8A2CtBN
dxOd+BuKc5Q3uS3iw208pgmkXuS3DdhoSHVUkrR5DYc7alZZctPYmK4Al0/U
sSUelcUFirTsTDyx5rjMjQc1MQ3u7ymj1LP96rDVuKO1ob2OtQuMdT6Owoxh
LTBbEY3g0b9f1u8T0IShjYplTfAl5LDHzr9q7Rhj4wJwEsVs6SrLYrrHXDoK
2ILemwE2eqPUC34oF0a34jk9gMgQDe+zqZOUFIx8nIeRMSNkq9uW5C5FfMM3
rEwnTZzsDLV5qDt28E6GnU0KT6agL1xg7YTCXvxW3sOlCMBxbCO70tjaoG1w
rg4UceLfCOL31AG5euOaJBURZjLZ7wqPhNeWcjB4lszYN6lFx5V+K7hBvYRn
DAyoyWpKkTbzfZPpbKvEpcndSKblu7zQQHrg0pFXcClcJVMt8jr23EfLntKt
q5lkyT01p8CXWHX7skZdIKdifqKKxk5Qb523jiCHfQFwW5clhiGUlLOqp8Xm
W0K1p5rOdU7yyLJKH7vDJbu8Jm0xclXmkAFRzo0IHMiTby2bx7Nm+iJebrEv
QJKG1zgzeL9yCCB363axctsz2WXUtxKQqvbcB3orGwQUVwME4Hz/hZPMPc/j
dvSOP6rdZyVUY/bZE7g7MJRL9yPHQp6mc5zMDlGxxbh4Or3A76xHSnLYZtwL
dk1nbZZgWdEXJxt5xw+ouSc1nlkc2c7XqPEpz/3F+fjyYwG1/lSpdPoRoJ2m
z44/5EA3k06hZONr59gn151iKw7lLdTBZHKbWlgsavAtV/GvzyFPUlQ60syO
0mjwVUkis6izrlJwDeBTKmq+2eTjb68MdqgEyxqrXviZAnXqKX/F52u/M1n7
stx1yy35/jg1VrtvGUCFWdm9PSd6PhupM51Wz2118bSNizTlnzhzbZH4XrFm
aRzlP4BAtPngXbLpBW3Oa8iDo1NcBoJQ55tJteU4h7INFQbi5RtBBUpTQzm2
fP7UkENArAb5yEXZc2SQVQs1cD2ph0Z35fiC/K/SBcGielu9bBNz4IqKCyyE
5BbzOQjKy9O4jzdB3sKgPOQuYvHJKJ5Zcq9eK8J2L6S8zgQopXRK9TO73USG
miFL9/mH4ooD8X7u4HA/rucaPcyrzrnVif75kZjCYdXnhQiRyaaYx0MJKulF
NcFbUVYpcuIs9ixfuqcztXBYfMgCt+mydlNlNHLYL0nQSRRJxus1LWZAZiKf
OUj5ee+JEfr9RsBYA9OqwrIMZXAa7VVnUyFHLhViBGnBs8ofJvv1qDSs0rm/
KtwY1ooxJeGVLOyu6B8J6HgMyALYItsfgE8bMhEx4GBuI0PO7xoGOvrQlzLg
ehiV9pduDS/1QGnlz7OATiM4KyCv9CFfNiQUMkM0MCABxuapXZjDwc3aLdAK
olWm+uedDK6ufjMoWHG7e1rr5WcNwzlSEx4WSXG6zV5sUt8eQu97p93bTIJj
RBQ78PFplsqR2DQ7twyDBOuN3hDmYyeYhOSGfanYMhrGyvF6W7C+Dh6820QQ
0/1VNFW7o0w5R7ol5ozfb/jJ+Ue+2948KNwc1u+dNKFWQ3AfmWgHURIQG9mz
Bad1+OBLC/JSLuVFysZzVq4+j7W0Ldmz1fJslUr4cKz18ascuqYakBqwZv2l
ii+U9OESipi8dCWqBss2d/JC9OKyyCLjtwWH/wJmeKBC1WT1rIBOz/D+4UGQ
1b4VZCj6CSAR/BxqXOdEEPWUUAxZJqGSHFFDLg/4rzkhcoIMUzKsYEd9gaXL
IXTj4Jzk0e3IkywCeNbhGGmhS9zDjIbgGH9QDTaeLMcbBzL+wdpXDHLxJaZb
bddugsB3VIuifDEvGbsoqwQ14x8VJGNUQvEnNqXW4ZWOG9tE5RZkyOca6NhN
nnWlco/0jW12Ounymt+PTrspFKc+YL3Pu0x8kYF0tx9nse9XaHPbkOXWTTEd
SDEkjaH8uxdUZYYOcAnaiybq/cl6WRdpdaToV7yHXrMnhwo+oa/FMu4EDWWo
39i3kqJnR/YekHfDEcNKn6AS5Tr3WzLuw4HkjucS5NuzznGi5x4KzhVkiO0H
wMusiLiCee8uCTOfH5yKl9kvJbn9KMnSH2+9yrdUvHT9gmPBRUgPqOKYQ0go
Q35fisVMN8hqWLiXu6LB2xu2V5RcnJFPUS+eIiaGInABGXWoY0DWejbKjBOf
4PvK7ZCniQzUU1qotspMl1oWOxxN3Htym1B9eKj1cmm+0vd8RmoJC6TSEHbh
t05pfkYrDQE8OA0YqbEvQcT7SfiLjnTb32dZyKGspQNMPVSF5VZPGVkBL6/Z
WkAmRyt0oTbrNg8+UdQhys5lMK59xym/5oXIT2qS5rYwoIJyqfFEdTk3Ucks
FAhJfhUJPtb9OHASQkYxSZKGyUpbiQ6v0GWpXVCbPC/Nuha4QZORyee8oDIF
ZY8nc41STMRvZ15cEFyyKxZoBIrjc2/T0cPsd6a18D57v9DOOPl6Y4mUZU4Z
sXJV7u5J8cB6a5Yh8BwZOnmAfk8vLJIRh7b/ewD+QF/mWl0ZhvNlJegTg58j
YJOHoC8r+k9ZxA+dPV3S3G5/jVoX2qQnZJmt/xTaKL3net49XTxzlmv4Qy/b
qsXLvq7cSdxo8rnNf3cyxASefajJKJgSNct+cwS3wFMEWcqmixZ+86tCQJRG
q6rAfPWIwKffaW0FtYpkik8jjNB5fXfEhdYXBVBZjL4vTeIz3Z38++yXCodN
wMgcdsRpmC3KbzN3H5rkDGymDHOfmqgqSUTMK6K7CieFGcv/S4g2Vs6tD61Z
AxbzfwG2mJU975KH7LoMusZBuaAS9h786Z6cySrLPgjWMNW548dCGq0P5ogl
Pk4osRRkiY120JaAY0J90fmS5LrNVp3u2JSL42oDO0vE1akZzAA6pFwNYOo4
HPQYFkb0CulMSVtyc3RPHbDtVMLoh+/keFqkTEYxkic6MObLWXOjpZyCTjJZ
5dhe26/Xx3f5e4VZwz/PGTROT6BFqz1Y1f2RTgj1H3Om1qolD8HO2BoiKOLK
0CyW2onagtJWAClcvFA4RrPE/8oSD7RGbJxJ1vdWe8hFTQtT5qynia8lB0wR
DoZJBK0nAUxqtA4mKQ4RxIaLUDXLhqZimtE9mZ6OKC1zaYUKaHtKnxmFOUew
EEGDypHo3gLrOkXjynK6VbkOjrTTiglB9yRJ3Yyg8YTwIUFXiBnZtXpIt1eL
DQfcB6wS064rN/bDKBs1xPkM8hvCHReRnvR/69iDyzEOeqUFvech9v+hQbLn
cgH74EQs0c8EruFmC58jzlDWxG4OG9y8l42osTqwOa5sNdBVfERMokZP1WeC
PGIcEcSGR4ACWHoe8PiZ4WWJT1DVU0wzlsKuQk+bh4fuhMoCjHG5FxehanVA
xb9m6BptaHXVWSPa+Y54AIj71jWiES56kM9/VTaT4q+5pC3UNbtmMKHfSLpw
tpUcbDjhe4+Hm9gor0BMcar86AHYBUO0RvWzMgNEA10Xp0gUwKXZe5+N62mH
51TdFi1a75lc3tN3XpGa9EP65NxoaBbzKgQv7fdB9PNGkLMX8IZETVtxHvzx
ZuXBfWtIPlEIviJjI4Srub4JeCDRr1KcnVByW478yzUhkmZlmwY1pY2cSgQa
xlb6/H2y3xRtUvOgWrQAxYegMf+Vhua2wLgRP2pCnHMQ1KopBoDJM6D6KBc/
P6zucsyuPbKdVGO1nwitNTWrxPzi9QnkkRaHvoV2yZ2GzZFjrz4/USSvln4Y
7qsDdIrLE1ZOv/SnWONHsAxpfq2pHsIFoilNjFghKzVu1DCPxguGBBYhOzHx
mHC5EaibqRhUQPpdOo87A/E2pqUc+Vkx5ZERYd+xbeFuEo3od3H9f+WnGDAR
RrMQRUUrTR/q9jjQortXXv6alJ9QhtoN/fvW4c5kVjyTeR3EdmNyuPkm+Lb8
GzrVLNRrSX3+whqIfecXNJsyKTkyGBMr4iTwIE2iMitaKskjlMwNZ8ySbA4v
GPfyGVGZceE39LBuWHeFx5tdXT3LQsiWie9w2GX3TSa6o4qlaFmuqpuXw9uH
Zp1VoEKR8DHMgPM9MryFDN7iL8W6MnN70JI8D+1m9tX3YEoZ+15taWztkcZn
sU+vf9rzGZ3NWgcbHVbR/+FFn0osHITN2dZPM1PI4QFxBkffzH8CR4FmMbfe
l1VSg4f6lzBZc2oYXE8P8PDrMXnK44bFhMHow5XIWtrM1iYoOhsJD+zoFoFK
Qswx+f22VYxsYYePbhf26wAgdboPTVSqic0caCGOjaUOtOqVu81r2yd5g+p8
syxcaPZVnDHI7k5H8CDIk5q5/l/+U750zHvy/MN/76S38sFk3WfFBajJPd0K
8r9/aWPrk5AEt9SY7KNGHqynfQyPZcAub6ywMg0ipByRHxCiQS7Vv5WSALgf
EvgpbnI0/eIrJ/RRlMaDQzEm4Szqds1L5PpU9iwsF1H7jhZ+fdDKJIOR3Pwi
AJ8I8SO4XxKqi/jQdql/AHLY3cHNVGG2k/N2N+wem1xfO4BYQWxuQoWTaw+U
nXV/x4k/ecuC7t0viBjyzSy8oFhwuyq+HVySi+y8RnQw4TN5gKfbcd7ZMtir
1E0D2GSXElB5RJSCGwkI6x8z/edDDCs+9VgcztN1FikM+fklUVv/24EyZV+7
8AAu/nMYereSEPUn2BT8e6uoAkaJTxkY4Jxz6TylvqNE03mS0bA3QfkizzFu
Hh0onktkwyCZ41ffPFRcdKeBFeSCNuwahSM1Yz6fGBKpHM/DZI5+vbSXpwAi
PX2Z3v6lkFxcvhTqATHF5O9rwg+O/WJcN0ymxD9hVdnqJWELwEmoNRZBG2K+
PIATnRUX5s/9Qvpu46zn87vJfEQz6hJ1AOLDXXdo31jheGct4lQwEh9D/xxN
wRERX7E/5P54hb5MteKzj4iwAp7LXlhAwXmJMP80aQeETB8dyIBghow7F75C
cjuShxMuN3NZUmqDZ1HNi41kMV792rM/c926KOB5iaT+8hY5jt+3b3R+RSha
XBSkPsI5KtZZRtRSxm/wRQSwhvdbvnvsHJeHkNiix6JnRyWxrMLAI9/I+nhc
aINXUh3KG2qhsortSuV54rudjNjJ23rQwE3EJGMRT49mDP1me4IlI4RGg7eP
qttX+jGuFGlUneZY0p9lwMjDmwqTWq6gTvJfgs7Ed+Ob2sjpJ6RaOfBRWRJj
DCYZm0l3bov6aTFirnbjoi8rImojDMqB8u0PmJ6HHau+WgYKYTQMaNefar/w
4QBvmBZ4FOWHfMQFQLlE3fjQXhs3diySAEjDeLjtJ6edGyqV5zyRFh1jMbhv
4YtlDBuUxrOn3WjCc1V0Ack1/4PsOQsRTOqMF3N9Lmx4U5pBRzkSupQWP4Iq
yNHEc5bzcbfMo6qrbSAL2hvPGDb7ZDAXCkmQsYQiu7Jd9fNWqNNGxoZNMKy3
e7q5uI0kjlQwiHLR3GRqGTHz6E1QYU3MeTAw/jtL1uWQYuxtfdzSCvEAHgj+
8TjYUqHVWAS+Mcda0bRxsObBHzNOLHeIzll8X9fv6bEQjeNqCBirW5rBBqAF
BbDmtbvbHuQebu22J8dxdyertfKTGSOs+7nmKw0+eee6x2un2BOcFc1rSoWj
UbQuC3CbyOPSDQUHkJQIlBbrmz6gu6oA481nw9+fQulxcAZSjPlTyOYajUrZ
IOOaaHegk1NU1MrvDazPuzDm5yWa6Ady+bE0K3C8BqjAjt9Spc8dduKaah5o
1M4j59Y70/jo+wICS0YqMHdqYVv+Q0optLdjstbeffW4PZ+CkVSVjFkPxh8n
TYCYmU3vlxTwLfqjUcWskqJh3P2tdO1p2OvHOi0Xskqk6PCalAciPsPb8g8i
UVyx7kt3kc/p0wHrs3ek5QAEfPD0MRJA4hakB16YziISAL3ZXZWk/V1Hl4M5
3/EM2095A1ugZB8avEHXjemi9jEH5GpeN7hJ/L9gQLXVZ1AAPRZGdoK+ilI5
HGOC2uoWWl4GJnyx2xAthJhAzXRQ2NhyI6xGSteU8vo9l+DkoqXp94UKeHwA
ZOa+f0tJJ9f0WxMjUmk/WPgT5BfBOoISJSgKdUK4ZI6dfeYoT/2m0JlVZ2ea
ZnbkMLkLUGpABKIp8eG74QYECkPLN+C8ATM5U0USH1CsJtZ5MhAK3r/11wkC
gatbpUiJJRt61fmpX757Q7gnDUpOOwnYuClhTRTD5sWOZ4P30wKIalsOR+Ts
crkrzBDob5o9S6bfma66lw9CeYl4THrrNmOyF9U1Vrh+yAGAyQ9KHEv8dhk+
x4tCFp0vNqoBr9ytNWFmuy6Gpv8XmOob2OvndL2wz91Fo/Bc0+u1DgXTGSdS
NSK5LS4A1vkMl9lR5GOck+PwIByvqsyRT/T+sfMsKTKjAEbS42Z/kf4VLlOX
vsAZDrGjAhyuUedjQF0g8kOybKsfPCPDzrWuWL4fEJ0/Xofcw4ebBJ9vjPHr
NoPttfn3Tr7qXP9KvdS7xSPq+v5ETBiYrtiherhVl4BiX/OvC4qdZKaYiT5R
bdw8f/IMYHq23um8oA2EOcNdWYR93WHfFwQC6fvcJWJjvmOe60aYDXHWJnAU
H4V+ISeYk9ESB/L/jKViIr47VwTxGx3183ydkSdsi+Yd4gufMJDzqqFGSVj3
THjn+AG54nbsVmtjkcEqFFgauYQ7hWtMkMfJWXyRp9cgXUs46b93i/siLFZO
a4F/vwTsNnLycW4lprrmSq+kSB3ZORijUX3PkmIAg6tBQeajVcDvIX7KxHHC
Fu/v5UnB6XSn4k2Aox3M5XuqQ0qh6liQ2TyFP0kNfQdElSlyBzrCk8gqZX4n
cR8+/XR66wSPTZE92lZ7C2b1jpyidrk902HQ1smEKzC0JYYoVXUaLjYKbW8e
HMyUJ3c8Ryk+/cn69ja5vwN5ScbbcDH4uwQK0bX1f1jZ8PYf2OKjsk1xKvc0
ItxfjjjCK0GHPemGNFYYH4RxUUY5kkLwgX20kMNg0C0LFiR7SRSdATTeqHFb
JyrJ+ZE6lcMSYZOMn4hxrcr2mohdSoZtmoZb+kVo4TpFLkMvRdX9Gf9uFHSv
eHW3MMuhEMHJYMcUxB30eHy4OrqT1J00DjBIY2LRWyYguB0UMN355pIx5kET
A95QcZX8Z1J0oVlvsGwFxTXtQXRrmTb4Uw8jfKqDDf7x8JfiMUH5HkL33gY9
+V0Vq+fyFMf03i21ol0+ZOkdemXObIVZOf2w8R68Xkj5lvNPslIlF7jfrMwi
Meg25ULyZL1L5Fo4yLwuMUNu6vqWLgMQjnY/6KlngDhUSDU2mjMhd5yv9f80
OeGSzVqIdKWPIxKFuPwpuoB6W0og9BJUdYR4vA7bhLw5L05x3jXYdUqh64tn
4lPMprd4OCUcnCxxSiYVB0uW2J4CioYsjTmWwJVOfAYeyk8Ke44AhpcPOLwo
Xf/ApKLvIQQLrHTsE3iY96McQEckraTKnsT+lCTNB1eTz5IJsrja3+Bto2Zs
BH879tuK1taCVhd5CaEjZEOP4D84m4g5IgwTz+ll2fLo83kpNvt9sa0qtzfS
peOs8UkkcpunC03agUzV+Y0yniTIe3km85sRSavGNi+jD9G5XpGblu8aQCU4
gDmQG9mrxOheZcpe7/K/8nFvlCv2BUJ2Cd7TgEfMr2SLyIwi2boeM0G7pRqQ
NQHc+91f+ytcQkv0jKMXIq6qvgLBMyBPJbacCluRfolhvWJFWKDijg0c3BmG
B5+OBejfGijvOrzZM9hoITjiLTGwfltC4h3orAuODcE7EjTMDwKkEwDmVE/9
qFmiuBe0jNMgLZnxBrfVKKPQS0CXLloYsps6YecvZwfHQWQhx+ikx6DqCTBx
ltQhBYiWizunEdIzuGmDDMTA+WFvPhUvYs9YsLY5Xyc9plg66keHWCgNQ373
TxIIkpgM/JBmSCVcxKv+QEm3xS8KjuJ22gI/0I4BdhNv02VoudJjOeeKtw+2
pFp8NUPTVQfAhlzRTFWHRMMXNSnSk0TPQe3LONoCgLsTW4FXk493MWgVV5d5
FIoNcmVPSOE2QA6UxuFfFNub+nSnUIUNDrTt6X3ImxMG4wQQ2T66MRPmD2s1
F/rDx9KXbc/KN9XjFRJepAtbq9U5V8VADG6q+obgSr1p04GtjFmRRAdlVZ2p
H1lBn6zFEChHtfbaEPSz/Z1Ci9s+vaMIpJFqUdYfdCCRpmc70qPUzqGEryf3
hJznpVsT/Da31WS1VKLVzbeTFjdCRWVbh01gsq0EDxEyOOz1Ngrd5a+3jh46
Ak5qH7N2aUv20rgPv/FdmA8AZV3xRJh+VbBaj0Rqyd48UaL6HnQUeNV5NaWp
TscyCcNU42eF9AQWSofiYwPOLnFaNT7TmzmgBqLy61V9OiakpoJzmYagSgy0
zTGzvPXaYVwGMNIgBLC+QTK1nODrYhW5u6uWxpb+fe8FfBbWaLVs5GvDcmdu
gLF4kYqI2llm3ch31zCrQvNAl/x6dgVxJElasH7Fw26WeFWNSLAYHA6V3iYy
U7Kh3wMScurPhoJ/LVDiyYtyGh0ra+CAFVhvi8sc25wEyoxVJttfcl1VlVCS
sSZIT1lFA6cYqKFS9AtmxapLVMPDRy/zmoG51nGlSPgcmsoIYJPP7UvV45lW
+4xBmOu6Q7ER3jLD1DrwPmplREUQq9435QpOntRGaVyCbCmu1iER4GvctIYp
8B3ohlreiRHQ1ENDBqbVHAQ9koKsWLp9gVFkocVWCi95Y9z4TNGbzSoMhSMc
Yu3WsFYaDHWemq21YF8icw1w6HYXsc9edz9dCGcozCozi5fOHCzp046MuNIG
Xs5FO+Rh49mLKyQ4gflUO2ZW+eRV+ABq/bKKqbVzcl1U8qzKeBhW4sg9zYSj
4yZwrd9BqTJ641zYUWjhqXsKthB9R3HSU0VaPQLOgB0O0WhFzomNAx3UIjoe
F20/oFO5aML1MiU0DEhlDsDJ+GkoGPsIfN/IqcHJpGAvRjwhO12NZ7q/0oox
9a6wqW2s94A0mdbz+G6dSc0Geqlepd0iR3HsecG21oiIjhePvfKCeFhkxWR7
QPcn5gFCehxSkJioYKOwX4wM3zNHk+n6pkK1rz8qpeV0eTp4JpczD0yFub3m
IfO0AJzPN/LjUF9l+TgDvmQH7rjAPVz0XGO4pKlS9zClL4g5pDxYzVIEfunX
BPdqCSrRpJOrYs5f0fbUw60u3gPtLNRlkxwEYwhlLWcqU4AEX5RE0D7sZWIo
3U76HhwewSwKBbpxpqTChFz5mUXeqeRayxuNuo3f0mEEQ0RqsSGKsv87w2aV
oCwLk9+kokONLMkedevmHO+wHQA+Akpo8vweKkN83ujkUYSq6VkjQ+Ko3foX
QEskLN0eLa0jtdTaC5Lfc6WUBHTrZs0pF26ma744GvKETjY+4fOwL2UnV36p
I1w18HXLWBHY1y8gqaeXfU74InHOUfw5ED8lELJRcdxjItv9lNIeeUoK7UAh
PzhaTXG5JfcI/7WSJrThT1BkpNy3kI196gJtsT8QeIvxVtNq/qipCGdDwCMq
nztGeLyjZMCydpCfGdPFioS9MerFiN0sju4f4IXjhdHFX8dIriZcDkCIDviv
7utg+j1Rsb0d51AymIFXQfohVnAVjz/WsM7pSGijd3ZiJ/G16XpgpN1Y+CDs
tLXHumTktEoLLDZQR1atKKR3auvV23MhoP9Nv8xxHvilrdV0zZvi6MQJFO10
pDkMLfWhrMk7qz82IOPGqom4gHetwLT10OMaBVIP6qn77I977qHPnVK2IAAo
nbmZUk+m4qA5xG5UKYiOcuUf9Zsnzvt97vXZo9XQmLiEW4X5WgnTDJcvOnpG
bKf7yNt9ZXjz+KYMPhoDj/g8StTmwaYSAxnCpnp15c98/IYXTL4NlE9EtDad
xiDpVG72teq1s5UujzMWIEILnmsSJlbhq5bw0OcyPrSifOozvoqe+LIu+yoC
BRsw2X/VmOJvvwmd5fEuny2Jc+FZz7jiNJBz4foqSHzgloc2VFD5P/FJkw0Y
gL8Kk2zjh824SvFmkAduGcmV1OGp2E5mQHoM0Arruu948nqeSVUOQuOgZ337
KKjDv69lLWDJ+K+uu5Q9FvZEi82a7dC5vQpcHIgXRrdYbtqCbd6fnU34VOJL
EGPnVjLIx+vWc1BFxR2U+KRVp23pUuBZP2UWKBQPXoLs1mAXruY9tOPyH6PY
Yaqy8hnmyi6i5GhrG1VDnUHS5o933zxkN4sND0sqkJobe1oOgwftza/Q3boV
tN7CzSUigMdT+y81FOFLWJ803UWpALFcqnUJrDqP+t36rSKqRWIz9I3eC6s6
bAxzpzVFanpHnuIuU+4QbJIlisZpNKd812sd8lRMi5SzRKONDWIFWicLnp3f
dyoG0C6Lho0mSPbC/xfnx9nP9EpPgDefxH8WyK2YU3qNppx6F6xDd8uiphM1
pW0e7WIHMEP5UlVxtYZIpX8n84mX/h2QUJET4TvDM20eOvNkxyx4WEEe+EyJ
n2rz1UJtCLO8G/KolANqMlRqVbutks5hielegmJtHQQ+NptzKRj4slGm5MLi
yWXbEngqx8znclKeHoxpTNcVegtQhnCPjORFKDnmcV0RIAe72FwtN2Juu+mk
i/zEEgJCP47UVewvDTiYrmEzcITQWGMZMaP/5QJynjui1IVvw9LArPckULTC
TwKzBd/r+TsJpLIwLlF5bMNnx7KOhCyKyR7X0HVEiXSmo8gZoIIrro+6TNho
YScKFEObcJJQjMwWpP/O3qVFkNf2SCHctW7BwUnouvlNQsm9WO6blm3JjUSk
xXXxaPeMcZqd3bCiyM7EmagTphy4Yci2u4fZBqV6ydkO6FkCDdR8W4cVi4i9
9rAtHsSVBxKOTaIjmLvfZ0UjKljoVG8D0z5FV6WPk57MLmcouvFpbONBmFXA
9uuny4+PKb8E1Ryr99Ug4XwPsA/hAikrQSoGJG0pLadxz6iyLdtUBLqKaaDf
SZcz2lahlVo1htBlbahrw4QZ26eW5RTAoA0KkJ7J9G0TjVuHlde0KXG8p6cu
TtoLWsaMYPTWPwm49f0Xx6AHvAMD4PkRjrwVYcMCYVvhzPQBGMz79pZHNHAK
j4NtDwcMymo9apxh/42HeheXzVwILVhWcWiK2d9AGbUPpvx+K4NLPN8Uff/7
6/ZkA0TXRNbYYCCCfFz2h4wdYrNLgJQiaHIbWpQBPtGMXJf/3uXQREvzxzFa
8OFbbME5ritI0HrR4IKFmQW5mGAzoiFJIUBc3uO2cwmiGDEfQutMaU3rzsHo
fL1alPRUjrpknl8BRq3nv4ln/fEG6FNyQugZsc5sVhOmeEaTxMsgofRcdz+A
ApW2H7+0rNbloGaPfMz6BO1DHW81/4Quyxe31T/GguibSfFGv7BMX37E3g2z
p0VtlCZ2O9mCTytjE4ZnVpDgnp2AbS0Z0lyoFvktsy4XiVVa4uznu1cP4m8f
D3PPmgooGhe83ThCLtxWGcX96bval78L12hkqqUy+HU7/cFc9juabOsW+rDW
lltRYJOGxUfY4NHH0IHf34d60PGMoCc9uYOm5AqTNiZKmcVYQyu/A4sCJHYT
X8ypbZwI4fi5R19NG0fS9Jeufc1QHSR+9qVxoC7BtGEhpsq7IyyjzNQl33ae
xafho7fM+7OjZAJtwE0aX9pz9LUhPW/CEQ+GYFkzGjIcRMnVNa8vnWJPlx8z
uQi7QPdJgA3cLXsYHurvi6dPiQPHot+3n8V2gEPuVBZgfUAvcqGRpMGkJPRB
G9P4H2ZkWrwa8LkBZHEO6ts3JGo6YwejZKzFLrww0yI1E+CysS0tH5BkS7Fx
K+b3gufBTAZQ4Riqcs4E+rwO5YRVrpMLTLjHTKw8U4VqeJLRbPdleHcjGmv4
Y3xGLsp1FLe1rbWeqihhWRNLn6TFhrwcR0kWt8CegixU7LPRVULW+rYnK8uF
FibIDYEbkDQbrci9GMzYSx8JbAPi99JbnKgp9NFHqclM4MmtDGrZDj48+kEq
ALKhhebGatNbWs79/7mY4mFvfKxY4wSocKMuIgz5ZgvpEYHiI5laz0B2yGeE
95G1Dga7EfJTTVZ9XB/2EtXKc3JPTh3yoghVQA0IMeyxhmha9Kn3L8AaSMQb
74Z5IRfx7iGHmEH9+NYrLF2odWzqdOl+/EaNno/AOIyGczbjLaxJoVjT9gMz
ZsHzWfpv298fCZyUKz3PIYvb4glx5NHDzyfNn6crQnu/UGKv88M2Z1CCTSJp
qMHM48uisMd9p9J2ixRXpokSqjUiik22+wenstfqUl+EuEcyZ8BPz1vr1pB7
oW2V+IcqKHlWqrfKSQ/8VmlVFEkvhDb5Hu2U2g/w/Z/r29V3dTYEV+YM/Fkn
VJYegQt6bW9Pcm+DxM3ZRcxdsifNEIXmoVbbpLlCvNCvDb2+hqk0rV/jZvHU
1lGq+jtyxzbrhdTixPAhPNywb5J8DENnV8VhQV+Xy9985RG2oEJKjHnTDK0W
BayCnA6LWFhVuj5j6bleNi5hqUDuH4u2TrX5CiH5+QuCWkc8oehWiXy80N/2
OQpt4yG3hSafsVjRPyahnuYOo0oseq96WSV5wtrE4Js5ArxEGR1ebbbc3txT
Oz4+Ykhjf7S3QBnb9QgCleu6N+UfXWDFDo6GOriaLdwbAx7z1z1HlGwKJmOs
MT9Ii9rnKQBiAZDtasUZ+nxLBqKT0YUFLzf2A/3EO9oDrVtgNsy6ePCSA1fJ
c23WLq06kuRmx2MqAEgqS8EG5piOLJJo/duq2CBLpc44MOGr1SI6A/UGiVUz
dlfI4Jbd6/uKUic9Y1bZxy6OLwPid/5umWZcGtCyaXIhWdQJ1IDPC/KRRThZ
XB1te1F2VXDum5/8DGojjMaXY9/dhKW9Pn+l27cW4CfhCaLYKdwtxVZamNmV
Kmnx3owrphxvV2U7266QYlY/rJvyxB8E+GOhlLLkzKDTmYe8iKGngC+pc49S
n4hSkXjN/iD9s1meHAovS1Y72VJd/yPtziu0AatCpMBJ72t5PemrtMEzBc1l
vWdI4ibZM1U0X6+Mvl/m6fPxuRT+o4qQsyU227KLTlyUr2MLHlm7s0uOnoZg
W6ZS/YnYdSqLMZ+sYN5FewP7StFgjK49HbghAv2G3XzmgdmqP/bef32d4Hoj
8S2hya/8FwfuDoeEZ8Wxj69p1AXsxXZPzgXUl1iRmTOW0QNzo+8qGK1LA7AE
NHwrAqTD3ZewNFe7mkmHjoEuRsTuH7cgLfP5tOGqX/okKMOsKCdeKnVmyx45
ayDSPnwi437YM7msJG95IYXmyJkdQ5fypibvIhx0Tw6Oa/TOs4VmbsCVjfut
a3LedVB1Ud5oaOd2DwMKKVb/NUBkV0KPc3uMVQ0WUhsGSYm/yiY2ZuanNp9h
ZtqsMJx+QcGBIPf23RTs7x06f2GTG6MLuOrm49pZEs/zw9fWFcT9tSIFsZBO
C57hmzCtt31g/Se/Dy9ehPfOgiZfVOcA0oPwJ44sOS/ZnFXjIerS+dahnzyF
HZxepsN7d6B8CJOkWEFudCp53pRESLD7wLgjv3NaqCQXjDT5lzGb+EovFRoy
DT+xAv8Y3o6zFzIIWaAfdns85bqMkjQ68a8kWfEGdTs6efgO056qKQipLSmK
GmV14CVMGbJL5ZIOjPleJW5+u5giPxKTgwyR35trNKxgApQ1am0XZx7HR3dU
ivpEFjPek+YiWwtGkiv9Y6Bdwr0wZFRvomAtA9NNnIKQOTIJDO2njqBKCnes
gtlmQJZj6tMChy++rIoSCNshD0T/JWEf+c6V17M4/7Ty5kX+81vpTNwBxt8W
GtU3ZMy5G8DSDPJ5Fgv2VJ92pnfDYLVS41QpvYmc0mw28XTearYVRVYPkdPa
Nn7tQfwfpzBLZr/gWnHZZBFMS6FPz4e/rS2l2bocZJPBb/Ftt+WNQdVEjWgU
t25XAJkIuw76GgI+UB0tQHuGMWA2BQzHrYkq1nIMwIpRWjWvF8ImMzZGuFUN
FMGaLfltclwe/pJ10iyEIfs0VuIT9Ba9X7EPEuWJpBa7YP9Tn6s7f1B4iWoB
8jeI4VJ+kutfPb8U7Rnjc6YP/DAaDu09T06xuQUoO3klssf+TjSEjEo4yELO
sUO30h3Y14J1wTLZ/0GnePLnCMO/yhKlOy/NTUPfIwq3zmzq0oSPV9sBzEmd
BuyQrenfI+5iNRadY+r5O52BGaZPQb4eCMy/xXCL38udY8pDvwoM7C9DHEas
u7JSpow/nLdZB+9ylYwtFE9J+zZX/TTZ5j/8geh/G9tac8EOMUurgfXyXSEj
Ol7D7eZm1ERVaMgOAc0xRtbboQnWW2mwcw2qU8LAprpIqkLBiITJQcDDqY4c
5PiUmIehh0WcYbmCfeQWU0qp8mpO1V/StOahoouYbVq4M2eC3/VKkYdwoD2r
0IikL4SbdAZnUZuDkQHVKzPCDmWCXlxZOmW4lx+5oIwO6wch36W3Ljdr+0H/
FPid5RzHWGJqilsx1zvMAwxOPMOucV/LWEwLjHOn8+JmIXSABcFWSlSfu8BX
JGw2mJRFHYecOO/sn+iOA9Cy90HH1V/RkjAc0X4SkVSV4exOC0tO7F5bs5TZ
iDlaPXV1qwYSr4yb471YhlKZRz1A/cbzfNYmDOv4Vjkb/4ynH1xCFaqj9ZeM
Cdb5jKJVsgVpgOrMyB+c48aapwR47UpIQ3FMPrqB1BnJ5atyJOaVEj0YwRfT
1db2imW/KUEG5recRXoANygqwDC1rL6kqDgtfMsgN1Dmt0E8txk12nT2ZmPu
BoLkXEXoStxeooysH0npXxdwzUT7L5yDg4uEUSk1dVUDI5uTPBCuTtZttBtt
CpTUxC1zIkTlNl+3iuS/kRC441s8/WAW4Iqh1G3Ftbk5h8qc4I9BrArxM2CU
HusWLRFGpsPGeefATOnYI3DmKqdqPLgBK7gN3evgA/xgDOPb3ZsMOk/ekuSH
O3BTEhR79nnzAmEXRHavbwkaHNDa1jHD9RanQDu6NOuy3LQFBJxF9xtYP8EM
ogqWalWSTpZAZ9oLblquJzQJUACWTG1+aAIBbEgrJM0QVxZQvzkLtvo4ACcd
3JfD8446t4InmDk2Fv9hHuY72PMoDfpttw67kNQx/YLaTXJ/qTn+pU3c4eWi
F6uoNgqvjDz/gOuhtOeHjvmBpmEWR3j3uMX8WXttjE6rO6+5t0qQ35mU+J2O
57DqLgkDXkFuG09HmiW1dl+DEQezgWKeNnSonfU8PTZ9cNYzOMvmjWHNjEHU
ZTXpIy6ypZh3El2N68tzV2FaU95Yt9jMwplrKIGnhJjfUyB+DnUB9jXHVFyL
eLia+vNefoI0FmZoyVElj2v8FnYJeXrLZjirgrIlG+Uaherobf1GdoGqytR/
B4s1KZpekB3KqX7jQsEkm3zNPMEpxOo7pDc6HlLwoQPqeyUe6VVc143xSU9m
y9+utq5CWce7ufNlEqXPH+V/p3/yLB7RBnvhTXI8PhlZUgPGe2rrMEES8wm8
fbRE6TVtLxV15DOQ8L5vghR+39RvGAxmNoN+VS9wyevCQ5WkOfysjDWoModA
JX+Yp3AaFCGGMJsagRiUqbLlgqiNcEnrEcY0DhjNdFO9o2EgVcdTWk18yJjX
beF8BaGNMa9riNwj0ZTZFiSYVMyixfGwHmoqQlS2TWjzoKjQTfDHPYhDOvcw
K4fCpl1aMRR4YWEABPxzD+Ad9BY/KXqhjZ0k32oFysdG7p6mX7m/Yvh/dCjw
MjHq4bBuOMkv83bX+nXpXaaRJIuFCANnIgbdBuHdDZUgoR8EZD15GGcUz2yO
lTdJrR6q2Y6hZwWIoxwIooVWL+zyFHHZ0UhiTH9EixkYNO9SD8zpmu+PqTf8
mN5QD2l/iyCz3AjQJ6CmSvWo3AqgIuYYYDt9xy0djTexY75r9quLZAcSdOf/
jCUAAEaFs/AZEhyjSBSOxdGmuwWFCkPTNWaKXt8uPqF2BwUEFj3inDRJ3yls
OpgLf/cyr+9GatY5zRMiicy7z6PNNaVKOtKS+fOHQYDCSlAPLZjTqxxapIys
hx28A5s6xcaVzqjtd2D99lDrPzM9pJyU6RgzK2FF/6unE035chc15mTTUKyx
dUnGtzn/+Ue7nv9YX1bVV7iSli4tPv2iO+YYjybQltJ8UXPY8iTqxHBefDEn
ieKaZW+0j08b6I80ep+wSXoYgJCKx63TDxwH76w2SX/ilTJyNiCnCm0jrIAw
dNgEQKGRCWBVbtA3Bnzu1QMeqKRAbPdhscNqCxvFESKxgCTVzhRMtaKEsmaX
AVByDMUcxW3AR52oymD4M70XALG/Lqy/CQLGMvatwZir8qHRol2/0XdjGxOU
LTyDTdB1oMaFpa+Ml1r32BfvSbUzXEppBncK6RoGcynSZ6+aaR7Q0iLVKz3q
g6yzX0fi6jYfCtWpNDhaAa7QhuGnOVS+k+PdpHrbrsv/NwzrHJb1+Y12CZAE
GzkOtDPAjXoWr+2ktWulfY3hxc6Gl3bd857K2uEJaKM1rTF5ZhN00bUFeVxT
jb9L6HB4CZRVCmyTvorPYHnXNCQb6eMiDuE2kRyb5LM/L79pxyIT+PqLsqIr
4ZBu3fvtBLPMQxhCs4u2nDUFnX9Fbpiozs1n6aDtkJt/PgZM5DuR/IKiL/j8
0Y8LWk7akSbQxts2GQ1DSOw3yIP+7m3MlsQdF7GNjcLrAtJIsf5NVSR7ps7Q
5pc7aPvn3Fx1YzcVOoOlsJhCfsqO/lspnZ6uDBfxe1ovs+wWxUrMMFwm6iIc
xM/MQv6vTjmOVHacItMtU65X8Lfwx8ftKPKI8RmktsH7XPCBKJgXpufyHLEy
EcX8tDKaR7q+gFqNatSNzB/XaaBcRKh8mSkqgCgVo2D5dFTzZidLXRDeuwYb
yXOrhsXV+3QCb7uuB6HN3VZpqkFPF5o8mRE8aQHAn/1QAhPxu6M+t6L/+ng9
GKbfjKmUofJmZ2GiS2oeXP1trbZ9a0qlbU2q0txIkHj043QdOYLJw43TO+oD
hfqX3sEuV8onMFwAt2G1BK79Y/9W1jLnhd3Asb3BDHCiR6HHfxNAEvqBggAE
gGqsn6b2/enxdHJ9hta2JDp2RfS0LVi+EWr+ieaAZIQY2KgJlKNaFjZp809R
BC/uS6ce8k4qdZuucfvV0Pc4frrqO95jSJpCJQbCNmjTsizf1ncjI+bY83ME
lbRz+IyxJ12P8koF0oHDCvdZK8/XG0kI1R02EWqvSHm7tt2bggFGffxmQzx8
eoQ3UvTkAXUYf+ZCtf/abCxBL62nMx3hf64lw9f/q38yXyHOIB+BU3HMSbOC
23KtXTRiN5OiAX1G7QMF+FACFAxSgcwWAwVfJr9vdX6Xwrz1wcdOHZ6S+Mb7
OtcUVTthnbANPjo01ENQcUR3jJzzAylFW9a0B2RYv+EMTQ/iKIS0Z/UjlwTk
wnwyItZztnNZAM89fRJNjKODHr7hHRzf104EBt9BkevRPVWIETEZR0Kh1coo
rwIdgK8Na6UvVOQwhV2wolpOpWlCTw+b75oexAt1Om2WNchaMYvHFQ3+hHk3
ExN3XLnnQxuD+6Fsu2SCTDAwq1Ns4jRivhO4OqvwihqZJmWu9H4eJBwSjrXV
G1lFQFKxunnOKghhsx2EFQehbxa4+rtsBhUM3Z25QX9pFyBabp7Wgas3mLQk
YUKpena+lfFNiZfbzXGD5NdK0Xbt+Pqh9FGPQLGfL/SlrNDMswUP2Gqo9jkS
YdF5cF+igzfKPF9+LHaK7X/MtxYBj0jKUi4Zjh2aDgUgzFP8DMMnM9gZJNfL
ZrUlKijEAbI3UJuqlE4Z4uC7XsBNdJoDZP1ds+qtmVVhd+CTLQ/acVkJdQyb
bnRWLOym13XXG5+3Fja/0ExsTqDSmrf0bD7hMKaaIGqZ7sNd3HemYMIqFjly
4lYBQKgW2TLsEhgstIxUPEFW6XAn665sKMvuEl0YOpnceIo8fCfbyM6vL883
K2z0Ft/eaOQmT5hkCmQYeJrYaFUkEykECflc9An9GlfkwDJIix3NeJ9ZCTe2
VuKfpTZsmwU44JMOoIZb4RmP6JCRQBw0uhbtewpUuPRj0wFIFnHb3TezfLI8
fWTwdJExTTMEt/U5cpAm7NSG1KkTaIDu9kvob9v1Imk9VAfO52cgkXVVjCch
5wlTlAGSRfLY+ejQQryRdxahA4IrhaXScRokAh/fDpzCWlqI1897SksDLIVA
PMLpCsKvCzD9CL62Bzmo15Jjym2smNzZX9bENndXxBTW/+FyFHQSJ/feyPA0
s8dCeRpr4n8irdd+42Ji7naD7V0FGUptNiXSE0a//1+LKaKt1BDQolbMdxkS
JnYafYstu5SPqicoETscq6VRWZQxMtThiK17P9PcFpRJ935msEKu1+vxkeUK
PKq6gqk3XD9woHrBQisgvRjJtga0XgxfCvqzk4hFzmDZWmn3NFVRXmQw2e38
Ia+uYF29l4wyDRwq53d7f3wD0CmYGUJo9oqBnQdAKERVMqTXE1WOYN665UUE
Cv0d0G5qOYWzwzaOfvr99ikCfIsEIoe/DZHbRht+jKH32UOpA0wbStjRIA3O
XTbRhvjR2K/NgnAb3Z4BvhRL+P6bwPDFOZIhqMwlCeQAhF3bzdWpmNoEi6uR
dIk2g/DCohtA6DabCXD+P+AQUpxGZ+IrMavnisQxCmBm5sKChRCxpET2O5hr
BaWF7R3xSdOf+Akrd/utILBi7+4/eTCiIWRb48mrSxi6W1Xq1Vx+bQmMhOov
8jG5U1e4n0gBjojBnvR4j1GVtwrS+je/Np4SSfwtyorhWHKmRRSoBgoZAi+1
5RkV2ke9obhfP1PIM3WQ6lUnTNA8t1i709v0vjkhx6FHiRd1Z/V/xgAffw2c
8t6oJzpeRhPWggvHmp3JiFyXgCyYfSbBvqoZgKjpbg7/ej8bGvKaIZbh+LJf
dkhA/lyzpoPHUBf5JwkDtMlLvhS67FjQvU008w9yX+jccYeOfIpOIYcQavgN
F98TGjA+uqpVb8ofrNAGNZsaaPt1jAGVjQeuZ9ytEqhkNiKWeTlR3bYqDKhA
PtBvnqblMoJLfzrYuzJRFxy0jpX62LzbnudUwTnyAQ05TcY3wvERtW6eyPaH
DWIHvvOh0DC0+oK8VRgI2iQF2Sc4zh+dlQCMGzNfabD+CgH281DuL/uWAavd
J5Ft+4yd6JGvHrNlVOxZzNpKswDwTSxHM8xrWuaKlYveT4bxZH7dnWm+oygc
RKKOKOb7ie8GtnjL1zpkGbQWHbL2NKWVvtxFWiaq3NwVivXRjbYERyDzf3HN
xeuD1lWQ+V32glDttxQgBkvere81O0zrzfp8KrMkrWkXu0QJkMhuVu1jgxNk
GE8MgpFO3xW+LKI8fDzAin4VgWfAzZV/CRbi0VDPau/V1H7bMd9OEn0CjYUu
eKeC3x254fbqJF2/SRQrlc95DKfmfGoQ9OSGdhofVLqOFBn8bLwaHBIGQm//
MWzwJvZVi68JzeGNX1YAuzj+iBvBc3j08Nnig2DEQVmnR38HfgQIdyYC0gbA
TmIEL7wsJ5FtfGjjcBh/I7pTycvznt6zc3662h5OmnVGHv2e/Kip3erSzbZu
LskHuUF/NcaRzpOo0DUJlNzk/VTmnP28iDDOB7w0Dyd+hIGGzpVQ+EMA7x0Q
L+eaGd7qwG3uUp26aEXQVoMdrZDiHVNZAX6EBn7A1eR2/ZxT/Z4RUXhaMxIO
HRyYAohPkyAmU8WjmoLhOD6TpbkXS5L7cdTW17xs+n2pLHQn+9eiRIpafBgv
ERSjmmAzegafdsqSB1iXm+js2RPjusU03qVypA46QimnqcS7Lm1XzP4JCnk7
qCUegWBQGfo2gOhXCANmssIo4VssXPYe5atjI6W19a7iMmY49r15w4XzSO/I
az5mo1hx1UntkTP0GveI3/4yIjYMf8wW0McqLOlY7Xiv8EwCIW7UzXhzFxEE
0cYt+zczmkVUbFILSQBCjmYl+GRiSJK0eHCazuW1o69CCXuZ3AqR9DfDr6Jm
QoTJ11LchqcDD086p8T1/qe/9H7OJTvKMCcEIK36KdqMaBEywe+ChTYs+iqr
T826n39Zi29uFWSG1frL5/ApSUxj/vvejhS0Xk+PALR9rjwVWSAoe2TtsVe5
AskCWv8RIdbg3lBipVlrYfQRJFGnJzpnDqZ6ZcePYc/AYxD7PU005SBzpmqc
r91zBnKXB7Im2g7XLKRk1DQmoqV17CiAmdL92YBZ7DkmdcIgMPUHLruAFETe
9EtWzOb/er/QLJA/h+MC4Jj81RD+9EoQrgGSZH4VIoUxQFRqI6Mf73XrVW0+
5QvXvvBlNEwDEbIn4iE3eC+oWtOEo6mDzWeNZ/SwuP/uRdDW+9x/r/RhWFk+
4wkz2Qk+r9NVN1LjlGtp59+LUzYPoGwzOOO/ti+WAOoISP4OkwKViKLLvwAX
KkepC/bCDJckqFHtM7r+Bv4ez6pgYblVSqYQwYikWFFU5O3qFOeQyKi46a9w
MCahB0f9c/Xr5BiHyWTFecTxJOHzV50v76+qd1nAK3tCUpAcGP/UjZKJcEEK
8iMLX1yJgcvngnYgClX49/qvHieyNRmGULFokfH0nAj7IkHuCFS5+gRmtmf/
sUaefl1C87jQK+EUJyxjv6c+Mtd2jenlOBYdiwNi6YmjBTzCn3S4PBdm9N8t
3gudLZ1VP7nxLpgfJAcCE9iGNaEv8A5oKMbwAoqc30LLd7YrvBs08zvwbGOk
0XAjYIGOiGRLrbLfVa4BkgfpadQwpZj4avCChkmc0BmIBahG/SIgXsZch7Kd
c6j6eVb8EhLdnN+WiEO4Nfre/WlMxV9v9UzTNnDUzmrMUoFHON0mnO1szw4D
PekMSWknjdIPPGD2F84/iYDtsyAh+rJ0JfWvTa02dyq/XtnlxdiD//tOqogN
R4nnLymXs5y2k6Nm8ORsxzvlGFNggHnxOao0URFWiXmfbeQSkehJOVTRBi6M
dZS/QUBsgueuEA2W/zjuc6LE6aco+xDb+vBg+c4w2ejHkHswGCF2ERrKZv2b
WULCCl+2oxbXEyz8+okpTxNA7ALpYMdPLfjKJQzCGL8uqGA+kzXZv0WkZwwx
Y0P2iHkh/eTU8okFh88MIk4tgK7r+fz76r2EFhu23um4SkmMAKohXxBDGBCu
MHTr54DSsJhHvPrMnNGV24stXU0stkPiQjjSPyWJQ15LTl5xY5bkaAP1lhht
kSBmMDyinp3AqlYJbXTTvReaUMvA+McuI2tPswgvd+K1gBNc8JyvyxYjEyes
4lPGv4z8S//EOmBwzlJax3K//q9iy28PXDWjKxgHGJXTTBAEToQm6l8Opgpe
MdP9KN8woHTL1eELEBwK9fBUQbrxgkQCd/TIMHxDpJqQ2SGxXoK+gR5j6mM8
Q9SoRyRmcurp+sn0hzXNCzh67HUSfpXnfcqJzX13p7lYTtKwQ8L8i4Z0FFLQ
b+zxoPQF49l2C9971Re87xo+a6KSj27R37gJr6svVd9ogaxysYHOXtiXazHy
uxMJzseRdD0Q2/6ss2ms8dWl7fKtRqClYbpFysHK69zK3WNCg0KgcEopjXiN
3gLJUOvSXTGbNcY9WekfcEMRdl6t5jITLXsycOMyyZof4MUu1jAQaBYqhBul
OmtlRbWcTboMb2v7w6wBwjr7GwI8yfxDzc+wvdk5U5nNaztE2t7pYsPBOIEV
bv/Kax3Z6jEDSufkbDWP5rCzLkULHOUvc0fM1dYcmZOAIJfuwPZ59Ey5ldis
nOjXjGYQjqBQt4mHTqzomyo+CEB4RE0FrvxVjijKvnnwu9XpAzta3LdOsIOq
8YX769cjtX115tSdQ8WapaXDlTkHm1qFRkMDa5qONDOb44MLQ29RhkNyUazK
+2YrsXL3UvW3VXCkZnHLqzsw2pPsn4j6y+3I1BnVIdUjHwjcZfKPxHybucQ5
pSCqnZZ3Dh8BXUXO1dH+TQ2iabY0d4SvtuiXqBWfJeAdBEIOiY0nBlRDszWx
suMvOmKxlyFTR8nMyQfqOKkQdNcA2NRrCT4+9pJbQykUJ5S9rjn2Jd3R5rTs
qfoV/zv8Huu+Ghcr/9w/UbFVR8Q7i4ahD0XO+2/5OpZaqyXkAPWH9HC4S/6J
alO464MFHVmfZ6IfbMz0zPLY3ou7TJCZMHlrTBlHxNUZlFIlVVKdpxHPpYLt
JaOuJ5//bv89jY//Zd4WKZP/KwmAGpyY03a8z/HXZBtethOGFb07Qj3/z2T9
WSBF054bwSlLJ8da4NmJnzIc2KJi4PRxptwfDP5xOfp5ocs5bRBaGLLn4s/m
LAkTKU7Ima7K1nhHZ35vUU2yHteIkBM2N8PdQTatGKUSEiGaA9Gbaigrcyfu
ZkffBgmO3M9RR8DKJd7uOBRuBsl7VBFXvL+SaqJeoILOsPEwzF0YRlsKtW9a
HAhZLbmyia18YD1P9fjwUFstH9H8tIUDD+4D8zauwVuiec0Sn3a7nrcmv3np
Day49KPWwERb1KNsPUtQZqd1uHbRki9ogABk4kKO2t96j2tmbC8y56C8aPWn
Vg14jdEXDvrrLUnnk1ssFEpG9SA8rUvpzk6ucGLIISxLSvo4rEPxfFe7vupK
9ASUmSVR6ef/VK4yTk4ffvWTG543kqiZeypKD1x2UV6WPjQfQGXSmFn6KQc9
jFuOztyPRRbLA6DQMU7GVNQLvs1SgGDNMrT77VEDtAWxPShJQErzk7RisjKF
S+dT9dxB5LMcLKyOOyefv7bC2ykEuZVBi6ibH92++MLnXNZn7LHSwFu0piIC
8ORLE9NyVYbbeor6ESNoTqdC0AgZEPaKQpywbd8Af01VLDF/uE32kAb8zHm8
8a278+QejGoytHqKd6YV1CS5SH/JpZRUSkQLFg2Q7sb66qt9nBtCFKtWydyy
MWS5ePvYiVcAW2N6lwiz1DRV46fEgYTC+zuuBuZLZ6XmtD2t31wA/sKFmUsk
iKGkcQyjF2/tRz7dgfD/sK1gbFvKza+RCTgqqaJru5AvBYJn6uDZTrlHCKrr
yGPmw/SEhy1LurN0L65mxJ4YhJUG8np59M/i+0Z8K95a2jbiHIskcUXTEeza
TvxaG81dM2kXVvVrsBubLebKXh5kaLRP7m0DCe86so8fVbFVnhjGGL7dvPVP
GbucRc+SPmcPCXQwenRQqBqeQE46KmxJDnXrHZ70G/FaMA583S89udjkwwvj
IcwZG7dZpBzWMGWolR3uDlCYtqMzml/av5fw2SY/LBf/w16JbmlvAoqSkKsJ
XUSmG24DWzuxjQQWm6DXkxmE/pNngwvoWsa0nF3GlhKcAOlJsZgtMO2rxKwe
G+XEpYEXNdCOQH2AFqXQ0CEzvaH87t1xt0l4k0eqr62WfO7f2Gr1fVffQP12
Rgq0znDqO8BcnqalYdq7hYOD0y4j39ybhe1J4ZbJd7PCZqob62YIPEUA8QDo
rwzFQSahYPRRXMIhTXGAW63jvU1LU2e15FCrkEAom5jxCR/XK9Iq8NS/Q7e2
IndyYPIH9k2PHngX56jowh8ThXW2TZmGnmrYz2pgeZ9xar3Cc7NPubv9ldAA
v91EZaUwQynfG4sRfl/6rWJTb4g3Vm+zuIwxTGz2OLtcNzZ8GaqfM513Mo3y
ApWhNy0/socum2/hUpPjtaikfm9d7yPuAchd4nkUr3sLPrgKqn06CDjs/HDb
LyttAgg7w5GxjSczTu7LW+jsG7KvS/Wb8wHG1Ou5XhnvXdkojCRFyN3Jo3/L
NgbkvIPva3CmWzw4xY2IcTBtxw/P4HfknCfTEhlXceUFJ2ljOmyDz2OAltw7
hlo46W7tPBsiMnPyTbPD2Ktgei5Wwns7ZLdTEcNysTy0mACAWNcZP/dTDRj1
oHXgELU1s1gj+6L+qOK/loM4WpoNY9c1gPgNqQE8M5yxaP+Aa/wJDnCtIvJ9
QORvSUZawt7y+KPRqskB0L65w4IldNq+TmHQvhrsE21HQsFVzdGjN/MrYon2
J65OldPT6GzeoaEdMPJiNMsUOR9BT3AySzk/Wr/kkhiuip9gzdzHUZ5uaE2O
5/XyA8REbFXbds7NAdjE16cd1p3JVWYuZ2D844sjZSRm/CwwWXdf6VgKOZi5
1UxQTsZOWZjBOnzsySFH2XdqU8ubYL8aD0xerA6TDolEs+0xNK/mj8Nv8VFO
xji32/cI21xP2Kgf/J81glEG/E4YtA+tztrzgG9yD9xckQDZmYnXZn9wJHrZ
EVU23Tg1o0M2lf52e+xgj/s/vuN78lriaQTXB32TrcBS2OSyn4C87usZXDrk
ulZWzw5i1vTeD11mhhJkruySx+Kn+i8kwYSZUuV289MLnhtv8L8WG34gTNur
UlflwfL0pvdm+LEwuKlN2L2wu1FncGY6ETzmrE8IRSoL/6VPI+svq0UT/GJO
P9TqstFCsfOhiNi4Q9dDKqAaduBfQBz2x/SeguaZQ5lCkDw3bGWcaUoKNOhf
BrpCtYaPdxSiQPH+PK4OQ9ga1Z/Da9PdOvwBS3k78xLQSwf22HVvvbokkrYB
D3mzYUxMSocpYUfowDO/sr17gHEuNL/JUXO5II4++iXNRFd38lMrJpr+tDnj
XNNx7zQmzrO1ATGrg/9pkhX9q4A8ltZobggItCz1Y9QrZwf89UYgSxBI897F
mSjVI8UxZ2f0PoEOwRn25xDzB+NWhN5lkoA7t9dg1yBigncwYVn8I6/HU7u4
BCiUFR1538K/WL9LRxGDFvVynBnGalwqHOO1odckaVBGOJowL5mdnEKhbbBd
dVQkclE6VW4OemVzkGFy844LnLLeC9RobqBph8IpoIl5bdF09RXvbPchW0kW
KYqn+nljSv/X5gkDbtOZZHf9Z4eE2X2v3xJ8RL2I072c8Uehh+PJykf20jaE
0ifj1TxBbchdRvFV5w3gSGMNwMemBMipgyN7sEjxgpvsHk8B2xYoY/hMyNpt
xBuC70Rkw+RaLUC9YWOpSS8demU4+XhjkYLDYxQr88alMYP4s6KNtPXSpGXK
6LlSJnbAZ7Cx36wlPvs1H/5PcrvYyYmwVFoUOeqzz/OJaKP26DDK90zE3flg
gYjRuaObd5k03lIVThD7LIO45xDN1Ok8SMKmnQV5eMKbrfcr9bjz42EOqLv7
iD2WA9bnPEaIzdZbcRJ2vLBSB5MmGpUZYRgcz9owFLq1f6pZlHm03iNNvKpj
gg2Eu5zbvVKmxWKxwB3+V/YcVoiQfzNvqZiZREWpQYQ0wvPZPfEpu1H8ezsj
TJ1auEU4IT2sTFKrDACgygUrBQl9kr8m6ERod3fyf9AY0hyumsJYcrCo2syC
QzL/ZQjx5t3pTZUwfWbO9cD2RaK2kJnRS+pPjyhUFadmwDbzutC3Y4fEIZXk
kaab0GiiLAg0LN+Ve5DNPqS2CHobAE1NkZvuY/O2BB/CfppRDUaYmiECywY7
RUSVgAIBPi5wmHz2jfgET2U5VSzDp31rqzSkap+MKI5jCG3I7QXd8uLTTcY9
MIraiPWer6Uas9zNbjs2GANV2BJOTq5z4NFLXzQUjmFoZuxxicoTcdoUtXFM
BeA+zlmKFXdvpgczzk94ipP8b0O/3ZMti6kQ3zT4/Z35qHhOe2+T3EmEVzXp
MmCnObU43LDM88c4CaTeAU5vVd3jz//Gklyrt+K65UUayxSVCFqusOCKoez1
EfFTK+oM8Tq1xg14Pw5eMPFB2M86hKA3fQe6FrhedRNaPDOoMdYPzp6wurpl
LM+QGoA2XJ7Svc3TU1UbGLyvPzJpGem3GF6Jnrub96qW13emW9qFgjBJqYmu
+EbEAojvhSqc6VsDt7lPjazIttTsdk2sCYIuyNzvCu9w0JsvjoqBDgOQ8FRU
/x1JvaISeA8l+QmooTls4t8tM/rJoXomRE5HOG1ifoccCUNA8A8xUzVY7TnG
DdsDjSsiwr8gQoAFLcyUAjV98lIqrs1aFE2dsOFOuWhAQbPGCtnJtKgDlE6T
Ar1XAboTXG+IYCN8TGtgh1Bya1eT1LOTnCYvsn9PmttKHCOP3BjCHM33/6ev
wETNWLgf61xCsXE/N/7PutECoy98nmHuhP40mjg7D2puTAKa317ZbIAUBx1+
R8UDg/0xY45shb5CUZcxjIKClYx4xaC4IAX42KIg0/Og6Fnzg9bYavte5kpY
3g5NKF4SWrIbiHSv80jfss1NS7fRLsViM+lqU15BU53nmMqjra4awCjWB42w
tRPP09HsgyY23Si5/8eb4nEJ7JS1X0/mhfkNjO2Bh4mj0rWqOllDDQ88jVt2
QHFYN0yId5I7b594hC9Tcac0YBMsx81wwo7Klj/ryjVVLKor4KOtzo+zAERU
CmeeXDWUzt0cUEqLSq3o0sAfkR6W8T57iXvBRjz648C99EkGVrl1BLgvRfGY
GuGZ2QCt3vBKgXKCxD7wt1K/vPvkEYzIWYcVB5pplpgqMdCIll6UFcDMmuZ1
6b/Ufn3i+M+8QA6B6aLMf/P6OlnGdA8kpJ9dULmoR4rfQjMp4RUmTY1JVPSR
K5jS7DS8wO8vUbOdNmKDNNjHUmDb+UZPXwzQtHncas54M48RW7uD1/Oh3192
Skj5zgRDO2Y/7I4XETUNgxvnQdiJcKigum28OaFdnB8Q8t4yGrkYrV3oriAH
VDKfKWJxoEgWNJzc2hJo3ruB08KVgfqi59LHHahcch0r3NiZQX9B1wj5AUSH
Mg1NnjBmOemm3S4ILm77pEkerECjnEYr6T4FGe2u7nPK3+U/Got7wTAwTH89
7+ETiZyOulNtyKPWjJpnceXcfwV4LI+1snF7KFvPlnhXWPPhn9Y6h7rHzLyM
Gwk2SI8stijyUDaWpDryD5mJ93n5Rq+HnE9288J0lcZwVdIRsmSdaZsFlSzH
JBQJgkSSaO2DQZIHmrm1+2mC2uoicvbswVEz7KhD/bsdI9A7dP0dLp7LvkD/
AQadYDGXu3IQ7xM9tcNUPRMBiDqeRH4o57IBevGG1hpS63wtPi2d/uBAaYTW
fk97xr4uKKJuH8+Ch3kjrrcZ0oAEt2f2g4nquTTQvVdCwxGm5nK8Pk7UUR6s
e6xnOz1n+OfyA2vUQGmZjnNZJ80x+wgqHywWFOl4m2jgjoglifJXduwCm+8o
ovPvoCMQ2zAF5yI/RULvuNTn4JV1ksNE94y9nqjlpXL/IclaXMlLo03dl/vr
YZM6eQ7wokk8rMLRbKWaVMwm58xvFNCk91Xl/jq1o+TDX8dUyFHCnonbxvTI
nfipYSIeDP2UQWZ7t5FR8wIoy6iHNtpKuUInQomnXnvvOk5fsW/NtYbdA03M
Yx/8UgD5V5Zp0jwn7mnQOap2qEPbW006qVrC8ce5TS9DPkpdrc7lMNx7HHra
5jNQPoAG0VLFxIxswfRFN9bve3la3u0usQzWSA4z0IHfqYsQEmByy38GwHyx
1g0pYfOfwlQn5aoLX5T6G10iONAhb85me8CXP2PNkpSZ3OLKP8zoIl8UYiZI
hhC9mp3mDsl6b2rFJ4nNMY80spHhVI7Ej7ol+qTu+Yp445u+O6cEOarbihJN
/pYCU6XQhUWqrlfTZod379X1j7kCkDqC4gv3GbS8678EDXzYUKc0Q72ChP4B
HwCYb1ocm2tmlQ1+oWzPSwtN7PyALLxdFM9r0k2VbA3tOw5hf1p8Wo0230hc
ZUJBvjOzhb01McZ/jAhyPfboSjMPg0RHGye1iaTPvx7lOPd+OvGu+cumOo5E
Gacs5OT++Dy8qIX4Fq3wGDyZxdwmcQomNJIvqn+Bnwb1vzopUCYlwjP1oSRq
rw8GsFuUwziroNfW/w/KeAC0UzRJW+VcCmyxf/JfsEE/JY6eVlVooRJpgoLO
LvASFYdR4bqRu8Mwme0Ik9XdPkXCd5Jse3zVkb1ryHqrQ9zO9ZFJX5nZhHe+
vvQWwSpRfzAl+TLKGr9pdzqbRrbmFN9ps32NUSbRIVOlkDPrWf/9pwkoioXq
WS+tNyhVBqy9SUmjG9J+T7Y2j+BISBtL7T7C8ipOjEdMRFKILblHy289aT0o
NcNHsAgN68Dh7muy+dBUbCjb56Wonc+6CaogXjzsnlF89W4ptvuO7bzFQR8o
ogSTKHFIDhkZT2Yd7CAqo/90A+oFhSJlzYQ5PJn9gpN1cGac5di4WjY1gCOK
qRKW3WUeFIPEtaj9pMrHuzh+68KfE4ZwQL9prngSKn1pCV4B34EWIta2rflV
dhPkebMSoi1yezEeF1QQbNYJpvcKVdY+BxVdKEUWVYHSBihvsy2K6OmLqr4Y
ai4MBZ0q0h16FveD4dTOXJbVMLsggbWwCaiFZ8bT2p7cuvbttA2vy50dVYqW
SQNOlda8QclL3EJG2hx5ngScjp1iB85+rv0dDWwGJZd2dpfWD3UZJeLqAtt9
HyjLuurDMYMHcPjppnjAEcO17Eyzj2aXezyupb6UMuEuzQc+YCInrvS77YWf
RYZSX2VdBXf2gzU+mDFkeMZtmEDcp9uL6Z9rZiRjX7/4zvkWsTveYpG+c4C+
Ghhp4YhPWWKhJe44thep0imjx0gjExWa/7XrKfjQ2CtijDmKEh4zUbR6cHcg
koxnRNAlXEvuwVYcL5lFuxYYFbfBqfsYgTW51h8IA8q6Us+PIeycq199pYb6
F8fF1leC4Kxa5/xXsy7WNgBd9aBrkRH9Xh8omO1hjOdzJ2aVt8/bfYzEI5XV
2G7Lpy3jICf2F3C8kNTxOrevUGFtHGjuAEGlxrjdm+2OyzqcmEyp5YCEK8nw
iPZ9/Wi2vM9hLS/0A4E4DecKcxjWawPqFWWvWWn0H1C3LgaJI0ZJYz4lFtLB
m8I4Gy29w5qGWjzuPe4Suf81DV2m8T5VFBHJkTWnFte7zRgeR6rWKKwqxwrT
EdpvCDxR7aQ/Qz0UPBcbVjemykQmIJLT+d4vu0plsaeDAOD2s78YraXGO6ke
juhGIBpASTjF1vzJhADEPY3WtqZISvcuhI0u0pwD85kEkIOXBhLt/DT265MQ
iywRslZklNZHule1zFvGPZJ0Xt/NyPSi4v0viI9jI0EY6nmcvQ6d6MbxrKS6
aPQis6/QqQnrPzqtKDwg/Pwk2XD8ziXIY1bQwHlNBeGBppn7HtIAOzJOo4jc
njJ/WSIc6+3PsioJRCrDjGPdCccImSQcWsU7Bvrbcodejm3lQig6c/X1FM93
H8h8H+IlP0sdBHycBkTcGbKzf8RLbiZJvyHVyvL5w2iUQobj4GeNMPrtPlTJ
9hzG74fc39i88mWU8rDDOceMwxoQbjFsv0Lk1MgbbUT0GFCYqibdAwOVpBIW
XeEj3Y93LQs4gUHvxUqD9ZoNrzWpvTtyPkgagrI5tn7M6tfpfQdDT1Pt2skQ
QzbF9ws+pPpRBsHPXOPC+yjZWwIvRXCJj+ZIHurMzzm3zepLZ/ph4k6VB3bz
nRA3Y1vs4r87UkCF7SEgMI7Vr/JivUQem8FMubLrkzxaUCYIxLcaxxKowMF1
GMOC+aB77XXZAGJihHtP8CfgZrkpjEYixDcejG+gOB/SP/jmMUY8qCWgvm6B
uyFy29BiO6n/STJ4Fe4khVS4Wz8t3zMdlMBN1jv3w5NXgVSOU14WgulxbD+T
qYi4qfS0dt7TXTeFcgyiC73oTq9PTkM0QonEtVuTdj1ybKXtMf14TNcDpKD2
aaNIuEtqHDlrtpWGfLlPs5g5qmZEn1lkasfIzFChNP0dIJsIqPaMRmfVpJYd
vU/LU+pTXmoOHAjpR6+REBkKCurzapANV75JPA61g8tAzxqc42Iz+fZeXRiL
snWKsaCOIUhLRKtxEn3oEupgb2lsy/X8qRIH42wSX91V30Z/mqNoWQRaBiXH
mm3lQtt1CABr8NAvh1dAsYWiM7Td06Ojk9rerdB9xc1gcCkBhPzthNI86Cgp
G4mFq0MdutpKTqk/cKINyFaa3Xb3aAtd+0OjxUh2wTC/UG5GApZkTHBzqfsm
6yXeLqgu/gobk9CBFtnD+YGHThFGwddMfpSZX1afLmleKJXr9QQSTL1k3/e8
t/HdAfsECx2j4LphSN3FTv34KPcDgKuC10y+Xl0HxQQEbJ9F2lNNqg2iViza
fnstlZ9zgun2xRUuQYQGpVVxa4c2DlKGhSiLfG6KVi3Iz3O+B0+AbpQDf3FL
eimw1wOzqWheagtptezxiimEq1xtIQYqwMZzve2ognM/HCDj2suIpxQgWpBO
OaIrDYH24a/my+J6HgBd6N5sV6Vyyy7Eu3+15buvGTn23IN4FzXK+07QY2Rb
SKAGrLw1//qHY72O8nE1TM8InaiZbD5s+f0Ift4f5ak2DXleLY5oTSIjWaSi
pF1G1MDNifEhYLzOqZj2y6W7wU9cb+U0WnVaeJ6k7QYsRUe4jmy0UVf+av0P
LHMqZDBcamXwpk5WoxoynMHqH/yVazOOmTyLYALjSfuUP4ZAAmhUN9zolpmB
lGwCjwXUNchnPlssintyhIpHqMZ5ua8ktsSJQE2MHi436F119zieYDpmxt/0
1FmJnokjIuyJw6lZvAp+KW5H0Dmhdb3HVF4R9v3TQo+oumGO90lOxt119LqI
Y4cMIp0+u2hatzfemf3s6yHu0zpPZrvYyfjqULS+0wMFt4UwTKe+i8hAVFvh
pu88zwFxW5wB3zPCCPFIO/Szu3FtC5jhQSV6Amg6/CzwShnXrYgyetvjKT95
IPBJA4Y5UYZIGcDMqJnxWrnnI8pCoJynwFmJOxytYWhaCeGK4CyrT/zVT+xN
yMnhAbr8+B8NIrsDLudDhY7+YHVlUjlA9lmPyk0bHrdd4SVGtT68ayJ9lOVW
UUAm4ZZ0LoPFT0t81jlVgziPnrhmvVH+8iUb4Cnnsj9AVPOaBQVY0sz9E/5H
hmj5oWOfYPSfnxEowC4aliLo0O4JyOjVCzJ+aEhmqk09NTIxbC0vnyomIIWH
nCpuUTK7bvMc+XmBLKQ9QMwJJXimNCKheRlEk1qsSXWtnacYuSijV7QMd231
NgobNXC21BQn2ubN2zRrHo9w6cjH+uxv0hqtcNnV5u94IeLQBUhkputmEAUR
NPm+2Fu6UZpj9NY7PP1cY9oznZa1FS5QTFrsQm9Cn9RMnOLFi359hbCjExl2
JhSl/yAUdYF6pJlH2y+546vWyS2GzYUQuMOka61QcVQ2t5YjMx6o8hYGskj9
3oGIkhbPdwBrbVc53tHysv7kZneh46oH80umg43Zh90MxpCMywtfvv+8C6M2
+zdrmkvMBXXBkUZPTjo3yWyJWixqe2v1TFxGSymxbDgJYGa2fKtDA4d0BrM9
fIvGvmvd20w7EPPa4qKYDF3NEPnhisfUATkyK4vUhucdzLkAGNKrbwU5efKe
HpvNm9147inYs8E2dkcXM/Klr90FtXBGA0do/erVM3UcIiWRgAgGTE+JLcgF
e5ockXxsf8Vh+UxtObbr77HPbJZFEAVJ49974RwuTraq8V5RIqQav4OOQ2Rw
vZIwGbcyOx4ENY6qQeZT3Bw1SLt2DeFNhiQkgd7nC8vDC9cCZSWgvv7gWNmq
gOpzkeB8uDMmiEygJq2ta3AuqkUSQZ61rKaqzL34WSYrHiZNoz4UihCONFX2
V129bBm8/GLBj1wrKWFv83ye+mTFlQv3V/pYIO4lk3FX7A4G4W17GeSUc8iT
UhtSQNqC0g550nnPZ2An5l0TNUSZD4tNq2QE0vVfRUvlaTeGNNf4Xjp1/TTN
tDS2qibiqqsiUN5OnhfJ61gh6DQer1smejscki6PR8jRkzwwCANEeEivJVYW
GPDMuTBNqsD+/vOlIMk5pktzRgYLdTulX6/tPvesel1rIg3oaVzfDU4NbH+9
aQa9HFsYdTTltv7QcY5a3uXH9izXe8z2VFdZbgqREz6uXAObHDE0Rx2fnVo2
1H+QdJDdZgx7zBd9CRfWabW4UZcCMOSle4t5mhM3/9Wq9gptgZHKjExYbDe4
5x2Yt+TydDh1qu0v1U8mdOGK9GgzT185kY5MKd/Q87IpGSF/ihpu3u3b/MaJ
Rxu/lRBe73BFfV9ZwAudwc/erxXhlyoPFfVDHu6fH/a6BI6m/p+85TCnPk7Y
Ijh63kjKujkU2onyU7ZmqP52DiMmNLB+85uhH5/G4aB7otsdQI/NujwfZyA4
4Yjj2NLM51k6FjbRCvlgid27pQfWbz7rOWGuY6WjFHxXZ6zR0hW6kzOTLW84
A2cCrexlIjX6afEcf6Jd/qbPTmYPqOyNjX7v1ZdeToY74Z9HU2IZaCa6KkfA
2HNvCT1DAJty1GyGFKjvXMBuufXLAGcbWOZh55cnz52nFeoqSnMPlcj+O6QU
8ukn7LjLK5gQ02nzG2nIGEIrjlwPQwGSaKo5XMh77NTv2YyjhZ1pmzn45VwP
DEL40jE+f20fGI03hXPGSj0jkyMsQehihgBJzFQhlDG2q+bLF3IaR5PzF3zl
StsP4MfDoPka1yOdpchFyOJZKiOZXr8RPp1ecKqbvAZqO5MT+mDp8+i2SNeT
p4uSwiDMR1nCasfJiEKcMaJfhktAL5VK6N5lo/ZpTEf6Id9IuEJWfjV7DVlP
eud8g9baCbJSsE0qX4lLVwUeDgXTgYu95uTY6Mao/jOchBMWmGeUmvyl9Ah0
zLWfGiPdlaKVRRnVdXve+Wc4TGPimuRWo4eh5UC5YovJhTvNexBaaqpMVH2t
XLKh9kbf8Zbfc8s8SMnZrh96nZ72F2ESU1f1aF3htoxzF4K7sFpFwC8krnaH
gNLPemr+In6OItBPuX8Ole+eUwPO7G4F/Z0t3993vPul428aNTZgBdxSuv81
VqXDkvVGMugTlDrbSpP8UhpZq3uSjI9Eg0ufzoxzlL56IwRe717Tm9qbuDAx
0n8H/5wRC9iseTWRFENq9xAAbDMm3bh0xwWO6/BtMPG84VYKKe8wcir4I5Dm
TCCEFqL9xCS1o/hox9Q36NOMevDqpo7Zi1Za0zV0lDnU20eTJ9QtVmgboLnf
LeP0KIqS1u3yXhNjnPTQ/uG48fpCItycWwO1hNQ82urliAWgGv3CEIOMbjUc
emfFs9u1I7uqTHfqqxXDawtZ5sRQPG7+SP1pLQE0zP0hA6+kEqMLgOI6NsUr
teD/O+d4bmGwCF/wbgZwYy2mbrzwrqO9X+8z0mq43tftokYJWV9RWJ5DPp13
F6T4LrXjoEL9R2sItC6AFm45+r1/1WbyqpKir4HIjKvVU0DZajuXTnKPzIIP
CKPdLh/hf6NEyPdqvGWfmStSnqAZLw4lXDUTmDuafCMOyfKBqi9uovTU45j3
GbHIAH+IJ36GQuAomYQI07zXJwtDZ97ikLX5539KObQ44NJky1X9O5rSGI+J
iq4h84sNgS01iTuUd5axYhwxtt1Ej+kyOQXxJ8ucKz1aOWja4ajNxC+0uDwr
Jb+wTkTNtFEPfonpoK93Ahr1tayEoshBj7pqmmc921nkxM8nILIy0rm4ugLy
MD2Lqmuc5LX7wPVgcv/+gf8DRDItQUto0XAWUpvZmBTNgS2J4tuaPesn3kVI
WwwjVM5UUecT0AjF0svMQh8vd5XsTBK92LK6IJi26PgOjhZTZ3bZSSo/ZwPo
S9JIjZgoMhDJ871/7NsE/54RirDD5tvgZCVkjUJrkgoZM/cBWqo0w5q8QQSW
P/Loy/iYAIMEWdo+gGVgUdnh04gu4zx6bHV6uIOttqbd1AR5IL04PiJCkRzE
t+hXSgW6WgG8uKIjO90M6C1DEJqgGW0/+qmlS8SX3hecCracoJgaZaiwW+sE
xyd3a4lXmKM9R11sA505Yj7cjZw1I7Da40/xD5NMJyEldP8vyubylZSeNDQh
3qeEmHzJngNe3CR2tsX/qo9aMBi+3ngIZvqw1LHZvQIlMD90sGd5eRnlq002
NlJnGCBsQNP8eb+ye+7RD/sNBTNmjA/azvh5JTLiworet5Ylwpz4ID6rBmbT
tXCnnVHMTmvefGf1gL6W/ZLfL3lrveLNb7t+8gUZKXj/dw6+ot26NMKo+AfS
+vSGoVWOO5ca52JLkmDWavZkQuw75dDc8q8fGb5AlRlQCSRMBggFWxTfH5N7
AtGBo/bMj/eLQC02CSV6/OsTuffjfB7t6kW55K4uP/vNHSwvMYXLD1gYSYV8
HxPmAA0ZvY2he6wvjU7M3mAN1WDqWdavau4n3h2H7t+yLoaeuIQIkzSALBI2
+eqPN2GUsJNS1WP+ORYod9UPRT4zcC79+J2MIDQ5N9AuekiJfnCjK9CXSM/Y
8Ug8YlRNvhi/zZ3cCp3dgPera4x1QFw/R8wBaeUxKUqRzlvu0QXtr24km7JL
JTREFRUA1+eC/5z3camo7auLoWZNyQUDdvTj++g1aytadStBKkAeJd5RzKcW
jyYCUFACMztiO62blw5PqiEjUTkXXv8EfDsKKSGZaQcyJRs//JwyMabzxQzP
SjxwtWKh3WpMbr8OzX5iaUKbfDosxLNswbsWURNhp63GrPa8QmxK2huQXNut
dlkqPg4PwHPjRlrztsspN4Vpb984KhsA1Q6FKVTSKrC8HIR57IdV/6m4ErNG
P9ucjKId2gbbRQM89Mvx4wgGsR3do/amUXLPSkGrNI0cVh3Dm1ZkOt73AJ3G
lclU5LLmZsYzJQdzySp7RL7lYOWCP2MHmRI9wfjeI0oxXjRSPJ8sEy0uLPd0
GWjVO+vPhJsdYSS/mnpVrhdeLcCekhiSKgFggRUGqDh4xrsisuS+BUg8mOjD
9OOr6pi+tzGu7o2cGfzGAY80Cyym3Up5SJPc7e+0bGQBLizYq9OIko9e+PhB
M2y6eJU5DybXXs3rxVfasVi11xBYYD+imiSICAhT7tKt8Rk1Utb8izUaE9Rj
FEiFbu0mWb+mFEvJmxzFWI2F5HOBmolzZ3+KDilbuQUPKRJuOPIXk5FryPCT
m21KRIC/m0P2uZ1exaQW+eZQ1HjZVsMsZtkWhSDh4LILaFZzKcRAlGqdRs8v
2JGkRwhGL6PmysZIJBTngMhPvCO5yD3WRD+ud+adMdyWOGeLkmtF4yLT95C7
UCXoaYFMFK6kD/K6hFWMTn58iy5Wc5lZN3ouiijK5hm6m/ole2RW6z/mG3wj
+Cn4zsWLJ1aXTWety7XfYCHA8PF+qYsgOttp+9kiGie4OP13mjq3O3PRv9C3
L5qPIqkaTzvXWKXc+A/wNFg3SqyeYk6SXjoxz7JN6xG0KUFNHSZOz8RtRbr0
RplwFtlDE3OMRRUaqOEV1ae+V1uWaS/llY3ukfk1cMAdxPM7cAvpjubavesq
HJ5wbh3puLAQu9WDBNFRBLuzCY82QJryKp/KSE01qYzxL246p8FC6pcvdA/c
1M5s77sGvgA880kYuJjfYImkr/Owx9E8S+ukZPyrw32afZC1uD0aoA7aDTm0
5vxc8hwie5qGEFxTU5/eJLc2er3GGT2SeAXY0XhYadDKu2SJNEUXKJjIBFWM
/YMT/cmaPUJbG/9XfWMnfJD5uS/tenrihWjX+dxxvz/Y2uPUSplFzDJVpONL
+sDYI85n0iRn27GLDnDwryhDeScuIoTxOnpxm82z8zS0GXcB8l7TZSIWf6SY
yL09YWLRpu5RwPT+XoKiPPb8zSdv++KLOp8pS3kbEdPEYTmKMDWtWaWmjhQn
LZlKS15/uN2QFTiNQy+aDF2KUywJpQDfXXKf7dq7LqxkJ8cC1NlLNZY+fwrA
A1qzU3pC057Ca/yR8ZoTBkDEUqui5nz4nNra/p0tbXp7oE/28mmv+Znxv485
34BKNkV277T5gxUuH4U/aEcVIyKyJ6zFpCGsJGf86mEe06+kvF9p4fatLlOF
yTIYiY9Uca5U8AWcXtZt4lFIqJs3xsZrrPMYP1M0M9lzfWO+Bbjz22+AogRq
VTsvj4doNubD/cu3ZE7XnSsPE9mLbkz65UTMLIBD2IDvwZYbUcQl/6Uk6P/a
HfA2FSQMDJC7dwN3JzBJIZQ9AMouCBiByyPOKvriC0VEW7PfguUCXjet/12t
sjZonRzEFq11VAWrRHCJ+TXj/7cwwx147xLaXq0nkuNpCKK1hjo7Ou6XUXIU
lIfPrU6mxgQ8ho8G6mQybvWjAlGfXIyEKb8P9Iy/V2MWuP7VJ4jObDRuVYDD
5rurvoQNSHdBQYCfUcowrvH6GFhmEAwLoY7hceDpah1CuBGy2bGz8hkReRg3
4oy5G3WKNan0D/nH6jcwswWSGt6Hxo5j1G5/NaEOBr5IKEnX/YNymIEaG9Di
xkaYAUt6VTSvvFmXenlxpS5D7pNYDxUZuuHUksN9S8aid0iKU1vH0IrvuVMK
Yc6nkq0pmYN/dKq/evqof7P8QpYNx3rH9B+DwD3Hruof+NXz6TtfPwgQ+lkU
RZo/p/DbglDvqlsTIaMEj8wGCzY4Dwv0RpKuu1WrLwgUuzc4wOeBAkXhbJA9
YC183XFvz1ymMxD2kYUZEWwNhj0CiifLmF1bnsn69AnDd8wq5p1T68pfT8Kx
logMfeLDtczKQd1rllZiFvGq9LRLvZ0AMGv/RC1uZ+WeAl7zMWMI/b/6UT6I
R8vmKqhLXlslX9eAy1dQtbUjvGH7AACFNTaMOYH3D9+CNYOk07JlA0+9L8C+
fV/aYDvXPUoI6DQOQ5CvfH5nVnJdACe/7mxzaXgkWh0YYEOpr1l4XhIPZUZ6
Q2IizJHLW/iTsKpmB0zLmzjR3HcD4O5X6qphVyEVyDLO6oVLg2587f289vMV
7cAs6t2KUpacxMVu1v+BYXhwvKuPcvzFRzouu2P0esv5A7xro8ZvEDcXhv+T
JjNg4zb369h5+FLQ1APs+CWJvkjWZWjrEIO/JSxvvi5Cimj5TNlww8mwMZYU
MU7oV2oUxohi0J3kwxSqyaHvaQQlZ46hZxmfUpNOTPvv4B6Igm8JC4Yob1mD
G2yq2rAyJ0s7rjY0Nd4RXwxchAfqbakUpF6/lg3D1mqI8zSejNQVfVr2e6f/
C+Tme3IcNjmCehhe/9Gnep1b8mfa3r15FeLcziblg/80mY3fHMs4qvzbvuuW
ByK+GfPSePffQUAE8bRHcL8JNacSd81yL9NhUn/LKt0dIUq7JThV/v7loE4/
bv8p4pq43FQuwPbNe2rLCHEOMW+aUGDsWAfnvxkJiOV0c3jOyWfKMzp7ePF6
IkOdYA/JVg/RwMSKkZQHLxwsM73tIK0giNFZH7xFPHn7p4fBxzRGL+R/L6++
sf2jkH2EuU0MCxBicmkzAeftQeecLjommEh5sIInVrIlnpR2r6b5ruuF4fzF
P0jOsnC0Ta3mm8YbqgYW5kg9rYaIy6Dv3GKf2fDLdqUqEOFXXyBvPHkLdt7q
2kxHLBgt2RVdpt3gaJ0IzMRP3JpvPfPWZySBV1WKbLP4MyaXpBmsrn/wpaxS
eACdDI5Sn23+Gi0ydWiOHab3T9PWlHJeDNKluJ59O103jwCziDpxdtf20sbL
YPTEkKhvJDBDk7M+Y+KUeYKjikFhIDzG4/0A29W/PTbjTy6epJYvE3RpQda0
1R2jxMZodFRx3drikziGz6mQzHQ0p20nj9xcsgpLO7X1TUvTwKSf29muSJ5E
LdzkwDl7Ch8NiWuKx0QPRQTZkoub2U3JcT28J+96cE3BzRziRzYlEAkn+Kkd
vxTKb7Eh6ZvT5Kx4x08fSdH3Abpto/7sX2EaaNYA2EjBxokEKbHNRmV5P2Ql
2hCmmLF+DDjnYcT5FGXY2CB0aiip5Y0ZrB1ohBwmAxp/H1vNYAjTIark+BLF
peYy/jvmTtFnnHA1qZs3L4P1kXxtFqSp3XW+RuGdOtCWiqXRAmJF0o4rlf7T
LeMWDSzV5DqWiGglWiw298KsHLSd3CvWxO1K4SADO4Qa5YiTz7WQXzbpDEXq
qKsSj8P39Tx+QKgg8Kp3sUcb3RYtimqCucWff9g0AMAcLpEd4wfoRWpRfqFw
lVEesp+al/mjxvPmucYMALR7nABsAj2ylGq+C+RTptOkg1iJ0aXLODgxWhOc
sJGk3tSOuhYRkiQzepEFMD8zddloWl48GFhKDivtJLS5/2RUROY//MwQxQsb
oBv3Jj61sk2SA57PQXNSLIazmOGA5T7Z+exStZnW6ZsRttIHviXYdCppympD
ftC0FINjzWSG80zlaeDCgN4WRFmIZGgunuw2ArW6D2at2AnpRBUa3ihDqFwE
8n61Ur/qu3Gng7AxBDEdP528pZvThYUyumVULQHMSIZB7RzyubIMso/3LmsO
Slpg1q3t6wv2Lssa2VEc+B0qYMlouZ81KyJXSRP7A9jTVU7Mwe5Oi7azVCv5
YlMfyZc4DHhqRxwMfWXUOrG//MY+yKi0hj3bnxYVxXgnhM8acn4Wm6Syv+Kq
mgXnJ+WD+hw/MstijMUMvikMJScHzJFe1POPFaX/m+S6ZRDdoEa8hakK2ub/
S20gT6Uy/OKGy1OuWDa0wsh81sDzP63I/H4aPJBRP0OSjBAo5VfaRl/TrVB6
0EhkF0/3uF0ROS02TxSPIxloBg2f0IqllxU1pic/Hff055jYpNxJJv8JpcEq
6+GxH2jWJZZ0HZJoFuhC4sK2bSMPiC/QGLoUJnw8BvMQmVAyiz0rrVEINwcK
PTwMFqftleSYxggoCURThtnAcSjJKCMH6dAXnmNVAG8TSfXP9fLhgt5TtaFX
dAeUug/6bZ+YOaO9orglQTBMHWpkc71/z5aolCo09LP4zYYPGQVWf0Ew5Ml7
dPNgC62Ow5BcFoLZ3okLWcO8X3xRobyZ+Kfwvi7Y8BiccDiDFB4gahxwFnnl
8Y3VyazfQuOJRXL+84d7qlaD9ATe2vUWYx6kJyJ8Gdl0Oths+1K5PpujkXxN
lj9nwTVmMhDmzXwCDhINfkkuUykRutNpdonP2IvLBw7SKq+X2CE3Zww/nLJo
GQRaCE2mFjzVupIWKug0ofYJT2GBDvwnYlwoGyCNL0OnI7XNJJmHzIaG193n
OkK3dbgbjwPMM7+czHtbXNtDU5R+fK9dewPmRgXriYBdqDxYI1+g0poOCsvk
tq6uJPvlK6veDSz3NpUfsklEht1Epv+HQhzQehIQUaVghEwKZxevJEM2aIC9
LzPoa3cMFaK06XLLfkUl7xe2x07LqyaE7LCpD1I0umkoiQDeiLKp5ZbZICye
EDLkDEJsd/JAfoY6Wx4d8q53WgILOv3FCkoIKg3A+nmoAVK2mPHx9tVKnRFf
IJtA+/J0OpoGp3l6UBEjQtHGh2mqBl84++L6zGs8YxMGMzVZlTfoI4GZk0FU
Ps6aK2ZTFsOYkbgZLBYGZGefq2N4lz6KqigVld+qxe95AYvX4kt4c6QxawYA
OG9t+yM+x6BpDoaP8WJmX6GInMuF0yXRoHJ5tGoslcjPcgvmPQ9+h5/vVBxr
ZlqFdBVna9ucOVBZwfOBJqIxokjAdcvnpI5NrK7xbjUkVSYwrZYd2ugEV3rn
1Wrb/rgAp3XNyb9gRuEA/C4szES8m98KccUTeQd5VNFqC2wUByTyaRQ0ZIeg
0NwCQEbCHw+F17SM3wOcDDzWljfUaVNHrDlUNa/lsp9EURCJQua37BEGeKxs
g1epfzJl3qj9jflGxQpgsundi2T9i0iEsAnj0SbUksbQqCvcwf3wrXw5UDmP
pZ12hy9p66ZqB5egwAxl8FxX+EjjkE7xozbCt/t2rZBHcDVrPYQgbDcTeZ2j
3whtFQb9C4nkSzZuZwbo7lJfusvdRujLFvEEzxgJ3jQlnZ7k/D0dtex8RN+e
xReuwu+ENBGhHKrah4+uzjPoES6tGqVcmWeGn6KHPo5oztQNk21+qnzyi+vh
AInnRQqcL6g236TD243rvDJOHcYx5bhJ76N7cgdCGQVaWEwJGlKBpoHAnXD+
Vz3OLouE4Ix7R3HtMHo8FOc91ERWm00men4xGdw3kzuyl1gPWjb2PT9KVAMH
8JkvFqjkk8xbZ4mYjq3EuNyD+5NxMmvW3LTCP9F94Kkk0x3G9KDeGCEN613p
jx/znm8DQuLzzn9+f/ZctDJQVVqGE96zQEYU2efuJNX5NSeLzjEMroSQ52UV
w2yRljDjOC5KCj/HDvPTDjfUo9LNA4GmQXbAJEeqJ0Pi78ozFTFVuOuUuzX5
sJGrp7NZdDwdqRVZ2T8qa2mkF3A2jSXZo2kLDBlmKD97NktEKQbkDdRRztWc
JqTENn0CfBep4cxnFh+96x8xqK/XSwQZeuZtxaXZYLDa1+qMNq5qAsXcV53p
r2azXl5axgcQoolu1aRfmQZtQIGIzvvZygbZrkumZa3jHThLfF9tG4AKroYZ
Bb3QOYO/1de3p3IXqurk+fHPdeVmJpL5HJ9VnZa3aAVL5lY0Ev39as4eI5nP
k/R9UykoVGqSDJ+r0sW20FoUOtge+4BTzviGv1KILUyy6pT9qAnQEdhHPvVE
44tVlll6dGNrqn0iZrv2e7desUEiD/H9KUgFm77J/PaUVpOAj+8ayg4gsHY+
rPM4FPfYaCyojTupRtbZlAzhPUBUTwOPegMmvxyOSM4hUeth76wXMOKc3Orp
HfobDwtMfyXmceHCsly3mgsO3U6COAO5ceMYIlVgSbOgs+xyFol0sWobv0rL
zaEQZQUzJk1QmVlrhGzK2uv6eJslBHPFxM8g0mzKKdPK+ksTO/LU3xcZ/O9E
4mxXdstRbKq1aEgKeU59xXZ+uCMZEnHbrKAGsbHlRI8TfmKVEat18vwoo7/R
89BhQVmy6HI8ca2qkhKXHcDxO6Aw/TRl4+Tu8+NzLtjKGawDc/sHuBjFKKDK
H0DcZoZJGgIS/PVwsOYuytvvato5w+oAB1QFMYp+gpIB4SaH74hVzWx0qXlq
6bp3xsB982HGZo//4pFqKX//L+a3kEaw5tfm/l0M+iRpmWAwhMCnj0/WBcWo
fRrFXNiSz+OdgE9c2D1OX6iPZBeS0JAQEQKxHUrfhtxsjpr5H04Q+Zdagu/m
i+/2aLcPf+BlhHIx/hp1l+Zkb1xkZNN2+KLvhgzQC4jGGnQfOijOn9mblJuK
TcaC/yo5NMgMAxfIwV8tmbYBeiZy3YwDDfjRx7fE6FJk1fm1jtC37+qtpLHT
POH3dud+Pr5+8+6eE/cD5FcAzX4sRCynELPvOZisrUmRLdewDg2B8UFWlyGu
62f/4/4o1OlXMPAWkAWMMbDoyiihU62gj3FULpRoqG4sxyUsMPStlpxchX9F
ohnjUsgF149Pws6k4+059hBav0WOIXGSbX5Ea9+Mw0JUM9HOeYNZsmWoOp+B
bkxynAoTxeWlQOFKBoTDtrRUr6YNCZmtKQxKsPwHpDDamw/1/rhR/mweqBkY
ywS0jACAIVW1t/E0VWOyEhSQDjWAR99Bus9EkTbeOQ8rinB4jxIA7ZMNn+gx
DKU/3UsE9nvyeNXm40s3xl+Po9fmoOAVGoDiFV+OTCzPoAexkjbcCxb/0/mY
ESCf9+kyXuS6MAWeOSyQexfJecOls6A3C1G+2Fnd471H/goRFSttJGePffU4
3qIynXGepYmFr15mQ91B6GXPGhPn8kO2LtdR/T9jfxovdFBmxfiAhw+1hyJX
DSeFZNJaOkqkGyY++foXNvHBDctDrbCQw1auizy7WJuuXzhTH88Vr+z4zOqs
BuFvtnxqYe/2vBcvGz3nZNdFQFevmh2QuyouVc2wT9fPGUJ1nK4877DmCrjd
SGzfPyQJE6r7LAzuPIelYLyOJjCEZWtUA8YTsQcxV/OtKsHFcjXTZvsnTA+I
0KIkVl0sDivIeC1NpUWpKweDqaVIpUOsEBz8fGjiRTsInd+4xWy5bc+Ux3xg
JpPaTbJb2ZEzOFFPOXY8BMvmUhLX9HrSbMDFn0b4LLjR4xwCeJxthikRQ0yd
/vChRtNIs2wuDXFgUEicyveQpaMVs3Awbnp946vxfAJY4i1fw4RnVAclY7j8
1/wzqYhuQjwNXaHzia3MD7gMFhOgsbAQw6UcRtLJgG9fOMq4RJH4mhC04q3Y
9+29Wpv2jUES/X7aGNJioiLg37p0i9lTXXIzkcBAfmUdxz5mueGt88TwKXTh
IXx8feZSMyAopoFtBG1Yv31gkGNeoD+WgSo9t9mYDNx+WYexjGDePqhGVgsi
6IGkPw5Kb9C8FeMF0t4xIqdTKWFXv0wDU+r30BZwZIlisHJiuydqC/xxqVjm
yJYab8PyAPlqElkrwvCx8B9LiZfbvGr2PyhrB2aqVuV8t+up9UOxLI5X0CpC
nF6tCmTZRWUimx9CmYnv/2vH3OeWgesX5RiPXC11EpJXc5doPBdPj7Hjz5Vl
soAl0q0ibxzhlpLyk639ZjAs732fWM8HQTLeFRe/Zmm0Dpl1jAHcxzHLf39W
r1NnfNJkyi/W7S0qRRgefSOjnsEj7EXjkkI8797Vjnmf2LWi8gFwcnPNLigI
qmQN1kqmjsFOaSSDdlT8WhnubK3WISiNwTicx4Qgp7BRcVGju3i1CZy69O3V
XIbbbgAtOmKB+Lv5/OOFHjcdQCvQJyAvR37QOMCKK5c5/Z8f5YIVAYj+L+6I
H6OFJSAGWOASLKjoLVPpQLxY+SEUDQoqzlY4mPeREGHJ59Vdln0A/b26LXmI
w48LwxvMnfuIQUce8r5eClU5cT+RW6YXU48SeiR3esAwUy5UAuy8ok8BAeDI
O37xk7GFptKPcP66aGLRcMmX4IYPwO+aDtIwiEUaD7Rn7yli5RaOJzOEw2tv
mCviQ9YptXQTNPBGNB15hs1RurT6sHG7DfH6lO0W5bNDOGXOftZqwesaGEQv
JwCbqySqqoe1WG7W9YHY++XqJo8jG0xDB9jIVi1/R2ZDFcPZYUzsxyA94HyM
USO5M5rXiSp6X4pWQD0yuEZWLjPXKYXapoqEH+79CS+JaFWbfk4QHm2Rgm3L
zYsRW50WSRhl3UQTtOqtdctbavMFsU6vnkUf205X0ErlG3zWC5lXJjHJBbB4
P0jwz0/v0OnFOEL9gZwGdpPllUhsRLXYzJa/qNWoAjdAXCVOeyAB5MFm+V9p
IIBot2mWfBNPbWqhNAbdZ+YyMxKFhTkJijhDsF9gjx6mQl2vMoyijWsB6A5p
k8pGVhhP2cmqkETtxsOmOgQtmY3rUWaNpBV9nAnuvLDWuUWU9lFzfkQapN+L
3Q41jR9Mq6FAGShP3ayXmWlIJkTZpdAYMz2PYpVooBbFWgQpiGy64eodf6vc
NRi1UYMo5A0L5n8ctB7zqsQHW6BUEhFFSJbSd8SN+7XY6GMcAeHjU0ZlvPUE
6obwogxqOztFiACD258sWnym9qr99w/EA4UEspBOYZS1/t6bJzr4MYbbZ2H2
ih7nfqca/+hMQkoYGzhejCIhGX3kj2WN6QQaMH7tnhZQolE6MMBdW2ziZbsm
6LCNpMbhw6lmuFtheQl9+MMAA7LmK+IerJIwe66IqOBWEAXfFZcvDCW0IG/P
If/KVFuDmf96UnwvUvtqqGnr6FtEuhctaqc/XHakSbmkk+YekzXpCx2qugCH
IiLn9zpwc+vxVZ+VVtHjeg1S1AkWdHKeTYglkl/IOnBRhe9Pj61P3eze0Dpz
T7LegARhsdjM9CT/iHaNMQYepqDrn3jL0uGQUrKLS40VP4CoAltYYWnr7JWz
bC+NCgJeeIeUzTp36e5DeHbNy3IgIK0YkRSxpGHlevyxWciLtozfi4Xu9s2+
kdQFKi4ctibCjHwCil6lL0DkN25WG4iHIzIr54Lxikh4lGv7w9KcQj5ISbKd
SbSt/AVU4Oiu7K+ODkMzek+EeUsYcWu1QjGrP2GexHUiMA6DhEZ3f7uBm3xO
qvFr6blzc+3gs8ys2oRLwhLdGkrUtZbtdplJ6Gg1muMc6lurWsCHNJUhbsZ9
a2wTmt7AO13ZY+NwV2wLUa768L9Re1tui6LqK4lsODxTxGwl9tVohh0MjNUt
/zTKNrDRBX8gElTAFwRIXwv0C3I2ANXc+nCg4ocJ1cFN5G6noRMR2JWbX9ri
R3OOJ8qfkIPxJ2SKC90Ix6XMrWal1+/7jIg5jty2eqM2IrVVQbOgf8CwaMqQ
upp4e/Zw9BcNk7UGJFPt2Dv5KjR+3oxKk8ibe66nMKjbeuvUZ+x5gMO5UIf4
NWW8g23Mne3VFM/RAPWoFgjbe+2SwDTkL3qn9ZXVF3xMVL/7s3AfAdAC0mpb
Sw0V4JQ/2LAh95C+k9LTB8XVDG6DgWuLPbRcwM8FWcYDYtzCP9eXm7jEcvOs
UpXRVbp9LRmcaFLk8vNwOdFGmeqk2LDC8NvexXa6pBkSeIXFG5J+jjQXNp0i
5yjRPxN1vl9nnqLwb9ebW2lWh8DFizwXdNx6DTw4aXX+jbgXLp02/ek4g72W
t01Lcqdrx+LF/ZMuHWuI4uQS6bjMpVKnsUBd7frLmqJyhHG2Yjd0OaaazNw9
3Rn4PAE/iUiGPP1YYCA3gPAVBReguVw85Ejj72BN5SucPJAogTn6LVCSRrj2
UF7KDw37b9AerXIDlqq04bwDL2w5pS1Jj9howrz1WjfxecxTjabNPuA9LR1Y
3TqCSMP2qQzuAIHMNeSM9QvYsIt4/BQBBgq7zRl2PeO8IXXnG/FdfvPZNT1i
9YIGY5FX6uFQw7oUAlZZ3jGc4+xev98yrtLEsqaHwP1VEqJexCSzk3uf+fPQ
1U0tR3Sn3Nyzj1+aYy6X8Dw6XLicudEuEpuUMEkFz2i5SA9jOh+srvRkLsn1
T9VZ9/+689DUWST39lyw0DeX3hOnItMk05K62tApdD0z4+PT1VjJ+h5nK+DO
UyDEYQpytZvjOA94LtAQ3+Nn94EHENsD3jSpfvqfGhvnhf0AMpnBEhz6yq4f
VrQeoRvKVdYsJXog7qgPXZHSZfatA6iNRv0hT7t9mpc0hI/7cQ/T4tgrsnK+
+d7ZdwvNRkPsBQdrcOcLjvLorZBBbZsmgtvLlIzgRALvAFhzArCxnmn+vTeC
YX6D7oAWLv2CWrZ7WyjTIcdv3097Pn51iZCcZX2v1ciUBqx6ZMmZhhrskJ/3
wtpC1+Zq0rR/3JHxAQOmR7iCAW1wYpXTuf5rrKd2IJXRO2B1gRXkhDwR/1xB
sc4Ysz0/MymXn0lrpYfVwhQcb/r/ULkdVrY3WixQVSb2lvlNDclqerGiczZa
6hzW9aqlQ5QBYYMeHOhQB5ybDEV8uMRLfjG8v6Z5rdfufXYulh/EieeKbrTh
yloNj8BpNBels1hWarUcXLcysvN8FlEkKyqhUdaobV0SCCSdETyoou6+Eqyh
kWy5CAdc0ch2TFb5W9Fk07n5/HdL8+W1Yy8o7B9DC//64JZMuj9iwEpKSi/h
fano0VranB8GlIUxnTROdNMHXUux5fJKLmKzNosuOcy1v+Vn8ClVSml/soup
+q7zS+O2uC0S/AZVvVRBxxcwRXcfTyHW9GLYXWXQIi2QsstnU3yd0yRSXMVg
ZXLO4CCQel6PmAgVgsjKKiJTuufwU8Yd9CQ3GVir2/yy21jcMVzBjkjYfxNv
XmPwlTItW8xqwF+MMViCu+F7OAPzbwfYgeft1cfh+H56RNqdx1NsJ12qWn1f
JmpSqSOI+bGzNA7LUZiUsc7SNDDjeq0hINi+32G3VpAeCmMiOJvjRWNrijLF
Gmw1hrwFlqj37TDs9Vs8S+gvpsDPPklgwdedZzF0e4uunyHOAxSMpSysmZGY
llR5e/ppHR58ia54JDkDPk4MM415m7WmMi6pHS4t1S+16wIjt54Q29wwS5VL
/d1VpDRwPHqeRTTc2Mnel4lOPDWScWr/W2Cu2ofo6gp00YV8YEhhsa5452/I
aq+0RFCXiX3T5610YT0FP27+H/3AbvKxK83kSDMAYdmZnus+h+xbcyZKC9YJ
doWZhPf2L02/cgQrrlLiZTQszZI+lT2U54fkl8nfDwKOx0moL3ihm3JyyY5D
/gF6oQjEOiI/N+MOjaFJIuWchzxJNEY/yzw3tJyrFiUvBMnHT3kEWoairly0
f/gGlhQa41cu9AcywcNVs592FxYAfQEJ7zk6Sv8OmBoOURzCASncujieF/S+
mwxsnhrB4ak1+ZPceLBSHbgaRgHTE2cWUn5LKS2YqZPn4qcWZJUsk8y//8+5
GjUSMBSl25XIMxXdYvGzTHn6wWBg9vpfHhu/1XEDSfCmQsxVOGkGIdcWBRh4
hYKnucrAXtPkIKFJlBIKsTh6cwNI7UO5ZrTbcJYclHQkZOlxJfvoHRz1EHcD
W6mNIgnTgWHPZfqj0ic8F45F1RTN5f6GWBLGIQZQQ2hpWDe1wwkaB+j6b8ba
L0IzJ+21xyzQe773vLBU/RWtlhDAkRMBREHKIEO9EBEcEMFN65SKk73+YrIY
mdauqlOF4J0Cpj0iWfAbprQD1vHzDSyHppheUucvK5y5XLm24+fz6OM1DIH4
BB1dZ6l23ANReAvnzlTU+7pGWTOzso+h2+UIkKrF1AFs8LxePbf1c1xtSNaH
amr0NHr+csk3IdV+NvzbmD3r4jKJgM+wMp5MunCf1+vHc7n32hiEnpMWWTg2
9ERyJ7kjFKaut0ZgIy6IHs4F6TEdvc6luhkHvt2Mcn6hyFSV5FqN54Xopxgb
v+WxjGBLkieiS1NOeClO4jQ8dW2GxspPhn4W/B/1n3MOv5i+oYkWE01UdQHh
ShGxZhHQjLEOnD/rmKKpxuEspqFInFHE8V+9GQDD4KVvA6JW6Dt0O6mnXnCy
3CYOq5hBHVc7QW6yOQRN+I15fET6MD0gkIQcGdLaeQ7XGh5sGIHo7438UO5p
P6lKAry23+McNL8/pjaHq8+Ry8JAb8ey4qVB1TomIMjmxQpc0WAeLYniF8sg
rtPXZYu5cWGT/0St+g+EH3f0DAxzhmhUz6XF1Kj3v3eRIitYzA2JluVWhMlS
tZ0XZVhsSyCpSIQQCkhx591n/yMYZ10obVj9JV5QHQdlKhX3K1Ygybn2RCon
wnPtvdBtzJqdghUL8TOat7gzm24GRZj4nYQejLVxQzPiulcPXAqdKVkcCyv4
opOLLCJ0hytT/eO9esObc3G2mST5fPZqdFdir8F7RaG1aUTF0yuW2nTNHRSv
vbcWGRuzdMZ33YYHedAsTyMCJXnFxis6bNaQHhPVeIJXK204bZeS6FgrDwda
DFzefrxxvUwILJ+qfx2jt9QzkMfIPKq0cpK1jCbsOlaeVlBAfRAEWaouIh5H
FLau65vbspo/myD0VvNJKi1k7cWWqYSej7f7QCD4LkmmaYJdDGCuw5ADrmgh
R3HtRd4cWNLi6gCcbDrju7eeKhi4rzZ5vNBOr3t79uSro9e3/IhunPQ2Wd1H
CahZG/mwJUF2WvgN8rsGxyUKiWTzcivRyUcs86Um4AK6tv+O4i2L5T33lKW4
mJuSx0nQ10LbIer0Y+7EChOQktnJVXsq/wJcm3WtlCw6M7AwbxUtCO6CZZA/
/xyPM/INfGwS1umYCMyrvR1A+8fj7p/pd7mNllMaxt3T+FKRmwaO5m6gElYX
9EidDk0GS94NE0qaL6bi+bJlWn6y69ZU9tuJCY54YYr5jzeHER03c36VqU97
ILZDVmkezHnWZTSlbRzCyyTohoDPgpWpLhuzEo4jzMayAJNgzqXJuOU/9tz/
2baWclL/joxqPbFOwr7ygkyuJmmsMowMHmBAYDleSY+lLplNq7F13xJBH/M8
bi/EHMLm7iww9xPxOcdHSqHQfOSrBDuJ4zX5N/vJ4lJ3bvx3UiMc6wxLL5uS
DW2vf6W9AumMMoA6fmlp0zyyIQE3LEv2MwZ3VY4jHg8+kQWZ+PMhfceqYc8s
Cv8+XKDbKvOeqe1754p2N2on9KV4n1T2g9ts2R8ydYWfv+1l6Bt/AlQ8pFCN
F0cQXgaYlrM35fjAj2Q3H6UkdGy6dCbEDq00e4cMQ/zIKM1+1k7bXSzMDDlq
yseAacMIk0Z6XUyk/IzArJ3XsVi9PrMMj7kbtj5g9gOJxU4oR8XMkGvZzx9Z
Cxnt0ui2UjvYpoLqBj7hDVOQAVl2D7Vl719/0sqTiBo2YkQ/3aLFoCn8y4lT
AvsHuagS3I8b+jl0i80+Arc+4oHsOtHn3+Wwm/lO3Qfshnt/U6XidRqnDTIM
ZjUGDTp/CBVVxJALQ48171HEvtousqBVO+9t4W/a9E8z82YgjoZGk5+lbL2s
WU/NDTdrQdBDptegH2Plx1bT20fpuB4C1djezNoB1dIHWusryVC0eTf2vn6u
4OMPhLPB4+NYGYRtmz4b3Iyuneuqa6ovLtiaKYRYJOgNZ+tdpaqgAakC0yWT
gBhYHvZ26e3w9JVQE91RR/xQYKsiLSk0yw5DQFiNevChBPn7VwRl4AWuJFpV
fc3D36ElFqKF79AjeU+K2mNUhB6xTY/LpqSYshxvOKDlASC7TbTYwaag7tX2
OWcyyujri33hjlB99z+SKs2lMX0GenzTdHAaCMLw3gg9nMqroAMKOS+LQvDk
B0dNo6OW/diUcw+gN2xm+rzA4JwA/u6iaBj2L5a6XM4whB/cTF9T4oLzyeFN
LCvHoXQzDEklC6tHJuoHYulZ+zNkuBpZfqA8niRQCezODl/tYIJeO+gbtm4o
/M0pH4Cq6rO3Ne0pF/tilWV/vL9vYQO7cvkNe8tkNYtPyPvByjuEoWrOWahh
Ra4U+TDzmYcP0mG7y0BfIYZIZaYwwpJHp/JjPJnW7B173IGNFnZ5ixix5Ah+
eS8dFNw5eu9E8GB20orFfY1Oa/eZc6d4Ah9ggsMFwdNy++9ywQUnsx5damHF
TCjfS2hyoNeNrzwiZbm3lGJsmA1rqP2MYX6o9harHxIEyD/1i66tZaIMs3XY
lZdrAWID9PRJs8NHJCuKekRehxKMqozFT67U5kLXkwDUDcZHGhGjvI3CVd0o
VCIcgcr8MAxYbF72XyeKEW/Vflrsh57qXo4dbUCZmT19sM37mxpyqsL2KWOe
l/0EGQuNB3snnNEv5wT6BFX5R22hqNZi4L2jlMSBRJn+gYxsc5PS0lB6f2Uj
lDmmEjw41Dku6hKi7UPraA1LVXQghuu6IGj3koj6R77Ha/IDsQBuoSgEvkVS
iJ9wTwzf1fawz7Rbtvdp23WhfdcEHhnJqSLsH7WM/6gsyrm1eH7XxJDcDx5Z
wgoyE5caVyI5EST4hGGp6fr8PHchr6B45nPZ9SezT9ps2BZ15xn/O4gwpSee
ZX9+hlJvLjO3dKRDrBY3mPOsx4IbWQ0q+kZDe7nomFCWt0qGI+uWMAUETR07
EcghTgsP+e1tDl0hkQTUpKxkvkq/2zqYz9zx/cKMS135VzL52DTOMtFcjL6L
coVyyE3pg5fv3ylwT+FXt4zPNebaXHDSxxv9NX2khCycaTTl9ywuQOSSkttU
y7CQcCAda04q0X36PJIAUhrakF8/kjI9brzhyoFSawSPcLgKZ+qeAsvCdtBi
B1hnM1sDyupgvAZjOVhn8IDye++rBYebCrfdm798pexEepubxowv6LNeQ6Ig
2wGYjyiU96aRieoYOn3nc2E0BAAuxUrmH6R82DFyIT0e6v5U70Uu4xYv4A80
szP0qDJB9LdnDiKYiF6aeQk3vkFeEHm305cf2KB1mPCNNuZMa4OhZJV0YWZ8
ypPzf2Fw3e83EWn3gPN6xKvhbeXjZwEcImpMRA9y+DA8R/dgE3EaAErdWkR7
ZZWgu82bxGCC59yxBp87qHsmZ8oercypXGpaY8ZniC5p/KkvAlAR4t0/FYz3
GJrVaDbWIQjeBoBgte1NxgimEEPXY4hVQX2y+kUUB8AcNyQIVVb4DY238LDe
B8wMSd6bQtN3AMgIISgSckJD4GSaQKn2j2WQKSF07FP+OUGeg6rb2ihR9lfC
coyliKhwIDTcGKUc/GfyYuWxlokIy/otYfCrStJeIjwPAnKehjhXwpdpD1Pt
nQfAQDSDTwsInCKwM+S0EqbcTiJL8O0bBcwiEEO1PKgJvABdHEekLMFWW3n3
/5+mp9MqPk36q9WYqwC8d4+4J1QyXdOmmZ4gOisadPLwq8dO0/8Bbw2abzUj
vT+ft1sZlXNAvKE8BmeSqp4fOmXzv8iVnYVg/WCfx5DCUu/36UOgdJJURzFT
ud79LEyxzhWLRCZWjX6XOIOVYjlq2Zz3p9gMsgDbhyYLoAOgNs4K9hnyxNq/
gV4APxKQN4vn1U2kOKkccrJnzdCHGog0+M26rA0cemoCf/s6dZLethXAPHAI
yHguMLRbqrxlFQrgO0fpFgJ0Bjl0AsCDmTk9GlsdQcyuoiptcW7QbzsEvi36
8Aq8K7RGknenDzkbPIPWkzQvvJgoII2yP5jbvP90zCvy/1pTzxkQCmDrFiBV
ofkoq2Y0//D4dJLCeV79fcer0Ae2YpzQpyyVDGo6VPQthTQmE9I1WPCDtvrR
gA6k9wAH5WhXESuL9tTzGK6jr339cUI52fsJZ5iwW5EDlDrgrDs7HNtZaOHI
WXrjbrtUSplfbhQWX7bh1JMtO9P3rNuEpiW4HPDp0KNPWMNERfpO29UByxMn
8Q7hFIzcGlWfaNw7AsWvAMLubpy3gHgqRi5KA+H/0WdqIUWmaYG51+NGR8k+
3mPhtmP1OELTe220wbKO9ByXiVzbbRpIE84XwTAISV9LX8B8k1OD9E9b+kgC
bEb21/C9iCZ1UDFdN8E9QLdDw/onzRvYnPp4msekcIsiInuDhAZ66/BGUQYB
z3siislEvZQoiia4tqZUkJ6GCZOn0UJ7y4t1Cz/5kTvK0GY86g5L6G+nty/B
Thi9nUolPHlHRfMAhgqSdHWDmfdn4NEqttHyNS8RwuRry16DuSMonIA0xUCv
9gjvP0qqXvAW6ngRQTEb647903xYcLmF+hCvIjrsCpE+/a/d6XpL1LcrBz1C
hh9Irh6b0nZ7qknCNAJH21RF0T0ugv+YvndrhOb2Sp8gJrqLsgcYvLs0FlmH
rHs6McHMxrJ5Mpq4J9d4SUOLsk86Kjb43AoLKW/jLRo6v+Qb6LJ1kKqlUV/n
XlA0U+pgHa8oZuBkYAjDisPEOkY88ciXos8G+CJIe39CYVnCPMa53jKfQu1m
PtCOCEbfCSACPh2PnOkNmdGsh68Q0keq7fQgxvhbdG2NePSfX1k8ZF47tyHZ
XjtQ+tdTPA9xOsAO+Q5Twrq1b+Sc4r8avIUMA9ygzKviAN04bvK7Dov8Tezs
OODqgP+iYAONZWFXUK7cIKuOL7kEbf3HmEUjVSt26ISWkshINDwshaGMaD2g
+OblHwSgw95r3RF2WAYmthq/S1dnvVH7DO8zfaKWsotXn2x7mDaezueeFLmo
RHEirGGXvxXMA/phbnfHc7q1aIUhWcJmkCSzZD2vtVCGHNcY5o5wFCxL+0lT
pcqa1He0qChfRxFLzNRuCqqxtmPGIS9V6yjVVMPNSXRG39h0KZ28sHOl6mqQ
Mgczpc1kyGi9WSQA6v+IYwxan0PlcCI6Az2C0OWunKE422eo00Z602+PmQgr
S117PC4vY1zEcIV/nibOjIrh3nOahCiSszX4KpqzlJ7dDNJUgsH/8cStMVmi
dHoUBaQvIkhv/9xS3hNnqB+R2tnA5dpU9V8shaOcvMPBHbh7MG3vrTvDqRY5
RmOX7zw/IZeiCyvKKA8NiV3GIAWWh6FnnQUE6e4E7VhpTzvFzlahfa2VuqEl
U/wJ+MZn0mD+YQPM6/qWgLFR0TN4uz4b251wuyt04LIS9OkH2OprFKZVUveV
P68A1l424KqhJ+k=

`pragma protect end_protected
