// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
uV/nqNdmTxAK0LQWFiMpP7IMrKcs8tCd9trRA7AzhzvyE+7f5HuAosWJboiVFILb
zIpIqSnWG7S12f2aXB3jMMumBB82Jb8MZOtK3W22+nRFy0TGTY2SRx/YWQ8tlGi+
VLAZZ2ytZm8HQ0VKoxMzcXMlCZbY24T+slkM1TUKwn6Q0GnUs1Mjuw==
//pragma protect end_key_block
//pragma protect digest_block
GSsLf18hIfuDvnZBbNy37Ryl2FI=
//pragma protect end_digest_block
//pragma protect data_block
FtRMlHEXxMj74ki8le2Gdc1epgXGM4QDT6yT3fFi8xNEViNstIC7dLASelinm8dY
n7H7GfH46Z8UcDtpf3EbCvmpKhQVxoFg7lTm9Hy/2uyS23p0AqZpzpAEVbgOEYgX
i4NYHJbHwc8TUHyiUcPNct9tHlV4YiTxU4v7+sqinsdX9pIh62Jsb+1IYS3H/3ES
+vs/20Q/XIZLpJXFFLGru22ev33pdqCgKcInjKwqesA/379+xra1ZjgoMrldYPek
B/T1a8JJ8XJAWD2pCQatLcIjRDPWWdvOmuyG4i96gmxC8Qnt4ncl72lYnt+hOtHz
M0OhYXGgtRLgoBk72AZySOel9vEC78x21udCShT8HjfOQEryqls46dB2/lcJ2/R/
KHdmGF0NquSSFMongK3Xf8iWgcbSLGLE/Fde95jaTmPdnrKULJTlED0m0NC26vF+
HVrglpSE3wXvFIKPhXvCJBmlamW8ywjY8psXqAcRI52xpFjiRkf1eCYIjMk7RTE/
6A4Dq/HpnNky49LoHnS2mfOmYN2kvIrBg7M7ihd6q7FqhQxeflQxWD2QxxIzLiRz
0l12ahFQOITLCW4hKddgWYn6EYnCMd0bSaeLBnDCqJ6idyyP5RHn4AGA9FmGGOec
GIppdiz9y54bVHNVH54oAZpFPkeCx40RA9sMMvouP2KxDxwY3wru5+QHiK3BUmbt
QCid5FP9m3xjsbhGADGVz5Vk/MWaMW63Tt6mtzEqEsd9eIWBGFvot0fq/v29Uagl
2vz8YUqmlbNEE9wb9nILjMzuwpg4ZKpbRUfMpevrG/AsE8OOywWOgOv3ZpNQJkGH
wHn10E4fu+CjDT+SYFumreVnocZQxwrA8TnWTteb+Ifw7QUgT7ypc1zDxALvLyiC
g/Ck/Hlr8tD3hp24sAsojBoKA7RW77jxYxfvxgoWQSN1aDgNOBwUGPG+aY0Eh6VY
xyVUY+tUcG4Tcfizyh/mSdYkI0FumK+YAZwf6VV7X1loj3dEFvot7Yg8bQtXNBiG
9AvdYeDhADOrJ+NlfKF3E4Y7MwIunzP8xJXnMahWXpAOSKjQR9aN5lzjGPr0PLz7
tKIrZ1qeuB9HhCjizfLacTTaU8jQ3PCDPijGYAHcxLTwDr65NMv1vLQIq+qPxn7k
LNRykaqp4U+jIrG907yOHd7lbYvZtiFOZWikEh8d1fyEzVm1vxP+ZEoZhV8QA9Cp
G3t8UxTLS+zxqDaRFXT0UDkCjPyttfgne2Hp4BEkHQVfwzJJcA5W+MlpTmom/+Q2
F92LAAH5JggYBJ4rYqxOP0x0FI48RbB7qEnYMrBCEP0Wsj585w8RI3DWRFJ4NkaR
RMlQV/dTlWTIoEQW5xtCKr/trkFQC1RsYCzbsQTBAmlmrJ7qNc1U6wWcCbamtXzO
lLdM+NylZYIvV0+QkslEX0B/IZwXt8/DOC7XVzkhR05zFrBK2U7J8WajBNI2jQoQ
RlLWPbHx8mJeWzJ/0hkcXARlD1gFuxutGUXgKgz/iR7WK46z6WgOuj9i8iqI+Ch7
Cwp9JW03n59JWcJSfmB83zBUaCPurCfS6NDJoQCi4QNlBp1EWajUZJmRznteQu0H
w+SdocQLXcHVG0IoRZKRUCR6fLC9Qh7Kjk/zHjSOdVtc7gZM0Q6fO958LiiB4FQf
IY19KC7gv/b90UnTkVIiY/xOd2xFo9fIui2Y2XedofiBCbcnYul6GkaOuUEk8jkR
evSpaSxfEcmw1vCKt13uDUlF8CLmT41fOEZ7dzRuATY/MCzvbh+ZtzAN6IiuTNp1
Kbln1EByTzGkgVbCLTCgQSeXXwmOLyhVRpYillawnWA+CCmveM+/tYJzXSjD7SHw
uRO51rFTLBz6B0co8DJPpFmW0o1PHvvBpHM6Miq3EsPzsHu01NdtwCY4npuswQ8j
4cLvh0xe5ayHgBQBZbwd+HPx6cafEbRKOuFqDL6SvsUZFLXS+wpxcNpBYR2deHJQ
UuN6BoVUOXyBfkXwlVwHTP/KfkT0FDmRKxY7VEyWl6Qcb/wJZDfAsSckI5k6/M9Z
30CTMSTFHoeVfjogEfQHJu7OteET1Zo1Cv1//kPNvGSGc/qB2YFlvlWW4+i1G29A
NnneA8QzCRAoWFI4KOVgl+VjuvXfNZdJ7eHOPqzGkBattfHF5lDwOLXXin61mhFX
65Y9GBzwRBgNPOXWbN4/jdUrDDs0oDSYR+2+oiiYlSaJbDVoRdbez9gs3XMOH70S
nnyu9+DOzDI4T4RtP9xYFmcYTcrCNSddHrWEwdtQxvyWuyiAxgPO0V69JV2lU5pV
mxyffkv9PhTizkY8hYTU2h0EOTOKqFyDnxrtUpA2MhUFA5T+YhSpBVYpZmdafdgz
s/o3Ry75B4klqqKbPHE/0bAJwrF1s1l9FEGRMI+0iu1kwGHUpvX3fzTLvF0IPxC8
to5mPBHQHAkDXMPyVFSTK6LvJn7ELNvX38qXw/HgU1z1uK5k/w94e8d4YViTUlWz
h3DRCCF2SJwO06w5XRTuDdHRRH+n7Pm9lprXN89JGT5v9aGUg5hCZIhl0eQBD6Al
/6YjBYgcr9ct0L0iaA9kPFIPCCY0cCAucVdnMhmzqj7pUD2ByfN2GG5SV3mRTfzI
5kDbxpQ8R4cgNpSCryNUxCI5AEwW9NuF0AeAQBYGTdzjiJec/wMdJqcEE3VAwrSw
zobRsQABkq6MJm/3cvneCAiSVOtysWDYL/iW6wwIpN22cwovBHSgTulBM3LPVdbU
dS5/VO/NaWDLxCffZDftmqceCLQRK8CCITpL9IpneClJxRf3oQFUMVPp5A6ROJib
dZmSFXQK+7UifjURiFBEoen4dlzOYFfGeiAybYWX3FBhqJ5gjm5Fdv5Z53FB0Qo3
aE1BJc5Rrjo3UdwReWSpvDljXHuNBeuMXfm5+IlxivJ3dq8UaK3aHsle6+kQ9nJe
+f8uvqUrHzGs97c++/Pmvtpr3w3We2BdX7s/VrrMTk6dbH1kVXckzwfE1AdIfuD3
YrDdr8kS4QOmQzGsQ3OddSKeqy/7g+xRz6tweB8K7sM/8FGLi00JbkZQ5NSsOn+k
h6fDo1cjEqvkaVqlGPq3L+DQ+C/PMiKxpYtkIBuDllDxNbRz6iI7jgNgHi9LVQXj
8zhQaPy+pK54usvonXsxRA7Payf5qlFeSpCl+Q+nIrjecKP3gCFQFF1BPpR403bb
5w9XvyTEPJje3A4L8gnbqfcsrwkYR5k1XL35DWapzQCOzyeVsm7lW7kLH57EyC95
qW0DUPWBNqSVlrz0fM9ajXTJfmqOWcx/33K2H3zHYmBAq9gY6AZiSgu9Df18SHIB
iJepMAZTpRB5F4sgJczwvr0eqTE4iar0/6uFe4dckMp7oJtnnxUiUJyZR0eh9H1y
Dza+csvm/jVzt8dlUH/6xtmNTsvTBWfJSffyDPqy+/2dRmsZEwb4ZY1KAqs7eRQw
vwJ8d2QyVW0Vz1EfGqZU2rat2NR7miTiA2ebW5fmxtSHIOi9Hv25nFkUCiXp63hc
Z2mfL2218xmIi7fSZ4AAyLC8lVPtueRNOoFpoFXamZbJO4yKQ3avgnuhMx2ruqtm
CZbJ4oBKRWHhxRkiVzXBqziLuSLwWnGBAYDB4xixNJkxOW5drsR96h1p66iJn/7Q
qDQQv+UrpZjomAtKo4wRU6D4QyEpMGsZGxreorJUyY8cg6u+giX4T4xxroB29piA
s6n0rcEGIiqlGeIbBcDH2G1hincNooqDhp0W2ltEk74MURLxrzDBJbh1sJcScHqD
S20KiUurALBwAQUupkG5e2L5F0oI0zfdr2igLa76UyujUypVPKEQQwtRKGmBH3YL
4E0efiw0uZcP6J4a06MONON/NxwdgtujJ0ByjlRelfMpZJp0modppDEACgMZYYiO
9uUEQzCHG1H2zcDEXsiLUis/rWV50R7d+lmxUumw/NLaWAg4Bmc1/EjHEpQ9fNiy
sOomdtCLgZs+XtITtuM9vQxK9n5KVS49FhsswKT6wLXpRvE+/oOR34FI5GdDLf8b
254/eF5qVOUTY3mfH/g+PkmrWdQ8UJ2hHXKhWK3ResL3whQUA7cUqO2HoywKU1bH
vn021bocFhLZv4IAd8OQXdLc3nYlUGiTX9p9PrwpTpR5iIsdvcsgeQN/eIorU1Ws
I9l6boGp7up+V1wklSjpCTerDlbfd3RvDIp3htFqKWjA8QworwgJ8JBKX+UusK49
wAdAE7IK2T7EAPjOFndGLGGSGNYadh1X3bqC1oriJfb6SA+cRPVTD0EJ0azwq4+l
QC6vDMoshiW7CHQ1/uROGsaQgiJ21mh+UsXZjg8yfa61vWhxldi0nQu7SW61PcTE
lY9ZPd+A/3Y9yWVsd8RJgW/yUT1rbH5gMdiKD7+H3Sc6g81UJO9qmKiTFC36x0mr
AUxxD3/3YNp8SCitGMiSvsb4jdg8Qk7JQj9WJTTNZg9gaX5TNtXKyS8yEiz0/0VB
MvtAfYnEVIgJOzIT2f3IZ7Arxq5zYfGcIc8s3DMnJMWq8NvDC+9R/Hm0vfbBF249
gSDfiXmeoJBdFelH1RVc96id6/caofZZuGRjIcA2mbEGX1ewP25z5iOq3XLa8Wr0
DCzClXoLX8nzoeCmvXAJNkweF0CAukAgW1LdW5aBQqadrjvBn2JOEHHcVJma9vH6
8vvgm6junjdSwkdIRIld8GsWDXb2+95DWZxdyR/DVqm9tinxTt7AUCYG11XKj4pg
9y/rnxuGhUXqUmeQpkVkJnoQsOL/4uKFV02opmNYp4qhmhm1hHSIZ0THPVN1FMg9
1dVNtSaie6ovU6ebYh2E+wGmornMRG74klbdkIaAHpTI4phOs/zRi/JRh0OoPxCL
sWnVgdBkVRi0FRp9V8iS08NitbP7FF17/bPf/LIOHr2KLM7+Oxgj3o72sZeNGNkG
aBoRKK1AclGrRsEgIs5+ejewr2g1NA1FS2G50SGZIbZcMw7VYGAHjBHoucgjYsqC
yTuRQwLTXqHiT2TiMppEyDLpZNeX3UaIBerJcQDd2wfcumE9bxbifzxxFPgducXD
pVJHQr1SR4y3jjuOfPW/Bcfw4sl6xqBtuz/wA+CCz8YVN9QVpHG5+xAbB3cNAt2y
oAyz9eeyjeSQFKwLWvl63INbsZ5H8mPl4GXK926pRYRiOIrbyZbpqBjwVRMpIV0+
suPHb3JZJw9+EKEoPLLFaBnySw4nRGQU5kKl+dssHds2tApKeOrAD6Mh5g14+XVP
k5Pncq3v6/UOyDeStCd9MGZn/5zYQXOwTz7plELnbtOR5drdJhUz+fH6gVn4Kd9i
fTi+w8k3QSA2tCCmrptkiL2veOTx5hPfwq/yuui72qPYhdlZgzgJAqcYJeSRSmpE
wkSZ7q8T/mvi6zsYDmaC+ZSuC2ZcA1bAcRPXJKr5+xzl618khVAkSxEDuBVktYaa
F5Us9qslS38H8z3lJwQv3biTXVE1uDgTrvHrflh+2NahVOxALMpat/C33x9H/Vg2
7bQ4jJUl/f6JGT8DWKDGcttXEoOlsxWg5nzzmQ/HCoi6N+k25Mnu3oRuSFksrObA
kH13nigxSCtQbjxIL8k3PqS3i91sEax3dEspyiJ2zaKwpVwWFT10OX/hmAi2GPBC
81sOj+g5D1OvK2IHEEVNg2oXfzF5rvTwwRZeZLhb+uPSlamo3niptzKnM272Mr1w
fDbeq4IFXB7FGS6RY7NS47x61D0slj90tujfXctlh7e75TLtH4mMEv6/3WQ93/XD
levHReS4Njq6wdY1wBe8SkVvEDFfrNn41vS7aBEMNPgxsyrz6R8d6a13o2mCdrlW
FEk0Pcajgx72nH5CF0bwVqFfiSuaJ8wAXY2+zGfrZ+qls1FUVyzbbwualapNggFx
KDw1Ebak25qFhODmPqr32GxdUEDqu25kl1hXk3x7d0M9/mS1hKVRB4s3cX34xCmx
PCw8OHOzSH6F4gwwFStn4JIsSIeuzfb4FNmalJqEleJXWWaldNNWwqlwCL1S3Onr
I7s/OJGveH61ROV8eaXjN6QRDFb641f1r0m+CCUgvqluxXyu1NEf4qnRkHgltqa4
2WTyG3qlD9MlvUY1+aPEk8VPw60DnEiyS08OnYEy8KfCI3xSNQrF5w2ppWzOtuO4
u26TyA5tElcs+QeZNqoA9w7ACPrvLZ72TEeE5AZlTNTOPbq0VoPuULyQxUmw+ksR
P8HffwEDISPVNKhHIgjl7aHSGqLH4vfcNDzb1hh4q2IL1NuQ8TiIoaWGAJwDvuFD
dc8Ai3FnKqrc+Kk8hlQA3MIs6HnmP/t3PGnkzum0uc+qvl6VaqL339ngMXcJLktc
bBg3CXwHv0tmsYzK0PNCEptGAtQ995DqJTPJg9HA79Jo039kcqaPg7EdEhw8+7hk
YeB1yunhKCRcvT99scvUl72K9DKeO6g+mMbCQMRO8aW4jcBJjc7BFSX7q/eGT1UB
LgldO3BrZ+/SMGaDvhaC57mgiIpNSftU2XyypmIyMsB2pt9DdaCZij07djZCYcSK
dznxM1GCqrzZiNBqirn//E39VdDFDU+sw8ITkUvtXeKOrkYefp2sG9rlnH6hvn23
dLwxdGOsyExoVZg+WubIbtyGUXa/F33aLsnDGYFhBQWx8R5LZvi3g4zQbNiYCvPd
rOuPMHQz/07T7J4GIr7M0+v+sKZIDUUdcGnGx5/KvDr+RITKb7a0IRdM6jU2peq8
ex+TiLrO/j+Oz1zEbjR6/pTKvbwpRXNLTuvSwU99UD4vb+sH931i7Q+a8NKrKpQb
iJY/u//A0XsZADnjOmSOoRMZB1U9rZnE4442skBJcFTDO/API7x3M8YZVwQEPUcA
MPNiMnplvTBO0AYgsl97ySfe/ab0VY7kVhOlQF1yg4wH3mmKVIN9TAwy1Seu6BjE
CUjNG/dWKcmV6x8NrJ8vMZMHh1bd3/UA1irdxOvPiSlliNXQOXBMVglsDJLPeNvG
XKpYJOLmyfG4w4yttejOWhqWn8LfWZO1vBZ5JNz3LFPOjakpDVYnle5gY4kDgh1Y
6vEJbbzDM3FM9ZJPe1kN0iO6VSTnp1b4do4+zu5Clt06R1b1tWaof6GH2Z0HiQxv
ot7aJag/Xo3FlIrnoaig+ho8mDkLyonqHo9At/dwaY72rDf7MM+kckSgWkVYGQx4
u97nMZny7o8V+HvF1+O7kcRFsuimOOV3SF5DLAM5X0zjjbRSMjcLlKTKCHQtvfSu
5yVdC4wwFFRuI/dlcEz4W989uRtMZJocrJ+cgKuV/i2Eqt+tM1czLUJaPrnoz6mi
VG6St1UjBJCorCsBZ+e04CRgGm1dccOUlbPnFrTCS7+RZtJ9YzLs7B1FE5Au9dnI
48HJivrgK5WQn+aWc+45HLZFeRqTKxUNZlVEZNDrvDN7p3ixCcNUUkshqeyQBwaA
NiU1PDrNxngY3jSXXwODpstfCR0rYlwIZYvvjzsPbq2HAKY3IbZawMSfK5NWhCFE
I0x3ZX02THZWMb9aIsD16h5XM/6svs5nk1eEAMKvaVkR1Qny+6sexWDsZDCm96pX
vKp3mHN2qNPTwVbhsEFJ4ox8HTOQlxyL8GyCDpb3N25QfXHHfZzeHzdvun/AYPnN
R6794y8XxP5ChPC5hz4l6J2vQ1t0h08nWa9O91tdah5MnT/2r0TUBGM7j9OC3di9
rSrId0Jpsw7BXmUgry/ve8n1Zv5CT6S4HYNGFRT5WWaalvj9eJU/v4uqHMpcaXlo
rgTgBLBG6GeZvOIgBZNeIGgdZR0VzXL39WpMJ//8ph4zj2QeBitmvIQ2jE2ao8rg
uyMoVkiZuGoCmIqhQeoT38aFM6eZ8di3Ao38GIaw4UAUAkZ/RnILJ+T5K/LE6wR3
jEykNqfiVhPQp2OSiM/h2QDL2JOrsrsvFjkfLpMoKlI1JaMna3hlUOBwh8tP46D/
FjZTezIiBLo4MRmn+UGEe797NndT6GPIfN0BEc2r59BnCtW+woaGsw3pMBUsdQQ5
VRVflttTx1bs9hNbkccMeavljZjfSCI9KBMMSIsSl2+UEI+NXelAL16xquXmIPsz
wA+s6Ebrrt/P22kXspRuE6vBvVMKmht0cuDTUUoNPN1NGrm8JSyqI4XORl4EI1j7
5axAg/Rka62EFfVQYFc+Z09VqQ9Jx7KNkXIFlXxxmRQmmAQfaDndEmhDsbxt7SNu
RTu0CXrOXOdv6JIexNrnJN3a/JbqK66Hp7rYKbsXJ3iZeLuz+oAMdCNx1Bxo1Tgt
r1mV/yee3SCbkICpYIuzERuhZKSNaAl6FoVYntSx2dJ1gDlHUuOAcduPMzbTl5l+
085ZHVA4vQL3XtK6gPE+f/uuVnNEaUJtXR6wr+0vPq8NxCz6Now7y1xcD3P+NgZp
a5dij5CT4EIbPCCA/z/Y1lLZXZOlO6vqv0yqwUU7OxGYKqsjNQyWrAI7zru4y/04
zP9wZ9zQC2RRZv4L23ENPDv9VV+8MkUaWXzOKyKxbmnuggG8EwMM0TwFMBQxEEXV
VZFsusBs9a9F/QV5pG0Gk6B+McI25AdiSZVsHIFibvOQSBz94s2NNqlL8TkuNGRJ
n68dHpQPgNHtg3egmPNiJDw/MvfWm+if+UZl3eM6b3K9sAY3JEMdguMMH6eEYIQ8
+XB6zT9mChKwmUdyY4Ptu1NtN9BW/tEEVDaeZW/L3XI5rxgTW5BAKQuqMIDM1Db8
ZbclvqYLDynsh2AmoMZqGTyxSPXDUMEk8eyEUa+Wa/Dk782qm11vLzoHYKkU2gDj
Q1uOwQXysCwUVXYVzNNQWkkBUG70qnr4Dy6++eHsGR7NMa7jYReTslAai8S2o/3B
9gP1JcJoDeQaqS1tSPBE6iRAUjiKCp5e76v7cKmm9H3k/LoxSs8PRLYpfU3qhEKp
C1J9tmkNI//M8jiZ7kEBoZe9ImjeVxvKD2KxKs7xVDsdc7Z1unYXnY1srbz1mR6G
alvCvEAnmhmCHatL/vxmqXjScjlbJiVEm54s8CcOp7m1FuBbRcXK7BUqplHgVeN6
11GTUzl64Y5hFhCo3xc/aPsNkrab2YJqM2eFJ7GfGblYMMSfC8sQagjQqt6fwXCa
ArL5jisCIgD5mfli1IG3O8Q7/eTspECsKi6EtZmcksombM6rCVrRR3c5JwdOMsZG
pFQJbk1TT02gcNZeOK8tE5v41K6PYnzQMCjaQ+CP3CD1sVVNm4rimVR0UMl3Ujo/
Sv9K+5KP7A0on69/QOLGzaKc4KH/B3h2K2VDCos26agjhys+4uCWgNBjqpRsUgP+
W6l7/eEMpvBzQ4AIt7/I5e1wlylRUPhWAHirm0tPow5oOV96OfB4Gm2xa8PB8J9e
kFdjo4O9h9y27/JyhKVApPiGnPJGPMLHJRN3sIs4pJwQo/SvgijkFdDUS6Fl4w1J
KdbiehEvMEapeeX576x6bhljHvxAo45BKrzi9PO1LjSyBkVkmK1WTUrWdTtYVg69
XQEo1RSwUM52LRS3J8bX/A==
//pragma protect end_data_block
//pragma protect digest_block
9fehLWH40Qm9K8xTzSSAFr8WrDc=
//pragma protect end_digest_block
//pragma protect end_protected
