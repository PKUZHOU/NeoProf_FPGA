`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
Fb8cA3rqqEGNHTMqESj/PQF88qqElaVVIAvBB4j8rLDoIC4qyWQcYg/k0BDTYl86
gLzHpiA8pcJUF4NuM9xffLHDUBXeaU33ips16YdU5KkCIYmmT5MWnpU9xSF1JdxS
rtZjR8MEPOw9mMHvHsd/7C0p61DoNN0sGP1bLRC0RDk=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 6224), data_block
Ouv5PpvFv1cVyQWD1z34gAzkb7P+d84bEnz0+6NBcKFSh9jGDcdDBtdBHFOzjxod
WE9e8UmElVnjG3whfxqfnA9NCl3DttMVbR9zWqcP6UUVN3NHpkV5W3p8CLRvV1jT
DS5syaKNOYk2+g2rbn/534fhoca5R5Zyhui/M2uynPCBylfuqG/i5lmz0rd4ONAf
yBqXWKnl2qIV/p2XxGL+aBuQGYx/CEi9xS6xPy2i0iA+Mda+p2csSw0k/h0TOtbk
vKUx+gAHLdSgjtk1wO2ShxQG6oX/yR+29/Og7d+lCNs24/SbCMqBy1USdd26joGv
RUISse4MnA9st+tWyYe2sW01Yg7kS0iMmkuC9NbUM3fDgAW5ulRs2IdrZ6O5UhIi
e6/X8v1met7rBUFRbLhSxXTkxONCl4qapUwFW3HzXNDpOXueSlnLvsB+KxzMgMtm
rNAll8KpOilXTIDgQ/jU26JXERgTp+fnDy/Fav4Ih5z3+N3yHN11FVsjpzZn33ZO
xFbQQakusZAl6vAz2OY0RcU/65sE+GtSiuNItXMjBb8iGXF2u/NXTWeRIrRAXRQT
odoij9JQ2B1rYVjHaslt+uGMpX2al4dxkvjlaZMwARqzP8JjhdHgWVDWBqkNVZer
3URqs2xzlxcpSMBSjTsbUbgS0lsyBqiJv+yH8WJXwNmoZ0RvlTUd5tk622Cp4xA1
AmK/nUkYkB5ci+4Qmj8Lw+ikcBzYsN/LBI7SsPr6p84H2e/WqyDI8httqxhZJ+AD
SvIn2alP3zaoBA0os8Pq2GLlRwWj+1yXOxQ7kXGowny2fjqt+dIsSwc89GZbfxk9
6I2nUi1h8IqUmkqu9GKcHUWUI+KLD3oIJd3XPDkpZQOQv/O/jQxS6hMd98Lp8yin
6TzxuF6K0h4yz11Kyg9+qLz/BbMyLqp1OHoKOaQ/wlPAmZ92aJJ9N0KBs32P2f6g
gPb7stPDIxV95JdMzJhaYughseVdCLCeUpeJvmVAxbhfqnn04pwIrdh341eTTmV4
LHiqaph03v3+l1Egvi86CTiKw9otNO1Bqigosyu0W4OG48eZ1Njv+EtrmBf1SvdH
Lg68Du55Lo91TmNYuI5FY9NR6sUbFpTKyNgaqeTCj4s/gMiuY+AyWv49XH59f2T6
7wfDAcg+qZyemnkYXxPGoIu2JMRE7EHh9kGPyZIFSz7zIV4r8lbA1Vnh3fEw0jc5
fOuh7i+J0drCRYpLwT9A32iynacKbxwTE/eirjt62YQ62w3sF2QeRr3EpYO3Hgc/
8d7YFWhHcGhdfULe7eBcFU81cPPTQ/H4CKkEXnnvaYE7d3134Cc6OoRs/87N6f+J
5dnYFs6eIQWcRB2De9qalSpzAeDQaL14DkFycgzkoQ1gsXurZGLyZZcldPa2olZW
nPvIYvUhXeePB41iMpbGnn37goFqnB//T2Cte67mlFBBEICJUzRwlTmG4aNhwlia
+8M3G2H37aXP9jiGOhBe769VUVlBnfrng5NA+DyfvVj57hneCECSsUB9GjHmiXMY
b92hSNHnpjBTUpwrKzFOzMNOnm5SmcvOZ4SlHvQ7dixAk9dDPCv2Wl4VjxSZ3qqX
9SfN269GDYhdZC7djAU6yWP9fEhGLljAvadmjDM65JxuogHjOqw+Sjipx8g7O13u
ZhEJg+MBhH2c00c0UAfsONIEwmLRwE97BLuRaoO/hXGGOQG4LfZAukXoyksZzl7R
2BL4JuKkTilUgJhVeFqJy8Q+qBWy2oB5qYztqSGHihRRPXr9Br+isV+nVz/HznDs
/BUUJ/QH/6pw5ownoF5RkdVMpLg1Dt93i3o9pz+t9X5YXtnMQDfNyCJZlTIoD7ht
bhtsrfJ9FpbPTpnW1w1JXHMitcdf3P6IWD9NA/QH0JHpBvWtjYUt4leGAD/rL69e
HO2u0Od11oKcJwmxBikQ0Gp9oJ6xXDcrsE/kQgmekheuLN2wkVO+zu16JZStTKip
X6Zh4A0Nhb3T8i58kLkPqjORntsFNWCT7ydvDsM7FT9zwoASb8NrVjwynTewmeqk
zLXImIqaAStNX9wZaFucrT4Ch6HMB5rKMCqOfTGXTCDs6hfCm88/eXMC+M/CjfhW
WEYPF5ICCQ2yrmzz2SbFV4u2B5l3u5EVrjq4miDrQZRMFAySE8RxaoTKvedYOxFG
PjEcvjiSrCcQgkCISslA5+FIaQt8mnf2wohu05UzriHh3udJNjxv8R1d6Y8zTJAk
FyTULxXBttythwIzJG1tUYZkeoZdmgSOPmclVZSpnec2SK3O0agWXeyQHJMYrcQe
pBLNiuydudCt7n1QCdsFVdIpeZopxmGwMsQ7fZKkXkLykmTjx0ys0RVM2nCB351s
1+LBO5E+sfWmazmoAZO/n7gt/yleBUA/KkN2tyq1axkCWHvMp9FcqWnyu4hGnAIP
MRteymr+wOjRQsMcWKV7TmtG520+FM1QOU2OumCXFMWQYLYeI7d6m5w1CiMFU4hU
g0A33/7MRbVwkDcsCQiF0HYw3x5uBooHtaoeTm94QmuoBca9C+ykEDLWvtj9twyP
6Fl6r6o9neANCL9qB+LkE/WkRtV3vMaF/NVYHp/7KxAVwPq9L+qnZI+C2loBkuL2
zLvJkFwZNFUmvP4Kcqi3N65U948CERyZuMbpyoYTlUJxFvSSes7QplL6rbQIECxz
/PwP5IoGCgDpalsOqHXBx1lAX7R5UjqyYkrraE5u6qCCKRZLEVkSx3qijJNBKU5o
2scZ1/5cELXTdtXh+fIxpg7zdKMmR9DfojXSf7VhU0T3kVSdy9WJ6nGTPhJOabNz
GeXZv912nKSfotcV1o1Fp76Jo3okNH0Vje5bGU9yVR9z9DH6CiWoUu//9PwwF2Y1
D/3FjX0GN8Vwf4rr2t0FEQM+OvCMCme0XXOKeEbT9xAf0hGk+4SiYLgRY0UNs10h
Er8N/ACcUUyVfCatkLosa5PQFjMP3salQq+/n6+jtAH5KVSAzUeIOptjUR4Q9zuR
APoeZWJ1sb8P9YyvZM6P3bUpjdvIaAZyiZTOLhUcceQ1yg9wMnjxsDGUo3qroynH
9giAc8kRcLu6fH5NXdkAjwnJ0fU3bEpwnKEDNw84zJauF+Y9Pdx02EHyl1JrcX8U
A7xHgrDz/oBqtAMN36XChRwYwdkqICg/0zVvSsL5BPiS3E/hYUeYLQ7pi8dFoIwE
wJFcdjYmUbFvh70/vmKatnRIymB6Ljz2vgw2z+FHC6Y/rrnQ1FGqAyJHHG819UiZ
ubUcMNXVSNuYcqm3R/EZhR/r6fHIJWOdEWWpZozw+HRx82dR//vrZkqPFvHGy764
C1NceinECyuiDsXrK3SUAHtC733iJVwoLvHaNEynbhziLU0CwIUiD2eW5aLxbFb3
fRV1vJgmmepuFmWB2dQ1Nxa31PLmCYRsOkK/VbuHIfrCq5XsbixS40oSKWWJrNqp
0qhlaA3BnhPaRjaVghQzBCKW3usoLVflsZvVind1vWoX1sYPEyFe6VJFCDykoRcj
zDH7GM1pID3YXOZXRmF8KdDrNwiYDDKL4sK8GfAd0lh4WXOwpmd8fFWoZUD2zu+7
GQEoYEZuVzwSWIas6kA1VinCULg3/WRBNTfesGUcLW5haw+qmxbpPdA0JazP5vef
L5Ut4yLcwsyWbIvQyWfyBm+a2T3vj6W+0tjff/XPeYoehJlrpTIVUeire79V7h2D
9YNBARbAu2uPaRDKRpfNxYOmkXh6ZWB3z3B8FsI+RiMbe3VdpvQcKdbnYzSj3i1s
zoodCH1o0s3iVuwblN9MelTwNect1ZoE9qWXhlRa7arVTe1lhCD0a1Eq2HTzqqCg
G6/NWCtIOJTXiPYG6hAtqOSCdhiezakgqN7TsB9N1paaAnLwdXS7h4iKUOcMtyNh
9JTdoNull/RwmvWIQ2lFENCAPdggo8JrCwlcKEnFzh2gXD3VyS/jpRWNbF6tMXJS
QiG88sfmgE2MX2R8efREWlgOJ7RVr8/8LW4jEf4b5fWsRCjbGW9MFsFdJCDRLNFE
zxZOnxUJSV2oENoPCUSSkvM1Jl1leCZzj69Vu0E9NElwekoDbWGGxv/J6mHMWMLr
qWCtv2ocqDN9BJZk3i22m4Kewb597J5Q8pfkX/p3bie4HVSLNU2nVXKOHfSkZUy9
mJZXpWISbdo946AxLwd9QMgfWLm4QIOfitNBWnkiXAKr2HGtZgDBNbtePYqofuxE
pGsMHs50FJLLRp8v9CsoCmb+Rs6kpiaIYzz4pXr9Qnpso53HivEqgUnS6GJw3XLK
AAYMbvcJajr2eDfOBfYOcAagzOdT6j71B9qETpCRb7yHG+1t4Spm7qnapxRNs5pT
XFrLizYqjrWyChHMGwOh9iZ1bDkxcEsOGIaBw/vRZwMEIC9j3s3CSP1umGLHHZKk
gvgflDHAcSxnu3fxmqxSY1tX+qlQUgELxQenk4db2dXZ253cN8k6+o2Nhylk/D9G
MfmsYswh5oOKVQOFWkAp28MdPxBXkgqAYULGCLNARyxFXtUaSz3uQPvon8aUciaG
vk0LKkvXhhGOZc6rsQE5UfqsP3Je/m2zitOlsw5BlaE5rvH4KvKmqOyG+lcbPEMU
+SwploTDNy5VgQheH0OFCMRErFcD3WYDdLWdPuyYl9U+z1Ba8CLYJZsgEunWEUUq
ezqFZAwjEMFHyKDK0C+VyD+nrJfa29YMHdq36Nwy0wA+CkCL1k7jZceBz4Pttemd
SpVighjI/+gDI1es4zLjGAx4FCaK4cpN3/dS3VopAhBc28r1WLasvNWCTWLa1gka
3QBuTqFCf5+4MC+3KmhhMhtzGcfnuTezMtnU3wACSR17rVz/Z8cRqtHYAwRW6RP9
aXt4bK3mvlLihcL4dma33VD/g8cfS2NZr4jGWQze+00GNu67ioPTTGrHVgh1P2Et
bqJ/zPFeBztREeBrmpfPcAmDyHtnwcTi+qPbTgNjn+Q/3jM4xzNgCJFEP73z9tpG
gWi8CFL14ATI25w+bjkLSqGZ2HqqZ6jZlvy+/OjERgM1H45pfk8KY24IdAXsC9nI
KLEdF+jIObJLyx8QEWsBy4nMlqyfXj7Br8r4bWL7KRgvOvI0vswwaZqS7flNIXho
OpiRb7sIs+Pst99mtbJAZzyVMT3JhzFeesdfDmCcsKNdwAjKUQ/IybtTRc7ozTUm
w3siauNqlbbQpMmJRTVuR4+7LnMC+oBLB501EzKvJk/QZEqB71SOhEEbPvKgBn8K
W+H5fKdvL7T52uaZgbn8sDTX/xHe/O39QFx7LpxW7JgvQY6lN1d1GmJ+IOL+La4f
J86AREaRwkG9/XCcPzfVixl4lDnBbWODgFoUR2/nXG3aQZocfz5io4yw9uw/1Bdr
zYgZgW3MntSoAg3JsU++8k+lMr6nuDRlMMI3ujFNAAbx/GCtYkrQAt4NfJPRThoq
Y6WzxA+9AIz1BiRXa7fySzIFbA7ZqnvaRznqLRmfoIa0fZ3Df5Ol7VXTj02KD+L4
LluiysRyPhStDy7wPWoZN9SMDdCNo7f2GO/C81KCoZAJXIiwH6gyP9unk7mfBVLx
UhYtBS6EV3jCSsbub2OJMOrEKAVnGndEWdWX4nc7AgYMLI1jOyK8Jp/ABiUVDVYN
TG8p4gnyJP7AgYVapr4Xek3YLv+4rD7OqQAndi+Rlak1h8nFJW741i8uji3fSB8D
zCeiXMN+Rn3l4NuHzrtbdElNf3khYyeMtrX5R8MjQs9Q/PNWUeRJsB3aRozMpJS8
XphpxR03rCSuoDGU7spfwBWbFT1GoHUbHiouo1Qc/ijHhuHYbwDiIsOZiresnq47
BfZ5fI9TNRFlPKtYKSlH24mIeAOhQj8it6dO2k36yaQ4wVSxxYyUfnshN4LPjqtf
3b+V9EoGzkAQRVJHcr01odANuCUSqCp2nxzLkXZcY7m/djg2dFiDImTSINWzZnLP
QsLMYFXxPXQ6HbVdSoqELrjO6TshWmGw3nODCDuMlXRPHx40zmyp7c/LwcGGG6/J
neyogjstMqLpLPBuT8omhpgpqrKi/xlkUaCHRZEtVnbCPRlcOgoVDnLaS/qi1pYW
7zYDAeT7Xu2ZbWqXZfS0zWM8wI5kgA+uju1JllzKjeY8ug4s1G2qeY6M18GZc466
OtyIrerSfIgiFbFrpGjDQriWcMeT6ojZ5SiHU9ak6vMDlQ0DVgI6W/6Ez/cSSfaG
W+56N+ZgX8n4vXazd5rWGST4J/np1UBOjhoh9FXScbL5hDm40wMVv5QyhvhIO5WK
LMIVii1Khdy7zkMh26iLKGf3AO2Zy05HExl/gKHoDJZ5lQ2vnqRbEJtt0u+V3rki
4x/DKjzNZbLXrijvuzrfbwNQCgv1W1m9uxm+lc9O/F226PsfyzJSOkupqSRU5aBS
+Yo6wa7rfdkbqmAV0IuOZEzag/38ydNwxmxmVI9lZZBncJK72+ma1/6QHj+8aLt9
26MEcWzfej8XTdnk7kAKsxDPCBVKtaeRh+PR5RWOVYHjV17IaIn1dUhil2IoPNXS
MhmJ3Di6GkLi0GRdhDaW3RXnizWSLtO5fTiCSbJ4+W8deCsd4wTVxkmVEgOV9F0R
yZxUUADCt1TfpGLXG+bSagqiWNH5Ody8TvGJg+T5L97ejV9Ay6ZQZ1WgMw3JUJyx
0CxihWzISH25fatPelgx3NvTHrSMRsWXdzo/L+H/NolBArq1SGtkEQyIsNrWpt0z
obotS87q3S4tmUVr4RZVEGH354BCt2Zy3wRBNqOrNB81eSTVLLh7CHlTiZqwp1QG
V/UYYBku6rqPNOebZhjRcy5So/KX+VyUCkj0PWXakx6tjZuvSHKXCN705po0iNsz
2oH8QvZliyd3o1BwAWclS+7gR042WhYa0cUF0Kw8gzvW+rSlJlzDZjvprj5yo1hv
SVzrEITLv1wtFJb89AzDeBI5G0C/cYQ6nAMz5PCOf0sfI6nIK92m3QID11ejmRL6
m7rUTvuHBKvD3tlQRPBdg3u1vfW43k1ElpzdQS4RqeQ8Cz10/0Eeyb81vRo1lcGM
Og45tycp5h8o7Czle+jHLj73flTpUu8oUvc2Kb/ZxaxDkpSvwxszzXoZuLplppu+
hnKzMdTmg7w5WqdFqaGu1dWiVTbWAnt51F17WMhh0vp7Fnd8KO/Tipd8dyCnKZFE
lwi2jvwVPuVko2kfFA8ccn4o0aZizHks1cQBFrYK+lGzwQo+McLXblwYTlyagzfF
6VLZWBXyj55OGaOXDSLBsgYIrZj36t+u9Oxcba6KvWcvr1aPdcNhk8HFrGXBtNyZ
8DX/BK8E9/VzfOb05l7cWcNWiaAr4EjZvoVH2nfigpkA5tlMRdmCbEmUge5PbWZJ
YjDtZpQHeLxwOIc28NqqyggU310NG1Eo6TxT33vk1AcChnb9VR4DA4kL+k+UWDVb
qbWY5w9ITiaIDt9AOV8r073MQRwAUK6BYN85fmdF4aQR3YIEPjL/+DwxE9EAzRt1
YqLY43I/s9y5+YVmMLQdzAl/V6O+vlm1N+oxScOBLtAEbr9Mzu06IY5Lfe8duQAv
3NqbLuglErOVgwTKzavicb+1FLx/H6MzCQh2wDx2TROts8YCSwMLp0zBI5ne99ix
pSEErg+vATypJZwNIYOW9sqLSk9x5iUpQsLmyACGRM+UoBecgdl+5ub8wiw9YUc0
GyxxQbmWiGreB6Qn6mcov7FCOdJnY5sPKWVYmeAT+1Se3B6EuSg1/hMGRCyKhlQx
LMngJs1ZXysvqexiCtpxz0hoK61K/qzNszGmaHz2pA4nfv26T1+mn4e+6aNNpGV2
aIqxnwXZvuE0JIWirNYcoSSvXKdtxTBCzp/jgRif68IEQvbgTu1dHmxtu4drlPji
Za3Ld7JjilnprX87eZwdjB9oEODma7//T8fhS0eVZT4omb+ZK70/g8a7KfKe6Xgn
s6ap5S4Tl7tLifDz4EgRg/jPZaXYYbmV7qIbH+7LxDlv8FQspRTYrRU09rRVlMPb
WrGYJBxysvTJdjNqR2ukus2PAOYmxDh8QYsNxlXIXRqDdNInwq16WoW5GO7M+djJ
heqb5NvdQIld1qOUgIY1WANlhUbWtRyW47gVxrg1mTjsMs/8XN6LFXwmegNQeV8P
81+WTDD/MYJrwGzfWC2zq6cAKvCWcLvcc+xjezkxrpsXgVcR4KE/FsXfxO5MCrBc
lM+bJAuHGOZFkFP/652R9X7JBjsiH97wWht1A02Sok0qthnWJ1QvKETa027kDBt9
Nqab/0ddqtoa681wQgw66pH6AAplA9HPQrSIPWodbMk=
`pragma protect end_protected
