// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
DvDQz+dY8XsU5AnUCtS7w3n0IMVtoH4bu8gb+UK1PBiN1Yt6uMZWFGt+AGBq
qgJaWcXenpBW6+aRLDkw1PNeJ8V6b//n/frDzV/KymqiYW+vqYvngwoWS5E4
xBnda/QNmPrKe09xVaM9+oiJF+wOJBqcQ5Ws7tJVhfEEx13F45X+A3BLlbbY
M7v9mFQFfO1YW0b6sFekbIT+G0uWFGLEJKYwGd5cgFpw7lJ4Mu7kpi99XZaf
ieAALHlUcKyTwJ16AwRUw89P+pdPICYzIW2FomdM2Bwn1VjIE/uW6tThWgvL
DdTpoicTqrN17uRnrHn7egO5FknomEvKL2aG4/p2Ww==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Tgw6ffW3qYLGhKLnwVnW4GVr23Jb4aDdyxrNIPNaSXD/J9ttAdk1VwnW+zm7
ECjft4jXoQBUUMHR0EoMFSxf96tKo0VJxa+wL4QrN6BK9IDozFLGSluRNV+W
H5rXr+DX6YtDHwRr2HWH1cAQ4MOcaEtSBn00WCfv4l5eRKxzCrTOGCOnxj3n
lsCAtv8HgZAqvibWoFndgYg/bYuzgnxqljhB0EoOW7WQgXa6ExvxDz1wu2iz
+sjail7iEgGogL5VAyCLZUNeEW1Q2wSWCgXeBj/1PALKb+iLRgc84kOVN2nj
kQ3JT1F8IbgsC3dOWQTUXpRV2/oqFRANepw5pj4uNg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KLAOPoehSPMEh4BjDT261KrJqrDIuXaQcJNYgK5CPaljjzsdf4ipNCkXrqbA
fUhaq8f3KDnNOMHFAwW/Kc0evjY8YJoByZrtLZxxTpfXymavGOhosYe9c2C5
gBC9cVuvWolAWlPMszzs1Q3WHXhu2VCL/KYklDsbmwgxcxY6xXTawxzrb3L+
V9/JxHbDXIkgbLHr0ezHwBHduikN29nBq6Xk39xnSTNiCABnhEBvSQu8W1O2
Ov+F8pgvhMIB5h7+4qooXJnIPPrqZzLjiPvw3300EWkZV38ELUIK75rhatm1
WZNk+2COwwlmuEj3MiL4cQmcW0ri89XlvWwzsWdkIg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
geNq7nNPpD3AkUPUED49D9eSX0FvpO9MoNODVmYhgNJzbl5XIbT6h4gp9iN6
n58L4kDO7z63WShZeDWrz3tk/Q3IcewoSF8zyNaFN3bgyf5RbEM7SUeYPJ+0
acHl6TtEbOliHezKi87rHlc1M/pplcFcXm2FnD6Rymu8eRpEZ9I=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
PQBtBm8XfAXbnIO94GH5C5EqZIzHmyMaJPkZoHnRfSq5P/6rTkIj3bFTaKKZ
8EY2AI4htEmY/HaZc/tRK7Rdjw690eQXTEL31VrreXLIPin0bup/hZLa4ObX
+ejMmDtSpmjjCjYH9j6MjKWyIc40B7ng6tG2pcWjT/gGDIV3IBoeWm4FUCJ0
37gmLSWQd5w5IHVPW8WJwnOIctYbscdLN3DyL4vPgVUQU34xatQQ5B2SRLqC
G9Vsp8eSEqBYuoCUpa+W/AiwWcMylL2UCVvAlta7wZ9fjuLGafvdP51lr1EZ
jILDybQv5Z1JQNHfrvey084H3iU/wa483pJ44MjQAu9j8YrF1QIKhSaFwHGo
uOjBlmNUkDurn9tQHzkjk98l0TRdspXH5esoqsoBBU2z/H5CEFE2woeBdMbc
gETAN+ZTKawqP0FfL0+9x8OZQDgVpD7qW5nLtGUnKO/mQhS8F6HQHE7V+Ewa
AxTrBs+C7+Ws5toDu8U9fmIEGvFV/qRn


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Zt113lgiFbPowLx0UEskX4oOcl3AzSCifuqRPqCWSKrrwMXOwTLeaE1D6X3P
dXTUo8ZwSUzH89g91qFPoGOC24APyCSEJHSh0Tje8LSCFymppkegdVh31xPJ
5LnDLUImTfIjDwlnkiLeztqwqFZZZ/8K5eWfUqa2+27BVShTfac=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
DQ9cfGeBMvLJ7DezfUnCTe/VCdH70HQvadDSAZEly9lEGQ4UpFzQ75ty5Oss
xiZJiLVBYtNecCHH15odfGmhKZwjvuVGt1nEAMJFAbXPuL6lZ5XIi9hHZlEj
uMSBBpTZ+vzklJJpkcku4Os8lzvrUjYVzARF+nsWNNmEc0HD7PA=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 25760)
`pragma protect data_block
ckcEuXUiYaxXEgtAjYevCqRdwxUN/6vFSUJqwQYfA11veuYIFsYfbwP4UxjK
LzkDQmdNoCtGPnWRkz5rlvBHowMETyRCZ0lPjCMhJYf/UN5JJfnDTmgt5WHz
SxdjkQdTj4TZnLph7CDoBwDNBfusJgfIZLjyJhKKMhsquk5LYQtsuY/HEQQG
ITJOXYjXvwX5xwoB7pAjIhKTqQm2hGUUPTF0qk418XMXfGq09gA1GfiFBpOz
uch+bjEIs4Rri/2hnrKE14kVBGmKpthXJ4Fkyczz8yaxdXfiEhIWSHbuMsVP
3YQCVL+12j+r1bIK7WwGu2UdsGJxoogOlror0Vjm+wKMg2qVGlhqzOqXZXaI
4j+lES1RuUuSwMib0D/US8QbJSy2mzEdw2XnlpGipQumuagFM9mBnu3aw07q
07pSfJkR0lfAHJH56B68SHgfpxcgH02MZRI15nUQLPCgLrkPyvPRac8lbkve
qY9m2/0NMdzR2YnU5OlWI2qIzG1AIb3edYhhidHjn5md8hUNq7eyI5NHWyxk
Y5S4MGhrAdAVMFK4JhjG4a4HIHYBibM0auRj8qw8hYHaeMpnS5Vh6ukIyrzX
mnc/RHjsWQYfJb9oZbu3S8hYNHdS7P/0yuk9/JR6W7UacjMhzazelXxnQGfi
wctumWerWn8e5Ip99j7RzbGkL6xCSG+GGvbBn8rUGN8Q5XLK8OxPVkNPj8wF
ff/5ct4g8l2J379zWhD2Uks8+p5Ti6UFrSfQw42ZlzKPRwKFL+M2wd3hHQKf
fa0eVdmLHCEEp8BlOHBbsPrRti5M0QSonr5sJJ/uGHh4wodD3AaOIQVK6zIg
LmTiH0qTE0pVGtS2fRk/JuR4ni7seI4DNW6q77p4Rp1hS9kx8MWaoH3eX/Wq
qPM2+V33O6x/DAZXkA5claBNSxNVqv7KGd4J6UhO77SwrvpPoKTPq5b3SJmn
4I5d/Ya5S3GhYjw2Z8S8RP/a0UFT9b9OHvfLleCqqyIrUZQhKI/WSFud1jET
Kso0rhDcqcvhRQhCHvKlybLj/lmbW2KfRK1upzgXl3Fk86nBz+0YgZnz5aUA
a9PBovN0ffpE1dzTdYl9mgcwK6YU8TYvWY6vo6dIu5L+6DLNGLNTdfSBIt27
SFfgjy0BDhssPfwhuWMcpWlbxUpkuxynepXNPNgZcWQ6dIgWpq5uuIK5lx4X
MvSvB70Y+JCawpUMVVuGmxRG+6EnIGwnJaf1ZETXobcmtqfs1ZzzZpFUotkI
+aezpWK9ERhs02n12EeCl0eOhAvussAwjO2etEC/y6Lq7zcRRKU9V36Bu8qv
JAwTNUClzbdmQ0BvgKX7gbQ2xBkERPHaMxi8DV1TTRYeTo32Cc+pdD9/fJb1
1uBTCHrdWVRg8EeeJTIOeB8AyXCikWsVXA0OPrfmN0+vtS5Q+U2/5LZqxt1Z
k88NlITjfcgd5pBvnrixnYIF0ky2CFWL5491aTrq1tSNQCfKfOcdlzOeaNjY
zg5YfBB6XxtegpgojQN2czClLWbLEwoZnGZeCK7I6uQjXlmEDQNamY93cN6T
+ZHGFVwDXM8AiCVDeF9C3Ab2lqNZWuaBX0tCX95XIqUJFZIXA/r24IaLie7P
ns6UxxIibcI3HxysXVhNucfs+IXIKfLLdvZaR809uuMcWrxP/Ui+qqVwiTmP
tI7z2JKbNt6N5DsppK6ZD8MkUgJDNRlv27tzorCrvQH4cq9c5TfwUr2AXxnn
/jviTaFRnHLzFizto2K9JuVA9COSSwSk6/1SAuObICElhfY/b82ZhF5xKzpF
29UJ8/gn3ckstyxoeNiGYm5huE5rdYGKc/6jgXao7qq++emNp6AEEOfZ6Jxx
n7VI4+Rx9cg1lqd3JspxbRmJnkBepPrS/6Zkk/ZU/USKYZWH7Xl9ipVHRgbA
pFCFt8Z/BAQW5cGx65Pk+Cj4Fv4Y73H0jcP1RTW6JTj/pfL8pq7Lu5Hg3KJ0
9EAwDPQZLCrkwJ6XhCuXpE58w4+VChpkZugHOntShB/AokfwpuFonRPcjRDv
Ho6WrbmV96wORn/O879Dnby8mx8afTiRCJPZw6xTgEziHVnP2gSjBWMw3179
61YSwsSy9eceXqM71g1hHuyjDv+Ws0HBlnswZSH1W+7nbxCI6/dd2Wocu4mI
2L34tvzDk5xOtr5DI/pI4ry64p22od/yT6+6f8RmK9FT9UxO038DeM04XkWZ
I05Fra+vrKOxWCooRZcBKJGXn72xCaug/4LfXQkZJzPDN2nL5bJJpYJvxXYe
9XAIhrvYjEEFNnLvCbruO3UNVTYPT3rs5VaJp+nAoyhfxVRGF++9liKbJSNn
oVuDQgoDDS4NKlMcCHHpJSpY1W3GOAT5EcogQsWaYSWYk05uCQLZReC+KRDK
fpMruR+OaZ5KqvBRZyHkGaFMRlpg+fdIGttgX7XFeBlv0APUluH2kPZUJHbs
TwkMHNxIh/IripVBL4ROwgyOwda/nn8J+0YbRNvfuLMan57ppkjKBEQPD+3Y
4Qo1+462/JC9Ty+1olaD0rG6UNZY4c6fXNt/JXZXfnXYxzONuCsbJmddlYCi
1pMNZTpppjj6poYhAgPc8Nhhvp8hJ4G+YHFwU45bzpHXZCCYqBZy0XxoGke+
UZv1bh7ibhsWNVM2kmGDjmgZx1vd0ys3+TchkMCPQXQKX0P9UIhVknsgyfZs
slkhSCNG1jrvR7spDUNKOEomyI9vXf5gxgaL0Ze7WTpI1U0HiLeAUUp2EfPX
i1vvzBdIF2V9YHaMM+BJ0YEiinN68n4ROHHw++UDaVF0r++IHy5Mx4QHaF0V
Px0U41vvEPa9UD/kkSr2ey33O16ODcuLQEwe48Dx9LRsUNNisRY4koezl/sm
xmqi7f81JTlqjFn0s0vqqGwHxOw5J0fi5j2l8qT+zJ+k0XpxI5hyAZyIuz0U
N4TFCdQ8gSIyg4B3QaKr+6aowkziU5VEdgle7wl2Xq8tlwN3IMHR1fq4Pmw8
4iz/KiiLf17ATvUY9oJpU6HIQJLhPA1AL2VYGGbslDRDYHBujrAJ5M+NCcVF
gj7/OiPlZ/pRhzbGo+W0knIi092xyIkY1LNusddWOicIDTEzGBcQPOn4jf1n
Tsadegi+g69oYvrZXfbkK+4pYBz65Xl+O+qrMjrZyx4rUJIWytFQFzojoAIZ
3n6dT69PUT2NN2F/yD3kcU7gDXGR+7wNQGhbpHEnmjNOIrbtWo8U1B+Jfzmv
L1lBV+b8ALVRmlFmFWfZAquFR8/SpdLnCiJ1pq6QRo29+J294QGwiWdrcief
a7DcqWiNwHQH8K5lNxDaaU8SCEqYUUA54GEKqEs0lsb/mz+b15W89zoo7mlm
a1f3u6/if2cLhQccKcAE4QzLsagxZ+/KG6WHng9rcjskE66+VlQN3TbE18uh
IGo+EPZXBvCsWbTO2yIz56e0xMYwuqhruJ6Oc2Nr5r+4Np4YId7T9FxBvnyQ
8MDL3gA2wn7PoJzkhx1Q4aXHFsamRbA/YS33t6d8i5pKqTEoQrp9mW4fkbbr
4xnjhMQZlLAvLQKtrBQctQf/apT4oEvODx6ewfaA9Y2uCEYO4JemGur0WS1V
grCWT7LR90rcwS2OPXAq0u5SkLxIhJFEwf4o67vz0T2/fyNEaN0wy0yB9Rbx
i9eMiRxeQP8vX5l6dfup14p6QMgug0ZGBMPfoFGc7WFZxMt2Tc3hN2ebMPQJ
I88opQt1yowyBlNNy94M0Yjz9TTZ0L9xfYKA2HwAitWXamHd27kiM0ee2I4z
gctn9V4zS5ZW/CPY9Lm9EsxIRRtwLY2wRkFBL7T6w0VyZo+h4SUPj+vyv8sz
XhqqCWxBbIWbby5EIpAuFs50vuxARLX/hpLohfSY/w9zS4293S1S35Eodr5s
scpt2Kqv8qNU0WGdUsQZ8N8Vtmt1pr5rjXhGrXpU23b7qKB0kZ8G4HSTFCSc
dTk1NAtQBjWibZI6ysEdrisyiZX15Ovy+ip46Sva7m+Ft6z4ZFN++DL2tM1i
qDILmwPuMpoWFEkXAUseNqggtUo2e+6RgN1QhMfPd0cELIXvQD/SSwTtr+Hs
/zFbKqYxyn2Vd21oL6uMzcEmEWxIS3nywxXpqVMmnh2XzbmGmmN/Js69JGLr
muWNX9ZO49tWAz6HvPifJ+SLK+rlx4P+JLBf/m4gyIcctWVGZ7jEkXez1u1S
3+MS63PtmVIYlziQ4Wq6pejFTpccQnf5domWws157fgKoykwTObE25AEdvIN
IjeEF8+YUiJB598aHKlAlx0kMr3exhD8uDyubIOpkH0XdhLtl3kOXQJDfM2R
W7qGXobFL8U0Mz5KRTfEJ7gcuY65/UsQV8byVj9mVf9x+8Jf2DVx/OxpkbbJ
rEKW4FPI9wKH8RlWwlR82mC73mKPoBOynRZWAZLF4p36246k1JO1/jMtii4y
Qljcn1CAw5MfmhVTzMHTX0v0fJmP3naNj9tqlCvWJ3CgwgikKoCE1y9gV4n6
cBG//OXJpP557Xf3a0fE0PgVcUjqzUL8zteGrLdceXG7eDVGEYkNPm423V0I
6Ek+7Ua8+oTPsa6b+01uXsboaMArxnjA2qAO2kS1oWNas/djWvHcxdwsCvx0
zN3F4LM3S4O1jqLpPx7BL8tCz4x4a8CPFbCxdaCNVchN4IbKIyaFAE7K8lJ4
XkRiHRBgTMQtQoVAwh4OG3cy5Zq7BrvFN05O/SMYyccZA48whRNNjpOgmJee
7Si6wvLOwqa5/pIEM/mBl0sesMgJbJTOhM5Xgb9OLsYW2s0NQJr0cAlbZgPK
FXwu4bzq2jZ0O3p472CC56+FcMo4WecRAzo4oMueHOBju3PJhyJ0UJIQvTjR
IeozLmrsnFzePrN6P71d8OkiuGQ1ZTTQgxAlHxqOMyVA47har5qAKjlvSJLr
+rkW6SjAoSNXUtbM+QWwg1tZ20Z7H8xMwgOiiaiiYffIwCfDXSlnC9Qau4x2
V3aB9LNtnnB9lX3lkQgEfTMvsQRgW7nADzosjzmIK9+CKN0w3NpSmDX89pJe
Sf5bZRFkzSj/wS6tfkhTti7kzYt10s0voMK1gKF0SO3PpbRJR3AaggNQDY6S
i4MXXmGb1MZ/lEUZeEx20oVg5kKOzba3OdBcUTjsuPNs0e97cDXno+SQowxV
xlRrhllVcADjtFiu76FGtytEhhBnj9x/TieQZHlSXasacbu+tQ1c12fRzGyJ
kuegOiwuUW/qf4rBE7JwD13VwpbmZs4s8tsHOTgvHGBDau6UrNpNOEj4D/lt
KYwJEhFIp4IGeTin6dm0O1Gkz5A44/jHNJK4k2RiodpHInN54lyrODSbYcnx
uJ53jpr3465MRyzfEvfuD78NjvEaJ1I7wBdBPKb6ZzfmXA25JvYgP54bPLTn
07wbnw81FbusR9B51+256iCnXB1gLSsuOhaejQGUQkcZDEhdwE1MoWe8o5Im
D7CzJRt6K6uXtL0D6jDmgQKDyQzNbplYkBTZMnlT1h09teWP/1FgAhFAYFv7
nHNW6qzfwzHQqfZrTuxMciM8pacSDRu3Wn8S3+XSIhbabWA/VKVQPDpvtdpD
Zc30Hx30GLXyNvh66GYLE1k+TCXFKcS1Zbvl/nwW+VCvAc632bqZfW3w5jgU
0+PzPEAtC4GTT6Nw9yVliA10xAGC6xWb0Da9kIGtCB/YzItRbGCNG+qO1S3/
QmyKG5LwAP0Kq5exmkY3h15kqIo0VPTP/Hssi6L911HJHc5SUYzDycxyLxU8
H2ZCjqA+EdZHqyzDXFjvJPZB2+rnl64uY1BxOw9k1SHSDn1o8K9DZA8lpCZb
S37y83hGdt6gffaydcIAQBCdkIaRGT3h1F3xHVifgWuv75a0dcvTormz+UJQ
6TYm4RkiPGA0Cx6a/aKqecM938ol5IDdX4TlgTW+xcqRHvgI334Xy63p1Ahn
48Eyf8cLvow7HGnEomtow5TSr6s5UsJIpwGkgJAlSGjP65akgSk9LSm30Ir9
KW7/vYoIAkLXEbsmcIwmeruItPuOrK0XFYUfoOtJU5pFaY2LS61pReN4r4Vo
0VDOlsdMKPdcm4fUr3MkEwyaTlQGoyLYcxudtxllUvTWS9+LC3HCC7fZ3hRd
0Z26MNIl7xZD8IGX43Ue5NIVv8A+wFbLsuI5ELz6K/swtsFP/Xoi54eVQZ4w
2bO9JBw2afwU0X4vc3mujqfMrY4lwYRcLowOze/0n4arjnslyhHAgOvQqRVz
/Riqvb8y7355+dxOznIWb/CMVwuunRXfSyGMSEl5Abnoe+1B1THEcLSSqUCY
31Bqg86bEnZqU3f5MqzzIwh7pV4Bbh3mw7n4MkLT9KC7ZssZlqLmrqkfOBJO
j+OZ1s1kkaei1zXJlxfBzSOLa0gLHt+s007PFRdMtW6yqJOhcngO7IVkWQZM
izPVDuV43cbg92G74sZEEA+OmEhgw7yUCQh7nhkuCrtH4Ks12+kZ/KiqchAn
znTIbWq08UVVv3NY2veRXPZXSrMI6OLxjCGWD6vB2iWmDvY/Atft/NHZyeHC
Ybws7BjXd5llx9DErUN7TwwAqqHfhS012+UvZSMrWQnbtMxPmFTHmGtdNWzN
Iev5RTa9T+R2Dl+U1hdZZINJE/EsNbtsshhRBBckUQ13eLnfW5/fnJM1P8jq
/p051Gdb9Pbprkphy9RmWWc2Aa0j12ZkVm5rD2+CbLoUtC8+Kzc5HpnmMUJ3
BA0hdeiu/H1AXPDEfSJiZ84CHVipcbJFNz6E2MGZICeZVQ53+AR5giFex+pC
E+yxmHurtawi9YRNxK4gmdDKYLtORqUTOjy1kv9M3pWl5pixQJpvudz+8QvM
SzF4PXJ646MwB3N2FCro0OxOC3B/IMiZpn6yGty5DYcKzF7w4+tL+Nln8TMz
2P+bf9/cNXWJRH8t/+xXS/nCpYHh+ZV+7QGphdMCTRp0WGouG6m5q/3zxIvY
moNPBJznLQltOCxkaZ63GDqas2kzLgUE/jHISiGWl4++M5sOULw884/K8rKG
VSadOMx1j1EmsBYO4pCWHPaieo752JsVhx2wHYE6p49wtFkHK1HGDesUnO67
RuznDPD0T49AYA1jcFFpdefBCZNLRwQRMIuTV6eUb4AYUKJj+xGbtr/npo8q
hDbl2Awdbu9sGKNbwAErGjaSaeagVdCMhUEDOw1113SdZvxnyas0wZ/FGx0B
XLZtnDPvALEDkMAgWVutCeB+ug/md6Od+8ToPmbdFvg635H/QiKHxJfUtQNe
jmXOZvrmrYKbujDbriYAQHkK8ZytMfOu7eg+XNaWERJ97wQbsdqbmFY7ByHN
+N5UggRa8nC0pPdQzuFDN2EZjzjp+DGxpvSAE4R+Ebhl16VNnCizz7ooD4S2
JnS2AQGYtx4EP4o0N904ZbDLm/J89tn0ubc/d9bqXJhSEt3K7jnYZ8ni7tR1
Q6Mcl1zz3qARUJdXVaa+JWjZMi4PWISXyDPiYRFbZ3C8nnogFSuoLFdhfi4q
KmaMJHPG4pNJN4YY6cToIpUnOVA+ZkdqWg6tJmmrCDQvAIgVCwTRUzAVQgwC
G6ZEkwmLTV82k+rFvgi/sZn+vzwWV0aZQHyIee/Gr7q/AMHP7EPH5G0o+gtL
4sxrqqOgYu5mi1gXnZm+UzRUzGHf1KsGf2hrU5iL5bafzvXijmyHhm3VXHmZ
n3LdkoCsOfKDCYTeeGnpKQpxyTj14ykvC/EZbDdAUNKqswEMiA4lZ2PbC22f
2VlQV7OsQpVNntB4EVttQTyROK0k1Q7ZetTIya57bmQWXgCYaHFitisvbtBz
xFtiN0tCVtgJA7EMmBVI3N9NXOj+XjJltazBZ8OzbXKHi6g/ZQs+jV1MFlCM
UQXj1llBAjjVqVqhxeC0Z0gJ5fqQrz8JQRDyF+3VE39GAHcfbsV60bQzNnfH
5Z6tKACEucsBoJZNelxepKOFDkakOkfn71sVso+iBwmPfBwzzSI5BiMKGHN6
OM5SUd0dmb0Ek5Q9EaYxxLfmLJpJxnJ7mv4Vdzu2gQFPTAytDrjaVvJJw0PO
E8dhl3xIJ7E3cPotjpwFmSYJCaCt7Qzfh60O90TqQ661QHkwioji+BVB61Ko
+GssP65BwBXwNHItw8vm/OzrlMNO9mY5XOCk+F8eOjSAcENXbKGg6+GBMQkQ
I/GqFm8EbindEwYdpXxAkgi7o/oHSQ3Bg+x4XZKkjiINjJFFSCW1Xhw2R5Pb
J7TaBdhjaVYR1yVrMcTMT8f4aK4gEa0AmKyi/iKdUyCsp408D2h+s6E7oXbD
ziycmM/V1ikB3FgjuH5touC6pWoQxwv2ed7gt9om0f84hECcCTjGyQhRgmW6
Gw1E4MSpiGXVig8De3pfzpiue8a0lpXdoMtypsqiTE3mUw+phkk/H/dnv00I
5t+cUmePwUDhc4Wt/HlSABrVTuZKg2v0FlRPJZ4ygFvrf0eaQYmFGugNCNhN
SFnOKT3YfkHX24Oh3Fbmwg7pYpKOfncFIyGbsipng2Hs7lEtkCP9MbiYmajZ
79GuU+lTr8wiOXxR256Gdk4tBdgfo0lvCxQCi85IXYpT1QhTvZjCaDRk1nVy
K5eiUQIQnDFWULUqrRGkrfGkDceEeK961860/51yRxigyVVzvkOztSS+52k8
STYV62caVnU0NlxuA3L7McaEN15kSqR7skbxEz+J1wJTCEZsiozmNlsnegQq
S5Hs0XzCObd5uMz3SMIMe/mssdCisrQCV66mlpCMPV4E/3wTllgvENVEd3Qj
ypEHiw6yOWHrFtjfsc5DUA0RAzOqWyGxmhEa3Q0hYQU+mOSucz2NGzwF28fy
jTSbaNqE1D9/cBrMl7bomZOkptc1T6bf85Fo1iCIz80x9HFDIax4O9EPc67T
0FMefvLrvNhEHkU2qQ+mF/ABhxu4O77Cvm51Xqiwt2au4d1wywjS6+949ocQ
T+sO+NfqKlTI9DMWtNNfki1kpML7vVS5Z0RclqGl1Ae43AMDzds0SvDGK3Af
dpGJDRJv/bIIDfuRnYwG2BGDrA2RNomFTsksnmOvGsuWt+3yktVQqoyDTAyS
GzIy4BfOmOFRb07k1mnXvEPqOvevof1oKvC7zCWQN3vZxyujlah0vFmpEOse
s+Y1d0cnId59bZvCizAZOit3J5c2AIL5VBEgewavUmcRqHkLswjpYusDL2Qn
OxYJ4XbtIciITQBFy0StmV5YMiDERql4JtD1Azp1ZfCzLhTu0qAhtU9aWMhK
UHQQZ1s2ppLU2Tgkwe8HSo8a8JX/DOfAHhT1Lt1cybcsymqRBL5m+lSZguAd
1lnildAYYNkFSV67yyd4g5tiE6LQ4L8Enimsjw3oiSdBpz1s7DntA1acml6c
IS2PokKVJzjZRbR741rLws9lfkS1j0/SgZOirGtUA2dDIQaw2Pj1JyxEills
qUPeSg14M+jQotqjkf3IbyNhqNkjuQGb9xwYVWwWMUPKpQOu1fheWXVIF0n9
53IUz04xJCllhD6eyu8JlAuU3XL308RAyRwHrm8aY+r/osNsqH66LsemuUHD
SHE9khvLg2Z8ekPLTWw7R7blgQggRlkclVDyLX9rhk3h1zlXQNOGXQmskgBj
UgAwNXev+kR5EF6l0S8gXUfLrGethURF4J1JkpXfpGTrk/WnpsBXrwv2kC0U
d51OgMCJm8xPL+lUD3CT85ngfd6W7+IeIEdJshZgtN0HtJhDSIe/wcebFgEA
y9+u6ZFZGCAQXSHS87NwIrO21oXaInheV9Ucl6k0y0qCpm7x57Kz2RvA2n9x
qHQBHmaXtjTVC/WiCCjVqr4bSK1XE61FUvOpfrJ1tEcVEos4y3c8CxZI7AH0
koJM3IQIylI942FzExD68mpKM7URBeEA/1+n0dZmo1RCLJanjDb47w508G3Z
22vuoaNrSnXnPMkApVn8esJDRTzM+fw9LtIAGDIQgsq4J41Upi+6tvadyhSO
mPhVkGIbZ50MXE2O1E7oUojsxpXy1kD7SRlggeVBgi1I4Ut3hR3ne/SW4P6I
c/p6wEESHS8I9pPrdmrfGBfnVRtU753h9KBTnjCZz4CUd2fp+jweJ9uXGLdl
hnIjyHJQt8SKpS5/aicpsqD+AMWjfHeTJVD5c4feqRqiRqppoOSo/aEXrlad
RuaJ4DwOfYYxx0VQgE4lx1tqH5Uidi01e3BQSZtFwH7RV0tDwzff8VuNU2Ti
huBkyje9dtiJj1ECV7txpBfvB9oh38EI/8oizr8wK46tXKzen8J6HrY2m28j
s1LYI1S9MnZcZmZLnRzp03BSlwNeWLNxqMXTWRb1+15/j5pWsK6P2iVbtn36
YilOgPhBZ5RCpPq8KRTB/vDmLsQt1SWRtULmaga2+hQzeO5aMBAnNe9dzDPU
QEghDpQY56rh74QEv4W1GfcR1ny6I6zgdn1L2A6GtwDhAJ2rBB8y80v9K1Lc
+3cXIWygNWp4bjRLJG+mVYvC+SQCN+e3oVf7si5LtR8SPA+PxFRZ1KYbQm8v
zvUSXlw/i8huna4RYcQxb52GMiQOXa3Ohi+jam+T3m9w35b7grQCRPtyzfme
zr3UKnVtcbxTz8igvSG+DDZEsDU+aq12AAaKb+8xJzKUXT6WH9dfV1Rx+ycP
g9gm0/4TJOLPdQutISuttUNBBs/3zbh1wLtOGjG/0Uqf3O1uFPeWS0yvZger
6T53G7DZO1GAqe+WkWK1K4CAxS6c0dkDBOZvvNRe9OvPQBGAf2VaKp6kgv+P
pxiH+K+S4rw/DSmOG408bL/Mdc00F4zv/mmSVUsKYU/duHtfcjAJWhaazlRb
oAok0W7JcDpCvVCLoKZgfRfns1IVYzgLf0r304eW4R6HvbJsQAZP+NWXfLF2
T1epDu9ufcNWqEVbB673xicWBKj4gJn095WxHcvOVmlystWSOFJTNWI0gDUU
ZfK7MAR0ZMEMwj9O5zjhVMg6th8pbDPpJ+ZPETchk4ME5KkNQWL4pl9MDsji
DBlL2oGZB6BRpRrXnMTjqNbh2L1pUxV0yQ/FGZar9r71ahGqxF9qWJGEu06j
Dc68Kx1fz0RdNIBO74OhDSt82PbwGpNAhUNV+oUUlmPJAwvz1WTw/6cHHIs2
4B9IUxi+TNiC/vtNX3CTAQGWEgn6xsxB6Nqfy3j+U6Qe3qYwSD23DBa7ZCFo
CMXSGe91C1abRaNtvgITH9T+c89Ajqnt7Zi3ct5HfQdr7Lu9awh2pTQe21ik
q3ACUm5s9GY+zgaWphhShTNKk0OPs6OMpRLaQ2i7m9wgxPccgZnWUh61KWKW
gnjiXb3ywLufPIQVovNaoD+SFOC8nWVkfAVMVYwSPX5H2cKmYgOzmstjCJlm
XAIOkTe6OSaIfHa7b151XZuXLAuBqT/yXpt4HkFeAVFMs0MyYpfOQy5FsZvW
Zww9ITQqTlpI6/qsasVrNLLvN2myN/nLvqU16oocUfrguHOdCRCno1B1uHsP
+CQfsP2MVQqZQiWcadPkaLGG01CVyx/Z13kTmFDdKma0u5t8qA/8A8kQY9TW
E1c2sd9TmEJCR7aHTkTB4FNenRX6939kMApLwBKWi61nOQ2uiVt8S1ikObDY
dJtadE+JYvYQaPzgwmjl0uK6rTZIHR6Uqz6d9zYddaoLKVhWw8EtsVXI9Agw
c5VCpOtx1otD4TQJXowkE/XHLV4u8lwJzDdLi8MTq6Xn5K+sQa0ATajh+QSm
vgpQiyI8JHVK9tE6PPrSA6PQrDo1I+LpOOIj7Ea8kCznLs9VJ4NOH2a9rFQf
6rRvigVJ2sFh6aL0d6AkM242fpWWHcenNPCXOewAjVUAiwQ4XWJiy8Tk6A8u
TFY7Ju0SjKxYJlrUhbWIC/63KYN/ISRN5EukeyUNY5eu7M9Gigq271rr90C5
k8PQcsy9mmaU6T3UYkO+QtUfQMJCCQw6wI/5lJq0zbxWTvYYI3Z2q9jspEIl
qo++0kenqabM4m0A1QWqc3tNNO36B1T1fmrKEOImm3x470NE6VlDvxYQMS/R
914oJDSzKzzCVKswEKZiZNMU9atsMcuyPKGeofHTgiCLqUd5NFuWjGogbx6L
f7ysWIerNgAm6Es1zdT4S1JvxMhuP49NtW6k20gksZ+8Jf1KQ/RzLbpoaC9M
RDDMPJZWzVZ7A2ohO8O0/kv/LRQN+GaLAKZs3UyTNbTeFCx13MkYWOpHLgwt
tslHUqJRmi927IurEutTBVa8DJwmocVbJ7p8SU1Ts9J16tj96toCnio6fhRK
WWeRiD5i8kyQneLLmh3dnU17zWeitKH9Y3Xn9P4k/Gmms4R1D+el58rmnhOb
0KqlKoMXSILBwvvU0tciXzUkt81NWWdehoA1NHqqH0/txe2Lzd+ltyWIrWV5
TwM07woqYsnUglBzKQgzBPuvT6MKZw0+HklLtYkueH5gXLIMfFePACaHn2c5
PMzuNFt52g+SHV+8EKOWtTIUOHWItrHEZihVN/uq7NbKSCe2zGhp6i2Emquh
NplwaaMf8KiritsV1ZI8+yi/+RCMkQePq5TPi1n9epLZ5PK9sAywInknCUXk
uim6GHY3CghKzhPWRksokUEwkR3tSPHeHTcz7IMJvo7lMoixBHC3NEKqgZJm
ECB/YTDlzLnQ0/bFJAeeltD3/9WqpWBoyYySh6qqewYZRxYBFaNBOjsxseKF
vCLlLMBfk4qUOaob7p6tegdH1HL6r6Ctkx2Pob9jfQYQm0dcj3KWTLM6I87d
qSEkxbvlAWulLidp8rzehXxQPA9wMVNS4lk1oOcz0G1cFUkSsA8orjpeU0nf
OX97r8wSLL5SNypoTq4j2HXui7hbJPYAo5+RMqPPJa7m/VuvMQPkhEunpXkJ
0Y/Ki3DCro01dZQUag7ft869wO6es7XPMMr/twyU1w2UDcQlla2c8QVtn+Dx
RLPQWErz1tbYA0t/zNKdEGXoxWRPTr8lRMKDiMR/ECJZLOYoMccn9mWf1VPe
zXdCP++c+v8ahFq3VioWqq4WCplJprnGqbmIL6lcCbXbGruZj/IJdEmeSOzu
VbeZjN1jOAhOFU5Nohzyn2hNvg2i5dorn+Rm1uKfCqlLHrsdt9XOdTxDyWP/
4/T3olwsGB0jZGWDdAlRpgxH/VVX1NgOyRm2+dyE3NytqduedKTbXNdNUqJ2
sib9S6ByyhCPbP8H70aI5Q8mytXBCvbO1rrqh6oruWJ6GdKygfLycHA/CmAf
94WKGP9qkWLV2nFKO2/S+ZXf1e1QA7CjVlIHZ3zjAAG47WUV8u9N/ScCivop
opUj1LZ3d2K8JuHbL4L6o8LiN4+oNCaADikk8Ia9P4ss9Z/0GOiy3y84SHC+
Turw31QskO86JH2kRtOiMidVzlPyqI7ewYZ31yPbjXComdLp8QxwUdHLevs6
KDo5Ciw+cMbGJVO2Spif1kZIdQ7MZQs4LqInW1YkrJwEHxP/BWHEjMbXrEjs
jioOJ2+reH9dafznUarBS95O13KhItfApyzEMJ3nE2WQh3W2N+se0EMv4XoX
AGzbTQ4t2wpT72EniRjFe8CmrqjeSBxVGEZqH8lYOjyd4nM50l2gXs9RZYx3
hEOrJiyupn9iV7jvBsvWIvCvywYQx3yFHpwRFD1bRW9qbfvxIK+AJDe5Cl02
d96Ut9xULrc3etMyKH2A31gOioug2JyvyXRPildqJEkVkH9BUv7zJKmOY5Ye
ewijXiB3aIAdmYclUzq/+uOyOLlT6ssASUdYnVxT6U3tAz/V4olW9qCLuwhV
rckibpkMMxCiaB+YxOynH+Yi3GmawgxuK6aYhF+mmNTumCQwN5NdD6x723LA
GRFggyhHGVZSyINlQtYuR8h31CtiM1ClEhPit8+C1NPJf3tV38jdY1P1O0AX
yujd9mhTltyqpIBB1urd7NR/l/7Ed+1t596xR1qNC5Vej01orT1MGSTWJa80
khUMhPH09wweQHKWdI7Mmffoyi30PDZU5qtrIZ1wXMqW62M23Ssw8HThsA4G
S8y+HbwzJN9AewKV+TJY6v2mW+ZtBtAcyTQWKboG+AiM7jK5XOVaSEhoqh0y
ja0h1fuooqczb4qJvmqDu1HNhNsTfHzvkATU21P4LaM4T04g/iwr/+TynHpu
GuRAKp2qOTHWId0l5xnj69DQpxODO5RoR++GqiPnYT/NDrs8ZjxBo/V/8T96
vR5KK9KsUt9muMZ4iJCu5NGh5ony4DZQ+DKw8w8euNdJgTYpWt/MhDeamX9S
taJ2iHlaPFWivzgGB4+6pfulFGRGZqE7+gdcjVk0vSCYmzpyznBUtysOKhxf
P1LFfiO1K+8mnMzJkR5Xs/WJVuQd9v1StGqaJrJz0kOrk03Lx61rElbLZexs
TSYGEaHSENGGbDwH/mQHylnEiiwu/IqCd/v27fky2xC0kIssNpW2di+NSetB
w+wP+lQMXj3y8V7g5Em3WH9zDnh+X0vqKAMABhAGgLfRkhGnX0GvJTTOTrgw
Qennp4+PmctROPtld62anqXwzAalroLnfFIky7y+0qRuqn5G0ozUDjAYubFr
tLYLRVxzjGxjB9y9SyhO/PJ9t23sZAKSmfw+oOWUZGHvNnigZovRBcXa7typ
tDxRGin8KoUcgba4VLD17zQKA9fPD4nitrTzjZ2hvJyBoQwGy3kU4tE/Ox5f
KxucZfsmoSN4Eiw9aDoLM1vEG5+okDpqsBpeJl+tL2hQpfP8s0hy2uFyVZxM
vQoe4ThX4lTdAIMxE67ALOuxVkf/1ilc/9sI11B5pl/IDkFiJp+LuV5C1mTi
HhLNPZ/Y2XFr+KSCFwI9Ty3XkOevcaeUfDTSkCCdRwPiGFF0Fc2kwXBMqstZ
mvTm85yGEYsOz9EzL6NP3ZvlKQwQLwHO18t/k0nLXcGLaeOT/hzxHnZL5gnM
VJc/hiFnJ20/cNWo8ZeTUG9hrbkGDlfe7J+7ZCG4g4Ot1NSFAjbrZNgbP0ud
HkitPL61EpzOE5QKR4da25xcXKLSPCz6zgYEG6DFj2NWOEpvViSFxf7CcPjC
BUymgXO3OByqQDorPrzKp5lOdEIMg0QXR/s4yuvHAvF7iKVppd2TMzp9brfu
0Ql4lGYc7AjCS2nZ+XTW4vh0g8Oy+pd0oQwhNYGsdNrv1wrROvsM4ts9xL/Q
pVYQ/V+D5Axk972LSAnqKTIWOQsRDtyu0GtTwuQ81EcPW9+dJDttmlK5EYK3
Jg1Yj1pstqmdhpU8BKvChe/MAvCMVxwpVezQbucWaIisQ0gnkgGdegBKsxBA
xCZp47cziAdBqa4pqxipThET+qQPYHTocNsgj6BKZ3Oao6UWzZch0ubdSAX5
BdL3RIAwMhRMW2aClvrGcW5Qfrze0qBr4wSPaispL7tu+fy+heKiREqdoxhh
IPuGEyLe6pyBrbMMb/1I3ZHy6BEwu+8QCoKCeAReMYT2hV8qFBNlgJHCw3Qb
jyMWVNVqUf8tcOkRIqf2dVkjEEJBO8UvnfNpJyVEnGlv/Du4Lp05C2XasqcU
z/bHCkcuwIDb4zqk89vCGeWOn6uczfls4112MgHckDaj29yR8XhZgOksjVCP
xbFNoeAFRwf9p+0T4w3YRJd5rznriWWNhcQ0uDpIKLm6PiJ0XUZtTWhpiRMB
6xFQQ0ecvvo0dFzxqMCmn+kGSfecGWMHFCtu0kxELobskOgtr7K+0g6uxM8Z
4w807DQwAvcheM6QlQOlYGgs56r3C3RHPpO8IlGq853Ihfc9hC41qpgasCX7
UctbsK2noUt8QCzTIv11oMhVBfSV6J/1BAUBkCRA56ljqzFYjJL+n9Fr02H0
B1c6SJ/MD5opyjyrHS0bgvnCg/RJA1wwCA5seoiEid1HCCdRFwB0gULz5Yhu
JW/GbFhHJCGmHSiHN49SswrG1K/sKNmE1dq51WLgsAvcQdYmLx0/j7kKtxzT
Mvr/gTFPtHtecT3XCOBhKiN7AxsorGotVZ/GaRikhoanW8H37Lx4AV7ESyQ8
oXorEh1mGy6mWGKwsCSPp//HXof6mkUjQfakpLe3PiHDXN4FpmHc5OFc4gon
1ylk6WbOXgqJbveST1FWHV8cdF3F2tchOtLqXaQ2dD9InbiKdSpsugQwKQgA
aQjMwLHW1Nz244GHookMbgYP+hkUvcnmeqA1EKD9NvIfyDe7b7ejrLwBRXaG
1DIpvD3spZYEwqAU9EXIgyvxYspI8/wsqfhcdDzgo6Vk+jXC4crfbCpibEsu
qN+JMN9Bydbdhyl1NjwYDrIVQXNxHen+lziqLgmFjoydOpC/VamC6a06dIj+
jR8XKPZCVG4fUIgLr0VIi4ZC5hAppYYqxLX8nRzeZnGXcbHy/GGlAgQFnxj4
HaEcnuVSr6BC39OHN7iurS6kz9eLRmBcI5uBFnTSzmRluBfqBs8oavzDjy6s
CBx7NV+B9vV8hB8XECMoz+Z+dQ7vibBdRR5vQbfmhJg2cgywHzhJe+tu1xQR
unubpX504hxskLK9VxKzyC0QE6zp5hsNvTBUcooh7I4bHywB+1kbubUDY15V
YWxeeZdJxnbwVqh9c0pUNIlYh67ZNLDE63AHPCjhrGQmwbT0W6dTw1dgtk/0
uagrUJTO9uOfkw3Ps0JSz9S+XF4AWhaRe7iZhIIF3qOboQIxqIADstGyM+Qd
xQvF98ceOhRmFCjpcUOJEwOHDnhbuV1NUUz2RtDPY6U7YTUyRkhG5LGd7dDN
8Y1Jz4409aRd5ybMh+bE4k5KuXgVkD7FMmM+O9X8G/QeWbv+d9a7O9A9k5rD
QotpcftYkpiIbP+ohS6/96IYOClRuLqeX183qPqk/IJkRveUQ/bsDl2OW+wA
srLEJQSGP3mIGKIwwFmGTA+VPOxo9ZC10Gqb737+UQj7ucbFILFQQOhzrerr
MqSMaOjb47Tylrfspwj+ijAbjhs2PDIAQ96qBxu/q0cJUr90qT4Z5qn7i9mr
xUhC46A58fFcEasKbmXFUJrx63KLL0fMEeEZF2rwtra7IGf7aCjvlC6H8yuS
dksHlM3hQzAzroWYbo16htX0QdQ9t1TxBZVmeKkEmhmCL0r1IrBAIzsHihkw
fZiFektuvYCj3D6ShQFHctoykMuq4AXKTlZrIKTJGbuQ81pJxG9YB8iqYPh5
huitF2COzb1UKd3zVIl317wDIJt8tHpIefOKMVtyE8CjaWdJgPli75G1gKmy
UXNm288yu6SrZ+QN3kAgjnRqIHhhuiJjcZnPRorpHpgUNkAJerHiIvJcE4WZ
zdba4iyrPxXewic+nH2L1GNFVc4PB1JXbXX07MMfhWUsQhqeJAVg6Iu6dlLh
r/VFgF/taIfaSVMVLGYKkbc6sseqOnUuIQYr1w0uO3TdfEnZNlspja9q07f8
A79WMVrNmlqAZ+pvy7u5fdTkoFGeqG9lfShjDbyRS/mc0SxW3Jobv83bKbw1
OSEgXyQcjQIxq+CHe+wLhDXb5n+bXVU3qF/4leojNE5lAq9uMta2QX2W/tWH
1ORjO1b9qVQRBRh+xNzgP8GHQ+nzfFNgniuxV6dpAwu6eIRAGOlEQfdtXDXn
LC5LK5uhaxY+yHhIFBnf6uvoAM4n0+6ADiMFzPM9JN+1vv5vcUKT3g6VQCoR
oh1OoPTFnkPmtDnPhEMzTSknyyvExB7MbB+Ny0f5P4sO2wVneUVqGiLECxp9
+v9IH+y+85VU3/RHgJmaSyoq0SrHU5esKxWr42kGaWG5G5ggwf/BqBBYdx0p
GnQvYYQjS+qxOT8CTZGwFlChuRvNscXACtAX4bMQYT1vcjdvZXGNuerJ3aQZ
hPodyi2BLLTlBvwq+LbC98MG67XOvVvomKdYbd5DkpxPJM4TCQoN4xNylH59
nTLNRL0BNy4wiJTrr1y49bG0xoWT7xjNLDUCV5JGWYljSBbs2Bygga8WdigV
xx+ofe09ppCbyE7gSv5iEBcUI27YnjB/vuPMk8OQ2lRwH5GJ8dBJh/HOL7B8
o0rvRErFemU9QEJpNQ73zGxbPZK6cchgjkCN8Ho7v/jQgx8PRFhQ53ZsV8cv
mvaUI45yTwnHA9TOZkTRhhHLDYv72s+WsjO2QHDqQZT7iZRL07zXD/u4P65Z
d4ycyxZMtcnbCutoEToxzseTKUzBkba0hTga1+6XpQLnCvClL9yW5ERfya3f
uRG/1ePTKrHtq1bA1BV5KwLB2ok5IPKYyJ9Ck57ftsSsoskSf34GaBVafaIS
j36vf5Kboe3DFtcvkNapTu6Vgc+dPCv52iFyFaVM6eM7jI9xDXNnrQfRjHPl
mcMMcAUUJ34Ltf0ZZ9tvLflwR1k80leEIL1yxU/4Q6pXRrGkaf0hV37QpCXM
kyU82MlRKyifXcSlqtj8uWyRo1SGntb2+fO+hDnLptdhJ6qkH3zmyoq7yGSq
v8kX7V+uwpPqX070UEV1s71QYsAuOdiNWZ/YLNTlTmWu8nuknHE7ruO6f+QW
wB/gCDIVQBSD8HQKLowPA1lQbS7dVulm9mEDef4Z0tLP8Z8LnaHetzL8hwnM
dLOypNlmGwO8xvM8SMc/ECeFPpjpzYUjh0Q938/ZWL7G1WRdplv4MjolBGcw
pZPWHLNstHPZgiqaHweAYngsnPbkLprgIJ5Q28+tS2NMfa4D/u7oRZ2/nmFc
ZD68pKUcK4NZOhh3oQU0GMug19aoLpYoTYJQzDmTqLIDtvzDElqbo7O1o8+j
W7xsvfD0+YJ2y/YhKPv9lXIB+eYyLlXm0BcujUo6C6pqj64DtFr2ApHLZejy
wv3IVEPDxfQdpJ1MRNiX/LJ41iYA9YfH61McIsiPxQE/B75/VjrLQ0XddvIy
NV9fRy3bZ2YFaO+XlSadPzyvE/yx81TFsUx7u0HHorbaJ9RVdFOJoN/+Dc9j
QYKaRn44HY/ZM0FGcQ2J+J77C6aDjsMJVqFPMeuxT18rywga5V0ZJZJb18+Q
hu4FPTogWNJhykGc5XigajLgK6ce7cYYJhwfA9NH51JR/tDaZmNrrw8PdqVg
C+LOm1jLNJIsqFjoDz/bjt7pqaswUVlBrere7rRAyia+cTtwYiS86v36ONQ9
Z5vMIKYOYXNifl89b3w91RhNjVe+Kx5x/k1QwjNxCDcis6WSvNslAu3+V1Ux
81KCvAO2/qIlwNFIzLInVvkYzJthpGv15n5XPh9s6fV6yjtRuy9dLAzS9L6f
DNLV8N9OCIsfETxzC+lMBIEgd+ef97LmKmd0FqJ8DAjhCGeA5Gwtewm5hEkD
6VoAnsgwp95V3zZ6qJrx0IUIQqX8KDDamJvK5ojS6ss7AYx1o4KqR4DiZzjd
dT7IUWoXl2s69GinMsSfMn82lpI2Ab+Jrb2NebMTFzvbsU8P1iCkp9TM1TWl
m2uLc6mH/GBtHxdVHordTtL7IQgBgI8+bwL9ShJ/GYyp+ax+qaTgxGyCFvpM
HZLEsVspHTuJknQbURBXFMUc/sNOcp3oYpqW1YLfxWss+rE+CwEGK38+N8+A
CM857VaLX0fASA6+w89ak0lbqjgRccUDWyaqdaMoWnRWFhiwcGoNqEdAtQYK
4L44v6xABCw7+Jy5hY0BS6tEtOTzTeh5jJXAdWWOitxEfCNJ1zVrwUPqJdHn
kD2pBXi2TsYgcCGpyVKSF9VR8b55ax8Njy05fMHAd2CIpXeNCixsfkpNsnOV
Ilpqr5kuCmpOl/gCJJqgiGyTnfbI3HHtpdSB907r+/BVJy0/EwX+Zqm1GhvS
lGewP7kAbEdLqIzMgR8O7GU/7EVDlUAdjWzRm9hLfsI9nERo+f84pq+ADWrR
hHfpj5TKSdMhJmRisS8u/6ZWVDxOZRT37U3/nMXSYFolclVgZerYVM6WAx1Y
fJgaw81FrIYPdKEjeG4BtNs+DzKh7uImWeANjaxubrDJF6CRu+jG5RLLswYf
sFGYa7o5t/GUHaR5BnR1vvNWx4dbQgirxpM1MnAurfup/kKrq9kEbqZN5/+G
Q/Ergb+RMJnr1FA8kjleAHRdEXz9MNkmHBCPtMyAGh7SyGEeIE+mpgmwHgnJ
E32WPjaPRz0LtFAJHAree7FXnGr+d0PYtbqM0WqxYVbZpzoI5vW76QiRicnd
oIm+573sejqLj9DDPOghHeooZ8iFfwuWkqNMe6PPCMt7MQBQ2Vnmz4jVCBh4
wHJ5tiY/GpSATXtAuWg5r5aQBE+jKbq+y3Xtjnn4HniS2oPzNhoq/mWZHyL0
C4xaV5EfeQSlW9ZMsulMwUXuznNH5qusKpKtH0EuP6c3yjqzB+MIbs1LghoK
SOoGSB+x7aMx0+K6fEQR/XkU2McC1zv5WT/fSFZXacdypC4gx4xkW0CHjL+h
5pSnAUFy383aj0jjacC5azeUXcfMVf5r6k2wL/N69sGgSrqAnmbeRz6P+NCm
u9QMHVzy7aJSVQxaENDgmcgv84+U4MXFIxMtcYVvNwNk3xH+ZnW+9ZiR+S7G
eRrwqaUMVdpYWEbaZW/I1f+Rmstccw8NP0Sx157NdOJKTNpJINS4zhMrusGe
CCX62gqtZi9NyuB1YO0DViW5sqjmAxrLP5HJTJN4jJ7HAoALfc8E0eTF/tVE
3Me+PWj3yEiByutQEq9XmaAwyzPXg8LsHKVbL7ntzhBD+/kX939Meuuj59I0
IbqG40HXMtQ14ZEPNnBJ1f34mcPYqhxSeWkX/yGd7f5KJCthj7wD1jzLPdHQ
MKl8WGt2mnVRyzUsUATcXZHLhoacf6aig0wxkAtGIjXHT7iQwwmvuv2zcaO0
1Km3qX4dccLBdw1tAjDDh6l4rJD4wkg8rWDUG31jo5n4yHmfekL2w46Y7Hy0
P1PEPqRaq3AwNUCbbEoQTWUsxmDL7V1HKmHD/G9M/ouqrgK6g1KhGeQe48q7
oLWlKJj/DxhoKcqbSbbULrJLg+Hnbg/FEv1S0SdVYH717PYHUXslkb3JiSjO
fG0h9Iuzs8ltQPgHWBthRFmK+kDTq6jkB0iGL9KfY07sc5eLeIXOpEXmSTeL
xu0X0nWgpRQmptg+xwuxu1uhr0xh9S2Loqd7cEjLxqnpDvN94hXxAa0mXeY1
JxMjknBD5j5lUupvSjFEKgBm1jQGGcf6NcdGviIJCSui9KrZ7zT8EZNlKnvN
iY6DK20KBVI6tKdBD/h7ZISiLTh1ACRG8wqw75QpK2jeLpqOlmA4HrHdTvxz
0/x6z3RnM9xd5vfG6M/8FIrHXU7FBlZHlugTiegVJc0ieFkNXn/kIeUl9viP
qwwjFYZ1/ldhHCCrt+IBBxnz3pY9VlspoMlX7u3lpgnSQsayG3D72Oaf1Efj
lJmJPXwBO5DvK+jtAkoSMdVEHauKTiJy+56xFBIBNawnTw6glFyqda930Q5A
xIkwR7g4sQKs3f+O4x4l1xucEqKaVblI+54e+veCvTmvu2pGZ9SVWTsoPOoQ
V4nZa8iLQywA0DafbtX4aprcZeK+W+J5JCvN860OLRmFjlfO/b2lDI/9P8IN
BoEsN/ySe1df6+4VILdSY3UBVjTvcVJ0sq/12s1/hjx0qknoTSj5MLLga6+n
/xuTlwwJ8tuw3W8AHny/NsBb2vTYcZ5JIbetL4w1kKIUd4CDIv7tEW6uPNg+
+gR06qUTXMauKiS/5TgsEkF5E2BCQlwAhrMYgovbF/NpONWs7l8WRVU6ZixS
FRZmGRBGUn52GluQ8f7AwMO2z+p7Gn6cHK3lKECCucyRrrzSfde91IXGQkUU
OSmaN9aOSX+rBP7iM9nQgmrOfwocuvC4tVADl25klRTTqv0juq2i/rKlfQtq
Xg4n+pM0aL+JMycWJwjMbzyrmS0JgyDY3tHMDG/QOH7jsXCMmhWBIhvrITmA
GDPoneR71g4ZgefG9ponNInngmRBSrESl/0iMuIarS3DyFghclLX5FPrVeB/
wgLvH9uMMXSKIhNGUjKM76xLnfdijczNAgc5ZO64Rrra2P/02Iir25XsPrc8
VAcQa/TkHgSvc1mRVzfLcWtZiizmdOpq6nuHeJ4NHzZhvLyRTdQoC/ZbsDxy
FE4ipSFEb/m2bSlwrLxZ+U/DeDPZxxV24cMxblp2eEB4CxNNC1Lb5iYK/8/Z
6YqEunTZ8wWr8zLEO8DH+8qaVPDJBUip9qQrO/n5jIyv9KwfVqNd0xGYXrvV
0bp40WZ26pHGxArP5XE3IxwjxTBB/ObiawMsuMIF2F8XetcNHx/zC4fMC03z
rKwWg9xrbTZvqakUhoiR+X+ldSaDllXZtXkNWOTUBphCy65lPU2/LCM736jP
rRGd3l/x6EBihhQGtoinKCQKA3YcVcKeUgVPmEnK7GOhuPLGQDPsnqR9q5CN
zRRmDfHCglfA+g8FFHH8V35hsVh9Sd1Bli1uHxVSDaIXFzr3VXSi5lvH9n4V
lNJe77W2a+X0cUG5nEBxqPHbWx8Km3ktEbY96ZHnooaSkh1xufKElC5f3Ko/
3WYGqbc2APdPfYBVnAuOCQO9RFc2YYC4mC+fSjVessY0vkjFk/m8BroT4CQk
TJ6SFdr97fsD0jrZkWGoQI+8d8s0bcokdFUC0d4pAZ2BQ788GcASGldXfngs
0Bc/xmuhOvEnYvtye4FjFNr5nATTprCNRDw/J56aBtDAig3O4kEvC6r8inBW
GLYBdqyr50zem6sxz4UK4i62H+hED4MVt9Sd3MNaT9I+HFBfdm+5HJeXoMsQ
PGwYDuJ/QBIkj8dbnOO9LTlI41FDoq0wL3CI9le6B6sRhoPiJZ0sdhly/yNS
rjG0JMLZoZGIAB8+gy9XnYMZ4ByBrya8UHixSWUjdpQN3ra0RjWBC5BaVh1n
f365hjshjmzbSq4yGWkqXtwqCgF5AQGOzUA/bzOajh0/9dNNwS8VPxEzfIZj
BfQudaAQ/Nsd5BSa737pSN+FWmI2FNvSZO5Z23iQA05Df6TiFNwDlmx49g06
egn/ZbvcVPaCn+ufLq/2CClZLahAp4o8+hBEVPfYTjLLs4d3Fli0G1E9cne+
jX86gES/AbqapkE1qGfPAWNoWyBr1Mhg02aeWORf2dgA5ao3h+lSmgKsSbqn
iCro+86vXl+zuaclK/VznskdX05psnuAFuk/MCqVSDnWLFrxsSb8+bGOjPCb
BY1D/zdrNfJ1acp75zo2Gsa31M2JjqMkjYSTio7CMMfyOhqQlJvhQ5n/eSat
V7jVKm9NL8YEOS+Hy1A3y6fCbOuv6AFY8h/kdOh3qeP3r9LrlTIPTZAV5Q2/
WkvqJWE4Uq9jT9PS5a+d7YthWxLAjHxd2vFsPrHJPYXxQqrzdvlnU2fvOb50
IvyEzc8CLmow5Dj2boreWpZHGUZzy5YRytjeq5qkh0BmwvAAW4gUjaPJc4sn
f12BNEsMxyA0H8M4l5h//MS2uxJ6imL+IbEZx5Db+O20ev4JscrYSuwW2WS0
MYQRS5HUbVsVGW5l2D429U2tqv7CpBrMuYYwqQ7TP45fFQ9kDg6zlCGnCXFr
WWtgwg61ybUJMtXICk5hzpdX+K+e/Jq7wCR+1cPV4/4ybGBXi7K2lUnHsMoN
VgfmgM1wjlqkmFVZxBvOH6WHUNzfZjAsvwBaveRXZfKrxDTzGHvX8csYON3m
tWfnQkrxmyfLZ7yljnp86RPi/TkibkdfHDNbXABANchvotItm5j+H2hWZhJc
zUay+Mg/9FOJCdjbMl479+cZcDBoSyewP1UwE4QkQQI2s/jfQI6oEbxCWeGC
iiikYdKGhubBrtpIy4BMBQvLkCaONSNQWabYl1T6PWxiwlnCz8z3M5MM42q5
6Pc9FuXZH+i1jWJLEQzTq5FCZbRuL2l6N1ObhuJ4eZzu6pT/XzF3zCZzlPCl
zklO1oyjgrTec91YR8rx/tzgTf2v5cnDjt1jIOI9lErk+AVRpdxsRH98s86X
m1dlvHtiyG35UI0+rMgjUtM4bt05N3jCzk9fi6h6EEE/ZzMXrdBUuMbFqgno
JxP3ywe+1UcX4UbFxm8+eAsth/+ZXovewWN+V14Tk9cdQ8UfUsOLv6Vn2zdF
TgBDGFKYC6jNiRmgHsTYWAxPWLoeVhAtGxeCcJ9xtrULedwdE1vMOR/sLjX/
mdfpH0GFGDhK234naIyV/Jnt69QeuG3RehFhG5rvQ82RIHjaiEYwLNiTmbOV
S7rMxCkmo5MFkvXclkRwksgQIL97oZKgBlE3BWBHimf4KnIZP3r/WmIRNiRY
SA9a7gn3SmCoysYyWj6qgXDWQTHnvAf7LE/fEAdpLkKCS5uk870QlSHKbJtZ
8ux0j8wk9km5CdmZVi5TCSsvH2aIoqvRFP3GrkPkaQHnkxvKCJiFH9JDvh0+
I/lmcVln/h18B4yQfKGkleE0MCRDx+eJt1ezkfUynuVIcmCONVzmQzShjjnG
zE79tdf2fFFwvdTjhQbRBciaR/P1o+UKD01ZEKpKq/m3f8zhVF7HomYDT+8u
VBu24eETzXTcCrOHaDkTTB9lKSnCKCfxdjUtuUUAto6B0KBVzyQ+NqFz635O
YHoa2oeKVvdILawYKNoL5ypLWbYPFleyVa+DhN/Sx5JwFv7siRxsNqFjhxiv
t17/k3x8s7iRJkC8TGi2yG25Um86AtSoKzWv1qRQccUcMQB7X4peBQhCKsrd
5QLezBrPv357fEe/s2AuNlGcvyD1P/ESGTNvNW2QXGTPCacPVQYAI1VFOoLk
LRe4qWlkbIPmojTPQmPK1xEFW+Y0UuNtIzwc0/bvnY75pU2ufZrswUkmGdWq
j/LCYsPFI5LH03hHZZgg0mkwcChsEjKNi2NK3T26ihtCUHMhGTBAZ0i4G7DI
iGy+fWHrpiul4ruwdAzlvut2nGfClsiWwEpahvcaFOwLVbY//E5LJyJIZjlN
m9Rv6oP6gqd4gr3+Oabmn2gdiIOyHGwdRCid2kBIK9OCDpU97qCetuKPGbCk
M7dCp//nJabk/TI/sDELd+UQRcxhgSI1EmcnWWOGNdvpcb/T1vrqfgAK1N/g
5XPGKr6F+KFPwGdDTLTfvQB5F1Lm3vH2lLk3nZQJZvzzO+UA/kX9kMzsFB1x
/aFIwZMbGJt4W24KdHNoz6B6p+3VniNJz0lgo0npdEljnmBYpCfzyuGVFUIC
T49YJmcx2szUFcKhBdn6qAqVJwd9ldhpA+qBgaDQt8tqKATHYVJEsCo0Bflb
53E3JlcVtzEneeyNYOBwbOt1Q/M+MJS++urSy3/pAK1QL1vYmDfivGISPHb9
aZ8JvCFONfri9IeWbbbYnXVpZNWH2/zA36cbZNarj9r6ol9l06WAgChOIYmF
VVW7CWXaoickRevRb7tbXFLwRNkmkGYrQmQBsJfNlHCVpDMunryU9tm75MhR
Te/V+oPLBtaoTrdRxdiGk6IiTert09lbQHmKYILiQaU3ft5Sx0nuOQhvD+Vy
HViODPQNfEOlDzmpVxcRCr65hWHhltXv/hL6IYkrc8XRTrEBVI9HyXyB+OAA
TjlcVOnYimyAn0mIkfpjwvP2tZZLwH32/szC1Kfa44yqcsCGkXTrGc1o7Z0Y
feh0bgVak/aD9upEsiiErTjh6htFpLBbQos9PGwoOksT4JCL0/vaGr5EXUBU
LxvzTYE162Jcx8wowiKRA5NqfeuJp0IOSWP25I+8qQVqKrPpXBExhkpqIZrp
BxwST6RDBlO3cGrFE35iYqiscMPr0RSP29geppe9rkcK1qxzO+qzF71MTynE
BcmBXY9Zco0KVhxxd1FOhm+9srD7bStKbMlQNZ4aFc+v640p0pvyg+v1+i+u
6je/zRfF846tb/dtF2iabiYRARJbaQbahNyJrk/j4NEWXLakE48+pZZB5Apf
i5AI+DHy3Whaaz9emEkLU0bJ3EeW19R11YFriQ8Gyssod04PblcKXvlfx508
oC+yvbL5jL0ytucDypCUK2b4pz45EEjnDgclx9HTGJebK5cJfxGW5OeLIjT7
qZHV3IOXVLhVHTkBZK1bNBZO3vY49XL+PxvTqFFd8uafqlE0jZwToNoBsOdr
iW9NN+iVirc0oTOQFwpKM6ziSzdCBzi2AQj7VhmAciYA9V7FSBe1HjR9gLPo
vPlCLgtPRubG+PAmQxYoti+ty8o4dZSx7yHq1QXLXUrxZWXUe+1aieWiwRn3
CVLdeoE5X3eGIdPq5mmo68jq119CEZ72k8+ePkSRFUkftwYicJWq3cAEARWB
zM9Ny7h4pLmpP1/16Uy6PCt/FppN7M3rqYG2ngg3o5hKSYvrK4i0TY87ejNr
DiMfS+nUqLu6HTtSMVINyA6ZXlAbaa7B0JOrl2AP/YVh/iTWrLALnbEx59zQ
BI2l5gnn+ZF/L15GuZoR7OOdcteGXOzOl6gco65AGbt5c7Ik7E/2tc4BMx6B
wUPltJqsQ8VY21rE/tH1U8dmQj6Ss7JkBsoXq48VVIz5PuxU+OY6g48vAeux
kbH3lDpLbUqx1LdHRVOLIPw1tVK+cyrAV5K1w+itcorIfiLkHK4y+cwIJhjE
apTuKQqNzW2Y9Fu6/Db60DuEOXqAfVBV1eEH1hOzcjm8ZPXUFqF0uSKO5dqn
JLiansKMILlHAYWJE5KbZab+LbLTzrgj3FK+IhAwfw6t12/7QEBnt1a07EMS
OLoNeEg2qGDVTQiTrywnaKKHVAtjpEYWM6qgRsVda6grBNq+73zVWhUPQMl+
B2dO8xWrgoY7H4lS5Q/VdvEVrURg+sbNoXvwAiuEzk9p4HZCxnpt/tMWkV/w
VBb9i2XbbPWQ+bHWlu+vyAIiEppggByw3GLDsO2sBEWYOEzxC2lYmy2/bBZv
ODcP582Gg24s7lkhDuNUE81rQq5Sf43d0P6RKGBYIUyLI2VPkvSWeiKg5hiy
YLMfwXs4rqgLbfjcT6YEgXMcMDzV6ix9xD2xvsH5tcLdTZUmXiG460tgABXl
3AqXrKsjZHoSz8g+OahXBfxAT1U7gYKVqHUIx7oCZnI0nMv2vskbSkwKenpo
eqoQZ2f0pimlcUOMfuj+mL8tN2X9AkADOuvHYfKXjdGfxdZ58CPT+CoexqxE
Ubmy6HCgO6zuBDpsZzR3jyNz9jK0I6FYc0s38IYnAF/0LM1haebqOJh+RAUb
S0wshZtX97P+c8UHQMJ1b2Q1tzOFIjhDcg7UbMrJ7kE/xlubSGwwkTdcUWzF
EX0zJcb4At4CwWDjXc1ocQ/I5TkHBScA8q86BqB64C1jubGg9iYII/hLLrcp
5zWMGG2N+LoE1S+1wNiZPI0snrIQD8cqJqrG8Grlz5O0ryplrTLNTwAAlDP2
VeY1RnJSk0Qr0vfcxohCEGXhJeZXHwRcCF/iPsxs2DGWTV8MOAWt1Q4yKFZU
7AO4aGzddLX30YGeUY2ZM1cEZb0PH5Tth/qP+FCY5+W0jmmZKsVE4O6K4CD1
7Qez1eGvJj1RI0goBkzJ5LuHDmfecLIr16UIYHajzK1io1zcOY3c4gw+i8oh
Pk9s9pNRgTLp5Q56HcF2BSSGQJxvJ2SKub0TthK45xDA+5OErh+wii4z+f1M
Esx80I2a3HL+RS4vRAa6Vxna1va3J0Zw0ZZnuqOWMpCDzmzk6ZZyKhd0z3Zf
C0FcOJJ5KRVVHOuzhA9N6KibWXWC0Muk+KIx2htXb99ostERiEEzFRHHcCTV
mO2g37cx3liBH9xjuXT4zFxd4agP1PVSyUhwCloHBM3TTOwsTImmfr+PxgMa
bYPTwlfIH4BfH253xafTJPIlXamNFB4MTlbhCSWxooM61hJITqpenrbsU+PL
U48GBNwSrqA6IQCvxpMov3RdKFC2mI+h0OtccX5KdYZcSpVemksQOghT589g
knMxXXeD9iZoawIs+/fP8hOY0tgnD05CfEJzWJj8FYjIvJ+6h4Sul0OskrQQ
qDEKmwGQ0lMMgiBR1HwQ+m2xf2Tf+cW34unkiJKvmW5hZnuGGWp93ejcKhzY
3+QWBwEFtbnC/5B8FcHnUQll9Ab/p8sQLWtbStGv2XPBf22IFZm0hCwUaaks
Clg5NZSUvkHwShY32btJt17FDjNNpIt0Jp8Jwbjb6QPD/5xrjwi+VRqF56mY
mMGLvQPxr2U4BULDRduabQ/DU5A1X/ROFpqK18VmJMhXYZ2+Hju8VGwk3RU/
W0+q56Yb0xIvs8XjUn4uV/2S0XoLQ4SD3QQS61M5FV0fE+OWmtbjO8i4Du0k
i72nd+6SCR2GCGuxIqAHkjUqjoCO5jVL/UKpKxcEla9BoSZNeWdjA79jN2NN
3IETyOUW867wGc4cSJJSU54Ep52ghVJG9ugPXr7tGVmJVPQayL8Z5PxG8a5G
0jXZS92uhjjoGOT0ZClsoKqgCAwn/i3y2+rHZElWjDn1/LHAFeENeBVgbpvN
Bmn53hHI2Mf5wLoAlqvZbQlFZD1nZ4CwzmlOQFa2oax2P3rdIbq+1y6T2ON1
AX3uIwhFRJksQNzW9Ay20RFCajLufV9DVy/KC54BAOb2fXRpL5j87Uz79ANQ
kzqzzfi93Yu6CkZzOBIp4T+mOFH8xiTzp37KsLTRVw5mw0Fk05eA6UFgLsUo
DuEJPe2+ooK/p1CUQ+7EPWH4PpMfJbjo1Bj3RFvUDa5pCefN1W2BZQrcVVe2
VtB4HIik1L0nfzKnwK8BbCKkmqJSo+Pg+1alk0s5C26I0uTqhaEgcfVF2pHE
9X9aq74WaVO7Fj9QC8ol3NG+6D6kSKTgNeCKQKOol90ax3+y1qR8CmVklMYw
NqvH6O83eYU1QXtu0Ld9ddDBDhXXWebG/0pRqt5J0oVTJE+eRnGzE3YZbbyc
KrfPIII62AiL1u6zNKFuG7f6DjwTXUsPOQ7gq5rvJyIlC9tkxQR9kGcxGH88
pHFpJqnB20gEj5D3GAFbTSJqbjea052CPUjE9BnVc18XE74yeKLGk+oSpsl3
ouYoHZaQ/qsjZRol3DLUIP/eCdtJa6UJW8WGXmHDBN7Gko6pjlm3hD8y1ZK/
mHlrZaH+1a6L5AjtIO6BPW77xAFo80rSnsfhr5mFGVQbRq0LO45yMcOlUzsL
yPF/RkJFlinMPI2TYxeVOXYCWqO6kl/b6Sou77myj50e5TA1QCiAPJlq2Rmy
uqAIwDW15L8yrgkfSyKAGdCSok6X04iUF0ZZ5uSCedrYqILakpp2deSOQZSi
PjDyhphT/CeeFp3YUpx3GfI+h0phtSwYD4LAYN1izEZQrUEOorPqosxeNezv
j/Qg/lifJpBcdVMLQw05PayYr65YlWD16K8UCykuHYbBMRr3pUdsxBmK2v+5
l/gq+crn1FatqVve8MEe8GiU1eHKAtgEvsLO7RtkWT3vXOHuNQjNH0ItLGYc
BjGj8Xzl/tHZp5lOgy0lmTjap2eSGCifinN3+wm6RFaK9ZjyK2OFKT/f8uRs
CaWpRPbvN7lN44tupKFJJN5ptrZgsHib4WPk8mIXr8/3ZRuEb4e3eKFS0Qzc
4j3qfQo5oTRTUfvccr+HXoy0CzCTnxk/wofqHzLUlPfJwpiKTxf/FKsH2GB4
Kp/eWltlam1E4SHv3v7cscjj/L9sbIeiKbEn17Vx0ANrJn7S7z2i1QZ1inGR
wTzEYTSO32DKrEhWGBmmY+7Aog5+XNxHrdM7/SpZmOygR5fV7mSiW0la37yH
9/3ekdMY+1BJJ9OLsx5GzAVQdVVi4dfbo++yG5vjP3eBUlK3mjRkWDXgpx5M
Y/gSOk7e/Ojm+aOCfUsyD2EalpXsNpwtJxASqZMddhu8HqDINDO9rvE2q/QY
1lrxXADV2xUG2GX4EzI5jSq3LtNiy0904D1yT+eZQIKPBklStYrrfYnOpoJf
DI/FhCFnbBVGsQ1imTq+rhdyRoSa94VF0ayxh5uLwStJigdFfcLpt7m6YtvB
o/m2e9exWtDw63hiiE0Fp6lCtTDuHKcZIiW3BO7m7hWzYz8uuBniNEVid+ej
2bcjYfZuTDplTxguwyeZ3sO0kxHVQBMTsq51v15ZG4go+sBw4+MQmBXxOY1K
6tzEEsyvxze89ELv/QcyS2tmQlfd0CZwAvBBYcbIosh4wX4AVg25OcxWh3r9
SaymgyyYoFdZ1kdHMbtRnSgWrLca8BjAl0mAtfDLLxOd3opLxpaEmkAY6EgU
GHw3eQXMq2xKVD6mNkSIRCNPOTxKM1L/DOx+PR5O/sls16tKsry/uY/lB70m
3GDXyHFoiCAjIHrLwlZ/0Cm+CJ9qSrDHG6xK1ZMLJEg3/341IdtVktaEG7dh
IwfrnNPW3+rWA4UR/BUENhIGqzj2cXT/3W2LMoLgTrX9EEDXLMDlzY23yoHM
RzkOOM8sfbYoYTgn/I8iG6sF1YHXeiFhm7aKzp8LkVAifDjmgzZ3GjqDMa0R
I3rf57kGSBZgZNoXGSTU20DTgrVwMG9OLMlA6CESRagnw+MIOwGMol3OZ0Aq
kSC3hfUrNJ2/wo2BJ9dXAH4AyZIMAI/FW3IAIEDaGVahrOj+WbaQmnob66yV
S06v6qDZUA88UKz1zwEl9GL6uUtXdJC+ay4LTCAbbbLQ+P/SRLLzegvI9jUr
PE15TPMiJz/7q3R3Scsrhbr6NyCHA+1S8q9w376E7a712Mfzwp/kE3YpWfSI
25kRvz5Q9f1z8L7jDuKBGBCoUJiK/EqrASLPiaS6cDl9tJKi8at1ntIUKGpk
yHvfnYpcLMWOFiPzh3KHM4mZc99ABxgOuCsePXw+GxmQUH5wxPRgx/jMczrJ
aliuFlEZEsSN0Ov4338aIKQbgVrCEpVVv3eQEIuhuU+ml5zZ7TQaz0GdxWZz
xbJqjnSw8H0s18dLVzoO5fgZEy0ieOrxQzWzHSKtU9/j4zlLIFGp1d/Uruvc
1ge7prhETxywtWgBLhwWlrmm1J1xwTiP+YQOyZpfOUSC4OA/QygJRoGAlUVh
L6p8pF+Ue/8YJqulDJoPwO7vCnphUimeS86zsjcUVMuh2NZ6q6d3aBP591/j
NGaAHZNrDuxdmii7oR8PNa6i5EjOmO/IlCJdv+WFCjBKPLkTrf9+cX/XTbPw
pcr46ozK7qG30qJtqWM7RnxmOZJyipA7EmQH652CQh6uH1AJrNyVQMq2oCFz
9GylCBeXgzRodoCi56sHMB/CuNuZQdK21Z1rtbjRrW+4Ndr6fMX+PNeHmhAS
llSAnKIRSC78Nl03LoTJIxfmZPxp0+n3U3vPJezecQBpeUhx5kzGMT+S6ztT
O7cs5yIYD0qBt4Av2M22eOe+zDrYGA5JOwCPXP6SoVTK91Hy2O+mGlMNwV9Q
BuP60VgztJacQZoaKGOC2q6ONEx6XZ5qBZp4x3JHMiaJREqu1fP0nzuqDvWa
RMuuSZ3IOTYRM9r8VoH39j/MwsGTKVps3bcy6qEEZmsMP/P73SEQJ+okaZ0r
/+eDAtKKNcxFJpWWy0V+W0rhwgLDDjcdGZSeH8/QdSuuOo4aWHD7Pk/uhgq8
KvWsWXFHSxE/siCgZQnkqZBCkAW6i0nSgCwE9M6v9c0uxDi/OxEaDivHuV2w
blQTRpzWPpKBNFwwKUh8GEZzwemj1EQA4LjshQngOitC5v5e6Ie8qeFqhs0q
HAWNnGu28zpSQEX/nIr2RINqhqPp95pu0u3ZPRYyaxyhTzaZgGttIz2thMnR
+Rbxb83B3a8qbEyqZIH99Q/s2VpsFTevnfA6PlVmxXo2vNGrQaq9AtS1v5RF
qnyPxcSWw3oPYZET98kGggXJKvVpj/G4LaEuI051a2c0Bfu/ZWv6wAu0pVY1
OM3kG9bNrlNmpBwnzh4MAVSybz4HEmq1TWF2Kvso+0OluAzl4KO6gdUHCm78
jGPgtVW7ZUM/PaHjYFt7I2Qm5z4oimCLhGHm38XdaV/vXAnGxfrXEe8O/8dw
OlArmPQiCYIZXj1Dd608+Iu0dLe0DUmP2FTISebVjG7gkmcEJq70U5TAPoWS
1i2xxxHlqriwybyXS1RO+TuL838731oFU0OFO1VjOVrgY7kPmrq6pPXDPkO6
XCB32GgMwE9vB+a3Wzy2vCBOfhNwRNAW9JAJ6fsWdAyacJYIqf30DL7dK0m4
KO71QbwsS1FHh05QTw1LOtSGvEaCIoN5BuVCcXtPgouIMYhdZwlTsnPgk+sH
EXzQgpMTEX0XtjDigdFgp5HgJWmO1pOAYXPqwPfO1fNIP7y/7Mr5FiErORT0
Y9XW2fEIVVpIkt8TY14u+5YMj3uFHvuyQQalm+D86hNdbOE1jcimHM+QlbXl
/LssrnbIUO3U1lt16Sz29lU2Z77lwQrlBu//CSdkBL3akr8NZyzVJrUc6CAC
ms9+d/soDXwz9M3FMlWV84YDc0LqkQhB8gQOThLuiU0QiRjG2AbZvQoL4YA5
4AUval1beKvGCflHFs4dZMf+47XLtNr680euw22oWmxlqTQCrW5mn/DqL0zt
ChCeUWXP+VIpwPTjmG4ZATPiBen6yh4k2SPxiWXPLpIPzzMAz3JGEgLA3fs2
/0h8vkbJJYftS1z0+MX+NHO437SZ24lbg/nQAYlAc70aEEZqlT1lJhJ/2kOd
Sm5xs3/753QcIHiQ6Yo04EdUfJrj4Q9VslXSb2QPLza0Nrhz/8dUE8AyIWXC
iByoPC8QD2+matRaiP3a7JOvMatu3Oe4teVaoigvEsbS5bQwM8eNZZfgsDDy
o63+pafPGnEew6O9jgss0zykeE/vgZa2DEBiBUAaWq/ExiTIeDQ1AxlTF+tF
EKIeKB1ZKMiUV6MrnxFtoD7H78O7W/LYMRhzvJ0tdvfuG0k7S20MaCs3LRHR
yVuBntTn8SmDmODnXlrVQF0otfi8ZSSZ3i8mPSzimBZINONatNeep+yhCIAh
UtOrFn58fpCWP4NVHV4nNK6VeC3sMoTl0DvFhjvYvAHsMw1VfmF3VTxN4L65
VmsLCSJAMw54+WDWJ3yo9SLbZ24QSCuL3YlymlWF5jG2lH1u8R0vBBb5PT2B
8em41BpJRUyz8kibppu5JIm2kKAXGNzyrgdvGHeyjmaFZxNoSS9lZWqk9HD1
pJRFLvwprtu4nYRjbTYcyUTeXeoEyBuPpBJGJq3myhuoUOfcN4E/z1iYUG63
DC5zG9gIvG0n/Bf0wRP7ecYYhmx6RLNz7hlyHtra49QIEZo4hN/253NmYA4e
q1OqjIQHOoBGytNndt9wElYU97BaQ+LinoAwzRTVvTH7yVIg4JriBOnAMhhF
Z4ePgs5n6qEvAfXWHnK4Wzkiy9Wv08vyY7+wky1N24fn72cyCic8nW7TewPP
6nrVBGFgFQICJXncjZcAGN7L/4Fa1GcWFXIJgoJvg8/WSug2c+A5/MG2YXxA
XlYh6/+8xTMGHanRJxGwMfXmYvBoLLhhM45UW7Nk7rKmzjm8+ij/yTzKb0th
BEQ0RNsakZ7mCqYBire5pMJjJWxBrD0cbGgX05GHgjXoT+jf7IXHBvnT7i1M
LT0R5LbTRhckH8QaLGU7NkXgMnRnja2y+PYrp5HxxlIYDLJd89BT4Sy8/9wc
ChptmsAJ8Q7ySfW68srRDpHDdHXWMDvhYnGUQ0S+Spp+aUhdMNlsRhqeXfFD
/3ta3W3JG0OJb8g2qGOG/8aDwzDS6ayoHOC2oJ/PfwDPbiRTXHqOFvAqXxcs
xWPn4+O+JoBhCRooYlva1O9/q/nl4czYfb+ZPcKRhdlNtLQz+6gZBa67hKj6
O3xkZ4NOoSei1vlf02RKpFtBCrX6f6/9is74IZfAgUa3Zag56AQ8FIPQ7z+Y
7ObbzpfnzOCmeuSVFUXhfCG6JF5aSFi02enJ9f4+fdYMw4NcjcEbUXx6HcJb
BFUvcwUwCnKwEgSNvos/Fo7kpQwhFQM8HX8JNGKn2PUXSkDnGmgz/mmZTVZ3
klfXcLObNe7PiJm7ZEpp4tHzOAi7NQDmLP+Yrfm5DfDroZjb7/SjBge5CLDw
rIZGaDq3QgYBF+Ox62R0Mh2J1DrHpCJsej4PAQmtHhURQcVJ2N9mgi2jm0If
J/Pz8QZ4wr4Z22An/YTAbauu/cWQQY/rC/08Nyb01p0seBlS/YZzhVRuFxGq
tt8s4d4GsJwZ3OJaWdI56D29V4FJdXU6bWYCexUVm2eyQB8MYeUvHTU2VWHV
4/wZvcP11mtwf0DBRyZ+UgDDRexX5tx74vYC+dYGx8UiliAIlWce1+U2WUo1
jisgBBsZ6uvCM3Dv5QgluEK4qKGv+wgP1+HO2iECtwBvdTs1QLHR1yVlWteU
WPFQ8qVfSi4IRCnXL7DvfNASZWwEyIff2W9CFK1DcKdpaFw0OiqtsHuPOlcw
EDIT4+eUR5x4DZTK2XjT4Yv/vy/waUuf9KXh4EflcC4jiEb9ihuSULaq7BOx
A5M3ndb/NmAiTYipf5w0zM0BX1CbUd235AwWfs0OEVt9ehngOhrjumbldUAa
rXCP1OR3fvyvzGa9KMMhhwA3gGMlchC2eAO1498YHs8CdST1J9fsFsb/BCb+
YT9PVrEl4fRBGo7yZrmj3yr1kcY=

`pragma protect end_protected
