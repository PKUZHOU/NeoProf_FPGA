// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
hxD5YM3av+cCnmkYehFZC99JE188A7LI1kD5Gje40HeiwOCC/fdfRMO78Cx5Zi/9
CSYtRrJVj6bNRqjkQBMDS+h6Ej2sfSUZFm7xSTuszo8IvxEP2VTFDUS6mzn4LJNd
k+ahSTIiiiEK67EeMYNrCsyii/npGbXuVJGsch1GL80=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 12272 )
`pragma protect data_block
iX1Riuk5ThxTOnPK/JEJ79ZAjZ8s6Xdwvw2C5X/oMJtrvgwBw4ulMZRtubyMekwp
2iEBRDiD1abrFsNGaX/5jcGiB2VoLuvraTXrykFYcB81phlYiu3sH3DjKzZ2g/VJ
Q/Erhyls3jBz/m9kurrnKN80V1T1abNpHtP3JPRPfNTBUMHNAmQOU1HH7S6CRO4V
4AhiM3o9cyquYfYqvfnK5NQ3M2MvVxzI8NcSYPXmwuPn2zgwpyrf4qLV1GjPhzxA
plsdstN/h6OBPGFexFtnY2fcHljV+UiHUUce2i4vpFU5QvZM/3CYpWTldYdMvmyl
N92/AoUlb7PwgjL4WNCHFJ6j34bMQAWRou4WB//n6A4H/1RTLTwA7CFPvj62pIAH
xlCXBbPuhEzXrzPLXSZG9HzPZscvTnBSsneXlKRxLBrGAy0H5RxUnD9fqFZlhFmj
0p9JoW4fH/cSTlCJdGl4J8PBYio3IRmdoRsPSqiagSsbFA+EsAL8aiEfX71RxqT7
livlTAHdgRx57KJdT7vCZp2i7UddkdM8W6JsG7AGuiQrB9pWroIpCFB9//sWPJcQ
kHjM6d8J6ytWMAHgOqAQ1GfEKNKtrVLyD96kgnYGdr0xfU1GKg9VK6oIHsT2IOJ6
Qus1aiVCqX8bdjGP2N9IPgP0RHaQ0rHN5eyAJ10AXPyKiU8eiLRLvNc4oUe/P+Hk
zh67eDQi7fnI+H80B1QjSQ1z2QBFjn7dpXSz/EMZys1gsBBG68dlpziEZ+DX+Hq7
g+bC1gomRJjQqr4ucghyC4nD+OcOte95UUF8Rwn9KjjVB0K4COJtd4yQ9YveIKZe
n68JUkKD25OdZnZz14dZtaJeT01jfI7PL+uP19bG0Hzmm/Isoh/NtJSljBCMVuHE
rxEwnjO0miWVZResRrirSwX+Cma5yO0w+I9sB+GHzz7ATLuuHUp4RWi1MviG6uIk
IpqmmyQ9C2iLvEt1iYiTJ79yjH92e2HxyQw/njS0ZrdahIR5KBst3QGiULA47H2S
gGY36t3++l5SGHyrWriqwH6ZCOFVo/eHWtmg2XatF4+zb905SMJzu1WkegEp1WG9
sSGHSUb0UKE7+cm/jD8BFx8PUe3/5B2MFB4oJmUgiUtLChIAnnBYgszMBkaxNQbB
uM8uEzo/i6LqmsOnuxk+BRfFAmEPO/2oE446Dz06jlLSWq0vaTh0SgCUGEC5inMG
CV20ehjIk/r9u5VKrtf5JL2ImZNIJggo2ofMwpyZkDQaVe5Uztm9KZ2R+C8OlM6K
4ASubFMx89knujULFxsadEMMgUA4I+857zk40tuWPLIN9BciFLerO4yTdp3C9e9W
i8XrUH31oCCE92Md0GtHD8m9OqWyur3BGpOLJBpQawrSAxBKY/aFmebFq8vrnJIU
mtp9ewTHZTvbAWF7f5/hWYdd/TdbLHoifstBVBDYFldd8Nl7uHzC3W65m7iyQE+V
XK+blcDqlkCJ14PIXy3gR7hSKWXU7G9rD7Gr0ngXsxIt7hgewYKqbYrwZzJCKJP5
PGyE+bhFCMf89FBZsFSglpMNLt6cs7MxJC4xnHRVUEWCkZ9Ir9U8yVNy+6CZ10e0
hbJDy01Dy1gp/b/b00azr9o8J1BZYJ1tmQHC1+7NhLB8tjI7A7SrXN0QdRdei9ZV
M3VbjVTp4TxWrLkw+iGMtx2V6TMMIYpAs/ueh1mvl9LrYMBQk9rqdmu0A8MRYWae
ofv28qytJ12Jw1jUwUI5MNnyG3T5QN6BwV4acCEw0tejdFRPTThz/iExW8fZJCty
VVGogjVNS7gjSNLzhita9YU/neUwy6huqakMu9litHlPKt3TkaTu4EOt20QUl4t/
PjglcwI8rhnqZBWvAHuXnzifW16d8dUUSWz2GytHVt0WDQXz5d+STc2UweGvioZ+
hrn8G1/u/ePpYD3EUhoZDzC8SW2WWtuLJlSMzKbzvG9Bgqr1CEAwm6fs7KTY+aVZ
S/QfXpOGChnzjh5dpgF1iJOZqZ0mlUuiH9mY0M9SXQV7gQCGVAxebOL2ldm+rVsg
rvv2AsOb8EA49v33ACHQTwAsyeo5AbuAzdI5iaEedTloNtN8Hjd/nH8aX17Rh3L0
JNin2+11UHClUAF0xqzPDUe/r/jcazjW8yr3edaDvi3TFUSznkA3PMK9So67e6TV
dJpDo0XJctYgqYQQfvWdiscwo4XBySL3iyNb85T2zP2gMgN1Knjd6w29KvDOI/c9
qzLaOTYp6bu67s8AnhJf8RE8DzYPrNygNDI1RVNc65wEEIcGLZUqs0zj16n+G2tS
8CRRYCNsiOu5gRrEPolVuheOzaPtYdfGiaoC12Xa3yALSuvPiqyJonATdZiT/+93
3cDw9Vo6oyYz0ExAzyciWDHpgITGDk/f2tfuZJvvJZvNGNNpV8QBzioODKbUdTn4
goqTiNEd3eoHsqjSk0zJc6P4du+m6ZZUhvTp7wt1cO+SXn4HN6GkEnyk7qRGAZSX
9qLEOjgY9AM9sQOBehXuCAZ3Qy6qMsiHbwuktc5/zZz/rQpWHeAmzf+kwUrvDOEb
wJZB7XXdlF5YjVE3beD57ZwkpgLWATsO+1C8m7TC20UAuu+5AfDYbymYrliBGjxq
TuouCBFXqU4JMdW4ICm++cnPOr+Pr+lQHTYF4YdBWaYxj5mJxNlMRCoPrB8xsgTH
KcFhT/QilorISV0uvPWTv7SEJlIa3cpJmBQjX5JL2FOAysBrVJB/ERkyG7k5vCpM
iTve+qmP7vHXcoQ9+pc3DtTEri9BcIGoKX8K0Ig9xVoFNSfiJCL3srwxdk8yNWPM
Gfpfgb8C2kFFbSN30oiM99LPzBdJi3vgLv3cXW71p5zeWNC5E7obXOGs0qpJtCRy
23aUGQSQ5flGpIRNqrYd0ACC+YThj2eMK7X9voF+oqRTbQxoeqXr9gdJB7dIj0Te
f8pq991/gLuoLDEqrBCZhcFiGIsILXDfb8R1PItzwBWpkhFczGBwYOMCLXEHn8Y7
h4BzR+7mFM6fgvSJuJSnGJeh0IMUUT++1T/ReXXLz+GHY1D/7P+TEHi5ek3YG2Fo
/+TWIS+eHTbQ6LkrpzMLgBcGPIyvoAYWQAOCIePG7US19gFMnFp/H7m50DUPuml2
ElGrZZBiUOh0DUjJNJip1PpOtT9X6dGAluKgR8svmcdQDp9uLuH4HnLgOXg6vKYe
dx41BtH0byWfx8zu8bbqeeyPXo0XDc/F+PFdUkt9PNegWzOIZcZZilOPApxkxann
FMH9700g+DA/65lWax2G+oj8+hDeGwKF8O7W8LL2kGRBvtRGpSwQeNOc4xoLm3mv
deVu6m+oEuhh2YBtsKqBCusFhnwG1zS7zUGI3bCTfphEDH2Jfb84HN1/PAHeFd4v
kAtFWXL2t4x7Ud6NAHawSG9aH62RnZyoa6I5E/w6VOhekzzAQjk+gCWkgbAcXQgU
uemEXcviQGMhyt3zrJEG/gj8Ka7YhAFMu/ROptX47gtrnwKZL+ImX+rr4v2ykq0n
R0wYowtNfa18GFb77PVdXFUyVPT5OdciBV+shujnrbDfDYOlTvEUVzg4bLvOwdbQ
C2Xc1QTUv70qBtNodOR2vI9f5wNnxF+xZ7bD3hz2GClBFYPIIev3QvQLh78MuvR4
LYWmCY1tUkteYxEetYVkQKymuX3P6I+Jm4TpKkPNP1DiBrdoHlePPn6z5sAXJ5n2
7EpOqgKAjpJvbHlfVYB0E2CtuPqZ/4zMU6JfEOKuPg17DSeJzSBIESNvpgMXQ3xU
K8X5tYi18xF5rBVb5n/OM6NRzwV/jn5sO/gIO8mTbAEnPKYAP9L3o6xSX/nz/Oqz
tj/jP54fDGIurdwH/CrcTZJPESxEBKcOBfnpKBuOYIfTRIP1I52w1lSSVsRU+wWT
yKpn0pyPQSXsBzjB7NMf1pO/U311FB6Omim3axTsBNfF/2CUHMGOFMboGK2Tx/np
1/KZS8kaLiONXcO20xEkLejXBE4E8Ri/UlTTJtHcHLsHmGF32VNJk3W6sFef3ELw
S2w3MIcYMjFqby3QklHd+1u9/bt5mtrDT+xd+08Q+inTu0G2vQ8Z4Fh2XQCw7zHO
VaESTXsjmJE7Mxty8ERo5TO6zikFAY0OXzRm7gXggVNgcoiViQ1RQUTHEH78eb7e
HQRgeOJLiXTc7jrD1womJoY9pjm3vEusia8+nMwqwOJ+HRyKgAUPCLDBTsuLcpVC
Oxs40f7915tui4sk1Cu7jtaQLvLsyaJKLQEi4Q9ShwRwhLy07YmWOCQpYj5qrG3b
W0fIpR9CBmRlPgabHC1WMkLOXmHxNDOd/zCNWK3X6Mrlvb2iAsRlOLAHbFamf3wf
yzfmQz0kUM4gJuFhA91OalrEhOrEEQ4BfiU0my82NYb86vfBChSiprJ4eESuS2yo
HYsSCipv5cJiVHLFw5YeET0bXoJ9NOEccgizWXOZMjuDaS06+1JyWEyky+Wf1DK0
58RazQINQ8ATtJMaxHhYyuGpNF4/sAyJi2WgN9Z5ChrSoWTOUujrV6wZdHFbaFYq
fo4bs4JsLPugX0GF2w6V4OXsrCLdnOloaqvD81fSq1+0UVczH02QSWKr908+O/qx
ha93rfuiFsbP1xeh41c6aidXF0rOK6KbhMa+Whax/2Q16+0mnoIGwMxXg+kaUK9Y
bJ8cUVuYFC2Fz72q+tV98KTerf8haB6hI2ZRSlgPz416+syXoNNa4o0TsfAw+/Tw
qC+Kr3ZOryRdYEQ5HCoik2NH+wSReUsj6FyWeDzO30Y2ubDfN0ZTApmma7GRFeRw
1QCSGqrXQVGrZRkZq2vDNm58Gxil+KDhlmuZV8GXRdVXnLAo4j87X5EOOTEZPOkK
81+O98sZro4jn1UY6FXOJr6GwS+PaHsU4pXaA8+JodH7S1S2IV0Hc4ZvgbfPATrn
rs916PCgS5pMOCP786JClV0YpTe5XHNZadVUtQXY9qHGAkK3NTSQWA/2in7JAZTp
7l4dDlRhieX7nduIMhxKMxAhn6vGxvsDeq5wcPSn1jlIt4f/CfaHrriPFs/MComA
eYiGA+2X1712i4dH7dTi5q4/5rkuaWtcRodsJPwSnP8bFSs2UbQZs1ZhuwSUdWk8
FMbobj1GdX0Mh+bUaS6PZiFy97i8RDiJ3SalJ28CXjwjdX2wvXBZVQzK6QNS1UGT
2iG4Td3l2DI63wxS8bFQbi+UqIygVc0w01/kLjmZXe+g4Pf6oh9bpxlDQ4eppidr
WQF5ii6bGwUMuHitjJNZHfBpQHHMVxwbR8HAq3Ku9RakPUwjc6/+X+yr14tsDcKa
x3FbcpV8qR+iKEwxQqH3sAgMV6HadmlWu+JLwMKw7PPgTL9Lgk6LJfwdKI8vv25k
GmIWm74iT10YgSpIyrAiz/N4ODPhRFniPsMBAx8QU1WtbpjcZL2iUWOyWtaUHEh8
Sgixat7LuPX2cbnNOnYxWFOTxJNz9ff541hMwBPdl65viZ+Mi3ncdc1UegLqspjq
2ItO/CV+S5Ws2EAre1fs6EdQ53uUbaFAc1oHVUEIab/tQHpVUQxE/pKIg5ZjyWEg
YDcOnI/5q5r8Ty2FKCFlGs9yuhBB17L90pvgfZ/dJ56G9huXKuIikIribjD8L4Oe
0p4Dbqo0T30Zv/x0Q/2Aw8DwCoskpWFpbfMJguqiQin2fNDacMbxgGFxz1jbIHQT
hxViqIjS/aT1Auivjvdg0ZAxEV8MrLB1PGQuxRKDupOKcDxWFSJDZvjL0ForDP4T
UHOcqTaC9/cIidHc7UvufQEtzapAVt6vZ2OHE6lHNXVPa3HXchLlbcKDcPOUYhmo
ZbUlbi1eq648SOs7Jn3LXBbYKyiZdqAGgRBamKCDZb3/g2WLHIZSjVMj0ThA8KnL
PbdjM4qTfMUV083Du8uHVQDrhqWInxaOcglxvJUXrV6VIP/y21vZwa5h9n37MEkj
qGQwaKoxw1478MuI78UpE21efJ+uytH37l2HVmkQEuRobll43U1xzFtaZdSrzlqu
OZetY2KjhZ+Q/7kw+JuB6OoBgx5CjEdsJLJOm6oLtnmmjGxdGOk9AhR//1CCkaLx
fR6U5vcUAi1ENWzyU12RcXp/mTCdT2siJkKDzspR3xf6epjp1J88unLO/AYyrqH/
fovGP47OE9aUyYlUhnKkkHq7IZH49A8+7ipCOHMPPSYb/AdgHt6r5WE7UZsLhFoJ
6Q0DKb7YuSnj+pmVLvkw7YZVdehcmmoZEUpzF4knGsg6oiz5nV1YhwYbKJs1QOOr
lxmNtETaI5h0zbHc7L8veDZhh5AdZKhblKMK+3XuUi5ZaL7DWzRyfvrPJHa3sNTj
lgGFvnZRisPE+V7o6Wf/40bWRcYTWm6OcHAiNu7gehmcRJWEduGGbh4dKLZLYBTM
mPDxo29KZ/faC8cYzcsgUBCweX/KW2Knh/fdnRPEMI8Azu3NVDOAH8jfWgQ6MCVQ
aw8+jODUyD/bTt9kUVBK7oCwx6YV7BiKGuOyWrn0m8mdZGPNJ1fSZ7nv466h0J+U
Rz7fnSr99uuGVhZ7n7ZH+e+e2FOSP8K15j5YmzPJ4txnDWHnxgpbhA+AhKisEkPr
u7A3La/R4q0gehk6wKgEbKPy/Tmzd0Oi6/n8kvRIaA7dYDKk02VZUhFtZ0nyeZse
1ZVEFkdVGcR/Qq7Klnr3pUZjOg1zF2uS5EN+CKgXAjsSsUixwbIRHhDJDvDqUNEf
D5MkM5pN2pTwV07Z7l5Ax1zoj6qyonp6C6pgfMCHUekbz6jF4Q4Op3/6QvYDa/v2
HcIXIEaK2FeV7PTtyumw51GQYVH+JaEqVESRF6qfFzf+NBc8Upq4BlRYblH3QChA
CrD9vvXSH7MjDESYjB2O4pZuo/VWLXF9Auy04BWz/d/qEgk4Kk/TxIxIRX0E8qUN
kDNl9u7Nu1s+LKCp84+nFU8PhNWXx0AwlGcOIP1JqA5DsDAIJnjM5M+wfls0q+Su
avxqD7C+9TdFc2Utl60Kwx877TAyZ4EIyINf+eAjHXXivt7IAvFu6mR+wFK6A4yk
0LR5jG+vhWqY+ch2REjXUzJtWVP77smR+iiC7QGSIZlylC7LPEHXJa2yjkqycgfr
WnrCMOf8qOvlCE4zgdoGTVmoUzaH4YkunoXRoXlUVbk6eLreUsVE0x0iJX0VdNVJ
K8BwRz41H54RXU7XcYP9RSCsPWNBjNDkHljWPgnSrYkpwOKSXuJmHy9hoUfzr8xe
If3ANOSJJuoEf65T1wjV50YiFMvRt9nBnqlvUesuVGyr+dI6Vey4JO+wm6+OHTTu
koqZf1sxvbOOf9DBLwvt6lwrj4vxyNljZKSd3aMCce18yIlA6cZ2OCwjHUkEeqY3
FZMXQTREeJmKh7d+gsxLNPFWQ34+4V7egPJS0a8CvxKBGhqmaLpd8Vth7ViH41+r
hjajbspajGKx5w/1XeXKUiFJ5W8R6TZLoqUDQrGORVmDeujhitTaypFW3ob8CZVt
1MDcMwPQR5L6WcgtMscGo+zr3znK6mVB2B8er1H5ohtYuEed0DLZuKvFLObhGKg+
muiZzI9n/tJPRQUOm5tXpJdfxdFrheg+JXQTmPE8oqC8Qr0lBbgscfR7tj2LraGx
gsvCOCNTRjEjqmqO9DyOSxGymDyy537j7NNbkWGP8fI/ozleJml/a90lJYklmY2X
t8MVtH2W/ZS/NTVxKY0uVu8sG7pArc4ft74RhrT8C2rn7GUKUpdkVjJ71+Ay16MG
WUX/0p1rtN8Uv3ofj9YrOgOwIvDtNLflM4VRRlLcGXhZw8ghUyC3Hc6UKhIKoMLh
+F8d+ss45tW103sznPjI8bmEp37FertUz8G31Ho9kznEbAe/6XIAgAOuuihJ1naD
qIGqxzIUKQgHqeyAnHdzoun90ssUpmDpFB/VWKp0hwZvsBTZ94HolK1cZQ0cXpGu
PJL5q0KHyZxw4NV2IgkW0rFQEqwZEV+5K+juCR354llVC6A9btNjhPNyanClZQCA
Q3hN5KjFmmZtkUjC6lSr5NkQd58KbbDvLEuWR/cW5tuxjDj9B3bn7YMmFxyI4cb3
z1bE8UVpUjCq5BK+IAW5qlK0rLiI8xE3e8BAU9xL7A0/gdobpnZJOljF9b/VZxXL
YU3pxtpoZc/Q2UJfnaxYSqmOEN93i6PQWkA4M00wgnD2hFcjITGEZLsayhuE8uko
PrchNzZydpomzKpRfp1GCyr3a7oGapdCnL8gAvbo9/yTzqmPV3drGUmJ4q47Idb3
pCgX3riA4glCo0FApXisB7/qJhn0LL1+5+jTiuLDD/N5ogKpwiEHzgpBbxUsqjvo
2qSxXEYQmwWTXjlkNjjwyCPcNPIX1zBr/7q3nhOxV2Z1dJxMPsCaS6iIOrpQoh7w
iZ5mspCHXtdRZ23IUVeLYmBOy4qItj76WcPq0RvDpKtbiEDUcYDNVk0e/oF7VaVT
KA3DqyipQAWp93dJVzSijaQP5thvW+AEkobe6UJJwxEhMU3ZzhynrFC68vos7yCY
5cPW+SDY466sAD2bhqKb+M84hXC1CplAVV7mT8vn9+PhXvRQHns5aCwo5+8rQlpp
dnYokP2Oo6RftV7n9l/ZAqAUZZF4/b4nsqX/ZkjJKiC/b1v2R46daHFHsvpkIG/N
h2l8DSR9Z4TpmZrBdcO3zQDdIPGGFCcaMYKnarAdWQ1uPggAkk4VLP6GNq39RoP3
PYWzZcr6ucFUgJ1GZbSV/weBUG0vdo29ElE1MmJgsddoH2BEynol0y/FnKMpTn2e
yCUbNVHWes86cQEDZqLEVe2d06kXgIFT2Bw+Rt877J4Ghd4vV+5cpCpH4q1YOvLz
TIB9/ylFJIGA5Ai73Xn8x42OgBBFIg45xn/AElNpkSCzwURn1mwlnoVYOwFWMgE+
LFS2u/wfBgQBpUrA/8G4I3KdQKtVtaItpMgOgp0+scENUvqh2HZSyj/Zf4KdNNaX
cbJzRyZmjJxPcMXKB8pDcfVZr1dg8NSPq0jZvXURa4IOFgOKFTnOGgBBDskcZpQo
qJVsTzG5xouDHWUeDWTovwnQwDke6OD/CCuR4BYdMEN1MBoSsE2n337ji4+lmoxG
WAIoxoqI+EfuiQ3LTanVFwU/Hqp7MxOPbMWtF2RbdNGqfLhLV2f5YPOiz6azUqZu
PsmCScowvtUp5nYPoj5oZtS3nanWo/LndPyQp6joXn230/jKWl+kXb0JR/JQu0K+
lGrxmtAqj0gMLwNEBFOEs8UnEI9ZF6SuQfvY4enQV8kNk+2dB6TpCxXPFnkCNOPz
neYt+NLWNsSzHFtTKwU775V1xheyxIdhriUo8FIyvvQSXLJnbqt4wZ9J68PReno9
Narnk87NB9YSDtH0FO2N+49mCrmZO2fAUh7gl+9tNNP4RirQY/Fdg5EZHzEtFSpr
oBLltaKyyeurrieTGS2vAUegylE7Z4dGsqMsZ8wcinCv5eD72EbtbBKE4T4fMw36
af1kp5fZb/5NRPDkU1JOVWRDWhnraQVKiILRAN9G3nFzZTXDcZaTscMlsOpg3pPZ
cW4KvV2u2AKifvm3xB71WjcWz/Rv6AqJ02B8Sbisrsd9xY0htZfeSS0jrFko2guA
I6CN/EIG9Mv+zzdLxe177e55R6JgHB87RK1PlN2YP49hGAFERya1J/zKyZp9Y3TR
qTjIFxvmiLq7gwAKA8LNM6Oso22AM9FGDmXuYYqWK1r0PzxDm9T2/N9jV6qUvMi6
kpQQT8FrKrzfu1c2LBGwt1BJYJey61QhX3dMRfxQktCk9Abg6fUQeNvQb8gK1bLj
kBMy/VOObEw4htpPJdp9wMGiyIHNmtDC+wPUYT+adjK/ctPUX7f54bC22MjXVyLc
JDPTPpNSoWjZgoaSOPQzS35A1EmgCCA/GEZJVIdH9G+oOcEs8dyy142uRWsHIH6G
AeFU81PGTKRAfCv/Tr3wKrFf4VeSdWKB+wNO/whrc5onbC/6ekpso/8m2m4R9jAo
zKrOmWly1NzMM6mKIml9w7xbltiTrem3OVnce68J9UOd2G3Ns1P6FbkLOl0r6asd
AVnVqr+Zesz454pW8ucqBsKtFLyuPmHkRRPRt4tnY+z84tP0ZwThcFrjORwLmzdo
41o4reoQosi+OWVTL1Palym7Rtcc+w7qFOkYe4fSlzcjAKPAUwNz/tWk42dnx//n
xQmUN9cfmTTVJ3aezWs5bWKiaD3+eGBUnI6KwriPT76wUFuIJTXB3Q9X8AscepTS
11R2QQ3eSJPZGUaeNesoAbtQEMfj8GGkxoH1eCw4a14q+YvpNIHmN8hPryRh2yiZ
9YyPZKWn5a4A1cQua9ClGkI2F1vhnaeAXaou7p6V9A1M+NzDc2bxentRTZji9vTQ
BjT6qEK8y1ucscIMYH/sVU/pOwa6E1wYk/so6/ce6SKVndSL/MdQATSMvl5DP+2r
yVNT/XLCjHjZIYh+OhfLZk0wXU7MI2kv+Xr/DSKpo8arZCO3NbZF/EVJ/Ucjelcr
QEln75kYZzabI/a1szxzL64+owVPXT+IN9plv2/BkK78BsHxFQg0hS/QwKBVCeB2
l43qfqUenXHP9fFjkYEbLApBhR1vs2XfnmUrzs+Z7GqzKftskDgJEozSGVNgf0OB
9kAD6bcWJtHhf+KNrFleUVVQsEW9XuZxFan36hXJpnMzrQbAo7XBHoCg9mn4nYnM
gRc5as1kecQDiNiyyvluB5ZQBA73JQrPHaEHvjOW7wU86/jXg6x6TYCfAeI26Ntb
5V8zxn+JV3r9ZHsIMoy3KhqXWdksQaOL9nJDjsHTxtlmJ3wfpZwwIHT7/QTfeYMb
MtpbbIPFsOrZVyi7WURqwCeJi3CTbzjG4wMIoRF3yNkSdQn1hmMF88hyLzbd1bZl
FW6/PxQOvSuoMn2IqnaGYwBPjizUtqcTZo5Clb2QS8cR3h6kTLnC54kCRUsXW/1X
MdNbqlGzBcdDC4Sm7wt4VQvMcDqQCUMOLUHGfPu01eIE0q6JlUfK+xp9bvHaulf3
eSqcKXY0I7+/w3RwjzT2XvKRwJI1Spe9vsfcVYVItcYmHW2tqisPIitsyvi82Qn8
viAWg5q5CS5vO+OG4JgsbYAhT5uKA4Eg6mcQqxal/vLL6dPJWQhk+gVkLJNp8Q17
rS0jN/uKgKbjVL+809jlIeajx9e44wmMIZj2oTngO0EwO84TTs1sfTYFcTbQvPpQ
j1E0td5NzmctQ64Wl85nta7XrQjItxRF/vx2IgSLhEOmfo6HNexd4YHYLfAkAFyY
Wnm0h+5TX281OdXvjD/jWu8jNT7jobOuwx2aHbzOKM1rMzhRotwXTyzf6aSYJZ4H
aoF+8d2vLYx+OxdhdxxRtMsZGfbl5rvU8aO1KRCvrzN22IxYVfWMwwPcDt6I43Cd
2R9UBd/Nt44/8Wqwhvlq0EhIFRc13fHY7onHvUTzBxPjb8DcS4w8NstxJXgZ5dT0
kG+3pcDRCISp4KLkzU0NbSgEKNzBWIBRA7ug913MB0xy48yu87ryEjll9cl93DSC
5QbdJNbuzdu8mlmEvLX1XnvMOBOhRw4zgrzKH5mZg/T/43t+/XG+i0qxwHnGEcL1
brgNBeyUYoNwIwlpEKp59foN1Fgh/GKR3dYqaCosYA1UuI7nKbGjHGLCkae5Ni5g
91GgVtuvVo6ec+EIv4Sl8CSA7NB5J8D3ulG6nIwc+NPZpZLI7o9S3ujz+c25VbOZ
fNpMZJiVXELN+mPjqBORoXs4XPKv1auEccuAJpY1bClFsZCCc6v+17ezG9td3w5q
0bO2DOFLH7dPwJgyMFzah09EKJId0zaCKzs2mG/aIlzv2wpZI/PfVrW31r6OuI1c
REhNnxGyz0IB+2rgZtAUQJZrPT3dUoBahj8yBQJ+rs5B8QILk8jrPczrzm0iLVN7
wckIaO+Xcizx1HU1WOD2vgHV81NQniRuVgMImj3wLFde2lLomoYvgrZKN4P5zRx4
lt65O53OWj+8yLcxu24/PVxO7XSpOIdlT2oU4rGbqQL8Jb5mZEG9NOLFpz4IoC1v
QP17auXwKe1ZGXgd5bl96L/IQP16u87/aafRWZ2a75CLbXsqkjElwYqShv00xd9C
v6RD56TeMrYYuLwRRn2J6b+EnulsgF/40wABPFQxL7vxlE80Fkm/NVYkjGQg7sXz
HEv83yUAoQQxFiFFJykCvtrBb1NfZ6MaUxLzz+iQyq8ggS/l5ILEnPu6X+v5I/6F
sAUz9C+JyVsaTjE5BIX0D3/6THh3v5S/oaO5539xssqyEjjNdCHhFOZWhXw1b6wu
yex2C2tzp6eid6vMwfWqA8nz+QJ0tHHodGKApqcDVP55GDWYjr7d2lC3+6NIZyH+
A5kkvQU+1MTtOLmsKF4Kf7ZMODmBV9CfjyduoiQ2dsKixwL5mSRwZnwI5+hBSLJs
kbha0XiDqM3IjV1wKBrPmevv8wJDVNjmkegYIK6vo7rnaW3gVNlkkD5HWBYRbQGU
V+gnotLV76d7XAPUuaDiOiX3cikJ/a8jmiPAziULx+u9SR+Ub8QZfjU1vzAsgDEl
6c8wTCCNcnXotNu8hZmUVQJsQhjErRH2F3PSlg/9pYO87sPXzvPgwbO/UfgEZDpB
UkZY+lkFKrcDbk/5khaNFCeL1NupiPnhOV/Rr+LL9jsevlDUqHHoOwZhnAsmG/aK
Idj0rXQ2ELy5VQfK+SDoTwssfSjyfcl0OsFfxKUtmoK2j8ukStuLC2kT4SJ3xZcU
Nqfdr+NA61aZFR9O9wnLWJxL+dcbfzVq+cRkQBJVPOgTRe61YpygtH8kn4qukIAM
rVIusMs72oXRS0emZftWAvG3DacKLWNfnCs6pHj4NPmuyYSSRKs8L0aCAm7nKQlJ
Ndkz+nvLWBukSbPg/VhLptOJbIxXHGXqF0PpA7wdX3GELZE89+5/ekYx6JzhslGd
4iGDWyNeCcDkQPGHXAC8XJnhKIAGVTOWXEiRRc6/7WSNUlRGNZP6ReO/9ynF7SK9
HS6lt1nJ7FgvNxwdYZ/Tp74PXICAsYnoumw3Y+CL73Rw47jq1P0DYcXMCD/G9SEU
UUZ9wmDxVALLFlZMIn2hYC01u0UGdCUEp2X4OqqzyHQA4TmtzdHa61g+KTiNeuRL
MIR0Q1FZLcRLaXE4P7R6VDE2DStm4MUcVu1WILnJSp/K/wgCfoygSN/c7m2nIzu7
5UsXFrg3Ymb95EwzOxVk/zC0g/psSp04FQ+yffsMIgYVbEymf+zPH8ZX65mXlpMe
A9Cf/C+du0Y+BR2HWq9yKqYF4MIWPn9Me8rSbVeMcEymwmONxRbd4+Hwe3wXoGQ1
BWcXut3ceOmH3dIg7K8Y/Ru2iIPii5VMk6vROCSeR8GZf0tmQHiPYI8MxbxKWW54
/J13b7c2tteInKsCziUZM7OCtNRHczov3eXpLgQMaX2JMwo04SkUy1CEL5nlsalw
ewOFSKLIUuKH44vjQsS4V646go8CoFbGFEtQmmjVfOtKzHG1+879HVM4dAIoaloe
6/Q/TUmigItVRhVWXDxcKHOF/pmXEspGx5JTVDY5i/33eDrBsBqm6hFCa+djRhAO
Rdc0Spqmp+cpuBWde+I+hNnVVLsFwwZmBZvb5eMGdUDi8mIc1doKaELwG3AArn++
FAqB8PTxvYb6NSbUugeigwsdBXARupGt+bQCHsMWrXpAFcgxGz1n4U5lJPzfHxNQ
94tW2so9OVXWN+npzND6sx5y+HYmE2hjPrFaqyBkGlYb7z0Gdn2rOcTyLC2jXVsN
FPeOhUC5abk8wiWLLLifUTA5mjbPE3UNEOu/X2IAN9f3BFNJZecmkPofbolWWbJO
Ss2JFOGRZokQVT2bSLOBv5fzu6VHWq0sh4h+q3H4EuJOu7KSD0SorGDxaZK1oFb/
y+nE9S32mXuo2eUMkydsATXVCKWD4W0hgVcMAPxD4jhuG9YAHzAJ01LpZWCnqeY+
L0vl4U657kgFPTRZrMdX85n2V+OI8j3ocl53XKsn6XcdW9XB8eYWmrT4Epx07WLc
WPJ4U+FCXBzkn9AFB3Ii4mJasK5d/dfMnf6NuyPjXLS+p2cc8GRDb/b4UFvwNTTM
RI04LdXmyDHHC51tMl22uuar6eG+7aC82zsGECuqs9Ck9yJBXHZYU7zLp4vO4gXL
4Hb6YCZi14+c7DHGAk6QgCl5Nk++dZj01HKBp3BID8TLOUjfoYYmbwruNFk6u+qY
yRjL/D1Evx2R0nm+V7Q2bI7zF6F/fMm6QGz2TxQE6Al5gq3dNGbZsIBsTwPBGLRn
DuuWeDkYiZrgzhS83bRA2l1FkMiRPaAHfUQAK61ZN0hpPi+2uTyg2IsFVMqMJEtJ
cq0N9DudJNGuE2vqUiAAFHA7Nw9xolBtc6YDwb42VSv2UjpU2i4a9vjyb9gfBeaL
JrkCKaoQuaZ2hWg0kmAF01uLFlJ1WVz3j/2DoXxDcYKwv3n5EUJtZZrF+Pyl2N3o
by6O5wM6byPU2vINup3MxJjwrOPbb3VEGPoDKgCv0g7hi0oAVA6LYNf4UBUK9Wc9
7G7T9ESRtOwNbzxMdj6Ek7qfwPVfp8C2yIB8EGuvLgz4jznqySH24lwYYH8qvfnj
wycRtHMfysTPl6tJ3F0+bNcasIeNL9miFXvKZOFfSKfelSJCbhYzEYvmO003Mtbe
Ne95oiLq1Y61RR/AkBZLXAqSR6yM9eG1a/TlThv0cdv4NsJJrlDwWXknS+mp5/M3
7ntwkcp0Hbfj3k9R9tH7WWFlM308+a0jusBccE9OqX+xp9kYuztzqVy8v8RgXFoC
K3eafpOoav7nZGD5pEPFlyphRJXQUK1L7McgU5JMq4dI2vdERFk2gqH87S6nOndx
DlkAWSuGvxex5jR7BxRbGB5d+ki5qSqU7N9HI1ihzZebGc67Q4v7Lim/6eGl9KJi
ZA4fn8hcKBgfEcBaRFl2MwW2FaVrvkawBN950QBIH7qCG3Rb5EZERqIrr7hd5fr0
h8roRBY4fpIb88WXqgdzqnghbKSV/O7GG+2E/CUxqATrEmNk6mxp7LQ13X3rxlQq
fGddxVuAfjDC2NmKYZ8bbK9Hnti/QS51XvTLcsGFnCmAC6PWA5yTUqMiYRvlK385
BwK/xdHln2/pA6ionVnRdr/WFeDMUxD3Y4lznDm+KpRc/YC5XVjjSopouZya2nJM
8n+/A/z6i/+aFlhA5I0pgrEPssdFuQshTFiPUdPQ7DQ6y6wgMvj2dQ/yvmfi2RdH
YJpTWWb3Ie7yKYWV0VgFgR1MnMQNE3vpmeuKrmkim+78fl8PIRp8TfpfGpsZKHjU
83CsKeoonTssInD+pB41PfeGqn7UhcV0xidw7EKy8amUjUQKYtLZX1JuR1yVyovq
e1zKXa45xihYtZp0TMHB1UumAvuvUbXetfSYL2wRhmQwVJKHdkFuIYKfE6Me1OzR
aqw+ZuqQBBzEbL+hvILBN6k5BtqO84lAKZ7PPJd4le/EiBbpSHHOa1kw5zAQs+cz
SAY8TEErxDip0aREgLndB/z6KBe65STVB8cukcJ6MxfpsOz3mFWGAESIqGSBNpRR
mjio4KMCanNZSi2w7fzXqdFa8d11QpakLjlaAFaRuTCh85ypwcuPqpRdIa/+MRnr
9x2Q3Q3eWx0bBDouDZT9ZMr97xf2ZS7ITMpl3KFuAU9nn+kJi+5Grh81bEDiPS7r
BD9lnaJ8shy5oQN+jPxsD7iHH17iRfSLUmUqsuJ78dMWzGI9OClzcg6UZgUdCHWu
NgeAtvicKWYiQAujgSh8mF3YNnGi3VLuijhanyhNg9mzWJHKS1MfOuXfXAHlc+ba
VGfUQbduwCj53acR6zfnqOJtIxSSRYW9mSq6aQc5lIZ/GHPH6a9MVhKZmdx09wnZ
th7bbemgB/2iuIm5J6WdvDuITE5AgjhZrK7iNYCNDQzdCkE4ZY4x7RWCDoQSacui
/JE7NydFdp/8pHB8/QHSgr8YZ0UExLYhLtpKdKh6xzPmsJx+p0TDTtc+ICXVVXb7
f2xEWXxTDhpctBTP4F/nKanzSpa9KZjUN5H3MH4JbX2RyQb6zq8eO1Tg9qPIQGm/
zjQxw+7LAPElBs0ncmKbuIcCqFMAT84DHAeUkXKSVxz0tmCrLN6vTzf7yUR5Mbk7
1HO+FhfGBl14zde8amzdiv1o23lFBvxUa8oWoRiebzR8wHEy1ibsjXM5uVGHFqMQ
TgNbgZHmt7RCoeYIMESHas+5+rfVvSnLxoZa/W7xXah7gJUQdQq1lbr6jqIXjnxW
HJux2ujUot2TtSwD7rDhexyhv4hLCAyY4Q7EVpqQ+j179loZRciJ/kLOq/5495V7
MqjRzFnBLn2NBQ02bnc993Sya+PLItzbUkUD+KyMKk0=

`pragma protect end_protected
