// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
vHuMofcT8UomPmwvgq9d9yCqvO1W46hDcqjuKaDqiCJ6X4s2jehmFePvoIMULkizJhHMNtW3Evvg
5dP+iLSfjWoOI50sPYtnvNdsVbcyFFEBBlp1NCRaQ6WxBmln9NfcpvUXAhdekJfLmli7x4j/rG4v
Rk2RLv9meSJxuJRomfrLnqYSij/ULPrCO5a0x96goV5WG0ntvRwD0VWhq2mEI10wDNfEhv8Afe5v
M02qYCNE62jta0jDmrXCM0bmdL6zEyoJJFA4Y5y7jDUP29lxaZhHi6/WUyEeXciTp6kqYDBgv+2n
lLt1q4EuQsB79ai92sOjeJb9dL84M/Y4CXKYKA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 8640)
Mk2D2eI22apW67iKS4qIfumdApGP+4mPO6FATC2kIeAxsfoOuOMe5EnY5bxF7/O7b2ESpUriWUFj
Y0lTnjBLEeBiOQAmcyS393BGsi5aWWBnxCCeT+2UzK8DsoHXDVx60M70ayGR20uZj9A+BJflmMCv
40x/dUMcC5toN+dHsdN3Mq2h41Fgs2U15y/K+eocgn4UXf5AmQa+yZUbbfbe7VxeodxumyQwvL1g
iZBSIbgXIhsjRv2iY78kE+ljyivLAkGg7rQk5NvOliis8kZS+JFPPcRnsvIW23+B1XfvsH344b4g
mhTOBZDbecH8bfHdWQ2u2tbApV7bND/ZFWcmZoU2e69qAufiAcjay0j81Ngttb5ex+mZiSlzIq8m
r1AWMN2jFvWn0angcXpMRzVwz877HCsbuWSAmt1fRZh0yb638L6Z3sTzwMgwkQlXw0JKytLG2VZD
ePL/7n1qHKb1/7AOV+0NO0LYRgqacDSFLVh/4rJur/h6uujcXX0BxKS0t1hjOP9EAzNDmJqk9t7F
A2zHgSZMN0WCrCuLFVIKktxgDxrGJM6cskCvVDHJyrqP56Gsd9cUQ1LHiwvPnrOYw5pYk+DHCNEs
sNJ+J+1L+zOeYecw8lX8fGE83B9eKVCnJFdJlSRNU5rZU4jn1FUySn9zImIq8Nwzxiue/iD/In2H
40G4L11d6vdsO3V3GhwTsIQocbpSWpKCyKKE6bL1WAgv3shO7ngwUyJbxn4tJjS06etmhKxKqYWk
NBaRr4Yf+U896dRizoi7mfvCqg+R+KGA1Ffzjd5x++Hz6FZAoKlV4Fv9O6KalQ7BVWrq3p1olFGq
UVEPkpAJkvKb0DzYpRFEenP7GuX0DXEZVBmiiLmIg6SMDrjNPG0TMdF9zVKwa27O8ns/K00yftsC
9/j22ba+3V2m85Py9Zo+U+iFxQHZoxICVOoZ6+rf7lYnDzVPbSEIF7VSkymHE0ve83lQlamNQBtY
iKS3q7BA2cxO0nNDqy4ARddUUu0FZ0OxQrmX/bPYMOvPn631cPZcfe0gG+EmXLg4hZs+Jn195RU2
xdTUnNJKywaLEgocMh1NOwKPmf1+wpWd3rhnWpwtJ2wMZhOB+MPw8XAdSuJN/9yj7XH2FIxq7jKv
HjCgkxNRSmg8tsLPFa7G86GnJvprNMWHm4XF2oL/o0DsHvyQY9+xoHSG1MwAuVHL9OZttMy6TFyw
PFtuxZkU1I7H+m9xn/kMvRSVacifOgc1P3gIatN6bt9fBrW41ukX8oTJ9q3I1lSMiiiICzcJqTH0
avggbskmy6sTcMh+6ShhFhrCu3MbITpF0GPXm/vw4oGCIy6J/zqikaoIPhvxXgWR7K6vypQYr8Gg
VxM/eqgB8qrSqaYUVKGeVJxqiqCrEeVjTe8ep4BQ99MJC0nX4HeBoWGto5IxhnPTb59O/N+qPkTw
vkWfUHR8rpIknMHVrlxCK8mSRDZQDJjt5rHWFXy4RI/c9QZvQIyLHI0DPdLs8CpplNbMtZjlOpJv
TG2zOOUYUCsTdITE73yc+7pss3LeYzRj9hNwWUpwFZazGPMhgGR+Yy4XJ0DgVe5GxNJORfa7ALPB
bmWN2nFx0njs5o6uw4BjZBTSwueOw5ZWf3W7dRwFFI5yxnmAnB5yc9S4d5AQn6B304qHfpFCwlXn
2U0O6VpeBEXbaF/S6fgbEr70wyaifL3pVTGSNHKqGvA1V3CYuytOyZmQ/1crtj7K0LnuAmDpOoUy
28IavaW9Rkw1D657p1anHo/wEwiMPOBBW+VIA6+Zr39E5Ot53N373Ks8DHqrXlymL15tmvawobPY
nQJ2+sKWECspWRMw11PfPwzdfQdxlVoVDuEvXsM6uGZviG7W+uhw5coSZDR87PAuDEeqCHu9JojZ
F/4iwqx2lsOOCoMe7xNVFksbba/ExdL7OTfnJCAHjJfmkvqbwOgZRFJ/UHLoI705+3ukcKJHYb++
Fv1D9YFwgizCrurUU8wGMfw0um/yIZsJIFYBuqiuLlNKc/tUIEtzVVa1Jz0FfpzmeWVQmJQex8jH
ahlZkoB6M0BmDqPBPxrHtz2oDlSiVXscoPjCQsnUfUdiVJqhnwiVc+/DPxjvPsXAF4PwTGUGucQa
EoFZRANfDQtIOM9lFuXD9eUPfVNGwKhzaWQi0CfwqDz4Cx5Y+ZtlLVhM5xARP3L6JuBoO20jcpvj
Cr2TuODhjm5vmcoq/a21QmW0/E+4yf+wQB8iK2T6eJy6MFGGcPObM6Fc8M4RgsDYEN86RigTfz70
z+G9KY7MhkROr5SjQIlIO4zH9IQNQa10ZJsXOBX5cgUfFFJBkKomDlx0HKfIRJGPhkXesR1PvBQa
EIjLKW/w0feBK78+fGgtcgIC6xqnMJN7DoXdWr3S8d92Ur51dXPhjo/iDWj73me6sCCicKinOrrL
7ALlcqIbI8H+Sh60nSsVaF72ugLGNkRoD07ySNhXLvzFtE3uqajd8vFmG/0XbGP24+YmQQ5oAys+
Ttl8bg7+io2ns/jpx3Wdxff7wzVOJwYqPEOOQ88xlDWRoEoF6h1/GC3vZPmjn8pyUs1M3l2iyEOn
1a/DoDwVYMmOjB0aREswkKipz9khKFBhbIo6AbUDuW4fQrzsoQAZ8D5PD4IoYlbycQppFmaAodC0
bemgKU5MtKShaOG1cHStUJIDGuKjj98NfJrQv/p4twNf5iMKeimT0Qz0yKJpCcQnSbA9cDWEPe4c
08rcTBfNkN8aIoLT5v1cVrLR3OoeAXu0yQ1h6axxX3HpGY57KRglmN4kyJvfmG/6drU+eaT9JuY9
BprbVnt/BbmuM7RlcDfHt222BBN7IaiCyGFiC7x7O4zMoQREhToPMuFedttxmBJR03od8XPZl3Ha
DWzc0g7t/xLLPqK07JV6Z5NyWQVsLfvQMOE7mPARtHw+fLF/BOi+36g3h4pfOZV/p2KptwpYSev1
Dp5hvC8pMNR8AVCXt5q+ZFmEmlHT0WczY4ywoa8snQ5JxNw3/gAVx/fobL/Ypx6NNrCuSTF9naYf
u9WKIu6VAkLBybqOIJ5oLhBRpT0n3vYg3q5dpy7mlqxvGV5WpX5aVlRzCTz7e49TvzWeOJ9X6Ra5
1fSm3aasw9BpkkqdmHD178mrO3QZh2pd88aWme/w0PSj77gAtUFBg3gaSSZb3y/91Kfkitp2No8l
XqCBCkqscqBvK0s5gb1vEC772ZwVil+5AbeP96ZpU9IhUuAZblpUhic5Vx5Mphco9jGn8va7oGbO
yNUISF+Gjh0REeOygJap8EPuOXyAt5eBI4CFc+sQla0hDCHDN3VUhrRtS/lCrK0zsXQ0HpFr7p07
w3mhICVHLk646pelS1BAWmfSHgVGuGlcxvTwSD6HGbOlnVm6f/gqBBA3JLvk1JgitE2nzesE2Qzs
zWTxa12IjO3EKyCzmrsseYJCXV89L7cxGmOABw3LuStxvlDVx1B4GCe+DlbedE1ZAMFzkBUX+FW5
yIc7KeMhfyKZZQanTewLwICmI4WBpLog4rpcfQ5qo2aoXmSi7xfGlquj7Od6tFpwQkpu49rbxpVu
vUVJU2wxIR2+6nqMBsRnlThaFW48Dso210du12zSSSgF58vFTsdb7O892qw6imF88LKaETHhhIXm
Es7xlEKHhUIkvMj5y3TEMsYGpDgGIBYw+fIIhncUFQXt2fARBAZakniK5e9e9lOFIRwNa1SMNT9n
85wWneFa51bTB/FYopb86fyyrXwt8qN+0maJeujhjzcCFAw4FOlIpQRWABeLx/l/GHSLf+1ZsMPE
CacFuNgLsSouqlnhg54iT9y/K7gBMbKjpce2bVR/UonEOLnqrGcqjn6dOKnfxhxUgjz9+/0P18YW
7tFxFgqyVgbwuIOTNfrYvVch6c+d4L+2KRuO+f8tTxJCbwWoiEZGrkUBG0KKJg95QOkoL3ybbkBl
AT5H+EA1fNgKdZ6kkkvQ3SR1styZDPueptDSIYqV6dLT18Th559eVAY6sM8qSx1RU2mwoTc0pbno
BJoXjqibHhw0g+EUQs8WPrGT6pYX9bJTy4PGRmyVm3GcPZMd5ewIB0xnkIzLbw7ErSNOKC2S6Tng
07DDPf3XRxXJDUEX/FZ778Z/JUQqru9RuV/WvleaBpTN7Vhfe9qXzh6+KdVOKvIi3HdGyB6YATl/
TdINZj2tfvhZjsSOJRI4yfHMZDgOsK1JlQNXF+lm9ycNFamRcOJQOGblFi/1RBwbcqeBnYwQbfEY
7BYERpDbqSryw8EtzSKmMPJljNxiFq6v3GAz0RE3j7tYug3dKnSetw5jjtq/an9un+r74z16/h6v
/MRL5xx2UF1vEnjgrlPAB4+a8isZKzo6dLMnLCU2EDYZASs9GofOE9l+WEkn/aHkbDylClYtbXep
NrTHrl3MyOB7gLrw0aTKuFEd0+x5viG6pfCRXvuA48Ks0SJlemh6c6vNcvcR811veXIHhAzkxx9S
CO9JHuSx6uJ164zNmx8cY+ftW3lGT0OloQnZ6KWP6WZDpesSNnbdHyTR+v+A3gnDXII2DYNzrKvM
HQilN7rN/6xBUzbc+9t+kQz7pxNawoKseTKEsbav0Ap4byhgh4cJ39XBYHS4ZI9BvabLyq5+rsLy
a3vDatSgfqojCcisgAH+K66hGDt5UM3mkeWBJcgDt1hr52oOGf/4n4GG1c1+ODD54aJaIAPVOHm8
vayAy3TOj+2w8aSrCChAh3laYArJDFq5+vK7BJArBHMmUP00D3H0ptc6Ev81nv3oc7mW5VShhQDt
Js6uiUCBBY0yOKEntPyeJarDrAK3ut2dMaw4cBOmHrqay5KigS5cwYsCAFGO2CLjGyt/r9lBrhGY
pitBer4EUHvV1JZoQRF4joWcPi0un8wXrC1gaBOquVxJJEv9t45SEQ+OExnmnbgbVCsu4ED41aCj
apePCH59PqyBKe7mjry9crs6Z9IdiKsqMbCCtLlNun2FPdS6tuPKObQ4d3tsMMF0MacV93wvLRgL
dd1O2u4KTeZz81MDvjekgT9XSJi2fCg5sDSXIWrbwgNyM9HoKgEC5OuTO/lAEP8nYYG+5EXIXbif
Mul28duumMHXcyYTe/LCMZ7efrxO0bX1ekqsEtNSuU5akiks1q1OBvoc2NqpBJC5P2KISpuuW63/
FV0wXs1xtqU56D5fsWLeZe65fdtbNJohzeohjPJpwb+h8DNrbkDW9TWXb3ppXOKCPrGnetaTT25p
S+sQCBq2k4WqJ1RwHUbdaFbDpJUFnFoJobIWUzuIU78bhjphSZUkKA/QOukQbDtHJgLLwgQWiG5Z
z2IFneiI0QFWWPk0betmSMthGCKurj2IWHDfUY6hCXmI8cYlRd0gHGkZghCGefBP3M/Q8JPC2dvV
5DZkd21Iv5vDE3XLbmq0Km/8xzRCz4JwjKE6aXN762tagZkDj+RKi/g/PTuZV80F5yCqz96k2CRd
Pb3k+lNhzNySrQex990LU4J64ablf8hJRVAwiJDbOfK+05vzJ1IeWWnVXUFytJ4pFWqbxe0MwNyk
SH0i9Err8B3DCHhUtverodgSbVzxA/b9lEZ5MoUGsoRPvw2ATOQUod+fBv/hXE/OzGCGnwv4mxfU
8Bkqo50FucyZAwJwlWW4WU4z/cM/4ddB4exl4t4vblZwniouhJXSmj0saYVI7+OKhFCiEcWyR4fE
1JqXT9jiNWJs7zd3gPkc5FODaIC6S/KROvzIC2Zff8604/q1orCJHxrztEwQ5GubMEE7WUe+hQ3h
24MZFk2kQGIuX6MfgxMAtIeQg694XHBHwN/W2pHKfuFBFLIvNq9ugXoj+wuu/T8od4vkv0iIlLZ7
+oKsiVSDpkeZxuwqioGbYgcytIAtr9m5VocLLtKe9iK+tGAPAdV/+m5125s+FuW2doeXnSTiQygS
gcfXWBveBeklsYyJT95P5CN1IyQ7kyX51fgmMA1TzdNaL6SQvxunl6qfE8ZxXLonTOWw5cmh2yTT
eimCj2taPdQNWVo+w2CMMOI7THqe4CM5bWfYCMnHQIAFkbHwFFteZz+Ywe4FuYorjOITdLpd9suU
Ed1tVaIXwCXiK4XiekEikMcd8ieYIaccd6fL7PcQAxoyGAa4hciQMbu6CCtLVopj2k110kLNiJgt
Qag3Jgn2VPCLsCNaNZsjjoQh3Asft/TTlKVzvBqG5hqZrCvk1N8SBHe0lQvLDkq+zyb7GhOISqMY
QM/SDOTGT8A+2dEfCSOUqWHYS36yUuXwyNEIGLdUGNRLUCXl2/DvjsM0O7Y0sru9k1gftjT6GqFk
GgIhO4WNHthdEjpDgqP14xVJE5rEiR1XajtNBShD1RiuY7ym02aldXSOE0NEWGm2yhkKYi2j3CaD
02urEUFzpJ3DR0kG2Pjg4CXUavNFP0JSZm8YDeYqXiiCDhftligoBD5cbIjmHEpnQ1UavXQ+ZZlE
Ude51GLR6MjhxUZMehwp36ATT5fDkBMhDgpK0Btc8D3iDIRIW440SfrmGxfvinoaBRSqYaC1YvA7
VRrmjmyx5WK+7Q/i/xDEAU5BieHmVZR9aQKb+yFlxiuhmCvUBRvePNq053xk+QZ0VMyzmk3jsDHs
M7+MyMSeGpd+yRETvHm15PM7kx9nPd4O0/ljHtdGxBTXp6gLCb3HvQ9JwGxfHEswzM4khHnqf/ma
j+tTlPEuaEdKW8FgHzRP7FkfUvVluP+HAH1DZ++X8/M1GAA7dqTeRFT0sQyV5ksV485xxLMgY2y/
sv3xhtws0zg+voxol5BUGMIXwFIrH7Ct6PE8Okh8AX2cqlmN0PK3+CiDXCLmYE1RVvOJ72Lzwp1i
UpVQ+MzwaC9vvmnK7vbVTopjUJ9oUVtURlVDEhRwVvlzqEkC7i7zUw2m9deG9VNzOm8WXomgaxIZ
Z4jok1Vr9QNAG2w5uE87WHaUyLjxPaSbVwATs3QFqFhRPsiblSTOgsUh2WYgpeVUwg+3AzNjOxdV
YNinGxIIvMZGq7XpkpsBuqs9U3Pp7zdlDYHbMC9Ju+zumfiktgWXuwE4Y8Hf/Qzsy9GEZvQHzD/1
QZGfTHTLTwClhmglT+Rd8zR9cTd+tu1gu4t0UMKLKA50e8gXOj7OOEw5izF+jzVWHkFXZezfrZwb
hW5doFKtAhz1gLZ9nzqhZiIbX0FpMBihU2GcBFvoNBDP0j7BFrNEYQsMDoOcTjM7zRxHyRzzCA6y
eaHnFtwqXVKYe3vDeEaYYu4td+TF37Pv8GY3aE4fjrir7sQ5mjvrWyB/z55VZEMPqp2C5S7eUTg5
FlEmPM7J2UFR7rE+lU1tO3SypBisLYQLYFgm+lbBz2OIvVyRoRlXOirP8V4CBe0k8upsnnho1xf3
t5Hj5qwKmbdlgvrDA/pFnDqlGNMMuPWRz+uISvQbYDFguyMBHQV3LBk+iuGpIQCqwvDZIR8L6BDy
TcTVylvVCRLWaMOMF4r/Xgp17lUha4kC8xQ/cEvOUccEzF4LdLq5SJJ2/rXcTC53SqscO0b3OzMR
q4onX7vvyj0JGVoUAddtDNrJQob1nLRa7rS7Dl7QroWPsJxHvXiZoBK9Ac6US7MG9c6zYvI8yllH
NfNHlPxJEcrnv50M4kNTi3CFrv5ndvViBwxlEkvGB/SRyjMMRT30CqE9+lfGZVp0T0Tg4i3zWJwy
U98AHyZReCPruLrvnevusr7Sf25TXtZp0vCPysAzNDyKSPF+Bf6Teom6qGh87m/duZSLMC+BYThg
YE2sTiK3HHyrj+pmHRtHTD4STkviG8KGERYgC5iU9YbK97V6jnRJb5wZegHBp+aI9jgw9hG0sH65
L/KKux8dxC1caNsViIDyEv+v+pLGP2iSuZ/Gw0LJcHjy+kQ4Lv0lxRBLf7lf2Lzt/cWS/sbxB+AD
SspMDWrqdLR28acCTwPBmC25KJDPf9INblSS8CMCEOQX0Jp2xw9mfQA6wqt9t9p+5rwR64mQ2iTO
vcjxnAGLzxhIByS0Vp9IesiLOoppJbBc4TR457sG4CMkqCsJU3QX5JIVeBwNyTvX0EUSwvvfUKlh
yxKXTeMwG8egxYkHQpumk9A7Wet5Mig6ZxcwWmnMHpMqrUynd0CJt7CUNeEO4VFBHy9ibH+gYnez
tdYqJrNHyJpR8vZyv1oetzgWG0EzWRicpqcLi0EXsxiD/bQjUqrxlXvcLpMkb++UnfD3Xs72bxH/
np/0IK999gSmdbQxoQoq/vhoYBVw/fbcocj32CLK27MxGbEch9Sjk8+mCEtd7EhPGgi3qld/RmhO
YOBmURPGJNJ3C+5IA1mtmC/VODCeKariplESZM8VN1dUjc3H0mM7eurXaH9NLZ4b07ErikKmz24T
Fjxb0svZ0I2K4Z2vri0XDtQmPWHtS8z0OVCSaPa4/hKaolQeP338krJ6JpbAN5uX4+LKz4io/mS3
mOf48h7XG1nwb5zQCUejtm3n1fq1lHI+QpDrYzFYO2N7OSOmuOdEd/JorVYlZSsFhT/cI2BtLzTJ
yyu9CHLizh6hbb/J/a3Rnprod4jujUpqU+RKhvmiZxICv0w4yAX4TW32/LkZ4zlEh8pROWBb6EwR
qJJT1wsacScGFIrGfiIhExg6KI88RppomeiLuy6/V5SaDKab8hFPYP0t5aRMuh18biH6hwGYNiXg
h0ZBHQPlQU+112EMvOOe6MjlLiLdFjBhB5bXLnOiT2M/kNhBNU4YUTWR++Pwunl/HOpjvRphNG63
kiF2cDwu9Ju8cpWp9oM4EhZ3GA27tu4IL/SKru5f7l8w4/3cKV1U7JhjnQhz7TOciIX8lJfCIIqD
oR87WcfpM6PGGOugXxlhJKYXCt/+ED5Uy8u8FCFKFWLzIVJ3GXmZriUz4Bzq6DAf5hQUgXCKTHOH
S7j4M6yXCRmcC4btJdkYNzAAGrxQDRqr3GREa2mIh54NoiwxEqCOP/+6RT8Cn12Lm8bw57zyKWqs
LM83slK0K2dsztm3ItW/qtZ5BSidwpSd0Is4yZ2QvCso/gqrTP+mj0IjAjcSzI56lNtM/UVpjhzd
w7W1vVofjKPGWPez8i9+Z4cDzDyU1vO6hk8kdu9MSKWVzQmePleQXszdqKZc7bzq6bnq8N/srpAI
eaejSqFCCc1QzBiMMhCnTG2YrTiFEcWeqT9EMSt1lCoeCCkf2ESUNmhvseacaAYS3Kk3KBUbbGxS
yX1zpmt6elIo5PtZzGmdpG2+t95vTg+Tqhl8b3/iT94K8KrTpia0SYFe5IPJGAcsvShmH1CP+ahE
jMZ69VnaSRN+Kzin8Ipe0OUsgJH5W5fLHg1TmsHvUn4xSv8LE06W8gw1aDiuhlpFkUpsOp4x4osK
KnKUluyNpSKLFUjIPVfxFRU0T2lfwokEI9kuLPtoN6Wf9wffyhFvydszWovcTa/YdiRTEyvQTghx
PMy1zy4e2SCrk2/PJnqBXl66+wviEtFrdcMylmrayU36SDBOX6ZC7cwf+6T10ikcqJeafRIQvraR
Bi85v/Yand9xwKvBoloY5qCZ0esTB1JQ/4aQD17Am9aOJESFq6TD5bJc2JjdQtZ0lrzakPgXQeGv
1qebPuBDworXXm0fWkz9Md590U/WfE+0g5I6Zm3Tjc8ioIFiCPQUWDN7vJ81HT46K5c3EB27Ryth
HwhCerTDuzoL6v17Av3zSammdV5vAfsYIlkb4ayAdqC2EHV5KPFXKIh07rda5scfFAJ4bkrkelLY
GsNjPhPbD9bvJnB9x8HSRnx9clMMOtq6lRzt8wloytdH34Gcvy25LD25drjd4HXZ3DfBwUMTPxc4
rtUthF1JQs7TuENZCKg/WSEeF4+X2drqhffa9nmOxF/a4oUD6xRngIF4EPBS5EjAD973TAz4ey23
MBo70av7KiNB/64YVJUK4KBGOTRcVxNz3I/U+NtHL7ecymPJEcq8N05yyf1Bv6y8rLTDbR4osKRD
+u8tQ9qu0vU7HoghqBnP+nbPU/uDaDtyAxhBRAsEQ/C02zuX/dnHt8EXC8o4CH/MODABaFUWjUp8
Fo+n+xcjG7B5w3kFHKniP0WebBqqyg02NLSPt7RAPnkXiAjJFZgoW1mmx4vWq4UezzzS/l6TIW/W
jdYUJ565sj5jxqwvT8BsbFsf8KVt+9oh4vn2VW0Gf9lNhGiArDaXFSrohP9Rl4zeD9qJ77CTUpT7
b2dMbn7t8pfGR8dcQCidjVZvQu4IaSGy5YvPEP5cnIx2WhLxBPrc8gRdeo/UTkK384CsKLzoc7Qu
phUf5VOOPzNeRE/trdErXD4ng4GWcfFLqAPJOu4PCOvThuszdfFnqyHfgnfUgtJwpi9CjPiyoFpE
yhvXz1F8okDh6YoDv3E7B9qka7wARKUlZHedyiOrdXa7ysqp5uPsRwlJ/8xZp43JOhyJGWsD+74K
iJLC+wYVQ8WZtliVOKmpR+Amogx4PuNGr9z1smmj0o1DD2cRt7NmGqlkWFr4cp7dAUYdqGIUWEuE
ojcQR+PtpiAM8sv2CUhv1fjmhlOSOrF0NGXlNA8HwWf0oUgliru1v2ulbmh2scljLFU7ZDnQ+NTI
pnHFGHirnOqD9EmtrpTkCzva+aWHQBcZLaq1j9RU83M+apVafyQxCiFIwzzPKGUo16ed/rhaAzpy
Yj2oxQA3P/YKpb9YBGDzgdQYrPqFzHwac6N+M7PQ+DaKwpC2HRqTZo5U88gky+T908icUg0ze8No
+WyEA30CUPkSDuH8VzXpJcE45RpqLzHB4+ZL86DRJ5R1Bf839Ff2NEcrCBN9xgE5O5i2DfD/UIs4
OZtMmOO5epoYXuRW9Tyr9xT801Gm43xuntaHVnDktdHT41d3CTdKSa7qYPYp8psbBzwD9mzpwaYh
CDmm+6ervSCDpmU2WG3R1G+OVzHO4QCJ7UeheIid2Y35KelAy0ol+yBxPpr+zQjkIy+yIFiNBYSL
RyX/MPlZ/4pw1JUPYYKFZVDZh0sxYPv0R4ypR00HBsnSMxk+pZFGyLty+1LmHH8wgZEesSANzU7c
lSN3d8oHCu65IQvjVRYkRerOgFUQ+YceROMcvIB/uKTwJaIA1QYDjie4hYkEo/DvxYpUr8qDayxN
VssdXfYXPrye9KftHr1GNjXZch1dlcfD04HhosoruMCFYFBk/8/wVTkLKJWo+YUeKOgL05pxEh52
ugnY+O0mWxVENm0v/7+V/n6EY+LSlDSJ4/03vVSLUde0IhnNudDFyMmOPwGf7YBJ6S7IOm2jumw8
RUr+z6yprJFPv39QOfp9rnVu/N3zHW3coorUleNkRbxyhi671tEtm9eotKIWTg76zYg9RCaXK+Yf
IPLHYfoG3Xi/TYTWtW9ktRDxZ5ro+ocb/5S3JS2cr8P3gbUGpdQwJ4ADgYLMULS/TcMLgnl6cVNX
M7Sh69PBL/1myDOmas/p5oqQ2NaIrcZJkL41C4jc9tlOsAHdiX2RJVUkX+69VjjHWi0+USf3ElVN
Ea7CNi9PfoM+5iwjQ2OGT3qjSRkpgEOuYEVdWBJDDeuM
`pragma protect end_protected
