// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
TRf/aUsYuxkNGmpl7CPE/gUBwlQW/sk+AiVAewnCX+AXD8zpY9HR3TyQDX07O6+9L4dE5Z5zLsP6
Hv+of2csFBTwTMU9ee4kaCRFnkhL4QROWE1i2OnODHtiX9+WDq9b6JIngcwjK9lz1cjxdSoas3Qd
kFNA7Rym4ZpfgbJKpDHxucgHjozNevjhDHrgzY1CRz3YckkCBYdCPWl4VDzu5kUqq7DtTY2Ap+3M
tRxf771dMygeVdhh/qPMxjXCaufAt8k0J+O4N74qje5d9xgniIhCXlM1LgYRj+1xGpS5xTcnehhK
XE/AqcLirDI79s6RcPZc8yPNln1a/SSt+Y1rNQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 8496)
OkE2ULh/+V7Ls1trUXME3slku8ImznShZHHGVHYZ6NFe+z4cj1Nbq6x71iLidxEXXR63a8lwBCc2
PJ6KdClUaHzZW+OVu53wKwQmYwmUDDQ8SXjdrpIXT2k9Dp4civHohjbyoJhnHHlJE4nvSNHvpGGg
Zg1/AhuUzZmwwkCEoNYKvyRgK+Y43rebUxJFzcPgi45zmXFVVxDoBRuvZ3v8GffQBgM04c9uvdPD
5D1hpSrKuBEyaRtr36Hvki03h6uP/+X1chBt8KWr15LmLyFfVQK+KVUvzrG92BTAd8WjtrI9lm0H
1Cmtvf/Pw+ryRO+q2bdSskrk5rBVbOAc/NA3Nn29bQNzJd97OAF4Pp5QHLAlpekXiJXA5MPcMHMD
+RNUq1Ygr7umh2yuxYZMAnGl1xrnOedG5/g/bvl3+mKTy44z8gdaPa/vWWAvN0C2SmnUwRz+8M+5
MkBr6dNp1mM8OmqR2i96jZ5MK4QZEiCT0Q/Hv1mjvvXyQ+nfM4bXDTZ4gfxZzbS8awCpORVkigcH
Nmkfyu0fmBJoApJS3bq5Ww0jfco3Dar1a+ZQMOfyMKZFgGjrYUDR+4MWwWGSi3ZtFwolJm5jOC4x
saz7iBFABuCKrWq7QgLbI14+FXUtLiJ3vgVQ07hUiLxplzNC84uJSzkMfk2pxOWBzcAlwtk25eXg
D/VyI0Q07kNfA//VAVMPJ6LsANq/h/uRQHMZFc0cgtt4bHdO1weYn6XY+AVUiEqdn1/OyboxERt6
fUCVcQdmSEBTeYPpnm5g7T8fIIozAUvyyfHT2O28WuA8zwUvz2QB9jXeP+ruwTMlCiTEEoo83CxJ
cqH36hrXoB2DchIzLmDyHxNgQHXLWhu433I5H9AQ8m4z0qB/MjqlJDKOK111Y1nMt9wLwKiJgjpk
xI5YrCxms447q/GDwYJbXRqOyfK+gEHGCn5ktWsJib1F38cTHYfqUVyJiouJmMTmYDJQwZYdrQDh
xom+TaYuJi8EONmVMwdNrYwf9x3S5nhd2eDPKw+s/bp3oz67gHZMK9a8agQplAb5RHsWCgSHYeSt
ByH5qVAKkAB49N/3bwnsy9kjLVorSAAxkPIGPaWZ9THvklD4pUN8nCdDsV3jfPW9DScQsEaayfex
9wxiD8G4x8TsXTAHk3bjfaWlyn+ZpDhibS+btFgyy82U2hY3x9t04GgHbVeS0ZDgO+3h3mnfunZp
M5nJrw1YUh+BZEuAorRjm8gU7aqv6BHw/2VgyeIIves7LsaZlJGTd/vcJ29/E0BBGErjIBkqgCMk
T5r2YVp7liw78W0Q1MCKkU/STnD75n+/aodvkaHSOuylb93kNv8OCA4yU9X5ThB6PXJYK7bAQDUK
fMW4HlU6+OKAYYyQp8RSKdaY2V+TNg7eEZmxMa0W5Vss3PEXMkVfMrcxguAL8j0PGhuOszmZyCk7
velIfT8GlIeeQTRkAtJpT8mj60sGvjpZnDaaVb3B+8qY8VMDqT4Ct2nTCdtYlbub0eHpveGXcMiL
gNDZQgaqSXEFVZUT3MIOYtUxAGrm/BlJSQPwDPCGTaj8IiafgWfhRYYMTdx7QGd/B5bZAQPwqQ5r
IvRR0/EiRAYLPlbJCcM5+ZDthubKKcXfge8OjwQ/ZL6WYuURiF99MUfbaZUD6eU4Xs6hAcNd8ECs
BSCp7n24yh5q5E4kluyV45z/pb9FU+nriUufjGQ/iq/+Cjv8U2j0fnoAFm8u80HT/tmugAVGHFMt
EhXGLtcDix77oQlzmuFdYsn4rfcnhoNXCMUb3wTNyrELD1Qug7iNFlfINAyfQRvKpDZqr/PEF7eV
0ROQoSS6x8kF2kxTD97PZylPIgVs16Bbdj854/BcW51/P4xMg7kdPSiyRXn/Aq7UWB9wnEwsfvnd
f5gIk4KQY18GqVWynlmcT1+dOSltHDTE91DoRaRSTpmyw2wcO4ohlVNUO0wKQhgyC10aWAySr7y7
4TsWqVsTa1f+yv1yDGtRYUjkUH5jg0Pr9mXRw1r4brxyh/unHm97Qvpv6na1SQShEsS5qKB+xvY3
ATppibii4Mq7+u9iKkOhURmGl2OTGJeNLOE601wtYNIPUIzQYh/ohIv+O1WhkxhCC7qWcjcw9sHV
FklHEDykW2Tp7YDMQZv2FzGlcMb6EmsS3R4YSdmJi1Zwc6wl2ohpQssDXf2hOGaScvCJhvJFT7vQ
u7L38gQnX8VqauU3uTXVZYIUIw3LvbBGYmzjxzyS/oMWWRDFnJ7oA6Ua/SjiXJ8JYWOkZ8Yhiju7
773Gl16sZvd0f6RQs0mX1ylIxioCi7/GbXHRtaIWm4mVeGDXn8zJAvj0aVlZAFPRF+mfNiEaXDXO
7tzS0lntyq0I+9Iy0I2AGxfL19mlEIvnhzEZ352rxd1gBoVG9Tw9wQaFTanAyPYpc+Hl0bRB0F1n
SL7AdN6bg2zYWYHAgIkFTFYsVVS0U+yAAGO9hfxujAHHSktx0eHIFxdf6u1L1RkUb8IfpEz55x/I
2Z2pq9TcO2SgxAvfUU0yQjMYS3LbnqTqEQ6JdrPccKlw+vM1pLpcLGDX6mYewDiKPZTS4oOV+43B
O6b6oNLUkpCzqXKQE4BbPf0KzCpbPbw0dHMKenpdAu4nnGAVBK7++4+rHBdyrZeF47otve9EFS6e
xPPJTwyWnJ2IsmTCBlaw7yB9pj1D0o/uDVUcB+CnpluRUSZShzivIimlguSo4Ncwb/0w2Kv4gNUK
pu2oMBLtL4B8s6ZgkrKXxuySNNFoDQni/4UScIquyM84VQifCGokiO1nHh/XZneFnQYxmYOY9O1U
i9FvvKagPJJ9h+HoMaqkpNtGmoUCvQMO/jQENbmL3pfvFSf5z5hMCeHVbk1Gy+NR+MN4HrBiHaE9
2nWICNsjv8P+Yoox6TNkBSCFd6TOl6iOgakp9/xEOtQu7scQismoqO3azVnEDjP8UaszlMnNOvKJ
UoGxiiC6BxE47lQXO8kSeYbNlvcfHXRlbyxWnmKBeixRb6HwKwPaFeaq4zzPyMV0JXKvENQcGMEM
Dw5N1yB91nL+2UIPt9JbuHIGUKQ6HzweyEnoVqt6Zivl2AyEES86DjB8B2ahqS8/NDtT4ht2kJHv
MvXNBDgHUBY9g/RxMy5KaZA4O2NdhVuRhTt6N3vYe39ROjKRSvWlB2Fi5/jgYv2CYvcv6IphOcbK
S+8rZ8QGnpgH2eJqW/LmzV6JOwK55P/VCoJZlYN9aLvPderxKBqrFa/u4dFQLJbFhIKWdnhaenCX
VAQEyWXP+wQhTiW6aCM46VkQT92nuWv2XslxN3aaTI5v1I9cjn3zRYnZ5aEuUHyfO0Rb4NmnnnRl
Sja1gCbzkKsOGGZV8JAZVlmc1UoBclWXcYgp+4QdU4MVSHexLFpkry76hS/54jM8calbzIdUncLS
h1qbvh+3gjNY6ElMs9NdhKD0WJowqvFJGoo0jIhLiT4oBMgmmesmSUEePbjobPRS0gF6bu6wO6dc
wZ6wMRi4+C8A2bt9WepniIjOQGRDGvgtk9xR8dFk/Mk3lOnr9MjuWvDld8zKoTU0PGHFoc5VZK+o
D6sYVmQWqcRESUwZXGq6dDcJ71Wj8fVbA9XBxgdM6qKV4PszuIiyUV2+jBWMLOhgll7aglk4MmAB
FodK2p2NvZMXtChGezmwNLB86xXkMgMuGSBkvFXYWHARFyVHMfRZ8+OSWe3UEWaBq4aKuqm7rHZA
Z+HUHgglaJgv1R8m+LjHAL4xUwjcmyKApy6hf3YLpSsnqSNmK8G3McKpvaCCeBAt5/uDkwdTZWCO
HOM5CsyUoVVRoX3su7yt+UjtWXDVVLDC9vStXynhFMIvB4O3ut08k8JdXHC4Gh1Wngl4jJ/b7SeY
6tL7o4DgXoMrs9oPrLu3oDD4RmEU/Jjh4u1jLFTFvrTC78iMc5nniwwMC0Fk6Rqlg952FOCOxpdc
gWjYpdnWtN7HrgXQJH+oL2YjhoJwoqrZMj639Acmzxg9VqV3GzxS9u0BE8spfKtGaIsj96awkXpp
h6YCvT1mBJmn2xBxU8mSIC9zv4kWKZAac0uf9BGpRhQqIvPZK0maLVd1GIkNPNGW4N0UZXUde23d
JeKP7+704nC+mAJs9AJfvMimXQEmaqmlVqWuKk1GC6F+hrvuw2QafVbmqllsBECvxdjidCurUSs3
JNF6FZdrROFr4QSTsf97jnZ/UkU0D1bxRYyONhnyl1PiYeH4AUkYFopmuOJyK+3z+RlN1O8FHoOV
aTYiKkaRd1YdaZgbf2bsH1f9UArOQmm1bEMVHuQj+KjBZsgZQ8WNYCh01P7YEMNgV4+yi63yKgP6
Q+yuK/U2avL2LLIzfmLOfSmFQtzVVb2yO+ayal9oxDVEUws2UcECZQyrXq73P69Lczrd9K4h5L9r
spvWRL1YTtmdN97P+VSb6PXwohlfSmXh2/F8RWcZOhUlKeLPmm0uF7lOHeRaSOtfqE7yRzaGF/L0
5vFHbVxTVSNZHQE2NhxQTEjt30eiIXsYS+uko2OZ7B331F+XdNeGmEBhmk1ZnSvkXqD/TituLgV1
A9Q5RFmSXf3E2Pci+09eW6IgYSJcYxou+CGKbitEYJF1T3IT0TFjIyJ/Vg485exrBzK2f4/xvOg/
fucLH9kvXayrtz5/0FNAINGlPLSOOd+smafrl/xergmSHqOA/n5Xmf/zT6oowc/AL69dKmL1anQn
rYIRtYzfMasD+8QerXPqNH0QiCsNUxkcZf2l4Bw8N8SwcnmTQHGUZ/7QIf/W5X6j7hy39ly+kfc0
ksCSVYTecZKaThH+J2mIewuVtoL3ovqh4zJHFl2jXD17sJwul2DHi0i9xEhrYHMvEa1JRARE9JHf
gQTfOEOBYjpcOp/HXt2aViFU7+8th3HJJ07QiFF3WkjI4UiVgFED52yTYhQ7RJwpD3C9eliP8eKY
CzDcX8G8JFblKpDi1Z96uuB2LcRidy4TIaeU9Rz996Qm9/Pi7B+TWDETmeSusn2UT29a73sPUY+K
DzP4rfSinsuxGkyxIJZSXMz7EyDnKVDwkEiu+g5JsQrQoMDdvpZB8dN6XyXELdn2s0OLabDRSQ+Q
L2HpAm4RrjoEyyFp2KMlnpEssPAqTgAcn40AaxwKn9/KNeNYL4qIvJY0O8eXeN4xIPZqg2atWa5z
lXwNDnegGxoIAc6D98SkaxZSF3cru72DF+ek/PCbWd+df+a2id48/IZG1+aiNO252Qb9j6EXDGmH
hc+gKTNqLxQ6iTqPJIHOo/cgQbaNuXMB4fMm10hOaOrXyCxn0uVQLki0JRz+AKb/+yBuE0TqhehQ
UIs14bxWi35oOIOxLofEVRX1K1F3fq5ODYPGYHWYRDQ+Jw+k3np7AaE+li+EtL9+Fo7Tydo5t5ep
z3j7OF9oJrWheZg+/SKGJtGt2yMLg07U5Ko565mjtL24K6r7muHQpcMjfojkQ4oqcSUIS+zicJCg
xxemTvbKhEoG4Nljqi8r5u3zsqmlhDzZe1W79TBp87DJybrrDcGh6ZGzc8iZKhAsfXOnIS4LjzuU
UmYmKCaFzFytX+tbDkhPXOXYxlvsXNC3R8hwf2qRMoxaZOnk+VIehTkoONl0b6AC0RN5bre1ucVn
Bk2aZXYyvAxE7lzW9BvlHXFDI1FIgaxFV0eGpYdv5spsxSCGKXJFHXVQ6BwqCgNamtOGhs+SN04h
P2vIT6CiriDI9TOVlhdVjj3YBuqcvqwOtTsP/WwaEV+RMC+e2VPxVHFbSluYm8FZWIpY+Rq78jMQ
lADmDOEdYjXEpwj33xYCus1SPty+AGPdBSU5mzLQ/7C1bgwERKouEQeYQgJUPrucGcjBaqI41lKv
NUoD98r5ZqTUk23K4QF2XQAwC1gltoiQ8fFP3MISmcldPxDCgxbSSlcPKszUPp/K3x+MOS4zn0gJ
1j87vB/0RcKLHHSnZ91TKle02OQJzSBYJ1QxIbBgSBRybS9WxfSi7MUr6Bw4+LgTP1QifVZzqDu6
HdZXfER6tlc6byfSsVCJwTrTpNR0TLpC/fxqS4HrPV+/GrgYjsW8yh6dO6ls61lOzptkfBEfgsqG
lYfCqxVZatfIzroZ872um07Qfou6cRo0/CL+NitW1+cWmFORi4M4lATVAuQLUNCpb8nyR67Eb9Ej
ThNoSWoMWWYXHAfqySvk5umJF9kIOj6Mi2WdH12EBBVEOmXgQcV/M/pz2alfi/sYQnqCGHU05yo3
6L2kEfzYN6L7D6YcBAw0y/X8p0s++DJoqDZYskE7ekGysoyKvJ8ENEOTqWnBN5Bn97+DGHQouD1F
YA8LuyD6iyhZdw1XHxS1IgMFASqJOL2SJO67rJ0kpm7KoKIhvd/FYo+kZwJ7VT1nJOxlzTfHobta
WNJcVFbqh7Kubds33gpSFqC+A2wbBr8p4wlmMm5rwdZ2eAH1n7jY6y2LstFrW1D8QomgxlRONO77
a7KObyGG8eZL/lg5YggA6WEFlaNEESvMU9RhpUpIVRRonTAqt4ocDW12CYTS0GugrhERUx84100w
B06yav3CZvko06kf6n32QV1Gcxr7MqSyLsIPB2d+RuXbAZ5Sl+c4NwG+PDSF/ILR5IA5wSWNidfO
gYbQnqGs3/CjK7j3Y8LHPzCq1tz2JnZlw/X+wsHzzjLMZGEw0LkD8vGwERrF6DxKulibkOuSdA6r
LM46Aj7IaF/jomh+yXG/gjTqritWmF+bxCi4ZOQEegZEuiNU5246UzW6AiEriklNUP+qwECyNIFR
V/YRgG1tyEdeVsDax6uNTqU1KUE5HvxixtstCGD2IuaSJThOh8Oek17TLD/sv2AMngT0wG47UWHT
BdDA2ZNIJoij8srCIVrmmQETjhwRl81ouo6rUsM+bHXPlz5pvY+4UDN9koRBL6iNmH6ymc4X5hCh
CHtg9cqa1iIA8xAo2yHy8k0OcVpT1hO6I4xOc1gNDlc6UGQazBDJ8lM/e4rGj3aELmsVHIsjm69A
Snn4XLuicEDFCbGILrLRjiMwnUq3k4+3fkxjdXD3mVXWhiiy7KT8J3y4EIsv6Coo//UAbR2KV9d6
gmd4QKc2E5Qapl7f/l6I6aUywbAPmVMdIunrfe8FFGkDceE4MXWj7EUtpDCZQQMgCv9dP6ifa/uT
uxQZDRgRFfmOg9K8e3CE+s2a5D66649QarRBHo34MJqHtGsBiV5u+NcDXLKuxN/ugqXZLvDyTWhU
UcKWeVONTwZdCvWpJmW/f/K42eo6O4Zh15uIrt+GTfME86ch2Zl/6SJZ3CMu81HMkQl4V0e1A16s
er4PsL99/Oag4xyfNX2NjdpJdCYt/wOkzcOs55D8zYLhVi4WUrBdPUWdQz3b55qxNeSIpePDgxo4
cHWDj0AUgNTnyfSm8zq1aBvGIR7uYs/lPgNBqcmNIEkWqP3Z2feTreFftp5hCyoz7vzAMheKZRUk
T9DM76+Gy+WD3TjXWVLxQ6Qxqx5lE44HnVxzyEv9gOFhsU/448MLp9Fx66qKnG6QEUdIP2kJsp9I
pytO9DpsX5L6VuZS3oiVx/4MDfRmV9vEbvnODmDrujiM9W5jOfMjHUkGRKhOEZAusp5wKIOlFrLW
Jv9FkCApR+Mgj8rGsSOOmd9QiuIMI+lrOpI70vwnU0Tzq/aSIzBdJTYS4xMyVNi8Hvz6/p3AVwK0
5ONmb2C0kvfZgNsqYH1oS05xgS/pFizBdcLp+c/WJsOYDVdRx813BNEWRWLc40VpS2ebsgsWYDXe
O4czXT3/qilVklatzc18VUCbTmRw8Hjk+P6gWEF2/RfmwOYdAkUCUKzYGe94RrE4G7TI2JNNMI01
nPvsY20uyxmAAsG0woQgBLjZvryTv+mjA4fDIdSJpFimNMpKmeXFhlmVU7EfPfBegUO7j/4PSmE5
dMEERXLV7Z2Z4c/vSW1d6qjUIkTsyBr3R8mNyXDvSTMXz02mCY4b6jrmnzxNW8r4zOhM7eLw+fLC
QttPubpc6Ix8omsIex5pSZCyr1ZnIkwA1M8/DbASB21RD+48bO8y7/LAO8stLyey/y5IgyhCP22L
Oi9V0E+e5oCau7ZnKPkHALlQTIm1pCSk4X49DXUN8UzrWBkw2/w+laHbZSQe6uebPVlmGRGxV0rC
+LSvn20CPmmiwae85cDqScebj2fXKCE5bMu8BJiRKxiilHqExQWdy6yYs4vKzUqKZMmylYtO614P
UDtC19W0erd2m/kgfq1V0vTakIVMx+bNWIzeYWGfjyGu8buSoZypnXzOPG4VX0a2XUfQyACzFqf8
DqYRqgZMUKhlyJ1CTpsN2SkEdiHg2VaOaQlzN8FoxMt2V77wI5G1KIG39hhPfkN2NHMRohjR34XW
n21HryS1sbDh+oeRdIc6BGNuxtHkBsTOSoFTZgs4hgOlMy3GziaK2eyiOJ73OOfquM+UKHKy5fwU
eo/1ibPUwwtMpNzX3q7SF1SZVzxrXG9XdF9EEO7XqwrQHZshaobAITmLR9B8tBE5J8nL4DRT3w/S
qkd7tBZrv9Hu9p/fcYi+Sb44trbcGwPGDpYWZwU/Rn4UTa2L1n8+jgfj27EsPBrzP4P1iUEgK27a
nh1QSsGvx7UvgrIs4+atnDEwMgf8Dx4w0GA2i/y3nnJ3wcUcbxJ+rOpFwvDaDRZGLPLrOwpuP28k
43E6J5QU3tDtnqxk2InrYmK4IWLWGtg5BC5wLac3BVnzo+PY80IHiqQuOcDl8hCx1xXo83p/ZqFv
+RngylyE5s8wgH5iKqxyRfv8loPV26Xg3K1IvbTBAobYiYzkHVqY+YFPshZVQYIXFp3wlKP9+bQD
DM07i+TqY0kfy0H/kwcrE0XgxbelowRRY1XOwW3pBZnnWxRtiZEpZ7Owi7NfWv88NCF9ZN5bsYay
aErpHmxN0hNIGhwS8tBS/rcFmynpp2nL6jy4fk8jWyXtMeGa6ZFmh0AMmGTPemk23gqhtg21ZgLJ
3v8LI4UlPdYEn2pw7Dvsfy1RU91Kh2/ykCRpmC5Mj9bPOEQOC9R7DQDwDrpidx6JkMNWdpJIxLMH
gxFshwonD+oBV+CkNRF+i4Qr2/mNnB2OqtrKBzyB5yU+oTt67bK3yr2OGff2eLQEc8CUEVrrHamA
djbfufWMB/FvftGds0SSEsnO/60BVGcYoD+bgj3JxoPIim7jl4Xp5TXBMOsOE6WzVxdbLRgY0sn0
dNW6sT4OYVD8FxaijgC/ACddT8Ll4RvKGk1GNY85Jk6I5iWQPdPFnsAM64gQNvb54Xz1oFCV86iL
t968lB1cD4jnkek83w7qWW0+d56Ul12/VrtHkIgEYqZKzDutQEfQ6/xwPAurjF5dgPPhdwPHR5w2
48bVwcGaJA1eEnFGajGLGyiTOw47sRFn5lKO2Qs0klaP5IRqJaHp8w7Mz0WzD816YhPDDS2UIdig
Bu82dXP4HtFyt6ZJDm9x+7TVuEct846k8W58hs7RmnInpjkJfL/YKA3wgO++6mDWZoCzfCm31z95
14yHxsbMPVPq5PMR0fJU4CEA1s8ZpxVSz49Bw1tmi+amjlz0Dw/k5bA/YMSS3Zg8BNLKutGf28do
Rr/KQKngLhkTMiCPY98TTfY9eIZjtTqvxlq+D8Q0CsWOxxALc3r/ZgjrnwjSsaASXs7kO5a2RzfY
62lE0QDcRkHp7zCNFz288GUMRfqVsBZNWw7WBG65pIfQDY17sQZ0lG9X64Vl27Ae5m/T8HSuwyUk
ny5vMfp9rcHp2DoFEY6RWgD4zJgv2QwgoWSL8uFO8ceX8sdQrWpsJwaEzm8eUBdubinoJZd00ug9
hRkmKhtwREnnvPnTUo2HFrcwCGKsbxKfjEpDjFsF+7Zb2TlYNHwmzVvnFIFbDttMOLqGVdFPRvZ3
M9fRxyRRDrN8Jg7m6TEZgdmBrII+WqXtkXjg98bqXJGGkJkEFYWPwv1NR+SiwkTcOu/Hq/H6+UQK
3lp7JbaldrvW3FntAH96eUEgdh06KsCpH8vWWlnw78CEL+OoRRWwlO3Z6sjknGChB3tDjCdxUPbQ
0AEXNtjdF2xMa7OhP5sc28mlXX6YTUNy0vGqnoUxmoiLRwsPELwnKIeuiXrjol8GCgPVXKgE49m4
fUFEEiFp3Wo2ivUVUM4BJCzsAQ1YzLZLOqjwRzeWXdPJPVzdIa3NHcIuBl3a9U7KiHQEc6Sbu/w8
4m0WjMRnV9OLtfS3p3PBHQwYiAetuS7p1NszE8wMZZd/mIErJvbm6bXBkq7M8BSDSppbIkpWaOHe
AbKpplbTMgUUccWjsFsLSFqtwxWarN2aCbrJ8RuiO2HwnDFSmdNmCr0b0/Fec9LkuOh9ex38uZ1e
joIb9qj54oL4rYnhXRm11c81i9LkLHARD42TnXIciXfhn76VM0gl107YJkSiN8400kyF/8VGD9D8
Bt90kk1t7X8kpixpnRl9Mdanhq6oYzZOmdVyvGCUXQChbNIZg+WhD3RF6KpikYfRw3TgRZxtEjCp
sUMPedJZgPTtRtwzaLupLxQjDfNtpHZHsbOCpUiCpzq0KFQQ0Kj50WNDLwz2Pkqgl9nO4Xu+C05I
iMy4JEyBa6mhi+CSVZBq6pF5F/Mm12xN10SG2AgS0G5o4kqw77NbPGqvAYIOTdmUSMi/RnrczqUN
Ccrz30G1eNOBtOypmWfx+TARK/yM6RViz/V+OAuJ5/p7snvMb2CLk2V6jNwgGMPKNsiiB2AX/xDW
0iak0K1u2llEXPMYgG/7XKurXkWNKDrGg52O/1poknlRcBMrFgLg/v6YTiL4cGX0A3sY5PXmQliU
XR+zibhLTlFb7j802MGDgHND0dn5xDF0unaJXd7bw+r//ADDpAQ/4pbrctr0VjsdAlMh9aRnOhvs
MEUsjO8luRVBhefTMQtt5IoG3mR2lVolBj+XuWekk1snF1rbq7Q3egFdisTDqE+nbYlxtkElh4i+
EYd/N5xfv4S4wKhOpg4wtk1liQkG3MuhcTdeRv7NgLzXyNvCdhJ+bV5nNz19050PGhbj2QjGKU1p
ltRnxW02r6dY0hZAogW4+Vh/b1ZXfggp2RMfqt6Pmepvh6NsckUL/YcoARM4goiuXECVy+NLCYxf
gDXBDvglUCXFquragaA8ROomJ1p/QbwtuqwVVULIu6nfjhDBC94gLF8YexYNL1C7RmtIGDDXQovt
t6XStvEtXBLR7KnaQrx3ekrvly7q1Ejhxq0/4pfirgpYPoInJmfhnmXAgYtEenjKl52fOCjnW8mq
ZNrB9I1GEJ35mIbGrU7iyVrTVBV6Og49zWCVx/7pO3X993Uflzp7ZioIfaOaebN8/QpWxCs37IH2
Z4RF
`pragma protect end_protected
