`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
hIjVpEJe2jjqMBgUMxmqpaKw3XH4eU9FbfhUes1IkupwSgb3AmIv3SHQS3PMorkY
FR1X7ZEJA5c4UWbrR8o7MYZDCi9l/rxUu2Jg5VO+gxOrUDiHbQJsrmRkT9vsLjCu
RB2F2axoirfTaNYUn4BqNzJX2YTgydA+dkj3zS0eeE0=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 4816), data_block
Eo5+aEmZAs9DvKI4cGWgOfJAVDp+4Ge8SYxg8OhYAagKJidZ+1rlGdzUgqlVktGB
gjupMqu8p+SPuWpsfsKR7EOsR3oPwNoZzHs/5G7mXHNwY0V6z35kDu55Y15zUche
802CVPxcuOXlu/ifczgbXbY18KYl11aQWRi8ndsddnFGIu7pmqw7Kx2+Hu0Civ7N
hzuW8GZzpCJcNW6ViR9tmHfvj/Txh9GReAiwabVB179XxzgDz5GJZVErGvBVvY+F
MmQVGe5w6RtQGOUH21bJ6e95vxWmj4/OtmHju5SeHHYhkVEC+jpI0fqi6IHR7PEz
LEEtygpBhYn2QijVW4nIOWz058gaIcNz9ODGahK2MzPFZiO+qrpSfLYzvfMgDm9m
80VJWXqTz4QpF0SRX1bPeznTsQEew9IsgXuojVbzHbHVBjNziGhGbDfl/jzRuDfq
dvDUJCZgIMjYYNMTC+ZoUgg7UwunA9ri80ixX8LW96oXmLjGxBXR98Jrt+opsQpW
r6tQV/Grtmg6AvC8lx7Z1yTT7AmyFtRxvkqkJ/YMAtevpDkJpjNIvVtAIGBaf6tk
7T3BSpCvIIjtrLFwT+6SHk9EibkSbaUy6ESJX0IUftvPh6JClRUBvTiKkvIB6zHo
x1ysSQ4akpq/2NFI5RG0ihsyNmfYqRfEoFyV0h5x3kYTDyaNOc6EgZmOANSyHNQp
q6qgDhbJJZfrOG9e5ly7ivUuxj1kivVlw6GP5E2Sf62rbrd5MargyjqBNi9P7ZL3
ksXIzkCInb9tWWkR6cYqD3HMnI8bg0G+ziv0qB3Aczox12l96/7d37RzRIkriR1u
erfRRg6gKgvmGoLbj7k+ZaFBGXpcltGtfQY6GlVCulomWPjxlJM62Hkd9XdACwT+
+UkkDInkZmzW8SkAA1WKJhZaRLpmVV81qnKVA9KQn2nbKQWAHqUu/JR50SGuePBe
fTIrw7OKI6rIR+I/B81TGU1sQI7DtSwh/skj4n44jiCuQweXyxZr1k/6wWyn7Q1N
kjelZqcVfTc3QoMyN3udYqj7+0yoj57YwLfJUNvJd4J/fGTsfSLfHrHxfOsz4EdD
69CgyDNEOZc4InU1OYSMUGNFVvnL27mdo/nTuCYeDaTnuhxcJc0gbQZkiUHsIECA
2bAVYUvQfr088rIzhJ7xkZAk4CmloJy61JFALOK5VnujsTlXPBLffF3G0hQV52z1
vVczOr6/3xCpIf88Sj3zMOMaV3BJDt+OuKe+/Fm6v14Fw9sNz+FRteJOItE7H97Y
gb0JvS47EJFGpN5JR+FHiY3Zg54SOyELcgoxwLysS2ajphPDRiS57IGt9DvRZdCx
myafrEY1kGY5tonEo8vzo+yjgyzNrUCvnMVjRGEfOPLAqaooVvtKHroe2jDYEJYL
VKoCvmHd1KbUg846E9xQXEboUnA0KjpwA6iJ1icwcB81LFvxDahmLbwFSfKgGlq9
jxhzh3bo9flJwKlEm5Kt0EKj4D4Pg/lbmTqxCC5U+apnqEz0L5bfdCbdpOCKLWeS
9vLKxuAFsdQikicBZ3Z3yR2CnyrqzneBHbo3hBg6Sd/oP4J6t1C/zgGsCnUi/qW8
duBfp4HynCM/f24OpB2KizNDzuV4b76WGe0Q/MDI0t/XiDK+kHH5rwEShbN3NPZM
cVHGKhJabRUgO52cjtyi/PnC17FLv96L5qz09+YuU07d4QeRVb+aQmzRgcds+SJF
25G/FFkJluLF+XgjXoyuSTeWBAfwtFTNPYGL/EQqmMDT0LZsl9+TS5zaJ/ZZKk9N
ZeAj0ghwIwbRk7kIlLDo/dXzxKY3gP6KLe3tRTg40rmxza/Qs5jVBVwnGnwKHgJZ
oMHtiwIVxmZ6p4kKvo47QNJVZM1VmfLsdE2j9b47ozITzB4d59AJev3LWeazVhJL
bLtfT+T3hU9E9YiNoIDGIRbmbvhhZDgLaHysi9z3ujezrn4NwKzuZbzji2LrCdot
/GzKkeiJQ/pmBUskrQJ0eAfHxP+usZ8DJQZW/T89UQIFtyDMcnAbHUmtc9UTCIUd
knZGacuFAWX7cDZ+WptpEOtrphtIUpigZr9EAGhXrhSlhaBkz3aMQVCGETIDBQ7V
OtJgZ7SCqc/NnJBYYbW7zb8DVYPz3noLaiIlH9o/Ps8sMZyQChE8Nk/YVnZ0eb91
iMQQ5OdKnXyii+u/hiOzGd7Wzb/zSIFYFfOBC8WHS/7yGJG3S5rt789ZnOcuLWWT
KaVK1kCh1KBMdPJcav1zanJ9eFCg3w5jf3UtkeO8ma/j9UJH4CrPW2wv9SX0fgFr
dxiGjhCTfYYgJU5Kk/Em2p/xJURBFyPf0LcReqGVBEEYtJlBKVYibo1Qdimrg7du
MX5yCB4BBMzq5k9Jpl3vJXRIERCyW9VCgA8KTsA19sqbJ1z+MC6kGyH+LnXvId6q
SIfdUTOe/HceCAe5BwifFmKgImWkQiG25sK/Y7SFPiJPk8Mq2esx7yN7idYWGUtv
3SeWpUigWpNgErWbAHOAQUXruj0V/Eh+zmTJdvzuPYa6rpXzSzu/ZXUrZe+WFx4Y
BRwsEqL9nfJCZDBYZgeEjCji0dWQpQbhsvvqc2OQfKuHju17SJj5sZT5t6fAD1au
ZnUh4mOUBnchrvN0x3nZ36/wYiIqbXNmOZZS9avOB4hGnvp0FQzPU1e1GrOWrJup
mvTZDHcS2Wbvvl7avwLMpIKX6hWodCSh2vYfEc5yzzZ37uzxMRESKS5oLoPnonkU
qRxOJ/icoObHxzikS6EiuK2OTIWqhs72lKMsuuCjPQwjK7k3MKXejynydOEGOJcW
wh2unms4ZHoyCSBecEtHAfPPulrlU/vBCFCsaeCtNPMXwdFWYKtkH8TVfCeN75Ja
qoa9wuf+wXFGXqhjzAah1Lj+Sm7VVeT7nOFzLtPi5GqHBNPciw44mWK8xXh810s4
HhlVlRspPjTyONV8MlOQv9WQir69b4GaAaWqXb2F9LyKLykayt4/wd3ZRmQdjUXa
1LWmn05rRX7qIBJw4zUkBaFdSqTuQKLLHcmI8HWBJMtZVFmFwLNwoM058F5vFHeL
GGR603MHD07aBsNEduVMRF3lfxNlGWHeeT8qxITs1DOtFqeviQaVN4lF7phOcPI5
ePJ7VcyP8IpzggDvHZqy/Q1O4hcVCz1Ca1u1uSWhlTM0MB7XeOD6YbsW7ZQYvL4H
Xkw7w3zeTrAjeuS3PX2ich00NKZjWyk7hOybUJopMXnBMYqQSheuKNnJrZERENTz
Vn1uxe/R6njDxErOlg3GLxi0r6o0Daa4ed8J5+P1Q/A73v4J8i86RD/fSoiaCp+l
V4P7RWwSZ4eZ0Vha9OxRlU4HOt3BGjhaIllgdpzTwFbZstFnsArAI0Gkk1OM2yln
C9VeQs/TVKkmWf7yCgvdxZnDRAZDm64tn7tkr9S6Vtodq5pPD1VqfGpgiQ3yo0Z6
r3c9yZ76Zr1f1NyeZfyQ1KwgpTYlfoFIzF0JOPDk38sVFROgHnhkzQQpFWOY3TZT
SaNfHGj3zsgfDeWggrJvtA+wjduJc4zy67ok5ItUS6P76ilyuOvun7qwGVnxWcM/
sJNYLeMdF4tPYkgsHC7IlAMaQGBLUw6S/bkdCpwdnTvh8jyXHeabO2OE0bok+SDO
9wiiEnIi5n/16Hq340pWOfkLqWWQldxcMTH+jFvmfB00/VU+El/mbdSkKaXrK6Kk
rN5JKdDM6U4HXE3i/lstU4L7wiDO0aqvJwLMTpCJVqBdRFO7ajf+WdtYI4cgdYYd
tAjgdFhmzcmt/D4FKR6DPCL9D+CPrLUNB7EDew0EqOsrARmlaQ5Cmy8sWwsI+Y4V
oIK5yX/OTGDbUa+eGDW4QNHR+bbp9ryhIta3UnbBDOCiEzLUmWuespmrPNznuDJo
bx4WlzxrmTANeGN9QVkyOv3t4/WL+B0DXw8oayfC3wbrrYhp7Ao2ySSXbbluaitz
m87S/bZEuooWphpMsEYi/PjWeUH7jBJU4ClCOemReqi2EeeqpenqgIoG58dDv7HO
udOuHksLiGsVfU25KZFmYwWaxPA+ooZDq6Qm31BwnaucKbHw1ZZISeA7So69NftE
pT8M8JGAvtxhF3zQ1fldhKS71uiG43OEKQK8WHYk3pZLpWrHCHPWN1XrycYQGlUs
sHphf71eSa8gqhnvJqc0xYqw60vz57TPXk7qaT+XHJIWnMgEOWadUvkmuISRN3Uc
EQnA61tw0U7RywwwB9H97Iw9COGQheJ20uTMkjNtp1lrCrOGlE5q+qb7OWPnS6QE
DDSAuZHR6owLyMIkm3TP+oS+CozNIT02nrd/un2zEqKfw7J9FusO3vtikpl8rtEu
0wn22/ZK/VSLyGvDKx2t6cGfl1WC3f30O0M1I9QejN3nd7w6Rspms/zUHa6vP9xs
xo+BMjdUMwk6cFERadwI4riIvOeXpAXVBCjuqgvqQJYG/qcNlbmKGQUFylQ/rtKk
UGeTpnwk/7v2jB32eloL4P/VxO/7bDmQ1MQCAxFZxh79gH61JhEtXXxL3nJRgU6W
zhdlLSaQ0UTnJwgp4GNti7RF0bBFFMbEXUG27AmckSqarjvW1v6qYWtOhdmf4lgE
DvdzyyUTNPPxoywecRQgZ366PWFbYQoPQchJqYYwQrzc5M8tUIkT2s1fCi8w92Jx
Gp6miF+f13F8Eqpm1p/YTDTWg8tT3ipk1gB6QS4aeBnHO5IT0jX/gqUzJOxQNVkN
F0wxUSMJLgkhDr0Yf8fTVFJ/YhasgSBHUKFRXfJq6LZOIW0Kuh/22lQP1B1ydgy/
8cpEnQKIQhTOAkBT9uGm9SRg//ck4Ro9KOa9ge55pzfMInlElGB3QPnxnks+dHy5
Pqn97EXWLI25k2nOphjg2eOwCM7h5cMQX2OpgEmvTw4j/LNTCmrdAa/0ioi29TRk
1WZdDZOGnjoAp7OlPkn8mBRYhIIRb9mcd5LcIFA7pha9JbaYIWlydmrUDL7ug8m0
uXp2RLIPIZ8+OPjNelKat92Bw8hcU7HUM5J3ZJiB5pwqAXWgZr+zaVmreCgP+FyC
sbcZLdqj9KXy53QBm1+T0INN1VKQ4hEPjJ/ba47yP5adyDrYHEiJlYDulAyNxfpz
AwZB2rYS2h1/otrbhCvGEJRSNHgEw2W+xmCWkhJEqbJ47bebcroYoD/xch9x8QCz
TjDzObQaLTZApt8Yp4I5jQes+59QOqa0R8RNq9f6hwltCy5RiNomaG5Ni68PUbAo
cPg8UjXrShzJUW59m4g1/4ONCoCULb/TyBpEEb1H+iWMs65XWsv0QRmV9HgprEyM
cNloX23eYO8LFgtTDjnRc9NwLTX8xgdQQeBqsj6ZKmuMDHxjSBROeEzI3nc1qOms
bvHZLimuvskii811aGvZXlOIL8G+3fe+QdvwTPLS/y9Iv8B0ExNVUv1AxvxiZRZU
T41iQ8G0qMxt9s8EiyMzm8GMFwaxuvvSOxeQEWo/oa+MxfcEW7nmEKeDsk/zmVuc
AySzFSaPiPfx6dD3MOM+g2Fa+3dvRB73K/mOqRamf3F1GPJnCUw582hYnJikBBAL
1DXi5ZR7mqzDAr9h2EgIYSAlnS/n8vflucc+9M5tUZPWrkADfV071OVI/e7sogx1
nB4+y6MmFt8NlYtkG4RYQFzK1Q0O0wXPnFy3ZNr70iUSLdGZ5+7iMoXPIwts30+I
1NL0TACHlb/oxLQx9/bqpCwjftq9OGs1pzhpYNOcEvZY69HtLvZOJSe2or9R6nA7
CH3CPa+9S2vJoEQD9vScENtl3y5vCxRinQORhefRVf4RuWhJGCENJLut14io0r5/
wmE/ayEgoTe1+zA2AxCjegNXwm0AmygoGMNzIV03zJCHtznjPQUB+1cQ3pRcgU9x
bZw8+enwqSh+3ZUifgoU03/VYByCP1pzLg6WUioyw6molKvddwgVfcJlZhBG5UXJ
JTucqGM3Le3JzzGi2Zc3LFiqxopecJ/VUQluGkF+6wNkUQwK8NIHw+EM+OUgsqcV
pY2XJro1K420jcU3lAH/nLmEho9j+lL8D1cnyYFi0purF5ovpLC0mTn6eI1/k4EH
UJoP64c0kJ3m3LsOLx7Zt2PpguhvOYvpc4amhL6LWSL9DsbJ89VwXAVK7EkjOVRq
FGxyzdmChxMyVa4nVCTQqhJ3ek1LpZ1WJ9ORYiy/wl6EeFbNjP3K1APJ17Ca6HXd
wndjUek+DwqCNWkECsohMKUbvFcG1yHtuJugnb7sjqx18GkX0W21K/2KGKB9qOsW
ur2wECY/I1bIUasDpQUyJwkivRbDhDdUOI+RQe/ep7gUD7VTeT32STGE+aYYEWMh
iSFrKLBNlF8CNixaCRSRO4EpCNU9rVzQe8uhIliN7rSWvvOVcJ++4tQwf5DrX7JE
/J7AuF/Yb79tIjwh4O0h2Q==
`pragma protect end_protected
