// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
b7s7HGUcmesAfnJ8Zh+jKv1boTYRhjStDmY/DkUF3XfIeMqWelJ7OdbAK9oZV9mf
fsL8vEEy7tPCIICEbYGH/Pnm38TQZbXRsPLnpKXXQNVBHr6lh+s4Z4184hBd33PA
w5cQBhDPfE4lZ/cYyoSZ+oktSzcyvmlUkixfzvCM3kg=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 5040 )
`pragma protect data_block
Z2XwDnMC61K59XLIfUWN8SG/c+vI37DLF1m3uaGsGE7X68wAwQMzOtZCPcbQmCfm
ZCkGc9yOioiueDDUSJQWKNljolKWJ9DfK4OWMLXvedADkcgFVVizBNj4JdyV4thx
fdMFV4pDga7apUOLvMVfJiffCF11xBlPwgjdK2Bwy5lB/w7e5hKBkiRKL8110Xq/
HwG/scAByXoTaqTOmn4sOzSKvXJL9vrpmeKtEWBQ5S6aoErRQaT+7Wyj3xDHfDHv
rhb82S17tpGdqWPlTCCXPpeU57J1Fj9Lqt4hOLPLXD8iIzpepDwc8wsfUu2ER8Ex
e5zpJTu3fJn/9JWVesHJfm1RbHOdgxuWCboh4fKHz78n9GWRghcWLWUz+mJmdDQh
+yNlZyNpBbBQ69Gp1F3pucN9ea4Al0ieJOaIe23lT4HkZIYIeTMkVxOf+BSGDLCY
9vs8VSBHYNTd9xlNJkj5sM2rcNp2pypHATB/d7F/SX4lrDphesPX0puFhP/hxcFB
uCw11d6viLXaC5vD0TPsjsFkJuoFv7pFWZMohFntYwA2qb75JFFPM+4E4IJbY4Nk
9SGVOHTOcHuwOxygVUIDZsbPriKkRAbUhXNqGy9I7HzsOzcnsNDqXssiWvhrJLZu
JWPRDfZjrCKj2EQ6onvMNwzkF6rodCdZ1QQLD4lyDF1Fz2fXdXe4FCyXglbqBcIN
jnC4viMDGufLihpYsiOiM5yUOYLUNRKskLudPLnY0eynVamXkKEBhvJkGYI5hrVj
s4Rdq4Z26R8ce2XH/xVefWTEDh0WjYc6cMZO6pMBdhKjFGZQUxqJUektvadp1kEX
bRTqFNAx2ceFNiT2eEICLTfHV76eQH2KsPVACQ7ogdIlcnt05rwRbf96lmQ7Rqiv
a/+sU1RwtqOA8feXh8RHPWeiV5YH1zdSY6hwWqKc2ua3dAojjjI+kRdhiVGAJflU
qebJRgrM8a953g3iK2ruCbxddhLLdGeVkc6xqmrLJiC0Iur1rwoF8KOaGbvGqKVi
kcH67ukUDOWHO0CnSFJ4FIm/eHSQW6twoNh4Qjp2JOBRKCjWFeo8uKtM09+0vyPz
IEBEmPLN72ZqvouH2kqIIr/rxLKjAsp/pCa9DgAgWdl9+4ob2vC9jKuYmtP7Fiye
6cwAKAKNwnD3uz3DUJUp0yrAbE8qyQH+v4++zLSE08YxFc/Z8NRM6lqFd/pCcqdV
0hBRkzU4g8QrQfeREtSU40WMA3CrWkdvXVZntxycZR3Txl8R+qPkiYcGHfijxyXH
YqVZWGvlKe5vQi3U0D7jQ1u+1rIaF+0TNGdZoo98uSP6YZVuzSn3Zp+5dhufGhES
mhhLxr3HQbuSPhEn13j56HphSQ8SdG/2qS7PGfFH3fUJ7GfviCbCmatUpF2vkw/k
fzFSABbd5E8pCPzZS8Nz25OLQ+dCi4Iy9VMrZT78O2wltfJRJDu4Af37EpsYOdZb
QBYTUk3cdsW9hYYTU2HtinvrFiUcEAFpkVJQj88kbEZod6I33NDbIhXYoN/mrbzj
DV1VLrQ9ogRQ6B3PRp0Ozlg7TUS0t/SJ4Wscg+jjyqTaBl64jPJUoUclFc8Jijfx
2WBbIcATi93srMB0fj4F24RaXHWu4VRS8l8KSgvNfkD3PTY31tGKnqHV3dyHHVtK
NUuPudRTGP6FMK1YcuOp1MqqkkSGbETMf7/7OCw2dcMMYLELXNg4DVxvouZBVAqK
FfSRahbTXnYG/aRykTR5NWrua4tKQ3e4i9W9Z5/uHL9ZHM3HtMPRB+RDuBmewQEq
wZqfIvCxkKNfG0blsTDhmgJyA7lmiL7eEQsKiwFGa7OBQQhiHFWUTEOU+rC0byXi
Og0eCyBYEy3Lp6a+MaRZ2QMeJyDcjDdahlPGEX9eRabhy1mQuYfSazzpoMpifrJH
puOlh6eXRHK2/01bJOFkmnDGx+SWICiGrmDHGViOD7cHvITpIxExfvsiWRgdN1lg
KAtkcuJOzXW43E1PP8vyC6X/fRN5xCkn9hBLbO4ib1riiXGGqYaEDTVzNAipZ+LC
iKMHIcSkU2BisXbZPGUBV9NWrzUdd3uPK65gq4Ws1gE6wEd/PqtUYIYrBFGMxx57
v+PpRr+iVKuWt75EkahP0gp891sTdME0Z18VN0EgFMQXmd/A50icuRmsYFWM4Jg3
0Kx5/FQNYpsnG+YfGnp57EUBtUfXz7d8VKPtu/ugzr7F8x8N+CV+vI/UWn5h00YF
aQSVoWHsVyYkH7Ux9Ts2HufIfMhi2yqzzMESN/c/Ee0wUvFlaIAABxGX7b84EsMy
RGsomVu6VfwH7tOz3Rw1elk4AjgU3pOHpCEur4nfeV5MMmSuhzpTH6P03MHovlo5
kQOo6uo5oUv7cs0ZzM/vRg/1ivzIvBdSW1YUgmVayJVOt1w+xlKbEMknls+wgPKp
jmYDdZbVFT0Qh1mjhV9/v9AZUh8OWh4J2omjF8qUcfCujrgdostDBYDKef4lGLIr
kTlnR0WuXa2ybSZldi8ETfTqnCKDBxHBarjPUVqNpHKiQ5iwNDAUtIo+5T49He0o
gkleMKdyLHyfDPL0mFREv49vU3XFCfA08/BrqjP3wcw4fwSl3B0o0cxwcgpIergC
5WyXfsKrvM9gmSKrTe87AmgfysgQqq9KgYf9ol3Ozp9Lt0lfiHagovit6K2MmiZp
8cIZ3oOAOGni+zOaOQ07SdMVfFpfI0tbl9q+KMKkdnLlQG8sNiXh4IJrdcNy23U4
mi3T0V4TwbMccr8p4bx58G8URrEEgmf530xxoDEFEPcwki+FrsFiuRmXCAK2TZ6M
fb0dT3OzcbzUuQhgB/WFWf4+LzmjLnz9J+dCie9n5d0T6X6Lsf/Z/p8jSh3H0X/v
UmgQgjoeBiaRn0RUd0LVxoNBPQE9RM3lmVLQZjZBgGIIsV4L4ei3923rdnToaymJ
B6ws9c/PlS0A+c74r60wlOldknoLccxI3WAZhLuu1TuQwjB8SL+lzaxLhQ+naCA+
DjZUCm0D7lqB7qK9OAT9l9v8vEZHxehB3/emcMckON4s6QAzFs25sy89QNHlSSMJ
AjmvOuIXfDKQG0ZRKBydQPehFaYrC1cNOSfWTw4kY2f302H94+qasR8sBPzf1efr
CiRxCqP5jJpdtwdmlFGePkyBQNck9mA3n1+JqgvQgIQ/QBR5Blm0h0i08v+Yp4Ht
N5RNOwQYtHnhLJqr4JxmKK4puZBNFFjQymyTYEoG2uqTieOxaVgHLo5S4MPJk0xS
KqZku0cIPwIIBfbSqYgfvCmwv/oYwygWnYT12KubCe+djrtb4xRmMJq0pwY0OXln
+f0G6gAAJ4kAlEAWyBpOIWC7gHdxPje4Q+70OXNVtSAhOBwKnX3ZljdonY53A1B8
nHKsA3FTzyBAh/SnUtFnicaBO6PCKfp1gE3fllBhexHuOfSv1bg3ukYh10OY68s5
xOMb2hqesWCJvLQSV8/dhqeu7RcUT74nK/kzkWLlK3S5eH4uQh3h5jbdKCIyxkJq
gwC+2mUhIJIEfTU28cMxIDHszGYp1ZttofVNyFncY+zIiypBiXURdRAeo6fuUyKq
JtnS1Z1/jgngOufRbn3O/6uCbsYyuKuFhzzNA0YYxaDIItDiZjGg/Dg7+Hx9/TjV
jn4ENabRc4eo0FzynIsN4dnsQIOB0M9dYVJlp8cIw0NmkTSUEtbHaOQVf3HiDSfz
1Cl3Ph04e1uprjVDV1ZX1MbR17X5xxm172VwQKndIBBI+lEOfGzFCKbzcwipuwVw
HxtC/AIo++k/ieZfkISWLU8MNKFw6i/qx32iaEH79nG81e+bP5ccN9uAj/JxbVsS
xOWfkegFMWB8KTPMPSBrRStvbGNdjENHck0OI0bIvK1RcI8YATo5xxPCOCOscg6S
3K+2jNSh9QSRRrFuXnkoUtEMUiFOj8QBHi+GBIxgdx2I9dzbgf18EAsuYH/rEQhD
oCb1a/co1GKgYIPPGcAImMx1WyOKun8MuPbNKMTDo97LinZa/xbBt6xJ5elMLH+0
ImUO0SUqWyKsWSqhWfd6TEM2I0aDVoLgFUYOPDTAvkXyh9dR5W4atM/piijBmA+m
ZQLgUQ+BQN5t56uFvKe2HUCxmxHFnq3MYsRWdLYAeeRPkBaAk+VfU9o64jk1Cffd
Cd3kG4ZvC90wBpFjkjwpP+G+WYD1Ow0uot3MnF4uuAth1Sk3YyfeyoykQCYe2aOV
RY+rrkGypvDXlLt8KgDV6/rLD0UWpvi9WScM29KqPfw4DWtgOU3jYDQWcg18/F7f
IdGxV0OXG+zIjoG+WnjWav+bv1GXmeaHu2pTvyQvvrwsnV8cxI8CKUU76qwAdkWR
msIdrqbsq9Ldhv+tjx2V1RHug07GMf7BIs6D2xLFF5sxdaNnsELUE3YCjthwhyHw
nZM2CMvm2BmKbYkm4DrqU5zNnLiTNYtzyXEqO5YLcm4Kt7YeYtY7hsSa+qNdCnpZ
OhjI7pfhLaoMDNfCdlrizn6wDJLifjsR+O7J5bhHWtCyBmugvpTUXNuCqkhHA/02
T9s33D2FtHLC/foyXJo5Xhcq0XWxrJGG7YE+2OLtHP/XPlvFoSLs96JkctPpvdg2
UojjS2qdtIfWD7/8Fnh/h4SSD69my3tKV7g7pzKZ/dsk21ArVLlnufHrlbkin4VI
GPzEw0hJOm3w+71N3b/b3OGzRGOtBtpJPTGb8F7p+57yF68eqzzMI4RLY/LGudar
pthV+zg2hIfdmr8Ai27i2y24kF7bH/lgyjelTLnFMIjdKHCwm6HHuNqpeJGwp8+U
gcFPsQvfOEA3BFggtuUSIT0k9vMowEKaelq32v/ZQBmNpR9dcv6LQWrfUX21rjWb
/iHHfOiHUQzCELpF2jjCukpUFpGS1ngJcgtdgeLIvXzFOUmQQtZH3F58HzWTDs0C
KO1r4nrNyjsQ1knJR7Q8uLzwUFf56cz9FPwf1Dmg1ZYjKyqa9vzKGBqe1/j9YzJr
JtPFJOqjhXHhvdYKoH1PF4T+dSZE0+ZhEx6PSHXjXALbu4+i+38GHGth/t9+MbB8
7UJYcIQRqC77orULKl6iJpxNc5+psYQ54CwUNFfOg3Kpn1kZrwJEHFqBS9NrsOzZ
8ytIlLWOoeQoVK+3Ivyr0ruYhTnhQAsqB94XT7Jrr6ZlT3G7F3t3MwFYCXXjvF+i
Zsf+W9ZBTJxda6CDvNTi19Kv8Ai5tu/jITMok1P1v7O042LfBXPqbDGBLDP27ENQ
BVttRadJghZaKPFPDqbxGSmwoNLeqZf06Ke8d3go+vMnsbGcUSKu8W2MAHReKAjt
y0jjIg4wx7eS/RIjgn5/VxsRMtbUM0Ak3LnD29Tn+OsZxhwIAl/ngIz0pFz5Ir6a
1wD12Laau8Q7d0cBqt85l3/2//HPUxuo0+AyFDSowv5FxPhBs8oy3qDuGZ3RUaQF
piUlgUwoX4DXk2vemyPz9RyR0LNLy2cVrOEaR6kTNJCHChLPEefW5KafdIifGyJ0
PDdGGpJ/zwo7/2js2iSbxT2NBTF+fOEOWuk0FOwWhIBx2yTA9vhO1vcA04Jjjl6W
x5z5iTOORtKIjTw5r8PpfPSarTnztyUgHso0pKUxHzpMuidKcLSVySdGgOEzDqt5
t5v+EEeDycCiMRKnq7IX1PNZoDADEDJGWe180aNo7xM3xQ0DxsEzWPXYj8bqpzSe
GRcD3D+cowC52Tvz6VfeutReR3hlnje92VNsLF2UEdBwfM4Lciu4q/MW9nNqUMgB
GvtGEfKEWZfq+AFVAfjJCKDxZ9+2cJm9eCU+YCJrTvM9s0vUt+DnvDFAz6p4aipv
up+Pd5AWZ9P8/yWrJDMeJgoQxx0OvAeue0RIwas9FPjUi0emUWnt0/HMzp7wvp8b
uZJyytyFgu+FcN2WRO+U3NrIYSi+3vOFeplY8OF8G/ZdhVL8E2TN9382fxnR6f5f
Q0w9dh7zMdfbl2aV9GcLdUWTWIa2fVf/xIG26BzBU57oAcrilhXvbRcNEDmylN7A
k3jxXFd4/8nXiCaxoo7Ym9dNFbRISpFjOIexaI5oBELNa1sEyoi7kjThob8Dgpkr
/GePaL6INkLCxUhyhm7LF3EimnFBzrSp+TpEfEnHUtBWE1zEpw9aP1xBwM8oYT/1
PGKjfUpUxdSkk1OgASwD4+xGmhZHoks8yl14ErbYFailHlwC49uuJlbGoV2QoLS6
B/vTBL9SmazMKcFv3Nx4XWLFP4JA7mgt4H2mVFzmNunDM/ohyX+0/YMZjUBNOPk/
c77wyU6fj8cw5paOY0pzqwKJPxwfWw4Tq3fYVZiXui9QyssT7P0p7mjWA/t2gFyc
5PeCL/Ecnny4zM5lWuu7XRS4dAhrmQCc1KYHHE3swjO1W2Zuks19U3SRRQcAKkHb
GqT1MvsNiURy75tNdJ6D1fGQ97k86Sf2TryYBads3SlhbOnm6Gai9kobtanOnkIH
sye6q1ymG3w/EXsCHCwZhUGF6o0CgLZ4slyvaq98qASrGvYlX8nZg+cAd3BukLxL
Fn6WRwV+P76ee6M7aTaCB3efaaBV0aeSHYf+idGP72h84myzoK5YoUJTEe1WNWrk
qujdvTakU43Z5I64RN67pcL/eLmoTFnVzZM8+yb3cNVBF7b4k0CkEdRcdoPuGvfu
97puEx8rKvKoCSXSwlPwL4vLs7U9KfaATSR0nB85C2FhugKOLHC6wesuoy2YAuAv

`pragma protect end_protected
