// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
cMhuIiuGjdBg9fiT0jgnT67Ec/8HSCuLNc4Cj+fwLVNSZoa/7NG8Swr+LXiH1ei1kKf69VMVIiDP
WRSfb14eycDitXmLxLy9Y7RxwMYVHlk23IYjPkF1EVz2dWEiyGSr4ssR/O1ppI1gCh2yF9i2BXOm
YtrDPevDmZbaj7wU3EOt0BRV6Y2pKjwbmAtoG4aFbZn/D/DljTybc1oThC0z+iJ9l490MIFzCsA7
4PxnJEXa91DoTjdBNNQFTfFKzzC0NTU1Vn9BCUZ+xwHs92aE4wdX1tO0WO+7h9iKnlbEZ28zMGIp
mtDZ0SawQFXqq0NdWl4GxmiS6YTJ/khZN+dzwQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 8496)
REMvS7A5gf3KEobB7e7RXDb5TBcNY2YkUhO2IIvtjBAsEb2PFydYOXKtOLJC0ZwiMOd0+5kJi9HS
KJ4SK6dQnx+bfdqcx895obkK6GdfhY8Mz7ksrewJq4U3dSBooeC6DHosZpjVkjLRriMGCycs5qjp
T3f1XTNuemgbsSQHGTLZeREpAa/bPxqYFJ4gz+4sv0RpVnHLupJa0V/nRD8UR7WUes/hKHXIdOZh
3MnDXihhFP/w6hC+qH26Gd5UnHODMj3Z+EaibMhBEsVIyBvpN11IFhyPeaVGInMyM1ZjJUoY+ZvS
6X/ldotE/JlRZCwBhlw3xRD6Sb273vio93CY+IOWkdvCf2UnUn7kqMyAg7mAq4xmjn3x0mwBNhoy
FZ4BlY8DIpOzn1ReMtVt939P8XPxr+F+rRmyi0SSq7kA9GmApu5YIjmUEiiqu3EDwMr/yNR1olDl
/EFBYUqgiX+LVvyrobhqf1BwBfNOhtZmwIWpEuzTuSSUi26frloXA10INMzAiTlyhuYLTXRCsvdp
Pi7mAU0QBMrG9D/J+8rBZtwLB87z31ImDfYl6emH7thoBGbYptFVp+wsI/ktkgwOeeQ4Z3/iKfMH
DmDWx7aPLX+IVqfhElfsozdwhrbpIP/fZJy6Nl46ZbjDyAKlSEELfX+F8FhoiiKPhrI5MkuijSJj
sPXsCswz62ZACvnluxe63+/5K9NCE9HvBb/9xEot+hkerXOUzxBFI30/Lc2TI5u8EbAVLevXH7qc
mpBA+pu182lrj9M5xMnGZHQ33dCkJ88EzTdM1xXomUrTF2uwQmMoW+4bDgDzyU5797uNgRyYGT6z
qSaXYugqQrmssEfaWFuUo8gdsHbQUfo0kEZHW6wtve4XTNZr+0AVRz+Hw8EjvucBnEUZoT8FDsI6
gvRVLnjIBqg7yBTR0pqEv+pO2S6miDjNH+u6psIcmsEJqY5+6oa/HdpelrCtbM2sx/umQUciZ8L3
F1EdF23CVedLd8mZ+Opto6vATM7sHmwR472z3rXtdBFcE1SpRmayAAj8uoLRqftwAW2Kz9s03bn2
B27/2nyuaER2fjmKZfHnlhLEVWe1gq3t2OSBxo2KtIcgJ9tFBTICALnb5/R+vYXoDuI4DXEBADc3
DqD85/ML54a/mbQfFcHEOolIW4744RNO5q0S/b+wtl1MLurDLrAdZbtRzw4zq2zziiN0H2bUy0Fx
0Q3vCdOrkNqaMaZMooOFF7LIp9vf28YkYFWAOYEXTBnAXjpldx+ND2scahLpXcpgU1v+XTuJa0if
vT+bYiw+g7Wun+93EPKJups+1MVFEoSTfKjLSk0seuxBajawB5wIrToC6oxEoCX5WRtihWhBJB1U
+YSNsAp4d00WDfxM1DZNq0SqbcBCndxBva2qP4sdvdlPKxiZTlt/Cy2wzOcVFDSnx9oEOjulJtXA
l/r/+nR2PePJKvFWQe0MgfBdyHtsb8AzwMJcf3YCc2EP0brYLYr121ZIq32XiAgsEdcftlqPf1El
MJaFMjwOz4JH3fz3O7PGOEzqkLK/fgoEG8PmtzeF/dlGSPvqtNIkNIra86kYuKnEWQpNXLGpF6XV
qv3pYTzpXCbcMDLwvhAeO7vZK5hQZ6aqK1eyvHb9L91Zi2tIulGhqK6FmEpdJkJYprsPTzHaurxU
zeO23opievJzwbhMsQopELF4OXPTjzDqcmyVewsaIeH7cDuW4f+b9/xMV/W+XF0LG1vO1VkPK9gK
O0hJXOkpvsJ84HAKtNU9AhTJr/ks/PzlglKYZTbcpr7ILexCQbftXTvQiR6z5elWy3z6BfaH2/NZ
/qe7WNX9Ggw6r4PF5LWYyvtAq1CZP5HPDAiRPw+VoW5ERDz/+iDEHpf+Joq3RqRVfZnrGSzRFn9o
K6H/laC5nydSmhENojhcbJ0A7X8m3f+VTRcS1COHCECq6gK1gejjkZ3yhzS5sKTh2+DFkmXhFEoL
KWXcQriBBvM/O6xWrGVq3Dq3CbnSUdlZnxcgGxNGCYZny+OBudz6FXNKmLo52o64vWc6GUI8+bFc
cRlqjRmotCNAk1QxvMmaBcSJGPKiNE+mkDKGS6mAs1I5xrzoQjt/AB08mcL639WuCtdlPUqFXmEh
YAX8EHe0yEFTiFfC08gonEymwCQPdDICf6UxznNnZdFJOveOEalwArRtrE4ia3B/G8GdU0WRWvLG
1ju/xetuuSSbOCSbo2YxqSga7qqGnYKqhkxdfbtDDOuHtiNer5RnaFX8gbcZOWURqy5/mU9aIN8F
3zPARYEzZr3uHJTe0J9azxYwDfa4TVix3sko+JiwfyhmlPMzT/v1FaaWmpo5Fw0B0Q0PA5TKkpxt
bChHjzMB4U651vk1zxA5+Nc9JaGrFsdXuXcE9VJr9PaN0lU+1Odt351WLIyZyliMZ+EOBkVhdvu3
ZmNw7NAyyRdL0OICSzsGnfkN6lF7wwNZZAaWN4S7A26w5QI143xXAD1WJgq6aZoiHzum/A8dA6o6
rR9si8hDUn4ff5Fb/YWSnJLdTyehEgqsxRVjvsScDKymNMA8WrYmX518+TwjE2S0WaMu5dVld5xz
ZEbJDVlGYlgk9vxKvKywNAClmTFZLHN1t6UtjQQvswWxDfTIC2HFc2+bbDTnXYUvt/oXSAsV/J4d
AZRBI2BsZB220tCqi+JPFe7V/lELyE3/XpvEIoT5Qo2QYPXpGteeNdXfkrlTmauH+Rabzl19lltd
g+as4iL7ae6AP6zP3ps5Kdr7pCpLoN04fMpVBgW5+ZrLHj3lWAPbVW+gwePtyTeVByHs0QdoSN/l
WFStL9sH929wz88RRDVZObSrTQg28CHJIcvK6hD/lxdDP16WjghdlfX2TkVUfNo6W6m9WyqnVwxY
MbYzEXU8l5dc0vNIhFW/c3IkwS0DfzawSSFO3aiAH4YPkuD/ZQmvEvzV8HMtlesPK4VKc+6Yg/D0
0UBNH9uwLVtymmBbXdU6XBu7VXE2aZ7w2Ws3wypUgyZvwa8f5JKkQxeGdtb2/fP8/H5Jichi5kbC
CKGJeq/n2vUhASjp3nDKHYt4jozTwcvv6RbUnFAc1E24cf6upFcXeyA5jPXssBSkrCq6uWzqp+W8
CgIPYo4BxzEP7a1HW3i0sG+IU4QQeXclUcCwD74cfVU3VFmY4sHUPlI8kwRD7shUKhqz0Ohazvm1
hLbJwDki2HBepuxKOFGRltFnBmXtm9qX0+Sfn/mq9eGz0HyG/0gbu8vCvvfHJHw4ZzRFK/IQXcfZ
qr7/T2WpPvkP667v2V9xv0bIVUyHv9+CKzb2AdCuppDP7Ufncd4HUHwLNPRe8P8CgNuZ/PhZO9cR
VOYoDdi5hzny5KMfN7/PfJMTBolyszHIYcEVAj2UIY4Sf/Tj9fQFyiyhcAW1S2hIcqiWwc7QaCOf
+DRICEieI3Z0F3fest1xEIChCaTRTpamOJq5z1MsPN3UJuNMzq/E+lOL1AH/+N7+kaOijWLp38el
tsDYverrOxsBuFWwmMbEU8JrduVOkrLa4ou84Fonerhe6OFfGa5k9jzuWE7ArtBYWKe+tBhdKuDo
GIBAyZybFcd7KmFeafw9+LyqZbXYgnucfD4sj+v/BAz0YMux/8/hMXbTrkIKNcBLbOCWafisu0jz
1dTZU1gBb0Xn8l8qDTpuF5nfGYm5vzEHx0qotXa65U/s300+mWek3SCGe4ioBIvqUqiZjW8SU/NU
GvPT0C5vokeFM0AQTg4ebz+vs897Rua11ptVXGGgQg4uyDwa7NyuXSWoafoT23aiE450djejAwuc
NLY+Nq9+G7yTGckYLdXtR+DfJ5ew8ievgHN2F/dvHz5Lm2l6HwnHb1ieYe97JDAB4024RDi5Deyc
iQ/Kd9ZSkAK7hN9FanTrT9MkGY1pHyxrH8+hCvLG/7W7pgVu88Wjq2z7YHIsmYZf1KNcN13B7mv7
MYOOR6hFFA7NOskH7UZXQjaru3YJsB3+2LhselVDKtrWCSyrc6I7Yp7f23MbmUqY97di+ttfG92q
Z4pKA/WyFxatcGfv42ExhvB9YIgDxTWdlK/PUjS+mYae7CGTHlQnlu7j6xxq9Ttvs3Gn8dpzeE7H
TxZy3OC2VjhTNXAi6y3KZ54YQsoeoILcPrDGcDuy/adHapff82TMGH+OXdZmIS2pF2lpY2Ivo8RG
lIrNpfDIPXz0oBrWWGUB6NMCY1L7qrgWZCZxNTAth1oX7+2eol4hjvifAbIOyP2twr/jI68vmVrM
oLi06QjDl6S6Dyxq06s2zA9z69Lo3QCz+JEPmmnCR907LpVDqiI88NNxISCpPfYBxOKq/nrPjBHJ
jOGCTuoeNQCI9Ow7zBImkgdIHSd2LWtN+DKZ6c2CFY7EcH90lj8VWAohMPShvr6dKyMLVfTWxRn6
w5drWjmvgfB2HXSTciFgaqrvpM8IW56DlsqFt7IGwLxQ/oHNQLpvmPrNfAyXmvR6l7Cjat+R2v/J
VRooJFKoi9PUmR0rYnQ9i8LHNI0vXjTGqcvPeWuFdSwQvZDSHm0eqn3gySxlLGJolQ2/LUwyIySE
0g2cnYdN2JpijarjtFRBCN+zMu/7taMtA9On+3mXSJODPU2J7vB8bJBLXPRDUvlXZzxpQJdqSKm0
K8RhNIxZKpkncYjp747W6mYsISgbLgoayifAWU9YHAESidrasq8Qlr+s5QtJFpiLF5KSKz/ZFLKC
lopUYHkRFrCMAquSXPXgbf+6dxlvq4xDjvkTo6njWM4jJlCE8rZ/QWM4SwL5QEtiatZOPAefum1d
Df1Ez3K2PYX6/camoq6zuKMvQBskYvFhnGCz35x7GtTsllH6UCo/wGEdngr151AFOhP5761ZzqL5
Xz7Srdd3RknxVgzkyleA6FcZGgeOiedXfVMSAx0zE4GrCEjMmejPSZ9OJPCa+vabLPzamtXR/lSd
b4mDD+iHL7I5ZtUU8tpKtT+Ne2FlxKw0ijl0mDKbpaVc1TSDLoNytBt2Xvshh/zEmaYT+EkN9ZwJ
Zq7M70m/alt++yTrFwSedg6J0U2FvKo4cP9RJDScnQPwMCQviPiegEnmdvh6tfXGhHS3cg/HfXd1
SyZ3ZD50kgtTdwrFCHZe2bdfzQ818wzYg+gfF54a5TPYoQvkriEsi4yt04IJvnLTZ8WTUktKplAq
aKJ6tXb/jktV7Rbmim2SAOPjotXDO7WRNn4nNGMhaLXdv0OUiiONQhHN089+gt7LYz0CI4Yt6cCn
VtIWtQ5eUVAH/3VNgPcmOavuJvBxKeANQor8wEcsH2uHLdYVlG6AzqU+G0Po5mKS9tCKF4d0fQlM
onHrndPpmGeVeodbT6f8AC2b7BrcOX7FxGIBnLhiGuBpFVu/ojcqgSgYP6BlAdgrHoq+jTveEZmh
E0VjEzBRl+VUb1+cW4D5KFV4Sod61LAZpd3oSuWq7JwdaBDLamnVQTy4T52paIkufYpWBaVLX+dH
Ee8EHxzJxNraB0NmZVUtKQ7t7TgtsygjqLxHbRtcAKv6UgOvFt6q6fLM82w3tkD1Mx0IkiHVn57O
XNgJK+pSYVMDbq9nd5FxxXPZsfY+/S52l7OC67adjuMF94OBD+0drUm/2bDdlImATrvItsuV/Ill
rVIKFQHMOgJf1UbuqLww/QI/RejEtqmi3tp744aE1ifnlsf5Rn5+SUNaZDeaEgiRsE6ErNR3jvep
RQDhacWcAMRlUtaZhts58FE1LKuvz4ydbV4ETQgxcGRvIShiA1pRcFJiFCEO5CG12Y1D4lKnxo+8
QEMjTSJmyBsDw22MzmBdHAd1wROnEgWggDLTC5IWhOj87xMe21mExNN1AEwUNYRYf5A6ePVlhg19
+MAF6kl9iMu4w3CKzSO5Ir2cB+EgBsdjgPn0+nhWlP6w6/tHAWrMcsNRZiEPtEcRrA1CYRPdayHR
8zQs/jFycUoMaMM1a0ZQO1UFh/wBww3joOwMRhO0CrwytyHhFQu6eettIYav9Lr/ONhR6Z0ah+jy
FhiyOBe4f5L0ZUmueK9S6ooUpBXjDZi1D8Az22SW/Dir5Y5AnqjeSwdtQt2nnfeP/9FbK4HxzEZn
Dzh/NBRrgeWwXZE/ALAnYgcrCMcrM7N9DUjHJXiVRVTKk5H6AeIgGnzed/7t6nw1MRBcmR6qJ7G+
DvmSz1/ZAJ8Lo3NeYQlVOtd2l0Kh03ct8Q+nVLHRllpZsO78OxCxA7Lk/9jk8/V+p2MAkaJsC1uv
o+RHz8uRneyASpMKG9CkcCrN5vheauPxzA3k7m2rAEToXtOv1gNJXS5l1Myg/DF61imJV2x8fF+D
pplWYqHbBxCcs7YXVmymgCRZdYdg84P3Ip0CKUDAY5c0xd21SfRNRGQxAa6TdeVtRpFlwkHeh8/L
M/hc7u9cSvGnXAoLs4fEYY9IIWpFCgeF+rBMjwVNSKIHW29mtzaMp9Iswf35zplZwTSpJnjFPG9+
EthRcFt66j5QBGCcb4crJQYZzxLwx4liqLvFVvyB7RHKJcwEO1msXVJHZy8HXd0hQUZEw5r/AMhb
uL4/s6EDV8N5AZRXIauFUTlLQy2EMx/5e0BqlmzbNw+zXgoVQd7pSZVitK/hXFmJ8OjXlTDUvEOM
6AceuNtlM6coJBURabrCbHjSF8ClI7WiTlI/BjsdpImCs/8CprzkADtPkhlzSTUZWDg+eqbh5jzg
ggrNrd6lbGxlLGBZrVDZGkbTWKhjTrM8RD/EvjEqXVhbaq2jjbuu97sHpXGuAy20t0uBmEhvsrUr
NUlC26+HzfWREX8cOMmc+V2CzMcRiLsShFPHHqoF9XuNesDH4V5FJshfXEup0eMk4Bch/lGAr0dr
a2Al+LlZ4VEQoeFLcqH5A4Z+DdaMjh381LERcCogCe574N87ibQcLpeZN7WbpF4AlqrtjbZxOX2/
Vp/sCx/8IfFQ7yz/uY9EP1G7ZFcfGOTpfsbzIJ9F2QM41iUuBN68u3Hrb3GhvvXAoaIodffc87W4
HOHi1Us6GyUAPG+fX8g59Lck/GJYt4Z/a3JF6F1bdTUOUS3t2OdD6laVJQl1Bd0YLd++Pi23t6qW
vQeXcm9kUsS7M7AskMWSeKJ/FXtqTpEjgAGGYL+CM2MOE7NYaESIigZQa/lt/Zg7qERoaq/ZTW08
lT86q3JIuK+DL+/fAnuHXu4VbWoLrd0GL2RPgGxF6IrPBwrLhx4aCwoXq9yNYNfNh/JjRm3rTuSu
GqhelRWjRTDPSuEDv91NuWZkTbAvAfY2L5F0rtxpheU44aUJo8lRhFqoi7BaFoGbF4x5hF7q7meP
BQr7YcT77ObaXp1NK8HrK2JK/cFpB7MOPCJJIJ7FGSkgo/45ZR/j7Na6CJMXkvhKJG3nXR9j4YlM
/P9ueC93K5joInhmdPXjL+IAR2nGu7nbdup6ub8fw1OzFwsP19Fkk9mBx6DcEHQI3kzNSNB0u3dH
lFru3GmWXbZY5zLOiBDYNYQT0ZOvbcaD7Xo8XuJaQSmXqQ27vwYJEZ+8z8sIeoZ3kEWnV1qi8/Mp
DlB+thacrhVFd4SZ34a5PxQohz/JKh5YzhSl14yLorQIe4zYabOGVpkdoShnr+AUa7joAEAslCXA
jfo45oHQ/H0Y/W1awQxj5j9rfjL2vtph/REpkJGyZ/i+vtZmziM/+u9QsmblZuwfeZB8K+DV2Bjm
SR5jtdMg5Ac0/XG1MHLwMMNPNJZNm5Lf4CXoib2vMnvJHippCI70DEM6Pa4jnJy5o6otrG7B5D7f
VV9BW5sVADGm8N/nb7O2Lugjpd0XhDqZI48o8nls0TdUvuI+H19NAA2fgUxE7fBPtoIzNIrqw2my
/K6QWZpR38i9kfaye1i8E0p/Lzk/zyGNmjpr2dYR2KwMRG+SqOebDQylA2gBXd6AqKaxPITerBOE
w2fkHksG2CeBT7+Ho++cDMwcxAGBnfKymbfG3iwz0dfZ/d6YyYJ4nBGmPbHcllqZsMYcV/x5TR/n
tIkOxT0LjTxEprC/hCzhiknvqY0EpwIULdsDLjNaGC8ovN/MNzeQ6KqM1jo7jFwdqQaga3YUYi86
jynOoUtN5OW0zfVVoKb8hXsQiAPd/28OE4vi+NbO06K36DT50m8sRip30Cu1UwewJCkxg1dxMFiF
oDcE1MrQ1cWSN60Jo9TzyfJBfP2ljNFajnjL7mpb8Q/Wel0ZgI9AdxZcF85H5eEmul0APGdht2F6
dBEcF1l4X3byg62y8KyvYYWFi/E1zYhJ9vBUMABFtio+I8Fzy6b/xAh7kYrrV12OZkXDIH1/ELQC
muQkgr3ydkm5NujZ6770I6yYAdY5mYQLae0K7XI1R5+6G2VF+c6xPkEL9k8pRgKUGJJ/ydP2ZQ+V
vqBTRaQGFjMOrr0YQH/eQL3vxnN4eqtMRUl1cWbs2dqJnZWzcVWAUfe1jzNR9NwEfOw3zkCxHNnJ
h3FulpMnFxajGiMri3gkcGxkJPqqWX2Bc8rUnyo01uOaajx8fcBKawjZBO+hBEQY49JLWUkdpnD6
QCViYfzZj4L++s8+0Lys5zcLCPMhmwX17ZcLbe9Zv4LCu2KRpc/iE+MTVl9nWCSpWRtZoogrmEWu
3FFOozZYA43VkMnwK1NMg4q/0XTpoSRfrU5NfcnuML81jc+ewHpCLeRWdYYVHwaIetGGUC2YVRxJ
/AO+MI6GkF314ivG1XnTXUFY6cL/ca8TvBZSWmrWqCzeJGttn2+7F2ZLrctaSe9MYH5kzznJLe4x
kSASZcVUl6atOLSmcLcr+ZXuQ29ooVIgMJIL8hfVVyfplLWbbT5PCPTPI+ani7UhTIWo7wcOfuP3
yR0BkykQ5h4k2owOIRN756F+0RzRcS2OZh5376lJhuZCo0FDpGAHY7SA80WSruDZpkQqBQtkciuK
5jGpRRchOwKZxrkfOVMkp6Xz6GGYOB9OoKuQuiHNmdyaZMYDVMhLLdLRsZrD0+AbGmlI7S9SD0sJ
mWKJgo65nh8oRacxQGFJpivIOW6t5FtPbXiABYGtFVx1WUjpgz8cg4x+Tp0OCAY/clGfRob0Voi3
YltP4l8ye61X3hviJ9BHe8bOAwvhQXSu/bSqzHvhQj0ZLFvnRpTGs4q++Qx+gCSSLhVXaYScZLEd
y3GMAufpkKCNPj0W1YXYPUwcPW+exkpZHShcRSpbTSXlaCDIUDHQiZ1Mr5Lon0GPDkTGpS+NdntC
ZBLa/DHU/cDCpsAjPQ6zHlU/7+F6ykd41MVufsEXGhlTtQAANF9vT2btQjz0yi4Ecbj4+mBI/5ML
K7rLq7aPqVqrHq+YMTBFWxAjr+v/1kkcg8xNUbZPXOS2izTZm8wZ0vrp4almAHGEKbiWiIqajcD9
laMkS9UWVXGm5UvGFh39ywzsIh/t5goQYB342Cioku1YxS7ukBVpnpO9aap5BmNe+a/PWvxiBVPM
GUxvwbyvoNFnfO2KGOky5pI+cQ+yEm1dZf+9g1Qxj1jqnQfUXrvtjx47T1TS6UHIF3PhllmH5VXf
6epfoOYkRV40nXaB5k7AiSq8frfQxWLFYfJeAumknAyCoySkjnXfNcJ1U2ElyKNIGd3G0brxowTc
vLXedEhMAfN7CHOc6P5OoY6gV1op9sBPRMzT9cQSOCNO+dBt2FlG8Ex4TrXEY0gozaK4DOeTLFVh
RA33Cx13D46ju4rhqR/qHZdZ3Zv1bv/H94VSBdo1h50348XIE56crj9/6Fddm5ousPNFfzQZRF70
ptC0F8GIQ8yBaIR3Z/jBtkDzNT2bbRwRgtiqExD/nML2xUpyeCewSuaJCp4sAt9vMYg3yp+3MK8L
1Szck4ueG8phJs1vL6+Zz5gPXG05fLOVDyMmplfPXSKE9a6ws1XV4A+7+cjZfogdyuvg+v/DMy5D
bFnOmmuTU3Hj1GB4bHKvshhq5tt3UmJ/XnZJQ71Fymi/GK1L66NRY6hPGmeXTJLxKy2KZVAIhwW5
0pyskM1uguNxOFDAkJObiEMWT+qzCA7cfz4ETr87nCnDt+cgqQK/2ay6JFAk7gOZHFEvz4XGO7ok
kiKgNb/ZNVqoXz5EGl9jcWPWIp8Vmq36woRkBbstyxzqlf69WG/6zXZDQ9Xo7toQA1pAW6Nhh4y4
9MYgIv/BicDipRUpkduwSIVB3T5QlDdgxBIeRaPRRTiqJeP5yDwFR+O1D8YivxN/sIvRFNddpPY2
f0FeKUff7Pq+aWW1jFDICmuJ83oleO8+kjxOYj32Nia9KgQxti73mMmJM9dymgnSkiSIOE6h4rKJ
D5j22A7HaekAJTq9L8WXOTQKANMN0B1Wr/a/lLe246sajdIvL7eWXmJOdZuu8C8cSkBHg3lJ5yyI
TnEjNCqrSzvCMv/w9xd6JHBIQ+/GTKKpdld0FUKim7mAr06OI1JTnbHMhRuW23epG+Hkv/4xeauN
VM6LS69yaALoBNYJ4fq7Vw5Q8J/Yur40H3ABBEyC1JcUWr5FxyuZ20/WhIbqvLoRtNd1UE+0Zpp/
3J05M0aU9oMnkMhx8/LsTRYhWKa2tGjE92nyqqDIm3rAHVvip8MKHKhaQKUnzngjCCvN6yEuB0/p
6EBoWheXH3eTSWZnhhud9VkAmZLjIDlzAlF9KH71DDlfDeeQJTUa8p+h/VnbSstby/uofSUvBXDg
QHd39kQF50pou6kfRl5j+/iBzD/hO9xMXbeGiniizd1HYoL3JnKAgWQz4z1JPohConCfC3+nanAJ
DwSodd1AkUo30TsmWomgKggJhwrdvIfGqfSRTcYx43q5pmeFZY3FmCSR1wrYnEQ8273WIfGIkGkM
LpcZEml1MZfH3C/yA7SJyjON3b+jWg5fPmrMtFuJj7DTJy5l6U4FJqQEjcCfFk0A54y6vV2uQ1HL
b6gvTz8vzeR5M1LohjRn++/E+Fc7W0RBUmhju8/3BLs7hdaCZEod3BcSmXO3K2Th+UbG5aNAmvv+
WbJ87I0abDKJPYLkNeP8NBReUgGel4T9DIvmVGBf65IgpLycmRu+GadyQXMRRBsCcqsPYVfIWQ0v
W8nn8zCgNZdmFKxIbAy9kxMYd1cs4MVmT4udc6HTuLBeNZucNOdArX9jdvYJ2ZSmaHrCfIpXZPdb
4Sax8YPTwq6o6aPfljzfwzfyHul8q8eFCqxZLxuSa4KandudaQeXjzDHfpreoIODZfyzrM0gBTJm
mdt/YPYP7VYY0hwcZHQzY6ENoGw0phHmYCP7AtUASAeZNW2/7iCiORCmUB1OOYpS99bnRFvy8FyA
/K27suEyqYNdKiCj/FOLr2gop5v/7PizkpFecNrEYvfNOg5WswuWZ7uyKrKJJue/oVewVPlUzZEC
023e
`pragma protect end_protected
