// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
W5PhHYykMHhNqqiGOB60I0TvnBb8HGu3D6T5IwviZcJprQrUkPiGmK8H9g3A
NjC96QKisNPMVsb6N/Xz7GUw4zWrKMmmwORl06guiK3fVEhituDJ+Kb4TWq4
bLuHStnBznwyXQpSE8z5yOj7OQvcOJA2F3cuN6QBnrsJm6zup4/fyS3cZ+3f
jCwaNZrBkNKlZmRF4MbbEhFm5OyQn4SNe3J75dKDSDxBgLwGwrv9nt0h8CVJ
SLyg53WvHAZde1Ce9cmptboYn1R2hCvR0tDXi2tIuN2KwrPprFRV5FySvhBH
wFQyaop9ieSAyA2shP0feMSLCJ1hEQeqhDEFp0b3rw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
NK+AiFXZqfXvAF8mqa8ruULVHfdLtiVJOFolaJL1mGle54EU39uDRTsaChiy
ldEYTmPD4zQxaGKnR0x36vTWPyHd4QsPjLLw9xvhh5otOJbtFdWpRelQ+kRm
PVNE3oeu0qbUSKNUl0je7KkakKHxYpxjPJ9LWDWLioRTGc4R7EiuGPQPeYXA
qV9zT05wIL6n59ZiGyMYMbS2TZBlm7ttcpMwVzYI1poZdWTZ9Fszmhk5Tqvc
s4WhojJwLUjm32LVSLMiaaJ/kzHZYFPUzuyLrdUXiGEqeDg6BRPdJ/V53/A9
Ku25Dr+BZo0Kixw8XBbqtQp3Qh6vOqys8cloe2tffQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qvRxFDFfSpW1OvWuGIJ6XE9Hjzi12cIQH9/M0XJExACdT80Tiw1MQR4jEDqh
tNpTw0KYtPGhxzZ33+HGk1fTRmfqDngvNK02q6iS95NS+lZ6D/nGEZeWhpVm
DCjVKiAs9txrkVBx3dQWKOSIU8InkPlGCQrx+eYrPKuYR7y5a/ICMqSLW1Er
2kBuKGoIJPm+1FTEsLCqhAmjFIEXwYaJvI1Z9l7iowGG2XWhdiUoOnGCPqJt
yud5s8eunAAx8CYZ9Y6kMp9As3SyrJtC9nKxArMYFZiOFwGhdt+ZiO4JPz2v
TKXo2BdGflKpnkjINmpA8tyatT8ipbkKTggI7ZM07g==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
mQWB5Gqa29H3paXVTEi08flL5/l9U34qFVDqCw6egFyzKMl5mmVmyIWpwT8d
7yQ6xC2jYCYMCBFd3eAY6loX7HyXqF2MWjVLzisixOrLZC5w/J+9Qx1Cr1HS
2qolFcNpTLQcVpOAzKuRazAKgCEqJ+7qohnxJJLlAhcefmd+Hjc=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
pSBt8eR45SSuNsVRlpK/GVhTZcPBOsdYPxS+xnIJYnXhlk4eKp7IxTYU05ZB
ucT/RqoEYlbXNLUlgel7s4idsiUqgoC5VoynE/BUL3kkFN+qK9HnSwmh/0AX
SyYsGLNQoM+KAwAIKx1HmR/TRfZshRNGaUJDUAMtXhqQSz957Oux5tFGPRRG
i0gRc3GuznYy3r+sx6ATrXdpYgmGtvqmTbltC0LaXN8sTBx8/xiEPjatX7l5
ZOaB0S+Ge2fBTdUbfCW0tJJs8hHOkwYNHGHFYWbMbFVotgolnSIJM4H+oLzP
y4DBdvmwaVR7KIy+lU5qeeW9zoWHXMa4BUhAuSSirO6mRVqRDITaCWwEFUnx
eeEujO3O1fTr8JKMz9wIzOqu3o8xAhE+cLjX7ay14VrWkVoN14KVEaGSAV4z
dWgzq+sURf8lK45Ct++VFLe37uMjUfqn8wQml3GtsktvmVeaO1mkZHOI+zXk
ts2K3aZf/87Vs2vJxlZZyjfEm3VCUSxE


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
XCge+jI7qW7JAeGFzMFNnsJ2WIFInEXm/1lh4xBDsnVQ+Dp4RwGYtLPfRxK8
tcY/cZLAVQJBsMU5S69djvwFtmKPNbzLXB5vOxD8+BCqBggtRWtph4E+DIA6
r6fWSFqIjoYHeK+C67iZ8oyzCDoUJfZuBIHbJu0ueB/b+pdqsTo=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
rV7xohfpfHsvGfAXE/QFYhIETJsrWGxF0FMwc4SkL0ZKCjWIZjDV4d8GxySc
/jHCwhHtKq696MhDKBbGXdDWpdlJ6A/dSPK40/mGoW+5wUbvEbzym66yR+O/
dJ7GUgBVz5UKwyR2eZmQazj1HdXX85sxas/chJbEutrj+GzMHDs=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 27680)
`pragma protect data_block
OL+mR5skqAKfOkDwUNl4Pbb3R30JplUyqUf5XhgxuY8o3MIOyb3H6TMnx27W
jRStYv6KVkRj8wsV6O1DYYnAF2fF6seb7L+zAb7qvE35MTcLBVnbZHMVeioK
kmKMhtNVdELYJMuW2gzhXV0fcnagcslCAqJHU0cjmT6vFY7FG3cyk6V+rP3E
lzwHMRgLtHIYVCpgWBQEIUdQ1R0HUAJs2WZOaqL6hp+EHXWR4Ta04+1uOIgz
zndE0mJAuPmj4/dbXTiWRNRbWfz5aEU7VZs7Brp/tuZaBoik2vEcuKI1W1TI
FD4INrf14D/ofZkiu0d2kgIevJptPmacjumIN/eYVTrnS42aUF6sf5m24MtE
0FJFAe5YktaE0oK2DzVr2sc3LYL1sV238vSxUPVW2pVSNMHvgxUwxFrd+lps
T3q0rC1PmsHwijFB21HJZFi3Omz34BnoIIeHTX8lTGiVEP3waijXtDrD68Db
h/KVee9X4UBWAfk2G/Ksm3V7lwbYACxvWjelEGMWBPHBaBNv2IcuGrKdJprx
kpbmYXR9ZoEezNEce/q5BumaDnbe98jIiBPUdjxYSPBcX2F8yoaTd+5FbZdO
zB3cQFRpAju4wpjprezRYATyYH/QHr5R2TjPsLB6q6q76dwMLCTtCJz7IcHX
fx8wWTTn2/0Yta/EvFhPakQRBKclTOPdQ5nD558thUvJW6R0rGVRIGGacqfZ
Pd7ar+EH9mLO/ZyPSDDb1b1hJ3E2unTxvz/uHXVJsiZdB3cTI+i5/atvU71S
SwbWw0UTY1cvHmHvTj3EJ31TCTM7ku3SAgSMDtOK9bNNNDLLs0pC4AUIY+N3
qa6toJz+lyLog7HUMPc2SiawNa4dOw1KsX4SQUlCKGwYQBHjb7L58FnkXzJb
s+gFPSeJ236N1wkZwRcpm7eWGpOMyKoWAkKeIS6k9OmtIDBOYNDS2KFnvP2Q
wDO4KaWGzw47EgQZgrfVc3TJ7DvrZ2vjavu8oYHyFyyBWnFVXTV0Bi7kZTsD
CZv+fgx9/30OzHLjA7fnehSAyZx12OvnOwjWjn2wUSfMTF6Ee8sgqZPvx/CF
GjVdxnjls/Sevh+PeDx+LviE/P/87kwMOw7+Ko9C/3qTLOqKDHEjOoqJP6QZ
n2FgnHjvd0inUiFpIqhcEoWWikjHl+AdNWV9Ogu8YA9dpI70YZJD9W4ZGK8a
tTJD5HBr3Py8iC5/YsPAPmNczuVVV53z8g8eKPBCNze7VVNmX5/+LTKCEjZT
LWpFIStatIOp7URMHp9uLk89GoYf5Sb5jsDO4CTlREwitXtYGk7XLFd/fqFN
lurBV87XerGPGePK8H/KrzmVnRCNnAZEVWEZGTlGQbOmEeBIAGiXMY9lF2EW
RJhRiqBqR6x5di59RXf2zKd4bBIhp9+7SToIwtd0ALPDvwfglLaFE6OSdh4M
0MyMK463rcqneroKRDWLgj6Wd+/rRt4QHQQIUR942HpTljDo/jzRRIdV9g65
j+rtCz4NI4OQvFerYbBJvJHcTdmj5k+MOctwGq5JsW7a0gMBaWB9AeykNCDS
3R3bHDiT/7OgrDEUoNUkeq4FwpaCdWED0P5zHvj2IfrBCyyQd5to+ESLQh9K
5KuFeSlkprj0ybqEhfK5xzuBsfbYPHuqmQErBIVcP3VjF/EZ4pAmnFC7rbXH
DK4ucuGXndOixzRC+22yeqDXLB0LyIz21lKGuhXJdnZk8k3ChpaMlDNa9Ufz
YMhYLZpr6l2LiEC4LLo/HfDdz60iksTt92L+fUAcIMkOI3Gc6tRDzUyp1iHO
6QKOu418aofsrglC8fvL4HRpjnt/hlJauO1lRUnnrjhfQ6S6qLuDPo0y/xO1
AT/9f+wNO2WHZzfVqyTtb292f3t9N+jWh7EoN1is/fUkKrGIgllrtOWDqZSm
nB2E4DFbknGyR7/QSckT23oo3nJ0LF67Pa1iZgWwZZ2l7GnVshuMfU9ywmuP
3JGNBn9rFcERqL92pm2JwZ2maBgPkzlEPh/M1M57IrPAXMFfDBGETBGN58Vl
7Q5TdxIE49xsB9YeijUgl4OGQkVYdmyi9slBHBSrDkKJnks2O+SGlIHlBUcH
L7fWEnSgj5S8wdgn/cPTgFBVfH0BRseRS/x5DamGYVDNwJwIA/WiOQy7GX7E
RGKu03C8mcvxVW3Xha79LEC/pYLLtQ4Lthukh3dSTCjRU7BkMD5o/AnRrinq
Bwzi5SDvYMatHlUcbmhn4Cmxg3os3CuKC45j4M4xUSCcrCPFoY0TYdXgt/jj
j7Sdmfj3PeMjyWrbO1b36A8IQW+4Ll323AMoJ+wazReeqkoxJVc2we1/o6xf
tu/tZvpljfl3oFC5QSyK62UOqQhKf7hRI5yVNOdWTTuzHlbyr7mvDMfBrTU5
jTBivdfMgnTB3nLnkXmf4dov119Yswbo/xrffPg6hPjpmCq6kwcUTbMiSudP
jo3d1091e8j1GEPIzTBx48uT2bjHQr2GUj43088z2XHe94Ne2lb60w+XFi2F
T9vDFeT2KZBM8FQYFIXMuYrVE6zHM6Kvk5UXyQnuik7H3IikLFcmRp23V9SZ
nZKKbiCWY0V858vEB/e5yUx7GQkiG53KGaZNkuVjyRO3dEDh+B1MSdf1buHl
0TaEzhwyy4GA2iXxwzTgYYjqGKFMeKaecnisFkPh91Vrljrv/bpI/B3e35IK
9axhwDBHWnm74IMYMLUjeaGnafRtoWpeyjYANTiUyABFKWJpEotTzQIwdZZe
H9ba0SyOO+pmSVxAY1RkSFf0eCqBztBR2zLUubyzDoBS5M5NajTznj/s2kjY
EE3R4ZtnSvOmmPEmrkov4Q2BqOv8f2jP6bABR5Ue0q02e3qN5tpjZnwTSkPw
LgIjcsES35cXp5HQEEmZg/qt0HQh1vIP4M8l/+8po6cfB4tf86suJnBHibOl
yu/83YIUHwc2IN6xyfH5NiWkTQTcCavsgHzfISKpoRsEu1SFcPrMhWXzDYLx
wmPopkh7t1IRDQusOn4Zct/+zxTxv9AOiQeR5MPN7CHSNtoHxd+z/RDa/ECy
lNSDVCqOjFQKPgq5/I550r4hfPjBGy7ONr+PAkrXByGCKhheeGUoMssgFrYo
M3HP3OURSd2YakC+Ykh5cuiFMtoMb+tg8R+p9lcwzxCUIsNgxME2xLfo9z2Y
ViWBclAIBTQnr5jkHGYFGuh4hitiu4kDGMGCbUpSQOP0J2vbvDd8AzZ9V+Q1
8wppWYSODT3MUOzO2Xdwt2T6QpBuyveYGmD2lZl0Qr9mB3YCsTPxkdgsoGHx
eRcEUI13T31MKjLtrp6ZThhx1VfRuqacrZrV3RT8D8XWawUPF1MGevIV70Hh
6nAIiTvYktnMdpRTOpU1loPnAIW1AXiive9hPoVa9mfRgdf8btjvXSOU+5r5
8SWSlGtfSapmE/0Idfwga/daf60f0mKAOIVJhsGiUNKYV0sQKnkBkDGjSTWU
xxn6anFvj4Q9mqImbP1nYGlmDUQVKnkvgET2T0v6K4rwpkp56dl2G8wG4Ugd
20+YvwVA2fxgdTWfetzws4J04x1PQTeRMtPL+0F6bAqz7dbt6mPZ5ynq4YWm
7TBipBqtyR9j+MQ9RDvx7OiXLrkGOyXIJL9MbPnauZbC5FbxaWgXKr5gJJtz
Wq2XyarS5LxuAcdmGQcW9BlaDHo+7uoZZyubh2hkiJAMv2zltoXqDrOiT+HE
kNezMbM60Wzbit2xtC7EdKPEiA4VY8dSfazNPkIeFJeC1DGQ+KBSHdlJ0vSZ
3XGTCyOUWhNPgYnj94N4qyQBRDY/kBKadY07X8HV/VLr4UrkSzkCTRlvSWIu
ilRZE5iXQqeVWxfL3E76wafvMzw4V6XoLr3pCWeKhyE27rGW5pa/yNwgtzlg
tlF2w+cYS5VwQ5CaSb4wSxgl3ePNENtYMdC2eC3Cwm11LsCSoc2vYnU1Rvnw
BRKo6jO58eqeRsLTEu01q7GgypX7mfW1Jc7p+DTJcWMn0z6IMIWsB+/zKtEH
XMO18GptPjLePdWGN5WVTPdabeuJemjAt+1SXhqEpjBRdjANlc9v3CJkwfMI
LocclSaYgb49Lgn8A5PxaOgXEgL6QDJQ5dsXhBKQm535cCnPJeQez7T4gKzu
wwWDJkdsrE/sa7an90w+AbhN/sgBk/qyGyGb/eeEMN/apcdcqZs736tkB0J+
r0SCnyPBKRMq79SzjoNa25jZiZIQ+9Ex+4ypwLHGp9bRLg05JqDeqnyGDo1M
MJGwbLEY+oAvHequ8f5yBMNbVLwHXG4lFyQo4nBYr45vM57tj6ACQTI1dplw
cwvxju4WHAh/rf+QIExX9jDzTLPL0pHj5n0u5G4T4YeCVwP6Eb27G7223i46
O8q+imOEdhJ6lM+UfC9Mu2Tnr0ZyxCZrCL354v5PoKV0qOHNZ3J1wMG5B4JC
7R6hNlRzDhkDamnXM6C/6r5S+wWz9Kmhc4odqX+OcrgDa0HySnEpKdeU4qaN
P+2Cr6POeh4FX5FuuRzqKSPPGCPxAPPzdMjSWiyZhB5bXpR3iu6SPBWuV29Q
Kfx14rZrpP9+Re7xxZoVUjHbIrFXgUE/u/tLhfOFRplv+YM4InD4soVIEWfw
ck+MgL9vTp/LVB+mNr8Wv8wQMcaCvzGj+nm2iNEarnXq1WK7QyTONlbfzdzH
X0QdWUuyERZdYPUsL0AIQhBJJV90uujiBjm4qPSllUv7fdl2wlzt8XCvLchw
yXSWA3cd+dHJsNwV/2xf7nEhswdduo4yYHJu+2VYyXH7j5E21IvLAulYMjXk
Qkld87WgIhHZXJ3lewk0xuVzgPCjd1He405XnEoiJoehjcoCoJzX0Alm5QkG
PjBnIenNECctTIwSSWo3cp0w76vqeSO62kZ1HjiqbeQ3R3XvkI5acLVz7Om7
d1oiu1Oru84W3AjhVlMwPFHuXnbhtrYOxnB+Of34w9N0yt3Sf/W7MZK0cHl7
hqLjHM2BYZvrShWnpsEby4O/kyKEbkEP9QctYlo7uWBctqsApAwfthCouwqY
MKnKStncXr88ZBUGPRDV3Md0iLHyKlXmlUSvCjzAEJq3oZkGrfp6fLsABlq2
MGtdBGH1xaum5zuY+1lQr5ap3g4nu0dxKlEg4bhKrhWUpnCly0VWOfQiaeZx
QHfkaC68btdKPEGlG9hkRDWru6KS9+R/KatrmB+e8zIU6h8fbKh2KAlu2naj
YjmTtAyqxZOF3NrUaNKy43IFJeqlDshgqClig3v4Zeg4525EylXHELE3BrWS
2gOPDciNCslIGDdiJFdJnXMnt3JZE3tFZIFnGVwP8cgwty83EfRp0DAIMbJG
VLEK2PGfDWok5NbrRfFQdciy56kt7pCI8nRrfNJZF495GblPSovhTV/i8mxb
JMcI98BY2qB48j5nfb9MM+SLE/7+wAJcAA9ZMl2l7ktH+5QXii7ghCifpWHc
y/JoVWoPJej7LlEgpwPDDcZrvSRi2g7AjyNN4QUmqBvoIrjUceQKHL/fiABh
HcRmj5Nw5XdJ5ga8REoQDx0wBGIjCrcGxdJghjvW0HW0N5dpmPuZWp54vynC
wh5UOcv+yo4OBNniek202vR4IF9y3X8h7PP289ppA3YDMoKuqBwaQw0w5+rK
OYjaB2hBCDcEIUtOP8KArxK1PhZJwCnQ+ZhAKhKwHsv9kFgoGnYmumHJq/SF
P3zY6Sj+hNpt4If2y34HrNg3K88TtG+MHA5tvvr61sknUbCCW14Y2mGA7TWk
ml7GOUABi2EwAu9UGUlEu+AXas8cnvODjwIXrRrn6djqzMLC2s9VwQAVliJQ
u7bx38N/elzdGMVLX+2bt18cgkwWfhgCbGx//68mtzi9fjI/c+6c1ApZzYbA
C1C6FRNL7SIUr5C4qidb/URxqTta3vi6SPtdInMdxaFDksLmvhKFKIfkLOh4
MOt55Ci6rjbIuBkojdgXs+CdEaJ1LK8jo3LsHm9TP+fVOCDao4cybKWpiUNN
jtPbK6uLEkhPAfaEcxrzdk9xzJYINOhdalfoxF8doCS4CJKytDtclXoYZqgj
B0mkxi/ECsY/NxxJRLffYmD8xd6hHh1GwVdTxspDvXEZ8DIt/Y1ba608PGUB
AG0tLU56xqFJDlmSoYQSRjfPlRSN3O4c/Ir7l/6+WG7mrjIcGKiWrobX4nfU
PlmOWJGyiFYJrpqEeXNqEzxcknSsX7bPyDbwFNW+x3JPCnJ/hZe2IdPUH9q+
6LRY9PN5DUesyndsCGGhFwFOozChY1q7dOEGiH8xS1OmRL+kbQoojb6lrMM4
55a1eylYSK3QodJXm+yWQkPLz6CziFGSRt3iBXcSObJN//6v8991oUmMGSMB
+rMlLrgAoinP4QlB+7GtCTF0vz9eWOUzHXRtTfgNTw0KHOZ5kj5IqWg1qvfw
TNaRfs7A+OpmbbekPMCxu/6hSNFHFLaMPU29TafEI3juze36A44pexdvPuwy
4XB2USdqJ5dLprmiGuZ57NaM+CNJf9GaEOpqH8WkHwC+fF8Ak+nkspJOjyPe
AQ0MtRCadn4OIJc1ik9DymXxZkDbPuxJUCQTDgdTtB0NeSuNPIQHBnNZnUPg
kS4NaWTTmsHd0aDZ997xrd0I/GLFZr9+4SNSQwXHspZ7lMAE+dqyp1ugZlIK
Pg0Cqm673BCFuNuYRgQ6OUxkbU7bBFI78jWcBO5Ccc9jrJc97YwN3DIlWDHU
IjPgKANA57ph3iMomoUbqQNsuBW1h14UDlsY1HO3rmemCr96X1oCoKU54Dyi
YW8avc4ICOxye8DHUp1EgYeE/aNIYw8lneZKHc3BA9VoDFXU3L9TMCCeFLws
cJNjwGQdKJDp433kpD8MTWi5yJguxML7PaOz1twDDbK4i1D3XlR6Eg6GuORv
yhl24dG/fAdRAAsQnO3B8sLNy8qT/3ZZbGPFv9ez7LmmCA1tkJ+KM3fQzSho
X53BhEgT0trN8X6u5Qw8X74fccpRd+e2nAAz3O86mxPozaoQTE+lRX/JjgDh
Eqlp6EkAjTlVrpLGJ+GdD2K3LOHkPAA0qLzl280AbVu7Hvep36vw8J++xk2V
PKC4l0LuAfYqfHleTArFW5A2FJzL0rE2gwQ3uX/86FiUGSEQrLdnIDByLBi6
Si8pbax+3ttv6ob9BZuOHa5DTf+sVl4RcdRa7AUZyTUPpPxRzOQ3cMW0CoRr
WwbsbCOfVNt0RT6mshmMncifr+QCrAe7DJUN9UXl7KadIrodRb4I/PeD1LhD
rmxz6R4ZYLyRryjsL6TqHH4A7UweYlh7PLXomoHNh3JEvzUh7krWBHViGFph
6hp0YEDBMQ88vSM1PS5BSBzO3MKa0QCX+LxB45iyUwhqpSy5BShiCEMZIv2Q
CX38M4VhjebXh1OdPndunHWz4UATFlR0WUYBfYHfauxnu5LPkB8QlyQ9JQ4S
KJ1nO9AUnIj5YOWh9zo1IpzyoeXsxJUG6y0hzzKbjTohOzpdmmLEQ0B5DnS8
OlFmUsJYsLtPjB+z96pTNa542k7FBHq76dhddEi+lKuTL4ZroEyGWpu2YdWZ
UCuk68jKrjUftLAulDx/SzE5ASv+N39w4SPkxcy1cc1lRyRBEsbdxfh0Nv7A
sR6ebTtO8UvqV5W2lNDoXIVMr2WhEmFTbkbBMKmAB5cmWXGuJL8F2/CPnOPR
EWDPN15K0i60aVRJC9jrOUeqAPK9YC0/3Qoc6Xd2NpOQ19toSQNBsXn+cS1m
0fXNJbSBT+5UMFjC9cSFFEy65M9ZVAByxUD3hjMxnRgkx/tIf5WZ4Arf6kz1
2wVujfIVorSJ5U8Nuj3fGe9OKPTbZqXVK2HckFnetHxgCXVnOrzgf2jy/X94
vyFLeQ6JRDQmxzYW9gXMYnW1FRLDFw1K3otJHMzrPsqsbuMioSXQxVRQ6Bn/
ygGgzOqozQSL7S/R33e6TLYSNBY44h+7qJC+RqDLVZplYAys6hqk6isjU/sN
Hfc57Ac19cRGyfxx4GqTk1mEP2lWAQPdiTE9A4QpVsemxghI3/waqaS3sQyh
bVk7BR3JrMGIX8QM+3UHZ7ZxF1dFZ1abKF6poCkC2edDxmdwsun4V9AsOSgS
Yxk+IGC1ham5psAEaKvY0xxnqZ/8B4aJA6BIYHCtbsE4KUkqLKEr3GCOKsVJ
zVQIfpjmNj663yPRK/FARdVkGV10mj5oR3K+GXhRt17lmZkuUTVmEjUTkfhU
8E5aJ6BQDdadBfl0kPGGMDZwW/VQjItd6Rpoo4wcQhRMBAZt0sfKU3wgSK/0
/Fmv00qSW12SM5kD+GHXhe/9CVMac93qpD0Qfys67pNs/IMAd6/jOZCMLQGi
JW8/E85ZpBElJAu82XC2PSZ6egYic6be+22HixfpHzm7rShPoDgNPGD6+J4p
4ik2F/dVuvXTC8dGN4s+vTtSYRvT/SyA8y9ge2grGll0Ko81ThXHlw5yuljz
jgbgTKhzSv1dJN7RApZJcv75gEq24tJJSW6alt1oW/ITcP2SuQsOBcI92awt
VY2WzHZQD7EPrpd+Dzg63UyYbM/GdvG5D1Ilf6GhGTawY8vJSzLIZBDdQGLI
9/r742mwLIGEDdVSeGH81Fg4Sz+ozL/+jdo1qmINj7Fk1MRvFKAniKTxrISA
kpM/dvhgedaYBIzq2XD1yr7UPEXYVObF4rbBxgMgpY1kPmRP2kH7H5qjI7HD
cm0e1OIZiDa6p1qX4TkLc9QRGxOXn2e9yB87mZ810AV9gi43Dsez2KHZE9cX
kTpgqyK6DuSw9aPJnrQoP5qciAjKChoRmuoxqTJw9E5ajYDRBW3M740ajUZc
EFhKnFZxAjBZWGN2Xtfk05+1p1Q7dAtXGZbM5FsDDkwdGNpfEG59+y7DmJPL
5oTN3mSPSG5sGrRTnq8zBZV4LSJNVFlVnHcScT7PuXqx+IIHhrPa95cqHsnM
4pZ4AayoTs89I6PV1TbPsik6IU7ZeWJkjjSMeJrgGe5pUlRRfDb1hVxicl65
nUOm/I9ySam2n+GCqsknt/nZZctsvFZjx2mTYJqRbTwZqZ8jCoimPxAnYwaE
Rdu1n8zuwmCnuY/vRoFzyuMOTXgviVY/zG5vks/HtG79kWY18gukpkexj2OT
EZwkHwdXXLf3d3YK5Xc/KGGfAcGHa3ho0pYDS8IW6gGuvLKVEVNuXfVSeGyK
pMRgjqSTsS0k60P+lNMUrM9VFEOu1jxVBvqblBMCU/bUAD0dlpGzRqa9llmW
7y4btGbqok9xCSiu2OAJjbxAL3HNDKDZ1wFQH5+tQsOHz+JYAIuOtFLXCd4M
MubDYOfDEwiCteguUUqyljC61uSxGIYkt9qUtyZq6Bf37Z+R7Orm5+TGObjA
05z9ajY0XCYEWc5rJlPmz2LfJ+bgR8UR7RJhjSuueZE2yZgvarUdPSn60GZ0
5wes3Khk/oaUV1zqMP7VCKuCAk963z5DK0xzw5Hfpl21hUkRfNen/hXtoFUE
crWyebKl4tYhaqjJgDPeTX+DKR/CbU4tXusxLGmQHuAR3b+PyCLvdv+7H5/G
8I3nDsVewRO3FdkZwsOXj/ljakdBd0+k2tuc/lFc1s/ymqSJGWGaps1i1TfL
D8GxV38BWnColdIFdkMjZJxxadeYw74PVrBvd30JkKT0+6AmksZ5zXMcyPDa
SLWBc0HtTQd17FPGQMOKCMCT3VmGOHs4RzmLD4GFncrkdIkcMauAnp2kir/l
wYDxzV2k6JxM8oRovyMjKvOotxPLAvsR7LNvBM7Ygu9DKU9wLWg3go9W35jw
pWvTCkbyN+y8vcaTS+Y9OsgdUFjaz4FHon9gF+iUOZOt07rIy9Wr9lEYxG9E
ZBRHiPNsBehi/Lac2ov+u9eHWl2lmJ6MDbCUx/sYLvQaLZGsWkSUwdEXGN9y
M6YaETOEvqFZ+pdlpz8ixBL24NakuqOgBAAVyklzVsrSe9I+E54sZnkAKtMw
eTZ1VHdsdxGdxs6S8vCgFCNq5rSX3T2PB3WlLoq1eMrJB7cN+lvmSDLVAbOq
1/JrEeb2hlsl3DOQttpaRWvNkCueaC5GrHu5QGmWY/wpeyr+h+tal/E/Ax7p
bTcOGof09qffxJE4YnqlWPKsW0aKoMIfsgHNv2xgCOA7AhBiUt0p/Whrmis3
geO/hGBiynMKe5QhNiq1By96xnlOujO9R2HM+2L46TRu09GMwAHh3DHwzEx3
mn2ltTWgHtA35mKdH8m4m4qQItHVIjgMBVdUARXW/3BftSUzOnZpjoEA9iTq
EwllrVh1tf3UzM9E093WKWGfCLWa2cmjB+J3HLma7HsExeCFJPcSb5lD1QLZ
hnJQVlDrC6/TZ9oCWTC+T4o6n/IEi1pfV6Y2d7r03NXYcTf3eBjJuJzKX/JQ
cgCsp9Ii4hZ7jT9Opi8Ke4RvoHnxHrJOY6kMIPxMMWWJGse0fkKFY2YVbHQ+
M2M+kxjMm1dqViWiCZ7ceS+gvAeKxYLs9foxTrZI7L11F4SIDYlVUXssHGru
iWTt5vAyR9Sn/FqCNuHodlm7BDafqCPTYz9LUQoQb89vTH6ztQdO1YjDoLp3
9WNFyRqH8N7tZntLWAL+0UNUdaUYey4F31y9kwFac1r4Kg8o+udMKgikzkP7
EQVB9A/5N8e8Iiiid2JOViRJs8DW3nOcuVr6KP+dkMcrA++DNA2vy9+Yk2ux
sbsX/nCA6S1nInoIaTjljX/swbEH5vD14MR5EC54eTPzXO32VB5BYSgRHrDM
QmlQ/5/0S/GgChH92k0R4yJ5YbnzKXu/H1DLIqTTslPt0qr8vm1LZ/wUjd1u
RVNTuyhaxuw8orpwxoADpeedu+AWGMdGyyb7roqfO8SKTF9cvmRjjlPP67Xy
DWtv5mzTCYZfNHQHS0oSQPKTogb+RF7e6RsKO4cHPXsJPPn4luM9M/eSnldN
LL56fV6+B68I4+ATlG1ww+p1wsB+bEIvcZ2/E4RLacEZBE4+M+FEEN1Q1BuO
s3NSomNBRrK0RH3GPUealUNwfdQnqUsaq1+zSPB5s1laGJ15GdLxYf+Tia/+
z+d2T44Ksvn64X77w9V2itVXVloO7sVW7o/hulHrSFj7Y3zXdnLYcEIiqfA+
xFz5ISah1kKG1vlt15OE6Y/ltNFgoIizY/3kabjQry9cr+Nh4A35bU2THUhZ
OrAE563FkCQqjFhffNOSpmRlFxS/GqBTZDrEp7Mos4i7NBAQFyumAIBIt8Aj
PK1sWypHkYfjsaMriYbKU1oGKCO4HZPNI9MRN7s62Kk4YZyhOQMct50p7RA6
fcVrOYF7mlkjC3t2Dju8SnZ6AkKOdhbq05DspuyCueStlwMx7iG6FAoAC2LU
LlDhznxm+CXDunApnOaJ8U+3+oxGpiSefWKiAtctT2ki40F31RAOMiFvdZpG
ts/XtwO3LWYflug/7CN5A/YzEVymj5F7hjkTgXj+P5nuubnmas47BZlFKmec
+kWGu8H/U+teRuSy7v2w8EhBEVitkh7r95HTo8MzhUVhgHmskzY9248o47tN
LK9uZOoD63r7aEhHijFd1/NDTRaLNeDOLsoJ6BFc1flO0boCPove3PBSZELb
ueMczE6RY+eam9Uqk6O5a/pe6LBgEdwW5WwAdc7umYuzWXsruNLDXqR33DV0
LzsjtHY2jlaFkFTACU6riRt1uDpyaA60NMuhbNQ/uRmLYs28texCAw2d7e/Q
BujCttk9X0q62qzXLnHxfKvSwP7MhMGatkJB0iQWVhGwhbna6x2WGhq3Slml
9/xTYjLsP2upT5zOPVaGw46LWHuiQqPkroRodtWLyHXVRV9b/S+8bScA0tuA
4din/uR/YS8dHNcxgLMeleStuu5uBW7KxGEx3zQolooZFDQNZkVi2pUnURTM
iML17qb0+w2z3akyTdfycXvBJjuqcGi0wxqfx9dJPjbbS+seDJt0q6lnG61K
5R6o0eAyCOKgqXumrxS1exZuNwV5xlW45GqVK5fAoaZ+kkWyMB3raWCZGEX2
GzKRmGcwGyVLrDpcOvUZhR/YWEey0t35lHGaDe7rGpc6WcWitxsulSqiMio0
+wKeQB6w6gGdB3DFk4FQVhRPI7Ssgcy4/SV3JDxDgj1kJZN227GpLUJ+fwc1
gcFRfLIZLq/1TfFFx/Maxzt9ZGIV0E4pTnJuQfkBo0v73fTu8luGJJaYdFUV
1IlwSh1JBQRRahKlFXp7DlSTJ9snOqFwr5eurd9ueibLQYr/1lUHLZ2ft4vO
xzGRyqSW0Vw1OCcgF7gMtM78CFAmhbzpAfF7TXNuGOMUD6iH/V/fH+Yby4fs
2XBlqmnRRKREe37rJ4Y5qu2U0T4TtUoX6c0lC0F8/01YFsUUikBNVRYePjuS
2ijfPxa6cvKyuHD8rsF1dzdJS6pbJMD5cDAtzNEuyjepOwpvw9kMLp4SXW0a
7pY9f3kusBJCk0vXVAZ0uSA4ETbEfKY4CW8URBtg0S2ZlKZTLjfkJkHnchtp
Vb4WuOSoJBELd/WoYiryV5a1kcrBHXdNag/6E3XDq9upY2Zj99Q32rFmyw3d
HpuCQbAD1WK/NVRdCbhNvlrZ4yEEdivZYBMJacVCdiHza5SP0n+MHVKI5kEO
9/FPbf6x3ofP3LBcDDdknqC34ELBpSUza2QJu5Gtd9d1jMjcsCtqxYiLUVJ5
nZ1f5kTc+NsszPecCounnmPeuiMW2ruGxI1UF19ZxevPQJEc6nxDRAiFQtKN
x7CLET4OUBZ/do2jexiiAf4oOOBwvovxZx4M6O01qQy7Ikh8tisS53hDMryE
uJgSxbekTi9mhCoP0WMqS155KhdtxWPVXLTzdn4Re72uesckykmMZBqy8/yv
cl6GCD0Qppcnblhkn/kz0W3ufoYQhFJ8aRdsq6qxkt5DXL06I2fgSXckTR0A
FhO85bYZDL1Xm1PBgF9WqAGp5Yrng++VFY3Lp39UPO8XlaFltz0YZXOkO9eQ
YyZ4fC/jlW7vg9aWBHjDgBcwX8A2UTCubKt2tOgaxtyvHViZQveXvTYnAj/H
W0PU1T52KNvXgqNiTGcpJG3+d+doQvGvChGK2dwzcdwjrqoyPZrvY207Be+8
cCRYvLrktbQdATn/IUdTm4GjOGry4zGhyDc707a2WTrQxk4ZdH8yAGMnvyH0
/NpcUtTN/E3uJowKpSRL9a75oDuk/oaIOqBIuP3i7TX05CV2s872oXdKvLzg
DnDq9tRDHoWjsyRAoar5DeWzmKKLKEX6wt/tpK8TBo2Yahzv2XLDUTqAA97T
f+BsnxfuLvHrdjxz0VenwbzGd7cD3YTv1ROcYSs3jOssdRyCsDZKHDTwIrm7
RUnojqzDXR4wMCKDq0OCjNRLUnjud5xbdxi47NmXeFPDKWMUTVYWEQdvLwy2
eFTqk3KPAvMHbVy2w0faPk7vUDujrgUyY/cfOfF9ttsMnTsej1jcaEbC2lyV
pBcd0m/9LkX+/6/FZzc/o/jq2AuPuoiyyyQwAhCBzVFkj+3PJd+H2B9aORU9
imh6Cg4NZ1Mdv1YGChxSAhd0TTkEo6qQj1+YWQCW+CZVGi3kdOV6QKSloFkA
Tmbdmss5YoYuHgRWcf7We9NGll8tbtX2SIOAgJYGeYmnY7IL4VLYhKJnOGRN
qRFHL/KuPCfCWQAFizw+902iLJvknm0gLhATipUM0mgfkiRj9jrfvYLC4oqI
3AGTx9+NAEqavJ97ERL/VRLijUQVKSg7zFvKVZZ3fzXBrJyfBUpQX8PVg5XI
I5rOrj5wNBLgd7fjIt+y1GCnTISasppxHmfLfHC8D6NEzqz8xF2/EVMZQjOV
BrOMgS1Pw/n/vwNoacZvm5WgrNKq3gb+n07puRFTO3iUELec8abLWGqE6spg
tzDpM0i1h32cyR8Ez+lPcylliw7x+ag3h+VrrEFE/Tp72vCIzg2yEHuNWFh3
kasF+3K+Bc4OTsTCE2gxv5+8phNOhbenFsemBJUX1SNjwjAYvo7yAli/fsFT
EY2XUjTvLfaonYJU5ApZQaTqiXLf+jg+6J0hMSSxsoAnGZUBb468u2oekgtT
NUXXVNMinHGR/yW9xMICl9ew22FIs/1wlGQAfadzRcGoCySaZwKQhES+uFcC
O2VOv/4p75VbS/bhJ4dNRtlAO/lQ5/+xrqClUGaLMU/H/1lTGDWD/4kBypFx
x7w8f8VEkA0HizIOszaC4Zbq9MtxrXoD95ZD1XRQyT/DF80K/0QXLA+VHfwd
SHeSxPBP2afV3lYujsWJoB3MIidyFdM2tRpZvyBpdUIpvzyUV7Fh4bVQcYFG
xJnFXaLK8l9XcMCetiBYWLIwI5m225f7b9L8LbNfM2klM9mu+QYpp57nRlfm
wQ0msKi4OBjVqINjHSZhpDn6SrBNPXZJqmn0LJY3B5CmMvWeRYyqMVe8GP+U
9Vhjl6cgY+EEdW934SL3Uscr+mIbcmEkXEjNToOha44Cjrztrn2UQ46hIFF5
2dFjmu029QDTfkhcUK0flXh7nRsMMmtBqfNp3Mdwfy2BtkJIBikOTZsO7s8y
cRqtzT0mbF52lc4z1WfCR/WAf1cdWxCEHs7Y4QC+kEK7H/xdA7G14ubbh1JI
+KmudrOpx91/86+unvdr74x0xfsV5+G3XYKwj6p/rOhM6F44+J4f4oQRoy2h
K7cyeRWcwwKY1aFvscO9MCo8Pt4WF5rnLnwtNf4vrwAR4v3+lQMkjBCycHGu
W5Yf+4ZBPRVj8lDzMAgEuYf8hM6VoE9YN+08cfOeWMMVi4NnyRcIBXAvhBey
HEx+zkQ075mmCGozrbWlpE7g28QY34NzSe1fH8CcnSkrVJ94R0+ZdvsfdSWH
/iEMY+0o+Y+rr4jUc/tehfdaHCZSCg5E6gVMzKOQKWRHJ0PwuKEmWgEbr6kl
/voZL+ZiLlTBUlXshH3RBd9zd4RetID+dW4bmv+CKs9Q5lSfY3Nj9XGU9ZKN
97ZtnMMW+z4sz429mI6DgjslvWX7PoXaZ9xm4HuGn49qaf0OcAJ6ij4vL4Lv
lAlEuzvOf0asW4LXliAlM/G8A4TN88yInL4BgEFGWNvSo99626Au1GkPxLaL
TQcW0/FZe7vByKf9ADaY4DFvn6FN0PZRnOU3YVE9PA9DiVa/PriRDAHiuaZm
Ygq6AhrdtN5VMTYsJu59misXXX+IBQK/9dod3evnFANNo2Z9zGKOHlf1O2n6
pl5vETjIm/0Z31Ih0spxVuyps80ULDFjTHT8hP4F+XSsrFSc+neE38wwkxm7
BRSjZNNQ6ii0ceBMO6UwGHXZzG2UcTnKOSludjgcqWGgkTQgPj79PP3qbw3H
OV/kd3uzQR+qtc6eOrvmUoBNtQsM9t678dp6aTAOIIDIzG5LpSkuaiF+8orc
olJ1RI/m1LyS/XJWIHR/qQgLNZYbzc6WABG5XPnjzgTnfN9RgToK6IHYU2H4
2VYM7+RJjfI3zGSy56HHQkh3ijm5+IBMZnqr1XX+6SVbJ3ghfyb4uNHjHWA1
klTuc/Jl/jjgYt9Yi0F9C/3A6MYaqFZOIvEoaY/jsLuUU6il77K9JjGl4fE1
OgNPZoqk9ZwHQNqGcJza86Nt0CZoC4gtvLjdCXrudeSL3BwmTP79BjIG4ISy
8U2DUHnsKY6DnwJtkhlCC6sMeLSaSvQVjZkoouDbuHsidNFn/Q8zeZOE/C8h
hfz4LPg8jEjjHQrCDmO6z4fPYyXrABsIDLfKiGXRAiJFeimDLRkyBuD4WwVp
OeeXAqDuLJGg/3aq/qk1Kmn0pTttBUbfzNyIJFcPV96JNUwn6Stwl579kiY1
NWtKVU9VYwQU6yAMLWC7iZQr1xNhDpAQ2t/zppZQZRvS5O9WKfXFioortvG2
gxPGMU9ntf+aNHJIR38wcB0jEKFFF04CXroQyVFRNIMbYnn9+hYrfpE5Dh3e
xHa7N02l22fzqT6Wu0kDPiDLSfLoWU+xHsZwL29j3+gO0SKTOmGeANTctsS6
GBMCFxJEGhEKWbEODro2t65eGpWsqjqwZSmFGq8EnYGgm66HUbuUm+NAOm36
NHQ388J4LgNPcJMoINLc9sliz/5oMkYX75HzIJUSs3/UhcrHSZGyoUMgqREU
WBb9DWqubtOXDvX1QkNXx3oItjWaMnrouXDmBmr0Z5mfuNGb0ymJ9kD9X5tU
fLt4ye8lPof8EYXSXSstN38wbzWYffSCuVSfLYK8PU40nfVjGveIFdF81GBC
YBYhetFRVI5wzQkkdfZhNj/dFD3aUx2f6cuyBAtPZK+GCM0yhmqbbHkzmhrS
kTzZl9uO1of0ygDfrPa2pkjLoK+29/vuWW1dw0MNain9WYlsU+XjpfzVFgiA
Jv2jCBq1g9kUUhYgHHoQlXeX2Wp2gharSvjuFKQxkyowsmnso4zTBC+ZUZlp
tZYeJxM38ch3gMqHcFhLjmAdKQ7ZbL3fAMFsi52vt/z1gfxxSHTW8TW7jp0H
trRfKWX1IjtnEOhkOc+5WQJL5SYxmFrlLENrMbLmcvGWJWK6uY0OUcur+AkA
wLHLzC1w13rHOL+mFUSQrCt+XQ0JdypHRUDjAcJtL20KInxvhR66Web0+Bce
swKQdCpjtDaKdcoVVXn6pcDoRBLz/IeCsQrLzU7ZkWFiyKW5NVinG67Jq+w8
6o1Yz2i2FgvzFJ7paVmDDDCyay6kK4acPeXaemL5z4UfbtXrr91b5VNgBSqD
KyzWSSimyHpVDLuD4H2gKRp9jtOzFmHrwukO5/J+zYoIBOqkrdyQyfF9/lHA
fqI/ZTbg356rRzKL7F2kbhSc/m27Pgt5lnrYmEorjVoKCd+eFAQ/rF9LQbAN
vlZUbDXz8mLLaU7TUn9vJR6vA6iZIVOkmsiqkIhIofiNokn27InHyHk8VxCg
zO9YkR8C3sVUBGA6DrU/F2mqjjtrzfY8uyzFA+0Z/V0LgNu3zCyy5qELQy7G
ESGuHftbnBLZu8gaY46VAToHNd+VuSsy/HohA/3avwGIbf5YtcjxS10+dCV7
Qg8WIPwUX0VrU5rtm4RokRCXSqb6KzhKTDIy9Y0ErsROx2h8kykl8YRpsTY1
iErbqsS7Pqqbwh8o9btCwQl51RSkLYLvA1xWgi5ifJM68JmNTsNKGGalvl/g
6Oe0i5cKNdwfeA1Y6wF6StuY/AFeW1F5PcY3Odn7eRTF7y8rTcZF1oWUIDd3
ilkJphKiVNqRayJLHPo5G3gRl+R78G/RmeUQzlRmRdrkVghS9icljZslfScc
iLP5IyZd1D8iVr6htavKIz5gLeH0cykiqB8K3SdFDmly60/AaTnp0dOLIQJQ
sueHWzCEGG8OP98Mg4X5f93sZwEe+nv4I8+NGyk0nAoHmwPs17DCNjzMWoms
q1sNpypqRdUCK+5IiK28lRkqJDsMYJY+h5BQgHFz0E5Ps64YXGbwnwInGobp
avyes0ZqkEPRRq88Djedj0YU8z9StFnJIXYQtWuwcRm3W2BqCWnxwKApuwb2
g4le2NRl9OxMTdn15NnTxZuct6al5o/BBqo8WSEA8tkwAsmx69sIu2tlh/jn
l0wkMY63Zjc7b+Bigckqzg/bbdvjKxf7I5t80Msnv2988eaN3Z6yC/1ChHGI
q4iTe10yDjUYpnpfoovColw7cDmPD0+ShtzK+y0DDxqNPynpmgiSwJ427mPs
+CUsMKKuLuzDFBsaUCl+5l7X+yRdwef+3pGBQJtAcEKw4Twv+wzUac9mKObl
XiWE2jq6cgOV42qt0pWmgux/6BVi8pptJmCjs0dY8k0vQEJK4ymGLHtBwNQw
YvSOIMhF/th+cm9OsUWqGz1+MJIgGN5Q+1kEISGJWMfyHK8hHNd+COUzhb+A
M2ciE2D3nS1wSREgmh69gB53tSp0Ez+/mOuxs0xgj8zN0mBImnWci25qir8O
AEv9lYCeUqsdqIdGHHIQYfuPQlkQpenJA3tjUYWKMYULhwI0BP5STh8e6u6+
OAtMnOWjGW+sJYeICAuVMIofkFPVS7rxDBH0aG+9/+T4GISRTJ1XYio+zkh6
cSTBUWmUDLcz3DQRTvNIZj+LoCRHJJn/t0zWPWbIllAfG0rai/EKrCKJoBEN
aiwdz60ibAenV992prxmNA/Yron3cGJCSLrfdSGq/w9IShdhooDc8ndBw/J2
XlDvD3e3lP/2kkpwQC6bc2PP8RWiJ3ocUuiNAXPVPvRSdViGVdYYFB3hKrwr
Z1pqDF3JAQCJGsDAdTsK0N8wZU+yJBGxHZR9a/8c/fCIGEHVJQKlVbxOVRJV
M1eUz8Q/2KjMRe2iJqT6WBB2BcwAZjco74irDSNP5T3OtCdmyQTIxPvhZ5s4
E0egvlgVUOHe5yZuerBSPD6Wi1UIzQnn7Yh7jeIXiDXG/sWPwsp70spyzxN3
RPDDorRGhxiT1UEv7cAwx9ARmWExRr6doeo59eaSdfakqFJZtDB+mHpW79rX
KNr5nhCFCyeqYX4cAi/vBXSnFRXXA9BYWAoF0puhHwZrx/vQECmnmPAbW38b
d6RxXIePlnqmQvGB0lScebo4V0b40TdMM/c0p9ZbDAnr6xSm7I1HrvMRM6wR
1/odiowmQNo25HoElQkrQOFrmht6TgINfdCLp8HbelNIDYLo8VhyCgI5P0y2
FBXQQb9AHLfKTEFOijOcHL2mRpXaf7U8ad/1eiJPruQ6qhTD8CIxxPUwLfhy
8wyAburGVYH6j2vnN14ErlbQPZceRXeAGm+mKj8Bag9RxGPOBltAVBB5juO8
GPdGRT5fPFPvDcdW9SXi2P8P/aPZeBdmPghu15SxgAmnHkpR/e6fqGw7R1Oe
Lr1y6k0RPxfHC0c6SKLJDj/cB6p9EyIEL3afTnZcC+S+UokTQj6m8KukCMlg
uzRm/W8Pn9Pl9ZaZ173tfgZqjvnNzS5qENfKBzoBtWd18pqfyHT53lMiPvbp
vZza31ZArI1RS7qcfhAL9AEl8IEd9vN+UvYyqkrKjLLlIw5LNATEi+l8ZoUY
r6zmUy4ODm0QJNrDD6k6cIvCmwsMmozPpYydww2k7gCM/4XNwxaVGn9s42oE
p0xyh2CWyKQP06KzC5NMY0TNbtSdM02jC0H4cqX7DlzlEUJ5tdzhJKZ3qwy7
72RXrCMqW2CkRKewu6ucgOXKG1OQMbNnW2ncnBn2m8mL2f69RaXWW9uBwHei
944LkzTH8/OqYnOzjmjZmDowvxFFt60zC/HW++xT8c3Xk574v9JZ/OFAOVD3
P5kHiNEDs6pz2WbXwqM3Pc9roBPPruWf6fRoeX/hLnaIcigNw72Yi4ZvqOGn
smGjwB9stT9NFrr/2pljNX9d7GIB3Y/ct0kZbLWZcL533yVjCluHPDmyPM1X
BQ6u4yeNDWclIZAlE5PJQ7a86qfOfc737HqJwivpzuZr5+ARWlniSSCfHkAB
cIuExxrT3FPc51KarUCDV9++Un4bPO1symtjGeyw8IqaInRjbLdovCKA2gdH
Zt4rlBX7iAsNioh6J0OqONJNPqNGtYlpPwXnLOrjQAQdGdjBcrG/jL0SeEAu
+KVl86CG8wIR9wUsIPInvPgU+OCTNcFpOSfqVP/W65rGYMUIq2eSYR5yetfP
dStNJmKIzvGW554xy1jM0fmq6eXGSIB8F/PHbGcpUIn3qy033Ij73WKQBZq/
7EHwwzIso5r1pfC6ydE9qZV9Av+xlTICDVAvDdM7m6B7h0eesKLG4/LMbQ7g
Beleom7GRMdarsDhHFhFxjql6yJCFeqJ4cA14HSboXFfj291bh8vxxGTUFhl
KoT/YxvyxPe0x4O543WMZVO/UN4sXVZORaKY7y/CzH1QFvUOkTEPj+YQywon
5yy0/Om0RCcQ5AS1jOaufGhJnf3bBhnR+qKDzoS1gTT1nBAOwZ8YVbcJIwrg
estm2jqvD6vvDdDTx6M/cAUooQ1p1oRR/2zMevEDe1JMcwv4xUxkz1s6jpww
ciDhNiK3bRoMb0Hf6xZfz+oCd2mnQENy7mOQ/yBWn+YjsH85iwLUNdQPf9Jm
vl3MRl2qvn5aKQqzO5FiuasSy+87Tu/Ey17pZiBD5nBSK7UVvtTE3JUmBPOo
f17Ss91qJqJRDDIq4rWT+p490vgP4B8WNoDDPbP8ZBddDwzTk/p4CoLK9DC+
kB2VFk2cJ2G8uS4XqQjAfyE8c9N1MpX50qO8gRz3NNERPviasvDzbxzUBcqm
wNvO/5rvWW5oFrRZaV5aTk4E9D/X/IbGBX5aeBOeLuFav9KpVrH3ukviZhEv
LWP/ZY9wQ6fduhKVRvWc1lOBTi0uC+68vqfd+SPceb9Q9yXPyrlM721b+ffg
3PkE0kzDi9lPezHNE3pYv7bWw4sIEovbmio3aPvMvUPHGRAUTkgKG5cGDfzc
3d+dMjxtKoVC+4jK2V4FLRvBeUjg+DTMCOZITI2275E8LxKMEAt0v7nUxeG8
r4WWz+LLq1ov2yoChvmh4no1uSQzhlU30Vl3UJ5HdtztGDFdC+L0+tVchimp
PlC1r9WH2P3Sm6Rwyv5f839IBp7oS5Z6gJNOfLM6GAeVoCNC/vmQxSRVtmbX
Cq9kmtABn3fpS7dle/aNpWuXi0NLPzdTsFLFMBGa4dD6dG7L23KYa3ZRpI+w
Y5pZVg2RA0vzZcs5P9uoGb+z8PvJB2aYt1WC8O52hp7faGSFO9C7hHYbnr1u
qryesENxyDjQwobcqVtwgQLUtNDuviw5z2fKIPIp08Mr9TIT7XvL5MpnNBdt
PD3UqCO28MJearKzD5S0UVgUKeRtiqdCSjiDexcLNz1SgdLwh+w8GrX/P9Xn
GMI4xtBZ/6ZxGxqUBnZ65DLUQA8mqaWh1hEEHzlqT6Qq8YH8hZl34OuRZCa3
1KSirsdrEL6ag59NLYrH/iUBJ6uh/YV+NrlLErImFgEduVcOPoX1KTBUvcAg
6XAMV5Js/it7F3khVXkHdcFGkFHyKTrhEQ3FyA1gZRNl/t14urvCmMI+si6C
hZ7f6qW1pWUEWJQFRRLVJsKUPTh4ZAzKtrybuxh/ZKinDS9GfOu5ecXHysqA
gSWaahE4yDH6yC8WMcUcTavG3M5e7FM+LHpyLI3MaQjGzPnLdPzl/vlIraeb
xCzdNjTBRPUSIbUKuXVNK1d2NJaLOrL0kCeHzwkOE7MPnHq1mLeROI5jF6k1
DOCGx6Bllj6cyzumHiUnJlVe3tTAf42BOfsvFlGJnwfasRRLo+XnrXVFBRyT
amc4gQBNlbTR0G+f12b6bC+BumywkOC+wg98p1ln/UJDh9CnW5WlyYQWEVt3
iA3VS3tmlA6ScWo9LLbFsqT7DaM1OC+TcXkIbrfpROEs7Yx+/XkjzvNYML9o
RdB0C2gLvZTJfbkCdWTrYdA932L/D9lpKo1UGaLKv/2bXEYTvK65dt3N0cc3
o4PQg3rSVPjkAyuuTl8u6d0yu99aaIvVhQG/SP33UcEB16UBvMCROmVeKdon
Elw2LQbOVVS8P46C5VjmadIoLNIcvZVUNfFQFLwCrmC56zdhDxqzg5lxvO7t
PPorXKg7loyOy4s1GEHBDnia/kSKE1NdIJVwl544vGMxc8/lS649x5V9CcFe
TFoTRjv9bS/YzbQ1Z6DeHIzi3mk2JpZLK2PjT6sGwDkte12abMPasEMX5Yqu
Nt1GUzx/Z66KWxma3bwF93Ayp2s22/OlkCY5n0fEGvtNAFf+Brlp0Ao6DW9P
4XhoM52tHKB3vXNHP4i95Cc6iZC6reHwtrof+7iDTH5vwYwubQeQSnA2VEGT
yHIIq3oCHF87HLnVpwbL3pR3kESRyMF+Iiy70sQ7oSaoPiyS2tQuIVB/iknl
mO1ax/sDWNNkYvlID4k6re+lzzlL5L2hhyxnc6Gr4kmJPBeShJnAfhPt/xbX
usbzPOVycaA+5tADHdJLoD5TTjYFJM6zkM8Ygsf7EdKwyonToNCXtysTf2Qk
kJ3v05Gl0aIrrEB3vnjEU7PsyfmB5uxsG7NH6qKzLViyH5OADxMBDhYUYWMP
NTUxKZURK0h9WXXNxWZhCTq9tD86SyTw+6T0GJhX3qVaq57FLe5C67rIjLYt
a5rJhnVqhrHqNypmfT34ljQJbm2phQm2MNrhjUhz50e/8q9ERs+lhfPsyBoK
h9tjGo+Dpc1e13D4gpusT3bx9M2Hdo8aMfN7JnVzzmGSAxTp6PRwDeaH4H2y
di89YpQjNxXUZmYg/Y8F0bmkesa1OYb1OQhqsWCVcnpmIn9EGl76sRZ50gyl
sETntu5hT8RnADwAnLdwU3tluZDolZXhufpJ7OvYWgsfckz9ut26zijmpZ7B
uCQI5Payge64Qst8lyBqBvz50psX5m6Mwmw2YhMxJC8mDogndAJ8c0RRtHct
w6DBJHMG3XU++fWvr7JRDykSw98IumC/GfRYWD6pRnUW0ldSdWCZ60kM4IJY
khokoA0XrpvGOB7f/ZUJCU82ZWBHicq3X3/fcl96c5S6x14YdB9sH1QniEsI
MMmPDA8GC+l2BD3rfAs3yIgkjw6yJQvQMDtzOexYw//sooQdwgzvA8XyNz9M
MzpFgd3j49jauCsarOVC7V3j3o9dgUzEGg4sUu7Yq+GdSQxYc0LgzT25VM9G
OnfG8ZKHkBAoUycgma2e6cZuy8MGtu+CeEbg7VFn3kZT/OpwfdlDlO+4GqLL
6e76/hkmM7Oik7FBklXJcrjxF8J6NgXPN1AacKBxgvN1TbBmU23dUSPLWTfz
LMlIkE7g0+ZnG1FaCQmai6T9srKckQbl+CtFrvS2kZlUlpMVNA6IiB3YWTV/
uNgsBtIt5d40O0MRfSAwfWb+M/KxEd8kLNsYBPCm6BFaTv8WjtCdzPOV7VCa
jaFH5Ejkv3hdFEvDRfBA95a3uWQd3QCsLSaqfsLZVGe6Fcj4HFV+w0K8P4IW
7UlCVg+b3twDM0gN3iu2c8eEUzb4lO1A7Dmg/qDpCBhmu2QXImq2zx8ykb03
co9lNqiFcKSTUyyS6s3OawNuRDo44UfYMNnzsJExRiecio+lLUUf9I2eOigD
jtC4qyIILR3ZCfmWIvTluHHr1ggmzfg3W/T16apPRFA4fVMJgphliWmUFtmr
NrEJrg2Ojse6MaehDgRmaSPjK5vv99pRPqFuhDRWx/bIiwRWeYhKhSPKNMZz
13qsuZi0iVnbpZiiFDYu+b+vNnxTlGbjo+bFYiF/KJll/pti/JaFiRyo+h4L
Paxqy7lrHzBG2f2L4uuP/Du7OZWhrVz/oRlUPB5jIMmdqnQ8DR/jTyjivOKb
/x3zzrP+n9zSP9Wbaswx097Gcmp/MGjRbgx7w0d3xzbkLxW6F/W60St7tN3A
38p7fctDExDIODV/VXh8Fy0dQVZmA2IglNaWr2PVRVBPJffWLanIRrvBhTTr
kvkOoNrNGeuo3AukVK+YPS6WeCzwI2t9k/ZCCnDrJXbIMe7gtxVE/finZauD
Q+sUIJ8VSya9scdXYQ7IrA6UaByrM4D9mEn89Az2ZfyWjqkMyCKuHj3rx8mT
KPYUw6DFZUye9AvjcOsH8uoxh7pkO9QrKp/CZKuCMoFAohOZxDw9ryH+V1KY
J9Jc8mQiXRfRxafKQr3psrk7IIS0lWoeJsteEJlxAL1fid4JnctJkJXGNknP
GTMpKQegZwdHVcVVU1xpbl+rg3jBbnfVoBVjxzWhc+ymyC11XmptcZMtF6K9
KU8E9iN4Hx3nBsXOyXAFbOkwfDA+H2AVcEWqz0GDE9BF9xWfLkSqaQtjwWkH
be5qPK6tPBLlUvgQWR0Ft0Ymaf97N0bxy5XL2rtPh0r+kVOetjddNpSKDDI/
J1F2sR2Gxt51ftSSSIxmQF3yqIKILIOzxTbQZOYP4bveY8oyLeegy2eP0JHB
MrHxzyfhYj45RdHgLvjvz+fxh1kFSUrUGIwCLqO6Ii2BsR0KFQ0xFR8xxdzA
mtvaACmxolllN9DPXnTaQne97ZBSVXtaBGx2GRTqZR/RsDbEKqCdFMBuBwwm
tTgSkecaoeAxlA4uxoXkzSO4th4ZkOf+TuHTJqGYuYXMqAzgu1Ld4mBtJ04/
Fr1DgRQMfSVNs20hcF1m5YZXF5edKRUblIhf6EsrJ90CPBt8L6AU4Y9uzNFZ
7JXFzNgg6jb0xWiza7immQZ7YWBDzUTafeetVVLySzaKZmRn/j48zJL0RTIy
/7Rfkt3Fgw0TR8FdQEVQfHkJ94kUAbGJyB3/xJOI6pO2msCii8ELn3mZ+9Iy
hNW4sjTiE22q8qskqtpwmcT5jXcAJdP1vPcP9a1+zQojOtI+csCbL1v9w8Kj
BD828cLfrZavGbvYKQFcCompJD/5XLnVcrl0pfnEFsH0xaT34r2cM9TnoKUi
7OQs9O1WMJvIqegA5M4r9t05q/meBe7MFNj+7D/hnL2Wl+nDe9NPGuxwtTtp
slLSdPUXfgBoZZDQc3fgqOzGx0v/SGsr3NhJ9rTS8yQ852z63C7eWnLimAlA
IAbLeIy+6CW6mom5hEpsZDHqmRyDt984TQ7A/XMwsKLufKJvSUPzpP6c4cQg
pGNo7qAA+e46pSLKpMW/e70/DsgtY2AQ6bdhuGIcQbgoVeNuH5Ys/axNc2A6
4onWYy1UNDc/8gTGYfHFH0e8AtXRR+b4Xp7aBlA6aAhqnqU0UbNBo9GkSDml
xaNHltcUoM6WqVQiICa5TzjsXRwjmeJ/hDy8If+F1o7q2ELeeJX99N3Jw7XI
qmsCDBFSEwXF0nn4q7i0joYHT8XMGYs9hTA0JQdXl2H5i0K/5Rxs7fMELBqM
P+g1wOSYU44YF8tIZscTGvwXNF708uyFN+uSjl9sRuB9c4z7rSQ+B3mYCXl1
wrakwAYx1JWLg1uHVAFMA0fQeD1sv5kMr0AYMOB8GnDtjG37md2WjKdokLKU
XtL7umUvANzG7wX6cJk+K2PiiiIKCbqDjAoSJ1s9uD4Qjyp/3LhlTxqBvr0q
lmwrXf9Pve3Q8Ht67O8vWZUslGj6kpR/bAFY7kOabL6l/kCqotVbBxZ6NmVM
hGAqvua3mN6giU+LSZwuAou5LA1ObBFm7Kxiu+P1UYyh6oHYTkyjoIncPhyb
oTN6iBQ8ERrTSQZmrJ/mS1/LwmvpHRsiURb7aosovZjQ5KV3sxMUkHgTaqh+
zILJ4LTvaV60OeFkZTUTr8d7npw4S2GAsuhkC63GvNcw9nT4m5td2djO4IOa
Oa3pyeHqCeNQtYYoVUwTWcXNykSvRhioI1xruvZcVlrknhLbJcgmAXTN/enJ
4wB0Nce6zJpm+Q4XGnMyzJckeNrOvxBwPNT6OMl9YS4rAroHtuhhm/CRnXwX
pujBykc+hAg04d6kwoxStgr8kueF1RliJiFg5IgZ9JTHd3czlZE4T8ooh69E
5Io0FmILS7JzmIt51ecfpmtbWZp2aca9duqQfKzqzS9ojT+nLIQeRoEe5hPj
lnCTdYrnPefgf4KjlKFMb9PFUVbaCMeCddghk3AbQzd8XJ6sfkajY2dsTF4F
bM2XUnXHHwO3EN4wQjkFI1Ex0pdN7RPLiDR6uTFsa/Euy+WPTxlFAB9IE6Pb
FG2N0iNUBgFmSCSq/zHIG1uSJ/HCLE6dntmi+RHepx85t3Hu7iGz8uMGrY+/
a52Y7IgrjrF1Kh2immDDISIp0YHZQvv1/ptn69TaZZi8/ewQJkNO35p2OqL6
O5KFqBjGKnKIcZOL8N1PiORdEh0EiajKvcYQFEVZ454/jmVF8k9th4KLAX22
g9qjp9eolAIO2Vb/oLIg9q6UaotdxbeYf9Q0PAC+yzA6J2Syn1wfvo3saT1f
t4lTQoyYO+WxmnT4685kzpfffXzeHZ93AVomqxVnIDZuIxQj3LJ/Nct1r7pu
ciNi+NtWpKlMTPcfR01QLj6nQd+BeXjbUSgHICem5GfTmI3vTqVUa2eJN5Ar
CbDhdqHOfpXSNIwIOd2yof3RUNCXYvjbm89GIho2fCkTATcJbBhJ2qBJ1Atg
HJOH4J/t6OtAbR8kOxMszpUV30V+AP1k7Lky58qfcs3oHoTE2s5HTQG7e73R
ElenWGZZ/3kzU7L2THtj7o2hd3nVLGRi7zpJl76yVX3/cF6cX3uRpgq19+Uu
DYveAEpF67sVtyobG3YV9p3pkXgmz/5uHyb6QedaXaescjz+rCZV/4VM9Ngo
mb82zLqq0MQ2Zqra+UH6xWuX06SicFMONrWAzkmQdgMqr3JuK0yl/o3qvHuA
YkGqC4CJba4YeGLZvyAIm4Mh+WpT3Tg/AfcQntQ0J5cQJBjjdMD7N+Xs2ZyG
13plrZqbj/357kgKIyXZKruY6H5k00oL4sxHHEWl22L05JLw3ygRCrZAIhXL
SnoU9rBlogmMvfTNgWX7U5Mir8LH3qQPgiNVy7Z1q8PD/DuQ0rVp432hvJuf
dk+uVX96MySaNeN2ODbZXn+L02ZlKupfLNUUh3zYaq+lcrQQPXgb+LJY2bSM
CZRbc0q3r5XSt2rX5zTdhtUkuv3070EHk6S9KcbiMz0ywXq3/QMrqka6nq9P
NzpFWFSM8gYwK4Fw00zNL2XgoQ7qY9iTDj/rCpzucPunCdVh9Qhvvxlx+thf
AbK5dHReYVdRmvy8XaESYhi8reC05rFYYCh6il7YTLtZl9DtKRDjYtteSTG1
ZY02biJ+OgzKksNF9Lm5diK7YB91GxV0IIN0jnM9dV+jLcyAEHm9LSSba+gq
ThI6JJ0lA1wRnyD9Zi6tt62imGGjqsxUHL96ZnnMKYl2KjnmpnHvjZm94MkD
iDWBNQZY14t96DAsnWRseaMx92sbrb296yGGWdaRYvSOYLAVlH/KRsnF9Rn1
SmqhdT5r2acIkhrbnKeo3GdeQGr3xsP2WhQVf+KEoa2/9uuG1zvZ/mpZtoru
BtdH7udB/54jxr0iMktGKsQvuEN8HflD+7x6Uq4cV59hLsyRGspVcv2PuGSB
xevUwbce3LYzEbQdnA32C0Yy3+nPUu/AD8DXmN+ftSMoger7uPd2SEt8z/Mc
CsDksj0ul8OcQwio7lbNcNi3NaRwyWCZeW1KZXYgo1+Eo1kcEUWtbvfUYX0c
vurBVNkYipSUDfsiCGnZFtDc6DJfDsjc3NyivNR4WW9j34sKHcPyaWal2yuI
aU+pOgXwN+iJqvlxM3RUQ5tu6jZdaA6T97TuRnDJQtUJw5PDSYDM8L/JswtX
FZirjeE8hd8S0KZdKy0iLpy1WDrJFebuZCcYdfBW1+Hmgn1raUBV8bllKprQ
7t1JUcHt0cDjSnQIE3tmd6pZPeEZ6JDIGE0QBEDLyCwB+iQ/aL9pnDGD4g3C
31PzIBOKdQ0jcKnmBJFhILdjpR76pFNad/NlCc8b8R/0UlYKr249jAfeWNIh
d0sAe2K4oolIjaWkzAWY4EiPE6GegQOgaDKHHywOHqjqHiUQkwGR9MCMXRgw
Y+8faiiEp7O2jRrQw8ZCJNqxwwJhHGNwACy/utuhQBxTPMRpRitnMH5bj8km
JSB3yMKt0z76KcJDiITbIzA0XiVjjrszZczrtfEoPTh+Z2Wi92k/XTfWnOug
+/lP8bIPGPkRxszD+Fi8Aifdsi3B/b7lsyE3Nxp4QEdWGHYJggfFnHFM3zPR
hAwJgaCdNHmsLriLLErA129zP4I28Fk39b5m/rnkfpmrWeDsxjUqh+vToLpW
qrBahzW3To2XtC5GMoLReiNvaV5Gfiic9mcpxOIQTtt6qvENmOGfZz8CWt7H
vJBzQ7+1FoZ9rSr0aFcYpThIg/rZigTRx/gFl/Xl8JNOfjqiPf7GnXh9m//H
ABa0NAKo1vep/K8wQ5xn09aLOItOwo+ILym6AJLrEm+5cf2yxar53bSRHjGw
SvvyRrWsD3UhSy4zz06SgfLwpRRrpZ3NA5RenApn6Vcpen1S68RsjcMIZd8t
xNZwRXXHb5DBAoieyIMk9MSYYU3/DEhK14i6YNUeKTnFSUXZ721DdI2xNZtl
tHGMT/kif/nvAKOxkch9tZpnST9MBK+TXMQbJEzf6E+ut7RhGBa/TbRahdQt
cxCXhDIdA4qCpI74P9eI+LtmucBp3mHc8uv0QUH7LXb3xiNRGxWSo6Sxqsbc
s+5NbavAgJwFszJEHM/bSe0Fce70trOmIECms/Dvi0G9k3NZ3Usi+Hmxws2W
/T8VHZ9qwLZNQ2V4RgdQo5gzkx1TUouwlx2uBXiql5o8zdgH3WoiVfi3AB8A
PAFfSf9IGWT3WDPLrMxUfCdCnKDQBAi6NNDBhL4RvXKuVV+DVNXj2Xgun+NA
siaj6dxHbsKogLK0HQZA4Xoe3hSfCDRxoLAF8bO5y9KiJ5BDra5IXeJ38Kcm
WmDQLWyHpujbYIFWOqOY1DLBtC2++lqBFFapEOZOFQ4WyvgyouaPXQUQg0K+
9Dff66aosaQDwwnEFvDTvcFe7cHXNixsWaCgE3b4iZ9eEA/14sxrW8fPZjSx
gxuPXu+0q01cYp/cj5RU1zDddc41tYRdFCFGAHxOsCROoVkQqbjgzl2AVLFf
L7OKC/r4+42IfEgi5ct/zQzae+d80xoNf3HkP/B+ozMEKBKPHEGiOZ3r54tK
UQa2n9dSMbt3N0NBc928wpBzMnsXKnH9EB81pgC6Yr4FKl/EiEdw9G8PX4PL
xWZCkZBno17t4Bsr8WbLAtGiWK6AHmbqGuqzW3U6Pyu3/XzksaKHw1y53+tc
ekj3yKGByLyz9udj0FsNMzjuo+EfXdCwZOdkYpbvSYD09t2Wnz5j8xARNS+i
REycP9MARFTD70Ow5uZo3gqHwfYgAoF0NAIwfPZCIBz5Qrzdwfe05t79DwDK
vbUcdSafvSmJ2AA81ev0r2Q5QnghgnVJx4DRNBM2uaghGZLjEXBv6ZVjFG1S
zz4H/C0C2Rz05f7+LFHblvp9wQYkg6q2FolJ2fP5SALQdHMnrnRq3ZUeajtP
7aZ5X3LOtCNnoJjTP6ms468oOpjScFuhfqsdoBDGOEHYVSAbzfAXXA5ukZw7
oX2Xxdt1WaKUU+oBK9h+7olk3xlyVH9DHW2sW3oGtyhClr7sPnCoUKbZX15Z
rUcvN/A05HQNtD0ZbvAkIkiriZKnAW7JXPAY9crxN/9teeOEzd6V2Bc1gAwa
jRga72xK7FqDdlZQX42K47hl3DNBbvk8a82z4SkjpJjwjOPVyzGtWk3gEbOB
Aix+iBl7z1Cw1Um4pRzpKI2/edK3U54nCb8zSMvbyOMM6NHeZMY2+j25olyk
nOjPl63/qUX1cpy34ZL2ZJP1VwcgCwApwztwuk0qQ1+qwrI4EyVkEE9bLKKI
O7/qIItjACzhYtPogoGbfyDhcrfucLkTSunfMO3j7MsrWjdtGvtnvANZKRkG
+tmo+DfZNQF+LgCPiHtGDVxmuXrL4FWOVXWFzLeX57WIAmDVdYeOMzaWKEmF
RKOcIAispuueoRAjFskFbNXI/+zbJzdYKjnl5iJOB1eRAmGySlgl4qOnV9K/
9OGIHFkeAWLvpmE7iRI0efLGsSJELIY2M7SVkkzKqaTBejnCMseOmktBZXSa
y6hBUKacIMUZZizj48JMTGWPQ5zLRog6qqQBcZ2N3AFUYYCTGj9EAOd2DBXL
jB3wI+HW7c78+hdy/ifX8vW50eOBp+SbWGIpY3be6pN7IYG2S5sWFtbHj3Lv
f2DQG33jpRu6tZdpKdSnKfARiynjPLLqMhM5rP3TeOSwXVjeiTFCTMvw57FJ
+F/Z3T7IOQfYFwZ0JA1J1Hz8k4y8VUP1nrWTHVusQusDsR8VFhHMhKmHpRsq
dcGuPnewxEy18wy/qLSjm9r1wY2x0/9IcYg9WDlzmY8GPflXuikkAgxYMxXX
+AAwvBgbqhy7OJjHNnsCwr8EMz/aZmhFq57P6ehlPgnVET/d7vyfzb8sr5Bg
h8CLJRMnfRhizBRjMB0A04Z5xuQFkX+NTJjhRByYbePK8KQbqf0OQQ3fPfUs
eIpEZiq72jj40Qr/vFi+qEyIGRll+SGOsG4acPK1SI/lrt1/SnPxCiV5JPu1
NNw1HVTwBcTs35uEjwGtZDCaD26Yqlc5v1qdwdQzmdE6NM4hQDt6pww4ihVY
85cYiG/LAZr+q4Wdu2QxrG89ZydUPc+Z6G8Rg/BwhPKDQItmE5Inw1DKvuyV
CDWlFcyrPLz35s8VQikl0wT3ZKoptkpzmiIGynXVWwVJe8YtsDS+456eXoRC
BugbU3qYmTMc9pX6W+Aog46fLexTl6hkne5DsQkSbevYCAU55dmynIdiyxOk
y3FV2U+2tD1IGO9fWAFPvCv/sSUetxielgnlhwtFIHikgLdJL8ap7QU+vUW3
0ZOk2eaSXLG1JhJYJCt5JMztRrAz4100zdSmQ/gi7NqL/Vbtk2200qYNvhGm
u+WIwwKtB+F8FLYdKG4V24sgHJFHSGbpGrbvd+7U4rhda0G8+PRpIN38JY3N
JCSYaa3I9mDlfJCsR/98CXw4um5+OZmp+7AWUOWWrKUV5dkCDXDuZgJ3uat1
pfDFvAdYx5LsAb1c4HOwTavxhhaoHDqX07I0B69t/y4dNDZ6rm4NuYC97n5n
LR18scExEQkviTWFKNJ6ihHJf0pPt3P8PibQ3Awa8o4BAUxPDXw9CXvKGS4e
qP+Qoy2Wpo0LtSA/AGQe9mma0ljnq/fdYpgXJz8fP13q+jsn546GvxzyKwXv
OLhbuQcnNYIG4fcvXswUIZ+oFYUCRk+RrtzWBsqTtkzwWqR6zDdhDNiPcn5A
odFBjwulQl/AYF9nz+aE49OC5KuDPRSK3REWCFVKELUBhh0R2bRyUP+SJa8i
YBr9ouz/NTDa/ivBAamo7Dfjya1Wjvc4gz6Nj3nXD5LDjAXd6Ak0Ro2KMpTq
1PYg8n+6vAQp1wEmxQkiiAWZDqO4H9wzmMBgmdiyMsnihudX9NniR5MM7Y3T
R9JqV12c3NbBKztCAuRtzZR5GRHiG4i8aJ0WcNJaatcS4cJ/XZJJrg1qE2RA
1MIYHA3l88VDbfi7GqaYvoXVcapNGHKzxNz4U4utxRf+xhl75VAPl/yDzBai
EVm44Dz7fMBNd2ZUURjR2qpac3AQtIssMn5T5Hv5TN9gfNleBX79XGp4vGYB
OVwJzZTFndKcKiVxIfQ5iJJ9AtlOzy2AtPJbUKWIfbI5j0S83ZRRnDHFKjRG
ugxuIeJEJDuFbbs3uOmlobTSyLrn5KdS9mFCVH5CM/9GANfLug3eETN2AnYH
VcmKVXNWAYCKqaSiC0TEcRlmVeacYnWyvwHSV44HnswNGsFcaY6N6qLiNDyC
QtUwFqS0RFgqiyxjXV9ZyG+t6YsA3r6Lu8QVBxgGkfvzIyMKDfkEJtwOJyE9
BAkKBChCMK1yKu3w+U417RC/K8zh+Vbh8Uf3yD4TaKvklqycvHrhxUWzw/bx
7ypMvJLXA9JDMTHY4hqbtZJY73PzoyN0dMVeNpitYGNCxfvDVaiFKO6NFpeV
UF6hBRAfbYUfFyHBkVDnQ4f48hSjIDauamNslelKO2GrhvF/5xwCsrmLDTVh
IT2JSVpt07KYXSneoqIRFRKcBZ9x4LZUJNgdbJeuRZO1eQsxUYsTrQv7V5eh
37B4y+ABxFgeX2hRQmWa6Jop5TM5nEiRygUNLjQIgDsmWGjOAQyHRzt79n/U
zD7XhKWuNxeBYXx7YBXzKXqtmeEc8SnQjcNuzB0+uLUptN/ClHqItgBZIwnB
0WGqfUHcmioYsOXpOnv8kkuMsC4qqonGVLfGuP5Z3bBOQapcDl5XhOa/xi/6
AHy06mv+t9cHiwAFi1owEqTEJpJCvFKcsj0MLtW+HQ+YjPUffKwtuXY8OhhR
ahxxMUThkCUluqOLxt0Xmxq0peiHl1BA4MKdm+vISX+2b7lAZ+hEcYdD4gPY
sAzINfW6mdC1DzWJ6bqj347ztWmu/GwDDsBoEprsDIfw5RtMsWzZnr1QFqE4
66aYOYLTyyElijvOrH5mAAb1T4tOu7QQ58nBpcsiP3iY2Tic0xavUVuu7x+V
tcTcFwvScKoXjOBQcgQxANFX6H+zaYE69B3N43ic/L3IcpfHDnrhFkGogMis
SJgDohg3xt2qoonh0nwYFJ5dklCcawDUqNMS0tYR140pbWoF9/QeQwXqpePb
O3LgvS3ySrRXN48TUpxeCNxgXgr/YKISAns44vDYVbfLRzX5Fu60sOwyDUxS
r3PDHf/QXKe0Mk3A3P1zfWj1YoIgWrnu+plKqsjrMsZYcAH6g24tqAVbGdCS
GeUWizxL0EI3V0Pwp2mlSUg2xHSISXpmbZ2VI/OWfruzcXOdviK7zKDu8QF+
wIe8wjtb6Di775StNS83+X5LIYvqP9+T5cC5/PqRV5a686cPT0++eh5a12vR
I5J0vdo7xuagnD1PQdx1vWfnQTsKjBhas1gjH6A+c5SEVO+HBelIwa2fCchD
zD/fnAU1OviHpJK+apcgjbPfG8JRzP7gq0NBjxlIOsMoRCfpYQTl5zVI4eep
J8uoRSJNifkASBR2nIsi9BZEAdo05aEgc7eAGRrxEsf6Urb+pGDQNp+6eGI5
/0osGmhITCJulC5xcYBPVMDjlZOaQLTJ3uCo2J/JbfW/lTDealcRy+Q6dreU
Q7rFai+fAd7aHJoOA5whCon5O8QqZ9IQhcdQMSaXaMg+X/p/CV9VI6JUKVjS
b+JzNrv8bON7fSaJ6MKMSeIiYEV+cPUAFbRCulK0gk1uxbbQFnS1Ik9ubFCc
4BknwHr1ov88YhFHknTchVrSz0/T0UhCCZTWNdEranDBILF+TmyTcU42Weq/
m+MkXN41Xawmaml4IVLqLmdXC3pJMsxQngfPkAjpNCFeVq9WCih7OONt3SPr
RqBWsSuhqniRkY7Cs6HjGYpu77pRf/uutE2wbxaY0ZvcY9oLGi4vT90/pjOX
OFJyUT4wq4DcyqMMhf7+FMQ8+YkdiH+VpOA0m+2TZpe5aaIr9CAqPXtCmtnc
I6Jc5MkHUPB4yTqU2rvA31W9NlTq7xkJ/HURC4QJL/iVsG1xzV6mt52AYs4N
xloBEBiEkrUB+i2n6xWZ3cfRaRlJ/hPRRHcUpHV7M8GD76mHC/m9L1QVspXP
GdIHDw524d8lj+abXQJLDdHrTT7X7BhyINI3FnYFc9bVW8GPqPkDTM2iFdXr
XJN9VNijTd2g/jRiJ+74w2ETfvHJuz7l/mg55NvMT4OLOOCL1Vk2ERAcvtn7
xdjQjvcNtmFE7I4E3zl1umFjC5vSVIiFhbi3idTaUYqhYfxNfyFkbqZeUn1s
U8r4UUe3CGMN81er37zfD7V39iKB0m6ufmnj0NG7kjU/Ml37MvEciJ/ZMsJ/
T50fG3FgmuoMGCW9rHC6TRmJvpftEpZbTjJpB23PtPLUmRgkD20hExsDq8RS
TMr38OxIW/spcQjSn/fr/UD0ujsIRHoRdEBntUVFa8T+RXfwjn2PAXI/3ii2
/AF0Mt1SARTQGInQrZA6fSdxZ6VkxxqXJjv9fS4zNqK86Ep7jKcpogn4Clp8
din1hmKIjv8br9fmWATODE5DMv/1nSaxjA0acDrVbLRxq7QF4Wlqmx+J36nY
ch/tlC/nBbRkWdtDEg1WqFJ+2W7Mdg+OuSYTXxMRcO4J0qN97CgZHNPPdlZJ
tNYeSnh/ICwXQ9UiKlrLQ/3OrftoFLcb2Zf/YsMtR7IV3QVaOjvJMLHeAEin
wYqhbYlFO5aFMYzUNJuKe1eRmc4k6nVEbNJNzIQsLlwR1Iwux2qZljU+/XkQ
HEEBJp7fZVopr3edjladCjEWQF7woAS41vsswHmoYYMyTx2RoY7dJJQGHo/x
Sg3Ys6x9vfBWZKFNTgP2uDKSxksozXKohRUuijCu61dSPVZv20+lLnTQlsbt
G1F9pa6cVT2UKYLWcvLzLsbgOvVpQcFB9yHebqSIzkE3yohWVFlO+Y6ntXx8
JuJE3OKHP3YbgtPNJqzf1DQ2CQS4TJvH08IH0PcFtg+mWMr9PR9LrXwczHzL
l2i1M6EowZ00msUvGIYX9r5iPU31n0H91SsQ+Gi3LA2QiobUnqvCzH6gftSm
CYVkNxcXmzRZuQYE7qJNWr0hdUgQdgVraOvfMVQt6qB4+Du+L+BXm2AGe05I
A/1yby7DhWRelM6IFc5BcYqmbKQcS2KLtEZq4/WgiWeyd4ThNkJCvKL7tBBp
rrDC6LQvrBs0NOwbhRrLpbAZiQvowvpnJX5yaUd5rdr05PIlcD/GGe2MHZ4D
WnKQO5xs+C+/UExhVBnzE0A1GUI2FvegEzy/JxVjnUNAnmFa6YOPSlKGtcLu
FfI3fWkCtZlWIdAwmDxG8I7WxpmF0yyKTrqE+9J9LeC0oUqh2lfecwDyNc6i
/0ByOwkDoHVPz+nYCgYLPDrzUMbuqn90O3qytoD9IeTMbVgbBY+miBPYxsNg
UhAg/yw8/sEF0pBqFBxp3TXxDICPpqgJkkdGQDBPFm+xYagvp4Y8dwvmGZjv
UZiMjh77zRF/akJZEfKVEP/+J4cCm/2QEGEdZarI7AjBQE6HuvQH+0jWhaaN
43TuGEZZ7xdjdc5IguREqsgG0eHvHj4MbZNc80HY1pqg5ball+FSeoA0gyFP
XaHhM8VtI0/5qa+4g/oIASprd8UFs7uJwz6pIU7zmZ0kUKAvKdn6AQu8p7uo
EDzSP3DVpBSdlQ+c5AeqS3hheryIVU6XOAM6MK0AAoJwJYlfhwXe2Ekfel4P
Dw9ElnH+p53r1yD7C0O/lBSG5eJIHlSXnl+yayK2g5qO8yzuoDMnE8/RXexr
843C1/HA1ue1FcqsXZ5ejOZD8zPXzaFgdEjATCD26hiWSTCH+h8YRNDJCw3x
BUAjN9xvDy34jLTi1yVmMvMGI0+ryRt+EsZHPTdovzK7K06duFIw+aT5yYec
370bXzvd5YeTMDZ6Hz1DaMWuMJ9BzTMruyFj7w+6lLB8DhMDvdgFQ7QfrmXX
6H0OAJOX3HWu3QyhQSUEHVT7Po0sryftKvqtTJGkbh+6B95VZcKKf8QyHGeA
tbAZA3kyiKh95GWtlfA6uuwp2zj1k2SiRhWkY0miVbLZLbGyGGZvx/WaCiqW
T3REzz3bJBBT3hp/tjnpETiMFV7LcOJbOrq9Halvb+3YTF1x534B99drPvi6
GCIhToUuPbp75XZ/HvxCF91JV6pclpyo4/A0hHGGe/hUSt1pueXPsMsXo4RR
QQtL1JeGUv9/gAnTTyxTkO29zLPDeX+4QthZ7bpOIYu2eMUtK/y/Vjwctsin
Bx91M/Ij9w2xZsq5ku9+SZa4ZVBLBDCIEp8JosiWhR22Gue0pQ9l23h5FPWH
kTxSj0vwPcWPY+bmcG0AryjCX1boOGNW/3DZtTZzNzHFPrTI0SicTP3yU0op
yIA7F1JbpcpnikULOjhRPR4fpbL6MaoHDxRbZDCc5WZ/45/2EA/VYEtiNcwW
hO3IS5tlOfs1KILW1mdTQRybr5M8GBfQSZNYlDt4QnyKUN6APQVfT0tqUoCp
r7nO95/FVEUHpeueaAIAj4OFuEqq6ISWReTYJ8c50KjkkMBMjd18u40aVMBM
VhmO128MaLP96gJXqh8G+DMM+9qc45zc+wRmv2dq5u8kR8k83cygRrVMK3ld
VVV4WXVDIL9EDlsVTxtbCmaz/eTvoyCBlNkCktGC8r1t9x9DSpAD2WmyW4Bo
cYATD5heExLGXJR3HqS2D/+m3oQNgNZJDJYFc1sXmS7dXg3kVxTcNhBLrrYm
HgM0mV1pjjJmfqMwyd1lPC7A8V9Ab8U3vFJjwWAyskRT8pATKazwPMFzFue4
c99gjVgp2e5bqxqo975JDVcqafRXm4sknUBkXvKXf1Ai3xQfA6P3P6F6hWtK
rgSIgkSiq0lZUYOIHGcCQnI7B0SSL+YL1DSgHnQ5pyjVxP2ulilRp2sM5Up3
2cyIpfb38wCtE3IGDzH7OLXOlMDxbJzCNEoccVPW7bEuLcGgjDoY4+/pgZ02
lFUpbHfrzBmS1A7FN5XPDGCXldCk/DSnYbGx1lNHM/qGZvvUKkCzZ8CYCGte
BVDFAXKbBJ5k+Av8ixDC7vXDoVwMAU5kzVVzkqlxhEZuuD0PtTawMS6TvD2u
x7LSetZ7SDhByFf7ur2uD1zMdV4Tsf4tDwPWVMWJy2OkdqOBqaPLRCylYvU+
M1uBqOKQvRGZdIeXb9TWFmTW1ZZfM+bcdhHoETaM1P5d9jvMA+Xp7vA3lmOF
iyD9/hltjKS38tyw+L7P8M1Q7fef+WNcfaSDoHUgzdlnlqbj+eIfdkvyd/TX
YtkHIDrUsTFQiRSPEvx/TbXwwvVAMbWjijB0r9oyjk2jMQxupWW4myZdI5Y5
KZ8BiMXinQrH5jnVybkuJ+uSuOHoJYubkSdrWTege1iO1wGV6IFOFXkUEi2h
SQIFcsVKGtg+OiJl9qG6JWD0CBmi+uLHNoSP/sj7FkiyDSo1V1e4gxeO9jGp
+3Mdp+XOLrN6pkFG2R2b1GLpE8+Gkfs3tIaoV1ZkojWMh1goO7lb9s41iBBE
4kfs6tal8nZUjLMTltaq+hMX2i4nSN8U4ap80A7M3CPi0eeXdtqRCt3DeOrn
pHtfnTkPRb9io2Sga0mqIb0xQqwo9rAfgrY+J4zT9tzYV7pIoYpE6rHybWTL
IPavZYberXFMBroST5pFu9Bv79T6De2yIBv5xyFvIlhdfm+L9AiVbFkiTe8w
v8uwH/3aOLkV5P8fD5zS28DNdzp0HGc9ahQzTrxKDd52GWzeTVG0+XoodRyc
fbqpHCDZde8OdB4qODxEbR+Gjca1jiVwtRv02pFpqEzsZXiqMQ6xedYubx6L
0LnN+z7ueN9cL5G983/ZroKMzK7eJOdNAowPG7MoTuoc1LcAKg5JmlruVL2J
0lwGK89dGh6d0JMthectbJ0pUSP+P5SYe3yPnKcivMVUHGYTj24qb2Tl1cEl
jSDnVE3KXXbDidIaTRMAEz3503k2XTI/L4PwOXFs6yS4cWHC2min7gZ/Ja0r
MQvcCMs=

`pragma protect end_protected
