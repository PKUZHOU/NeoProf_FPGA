// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
0aPKz/IMOeE/ZCGpeiBh424a+cD+ROWw/UBDToFyR+11g+nXdQWhWin6T2j86ZnV
pjcB4rnfeNRkPzRfB6hpd4OZivAtMwR3Ze1MrrU7W+mB4tLm3I9myiwn0rCK3ZEd
pDMEooQFJH24D9uMl/uKCLlBzxe40VsQcBp+d9nWKe4=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 1152 )
`pragma protect data_block
orBzucaW1jx6N2YMQNTU9llSsPlXezuwZjFBI6PjVXROYsj879EnDsCXt5PrgK/Y
FG2nNjMc7OcU994Ixlp+Py2GYIrFcbUdi4Y6WZ4J7tbGgBOH/DWErxSDjYP3v43a
aygyPZUeC4x8QV3XdBWRqGtduAONGJ3BRN4WLfeierW1ocotv3sbl1xLooRpFrR+
O4XQa+FrRixQnlU2CMSfRZrnfdKg7OqkMY5mL3nunxXsm4HUQXtbBYqcSZPe2QJG
/2sUJtqSgLjs4AdE7bhhv4hf1p2JUYMlsRNOAz+PsnWNKDa4tpyTN5WN5QToPMDs
D0hFD77dPGHygYClzeCxQsYncrYiNNzOWU6/SmlPTEdVeLAsi4evmUTHH1XuWLe3
ZhucKbs8oLTjean0MtdOqo55N29fiFAySrYr2m4+XujOwMU6gfoNyq7VNN4UfT6K
XUjrTRga11ECsfMZ+UQ2cViCf3QJzGxP5/YlbMLwUlpDoWE6nP5Hifr64MOEkcPI
sLMHW5D030zrtcXbuDKGBIDNgq7uUrVzNkBqvgfelRyOAR/3Fuk3c1uf/LzcEEMy
V2wnPmCnjvHsLhHoegiNI6Mk/QW7J9phWGgAfpNRBE+RCcElnic7dHvNxSNamQcR
qgs4zbj/88BO35d7PVSeyvJFt0qZQqukCDvieLCzwLcYBK1K3BzNsCtszQaw0a3F
6oTOtjXy07PC0GuoEONDsLAKz7alfcyySmXVg5+YtpYqC2gei8GPAREZNf+fKUCS
qzm/ol8KL/OW3NujH4iN67UteuE8zuNy1aj3lXHtHtm6kEeZDyy8fUhHyZExDpNb
sw9pAWCgksQ8PMzAnLxUhPnLhiuP+CsrpuxQXM8JlEkL/nc3pc6yIrOzuw9qZY9G
srHrrdSxhs48Tj5TiI6n0IN5UHYKQ7hJHN9nLusR0DzbcoyMpZQ+KSg/LlIQKM7H
Ls5qV/9pcohW9/fHfiacFp6XdpZ6h8g8ElWsxYV7jCcxhNNR5gQSvYKoEJ5aPHa/
P41ezRndinsDu8UNtt57l30bzT0HXplkjpF+znIjI1Wz8hv8I3NZfUrgIOhoZbY5
bFo3XRiSd9GzKMNAGMzObPCjrqmLZoPV2SXrr3FaoBKYKnwCjqlgnk6k254RL0uj
OCQ24gh5aj9U29rHDD2dxqWNqrX0Urmvi/9UW6lAh6v9iW64Dcc9NnBRZk3/xyKF
BT5PZFfjq15473kWHHT0AoqDFtcOHhNfngUCNB1BBc0VMD43ppNw8rHVpxH+7R9t
aKqJHzxvqj4Xmf83o2bDfQGKMZtUxgARPOzmJz5qftr8zujVU25ZDbeRN9HqFODn
VndE1BDcVG4QhQKPauOq2ZIxLK83VPT9WY/h1UUhrKw+vjxhkH4U6BWhHWpm4AQ4
NEszy7qWd4liJnwevs3iABi54fh5ulOgu7ZmzN5fKkpLk7G4TfyCt1FX22pyDZoG
LKihv1oNKj/GrRc2wBi4Bw08ofx7EdE4W1OgjgC/KlNGiJF0YVgkhZUL0+ggETKD

`pragma protect end_protected
