// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
wH+riZlKnj4v2Wi+LpY1uOP8OmncsWLwhoIwciP+EjMD7W0vrjpS9WCRb0T4dtoo
rdrug7hyIGnA7BX7Purl0v8kja/aOUN6n7y4C4G4BL7XuTK4JsZ9sb7o1EIYtOHi
fQjBb7Sc5/7tdAeAKpmsP16XGH3p6J9uo3gSDKpGO2M=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 15472 )
`pragma protect data_block
loNHoa+fM2FhFoFNv8K9RDla8EZ6N7Qgg32g1qwkw6jnKsfCyNDzBqZI+eIDKCvk
b8Ml6ShL5AEvJKZZbe9wdvfX9n/60LlTTwzuLcgUuMVfVZjUFDillKSPzqGcCFRG
Nqnu0dkIt3AZB0HM4qzuC+28olMeKQWCyMmmynMIKdpcsRoZiQrVyMHtQG/qI64g
SzG50/3yU2JnzgErw5xAX09RVi53j3C+ixQCZ4DGeYz2Kd/hKWBwXYXtGMfPUxT+
06rhfQMtC+k3ZPDpC9fPjdX7loxc8Zj7fhV7yFKC8LGKxzu2CC3UcJZLaSjtDmZV
tp6kI1AnrkS82BA6OrGEQrsgOUHwfkMxNvJJK4mvE4xcepIgrciw8EqJtRL8xEAt
9HAi+NX9Qk5ctVecIATlH6om+tLOys7f7ji6gausXQNHk3iMX773dvFJNqt/oHo5
jda4hTlaVfuzsamaSv5hx3Aom2DeRC69xtFb8J1zuwY8Sg67yG1FrKInTf1kzFGc
Vqq3TPt7RVyGEnHLxtpkJHUPO6x7BdFVIlrGnXXV2gUSLexb8+cbWUtiyMGn/bn4
4Yp7tmI9Dxkpg4habjqp8+NVEKihO3NHGiL+37BBA5c2KpKNSiUB59VicBThfJQn
J4K3MlbDykl7u6tRyIb2DBOlCsxzW99jyfED+nhX4SrtKAo4LdShfOxKtWZOG2lS
kOM1NCrgHNsEGXE/5FqSyfoX6YQo8oigj3bZQzfIgYfEYp/SUXeljXMgX3UqPBfA
QYO8qCtMVL+ZwMCQbSczeu/fwkpZ2uOL54IkMA9r+x5CalVNcF42s9mpGxqfyws2
JWgL8bnEouMQwN9/A1e/ydatulP+oh4rJs78rZG0/M2Td3d7SH2sKO7nIyc+3DLT
csddcEETpcuao9BgPQv/1JmjQSRYVVaISjiIZXkXoX/V9CptnY9LxibvLPmZElJR
9Q37a66N9FcU6zZkcrM8PguFb+CevXaxqXYJfpCInISKW4jL4sG9YIwdKU2uPn2U
JWHLHZf9cXy4WKgv6Y641qPfLQVyG1af+doSMOX4xJSN15nMdH0Ntoh9ZV6Je67A
Sgxb5admuia2on0N+mM92o6/RP+DYwu8UD3u4kJbRklhXJzfWGpuYmpYbj2FlLoa
zeB2l+D5QqB4DbN9SOel7AYPb3usnevzpQFeEqefFsHZbg4eiXDxh4nFY3pmQ2EW
4ux+w9EYjHEnkvuCCkUcT9BocoRHbx+lfUToRF6zOmB4FYDxu+Va9z4lZZjX1lll
3opMr/8WXci3alC684s/IBi3Nh8SvJ5Mb4DE99248+TIhuU5/3nBHLfFkbmvsijd
Hal7+btKLC5/4kwXFsPxe/aW1b53LISD9TAX8gCVvyIHBk4wVb/fVVr3OqnUoRr9
qq3gWrTLV3f3YX2bHzSf4okHgSSgkanF5YqlGeQTnsbhjncuHbteB/gCElfq+G8a
tgOAQpz5X23cijegyOhrRDL4h8bvrfViAjyN6CofwrSXXfdf2+pZJTj1sr3HSs1G
xfbf+T2s/jzZPMW29ZQpr32GmOk75e2kHPcEbOTESwJPIPJkhNwQ2o+CXpfTjRE5
EQMXFZduSkTpwkiQKAag3ojBR7Tim1UR5reamaxbX5NlHH46Lvc5JbhK1Bk3lcEk
RH0b1aSnAidEr0/6Ud3qWuKY+yiKBcejq9nHD19oSVlWuHwVcWOrVjnxUdsVrG5l
5QbGiMhNF6aF8Nv7MbRvTM3tFSbjIy5j+rhgIE/0Id+ntPMqyz7M5zJy+S+yOKnN
sSsEg3qz+AiBUpqzHN2aCRFV+ZsD2JQZLsMpP/7abJ41Gkz1CfnNA09DUnRXcuVh
KTjHQlx5RVRiKr9E02J1bqe5/imJu+phDY1VJYAUpX+85ce+63EY72q2uoBmhBTq
SzIOKKPrEKpmhnFZNe+hTRWYa8MPPbL19m08QcXN8HA+iZ2ovCH5p/xHZa3RenqG
wkh8jCXGPQd9G7CkxxymD8Q4onW0yNGT02MjYLr9BXs5n+W2MOHYOA1soRfvh5UT
c41vsrNJeow/tPsVxdCFhtzSQe0FThHiLmlW1WmFEgQATa55wR8kgXuSaXm1iOj0
wWqpTKXVEW0o+wmkjTjZPzf0IBuIMkST7Rp8CRvXIGEx29hjY+/K3Fvie1/XiIN+
IyHxseg+qGYNPeqMWBMpmbv8V25CGm3adc54VcDkqx90VTPHZsVRD1LjzNfTdFoa
xE4hEG6U6Mg0sJFzyBgKahh2jG2Qt2xCLBKmac/2ZYhNFVIhwwuhh9qR1w5pkQ7j
mCS31TI9U1/V12vOssOUgmwD/k/t0j6rBURYMMF8cAsO7MtVXKGW7W1VwMqMAqfE
fghklZWeDpPblbpp3lJ8DyR+EE+nTtf2+kY7M7RN2d3+s6dMxZdrgYVgHsVXlkkv
1PMpaq3+cAA9EL1MzDKJS6eGsXD/3eMHhciS6KumPAjqI4lgaEFQM9C45wxn3ihW
P7uSdT4S6BGvCdkycXFUqH4OcvyU3YquUVZUrST944hu2kTOvbIsRvgBv62koOXt
ey8N6Z1cvT0DzddfRBg+J+cIdg49ur2zYX/lDr1qRg3TCZYicQs7rcseBt76+Xqu
mH+4s7GGasy9vzixDexudN4NAzNePzRvWuD1XwvMFJOq32L72QyUOmOsEI+6US0G
abRr4RcMAgHlQ8Vl5wN5sjbTYjEFPbfXgl8hJxzKFaDkXJ4rFnBx4L/BzHTNa2L7
AvEfYQlke0dEf9J/zsAlbvelEdDTBorWw0MfrvPiXDXtwTEhH9yyPdedh2GQI1GQ
s/ArgcA49kzWAxPcHeaK7kpGseI0cMTaqiVqQO2B3mBZtXoGChQZweVIsbVIDcEp
fh7i/c3Hz7Yu6NgVwB5bLq+rxp2iXuIHnH6CNMxMSsVKTZDCyuPM62jmOUe+kcTj
Wof1o+mmaEPi9MHkzRg+oDkfl717ilWBM/lXSOBVYz0mZYpqNk4K5DFW73NPxX4K
vZjshytAY5ZMnRAfd3DpWg4sFCbubbQjH3b3XFmxPJUqMdvLv0m4tqrtfGE+cpvj
QtoT6z44W7kVizpua4vVCGef/T2Bhm/aOOsqR47wzoCYcQpwXanuCBbad0c6jPgk
f/V//bdGTTbs5Devuoxt+Cuqnvol0k+4XS1iUcDtvbuR5DtTvu7EAIf30mZbVhzm
6h8Tv+MyU1DCio2OPI0moSQafqKXoQ831kAeSQqx4y9byJJmU0EczAXlpLDxPEpG
xi2sALidsAPLXx7k6hLnW/4FAXRganTkkH808DEf+YZora7Xdol1WTtVrUQwVEPe
swXjqUdLGMKVaWsw7piD749PjjfmwpOSbrOZc2pyEpGk1AKAWVOzu3Z/tCGoXWjX
VX0mx0ImNwb9GoNBLJlHt6L0iyRVul4/oYLK86w/iKUc9lsTdsjvhqnuNQuYr8m3
krUH9fr1V0Nozsd3CKxxGfuY+njoI9T8BYyP/qnCHn7C1gdL7ayd9Ak8ht5b2twd
irxVjUBKH03rUUwAdIwKhU3jGiwVnWHsGIVXIvSoCdFcSvcH9eIvuV7/8cT0ymch
HjrkocpjYBK+jDyG2EvM0LZw38a53Vtp25NWSNaufK38h31RweJFfiWztvK07Rw5
T5+BzLXwHe6Ajj0EUWX0bueak2ubDZLn4nVq/8tSfIy5YBJs6CdOVpcdCb/hnIqK
JMo2ET29aOY7xlz48fpiKRz94m8FGKMI3diSd+BFi53vl/saWZils88uxZqLPQvn
SxqhMS7SFBP1p34jStmTOyrda8louUCTPUOHgrgLXmbJfWW0lNMReXH3rIdM8OgD
Mx0DNH3otc/4eXAf+dUtjZDVxZKajyYuhxmlrd2Lp6BB0o3w0spXsFNTIPKUPxdR
wFGdTjO6bcQAKeKuIFB2F3jLXE4wyT5vaLvMER//3Sx/FhfcbhWt21m4Efh/qf8H
Dpmr7OfN6AVXQaLKpeiUgCUZqlH9RIaSvJhP6tHNtlYJeVMroA+EnP0e6S4A3Orp
jv6oNIixKTLr9UQ2uKqU4Ysu6WESs5uGGwNeFJTgmdIifE3f5MP8G1JsUnla0cfh
0vWLflrfLTfHjjxuhavWPR7njhqxYLgzoDIi3XgNQy4z0HysbcAFUZUGRGkOK1VC
+rLTcQmp3MykLaRRCvTs5Nw7JWCK+TJSSOfmpy6Sl/1GhL3V/Y41qKstZs4ijfN+
HC4O+By3v1+jawWPSM0LM9oM0WxRqz3klQYe37k2gPs77qUfYpl7caamf4bgWC4e
dT3luwRzobJth3N2j/X+MfwbnTbJ2wn5liE8f/XJGwHUOCg+Q3yZ3B6evq/keYoL
lu5XHI9z7fVmlSydLyRfo3GFDACrBXmpBWNR5l+qsYlbgfDQy7GJlH4Eewt86BlH
cfaT/2SfoCXrdghWirQaQsx9raTuzkaGt3BcstbcHNQM+YeWEfxpolaozB7JPLrP
1ACrHR1kMZQQ6MAtsvv2iOiVPTfMdg+Hp8HL7RhS+lrkNqXaVo9dTrnqB9BCAFQH
oajPOj/hSZI8GFbXgBN+cer8HdAaHUfDCEYSIaQgDgLCEYsVfVNDf88WOh52MVqG
fisEO7BwNYyEp+SmoRRm95+BxgotsZpz6PvcSbL4AwtO9lv6lBBEbGAb3IV5qqHN
fj6PsyW/nTiNiUh8OYGqg/HKRNObFqhHRHcshEW/lDRKzo1OcqYls0ZbeX4CGQUd
mh6V0ODOLZvtLxEJVqsAOK3Zkh83n5MZoqJsRIcT+u53vZQlxv1uukQmEJrP4s+c
LRQFUOacU9PN0XcdRdkJ8FddBJUcjTdO7l+ppPV46NLAcmdyRyxtkfgYM/ZopHLB
gG4b4VdQRvAKYjwHTuYye2oj+qpx8in4cY7dw7Tf0MXotI/VVwQ4273arhH32NN4
7WdqJ6mibtxrmxsFPaIV5zp0IMftH+D1VyiVt/akqVosv3u1UCUxFw/Z3yHMvMY9
QBVqeN9Bi+idJQTdwJR+V2Bc1PO/G5b0n91o7ZWprfTku47wVUp6hbbqRWaz52n5
voZwgaYFZI+LrIV9pEH7bco6V6myVYcRYYwv8CwK5eI6h0WsLVUsBDuZbiDW45hy
kCtuJTatGtNAXuSPykPzY6dLw0qNiCjlaazwxbMUUZw8ofhih7BYII030ZNBcEnH
QPIdEN931w1F16wrPghsACzL3eZHf24L+t+Y7wtbla1ATkDX9ORiwuy22Z3X1RDD
oXVMP+CdUWWcXo5a9ig0BgnOXQlf7Rf9vvNturxFCPJTq3Tpe+SnSOp7cMfMXpd3
pBFPReQbN1AOTn5sk5n8453GSA5eXCVk3ystXiG6m/tUH0PZoqp7qZxOkPF5HR5f
pTC3un0+THTeSU1PA5VbKxnSmqkxPNtCpO1M55farZK45vJ+nu9dFWJUMXb2xPma
1ukUTOI3QXA9zSbKIf/RUtYzX0slh3CUj1EnCiwG8WxhqQdNMkISgx/UfsYgBz9m
LEf8CPryVllXUEy1cKFOWGOWMPO204mOMOEqw099y73EgY/vCjwKME4YmoPA7kiQ
Vu8OQQ8l7kdu0TNmG9G8G2IVH6I5B302bapRLMvKSempY3YFsPK1knUG0CqYCPgZ
nDUVw9yvCFF4rYyb5mcKo34FSBY5slFD2bccnve+gi36SIPhQ76fY9WHyQA70u5q
Lx5yGuNx4YSIiO2WFTcddLTuyygA3Dl9PbI7YsWWaUc0HKpiYcIHnlat61NaO//t
O0P6hahf17UG7D+Kp6w+Q/Jp03uQPD8bEbg/tPfuMC196JBv//DYobCNyrdmbC2a
YXyknd0C8Sm/lLXKwM9ovF6qxxlnQ98HYliR/3zV77fqwJt0velRZfR6w2R7Ikcf
9vo732Y4/i6lvuSfvbNwkSPvEjWuDd+9uegAUjTSN2iPHONopwE7EksvOGY+tgYK
Ex5XQH587QY1Ch1s32FcK/YHFn8gLcJNjv6Mtakz5Te5WHN0WEcY1gKX7ks7F6Au
Ufg85E3p+5Q/Cj6YOQ1GodnmwiN8goMibLcOurIFN5sL67YSOz+OKUDgMT3bklx5
MaIa3iV0Yi7Idx+W7hFA8KLPaC3o1Z2C/DaEmE/XeZoOsPYOCYt3SLIxZKau9Tz2
P8UUKM6R8jcQ303G5A/I3jghMref9dfK7db/RIU7/lbAc0xTpVHIlGmSNPDRQb4s
YPx6VlaAZ4vJsNDJzI9lZASb9MNyyRdEGLnFPEWT/lbbX6QkukULU+gdCoRgH6P7
8EypExPy9bPlwnFGJ0TvO3rWMc+OC9KtT3m5mfBz7SrvpDpEgDM/KdH3Q8aBmvnk
fvQ1yqmNyZfnJvjtL5JiZx4ccq6zRioRwklJ1iOOZuHnmhRT1BmSQmsOovEuBs3k
RJpoZOIJU25+ctQxuqhw10tHYXP60z9HBflE0iESReNuEMHlzUmwfTJZPhcogPzp
+Dmj+tB/MzU7ots4nuXW4zRoArm9Xedu3VMu2fEBk840rvgiOboinOkIgcn1oP/D
Ur8u5n8Pj770zzIN9CTHBp+D0Rtlb8ShMy2J7H5jJElx9y5QJ7ghnj6CUA/aK5ze
IjzsZeIEXbUgQAmT4482kk7iZY5Lno895q4Z1PxXu+mhDEQw9NXUU4o2w9UG6BEO
KB/grMq+ZLL+qa97tOQPOJvhYBmIbvLjj0jSD2lbEjdIjAwPRKbZIfw9oXK+WIlc
rS+ti20uPU8VUAr/+GhDA1mGBgrSIddKa/7BK5lr84q78OpnSBzwp8NCiX/aYSOP
EEq/Fp/ucolbHDRnoLcCB5dIL8vQ4p7l6nl+QYX7c7IPYn7j0vZ9KzZrBybbYn2s
s42/zC5NQeEyd8Dy/NjB967L5eh+awPxeyKPc9uqivVzxmTmU7AdBo7cBqrtIvgf
fFzlt0u1VzaQ7RtvZCFlUlxWlIOYVP0Ktj+57IGUZw23hkDlzzi9A2ai5I+dNkHa
mMvQyUPdVk9XTRZqRBcNjsvFXl3yHAF8Q6yFczwatWBi/fAjlIfXjEViI2/qlzjm
QKm33XkPmPmvYUX21AzG54vNe7xNhdkLt3METfyFtoMN8BwCeeiJmTopLniopl89
lWDMsirUg35/du0p8zvpFDkTfk9zAQQhy2QZlIuc94i3LfrlNuKyBgLY1MneS1Wc
Mtz+5QSw8Vwsriyet3X1c4I8x6M6USc+C7Owd0aX6DQBlAVLpqOEXuhQ9zujyob/
hTDXeiNSYx9dEOzzcW5DMm7vLYgxvfU8Hx0KlECRXHaZm8pKBs49Byb/xeWJ/aVv
btFjgg9dwhdVzrHXh9KpJhqG1YkcLqizXL4/40XwIkstJfHDADLDrHDrIOqySahs
QdEUq0ORJ2KsxK/0kMra6Ju5txzzeo7c1MYimkH98mCvkO1Csn502buhuuThRoJS
i46FqTLPR8bxD+3Krj/QLIwtur3YZfsH8YOO9UhiTrxSH61GlgumQh1wL8BhtdHi
Q9TipWbpaPEp8GIKIEG/rmxOBAt/YB4MFPiAIAZdhAb0vnAoUDhz2XxWSAicASxf
/Zzxg48EwdzzPj3lF+4fgHkb+MMIq2l05dKgo7UrvZXyXfNSyvre4YRgi0dmS5lJ
r89d5p5qi6KV5lxbIU8Kjk5IFHFUpjJm4n/o7gul9rsEzj8HSyFufbrRi0iWzGJy
aSe3CKiX1xLvwC2f5bghvjqGNWcU+mN8CNBKRjQoe/qtqKxtCrlHBloE2o30oBbb
DyoMM981QSEpvrlXjQc3ohM1cr6VbvIpszHjWf/pOCgaVlUxCagEfw13JukE3M8y
x3B7kl+Cw43qq+zacBEP2q69K3UZo+1g2JQ0ltndHNSyPexG0eg8ePtLKrE0sT0W
6q1SCvQCF3RZAmqxrTMJcFNWK2pwT6AEikPgAZpzzRUvfXKXE7F+PlIdh8t3lOM4
zlbXDQ/YawjUwfeTybYoeIVuceFAdQhJl4GKqoEfEbUecc3SqqaHZQlSVXEqOdAD
kmqfAz3q17llgZcfqEYytaB1oNSxzHSQR4xXagJkBfSyfHTNf+yYFfz8+lh4X5pP
0JgtPITA5ZSwmSKdVBPmrd3PrKSCnVEt8LBKQ4PeL0IvcOJzkHcMgKg4s4BLxMgm
DLNDA+b8hN+CUx5oaTSkB6uvMjU4CwtUp8p5JACVJo55Ysj9Wj+ppzBKjMCgt9bm
wXT1SBM/C8duydN8L9GKqoCxqiUI5nDYNu2i/tSyROlHRU2lsaQkkp8Bwm3fWzdW
hhupuH6XoNQcBRoZdtmfpyMYQG+pxOwfTgexEq10Hd7TgLVNB1aP18bj0HnDjWfb
Uk5E90wx2Z4QAziAeg3nsVzBJ2FDdr9PuIBxAAKczUyr4GHYLMc5+ipwifq3W4e9
ESZTlVW/vWs0r/hQZtyoBfqmCPjfGonkcGzHsnM1MVQPGi9RQRJl9IPSJ34WWArP
yNEgAYnM4hVCu2pWjd0Wc/Agmh4Co6j9/0zKO79sKu35DbtG7Pz9YHYI07dIFGLa
5rBhkCFBtN3crUSyQWlZU+91Y4HpWRy33ElZkHA4JqbyzLpQHioSHGRg1I/jDAsC
zbfEoiyjPYIWD02/VVHtC+j34Z/NhEJWZ9wLf0gWka+yF+gCSGkJ4YnPJ8Dpjzl/
kjomEhS/ekb3Wmc/Izi9dUWnIqasK5BeQczkJne7naRUx7ASbuMCQM7mM0BM18L0
70Q9OcK1T+hkb6Kjvt9BVo1FDL4XkJNzwLUnNnmbMzaEYI/B7xS4/cdUvFcIVzXR
DGz+dYT8ntdAjHCw7qOukcrMKdA0Hwroj9LOAXygCY19fR6NN8lvPH5uAMk1weem
1SLIWssuQFawosCDTsFXYTQC77AbwimpW6r3iJDdCh1eVziZBBXYTT3F+wLAOSkk
sU7oBpA4fak9xiz1fB+yes/2ZOzhp1LrQlBqXnVtOiSA5FwEll7zTtQoWGoTgyqe
65jzUn+MqaE5Bm5AyCsKIEtd+T7QLTVc8PYSro5nsxeFxv2iZ11xZa6JG9q1Ggom
xuHtUTn0pWJvbA6ehuzFR9wldaFLD9jU19juoL6hwHRQolqWIUUc7fZ5NdCqk/5s
Hs0Zp0EEYlqyMpGw04WZVzMxp3QubSp1N2Ar4FhQV29iG1/1busCg4+ijBELgzr+
gvKAGauteeS51LgP7499ynAr1gkNf3kbRzARDvACnx4k+GtQHQaxm23BsTAClzF4
zVDINfHWyHQOBEs2cfHALsZTYpRLYSg0DlSCq8c+P+6b5otvF1b2AbSTloMyptqN
OfV0F63nGDIIm7KnMfc8hyTdmweFpsKZTGomZRpXX/QBJTZg9lVMLV3xdJXxEPpd
Btp9Yi51eA8dAOxW0vETADP8MAHAYzXWHeGEi2T57XUR/Qoa2ztHOLI/Q6t4CdzE
w5Osq5gW0V2gvI7rs9CETG1WTjPG7G8DTBFFc7mDemJoN041Tt6jRJHG0aU9zok3
nB/44lDHH83d7nAdKrV7A2H/T0SOK9skC7GT9QD7GnKc27h327oaa4UBcG22j+/L
xkntWESXRv/3H1t4lt23P5rjs3DFtuGvgWPvCHjOlDneRl8ovwfH7kRJU2YGUwMt
7r3YiUck7aYLd3lmCShWsDYQQQGFkJXeND/YyZNzt1d3e9Aab76mWKzjwygQlGyT
kYoR95YiocjYmAdIymitr0ecT2GFKwNu+vXkTbEJsVS2b4MRTKQal7GLMo3nJ58P
6x/Pkp2r8+QGbR0fHv7zI07NGW+7gjI4E2K5TqV9Ut+Kn3x2osnoIBfaU3mN81/i
5yHKAW14rIzBqdlrMdxRwlL2kKxafLidJGfJ0MsfmIhHR4sPYJ3hop7yww2PJTgd
vq6YuA0PrYQJ641IoqUdZEmZyXXE/j50ROkfQqLHF7yE0Avi1AGRip2PkLHqmsNb
F6twqIkj2SyTibV8mQC7iIT3ltT51X121sgQSAI2U7aFd45zWlmoDhwr1lmpRexM
IPqhnDmWbVkQ+D7jF1s/aFMoKd7oUtZOqDxGlootyjOcKzydCq7eDJiAn+OmbiiZ
iZ2KloiK2C5g/4ibm5AnzfvmHY3QY0Yibkx5q7JeJ9HZq6Ush+MelYTO3Tw8r+d+
ezSKqBnKVMeRx+jwZEWbBd3lVPrttTQ7w+LW50jLuHYGKuYOb7eIMK4670hqb+cv
0NPQcXwaj4+sI/T0Ze8Yxj8BXxphAyPYcuxNqNMsxJDg8oQZW00nnJUhqAdZ47rb
nIl96HuqZUvU9Zcv6PFfPZ/mZstFArtVHYOjkjBO7MNsizILhbFLv16cvS+B3tvI
d+7hyO50LWTwdJc0PXkd0Kqm+WYW3Iy2lPXEdNGkBgrsEhw9U/Jtj+BQFd9Scggc
ieFILP0C9FDSUMb1CtAfjwBtrP2TXojnAT1CYsikOCA61UVnpMFVjg5oZODdDIEz
cLVIek9w69+G5Z7iNFZBTlQTunhGTj42Hvg3vTAsZO7iQg5QfcFsxL3w0dxn2TQ9
r0WqTaXqxYnfGUf5SBUeGamL9JFBttZIixChq/7V8TKCMo91TerUg2NMVoxkfvnj
k4r9lPUvs/tp3eo12xilIV4PHco6lTQx1tBSfZuqoLrM50A7vvzXNVJsJdfDxQB/
aSQ2202LojW5ynetJAtOnNsEvaePs5JCMQG6+7a4jnQ03r2s5Nr9b22q2ZXvbY/h
U5GW8Jz/VayVxuound96iHDgHgthkJU79lrYw8J6CqM0gvwb12o+/sauLj5sA/yP
haMgkZzDUwOc4l3vSI1ZcYfzIWlO+FT0ODcs7GkypFxHDLPxs/y1uQ0aAWAzrYs8
AGT1fpObogKtW4jw9Z7JGLECrYhz8h4iEy+z31OzvWjiZv55NXekIHU65JVCVqD2
6bboJQSFTkd48zdYzleKfc9C7ccttHMAs27bA0VP5DXagMIFWQhM7DEkHv0GXNP0
k+UOw/SuzVGoxnevFWr5FAeik6mhbXCBrlVzsMAyx2qJZz0QjN2EL8x3bg+s0m6q
OrLWiC0fXlaey8DwxNqmdXrxUJ1o5PhDAW2icGHXP3VEmlnIgDFKN1ZOThx9164d
95uNPaEzb3k13x1JNLbHxFCUeecIclMtsRkpQHH10SLEVZtB9SEZgf+F1cuUfKow
Wlj93RjmPc0xrKpqlbQBIReLu2ajKPOXR8Jsbla4m4TY5R1vAuJpeAZNzD7awLXe
MGAh2OPW4aDsvdmYrQlFkk3US9CyJdhn7wzm9klqx/RCP365IcTcu4fBlU9ZWlw3
1Q08dosG3ZZSdeeyl27pYz2k8x0RhDAiotTbvrps7APx3fM/tKPR9ysi2yOlUirE
5nctWY0Wl+SJ3HQ/q3x67VINmhJuGs8I5M5a+9HJ5QZakI4t/787EcLN3NT1NxWB
CFXrsBgXkaEcH8t2AHS3SG2TOcKaadabtKBvApXbs4+eqPsnN0eVYKFfVuvJMNs+
PbkY5wsrsbrfzNp23qAUF8/zy0kPXGn62bbhVOVOQlVDyMDJxERo4+OGtAuL2ccU
uiX0NbB6Y3fvf+nEG7X/Z0U3nLVP6NkDy3FmpjFtT22+sOmAai8VXWlzkR1+jmok
eq7WtO4E7FSEXvoVZbwQK4jSFkCTOc9NDX4pXoHy7yklTJT7pJ08Qbi6FebFM7xb
Z2dnM5ANGWECtJBjItj8IFypO8ok9IHup+/EUZEpieCIHrm4kisq7qHtpjK7wG+Q
h4xOVbTLjLov7O3UyxlDQETkR56AsaBhfx24UcHQULrI4xdX1LLs6SSAVSnojBfq
Zl1MxXLnuvGXfVFSAGetLRqgaaK4bm3zznErbubxbZv1eZRVEs1BCqOOa4UIkv0j
PZgFJ0RA/L1k+CmP1DEWD5NwFw3JlwCRjPPAyN2Mjxx0xmdMskHI13XmuI8ld5J4
fSYHfFWaKXvdbJ10R79zvvbAiiC9ayt16e9GN+x5mhWG+AG9JGL1B9ZadIhYP6L6
fEkVpMQBtnJyj1f4DN9gi/u6FvPqr+GThfzT9ewZs7sMvbobsxQwiokd3Py2F/gs
GYRPsm9jjCVM4NUEM+3xefX1onma5eJwJob6O/DOq2Ev6uDHFDYJ/GyWB9kIlSs8
IzZiWiltMOQo7LLtNWjdoiBb/wjaLb+bjK7qor2avrPt6n0TbbIPF/mAlozUqSu3
WP53mX8DMqSOhP/+qNE92hy3u7+dq/VogQEmCBst4yRCfbRTma1S0NefNN+AYIYB
KpfLJUZIJWZCB8Dc+gQs0JxhL1Kr3LJj+JBqGJ7E/Vm5GL6UPggTP9N0oiMAuRYD
azwgtsmx/DOLPyFMTOIIMWRtAl7P5h9QwSjx6h38RoC/1O5gq/0fcnnHpZZS4S59
WmGmE573pmOLlKgIIBlk7Q1BtP1Ucc0oxVnjcAkVgWEjvSOTOC952lJ2/44o9mxC
nbhau35tvsUN/F91Ct7cymVXt43237/04phnjJ3e5QvpOBHSP5GpM+gyo2MVC1wu
Z9ke1eni0iCwvzGDzhU/AKfgTgwJRuJB1rMHxjwN6kTszyBz2mO1RRD2VuBOUHfr
zQE5OWalqZ7HgA4T+lvu8p7kgbUW/YCppQ1hb6nNMQ4FmfPXgwEEEJWSyxrkcZIA
tHldijZjcwwOmI34nrE2T5yAWHJIIJcRbAQq6URRj0CU3HuqjAODokz9Fhh9NPcc
iG+gfjenN0AuvXW23/XOm4X1dKUOiKdH3OcLN9d1SfE67Lk6c/prWKZdZyqu43hx
5mp0a/p5zQw+qM15E8lSElbFndRSJ7Msk1/6vplwcraIcQ7OVrGMW3w7AZTI0Yxz
TsH6lrzhF1oZazuBZl5OJ8z4QToWMt/6aLti4Ta+EU1UDzQAdgQOfaAAR2MUZCL9
FJrxBNDPvrk5B4cLYsp780IGOJ2WJjchKUxsKlRUG3Gk7oMlO1+0tNg0pfxrZz2c
AYAwFLqCEkv6kIz1YZ1izDJiBLYYcxCc9vbcnywtzs75DbpsQ0JfPu2tPu0Ldi7k
qkwuZ2ZosZiMYa2iwgset5XYheEVpwrZBbiSmljEnzLMYTlHS7PC08/Qooo6KqLs
6PSXNUB/8jT8SvwgetBsJkIgfNEHUulx8ne7aVK5ptIoI2L+UBz3fYTF24yR+F2L
lq+JUxmTKUUOlC+qEnBuIk/0ROvwW9//Gu4r8geUJWX69uPExoEXMdFhk/KJEOji
Z3rvsir8rwFcakVbqXIMRKkPQ9k2ueAYuZcmKxpDyLsXAKAkfqAWwTXdGKuVEwxu
if5GOkW90l4jK8r8/ONuxeV13UgNMLWof2uXLlTaRZXS15vUwUBMqHt0lJvXOBwL
8qMZcVQxwHtfbBA0jnTbY5+YruApq4rBgE0WIZHolhK3F/et3oQ/8iXPdI6UEGbV
gHl/1/7DyMhdvgdVBaxS1p5heyOU282bNm/jLRVVIuNpbbYEUp8+QO08EIWNexSY
ae2wC72GSbAsH0Soe5LivyCvnxogOnNArdumPhyxF/4UQEm4rQW1Vhf8TIevrR0j
fRts4hbPaos+33Q5vknDQC7L0grVx1z07I2vi5eXfi/stnsJklUid6U9Psaz2gle
LTWJsZ72ziGDcEpnUYUkIKvUHikM5poUkXm4BomS4MAQPlFdCdl12xTezn2RUmyY
xvUSX5YTcO5Q5pdP6TjOrgtrWd4axY/me/lete0lz3MNf7sR7+yoKzOvJCefdNZC
mJKoYmfZia0i2ZqzTujns0uIiFhVGFEQ7H7XGrMzF+daXiRoyPFVyHDlcnelEvN0
QrbGzmWHvCy842iH42vF6/ZOQxN7ROO4bj0ZCgBKcyMbT+paLEFyS7FLKXO7EbiW
O8rzuCg/XEnkJHIvuCwWp2CYBU4nr6gC16kFcX9MDOnBs0kdQSFRD7irDRqg9oc3
N9fnsdN6nJSiOKbwYs0Jx2D6BdO/jccHKM4RJVFNtpXhYTROeCMfGn8KOjIuDGkt
KW9bxrmeD7AVUfyOx1cZ7b4n8bcEKYwIhKBGEq8mfkrd0UVNvbJKU9b0FsfUWGsy
WBjjoJ3539SA4KjDdwnyyWpSEl/ocy81IsGKyRD+nFUHwKtqmJQo0W2hzG/vYf83
TUGZYToTOHNz5VeiuFUsJaWhh9FgaqukHXmFhUmLBVlzC+PNcVfrDflPhFZ27DVD
8YC1jEfGJPWGvFlz0EmUsUViOi30UvpHEQE0OFCyBIuvGMcShb31nPbI2lZi3sE5
VoOMYsevdPGR5LjMP1LNyXYiYK+2j6TAcLWnzE1cQ40vkEfTFIU/r2SM3RLPJ6FM
RWMUXD0IestAs6ykBCN2InX55TbNPRQXT3Vrb29gJh/S60FnhP//CLsktdPDENtH
H1zX1A01zNBOxj5ET/0iKFNR9KyJjrhYaSn1jacIwxFnQPaWwm/gcfq7KUkWWmQi
xwvAW4tVT9lLHyHpG3VwuIEn7rJhl61W+Lud9RlVOCQ/r24oSlgDXeYgW97lBfS5
TSici6xbR9jMKky1V4atZDw6AJElVQLNUy1LDUnLHkpoiKNcEU2ox0fLwojQGk9t
zyaNFdwjix1vzECcpXuZJteMudxJvde0rpyRZAQ+yT1KPSYqzCUXfZuQ8srOUyJj
hIUrfqcXVOYk1saeQmJ51ISDJ+BW2n6r4bd++hTKUg6YJIXEM8SJmbQBEkxt03sx
T/bfZXy7na4S/Bmct8+NJmdMCIaP2Jf9q+mJmAJSpaQ5epOejxHUbVIgey+YM51Z
y2U/aaTpV/IulosesOSa0QLO87nE5R96NExD0nPzdjo2XZOGmrJmQ8E+FfrtCa4F
xlTR/whGGzacUzhMFRQK361PYtS8WVaXGez9YGqEC05Dkd6JFyhcf40028LKNmYB
pDh8+8nhJcZbrXjTJ3QmwZDSjqchSDWiZ40kCVVaiQXVg7uP+Nx1GkgR9C/Dn6oe
O2eGQIBj1g6hthMZKpvzCKKMLtD4SeC+mwx5iqA8onY8uWl4JLEnpXqMjZ7FOtKd
QI2S1mh42lIneqHWevEb/GcrektdQYTyALTaCqP7l7B1eakAZeaijxDNj8AgukCP
X2DDKy3ugBwNb2nAr39z9nJSmX3oSK+TTH++238TgpBfollZ8jG1ceg3jQ6FIhEz
+Ainqr3U+Ch5qbnm9rDVSX34XhInq7TXF9rWS80H+eZLrdERAyg/PMz5WQjLWlZD
XChMdzbG1bkPK23B+cC6deUVsULW1alpo3WDjm8+rUkvthvl1vf5aLfzsfzhM6Xl
asJRgsZ/+IpM2ZS5xJuZqXwe2zb3zRSW5ojc0lNAyqU3GUW6VsjFFRyRFoJSeWM2
awEqJnqPzjGfQTnLvtJWdoZhl7GUThE+M0zbCWR8xF97crA/2ZQwHeHX+mTCEK+p
TKgIttheNUGzeNeEZmp7Z8wcNWe0YNA8ZbVe3PwMMvb/KYqdlrCmytj28TFR7jjy
Ez/Qg+7R/5UsANE4Wpo8Taf9pCOBRcMVY8WQkTP5CHolmZYSOg/RyPQ2Mx9+Ns+t
j7S3NuwamX4m4HuNVrpHqQXfazoYxnf1VwAizSGGhg8bNQJmbzH/4uF9cLwNyGYk
FnlI12/W0ZDF1oacszzIx9v98BwmaFVg9hdDUMpWMfsXMNUUoZtCVE+HplebloU6
B6GT59A39b3TC6ZKD9WDy/GZ3LDOXEtq8kDlv1yaT1ei0LURy6Ri9Qu1SRfnw1AL
ydwseOgCU/Lmre0f2Om222pKgvJa1KJI2HB4PJigDlbXVxj4CylnderI0UOuILaX
uBU0/tvPC0rI5UYPac1Xxx7alU8QAGGf8jl1o4KplsB/7g2mxPC6rnc0VZiYuT8d
W2Z4MG8nk7aOnjDc9VY+ElMzAkRkBz1LST9tLRZq6je2p3emSuwoyDnyzEaKdTLn
8APrnu7LqHovG8kWzoxpipKxVbgiBq6lXQZbVoxfBsy4lzN3k+dguZmRlZoCixvk
vhn2wrHeqioUGCkipmu53GYTatp0iQ3KQzQTa3M8L5tgNmUwWVYTXWM/igSB0+xK
qD8qDMSwR39OMAYadfCwqX/EWHW3jeFdzxjtarP1Bwh1XLneXdjXI5N64SJBrSBg
wJRlVb2EPbDcl0cQ+psph4s4UjP1P1F9AL4PUIkItTmGQdfFgWRu3cnm80PEF0LS
ct+HwLUNGssGTlEuKk3zEmFQUoI1GEWVAsvjhMRcKZa0ADsH8r0So7xLjSrOEopP
UWbRvDYijwoHKpN5xcx0dBZdhRuZTyD4ICj2gQOtNNMm0NOcTP3YnrM8K+HBx9qZ
TA9HR7o/nACTGCUS2krHEfDcf77sAZ9P0sJDkxkeV75PAEmIhhE02oeJPNoWwW6s
lwJfVQ2y8x3EO9OQLNljUg7vCw6H2+Jzt/9CEFR/zmwss0nAsNRnDmChkche+Qak
WIzE089r44jDqy9aMATJJv0l/ByBjVO8kpVIbFZpcaEadoCqM8kFQtUUj+OYTmE0
hQQnZUYTWsgwJx6O5iQL1K6BU1Xo7sToJdqXXY8S6F/+LR8rj46t6OFknrMjQY0W
blaEFjAbpDpb3Pj/kDY3+TYuqjsxwz6xYSHutYA7u4zX5bSHGoko3mV66KQiqbGC
IeaBDWZ12trb07rykHb66Z54OICHZBtA24cKu0VMS4qSwmbGAC+dzMXtPvxDnz0N
TuAkBpXG+OdrHgv53u45M4vQJAURfUjhPMC7RdpfXKqwr5OhL7arAgFDXE1cRGse
jqKn7HGf1X3ITG6e1bLIm0ES4m0RV1hPRh7Ro7BznIFG8tkPG042qfWRMqeag8Cw
WOX2WlWHN1Rb9eAlJunXsq/I/TaA00hcCGqGPw23I3E941ZoYuFh2G8JlaIHKO2e
3JoaDfWVHA9kMUOzOqfInL2NONO7vyap9QC0R7GsZL0+FfKjFf863t8c1INke+Tf
JdRs2PJmycOcdVNVPKnvFKQQUqkWG8KztG8K3SOZNAKxO3sgK8gaS0dcfR26Y+Fk
++6sz7CeyVziKKj2hy0UVEZqH0vKDZa3kNvkfOrJdyQ/YQTuFsOQUt2LCpCWaKmA
fsnL+cO8oYSpsk2HK+V8QqvO6Qtd1sxyMpNB11TpdyeUz3dDGX9TtpSSmrYfcSOk
53UspDivlfgOKR8wnIDjQFyddmAAQbAc1ZMeMD28YG6T9yq7dobFFzLjpbR09SDT
+aAZsK1DC27PQVHyqdsBd0zyxsJVEmxnRxX1pi27pENcxiXfY7YHZygpK3sI+0SC
eEWJoEcFqdshrlrgAokskmprzVNdViwBJFBwC0ondj/BnbijdsGUILzJEJ6XmP7x
Gkox+j3OzVCL9qkjcZuZgPJER3OcUZTMRtZBwAOLcH69uKP2rlBT0zld5zycyjhc
9uDnFNNReOk3t7ifhaVKjE/Z8vqEnzyAmAiNza8jF817UIt9BJduRhJ0OpKc6OOd
am/M7ed0u9jI0iEE6EnOXsOjirSIRhcZmhYajTXlejnf+eV4mg7QUIMQsTNeZKPD
bzcxppgWkVEJvvuRJpBVoft67TqbZptELbTRiZ2STppIObB5PnmBaGQW9j2dyW+8
Uaur9OlpybjV7fG2isSc7YgZp2bakQ/Rvyauf0JBN98R+0mvGvMQ1oYtRtMc3So5
WR0T4HKCdxfk48iPTb9G8ctybQ1rjIyMZLi5yHqItdSfIBQBnU4BNCFaXD/wLF8f
PkJnZ2xbnN8Hz6l36huRhLnnzpgx3+uiEnZB9ssVjD0i2x7/BYoey5wc/drAoNq+
1369hWUce8f0NC7sXHvx+F41XXz63GIUmRbauLGnVVJSHmT62WulUWJ6XqGDUf49
HqiyHvE5vVa/gdwbOdG82bQdoX2vrdc8PhozrkWu86D2WcynfwCSVNMD8QBijWDo
YjE9r9E+hTtCkSMyD6FOPSGjrH9cQzFg4q8wgAXYKl6EXrILNUHpKJ17k/ejZuDJ
UznEpKr9CThI722AB+8jYapAP/45FhivKFYmvTeC61SN8st9/SLUpqDDFqZHk84O
CmOiakVlFEE5HXB++ok8ZdAtwjgxUcfuBvkfeyw3rGnxXfAa/6ur5d3STjwnX4DK
pQgXHeQBPlcdxoheaxRxPkYHldmaPbsWwv8GEeVsTDTyuo5wcUOltTxLZhffoXo/
V8Mi06D8kxvzLccfQO4sMRgFvLG9ZWCeLd4AZx3/Lu1mGPmPD1RcA/NyhjUIzHvW
Dh6dkH8U9791p1r+E9sE41NMU1ysMvP0OkjGswFPbPGQS00xRhgqcEf48Ii4hm6B
/L30wuBGooUrUXNgLXlIenELDFBvCz5TZCqQELXpwSb8BCjOhXjo6sJAB0OP2nAf
JkyfGjbwhBM65VMqY6mGApNgCggG7RNffgbqUT3Db8vIeFSWS2fesDA+jB55ToPT
B6UfUadmbQ/c+P68jesi8q9z6VxEUqtq6tSMwM9Zx45IDSfOeKt470IX7ZUa+Ja6
g2xFFgb6aaRh7TI9dYDo/rBNKcocBIrAN0RrT/CqAMI5AVTVfqNx8vcPyjJyhYFO
wPRG7jAv0xd1H2Oku28jSp6eJ/aJcnL/Do0lRiJWO/+91z6QkiVUnaIjbk7fCjwa
grqPN5GQbZ97/6Ovf2bpTFsRr3ucpxKwVP2/bthEiJs9pm2b7akJvDO82Zephyz2
elzZAhAhVIsOYIoB4WZoIPIUePCX5SYSBOdgj2F9sUL0QpxFHPzAgmYfL3ygUw32
kBz7+vr5sO9VsG0+uu1zbexFb9G0e6qZlBSAzPEaOG6n/Hq4jeP51e0ndVDLBGL1
AXIxd9XPc/vqwTW9tgrJGiHoTvJcY0N0me3qbsyCNcvKWHVoA5v4Zb4HXGuH4maE
T5JKfn9LP4DcHnQWSrT5e7zwfKFvlkEkL8FrpLkheb2izso0WUx3UTLuPyb+C1fO
CWG54lUf+6qTRXh8COyeEt+0HUZl4lEhPPc54f+Lh7IJeHLd6mMmlrRgKaKExCXs
FhX8onBEnQDAiyYlvKpf+o4iwv5QbvAX77UM1/WzRkc0kRO558yVOQB0PJawh9f2
zq4ovN5bxFqHmfSzJ9DQNUlXhSEr/0gqBmk3cUq66k1iH86xNhlj0vXrS4jHjwUu
FI/CMnZ+Gx8v3A7UEcDz2Fd7GXdXXYy0DLSvXFhaHLfIwUQa6hX+RiIls403H5fY
rC77SvXROd/sue+OVNUA97xv+AuFPk9EGG42aHfcrbi7VXJV0nLnJqEmFYyPfRFU
uFp/g7BhOEkbjeUJwW4t/HIy1sIZ6penxruLwvOMXYbX9c2Vc8VBS8FCyjUaoJas
lDkUYxweZNXNX0yfs8OP3yXBMz0HMKZ0hmOKBVN7gnp4ktgorBYcFnlKW6B4QnCI
BGV36oVc2ozuHjY+/IBjCDv+EuKR0K4YxAexhQe9cuH5ba038yDCqpF0LLdIcwPR
1QZNEnsjflOn4xqv8PvudCoHaoUb2zPXMvYL5Aqzb0ZhedyGKF8+xF7CKJxXcM1o
I6ViAKMLu2LW2B2PLi6yNrEf1olyLidTYaW9nFJFGIvEhlPTma3dzZjil6hZvvav
w0cuTuTafLdqrBCpoF1Y4SXqw2uhlAoSMMLYus6tRKvrQvCTFqr+ws4guBBRRWT3
7UkkaRxNM1LXFW1eNGcH3S99BL5KfIKXdE9eFTHzVKJoxVS0WjTIodFioeBzIvDR
2VnY19FCz++NRPr6As/6Rij9/GNkGW6Cn1SQ9ffFQFWOuuQudDAaUHV3jT9Ir59/
jqIHe/DwZwz5swBPjAif87eE8+l7wkE9UtJyRHMo5as6l5ITtxvTe7+txCCctdgX
McgJa8Gq8vo9Gcd+NJRPWX/F9/DjIGnaxhP+aMsJkZQQBfxrOVY6NjRf9RqLT/CR
Stg10LysHVRCAiUQTnu4xACYYcN4yLAtG4WtnpjCBbEPKhrzzoJLzofvk59R+APM
uKTZLDq1IqajbQCJDALg6qgITbDtvNoq29RnqEoj9MkPRPoy792YxouzHTEa1HDx
X7jSj9nsYS/G0Jk1+hD3nJ5l5Q7BzTZND3y9ROAIm/MVZ2oiPmG8onyTlJ9C2shS
X/fgNqCWcoer77ND8JFso6wp/Lm9SjwAoncVJ0bhodZTRIle+A77FWsc3K2I5TmX
tzUsxHILvAdqsQsDKqZdPPiOxPDZFptej0QLwP5dJPGvClv+7LZe5Ch1QikQL12J
WywOaZ0aYDCfGkS7PRGSa9t/z1CKhr4t4NiLD5FftFKLNhEG1Dyn8wwL2xbGeYZy
2SYXYyWTlo5g6Gtlcew+mxe/A9MNdsbQp2xj9mDu8EbP/s3UyEH3x/cNlWJcWPY5
O5+mCtAKMIvnzxX5+ScfqYGw9YdwmRv7mIm5ox8eRbqmF1gDwTgkOgmwAniuijom
BwCvKAM+s0y/psEfuuBUhGzSYJAbhEkIlM3Q9LkZeuIdSisExWPWuZzRXc6tN7w+
HjxmPamSW6NDGDnrm/nckVyNMkiJ6j0Hfp0b/BxdzHurJNAqOAkfZA5llKgA54FF
o/PEaDSl1WXXLqbljLegEcO54Y0xdGLD6J0LLb9K6G2fvhkfD4Vz3VjHiGqgzrMk
DMIgK8gDAAlV2M73xVNIF2Kvq6pMWaP8cM+l4Xh/09swlyGN3zZ4IWGdc8J5kbxz
iQWlZayPKGe2WGpj3gnT9g==

`pragma protect end_protected
