// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qp8V3oNrIMw6xojy7idZ21KpVVWbsX27X+YBrVn47n+xU82JlFeBN6jUy1ea
BhS4EdbhOdi3rbAhTRFHPigTvkNxQq8e6e+doIUMfAZrOLqwCa6hxOowKm7r
4MXWMSC/wpPacXSuStaZO4+x/EvQEOsJwskiqUZnhoRdSSlmiz7S9Dd/gLs+
MBhMgi4yPyL4ZRALlfJ6YBV6LZ67eibtkk7Q7/5pU8rTGH+Ni0Qdg56APsZr
htJFdUPquvhv1YAIrmRDj3BMj/H8FyRxMBRyajoR2qFu8N+8JM3wpjuFaqnt
sLOaeiAK0FOMT3GAWPZpQiXaE3d2brhPM2ha4YxoEg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZWwWRD7d1J3WmqHkSnvINrps1Oa9QnXJisuiH0P4NfO+KFJXIjqS1YkkKCCh
ZWB5q0uqsqmzK78yJ3Ecu3D9qAV49TKpJCha5cbnAgcSlK5puXUHXFienJr9
Nd4Uybr9wV7q4NNKUSG1XDAfbo34AkTXdo0wk66iGWKx4/+urJGnSBWSk1pL
Ow3jXizoOPBxiUf+vOxrQ5fFMPXhbVtv4Bfz0NfDs7ZXAvqr5aTYtW8LdD13
DgicUibJOlfk93wqMhNZ3bRYQqwSvpANRDuJ7jBU7u76Y5gaqhzGHatOPIL6
Gb9up1gEC5EqntFL+9ZA2oJOF5SOEtJ3YSenV2mltQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
eNVNYGLOTLh+S1zxWJXLpsUZS3NqH/tBxJLrb71rxhpL1iTXq+fl6PErvqvU
+v5hTAn7tQ/Dp54AWbGX8GM1ZkSxQUVHgi7GeHr+9z20Lb3juG+zAwBN0L3/
LIa0upx9ZD0KVJUs0qntIXNwkLAFse6fTo7ykwXWxIphCfXR6EmLFpcRO7Sw
cV4y+inlFAnGHxVPXj6hUWl2+DJ/wd1kzePbIYuvya+DLLTi8/AUMq7Wut+p
rPruXGN/X6X+bMSjY1bRCqnmM/Nh8o+79A3zEPojO2PGnoit3JeK9m5mOdGr
Zk8tMXBQLLHla2dGx8i4ZG8nTDdOgVZtXmmVnwRu6A==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
UN26oyzbA51pVuG8HtpnzbLmwXOYmnCgviq9iQ1lcEYxPC6ROdkZAYDq2kIb
F38PQ7tgPlS0qa5WI6QqPTxlg0L9E4GSbqFxU+wLoJIiwCA2sPrcUSQMjT8A
A2p7U+uf/SVKxQ0kk7kGfjnohdOJ/NVuXPcdUrvSVWxjyx5ZQBA=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
HMBxc1ZBXbFIFCCsk0Jkb/YCMQ/9AnNi7K78jDWz6qFo5rEkQ5BjfAPZ2okl
4aEKnZtpOWAAOGu6l8+qxnzZ/0O/lBUZaukPUHyWdeUglCh8QPulg1OSPtTr
xNmhi4dJgaTwQIBTGny0houZGIwQ3cNmb1n5dHjQi9Y6zsUrM9Aau0nk5Qpx
hMFZAR3rI9dcg5qhSs09e/HLYjllNcTU5OvfhaYW+YOeUHY/Fkn9+CWMehgw
zEUzrWaPbDeCuH0AiXrJymErkSfMQDDR3SNAso8xOBOS239HnWswNu+mMm/9
Xv7KVXWVlSqhZniv1ZpP7N81hnU7j7FaytZ9ggGxMyCCC9AgjVzCm3266Zc9
Hi+MLKkUHokt7QwFzIYguivB2NpXfI44hSsAhf5nFSR35oSJEsWhIpMpEoLu
pwQXkeOQAviumbXqt9R1bYIITg9ynWW1HC8lprv2vKTtFgKirAHaJHNF3JnI
sYEwUWtJnt8AEPYUMa862JdIN4g74U0x


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
jpoPb7MuENn5gWvey31GhseL5EyUkyyobq+HitdE0mmKHkS3Wu4zHU5tVqC8
Xiqw59wLG+PoDU/X4/oFNrXwo0Mwqd56IwQuEvYx7mcjNOqa5r83Ycm4Y+Gs
m0G5WCXuhL+t1cIZ/dYwLB97txQDkgYTnmK3SGqdG7Fgx09PpDg=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
k0chjw0gb6ropaWxU7ThUv4YebfGjTkBt6QRGO8KhhX+j6qSzbbQQ8E5mxYB
u+jbVjrOocLAeBn1OLazx+cm8udegXYy8Q2++EESEqDk/wFzxdPvyJqveRi1
bE9dlkKH59a8ITH1qzcMl/OJLsLuBfFJd24fX1iuNw1GFTjKWss=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 9856)
`pragma protect data_block
UJnSK7fhtPPxq4uha7HXGhGqpI7fL6qCRHkNYdecyebQZUhfimnGCU8edLQ/
a5kzipHTsEKmz+uIeOFCEdNQA1xWrNuzcl60jVjTo1Mm1lJnRX6QOoXHaGav
agPjbT3QDDBWA+z4UdxJ6Q6A7EtFtjZc4r1t41knh4RedepY9ax5A5OFnVPw
8P2e2vqW81W/H+Jbbcwm0Y6h1yaAok3qbjrpabvLfutL3jsvTAn9AOwc6qKI
Nc1p1gVRBaG785Y9o1tAz4qDAD8BHiIPuV17MM6eUeJG7GkjKX+drRaB6q2s
R7Xyt1H0GPz5HmUN93gxXUpsLnUTvqCEtzI3HJyCYDFAb/EXl1sqjJu+ahd4
wwlGFPaVqj2kmb1DbPF6oI/w0QT3RlAdFCLSf202jc4Y++oYPxhlU5NHCYt5
r0ndTdpu72hsJqBiQ/rYSV9sPn5nWOdOyHR12NPgQgbyLaSYJVFBB+hIeuTI
vPzs6RFIh7AqiH95qnWxk4HWpDQLxp+oXUf+7vcoVgXoIoS4RNPVWG6OXjIW
GF+mUMuCbmADFC0DIMtCDpIugX4VgBNdJbhow3C20BiXF7nu2Ovr/cq+BXom
XEloW/CXOaMhVXfxWENuXExbj+NeMJLhHwFa6k/WlAxaekkaI2yfQKJaaCTJ
/9R0a+YyBvNY7vzBzLiKUhafMP3tDNSIvRfhVjS60nFJhYh5en4NEFz+MCk1
tTPdmpxKPEkdczwwMEY5qreAQ0AGmheFOmam1QgN+9FXUoFfQS/kwmzKJpDL
xHPXt/g0+hvd94WeU7W+SadLxSqJ/CjdCabSA4kYOS4eZIF3nZD9iExZRtfa
MW1PaZc4+giniWGg///QbtilOnFDJHSjTVj+e+heyoaUoxGPYQsPQfHYDuUD
4SPPmLuKcoH7Enoh72V9VD1urOzQHA4zF4OSpfnoYBxjwNvPQpVNMsDSnGlZ
adcuz8T9dO2CVFUt5nZcNBDRLTrRd0YI2GcfNI0rygJyfJL4tHmR2NF4W1N7
6RZQXJOjx0LonTVJXXTAwDobOTRgd2bN/rRtgQcYLmmIV7oIIKLFSrFXNWYC
/phEojgTFv+LfglsINyTg34JgR4gDLLrZHbpP3f2/rg81g81x0U+0P0q93jN
S+zNzPEBrXl48K/P3XI613nKtx964YS41M4pXC6DlOAXzvow1Z21JO+SjjG2
rqbbiyU8egwJGlK19vtGAtbDjNes/RjA0njizCVd68wbR8d6DwBRE+XqfZRe
62//7WwwgTTovIWJsoMAwRkvZJBY6zAIDgkWZYR3ZS7kW9RI7kafaF9jh82b
HJo9IdHMgdwrss6uhOk7o3HQoBPjcDLoux/REiEcA5+Gmg25XzYQfToWFJRs
5w7R3Hfc7UXkjpxX64F51CV8ThWiFrZBasYFLwQdN124jt5C9jIBUQgKhIJi
kVblBak8uRzIMPFZ/G+aqn+QeuKYbH+J2OPMJEyCoT6D0hR9dEsXN7hAuXW0
xEV4BfonSJ7PAbjjrr0fbo4Mw+GOo2Z/gFuMc7iUQKU+1PPFAYdkYKMEbfb/
PSoxN14R9ah6XzjKCNpgqkkzyq+BHXFsj7PRZEh/2TAztV2asa/jDiUKeHLi
dYfmFoM5JHy2TYG5ieT0IIxzIQeyf2krpdwPDtoTMZUuVFhZo0nfBh5jEk51
XX77NAeSNXb/BI32xbgz7wSkvsTNEwFu6vI/H1KMI/y+iNxsVSDLRk3fq9Lr
KN8pT4FEAFFRkEJ98by/2i7tpbAizLArxsLXXsc7rVIPF0xBsitgG0jjHODf
nOTnka8C1Tf7BN4OqLTEF5AaDTZzD6xQvZRrAXz+On/9lI4/zpTdD1OL2qJY
IldkxYNQE1R7V+mJwayC9G2Y9ClIONx0MRsQr8EINpxUrLDLnyRp3ZvLdEkg
33PxiakocX+aczFnoeO8wgEpyzEzhO/r+piTQeQoO8oL0GPLPi60ItqZNo4R
vz2n0gyofq/77jcNhqufoCmzO54l/ZSbzGo7maF/GR7Lq1p89obN+aix98Ly
9dObnNLUtl5aG5vWxcc8VF/ymXvf3waJEbS2AT0YeQyOmJ0EWO8HDgz2djY8
80K6jX78i4QlaJZE7Z/ECknXMLWWEuUX3LUtwdIDIefXNuOyq7eoAvf6CcPm
PnW6ZGjGkGP7lXw7Cgj41M7qY5NcsG8lvnZIoT1EyoI/egB3DkJZqGbT9x6d
gTzpW15jQOkHYSUZWMFA+SKvzsMCMWyk8M0yKb/zUhXBrLdh54+mELbQJAWh
75Z5bg1b9kUCijiPlL48Qiik05PHWWLer6ZTKFGdUesu8yeMsHJCjPwHtADu
f9Ii/s3mnMVsEAK6Pj/8T6S8Fy6uga2yRPF7LAgLBhJcRvcsKP2/yUwsJZ5j
IsmobOVqL0GwVXRuhRC5TEc4AgIJj9WS5Ww8CfBgTcJ7y1AvrjesBtdSaGI/
Rse1ppBNo/o6QJqQ/vyBlPEia7niZScaW+dVFpcG/V3RiNnfEaR0FVUz7st8
MG4UJcD31QxhLmtOlPWWtdG0eogt20CbsIJAzug/cU5qVVhexDyEm9lzy0rt
tcXFzumeGXBHC9dWRnl25xKzs3NtRAcZ1uFV1xZk7lj17vwMPNbhwxDXiIoe
vgoLs4YWoapqBZFsI95Xr2Y6yT3KIbJq8KNQBtdy2bY8mMGkGc6Ews425UwD
P+AZotek2LrhnAGxVjjIW1bOWVVdIOtE/0m6IPgp3KNdDk16PcsaXBJBkviO
pML+Y2BcHi5xHnuMk7P8+/RYfN3h6Oi2A52y/zzYQIuXaIx+/tUxmAgyk8bI
Xvww502qJqaDILxkHu4BloXnfWaRkAz/FrpD2Uw+1c9VpSQLUw3ivBWeBL6F
qhNh62cqgo0TUrv6oYB5tudriRSBzdyNyLC4hUbXgVk+Xk2bEUPRauwgQtzm
dNWqSjvGMNwGojaiGcNe6vekVswyN7QwppTTv9/Kf7IasrJYzZmPdyaK0R+5
8bM/23WAUvt71Pe6Hc0kliNNnchLWocY8gz6wb6lf2Y6UFiDhnyOG6nKz+xR
lt/Ps2/cErtiVowtfOWZ7d6nR03TyzisLMQzUw/wBYykmJn157qWsN5AiaxA
XhiuPHvSwriVqv1Y31czg3WqUCwSPRwLfZ8rsMGMQAB1j3HDqXsv63hpJG0e
ufccUDxPzFMos5E7eAwLvn8kckJ8ujh6WUizMcwupwIQNNFJiO/6bSCMJgxM
FGsQo/thD8kJ/RXEiohsCpC7HCfWrb0wnfTmeUsEfLNVC6UGvflSaoKCUQrJ
K2xl7KiPuIL8anJuJH2a7WhVREvpSQTSvk7EZx3BeoDFKStYAR/8RMOrwB+e
yHPjepXYbZrMmLk6a9rs6sjnPXtwJnIraaPzibB4rf0nr79RKW22imydcLhU
Oq1g/yqO1VB0cfURhcnjcDygfNQ/oxCFvlm2p//jZRkNe52JdaIRrazi5uF6
xaxaEnpwL6hMv3WtYkeuq3XwXD4DTmcjywWeQ/Fx3/wC11/hqmHoCWcfXpz0
ly4xykfLclbTHuHoTpvXAhfIeD+plZNxcQgnfh9COKDUWeF+shpvm4eEApOK
ozx2q8qF28Cc/tqqbvTod633szt7Fr5IsVefRpwWtDEJzRAPxMejUiI336rK
ZQcwoGqD9dNfuZE3ebd2JppkLKRIlHrXF4yX60wPEnDlHIg3GlUrEj1jmW/J
/aYm0moV2R0QkDz6zniPx9+UK3i8EcK6c4msHrLvWMD0u3kFY4CqoWtLhJXt
2jpUFs/ehr9ji3Gu6ZP741bArQYCUDt5ul1n/X2uobUKyzgzFz/x3ucOax2k
HQpmNpvck77tE6Wvu5srbFI6jpIQ4H8SHUSwAsBmaLbfxTWPGZkVkz9DymoX
Q6an0gNCvYa3l5Ks2pz5r/V5DocnO1Z2vt19+NgK7pP2PF+XvD/aJadNyAMi
ACs8MzOjG879azfIn7zKoaBexpKbRhLqSsE4lG+f8T06s39yVWeWkxOZtlDv
WEQBF46m26IfwqRvFBb6JPGmdK9MId8I2UChGroGLlBjHPGaVLnuLYKyhyvn
p0GsOn6EzmREKYLm2avET8p12v0Si0hoZT0GE3yscp/G8qrun9w8r8cKp0eo
dA5DG75saFBjiRad6QkS3/a0iCrXDwzEk9AVEh3YewT5SDUl6J57+ACCZwx+
yfa2aKyxMvcfPsvkyVmTG2na2RJAV61tUDPY1rW1BmPmHpntuwO7VHN67dDw
GK5PqSFHGC+k3RcI1+OYHswuSe2zr84EXCHIe7u3wKpjnayHrfmHrFcLCjW7
RzK6/bsv+2t4GRLaFNYEjmAMF3hmFXRzTZDlPmQqTtlq7oM4xd3VxGscVDZ/
/k7/uvS9GZFTmi3T+CbtBrrseXnd159hhn2EHYVV2n7+bhqGNgaKvKdXgMbE
f05/20lh6SoRBmdrNN7dSoMrcxGiIk9YXMNwGJ2BLqBns5DB1u/6w04iOar6
sZSdR2VuFuz3CAA05uwnlq8jP/TWO1qnKzxZpgPpVihtuyi7sX7lckAC3uhM
dWXOOlFbbWi0ZqmdNB56vbgglC3iIJlXzbYJB+W1rhOlxbLyLZ+gRz/S5v0E
AaeP7SR29X3+vo3YLANJ1kN23BAUEaKaIOqiyrbGeIGsijmbQFwopBaTqcl/
+6QuVZvjN6+YLHJqOxij2pUTw2jsT0IX8JzLTkyoR65QQePHj9MFs4qzF2ov
43QWUm2LzdBMzUO5wquYHBic7og2VXD15yLtRx2OQHBuMeP2YFaSq9PXWq4h
RDLNRAxLDPpoX2Zzy7Y+AsOAJhv1xfLmglVnGSWp64UiQJ+3br22aUi+ZrvZ
InshZ5vvju/dBJaxUHSwJCH/jNWhtu0ckILU4PgEjDkg0Lcl8AdmAP3/MU9z
2fMBnvJRFO49jqToTFSdCAeVvGEZaIhM7zfDqy4pUXndDd7IQwM/LPlOMQDI
57owb/IVb7zmO/c5ZOfs5MC6Yhpn7iiavbSCCGueI+q6Dq7iCCuOzMR1meaF
gxIvQiMjyUBBQx45FftV857P0rIKKd3sGQwR8wCwRt3JP2Kjx6mcp5PZo9S1
z5ldKC0FmuBTUQ4TdN2Uih2Q9zpc8s37R9C4JWzgYP15UMr18gqVZB7WI/jE
85gv0+bNpFr7rxgrTHegHBLkc9DutSz/ADx4uKN8Adxg8TEL/sarJnQTyold
gGf7QkB/ik8eAumhBR+b98rg59aWTLEyqtmh1OH98k5jdVieyC6QmcMCTKzs
Ln+ah8SlGUpWcwSCibpRArZaRD00huugF0Y1K9BPl7qWxa607qZCMqgS8o2h
x2TkDuMEEbkUOXf7pk8Cb244EwpZ491il0TYX1y1n/hhNkDXgiZA7qr9gWGw
sBBHL0AaUyOn8GKBSVymVICYNLZB/1s2LPehS6ORYcsVoNZF7z77RfMGPFQk
BKgKxu6QQMryyWEAxre86np/qW0PisHlpqHHKev5BC2w86P0/FmMLooObDki
bxCmOqpJB64+BcFgniVn668FL2Qm5C40uxDFiXbXBq3tNh6s8OUt+nl29MoC
O0fBak4KPuVEyEPmcoqfGxCESslOYjlCmqLvJBGLwCCRqIV8Rq4GKEfWWQmW
ORib78ArvR1+ZDB/GjizOE1IDXTjOfYvizgcKF9QAXgL6N+ibfxDizVQw4Hj
xylutnKcSw98O3oPjE0Iys2uQzF7Hzw+JbdKseekWgoHX+jT932oKssczVhk
2ZPkoOzW5KZI2Tgh3nrHew9SXCX5AbKOtF9tj0kVo0wimsXEtq3GduyB9Ky8
w7i6ELRsHAmPsPwX+BGeYSnPbFN1MJ6wjdWWuFAat6EchAErtpl5FVrSgCLQ
eDNCXDACkE4ecazqog2IentApXuO8Zu+90Z+su5spaS4ST1aZmNx2s/6du7u
iK/+jyoL8/9PnblRLRX95zla/1dZgu1xBUPEbvPALWmSMJXUyTrF3quj1iVZ
E7xNJ46QGupK33/DxF6q6rWqpumXxgO+ab/vu+5g1Iuc2XJX5nLJ54s/GhHK
0x6bHveaXQH4krGYsmGdlZCYtR4OeLYF+fCUphjqgAo9sYFfOR899ASarPpx
GfiMmI3xAM0hEF0yaK9rC5wZWQf834VFW98RTlwnoxi8UYOeoAEXsFMqm/XH
PrX5RUVOitArR1trNuMAiZsdSGmvsJd07F8wbxSBbLYhvNnBIbWG9a93qR9J
aGx9A/oaEfDXp6Azj9w7Z0gy0+RKJPfBqpbAL8B/h4K75an9syw1MezjJpiE
A3QTwHK6T+I7wf0AKkxVq8+X1xzeiQkeuSX0EjSvdTzfSkCfs8yy+Cf1y7Ef
UjJCBMzFrZ6MAzERsKex+q9KXB0H8Ua8GvjjXQG2lKw+vIBydA0+PcDXMmOx
RStV0Ffw3oTUzcPOteoDWDROTBtEYe/48CC66ya8cHYEwwngkkQNLcfXkHl6
9dps6Nai2pee5viETMStn9pKyQc4WWqaV4vGOBzyen0w7Eji7lx1nkmrg4Cf
dtrZASjzk5hLwu5i/isDw5uu7TvwWqOvYD9yHdkAVCq1Ip+PKMJ/HN+LcYDT
5H1kRD0G3V14dXTEW7eu9dHgK9lSEyO1pLH4Goa9JX2DfjTXAfQZSakMl7cQ
kBKXemgDabobVUzjc8L1eZZFvxYVzijEHBrF7Tua/i+ajzKTtWmtUNGmH64g
RWO7O+trN7uDuNeMYdSebkNr+tt1UlVyA4W0hV5RbS0E0qS9++H7+FSUVnvi
gztyKPOpfOhnThf4OydgtP3jNz9fUwqisPMpMWQU3A/EPkOHD5w3hm7QfX3C
uf9nbhtPu6OtYL/AhKKGkQli2KpsC7KZbcvEE6N4vodMh4h1o8KtOCeeZTUC
LKk/TeHY9dPQuBflBTzfmD3lk//u5DR2OiJDwwIklBZjcQmQQ81eJc/LdTVg
o2xRU5QzxykQsnOi0BkO6qjttAdg9XiVqoyVLl3RkCfha+IwvEjbEgCZDgJp
Fj2LqPir4vwLePT30Ze2DZlRdM8W+0CnA7nlieMYce5tnXRPNGUbbrkcGRkM
KdcnSZ26tCRm7tX8ZLmrle+KSSRwbnhP8wxfefSTYsmBLe9xEegN3NwfCiRz
Msibd5Jbh/724KIGrys9/eXFtCOsrnF4a5bMVDxqFfMxsKhE516uysM9U05l
VgumzdQz+KUeyKoNTST1tmh+otAfUQdhSyECxR/1nqTM7QTbOMEIDyzSfMhl
jblI37JuVq4XlWuNXC3Nh0d1p5DR4xzHe0KXUPczZ4MZkD7w9RgJqUYmhgAZ
Znda0Z3gvqmfiQHPJs4Xvfdrx6J0zm77pmOKwp7IfP+z75Nhuzuf5Rxh+MHX
2wTdt+Di2NXyIGQ7oQz34rVcdVtNK1x7l/dxxF/M8IbqGYzH9gETxELVRyDQ
45J2agJ+GqbRRfNC4NSgHI/e0yL2LnHZnKXlA9lhSHalrrXsZ8y7z/fKv/G6
6V6G5wWrxn9jfPUw0fdF+oviQkT8tmiNrz3UoNjubaDJX8OcoMpjtsL82Afs
y+rM6pL62S8kvomvU2pF4od51VcdYl3vRfo4Bd2YmdvYQw9cKGC8s5uJ0ups
+4q64CzCktY4BJkeFjOZM8JP8GEnCNUT1AgoeI5IBYAiGc3v5uTqgAyh9IIJ
pY0w1s04yt7auLChowmjRI5FfpPdHhBT1BMUC20Hyw6dXN6D3RKfxAShTNys
t2IOPj8sWhMSRmTyT/AY4pPIlcAKTx5GA9QnOQvTH2Y1Lm8517vfH9jHBRso
xkQTtSWM5RGcP8mm7kQNHiH3hgdJcXdRnIdMrmcpc4bvqjk1QMTlnfeUqW4J
zIDw90Whj5u4gCv2hJWJ4bPEccuW42O+LxM8QSFcM2BS6mp89DYRYNSdAe9j
pN72HGIzwu80f3+Gkzdlf7gw+eReKzHEuFhgt7iIcsVjGqbmMcYdhNgzFzk0
Uqp0SB6O9LJpLmTgxZAVRGhmsx2Q9czrK9EkhIZ0RUTh9FUeMCM+quHKBhtB
Cbr6zIcOOS5RCqmrnjU9tFpeR5dAVXwHdDCH1APPfKPhp4lQboVAMkq1MV3v
5uiPXjYna9A+20j7FERoEiqmSC4gTOAK3zoQODF1z1rOjH+Pfi6T7sQtBRi5
yzt/fX7mKwDuQZY12wwmtYPY7Gebej62XnrfH0tNEUtyPxcrI22TWi8UOJRy
KNjAcxW7YiBM2kg4SRVZ8W2O4hNvGNnounZY3YAIHQXFf2rJd4PALHBYZM7N
ceiSzg9jw6a1iDib8ZQRuPlzeYnQ2TP85t29Bi6Ge5oJkJOK4NC4FKDroE55
dIqrAHQ/nlYM9O/jl/C3axrQSqHkhAek4oZjzryAQ+KWL6PZkEcMX5DkNoT7
tRFAuY7DDRLs4L+qm/zKsfQc/YFUql7k2WC0G0Gr+N7zFw8iTt/yNowFi9xU
DvO1M23ztwiqUvqwl0WOVFIVaDwyBEIQs3WmbNx+xWDILA3llg2SFDZFIodO
Ed1BEZj0PEGb4axr2dx98qYgzk7lbh4yRZ9UaBMAcczZYkb/UTahSYoIJ4g6
plSywBo8rMOu324Nity0Gmi8ipKaa7ihYpvZRBdmexRf+ZmAPWrJpW5plyUp
rbBsWa1mW4E6N/7zWN7CQWH6ZeJ01EBL+iiJQfc6MSPEwQgZLn0pm3snWd10
w5KbWoaE7MwNFi+eMXN3Z4NtC/Ej61BnPIODaTNfkH4CeMJ3FMGf+6k1kSL3
fQgRYVNlwjmIMPg39uSkxYvi7qrLUd2CzIIQaUjt/eJeuFB7wFouMvgW2qa4
BTrybfjDiRj48T23KZjwV6ZpTVcL74slBrdkxrOy8xBMrmXV5DW07Mt7UYI5
w1Fw9l6VClBH+ZvJbQyfwIwdDTM4Wil/+tuapfnWzfXYkCN/UznB8ZSa4agw
Ee4piNX4KFrcZx0oX4m2ETWP5n5/TnwvZhr2TnsiG5sI9OM/rMjgJgjyIfno
nB3PShqhCKBlxtSnnwiKRyLA7ryWiFD9DZDGcfBwVTtv2+HhXkf+XZGVXalq
Z3fDHHNJzpWj70ezMqWdtGzfKQvSXPse12hjbhz7U4q8fzohd2aZ7gcBzlOx
aU4NJl/K3zv+KqKM6rG1vi+LS887wKyA4D80CQr6MNAtdoYehaVY78Rpkpwb
u3kuqnV+Rz2AchCbOMHGU8l12GSqjCj8xZ3HNagtk7+eiol0LccG2bFsF5Pv
oniGZKidwsWSreKALYCjHh2sCVlLNo8WKT7h0/osXcpYwCzTvVPIcnHT2fap
jUHHSjgT2Nk6mkXmq872ntvBXDUQyC0RRRUNpBJrAvn4ZoHGYAXer44QdVl9
pEVhXujZxH5wMUSij83z5z6lymQ5ump4IqP1mV4srjV58RUknbANrjF1reM5
6pR5jGMkUn59d+Mv7Zp8WEFF4iM5cKq2XEHqpL4lbwdL3p5kEK4gzhM+OASy
0HvwuLDrS9YOeWzwwvVYAN1OIzY9+NGUXriXIpUjLrTcWMbLAlIqtTiMhjc9
4pSOSZP4fIsxJmGaR2rJ3cAIfyVD+4M0p4F6dNaStWcFVy1QIEQr1uM+Mnra
1+Aay5hBlQZ6pwdimRxWTfTDFyhMVOKIGR0mIjxOjCJYsJp/mgsNiCTu+GnO
MNJ07NYXVsi6lGznizp0Hz/YkB1qlTcwdFWpwmzUfLrn9w+vr/C+y6Uzfuhs
qbQeKLGunGo84wev6LmlqbdaNmWWOEQZld5Kw5txoSweFFMALNgZ4Aft3K7/
fvP4nNzUwBrJ6614hbfEPeZOx7G7vgPNnD9TJlNPf1vN2iULwYD6clg8tdYn
RA/8UzH0WJiMil1Jmv4wjI0kJ7J1SwyyeRoM9yDoWE5BmhAhlgGBWuXWKptg
3cfLa8GzUmBc3nJZKBk8ZC79ZO3Kn7jigBZG3kDgzaTeMwaU22ZXxzABqybB
3sgoMVv24qIwm53FuyNIRyDG1XFl8ov00rSNhjLXwK+z4x12e4n0L6Fzi3/V
oEnnITBsCSOvKLoKp7qiV48g1N2BIf2J3VUFNsO5njUhHBQ4/Nx2BjNLVA7y
tP/iwJo3lUKB14VNO1o4/PS1dn7HKUHitetMyeMw44rRawsm7eFPza6ZTrh2
rjLPLjWtyfe7n4324OpxTc91+rSdGMaIAr8E9pKsM4zDxWu4s2D8mL4uBts9
x6q6h2N3mrFp2K7UGrp4K8sOPQAS7sFZA5LuNg77URfB4kBZ3tXTw+6i1MPW
ylldUUUDtGHuthpf8+HNpcapClUz0YFCglTNibIkE5s4sZal+NPhBrD4Td8f
Eaz99EG4DENTilIBikk9m1vt+99F16dA/HPHPApYVNvUswAHhmerYcYZ34Hf
AwduIQD0+kC55rWCEnsDm0/dFTP5ho5yHgu+8I9plgPHE54eJMvmiRFNj7sS
n4K7Nn4O3CUhltvkCl8nybL2mO43z4pdEmO+Hiwvx85KToszctZ9Mp3riRTk
yy3iV/y3R4cojxuKnj2HDgTq127xvAd0JVfHYM0mTVmqI28jCo59rWqT1FZ8
NSm9ZNggCruXqTQWFxV0YHW8A9JGQy/CVD/lFZ1OsaalfUMB/0VuN29yDv3Y
A8oHZ8Yz2OJEzvSU03FepFPDKdZ4nxdeC6D8AOmBtbIZBW1FPdizJaTlwFS4
qA4fUlX+paA136U2hAPB4dBZbFZ6twopJcuQXv2oHWh4VK+buzUvMidA9u9T
FWrAnpNxRR+GYca1bqh2xbxvExz3W9/AJswhCs8unJQXba3WYCzYBwoJNqw+
eimye8XZaGETNJsdC+LAsfAl3+5LjmYqgfl9ty2Om4jkGkkmlzQWlXGC9QEa
CNwZfGa9xJsoBqAsgXpa7TVVRfUnt/ztIokWIXiVbBtDgJ6iUrzJ9MNXoCKn
Al1xaTR/9fDfGYIL5r5jdxqAvORh7wXGR1n0Flc1xnT6XqbAPapgh96MvkgS
mnqVd07bwB2h31j3hFZLEVVg5NhO+BqtPuppbgUI7P2yEkBQFfb3s1B9s47j
JZDW4vMlgxKnfEIeYiGlt0EwwGYtdo5YY1rAhwoN/fBOO1OqP7b4t1ZEatjz
6tHOjHyPNLg+It6VDvYo8JQRTeup2Mu2XE2Pl9juDEGCn7YiX9TkdbAWUOL7
bkQRPlc0STfPYoe2/VFY3ssSajLmuFliM29QJRjqqUY/fNmZ53luzdh0Plbs
Lrv5txhcSN9PPvfPE21u63Nx3syPmPSPCQdbmVLC28R/0SypT1zNuDUYr6AC
X6KkQzw5krDFK0AjZr0TNHCddRMoPZZZTjG4qpyAedUnDlHKwC/p++BTMNha
MviZfvmbHSJd8JC//qK7uc6/m9K3jP+KEdnQGJONDc4jbXZ19SK+l0XfRvoU
oNJnMkx8TdyQlSaUyrQmZa6BesGTH+ulFDCbl1twwtL7so2SFbASOCAP8rRe
mMCoqCFak9d12Eqw2tq527crWIpDacAKA09S67dWIQY6yHFIlL51UX0G+0in
4i5Xw24QveUDl+BCDh4zjO3u5jQUz9T0AFi1/3/ctPFGoSD4kWbA0lGVXv1q
luW7w/uXIMd0lS+5f8m0FGsX9aHzjJSGrzXKl4UVRuYe/vEAfQVTNOnATcwl
zHC16r5N4tpx1rSTmuEQ+oInxq9/JUphR94tREbGgyfDUW1AZspDFCGinGPi
7xRaJuKWIQqBtwiURgYKRkRFETB1ji76PQZBGo2nFlq1hQeQhjX6rrZ++3Kp
UhuZCive1r95JMk1toxoZ4s1JLrGKxAJ9oQktH33le41TfL2BensgDK1atJD
0lbsd77QiaBxNJpVTlmNFuvdB3q0L1XzEMRTU3yKRTk9budNfrJUTZHl4lay
k+dRx2rGPBr8ozT0MJkkNsMk4A5kB+JUSFH96IJ+O3l8bG6MWTn2HwOYgyu+
4i5DoFAPuB6Alwc8fEVJEv3+TZV7oLhc199xrMiy3UKqfU/vxTXn1EMK+LkH
poQlx4sHALoqd06pGnh+wyZMXtygDnq8vSqFKuh0VVGe6QMCwAMzrYLcGFCW
5aJF8uJ29tI4DpDMDwDzKCaspgEZI+xW9t4ajL3CTG7hZ5lh6usMWD1Y5e15
eLwB2pElAO53uNDnkyu3hXI+SEPpMxWMgiq3/assotjHBgDwqVDtvTkCvA5I
4kRxOlsTj1mvF/+W8+it1TRWLBJwJOQU9c59i2TJF4GY1ni6IVLZL/eGlhal
JJCBVEw1FpN0vUcFXaTIKMsUfyIF7PReqqm1AYffBwgTV0Nnf/xtl6YsM6yf
MkTQMLP1CCmE3FkYcfsI2JsnBPv/xoblXQCBI4b4IWFoI5DwdIriea5EDaj1
2/ayxmO+4uL1NcpFq+bWpgBNUNwLoyDicMLzs5/QxndZhU6aTRPpqyPh3BzF
jKAKEJzHlWzZw/KonJBDNRWzcAmLsI45+poL2ciSugZY7iwoAktWuRh/Fz5Y
PYo84AAKaiPOO0/jHw6PPSsILJMZliM5vDBqBr/AHimiIRmUNeop/l6xfuyP
dE4ButsdrfEaiFVK5EsiwMvzbCrDcH1bSgzgesP0T17nJL8J2BIu2M7EjHJs
YnzFoIvhkE921Lz6CDULR/bylvx9SHT2jVLOJYbNyJKWzvW1vBLzSSyW7iq5
egZKMi2Yh8yLuYK1Kr2c/3mxM2EFkQeLcAYVuVC3tuWC0dgQNWKwqo8kl4K6
zDoDYCUOe+SbDKV95WKb1kcWFUbiEfiM3lxzdZbs6QvgShX8498Q9evIBajh
FzXt0b/Kf6O2P2f02S6+3Q84mppMzyFinvULD1Ga7/zKu5nVhEFLZYlo1GWo
PrTlp+FeouYw/FaY9RLz+9rmgLUXwAZ2E6hOjCtycnafDDM+sR4YYQaLhSKZ
s+uxz7jVhper1jf6nRtvaXRZgJ0RktKLplNiIr+uOe7T1Xhw4yQ8jjZU0EcG
4nDDhyLfwxnQ2DejipYl3P/FSEidvwmXRO6/NUX7RCU9okbxYKjKwFn6+NP7
5KSchYUfb27S3qJA+fzIFJ+l3gLAZ3qNyH1gJ2Ex2u3iyzVfRmc4IK8xN9PX
jHrz0dTsHTJMr+/MPscQdE9FStUTCD3JfHX97OSfVuAPuz3iDvwAx7s8MI+b
7g==

`pragma protect end_protected
