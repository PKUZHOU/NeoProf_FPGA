// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
yz7b37YyiWs8P5Z/NrL9oZTJUp2Ec1K/o9fvcDKp8jaq2a3r6EOxUMPcZ8t9j0fJ
vWz41J0z87xlYV5RHXGXPtY4blh79j1sbx2+QtdTPG9rvZ7WJAKbC788Foxnooe+
xruItqGq4AlqhurzGyiIaNjxPJh8L2WpJyEcPRnasPm8Z0mFOxW8iA==
//pragma protect end_key_block
//pragma protect digest_block
ydUqJ/bmCasFOxnGaLYsujAmAHY=
//pragma protect end_digest_block
//pragma protect data_block
VUVtJhoDIlJ3XvCoOEbZjqXxgS7bDO+2DG/1ztdeXmm7+gmwiTcSlHRgblbAnrRG
MoJY1QRO/E07kALY7LBWEOt0pM7nhS6cnfnzOL/73ovgLTbl55KqQhFjoY2aXQ3v
/cp26sVndDDJ38QL7XUGRZ+4AzBwxcJXUCnZWgDpWYudkEC8ZxgTvOKtijAV6icX
JNc1ayxygyZ7406rMgMOjst99GTTf8tv+sph55fPg0dzwDoaMdLe1xHgTY42KKeo
aff/KuCc2i4DtYtuew9l41LB2aRB3yE0+ydXM5IPszfteBYN2iNx61UXZq6c0e4/
Dg4r7gUsmzEuzfbvvUrDjVh5ZWV+vtyNjzzLqPKvUNvuGA8x0jonO+KV+nt0mUZ1
RTTZWAeIgPY1SXQ89lnS5H30b1nZf9ApF3y2oofHU04cz7/JbL1mV7rF6XAzGbS4
D/Lyog+BGBxryyDyolXQqOoMVn0bTI6BdHwPmJfyA9x5nsLLC0MlwOJGdjfxHi89
YU6ln0mCkq/+6sARW44GtK6iPc4eg93C7fXawvFY4237tlmOkoJO+sHGGfadJQR6
ErYpCZTSMNgDjXG9VIBMyLe/0LRIk85wRKFbUrpq1JH92wK0Jm7axrRhU2pVZ1kl
EWyKyo8VMcL1E9N/EY/1q5Y3xPULF9ma38ijlmpJZ3qVkiNY7SQwaP+soMav78zd
La05qtrjIlF4aXBTCqKrPCX3jtOaCTAYpaeR7TKZQXTjUxtQJWdU+WHiClg/rB8C
f+B/n02Pcs5T4YB7USObHWjXLxnlNSLcRzMiIfV/4f9RzXJJh9Lfzdgz7ij9S6LA
pHS2iCzBQmRmSr4HqospwDKe7z8eFp56N5TqYDpAvJ20AoYuxCRiHuVNqu1BKaBT
TTFIBe0pH+un2b3QyI1hwJvzYu8Naf32yf228T/Sc7O+ThcAq/oRBkEW7ynfmERS
PiMHWfQi+RO7Ql5KRfihp3lEEG+PFIXb4DBTnhutTHcSsM54VrTe45LBBnK75dS2
XXrrVsxyl2aw8EbOctfsVZyFefEd1/YluPhRx8jYADT9QIwgUOizj94QGZf5KhV3
lbvB1ABefbVF4i/ELjcPebg1FTLAFnkt+T/6kQX2fmZUlsiCD0npodtyxWrGSUlc
aq0Xp2xFTiZqM4Wm0qT/rN82auWQ56mQJUwluTGKIs9fmX7Brr4G4mIoOD3emm/7
8TUhRAhSeUjkuCaoU7WbMtOBOclRIdGuyhuAh2HDrmrpynRdYDZB2XJR1VAelgIg
HL3F8qucc6lntU0XOgs7bHFvS5Q+alcMQt84PRJjcrjF6iSU7htBt93ZYfbGtzZf
WiPKHiRML5LfvCID9B/5z005OKJUdZWytT0hsXtykRPW/o6GqVF9bzR+w43EIxuJ
nTc5gfxNNnhNk6RB1gmM7qnuBuC99P9QZSFsAjdspfiLE7mpCeSM9at4pzs5u/qa
LCmE+BlR4PMC5CfISzDhr6ugI+kzM6qbtdBIrKWYp/XFv0uplqPkPcOKs+cJaW99
pFI/pbFyAgNcQV3liayMp10M9wt0d44ISKv31a09g6b8Ep2pA9Vu36nld4c4BM17
GR+5iEnm9qu4FkjXfhvjG66fvgBEzHUg6bVhyA+Mt7jNOSlSYQdoZ22O2t4r8S90
+WvKu2bsMR6dSP45vmieJvhVFOf1uHhqEvz3pMAeAQ0jJ7St6KK6VcAiEmhlJMuH
Z8VywihGvpqiOxzkk89RjWpNsdIOEoaFqaq2hQax4fSQV2nCgvsFrweGG+J0aWZd
ouBCw/I6M/zSkVX8e9KvT6BDTlGbqwAnAyq2d9B+Q1Dp60YZtSzvhwdFcf2Gj4kK
lCB8hmgCLg1Nvuz8VkNNXJ3n1k2a6d+tUaa1CoyKPgndF5eNsCLkEZ8nzpqEzcJy
7v1HGbS/S4sVQNBm6NJ0cHZJcO2LEqqD7hTnByziQYWfDgpcZPtqaf9ibZtfxwO0
faqMBP2CjYShnR6OJkpplCem4+S896BMQPEnuJaUVvVne2HYcvsFESTjXyaYRqvj
xOi19vnmVm6mQva7Bbv1CxHyrH45LLa4RDabyInBvsLVc7Q+8i1aIRphGckpFNKL
pmONExavL6l6HjqIdJMq4gGooV1p2XsLz/qHDaxnIb23+0q4WYideQM3NpO+gGCq
Op34nldcSdBWAJdcGrHqKhoBaTb9g7gj98f0XSXXdiAPgFH49OOfcb/jMJAi1SDN
n16pT3x10Yel6u95RudTBi1npkeaUjSESOWLhH1brhUoeTTwFTLZ6ccaK79spDZu
KnH1XZIjWm94EAPV887oerfffRM3SRfM12MDsdRjCtI1xOEze8hHagGw12RyDDbi
NS/LmBJUoAAojLfpth6kMup2veq+FKExuiCKcG3xEFP6+QK1Z489HsT75R6V1JlU
z+jZ9bt4FgnvOfCT/ToKke/C0eKNrRPrjpSGg5ESg1yxuO9xAS8wdhh5Xeqljqn/
xvIxcQrm2Kcgwtl5b7qWKNeiFmDA0/Jw15yrCZyK+JAzLnvDVEcSBy+BHKVukODd
ko6m53nPizAxXuMoR27cUaAhZDyt/sQovzMad3P7MYQIj9FPIqMjSj4PuQkKb0U6
h4MhZQqt68gRy4nNMETQ74xlwIFgWqCcWV9U8qb7qkPEC3weZXm76tQXboDsKINe
sbMO4iXCb14NAM6xOlTcky1g2gyUyLcfTya5VoRHaqE0vbbx48Bk/rFapWK8NEzd
woepbgMAX6gL6JQbYXL1emHA4GQDVBzbKx8JYE3wCrSWJNzHzRexeEpPRasnTMoZ
jk/++l4uO8TAG6t1qYQZcAZbg1F6fU5k41QfiBDi4CBg+GGVtDuJqzc4sGUseMN9
KLgSoJBDhbVpbrPKtPV48MjDslM6R7RtMXARkX9gMevBSZwo433jq7yutp5Oxk7l
hAiC1FxkVOphxEXyjQ9uck5YaxrVgXSHe7plKoi/nSc7K0wcbtZYZzr4bFDxzPHC
x8pFjrXHNa+xknPLiw3iP35X39U1DNQZxm+POis2pHNuJI7SFVjZqFbk3hNuhiWo
o+81FgWue9iS8U1mkPKWrQmA9SfxVrfGooKjrV/jitey2EfP/ng5dscwcUUVrnas
XB2bDOZiJskMNoI1+G7Husy73UngO6DpLSObQOmg5YXyRaPEA3HLVFrF0lurt0j7
AA4TYcK0Hk8mwynj0TyN7JgdnALEveyZwQn3hZ60j7WCpV+bWHb4aItLVSzVV6oy
4uo1ZiojgaTXIcY5NmG2NuYkaVa8kfuKpI3UVXt/sGCKQfuOP5GvoN55LM5Sf2r/
qP0K/61tTLW+azVrsjffiGwPBdC4gbB51wD+ezbWvtToWN9Y5TjDIr4qXTOR0PO8
eRZf2a4uP9ufoxJZjH4YOdzc/2dh0C1xdJCRc6ksW4wFsSR6PjzeASXLSLSNF8P4
qdvnOJSatkdXDOgucmptJnleRN35KSDOOcVEnMcln0mG/bhFtvnvwEJiH46+zcWI
z4KQij4zp11BvgmsFCMQ83T/1PNWxla+S6fRzOj2BBkmwvDCDXcoBMJJBEreZUhf
nsqS/wzBq8IsSGMBefnyszST5y3cQZBAI44N+BpYfwUbKJovlUPDBP6YnE2TljeY
AI0wICzWdbWUn5YdJ3Dwr3JojA6vA08TG170cVI3zgEbBxoEUt2n31rzFZ33gUw3
b8ej4xo3oHw2gNsf3KBjH5oSDglZkEN7co3fbBll9b1Jebes92Jezt0D3NUkxD2K
VzdLiy02oCt//LWf4SFw/mIVrvjsOemGungYA6GaYDSSmznP/j6hcmI0+senHwN9
9fAqq6D56YErAdfdDL4Esu6v/VeAOxm0OkIEd0bhle41QL2s7sziRsulVD7ipwX7
yaf3xI94Ek8OtxMHNYohY366CBs9ceRNIQSOqGUIrDElng4rabNjljdRfLZqkirj
fIE4vqgqqy6DYKQih7Q1RpHLsq2XR5tbZmJD9pyyfBp/+KvUlpslXBoQ7EBxZPiw
P31+aTUVtRWicHbBCNLVs3Z1y+D1a3Ab2ygwLbiWJHECpKhKSjS3DZsehq2u4Inb
eCM2iUDQo5ec6kr6OylhkmbfpAxEx4Hv+xSN1MYTcZfGgfmMDn3Falw+qTSpJfrM
RnLeJU9A1/6CWrf5aekoXJV2pDgCtlS2VdvgVJkSXftrO9vBDadMS37J62daKnvm
ASqOmozV4Rsnv8cL1N8IfZCL8QIeP1tKnHGxGyz37GfqOQAEt7mLzItWbNWJUbme
6vgf/o7gIEpa6gWMUuKYJ6EzO4M1h2+eFFUUDLGcN2yabWejw6RJMG5GUxRwlBBd
1+TalKmvHSHnACYJEZCNR+Lc8bFgeAaw/OXMV7ehwPoAu77JPeicyBZtXfrFFmIX
8sGGGaT4CMgkoy4fMFOwF1Zn1FdjJFy28FXYL6eXDgSHdbE0JEUOSxqyAaNGg5nD
rdQdzxB3ksfigyDDF0nT4xw1WHswCPnDJhyKocxmas9ye2kJYSWOFBdU4kvZjcH0
Pv7gxJXqjxCUFkYBYfajOpVkgH9DomWwIEV7EuXWGSqDrXTNyzca/+uXE3IxPyZ0
6quFw/hS3pPiRAKRiql2W6Z1QF9nif2uVn8bT/oAoGjQ2b3qUr2gJK861KQ52RmR
sUjnzaH739YxEaf81ZSMhla+xzUYQJSwEPiv3UE01f7DokcdI0XdTvUuNOtx0r5m
Ja5E90VlusdvLGWt4yRqrTyIfBhJvoTQ6jYgtFiG4cX4ifITY1ZhSPoPUjx7ppdZ
8hQ0iMvOGID3PVqT82mV047XGnfXQnlTnjHJQh08ZbDIOjFlzpn7vnrK42AxMFVS
+edOP8hoLqtn2PF1wiU3lb1El+HMxg6h3wzNqImQCv2xoj5nTa8udZHktrWkqQLI
NWRue0JVp8kmAMa2SkqaZ4bUfdO6IIOZbAy65qdzTRaSFQt/Sn8X0qzFJJxCMHTK
LXr+40Ogu0o2WCZNBhjgnjgrWqUySl9eIXEKiXoNOn48dTS/yyOzhbYk9Cn1Dll/
tsZo3k3FvLXq7vYhfBP1xs4Mf2vsvMYmqSUB9Ape2ZLHGsaV8gCJRPYQ02ipaZ+x
ezyl9ehUZVg5FV+wnTO1Is1phOuV/IUAupOK3x/4c5yhf/5fbthpl+vCdOiSf4tj
NCrx7iWjjWwIvDMw4BlDuuXym9STTW1ZwX38IpMtArf98uU6nQw3KXts2XQT9xnj
51tLnHtv0UOyP8JfRR1KUNvTGS/Cz9BR6WtD5qIoChi8gYPjarpgv29VNOJFFrwF
FztV/BUSql9rxYypKNfrdRaDAeE6t9JHkMlJx09n9ZGVjGpxUn6SDAqXGr1Em3Me
ZjYTSD0Yoo/vAmMqcfYfOuiEr1ypOR7/wnCSgUT50xnilWpbVw7Opk+whVluH7tc
ISkdctYrL5KBijAOJRVy01dhnztwdfaGBvVc931FeqKuQpA5g4Ra/04wAhWs3DU6
x3moZaP0TxyKnw+J3yim0Q2D06kwuJQCxSzckplQCJsEmvQ1DtRRwNFVXidjc+Ci
RywkgeLaempgMQnvnVQGA9QLbqn+vYF0a9kxEh/S173eBNha3wsVqbasDfnTuKYK
KIdxjU+EurPep1DPfciXvm5G+neY/HpKDNM/ezqRz4Q1YMRU/jaDDqa1trfqwMnH
Gzo/4uxGpDiwpGeOBGhcSkowDj8uCyodXyxoTMF6EWKFrhNBE4CntNK6TS6/AIO3
hY1+XV897MtNFxH5u60Ml/wu3rbWPfZTXbq9VZVcBNwDCte80qIW/Ih6TnPimmrW
yl7zKdHBhZmLb+/1spnenbcuSr3zs9XnXsP1fPW6cPGndrMjhlsPwSldLZJtFBj5
NTvD+M/8VyLSstpPEyd4nIPoaYVnUmqSx5h5pvF4a/LO9b95D2L4MOyxemSP4F94
PdSQLcdK+MHUwMYD7etvEQoSHBrhfPvUBMXbfFat8fQDJZmNH0zYRWjXda5oJ+TL
d4ViS5RiKsYCuFq8N9QjLxZJnSLqxnlXyIq5kSKbsOQfld+97Lvy7jNWXmk4RQCM
bcCveacpQ8YqCqSACJPcVScuJxi/mhrvCMAbUNb9BAryQBPffpeRaKgenQ+3FMgp
EzFG+1/Jrp6DIPeGAa+Wez/+N4PhIQwe5ly22jBaFEEpU8OxthOQVOKDUJi9s4ao
+qK4eBFTfdL1MlBFvGMWFJt+iEaga+HpDFz52eEF96cU0z9pRfG9jiBDJi4qZHj0
4Me0iHLp5hN1A+MeyvgnztyPCimkbksAT4DNjlJxNYXmIM8tYxJ67TIe2jSQEppv
5GirPgvRhM2hrwreBaT/+QGGk44CU7Gj3ioYCM+e0OhF1lRCnSPX5RzFy+sEXONJ
gyk7Eu9MiCjLnUjcRT160UN6NI9rLA33nmdHgcuHLQUTYguamqv4A5+HPIuLwJ7O
6dkLJOXf5JGlwHOMChvIly1OJd54cKr4taZBo9e1sUuMU4Vnns1AYupK9TnQcLsS
fVeia7zpprV47WU57r4ikddsUqfgGnj9A7VU44FjA2I7hS3T8CcQUTwe816f44eK
xkmNWAYhuaP7bhqIwIVMXS4aXmnetWB4ytJ97myPZfkpbZTGTrTdiASBVIIXvC5Q
Xgex8Tj2/g08TyvbszV31VsWZowgoqKIeiT5nElrFv5wju7BJZDwlYPhpqPE7DQ9
cnFmjDTH1K5sd89BeFg235HVb8YiQZt+teyCBSZwZKfNFS5OV9WfVGyv6VPMnwx9
rsM+3Q9X1XZt8/LCZow4ZnEr6i0T7DpNCGHqLaBTxadCHzpUfyuskcEtTalXRlWX
5BLB7TW6T1/SZdL9EFj7AkWGkusuD60/6WRBX/XuBzCCZrD+pNZiK2bAt2+mTKyy
9WU1T89Qyckw++10bjdLzASiwbSgb3yDNv/gzOqwLKTN1H0wYNv0S2U8XtSKQIhR
4jhiBv8BBQAA0dtBHkLcWBN4wPuDoSLGxuCfnsSICAgn8XjVgUE7e3T6BCN6Ky6D
F8AbFKhBHfd+1rMkQP/PcK5sP+zjj+qASFcBQEd35jSE3F7YLRAinK8YQ1IjX7CG
hwBv7scNf1G+eOOnUbGtFDH9XhIoaq5275p3z6DKtw1xVK7XSJ3qwBGOrDNLaFdu
ea2jAnAn7h9vJNaBFAOkQKnk552zuLowI9TjKwh7D/SmnHjIjHIvorBSmFiXR6QM
4/UMJIjjWmARlC+nKplXvQSbbjuwTi8nfYVEVtVrUQjHhtuUjfrmABOpF9z1agzi
tzk9E+v1ECLktP7o802y5DPAEEPdnMnd71JjNWpSBK2aZfxW5xppgyIPqOdcU5Ve
zUyIUHxYEzL0ZK3YtIoc+sP/al5DIWwZgaxxN4xavLeBzKc9oRfJUXajTZPzQRrj
MrHu7OmkzXwOZ6KdPVKJeOvJpGD6993dDRwNDFHBGwNKykbef4gu2SneD3zxtbuo
9A4hPxkrLgTvsZ6n5IOd8s7S/l2iJCyBbB7eWMArVT7irdI2ue0F4o2vlik21Re+
vkyh+rya9Lp/i/dfaLq+98euQApViFdoN/EQFIvaxgSjSt0or1uJM8y6nJHD7hp8
W4C3L7Hp9tdsUXe2B/Vd25o+WZXvJCBvvOoXWz9AG0Ex+MucoasQMUQjfu0IB0cd
2jk5A3dVcLk1XIyyMwuP0s3kyN2Pi54iDI0k76Ny6H2a19TkFgDuVmdK/N9TTmoB
nyYJ9eoXo9fvEzPmVqLVSdfX3m/J4OjGJq53M35CZGe/nkK4bBPDSqtDkbPJCq8U
fzxt/p/v2CPwFDUVKybpCfGpBImpULX5Zdfx2jmKW/mqnizFYjuTTaxG8cz/fJRd
vrrRy+LINrOzl3O70PJYjoORSstrXynpEKjuyWJYhPef5HSPQguQOCaFnpWRr1fu
xBA+DZjc1z7RURx4wuUjgrBKJCO5I4rnGhwXeBIku3/ktOIWfqKYZV9MvXLlEFw/
o3iNTS9XEocRiWd7DMr1FL8HspQTBKRG716Py5aAfGzM4VDSLP5pGsAC+ePT1Kl/
XvpEieH5C+acSKz/lSRcipKBZGga0Y77fqROOxDODsENFjXHK56qLdpmd2LR7mBu
ItWh/VVfiRJ5PFZp0KsJxqDHWtfzfDlUDIorpcpHucT2vSpbKLbPSxBa+DVJpLv9
gtv6VKjbKmJDQjeqiZwEtqnPvOQd41gKTCkJRaImAt/J8VQ7yPvDsx80fXyFaPwt
twfEFI+ty2n1+Xzs7PYIIGAZu36K5spOlgKGjMyOUJSTHxadmbyg+WEBdydLPE1e
SJ3Q53EpqCK0pwt4iSyghkUUXRTY3qNfUDEqLh1tsjDCQcEZoEwl1+fhgJ/X4n90
vAZxgYUwkG4uMVRMclPPHW8wzoofGqGxGfdiO8mmkuZS9FUrQ1qCF264XGyZ7gam
rZsWlB0KkoskIce2Uu1qMljK7Yle0si6o52uzaOcmj/yrtldranXfVcyNUae4gmA
yMUUqhFv0pUYUCY8CCFaakSiYrdIxBrAaiYo1azvx+GfwCdtfaYUMrzt4zy189mh
X4HzAfL6V5r8t9O6wkAZnHVX0yCMiOjSSBO2yrqzZqKnkRscuM4xTb27UUe1nRya
fDhsABpL/f7ukhSuVkGyQYXyyPrpO1R/5TJkcsVZyVTGvx6gaGOMQY42DW7InlcG
fmm/RVtFuErWNQP4ngIaaAgnwkM08zdOryxdZTKtGKasJxmEwWRGUY+d0IAJORif
IVh9a40bbNO9wBlzvqRgIRRv3gEdNuSzp8xOeQC3aERDg0pTj0E8DSU8rcmgrzl4
RtiidUxY7HfKJdtxJncNSvK5yX+E4lz6ThzKbwcGHvpFjRQZa7kF5ApCJ7KPvADt
STwcyX9aUvnJxj70suTWlQ4TrDCcXtcHHl5E8tizWTegenLzv28j+rNMfSuiIdDB
kqXu2rGFRirjpocfPVILLgcO+8X/jWAWphY4bNdy1CTijn6awT36T/EwlcvystEz
jiJJpqENXSpAMApbccez4VGg0Mhc6mUkGp1U52mlL+Dp0eZfULu3vgcsjoAcXKpz
F2211lgql7wUuunuvC3vIV/wsg6D7Depn38f9DkS3sfrhdDOPBRtabcjwd+4CkRm
2JonKwigqyRG60uSKlM4jS8RQyPC1g0IWgQm22d3lKNI1TJhWLyIuvt1pLTnB9EB
t77E/Cg+aeSQkPcj6bVzkiXjXmQ0PNquG4S6us4mstoCifswHSizaoB9YDBX3OLu
qvmILI9T1YlRBL8QJsHv2HF7uf8gX0P8S6TfTAjBeyRynJHKe/fkndDtSST+fFuB
71XQ0AFcET2ZjE5YXsVpDb2NTzoUdl67+0oV+DIiY+nQG2LgL/ulLBlNmgXGa/qi
jAA+o50nG2dUF9CxtRGwhhJaLb80oVsEBFaSTt8j/GGda0p6xe+iBiiSA1HzOhrY
QhjpQaSlGoLLuU+c4Ki05NSOAOeBKaZ7jyRdIn5T/gD2e8ESER24FWyjZfWhJzQy
ngNaoWcUfjONpeTS5ZVKMH10TcaH48gd1puuIdoXv18d7UkQl/G55DSPCn2bnMSJ
IkGE1s8MTiSWS6sjmyKUUxdN27ArtonVYaPyJUIYqOl2SGG65lUUpMwfbQtAlPtE
LCB04BUiEcD8Qy/+XNRpGB1Du2/2iOZMQSh259iIwLRKZXaF1CBC18mcrtvJ4W6y
Rrc1IAzVf3xg/aWgO4ZcxzE68WjocKpIXBTVP4JEsYj8mCBTEAeHm/bQaVQIUj1i
XqQXUt01dbU0QaWHaT+azfX5GHkT79S/5nNUFDEJ1JVimrd0IsRqekG9HvemSAP5
5vsawMmGqYDqEegI4BoihAs569uMx5FdhAb6wlZ8H9o6+DEnqPZi3aFFvEF9rjaB
U+rpA1r8yq5Zmk3Wtw8fZitSPI+epL5Suz0RtuN/3pse920Hl5N3tAaIThD9S4wX
hzb0zTDVEtyNvIJL3MJ0QTnMtk5wn28A9fK9xwCpqYCO2MIfabvRSTSdQd0I4WWs
3UYovtU5xOQ2luNoWwshA+pWPVQyCOw9hTnJ8GBpJnZW6fM9I2rhGhAeQrWIifSB
doA2IZrcL9IFcFWdO2P1PmIP69KN7jh3vQNSq6rYXcfSHsx2Ae9azMVUSUWIuUkP
Dts7ahCEcJU5ZbQBz9QQJSh25x8De/2wuDlsgvkZroifjO0Go0psmdRcF8k49FAe
2NzLTb6psUOBFi5pv+/3tzuY1wQuACHiwFKKV6+K+cDfXNdrH1yz7OkAzQM0neYP
qwSHYptvqRxJLJrm9hFasMbPmOL46JrMrXkMykfTX3XMViQdxG8/SjnM3acIZyD6
bwZLlsMNLtFCkXSiELCRmPsFfPJJtqxNZ6B+V+cNO4gcPClk9+ghNxcXPeubal0y
v7POcN/c0yMIR9lg7oS91k7P9We2dCYgejqp+VaCWkrg9qbem2lvJt4z2gUOrC8z
gUlzJQv8f9mwuyI8ztb7/cu2m1X08ILoUL1koR59X7H+3hSsRnDWohqwz5t6qYak
rQqUXBPAfecZfoJG7jiJoRtqynhc9o3uZ/CndJVvfq0TD0yo5v2JrJrTQ0oo/5tl
oHjOMoPj8JHpvk/T2OsxlF902hJL+Rpk0KGiKDtT6VDr4rc89m8eZWFI8gadVylo
uOkON0HiFcE34o1iNiWFY5Y3laWhn9X4vF8w9TvZAYN34Teg6GELeu1MhOQx5D7m
u9LSfP/+SagqW6GLFNemOIvGc5TkNJWTySWp5orc/rHJiCAOIMcWfTeqyUYRMga6
2MHWXMcpkfi3uhWbM5EakwzxTi4mESxgq5LaPt0iDwezoRh5J9xBbb88wm3Wyy9Y
o6D6nrXock/vVm2ucjSOMAEde5X9TmFVHjnd5h9Pe8LiMZtF6XrgINHiRyDPuNh5
RcTCjhk4lib/IT9xkTWSMMehum5EoHRITgS8gxD0YmHtRtqFSqNYtAH1KLfd7UQC
JDNro3KCVOVQxY8Wr/0luVXJbo5Un3dZFt532BOf8OUpkStbQt8qbVrnZd94SOc1
Ti6Ws+WrLRu4X9X8kyoC/oI+P+kEZl4ThtkkPOj6ZPNYTzLd6rdzYfkcCLUkKdxb
yhkFYCAZuDw7kOK1hkqIq3EjC2WAFmsS0e87D9B3X/gLaeIwPcraZ858i2crVgbP
NA3fXOynhgABQtnNh0h5c3WNYYcd3tR9oDD7kM2mJOJkmRkHBG9mTxTEYbfDnbwQ
IdTF1z0071FONCZaC+c5WWtxs7EF2iCU4uKghmEHHFMEKxa4N4l0mzAHxm5M4RsF
Jnw1JkUEQ5ZEOcLoLjScnUHMZ2wUS7PefAbzVMMdVX3cc3upnSDrC0vYToK6YFj8
/sREspoxwOFl+x0QD3USscNlj8Z4YUv2Ss+/wFnCWCnOAVtMotXialSrOi9as35w
n+ZoPcssYJP8AO6KSjOTNOsZQhp7ugtyOklKvHNMBDgdFkERYlz5jucBqhJSVCfe
C68gZnvhhCCBszjni9o4K4EGvJN5hDL857TSObIXQ70TOwFTeesRP14mKKsPVP/2
6R7uWdi+Ke6CGvubrdknqgV3qZbjkbEOV+VOL+6gSJ5Vw+d8Wm9k4kF9+R8E2Rkd
B7hi7zhvtlPcmQS/ygskodrQRJmxULQc+oDJmTBI49EeMratCUQc0A0bTtXLEZMP
cWo684Rliv2KIsIUSmbYiubICKQYoGDih7SeOtzPMk6lPQ3zz1e4yY1lwWgTN0kY
8sfOhpoWo2pdT44Lrw645AQMTpmkLDM1hsRcs8dw6ut2oAHq9Qjp8WyaBSlojnaK
e62T/BOSDRYM8S2Iz4baZmdzg4mCtfVXwACmbf9T9/iwmsIWOBW/GhHxRqxy1VYk
GRvJWY57fLHYSGZF5T984vsruPtgg1n03aXnH7HWgbk6hP63Sjw+IXiSAcYu8m4W
zU351vRpfpHDiVK45HHyS13fugCC/TrJXJQ95zviFPUQE9fSmoPdILpJLQFRgbrH
bGnU5V+v8pj2wn+eom/m0ph3Q0ZI1tUVMNpPbW9gS78BFskVwDV0Z/63nzHuOpdX
5IkNOUT3E4nhVKe2Xeq7S0Hsk6yoeOet2mCfutMfFERpKnbk7Ua7It9wMv+SDCH/
G4ITm9/Ie15yR5SPVkL36XKyz0hdonhndXcUBkxL76rbSlI9iasXgqER6LMK4KKg
0yEeyLloeloYG0nl5bGIMDtMEtvBU3LE65sVfC9Whr5v3IuEqwBoeCvq9UmWm84g
FExNzoLkaFAgEBLJXBSaYgmsZ7f4bZ0lcA4pVZ5J5dzFzPYOOnpsPfnf66menS/U
LsUmtXFu+dl+iKjQO6ttuFw8nwFhvghLNXnqyp4i2BusQcKYqaxf4frsOozBFXGc
JDIf1piGnkbLPwzlXVWRy/jKMJAHpmFYcsxaBwltji1swxX7fG87r6x0lI1Ebcwz
DlPZGIrUORwgpJbo0y7eR3YWjqvLq6ABPJgAd+O/Dg0qhVq0QyMjYpOmFasiMbbm
NeF+1mtAu9ewize1Oe+fmS/N/0n0k6HdJ+T9/aOC6T6nUmjEN4mwpAl3/x50pMf2
SZs0vX5B+8x6RKhz8WHpyNAB7SZdmaj2hqVgna/MyxNbHbiEmnvHTWiP6k06xSlY
ESA/B1+7t0bIWls+XvjtvHZxSgIjHO0G/WEVT2p4zsMZy2crv9F2b5UebMlB8l5r
2fcNphZ8ACjk6Nah2Dk2aM3n1H7r1ly172mcfB6gxuc3ILdzXUiPI2cfEDxUQp4b
piJYnk48bO8E2IprdbHyShbtQolRbaGKkQrhaJaEZ1ZY2mhZ9EFaWVYCyigl3m7Y
VZuoPd3eLnDtm9+gKFfk2cEhSc2q1oEJUtPnrxFGtRDNlVocGUcCVujUgSjBbDDU
5GPQVjt//FwhpBStES3D6cV2QOMtJusLBOd4vN+waBZQxktmhPX34ej0Si1nLxN5
pKWoxzzumabqlV3mRUOcX3vrnZTkKznX+o7+ZP0/fg1JzDuIZ4dbbyMdGlj2XmgE
ixUs4PAJP/E4e0K9zy1IeAEwCecxarziKpF1Wfs32pBcC7/ZENWD7mR1bYYkKNAK
DpHxfWoH/O6mUfIIujQFFRn6mAkcTAV5GvIT+YN2wjn+SaflvLcU5IwsYzabaEXH
SbdqCaMjhIBbKXJl4bdnEakY177/E3RXMRrKDOAxZmJAztkatBxyB6XQ6hV0oqm3
W7ei2N8kADGdtOqX7rgpEJf1QXvrSDUvHZR0zAsGQZM+Yn6NBIDAEPPQ539qG/hX
OX19lRWka/DHkcwZ8Yw7OsK6WEpcR8K1gAxAFUu5TUJuhhB8JX9J33gKAD089eHy
Avl5s2eMkvK/XIopsOGzmmuofBdWAHwJm0mdze8TrP8xJpvOnEUD3R69vzLl+iy1
T6tjr/Ey0Te8aePG/XKBRHGvCKFc3509Uqs7uWzDRPz86NIVCa6Gvz7I1NSxfn86
kYo+GUdXpsUZwPi/BbuZy8THCPO+j6ZvcmAl3iiW66PGPYfoTALUlLsCcdvyq3Db
eJTZi3i9EjUMySghYw2Fj2iXBsTan5lfciNE54gNy9+wtac+xcC4sudd1HzIzj4V
a8FP++/5q+6yzVgFqpbC3JrSfPGQpizw9e0xiEpZDq1Vg9IqAZR7ihDU53BrvYc+
2yvj3BseTKBlNFM8dOwuKDkEZTwefUXBN7kZzqkWt+GoUY6/D4ZhAPpeKLtYc1lo
gujjeXsHt4MKLrxDNC9XnoX1+Jrhnl7VEfhAnp3qxiw5tjT4otTPdxT0JkdYFBOM
C1sZ/iwRTC7U9bdxBk0VCv1PSf5o3X2NLai6pDflPrAl7iBI9ZIQsFc2ssELlE6B
hY1D5gFF5WEuiLA76jRSvcOSErkb1nIohS9KlTiUTCBihlOIOIHUnAJc/uup+5T6
SgtrUoou9i7y7QJyl72UlVSJa/h5cGDjuj2V74hxgG2LthAvVSEEMbD61PfzPlXC
StuV7yKt4phieklPMhzuea8Tz/NHK/hhTlWmaW/XHB5ZG2KItnEaOhpo3ZxKEPjr
afLueMbSqhebCL6Be8rKGuEwnSiHHu1dAr5E7swc7dWhWAX4igHFcG6BkaWEQZpO
Y+ebiSOXXLIB3aHb3kA1Imp2czt1BOv0YPcWTl0oJLT9cEzDmno7oiyMwG1/ucQ6
tk9NBsgLojeg0ZMfBdVJTIGDerHJxpMcw3wECw8nVh4F6dyJG6upG7RYe20wGc3L
3p0HvY8kBoyJFniHyoprpOLOLz5njGN+jLUve+LhrtWqWzFFnt+NDHrWQ0BPOgGc
DqvXhK6xPSm0dhauhAs5OajzfwlSy57yz8xJKuFp7H5Kqk7E+LwCZ6YGUhOx0xfe
AxZafKBIXrob7J9B0ukHa9UKLw7kG7J1ntTJKZnCSP0JIMmPToBEa0AwfNSlXnOk
YyDW/AeFTsIm5JjNJdtA4xl294FC4WHlq+3DaP+ow61ThG85MxpGXefXYiDkd+b2
C+Ca0xXGytmJtsN4riHaPqGZZys6IMY7TLUY2S/GR3jSPJpiWLJJ7XVn4nnKf4mP
ccxzycbjv2t61KePE0CjVRtb2GznSV9vRnUMczNBHEXxmGl42d0S13RtMSobdl04
pmfTWI4NsDVTtELUbtLCo4nc6zFPHfrGhxV46dMhiJL2xC5rDTSTgO0SrIkuBRh5
l24R/a+lKSmpUsTzJyJIwmLVxrTpwkefbHgDtKhyma8SjDW/3qWXuG9lsvI16u/w
mk41jPMCvnOJH9hZyCSYdzquAlFYOgYUsYhdh9f2TEKTVVkd+ohu3Z8Y3uVQ1XfR
2X9Xz1UrOMesQtZeJjkHb77PgefD2n4Kq5s9SSOf6b1Hd4hWddyqFfqPopEhpGNM
77uiAJQ/aZAzGOHxK8s265GCiA+agKXUkUAPB8GpBa597Vnc65Njj5/XPFK4MV1a
q8G8yHuwRNNFDp80nslKccJC4w3SUqWdG1wvSlGMHu5S9o1u7jW7u0St4frxTTI4
O6S9305tX9f5BWBDCzi15XgpK/uY+FmPQTDhc07kZ/UjSwVowSp1vNA+xQCdPVy9
menfCabV0Ew3NCNvh+q3H0twSZHhfaa8GfdhB7zEn4Fk6bx6jAgVa2zVXwPZhNiG
y5h3CkM2J24026p5LQrFLRcUgj1Dar8Td8qO6EwfHhFk0cOj/XmFwIcCrRu9kr9K
kUVLXcuPkJB3KnoBXhEZM4sWyNasfES02b7LrdQ/2Y0Jb6E5F9QcDZLnqmInI+e6
2HWUZdP8S8c+tqgSY1y5L4epm23cIB/14uRSUs70x83P7W9TxW2SIA876Um+C23l
5wr5OgN2EqgdqYj0eFeAcUdTLGW6OB1Wi84qkF6H9woU9fFbvHKOSds/aFlkk955
V/BSqOXX/Hxlr2E0un/FeHlCuqkfUzSApGt6+F+V2my4JgzFD784JsnVxmiAObGv
5Ov1NfO68c3I/xYLsbLOspt/j8u+Yqy9EZIT1H/iQHyvCU7QYxoPdtNdANg5jUQY
wCeNyNQF8hm+C6pH8GeQUwzCyMQs/5R2XXo6i02/ETMexmL5sEBISNuFlt+KDniN
duzivh7wrBVgy89smpSZsLHGwfYjcCmoHa9nsOHelYI/75aVGp+dOSJHZEGoKEtx
qHzJLziNI1AYNTpRrlMvyx6hhC6WvgNt8scvZ2Yd2waVLp7ZSEfQACaH8QCTXr1I
CwtcAX9PHAr2WmDuYTHVo3z7/4etiNRt+YQZccIbxMQ22B85ZrU/BFLyfUkORVHx
/LigJoxLnwngUS0Ehmnlowaulp0yo0hZOXzBu8Jp84CeBA7YEY21ViOn+RdAII0r
BeILCMQM/OK1P1YzDpLQjgqvtHnc21pq0IFTvqJTTvL7YJ+Rp1T7BasNIWt15qHn
0+s0qYIr7WCUimLx+iji8DEkN9NcPPbQI7eXC2DsCb3L+SSDDuktA+DnpNHzqYas
sN7cVjgS90mo5b8ujeBs4bEPEGlJpqgm+McJNVVhMT/0TxO/PDjs8cFUeg3plb3L
q+qAAQ7nVPvBVUUyFUGS8olExT6UdF0s8FoNy2/WW6lfVQCDMUzI+ojcoWEGEr5V
EPhcsNXUFhd5Bext1vlfVEPokiSdcKZGjyesWNYbUO8LVMGl1jyO7avMzF0cYKkY
n7qOV8mFpETMEZcQL7LNLgO9VYjamPM83hNAZwYwVXfbEZolDhd5Ad3t70eoEo8i
S2TsVFTRWtRHxqPQNu8aiVIRk7NGWbn2+dkuHv7+g+yeoOvHLy+t8CVhIDK3qvlG
XoMVd8yWgBuL8IYIkkwk3ozaC3rXD5r3b+MdfOHYURDSHdrPqcOwQ90eP5cI1UK/
jin4qyoTkljj0U5iI0k1OZY3lk+dciE1AJkMnOo7FMr1Fj1Lg1O/XYc1vmVSXX5f
pa7qDhAWg4URwefpXbt/mAx4VcSEolWiZ43eXL036LKJkAlbmbJ30UmlonUdZdPD
E+9ibWOZA3b9cuXc/4jAKXammH+WtCjfE/YJSqTe8GGvBkjLoVioeL+Ncf2wpJhz
gCHB2e9sNWlyhiUFVBwTw0g/dNIXKwRkW4xtEuamOJldEodHUGWRkPw9cddZvazj
W7TTUuRSndXi43IZxz4cuIBZgWDktaPWiRWzrhGfTo/dE/Wn3CXYu4aDSXWt6xMZ
P4IoILpL6VUYzuZP5P1jn7rQVDXv4hqh/hw3tHrbUHj3HkmrCeB1N1S12g/wm88p
uLI4bPY9Y5Wefe0+zitsWSKnLNCn46BS7gU7phoumIJjo+5OHWIsSbxQm8RhJ6q6
QsxG3SM61HG1PoSEOT1qK/au4I8fRvNQ2O85yxY4kfQJd2syhFsj9//BzYjsFoLo
4eYG3dstGegsad8TJ/Dl2C+v+yjcEm6XAMKbMceKVJvC3OAE2rmVwcemTV1lmMoy
aH1UzrXgbh09I+pLij5PDvDGdldtxe/twg3tlQbFQN97mQ/Rlq2h10R5sGHZEijU
dLgSUXx/KHsu697Rtn1O79nWXoRqjDG97ccrxTF+QhdbYtn1Ml57/3iWzyllAfhP
XwqsskfkPvpLUp3YMEpGKJAFXOgXA5zDorVIOF1rmxvFOLa9atZzh5knl3GX8bh9
58ePviAqBQSro8zy6Rr1uW6djlmwaUeXkLnLzK7eZ+eaPs7kiHNFvUJ+FpiKIEN2
8CsgBXyL52MP53JcxzwFBLAQJlzyjsCqJZ+C9qWR0nCsALDxHL6j/q+h2rTgEmWc
T2GupIqdAKTODRSC06zskktLkwlEuVhbP8c5N6hkCSr5SOZpj75obHxldC7YTj3R
UIkTgKK8AEY3vmKgcGn2634DUgEtKAsCudOkbpQ/pDw8y7i7Ugini3dvJb6ghhyp
s9Fneo0bsjxUXJfThkftFCqoEUeSxPC7YjcnpHuL+zVhMM/LcrT3CJl91LEc9zl6
5X2ebu/RbST7Rr/2XiAti43ycSAqmCeyttCV/TZ6i6d7+pP1MF5t4Pmqry4rYm9S
l4dyhg2mbrla4xi/nh6ToHgfWr1YwTvJZ6ydT6Dy/0sYn5/BH6ED7/CqHzItszsF
D6TqHz+u4UJ9iLmxDdtM5TK+LVkm3MSius2XR748MCniRopa1dqAw2YJVcAOreWR
Iloa4jiySBlVtJAmcWepZsbM0egcWdTNoPhYoCSXnlRfLuHGC5BaGKcIadaIXXdr
JUtS6boAvKfjbc93UIgCiMxUPoK7E1UcY/483v9mOYNNvWCaYID5bqKRvfKCaYVC
Hr3eYM1guMuyQcrOTyLOqlnwqYJHCs82RXgJPkERtMA+HqVv91d3emoNZkcD2zy0
+0oLAvG9R72JwQf9yi5jqyee5Nlaxu9IrvcqRYhpNnS1NFLKpINh62t03ypIIEHn
nZVkLQxC7Jz2vBEywkorrr28lZzD2yY164K3NghmF/0zW0XzYJKQoSBpKF/kLHIw
QlqFJ5j+3yLCeOZvSwAGXl0kMK599lkYwqK/3QDkQ/8oYSDXR7RSzXgiGHBznNbE
mye0lAK1LyobIhL6mh8K15HBhWZMXToNJqP/gFRBLKDKcTxph1RwzWQsF0zfkOAs
jrUYjhuVvJeks4uYP7PhjUZllcMMJIdNn9dKF37LLKQxDmmHh4k8VFWqgaSWV8H2
Zgr5jJ5ndWIPzES75aBLe4fs6UtRkUVBBBReX5KIMLmYPE/wW3DyCJPeHkTbHWx4
iCVAXib13ghx73MtaeDPy5078BUN1iFNovYEjBQazd6qQxn1lGuEu1ywxu5647EV
rUBm0HOr6HTX2AMkPU6jO6Jz90hCn7F1G35npeGfP5DXUjpbnjafAXSQJkZqzcja
Zx/kWmHTpEsgQd1xdt5YINb80qH1VXZ9Adbs+6iYhBq1abxE0RLWZzxV7Xkxx8Xr
eykWLnwCdnbN5BfH8yqA6qqyITMHKlhjkD2/YdP3h9lj6B+re75CB/JIgPOFqp0h
N+UzIPzcOdL/8KCL1f4NRK4xXvxXhRABqGkFFPIMJXT2Vg42bWqmeAEztNTVvYwU
Q9Z8aMJMvIr3mASmWn19+iCRd52cQuL/GHS0wkifrH9fGJKP3xWEA91Tqi3xDgv2
hoPqso0vwR9XTd+qH/zG14ewVlo6VVManPI0qxmHOPvxMrZGuTk6ItFNc66CaWNw
Q2P9U/FJi78offJ28KUXegVkczoHcusKsVUst9aG2imzyhyuX2NKGXLyhtNb90hd
0woYtHXKASK/QFbmmSTX2P8980FsrxrXUS1PYKwIwb6eVfvLXxrovBKsKIbujbfT
WvMOc4oym3P83Yts8gPkYyKqtHPtGnNtWDeGwuquOoiMtdvh2SSfnqlCj4G52LNY
Rq9XumIeivOALnXbKkYP15jv+3HRJcNqXZ1GH5I56/YdUh41aLrx2ZcA0LcHhH6R
ftvy+A+msIsjJvmbCJ8AgW8i9P8IIbMRBWEQex+Wf1142LEsuQPVmSwotXNBEDYJ
GtVNw8VlHBQ6ryvtFgEYaOCb5g0C1wwW25dm1DXpZi4gBc/aEjjMncBkwVdzvcpJ
YXStCEf4tVy4V3s/yxqnwdYIDMe9xAcXfNWqT8Pyp6+siCGRh5FMRkN62c1X9lfI
iLx47j2/nO3vd1UE9orAjdu4fEDtSEnJLBLj/VaxwVqj5jDLAPlvqNexO1UnEPw/
ep+Vp+dazCsDfmEakvtToJ6GvIkmSERtgZhuxs2i4VFj+69Fou3/FqL7TQqBBDUd
jlCU1e1BTx3LCnx6wrHVPB9nn9E5ZErClW/eBsiEQUuvQLnCQYpc1MupSjhCfcAS
Ab96ZO19sEvxBJQ8HtOrGx976QtJui2bSc20GEwkFAYkmDWx5r9Y0H2PdiFgr7R0
t8477vTMhOjzEkFX18VyUpUN00eRJ8tSFwwrlyaL3NoShajIV2syxlYnTTcUxrbU
n/0WHe/t8g+r5/quOIKBz/5tFet4s4AJmqYLY1+6tuO59QPWxldcbhofjuwVdVfj
PFNgWuzgI7lLrP4BxgiRFcXBNXzmsyqZExxoFcwfYChVlNN7sYR+jhHlBxuGd1VN
U1wAIjvqrejfR2B6mE5LyT6+rcWTSUWPtvY2MFQrwvo9D5nZxSTemfGYnDM2yNPF
wkkw4NwvrDLt/NmeuzeFvfJg7QT54E/lHhyNYGNSqIq3aqwCXrMK9hej0tL+KLug
Nov6PNL/v6C1PZ9loZAvl+lwNAWjnqPSK2kNjQc1oODZvcs7jAPcDdVs0yRAFVSG
YbPNc4MYPRzh2IOo+uajrlhfo8W/dkQjg5OQpK0Nt7VDbcf3CWTcKNh6L8CL7BPP
ooCM8yQyfWXh93a6+hMAqKTbw770XraxGOBQLlfs49zm0EHhFEPvDxRis8gAVgKZ
TmH7vb/Uhz/aJYMorBLqD6ri3vvSuTy33UEmTGU0sLKWh7J0Q1/C4vriV4q0fgeI
VP9TFGaU3DRsqtXdGsrb6WOJ1AGUk/jk3Y72HLnPrtZ+7RVwHW8w24Vq5YPDshts
fsq/G5Yi9rRftRKJdcHWp2B30XFuKRYmAD66jMn8be1f4c1i4QKa16TvhOF2lqln

//pragma protect end_data_block
//pragma protect digest_block
dzADZu9Bz/Sj8cRoKQbyBwnedLU=
//pragma protect end_digest_block
//pragma protect end_protected
