// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
y0x4vAsiPeFLvhOLVskmwlA7D/Dm2PqvOdhD/KEeqpM+eNQZWFCQcv2HFY/Ts74yL//MVLqf8qUe
QCvTpQHrkpEjLojCBfwJHSu//1ZGWl5VecaKB+JsVtgIGr3/NS9ttA9gSjTGECIf6QjoQGdfOPII
FxoLcpC56gf+b5bAXvCuyJnUghFRyoKhm4B1NcF6tiwcFlCjIdmDzxbCzP6v2ARX/p+Hj0uWya0g
fAoGQraUuZmQ/eR0Uah8Qcc//d6v/2I4AfFyFpEkB+WdoYKM+jSX1MuXjifMfi9qIaug9u6Bz3eP
pLm5Xky3/oyHllAe/9S4vDAYF4i6po1ZfJPaCw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 13008)
gsOvS7lKCxRTtjYkDNITBoW/E6JqLzMp/ehlEnK1PGnK6IhJkz6JjGAt2DanrL3sCWx7mkHMY2UW
4D62/WAXM4UzRiRrsqsP56SHulIEqwVTv9ewO8lF3e+xBWKdY4L3Q8u0Ajt6Ua+qCCHq86FxXHaM
vWD718wEAW7FCOI38SuYHJNbWiV9FdmFm1OjTcbZrKPAJ6sJIyEfmdX/tPVnEgflIdjDBV3at1dW
LjCz8bQJ/P9nTb4mjwR7GW1MTmYSvrnH5svcUeOQ7C4sbsRFPZjVBeqLZP6acCnxfXH8EoVWjLGi
rxGBjRaz9HXN5kr/0Uy2BRhoGuE9D5FiXqDJHJplyK+Eg3LVUaOTNrwSGOBww1j9CAU8KvjkKkfu
funfsLoGiNeuRwbFjDklVkqfSCfhgGeESHX1gGdzUJt+KiyvSbHw7RMW8XgiNhnVQq2GDRQ2CIlv
CCqfAyVmvzMlIRAeukSudeHMnXzFKgvB1vSWpXfCqWEwmxuLY4iB4V9DA+xBD4iEBoxx3v8a0kUK
zVLcI+XeXX2EA2F9vg44RcOYTzPcLuveZKlELOXwZgJvDWbvk1Si0VpQUJRDU5re5Eva95Lo8bYH
KEJ0P6GbnwIIyBAAU6BVZXEFE3lI94s67XRaifUPj66Aer5J6cx1+AmAiMFl1KG9zYVQ4lFEUdOd
xMYYVAGLjCR3A/fH30WbauV447po8mqsNCGTlRgqEkEAi009h6ZnMn71idaPuwZUgsQ1J/3LBQ4u
A6JQt90g8xeYP22JAZRFgYe1MMyZe8K3N6yHh2f+yx1HUWDuBQRWDz37ohg80ph+ODVh8NKHFQCy
FkLC5367df93I1M2ivbh8/XldfN97JztswrQMs7BMu8eI+lX6RVcLBg7IKn+nubhGrSn5lOFiosf
rGAR/T/UwUhdXn0Y7Kr5jC6M7rBgaolxONJMzVEKuBQ/7wPqBLZ64NxldLPsC1wdG6ShRpZYmG6O
CoBN7x6NEa7ziePPrHhg8REaH/f6uYytg7PEzVIYkngA48IXr8wJexT60G89FWG3sEZhWs5+WTcQ
Fr9uJ/97oS09rwKbuFBP35cDEfN48qAH7Zs52wH5Fw35+77/PAxOgidKAIRM/ukcF/+rtbL7Gnn6
iyLWbaqTHWiK6lHIRSbSj6BEkak22MQ5BZ8ExkqLIoJvIIdFJHnRMbhF//g5SD/VvWVOV9GIg3hS
ChHGdqMm7q33hV8BFMUPndk5clQWqq08Uw+cgKLCbqS7QX3MFYHrAqhEUD6XbmBteBcKMbON5Gu3
hBlp7hLPUX0glxvoRxLw/TQ02rzEAqsiMhg0/eh/qOST3MNQpUn1ydN0m0JcHiTdcRD7+FA6aKNV
V3gWNSr1c//x/9scIGt6P18BIb+iZTFQ9bLUuc61cqJumR2iJK9up46HHMHEVYUa/I9dTlRXOYbY
zaKY2gxAXgy5/B0hnnziAjlFsgJEB5DbPERpNqQJu0B2YqGpEN1Ob+jPYGxmQT5jFXJGOropCWKi
eG89QaXwBZL51aek8zPsptbKHIoR+LQoE+DAxPjBnWjuvM/Kq+06dPzBrCe31BjzSaGUFV84yfn3
UeV1hAPUDJy23qgIW12fCCOzsC7TVJslzaYBPJPMMFQK7ZSidSdwFX9Mt6YFJPHYvn7M2yvB0H0J
ROw0CO8YklsoOTikfzETw+tf4dWtCwCfzCcUvyaULUhzBnbP5byOLPkRlg9GgVtwLlz5EayQoZoc
uFHYa1UFec0MjWEE/iedriPavSQPU8hIO/k/B7G8u7wP8pg45KvSzUx7+zTk3TMNg32DkGlFTy6O
n30RwY9VB6rT3yqrj/1PtBn5RkRO3YSSWXwyRYN0225fvfISgwWRrGCNRYak/uM8+UHAJwOg+oZ8
y5hxtqDoteeKjFkR1pLB/tBEYF1sQrxORQFxmDtthRQ7QUJG5mgO1YPk90woXZkBIeD//m4MWRPW
dlvJKeTuklaGSFhFvkXLIlE16TF+UpvgfAypuDiDLWYih0kyOCTDvFbImgxEFB/WYfOcLBe/Mlt4
dD9dOjRPLptWH2uP48DFcotIUSTBjYFLKa2Yl5xisTDuAcM90lT3X6XeYmjLNqandzuyzGJj7/rx
iuQfpJcFmK0jvMcJy50geh2WnLMNI6YXgNaArQBGuEnji+pSOICK5zTyOu+Q4OAuDwM+CeDMV9Tl
CAXjGk9SR/nDlUl1ozZbgKlIZs+nUsNe7vVcPk1cp3lWNUL9TK9M1vZaRTT9iEG5yhV4X7zYvhwL
LJ/Fylz8qNDFzZMdSh49rXblh5L+kpRQHpLYnxR451zWCj3x2DgysE5eZ01lpxsbudBh8qDFRmDY
fQvaETbQls2sigC9FzUbODE5N+13QTzwSBiYelWRHVTc2GYX4WV8S47eJu5Bg+gV5IY82ffu16vh
9mCgBPZ0/tRHYKuk+CBIZMqk/lgoW+nhyzXUaoaDR8wo+oe/nHka5q8OH5UKiYQX4tS58epdSOI0
Al3I0L90/7wASO3yj9J9+AstEv7F60pBm+uefs8H6lfL3Gu+iDBkilFFLerZclM2VVcRu5vMuUOf
APXNdQRmA03C9UTVs+dj4qc5fz6bioB5jLJySJWatwz7d/QDDOhnVCzfDb+OACFFKBInZbHxekf9
HADLLWnIRhVzc/MYPckN7SESuZ8G9qlNzIEmcIC4fwSq2XgJxrc8oYZCCyNCvfb7nHPEwESxNC1F
+JzBNgM5FW4CPkJmKTFIEMgpdzn6XYUoQQ5RPk9h69lkubNGuypWoJWcH8eqjdHQ8L4UMHU4wtvY
eC2tqfEbWyznaPu7NKINduqMhBBnc1IYgMUCXbh87+NESnY6G9QbrBh+VY5sielSS1LSbUtWYEuX
J9ywB2cyGZ3uExYccZJpXlsdr175L+xllOGsxLA/WEkV3nJ/pp/8RjdiDgfmuXrgGbmLzizijacf
e764uVciHJVfEKwa4oDPCI/w3HLuf9zeiLAg+sn9jIDE4320V3N1kVx58I5m6Bx9AQ85islnh/Jn
dk9MW6azt7W8jmAOGeklupgRTrhcKN5WD34t4NTQCksBifmd7PGv239jYjkNgeTS579uYRqGrZ2B
KYGqk3sa94uf2wQ/TQ02Kv1o4tkICiPPlDowa1HYDBMRmKJEC2G82kc9TSnLpWb2+e63JkP2w02B
Oo+w+rT7A5hI17sTBSeoSac4Cih+0XhcesDAzPaFPFYkkcT59BYdB9J2jtgGSs+VlTty2lUXcgQl
EQvURQj5arvpydCFrRuhIkNSlwamF0dHxU0dCY0nNhDctJtEh+wi12sMlbT8W0/PCniqY60mPoks
zOR17FvRhH9OJaNbOZRKWjpazcieTYhmFssO5nDLdd8eemqcxiAJhn6yQeC4FO2twWyEO4vWRfDU
O05powkpSUtYEVxEesS+al8fQkwXaJ29n39u7FB0EN4YefxjLaLkNVGbnooND20EKmk0DaQSFq/i
VE/Rn82iH+uMGRSjb2B9KewcuerSsLw2br2VP/0iTljkuDPD7XNinxeYOZkwM9BAQjS7C5fWyER1
v49K3yzW5DZ9lO8lzrvFt/RNmU/Is1HHzFQhZwah3MhU1973pjdC4iQUsftD31dAokRyVto/+yuI
3fsJdnle3anZEMw5urisDzqgbsu98C7w3nbxy7RcQXguNvUy0wuleBZOWWGyIDf0FNHDdZM5ZvQQ
Bonajoop2uhkxLyf8MxTarhogU2RB89IRdg54jkW9z141OiuNKEjXDPdB6h0KNV4Yo3RNIVddB6c
dDGYM+SNZpZmfZ7+oQ01MfeWYML+iTZFxY0A3mu2mwAETm4c7Po0tqRRNLTmIDF61JHTgo2ADkf3
jBwwodZ1d8HljMXbKs948ODMzy0qDhGgKCPIcI/mKDCrF+VvH6T9zWk/I3y2MDy71BRE4TnwzuL2
Dx+loPdQq7JhqAdlQ9pwog8e/fuAjBBuGLHvHFhJI+hr/bxmPaXDnlZoo4AT59kKOOxycpHQFlfJ
Rv//qKDJLy1F1bptSrJkeScLBp7Y87ntQA3xYMrMcHk8j5PUc0mUX6XLpbv2TKE5xqAIgdEHxJ6P
j5VkkeEyhmsEVyO1YoXyYOABR0i7wUNzh6V+QVY25gGAmOe6ObidOz8RYzWYAFW6FI/qEPzTpmDI
5j/lbKBuDkH3vb3LxsdwSwk4ga3kzvhxXVTiSEGKx53wwO15k4sytdgaEDZXS6EAquxXHkTzEx0W
TRy9jXB3pe2UwVIRV/sYl+TYloKCJwVyixoCQ6o6b/Fd716+3uwfFLGT0N+GKQ31lohAhd32UxrV
BlW6abgM04oZRa6KqxR/UjZ3GMnNBsnewPpocguIQ/18tFM0KsHMR98YvJEAfo/5i/UpQPwbTZ3R
nGFnq8hfDFMGkm++XntMwoEmOIBVQXkEFbyDgWrn0w9OgLn8Oq8uM4FXm3lbF8QoJyiGTI/duH3p
WdGwq/HeeHxEfJ1aDwnnoA0XItHdUeLttK+kRcew4jHovEpOB5aTsWIUNQVCNNWI7yxINvWGkjtD
HtxlcFH7RcYg2DWyHc8epVGa27rt+B9RvJw5Wkt+3dFhLkjTeNnFGT3VtOY6OYxrRrBGiJLe/bIT
ZWMN5xJ1EUr5rz3rKoG8pFYLNWEosVYppetsgnEvqPQI7uC4ezIqBLY0/pwZ56RhmwpM+cZL2Zxu
BPDUYsQ1IZ7PbokyRlXLKlkHyRUQ4aASoYuGMwWdGia+m5p7t2S2w2P2R2OLYt6ZNrSVrqN8woj7
/GoQ4GkMpzm/IDdXLAU5EH7H+LjtDDswFBl5MYW0ja8WHYjrYJq2/NImxDiqdh7CkP8wic5pKfQz
UG4No+kHxpiqtvSxG8Q0tieupbB0upwFy+zsG3tAFdzOklPj7zIC/3xNoRNJs0itXYap5eqs7u9z
uIZhZlo/ngbfy0/SuoRFaPTZj5Mgf+mMxWQ7j8Kh7PsN7eHFyvhhT/am5s4u2XdGSi+aUIFJYXn4
BKcTuhEg8VlokMmDwCTqlzcASpvdzoyM7aEzfMssFTySqD85VDzMZ6UTh66qx9+4rbClcN2Xndev
LSK5eh36JfD2q98/s/uf59AfDnLrg5EOl0MtPm2OaCckXyQVFYp7RqKxZZ5dTxGevwsrE9tRfcZk
DmncVNlZ/uw3WVcI7ohhFDErxKlIOb9qdcjh56higuXzON8XE1gshNpndW5BDRCedWxk2YRpoiOs
aUCWlJDx2bB9/O7wUBOVFPwk5Gi5A2xLhII7yfMVVYiaOQnKM2XQsnNZ7moK5N+XjnkamXP3sj1U
tEDLD4AYmdf9cTCfb6wcyBEEpr/b+OUfrApGqAxd/1Nczz3+Ta4dwEnTj94DRVzbl5iAQJ4ZUYuU
17+VRYj+l49o9PfPzLg9S95XDdTUdZ6e3aRj2656xwFAO7/aW2Fhz/xceeOh8ODy+N+X3ccwfNs0
JtzFCgrHCp4KAaxsVaEF2BETpiBSK93Fywiqs6vuw9cd5Raw73S3mUuRyB9invdkSEfuYSybCSDU
xZkkjahb2xRMKjQKaESYZ7sxSJJuHaZHzW0K+zL+0IFQ2HBocpXeh5SpNgCm79SuJPEOdmtzmN3D
0PIUlIvBXdwE5DSp7g4+k+y2WNRlzTzp4DrFGWfVYAQ4NPl/aru1l4DVF9xGG4kGgR/u4Ha0dkLT
J6mJE36SSs8HknshuMKpN+Jev6b8TluJ+h4V5xy2S/Z0P4Rf5pwBxwSBpcV+Gwo5QQGuVP3oChQq
2pc35PFJnKCCzBs+RBnIYeq6xmmu9pk08xQAe+o8AJNE/3cNu6lW/shi+rCttfjSSQXSwzFY6L3V
zZsrNQKzGFbG0HWPmoH1xOuLrXrNfXy9dJUm1nSsy1LRYaG2H3/IchBGXis75DAx5cdi3ZRMxRlH
UCMmjjbCl0883ymBtd60nLs3x2VL+jKtpGjlGPSZPvworT9FeoSF4EncTS/hg1Ncs25roKNW7Vge
gKCCqtg+PHXnYn6NLkBj8HvTKYOctRyK3HN/7Ku8SwdNydHSjsZcYmwb83ZHCzDoavIc24/q1oww
Nu1K4WlFrehYI/3DYEubJFXaOs1xm4iSux0Pe1ofDepHSf4QcDm0YfbIKg4eb0boT9HfFbFQ9Miw
WAPAXJ2yBelJoV1iXt4b5FU38jleLUKgP7UaCZ/8UWIim11HvLArNHeYfmx+5twn7yYmixuBcrtR
peo1kNUKJGzK9E/uGsqyzyCHCw8kSQTW5rX8oMNVryZ+PgKWz+0l4M4UInHaPeBHCuA91LclFzi+
rL+yLEvYO6NC2xKqBEr0OqYkqT7DE4qbp+2Yy1iBt/ZBZ1eRklaFM9aRjMmtQKf5eCR6MxOz1z4h
sJwbgJQ7r3myM9nQKjHyrgLiqAi6boIePVP0iZ3IrU3p2WON1tnVnfzUkcsIX9F1r0RV4op2cXoR
kXRpF9+XykzdwTqAD18lVgpaZZzFr6E9D2teqOz0AaYy4QwDzfnyBeXYyiFI9n0R8MoIQ+k+aYkv
YpkdMHjLqbs3GcsTzZFsK7DR7aDhqSwn9yZ8I2Ov1HDKu2Hv3KutH7VE9MqT1lrU/P6MeBUDqX3L
Gg2pK3t3Eh0mRVkYfNM6OAVYUTes2TBGNlqk41DdXmeFHQ7yLwYJYZfgXdL3gqn7ruw0YDo07Aib
XUKl9Sf1WzlobGjCytnoyHFwx10EXXk/0wnbXzaEauZROozXp0/CVaAMVcw1W8VW74qMxFBQO3An
ND4Uzum2HUMji+eHxk08K56Su0jtL2CvXuu0frdN4zaobdTEzoERLWJNIAfflcup7sYMsMkGQhBw
hCzMLeMJaJWqaPxNCKX3gBiyCjV8VGNfrITvMZpSN1vIc2er5oHPA5bfCMBsoelKM2ckry3y0OXv
RRGDTum/2KG4TV05xFljRb2BL5aiQLzmu/wqLzfIn6S+OYX5VX/eZdQCfP7SstrJ/zTeU7prZ8H1
svS4WqD7G0pZUO3ayUjyPRPJxBm+X6OpeRqLmWCBtvw4niwlqjqwBSfQGZLDFSNc9H2iZM6n0E4+
BLFNlkcBgBid1xedjO59LW7pf41mMe/nB4YwTC/6eTw3/n24VGVm2t+dorBt83RLe27v82Dzfk/X
tUwhiCPmyzxygbTAB/VCSVx6hRsGFgt3Pspd7fzoykX6ex66rVfVt5ukKPJKpwF7ZAueBeSGWZ1l
BFg60gZZP96gHCmGdlNQtMJwx7z3XTF423uCm7fZ9O2o+57q483IXYKDbotn8p+rTt47DniviSap
zoSgJuBC+vg1XtOD6lPt8Ee2ojGkPp7dTUfnUqFcd83sNhtIOGPTVwo3/PIwoOT+oKHrAmTbkvEP
gQMcDcsGF1nUrLcmjWyXclRVGj1v7awP9Lqt0idjnHRPh5I5kvohtT7RRyXReDOwgRggIXe/ufJN
E+4xmLCL1nbJ0Ikp9mCgBxRSNDl0+ZlhWK2R+VR0lnNCX8+lZoiDX4Y5Wy3l140LQR8hN/G4/r0d
GVfzdlO7ifIQiiWIlH7OIAgdHB922n2FES5JcLbiX/N+MGYFzdwh2bz3aRTRBQZREpsnX+2O79FL
QFAHbWFZBUV3RahBfxZvSIZ3MpJnCmo0eHyUgRbfkFwC4WJckSt4D8FwIti2G862eTEJbU87Vyt6
X8GBGp/ViugXIPnstFEknQh7JIqXMPNz3zfzvfuULZPQAuUylv3JqDl6JZeFxJC6L+K4ajFgQq2u
fhV05CDDGta7/eJhfte3i6chLsDnyJ4cG2mCDpa73tQFl0dSRi4/5Ag79VdtJw20httcRwPaX+ar
E+wB6gM5KU8E6qqXB2qviQ6EmYdXYsXzxqZDwEvvwgMlawv5w/PkhJ6pOHfnVjWhoRl7J9GIyBSv
0hET0t4Ozpqil1wqG0X5iGuDCiiwJvNyH6qe4H7asbpQcofFmlDDzX+XuGQnktlhpNf5s8yDb8gp
Lcof2e9Bk4uTcFrN7j9I3Fz2iFWK0dQLHbN3bGmTO1cSvivTJbH7lT73Xc9UtAxsxNMAfAar04/G
0sXkEHAcfCHXawgBKno/ouuboHu2dG49VD1dhXlJ/NL4HkAL+mM8SkMLbOvDEu7CfxMg8PqjcdnW
b3rhNQYYtRS3DhuGDNlLFRK6SxYecFVoVkqzeFkefiO2JCE27ihdP6cSoo7HoiHu5MPh+XT9oG5X
rkiFGSQGYKtJICDZ4XMO4TEzk2gBZJgh/2Dt114bVEtg82ZuMacVRUrWIXfrbgV55WzibcTK26rd
cmB++sZwrhVnCV/jXkC4UNE9RN2DR4QZ5KOxCGPdUkTjtChACK+Pam+iH42WyyDKsXm//cR6LeN3
rf5q//koSOZGv2JZPRBFA8GSaKlOvPIDADFEvBatHFIa99P61NNeIl14176va3B3djVrOCVZnPD2
xq1NXRqfq18EpJPkVvJoG55IISzNuPCkCmtso4NXIXRXgXXRLIIZQoc1dwQxXA2xXypn62JYYlhj
hY9VM1YzdclCGhvsgexW60yXHuEWxnm8sjygsgTR316s88HcL8lQ7pie094KaeqIcUkeoyXVJjW3
uAycMUbaYuxOWnYP7eeMkQHM+E3DBLsmIjhEDiY2WddaWrek3aukC3bdY38gkv4jfrl1VYh9N1Zn
Aqkum/qPdKIfRZI4U2qESPOkP8zwdCAkT7e7a1ijND4IfIS/5jYayakJZA70UoreqWmnqWiM6aiw
d+4Gs5TCYdcFOcgsxG7LRr0vWxxWhvmp9KLSGQG4OTrkBGa3j5Dstn6IgW/IKtKXyDhoJlY4zf2m
UfI+zV3WE0Wr4HN/0d5HheUduCssLTZ+QpqSmJU+jevyXW2+DivDguDIanplsXHPwKZe8ma6y3PZ
2VYFRij0HAlvfbPBVwXwM+cUKnrcNlTYq0O8k7UGmJVVw8WvGT9pRJLcPs/94WcSAuKSgKc8Z7MX
F+uFygjToB0vv0sLEY8bIu1GwPCPupM5h0aqjl4USJTYLHlePMs34KTYQOeRd3iWdvj+ye5OJEsq
7DfdWwt9dpj68YALYBy3hOUwekyvbBd0UX26IclpD8teZp/PAf5WK2UFrZMDzsmhOf9MjcJZ63J9
1J6r1zxLZ4OyZGfQWpGh8iIiT5vrbYTl9/Mw5Ui2MSxiA2kSSZYPEChhXyn7jXDU6sSp5gJUe+ZO
im53CkBOIVFa/CUxSmyUdXe7ZUVFukE+Sv1bGF/5pDLMWwHBZGlIikkIXGjdbn1rcCBFgBqPbZGe
42rE9nhqFgF3p5r8lAcO1QSVZTM+F58fIsg/dCL7/M3d5xE8ebdu+YcTfoXftuP2HMAEmi9EJR61
HkdxvQezm8LvsUn63rjhtGWMr+xUpXgBhe6DZlBALAP/kBpvWW9vdiXG5NFHtSTohNp8qluWj2Zv
voVKvRh07uortgLSE+nks9lGxAgF0TA9TLUEwnxe/DMQ4KPctesKK6nO5FoK32H7dxfzALV7GVHv
9yAVXJC8zLcdkVAkaJk9os+TaPhDo5d6DehvRkFDqA62mr/mWjzUi2h0fbG+clXxYsyWhSqPzVBE
oi7y9egeiRk/ELSRlsA+S9hIokj9pOLwolx473rWCcQXKJMzlRGwoLfKa6c6BlofOQKdP4d5Wfj2
9c1i5n3FwTK1Bom+44YASZzQjZhJqpmCvOLVZp+tD3cjsJ+XKARVNRbAhSQ/YxuXQ7kmMTRBgJJT
CLj2s00TF0lQTB8r6+Sr6cu/vpxQW0ivScCS7VOT3EDPi5kKDScA0gmXrikDwGgMsCNTqnAgqB00
OGrEfZjn2dX+d/YT2t3WiNzw0maPzEs1e7M5Ej3OTkgP0f22W/oGOab1IbhA+Xp8WHPcarQVuPFM
vP8E5bWez0hbpNq07z2+/eytnWgO3gBllEYkC2XInXsI0YcnKxi0FaqYrs0OFDO1hY3L4naw4m2f
W1+ra3xyf8WMOJtLtHIQigQ0/KjSons5p0J3Gb7ZF5Kma3Bf832Jkq/oQQSDRH9UScUe3GizwKF0
dEekXJ6HSp1JrRJaJickUBlWnN9n40ggpDq/v18Pa03wTSbRAjf+qDcotuh+DspKaxNb6imvmV42
DoI6C5s7+0oez+xzJPYV7qUzYY6hQf7arEI9jMnzHIivOz6gTb7YxJQ+BIMVSHYredIJjklj9vZX
wfVRCt5yDh4vgQ/WlOz0sskva6jETx6e9XkGQ17keAvUho8i7EbTGITu4MWP8dXyUkuNu8GU+s5D
i5JyrRSTEk6sX6f+mNrFrLv21kes61+kqd45rS0SVu685QOc6yXqPRY/vYmsgrFgEdKeblg634nE
Gn8aXmXkt7W1vTfEoKM+3wVXAMY2U2Y8ESXKG+DhSpPri+WK+8Nfu/YGBygk0XW5irf0mniN8zmo
HqEJHBmWyACxgFgn0T+aAJX7CE0lVbdgne87EL+W55oL7rQy2AgGJvhGR9lj3yaKq9Z6H8uh+ACs
4Q+XM4Aj9NN2eajjWYBg60VmwK9165m9vNQrrTR0+yrmnaZnZCfNTm0I3nfqOZzKqSqrwwzG9cCc
HA5Nrhib4vNgpsrzKxj3dGUGUPYh1uv6Fr0Rik9PnW5wePKm9nfL9ZF343gRv5QoGRmjNlSE9jrr
lxCgxcCnVgedExu2TERnN+BDcHOpNjGRaBdlJVR0jx9rlwRt8RLLNe/YQTT4u+QeGVMxzkuITXLW
parIrq0p5P5Cn5bVfFjGrgF+z1qp9Z3m+oaTEWHTZ92ExJzRAvSmbXYcjR+OfC4eAs3D3INW1YKC
iK83GZcOVBC6UjAvWWGX7aosF4b2CwKL59q7IxI0s3mW2QcBDLrexbtjYj5SA+uroqNlBMA17SJ5
iDB6fyZthS4FRuhzE8vQQwaOlrgBiJnsDX4K85oFiQVLDGhK0DIaAlnICHl91P5ab3GqZR7OJCaM
ty/YoCi7t2af7A11AHk6uh5cc74ibYHgbq1/7Tvt9kHFohc7SE9/4lIpx2e2c0oOVFYsL3zPckgZ
H3bcyS3WA9Y8v3NSdkvVj0L0NBVRabaVHMOXX/f2rUD/MRwaLKtc2KD4nygHCYqdOsB6zZOga2zN
RxDQz96AIonzeCyzH0j/xqCOBueOkaHMJ23GtDFBCKRdaSNoAot0dGtFYib1Syg/nHDPffBQN/BQ
ifEFkyvKM8dX87jTiyYWg3f3tUcBm8Yhrzyx7rrKTWJSzEcTWANjmxp+GKSyjJozyvwA09eyW/l1
+gBmG66SSB5HJ7/LjIR9saeY7AiidlJ+yPM40+RpWvyQOS1Lav6V4/BHAtEarGKtCHwCyqqTgI8B
SQDp1cADF6WlJlmI8m0IIlB/ps2b+2HqMO+x1d0SQ1HtQpef2R4kTs5M8dHZr90XauXbjGpIpotU
P1jdhbzyvQ6J4cLPetawzvPIvw2H0c7xlWVPZ4FAp1k75ppU5XZkCW34ML/bDAX/xWL7DcMUx2mh
BKWV3W2dN+JjY7tJdaFfzUzAXVdnUiB+UWSnrQt1PlivVE5rEiRidtepb9ubcKBTy6uBqlt5KyIQ
nx3F9xZPN+d8uYHuTJT/4dEm7z3S1Gv9lTAcl5JS7IS+AmlNAdhxMwGGDiEm768Y8k/jyjCTHYuG
2otKGOyMVrUe7mu6voDVkVq9XgQ18Buwic4MfbO1B0cHUZOI9B7jCMFxQxzWpR/xlSRXnqhFSFJf
lmEoDLnNZzx4qvANGmGqBnlvUIEAVuipOVJb4boj61WjYegjO4UX0UZuQZEzBV3AHJJJnNkqAxgK
+c7tpnVOjeNMvX4xciuaBhnWnJ+JzQAZx8pDLSsk8JZ4wpHlZLJztIzIZUbqwDoRU20eq+vrN1GQ
xsytjCqomCVFqgUzH2OPc1OgviODchmOXcztJOrFDYy/jD6+sECoKNVorOMoHfq6jfUPb3bZoivs
HP9zoemFNY7q86rSQHQbLuR34bND06Fdo4FdrOGzemq3ZuNYQl9DzmS0LpTRlyMYSd/5tGZOovJ4
5DyDZcZgni+EEDMLin4XMFZvVyqbL2tyBhzHnrSAkwAw6iGaWhKjmwJltabwfkjR0zPAjviEdJIN
+ZUHR4Wea0dU6uX9mi0eIryVnj1srGg/UTUE4tyxaH6bXS0HIKWDfrJIQkGjR+5g8RlrIaLipyc0
1QBLRFl17FLAkpVSFjKww7ivZH2jsjx+WOUzITtWg3lxBZruSdpWwYH9w80aBRHDOLUsQJPS5H1o
wjxxorYbIDh+NmS+eBv0gafAqv1PfwmNYhGNuljM2gnNgN8DghYDRzIPhe6/f+irsKLLw2Xb6BMv
MxWZhLvEvaqsS4SU9x+QweOgzbDuMX9GOXVdbloB+QoG7p7RwVwtqUvYQEZ7xXco5fbvsm1aKBs8
Yl7bXCm7dtL8zjfkRPk4f8h7TGnaH9sH9kC0x5e5K//ci9yn2tx52kmwt9D2UC9GFIAyaX632KeV
WFS6he14qq1HjzXQColMppT7S/sljJtGngKqcc86y5T8BfhkTnX7cxwRFL9wlHhdE4lnUwgtbQ2P
IGua21Qw66W2hOPJykV96fSjapOLc4fdxgqeTxPJRDW8HjralZE7JdfEq/qNHDN8YVVNVzN/nBag
7ol3ufqfECr//aSyDmqyZYzc/L7p76ZDmdeZCo01N9poXW29Zh7Okahx2T8JFI6h3841prmeWO6x
T/hdVTLSaSyFwoFd8NSXz07p3XUfNzWReUIwCqXgvuJpeHyz9rTQCjeHJF5nCZ0+R2tXHYAmaQLC
sQuMnx0Tpb+v/lwSrg/x03wFoqHnPNQqFZo0vJLGCm+qu9kjwgva/6mBTUVSjuffxQojbGfFqlUn
//WwlmCBAmjoEyguSpi/1KtLZKdHBKYQnJemjaqF4ROXFzrnffRGjRdGnAEj+2PRxardzxu9akCN
e36GueD5jmFjnYid5r4ed5mTcYVmNdssJsuEjRUlXQlWecVYXPMnyntDCknjABw7uNrb+sVMBvrv
CyiHmAsA038oTGNvQIDPltFU9cn7pRIHxauge/I1Ki9fBvaA8qWJcwKiEJeOeQrZRhvq1W7AJP5G
JxrsJcDYKCHafvuByUtyNlR4884CyrPS5sCes+KTdkIOV+jiqNjWq9ji8B2dc8JtUk7vVKICfrt5
NspckHEXuYT8JXgjIqpyj1W8h60kjcwpOg2J4tdd7BR7v7kYozy2W5OLcB24/FWLJjyx/vQ6mdGO
EY4Q4BujZuMx2pS22v6cV9YPmOUz4HebTvjyl7/v9o3gwlNpMY2Xqm34smQivS5vdA0G5d4kfEvD
+D+1ref/CZr9P1c6swPC+KJMmur1298UkLWn/ZQBXJlC5KcT2FIGM6fRr+sO0mAncHBhvGkyliyb
vHv/otSV6EG8mlatISQ7uNVq22G1eXUSw6RHzLHWUBtiJ7hW4OpZQ5m3aY2sa1kjBTIJTqEIAii4
mAeYbLoeGNyZri7b1pqm93Oal9k5VprzsFTfU5UDEQfy01c9QKrNcyCBp0MEHaBRQnKgW/e5giCM
jzYRIEmDr0qwZZu61Jhtk+varnWG/8EqqAdu/Hq3UMxcDFxuEhua3RiCJNj0U3a8LL/UOpayjbCF
o3hIGa71RnIZSD9y2W71f2xRH2h61An+PQ6DA1fTqxMq13F1eYL92c/skkTPLFg69uGo/pEcKNIi
awP9g61x4V7oC3oB1MLeP629EcS+lYsDPzd3a6hXJ13L5mNhu0dOFv5ZbW7KHe13H2V+VA16zmFr
HRklIbHN+uRE1PlX/xv+LCka7CvWxCfzH9hj0vdmORgz6W879eUkBbPGs0jewMgOfjOfjssCkxj3
d2nMUNFJkR35H/KheAkGGmbRUT0fiLc2H4CTcy1vhsdBBvSQCS+p1RWfb17JZ9uo1JOf0TFN3mKS
FU4xh8pJAdIojviqXMygVFSeJ0kqAD8LvvYQ4oeXfDY/BX9A9YRX1ZMuYajxX92Rtszr2xFDR2E9
xmebFbLBi3O8Lxn2Wpb6paMyc2IYonDUGeBBdSGpVSc65eFn/SVoIkzmJrThK41/DTQlEoMUuO9o
5yfqwyrMvL2WMOFZ+zASOcEAgQvNQu9feH++I5oBfkQhEwM6NVPh8Ic4KX76BUnriPQ+jMwuoBzu
sSgBA/Ls5SV9tZ077dfIVj+BxIhstsbXeYIE9xpOolv11ULIhYvMw7GN9tWw+mxjv1drQ4xxeWt/
Wpz3UMshmqhxn49+WYt3eqWYMHf5ZQrBwzV1+UvIrX8EwSAZwjd2KrRm+gDZuhLOokhzqUYW6RM2
iHHmf0DRMvftqqfRhxN6jCpgbu4fdWx2s9iVwNb2jt5OvPJKTkXFvxw9mNop+GmkDjkgzot/G3Uh
h3nw0IReiAE2TrN//hagYMe4p7jB8EsUk8i0BMNOLffSeBCH2ySdEy28j9dg3YHvSmVth0ZP2f4f
WU/y/C3V05emfBmLS/UqnlEocjuUWd63j2ZMo9PdYhGBPsddRIzuBXE3EORNN6LOVLsZQ6WJM/H3
yZsCzv0PdIEI0h7ipk8bokwZ1Nwj3n3gm/5UfkoGdVhej4qYSSjmDzaWBxIh6IBpY7N8+1zuG6KG
b3ND8Mx9Sf70caCNir4Frt7Px9d1a9T8UCo/rKft8s+x63TwHxAo/sj24Nfl9t2H9KNvXBSqXi/d
EBPjUv9jNosCR9o+N8DYLcY4ezOaxuwbaAYSEtE3CHnRkf9G5lAfXncw+pKBRElV6ou/5Bd05K5d
SZ/W24k+o2jzO/F9r5925GqyMwj8jL+vd384GTuiPWF+zInf7qvbn6QxofMALoOqy28YmCpkCpvK
G+akeasnQKjip3og80+ayBf0O3RxDOmLRVi9PokEtAMFYP6zG994YtdBcofHghSnHZLHwEgkA+BS
R1t+zwwTeu0p7yu/OZLvN1IlEBCLoaXTB7HpP9l7M3rq4PgmNnDAVZR2F0RvwzZlTQs9g0kp9AQu
yLBNCTH46+Ydf575yC4VcwqirGSbb4GhfBCP2dy08bSJSZonlE5/tafNn+gOHXDq/O8NThB5d1Zm
6zmrKI9yclOTGcHENN3FBpYqC0UHNDhP/zIzUCKOfvAFCMRvfK0yDdcmdPZsHM0K4lrOM2tDsNUr
myJ5Fw4HWZFiN+st1hgPqeIpzpgJpshQQe26BGMgJVx7VbfRRYAHLhi7c705lEFKdq+lCTnLWDSi
cUm256C+RaQwRYp5MS8XeoO2vP3u7OnT0c1oRldkON4FnSWcuTlH0rvnqH5EP+6M9y/t34jrkq6q
aTVg4eknds4HvLeNEqQgM4z0uDif9rcV7+jyETWay0bflcvxkbTzq/6GVS40cXTngsq3bEbYp24g
SXkSwl3YUg/udAORHEc9Ltj3SU6kZth/kE2cIU9a6L25LfeOnEykYJVk9er1krkpIjYwzFsJ+7Nn
59Acf+cGSWm5wQjIBiGDqcojB60ekIfSp8FBXwl88ewYuBDZkAU0eGG6L2bCKT3zII73F/iJk4mn
Y/zKr95a3gfeDodYn/oYKhSxbqs/38Jp8gVhHsuARR0pwBSdkXup7SvxXqNA6pwc95z1+efwe0Qq
7YRmfJMD/wpESABec2eFpAzYmN2mDWnKwSa66vJK0PK06/FPWQMb60W2CbEeBFRHLka60Tzp0xVl
vrDxZx7P7B/pcJhtGixpoSqDEXgh6EOim17lJ7ft3YaJeETxSlFStNPDsI+fw3P3JTWWx4oTWc87
Tl6DYRMaeyPfRmfrC99A7GBte0fCovsgf79rcJdAVHHc3GcbIzUgKoUI0W2sJzTA3cUaC96vewcL
v3GWAkc5cc6iqd86OK6dVLW3vP4pHwEh7SV6buJdLozjcVMFtwcmCowtSH/bEPurL4qWzuZmPfev
GTfgdu80WRjvRZgiSgwvpIjkLQYMPfenP4CO+lm/e3MWVdFQXkVKcLui6yny5TQuBm/YnUWCk9VW
85lz1lIAvVkZKMb8zNFYvrEUEcpKr2H4NghGXMBFqVltByumvXBht85558RP5IJNCVxG0U5eCWND
QULLaoTK/BtWzlTd3lURN127CO7MNL6+MdYtieeJUTzCoTXelKr8BmhHj7fwXdea4OmS/gbadgD1
UuQ7nMqc+CVgKbEIRgvESXAJaAh66kowapFUZ/cHQ8F73bF4E7t6zlFXTMhHGnPXBqlC9pbO67wy
9L2WN/Vdf/xHzVjW49Vno26Z1suopW3+9gWLIfCUadDVJubKsUwPGF/NzuNHSt1k5OTU0T98M7Aq
4fNorqcx4GOGSxa8zVjrOjSdoxPLEXWLlXc4Jr3CJFbXll+6mqUa+YZXbv8Jn9sOydyJutwWRHf1
TnAdHUF+fTL4NwRd0bK61CY7YocWzKcmU2B8ZHAKLR0ueOwWb2zIyhQ4UTYxRlquhzOA7XGXhoIo
OTTcP4VVqviH3aVIRE5EtFX/3OOozaz89jxNzi44UzydgJgcX9NuUQk/cdvDLX+XJCiFUG5Ybr75
53S81sj5qk9ZC1VHwP6EiceFIlmd2Jd0qVY3zKXsVjXGKabltOMmsa4UAE0ugjVbc/Ug3b6v6BSz
m7XZ8hhR0vZHXPiTNKH6YmqnyFpTxuUahJ5Ezhy75TpjApFZF4jIcR8yiE243XTDifyw21XHxHvu
5v+t+EeQ/g8lZN4lp0uhKrs9UparPJbZPjGBS1foFwYr53DS1BWXRnFwLwqzq9MmpGFuyNphTBux
S/xhhS5JaX5iPKiYPvSHwvxJODbtbiLQqJkM3irKFiz2ZfzxG/ES7ow5G8U5Hc5CAcfySkxtBwl8
+y4jadui35NBfoJujqj8/xdjTASGkmSSPrbhG4jP2mYD7CPyAtJyCLelE1EUMLlYkVcF2QMhPDPl
CdRKGH4RJaQUlfsypEWKH6DwzZuvxeZS3pVyFpPgBi6XFQXVynlAplbhDyqRzP8ivggcwNOHGaBj
VxRTKt/W0IS4yAKvAnOFXy49wWzhDUDrQFjpXeSzG/ZkhSH8Kn3JHxPFlSKFs6VOzhopaEhq4l/K
kvGxHnsQKZLD9qKhz1zrWdMOCL8OK3eKgn2PWVsydhko338607chJ7nbx+EpLWAUo3g5xywQLiD3
VwEYV5C8wnZlzjTR1QRRyVDZ6QeyqyEtCTWx4+xKcZKo/09DYJqelnnf/n8CqjqKscC6JAPWrpmW
UhbPMgdzgZd3yAmXrsQ3FuU6G6GK19XSlYaHH/HIavbKDFWMkhVDbdesQ98cTBOIEmzpYnUgTPZ8
2AmW1dN+TqVjkO/+Bq0GCK+h9t9qoPpbqvDK6bpTUDszvwPHafN1O8gOeQvMtG1JXra+9UkfJrxQ
VuWjOke1/ssAFc9P
`pragma protect end_protected
