// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
RBhMTLtTE7aiL9Xrlt6RWqnFnkdFJEEeRhiGmdolTrqtlFz0gvllbMMgC1ZL
JdvbktdLnXf84O7Q9/ZwkfdyTaLANFHAiqQvO66GRDTyXJUqL8ZlLfFwAHyu
/6PdBsGVFge5tRAxFRNfEYDunVryK1qPA8Wlq0/HKzFh+s3zTRS/VgTf6sRZ
L2O+4g+6AqEQS8VsRLoJEoqWEx49lzO06Ukb5zOuV1bomuovWz3r4S0Nn54k
xck4H1GhsOMSxHW0Q13fIRSkm2tZb4FENN5NXpokAYPgOz7QrFmvu/YLzlSP
CUNQS5D8DKCIupd6W0ARlpN2gev+JMrWITtEYOj+BQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
QQ9eAYAV5LqCDhjeDQCftLRTA163n47fdbhcdfOf5cWLddEMuLpeVLjpyfav
ycyVoAtj2g7mhid4B6gQdc1PY/WoEX2nHjiwNM6aZxc9H34Ur6gaz9L4uXHF
pdpFMNIhJGbrnB2lTi69iPyp3I7nzxtGw8xqFm56Kl6PPaQg9t6WVDZdZoK3
P00TZiBt653OCFd2VjsP6t9zYdfFRp/35omTtMJETogwL2XxJQ1S1bkFKdNU
KvNBAdFa/PbPA0HUfAFLcYC4KbHxbLuTypkMIXeZEOYggrWjcx0k81B9YmON
3Om5O0i2MeBORsTeIiFuQ5LZpe1vDG/zpDhP+QFIzw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Ah9Nht0/8b16FAjuaipBJ67xSbZ8jrF98w2MiOyvIPPIQRF+MOoUHpa+PC4q
fa2G+L3Jc4QAjbJq4dnG3lredM1j845kHgcbMS5f/LSAYV7G8Z80oegc31cH
eoA3YmsGaLsuOtxNEDRbzPokPLDXQolm3oL/ShElDWNKuseek+zHlxbgwh7/
UpUotdZCAo2chdjrEcnsm6rtPLkTXBN/M+lUqx78UuKCgPrllmzcBve/+XX7
KfCjFSdqhgFFV7KNMilBZuj+qoQLRoH4G2fRWgbYCbAe123R6bTtivusPasG
e6TuGfNs8yCFROGWaKncIeL4uPeMTKcNyqm5iMzylA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
MTIhpQyWEpzn9wXZKtdOQUC12hhU/FiokhXKQxYZoi4EkSOBm0H6Vp3wC+Fj
92PKj/VgTBEW95pGoJ08NidWGpfXV5B3Hr2Ea0aKadCpVlCy6z2wHyOOMCOv
I7o2sHhz2wkApA5nojpBOYNaXf/ujxmHY2Dt2bAsfpNLZakUaEQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
dLnlQC7tHX81bkzx6gaSgX5AZOdt+x1riSGOxZrNOJH+z5xOl0BR1d38pvBS
DEJB2MfTdr8kkUnqN5o9UYUuN2qANgwvNLDq/KBUGOQSuwqg7Y4yneBC8xFI
Gd6mVz5deDrKIgK7K+Rz7mO7qpBOC4MHu9oln6BK90uq8LU/wSbegGOBoHiE
lYMe/YgVsHNyCYXoGNZDpjr73ppy5st4OmJ3oVIqr9omrQHSH0tphljzJjep
B7e6q8t30JCMyGmVtK5rOAUwBFCc/zV3fWTUvodgdTPRj4pZ5SRPYmtEM/sK
4EC2KmbIz5tKg2ZGZRDdPaNcHCUp3SLRRnjpUYijubBVbEeLoEXe6xyTgYW8
Kq6IjXVYK1xn0Bpd+1pZFBfU1Gt7pjLpaLkGbhozSrxRZEjsDXlPFinmfmid
hEpUzHO5T3+V00ll/GpftP0hBZUAT2iqmd2pw4UZ9q3UZHgln6yx/UGctI3U
5N5jfUnSJCkwtdahEgD1u1iTf2forvkd


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Ehau5UdZJJAm8Yh1RNSCCQuCiHBeKhOI3jFhuE5x0S2gkulw5fEbVMBW0S++
cY97Mllik7tKoqV/uod0FMLw0ZUaHBw4Y6SijTTLntmncpUPIKJJHuvZrbAg
VCv8VXvfWpTuTvt+SUSxlaJAQTkNswbrsEdr1bCVFVtnp3zlcEM=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Zv0tBQOP2NjWFszH9pPKEeS28NsbgZDbt1tLgaQg1qz1Y9x/fPSe6Up+KYiX
xttGzy3oTwxRI2HYicqKmKfu73VaP0kwtkEUHOGD1QwS08sPZLplYpZJGAzj
kXqPs6neA9mlPy9pGkdjTNsTgTFoLWvcKGlQVAJKH+/qrLBmiwY=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 71360)
`pragma protect data_block
Wfsh4AAy+lfo7iaZ7E97GJ2Na9vxeX91qm+6axwfAJ84f3ugg9CKFn6SKao1
E/tYpELiYD27lckMqdNQIhszBZWT/s6nniv3raBbmqGChijF/ZWEaLBZmC5F
plSF5FIrMfeN0DsV7U5xYctMBm4u47tQ+kbWPAgTYnw0D7LgnXZknGP9Es9m
RZDTsB0Lmqy2O4r82g0s8M+9FTWAQWlLPrN/pTqrGIYXsjFbRY6QoCuNRNFt
LvRj0+SLcW9VQ3pFx03Jpc9h/7mRWfs3rQqhG3sk+G5MHqQbtaMOYfRQbi3t
wWrmKezWvOwFVMNz90I4V8RAdaPO0PmrNpCWOSRWldUAz8oDWCazHOcEokRl
9riOHX16wVcN/4TiB/REkFD6q5cR7knrKQb8aJ3xU/h02cQ2PM5uwOzePK3h
dYHMdSTQute+aiVixqRROED1n/kP6c9q/HL1kDCnGKi7zjHj7279f7NWVtej
MvWHfzcUA4Kx8fq/pvTu4LKEWtjq8GgvHl0WpdLdrbzPtU49T1834A7JJAIG
GAk4jmqJW0LRNWI3MwHjK3VPvt5knWjXLLxJoQNcLg/w2E3QssjFUWDZTKr4
nK33xooFCKW4UKKtsrLvrcd4GbgFQcdR6Nl61n1StEmkjJ5vfkwHH5PCe5SR
TXU171Zoy4uFk2szQQyEbtyiT8rHOrH2Z+SCUVpxFupWpGW8Au5Ol3euZEAQ
WTk/X0QvXOXUFLD7tjqQGxxBgb/wMyERdefttacw2oqRcJ84c0jFtcmdEdSd
Lq+JExYlO57ujdMB9nWBf1zUex0Dk6m9/NT7ugyXqSxslUiGgLhcuSw2dWJV
5BalcXsu108oklrETsncPJEHH4Ohr0axHUvqVAGXQu2UZo7u9PCCGDQnFTPH
YD6z6LWi36Uh4wApbNqyZ2z0iYbD7QpqnTY8U+EqOVuzy/zzvIxavFeiRtmr
piLlNHaIwtXsLlbds8+YiRY4W9gMlfnrQXaQbqYFftdUKNme6Ml8BS46rjcd
8a/8PT2c62Jo07A7MJHLXpuYhf1My7fMJd7iD4juHdqQupx4wtn5g7aZhbtp
7EkOTNfCDhKCVi40ZkqrgxxTVZlqbmzRTGJIP0gdQm6L4jxOwITyB11gqmKd
R8w6zRluxdUgbEMjknY6O83sbWLkqLI11TJHOT1P7WaZWNaiYN+1Timuo8/4
Uwv5tUXnwetbcgQ1iecOL7ZRH6a3DVcZr3Y5WVs/bRE8LF6d6XQU+C6C1p3n
ci+9cUS3F4ZKHn7gfRzXa8AXCZdT3GxGnOmwep8Go9h311F9fYWsH9JnUNuK
W5IFAkOvQH3KQyxUxFryAlnCguHf+2JWsc0yPlvRa26T1wkKJmEWFOY1Es4T
k2i08kc89pCK+de/sdVQskWFpJKHNbPDt/wdoecvPRSIgh/Q30+5Bqnqoh6J
a18UYHfd/mdhh9KGzU55LT3mjwLwCyLvMD3bd0hbhhjq9YLiCxQ+ktBNrOi0
L0LAOZTu+nNGwUAUHOQHwEySlIzBKV++PqWUIRjDMJgDbiuA0/fAwGnZ72TM
9HoVUhjkbvLfeNLpBLioUmdEAMjSEHSgoHdKxzz46d3eNBlPHaaI4Z3t34xR
XYYzku2H30iPdo3BxkzIriUuUMuN5/So23iBxWS0sJW6iFqYvo2Lcxa665/l
fNVwAC/svxveY5TB4NDROrPgY6WDFgV/nDRHsqIys4Ijkb07VQdVrLPP/O3c
3kVV/c0e2qbi6Zh/8LnvSV2yvKrWRBRKQ3fzR3kvaMw7xbg/NZs9Rj8RwM4F
2A8yTsLzoMDy303Dg0eqSJEiVmpsbdHoHco3yCM/9jnPrJALmQcuYmxlkCRn
rtbWFQN+Q1Qg7XJVE1vbPFi0UeQihl7+PNw6rVNLCVKul9h7gjeldL5N+h7T
ZWEV/MtHQPf7iQmJnoiF0jpQNRn7D32mGyIsmoDFNoliafEdG407eyA9AF7s
LmmxEtJN6G30h3JDJLB6crAYFO7TeQfNbTeLF4gGN3jcFaqAAXcmI0KpaeHl
XT9lhQJ7swtmm0dTQy4HE+YS/ndwmj5/qJTad83DZAF1k8VyI4wHKuySDUKE
xplu8saXLeoS6ot/gK9jJAru3Lf6VoYx+J2a3LujyO0ZJ60xw+dlUJ8zUArZ
WvUZz2mjkvCX0tQH91wWOgN+xCHUWWveXTfdQx0YB1bK8BFLWiOxeKkTZhUE
Ixv1tPCAKKg1pSdzcror9exFDaMXDnEamiLP0X9ode2DaPkMpuc1w/bT1Z5f
KWT8vANr5H+qUZ1ANe1fgVDAwnyyxWO6sTjCogDodV9kAxM+eAz1OS0LELi0
uGXDrpAYibs2ljSewGx/3vvmnTUWuI0Yq2uLJtRJm09RfTjrRDObrkfHQ3Pc
zGxth6jAKJyWwOxcfKhL/1va0SQFfRFtb0eN2lgQ8jCgR+4vjRu5RVTHVr5y
Mt/DBzYJVp0NIek7nH2Oxr0sGefwMNVyB3Kadx7iYJA6ml5QYI5oKRWEjRhz
e5rL9kkCHgpnkDIYjOhmn1tnlp+V6ItjihNcDM2kV/Zm4/reEBfIHOQWEzAx
BRaLcNK0U3p8D938sGIZpupgh0xOhyJcm5ocxrMaIeWRxMwJPLILgMjCXr3c
pNOzEc+qh/FAEFH9M/4sT9V/XH6thJ1NaDMU4Dnu+1VbWr7zUctPN1LUePFP
dEClDW8pTGq0Wul4Gz63Bb9VRsNUwrqx1XqYpMnX8ieIzSS/JlNCRpkB7NX6
mW246zYNIVOfOxivKQ/mXw6PU+ibYYYjMkDNO6YdvoeaGMRB3y2jNCpmlYhL
eju6hvkOhBcodAfrIWmkIZH9Mo8vRqMPNsKE/2O43ZkEyYkRadyDUQrGF4Zw
iIOn3ia1mugssyeT7XGaPyQ2Rs8OtbrmVGk2Q1ug/FPPk0N7ghJBVk0BRPt4
RrAd8vwz2+6V5PNQavziskiYkOSa1Yp2lPeTgwOTU+NHG6g+l20CzU8SzLDc
rQUNfJEf5m53E68i5532Zl5cwlmllxyo9RckzM8SsI8ZQ7qYOI3tjaZ5KyWQ
tBxhNCjoepkNz6T4su+OEeD/QyhkGz86IKlObhSEFpt3kZQ3MrrlEyg8ALxL
zt44+j5OtZK7DWEvy2rICk9kWtosRm2vhHUmGC5S7ZO5/e9VAy31qpthz1AV
Q5S14oSj004GAdIZWhbFcYMu+Zu6qmn0qQ49o4X43Fcg2lPyKzixkfttsHnj
a5o53TSXdK/mruobqTwROnJujdOeHcgTjeysTy6kk3ToJIdQA6zjGD1Anxqi
K5Q8GcFxQjYXBMAsUBm6XSBao8yebs6Ns3D7kTsKf7RmtcmkhSyowMqCmJ+n
cEcNiGV6oJV0kg6e4olXuI6HUYiaKjae4kfNBx1vFyk/c9C7nT6kco4sAUZw
xZcc8IEJdHMpODZptHvskPU7C28RztmRkbdZP4UX9tkEp4iKCjhQui9HfKLD
RoGmQv63bjotPeZJJp+sSHkR6KwPfR9/561A69R+eLCuM9Loq/XcPdA/WIGe
7zWwb+t40vjVtng8dVFxCm2+un1y6fLQHmIsDZ52ggDzlWrqf/C9KZD7n62Q
xjJz8tNGOqSxNdk2bnpRsUje8Ihv8ygDBv6NvAgiVK5a9rr2c0VbQfXXMG2J
7KsRz4VU9+lT1E7tarQ2aOkI+zGanvWH1iHsSqDNfqiYT0uRUdAc//Qa6bG3
wn8sYRMuwPFOOmE1MYqmNU2SiGnsNkflAY/wqT+8RxGyPBAPzj22GbqhM1IH
AnfAcsD3RnfvZuq4tj8sm9K9Vhdy5gOHY2HlgrBfnn+ol9QgbcggKiSWf1Hr
D081Q3iPso4Gp0+dB9/peZFHDNYGPzdzoWffecVTTkHdfS9k76YE7RdhnmMf
1dO6jvhcYiZSuLEEzaA5iag4jbkPVD7WNiD4TjRw/RknA/4mo+uqqamx/po6
IucK8h71xQpq7lx1lPh8F+ialCkunXhDi7JIv3tl8A6EOLu6zsIQTtL8XaRt
Zt/2y+s6VUH1lHzagjaxsLkPm3lmtZ8an8RmIGaV0MCiOLG6LjAF4K3sQ8/5
ph0OtcxwUhNJwzLQ8H2CdlBNOsikgXWUZI1faIm28EBcQfX+Fg8mhamWPp4+
p16MX6S1vYAWh1FfnpVhrlS4U02rnRZm8/F41UZeaq4W8GBH8RntI/Yq2O8f
FeLJ3y1Pv4Gv2RSwBKaGShZZ3Gm86XiLYThMYObSlTDYmodv5lycPy0xfJZF
dW/8QpDk/BnR7erb9yU4lCC8f1d72Jn30WKgYaQTc/cPOZe5nvyatDOzrM0d
T4bkxzct8PApaDRyGzuF5pSZFmoynPlYbft3yQntDXFf5aETKHxJYO1zPCIP
mkN76kq0ZT3V+MU4mZnzUjizRu5BtPrZU7jeggWAdQRndtn88+PM2hWfWuLM
WyOAezbPBrHNe96iQuYE8fJ8RZ81tZwvLWeMvCFW0HMZttTVNpEtZUrVPx0H
B42Oh9SjedEhz1+b2l1zQuYkoyos2wH2D3VQm+kvkgk+ktuL1R5V6KwslT9V
oJ7yNmQoBMXOAodJ8JLl0SgzgNIwaoDOV0TQC3mrJFrcQDXqiHQcc9ZAgWDH
Mx/RzrYcQ74tB5P86NrOlI/+qof1tpcdcko2GCQALr2AyQJ1oXMysuddnuMP
k/9foMizHbk4f0PO5Ty1urCMJNz1ifXdz8qHh9xOwo11sopzLCcIVSqfmLM0
CPWpWTad0uevezWZPyxDe5rgTbRdZUUZkZ+omkZmMZ5PVYsm1ffPCTawek5R
y3Hl52kL/djW+K8RNU19ZuIZsWJxX3hMY1kXUZNdLb+Par4ULVQDMr6wvxIQ
TITuQmVPRHVHSJifvggnK/A13H0pI4GOWU1Z3POftG3xIpaacrAU0zWwLQrp
CJdL/2eHLNvdP/NcefUi+e5fu7fRnNI6oZcBdiJC7XxDMniwnFhN4GWwNqCu
httw14g8IC5ht3NC6afsZx0WqlFYFxEm4WlooUni0M23NnZ8eofayz312ot5
lwvJINUJvLGVv4xvh8x0lnhy80vtsCZ34kQ1CZcXjYggQjlsiYqmTEE3cdYm
i5dvPD7PeGjKYv+JCNTalXZlbRg7VBfvTr/fTPITRTSRDjaFrl8Fspk2CwIQ
EO5Ct/fULcEcEIk80D+bz+lYrpsnH6/C76KGZw2wpm7G7dnQcXH3d3gAmN9f
L4sJglPs4JbPAdgrHUHuCntY1iEkxSXmZWj8/gDDDpXzlzC5YmgWIWOjb1h8
JU0eBl55KZUXma8vUb1Zx/Mbv8dqJX5rwj+L0qXOp4P6bYRuvws42Q8EvPtO
snQKQdrdafyHRuzZd0NzaxVBm5FcJn4iWWPOM9uFlWHtUO2GSeDnSMCwSMvB
eSccrCMHceExtCi/LSEd8dOHjNdAR767FcAwwW629Lv4PsHrbJJ0WZiSONGr
a30nM5kDbjS0+wPRNSOPLuSoW0OLjOH4+oco6r6d/8ijsBD25iblGW69mdnL
WMD21dbhLanMeYIJyJHNvz9BLiUNkufr8gz83R6RV7NNApmD7aSPgugQkuRS
jFiHc3atoqPgXXWrQJxwWqtTbDIQTgvPMUdXG4HvqPvJpxcz+9WOPoCQSo5D
LPkY3waDxhUxmHUuNBJKyKBiNa1J+cD3ncx5QA/RlA0RP2gihuvzQqdyFBJz
IL/jL1OWKCMphwWlNi5VIX8FnPnHKVlw8Jy+Ug37N0mEfApe4RM9fFgtrzS3
NSE8rVGAIh8XGTTVBOn2c2c4Fa/64eCBkjt/bljXsDZpq5f7bgR7of2KKV3/
WBZFRwaxrUs7oqUWzIwJHm67/6Agw7rJ/n7yUGZoFnA4Z7nmCi7pZDkAnXer
U4vt77HKq0C32XFkJKa77TvcZShV1D4DeWHlORJC8r0tW8csBlFYZrRZZ0yG
g3xDR7CPASlMCjCzSpDx/Wy1k1kSAvMNEs6U7/g76VhrYadizrZAm6xeJCgj
0AKXzDLXmpF/Zsl9jpRheC+W6ME6k60ONfzsWqqpBcqadwayaG/c3mA/3Ula
hgXhm6uNZxFD8FxiWEsPJ4fqBh+txZ2gLMvH2v+YsMGBEkbziTOtzHYpNBnA
ePFS9r0/iFxCUjHHYf1PFkEsT31uew8KPufdVWvAlJnq0wsWAyWCLoi11RGP
b7+MbJijmtCZOqViuuTB8K4H49QPhs42nIWOGetXt7lQHTpyp0DDldN1+8Ma
EX2tk18MsQM1kNo7CV+7LXLEJQgdbYcwBLyyRBl+mpEmxe9PkCR1UTT/rX+3
Qo6NA1BtpodmqlxGMGuz5lDZ73rUrWYLGaRIL/9Nssd30E4x9/jhSxCAFAqK
jw685RMtIesjue6gjwETGd7IT8F1vgngqdcGFIMaQYeMptEqt9exLw6FpuqW
LNMxealI/s+H4zyN/9FNuPReXE7DeouLuKEgJwGITs4x9UEgSoGViSeyQ520
iCOEoIUaZGvEb91f4fnQAHWXRgifR0JkqDS+sWF/0SFfgdYYCx7GGnKytBMj
/fLmzFEVki0NhsEzZcJNAzSah9bA46+5dyLrU6TvAMsu3XSCpWwl6Nh/v7Cf
CkNWq5E+GD6CmSNxUvArPTLxxn5xt5JdnT3A3/bxyUuZk96r9qPz1AiIh6nz
diK+u3lAKjNgdhJXpSJoKafJn8yROALHZBSmxA4MB1hMZfMjxg9XMQIeIGny
Drasex+I+OVVAwD0Ow0vMeC9g7CwD9+/GoH8D1gepPbSW6e3v3Ixi8Wyoz4d
yAepBb2PiMcqyOfRwkaBxiXxAhJCXYlBAh7NPBPIkkvV3HA86d2mnDUGspFH
vxnbyLWV8rD63csASgvVOFkjAD8nzYFyn36HMQM27NhgT2//lI8hV5Yw9S+6
l8bePsGDlotLmv3M54Ha6oFEyf3b4TJ9YAHlmYUpvZ2yrmlk6jRSqdlJDcYj
wuYDx8UCgSpvRiq5RYyy+LLmVtmDTc7JjbTbNlwj0u3cpZlSgW11AWg//9XG
WEUbFrxMAkxMdXfRmJJjmewVEygH6MhFNcqjAgJaw2nBcqO1h83N9Kgx7ji1
ewCVliM545d0PvMVmoiPQ0dg7q+D2VK8T7L39o+YjG2MWnftIvxRY3nx+jqW
e1BhsQa4c4Ev90wrhSZTV9qUW2qL5IbT2aY3IOPXPbnHq9Z/pHQ8RTnhWcAM
trLN/L9uKeTIMsJAZyWRX52yJiW3+LW/CtQhVu1AgkUMZ57/eGy3EqjM6rzh
qAAzVouxGnsuldddwkQ72LvGfDlow+z0yC1tQJGesmg+uy+1m5wd4d42XDfY
iZZE04u2Np1AcCPEPByS2EBqYRaI3dDSXnncZdJ2kJX9OnU+O4XQ1lC9b9Ub
H/jaVfcTlnuiPsU5bU/mrrqckt2i9I4Puo6YLsSKwbdlAQmnW8uy5pwXrCCs
r198iI737o6iWCEa7MR2TsEYUkcJECcmrBA4PVesKBHSgi3QrDYEJfQdpRri
nO/LAJm8h9CRG+sLIyMJQ3QsUcukz6awsbpeuP9Yy/Yy5hCVj+OrGrovVSfH
5esY0+dubCRiLN93TvFJQOTnOwzhuJQf1SAkE8XcDnLWcAKaoIpLBT1UneKz
ec+ek5whHbQ6EgGxnbeC61Ds8KALCqWHIaY4FHod1dS60rRBnq4Z366LOImk
O8Mpb9QlzUQXxoODKRpCD1Pt5OYhuGk32RjJIW0xzSZ5iSlrEPAas7D7eKZS
8NTTvHuHOUazrcE1uLIE8y5vXWtj+s52dbOmlb5bcRsImeC43SgDZ3/DZfW9
RpqJVcp36DCsDd+9R/UFH/i2xIJkhpThiHVqa4F8RIGzbsAKAdzQWIX6XeQX
cXUnECM/Vwgl6l5h136po26oJwldNOyUwdF6JP6Bo55eVtDjzEuAtu4rCk09
EPxfAkYuay7MEsnVFS+AwP3ax0iFhujSlOZjqNFt69UZG32bbHUX4R2LD2bk
wXq81m4eKWB4rENYg2fjX7tUx98J4zvXHmAxDcKieB9JFV+HO6uemNSE1aup
1JWN5ou7twiMl2YpGR+0bkewL7eItuW1KFsWKtYaC/Vzm9HqgDPBAPeOgS6L
MRsvEHHmEDu6SLDOVPlKJbJaYEls8TFgKQfHeKtVufZlBEGhLjUmJ1MVDLcx
jtn//1wRH4XsItkokZG3yUNRhtTDiULO38Q2edHMsGYhO0W0bWdaekHXd3ws
5qW4RVis+SRExgGOTDOl/jAzIwhhJEoR/UnAUWwz4rM1a4ywTON/+YOKmZHs
B3298sSCDd32w8Z9d6vmE50kxVY+I7k5X8XG8MEEJD8N4SNNUIV1Ojwc3WXB
grRXlW6BGrPh4gMXRxvljdvBWP/7ApGTGERLsU2fjAns+fWF2RSwu0TY6r9F
PX9l928hxOW2E+l82GZM4HX6wE+SG+6tEcqLP8QrrYwROIMmQoErK2VpCqk8
mKkOYxasLMrW89qi4RhSS8ZdD+JiREJ9QwC3KFvj6MAZ9jODMG2cegwY+1l9
KheUTtVlnLVC8e+xt0gr/8gVWlMVBKPnINgAcPX25bC+ban2bOrwfBmAiaVl
/VolNikG58ZmY4VN+dgD6szJxJmfxbEJtA4Su1X1kWKwqVFf3A9ENzn4rZwi
x9YMD4i4BGVahDWde15/tV3USFdtPITORmq83ATBprjNI5dBrWBLhXKKX4iF
gUdsi+X9KC+pXwFrlKG26OqTZo9sof781yFP2MZdsdjsZBppRv8OuzXxyhVl
hC6EbSceISNAOIHpynIwbiJzqFWFrRL/ze+p87CZjqMQkXktMkrdchkS+LpH
raAzr2fA27VxOPiFZitddifOQDoCoYOgps17DuW3EoNEitbt4531mU5c5WpV
vepVzoHSPNBF/hkuYjeywQ+WDDq0OwYXWa5WWDm2reKUNiMnx0y98PIPyv1+
2wUDcuJpP3bfZ0xVUO7SIS+7Km568qKQhMigQCFSgt9TzoPk/UxJgGVhe4MG
RNAEP/Jj0Q4bf3s2/wzLLolt09/ycoFiRolDJb841kmYaErLJ9XVfL7EoURb
Ej/OWgN1CXwMxYEB9jEu2ymGGuu86qTa4gyXtakwpFQ6jmBmtgFVnfC6+19o
l2f1cX1rHCEZRIyliD4mPzn0qE+xrxDa7V+ut+Hen3rLNcF4mo/oD30TdN1F
tmg0i66RYIe7/btyJV6wpTCNrACYJ0EtnBVuEPV20lJMYUiZEuwJ9rhdT2PI
bwq4a6xt2APJ4Z4e5w1w120wqVMxx44Qvrn6RMbEunK9024VQQt3me8Q1wR/
oyXyUvit0OYLQvI2Qf/kvPxZFncpQN66iG1x1W50bwqY46ZG7kMI1Am/z1oZ
tRix2+Ht04G3FgLpzlMbYfQEsAqkI6Z7zbfAml7mc0bsAk5Uqrqu9RbH0n24
1pAFYwxv3Sli7IZoeD8OAjmni9m7/wQlOsZUejzsyAagVxGaBxu+XolB2nSl
99Q0wblIMKN1DcDPZltyY8v9C5lgry3gWnpiY2USX2fYJ3yE6q6INZ3jbpP2
T+NDjE/C0OIOHMQjD2gSh+DokltNZ1vLPUJiRUSDln00aePtFs3LNyUxrhaU
4+UItXrXqGLKLdrZsDzG4MROsSWCAx4frQe8OISeVFw6CcqmD3nv+CJKYKif
r5Q1Da+0dTLsHF0y0U7ir/7WD0LvhMkwMJrj2GeQO597fot5tg1m97VjiQAX
YTSRDa9w/eQtHICcWnWwOm1YoHymot32RdIqGQ1ciMz0i42BE2jfCT3dp6mv
u6axLMtZI8NCjL6Ffyzb6VeGhXqI/VXAwEZ1Rt2iUqL+XUOpTiFH5LFoNEnV
48yrjpIOQ98ufiLopgPBdp/7FqNxVzpUtrSQ3egmI4OlRcgDqKovq7mNxShg
JJMdHYjGMDLYBmf5pgAp59XAbteS7B5iejHuHdjrwvz43G8chujl8TGqqvta
mLfk1Fzx9Wl7RD2E652zN5OgLN37MZPzb0Wa/nSY+hPbod1ZB/KextlDOVlw
qXPyr12hyito6m8J5kGXfWkJl8/DeqKxMCCPeUCv8RL0KfjWtMmWPS+kmtsL
PgyM6N5Wx3j3tDR+FGoy2ZVyBDgwq1p9nvYHpUSrvnDR9hRPYfAQhV5FzdvV
sUbfYQ+9JMAXT3taXOJdZ2SbTw8irkuBZHxRhQ3hQnV5bq7hsitUti1xqfTp
5Yb++CnTXtO6uKZlKVnJTuIHhqOEABoWy/ZAaDg1iK321b4/hgbhPWqVxCOk
D1QAPx412/Wj8a5jB0EDPqYvzgT6dkfhJqp8iWTUBf90ZfEqufKDCHnh/xZn
5BatpUop9CIZDrxeBRKP9B407iWdZGBlwLj9DPeNmOb0DJHATU+paqtgWgfD
wVhKSvF1+LjB2DO4xmiHiDXNNnDaPpxm6ZK7c6jmW+g8yfJ14bcaU96oEEFB
tFXf4qj1gNwoXC3+F5zOg/DKPwV8fZU21wXYMcYV+g57kRsZmrhIbtsUsUmE
GmXL0SWmWfjmJdEcR8qsuaAbxoDHqUDCX/FqAw6d4Ik8V6PbKFWQ/4/qO8Ix
5vcPBK+IXK3bvVaaAkgUGE/zYqe5HsMMtpoDWs0IgUWkGK7Jkq5cdHWfGQx0
JPO8LXrT5Uncd2jIACJlV/08LBsJMEWvYlYckfvhCmnaDhNG/+aJ/dOqcO5C
4ZU68Hmv/5NXOrjNmB3BD/qFQABSoGGOwfcrUwtxKH7Z9cwKqVEcfQDuojWY
frMZ3/jjGjanwU8RDIkfR3zxV16FziRq9EoT6BqYC34O9DgWh90tjrVU38eC
TQwCZbk4B5D+xYvifrlSjIu4m/eaIeE1Ar+K8nfP0xasIv8xz+JB8+Siga8D
dOEWTG+s5iDD91VUXjOFSZDwEBDT0VfFCkaW6GmTAvGkWtG1p03AqfVP96Fl
s+7V0hxIv1jLkdswQemAtyr8l1jLKw4uXrtAHDbd+rolUI2CjpYgtaxMDdKB
RwzOdfJ1fXoQn/ELGR5P850/OjBUwtUGW5lP6w+by8q40mzKYHV+dfEs3mgh
iPAbYZ22lO7242E15azGXzN8LukcCde0TRWcKAbdykff38RuXF6TsUoO+U4H
DtqGosF48WQHRPTW7446QKDp2hLENrdvf5n6CqBCCn07og/4S4GFFqXy6SE/
iv+rUJUhIA0087SEr901LCiwRFBdpT8ou7KtkIg1z+N65oXOtlHrFJnJIhV6
Q/tW0wJ/LoTdWfxPa7Z2dWXJxlpNSAFn3ohBz1cKzdp1GkP85lmVkaHX0CeW
P0tuB/Tb/Kf21f19tgYJn0+Sp7i95op6ac5opft16HnIgCqSd3pcyxQ8oAeH
2O4czZFNg2YglT2HRA+7GSHAthT49qCI+puWI1X/KTHnrnFj95n7CDpZcmyw
WybvCAfl8KQfwOv5qyL0Lz3pbwT40lfDXGj1gP2xftgjFCC+enUONpWTaVjp
ZLztHIMEhoruJ5L2LIvYXvhGcB+Kua/iTsny3qH8sllpj162/hU4VM00g6yc
vklzOHnoRyDjU/L4iXWxnrZcv9eZQQD9wJtpHbiNv8hpIgDpRH5zSfqlAYZY
g2cdRy+dy+ie07z2KPusuFEQRKIm4W6IA05Cvh363Om8BvV0k6qjDyTgqLzg
Y92IVdMrhXErOVzeIzDEqr6B9XSuqnJjqAmK75dssYOt/8uzwe4sm6bl3c2n
UzFzcP1qoa1sv0nh/5WhTBLnElUbs535zfF6FeuKtv+0jMiwxH9DHlE/DNJX
PUAHiURBSGk84uyghCVHjyRfVMgkhcI+naB6LtFdXOOfUzCdjVGaFmGyOh3u
vJC8DT32yr72dltWHYCiex5eDcwqRUbsmg7ksBSrFtHXhcdcABD0of2jw0JN
0UpnLxMsF0O0Mtf2Rn21/YNnAE2feUm1JDbkHP/3dnFyw3TgxsDc2/n9uiMm
/coxktxOImd4K5cwp7RO2I0zhT8AfUGFdMlAtOhMajbKqZOnezrsr4BPlRcu
PeHl9oBi8z9GzyfEKHijABx9a2+D3bV4y41Zu5CKuB4Ogxq26ejBJdH/mqFm
9ikakECckFqb9cWB4thX7huC4WH+zPoSIcnbbFIEl9yPi494n1dcx4UQPWYl
7LeABBaY0CP0cLOA1S0Oi19Q8zkg7NRaQJ6OmYaVtHZEtYraSYiSZdVud1uM
A44PzxSQfvgwIWV2KEA1tNjp3rk/Ys1WmBsYA5hq8M5VWmhvFiKxYjQSR4nZ
qwUCzNbBL0rnI4a0fGwHTKQwEUw+SumS4F0D+zjASJaI1D138ZOo3UkFpf8N
dzoX7VZzvPAglNesFPvnj+O+z2DDu0D1D7biBi6981RHv908+hRMhfn5AI8o
oya2ACAw5+QWiryLTHb7LSrje+vUQhR3hikyOBL464DiVH5gQ79o7eAJlzGv
jiNKtbNREg1kj99AUHOsfDKrEQNRZmeIeaJlssMnldr9teIG74ie5D+B0qP7
+oihM8hTCm3K8raX3xgvUXO9EUt9vxBqu1EtrgFYB1ZvyM2ed1uPuQhU9oDa
1xHqLtxrdTkTR3P9w6VsG8iyxHsfulH0XUTa3EOjJmPVBKluG7GREdFCOq+V
/o9+ziFpXzGRsUUigksi6L/v1Fo3NWHbOOI74HLWO+l4r3G/j1Ee6jkEoBdt
RYdPk4hBfgGYUw7a5cTlhfROKR2K9tcTGlFVvcj8jRgnuj+cpZnRI8qsKSrj
8NpiAnpQtPC/2ydue3a0/GmvogNUl9EprKsp/GjEOnLE4XfAlhZs1KK7YHsp
7O91JlWqfGceNjjmcbKYeq3vOkC7O4FuW2klBt2VuIIokpTLp7yP/Jztvh2F
tUHwDpRPy1Iro7XnJ8rB5nWKW8hphapaiVsEhaX8+wAxuvjuz1MdPti4CU5w
n+/LscTBpVBMfhEEh35DXLNDgT6i+DUkfU9KyTqsTb8ITf5drzv7LpwB90uE
lm2IOCLQYAVSa2kcO54oI8G5Sv1Etk9HC3TKfNr66AIU/qeasZvayI/qr4Dg
iSqicM0Lttvil4RfvFoChv2aExKsquZRom+d6+sw/spFiw8VPE68fvmMfDXf
p5Nl++26818Kp2jU3+CvP3IBnfcI5w3RacZNhNinBhg7UOVHVTfEAL57MEa1
yc6A5tW8fp3+tjfbqfA5082RoX831Jz7FCwYU/YLSRuTm6S2WhFBdWXspp7A
LM+3yAvqrNzf963HFPn+J7f3yEswRD+C8dIbG8w8XI0CnheBq/O5LXSPlQSk
EHtyKBrWgopGGfBrfVmlZdTZFOqL5oYbZKAsXTFYx2w4y1rj7BeglHLeGurG
civjOgZs38p7WV0OWUtsMuKM2HhKjzowJJmCunZDMg/Mh09HZu03+BDXkJBK
PKxCBC8AltcFyUxRXZfVVZ+gDQgcgljo3PLSPN5Od9OUcVq4NBvgV4TzCtSe
hyN/Sx3Y+UTCgOHyn0O3UAfI6hy2V/h3fT3E2JKfd+ut7USxj4hTGEWQwmtj
Z+54fHjydrtcgGcN8YoYfImIcw/Vj/W0Fpo9rgbNRbqFaSdJ8/ZVWKsQgAoV
5rIsCpHOgoIMqwlIqH0vGlxnu5zo4yf3UMeNqanHeDV8zUHEhrtWZRJIugY0
BUep58YJB7thRZ/NLt89GsbJRgg7bo44/G+lOh3Ri3JlF6dtU+6MlhBpn56X
BLu76ln8yq82hONOuzd5E1CWRS0i/jdxyZKdwmU/QjeLbx0qKU6814ChFdeO
hQQPgQ4bvVKAI0aLbJ17YSFdeAWflzKxBzKelGs9ODdV9ZqA15QFk4KFCJ6r
ojNDybLzStgs3ffmdsoz6/cojXiX4q+jUenVd9mTTBdVJg0bbOpbJqKrImc+
DhXMtL/QCDphaBJBt/vZPt4Wk4uN0MhugpFsqMog90Gt0naxuoaX2pM37hHN
h/D3fVrk8lbqQ9MqSG6MGc1mmiewS3ofYhbfZ2yjp+UHiTWCzKRTlzcX/cIA
UxGoYbCs4fI4JTSxWWE/ff0EWOA04HDWSA0hG5D+qtdwPo+Lkn1/e73i0Ija
z7UGHHlkpPzUW62Ij61Y3A1Us8ColKRgRjilKxrvvBYAIgcH7QorPYVYLHXF
ocnLGjmiXzoorZ5fK73UBni6xfCmIZi55/INVGxAw1SSRAxAvtM6ZND5pXG+
eIPKQhLnbMeSeXYu9q0XJ0C4e2VxOdKz8/eQafaQo5EDWfot0Fi2Jowf1jVr
ssHUj53s6bJwRGniGeClCliMxvxoKwUdPUIJYMelPdoklzPbb48jw+EzNGVB
/N5a6lzcAPSitjN5BmFZFFXu7z7wpTbcKNZrj1xcIjK8+NCJ/Z/XqUotW+8X
EIApHJgNepbxQu7JXqLMFX08Bm7H0Y4tgaWbtalPutiwOV3PaZ5AZXR6i6kL
1t/RKJTyxPhInDcOKWUt60b4/lS8uf5UH+DtyqFQmc6FaX8cy8+jVOQiWD5Q
hvWsodCgLNMgagKSTkH6qWCn+lfwatXiGyCWv3dGBcb3n8d4hE9UP5WqfQK3
2OCNLXwFEeH6qRraDL8y+ZZ9wXFJLkmpRcArTp1p6r++aYYt9I5Q5a3pA2QT
CtPN63Qwg6FOU0QQ30Kbt4UqrOQQCRifpU2MtTFmo7zrigDpUSZHY5y4KIFA
RFRKysJ1d2zZSNetMv7p5YxNOi7UaknCtfYDBUtzsSvdsp6BwVzTn5Hgt19Q
imUiW+XgvsmZBn6GX2X+kVSalPFAw003mxI3nDpkKyaUuc+idcdgncan38ry
sKN53IJ0/RwLeQ3iM1guAut9U6EsbWSxK+T+ofdwuSG8ROJg4PzSJXNcvPNl
d3nusXB1AcIFwcnz80G4ut4Rf4zWpIjh5CUFUue6HSf03f7IEZPccOH0YAqV
11CRgyC+WVVqB41nVsEvYYUlresBpuoa6F48ut8xb5poXrxFGLcNNfY+643O
dJ8CjLpIcYnfw1XDFuBdAl1uorUt/eH4KJix251+kPzhhXNsPEf6H5vgJmwH
0urP+iig0XLNvkUEffN5PfnYzBhsyBTy0zphaqygQXKXrOaWJ5vBHQH5xj2Q
bBEboIiz4pyfYHwq0a21H0O/N43VNAQvBUrc+1hCaNp6JOvlqMW88meLIjSn
Q+jDpjiBK4GQ753voEY9D6Q0bN9xxsw/K9oOo4z8fEailjgLeQl5CXCQWcDa
1Ydo6hAIEvDx5l8Oyoz7PkLmX1AMyr/leS386aZUHCZIxCgEEyZXPSm4a7Kv
srW+F5O6zkzR5k4BBp0x3IuR68sAXevp0NggB9IyfimClDwtyhVztyGMrNvD
p661OoMDy+UrNBEQJQnbN26tSCHCEDiRaoOpxnY3KPwFz31PAqoWSoil1MJQ
lSawIFunooBPLDeCngjj1pA2w0iJ8Yo0pGPUkjgNGfrVIYbGKRsLCxAp6x1M
qz76RzLFNeaWLb6576TMjRf1SoZdRbZzxNJfkbpLsjN9dDZCPIALAW/gWcee
zypmXy/KBW3qnHvK983Vwg+vBv3dN31Lz5DKZd9iJHtb/FmIOvoeivLoUGNX
iF3PxyTyC+4LD8Ar+oo8YnKzLnSSFAt7s9RWs3p+seZeH0ktcoKCI4TZOguk
nW4tJrvI9ehZISSuN5FFKu3191dp7EcimfTpZA1I3ESdBQL91lf/bSjAwTAp
ieU9tB13q1bpDOA1OP7EnI6+1m5gizm/NviowR4+flP9YBUykK0AYpLE3MWJ
GFwDxKCQQTSvEBztlvt5oBwA0TWiUW2vvyf6ZwdphgmrXz8yYmD36110A3gV
V7jlM0rmln68Ew+H3zmyv9tHN2FNDtLkuk8KnQd0aQtwhuFtxR/+eKqDVfJp
jhRt50+JwXvjg2gnu+cXlD0CoS/ndglPn/cdtkCsM46T66Oej+8v5M+FJXEf
Ci1qWWAVeXxgHXrBOTLgLD2ADTSvh6QSNAfh9dezGW/vmfNRcxtw+a9RBRHn
WobjT6RihmCAqKKUtdPRVdK4TJ3xvU0n6faQ6V07V0/cdS+VrywW+ZNa+HxW
7N3oqOKEKSBgkZOZ0sDu+lumUWe4HHhwnCvpsTAGiV+XpzaJ2WnsJlS4FArs
lqwo2+fj6L195eckX2EVBon9eAzpEN59/8rDRYKaX3enddltKj+QXxp3sB8c
DDWZyfgp/TqbKIxrj3U28Ryo8hf7rFIEIcgYyMiy0DSrN7TI5pHt5vSTb268
CV/Km1LREbSrYno5Ro66ln+QTW+YkJASGxVfaTj+oRBgiqHJVbhs8KP6wXVB
NtCKCGN2fb/0WraAs9IZ+/W54Ur7q0HbJ1f25Tv81pG6oVwfByICs1EvP0au
Xl2cWyHfA+cJxy+ZN00341KV5fMaY4rK/gl03+rpN68mBKb43kkhmkI16HI0
SzFDTeJBSiMtXRcVE0qzAk6OswAIB8ML8IQBI12FyZeSmRreJaLvMx3p0GQG
UdOnTS8sZVR7BLuWYWeM+e4v82Jt8aNHBYO65SRJOM9IWGLhM/ASliVb7/60
eWLe4mXDn5qZPGSd57nwSTYt6dRx5NnivfwUKwv0YUrNTQlPGh2iUKqSC1UJ
aVdmVPHT+A04rJVC+XWi0lqM6VGii/04/v3nS6zm71puhaXGLBa/lmbJEgbr
LbybS36OJK1sL9zaNqTg0HYp9tlJpW29Pk8NLuV0LjRKbpN8/sLkVrz78kyI
jP2OjMhPY/0MU7e0h1ZOfz0NwMBjCu1+OO1ZpdrZek/6qPr6wOPbmkOXC+mP
+yTXM5JVfCNKxESlhcEVgksZKSzu+Wf031Uo5IJEVujom2N6fcJiPdHeo2uO
woycn1VaxEF3YNbUzY2NKLRDZjDcG2YQT9R2M+aJY04Tui9F5Xah1BtUR9TP
XmjuYLj1CU0jOgUH+X0xEuJGW0kxzN0GGanujJK0MRHguDxhzqCkO1ep9fdZ
AS/oo43yzU3GWeiRnLZQWSbAKc7V2vudeuv2Wuj4N6OElkKn6Sb2h+FHxqK8
oZKc8V2hGmCCTsnchowiSFt2cgLLQcJLaOtR4mOgp1gPxM/I+Z4t6zJWgh//
YGUwKVtXndH9bw5MpuJnsNgNPB8r1DMpdq7c2DjlJfQ6NZaYCxq3bdvImULC
XPl5VSU9bH+yPF8hqkSTHPpRqn4N0iRGRweGGZfpP21DMgDnCJ+kwqFTonI7
k93WV+ZRzrPgmksulUOqZsGN5HpMj/zjmdD8+dBdzc698rhkUEHznIdHTZF4
M6RRSGbS1VfQL2MVIE4DT08InGvWkf32+NIQB/A7qBoRKsmIBhoWb3UebrEs
Ci3w5MHHAOXD7jU4YouL515fT8edHkjuETVC0wIxYxIt2l2I292KOqLfWnbj
w2Pa74AmZ60anmi3UH929x09IyGJ2+8jmF+syEccs0ExPPGc8KXF3GeJj1Q+
PsklEIO+kwlg9kVZEUB2suITsB+0jUDPXFqNi69xxmtXLtoV2zfQ7fVIPhjI
+SepgIUPPeibapYqJNZrL7sZYfy4hsztAh/JHzF+FSvZKAYP+eL4hvOplfhq
bp/xP4jpfdrsgu/3zzDrAJBHmyuLojY/iagdm7tPtJIo49ic/9K9ciQ87YpY
5QHrrKY4qvhhKrgHdhCMjvHDsNaU0QcSm7ohutrY2N2ZsCre0lsicybPEoJI
ZvlHRGUX1jUc3/DuAUJhauMX59hkWCCwkW8tVq1VhpHLMMhHgMyv1hMrlbMk
BkUcdbSls+6cy6sgkO/D1sfTpVLlKRwdgTtNoxVkGQ/v61iwCqtLqC3gSO8I
dd2UGk2//1FYA9xQU2cxgIlfAebDasX7yYZ+VLTalnsKKcBFpoLdmXxYudFX
tjb+NNj9fodoae5BzHrV/13bW5v5CoFvpHQawiBgkmp/+VNeEtao+R7vA35l
h02TSYdZWRuWc4kcYCrtBAOZw88OSyireaUSgrlbSzRrj22bWdt4eUDyOAzF
f3giTG6n8c4tQ+fMbNJFSk5tinU+7vaNL7n64iiIowklhjxemEwtcRWqIkxM
1jm52QAxQdJRRj2bUluDGiAvDZp7/94vwuMFrentmLwWlFDjl11GFwgIIqGA
DqMKYhi9mH8deyJOm+TPtXFo8aplNAdNXIwhqFP3qaCxFeuOhN3HtA93lbyV
OMq0BQ/2z50AonO0CSOvpN5MWCW0KRFckEFtEfJ3CJYT7CH6APiPj0peaDiv
GVTxFr5Du1+oAeBCHHC0M0oB/2dYKNa3fly1sTNA0qqVHNVIUF5sp8mA8l+S
CPLr1Al3Q8lOR+Wt9BlvYzvwSZDJZVEqqC48tPVw61yGeQnvzafdkChOU14k
Vjg+p7ZmSSNy/QvT+aLpkRyT6CX6KQyBEZ5rZIHi5hrL9zViucIpgC6k0pKP
eEPXIg9FgcFdx8uZDXHlI9QebFwzXTI5RjjQUGmScZVQSkvZa5GureLTlVld
gLpR6euovyWGhXFqSdV7dHdrJzS70p687wFQyIbmELGDGYfqx8YJv5HFRBwe
Ctn3lZnXGTWNCiJB8u2vaimZvvBo+6X8UIhcYaoVE5ujq2xAz0iRLR5xvDr0
d4s8FF0WlrB5qWqDRZZoLCTotabcM+DLqSQzu3CxrL12WpoPxeg/P+GsC4pE
cTolfU/6ZXjL6jcqbJSGLTx+db7HTsLkdnXohjlYG334Ksqu12f3WRiSUJ0c
AzdmpUYHpm9SanL+10OaHCLJlRHuaIhHMX/7uXpO1F29M3pG+UpUys1x83kJ
t5Jho4Bz8j1NgLayVTyQWD5Oe0/wYXMeAgfF259m1ItfdbJQP9E7BnvEIdHK
FrJPulr2CdF14l0JrMA35Z3YCBQXb7Tkk+471KCfrII09CiODuRheJsVRMxK
6nRV0R7hWPrI2gDr2sapuFZ71Di/gyhQiLwVer8JVMUaH6P3TXZlriCbDuyG
sPDqibgpLM3AJcFJJt+6Bl7saUnbuiBCuKdaH2oP1QVK01ojfzxDdc93Hm83
SAtq9mWu7A/mNpy2eT4FQF7Sr2CHfpXhzS6dF7navQJrrqWBXXDfVDLmmY9x
HNlTL4IL9eDy6nqkrQe2gwRx6hkn9Db3gzIp3XV1jdqf3428zMayUjBllhRE
29FeUDDi0O7kkxOBBrXhfvD1K5P2pe8tLQEkx4Ubita2usRQWi8UrHWD2zqy
NZlvnCuzZ4yhqN5HaVNElyLZHxHJoEjaf8LfPwKN8V0HqAZ3w91VSeUqQa6g
FbUXu2qIYGUpV5QCEkmmrUjJ2R7jJPKQqMOU43sSE6CcIVOrtqq5Lisa3xSF
wXfmMdlH5lCIWUV4ze3SYOKbLgQnZveslfIk1+nCg1BYMXwQx/zOUw+gz7S8
1T4JUrMNEsM5yibb7dBnS+0p4ij4pKMDdA8T8Ji0yBZRQil0ATRriCb0zLgm
QLBG+janG4EHVbKCfl5+qmtX5SRBrPIGPzZXbdaTCa3TAsinWaxhOXawM5WN
5AUvB8J3PryO5UopRgiqSOG0Fb7ODO+YHFUCRiXAtCuZXxAxKxD1PJSNEVXE
umX2tJkZXoVQhmwXUqgbSK8dWkpDYt71b2EWBOwIuVMfIgyszBlrjjuPZg+p
FFVgKebbslSVsoqXnQlOsyXHjkV0alZ752qOiZ+D9uVyvIbXl72mgsLHeOqB
qSp7hJSs7mDxDO/SR79rjhLESkaJECQ3Ev0bQYPe01tkTx0KD0qqLhXxe1RB
aTu5M7sGKvmD57gUCPMzlcU2pVIHIQp4tUWwv4JSRHYvW7atg7hRvt0j2J5K
koQkQX79W7I1Cq7Z4szJtXson3IvHzB/ilh0Rp4zNTBr+rNQYZzMQBe9I7Ft
cpkHuwD+DCT2pFZEFHjxCjSzMUt1geZJwROgoEPhUpvm3qcNChUSzOkSwhrn
nRWE4Q6hTsIRSAfPeaAKHEMZWRQbtyLaViwD/3cImQ8L7DMIIyZ3Vx6GB+uQ
4C00kxFDPxujcl+5WSWKuKu5nP+UDZ+9G3woYuci7xOpdc8pMk2M1qYjNEnq
Eb99dRORqVO5fC+gHHBi/mWcr3R1t5Mzm+X9fAX2lB8Qs9xqfuPbhiOhlvrI
NQlngKDT1/dnNir6LvRkQgTf0LyZWKheEOdqAsCTeecrgIfelpfXmt8W1f7X
HfpmTgZ1+pdv7fI4uYSVEMQNXGCVh/yCKsNqi4Uz21jpVTcknhh51BHX/k+/
yyp7qq+m+CvOQS8rInZZ47Lnor8qeB03voEjW/w3AA3TgzFC6P3gW/qeEa48
69OkC1f+VKx7aaDJ8CKsSqHc8TWA/4PsW4ISiWMsalcTHUxvwFgNjvVadbWy
6Az2akLohwmyi2E5QMx/O6koCao8Die25DG7DeoPgNOUofrROtJTQLtTi6iI
D27R3YbuqVUg274B3vWL4tHELZu9+nLKVcnhdZWWHuKO7z5MQSc9DMZeW8kh
ROATs4hd2e3N5uL9Ri1Cv3UqLc5GEq6jH6/fBgobHlbUA5Gaai/rAegrJtr+
U99ienOnYsyCicSYG2mp+ToJ4JpScL7yihHXh9mG0IPf0w3dpDSKSDgMBaWr
1AtPXfIXVS5pxSQZxQ+3UsK392QiwRz0MMcFgfcCAU7b0s9/FNx+24ralHIA
ZN8KdauteWQx7KM/zKrcOSEQSVaccWO6n9aPjg/0jantTvw5RUJ9gcXDfsfH
w28ocUHo29wMxbZ6tx2O/3ic4urEl3ZrMO8o/+K7aAT9X+uSof65jPrsCsUo
op5qpMckWcGVrfIyKpIW1yxvyfYmyhv44rxv45Mw/Tn6jd+XXyNAoBztR09M
h9GAN6sjepSP1Fdkp/S+sxTqw/en1IeSSL6xwkNCdCYXBfu38iOk0Il/N14w
YJgOZHptkPeUi0c3ALLtPNi2dm5SjvaYG+7Fmocy9ED64AU1AQjQxcw0b852
c2GNuXVwIZGHDGcKfrqpaMuP1pRjSgsRdxRWocXhEBKQbM/ksbFcm6GRS0n/
dfcsSz/aknzoopo5U1drEPjhsdRAc7m1GSD46D0Zj2RMd21VeTiZQ9aXrqie
1a3eBrzkoblwuCa3dbU3wiAR31nFdyUyeL1MY1Y2auYoolI9tYJAljLvbAg5
DJNbloCr/w3FnZRhhKsC9BLFtMJMKYY4yw5EOvWIPrWzIeGYSHxR5ezltb3a
J4fP5q/5ozcbuwrzeSzLfeg678v2il32r66pOVBIKRT9L2cBMqVX9BjnfPrR
iq/YqOO0FMX1DQVrgJvSuDbqtAScGuKlW4Uy75mFanlXQVDCR2BSM51fd/4M
Ffk8sfok3th1aTgxlG/KlY2G/LLzX9Wa7e03xspH0Y1PCpk6/O+CHcCHwsUB
AFeiQyk6h+5Z49jaduQJ+2wQ+dAFXIg2i5CMH0kItokPEaYsRnvm/HGweynw
9ZgE6ZMGq386YJnJ4G7A8e/aUraB/HKynb8ggXKDKnuxWfjuWPd6LdbzPYRu
kdR2QXzhBxyqC6LyKYX7fxRu5zn9+VsdgCUd2+VQaemRiethduu71P90JXMg
NTwRh3wU1ebtKBfEFuasTEG4Adqpq2Msxfj6qW5eeCBqtYHnrPllvjqUBDYW
0HNCOccDu9AY+YGui7JugoOk+JrUGokhudbqxIL5BNRmeLJFTJ68nQjU8bKo
ddFkT+Wn56/+sL8CeNHc1R0B27hrTh0sMHYbzvh0yn7xGRJqvrksVeZKsxkV
AG8HauesJC4KE1TYUJ+xT+aGTnslGckt2cNPR0/Nhey7/WVKbJ8S3DyvKXFX
tBwNR9rON5Hnwmklh9EhX6nYwX/XXtIlSy1ked4VtIfLd3MbdTE9nhRpE78E
Qt2ULD/iz2YXDJGF4fo4OR7QUHxqM58Ncn/ysgx2kKDQyF7uqq2pDYv+5YEC
eOoToA+V1g6cOFiNHfkqSrF+AkdOkodpvGrJwtoEeTuIdWX59e1OXMsPPOXT
dadnB48p+ocRvY9TVpbeSP5Hm4BFzuLuF2uqdkQBzH8bty4tj+dWtn7oSJPb
Tx/x+//hdCfpAtRaMFdRwB2z/NdG987L2hynqti9Kq44SKF8lOl/Q3UhqxvH
hW/lpL7vj3a/4vQe8W7K+J3QyvLkMgFu0DAu25XK6IaLE1BgFrNcVf5KMrxh
XklXMoKtoTD6R8D14rsV6JTSzD9OrKS9QnkWWk5kcvwzBQ1UYur7RxZ9DjYA
N8dfzaJWBqsg4EdWTajebFRjphVdyQFAgyrlW0qaw9e63jj7rj/SfsnXfxQE
NOKlWnVetUfrZUsPoIniq5uvohDrI2yCoPj2Fw8s00FtAtXNRLIICbiUfuB6
tINrxTJC/mBi977m6UdmTukS76y2ScGikCTI/fZo+L9W+sGR3JAE9uKvKrhm
tNN+jKpVv4xN44xKp5/6ZLETFPRJe49xv5e6cncs0GmRJqdZl4vRwdveWgAM
rMh993Nq61CuGa+WjxEzI/u4fy1sZecbQiBah2CTGExdqljmf0fWJkaSAzu7
44mFQhuyXxaaQkEBmp6w9jiA0g+X9UEj/c4A4VkhVPVbNJL/kPm2ttnjGUyb
y8VCwpxpczr99/UDiEzjz958CfguQVpmQN+4m41+fAN8NseM0VoiLzZA4JHU
RXMXsI9mA4E374tNS1S2JoYgMzuqOw87iiynwdUDd0ifMgZ0sQvw3c1aXour
/0lh2W52gROjVEtqSJ4Fk+gToll5f3aAatkoPZfQVcIWI+yOR5nyKmrDbkka
+QmTePHZyjhF13QHbZeeYvqlJSzeEsn1Mb9jJG/FZC9S92TaMU09/5RnP5aq
MNJBxVPtvmdS3P69Lm1DkFyzYU+f3q60jTxnsPIVdTkgH4vWE+P2uE3PRwjH
FEvRhjq27PPmKy2zdNvO3t9iJDYsTCrgYnhm6CJF9y1uYwSuZRTQFxuQ3NeZ
FTI4eyvAudQEn+6Yl6FKrf2MubAFK4C6ure6phxcLpuRAo2aa31g0KYbm9JQ
3jEmX/yN5DD5HImBM41e1B0H+kIhdWVpNrfO82uCMXtaLEagSFGWvH7wgDdt
ZDkYpHOD3kSQBibDv93GYVJVChrtjpvy/I2HadlaMSTyDPjBKtOVLp4vdkKQ
J412JmN61DbpYNRJnmf7lsl+0V0fP7VCDb0UTd3yZWhEKGQlHsY55prZcIMf
PXF3a3snmbmv/RLvl/u0YeNM++3kw/Cdw3YkjOv4qB6quUpSCQvi5FMkT/VJ
EbBjeeFrdXTIWLwrir9AZzeOVZ8AsoYrJweiIlvcNi+MKKMLfpwLGn34l3NO
Nuqj9TnpCafzJEXnWnA73qS4rRA57jVK1kqaHQF5dDNz9B7TWVOp0Atb9P7G
XHfa2CKq5iyEfTrBigUFMpUb9flDv71hJAo1vW7EOVHlbvLjEE4MpTMlHxsi
Ni0VGTcGFZfevWAyAAgdD0fR9zoXxeeddI0MF1I1PvCKYquPdwv7ChMNg3DA
BFpS+VaPR7YGRpvHjNgSToMw0R14sjGGmWsWF7MWZYiimj1SpJ9LY2dU9mIL
hPHiel22mN98xnDbMbkcJoyXuUYWAI7ScchWwarRnElA+l+N7R3hshoZu7Nd
SMgiW3AB3dVZ9Zsrc5ArXyfx18FBSOfssJbOdRVSFf3CWmCznVcdytruGfEw
syVGiWpiocXyMRDweUpnUeJreaI4XVQnJfCDkitHfH043osJG6fgcog318jp
RjVlv5KwzE1VL7AQO6DxopoxT+oEmX5Z5MUMWEym/eOYP+jnHoWTOg/cknm+
9s2kRx7sKXdZo7CMQF/I42kfRhAknzp/pHOMpwhn/KRFu0xNlmGuEeOS0TLa
M3zML7LFt7H1LeZaowJg6zNM2mAz7MNUxv9JmEyIeJCMTh1ca3SbKCe+Zz0d
yvNJ6sT+M8jQ5p+vy+xphxCTV+/IkDTDzk+TeP/jYGPUtHVwUzxNwgKdEMh6
wbBZX3u4YYSeCMCARZFDEF+QPChRbTv8MIgRIUNwyPDUwVQKEUufHsr2QBkR
B8ekMN6/KvN58NMHS4InHL4YRp6lxfbuhGvMFmguG4LrNw9mg2SkZwwn0Hll
eGgEhg0d+24I7pquLY+FU+ALO/RIVrQa6lV50kzt1GuO6O3TWD5lW/s7xjEI
xCAFJSBgQ+yu3olPQKan/w9RTQiiuCXE8ekMEMrWDepatHa9na4piBO9X4No
7shBYyXnw41zFOposyurqFYzxPeM4gMcfbOtOXrkcquHXU3i/erGfMLfFBWL
Mpb/kdf9PGeBB6gcUam7AAF9iZIRxNd+V9btCQKJANXXlqswgeqAVm/Mpz0E
kD9y5+OoReFvEhHxLrmdnajEzpm9HX+ZG7Bi26+j2AtiFrcvX+Xwt4qIkpFN
rvxV+fnU84k+k3shCb4rsWSYW8c6gBZecDSUUkfvthCtouO/6Hwv8usVdsBv
8VNBRzn1bIVeXzz6dVG7crRfcORGZLz8RQ2kmRcKgP2+wrHcGSRv4HLDYNrJ
Yn3kkn19sYucFm4HMeTYO0KdBmwRk/acoFFolr8GHGNhruA+xuXI+1WKGMpF
7QFo3ll6JEwWVVEimsLBzpWtL7e2Rc4Bd+FrRCXj1C273Z9PhTcH2v2fEGEP
8ELpXlmD43sEf/cjidAKBUlf63yhUMyBF/Hrj4Sit97uxmzddTItkxSdIRkt
QON9p5xV6ngsMNivJyrtMaKD42hl16AGXlWAmFGH4hHXiTH/TOvFkxqPy6Hd
tYr60lzrBT0eEYdGwjxPej4MgJzFrYrIHv1s9IY1P+bMYBmE+6J65jbsztbO
syLDZxNNChTm/6HksCsUWA1ayzWcoQ+Eh68pAAJRhW+KnPLq0R5mcxUAYqAn
9eRuVyGurbAjF/EY/RZhRL4hRljrrHGYDq9mapdhUTnbQIrrkb6pWqQyNuSu
9Pn69rapDDlP5bCIa4A04kKdYOjIB6G2xV23XnNe/oDzF/ea9RpLFUCvuZHm
aRCtkpjpUJvTB2ssQAX0aNrirso+8/93uhh/6EO8pG01dbrsG29+I6TZNhrY
LCORu4cQfRgZZrMFexkDyJoWkkCTEQQEGnSO+Zvoyin8VOSz2Wu5ukm4XkI7
kUHXtmtp2LkWSCnQO9+TPXbbrqE1EMJPXsEfe0OY/+kaB4IV8JQuTeCMa567
CaoSb564NxwutAxJwLK+MBb2rGcJQ/1mP9tzyXvM+fBp+Ykn8v02yP887LIX
TQ5AsLl8eusUxmEFILJlkGPBoC5K095lygYAya2/yVpnyxgT8EYE24hL2J52
++dN6/ZAA76pmo9Zy3wBOO3TJqN6A0xlikapzJ+KPyBm5uRhxqpfmDbS3gYa
12wkN3R6I/591ibClyl6krpRuAgXto8fsi/cj1V00rqd8//zDXGjHe0HNuGw
iglTnW3bLZJpPRQOiWmdKEfaKdxNK9JrHjXFPcRY4GfLQ4Jpi9nasoKtO8EH
e/RQy5o1O80Q9EjQsitq6yisS7CTzhNkqf9INJLtzCw6x43fEU9CJL7ideUe
qjCL/LT8AtnEXGhcPPY/nU20cWwG+HWvwCd3h9n8lKN2l+iOzDeWNruIj1xS
ZbH6XHCBaGInCCpqrMpwNK3uOw63loQRQPvQYx1CLNtBOrMLMfhPbIXfkmUm
YGqdszfw2nEp5NZr9cMK2bD9wQYvFC+YeZvbEtgdjTaqVwvEuPveKPBdEghl
LQg4S07S+Obuwb8KXREjkfq0jOZlPVDKmB9iomwyVO5tCaWi7WDxn5eTNdx1
uZPsaLSHFDODSdDzxyFLlYn+S2n1uIHkMffhibYGLjjbRxD9mAd4AMwJf73G
yKTI1CbF3MA/KgvhHOlnsoQa7JxvaFKQga3rR2XaR3aRUYLfbYu6ZRaInYlA
MFLal8gUY7gzJLOeKiFpLfltl7Fzla3AA9DIyK/btHl5yeVH1Lpp/avljrkQ
Cq10iJUbfRVf35L1CRyPoipbsZRW5G0Qq1tdJZc4gpiHJNKYTrE+0SbyE6PQ
EmjtMck0dDGGPmbLivvIjUNjF8vFl1e69mGztMCotHW+HVaCNh4qlBd1Baqo
1+7PaX66Y/85cRcGP0c9looFIrDHRkSJL05No8WFD2EaplNkDxwCOnipNOFk
mGTKama72FHLNE4/R9s1uB6nxYCqsSt42jGrGuG/n1sMeL/WRV45Umou7jph
Z56vS6GKNuSbkLOPJasXI8597/LwdWr2H/RjKM2ISg8HVm2zPyz7oTyUl3KC
vFJWKizS3rNsn6rT0SVX0dlAldI8tyJOJeH8zww6BmxXcu596rvpEaxDjNCz
LSqQV03xeLxjT+oKBOuonwsGfNipSLaMp8gZIznoajztmtqJRVf5hf+ni8gD
a1BYSxRkgLyxD6OaCRNa228LUPGzjUbAnjGFaqAQrbnugY9vZgjvGvAWN57W
sOxfHAMI2C1m9HqZONXJWa4k14Q1njYXMn3y7MexoX3Wy5DYShyTspaq/Vlm
iVNpxhHos4AZLvk2lljSSSGyTOKxr1K0X00N+UqmRl5TySt/2O9OeWscUcVl
93LYDF4UzN6vJwH2nO0Or/USxoUHCo0P6NQ2gkqowfcSudGDBSPHEHBYZ7No
6D/C7UHuCjlasaocjs6TDiHNBT9PpPQ/zYiIapaqFg09uv9xfByYqibTAYC3
wqpigKF6KAaI1dlk9JJu9oO5Q9ghjrYPrw31CqXbXWoNznNbKKKqm3T/t74Y
0Q7+R7xQEPWfQGP/0cSCpkCJUVL6ou8SuTTg+VJs3321Kp/ebRTx0gkr6cA1
fwAFEmFpfIRl6372J72k0cNvBFE6XgKSAtrag/MC3LURn5j1kVqU+rbwiAUO
62tkelpOKyX4iH1WVnwey/Zj/zilMh50AgGs82h14VQgXpecM1FquOlNgi/O
/pSD+3lCDSUBav9VyORKNJV4RiDOxOJLJVje2kPmuyIdRbpboH2bJlqydP5F
Xx5j3GcOhN6cqQFiMONWfh95ecgS18OczcQNGL0zzGiOBRwzPvn2E95LHGt1
CeRGNDcoffT3sos/Tbo/M/wFnvj8ycdE9wGE4Qfko1A8d6CDUrRcG4NzSrIV
F2b1i7AySWJgqC44SgwA4NDAmGhy7TZriJSe/fC+JFjbmTooYEJGCQK8VUbG
VbDGu6hWyJip68zO5Tc8snuJpXh1bYMFFUCIA6Vluep1dsKO4eG5sr3NaT/J
cB4+k2UtQgIV/9Kii22ht5+9TRuJKx68gn7N60vsD60JJjsTCVvgULwBZTB9
kD8sF4jLI+rcZk0b1tiLalfaG7kGWSTgNEvpkNfdz5D6sMysMHPf4anKO2i8
l3KEkwoE8n2Ke8GanTwF6MIEItUtPdlbpHNW/meFTyq3B9+MzMfXipQhZk0V
5Sp/VNFoIl5ssweQNKPNL/R3yXQsyFe2YkN4zJimslSZTT1EjuyjUY93cr79
2T5FMwKkJxFMHI4AlbUmiZafR3SMsuECVwSIK/h5ZNm0Kx9S0ATXAPDL91rG
KKlnMTX4FJJPkerTxcyw5sJDbZcZou/syZOF7WOERR0NTQvlkcpegfu8TeTO
Nocio5EqZqRsXDFQw4CCY1pCudOWG4woZaqamGITycljsWSXiyqIPaHgg1oq
TcFsmUjoiEAuXVGnxjdKiugJwnwM4jaXiNmHaXlWv1+YG/J0tKfFriyAHIuY
YRH1XGRZzlawa2NMz2oTX7o0Id04Q+W6uiMI8K8HbidK3qmrBJNHwJPDHlKV
yt41ZwVZsmfEsC8BMdAeWB9YiGpldT5w5DDkWblJI1J1X32lp/rSNQEagiu3
0phG/ZGr+D7gpFCoZJRQ5ztXkHMTyYQzq3mxT4cRgtX5x8phnfb66Ig74NLd
eYb2wQc3iuTq4RXoI1YIvAP02qwZRTlPGwB+sbgRhzX8j8DCGDCIZVlkIdt5
Sy5O3GUFWjfBaWHFPcjQ1p6Iv5uXSSh2kMYuYuqlGGohM/qmLP1MhFcdyahz
/hHXmVyb3EUFGBjcl7vs2mwbKi2n2oRpHo4u+QueSgOwBXRcv/G3f+5grnAz
fx6Bh1xLlxVV4TqlO+9GvyUFZNn2CloVTLCMSPXCBknwlZNRjqYAGCT6NjtT
FzwihNu+FqYtL7q0ykX7WSOfGtXoimsnzREvX0ZZWzHfS8k7rQGXSI6OOxpM
2BdEwo00u4T/oM6sUcuANG6YEQf2Tg63ijYQ9G2kFF9eDc9ACucWUg5cra5u
g+epsW1r/vL16wIgJG+vhWFFojtM72KlhNATyywT1zrxn2vjwgGNSxaT7sFJ
cnIoH/hLCpMowR32beNT/UlIdD7AQijep308n79pl/XsT6u6Kl4abfZbSXmm
gea9RheXFtc6JefICKBDSY46Z4UYDA7kdiWG35rOlISCpj0tWPyyBhIzJI9l
54gK7ugWYXMIuSGfw3afHwUmDEeOZ1u6s7IItyuUNAs/EcaBCOgu82kQxKu/
jF5fJkIFD9dpEbiYgzci6bZmSxY5lHEq/P+CCDIBWr4aivUlawaV/IRMpkmT
VPizrHB0khFUdfgcXPxXZiBCs+e/NAD9vkQivEIe4acHgmiu6xdZ+QEUOBHU
RS7Y1xhnVGPHXzAuV2kl+BZeOB8LoRVZoJtuTdTEaU8nOR8jjOZE3PM1RG9g
qxdBJK5R7CroRTGJFIWE4RNIDMPjd2hn8QalGfrVAy3Ts/r6fivso7xokYO2
nRen0sVMpOHuQlTXCWmGrMUPJ9U4MVMHHoRSenneosrJYKes5zRyAOvkoLTs
4LFOPkqfTA4bL2cSOSh4/PVUv6sUtNSxfNXXNeEgYFyy+hOdDWS5uaEe5kqI
Ete3C2R42Ols4inoY9zZ+O8I3QTs2KvkaFhEQCOa68u4qlfIN3LCNYO7/KGc
b8jCadX5W/mtCJFZw0QwVRAKANWIo52hvxdji6so49aEgZ5AKldM7xE717zS
Vk5Foqh3TI9g1RXWDmXRdB9LKIeVnVPAH7NzoQHSqpIAFpda8fOJuTsV4tIv
gCiCcAWhieCjb1MUzI5updWhfwSCAuNvdIljZVWkozklTbuefs2tx06f5CLK
ZyZOPsLSc56muYUs31RGWcDPQGj6nzTkuAQ+m3LGaxEv6+0+MrCVhZFHVauL
UN3tjuOmHVqc0pAqLP+f0BlZISwtA2J7bMlJly4NdhOo16UytZfLJcGey0S2
Q12VxjxaxGgmTF9x92Xwn4T/BqL3BlFB9pRn1d8FQSurG2LEIlTlaF4/HSc1
iPMax7k4IF9G8gkuvHMobHaQSH4dd6R3THkfjvdPKkJJQ9IM3UYj7JaeCRsY
PVYXLYzijL1/Zov1RxVZ38UmPdEMDdEHi1YjDU59Gk8vEsBE+j81415xGzqb
xGN9PiW0rTYZY1I0yZoDX8bZv9IkxARl9nbwfpEcS1v+xuepm0eD04YCTJnn
hDkmTGJaNOUbo/q0AILUSPvSkm0Mne0u3vw1ixGXPZpt1Xw709eU7+caAFup
l18A6ucen7h86O4uqHkLeyDPh8AWlP8Uj+upqVGwE+Yb7fYK0LQUBEGGqI1d
MolZLnRay0KhQsAu2q50hoNEt8RmsI/PRPzEs0ejpzSPq3PbbziEWh/YJ1P6
EzJKYPGPBYUHuH4U5eBDOzqOiTAS+zABDAeJdjb4IVQMiqGDY8N3No7Zicyo
e8iyb8oVwm3au7iqbWKg+jADephdCVp0bVE2Gq4jP3w51jHo3ZnJSuwncMRe
Mp6vzAJizT5AhAbfccB3mxTdzaWcagFxKOD5y25+Tl545EZTAXUEP13IOX6z
09d1CdKFHEJL+uT4l5ty/6xYItzb6Jm0+Zly+K6TcGug54spnCkmIh6nf6/U
AHnJGJWLh3QRuOFS5XvQsBxn2G2n/UmKwCZCcO/5OH4goUklN4ONIRNeoG/A
4M5WUP5B3zragR9XU73iRVcx8zUyk+V/6dw/3oirZRu40av0KASzi1lty0nY
1zVXZi+xmh6wskxXveofkXY1mysYuPK8hwNDsvOKQ4ZW4vUHMhuQWO1kYmgI
sEHbl9GmvjwgG3o+RuJ68GA6TOYur/EIfn7OZ4sBx+wvcCiSXvfnIfAMg1LS
5fYjw1Os3K9JEAX8paXdo0YqAisrskA13ihn5zWKb9WZubOnEF0WMww5AaG3
Et/yT2b+GW/rxGjU//6aWqlNGUZ4kC0xy3KoK1l+bpACfMcWuloWbTD9pzJP
rXckUk9/IZoBvpj5Q4XTC67rl2QEcuKXTC7bzRLhxSlhovTMqIwJ7BX3800D
e/XdzdngZaDOH5hFh00Ru8ADwjx/tStxYS4AOlSmYHbOTDFWTxdd0qp0rSAe
hb+OvfNyxIXUamA7B55fZPdR7TgXJ2Oft6Ol2gv9tdlkxDYIWSXWMoVOyMix
mwKwJVs0S5WUkdw9PeauqECeLfWu6vURi3gC8LROhH5O8RCbZ5AOOBwxU1K/
p5+PZH8ZqRhvYRKooif9rb1VHz7AcdGwVyQ5yD2TtanOC4PwZI48bAYrW9he
X/mWDwE2XWy3Ifa9IxxmTD0mMY8SVaJQsLiKh9I5V8AkaGEpuwPyD60FfZwn
94rjpQVZF2SXoQBTy+s9MAZIDQTDf/KXh4VurOcAYklNYWc73qwpb0k43zoM
xKcLTEFs9kiOCdPCgWNrKz8BhwxrJkWpk+DwVJH0nBkea2ReKJsz0q+DI7fJ
hFxIe1Zfrc6s5QKG4cxSp0itmpnX7C1VhGw2owPbd5c8zXGzPgqRstas+aFr
RBN47k6XJ0XBE2wiw/kOdcjcwZTMbGYhqoKmnOb0d4vnlOJpgvepOQJqs6Rg
5VuuFMsy5i5pqBAvXLMdqakKG+eF3lAvix3GWRxWc10ONtWLSlmxVLnjWgRN
lnCecj7P5ZRtM+NvGEJ6WwGPcEExAXHGLsgQ9EaoEd7oSrwnNQSqU031s+8S
yLt9QaVtV/1B0isA0pdI5HDM8p2KBQanvUNSK8cE7hJghDXEm6XretnM6OEt
iyQEXsL2Xd0uAOBoB8GJ3WoyP7FoyBxuByJB/W+B68QVDM+c2nTEiGpbfs8g
n34Xn7MBIBtdvqUYpJv0ctRFNawPctdzbj9Z6NnAAdgqjiaRjFo3fSa1i67L
7SNDbJ+Gr99IOj/vd7kWyXj15tUiZx6x9qT2xjZObeYQv09oanDUDrJmXVqy
d9qfTEfQ8cJHCcT1H9ypR7Fv+Fkjv7oZ1fRyIyPnAJw44F/fDbXsGAfys1KS
ARcrTIuwg15QEWeChB8fm5i1R1Malw7kyxDVrKyzpM0Q8k/iG8FrsGM8ufgl
KotM7Z04PjLgiSiP/pTgiXeQ47zts6bhoiLTPgLhzYtguwpTNKHcfnO55SR7
GW263iJXF8S5v0LTKFWn+EG9dygKJ0c799oJD6n3/xviKSxcvJte01R215r2
dC0zxUUNuVu3trF1TlVcopZgCe4P+OclLhQ2w0OeuqpIF/TBsIPOtIhMP3eT
q3v/LZn5kUf2a7AshqGzCx1TR8FO9OO2na1oo9y8bEEeyXZuIgg+sXGeAvlS
GOfLTl+6YStDbFcHBBoNYsTVGrHCzQbVr3I166DMGSWh6Sk84RLSAzPacsc7
ysYjnzEtDgKGrwMQQ18VfRJkE/1rA2s1NLOcOSMc7aQcNtcOKQMHBMvnX9cO
TR/ic/Jsb9aohqrM7YJJXTGdG8sh1kvSineX9OgiT/scBdWe73tjiWu2Io4e
K89OKXwgyK2kjYqbtunu1JdFCOhX9RQNHWWYXfABatFC/4kZD4L3iJZEZYzN
l65heQ2wQvvfQC9BE0qN7Mx/MHAethDczRYtMglPU3RU7zcl6VKCEqjSQzng
5oDM4lfBPy2aVHYiLB5jlqCk0Bv9wvZPvTNK2UUj89hyZ+JAeZsb/yOAg5AM
wSZzLpOI1LvKOwSz5sOy2OAMrLfbgBBwAk2tGWN7M/8CqwhNeV2ylGJZOOus
wH4lwloEYdubEF+aHMozmT4Z0jzJhgQ5OrX1YTchqj2u4a+vteK066psWCjk
8tNTXJivQS9HbjIyDuUHHPLEw4K25ttOd+9i9JnPeodljKEA6df5FZ0J1bJt
jUagaRAoK6koCuaGwTxuj1fk4yBQzi8BlhSutoUFFlg2+ohaLy0lZyhApBVD
9/JShxiTJ0aZ7mChNvwFZoicsZYPU072zwj0Xt+cA7cO8DstkRlCxnVWq0A8
TPJ8A9+5SSX1yEQniDNqWJQGQUgMHICe7DHLaV9L6KKp2OjcxrKqavubVY7G
4EmPlzWQuRsDBz0Azf3TO6/4vvGSV/6NRf+3t1VmRvR9BhCEMbYWzqPiLKHE
bTahJqxLx1pJW9V/AqatBXXMPUG6FTXpcvyvhUyQpL85xRONRyCKh/3A6Zy0
/PUFc+8gfwZecQ57xaCVSi8pKU2fQAxs/JsQyUQxtu8G7K5f41y8bXYGDraY
m1M4gHOxl3QsuqNOcWuiJIUPPNzg2r2Aypv8Pj0JGkLyB9W7H1PdI8//sRnU
VeTcIRr7hGmYibtS3cL/D3YZnWK3aQfOpRoGPasd/xog4Q+uloDq0sY+qRJz
YshP3+9GHfjI+edRAMV+K83e8hfyD2q2OUBjkNT1zFBduH4pFxlg48X7b8MH
QkG1ecp+PwD5l+zukO+htR2ajj8F163HqfnPG3a3N9eTsxzf7fKlqkTGQsUS
Ct8aMgYoSnHQC39KvTpnCnex4qkAMpG5hX011GYKDMfz3OxRhn0q5wdueZfE
3Ii0rG9JF5NCz/2pO+DBr5Q8nhaT9MJpzHIzxK3npaqmQYsYQeJC56Nv2Xvx
C+yi10LDizKIPVErIDWe3hiR4xyeJhFpmPDM0ussRE00BV++EHY96PQPcRMJ
aIw/eDMS2H6lrayNLJQm2G396TyIPlNYq65LTJs9Xo8Ha3CQiKu+jW5h4khk
yo3ZzXdEPLgjfaQ9FVSUaF3VtNUr1zgGAGVKlMABJ7MB/3bMkD8UhswUa+Yz
kSjGvndpFqg0gpUoCJf6So7hLs/gh0xa89vjj/n6mIAS0+s4eA0d7VxS31Vh
78bjKVzqlzrDFlas/UHFJ2klCKuYvZ1wJ9os2FOgkEP5XCUFZcRMp9If+UwC
+j5gFt7r0bx2cowjiTI0KMSN+YizdNzif2IAb+612xO8zF1kkgS1oFsuCRy/
PsnU6cWuDExNBYNAd5VMlNXBPWuOVDI2yp/tM1lVvzv2eohWscY5JmyxEEqe
3+vJv16RXisB5mp9LAN5N1EUdxOtgkzTpTjeFC10+ymreduQkB6FJvHUwCM6
QEbcEvusDdkfn9VOGAjnTG9hJv+KGQiDVl3G5WkLRoBYvq9exx96Cay6NACF
sUF26m6akEbkKOo4TawC/1iK5Jep+86CFqqr0fht+qTnJx87BrNhFQLFMdlP
zf/XjZ/mIkRIyU5usjCjB+83rH2JNLSfQ+J1xSLODGBGT2lTpiot9vVCjSWc
Yw/Oc8OV5pZvJmyXxclcbHTi4SOEAFWCr6YaFkt4WTswZmU+e/H7RiLdqqLl
3vPpbAfFs6gPfVOwT34sy21xRg01DKuKR6h/+Aj+XugCfIAFSRcr4kiq4PNz
zX+wvEmXalcGS+6BEF37RTEknsH11j0p04/Jw8OF2BBThWCq8/lb75bHygQq
esGJzElw+M5rnPAsT5PtbJ0/VuS3ProBYHV+tYQ8yd+w1P16bQfDZLo5LNa1
94fM3ubNjGmL1TVs96UeVnJWjB0Kc28CNp6tZRMucxm6rI3Ch4pb4qB1HTzA
TltFEYF169f0vU3+xAy+ecL8GViIRaOxE7eSXjHCRARMo0WiXxS7JIJTyliS
4g8+5nIdaRmwEtvxLtwX0SXGvQ1MeUlex+KvaEIhYyHxxeqcJEf88KoQZ1rF
zMQzyNTq7cd4DOG3JPSVU9M2rUwhj9CuIKLC2WzLC9cRa0CsLKkyh0Lfn1pf
eUhbFCFVXtHJ5h+uQ3iOhkFc75AKYV0yDztHhhjfX0K1QGuIFp+d6JeFHJqM
MKcUUN0ZfBU126dK09fpsOA2yrYRr2QniM4kg4RvSvlGwwnzeKh2k9s3fTCL
6WZ7NafbTf6u7pRuJfUDZUZtBjHj5ETtiFKIDgBL5WI2Jmqk6Rli7KnPJ8d9
N4yKVqBDnlv2QqKuyTytN1MyFCE9FL1jjZyQi63AHEUV5MgTOAYcdSMy9IE/
uZSR2qf0wVNUJdgpEUyJjWgNtV4JxcCGQGFKkqE5UXnzuMWxtmqV0cvXBW0E
7GpI+pIJvkidPMZp4UKcCjvuQ6N9WqMqE3qJGccIXTcWtBsfLPCIn1nz00cv
0GMVITTaPEPAfZDn+zMVEziJ99rjXGQrxPnDRRvTzXMzREefvhZu+VmOOseH
cMQ4wSXowC5eoizRS4J64+T9FDs6isQxPEncYB7x45JyOEGmeKd4oiS11qGi
iCs+t9yPlh2deeyb2pZ+yv3sNYOfVOLf9jN0sFZ3W5K+s31AkEt47QjKNKwy
3hZBurkJzkesAYGdoNCd1z6QoVDDaYM88iPwv12ShqJeK+XtIq9v2Bpcwx+c
mfR0gGZQqePSSkSuOhND2Oza2HjsZM+RPypTt8czMLsohCH/f+bOhCJyr6ma
wlyg4TrMo+vdSYm1F/hIr9Fl7f4dVaWv+zoo/SLLnX0KSReVtJjh45H2/iD4
Cn35jLnxPGu5tJ0GzJnHSCyrSyyGkfWgBrE+lAzsQeBI0pagJ6DisSOarrMB
AC65YxsAHnnFYeE7V5cM6jCJ3i0C0MfUlT7Kj4T5DRGqEYDsQtfcAJQly4qU
ifHnBsn4nTe+xIemb1JsnNlys2bZnlHccwb8XMkrHoIndgTQPXo5zeZGxWW8
ScyuJHVa+0dK/Qvz8NgN4kuaXJypmBqrM3yA9j4uj4e0KjHXe+4bHac3Q4fn
qfK6HgqtAHKMnXo6/FzVGX1x6FvM7Mjs8IsLtLaM/YsDLxDGvHbd92LZmVpz
Shp8agMj/SlAaJ+y4JD6hOOJ7ecM86Z0razT2ur0ci3M2x9ZCHcOl8O/mh1B
VIfBVOMB4H2TCDVqrcyXNBdXTfEGBhphLvlcGUbmNyehHNaVts/a1rwmWnLO
Y8gmra/c1jbuADSOY4XcgaZNj/YDUnkySM1/L8zoE1vElnoOeBvm1igvix3z
1sxZIsXeVRVm0ZQmnMUnECxZvEN3ClkHzK5sA/PjAvr6LOa/XhPj18+JJdL8
jzj0QzIfcIHp2PX/gU6bRSnzeyQIkw1grqmCcmCO40TkKEhHvsVBm1L9PEAS
i691/GmGp/W/N9klUiRqx0yTNbkOJO+9J9TGK+3ob4bBVBIOjC/lFV2R28IO
SJmakz8U1Rn7eJgxSLSbbMuTZv6i9X+LZMfXc9PyHXq6hvECt6WAb6v3Wdzs
qdrd0UdTKrDc1nYoFRFA3NahoH1VBCxPxycXB/RBkLpXyYe7dgd/FbM2SH3Q
IVA3eRVIIy7ugFbZXmBxLD/KB6vG5dObnA/dXyf5i58lpbRVBhOc2dPvKXeP
36/lRFBhrSDLo/tG8kI9KVpmX39ZwJrvcoKjEveUHf3Ek+72G3pTFlEj9y36
Qq78pitimVfnHkk8qoKN1YGi6uWAXUO9W9x0RfXksPMoGbbOjAdJ257/r6zG
9IAtOzqQrMLi4TeZx+ltZN+MUuXNw9xfxo0/dmVp8ukGEgbvgcOJvXwi93Ax
s27mtJ5D1eB7+AyqzQQnIaQ5VVJpYTAmicWXlkIfVXKpMc1XaCI5LpL+DpWA
1cBHwk0Z5vsU7j8z0xiL0SqvR8UHOThIeooYDzD9LJl0nitTCAkM9ZOPXK79
LdGGtpOsjPlrmEJ1TgfUZMQNt1igfiMzF9LMShA792GoCgDVdK/RE+yXGgZS
BCs6NpNLuFU7MENUGY6N+3XdhdPdFyMq/E2byEiSfT5QO3AVHrJAABhF8X78
snVMlM+12jCbJaM/zpk4aoOUBzV3AMljz20OZnRoqwDhqa19IogPhIM/GJ7x
hbmx8NG8NiH3+FQmfe0EcryW78TM+9pvt3ZBw9iAU7iXYclvUzAusWM1PXUo
LllIwCB8vbC2nG3y6hr0zn9FDeDi8sY9/F0gHREkUhEP1qg5ip2XtFLg5vKi
z1O+ahPTxABY27Dx/0POy3QEe8KCeUCVSARN0yG3pQz+JWh93JePMU0GAeJI
/h7P2wkyIejEWwERYgx1hEU4Poou6Wcq+Kgkqd2M9wnq20X5MXHFB3uWTEpZ
rfs+BHp03IgFqhkLy4A91WReKw3vsPjyedwmydXKt7Y6UNG+3XM+A1LTQU01
zdYD2PkKS6Vi8cGd7NVzNomai8wiKcIRozShPz3sM+kc+XZQLrKVUO89QR0H
pg3VsYZrCiFN9vZjWlHCXy4bZ6UzrnAz8OeTGrRmHzCryczAlaHH2daGualX
Cj8Ubz9K2w2GPf6eiZTDZr+wmPde/MTzXrdm8gKf8FXUii6PnV1lu2aR6A1L
aBJcgcNqytKFLmqbvZ/aq2LTiq+1b8Qs2ZqOe+v954kyrHftNd0NKU/Wm6dx
7ycP8HlsIz4BZv5PCZCXaZioH1MYrNxpNmmTIr3YW+EWADVbCdo2jJGIQNls
y3gvjUbt0CHajlTzKpK5yqsCBCjsDlqfJXmbsqIuGcsfUxGdidw4BYDf6qYG
koE3H7JJnW3LkTJdvqMX53V6hgodC/THPmd5AlCZ/r6+9DNYE9Cz2B6K0kmC
L6DpmY59H4Er25NNVxuPLbtT03CUqK7FtUxiZAQUO/phV+Fv7MBHfB21iwIi
YiPuv8V1WndVyWzCi3LChPrGYfFRtF/x5HwtdkrkIaJyJdVQlgwGj6aF9ETv
LuEzPCipUziLSaMGuwi3xbhaBowiYkerbUBMQTHNtl9NmeGAIl3J2QVdXPnQ
qEk6HLe8o1RNbM8n3CXmQhaFvBxVrxOYnyKFJIXGqDnDz6idQ32jzIeX5D8q
eKrHxiLiGzc1Y3k2LQRQzZ+A1NTserDoTF5ZbTEZRGdEqtQyb4c/gUvZOcyy
6GN3JEgXOLmP0KMAVYhyOMOHGsxKnVIjXn688m5ry52zrsXKu9ZP5jk8yx/g
Zd1HX0uYdDCI51VOhmISdYkyvr2XuFeAxNOI8zgUfYxcNjR4ptSaUE3c6Or4
853Zg+QlZznNGQSVR4mIFmC6FaLyAkC8X8AV2CUgm4pyHw5L0QA+JCGrxido
Wdyyni3+Qn4RyZ7CzwLBv9IuPdVdLiuSi2MnegY31p9YNwZwFzEqKF5s2hn+
DrKNvVWgKPX7L0Y+H/qVO4tFgYZvvVriwnjmZ+UAJLmA5PZYR/5Bl+mjcLpL
TjtY0Wf3bFh5aENgnh9Wkzvk320nZuY40SgzkKdTMzwnUVpcT/Vxdm4gDoQy
uW3Zp8cDLTRnt9G2GFqWJULLBQJcn+3xXgmVrD2bUY+x+bjqUwMnP+6L7Fij
b6IxZx0Q3HHJk2SmrjNlG8zV9FGEZyki50vwcZAT4AWrxBBKQtvSp9oBVFg/
nzMwAcNY4HSxximI3yPFwRkCmtzdpPUtkdkJJXk94hRnSc+BfjIvWglxAUTE
NUKQoI2NmFlJG9SZj38VgJRbUDiyqy1wlyLMih4Ml3dN7p2kolVU162SyQ3p
s0tk8yBp4MSSgkNLOLc+lS+bDJAvhxKE/Ch24q75kSmLRDY+jxucM3dsoVjz
PEeTqCAFcUQfWrsw7ixzZ4pCnix7thYnhe5sgFIs3KAXvS6YXwBkENNFH2Hw
jbP3gvROOjSQ84+cTpJVUxLal3PLVl/qIONOWQX7GHwi7oUENd49edphyrv1
YgTvoLxzGjoOkVcJo3LRUrVliB0WHdOJPvQpZIe6ESZB7hA3gmlEj7wqOR5p
NHESUGBhYnII2md9YuR2KxgASiu6CSTuCLb78pWA5JA8ph2jm9cGb7XaXRSf
ZS4W5fOdf0JIw0ixaGC6VVBNofLYA0mZnUtI32Vdx/gvbbDoQpm5sBwsgsJN
pYuYS4qGSMhsjurPSmQvLcZXZ9mWFt2YUvnfslAp6/oiQbswqnTfhej6v9ZT
+Ok2OVsNHAYqp9OFX+Mtu7zVY5o/lbgvkAawGRjfDAGnU1v/iYQrEk0bjJMW
XV9kcD4tTYUGUBr7K+K00FOILWnq8drh7DiO5/TdMPrQf4HFFetq9cUqEdH+
lGSjBiojTchzBu1W89yrhumVUOM63KKwG3jhsT7SgfLaXzF2cVc5BxxlNN79
QLf0UYu/5EhRRrd95y1vYQ6vML7VHH8mVj/pdfgnBNtUfIPXotMwfsYY7dk7
vPQ298ZTYQSmfMOUB4MI70ffFeByYCjrgemHfyhGEli0wRN3cwUJ/k7oARNP
6lj75xeCewJL5zov6P7u93UoNvJD63lW2sMckoJxZih96q20iTq7P+ysz7pN
C+AGtGBmFj5QlleYty+PJQfwuyFdsjvzpNRtHZOWvFnLcUPD5H01VeKc4aqU
HLXXIoiqnTcNcGvwiqlNk4ts4SMAzyM4eKvDAFC68SaPxux9D4hz/3P5IwVH
X9sYLH37w9PSLjjHIRQLWR3RoKLZP0g4UmN534kVVeRmjJbaMeVKzP5aVqC/
Dg62lDEHPyZ/0l3nUqeX/gihi3v4Bzom1DBYYgsWrNLWHZha0/Kq3pkBCaax
VSriYI922f+3aTSwyVpQZTlBOJo3HbC7fj4Rl4JikIWEWYAnNi6CRbhWuM/J
iQTq12GmwfNK6PMR0MURSCFJJhNSp/o8hhhAq0aHDo2fq6TjuBFnk7JTxoHJ
qSO4CG51ZPM6hCHSrMfE+Oag3ofCC+axreTHStR/Y00cX9gF77UOs6ds88XL
deYEG5JgHBKuSEklgKh4D29wALT3EaqbCTHpOkaHVhKTJPngS4B7iFvS5Jf6
tTzKMC49QZOFdxiYvAksJ9ULH0/wb3zW49aCEva8HqLSLpZpWl41uK1YaCNG
zLYhCu+ZHkvtcReG6j6CG4B19FokBQ20VZ9P/IPJRuIe4qBGREV5uEDBkuI+
bwPocuC42jEKTW6jJn0qoa73xzt7jJDdXiQWhLDHszcRqC9sckFr5UguFoMJ
CBxQ1SLWBYeCTCsJySurU3J+kQSpDGV08B5YP8RD3/4BnKKkBC6hLFgDXuPg
S7nsa910ojSPVyQ25Hbojd5Uz/WhqwmUSjwZ/TFKPFJNRRGYYYA3J/0S2lYA
bvJCytGVdszj+j/1C8a6E70eRGUN2QCjOwvU6x+YiEAb0nqEIBviO0ursrYS
1a5Fe1gtPP89URZOtG+HMP612vE2BcbHCrx2gccIw7AZSNL7HPkA35VCxiEC
cUs7ZEV+aKdpw/yjl6ZSUrZRV/94/fUPWLmKKMBGUohQYa6kolrhXb6h1eeZ
14blxAHdUuEBQh+XLMBJ1C7JLBCj3BSylFsYDpWL0vsHKfew7UK/TMgaBTds
7Hh8567IJL3lRPsnWcOSF4zO3oABOxG0/oJx3pTqLg/f9BqmWC4hK9gZg0YL
vENWWMrvOoxGo4WT7NhNdIiHT2+iABeuEQQ+skJod0jlsO3lwb4glzHt+54h
lTMcKxv0bTvhrWd+d26VytsWcEMBx/edWEKd5lWL6t/JbLBK3pJA2YkaySxN
v4r7uHvQfvBSI7ivJVTZs9s+FjVXgNIeDCNBfRst60mWPtOCtRCVm/wPWHD6
5cdvAUobw1Xywlawn1fpkqLZhcbq36eGSmQ6ZtAhGOO+v5ZdPrfyG/c1ZojD
/SxmOK6N3SacLhSzPOrmGlEaYl2sGdCpNlJPFbkLGInbUjPYZ5q3D4cGDjEl
/r9vOyJi6VtAHVG6nMx3gNtV1aZLSIG/KYO1roYhF9cqx9Wg9JS5UeAhemSt
0bt6xAJSWj0cSrGQNFVVNC3BqBesjonpPMwfYFebGCLvP6i5yE+aZdOOT62r
CWF5haTWlyGKlA4lOwC2313c29xw7nM6rzn2LCgPcDh8js/NAIY5uB0xqhtv
lWyepFzJNJ1+ojUHdR3kYb/Ujevo3kdcmAvSYddcmo+W71oRN9bj9fWWfSTF
SXToZLq8eCt+HCxscCbhPV5ViPFK3MkrC7NjSRU3FaaafhgqefFI6YmFa57W
Q0JcDxsRJLwuTHQ6oUhJXgEd2DHybSpnp2oUufnDYXdAXWMapsaKmZwfHgX6
kbv8grfCUThAPr7oeMlmXhrXvcdcYcta23I/2fA/K0SXfPPx9JHVqKgdnxTw
STd3Tnq2bPIDILLVuWkcTswfVjfLzA3fXqvAfJbScwDRy9XuSiWjFx8oCJ0A
LYdBLl6QC8OKmie6SGBEtUiUs5Ii8McejxMzJ/652iwcYwfv0zWquNgO6NY/
FDk8ZPp9NOfq1wnZ44CBRARMryuvjQnfCgVVobcitU6ciHrByUfKuzctcXHU
ztdTgSluIhbvYRNlY92XBKK2Cq6eWmHk7fJTOBkfmxxy4dFf2cZoN7sOQDzr
/IRkvqsBQZqV5AIGQl4TEieSnH0NhHqSYpdT0mPLk9gXCDiTySg/4hNHA7To
P75yFfhFM9Xnr23IrHzD9f12R1pdm8D1Wbjc9KV0rC1oNSfNQUiWpAxbNy2r
7v4Y5sF/ts3gChT5BesdZdUYE5iKmZMcM1wt9JTGsqIBiuK95bAIh8PaK8+T
ca5TtL+WcfhaV/wB3MsD3GA3PIVSDHPd+4EINC/nvNzR/VCLXEHZGJI3Bu22
z3Rl5GRvKtcWmH4yVgdIklgVgKCTjCs1w4hZC2NmnyuOqPWMqua+8aBTef3H
eyHCkBKd/xeLAcA7e21bNzhXQR03xlLKMnfR5dU7JhmNLLIkbiNH04HkhEAv
F7zNhf+fbE+rA07/riTSPrAVWzDU9q/LCNHrAaiIMIJcGdW+Tp52Y+Ctny8L
+WIixmfEX7MAERvc8KxB86O3WaFqkqFQw+atNBvUdf7ZVZIXV0Up8c+d0Fmy
yoFKrduinlPifwFkULzgO8DpNoXTNoy8D2BxkO38HcPtwEEgcPb5L41ZRI0I
6l+tM7AsCXR4KSrP7qSuThFJVQLKuXRDml2CA9QBy9h0JKPfaFd0oE8NXsFh
jpq+B2vBwlZR/k/JYiZ7P6OgCk6B2Kzd8dF5Zkp74wzwMXQGQnMld83lOgIw
3zNP7KIphh9YPumtsLi8dDN16NI+ivceME0JYAy+aCffzDiDLbHVK6ZsxgsB
4U0LjSngTymbAh/XZLqQmn/ugRUF6+76jTyVplhuLIS8hXsnwD1XVKd9FfQH
wAYRM165NtebtJEqUvg/pAVNnbOeAaf2zzDNXmQD+Mo09O2KArcrsaRu7c2R
8jT6k6/V60GoZGoFPByfPS89O7/0E146pVofnoXlB4emUkmcbpjHXXVcGUnI
dh3nDNzelBXczYtxv8kHni7RSMCXRZKdSve/gl96xzlK8eqDurW17hHZ1iAS
OIKi1/uDAyE4fK2zQ/uAcUVALsHITucnB4LbE8I2uuybItD5suV8qPtrhcU1
i+Rz6HyYKT8Z2iMMOSGQXDwIggZyRmvC4m7TzATyjUuBTF4Ey1HSLpl9Dl2K
s1AOmghwrzxSkboCcjfMNr2z93qco5yHLhltpg5h2oz+T1NtZvtnbpkNWaF4
FxKB3xJBRj7U8YRs/I00k5omRho4lW4o+OOIEmDokrJXoz8U354hqNAfKNXq
HBfXtzg05QhcD6xTxMpIc1FVM+dToaOJyrrUAirYRMKG0h2xob/GXmMU1dQ5
UPYmws76Vs/Zc45ou3Lu++hQECS6bc3HD2vBwhvmGhyN5EL9uqYWxMUC1y1m
GzczTHLbzor+d/g27EIXWA9fKObwqdYMJmsdFAEQXwi9j80bvcDZrX2gQ+tl
rurUxyez1omYIW7yJdipGxf51CqSnbrTF5HvcKD8PUsyi/ONrID0prBeiIg7
2JtnuaUBVLO9s4/H1gf2JIx5CyBUhOTXPgTjm7jUuHsY5lXME+6VsBY7F/xk
UCXULBhoiCNngPCd5wLcsobYXQhLROKVqtaKXjwSbo6x+P42PpJIaEPxWbI1
jjzraBMSqnvVckVp7idMIzr2Zg7A28bGMWMLAWsRxCqzf5SRiYGVv4Mn2nkR
drZe7UNmORzC37ZyQN2yca2XbEbubKlnzVvgUyG88wEfsl/CtiLRjHIoLRDs
MRLbreeMD5l4Ot0iRR3nFTpfqntk6mxAjMVnSgGSpJySfVORMvC89+syPPiw
zuf2lllDzuWkAAwTPSjg8fIbKPwuUPHkjEIQs+0PLXX/gPjESwIUJz8chG87
5VS/mt8vVaxQe8MjV1RvO8zycsAivYJ0jt0Hqmfare1qnUpCYea0O7wRkZYP
xoeEmF12M4DG4Tl2bUKJ8eI1NsBw4GGuJ/9JGWukIcXjCxZWrY7JUkQ/fjnE
OvVv7uI3mv/GRdxkh5Mb8/+FX10FTmYhIPHUP5WTQY1o9Tm/2qmC4EphsGWq
ybx+701S+BDDfFlg2iDq+OnaK4f3blNkNY5/qOG1WhPkqiOiQY2qmToHQH//
Ww0sARb/6Ue6ajeGT+zDqS9hKL1coeiCMwJcih0aVYtffPqcI2gErM6ul1Ot
/7G0BPaP2XBO4ktw6XpDCs0Jr7csBkbrhkDdwM/BF3WppBVT0CMfyRaErdEE
fNHZtywoULhnHJ5uWXmEgkKVnCRutd16gR11kdM4ibCxhXjYFtoQPIUKytZn
6Qh1xZaaQ5nArmn5PagxBdN2xis5xgBkuXCN5RUBQhrCRcFXhVYw43DVQvgS
UgfCPXGTvafnW23tAbsvTU9tEXDZm2PdIdqtcxR0/SOdCUn60kOcRQRvaAxe
jmejrriugctCQICeUZvTDSEkZ4baEPL+Kfv5OI5tJREExVaPnA49qf/hUIxj
JZEzdBxNSsq8WC/5FFM9l3uzVKcBUuBWaRhCAv3QyP77OsbiSK5Km2ovD5FY
aPbXv7V8DRjnOckWwrlGKkX8ZMZ4tcVbVn6nfXkIEFBkeU/IWudugOspM3dd
SHr3FwwXtcpmpp4hDZcgrlbwNMWF9Evr8tTk5Sldold7tCtDclpWGnout3U4
b5iPRgL8MhPSRlb7vRAtKIDbIGAR7WHl5HC7NOJqA2YSb5c1c8mDTbLm7Y1C
p7XgJF3Qaon+IITPL0Z6zqNOP9MdVZWpQVyQ9EfZKfrPQlyZ6Kdu+kikFw5b
xAI8k4cy273kRFioaGKTTnkPVWncTyvlqwN9QJ16dMXxYMZI+NpnatmyGuYS
E5PqZmiK64OQRAbu0PKAqDw1QrwgyXcRohrXrKlc6PB8WpJD4fcxj8zyHyNG
xnnw1T2RfVq8rMTQbjzMcTTIiOL7JK0JQ7b0aboB6Q0g7NiA9fh4AjwK0iZO
fiNJ2SCRj10uKlJb+OzcnkDfTDhYC5IAaIGaoaPcP/MU+KyCfblvU6YoyKNv
oVN+vnET+Z78hMrblDqIKm2IuazFf/2JOPMZ4YDU7S/tY1FBFqwK2YomYMz6
ANY6S7LjgRrCDlMO0mytxsBSZ8liDtAvwVp1+cyJ8TLQJmZomo0luuaUwVhB
Iu+c19FnSlLLr3WPAitjCOZbY5k9jVtWBCO+PgOL+Bqq4dJ8cr599pxDS6Ao
x6lVKkQhC5SKyc91IYNoLu22Yv1qWfzqt8++vBRhN8QMgWXgP5pRoXWduBSC
FAT0UNeAgjYJUoyNJ8AxjD7fQO1FTSt/HxG96/yocgcnJuSsIn74ADF9FyIR
J7X4ugpG3s7bOAdXrFxTG4QcUkMxcBN181w324W3JyYKpRc1C25E8uZCCRav
JTvSkNMhP+s6Md4cPIb9tCH64srp7b2JtW0hjbAY6D8XwFPid+NrDYSGBNWZ
xUXXf8ErdAgv28/dzMryFPQ50qTg7WqE08K6+54VriFdhiEJ2zksYYpLQ+v7
PrBPVp/cD2SJ/C55dkH4nTmyH+XxMVJXH91fmBFddhJig8DnpG4jNVnqAfdg
f+JoGdVV79TAptfP99x9G8WnysjMBUv1x5xcFgBXPfoj74E131DvHXfZdMR9
MwtlbiKrTnmu7mZ/iJLRRL3ZnliYzihS5A10m9NHYyrNDpBGDMM1R6mX6x1m
19fYAoImCoHUKrRIBsibecBF0ZgpKMNneTE/7caxk/lGloNCzyKLaVjuNiDZ
4Ox1pvsxBlXzNduMyLDNp3bSyPhfHSLMbuHvHrFSV5WOWhxr7M8TU3/aQC0Z
KFx2DSraOqkrbWxh1I7dh27BRO6YQH3jSqmoVr2qr1cXYwrtplHF3GTmuQk3
C+I6jejRTbrhWcmHRgiJAhbmK11CCZx4iMJFrGES6vO0mmzu6cNUfH4FZaYI
uaX/PL/P7gJVTFH8iUaWsjNyQeIsO2II/954RZGvK8R/DC1Ea8dzHao2jG7N
JciR0rgSQGZFutI3jwGc/N68LD7TjPOt2gyiXhw8UyYf5KwrKFXyvmiLExNq
H2QRkQDEW2pBoU2mb/rMsLji/+22USmlXSVYaUv0U0/yGWHbORG+FI4AQauU
y108LU9luE6gHwbAsPp6bPN61QZd4u2FGUku6G2xihXK8AFAxXK6XRxP7LYG
tR69ZsBj2LRgi4aBMpngxJqvmHU4rCAOdAOc1xddfIj2uJb7ReNKWQem4Rd+
N/9KQPhmt4ZOT65/UqSvpm2fbnEExVYN+lb3BWBKHbhS2lvqgKeZhhq6xaaX
emCvf8iuqutiJtVwjonvoghTuTO0scUc3BtYQblQ/EVX/FRmy6fqlp8throd
V9WhXvqhJB/TdSaw3i+kTyKUkrhGT3zTEXUFJfcpLEnMS4V27aFLp+sfe/RH
zsTWlVDm83JuQgfH0z5arcpLJ2Y6BujRNAh+TqxbEMBMcMCZGKUppv2Ouq60
LLtWLp7/2pTZih341oiLtAtOKS7YDLpbX1lBfCoOynBPJUMN02o7KWXA6tmf
ipaEB49qBgW3fZDrSbppa7hX9Oy4KtEoXqeJU11G3985ShaXNw84wXe9hTKD
cjcdWRE6HvFKB4582rBP4TBdnZDIM9YmAyLy1aBfVnh1Kp7a6r6KJ7ntTxGq
QuDZle3Yd6Brgz2AWFX8fUE5Co1VgS4vWUpjlsUflpHhdC7adwRDUMb7mdP7
8S8a1ks/oY8t0YjVfKbtc5RujyCqFOT8qmiLSgSa7m8db8qf8uOBRNn8ep5P
UxpINPhVqyJGj4rSPh4tm9uVOFPipLoinqHTjIXMqS+R/iZWalBfNTckaz+K
t0wa+O/H0Mbcfu23nJT/5GIkMc3AO6uWPSSCQX4fqS+VYKUXUKEr4v9ZfgG6
fcetRPQE04GmPdFYgnePR1jZe+K1UFUzwnMOn4Tg728PvS6CJeXPKzEK69/A
nWSBEVFunQHiD7dhYISbvai+/BbU85nw4RIy9/MKkH9qWmHpYce7lLM+IdBN
9BjY+XXBjAonZrlxSNHPDyNOqkatqMudc5e7Ei1CoziDOy4AUQcsph6cpn0/
W7mtbtToFntNM2awYQab3Z7oDcfNlPvrLWo5r7luIVCqU87QabMmJcCZ1EsC
MyUpYqpf2p9ozkb70VrfavJphO5amQZ75iRujTdfhtr+YBO8O0ROTsNEglhf
c4GuWqRYbaljYVBhT9/NTcYzrqKLmx3i9m0cgHyIJsLfIkmfkwSrS2mhzLXY
/qKZG6IZxt6BkyXr+0C/cD4yrtvpYGprpto3XwK7mfdaSDEbQ1XgX4jeIFf3
4MIu/2gijG1K9MrxPkTRdRUMmDt+TDQkX1Iu+W1Kb6ZHw9rHYKGad5I8HOJA
jyf9M5eB4fBvq1vbH5pE/881qCPde+bWypnlOlOyp8B0d38wSIqdA3QFWGAq
dzq1fvO7Gj2sE64vIABQ9s84qeT4w376K0qpidxaEVVnXZzHNE/nSQDkUDCb
Y7y9qMxGibkxIlbquJqchhRISd2jBCn9gV+or5AgMr2+r8Q52NbURIQuPKhk
7ZOFhYYLWLMFxTJ3kS6kCn7uqoU3/uW+ohkOFgj9tDfLTF/Qr8JJWZI0ZE7d
rjIkDxBZe8PEaZxbJ5mu+UFVQWjbwyzLoUtcGk+y3pgEQKV0+4FFLCiVT88q
h/4BDouBbuh5ClcGVEpAvMyXrYbQttnGBIN+39gbQZT853wIDS7fiN8Z2ke1
LdIHIy2LsgiQFp1aRwH5zx4AXIn5gcuRwkarPLrM36X/96DW2rG3Y3f7+YsS
FzuGoawi4jR8WihiaHJXMFHuVxFfDkZ+X+Ok9fhxHvys2u9NvIjbFVkSX/uq
tloyvsTyfhCF7Xgc7XQpzcgHHfiwzI6dIO76uPZa3UisjcJo75HUuSojNjRw
WuJNC8NG380l1Fea4WBCJT8Vsp3lfJgJLuGrX6XJH4ioTK0cp5ljcVK2meSi
sptMxfhM/mp09bPCt/ZPnpgndAnFfLjGDAJyBnHcm/9Xasm/2ZOHVzIZI4f/
JaxC5/YAxCBmtFotxpifWnRlG8CPGoB/ENBMtCOUN88hjA5Xoq+yA0qYnVHs
tpxpLN5rYbM4DDmxyJl39rusGdyNsFaTyk56S10JBp0uuNo2jbnE+sveBhGb
V6CBsSrY8Epqs98zvCZTEHZIPZfsQjNVT7vCLN8cMb6zRxDEpUxDJYfoOZnt
J5N/IoMrecl5xaE2T5DSRtZpJ5NHNR5lCBiB69zNnDIOnTwkWxA8gcwGENEf
kCSv/B69tBsCHArrzfcHZGF74JiXE/3vxcJ+61j8C5jcUSuQ1bgUn695l9Db
K6y2H6amcH2cgAMWhECuhMIdOewLIYpJV82kXC/rOBVd+yaO+bAtwTAnxSu3
XVbeebocIxXRMUiIokgWc7UfLW9a6odHw4FTiuDtD69FSK9n1sNCuCEUvf7e
P1Lrwc8l3Y99qU/k2R2HENXT7eS8moOmGzE3ml9qhii3aMrNJuldrb4wmnWD
yl1dtsKqw/uRu9JgBgeu4e2WOdHJ0buVK+zGHP8Kg5pok3uoAnIQs+Ohqhhw
LwUYHtymNtxjroPTUejxi2jodiSa1QarpGy1PucFhyJZeLl7dNW2lG8PsoQ1
onDbx0Zhiquy2XV7McAA6G1xnIfuyoel5Xsz5r3OTOm+csHjwuvf9su4NvFR
yoIBlvhBER9qu7qUQUHDtdLRx3chrqyo/jnFSH4SmIDoDOKGtP2wcsLovk+o
C417rlVsUYjNFZIVCPqdAWqXmX+c1wCEnRs9I0gdT82/r3WFkf7sbyd5/NWZ
B8LPMjhcAIDjUFAVtfZtYtfryhWoOfwmArSLvDBLROkESZIhChwTqEcEhmbI
XmA56J8k4Z6+se5dfyuJyMkm9HVCjSMYAl8xM2c1LcTIYzcxrHU47iC4bE9e
NgQuB0gOK8af2puNFfRFwRLc3X41aiu5szpXXnFuxrYf4jikgtkPnjvMZtZp
r6n+ASK6maAiRHhcpKidaQudu0IDoKvZscU0yA68K/FcTIPzcht+Qvb7bT0M
oRcGBoFcxaNn28HXaMMowva410hQ0T6PbgOXROfNiu+PU4+KU02cX+zMkW9G
J9e6BvgIfGHqfuDc6XWq7sItCoqTuPz5zlRKIXx5uKSgWvG0Zj8hXgNOV31U
kkC7dDs4Fq/nlcTYKv45PLTak0TsTJZkJ99Oo2CawDDd0C6mq3T7BLGMEm3M
yj0Madyx5SXDj5pmUIQbKpNp1jI/NSSsVMAlBhLbhRWRIz6/deEYVRRFqbSV
e5pcIiE5miqDyYuErp6BZUkUnDOUbCpzTYk2zmwd+i+wlFiSfFpDON0oUnp3
osWICu4ObMNzWRrudAHWG9RHtssUQYmlp4Rzm4daLkf0/3oZNINBb3T0eTCl
XFljhwxucKRhaoWMqu0aT150EtHeF8IQMdnp2MeU+StJaKqxDGnVWD4hcN96
QYm9WSvvxcFHDQrSTmDSBf99C1T4uCLjfIri5PPGokCGQVPMHdeFRldvHaE0
aNR49Mhogf2UqbxLjYVLwPsiBIn+7aIEo8tmkl8/pEuY0jZ0FCOg6IMN4ZSy
93w4CgLJ2p/mEkU/H5nACReExrkRiU5sbbTLceAFRV14jek8POOyayVR7cRB
TR32cqfB+ezZ5dYN22vPeSksFr1dT1Nr8GOdbjYY60gD1kwyRfi4gX5pIYnC
QiXOt5hYAg2obOcKtk2oyzJE2HdXZEzLYaiIGU0wWhEBoJpD58SgBMNTxN3F
dmqcK5cxhVHwnanB05RYPq4nqmJpvh8Cc6knZB7YBw096RMlcUo1fdWShvEU
p8jjZHECdSASH1QFh1eH5dretmqQ8I5vCaGpiTqel8OhQU22GrpS2egUy4Tj
I15mcssFzrxtSHs/LHLb7VTvntlr/EKushJgvq+IPihURGdILff2rY/VpOiF
d0a9y5Yz5JTrK2jW95yOb8l9Rh6CeK+g1lFmIwY2zaXazflZ+RRBABs5r3z6
88LZkyZ0GCrqJuPte/XX3zzEK4F9JLXb8MChADjBuVGGVyEja8ShAK3eZUVC
JkL8SoqY7PvXQDcdZQzIA9FvphT7Kk+AdPADaTUN0v0+d/GKWa3NvD8O2rEb
1vdMXl/XZQ/nqPNC+oE/gu/PLYWsyBH49WDRFJx7bINMVC7xfw/A1gq8yn+Z
tk3XEGSNWwiIHsOMmfACRuQ4YdQBk/eV8FReEp7U5B0/5/f93VaMX6VkoCI+
hdqGmDjOkL+xmyYKaK7aNXAhFVJ053SLwdfE56KX94lPOmyyCenfWPFK5vLI
R8aQ1ZvNMWg1nAK4o+xIQCLP1vIhkrhECeqmWbwWqLfEoxWEMbnI0gMC9BPZ
Kd0JZLtM32p7PnNP1/CBuqnNMwvCIFiEt3nBpY4kuJZAQ94jvTEcDcTC6yRu
Dfj7a5pvsEfet8IxLGB4e/D2bI85062EUxTMo2prMIdVsbmJ0jbvn/7m1/No
0SFi9ebIGfmByK0hgTMYGdJiD9Xk1X5FizQZEtZm1u5OsZpd9blp87noSl20
Bfm1tSBhS3lSyYuJDFzmYcuxYe/+vrmHMwAxAVpSBS/J54jNFpL37tNclDGk
8XuOgLg1g+cnlDPOwsk5sYpLauTLD4WYkhn/Bj6Qv/r5eUMMuebgDhxbC/9H
Z43RkbPIAzfMvLiJGcHeAf5s6I+Nq+MPIJezPV1Pn4Q/fAqK2aAh16L+LRS2
nUFFkAtjRwP6hvVZJIBuiuPYdmvBZtGvEigCNs0k2H8b+VhD9B6ZmuKIfQrq
yk45mGixeQPnYofyK57L8rtuSDDqeSL8jJGnAyHI6hEXZ/wuaL1Qs8iMb2z7
wmprxM5v4/OgLmZD9KwsNjVyq8WV5P7r/ZDrmU2q3pu+4PfP/mab9vo7pqF9
DCHVdR8jNz8WULK5Qx5/Cop+rRU138B9ald5CYTpAANuUOaw0w7fFK2kD66v
3hhIApdzhfvhSTj5z+hZOD8F9bJXx1YxRyAr7ibaccEVj6a1ur/SqWqivDcS
QjOQXYl+szRyu5TUZiiBmBU0MiMrtwN9N0Gsu4JkN+NVEb+LpDK+uhvuQU7i
iNnv9sah568snbrt0SUtCxKZRS4mx94AnbmQsSugBxMnZpVbEobrfrqmny3p
1GCG4GG6OfNvLfivQjz8bOm845Yzs7SxqoeSMwGNMPa1H+kjo8iVFfBNcgpt
+gHWdJ0FUkljXcR8wwMHC8/NW2JsT5i9B+yqQPnF2OgO1lgy/XUkE4klFEyI
Til/8rpyOBOuEcXnZj5aIurtPM30g2Ki/7oZYujSF7DVfjNw3EY/jdaFCbjM
mxHCmtFAzlWY+G7QTgnX1C8qFzaDPRxm5NJcFxxBXlaCENmef4d7Vx41NUsc
7gydmK+mIeEfeUW1lxHhqrOLlmhchNCbwcAaOQH5SCtFXGBU/OjnXvae9QuA
bL881H/BPm4fFvJif7/ABwDPOZNZHLjtgqT4BYJcFtjdn14qzqenspL1mN2r
DBnEPFjAIyOJqDaqnFv3ZEiHHhXah4KxLxX7O3EJgevko/zOVKx/Fyt6W5MS
yGsXZ7KGLWUFAKAstWekYtln7TATX4sT+Ndlcd0jcaTt6+qRBhCJ+qsYFv2S
KXE6DwO1x3TLiUlE6Q+/L6SoNuh7gWw+WrM0FT51YKP282FW03BCByM4FLwk
ZKyxMuqEBhQ7K+KFz/wOp3N5csTpSV2HloD9l+R8dWI5SFPJsjuNC9LqB2GL
OXeSYWXyFHvgXB6dj0l6mTgMCMMTqBLPkmaxNeubmACPFuXqo7DNME9K586r
y2K5FDa/skx3KHRBlu1FuySgbsJtj6Q60gLNqeMrVhPY6TonqWzijKXwsf66
v5L49Bi/57UH7hXU6LH4REJN9YknNmuOAUyR2ZlkWBvtpGBEO/dmATfE6h4O
r21Z9/OaIgKr88wQcmCmT9DTMCP7fYKzWkL8N+lHJtYKnM1IJ/l12Z3JPll9
jaowFGee/PXApLcgrIO2Qz3WSVc5RxvctRvwhdGEuTmPJEWOY+O6RBfiiymt
r6COltE3C8ER3S04td0wg2Hky3YMa3uLquo4WaRLYlTja67N8HDtyXHkOwwt
/CwIh/BSqC3z6kiTCtM8Yl863JGXUcXJIgjJtHwWVBT3fW57QmlR23UchVnm
YjgfVpKiakHl4yT8ArnS3pLNaGlVKAo0sGfBkfYewlkA7R+rPkuHTfgzkDdN
iBhSMqwMf3ZModjhySCMdAC0eAMIElZqlAO9l7bvMe6lNPYQetyS49w4JBjK
A3WZNPV152Ubtqm3jeW9VHbKK0kgCpx0PY0tY4VulN1xXTthd07w5VJURA9S
mqZXlVaWfZeX7uJto4rx8TVI2N8sw4XR2e6TDq+P6CQ1LqpmWhvtRyPvM+dz
C6GRbXdf3KJ1YBeD0n1N6JcwXiQKUK8oxcLCCVqO/ZLCZlUz/FEVF+D/ExNc
z/HysGBWwez7N8wL+SxK1hB8xgsMKxmcSmEPP7zipn2dlce5DTiNAYSN8Enz
qcwPb5Dia45E8gASk7TNuQQEQoXJQ8m89a09po80tAkjhxDG3rYouTEPRoLo
tVwc06P2Pxhjw5trTs+szwGFv3lo9wkG42vW0qdiWOGtrBuOpI1NEnSBVuNF
Sc5uos68hx8pQnJ0TGRyizzRxz7OLj3PVUzMHY1Ze6Cv2TJQFMDudz9em3QZ
v964yW9P2+VjFP74CTVTxH574IE0KphQoN7jWUkuBALcE8sQxwcMDIvNUtJC
D3CtYNHwg83rucbsg3E+274xOu6PlG0PLIqMKxKsE3Haj5lco+kehQjvSWIU
bcR2aTW4udiaX0mVUJyuJrrrKwuaQgkGRlmughg+xHYHrHcug4HpUxqcOTdY
cZ53Clfv0lSN54/a2Y7VVgzBNRd28CaXUWwpNp7J2rdsUzV9+WpJoKbAYaag
FOTBQMZy+aZ0E4z0Zx0lSkiOwos0l8VJOCbvCCVrWg95ZUq95ifEWtpuzkRw
JznwusDsqAVkJpIWYmqmmUHzLbXXyd4fy+tekfmbFnOHVKoaYti2J/4adgfu
ti66P1ntPLZ+6vAJZhuD+/vQbkhLloD/nyuXdpEvTe9QxxUva+1bNVyQoB3X
bihdV9Jb9lT//3T5NZHrHhISg8w7p1rFuJs+BtRR91j57ayuD5Dbyak8q68v
3KHsg4al0ANHeV3A3IgaNkhjkRNn/to6m+SKnTAEQwsAkDFTPm7e13Fkenft
Xfy/W+WDeRt8CNO3aNo61kfkGG24goqQEc0dS8U3QZ1rD6NE88GXCdP+YHTc
UaloFoyQeSMjHuQdhwTzCo+lgjgJGddBc2nrw2kpQJAuCCM/RTtOtG7KGf5u
5l5KgbsQxA/HNp5nR4OCGijEgeNIaSJJuqfPbVhH4bHUbLjHiJKKDYNDAjFs
PLNIhfnSMkxpLA4H9IK3qtd62cM0esjwW7Ou2K2y4rDsGuf/BC2TsTwK9ohZ
vwWOPFd2HAspuxe7C821HRHmyvQTuQvkzcM5XJR7BCQ4c6WlsltDLqXM7mda
2nd8rCoUTKQWCjMnPai5jrddQKph6f9n5/9oPWDAGLz1ovAVS/G+g93ne2lD
Hm0Fkg2qrKGQ2MnqnbMSQBKu61w4S3gQSEkRft/zuqf66revFbInW+oOJu8V
977DDh1m/yuC8GhtOFBi97NDmv349H23N9Hj88f4DxQptIu8XAg6SCymk9Ls
DYTh8ObwlX4/Tyfn14tScXEkiorRcEkrqBM7xlUJtPhXIb3dg0y2BbHq6NEe
dAolRz/KDOmQLBdc42WO+VJdJQC6q1p690G7ZZ/GvlkPsgc2HNPdpoZDwsAO
4UxFX14Yi3uVTkuVAFnBoreyW27eT5j63aI0DHQHSDEJ/6L1J09cgXf56n8Q
Kz0pSVZnVy+smi9RcDas12k2S3xDwK66FtyTwIc+PKZqgEAL/G4odjxmujAp
cnS3511kkLwV1aCfIiUnsrGZdchUCwm8dr6kofQs1h7IuHOA+TlqBGQ1YiU8
+vupSyx31XSCrNXDMasAUDXYBJWRM5WhPoxL8Lb1eAbbMzYG/P29/uZoYHPU
hxqtMoZZV7L5gvyPc+eMmHuTZeDuEEKqGxmjNm+uSygzEwvv5CIapi+fA+Np
fAkKaBT08VfHB0Rcf1ifCo0ENG7P3owP87NAwEpojJHH7Fh9ZfvvJP+tZ3Ue
je2N6IF7/ahgEaheGPxJ5t1Aiqjy8H7t29N0qQq+z8G1LiIOCMl0RutmOG2J
O1o7j3yRR/Noji9AqqkN2CY84Osa+beAD9YdB2D374AFjqb3Fdm3RV8gBntP
oJZ12Y8DJP18KF+PF7A7KOoKJ5+C1KIFWGg093ZN0I5XcFdjFpuN4DKhoh3d
SyQTILeGaacWmx9eclO1nOxwzt2n4xeF3tu6Nzuji4zzc0VcE1wUKiZGua99
EDrzyx9HqaTrW+Wwh6Vs5SOG4SWWegFsuEQlDaD3hSLJz+JLVFEHAUxLrUSN
7BTNCdQrkrXC8mIUMQUBVnILUx8IpGTnk3obFhmJDajrCQIVTe3N3VXAwfXj
bLRHCsuGt6lpuRFYBrSSHAYybTdk2q8t1HXeDzfHJE8NUDhOtjfO5yw4R+FR
nWeIS+Cc2nTbA5mUGhDZZJRBJYWVec2MDlnktdWB8gf/v0/6s82/TVNqlqtN
Jy2yaNj9vaqWSzCkD7vm6i6HEsaD957CBvnj82f1jO+rqbGOR10PvlajKEPC
zf+Rz8hKlb0jgyWk6AD7GTnrGxZO8vzZ51I1u8OJT+H1cZ9Wpiicny6Iy6Qv
Dz5RcekrtlV8He6pXyKwtd+Ry5Ll2L3q2c+BEZyy3n8lo05ZzDFFch/ePqWb
l0W8szhsfgm3Hkt8m8mbHcCAxXq4AzHNZlGujZvfwydtFkskrtrp09U3iDUU
IHkjmWVWmGzAKwCN9ho8CZrY3APwCd3HsrQAkN9UjiE/JWwvZIpBUHel2KDM
CqgZevriy9XOcIjo9X47Ut5/k+S9IFgBeRMgR0OlNBieIfFZBxT5/0Nne3Nb
xD+UhQwOx2rLWBLAl5F0fmBumTEuTGGttcm9I/d5B10Rpv8uOVWfxpGHKcSf
FBbgxNj97HPVV9M1/HoDC/nIDGgRe+iWP9XRMbC5jloYwvFD0HOeNgF+iR2A
vqnqrmfjNJ+oIhT9LA5g5QnH7B1H6xim2ISrHTpN5Aga6llAOxLBCVdd8PHh
GGguM4qzmGES4eEpIOuzeiFBUE63cxJodlfahTxqxxSoimWx+j5lBjSuuTc9
R4knel0DKW7He7mRhjueHm4r5EPhUxbL4gIdznSUlLVpXkIjZeuFLm0eFypY
eq5gli9QQncOmYel5PLixeaN5THoVOyXz2Aws+NOFx1P9aMxChzXBnhG8/aj
T7X6Ud+lM7FuITZV1VdiYHkCQl+SYwgfVcqa5yuoDsGBxJqnxVrl5epBtceb
ztEWl/07Q9661h23ngxSSFWJzvj4WdJiyggwHdP8IwvT/hJguo/hu3ZfyM7n
69N2jZLCJT+r0Momfz7nPmr4EFPstDcXE+zUT3vV+p2GGX6rS3pM86NAb4WZ
VV6QcmLzwWyryhqy/Wjl7q4ZgRsCl7J3hd+5lCsX+/2jJW+A15r0KUIuTRlD
IsJFhaAstprfVY2PRT70bWX2nnzMkB0Qnmg5B0kl5DP1gKnSkQiksFo+sajq
TBYhewk60BaaqvTOaFx/UX2knEqluIJwCFW7Lt/3+cAS44vZZXE+qRMeDrEi
NZbidpt5yGcD9XTbOVeD38ncUlDljpwLD6cvfmLdMOBIZ/7zCPmQ+UTecJq7
cC6t59/UZSkECLdsuTpnTDoxDUNR3ZtskbZhcpF1qBxIePsBSbIMCwo3+n7h
lpgdll6vgaugjzNL1vAN0BDVrVkaitKzzpGQwJ6sJDnvpyJoXuwzQRXeZ+TS
+5qA8ct7qkx3ac4zw6eeN1UBjjiwK/Q6tVKGR8fgCZTr1j9DFUVRIrZy0QFs
uIvh9V4PV5t/D6UGVkBz7frZfRzCHM8SU3yhwZ3OgespjUHHCSJ3Q74Gyxe0
yKLN2bfqzAbAYBz8Q47f2TQAtic9wylr48KgoFWo6jZy4U8m8T21R7wtGvpP
av852fPlX1cyJjuooCJyVytYB8tQKuK1+uHtjlgxGuUAPnk4ygOu7JYGEnC+
8vUeD9vCjfhtHzOKws41CujpxilG9WGAsDu12APVM3EBtd0gGYoe8d3SuJrY
+nFDFap2mwzLPbSItTIV56sadwzxuLH9gghYXPk+oGnah8FbdSabWnSO2tdL
BCLz5eoG3nGOxu9h786PzDBdRJtkpcAEdQ3IT1aC5vtPIR8Q1aqTjWtjHTvw
05Mk1+QcG1uVAPObKBw5yHZm1Y5fL0OqHj2XGPmv7UMnwiSG7zvZshWqgde7
sYQODAefNFnVyUqOjErD4WdiJkPjccrq6FpiuYuQjhaidB/jd/rEOxstRuE7
R3zwUMFCiVaVuF/ftscumD33FwaLgy4pOBKTES/9Gg8mRMee4Dm4cjduqX7u
5CLYg4cg3y8vqRXBy8bdmxlz3y/nXcvCIJjieDIspGXye2fSrqratX/3jAYh
KXicoitjmt2vlu1ijWjBKUQ0XFQsZzFWlqGlm8iyk6C1kGrbq53Ex3UsJNXt
vGUBXw1hysjh99yCVmLSZAIvdv8SVZsvuXFYLqb3wLr7nXGnL0j31txqwlJa
H7neiPCtEHLwU8WduuSXoxu6juq7vpR1f5c51j6+3fddg83FYLYcBOEEuT3/
rNNBsqKMAUnRPeUY3+DVprgKXo28w0KxELP79+FEfWmPgrmyo4F8bfEvEpH3
dXP06bS5z/0HZ4SwM1i8N04YFC+iNJMuEQwMra5FS+mR/MTaqYK8FQfwhPX6
wvkOT6UH6HVUI6XlR0eqyFJWg+mONR9MKd2G4WhWaMwD50ZKdey7yFVqCCCZ
7gJn2GY/CtjOeXqMhMN39O5x3jvRejJTgFEJxpwvmL4BE4yFs7DCkSzK5+7o
EWgOwT9oKET0Qg/y2AXS5uBQcwS25uk7osBv5xBHm22Be9bzyVPh1M/ZyNsO
BSgivnd/2JJlOKdX1cGaOznEutrOv8aHOnWonNqawbCfjTWLB9vK67oD3UNx
BlOTP0KY8gy+PEGiZqf/aIEJG6GBGXY1SQXG/VQMoKFlhtAKOMvYldqpEwd1
0Z2IUPryEF396dGcaXsbTFEnWQ+DiooIXLj02Smr6mD0fTrPizPezw/jGy0H
TYsSVcDS3WhTJIYq6DlpDmgoGW8/B95DedJPbhgFiDjPAwbBWBCXwRiWTiuY
zHWD96u7z2V/NfVxOivN9uMlPx/i+jOUF0oZEBAOgrbQl78WyWxLU7FOXjkR
ctdkOf5dEZk6emR0pKhiJgesbopSIpu/JuHUTQKH66op0CM3gEJiXcphTnHm
qgq8Uc0+JFgwesn3tSOkae9a1dOaKyxUEmlcs59yHACZSRmXe4glauOSHUC9
ddFGRz3EkLp65ZaYU+jYKaRTT6jw7k4tU9DpwMj8j+4tHs711Hw4nio4MnIT
RGV5NKQezoMdjmdn6z5w6FZ4mh9YxoAOcX3iNd+rQzZ2SAm2wx0pQ2pciWyy
KsuUsBsVNjslmXJAtRXQalh58Fw8Sv3V8R+D+nNZAzV3+u/IRxx59yIB5Z3s
18Du5vwIY66DvGgAI3Z1THxy61UQh7b/7H+mqZ0p6hCowcNdWMtLYAotRsUe
d/83A9jMA+t16lJUPLNmFGFqgv2J1OsEv97heRJitnfwuH0wsMmq9Mi3bp1E
3zQGFyelknr9XWaktxeueazNg38lsMwBoKDu7PzIUFKpC1r2sPdcsN8mfy2N
PubPerdD/9ppUML0ax4d3QM1A0wKzX+q7b6qIvZGCdjQ+8+NYMb9rn3J0X+e
vVSgDiiKLqjX57CWgOff4vriXS0sRg3TJOvFAmDUt2z7NQvAUu7VJ2zDPuuS
yvxx8nQ0Y+YxValni/qS1vM3Ncrglk98IHQjx3QT6DWKRsRCDHtPN+D1CP57
waPBjtK+9bRsvDYx+dKAkmvoRFuKhpipCUI/0V3fulNzaWIMaqIQ/Af/pbou
6AB8nnVlbvVym+aPuQqljpczrP6bsAT7FPPqGOzxn6a1+zZ5VcFsq1+5w4bd
z7jWedRI2QxQ2N6RmYtTopfSN2RIrcy+PrCE90cwGySg0/QRU6YFwIIXup2y
FzM15bQY78IPj4S4wdkcKMMNwDm1JgDSBbmXvTr5H3yJ9vaJ4M6uytAJjcuJ
6rrx3bw94mZqzjHJwqIcqDd5lMgYc8Q9GLUUm4/KhZdPn6lIZK5QPJl20t7N
8r8LdsPxVmrbtU8dXcdHNPvKBbb0GJMSnWb34Iw7FRJ2ZXKiVHou6GmewoKq
Opn3x8gK0mRN9WnlqJEiJMuoxpR565paFAx0RFo1b/UkC/6LFsN8XNevvRQo
MKLV9txKRcWzaVIkyaplurQQ5va2Bqymq20rZFdS64ox11oLSEa9L7fNblPA
gxgiAmvwIWB6bKwBTo5J6N0v57q8A6x1zJlMfRIcUzSXDJWqEDJFA44w4bT4
YNMVqk3oeVXZzJLrdhPN1cmG9XD1FkQSk8Flz2YL5Sv5Bzb0idORlAWAFt3Z
K3/BRrwjBkGnTZv2/qwEX+Vk74RqAMakx3fKbhyAZiAvPQB4NB6HndPytKKi
IYPt2TzVoaIGqHoyrlQnefTueEHqGw9VyxxdBr6/7EnOncWSEIWQ3KkwcktX
R+C+4RilHIWANWrE/Q6I75RsLXdd70akSVjnZMk8CXdEPH5+R3uguMa5RRWt
gf5JnON/0s+eimIbXdC1+IC6OM53DPO4pXyJYWItpK9o1yYGyJiy+hXO28gn
my/aUkM+nnPfrE1bQmJyZANZqIvoRg8SuM4MkyvlfDrGyUsaAMHwWSxHC2qO
WGAkNMo3z8k6KLOXyHgSaDgGRBKkHSeLI9Irxal03Y0E6knIvawKyk4YW8TF
uydnOqeZgMiqb5t0gsXrzTNtivbF9OCya2hMf8/2uBPdvgJeTr7A2of9Sh7Z
qTxmxaRvsM7dou17I87iEE6uN9+u4+vobz+BaT8ce0kCSShXoLfRDxragtU8
CLTtCwMsiCjIHP3UStWtmxR8CaSG0ME4eRa1fuSXvXfYXJVU9BJ8dpceaPdD
+HhvXSiyE++r3mXCRY9VUoVvIU03hQ+83k3M9FD8CW4DF8Q0kX04RV6sTFsz
iW5uaWcHD3xhYzj8lbGKkTvekxUcNaICGThJYUmsuup3llepsikiaC9l7Pqe
VANSg7wJqVWo5YN3+ut6CaK8p5Zu2dqkKSpj2UovOF2JNGRjfEF/CL7w1266
d283zkcCAFmq9V2B3TXELFBf8YLO5TT4VbFS4KcIJrhu6+ESgB9plbAtexl7
5HjXtV4MVBgekt1AX/hnByRlxRNvMDGUGqdGN3JnThSQsNnXezRqr19FuThB
Z5I/bgVHW1+bdrrswOv5n3sbxjNfnkeiptCUBvnymR2+kIE5QlF2dTuQRc+u
0/3Pk9776shN7KDjXe6IgceKnIGCdJ6A+0iRNjqoDE9IB0kubvm0WxxnlF/8
V+Vbp87pnQcSg+kJZ4e8JJEs3Mrk6dqFT24SrIUV5WbGor5jur1pg6VxDP+b
VPzm234q6RW7+qnuDu0VLmltK1KhqznirFL8bSKuTdRy0vgMG7ZYIi6dTg94
cg6/ZzI7KJxk43NegHx/Zdc9iEcVX7ia3lRgRFugrpXA/EHGKo/bgL4YVQSD
ub56QxNwmb/uXTtNMFPGY+gW4HioRsyw4YgjBeneCiavfA0bj9LD1++NXr1g
V06mZbUbQk4+RJkA6dTn+L7TFhU9D2RVSY7wU7RbGKchhiIWE7NH+Te2PkMp
gH2SU1u+YKr28o9lmAdNok3PalAFmwwOXJ5/1e94JnvfFzWDeZ5fSJ+fSPaF
kx6DTGAO6AVo+fBhxdiBShes3mV1sjJtC+Lf0zAYTx1EDTCQcRToOv+kGWzs
CdRFxkEEAksbvpuE7KvmwmxcIACDJ+dfSmlRpRH7j1ke+FIMZNSmgfWu8bEs
plaqTW9IkP57UxEobM3aOoINbEduaUKb+6NpsabhFY8Ha2l/cqiuLP4z6FCi
+KcUNe4OgF/qtlfpVQ+oLig50QurMwGZChjJzNN7dCrpBzvjmmspnLNgz79y
ZgVUnVawTLwWs5+XZna1rOx/OVI+GZfhfl4r2WX0C5eK/k3FLRfBHKE+Pf4B
6bLwjRrVev3wpAPt1UFvL/ThDocoxh7r7U1IrlMk2wbY/rUajEgH4bfm7s+9
0oXCwUBNnL3GFNHP8JTKDVXL5IqmayO7RzMSeA2ZPFyt3hpCXpba5Ah/iPdN
rrBdfiN0M+eo2WGdDJwDKD1U0UkZqL/S9XDKATMR+vAF062rDQXQmSr6jvy/
TR5IGMwToeRgllT5f0yoQOHNUcAMsvgygeOMjhmj/8ddohhuUeR/YlvVH+HI
RU6rmi78ETeuUHYsSFltO9pNSiba8NRtverO3eHcl8Ac5HQIZ8HC+hdtYHXF
9h9yQGZ6tNTBxTu4rfzzVmO72mGtKfWabVR1/3pvkIwdI3Ay2M9WBSmoPSXL
1WvX11GSsn6+uRTinxwsMA+gVRI5ujUysHIup0cqqMHhRplOY97Gk2CwfGkJ
3tpDiUlAATSodYfZMVtJAg7//PI7XOGwo16o0L26zRtrh4wigKgl494jspC9
2frwP3PrKC9SKheIT6x8gGTLryWeRBfwLIFObEWxb/FkALzLSPjvPuppShi0
M94KjprF8AF3N26AV5R7Qo4x6QuCAVOr+sNt3kqeS5PKEsV4mxXqOCOtFEJr
TVG/m45ksbPKZgqRVSEYPJ72xWSTCvhca/yl+cgtnxaSj9KXVKEbjc/ZDHT5
KoCzh3Yl6zaPxq+9Jb4aUcOArFi7WGowP4lWT2ikvTFqB/PcLvmf5mKZtVH9
GTPCWhVBVj5YSTGa6hvd09pZ3VBsvUsjO5mcXpGxLdYXUzU/eKkzQCYy8ZFU
GSYbEm2j9b1dNAoS+nSosci3HJhIu+ViINPqCLgcwgl+fteemmUK0Ar3t2qV
SQEOxeg/d+UZsQBzX69uE8Pyb0m60oSfKVZSZKT5bokAyJvfQhR5RfZJZpFS
5hewjjkt875hBO4ppoEFBGFYCht/3TO3UlRedBYWYZ/kd62jsL63jBPE7pHQ
11nHvDz+TaBCnKe10foNXPwp5FVing+K2DQKLLWrG745zlNp4xYD3mmbX4TG
Td26NSRVj+jUf26/rlWe9fenMX9rjebGnlS2RGOLMDpUHuJeoLrrKRSw4PVu
6Tv8trHDiVUAiLs8UEAx+qRaxWltaRYP9ofp6w8Fxli9oOM+3Yh4htOCHFq4
CVT9RczOYzcyQiCwVsHJnpKLk7hbj+CceDIESCvojltjz1p5CAY/JXSEC19u
d0BWNiSu/LDsDzFkz1ocKubfafCFkiS4yMv58RvNe3aenW1oxlrXbQIRCXw7
3pv8HNY0UiZyRHkvfErClH1QjpeBmQ7s8dD1mz+mmz6OIWcROFOWsQsfEtyu
PwP2bLDoIf9O5jQgZTyNiGh3YhvOwz8kchQBkg2r0sracFj8lrvkunwyOxU7
GEDW8ar2byXdnvFkHDBmveGjS/MiqU+Y4m1YgTJgdGmmn4ZqonE+1SUtFZWD
sfIUxAr3VTdBS+VnRWEDweYO8rslSYJXuHYIa/68/kbHcXQUyiH32Xsrqn9M
4qGyia1RUAW4FlyVYqRtmDmP9TC1XNvKZoQsnLRZwiHyNqaBlXIqEXdbqdCz
X8W6mJzgkEjIZV/THxghs7WyecihyGYGPKAPmNajrDCmHKZldNH7j/PrLJmV
LKPupsR6Im6KeH1VVlO0WOZgkuzDoaaW0YprvJGwzZ2RLFvhZVcPFIIC2P2z
Y9ak5GewFd11+wdr07qrT59R/D6ZlFPjNkHlIh8H8tn5Bzayt+r+BZRtvD4f
gnL/ChBUC+MEK0egXdfxyXWXh37HgunESWOfepZJzbvEVHDudlgWGya+TgWN
4wVtUTC8As081wfj9u2xD46foNruOHTy2yMhAacWW+cQ05xbmLm/piNMqk/b
u8knOX3IHElWFm2VllvkfNo5nI+nzjyl5TC9iW81PK+Zf/KWTckNGxMp3VHP
XBOQxX4RhSeq7dkMqhIIaTAXdy8VZ3lyqq5PA3Bl9OpkbvDBAnURsNX1aXZy
Nkeu/tY41LxYotiuSkjVS8K9hQySX/IX6d2H2LnCukm5VAjEGvMu8dqXillr
QlA1K2620DJZPHOmEvgANuTmwPf3rV+BZckRXGk86xCAri6Y6gwIej51liA4
+TxhYrfu+M8spZtrZuUOnAfkNGlORpuWWnQmh6wJBwLrkBJ4mcEqaNCn3Jm4
75PifEXrEr5W0dhzQtRdey8W7cTQqFDRpx7k/0WM+M0MPJYIFCfhSqyBcHQu
h1U3XLH9zYnnDsUVyZTZpSO1YxXSJ90xa9c1uP89SY+MRcnLXywXJujHNTV1
5PZQy6jwWTzG2y/Wn0DNDNNrUpUblipAdCsVPUhbBHUhhSMY5V3jiBEcJIoj
VNZQ1l9+jAwzYkXlOSrTFOGFdn2/AKP0xlwGnNutUs+1O6PP44HjBxQRzS59
R1QnQw6QR16oFq0RYN+HeYn1pQXTLfE+Aq731DrMD5DNwv1Z5vLXMhSQIwoQ
e4o5Yau/+U3LweIvrO4kkXuMZkVbY2uKfBGLvTz5/Fk6sTUf8SdQ052WXLIs
7yppDf8TyLi7DI1AxlONpu5ptBNEY+19mE+s5Cn3tZlrA1sOtkIwQSqEci/A
0jexvdEOUzrMur5TdnP2E/MAu3gt61HeOtgfcnKJlQ6hUAIsO9eOcqLVyv3/
evGx3gzHoxQPh38Ta9jCPIPEBJuVjgrSh2kn9soZXlQn0wwHNo3i9g1SC+3w
wSyrSazCRP5Kov+S0oM8fpUPtsAeqfVUS/qqY2B53BRn5jSBUsb4fwxHF310
gfYZS/dkUz4fDmjTKnbOiQQySHFFwBUNk1zTBfaZqApxqwLuSL5DmQ465Gcp
fQcBPdT2Y2Qe8DH7a9bEEQUROkkzARiNYOfrvG6KYSm9N5nBxlHRAvy5RH3L
rENWSSz+MCK/IVWPoN4/SVEF3f6DbNHxXEyXODpdZhcE/rQUnk+waGs/Wa3h
r9YDA5NETpqFxlVx26loMddXBmtUNAC3tKjFLbvDEpaB+O3JSqVPvhULi4jy
W+NAxbg7hUEuofBzdBoukIbsELiSXiVE5lGDYtIZ/Fu1+mWR7Aq0oGDrvhih
86Cs0qe5ByJs95d8Ie6caePhCyxj703BzRMKD1A40PCxLvHRjvxkqb1FzV8P
avznupH6sLfhz5NJYCGmjR5tysybit3T727S1RbyViSvYWMixZbsgADN4A0D
3dWnp1sYmhvjUSXOtxjDc/TZvIj1wZjb6UzCkPTkVBj8mZ1oIOU22vS2Y48E
3QAcbNpRbQxX9TjzXdzh2gtw1Hrrb7ZtV+uM2BmG/awwekQ3EKExCcCUN6cp
D88r+ej+Joj4MbDJ2r43CIv7ij8lxEi3Y9StcxFgVFs7JJkohxGnFlw2JYsK
7fYc1xes3E+RNcW295JUaz4y7jePGTw/ylv8K90QkvcbsJBIY48K5CCJhPJl
O2bGfZPmWEMiHyO2sy/FsbRZ86CnufwsBA8BsvnG2jNuEvcys/HZe1+hycAa
8i08jAq9WNo1uYlPcZNEqSLQDBETfWJNQafZU2ISXvIh9COGdzs+lqsDL95k
eLFUY8X3bhg2IyL8R8ywQxZC5v65kgumwPjuzYZ4xeD+MNOb/5B6cTjluOBA
gcWPx5fn+IWa9ZWJK3pn8Fi6zytYJjCQ4wLRXN9JgrKcso8PMHt13y8vYHWH
kFIFJJi4RI3F2yWi1d8UA7b5ZmVpzgt9/nivxGYNsKvBJm52vLjnGqk5K1Nf
sGG9O5TepGL9SJDyIAkrKaHrgyTGLSZZ8Tq/tknq481d3OWV9csCBOCyxeXO
UX4MrrzFOrXkEngNhxx7+aLNlXm3zYKEnu1odrKRJuq914ZJgG8CFTKHJv7w
jARRZiYz8KFoQSr58v4iKUPO5zms3HZzMIsrfPwR0vj1ncv1d8ikmwBmdmwK
bvyZWES5ysqFwYayAuRJ537EByFPRTocjPiok/jGsO/3JJv+tRv+dFln/4dD
q3aahX6n3Gg3yLedbRLFvBHRiMmpJ1NEmPUhWinPVyh61dDEt8kh7gQqkb/R
RDWDE5xkHFQbpxSfMnrk8J8gmMrLULoHvWQUwE0A1SLoBM0C9ZJyvRTanr9c
rQhpqpilCJ8egdnUKnL+3y134B7f0iCDLbEI7WrkHdC0j036t1PRf77a0ixX
Qly/nfEKUHInpcGsARoIvq1ckkbpTw5gWhE506+JAkGt7GuReemqY3NXNAYa
lafyqbdE03KTCGNz5N74tvcUUekLo0jevaJTHQ6jW9gDruxq11uaK5xBF9l+
D+OsfzYKvJEldVylS8QYLtMZXSk2wh4kaRpbONc3XTu6fZkBJ8ElOdW0cMkd
GCLGojmm3157SIUNpfgMI+B3dq3KjLJi2dGDbHKB8wHYi/bEzEgPFYn9pGGH
6OHek0gP3xDDA+i5rEAB1kVDTrzRDSqcZ87YBDLJ4xkn387VSz4H8v5mOcBL
wocw0JoZttXZ4MDdhlikWeNEkYDdeAV2zIyU4xOvQkXR2QysvYg7ls2WXN6O
trCuNSKp//ldKpoN458UIpcTB+5WUequ6U51ZQF1BSq4eUbwtGb3FU6sM1B2
fAtZcDVBwUP8nW+lX0EVzaytJUx31yotnbUqsJAEGJXmeEIV8W5g0Io8SsGV
hVs7CXq0py1euZULR8BQ4Y4cu0VaVMqg+c1VvodS6EMnaK8M9/fg7sykfSwU
AtG3F/KdU59NJok9IggkWWDiZNSCR81OtbB+kY5KaFyfbTd/sts7jWnDahh4
S6KYoNCb6AENvqKlBhgEWQAixKhXKWK3ojzyCl4pRLF0KaKiu1sgaaZUP4sJ
t3vSYSr4q7Bz3wigVFhJgZgm29c14qWD63GxO5JPdTDJbJ/JFsLjQgqDwvwX
J3TW3ZpkZOEsxwzijS/IYo0w1rIxIO6cuUTaGNYkl/WEUF90plX9aE+Eu03q
cu6mF99kOpazFP0rsTCwvGoFBiEKEH+45N13ZqsmUiqI+K+Cgd9DRKqliDM3
U0L+pLI0d8WVL2W2A6rzKQBjTVREKS52xgPCbEyXEI2DkKUBpLN92aq0GJee
KFo4WOURnkrBu341K92AuThdjcf6YalM+bLiltpScCweJz1rDlok8vOiBMZF
nepY3/+LiASqc1l7CGisJnIutgPBdN46rnLL1IIhx68dEhxeeurVchecRFu/
9qvtG7J9ok3AAZS8JKIgQGVEgfpWOwhp6DeZLPxjQMkXp3jmwA6pYPDy65uz
O2bue3VjwjGcMky1PhKvwBrQ22WchmnMohxyh6BkVjkIFWBUR0i2htYU836L
QCnbVmZeWFzW+eZdsWrMo5SmvLBSIbqF1a9B8U2cQLm6PDUrHNwkhZVQ+pJn
Qa/n/tX2xIdgr/ZlIhkOmbO3wwo0yyqk59K1FSkSMfgfaSY9rxdlbVTWr/y3
rKfJnhecJow9ApOVwBu6xiBjnJ+aYl2mtYVLXk9Cjy7i15Afg7ypfzWFilp8
65FahecZv8V5PBayCG5sH4mCccZkUid3HE30RJFdA0nbh96vGxkDTIUMSRpc
f5nRTA8m+mCtxtt6fLuZiXkqHSwbkWPbTOkYEOT5Nad7Jh0BO6ZQyIgnZJxB
OmDR2gFeF9KV6HIO5u75gFraGccJodhq/EhRlZnf6TOm4VjBCyz2a1HFDNrV
osuyhGl2c663rHzMd4oDhcyZwIWkBC/OY7fbwjv1j2zMrBqUCPU4e4/RTd/1
tu3tFTXOC+kaPoTBmqON5qTKAa4dTGB7wY9SgkzrHUjyuUJEqLVx9mmFyaQC
UFmHtnvBG18D/g+9uPnldd7RvPNVYr3gfuF5L8rrmzX/pmIx6JiMlEyvH4V1
sQTi/ZqL+DNG2XeSmOkfCNJbsALQ7N9tAyOIWOX8nIp+kBaLXj8l/qu/z7xh
+ofDszV/333YZkuWGL7+s1m2CKL2jkyG4HaKvuqKd+OJ3kevO+4J/NubsYuS
WFoHEsQSRBE7I0iYpB/ToaspuvvbRTskK/I9TgRtcs0HyY94MlAIxzFjybvp
THrUAfKAgRc/UnU0piWWclB4K7M9AvCk+JwiqtKrg+7lT9w5Qp5o8JqT4AmD
LQtesBGi0HqTZBLkeFwj+2/y6w9DBXdWGXNYSpKn4lk+T4iA0YKEI/sHQ4RC
dPMlFthN2hWHkUbdl/flsRR+bdb68tCgb9rr1VuPFsuwth7Ni50m7j+y9/p1
am/7q8SmrgTxVme7jaqxPmXWkRK/r9CzpR6g4sMSpDP6VWNxjYLf05q0TiTC
/bmKv5DGw/GCOy4RZbOCcpIEhlTGRf56T9Rqf8TltDhOLukLGGWd7liXzjae
Ke/kpdN53uyec/l0QoBjTAM2euTFjJ9HZUCGIJrzBpAW3WDa2fSC7Pk2bIQ4
Jb474lkmmdNVE8oITAAiEbhjLdSCAeuOHZjDQaYRDt+Qu9dIT2n0qinQUeFW
vTLpc2o4v92DrCWoAck2rQA7SxB8pEmNS11JKv7nDrPfRVSZ4+b7gE0WPgA3
ckId0zTnVFL6/3nbPYNnMQgcdFNHne7pMnODR3TKZX06WCHUEE22NwcRyOJe
Oh8oGaZIYeJDPwVwoP4q8UyE0rZ/BfNF/Y7xdkJOyIclIFMBTmtZuOtIp7Jy
lSBmbKpuB7QraTB1cB4KGkwsZ4aqFliy+rPIJnpTmBvswCakXhNGe+M/bfFa
xkmsIie2UKT1cEHGmnoJYPN68M9MqgcJWYAfuB7hUdVk+IEo0PVyHhqWhlRV
/RNQG83MNS0iMwo3aJ7l5ncwE6u8aGwRvKJbCyn/9qlEL2DZEx8N+mYSKFfr
6Pxyts2Ecv1F5wWTbR8pCRFDC3EX0ijfuwnRYoA2sqOtl+zBa/j8J9sJjR7A
3Z4llDxO6q1WRj/IiEBwMPyJOnqTkmwibJ2qV5M54+Nwako/02YLX0RUt6V8
PwMSCeGtjVykhztV897TToj6h4VyBkUVIm6Tmkt3LWbUoddguugUmKKaMoOL
2tCMeBW3GQc2POoKGfWtEi6qgdPZZaMKr0BwRrIaL13sl5wM/9KlKtWP4D6G
F07O+JkB24liDDVMMmEnL8iM8Jm3Q3d3xk/Ff3mqconRMG4rIGGnw88dPGR5
FLESd3UGtfkrpGgIRGjOaNCdmDSVk3jtWhr0YkEqs5ER68OFYK66arAQ1E1V
iXHy5SE6Duy3KdKsWiNA3SiRYyjnlKSTC3g/cYB9TUhYHXfF1n9ZQeJhM/Gi
xkAUZgaaRNhEWVtTkDNKVwWtbXjzBuXMV6AzXMelC9cA0L2jhBIFH1e5s5Zw
7Xozvb0fX4ylDEvXWMZjo0YPHrvTmGzAEeo//ocqkn2c7RLOFYlx9O4GQLkR
A9K68LiWjHinAeuxy62aM9Crme5iSXASRojmdQzJxXaPlGayz7HnGWuhnFYS
O8+gq4BjFazopV9s1yq79ns6aVu5P1ZSXJLhuhDIWmWs5XwGlv7vpST4KaTV
YUceQHqZL5dna64RTVKlXPA4G/fAk7IzOIRSxQBQ/KV9BD3ZkFIceA46xnVF
FIqkEyVr7nQ55a4Q4kgnkIfhFmozKfaHI3NC78LbxhWDaKgA/aH+kQefd507
soysl8ctw3SVCm6pz6pLEBw4riAwvAYkml8VfrPD2e+iZQ+5wiHiwIvDMYpZ
1csjaxMB4JPxRbGlvOWlyZx3EuANuxcVEgL3oMqCFjCOqy8BPWKlbQp7rXgZ
4t7AJKlnoJ5YHeKY81ffYlrSTsuN5cPE91pP9oWfGsnFYQ7ZQ7nlpQznjGIh
LojPMx4I+74REqcG3sIODFimyeMtWSJ3xuAfFv/lX6VxY1AY+rU/GzqZfNYZ
LIpkkSqPykS97LriRGSE72OMl7J4ymbTbbn/RmnT0ryYmO3wxMfLTRvNFGee
uBFbTrsPJ/zn/GL9fq5SxyXbC6bfF+VBsk4UlDjDIk/FX6JQ2r9dz4aSQW/O
F8QkdB0Ktp2AKxafjcjLbvQiDmCFkS1WPW2Q5QbLiQ60fkHgLF8ppuez37KF
LOtB86hApdsUFExftqJbGskd3dozC5GhgooIk4AEjyu5kV2zSW0By0f+BBVK
v8nT0oH8oF2S93gMnnQP/TXtoWKzPdu7Hxh3D4Lj3ytxr4RShvSRXAnj7kKY
pUas3QrE4WXsfeuwZYLIKaUy1hncfkTrsi2SHQfJVJZ1V9RoFRumgjOybGDb
gv0J6MKtEDBq2Qsp502cL5yJ6Trfn+bW0JKY4vJEmpbzZqD//szT05yt3Qca
mr325dETiONlayPTj06tXzQ4qcyWPnK3S4S6QMY2+Z7LLX+Yj2qfJI/L7cJ5
bHx7/pIId6nUFiEjzbqXqBMHzXbTAGJtfI6OsLIUTtl56ctLDzHAY6GZYGuy
gDqZ2Q4CQZr/awleTI8G6mQ9QOOJZX/YXJ11pCy209e9thChBSFo3gSnMCsN
Dm6gu9VZk4Yn4RQLm9MVLJljvttn4OO12MqsM/mgLQccsohRRUK3hxZuAwh4
Joyetg358d/P7RJZG+j/bKrQuCZidQGp1+DUos7REavrY0nrflj4kONacDVp
mSeVHwZlekWjng+aseACjo7EvvfR9ZfvBZCB7vEd8uqH75PNTN4tLOGw7b6D
PE2yD1P4nH0yKJZ5wy7aGTYzqSFCw4dRaDE978mVco44U9zo4prcPEM0EuIQ
1KN7CIqqyQnE8Zvw/joqeQ5oqdYdEbVzGZrYPPEj1430L1qBZQ00sB7Up62Z
mXeWr4riYVO9FMi2t26DUOs9yInBR3CW81CEpEIKmMPaOznGVT7Hmiokana2
bCnr5VCufG4Nz6SXvuVOMEIjw6gdTqo1jb7R2fJNIuX31k6xUa5gBYPXHpaw
csKLrN9jmAQYKY/df713mAFaE21IPkFRxXSRfReIj8KcQ6sbJgFt0HZ5EdVu
POaPzkwDl5pjkjxuON3ZY6xDZGizWCt22c+gCt+a07pbF/Vamj0b7/rbzNdw
mhH/KCjvv+jyxWnbCNl6HMxWKfrdSYZ4FUbP+a/TuinBf/lFqUBTeWzxi4vw
2oFAM+hsEVCwJnDQE+E7bLEEavW3IFjZHpPIqL/dyLNNpq6npjEv/JGFfj9Z
LkTnyyJYuhWWQwzYT/pcMLcyMvQfi5SaNogOYnttMoN0L0WX9X72S8OvcK4f
7qR3C40i2SdWUEOjzMaLA+yMMNcBx6fL4ZqIfSgbIeRpo2Wmp9KvL4/6Hqy6
bMmtl2FBZsFXOxM+NI3zqt6fynAA6tHx/aZK4xGTE+k+jGmcHly4NxfJ/qc2
YEFwMn/ArTu0ltnLW+r2YmLD2PGtrPFhf87fNxkix5XfrKLP09oVg6VRTCqV
jqXdPb35Nk/zHfFHy87qvh3GzqruJoEFlMb1qIey+64pbP62szufMUkH2CDS
QxT94D/qT2yJqwcJGDoj1wuJw9svt/ty63gEzvihsId0xLhjnDv6EE5CHPKi
QQ6j2+p8V4shV+y77vQr0T21r6OtpaLCuGhd9+aAq1PYRtD/GFBbKOP1MY25
G1rjhlIrSImhwEqAR+xI9DS39WB7ZtJJM5FO8g4TmZTj3mm9a2a2rb/63Hiy
OrGTzMivZEcyNBvZn2EmXoN3LrxfJWgBn7KEDq9b7Z/JmzIfNHcHTLGNuzgS
VpNBTI0BfHVxh28bjsHlBJoY03ZFPLHI3FqE1esfalczNBRMZUahl7CGvBMv
maEgQr6ZAKqMvCut1/0SQynJAYNNwMb6KWnDOYNUHshZodm/vjaNSQzevb8a
XQ4oMgyKAQnzx6pvBIWtMROCs21KHgtG4ZtxwOu9r90MV+SLZ0aOa5mX7dwE
zbd1ez45rf1Db5r0JKe6WDiaX0bSxz/j6nzh9gFVWqt/m5iWUCEhG2/07b+5
QMl+dUGTIs/8dfIFObtWd8pkuAqndxtP8m9L3//7rFTQh/iJ/C24Xrgp1Xfz
h3Q4reXVrpeGl+Gsun5+j50JWqp+//RgguFeeTcAX6b8JgOrDpwjt/tZqw0C
7/y8chuHJzpwrPDjIma+u6IwId+dg7l0baBvheNKqOGVsoe6OVD4L7UnIAWN
l748nLN0ZJLmDcS3bvrKEX1cav9ShqjBbf263yJgEudodcUmnqNyg+w+kU8n
97YL3bxiHjnIfKQQ4RFJZVdlPSbuKYPCCBNQsqAxKC37U0F2wZeuLzsM68gP
qgLMxUlL+2y4GRa8jtvovMQK6tm33qs+tLsRFIVHbYXF9cPp0FZzIxNVon+K
Gwu9tDUODaQ1FvWfJx8o5k3isyLmSMJlDEDdrWiNGlkB94TiLxstpHMyKr23
wDAojiDiBWz0imm7R3X4Fk6xkEmbvIg70ON73liq+d6QmqK31NxZKd8b2O54
Z8JPJ0vQgHytDN3OrrUYTuoyicPRzUPJHd3LhwStzHf0gGZ6V6H6aV5Gx4dB
C3Tp1RuVEIfxw4HEjPhGoSs7izm/eBqlVu6t2LSwP76obrrLtf3TxRwXfGoi
vIOPxigyKsQ1bOJjBqK5hS1gLw9JNisb66NO2+MRi8hRoFWy/GDBFOPM43M/
neDkAY0Wwk9CaUKUr3ToJtv6xlnQgtaTsO1RqqbTbtH4IzPr5Yucd0lJqdzc
hsnDJ7Ll/ttywV3IHgbor8iSOcQYOeX8hK5WpXVZYWMnuyh4/UmRN86Uru5u
Zy0AgnKONZI3hiWmb2AbtjzPqFT00gx3597hWKW4gwShqI20p8b1nqQ9zvEC
3uOXX99oP7GqRpPEIkJzmZw77lPfy+iSneNa80xi63Z71xngZjmgxD8fNXt9
qciO/n7ixmrRij/Vc8NsQUMVaHieKYqfKfLSCjL4Gi4G9+PSxvRU+9a1psSa
7i95ZPLYKwoxw6qiDYhWw39w47+7dRQGhlgaVLbFeDwzjBiXyo9N/Ejt54Lx
0sy076dZ8eQQsLp72uP4JW1Y57BBl70ARuj0MNQroJ0tL24M7v8wngrDu/OI
I2N+G/ogOYtQsz9fBK9scmaz8LqtBm2bYNmoK95r1fXbgWh1Bzz8yMSkOiPk
lt5rhYoXP8vV/WNlyshUVynZoFWmi3Eeh1msYDpXYetPqWNnQrVHABWZWkGM
pSI/xpTIO8YPFME78ZFQa4xsBJS+CWEQcNfVgAU9WdACE2twRw2RnwLDudp2
fq1DpY/lixXjc1V8RhQqjIZg9qTS9gmgNc08aRWhy+aET8eOxyLY2w8gBXRz
7IdKfOc2ypt81jhQMc3aQMluVuq0H/LttQE4xyclpu5EsU6G7JwBryxWwVQm
aq/X0PItVULrjwb8PUEvGYht97Lzmyay/95DljA8fi+u1EyTw/LSPR9f8Z5p
DzZeqostiBc1BmxpREqqJRuQmjG4an2BFFsSQOTy7T4/BP9Mlr1Ihkusp71a
IbNQ4OP/egu1rln8QDTr1HOU7iBESBJw4uXw1Z7UUKE4DsWhiV7kSXx1HNH3
DQ/mne8AugxuNFeWrgVvFGCpUg8tocd2YJeofmIQXghxbaZjxowfvBdj+rp0
+fFADJweuYB97as/QrldQh81irJy8qwRD9SylPn2e+CpzeLss4husrnXBeEN
SGpkzjU1XkbOtdAKrUbx2ttVDTmvjr/LhybP/yyUy1iVrZzs8rvSG9abuitv
rz1ZGP4IdPp7PhsoxN9pYO+VGyvXlU7NsSWS7TBFtW3sh1Ub8c9s4dr1pGFR
dxElrGjnaK7csZtJzSNM5/Ef6DgwtsjyUeTe8P1iDeVSh38iCQwLXKtxb1ve
tOXGXiVGNUuZLTRFyKkR9Oj0McKt5Y6inkBf6cF+kbQtzHm3jqePwwUQfjNT
v3zfsgaLz+ACwnNI2qU7BuyQn8mKjmXmfLc2uHsaS2DmhaaL0KTOjg4Dz1nb
tbHqsN6jJTsnOvUSpi7HNIddeoTkjX+mFr8S01iU2TfYGIWNdW5W0QEYfi8N
npjYvymoBdCUtyhgOfRIfDuruejUiDMEscu2GSHrhyf4ek6cpU743v4B4wdk
dLI4rETbrOljsoo/klp/jL+f5oXz6IjUo2yVmrtnQrDfjX49ZX8psgqXEwEd
Xvc4Jo+0dVki5NmnsiC3SpqiCLsm937/dCjxCHcOl49mOOmW1jIIWbDVXuhE
tm8n1lz8N+V7slG4MZeOhZSEY6faoVOZrbgUwWPw9pA8nSm4R5J3cYqdGltG
ya0BL6E/xMmpaRydaAZSauSpdlSCvnmKWuMbJAI+Thr4DLlLf1ZVCDIoxjM3
QgQsp+l43c8XPNcva6kp8lHb1OfdIa3Qq+/FpkpiJ8nat4OhWiDYffpCbY6Z
qmophUmDJzp/OgDjAbj2ngr8Iu9jfbym3AqHtIILrUrCmIEGtR3d083GFMya
1z87F3gtoTdretGN3zcMG3aQL3TFGn1om7ZXIHd9D9WRjeC/SuQF9pHd9LHL
+lo97xMB+Yaxoc21hV77VtBziqkAKCyRpkNKiDMQb7xCYuZ2CvFn/ujphauJ
VYT+sA74IfRtDQ9th1pocQYAwFdFldeB31IGKPjskb7zg06OUM5+4p8Lcvgu
20mQZ1iVy7bu5BNPOIbmO+6AgsMVEJxgLdtXiHsO1BRIZP/jOna4FvIpkjGm
m3vEWeGNepqtNEuN8Lm0je6lyigpxk06eIlNKWo0/5bs2UyZajx4uWe8O3Ju
bRofslN5YRfwA7I1AQxtnzriPgW2wo3F311t7/RENfpiujVCQNpSio844Oe+
cBHSIraqFSOpndnkJSo6OsEsseIUM67X4bWIxXutjGTEfplI0WREH9Fzf46C
mxqxEI4nt0oylvcdyTGFs79EtsmF1bezpThiJtzB+PMtTTPqBtxodFSxc9m3
CT9U7cksSaWRAaGLk6+SAu4tgAWf+KsuTCzI5i5+2i2OK8ODDuDuDqKMEMtg
k42YEy+DO31Hjfcgyx2Zb8J6odiFDrkTU2Y9/YMA9eOpd4R4x4/zis19vFEq
SuxhjoVAZiueNYZlNt9ihkcEuHPXJnAtQeuzsi3eliYRnhG9iGMruSUDkbh5
hBXMWh4K5mvICLZqlrfp00nV19NzGnlZ3+uROdNG+lAePWt8+z+8gjSoGNNW
IYmgRpaDYQ0Q0XSQCgH0jGz9uAmez8CkyTGlqQiorOLBEndAN09qnkSdLj7f
uUg0/d+GfEt82B3zh6dVIPOkoqmyDIuOt0JAc4lHEeTF2q5+JkjqzGJBsu0s
k9AOLKsVuHJzHafW+/Y1ik46B1mWWOvDqgMSMoMIXYPO9LaEO0EwvEUh8LtV
PK/8K2w7RyjH3ol6I8LkmMyuSQarsodBPLGLRQJGnuWEV4lzf5gRcDW9I2Su
0cQin1LorTlTBuz09SlD+8AJOpqpjxDG47fU2KNOTJ16YsBIv9rP9wIaXmOU
vXX2Irf9LUNnwUuuttDxYO+VGa7/UPozpFJnUyl9G8yApig6hwiCuS6V/jmB
z2nghVaDkGgiPdxFGChmlKLb7IWis/S6Dvkqgb7BpSBXxWLODUsrxSe7elTg
9nbpx2o3yJ4n2kq58kyZ06KFKIwBos4aZ4uT0BPWcGI0knTG+mXOH613UPqL
Bzo3ep7NDpJOMDduvJhHKMF5QeLYYf4q1aKR8zMv0NVQcLI4J3vnXdZwP/zZ
ZV/1W7hXRnm+/L9jPx6RIGzOxrXZJoAvm48Cy8t9YdB+3CMP9yjjiahxiZTb
HqKLhhHRByRPJfnEsar/I4uL0L2wm/vqLaWMD8FbvFE0mYkFtPLgnicSALZ4
fgIKMpSu5/Jg/t1kc7NWVl4q3+0eql2oOoT9ZH8Ffqqj92dln5UOWg/H6GWq
CdquNFnAY4MJC/P7qS/G5S8IHpgTCfkY8RN1EveMaAA++bN0+VrarvmJa12R
66ker8asbVYg9VJXS4kwBFKBf8qgYor0s72yHKIazOfBLfBwcybnsq2eOgrE
00hjsOrg+TbZNi7oLdMB51QzgM2LHVHmj36VwxGdqwaKGw0BzU4HhpMHGpGK
XTlus1tD2a/qO0jcPXvUylhemWBccVpHh9EWuBxS79c21x43B/MCB4saTLC9
4eZSXpkur/XVlEBHiwnDt0sgsOXKS45kx0qfcKUovlAGHiHP7UIZVGrL0JRu
yrTurlJYyMTbfRfKIEEgbfUYyQwAxsiFYKDeO30fqaeatKXmtjiCjOaa8d30
a4/nD3rAiY9FyEXCKYcq43ELEs3dRCfgj1dmFOCviwc9irjm1O0TayJF93HZ
yLNYpobmCxanbelEQcH7qehsq6/hBtfwTD6GCSHnZOv0dAKomQycA/NhFpnf
z50VfOBMnxX+16WOSu3YYsIW9helG25EO9RB+R3YoEEQFv9c+cy2g1yKWL5t
Da+RwYx1wKKsuK6huvaeryXHPI+OzEKJjo4qkpqkl0R+n2TNCh86AU3Qy4Ei
5uDYe857k7PAtAV+A/X66sFxF3CrJVHKCjcMC3KGfe9SPjozNvW6eSgEHZXT
fdaJTGwx/CD3yQG//wOz4fq2a2RLjsMI2Osu50+mcNU+ruF8PGu/ZolFfN69
UC5TjWXc17bIJjD1AefFqqsl/9ia7K0X0+yX9sxc+u3H4lm04H40GbXF9LvA
CHrkJbr6NvLyzG4o7sOQMTqBm+PzlA3Uw6L3m9/rR7XEmoKmqKY1DGieGXmd
quEbqAzMpHkf2is8IeQvjA12DWUGFtmRUq4PVuFicyCoZ9SD6D51Tsylnp1u
sMKvZz2vA2BDr/wlav0XmQeb2Lan4+InHEGzYZ/o5Z+1Iy9ntJs1BXT9yIk6
mbVvrmyestE0ztX61cRY/YRFDYxwReaxRun5K78XmOys06FWg0Qmk/cLw1OO
G8TBT6TRnVxh/mRQXi59v6fIOrZ6s3aXvil+oHhY/ingIAgtZD65so9p/UYJ
H88IsPR0DjySA4Nw87YYE2DqSdis8qC/D9LjIuONuYVIeOdMsSkf+bEWcD+0
1yYRaeRGqRaDmUgQ8cNrFjTo7LKEeo7SUo63+M0hvrNC8FugzzvY2WBrzwv/
3ltZy/Orng8yTOKikymgnasLKyO+8ZM3wWGCTmTUbAnlhf3Wl4d/TQ6TfOJe
uIG+EBY0D0G2AR2SzR83Bd8L+RMPgoGAhQxNXH56WN4R8qY3NedZTXNj36vA
Cw/e+pUTKU1dpktWpsuMiE6JfP1khqFETxTj/1IVBJFSczLDxZWDW+yeUgnY
YuipwOaoswmkdquTOPdDLyeqwkQdm8/11PurRTuxeatDxsCKMglcABTazf2d
L0tCoV7j1/VyJIU489oRNIXB/vW7kavsEAzVpkdRL46gQ9xzP2cHLVW3e/9M
sdvy3L/PFNlpVaPu/yiQgrybTUQTkBkRiAUFX/KR+u2X5LsXxADUbS4PFfq2
O03IUQb9/93ZoOJNudw8qje0wbZ742wo3HG+vAHt67tLVta0wh4GFb3+uHoP
fRex3vCp1bOmly4x9h6yv6iNxClCsCP8F65OOzFGOdvuF30BjSjCWRJM5pbd
QXzebDAQYKMjUX/h2VRAMPsfuk0W+Cff1OfiLVpwDzhVRbnuPXDagOEc6vYw
XlQNnIUePRUMIBGjyxG1Tv67k3TywbxQRmj7Ucmqzueo0Ug0xCj14CQ7Q20H
O/zaGZAhOKlUaCW071uvlomYSndqdFSQTMqbzZB0Shh2Ezodtx9nzVdUjF7C
yWDi62/6OtrfJAjnWU8VzLniVDWJmJmZISU1vfZ8YwpLTDZ8HE8GUlUFhi9W
iOVz6g4GGm95MxP6ps1xAwmz3hvbx6/QjLn2xGsj7ukE+zttTv0KKweZ/0Pp
eOixJILUSpsdgrdEY7wtZN6P0rMvk6Pu7h57SfhBsR1uhI0898Rco+IvVG+I
DF9vBS9fNesb43fhnIXfg0ubOTz2m8mPEetiwtKVwpzwZrhmbjXMt0Cq0veb
KXSmd+zC6NauTHInsYbE0VSKU7zmWrc9QK6/73NewKgY0FNCQykJez+CEim3
tiBUKJLZSuzUV4pMoLnANEQbeavqIhCIVMWL3GMOniCK5zq9ws95HWCS+ovB
0vXPXko5Tbqy9CwsdpIrRCvJZHEmrg7ZkwbbhC9ekW/itV2puzUmyFKzz++Y
O5z16e1Wukk3fRR5M8+aKhQ+Zm5xxvP/sGGUPHsB4dE5W1bULCOiV/64xmVs
WOIEU8K/FUxk9wLDqQbZSm/OnxgzKP4hKIcFRuQ7qCrhOo2TypcjUdamhZIX
N983PxVWv44SrxPmd/ubZnKO6xq88L1uKf9cC/Iv7xJ3nS5fuQgrvT7ciu9Z
HjAcjAvTS0ULvVnib9ffhqOlWineqTHhnpMjFrKgCDiC/rys8ZF31bu9E4KO
SkJ/hMMzV6cp4Q+2/cbfxnn6sxcU6FWXlW92Hxv4SYi0P7DBqR8kZnZWi88y
ocdJXaiQRi9SjHRy5noyRurtGfWdgG/oCb4HQU07OT3peIjYe3S6e9I5fvGL
YjhALw/hpPP7m2QpOdzSuzxPseuz+Tk4ZBVhP4ZAol9qEoTQZ/qxvXTeDlII
SYtrpLnBoAg3FLC9jd9bexe+XJyDVJaGzOQluIdyvPMSW/6VMjVKLSid7VFp
UZe5m9dIBpAbSV7SjY3ZVHB69WGkT+9a1+16Z/otJCPkXT8Bm+iqgNZ/rl7x
IkYTpIjB/6KHRIE4wQFGvnPu/Aayj+QiiIdfHk1zZh5wR5wlt9c0rR5WJU6H
V4X2BCc46nUUi4YfZavswlytd+3EbDLysUcMPppIsmN8boaal3ItGXJph5TS
8x9zm6yLFZRp8DvNpW0HVcDGL6kMJqpY92YKXLSH2JuiTjT4jaUC9nzuTVTe
x/ooR5M9W90dD+NLbOpQMQEdxSWBjAEp6270jO3Za5YM6VFCcPLKsvje1+Vp
Rr3Pg+z7H3RjgGu9GjUc2Aq4VUgYDlQvE4TNd2qlpULqk24Fr01dMkticF8J
hfPpPAJAbZQr3bKlW11XuaUx1dRajK80vGebjzAWd2Coh0hW/ROdYa7DNhfd
zpA7JFotW5PoXRTtkJ30DJlFOkb7nC4QY5AosfhCQtQ2ohPmj+qXvzHPSM3o
hY67pM7gqZvyFDtaE94Hw4edYjJ+KvHG1Y93Gw/qtG3ulq1c8TptWaDqach2
lEvoU5GVYZu6axur0c1gI8cS1loRzJcS6UmKE5g/W5N1HoPFBMQ3QM+v4bPk
p+4xVTqGm+NvwwGja/F38mM20NXeWjXUTAVPf5cMBpXdAL0ZNLfZaPYEQsoM
TY//MymOSaIVW1ngRSn2LL2qUlba0qYvu/S+Ia9cMlbAaCQqXcBlF2XMUt+g
KaG7IlO48XlZBI7rX8xIpOfg5t4OPL7T2ROZtnumnlah9TjHhxuZKDQcNP6x
0KyNlzUxJz4Lwz0ix4HydcPDHo/HHXUZHCHPYdMXNiv+V6HhlnuGZW7CJ4Zs
BVbEVe2+vTELsPpUHn7UlStYXGLPZ1/vB6ZBJFdLyN6fpEU57b4oJ3PlnkP8
kPgX99fyDrbyAx2cKsTgxyu2gC49yHUS82akGBvZ/eJx8par4qetk1Pl4fvo
CP6rAMJPqkyWWHqJL+DVixZ34SZXbRudS2ryb4XPlVIgE9IjBI7c3U9TLd14
HQbXtiM+KH0jdA65Hg+k/2i2flCYQN9/JjWEuTInF43IQ19cJP3IqaWftfnC
E+aR+EI1jJlonEh0cUeilVqtB2K0WAt9un3K3bhm+l3orfK/xrbbOtTRKsnX
nI5bnFfE/CGAv7BovQmNMxDVtxVXsjirxAyfc2Uh2vyQiWTAOrKzva+E9P84
ump0b4MfLm2oV6E3hArxtjEVGuObVLJL3sQSCs1L04wo4iJSrclYjXFVOK4g
gdfWy9zEtJmsXuTaEYxDDl50u/0fLYJCClpPLoZY79NZRf+NxBmkycQ+YO2M
bYpGSXTyx3dBgrSDNE0SQZD8h6Y+aSOjIWBeXNYbBFo1R/2uAMcBdfuoPGS5
y/3mfPhZ28vVv/K40QZ8nExaCWRIPAHM0uuirHrVrITzLqYtfBJxpBhPM6d+
m4eNn56gKL/J8qcR+eQWFBdT4SSLFQYr8FDgXx86GWTXUqei24NahlA6r1b6
AQfnbr+0ZY40lQKl4mks8x0faXPDYk7+wz+uZXhXSO+sCfKJR61chjG2dFYU
SRqeJ5O7ysvbcn+kQVM+J7jEyQ+XYf9Qlq/XG95LTkPvTlDz6Psn3jthRhYQ
c8/MwkXqhMPIwQIeBqedykS8JHLg4vwVzfIO3XWZhTULzpW1j/HBQA9FPdzk
82/w/CCzlEpIKtHR1r5cPDpSntw9EiFKsdN0l/3cwhbqZHrKArU7aWJZ+pcY
AUM2uugokFfrKJG/F7b4QmzNyd/3vP8EDo0mdc/TM+tAgSvWCqsVKfMDDCm4
ohiXozF3Ptl6LBE8bP1gaNjGrqfgGEjfOiB18dxUmu/L9XGjITL/+1ANLIMu
avJlE2PitdCC0OIfrQhVgTpAhCIt/AGwtGsHq1AykMj5HVYkQRJNiauv7jIb
tKLWEF/z5ppOz6nwYzlxY+3tDOnTeyxrvmHlJqF7xs/hDRDm+O9daH8R/Nr0
+suIXyEbIDzHPHuJRDVogOdanaWcxmAaIPTORiO4Q9L1XFfPrSltMtuBVaHJ
xqhKIPpnogRkE4Xyua3Zd6CR2RSgDB6A2nRYC4apaVIA4EecVFNMDmeIeBV7
H0+dxwKOiWh0lXLSDQ56eDRsb4ucDseQQyEIQU0E9oB1JnmoTMoBBcup4HVs
emvOgAZVjjvK7KZT2PW3d9Uo+qFn4rh8toNsIa9cvpEiamA1TTXqEOWkk4mT
Hu0Vubz89QgkmHfWO60S4DEcIMeLRkcFkaVRFILPYR+CS03buzIyMvBSTFb9
hPcEXauv4FBWlmT7ffy8juyD0NFjQ/573CGAH7SwPQUQOZ+1gKCIfqORoY9V
d6WirQ7tHiZdDqXP0wgNrvCMNAe0j22lf0Habfu4R+JXP94Ee40Bwf1TbA6Z
yA9/YOBURS7B3TuhbrhvFg0RdAgWyHcz4JMzkRGEef9aoPHdZtb6vF2Gx73N
Cpk4/uFgDHeSdRkxmJjZcwNm3qGF0PA7Ec9Fwv9IZKshKRGk2ESsPsje37rK
B8NvEnQkoLQoRVBrl+SLT/IopDFQZITgJ5kVwDgLZNhcYWnBmmKXw+5jIG7H
2U89kPTx0IZA79iZ1JTw7Kecr1YBq5OsXFw0ExyeX3YBTa3M5EeUqJs0xpVS
M5GEQ9e7i1yJ6KT3juavQs4TOOoII5coAt+OgU1XtaPCSD+LjMUHsF2dQP7w
tRqfwmK84rg5a6XPLOaLcFr538ZcJUdgqveYGSBgpdcpILgeHkp8BuG/BqhH
wkA9VdDmS07BLnso1WwJ+hHMZEglyhSdiC9CsYZcxc2Kgdc3GsTn7UwwbUGF
7sA5owCdJMbYx/kXCx6MPXPxOJj7ABOlAvbeQpv1fWR3XlkW5wS7yf2SOoU+
rgvqxqe6sNb4jPB8jYlmbqjPK22ragjPz+bs0azzNehwU2w4b+7Lq5rTU3CC
M/F4wGNVP9HKGu5EgeC8FdoAMJXAHKIg0VvYzixhQHqTjbBnQ+DvQu6q+5KO
RZon2j8aWh+tglVOKWqmvGTXOoFGrYdsbNFfOzl7VncWmRq73962U3xIsdgJ
f0ngT5PRHzigFv9zTUxXowx8xChrpsiyTNra8qQk/OwYsiRE3AwJ4DFbb0MT
C99C1YPDOI3QlctZ7kX3vinF+qfHRzVMpPwEgjqpev89BljC8HKija4qvJpH
flyOGUThVmwfZR6SVmji2dpuaRcjKKfnd7w+N4XdBhzgyKlU6jRIPZJab8+O
lzD4lWPyLE7nd+fZ41/BoDN/gbDSxO6yWTKCvsTlvhL19H+z+9e+THR8eZcD
ZMilmfgxyPTFenh3SPm2gxHm78QjOezeQjrU1WytpltKspIiPPAy33G5GUE9
54oA1oiz9CYfMVhTIlWMBAa9tgqlBnDaGYOp5H0HqVAKrVyM9sG9y3l7ziwi
HDVPSAI0rAMTnFwa3hXjbgB2NQrWEW9cGeDds2gFirCPqnuFPAV+5VNY02xh
ItBWr41PKt7bzrgsjOqbxOBPkW1YopFXpHkovSjzoCQLmJWYz/gOI1zuRT/A
HOYcCiu5WzbqielbCETK0BU78tAsGwssLJBt+RwejiY+FoFJvJYFnzU1GgD1
raIcj1fslcj6wYkOLkqm+9ChCwDrWHRhzea+mUc7iXbk/eSTVkm/qFwytMi2
tIeSvZvEOQ5bmcp6ICuyQXfnnmQ09sMDKt+YZKrHXvstw0c3uJ3EnxBkf0jc
qR92+haRQ4h6ucTsdf7nOL3sDoyiem+8s9OJJL/EUDU/TiBgrwBl2ccGRQMF
3pbXIiz6vRcaYgOk/9TQe7Y0W4dRTE4TnhmbUA3obUMi15SObVxaEPzCG7vv
J+bB+LU9KK270u0sZxdTcMAGenuifRJZB4xojxOeHz9Fxx/odZf84vSTCimG
Js+abizqxwg4PKKR9PDhAYwrbGiLJBMqrusTjUe23J+Olk0GvhxyDcGAvrAc
FwCImScGMxJxn75MutO1O/jsBS1OsWNSYicjaoX3ourPNWz4f2pYp51efvrK
6H8kMaaa/XeNd8dy1mu26RHIUBj1sMfsH2HgtRd6K76oF0fnc6olfUvsRDUY
iIYY5E9CaUsHwfpLYXzeLcRacywv8DN2PYKAH8mmbRUK/uPx9fxUsPXnQDIu
IGyOq+PpmCaFTFi5Ihwdx5rgjAaOl/+oEGe39XFbqbNSxlRS5HxvkGqAdoZt
2+JnBUynLTUerJVsmSjDnC0d+ZyTeL3lQNfWNHIWvpc7iaaenQUr2XG+4f4I
prGRmTchYtKMK6z2nWkRsnDWLpgpA1bqK06mKJnqbIGSAorwcg9zJolxFjep
94bLXMMURDapTKOZUMFvhHoIj3zoJqQEGL0RKCC5nCH7fMBpS36ZXiE9bVuo
qp/VFBbtD6J1kuHnnc9lIKd5+nVAraQ0oqsYbaksDft1tEaG81tuVc+3soqI
p1M7SvzmyR1DuU55GenRTuO4pw5mhVA3XkZdWCW0DqS63Wx+q87e9X2bJyPy
1hiQwsQXPvzY8Eaiz7j1jUMQow6cVM0F6YAUa/6QmTtBYAB05YVqgFg6jA+1
i6aBrqKf8SP+7ze4pbo83I+QZaVfM57Mp6jocmFv3vmmEW/EvuvP075gzjIb
QpsI8Qx6z9HKuiwvJtrIpRJHQSHp7P6M51pqihj9hSHK1yJ/aAym6WhY8WkA
17TLm/+Wl15DStIqbPwZfVBwphp+8MJHDnpHfEuD3tV/ntZ/yPczzc7+dR+R
s+CrPc8dMIdgPvTAZH280FduiVzWFEUXkoeHIgmWfeH4uze+oKftIk5x80i/
T3lk0R69bfCPWEROw8u7PqCN3onED5gyIp/foWRzVMkrwe1AA1ecnQKOP/Zd
w1I4JJXjqsJSFoP0YqGF7L6sKB5C179NNeN/+woPcAIAXn2GeZWnZgGZj/eR
YwP/t4D5qrkHQVCjFY2H2yx8u2RPCyPMlfcM5U9AWLlclBy31NY27y/i9XiN
AA/YewedJq0vLZR9ubEhBGJsivwXc6lKXhbJVEZ03V7DN0i65TGPCyY5q83T
idGSCuAtXUtW3/b3/KP6skBcb3TIc/hXz8xYEBeZrzPNZBD6JUMvLFXz3qVB
D03B6awvsq8tMJHTGOvBtWo0lUN6jde9fK7H2sEPOVFn89qBog4JyVPrFGub
rkK7uZvwRRH2VWLFiQd3jgNnPrVaWYM895JVeW9SOBrwfOz6qNsfzVX7+FSu
0t+2FOQiP5wnwLB8x9uXFdCWisKaAsR68DYhY3PuA1SC3ZQJgWcTd9Olv7lR
NX/zkMsNO0Ot09EcOJMp9sEtTSjmoSC2H0WCwTd6hlRG45w3ibSntIJEKJlY
ckQFNNSlmffuOCZkKx69J6Xvo4U+Ot552HPKAKgH884grfcl/2sosWJAbKuf
YIcsZK1hy37gyGupqC/f/7yJEyBYjGJDryOkZDjA856W7g/qLI/N/oBiT1JA
lzJCmIJi4t61Pd2RH2k79OgIHNdij0EYLXUfFyPgU2SGzopbEcjAg1fpXu4p
/NpT0vfynRovLYecPV74wB1MgUNVppCfGbGPYu+6/AYxgmeiy8HVFHCFogNi
M3b/kztNQJCx3IUFyF2OxKsTveWzmeKaood2Xa3Tt7lo7mB1FEDc8J93RRqN
xXRMhogBlGAi34qKnH7Fboad0sMNV6a1lcFK2DKRl78xFJMsYrFb73nOJ4DO
7/pALAR6hChNPUcCcD207u3keByz5tUhn0mBrBav+p3pnPKkHTbRrGCNMY2r
a5iJfHUIcD1U8MMuqwpVKVp8oKYmxROYBaHhIEZUGFgZ0Gx3QPxGrAWweA6u
aMs0LIuE/IBXbA29JASEroCWwaaF2U7ecNAcsruTFRcgZswoY7iceGHFWT+w
TuURQ8HnDDmK5WuXnMOhru+hNJNr2lsrSN1xk6HpvbDIdAj6SyaSFqXSyj1r
M8GGHvtVKOMAIdt1po3JBL2Iwcx8Nq+7TWbkV0unzZ+4IQ1WXrTz7wf69YnA
/CBcqIR6PONgDHiwuNKdl9ZlS1NfKw/BQPr+72zs83gmV+CDsxwF9rtrmKyx
mDoiHM5SDZ8XzGTYLdRjdfPJ5MsujeuffktFLvPGWzP4SyA09V0nQJvSTw/k
hnWPcMiV1pneSR43xyZpyHRGCiyUqwGNs4MuuvbtfbcpKceN4WQA+V03aSGA
DX5L1Q3KY0IayPDVQ7ahTYUW4IP3dfayNcvVTxcDl+MdpoeyCYDK7J2CmjjG
7Lxp3At6zuGgu20WDdOKDWjZv3FQPSszmsOTHnBr0AI3H+aAqeGkCaCZp0Ci
NsFumSuUfjh6Z6SET2mtST4a1YRD4Trvo4ecqqBgmECy8B2tWsKlgI+NRqNE
5M+eRopDB+2NXmzlvbU/CPy4DyLUUhbGsFpRkchcsDuyy0+AQ4RnJbQpOepe
0Tpj2RJBbgmQxn/gybj6HCo+ljQk6/Q129ExRJyESENq+r5yFbOZHw5qyDVH
KCrp6ioQhkxEI2/ow+xFYxe528lwwM7kIr9FCv1bIiDGr45AWZoJ1cpgYK3R
NbpLhgIG6pL3YhvM92s/AshS3KeRj07ow987dS4OfYaCF/PNm0dnGOl4MNRG
bc4rr0qYW56hom4nvoXHpHv5KjOEzKgTgCW2nHYLXWD9zQh55fhxaTqJ4q1u
GTZtx01WGWtQMeDL5gJWV+iBBvjIcToqfHX0G6YJltATg0U+kqo1TRNCbBzA
I9BFieBQapRSBVJG3clRtBKppzPSoFApCk7Oe1o5iGD29a/avTbO3EDuCQ0I
LhxE6ajtaBM7ep5V8F7PAH7CATTDQS1L0BaMLBlXq5XQAbA84FevM2S/7h2J
EwFin2cnQ44hrtvhuSQF+9e7DQtRewiFiFgk5gJ3GwQC49BkuBRemfc8wAKA
WkMFMiPVAzF9d0ZrXTPErlFx5UvVKnso9pVQRuKgKflSywqZFOX+LgNvKHE1
bHMticvl2SMCm8aSadK78OM1kN8TbV1QC3b34RgVXRd9/CgGV7Vxw4Cs2EcP
aCav0wJUmUX6IeHzA0nbFz4Iqv9IUHgxdPQYxOUlIJCr0KYVFX21L0/3+WQt
bYV7f4F8Rd2AO1so3N8NKrVAUkHuQJZgdOv5bP7Mcfjciuzb/cqrERlbtW8W
3DSLpZr5FBDP7yN8zOXLGGlWxOpB6VL0qCdIG2mVXpvgrIER5gQMZNBCPUCW
xX0vBqwAKVec8u6bakA3paFG0a0wPBgEef+hpc7LZ6Yq++9oEHdmmbYJe5z0
iHJ9w4IJjivkuOciXGJiK73VQZpvSHvVoj+rBA/qUT2pJ3zE53oElNhxYzdT
6yNR0ViuqCBjuSXPuxT4HNX70fpCzlzwXMXk2rtn21U9ufbpRjn22upM2Z0R
SBqKwlkawPPNKJedsfzcGmi8HxoFDnCBXeH0RJI+x0oIpBdEnCX0nHgXlBhf
ZbQ5q/LjBzqp0rb4yZiSr/F7zsluPlXtu4X0sBJk6g1fmexl5wQEnuvDmi5P
Csyy90txF+D1nhSDBmEPeOn1NnAVEeC59RpsOmcWwPzf84H/C40mLGmHU1PW
KJr1Dbc3nNHKlQ4GFtUBSgCi04ILM9Vwej9vhYQxnzsvcrJoZBGlilfojVyT
qvSRonWFqSBXfPrWM/1vkVWoCTlXcP1aqlXujETohsaVVJtvpxbFP7QfLXmB
H44/EzqHqejBBhx9Nv9Fw3+loy9sGXY44eqW1VT/cjYP5OYcZ63hDwiQ0UgT
qaP9PFEF1MzElj/vAf14qmXVmlR1HW6bdgY8V6naC8kRaL4DBzpXvy4HzDoV
InKZDRl6+NvBwXWQW/sqptuD+3AYl2DtXi2swQQV0nXLN+XZw7cSXhxqpXx0
WK7POtK2yPPnQLifDcCP1degP+Zj2kSIfoMuXJWpmcoYAHu24cLSrgtDDoKk
pRnxw/Ie5NSGGdkTmlkthdmXRXTWNS8cvlbXRPPrKBz1V9y+Pd96FBqD99fE
pFi+62BbUS+RBSY4if/h3rma3BuMFz8zNXt/4VQ/A6XBZyC7ba+qmNc6FNk9
uoGSPpA8RZ1lEZl9jQ6Lza/Mjol1rsE9akk98VTaZmOK7stucDPbO5so6ijQ
LiIJxYow4AutaOv6gRDWsVf37eK86kHrL5VkbNLATgMiKqMrhnLnDr/SzkOu
maJL7i6v+EZz4khnOuKBzAvUF8iNNOVzfxN23tDnu3exG1zh1dUZ1wX6Tjop
6gOg/d1gvqbYAN1eQjcuzE03xARcT5hqnuiLprX3zZY/swvd74jOUjCiEgtA
qHEsyzyOIRq6puPJCO3YxDv75VyW2E+CgysJdQTWlo9rS3HYD7P46X6q9fRc
mN15DqAitjDdrugtKmcKyfrWxfh41Ps5FXF/ZIn0ciMldq+nmia7IbyCxGit
w6ZVPh9kd6dgcDYFZ6b/9pi6fc2/9qSVz+l3t/T/L/tCw2h2Si2cL9/W91QI
z9OciwBPqXK96RLqtnK4XzWKR+98LkPpQGf/IzjXfrmTAlk943C2EYSq8vsj
f+e1e98D4sIphln/34/N01+D2XNW63deAEho55DyqJ+aQ5fE/ydT1NmK9wwI
DtdrJF6aK8RvxB09aIurwoIbg1x6tCYPgi8f35rghPDuiMYi5lusmuTOTCOi
ac9voJra+YAiggSKF/GZOPYpdqUtvIpnvQM3wT2uSKD6wirnnTmfbsoNQlIC
fqVAZ/Boi232NIcW6nSkIKv1K7qIcK7hdKLVsNNd4hFpGCggzu3J6Eeamyze
SliWLNQSzIB1rStvjwswmNuuHWSM6QAIHiw29pSu7Tv42dFJTPtfISr8rdnp
QJrd7aNKrHxq2Mew3gCtr6SH1/tfewjUQ7s0nGSPlPy5PEpAXzVqjhoIoReX
uXkCJRw6GvS+3L0RI3OgiPQoL00KFRuRkMnM8fEU1nDPk/Mu+eryoAml/q9r
yD/jdJQrH97p/EE5wZ0pTFlCJGOMXdqD1XND0g76ssIAE56qBPayoM70P4lZ
3KWj3l0SiKjj1nhRQj+yIsOFqIx1Cwwu7UIlCdEB+ZRyA9VyH0LWqus1hbdF
I2O8CzBYeQDOOkdO54vG9E/Mu1sLX0IFukQ9YC0Woq4l5LojEeHy0L3jb/+t
tp0XC5+7SoJ3xxhnR7q+JIY15VGr5agbZxP0YLNFvkNVFQ2DAGFV1iefAuO8
2l3M83XdUJ3r9uRiDBe2q/bIUjiwwS5JcaB/T77wM33cp15vWBzwtWoK+Aet
zYfDaVCS0DDEfx1nZM0tNbyeo5any0Vl6Qu2ZPL9IrBAAa+UZ6gTFChlUjhe
E3d16PG8uVMsNiQrmmU16IFoLSTuB4ORSe8mlkZA1KomnOvuXl4Klp9cEj6M
Gi/k7p2/M1Ar/f3wm4+7/S7cJXCvdOzAzgl2sd3i3w68e7vbzoIaJ4SWCi3V
zk4GJDhJ2XAWfWDYhfOPPGviU1kzXtDdSClu56pf+C1QK8vE1BECyJLA5JZV
ikyvFLnOpMesJinOI/kYTyndmGJXOEq1jO6mY72/wgzARx8lXYqKWPDmd+M9
Nm5qOyDGW7eu2qm8x155c+6cL16wRhd4q68zGvMsw7DyFbm3D9Nck++kd4bU
G7m/rrXLTDAMEc3S93NRUyuNkHaC4y/9a4StWKV1VB1R9irHul4G0dJfQ6qv
J0FdOgLaEtwCgPJ9I+MVaPoycVBTXI0aX80w0USO9Q7P453LFFBz+7hJjgqm
q3cUBfiQS/7gd5QxqluC23VOZ/yYMCcDZL4rbx1MAVREALay0JWS1HQR0N30
S0KqAjUsIW1wj4Rkb1CAI+w9/iTiOg+3CWW/ptR3Bl9A9ZCq2F9V37ShMLFo
HBuY6Wh48TQXIYsefUjw74tFRSqOhYJcfA7pB3gqz63J0roWBAMLnWXLcott
svhWD/OXJYjPTgJy8qywib4SbrYzB37xXhZtKIZLJ09S4u9VEzOPVgFsPCbi
a3srnTeixuDerftlOP/KHZG1m6kgEqkFEjnZRZCb1yUyU6uRiNGuIN0xQT8M
UUbOdeD9eo+0MW66l+fH3OL3xds22Gd2X5Jp+UbqdpS0ExZe2UF5bS8Wj0lz
O92vtxEF22/jbivUIGLJE9li8zlSBWDVMh24RVQ45ER6b6CjYOJflr99u4PF
a7qHc6NEXgoeKKYKo5uKdzwvDFUjYgHKZkmCJYeKJvIyGjOaldo1ONAcFe8w
EbT5Jora8ScSKoifTNteL8NGD1AlCJPoeD9UC8PoW2R5Ox7dQ9Vc8RV10BIg
qqEh3N67lhoL31F3n7jyygKEZ0FwTEA6lFrXlxKdMlDCK1uVcWHEHV4Nb1Rv
8rFj0hKExXizIFxGBGjIuqK2D2b4fEf+1Y0O/Nvl+7QlDq0ufzM7Gzye8jmt
kl3gBsUlrVpIbyvu/GINHSU8pmnttSYGJoqzs5pWfBQpT6+ZZXUysXg/u+ub
wxWRjj60GHwcpr2xl7Jn89bqv9ucyfaC+mplwQ3+I3X8qcMRgGj3J6J6iBQG
I75McYurXZrNxKk5a5TupA6Y+fI4nQyFh0R5lR9ruGkCphLVumxtlGNopEGa
NwrNH3JnpqTckgm7/RlI8MJChdtRJhA5j+oaTKttq5zoV2SjLSClz7gzU6pM
lGxBcsCYxgPqxhYn4o6fnQ6ku5nLwRHNrjX9t2J5yiHuHMYNZ0CgA8RPdHij
icmPOBYjHZcbVBdVDUvrjGJYegDE4s3Gzzd/CUHhDbbJWPjMXKSGFBB9G0VE
N3w3JCrjEpPVRnNVZQwUS17e1MjOb7S+JgTHgDk/Ja9iibZ44ht6wl7UTdWx
4HLfpp3HBm94pho5UM57jVmicDglxh5xxyDfOZtHM/RwBWezcPFTP7950A8d
M196gN+tKo+JllL9QhXdxZzDnKCwM+Y33Tl4epOULSsNWwGo+IxIZKpxXFao
Dbkb97dv0YE6dTShGUvAKfOsTVCNceLBjAftvJLK4tnB8gV3zgNzsAlgamKi
DArEdMDp2JaEndyOVZViyCkfcEbDZVOQBgeaOV7jbwIl0sYMI0FRnO5imTvR
bTbfgkw+bZcfWJPSF0McuUdQy5S0WiM0t7rOna4+qnY7TptCCjJX4VeiO6C1
FlLpUUaFnn+1aLnccx/obAn/3blHiWYZgJsLJ++mUbFV2uScal5evjloMCJM
pjne2JqAlnL2UKvXUDQ+hSe3EWDwWG0z2ysohA4Nq+czI0Gs1KSGh4oHJo9a
R3X1yR5DcWT8Qq11BQsQCI/LDG+gN5Q6Rr3Il6TenE2zpAMdfF1cdNX4k1zR
ymZVV8qrz02aWqtuaeLJ/MoJ8YXaZbH3sCyF4s0u21X5WBfsaUFPoZZYNPgK
uhUSAcrp6yy7gQA1HZ0CKRJBOA4BmFZrQ/TdW1l5nTdVjTvskcRrBXmZgwNn
sia7SwGPA6j7fW6koQJy7v0V0MqvqsSDTi5vUsBt4Wb4UNk37AFLNDkSqW4H
qUNryDOH0ozjJteKxg/VjrXyBTymWgbA7bKG1R7Udo2tTdkERbnjdIodlaAA
DQrKI1FUXDDHst+lwJbqyISng8TOKcETV6rtnvutGUXgxoJOTrq6aHzUf2Em
ZvHIxvaMpl9q4I2U9e9ugzb/JRVVvXeY4H3xCi3Jb8thK6gxF/zBvBTWEzk0
kcR19JUxJXz72hdETuBcF+nSEI+wEl5IygHNHekVhxL29lFwBXrS7osXE55+
Ft2zKar0RsjUi/+kGQw2WfPp/Nthna5aFuOclF3GAyahSZ00RVWJTUANd9Bh
w3ZPDPQ5K5Ml4XV4vL/5hkID4mVZ5M21C1o1G0+Gv7N//hwk9CGBkhlRfUsy
9IO1HSOc2XzBV27Eo0gyl8kTFPB9rq48fzZOWzMsGvf/4gUecsoDXTv5JMZD
/IAaA0lAjBl1l3OGy3kJuUmMemEr/5S3LkJ+IyQ2ctAeBA4Se3TUIhBo/IOL
+15dEhvoMn0Rjsgb2ZD6mrq+lAjLn4wKDti1vQsAampUA2QCnnWNEmvtVag0
rcYqhDQ3taUV7xNPVubCjq6PCjTATJJdYoC3DJM4vyT+0PcWSldHZRPbsLW6
msLJ18KWLxVKzmcvlDolnl626XORyTsQcHe62rBA2Tf+U6JvvhyjF6W/t4s1
qu76IEeMOi+aK910tjKAemt7d/mjsKgHDQXqW7gG6ky3gobk26OBBzMeL6IJ
/bpLY6f5iIvs3iQLRd3/8FEmpf6NjjdIFkweDjkhmYhT7obFefUWtIS2T9r3
1i5dc/T9dVZ2GaLhm8VcKuPt2tpdsQe+ZCwyTC01uuXhP8dRtQPWMXs/DQxL
e/Y/ZPi0qpCIBACwci3IZ9GTnp9PsIMAIDIaRRFAiCH4d9FF8tPABE91D6Fr
tYUCgoow1xrAxoy1wguFvDra7iwIY9k1ZzvWZ/0AsZAocQnXMcMFuK+yXMhA
5vVSEgFGkvl6zG15SKgzDZEBmlf2GrwQQTG6kYBhIeX0GXl4hoTMsZRWBm+X
ahWtCi+odGrM7Xr7Q55ULz7UMVghEaUcuXtGWc4fr1lJZ3hPg5D/O9iiepJF
FFzGIUHyLdU39YIC+cZZkHO5FTu2GaCxLSg2f9X8TGzJylitVbquFpiqf41y
NeCd8rQ5HO9OrmkpqR9xxZPrId88YUpP8zINO705h4HTyOGmMjqrCWPAr8de
TeSu5KktkpSKHQj2jQShl4Xs2bkGRFn5vKytu38qQEIoJJYu1WEewRZ9klXt
7BQh/Sng2eNfeWGArm2/KkS4DFXtYLqsReUrNv3is6UA2aC9Oqi5DuicVbaK
Hq/Z61qF+lOCQqyHPj145/GY34IWzhDzPLxsQh4FTezwyRMn0Uc0IQW7T8+n
Vpinq5kzVLw6mkNCxtG9iFD0ho4fjCsgx2h445AWdY8zmh9iv20Ln88JS/Fa
AvM1x2cqzGVTjT/WNXwFAp30Qz83B5rPFOCC+VPNTl4LX/flH/gqcl1+AasR
b3NYZYA7xqtw1fOakIPH2/tmO8jsy6i0tinof77vNHKReSO3+uDiozjVmhRH
Jj9PAMFJeq42fnWsUcBNfcF20AyFDqzYV5zYME3cPL2y/pSdwtRgbfSULL7F
sfOGgdnD8lR+lcKfOKY1O/mnJAnfAnHh3lGDsiFp9x9ahjZvilwXk38GBetg
TMoq8f8x/YBYOueegcmPE9YDuiMa1QsCbrnCrKA0MyxkLHvhKVKnLpHzkc26
5K+EqVGinXRPf8DORYbvPDVVZ0q5Y5Qf45LL4SZQClk+Mir1czSu+qeAKAuh
3JxiunzBE+BEKR3SnucHuiB9hg8m1+K/oomoctJAcVk+QwawRnVF9ExZba/A
r65PCs+n1yBEvx8gMmL3JPWLLWZEmvVpsAKvio4FQjk9QmPRAJV13f1ioeJx
CKEZTFuP6c4jnZ73RwnuF9PKjDTTFbRJoFt8y+uJbX5DWFkq8KE0c8U+seII
vyon8h6YCNgH4bTwV8slXFoJ8ER6XHr4SgVO8j62nZpmHQWMfz8A0Bj67Dnr
OUPBcp+dfr3dPRmxRHi39ZKujHqTKmx6Js4fbjJ1TdGckHzt5xQneyT+bRbH
ItAMP61PWDE7Eo94LWlPsrbntlXY0KiiIL/CoYyry5+V73u8chB8SpyoIZYV
xedKQE/ma0LvQn05u7ZEerJb9k1Yr3q5sg8sVH5gS93FPHM1xtL11lBtWDZW
LaVcMtTYmzs4sddMfz5V9MScVWq5qu/S0xYZ3zLlT1GyzMOKC9X3GJi0I2vR
Fmsqd2cvjTAbm7UKtsmYT3+er4UTfL+2DEfPrM9k/Wx1RSHC4fkeffcFsbZo
8d6W5w1JG5kqMqU3tqayAP5nDvk4rzul1uXcEVPkm3WT9dyHTMKI3i3f4KMh
9ZYyR874Xgly41+wiolT7vxtNfJzpm1tdsuURSb7GiBIb6BjrMgPePgH8d/z
V9bulWo7AXqtrvFU+8UVP57ccaqS/zK6/ytsNGtt540GeAgBCVsmSetGQCku
mtkWB/jC9mwVmRulu7fMIFAFaC5CIEC3ATJ1ECoTYC/FGciZnSOgkCtQEBdn
vW1xnT+y1Y1I/so0UVIPw3epWn8dtWNjilDw870kxQaN5uLJKA+eQyQqDNQB
nojzROXPW8+Z5Ujgw91kH3qYc2HyFTvlqtnFzUB5kOasyvxsXaQL5qJ00yi0
j1/JxuKnCDXKX89wZWdm6sQt4HjMql6tDdU8+1n9BbGpaonghJ6/U2+1yeWh
zRX5TpZsW1L6+q41f7ICUXzXTahtYoN8Gz3lSNQUGaYo9zbMP06yu7C/nu8B
v+tJBhVpnwXCznRFo2VU6AhtxSyeUBBj9LkQdVdP0cwqEVx50mfqDIxBZ0QV
xJZmvnXyeeG+nK0HEe1914w1HN+ZvUWSIu7IJXNSXocjqIvqGBpj34i9GVNY
uy1qy2ifHwk62l2swrliLBGvV2TTdnEbblQK1J4MG+FfRiSySwqx8yL2sSo3
RaFwX4tU9X5k8TiPIuY6lz4Ih9T+QDgso3738YBDMZuMKXglPrTT27VSJSWL
9Uuy3qbAdevmac1TBQRFtCB1O5sZN0na4FDipf1cV5MJ8ISR4SGUBDr2f1tb
OdTt7u7REMVM5F0Y2zTX3a51zeikrjjEGTo4wMMzhy9CJeaZURyCB33qTtBg
dFZanN7Tqct6cyQg8S5eJcM6guo4C4ertPgplpacA0avWjViXEFIKqGmAwU7
BQryP8IhXJSGPATgJJGjfzOGa67Q6K0sIRitix5dDsWe5k9S8rz/UuHMLCdo
quhSUOUxS7gA25WTrJllDY0L9EkSZPC6wxRDHKMo17r1zPIrsksFAhpG85yM
lKJGiEMnIQpPlLzz15FuTwSI8Yx3nJgdMFF6g8CAFLQksJTEdWr5RxytDz3o
qYXG302U9qPHnP8vxn+hxSHhQghnW5xBudLJaGw80/AD9SYqLb77Cskvkumj
8BHfdBGwysCg7OuC1+I0InaSW5JsSXfDDUL9YDwkW7KdnxkYvLhDe0zrVahA
lQqMNOoQuoZ1g76fzJZ43/Lb0NEiV9wBgM9o0swl3xyuXP5XFyp+VvdSEiRC
XgbepNbXRl+Pj0CUrnegk8nsW2MCc3T800OYlpOwG6/GoT04GpLVx0SzPpON
DXr20GZqALT900ywzvRI+2+yLooiazBqxYefpQ+eLhcSq/Vke/F8DCnGgsBN
QO+eKrvlGlwjrvzsGqddprrZdYpdnx1//8oW+pKqmUQxwQ+W3z0uhNCjGEZy
rYm4awozQKGW8Px6W7clpLQw296I6jMLkq58q0leFBSi95b409PhE1PXI6hw
rsZSpp4/AsxVoMeJWEa+X10ZEbdFFBTtrmfvBrOjFeu0UJpqcfv6bWxZjLGd
2M+stv3xLUSVVIgxWhQML2vbCShjU7cB39A6lId+7ICR97yofFvt/9lP+Sg7
WZo4Z/7dPwk2t4MFXtmsr7iiCrziKc2TJuRVtkF8YfzLTvfwKivC7l/KhmSF
c+r7PqYIlerriWI5eaKa5spowgXLEx6DtZOlUYorT+yTrJedMqOnvcaegz08
+SVLKqheMwyCG20XjyttC5CocZOL8A7LHH7njvxWmZfUvwgGx5xgDeEBCxNS
kzknLqZipP+73vAJ1bNO8VtiG/RctZQe7Bcl6bwFQ5B5NY7Fz0dsgmylKHY5
xvMc2iYfeLXwlbi5YK9FqJAUgMwjlikJhpMOlmAm6Mz7YMMrDb1CxHzkXJKf
nqRdGQK34mVPiFagShz0noOZkaLgjCHaWl3xN5dy6XDNLzGC3nuiwlS8vOlh
JiGAvZZjILvcmtlE+nNcXOsU2wDw/Eix1A2ueIklRa8WJ/Tw3h4X/jdNG3k2
FTa9XSfGsvdlCZ3Gp8WjK9Jz5jbWXLJZfa6HRw6nQOzlvHQiQSZwxY1LF8xG
AWITfOeMzqV/+vJrdtaHSbtSwDGetBNj2PgaZV89qekrPhT2tNOFe1o4IjEE
o2YBW2A0VFcvX4tKBOiwUTeIzCqnbBeIQo5YI8w5btcEIq3y166eYrEZjBVl
E/OXJC/p+eqBVg9IVtr7ut1V2kntZYYQpODysibce3Np/rmA2lXy1/tbnw0B
/KQKitrxr0pDYUKe36zpWhrjezlWtvcGs8pIWjNrh1DqjP/W6ho4rXwfFZMz
Q5qCMQjEI/mPCEuEEHEWl10oHA3MGB8iPbIA6PqNHcAiCsRASoWW4ASQXmOK
BPLYh/DLdOEqasxRSgOidg2UX0G+8pLtmJ9PGb1hlM6TWEIHFC/UOA8rwCVH
WHl2hMw42P9C1QnzFZ4xp2mSRnJVnPJtAaP4032VdZisrt2JZpQdQ1NRDob9
UIRp9QZmH4VUcRQTUFPogflhkvnkkANxEurc8nusg6081RD3mQIQ/KUVRaAY
j3DBS8yaMuRxQSrA8rvjL9H5Ci6IjhzWbI0a2JARJBPItTCs4nR/cf0RfZkB
v8u0CgFeHXXCHGT9/5XK+3fZ3xrz/lTvIvXOuhGtT2X9c+aWsqeG+aM/6n7C
pd9oA2/sxsJVgbOL4BtEV0FHV/qIvrb+ZQSDfK7V1GcA/YTDcQrzRZoRUkxf
ELNZO/Ewg5NV2FrultgYBEEmMnuPzBsJhs2hhZOMVZQk6Ty82g/9vJd0WM4t
Bw5oKhu1rrw2fzGiroRX1IZlkmIL4JewwRTbHUECCPE8vUavn2kGpkS3h3iV
V6eDn08YbODyXzfpvpYTq/zmZLdyomgx+fXjLQq9gjaz6GuB8r5BOJJ8fBS8
2tLZo5SU5zyWaXWglppcTigGda5puhMccgN3xSpB1sQ1Qs6f45TqedbM6lNp
MFaFhJvwcsUW4x3GadeD3dgQ93ULqfoE0bdBlSylVaDoTPL/nQXyjjMSXHSv
HaGgLEoO4C2DxKtjc7fKmQOfmXPB8DrN4bpGwuuXxqRgdtATMAK06B3MfE0F
ztXIFoLgqnpBELoGL/6bofGQTqqoiKFpptBHpcxQTxahHp1WcA/pzDwC1OHn
S+2EU9h/YxXLN2452bVoipvwB/XnNHGGu9Y+6ZCJMHar9lPx6CIsuA3QtV0/
LTIOE+I/Q846ICGoJmsyxUNZWB7l54Pr6pafCqrzlLT1KNA6EE7ji4yUu1+i
e26wask45Svse6FSoL2lAuSPZ+3tBQoawZgeU2ezzEtetlGSPMEFdvGL6TJ1
GMdZf1YxBeBHJztTu8dIZCi62gab4u6bhzFJ5Q1Ot3rBjwLqvC9P7eb1AQJN
+rpwM/A8kEw5DiYOciqqhr9fdYSngnJiph/8F6sRxm2BABXVydQYwbeDg4rA
QcxDqFk1oYRrOukhAz98yeR+IRsosEJ7MwxqWwCnW0MnUeYiu5mTQyQDjhzv
ifo8EfDuB/QvvxgMAxhASgYbycl1yHYeiE2HhcmnLsVflhW6OQODdxYCo+R7
SzpHE24Q1yhUoHQ3IAYSNM5iL9+n0BrPlStXZkPzeAubKhMSlqC0F5EkGXV4
I2Yd84+c2d9Hfj1EeBwzEyRYxVyRAEQZxzDu6NgQtiqI4B9iEWLZWs6OHTjf
Wc1FSfMAkVn+nTjDT0FhFMm4zOBNuvDldsCRnDAw9I/kJ9j1DAxqQzu5oBE2
aQC7V+QhktZvfrnmjKwJiKOQMCXrDHBfFjG3e/awGXsd3duwmMQghcgWHkzF
LuPVIZiao9+37+qAaNIeiR820cTGRJnZe4KvXpbb+vWIHHhiNUxritGh2hUO
TkVy30s4zqbFv2HxFzvG9lMG5+Lrl0Mel6kBE0gKO941MaM3cbu/zb8IgmYf
yeSe5pIWeDhLUISjQByVkgMEE2FyyF3PvrYrNelPT8eyXx+WaGIP09dyiij1
DlnHJADvi31vplSuCSH36/AoEiJ998E2F9CTIlIaSSwNA7lqf4flWGnyy6v4
Pchesrb07WeQ5s7p0QhNtwgcgg7sugg7v/uUCCkMiSMO0NzEiHrpmBQUMBa2
HlLPFrgCUrYhbklIUyo99wUAdua4lpYJ+h0+SOh3d2w6FlErqjY9uBnNMYqb
NzJF08kiWZFIFjIhcK0aSgK9CvnCUZ1Tqu4j9ALTpsy3aG228nnfUJVFm2bd
fjMeXkyl1k4w2X6GbmTTmdAL1IMZHlrAnBA5o0C52frAILrYkJcuX5lEKp+E
dUsT+FYU6mko13s4s7k+U+a8i7nLyHWxbkxNAPjuP34q1pjlOKLIHKcc3xaj
V2isKfoSqtHJILwLwtT7bdt/wdvts2sWiKfG7hCQrtywGQ8TxIxy2qkmuH5M
b4BzBc8EdG+StUe1FpwZVES0MUjJY17qwpoeWJXReZnLxwuzEo1H61AmYtGX
f+nijgyPlDh25kzczM2xGwl4zMsc+5XyBZmQNcTfvKvMASIYY89CY3af2JsR
yNrtXrlwGe/EDTUJUxU/Yf7YIvO0N3cqpwxZLIhKfiMHjbEWh3CRMfdLDiMb
K70i7Y1y2w7vYUup+UCR5YrvbhTZ/W/lSJpWiUf0PvFqLBaeC27qU9CBifTz
sMWRKoURQ/Az/ERtjVTX4+9i9/iqWizQ5C90GzmB8cwiptOTjriaZg0LhNxB
RB8HyuqqcL+ccOrhqTurMUt+QrBMvgjmmYw9hvCKT/j6Q5rCBZuSrAyXAYK7
/6JXGz1ykcTMo01BmBvkEsm3yzRFGFCRTj+wtA0PuEw+9AjWAjnwBGbeGDhw
eGT0SwfyRxqs8LFOCKc1OeKF3sCvfm/ORihKkZ+omSqP7SQgYKgWx4fFr71Z
gEo8o7+SbRBkJD0Oda35Sds7m5J++6GPmlm6bLNdc1gH6/nLI2CunZroSVBa
OhWmVQKsAMSwTX4KoiEIQtadjf5XNJUNC1ceevcdZ4qDrwrVC7w9HS+AkZ06
ZAHeBKeiBjl6MACsfek0PlJliqNmxTd9HngozU13aJa66bUgn7ndH9nrW061
VoqjV0tM2camfrSYpMPreulbmbLcaOFxu3Ucu5qfKFJd9aUb/s4uMBNRxVQ3
d3m2ew+Tfae794HaOxPPDfpOx9ooWEZolYScTyX/CfNgQwhITWbIi5mP3U2T
oeq9E6dfvplU54hs+crL5w8WYCc/zwtwXVe/xZlvmxqeu3Ox/20IwvSGrGUB
jE6+WrOesU9LF6CqUJOLVBEC1Mxxdl2R4r9Ao8LU+2GEl8lsGbUwpwPAIO9j
bF6kgliHQO4LNrAWMvemS8It5UUdhKUgvhc6VI+X7wZfImSsM8qZXmNZCjZm
VOzVoPjtMwoAQBKCMAZxQutCiPJHn3oQJqNKAUBRyz/rSpnjyHtnfcqGmzP7
zOgqOKTQ5KvpUpwimPjZK8+GDm6NGCnVschQWcy552gSJf1RzkVpzR5jTAHq
KZ740/kySl6w4QimQy4yzUiF4iqgqYEZNNZSPlsrxt00ljHoijrtSXCXxAoZ
NyW2U99DVBMhSzb9ydxPmYnOCFVosO4/hxg+Vw9wdzXf3WMts1GxIKnVDJL5
CJI3/nmcCgOMNiuwyGM0LwDW2qYHqByE/I9/puqnyu6Gcm7k1bswas05EJWC
cYRMZF2T9Sw0joujYbL1YP04oSy6cgvvAhjEZZbALuVw6zVHGuB90AOMDTSa
mj+DTYBHjI3+iktQIMXUBXwmooWTWrezyY3IGvnFJEZDL30xCpgMQYCVINuu
EwAgsUg6MKFP8TXrGIiwlr0zPSyGym9Q0b/lwbyFuwjOrQDp/5Fn4IQijHV1
uyA7rvL5oHMi+At0qDxhTDBeS2lqnZFa5tiD1AZ9vfEKsJmNtmWKeXFzhbMc
sekjUI6t943C1VT+Sk1kLgCHlkILA4+G/FdhkReEQ04LO56FkM+s4b5k0ajP
Bv/JsIK7NYQ39nD/eJ5ZE5GzgbOD8LreLHjRH1DICeSdGVmTqEcrnSAoPEaH
usEyKLhhcvCKiPTcYZ/Dx0CTTNpF8ih8fQYB+cz4/KCJh3Vgxrao4ywXmXBK
SecGAfgyyQbQY5iWMzqI1+X/AZcHVdXoQZ316Z7WHl7CxT7UFkVne5lw99pA
hTWQohQmVBZQwvoDn8TN8bkCHXlnh/yMEMyyRKSn1ppLfjHqJ3DUYab3yjlH
2ARFViIafmdWATxSSiNQDK+p7S8dB+yuVOyCjs+SUsh/+t2QajRHoVbmd1dv
DkSe7v2rFdEn6Tx4rGpDu6UA2wBl9AFWJZwGiI4R17X2iN8=

`pragma protect end_protected
