// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
Gd+BxbQx1y6/0M/krwgm3DMQ3LQqJBJEdAHmJM7lfJKTEsHpdyQwLBz2g2+zftgm
eoKEZK0D6WVswmHtxGm7xq3Mso7HpatmVcLUdyQtUc0DdhllBsK9r8Ooc6eR2Gb7
rkGdJnyFri153hHlvtSUkVoELuacNoxJwqYG27OStFnQMor6sBKDAg==
//pragma protect end_key_block
//pragma protect digest_block
ahNjK9zxM6hYEC5+gUwV1sqdfgo=
//pragma protect end_digest_block
//pragma protect data_block
M926klJ1PnMtnJUOZlnBC6eWoATcV+U3PJcf3xVJ8U4WtdJkoo9jVQ0RyzFXSaL0
EM6+SFLGxxfEt+NxkPfXgyIPc3fKSAB7HGcCw1EHUcBQK8nMPPDFIp1OpMRw5XWZ
iXFX+xPnGWvdGrTEbunhb3s4rD0n1Aqm4s0w6av4wA0oerg4kINIAS7xQMgy8Oww
F3JozYstyN3raTRhh6e+yxndWv0Xaucj0Zl79l9MXgMQYYwxm2f3dTlSdujuuTkm
KTRgMj++mlmBCn4NYLf7eyhVwN6O8I+sI3VzZi7wsbn/muCw5QhVeZ70/QfGf/M6
9STCpp+4rnEiVNjn6cXYNzzF3mPeF7ZYd8aLeeLwEzcaYucrHBZUeA0S7Zv2Mn27
222BO6a/1rTOUvsaN/khpB4SemXk1YUwSlhIqn8pcHTx99CRFS/fdQKkJ+hMogQX
PDw5DCjQyfR1k+Y0pYffSRYzR4FPydVDbpfRTegLFwzH60v6bGXRYO/ljfbmnSAH
B2TGn5wf+Orj4Rrco7mYRfH+2fPz5dyYzUmKf1ADeYuvZZ8AH0fTY7L4IlZgX7qu
tNqqW0+dxVE7R2pqsLzR7wjWei1J7B/RMKcNMyqbF5+27UxcJWxl3xUPiIbVw7CF
PYKHZLm56uuBqiq8W5CNyLdRm8yvr0+7X1OhHHjnG/evG8EMw5Qekk7RNmBNxQ1M
uNgb5MLfvM/2rDJBcdL3ibtQUItgu3eu9MXnww6FW7p7QoViC6LaxHIe+1CrNpDN
fUjNUxac1QOR5YaxTSP1OXwS1By5bp8U87m0Kkez0shLRjya5m+2ax8uiv1NP5zO
jFts5blu7tuVnZkVM03qFttO4XcekeskU5/zU5hyQ7j7AAHL8CnId7fOi93bs5f2
1rsq9Hbb2y/VX1RVPLB4dUlnve5XEK4Vr5Uw1FtI8oJsKiXQluE4d1Ko+H2aQTMh
Rqe7aCJpJs6YobFcuKwYdyVnEUi4WnZRsZI1kbJn1cuRlD+Fyl4r0QKa9eAxA/Ol
yrOggv9jsGyV9QYBzlcRMPRIL1TtnBfkytnVYH9ANHbgPJK69eATvyFJBnMhGEQz
Mo9tYjGwj1FHPTOJbkmowpyhHyKaE3xal/uNdmVUygFknC0AGpTnn5Ozv8fVJCzE
2BuyCGKDwH18mgyRou8njtYhI9aqR7eCmAqDcQZRdez0Hivz9CDD1SwF+KttplTd
dDXbcW1AJha220RlHj8zdQTXuZ8JL69pmvPLq3zA+8XnMLu7oEkRedpiMLjHFO+9
BoJd51m2VVUOlK6PI7hBw59W5JDZC/KQCebo/Bk8s/53UyL/LwML5PNnbliYr3AH
IhK13lmgvA4YiSaCLdkoAyuXo732zWBxtInmZk4XIAhJEFBwfBHLZ3KqWF6Fhtqx
2OCZdTTvXTDvpTderWRV4XqhHTzpZDtapgMTU+lbsL4if2dXHf74uqN+PoSWlTdk
c1cEwmliQyevkugZX/Fg+/HfJ84VxzqRfghK9wuJ5tuVE37HRT3u+ZadCINm0r8Y
DCwXl2RXyZmLn64YV8GRhXltJZBUKx7Di4lhP/GZ/iLxWyISxgdDZ1AkaWyjyRVV
Ob0CNRKkwD63r2HxAYm3oEuspWsNT6mHhpCiAOfNq+InpomEeQbAHK1ptxDytSlZ
+bufjqe1mw6RQvsjId10oXMch5hWvWAQe5Kxq4e0rawWFy6Zd6VTkdvE7tG18VoP
v2ACtlZIHMNyyFGp3jWxUtNnRvzziclNoUoJM5pHPVDhOQh/xPg85pEhB8ZfIhpm
advs2gtyVxNkv6QN7NJDxdJnSBrxWJsAbp4YNwcS5iHvyhujnxCF4B6GeMUcZPNM
nhs9VPOuTzKUcdNltvZ0qmpAWNZCJ2GtU1V8TPwzAFloJ52kCncg+cOb8iZwsf2l
UGpL0wYVPRlEDefFd83GKn8t1F3NnL40HLhtdPxs5X0GjeHeRmzqGOqUkKm8Sj57
gn4gdlQ1+lrGjUcDOcE9jd4+yNbQ6lyoyvsCKSQ1Ra9OMDKXcWNeRXHHX8c6k51p
tK1xTm7E3EQvO6wGaZJsoJDW5Fnc2daffTwaKVI25RM0q6hURijFm/dezNvV/lWy
csV2GjPGTSSO7WaePrhP5KS4tvOQrTWp56jle95XxqJz25Z8u4awJGi7mS+4REgA
YcyqUeuk3MX2QEuTnZVkbEjL+1n4WF1C0G6dU3i1UdrBWq9c6Z28xHOn3SCUVvK/
TPb+v20LmK9xwGWqf2kF181/Sdnz4BIpK4Ond156qZlFcAsWrXiMwnGfifVISMhi
6FuNB3l+H5b4csYUC16an0g6gsCNMIJhNAnw0+jSrgsceT8wvUhm7qN0RvmwZ+lI
yV8Uu6WoXLqT9+ctxhjn/XDcZJJXxagaaw2+PqlnxjfQYXr2XXPktXF+vDVHnu30
yP1jpZYbXAcRozulM0eVOIIqCeP/09eMgh7zcna21iRue7qCKg7hQ4zU7iZcZPVF
FhPkmCuifqMTH+hlQEt350HvvweaSbOLDecOpJjp5xPXvM01hwYCZgp9gB34zkDs
M3NR5mmf6oF7M/WATcL96mAinayduO24nqblrBTi1w4sRjzS3gfd+AoZSoZr+4ey
TZd6YGO792w3Frq1xCrBazbKRX51hf6wl+Mx3QjgquCjahIpoaOl0H9AWj9NRc18
V8MJWyjLHsTKYQDQT6ffHaCrDKOMaxCT0eLFD219X5TkKEV5Jljf2AZvlCFAf0zb
S7Yc0iI9A2wuxf4VoitGA6uu1GRiaNsjm9xeyH5Gwx/mPl89ijnoBiaUrc5nSO+X
ok2BqUVn3sBSTaS1nOYnVVNr9gWDtgOmYvj6f8xcPEyCGH2/87QYt9MgwiRFnMyA
0QOjMIAq3hdhhfL95TpI+cl52T1TVZENuzAUUzliXTo7Wg/wdH2do3brGmhIbIFO
QbCSxvzFs20cWiCrhdPmmqCPpVeJ86T3Xw/YeA/cTGuCiEp7r2/vowdTXx/E76Bb
0lbG+OuSPFzDBtG5Chs6vsWorH9V6643rvo6n0aaDuc9btBHm2nU7oNyV+3A3Yt6
hR/vg6rzMGfv83QPYmHqF/tkkTePdCi3HLfPNpx98jCK3JGqttaMYtRdJQ4kMv0g
bjdWhCGwsntjmt2q89GBA/uApfAiPlPESXTEY6e2Is7S041AhDU7dyxVUi74Vp3/
n5IzNZxl+oZa52t8PDPt/9t3PlMZtFtHIKi3Lx0phDfomyLQrWhQsJUhdCsrNMez
7IXfiJjvgd9ZgtiRB8xC3BTLIS3URm6DGiYVgdp0LhxyO0YarwjLpXrqCbtz3LXE
AQiWEWr3ExZZPiqrbYeXLDtLO/B9JeLgsGBif8guS95H7EWievDcJDXJcKoLB0Sr
AsgdxKiMDZFs1bjEntLgEeTJ/st0iOzP/v2HcxF1cW3xmzKVwtQBoVRol3MxNgQj
vPgUAXJvxXmJ75Xkkjp70ubVGPEeWgAhYYL5JRHKYdoNuGmcv+DQJlGAefWbMBtc
iceLtnroboH63Blhp+7o5rDSeDgjWTbOONq0aG1y8H05v3mV1sV4mkViJ7y2fsbq
1j9w2hfWOSTv/JfIeVka+Nj+MmzKxCRWlxjRaEZKNTQueHV/6zIyTlEbbyCXNOZd
rlIsZClu9JXlGGnaoRxVbYeLIyLJEbE6+F0ojLbpF7d41YwfVqoRESryit+kZ4+w
FVPWQoyc+iqummici2FZgdbeijUx8P23SPDjsDvPYjeUxq2pByUyl8o2Ur1X+1Jh
vhoeUQ7DHUaNp8+AP9UifX7ocJlCCVMrucTOV+OVIyBrNPC2l2lwaZnKx13WUrM8
uhciQYYIg79ZRH+gJwWg0DEay6NobZL/UFRJTRJcWY/oF1sM6jscqjCkUfaqHLgz
7iOwCdpeqq5Fhec4hdBNvTArVsZjZ5kyvw6wse6sXDIxG0xkoxcLBvsS0XSWT8G2
W3emf32oBr5rfb4RFbyYZMnMErM3vHUQL2T/8iMUgYgEKBj+TG9AbvrSJCYxjReU
7k2dUfvu/hVLXkKnFoHxqDv1zk2lJNCV/oyn99sKG+H3bd5WJ2TdetwtSx/xGJuZ
3Ydroe4Fo7jGnBLqKAZPEWbJJzjdQrx5Gbf0V0P4CuQaR99WgkJ12rJgopd3cRq1
qj7fAifn2p3CWuxUkNyWtTv6pcKcCJffnDIQE44DViXJKzAPVqKDX4nkgLYd30Ix
zNk71y44xgpHfWlL8nthQfSmet9TTI3Fu1c6HSY2Vqfvfu/uzVFB2dTMMRCNvlXF
egw/MG79lEEvuo1CVmCZQ3s7ncEcwlT5+5w1fv+UILheBUGN4o+kZL/DpKoAAkB7
50Af9EldMeQEQ55OyKjWFjK3bQ3l5MO0DmKtO8UghM90pbb2K5h2ADqXENt8B21a
EZNDrJQbl3FcsnBrCih20KQFucrC8m7LHy5nhRGndsLznKAxcz7PPukwQ5e1lijl
H+daE6wdHeg+r4YkDar6E29Wpz/Q9ZebhkrQCrPNFhf9RS3hzU/GlSW50OOQ2RsU
KUj2QFafPYwUZHL23cdi0txHs07+Bjez7BXftxjXzd0Qk18UZGlYCeWJyo70SZTT
Qb9uMWocBphykxnWbT8TLNfRHbgFxGDxxN/tUvBo/cqU5XsVABPDCyVWXPKsGo+o
rjZW6v3Z4c7BT9aqD651VQj9prCoHGhBRRVOdcZi7kGBla99ZgPS5gyjm/vWW51f
LYx6O1gI7Bu6seTaqBnkzzY4hRcSV+G+KBLyZpTgFJpcSDwyz9b2ZWgVnEjC257p
hv74V1Vgf/2VUyoYYMXchOx6iuZlwRbxgq2wHuhTqtjHlvWCLWFAJ4VgurXkfhMg
A8yCQLgmTWS8DLJYUxg0K8ahHsb6iUtnN+ueM9OKWoJE1auM9lWe8JUXC7nqCWzU
iDf4YxzUPd42T3SN7O6D1w+QCCCFxwWFdaHv2XgaOWpXjNsuO3ezTiC6/10RKP5P
hANras3kU5a+6VdY49pbyyr9NkiLivXsyQAA04LnEyIDaHJ18gzHrjzXNUu2YDue
4R9mDPCM1PhHDGScKENKqkeeO9aUObMfvXvQHvNO1BJTlM3NFFyuNDaJ28kDkyRi
B3GhkEzo7C6hLcuBxNwm94+GKt/UciDWqefTh8onlgCQpiSmIRTzq4E2kF9Xxpt2
u6d2pG30/itz7e8fWX4h8fsnHe8b3a8/IVYHSj2XfEmZvhXO2A3uf+/wRa1fbvw9
PdNx6+ANOvVAyxJ+dEvX92ngZT3vHh4ckSKiU9V906p/yWSmW+50vs7GwiIJHiSa
N4YZC0IIg7q6eDIInOjwNAO5VZwXE/V/KIUtYokwKHhjpMBW0uL++qG3v0oisFjD
9ah3l/4FIT9rxJQ8ER3Hxx7WvF1wndwzObBR47wH3cvM14b9RgI1JYSxZXGrjxXW
GbsxubgSrcVdPAsaRRY1NPx6Q5U4wBN3+vNw2xYYd+/HeEhwgPkTjwYl8TwMqvXT
IDj0/kz1jPGOfSyiLuiYUxKlzUGvJmIqt72GHSc9eiYXNo/TZ0Or9FHFu23+UofD
CKXqquXyhzr/JU6kSirv66iusgcBBkYSTd5dntoj8ohNt6LMQFXROBbkekkMyDWv
fqxaD/SHGNTnZYkK1GyAgLLZ7/ZmTlhbxAmQsGLsZNWapKkOKSQGFDe6oB9/d5pa
LiFFFldU6F3lNfATpYaFE63nJ2AX8TTAARIWExq97fDwVYGzDMjQiRBub2EtgyKu
BH2bZrCLM42AFLR9aUD5zmV6nBrJqyBfgpVzp2hR9soqiq0g9Jg+ibUOxGM61xM8
AH5HxoJzr/KzEerSLIIplmcEYOrMId/uvAWRqldXMjp8WNE/o96f9vP0SkSPtQcx
PyAOe4p3LSPryF5uZzYlYhpjx3bNKpaCH5rNDchxuIUCy2dVVeml4/8GIvUIsoHg
JHetw16pY8RxQ+UA2UI8/ec5fY9y6OYNLdzStWWPdM7NS1HQmHoc9ORxzL1AihUg
nJXSjhooRb/ceN1W5GQJbqhvO4vc9zy5eyeavmCMC0+kt7T0ZaVpuPsXQ7zznRv+
tlfyk2bhP/V2nLHlNMr53alwJnzQYmT9yyxjwKg6B3jTauLc+FfRuU6mk5lgZtU8
UcYqlGpQzpXl4/ARMB2oPdfHCvGuU1xrO9N9yjnVJJL8snYkDId2P4QzBsL/zLdt
0q3XQyE/Nl93H4lc+IFvwXvqqPNGJtUMmKq/i7tJdku5FnEHcBWSPjwlqNJpjdA3
b3UAyhONZGWPVIHiO2Icj6U+PGMl+nmDTUdTQYkhSvgWs4cyTM3pZ4BmpzwERHMK
CnhdtW8s3ts3lJh+8+Zc6nLAEpWzRFlTT6yldpWh4Md2oprkFvlobt6OPonbTC+O
xqimRCcW0rXz/2yONzoNJEkMDjSs8QDteNlIGPaDCxaxM24qWf+SD3mdVYsnt8QU
/AVcl3qW4tJMig1OwWCRp3xmy8vBUpvtBrNeWCo/QJ0McpSBzjd+tFWo+foX6W4u
hkni99yZz0wZHySFvhxLYbgMcFNz0Ewbn4e9S0q8OBLFP55QZU9RtZ1H+uga8C2f
quVYoZRZv7atIduC4KJcem5g5vOEGG9InJJ07asrcbnjcBIAREya0tOOkhvxIb3K
4QxdjhZ9zdFaeDMFR5tCEcZdliV28TMxLI/iXYmiXQjJn4EXAJufeRbDrwuNZTF3
JRiS4qLqQttvchE2yZiYqih/1ovwdYcdnksjfkd/3/2LIElAwQdqDwYCNsYzbq62
O2MrT5OAUM7pvPNj3Ri9qKd3xXcGEL7Qucbu2lnkX9XCLP4gwuFY5JVWqzqJ2pil
xSAQVgM4cPKweE0THOLgb9CP/gAVc50isLi2VmtP5Jse1fUMlIxAwihHBqZjcyGw
cCX/Gu5bDtRHqqhCIWty4p178mupzYP+8JD9XvhQOfwTmHIan22lw5sTvv7ycMMu
gJOqtGF5H+nwJzFf5hkzTkFcD8r+KmJ49zNFVtDZFNzyyHUnlp5D1czl3EXH6+B4
/Z15N56DwiuA1JxA2+6OMv10oPykDYmIVZ376Tzta4NrWddfNj2HSLKRHe6OyuAA
ZZCDFmgvToxBdY1wbbvL1psC7S6ss45LnVQPJaozdd9K1O8i7pSodase/9/Hdm3x
15l3ST+lvIp7xj3h2bUMQbolzUqFR+d5uJx4YTRRBXgDVmnhbFLXmVotntGC8acK
7IR+4uT9tzvscYv1+Ga20PuMKvPxnVYvFVph0m+vQ/kp0WSEGaSi3i3LO4e1QIJy
MUcKTbibe6CTsXQ46zq74c6xNCkrHBcvknKLlcxW71/HfSQX1G+JX7ccy40aeZqP
YjP3SOfPZZC9TbWj9wrAubb5GIJasVg/kKDxX9Ow+jshECXxU/N4xGyRJ7OgkPb7
zQmJRGBhZSDXtxkPNFj/28x4kYOX8/vDnMutycFwJWytPcZIRtw0H/ktMvWIOyFw
UcCzV7BWDsEMCNUj8tuuR/vKZqNiyUFr+K1m/zqmkYOso8SOr6MUettNIQGw8gdo
8fRCh8Dhe6HWPlv+WCgMW/9IbScbniRgIa6Ss4Hy/0VkPCon4dpATZjwnxLH09Pn
Jo8zBO5y+OfCV1BPqssdaQygx+u/rWjm69Khee+4KHg+OHXsXHkcQZkA36LquMde
g/s2R0MD0AoOSV2goaNVRfOgERyVtlGnO+guNmVdxLZf7CyKCdDy64WW7ch7zFKO
80LAKmVk+rmDYG6RvY3lsMChoOC8k3watU5+ZhOeP0GX60v5hOymeTtFSwwW+ax6
vqLPEYGi1D9eOZi6QHlnFLwdEKfVXPNRcf/P2K7SY/+m5tlAR/crmetM4XJbNFkW
SXxrL2//yGY8bO+73RGrP2YG5IrGyIsyJPEZHO+BA6GFmZCXTvpBhJ7oM67BKX4m
zHw9MT+5AMvhYCpCt8wiwayznM4YcR0xQI4DoW6b/CrRf/WTaMTC2UycNOPPvZOn
6z+DCrQ7bm3pSf+O70yVHC6N2uFEJyNVUOcLevWqRLobt3rR+X830p9zjBl0Pe4n
fF/4O+cMdN9K75gjdysJX+h54WEmbOnqlc601HhBX76n66aMG1EuNha9FeXF+8pu
H0y8EOC9tOJGzT+rAjCJAT2oW3UmqrvOQsBqFAYpwC/2Un+MP9Ry6f1GagrQlcJe
96mRDCiqc2Z8LNHiaQKNb32wdsnHi6k1NILr60RUS9RUVYXbmUWzjljbfLb4lkAO
QwsMSmfIaFx/Z2J+K2hsEdRXTjV1BSjsoAClCy/1WyJNcSmbFskOsVmqBr81u9em
wQKPQMc9sNbDJd1Xoy2FfzbXt/gqRnrqd+daDAr6MqT0gkhTHQYoNv1ZjNKTZ4sO
ymrNFRfvDLUmK+lADej2kiaVkLc1I3rvAJOCOmyoioV3JA7C+hP58jzDJwSPJDsa
6NlqFC58rObgvwuOCCwPCEG3Y1ZZbjeZj0GWRanEIo5qIHhtakIfZ6RrVbQgoQNm
IS57+YwJ3K8rLqi41/2KZURPfl07ISE0ACsHJi87jHlzsW6ZMLKNaBEEz4++8O4S
L5/UlGBscRoQ7E0fNELXHPTVKBr6vEop8O22m2+IGeu9PpLGt5cbcFrOWq7f1HMh
2VsQ23RNMcDjIDP767p5QXFpKhVKuitwo6equduQCmMOUraEx+plgEUiYXtoN5e1
czoa33AW3DHO0EZv4nz9+u0uaZM0X+4RGdcFGiL78N2RncwvdqkqmTyB4SnFSiha
7L7C/8flVjXAr149wioFkACFtu1yM8tyosSD1iDJ6EdOvMHksWtoneJY4IO4rmNK
OphGm3pti0PvmLxrkQ0dgOeUZSZ6j7YyAO3iIzKOMw+0eg4KeF8l7DdE836ZpeZp
wpa+PV+y2FlsaY/JWevbjApB+XOAsChkT+lF0ksfuMgpUfe0Vuw7oWvG3CVwcDg/
MFikNquLRwHp7kjFNK6GTuYTGKrSyJDe0DlbZuFpuPA7gyO6g1s5oZE8Wnl38nKN
IVNNupeqBfTj917kqRRyy/E0PMKzS9Vr2P84RDk1M6jSPpHet4ZkNRmo5DWdTCti
uJY+bb2XumuQL/6Z1VYvYbq1ii7MXiX0xDyKifNONAjFMs/d4QuZMve1PEVNgW2/
vjnySe6+ntjBPIo8Y1DiV+qPBY+13I0UWMo7vI20lFVldsFahUzBDtw6X5J8BWjE
WdQWzuAsaNOPD+YiLHvJvweP8abKhyxJ5pNldycj8nfuan8r2WeEyEKf6ZE8hmph
NUKlBkSThXgrM5OBz9ITrEGkHBRF9brP369RgcmFRoAAgL5vj46K7BGFUd77UFv4
FwFFJosc2/VcgP5Ewdtl3yQyJNfEgYqJ2nDM+RIEXKzn/BtUnkZ2y2ctEZY8A72m
zsZ67jUTgySw5SrRoATFSwcQjBSD3+cCFjxeYt+Iel5UYKuBKrzvFVr2ALkLIUTX
ngpvEjnLMoTnPlaXeRRmqaKuwgLRjZANMx07EgFsDiMyvNQRKgNuA2qU61q9mACp
yVPyQY+iqZAMvuwp5r33+XfjpDpwtzPFtgFjfRvCp8WE5CiFVCK5M15mqZJkpTDd
wZoAzGdoA8UiO4nZBvxM84s3B1ftBnB89bmR7op2tLsMMnTC7p2R406tvb/j6fIS
CynGBrerDtT5ZYJhA5gy9mMUL/qVLjG7CmMOSOGUOJXT2M9/kQV3EsNOmazx8wmO
VF3gFuEOlqMef20idwkOyr4tsEYR5gYuR8+YMjQi2pc8QQl8kyvqWwdVMpJRwGsA
fnm12iKPFIrVOl1WrYdnc5gzcBJoDLapRfUjMaP3rIKLQMBGinRkohFmoeOILbXD
vOTGxgnHDWRLRIhNzSCCKxIjviNlPx5TJxyHwGm0VHdcERSDsv2SbTquR9wv7CyC
VGwtJq8S4GqVP7RNRNz5gLngXi6R7hCw0TF50/fa4r46fvuXZmenzxRTWKR9Od1U
wF1vda507MM35Pn4w22ak0qwyff9i9WtFeC06xTkUCFTd79U8piz5GW8HTqzau3b
UivGfwXv6adN5CkhKz+NxcFV8iON80u+YLW7agO4JG0MxZOpztCfEDZQFFDhF/m3
6ufw7KTBS7VI3dfGYACBKFWOTqt6+PPaOMYiwc2HXqPx1glv24YEinvJZhIB4HGA
CFcrvq87CKkQGDfQoPMOUZ5Xxwmd0gwyd/7D8uFZfGhgwkbkVIevCza372gKjbTs
adDibPdBaRWEW+ZOMnr8z++FNEr3q9wSO7ZnvtYVhg7uKLBsqVUEI+qTn+hFxHV8
CumSBjDBUvp3tqq5/ot12DGUBaGQaWhOPwFgIx+Hbn4SRXwDzBF1BOFroXh5upkf
PKOqQ3lNT5W1jNPlaTvLtgpXlfAz2v0wfwSeoYHFpyU3Dp4OFFwwbk75/3WP6lLo
yZn1mhC28FgWDGIIOqiMJ4oML1MsptdHML8B/ekRuTJ/1nqymLDO1Zv3zqwwapxs
BtUh9cBMW2sAzMTcOKpCqVXtaJePK8x616EYz177eRTJOjJoMYVpvk7I+BfQxWkI
LIkAI6lgMhbaQaGtSph+cfyqJFFr5kPzUvoIJNgaB5YJm/6r55D2GMqWbzMeGknn
WBm8YlCQlGDSWrkvLqczpudPfqNYvXWn3vnsJbyvNWd2BdVOQbDZwzubzN6hlS1n
lRV269WPORa6XDaVFWdkQuizkyUosUzvAtiKm+cz+S8Pg0+C/Q7eMuOxkqtBo983
ZqsRIsovqcQTKiJrGufImgx0W+JPkZBjzEjJr4rfbaRWtiDZ6mB/HMh095iP9mS1
XhhRKa1u8nU++rbPHnd1n+a5Rv9Qazz6j9/cSD8qSJ0fM4s4h+BdbxG+lSFEzpER
HtGW8mbHC/kB954QNtt4VeqBJuA2WBi8veegHVtR4rwWuRbFcGGUyZp5aWydEwWY
BAYjTx6V0nzwo3Lx0zniTyDNCwDbMatKEA6+RF71zj92oCkbhueV3y2XIxXfpHz3
PMo5NGbeoierRMLq+nLSjNk6eu25P2b3vHj3VfB8+JSQ1oeZz5v8d48JHj/yv92X
jDUSpa6fzZQSeWDk+Mryw0BMtXM26XfSc1udU6zYKTJiQpnMIc0mMXk/66fv6jT1
R+MfpJBKAgW5FFYvSOgyGUBvXovuokTlL7YfMYwD+PJ1ep6O+QxL/qW2EX1lMXx+
zd+kPxcy8Q8VFhPhKBzBpyKOF1Z6zwf844fCNNBlS9WP7TDjppRzkF6qJIjGuZ3j
w+BcN6HUWkANAQJs6S67gpvwHFtVxJiUByPHkf1R9JrNzbwaccTpu/7ec2OjKOpL
dTNuzifpZw9T5yrbHqK7WqYoPgtH1GtDFRWe2JaYL282pBj6UnJjRQurmRl0tTON
/NUAkZplq9LsZ5KjiZqS+XhjCVURQhkmozzxWb04GM7nzdyLuhN2d6RnPWjKqyb8
ojX9lMAe4oz6K2Uo+pyZCkz3g4NQp3xma1SxuUzz9yhWktrx/ST4aAwjGMQu2qkQ
1YDuGG6blt0Pxtsp/svuXqRTSYa0vpNBpg4Ilr+pgvE28E0yNcFsvVgKstlrdQ1T
q87tI+KXY8SmBzyBaxiR5qQo0jPz6CmbAddwWY4pM3Pzek6hb4OmCmCvLYauE0zz
ccdsfNAL2lO/2AOt6+OqTyFp/Qm2OEJCrTxzKpuv+SNS49kzY63Pjq02N/TXPU60
gGA+QTe2zLqltVR7TeMhJ1xYaGMFV3A8M2UvjoBiXgkPACJvG8T1nYYkvjST91m5
jpTjCw2dzSzr5vj2hl1CX7rHpXclhk92X/hsLOfRxiZy6rLnjPgUJK8tKrbACvHv
23WAMn0TtJ6FnMkZZLmDtW0iK8DViNIKqAACJQxQEGutj9OOQLYKSR3rttSip017
2Z75FYTKXPIbBxYFmoruYS+qrwgNzcERAMQNqhgFPE4RNt9hEbmmx8W7Rg5fSG8V
3f6sA3b98e28U6TkHYVvTv3a+hFHsUCkbGS1peLZzosCsZih5Xlp1iduMWNvmaYn
XR1RxYCv5Jlm79p0ZFmpHQ04pz+ThuW8mE2eCnhikJCtsJWEVh9wrS5wc+pW3F6A
Vpc0kliTCCwvqAQFFlu1JdnnWRNKtZzRC3Qik7bmodBpoIYzl937CwiooUZ6NIFQ
/E4s1MRUF2fbdTXjqIYcGOHR2VF9u0LfIbG4aQ0WSdhWcojQKcMHkZ6jguHXv6RV
WapD+bIY7ZzjHK6V2gslG3B1y7WwYX8/8t7gyuBHTDK+oeO1Iomo+Db8YCgIsqHh
zOOd30F/KNMP5Sseg8SPVUp/FRENmy+GhOUo5DHMgqas/hYB3pXTZtJhuCUdiUoQ
R58j7XbNKa4rAMSIYWN4q1rVzZZggPI9C80vfDfLZ6VUj52LyT1HS1+HYp/KBfw3
n1uXPMRmAWpYnhM9crF1i7q/TuS+bLUjHrwuEcgQ9OBV2jXF+2s39K4E0u2BpWc4
gj670GVmZ7jFZQ2tKVZmzNggUYULGTUJUuBq0tW8OxYBFpocDpRwVnswVT3Yqj1d
Pfh1x4lFL+QNBFAjBs+ked/y2rdP+hyqjlqh39pd/3VUW4Bgx2T+XX2BZA5wuIRZ
Mfk4uxb+3VkzRoSUaydhkKZwN23K0u+Qc1B+SvETmpy1TC9xbved/vJsFqM5VxCC
yHSMqlIUEJkJHHah9e1Z9VF8+peucwugxWGCUM5CiuBG0bLjueokpXZt/U+QT2Ep
JC4lCFPZ4Y+sWKWszZ//09UZnyOyiGk7lV1xrIqeRqXwnHo/uIfnPCgxo+lTcFAa
CtKfDUxVtIFxR6GKBG0zhXULoz9cFDwAYR+14otgYDagh7v+ePJ3bJBws+1k7sxD
rLTfdXdcJzUtadoHsHO4ya8Y8nkoFFtfo51bPFANveYiQ3E7CMIBi2400WpPfGH3
l2p3tCJuWyhDfLMwaeTczdho4+jDPueUw5wcBnOkPk2/8xnLYZ+aAxCwnnVBG1ET
pF7M3JZHqoaXSnMn0TqvQ3BTsevv32yHkIZ83JRZkzMWrLkFM7WbJnHLEFz2t+KI
TpqcrJOlwREfnm/7lMF22KXV16rUdUpEItd2V4APw2fJmu2D85Tkre+O4iOtev3L
9yOKPTdi9gzE1zMfX43FxJSofGTGvB7LP90WuboUr/0rA6X23SfmvhkaQBqkzQWu
pkLUONlM2+Nk6zdvyK8KlCcsR2vAWSCo5xC99aR15nnwKKhrJJP9Ety+aDbMc+7v
Z8l2TGuSVo4dSwKhciAhZb3udMtxD8QO3kTxrh2A9VsdqPdtpQQJ9knAyxnKUU43
L6Xl8sB2Pjs0R7ZEQxN3N6rucNMrAU8J53Af1gIw6dwlgf1Nm0g7TfWTM2bOoRwl
NAex/VNNCzbXWNBiN7ESFn5WZHoyCgG1f4n3GBSGJEx72dNhhU6fKC/sPh09P72u
ugK09O0KuP41wTY9mDFj1cqoFL9ou07F5YP28zOXsMuvHJBPOf35r3fb37d0fwXI
CgxqwabrxpcoHy3v9ckKado6mv3AGz6KNuDiOjZiY4zEJkaKwNidqden7veuXOjB
psAEc/8LXfrVyLmFH45g7avGY9kPUTF48Gn686cemWyTe18Q0nyad18aIliKange
tvc6QioFijR9M6dQJcYIzqXuRDDwxMM8R9Dg3NrifAobNC1/AC/O+cR7pbeu5zva
7Kh7m/E2ibROFYxmxTOH0hAe3iSPoR8bPWwWCs5KMr5oQyJx0nXhLSahfRDoqe05
8NCWCCbYsV+Fw27q5G3x0PmMUsnR4WvLRIUlZbMPfrPpP+ggHY1f5s+KcyntctSw
61EeJn75IQ5tZv1Y80GXCpOTHwKsiVTkMeggbPlHfW3shbHNmYLZYV8CMoqP4lOk
rOJ3T8yXP5/fbTtGVIpirIIQQJh7cdZZ8fYozu58YJfSCdLv2iSpWnkXAxLEiJEl
nAi4ffqkVsq6cBEXkysP8t3Suv2YKk8anIoe/9iCbULsjZhd2l8e921SOBW3GpVX
q15aF+UzOBHafAESfDY0rKmfMP/rLRvQVRH4duBpiyEoCLKbLYP0+R9WsRyobbHJ
B619yswVZ11J8KUj0g6jucn4y8XGJX8a6gIUjcp7P+TG4TGHmQb2vMLtN1Z7Tx9i
jn9B8ba1FzkLWqzEys+3+axGNJ3qIPQO0sWACQXGs12IqDHSLXP08GNqXSS93xVG
B7zOVd4QFnWtoWO9ULyc8nSCYZZSYDybMLCvIVedOPV/A3MPwl5b7kM29NQ824jL
z7BdD3YtVktxxslDtTOYmf4l9Bfgnb5BPmkct/r25mkuKlNwfqgigj7hQatIncfE
Aj9gAtwJ4o1MQT3+SOERbYIzknr0hPO+R2atq7jx1nJ+rlqCOmzGdm1OE5BbSka4
PI4yMV9WvOyNcWw628XjRU7xGwCK/YKnDg7WCocv2lMxa2XZIu7VJOtrZZ2Guwqe
CIwhGjBtZi14+ckx3H5BJc5ahmE8VCWcdoPo6Sr2B5L7Q8Gk9BwO7qZrN845ZF5L
oqVGiMYyFkJ5GOJOjM0FQL5Hcu8Ztgyp0+pmyzSRGTddjFTMD2AaHS7ZB9PrD60T
O46kP0AdFVmy0I3F+HMgUSaM7WICcGTVd0Q3Rm3H/sYd9QTc9+M7az8536YVIx3B
bSAUraKDiF+M8X8Ezc0rwc+TPCwSi8Hn10Eo2TflEce9DHK7pMwyDhYXzrdrVFi4
DyDeLb+FyIk0kJrzhMXL1t+TvBLdsgC+uUCPhm/VZubQ+S5UdbfPqL4oZMVbtdCq
L4W0PR1vUkbC5M+R7a6HJt87rN2bprFLS6a7DYgpIod4kTZXYk+Y+Xrl+VmFtp+t
J/dL1hslqUB0YekaCa6kWCJKgZ3bvuWQ/kTx6XYb8IXecmRQqsFKNqpTIoctDbdW
z6UhUT7zcWMCiLV0BTWHKJYPK/PqHWwEhf/GZab0QlUPHq++QE4AB1Cx/7+jqidB
8elEe7RedRAFWAIegjCdHSLwIP0Hls1ry4iWbvwhb5u84GOuNpwaRAOHB4dITxiS
JVCNBn6d+zV8/by0Vlx2JMucNwb6VA+vgIl/J9a0MgdQjZak96EyOZFTxd0j/wU4
4JH5njt2bRBFspwY1PMBvfpJEG18va25RsQQBp6ScxgP7qTWAcAgNfxZmT4+Nyqd
imvGXvd8OaUC/Kp/ztlnJIiQwivPgcxJKVRqm+sPMhPo0Hb5QAohn81Jo32BOQE4
34AU4Vo95z83Bpx6uJHDf9KsVB3dFMWIOBbuCeQJAuFzarUP3oEQztn/GGcZIBHr
iChmvTUHUXkEqvSGUbXbRyfmbAQgvBUulSdz8RLgAilLXKyjmxZFzVSgRU0uhB5t
vbYnc46feF8byPBT2ffYtDPFQIfmxzHu/NNg5C1whpABzZEgE/LmYxUekkhZyZCB
9HwTR1FsttP7B+AGvUFfT1cVkomZAhkLJTkofCdndXa1bVC7wI0NiOfjuIEzDIFD
h52gGt/5WEu1szyjhLFIWj9eQLf7KR6jwBvBD+sJ1TsMZ+IgraEOZcqFGhZo6naN
EsOrSpmUf5Lh5T8vpcDOwyp1lQwrKd2CeCseifoWQavDRONrx8L17htOnnX+G0PC
n4l4lDqCVWQas58chDVV4ZR0OXNIKm9w5CoVa0y5FnRTEFA5lS9otiASqmVg8LdP
rzXwNXHPHp1QPmMHqxWESpOVko4vTL1NqTQCQCCscxAY9ANzfoBOocNSpe7+UIzL
T9BLmxAFRbGy4M9cvtPk/MBatu8leYICuef5ODwqo8KWlZRaUddV506wymgeYnoI
TbRJMmgqmeRCLBHv21aa4fFIgXHawXfqYCa1VxqYr2gV0VQHlEN8CQO5G3C1iGwH
UyxHrLOzTMA9o7D8pjG/OoTqh/bBPULRTctrP0u75mVyxzwes5/Ag9QUUPcd99jl
Sud21HVzIzZMb8wlL5D/wOJT1PL1khA7F3lbVEgH+jPlHNeX/YsSeyfLuaXQ39+z
l3NFGecFFSUnTCLfuPZzMhD+2P3Sr6Xqd6ny3bM+uJ6A/nm/rawUN5FSKyUOf8Z+
KxtjPj9JzlyGQw+Mk/88wKYsGYGgD9u5vB3LmMcVksE9xwKDDZ4M98GhI2hUym9V
mINf6LOZex689dY+7DLfhE/lZ9tVvKzXQksSBlgHAPyil7NE5CmsfyKzVzRM2j38
lG+D6CkLiuarSMfk66UIuVz882pMmHtqr6RfYo6+fqmGtanyoiikKBQHzeIhHrzc
Mnt8a++PhNZJAapjtxEDj3YbdyGKKGZ/pngeHf6e3dgzLgZB2DKwcSi9Pm3neCeT
JBFke0NeLcqPpO2cEyCP7D80eNIx8W0g0Gm5T8xUpfeI2uhNKK9JZw18RyxZIhnd
SbLZB4OYdNCwM0jyazVPWglApEYqLjd7xO9dcdUKRbnnYLkxO65tgOouMT6cTK/j
BawTgrMFZyXB3GyEKo/bOlnZO0joCzHdOXOXx9TEMvIYtGq0ins19MkEOB4SzWwm
80QG4O8eWg2qzuDSLS06eaAGrKpTD0ZevbLoSZgVKIAc+ZPqLolHhl8l30pCsnd5
YUevLuLlgXdeTU61rrHr0a/QujWJjYMjOX04QgiJyRh1wzYGgkMPXBDO7SmqahK9
GTC7tDgCyJkbS52t2rUgaS4QA/r6DXp5QSryr8VG4j5FTkG5mut83OY8kxuSTPKy
blE6nZjsmG+rhJk7xSXmKRKW2BQr/jx9AAOM3LlQIce/xgO4ppkHUufGfRqADlnb
Iaj+zaVyr3QxXPuXK4085CxAxhBxmk1amHs+dY0F6B4knLX4nlliiArbGG26UYen
sPcZ8TprRld5RUa3Vqb5m/LH1jFOx8puE18n/JR+nw5T3FXSWQ5kV0mF52o1VcBP
XNAocfHXEVMxmSdHz3ZLmDwUKU6tZsdoyDm7rCt9I3CvblW/nS6aWCNNqTwWwNtw
PuVxEr22OjzFqeIqjDWtGdBZfcxs/pPpyjr91165Qrp+Ewsyc3NPlNcXM23MZaAc
RDqhJaxG9va34edxh48KcOfWvT9OTxt6Tq9GuYd4ly1DDHZIHa7beoJ43QawtMqZ
yXxLPty1Ecj8O0glAAoII2FkN1tpfTEp9J9fmh5FbYNae7nnEGxIZ2hj8/R1sGmD
ZYWfmU/oxxAT4tdrh32mkLeYJN8ryjCHdT2eNQN7XNEm9sZoWY4HWMjf5Q9tFEN+
tn51cdal3H5ae49wgMNqFy70LMuTrvPlwgX6QGi9m3srj+OQp4Ca9dHE494Z/nmG
zIfOt/uvQDHSJZd3/vNgksxOB1wgxw9GeQUEkbDN1EYV/BYD21Rk0MTVSjbSkrAg
KUlZrG0xvDJWpwTSBuApxryEo+fjVQ6gQVIVfBl9vVbn7n2ecSuXRaq78KGvdHkH
ll1QfDfwvAl8htJRhA2whWjqSomStGtL0Kf6OzUDriHjgwNslrgAlqjPXsLCTBDg
4ptHe5pFNnErhoy9bbSmzYrjIViBx/pbUP/XrIt98BZNFa3FGDCvqFV8zBSL0nl5
vo9Bs/aG2YsGJXL5E1m91Y6GgxeiUFKCkc88XMk6Tv3o0iWLQCHbozP4rQQWwdBC
wEnQUrJnZE3w8V9Cr48n2hFHp4khOtXotSJYaC7ar3PIX+GcipHojTUxjBiCF89i
OBGGu08BXKX0teNuhuQR+pEShgC+FMfcdc40fiGr53leU4AojFyqAFti1f798C3K
5DPw2KRJKMcyomSnNgh4zCDSu50kjbHirpirynz96Y0ZmoAJ8sndVC71z4IcnXvE
FU0DBq5l5e3AZUEM5io2z0PAwFYs5y1j08DPc747wFuJd6qwgnxX1TzrEQtXbrKh
xMfe4Q6RCp7MpADopSnsLWlJUjTjTdlNAyRmQd2FM+9D4KgT/Ohs/FSQ/Akerkh1
C9M+BATVGt5qFY+UE/KsiogYK2rCM530T0bYIT69Lwtv8Od2PdiJcFwIv7dn6rLR
qoKER9QqDggDJCdprhafIL1V5XM7gwjhy21yESSflBqDRZsb9TRlBNSCJAAUeyyO
RgVhTYQrbwHsz5YWm2kVWLg0/blHRSVETy5Oypw6wRSTtG4wHxkmkF/n8RSkl8bl
/+RgtWOn3XuaVY3CVibahbv5SSPMtV+gQeQquJMH4Jpa2/3ZwbsrbgF0MBfIMHXM
9MEDLmPcwc6Q6NejhbZuaIdaG16BAMglb2O1sXOvAmIGI7RRhxX/9PrPjVWSoI5g
Rh71Ln1i35lX2XC28s4qVOpNo/RQkzMb1A9ttUBxFQ+9VL906A+JwyERdsWMLJR9
zZsPjap/eljY1bbpqmcQn7cFWUsjFaRsLoT7xEnRoCffkdUf8Hf5lgKASGt9VWfG
qYXl7Lr3RX0tHPkFy7YVMaRGKUlPYIvoVwhRQvK1iAAB0ZlCqiZh1MpHCXydnR5j
jgRTV4fK0eh0kkRjQvJ9m6qZdflf9Cbf8hzYfv4MVw+jOxx4nHJMVeDQVMd+9H6O
odNvKKPW7MQIkVFfxd6HLjU2SwJgEvYecYMTg8YBwcanb7w41QH7lpigj21fNW0X
16h7OHkpgF7fo9qweyVQ4Ykhi7O3BDK31YFipVUS0pF7YLd8Jh024lzvxpsxbjFF
23m/qAfHThxdXiOq8UC+rvt1N6q96wmJau5LBusy/VkcNFNjhBdHvFWduwjSc+w5
J1xdV9jMlE7GJifgJgK5JPCGjdjpox8QeOlPAI8OWT0qQvV3W3evw4KmMjJeCyzx
q38ClFpjnZ4feEyV8KbD0wBYJPK8tDrfoB4HBELU0jLgsxDcbHRK3H7laRcJx1P8
9jSd3AgaftXoZGVo+MJEMxRb/ubvw3skEGRa9zuXjQttQaFbM7buLhNMUkBY5sWR
bwSc1xSnQPZq6QsYgiRy5szWRpusE19J12BUssxFUVsPQ3rkqfZ5qZh8isHLxlx3
F6G7z7IH5hVttqTIyju8+PG3nYe6++pT0MHsFcRA+IoQYzaL1SRBUPji2lwM6df1
9b6oTawkcF60krLRaTvAoDYpiXFN1/6YqTDhIZ+jQ7+87YEzf+MHZSay3+drcgl6
epwU5+w4GcZPutqV2eiwbU+eCBkwT9Itb0OyS0XRJb/X6ePpyELGzCBJWrNwvx4H
8+05XNkFJaJW8T1GAariCCWH48m8xTy1bj3avG8EeFlf4zP7bAWFEbZWcHdG6PNW
92WrRGEOsa+1+9WlkA7mWUBqzzEOuHMC4PHAr+ze4YX8obu1dHO32deN7+bCs4Xv
3FfPjdq0zxDYrLGLxNE0FO20jLlELuB5EMavdYUocgmjmLryrlJwa9rEXS86Xc7k
XjIzY6J5vs0uAV0K/LY460lBQeS5YLN++ymalg/am7tBPIaqA2PFdNwCl9sRCbAj
TCwWu0kG8Ew9yFN72CQnNEWqO2v5+EwmphR47LIO7nwMZA00C0YGQaa9raFwXG6w
EZcTwPfUtKfHuNiJVWMFrksdnE+9w3P6zBnKg5xritgo4cqo9ViJwCvWes3YFTds
y+wAakZOVrqURBDxKMfw9Uzp5KP124vHfg+/ggpexqiUNfsgRJMFVvJwU/PRB03a
xSDtxjIujPcgrExbBnavlSNWiwi7ymqQrAhfHBngwPRYk64ORm6031ZnfxK4C3vb
xfkMcoTt1q0kgLVLb1vobOSsZGGus+kRYUsLYtuygffO9R82XKxGQQstxATe9UsV
oRKyWlsOWh0jecnLLHr+B0RnD7ULBEiccUbRR4ZF50eewLxOE7ltQN5Uhe3dpWbV
76UVXmQCSUZkEHVq4uy37cO90NJ1k0voUYUhblkM67Gpwhiuo97ANZjm0WZS3utV
vrtQLVPRnEg/Pn5CgAUlJq51YOmUSN7CJcfROI7Du88pzO5oaVDuqfZ/yfCImVtN
dcfcXBYlWuiWXpXHpfOQ6wE8cm10L3Sz+UWnq+WUlwnDB0fEDBEZY+/EttJtzCNc
ATIri1zVPRBRgIE9H6JkgroCCbPnHOHSgQaD72NkvOHtZATXmz47gR+Li8pr9YNu
tCZtwbtKRVzwhbrydYUPphEc9c8clkSN8jpm5SG/KB1kzfsVD8SbQCL5tiTBfy6F
zm+Mz+lYB9PxgJoeCheMZzyjVnFhRhGosUMRUguAns2SphVqEI01JWWe6IJfk6Dz
JShxWz92fFibwjpTFoSvqDB9sTqz13yGApk6KTSx73AQKH+jc/Msla67DBgceug0
Yv2xDwqOhX7wMoCUn0Eb4Mt6Ba2EgVogyrS02inZvnaao1YLKUXPKqMFkDE/M5jH
IOCZka2Wxibh70h0MynbsfWOO6x2/quUpGM8Rq24Oa6HfQDCvqWJyaULdMD9S6xX
n4Ylr1BnLakxMbKtAJ8XU/q0JZFXAMjVgim5K8S61NkmQ/ZyF9ZRES1OTpRjZdd9
MKUY/E4Ak+DLFPJRMX+y3OM5LJlHeiLnNRqxr4Lh1VJsd0z6raiYVm98S5e1Ep/F
4sHJBJ7O4RDspJlTDl6Dlxrl6K51Jxa9s6et2gQlWoZjOWcmUpkxtmmITCwUn9YA
IEfgi+hE6fyFZKk0tXa2uB7RbWDKrdDWUC1CCF9oi5LUuc2jC0DeoUozml/KBOVX
U7DO7kcoB6tSsVYRwyZQGgx8pONjzX9xyW+BtP5scRk4p5ijw0vtILWOO1tHDP5W
VglrfEB9Gw9rIRISgdLJZKG0CSvQCcoIBvgKPbYt5gUqYXtwWfpdMb7/NA/YYGD6
+6OtKZNIi+WSrzdLGW14cgJxT4rzqVPK/wWwpncZAqT6sQFY8rqDgJFkJJtj55Gq
nDu/PVt7o7uDaWxBxhsTvk9HovgPqVhTf6xkbgha3NVCkn/sRmBe4vt2Z3VUfy2V
cXDTZzJ+VMNrDpD0v8hm7W34LgpkIC7y6mPDT99B2Fsua9PuGDDKZnh/oksukHoA
6kfetlJwM8v6bVo8HHJkMFAlJJqXn5L+9I1w2vhIL3xaHnJ/zAl+B/12S7TawP6D
mruNbfwpuMetzk17MzUgflxwjs0FSexY+qxctXFqG2ws5O6sL++I65PM4Gjiqizf
2r1CsQNhhaM4as7dhA8CP0V2lwq8ipnxNR2SW5wR5zmCqEQJpRVCvJXOEMcS2zP3
GOna4LEMPc9J7qDTPdx31m7QvaKsZgGWYk2M43+EHw4azv+HexAFHbi4dE+9Cu2B
v9SK9T/+NrLzczGeIVx9xB8/zslWSEub6CmyYGNUjxWyxH4uvczG/IBXwcG0rSQj
QJZOGCsFre/27pGBezQxOxGVVY9868b/Ix0XgLmPCM8QnbjFyW1EzQd6c+N4HCH3
YqBM4fGigFgax4mcHGK8foe4qy8IfEn0E6/cgL3TcA67HXo5nwbPdS5gRoJw7wqp
IQOBlKpbvB77zMm2Xr08CbpSninIdGPJN1irb/1ATHO+EWlh441B5j+vHm61mFkM
8GLBx/YSd4ssUDJdlsu0Y0wHF+CJTFeIsd4PLW17tkR4V590hbOwgl6DaLjor4he
Bblti9fl0tQyS1Ml+zoh+s7wdoD/nwywb6DvIk4k/6EtHByanfJx1jRmv5S3IczB
2Td285JjoAmR2qBVOWmNzIZnsJx8qWCsXIiydfmhjhZvCsn3QfYhd2jMflmCCg5k
JLtgOX03bKGa1nZt7jdWpr9Lh3axxDk/dm/7GtAYaKw9+r041pfvqkkJQM4kFr+G
dFbN1o9cmU5And5/w+u+cFkGPmbwEz+zobvSFT4t+NRU1nDYmFPDG2Jr9or5YTpd
U3zpeNxRna+jRIabR3bzftZtbCeWwExiqvtDmMkmXBV8h8zOPt0S+S19YCnyfE2E
Fb29xtrgJRpHFGUmBkF+LOHiIvCqXCOcohn83/lflLbeGHS9wYUtV/l4Z3YOMuHO
iX1H4iRVx5YGo73jaJ6Ji0keRXqCfD4Tf3IGGX7okYoLWZ7YQbk4bX1jYe+60P9u
3sA6RyL67gJha5xFzdnTzgm+dyk0anCRYc/ojll4V5Px+WQKDfbEbvH9dLhzH9DH
dMOxzarz/Nyp2qaanueEX6pqh8tCWNgTa3AoitcW5Uo0YTeROoeCYQrY+Ab67LEh
8zXADLq6FrqpQb2EhuzCxypWnC7eGBwmUkypGPOkKEDGUmsfuodTr6OGPwgt1eF7
5B525n+4uld2Yhc4zA2eVByZvDATIfpdLSBAWE0yeMTRmXuObb9qk8jJc8e3hIYl
cdXqzchxjh491QHsGWzn3Y0iwhM+B/W20T13BJ1foWcZBSCpfq6f+TlnW2QqjkGV
gVyS4JRsjZoah070NN+TOG7lWLjQ6+RGUEyWuUxkFNJSMzDfAHwpAFnNDA3tyxJa
yQagp9aNeeaDo83TPgZuxImaZQaI6TitZcVU65HmWCUCQiibCIGZU/Yks6b801Xb
oDQW7QC5CwRTnLpJjIXGIt+BVili8vx869P/BZra0koCp9o4/nRxW3AfjBqu5hzJ
9G0fcbyrg5NT5pzfIFLJVV/towVuEFmmUig3OQfLQDFEarqLQY2drRCJCmqbxXOH
EkSHSxvULat5xmXEoc6S2kAewP8gPqkontFVTtRv4lsruYfD4k+Nj9MqkWGZhxTJ
Wc6SQATEK0+1jAGoEKStj9/siab1IrmH1hlH6i5Aa7K/nCEZqQ2k5Nr2HttitpYa
oiZMuFyTrD0hLKP7HpMcfaM/C1eT8kJ4qC2sgaN2I6RjN1YEGgmxDpAfQSZ2oVm9
XtOPl9gB/YyktLRew8CTBmMSrrrOE7pv1jgFf4mCON/j4pZWsUbmpz/p8hkik9af
tEtNX6yQioowLOsqfHTimRqhbbTmDGaYVRZ18p/tYbOyKqUJzDzi3SHl7ZheTrkR
6vBIIcOXoJFfKSnKjH0/HB8jokjv7xUmqU4nJjLoAky5YHrJrZAyd7q2E+kQN1eh
tP0VLf3S2ru/uGyQPt2VQ6I0+MApOmW43uXwyynTX8plRodrxOMW0SAW53O1Kdej
MRz9lupyshz3WHDf0PY3krU/eXC4AgZlJx5USEMLF448akg+u/KVGecTEKQtH5aU
ndUSubJVinfuLR4jdfvJES7Td6L8WnpOsTR6+XedBHWF7Pnd3pGwn+IjG0/wuFSd
BsANcbbhphmHRsYq7XlGebzVJEOrLW8vJA0rrPb7XzsJR61pSKZOSsaeka0nSXAq
yajklSy7HvLHC3Fm6xG7jZUC5WOkU6tbEkc+Gu0YMbAEgRwDZ3COqXsszDpsRx6Y
yaWAyjiupSD7ibQF9ZXKb0iNjEdpxoJmfFBKOyC5ZR6fkb6BL1OAc0BpsW33xOpT
Dea2QTkEAoUPri+vIchsnz9Ze0GWaqLJKeVKVT5EEu71sh77v6VP4KoSVsc1NKSZ
4FlisvHrltFF0nUUzTScmo/HyM5fgIkMxQN1x6rhnA/QIn/dQWI+/IFdchtJ5Vng
ypvWXHXG2HZF3MWt5Ao6Q/UP4p7CiD1fJ8TW874wS2ARvaoGaIU9ZG2zixOtE6+O
ME13108rK3EcPi74iGesLOgAELHWyzg6HhdGdkx/junkTWuQr7Ftl67qzW6RfEjW
nV9fj+TGJXZrO9j1b7mDmcJO/J6hGN4vwclLzu2oubtBKIOMJLD9Mtbq8Rmeoqk3
2wkT05wlGau7LDBxVl8GLI7+9PhCQfDTlgvW99KKRRW2coxEG2+doakvOuI5wc1f
dLkOsF12/R1OyeSRf/HzCbRYbGSEiyXKaDdixuY+z7Xa9bDN5dD9nUU2AqbQntcs
isRmJgi3seVVT/Dm+HdiEHC8QI5Gxws60DIHpDf2exNl3/meaB7u6hdW+mXKDduZ
wvEQzF54seh284UOCrhg2uOyEitY3Gm78oi3jFbEIHpajMvO7rTwheSjTly04bD5
RVFjakJ9fBn1LnfgVNnE+AKd+z+81fRVPmlMJbng7JOjfRMyGTaEpDH/5aMmh62G
e3sgV58sF55z/ZNcIbUuf64WOcxiyRvbbkujEbz95+rDdl6wIcdhqAZuFfQCjtRa
4SagpBFHvRJvUTdCjdNlrpzpKOzPLAEZI5fYv7831klNNajlCRgCPhDxfvIOKK1x
bwRLyNgp4AA0spBf2cu266Dr/+xyr1y449dBVVO0s1RLlMZgEgaeXNayJgYqsSxd
UKAexpow81LVua9RI9RqkZBb+1cpwoncmabfzOpLCHu8V68qrhkaiXfmQbX/iEDL
8StTLtMnIb4Fy4/5c8wBagtV+hKaHkBE0GTnu3gmnExFvfINdeMlgUXfzfYP4Fu6
6mrZ4HBlZFhnADNROr2vc9QGLSODa7cICy5LDHVDcPa9ncbstTcgWZf+6EKkJAzG
Rc6GBQkccU6E4mVzZrVA0JsziI0PtLykRw8vbGDvh4t+wKCHWI/5d7Fcox0rY2GF
ZducHoHzMfSPESdsOhHX+dscvAyjsajJ5POX1O6/xNNXG6RQ6KME8pCpJLEX5BT4
ROmmzH/88aLojhPxVRoqKhzXe2FbD4GZAFyZxsm9sGQpbz/k+lxktH/l9tYiHeoc
uh/T8hKz9JC7UoCNxR1hUd4zi8IL/1iEZwy2Yi+dKvcEIBOsEhlWdUKt/U1lpaiU
r/ZKnDLNRHL1QHDU6ocQscw6IcbeE6D23e3yPNmrKv1fkTBvqm2v7Skq+2GLALBh
+0k/lgyt+/Gr6bK2tygqF7gkAlWbt7sbijXadQsPQNTnbWLjbOPGTbBq0f+2R3LX
8aPXqVMVX3vEw8AnL4cIPytVf2GzphsnUj7JUfy04fpQ3zT3Ph8I75wgcMCiLMHb
mo7MYDwK3lwz0dzhR9B+esGGjPVRloh3qJIkQegnzd5Z0YPcWxqpfGFbeTFuaX1u
7D2IeDcLBDwO2ljHJ6NkYh35344S8EFvQlNZBO6uuSn/pJ0LC0sqEBvn97MAtjDs
eeghvbH4BWOxm/hpYPBeRnl2z2swrrpRl6KRDP/5YhuQCEINhTOBryERHFgALlO5
dyH5ZSChl2Nw88lxuabxMbyNDkxHhjbGs8EihkbyMuijNgBDwjm63nIYx3iAGEh0
u3YdBSsMllWh0V0A5Cqa+UVc+t8beTvMzCZ5xf8CX0/IeeZx1HuotxVWF/iCccvC
dTjBfIGNsaiZDUm6EqfWQ83HIepSK7hyzCiOcw8CcUklUgc01QXu1gE1LOeYm93b
PsiiKg9YJOaFJjlnCYYP4wH/pY+XXEzeO0ArsbEij3J4PdR8zH19WtYkKYvH89LY
q0J93gbZEskd+MQdc4DM3jCE4zR9Sm6laGXsR1plyWWxGtAVh9xBIZVDjGn9iH/J
ktd42hxyhROIn8MQmoiJy+DK0EcZvYcIeTNQeAjfuzWeffOmXnYTCP+I+J+YpLDg
mnn4snkSteAmt1JVLXdp+Ki5YhC/3rWLyl0Mq23MuJq45Uv73Zl17Gbe4F66gvGJ
gmeMYHNtWV+Ed+qOax9Kg4BAtNDrlxbPosUtvR1R9Sva1OsuaARN3WK3AbGs3n+D
ZZpxzNQrla4vcLudiTm7juMHxxTSxF6C4cMyUEIrMgA3ubaYHizegj/zO81woteY
KWa684E9k9tAI7TPUV7ngyZUd47/c+iszSRSGXqSIU5ELxPdhLfASWRyiyzzFWe5
oHrjnKSxfd7MSrfnVLlGG0T4VIJK50ShlhzOY/spY81e1wjxYo6LfHXkFiJxkO2M
2MTTBHHItBjf4c20gRpCSlmSnab0jvx8JlFw3a9Nw1q+zf16aDDKnb/QaB+1Dx7F
yd+NmnNa4YlJnwAy+DxGO9YRNSP7VkPOlw0XSWYUNLGH6oC4OksJXwuaTZQl4H6G
+/2Zydumte6/17MwLuR0XSsfTqGmcKMQCldHTpxrSBlPpscAqy7HFW8e+a3Z81em
/OxEeL43kzStGM83AiDJ/EeZDjWhhCSfIOSSxS+4TACA0P3IpbVTY4e2IoJlp3NC
3NZgZ+cqxaBIj0vN0oCBq9prQUKYm046Syo12//JRBc8HzcMVdOWr60aYL2iQWN8
BMzc5t2qrufqIEs+M5fmM4cYEEyVAYrNs78U8aAWpLJln9ihBiGc/8ViS/iuEJFq
XR7BcU+z3Wy3PFxDXu0xCTG/DAws5qSW3yUqk7FxhSsTaH44DKsCTi9EVyOnSL3b
sxb0AnvFzZzHkOkHBgutwts1xQ/IkhZAjz6gLSIB6GnNjDpkTn06w91GBW8RfL5V
zk5prhjkJE/CpB9KakEJeUVyjjXyK9JvO1zhidyc4FoIO+llZsLWJdSS/DIqG0xS
vyuJF1qWH7H7HRFZkMxUHNL6zMYnh+rbpjJdCaGJsmDHlV7Pb5m1lrlP4JeKV0jb
4N9n+i1RlXJbFWfYO4QC2zYn8IU+7Lmd/IE3XrZadJOeVTVhkOk8hR8CvOAxKxLi
wXQ/db1g94CkIeBrrjNqabpuoCZnf5DCS5ot9C4KXq0UdrdpnGWxRIRCqb3Z54j9
PPq38U/CTZ+b2FcrGQ+2RSgyhh/E5zWIYfqaxi9z8HsMBnYdG+X9NfBHswJWZNo4
9KCl+1/Qjmks32GxIn9N+XPBsdznRzBgot5PI//l24SHnMxFxvrkD6MCPi91lme7
0vk9lkr1YgZ9xvAJ0Tnmzbi1/2PgRxHrMNi1dbtGvLtagk+ntxON4HeFA9CmdAM2
PL5N0hQ88YmvTpPsbXRE6P2wCRVNCE0s5MiXHRiAtWjjZWIREiyN/NjeO+I+p+wE
fCK6K0ojXRbXNemWk5z4Fbn1o5TPyyF/Q2QKoNMPLvQuyh6fquf2LG0v/n+JF75q
UK34FrW4oaTY5ESWdrupK+t7/ZJKYA7dHrj1j2XkWo8XEzEzPW2e7bP9+A14mmdH
eJMCelr0WChfVUGI/eMMUIre+qI45O6M6+cK6iJhuTNDgDMSgWNPxeNW71QXxp3b
Sz7xWzTS1jME9fImIXr1n8L14jikUUPBPzWrNGq1rWwCB9T1wj66Rqvl+8j9RtsG
xOm1wEzEOvMCuKhV8eEI+voiA4ux10OtoXDiHB2IB//dOR6/qJeLupSovFhnCpzP
hCNR8zDkydMI+B+ii0nMtieBH/bxbRGrpIBi/VPqFSJfbBZbgBopTeYUKo51R8yH
bjguKSMkTX9SAsLqWSz2bdRiFZzhfcQXPAyA7L+JJswByNAIDd/h9X9tAQV9J/eW
wGixt6S6O3K4MYvOnLB3PouKjFsPgCvunLVcBo8cwkuQ4Pc6GR5SfgAu9MjjZ3I9
hcLivosp5p3tR88CRRq9s64R1xsnkW+Dwo5ol8jXvs/HZeSkMTXNUXoofd53Ub18
zuoeNcVx8TRhv6kkI2jpwjMJpbXzXCfC4jYuuzKvCc817IRwyiihsnlBkS/ZxKms
T4+Z0wfy4QqpadD1GPYhkyFKso8fuDds//j2YOSs7DYzN7soNBCX19PJ2UsWeKfj
agWK7e/b/Nz7d1RXq52OdCFNOoYHIC6xYF9cpBn+PiLYNK7Y7OfLQs8KqSuSgmUW
l5QkVF8WMfjXzWpTWcrpDzQtOW8gHovdnyAlixVnt1DyW9lFfXuAxtjPUsGF4hNn
aXQZK5vUMsd48n1POAehuNFbqh6VcqDTMnXU+DUEeYd6zjbxH82S5d4ilKR07Fwb
VefOAEJ/DJn0hAwUUXtPx/CY6TUa73bUqih073xhwSUMV6cWQDcwjoOTB2yBcZ2Y
LOHVy2cKwImS5kPAqhXU8TwDBwyZ9E6d2vLzQ1OZB7jpqV/qzQnGWR3UR0ieXlHJ
EFb23NCf3pjY8ch5N9HXZPbhoNHSas/PnlS3ZmVxm27P1AhYiNuPVcwMoQSzkIPY
EZLR41EWOBStUelMJgzNsTEXsrWBfRewGY4ryCs0uQOibVQKZopXdAectiz15yVu
FhoxKnfbGTVD/zvW3LQvLE+yqpVxeFl3zawpL1Ty77GJCvw6oqiHh2FmZKU5v/e7
2aYJimQverEegjcq9qrpyssZOgi8zxU3W9UjnmGP1Y/ptZ2ueKyU6dGYL5p7X0OY
Al4Bg8djhfWabE3w9OCUyXZ8oefcP4VoJV7xS840P672wGWw8SVcw+TcQ7JhJNEJ
UcbfKuvkrWaXhUGxsISIT6DbUEYf89lvH1BIx6f6bjrTx0a9YDpH/+bsMw5ZNbpY
KvDMblJ5qEEsOw+i6S9xsX/qKSPu3R7swYuzTAsRZpAX5rulUuP0JfWm+riFDu1a
Yse9+fCs0O/hejsJiEDZelrAWtvRdXbIBuLVQwgcR1SQKf22Zvo17iWceN5u+F4V
G1mbjxJEI5DuPmTAaGbp54oYinLh6KSqSw0LdyBLy25sUsVUBjuVzZ8DZEzqt4uv
4sPrF6ecXvBuZu3YHU+AuCKCl8649fdapZWS5g5iULF3jG+Wq45y7J7YlmXavFPR
SwewWFojP/9AK1XhvXTaq/Zaw+4AySYbpbSQSCUjmk4LkM5LNNmdXZeMYXGnm5MP
SDHd6/ezUcB2OBoa/TyLDKi18Vh+y76iZ8IgCIkP1Vvf3/8VsHiFSvrxOXB/T9BG
Y6Y7i0lXWy2PexsTTzRvcz99PZcEWHwiYXFEGezpKdc5b04wl0XDPbHbzrT7ymzE
Y0rrh9LPGl85Zu1D0PnmPbgCL2BNiUvlef04tbOUQUJcATrvAvedkUfiL3KAqlzG
S9F+AjLzBXOwP9ltsIE9+HzSDxGYvLT1/p7ZhwcD7lhqKS/kHAzRvmFbXv/CdcsC
GtgYLZhz1POlONLtZTXPVeFyYL6trs7iREGKqRknmdB1K2zxasfVKAY9FEkocSMH
jmnK0rc/lTYhzs+S20VSc2P91egKTMXmCoFtQrJqIa9K13iFlM3rb4ZTArvwsA/0
lPa6CNLOB/aerGSSjX5PoZGgnYYj02TOPrzJ8UwtVBGpFne+cb0tghLNI2JEwMT9
N+9Fru0EuvtyewVewTTZ3wtnFO9pn1SkOgPk3HT6Nx5acwtusMDN/Rc8lBI7Gqbi
RuTTmcBFMaX7TVL2lJMAx1Dvxzwxlw8s21/bfk7Mi2g8a/ge9lDkw/Ot2paTAOhO
9H42BQXiMQ1D24aN4/t/CRVTLLBxBCrOhLkqb627LPwr30WJZJNt6YIESK0j7vZ7
ySHoFN7wMsJHYzmJwM7/zxLW6Qat+jOMT4ku2cSZQVv2zeoOlDG2sI9+tYk+TnCU
veWGr7yViMzPk2TbpiBA7U2Gl62FIURoKEPPLpTgdknyZchFuBrlXaNWenrKvZgj
7ATtOOpT2VGrX2sedAYvqZ+FP+UswfsC4gRcifySnre3lJ5MDWc3g4NbqU7ODS7N
tP1Qv4o9KZlLOIQULZRJ1mOv+gSAc1xN6X4qbQ0Xf88EzKCtTImi/YJRSEpW6btX
aS9L3ypNGiy+YtILnoOmgqoibdOHNI0kwLMrRYI4puAOQAfTLjktrXxIDCtqO5BM
NIVc/8nT6ai/k36mAtXrw5Uw8t8RVp02+OZmWUdBYlIKRSCfpOEaRDBN4FfzOPxZ
M12bzSuwV3paSRY0bj3YnL9pFMAOlrUstalaxI5aobnKgpfPlnSpfVLLLiisyWBj
Baz1dqgFY/d0Sw2F4ttA9npb85s7m2F5VJL7p3MxtdUwxJlEbJIA+yMO2c998Kx3
o2PIkYMRKH8hD0V6/EN/BUmBFVczSeTDyTMpLNyo5JGJDpFaC3Rw/9Sp+C67xvrr
GOjzZLJasf4cgSNk2GoVsfXBIyfbKC6t5JXtZzAEX+wMuF7c8IbqokxlY2AdmD/L
w1P6tvH5ITjL8TD+dXtnijBNebVX1BUPLx2YyySJ7hW2K2V1W34CreMnP89oT5Jl
bkZJvck+yjia4x+S5fB9n1fn6PP2iqqVvcO7dn454J60Dth7wMWuuH97iSMF2vRo
6w46ataOt2IYnYMJSHic6QYT50hFYu3T/wRTyQSP0UR1G9TGh8uJZ4LwrXZY1Wzo
qowUZ5RtUQtBm47FpNinnawJZbL3OywWlMf9eE7TGeknjErIUi9mkWgupONJkv4B
5H/DgM6uh6b5ByBBnaYJ/Ge5xu66TpDxSmy3bEXkbzJn9aGzVsk8uQlvZhAH5tKE
E/jQpwgbyYiC+eC4AUjf3foNbEMNczvUYG2qxNrgjng5fOUTwsHfF+wVXZw2XG0k
ENuTdaYcI0QucqGPXvJDlX2KgBKvxg8I09k/yD174+tdeQgaFe21mZc8Wv0ZMQUU
rQ/4GEBHjtUbFn+Kl0Nrik0A1NOL+TunA67bcdltPZxQzb1fPuOqwC+bJpuD7XJn
Z8QO/DwE6wSgir+3nlNfASaVeP4spiOcrvXXA8CSc3k+iw8IHjef7thBkSzdldjk
6W8DxHPoRXbAxR4xJ2kHB6u5NKCZXfTThfv80DvA30HmeIHcu+uAWCqWfeqUwNiY
wV4D+W61Z4/RTimcWRTn+66M7iKCmpvufNowxOw0OZnT8riCCx5LKcfkrgdhAEYh
tANCUXbSoAOFPvHsqFN8leErbf59VzwS/WDMxevIlb9YPdJfCOGUJOjlxf7CrwtG
W2L9Scu47k7BZs62+csrleZYsXRjjZTbubvkoQUy5l/CtdrlaLJIcZxra2o+j4hp
EyIJ0gy0mzNXRVPoL3/P6vVNJd2FOhpFvbWtV7Q+JhRMfYvXqQzlgCNrqrLJ3pEt
/KY/Ny3ztrZLTLb4QE2vYVxRP5TxNfPMhOyqZ9oijvC+5c6vff8U8GpeMIe9PF/D
RrMUcUUyY5aEcws54HEy2CMsrWyXU9TX+NHRNdW0Pdoj7+srtC+WQT1E8vgjCPCd
UFD/jA1l3MIHNlDrF/TxQCS3VMFog4RY8O+Om7+hJQT//C2d8ltT5PR7+Zf4Ida/
ubxsqQKkTacOyauvB8IKDURX//ybrKclKt10rvkWdQtO5Bb4sCagMlnJcJYrRu64
WyWq/Hva1PEceC0b8gDZKb7PrNty2eCYdP8sPIZXCL93C2tvM8X/pdUUc+tHPLMA
mE8TQ70HmRMN9G4N7q6Sy117/ii+88jmA59mKuXWXHfcfkyyUQ3Pp3Qf1ow9J51z
InHBaafiA2FuIMeSoPX5VTPup8t/LhNgi039IOtOHAS6LcC9HiAvKBK5kyPBhVJH
OjvDLIZTPXUYiOY4riNGLkP17aRJnC4vA8mnDaDMBulN+1/Ue+2BEyRkOkt6gFaS
2ssKanlVh4AwkAm3QOCaw/yRoht01UYIA3CRQ6wmMhyOfCmUjED00Me6VW1Hhs77
wP6/0XbS+JfnAbp/3/00cHpkc6OPhpsu7cYGNwfEuylfuUX7eWOr8AsmUdJQoPzT
kYnmQV4++GLXbww2KTET9okz+2wivoTpchf0NcLaURdMWwy/xnSleKVxysLWIM/t
xqmSMLiXe1mt64J2xMNphm8BgYArLKjmKGghnLasHyuMkAtEOEalYisyxNzD2/DX
qh5liT2jJpGEBFk5S71ho6FFrucFZnRxyl6lX71PIlGCYsly7ycMUyd/ndOUHKgx
0WjVOH48Ei/Ts5ok4XkQZ4ysKglBXIVf5JI8ffUtXzc72+c5298adJkjF0miV/Oh
BJapwM0/vdzbcaFzdFTJ1jEIhcLA5io536owaS2k7MFkP8FS8DuEHP3J0ThFTCbI
nbXKaX7ta9YohssAwD+KeeRX/FtVdf2dqSvJ2dCXiTVeNppQwOI2mprBCVMMuOQP
uPgwgQcaIc3mLYE2OqLxkvvGJpnSsWp8YVBVivSBrwMyJdtLxyPSpnJZfFh84/1E
kijs1AWI+3/dsWvbeMLa7GqGx0xSrRXWAf64oT8hIlll+P+JnstjWglzQBpNQ9Ij
CB52qloMwz+MFn49gFKNhfxNouwoRjHlKl3FZHpNxuuYjYrXAJbHUfd+oh/QDAm9
GQaZV8UteY3yq5SRP8noEbkc+hPyY6Htv+jPPU21sr2iWMOM/q3JrfaueId59vOS
oOf1SrBLfYp/qwoiEAPHEj9KCfHgsz9cVjxr8BV4zgCXuWqB6EFD5qPqy7b0WWPX
6MDuTsk7fwFesbInm2YdO23oAM0fO8aSM8vMAH7tSLS/b2DGTPjjyPwQYjomVV8t
j+jVFwpY7oDGWtwCdjx1bbWhGq7MeSzH5JegWm4/bP1Us72YYiRzI13UKuk2/PpW
HLOwbTBCYI8gDKfu6CIQLQu+SnwshmIJQaciqApxuoV4SJ9HWgJfBan9Io0rdNQo
aLe7Vc/WUpG0+MP1QEiAULYrKYctwrRJtFgEto+5rTIuS2mUWfJbmyOfPj04F+Un
4MjAxG/5xSzfhyT66mOIEA3LsWP7CvJU8BW/bjYkhZXue7QQg7tenhpsOvPdSBrQ
3uqDYMoNKDDnBREHnM9gHETi7gYc3IjubYHDs9lISC0lh5uBsUhJ6YHJxNXAVV2A
PQjZZcoMXpcb4lMlLRjj34YASPC9CiYeVavCl6m+GwnezOzKvgZggsZIsgD6V5Qi
zllBVMPXkhpiHZ3GKXrbgFa/hTJUpCJWUm+WG+/L3pdRzdzwNSyzB+e4GjQYjOuP
gWqQE1lJpwNn+FTG84WkTbAimUbEc11knVhjdnhdgCaxnIDpXYCXwmWrbU89r/xC
C1sf0DZlUp82p0Er8CwknQE8QVVJUnSKk5Xv+DXrwIo86LKL3mABTKKoAbtGTtUd
xD4wMZN3ewAliGPVl0MeSW+Laxu3B4aIcCLgCPjvA2UlghnkwUk63bdYJNm9bUd3
eQSaEMyxpH+5AcVIJH7UdEvYvnsrTnkCsxA8ZJnjoA+9oyGWYOtHIO4GQzEUFUSs
VTPmbPYKt/zaQfZtmBb674dBboiXirZ9gU4WOOOSdQ7BYIdRPTextRLZ3EUkDYsg
hn40LqT/2IIQpj/LUbW0QjxxnIaDdugA9kERTRiuziaWfXimzYQRk0cObsbEVU2C
phoj4Va5s+LteJpMzMX+20m6ZRxpJvSNpfkjotBXtY5uVmzRb+mDQQB5t1McCb+u
AD6zYZQcCMURKhTZCss87kE5iAx75gdvSsYvZdtF8Vs3PyG+MZhUGexXVi6qn9Rg
TNmApXrw+uF7B4Kiu+HE3DjXZ8OgnVPUFC1IT8V3jMDvlQNJwteJlOBWrxAxZDRj
gueH0Wne3m+Ihf3dxy6HPzzAb640GvPGPuYgzDR8F2aWHQczLDoTt5AFB1Kl4umJ
UAKj7yefvfHmg46kX+K6VGRZ3XyhTHo7iqU2zgw62OzDihNbUoL/+GXbPQveYjyx
q1hpsENGel4/h1XtbP9hXoPYCy5HqyCs7d5TsaMlhiwmUBdZL5sQZYxoo/lAX+uF
fS9NDf5V+lKV4heuZwGn38vMvFuX9hWOzAliVZ1Fbs09NaiYR7Xe1Orma0O7N9lb
K4LiFir4zNmK8HZ0YRghNv9Kc9H+ei8nfeuoF8VGgHWJAYJdZIupc3yNsjiSb6Lt
Y281iPB4c9mPjLtHKWmXnK3miF3X2T4f3sjDVBdn6aDf0/4//gmNc9rOj4YpMuVi
k/4QepLptNpcY/NsCaRG4ATBydVN+04abpghejF3Az4Kpu5l2Add50PVQrvyeFTX
poMknh16R53XoJLFa5IkG/CBaL549W/7oIy4OQ6OwC3vkARTsgtJzWaNMePIPjbX
Wmy69lRMiNpxiawosQFfFozTSOwkadHmL6ccpwwkz9ogk1lUBZ2gy+D8AhbF5C5c
wx2pwg7q8IARuHiJ/R/xJv24AB95GuZgSdcVOgF6AAKgFJcFUJdLfAvIzy37Fc6+
pU9/KG6zFQJTbWmi02nLirNvoF0OsiDE1cEELtaZ5QsDV9PGsxeu/6pU/QQTR7mo
nn9Lb0b7+zDIp58dPCTdthJykeHrh7DjcmRiZC2ZQcxz2U7E/1ul/DizUaGZsXQZ
yYi4WjohGpP35b+wKKjsG7br2sEim7uCN7/upxUg6oqMWTsTRefHj3MyQJBv4Dke
Bg0r2czSIyDuJkoq5nO8OfLtFCEj44/mS/C0NiZ+DWq2xz/B8y4vzaHkKlrUlsVr
0xedDbWRiZw5YmQFk3D8wHebLn2dE3JOZTxh9buCZRoodUsOS4tqIYN/w8NZ+G2v
v2WPM1H13oCQeoln+w5XGLVJrCAN1EaU2i6H6DLnJg+smup13fSfBeH6iQmJD3No
BVAbokUb6mZD1SYaTnDFbTSBi8rvlkj4k1n0FEy6brgjpN32aIgFxIWxZGVp1yVA
LFbKkMpOUiItZyYEh9mGSlzbskNyRNHjKShGrdaBMU9Ot1TiDaT3yVXNzYqAspm5
Jptr8ycHV0bZ/kFVcVTA0XNeTAnIecpP1jpPjjYp5kCnpMofsq6O0OsUJn0d+TTf
XvG2nTi7WsIw0ps3+p6S67nslw8coL4Vzbw8vIvAsSL/IdK2mywD+st8U0Mpq83h
5PqukkkdKctWbjD8qLvCIEn+SXY7SGr1S2AFduPvfhOngGPZi2Llhosryounc0o3
P17Tk7N3Pnl55CSjWGuIaBcfiL4nMrmkqXJqwS9O3ZJz9nCWjYtIJvpPv4KYKFJV
f4Hiy0QnD84Bd+nIMm/4MoqduP45FoPrz2iK/Ho609PVA8q0KG65qNOKDphyRgcX
D/yi5T+jPuiQblEzfDcKcIdXqKqujUwCQsoXYiPaOpRuxHVYpf83WQJTkLcoSKsy
4oGmubHIB38OXe6RAyYzUatfFNmiVQ8QpvIOVReYWRZnXby9cFBzEnnNzHEpvG+/
hK5UDBQOxe4CYXxzXb9i6EFPQ1rF+qZu5lrtSuGIYJhyH7GIVPtWk11gZWyfVOqS
GrefNv3+q8rlQDzXZ8rZNWkL7SyIQoSFkjGSjG9G1CGm8+WyWKpLYU4VUSSHqmyu
iaTS+C8FLBYBcBKthg91Puz8/k7ZUYgDfh+MBlSC1rzxDSb0VX5a1OUKCZlWWd5r
//WnHHCyG22r5soQmmOq6MGyB5/9wg4epAVwMtyqSmQ9voBmj9V9sNgbVNorZv0j
kk3A00m9Q3QaRIdQFywXb+2qn8fTvHwqGMGhGHtmjxlvdYMzhZNSRkf5EFeqr486
3T86FlgiarhjZVkWk2mgXQrLgfjNYBNxTuGlyq4VS18DsnnVeOy1J77C2622DtwR
PWnXzbpfibgwiw11jQjwsQ73oYzgBDystfqDA3IgcluhxxrFX4PYwGK2mZnFSQ+m
4QZQQHw+u5qlilBWqWa+szRx8ZOmuw5soyBcRWFsjymOSo+ohsNo8V87E1lu5HrM
wexVqw8h1vFTFm3tpx01oAdGj6kcrD7xJdViNGE20dHRL3kS+XS1Us1dzpCs+mTr
t7daVQUHKMgDOY/afQIkyxQe1NlnPja+DGPxM4W56P7PF8L+3pPerAV9rN36WRNZ
Cval380g31+w2jVBto7Irh7iihFm6G0vRkG+mpwbwEpofyCErb7q0oOORYdvXWfR
40Be7ViwHS7TCuvBR9aS2/yA+rxXWZ390VjKF+RAQsM9Yn5kvLx+URfiRv6nzTM6
L4WrEgjIGVcCKofTfPNJ62KAJyVUJySARoWrnRyJjA2Uqa1KQDYF5c+l01gAi8Ot
cRwgW2+7+V22zP+CzJ5j637Hq2n0QD0qCkcYi7HgkHzwHnHEwhM3RS/DeqPxxPOT
ijnR4JMKpoY9GfzKN24EjMWfbmiaMXbpXcy1dRwazrZNvV2TXxOFvXazd7PgvolC
FHa+RDombxvjyDMJB2M2IW/g6mPQW+x07HQE4VQYhnMNA9PkmhzGPMYlR0la/COd
GTpDszbwZNpLd19t1+ec5l7VUj592IjfVNeF36YGU+nTNeNXrzny3Xkacy9KX9dZ
1PMg2sMOMMBBJolTvNYiAkAjo4xLmsPGweh0xGUpD59LFYsSKwRo7Lv8/ziOyZPS
pt3uGhj6uEjGpYhwUwGqTHwlKi43naB7myBZbn6TNBckPA8qOO3CIhf9Jlq6QFfz
Qm/xSALkjgMQtjTHiD8ryqHp+8cPdyblxZ//gxV679C7cRDxivrN0421LdYvTVVw
Y2P3uBiJVvk9M9oJFdQ0Lk97xyUx+AGMxc9m2AYaeNqF1D2N8iAqKYEiaqfuDVKJ
MTvWYapScbtiXfViHzy92mjzUzJjFTZ0dZXN7iS0B5vUapx+ny6LB0AJaUtYUiny
CY0TwrHHpgXmefi1gWjXJAqSHNl8/Dvhbuz0zeGIwrJ27FPgkH7V1ixP7UUcWu5a
ooZXv0YMXmJLTvGWxZKxJ7ldA2qlBlK0PpnMvyOKYdXFDls5zyScNcY749zVVb/X
2ri6/GOgmnPc4R4JVeEgaTkpHgh9uQ73+8RYY2G+K4EHkFDtpzPpw0dvY8pkkoTh
8DC8TGZhbXWdy1tjtbZ7EvGj2Wg0c9zB1GuTgAHJhyx1y+GyDQXXJxxV9rSjlx26
YVDDNSenUjZlXp0YiXtFtWfFJD8rxmD6Jcl53Mu6jcW34dp2D884F7XmQlsJVhS8
NLIlZDYqlPA4PG218q7IxyFiORa8XNbWK8C61X+xF+U2+eXZAFxxeWRcHfh9kKik
94DtcQ/Z7gMxeB6HAJE4ELL3e5H9xRvi/DmVglLUGbG1JgADVSHGuz+SNtK8a+CP
jGA/i8iiuCgP/1N7X454RUTIm5lWfl3w/X85vKtE6cBxZ6mOT06pm+5m2F9xarvi
XUrTjGgXGWzyfu+6ceZIb4EJ5jTxmlBc/0gq/aIwlXuwD+iB+CPn+zTbflDzb8Fu
ri+XXqIPA1NOWEcEEemQmBkeW4WMtVfCD8OQtJGGJW28JqXQUY73BJhsQzis9tG7
baULzdqECliW8RTuEqrfMph3fNQKzJTMlttnBsmmeBNRbBuet55yttrUjIp/iklg
pzhSf4NKYe7AgpV2UrJnKxnbJddxUYGwAZdh9IQse5wBEQdBtlN+kidYyseTeExv
LqSMpPvGFf0kRSY8lC+m6oWNyIg61HwZVJC5vTVYJ4LHcnROUniDJYCLz7XOQRT1
etDNC0ZmvgBajSG/x8xKQ9YT2+aNkDWSKesvGmbSmSzvRgr2JCK+OrKJTrXWkBHX
/UFFjKKUsF1807YBYYEiFdO/dCN082Z09nBJrgGHaCRkp8kLOg5XyMbCvFOuXlBr
dGqT8e/ZXkAGgUtHjnY1lmL/d712v2vNbXPIOUQF1T+DXMBqV5CpXFIanDerUhnP
zL8mO5Elp/zS6xBUSFBKF8qmBo/KOFZOIfT2ZAWF7eYum7VDk1oPDlLL9J+PD4Nm
xvmoOnG38hgGpcVxFsFTrdq3HkSRqk1VH6J+arfqIW2gcaR2ACFW//riApzD+LwO
drl8nvTXG9SJg/+JjLs2rsPsSp0w+/OzdyhkyR+QMtTXyKa7zVSB5LX0OVEjZVs3
PhhT3W3AHpqLO+mbQjt1tTCP/vOdkIA2D/Bg09wGNX1CYHYy2ApByfdlHk4ROKLS
s0XVor8nRHmpXrL84/AOuNRd+qCpEQIWKiJCcN/8PT0cgXlm20+gpsBvjZW4Vsci
BdgJVEraL9wvOBSzOvnr9GbxJVHqTrOVN8OJ0CmMvI1Yg4TjsWcnximkfYLWe3fY
RuQsgOIIqbPChjCXq51QJmbEZyjhTHQJ5v39VFjtLRLP0I7DQDUhX30y0GfPFpWx
fiM/+XpX62TbVudiBoB59BwJKNmHW89ryT+gAI0rkHMIeS24PzK2WZcXFFcgXCzr
/m2blcLH8vs+VADCSwzZax8wDxuqinzwCLCTdhQxd5puo+xMd4PZF+SjIk3npOmL
t0yu5gsFv7mW5yAXyBUZYEUzwKJquUjDm82tSDM4tH4Ec9rbYfzKwnorFgEZcmgr
+O0ELN68GmIIhoYw06pgPlb5klQ3rp5mZBT6oQJqzbwKsL8RPbuRDQYvW/Kmfa50
qlEEsPb6eRyqR2JGMCZ/I65NCxOEgpmvKRO8lIvp7+Z0UripnJOQKUlpFjctaE4n
b5hjAYG+vfpPYddUOOtV1Xz0Z0IslIBoshlivzexqlSN8XAYHXqRBBHVw83OvyIP
KGSN5apyrHpo/hakAtWW8SYuv8t54ZVWGnsjqNmX6kb9rDnyJpLxXwQKLulRVmIa
x1q65RT0vs0rTz9aEpxUHiZS2kgc8jUS+3Yy8WRKb8zCipR3O2T9O6CoL8mELThF
mP7Zp5+QK+Zkn26s1/7PVsjTkPXyrEA31PmiBzvvn03gbCiuaKT6z4DOhfIL6Zip
HJAYCiSXX76UG7hTKNv86x2F3XRyAJK/SN2WedyDZ2IsqsjiRluhuEKytthPY0hr
NgJT/DFBx7PN4+Jx4XTqnEBWIwZva/dpX1rLP0KC/fnqmC9kXF/DZDYZafV28uFX
th67JTXrskJ+R5SntdmVhAp6v6Tkc/MP1Of4ZTqmwtl0/kqIMWWAVIweJUU1ktfH
VDDoE7S3i/btQSu8Eb/ks/HVUBjWCSXC9g0wSwgfqTHehZ0dQAwMZdP0UZZTKyIB
b0Dr2VbX7uB5f4jgSPN8tJKpc89v9tK1UdV1AB6wrwo28jN1GJKEVjqGd6bwmzcb
LQBSIn2G7axZOl6GGWDgmOhd8RZR5zs8rAB5qVoHARe2rfRxhKB/7Ca5oWiV/lR9
CEl43r4IpoqYxZpsD8LwKyws4xTecitgGcXYQ45G3CM=
//pragma protect end_data_block
//pragma protect digest_block
lntgCns5EubxyFP2I6QB/KyXd0o=
//pragma protect end_digest_block
//pragma protect end_protected
