// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
llrVxcFit1XVxUEYx708g3Fttf91i5oYtPzrlNjH0nrFWegtTFUhqFRHTwWs
VAkQt/6dJZrHAdkoiZiD4+KgHMWkTzzT6ROZiyu5nZRsGEB4Czky1SNpJ+cv
yJWL0JiP3yWhI0AIHxIB9r2WrK9O451hqTcjMD+fDrRkx3Q9d/eE4UvCYe5C
6cSenCKdHofNMB1PMcNx+aINzNmOVP50lV1LALHDwYd0FdGlRhIe8NdITFbC
duqk5/Z5HL0ecqykdx9tmo7+JnJizGBZvuOGLxXBgZ4iZiGGLttxi9Hh+iiS
MdwX5o4a3YtMATYDCk2sOJadl+GcCGMUHgrkxJ6kJg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
oGc5nL6H0sUt+MqpN3obUXuYW7h9kKroSeMt/lKKQfHGakJLP63v/WfNqMje
0NzqUK8YxBO5fj1+aDoz8tgZ2hWs1ycUT4sjO0WYk4bfTcgGkEmQINJtQNRH
7uD4HNuG4jJw2JIYHiSHV93pqhloMUD5shhPX6ndFNCybE7ataEl5W0so1+e
ZjHHv1kT7+GNFziSalh4kg07VzDcSVqxjCOVLJg/XaDOHC+mrBNV7adt03kE
VqplfCl4O9YAfbV3k9GDM2611V4s7i7oTVU3EXEJEJKe9Viu4EQhr0PYy9+N
oKyvdhmJDeOMm9D2LMXDsKtrI1ugeNcs7f10qVXp+Q==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WADwYcV80V8tH2rqcQoTChzy0Oif9KhQfaM3PjCfRlSCOy3ImX0O+a7y1z0x
n5Pi90imijrHDtQikgIxdsXeKv11yeHFjs1zHIOg6ENeSJccq7JRc6IdA6LP
7CF6nRQa/H80IYrfaih/m+J8OEa5IZ6dpY4/mIHcFCAGvImHwC7SBr9MRdOV
pWWqm8/EDiMdVmLeXtGa6TpRP9wPfsbGvCnOv/5u7lQReuThgnYSHCYuNjtB
QXhPFVkVAldbrGr6AXZXWL2vtlJJKVarK+cPjjrh4cmwye319UMjrdnb4YHl
fFo/TbYbhiZ/XZDIRm/s9yWgDZQCvNkE4dVwNsfAww==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
SFXSzoPMG3C7RnGCLlvJFnx69ZPfV134P7o1tTK72m0kJtxoZ6Tpksjo1mIp
2OqbSTQms/N7Og+P9QB2WuyFodHAYn119pmMOPyE75I+w3k8PSJRVe5j7c79
EkYNG/Gq4RE6eHEKuHZA7yjr4UEIRNXT1u/XIJQPJHNxwDI+wkU=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Kll5Rxw3+cjY7z2eKolLxfjXmURk6CmQ+SNpSD3zJcvxZv1JMf0KzyXOKy6q
pxLznF4lrdrB8fRcxk6zFwpGuvAjBzqnN7vIrlKEWbFUHwDV4YuZvlpGE+ZD
QLI30ngKwIhRtSsfgcBY8yLN2/RTt5KTN/W/TfXWIJ9gKV2fmjLrZnbTtWW2
qJ0ln56xbspIQSPeSeOmL/On0ObGOXmzN3/qVMXiUEg2X7bvd6+juGSVaoiB
CU1egWL7ya+0/c82lT0xNNtaNpC10bk2Hg6BNQZAlRbN7Nh0gPu+X1z098ec
fmQZXQIqcgY4OQg0mEEVCN1wi3Mmq2OYeWejHIfE+oXW/dFiJRvl4TvWzWPv
RmJeTWQSlFlwsNozfZA7P4roL3XqLNhZkBSs+G+q1a0s+Yj5h1/wS1jpnR+C
pNE4GDWX/Ti063PBPFoQV8hQrdmGGxmVJiLvwlOl11yTna/DWveIRE+mB/HW
rOF9kmBDlwM5k9UAFp047mE7yd1Pd9tu


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
RRmSZSKhPRZeCemxL12bAN+nDWxcWrHq+dggD/73VIWrk5VpVkVvpUN7CxBn
B1iQcdxFDMK9zNswcVyBl+onrCoJfSpbZPD1hMOwSTsiqxvU3p+FqqSd5kHk
js+rs0XRZqLoJ8FoZUzhd9KUqoZL+qUZPJF7b7mh3rQpoi3PTcE=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
cyIo4j/90v54f71VOtrtQVoMtEG3bR0ilaUSLLoFxrkWKT+R7R3FXCkmzWzx
7rclpL0F5/GqVGnXySCiWNHGTCsQOmw39doAvQ2UFOPh3oyrgGhloIwoxFQo
DHtySUE5p2kOnZdMZqSxar+AyDtqecEQGO1dLndeMa7e6N2w4Pc=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 13184)
`pragma protect data_block
5DB1GfEvVTHiSMXFuGJEdM+fvsC9jPNVRZhioJHZTfYScd3oE0XOXoU/vyG9
mFnyjaIbASQiTDk/CZiOSmbVYVnNKPcMSa42NqJ2YlqISE8u5cs6tT9mputt
RkL0e9TMX0s2J+m0romJkp9wx4hBLvbk2hYgsebN6zxUQ1qfodyuaTcK/7QM
r7XNNs7TsMFJPpp+TuSDjjd87s/GTKe5ehpbDtgq6JuJJS+AAPre9QeefqAu
595gCUoVEazxWPCgTyL63xZ5cNvEbwmX3CnHGS83RR8A60knhvpQJknF1wFp
oAruaEzI8H0RN+/4DTss3ZOT+EmM+EUx0E7Umj43KZP5fOaHby7o3HH/3lMR
2orDgcda2+0keyaR7muzT5y9fzem76cbyxYGzfD/8cbhJjL5SLlT61vdArBB
xygdL1uHktCMLgdz86QTXghCX68SBJ+OqY6CFGOcCYMw+mtqqaG1Z7dXGAcB
5oEEbgokzjeKDIcUMgkRaDES6aLdLOtyA1mbG54s0NCVn4CH5vD+GXd3HcZu
ljeaKJRyxr2XsZMosH5cNUocpJ93p2NvV80Z3gqMHMXREGY1aAS5bk/goY+3
wE4jeuoOM/JJKhfEqHZdzoSHZg0zHmjCqlF3HlKGy0hnLSr9N3pKtilPzWaI
JeNh+K47NjOtew2GdxtBv1VLeR9yRPzH2Plh/bezsdP7NkkkWTYJ49KJAGOc
cFxyP0v6N1Ln9GTjlZk+bUDt2uqNmXIVfyRw/9kZ2W0Df5X1qXf26nwqU/Ao
PVIwv4NTV4Kf7bRkvb7wAMm4jTMKvdm7CSv4dmw/6rTXy5IhttFhGa8j6wzT
KbC1IOthWQzZLSegGC7Bmsmia23bKJCOHYCvhBX+/ccKPtvDEqmWbqfTd8b2
AhRNOBHqb7D/IxnjDNs0NhZ7SKEj734lBUWiOyRUMu+gmxEGu1iU7fr9UDQr
H6bRnHopnuW80Fam9actxdp4yhcpY8W7QNW6k071ukP01ECmED5izl8KrDWR
4ah7ZtbSOrGGI9Ah1EemRH9OvVwCvRCpkEhS4Z6ceZzcFiBQJKZ+77VFQWqN
CygD4urUPIeVj2oUQUw42vPbWYH0ltm7Cd38wesVIjCFSTskMtpvSNg5KYJl
wZF6ruUpMx9zDOFdXZ3ZCijk2DiPIqagCJ8k2GgkO2WcCBbZHCP+trrL5Ljs
fWWCBJUQMTSoveMyZmoiDzDSVCilDT+7JRg49Iw/LXSbV9KT60iSwADA72/7
ExYSi1+kIVWsw4a1Wth6gpU7/QVgDykMmnpUvNf57pWsxfOAo8Oh7k9bAo52
Mc4JrRB43Z/bMRGKdgPTiUFcyJUKIcq7QwfUfyFqVa1NhzBAf1o5UxmieE2Z
qkR/7ra8AYYE5LUGNrpdUe1Qns3j6aq+xzPo+rUjX4TU4M/1T5PVhVNqVHRG
LFz9F9dH5WWO1k7psNh6ElvqSEkA7qI3ZoGk+IERLi48Sm8yqL9SYsWZnWI7
y5jphiCgRAdP+11+nlp0PgNwfVcWpO/T3ZCRXT9+Lp2/zI4r751dOR6YtPSx
zjLLUNzm3dBIbR3xT91gjMkauqKmDGzfRqYETlTdnQJuzqNg09UYQLMQ365Q
Ii504GAMiAZ9vNkWYXZDAo1kx1NWpWTVYENetAwEvO7OoUIp2DdmpQhpnw7a
ncXmCGvjpapGYfha2MwCJhc1BzRN5udHTSZVeazu5O5lIVHnOQzctO2QXKoB
nBTPObHI903eFOd1T54Syz9E1UN4MOCBT/mCWBPl/vskvyA1GtnWU52aFMbc
uinA0ppddotyurJ3BiDTl2rnO6v4EDcAbVhruArm8K3+UGXU98o4JF1sPTmZ
Iy/cuJVmI33YC04aIv/shr/77NYC9UjgMZs3CZ2j+P43t/We9kNrNeoT36+P
lBtsVEZ1FeNzlPIb9c7b1dggI5cFC5C9Zd/xBKVQpui8/DfueAm3yleDiIpM
79JzUaLOtvgHBn9uOrNQzrXQ4tFbuZwP0fYMlARGW/H7ej8YHrtJFr8W+Xn8
9zfobjxnlU/01Zu94uXwwiCG3jmZt3olVz5sVIfnAednKB51UEp7ncqP+5Iy
KTVs64IEa3B1VIA75bK0Y6qMtQoebb6jj1dXzG3O8kMwO+//QT73W3M9/QW3
NulaZrM2xhZksSAuBlGE7uoUxE7qtpCRl5w3GSf6HmZvKLL1raahotcskpv3
5xncbHcrDUOcfMgEBr41eaRpIBrGNUAwzLMYHccfSKtIYfTDrMibDF+Pwovu
wTKDbDWHWWDac1xKktMnxVRYOEE7ZwrKhfIFdXllTRBQsvAHFPzu0go8llkE
OYnplHNEf9qvioxOirk+8EOnhM9JBK1DzUMqGyaj0ClhqieIQEqI/wGpZlfN
vLwM0owipSbF3aRqm+RC98OJAa6gcumxQrMQHQkWskSO2NhhN6lkJG9lebCK
bchv2v6sLwDQ0rLBwVB4zMJoN3G+P5efRl6oDkMPZ8bZoMWgCkY7jZXYNxy/
x4Z4Mwt9TpU9crDQeeGOmahnNw6EJCQanE5ynCtB1OxG2QUCw/qxgM76EJRP
cxn0nUprdO8gZKIpMKIv2C7P7KWR1SEjewtyXr90+UZasoW0vkF5qwh/kbxV
99ZHjIfXOTBZicJPuZOp5NR13kHl8o2W7TTO6ajh5kkkyQs6pA3rwQvCTbct
8IRQSkmk7Cvx/eO3DgCng+8BN0kbcMClo6J4bFm3TxVJPs1tTfq/D3B1QkWk
NQlQE7j+sqDjmt7cPA91I102Nf4p7x2Y/EkOgjSq+SeXVcGf5gwlT3cswdej
bceM70L6aQ8BP7ihmdbv/xPHlZYCVh24qWY59KWQ5+LwAsB3ng7+HwujfJgZ
IHOeaOJkzePRwTWHnVQxKW8PQWN6KY2oQgPaa34MfpxmpJeeWYL/SWemaNut
2Yu/gH1KTR5fCkZxcuqUPvTPGj0udXkDO8Ahj6ZYiigpJePI4SM9EkspU7NP
ihWLBfCml64ClSdeuVp2ovle924pSjNQAveyldRjkYoI5HVhirLGLeL3huQe
WQVYeHBJd+G/4WH9U6/dX+7kLwx0z06xviRtU6Q8c89y84wFCWxjbOMRYrbJ
16b3oAIjrTH6n8K/a97bq3Gf+HtGLBRggA09nH0JstQxr+tmYJ2xqnmkMoBk
j/Tr4ew/QxpdM1IuiOHtLdcsBuqiogUSt2LD4bbRgY9QHKChEcCwqDtZqTCy
aa8kATcjiqcbhPhy2GYIXcpLvM0Qe16m8/wjb9yLdZPwQeR63XC2R9DNkgxE
NQnmHzE0e03z2CVdJ1kDDAdnWGa2qtImgZhSeLDR+zwNEtw4P8t6aZhFHB+u
k6Rbx3ZcSWqAZqRyU/whhcJTe0/C5qQbIVBjfAY97xac4oaY0DO/2R+z+AS+
oXnKjCU0osTM4zkBgtFHSm7hPEQkJoLMijSBG8jVfEc+K84WRqW6sR975IEZ
aKbTBWup2TmPhoHx86afyYxcCPACRLUiSbi+tmiyeWsyrf4QkzGV3x5wUsxp
fp235VYydYuhPOD/gnoQX+xAbiek2mBTielplhg7KPZbK9PIp88gAa2+lL1R
4m7bUgV2zsojxUgQKZo8WpQq/QXfV9TnZtEOAQeYEWS272Tqq3QEvn2s0y1y
E0B0qpKDbBb7/mDMkeImXL9/ZHTnyjXh/BCedIBNuQWRTjs/3HWMRBXyS7dh
0p7YI1FqVvJBYdQJLBjL5dVi/jPme2qIi5Mbg0RC6FlgrWKnQN4gyFeJmIta
s5r8ZcTSsOMS9X7oKfKpLuSG9w2Lt5zTe9mE5s6roSg/GgSfgWdEyc4Nkbjo
2B4zvEqUopNikoiY6Kc86F3/+DBMtppXSR7E+4VI5B/G3CD7HmMm0DSvBPY9
CaForBPvw2n2T9WPiLejKbY5uJb9SE64JwTSDd8e9i4QVpPECIu99Dt+3+un
c72vg72qXKRbKuQTEXqTDIzW106d7/UuHjTxJf0vQIEKFAhpXWHMJD7YvrCD
A3mvF1TrCGhpyHkXE5+P2FkicHvyuJaHR3KYURHst26wqNkXhb6ofn03qX1m
eVhjLOisE+8cqR6aQjMTbYhJWfBHBEASYynd6WYT9PkufZljs2+n8u1fdu1K
truc2bZXW5rOLz2R+WxAhl9M5242D3m8HZGmsN4jRKN6kilEJ3rAULtLmG4B
jYS1gYqZnrUC5OTRVY+skiIpkzb18y625dNe7DgwVMWrSv0ma2a9sBhEPCMG
qEvsx37eMPEpnQzbnpyMG5U4hiJ9z+HUE9y+ScuBanWdjk0rEeFkcJhPDh4e
CPfu9ljy9bwR1f+0Wj2gFfjv6e6dqH3e/Qk8t924t/nCdBq/Vv1ZTj/qkx6G
b7LppJP8VXXc4aOnqJGkXBid51DnwoLh0+hAB2/ageMokrj41ZLA4Ml1klNT
5FUHC4yEPHbSc3gzWD7b3YfUpvPbsC0PbSoUAmerHYiGxfLeIP34ySyXuf3m
QyRI7BNuhQSRGYnm7E8CG0SQcuWiDEn5DttUts6cR5YXubK0SCYSPatUvlRa
KpKjt0g1tmBmV0gcBDNyz/AOYyGhMJBbfBLG8Hn+akrdg4drNVRb/F39mVS9
OSeXDi+caB5nLtA6ZEUvHXA7s/gXwiQmxfZMy03QLEb2zLFunoC5wHj1ACRn
T5x1TsYd/SqAZtHP5Gz8xdp8Wv6HqH1/HjHQYzoYigjiiovXvhKrS0pNP6f9
2uZYiw8j2g++ZiSUkZtg2EFEE9h+QVXVHDLPMlIVTV3bWS7PIsSgEetWRl96
GQqo/YaRvsqG/KEdEdkoC3eFKcr2muaP/IrQZ2xtzd3g06nt4Qb4tAyb+YZ0
XoW49kQKbP2PCO4FPy3Ybrf+OJN1iiwcun7rv8T1AIAqBGrM/61h1nA3o+rY
tXv2FbRVWUmyE8TIuT338X31IHA+tWCZ6mdOAFZ6qUg79YAnbrQotAku42sF
0w0JiPHxvtpxCIzX5/RS21MroVkjCBlqrIfEOlD93cySls6npyjj79QM7Bab
Py/imh33uJ0CYk8fboxopmOdLPiaKYJSjXrfCXifCpwfVtHSKtSi4rSaK/yM
SqUS+GK76NXtK1sn7OE2dVMq5fxLqo39226/WwOHYkxE5tClrkAKCs4FA5Gu
+42IQai6OfIQObxjSJYqWCp+XThq0o01a2vRY/3gyd6HiH/nROikllER48Xq
EOHtU6/9ByT70uUjdu5rvUGPH2jlkSWN/nJIlWmsfWAANqGONhkMWIzVuWrK
+nLa1hd7U3sRyUQ0D/EHyuBT5YXjOp+aY0TEzoutEwk4+KQeVwwJkIIuK8TF
pEA3QkXswScY465AAyPQj6J1wIg6I8l/q4l+z+WKQIpdihA1312kHKmD8seA
X8aHM92yNTx5F2zZP3P2pbdiYYCIbIGzynNEYlGFaGZk782nAZ/pWCtMFHH6
8JGJltw1YLpzdiq4/h/LTGOQS51rTKWVr71AA0PDGj4MkdEJYazSkfPFfIeY
sHt2eXgiQRoIfRWMmmbhcKMpfi/1Bbi02/Hbp7nGVO8iP/P2qCluEEaa6leW
r1tm/7kwQYtKU3L3XFuBjVUthTwmYwTEk4Vh5s22m7IYIpxtJBR4CNDkru8Y
Hsc2Pr/Ix4ldDDwV6iy0QbRkwDxa3qx/OuRxGtvNPwLqIbKFvn21SEKkFcqK
aBJvykm5fqUuyO2gL/dRe7a0vqsZ0pEs6IUmdRoXLvIexWubjuBKKA5WsJnz
IJboYV5CMTrNFl53APJiVzA2Ec89MQ1PO5xJJJ9oBeZU3xvdp/hvjUCyq4eJ
NrEMq301IUv4RaXu6aAO3s2W9fPqPtyqyI9UAoZLhPmHaj8YVOyeEDgrsBxn
l16OKgeGWAzCm9Bdyfi9StMwJgbN8abf6i3Yj401xKOhpLcyq1x3WkZ9oHem
Hidbh7hy1oAQqsB7C2PH3c+rECx+iCPpBDCzBwbL4rH7rUu0jSe/DXLCJxbg
ii0u7TyFCyPyOBzTYYT0OXCmT0nJHvfYHfe1/ba23jXn7R7MUHBDWevvvoV+
9okzBhqCB+UHAIIFOa3NNL0p1rOdWEyiIdfEXdhipXyjbb05voMTvdGmFRU1
t195j5m+q77klL6vgNOsgTwXoXfYf6UNoJW4hscelFfkW7mley0iD3Yj7nG+
xK4Zgz41vJyaBApRXLIN5mAF/1C/OBAAKWApf2pnc8QyL40x/fVBFSNhzStr
BbtCXYf3sa0a0pQU73dkr7Wgvcsv5r8AJnxsv+mSJOOPYyAlUng0l4ATkExR
Jffmntgwa7Q9mErgE/QGwNnJ/IAvzXlQk9JySWJMHvJqVXA4HRn1qZqbyAHf
V2BjMXD4/cVMt/zrNFloD4PaTwoiSdBRqQnFytCwieE1z5TpRK9DexUCZDp8
pLOhz9MuzAcWlkAveH7+TV50OYb8FcN9VRcS+j2hBBOVRezQbXK8zS7WCgoC
bFaclYiQJ101EvmiahDuOakeX9B1Xxx7HeymyUtyBKigvGEjXBtAR1KJ/9wK
zdNgEKYydASuT3SJXPPQ691mSHkDr6PFsH0/IKxobOcd3CFlMEd+FolcBQzu
pYxGMXa9bjHDQc+1R3i53cH/c8m6gu1+Qkcb6e0UFea7q9PiIsnooYH5ubuQ
M17XkLmivUmbTmWrw9ozQChAGOmRmaXkDrPq9PYg5voTotvb1D/00wLMCWPQ
9HJBZwlCgp94LwRljn2ky3R5duNtCpluHtiaZxpOpLD2j6IgANfLi2gG+rx/
odAPOjLBpezrO16lVxcWpWH71ARS1xFigDFldJXZLPGe3Ux34D4VF2ZyMa9x
Ac5aoUEdS3JjgrZ0ZHLbJl01vAXncDZyrb01jCHkhBz/XyJ9KrPkOCd7GzWD
n0HGMzZwSevxm+npDmsVvi6iUnTzmCdS9BLpM+VYop+mJ1mfF2icjITpLjiU
TywyZg5NDvs6gKpz8uOA4Z4foTkfRTAvAlh1wPpNM4qL5vrqQE9HfJPZLT6i
2WCGKEL1wIEeq579GYakejmgppPR/SxV687xCFS801jRQ4HtZI+2FsQiUlGx
j8Xf7e6k5/97duia7lhtizH3KRQUH2/6zlZvO5aHGzkW4BaAJnFw0Ec/ymiO
fBUZbjTfL/9IQIYW16DHdhO7nVDsmSBPXhr01mmOvceki8vU3WHq+didY8/f
NbKL67T15sp990vk4IdnwTO+qowZY98k/7tLcj0ncdbSObexEgx2dgatC0OA
1oiLyYQKIBY2Ym+oipstIKP7+MmA3zqNIL9IntDvQILbhSZ6UK8Lw/mXqWpa
7Cf0RppxvoS0P/tNkG87Axmv4Fw6AHYsbeXvG0w1sAkZMpF9i36T/5cW9lG9
Fkaqux0Alyd9qtIEyLJnJbVagEyC/S7uZynF3j2YEf3uh1mrFSgCxfEJjAaH
JhhkkhsYtPmHx1P9J8rn4vz4DoTEOhP3xd3+6P+l328mZHBYT0Ya1hnhMiJS
/xegdqe/W/JZKuzETAfZvhNIAYFhdgvZ1T/wstK89Pgwolx7rxU/Kt3xQV9A
Ulup5kHPYudGacGu7o5hZsgY7xn1wn+yP4VIhuaOierk0R5Jcjn+Gvwh+5Kw
tTbZaNA9lclr+D1tms8nhnKRpJCGDNehWdy3nP4DgoO46BffYQXWLhm8dDtM
P4UewPRxHozjjjpa075ovfgq6rFT6Fnkel16/44Vy5ZXEkGFPT+iEVySPqi9
cU4oXFiTA3OBYuU405BN/b8BWur6gqpyFyGXJwxUOkoWx7T0en/RVmxkvTYH
AthYS4mfsOsC5phSv3eWwY0xJ6z1urJKWJCGwqTIKZgwXEkXOyTTPlS5RQCO
llyrhZEpn+0+8u6Uf0W6F4tXJ19yeiTjqIVNz8eLaTc3sMDFAtwdUXMPqu+6
pfNSL6pPwrhRE94cZI1jdciyVBMe6HHdMeZSx9VTU0WYoRs8E3fT0VKgq7d7
rvyFa1J3yBX++3QxbO6dVskv6599m1hAVALZMOTLLbQb/R7cUm9G6ZdRQbYE
FMJfsDrsizgWNtD1qjoyxnGD/RlaeK7FNR6P+cL/VNvPpNxw37M5jiS/RGVq
alnBUgRxSf8ZvSEHd0bQanP1SVM4n+G4FSo+uIgLZkAuEN1Xr71DqyNugfX3
tMKqYj1cKSp/AK+iqjeWB+APeWE4izPMDVXRQmpMqPVMTjdYRzIkXdWyAyFd
TBzwkNhPrU48necr6BT/FJTgKAWHtP31Y/Hq/Cg98y1hb6I4csdKfV2YXYAR
+5xWwLgvy95k7wmz/djbuomyfPWoLESdhFWVbS2B2EFG9zpBvPZthCOrLd/v
GBtndJ/FA3gfU36Oudj2/5fiCqp3pwoNgzOIanqIOzTYJ/UD/WGnvwF9hcqA
2Js42Injv5A0kafx8CEj8U7n9SuU3COS7muWqa/CL1QatUMlGYp0gciC04i9
OWJ6M4WvQ7DeztLgu8RSQcHzJya37r4IFEoinVp44t0qOmQ4U1lwoThlW4mD
RwvY31/ucjL7mN0gRyl8VkMA5DVRJPo1LG9Xuu6aBnF7r4TvJhoJLY2uJ82H
2GI32vdx0ZqpXmdqyIT3GJ/Nn90refbiIB1whEM+HyX3mefxBnp6WIg9JAiH
vx+QZ31PpAbg61Z/hdjdRA7CGTXQWw1zR4Tpj1H6gJ3hk4W2qG1Vcg3IGa28
1Y+VmbQX0t/eXej0nwP+aORMdbFF1c7mvlrX29KZXUvFHfTC1i4hX8Hq8WJ5
IMul3BUPSBkAkhbBSjHNuj3FdzvSIH5mV0+L74h6P1vqf0308W/RvNaoYOMX
SHc2bU06oMFyuEY/rJlCoKnZJx983Ro0Qa90WJ2RlUYwlLwh4bucDwmq/7y1
UCipqAQeto0s2o4RC4CvFBIoOdhLiqxjmeScHxJl385nThTEwFtEJzc6MlXq
X69N1rcKUwLkmnJC2R0DZ8LKPXy0XfoGBs+z7RNuy4/XS9ohFn5G6VXAwygF
CvXgjCJVPjBiQBWTPoiyqhDAdQUVTEvOnt/by18S8zLwgzVX3HgFKoU8+HtA
q7/BiYL9Kx+20yezr0bnha+++jME7Wg0sAR5Dd47eKv0vXf0VEhyTxgzQFFY
/JV0JsRuEaloVext+NVW9cGfNFQolkI6MXbiebSCXmA7FmDCiuyMVh6WOUa9
Yg+tZ1NBqAapFDmE5+ZE8DnXnGRNS3EScetUgGEQPn1/+oSo4I/jhcjuEtou
vU06ud2IC0S1rg2OiAavUOJh0lxXHhBTkI7FmLNRxi6XC71jSbXvarWRlHAy
qVIMVJO4d1rBdTEi6ZDtNAdK1rXrK4FNVd8B0DD5p8zMZQ8QOw3e2iAQQmZ9
WWG5BxXtk8z1du7sT79JV1wZ4BJfH9Bxl8LCb+tAk96tTBlNswDMp88+Y07J
7Lo4GbdL5IcncsEYe1+TKyLT5ecUQurIZjJRZng3kR5tEhAIL5Adesg3nuGV
kD0CI44RC2xOBwjgEBR0tAkbNnVSUwGrxYyk93C57e7hmCDkE5FSVxWwOAiI
W2EbjRN+SSsWZliW4kf3MXfTb8MD4qfa277ToEzHSe1AM5NaphH7lk+7gQSr
t+lNa/TjOnIWnlWqJanH2/It/6k/PG+X5Y1UhkPMJTgU4kryPtlUnihs4lQ+
u5TWnoZbSS6e9TOxjZQSjtvItGVfaIaWU5SQZjUd4VOpWM6+8uEGC46GglN3
xehqIZPRqsO/RyygiXw9067qSqvm4SV+jBza9N8G3Rb35CpksKpE/ry9koau
h/y8PHYjVxlsTR+nLpOEd0tGzSndBSx/2DIw6+E/OvwsPhPQ4PByOJSY1EuF
O8B79Ztm4nW3gyYaq5bfQCeYA3Xw0sqMgtXv0FfGkwKnVG+XOOLkG6zVLRNe
r08xlBN+5VJJJ618Vu/IOQ1xLFfKwTJn0mV56/poxXvtohg5O/43fKkupw04
mtO3otQ6CeLjbQEL4s6Z2Uygpjm1MyoyggxCWgr0NIwbvkFGzjos4//mHosY
8Tt6eJrgY/GY4lKIAovATepMBbiC8sH+4ot55BkdoVWl5plmVQT9tFCLXqqS
3jmYguLIJFBlptTd6TevQzPGDMiYejY+HsFxOolFW6o+QIqdU76f1qMnMny5
w9YsmwrmwYRopNmeBD1A79c8+glVbBE7KuAUkOzsfFhqPsef99RWJHuyw0o0
gL1tKijR2gR0F+VQVTLXmHH9SqUPoXcdLKAbCeSeOkmc1vFgRAY486rc4KO6
dkXyOQ5h4TxlfTw7NF4uEHn7wDVpQlJN+VJDn+m7Fckle+O2yXTamdXCYKKy
pWGJ45XIgevRcjpubVHRnz0/catf/DZbAz81RgdsT3E42+PdEJydxGHSlIYN
JCThFfqSfy583n/9+PIqhAfknNvWGl8QFcqbwM8vQK44NLrOe9tjPTDsKIq6
QtMRBFTMFFwFSolx3p1puNvgjBPfJ/FiY/pDE5+iV0a2VbzAjpT2tdSmAzTw
+upPGGr0EspU+qBZxf2bbS+B7nza11R41guaNmUS+FPsE+5TtOmMpk0Ax0z/
wBcwJvfQ7g90Il2ul5/Q+Ypt3CN32ZmDs+sNxU2kJZ+baEKgvkrW9BXjXWvI
OLpnL8s7ouGtni6aGDI+XCst/2x3mLKD4yK8tmxB6OsHWC44f87jeqoMFwjF
BgQt3Kurplyq+jvLtDMzvLK33joOxk8GHPbViO/431tU259KaoDiGLDTcSSp
XSsLI4/ggdX4DGRmvuWLLA/wEyrVuOnoZZYa1QioVftucGOmqdNPnY28Q+Z8
Ju2GsAlX9KXQdH6iNFIhr6ZupCjKjWc5ImGJJ3nhiOORdsebf1/0EEXtfi+S
S2rcYxIxTCwfi0Kf364qfsEx3IQMkURtT27NtSTu1k4duIadzYsMPW5M+nsc
VMG9lB0m5FKvJWBNg9Sr7b8hq6n/K++9WJyHTas+Ivq+yL9WkS+w9o7gGA0t
sWWNZD935WrfYItLk8+6QQEkOyUy6NVMx97udC2m5IuKCEKZjSjZLls1pV0z
Z0FX4x1rA17oiS12tRfPx1mgIB3nGFL77A2cwjFHjoh0m8ggaur8dRJAdY4C
xK+wRV3j5kxTe2QmJB4rmj0qRjLIrSPDR1m4ZT0NQ5EoO8joT6tClko7dlu/
fv+UeRqdl7qbw0tvCHAPM2bdgWmfhLDCYN3+OnOE2u4ZXdkqSNJNL+inXuhY
S4QswpgtDqVWzH+MlNFAyy7Ab0kH0w5l5IKo7S50R34kjj3tmx9dnEDkgoGx
mWD6qPnVl2UPxhlxV7//qwT6/cR3whqxm0W6CJWzxXNkbXYc8Yj6Qr9dzF41
fgV9fMk6R2WId8ul26GhwLrk+Go4QNj0VqvWbo3y0bxTokUccDsHvfGlHXUd
i7oNMbY9J6i4frziQIYay5BSa+c/vsU+CIpLBzFQ1N+QvTNsYqOnGlsXKi0L
6LmmzR4U4O5ujF05tpQfoexCFg37zFddwSZG1Gux0Z9pBQwDhqHipaeGsvAv
TlutjBpMhnAp9nY0nKPbdVJY+o/aOqpQmuzia+rKwuujav7zoFE7FzC5GpJG
XBxN+Vw3Aw3XJNaErXQhzUj7p6kc+dVhjvdDNztuz2A+h5CpMHBj8WuAPvT3
Hm9ODQKqUPyCDi/F3sNVrZQJWhkGQ6DgH7zQjp1IP+XqwJD3gD938YSL3AJH
3MxOjpL7+jlPYwEUATIe9hG31I7bZc8kvCwFl5Zr+0n4BlUIm6s5MQeJgqqh
f9123YaqoqX9guuV0BMvv3ZGo6CgF90ug+VCuI0OqrMNmR0gwKNHwNnLeLYB
4GwDQ0MGCyi6Ssb8YrvrPldesjmtfHk8SU8f+vLmhgtwQfBpoiP5lOvg7zez
KpiP+hnwPksO9ol1lbQ0YHpKNvlyn9Vyp9RNPYbqpeJqORn6fawysZdfczaq
uPChiUIPqd8j9j4imeHXoDvcko5qFYhwtN5fO/wNLrKYs/Mp4+LO+6mOUWn9
yiZHo9ACV22ByCENgK8yUB16hbEjtW0/UZALYtKeISLWNot4CtARQsaoAo+p
LCjjbV1V8SMiD6Z8CEYOmn9HhfB6kq8LtC0jGdZvw+vd9JniHlzKq8Big5Sl
kdCrdpIPtLRPeabOb4POwWzLm7OBAcMGf+YuGVPBa2zw/IkJzufTrNSUBzrk
0Eau1Z8On8KgV+sn+3LS3OdbLsLpJSHBGlN5zP+nQ44n0/Oyq++t3r5QLPkC
uPI2rvW72vi4tOcgCCC4vd7BKAWoebaAhpbAurakZPo0S1IcPerBCpiYGn5S
QAHIJtqzROT3QylSXUw26TyCUR69gDy5sStm5pWiPQBXz8hEIHc3Cimm94Mq
K6UzXtUv2ES0MEZ8/Z1b/DPO4MxCiK0wOfKGcn0mg+72nE1ITXGdOzo2PEPU
l9w5RK9tRk09pfPL1yiNGlAJH6lLn/hL6fjMYPJJRjxwLGnAIHtNfBAgHWkP
bCyPYD932okU4uGUSNXVmlUUs7gZ/4IP+FyhusWS5y66V6ZHnxVuZpDlwzKt
5Etrj0Ysn9MDxLGS4/jc1hpzGv9v1uGIoglcdHcM7RINXwQaqVYc5LA1Dh4x
zIhpsshcF/ndccYdUa7garZ0hEw1mcFxGJGm3fTWw5vCLoslCC0ipWS3olYJ
v/Jz761Ps2/HKDzlnAOz2TS4NdUegEtumJJokhoO9hVGdQEP+mMtWOhR2cqV
/i8600Fwjyt3ukZSUotqaaqj/GCYF6bABGmrFZtcLksu6nV7EAJqqV4SVX+a
PfOW6lKXabA1/s6ZCOmlztwMx6O7W4ebkRgOzI5vhCFdvgUn1ODN6YkloMXu
+B+TWxGzTUCcFI7smF1vE2P7b09kHGJSzdkl5JEuzZHR+Y2cDdY53QpwexeN
K/ux63ch0EZX7x/EXrnsWCojmj1DNpO+52/3PhDzPL1TF08Gu+z+XilYHV3H
AVignq0Ve1OyYYWPt0SKrbf4sbPOTqwU4YM4+SN/a/TWb8qPp1UwVFBpd1GQ
0wc975liDApVI4ohJXFuHf9d2iMJMzHPxLnka340OsiwmdUSfI39ynVk9NxX
yAW1JiOlShdKYnyhWoT1qRUm7/TL4qMqM8S4f6nVfHousc6e103q6ALvBV2V
d4X7VXg2ODwYbBybP0f6zeSPwgafyBJE42yidJErj8LNvurghnf5/6lwJ4ts
OESwQsO0HoEJcGYOif2+Bx7/0+od2xFb2DP+gsuV4r7vGR0hYvjR9m3MNxoP
Y4HgUQvleSUtKXilG7yM29zIUsPz8ch8ckEwZDYEqiSBGTTax5lHOqi2Id6v
N+RxF4gZZwqwNDI9EDEjRoD/J3VGjhH3B29nLJZdSe+0Os4+dWmf8Dxm2yGg
B87rHMEE4TQYTJ6HV27Ttkm4ZqlJ5KgIAzKpbtzyohvEYq+VJdTwbhhWtmFK
QNMkCD5UO03Lz+lqGmsG0RH3GCOtkrBd5kTfCb8O5WoC6VAy8yzof7biq6ip
1GLDHGJaBoWUuDFXzwxIo+/0mfBZf1Sp0DQCptFoSrJ1aGZymnDUKrLPYp5Y
bla4O0RPWotT4RolaRI9nlrO1M+/hSASI3KeSh43lIZTX+uZuAEC1T/uSN6U
vr+1DiwVy0YrlghaeISt3w7jWEuaWhjj5+CmRMlyoCQYjMU5FMVe5nqFvYFX
Juy0bCEhS6G3y67OLxijan40kLrEom4RcZBUc2y8FOmxg60mgVyyHB3a9jD8
8xu0P61UpA0YJlCfm992zk/nxJBMkgKqD/DwVYVWrS0WTzsqecOCItbj9H9B
NBoSonhE3nRpak8yfEzt8wRjUNe51miF24o3wzSHiH5t6+SoO++Da7cjWn0K
dN0mnmPkQ9kEMDqiPGWYHsBM0xNrC0aZbd1IqGXR2hLk3SwP2egy+0EX/71J
gJAuamY1doPT3cAH12eJetLgYuiE/qPftcj8FPs8D9knYEOb6WId22t688e7
kK86y148nFtEeQPURGQ8/rwAp8Fq6Z/GM0Gw7VX/OzBvicniErT5zJqG2ZRe
a3V6zs6oE9nE5p9EaMzJ+9rj50nEjjFeKheZT9fMqjVhbLeYXZZWsHSIDkkC
CfaaRIcqCh9562IH8OPnd1ZbCR6FwelV5meBY7+878bcwlRqFnwK/z467tIQ
90zREGr2dNYaLA06eFa4J1LE9KBPuvTovU9nGwfgAYIlV/HLjxEZ8CeEnCLZ
PiNFeiEeIhb3txnmeN/N5k6fHq5IL9is9U/G09E6nkERBiROTcfXiLXZTFDS
QEaUbq706LGHOF43eV+XhWHoPMh2fG0NdjbNVyhO46dCsJlhdmCAPqA2eFB/
Xt+I7l2Uxq9wF55wT6/pq2ZCfuAEEVcpAi7JM3CM2OIiobRzHYyrXwuYpR/7
fs9lJc/XPXeIcKSD/gsNU6tDymLUK3kbe7jFWlmmQd3+gG9kbFx1Q86FOI4E
dnrE9LCUU0MRCx6XVeL6P8Sy+sq72GqXb5vx+0/zwea/cpv6HV+IGF6GjXpK
iT1keapmVaNCWcwM/It/ddbo8fEwHuxXZVQPcQoTvlyDIBBlAXmf9WHxDqPU
8APvbkppREYKW7xja0vPaTkKNemNqSyLKRPPC67jbDlSLsvNZwvwOE8ecPAs
Dz7rildvUQng1fOmkjRZJC7gP0voX4SyOCPdDQZ0c9djXyKJ9zJE0ZUXYqKv
PA2PN8tA7m5Xdh4DQTYEFuImVynLFch07HPVOOBHF4pfL8//AplBQGm4C+pm
qxdKIV9ImyszHPmhiGT2FtxcUigKC1QBGCZAgeSDPnXKn4LWVM72JthCE37t
4yH7ueMqf1oOYOgvEdMbc49KE6bBRhzVwD0oY0MH352vMf+kbqF2aUC/0L1o
Y77VAhQ7r8yiyL2CV5QXJNBdRWCUM6RCtjcxijdcxeQnj3Za74N3a4z1Resm
6g5yInADRiN3gp/yfwKF64BsKhriDMWqMmG41FkhZZhZJ1ZOcsSrlNLVqzAi
e6GY811kqDnxEChUgW2UVhEa5yFZz/olUyB4NnYrt16qbU3v9nGxAGnXotxn
aW06PDF2lPGMiF8KuCyEfp8xh+G6BDoHbCMayLNWtt9mf9LBCKIlu8aiZqdc
EtU21tPKpgtzz52iAZSZQUOj4GNVuz8SzDwMIwiiqL53KjmJkYPdSoWCEOUY
ayac/oR6CyQrWoWUiZK5C+jnAJaUgMpUx0CpUPtsy9iv36SyjbmfsVyOBZTf
aFcxrlmSkDuUp9WuOzmFqbxLldl2HAbcMupHvlH9g/YMemBYbHVDHwVN4kSO
Ng08Xis542WliYKxf6RnLN1AFrRtBcmRHdgr3/JBIXyqQdNJuAn53im6oSYB
AwHIHXgWkwgQ31/RnswDJc6SeChKf+iC6hfbAEwnWlXAcoC/hWrDnrmBERST
0qKiWimOKIdzboAV8+gAvYLA9i3/r8NPgImGGN1sI4Nt37FgRSKdQjXllFIB
FG3MWamld/k+mrQxqkXiNqxPIEEeeLuOZi2uA8J8IrEq+E/iTP7r7Kr/Cfb/
HM/CrbaX48dR+Z1DNeVe5rVtgJEPyYRBg7pFMDu7qxWsiiMDlTlJKseY8wll
a4WsCAnUyLCF1dNB9uhQJwDs5ENRrrLKUIAY6IctVn84MXxEUfvgp8iTNw4X
H2HSDZrmxCvkDA5HWL+GFDZq56O6fycgyhX9NE9cwfz3rkyYEbpOBXutECV/
6gcjms9KTL9YLSOip5AqKFJwSLBpJUygrOkMKohC7c1W83Db7anxw88yGA26
dA90I+j1QLLuz+Iglb4H09H2ARp27jNiaoU3fJdzr/jWz22ozzz7vAMBH9hr
JXBHyZJRcad6UqWupm1tcPhn1VWL3OP/o49kN6nh5YFkEWD1d4eof7n+T0NH
fORyuSoe+vP/lIr8ME1o1qWl08BeHjSAULofJ+cwcTCR+fGno0TeJ4sqq2az
M5hSZqBMBUU4Q14Ll1AbDaPblOwKL7oWXgvOYwwFqA3S/uH5+SPNkG3cO3sR
bukbOCjv0D/wWeOCcawJYoR2pCyGk5frjQ3meSCegPC2PmL7gdJKd1UbXUJ7
VKY5YBnwTVotbYyyNuOqChpzD7t/8ppRETqAADqsHr8oUqiTps7SY+TUgpMm
/kdWBQzxMSWtKZgSQ3+pqj07dly++4bgSEJz0xBjrS0u5U6lhCyfxbRp//6q
yeNZH3wXVg9n12cficVE68Ft2nTvlsxut81b4IdtyzuSs2u0dZYls7WALu2K
QZxyLOlcnpmGfkdHg7R0KiARNyFxrMaA46xj5jgVl6iiY9S2uXN7jJ9/2IEA
vePscSkA/61MzxiOQZtcVzvLkKIBGZAuNIHYRe6Udrk+OU3z2VY3qtHz0aMV
laUb4rsGjOv/bk3OkViym7V9a8k/D+ZqwdHW2uDNIyIzuHZm02IrWAmslU2Y
2w0JJk8etvHGzSlmkiSu6/timb1+BEBiwPDMDEjXyfI5m2QaCSTcw466YX3n
LqrBz2eeNwqW+eHjRXJY/L+X6Q+6ZlNSGEQGJVNly0pO464c1vaUq8CKcADB
PYtVeVuz541bxJ1MHrA+h9wLT+uK3ED6e2RSd4bSda7ElgduwYosjx9mVloc
u9eKLfNxZKnla69JtvWfK/ZB/5XD2c63QS6g6JXyxFSZGc5zvDwz3+D+32bm
BerN4PH12IBXb3sx6jrDNKf92wDBPvR8NJQLoG6fyrWZ9kTEHBanKb1044/r
b4PLU7TxJxaj+r/xFdM7oBiCh+0FTKy9VDTj5R/QeJrYAOWKFGiV0KbSZSjz
GpY6VEnr4lkR8ckAeTzGmJOao2gjcFIcvaEHagIKANwkBDs0zKy5lKHPY3dN
C9CevKpLwHpQXHx4KVNAjhzx1egVYCfnfg20pgKHizIx+SFHD+CCmNtzbRuL
zZ2samZXLV1nVk8RBH/3nTGQzD0a+DlA47uOsmxzxdIpCGVg6yqg5sHDPWFt
ZF4LOWnZkh8IwUfTBAGsFv3PAEff22zOGgPWkDyOCYzSFznCsYK3tTnNv4V6
fFILC4CY81f6/PSRdYZuX3sy4yB9OuRjnetQBw3NnE2trdiQOxWXE4o4RVOj
DcHjq/wIhRiXz5NwN1uWoEcxjAQnWAJUNJuWHp1h+IGlkxWkcBJH872qo3fs
vBznzYQfZnuKJGI60LhLJmF5REQj0gclKlJcRBSthFeteMA/hBHNpsK5eZ4d
C9E8KPri5msFr6aZnK/BqDpNkQaEhaRJYALDEyuI5rWRHeuCqwsfzo4vYapq
goUVniNvCfIR0NN1NErtCuDzvsc7oXll5tgYfvAR6ET0TooHsnI2Outbzevg
ja2fSanRCJeoG9HkMl/oW5p4b0UPwGPEoXhKqeWDMdgkj2GZ4fNhKs3wp5cE
fn0fcq1B2ypTn3ECIrxTDHrgbpRQskIq2HeOYVAPvarIQBmJ2UjY6lq8c8th
cGqJz7VYekxc0cgL5Qmrr8TLufo3AIEWXvkjnceBm2UvCuMu8KrDJnaETT0P
F+FbOEKhJliFnAmbmX4S62jkvMJGBTw4vWhm6Tcd36ytMsNV41GesU1YmeA=

`pragma protect end_protected
