// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
TpVhg4b9T+6JAlhgsyjI3lJPvrL/sZfp3HuBIpy370S/MTbGqtlOrsyL17xp8geO
9lulyppGbE2CRx6DzIw6Y9FdZf5iggdOnKqkWJTkhAy66fWOjGVpqAopz86Nzyf2
lNh96ttohACJBuVSuRWIS+kPM2q2vZQ+2kSOS43Qm6I=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 10512 )
`pragma protect data_block
Z6H+4W1nUUdlCyVn9u2gcbGrul1qf0dafjKDHkSZ7EOqy/x94GMlK7s4knhmNFZk
DwBkuuGq5hagVFq4rsNsbvoIcI4u4G4Gy5dc0Q3ISEY08P47IeAp5B34oypcJ6jw
xJndHzUEaGQVJwfgNgpTDmm2WAFoKExON0ipn0yt9ORigJVBgn4hv6MryHTM9MS1
P98GY7BFNGB3UW7WVkDsGr86/weaXube5cB0Icn/3nlJMP7V9TvSE6tryMQ0LpDB
Lynv3gUfOwVNSacdbw3MXf07A1Ygjn9nMvGuqungnZooVt24r2j1tzT6SfKgQ4D+
xnvUDQRFrfdojPKeAV5CiOT9lQObvolWn1OJPHuXgxAeB5gt0oBPtsZvyZB9r5OL
3oektspG/M8orCnBDJTAGOhonSDBBojc2EVUMRFxD5SPo7v1R88IRjQjWQS7CgYA
GB3S9a/ISxBb0fi4PxTyMxXSZuoj7KYZS5IB30t9ugOuuDneXlpgnnAZLoJRxviX
d50t+5IciwKx8aIjiDDPiPxNao92qN2s/0AO4gOijKIMtgL236tFVrDkFeuT5Wd9
aUQ2TwOzXXYhHAQ6pH8BUzp5aGEbsHGRNng6QIqW6Q0tASvc0I4iWWs+Xrd4iTbl
v9HQ3Gu4FyKGYYaezilVa7J/uD0rUqpMqb9wDxbPego28+PQpX8gRNwc6/ROSIHz
QHwdVL0wFceA+5kqtdt+Yeg5QpzUTVJ3VS0YrFMyesL14Isx/mNc+66BRt8sdYbb
0xu+LSsmz0j1yYxTdCfvWLOEIjk7rzgoHcz0/MaXjBlyDK+c/rwgObwBblAeGedf
vKlsqtd4EO8YlK+YAbM/OW2t/pCCJcme3GkHigeWVu69uFXPsgWSUcvcqBwPuNMx
6EBa1AHLEizhCTw0THoFgYDtPRyhrPa6WQlImYvpDf2LkA3JzUK2bXTz0vLHEz7p
BbrQQQsFCr5LmTc8PdFZgz5XSQeFAd/oE7Pm1dAKGbuiZa9N/Ne5wrfeBbLxnvRv
+TW366FdVgndHiER5O8n40M3404nR30MhjYtQwqg4dS0iz7XhERH0UrpmGUBsKbz
qDmXpO7qM3GfdD8K2hAqQcE7SWkifMKT7BDLIi7CQqbzi2YFZcOE/oJfxeIqpJEg
c/Fy1hCRi85At+I0LP3kEh/lpIP2vwucAYL0U82IrUpQfPKakOjilLkFMBYIYUfT
j4PQ2+zOlhDZb6o1igEw9w2ULax+cUCAKGlisfSFoZjHIK0xPCe8QWuzfvMqhibw
b4Bx5dUJWr8ltGBIu/3B+nq72EBMNAI0O1nEaGgk/FPEbtAUzDqd+BJ/A1+9KP5D
UqsVDQpTm2BqE/Azl9spNllOfcHdIsdhll0EdaRSpOlvTVVPHlJJvG5uH2j/64im
DhXAYyIfVei4IEkj8Co6KNP8UhdW3HtuObIKBVAzemhgxAaidn8jojN1+MI5znBV
9umtXagX/yjnBItIK0u8ApBLaXDWdt7iaQs9rBfr8aCtc8N9oq37kRSKFsf/nAko
dxL6mBVYCFB7V+GmTLvz6WFk1yq7gwkTRQpR39tMlQE+A50RnOoBnZXHxo8gdE5v
x+7bNV4rp6/S2104PN/mWFX6aeGbUMXGVOJ6qGHpN/gKyyrMXrefbP3TdglVuxwN
pyjEe/OipfnmefZamOaIpVX3VBh2ynKUtJUNUyHXaFhvhiHaJ/hI98x0xjFqL990
ZYAUlsed6YJN6cK/mMo/vjvCz+zHP2QGs7m41KIUlU2GlOBkB+zMfVFczyRSPMV4
em7WRbaiE/Gvek7flriAlEbuFrgnarXC8+B/GycAeF5kEXRC0MuPttNF3GqEEe0E
4u5Au5F5dT+/CWzpYbTqIVDNxNYjwCSgjJIsZKL8A7SPC3VrDtZ/FsyMvI51HzOp
ayT6YslZ5gO9ZjRmIa84tfU6cCWp1jcjNc87vZ07ltkN9bFaajtMkCkfm1ksC4UB
4EqQlttzNk9lLUVzb3A67276vhieeDvVx1KJvvlc2fEMUW+/4Az1copp1sTANGfX
TAXYf6bEUAjW+kxwG9aUe7tdHNEI43rYr/tzd6Vdmx/IieRgs10lA0SGPscroBD1
4bQyCM3g0g3a0zxYQmulr0jPy9DLwVlqkmAD8mtgP8K5kWK8kk0XBUR0u6W07dUK
HQnWfKATSIy1DteVgKoTnrHukpC70qcS7EZVV0qd8lIW16F9kVao0dGrusCRPPCt
YXldLUBAbRw9O0ojDoKyOTAbqrdUASPJ7Xe2XSXCNpv0rHw63pPvsDioysr8V/6F
jYkLkZkP1IrjF4xcElfQqB59DHo8JiJHatu4TgCcAIN3Ly4mv0wg4xtX9hnoQlM3
YJEfVtomvkWPXZv1RyNlELZdJ+UjhcI93Z9rqlnd1UB9PeyBpTZLXCu+EShQ69sJ
pkOQA5bAHqwXVhQLuOK0EFZmtDk0vvUK7y9nyZnxCQApi/21Fl+P4blVRvh7cjET
ym6jN8ZYeZR4aeiV2qF5eFDhUxPbS9040mIlq2xg6H/Wf/NJKVyFroP61Fe3DNSp
tSZiPwievWsdR8kKlOoj3ylkoAd0OfuWFgHpOcLpg6reaoZioWwoJojjjqjFNNTk
ZUcoLIoecMyvLyd7KF81N5HuEN0xTRE6HxMe9wqGM5n8P+bxT2egyi07fGn2jHsv
w5oRviAq+69+FKLioKU6Auhb3noStLdff7LLzhQRy68vGSg+zqAzo+FQK4WXo84h
DL66oabdCRStLTjNDsdqBSa9AduI16cy4uMQb6MOIUhuGvezITMCp1M8OLHlu6wa
jAU8mix3TfCBmv6BA7ijuH0eolFTVZvFOimF4AOrqNLhTLXsiSr64aEhCzw7mS6d
59y6YlGxTyj/HI5Xr8kdvNNuOWl1bsNkoJgdqRf9c9RXsGJ2GobmpAwx1I3mPc0W
tzQTSyyIt0JoRVXHqI0qh81+gTIdX2NcObAM2MP3TUg6O5NnnR+hJFPDKScKMO2T
KyLp1BcJQelr/7Wk1Iece46i7hL0VKLrd9mPJYP3gZKYbL/k61u1GopkyZNdicKO
ramcu54eAjyw1HL6V/jKk/LWFwi1Tuwf5y5Z66uQ+/DgAHue8CJvFWiQxy9Le9cG
A75u8Vq6NiIpZ++pXhQXySRxnLr+9Zb+UyHIqL6GpbzEiO8FnK3tW48gAe7F4ITp
/u7dE+XsAi4P1xNyRAVTl0aFvxW8wMVDVZioXEzOuj/b8BvGNCUNmL+vfEQeXb4w
GuJEFW+oFq+nyMxY73BDey/zCtaQVirmfslYXoCvIsmjp9DgnOrSf0mytCS+8qXX
oAK37HMMS3/wDnBIob3zNTv11m3b4arUNCf4o0nJR299n+vKQMPa9eEHaS9PWo+s
uOInEg643w2o2PAg6bjojjOwcypA3RkndNXsSZRFLIPrv6/OyTC4vrbNsP4xAJNA
r8wVbFt32iSUhYs+P2S9uLkrsKGYdsd6yipTX1ylzn9JTp1yTPanOjlB+M+EGK4c
k3H0wPCIqjBYk1MzW3EDG50hyjTguvS7jaxgss69RM4Q/ifvclC3cunRDWFmKvt+
4J7Pp8lfLNSuO5Kl+8f2QrZqk7R4b10dRE4RQLpNz/Sday9xk/b7UqrS1o029dJs
s7r1RT0nNKgCLi3XUzX8IcxutU0G1+3TrjxnrHll02d66pZXzr0CVDbcCey+XoSg
1PkKgk+An5hC0Hlp1+jSDrZJL69bcBdHOJGgJ1F5S+s+cpEqu9RN808UoX3qfog+
OzE5waVDSUdeOMeHBWLfaZb4palBKFBVyOD9TWpcMcOSWcdHbZWXDGmL3Kr/f1gI
2rQU1HNKt2W+vXV+HqQN5mZPU4+1ESP1fyyvLxIt61ocLKlYmOsNEF4nCjL5wWnh
ZdvlfBcUxd8n1ZeAvfaP7ccOdmqVTYhhiZCcH0Xvno/bs7Sc123DLFC5n5TJ/swb
30qj/Hke2n87a48lneVEVsIyGlH6AIMFQXsLLzJkpJqmYtLkJHAfMG9aYu55WlC/
uIOFlMEthEXfHxODVU96rlWan+zyLNGfEf8wdEKp6PlLCddTrJf2CCZfFSitnrjd
9SdEZm1vHk4YAbhagUI8CkSoY1U+pG1dj6ISKbsUOBr+tP3bKL0YWQpzkzebBkWs
pqZ8He7SdX28W/C+4mt6Nj3Sed3NORqLFEnew98Wm/hI3RFRoF1U/Q9zeYx0WCbb
g/XoeI+Jjy+l3om9xy/EIjq19iY5oXhfdRTo8SifcNKkZDd75qXhwybe8XRBmH8G
Sh0ppbCjWx7jx612e68LtfC9t6cgh2JZno2CZTxxNq5vJp8KeHyxiMzYE87Q/yeu
C1VpnaZIerewrQufeWQjnMHXwmdf8/BtrHXXo/yh3ShY1E82XUu3puZenqet9xFq
IEWCV1zCicARmwSPPHTpogFU5u+tpyeUVmrvutyXdvJ2y5GHEcMlUuNnVI3zMVPI
SihcvkUWWxuC+TzaQrsZI4ErE5N7FFNR/HRaT9VtmL/WcIlaOj16EDTsXsjqVyq1
aGbhxJtsQgZcJHx2U3h18KObkVtSSf1ymMtd6gBUrAFWTYhDJ5X8vrhdM/5YPXvW
rf19RADzTwUSXWnKwHJv/o3H+/SJ87ZnH1N++TdsRkmjLQ9VVabWqf3SFJ/vmvPW
eKnMribjAglDzCYWAY1H/8PzckXQXCdUjW3ySIsBKb9RP9i8wP2/SleFqdDwn5IP
6XUVmfEPiJ4cqajxWksKj3xAayAAUSWzr21o2PHLUQB9ABeOsn2rPgSVFm5DepHJ
KYxwLyhLcxbWZxSOofWIeE2hd29SlyTWi5ezTpLiYWdQ0xJN2cI0Bw8laTDWo8JX
lJUhiLmOZdGGjUXLceznVXQcT51nyAeDtkjxcsTIyG0KRuci3ztJCY4ZvcwJ3RYP
eyrMj57DcYK6Ghz0BKZlMdUrxPiydbhdqzmnCiEZ5sFiAUysvLOKC9qt6hvK5z3C
NgtLEvKOb5GxbC53wYAW9yxiuSA2rF4a1AlF1enGfBouuZaxAu5uC/AsfAAX3pXN
QkNy8xslR/y4A+hnPccb1fgFb1Pmw3P5MYSG/so3/ehipZIMu+c0x+a0InrhzBAa
OnVTP2OqFquqGaBdrUc5K8nHrNzrFEic1MSS6xqAuOwz6L5keKy3lfAwLGnmErs8
iwn3K0k8ZT2cHAi/LVtQtTdKw6Ub6mMXViYDoKESWeT+LHKKbgMSW4+Y/hlu+e0n
xPjgRO5t8xk+t1MWuAIR/FR4och87kVDLGwUugGqu2bWsEMtNus+uikyTpOdecg0
yDirTE8YjsMdunES+Eu9UirFYdcB+womPhzEPRVV9NDI3AhVfhZcCqybL+Zs9I1x
jKmg7pXuJ/gSNEDShB14G1OCIygMRFpXNS2kG9WyObm+PhKB+HbpwWszrL5/tbaL
hfONntHWOsgMZAYX6BgsvdPeBSnLuUNjFuukUPB7zixZG53jErfEIpcRABm6dZtM
vZJ7Zo7915nxph47TuiQ0qLPIkS0LoiT7ZUrQL340KY1C+FUKdoo8Xff2Hr80QmE
cy1y7/tZrXJvm0/YUUQBshCbZak+mj9SnjPJR4sm2faA+onmDI1N+ryq0SEUYLaz
i5E/pzm9Mihv2dbtAuwnW8SvAX1pDctEnC9cMFMFPC5/AoR7IuqTnShFQinetaKq
WIQcGKl+GC7n5RKKgPfBSDH3SI38rkIumbMt93Xp3XlYpe2b3G+m9P61OLoHOwR5
wwEj59maTaPZShsFN/9BVPsFAwdsaYhW4RN1LNjMM4fnb8Uo9gFcBO4AldmVjbj7
ZA7N1JGzbuUH+jac+g/VqXoyDCbeKMxNKAU3Fz/SO6CKnKpSYrfmygD+A0IMj2aK
3mqBj5vSbx5awb3RgdLTAlOzoWGGBaJERe5XurvCNPScIWS0tLrkD8cqi8Ige+qT
d8vcUEttArwwKkDmXbdpvMAxzhHo18Y5nrCE8aLEaAkyKf3I1omarqAwcCEd1yV9
s6zPIj3Qvy1TboScCbWhXJ4fRc45OUCMRDgF6psr7ABBk3lQFv2oQyIR0BdjgCyU
NLzAiC+cE7/WFX7t0WhW4T7VWl5QWYJLvBGID3C7ENr8adFOj2IZ/DwHkGX/9jVa
pPmWVXN/1yIwqSJvo2yv5oIkPhAe5F6IB5dWk7NeKp0JLHl5Zm13nUEK3xdZnWh5
JqZtV5aXkdivu9E+kY58woFFkdyOKEUw/u7A9nxJNxIBrtMpX6NPdWaoWkqcNkfP
IbIQ43sO0I+Senl53idKpS+LhLpPGT7syI0PGtrSZ9/IUQUyIPIw8Fbobp6s2ZUF
p0DrIKIgAoAy4PwDG3mLoF/Iz+Ms2Yul2J6lze3vE6u6YhMnJWbcmcqqjM6dZmNe
5t7DLg/wUR21jYDOZH03ysgWYsJ0/cy6y4qLvtgTbko+aWCz3cZNVqVfS3hhNoTA
DR3bWUyCbD3nKL3Ij4ooGrqgZ7CwdZ/2eOrtfK1vttefX8rxbWteS8iT9/CePrj0
TOVynLbyBG8PkvQAqjwI/WpUcKg7kyQfL0iGJO2KldwEpZi3DPn0g/BKnVGqnMw+
Srawf93rghHDwnexMe6MtaJwFOUFUu/0/D+NaNMCP3qbUhb9eD5GOV8kPo+QyYBN
21c9eavwgUSHi/knZg77KCXmq0PaqCpdv10g4l0HKw2r/9HMPbzZWd1vejMtSKQh
QA7ifJCmKNUsthSx4VBU753leMju3SzONSG+JzOytCj48RzAt1ky4qC8UnHSbrwv
uaQRWAfZq3xfxXFcanHclTyCkoUDMkoy4fSSX5oAPs4Cu6bIgd9EbQ50WLatO6Xp
Wl3PmpTygFUqrx/ytvNoKW/ncZErm3K7NZ6F7s+RSYjtfU02bEqPavYMaGNult5S
qHzAgkeLNu8Pc2AgrprrKQyHNFav8K47GAD7P5B9Ac6/iCIWiLJT3tnvfyQcjeIT
IneykpRy95TPcwrMnb3OcMqkOvNNeoVeiUPpwsuwLtePNNEe9sKAfaUWYaqyKQDi
8batBPVsVT+jhrj5eL76F+u1fWzeGN5n2nkJaNUYfLBhCw5OxMh2sPZ1iOqDNPPF
i/qIYRAPfiLD4QFPSxGa9SAQTbj+ywrh95IJ3QAPWibFCyHgGcE6uduOfLou3JMl
h66hlc/XgwmZt9RuXpcg+dsFXG/GT22PRFLHkIYxhDFcSlLALNSJByxnCx4Slpxz
bccIjriVQHaQMAlZPiymX/GoqxCC5bZiGRI+4tA4NhyRaWGMFa1K1R1gQsmQaqyy
1mgr+feVwVYNc9/Sa3MsAYQbnJavbR6vPq04E0P03S8HfxvAmHruBOk9KuOTflWI
dgc5H26419Pu1iY0bkBV8tuquGUMD1RMoIuonp4surygb+PypLaRVKdNAJa2ZT8x
XZyQnHpV8+HUKx44+bNcCt4iqzBdDcc6JrvXdo3oOPx6KA5ZN+1CWfMIqCNWSht9
iW7H+zM0K0YqCUpvnB0zgdTyPVzhjqtvIFJwSVzLrReFgTB2R6bOcAWP/yDq2o/o
cBXZSCljtRZoSpdiwY+lNknBziB3sAzQh45OFUWlSMiBkvhZxRku/PxpzIwv5EMo
C48fPLzaFOpJYpvhJs8TTTdll/sZQ1LRs/sWUxa3EP7kUHPUZ2AR5X+5HpowSha7
N+IyxIIJ2cMtVHFhZ8qI/B6Aig7UIy2DrwTPPEdpW7p01MmYpep6Flet7+dIC1tl
IUhE3R2Voe46Qz2kftQ+/gsqN7P07l+EJd+nfWtls9ZxrEjV8Zy/T355MRjs+aHg
Fp72ZFwx4Dsjn7u13/vnyAIN0L0e7CTVtzHDvHUQFHIjbu/NHP+Z0QO7OHIiWlMB
Z99auEadrQ4uJOV+PV2Qd2G2/e5M6pGChnEieOWiKCvGSjvoe3VDLt6I9KbDj4PR
MV3SV9HyWMJg1JpK61UaCGpoO/o+RM5rkpOjxfAeAkeXqMl0rCwQXjgPHA+gM34Y
P6aka1fWpAcXQnasm6Xz5l2uZ7lhvL+javjurp7J9mw9UbU7UaC9CsObhQVzAF6x
56qQeAFRveb0/wBLUMtOqX0BokoABgGO+6cdK1yKXaq0Qe3uHTmuc3pE4EyNTAbJ
M/6RpHMK2wnjJeX39xkkwKEmgjUGLqf/PUKHt4X/4i9qWQn2rdk2so84hO18AQEQ
IoHVrGiNpUYPacF0nJj2ZFcHBlNcCiNUAhtHyRmm7RlwymdnnVzpBKbr/GZx3gkR
BZjwq68w/Qjn9Rbt0jSTZuAsPwYx+xZIKsMX7p41uscvTd1SefQ+2PHpZ36gkXgr
G+pSxDOlNvwQZ92ldt0nFsrHcGYGp7Rqgab7h/Xze7vsgE8CEk7VIQjIIjujhaWe
ttS35vFRfcwvU7Un+/0tv95mKXjcbe+4tfb5AG3K1kdYmU17PpAFcalwkPxeMsyz
dWIiPHvXfNzzDeQaad15i+6/T+qyZ7lHiHeWPbHimc+Vejnkw3HzR4TOVUNlbDhJ
2FU901Jn0nj+kj8zbEY8Y3rMU7w0AgwnkVBQn0gfUNFiPeCp4kAA+bUJ5cT9Msg5
Sob3wZXFspeObQ2I3SiVo/zfn6IGvjyHeqZcH9CTvyPDRs2tKnutXkDnoD7xufme
eZKOzcdB8JW0ysCbMkjrK0wKh/bxIDrO9HcTA1vN7SjmStnI7Sd0G9Ob3aiUXP/k
9dtve7qfWBn9WdTANhnamu2pkt7qmKzLVgv9kInCZvHMnIaAaszGPJ5aLUJ7nKPI
ltEFNVHJefFlKt3D73cJQIupy6J7DV0/2lrghGkYGE2LH/GQX2E01pTKF/dcAfdd
0R33CCQhgGtwGjJ08lvdew9MeY4hfvQSA34cBDcjnoQ4FzQ9CBOLfyQf7pj499gM
uRsXwOw+iZ1LAv0IbdkUUAbrajfO5ChiVNEyzLQp6/r6S8Lef8d7L9x9fMaoaDm/
VxYUPWBs5KGGTaVwH84n5LETkan9uaxoGfy1EOKIzUGKGDC6Yxtm5htt+bHbiEaa
yLsktsVeo0EM21SSR95s09RtnUtH3cyv6S62HItw0Ul0BUMGbbTzQr873xMvTniE
oJYjA20ZhsfdB87Sn44IQTgIfPOXxT82OJmuWBoEkuFLhoXFhvCtxYw8jxiUdliq
vO0496ps01s9VTxgyaZAGu2rsXgd8sEwwta4T8db+C3+dScCKPv4ITRzHJoHLATa
LwQHKSD/rxQ9rsxpV4jBzMMwdUdu19Z7CmSsCIwum3uBOvXthnRL5QasUGiOwCB+
wc9M3toRwiiKx1M61LKcK00mdgU5xeTkmhfGVjHCpZL7vwEpCgKHpEUtZKqeuq9A
QV2qfHnil90rYrrhwisOgzSNtXljRepOkDRhwXV5QiUHnWH8bzlGjMCzx8vXxhJs
s9/IJwGkM2DLMJRZS3TFEQFDURrfq185+xO//TqEdyApY7nlkmpensuuxRA+YpAN
xEcUfwAG2tslvvOl6Phgc3YNjcc7bs0PMHLvQAT1E/5/ATWjht6N2abM7fewEKjS
zZYTNjSX4x3YVN5APpIH9glYk8DDqixsggJCbYc9W4Vo0Rd1/0hqFedtghUfKZyL
gJ+9AndyNcZpz4n08cNcCOs2tFmgsaqCsD7RFlkaG4B9rpiCDp70U0DPPq1o3CIR
iSFGb+UsDXDVqoaVaukCoU7LcxrFWBM4R+uRXtcSKiigtJrbvJ22Xcl1PKK+js6c
/yHdS/X3spmi/2/WfFrKrTKNvbnalCmw9dvxg6jFfQTCszGFRbHLm5dNf2MF/n2c
Rb92b9/5OCvl5IncRcBq9b52CxqPSb64/Eas/ZrbQvdUVFVsh6EptgM7JjUHNI3H
IaGCD7CMSZb+ckpYnDhKCgo+KcETnFy2Oy+AhEo9QDTMG+j8yMdVmEZ4iLJmDT5H
yt7ipKf+sFSrYdSzzv1DLyxoYjNhrxTTfUkrnU+rZsH4YyclMcjZETN9caoaQLW3
5szhcrNFNA2GPIuJUpTsZd7ijJE5VeyQgZAdY+Kon+LbGNGJ0fvymtsbIUOp62qu
Nd1sxLPhfxug2jrqWgjHrkRisM+M1CFo2XtpXVc/YPlMpE7EuZTX0qR7lseu/wNu
cDoMS9agA3nNYlDqT0MsPcvnQU1r8+0NqQPDUjZDXxnI+XA8Q5sQqKOCMUYlG7B2
HEFTPC04MqnIvs2BCfHfW+9qJCiAaWNghxXCofqTf/TGVmqsIIRiEPuofuAkaO9L
u24L0Iwb/Cha+wdA7iq4WRJSUEb4fR4E73OE19BXRTLk7FaG+/kFr6V9hVhKnYvm
IaxkzkZaqFYKjwW365T5rzWomM4+24BgIpJGebFTJF01Nske1pX/3iE6nm9Ccr8A
n3qK/2HwUVuuI9TRbOE3mKs1YO/6FH0usDqJyQQTOsSUkO0YAyllZhpy2rFsy3Xg
oBJ8ET/rH4JUN1dV/KIQ1MH9OqecDGqM4CRskAndJNg0F6q7P5F/4iQ13PQkeOXa
iEpRK8CWvP6WQLD8Vdr50Clw73Z/RfgWWvIijkN/QuTRNZnQ7VJ1p4F8PqF/Vz7v
Lc5mA69QSw2BEeUmZeIdbbG0mdz7R5s/YuUSt/So4vioHqKpT8NXyAp8Ya4+Muwt
E/D1pnvnZsKGq+OyUCe3Tlp3munS6e897RLKhf7oxMyHvHS9oM4Dhl5h0vyqNkNX
6NvbB7w6HpizFmz2MrRC3/BvTkcZuzzsT++Fcp8dSfWHf5ZpUVswlPSY3d4i05mA
/BMlu61JiceX4RUYLa8oaowdOp8MbxMxVXxnDH0CoIRWppVPlZuTN8DuSjbrB+5g
QGFEUuDTPbFCHALYgXnRjVclWsGVUa06vP9coq6f7U60bxnnN3+MpEzq0LdUXaQe
0uYZZ4elMM2mSq6JRwG1qAhcZP9JQgrOrkudEQP0YhoGF+B4QcgCSgaw/Od5Dke5
CjSmr/K0riHmctP46i2XASUGEmtBkIF7Y6/1VPyHqlipsnnYoSmlRv4BEZA3JstV
eejt8/TdKrvD3qmWO+DDBmr7CrRGhuNp/IrkO70ipsUTH9WQSLwpzknNY/e3Pt1s
dFWRyjED66xGfGaeNNTfelPdHj7Me8y6pH52wOulPMPd91q0Z4aem5ZM+2cMjjtO
795krm1/qDzuuMtE9EJTmFRpk4iv8WYZPzlwd1ibjOIkia11m+CoP0o3Nk7IKteZ
aPAEr7DzAQEmqT6PdD9YHSSvq45FyLckR6byEDqyHaKbpcQNJDF+8myuTFBR66wc
wpFHeXQjRXejTaG2D9muul0w2WGJvplZghl2DzCry90PLRy6be2H+oVLchW8JAUD
GcHzcfxHi2bE993s1OOV2KGDYpAdzK74kDkrpI/7zqoBwt9alBQ2d91sknhKIuop
2v7CBTmLvYtO3fEKk5/x9OAQnNE+BcIp30V8OiaxIyAz+sHrH9M+kltOLg/j3yZe
KOjQ8bunXLnlVYm144/itpW6Hk1YHGLVgYjQp6xQceomfZFqKQghIeGkH4uoDwW4
k11RjgC6Mz7pj43Si4dxnKP30ICi48jHU5PWi4xK3eyNHzyRSBJPKm05oUw4mJyX
voj9ga3JLjkpsu+qOKruOeaDRLuUWkYXckPXYvry4YwZjfFh4ke3nVGQ5b35p41y
iY7A7bC9LaHlXXZqtpmUzoaF8j2+UKAhpRhICCWDGH/J9CjCba21Q5e/5AWhDXs1
b31sDqn80HRRzax8mPjriwPysr4rjs7rCDizkGyBTEp3SI25/3lQlOmBHzsHJHbA
UKeYtvDlL2bfmLWKxqCokW5mkTrpzSHGSpDJ0FKSUg6fStHEyHpCXRfWaoT1InPM
DgdZzvbksIL5sjTb3iIO6U7+kdqrS0ekEeP5+bJbwezEnbQOOuouSUfNbNAnWEM4
IjkbmcPoUhWpHXPIqTV12TeAOr6xZ9mlDyXna7urcFt09z++VpD87pPsI0H8nMAF
Yntt5RVkzTXBBCeZUQqIxzqrbzjODr6dyZ9yM0rcKBDUFCMmCeud8xsh9PNL1dF0
/WiaOA06sLFzflHPsFgbMLcqyf2AY1faGWd3cjTEhmSS8maYVlRBSMf4scET4QP2
1JmG+/oIAaitDGWjpVp/I42E8ibSu72q666TKzDfcrFkT/A5Kj/8w8bOYZSCEBTn
qXcBU6HGqcCjSQ9hQhLdhCmgV6kcrUN14yZudjzSF12vZHfbK36Og5DAoj7mr8It
D9pwRHbjZc+koPh5kFN3hDasZW3AJHWdTmEMfjUTC3Jamc9HyQogTXVFRTuxwESz
Aa6R9ZzgFqJiXL+PS5xAD77KpQp9BKXPw91CFfzEcqLR4U/1BXCHxy4EWxYfQmm0
7EaYaBe6RokUfB4RoYyYLz8KkGbiHiQFz/lQ/XADcUcXD9AdN+fP28hdmulRnHEO
Qc8F0Gb7jgR0AfyHNdoIAeNcAuzD3D2SFM3GnXZCMAf5ILjyXdhbiL82my2V4LUe
Efuyuz2rmttii5cM8ZfKbZPZQykcaSbb4J5OIb/G/DbDnijpfux0/vxHgq7Camfs
7OyLkdUKDYntlr0fnlNfhLTk+3RieYBF8dVNRbkq8ymGLALMHs/qhzpoBqU5qJ1p
sV40Uh7blPXBQulOZMKdkR1SJDLxwPMQrKPIYmZaw4BhzdS0vdKJnIERwt5yN/vS
a+zlfYZzUg0IEZ6vx1Esg7ScJ4SXq4wRM2xDIli+xomd/8z4lUj5dgn3YnFsUgDn
PnYRSt00v1GUOD8UegN3K9b5iPYOYPdeFPXBGRReSWQiqlPHwiedM7L5UC9pej14
Lt/tB/zy7oHA87f0VnggFIYAityG+gJRuFbr4iSy0NHQzFOXq5Bs3jD+iIE+ftWI
gMBx0b4azkPDAQamqCZqeN+SbiytF2uh0P4gwUAiS8JIp0OMsihtmH/Z3wVhM6hs
3ZquHsJGnXdRkteu2jvlFTsQtQyTEX3pmdNqy8C+8JuWNmHuml78JDMXX/nINO9T
aNZhW7fbBaNA4cvFrrbQycSeM5+R+Qx0ZpQJtDW0U6/Y9Qfy6lBRu43VxvHRpQT3
DkPe1gPSnyfamjlY6yPNZwszUkLjtzhxvVMS8sjJB/mrg77j1xA42qTdgPJ2cJZI
ZMvTpJfo6Sm79y4lBju4iQdmpRsR4UxAP9oGGWAHN8lDCW8I7mac4V9IB5cQPpf2
J3t1p4LoEsOtrSKsJCZbs7NdKzsi+kURsL81i+nD7hYCZCNsjON2cz8HUwNB0Uxw
SKTiyerklDO1gNwHgnqPolCi3s4TUr8xgUAesQa+5wSX1Jm3phQZ4OwKHEVvlk41
4fqF4P/rZZzctDVMlmRCrv6h/TxG3MnOZs4U4OMNjKaQ1dad24vPT41RBaR2yN0A
+/R4MxYcVzTqVVKlS7PuAUx9rm2Z07HrwqWvsEiSAP44xYRanxxVTujdZBn0e1uU
K0Jaoctt62QLn+fb6Sf2zjJWqmoT6paimz32+WxBxSQLnoX0kcnsUfBKdkzW2El8
Q8C81ZDHe1W1/1w8tVilCjz4NGQoAhUCFPs8CkCWM1S9+weCURst+Bc75Z9qU4f8
yN81PYlcJtgDhLj2WIagtRseJTsHq5H1qkgNvudxZAh8LwuqOQcZOEGSISleAzq/
JwHw2oCLXWRIxwM/ajnaPpVSK7/QFVT4/RGP/eM5Rehw/HSnKVjpLr5BK6y3BFk2
UrOpq3T/Lz4AAd/3SMavOl4Ohn+Oo/Lm3YSwHuRS3bWBE1O72hHxJJ0zSirxwoYO
vt40uRJ5tbkEOxvAleZF2CS2U7rjS9xK8mohp6iWPuHLolw23lE7/GMDGakZOS2P
pWpC5oqx502mPb4w+K/sMcRWj92NR8xBX0YNcoODA7gdPHBq6Prf91eK98iaZKSG
BQ63bzVGzP+Ldmd6obkt+NX+vLFH/azG3Mp1BM1taI/MzPCrbRQqNtJ9SJaDrLfT
LeZFSHoG2Mxo4dhRpYJdi4VD4uhwkEA7sTrFpmngnoCDQyUM5dIDUut9k/whLG5k

`pragma protect end_protected
