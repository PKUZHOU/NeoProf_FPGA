// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
4azlZgK5XVTMjw+002TdWy6ntyn5i1vOaHrS6DQUvgRQNg47ZB4H6xEJZciIx5Kg
Vlx0tNcII5ttI6Ul1tZdCZVQZqWx8LHxPVaTaO+kySs/VIIjp9KhXerZnQOkZQRe
DxO7VG+LTzq9n09z619qxdHf2Qgx60/NiWaV7l7UqSY=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 8496 )
`pragma protect data_block
uDaNsSenLWJz6zoFZ2cYeWEf2QZIPEic7jTKrk1ANg4wv22L5Fqp/bV0gTGQcU6O
eyQw4i28R0WtaervOYtyYTzDXCYUEmiV7kyFbwS3EWZfc35S92cT0g5UoyWZcGTA
+Y5F45Ej42g1G5fumUwqOBEVkCm0oP98RAfZDtbP1H3/KxSKOC/dt7oe/kqynWi7
SkG0utkRl0k95SY38Yc/DqZ4gx8slPD8qSlRaST7kxc1/M0FnwmBCbT6TRcAuw4+
qjx4VbFEydqrdpG1MW2RcKxwwoDui9x+hklAQXS7YHxDibfoPqpPIpJtlvFKf96g
jIXXB2YfZxx4Xrxwo1NbgTQvxnciK7i3bZ1EJnLEzcUFM6KW7OoKW/QGh+HK8f+8
Sp2Zh+hYTQSEEFJNcpSAOxQd04yV6zSKSuxkcN6Hpw5p6Yh6SE4UAaV/7wTOxzJu
qS66AGwpCLfbMrFCtiwBLl9yr3rR4fs6i7okrgXLtoEemOTkBbjPNRNLuHqq4wAl
ks6kK9OUr7sSyq8to4BzmREI8HWsH89ICr7KDe/zgRrUh+KxqtklDRMWaWH6YtF4
jTeUklT4UUE1f3Ao6uFFsvM+OUwCC0UVl3RoFTfdG2+OOzVbSQp2398dmNOFPapz
r6bDgDgJBiPTmCqtL9UDWmPkjkZZyDHsyGF1T+kC3HLK+jHYbETeR0zUBsWN70ku
thKFbyzqv8UlJK3OCHRA6qYIQ6cPWXUDZZ8YA7QG1e4FYPOp7/Dvs6qwjA30f1YD
lc/NJFjK630Cxza3R1KCZLej6YxRAD06ied4axC7JF4tAS0Nj/zgkXYvAf5grD++
n+DFQast8WPeV/3JC7TsCt7F5+5MygIAyoSyc7ZYTzkXSoc4klF+1ABMwcHOcW1s
aaElIVrb1aoJ7fFbK5vN1TOXqKEb8N4ncJUzUFZ/kGjNECeI9uCGh9Kr1dqxsZx2
GN02kobi/WDDd7w/o52bx97SiSv2FY/5Q2y/mkJ2iujVczNQJTYkwT9Dy5LfFgWI
L9Wqc1KIEApzl5F66Q1IQlA7A+xDWCzZD26LnLoWiauWG2FCgMulRQ5e48rRVoGq
7jbrCQtzhM6i8+UCgREHPO9wtPUSARO2+/bXrzT1B98Oo6IdcpzdahUDvVPxemp/
pTaTlz/X3hPtF9Ve7D/8NdX9yOdUPOCSK66FMYHrKgOXLsiFGN3ascxgn/F1w0UA
yfx5ERvqMoFRNdiHpXV7pMlmjBrAPlw1OOHVZu6VKrYDspOMESQZphwWH7v8frQa
xTwRcGat2cJs3Lth899QBa4JlcPJ+AOGObecz1yq5D/gMVNell0tvTE6qVRq9680
i0GcjkiAaKvrMG37Enf14/Vzgy6OjIWZs17q8rUe16OU3XN7Cyz7IcezFmtpychd
7BK2OK4TnKpKDkICFXLEGmYDVHDFY7V6E7zygT9zhvgJipJjzJuonsTun27M4An+
Z98Y8La6f6U/awZyndKnY+r602aI2wKqCQ28by1KUiALuJ1YDRuMqTgRyDlyMjlE
kejPaBQIf9kxxGJP+MMdZ0gxWoBB0YuXIEeM9F3X+DbN3KAovjmYY9rSVp2x4WQm
Qe6ZvUlTpSF8i31ncEy0dxNWpQjfJNxXKd70gTKHDdpzUo6ARMExLj36rBepOWnC
YuWrsCvcqH7iTvhAhFCfE/aEE8LM3gtsPCsi72di7apxcAlVE4/X5rMhWTnp4W5x
3rxSahPzF0SxT05bCqusQnLBJk5X6nynZD1oims56Ddt+0fXU9TpFknWDHqLji7j
ikAmrczazkt+jhtX6ahDxDwPbmSb76Z92CB/RmJdPVpTHH74tZfYy+ERuAvkviAG
ZjyiGv2swmMzhw6nXtycjQwbo6IiOsqqLLAIXPcJYYPzxU2nFozTQvZmYr9BJLIm
Z5QzLKGMptNEQKWG1tc7UYaoIm7DiFVPjsTFxiyeK9MUrW5UgjplxRlTkQF2mAYQ
LR9EyiyT7FWgnPx8z+Xdtgc2ePxXsa3T/tjCS/B0Ke0UGZWDTTmcW5bxmiGTQ23T
AnCyhtBNK8rogbIsnk++jD8BD8BNy9Jn/z8MBLxLf/32WzebDLpFVrcBZY74Antm
PszIGKMYfWzkdzzXyD4thOe9mVLiwoBNxo7RpWkf12SzOQtPSq9UNmTuRRebbNfc
Fbru8l86Nsp+AjgDtzwdDB6eiujoVuIcYxwPRCw8UiXFb+Y4UQ141FFyR8q+9fSW
CTnKKAXw93Aw9EQaxMJzQgYzWjdIFAxyGDyUHILWy/GOqtBLmixqVj9coz6y7wu6
HuRdOhutmM+ieoEaPQJhNEQbPLUJaGyI354mefFAy9AF8hWfBgTlydm+Unjiiy7s
Z7TSsjOZGsYAh/t6wWGgn7SN4sP1tB0qFCZIjZbjYFKp21fXuH16Kq0IVWpUe3QP
HAF25k9fM55iti7u5nS0vSlqjCeY5JM6qYcMk+cWIHZjJjDDFE434HOZlX3aC8NF
kY9kr86+NWAdtn2AfoFBAPbgM3BjOhutvYD9gnpM7uQIaCmQoEG2gyHtUTy1Ty0v
nYzA0gjggsI3mSJF+MM1mxkewtitU2R9ujFNYJXwYOdlkvxq2D0ZCu+56rGoHvxa
cPGnT7/Rt93N7YXNhD5C5qmcQHuhIJRJYtSl8vcU1ZG6VuT7fC/6sMLzYvxlVNFe
sBXaxaOU5WNSzO8HCr/edyFuRF4jOlydIdCE7hKJEwvC0bVt5+GciX+aIqtIyBTV
4+jsxyeGNNFpjHQrLXx/X3mWjh9DrmKnmnzWtrJwm7cw6p9GrnwYBlrA5NLTpd9I
VSHv052xSB+Tj+wS0eQ9ii0OqaUdsugEJ72yoUTVfoDSiWIaaYsXzeZ786olwYA5
Iwefpj3lPZeE2U53wq0adk1hX6VY35uDv8l3WbJAUfuYXguBAcmKPpyiZw6AdE++
Y7kuKpHQXIJ3lQodyyUDDdvgEJJJtpA/mtilmZZnByKRayJi9eehHB4JNtVnaTs1
flHQcFw9LYfawsMTgilqgbvVmwNZC1eDkSwjAENqBtmWFkL4Bpz/18KnkXigjyol
tsyklfwJEyLT3u3j8ZqCCdr5/MbbDt8jp2GlK/3Ss83NHHvWJtzklZPjD2B+RXVN
HDK/Clngo46JjTtvgHyL0gy84dDFRMVesD3PEv2191zcQrHuajdMzhYcGeshWJpR
eLIwfUXpBtVfoveZ78r72uCW+rOKp7rEG9m8AX2dVIyq1exaNvN3ktNgEurKOI+i
5sDKcSGXloZ1D7XuoyVZhxtKxRn+Lzd7cKJmq2Fvw/Ag5J9Mi8r7S56MAEV6hkCz
m6A7SqKPv7TeJD92urwzOcEVscb09h27hvNYPbhszJ+zP3VTlJxuOlS1v6PSEAKp
2zroppxa61fSJ8ZADQPvaoeAawWwoSVmEs8zPsZ8nZaiWVItXc1b+zi74RW5Df4z
Z/ivZRo35Vpk6xbpaoT/hwDOwgGOCYfasszJlDSb2pzn1D9ilqqZCROKKpfx4Li6
v9djzKzaaNSVz7ssy/K2cBdZP+I61KDF/aVZl42AVzkWzz3nScQYDs08PgGEmW2c
S1mY5C1Q0hHaCx75n2UYM0BM+kRNyTjh3oe08x9eyJz3918HhTNxl7pa9z6tJy5f
qXRVZ8yzjpjaG5YvMBD8QdDqdcXXcl7Tsz5KM6A3va0ps36p1kNKW6pvnZjsUoxe
dtwFGtcaUkhGoHVJSe/hQ8fX7u11/pF/UPYM6aPRcKrHvrGAv29sbRWfcf+fX6P+
jwx2xPaeTtY1EE9/Djs1Gf8r3je1e5fKjUfyZO6Zp++v4vdDelAv0eSorFyA0IgU
aDzgUNGDe8jM3v0CyuBlO33Q83sIg4Qx4yWvEMexSwTGv4jf2J3I6UjJIr5XODIv
6KqgEaifD/tTctOgVN1QwmSfJ9K1wzMQLXCpgPLvqb4NaG8vl4zvGTgQNXYxmrSO
iVCDDGifYDan6RxJegacmfpdqyS6PLU9p2WtHETzpLvfOreDzK2PfYTphZEZOgqh
w9fDQrBFbvBIk6MWxXatgvijxUtoroOGCXiN9gOG8/jRNijrB7AeUpclTfq+ufqd
Qc2Xe836lwZuxXQUd68IKgK8fH1W0xdgIEiccnfF21iTqt1AX4IWUQgEsymxar4l
55Ui7YF5Jv2Db7aLIrDF9S7yLzrjV3N5aW4cVCIx66uDZO9nvZ/fxdZjMKMq0tNX
HD/fsksGDC9bfRHpSYVSlAt7J1v38PApEBzJz4bS+Dh4kHQr9ZPLWtXrnqXUUpma
VHd2Rm0Wjw0VxdegpAEzWs7gMC7CN7dOQM2HCzTbEqb0MF1bOjBH0VWRv0qprL5/
5WNZCKyzAbiQidmyX0fpwfiEuye9J50GP3pH2i4fbidnjchGcb1ww+FljlA9n55G
/ZE/xX2CkNAVmhfREe+C5iv74+vtC+1ELMggLjGOS2eAt14Ou3HjDj3wZSKLBSxB
dOJHfCOjUNlGMyvppaETaVDHiak/rk+mA6OVvxQ0oOp7zUwTdUAAvLLMRuA4oH/8
GSbYL7iYbZCueqJjPO032LtWCvr3Vy64BneP0UsNsq5sdhGS83jdW+lTB0enbtCR
z8DdpfkDfL4IAZ3wd3p8gegTrJXzQZUM0GxnVU5BgV/x1WhiYpAFY8XxuRn1AlpF
rrgzKyEuMzkUwx9485ptS1q4N//YmscN7QeOMX14kNt/ihtEjp8UXZpyI81aX2ap
5sFt7EiVtO7WEUbnpagozz1tt6zyJud1FbkxYQxSPUWMkNlvTlaDSgSBt5I834eH
RGBoSCub8Zgnt+S2Dt1jG3GSUa8aHKLK+/G01EJr/2vohjDKlgt3hogOuOZ65i9f
jCh4Zp7JuGQ2ggyvyWN6LLpy5T8IlP9SL1myfWQ2q7rXNc5oAAyjKcXey6XM8d+e
QGvzEJbX5G3urV1Z3lu9pI2JNSpE9WenyuEt7WoLxqyneZJCHJXsZJNjPqq/ru8V
DNuy4iSXiBroNZ8y7y7ZFj919wIx6zKM0w/K7UMns7uLMmETtIoQAqdNmJ5WpIYR
tcDWcGn4tS+9awGm99IAQN4Ot1W8kpMiETKXJb1SmrfS3zkd7omKv/t0a/o3r2fY
MaGlNoIQRURuFrroKXgjmlToSSMd/MuzFhPxGq6AJaf4wUh0hqKeBW8RNWl89OyM
hAUBKLBC2TxUQksW99LLLp8nchTKr6nbVCnD50UQcjMFvQBsdyABfCvducKedBfy
XdUkT2lu5sFLrJh6S0Glqj4Pt5VAszQMBxBEE5eCp5VUNFvfQHNjpjuWYA2MJ0Qd
gPxu1Iof/3nDQ//X0KHHkvAC4RieYP1zaiIlFyuypxdf4b+pvVGh/INNr0Kcr1v8
ViYKbfpLKuLGoZzlRjBhJW6lsosFBJF9OdEDcVAPESl8fJ34voDJIwagRbU+I7gW
ypskMM0KKx6kEo8RgrQib4WzxFOh5jQ2IxDBRy+TPoTQrAuUEgNovtq6+So9F4S7
YsgAdoGwRsTFDfTaKnhhbNFaKNFW40nn5+nR1iQb0TMeYaMYR086G8t/l0mW6gfK
eFoxJuvKFz+tEAPcGX5gUlUDyLveJmbkIJW/+xklBu7+q0MxOQjm5FRPu0ixvwIR
CxQubFGMB1FEtyDoeP6yNn2n/w33GUpf5itE9a6hZ69Ji8bziRQeta/1AKl4qFYU
fBTdJSPTQYPnGMHDOS5eXJTgXiQJvlwx3B1Dh9Zn1L7cQAVt2OlhdybIVNaCw3oF
oQFrJnfGWmK8KuzCIB5E6X8JGrq0ppBbXwYZIR5efBDHgWlmLBYtiKRDWNOfmeDc
RQaffYlAKN2ldjVZ+o8Cbi1sssN8qb+gsTb0M5FtM55+ZMjJpcVaDGzztGA1HyUf
1H5cOiRicFJleu1boP+07/JLwDhMDPVoYvowzA3lOrU+pZwYQpIq+IZArawPJIDk
96gWfyYa6WmiZqDrAH7Kjax85CAa2iaFDuYSjmyv3geLxRL94AWyH0QXyKT3Ghb2
ZNVL842fporhxQn5TtHZcWafTegCgLxTUZ4/QrqqF6podgu8WU1ojRAutqAlqOgm
ohdhnnqBtxtFb2mvfZZ7g131bSTM2QwMN8WI7duKf0L/YzOyVUOmFX+lV0RDcjkX
6fWv8U8IUyf+BU9gDyGwBw2xthPhl3xbXxJVRzk2sa9WoDDC8NFJ7lcnwX1+yz96
Oi3dvXLMOn2J1Alzb9Gm2JDjRDg27u75jKjXz2xay76feXRRHXqnrsKbD+pHLEC+
/Pne2J1aqmZWhTQF12fuln92ynM9BGR+HPCOxpZNxdE9yUZ+ULmYjZujb4KaFq3F
EgjqjpBJvFyYRBte9bPuYTYa/HSLV3Y65Hf9dLVFl3usVVCzlrUbhWw9nXHZ93vj
uWwMxwRLcghXMv7+y0IXgRWKIBojaHg2uIUNENd1uhvPq1zIcjjzXHugNMUydAAy
v1ntjw083Y1IxT46t5tBUBHUWnG2HA1b0z5cSBnvKeAV2Nys5jpyXoqmxMUZP4AI
VOGNbzJ30ViTjSyVEPTC5dMSB2eIlfM9baI9OY2kRayoyoQabTZtWDiM79VMpaks
OF3ySfI2osXOBqt6otw0my7szyzSjXIZd3mTeI8uL1IGHrmYIEmDcipuCuu5WoQu
+Xhafb4XtyHxrHxtJ0GWl9ht8GoSdNlcia170iXokZ4HcEtk/tJwT9aqftj/IIbR
E1iihI4S2iiJPT8xAeruWlLi9vae4tTG90Etg3AsFyh/1EXfoccmt9z2VbjuUX4q
M3+ApRNVnllPWunxmfyaH/79IVCvUbRnNp1movhuWmnIqP2J+9BK6f16+DV0GRnx
YBrOjEqdFoR/wlrec9BEqRAgvXJTGGK0I1t/meG5jOJubSJJDDJlE+BmSt65zCrv
N68KI1Quk6EV9k0WOPNuTEwut2NHvVKVc17wNzMGB9TbMHCgE8MiBV0naWYzlenM
GhdZZHklm6n+OG0HZphQ+MErfZlTQzT0UlqHvFVbfQ+84GSmODI61ndbqFQogAvH
cwpEdM9BJQqiJSosRHoEAaFVUJP7h9qbB0+7KAYbO9guECwWyzemFyTulU6VwvyE
yQIWoxi2hkUyYs/RJDx3lCH5EyWQvecJOV3FrRdF7EyEMqorgvHIH5GPqHKOQl1P
orJA4bq3dwT/qvjmNo3CKDoZ5DIiG4kjKBA64/3eH28SNYL6gi51FNgOBoICslrU
Ur92s9xD8wV47Guhz2SE7LoLFsVOgDMDTjEh5UsEUv1yrLtxZF7W3jxULcsGmx9p
OvR80GOF6px64gzkCdRlw4NBktVQ6fKmUZjyly5oeJGaCTj9lU6pyb5D1YLG7C5n
tIJSO7maSaoXflxtiKnyTVXUCNlp9i/MZCFRhSAqar2Fke9zBq4F13Bw/iHtVIXO
QRqsCdm7wi1+16RJvTdEXSmm9hOTGxTVVQeWmOXVcwOwsqoJcRUq3Dy0FgD9Nakb
K9l2UKtf8ys0iw9JxtaW+km0s3N5rudfZbbT0e0R0fcLDpFt6Bxsnfme1cgiU1Yz
IpgpKEGOQ4KraBSLI+KTpCQHv9UHtQ2CPqrnnxl0Ex04qb7Mn4cCUGtHSP8Tf2Ld
58fE+Q/QvoI7dyy6GOOwpDwZ0N/84h1sFjPnpT3WTBc9udpxIRtjE7+YuPdAeYlG
FKfi8QPH3gryvncXRFVW7oDdEA8Pc/CPyLsFTBIU9FKF25bWRY20cmyZfMrctu5c
STwmwKsy7qGYpXf86g/K8TAE6rm87rPKEENCmEWyFFjv4t8B16qEnRP3G9WlXC66
2lTRpBVRPxmcfPWGj/OHLAA38W7cCZQumrAoZ6CoPN64j6zZFLsaL904EQnBPqN2
FVz+i2a9YRcdMf5pYEoHskvep2dDSO8OjhlZAU1U4K8RBCFsN90SBJvdpVo9eA17
3/fO6nonMQV754OgD+wE4NomqQo95aHUApdfTi+ctA316pQbkXYQ2pYnXp/wuYC0
m3VWzbUWujSHVAAwjtCdWGfXVyVdfNW/FxuTHndIb11hgCsWRp5Py8R5EOfzMF7T
knQF+zWJGDbFHMbCDnrIVss4oV+1GOYoM0v2+6pl7t52D9O7tLmQR3sACOcP4ddM
vutI8D0ycENx+2QVOPnKZ73GwtYn6RJjIOEu317xA/PWx5QtxVXoG6icRgMi4LgT
D35qjvtwq/24divTxosy3tX/c87S88EbzTeLWb3sWXI3mqhFbz6Es+G8dXaGrnKL
fejR6+uJNDaH7UO00+F4veYPLyQEw5DPH9q1ntqgQqT7BCHJApeIuw0pQ5qO2xkT
X+iCxRqqp5FUU2ajMk7u3rQQ92yRZJfnyI5/5Is+eV+DCULAJpRZamDwsTB4T1n4
hBmYYMSvJFc87J1WnNYLxfCdngD8v5TvIVUp1N44+PrK5tr2Xo9NETf+Cs6CvaJB
jnVh9PZJ7Xv+2yzIUPt3A6uUIuWgG7p+iHI5tqQhMSl8lUpsbMP5elnhgQOF3TqH
3TLbHUSYcIS7thq0/MEiUKKWPGIQfTCpjJHiAY+pLO76nYEBtXhxzXvNzUkfcj5L
s9CF8yY9LXNuRzycc2EtHAcTQebtKxLIWo05sA2jLzdwctc0qKifAGNryg0EQq0z
v0ub80gc56rgbsP5qDfErqrtM1N+BNmMKN+oQ1HB+yRxxWujnKhNBn4b1N55HGyO
YfkLarWq5X1spMhFp0zDM7HTdo/CKfmCFFMWt5dNli5vMnxka7OgoeBg4HX3PSNy
2EV376kgnBbMwZx8Xr3a3t2g4F1bmKE7RuI7zlZLIXcbbWJJx/QLQFHIQ+71wsP3
d8Hp/97s3D7pqcBTBtUEhPlWRwjXefBEnSOyYtWAOSjQoEcwoYSZxMchCHwf+b3e
sGBh8Rz01o+pj4IJhseMdXqeYgOJy6P/m/dyIOfNnSKC9twtNXI0NP6VMWYYB5fi
thyzx9zrzM5bdDjt1bNZkqIpdRGcJIq/fK01YYnGZ27OkMDi9b5i2eRzNpeqViPR
pjUsKC7MjNatTQ9Fd10ZKemfvKJuPsxx2oMOZE9fKMG3eaK7vTRjBDu7aOOs3Die
lHZ8rNvvivph3Aja5oQG/7FZnaVLlakWGWcOuV78NT74y6jtiq1iV5CqDqH8wQ2B
nVzc+9gzyqEdNf/Eg/KVykgtpViJrQfsQje78d1uplj4xH8RgYyZwKZVpa9fvPrV
Mc0rHhMHmHPUlvYWB6ua6MMecLi3cbtgPVnzVfUZlKU+j7D3R3CfA/sS9Bt5NcFO
ITSrNTFAraEFuWd5uCef/Zgii+c6HySuIXV+kBkYntq2pVjNhPTi9YBZsH72qQWA
6FbHIQZGISe7LFkytzfmnvrbLxMlN+7SoOcpvNkbo4IBYQckqVDwVxA9iTDdWPY1
32eZO0BT+B5BXXUQwWhyglzmiceTTfFjdJTB2xfouoAw8j8Um/NjoDC2LQKonWjE
sWUib1Wbk4bwKHAiTzC3YRDHFS5iiVgbCyTfTvxbwH4RQNNTQwiSqVnqzUGOe6Lk
boCt1vCPO972zVDuR/U5T36EzMWRu0ks4NLF2a847XnYEDPpySSVmSpuVvhLrcDf
s4XtNLUKkca5/eCtBzKMbOEh8bdDHEVgWbjd9Ah3e5SMId9WrhVLuMTM78Z+fpgd
dcrSMOgXirt9633Qykdw575yNwuTdZ15XXz8HwbqW+P12yiMQ85MY/+lZm9pTseW
a1P9aOr9BkzYUXiKfzeVtMWnQCJpZseJ1TUP/9xP8BFc6WIHv5PCCeSPSrKkNbq7
9/H/qMUEVao040T6UFZ2RUDp0Oktp0Gzqqhv+DSGnOtBlfjgo6wGLGVRNCMOR+dS
EobbJ3XmunFYxXDdXSC54lUqUWHJ4QRHsEoRd8+ES5IgbcHBXXmmwm7O/ZQiy/NK
XNUACYG5pIDb3syHTP9G0Q+zfZtIp9/tvM214d6nTDLmNUrnzyHL1UyPxQsLoKBH
rA6hfBWDowvwZK35KZI1t/x2YmccljU3Lqdzau3heKcC8K/aqzGVukfg7hHNzZ+a
oek/XMH6e8MhT/PSsfsLxBu4KltTBAT5bamz8xFTj865KSF4Q+79rY5MNeCcaJ3S
pmYIiV8fkmHGI9+imC4ZtgqaSFGzTHaHdlODCRofb80sK2HbcVV4qyPnYfaZT0VU
EprrzaDD/YtDkQ5+0Yd+v1VjsAuv3y+HLWUH7IWaU44OsGrrv5aTHHom9/wpM5ba
r0gELK9V1Evp9ofFHUAwAlxhCDZ82M5ms/5wqWvW+yHe4rSXH83mQz8PAbPykRkV
4d19Q4HzbrfAzaw/0VJoUECOdbZa0Xc5EIKQ/ily9x2UthfxfGArKeElTSEbsbYk
M+9Uav8eoYyqZth8yy7JOZitcnE6XW7dYZlS2cUVez4EW3IdOWcBhrxMyefJtrT0
pQ4EawFdmrFpc8xNPsmLw3lEgPVRX25OVHXYAwB4KqPCxwLWtwoT5y6+nNOEQWqD
mceXtUty9JZNFo0r+pwN3ZC0tZkOcPiKDBQNL4ggbKwUTtgfn8bwhm1TaQnSDHoH
+3FxkO52+a0gb2JdXwQHVyDgqItnmi15UY5+0Gp+a92/diB4hPE/GAXX7fPW2ILZ
gpcwI3dGbm8DHrx40lqYiwXVd3u/FnNjozT9Wo027eRM232WHDYQGG+GNfigdWaD
emdFGfxwR/CSEnaH9CRZXKHxp/pMfUjvYqDHaLm+jRkkdvjwOyBdvBvc2FcX08Fg
hlDqzX404mGOq/bryr4SA6KqHAmA1klC6iNEdKwIn/5QJuu1sUxc7bUluKdbUhXi
+JZtRBfLpW1ye/Brhy5u80elsatVLUqNXQV7UXNxl0GtG851XgDqrQ9IaJw5nUHA
0gil+TFtI47MwxbrCjTgjIgJ2iB1CMU+HOmbvajuNIq7IDnzqnyCS/X9K6eU7Ww9
TDeRNyytJJLx+A+5k8tGljXDynyJNHUebjWEFnE/2TmwiL62je5gPKPfHNQzg0tg
61sMEgggEJVZzSfxkpuDcSpY74n314Klw5DPDXq0gvdSsyV3xyiVUHuJJDeaNHXk
ToRK8eFayaOVRQq9+zbmMm8f6siLWcy1GbGRGc8Qa26eG8sUhvOL14TYAXDUdVUR
ruHt1/2SnEKfAsqzJWVDs2O5/+4j10v1pFd4XetODpupZlvl4z/7C3+Ru2eQDhyF
zLoKcQ1RcBvUsUAcv9TVzLqy5gIrbrBaPASl+GAUDJOFuyEu+lgkExpYf7AINKyn
QW0WFNtvpt4O+L874aMwGpyp+aDwBTZSsORo6vZZarh4S5FHEmuzHLbJ1t6q7iTg

`pragma protect end_protected
