// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
fN0uS/QuUZKoe1k4bqUL7H2lVN7P+eYNYe68YgqPBMPyD1n38knnM1o7Qyqy2Pt+YAhWMLv5pjcl
AtwHC/aeNvjsOiLUimwAw0sJy1z6brEJebEfREJrJ/hKI65AGVlcjwGqMVUqusGbwUZesiECG832
DyxP6jkjH0IFMS2Gv1ag2UHnrFh1tRhmrLQL5U5HcNPlg2VFeIICE1P0FD9TZqpKZQ3cVRPP8OkU
gHgGj737UtP2+x3REyO8nilceaQ0nJ7hTP2xGphaL/9L21OCkqR8wXec5FtB8RHeXCQhaUa4jWkV
xkLNuAT948jjO1B/MDXzS6FG9rbPcnd9ZSHxuA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 57664)
OOzMDMmDt4EAr7XzrUc/MzC070Uj9hFLSECX3YQx8uEi+c+dIMOO4nQLv+gWwqAeifhtnTkqeYjY
wHMH+WtpLYqpGb9Duqw3EK21bsBWxFlcHzeNBL/RvkiQ5XVBFAf9QDcfTYqxTeaGJCC5f+ux/Ftm
hs0g+Vy6mKM/xlHQ2mTn44VznJ0d9dr0ModM+G5qGLYtlczkIvT5Noq0ybL9ywXJ8b9RDFnLzb2i
XfjdbgxNTWTwrry0W3EwGrctlS5LvUsR46J+KAEnXOvUuf91iqBzP4coPpsta3uexSLB4m7EFPAs
JTp900WuvLH3234tS8kmZfQDKrUEwNheLAPFM8L8eeC3917Br+TSKaLfr5vpwhYZrm5a2h9CfFn9
ozTCHNwN3cBz+jK42IU4n4jsP/ni/tTvcO4DeXazJ4F26iEFPw1BrmY5ck+HM1YBqhN2UZB9TNM0
07x8nrj9Qt45jSubzPfD5/fnKM4xrTgrLFB0TknIqZpFjc4vxYv+6D1D741ElD/aOKhndcGR42m3
a0bk8FIQnr/Mg2ea1+bc/gisy0dPGOXmIQa5BKnNDBNxVG2c0ol5sZ22E1H9DYpHuU7HZ767Zluy
3F5nN20vX6F37NjF6i9YnJgY24JPo46BA9lSin0kN+wHPjmxobbVlVT8vqVHI6Pq89WhD+bAeORR
HRGZqwak04tBL2kTwqu8HL4UX73fhbM+ikrYITwQElfEJ37jsWBCgovvXFSvzYf03XKX2yvfolYd
XIBGg381CyE7DphpSe6y9PAA3IuSOlBmI14s+xq7Vme/11yf5alH26KkITKARD+YtVj05p214xdV
jzGJi79qkvnw7L+buS7pnT/5hHpOHsDrC/bPBYlBjyxJ2ko2qDON/ClpPslh8XAanE2+W6jrMiYJ
4h6XWFjovTn4bCkjfdTY52VeBkvyiEMzdkkfb0RMuAIFsN5FTI1nBXnLVsEbuxGJAol/df9XUNfH
PffeoOIb1mWYNpxBY3GXObdqB0Sz2ofMdSC1UcwclH+uuBPXLNtlKXFPuiPF1ps/ynaHVAbMzVEi
JAj/Ks1QceuVml0dwuATI0zKlk29P9voyuk4jxc9TWTshbBJTdIYy0iRyEAdkjiXWhJIseIUAy4J
30XBjnQ2ZiRlB870ZasqwRshz+DYFumCyeT84EQjxY/3SBdtqSnT+tFErvS1EHoGcM3Vys6pjPij
DtyhapQZwoEXJszOKlwCmlmPy1Ack0VPM/b4twosWLTPiVvAIfwJ2ziY9eL7V/lRiHHfXCqe/9Wb
d/ghSVyKWkTVGFJhs+0NMdcg3PacvAnVv8liL6+wO+s2ZuAVFoLC8gg8x/yXw2MfAO99iRDE13bg
GBXZrF8OX5H2CUB9lTnvsGN6jnGlufNJy7kwUeD4hHlkai3ZWNQ4O8Q5qiegFGjVRGzv7J12iBpm
UQASuX+WucKvMwHoSMiCqzjEJ/tGtZZPoLiFvX4P/5ad2+TIw4YxVccOTNIgKEAhxRC9RSGv/Pli
FC9qlt6iaRutYl49mLzbcB2sCA128XMSrvphLzZrFbaMZWqGAISvSflZHuZQWRQWqE9CnqliMVzM
qFLv6mOhvM+gwMf7ntSOF6u/d4znyvrd9YsJ+9z7k4Z/QiTVFq24uwFA06A/3CjMP4Tt+w+mE5WG
g9Mv7VmUcxnTPYJuJ3EkD3VA8CRIPaugx3aTIIpeXLNln0PDJQpy0cLP8w/k9/6t1QC64CdPzFiW
5jvL9jZpKGAej4ynUeaYRllmPKl3RkDWeevClOHvQ18+R1P7vwQYN8WQvT86BxFTNykRq02lSMDp
1Fmw/F/bB1TR+BYI/nOVqJ/UhUo9dFWUUAzT8TwbpsHbKzqv7naeGIAm27ta66MpVyCtkbWcCDEr
6SdieZ4kltQQUWJ82oz3k1ngkTVgisTdHN63K/h9vF+HfVjSDwUVry06yBcCyMfaKlmn3XgEuggq
ImkPlrL4sUWiSRWMz/ouS24CjqT83QBOHDac3zl0SFSmO/Fa2YkiqbalC/G5j5x7H3T1hPRR2A9v
V2ZJ3Fvt1pyKIaJo9dBYgd7EvSXMjs2ANelXbBgsoFjcuEiOLFDkVuiBEEnUbO2NBp/apKvlIVUJ
f/3/+X5TR0j5u01/egV+rsEc2XKoBlPzoTw75i7F4wdRmtMuh5B0qURqU+269r6GSU3QxPKPbr2u
3aOjCtH9NizJ513G6UnzLcvfi08l+2t/nM8OPiPqfdjm1VhG+TDSZ12DNbDwpmXYsgob5il5E9je
HUaRZBa9LFUwwvQu10HZYNTe4hBeXagSa1Q9p6q03Q2uRgtp5/60LPnCY5pLYo9sLss4qiluC7us
kuljqoSskZOaugpkVDtUldGlwuBOo1CHBm7zz5tXlPYYVVQTfe77TlEdG6BlsWUGRnYYhyctpgrh
3kDh7+srZRDAeEYGdd1IU+5vExFTd6AIsbFsa3CM7lUI80pTd6Hak6pNDzDB94Ba8b01+EzfaZN4
eQMD4dd3mB+k4vFECgvdDKCW0F5qgttPK/V4GG8naNNEZEWxSjDNv0tvEJPTMXMzdWy/SVZCuKZD
Xj/weQ6cvnhbz5raZ16HgpN0CpnfgDbvSpQjc/2bNMWd84xctxwQwPKwNavYZZPlD8X259pqJPTQ
rsN3lcoIkdieheH40hVicV8ReZ1w4FSkXNgEdR4yuWcGsYIJ6WTbDKczczjIviPOFOcHvUb87uga
Nx3FqcyZvFfz4YCz16Amkb0oNRFXd5uqbjwtYya1o3ZQhigNSWkmFZEoc5tQ+BSve7salMs/8FD1
5OESmY0B5UUqj3JzX0ARPhY4Qb4PExgxCgr640QcdEiKK373LP/DOCC5XjVzPiCrHoJCQhe4IcsC
WeEZzCEmSVVRpdMRMz45n8UbNs4/XLg41L7p0u76TpTr+vkmtN4vuHYQepKkR7NKzKQsWqyx226O
u2TldayMi/9cYtGLsGO/aj8HaF9rJ3zqO/kcCeHa6XgYxhMUZBSEfDal+IhwP7gHUyay+4jgwAzC
xOAdEunGh8EjKjSlDKIaiGAMjeH1kfPNFeznJvGcIdftMR99hH+CLo8ISaWggRzT/dXVUGkEjCC7
+V7S8n05KhbajmGno7etrAI0RsRTWQrQkVR2rcxF1Gdpp7/nlUxsu0OXEUtMvtcPnktMai4V7CkL
TcJv/KeAVQ+rebY3TBeiF3KTRhzze8b2OFl19ZW+HQQ3q4ehd46TwZJZfW5LaQ8RjOWiCoI97l4A
JeIFKB6xm2UAb2EoTlg7ukYOmT/P+AlMOvCdXedkUEOsd1Dm8O8kZnzw/U2p3v2Wnt3wJFQQm/v4
Sg9YQttVCDZdqtlRtdRC0YIgcq9mGYAbUsXch6ZISG7azpJepVTA8sE9o3CPj5cy4J/vIuk4RPWA
fvYivWUwUrXvPHL3+OJVaCF8gUgkvGirEiWR6LN0jN8SWNhifJwR2CACe+ow/BLuXlODSRsOHwmW
YfT9ZtINpBQj/tRTvA9KfZlfbGf9Rp121bkcwLmAmWs04Gv4QohjkooLN4lA580KdQ/9ozNXja5M
Ocda2ipXYb2RuWliKm5ZAejcPgiFyuz88eLxhA7r71p8kuawtgS7Dbx8paHsLRPHypSf3Z3t5x/s
PUCgbNhFWWATceH0NYWZtnuP93ZzppVIzIT5QdqmpbFIkqPm0YTkPfKGUkRKgpm9Xkxv/fsd9tNX
f61EBGSMaxOmPkMDIRTihrwi97b2yqQJ9PZbOagVEzYDenAxlaFvMNjcgL+wOmnxbMCie/gdJ5zB
eRDcp3CinBc1M8gk+JelM3FlYdg7Cux2rkEJiKh+aMyjSSE5nRMpUk/YYdRT5q2lrUSEc0r03pvj
GicFaC3pFJlWFZLZbIvsIlHKrlOKhh00S4cTGX/AFdqoozPBPrgAD2pFXEhDNHN3kS2GDrp+qe6q
ZzYgk9ZAwi0BxyoPIASmswTUAFHBDTPDxLxooUJAtFViw62CCBWf2GRs1j8gU2x1CSQgJmaRE2Jh
td3dBJ3WluIWTn1wqPZAolA1XWh6nwQHw8HrRAQqiNDET69+0PVNJiO3b9nzuxVbW892XmqWeE6Z
RdjIcG0wVbj1hnJslyre+edRoTkRaNVTfMzlxM2Yi9zxYiGaGKMOtih4jcsqcO1qWaL5SKUnwhvj
VTKO5IsCVpmnRlmRRW6HHmsJzOd9943+25xZ+gPEOM3ML7G3J6S1FTyFYNJX+Scuz1qOmstuDPX7
AwsyikuQV10EaEFWkLITwL7OhACoGIuMlklfu7R0Nu9nURIFtiLqfdJ+myZqmmpKTTQ4+RyHasKM
8deKE9tJgD4WU8ryf2u7mar92mo/0lCzytklKgha9moeVexFs1KkAZk+YI2uTO5o1QraN+HW3awj
1Pn7iVoQDjPdXbN9gZgS7nke52UhR1VZqLix2FTrFDGDnQ+EsZysxnhLeDRIyqc8oVJbCS1dtHcp
SyjvPx7rLy9phsQYbgxOL8IdTwqE+cH6lTFvE5nSb//xGNGkQUd7I1EYvXMH45FiskroNyqs66tH
RdYPMhE10fUBwdIZueGwkfP2I0zsw/mU7Z5vI9KWIyl04K6Y1kk1CRU20Ge5oVThWMfE9uVMpqr1
5ez0lLALfZgl5+XZUfgE6qZmfHIuQB08eCioV+kZ7Qh5VsXelaxZDze4jdSPRYxedyCi+Gfu7H3d
iFUY+9PVqWv5dBPRh8NMpxHQA0dhwUiBhLIqM4aRkZ+Sra2B76KGOUznRm5DCiyX4zxflIjARRoP
cASGMd2bNL3tyI5W/GVoHfnDa+BYjqQ87+GPBSjT78G6SxI5pWkVnW+1PxGdLKw71rZc/jE4oEO3
pWPqAurpO3bPotpHPmZFAPOJAPWBvl0yxOojuJ4EiIS2Zv6ulZAc4EdvWaqAtxT6VZsnBhGvtWJt
uo+uNeuXP87qWE9tbA9h/7YoUrvuZRDDSLlqAJ652qdtaef1tyLbl0ufhPqf70ysQY3ddHzzkNUo
AvwNlQo8JtDs4Uljk39fmZj85yAnTKMWhhzZVMORsp+aZvb8W/Vy36j727lFgCvm0/HRQ+oB0n/r
wPgrTvnbqWEmt5OIy/fkm0fnV+yplqyMywfM6brhR+R7yQP6b8AqE4Z+VjslYFhB/4/umYswJ82C
tYpLXb+eN1szUgz1JxzqVLK3KWfXaoCHB48ta1V/eFmHFgcsl32sKEQmtACyZb3w1W1cc+YyY/X2
0Xx4ntqDm8pImBOxPFsOcVsG7Z5chVrP8alOxfvpZohTtmL/QCAzRuncooTY/QNllKB99ZUix5ma
nenznySBP3nu5eKlB8LpBqvjTQ5eghcdP0b/tMhwecKj59WHu2emsaKzXOQi55eU6HYQcB2Liz1K
T6gJFC3o5ORWq9BPN86KhUvP1g5qseThS9xSJsMi32onAq06afzwyjMMuoHxf5Mq+KGArTTCFYkA
15e319U5fwsxGUjC9UlTdhgoff/Z6JOMYlyYM4YyCy92jg8yk+DLnwHKLCcJZp9gbES1H5+Vgwsz
mGCeqxt11JXhM2d/DdYnmqyp/8f24Xo7UTx13pfmbUPyPAC75fMFFHs5idQpue/iJVlo6wffDCII
6xg9FKCR2j9omcOphAS6IjeZdCaPu1Xa/DBoO46uszMUblCpOT7yM0Cio9+WzFDTLzLbnRlLrSVL
kVV//tnuCbMDTWbLesSYG1w0YNUe5B+g/vi+eaDT+Y1rMhBsCmCxSeLkqZvkkJcFFPwkkBmGnSl0
qM4G4tjj3cINMJJBH0U+2xoLuRyYFSGJh55GqkuMpOEXH8IGyFyVkMZ+I+T0QqGGRfLNPb8tz89y
s+JzZ26Aw+4dHOiH754YSMmm0j7NfvyNEnzN1e5MYRiDDDDuyzXn0e3496G3Ko7FJM+reUGTbtlQ
iRyPSGkJe7aeP9wKPFk90i4Br1Us4jBytQ2kWmpc3c6vGKluL7p0O1YguWK1n7WXcN2SRgKom/k8
cK9c1njsDs3SbU4ULLPIcUIB+/sXGAHzSwTgIW8xgrh3MkQDI/NZZWtncE9EnBWmuLWf2xcqvLtQ
KaLymYNnkUKz1yFJgYmVNQQlro5CanuBwgmynLJAs7oyWMhI8uBaE1asOKdg51PlxWXjOtj26o3/
OVZl0yQ2BASkk3LJZKzFVA7GSA80RQKNSbXNRwauvRKmUK8Gr9k222h3mTmRQXPUVzeVmoWiJ5Sf
tSCuMhJRYtIp5GrAF3yokuOXkKCRS4LethfvfXC8EdZdDhvf6JAXfYad/sPCAGgjMSDmt5QHhp0e
WEZjwR6Nq7ZxyXLQTt+ZDg0fHta5/T9PjiihZMCGZkhn1J2tkJEMNjdXSNOqLfaaQXRzLgLCXH1X
RTzghnQzjB6Wv7jBzawEe5xnlrh8Tex7vtq14c28xNl4XjTKPZy9Tb4CUxqArKPx+o/AxXVZ60BB
2yi6lLpeS5F9ernPaBe5LqPzwMTzSTl/LkwuDgwgmlZODMcEfeUN0/hb7qWefSCBqiYCoSR4x/Ma
chtd9l9podOxLCsu/0o3NpD/1n4Ro7w0kH9+qSexvSz/DCudGtng/5jlOHnjYhu1kVQBO6zn2Kz3
/HxwEDL1x0UwVVrNjVEQO8WflDWwOfJ/NfI9QkG2xHnb1aB+4kFL6AhBgmR3A/sts6VN5da8b5fP
GxRgzmjJD9Q6cBc7irPzyjnnWY5pAPwpqfkfRF5vDeClOVqumTFi1mJu+dS7eamrfKJBZR77W4td
fzitoUtXP04sGrbGklb4Q6mNP+ywvJsAHsTlAhJG6mr/pPgUDvLn3iIx6lBJkCl4mNuUxtr2HXnx
wJGhZU5CEQ3rTuoLVapQH0WzY/fxtVN1CxaaJnVe2xn2mqeRZrpHtcI8eI4YdTmpqIedwfp608uv
YtUZhcyTW0oo4nbPjO4Xyi4/F6Rljg9r1Xo+jIsk0BXiw+ggtiBumq+6jXeOX6AEy/Iqi67CNVNv
M11ZxX7r/olLsaawWLyr1FDjeztJjk6u54dZXBfEee/VGAd9bmfPvtxhNBNBvokMDN43NxeGsRpg
araU8L7liJJcTXqwHSETjhIrmIjcwk1DMv9dWbgw7oFT35k4PNgTYvW9FYqJmqfRd9BB7DzQbH/N
6/wPjxMd5R82GLvgh8CWE8S3VfKETaIA+cAyTRp20CrIx+77IvbQ2kU4e5A86hV0JKoeDp5QfmQW
TYslQLG8/pOlc/bkVmzKXyzokIoL8+kQvjfOLYL3IEZrK4yczIG5f7VIX0At54/xDRY7EAl2LZcj
iOityIw/Xcn3oCXTRoENIaC98V0dIVTc0kBaYlu5G3Z0eDI8RJGB7gFjhaoFmKpVV8y0JL+PL37k
irQBtQE17L4YvuW/sIXiZUpTME4vMQHnU0Je+oFHWhcb5LKf6RWreotOu2frQH009txlPBKqAPsI
MvwF3rkGXxVPQFTs8klMvxoNCmYLqHOA8gHNeIIcVlpgOKoN51JOw8BQXJ8xjwVS9BVpVgqIGZWT
03gwf/+GoNgv/qDsNR48q7X9FGYxL1UIZgcy+r9TCzicHOURi2K1/QkGl3JG7q4sluyTD3WQ43rQ
U8h7nV4eNo68Rn+dymWIJtuf+JRN/M7tBW82rs8bDJOY17po0Ie0S//vl33N7z6T6VvV4o56cPKS
+dV8E//XjmiUKZ35QqcBwkdukRrT7Ru8khWOVU3RR3vVruYfzLg26ISkRZcqUC9+Lqei7JI4bSDz
Qh6V1GNhFr3MnBJzjrRlVZsHGGe+nmNK1EgRy0TrQVdbi1x2XFQBzhpjghM9GH6ejnCKc2It1mVW
kef1uc+UlFLvOdYhPHQEYL6j0/6+C7mrMbP3B1fa+90IxIQkNS6ybuxlGsHNqbpHcUNQ95QjGy1j
ynyTkrr3zpUwf2zcP+IPHDhN7D7QMtQigHs+Sehf9OU2bB2GkXOyxc5hMpUH5tbg8/Df+IjE97+c
4/yl2P6jEqh4C1buFcfW/WNFdrg9bw9kF4ifKxfBLLcwwvxvtxh3nYIrMGPhEo3Dl+WYvnBMP9/X
L+/lSYXXHTOJmkdHNRLz7W4J8quB/Q+uuEt3WmWPQcyYwCGBfgjdc0FKrXHaNXMpJxnHnek4OFbS
Oo4KfwpAV0tNL4Y/Q5dF4Y33bKM0K5ENZg3FhFCNQ9pSdi5V59BLeTmyPXt+UiRg2Opct6LmFk0M
la6DpqjsYV3zl99qWcvqJTYawMd6N/cXDFSHVbdjyaRYvgeGvP/LqRwLR4R2IIJ+q0ro0GKKmRWr
93qWymV+PAZraZKkVphyzd+RkueOkmiLDh4hWIdAnBdoM3uVxubCYZvD+HbHBcdHyZRhxWdmZhN3
KopnI3V9rY9NdnbzQ+AOptw5ITSU+1p8l5ywKKKPyIiMvJU136oSxhT9XPHm9+09mY7LkvMWBiaj
VqvwJ88H2pRjpGn5zFMKmiDQLlKFQf1V1aRDXJkE9wsfiqZJ8iB6WLdF790JBovFLbSGs60P2WAy
ZZ8iP9SKL4GEc8cORlsbmGCDpHRRDY7z3mUUiozQ3JCpSWMiJEREXQt8wk1znzbbG5N4ess9WHsv
6OM/DWTcIJ0QIBNByUWzwc82jhlFCpN1CkwWbxYZSLBBFybcasb5o4UdOJZd4IvLayiTxS7eP8qy
grYIih4VLKhmzvNcNPXfUu5+JFJ6tj35ltoUq6NPtIQBpAYHOfnrgBvkT6XEWNfm6DnmPFWdhX+w
yW6J4O1GV8KROOyrh13cd44LVyZMsBWiUYsUONMgMUe8P3kUWhzFZEuRJd+MTq4zLSQYRXSrDvMP
oiZymhopj+w4qJTcSr39LlD8M0M3jThP/xpRiKXLCev7F/yWzB4B5XG+wvzOo0Md8XKDLSTyyqbg
8NqPL8WALMoHnwuzCRDkbMG4KGAuNZ9VEGUd/rOw4hFRnu3eEwG/Tk3yuyekUY6eF/PKH/Zek35+
mHV1KkrnJ9pgxJYknIH7ndEYOtwDx1MdA763nBzV6YCUIcZFenF235cHqLJ7Hw7QPMp3BBjxw+IK
x2nTm9vcKIR06/ygr089V/0amhjL2PEHgEYYSKSk/w6R3GCijtbKEDab0EklvwtWvEu/Lu9eRYzY
vC0xi9mahyRY8/EUr0GSlB4aUH1j2Dp81oBB1FYRYoIQF2ELNLjeJaz6p8BWyf3GGPSJ+6S1CdMo
XJ8JpA3br/cU26WEwgMH+1I0vQAfFfsl3xbW0MWRsRkW/Wie/6+tT56VhpeiSKCONkrrXiX4alc+
RS26HC5Ig/FVgBpF74ejTElFrt5glzC/W2jE9D+uQEpEVhltkCOd0wmBzM70fuvCZa/RpxAzB9Dx
QBSubedi2oNvsanSVYtbkpLtL7C5OGY0ji6EIGP4RstBzlThovso2jFvcdbY6JLe56dvqTCNepd9
a6l2mr3OjNeUTnMa2NJz1626AIFJSQd8RPqPTfNMC2guC1vXC0kUWn211DN3cDoDkfWnwYSFKU9G
UTLHfCXvK6ynAK7xw78IoAaQX9b/CnSCR766zbqDC0hTZk1SOCXsG7RpR1Uc6QqSAGmqML3PDuZD
k7G3gisHn0tV+YdKSp5W0hRaS8e5N+V9i+AXI/QKVYmMkfnJGUVeaceoyJq9jGRNwtOvOXAKfQmF
ERkExPmDqTD8Odzfi13GEdNg19l0O0H7ajOHxT4u4Xf76hQXHVLhelBOTaCgur1PXcXQzo7GsU/j
ufNsjJiaMsNsr1wRLDuRAVMFSq+5BdglN5Nf/1fpt+Hrr+SGATsKwnVUYHPVegVooMLXMgNJmEOI
B56P69SkES/A20t2xGggxIv12Y9s39bMudUX45OrR92v9/v2VgQBlN5hg1yDF/2JPAqpV1KevcYA
Es5WC1qIEv9Yk9GrPPGon62oX8Hs0ZZO7pgao5O4bGuJK8jwS4ERZPbaPk4iFMauwXfyCOOGjmPV
XhkFF5ea0YGQU4oFAGZdVGDSjhfY5OP2e3ONK7zClEeTiarwxKVz1NE8VZYlHuc+0uitpPelvTlT
DFNNMVCLiGGlDq7GotC+iobYnWTzo/GTb42Novny/UHuumnhkvs5CfhemmIgtWM1UmufG8yVK88X
AhkC8SIAiKhNRpnGbE/BU4kM+0zmciM5gzm1Xa7bOH4bHmJ+HHM+noB04iQHVIQZO4uVRseWcAA6
j/tE51Ac6RM+M7WERR7H9ujStXxca0Ri3QCm9h0z/lt4rCOl6ZFwPpo9j+Wu/CsLdYHiE/mn02gJ
kTHOyVr6NV6mv06GWby5PLvTwjhIMCjieYDzUBjnuQlyG65K/pYM7A98h0byWmKa0qU6tEoEDcc/
jK3GbdcTsag5c9iZXkOxCoUCfWZg3shHKd00hk4gcw90al8jrH/P0XUYpOcqDYyTkFnb6nTS10TL
H+PiH0o+qXVVokVv6EPrxityaJTzICTxjV8LLkKF4CL6DRoQWM70hQg3V+LxUZq9d0C9a1AEu4CO
bN8fcOrlkcXxKZ6BQAaJEdvpaVHQraFZ6FXFDV0E8rn38wW52bMNkV7PeTFL62Gt+g726n5w7Lp/
RFneHtiUjFKRH/B6niR4j9rN11vzE5/hzeALQLAklHOYm02eTRIK8vcO9IqM6ZZYbS3kdsaQGfYT
aK7lD+/CL6fD2nm7LM/t7gVMgG28Ji9v8LCK3KI/OBXlAPvjnRjSPotHaAaB/jyJ2HBTJV0G+dL8
7wVWkX0P9dQB+lP+mM2d29fp2TPP+WR7hx5i8l5p4iN2fIGN/D9PrX4lBFmAISn+4kzf4oUdcOhz
Yxt15gHQYCVVaoJx7L5H5xRbsaecdamtsu0QhQVYuYeKCZAenSYUuYS7Rf676quInrh+DW7A7j0H
0znD4dc0aofYLJYK7KeWDyveB+alaHqDRwfgZxdP2LcvHJrkRdKOYZws2V8iUBNvGkm8OAhHSIx4
iU+yO+/lkoBGOFBW8uho+BTZABUOkq+2WOjh1t9t+3tmsg3MX2NT0GhztB5XcvZR5OTdkvVMpWby
LPog4Kn8ND6fIZcPPGGVTd4Au4HoEXRVqlvNXI0ytHmihSzOJYJCm9P+FWWDCJzjQ1Qpme29qQU8
omuQ5kHKxu2sPT7q1BFIY1DUcfER1UsfWkSDrwZ0dCN/19oeqdcsbZ+j8gCpgV4SPlHgh7jKJxK7
e2DRPyh6vkkFAn7sUFuwS9oNDLYxTHScJQbfpQUhb3LQM82RVSdo4v79B9cNoQYAsxRCNIi4Nts2
Vc7g5QeKISSg7qDKT5te7hvanx4agZnQgueaBiVgTDfe6f7EaXLpVe4X0cDJUzF70+IgrXe3FDGp
rQJ0YaUS243P+HaK3adiq4CR5uydob4ADmjhQGMU3J8KCi+n4zdj4TlWwjBd3B55uOxCVsEKZXxM
VcpMiVie5fOz2LD3T0ZJoOp+FNCvU8rnGmxxb09ytfOCsUOqzo/aRoY8eCfb0Mxp47c/uJkB3t67
yujkK6BlJb5VUItMdGjp6IyK1wG1nhQjqI/YNRVqZ3KXsfTtPkUBZYCi4od/qZ1irO/WHtiTPYqD
LDWwIcgQhKMImSWKhh8b4qNRasDBvz+nnOfnOkam8K2Pb9D9a3tPahuNWDO/n+pauhwng+/ZTH3m
2GdvVFakGzAGyrIXk4RcU7bqu/stN3TzYkrPcI/du1BHMl3Rl2lzdqMnK2AjmbjqpjJWPq2N6+77
daLzyF249f/gbx5wjOmlNfwoocpGm9wtfaEHDGlDYTq7Bj4VEJ4LeKwn/qsSh3IRTRJ6xHcTL5qt
N75yECW3b/jJnzt+EgZG8S3a4CpLIzjAiYW8eVitOruti+ACwOzq/d4D2R4bojCXqGsw/aeabs2s
tZamf9UYdKL4cqJbCBCS9zCNhmIfrd/iyVIXdD4oZpbTp6uqSTJJN3LBRHQciK1KImqRbh2rLfm7
zqN/v2iMi2iLJw/WQfS61T4LUjgyx1VKeaxsm+G92f9qecmDG5c494EPiOwqI8LUz/otwbz77AsW
etXdkLBnwGB+Yz0XWPBLpeaK+rhJF92SE4OLf/p5GvdxJGsKjrXL5CSBfFPnHK4oet6pYILRSgoA
XrKQSRiAzzZJgJoBvgNSufNvbE6uzlgqMFMg1AGGC6fQPcDIuozrY5cETh3xxz2A+MND2dukYeoR
A2+OYUH3ZHU6pjEG63RV7CJgq9pud0Xb2dQRRVGhc4Ptkc+lI/OFAX5rM/9RkJhLJFNzzgRJTTQT
zt7XGB/PPCJoP/aN2wghOYTuZArsRiNt/Vf5myX6w1UCg0XDj1sASqPZ+915UPcm0gaovsjEntSm
lDRsawGHIuYQL11xE2CmL9N/WxTSnDTDmN7ks5aeihbSOgTMKtwpjYk8ZeCGIFNERVkI3FhLqgY1
dy/sGpbBwb419pFAo/+zUuc6i345FkzYG7RCKsLO+aNiXpkt0wv2/+1htzBiAIL03GMzaKIPl7XJ
V6q6+3qhgg2BojJsHdhtJIWV7DZ7e1VDupt5fgduZe4lAxQ23hiSs+ydCwx9X8t8oaJ3E9wLptOi
tmUOBz3MPWczXBJcMnygWNiPmghfGwo7oebUtPKFJj5GSCfPoFMQBFA5OqONiDEL54FYsgVjBTel
rH0Oi+z/8PihBd/lzCe42+2wr0K/04xojlOidyoDdhtaaaHj8sGcNozuEBSfgMmZkZfrgw6/Jjei
4KDGEHOtohXA5QGspPQIcmpPkL5n7lTx34zWmgzXCNbXUdCjRtjhqmtLCBeC3qRt4UcJ1QPnUXnd
nXrYMyNozUivDoXHdmGK4kDKSV4XZV5RUDknHHMjL7S20kDxZeKGOkbdU22PidqEaoRa3r1PxHG9
JR82dG970v8A+/nEuU4Vup8lGjq3F8E7+Cmwa1EAtcmq8gCxvTjPwrAuUYOYU2ujMaNKa4i1CIjt
Fbly96qXSk7udfwilshVxPc5vRyzJ6lAOmLojhhzR8fAeQR7bZiaSVMkU0PrNjf8rQ3IYGzUNnk1
IZZYNfKjRmUBUBTQJ6yxWxZwlQ8Lh3LJTTwLkzHGttZf5zn1KuZp1OncpGxWFojjgQ0kVeHZKxJb
ywmeoRYxj9FqSVU2A9bqLARkxLpad3SIQuz4u1TmWsBE4Sj6x7dMHbRxv5bER3/uuN5XVxSF2din
SPyICEZG3YaxwQMZ0MoBpj1khZS1hC0c6dCoSRRqnH+1utBzJEh8xw/TolnS6bis8uhhCJT8fdWN
rTHEaf3eP8MudEWC+NQzy/7BG+C+xkVITd71xOwJYwIlJW4p1Qs3lQWOYD/IHJeTUiPqIS+Mp6qI
Ju0Jff0YK9A1sYRMjEuRMzkyMLeLGdeU+ZZMSkPtdQpnXK2ofD/b9Wxl8mOvSuAzwsJ8miJho811
eFiVB/4vC3kWGnC87Ao7nXe8bFkhThGHtX2C2APyfNSzoeIDG/mxFGYQBDBxv1ErIJJaeiMnW1qR
aHP68lHPk+/6HLGm8/leM2KJd6GeECRrZjKaA0GoEwnNpm1Muz8Mn7SeiaWpTuIwLcrcMo/ZrgZh
PPhRlZXxUCUw8pwdfdJXG2ZYaTID+lMiZgnPj8iKYQNgqDoqgdaVBWiifDCr1FbzLSpOnuuyDZRd
igukrveiRsj9Ei4giRxwnVYPWaeRLkmH5rgMcMQZSWkUoOh3YWJCJOQBc+bv4MzFTfEkdRMfwxIH
DHW6HbLMclOtrYGe94XgpFLsd0MxI8zuQv1e3ljk0vhg+kG5rhrT+oiGt7YJJfb5EHzSU5pjxRQN
OReQuWZQTxm3/IE48pGUN2IbMz9Ii3SsOuhpNiRl9nkxCHznu71gZYKCEV/C+qJixC+uEKIJ1wWD
wO76Yj/BoL00fDWvhHoO2zYRr7DS5HM/WEJBiWWGFyqVmk+avavfR+KNuWhad1mzrCChQoGVHwZT
VBqSGawwc0RNOryXavbLvyAFMmk7N8EjGNvTkKIh89WURIcZZ3BT3SOPJe+WgUt5XPLyZDu0N6f2
gj91Cqs4rVBlhTPUFkEGSt1BtlVoOmu2+nIAFe5/L8de3nNNyWjntCEa/PMVfA/qrGLIah0tsdRu
34f6CWCx76s6xlWszi6UUwQxbIpm5G23veTfvXpAXrnAkr7GtUFf+ktbwaHOGZC9JHu9unft4iOb
E12O/5QaPvWl3QXHkH9L8yr58yK+uY78CrmUHovY6a+o70bo7TkI0LxhVjsSIpN1nPGoD8dH19Wi
g8DPT08Mc9vBicmzwEHtkaLvBulwQl1BWCAJ1CosfA9DDXxvHg7z08Q5qLdEhCPNq4d8k7XctUHP
Qz2oz8Z0lI7aMwFXJ9ti8DbaKXdukjGTVpl5j6N1m03XnuZLl3p6fipdr0eWY95Dr4TR4+gymVW0
P0i+/7ZBTeK+pelozX9wNN6hla1Jx9/3/O6TOKcd0w9c7SuL/+l2xEd81TUuuZ10Z5aFyBoK0lL/
7jQqdeBfckttxyUYiqBAidt9hAP9g+lfdc6Vj6y5dwhHr+LG/5QBGFnFfe32l0HWolIFmbzhrzS2
VRBJROv2WqdHKDn9ZWLo6boXxL2dQACUI1XTjrOf9fwE8kr5S0R8aQxa6pPqHozwUDHRdzYf0t7k
gKPIEgo6uTFUaKZf0tPhokxDSz+H4FfNfAwMRFUbEw6R9M96Tew4F8yCARyFjpkn1HKzgi7po7RV
aFlfAao8Q4d4ZAAdmvmuvyZdSkgrFyWz5C1XYK5xftUnU06CLyjeHdWvvOLVNtkSPZFnTyap+Bug
+6Y5SD0RfIsMTemX5QN+CTf3Kcz6wUORFa8c7pABoYayl2wEPDhNLBs4rVKkk+5sG7xeO5+ScwEJ
W1uOvs82o48w8SPxBQ7ak0KW4kSwRC/fgxObaeygv35CfRYAf6WXJwlpLstp4PV3X3R/m7vN9xv1
MD3n06aZLYA3u0RaBXBDe69s+CFmsu26oI09Egs1TVuCcb0TNRsSifkTopCwi2zY5wfaWIMCD7os
so1vfexdu/yve6+E2Td+isP5r3llODpgTpNQ0+7HODrW5KaBuhmDN5CcrSDvjTd1ZltfZGC5rtWg
Yig6H0oxFrl00OWUI3LNniMF77TF8KaJsTY38DDa8rR4BK5TsnWwb7yBMu5ciU9a09VZ0r+1/UMR
zZylGxUkMepZFhs95tHnCVBY1ODC+rnm35LaMT6NIUTVNZBPAZOITYxo+9xzd++6VMWVhz5srgpj
HC+KnHVGMBxGERRrUb047i+AoT6D0NNPPCFduikvOkUW7Zf88vwfjuYb0J3GCRENhw+rgvDUXjx3
ThbSknEHbhA0JfQhmaf3qHAnkbKslbAbB3rX+lBU6uakb5rmHVFXz/yUgKLInN1uJjVsg9smbFoQ
/pUO9QGIEv1ZI2pj6VL/Cczvnjx9H9O4ll+RIe0/4dZLtF5WMP4s5GoGj4BQ3jvCnCbZZ33ivK16
4HJFxk0ijrz2YutgiDRLMtAwO8FScs6Ac/XI3jBw/9SKk2H02hckzbevjPEpbI7SysN6R92KRS/h
GAEX/r/e8OvubGo0etzHNHT7lrffu1iB3cVqeSvVhzXZFzZIUosvKkZuYtYZA8H8PicHsewQuCzR
wkQoGbydcxuSqsqdSoYAOx7pR6Q0uOK0woo7MgplvxKPNJ7RYgoIkIKTE3Lbs6yatv/5yTAd6Ul7
mUxkE4AfrMFXerEM195+p3Hrk0arb2RAR3vfEVJ98U7YaGIWc2dr9lwow93hDSlRfVMxhRPr0Ac6
C0heYhkakS4r5NgR7PrfN6F5gvJW3oUhQBdF2398nfozAQQbq6gPVZ/ZJg1VHOhO1Kilhih+fFzI
aWpFQ2WqDH28639mTGUJsmgx6cTsoyjfNQeOuomNDG0xtJD4vr3M3th2I1OgCa0m2DSRoBN3Il/V
tVUkuvNH41eZCJz9VfnMiXFQvAuIE9hefqzTsSwSfxFtDUZSitrHD8iKR+C7Wj0A3MJIz1IwRY/J
xoVgVVF4eBn1b88RUfjCrBBGo/3aRSa1Mjg8MS2gfSZFWNPFGrw4chZQnOY4puGJtwjgBEbkvL8l
eOEvmbg9Ug9St4I9yz6RsWgViKKY3Ap13qQ1qrMVu6FWpNCv/M8YOSRhXMBj3Ta+nVpY5nKT9taE
j2SoKnTHz1jchIETwSHvlQhlHdBVHbdYV5SKlgRFgLJTtBvU4zKVNHhl5QNQfGUO8iLe/+2c8cnL
aRDdiJ1n+khgbHDm1RsqyPOU3pNmm6QbyDJjVg3Y8eEAlUbEKpCFxu5tfY86A/U8QOHRUPGFXTal
X4jFLTZLRJW7ngnfmodiHdxnmSsy4e8LhoM7RdEQ+2emsQPSxDDyjsIpLzuqYayctlYGq2ymN/es
2XiwgJFtNRd48h1ZOEQAQoW06quYpYLQgk4gQX97rpgsFNpbi0CmnV6iAkBfwcp236wojsoSE5Bz
YEo4fs8WYQqd6m7tvJHm9jZOSOJsA37XxnJbBmNXNFaU1ZbA1kq4inekuwCT36YZpvz83SUfLie7
1DVOgjvOMvZD8NF3XxWcn+5GJmN4wKTWxTWf1DfqJfMxLyuX3Od3Rc33lcU4b76hQ5xSedCJYW97
y/FmUSuW6o1vL/1MFKud+FpvJ8AEctps4QjiqUlMfYxhAU7RtWzljMCZszFcIPpWZ0AzgAcochda
RupVBkAdtFsDa/q3yh0IDc/jxDV9nL0/xZFE8V4+1kSJsvIPo1IYdsKqPPtDihlGS/SN8U1AFMNE
YFKBdhadi8S8329knAJYbcgzZsDuJvWbLdMxhoVyKx4tzU7LrT2gnC1GVEEqhq28GpztCsFqA6Zf
TJ7RIs7YZv9p5ai9F+wsczQEs8jyzjMWPjSjqy6uDYuJpCRSsu4pRWjgtroztWw2IMjnF+mXNk6s
oDolYxRmjHhqfdxo0ldqhJ+bX0+KhgUsUiEv4W0yE6pGTkgpSriQnewRXCFJ9NPZxk/jEnPZY5kV
pdMQcJCd7epn3injx86yivdNMhzjx9G04+7ZO/+aPH4Ceq+yaue3kJAUEMPBoaRWWZUMzxA2zFNF
IIiWbVvbs1PI+cGhfdv1cG9Z9+cN7yr+TghyzdBPfdj1aA1y7z8aneyyeEWhN/C2t+lFIjAPnolP
6g1TjMZKZmHPI5KBM9pZfCIAcHp/M9vag9Vy5Pupb5ECwh28OtejQyIL7hcZ4+jGiS6tku3GlwP7
KjovTxrVbo03B5tX2e5U6mXzDwRKaYqm9+oXPEpKyRB6AMxOwtLacmag9AgEF8/PXlK8XxYcWdew
+7ZxNeOZMROrJSj3TYfPFbUc5Au2HELmPekeTcPPKBUEDBA2WPL+DwceqfZAAJr4lep4DZFu6fN9
5I2Y6oeuivEOnEiFJImtthnYS2zWcU0pnMvixVBgpiOKSPnjf1+8tYJy+Yv7ZzOBjajIhQ83SvmL
ystbKW+/Vfw3KCCnhMqJ6dN1rp6wfYBrFpCtcYepIMD7xDE3+duZpmzS1AqeD1I7MwNMcPveYRcP
VQLbp342BPK+SR67owBohccKhgMpWkJTRKSI012N/TF2uMOqcHYHBfuiwDxAqvddw8KG/sRYxYLA
YRWtiSc9/NurJJBHwxOhP2oiBicYTuK9/O8Ejj5zSybcVGCrj+TP6zlHhsD7tsMCZhuQ9hGaGsNN
5flLpH0Hv+48Rw1PRM26fNpj14tlJDTcV5g4rxZhuJwDSffguInUjwp4RnL/Uqn1yieQWw3c6JEo
YrhWuZJC0qKf6INKXZeqviGstCA2DnKDBVtCTOs8Xkibnsed9enfcSxSqdWul9WhCK7pApHqke/Q
zQ+kyOMUVuaKDN1zLZ1wIYNfP8lUKoXRYs/MtaJ9oZMRTQNbHrBuHPUr/WBjZbKuJKO0r+w+R/qs
baWxDZSEFozxZdoc9Bu4PGcX1R9K+CWXRMo5plr8+ZUYAYDFkjghU5OINwq9sFYqyj+mOGsMEpWZ
UyOHyJ95THefMkiICxoaC3P6LCs+aiPoFBclR94GFilSVGLgdMoLDIUvENuc3PEKIwcOrlu0GUIT
FCGGTw31Xp0bOl6eIKc0z2ejkHMopWYOsQdqxoBvuXuN8I5jKcfece9lH8Q3nDXsk0U5tSRUSJSq
v5HPs5wZOOqr1GqFJ4dVfg42N/+hACqstWjqowMBMq72D6emotGoGUVO42r+6JS764u3HP7ayA0S
yW8Vi9zykh/H4sD7yWDHn8DJN2/xVjgNoIBt2ppTgmSlJjiCbJwjvJ1QxEEV+ZLqjvn9uL3Xy2Ag
CKOwHEXkHDRHvizvjMldxbkbKhth6N00sLJBFj1Eq+1AGqG5hQZt1c3TZhNGeOEndZDbNAG52RWk
hac9PL6OKJl+SbvU8yJwfjzNJTHitty7HrWDziGpN+FeGvBvkOap8pVXjU5URbI5JQkKTi9hyIdv
H/f51Mzz04bSUh7CN+LVOBGOWqCnjaEIRVRZLjs/RlbtreHkUNNxDi0CCE9kCNUmG+sBkzjxtA/V
gPDWT105UL2YbbHqIz9xFfpiveDq/I3A9hgEtlVgeCnjcH3NTNzTEMvfN78fiGk4DgmENJ/BExxq
lOAfDqXqgm5/ruALexHfYT/rpd1p2rSrwPLxsNklBjuG1tz+vzXb0exvh6voIISewNuSTc1bKJWW
+7VEdlKkAj6VSzA4NnVjnzC+mj5vhAmHW1PiPo08tZsgFS7jmsT+Po4+mFacu4PAXMB6Yw8RN8Sj
k9QuIQOXaoUGFUBg50scZzcD9on1ebK//j+gLXh9axo5YqkW4wLiPRMJ4/T+KZPd4yUzfB/EmhgJ
jDsDQt9GPFn54p1k112GKwY+nVAghivlibXJqx/rHBqkFTuP/RA5TzPRBLietnN9inR/SuwRpPSx
+DkUxvG/AbS7l1KQ0S2Bz7+TepmjwXVvACv7OCgY4IFJ9HKFc2e/C8DdFgU8ehEFPGEvW+/5hqHX
UY5u8jq6CIFsQQdSeXdwHJqB47252khJPvIyNRVQ4wwnFQ5R1C5TAGNv599hWUpxU92mKmCUvL66
EloVr9+xyVg7BP+61CtXIxFT5ra1N3HNfrH0dNrCzh7yoev+tWsdRbyEOGVI+jqaBJKTmeh3Zhwy
VlVrdldVjwHifqlIFjf4dQxWNbH55OOb4KwqDaQAgiwnsERzpAFTTGFisOAMBLpzKPt0AaEdtAoR
fXa5IeeQbU8Uux3HzsYKeQjqxEjzZov9xUhlR9sU96RwbOlfiTRWiOoJBM9P6IWBglGe8KPdC7yz
b+9YQnBsrZL0hSljmugAREf9lycA/G3Cr0L7pIOP6dEZ30wvs57RoIpoGii83W0LEyH8DOz05ogX
C2l7EPJOs0evRbq7tZjzn4Gp3EPNKkak7Qb2Bct6A4hEKGBlvakHD7qmu0pzvpD6Pe66HGJUM7hI
qkC345y0uhfTkXSjGd2FLjORhtxpxExRnBcogf37vLty0j+MnY4/NYxvKNK3Gp6VgdgTYaeaJuIw
ugHCBJXvNEJDMYBIG8dOk3H8RT77Kh6OW5yMtNxhu5ITWFxySitK7NB7YM5USODGERp65axrxT7I
5/LxyqEIrT8+0wzVzOhHcOzSq0e2q7+MIk+sDyBQDFVmgHbR6tVKt7TNx5Z38Y6k1lqSxSaApUup
GXoyiu8fQPRsmB3GT5t/8sD7agtbg0+t9SdwT/jZLplRGJ+zfx1UqtSqPty5rY+DsChUB9exvHmu
V+UN0CI6iK9cM4eSm0/Zrs2WEN2Dw+Vzt4TckBa4cofzrKw1AJhpK3zbu7rz+gRrcoYDwPyivOPJ
Nf8fGBOzrXYoxOP4loTjNsZZLkooG8sL9XG+lMqzc7YSuMzHmjmkVgUlV28F4fb+UB5tV15ZiELe
dtDfIQox0qk/yrbAi8qA55lxpbfy47M3JqFWseFM0NdY85sC7945HqC/l5ShVgpanba7ge70x4hs
dHpITcypITFR7WyBVFL5YXhq3Beg4vP36/AWpIvTbNpO14Wfl+1TRKBFEc62r7sND6wJofZ4bhyD
++aNudQKi/fxOklUMi0lto24F/yLHK5eclmrmF8E1i3f6+TE8Kt0SHWwjza80fJrx7aMCDP/XKpm
C6vjdberXA7dL46xsUIEomEO5Ab4E0c0u1hujdIoAysPPPIJP+YdVVnVSlry2wi/CfxCNDcvKi8g
g6dH/T+ZUlp1YKusOGV2ZISPKHBUcapTLmXjhDCl8cciJ9ji90MQ0lZYcl6SkACRE8lp/8bHOxVn
EVTvtGHy22mnUm926pstxk4Qc1YPGXSx8SuXG+2i9gxH4R8Z+zUIWznNQ8+aY0f5d2mvP4SBEFA1
M419GoIrSDd5NSNcmNlh4m/mjLNtwpbkUm8hFEyItwZ14I3mjhTJnwIVWkUhz6PrOkX/4PbABsC9
71Ly50kQepXBNqZKeRFDlr0LbcUKqh8wKNA/guFcLoyf41CMc6k9fPfSkCjRhtLxokMVfQa45+AG
JcscycBbZsD5s8Ut82J/++kXjx3+M+gYGK0Gtz3ItU87v7Ifo1+JJAPfrVAG6mkbkwG9diMzcqbZ
fOsAYeXWUnC56cfMaPSudezbEMIRUVxIRmhjS5IjfdqzJZpQnD1ig173XIoT0Jt2KSYyuVLly1Dk
oKEde0Dy9hJBbzr47EoQzRNoMmQJP1wf5WWQ+joOEHcZzO4iMiGdRRv6cH9kMXyut5ivUG2U39Gu
uHleyo2sqJImmdauT/+RDk2q9f0ZC9WfQpU45u9pu/vTYLHAga1t8I4VODseLwOqWGFs4xCYvujy
fTLJl06ytZNKHDe5Nu8wcx2NmAA5iw3IUoemAH6Ugp4LfdbZcLbsrh9Kjngxdso4DGE5ONLa+OmG
ljBgu/REeIZM+tJxrJfvO0hzqx7rrIeBotgbNJsfdZBfKmWRVx4FUqeKkmNuM6FPFIoQNcVgnZUb
8dlrNBnJ5TwZBG92kCk0VdCJq5vyBJQ8JQNSbtc+1a2BQA3oe9Z2yz+1NF8dQBYYpvNTMBF7HLO3
udA4XkJtgbX8ie6D1ovQ8AZPFuoARBRmaE5bxvgjRs7dvuM8C9xyFfSuLOEbdu4s0RF281//kyqa
bvkVOziraCr9roRQJ/3d2lsY74Q2AcBixcYFKnFQUUVHEhBZUSicivTXo3ZFdalgCcR3pJv+iwN/
L8Vivdol+nnlkUcULK6uDQ93JmhhkDm9jEygVqMJmuc+m0dAY8w4Fz2/roqts6tLiK16GUQmAvIs
xbjQlomTIcyDbfVPF93WFzcrrNf5Zvcg6Qx61ttiItZ8Xo/BtMyocGOxXKxSbL1NXMh+1Yvq/zDm
ZXnW1qQ3OyTOuSM6zCf9qe8b9UL7I2OGlwS1Y6WltjgzJ6qpDMNE++k57Ox1e1VacEaY8/akBd7K
TNm4fWDakM/BqZnFmjOCAezFEJvgHUARiLxgyNi1lM+ihMBXltqlXqDb17DPT4uZX1BCtxCM7rhO
WqzHUz3CSm81ZI++hEU1hCEprJxsSZBWG8I/AdXbUur793g5lZTe6Np80v/pM8yj6A73/lTJRqvI
z+7GwgCsuWPcx25U/T2jfgcNPIaZqjOn5hi0z5TgGH5JQY77272ki4PntlmDjcS9hhxclbiqUs78
bXS2sLhNU64xJ7IMw3JrNGGaRbyiobUp7oRgrK4Vzv2201xdMNfWf4NR7DwH9cWtZO2UQodGHwE9
kfGjSbvJg/eA9YKz8c+BqkpwwCGZnzoUADJchYPMCkEY7MMcuAPI2b4X0sC9rIHQK/upBarkCTsU
/Hm6hHo1SFmm6GZK+uexpzz6HWrd+Fda0zis+Pu+z/TPDbRemzP+KlVfSGd3yVQGZ8LK5R/pN+UH
d1JkFunMEOxPvFrx3T0xPW7RbjAJSJKNLgvL9PzsZAzCeY9faccsn2HwyCwFuJ1wkAVJLkXF0V/E
ih9w4li3+6HGjWtNqVeOfHy1eWHpulu5ASUtA0WL55m9sB3qDzTvaas6WdlO6E0Efup3KCuYai4a
ih/R/nRXGJ2VMqQ/qsZep0tEXP8gwdHu1jYXVskxks1tm9Z2YIspp4y2hI8hSDdsuAiY9byabK2V
Rfi2IgjIgviXyc7ZlFiE5kFN9HrKit+d9th7CXZNv36D8ZkOIXkq/3nAqbU2PO+P3dxKLIG+yblb
GDEzNXK9RHhBMyJplC7kGzl1YVfV2HR72laJP1ud5nP5+qES2z1UL3sG1YMXbA/Cr5EEUykbuFd5
URWRiW+WYWZRwhKeTm3TxAVYGHqs6Qgj7PmSkn5ifMnVA2yuDAHlfCXD4sdGX6swpcQSK9r59+R8
PT21HIqGYkevubosTdH4qY3aR/pjDTmYXUWbD4ahtVgCiS8dFTxiyDq20q4LitJv6if46Px3XOHy
TztqvLiazXwyKP/gBdeaNBC2bzepabxeSwneyNPPRZs0A30Mgu6QU+a+V21xCPDLSSxoT7x4fgJp
0k9+RpBW/gkqFKM6ZT22U4EAtfP1RwM5d+Y93qj2qXvLgsvUY0fIrsHXQH1Wb03RKVyt2l1V3h5a
IklljSL0VjItx8SyKSYnH0G+ZMdZALm35f4XDn4l4aiacILb0Xjwt9edvx6ieFOoONczbN7AFQ1q
w7LhHsokXMA3J+MfuQQyJ5VRxCfQkQs2wm6P1OQqRu9+B3l9HYep9NDwpCNZzQo7BjwzH4MWn+/c
FXxoh4yY3ZaKmNL/3RxSZrYUqJ5oFg+y8ra3OWZZFCDL4eTNm/ahWkAluZjhMBxX7P5H1Ozjvwf3
My0dJAV2B0ZTBJzihbyExAqmp7kfeRYCedc4iiGCxWtsylOTwRgI5IIBvWT3vgdbgWjG4ToVd7O7
uL/b/Mdwsyk4J/FOa0fQfEQYpLZekaZFPzv+WhNrYenNjvqfZIwPD0HxJWYLDmHL6s79p6CVv2H1
VbseuOGaueG0Fp+XYYrbd4RzBz8x8jZkF5hvURAE9Hq6meatkTD9dUNskcbjdCcepjOv8KmOsKMP
yzcdnHYXFwXDADjyIiOzdd2gwSRAqSvbygOHQCIM9RLuldw450F0FKysLzWvHUwng7wngXQjvll6
MTdSorjIRRElYjOZsMqziHwgKLxE63hJvg0So0NWmrsaBcRLw5KmCVQQJ37pJVxOCWWAtPSRRz2+
3RIBh9ka5bbqRCQNI8v2bhW1vTZXkPxbPcqdHgGXmlgsbX8zonHpWP54EB5WYEaz3OcVQOdv2GVA
Ay+pCQgg2Vv4uPzLRLfZ9IwdcqApvUc3DbnMxfAZTZlLhrmbql4DwoiyXa2vMfvc9VLQ/bNWsa6+
Qh6xrnPOiepqjCsQu2Rm2dU5WD8bjPUg/nGgHNs7hFxYcnQnBz60OyrUDU6uSYgLwpvdQV7TF0n3
2R6ntCkoEfFXE5VncqEL5dirp1qe6JK4ejt0zie2sJcSHxlnlkcqgg8Mgu0562iulsvs93b5jovD
mZEhHhUzh1K4andgfZDfQ6ASjJANAWor5LGtRLoGQbSfx2lPgDtBjz0Tebe5z7dnoVow2gto07EN
hMANW0JgJOgA7KHGjkPo9dPLgVoIbXkv2CIQWhOV4MdhW/9Bus0TYwbEdXomvlN9KGixY6PEdk+s
UBNcFGBifS0A0GQK/cPyZ6QrNsfRglamdaTJmRfFb5J3w0QDaGIwaS50/pncygg/htOKe7VPQR2r
atXZRY0BRk5jiwxTrT8cbEEJIKOgR9HJ7MzrCmi9UGf3qnr3IN5mqIc+z+9rJgoDdze9lZZLEekk
S21CK2CS2Svz0WQWJgVcjb7VGEUsMb0uf9s2WzT5NyaU7h5PEYTtWIxmMgUgZArPlTDM0oDfQuep
UAsSSR+yPPFHy6nuyZZe28yL01smqT8/VOeSC47q5tXSS+kMZE7ldvb7cNMy4ON4PrfJ3ZaOMUy5
ANhHJMXWgQaZuStkc/LUqEKP6TLVsAHKmUpPZ2Fmjb6cRyHfuTZaWE+rAYNsucy6rzS6Ll1fFhzr
gHOsSBmsn2U7uoKOLoC8jLXJwLPK+eQbnqWy3nVVlob4P/8SLvAQGvJ9xZ7Nl25PxARVcxrncor9
FigdAxF83M9rlweL8hbSUkuoz4Z1xEdWDNhfaLd7f39KYPXsDFSkTj7nn+++/V1fvMweNVWNSVHz
qC82/OkCp4FwG0u54Uwyh45rKujp+iq4TsoUgKaXpj6g8IfiHeUOHCE16j8q75HdNnJA2/gCjZyV
guvkrcoV6OWhJKnwM7ZPqWbllYiJtNLWJ+g7+pqnkuIaAbzqRT6yLNxTdnfB3KSofzvgQ4j+Rhv6
UwfPfPK7/wstWJ+ncdVxqnxesLaXWF/u0QA6P3JkpG780LULU7cHniS0AFxe/rp67Rg9eqH2pIHm
pobra62Wf+EMl1ehU+1GHaCFMSwcIYGxi8DxHBxX8i+vb3reZ+hXy0M0l6GEJ7QjAfTWNKF6MESe
gtHaB8Nc351OxpvgLT9NuOLjakRzsam+gz8WKOkMTMAc7UgIB5Y+vlyHu9SMFttFveV266JR8Rbf
wjjmUW6ynwyEzu8mumrj+pRf2YLwEJ88DA2c8tp3O4WWMU6mBJVdqGRBatzQV4Wr1Dn3qJUY6kLD
Qrkd/9ivak016RKuYIGM0lT8AMpCABGHVA5bcFCHVoIW3ZfXO6XePfyaI4OuwLzQ2AdToJ9gJyNQ
eLf6qYU6PmKY/81Iz0maRpNF+TbTbbJR4DSrh7pVomxHyM7Kxi/UF6bSGEH2kAQF5ImTwrdqS4nF
mWOSCBvLrxfhxgycOLFilJ0XCry3wn5xYTSJIgnJSyJXuxa9qXIAJNKPTm0a2Xd2zT2QBDUY09dI
U3sQahKbD0C7VugBJ3aq+NvvkPsuipWSAqoj/CKEiCxFEXMD/zCHqDk6vbr3cxDtxqgR5eDegCjZ
uGGk7qll0eqKrCfMRaH3fmC0xhXOMSUXqMVnnKHHDpgEnuVwrO1xVU4jgbQ1xTj9GkCk2fr+A2jT
YfcXhFByxsZs6GAM53NRVkUc0AKGCUApOaoIdQddihJtGI0F6W12s978gOb/wUVWhBsDw5wryX5g
3c3OsNxgrkK1N1vZyV/Tq3Ev8O6h5bWWhUDr9pnbg5DnudCIDTae5vVIvnfBcQtCNdVQP6Qyu6lY
DHFhX6uWZtR0CxN635GN1CP5zl3VOk5kRojmvMf/vbwx6OH5NEkEKR9XwmDkIG7HYd7fx7jkZ/43
s/Gib0Ecl1kzZjbMxGPu5wUddrX/RAkHeXfzaOAubh9C3JS/3k5PdQUJ4ekU5xscett1GyqB01f5
D7dn4eOIoyFbJo8A5rsfX0i2m8Xo+0F5ir5TrGWNM/mu74F0e+W/sNn+3UEt6inRm9XFRkjN25rc
QZ1nSqs6xYlVf/OswEK9W7ZOd9e27yjUoPfcj8u/dow0ODBIg0RrSS63uHLhgIJW/LcZI1vN979Y
pbTyGzi7GaHWWoJ0RhvyNi0iG0DHkkid6R3F5mlOsavRZY+m/Prtfx0Vx10KgnpgVtQJvbt7V738
h9Pla2z78LFD0LJJLVFaTCekJCr7P52GY5ZMveBxcOTGiLaKbvTBjzlAXn8T9vxLZTHEd0H6sCNQ
STdxSAIEQ6bYk6mKoBRwuVApsRA4AteCF7OXJXdw8BamATGxHM0gS1JBE7gU6on/ww3dlyLN4McZ
ojbntfRbA0YU43il3O1zATXgk7lrc/osKmKDOCJ27HQRdAqqsjJbNCZTgkHp5wqRpJWb20VgqANp
XQM9/brQJ5wmHgJRcH/O3VJ2bEZVLvujX4bwCjjrv2O7XPJKF4a0pv4kf0TK37CqS5iE8PNQtacB
MTBwTPOyneXvX+TDnD7aWSHuxKDZZYOM5bAF+VodOaHyy7DM1fTIn2SmyDvnh7fKITrsTTTVYEp5
ShWWA0NnQwOGZ8nZrBq9A84ftNrkGV6GW1nTB1jGAHjwwi6zO7fK/jQHKhMXU3saxD49J+JeUJT/
ylhP1TJfaz2jI5lK8Eumuj1Uxnj1Ks2GkW+uaukvy+B3DDhK7OXqyaw7r6kMyTP45Y0m0njn4JNF
uklE/rrZz6aEBlq6rjhS6CwmKnHtMDOzHYU3l0iYzVvtotJUG1GaDp8kGnUTmtdy5iajyr8em/NI
XvJegzz+Lpv8ahwC53TlLXQPQgc/rfRf5bNF9HGVInTR724y9C9Nitc2ssEjr3+xCqgeBSa0YocK
NNBZhcyc9v6/PkaUfemO1zHoNsoDCOroczK9IgiBMCf80PpGhmBMxFMB8ZotbD6t5a1PLf7+UW63
IqYRZxGRc31AR6IkBooGwK+8vrDPuFToHiLwLvPFjmjNQiLPKz4f8A88l9e3Zb2hLlLlVJ9rLlZv
fufjHjIXqva/6g/94WrFbJSNJfkiiDFor2hEV/28Kpjo0ZJS0JIkE7ZVa5ZngfGVXc1tHVGxTnq5
TJAXEOnZzMlN6BdG99IpYfWagwf9DpTJ9xehblOK41kE/+VrNckWo6A4K7zajm6FXrD3aNo2mPHF
0b39xTPe3icHBY/0XsZmi08ga/6xhcnFNCjiTdGowbFUf86ejNcPSyYTklYmW7i0l1CxtvN+jDk5
OOE/w9aauLz1ZC0c4tSjMXu4k2vhZJcRxYhlQSndLrQz6vsmBIIE/pKP66zXD9YjiZ9yzXZTPiCi
ZpFTXm6ZseFeqqAKGOTTNgA27MCXxZDd4h4uBqT19SqE1u+9TRW76bgV+9i8wMfMjOWTH6oLJw2v
RW1PWV1XR5xy84YoR3Fu/4/ar72BmHy9wVzA8zdTrxQIZ1OkyQzR1vam4XnKXJTLtiRClxkwAZ4e
9/7AE6d90jeTSuQOxODCPwtWFyyc+vd6dM68wIoudNKXMukIBnB4S3dcXn5pI6YvJr2YnSViPc74
43nqQkQmUfH4sXMWSeZPy8Na+lwIcYpgClMIkaewI26SOPbnFN1oA7N1ieu2QfWaVg9l8LOsRoi2
Vcfc1FqKRmaqjpmMTBITmdfZA4s1jSyvyNix6cIG9vVyLUnQfMiX2velQAga+pPpHoNDfL6apFuA
7TW7W4iBKjla2/Wrdu7+d/t8igEFsVDZ4dk9BS/RuISQJ94WIODTphh/pAnxMOPR0d3f+YowLt7C
mDo8UZ7Ce9X47R1v8uC/Bm/i5jRsBkHx67eDs6KBQ/yj85iqlWtmYNKggjYb0tUbk7Rn3wHPNOWH
Feb0PTqDIWsMlM/i/WYttahmVKQW66LxqJcJMcOBo75Iq7TuvNQIuePRpWjeA+GjguIzHQuq1SZW
Vw+9sEX8qv8bVdY4KXKQ4IodGbA+RtT5LMuJvIq8z1MXZ8Icgz+BCLqzADGRaMEYY0d1wGTKLzPx
ZOunK08rc5ILqxbD4jezdolI5AsHMCpctVgUO7OfAGruJKVej+7bQce2GeTnNeGgJ/7/TuEQ8/Hu
4R5fiqsPa2fWg+1ts8OGExGAB/LZhA8o3vWTzs5cMWBJlB0UyI1d5hjCjajIZHyxirwSxK/+azIr
WVyIYT7ZpKfa20tIAMIOP6cc41PTZoRpRPQkgmozXKqGPMpFQvG4/e6ux0TolikG06xiWbp5xjfj
Vivzi9IiAFhEYVw1HBKnx3zXgmdYlxu2W7y+HRxW/NLwWpQnBfKtxRbwoxAyZxAz+BPtOJhCf8Nu
Ju+wQhfkpn264kOoIEEImR0RFCIb3u7d7nGdcozJbKDN24ULjKMMCuk/WQs0mFAUf6AYHKEcutXn
C/T7KMTyt+v28v1HGvfgjit4p+0JgWfHiCqggcSeg/GKeCVdT/9ox97o8/afZ7agvdVSzNOi3PcJ
YeAvTjy3QkXI2gThTKwnnSDAoSj4uHNSO7IDQJQQ8RqsZFTr6dV1rXsxxdKpwcZbl/gZU/Ciwv8Y
uewo+osbQN8kZSHjRj1MFCle9Wuor8JI8CKNpiZJOFGJsMzzW5jSy5zcg/mz38rPma8HfYkTGvX4
OsOgsZmJepw37TYsfvI1a8O2HUrijdZ2GF6lo3vu6tDovXWTdhEsEuZi2NrpxJr/eTT4UcsNtWxx
qKjIQeVIyIGXv+QbmUK+oFGkzWt51U7GDClDhNnWsW+rg9SP8S8M5Nl3niP9TJ6PWm2mwkDTwRgq
eU+EQlfxa7ws7TimtuIZyBE4CpT1/9pF3cICT8cx2whPT7afYoPj8012BU/HG+CZoHt5jRAjjcMv
GLI5hflndXRF09aFdkDTFpkV63QL0IFb2kwzdEizthBfo+Y33loOs1BVrfjo5djmiESxH26CvBAi
2x5MgBApgWlIVEQDRGA+tGSHTJJQDFM+O7Mxd6p5/69JinsV4VKIuJrQlcwNkrIJynngWExDd/M+
OyOOeXR8ASAiiitF0SD0BXQkGmRJR+nImesHcktHANpcWd1GFBNeQGFHTGbHpAGuzd3Pwkbo6Gn9
qRu8qcfwLjpyd1QL2eFie4mFYPtjYdWjNd6EJ6lXGg/Kfg7UZJCR3ViuvP5ftrHSKgBPmSAFY5fV
zeCATCYiwBqvr5557QG7IUPKVwy7R7L9eFJx3+vRoWNgZj2Lne3a8UY48tcCJsDrAUDTYJuRIYAm
SV3Yvi5ewdInT32busAt1doO6gK8C1Y55mOKIEf6hUypcapwBTGqDewZWU4uv66owNF2kh6Zd/FP
H4+NDmpIOXgPkhDUbIpOpYaOC/2mLOr1osuIdyxDTcDqV8+3O0wfv2NgXhr0VDFoLXg9JqfuzNHT
6kmqcZobOR1f+m+5u9t6OOf5S5lsbUuYruhV10w2jjdxQDfwQayDnQkv+XaCjkmEzXHMZHCJYzWf
8zeW6gw2pCHKvk3Ne6hCAyDKyY8ljyVOG8tWPx20tQqGjBCcT2rc7UycXUZu+x02b+Xi2kkTRA4X
LMOXjGVpSMitpu8MgoU3edx6VIQ9IO+h1J92fdfSfy4xEMCwdX09X81QjAPd0K2m6Hn6qxhEHqYZ
6QSq0TgH1YPq93HtMGkPxwNBsxXY8jihcS1+WWuIe7YvpyufqIZvDP4OmQyReQFMpmgHsEIr/ivA
W6jR46QhQ2B6Zunyl9DNasEhE513x/mdX29wXN4W7nbQxkJMd/t4l26lZzyUOkQYYibZ/5EOvwR5
Ye7+qMw6+rJLxAWLk51p4/LS4t+iA63BYqayaV4jQkWWeugg+gORZJ0sPqv7N+0NAb/rnBWxJgL3
5IVFADlEQO1vVXdqR7WMWNhPiJJOB4EkqbtOzjIZsMVe6rvxjyi9YTrztNE4vipTqcCYhX/836Wg
Pu5W4ShDA9+dZ6qACm4LdDWOBr2Jgy+l6MwohN1UXNlr7zUHoDK8qbGbFn0I1BsessQ7UkJc3koW
5z+v0ybYAa7WHTq01PtTjXGdl8PU41rWf0OfsdvTzspW+P8rbQZKsEJ8A/vd/eabbhMnzLXjxmiF
tL9YmGxE6HY36a+mDt+YbForHd5fzExkIH9qdS5w060ULaFufCCBSwWBbpsC7CgswLjwmbU26y5z
Y8Lr0+htqMtw3M++WYBQ89t+h1G6k5q/HDKkIBx3ktRl8KDJrs3vI9PsqUQdk9rBtna+gfu6w6E9
I0XekHkOIFLeAOAscuCoF0GPI5etRO28C2PFSbk20eGzSQwKzCk092NUw+tRDjJH9GFBSxTxeSq/
xMGufRYCH7QYoN8YGpqL7tKyDg8MmFvNhYaoaL9KV7Efe2OYr2zuYE3fqpHb6+EZjaXPnqms/cy9
0PDQlUYLpfEz1Dmz8sgdsJY9sDcfBJGLdW4Owddczg+D9lN0XMEXGjIhA4cEAnqIiJ1lpbuSt71j
4Cwn3xZnsojkkqxKAvRuRHn9QoiKRA6LwMwHIJyJl+Dq0PqQZj+8H+vuTbFQj02aQikaHjt/iC+6
sf+mSbAsIcwYxq6ueDG4Hr6oS2Jg63gsRQU9vYYJpkVGmjDTyzovH/CPTzjrEO34kYemXtilIcjr
NscKEwlPAhBpW6nxN8Hmcb0+hRavffh9XfNMagISkBbCvnYjVzKq6VZ18qivjrt7/nML93HEb6+k
he8inkA7b3EB/e3T7uswPkcTM1MTKTb5Su6ug/4YuPdzr6w/AvkUlDN0zVUUNDryj5eu0oImwSEP
DqfhO+4R+1UErbowxBdF/tJriWjDNHnW+eB8y/qpx9/a581s8hb7jXZWLLhbEAQ6iYHYBGGbL+OG
FksbA0Z+yvli5jRgENHtQe8618i75NdOXXYdWbFYlMbnr6R74KXcAcwfSI7j9Ra5uEFyMqCM+Y1M
bLzo1e53mN+NcPP2TrQi5Ach3m4Jwvi6oVjClxQfIEWr0te6qhy7WHhJeGSNnZfSoh7NFDMMl8pu
3kwcu25keQnMV66RO/Z8wanfKTUUPMulZYvM/inp83GsCo5yJGYqZxnWZ2T9izs8l8KyHWefSomu
xYjtkvYcGzR8cnkS6g3aGb8Vv8gDCJt3da/LfTL3RrC/RW0nqvIMomVJlUhnCtC/UavtY53M1MrX
ZpgS6x1EqIFigHFn9HZEiuY5RsQfny2z50VpJ1kgzQ2U7lyL8JPYeCAAZQXg8jizjjcTe2jmVyZy
P5nLZ5t8mDqK0GpTCpV0hLd5STRUfpkeYKQl4ChhJvPWIUz1T/Dv0xMzZKs74xdpID4byQUMCGdq
dTvZReg6hiSSlO+g7Nl+UGfrsbMpZasChSjEivWgWH1GgLs0fi3NMtt6AZGRuGkCAHKJd/OlULGa
nxNljeBy5nOBr732fJogcQhtcg+cDswQ33vm/nfRrJ4uWQ3suFHSStRHl4vU0j4eJhRtlsvuIlW4
bI+OhCcV2tAq8i+yOLaGtrJsCTc8qgpNgqdKm7wtdd56UmK+5LzqhzP3c6yhHWZb2FNf5J37/Hlp
dMzi1526jQCS0KlmUlNyuYXXld9q5bf4fR1qYME/XI2FKhp3TtDAQbSmira6yfopb1LmC7OnnDCN
WLdZpOQ0DtsDraJe427CHCsFfarA1FXvysS2zmJmZSFtRF/77iwNlnARL9pm2E9l+cz3TrkMPEn6
7dM7NQU6Hf7dM4RtjqPYyWp83oXOwdrk9f5kf9m0f2P94ENHf3Mr+sZDubp5xKkRnlqrgo2nQeNo
PbL8irhviMARWrs/QdlZXoyG13WY2CTr8WFv49SDwPySNcdSlkUsmQ++UwJ8bgyLDxOZH1E0G9AN
592WAOCFIDScLvlnpFOH1UpsK60DlwCci3KM7w7nCq9IYTWX7bJHEA6QRGM1NysUnl/R4cxpc2IG
YxxPZFAdqUNop9SVCu3cyVnOB/3Txo2+EQHphJ5/xReFCqP/7Ekzjfon/QwZ9JUdFmYOaq1JlJhl
8GL0HuEHsqAFESZMr8QYDtdGAX3p67qrpH9cmtwB3swoeqKOd674xln5oEPlpeinOmDOrMsMvYbg
WU9kr+zar/dBMB2J4e3lBIjVGmpvKV+qEQPxj2YKHgx4bTNCzgjfq0bbfsx4OQmcBmOn6MlDT4wA
blqKKW7BkTP3iUbtEYSaZMacC025Qg4Pmw4hPHfdV6abVX6Ms8P0k8TpMirwKeGYUUyMELMps0KD
tXCacaPu/up46F7Q0VSkMRBYIXCUm+8JaaRzcENDc9k6cFjErtyaUZXPYyCF2DcHfDEOEI2Vkrnd
j4o/j5ZajMlttsWJqfio98/lEhTDWGT/v+GSwrPKV+JdJomCA0OuCNw4RwVRR/eY1zv+dqUEGZbF
Yndqp53Gwy8WCuKw8C5EKaA0NHBaIkFnVguwDb/SFGyd+ZcEjheIGukUiYBuKFMJd/iwCkG345bf
CJCVBgI6blxM/pyWLsy4M/tZ1LhV3wVhBHNn8sryWTmthXVxC9wEBafDV6QKDgauVEfTJyKaaxGj
2xhKd2xet/nBflSkqtlNLcLxDatsSDxQIr2EKXo9wvag4Web7jd54wBi7T8aiACfiLqR/r2+vkgW
P7rLDoOWpXRmvFBRCEMlwhXJVw5PIAjBcEGkXZAQYB8pNCqWLWoxiMoG9A1OvBz72HZI9zSIDSug
vT8MMgKj+kWWzfwymTM8vZYn+Xfga+GT/dGUMuLL3m43+iUcB6zBdunI3mcPl7cF8stXlAi1/pwj
9wK5rCRT6NTPlL/Ngvl1NMjakhHgYaiF1MVFYROk5N08dNKP5CYfS9sPYf+HURkYT33sTDOnUeJP
iyQ2ZcEJcQY+/FwyoeZTOEgH7JhC+vMPnn5XbGMD2vr3WskgqPXQEmG8aINMCLTw8FaJxEUMMCKS
Zg109AEukW16WCHF8yXJ3fB8qhObVlT46PaxvyZ7DLKX5x02Q04tOEWZdu1/H4UWXsiXrIlIXbiv
Rr1MamYNRyZ8XPrcdOdqMQyVU/xqrW+tei0QXDrBq8+Yu6PhfJtE/mpJpmSBKQlhSIu+HkY6bhnm
6JywAkyjVgSq122f1scGgyUrcS00P2Ec4bV7PG0BCIRMOPWwSeP2wQ4shKCXSdtAZByOk5qIrFFZ
jtVLTRQbkXizDfLQ4zmnpmnPOqK7MP4zK5FPoeFOFOwmoDmwI+I83AysAligtRVaAErizLzkcExu
Lp+Hmfn4h1GNE/DzrU4TGu8tGaV3rjxk6pmlfmXjhmuckm2l/oLcdDMFohSE1OoqPJJNehV81B+s
zkOin2H/+tIzyyz4eMKm037uNKToV+HXfusz4mnLfg7CxHCbedTk3pZ7SB6T4/c4c8k+fIW3AUNG
Gyu3rv7mrlMfi2trnpCPeW2Zn1S9RdS+dOZ7n35W/hDllwy1tb7oUU1HBLXzYqF7f802TJasH+Z6
eLo0+DbCI7w2gqyICV36JBonK03EFSy+mtgz6BLP+XrcSlL3RBaQqxPioXnd8mVk3DwiKs8LNYDV
tjba/asik7rboJwB2a7N0k8H9DdfrMfFEomCylFPnPyIOWwx+Dwm5jelldBy/fhdPdOytKbMp+wL
pxC444E4taKWzp+SGhbIUj/0wONGGdg0rz0MJ6x/6nr3MADxe/3V9IH6RgDpR+Wkz0KwEWznvCgW
Qjpk/wvEVxEn1dYKu+q6YHUb5waQ0OxdRT4zWjYOV8Tnr3X4QaEVK/khYzmjeE4FRRDNW47Yo+5S
uhvIcJFczEimIksw+WyOVU70XdskUzhoKnBY0wWj6q27/dm7/dTQiI5Uxw/8HILAGOBnvCxbhOk2
PW3ZMlp9l3YwhO5h5P8PouCz5EC/uUMMe4qW7J4f8O/PvuXIR6X/QMNxWD/lNTPjN9RLn8mFg1eT
x0OeRCf2OZz7GmX6NKxcpNpw1MOSRggzL2TekRQfHT18g9ab9/q6LQkjnQ8/DNA/5I7X35uZEypv
wlXTqTiq+kX/QCTzbzhIPKkWz3wzVsEUY3XWmmisCUTnHBVqkYXYH+rLYUjCNG7Y7f6Q9M4tmXdb
3NDtQPOrgI/jG8tBXdAvOQoo6VrU7zKw+Forxhww4sRboMjvkN4qBmddeOgB8l3XLTmR4C2MMFLS
WSSKCWeqlLdIW+dPkJWKyBzyMb37zYGsSi4qk8KtxvEOkzOXW47M9TFqLtrDPdKnHgIFNZh3iGoa
l9/1VTOpljk4ZS1dy7piSWNiZlaJtsYDfhaw+HPpXp3ztdDsh8OC+SeOwWE7/tIC9t4NsFBDwBhN
HlM4EUirYJFIgUZ0HoMCwtdurMMpvRag8ahsseNGnPPM+IoFzn/i67x3Wmi1r3d+TXinhPswt9TW
/aEFT+7oaA2xGH4UkqjCQdt5Oh5ttf3hNX2CyiJjGl0+KuQq7tC8PnzBenEnq14MMB1CCWpQef/F
UvBItSynyw7Uj6+hSthpWWrc5tx9if5ZsjdTyuyZb4Vlp8cLW6VlsbxikyXg6PeTBi2AkhxvAgb3
zEA5fkLbehGC8GgVYu1xvHVw/bJX8PbayuAzCCy0I8dkHQ/o3oyC3ryJF9BC85PBjwVnfCfl6m77
lQKgsteZG+Xqi74U8i+V/FQqn93KZoYTznHyGvmilKhIdbXIX34JFw2PykoasWkfhAamkf9LEQEJ
AN1SLg29c0z7GjvufZm7sGCsucQ1ngoObW5n/pdVCH2TwUXQk2aiJZNT8K4yV1kStGXSAtJ1AEOB
dCzj1E4tMoBX2uVxAIMMQaPua3OhG0jYyXEzBivshYdkfNoXSFjo29NDLhRFp4v+PnTo0BSZPBzc
ESDKeRJb1+7UBObMOoD0fAWn0DN2iVDyWzhuVIH37kseL15hJkXC7I1QRqSWJiLNezNQ9jNKlq2b
+xP2wpcJxgbuSdkGDL2fFi3ShvGL8wBYIFilZWzn7//pE6Rs14qLO/yP7kmHEhoLAW47xdL9gRAv
blAWD8GDXEAnkMQsSP4w551HfWzacoUA0lg6cfOjtAxvQLyLScay9X0YmSVvxukOeTmk75ku+g8k
W8L1dWdlMFWkWOxSC7A9fGNscdgSpViegNyOP7oISoA5Cyls/z8n5snb9ORzw7VDyCbhhSgjmg3V
Z18pAIkkwl2o8yiZPFwuY3XSpeMrsm8FpQ2WMk2dCQHrFCzoJ+TvJn2YyLma/0w4yu3c4g6gf+lp
j9UyBhyoM5513W9QWe53p26Cqi01+mlUnmCZqQHWDLgqNCkbx6RxXl2sPL1fFn9Ymp21CoGNv5L6
aiyjBUbPAecOKMVGgcEMHDsyilk93UIhATUAk1XbUgU1uCDU5mjxa/n+eHiRppU0k+CwQ3kODsEp
CezWST/yh1ZgNC47K5D/eGlfLVA+3ZhVFMqopD9tKAlJrvD2ylNHputgGFMa44T0c01AvC5tYncs
/C5UoFky9gYfhZ+9Ya3bWGdqUg+Gxa8hI8g5iO+Z4Hsc+Cchy1eoqGlRom2bdhoKIwjy6TGB2Nf+
7m96i+GobZ3Y1A7ZyP3k1K4UanHY45mcJggxNL0DKzWHhJsDkp9npzcQ46BPZA9VkCqrG/eMG8Ij
8+ttjQanv8UmUS0mc/znIah+0aomiNc5k3y+Ylj3eXzYfJ/n68wIOzKUrox3tk2tKQCaY3dAIgoC
Db43aLgkdY/8U9E9ZLT6BUGo8yrwzilorDe8spxzcnNedvmQtrLLdZo8KrG/ohbqyXHPwhhumDMv
6EjnWhTkPxDfJe2o5XfG+R0tVhikX+UdA3JeaMU3z22YXX+Ne8glhNAxsH2tSoOVW7a9pXb6OjyR
EfpZXZRY4E66Q1EJtvwY0DMTzKPQjhkht4wHxzlgqnjArC2Fg4tTUBUczvlcBE+OSL3HsHGxJb3e
TnP2Z5XCe4bULWt+G9TzGiDbK1jBSNOpFDZWRJPu0Nu1bWlrPp2qdtDc7R5n37IYUU3ddYuMfnd5
QwLfg/0zBIRQ5rlvPm1ByKZpjovSs0DtEAiPNStJQdUXtG2Pa+mwPLY7hCkHHM0uEjZLKyPTW10+
coaIHUbuRUSzp1Ta83V9vdMArLFzhoG1SUgjge9bHV4iqzv4e4svacNiBjRN2njy3jaq6WbepcJz
3fbt7cijCwKv6g3QhmbqiBnL5fkHEjziIK/RQ49lI7fOK0kTGNcyDlWyrRJCeD/CEzDoqydObILC
ahS8j1p7hTPLaD2yXHIMVmpbZmYHnu34uoZnRXIGtsCoJisfhAxjk2XQtQl/c/+m5Xt6oqr7lLcL
ENLKnYqwrUm/a6c0YftUKespZupapBcKenvR3HGwiV0bsCfh3BG8vV75ReqFkrp5wNz25++ARm2F
iuWG/UKhjvd2zQ2JgydPe8W3C5lzCRlhPrKRjNSKihM0UoKVvDwc76Q0T0dmN+n9941eY9HeqbDv
WQWiFhy0k6eNPIhhhlDOBRBXxwSahgK9PnhFyzDRxBIR7BJ/91Cj3e4jvbcbTCN8eQPmFXu8oZg2
oB4R5blLw+15Q7eiIGZn1UtFd+MwHmG2Q3EZwPOJRsfIhldGbJvJGs1no6wEpqdVFt4I1BJ2rKHg
h8UOhfZOSAvwSQY6CtYJ1v38crWf1harc9H+U5SOwNDlRovMDe3Xu5DUm3SzuuzTSBNE49nbFJTH
/2xn6KgGxoecJ7ild3XXzP94Jenk7nTWIwG6ndu91qApQDq15S6M6BPnGsUcke4lyo+RVGy0Nw4m
q1KwaRQ/r1ijzpE51ws6/V9NKso4wX+Vw8jDrhdE9BDVifCnOuBsSfVmEetS1kCpOnbSrfnhbwPp
UOU+Gu/2afsxlOEJ2+TH+n9YntVeMb0fpgqDStLhXCAdJTZFdCVttuZx/iHmo1fz7jZvmid9di3i
QxGjqSw1/vNPo33Ch6ws2p+LYFATIjcYh7HXYr+FCjsfGRD7xOUpm0hHH47c45UEpNOCB/Dg6NnQ
JhlleiDN+UZrGtZVoRljFBx9XAqRwIlpaX6tPfJYUr6b9dsDwTZ3xB2PFWemVC/cvWVNKrW5+2sG
XjrZ0ZZQOJtX90FjeWI5rCEKHbLNfrec+JMwbxGw0NcGT1u59olwGv+d7BM1sUU96GzOd1uCIsH6
bb7Uv527ltR7MHZkI0IHUYrs1L2Ju10J33GhkYoJB2m/el6lCI8SqBiLpOnXZyIk912jF9C+LN0b
3XY2bgDBm6a/n7Ah/3sWOWCf7NsvynV5c+ywK0rshzWSHItThNcDKvqqVv3bso6U+DgyfAIPtlB8
k3nzrN9/4EIan6FiJWeiDhLdvmydemwGub+S8zYouMQttKInzG5IqTwgLZ0jWluDy8bNVqhlispA
49MBrjVyYtgMWR8/+RwKZihbBvFHRzMICUo/m1UW6CT1GZn9vZa6faGe1gGuxtgR+92fXBUI5jm2
ELVypyfdIEjAAqLTwpxgq8MkvR/mJ0ZATnx3t76XY4aw4kseqk7HhwkFq+DC6S1TCLsnmntWdIWC
l4otgIjQ3A1OXpG7Oau4cWxhELWj5HZvjpDi19OrghTOh39ik7jb0mu6w6xyH2sKzHMoZ8ce2qpS
jCsZFqLrXHIPbLZmE/3ZwleCHnQwBkFzbZKM49kggV+0ByJeOjmFCb2ZHgmgZ1QtPzIGSD8EPgYR
8cQeBi5fO4ZVy+GN2Z6oQ/hUuLmqVEc37MtlJHLq4P2SA2Vwy68w0y9G7ELnRagxBfQgolPw3QTc
5yqvyfGeiYlKW9ulvAPSQ+m4v3pC9UMz5EDSvPr13eUrv4cwq0bn9d5roJmAxOFhOm/LaY770rqN
k8jGOiwUFdRBnBsIBLB/oRz3RT8zi3Ck96LmacsHXbWJbd17PgfbQhsdT16mK6+F8rz3tgK2M7DH
YP46THIptSzhNpFvg/DnFZG0ghYgLIw8idS3i7NXyTDA/ATB+gBylANAJAw+7XopY3Xc5ZpM/1JK
CzlYX4wz5Lgu00KOJgZroKR7jJawLwihiK6krHd0KWo4640p12SFluFyAi3fO/NwOEJyF1XLt93T
PNNDwfj+g0MFr21UsYBhh/03+/50kAV4mpL8Z+qo1ITAsv+YjYkEfaAo7/0Gk+JVnhhAd07QMXdc
CrdtyU0D176aCf3gNNOMWne5o+XYrJuWX1Ato6eJB+R2gwIdmOX6l3lHHcuLUMP6Wcb7MG55bsBE
6NiuMq0EXIZVWiXMB30F4u6SlWa373QzQd75hak5c9MoGwAxA1ln+dnuLKMzRqcJVp0wsEy3g6a/
MszDAIIW8U4JIhWvdbXodw/eWeBc0juyKjoE1tJN9B5ez67HzsxE/s4+I12vTRRZPvM5k+gz1zY/
uQoilrCbAertKQKFyDvcxX4BhweaJZxfDec9AKousnnfS16XO1Z9TamEaWXT1wT5UK9BRbok19r/
svkE8bHrL0fqESGedgFDEwGSYG8UpjSl87S2GI0lpzNGbpgwa/8P3rNJzM66IbGXCxPPHieipXw2
f5XZMlrZlgULwOFzLLqw0pHXs6xyfrdoGbHRuwg3qehoGY2lCaHx+HV27VqwZ+f7+J2vX6Jqu2q2
agJQKByrff1kkUzBxq+ATaMI+BApcMiD8SAUl0XTEMkJozAoTs3wAkAT9jA1LzpJ1CBTzqCzP2S/
14F6gaTBbiGMg1dVxnAwJR274US11D1H+kMcxxoCNLGtjapt9iiZ73lSJIRXYWtpz1Ev57avQFvL
kPwsWjfxHRJhmA2kjcfCMT2IJdjqhR0Gt43qYUf3rdOhYSR8dHyw1qaHSZKhse12aRoukfbpWOrw
rNrks5HlgRXyWP6sek4ISYxnXIIXL0hKhShnd8bc3VpzgwvC1o2wLrY1YVuDu2/2p9ZzatVPAI4W
aD8YbNSuUrMQAVmwUQpxDHo3YwZp9bvo4qbMhTLHAdtOsBne6+A0Ny14dLiqunM945HwUz9NTIJh
XXa+r5aqGOG9Yxz8lNDsnu0bk4LM7wAKWJCINP4/3ckgPpVs9JCiYRHRSlIZgKP+dzpj7lovuQLN
TK91OOInFXuTv1Npr1FnVgySDF4YIrhp3YO4HXhowcSj/TlcnWhf0YSUpzLXF1DHURL/8DPvz/Pk
tvqGsnkbir3gOirRvQPbLddzPgbHXhd25Bp6ARMnL30JvyHs3OHecsy+TIhmOovSb2nkUAEZKJTs
aLlmIzhook1pVKZvzHd7MEOE3u3WP9G4erzeUtJ+f5tJAUWBETXlv2jtiuDrsFIuhQc2stO0fpQR
ni+jen76flW9sVx2Oudhc2COyH5CTIp0Hno5jLRzXthWa2paEHMhTO/MmkuunOhF0xdT9gmJ+Yhe
/gndDzNm/LvCEN6Z031feZfDK39XpCzkuGxcs9FTiSmLjYuivVAbONevb58Z7CQ0gdgm2M92KJfI
qOd7FKdYnPpSvm6Fc37xEjpug6APLS14TLOF2cc5tuQzWUDNsBTwMNXopSk1Iam1dMDRYCl7EmEZ
4Hf2AqJ0prCG0hY1Uq4OnuRjE7rqbPWjbZN4p5TDoiQ9X5us/LUlW5o8IbwGLsm9GpBGan+tDiBf
pclO8kZMxx94mgBdYvS3PiAjBcktqrAvLXIpnIhs1np0fIsvCNMyGHripFWb8alOWAnSXfEYWVcQ
i6GbpuuJbV2BxSCXKtBg188MnzHVnnAG3RMG4Czr+dQETXNqQ1F8QWhoZWvGwAA1lu2d88E4KOV1
xFofNdsvgJAUvXZDZzEKpAApSxONPOx/na8t4cGzMzZgk7qf93lD2jO2Ozwzd1F6Xv4dQFmb/PC5
3HsH1ar5m4lPY6KX+C/sVBMPsvB1VQVXspOjUBz1sIqQ+ARXwIZNf56mlJ6u3gUjm0Rk22tgXhsr
TjwHFX/Y3yJnP5LsOhAflP/ikYLC1urk+t2Cqhx3dDtcx58ffXIIwoHygYkqlrmvTIH+z85QI/23
0AJGDtcC5R8oC7J57gJo13qiOq/8HqwEpsOR8FPerEKHs2n9QS5iWC8QfjAHMyEi3GluH6pMsJJl
WXXVvSqbCB/57MXB8Us8ydeYTm6K1H/jzsJLutpkgy36hCCEsQ8fS9zcZeBumsQ1fzlAnHwzurNF
63xH2lixYRjF/7dLmeDODQED/Edprll9noyV/HIzen+fxtAamrTApeaAqQYmdObBrlV6/x1su83z
lwtEXkp+G0Q+dmn8gobKNBBXR4P4l7GKm+7Oz/P4urMpaTqjaB1fQaQH2Wfg3xuEgmmYBjCIABxU
5FW1NWN/OrZLm7BlHjE+FjEM+i/bw72t66HiSLD3nskRTp2N9VFYwtFiGWToJBWVo+TLndpxuVZ6
wINI1ZbLz9OhbHkuVPIoIm0YlF6onIlWLpt9fpEj1fmWMFNItkpVF8N9Op749XQR8I9TXVSv4b4x
vxDkrGeLw3kZsDrhYQ16RV/WpWlkLumVoUszlIMCG48nDSjpHnfVnvA+Hy80zAAhJwcsizuKSr+t
T7VULROK7BDJ/O0xtjYVXZ16Ckxf+arBh6GP67nAWLff/rpraQj1cUideteDL6Ku5bOLRml3nt8C
KTl/s52nlBTKGQZhTAMX0qMfztrD5ZtrjSmwaLo1P1q5R5ttItKuf0JsSUiWizrDzrzSzO9QbCHR
tt2B0bFAnAQIWqIRXdxJZ4xS+njf7jOvjVlZ5lz7SRzzOkVZzaRGh5NuyWydr14YUWmY5e1EfwQN
CzcftPSnWdv3cjMlpM8bYVL45rVJBVhzX6lwUhXYYmXYLpcxPGWTftNeqVet5xEO6/2E4AkhsdiG
p0688s/hTSXG8PrCguhtQuF8nqHDKWdbTbCnH4r6kWKogseHDe5LdY9NzbBdLvDJHeTVxLtKWXZG
sU33UjF6cIJrJl+tK8nD0TpuNPABRZaoOonwaLAfCaJW9PpLool5CRS2z2MBCsN48o6qaB9GB/i0
Z44FNtRAF/NT730JCAddtiQ5AgmCWRr+vO+539Y+tyFaXVm6sGP4ieykO96T/hUSy/zDOR+2dT04
BEwtcMjzTD8XVg8xJKYFjOMMYIRRgdMsnxetf7TQ2c+nwb6FIMJGu/XWjNCebbxcuqy0jzsBqmHi
eQiwuwHKcCpA0wHSK6eRZSwLbkEgvNjA9WjfY02/uSLDQVYZXN64CTnPMjAigUA8HiFLdE2Pvjg2
K5WstVeFC/VP/IMYaPx1jV2PCwLPO1H3QYzq3h++/uARcqxchyOhW8CgnELapIw6Le3O5WGYJeN7
oikK/H/voSpHq0o/JrfhYkDqqbGYAybiNPu1/WWaPxeE65sqclhDSLpLrmYuAAj7RRzvHnfYSUyS
yZEcACduoATLNtut+fsJuKWhcWRWehF8FM1KTtBrHqUAR37wRtccVYY3kKzYwCh33D3Q3+bPrK4d
8Kxn9EIyBU5NNrY4f2UBltpRgUAbMX0jqrs/ovyb8s3i8AKZRMm55jI8mcxS/3nbqhfJa20AC+m5
YT9Q2hpSOxHCOzYk2KkP3xY8NDPGatcv8oRQjZqa5CyjDwWF2YpZ0RuYbupLpTBr0ROAbk//tThz
6slGFW01ip91NiweULF/C+a7haCawauPLqpdlUH+qjT9qbd0MbHVZxjGC3TDJ4iAi5ZMUU6r0KGt
CiVNwhUHI/CYJBrDc9/Y65oMkaHFjrp5AF/EfSti6I1UYYXX7F0Yx2K5ffhIa+OqxbARymVdiFCh
IlT+rzaiwarGAE4rTDv/sJ+zo71we9DXwiKHtGAs0OxX57jgWWy+UZ7Su55i4r5OOTgjvfNGeLB7
DAoDKaUVFhB3QT/SGAXs8XhIz0yc+V3wlNCHlL0FENKAq1m9dJjJiSlGH9LMgIGuF9ECPZItdqpg
n6m+sAYUZ6AUXw8s+YSlZkxCjmKEBOyCCp0mN7ysDgCdpsNrnYyBFIMD+N9+8tSwAZFkQvzPTUcF
Twp8P7te5kujWokIu7ByeiEfDwP0Lzn3Di3Pckk1/VRCHp8RRZUxkNs6SYX3v/03Y3tolLH7szaL
yfjx5Gv4JSY8d8oKOKsOVNqJWnCjpxtO5d5ETjg9wbh6X1xGJgEBDWl4il7SdMakjlrQGKr79MFM
nLMsAQcFQA9zyplKYNqlGKH5MnMG3n7t3kyOgA8v6QGhfQYSwSGW327FZ3gAL9lCTBVCgycAQy3g
t+19Gdei3lHKvoSKX5vMaawvGB/f+KXvgFfSSOSNBH47+DGQfG255/4AIzLuW3PEw0vsPn/+JhIs
jrpDXgLTFOYbIoOzh04zrp8Ql/YSvUipAOjsUG+Z6VAFR6SyonY5m+nUnLq9P8n5rqvjoVLZCO0A
0ngVVDUsNNCspppTFsShqsVYl1GT6Z1XYCqqLTjtYkVZ/TVysmX4pLmV7LOXMRmQbJpCnVKlNyTA
blVxNso+LBlCdqr2isvgGvEXY7b20XF4ehIPj5BZVjpVZoEoaSRh5OiLlYhJ1hUEUa5mRUzGHR2z
7c9A3wrAgPmJYFVup6CXT2kjOQWUsBC/cW6853J30Xk1E4UXURAptYiU2gY+4mne87nfF1bVQUWL
M6tR4+QKTF1UQBohBbtMUQOVUtkQRyNdHFpGRItFeIO2ngehWt3iLmUrksbz0jqqpoN1F+BgsaUL
P6eLBgGnvYGFsJWGQe/PSPwnBoF7nqCRcxZ2dap87YJiiWN59Kd8rs8r+eDgWv/2RXehU+HpBw5o
uZPudGqB89iZjTKk+2ePC+Lx1y+z6Lhb0tg+l1ZKXKUyyNcJLWxKOKdiH1cUeZ/6Uet9AbbQTJ4m
CsmZULqpZf0sIBag1cZHooIPUkJ8/ISJz1dntNcmbjlwp1BUpbpV6oi6G2ud/7izYDZVyqS7Sr14
NewAO2oLHH+HbvwoHBmFj1H9ukUl/fwFE35W7AXAwL1QL47tu8ZyKS8bua5K6hCNFPfU3RHG+Aio
AD5juo+LY43uMcTCT6720QzxnSRgqt2g0cx1eUInh4lh2M2Z9gzrLi5ch+K3x05gv3P5fLLp0EBz
AzgoATjUhhlQH6GSzVpRTI5DwJsn2mLPGLl4pEvChh4p0m3z1Chv7vmVwWtGHUfm/wY3MD+rWzHi
GeE5TgUO7U2Gxd0RKqF8PnAqqT+kSKfGF2xA6OYDBRPHHtkPehfFPlAq09nAMRHNUHktNypepL9j
SECOFotJDvP90axRTvgQbRoZXky7/kyF55unVbPsMIZk+4KzUKfKIcFUib0BocN/Hn5MyUjHo9A/
cuBidqrbco7fXj2NiVzSabIjtLFNlQEAOxEJjT6VCecx0vA/BEKWcZYzDr9vuChEOuQOnAL0w9Bi
juEtXdJZfQm/Wp9/E4DDZqjS4+1ExO8CakhW4qYoeNYYodNeO2qPteR4iEtOp0DtqbcGZcJPSXlQ
JyF1PFQuX9vR7vL9SlMpI1tssayLO0GwsPsH8JCtfd/xCR657ig/K4Ni8KGDJJdDP3JBscd2hren
EDec6yDYReqvfC0Rb5vU6x/qtY5/AWbtlYjenHaglm0p9q1kkMXJWqxju4i5JekxGUP5GcdBb2kA
bmxhers39c/qPXTNlfV3FXthzE74qUZykk+gbm0oCtWiifGxngeFXgfZ8Xaa/3sWwHU3p+DMiADN
zTCXxRlugaYffcz0kcKfpFwpQcdLlbFEwLIDzzpQC3wNoLHNaoJIjI7v4G9Wp3Htgf1QEuVwtDlS
coS4MDwOrcfxxKNxL+EVKJbYp7PT9cfr0Wrp+LMcvKSl3wJ5V9uRpOUYiYCpPOGvhrwzUCAgBrMf
/V9/1mY//be44M+8GaG2XU7DLfCE5yHmxSmyz3FTR3RbGROBqK8KMMPe46MdBgM3lXflYUrKTitP
OXcAwNbsrfP2CnWWsm2NlQrHximV3b/LF45zw5uEyerGeZfy1kwImbw+hgF5tcPVHv1So9dsrhGS
EbIe4ozXCdmnmw1eLYpjFzIh0Ano7e3MNbe6TlJzqz+2vm5DtTSgokPDYqzdU7txWAyMgOypsjHg
HVU/lltDeTr6HpxS/geapLxEIzseku65W+SST1wV/4G+Stxqdgu2/F0NZDbfb6Ev0XYgZGwTmAeG
nn9lQMGa6iAsXdEfNm+3HfTrlwtnDxOBYAPLkGjpIjCTJeObuPkkJCdXqrrHZ3vZ4NqHn6E99riF
i39euu2uSX4VKE+90XFxMwzEpJ3TsDEk8HiKAZ9txcQ3P4mZL5kALqfiylQbvKPoGIESTXvaUSLb
//5JCJlgJ/nAAdUBJdYtsuEtzfQVzw+y6cJ8bLKv6ZqBxgSUbmHi/KHygBD1gszaYd55PqdSv+Ox
lLlUKGuHja2Zj7dxPqIIEH5dJ4jSIE3Td9Mru9F0z7alHqHyw+e0elhtPjs6RW7uvsVs0pxCOE8d
GKehQ/q4GEnd6IXpo4ywta4kIems4YsH4AG8PUuHL/J4fyv6+uNLb6OQkl24b/1hibw8c6lps2/j
hH3OX+V9/4rv5TcfZiWNIQBWMUcZG4ZZpYWKb/YKdV8PKjhcPtS3Fdrh5Rrfu4iUPA6khINijmoL
TFuDiZ1bgMciFTUmqhmoOlJDwFU/GPnqLpcciFzO7YYHUXkvnFiWBLHte5ltIncMmQSnV8/TeDh7
GAUbIwXa6/tSPoPXK1js4eOVL5gCYSnUDEzOEGTSahuUYpzblUt7Mc7kr4J5Gx3SVrwexHjoTjLN
fNf6Sz2DTvW9p0vTG+QsSlF5bzG9SF8+/NOU1VLfJBN+GebhBBKRLE/tv6dUymZQclf0BvjNvQxK
m7MR420WsAa/JLh//6UZbjbe4zRFLlMLqBQTgalW3tJew5qhmwHWyzJI5MnMQAlrhuU2EKZgZrRL
m9cg+UBHv8vbqYmNFkN7pVgsxmCGcLbCr0onqTgPN7mNiGk1GQiBZ/dblkpjKGpkazbFoN5qmpOW
8+CyOwk7Q6j2NWnMczS+4Ug65reGujx1d9qydEeIMZWN9I0zsHnVpJt75kHhvLSVOe5uE/Pf2h8h
Fg4KMTJgdVOHgjRJXG9kxiRJMSZKTQkP5onGeLB4x23k/JpWC3U5fn6nLcvHlE7LuxJ94ny7OLnR
2Zxo9/hT+rhja2nJwFbYlDltFn8KC/MmNpdP/HZA42PhAp0yGJz39e/y9rX7+l6pbe0vJ26zNknH
8Jlq/kU1eVW5XseCY/FipCFMbURHDA/oQwtgB5A7Mjs2x4KTVxtK6EBKcCB5INJngFJydzU2wajQ
+2MHMx8TLf2GtroKBp/pX0JbBerwKmoqANSrDwPY+/eWHi2M1iikeJBQubxRWWfC/rh0ShvUTiI7
g/w4BiphVjiOOSWfqOa1x45v27BiMT9gKFHDdqbpEiHWZhE4xt3zRZ1I3zE2OTA6bpwAoDxt2QVZ
pXkO8XWmsL6Sj3xINsYKC+16Q+BM4gZaixcGWEEA5OVuMY0jNkOsvWcx9AyBo/jHNBedcn8MuE/Y
R0lHjGbbE8vC7c1Zr51Q2VTH2bdZ1x1A8Pk59v03Vik/YlsM4ABc7REo2oJLdqXDkcVL1PVgYQpY
cmNArdjlkJCYNqe5i/setvbPhwNZhbjcGrX1bIIzDFtaq4UbgRgtzTm6Gs3/PD8+IfWi0DZX0PO3
0et4+g5Dv0g1DbuduuyQ/BN/jawLXuYEU9oc+sbWs4t2DzL9J+BwaXsZY5xbnNs6WU0TKfvdKums
CVr/DxCWBVmkQUvr1aENPasYr0oZCtiA70da+892pGMTAQYyRAtGKrlKifXA0PynDGqZ9iNTCzDt
dUkLoiASbF2edybGDAkAvY+vChUefpnUFclHuKJQXIihMgZ7qh3L9oariCAKha4y2KR7NxvUkq/w
3aUYePWrkM7nPJ68u027awyLoSV13tIf0mFgawJwcDKmWlG0hhTXVApShkzv9mg5DaxcZGpQJl45
lzdshXBC50DYaE4YKn9vpx06h/oHiI0jp1dBP9R/zWrMaKS5ItbigI3zsxNhWA28buUhozrenx6e
TlCTgGbHFOyEmwlUP03hJExdwFNmLn8OXxjUlGf7T/at5mRomB/P/k2o9py1IdXrCXEmB1s/8bJK
rHBkGi/NMSvSFguzhF5+INzLkRpIgS78M5udF+gXsK6BO4USaXMqfhAfwvDmOgOIX6IPMjX+yzrv
zvnzPzemP9yvKpTwlAmePA8JZUTp71yqRRTBdovkcuygLduC48gQ2tOMiMHtLxa61S12WDQB1H7y
QnYkPcZgVGLOu3bTxXx4lcPgWTz4xqOvXwE7+brPr/L7+FJ86j9qL3FNlft1ARr2VJ2vF9cRbf/A
nObCzcYp17LOpmLyBo7KPjBtHNPmKJQdXyZwhAkS+PaIIxfKgmoSccOnixilqSUGk++4yVi2RHib
cP40CBI+8zgp2u8GMADM26cJYtuwofkszYXnMF52bsSFyhdaGTivLEz2diI02vVaKEIRSXyuIEJ9
QUPTsF5GdgOe37S5ZBxKaU12+Bwzhsr17Q7JMFTIggIrl0jY9gFvyHlmJl1WsxGlm6K+UyEXKpYZ
CgV/C5ECYQtsiOpx5GFBgF9FRgITWOdx5uiEwiB6/d1LD1gZP9Hs4z+sDzBDUSQ2oz99mCavP7ek
JvpaMkpwA5I8yO5GxDjJXiouJBCh4BobVbPshGaHxjQ9Po+46UZ1OSmN8FPoWk6ANfSmMbVOAmfB
nYUys41ovA23PE+NluiBZovkX8mX8Qm/ooIb0JhfU2VcUvVi9BnddNkVc5jFuyu2qzCFobDhvDoS
uXQJO/I7Vuuv8JM1opIQBJby7vyS0uF1fWpVMQ36hrHSK4e5ujufT/PQMxolxQkxo0T723CtXWAc
qDeOU3MXI7O0gv6EZ9kPcYmYwv5qsPfj27oT4E88NQb7nCxC43V4l2atvLLb4NajUXBMxpBM7yce
l3G2qtaGE0ep58/I7M3Tqjexc8VFXySOxbxxCMR/UnTEyMIAFwnGQpMgkpqzl66sA/eHUqxDTueb
1Fe76b+8/x7d3ty2vwW7gNZmTYqkU3GVbvUW+tcKkC94dsEP3Io0Y0ghLzPqY0ej29zRxZaRX2+r
84b/IUXS3aMvRLzCtMnmoNmpFt2ayU8kNKmcDbKd8e8XVrW6wwJgZsXCT1LDcSSCmiAdA7WMpA8V
C8oIVsODfTS5Ar3WMV7fOqJTnJzJZdTquZprg1b5mNNcM+TC9wX/A1vXHb2rZoqqDOAgD9HnbeUP
IDYZ3inFtpYu8hwjEvdkFUowW7mgpsvZIH0WgqTnfbV33k0h4BthpjUlwsPdrVkTyXuxIT7mQk0k
qV9yh6yUbZwfNWmHJwpnrCD3uBWhQBRezjP3m7mIFbrxqRc8HY9n7Y15upc9v4tkm8sICewGRed0
xs6csCNf8b/irWEeIL4dI0R7IY0GhS+Hnb1qcM/TRchv6sNrsdzp7YtPEaQNTDZHSTQXGbIRbaWd
bLwBfdeiNrQrzaZT6Vdh8M+1nV72zaemGYBxbrIfdFP6vt4oaQMi7DLwWLeYGeNktJaVJ9s+3jq7
QZYF8xRPxjbc340URMwsk8UaVuMLyiVXCViZ/UjYFVJXtI2659ueAu8fP7FJfGLU+u6sw7FCs/3n
cUMI+TD42XJg5kPskhLawJxRDQCM8uEFNayNYZvuEMKFSvqjap7kSUj1C6pkSPrA2BeIoDC4yZYi
vHAzYETNfueJSBYlhC7F9iWTRxN+8cSucFtg6qlJ/cjySyy8r1AIgLzh1AOVRAoVogWiOk+xtvPl
w1OLE7TnwPQiyqVgEnqW3aM9jIwUmw0yfT/xZ9ycNDTEZuF1IvOHAxvPVd+vYWbC9au1zATpvabj
jZ2d3OTZbcH/BCqdkuu5DlmUZkkg/0O+VVscACB5rDddRG7Wa1GjmO5No09IB31RpAlobZOk6Ilt
wLRPhyE9uPu6t1qrOaFbU4IVeypv26Z0Lpq+sSF2P6qwItCK5UitggzbfWIiHeoZ4C5vAtk7zut5
btHAl5Qz1/Pl2o97gbW9kjGu57995toldRootrw4xNwFZRUhArRqDdTDuios5ZdKMx5a3D2LfX7P
FRhtKgik455qyIDLbIksS+YulFEEMd7cGxsbmWnlJqMouxeLx5Y3hwfbLVugfHxC64Ed3Lt0CsUv
ZSrVOZDtWan3/KliS3CVGF32+O86PvQIPR7zekbS1QednJqQfAFAEXvXb+sudfnPP8YkhOWmltMm
FAQf7pRwIZuAebhz3M/F4fz5C6Z55jDIACd+FO0PPoaMnnTIknllhIzsy7xRqECU+1RcN/b1L5ET
fb4Ot36kSFdknYOmP4cQaGN1D4XWx2IvBu9DIOL84gjndE47dqmMMo2OJPNCwDMmUBn2Y279hM+7
H4oc53xlmdnSbrwx7ZYJD8TLA+fWjw0MKgn0MtRY+jg5JmDenSuopLpvylkE/aLwosbqQVHhNedI
+UqB7Swh7iz6BbY+tArGbsRU85p8zdTvgglbSQPSrRnnDJJGiPVoEKSFFPE3AV8RvvBlQGRxrxiI
/t9vVSEGU6gLCVUMMiNpMM8cKzUV/pLvek6tiOk5TUQdWtuOQg83Ia+1nmO+q0Phbd9I9HJXJ+KP
JDlPdAFoNjJ6cowpZjKqhdXNYTupmhLiy5VerR2chOJREO/EYxIQ3jb8Vw/JSLMYQUv4LTM2MajP
12MH5YACaDp5q1F30t27IHP8YXtPhX/qC9bbtYVjnSLmvXYe4nqF0u41EZ+czbfZomWAufiqyDoY
IaKaz95mpcHmFBuu7HObM4lwH2QKbIZhydP0C7U9zWq0jjAgAudnnce0Dgfas7KRm46CNhmZvzZn
V/Zv85fcHlhd6cNRJBQXM9qUcN3W4QESTJZYGejGK9j/kODtUjhQJziYJ4JG6pXyAGNCM42uiMXd
+w4yMMU0M3zwLJVGefURQnXlPbbWjoMdyccvo+I9CMsxMGhGd6yVaGDzRfMZpoXWfKEbMA3oF9OR
5Llv4q3aRGdnOElHWBcKHU65o57yDLC8vW/eEy+Ma361NOpJomYlARRodY2XZJnENDoR94IDqPU5
pE6tQ5XqMoPr2XkX7hT19/rymowdrcYVNCpIGItXltlZ+SdBkqjZIaK3gkbeBOipkzwa81+7zneb
qRjXtQSV3GHUDu044cHJzNSYTggx6ZVL60+uPssQuk3V8z0yYbywA1tTrZmOBBJ0WnlmgQ9k60f8
3e2Deq43l4qrumuakJNpAN99Tvs5KNRXamVcC+jhwhEqI8FBHRe1Mo+CkDhjxOUixNjn+1J3BB3q
kc1kp1Sa3yOJNAcsdENMqk36qeuoadZVcHTUZbpoUsfxnkRIU7PSIqrvQ5P7+Y5jaJgxAAm8/jsy
xODkzFoIL/98LRXolvXIp/ncMnRFNcLdsl0XOpYkj5uCh5hCLczb3SfuHA69ZDHSGZWKhJm1JFfW
GZ3VPutkAdtgkfhCTRj9CzJk0va18aC482TL864kXGCrSpWreUj8qd2CyoBDjqUh4P1k3DCoXr/b
A0FhiGMjFbEggzAi+3RZX/xRqW2dz2TGBJ0J5Ya561usggq9A0ITUf8gSaKRHhpIi8WaLG0Qsc3x
cVOkxDVZCYlZPgEBXbgrACefmJgoOSeI2E263IUonIohaEWkEk7uZ1qXxsbHVPlnlas+e0EsUtwV
bBXUmRbttqGUYR/OtU4vcOKU4RdVCSclYmWI4Go2KktAE//8rsipJtrxneafdKJdhGQzlUKENi7N
ng4b4ZWtRAyuMoy7zJ8PjmRjU09aL5eVLrKK1FQpecq66GdnQUxO6ANcR07U2j4PlAQSfHmg2xoo
8FkBcVWthWWRtmLDhkyRPDYF8hx8HeyUgxDcIMkXyeL2IF4IR0OxPnbzbMsOmAUlTNEkanTj9Qwr
jciGrsZSuk6safy3vkNw5s5d8KcG6BjvXBOTSm8ZWNsmUIAxKAVfXAH/PUDKEOt3pe52f8xJqYjD
cdMhwjBTn3UgmQQ5+aQfuyldzQZgCDOVDSTSowd+ft6qu6SvRMngPQeus7ZDlXagboSuIPXErIHQ
I8eu5hzxpFsHVEFfE5uqN1sonHcVTwRbBI5KyHDijpkGyxqwiLJmrVC9lbPXQV97uVhaFFDuXZFb
K3RyOkwB4rGusEVyTDkwimChYTI3BH6sEBe3TfW+pXkvcIgrwAil6bsm1l2g1+cy159SLpwoDFYO
g5xXHgeRIcrpT49sofPTsg/7y22xoWlREnH0xU2O37IOohGhDtqF9SZd2I/VbDS8znWTXP8zi+1a
7OJedrboTRND/kCCw6jdOzsukMxKn3Dw99py8kD6qCrlbV+V1AT580PEWib3d70f2/NGhdqh04c6
/DIRPc1NYSuNwFCmNXfFi+zkUtB6YFEyma9ue4QaY6GS9QWU6UUouwmnZuWYpjknHsYqrPWkVCX5
T4f00gkEylTdAezQKzoex227Y+Xtvf2FwJL3Egm4utaui5hd8RmszrJDdWyeU7Jo3pzxok1lamQ9
uDDwtx5jwmeiTQKApoXEAyR8ZgwRuWBgZntffaZXWnsLrS72Hws9Xz7OAw8btNK6HL59K0duNlNd
BuVmTC7F9Au3c1J+wYL2RdbRek0JAh+Yhg6nzsKCgERA+4VtKP2Tt1wbv8sC0LDRCKtNujn4jJrq
KVmqVykD1H38ykFBkwnMl1HowjdoUyc/MhI9XKpAge/lHnj2jWIC5h2p7J/Murpr/21nSodGs1Hw
gMX6NvVoSzvz/Z6Qe/n4irwHjevCeu+8Tn4QzBDBG7YU8n2GyXIt2mghMoUsiZg+DTa2xpFwF9kD
ceOHE19C2SabOovE77RLNluMgrUnadJPC/+BwST+hJha5YMt0jIx/qq5rOf2kNtPloObTUC1tFMs
08aEXXwYC7qsKPg1Bb6h20DXo4GIstTFODL1vdBNpfQVFezi6yjlehpZ00zgrgPPeAIBuqaUVTdI
2M73TsfomH5aKX5Ew5g6ph37lCs6GCw6fGsUqezSem6QT4fAA0HNRmuz5oZ/ZfxtGtkMF9yENOIw
XdiGvPtZtyCjkFDcNobBXsDNvrJUsqYECBHxMkqbxPrCnDO87gVL8rKkgFcIYxXQKtVq4IAdDYdT
/EX1L9On7Do+etmIPASglY+GrCv3W/b83qt/sWN1Yolxei7XXtBZCXPcmCamB9j/q6onSm3sakML
jkFzCzAvQSgfWSF4+ODDtv+wL4sgJqMfUa14e9OzQYzFT+U1ZF+53UkiCBTRE7ksfhb9B+6NxJGF
Pxxjxvi/WlvriZKwtMT02Uw3BGoI9YLVpAf6mjb1kOgHedtC3HF2rBr8roBS2BbLNi8mqe0BueKO
a2SE8i8NlmPd6BrGmvZQTOTaSEtJR++7dIFmJCTnT7AP4qXJAxgLzh6DefuUX0a894bpjkBEMY+f
7PUJJSlFvic/zXm3Vjb+RsrZTYO4gCNpSmqff2vsyCw6RutKEygmG3QOcUMVR6clMqE9Uklxp1P1
7KSyACfZd7cTgcskWrWaaOwn3VriVN/94xgHI0g0thk+543jF4n6uHHoi60HgT3fro5PSQnHbj0/
ySSnS19g6bZ9IidvSPVyFn6rE1TPnpM/YRzLxAlI9xJf/+aF1lbnrK88hsUSpcWDWo6xGcvfQ7QB
6/Q8Fwq5oRUO3ma6FEuRdAnEiHbkqP2IEKDt6XibW3nkw0JVFICsf/LLQiJemJxeCR769Z1OCxig
CjA7JRBdNAUO3quihYULWgR18pEt8b1Adldnn9VI8iq1sYFHRpWTXlk9sRHeGA6oSVDZ2G8YxsLh
xKfYjmQn2Ff+beWk5V1Ii/4Jg2gQvTaOBdmo3P6vS49iqqs5X2CuLqRpoAZK+GDGOnsfA/xC4sgD
tFGK9NC+0I8FF9fCxo9GLzrtYH/UWz67msyRU2HsUXppnQWMVFORBLUd9phwJzVw30nZEDaHUOIC
/Erup+jFObns2LfrxPvvjrMa9uT8rEFst3lq0ylVmZqQeUl2JRkK/7Xm8TDTSi++DlpzOGIAfEVr
j0CUOJPRYKNHJGh/Lu6gI3/UM4xaGV6vKyZP2veqFDCRcK2UPhBidAP466Fx7zykpX3sQusrmep2
LC7J7dnsZd8VqQ1cfWupnoi/x6N6vpNuz9RZLv129D232I7DpkHMVpxJepjeSDKQvB9hl9Du3F4g
NuGpJIumZiPyFqu2486bMmSJVcixNd7rHQSkftia+Xm/ZdNSrlxGly9ltPhFDGrDosQMnzwFkqRB
6ZD2Vf8N5gLeASv3dN1Ld6fBZ0HSJzglgm/70grMfgIyUAESupOJbMP0/HbdatA9PDuOR6z8nmFJ
7yHlou4MNOaqt76/5Cg2GnZIDOVRGILc02oYqSo6T8URxZbYWiINU7ghq8iaDdG6JK4ASekG+lYy
yFaKsZJxkBiWXi6Z3w5eTzvyJ6VJJdoxQWwiGuip9K4LFEntFT1iT5WHkibRjuP719KC1p3iSHYi
n4+MeJXjvQxq6OscQHg6wYtdex9/cVGXig+IDvxVbt9sDGPA2Vb5QGvdjOxWBRx2iW+h5FdiGPxv
UESJE0zfdLFiudK8j8P/lewe3coPOIbO3mme+AEdKUB3FnWt+suEtsQTBAfkOcZ8bzVPBikX5wCQ
TnJecJr9jgo/vj+RyWMgPnIvDEUDARo62GQ4dqmxdRNXIPW95pNAyLdzU5sbbKnqI+mizZtxpOOd
/rE7QZBCPXFnzQ0Ea7OKXgbFkzDZdbzeZf2/BgHL40Xl9e81rAl9cz8R4FH6EenEAPK5Z+7mn1ID
Xdp8sYeDHqBNMxEVExkmWwTVsp/OGYsx189yw9OJJkjjpYHNgRPpVfR4TJP2G6E81FdPKFrQ/WpB
9dMNH0jLum3LOEtDk4Jore8anNcClKxqL7KqHFYiXtSCfsl0UwlZpuCsY9bXj+i5eBCzBnNTK/sE
2/Dj8f7qPc7rYjyMozhvhdpjrYwpA9D4hMzr6qBuZn5KCdC7cnCDMoeelO5Y2lrGBxoPSq8wKeis
GuyQrZPFzBYQFM/NbPMv6BvIk8TvCeXIhsQXHQEnwkNVQdxHgn93RnCzokMzPyCvYZUhNThgIU4T
cPAfRTzTrfxdwjoeEriNPrNXFWL2bg0vb2me51jSzxulJ2y1kahlD1fep5oEnLLawB6XqJSWMHj4
hk/mpfMkLZGNyh+vavTEJvPJ+rpqxmJlm/iPrrLgVrNjxHBfohxta+JeGpYkM+k082jwQb74QYkj
8i6YfC+3gBTtMgjw34XZNH0ixJrRr+sXIhIWOJyJx3ZvBjJi6dPLCSmsSyhbEudixbckOiYuNyhc
gmipoAfSY5y8jjUyVLJMioBmYhven4tE0CDEnDCGpOc0xL6rYhkoms5RN3cFpbgpeulhgGgq2GyN
9SBnmMl6fD6rF8kfjnywL0Fl/40Gw2dlAwEP7CRlIujEBPbTY2lSeEUAVQnouq++8fopmqnyMxyu
3cS4+CpPj+hxXYK5I6FJm7mySTgU1fEgcTcXFqeVw3WGWefXo3LBRKW8RiE5SDQsQzpKI+/jTWYe
BsXyTXSVZpgZ4p2b8wRWYgD7XchOBgkmh+STzq5t7k1z2tqoLTczjyzpQL3Lu2qJ7EDgiKodNKnv
AflQNtYkIHG+Q/m30B94F9OhqVw3U0ITJEvzyceBSzXUdhwow8n7JeysTeDCUmXWsdjlbHQcQj0V
V/6NAlmisyepitrlfQ0ZQEKFa+wCHNLlR1bEhp0IMZXOiLAzYPdOklD3RBGy+tqGCMuqS2uS25sE
+TcvBAo/ph1gtSSH86MDm/CcqzKT+t3CohYq0loQkJlHrEqScagbuwPc02Bj6QaUj8aU3viAcScD
KTtK9t48+QKLELqSY2lCIIKBMW3tuoB0vQBk21/TG694kzIbPR0E2Qchx9Plufk7fBxkQVTC1Y1W
1g/4ixI6f+HBwc+ME0Rw8iuR2XrIHja4ZS2JxO581BU+rI/WnEKtSXEa42Ns6hqaVyFMKhvr+b40
ssz62AiQLIb3qZ88wcteu9E7FTR7kNLRASH3n4eEP/ju/7hiIpoQmDCVGWmgp4bjLDsgtQS+78Vu
zOJz+Ll3D65L0EtK8HDkbSajRoO+3luOb3iBIAqV1tW1h2W8iL5mc3wx92i3Ans6yf2tclhCqCup
qK5vjLZQmDxFlV8WUZbALbEPa2h+r1zWLc4wn4ibrAIAe9o4X58QyriOl2IDEY9AV4yUmjT/44Nv
qTkx7D2m5P12jLbfyJb77/YcPbmPpRY+BRQy/N+bSB1jaYdej1jw1+Zyp2UXi8pTxwyrOsC4fxJT
yHQI8RXiIC95d5+SqFudCvOrg6R1o2JErJ+F277Jjir6ucpt/sKdzoxuR0n2YJrhPbTdTCcJILDP
3CI7peWgtQ2JSpG8aO6nK1CsRUhmiZfNap7FOh9oPHdP9P5piMC1LJlc921xMt5TmH8EaPmZQEJt
+LK9Py7MX5oiOTcnIyVhMFxjmAzGR3B1/P4kM2CaNTStKfC0tisREF+PzA7/JycBTjbnKUnmxcls
7wK8ITmaUnUp3pKwSxVbzfkQZbJtlZcqHTDMWd3HaNbCD6oN0ZgXK+724pEVB6BInvhvKr0Ccm80
ETKcukAkFacYZ5b7v20hUIYlJt44pMPhBoD2esjd0DxKHJGuTBM3MSHurBaW9EqnpqSRH4M9CdWk
u45K+D0/S4TSJjyIKY4znxbtIYGSt5cM0fsRMgWS4q36MbmsETJEdjhoRhHjzTyogANROAriq5yy
beAavvULVdOQEH2saq8DdjJX5A+bg0Z4LjRVSKwATHzw5zO11yW2vpZKC/mFuE7sqVSR0R5AYXxD
BoGZkNBStOYOc+pv2HvaADIkyGzBNJNVX+/2Vv3jw+9kXwl9rMcMPkqWYXCaZoFB4+BZvR8p81p+
WRLFMMhUGXGugNQ/a1rUHu71qeFZ0huxhMWrp97fWpohSCNXOVBlUoANtF/ULThMR0vPY0CqQNTB
H4QM3POCpDSL42RGkVKuuy61Q82ijBPq2UgbHu2u+iX822RWdE1U1Pd6Pc97uESHzPvzRFr6vwkM
khFo/Bn/btP7jLnerjpw36MCssCPl75u/vCqCK66l78GBXSEbEYZcLkD+EZ0B0t9b+lnByW9aHMX
V2MIEp4pDuw7I0AwF05g+kb8A05G5nZnDLMMN/Pl7Qx9Texi9VsQLgyRLXrQZxSunZ4cQi8bP2fO
m5FZuEsSMA7GDWBgjCxDhMR/71pRPKMsBPXNWtba/I/k8nmD4pujcVJY2gQoW675mOWvC3sUCURq
9YJho+HRF+9LDC4wD3/5RZnJso7LoyGx8HpCtx5ilPhh39wljQXSV+vnJIe783YI4NM1NqhYdhPC
uC9tQrlMAWQ65aAasrt1Uv9hJBWAz+WO6Ar73u2kaANVGZ9w+V7QCwKmn066AB4IB3Lrs816K/yz
I4+pR8w2IKEEAUCSUn+DT1fPlJN3KV9EMUTvfO5Mz85eoFtI7hnFzoux0ctU2AbTIgZKHCead96P
snZoeB+M5B/4N29SZIfFswjSxpT9raTdJIDd3ZZ5IyjTX3IWmw6QVI+Sf15PplDAghBweNaYuslE
IdQvhD27XlYARcP2O3GOHjxaESXXgoA8t0biCXapiaHOUD4nM87WZU6l+0+HNVFBunOuAe1Xh9da
CQfQC2DYNmO+bHfYlxDQ/2kKQ2HF36x16xalX7sDeFTllz4Lp/zND2bjl48b4E82w2DhPMVvs/rZ
Ipm+Mosc+h8iY2WXUTZ2W/lOWPMxQn0axC6cGmjIoXT6qr4g9um/da6y70QzzeA20qwPuFmAKZKu
mJAB/EimJaknYCKeFqpcIjI0GiU8CiuDGjFRXmUDgIFf0aj3k7jdkM1NnX78dbERWLZwOBaQTlaa
+tmVvucKhMLtm9iRw+mLZdUg9+1j0iRgLaLH3CUHU9/BYXDq9H3kA/yM6cbOjGP030tTNLYbkdsl
SFTqzbnX6Fb0zDpNj5qN+tO5bw6kbmmMUoLkBJWiNcSO8X4O8KoipXQG+gLqqI8pnu62dg03upkF
iVQhFmZbqqH41Uq3mSo1M+C7higrIJAK1bNUnPD1LkY/HM+l1IqsXi5YUYXz4GMYAKUx3o+kFuij
X14Ml5Xw01hEnL6O+Djck4YC2qJbyXGF2fbZsqsxcmxQ0GfXdVv5Y9XCx56WyE/P1gPII5BNi0t1
vvCoCo7pOpqUv+mxnpQVI4A3t3++m55beYiT8S6A30do/xNCwIDoP75SGjuBbG/1HFdbEjkWDkc3
/zSuYBrhFb2JszObrtWe1pm/T6OQ8mKd5FIqN7zNanHqFmXQ5Fa8PxW5zGIb7g5x68u0Klny88qj
qn7NQpB/z250hMauWZ/BlllxgDgv6XvQRruQ1pQ58j5j0IuThXgoszS29tmg9n0QVH2aaHtu7j20
XQbhmH/bvOhiD/B7WTiyXX4DO23rvVlUAESYBsIoubXUGoK/nUYIPaKJgz3MhHsvv4PV95+V43eN
cPALsOK0hWMUvqTXUsT4c9LtKw6NPXs1g3JwRmlcyx8NH7h0ld5oRFbG3+IQzN3ZA33HKUlW24J/
LyfQvtdRJUbjlTPq0zQGFK5e+N/2tkUcp/2cKJ7HgYYR5ORPOd/jBLrrmTu5VRGRnjigrQ/EkqjX
gKGw6GhCTG6yX2iE7MAE/50mLFh7cBjxOUUF1RdNf5z1Wlzlex9zj6HhGPb8dq2ycujueu6ITZIn
gt10/AUoKUEmXM6lXwOdINeb+onA65ehkwTQFMsqK5/eZ4nt6LqooDUxr+SGTcULNwg5rUQ8CMOa
F36Z/ltONVUJ9yEMOnN41psBJ581qJrU0j2SDNT8p7E6+gE7t8u1+cTwS7JWdGcbCoQHJBQ2Y/wp
pQLmVRgD8NgCCt/1dYIYPUNKMLTiMalQ7xW1exBrDKJAazHNvxtI+TdcZI1q1ac2e+kGEnXDgpsm
j3cWklR9lfiP2T3CyOVHlDoN82shNuldjWsgFbUPTxWx3vhDsLYJEi8ZsfKCHfOsLaIGm1Rxmg2Y
eKsb3zL5wesdPmKebF71DdbujFT1PS6qc7MZtppKnLFbTwpleJflDaVsO0TIsDaKfAAwFeM3ODFB
H0+N80vWBlMf9PU8VjioKoh22sIsfTtYycm40h+7qNOlqimpF+qEsHG0UX2/5wIy2ZlAktW1nja3
oABchOAYhrO1Zqh096AUB5IwsgvdsTvZ/U5h7Tuo9wD8q37m0eRlTnKaI2MrAMaaE4VBmA7SojUm
K8JSgTdPKUXIK2Sb6vwo9GB45cS2J7VSNrVmO2SELjcfX/n8Ue38ru5J2davYvsBtUUI5Hj0ZiMa
dNOOdgrWyQq2vxKeYkiLx6Qp+wWSCYGSWKn4ePf8r/dbsEYlzAW/7tRwOsacowTMQpH1Zvo4dFpO
ae2BNGtwM4fyZW7Se0Lj5WHrkGaCYL9dFeH9uhHRPq60mRVLDkIXGPUmhWOo19t+YjHHqbqNT+IZ
4/pGG6zY0Y/z9pX7azkJYoR0GBXa08QRwnD88AD2YHpEbeKVKD1AvN9656kRMV0VPrBb9+tDKi5V
K7dsjmu7PY1rQeftVRuGZSxO05xDCozQH+LgfP/tx31b9yJbSekrLNWfWXdMbc49m/fEuNfEpXmc
JOw1ZAc59pWCI5Qb78UbUV082bXRXar4KMz0uAmJPuPMRfwrSD0I/OMj9ARitZQ6i1seESlz7NK6
491GHyf2ud10fUETI39RwFt2DvYw1I84GbOVCXNfvq/8ERnrC7cJtUAoMLkCCcAPbivPDaTgXHrX
uD2fO1p0SBVhIhNxTma5hwjWNaLT/lWz98a5Rp0opKO1wpoIBXqY1JPFqRuBUNQ3fFBV9oFlR6ZS
y4sgl5M3FIlwnFW3UIRVj1lzImCaS5D2WplDmXISJsY1aFXpXy69ElnuEcaGFdVufiWjHGNiwwXI
1mkuzdN0NXjRaCvEwz3OypANHdAefrB/k+r4kMxvsjG+rieH+T0t6jrXHW+/uyJVtV+ira9MlP1W
gx3w2GpvFwfjAYetVJzYyj/3TWSdjCuaYL5MoEw2tX3k02g1T6TZkLmdHzeI/4sHo1o10pZUzo1r
+FYvF18MK8ihAXykkAoznipmuqR3N9p60MTXqfhm0/uzxeFJN8yut1214kvonZCEdOmaNtjU9EMf
I5A2jjs1+Rw+MnBphv8Njxun/l9fXB0BoEoAiBO3Uds6gAMvY+uIOEEykoWBAr8CczlNm35F1KfO
+7LmXNJXrO6+i127j4opgScPrUyDtCjrnuLL3iLr6unitR6yko3Wl6g5dTr7NGwKTKO0ZlanV501
od/KyOrMPReodNisZm0iHy8GA6ukBL6MqpXuSHhWzWCASvp4miesZ9q+R0MP6RRc6D1X5C4WluEI
tjWzfdvt3FnMRSyNvQEbpJx7XGmOxCQWJkmalbnJZV1L+xwJcUvjt9HYm6W7YqmaQOBucDQpUHRf
s3ZKRhBit2+xLM1ptnpRW/ABffOd7ZG3qn7PeZrVFt/LG9vRI1BX6dI74CamG8BwyBPerKstOFqs
+26KrC9lmENujp19oDEw2rFOOo2gPB1Lapso9YjpUJ/L+S5rsRVfQ8TkcV7AuMfheI+r6msCXSgz
SegOGM1Ub8SMWnGUJKruC1oen4Xa64jJ83oAfqMhugk5FrG52WOhNPVMok8dHzqRMYwWVeF5rSEO
E3NCZ0tsnddIrsCHQSXrtkfvJP00crilPNQwJZVRO3O9IKFo4U9BTsnGdlblweS3NDuYUL82wZU4
MO2f1HJuExRyD2uMQbemn7YjznNWcu57xbowV8nWgKUo1HYbIY0RqzAKZlOOn+pxbT/nLpRZl0Lj
imO5/sci6rd40Nb96EsJXcDBu68WLRXO1r0TqDGNuc4to5GU9OI9bTccyAU9r81IYjsSSIoMx3A/
NiXOwsvSsCzQJWtHmcSp42cxrxswHIOri8MMVvUZA8RyRDWB/RcVs49O5lzx6/nNBALygwzhR8Ps
54NpxRZvxGPQbST5NFrjN/OlVF00e05r8rsDNupBwcsNz4iW7qtiDhR8LVZGYyKZDWlc7ITo/AyW
RJDyi6ltb7DwzJDL4w7X2FASKEuvasJ36rRs9Gyonn7mrVc56tcPE7UIAjv5iLf7UDfheQMYM/Vq
tD/3J3MhOSDGYRLvud07VqEzvQjX2yW7kjPNYecUOAX8GdCO8TU3NviK4TCtBXDrqwVdCWmSV0qj
5bsA59vWk7ettlL92G7rdrxvbThcec4P29oVBY1JyRHgAFh64b8SrwdSsLm6QGqG4bJp5OFldeQo
a4ggDUUdt2Ay74PYrXp3kH8V5BUxrRwCNpJSx2N0J8ahp8SP1T2CoNwII5IyGnwijrA3fT+ddp0H
H9YEMOu8ioDmWnwuLDXlE2b3bheJdBmknzaHTrZ2zRXZAsRXAyKlZSbhtiR13PL1dzVj8oEJWBvP
C4g0KJViOepg9tF3vscAGWpOT3s1ZOKMoiJPndr0hButXpp+LN5iYsEXM2Fi494QV5cZ2xVUcdeX
GSa4i6byUdecB0hrgg+el4P9DvaNtsrVG2jaRxAoE7lx8b20HNsSCGRERIDTgwKF/cZCsNTJ8dcj
u8eGAkuk++WCpZbwJWzVY9iHBhEqqb+gzL//FNL8NCEYPimwjY8bScKLfBqcYE7A7jSDPL6J7aya
LxmlXRR0Sh4G8TZFmMwnRbZWXaijARt295JrKhAD7KzKBZKB2vi7L8ThcGvDmGGp1QlApaiKnFtx
n0WZQPvht1XINQJ8ioqkK8j4U43sT7ON8BGunWQjOjw2FbEMVnwghFM/IlWGtmCowwruNdHgxFVO
Jxn8BigKKGEBSCS36MI+Gh8umbo/piwpLos9d5djcgwZGNHv9qQT5J387qEbktiRKh9bDxTlc+yO
6NRXRs9enzTP54kcCdIp+siAWR/3TyfZO6NJe10BPtSokBhKeEQd+xg1DiKUJMk3hxuBk7VTI8Ov
P4W8iSOImwqeFEsVeM10KpFb9xh26c0ahM8AjlkO8h0AnIoc34ktF6y6cCpCkX9jhOSBhzEJD0jD
2rkDUYax73mJfz75GEMB1rBP6pM9ftRdrREBPA2HdW4Q6w0OQyAazvw0p18OpO58jiyJow5DPBx6
Ax1dTJktKV32Zl4s7NSakULD7aBOehKMGwDLyKASM8u9JpJsptRN5J24A3ubaiPndWyWmnMcv956
pdvjdfh0QsJ5k4kmkMe/TylIcuIFcH9d6FAtV6rVClasZutTcGsoOzyFCKXgX0rUUm++Ae/qn6YT
yYx+e73F0QPkQLxbviH2I08pSrotsSf++xyZBE2aaHg1cFJ3TIQjjVJkQWbbXlFe2xpFFSnZN8Of
Yr85or/WbHR0Y6RYD1iG7tTvWyCVg1C1HuoxueSyrKNuwoo6wzbe4awdyRlYAym4JbXTdHuWWppt
fDpC+qsJgPDP3KZBwR1zSGA3BVPjouaCaRMzYwMgFVywc0qE44hCGw13gFLOO4goo2z6oLTT9LJ6
XFTuctAxPT0vmK/Ao1wgDGP6ync3PiaQyUrw43NPSD/NvjULrhJ4qAJ3cJt+Sk3EdhefT1Byk3xB
ds0CbhxhYHf87/xOMFPuIlOG56D/kuAKfXOF+QG5Ydbl6gQ8HXylKr7ia7gO1PtHQ7E7fgNS+1bu
mB3ycu1fS+OLhioNJqJS8mBrQTM6ZiDPpby7CSXKXizg0xwg+lAgIV+zHiLbhwpsFXDYg5tI/+SQ
0NWTS/v6+OLtL4AO0OZIplbbneGoRe1U3ROK1Qx/sr0f3JBTy++WLt9aJwEHeEwmLywqLKfuQ+IW
t7mwqKNJ0MVt2A1u+7oz8XPe1gIcHb9UyAUSBikOTPHgT9erbAe3V7JbBXLuCjvWBYFttSKZSnOs
ArKX3QacdSWWJCPAtp3JiBtU7gzOJ51KxnmkhQXO1oiu2L7TCGUET5CJM+CkT2Qn/vXFgb1vO5Pg
zIqbSItsdJvD71L3ZHLpbIBWcuK2BwG0lYYkM5Y/dqPnvxhBP+f9fVVmOeNzyRow8hDgH0UFmwB8
T3OiTcwuHbFUprT+INsKG0cTv8F7LQ/62lP09YbxXf954m8aJRhuccBq3JdFRrAnAH7cgeA6U0i9
LXFgUTtydv3Rimz9HlPXHYrPq9f4hin8epdiEIqfcTiZh3Ar+yN2SzPE89YqY2JgjAEKOWxXLP03
0xBryN03b6n8St6vdUgmuzw8iEiKL46AKPoheoCW6G0WRc+NMSUwaE3bq4ss707Sro+5HrSjtVws
O25JHH+V6Ad7jqPHalfHoasoaUF/Jx4NzNER6qdNaJ5KgSluWbcwq2iDuU47r7LDD6ChIzBYQ4kk
SKARzFq+HM6pm+ohh1yG03+tXqjAEqIFWYYwZ3Wz0avkAyvLkcOML5xF0uvx/iILoTkyyF1vm4NP
Cw6WmmZb2/qIE5SHZvUmrymiCV0MdbK3x8MUex+Vxr6skmpdqrSEyIFFRiuO3ZiHHPpt5Wmyo0Or
EK5/nIXLDXdyoJ2b6PnNgCFE8szof29q7zmo7oz/R3SVCzCeBMbgMijADDr4XFRKw2UKOLg0km9D
4PH2oeQOpFy/KsupOqgkrubGA9WF0FJ+o80T63FSHd+QnDpIqrcBBx1dPAJldIXXyNTrslD+m6s6
lHIfH8lLM4X9ZBK0yh3DPWOVgL5wMZCXJezUZWN6gufaPhF6Hs/Zgjmu8UQb0dUNSHm4i+3KG7Rk
Ssca9qQhDmD02m+VXbSzrTr3xtMY+QA1eqZBOgMctWYCKd22CyMkQTmbf624Em3JtK+L7bwzJSAM
WpPZyKjc36JKBP8f6XyoFrLnQizT/+L3PqqZddv/ZHq05T7FmU7KK6PZX7luMfMYrZ4PlTt8XSDy
/ofgIfjG+zZG7Bib4qLOF0tgRZ5EHxQ9YJdm5uRkfhCrzLaJ640XGC5s3sn8VWFF7c/UlM7NThBa
6dWbah2FwTk2DOrQg5eEjhPYfZ5NE2bKS3asl9ae7IVUliV0ljDubSOVu7wYYwxgP+2AcLIM2THQ
GcuYeN3tOgtgFRp26oqaPl4ZqBr3rleHqu/sQFqK6kIqpg+Cm7PEPyKXhjvbvcLw3r9o4goj53uI
Lj+D/DJI8bBFhND3JL4QRKWqBnduujQQozDHNrzm2TgIq6t3YY5k9Gv5dPer8MUkurD4p6+xAIXX
KzJdyxWeZ9lmn1ngNuWE8AaihF7xbq0hv/zI8JlFnyo9isZo9IJUNdrV0y9VrzNPIu09smYNeKHO
bVQK63dCeWSRYAmbARf1BAmufeMuhWYkj/ZiDWzgZ/Q5R3uAW+d7p4z7Hx+T0zJ1cxdump9ivK2r
EK0j1KqIXfyonEZhNMq5qcwiTisWrAWZFhEdPz5CSyHtlViFNV5TaEkkCGIg+7uoE9r43Cqo0x9q
TCeb2FtyDFbdxc2vvW2qZ3lspHE70D3Z14KUDTIrNTViHd3moOfKmN1ljuvkZXol4083XOICOqt1
9r2qk3soA/UewQm1jKwrdj4EsOMhdJz/RVnY0RPY5chp1LXgoqwcba7M1j1prfqzgQRvE9Y7Pld3
w3LOGRMA8u7NRIFIVTyxt4xxh+DmVF5B/8pTbZF9gITOMgTMBMqLw+6WCOD6KxXniP6/xPgp+mjw
eSz2A5SjlJIS7nLOanYnesy+QkI4zlbgFMG+8aT1PZ5C/7DXruGhEBOQYePsdvPAQYwDlymy7sz9
B1lEjBDFYNzW0jcXFsY2Bdd3vK3PCVbCAFwSnFamSaS64EZhfeVaIuB6NuF3nQ7lqQo2gevyvgaQ
hnyP84ywiUVXIYaa/aCZPHXfU1Qzi7m8GLrNJwgnzdBriCRfj8uJpKJGPXvD47p3A43JVDZ3WxvK
9vVb5bbBYp9zBAUUDR94D9A8IQ+OEiXH6GnK351NbO6DyaHYU05liaJ8yg89ZLSvIWF14UZs9Wob
yKE7WLRfLgAhCDh8VuIyxN9Kq9mF4DKOEgqmiFJPbKQ+7FjBe74C8w0MkqFgTb44MB/25KSudd6/
91duSwBCAK3mBiFUvAl9wSqFncoaBxxu5/LtJWZE0YhemI7xM/9HMlcRNNTGItSLRSzEUZ9kqyIH
pFG8wbMErqgRIdc0qjS1vjL865fxmKdH6Fx3k3eYo9VDOVDRPE+qYUwQku17TChPSpvkEITqn1k5
MpfxWj58eBPKR9KImhrCjWmVsckVO67qNR6G55oXUqw+0nowvNViHBGnC67dVLtm9D8Z/qWhHyFp
AhUpvGsA889yQV2JtC3ELzYRaCaDWWIf2zcm/N3qTysRx9B4rmVlauQRbNrQ7r5CRvLNap0yLFWN
BiuCYl5UVZRyKsyLrHxfh+svPlPVuYiM+yn7u3bA4VE/J1NS1faqZWCpjznwwbbbXMvDE2FvQ3fa
LVn6WspVIjIv0y0jzmLIF5iJlQvyu6SfGBSluP41gkWsPpB+FZiuF5SH25c+BmAXW6t6TfRPE0x2
ziUJBj4XpQalmYgV/GLpNkjF/yQZQGjmqKTpxEymJqyuc3IenLY/ZbfPDNaHQ7XMmITXxVaDJiC+
ckSGTbrFinBZdj1JyEYDxJ6UEaWDVh3FIXL/3HMsnCw6KJcQ888pfiBCFnha5ReanVKKam09uYv3
y5TqdOVKB3SxYjbBZ4D5Xxb58rBl1+q0VB2HsZNvkfpcaX28kgJp+Jp9W5/ahRQGTu2Fr2dzIB1s
wJzV7qq1kmOxg5RwlzXDUYDjrw0KFMGwZQzyLiacyr1JRpq0LKpR9mFBqreBtcu5/ydhLfnS2auW
NyNoz/vWsHN/9QBwK/Tj1YqrNUTXpUYAHY+agTg2sYXnRW8T7D75wKPnfYEwqY98ZeBrffcleTzX
JiqChBDEfUCuMeUQvkOzcw4NQCRn1melLhQl+uFxVvNbmY+/7tgTW1dJ88OPEG1UAEo9MKn7xt6l
R4zbBtvUkOLhP65140ofJDr1hxmDOi848pmh9dAePydLRTQcwOxQ6307lOtx/algJhuf1uZt+WI1
u/m4UD8cyMhJrh9nqHFDQ7ZjGBeXtXAJhQtfVAZoGPHMpEr7UpfayEiF8q8/tXBEYsMHgnU9f7FW
/j8WR+pk+B0c0pgQq0MlT8sziJDmaSmUFkMOyVX5Jo3MaQnnClmNkvfpYvRLkdV+R6cKStSPr3tB
c7AILkoeVTsC7qXcpBb7ajpz4KFqR4m02PLIhlWRzywwNWnAeUVhm6nPSTywp14+4G5FtNFBOZ23
RUapzkp87gqvxJEuffwnYSxTlaJgsOuKSu2aZDOlS3UI6ntt7yuuTtohAgjVq+nrVOQaA9Jq6196
suWUfbBUi1UMlajD+KM+1P7fOzc9UZKRBakdnriu9g6eO0ohfRvPwdP2KX33w0JVyxmgEzp66B9h
YZ1DetlEZxynjI5ehgayVsQ/IKBWm1TSetMiPo+m6KVDbAN4U8BG9sHVhjHeUj0MHJUxBtIlFqNz
vVK+Qq9abAWnajrgrTdxP5zs9tF4sV6zQIekcdmChw+aGSVBpH0d8PS1pgRXM0LulSTgvqOcfTZC
KIfvWq7OsE8BoYRpNlqwXDh9AVHLXAiFAzB4JOanpkKXxH22VmR//CdixuuOMBDP0mIN9C2qjHT/
AzdIJmFqB29OMYYLsghy4LCYdNmOtBNruA/Lb91xZfnhrXUYpossO2CU1+/fT9d5XGQ0T28avuhd
YaI6Z/EtC86xobDey1S2fw+2RKDM08A7jPo3tAzqhif7qZg9f0Viw/snT65KsJvHS76T1hix1vTW
mFeojfMcv/1p6xOoiH/uN/hp6YgpCtH81z3UmyoPsa2FHHoxfy+VP4DEzxHyAMT5dhOeOorRe5r3
7QEeDXIc8UwqH5HHNI7VNgSRHhXQHQt3crfrlG8kAc/hDfgEtYCGVx4pRgqsDeObI0Qac9Nu5Mow
tpl5+LF3lPAlB9yliw5E+nV59HHP+KyIOu4Rr5aFlUr74qrtxHXrESrPzvQyGPH+q3uFt+nWFea0
6TgZlsVd3pKB//9O1EYlKbwCPUVfChe0sJlJpRTHuRc4UOXHqSjgU5qo5jU3lWYnb9dxhOSqSyqR
UTxHICcPq4qvYYQkBQzXd7SMjYj3dQM2tVbWqXIEcmIrb8jBkiDmTV7Qt4ZTOWJBkleQ2AUdnR5+
I3BIANpJE5kZ446lPW1mIMPWvrInh/PB2oD6QUPoqvYuAwDxJJPQT/4I9lHVCIwk/u8upS8awPvg
qbA50QlpykXTnxeORw3Lj+3BHng7/MzbfunQUVI8dm7zT4kX4fuCq8VGQH4v+nPTZ0pxXAIERy4u
W8+FliD1yPdBmxIr6U3USXYRAEbkJ7xl2MHbqGV0iX/DwLj2etFaOyzjon9DNWsI0KSchtCODSwa
SQ22svqVm43petvNOFITVK//E0ctI4WSv97pFfbXdZ03Jecozc81ggOLH/xX6kilQ7aIBqTuwRXa
bDLM91WK1ZRfg5o3Fc7AlxzQWDgFHwoQZpM+Jg+pPkeMAohoAA6vUHA+2by7zNeA0Yw9mD8xTZJD
ffHSRGdi229syqEfeFQi46W0FtCxb7GQL+C28Uw22bz+/XODTGD7DC17fa2F4gGN4W5FHrQdaiJq
1gg9myysAICT+wsVcIqCj6E5VMGCrrLwI6H8kT2AIcSZpKbMCqY8Y9cGKTnst3z15Wc/mvIXEqG8
+htlPfsjlwBQI95CDZCRARO//PEjMg5pJnIXz67l7AR25chjSOjnx2Ts8i9U4OtIGg7VH3WTi7tR
aL35jOfCcUMltNS2+vqFZStkJYfrxNUxvjIMAfGU8XnQ6+nUmvBOkrwO56vXqBnBtRr/6QXODYlJ
0CRBKHGSu1lDQbG/jV9Nf+SLfCO/ZDGkAcDYdNqg2tjOoW4agZ1EaloInPDZqzIl3Q6BnZU5UuWo
elNwHFW9IpPN173YuwwHYfMdRnbbgZHDF0rkABSkW5bn0vNQU9j4CGYrd29AOJaf9kCLPRU7I/jb
pMRv1UzlafCe0CTLnVIPCBWuPFSTRTfRKU+AII99Rg1PguNNXvDXDf2wpWmH4ba91c0OcRlFYtQY
27rOGiJgp929PT30uMyFVDuz8zlrZ2HpOthn2krPFwdMFkL+4aU5aDr6OCx6dOhOWODsnSIq7at1
H+HFvA0JYvXvxF995aObdcxbCXSF1n2ecm+6vxZ05PUK4LM9NoxywGKb0yx+Nh9WGw+Xsraza8zC
1WHcQqlVssv9wRxDI8OTUyC/31niuzs5T+AiRShP1RzCuHZwJv4jTc8i11jm7zmk5tdjRjQbfBkk
Q8ymEWBFnTRotd6aYfo7H3+iw153btJg5TBDCt1Yuwt7FHDHVmyAd09WpLD7fW9hDLJdMcLtI087
Hpz9AAs1uRwWnysHkzKXS671oo4mF5k1jYx75gHvHV+J5jSOvgqihO2T677VsKPHZxrntABfVPwr
Yy5IyvY7QtuKc0Rd7tTybrez4BnkbpsLaUT3tjnYhIpPEzstjEmBEH64bMZTregQpC2BeCRQmL9y
F5h+c7WMn84JSGdLy/SKXfV3lQn1R90O4gTkpk6MbuV8kBqRIGmDTtEdsYRi6Ixl4kREAfXhNlD7
MgrKHmx7yRJEsUZRva44TJp5bA2FfHGbC21DZzLllp8tZ2KHYy/ZjRc7ETOexOvYD3CVn6b9+7bh
t0VXY4v6fwM7b7pdZEA7IzTTsFoccFtQ7r7uvcul6JxLQGRhCxp0jhUrUJx7ouhGUoHQpgLisXZW
ogA/IjdzHFXB1FhcJ7qQ3Xs/zKvP+xjW6DS3seBov+vTS0weHngpalRx1vFoQx809bt+sssu+nT0
lB8UM0wkxFePuVzXTOWFf8+pgGJGHR5XXT1vcA9r3d1L87X5GVeSVnP8OgV4PcViXZsGoxbVXZWB
Mvj1j36DFQ66YA9yn6k5sn7NLKarvNuzQN8A50iAFfQFKxYUrD12UZxDBHyq9DgyeNT1YJaUkigJ
C7UhBWZiWv73LTGjbs0U2AOgx1iyhq9/GUmUawQdhI7qC4YlU8MpkWFl8ckcAFZ0rTNxaJ43P8GQ
OrN58/08q0u1s+I0CIs8MFlmpnPMIHLx5DpjALQXGj/pa5TpuLk4GmEZX9baKr/83ktRKpVb7XLD
23BxyzG+y+Bx2S5Zq0QwEkPqlChzIXhmbojfzQw27bg/EKM79nvF4t+x/Kf33DkHrE2AYksLcwg/
lITEKMSEoBtOIJYAII+rTYJiKv9Z4cI3J7Gb2fMvtCcpCqaWa2I3THCEoLy2O1GWEh2RGe4wGaBT
ZiBxygS3Wg9s+2wH19nBvuMAjEFmD7JaK17FV2qppXJ0r98Up/3fMvEocD2lNAbROvr7OxgTBQf/
h9c4gmgv4x4LWJ4py6PNl4r3MdV07nKvdQ/8KK3XhTsVA1Tq5IOvBtFY51aenYGqJCDo3cXyd4SN
DZsp3mk7YMijcJy5zdETevAwfMyH1s6DkqxLdtDbgv5czgqi/+zTDI+UmgVFVhm329CmbbCwaZll
okVkfYZSPYwuDD6UpFQji7tSA2Iafk+NVjCreVyhwpZkfUmZcDP2niY863eOAD1bkubm1Huo1FTj
2O/B8lGGpIobehejH65v7Y/Ge5Y3T8GwHwah8tp9u/6rqOVRSCcJ2lmmlCZuX3t6q9uZXMO37/+V
UyVrlAIGbG7THRr5utaP5mYC0UBpkKLz8RgCMvQ1MPaUcGXeXER2uMmodUC+Z1vk/0T9k5Jnnx0d
Tg9VQ/XrzDhZMl9vE92fO9MQsaLc/8UjMPtBdQ5l1qxDH6y1yqAfM+8+MIWH7dvaXbf6qc12su9k
FkUZoYFNTwCnu17N24glnITkkIgthiDQ5aH5yztzr5J1M6GTSUlmLVwAE8m2Ns3CflgiTZmnqihk
g0vTDH2EeYNKBRUyAZ+FLUbFcqNlDKwKRoGKyFLBq7iBDswYDrZTMT6aiUbCAiVRmkpP2tAQOHL4
HXAo6Aa4rLncPewm5DtmSqqF9iK7VhAd9P2Hi6VYdOlC6lz1HiEJvRkJ0FQwoQwyoeMWNnG77w39
Nx4cwzK0qqfFCFe2HR1TYUucx4hugBJvGdVeaaioxRNwURO8XmyaqvvAErM5ZaaNp5q7C2eWAbEc
+hYMD8txKqhG0Q5Qa9j0SVXJUKP3Qhj3v6izvFBSz2OGGR4T/Hztn00YEHrV5esYVruEurj9djok
FcU/Z46Xu0KpWIQxOzbD5Wn6iv8/O66hoVnc0zl7DOMD63aE/73hTLHNey8cBCwL1jpz9H/kZu0c
rgqU/89EG+Aeeahf7csOmDfrPA0MEiALP8L1lkSdKsejpDppm7ChDeRE697ke4p+RidroPbAE2xO
Ztvx3JNKXsJcNCnvZOaSIxCgrgxotTpPFMiFs/nY9rUL3WHzm5zpjklgtmPwDwdbMnOKDUdhPG3T
rS5FJ4g8lOhP7VEgqLx3rPfHoayNlTYk7xWmzinw1Z1o+PFK6p5Y3nZMgjJoembtVVAGz3G47TGh
MRZhOt49LjLAY1OenQ4WZSN1EZRs2Eb5/kxZR34tXKVBzmgdDIhL8jVwZ4v0mzXozNyVrM5posyo
j7gWsutV/MWa2+KnVz/G+AVGCzq6x8f/TmtQC2EHNRiw2bsr8fHSP5BX2Ef8AOG/uCd8wBvzp6RB
H2j9RzL8rQJ0ouZoIlHU7SbvTmM4gGUJqEIInvRygrl7muDjIxdzSgSUsyJkqAFxV8F3iFMNehTu
HETNLJtBq8m0k+2GFGuY+tkEhfLLIIX752MporNin/E76+d6uuevNlyHl32k0ckfT7xSwypTvkpQ
2QB+Fowm23UeaMLH8FbahkrKpkm1lcd+yR+8K7U+FhxXjDEw2qPAAAw3dvAx08zD0/k30XCMWwco
w8VnZMzrxGH4WneN8/1mU/+FQII1/FM6QlxVibpAdXy2L5Y7/gLHtRAATBF+4KyGP6ngT/Fo5XiI
sCkByBTVo15xQQskNKy3D4+NAYAPEk6GSHQ1hGdWmVGo/yuuCbGZzb8npnLqJMnRjv+xqTz25X7z
XLYe/ZyoY6LcYr+oujxpqDZ2J6J9jSCVPmwOjBaLiwPBo7GZUwVNlEazlnmyoYaeYjui79OWyqAU
nZJai2Q9LVxo50ZOsXJWs29Mr/Gi3J9gS9dH2u7PgMN8uGYzLMcTLEJ6FM6sPoNuhKHMNowxFYMy
8lZ14VKrC33EwGevqUbcXx9NM+Pvr7KgAhUKd9C17CEmCSig0tqJEI2Vb0z8BbF++kmPIeyrFOHq
0OFooeqESln+9qJAAl4zVsGLza0tjl5tmQFjqDQWVs6zyzCRXb9ASxv25EcD+EKvSC1/xDtYcu49
IiSJ3Eh+QEVJq2UUQvcmaN6jd7wIWKQ7mfNNiBN3+lnsKOJx6GEY4iBQIjLFF3qfoHeDF94J2wnM
WRFkxBckmLnOvo1Uoz1i76L5LQvc3rGER8ssr+qKyVtyfPA7N7NGpphiRvfminkPYspa2uwteM6Q
tZ52n3zq5ayQ7+i/jcNZtFLsUhS7tngch9M5giEGTuhXdgxdp1fiZhYDdzeis/Blys2tz9BQ2ARN
q21CNqd5C6EwlFYt/OTDqFTkPlFtphHla1MwaM3MrjOHXF8UIOq36xl7fmsEyu+ogQTLG2H1PTje
pMIv3wqLgvnbUbniG4oaP6Pn+nyyXgfOJevcYSiG/djpErqZiH63t2LynRmT/js1W4waQG9jgha6
tzUlMGb7ggM0bkSQB5XO8WU+lmB1Kr6HIDZOlLyrJGvhfLY7dkFA+wzMxfBpoWRf1pUN45ggOSu5
+/9iTnuNmDrUAEOHS++vuryWDyhpYRZUn7vRg1c/0v++rdePKe3GyWpchZrZl1aJE7Bgnb2MVKw4
iD4qAtvrb8cpQ2OrQfRaqZFz7vO02RUVbyqSDc4yjlXM1LfCU68nKmGPfWdCBi2MMCqrCCQf5U4w
CBzsXq1qDAZE1GdHlvkucbCccV31BY0bdGCEH8QfLrGBqIYzBs9mToUmrHP1LMiO+tYASvzv7Xb5
gzzPyjUC0BEzAm4yqotrqjKtYN/ydCh3AR0msD950zPtoOrkEEu7Lon5g+nXOM4BznGb95Up+Efv
JwsRMhrEFPEWp3shxFNbN2v6RjMBoTEBNTlAWOVD4Kq2y1hjUnEL1sB9SqnKfBlFKZY00dgs8E6K
RrjJxm9fbBufuPbKEUUgeANt1uJlIiGzReJpVPwiVmJdb3Y3w0Ojsz5Cw/CcMHTwGIwLB35NLaqD
Si/kPUhYQBIyhH43BpIAuquW+kNx32EPeVnANLicA4TDErvJ2U/GDGfHQegMK4377lqVVWC6NE4s
Ii40hnOWMVPIW9KsvFDez4x+eciWWc1fOw4TWNHrXfnmJRb8Oa/rMBayceVaRbqnjzvz4A1BhfdP
+SkARhYSEvT1zdNqWi4bg/P6AONISsoOxv18EygQ6QbjdWQpMrfCbfx/bGOAyK4Blv3/Vu7Kam5H
Zfi6q7UqZHDQ/w94spQbOdWtZFRbo/W84Niib4+czm7XUfi+vkbYUiSMaMmyjQoAhhbMP2oyw6DX
ltZBNI6nLzaGkUZphxKJ2Tak5PAXDIMAaAvauPhLhbwQSuZLkGAqVf2ijPX0vswoQQ45Rnm+NCLa
iOKP9UISTr5DV71i6V5sikSacqj+lgBfEUFfZUS0Sd4BdqquV0X+sY1AXKHDLPA9+A3XywrNwcxZ
80OWZl0+WZG2slK7R9ufsVSbrsDp4AZ1dsW5UyRpKK4JbgYrfkM+R1ZsfHa7amintjS4hYtDIt32
gU5A7kxan48fOQvzrGmOMF8mUqRxzw9QZFN0NVgu2yy90wYyo50oW29dSvRXnFCKbkFJAPYaJTHZ
zITi4cVyvLzZOjBz/Hs16r0B0inWnIehjvlAF+Ar84j3PtjebPwihNXa1nHbg+3Tk+2TEATKAb4a
X7a9VXdWSWW39WC3/uOiQkuEQz8GhhLPxwKUhtrPDC8e6yikA+OAsVoaU1rPaZlbQeGHHZ05kIwM
3DwKu0IhdXAEfaS8FFUQZ6h7JrrPtXRIIflcuI77/EfU59Q9A7cBvLV0BRCJfOXw69pXJin9koG8
fcwY/FjIQBDJ7DGyvvkgeIzUOJmh24821J8h82zB98npSNZeCnHNxhQ0UDMVI12XFGYS8R+Vc3zj
3XX6GNpefJ/PmiNiP0QDpRRi+ku5qBGEw7pepSDAQx1rr6TnFYzXpb56u2PaHtRmdo0SpfSanvyH
vVDKAK0lQ0sD7NAJRsayCCyzamk9tnlVhDaPdLe6QqoHpBFqyx3UKohPgA6LqIkYz1cynegO2RE8
meOgl3Ryfeg4F8tCp793MYR+K4D0DoK0yZxcb1k653gETC5Kn9GcjypvSfBLmLIhLsnZFToe779S
aTHuXKHCFrzruMLg1nseeLu7n4SWRtITG82BHsGSX/igWd9w5iYGvvG/mLuU0C1t9GRMP6j1l0tK
NyRbBxZDrIsWZrdnV1CF6z59px3WIQdkFJBxwndaMckfo8n0Oelcp84kYoU+Tu4O6Y0h5UKD5qGL
bRUg1S9LQCSHU9Dn2nf8b8yWqTcbf382H0YNyRA24P8RdIca5GFjnVqzZXbZVtQJSrqrJkKMmFPS
B0IIPq9e2hRwIBG+pTLvfJzMIDfvMoFnqzG9Y0chhH1fMRUNdGX5uRm44/DCk+pskMauOLw9iwCT
ODn0FRR0oenYS1qk7SaRt8U4p6X6CyUXSjQqOjW65U0GsWKLcB2IimwKsUqHL0qJsGj4tu8+w8MV
eH5ULLmjRndQ/JP1bZfexqHM4XFmN4ne5L0EGkdE1Xmbu9CF2ZSj6W8d3LmDYQPjWMEwLdF7qLmB
yXDzdYVXihRAJzaTJHHYg/oMUswfDIMik70LxOuzzCWpgrN8npcWQZOz/P1mPlLoGox/3Hjxwu2w
f1M5Q+DOkd4rea2uodjZnZokHQPu64QJqrWPTe893/5ybwNXqT2nqFeFa0hLBdc8c8GAB5lX9fYJ
mjGHgq+VNv1F+LmtLc48OfB4zVC6umDyWE79FEP/EPBbAmaVFIW5q3kfekFhtkGtn+qPzZ96m8zR
7396EJ/bNjbGfSGzHAQRg9cUdA8+Oe133cjmxDxnSwUpgp3Y2QrqAKfPADQlHRPtcqZTI4fbH/Ug
xIK7iA8x3hZNNESf6103bC+RzzT6ECfuhY6lMA6qmeenuKGO+vlyDZ/OYBEAkSPwtKUw1aiQ8q7a
9i1bWMXqKclt+oH1xK2bNa7jWc05wPjfKB6Z7bBQ/Nocv/ClK5j1KM7kuu+TPvPbkOkoEjOYk/cR
6IkopLCWmVqUEDATJhDiM2pIxTxB5Zsek9vl5EfZMjvndUvxkp60L2koYX8VHSJtZirMenBiZHCG
1OL27duLiExXMhwcv8D3IWfyQoD//R1rSeCew2L03iUD0GRVvQEeiQpC+9BUmHJSHu/egY27lh7l
vE2NukvoX18YsuqgD6MOobbKAoZcbLBe58NtrjRBGRWsVa6/mWmWE3S+kNez25i8itqPEd7zVsjD
vs+mik1tP05wIctJiaYXSaqyNLdEWSWuCMcl9hsKXNcYFPJNFXpAdOPhKilTDtAk/OZ+JbxDLlrq
C1ppzDs/2aApHlvWk1Q3R2FvU4dswfO9OGlpZ04rbDIjj5Px8QryGkeZIgkcSayRbgmKuJ50h9El
UOTxy/IoxSqyzprHO8Xmga4OHVwSa5IqcxoiNY5NiFfIEa3jauZOpu283I5I+tBw6FJQs4ugi4R+
ZorjAdva2OKv5OwlV305YFz31iqC6ciiPa3EcXSvTqQp4R+0hF4bBPBGD9x2CcTzrPKJ8s4RQKoG
a/PLgFsizOmYNwdNwlvy2FsdzOng6Xy/XNduVmNXueP9EXeqNa0KmDEnZlittF4kkkDrdwXyY+2M
iXRNaI9tUfQshbhzEBZgngKEN7C/RzBU7Jn09R+18kz5YMlVnyPtKxcJW2zeMBCrFHZ2I+xr0IHa
o1I2LW2MPiOwLDhS0vmDvTLpzoKF8aUXe1swUZ7mP03DI/Wq1YsIWI/lezDNvb9+tsbXhwuYAWIO
KmC7HvGiNlxR7ASOMt66rmw761IfVqlaUr+t7LNliBV5NyhVaNF8F0eDM542+NSc3zybI5T/8/Rj
jXOSyolW6BtfXCdN+xSclaR/91vT6vkuJYbjFYxt1fDcyze2ebbywKHEgaOraWLtmaG+KuZd0S+f
1huJKseZ3pHswZ3QSXQXHsNfpFseCatqQv/yqipiLLMyCJrccuq3td4beBXsTNFcbesLx9468erN
mQ5YvNoQZeYjleIAZ8o/Xz0lIFO9LdSCOVFD6o4X1cWT91I/UD9nlv5ZXkwd8bQAfcq0RpV+YzFt
aFMxc4tpJP//PgzZO5BpISojNizQQIQgjZ50z+Vy9KggUGtZ4HuivkAyz7NvKK8cv1sbIzJgRyCW
b12Imdkroqcjt5Fbdlwj/fLfjQGCEsLaHJsawPtp6GyFKQhxEjvVOGKTsRbXWw9T9uPCSRD6dEI/
flGqto1db2WyAYfko4ky45KSwpGAK8FMmoqtjyvAyIRlaEEQ44duA4wmdp6bhmoVZYLw7I0s8MoN
Xmfo7HJOlIIvKHBGCxtGYCPRAQc9Zh9oHsVGiu9c6s7N+ljlSWd0EEReeTgzLoWVUBExQR/uWNpu
XAA4JB5p299g68LZ/KqZQe7UoHQriQs66XyY2NZP/3i72XDHiWVTbM560f0Vv7NNTRSZKDGhiu9v
5T7ueXe98GKqB8GSjTxsPotTyFz/WtCzQJjhw6X+uaHV2LMYylfe6gpqRBgDu+3p+Qyo01gEVjfP
5yVJ73xd2c6x36mnugl4IJqTly0IhRXwCIfmHZ0WS81TYGioobJmeANUAVVpxMAZaMTxoMaITTYd
29YJvgp2qRqK9o2DdC7ZIrww8lU9Sg0JwGE0jlFhZsaMxyUav7ZKU8bGpEj/R1DEinlcm/nLZJNM
oekHm3wPqJc1uLUSWt2ZrM/Ch8m6kVuryeu1aLjChAyk2GUuYs+LVbJ6swapOIFCyZqozK4C5+B0
H4/4L2ES0U6eTEFGkf68ZUkMvZkKtzKvMVF5Q964FZfWYEdgwfesnU9bswovBNCjKQ7UeytvcEfe
qE9s5QMO/LrUGRCgpuAlDLweWASidtNlqI0VoSfM99xHypNbMFBSgIW9CG9UhAqHbA/Fu5SPWh8N
h3Qk9LXYgC/pqYpn8mt6NhdRfUv0gHBMYiZ5/fghYh1zh47LJLrbk3GqyIddNLkCfAksVQRQaB8q
MrAQEqxKRVl0K14+cekS1fvG8NOaB2/pM460hMLIkOR8iKeiYb6VLA/6B9oN8lmLq54sVuf60p0V
EuU6nkZCAYSZrSNuC3O5chNMArCxe9ExSlEX9SmY3eVU18n8rPXqweASWzwQjhKvqVQtSl+P9gE4
CySJwZiPosXpJjLS62jwwQJ5rmPHOCXKprDMhkTVTHCenGLJapenij1mwp+Pi9UzaVKpJ40Xpvs5
UjKvhB+llzAJleuPzf4TVVxYPWHQnZI+KdjxlGMW/1IX9plePLdL/WkvTSyH3G2d/G9N9SbGs2zF
RqUfCF70XEFrZq7lZ8jcGJs5eKmEHZEGGcn1g+/dMG+MTWPJaLrfemIabYdYY0G6ENMo3fn1VHK8
iBWFA5bKTncEh6ez0VmSRcgO6fgYt47Uvm713Nue2hHd3bFccjOCzyA2VotQ3hclfJT30N4NALtj
eSbo1j9PqjfOLTVupGBjx3562wTTtTb/BxBcBhLZwt4ChnhAvr4k7fAu9gMzC223aPW5mqZiVE4X
TX0RC4GEjbYF9xVrArYj/12XHjo8hgDt+vTBjvLYbxds/oJsOO7VnyKpRvr4COyoralqLcKKtcU5
+pXvftiHCWpgiP/ABq+Yp2HEDqrU+FzJpqjHGYGX5UMgUyPwAxjqpsC8VGdjcDyzjlXz+nuBAftx
exxlVmPVEWAtqEF5mO4pOg3wJbUwW4JiAkhb3IBOEpSREOKBQ81Vu+slVcn0Ig0lCEgN+O5c2ZDm
dv9pXBTSQESQE81LIOcgwP1GVKAUMKeeeVFLXJeK2WJc+5+iytTrHWLGXkRsc6O1iqPhhtJ/wAu8
lIBwONk+91P8zDjVboIxWKmciDWshMK2foG0/dP9RUgujPZcZRC4oXKWOBkQ3Z2dupnCu9aQOzY8
IqGDBtySK7YMa/41bq5BBzqxj6NcIriaw6mulCQHjPwL9IS1dLiIq0TCbCGzt/jMBT6HSTUqHzNy
0euGszMRvEnnHJajOpR/ZzzAi9AohO5UH2VFWlcnrUb/jpJ59AnhpK1U7YSG1o9HvuQ2NrEvZKMj
7Jw89MJPscVS5L0pOtr83LeylPLZB5qOtHEPiQO/4PocOy88p+3MrAUtqOp5w8NxYn5v/svov8HN
t2p7lbnxxUpZbSXggBK3B/tkmTb6MzqtNSEoHzgXqy79V98tvHK+usT9xpxMngu51hSUbKe+7CUs
FghArBT8Xp1aeU5wx5GDK2/rH7TUdPqwXOM3LtpP+zTkncGaF6rHUUUGogulmGlQQk3U0BhxMnme
WBXrRjpWpTBkpxkHmNf+DvAZwmY7ptr1Ft1G//LXujy4vpcezSSBiK+adoSD5rZ5ZabnMFnBlNWb
hda2EgmMh5xlrHyqn8EV1c3lPrCRPVXQLmPnoExD4Gzqqj9gEGlpeuRWbfwBGncrKt5IRZzxm++c
ZWkjim/gO+nnKQyrlbEdqk3S31d/HEhPz/VmFENRM8rhbpvIoDkLujb8mI4hAzYHNIqvPDWw8qis
mSx8MniyRUf2xwOQM4bIyh6u2/3MUqPhahOBjyhlJ1A7oaBqR5kovCRN/tUZZlKTSYUCs4G4MBMQ
xKGwThL3sCfT+cVdZWLhV3MRW7aYXH1FuRtWFrBFuUtVZTatEQGLpgFJEWRysEcHxq+2GnUa024c
RPSv0Szmz5Js9c/rtmLkRFD0lk8t70N62t48R5K1YMrXe0an2L+FxFKQsoSeDakSN7m7DasXFXU4
aqbZX42Wd/Cn/eKEYqkqojkfk7aY1ztxCZ8iyI9Jh4gXJUiIPZPUsH4zssBebvB6KsQUkJY4qoS2
8hyrsx4VjZBu01rFuKRZUOMrQpReGoRmZtdjk4h/2K4da2ndF+Q+42dBdHGBFciV5PC5EixAfW0e
riKytAWH64mXNOrE8ncvP5aqSrYJbsA6S2PpB8eD5s0EVkzTwz6qzmB8kIOBF3TCTuBbxsYl7o4W
ZO3Dxn1CV/7Gupmt73BDgbcedTK/GGIijqhhS7bJexExQ8GoOC7qt4jCieIGqM/lfB+v3hMqCZbS
iduJ7SkBsuJrQrpAImDVAxmskQE1eayKOVJcUC7LF3/R+BIwhAJsAtFMBc4pXTX1rRAMoid+CM4w
tLlqeyQ5ZkLfILeQO5ecdpNTPYXOThEhO+/4HBfbSayNPvZejL6RBOBx6BTWJ/QvP51lHTQJemlF
rVNU9Cy8DvQlfhOGIXApiSY6r3VEDpI/lLyzoalFw3oWLZDVTHp+lQOrkqMF7MULw0I06JoILHqs
7SKyOQxDHIOEtm1BalEN+6+n30dvLdNiyTcpajbiFznNb29IosXpCpbqZcGy93iv+pL7+dt1OKLR
CQZyjUcGFxstvFei6rqqtgolWn0EDBtxkoSdeAgXcOrZwmwIb7RXxCseG5RK9dJVCKMqElJVpEl5
khtJchN/GqpEECeOjGQGQoTf+OvdvbA/ayJIAUG3MWcVPyOK+KbmZtHlqP0CnwK6/SZ18hcb5OJ+
1u7WZz38wzkTlgr7ZSOLgkzlIr0YzHzgtSDKhvo4kyK9OKEj6eRvj5r3U4YCxPI3IL5wGgp4k/4+
RlbScOfn0cAZ3y67CFT732J+HWzzfRtuZjEWc52ZUmMjauray8N5JH9t18vaeUeFxQ3Z53HHsLyC
aaPC3yz/iURo5YLbYGFL8SwBGQYugfXxb+i4zzu55JXS9hmOoxIEElHRag/iGfWtsu0ENWp3Zco9
mzSE+IAeHVDzgIC7N9f/MK3tB9V1UdxEBRhmJg4fmEwoJg9rbXnA/UfOoehAuGBydxMVVTYbt3cR
NBIawxTgipl7yZ+CT2f9oHNLc6jQ1WEzbqlRLdraZO/P3I+7t5aJbglwumWzb+kPItWJOP2bNdwo
ryRAtRaPXLEjO67a6GHM3+GmAEvm2EQIFEl5H32ebI1vo+2t9HgK8F2RNFlJv1U5ZLbKblreibMj
6is5TdaHEIDnUApChUnSaANPZ8uZSYwCf0PW0eEcOZ1t/+iK9v03jTvGxdjRO7qd7LQVnqY5kEnL
H/phOMl1NKGiPl6EKL21AKiH1e3V3Ghvf60CngCIjMG6LQncFl29EVjkVkRjBXYfUOfFCcJN+LK8
GmIZMFeUyE6ydvLn9mtEbEHVYWSOZdEliQqXbnAVvYMk+w0oM+zZN9R5A1nWFVnJ2xm1xojLO8+L
prFzk+mcfhYz9lDS1/CS+60rECdpwHPTNV5RWi/OyMD0O25H68Si3ClQG727CJ9sWnwTher3DrRt
s4CXdvJS+eX95vuwZ8ka0pAnBl26ZKsmrXKz+xPk4PPAV0xs55s1bvfLorKC2CTSscyEqXFXColK
upx8zAIA7lOtnvZhcf/V1P6XQgM6eraZUFTUTzdooyfgEi71FVAQ+Juy1Y5Hx2Vutkv/2wvWZEOV
loK4lwlpLtRDPjEjp6lTOYU1F20fpVj7UFvFJWFOTp+v+hwEAQ==
`pragma protect end_protected
