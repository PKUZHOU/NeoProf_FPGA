// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kIAzyDA1tt4n2BOm44Ow37rfmOe+6tIde50iLbnu2/cfOZLxRRpZ+746iUrL
zdkTV1iJLsWj/JZl+kldEqaXn0Mc3LeodubdRUpHzycevkbhU8NNNGAEHRkJ
60/ZZiPwAEYLWgwsBJ3sqdaz2cbi+eACNqZQOKlO72Pbp5vWucH42nZX4gjw
HvdkOIHkOJLTVdjUHwN0fEzzwrqgbQXAfFaWba88A+4Sgbc5ccu29OCnz+nP
p4QuNPZK6rISnbWMcvSvvAMP32yL1yhPSutvDVW8LmD82hirtfSw2iKDCBHf
jDHGKs4GORXb8FSsx1MRiCj+65oCxF+0ugv5r8P3+w==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WoGu38M0iHJvNGsG0uVrOvz5k7FxzuScsDaJA23SAGY2ZRxUZsxdte0Y8OFI
5n06aB1P92XyKCQ1L3b/KUnNtIWZgCM4O4t+Cw5xmX60T4olq/MyLZUS8FBR
Tyhy1n3YI9z3ydKKYJy8B/fz3QH74a1tc6P2tuWn0bb2HPNfIVBWOoJoUqQG
pwdWUC7balOfnXOWqvaYLAELCZlNK5Vl9iY0vheLYdHAAteZafKHLwq/xi5l
G+lbdNKkfe5FnHj8BHdh5GqTLcOBYttgmnxLbAmin+J5RDbys+NyZ4bRZrww
IgYE4kDcSkYdGTHp9RWpvECoEOP8N82dauRf8FWIag==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
UkGY4ThmjwQlrR4IahDUHszkeoC2nDLqNIoq/9Ryn7pdCF599MT+Y5egLzo1
XHcaDGZiA2WwPJfjBYJ/naLobTY40Nahy80GeDVh9nc5hWScsozGxSD7VSZo
E8HNBwVjRZu/KROPItAM0TSu4jc/D/QD+E/TwkTtvRAM5nPNPIsbv3GhaJr+
4I4dNvYjze/JB2OHM3nsCX0JFJQaBQJfGGClRY3PRJUZ5kL/cDfq8Mu/5Ct0
AlupurYdo/ovGppZUGsrFsxEnaos9pq5OXkBYgWKCRU33Q8AYDqaxWQKrHjH
/FtNke25v4o0uicWsgNvQ7PbtqlnuSnMaTL0LW3N3A==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qsgin3P6nl6NUJZ6pQ7Cjxsv7/R27Hp95FgfZamdRcRjACpjZuGwyuVoml2i
OfZj6YGcszxFEkjDWJipDAL4ACrPgxKAX0dKPICX3HMW2Xd/NFuXaBtr6TOe
xlvDgZWqI3cI31UrcubvQU41E4IDtV2ae4Jx+iefGFfiAiGbhHQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
utRTefGHhsCFofT5IpHw+CzAy6zgojync9cQnyXspZ+MhclaisuxeetbFz9N
eeUAy9JXDFEMSlU+lm/w79EWnHJWkIWhY1B8aOdMWdaMGB76OHm8YV9HYXYA
68NMWmokPt4dx9cVmJIpjq0qSWIgU6mnm428YCYRNdZUS8AIwcAMqj2KyGZK
5xpn8NSW8VrWYJGuAasqNQc0bjvG408AQHRoZvY3SD48Bgw9FEsjYj2N0ZOf
W2XBZwCVIsOLWQnHZAbJUGINF0IT6j/TiDeTjYKudHvjohhcxCHUB4Lw3yth
CkX5LesTfoSD4rY1fiGRCnGsUaMrYVUNJdQ9mqKJBw5WwOxxpRmyYPZigvcw
i8s9wZlAJD5L0bU2XK1gSLV9LMX6HC6E3xw45ccskozbSI1vuB5WBoXDRcT4
oESbgsJrjZrq6L+YivO0IvnRt+tAND8+wqKoVKkCJeM9hGKKx8I9yG6Jq0fq
DIz8tZ0VTOR4PoLNpxgkMLa/y9ChmH9t


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
lJuTyxf+YwV9MN+X44OhMRa8x1cKN19wsQvn7WW0hwF+oEeXxcZzolWTkRlR
Z1cJT5/3zdMGQcfWsy5KpLpdfjkILFb1oCTeJ/2zn+2mWg1EtarUN3sJVeOa
usTC/L+mJQk0M/39lSunsdngbzWRVoHZrLAlZw7GE5fRkSUZUOU=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
QXDdPMS1Za3+mej8el1CPvv56CIbMn6u16meOaLrrwv01nj39wC3hPXYGxbX
4O4byivvYdEBogPLSl4Dt38czIQ//+FRQxP6TUcFmeYvmaezjuyhnUbDaDAJ
KEJenNuBSxjfHaIZt6BsizFlruVHoL5SJBESW+oXp7b5PvyXclQ=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 46944)
`pragma protect data_block
KfC9ucgQVdFFHSAejjEVEkmauuW8Ea1eC/uui3uQS0VuDeRsxL+o0NIMV1Em
MR5Ek6fjX+6iK7b/nYYJZbqf2Wuk+FDpKL8q1pwkF2k2wpaEw3u/PQNVjMDZ
vywjL0kBPCNzlT6CuyHAjS14xOvX0DQXeP5GsAoIaRsstIxUhtieUTNTjpBO
/rgtHknjkRHI0ZT3cOOd3JjiirGG5y0FCRTHYu9l8EyRfFcqA8zKQoS+Ne28
IIMznzVhY6LythU5olB0RbDZyth7t24rOGFlxrFOauaaFouFXab616JJIm/m
yk6uEZP2ngy/l0Fo1bHj7/iQQ+AKwB1dxOwkltCKu10AkF6WUFfkQkPk+K5X
dTUDrjpIegYSy9/Prrq9c7VjHa7h97ypmDsRYrN/o8abJCq9LzuhYg2bn+46
bsTin9sEsa+5sDBvNoCxWoJ75Z3AuRf6r12CZ8OA9TWT2kCtNNhmsSX/AEFe
zK1e1Bj3pJf2rrB7RLx0XV4uhcCMnJJ4m6jxaqWOXHAFyO++PvhX5xuOqs5g
HmAgOeOihql0fojTN0L0g0QZEoblJm70BYjQhqQWVRPfTFJyILVO+aXvyjF+
bdFO2oHqTyuAbF8DPb27rfrJmrHvMh+uWjoVKvpnjxTgt7J1IgSLo0NBKjsV
XAFwvNoEGN13Ybjq9bOR65rSnU49Jw5vK1+kOOihmQ4W6Yimlnkn9OEwxe82
DkZo+cYRmWN98gVlPJ+VuuD9J4qJ/klggVKSGDZp8Rgv51B7JNL//6UL/i0M
h2es0VrNl4hwCN+YudXgMS/aAXtfqlfbKBdsNYk5Ro2bwg7qUVa+eZODq3Om
vYirc2HigkNX8A+TY+TMc2l10PX6bwwSw40b9xSy7eWd41tf+rq5Pa8zx+XK
WFODxvx8SrobcCc6DJO1TXdL4KBN4bzf0ny/Y6Le+soOTmHxc0h7l90k9M9f
nU2ytD00imaZexeb2nx23vaZdeVr328RjfZmOyYb/TgHsxuxA754lwTBhrOx
TFC2vpbp6AVYh0+QyEXbWwH7ggqF5WiRYE6NRjR2BmO1gMvj4w17YfJiuGkc
IcAMOsvf5KbW5kzAKIVZ7B7SbGI9o3N2NV5neofTWAXVvMb45CDtz572PiDk
2/nnY5mwHsOu/zRM/MHcnUioI9M2Aja7sTwpTKKhSUvtttwQAtW/jDlmGOVC
ZtOfUNxrPBHXOKLYf17FisnkqWXaJ28RmqLLeyzeIpBaMjNwGrO7iDz//X6S
btUHq/qu6OsW0zTTEPSIqtSYqQBw0VX6E19yo3YsNGBqh/HqiS/AVELS3x16
2Im+waXXg+vBNqYWn7FQKapet2BZg8ZPz/o89xcuixKbJLIKhcxXOnFdB7Ma
1Xl1NYWu26Zs2vON9VkVQ2nlihCE3rpifmnQEivp5YPBYCQUfMELLvmS5m8i
pHRKXsPLazrZ8vTdiGzKZ3iTdXDBMTwm8MrEMZtYJHIzXjnY2AiU9J50ofrs
tPf5CtvkvDK4HwzdwWowL87JnJ90iUxVX94VUPij6hZ9yJsZnFRUdGKpAq1+
xmqtGq9TCam+vy14BbfLDR3VnokYhmtMIJZLgZXou0+q+S/HRdRLBhk/+z78
rV9Mz/o0YxH7s3Iv/dFLuaX3CZU8776GDo2uCyV37UQd2NfGjeltOmHCVgjN
/fSy+eiTeEq7WdCDt2NA7QWSK9oM2/SuUXU+pDdbCuDXEvxdysyXwV2VMJnE
MpIyPUBvs78nP9p4u/zmEX+ec7WbG2RKqB6ZxCIWrDRKrjevsToXbghZC5dA
KwmST9v2VwcHMz1VfjKNLlDlHGy7q1hHjKQE90Tqqvwf52IfqtEiXrX4Picp
QkE41T8fw1X/vM4D5TIFDO2okfgDM0w196acQ5ynRgcTJ8CxRmJxwgMgBTx/
9DcJNY1AJsu4MecK3NMl1so/Hsshfq1PyLNIR5Tew4lf7tjW2YpnS8MahzV3
Rhr9PWrEFrqxA8OnKvDN748YhdgIoT7qDasbps9+hk6aYuib0z/HdFfpRaG5
gp5jJ5y1UNbEy/E591qdcyLqOjEAi5o9oiEfTo471wwpmh7kksiKZ+zs4v5i
tsMmHnhudj3mvIByD1sfV3d/WRwYiA0DY3OxR/XNLWIDkxDEnrsbBiN5IbiV
kfkbI9BA3+0sstsFxWY4kOzyyLSldKjWWqHlLPYwazCM3ChyRe9zA/+Fg5Pn
rTLiLI+gLiAzZLg2H0HFWi46wNZtMdWmgKMk+n0rLy/TzSUncxUjWAJ9ustG
Cdm5nQnFhHmapMtA7Zf7rVc3vu1tKhLTF3DxwNnnCKJLbOZLY+p5I3K0TKJd
K9jFhEl6MQVXSC1NxeofG8Sr9CaM6rAgCSJfAaNrwTFAFsVf7yy4bHwiTGpg
59ZqvjHfpwwTMMT+Dl7R6reGqH/RDLh7K9xRE6mMTVHwuhGfyW0FXxWfKFpv
b3FEaF7TGuLLMA3sp02Ys9WV/WABUioflQSJMlVWIhmPxRVEjbXGoUSO1zvX
4qZq7gchBSJWwtzJU9tB3YN4IbyjVe1R+CoyOUzy25iKMHBsgreh/FI92Gwn
0cZakTuINMZjW1eqyD/WoINI0DP987mDkaUgVDlNZtJEZXmhRbf/oPKVYbCC
bEtQeH38CkQc3yQ8CXtCY8BqsKSaIF096h3ZNHiNftp5SYKS+hZQP8P3gX2y
3QEEm4osBEjwhYgFiSSD0WlVjNFF+xqS87tQelZqsH1JguGTNKb9A3/aOxn1
jrqWDHVN/6H9lS153gMMQfxqQiWmhwspKUTkhLq8xFVrQx/bzb62PwocOH4u
/oEZat8nD/IVmoEGg/J2wBD3qBs6HbyXr/tSwJbg58lEdo7pEOHBecSZdLl1
C35/H8TR4zf/3xAsbFlhuxrGnp4K4aACEPkR4Aw9xGbeossG3s0oUIpMjlNw
Qbsj68QnVykMYX6is540Pl9KsX8f6zPaMYgxtii59C1XD8k/GCQMODhd+H1H
SAQTTjJ0JPVDqqdG/fkHqKbq4ldap+HXcln37wWeEmzG9hjVAWsvCLPFsmww
/sJzVtC+vbCEXy95ReMfEDAfPRRrBQWbofwIAPqdZkECN3wEtxPTH8kjHgN/
R9kPzva92BRI4xl4v3zTPEnFIgF1QXAxo5hdBAFaanz9UBoXMPlcXkyK3Fjk
9Se91EGJT6zqXPtx1iJ/oOjk7yZRM2xz48+t2tHntsvHhBMINY1vlqBPJ13b
ym4yuCx2jVoXLAplLSr8ZXeE5ypuN8mpQCbCXp6gBhxYhFGGb1lIXRspnJ/p
Bsyy3AWfI4/Cg623NuKgM3Ljm2Hw0voXnshwOHNl8Rwx5O84G8OFjAWXvr/I
dzQ5ffM58fhthkwTO1qLnA4nbZd8ZReRaVTDTK7vD9V1G1r9yjQzPXZ+bqFF
+Ptkvo/tR4j+4Na3F+c3Z6091ivL2x68nTRQkZ5WX/DvJskYAVLj/4jspXLq
FieZHjiwk2qv+5keLIkgTNnAVpgEM5jX+Y09hRbTi04/65+PEnSRH4vQ02qI
mkYlrAsS0PgufK277mlGN9NXavwN30t5JPy+Jzzkm19F0Rrz4iRF46a0V8B5
abJD1+uU7cdOAHds2JYJKu1pIRUCYHrwknRoLNowVNOF3gKsOesounKS6gxD
+Iwu6nYIvMGXHfIjkbhcrJaGAbDu2lp5PLMLQG537xfMaByUvknPgpmdgOP/
3LxvG0d81MUGcLRHq+9dabMdEM0LBhIPKWwD5LalFk54LSJx1cFw5idY421C
U2SGDPnRmR5kTNbTHXNU+Y9c0enrjnDphHZ24S/fqnpCRBdcw0bgvQNKMisy
k5CrW9DyFZ8DFSBJdvOiwGzOwRvQ2flXivjvXT4rGOHI1f8CjSIhHBGMnBgg
nXtc/mnNWLYdnct5bXG2PkY0MdCnPCcUDtgrq9NRYQD6iPdYWELcbf3JfdPk
uE7s2YhIFpaCPu02RVCz3g8r/L6KrmARcH1Bi12L3QbxWNRLsX5EDzDEDVrR
d0Lc4N0tkZkbnRTvi+NHmHfClwCW8tHIbohTYAM8bAM7uihWCi66YtowefqJ
d1mrWpbvzE8rhurVq8awfF0kAxNmwseIZANP7noVq0eCVLmm6D7sym5pZuNC
rNgh6CCq3VK0uJhFw+l48l4ZZgRt2GK4s69l9FsDo0uh47OERvSKMMyrrC0V
32aEodJ4GitDSJhXx6/fYjLsIIaPDFgVWWkCHnaw+/Yoqo2LXeT466EtDqGl
90GBN8fFy2zUQDbmPlZcdkTOMHShEu+ilohpkiCvfZ50PwoyP2Yo7YCOHKiA
Pp1od30cgp2OE6Tp5yHLkLhMz4mKmp0rIvmG2XfAHpUJVBkAboge4UlByxue
8HrgGf0UNSE9wE01inaUvKnK2CH3PuwsW8SkJeewDORXisAyUFPHKlit0u1i
LEQNHmRcjOsX98QwLLQsgxTPs4UKCocvGAD0NbgIdLysGnyO7RsxkPmAHP6Q
z3EYwYc20HAtgCsKbnMrFWfADETxol5YSCQnm0CNsLPQ8aBUKEdTx46NPb3A
FJJwUXr6s3oHQC/cKAyaCR8QiGT3FZ39LBnQnrw55isdndPac67jKDf51mXB
7duAqCTvy+4ZRkwF2gPKRoHwmdMhajePliC8OXmN2Hr028/YMrmFfn7HcT02
MfIiiC0yY+Fylq70KIKWwyamzWADLymCwJKb9GFIcfs77fWlmGoLl+flLpAL
OwWwJPZRcqHHggI6WMEEGD805tUFLfjOusrpC38b5w0qv8ka38MkP1bru+NJ
gk9C5SOs9y90Gju6RQZ1dV9lN5PBb8YMH+AZahjP1gy9UZWOOLcI3mkax4yb
nvpiFyZBnPvWdwLWQo/ayNewT9djVRqshPas8lknJQCRXjIbl8CsYCwkKC0q
Pt38shYfG+cPogY3E5McaisJXNvXKp4KU7tTkM+/GPw9OknmMcVUsC6ji2aR
9JI8nhBGKiauCI1QQNvR2lTn7Se5OhzaKgPL9gnSMJ0sQ3ybIgkONF1WGWBS
neOmV0lrCeFfIm9eG+YfGrOUj6fm8o8sz29nXpufEEiXUs0J16dKlMAP3TaX
Ll873XYbRMBxIbdmlNvMnjJCw76O3FNS9iE/T7hYakz7KxPlblaqIpkH4cdk
ZOOjxFt8KnvCymN/4MjlO5yD7oKw9ds/KgtEU+hkhHVfGxrMi9p2anWZYQvJ
I5zJamJ36L0C03fI+w1lLDdF6hGJLIe1ciXV1IfiPORAqV2AqVhBpeCzXIE4
HJaR9YctK/VNFPhcxqd+iNefQA6GVkKOGir83mU7kKHa61l52eSScFuG9N9V
4CEN3+sC4hHsE/phZ2Bs+cASSmA8lgeUbUGVq4Yq/0eIXATyAfD1ngziIkw0
OrUw3xvlvq8M6RvGPkboW0J+G+eu9DkOIwVNR2b3SQ9DbRHH6KVwgiTKenrQ
t5c/BuipFOQVS3qLTfqw1TJ6VEFViHHk/EN4MHfmybyT/QJK3ex/pUsCctkl
rsQdouNmaM8I9q4qfypuLsudgOxRhRisVuKw/Jg+6mD5OykmMJYifUYqbsfx
hHTNtke5Ax1+lxc+U8RFqrf0hrWgZVjfofm/4Fv2Zw3iY9Gce8OTNFmR4pYt
AWX1xru2kcaHKetYiNyWaRonXpVsdRrFfbgBaroALhqfK1RQhksJz3pHfObY
jFNx9a0riAx2+aKpNwqVp/oshvhF+C/p0V9TKoH9ssoOUhVgxoUaB2jbrM3L
1I7foaxkw+OdPMIYY7qsFTSvOziecd31lMLe0EbgCXgsquuVQvuo+LYMN/rG
OYSTd/zFbj4dR+MDxyyma1cyHRd7SWgzGhVdP+9Bjy1TDvouwSYRY/dMZnrF
+ysQqTNk/aq577IpWIFmeqxnkzH4D/2WF3JeIgqGMLPFSfrYB4dj7029AQSI
5f5gmkZMKZSa5tFiH+tVc1VTCqPd6OLM01m7VZnyflV5z5kgCn1R9OBIiivF
kc8wyN9Oa4PncRFH5FPFoA1rbiO6Q75ftC5ze9sgJnFjcbghN4iGMT+cHbpY
cMeFbeDERjDzzNshoro+GxJ3bmPiUFe7uxq0bUtvRObpCl6TTvQByTedoX67
QLYMU81J6M6sxfO4f52lTjD+NKji9B8a16E62poLvVdp+/VcOsI1+qSp171G
W/bHJ4gUs+JX2nHojLBrB/z8b4LB2bujaED2OTNmIxuMyOPTa3Sva78AtNgl
wmjoniIndvsofA1lhRRtPG27gUN+lcgVc1ecSwfNGNXpkmZQmvI33RjWPoGA
E2WiaD3q9ItF09iqNZm2fIsN6/3IJxS6fbVQGgoAKNhYECyoB5nrRkZruQAe
zE7gNBwP5ZHHLO7mrLEwS3Jh89PwUcjRLHYEDv37haJLIUCnB+kps8CBOSg+
xlQ0561ytFs+GKJpMPpaH0H10/F119+0dW43HGxFWYzLU/2QIZjMAETD9jZA
fEMHpx8YfpQ4jEPVUTFhp5ytOkmqdxTOIZi8JbEZCHV701C6MI62dY9XwR4R
Nki1pXIO3p/IUz2dcG5MOxdhfqvEmiUPZDnt0/JvOjOMp49bvjmNxxWCfDeT
zA/0ATqULKKS+6AQ6LQQi1I/DdpSMx4y0Znqr6IbYv9KxcfpdOoXVuvU8xgt
0/HLCYHSciEMOaOql7tY1+MmxtVvIBVhQKdlvm/2DEQFKfOf0hiRnjv7v9z2
swZOsIMpAFjH+5EmHzAhpOyUBoyRPDpWNy7ylDAvRMDsgJZFhbg/PFxjckty
CHnew45r9DLOn8fd/+kwxYvW4LzhxAAKVMY235Jveuc0hKnonWSrD3qt+BSE
UfpTJLtnziiZ3TfVHZy6/WJPNj6QDkkUESfWkLSPeNDLS3AIlz3SeKk3Xe9J
dizTPmTuaf8o+8rljOjYws4ML1EllVIZeUVRL+nmhfcNDktz5IOssEybBtkD
rPQoArxWfPlxRSupmmaDxadwpsV3L8gRytUBewqTsHAqgUtrGziqrqdBmD6J
yuV5EF7A/JBgsDfrFt0ywJhAhHZuhU7f7U5jmFFVZWr6/11IxnEebmn1gQQX
qrud2oJmsKhWyF52SaOuN0o21w51LS2LKLuJzjtNGUjACDVVvBDdYktT7uFP
078uKhDNAXb+ickVrQPpUyvQIATFQ6XLfaQSjS3TyLG/opornT2HO+uPAOnF
54JgX1vwV8qVGFov7qK0NmxvkKpbuYpb/pI+KUDERAL9Zxbsq3FnNPYZiLaw
S1WaJdXawvl4z/b15HWyQY+dfbTC1KrvbaJ2AbcYRfvQqQzI6LnWINnVUhMl
8yFXpj5rEbyo6yDS1plXLYESzyvqsiUrjmD5oXUsxUU0gIIKuUmg+KiyPkfZ
GjJVqK0UIgHIzBlixCtobP692b/VgTQNCDE7OMJ1gw6zUxtEKdI8q3ANUrtu
AcHH8ALvPIijHllSuAulCHZF516p4UBQTW3wJpj8i8nW/VioZ1LmtS6xN3pD
lth5e6ud/WbeWSAnMUOBxY2lxNjVmj66ChZ7aiiemKmEcrKhwnwe5hDIwy9Q
yLUJXrJoJybb7VfApHwAQW0jQK2Y8d1fN0TEawUFiNyjmxTuHiV2UuFxqQVA
Y6xlUwwwsOqNH4Ux09nOxECrRwnPrA7cNZ8IWVScJSbR8EYEplpAQeSi1CF2
qPrbAQMtTJX5+AbKsMGSo9QHxmIZHdTZaWx2Rgs+gVA70KcbKIAuA9iEJy0+
sdOIiMaDWcTOgvJRdnyI9C37Gzyj/GjQZER1P9zHDpZuzjv86KNSqcXA9rrF
nmapFaaD9fCyn4f2EnehjF0hU7oM1WKZ0lW889bJbvlfOWo97/LkzYXHBmIV
O+tjb39miljpUV5cqxcpM91A1L7fGI8rg86/Tp6Hk7mMwvxSMbmOZc5yvK68
2AsxzIMKdXfQDcltxKREGCi84ZnTrRt/32c9n7Y2+mj8wtM7RVnBpG0bR9xc
vXfnIHC6GDWwDOnR1HB6x9DSDS3k/BVBnc0u99DuDAWXhz8QVWs0/9ItsHUT
IiqAutzUJhcSJktsDt7dtV6iQatzLC6UjTvuXSkCEOnQj6TLdBU/CzsseZJa
kMFNeQKY4b90XKWE2WYzxRFs/dRNjBC5/yBj2QP6Y4/BwzbPmcQfvsBOCNOk
UA8x9RFNR0PvGDwO2wY70DLjwKx02kR0DacitnU5mJVd6Hj/A7IgsKPkydqi
CFNtvShgXfNyXIoCS8U0ZsF5uPBf51y+GPtJnFxlLQy23wlDhvkgAKAy7dcc
v+g1XrhN95VKyXSXksGROASBM5ASq2+xqhUfHaKN+Ao2H8SWikc43SP46GCE
Oztca0gq6w6lxKbjbHMHfXF5JxNKtGjGDHRqBkW2qLxww6PujthyEGUTXY42
2ll+3mWe40Q9XRyTGrBEQEz1sbYQHTRDyQEkmR6y78IG8Eztxs8a+ZeAUVJD
XlD7C+fyY5ufDTt4/AYKoZ5DMWV5nmcu2SmDJiTzEti3YuKojDJp4W8YSLVo
zuiV2KAX7tXoEyJcNKKJ/enMjhGmpH0Naz1fEwj7MrZWKyCol0eDWihy4fNH
Bfu6AlTafq6aBpV7EfUxKhD3Sc22pgPHKcAOGtDCW1sC3JZkUQ04kpJfyCEC
gxtr41NPBY5GKxLnOGsuNHGw6Cej+MmH4jgEKn3x3nJOvE26TmV26MFlEPrJ
UqyWFgaZhXfsErvjD65j7oWYneUOat54KAlefd9MLl7MYktYnScTJ2DP34lx
Pxn7Ur5Vjr8etnPE856jCf3tCLomt3BPvqhvCrFJn1B/1U9A5c7tsOGXn1qS
uTUFB4wEW/BsDYKCIVTbyTWiU8Gup8D1C14YxBYO5rkXcm1ge60DXGSX3SE/
uTihQ+v025QrN7V1J2TfAG4YCy8ObnSi5QIjag7s0ghSxm5dbXNV7CNUG8ae
zFlRs/Tst/xD+EryOF6fPCDAqjf2AOycWPuy1SdKM6z7kuZ5afDNz124u+ci
m13n4yStJQ/AkuPtpjgZKrtuBdyhK1hhZayFkNKVzWslhO6J5/esmN8eQV4v
c8GdsfAp+2+6z5avEM0jApdiMTwbnvSpe/lXc6p2adIjmMuPkjsa2i5suvkO
eizsZMt5CpCTKhT88Wu7rKVySoE47HuegbgXb5Tjwc9juLKB8Ok6Fjm/7fZL
DO60PY0AgRp3elABTMMhb8bloNUT9kumyONljFimdsUvvJca2Rnn4spBEj7k
000a4Jz+KGN1bXrqkUkhtT2DIRAVLvuuwiazCfaGoSk8lbIzlU7EGIZQJdxD
gOd4faEfb3KVCoCCYGbI6cbfUiL4CL549beWAGD/LbOk1YHhyQuFBRmQwtOD
azB8zbmbguItFavjtXdWbDMhRmjyJ34n+Lof2qnqyvvpzLbii8blGEoJbZvn
Wux2HSX0Vn7T74usepmq2Zgqto72Q/RQULH0wElSs7BInjqfuE/kF1AJreiK
8AwykmgkK2n/zhum997aZBkoQFgIM/02osOPQ3YaaG7qHjfDGrjbptTR/C06
zL9ysrwiql3vR41OVzsomv0Ro0keIsPkCp35q22lSbC8DV4beDgZNow5dcxn
aqQiSI+4W87jY3RZwAoTRKoAsfJLfqtbb8ka9pptdJ+RyqoD72LBeWPneanr
dqVmpYQhiYPis0Yo4Oftc6mOSw28oK8RHDNUygeJJm1vgfxT8+KXTWAmZAPx
qSwKc+jqtrbrmqjLaMOofVE5X+8Z/uBGJ7q6w4y2ZypIlRv8kuTZWQ3kcipj
MVdKayTPXl2nD/aqoX290kS93xLyrNrsZl6i0cyh/6XBQnPsTACk+IMQpgJ7
D+xR0gNici9dLmjA8mE6e+905lEMLlFYoKHd6NdvCv3oIKxL3s807ATh4Dh7
fARC53bruT+B0ZSU3b9OMMqPW1v2rknWsMiJ7lnnsqBpDsYm1ab82qvoAzub
QsX6g8cwvPH6cXH0Ame6m7pjGkzlErKbSugDmYRi2nmgcOl3hTMDJHVqQuCk
9D8eVuRX/NXASa0gKG1PER0FM1KzTzA+UVUQ204QlXQa3kUi0NEpWLCfgo0c
z7gu+JzneSNqyqXQRAeM2o+I5c/x1Fq3SfjNxxCsQHvhxc5ZxqhNM4cNlutE
Gg0RT4ew7pvDxgbM56IDHDJ1lNkJn5ghb0U5wjSOI/oPq3aZB8Bf8U0zHfEL
ZYtAVggkJGT9jjyCzXdAgGiAznBbZzXilxPmHG+wL/etw6cBPp7Tfj/JFYhH
v3rnmNzH+uzNxxP/dXsfUXKpAZ7KaJfrC548i7siLue9YidIiX18YL1K+V1G
bozym0WDH7qEkrML/eCy3VHmsjlJH0BXfeIXwHbb0Vk3gDcgJZyMiT0OKd6B
tNpj9vj8aPnCptVxv9EWCdgfWFsmd8k8+TISeNWJBQRDVtNI0K1yDUXjQ5GS
28U6kgAyqPKsXdlHLGdMHpPOBaDmpit2/lPs2z5V065YL62p6hfIsEFWC0m9
N0dYlRcr+1F1da0QxEg7/F83IE0EtbcOeE1gKVX7HJK+5qw6Mc4Eov6aTQay
y7Hv/xIuxW80vAnMT+p45VXRl64J2EuUiS0sNLng7HBwIfQ0gshbY7vwlhFc
LxxyfptZX/lf2wqUxHEnFzlbWy7z9sb541n/XQ1iYba8lQLxzaDEDpbHpKQ1
LCiFTvjPRKPtNPXgN21ag/SK56Znqdxa8GQSf2H9rIy0LL7UR6rLVWdiNkTa
KPu/CmlAqaTVXE+hCRqi5Ol2C3z/vpA+phk+g25MtC6rmltpQKAmAKvwXnV8
MraGZkO8pNtpRD8y8DRT1EsmXT/TjBgnb2Rwxc02r9ORuxUKr8Vm1KGCFGCl
iJ03taXOS+EQW6x4bG5ScYgqvUCg1JbwgS+vaNe81xE57lxtNKQzYd2VyInA
wjX2Y0IRGH1UcQq1E1WeW2F9DhHooFooWhVOFeb7XoQbMJp1izFij3fpiPSR
wE3XpLL9WwXNFYBRXB5wxGzy3CXopP+GCD4jGqFfL53uk93Tg4ro7iA4EY+h
XPlbCn3ToYOhLTgnTrXc0TyaDr6OSP6uO1qSKxIsOzbsWZEfp+cah84htJGR
0m/pjC0PlrXQ7lH0r01pe+3ghhgy9zlf/RIkhT+ULg80lMWZrefnolNKtMUc
qwnMgM1nBDah/v96sBcaEqpeDTZpRzR9YXToQbwBAlt2661y4G8Pa0UiIqcR
fzLdNg+20/wTdEMZHu9UMwxfywRCI/8YutHjewTvYvn/Qemw60pTRJvmkcI0
MlOKb+y/qhQIq437OwWk/sgmEQqgiNnZxviSiBXNCmi96/SzN2/Omyedk7B/
DnOr6G7Bq9ZtzDyauSs9kTAGTr2P01RBU90vU9AxkfNT34VyIUfXC8lbJADy
FVVB7l2G9/zZgZYcB+Y5L2YmECXOB8rY0QcPDwdCU30EJ2SK9JiZZVyoMkgD
rHX87Kbmr8mf/e179+ohtbpTic+7xw4ZrvxBLID9MpYAtPX+2o6d0mBUDoMI
xoq+L9YZfTTKKsugp5Dx5ps9ksGo9Dwy8MGntEHxM9pQvgrd7ZTkibK8Mszu
eGOfYUk47261TETIwuQypBkv/eYxpPVSUdCB5kmp2W4WyhxQQYR4zzzKHs4u
ghRK0h7zGjzhvLtOV32ON1C/lUo7Tfp2+WeYiMjZqYz6lT/1fk1hJw+ux1k7
i4dhE98/p0I+kDTbTe/+RJIGswr5abGHR0yxJTjCpUN3KVrQjRokhFF0VqG0
MLdVR6jkknUHBXd8ZHVU3W80EFfWFbF9sWsTEDRXXZBxZoGjYP9Jb94HyIQM
24UTt4G9C8bVKzLeE6jW7YV/J+oDCAqtZ527KbaE2YHynp5K3V2XTLDQgO1r
hR9cPakDiCAXlxpbnTuAcWcHoBohAx7WBWviP00xWJPLg4F9ajBf+gtLvxCr
JIoJoj9CyzEt3xmZH1MPpRWNZWKwuB4thKBJjwqFgPC2+khO4NHHk/xciRsz
OiHnHDsUOd7pUPWFS87SJZKCtSGwtI41XjOk6vxXPZB7SEQUTt8SrCJd3MS5
yXzMUd69WaILfcapcqdiFrQBYSy8EGBkzQpJQTJiBf2Y2Own00dUsUckaOSN
HtvqqQKMuxAx87VLX+UoJ60ScFL5u4JBR+/5sFkQBYjNhRgT/qaig8k1bzOo
Wa7KGRmMd3AOFSvKjWTICsBr6ifAlsw1OGHvjgEo8ov+y48Jm+nZeDhSz3yt
ZBzBV998wqIItV4PU/cflB/rfeV76G6VGS5LmRLh8v0Q6SlD5Y2q9Sh4way8
nR/PhMtU5YY6usk90R2OPxgiEc1JZnxGuzrNixLtX9pLoBrNLzMblIHvfHzH
KvO+bddi14MowwKb9XVwVdgrw+tTTgPzBcMVGoGXpVOcfChwXm6Mi7E9VZJR
ESYo0VgSUqscGVfLVg2MMRx6nS1xQt+0W8s4xR9wNgRZNV/zl0bCLQZZkzLM
zwEpewwPaN5jqXMFHDfDCu07pHtwr3/BkNYS05cPHCPvi5bHkIQkXWbYcpi8
yx7TVMtN2il1upR8MLgyB0nw9YLXWl0pOMpvNzNrU6iqqHIaq8r/fyQVnghp
P5I8rpYB1HbkJNpZFfv2gjbpg6lS7Xm4T6T5AKUtpjSBMkuSX98UGiu/T5Bi
cF2TuLINE0kn7UQj1T3h6+y+BpwgipXM3uuMo/LLSHdwuU+TBSo7rGzY67hg
4D5etq32XScS+rUYskuxgecuAgP2crdVkLwjwS8vXcKCLKwCfOMUUx/ZP8nW
Z7iqEWd35qHlyO0wcHakw5MjybIpedSZB0KvdmRvoZagkIZbSOP1gxFSbwjk
FF3Eq8XSkyAzyvWIr7pdSI5yRh+859XOZpWE6F9u0n4B4n68U1OgVnIwShic
GtM+A5kXvNq7sROjv2CCEeQ6xrnylEHRqOfubVT9cxDsHJW627qOEI2Hny0S
9PLppYBvQm9cEOJ+HMJJd6DzyGlpJ8vS4DelmVwXKuqvq/e4KmJjgAQkDK9K
hywapE20ZlUCAMoBo+VHoz0z+hnQRUltg7qYMKdu9lZbbOTgT4QuvMrfF+n/
vqr7kDaMIDAgb40p+CQ0Pn3p2cev5EiBSQaYygIab68Q2OLHBjimbgTk9zT6
mNFYECRZ9mlKSVPhoWS+eCGGUMSDcJ24HXflXetj+0pEaK1K8iD1IOAh2gob
Zx33S0cVbHSGnUZO5weaLr3dEuqZalg/r2lxPK5Xd/E2n9l9CDkqU3RRh27P
9aGHTpMCTMLy6dMSbjxcTjdmNPfOFe9fl2a/5cbNWAJy8Rw6iR0WhaIYc7An
WyZ6DveTfuKV6JWvzrbAdZskld0ZB3QcMHWWvsGr4sZ3IL4E0a5N76P+5D3M
OnNiXHejWY6h+DoVS6MQm0mw4F04efaQ8JNUvWYg7hv0w7OMPRZckpqHJQz5
xl7f5/EoKn4P+sjS252jbV6MDCZw6UzJim3xaLilTi4EkwotuBHdfSjD5Dd6
xye/oNdo7/2XkIVynEF/qDqjUeXuyl6T8b+Nmuwq6MTCAeFAniSenk7YPFdE
KDZPO5URAgiFJy0kdymhPAOE42eGoYKLtEeuWdPuIIs6qzEeXTCJiWMFfN69
m7kFTWZY8gQDEItdf/NNhSs5G/N3EZhte9gZjbTZl4D0HRTFM6ulth+dJBFq
XYsDzzD2NPsQ8HML3iukYMtMkOlpyZkTAA+OmSzwXmaeumS+gLk/nl/PRrmr
sztSK+0sdyIBhUykWUYnlNr+m7IjFfMof9Z2UuQ36OGGNaRUTMqG9J8gXyKA
9OHMov5DTb9PY8iX373iqElmH/9jfY4rIZu9ad5MrUnMQULxYQgU2Is/h+Kd
Sv/UeWa+8jWoHuLDp8Ucy8kKO5HODExAaXSlrsWYA0zk0U1zoFTnF4vmEU+a
Ix9CJ3yVt4jdrh6cT5taQy4Syo1MNN4xem0lCnAtJq6NN7HZq3P0iUl/jC7o
e/OZe9nG3eP89AsZidI+gwFm+lUk/sYkmTwQ2Ue7/7n3M3oGZHSV54gK7cmc
nyV50rj5OGtBIiZKbJ735wd880J5WTmX3l71KmSKXSaScljkI4Wie/JyUEKd
fYrE3RgSJoexCAV1FLVQY1lfkal3dReApRret36XCVYJeUhz3Kyhc2Y8X4Nu
P8d880t2RtU+dvm+mLqY6fJuO/MEg7TwfmKbMqYSxyfit9QtbaxLo9ZRl7kp
q90JQ2j4Fd52q41FvvPASXYYYttTVboVvDd3Pr2+ZUN6gm5JwjVQoPJxJkVP
ynVNkKMkR/eeoaxgFJOUqSs+ktCg+FhY077PnLKg+XUIfMUP3ZHD51vxie9q
1uejMO1++6cpL/NUs/vC19cK6xuoIQ8ALfo9P98nm8f1Oo67Miuhod+brJ1K
2WKH9idSGiAL/WP/L9U2DS+YGG0Y5F7SwYZBMI/XqkC2JSzog3Qv8tQM6HnU
Qq7iOxCQs/tirWbzv1hHkOB/9sPD5PfBSAbVVYhzFcqBp5cnh/fpxGPABsP1
fMbPkjiSOXxBZ9Qaobz9NfYrQy4fSgj3A59dRaf05X28OMJHeBe8tMu7GE/t
9dJJIvaNOPkvOEFvM+91nHH1srMwsawqWNfjZX83mf6jRJ/pxvx7hehOaZp8
enFKUh6Sb7Xn8ciPqLU0T5tt1enDNJWqXk0Jvswsl9FYUGkxPupWZ2/6mx49
/ToxfHrmgAjo4Rt2ElHKko+oljx7U5MST/XOLYJUOoLoZ2GnjmNc0QI7QjTG
zso60zUw9tSsVFzpC5abSFuFWOUVXgJBY5b5ezK2MXV1lbnDIuRNHThMNvB1
WsEHg3THzAqT2BVeCgVBusz1IyAuTPygeP9otiwbQjiL0n/Vf44CLt0O1fGX
p8EArmEk3IZiy/OzeLfRbfnJUtgNXvzM8TL1pU1ClqWqJPBkqaKkku5fKv2r
9b+m12YcX99fRJI03a7E3LhX3MBUQ3w1r8odNgV5lgDhiTQ6qtB8sFzq+Itq
XY1NO6hJrOoAm63QqRBpNiCSeTt5Mr3sSM/+SVgyT8jPBBhQZ1w26TIcPnkj
fCPfSX1Nmu2Bg5YUKmc4WCe59PnoAogtYNDeIhSiRb3XlBz2eCpJ03p1i3dq
okhkwxuze+RlyEN/ao2Tij2mfMbeLkG03dnzqyNwPbHUKcSw4cp9dP5tDh+a
lfx8Zp10OUHFyAEoL7lopaIVprWUNhD7/d5xLDTVjF5AiPlR9ebJslisyY3H
D+lO5hZ36uZiJtZx/HqF5zE8WN4HZavjUpLjkMlJ53npHzb11X5q3QKK5dhP
rlZlUhW1sOx1myHBKdwb804CS/GMgZ5WPy8ANQxqaTIJairCgK4v6pJqFAxW
xzZwe9mcWDctyqOt+cBbvDIEPUMhpWzT1wKuaualOnf4kNVdV6123T367bFO
GAacxQwWn2/lE6WwxWlNtlfsETgwXzq5vKSyBhXznTsslzPUEtdPgy44XZNt
4mHFhWWKqBfnuyHwrraApXKbLcaMNUbV8faSm+Bvg758pch9K/P3PxA232ls
ZUWTVSAbIu1kG1M8mED9cIV79dk3tsH5NbsVkH352hDTqzAB8vmnxqvsEeZV
KpmnRF0Hul9uf2ZKOT+erN2QVf1b6nQFwyufHfJtpMoVn5RXnGMHr4KaRZ/t
KMqL1lPvziOSXO8NEDHZ8vfU/Hd3k5cUD70QFMHtBDKkhrL2NwZrumLASxdZ
A4MUYz/qMqklttXj6nTv3CAc18PW3+Sz18vzZqz1lzIzXeJJfVkNS67tgy9Z
JLT7luYKt+iGMe9Ebfkd0RIp5KNLDlpyUSrzcet9gc8IAWAEw5HdR4nS/40Q
NWNFUxjUsGbaUyoIUSn3JYz5UM4OVaUiP6/+cPJaBGmbFuzXRBdEHk4hBGfX
r4gd2LXdO580+g1zVKHVFLhrKg2ki4FBL0LpULoM4cXU7qjrgm02lQ/ShkHf
6SoqBhrAHNHPP/O9pummJYaVJCPaEL18JpURZhNj+9blK4vXYNENa4gK1Qn3
KmpMDYvKzpfMobfnDP6jc90jxng7YcIQ2arW29wHYnisxsAV3St4f11Eedr+
oHczBHSTOBAXd6lk7ehwHz7q8/dG+MsNk0O3nHI0xQB4myXuH7bJVnNrJoA3
qClKHI4DI2iz5mWK2OLBeRggkpDkUpLKRsLu3ncmKZ/KbgMvszN+vQwk7YWZ
MRI09Xcm5/uFjTLaFdaUuCCV/vBSSj8VtAVBEhZYHtXtrfeGYbgq345dzNyC
He8qBYk5CfP9Sv4iVnj441ItoSyu+EdGYVN+OmNY6lTHIhLMHfQM4XxHwQ0n
+ss3/eWnmbHAuI5YAXWxnTVi0RklJSfTtscxayIrkq3nnt5MJrOQKiK+FSfl
BOG/lgVvYIL4udufO8m0KNwxgN+Fh4exHNHt4VHjzlyRiz9yk2CwNvRfPipX
SDjh/w36fiL/e39QF+5oQOi7JXO9j7pHmahddkd2Hpb9ZnXoTfTEXf9rW3xt
CbDJNuVj0YvJmtnX9M7oJ6xbGvcOUP39T6PrLqlXsA08+gnZqiTBnIhXYsm6
UonhsJziGG9Q1Yxl98vqcms7bzkvEZTaLCLkwjevZIqoMFqe0eoA1Ork9uSX
cJFx3Y6vSkiGW0WujeQxX73H91q1H0RqhGGyq7tYO4JOJX/KXjO0AidU53lC
muO4+N4ZLboDY/3szPa3xDKbmF+24iT3RVadbTujtQwoAifhQKwLbmUTazNE
oOFvBWc/l6nXEjMKnFYZaFdGdqcvvrEJRd+t04rmiPhoWuFvzw9UGIZgaIIL
KSfyJhdS5ANsWCUUsog9Zkbf3e9Pb7p23OV/AdtljD7jO2KBS+QwGppP33xQ
oZ2LhFAFNYvudd5/pliP6nbGzXk4fF6FDchvEtl7dUHLB71k6ifunLjlNyRi
nso44W43tdVqHnBihGCLBNftEqbnghe94Lb+qqjLgGEbLj2LT0WwiUS1IhFn
UPN7IYL8MiI496hN+ECCCDiuVoZO0wZv2HEP/yP8SrJ7QSlhbwHXFlXeIKD8
aLXbyZTszJCmPz9tsuF0Rum3kaeKlGmhr8KOaFWDrsp1Mde/1PIBA27vOJTX
82YL/yz4e2Z/6QGsFGk8OSuCgVsM4aX0BW5TSweSGTNy9kYDAa11ZBVXAMZt
q+XZXk8An1Ye+TUPGDsfBsrTml8R/CjADBoWJkw0/ShdDGeivutaemytYNLe
8wVdW2jhtxIZBVhMc8s2AERXd0XOOaXO7yiRcN8irW1nFpGQLC5PE8N7icns
rNSztCg1vbrnCACOkFKeX6ODSTcKxiOrczeK4z4SBfRgOQgOFsx88QExyFbU
06bx2Lwjyed9g4sJ0JF9PkPnX7pOkXHpo9tokxR4lQDIpdBkBoOfGXBTy5oL
9rPhxRHT7Wrck8d5ZP6+P3tmp5mCgEMUwrHSg62h57mise5g6SrgflW1id+m
53yS7W8EjQvaGLcPnBfoGVLJP4yrM98abjwSiKkEgMOCm5LElZn69k0X2k+q
y2mw40oePT7g48o9rYHaKf/CDMsnSWFmPlC2+t1dMlcLraLIC6IM5xbN48Bc
RLay1I4JeeSIeHrT4rUdobS6+0Vox0OtZ7Yw+caJ6iWtMDmjrvo6hPUOOtqM
qThQUL3q6lBcomYYpgvg1ewl7H23Jg8pzzFRZ9xVE+n9CQ17qjzTJN4+fcww
8utRIb4AQOBvEJBIwMUi+d2yp9DOt8OEcbfx4Ie1oiAQyo9dCF5zpx50XQZo
KZqeCN2sRD+KG3yYnUvh2jN/U5BNYzZ4/EKDYfIbvgJMXt4bgPEcCdWwMJNe
/Be0C8admcLjNoyxOflx7IJJHfzgqpe1ZdDF/jAIN7GXxkU2aWUIwHvU9MRt
HfHHCibH3O/dmuCQulFj7D01ijf8GhO4NIWjaCRuJ4WizPcOfRmhkL/8B+Pt
xdMwkce6Kdobww6I3hNBdrSK1OZ1r8Cu3DkSy9aE1gCrLwO/yIhmu2rmJgBN
NeZki1f585PJRlSF8YOEZYyNcrpGnaECPefkdzxqUV8C/VhiMpMSzJKMoUf4
FpnGXIEhT1aVEun2+zFuijnS0Yi+HbjoFKwnvasl1I1b3ZmjWiFPekR/zoVg
xYmu1uSeWV8pIAV72rvhfj26uM1cXVS4U7SiXCbjXZnzMZDgdX65AIJXXijT
tyDJNe0igyAkB8d82hyBXDeJ8c8gunLQBf65/f3qFHAKLSfr/fgAdGzi20dp
4n5AzRsd6ElgK5qrC/SmTrXzw7uGZ6S8wbrjhFonWE8m8UymBIBUHSROKa6J
Hyy+xVvf+J4QxSjqIRBz45tpQAt4ChbYHjOtM1YwC7dh1OlOp2vBHE5zUWPd
UdC6n1YcopWqvZI6KXHcaVIYoKgdbBcRp8setATy6WwyC9XgcUfJESuTd0/S
QgsTH86kE9RejkoImQTjfoD3pU/nBJuZwzx7SDCmR9ETSFIQAZ8dGAiqGeS5
jkvYMpWxSRGtaBFi8u0d8lQL5nPJgWCxxVvgK9mtTPXopNBTvGY9fVCN/fDz
O9QeXKledC3dMfqBOU90eEI/HxgzJswyeF4tLJU3pdviGwCCFudkE7nIcPi/
qUqUqMqoBcAMcdl4+6tD/MuRjnyI9s1Fbaxhs2bnFqscFxmk1aYaiwgOqn4Q
no1sEYlsEQzgL2TgH+i4KK1PttLbfkgc48cHHcVRf9MU6UcoJ9QOEy4r6Uhh
JLmIMJuFJ2fjt0BkaGkT/l+BVnDPY9IM/IKLL1yamNMta7RVWiPbE5yKV6Z6
LjUc9mnfU+JcGbaXbtcC/LqHTliqfmaKk8zi0ZZ8VckQmHnHEuOmtrTjIv47
scp7jE7acEg++uFO2dxO/4UG8brN+KIbyK5/D01/rb3dKfMEubpkw/k++JZc
viM6J0sdBLvyEDR7q9n7YMTVsGHChEhG7Oqeu47iEqpC0Sr387oyoOo/5BuH
AEjxEKhruKXB9aMTJ41ZmMj4dcpmq7No7BhKsyxpT/qQQfnbYgnRLo9KUGyO
BeXmfYq4714RaRUfRKXmU8D6ta4cR2R/pYR+6IJxf6P8ttx9X09lPdswEN3X
YhdB4aMA7H6SwJdaUcCiCc6psf+jLrJTkqM1XGekxrGmh5Kvvm6HiNCZHanZ
7W9irKAK0UNAbshYLmY1mPKz7E2ynzKe7LKwdrNm/0ckaXEa/38nSVI11aQL
a4zDtR2PRwpe41yAV7A82hi9sfFA+FO2UOuzpu9EAGwI+3SgkhGiQQngZDU6
k2Ppu6aQ3/Mh9NJT7HS48kKi8Q558naD95QJUrPumgrY+uqkg9Yp2TttGJ7z
hLOYqohC+OqsplrYJBMPeL2u8q3EnkzMZJ/95hb5MSh8TeI68XG9S017Fj9c
Wnh+N5SsoTrtInEFwn0Hv2sh8ZkePYfYAU4Et9kR3lGafgnX6NtljfUp2uTP
2jVPGAn2e6KUT8d0L1L5r414FUXMHmlN/9YqqDF+nwl4ZWriKv+9F7foMHPa
rmnPK2gue05cGYBLucCJZJ7+AkGlkDg2yhBolzdfiBaZF1OatEK9RPRLdoUK
xQOffRiGX5s3SkAV4SViXLfSe0O8uLcHinvSln7q2asAHrNAWExeWjxe/Ei0
Fyg+zrdEfYOuOsx3ByhR1QSMC6wAHE5Xb0YX6scRltdaADdDHUClC7vTy2lt
bkg56HhNLVVUcK9N7SihQ/Cvv2YXP0dDD/X2LBqikKBVBruKP7ZxIQ6XI0Nv
RmyzvPStjYU6p2eciiDYUMEFgjNUqV331d9sdK7FyFsLGsB56XmwxidvQV5q
rqAlyKkZ3gyrXVKTfy8ykRghTyPAbpCIqRjASuqOLU+SgjRYwaW34Apg+pUg
HeYzdAO5D5Ddyrzk+yIdlVWPATA6NxOIOXi2rov+q2JfqziZqJ5i+Udj2saz
TrppDNwATo4QgGrC8Eh7Bwyb48kDPXXzRsvzRAbnoJpwKTLNjRsn1+gQqMdL
bVBz5J+9/dFSNnoPYy41pzy4Ke6Lp49gn/3lt5e2AOKfhAc5nMwZmnEzf5Jv
qghTRyJGoNMIp/45VC8TmM89Kjq+ikh5QKiwh/sk8lvKOkqhicISiLzbgpz6
lo0B6lTM+24KhVhkbF9AaO2Y38tNjwwnBOmpSCa3HI2DtVQWuArv6dqxx83+
P+OEDWeo5hsviYCiJWxJkukEF/UHAGzwwTf5XlFcw1kKnwhQvDuhQ5Hg2bFC
Xsx2bMbuaWYVaojag6xKu6+lCE5+BjsRnlUb8chP95sisvJw3zauCE7/3DfJ
tXv5NZTP24E5l7TbAmHjvJK8OT1c91FE5DvnEN/q1ECzNPEtOhaN4A9rwMip
anG55a4u5zym4VknLIffDvAyT5ZR8aROGAO9FzZow8dyZxcn9iYh+SC3zoKV
KF36ChwJvS0zeF1kG3dP0Yy3Sxf/eo+4uob1OFaj2NTka8ILKw3hmRTj8m04
NReafahOcp958QIKAlGP/CvHx5sLqIsPj8gBdtValRR68ht0RuE97qr8ahLw
wx2aOUKHjhh3lMsBrGRecVoLc0jk5bmbzYzlyzhtc8yza0hnSY2M3wE2EsjG
EAX+ue3ygSbF5Rdn6dU6G2ZuNZeof1sa52uMs7B3wkegm7do0c7RJkhRNmUs
rSYy2V+9ocNLpPc1t7vtz8QcgPxKGG1ZaDM/okEgbeFz7MagClRfDT7ur4gJ
ibxLi290WJh/jokQyglSd+bu3GiY8ALmqYUBVrMU/NsUEknFHyXbcQNy+5tj
4FOaysCYIuIlYo//TL48owAp4X4bj7lZX982LIg7TtmCwYjNA6T8Xp0GSnnC
HsVyMSXnNDuBwQZ+7DW2oVbgluk6GJoeiu9c8HllRAMg0ITjtGwrHOyy7f3y
gHpN9DTG4VQcM80c87kEGcLvVvVBevOxoxVLMz28jCeTBPLoo4Rywk0+fMMS
Yifg9sLIym1KW0L/1D5eOLirTYNklvlleXBJa93pElfFkrprm48MQW4HjKH7
AP6MRp/sqGmirxUsfLjIxykF8m8P2fkX6gsT5wcY7XwBUpjzTg+4O/W9Tgmi
nLObfXHlBeRn5214AVaKir5s8E6cr27gdghqgwHXIvbym0jiO4inINpiBc1w
S0WzICu6aaMsvQSPH/1+AL4K6DB8g1UdncM0WWXVa+YXenHRwMYQWoWb8Ei3
GAGA+7i4/INbCfCEHF+I4EIV7l99Yl1AyXlEOgvGA4xJCgXiI7+ScFIvaA9W
8vDUi0lyQEzau0hPUOgSXY0YmHwlUFBq4jKJSKWbAb64BuI5ansPafb9+bP+
DPYywXm0HRvI5OQSW1ObAc74qlpvzLTXm7pY1mJxkmg3Cum5XoQPpbpbruhx
nc/2vUlx1JZs1mLUUBc1aCAtgbyG0fww72HQ1DYypHc9miNwGsiM3y6bIQed
mKBxyoHei6xWDLEYr9rmOFgDa5Baul8+EwzPRdRka9RvIAkMuHsh5uV1JiTT
nVbFDPzlnv1MNEM4TkIpDHPZ4AJMVe1HQEELeCJY71jZfTiKIFlaYUCGDr6L
R7BPdeoB/GLV9lNf+VBKPHfE2V17CuNp1M7VJis4lCdRWIcQoxDln3P9K9/j
eoaivmCmImKgFSJUjUS/sXG/eLsUkCrEIvLpd7P0cuG/dqdbar1XSlqyfLrh
FFZI61pt1jIUs5q8oYj3BgfS35oIFH2veMVqTQLdnrandQcLDzoGtmv+2OEk
aDUmMjhlgMj4aDRsaFZLFDPQ1IXsgnrhqsAvTbff8YmNMLl52lVSeaIFREFY
zU+TqNMF+YEz+Dyo+QJWvdF6OTV9UELJWtfU/DhbNV1iAzbyOzJN4GpUMdyz
02+Xj3hNy+bhdF1ZY6QU/1rIK0QLQH3fJHxi9Jp7IDapKZTFZD688aObzvmP
V1ASNgKOBvuEE1So6dwNBxfprK6Jzz+xzWRPAAIMslzlBSGLdOQ94mrP1+pC
BvbBHDljyyDP+7mTR/s0FvPA12o5J/FkLstHXi8/xw2p3edM0p+PikpBKfTV
2NZwfibrpi5YXRc5DLAF2IaoyWiX8J5YZWlYpkVtxp/15RjPRnpB5iDuPAmX
68Qg+6n/7EvZV9yibjJY6+pJjLYFR9MJQa6Vn4hyxipQrjZ2Maw+y7UTbChp
0hT//z5Ibt5TK0pQ2U9F2BCU1Zpj4tV0WHGaW0N8KeDmd6PzWqW9088ezNvU
kopaYhqSD/ieRBvJMFATlmpFi/QGzU68CK/BQaYZloNmPPXsfri49Tq3ST3G
GLSLm7C4EcKI8ATRqLS5YCLTzRFaPinVRu4xOdO5+zLKDRBzoR13Q9pEgudH
pBV2q+y3com0CwEK7tnD9DcKthrpw4NkdL3tOA1czuh+vjGmo8wBVQ/0fiAJ
on4EZiyXGjzkrP2/2Eb3oBJiOKJLc/pWlg+wJw70XLXZcK+PzW+fSqGxr2Os
KNn8dZbJGyW1o/mSKkuwvr1w3dAlF6lSrZTn7YnpG9vpOF7oTwl2QyO99NxQ
dRnAPehOwGJ2e+FjRsevKdjTUmTTNltlXZ2qUL/9vqBqiGq69DYkibLaV8VH
LYALVmUfGexxiou0pr/SFn2MK8By3eVncu4YfjyXe1hwB5rUXE7y1IyrQkgI
+F9HthRMB31z7f1o7Kvf/t31q353At7ztVEbdIvVBKpy0Qaz99nekC9Y9j+j
NfpJ760cnFPccw/0Sj/hEtekiv1QLnJfZdl52zX0xZZJnRAL9UVwnHw3aOzZ
mcNXMZzoPKwwdpWlFn9PfWD01lzhW62yZUnDBZ1Pi/8BhwvkMp0/DILduz5m
JakgZELHui+Rts0irnJKCEZoNzZ7HQDRlRGbcQUAXnzzGueGl6oICXWquNV4
Qt95T8aGQUVzdGAzCw66nGMIXSBGWpvH+aT1/p/qKNI5JbZPvvVtNXuyHaao
PGKklIgD0VLpG9KIkyql9gTTy8HjGWOzBwOCyZK43Z2EIgev9nc4SbVG4mAx
VemtMzg/ns/4GfCnQb3GbWkn2FB0cers9jXs4lRf4w3l9mGjkWRhN7z5y/1b
w6bJVaJ0YcSQtU1OilpYWR2lPivTJ3SY/ZZD0AxCSNRCWxgSeC1Gql97KH2V
jFzpyPyTsEuzkMQf3adwGFhXmVmE+1LckzjF0WR+0PY9IS69eI5WfGhWFKjc
EaXEy4jpQ00o4EIEOO3irej9Ro9suPqT+VzWN+0MqocIhO/vGmyNwq4+2FhP
LdNyd7vsCC0aMODrBbNO6Nrv7uM7rA/BZQV6HIH++IFJkl0L+dM8Qyd+G10/
rkEvPt7KOEBuTlkf3gD37D9OhitnxBkUEFIAUcA2VXt02duq6Udeu5aoUVa+
tUmY3M4/Vu6HYdJDHPptbbpmDSWvdttW4vskA7IKtjG+X21jm1yKt0mbWVYY
aQ7eR+dNZ3L1PS40kH1UFpuQe864XEC7lK0+ArBfGvM/XOMF2oHRN1ITgQt1
CQxINZ5jAD9qxNQ1d4pQ4U3vPd+slHMy3L91YGXGH/yR/eFAsUX4h2IozNJ4
nTI2ddoNGTHUB2U01qBzP/8E3oK3z2oO2Y9K2X9OXgZaJrxVLW2RmcY1NM4F
5AKw0OeX2K51fUeXFBzhWLhfEpnkV1eBcyPPfKmaPRAWSe0kL4HsqeSLJFeX
8WONVwae469KEIAuQLG9tRd9oiZQ7GqMs0KuPUgDzA3UP8MyQ2wBXxrBkYJQ
hqpErZ8lT3EAi68jN0VdrljJ4EFtbKSuP6W/7nLrisgXPqa8oexa/d80wOSr
pX5OwvRfu8UPjyU47b6gwxdmTG4zM0lK9ByfnpGpFYfw4ShSiYWl08RaUNn2
Ja25gVth3bc6Z+vsRZbSwRmwUoEt0i9j/ByiDhWuZnDubtaeNIIyAkQWRvz9
I3T+AphdD2bQwe/52rGUz32P023Qx51Z2XYHn4O5TGbkXWr7RwP7e3k5N9WV
+AurVow6PGMeIQgAzk6bDyn8EOCPZe2rSjE7O/1swfLk0EvkKJV0T2LhxTUZ
VTr2ECDZH1KCYdYOB2/7M9r50bDHDjzqugoMdKn9yIP496ElS75shkXDxp8X
NjLa7gPpGUX+necURdJHKlYMXCfGK4W8Ht4eCrEp4DOOXmk+MjPGgLz+rlQC
VBxDyVUcPnDE9MEnUFJnvVhHc/nSoCRPOMI5w2UCYiZ17Xrws7gDo2S5iuQ8
RwG0HDhlQB37wxBVbRYTXXzK68TTTCWPoKFnaos+UsrTjhjQoCSZhasef3II
DMVG4kBRiTfkwg6tYqZhArrPDJzSJSuC7dZ675novx/Z0gRPYiG77mCFME1W
af0+4/506YG97kZ7V/hzVoTwV1sbd9eDoKVLpfqVv4Rv/DTZ4ztDk6C9hXAJ
pKYjF7/WAV86uwus2v4mz9O5t2fyNq6YUtR04dpZpJF2x0y3fOSR9PwWnPMF
Y4yd8iEsQ9xni9VAgRNmjngySfiazJOFb8PPibG704bwMN0/iqjWPf3oY7LC
QK2DZDMJ+aa3GWvifcs761krlxs5ZCDW4Nap2wzfbqkcrg/LHexPZh4AqD5N
31bvFEeOVARI2H1McAaiDd7b2HTvQdMC29MXcNT3JQOozRXlDO7qU3XtgWee
d2BTlSyNNYC3mp/9ITiR7DHZByF0jq9VSv7MxzSWW22aJQdf0nlphRFd4vuF
4jXMsR9l6piM+AfcocplyIOblY/pwkpohZRGpQ+aqKfNvwjrItaZ//uDkIO/
qDdgeK3lpVa8ISlmvOokjNby0T45wTkA0n+KqdJSeeldiKSyXqpIez9npZAr
CO4AAQvz5ENsqDNBbpOYRn7Y+55oMHSCFw+cP7QBv+uVEojT7x9Si/J47jPQ
7A8OEOD0Mp5ojI+DeYdgJ4XybT0TXFn8N+IKuj0XbeyUHvfL7ltoJJTTA5BQ
/BuLGUPkFYAb/otPBLUg+GjFE85rA6rZbpGntOLuZji59DyGwIrMMItaqUmm
eD64ClY0QZ1V+39XVtsywks5teoN63a47sDYV54/PVyT+tKQOxLP9II18U6Z
uJcbM15xW/G1KMIAT8LvRavz/rY3gX/PhFcRA9ZRkv762u9rPpa52eBeaSoH
KdaRF1sLA74ZWesQLSea4LHTL4syeVxEy+4JOgepf2PQ+X5DuMQhQciwCM7s
qOKGaJNAPHW0HIMlyMZYNFrKmuZJ7AUBBfBlAxE30Sv89f//Jtcqoj9eM1xO
r/JuvODtvYWboy1bhoEoShfkCMz2PFLE6DfH6wZHnAe/QVoLPdsgnGF49ZBi
rdjyN5dqA180Ohaub/lzXht5r5WU4npy5jLoRIOh7F8z4zLmM6k0hYTgUmo7
a6OqNoqSuICAoUJxqrM9aQgqLIg8ZEnhI8q9LbHmXJq7prGA2l7y2gDpCJyz
a0oELqRoh2+vLdcN6TASHtPNJlPhFIiMDE6ZwY2H3PhEgMDvf8yKErcHwz0Q
/TLuM7A3G1/zRivQnMPRTRd3aR+Kit5FtVd/TKbNjQVvWdD7DoztdWWk7xMt
FQ0XsA1Xthf+55vRHobCKOSGFVJEAqwSFqla2BGMqY+jRAE6fD2PeAhT9ni8
mfMvIId/d2TUHnhkpFfxKmBM/onjZG2NX0bZk3ruHpujsiWmd57fsMDJCXF5
BLIJQBBedVE78x5vhxniNArPaLczEIA0ql4MC0f5RBYJnZRbd+KOmX3F/Mbx
QsZdd88WHrCYurWFXCzVO/dJZtE6iisTSUW/bSkL49jIs178OGYvoteB509z
OSXaKhE66aDXXGrb3XEnkfCYFqbBR5wVVQoDzdMG4qBu7QpcS8fTHqNKxxSG
Ktn/ly0L+YXwQakpCmjVSrbmSKtKI+HtwsWyAXcXQl7knaWHgTrQMvHA+hwO
moDGP7eZ8t7qqcfwqdUNl98XyWHuFfVqm32sXKYxi28cjEOfQ/st0OgpEQGC
3+89cpCk1E0vyF59k+10QzsD1vE5ILtZTiP1K3P+8oiBFWkFgwvqMJAGiMQ6
No6VQhwvO5le47zDgDg/qQYl4BCAIR402e+aSqenKSWPWx1eJb8KpvgGVpDS
kpdNSQnGsptvHV9QjSoVCkSHFQCVGkK2nOyUiyuGaBR+NP9mpJ696P7mHYp3
04ND/AItXLC2ZqXpe/nXDDfyHIjWwc6QEzYGXJPss060N9w5fZo0M6rpTBB/
RzxSA9uMucC3mSWc5sque1EAIMQvhwTMSdV58V8WKxLk6UFV+yHHP2aSrMTr
Sg+KFVKZrDlVY4bPjyQg+aTBAMg/LJ550Ul+uG5PfoPtv8BxDRUvlH7D0xj6
rC2wd81upeNkV3LP6PBwWt7KDNph1uWrCsJYAYjG4bjtoHmEg+AuoUXBUbgz
UCb+ZmS/qm/VhmhXrgMY+d7u4giAZJuz1IYFWtQGdyOjpHi3m2z/SBbTDFKe
PDyf18Soruvb2RaBPKnzGa6H6m4704DcKd522oife3OIvvSVGzATGkzl3lLg
2zLelCwQSdGInjvf3oxoqr6mtZChhgbfjPlGxkLeavnMUP9eqwRBHAPG59se
cnlzxgRbQeEfUWxIMSHHNFubx9ICPvQB4ghbZhLvTwNrVmLmquUSvTg42kGe
ulOdGP4F6Jsu4zEObUTL8qDe1GZlUDaJMKV9QPrhvV0JoVpYpP7T9ezWEzs5
m5mPEl7NOQAOM4jP2h/q8LwZXFZg/saOjtHndyeJYsWZ8ZwWLTgZDfmqttNT
2UtdlhUzK6eJ5smatFd63rIWKbkok6AgNfM1Q+zgC291/aBCNQriQX2ivYqN
iAGqZ6xqr37M03USIGdG4yGZpwhuxAc9p9FxhoW1R22T5yRyQzEuh5vgd0FY
lVFXgvF+6oxc1K7nzD8LSkjdUh5HGg1ve+Kz5E19MFmiVCUIUKyuCeGotOGY
abV3dLXVm5nINTUZ5jfmKBLCFMUSX6U1itqe64zLjbdqB/oeZc5kMl1HdzU0
oIVV9WOmc56lSfOtGmIK4K7PgeIMO+iuNwIfvU3DU4bjy/OeYRkjmE32xniR
nK6CHrSM4XTmdpr5cpdmMGr0rK86ZsKKa6XACShkb3iuuiz/MAB1fTgu00J8
zRjWE+aSDqyWY9Z7fWz5hcKasefDJzg1tIi+rKv51pPWY589yxeA1o7z1Jde
mD0u+gZ3+21FE8AfAfhrducoVrnrIymc1I5RwoYflltsq38ppR36oqOvfU7z
p0id5AM+YeMfpB6ebGT/yGTm7kcfMLAHm8189PyiO/pCkHOO/fom7uRdCIY1
WJQcEHBkEZVb+yMGmkXl7UmbfD4AOtuqwHADglZJPlA4l2T2l2+/wgn/ILHu
qmCxIktWAETCx6oFQEsKOd8zq88hEqUlGAPyQ/93vu2U7ZqdxQ29dGEYl6ii
P8WD4OgiENmBonX18ViZ57WbzCXfVQBHbnUy3rStxpOlgcfFJ5q/mWKsqx4l
c0pxUbh++Ot4HEaWRJQyHYup1vqziZuanWZXgoYEV5rfrezQl4QnfUENWcrV
tf4Nhh22XDb21zm3/w4H6WupzFaajd+G0XboZpCCRz6/Wjl0db91ceBYux1e
JMvakpEk45NyQgCpIDxs+eFYjd6jXrsQZv3dO9cIcrdlr6hffU3w+Tk/0H0Z
fdykl1IdFYKv1G4rUNnALLJ+CU0emoVt01ie3I7dsQQ+q9Oc5FgRO+Myr169
AmWf85YlS39ujGvtBNF4bxnEGtaPNLDNMFOdtveZLvGbmCMJlJMl9JpxVLa5
+QeImDL2bk7PpRSoJv64gk2gGrw5Obrs95E+yK9I6dJswDU4sE3jy2JkEBF8
VBi+V0MHi90WJoVcJfbj0ORVNpxzxoTkr/I8RJV04TB63JoBdHQCZ0f9nQKK
j4MJ51DlzXAVqdkpyNx1WRjpHum0ZogO7/zy0NiUR2Aatp008bJu85w5fsla
Y4rpkXTD8IEj9MOggyJGx2qsXCSEknD6FaarzJUGLpLmBqpuKQcK4r6VvF1K
hCTnpGWuPbBFREX02XH0dHSsPlls2/NAwaDRnOukb3uEh/U7ixUxalc/wgNA
HVDgkgvM/TTbzW3rqNAOrS+nEE22dNxSMJ3PFZxxwh8n6bsfL3CzCeAXoQZN
TVERL9B1+kAMnS64MufEuvx+JsRhMiwOiZuuoh64XRVW+jW908uyn0czAeQ3
E17moh0BAu+kgjXpBCKnydrhQ/JjWc5BMmNqks8EAUbNv9S/DaIY8Xtax8Dt
XbBsEMIDPo0ve3IrLesOgd0/RKuIiPqQgrFY4T9TiLQiRP1x1/tyj6Ip5lI6
olE6b+t0rGbBsBu/75t9IWDmhUET+wYFy9zavy/iQ0oNACLoYKznDJFOrdSS
lOGPkmWOFrHjLLWJ4iYW0lRpvudTyAi+HeJkbnFzHvbevkAPHKowjgZ9ALTZ
fNo1eMQV/HAvZ3HXIM94pDhfDbxTK9GeWNb91XUJQaGHdmYFMVMgY94UxhoY
+kiTmoIDQE9VQot/LX0O2xHqxfRpKdaOWXnBNqMHNFj4ztZvnrfcxGWvWVvf
2bfD+BCsur1Qptac8Nwkilczhom2YStfUtEWGFdT90FBqWEnOrUQwKfjhxWM
eMpnhYxW0pTi1/1SEbEUaCuHSLvv2+/WCCB7651Hwbx8MkhwqvDHZl3g07fC
ISNKzWa6t/VjDKm1lPGkP1FZXScUyE1mfocfjWjl6z9AOxKXkieG+WbIlsu9
E3MIR/anoxtYCMclUZ8RFQWNXqchWTCLDX0WiT73QoP6wET+lxGdoWyHD5Yn
BWB+3T+Y9YHsE+32QzamQK0uTIm2Y/juIXo/xn8chNNjwBcolBG5IKkRW9fF
zzPYZ7rFqAHJMHGRP63uIjKYTGfXrw5/tYJ7s8tfuoWQHvDYGNHvRSkJZLdG
poerIzRT2iBHO518HuIJU/U6qrViDEYL9+mu7hxbeAvNbraJ+0iBogyIaCjM
8TEQ7YSDjqNoyZOVSCTtbgbFykuh7WKBgT4jYAyBbwYeownsaF1tEdSUiMcJ
/U0YMbij0+95bUjteKpwKStj9Hchd1Ca6alyJ7uLSfTeq1x9ITzK/eN/x1X2
9gof5gqpg30WPcRxDVQRdcyCMeULhJyLiGI8FszQ11B+NINEuWRcfnsLWojC
42yd0sg+8JdYrWWjion2T1nlYYDXSNeG3+KNP7wjQS1VsoCAK1EwZAKQSAxG
2mP0FKVNQZ+MRDB9yu8dt6yenLXbQoEYmdJmrUH4PrqSwhjKLwGCOUuSNQZ4
KIiGcBhnf4y3KiLylmYxjdZUPIzBcWhJX5a9JRfSX9VlFgz8F65jMY5ObOD+
G++9e18KBn8bd9xrwzMdwCePbaoGaE1mO7wmvkf1tkMiMKZtZoj/8zMKnXwV
/a0vsqcJxvO+GqgZd8lTgPFwGUC4hmIw2Iv5bRbCwiKkL1O9YlpgXMMxx9XG
r/xgL8ZBY/FJHqep5MchQt+/624X6i4u/goZ53gvlxwY4kxhiOkF9F+DlXbZ
qDHBt4Aj2ocpPnjmY4ILEdRJWQRM9zzvigkwB7kcaIH0nfWEGtlDdHlEqEg/
QgdoM/W4kUMYpLS61uX4hv34wnmlnUKMx2OW2GOIA3AsvFdI1NQr45fAHWNX
7vnWK2Qnc0eQOMczVgAZVeT+VUNbrMbPOU5y+roU4xy98m3SjP1lgRO+n2UO
uB9j6nf3PnBWNTOPEzQ/e00hPQsw3H6IHR0dJ3npDQFNBwF2IPo5sM0xUD+N
Q3KwLyVhhngKlvfJuxifUH4vnEXUyqrzL1BpJlo6a4wcgiGoUT1t0vB4SP/0
+6V1aS9ML5u7wDjGbo8QFjJY7oDmE5rJIi9L5DoOZkygFG77tiFlzXxDCQTR
WUBriEq37JT950VYf2LDtmhw+UeyK0KY+Sci9iKYu0wUTclWeE5u9vaXwcUN
q5TG1hmEgXQGMSUndZ6TWRvMvzALl/9Puaj/NQE2J8V6Rv3ZeuBc8UU8FgoH
HtIoh0jiuh5gfTykjTno5jk8SGYvf2dtxFvPcxjXaA+N1ODTB4VUd7hZmHMQ
lDTk+8Ziqcr/BqQ4pl7Fm7NDA5J0r2y/UfxgIiHqlIx6ndvbTLz21D3pRfo8
zoytIkrLYu2/mD3s47OyCEuGILxL1QJgqWOrbE2kjiGcB7NXU5oSODQUOkGv
VcDDAvceXJ9HfTF2ZwrWuQ0Zu6dPj67pj6Gl/ReLSrCAP51tvtCBydELI+FD
TqTvU5O+jqzYmH9PbqCPgN6MUlaJQn19RKKzKmybN6NL+st39IzqciltoGnV
mKxvwVRvCxSueN327OdNlkHXrpxqXmN4xhbtb7KhXniqeiOnT9Y2zsAvUrlN
U/MEaq7bN1M0/htGLaxo7itbEh1dk6JGxBPF1eUUEHzqQdcxGoaGaHkD9Qw2
buodY/WuEXMQ/FxFnNd34qBfKXRaXFiG42ryQnKohDGWAjWa8bBsiS7Y33MZ
dgvbDT5srLipdHvo2KDv5v66FCr5AJNh64h/nLZEFuTsbfSISdwKyr01SusV
XIJ3VvO15DKbrbu4juuzy72GdkA2oGal+d8pHqvX7U1X1Z2a7BfQEk/FqgAU
fab8s7agcVJ9fri6hXlyzsNaZnECKB9A0lgvOkn6n4zcY9fPhQ4Pzp0xR6pr
/IQPuXdhuj58eDw9U+i0utzUOwVmDuX4p4BDER0m1eki4MlbAaSMQ64RZMzJ
JMTY4wKHKfNheIsFELfhG+2bnxLGXIxgMZUgKEdkCm59yniRVP7Q2ROtGXG2
E8uSBNutn1yTcpq30cjl76NkVkLAbu41w7EzdiQq8sAsohZIYuNLOqvutJE/
tGu4MMVF/W9dCOXbIMq+y5PJq6C5uzJQoBDXd3eKEqltrnDpjsMVYG/DOMT4
N/wwqYPsPFBr2UblwXOUU6hODdLw8VDywwlf8uS7jtcmxAqQNNvGjG/T+EzV
SjlzyXbJqiHYohJieWVwb16i2bA/u8CWBgEWrk0SgZrKrWPwnXYZYaF/noKH
mZjOEemwZfER9r5fBkAbSTHvIrjz5RTLsZ2z6g+IW9/wJDTWlxyG+VHzwGPz
agtEXYhD3t+bbug+TzOGD4SRs69uheqe6vgNEWMrR+dnNtz7RKA9B78K0Pky
ecf+3GVqJfDFNziqr+/DBwmIA+vCDfEOVx+TnidTkeYvBwpcnTvURLiqR1dq
vZVUKKY2El7JPBUPvRVbEMuqUzG74mPTXlH6Wm8cfq/vLdB2uyD49Ops2VV3
bP2jTx7Cuh80j29k91ad8SDbNecCddyOLDq5Oh029AUOlcUppVFG4G4zeLI4
JfWVk4p9B2h8Zq9lJ1jBeUWPy5h5eUu7AO6fB7alb4GoscHCsXmp6cJldzPC
2vTTuROkofj72nOOXR2NyfSULwLsYqcXVH7ftMS3UqxGwzgbJ0gkLYcoMNqb
VJTuAtq/7SQvbxdbF8h1i9MtBpObJ4/3a1jBP8cAJgMtACxIxS1Vyg1lGuHa
eZAF64uD4mjWh2wVnlnqfcfo4kLCXJeK2v1i/J3SIoXbUYG8WzE+/EgoF9KT
i1zD3QqXGYsnyLNJa2xQSTW/yQKSiD/n7n4z9wI4d9k9o/MdM6AyZK4R4M9x
yoFn54sp/vQ1nS03xNGwCE8ilUR1cFN1y2f9d6GKK31ANCVWANL+nmXLZAzZ
TiBIX953PRO5xK25WULhvud+64NQHaNa0Ic9H3LjvHAK7x3UQgIYYWHkU4Ti
t+TseE7+TWybE6s6+O+TK7yqyeByo+ZVwXjG8XzvsZYii/4PeRPex3WTj+zz
gGly+do25Wmk4WF0Ye1nzcRH4t2pFZnZCY4IeOAizorrb24jFpIvikID7pUl
RXbGPL5zb1bBNXUrh0/nYtLjalZ8SHZAGkSRh3L7ZQAL26uubpz6cGLZgOSa
itrkR66mEJabvzs8vFGMeL9ceIoGetiXd3YUPUGG6zBusQSrsVKQ3ranYo6H
TlKnu2BT3IsPX8bMGQ+uOzTZmASknv97TNUEjawpY8Ad+SS0uzTcIRtyw69O
yQqOTNuHN3r0Pj3g5q9Y74rVZbAA/l3BzOAwWIbcytcFOIlSoyK3MKOPZ4Gt
O1cjHEmo0Fhej7sEMBpJfK+/iahe9Wluy2//tW/+bWC0tgGqiN/+jR45KMsI
Lgu0xxmfi3BEcL0eBBLYtUsGHpyI31clGi67w1PToXaHIgdpK0MHRbsRTACG
FV8HyysRQ3gkCgv0QpLrGbRvFfh+DPbsc9MIdvVaJhEnqffB28RTVih2CMTw
//RwyQLqjuVMsru91dqvglYYAFhRpaedwmtY8OShKdURVQuwfKN5Woy2oP0+
4Xa9hi9/X3BaHBzFAft0SYMS4Mjbtxc05cx59aduhlXg0GtM8s6qh6KP+iYz
PDtU2Prc9KT+OdW/fjWDBKatd4HDowVTnKIMkkkHGDbaxYt9HH8DJYb81YuD
LiW/n+vc/QYPLrXKBHnrBVRom+UESBS2N1O5V5DQwiS51T9kiig/7Qu/mzm0
j9bSrOfN3PGvKoIoOGP844mwcaPXrbGBr/c4j8v8iCUGB0OUMzDMsCFHMmP6
gIlbUzzMocL/IC96j9FOQ1geawZLJsguqecVe3ki4bPa/2fbJk98sss2cN1v
BW3y4LE3g9CK7hFvYs4kbcttK+VkM72E8oZKAfhmqCi623SnIVh5Flp7RgMr
OVZsnyHNkYU22dfYobglSXKJfBbByNBKGTvxYPeuC0qJJyJQ2YZmt/FoU5Ce
K82dWh82CNrv4poqMfeVDaiQehjL9TQvGeMBc2akOBks9k1HsEFLXOgShTOc
0vY+FIoS6gsHu3BR+N8Znx+vF+5rSL8XXemO+7SbBkhQVKfOS+efatYZKWZG
1q5E25FVo0eoVD62kReVG3EKndYQnsa7JczOAalhVQsLuzWsnSmtWdAqdmxX
FUZntclNBI3ERG+QWJZGj4dIkFpvFCSpvtJC/SK/XMRBlfOF/GWEQdD1Llwq
+0RUb5UIQZUTpH0Jd2LChOeBgpZywFWMRhpg0ciiuFYTZdlUyx0IWSnF9di9
VsvECP0iYlPfn2QuwzphSq7q+yPrhbd2sEV8PS0dG6i6HSu2fcIxOtpEKOTa
sgoTacDEh4s7iL03BSEzP4Pue3Ef/zrn1C33CKT5lvWP2QSLkhU5KgoBiPh5
pAWFWXik9PEBFpPxHPWFTXQC1RvSad+0CLG/CZjUkFlw3w66j3lxKkj5Ou8r
yfIqWawPwswgWS7F3+Egv4S4W3jUiOyRcsebHZRFtvtF6AGbKXMhVlFGJSPY
annQFL8r0C8e156HCY4erLrnxvR544Nnh1dr9aEivb1DbMXlcEEHj9l/TvQU
SE3hMktBLqVIhW0ktu/p76G6oMI9hrWONjPw3Rje6ocvIIVI4olExVgH8Xh7
XDIsbGwZBJ2KGJr+x0iCe7z7C2nDHvX7FS5Elx/T7ri7vkbHRSBaXsTsUHjE
MOWvRc5wwTducD+dF5jvcsdYro1K8Y7JF79EiEf7bZHCGdKsRvO8ExXJpSZ8
6ckDEkTDmmOyaORmitAM9EZwgVs7ixMC+9I4YdoJnSRHs1TTqkmnJV6B3c0s
3dWFgWB5VdtcLFW2hB/Y4YpTG4WtYoL8GQ9GyCA5lzOzbcxYtblqPQ4SFwK/
BfaS5Uh32rrm9Bm6uHEx7Zzg3VNvBUbF42G8ctSt6VvcrykfmW64iG1DjLKC
lJH51ESAPR/p1UtVgQ4X4dcOsZXZpdo8AEXfAwAzOkaMlXc2Muo6Ry3ZoUMb
9EsZWhr4AMYEIAzuzFwKiBaPAhdP39P5lKF7h0BLth19aWwMjmvKmUIFxjNj
4DxX71bCQvZ2gS2wrfuYwulV0B6Ut+vJbi0bSTd6nqtVrucEBbOFHivBcaHk
i29GNQVXptaikhbmgnYw3/h/waWlj2TYz0BFtxPpCUO0o9Rjashp7a0WQ8xF
RyVe8eMNNxvcKntm5BpBRgQ4H6Yy7+f/qDwyxYht0DHDmH96VonpelaLeuvr
ghZ6uLC3JglHRYxAaDkx5ULZpDX/WdJ8RpIJOvWvl8yktEIplyo+aCYv1l2q
IS7IEhLOOPNBgXhkv0yq+CYAlUJ+1wzAerzVViiz2gePXkkwusSxcsOL+c8L
dgrTf4ZwoOObKukd1VJyroxYA2xp3lOx5qT7BXcpdAwAtm83OAJ8EBfo4ntJ
jgEJmGp7XIkgZJoLW3Ebi0ovXK3tsiJzCNfi1nuY/Qh+DENh5vIH3s6Zj/ch
O4jB819GNP32leRNoZ6+CKpgYmCWywjtDMGbhqdqNqBtEK38Pm+AYzeLxQyx
ByF1INNWgD7rm5956RNWLjR0y+gILmnxA9mMdwBAXkmucpdKYHi9xZHyhXvf
smly2pE8xsRD1qMtpOhPZhDHbWDycfv315qAwgcmaieNpB5O/YD0hQBIxgKq
YiNXCqoU+2GUgVb6vBzTBlxKuZfQOtkzlDJKRK56cvU4rRokIvl1AMBYA22e
VQ7/IPjSKVDUhLcI6bBz7WAfZ5P/dp/GpADMe3uLuW0/QoQtV6bnz3T3uCRg
kJcN5D7s/4skC4TTANjqlfAWI+gEWXCAotoPep9PcivwPdlOsz+VRd5MWPKQ
opwsA2BfCvKfKVsS9WzC6k2T05QPi+m2EkJ15Rv43Ivpj8Oce4MnV1MYsHOA
I6i9C4lvAqOyaArMFiyUDkvQi5YMiy849wtsGGhShxxcQWkux6e8EBPgTcnE
QQPfUcZhTiMska+9aZwxJz86X9tLr1nXc1T1U4HSGgdE62SRZ4r34i+lXzAm
I1wA/S/CCtbRa2VM9/ksfpzczrUPj1OXoPCTjzI7QNF/H6FG2thAsNwhaDr0
3KD3P/8+GJky3H0O1rsjxFAepwKHhJ25sEtoTTTJYxG/rXGS8tLQ7mTrFk7b
aig5tJScCJdt38jhDK1FuKH0O1I6y4uDsdHgbWYmQAMY+QOwMEKHfbmkiQl0
GRBQwFNVgLwEEmBBGw+39uLnsrw4jWfsurqVQPYyfPppNlMRzNP1cRb59Etx
gQxL5I2QzHQi1cCc/Lg1KqlFX93O7ixV4t5LKFMiFC8Y4wbSYunNNPaofhPF
HDpMHJqmYvZFfc90aChuekkMdTaGSrIChPMvtRZhph8hKLU7rMAZUpZW3A5n
lWh1/Wb6BX32x3KPW8X1T8DTju9mLDH3Z6lGWVDaen8mopKeiCAo2s5Nmfkc
heUkWUeeJCm98v4bEijlWovKz4Fo9hshhkY1UA3hcW7ttxNgMcRymne9beKr
5yRqBtxaMGGt3TfRN4UYMfADwJdU+z48nAFtlbhuuxKJ+oNoEiosyn0H1y7r
zYuvrJDg2uHf/5yFXksQxoOnRAWPcLDKQPeqEy0dr11Z8q30VIF3L0efP8fY
QhZjUQX1RtERoXpYW4R03qCYYHETq4z4XugQFdUNwPs//v8ML12pnZ2sfvzF
ikLS3oaUjONrSL+1yqZ9ZqThqJ9GOTXGkDo4RN0YWOT/Lht3B1cYxm4HXXtu
BsYw/gYTYR84R7bIEq1Zh0xqa0sLHfMtUCc4xq7AqdyT7B45ZK87db7KcRwA
jKklT7PMcuu4gX4D02xS1nz75XLAsmpW/hkgYnSAcZCaAQDnVQiAQGZtX8CS
rHwAN/Q6UNuludlBpP1DNPITiX05TW1gCtsUkqLSEtYhY3xIeCGC5O+HZmA+
pxpdVxQFUaXnTgLVUs6GBwDLb/IDFFxLxWZtkV5u963KduSAD+UNQbmiB2RH
wKVcCVXJUlNDdYNGT8bHnyi1RyDfKJWKGLAMGgq7+VKXTWbOX1i0y2f270MV
zDb/rozille+JYHlOCY3sTfaCVeSVN9uVok1KGDuB3qeGpLr8+cXLYzPBqPF
iBpL8s9QpWpMsOSkmKtFvdXGcySR0iUEjivIyoEDWxfDoEZ2X3fot2oyVu/l
hRIbKz30J7UYpVqb4vvPxQcyPPVs1ittLpaITRS5V7kO92gHFmbMO2Qgctqi
gMJ8ufAOkD7H6NxBEYNt5jzU2QVSarfzoL+S45D6DCs7r7DHIy++bWRIfWxJ
YsVM3fqPL1zTqG2pRT0UATXJ7wozkJH/Rh25oRijmGsa2ytVcYDU9H8nXhWh
OdgV1vZN9caZ8fBd2U6DL7/CLtZ4TpAnQu/dWfJr4CVd1XCCBNsMV98CsxEw
gkCxmiac4sCDZ4fgssuqZfvSYsOzhPF1LzUgPwpUbQhnRFo967MoCdWvebfn
tO/qpbIURjOHKdltlJAwTAcNvZ90mH8mfu8zKIr/SBDZZhszT43Lz/AUq/xl
7rWeWbQG89PwAygr41mGYCuzXkWfvQYGHbHKBGp1RmDhrZdhub2poUMx6Ll4
ld8m54aD7JWFfCUQVv6hH1jL8CgaDGeYaUny8rUtmN13Mtr6k4Cmq27ZQygD
FO+o1pCG2a/Yws7HyESPXnFSzUTxIm5+DmnvW1We7fzW6jgyecrbI2qbphYv
nMb7Ccy581bKf98xzENmw0bHCyn4/IF2CQm6fgsTQoqdcDfuGD/m9qXp5CFF
VeJT9lhxIyNuozy+KDSlAp2XR78IzeOrkOI6q5Xsj5wSRbWdEYMWaO7fZoFx
7Lx8az0EZLWgYgdoj4NKbV0fhod49sqEHPQTxewUZerZW6zq0nGbOF9prNjY
2Y74dPOfFWKA2YclHUx6q1Ck8Cdnv/vAsdEQ6QCwIOJiHg30vucG1HxmZo4D
xbO9Z/4Tg3bD2lRY9OACtUvDh+/b/HQaqg6/vV1kIffJOqPafJHY6yi/lf27
vWZHY6exgyEhWP8Wrc5M45OR2h8v/0InKgGWcuh7MoFanuABZzhg/bNQpe+4
4B608yXCicz3xOwpbJHA0hkzKmQZw68KNyJ8rds6m6ux3E5MsGm8VXt/xG/v
Hr11D/8RMH8biL6pVFAduTPIEra3Sj62H4j3f0rAQbXeabyrBkAAPZHvom8+
tmkWus0/QG+T2nEcxUc8T8ENTqLo1MVQGTlUIfaHJCQpyJIv1Ye3oo3KyZqo
2Y8mogZPX3iOe0SHqXywYDEsNWh/S8UALfSlErQzBjaB+BFwxwlcWdwkQ3XM
pzyMUt1lrpwiQfTbg030jbW9nSzlPnjhfgy5V0k12suo9Dy63Tt9EZL6YzIY
dg6pGt39C6BHqn69YplGKMggXz5FAT3zHeMBwpyQ+OG3yNYhijHo7d3ZyEMU
mMCIuJk99+M3pSFtCJdorkecSgmZv2S0JcHSW9tVDhHkQ2MjPSwrihQVN3fm
/STqzE7+Twz4FgNHM1kQvdl2zRaHbmJpbJfHiABjlS5iTAWQt6vFpPiXmSZQ
4snIeDvTnaI8QNXGSyc2jlTYa+Jj8GUjdvVTfu+UWHe67nqPDjEvZ2MPWObR
zSWyoBF7S7Z1kxdvgPe+beVcFYUEePiZeselsI1yLv3belnZqxq/MkKNuYCg
3Rz0FFYoK8pj/Uwzga+nO/DxUfSqwkn8zah3yEirXMnnNfOKNegN300GvbuF
ZRHJj0ce987TOqT2Z6puoIHulbxkU/i7byofyyg6AA5qa2h/jdW6nYbNIx0B
s2lA/M65oEtsXP8s3Ra3a/05LSJORB2vi4pd5omarFak/M3cD3kqAPAobqM6
TWeSKg9o5rpylLN5OtnDsqlh6J9rHlkgJ4B3tAw/S9M4JUWkG2OloQBoZLVT
FcyJjY3UDsjBMQuiNYyKuwE3tXzUyX6Vk2sWnI9ApSX0aPrh/v0LvXld1gjy
yo5Yr6QconxqdHbk+7g1fhvrArPKR4+hueSX4xViZXAjNQ1x4AHYn1U69CK/
SSExaxE3PPX/NI2sssP68Ji5+r9WfHJPYTM8zECDAnDvhRdFWTnMjEIXJ7vY
8m0wBbe9NEhFtUUsz2Qo/WLWYqNrIcj1wKjj/EVn2XySH/PLDTwcAtJKriHK
PmSHbt0LjlKwpOlSIc1uz8C81dec++lE+30/vdaB7xx3TbuJeAb4bL8XVYqu
hqjY6yjbnc1qF7NgAzpyKdRJycblRDOLSSQxHWvYsTPtpgq3oaPdk8ewWQLD
FSPbo1avZbyEdfXITA3j/9F0cS5L7lFCIJtEgQG+5o/Yk/cwmDB25DvIy7SR
E523UTFMq5yFU8PhqlpKYVS+otlTzp0bFcobMVoPwtixwXWAr2Ak98RAF+hA
BJH4jWYGsyTN+VVala+dSJBn9EjPdHtxpDyNdQau+kAB7WVqhDJZ8t1UYSCO
iCvyHcy3mdK/mG/mZpCV40CLomjsc5HuUAC5hGeeM40AdA+juGRq/WmW5A+0
cq+pHXUnUprD0zT4mu1Y08Qr7K1Bo3U98XEo3SHB5/9x3kwuZHc9LIun+i87
vcIEjRv8ENhcyPwJbT2oSWDfBvZjix772UBZgelAcUVKg/zmfEiEL+k1ybQh
f81DVuQGtmHl40rAphoceJ499Mmi06mg/OXUkWeBWr9aobeA56VIMFdY7Jr8
ZZKJ99LwRBTUAGwAsv9zalo7kBaro5QukZVzGLMt2o50jfE3BmnYdUalaibv
sYymozKga5V8V7Q6j1VG9tL7YIdxGZdzV3c3FVFT0O8e8FLCWDdxpV1yA2JA
NesiA5nj371ndn4JdLZMvgdyKRtJuvvOEDG19jUyEaC2eFre3v3K9tMCvdxb
jRLvD3R1O7WkDzuPGsB6SWOn41MeJtL0t6DdOEfnhCGp7/k1CMcFRAu2JhgH
nM18SZkIkkst9oHvixRt6A4+wgFLW5Jf0cuR82HANsDud9FmGPzC65oxtbBT
F3iD9pC9msU0HfJ/NDUg04N2FHMuZncAJZsugZ2luNRDpaqqU5/w8vO9a9ZU
HSUIT9W4Xo85JWOYVokr48iiR1l8o9q8iFa8X9CfpSCBs1+Gjvmy1VmT6Syb
b6Jy12kjvpncBNJFjLS6Eg+gyfmWulm/qlxnj/601i6gVPYYwZhPG9GFAUd3
JkY+ORPRol7vFSdbbM3aUY/mbL/ZiEhitlZC8D9h18heXrTq2YutDllfLwUJ
pp8zjb6ZTdxYx5KqHqssXKKpWMQwnO1HIFP7Sgiorr9R7/Fe89b26bstjtVY
s0DLWvB2+P98hsozPAwmYeMKMF0avt3CCD145tW89JZYs2J2xVdI2zyHa3au
DhDIkFC0q/QMOuQNCBMMCjOgcO2x97h8nJYOhysq/w2jWHk5JXbumcF7+3pi
MtvUY1D5kLkCqPbXaeJIMB35KE0G93VOKv5lkhPzpwa7LblwMvO0i6sma+is
886iPs51R70WoBSvF8jn4G6XrIQqo4e32zrJpAlHa/9kCGtEqAKo4e2MJHW0
CZdbW4UKhYQAvgUhXLs3p/UOAdJRFd7cR+4mUZM/kIoQbvUhuuwws0naX7xF
hrj6HnrGm7HLj3y1f+eVWcvHcIp+WHsRdM4uBjjmiJbL+MJ06r20kKjInOeU
027JQRskj0P18aS0oUq1IL663iwKaiA/e8XA37UcZjVFaseegF8u9z6l92pq
4LB8aypSpajV4H2MC2e2eRAnB9UHWQKZlL9pbTIXW7kKE8eOQ0hM3Pt35iXL
Lomlp372x+6fu2tW6BT938eM3QkgqoVZ/TWthAji0avmgSF86L6yg+PM+ghl
gM+ueoJ6/dCV6FLSdVzBR47f0yVw7A6hkw2/bMuIxkyZhToU2wn8HxIxc12O
4QvajTH7ssMSN8jXg8WYPMwJSwE2mX/XXWpojVYU82dHVacBblYi6z5gR5b9
xdHzl8gEGWJL2EFQ3XEu/sM0S+HzMHHP6So0sBeXyTqCfW2VNZA1pwWYvifT
Lj3+Y2HryICiwqUqG0VI1eeHSUtQVc89R9xWmyT4bFiOaS9V7fDXm8i74NGq
aop7qW3DFQqmL8KgbHERO6/7Z/FlU5E09lBZfsIWOcWTjVttdL15wgpTw70f
OdeD3znjPmyl+WQf01zyKWVMgG8tLjMji75p6lsOQ5++gsxhGO0GhxvN4Dt3
9AJ6LEYLSF0WrgHtq0DDPPuaMuFWsvDRULu0aUoHFCTHFOuteFvZpE+NwEUk
RgZLb5Jtsi9ySHlzlRPF2Cmuyk4s1hs1/ZSLwJ72f7ZQ1gfirGGDQEFS3o48
s/mTly6gFhv8Zku28YjwRO1MMp0y3Wo0RunIMsnzI0iHcI6KJk/8XT+6m6Hl
j8aTDC1ZIfHfssNWDTwtNAsbVjQ2qptwIGlOOpCpQzbkPGBxYy/bEd9sOXZo
7odX7jui4IIqQ0VzPybSN3EkxGHBqTyYHX8CpDRDTUEkeRU8FaVuT4obnTZc
ZGBNKho2pL6yxJMan/YLYOH7yuWfPMTJyVc4Q5H43wgx3dqA252MJ4UPPVoh
dk1a9isCItQ28v3mCVYXA4EOOIP+Drw7zy/gSJ5qmnS+IReBHFijyN/NlByr
pHoFqVM2naE3Q/Q8ePB/XBLeIsrGpy83wLjZn84Fzf6UrZrh+lOVy+k9lxrX
okHt256Z152G+iM4Nst0m/N2qGYqmzwiqGKVc2wj9jwSnOrHiebxEc1mgi/i
yuHWMUdqtDG7KUWnQw25HOtgLFgak9Re5a0F+WO7Vw4r7mR7HLvSq81FDe+u
iyz0dzxT66EXrYAJfmCvJXP9BnCjr1OPNwhdUx5Rl5YYvfxtFblBhDNip5bP
UkV7h2XiTJbeuotcg6tLdnM0itdh/bdfkleTBd7BGXG4kdnt+Z8Y5cVnzPmr
O8jZY+GAtZuWGMYFBRSyrP0Mvl+AtWwKtAgRzd5yQoppJw4AV3zAQBWnvHol
BSxtjmvYoZav5i/K4m/guP18c7I+K0nzOhoZrzUHy0v4x9vbtyZ+cnKKI8Dl
XVJGSDd6JL7r7Px3Z4zfKGciRECjv3wgZmjHOU2HupcOSgRbEaO6VCasq/3d
u42ky3/tp0sS+Bl+YNtGPMRmbvIhAfHdBIbKf2QKqaBVg/xm83aUMeTyi7nM
riwVndHgMTN3nxK2JUJ3nOJ8E/7wackpUPZJMlGKlNSxgZOj010AUEFbLjQx
vgFhxdsG+VxxHkUJkBIjjBwd96ol7V6rMR07ohXKpajQ13pHRTsTKPYCj6pO
1rZ4N9zrEiz0xVoOgor/l+/o6iHTJhjvHTfR6czpDKmp7nFbd3eqruxAv3Bv
we7yFzEpOYud6ZNowx93PwCTVgzMWG15ZBHn06QhHd2LzadLHolSRGRUAgLA
ReMtGB7tdMhYd1nVzVWH80CFqwQrKhH1ojZGCiWSSJIGD4UoISkXTRlxrHBI
tKLGskFVpAsTAhAoyGwB0au3OaFNbJWGjO+FsAgVepSsEunf9AHqCiG5bwzH
cLnFZgWzp0HzUI8hDGqHW1jiQtFtShqjjI9/vn79pnNzmK3R/PYcIqSVqUki
DfN7hPhS2KCZnsGx7yAE7MeJpvM/HkthidCOkbARv5D6oHGNi0V5SIT1n820
g8S0NiXXLnvXOOzY1qKfsf1nBb7MJ7jMbziW3H3kyvN238mokMrHMF9Mmm8A
s2CF2Cug/kxDdP1Vti57DFKCe6TnAWq6ZJIDyRZsZ23Q4X4uWdvgjivy3Sf/
SOAyaS72QfA2LqFiGrYzhb6WJ7hG1HllNsqncNboYOWH2i4CC4wIm/s7a+7R
DeMxTdeVdfvY0KVDLn0hAXjxpSOv3sa4P3NyMVFSVE6KSkG9QMOSsJh3jb7k
Pw9c0NnzYOQjrrug12WZofoOkGoE3Z8DTwB8uEvMetAOfvc+YItIR4iAsxlw
SWVdqfnj4hERUJY7XNMkK+vS8NUI5hAKl8+7Xfxb0159O0fQlGVkyY6kVS0n
8HOf6Zle+Za2S5jyuAv0uscKjCwUtLdABBYjiXDYN8aGPm5TMgY6O+P9M49K
TWYaubX6wGjPaPzlTNHHP+IhWH9OXmTZQLD2QxCkNaDrcqK/63GFnwk2sbhm
zvpKHvsdHiAO7LPPgy9yNWDkHvR/ShNfw0R7AUvAerEovYXbKpxNJtK+ORff
B61mWnL4diI3e/gwZfOzvAsS17t5jSlgiA1LsS2PEEqOO4/Q4ZbmPdZyB8Lx
LDpWCWQzFyuyfK6iX+aAGOdRCgBbi4HO4ELhgbF5DwUI23v6O1wAMlk6VOTD
8xuHUq3Zsrt00EFwMM1pWAgJctOShpYXkNJoyp3MoruQDu4kjmPdIv8mmRu+
PiST0M1jekpJqNEjnap4e5RfaoQPNsesaAoANgSjLL99f+KwF3QYa6tB+ixw
QeylM52cK+clWrSL5xBB7H8vY9oSfff48Pkq4qoatU2FfffbcDyO/rFi9x8R
77dN6r65BBoEm0uvyefT39pzIa/EGMaaHwp3YZov1t/LyTpvPORHXXviWsPm
WA6JwaGx5AYtXK73o+H7OAhEN3gJbfeBioCyNnP9yaIjqBC9ejymksdl0RCy
kCASm+BgX81wHh+fHsItS3H3J6rIOvK2JKvc/oY1ck1Zgk3fzddRR4LXgmH9
WwnHgYQn0ygkhV4VYw3B1IZ6afQm6iGKewWi+RfhQT+Jnr8BRsRbBcpd6VC9
qnSuATK3w2uD5ppK71TEaZVwmsYVE3ZpmmqjxRJ+imHVp3BT2xFyzgBhDLP0
BVgV6xUrze21SYSlUL0oPhi/z4FOR49hJ7RqoA9oyxmRIu9isfVMG8SC3aTX
YtZdHxL2g2T+MqCO2lbhIMQfxsZyATxYkqrqwg3fc58YiSEfCqmdK1sXY6qX
uKZvH3Fl5AV9NIoTi6dsjuFf1xlrFB+8S3s+stp3ErP0C4/mxNfd4wlXSliO
QPyuDCw1C/cEK/gAyzFt2tZxoQVhfrTjKKaiJjN80ty1tGh2LzLEloAK917r
vwAzuCzFAoK5NSNNVQZeET34kO6kWA9I09Kc8ftDTmz+aExbILBsJ8cfaS33
dkR8GP3vVp5PH0Ur8m55BXObeln8Z3b5Giry7W00BIGNtnANhTJKECo/cBkM
PRYgdpf+2LYvyJJUCTHeQ0fg2sFDEiLaA0BeC53D59MDgstELVhhxZuSV6T1
rgo+V/sycfFBUgKYTNJUirJXpR6XkWIRaAiPAFYprQHiQef397s+oFlRdPAc
jjzhCwJVLZzB1mnJ0YpSLxn6m9/wJ6aCAin2bHXEdUju1Il3K50dFAjxb6VI
8B7dqthRvklLRaqF3wV6QHdLS9rF+7Qc+IlAKZzYZJDU4MjCW/ICGkp6OMGC
KHW1ZaNTmgNthtJpMYQY42Lq1ZzgPgIzof2uJ7zwQVL4LYGQA6GrdgAQemSG
I386MTPFpOhpo7SFhsF/tm8ZoYfU3No6sqKQY+Ufg+wjOy7mnPyObKoCCb7x
ZLbux+caRf9e3dWUkoWBDvMiFGulNw4hG6Qm8XA5W4E1EJdS1mwRrgdIsJXL
vF7Q5kkrShulocjvSt38AjQP6glgmXiraZ4VTUDxibPUhLnq3IvFaqr8962Y
/ID3DLZsU7QwzQbuVQu8Kkwtr8rnxPa68636xZeFltL4ecpXPpeC/r581YTD
4iAL3fs+/Z054QiCn9WwNM/Lxm86/7bTXrNghbYD6naI9xI1ALU2D3XqJZ7E
E1w+txOdpseNcJRNRoXoRxMklDAW9f4b2ZMJjpKQF1NmkJIw8VPma20asXlV
bZFzaLbCdB+zH1ERzBPwi/V85FgEw7Rv0j9T67vzIb/pn5h5tsdDdcrbQwOs
NefebA5CVxy/3pQXlxPcr4g0kBpA9RzP+XzKxNjjtAMIbluWKP8ujQIENIxZ
EYjC8DE8TbceerkWNMaKj/a8z90CMNl+oeOu5V3cCamTZiqxVoLwm8VcVlGH
P37q8CmTC+CKCvVEPuC1tXdDSOxF4LDJ5LwOrIaHGNzPQ032AmgFcK/KOPNi
/hCxi9WouFHL0N6iLeE981b7CvSts50wsEpXaTx5GFtym+NhLbmY55Fj842H
3aJtxq/foEGA6BfPkUdg8I5C62unKR7zu0y7tVKeGUgelayjM/fTg3QeiCbc
O0wmvpVUByAkmP9ZenAr6xu9nh5lKZk9EljQXkbgiE77oRjbGveCTmimEobS
ZOBj5uInUBh7wyO7J6gAZYQIsggGPYgyWg+zj7x+L2cZXz+8tmCRtgiGVfyW
1PYVzEvau60/VwCuieLubnJG8YllItl5wO1sbQQ6UYlmrveQah1ecaPONKQH
A4gcfCXcnwcg7LQhqjrE9uM4CGnioCinvSzO58rqGWNj+zDZBE+lzfUaWwYp
xWpxqMvB4OdRqkvTyrrKBspEuwx8j4MZxek+IXts1mRm9AJvzYq6CaG7O4xr
8aJbKqbQypn8GsL0bgUQgtRST10IhJ8LDCLG4VUfL/lj4tPz0B2X0Ovvcpv/
uvRpApTWslRm3Oy0w/hueqEvWbp3ZgoVtBsdupPEFLpJu+FLH2RYfya3D6fx
yd+/NHgSe4dIALVgBBccaii3HypaX6ACnLu2ryXTfnjH9cjG9OSAUn/hAy9k
VwRdBbBekqnNgwOo1SFph5oiL6yFt8Hgk+ihyfEBSl4RKZ0zKpvKPyq0/BAS
9eRy66NbnkqnqQdlX0x+VbpgM+2Oopy51Puy9gGDrgEJ2XdrVdNY63N/cgiV
7LZ82zwL1sy0n9aGSamoywL2050oKYLcHP5OTCSI8xyeE19TqTN5N413S/se
a3v3NsqimzfH55IBCn2zPzZUtoB8nI4yKTjJzQveFVUIpueyYUA166ZiY3Y5
cWNCdUXJSGYCQ9s8Gn/bQS/+5nptvdSjC0JvYm3V0ngXZehDbIpUWOhAiAfG
4cRK3g0AGE01zWd6wbDckDsXRiAZq8Cj8QdWZHvyZ3Cf0AG1zbwHCpjMIgC6
YBsk8yx8Gbjpyjo86NlHMQ78vteWooUGHqrr7woEaoUDVWp74c2TtjZG1mOM
VQvyBrbMFXjJTaykJQb8pXebxZXqin/uOD9BcdIskJlrlSLB6T5huA6hjv8n
FNAlsL243Vs9uTkVZResrgjK25yGlLzcKUzd0qjk3+zKMsZQMV9S+txs+z8L
asdFMLuw0yR1UCyj8OyivaoVlOWpjTNORqLwvTWkfZrWyoVfijkHFwu1RNgL
wTuc08bv1gZdAXRYzukC9xuaTb7YgpdSmqwxodtEhAm16nJQLLnVUR4Z89by
46PvB3RvaF0GXLZkaw9+izwQAHFWNZZrsSkcxwccrtVgE5ioTIeW4Ne+IwO7
z77TQ2tHlcKakt2gx15Pm7Ile2s4/tV6HEb8M7TP6FXro0PaBt866T5joVcJ
U580/v2cn8C7MiWUhLY33XTU3/NhPFC0xD7F8td1kX98PRjJ0VlXKBo4tshh
duzAQJ9o6zSbI6b9EIy6gJDc9M6lo6UvMOf1Jdb6Yh1htGtpIn4oC8DSeBqy
QS7Q/240LbNLCLAcdMwSY1Bb+Tm3UFeyLE3vqN8ivteF2E0EnYxWmTh3CQrs
SsIeFDVf3jsdA5ZizrX41XMHb7QH5RhOQI8h1NJMiXyMa3wHUOdlywkou50P
7vq8HRJpF00/kgictjwfqB1sr/EKW7iinQjQ+I/mB48211kwDnEWzVYTBpjN
o0uDIwJR75sihlX7+nWavXKdbr1JSMzYA13C+J4hyGhiaBFt413SFWYqfgSk
e1ZjmHR+qINZeMa6F6xpKUnjjDIdDZm6JlsmvMvks0VNCsrg/PmM2PYId6S1
tsqZOAqL90vRJDtYalomGhjspeCRxD6+0oqe+j7QKcdH99bEei+oLzlIbTMQ
A0LUotVG3gL4X9zsLJoAVakY5e4oDoWrSb4SinZeNQkmPeEGdDDhVHGgpndn
gqPjtGRnTgmB2ArEnF5lK7ETySms012AEUoac9Q7OztooZVOzaGHnon3cCCu
Ap7NfWhhryJoFKnKmxv+dTjIMqkB9hHUpNzlpiMNPimepOxnBUMGrAu1WNEh
DwUwdVWeqXQ10a2ExfktJgxCD+gvcizAa2bq8rTFitrwmWai4/CFVApLFLdq
MoLZaqLygVrfC0ysEMgZ5kzfkhKomR8zvjMGTnkOHujzT4nAgn/NEajeDmmP
58k5QoPbu+AD7izGE6zSezXC8CZ5+ET1KK7an0SMYxkKr+oH1J+7PhLreF4+
MqWwTom6e+08WHbtBK2om50SSwpcd9D3PzKPSqZQ/OE3z40YGmcW29Z1oKPk
0D0e0X7+RcgszRh+vDaolEXbCHbVx8NLWFd85Rr8jyU0iILTwjTlIrOFu18n
I1tCi8z6cNXHhUtlB2cKgFATDrx39ZT0piCHk2p5IcTPKQ3WrXq76DhOW/hE
jcsm6pjpHqRST4oOCDz38UUbzYBmbe+MrrS6/h5ddZ1gQwycXyalFuPCAby9
tor2Q5e/ni5Mk4FnQMF0idhugD65/Gg7sTTL20SIX6hvJswAzvyIV2ur+nrT
fnkaRPq7qp9hhW7AtYODdDSCiBXIpCKighquch1jJpfFi1bdh7m3KhhB0tIj
6VYoNDjpRScgzdAW04muVzFP64/7EeMVLazbLIJZ8UnAH0UV+ARQe6HywcRk
l6UbclQvyWEz/s7uR8TUxLfTG7BOs536+MTFEhs89iq5KKstRpi0+S9+DpME
8jVkcDyuuZGTkzCvYNatFKHEoVWwKDpBq4xuXELQUbOd+MoFg7EG8zNsFcEN
00d1fWJl6TXkKA9BeJSCldEFQ+lAlFX6SnPbegGZJ/gpUskKUgsAkIyHpJxC
cgLdBYMcMkQANrdO68scxTmgBw2znPiLA0hcjq8UGywcI+ARodrlMjLS5BlZ
pELgmdgUdA2kzMjgHAj0u7SWSDXjdYcxziSfnzSfUzZT0mZxxKLjSIOCvLsA
6kATKHGBTWuoCtBBitHDfTglRhljImQKtRudVgAwMNd74g9fYo3CChizbOe4
Qt/5m/4Qd8CjtyzdzuXjK8umwbBogYFnS5+848AKiYiifrdNfiC+v+SuW6k7
ZMqbcof/cw6fL/5MWgFw2YHa5jAHthcsWFdEqF2MK6EIZOkq3N5q05Tum6w9
a40bSlmR5P5cCDmKVqczs33HYbeqUl73hTURWPOI4Ed1aW9oQz9+Qh2Ndzxw
ZkbaadnbkZCoReh2DplQ/XMvUH1+/Cp46EkCCXmZ9c/eYtFmOH9nHtoIzSVa
D25rmQ5Bf8ugZqaXT9zXMsHoP1DZJB+ZtuV0XmeZiL/AwD20bGKxkzVI/uU4
YZt5H/oqGPx4QxKgfbNg4CjEC3FwjeNQZ9HCX5plnoSXWagoI1aKPPHpmUvX
kBTAU7QF1WKZ140i5U08pOxdNdotBvrx2v8a+YJ5vzDZ8Eh9NH+46mBW7sPD
nyYqWKSKWmoMNUbXNB4mP5uFqi9g8ADDepbc6OhpFGleSsuRenJqgh/ZUdPO
KJ1vf6fuu20A4nzI/D5PWAYnQDfswaAKi9pJBXN7bszozrDrjqe8aeSzhygZ
g7BKBZk2UoXKsLeOabkbLQCFTWb0xIkLAzZL3OwUKA9zEUiIeJOW1U88Z9ew
5614hjDK6Gk4bk+ihnQZsF26famwwxq/Bnv1GTuM365R4MrLx0HU2+8tuGBs
PlYUdSQsVuyHEf6S1uVvtG/briukD47mc32FCJqerz09VplGaNRbIWl14PQE
zhMDoHNgIqqgoUUMfajldxgffaVvGEtr805cgge0lSa8dAZDo7AMmSuRdpeL
SlD22+vEFmwO3wkwp3Gsq2sPBh2hnVcWp/tRZ1qCepFIp+96Q1ZnD2LqxKmc
xx0TMuQRa2+Hh1ttj+NjMvQ2UeAO2sLKDEhRDwa8cAr9lw7xABMUtbyNZ5PV
KFkVxY4soSUvkKrrks1Cme2RqKe7i61FY+WC2J9l7MkP3f5jjmaTTOUHG1t8
wbu5BcmD6HBbUDydWdtHDFQimMiPaAox7iwZEw2jUcWPc2L99dV+nCTJwOOO
9xFH9oIKbkNBhXqlwXCU7VFZBRfSraM4+m6l8G4VSZcgWMRR5K7J/EZqgk+n
TH0FDhH16ceu5OgzIgBU2bjYs+eFuKMqeP2C7VlMuehF2+/qgCWeJxj6eNj2
8lxtFUv8H7yC9LhaW+BIqlKjo2NoJpbqMSNGmEtP6Nsu4X+H4JnDSVEHU+Bl
+U0wsrobbwDsx2ARHFcOWJxmTglduVDyrWyHMjKdgGIT86nwp3EFJ6l4K/Vd
K7n47gd4gCNwtg0m6qv1rDMwpmdYKa5AAlMztikchfJAy9SQDL6J0p7Notke
HNJ1vfnabOjDnjIFln+MHNgKJYmsH6rI7b8t1dBpnEFbqAR6BCONhFvSGrG0
J0l04f4diNsYac/IXs3kW3BdvQCkuP5BbrgJ2NW/uokgi8aGM+vLC+Tab9hw
IVYMoV7qxSXapRU6nHlCRsiI/l6II250q6JywY7UBy9+Pg+I3TyympXvYbS4
f92fhICoMyBzM7bmjmTarBgneH3J6+bOG1eW5RXCU99fFW6zSVU9zFIZYiE2
1/mY5gkCTdf1pF3v4MIkOEIPyDet2RCzOwTiTT5i8iY5rsZnSVyVOGinOrN4
wF7B3+jRSmA9JDqCEQR5TLeiCEcZ05uvgvrS651mga7sRbN1vpyOpjmDJjIm
ap4ZSN1K6oKEz3Xj+CWHfAZ1kO2S8ypRxNb5EXqqB+litYGaxeDlKmK2EPxC
DhKPAkjmKIDS2YcU+7qpguBWKOBNOtm6SyugPyxBJJBTzZy8H3J0FiZDr8hK
mGWsxdhZqjxtCRiewHudcRKgZdThljRFGxSPZvp0Rr3Ql5OXtgbm21bOzuSE
X4ZBWq7Yk/z8pcpQzZP2VxhUWoH2dpyqNoGHb/O4G68xoc0l7mMZEW/vF9I5
WCMroZqADm+RFKDI95So19XFFt6+vzbvDwFcCau2x7t6Vgf9PvC1U8LWq165
9ZZtNpvyo7fc5soEgw0cIK/H9mCZJ/7u7Entuv6WnAmkjv7Z95LWjBb8zmA1
9m7iX67EqxI3i2b6l0n5XPvVEufE8OEUl9Zh4etb1UJ+gC/+k61dAOBt/rhB
Ua9m19e5erRDiXK9JrVDS/HyX9een46pNRdLdyAr5uf9sNweBV8yqeM9w7kV
itaxArYFdqDe6+9HnG3ZbttgFVPBDpSpCZSatx0e/p2zZR3lQaI1d+GSkoxs
VMp4+M5usp8VUS8d/C/O2cAfEE1ifu2zAusIKW1t/rYnCCCxlv7sHDnK94v8
xGBF6AdZ3zC4rLjiykE/sCDD3hSxj7Xt0Rqfbz+nr24P7Q/EVc2LS0BxSbHS
A6vTF01s3qSHXUhhE1agBv9oycwFpTuN1RzItHpg5LrBpKPoxCGqcS6wQ71z
BoAFsj0j+tMoOwcmObThKkuhAODhyjKNPLWFa3jMdsxkLcJLwsLdYcr+pP3N
VRmnbbi4y6zbZCVRtbyiyOJTaSIFfIEI9P3hcTa73HpgzZpzkLQvKLwvdL7D
ZUvFkoWyTX1D5E86GdDwd8YMVlb6Ae1cA7qtzlLlZiKYAVOUNaBLYVNPQFNG
i+7A0WfGEIl5SSq9mdPV1TK4QdFKzfSQgoYRS1OxXY6uZTR4Ff7D5WYENMzW
EdME5+z5vDwoF9unRkIMzHdwNke45NJuU5CfHTZhc6L3hiX0aTx+IaDTeqYM
rOxEcSd9ulLTMwgbfzRNICL/DB3xXef6GcxI5dCjtfzfyQLJIs3fpdUqNp41
W4RAY4Eu27fKJBe7cAnLJBuN3hjL3RGxFQH/08pE7sEdXBJZl24n7Qqk1AbS
8PIs5y2j+LGV7O2MwfO5pPgJ8VMhVvsquVpQWCkLaaz78+taMg2nNVWoo6cO
zO8+aPttKQ+rESjIMxrFZqMTjtJl+3vle+MS91Tl82BC5ze5sToWfeUTIcWM
VKrejkQIva1xioYmT2t9k2+2L5hZ8PHcVrqJ5UXXMUW06BDXdA+DZZTn4gLC
POsxYoorA/HMlWxz5R+a0+QWDk5U9Lz2m5tF5rYx9/b970BKGAARNsrLHgUp
J4XNUX8YZvBi2y10EbvIdfLgtK2K/+f2FRgk0ocGfFv2lPK4zq/PbjTzvEVZ
+3VvqO+a36ORhR39rjJVGIcQ2hCIk8LK5WO+J2rXrn5x+3b123qldFjONHtu
myI7Sx96hgtD9JcWfU8RViNsNkTTj3gutFRfOFBT+doIuGDf3DdNc317iEU2
amXOUCJ96uDlLt/wjtuWdLt2ZhGurrIqBUUrWWvyYXHAEPhzzk7o19QdpAD6
lZ9VvfkvhpAKJbNeJme5xxHI9KkX6c8u3i/ToAcAj7HpKiZPwXDIcuv9/LPY
3acjbI9Fw7P/Wug7B1n2u7xp5YTKeeGytpdbindD5GcK8w3tYFR8n3fZH4qw
wxa/OX/cm/hkFJZYAQn8/Ke+/fVcRm8XUHLUPMm8PcztNJe/ui7ionFR/GiM
qZ9evF8bPq2SdXeBcQbXNn5VlFAp9UwmpDuz3dFfyyTZ8rtsQhmop+H+ywEO
BR3Tlt1iTEHoKLrQy2rXG6oS+aYgq76DAE3S2wr3990/fTBzs9apLvf4J31j
1m040FRk5VXUswgBrSz7XnfKR5+qi4bK3qo3nn4ovoQhxfJ/cStf3Vq/3CZX
s9GGIYntMpOmq4Bd48h5E9TlJbq7Uk1QQLUiWcGltW604qXq2czYFKVxoW0M
wmVoeUqxZkJBUHTzsCj2P5g91gTs0hEuBjecQXprWv0skaX3yzRj5WkLG9kP
2HrdhI92Lqh+60ckHcNVe3UXVGC4khiZ9Vc2gYvIi2Se75sDVfMGmPxdM7Wf
6w44NziBkoyQyrsl9JUM13LDCB0eGFSfalQElP2DzbwtTilkZ5A/N6LQUfmC
6Cdm3YnT3sHgUosyNO22mMG+qRqn19kU1MM7VzwfkIlbj+hCJOqwcZXDJTVM
nrXhFl56hR+AHdRbAoC61SKpDf+VuegXaCJjwV4c8Hm1Fen7LIHaM6WUe74N
BSQgMCCQb8FHdJgYibhV71JeFD/mZGb2SyEW8EvzXo7aza8XDcaKRVasWux6
H206M/MkknZSbRVl1wa0E/r+RHtJ5mS/5eGxeJjfsSphvKqKJ9tYJYTG1EVt
0vW4kQlTE6TD4W7ytotnb/VpXTGJQPUl3rszAb0jCPj6qDSLwzNs3F9ri6Uk
50SsxCfypeNb2tGmC+yPz3VRMQ+xheoISweN5OmVkI+LtT2lIHm/Kmt9YyG9
YPiTBst4A3/UyMc0Xcn35MqNRJj7AhOoeCcE90XQl9CtpPGM2xxPDqY15A3E
y00HYOE4s+90hwVdi4Olh8xYAJSgfDfOmpoooOxsv6a7bITdiZHQml+lv88D
aVsQB+3g7lC5OSgBwuw6VwkM7Vj7IkHewSCOwLVSp39GSWN2pZ6AkjLSFhNv
qSFTw0YRbB1nWLCS1TTmi8CvFCKqFGXSAtlMzMHADQdFEkx+UUu3wUMFu2Wf
jl3HcGjHm9bRjpU+Ycn0hfSi1yRuFGg8j0clUNdHQGO2lfu43ITrvou7YMJG
k47r9RMoT5RFGlHCY3Z6XEhWcjrbk/xh+lGhZf1pA4KRArzGTD/dQ0jP6VcD
CNh5E+FYFoyEo5o3p7ZL7/onbdWxC15R6HnRDezqspeoZ81+snYzuvnk3UbW
Sn8zYk8xQTShmqd13g62/mSeJjlUy4VARghimbfk0iG8/R1n/v19ghkRbM4S
phEBV3+dXa5jEE31HHvuIuyC/sTB9WzN64P2+WhtBlIUAcbQg1LcNjFMwyIR
d89ngA0T/Vuu+eVQ8VHybF6UmG+HU+GhWJ9V9UfMvksq+KzAZtN1eaLvF3Mn
FWLjRbeXxo9o9COARpEz4M+Yw21SBl8UsKiQdFfv9FXbEibTtffHs998drnO
Qvwb/UQZWBILdS/qRLjTuaZ35T6VHnZ3FnzSAOccyq9d/quAEDOPJSSI9U+I
aP2UE6BZwpDn+NYSc8r8WiYhWscNToK2zSwbEJGMSb+c6PHc+qPgj8KI+xLm
2i3lF7biXNqw+w7hpUcx78JEFqOJU5NS3dRg0HB2Ekjs+5tIeG6iMb77/dq4
XoCjDEZT0s2UBhLIDtsClglRM1zAoOAfuK17YTaycK3FwZkDBfRWzW/koKU9
UIHONYAZXNnEU0F/x2EeeWsnazKUJacG1alQQY+BGUqxFkozYuPooaZAQR7M
DjZNZwNEeTCsmRYrAgX9QJ37dBknFThhuKVGfn10DRuFJK0Pe6vd09tRbQt2
Yupu6ptAbrRnfhEeRs2kBJjbd4Wk79jLqlYR0xoRI9XesevOxBDVrmvE06TH
TZMRPj1iQD6A6b3Jct7A0LK2U/g/zsNVWegQsCYGyiE9PfX6gwkn3B3snh6F
jeWpplnzoQR1RcSOy04HsSfF7YWTIUdfQuoMnLUFrzhLQL+Sr3uEkln/31w9
M7RO944a7OUwqPx+haXq3/FryrIKCpvkIeuR4hrgyBF32wN4Qw4LCwXOfdnv
QuFoANnaDijbt9WBB2ZND9PE9H76p1bwDxUM+6punPM4CrJQmXOwIUolFG10
2XjjoicnraIsGz02vB5irHjj6n88BsPvwJxy8JuWbngpCcuyRJq/yHPHVGjl
N7PFrQKYFXlxbCl4YSLkFtwHNoxhnYkugOmDgU83l4QTCDxjC5G5o79vmSKb
NHlQWUQiMTtNlUTtomwVX4BhEHuLwa+8pqWmhy0SY+KA+TIKw99oDorI4yl1
pmlHM69001BXF8e2oPKcIauCJ8aSvF/xiF0xfF8YV4Kx0pI606if66aulnn4
+sJxIFudLLoaQz68NbLGMlcVFp1TnNZLbR5lSa1HEw/U0Rx3PKey9Wocv2en
atjancBCg4yZnxyP+gmI8UU5LUAZ0Dg22fGkdVUuz/7d8dILBaD1mnMyXtbV
xiKNBNWeBSlFmu5gneRoslw8HFN9MdmwIjjJEAxYN0YzTTMVQSq7UdBzZf21
CSB8aQc/1Dt0Fu2fwUwjEe71GASxhyO6wInPlgLSX8CIF+Mj9mQJBNPGGT6t
Tq6tnXSScBzgY9ZSaE2rHwOn0Rg68xxMpocCfNbu92UEipHcwK0rqImEnxOH
Um6bM5PGfFmcISJH9E7CzPTUI9MTKYScnlh7pPblBesjCMJcKGjbUecfpfJN
KX4UHR8gDc9BX/Fp3PtWRZMthUjGSj5KQdsqW6FjFvSrplb1xINVlmhALKNz
23wRpu+phZaBjfy3zxV7xu9/eVkd0g1iyYP7nEWth3YoU1JHMTychGUIyY5t
j3fivfPm4Nb9FcHOMmfv4TaXcwoH+OzhiyVls922lQkfsaNeARBBH2lLhWc+
5VxTzzLJ3v2uRfWeCNP/87iJh4L/vtmgmBkguP91EwMlCGv88Qt9yAx8FDbG
v7zOj98MS38D3bjPknjboyRVcrj4L/Cc0/x/xzKlTmDWL470uDhdT3dR6iXF
oQlDXpOMfzerJciY8bQPnfGr9JwrgrulQPAh3l3xOCXxI1YjbcuVs2t1dYW/
QIJoeGXZFDCiG1wLTvvyvf0ptw/wU390J7aFcx4/flrpnWR8Ejsrg8G6Zm0N
8zbFS1jN3HJ+N2c0GyoqPKcJPIVXXeOuS02SKIsMOyzfSNCXRhRQvFqCJTap
NpjKsEpQi4QSvWuReYSHcqvjIg7wteyGDaWno+/n49Q1CxDSoBKXxyw4bXVZ
nFixji9+NMSOfP2XQxkAHa4BUAYB7OKKmoVa365vG0ogvVYB+c3OipCIiGXa
beJo2qUvhXY+IS47O9HWCdOtyaQE0jIIHVq/7k3bo/37kSMSCttMYAuV/fB3
15qQWQLyQs3oIfi2l+WPwPz2MaVOcI9sC+eZPZY2uazeTPAaP8k0dvLwV+BR
FLlh2rGPpCPlx7eSFmGpiDO3JU0Re2skiZXZaujfxM5HTHN6ofXNEqO9Xji/
aidmdCYNbmsx0EmfIMeJwDQv6tvqyY1aRkgGN66z9GVKON+9g4f/uBqmPLBO
UITzMHAZPHEcPXmwkgSfTJpTbq8PsybOfghWqBNyEql75vk7nm2WJRc9e9cN
1Vy6U6ttnoZyeskrXaVIR2BtZTxWKZ7nLIpIqT+aiUzBAeYXBaSThuEpbHAO
wxRD0xvdOOuOzUmrlL3arQp2jKdS7QrsQKLlB5rvvAE+46S2Jk5mI1vaneaY
u7gjULNQyC7fBHZW3mC7Is71DimPtLgEtunnRRyvpx5HNjOpbtEQXzZlKu2U
8ulIMY93kOMqfhCTHhwA6t3y/CicPNtb6r7sZzxTVKLQPv4a5bgPJwpnH1EZ
LmkhKvEuaWrLN4oaTy7pf1XKAt/07IObt1+8VKJaHX4CZgKabdH9b3UWx7ch
TUazvOfLmBVUMfVoh9BI9V+ECoCoDTTx1MhS0p8MCryMlvW/3vPL6A7AR0LW
QZXJiLLCwYvCHSpgVRya2qijMaR2PzSFiOe6TISvpzPp9op9tOIZr6QnaumA
dW0Dh1tO8TBErrGBQKLEM6vrc87ijpeGLnkU70h3trUwlOzvidKN2kOzUVvA
4LzzoLJSoep5vyumxQr9H7M9lpB1hCJrIZJCgiRXQLpNA3MblHeoIBZFiTN6
yvwFK9nuGFyF3H/50/2T6O5IdhwDSujErmmfFs0eq8hHAoEcI2mj5Vs6Pqa3
qDYj7lNx+fxQ3phPTI0M6Qz2bcm1/vkIFxiIMN+qT0nusUvOswUpsQQCt4UY
Ou1gwEyXUvx/SXax7j4Gnf1CSlCQ7suDvLhD/am+anju4/m8lbzDGGNZ5nC6
r1vYQSxutwzFiWEBzirn6d2NBN8ZZlLJI9hS9Xlpi7cO0/VJq7c0zc3u60N4
58rFV7vm5Wr/hDuyS5g458XevrHOKMcH/zidTpeDlP01c4GdNgSgRIJLc4sh
2D9IVWeVizntl+GQqBx0YBLfASiDezOiRBhefmnvUr0bekGsopxcENJVm/5Z
UTh4zm44A+BWs7Cu/s/TDFInlPnqIjMJ9pkeHD8tuHPpDD0rlvkvULHia9yB
VaB666LOinq3phICa7q2AoK09nvarppIhDvooTr4lj96Cz1EKwfhjWaBFIlf
fQsz0i1GxMnH2xviFHSDIYQkGMa98OLYMN0ac7KK7J14hqGEtMZU9a6sFwe2
oezl95ERN/ai5NQKGt0AN8vigoBkGbw0NFh32DMQqRbXmQOIGqaQFwmg5VLo
IQd0hWAWK3nvhrcwmx2oNAfacAKM9Zq1H+31iD9J2zeDSk3PMiFH64MeCIyG
fNBU6QCGsp6WkzakFfR4Y1+jnA+wC8ef+FGBOiLtWUMhZyvvJ99Bissr4XXx
cCeNmmJ4z0V4yZbG6VJE89T1S7YLumLK41mrOWWyBEFdcbiY9P9vlXh/7rxf
iQCR0Zx5Ao/YCcqIPMBm9+jckwkHpQaQo4D0bQ/3x6yBQGBhf4vhSEtmYpHV
WDMubG8abV6pbjrmco0IvZPxKMuuFEktHEmKu9cLnslIA0dsTtwEEMRC5gnZ
fbcsoUXMZDc3Wt7RYl7zDnnL09NNSHVIOvcx/ad0ezMIn4pbV3PLyCS9p0DP
z7JkxAzhsWWEzy1/WGClpo0yJxYSZV9A/5qZ4PKORVKcwgToefCZsFu4fyDk
/o2kqJSXtgtptPZ6nBQtCrCQPDM0GMKfzZH8PAeRfK6NmL9IQq4EuMukx/Dp
vwnhbbxIX702CLUJ4GR6EpXSJi/0mKWs6KfR6V4FbdVGa9wIkXfePLKKo26k
FES9PfHcTvE1Eql16skKUPFjNedcQtoIQyeTu2ptTHGrhNdIL78aoJ9TEPLV
lNrpCNfuJbdnlz/+FbTSEFXKSK5d83p+g96udB5s+98hCA1o9KZLrSzUmO3x
r7R5ymwQettjy3XSsFa99GzlrRYXHbJnV2uqmataRj/Oo6BBpWsXK19YQu9b
wwCUZP+WYW7fSOZd1j/oHl6N9/iPJ3yllSJwHrGJKK8Ow4jgTL3R5KGJks4x
DvGi1+G6sETpb/AzMpzVm/M9cUxxogSCugW0+oGEpQMQFmdKZ0QaFHM+2F1A
A/hloXsf/zxxBSJI2HkbrdpaocjXTjtqJKV5Mv6rUgn7Xx7atqyS+r19g8Bv
nAKYCV6hVAYwq58ITFXAAz+UB59ScNPfW4FgwpwTBWfgmYcsvMTwTl8/WD2i
HLTINCGA08D76rwkNkMj6SOVgSc7OrCZYeCj01y63l5rhdVit9HnUGLl8u/y
L6jk6vCiG01RCdn5SaLMOgYXNs5P5oZVMkJigUT6qQ6EkhEpRif94I8z5VLt
IOuSTxqEDRimJxgJD6iMcKMp6+d1l7H0GciVrF4ID/SyKmg4CpEq99tfVGau
fCEX0dBibzxeLh2s637KfU7BWFfiJRk5OXzDApiuArK4gjTGthYaSP0cOQua
GQxCb+U0Vd2FQc3eBv5GHeSPwwCYM6OiaKlPyvdct8Zu5eOaKuHrj2H6KJEY
fe+8yJmevDTcZc9Z3VG79KeTwin3+6LUvVMFYmnDtEOmAS5+oXPc4g2dJtHB
l9rWjngPopZH1RW9Y0ozmQZ3S4FgHshwZZdK9WmNBZxYbVygozTKMg7c3z1a
Aj8K7ARsRIqcQvCSjksdrZ2NG/xUrd6UJyLrmBw9GGslYGC+xLCLa6SenaJ/
C22PkcJotWtASO8EnmKNJKXb68j2Wn3/zI9B4hxs2OEj9Me/vB/RoVLCLa4I
u0GFUKMB4lSXjbKW3Ow3/NZ3gHzCdkDC7HVkQ53ZJCdEK0hkZ8hxhnahtLMA
KRgoe8uvskf+tqhBO09H0QSkEuwqETxosEo5pyNQz7TWv1os+JXh2tCPoOLs
YB+6scplfOodCFtTMQtQnQ0IDwiJfoL7DCkARkMlP1TMoHVTVEZH7fj9iYKq
wrWx5WOYU+qftmohKLEGZhwmMHc3w8JeTDl+3ObuFziolvuhyF+6i4f2c9XX
gqVZc3WRb+2xVlx3cejwtwKjw0GnMtCVMdU6cHrHHlkRIde+NFdsdL8UOgtK
7fXFWVnuJLEnpF/G/AnaUXBXpAV4z1JgGsZ2m8efq0ZEWADccyeh+f7DkKcE
w+WkBoNNx4/qfsUvMC1cnPzBMwIeC7XeenW1bfV14dTATGFBNoQ+v304SOem
QOsTEXpP2kAheNJQu7lr8aKuGH6fZ9wQQNJZMGNxReKPrhFCJRvK7gfV4dr0
sgAD2nM8dyLLqlOzHFh/DB/NvS1+mMFObHti45DroKmHoIfQ87fhvCkDqLJM
ovSx3p3aEvfgDv6YOlBOvknanvbtuzzqvyRbDp8zBmX9QUewLZkm73N3Plrh
7MYrYs+FQ9vDb9gKgTKDu6gl267g1MVwVwrLxVGGN5+fusP39GrD3NQnEdlM
9W2/8u+ecvkABezHZdq8U+8Lu85xklOifTySOD/vRcp9LqePztimkZ8Nbw9I
9O/0TjtA6+cpEowQPKJrVhZze079MF/onOEWMqob7+pmsdoF2WCNTPpRlgFL
hoTKtmfUmWSFpSVSeMZ82TCQ/a6t9MxLR0BuhqrzDCVIEChz8OhvlBJ3Ratf
augzwPWbRavzm71D3vQ8NjRpkaReohtxNUk+t2WaDXwoHC7XrIopjcZYjE2q
OLRUnlyp1ft7rGkDPgqA4ChRPXh3hKr/xk9jXbe3QEjjkxeY3AJHEjJiP2en
IJQkpHQOcdf4h0vPKskddMl0O50Kad7wzSmhcxK8ge8Aa9v5tLiAyWWe9a1P
5ieTZ/wPZf1agdtE129vMZWjH4rEyYjgcXkMd4k3eXUhfPoA30BDEd/9cfUH
6bYIKmyxbqk1L76b8cVlgFwbMVg5Gf9b5Il6mXxdtmtOKcmuFgnZ1WXo+6K8
ru6sISGjzL/z1fJMrk/YhTGq8GC7jQ904axSCz3xGWlu2XCB57ArHnGyBR3R
3RjVM6x829YjpO+dFLS1DnuwswjRfhb+2/2ZUS8R2WRZmdmnd1AaM8JvO/np
CngofhHKDLad7ODg8KlWLdn+qrhzgKWGMUxzbA4vlt5ukxAakgPKRiOWdQT2
zR96ql8cv5VALT+UzegRGCzjkWeNRixopPpF+U1X3CKwbDpzQoGxE6qFJrcc
y9ovCIdNjUHX1vYFHlxX5IF7nsbXw3scDvu4Z7Z2JdH+kbUMiFy1bbCP4gLB
8HyVWuGU4apfMHFKNtN5MdToIRyxBV/KI6iYWIwKLHc1u4hqohiitKc5pS/6
Y0v3IrQ7J8FgUK7vVYi5pQ+OUMRtIfPaUj5jRToDhGMlnGFTJHtq+W3o0lmV
+dlJ7YQqpVoR32ohQr6nzbg3wOfaQh+4BBMSTSLhXy8hpmITOT3BBiQjyfEj
s1FEGCV/tfk/Jve5lbFr/x0mMZJg+kM/ZpdpIWQaVfT+oN5PP/90pFn2sv/r
Y5rt50Rvedsp7UNVjEhTbkqp/yfFWylDn4PNxO7NVAokz63LvWZoYn8E2AuT
/95nKqpR+lO8I4FiIbS/1OxfFnmi7KZpEJXXUAnLgPvz5FaZQ7HK0/uIl/a2
D+cGZwESV5yoQqSk/giwrErlw2I6Jyt1kFB+OiTq7Entg8KwP9glIugYEkbX
ENaJdHShyqv9BwPm8yb2ibDQew6rwJ5NE14o1s/YywGb2HArLXmKiH/WYSRG
9F6OcMLLS2n/xg0yAO4wbrmzURUXlJzfuH0LGWuZpRYEFIRBjNMDVzuZx3Bf
PywdLFICXXR6A/w7uT/0E2PzvxZgx9rgk2qXmiCPWMO5/rZ7GtyU2G8VP56G
cTdm98MEUUr42TQAFzWxBu6RR8kmmgiBa3PYe20/WsR8D8nsdEZ7KLrLqN/G
pbqiIucTO/PIFR3/VITWstmT1KzkQZnxRXu35nrbuf21atNiCzkGQxrM5DVx
1fptJCFXxxA4XcWHEe0ig0DkacwA0P2tTLfiULwUH1xrJbmT6CVJV5cvBfY3
6yudXqDsV9M2H/D+n2SnmgHXk/zCg3TG3JDuuFlPmoidlZH2u7D0YBDJekQc
4heOwCPrPR+/JP0RC6hEPYr89VfMjfouGVGQq3RhMOvIjQZEn+At6/m1dEkH
Sv7V+S5Iq5KgJS6e1U7zuWftrzMhG2Eg1UsXD0LaiRVIW+08WSB6UVyPmL17
8QjLBbTRxZPqmunXkH3AlnBp0mxCpf74ms3udhW0z+t03U02plANIBqsltk5
bllX0J3tyO5wHeLgycixcoJL6xsmyr+5j5HEI+O493vHCTCDwU1+JW67Z+md
2upaNI7HzP0PgCUR8+xRjJX/tP391qsLw4CQncYxau0H3hOJdBQYmIrr/lQp
NdRTmS+wk4UMkioQ6eNwXpMOTy29vwuB4Dc2GwZpw95uTkEaUh1ElwL1Y7l0
vAQJsHUItSJOkn5isRcQIiPFyEsIA0XjaPmO7gP7cvPcON+AxbiA6idfdhqd
RGgt28/z/E1MDUZ/ULDKA/WAIGOI0hUtJK+93iETnVdJ8uEWumeB89JcIO55
ZzOX8xjVF3MQW+BT3EULt4k+Xl9NkS1t1TD9+SBa+k/Q3LDWofe00d2y/l52
uQitvqaxH1uVmcPxH7CtK+tD9uz1r/NMi3MQm55lH9f5yK8gCeyzW8pKWVZu
ZJ4oU/kQB51ucjnnHkfCsTLtE3O/CxSnJuUHXFw6RKq5GK4t3IHRUOI9JfAA
vOV3hfNeWNbWZM5RQ/sM2MaHdWjvzrc6DXY50gzUXmtW1hcHFHYwuQEk4uJk
ksGFmu+6JVwIJOYWzqnwts/21i4tdO8DzReX/j6SlSsLCPpZ4wuxJV84Lbbg
fu8e5N8TxovqXu1wo9PerKrSkBlPCmzuig3A4/RFzomuEy233dx0z+jNOrE8
6e+1zMcIkeNBp2mDoztYnutEmPONsE7jDAc+IxpVnU1QidFZskOaRAhTglGi
669LQhD6kWfJNsj8P/9pTkYBUVYUUoRvs6C9E0cIPV2CJV9XQvAdpWWiI/ak
YIy/VkPQR4qQNz30CQSy13lkPqXw2CHpqegZ+jbo5xAzemU5sYxcmQlfcz7R
rofVj0ZNek3qu4XSekiJQO/F457wNrLEM2rEltF7pr4LOBdmwkiNXhfImCkx
IPi1CzXGeoq8nmCZNaJgqWmXyodL7Mxw27UKE58WEmRPt6KtX/UUcoTO9sWv
bobO4iIAd4OXCk0Ofkl4sE4EGDXxgDmcmK/c66SYM4v2DH+4YasLw6gB/E/C
XeaYQmAHZ4/9/KTBCA3AaepfI7uvgfhUzmmEVYSG1PiswQ6FUkXBNXTTZ4k3
eQ7MviPX8XjCXO4NBY9mOyvpF4I09sNLLKjIOBTUJnoCw0lNhwHOZ84Z0Zbu
2dJlXf5o+axXcGqmNzZnQdcTNXzNUEmRczC7XsO1P6HX9PrSJ4SUxWJKlh6d
IEnOsCm292HhxpHO4DsfD5VqEuFExZez0Q5WoMNEYSMoNt7CjgEkV315E52p
6P6Sxv2LLaJxVYwaJ8GQSbuuwXjJZWiIbHIHOU8Bjt8JRHgkS+D5Xd2PFduI
B8X6jdQnh25Bu4HB4vEKmLZ11pH5JKwbLZNTWb+OO1VWMlMtp9Fy2oWQ9Qpl
CqTntsFq3LxP6iRDfjI2VCxjO//t8xCAc/9wZjrAPwnXBaFqmDrqCCpjJHP3
WWVLkb8SoJj2TOGXUwiF77jjWGvr6s8zLV5D3fICRkyU9rkOtMEsVNDIfP0w
OELoL5QcNtPCQlKbldwI10zXmr2txH2/ytPunnRyYYDjR6rtnBjdT/jh/4at
7tcPl1wEGwYGtIVJFauAg9aZmZ9KFv+CTzHtitwAm2qTQuH5R/pztKrqTnv6
Vxjv39joaB3TMPPPF7yYelO4ZYpFtiZaRaroZkq5YC/PGRkS+1HiWoBK8tG5
1YxfWu2RzuRNOWBlV/kLWkVqEFRSZXGS8sixjRZgqLwJ4C5yTN45IzEEtzzD
lWFbzGb3XNUrlt4hWdPXZ2l8USX20uVfhf2/7Wzlx50+knbE058SWgATYt1a
dUijvB7KJrZLmm7meMdkWHXCI3EyVOc/RyqxZO8tl0k7x1d+RSHhGtlbzGtp
wVss/YoI21Ugs/IL9Ezdi+FWUbfQTsKpJ9I4QLj+Bka2xDPNyWu+F1RViEXw
qA1egrpCwum5bVMsPMoM9smRCuJoEhxAbH4ReFIvyg87IgmguR+xzzb/P6XE
gJPoItm4MBvi7fbTJGBH7Hjh0ikfezAvY3nxkPhKjsAe8DLjHaSPhSDUih5Y
RC/quIyB548Gcv+1GEwu9D/KKFDPju+PxdZKmvJno6Gj1SdNvuRAzkRjMLNy
sD1aNIeDctxcBBXtFp5tPzJdEJ4AFFQaVhDAyD7t6LUd3llfu0cDiIhcEH+p
p5rFbYUBeCQFLMIDpg2tjXh1VVs3WXN6fcnxZCWoLMKI3E2cLotZ48stVA+J
kKvrLBI0MP6/0shYuoiADIgwKHHQ7Hs/AeBWwcbRQgmEYDHzeZrORUN6TTha
oQZpUZKFKlHaQHDJOlWbqsem7W8cik9H5ToDpNcY5aVo54/qMojTiS64FnmU
T1NenTXRUdgLgdEwvUlNAEN9PVwzwbpx9+/z9JZk/bDKf3W1IIWMRJUd+aRY
dXpRSeF8pyd0/2azcRvbP2Y55NtvIE66LkJVh4Nv1uem+OMo1orSZVwVjbxi
d3Y7L86E2eZYomONDnaxI0Il5sLcXwFVSSvlZPMt3e92Tpng1JqyzCEIxIMM
orn4D9hmN4BtF2fqpdK/kgPG763O7uRGFWc4/y4pFg1cIYLcWDzWDFctFmG5
tvFjkBCesAB45QJ9zIxOD6ZAkd8PyGGao5SU6HSGHIkQiuK18HRqoT7GS6Ly
TnNELu4329Q/K6zfwYrzspFObGKT/iCJ/NZfo3DcNPKsVx+h1XI9TUibhbOc
9bdD432XQhhk4+BbdsIg/13gDsE1xD+kvEihFXALuwBq2QyOoqNcpXDYnwQ3
rdtUAetHrl2zHkxbh1YmOHkwsXmYs1BMq5wgPMnOuZiis4VwzPc+9WJcRlSo
nWS30owiCtLNS+sMyUMEpMb2xe3dTlyGdc/V3GQIaWKBR7LHBT0HSbdSdfCy
Hn/JJIqAeJHos9gMchxXdleHCbRnsS95l6GiP6SAvYqZokcqmzEiOXDejIhs
yCHvmLf7PtR7ZrmJ+FYMx4TApQJwv81/Xk7+wD2QlWXqhwo/CJTVpInyZAl0
UTjBig4F0p6dLAZ+6Rt31w7j0qH566KZIqfvajC0sg8vIOTELLqczj/bb+q5
WOtQKRzraro/mGjxLByTxoLvYTAjzbFhBjUW1xy9ZJBz8FIgia1W+25SWjMk
IbC5UN2i3imQS2UmdnOY0cP/zUG/Z1Z9V4XLb5wd0cyPao/Se1jKYKhaWozv
+9SES9xtpOg5HSVFGU92OYKHYf6wo1e2ApPjAzUiFIh0Kxd0kZH2R7iEAIbn
B4ls3mv9u/46ZbAhQbE9c2zYbizVQ0XKcFyDO/qNyWvvNULC/ATgUR8HqvSi
7NhAso6SBpwd4ImrNa/lK4gRXVkXtuRjS/Mil4eO8+Gl31iG5+2yh0itHBsI
9ZwVcPe7Px2MTWCBIh3zMcgMp6OLt9WJVOhYpb8A7QQXNOBAQle1OocLaKhB
Xpq5/m9wotfIRNx0vo9DpFdUrOnq77Gzq+YQ4yuy+3KHm3hvsnsHqEprneNa
DniS6hsbvChz7DXMoOalGNIsr0Cbhvyd/iwy4BUeTYLZwThPkImsrcgIZZOV
Mt1dznCxnn5DCTUjj5OIEZj6fGMj3sN82PEYMXhzSzEknjiyBAX1oLepUoyW
mtrVw1tSPk2hkFXpjXc2EJq9ewSYn9aS4bMMJUGJcAcZppxqsUuuHlLDPiav
ZoqRQbYWRhbC

`pragma protect end_protected
