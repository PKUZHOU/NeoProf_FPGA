// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
oSXpWzW8Attnh1K9ttBPjowNxFqaIHLdNkREKiO5vKO+U5f+rrt4A98jbvZX/KOa
VEFemrv4/PUW+BqgJGgl4cq9EmqhoIszV3RD3nhEYAi/3a3o85BalJA3h1B7CMFS
nGyBu7INPVFqeXJ2CDamHJpV6K8t8JgYA5K46Jm8TF8=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 74400 )
`pragma protect data_block
XyOToV1GT0MNVfBzthhTuKvLBsCZSDo49AmdgCYUDZ3PKAFJK7ov6mnjAy1bk2Yj
+37+AL4g2vY/SWN4TmIZOS98V6fTT9kC5Js1sjjTIfxNpKRYsaPbQjNjjgLzNnP7
XcCqHbDqbUC2OgWpRhtHky+dyRYj1iWOp1lCtI5hQVX8Dv6d3y8W2oSp/tFK64E/
sFaw6F86E3FbsZTtIiy58Bvg4KFMAImcXf52dP5yR09ujS+v8y76jn9bup8D+Sm+
DLNtZOKNcJoPilISezwdTKdIyE/Pc1FNZ99sqjZvPrVEtvnjDaIRALCSACREjYH4
dyR9CooB/lnUgQHKXP8Kut00pND07jajf3XTlNhkfQI/PndRwaO2GRIN9ePaiB2t
ocibxmxuYiq4ECxVBtK8dO1TbWNvsHswaRjucw8hishvGmwmX34GmdNoS/rgf7Jw
xojCEUEfTfVREh0yTInNoRkzdq2GhdD6O8BHgnWx3hxbp8q9ZHexLIexoCES7V4I
I+AusLmVApXfb73gTTQEd5KSt4aPIp/wCL/5kxVLklF0xgZ7YKK7ZzafgKV0WCsc
Jj777r6luloTyJzLqTdVGHqX9icsxu6u0MkwDCuEXh0Oc9guCN1hOagJ4m1zPSfB
qKHmeBmciDpWWJQwFo+xen/MrZ+CgV3hSKhd5cEVUd88BxeoAOVt+1Du22r49K+P
5FrSPAfrRiBF4tW4WaaRFQiZDl9fAzXKeydOG43+w54Iu6qHsPzugpMsfMofyVJv
Z4aBKacdd/0r8B8fT2/fH2n7w2cTRBCuYjN2ZzszgwCIXjsW5p527o3cxvbhzMa+
S6Ai9+WjSmyvkjVp9mwxVVXrkX/lbAP1cdwMcY/pzK5xMgsZBik1Ud61NOmHIhe4
KzzrMd7dZVvRdKbefPvIT4FYuaTTO//exMvL3YInzS4oj8qOUg7zMKxzFBAkkJuK
GG1lmr1gvXVPtXNs2vqjkHsAAIVtcjFMA954UlZyJY61SSiGTfay1TnQVBXK5xUf
BBh0Gn35XgxRcI/ULnPVm64ixyWidLH3D5bcNYd7KjIDCyU3SpfB4W6o3vNmOdQI
VC1UGza11gDwUF7wziRxzRswjZItfDCAeG8qCc0EvVnT07rdMvIRXo7Uocbo2zyJ
NQC/dau+QQxR6XAOrYDdFpxagWLZq0WM7eGi1gFwEg3SgZGJabaT3bHw5n0LFoFc
CVGYpuRVA/m5ieFlUtuNKr4HZf2ZpXHllpd3PGHZUI+L3M7IDkHUE7k7W++2uvza
PSdz/Cf+Dgzev9dhbiVHLmbrh+VO5KVUxcd9IEpgLlOKad8ZTRiLMNyElrRuZk0Q
2xrorvMZvg4HSwBWJLF2MOQSXHvfr5KNK/DhW8uS71pttCITGcONLNOHSwO7Yx6f
w+1Jt4BJGlFF/zde5VsazKiLjpXe91XEmgfjhQJULjnnekhf4b84UQUz3VksmU4E
Jn8igs6n0Z8w3/3zO0FVgtKcjbgjhtL9MGrolL9NMYrQGNo1aG1qA3PirKYTlczy
C9qIjDxE+1IB8VEZZ8PBYujF/aPIjffRdaFS7p6Z7z+/+9YZ1XKDPj8/XUOL2aX6
7lCw+GHRzfW4Jf+AhREgVrfTFNjayUcM1N46nFNFA4yRLa0qE3ef7WKb+1DU3dem
XbKaZutwiycnPIwgjlCMt+EM9GWNf/SJO9QsBige591RWIBl17bHiRC1dPQEPMMb
8AQIb969Ugm5K2J+hIGRcXO0Xavk+lO2F9tMHIz7El9Ho/5zvPijqJJLR0Q+Zcxf
bscfZvj3QmeHCteCqY0tn04g14+Xq5U0A52H9wqvGzklE6pAxcO3PFTZ1h4mQdjx
6ti71SqClro1DmIha3pkshk2NrXncpBBKOZjsxiyX3AV+sw+rRfDUTUL12IUsRyG
LZgmN/dGsqZ081qltbGOFqXO/KhRamlmpzObIf5DX4dquBa3douKyW3T1MKe6C79
BBzJQ1Ih1Zdb8nOBptZCuBY+s54zvyp8246Z/lmmYn+u2stUQVzngbIMxP/GihLj
2yQCu6/FMgHwUMFxQXoehUaKgg0hIGgr/Ytgrl7Uo2CiWXI2gFv8dto6MERQaVNe
h5bMMYXEX3Zt1FK1ywA8J3P3Mhq5b1aodndFPeBGRM01o4AEbHQaSso6aQqv3sk8
BP0nkcCmzXKAKpovNJQYixSGamutJlKopcQ66yXvxE2eDWG0LdSmyOGLDkuoPCnk
/volyATnRayGaVygIUAbzNkCB88EchOPdNfxYCX5UtiA0dMw2OTxUi2dSk1r9Q3C
FMnBjeYZsHjhOhUsmkPNXpTCj8BlGWQI5Gqwq78/UAQGLQqwyplpf3tgaR7znnel
5NRY/NnqPshqlgmta10nwosCJKE8UnfDRzCCEVhj7BawPLXSfM8QM2yXxv2ZQmpQ
fdp8qeWCXSwgVrT52ABBkDis+haBaGZ1vlaTpiZq6eZe/4ZYYPSp8mxam+u6QTdd
eyYvt6vfFnp0EEVYnUcX9feRT3VDaUsZD4QnD/CyptyR0qzPmdckicqhLWp/pNfx
89NeDStw7Lw7mo5WdxVGy/+FwOOVMZE72o0R8t6/6aWCuM564zXWfGhG2HUvZ3Oo
GjtbzzF36GhSVP/7zcAKnn9TlE9Z9KKABcFzgebiAmN6B6SYw2gdm7c/l21vbU4K
Q4LrTOyJOx5ZCUtnn4hCm+8tY2uNXDoe7h/qt9Hf0+9lkF4ies+4HSj518r2rSip
7sSMezxxUxfq1FhiB1P8Mv2GrZsL8tou34gjpJni2gVqaMl9On0RBNWVMBLPLURA
BqhMlYF7aD2GJcnaIADffrTIlcs1RBM3HlSUngHvKuH+ZvN0dSimDBPuR0wt1gbV
H2fZ18piScBLT+Z3Ju2jQ9+4lckwky96wqV1oG7DUwBL0AJ4ldJijaT8J+FiCQNN
96ovEecdFML5UEqDypTcNNqIO26AGp9GBh38jevq6zSWSxZ5JB8KVOQ+EtH9++JX
01KT3c48Zr5qVjR/odriEkpIzzIHJga1bgW0+5ShO2kk9UH2AIDf4R1aRJvZDiHz
MzkhvsdwAsUDGVHnmWDFpAS2V7PJSn8x4vPBiugeQp3psFlTj3DNFSMZVJCuBFVr
PbxjkZWSB12VV+CpACz1TQ2fUBFDMdXvI1EHQZ42Y6AiES5QqXboodZ9BEUkDJnq
ikrQObzQuaRXtySK8ougCJL8mEk7OtsZqGEJbQSONyusML6QnebuLjOGJPwa67mW
QoE1J4mo3j7boXKyL5JZVFf1PoRSJniUrs0d8D3nErkM6+iQcjx9Rf0rxcgJ38dP
mnKSqxwqjcnoCxx7uHRwrPYzlLLcNcDeBEUaHvz+98BDp0Qo2Xctz6p+nv80LLHK
j+5wEOb8XIHl5Z0ccBed/lRw3n5pTPwXsBKEO5bvjd90qRlgEaW1FauwKmx58lXi
ajng+EDBZvvvP2enSr9wSO/xzgF1E2N9Zh3tSa8RCxkZ1Er4/kOLHhBQm+r9FblO
efV2ho1vO0yNjhOttwhEaxamGPVrSdrv3A9QJxAELyPfvxHu+cGyR7FAhngQqphw
EG3U8FoK+WzAphEEP3SaAE3fH5UEA4j36ozzHDx/zw8/oYYi/X2TTboDwGBzHTea
XYV4D3KHjM5ki6VLQIx7Tg8Y/hTQj7OZhFif28fS6wTmxcSrIluR5CO/VLojpyRu
BWSfU3eUFnutonr4R8rgTe73KQoxd4rhytB+iRbjV4zkNud+VNL3ePZ7RFfHFzmN
CMuue1WY8PdoLkhnq/YmdKzDucun8o3q5ebSm2pVXDEsOoeoXjCSXc8mqg5YJ4A9
U5R2VqEuDPnPmU5+zWjLC7zRXmkbqcuhbafPPedJ1KEk3X+7XlD8SPj1sLpM3VD3
YnqCeLIPNGKyNqLIEQ0iQqMG1D4Su/aZDTml+LACpM987GHuuRvj/OAUWV78vt0x
cxubECCfB2kXqNh27gO+i2iuebXvHygKBKGQmMTom0wp+fDSQzDoibrFqIjPFNcs
Gzdb8w/2IrSF3xfvyp+epIZT8/+pRTxJE97qPHZVVXm+405mTGFlG434wvceIQoD
ETZwYWggrXnMzcXECjN4MUz3AH+K5BnXYZkBjdxcygFmHA5u2ZZGyPzeNv5FYTdL
ii7PToigQizoMhtCehQ8nXIUh41XyB8hidkhgu0FUpUUEqH3o551z80TmygCoZk1
SOdK5Ari09w5I3P41BlKA4cW8qwgUAkX2ynOVrdkDgu6jSR5phYhvrQ3W51EbsKa
O0trR+syoeJTyOVsG0wzRLffmgFfYFtPJjYS9oSf9RI+/9dhLw4cuKABKk7KYnl5
yZPke3WoEctHCxNQe/wa99FY2Co1Yw1hDlR013C5Fxwb1vXRpB/IBYm1O6ZNSZw3
wwbAvp9eNPyanQ+Fb0A4YXAjFQP3a37YEpzG44+LeMGmT+QpWHqYmMCaIA/b3MMm
EZ0H+bQruvNIsjHaEml/V9DYJoIAjbEHrSUrcJ917DxKM5plafI52RyO4eIUwW9V
rbLrcncecQQJuIL0wl0e284FIfIALCIkVtKFSD3RU1+VF03aa8jEFd/saTG3cTXy
SxBc6aCwqD1R400u9xdbO/Dv0JE020XPbjJFTBQekc7tci1BqRoo02evDq0AAleB
SRViYXQC7thWYUQKS1HlhrI2dNu7KC7y+av4m/izqoNan9L4Cuc2v3Z0HebF/QMW
eg0m9/NH5A92n6yfjOyr+h2Y97GoW7v3P5FrjuELb2rp+Am2xeqLJrgJHbvr37OB
53OR+thKy62GhxtgdkmziNdQzRcGp8/yZnC4YhquQSnTBvP0mlmGu5mQEdNFbvnm
wcjCmg5LkLK91AntSn9xNmI1vUsZi3ez59YSVIgknrJ+kqcr6mLAbFQvOq5BWgoG
O3WlscixH/pLP+Bkf4t0L3HTNV7J2fSnN5x1BQfV5FuzCU3qmZv+uFzbssgcFz+A
GUvKXcLrQ+vggmmje34rXaf4MrI8Y/kQBfYJXSYoE5HLuWgKIOKrtdvKqbkSZMHY
tO7ElWW/52ZHQAip1s9Ol7kLX3esI+wpHTZc2V9IHmSJcDJVDge+7ECYLdN0gloD
hqVSX3fX/jCNlguHPLzeSA8+8kZ4WB3Vc7Bh/rOuGxuqEvO/xzG1ApDw3X3T4wNR
1yA6o6b0spMwoLwubmWdjDnKhUK2out2H4sPcA82gbNRZxZdCY2FPDTjpGyIso1A
hBAlJSusP25nDtK1fGJzn5qaRcIIoNrJpaSMJ0w/9NhxCFtEoQa823E6xHBVIpat
RQfQP13+4MR0z5iLZfb9fvs+KoIEm9lZ/vj8A3fmM7ERFC7uDlk8W4u5XD5zavWY
qiAuuDdBiVQxBBeHHkkyYWlj3vr4XoAjXIeKAcXPYi0KLkA0xFedhsqTsHP1RGM7
7VCq4kBlGKIHdhpUjAuV0auCtkYaZUGd8hNPtczfBpyqTjCdX6sEJOoUPhwt7GZa
KWkhnI9k5SPFUF580PdChHHlcMLi47FGe03Onqu83x+toGGY/aGuaxoMBf2yqkN1
OKT2BjQqK5hDJX+QbM8FUS2MOWugE2N0BYwsx+ejTFgX7TtfDpAR00wQqwDD2JMl
AfLC6aIPsz6ZeBlgVJRPLfGCIWxngWsy/OuY1ZpnXKZrPMgx3n/Dcg1k+7yfGOpM
XjSfSCsrcpnwzKPoLGF5alQyshGosCqcqe5Vmm2zpjcU6/8CPRkM69FuQvjrdyfA
LO0VCErzlIZxhRf6mQPmZs0TQKKWba3X1+OKXQyKq857r5CGwQX5N6tSnEroK+8J
INRW6/PaS+Ffy6JObGD7R5iVC3qm275PBUpuop3OS7HmxPCRHnSOamxnGr6dho3g
BfIrpjuFJgsBi03PdE5KOkHgr2sCmdR7TWF8+tyaygzta4XmZJDtoaA7nV1PPvtZ
+t6GS9nZ58h60foaXttpt4yf/vvsNPbnrOXA8MStEhlEC5ycQ83NtlvHdWrCQpLm
cP5v8YfufMQYqHdSJegv4xgvbDS3iL74/o9K+DCEJ6gQnnVKqqGxWdREgvEpMTGx
2LAL4mFk2Og9rGelTyl4oCqKFTWvKuL7DDaZGNJ3soJcA9NaUDpN26aDEF+yWPEM
txTOKxiXBsQgKXPI+94K7GySNuDMN03tZyALXq3qdABKgJW/Zb//8ZSpX4Vga3J6
SgQIC1+TgKZMe8cAmHdQN0/ieHWJKr16yCvwDX6YlXFqXhLbXgev++yT5aNsox5J
79n5uk2eG2t38aNeW7GAtUO3JbdBRim3yl0XYpSmSajHRXAzJCkpHIZUdQDfLs3R
rnWy6/nfP9fJaWKDhdZXaddDGaisQjJzTbbrQ1jiCRKi2/pA4UhQuMZelh9lrnH1
AVfmSh76r2amMFII3nWfIXptP4PzV3Vbw1i4lbo+LXX2wG4aAwvkYIJ1CQKsOqPZ
1aCLuD9A124jSxnw+ivBqgmItdiCdo3B4Ko9QNI6uJKYxAlX4GJL9vjfffArefDz
oKUL1+5E9YoP0uPoS2QCTwKfQ5jEsq5E7wjRMVDAJSH9d59Ggy0SFTJKM3n5g5Bd
DevLfveVvqhpkAPHWyHjo9XsfX63mF4wdE0levqvrdN3EdjKMHSCkwMYQwlLSLZh
49l3YaWPUNR63cOyvj15Zqv4RIAp6x1DEUO5Tbx0a3aQNraFacIILjW4vNpVKGsx
LM1f7P5sRgSs5UR66SGG0aCtY81iuqM44TaSjdVn0buNINgdm2QJlWXVgPJm9CLh
exq+1ZZd7kxkeVw50rIM/CcQinXouDYbgbowpe7mGlUzhdwb1G7jPYYcPUxh7zZg
CT7fF+6/4SZVPzIEgARWSfxbV5gDFfTDPNB+NF/1+aW9/HwCFrmtQS/k8Ck9Gnh7
8OJpLzBq0+M2AaRIczyMwQEaEuhHjWyYq3bK2g9wkT5WVrY6W3/06TZ2BMsLEAWZ
8rKcta4TdvW6X72AEgrPdPcoSwoG3uzsy99564fme1XSrWJN6ycUWcF85BOB9xpt
GV3sE0rD20s30FBPLLefjhtMadZPim3bCshenun85wqrPDlnpc7I11HFeNxrAqjo
nvqNt+Qt8Zz6ETXQE8sFG0jtZfnL3JVknk/E0U4s/kKL1uIBKxjd9L9x1GAD5ONu
RNRFJAD3AJN+FRnDuHQQOTpd31uUXCRoaVrrDH7PyYiRWF8E3zBOaOb0g6ivGhEk
pK5EPWnXbCbGa3c5fwey5lYe9olZPcweBnB4mC89jNawFmO+fUKn1hTgYHm2fsmd
qztQE09KjZzdYqN/HhtHQ6b1CFen0D8aMueTASaJSqFmr7kl8gOuEYwYp7is+iuV
B/ZYzK2Onob+cVOGwDEKX+rkJd6PFB0C+vKXYhVQiDnLVOffCbQ1uQKXsFi4GIVr
uOFrsYUQyypXZ9lJ0CB/tmT8869zJPUIpKi4cTcJbHD+0TlEJdhm/LbsVLachCf+
Y9fk8uNG7WvblWbx8JxmWseTmv4XPqY6bU6YVCEGlADoz77Smtf1HLFJAdQDwofe
RryhKNluS8y82FRXz0U4KGzmufnXm3cnPq7NJXYdc1pKUuYZ+a2S8sWi5aydnjTM
IGIK5wCzmpt5kUbBx205rbNAgJ3OfaBqyRkOJalWECvgG21LLBE7J6N7oRCXkwUd
wpag+9S0xNdOVL5RTglxMdbutG4yu2uCBMJEUe9/9IpMu3ZZrnzGLns1NE1B+eiZ
UCAeJIGBPsib47gf0Dh1/M7ExzLt5ESnRknEfrNEnB8ZIU4ejBZoflQSUd/Pj6Lt
zuPmUfixnLBdTwpVETgsuKUImrRTEY4ynboHS0uPfYmFjA/xbAlxfGiSfYuVAI4e
wIRP7eN5R8Zy6uBU/fHwRJmfwTX+YYxoUBOStMiy6GRIcct3bzfRtazxrA8BREoI
XXKn5TiLmUDlzHubtQXjFbcKxZJ+6E1HmbmQyN50x/Iq5X/M1G5k5HijVfuqVEb1
4k/5CRC1C7NgvX5fUYwnGePeKO6hz/Li4p0WmRu5Us62dCXtBigMf2tpYGQ4QBE/
SGs31YcSrCgbkdxNH+6u2u28jekvJhAPXby3UnqZ14HYH2cYIeBENOAYuWQUckOz
xPqIpxwXpalNJ1l10l7Sr5JWbIqOVrIKsZB3skhaLsrGEDg9aO4OsxCSVXnZJKXQ
RjaGS3K9frZcl4rrF+0qKPJ4GladY1YStznk+7wuKgep8jDnqz4r3H4LRsEjd2ox
2qVX+kfWHWrNOVviPkASP4/IA0LyKe+l69MMDnmig0N1HK5pWzLzFNDXnIN8D+6e
38kz0j2tuIST68eRD1zEUZQ4TwjcQq5C82ZhYALo211IVw/mFZilL0yV+wPPXzzb
MkhZpc2S7d/mX1zK6YUlN7L2iSFQbmcspmU9bXR6IBu79R9xRcppXANK7fEL7cwm
80IQWf57MU6o1IvobVA3AppaYUw87Mq1dMigUfWfR4tX3dlwYemi3gtn3a28SmED
6NQ9LFK2qRoDTnRr/5u6zMA1TK5Nn/dT+qj/rDa4D995cP0KS+4yGklDRbtLJ0sZ
JSdjFd+7fzIKIngDVwZZfn+GxMpHmzGhOqTHpzEgPtBfAubazYpZQLgTcrNNr5ol
gYv4O+Wnqxz0O/IwT7YJMu5RRxBTakX91CyXaCc/hDLpHGzDo3KsvuKb3IU6DfXn
gMDdEd1WRXzyLcLJxyk1XYyv9lAQGAO+eXBGBcONxLtJ9R6lB+F7f3SNbSXMgMU6
TPtbo1CHDI+i5rFcqbvV8ZE74nboHdKJY54pxzSrizZ5MF2Q3yT9eTJhQ9qPDxrU
/WzNRmdidADrjmMQU6pcHyQTxdF0H3uzmAkj9pkw0Nfp4S93y3httNcSK1uX3Hcl
EX24LnBtMRQHF/eBHCdieDsqhV/7hGfJ1ru1plLAQu4Zd3IC8OOyMR+ehzMeiKHp
XhCufUBvO8dFG07Zwn+QbLh7NFxbc3n7KIfbSSw001yfQae0pqbPVHI/ttBooCbc
LoQgHle7ANM6GW+0isdjhGvjVIlTCK4VgT1Lp+Ri78g1Uc77xjrXcs6R4jpAgrFw
t75OL0GnaGpf30ZUt7vggYa0tf6rojcqZsEXbX6xsWOHCdBHlDCIcuu6LgnApLFF
mc/DquiszyjaYILyjuDOIvEW/7qQJhJn9d9DvbysyvrE8UsDK8lE5voaobg8p4FW
E980Kskh+FM/xuU4Day7uhVoOhQK7DZTz/MUcMNJuBXquRu3UMSWmSDhd68MO7Lr
qfPWSUCAuUSQbd5M9txEiH5WZ8Q5q+fuzgUFnZuu9h8ihKEs5EVGRu779w2zGnaN
TkB1VS4/1C3cDAwuZyMiyVP2aA8dvKu01fN5Q3E0QvlaUwZg5YBm5lgiySx2yyUl
0WyJzukvC8VpKc9VV3omZnYmv0l/uKx6J2nUHH1U4JlyPkWGtYW2Xvob4VOJ6V29
6r6YLSeP1gitMB7ZPFwcyRes8qNEZhUuT5KDBp0aQr+V+5hSwLuk9yWBsGR20C7o
7Mt0E33gpdRH/wh3ao0wEeYbBmE3lDwOQMu1yyNZTYA9wDcroHUfIZfeHWV3TO6o
C/9O+eNFN/7TgV9LCD1eNkZ4ezm9V9XbRbZ40Hn4aNMka3aJAW5rLVSPCVXqq6VQ
a9b/PbG2C+G+VmNFK5GrGl7YwH5avuSwJk1hROxFsrggQV92956Sr4ABmrjomO7Z
WZTUmR0ZB0ZFpYiVbFAdPfZQAb6qhfJYCUm61vzCb3VtPh/c3djWI8vQFiRikDLO
H6SvjnUMFKV/iJhI/fXEJVpT/oo9Fz2ZQTpGwVb7HZyCyzCotjz4qsCZ2A8vCOkO
FCrpiMCJpTH/afMbZRlpuPzM5zTomBhGreHw9M5RBpWfSbQkL3k+xKJApeZyBdX3
2rWPlBjAEi7aKiB8w+AZDstkR/GKxOq5vDzX73wiuQaq6yQ9/34KvRcvAz4IC9oO
Smmwrzmx6S64ay0mvbGTO39z36ss6FaaNB6dnMPB2aoYZxFCL3Bm7BpAv8pcVGNF
r7UcU+7VNRlNJJM7dAFhp4XWBnr+jeTk+JH488loZGEF3q20ASMcoOpdI1TU3Gf1
AREUGbAJpv8h0aF687fK1w/8w2sAz9ZRn1RJSaue1dAk1miRkFA1n5hByxwkuSfq
t7BxsGzXuQ59tx44kqPX1/Jtj4hIP9fZAJx6qvWQ0OFjVsh2eK/h7lY2W/nUHX20
ICCPkZ/XZgzAQMsH/excWOc672UcfPTJxB+Kfb4iJVeHcR7JT1fMpdAZyzhBs9iT
1M3gPPcP/ng92gTqCMNkEKkOjjuSgRotYi8h5EkYYgvvSPzbRJbnF7TMhgr/1L3S
oce88Q/lqb4o2HVoYLqzoiJ5eOJyZ14lQ8zfS383y0SCO1bhpmFzjYUFgh0lHQhu
DEpvqO5uoWmirjUmDEwsbd6G2NkpDQZ5T6AIuv5Za0K0rB9/a8rlOFfiWzYBMFEu
dmhowpitP7Y7yPJPgmF9aofhzjPkFzOpWyjllPFcXCUL4XfAyPbueoVpwZvitoWn
XQvuRYW56m2MTYfPuVuUXGwgYXQu2NZPIJ9Qy0yNI8d7w3xV+jqT+9d+eHDajj8q
K7jG1SP1ARF5Vbkbk0UgWx9MhAGHqNEvkdo2RdjcdFSi31Z4oGEZVjdOitwkUZUH
wawuBDA0cB8I2xi+51wy+Mq06Ox5hnXaCKAVby5Q4JiB+6KQSvunC1LX7aA03HmL
3msD34yCriMHWlROLKZcfYPFOMwMP59YJnDhY2jYQNaleXmDQN18QcvcCNEFS4JK
BVGajOH3GdEx41eZmsqiWf+sIrorVmrLfspxDDvDqDipOIn9YoxG81SVZ4ZELmnI
tf0I1ysav/4jpkggPGhEyl8Q5EYtPpR3vesp5ciqjrS6YrA6DX3PlJRB/x2lO+iS
WL29JJrUmUJt7UG4aHjQEeddGiuJbyyKTG4++nCJ4j0IA6taJ1luDVKSprgLh8u6
altfjq4H49iOjt5qOVz/4CgM7ndhBXkjetHIre0QJLB9JHYeGuYtXnqX8F3Cn73N
z5CyJ6KP1UG1ai7OEmhHFv1CcJXH3+1Z57i9ZF0mqNUPGu7ocM9CIcPx7LdJD6It
8mcFMr3oUgAo59cM+oHCrWqbgin0BNtPdtO4G+RG4ph3eliD98zVtp3MbcaVCSZy
FoEXfDGMXvt7HP6V5Xg4IUUd/hrtHQ+Wwv2PR21MRE0HAUz4b4pykPyM3XXIarpN
KokR6rUoEMHrjTa/7ukJ65KA0A0eGr54hksrfULc3CtRO2kEdDSSHkn9shcRGtcc
cUkrjE/Qf0JJsH1ECwR4TQnPjugophjswhiI7yreQHHNOXxm2bEdZRFVaWvlUK6u
Qa9YgNQ+YszfAFrP7F7jN9226cBzQYpYp/8D099QhbxDcrgLPrc0V47q0jcduIKL
70tumlMH3ce5T9yxveM2ENvw6f9+3OxyYE5NOt6x4Yk6Z+dsAlvnbAMrbKky8nET
wJrKwOgEoq9p13jcauy1mox2GnEDUdRGJJc/lgvjMlNrY5LHURb3doxbgc7FmhIZ
mG/wkV1uo6CSuRXZLYDsIRVpdztuHLdA4OEs3r2xAsm2CUx7QUy2VbOWPTz4yL7N
7ExaBHPu6aFEcNDYpzoZTAxEAtscTrQIVPvf3b9K9be3Jt+FazrrzfGB/1fFdbbL
Ve/Qv5bWEK3CwFnFXRe04STc5Lo5pc2wM+sXPbc8Qy6xHcgCLvkjzSN7BGmebmzA
vcfrXTBIeN3u7qcC0Di+Fk3zq9qL5VIr9SMcdaWPDnNlcjvgNOTsRKpE0S0S7YA1
CrsEB52ILwI+ZKtRHj6s6h9hX1u2DSFqlFxW7lPXsQCfLtLN4cGI8ufVmqE8uYb2
GpGMH1E2Yh2EyF/mRbwMBd0AtGAcgWiRoNd6YaRA7QW22MG2GgrsbgVWkBDjKQtn
Td6jrBq7yk8SoPYGkJJ2LQFWXhM7A4P18A87maCAXPjTlzEdIBpHXhuXrn1H4Wod
kJbRwCMobLG7PVWuuYKziK/gocsdblGnrMR/230Iljh+K43tv2vQBylgnyWim+CA
t3lLcYc8wDIIyu8Be2+hzUw2q/q4S08VlSGd2Jrup69V701HF6IjLGMMYNQIE5bZ
N697IT3SHV3jhP3f46mCeTxKv0kDAytzHN6fhXtQ3zb7Uf/8erHpZhVtYJq121xq
8o5kpW+pxesR/nFTiLE8WwQ/g1EzxUcOmV8iOgpBWr4DGxVxS+NYMmjnBb2AC2Rb
1e4e3v0rp4CA8miF9LDbhx3G3zo0LWilFn7DYC3mOm/FUsXVBKyGopobnqSndQm+
t6iG+8oBMhNl3f0Qs3r5NwbNIznvwDKFRjTMNY/4ArthoSHgC+7chLwS/3gB121t
PdjRLjia/rIWx4z0W0KEBf8Ot2QFp5m4DTx6tBYvkNfEaJ/olRbkmktKSSz6nBRS
WwThFwj0hX6eAFtkDcJnv+PS71o/TZrAY/5JVI28xNssKgOrb5ERj3iWCEV3ZeHj
g77TH2P8XBqQq2xpwAnQic6x+8hiuYAY7d/uk/kSupSKn2CsHyba4L+7ENd9YwcL
Z/4LFD5bxEaOWRVETn5mIoZAWdgnEUMqRRyS5fxfZWVNCzr7hyIRQgAYmwyCpn5O
onVjer1gvTZ2+U5yvLmxiWPJ0nhuaHy3gmCxXsdDTYKhf4Ouslfu5Cxw4C0bu72e
efbBA6fMQpLfODgoKz2hrTdq1r0MY5dO8E2ol2tB5Np1vOGlcLjZFMIsNBW2bDGS
pmdl69b/q0unF9taYCsT6jLigoc6JszLXBBVBW9rODwFUYMD1o1Ob3dA8M+GU5PF
9D45uTB8uXXc3UQKkwmxW91zYet5GoRUP2pKpDkQBfvt/5DCtGM1Wcgq6PrHFg1l
49rV/COrrhZzPAZVxEZ1u0f0Y6IsD37Y/xduzSyRuPMlAbiFq0EFFf6UXkEfgZOT
5nRXBWZ5NXM7PkzpCCkGB0kSu4rIfrfB9JTO/R023iW3WxZ4ZX8FljFut0p5FH2I
SvI+sDR0Wimp0wDkWusoNL4YfPjHs5+5z8Scd4cWThHLLx3cQdRVXC7GkjqrbsAz
A5VcTessxC9VHyfmAnT9HuAhzUHwxpcn5tjW7x1sMWtMQhrhyDynNeo+cuzeeSPB
PnBkMHJ2mIskCS1tSmX26qCVntUrkeCnV0b1HtGyjtaF99mKdz+Gw8GTZjVYjeFe
PUE7APdsEFZlohaExiET/ICw7czsHbKAMclidYnd0QCvog+86x1Zw309iqb+OXXc
c5MlsPb/Lp+E+xsNKEMD728po7vh/t7db+vxkvb0f+cpfRQyAVe3dfqbVcLiJz6M
j8KQvzb9TyJ53W1ry3qIFaLmd6k0bSfRDO6mKpPbwvRxY2EW/JbJWd6DjsGbRp6s
oKWKrBL1jNMvYj1rVhW2E/59IGjTcXIQtCgPMAqKh9ut/YQLxgChXq0b+qTXNdPz
U6PEAMJ8ozXi04qrUn7qRzT1lBbu6szLuQFhI7tet53ePYqA3vgVTb1guDcNoKUv
p9B/ali1NBjeEiX2cD3qcNIUqKNkt1aLL3Kbk1rqzQEa5KsHmPktbIqgFx1TtsMq
kveWK/z1mV5kaBZAIQRHBK+npiL1b9bNf+DmaKZ6uQXT9mRuY4iPfwvqhaUWu94+
eK+cXz55hQstVuistQvRZnzsRYsf4zvsAYPjx738FuWOeilLV2pd//jkVo9azhmt
NWavHEaO2WH4DGOTX6nb6J3Wlva/vcg3Wfum05+zVuPVrtIheGaKZLGyDwuCzsjF
YWNn7ChJCvrTOv6MCh7b3DjJowOJzFQkG/Sh1O7YaXAkYRuR0xgV6vFQk4KzHDNA
+6DINdrjzFEPkKPpQGgNjY2kXJyxxbHLwuQnCpcLM0TEYMzw3ujGvVFZJH8lT7Oe
tyl48ZReVwATMwb3QMK3WpM19nc1zYxOvBvIFWCe8vQc2E3a5/wz+YrVgWmpPZOe
R4BfDAADokkq4mk0xMY0TSWpziQldsZhksIc/q6iD1tm3SQO6J2Yevcod/Cx5tl0
eClNdURO3YKURcuPzj5WQ5lAiu74TYsNLesLeX1eAfMJOxEhOY+KO34/M9n3zx5J
G7T9c9kTql0S8aNEc9UHg2CNyD8lQsHgYqmvb7udzuIOcgFWekCOK6cgX/h53imi
6JxXddykntr2GcdQSGmCNG9EygdgZxgfSXbeKGbx8FkC9Op9NHMlykprNnn6iRKw
BauXdzhKSgeqmgSMN5Jneb947VkIllDl5lVK8qxjv5Ty7NrEs41Q8skWfMaFovWd
BQCl68WnrzD27IzVhOkz8KqdiFfnmK034ZjbnivV3crKEkcHDaZ6p4isn234Q1mR
dFlMF+EQvcIErwiasNTNTl4PQP+/jUED+R6zgCyGe9NmKPEda2E5IzcgtM+3HBWu
DfDsfYa2HL9q87/u6BhLM3AhFPp4tu+8Fyb98y6luaHJWNI2BPlJNZDRGJRppryX
u5HnbmCpicpj5QAbguZVwRDJvcuNMph3PuKghdSp0J1bydZCmX8B7XnynoQLOnF0
8pRF0ShWqwy+4dkvslxODAPVdxOE/ChGKKvHtz6nogKGiJmMyzH2FE3pFvt1zfST
U+ID3Lb2wBVKfLlhZxfzsLqBOwOH/huODW5fZbIeEsJ5KCuOxb7gfxCsvk3d3Wau
l+OQccbQWZfnZE8f5isbL8bqAGCSzYv1IJ2f+Vj+ROJKV2AcCqqQW5ublKslbCWy
IiWTB3S/zkJec2xPrEC6HsIX/EQkIUxrRuU/0R02ObXatViNdOLSUBKjBxU8awLs
VATslqfjws20GS36G2rjcMf1vIoax2/ZElhiTpmFugsmgua22KHY3H/+4ulaaI14
WlxM0LK1s6vjHzHfZFuaK/mtbFbjlf4s+MzSfYo0+jbFg/vKBVR0XdH6ze6/EVOP
TaN9SRuXywfpdw+Ud4LvFBVVj77bTz7gvwnm8idxTQqb8Mj7nXGLMbs5ez0Qh6lc
uJMm7RrmLsJdtkZCsZ9cWMj46dersCVbbANMgs5x85PFfnE8Imd/iYT0uqWJIql3
O9F3Zo1TbvCtxBWiPKn9+vZio+/pvFkIUrbBTi09hqtfhxIb95Qm2IRvDVSS0Wm2
arU/G4nIR/6seR/AIeB1KHhC72wiX8GSvzxe38MYBuqNkZVWP+5725UXevNVTI1c
CBy+lCGkdnmq6mIdSaYGykaH/W0q3Z9925W62YTrZtoDw4L+7IyWqlmqY22xGgeX
IaVobVFNvqFpLjO1kFWE5HeAXu8m9BRejoyvOgE3hIwAt9hCsBnl7y+66InroWiU
0WNqGMUWaLylt3Si9zwNBLM6Tfc03/bpuKgSG1Pd+gbRKMdW1IqdYsy3iXZWlo3w
RfDbT3A7z7IbIY1k+lZ9+Jx0vFUMB6KBBe933BMd8eezYQGujczI6jucF6IoR3JK
lu2FRxJDEQQAqh8Fhcb7jtcpvVhg74aZrkOha3NOHwRojyne6vPeq5ks6fftB0QH
KeHgTxbHtij+LLCYvYF0B211j3DE9PVEvWWErdZe0TIihnEIRqeKQW5Tew+QfNSU
/pYxnvFLKBcahfMy0RzTfy8lXRWyyV0coRpuI0jYh+3uUx5Ad3E/mmwaXlQ6iEVQ
OcqnxwZtTBvVqEfCoL4fC/t9zdD562/gnFIkCC/7Km4DKlmEEQXmVxInQHRyHGiE
GosNOMJq8bh7nceSfNxJ/sBoq7cQiQ8hoX7qCPHuxLtlW6NHXZ18iUjS1imL73Xc
KotQSHH88YCuDZv3cBCrmasv0TTUc9DhaP+yy2qrjwM8N/gJB5AU6P/Tgn03vdPf
nvrkjL9/0nbNVdxd0+i65v98yIrYnn+3FCEsAdM5ZsHccHt+HzKDarsoG1glNjHx
DqU0wV4I/1tOgcALtyc/biuocnDAxbOp7yfQQbrrEzDGPKiP1rftmEQRgZjZjJAS
VAqfbuakMB+AnxIQwvfx3/SqvUnmOc9auvIoJgnPO+1UgFdvhKStWRTFuuATZp5D
bqLe/Kz3A4UXxHEvYJYsuEoACIGxoWjLKmMA9nokDXCwP2rVLpuXzoGU+aTHvh5F
ZU7eUMToC3k7+ygtIxMlbEo5vCHRZIXId6a1NkHEPH45BuyuKYBxDhhXp4cYibLg
N4nkVU49brQqnPG6DvEgfFuk6jn3gfSNk2RP+w+lW9w1vBuPU3BDKqGeWrwOgotB
knRETw714rxSdA3LId3N3ZwRehkLRyy2958j+qK4lt3H0YU6NA19sHbdMyxbLTHz
S53+41iWySxribemgc6hhu1B1HS81bvyUQjebCoQtuhmwAUsUxefKJxotnPk6gZk
rN+JUw6XHdoj2VkYP8t6+vvE2Ai18ADIOVf1bxG4t22kz2bwNUEsILgxkFX8ba8B
0J84hQz8veu3KFgVauPxtGwUdf8SyF6/WlfJ7xomRnCcZfvkJaip3LpQ8CudfK+u
B33rCZlDqS952oVbXCg3EZi4IrDWlbJN3s/KfbzYccKdmzFKm4XBfp9YZHHPH4WH
xcFrgrz/nLK/3aIxzv+HrcZf/TXWq1PPOHdFp5AuUZLMcbCBNxeeTdGv15Y0r+QB
YvPohEiVr3XvH7br2gfezEqS1J1tXxHG8QOO5d+cUYiGj79OVIDRjubFndHDBpzm
AZsPWuO0xWlBv2HEKYSWTw4I6p3brdGo22rcDlr4OrXGnXEy+aZDyNrxYC1mKRyP
Hj/oRB02SewY3s46pabZFkCwv9E+e+NsORkRG3dnwm6zZ0ZLkUxHHTyz2uAk4XgI
6cXYsbib7MnOof82NSVKVWLyPNxZZyEhLH46i49wAeMWFI3vsvz40Si1st6BlzZX
vggs14+MDIcAxmTD1op9BQ6b3zVG0e6mGyogBaGzNzZTMdTg66O+80NMj1WlaPFs
J36g4gpg8b2izzMvhsd+SD3DSkKo0Ms4BH4ocbJVa9D8FCs+iX8mSpEbxZBJfXss
xi4ZhIJX35jn03gYtGxUOzGfMgkG3YhWcbMD6zBy04g2Kf1W6fm7RlhBwC3AKQTt
ss3QJq0/Xxr3fGbJCt5b3arklvieATP7WsqHoWhBxNEIqNjkOr4YA2Ge6siW1q13
PQzmRefDNJoBJJf5gj4y0BBb7Dc9EOZiimkPG2r/sEvADnxw3cBTI31OKQ7Jekny
NNrpSFQ+dMWMupS94PkBkQcpsMrxq2j4d3lE0jWoBkI/RWocimns5K3+tY5Xrhiu
f3nFsf7US7yuHR8Kl0JFG4/GcJgmoJnqpWe4mvMchfM9nrv5NWP+wKb+tqY+lIVF
jEr8jhmu1nVpwh4YmUWIJTKhqpjUMwyQptfMAVHEVxMb2LzuhWto5tWzLFvIiWWp
4qEq/4mbsD2a81shPvUYmPRzm8fCTZnfizwjpZpXPLJC6oiv+Pjj0oT53KoJQeHX
1mOE4+KP8b4rfuDAUBwlYGT9Esz2Jyk5wDhHI1ZAIEuJmC5oYEF3HZe5nu6peLh6
9jPE5/iCdPcsbYGxS3On9z82kKeE5tUjdeH99VeqHLI41ROffx0HUKFCc0C/6sv0
//bw6/t68c17ZME0+ZrOgtO+Hu1JBER8LFDb0BCHXb/cSjZ0f7G3zCE176sbU0IH
T6Y5y1x385JDg/iTAfdhFN8le3+6H73hlYvPpqGOm/t0bZWl6mw6ymrQT4A6+uAy
pZscZRy593dhLtsrPhgvBaIFGf4vg7KGuBy88utokYhdJAyAZHX8msRhOoXRKIVb
fhidtVPAjyaBiB28Atfyxarxd2kik8cOjtzz2rV+CNJgQ3Tn2bY6fTP3dv0eXjN7
3R3bo10aR3I4cWk5RR6Pkaa0Jg42V3Kewsdy3kY+thOvP54MuGIKx8z795mBfLgI
51TwUKnJfg8u6VmE0WOpGckii7Gfg5YPs/cND2ZC3wqT9wPNtG9xMec16FsWVZdw
qnodolARmwwViD18XvVfLOi90PzXJenzgZwidMaIxk/5yi1vzuHVfoVlaLIHZItW
zYunxN170HgG6i7B/LTnvVZke+JoAUWCjfUOR5e0kcMEFLPUP8gdv+E2PSJdSXn0
FntNEWZEirrwpVAyjIXFGP3HwiVJ/dm/yB2mWYD3qRsnv2bc+Lf9LX0zehGlqeGr
xUGv5qAiGikeLeomw4DtVNPmmqrHP8lFFQHh2G0tkwti0TvEmH9R6YmOY9vvEGyH
v6IK/aZoTXtaurxieYrnq4ymSVrXBN2kVeIhtqnc832QuyPJdY7CGoyWO7PMJ5SY
JYLBmgQ7U08ue9VbMNocORLS61Qu5NWkWmuSLzBWfjpNt9sEKDSVST8il/XJTOYn
lkyY99xqmPCw8d++/3dKF+AEz0ZjLhQUE1nGl51l+3jtCGh0VtRfLXeCUNvLKdeb
mFQ8lnjbCFP5szLpc0WxQEW9FSvcAq5OhWhjz2a4uPiByAeKudS9Gda/EiHQstZ+
qMJnWZdxa0fyAd1IUF9zXumN5/g8FLXmk/KTJ1x/m4BoAc41TKVEgFC0DwpC6ugV
JIIhoqFMQbFd+YOV6xCggfRjd4DbZWPlTl7Mh71D0Mpj4wmrEsLCBNdmtUdrNoFo
RpaI9Fepxr3SjyPsEMSAPyX1oAXMyTUnTzEBxVCh3eT4OCKZP3fy7Obti/v5oZst
n96yUsWtnlZi8XwDa+DJp6xmKR4a6qf7OpK37uJWWPDavoXOOdWsPiefprg+Ee4j
jcIYN499Rh+3QB2JTqYbliJHXg0X5UZmHam/2eYgRep+DPmSYm84gRHba484mjFZ
BSlHdKxPoskwr5OgweCRppy3JadLuUmz8qR8ukMsqe3zeM7FcCO5WpQELZdKGLB5
Vw5zVo/ulFrze4giuxAVNeCgKLAGXZz8J7+cErFbVesJjalQeY5aeHRFW0jRdiZB
d8LpRS9KP+jskvrPLXv99FaZ9x8bgWKO7x9oHiNQPTkXK+XW9AnfJJwS5LRwxiDc
31M0ZLPjJbuL7uSd85zxo30BfxTYeKWCl7k3L5UwDyPMSgNFSrlNl+k14bhxcoxn
xulsWW3Lz1Or7dvbbV51WIJdeTp5Kh1Apkx1Pug5Td5Wubkf77bCrBygLasynfv6
niqUm+ah2WxIW5c1ENlRfKVwzz8ArlE4bvukpa9mQmpSjrFZhx6WJ5wjL9VE3pl5
Ufv29RNR921pKBi0M419VWfIXQBkUvxY9Tjejq5iR1hBqUeSODFIxPAy6EN2g/fe
+Q1/ivGtuavJhD/0AyYtPyH0pVhfNgSpFFQhPsMvvlyQWIYssm1wCCq6+FnPE+0N
R7SWjDQFejaU/2Im4B5lBMotf3a5odWwgFG3J0bPxdoY9wgMVCohbugPtax1Blu2
XSqs3vPt1ibYneCitCOepOXimyeMIK8YsTi86eJDLqJ+2wQe7gBAf28xdgPVPdOv
d8d/2Qr1tzvbjC5/15gaMsdv6NR8wShFCiV15+6UlmHrfPhv1CYqXz2GRByb+hnF
msPz7wwitYG6/cfQ/lwikAjXbgLUl+Z3g0j4cIcMDqcj2qulmwEV89hpL6XTB03+
XO/MHqu12z8yQqZPRYy1XnldXQYNViNmWxRUHEb7rI6MNfBgth7bIPhXeFblCg9c
T0t0akVXCAWWd/1MTYpiAoxi9MmRpVm56VlIAmZbLAn3sQhNExJgmjc2dqpG5iaO
heIpTt86yQw8SSYDGjGVVUxWd6IgiLFC0PXdSvXVYipt4MZ0AKXS+XFflzMI0UDM
26nNnfEXWPT/6rNUvagFOwwuzLOSjG1sHYPAtquFVn+aEH+H8YZ/SlEdOxCVHcck
ApHoVPkLctLfmZYI3y6Ar69do0spVavK3HtLR1EmSt61agGkdzRiOB/UlsGXpev8
q2fdpEkEsr7+oQp4yV6XHLL+6J+bPTb37QHaNuJ/J7mItfC1aG/jlPYYrITAi8cA
AfBFJjtmWrf6jYW129bMq5AZZA2BBrfKrYcLcohico/EFDzmYJ/CVcWfZi2mgUu8
8d4NlwdMYqv7L22BWjf6+lRB4QZjKdBzt9+0FOxZr+Xl5MoBMsfYbEvyWEH5vGJw
mZO890dV1TK4BhFj+nZODSTObHtKc5MTH7gPGFL3uQ9lw1A2JuKsXfQJo14ckoQe
oxtOg39GNuGh5DQq2fSi/MoamkvnoeKcDDjzO9pNK/75WW3Bl3gbfsLZPmJh7Fc4
OOA1UKVWn/zjqbFQl9Cjp0ZuS45SDcxnZJLTkUdYmqUVgXjtEe7OOZ10vkDrcqZc
NMOfK/J5s31uJtKGmaWHXmc4y1CJnbrWEAN98p/x1t0EJZBsM5zb3pHsIX5Kp8Fq
xMPtapbRDzVf7Tx8pgIXW2sN+WM05BiI/fY6W5IqZhQgofU1EemTMCJj0P+3WO7K
+KS58/3DFcH6yklFcXzeQM8Cb8P8UVL7dm9/++PBULhLlRxCks2YYzycIH0UpOfT
uXy8LDwX+DAr1TKZpxWCOwqDJTbWMmPZFafaRz+0/krc9ZXplz4AsauSDHH0M0GL
1BF3cBS1aCqhrizGOUVnF6ps3Hum8giK9PexTPtTXMy9ywehtApBp8B2EtZDLjGm
jkXtrtTjQ1PikGVNC4OwdtUamwjPDakoO+WnMGj4qmiHq4Dj9TrGO15j/8nBJkpp
eM0yldVztuFvAKmnyzmlaOpQMr8DJ4WjfUN+812HKcCdMIt8WSPxYpbuF8KWE+Lj
Ti+C88An+BV67NT1nktQiLWiIyBfVYnCVfZ+SYZ15uMhq6o1omO4QVsB4XrGIQYd
KQ70fw3ZBrjBy/X3D09UG+1LUC2mahDZdpGwqTqTQMmsn4uaDjLhlJQJXopeG1hX
a1DZgWxWBeCkWNRd60ecHG9tuyxubdvLgRD6iasAbqZvjQc3D93kTPEoGoiTYaXN
URI2dILsGUGHZgn5nr1GqQgOpvTPZ63s8aK1W4fspjlXIc2UlsKf/cOoIZk3wQcc
vkHwt2Et4LRH6D7mScMakvERfQQ3sAy2JVXbm1ldOSSP7UBE/DdW+LUKQq2PYOCv
Fv4FdotGhuHkz++twfHak7XFH9aWbHjZUh0bReh4WLdxOGI/xRQsvjg2S0m8f5cU
3tdWpyQMZJJj2r+tvtMdnB9Eltk5OtP5awedXkreupmmjbWZhWHcUXiyrIZVaRlh
cpUuClpO8d5NzRbKcskQLb3/QCyAYzodSQepJD7Tkn6FMwJe8KZUwW+IMhg7QCr2
ANDTUfG1lv50ZptvOanIkuWi9R4w94uZTNV4r36H+ymxRHVxMcguU5Guw4DZZHF2
4UpOS7fuad8EgsMHdA72E37QtYSmgoVWYOcqdZjme5lCYsMFEYvwtJlGHL1SMSSZ
vgw69k+d3Z+Q/uW04av0FSnZrYKDbCVmuBLug1apXeP+tGDfNhjrj+cVk9ekD9wL
KBpHJjBb+UslWr+pSTWx3C7CdSiunXGN0vD3RfcGFLtvdICG6TgWmay02HKE3NkV
MjgRrZnUuqVmV8EgoaGYL5Ry2X1Onr2RdcdHW4dhdPJAthWQUf6iARxWnQi5tRyR
fohzrFaSS242FT3XqxfNl7NMBX/oFiGuZMS4vV047PnFPldDcdidwdvaLaTijEdi
EFPLz0Q9Mg5n7WtEmfnzMfuYMypTcQxIUedST1yprgjIbVZ4vyz84BcHVceYjDgm
GZCb5Xmt01P5BWEKv08KOn+/BURIJVmr5ZoxxCpb5Qlc+MCKQcXS2M/VaJL//bml
0B/z7wWqCwEukxqIS2aoRPr3CFYj3vTJLpy7ibXfl4LSozSWTIuW3h9NOASr9SR4
uILBYIJL4oQIdt1Jt/U/h5dg0H2ghwP0gM6XX+EY5TA9mmQ0AKfMWkGhzv6FAbMJ
HL/zhLtTEcpqzMKHVO10nv+IOUGF1V4BvzcAY4UJiCS7LNefMcjPcOxsClQ5Fb5M
2cqKPIqsXamBS8N9b8XU1/hifI1NDeqIS2w3BPUqg8Xd5Oy/VUCZ63rPGesXfN8p
hFRpiFgawCspQ/Jo1/NWOSbIZzMJbHN/ft70zB7mmq3ut1u0W5FQKj9zlwu5bgTN
7AV9DAOyKhfxnOcTQLPhjufGgqIzbgObMczsXKdzeQ+25NxKDzSY3rOEaiP6UR+9
TSqvNMbNAeFs/THB/eo8nzjpQc2+Yg+AxpMgOnSqnr0g2ymwr05G81MLdEsY1meX
1DCol+UyvdbatMyRJ42l0GquVlHccR3ZPUllqGOTbMFMSRk8ayVqknB75kfHjQu5
/Bm7q1LszTIxgnTV3qHr7dj0NPDdIRzXyhYLvSDNisWdnV9EFBVpD8Pqt9PvhwWc
38i9npRslI1EOMJSg+tJQbXKaD1zIcp1oMZvJuUWyvhCDRKaqczNJ2RCOjp0T1Jb
+BXPT18rwZ8jsG0kSFAX/AWCPsAi5uKJBwtOJm4D3ixaGiqjmiESPscA9OvSC+ar
5CcS77Mdx3RjHh3nMYzTDA7kFm8zySjTZb9GXVvlP0NA485Vo9e4V1qB7x43iHC9
98YHOM4a65hIr6eMZi3POdsQ/TPZRTZ+K4PLoEV5h+aezohRAtfvxZvdEuJAQhat
jo34P36JCSxwgMujZU88gPc0xRPdMvoj+Ygwz+y7umipb3wmffbKd/wa7mNw4Qr5
VqaE41ba6vq3ipedZbqaShxQDiwbvDP7PzzIPX1ADKgD3sNFyAABEiRxcUN0HOdP
CqXMOL4LtfNCJsahurqG1A6uIXz/RZwIzaWGHvvN8K9WKHxwUUMUc4oLpd5WWcDd
cmAHW7EX3kGwtDuFYRtYn5/wip5XJ+opjnbW4MYEo71o4yWVHoaiB4V7nxq/h1yq
P7MHIQGFZZs7aEWv52LxxrVjj6/Hyn5pcJaFqz8Q/D4XI69zQdWS56RyarIo/9Z2
3jS5rA+jOktlaa0lkT30KJA2Et9Ko8IjoanyQfPnYfKkBvkl2TPfTz8Nk3HbM0ro
UH9hOe7wsVjnqfZDjS91K96Q00kxNU1Q5MAsEGEosPg76GkQZo6JLfVuGjZPBIs5
Q6VeT55WqdCym0pFwsqoq4CzRzB1WOZHu4v/9tFGDHNGQdhQmeIagYvdKk2dRge/
gKTH6S4hHIQHR5nh1Pi15PEZz0IwFgA9a8Djs2Xh/6nVspZGvckGYNl9FRnEQ/gJ
VHMI8ktdrmG3oSKqvOShLR9KA4iE92yzFfg2wHNoU3KIo85VewFkrN9kG3xkTeXa
9wKOH+AJi6dQ8L4/+/IpYyE6TAuCpYPBxY0dU580SSHXY04cqldw31hnNJIdijme
oErKESvm/hEUPpVfmSprOOx3EU/NWV8aXbkNzPS4inHXTJdtruRHLeJy+z9uTP5z
nPbX+C4mVbM+7mcKd0z5R0L/ZHSlMevGXO19itHAdX/ZmqyizV1EvN1PCxZwgUZn
TAGSnLn08yqcG9uA82ooFXFri1NaWoWpnqPkp6J0MgwkLDcP49228UWsjTmsZ0fl
/wfb+2FOLJhHnQbPMzNBvFQrARPoVZyKy9o72WvKTkbsoARykJAcM4fdu3YpWLjX
oEgP8EwANy9+WR4c1AVNXMZwsLH+1CXxhGG0kkqxkL9WZ2Om2dzLKvdQOIU0dT0l
InMLX9JDVajEtUCKd/G1I8NA7aTR7mUoBpuBMMtsDNFJYYAiz3jQz3lHmPK0G5Tq
W5YYtAr3a71kiImKnydVdzvaULqZqKZSzKyADmOO/pXuRo9Mtl9yCzjYOet1FdPI
vN+DshqUxpA67RYdsX1kTq2tdLJcKo0NxF11/3MEG7czvaKl2o7dB7jIIdt7ogOa
k0Y+Wm25K8b/ruh7f369AaCnLiLr//BZe2TEphCZkMphrRgiSv3RyV2eHo0rJ//V
MgVsiiTIndoKZ/EfxzIiMEVY3e/RyZ2bNsLmlZ62wC+dPH9y2etq7pmJ1Z1JLyiq
frv0dIXRRX7mUbCGo848WFYUmlniIGe899X/cw33KmguYjK+8gSXE8pFqX1TvfDL
HhbwY0DKm87qA4KeADRNcQBvYENhfE6A4iC7T97OxGxNo88jv1/1E9Qf3otBJJrB
08uqdsb8JzkzreVg+jIjl8FWohtHN7cFu9w7mqhzzQDpffJ19n4r/7CHhp/8ZFna
8fglatIyzsIN0NnTP2nDZDDukCCut0WD0FkRTh5sHV9FqiGAfPh9OMJzIRjj82Rb
+9ne/KLkdVgd4zcOdezWVBD5nQUAb1TAjrUEe1M3NuX/eKTCeGpn6orBgVNWXU85
ZdjZCg6/67MoIZe/QRHDQ6q5fGvRUdc5NBkGFvqblaQGdh+oh0o4Ja/By1LIi6kZ
ADtCy43pWWa8pEfOQLZRpJW/kY6XGwtZ8xX/PRT+KSk6vSOzkS1Cfd1KqPFAosP5
nby7yRc6CmEz12ngV6x7EWRtnfnmRLbu1g3YmbK9tBlDTHn8vog3TUhpoiT0GO6G
Bkl2oei+Z3vgcD+QTUmmf2ZV0tmFgNPU3zcd9mg9GGrc0+gQuP42ACNP8GLoc1Tx
mhxzVTNquf1R765ztU19mV62VLc+5QYmbuQG+b+rr6ncRFa20tcBHiVKMSZWZhKl
tqszRmUOd0Nd5tRquq0tGamgQME1Qg3v03LceTnhYYKi+bAUVdzAo4Rl/zhB/evR
DSBzxkbCXoJR8r99fKHGJmr6+XwA3cRp7riJpbe2lGqhLV978mmOyjRgWVzWfoBl
XVH6pMwcHJ89BA9o1Ar9yKUwYFu0tC/IN1MAS9dfIQGX9XB0n7KrSoisgZHR8QOu
2kwTOij2upkausdQ9j53hbyNjF/jkAkvO14kgT+R9DIr8V/gspmkfDTe/AL1Pnev
57D20cUKiIjwrAoOGbNoubiR23xrX78s/Yi7kx+TNrBo57KC3BiMHNn0LXM5GRCt
+ApMfPOfB2s8ML5QdPy5V2dqpLe2MAKIIRsKpYTNZviUdv7h/pUvFkVlqT3o5vTS
6hQ+UeITCY3fquxSgLCK9xtNqZKXk7WvtsVFsyy3umw42V+uw9wJFCviGmQjnM48
qsuOZQ1QfC52hPE73Y7JGnZ5+lFdzdesTcHeWudFeoo/QqRtqXlQnIKT5kEABFxm
7o+AS+DJjh4rjiNef9nrkcZgOwbKwH973aI2G2s5GP+ucEA0RrJP50PHRX+EUFQy
KuY88YlyHuxrSa1WS69TpFQB2EegDJLMvP941vQ245GIIVxOjA/O+JIyV7qaYlny
gEwJtjTR6jTvTnKVhBfR1DuOQuOV9evbYuTYyDo7pFL1h3m4nCsutuO4CJFL/Krg
Qes7FuWreL0gWxsHDTUbnvMp8NwUQCPN6IO+BmI2ZucuHku8sdfYpvz3Hzmed78s
KSrD6X+ph5Yc6VSlD9LJm1+dSnobgzxYUPVR4crnn6pQ1VoHdc2vsw3Xscw3Uhz1
yoji6X4S4hs+2XdIdlm7SzGnY8OYh0Hl08SzTEIGP9ng0eX2r1irwsaKaRvc1YgS
nsCtX9F3H9H5v5XnKtsyrve4VITtf7ZGABfAlkCB7fUYR2yazXAXXrprJigWVnHF
wT+Gfb6VHSqNEgu4SCQl1hCn6/BXv/j42b081Fho+lC1pBprbN0uDLXsTj6CWcfE
1YgL1jxPAeG8vmEll3CgBbx2/soJBbivn+OlLKv3VdxRwCQidEnSZ+8H/bH7AHXt
xDTWpSqzU784to9N3cvzKyXLkTv9CTRDvSfOCIRpajmL38Z+lh6SIBPOWN2G+Ej3
WIAIGgPxcRWnPqMhXLlnMjX5CNFWBUlGj7YmMXKDYWJpBPjqp9xloX7plpd2HOr3
ktdRId9vgzxjt5o72dR7G7+vrK3RiRQZX+AXu3B/6UuZuqesBxlnfZxBqT7t7Pfy
wTJ7NvMk1kXZNdj2l5SZl53eOz+lj/aAJWzRRKuAVsLjIrDwPkUhz8otut/8Oqmu
JzV1HfC6OPw8Ym43W/c9hkjdWypIpJu8nDdMW6E1GG6LVaw0SkrB8wWIyhhn5v2L
kJ/dMu81+um1g54PvoxRd/pP3tpUsc1n+9Byu8F1ZiOIvv2yi4LdH62PbKjunW5S
NSvJlyBj9c2DlrqkISDKFqArxFOKWuWevum1rV2Tr/PffYxx2x9oKXV1SSFdEHDh
nofpivT3l95paRodhzqIFwJ6R8Y1wD7VBbuHogkbvwDtHdNqis3hkONqx6NIvIbN
WLeINi7NjLsbTu4ftgln1ldHAi3nRmCNJPe4n+KK6XCuWn+XW8RmwmBFo6U9F1qq
fyzBtn1iIlQg20DUn7SuHoOgWpLlnKzfjX4Ne6cTKpB8Vz27xh+nxmQklufN8zJ4
bYq5JzlL9T3w+srWbDVVtO4vm4ljPJ6PAb8/lkgSYudKNc+hFbN9DnCsOERdTN3i
/I+0PGOih6ofgsvnDAKKaC3+XZ2fXgWvfxZIdKYj4KhDTmGg3trvUJKK+ljvsX9k
ooW/BadHfT8JMMahhAkzc+EJgCKULpuQWoQ9zwiT4J5Kdo4qE5azZFZHyy8sEAjS
G3gF88mKy7a8AkNFT4cyFve/Ywk0QRavHEvZpPE/SektRkPh1sEls9UMDL7OhPPE
5BP2SQx6qBqFNd1KI1zqEVqwJ9aO/gC/lubpA9WiIVPGAoywscIMC//AVBPxUZpR
xijWrj7Tvkqb56A/b14Ax4hU3+GS/wWos0yYTF/Koc9YkioxCMoukELp2tXvgtAQ
ghCbci5k6dIzHI3O0kx7Z/q1wha2FkgBaAL2hlycqkkE9nXrTTsZQwjRi55Y4o4Y
fjOOyAnpu+YOLgPGLAWZaxzBJnQ4bt2m/2lFa583FnTvD6AiQrednOokMMNlROGb
KuYHb1w92LsYX7hWcgChtP3hUOsIGRqsEYIrnCE7jf+BDvWrmd40hpGR6B3nMB3v
UsyLt899gvReehY0JRmpzqsfm4PG5mUhE8uEg+KwDX4rSkHuXj0T755zjpAkNt/8
5islLYEHdeyhFiLuWr2vm+AiGC2e5p6+v2MWRGq0u4Xpbm8iAQeLQzfdgsWN/wFF
HYmM7/27CcEqoys4ayZYk98VcPNHgJgs8uWdGV1jrLYJ1sYthBF77fMiutT9750M
GU0/j97cu7RI2qwKyPG58ZBBlOU9w2ZMVKluMXp6S6RICort723iFMVyCgQuGXVB
fWcHLWyShJtzzxc8BYRiUUc8m7Nqr+meNjn+tr5fpuW5xTrSDnk8BqlPy/cw5mq4
BbdlCYZcfDHXMhp/xJelIg1Bg3qUAb970LW5dgGikbD094dA4X4ql8wbg09BjGfR
sUyiYKJstNwRphRmB5boIcIlu0HNdE0YjdjDiP/MgvvqsG/5SvYrE2SAh3IFrkpi
SSzH6L80utTgxy5AaczqmYXwyEz/gIJSl6ENMKTxxypnexQhZXNA/3qSf+25/Myc
4UCY6qsH6LY8b8TKZVakfjLxcZ1f5oNihxBaleg0YJjaG4GOAgy+nhPCIyeWQVol
qkNIyaUwxaJ5H2kXJmieFmyo+nkiGB4lkB92zcJ6d+fQqCp1lIYedOgEZmXPx06q
Dfow07fbWDppaCmAA3ed0SkBC+JwcXDcR5E3Lv30YwiKsBVXKphCJEAS0MIhc83E
YQOapMbsSlyfh6KaoiBMuERmf8zZ+R0NSEBDoM/aPSY2EVCxCFLDydRDIwipU33N
vLnVjpn8xgahDbHvyrX2wY4Uj+3pVLLqCya4HJhM3BiVs4amjSKsEGAr577kdy6c
Gt/S+DraT5oPt8hO8n9RsllydDM+zL2mZJrOkZI+4NFdrZfIqQGLAfx2gOO8A2gv
M3uEfo6ye/SjZaSW9xX1IxaGN1zJBCVSp2x3cIR5Q+VK/5+OykdyORMOYlL66POT
SsBJ6BX7sygJw5Bmz3B5YWnLPXggv+co2j7HehEFLioGPLn0IDXwoaaufIf1edI+
aoxb0jKq9ps5guRxZNn9htwmZrx3nFJIOr665o4eNdyhapwGek5aqtKjiylVougP
TN5qXabzqRm49FaQV6AvvsPGU7sT0amfulYSbtbklrsAQ34xVN5UjT1Z4fmkF7Za
D5PSiC0qFK9exOwlrDq8Agmt15Hj+TPkkj5pp4OswiR3Ei9mFnNeh93DQ5tAiiey
2ZbVtGLPrzE2W3taXTdpA3bN+4b14EB4ZOwcKFkMzO7YSquWFL+LXc5E507HGbJ3
QzInH3fDYiVIiVwyvkdazHlG5BfNGjMXLD3j0P7gMO0BwgYC1y5LLteFu4kcJ8U1
ddaIR6RQfv1vt2zUO8k1LyhxvghB600r/GTU05MYrexp1mOM8jdGYRye2gV5Wr5x
U/xX03Le97dsHKI+qDpaX7dMORE9C3/J36yHHcHh56DM+wuh+7nBsm7by3o/2q4M
9qmEOPMBYhXoYBtGc5zAw0ckWmJSMLtW3aSJNOJbvTOkhwAmOminwgu7eV/KAR+V
44+Eyp51vigdc1lz9oHSlEy36PBUdlG2EzL7lTTYBX+Kx6zhYAFIIQEqZ8riCXTL
/PTK5HPmY3pSOe2B1knYpunYdAYl6tUAOTsU4FXOYw7zJJihQKcc8/xlugLIG20g
49QIZYvp7c3OeNcBqZmW71lNEi/MVPcNhdu91SERKK71JUpUovvJoMGrPrWpkAXM
/+5YPx80f6fANtjiQMxHGvMBCIhSqVa4bKbPXeJTfzs3f1Pd3uZproUHST86Q+1d
saj47qUBCeQjpuqoGSYAbIgcjvzsB6+72jvdi+zQFRu2XcGnZt6Y889EocasNCb7
vGm3um5zsv32VljUOaSFydXApLLa1MVnUl7Y62qNd1cra6mlWRwRfqb2E13qOYSd
Im3pwCJJ5BExHILKJVJMzOewvqzXcfTWp+ZdTxPAlSXsRhSg7wMRB1/Ban0yiEkT
ACRrzzMB5M5dIIXNwHvtG1rWUFjV0BHLPCP+xoo+FDBwihOdxGy8gx8yCyyDnyKP
X5AdFQ2o8d7wDMrRtrOyUpKK00uxbWonNBM9To3s04OemwxIMBLf1Up1JGTwzEtq
6cXJOOjvD5pZ6GhoY+fwlTxeAdZ1sD+Wyi4PbUVG+h4jUcMaw1spgpGissqQjPD3
HTfeAFgobzHDfe4JTvR1Mysnz8MlluSKlReBP/1/OH+XuyPawL1Wv4cJf/xurOkr
W8C8v4hzn8LxSqUV7o/Fz1OY+HtlKhiSeKzQQWf2pKdAkabxBTfO0WtyEA/Lrpe9
ylETJxo2iUTKY1DULZnq2wEzbg3TCWBUmOh3MqPsu2p0rbKT81x+bZl146KQDWg9
I671ttXD45BQtNRg7J2R1tSh1XTU9+IGvB3wb4A5iJ739jEqLB36LDVE58/xTedy
aeAwVOE3gTVI5mjdcarr0DB7ELca71nVWubvMAGav/LM/dDzT7NV/4DEjqEKzgDo
P4XeG5zG2uMiz/j6HbXJG/Rk7eg/Ol/vqoVMkrD1dzuNyAt2wyaoe5gncfBHS53u
D8FyGIVQLNwHA9z/ruhHpIDNtx9niHheHF4DDIBrLvU7LIpabSF4OcI/zC+KIEKv
gPzdF3j60VI0qTYvWzEeNMF5gGLMKQvYiERqeLZYJvd3yBRMBid0nG4ikTw4pB1C
PdvJhiLkjlfl97U2Va7yzeZqzXOfFY9aAJQli8j2jYWaLJMTyx4nmIsR+rDKAsTQ
F0z0PRty+/DFUN8JF7+vDovKT1h1i6eeSNJxXWOuE5mdRCQ6ER5A+aAvhgSge5aY
zFgH8niIxwWFG05JDtkn0s9PKX3+8d42X98zPBLT7Oy0YdBUWcRMMa4WFpYqBoTL
iBKqL9Xki3s+r4cCZBjDzIDMnQVASXQvVaxIckT9Rl/ju/C00K0jGgxvQaisydPQ
Zr4KaQuFNXpr9geDA3G1hWI6CiqqKcfa1ustwqRTDuIX6eQslEl7R66ToR4yR8sb
BG+aTQr3DzQfglb0YCFS6cWrKg6tz7n5A/c8wlRuzSkHAnvxkmxHgn/640eFEgfh
RC5AV0Eyr4cmLxnIqgeCIaD2wsTn7UHDxkk6eCGkJ8uTVBnIIyMHWZC2VnoCtgK1
9KZy+DOdi1trEbRQeVZ8SzldVzUU6yr1Tpv0qJ2ODHyairoosxZtB8s+wVzqdCZe
6xp8CqtJdboWHO1uWyK7iLEjiQ2GPwDPihTCG3ONOGuLbBGa3Ou788x4VVgfSyYE
o+dyeH8QuSIjX1MSF5U6rh+mwf/GOgN5BKgSKWODGhMM0t2ez+EDOZG0wB1ihFPr
sb9gtqhEFfwVMHuFQl98ZellRdauGenTgDCAJUN9xCdM6/+oGJQS4IEwzlZ7cp0h
7JEwwzZmzRckz4B1p40iHYGUUsez9FT74BNNkb8PtTDMeO7VXxRD+9royCK68r4H
+lrLQNxmBrUkq+Xm9yijvoig8FFftFKIvcspR5YYfqsGhlRdmGKNgW1aly3gTzly
DPWnlBfQNkjDWhTAdbdVDzRudwAM4iQRNS/QWpVsq4Pt5o3WcfgTZBVYr3bjwRFI
1KLikfqk2UxbPXmC4qcaG43tvohQVicmj31WOppfz2FuYf+rPdZyA7XqxrdQ5CFb
oy8VfyE99dOPTQmYnrTOJibtuOHEc6pyaxrhu7eaHkiPjD+7PWstD8z6VdqkcH2u
3btpwnkCFSAeyLqvwmtWQGL1gxfIMaWtcciXbTCGMREXWKb0SCs/SGFn6sgvt8Yj
3s+QkN5l/8XkwqqApZQ8eqmn+U2d7zrPpzpBTpbZr/jAUzTEmsvpR44z1IjhkJSg
nVNtFN+EXb2pPQrevS7eqmhhz3gIR0P3p+OBseI5q3sPgZadZaOpPpQH9yoE5pNk
OPc9UXodp/itPkY6Zba/FBGGWbi/28C6UDeOKTehE+4p7VohnAbkqAE+OvgLmYg7
KmZwVtMm9XezDSCBq31KsoTNeGjHehqoKqTasXMGhnErbDTRq2yAhR1hzgKyGkh9
E+17yKEAtw1VmslpHjGLJ9fSDBlmFudD6HOz2YS7Q3jN/45M9hlnrBcP1aX0OJ0k
RA0to5LoMCPdURXAhCukNLryTBlyqKQEoUoA5JQmM3FeQ1UYSbE1rTvVqKOokjJk
5qnpzVcSlYh4zOERXvWmgEE432ymXQkK95eIKpJx0cC78J+jElRrygFTKFsXmgHN
BaRmGz+xrrnpm2LdobIplAD0HuTvVWEDSEc4t3+gSVf8sd+83wGfxPUjVPwrcwnn
FfmoX+7kNl0NiRqSsgobcnQez7VsDzvFHQ/0ligqIqwvxLKUZNrheDW9FtwnKtE6
L36L6rRW7JsSPkq15bLmPTQ+DxYIdtXk2Ew2wXqFQYOPvHDdLwEtm/UvhC34ZmXS
EnUxkp/D4kqsHSPUs74s69l/lEzT5BqxiOVN4M4ro6aT6ISRi5936K+/d/mwCO/E
4jlNyByBEhyW0OdJnOC0ncrUTFFNlBBPlTWGtX9EMd+m60FkaPsZAGCR0rUItfqh
yUFE6+uJmj2DrupG6Po3a5BmkV5P5WjPqCt6zj3mlmX4zfE+TZyhSgfoh9fAjgr3
bXF5pOinBi8f67SHd6y3+IASqDheDicJUxLmIixiImkPnLuViKM6KqHg21kT6T3u
l4mJ73jT9XAmQ0P2pQ+Fo5gLPDDLJSL0XfemD1EXlp0pQ6TSpFbinAXtLsG0AlLl
UfK18ww6aprQt9tch2Rle99QUAIxJTs+Q+JZ2rmJy6xpGADyfVEo90WDQDpk3uuP
TSUEWQmSL+TE1tmjn5ZlODxHgxbIcrmrW3mPwT3eqFpcZPnFkFgS5mz25fY/lTP8
SguRWCPFOEO2GtRD8lNu9oHOXb1KQKBCvnAbPFaKVgpxOPXEwBeegNGf3UR0/PS/
dZhbBhECObihVLddscTkT0uhkV+w0O4Zsrs/WUdnSx2v13toSClJ4Jr+BdEFjJb6
OkwjL9X3GkgnREBOYM+Z6/I7UYzERm+So0jfXyv3cry2N8zpTahUPXdFPkX2MZnF
YVtVYTdT89PvNztFFKXU1e4ynBuHaoeNVg/MuG4QXZQNqOL83beJlizPqQOVvyaY
Wn9sjhpLhOFfxe6C00eEbTvlxdpkKXmQPoyeuWZFIerxu8uInVZIY6eYTyg1i9u9
HdacYvZA4mPHDJMj9vK6i1NuzNJAMolwNX+Ry1qTfIrU8ymdSNQHDw/8KrxJ8s4g
VQxUvYO99WxSHI5aAEOdpYrKe6Va/lW4ICO4hVNk8lLlQWBmiMXyECi0MP/FUvxU
l4TmQpGLg4cCczXIh4nB/knCfB9ZWQXifndsbQliqidaT4IHBILCdR5QMntqqghH
A9C8+0HrrfgQI+2xPyxta5OJPPHTsvkctuxf8Rb7+vyrqFRm5Tuo5yWbFUC9/khj
K0AO/d6QuzaSxn45SeQTFANSuVpMxBaq7qNwPV0ooNU7hImcEaOkwYJ7NB7RUf8u
ejzv1rFUGpC+PQXWEb3c8I4+xsee7q/g0vIwRddnB7JFgg5/x/lcHkDwZ7g7lMHC
IYJrDGetx8svp5yFaVFk+ql/3IJxHkyIc5c2fvkVTOudjR3ZdAoE5btMkDroAmNR
N8Ks2Q1nX92SYs9sh7BZ1mfsXQmv1wrXxVadhtJEHhP2RcQP7dHGeY2F6SOemaei
M0NZTeRrYYC91U+qdlZ1pBsWOx0QR5KCbT811uFUeaSt4jEcknnAFhXFxa4Z7GqL
Nz66ZEa6BKHIzAnhhetUB6y8tbdzgUV9CRtcCl4u3HgQPMTtMOBrI/T/e+UmsLGQ
jCAr60X6PqbTIC6zziF+k2NpO1yZTXjDgNp4GrE0jvFOkKee335PmL3X02eSUAvc
WQwoq0wOkzevNRwpFcnI5j2GSe3amdSI7KLzywhfu7e4Pil0+yo7fgKLT5n/1I7N
MPQG1qJpIwxMCpqYtb7cNVDhhEdMjOm+EXs9I0HLh8O4YIZa3PSMUoX8ec4cy0aD
vjarIVbF19/ZjI4a30sK2U28OxWa3nbCn7Cf/Os4UuIpmYjIspuVrV+ZSeZkQpJA
9l2+el6M6GFwEk7ylYUC8cHb0RM3yUZsDcVl5JMycSP+WCfGlZMx21MbFyk/A7gi
y6MEqdEAdx3F8fiYPyWTntUhELp83qWk6IKTZxEIg1onK8/nh7zbZpJJfhFaPm2T
R4kOBXFmjLHCv48XRPxYDe02VHY39GiEDRz7pt7/GF5MpjcMkr6tHvQqC1QMHI92
F8QMSzl6A1mKIm8Ymy3JTgaWtrHyWH04tELhdWHkUoncahZx5ldfFR+bMcVZGLiU
u1uO8etEKtPaBsweUQeNWXBsffaCtC9kBZ4G9AJ+E8cuJeOVP84Fi/AFLXfUQtMV
3ht4s+v/vY5xXClCaGN7LUvMIN/cON2RQ0p2PXcMaCyyP1EU9nbJRqPGp7pZY7wb
VWr235hz1G60Br8QQS0nycDCuYe38aVRhVbrcHUOjVSMfHQrTPKKLAG22oen4QBy
JGeRH7OQYhykOjGV5z515gEYcVIVbiCfbSUlihcy7ECiykx1nF3aq6+1GDnS7oXT
/sF0RLu3GgX9tFJSPDsJ6Uuy9Sijdh0hMMCQC0RTBNbZ4bccZnUzhnjqUKPUmRy5
FaeiTUTuJp2mmBuzrjdErSyCeqo82dCClMRE0AIhtLhdALrJqUqQUMdRS6tRf1qo
yIrMiWGlVMazTaDHBfGXUqZsDS7eYkYK8nckCGR0CRyHnSdrZeX+kEWEoQtybKXj
/caoC/t/6qrb2+/1UBu8JAGYljID+aNBTkJhbttbySRHW2cQ42kjRGaem5gTwwPt
tmdv2YDkZ+qMxGDmReRrPquBEGvyNKNoSpQDBDBLlspMEaVVOymjpK9E89/6srW3
zoA9kb96jPZMr6ij6MFfjkVVQu9vtqIxH9y3vGmYbJzzzjcphu6fRVAHI4OJEDpL
xmkUniF9jfdb8tWn/GTy5Y4+xEkqstO1EnGa0DmcK3eDsIQRksS55oPX46g3fH1b
a9ySK57JYFlxSJDuBx0ATpBKrcPOigHnc4yaPErq2JpgpYHdwuPW8Ogt+fcQksq1
72D70fc/hNZe5x1/GTwPgygtFaCnhrn2lR/D4fgujsYoaL8gx1whn/WNFY62gCRA
DKWMCtjPMe1PUatt0dziGtqboKW5VapUxWUO7qd4qHCOcXC3rIcYt1ScHk6iCooT
Xc+O9I3oBPDgm+vmWKLuNAh4dPwz8Ef4a5jw9Ya3b6MI+QJsNwdoV2lYLqYOmnhc
qmOJIZyhMhmjB54HyfMb8wjjW3HX1E1yR1HmA03Q7sscG7+Ub4jD9UNWrV1iUk8t
+75TRSTksgF63KF/42OUrQo6Tskv9vGQVlGNKnvZNcyGyMAPa2G6lWIvulZCV0zA
QNYqD8heLK5FO/xKkC462g3NSj5jl+zi/4fCZ/Ava0gPHGFO1AQUFeMVEGQEexaG
SB9dxk9aGLbnuz0imDV55i9suO5FGCkRGkWq/so+FBcKr5TKJImXnRWhjlL/0KPL
OyBjxnydWFnBvWYAYUto1g/N+JaQCnb25Q75sQZ4OwTXMw9leSro8CehqbZwAw5m
Yetz3VHLPR6hkI8xHeZg41DPvlxzqke1jWJyEJhJIVvJdZ79R8gYn51AnkEuhFnm
BGFmWm9Q4PjOdQrVYkW+EclsRAPfMp1HFLRL4GvzQ2i0xfFNBFPLQx3/jn+y9Mnj
tVKrGunK1iSkFQXuzC12Giha7/Z1nBJlkwBfwD7GLBnCfTzZP8u/0fsIW2Lc3QCA
bdRVEv0cicC+rknatC/seBDnHqKz/yyjIRTQL5JSFUvm3UBl34HId8vaEIrgfiKR
cgLKVvOCxekCo1mWp6ukNBSioSzdXlP38hHqM7P04nzbscnnoZ5e4hOCXfbF4Nbw
Ag/l5C4rDb5u44zvENAjeKq7Qhv9bGa703nvEnCpEXibMFgbwCJLHs2IKSQei2az
kbkI5m4KaiDBVI10DuLzUciFQFt/D/8QW3Dpi1g4gTw8YxSKASQQ/w6gtlVS/AXy
ckGwHGrRwQSD9v9Ytp59MeyNQfjaYfChnR++gJuwvNFKwNyHzDTKLLQhPXyxvvGg
GM9asK68/kdP5/57dpCz652Zp4ID5g4usq3IR/LDWjG1bZxpcXW8gcLoexA12nYk
iYu836YSY71ERGkGrY4KHoXShcmAE2PN8+4rfxiQj0tyEq5gSEOMfXu15JElK9Cw
2EOXL2K/EFnLcP8tjlLPEUBMiVSddi95Q6AdJykL+1zGPJcD7qAhG582bGuPjMzL
Vdxmef+a5U/CrbPsMLv22H+nZb2hclKLJAOAPXA/tmCizaEgL5cnMmcl+HGRYxDV
EwCSYuBQEi4QSWVZ5uynDoz1Z5uWA/ur9jYmLnR/JJ1qb5M1H39PhDfX8t7MBWb2
z1w0Wz1NabU9R0/lQdngXWhRiop/yMOjIUQTl7ECc6lseCce9DQbPxo1EIIU43aN
2YoMBPdZNfdLpy6msT9pgnyk1l83cqUIr7ErcDCaF3HG8QVd+aSUq90hhYNb3c7Q
ETbn2s8Qe9dukTvL6hX6G2JhUu0aYpYX/Jnh9NIaCUXi2Ya11TxV8syR6Yvw816l
8RoTw6EvM4IS6QtbG/idNfb2OkfwaMEfM/D80qBP6+wn1yhQ2cGYsH74M20aWfVk
bJ1/bjRYUtaxpNtD+5WXqRew+9Eh5OImle+VketceQtS+jQjjbZD2P1NGVd/Ttjd
F4TXNzZWa0QMpnpNnXfYO9yOWoEjSg1/27vcthw/dMJDOQ9WzYWYD2k8D+ss8IsV
luDoCZTzqTLgjZfmbarovdLQ1ujz8rJiIODrLF4tOPARQLa8z+7CSUvzIxUbokSV
iUWD/z+Gg1AKyZaSRkOHfbhrTnw7mZoFRU1KGlnbVQfY/LVrkscZ9lJU6RANITNM
GLCViiYF5RmXq1g7wAhPLWicNJY9g1GaYYu9/QEox5Cln7Tr6xryqqRg3mHeCa49
VttGi3SQ5uC/Or1475Dj0FJQySUFQ7saHFhIU9GdQ4S0R6Rg0veH5fXQLceoTTb5
3rOhVOOmq/1EYPv/TJ4/+IaKpQGHGFva2I0MEw8QEhb3mZf/MA5Odmmx1rYy72zu
J0iak4dp0dD3V572wghJ1lT5uPU0/fgJUMtW/GN1Rgyd+Dd87pmktLwG6JIMp71h
s51MYK/lQ8h5d0SI+c+4M/bs3xMAINfHVGH3kImpwURf3nQw56VBe8l1mUBk3ndb
MvOV9P5R2Q6Bn0W41mw0yNGN0rWkMgdCdRodiV3J0C1jO41cIYp9pYqMELoAbkBu
ujxygp4jb1cepVRxtV5nMJEyjRQyoqdlt2mmPXDFvGPxjnp0qjtc2SwTV38YoVY2
xD/37PhYEpDJorTGEnzBawA9fpnEwp7+epImSaWl1vL37SouDzocv9Qaks3PGCwA
veNSxVpKkwodwctrKG+Knsp9t0ur9EEisEP5NNSE7zzMX6DBK6/UyHx1ByAxHzrE
GS2yye+lbsx65SFg0Ob4WvGVTuDAUZSnzX3xR4c4G2ogT1FUYyzdGE8enAP/qUGV
lLXSuJIB/A+iwu5JnN2Ad4udPKwlRePs4nGlv5dLABMYoKWHg92KlRXw1X0pBPjE
YLrSV4kOzoH3HL9UUJkD1uucvi5SW67FRGO8O9WipjadH2sLvlpWmoiA8+a13ujf
Qmc0JnSRorUfj5Se8Fjf+wG2QrlYNUJ45tfBuPjwTnA06ExZuaJrb6x/YrKHEWrr
/RKL+ZiKZMNd9Ny5a8reqZs8oeSQ+gM5yfvGa+Toc/3TelUN4QkWE6FWd7wWJD83
WhZ3znSMcrT8qxEUdG64csbauk/zNpzhh+IpX1+zzhN2Uo7tJmdJKO42AsCtowKu
Tqa8S6BLmvxBUYSK+JnMQftrM2R2sfWEqohTmmoE6D7f/5WvEC4mS+25coq25IKI
M6IQmcgkHF0d3ym7ThX9C10u0NmgZkG2P0S3WQVjeVzcG4wE7lxY0ptW+qyDg8EY
JtnYQxvshE3i9mOIcTVx+c8uJ017YAtmhopNw/FxiZa/aBtzYHfCUg4RbziX819A
5+BHvXQ6bePyvoMfjmz1UVfhbAdu+bQbCBc4JnqfO0AiXE8cOYFpZyzEAOZz+nLN
wptAQiQT/dY02zEhhm3Ys7A8Gsc0/HlvUPKYKsvjPlZKUY0pgH9Y/hA8FJ907+y7
j72uePAeZfctazpxX2Gi/rko1XZuLI48QvEmJpZdjysV2pmZd99FoBNJrIOR+aIr
nezAEeMbk3vXNw/kILCWe90baVhJ0mbijdW5wz2m+YGUjD7VbjZE5yCJPFUwRpWp
3GpFg9EUq8G15E2+bxL0tr+wIIEjZeFlNZvMJBSolH1Hu7uTPD5q/sL1zfrXzf32
RE9y+piDaBDcgzSneX4JS+ycdrpF5A1GsFXVDaveia8+/xXZyoLc1ajIanGtOxhr
99LeHyssD6+7QsEBaK+umnwZbV+DG+VG/dGLDFmwgchPPll13AnL8b8XL32TdcUY
Sz1BcP9sQz/Tb/k8B3PfEB0Rfyv6ZVAnRZiUe2/UJS9ylj9Iw2NHxQ3U9dzWO5a2
PIrIxWDsuJQ03xI2PVesumgxWxW53CaAPfSbBuS9pit0Y9FQ0UhG+qsEyo0yjXj7
ragJTedeUSBDpsbqOZsLb6aPOsvmWUmAk98wjalGFp9ZXaOL070/oupnyvNA1MGS
JgCioZBk24OIa0qa36xOFivwoBWFvrRsC8qrrzXoX+9FmpUtvScClkg2DNM1INwQ
pdYtaf0WV53+cHIYPjY1/C2jjJFCbfcKzs99g5OKTM9tsaZ3tJSrvT7dDePD7RMW
F3Ww8DMZzvlYByp7IPNiGLHpLB7PrZub1Ebf3V1wu/9gjELJ0wnMusTnjxiwP234
xR14uKKcmFImcYgGgYxyjnV+0YmTXfOJfe0dAxODcyynb91YHfJB8zei+hUW/5iD
bta+X4a+zOKVNcQIRYZMgutKjLePJmOF4rwPBimL4QzSr38c7W0k6QXmXhiN0ikN
DLDXy4wWeWCP+yVX08RGugCJCldphDKYWGKTxtDoWjPZHkbiaOKvtjtifRJpY0LI
QKgSe5xfEGpvl3MWpba80gPPPOxVnEr/2gmIQwDYdvoxlkB2KQvxIMECTfg4n1lc
3dIdwc0Q9ShFfrZJYmJ6VMPPwsBv1muAHt8mdGRdHE6CGO09jrXYkrAt5bPhc8j7
x60wqahciZMeaK1zAUQ4Il8imHd3fIKWZ3H+xS5tJTg9+ZCD5OjLDA0Z/LOg5mjD
iEtRKMr1D+7duDlklVuUGc6cUMdkPtzGc5mj3OrEkdf7ZNshu0wDTuzJbbmK8zk7
ioko72wKeqhgWiis7LxFIGw+UwBVs6GRyUbDMN2lvJx2hldzmf28H+SGVX9FQ0PM
LhtRZVZnBpp44qsBkD5CK8f6KwbCN8ZpAoKh1xNWRHXRzKPsw08RHjy8k3RCT6O7
kYNXOmmFIxXnDoWdTZuvZ0f+sjT7sZaoXA0YBris+K0lBYDF5dBBf/wHMgfVwYfH
0gC7O4JYwuz3qbS/1VfEwZM4bF/YVm8uVGOoIR6ag1Evoat7LXkGQvq0m3his21h
+wqtePWC5/eMzADS2R8v50gQzNRbUP2Hk/B9n1pkF1Qwvx+/5Oy1bCYNibx1/2SP
KHRg7fhgnv/bp5CgaUI9AH7EvxqD5DDJPVnbrwfusq4BcB4lo2NCdso3sKV43ZSR
87pEH0F+uiJW2UDAoS7JnOxlX4s//nn9AWZVCgk7M8IFqncM5e8MUfF5NN9FZ3x6
H3MdZhgrjU75gMl0p/hdno1uNRCp+qicKppM63nWEvr9rFAlHUqP/WnJn6cj21tn
oLPNhLkApv70So58oP+DTGWO34VV+WUTENDri89hLhXdlUb3F9dwXEPKqEX8+G20
KOptUyHoZEeNbEdqnCeClvFXilaM+jyZYQMQxAxipcJQ1nbtjq/z9fMCUFA8umBU
cxhiq8aMmsb3vaXzxS+FK4zvUDqj6BrAAz7IGOb/FIbnO8/LqHoiw5KHpAuRwu7o
qdRIZOIYaMPt/IjYjUhTxX6EFo5Y6bYg6bsAFP7PYGGTHRIj0MK2Lg3QKfaMzy5B
qQGmNkLBf43a1T8ssGUvcV9OMZG8kC6b1yz9gLCh/XWzwRfoCKxjGxz5mIMys9UO
ArgVWgi5JzmQTdNDnOwQzmAmIo+g/ldalOzdWqD1YX6bosQukgcD2ZfVFdlPtGjH
egQhFCvCsy/U2xi9cZBBwXBVAwklAIjirZhLn5pYr9Xggu47mo3ZTNW6WpsU9zzO
sYv7N6VeO5AM/f2gO9gyPBpPqOI2PjVpA84tLj0792tnBvq+xLS7/v9odW2abo65
PGiIYmNwobaWvfO1hPXDbTPizpl9SRe+XBMgnB1tD1Q7janx3mQWpWqhecqDLOSS
Dc39ckrvPhluzx5xAAYO2IxQwfqL0NzUQ64p6m0OavveXfCV/9puXUwI26nLQzCm
KVRGGgjQIrVNGML/a4HX/lQxMZSLniQ7codcP48fda7TSsN4qbn3tbbrDItGDK8+
M/BPDB2fffpf4uDXM3VGVbv/sMwlz2ygcu67HIKVLIFfE5MN4yTsd5wpeePIVcwe
RSOo4/4W+Oy0gJAetuT85HoNKqCu0nZxPPstfFnJGiSn5XXKbPAu6it31dFihK/9
2r/a+5XXjaSHoh8IBODlOmeOoDWxcjTgFaWxuKr0K/sRxX87rpsxQds25or1mHiS
yi9K6rcHzs/tKiQYAqjKyRXiQ6Q0LRhUTyfYRtpFosiigYDFtRyM6UYNyjQmy9nw
9TfHxAT4vpiROT3+V/0fy4YwA78fHx+HMwrlWdGdZWnF5us8Ju73dYErRuE0rldL
1UeTY2IqZDt9v1O4S5j6ODQw3jJG7ORRAC3uGUR9BboWT6ZtSTMtTJi4tWjhqp14
/mpfGsa/nN9FWu5ouw9dxHUrUYNPfth9rzhCOb5As/GTmvPv4fZF/nQVhwnGUQJV
A5KNiLPneMHgrXsXTM/Ty2QU657PFYgKQBxue6jxqBfCoAzHaXUiCgRtvusz4v9l
jGK1pJ0QZv4Yw4Zt36cAOS1durz01/GMTpd7WZvLfA1dwdngCjcwqhrsh4N4sHvB
PkaWAcNQrUitefdAsKgcjboqx4fLiuLcWNFj94CQKVDVxDl1XgjRQl6pUrHM0xTr
EGipZqEyL8F0SD9x2HQY5UIPHV0xRgWWENYuj5/jyVaRrLdRQpWAmq6AKSxwPuhD
Dyf4iilPHF0dhScq9FlHINTgrMg4dAjm2FlcToiW6Fx26R5OSG9B2/M5+S5iLR5w
5TsN06120DQXkmM9vQp/ZNk3eqP4vWTbkP9j3rbP1OZ2o+BsR+JRXBuRREpUXtgr
MSEUj4uvDyWNXk/lWiw/FfbO7ROzAZt68BoXrENxB9fsLBGhZrxuQRc/rVe3wB3e
M0suCVbdSzf/ppE2OILNXqy6DmR8aK8vb1zvJKd7M08s7MvXFz0zvgs04w/bGjBv
mGTtxVnhA6BHvRNwKJGOwQ0CeT+VB1L0UC2+V0Hdooc2Y4IRpqusy1xZIf4LDKzu
gLOid0VucW6xTosUt4+PWwbWsxxEQRyooTPSE3D4a5Yg4yp2ITvY7Ah5ukbE5ezF
T6R5Q07e81nRSWQX8w3vCBWH6HCSfMXIqLjYEeo5YnNB1v3Ko95cLxqMINIrXHmu
sc6hq0Or0ycxz2kCDemhhmXR9obIVNQF/Qam+E8sx3jM7nrQCKEvwDib6j7e8LEg
VDsIpYmgeKpLcItp7VYW/v7AsW+Oo7nEMth5OLzACQDT2lmpzqSxT7HOyv3cIzME
98gVDe1F3rjjvzKOV+BWsFHqW1mHtVLUs/BOLRhenfX9nYRR1l/JJl1+O5Xn+nH5
RJbQdqy9jN7tpyq9qzPOj/a2l7Jv+7MLe+cdAzfwnoOwhsAQwAmiOrEwn52V808f
+9SzVVIywkJChXKCxYDb3b/6KHIyTkV0N4CZSKEPFKgUuFgOsWRiQHjQxfqaO7So
dAEOQQGo2L8vb4ligR8kjDRb6Q7QixZpslDk4Kvzq34Ks4eVAS4Lj0+vjqLKpL2y
zvU/5iHxMGYtQllrpxkHaWgYx0kQgN3yfZ7i0KtFjXiHqYbePWwpsGWmB0JNYkyU
M2iLilHF4U+lrVqaEzRosCfjvx9LrmJBO3lSzc8KoS/oBrzxgabFe1YdMB97eStA
AMGPHHBi5nt8Ve0oz1pGb4lNTj3VMbCWQRhQDn9IXueZoPM0zN/nSHowxy90WXlH
f1kyvhIbZQ/wMrkdKkjmTm/Xcch9rrnPt9HQhz3kpjY6GF8z1hKbboWbUL3UbEbh
UWuie9/vZDu06OD8BNHmtTF7ORxHl7tG59DasTqKOcm9809ymmKV4dRM66jrg7z6
pLn7luhkoeijQFnF0dALBQywS8/yvCHQbJ7r/5vg+KBK+ROgaQtkd8O1T8BWqlrm
Cm8uf07IkzREvqbBscxT8QNUwjBV7n1wrUfulQrdpCbmm6k++01glhXfSTyoxsMM
UvgTfExTMATJhHnfGvD5plevnSRNEAhMUlLaPN1u4BFH8X/waAuQGOc+XZhKp69V
wC4oWJ3Ad8TaONaFzNUtJIwrVt4GRWvLnRnbyCtP/HdvUBzDTftxdsmd2wTpvXYJ
QAf7iTsX9AEbWKo4wGTzrP0ozxsRY5/deb3H2uAR7k0lY+kdVsemA2LYgFCbKoEB
6Ylo0PqMFCy1NsHWuRMcI9Kx6KluT5OsfvIxiGBtWcyCStGpt/zFxjPp2uN7W43v
BF6vqEqaAMX16EAdGN4mJx6jml2ha4j0FgpAAqHC/eKNzwWJUm5g2XVLAhWiRAvd
E+b5pTHpPBLcRQU0GG3mt1DXy0sDVxO0Vyc4aBQhNtvw10fbE0UZfuN+ZWc2e+Pw
vHiLwb16trpcJWHweYZIn8pCXoZ77Tciob21XS/0rXhtReunpUmiCtT+eItvp/tE
RZSDzKsRUnTJcAkKGvEYBWTH3E4QqtOBoA+XFJmY5tBANfucp/Rz3QfmRjujvgmx
tT8Hu1Ho6YwWGGVWrziKpX5oldb+PuwAl+0S9xR3WTZSi/oGzNJTbR3pvCIVJwYb
1ClcqMXLI4tIwv0hN/+8T1y3JPt60RnrOVADnUk7MYP3Sxc8olPSBwdCZmXr8WUQ
DzX6+Gh8H+8ZMIvHaZLzqPb/2/JN0rSiY0fbOsCOXeSOjtyjbbuo3oRXuMbaqROc
d4IhCon93Jdv5U6RycK2eEAW6kyh0FVkaIBIw0WIpR/pMmwC+LD9bVbD3x0F3JGO
Z+PFzJRaWUfOIFbs4nlX5IAaIr8SRX9f5JkPoR6ZhrCioRudXgDm4ZSrofb69k2h
erLan84xtwIIk5FrCiSkfetPbvDk6Rt+AVCMPvXsOMEM/fps+yUlXZMQtAgqvUpa
9lArU7EU/8svAmubryJt6Kj7G86sdK0FWWX42Bsv+OX02PV1vUhT6IWQeDPMBi9N
g5pMkH/UyFveB1xtaYRLVbilHR6GerLFtLsT54Pl4tnjp2JykCh35MD2NYTBwl/z
sSjAUV4SWloagSjkqbTwJSag3VDdrFGzDSWOQmgfHjfiZOnzubRm9NstD4XyPHml
unVRHvKVTVnJ4QWG6dqa1oECxzIwL80JGUGqsErTNBxBQodqslmCsv3GG9trFJdH
jh8WHGqHFkGuCtL4WtuhKqP5XjYg9mfPT2AtmZrnHsrSm2U/+4XHPSdwnd/XdXRh
thCo9OFRHJvoCjV4yTHtA8G423ncDMZ4vvXSHYi7f37cB70YntSithP0je9jGP2U
Q8RBgPaWQ9WCG6Min2TX48QCbWX/DLz2E27c/sNo/ot7ckZBle0HH0CV1EHPbyq0
RhNHBWTsZq5IDWTJ/b3/bbUH2NuDtsRrStYlOIirFZ1KfVUae13B4QLjKQyZrRSs
YnLt38GItAVf8QYlgW6Im+4NI3tg4ax/d6kpqOj8AUgRv1B8VTATs3WikuTtg5wM
JI8kd/i+DLnU5VdGaNPHcL0F9bVCdWxbQxFf/u2LopRtFsxS2CsMDce3HxynfaXE
mIPSTJdVHS0KAiqqDvvDYHapAP0ArdyF3VpAzatzM1ESd1DoHv83Vp5YHGC8HsTz
sljSg1i1LMt4HAJPizo1VSttTB5ZZAQg+gTIqUTUUJAwINZ0B4n+nRadmkA0nogd
vqIBUQ6X9eptq06/Zy/ZG/aHFoZb1Px7HIZ6qU0AW4SsIsNuJPv/DbK/V+pZfmtW
7RGgj8SILS9r6tsFCEKRGh2DerIDPNf2YOysP1Cq6PjcfRSSuCZJvcgGGBvMkNRu
REFvveRoFgbjk6CZOIVU68Zim10M8OUZA1SbtHJbzJvYik8moeAsFMY3Akj6Bw9X
7aBYr9b9qKwa0HfWfl4on2HzK+6equ+H75swrdVwa0iK83GNXLtylvrz9wMA3keT
Bmj/QmXAqWZHAEjqwM90jVV6c/4F+WxvjGkmRKNj58xv1BzHf/Mcps0r1BaGhxAO
RQttmBOLeeInxxjirlYGqg45j6pXHD/HlSuJFRvXVS2Ul4jP246iSpIdTJMftMPX
oK1xjPZ4QK604BNhU9PmjkCsR+qcQSoj2QmawdRmWsIfrsCDs06f9mg8JvSg2/I3
o8MQ4kzy/fc3NJTwkWX32qgJFdE/7BaMlAw/kwwOxkVkQFnnwCjM717uAj4879vM
wQz0Kxv4aJDt6hlRyqQh3vQq9Bit9FHauH4kqnF+4NqiVBWa/DjRNbpTiuSV8wCe
+qnFEER138tmLqKKl6v/JXvIJZg60LIDmQ0IUR1GZFsicxUwtEKAx1B+NRHu5iOi
K0ROCU5Fc+1CueBVeu8wtzMYG59ilGeEtZh2N56cdU2tdKMDm47NlEIlgWQeUHQm
YuiLF6057iYjJfNzCWBaSBNgw4IFZ+Mas2f//Xk2sZ9pTclDJniLTVOzxMqQ6wfF
A+FUtN8jmIa1p8Go+F05RfiB7TExkRouYyshop+9pdjtdVnyyT/4FwEIo9rGY0Of
QqIkufyl3nVaVy5t8bV3ephLWf5CMxSlZN61WeRgBv9crc8qurT6rrgoEqyRuyM1
zu4PATnM7dPq2eh8EpN8ysvqZUMYpvi1HzkugeZxRdJoH2ZU2HqFGy6T318qEYsG
A3rcckIifL41/+OwJrtoJW89McTPCzZlEONSf8KnJgbsepMWUZSxcOf1c2xh2pJj
UhEzcEYlNb9d6PbrMLpnG47cUkVlhewpjW6NXE2tjJRoLQLGVWervwScojjXRB8U
edagy1JhYXttj+03IEE1u81SWotDd6eyZctItZANycE1E2dpRSut4mKYvNNDE2Bk
7trK6ycAXdmJg/COCwzUdVosSJtCE4YrFx0o4EvkPKGvlWiWBcgjqRsfZQ9ifQol
ZBQ/p1osl9/CErlx3okjRQ1mGqPyCVF+3R1BRjjtadNDlAzh+83f6XK4R3JtKWoa
0DwpTvxjWkXpnbiWCB+uYPN5AqPGiw6emZtPxWV26G4+HMb14FAasx7Zz7bAAYd6
IQk1qqJ2Gs+TwhvvZI29ghbw6+Qvqo9JkgcaW8DVokobdvxoSDVuOd0PDeU03trj
ab3W8qdepUNrSl4W+J3rLie+iuAzd9u6jTQ8W5vPJPb1pElP4wvF1S30wYv/tTQB
tnMnjK1pv3yOc913ZY5iUT4Sd+rk1B6co1RC2BE+BUR2BsBgcyeza9ChEnB/0iDI
/7mNONFc8S4xQ5OO/iLEyVE/jxZLYwiHDkz8+w08c4UuJ/m/Bugwsw/3c19Ii2mz
CLNFLCZVlad2b4qG0M82HJmrDNCc56tdC1oy0bKOfPhZh+/IyU97JJIAEH36Ee9C
KefOyVE/3PiA9u+NWV/8mTvCCoLH05RMAkNM1FEer71pKHVyAlz5phHzpGAgcD6E
NsITmjVD42ZcurJnUWy8WkhaXDVYy++S2Yl7n5/o39sYZQ+cPB0sPHA+Xho1zQ1x
/yoOxYYUDssisoKcN/5983t/wF5ErhLSZdNQMhngTcGLYZBfSPqyiKNjR4jZ3U2W
T/T5WPdEI3Fs4Z3sxFDkSNGhE86dbGTOxqLqRng0JnJZCkkRlKLa6IiwkMbek5Qg
awjBeYDF++DDeSGbD7I1cXlB6I6jaf2IyvxPpeEbtflRuwIeSfM+T5yGZymRTr3R
0nlP5ix7oYl6sQiSMyx1a1GVw3fVz+03LvTjv7OM5PhwXHB0i9m5DeM8gGXe2Ckd
iskcHV1G29N4EP5paCTsGJRXHO9XGQ1QeSNF3d/jhh7N9x7QTHfRWQtRZkEERTb2
glR+jT2n2cFiXAAMBGUagCps4cHjAurotaPWEiqJrKYMQIEatgu29ZX2FWhV9HOi
fLD1D1JJJoNHtvmCJ+GPZ1keaQqI92WHGKoEzJXznjdzUREArdJz7INRWVCiaMyd
bn3OhJc4GEf+j/gtzZFhpgnLByKCbAc3h1oy5gEVKtCQn5LPC8opZ9cz2vJr2XUg
T5y3AV80URoHkiFKXvdFhBKKL+KQ3P5CNV1a+htDs1v5ZsNaNPUAyTs2SX/SP3Fy
7lVGhzdJB9Zji65gFO7Plf9T1lDkwCi8If0XYjUNy8oT0H5xaC39tGFs1H05/fqs
EmVvAIQ1icOHzo4ZNQyJ5Ki7ZYGuZiuQ78oEv4FOqe9BGRZQMcxWc3lb985ejSyv
6MtQp5qUCOHHl6hQFAm0HzcyxWNgtSqnxKc/DXVxPyEDokHWLQfy2ac2wGNkKUR1
JDwd02YZPIrEA9QcTjVPu/QP7E6GMwAVJlTt8QM7ikgnY2klba1I6gyJ8S/GQghM
4kWaeTztpLO40lhV+hezecg6t04SmVLg/qiaHKAavGAxzruQ6xAnWWb9/FLt58Yx
aUsAsT0XtVnGZkY1hNUfYLQtV1XeMw8iGHP3Ngfw6W/p2d+tUMbYlqFLh204sNW8
WDZDfVgQqIPA+n3pxXZ/z/GvZPTHOBfTLDBVZZqKRFZ9w9CPlSriHKLuPo/lapWB
dXG7vfnftpjhJ0d5SVSR3TpK58Wd82Ty/GJmYnGECh6Ts9JSeLQKwyp+UczEojRZ
JPQbhaZH1YF25z++aRvprQI4Uh3j5BbTSpMuOJ9B/dnrHsUgzAWBmXY8pow6Sv18
/EJLLltlZTcCI15bRJFBhUjbzmCpPoJCHwr+TZGVf6qsIyuDk7n1HYxVmaTkvrNg
/1Dde24gS1rGIEt4N78U07bxP0hEJmQlFW4A8Li+KVLckQuVOXW09hv4quaz+ek9
OVPBKxkpqbbz/o5ZQixDNTfstowGgd1NA+x+D723E/uJym7gs8SfJURm51V6Z6wX
uMO55wy0hqFkERa0A39u4Bsj2WAbsOfDMoe6JbYqTUsFkoIiaqF5yy+aoXtqWe1Q
W2TW8TADLgogw/rYz8Q9y8Ssd1fpWb1TgftkjmTCfOYean4pMcmGpuFKAmEEbXma
9X7Jpc6xGyHG9UeONTi7pJpn4u8z9fybkDWQ7FPQSa5943Kyf4Qk6m6CP/lMRe4H
HG68Wq9U0r2tIC/RXuErSY+ScjULspx5YTYxwfh97J40LwjgTAL1tGWVH4j8Zkg3
+sJKEMOQx4KQAscccqKyxfKwkzS6dABR+KBqpGfuzIKJDjC0+Lf/DtsR47ufF/Tp
MB8kBr2ra8S1sbRenPzaTpMynD3KjbD3s3tngN3lqxvJmpAAgufdH8QjPMHaUyTY
87nagHU6/ECNSsnyIBJFMyS3inrzsmxCpIBYx2lUJIkBqX5jfprZXwXI4rA0krCh
W88D0RFHJ+BvznJDbuED47Ru0eKn30GDIRGMBGLvNOGMoFgGYrF+V8Hbr8hTRfVm
1URMVQh60azXU8mmLQrTZb+FGDpa2SD/9aMnvQcc6BFbHLs/LWVlb8mp1Cxc4aY+
Bvm8H7SSP0XeeJjnLgFBYx8D1BXDxlh7Vj77tvd3KVvHLCGWolbY6SIyZ9SLtvz5
64QoK2KimWrBZqHYleK7CBEoUUSlTZZqRJ5nB+uKF9lUiz41jDQaKAEGIOTdrOnq
SEPm9y6gKRCXyhpVMoauvhjQpG63bbHv4G9vnhSuLmZxYEh/vZ34XECOy62TU19U
QeA87f06xK0BvY/Ayly/G4o8TlrvCc9kxe23SH9MA/930eVRzjVj7sk7c49ivWec
vQFnkWLFY6LWlLOYyesXKgkSOB47Lkn/ZiCj5lQCjFolKJQGDmsOEMsIPjTK0juu
thAm/IXjcyk+zTWYY3jhyRhQE0VbCOb3dErCigsSR4wOngN84II8CT0f4yszNKck
wgOPlkKUZhW+Yie631I19Zoh2H4FIbI0OTAYTjTUWghSXsmp01cQqR9AFaIKW67F
dZUjQ7aIN+95D1fmfznl/i8YIwgRi5aBGiUTamsMKS2hrP8MgqX3rQWIuMLMHufE
lxEjH0U/nod75wZiRKH1qBouVqBoBCtfPwaVzipuAbkP1gl6S/QyEvwIK73VAwr5
XqwSVoew03P7hzr6+JUsFVCqtRuEnbLmn+xAf3Q6CWj3Oqq+dAqKoiGZOq467COT
aN4I+nV1XNDueF6XJt+ABoOZsCXJh9J+6O191p1LUdOxQZEk1PKmPh8Wq8v+h7WI
mNGceY/sGBfN0N/wDzoZVljhph8CGrt7Ff7AxvzpO1KjJDektZbQz84m/uE2eDz9
3o5Q9CFCBEuoYJXJYOC5tZteChPQb4dykYrIK3IpVz4XhzlRVfAcQN2SuROrhd03
6niCnkWotRaqRdxdoMxBz+s7+Ji6/8pCrV2nDP5guSWI5ceFPrFAXwCOAQlsaFHM
uy1syE05hpm0/BXpddN2KMk3i5cUIc+8gCbWX8l4ln9BaQap9GIAWDVOTyMVDtjn
2RfRk0i939pr8vacPKTf+10XlxcrYF1Fku8jFCgksslxLbYqoDferWFqYyUfnAUQ
duRDZTsA4aFE5JxUkHp4J7iH1XPVzTHtgQ7/HV6/V5Fz2j1nXC7SSvzdHMpH/PnT
RTfjgIwZKmbLn3e3Ihhlfqb7bIM3zTpvH2tiP8PICK8MW+eibC6IaMiojYpXXUCC
Xsl97SMgkxH9s3ciJbjvacYc/elkQoFNGbSjJUiQZIA/qCqMqJ1RHOE1o9B38DWA
16NX57vNnNNdpkRuDUdrI6+m3uiGAADDWjOgvtLoJNQNI6HT+yyGgXdUDqnVeoMR
XedgrBc3rxO3DmxCwA9DQ+5U0ZTZ+Lmk0KalZASe9PvpAIh9yVHc9KzWWvdN6qGi
ZZX8Kj1JJpJ+s3+yM4nEwI69g/a60jln8qBED8W9B8y7SE5s0lYpdN6KKHSrOi2U
0957cdL5Yf+HUkEaLZKhB5LBxHXLsM3/Vb7g0FtwEYD1rjOxy7o9tXvMFeNKjv2C
EsHMr9dVm5qK32alPrkgTqsaimnrV3qD2+7jibMLv5ctqq8Vsb9coDEEvLyc2qvt
JRfdnhW3wZUMvX0y8sD3yYgVNPgODi3pOnPL3XvLr2JO4+2nFMzPS/I8tgnVf+A0
gB/0t86B8v7UE0lEmT7cxLxkGnKBkBxgGXZsZu3XptkGgbQAfXZ/kgjpdvJbPZRG
UkdqwQfe8p6qo26N62g51iXXzHIf+WIzjck8Oue9eAELViJMa05GOfMoqhJqgyKx
+8RgJbC7qvYy9A5BUETzYGAPafc+1wkaJ0tQ6F8Nl3yWU9w1Ot8Kls19DNJq2+Yd
fGLXG3V17xB3a4V7CQhR5+QG37i4Z8ZHEV4PiogE/itU/65Xa5hGuQNH0j9lnPJi
+FasGjM+oK/uTKoRulWAXCzqUrwgNDQ2IKDf1WaJCYdR7tMv+NHorn9dui0hLJT0
AZqzMyYX6ndWh79asPX4QBsd3A90bpNgCBL4gThJt+uQHPXlK5IOskZIdRo6vLuJ
L7JqMyJIxD/lNDs+uWQWkYbqg8JCVnfw920KjCU8zpW7dFdUx8ZdvgDj+bzNqt9H
0pCm5grp0JXGvqr0N82P4awX1QdK4oOMYmyfM84lJ7+EQXVj2/76TXoFTEYcLbTm
5IgikUrK7u+aJPMXuhTWL/accyYPkkWNs8qZSK8X1y94uRRyuB/r/SbGnZE8dR0/
eMIPgx0DAoybH6JwlQ7UdimVPK+S0bqYB863KuzucHZY/YMwztarS/8X+CINWdNn
hdQRxps7io0RvOL1dnubkpDORWtBCDdpwZUIIILkzcZ0weeGyvjOgOd8xse5Z9y1
ZThhy+1Hxy0EL0jjgZhwAvz/QFCGb4YtH31K9Ex0nPubm/Rxh3BMy5fdNLnqfazc
sDH/4TveeZUC5IYQu/qa8mP0KWPTqe0aSbEH0NzVRKWHv3Mar2Qol5kAxqUXcsyF
4DfvPNM+sN+2jeIFksS2H5V1zx9r1dwN/QPwKfx7/X+qqUG34zeAADiHH19kPdJh
2WM3i65EYxY+3MVjLJkIJkp4/In82zUGZH88J2DRyT3SMfdQd69MS3zOd8kNsaH8
QWGSo1Jyua2GhotxHrB0I2bQssl6UVT+qR5mJ7hSzwoVEJbgzCn+EEpzQJictmpC
FcOhwHYle4p4c3hrWX1QpMGz8ZjNj8KJOn35Sz5zyya2STo3qPemQ6M6b9KfEWvf
TtpraIhJz8oIrOrcROypaP7yn9eAAsgbiGFPebnCwpdSe+ndssPQoAKkeu0oRuqp
PJkH/ni4atoA3OCKlMZj0gdYeFQMHJqFaZlQ9wTP62jO0fBFGLCYFeQ3sMRqxS8Z
T9T2T6S+d2Dj7upVlfUit0e90PPL43vm/nDzSEqVyEHFnv46b+8e60J9Ian/2/Gq
wc2c9F1rfBFT77XlJmfa+v6YRn2xt5OjTs6VX+98i55YumbJQuH4xcTjizmA1xLK
kuUwUHEjRRDlFp61DguL5oJ24CoDIIa1bU1QKstXLdw/4PJChZi4EbqXG6A6XRD9
/p+VjyfYWMfvdO/WFadnU1mpzHdIeG2Qd1TvhFU6IDv5LewIptMy3di5B0/Oem1u
bvTvxbYsI7EnoV+nMlNEiGH9x1FJq6c9gmSjIqt+Fm1WzpnUs3KZQKUsnqUl13aW
+N9Bwa42+T2Yb97IdImR4wSha21spm0wsKOgU39Qm5EBCVtw0fB4h6UtRxrA8k+J
W7Hg7PFa654hnBT7a1BO6CTpmrkZ5ixziUTe/5iX9kdSC/Cq4biDRTUmzorF8QiH
gxjI1Fo6KrA4EBYFFjo2nHPcTLmkE8eeW2UHh2dg8IzmB8KsMxwQu+m+S1A6VehN
gSc6y5GRmia2yxD8wNIrzuuZRRgc7o2jDNXVKpOQXPhBNiYObt1ovD6WyNTby/S0
V6UDA4KChnibd7HTEmWSTfnhPHy5H2Vk0vuIR766OQ4iVQ4y9tgj8+hIUuLNHqMS
bWPqNIF2a1LXtqhbI3IOSNMNBG8n2m/NrJKsx8dM62b94MpVVpzL669zBFOOoGrQ
2gsh9vJ6zDfNzaJebmf+d0b3nwWcMV+jDvhmFn8jFESIhZ3BTBWXhXzr4cjdAlc1
C6lnIICIrR5wkPltWNNmRN2RzXNaKx0e802cZoRuXJwwLbWqGSBvvoq4tYGpZtjq
+0sdC/PYshJQjtR1P9WD+z33zyxHxdE41riyL2UB/rkueecw8Mui/3Sx+jzQtATi
SVki+MQUcXqgd07AMkDARvTNnvTqmWdempsIWB1nVajGAH5tyTJjolqgNCv0BYDi
+lvScW9N3AxLZ9MDfG/Dn2mvlPl8Gyd0IM6qp3GAXY1nVfJcZG8/I4MUske8Z0w0
HY7v7K9UAkpYmLPZckDhfPIAGXUG2YKCecfU4El2Ef4JHMw3mEKo9u7ZCTO1isb6
dPq+/lvua6Ffmz1KqPdvo5dq5F0XjULHtZyKGITjq00jr0J5RVlWEFBH1+TAOuK4
5eZoS3n4BDelYzDLz5K5SUYhbDNJQYKiyDeez0SDEBqWL84niCeFDuv31tVU7KnT
al8RlEQpvuwDfsfuWXsT4FdE8fB7nouN/Hlw6+/RtRu8rHeFzv8zX2q9qO20elSC
N5FgxGTPUvXpbALBECWIOnoNEmMvmFZlw9YVBfGy9dRVCF3BHCuScwIiePLiHiww
NvAHbULpJifDseis/+PRNwPR3bZQJdP2U3uj0uYIWpwWpmjqCrvb8cLx3oXFNAaF
U30tA6L4VGy881l0cT+Gd2X9rVNGERNt7rAYKwbVPrr6IXLfVzGemnCF0xUSYlvc
hzVLb9HgAm8gY4YN1bsWFNh4AIonYDAZcNVFw/FITfqoV/0jiqfxIr3KSgD3bfVm
VvqtDycNPogUMuhfv4MNj92LGI32NR/5OWG8GY1Sv/adbJa6pOs0jhHvmOWIageW
ND0+Sg2HzfO2levUwNGweh7MncLfL8kCrjHhtCDpGwqLin4RlzTR3Q6W6ei5860t
OxAMwSscJeZIgII6Su7I8aKmVQY+LfBjd1BP5cZ3lr5pqWpzQkdHUTR/roZ0ZlLc
NYb5g1yvKOJgnsTcpUgcJUTJNCG1b6+NWGhzpsP1r1PsQnPZYBIHTqoHQ2NS94Ni
hm7ha5rExm/3bcJG/eMRLWxhTuJEoGzc1InmGKXrpNKUO6HdHVQlAHjca6YgFVbb
b7DV9dELtSEcKftgQufPlKI0BM4GQ87FiP4UXHpTEd7/7y8EIagkMxE4UXs/aT4K
3kCkvGC/fSGl+Rwzdw4pBVFfphfLKObcP2zjkaO7j9v27fR4oPoPUs8mjWt71cTH
az4F8S3XH0KTlU9P/T3ysvah6OXyX8JI05+YskwBx6G46f8Ui2vZlmVkw86Vw5SQ
rf/lvmtajNciEm73rN1B/IhePLH3T2SSwV6vsnLUrkpsjqbGx0vr6mgLNlciRM/C
S1GSHdOj7c9q9jG36UCpoxuW0Oe8NkWojw6OsC7/+hxsRDaohgU7z0m9M4Vl5iph
bC/jLGsFqyQIag7ZR7L61NB+dSpHfDhRTz/iF6aeG9TkmbXHvUohsiXwtZ3RfOpi
+CSXc4Ual2UB8Cwdu1DHvUfjx0yI6vYYiabpiYYylE+S3NLbv6Z/2DFcq++0OELd
G2J1qsSnrT+kl68XXVOR1SaAUenaXnpBPqv5SbCqEJytkiwHXaKp4cAQdcvlTki6
dua9U3SXb0Nb6m9tFpnjFh3R+Xqd6QOY58WD+jbrgZ+BlBjY32NZfa0KJikwK3eI
bwQ+8fwDyuFhRpwTGNsH51d3OqSHjHHX5OtJXAQ5gMuJ6I7pDBc5mQsz9vKidQVT
67mQ654F3worCHVKFD396g1qwqpzG/djDPq25woECba9B6cl/SKGmzTXSM+w92A7
etq7nHQFVyK0TaqluTPRgz5Qg2a9Zd0aCWAQktpqljTzGnEysfRViZmeC5BO3QYk
3OBm05xeSH52iCJDXywqcd0EgsAwUh9o0Kg/Ws6wQVPldSx/XlYTAAKMPOujm5Df
7c/PEX7ehcVKGKEdPM8g2Y912Dw1xwW1IVvt1QpM+vzUpl2Q1IfI9VILoG3S49P3
SMo/u/ismx4mS7tcuOF2WhYH87JTBv2YCRlm3dU78rkNE2SnvuheWv7EQPzsLQ5j
iwyZlTB+2llzSUXu3IV9at1Ht+CzLawkeYUBcIid5nz8PutM/d6W3cfVouWindoF
Ukw3URP111iOhy1tnDvlqMme814NpDtttK3b4K4+32nIQoIWT+4SKXMD6Wd+aIIq
6zt6iDAA+Qa2ANcYJrEEEhgj9QPobEYcswXJv3JOFtWyESxIusVxBWYmoN3VaWUY
8FWY3TZplCihLAp+FaHynkGdzZfhk+qrjr28RZgyc+ZfWzKUgBbQrDSXeXkEL6Tf
4FKUtMoX5iTS7SH5AeMueWgHqh6EYz+4SCYARveUkZAPKatRQpoJI4TrQ1hLZHk4
thheWbn+hB1fKB3eYq1ryQRlTz1APV7BNbq3QMz1pS3exhIjoUyJcPrA3CTOv5ip
6inZA2bpQKGE+CdDcepf8R28JJ6pNvo+Y1lzoFVg3eKe4gdGX2PWBmj4wbS+QIh4
UdzOg/NTbloQuQQvWI+A4AwWWxUUwcS0VlkjXmEWKXqI1ExK3ZmmMIA66A7vIoBm
274U+Gw3EbwUyeM9uPlEOW4UoQ/C1Q73xasNhd8D2pODxWkXRfi/TZZKXrrciMiz
p5i7fwx1oYnIyuIHDTdlEYIj6mTU3EFDGNHcsKRYwgMR4kOfl86p2+TDywkFB5G4
7oY+rByNa7SHwusWKE378zDqJjC6mnmmLL1VlJt0pm+ZY+PRdRz/0FsNRgrCwXiO
qwzPBznDQrzCxhB3CqYG19Id8es5vPDM7TsdycXhjQXtFHQ2XESIq7Vpu7inJRda
n361qWrziX+DYlt+PZLrxYCpvRPI2swhMyRjAfv/TMwlwgBH7WN4ZLZF3YC1GL8J
qA56w8Cvit5pGLomKkrYpv0j4Ym80nunkCpex6afVduMDqdmd72KexNbUV5CI+CI
8d/WSwupKu/mYu6Q6qeBVZasKyJbfO7SlBYk90gFP8RawJCjuqG4WWL7Ttv/Bm5S
ZOCAxD+uuo+R9+Ptt3WFOT3i8U8LcSAqr4lMPJbe+x3XiPgwRWccvsSXMgo/FuaK
UrCX/teAZL/WUo+oKDWSXQqwMJfFsg0TgkI97D07suDV3Y+5RYeBOGNEtXClo7cf
STInllTzY+4s1Jz/raYh/t5LwEM/6tz5+LrJr8OKTdyu4GKew5ciVpA/2F/8LCUO
DjKl8sf+9jPcZepoK7cfPmGGPBXHiKn6PfQ4942ofZSyhB/h+N0WvZHa/eK8yazI
A9xWpe/cBNg1Djd0r0y8jCo1eklwctyavBH6gCZbb95Qb1+SDJOrHgZWc4zGhHfj
vwkQaWdrYHDpu3yj9ZXgcTeYeC4NzXLjXqaQ5w+7PKdkhDzCqBz6kA3Cakbp220H
KtoA+GLx4YNjoO5fr8p2EsvLB3SrrHwBkChsYjrTtjTyrPt5QzGYLnxIPuRRxXsa
ge8qBEP1jdvYyX231k4XcxSfaaONxUtl/btIRC4RRi+TMWwHji1bt2NrIOQqx6lB
JPz3tsnTqdunmHa09RppiM5bJ5Qh70Flsnk2ZxbGd9SeRr3tAJfk44sc7T2MDGFU
PUxGqQJ3QTMZhuTfjFBcJxhGRgK+ERxNv+NA8q0S22C0h4gRC4aowJX3fvVh84nc
ngLXNSWNcCFAOKkdRJcJa2YoEFv9fyEjiIDE45Y1sDmdKXTkb9V0bflQQaP2en/E
jLwr3LIGeKI0MzCxVVwIHx97v/dny32+2ax9CdRuU7Joi5BEqGwCA2mLm6cTa6C3
WdorreYByYQs3afbjOQdVNZZ46Sy2QyAoqO40UPT+ycsiagOYyGM2UbNck2vlfe5
+xUuVLD1jxbcroNlHvwgGxQjWeQZ2EnINuilu0YWwYfo8X0MZPAYPgRCcLJ5HVzv
izsuHPEr4ulnVrNk/SH7JCgNhJV0Cpaw1oIKkN7PiTWCbq9conFi54cijtA2s6Cn
KMc8JK0qFtCF4kXJO3uU+3lBlk9JeFLXcMvEnzI1XK87XoCdjKBwsx3bZXCzDObv
aDsXamr95YLiqqEbKyPV4I7vCA7iVAkWxq7EBqnJjHJkaAqSX0aDiyEpb2pnqPxu
ndJTqj9Lo7NSxIGuGOR+JvRMt6CeZFlKA63IqhCbiDIDkBlmJTo3j7sQODe2o1aR
nhsXjSJA1lB8FjQAgjsCp5vhGDWwQ1FWqGiMoZq+/FDHSmrRc6Yg2aQkMa+NRnoa
Ty9Mv2AZ8brqE1nN6m5RMI8uusW1edsq9KgzNzPVCbVFuua6AlK2P0NduiGQj/Ou
SdylAxXIVbG7g3OJtAU3dqEwKIliLgDCb0GETUeh6UVqHnC8cqA9C1/9KYpI9Zkq
0v8/9kWlIbvZB1zIs/J0H8q+i23kAX4wKTQbqMTlgtP9CO0Nlo6tyhxLlwBRmvYD
U10A2workEG4F4Dow5JXncSrReE2YpBi0LHgFO5912v13sCVza96UvBakJKZsOT4
lfAk9u8Va1HyefkCaUsnGxEyEzGvjxy6zvrdQaOm3nDX36TWwqaTeTe52LP+9KPz
0XnBDWAVq54VnGPFFYQqDYcCEsEa9HSLUPob3/6gO7mKBCzTuV2rmZ0GBwusmbZq
K7zyODi2Ecm4+dLCsZVWCe0B6RylPynY26rGhVlZiO8lhXtM931IQxx0IEN8zmdC
0My3cppPh819E/Qd4Wt9xTvh69tDTP8lHsGWW7HWQNrMMqPCqYgrCU5ChzeMhg8c
JZ8HnMiXb/CMqHj59/5W52DLd2AWMbDVad3E5CjZvzHxhHG0eg4Gl3eRLoCbNXkA
4iw0MP5UsZSB1zmvs3NN8sgDptJI0mVShlTE7vxb6TkV4MxIemKdKzhClLroRs3C
eND7QOC7eLCAb2dvwSunbnP+aJ7joLG9FSMpyvwVgpk5bwKML+vve0EkL4HtM6SI
21VFThEzqLmuKmEKpzEKfv/EVfSUxJIbtm5KwtgP+vnQ9AnlsVuCVGGxIrJQhP61
J8AFghY+8cPypVcn09d2igvM7dKh4PyiT2OG8uv8ov0TpUShk0aCKij7VgcUGGCT
BLlnro6JZh3LNLxH6xPSct2JgulwoZKQ6CfF+vYS3UDAljGSRtfTK/6jtX9PP2qk
iZTLJe8yjmM1Jcv5eXoYwKDlTG6Zgbd737BzBu0z1E1Zalg3askCxKTvSR6vYTST
fMZLyqQH3zjDu6FbLgsIcn19mI7W3VtYVeR7WC9KQnjSLl2AUFRWW5Y0DuG99Uzu
VTi3pm8c8p1NFbJRTIqf/QJXwHkdUfdKHBuPmHuhbS5iwidWWAprgHCC5JRZp1Hb
VvD2GUE6SyFuIKRrx6z79eEVcMaaqTqiIPz9wyBLtjfEFgLESYkctJiyEA8t0Bgf
oRuXhtA2uSmMg1pCJUZMHs5LgTEgPtIXotRTI0PKwyI1OF36euC8Gyh6SThChuR4
wHfnZFa7rmKffF2HWpMDuLKzADnp/LADYjShNmMTLjEFGQCIRFbbH63Sh/uT53y2
8OG90AIFTSGjWsdNDYN62htUXQlq4pBAqd/Bn1EtSU7khbT/fhkDagLge9OlYRUD
WxIZXm3XqlU7cL5ehBlfrQ/DuGa7BCEaX+n4JEjv+bWWEM99uIq93PjAoJUU9sVM
mU9//qS/vrNMZUgWVPQ9O+Nh6k9xSLRXV7YkpgXqzm4sL+1jP7hRt4CY+lvEUVkJ
ajY443QeB6ijY5z0gvlFpSVJs7emt/4nkCWVouL2tVW+buZzc7WJn5G4b/mC3Td/
y8sI/lJUAGAAbNG4znxI0eBY2wX3twsgGVKilLg1cVwrt29bhMi5nDakDXrD/Jwd
DLlz8AVr7FX7wAZmLj2ZRb6CZHG0yt0Y9RdvJxcgfXdsLkVLdislvWSxzf6ve1E1
vf1ysPetQcnXKMkpMGIHxyHA4wCyrIYro/t4tBcQ169HMSMaeA1bT6RWLwJaPMBY
AlBLncsUBMev0i1tKmj/62EOn1NudYbKiSZCePRkvLi/Wpmshd2CH47EpaxXmfQI
1CVCPws6hpOk8HsENVhNRLPxq4R6CYklpLCE014VdyWsI5YZ4BYh52iuGzI7bW4d
gMrJrMz+PlOjSHveVZijB9zaXoma+s+Mrf5j6FuivFDbSFdjifQAkZi/sMz46Fj3
a/UCZNu7kCG1aZfF28PmhR5kWPbax4jXIRrhy1125H9MeEhea5KvIzj2SdM36j8f
zXKLJBiMUsgmdpimxQScX1Bj8axkgSBb88/n3Ddqd0MRNcHw4ZtSeP7hNJ6/m5nX
TEiG18FOeih7bmSED/JseGCfrX0S/1fCo+/kVdjCZZy4RxOsw92NSc4DvxjbCtp5
UU0PVHjWOqx/KFOt1IwQ6oalezy1Mls5vmB6A2iQFzxbseWT2F+1z1A5LPhDVCa+
XZ6FAq/b2WJoyPZt/2/CTmx1bHCyGVKo8+VvJ7j3oF1aW7OGIzRLIqGGnmF96hSs
JhWXff+5IPOBAWVDxPORgU+TPPuIKbrkUalygYpd7GiBNmUbM6XbTzV7G79lNk/3
i8rtc5JykGTR12yqUR9sXnmrHv1Bk1HRxOy0xOJnaWAbQ5bVIlYFfaHbGI04P6mT
igym1/p3TBmh4+Gl4kDSuA5kVuCxLHhfYhdJIBd0uxVB+QRcUySf9VmZMUiHtrRx
esFttK1vbGMU9fXI5IQHHAPfrcRi5BvGe/t/Wyq2ySli1q3Pq4qw96mFcPGk0x+g
qydXFh7Q3zduV2gNxg88ALZSwwPS8qjbeJ8PkqLNSlDMpdlUE9EFpO6w7ccZbItf
rK7hvLxnJc4hynf7OYh2mAZvWHPA+eD458uabLQp9FxCBWgrN+691Nl/yoNnhINw
X1MLw6FzmhI0GEFs+aM2Y7m730cRohOVY5J3MhFcF2Ymv5RPrJCUFA0jz4HUh4eo
mmlI1WR+SR54lW8+wCQzJqCr2g9wjNaNcleGmqZiZQiIK9pW2nPc/9clzTYE9Jw5
zGCdjNBkZ4sVhU2qeL5l7fr812yO4q5E4jzN+dERbeUgHBmlimEHbSdUkp0cc+vt
yHQA8VVH3lWth9pAL9HTCO2y60naXdimotm0soOwGQYb9HjhMT8lXqnmecDS43sb
0PtEZ3kQPJgKNGzbSNptUOJxadD20KOz/BWilhpg8OtL2IGQhl8iUR5DNKnzbBax
o3lMXw45kRUz3A5vEOdaTgqLHOJbWqZnzX5R/hIeUY4bxPNWMyAoVKkA3SxBIwLF
VFnPLTsi7YvTDp4TMB59Gm0YICqhGp3nfjpQSQcgdhckCA7LgOifuzJTHU8Igu0/
QOMELZLYBbzuKxhTRH6vfHZ+mqi5CoLp+LTIke9Z3GYq5+YlgGAgGUlSjnqrpOBy
+KvM8a5LbIeABty/yGAteP4/zXl2IfZvaAT4LWhsjXRGFrhfqFWVfBfQYwr/dyCN
zJvsIcppnmEiMQKkYrw7x3/VZOhW/lPgRv9JHo4usxQz4w/9xZcH3YzFHrrarQGX
EyWoeQh2YAXo38CxFI4EL2fBp7XMQ+J4xmzQFegZgHts7CnRyzUjmUQ++xMStzzP
PLMr19cXn92nVm3x1vgFRN8BGji2VDH3a/Y9XwCgwEoBD3A1WiALPgBCQAMcJ15+
FYeA1bgK3nr1ybn3aa0Q9BXHZ6evXZFyuh2DcatHDTA/kV8RwEssuxFId/xFvoxH
+gJO+xx1hyIhylJmMdAJC1M2XKj53BpccHP1rENvTKwHwi/Ve/TxY5V0+IivZ1NV
cmbOMHx4pSmSbHHxZeYDpblKQiah11hanM0QIV62ULXXWga60afu1A88EUPWP9pz
ooevAUIp/aWnlACBo64K2EyQDU75TBH8odybtHwXUUZtNDO+fs7L95SxLCBMXW71
QQg+LL4HFOCDS52cHYPnAh5jNgfGBFZAIDDgy7HODFaZ2gOuNqefohAgaXGeYnPz
UGyqp8JAdB8AjAu6gR4W2GaIrbb8kubVsxVkCEi1NOVR2F3O/q/01Z9A5r8FCOsy
bblI6+n2D38KBw+VH3SbxodLrNrgd+mb93KCYypU1/2ZZhGc5TdbUPzZ6PzhEjYK
riz1Xalrp9Ksab/WNOPM0OwYlJTjPsyCG5IQjOO0O/GgOvLIlX/EOyZiKSaz5Arg
m7v+Yoa1jfbc8bKeKBNmj1eVe9h6l35oxMtj+mSOkqprY5l7x+vS6yK/KSKC1ouo
lE4yQiG/LHS2PscMeFy0HRK4qYw/X6OJ0rbwD5RV+Uhn1cRM9Cu7bcCEDe+pv/da
+N2uhwmLzlR+4wEN2nKnJMidHwatX7dO+iDsaT6mqteXkAryV1HiWSZUYgz2lk1G
mj0S2vN+PAkKZ+YOjynsDcw8+uK2uTwmLJ4ej6kdCMK4ybBYOixmiyKWDU+OW82n
0JUlob6wJgmL7eErPVvXuhBW2yfoBCHBtLTghPvnfR79+S184JDKtGox9BF0xY5l
GrK2GZdGcxi/3ybYPxueXakmwHXmBNqb3T047ZXRJZveLgAvhrC74Gn1ypFrfrff
bT5bBPLSqfIKDb9kn7KNC0rPRDQh+f+n07XEljfKcfB6+nF7ynsbVaqk/ILdVL9S
j518RCGKqT3sgEdpfSeigAPpYh7JDxtXxWId3py0+Nu+VbpOxBLZ9P/sGUiKXX11
M/4FsSZeuSGHIV9PBQzzKZleTDzgf1h8xvmaQr8hzbGsh44mVg54jVpVEScK47xc
OJDKqEcOIKoqcNy3/WHk8wRGVWMJWE0DHgRYUgj+KS1okCVO7F/yVnfifiqwJnPn
V/j1EFe62fC1IcZt+ETBxJlUOV1Sfw26a3RM8ej97TIaOj7knusF71U9yuaLwIpS
1p7CcOrvI3S8D0c8xSS4T7jI396g2+RpeKmfxRdat/IUmLiHlsg/aNEWZanUrqSN
PjgXHr2HyEkCSzsQ0pGuIwEVC5EhoozQN7iQEotYOh9sLNT0/diEYvNwDaejkGq1
fZUSSXIoM6HL7mc3h5MpMAsrO4cHnBdRphrcfjTH7kaM35unOwnsq+3J/P8Uiqik
BSiG4RZyozoS9L5U/NN67i/qbsu6ZDaWAEAsMeY9THQDd5eK9jfRKphlvQaaliP0
6U0g772nfyXYOKPjn1glPmDENK1o56BQeuDU8qbTBjU/m/U5llrpmtIZsmW9RoBg
ArQbJcnEG3knxMWR/SgTAiT5J6ycVQormBbS2vbqqXUhJURNyUu1I2yCoGYZv55g
IadjwZCawYVNngCke5/OI2OzsFzYBVU8NQSQHx+6MCRwaYbAVh4OtRqN5vtoGUVY
qwjn40eoWE2JHu4ezOp8FR6rxuts8N+vjqd1q7iN1yihzfYmkch3c1OfoGDtdAo1
Wc4CY5GOkoxuIuR4O80gYSg5+phPWgUJWnDA4ECBnj+muBDrrBilSoVIREwZmI9m
dqVqFCguXsohbRLKrv72jGjJCoDFvljKQCUBdGWkxVgERB/f6W4R7rHpBtFZsum1
N96N3KuBFicJLP8PJwI5E0YCI2aZNwkgTpSBu9C4TXVKMpqIDJQc8P1jJN1Wr81s
7G+6HBkpaqXjKag7pKbHHoN09cvBkLhx16cAFxbLKYR8681iEbjb/Ya9hiBBgZr2
y7KsMOQHw9I7iH9g4PVJKyd8brdGWmHmFzuKeWSZLzaa+rljJ0tmj23h04n3KdGb
wIcYja3SsfIX1M7+bVk1k23hOhVbwWOjzUrTxvQ2nOeGcY+PBZFhHzk9KMUngN4S
TlJqEujSRU6dIPg4XvlliOyP78z5AayUxaE7FmDbX7/rqUcAwc8Gu7eHET5DKjxH
66+ZvKmzYSQ88RYlPXZXhh4t51wyQzGv5+Qnn5bTNIYAPJwKfOYBDWFSeCLZKwdF
C57YBvNyz9FEs++GZ/KltodYipEaxG/fxR0E5zBQ/jdmCdjBykjazGz+nJxqsOSx
PjPoXi3bSmZzbIWJ2zZAgt59AWPaD9RB5ao3qGvg+d+ftpHLji0gnvs/ot76eygR
vu3FgWe3AWY+Cpul7FljUgJbG249B9wmz7BKX94/RTawJIs+HqPviNJpbpwvIBGZ
C+C9X8jlo0hioUGkehheVp0f/4/H/g7YnAU8R1FyClPPxXVsF+lE6Q/kiKTh9OTP
m1EStx98yGlqNGM+80oCcBftb6CnzjPC5CAqXAvQ1aa0QzmtQUSOlwgJUW3B2zto
eSe0gMOOGe1w7JUZr/La34v0an/6Q7J+y8h0/nCSMOg2dURQQt75/wIlMFxexXDR
5Kyto6mMqGeq7CeEg/zOR1/tS2nXtwZBkcxU/+csVWDYLP2Tic4fItwfXVr3hyeM
x9SjAV06HAOS2K81HM5nDTpaWfac8pZcG1njX0odGmSO8VY0TecOpDoRnXstx5ow
I+aKngNlRPu5pxeAy+munWd3Gi6pSfHjMZDOA6VMOciaUCmANvHjv2/qFnZMadMb
P//RlQJl4oU1/fBgO6oT6ZzZzmsALfRXNU20xrBGhIis4k39M+d2QLsuUCunS4QO
9HCSitVpegd8U3CgN1yALJYOtuqa7FZc1OOCwvKu3mx7rcwFBN88cvuVMcHgTL2g
UWQ62GleER0pcctOQPfv+ryKZATxJ2djKusKyb6AOMC9jtqlE+EtpLS4QMkacqh6
A1e2hlyMo96RwUeVr1uXVrKR3Tyiy6gADbKNiy8DicjeiGvd/heuIwEk6Nu9jNG+
bL/z+NT9omYgsj0Ma6fNnHlMdU7XOcfZImAN0qoLDKJJ/X4V+9xJXyRrMnSyt+dF
LUsJY6LUck7Ke9lih28hjOUXIH9opRxZOVjj47b1YzcKE1bSll+CRXjCEMVciVRl
z9CdiT2xI8MCY7MgR8XfxsxmLNq9DucQaN8uvb7R13PwpjOh7L+lY6dElzW2/4EV
Hy/SkFFOnFrlv/Fajpup74hvz6L33pAtsk9zeNfx+X9cB9vCO0JqwDMu7oRuyIFS
oB1EZH4g1KgzeQrUVWBCDBSYZpOxvRLTGLuKUvkUKCCJEBZESWO6i8MYuT2fS8qz
4vJbBm/nCrtyTmJdnpY+BoAxDqqBDTXRx2EWZ0W8pB8zF1nAB5+Xu1GOLt6hdV/m
Qx21ayXDw5iyPoisVRHH80Zwbj6iDkF5dhq938hE1TIPuqbSX293WgR1xrpxeeiM
Wx+QZHqMAM1twuOxSUM0OA3yeq5dU9xBk815JtXeYOTO7KFzXy5ZfoMKaEpwOzTP
ya6AhIrJZnvlug4cgDUGfHh2tkYZtAGOpeironqfaodVt/jRBcoP921xJwnFkiSS
M9nbmNTradfDLmm/UbyjjCZFRyTYseFbrOPO4Sy6jfNsOtoumALYuxOYSixj5Mns
VADNf7O+AWCb56eb2wA+/CeFrKX2ELIyV2fmf626rvOI1bwnebzm+yUum2jAWVgq
OrS9RWlW6eqSZHcDZBLq44W5CRI1Zp5+qwJ+cwrk8RyGiLCcyNXfGa+ccz9+LvUg
+1t+SBYnC2Rz6aPkXHJBjLwUT/rkHbvhCqypplV8OF3Ax9I7RTEWWYJQJR1BWDY7
bb2DRJWHc1Jgyc3uPHtEcirt0nnBoABOG8xrfU1IxvIj+zeTxVWE6XYXuEGQQKgP
jiz0l9sCnkCkOoys9EZM0jmuIKk/WTUlEaIuAMJSPz9QXBtnTkJtOPpLomHoQrJM
R0J5M85b9s8irU1bAM4aQd44NnY0gSZEzQfugADtlTWK94gZIEitfP/3EfbDs6a8
F6NzeRM13r0JbPl+Z6LOZ615hu6RFSQMQGK8U2udbWmpGsK8/ZeRe9gnme+qv9sR
douAe/v33sruwVqVDb1yHMYTUk2MC7bybDBapMPz+SaubpomsISe4HxuAde9FhxK
J6zHhKZY07cV9alqO19/mThUvpsljVlNStpjHrNBjSe4ncb+p3dh1HVdUiACMitl
X4WXl2fdJ5SCSuJFwn6D9Bu+GZbNCzP5IgYvr16HEoPLZBZJgaIAk/tgjd12kgEO
nOBZGY3hESrGlCdHA8iGYECukxU1cDPArkeoDLBmhyw1VWE3nc7biwysHE3Yfd3p
CmlmD8vDTA+e3zckQYpRWajhqtpZTiagbhr4C3RNoYI6KqyYiJFiq3XRPe5PIH0p
dRYqUqkyL46oJ8pmdKkNyvEgaCgtxXoB1/0jIuWzxDdCQTmvuhDIKNrJhnqlHiLl
uFCkSBKCUsVv8+KQSj3Swn46g0MkXRAc0B4a0o4ksYFxxGWbqTA+m96SG5FfuwFb
qLMP/+EhXdF0urt+J1Eym8pF3TEhNPQnGaVlMN+s0iUk8t0qgDoOrmF1A4h77tHd
YB1fG0g+zjWfw8iFdqYKz+Hho5C2ZwnMs/6d1OyACnkNgIV2evV+jS8c5tyLsUHH
J2GuB6DSMomtEeZ5R9AoMJG531f0PWvY13e6Oa75+rbbrUoTc5oinFUO159v/6jG
DoEp+GvuLm9x2V0Ith923//JXeh+XiQ7q6DdtaoOtDh7UKsfh9PbOfuURdkwiE74
gdHG9nzclKgtKU8LxuhpGSk0+zEmBWQZP1I0WiIbc20BlwIIiFZMUqAeXavT3kZP
VO/oljGwBCWcEAe0SsqYTEY1bGOTdcUZTVdYlgB/5EWSdmvDhSBiL9jelRPM6xXB
nHZvATkP6a3uN3NchuJvsqWUuJkbLSEYu6BtgZE2FFwqRDy4J+eh/cfl9hSga4yZ
UgxbA8kZ+nV54MSl5l/hk466Y/LEfIZAHOktpm7fRfXx+Vt3A4rF1HZund+RGQVW
ocb41iOpGMqvOmf3jH1oj5D47GqGTF2OWCQMNtIutbZzrOUEi+mCWFVfz5HGgjhC
q0FBU6jtVIVTWqQFtEB46MpLt+jDdc3QHb1qk6d4CY75waU2WOhfJtmHQI7oMczJ
Bd0m1LSF+3lU056KR5W4daCHymebJHjpEmspx2EX0Re0roQ1J7j2LGbKh7uOYcfE
2uSxqCrgNdmlT30gvqCBLC9R/XhkYCuefiCuCuTVThH2S993pt5U6fmvvN40ymea
51i96QTuUBTu+jSKOwNu5EBZ0GJO+0f9Iw8tfsPIR44VcKm3Ug8VirE9ZeT8F84D
f1FYvSITnmV38Eo1zAF58WDPnrzenRLzxPEPcPs8nZuZXT1yVn6TrnqJUzOv2Kxj
8dlT1XOKnYs+TSIcUd+nvtkgqMFrd6OO5vg1H0ec6un9n+H3TeNGj9MtK5zXiXMl
1OGU5YLNn4H8MOouLuCHfs9wFL0E7aSMBUzGPnYnTbG7ymfTk4IYW/ERQl8hzc+7
03Vt6+3Ux0tEDY8QzcVMdxMnQwJVIMMGvEYhAA9H2g3E+Xy+7F4rG/4oSHGrw3fT
PeXdzkkIDULiddao7tfW6rOzJYCBRGWFpJGLOFwR3AlaC68a+ilU1jmrdoJYlpOP
r4wqB4paesZXpLyXEroZx3iQfktxlcEUUZQ0d3sfVGWLQTaZY6sSHTJPtUC3jeow
jolgQ4wJ4GqcpSpoRyxH11TbLtp5i90dKSPlq8ZixCL6Y5U/ImuMm49Lvef334Ja
A61NDTO4SJHGXoxs1zEqrMW19aWYt4PhQcnNggYXOV6DHLVDNkvKpKx230taqEbU
Tl/4+IPSqDqoFw2yZU+vhraBlxzGbsxdVXWKJ3xM+oAJFRTAWlmy0+fwaZzXo36h
wrFjtsp9KicbX+hXVLHjl4firBbSC13AcbKgSBAxqMjUFlItu4iLM/3qZ5zzIgAN
azBrFY6OJLh4FBME5Jv5mhFibGQDJI6eL8GkySibGuQhI0Hl7NVKFkMaRybkCzWC
RfXG07l1WJH3GsPBy/Gt94Xt1JboMjrs+PoiedLU/zTXpCHVtxKkIGFWd5fLqme0
aLcUdS5BCIaNOzAofnP5M0pFFFltV0ZyLICqzAxP25Hj9n1q7PZJeJlOBKbABLgu
YYLDCK7n/vXoDEJkhZbT10E5zCro47x4dveaCZH8MlfOeh39SuIjurn4esp9dx2A
EwCWm6v1fk6HWQSZlUzjIIDyqOMlWqfyjyEfPEL20e+ugGkrZFg/cEvMGekxycOn
Tz4POD7zlYjA7g1u2ZXCLy1rQLFMRd0vKXberPZrZCOrU4Z0xZ5Oi2YNrboQ551U
jI9UdUVi0W4QwYWFq/fXgoyQYhSXmq9trZxFAfBXfth00IsU3ozLKtuCUpN6VJHR
eZevI932V9XpmN7MrsJdDsqxHIzJ/yo1Zvg1VY2FS2S/UFRjxKA28Xfs6ZgHlWBF
djuus0T7TuHZpnNgE+48kyBZaL4+iUJh772UsvftsZd0EnMMWvtb1wTYVF9Uz5qw
eFmA22ZBl0RusFKDXJfeNMJMs0qqrH5EIckBXOBo6cLHrMJTMr5bI2xh4/B1kZ0k
NuzzKpXOi2U4j4D3MfixTdKUOvDM28paDas5F4WQZ5zZru0MCRDjPVsBTnXUftzK
IDiswvDCLM5Ij0Uu6mUQqZgeXgG39tcGHpzssikpZgFZ8WvZiSRCOKDsToNuobCY
E0IUYtyt6JDjB72lw0XeAdaTwTMpGj45Yw9XPmo1y+drsY3TOoPiROgBZ7oGlcYu
gKSTHOMbuLL2kQQiG3wuf6sXxqL+SbKhXbLiSbPM+Yj8L/ZjSeJCATHj7qkrzlFu
LT0DUuxnO7hAgnMMVV8rPlicvbEE352vRo3jjAzX0G57BFJsV164dk22Hb3ykCsP
XFrDOtaUDvHbmmnlu5Q7tOKKJ6VKYeFC9uC5l/j6jQ7PbF+li8WqGMjqv0oey7OH
d2u9R5C7Pu3cWYlLsdZarKS1MICJ+9fZhu5pyqFXCQFpZp1ILOPAg9sO5xsefMhZ
QqA0QbrtUdqYMHC0cAg2PO/WNo8kjH5pEM4RT/0msAUZz2mahX/+5xn3iBgGWL4N
BaDR3uGcCFWPMGziCQA25VzhpzxSqi+62ttHUehvXtaQ2qI9oMBIIZ5kFwiJxiQ/
5986vRRAV23Lib30zmZ0YwN4xx1SKyRhTTt1nXo1wc5s/i2xNjm7DMsdKNys3hbs
s49J3ZhFCC0UCEGG+p7rJvo0p4B3XsWUh9R1rAjdjZwChx8bJnr5nrvgeizoHIu6
1uJ1/YfJU/1Dy+05hBMVzDbjgWdb4hADFyIxmmLlMOSe+PnrG29VwW1wVAVg4CDL
lxAyv2Gn1eCe+XdUSVqq3tJU0CDJYhY32nWILBr+6ECC680ZqfdaTtOjKlXRWYIs
vdw9CHNpOd7mTRWazuDw3SsdsdH6PtsM4YlvxnjqhJMGw9bTUUtb246VRnK3QaXL
pZAZpQpdhUV4bDRpR438mpvxF+ASIHqrB6TdiUYYQeLUuG6rYJSJCZ7dI9jF273b
K8BjoYM6v5mRjyhtrIqgZtXoS3oFxwjw8ypfF/FDfJhf/zHA3IOHmU4m8MG6HPaX
AiU45QY1v0ZD9KmuSjVmeEYzHGdkvrGIU5rsBE0Sgi6YayAAClKygrXhBuG4eTOm
FHi1LrisusX/pA0JpbLJPS04rt79S72F4u7J+xzOA+Q5M7/S5lvXdbO0KS844UQd
7/A6zXx3uOwiTsKHKe0cV7cblcnpNlF0OX0OlwDfv8MoF4u0gEHmFduQAXIRJgqz
EtO+0JmpdpwrCtgPS6uqgOvrTiJKfHgLX7jQAI/1fPMNELL5uVwsV0VtmZ3VfqIh
A17Z4a0ZxI8hKJgmolShUy5yqzf6+r8PURawPRbPPreMh5vjy7WjQ4Av3hxmvKkP
pr2d1KOQgpnw1WvCqxWS7+tIRnjA8Uysusk1qfPJQScvgBERlXbgD41atl4DKznR
A1jzAhBwfDlMvBzP3lcmFim2TQpQDd95rv1UrC3qzcCNtkQTOPailr01IdDgine4
Sn1EhsZiawzupJPHPiUCAoqLpwsO+BPWZi5fFHqvSoq2XnyAg9oXYiUr8jB9BJML
G1JaH+LumkPcBHQjphhcsVOu5tHZ59W+U+OgNz82AXHJxgb6jXnDrmfWxIDhV7Hq
gIvIXHirWqAePjV1C5rXweo73CMld3CtMseM4+p+IhMicVbM3s0grrJvTpzKk7BU
QmMy9wpaUH6EzhsPaTOV/r55ihERCMazSyB65Ffplwu10XABGrlfnKdQ3qbLGh3O
QXA5RbPuQsEng11I6Io+z2u8wvXwoxhREMbdgzJzlaSSARgmd+DiPjX/Gp++GffK
cS+tqqEePiqmXWh6JpnloKrzA5QuBwXR4nA/+VyihqDoL6ywV7f2YROHu4THFLLy
KxGlGGwk3uVWnvOV8nDpWE2jHdAovF0szAkaH+g6pojepMUz/b6PXPBCgZSQeTtQ
I5Y43Fue9siPZSMHi9zxPcQWIwq7ggQAXo0GJtkKQGK4eqspaRkdPTzx17iiys6m
AzHAzn7dQgB0zd8QrzQj6OT6MhO6LtAJ+WOn+Q0eit72GXlkMjmTR0PfqfPKeffq
TYLRAHGxg49eFrn0c8Mef+SIDHt876V19qL9jLrnFsGyZQ/Y/yyE7o/TO3PF+zJs
a3Hl61HUpPYEbWeqx7ZM9gbj/skmDHDlRuiGJgJ3ulwDmKk4mez/yhZFNCjrvU0G
bBqTSQ/vfwyUK/1nFWZHV/e5H4Uqe0bFUX5PfTagmX2gNNaCE+Y8oKOHl5Q18wwx
L0BoU3x6IqkdM4ZZmzIoJgjq09XpdewyVbgXkreaHHEUNBGsJ6d6E4BoSZDEpD6e
st5tYCTWmg5xJHlS8Ih8NMTXg8fTIlgVJoRnA0o9T9yEDvkhDFyeMFdDDzznU+rF
cLJ2B11czLIaUUX5lv3fC4ug2C2+oW+HAp1uXFmNtzHozFE1WRcRZUvSJdUN9ji4
EDOi8FGP+HEjohIjuoi3Z/zG2HmuxftHzvN2556MlsxN7um3C6vebKGW7SVo3I6H
eG4XafQN0fSAR0fG4MAWDQRFRnd1bznABA47H+02iaI78k5CR7HsAnaKgCC5zV/m
4zhl57aefk9cZGNkXvVh4Jn3hvBM1+WTJUN1zntdlq9e2x8RvDkNjdCxs+Fs3Wir
7M4MMeVfigRoWf34li8U2/L2vDsSrvIFNWRE33pG6v754gNxQih6kbzBrItefdm6
Hjg4b7xfTyaTgyvtoaj3mJRHxLJ6kKxPWlBiFq/sFR6Cnjwwl1ti/43cP/Uqslds
Hi+D/mRYQFZFSKv4cftmeqTrbo618JTENUKsMeZ+igS++djvC84LFH2m3zCJATDW
D41fySczIiz3zLOgJk1cOR0l5sD/G9qYozHNvyDoKMgbgSNoHuby3ASnnlv6kbut
tCs6SRYu3wrspdcTq1rRwMji5M94bsva5MNT4ZhHrDmFUyixitZaHezLbaGESb98
irCyzeTT0jx96DB7CFtgigmov27W7jIJjTsZzDdUssmXYNV6lzvcnZdHR4pWKeCv
xR3d12uqgbapzYUGnzoigvVtAJfA1oe7bIg/x1qhtjoGjJHhL0ISKk1Tcf+Q5KSp
FVZRN02be5yAaCQnReWGwE6ca8ltRIbAjiTi/X1lt2D96JuVKCWgVGg4fQM+XSpf
X0rb0f2EQ4xVtr0FbCmOUg2H2xBwrQnuKz77BILMfREalpJEa+mWKaOLmmCCM3EK
gDqJJDaneN0IkGDVO2FSXS0SvE20utRtKHEU0RWts6WN9PxI8cJxtHh5IgHs8UmS
hi9EJWg0kyjIxwelke0E6c0Y6JWQYY+r6wDHUiI380ds61dCsr1D2LRL+0t3PooH
/aCQoy4O/ulS79rUHZN6F0foZ6CVWHXsa5ku4DlGaU1fzAwLvhCv51Vpu5Snz7Yf
fbhPY3PxaJf7wjl657fCJFv1UgLvpG7D4SW7YvXPL2emTD0lR+AhCCTvExZYwdNt
YABOoqOvVWj4yAyAzCSiKH6kJ+6ozLpECMV/egcQQY0KnY41YLTYYYN17AQfUuwX
TI3YmJbLfN1xLUoe2yaYX9KwtCdPi3yAaV/rHgM4VvAJ+RbKr2hfnyJa/QZv1Anq
0xxuQ+MbMBJvrbcCKQ4NBKS3bOLfOxSSi50frrkHqCeFLn4dcKR+zL31Dh8qcx7Z
PCAxOz/83IDmTe++Z3+cB7DQYsrZt/bQeWGlNMn5EG3D6qlGDRihXKhcDDetwUBY
f/a8Qp7APv0g9qNL+x79Y/bavNJG1UlAee94JrBvj8wae04Z68jpYDeeGHbCm2jI
HMcVNY3tVQZR6l6eqV/ONXd/n35WaqoOuzVH1ABZBjiZnwIWU6ZbHq7GJ8rIFIGZ
P9Z0XR+EEIGRtDVnw2iR4oCcKyzX2u7fyDiOImdqn/IcV/5nhpW5dIi78bItjdr1
IFsU0Cd3TXbMzbua7o2YywW7n4w7ojgaH8mqOlvQl0EEkDiBQ9h9rY2EBq1X1ITa
jpMa77+5URaF1Q577mlTT1O2gMKhIKFXUfYLqst+ytZ9TBQNFojrIdcLsacurHyw
wVbpFavftzEBB/benAwVcwQ3tPSP+SaaAEk8B0GV7ZIR2ehWyGVUJbInlamIfl0K
h5B8yTa2wQT4nqnSkVnQfGB1T5IP51sd+SbPxZKEmS7nMzdR5Y2Sr2pLVQuV0C/8
DZnJp+fVqhhyA0i444+zhj7wkRmWE+/EbXXAlmEa0ST/lAPq504vHBiuwmrcv66k
BxVzFKGI0NMFBlt/yitvx2j38xyPEPOUs5os44yz+8UgBxny+i1oInoVnJp1tUHN
uv2Z4fF0kP07d3IL/vFGs3EPQg1UXYQ2I5r2g7175Rezxxo6Cj8IgB3atGDCIJTl
GDv1p17lfhCWUiCZ6fVAe7joQlp2/5+7Aaw2MXXczs+ZrbMF9mUQe6nutXxwrP5c
iSsuTpfxzxprTqtTcIJvzBfix5z44T5s+9lYnNEREo0BDlBFeTSD8yg4jE3JDGZu
quxbvREypaSjGlHnD0Le/eVHoyTCFj0FOMYlnEU5tDUF7EVPc67YXTt5pPCalvWr
MbvC391hhBWTkmJGNqdpTpfB3Az3SclNMkrJ631+lIjBErrATLf/W0M4a5T73kHW
rDPQwd3QMV7I94+cmfWZSkzlV4aEuRJEpWymsVHTVSMzWjFRYQ8L0uTagchXPoHt
bleEQAyQnhV+8Sg7DPboMTwPjH6Q8MzoVE9A8qYJgkRoKOjSIoZt+Hu9BEgS3xCc
NTOkClmvrtqnqMgdB8WSL1XSkRX/m4GqODWs9LQoL/ZxfOUdY2DOdYHaw4g9/1dv
gR06+CKFICQjnr0N5LpMxrTvmnf6KM5cJCPQKWp8Lu15dTMp9kQLfeepZ9pnK15t
WfxaOLV+BIoTbG9M+Yp9FPCuPDFIC4W+W+ZhIMjK1mrY8Ngh4PH/NlFbCk4wLOAE
B3RzWFQmBX7nfGOonwKUuENTF7oNnt8aV5MfasKhK/dlbc/k4jszQ71TyGdCghbu
BKcPKpJut/OyIOjrwfc37YF8kre9PJlWDpUnM13jEAFtwCc82vI/41w/cFWIOR5D
gBZd7I4Z/mFjbrkPLlFTgq/suKf89hhstKOrdVR3LbgeUpunuUvPbcN408QHuyci
iKzUQt70jqxBPsTZGT8FieaFsHLI2ZrH1i6HWEHKAICAHSr13tvtbulNO6GhUjSS
Fp29UUyCAMO14WzCwXMTu9w4Ud/haFMu81/j2El2w0XF1pByDSwjy9S4J34FDkih
2KN80FwuFrrKmeaF76KCUbCzcLqS2eOUb7ImlDmw31RMukQ7qg0k//LvzA0atXFZ
TnDz5T76SIBHb/AcYZ+OBPMv6jfvSHrCI3PXnhJ98nlaF5tDylib7MUoB3NO5B18
y8JlkWnKkv8ZfZCNwN333FTmkOjTZ3GiPGXlUUxNvCUZe/SpkN2JsZodgPIZmdfm
7cj1OEpFSIuDf3L+nhhJCovS0vWW5Frh3VEbRiA18XAbG/lDTI64oXKJE+ecNzsE
VjciF8U1BO7jk3rVAlYc9QDSPzrviR+iK9PySXku952BMK1E+y4rdK5dPGmrGdOP
cFAjrtk4330RqFmuqKY7lifjwMedPQyzOuP5eWLBE0lby/9seO8JpUAxRGuK5Z91
Zz4GF7c+PvgCjh+/QBQWDGJsMLvunOQiW67SMM6FEnLhrJQdVLwO06D5XKTnQ1ev
U+3qHWTv7hURbPrQ8OKqDgGetEaz6uKKC+/d2ayBxGAyoVETNoyLD7FEJu5xSq3k
sd8s8PCrEVlovbpc3uc4t5o5jzDIaShUfQEdUT/PgI8YoyBDFJSeKcIR3lw+Vbdy
mNnBjY4LaFEYtpMbuHubHa8Rfj2GNCJolGrf0dydGVaBn8N0I2HSfRSjmUHnaxaf
Ox08uxjx12qGw4QhGoZq59nLfaRNzoTF0Sd98tz7znPUQ/7pX/H7xZ+JikQFiJp/
nba7yVMTzHo7A90JZSPpBNzCC2UFHDWVwl8bAbWkayXfjfWf793pwkdAGRIik8Yk
ekchRWf1gTciehk1V9FApZokKxRKkrUfs/zfKRM7EeqyECsS/1b2OQD3X4P3WL78
V52ygNmtgpbrenSv3XuyFrWLdhULbJHui1NmIevbFd4Fpkhm8popURmHmsdAwPtz
y9RiCPKiruZfJGJAzWxgPz8DwQSljX+nH+adhnXelIcRjSnFMT2pDA1JWQCKiAw2
K5OHeHqi5/9X6AiIySDGRtVM56ayrqPdjVFEPBRBdBCLGDG/MkaNYvD1S2wAczxl
xW07pW9gCDBarBvzqbl9HO4akniZ1ujX1NSHxIAVhtHPOqlUwTgfQPrP5vyT7lOJ
cVjFBGPMCZgMJOS3Q/uiYOWct3us+nZ+P2Xvd6yXgPcrvRi4P5VmufuMaf0J7X/B
XhfBwmzjBw58X7G4N2KVpfHkS3qiyxLYjYa6xS5Qa5ndtWdviIBQns1cUPQn8iz3
hbz/DQx7RkbR6Q6pYj1KLO1PPfro1f8eVJB405HPkgKKBnXpmHbqJz2uhvJzhFEM
QDif6/Px/1atjhI9yqCEMqFoPhIyJXVfdNUNzGp4MjoggKmB4EjRGRipHtSNGlQ6
pkSq0aaLjq2L1woCc5jBff9BUVKWxib49Pp4oIF5JuGEfLQz2LciwwDL3gLg5+m9
E/mDNExvjJXQrqqvAzvNXvfpWy6eiPczxjhkvi3swincIUV/jCGmKMSxQ2Kby2mf
81aXIOiY8zPdgmTVpjYyq1XssiuScxbPreg0X74wBSp0CCpVVNEly7VZVdy0VJUH
WJoEJHkLdNCEeFZSlpuN1hHLbi0gOFSHYQXQvFkPZZNzZoAbd1Hff2GlHnHPm39x
Oo0/A9fvs0i3DSj4U5RlPvkcgbTgmPokO91ZnL2jXLcCRQRD/a1ij2VhkNiNL+6H
MEfqsp7o037RtrsjkgolL+b+jPT8FB+ZV8wRcnchJNOeXdSHgzH4EBM8OyT4yxi1
RlVQTB8jv+FIKJ1IjUNAeTKcLqgpPQljMliT/Ujyyqg2lGd+DGgYh/fI7HoQpYen
tSfbi9HNqfq8M8fOSqzE8kQfgz0dLS3cIhcJc02NvHHx1kHgtLcOpXoLEWWl4/DT
EKwHi1FZINNkZW7ZRWBkLT+17DkracTu7aUsh1Ub0T8Olb/Ur7sZ8750kuKZ28ET
0tgaRlT88lLon90G6GBOr+oSuSKBFb8+/YIsplXzqXnGTbUvWgGSVyuOZYY3BL9J
AfRVr/1USOjsqqjH5vn7ArUHx27TVr8IW0/e7X4E6mty3f8qYdkYpCA6sXHSEyw5
2heAhdlJgEHbA1I8zOa46ctvNcSsVL4nHCUr/T4oBx7L8uV6bs7CtRit+ksThSwa
b1ijsCNKz730UthP4+IewXqgGFp9JXOYOfklTEw3knlTr1dXTzdtHxpPx8jhxXoQ
R0P3S7WymHw+dDmM6iCkuoLuERighI8tvcv3SpydLJV2cSTlJVbTqR0R465r5d5I
0lKBXuizi1909bS/SlLiVaYHSpVvuJT04qpRbcjp3Ia8p625vwl6H9AWwh9gJScf
BXRjHuxr0+B5EWE7DlXhB4dFI6wkDtvqjgoNjY4ZPoJfmwbohUYaSs00jwmX6M57
1ZogdXcA4IVApYzAD+dSJICrwwvjPWBw2UxPFhHQg9JPLT4pnQihbbXWJ7gVWvMF
5SjGCPuWjlrp+6LTwvfm/vbgI3Mex4T2OgLwJUoG8bxMEag/xth7Iql6luJQ76Og
SqojGMG2WL/5g8V+U0bB3shHCfc5fBNQ/+m3gCoCDrb1JoXN5wHFaLvTOXcmelaW
mGKIELAR5un06+fkI9xdDUVFYMGV/5y3VpUxxVcyPC2XXV3AW0BQSD5aJApkYsFI
xDGXFT7NU5Lj7NFwOxYjVt7I5guVmWwLZ6z089P8d+euXEeEv20ODnSNRlz9xoja
VrujSUyOmj2/EVcSbf8ivGNFelan886OPHUEgIlSrmP/eP7yI709reruhpltBcSW
BOhkZsA/4vMy7e46j+t/EEwC7CwSv17Sd/bVAEgMr6acWgW9EdXYi08osrV6UJPo
OBMZMy7lnVranvrxTd/T43tp+NVobPL2k87FnfjaChk4X4C5NoD4YEF+av/bfpMl
P+GuU1aRRy1rmAdkM1SOgPVj2hFR0GTAAG0o8QCAYC1OPILQI+S/vGKPr2bELAVR
++nePzNYIEOpqYacTbBphHsyyUODeDprarCCXmK+99aAnnsTHGkkKvIM3n6nK3VQ
ka0ZqE65X5Kajpf/TUPLIAtnDcHBRFJ/ar5+3sss6nXQByVFGcyqy2UpX4vI21GN
FuOpQyqS3vZRymuH+qZcTkrEj6kmf7TK/d9caG/7IDQtxQxjMhz9a3N0ttjeHbAr
jlpGkEWaoel9t1WV58/8PULtDkhSnHYvRoTXkarKsWlWV62BUnD5FXCWJaHa8T5S
DwDH5Clk5AGyuBWqH2aNer1B8bTmLxatSgO71SoBShFJoBqx4HlfDrZCz0yBbqzP
lCmQEyAfKSBkHPtoU7iKmyGERTfE6ESHKeuaK/cx6mTdegbrm9teLkvCG1PVU7Av
r4mM0k63ZtnkqoJIv6oTXeLvsIIDWH1YxkbxIZp/2Re8a5gOVXqe9TgC5X+TIoEm
BXd+o/K1WaVCkQl22ui3n9vyqMZHa8A1In0UbtDdqnzE2QwCXBZKAaqbcEqwoVqz
yEVC4v9++w7QVkLXJpXscFkAPc3C0uldOCWm0/5ltpuiaKRdUBU40o24mbN76/V1
5hpj6fzroUq5p6bFAN4CGv9jMAGvyGNDXtSiLslrN2rZYBRhtTu7QfSG7G7N+uQg
6Qm5PiI1uUvTsfC3Eh5g7LZUjb4uKRckFL/8QZGYcDspLHcsL/zBzz7ldI2tDRXR
BSbl41bLWRSi2FjyyUUY60tgJMM6QeGBiulCqZ7UvjkStjHNg2B5g57YFF2psabV
YeotuzbXU5lorVunRc7ZyVsC1q297jUUEZBjDawTFUpmNB3ufKdnL3JlWhUT67Ur
yGz00dXv7o65OC8QFGBlLeqIDBAyNaKtlWFar+1KdBZySs2Lwyh02b1EOcxq178m
4aaWB34ij5rEitZGfg97QjrRpiPX2mzKK/2X43iJvoarwROrSh/HdutJbGS5hOAo
agHt8BiYKOY9vUEQYnySN9KPzpNIdhSKAKXDqiz5o4DYIeil/e5y3O+8CWt72fOx
2s8CepwEthL2s0BsehC/PcZJqppgjc1L9HG+g+WPOCg14586sM6JPkwCFr0NOWJ7
eN4YDg+dpXS4i4eaOLo3xzfv2+HkM4l7900p5ye4+GK8LM09OwFV+LVQgV7XFwwp
RiiDZdxZHGOAj1XZ3P0TXGMbNmHSmvVJ01RGPJhZolZQW4hWqjT70Gz2V6x1JSq0
lz3bYA3ULG3/5VDhy7N5PjdUPijUc8pvSaf0oIfH5lK+oRImRMUa2y3Qk/qlUe2j
GubhqpQtaFQCxAeRVXtgzOKUmA5Vqu8QXp0Oas+fkM9Tvg7TZMokS+NmE/htkzQA
EUX8yVU6wNhTk/tPVVlHg6YvQjKMyVN5ff3O2LRsn4UwlprdoeSK9SlgkVgSd2+K
j31wRg+1+R6rVzsiS39l8MVm1C8ZU8pqNFrKfKCPqp9ylR4W1r4db2RPVHyqouPV
Trc9/BHwYFiLlONkXGnYzlFOXjZ8HfcT2IlCGjZa8ebRntSO2ZZRoAIWn78RJhQc
gbq0OWjoQusjh9hzLEPINi/IvXhjh5ccUlCWLBvMe6l2umAvkRj29w3vaI9fstcP
2JNj/tEEuJdJPJGwo0ziH81wbDn2FWhNhorGvXlARx2m+bFEZrLqmqF8jVRwWjai
+poC57mskW9HopxqiW1+0e7WRzAfF5Oa9ZdSlwwPIcNf6N2xwke8TitO4C1STxjl
C/ZAR10wfKSohZENiAq+aKRos9GTnJkvJdMiYTmo3HKv2BOBy1+sj3ylUTwLTMuw
4iYs2yvAa/IWb8MJWqZUSpIyTblaCEHqHF8pM8yfu+0h303OyTU1DyRPtDHgooeD
QVMTO83DujoVWsQqJ7PgmU/yJTSBAoYt4gqe81uXx/whTNbEhvhJ9yMTG7HVnmCb
PxtUqKXiLzWWYGDILf1ozyPusqDUrluudoUMRNPT8s0Ou3cz9+gf2AAjmaUGIt9k
7ro/RQJBfV3bzxoi5QpTjti/+SejNkQd5Zs8KPOvzaY67td11DDq6eE/Qqr2kDF3
x2Z4QRZHxyE80HDn7zrW/TY9Khv1qssMuUWgBjyLIxUCNwmKvcrcTgu2v7Xe7nbV
OJgyOrG5wQnaX5gwjSKGKJdgj6CZvHaT/vjZKObT0jx3gHtzdboIldWbVGDK7m6g
UcN7rmKeyb0v5eLqgWNdVV7dDE29eYsfiBZykHUms0MQTIvsWbujXw3cVk/wSk/L
AkhEf1yrAmx1Dm7HSGsWoyu3fS61bBvUo8RJPi/3PyPEbU6GH3/s4o7veaz9R4q7
T4HBEiPj3/CYCIxEGDNPMtIq3Vz8jODdil/8iuIKek+DGfgFTKb/0fmZ/WRqIeLv
///L3yZeyZ9uc8sK7yyDbmpnWP/hYcCmzVTRx0J9RpnK7Xv+vGoBaCtQJDVk53Cy
MIlRj/4dJI8JvZbw++M1h2p0qUbhm2DcVyrZcnYHlt5JYoUHawoUsO0q/CKfwnMj
JfpE3HS7YoWURM8/NWQSyL1Fcz1EjfF+zOsJcRRdBvhRgsVqNNtm5RXBaJiiDS/E
LUYT9oL7J6mAVqT/Vog6TtecXwh5MTEPP+3R5/LSTMa/XVlpBV4xGdPLtpyMf68j
kLdWVIksXRSHc11v+GQq+o9Tw3V7qihcfwpO4BRkMlA/O3icXC2L1iRkr3duJfw9
S8EamvYx10xUzv4so33+0qRp67FFtUJXLTNiSXJoaNxZk9gQGnumuWh7+zuCxCTv
XlfjZpwAPrm/LEJx0K/0hj/zYLwEX9kh/SdvPkHPQjZe9+Y0PLPCQXcMfwNaTPSk
kiNwHGKdzJEcF+F8jkE0+okVtp0h63nj4vAUOZdy8n+f/3MHXeRqoxDur00cWSoK
Yd6a8F3Cr1FOOZGTF+Ij58SDwMSER7ZREDPvOxyUiSL1G/sJJAviqf6+9UnCSFqq
DsLlIwKSsz8ybKO+GbeMqPDe5IsfcxyHMhaQ/64N4azSsogb30xVQICBS0AG+e9f
GXjPabYIVGjmxhjUogDSRNCqjpJxySii/rfV2SyKR6yF6QQyQz4zFLYdj7YT3rrt
sDaq3pOlVNZNTvVkq+MdgRfOFCaTr3pLfd1jvZsfYPJ6+HmsdEU3hVcJWTpmDkF7
q0qpZZqa+21lian8Z5q7O+/BEN6H9/EL/ieUgX8YfhOyp8YH1KAduTiRCchIUxM8
YE9f6Hf7V2BRO9rdCxjJwqe5vIc+jUrAIF1/4zxFIdgQ9y0rmZWcyo3RTX9gX0bn
l1coK/iI14TDoYNvxbKxIRcd+HssumpFK+6R2jrAkT2CawrbDtTw5fWwxclQQHqv
cc3txmQwN2jhPMDkb7nQ95r3kWrgHJ/z4gnq0MBp/egNh94WEHOsGVWOcc6FOf/G
T1bCkSn5UUZX8EYbCIZ1ia0+HbJB3gxM6m43ZJiujxLkLEAqLDXHlcwc46esYDf2
6nzqwnefPiYhHi+qy1Wa+Wbtt1wLjuFEwbCTBYMWHm7wHSvK3QrDRyV9ATOeMxYs
LolUKquO6P+sFTWfP6bo3f5lHVKDfTnm81tq+WSauKQ5WB/7BVbPBtGC/LbGjVmG
iqmx65oJ08tiowTmOFZHRiQrcjqZo9i42evtAh/Bc6B/Mfzj+cI5CiniBj6dpBPN
jLi67pUqLKhaB5LNYZEqK2gTi0P+lagHSpFeb5X5utk0eNIsC8vw8JIColNtJf/L
RlKSfC+/P+3nZzmy37x4Eygk3DNgvah+XuRb0QNjc8sdDeJHhWQgyYHEYZupOdUE
R2qnvsQ1rw1ZyhzI5juTt/deU2ZTl4TqEEwO52KrXHjOo9+mDn5P0dTugXcwinXd
8AP3WJEmsQApuzMIfAzrMKOuQktKiQRJHtkeZ1ME+ycsYZbp2nNDhtrWT5IZAh4x
Mbd2REGH/s6URb0SGyT9m4Ebubi+3xq8kCC0+RwAmSAyVIdop0AWrXACsumm97mI
LHUQVOpWZuznUYitai6FjRKAkeUGkzRpma9dAoCgrL5AKxRLXROMXhZsylxqcyla
FPsVDV3yMidJOSE5mDwdBSh/q2fqTUKocVirnaHup7+IbrJFz/b53m0F4pWKvI/d
3zBGgGHKwDmxnHqxqDjXPrIbCgGFn5NgCYvL5lnsUqa2EQAhZczU3VwB+LJvDM5L
SwPNlx0mFqSvK6lHBcxOOVtULyL1kxHzn8MWIyfi1K/dUYsZhq0Pl0NTHVzTMYe+
Ek7KVz3LpWFz48gsA/TBdI7ZH7R0XtQjA8Xwd/+aUt/qML5phk/aILpDFxa5/pBG
OejtkEWA5A+sKlLA+SnheSvEiHok3gxquaRS3WHarbyDfjp6czeRbZfeIE3ZXN8P
SUF/NcdBd/6gymRa3tpIVN7tStmjtcq4JX5i1q390NdgG7aYvgC+JdVswPA3fpF6
AITDuXrVDvTmWc0shSZ6EJjI62xVrmiTE5OQ1ZK3pWQs3JLlBKqr9jwpV2i1I8vR
9TyQc+srtv0c31tggQfu4ZD3H0pV/0iw3X9m1subTIlIp3YLsK/vhnT++rHYptgq
ftPPZ4KlTLxk8XbpluvT5inLZepcJpcfebvVJCCdVGm3FXw/h83PEF0rkOOt1Uyj
XFkri1XTB9/y+tsEKlQefEA8jzfWstrDBwOS5XIiNiEhlq0xULtxLYIlQRmJhzZb
AoXdBHIGga88EOGknT3lV4JkgMdoUIF7asd5YFgw4ZYeZhxNMWFhAIOXSkfoW/Nk
PGWnWCm86Yo23T2+dITJekd65C0+QghbuQjjay5N8Ynyoe808DeEfmR2NR5sI79x
ZzQ5oaO0kvLWGCKT2/dyU8GwBuvM2jw1pRZ+/CdtmdQEzTVoUgZxum9QfesJEjQm
SitIXVW4RHvNHsbtm6kIuT7V71iPvDMYsf1pFWbN534vsQ4w6TPG+miJvBHQ94Mv
UmWC2vZMRvurDdA21xje1HHyb4Ul9sAhzzqXUDDk6zmvp7KyGzE62HdOj66Cjp9E
vOE4kpEIa2L86J3ShsHXOzH1pfnlYPr/B+Qo7I9wO8NkoCXqXSXo5YPlQxVTDAUW
sMknFBzM4wGYu9mE/4ZgOnRhvzjMj1Lp0VrOCrSsjXNmNUYfAkG8mwVQ3m7x5E0w
SB6TKrxhr5UbZTREYtDT5ntP5KXL9J8km4SXR6chF+2om+lOCirX20+sVs+Hx3rd
W+BvQ1p/LOpI0QJ7xAMiEEUlK2P90Klwt9YwbKjs4kRWp+GMDLYjUxMrhWnbQW7/
wsA2sE+FHCPY/+poU6f1mzoU5WTrnQ/1EMkQxavIzcuETfQefWodhAHx6cP1bj1i
eZTgxcrhfC8vNzjRbwbc/osI6QDLCz5G+UbE0gn++1VOEIeXFx2Qz9zHTsckSj1u
5RIRUKiEcKyCj/XChjIgjOjXpZc/R3VyW90kZ5Qah0KIrOH0DsqsY840e8qB/FEH
lUWfx91saDSbGKsx0spGlMun7NQrrjZZ7Bsf+rO2+qlGMNGsyYVLUgRcahffb4K/
GvlXipMsY9ieaFXvyuVfr0Gsno5SJTn4QkYPOcKXq/6HPNAQld2pABi0nikhMwzB
ETyerDasXa4+WBB0x3pS01dOQWMxO3CzzYBq63+fc9aWKi28rays7QPpQa6YxQAi
nTPtpQZCYXLAFxaA3ZF1Rt6OqV3wY33CADll5cawLGVMj8i+DRxUSV3taOgvjx7H
e1mVc5TYN/cEHDK46ZdwICa3NSbUO4G6vBl0uIZPvOq+4Yfd6WYfoYwxrpYCKcjH
/xKT4EHlS9XVIuCi2Ryt09/Trpgz8q0TxScFxCS2upMOjpLc1T9Ky11/ONIh1nuG
ej8tJVtm99RLVmk1Cfe3DjYmDRul35X95YoIyCVdd0riz97lrtk6ap1yzaNe1N7S
YPwKW1b383zCtvhu8liGGkvOOomT0Y2xduaLRo2oIRYeDEbUODQYbN3+BCTU/SdC
8tpItsTy7SRB2dun3eSgZ+ir+huPsmGdiiEpiuEHpYmZuYHWmvw35BTSJZZH833/
cQMrvS1y+Ze+nwjCKHs9K+fM6XTIVdsP3cRRKRYOEZIo7aDGK6d7FnLll9hHzBm4
DMs6fWIoRFwsKaJwjJ6IWDaOmqJN2AQ03vHf7+1ehdAIOO3DrINQtd6Ri1qnoRf0
30B6xx1RenL2NBjoVxYDA7/u3EpsJZ+5uBbW0kw4/Q6kaa9kpfiaAVIuo8U+tu/g
hn7i6cepCviQBrjD5HkFQ6VmfedwprgaeQCegE6/kj5gIPuEhJ0bpTUyPx/CVYXu
nACaQwJlm/qKZXwJHGXBfBX/3SgePRVXyGEdJYZ/LqOXMknVTOXDLjwHZVZqN90O
W1z2Iw9xA6Y8uQea25+fjZHv1/Ah3V1mLcqKEO/QH2x2d3pzMRYKaeRkiFmMjZSe
LlxnFJDUC5kW6wkt5cRtOWYJJOMplIUpAaP4clAa71poxEgSKXkj02zzbIafdzs/
t9yhAbyqwAfCrkHJOTxKEIP4JK4YpiUNNlzYQBnjkZL/udIFSRnxdZ9xkEBx1K7X
Zd8YuIMcmYc0/jjnYWFETPdG2PtmBbMG+cPjjiH6NZPLtIPXcsvEIeXjNJpyyUgb
gtwjXeuypZQU1QRBv5HqvclAyc+uJSUx+F2bLZ0gBBxO7KHmpS+E+5DnoAyxso2l
oj9AIxAj7NfBxdN+MduARds04GEBXJyfzvl4+5+W3WLJoqt/NvcI5tk0OKPOZTFQ
jjA3JkbCt2NK693gKmSrurVLrJ8Ra2seCFRAJaPFbQvik9ZmDo+nqJSVUbjvT/rb
BUrp/qp9nKVJw0n5nI1LhDz3GHqmYkhH+EoffVIVqzMNqbTzNXuwIAdTE3aHk726
f3Y9MZEsNTYpZg5VhgYRgKwUayoO0p06LNoH60+oEjeu0PSSJmx3MggOXd9cUwMl
s/xzcK6y1ML29AdaWJbfg1f4crnLOxapvuUcl29mCbYcAQ8/CQWN3iTFJRvr/Ga/
RZjamaYTFutr4A/QsX0JI9aAhWernrJnk5zNDSy0vYvtAKOwQjOjXnjdiF7yIsYQ
7kqdQ6rsC5X/kLqaEzmVkW1k5VgNng/yiqPKyPaAk+KYCYpHCdxRE/LjTBIc0dxy
f12zyR4wZiiPCPk1gUwqFiZ5kF3CDFyeSjEAEShbo+vB3ypbIYIVgwvn9c6gRE9P
hJTb8rLRMowAdsbpTmtWYts6Zd6kHixX2p0wwHn/FiRN3uL4mLQ1OmQGtERiCmol
Hyhj0NNB7zOY3Le2hVI1C3Q+IgyKbuu8zvhD8meihkxFcRB3M9L7JwcAJPyAo2lm
6hf+K34YnJAVe7bQd7v+vfuJveGut77R8+YU6sOh3DiWutecYY/DOg5hgOBQXhqZ
+Zvm3NLsG5vs1PSR5+MeWdMgIVIs//W63YlmGkNN9g+BVX9NpvtMhL3bgf8Tqd/3
kFTbTq1YLC5ggYczi70Ae4ai8+fq7XbbWpMWFgY9pb5fDAO5Nbi05iuW9HzQSTjS
p/7lv8eJzgFuPn8qPvQ+jL83exsogqTBLDjbzGNspPGyTT3QwUvJbSrSn3zvl4LR
6I4bFQ5wQADFWBXVOKv9z82Bo4ALY7MPnW6UOoVGAk923GEMvv5hFZdnigvzWlHx
y1IZ8a96XXv0jtscnjdPXd+38+MFi6x0U0bA3/wfT/Ztea9NfEVIMUGk67BZkUn/
vccoEBoPChg28pPGmeV5CeBbWeKNvTtLzrMuxSo+5vcPpNrY47OOFuTKZVp+vogw
GZ1LLRU8HLhcGbFA5sKSw0ol8bnFU7zq7ecmaP5eH28KK/QKEJZ4uZWBZHUZamMY
uTvaru3APDGOBzhqDq7HcF/HVUgLr1c17MKDhrsqeC1jA/czob9bqPoYnWiPgr5H
OoezLWJMyv0M2VvzfLUNERo9OKW14/TRgv3UOsilTQDhJ9KiojfiHKf3vxFHKo8u
jNVWHDCWRlzH4o31ireq2jyHkYQmIUqQKcxuQiWweae5P9dBK9g61XSkbZV3BTF3
6NQkzbu+bNRIKsv85Zx8ACaaCu8mNlM0Rin666nagsNROqFdEp9r63G32/PIgbpf
AZwdD8wdk2BpuQd9XdCN3K2SlkIFIMG0uHpG3Sxu545Q7PjvCd1lSatDTVONcOuk
7QtzJTukRWLqeTVHuGx5RjIuOPFVFgIpYGt/tgbUilAKEruS03N99nEnei6lh1XK
ilsYUzDMcYbcVeVoz98FojjvtRL52ciVZrHjlkQ9QQuigxzIniV1mSQpbTty3+fL
uc6yBbjAuAwcQ/KjZ/oS53r4rDXlf+OyhTuuf09ttcD+sQ3TtVUj6xOxXQMmEX+V
Vfd0T5fTYU/mNC79ux2eUnVBZxnwzGAa2XYEGHVZPbQCTXOc52a611VUxiY0mp5H
jwA6cZjLB1SIPMBgEpT1PgxCA5G5842goKRFLHmNSoetegou7HvTYPZcC+un/ikj
OylQgEmyMHkb+1DS+NvjPJfE/aE/TbBdsryTdsEsQwxsq5qzpxRbcOoU7/Se9VqP
lpCARutoNdC8NNTYn8xKVkUtOIta+J/JUT0pUVb7GcrpD/oAdJptgHn322aWxCo5
bAotwveMyIqFP5izu2qzdEcyJBs27HC2x0fz4Z7JTeyomV9cBdy+1qLyzzYUDXc8
gRrGMUctGRdI+ZICuGfpJnZybCa1kUp+Q0mdl3gj4SVZKapdC3OOnXOjSLxM/yLz
Migyl3eySUsFypXHb4AZsEvGJV7IBXEmtkeljmdZc4+l4eSldH5pCqGEv8ezcak0
GfQIley1oFSh+upM/kj+rO7ffYFJgntgiVLR/hkWL3qKawjTEfkxP9jnRGtFKSjO
zI3RZxp9SQm6NFZV+b+tWOsIddpOX8NaN/lRdsDT4UuZ3LOYAWXOMJiLDjRXeQYM
PcPmVq6SwUkXe5+OBTNVZaZtUgIZ+Nqt/RWpWAPx7eZY+Bu1CPe8PgsIW3g+dTh+
NvFU2+VM4VrZ8UCi0CGJ4LYIwcfLMb7WyYFh5otd2DTW1h2LvMPSofbQoRigl5Ci
s53Ma5non+uvdfhbvHsfVRrAsceyq2snaonCj+ZfSIwA1Kp1YNl6+o5kJsYPPJ6P
xvlVbzqv5K/fpFy+XSaVxHUXLvLbC71eo0jTcJoEO2sKFQihA9b18LdHwFHU7H/m
Rv/65qHj+gqlLpyAVpmkSwSgmd4FY/spGLsHj4MF3L1MzHM1Wvm0diVuiExpLVI3
tdekODSBPeDwSjxx7pN283rCCZEnHte7TnFqo37n6FRF2QBRI1HLnvvW8IWI4oia
p2X7WVVHEiZwLO8JwIuswYfxJeVbVwLDQhAysVwoD3PdfYVb10qbxkLKSziSaW6M
4kJ68EqnHVZfWs1rkd2egYqUTHmqldpwzpIcc0zur03xYgIOWwzyqJZ2JR/hLl32
038WTA3p+1goGNzLaAjhpAnpfExuxxRrnxb1NmxGs6uV18s3PB4QnNjKs3JM9SHO
4HNBf0WiSpxdgrTYl5XMUNVS1V2+UDu+R4Ojvs4tQzVrEC6fACncfLb1BAcXAacT
V+IiOR3NKCmT2n9lr2L11mmOH7o5cXmYSI+u8r8/XDJo5JUUTqTI+qjm9usGpwJD
H01aEQbbRm/wnwioQfroZlxwOQD4sAsgX/ECHMVj2Of4UB2D2VD0kqXY9kw1EVrx
vYzKN0y9C1/arawAIf4bsWW3bVV6O/rSw+/dgWpz8e+p6epQc0xLYNyBUA6cb6rJ
6qEdiEIGj6KV7DUvL6qj1mz5WktMC9i1LLPRWTktn5ylT13D/jMWI49GEJ2nIBML
4y/X78q8+MlABZAgEuAvKS231gPh30rOsbsv7B/sjfdixAdBp3muHHuqOVeGL+Nm
S3hOIwpjjojqQ/7aumECM/RSJhV0bpZ1uZAEtmcMCjiS9r64X5O1jmGP6xxkOoaF
+AHJOm48XjJMVRGSxBuTjec9eNfIsl05eLXWXS5TQvXTZzXUQhKAgYhev2r3iZXl
sDYE4Bo0RSA9NqylLuIcm0vOMwrRTP7WJQgyhcBvCieg/Y0yTrS5BZKr/bJC3a2p
QeiF5CRg2NNG4dFO0DNsmZiXI0PBGcW0/XqQhcTGXK3XHde1OXxY4qs7V8FdVoJw
+xeqeutsgHoQVsyxEobjRUXte1xav8NTQWhCs5PxO81WVHgQ10GSx4lsCNH6Ronu
1Rta++fmS7NkW+pL0aiJq2Lb/zzYan1MLP3SASQkZRW9do/B4IT3VOfOEkqHZ0HH
O/9AXKYQfNzrnqhrY51+P1VHd7/cpqe1z4F/gwpEv6r/XyE3SDS2El9hd52E4+Gx
M3UJrumg8fmFUARld5juQKnpdVXRbZemmlTLTr/xd6023fymOJVMAC915Y1WP4Ib
62c6dVjvmG8BQfb9PnZbpCI0H9lK5zWAWSQ0oec9HWRGMP76VVL4fR/cXvT+PEt5
nzH2gf83JDMl1DfN3NnA2Za/t/ZNEgaVjvvj01WcYFLm0R+2gUKWskpA6MqAD6V6
VAm4wyTIuG3mVK2uslbGjgcGcnVGHwr0dMBWyBq0FwN/oTBRG4nrnSKV71CTD0eT
fUqNWmtcPGyvbRxexQTKEPCh4K45CTPeq3gOCB+v8JDtD+Y7NdXtKp+madX1zoEg
uUehbuOwf/xG0uAl6xoinwoXtlnat6qgX+HSh8ZhnDp/LXEdajhl/oBH5sUV9N1v
MTc41/nFV1/0iNbHs2O0tgc4syca7N2YHjcm9LrUkvaMdoAp1hgaIbMxmJI+4Ua2
Z6ip6geaDqwJYu6YqOH6EFfSpWTi5M8Z21fQUKy8I3U52rRtmyMKF3V6J2LqzeJ2
/3vwbJDfrb+ygbyWQwL0aEfIdrBnKFZRcNDaFANU+Gsxpu8Ek1H3b4zXm/wyz0s5
RTpf70OIPOlNmctH2+1sWhc0anx8FWpFXi7UABi1aEM/ZYsOBYOKw2fRrDig1WTG
VNnNe+VTB9dr48sHUw73wjZDZ3XY/fTJzjcU2y9Aiqjh7Y6K6Sx086Nk3oJakmVi
OZn0JQQrrsPv5qC2HwHd34AuX3mRId8r0D5jiyyxotXEIQsg3nybUsOhH0aYzXde
I3RNiBSf1qv3Z2afpLHJmAvcyfKsAwFKTHZLpV++x0lGu8QZ/4dshs/2cpLS27uv
dmPM79WGomKWSGcj6vey8/B7GbbU26grGGq0zmwCRBsHrZ3798AuJLH40WJA5289
Idlqx++gJeVm4KagbVWyy85ceTY0ArGXtLN8b/YTOKJAOLGAiPEqIsAp4LBvmhc1
vuL2VP4/S5nKgu5ldZf6tfZVHV6Uq4RG1G1prBjW4/MDcYh8dzNSFXERBTZi3SNG
QFuBddLQVCq4OJMhTcTmmzar5un4KxCUWhgQ11QxKe617ptTRkiatuuUrSGqzUcn
Ehm4swoY6/kKIO+edtXAReQ0DLVcQ6yRFxetaMIATv8Y0WixGnN9AEgzTN7Wq+gs
Bqu8Q7583U7ZSEr6u32+C0LHYpxB2XcCPzopvKCsE7JFMAFAhux0GyX88YQhg7gn
vC4CwSzznxAwNvCu8kqHHdu+uUScaRTMoPnoJ/QtLyw+sBHzRBTKkgvBp4cAtFX1
zkKFg+VOo4dgREdr2d2PlhegcztGfr35nhCsQE53S7tS2HJ9rXv6LIvb/ftWVLOR
hvB82rKktVKfguyYm+A5hcc0otHAqZk8+fqkmWqmITaQvJ8yoCXpxuFjvNz8IB48
P7SbDmRMR5OvFmA8UWLHg88n+ddaTd/1qrM4J02q5my05ig6DCW5RSYleci59CtY
W9K7JQGA9GiymWW71PZvCAPVevjzjRN2RtLkfZAxdSy2M1bW+ADmXBC2BAmxkuLS
jpBYJYWsYL0PseSuEbNLMsdf+ByCoxjiee109jAn15z4WzFc9O0brx/R/G+dZG2d
qjI9m4D2KaEiXf/T0Bz25aIHXqDtfFcQeHQelsupnwHWuhqWzGX6YDlJzMMjF+yU
zRlT+AtabSkLbEPzJH+LYwqDxXH15DQixSXO+hjy4lYvvOkukEC8WbDYbsi7dIQY
+mq0F5SYK2SjhsDVpepLZ1U/ODFaOKgRqzkl23XeaGmftRdq/Z2qutGXjPCqsae4
5+ls0IZE4+uKup264xHCCzXCbupRcLc8p3q9rnx+xAUzqoq//rH7753ItEabZyOq
P8sZA8lnAwY3E1WQ0PP2eXzkYGLIV+9D+7WruzQNKpihK/5DnVFfcYj+7GOexXg7
9XLGJZqKHECrsZ+6ApEPeeYrboEEC1DKc6j3rolzRddzMWjSSJDQ9hD6K9f4Oxh0
wTZ71rdU9PJ86jt2AqxdG5O+mILrVVaM7SHEO+FAm+nZcDToxVijKOmi41tAdzmL
EtrbU2TrLryAE+gTN5/TNeymGE66xVDKuW6i1+ZOd985/95Xmc+CNhQYsodKb07O
ME5EuV3Pt3/xmw2OsH0S1y+Ley5Ll0LUdqsHmXv6/QHI/VHyuJah/Aq5mN7zAuSD
m9N23tooCbWDQCnkVWzm8sSkPnDpMxkVF8XOVvzMUN0muejxz0UhoSltihY92rKO
4mSRQJ+mPvvTQp+HnGbhXtrytTpIXijELhKS6HTbvz3EyPgTzz5qbB9SLF4dXboH
NMa1ebrLiKgAFknD+Fmpt2Ml1ktEsrn3iYknTA7Xd1xdwMY8ZFRfbiFHQLDvnShk
oIfzPsVz7tbSnRhIUuoMbYOuYR4jYEEejXX5s/kr+DEJpX6cNs2zMFEqH5gvZ8y+
6mwCzY4F1i3OVBr1mTbRvq2zLBLhJdsix10gjKwYe+xr1hqMc7uRf2CFJh1hbU1E
FvEsNeo+wrVOS18O+NfUCr+lNJrTfyzCTSQ9VsG3TrT4EYe1w/Gjy2G8uouVUthU
S51NKVukIQYwtl+DUurnEsgTL3038vyDBMeu94xMBdBPFm2A71i17sUJGEDHghrb
NZf7zKJ3YYFvFER0veMM8FNbcCgdPMEW8yWpTtYDUJrh/MVVi0KQadd8l+woVvsR
ONkEC4/zHzV7AagPa6DQ36Xx6Kyy3OjZ41AGI9nbuO6i8pUhG2hpUM6/KfeqMj+l
B3bc81OzQWOHi9rSrZffr6UctupnCQjtb/Ex1YpX2gTd/2Ho/A3zF7W0eLX53Z1P
xFrvP7y7UgyPM3VT17DlcwTLCFgBxvw30HQmc2ZHlgLq5eFwj82jZUtw2XQ/SCMC
I4NEdBjBJebbyybk8UlW3QESzD3L2ndiXewLysM7mfj7gOeAf6TXnlk34vx/LLHe
Enndpa1kzBPzh1yZkybgkDy2ucOn4rysK85jnQXDzKzhNj6909bAEOQBVJfyqNhO
v/Zz9ok2PDgRhjwKiC0lVjOcA6cFpEPsB028gV8rB0mG29v9WfaEn/Y0IKZSIEOs
clvTfQqgGJS01It77n5ehh4MUk8y3MooqUUgAf5rn6xKLKY6SgLen1b5pPibOMOQ
9hreX0rRU7+B0azG3/L8MVWhwNeRAtbZK1EmLMexiOkW+CMLjjpneUTsUZKkuREW
3VwfKIAs/QdSxK8Eb/i6uefT7sXNtwoKuVRnHI5k+OTyxBzaXDJL/VpVPEpcWnSO
5GYBNWjwE1vqDYLJ4S65LYzO4xy75Augehr5cdjPoh7FpzfcuFxyz824zrsUY7En
mRgWLrhQKxDMU19hKTRVeG34KHtEkA+XFmDwRIwzWJgLs1i+IiIeH1eTtV2xClGX
n7qVUbv/QGSmsXGaPMWbDAXHlrNlmDWB45aPSgyMs6EvvocxfNiSf3RsqWMcaxda
t1E/+TGZ78Yrnf460f3+jqCDAPCsIocji4GvnZj4Rx2B/pV6k5ZkVHaMfpHjKPFK
G/bkScO0mi92+fle0RHsYE3Y0m6oyhpP7MKW4DhtAwmYnQKr4aPzYD3V4pnXxZMq
qBSyeBXlF0YRUIWnayr97VDBAmjSXC5CUTpGOxQZ5PARIgXM/qrF8J02iahpibXg
6d3HeDMAs6A+v88KB38cGrbuGYlel40irWf7FuBULl/Dn0aEKzNrhKGrZ3yoPopq
ufcyTJYW0DewYghvFdXsDXLVo4qwsNr+gCvhVlqe13dENn7YiFsKhyssZbzfRBbE
RXfzlDlQCM2Qw3rmoDczBkLUwwO43ehF4DhdNkG6XYzcGLGZrITeUSKnKUm0HEFP
Vo37mgPeU2IoUnNdSvEMgbffJqgVymSQDybQp1P8aYQZ2gmBQ9CulCwor9ACavyY
exov6UCZhF3jo3AvReKYvlToaBqTRvKb1s/yQR5xEvidFPxsT/Uv6pF8XcuVeKyi
d0D3/r5lbzG+AlfS4vrn4OQxQT9sdn7CDQfc60WCf4TVlEv+Ye+RfjaIADIXPssQ
NO9wyxAAiIYzQiPq9OkpMO4e9d7f8SxAX688qxRUUvu/I0SO5X6Smkj5hugjW68T
CiR290i9xGb/GKugp5l2WHRhrdZAyKKFcT+3dox9hj8UsZi5tD2Z11KS64zCi/B5
dkxKFtbQq+ubOYm8rHwFPqdr7rIHKKm10QeipyxLLaizgDdXCgTwf0/Rtvz+C70j
rKq/psInTsSDbXInoipnvmxNp+tmAHrb9O7YKYPvgFboFseCguYw1ogJihqMmntB
j5Yvper7kYGNnEL/s4RWnO7Xl/29nnw08moNetYpJpj8eRXYWlh8EtlHd+B6UMhW
tsa2c2v4z81WZLXxeEX3qM/mkXzFeWpziz4c5Ka2H1OaZeYg/ArmoetN3jNvUi1U
HRm5nmS6U3rY7z89t15H4Y7CP4eDv+FvPO+sz4WnUYvPCwQ8sw0TFktwMmEgb+b9
RJNvA5w7sCzbO3iBpTQJO8GAmcF/hqg9jyR8JGOWO/pcEyxtksIGujyPOjaID+hh
D21BDBfR9IJBBPPzUYQiqIUEB0AAuntLE0zUG8/MgRvDdZwOItK8XjL44l/bu5tZ
knJdk7kC9Qm/YCujO2ICfDuZVNIQ/4tJN1DJe01JO9d+Amb1e8CpDB0zAnvQyWDn
DPacmGnybtGpcr++3Q5lYPfnQWSUAgG9YhLt6Ju0LwpjhCCwhJS+nxArptAMgzzt
SqdijQfAG4MZJ51nG3lbh55m6eFMURIA1O1NKy9lVNwpH0WxzpEY/tONJWZUpGTK
Gwi6L0Thxh9SUmKjo2x6uspU9HDKMIrtEA6sNEW9VJRsEBHRsxLl8BtxZQExp1L4
2b4CmeRHNhdpS9NPEHqw5tSTdz690kEAXGniGaGvCyPpMeEIBn/8A3SXXU3yIWc6
1bEU9lWsRkcPg29VrtHmlWobafX8kHC/AWv7gSo1S2Cd0YKfkjn3Qilyry+3mi/D
P9a1TmjQ539uLzXVqyFGpICt69w7g4WzvAJxiGZO86XyejuiXSj7W8AdFpxurTVj
/tQDY/zD15OFL0A3CcCsg20sf6gdh/BQA1bjFEWKF6G1NYNf3kYtxInUCyBO0ud7
EM4FPQM7hMhzRQjOdTuSGJUAs6zbKhrOODh+16SKuec0pAVkIwiBFYAWZU9kBFaf
ho7Kn9Y5aY4QCNf2OUp1Si86UnCXGgfnGd5BWWRfcjMIdou7hcaS1lHIRpujqA47
9fWS1oPKADTIXobz3JRQx0NxxK3MUKLH5fp/Nxd0L+g1khzLxjepLiLF9T8pGZHm
/6rJLO9+/5dfp95vmubFySe5REY+evpox6vJku17cHCmkrDkTVUbgmVf76oPi6BK
0BfKuXgu9dCzGxnwvWkmSV2VBCCEqr0K694raFpguY0/j0ATBlS66fYGoavy2xir
YaIcHCfl+GLFr4vzXtIgUd2p2HdN7CF4V+qpH6qzq898m1B7xta1ZJpxqWkRv1qi
XcSAPoeUdTSHE6XH2rdKeRJYxpuQHeF52V2DxMVeH/vUa/6dFGEBuRLJP+jKioJw
crkJ++aFQMYpuHqxzSkm5KkQqe0sVriKoYK43ZvNHytAl/WqCWFrfzSkIIT19Ai0
bY2diZpvD/wnoM6lxWaIXHWuYJvqYDpyFvvZnJ90NEU3c3EWWvivbYOsOZL5S1EQ
HQwtDF2cP/8gRQxkiK7rPAc381QlE24GJ2OBU2EfdwaAY2A/eufZI4RIUr5g8fs4
hm3SGNl7AA1PKM3b2xztSI/N/htAb1Yw4KA3tx6g/9Xk6SoS1vgbiJppYEH9S4GH
RmmYkdnabtO+VKb7vO7TvD8PW5JrDR6CjsN04TPRi81c3jxcQKVo+FVw899ICHz4
pm91xv/cIBrdO1ziUOq9zDyxIphZyqjWqatYMGlls5ySDPQ9H/hb6vrWobMQDZOy
X4bGHq8Onl3hJgzQaj21AQ2tRdR4AhiePc1FLZoUhVTD69Op69jI77R0MZaO4Cpe
DRkJf6TCcT6A+qBrVHJu/0EgWMlYJkeZkMD79JPHhZ4YN2wz6hV3UYohvTlckuGY
gdk4a31qTq/2Cp0cHvBcpk89bNeedxc9NDuMZ7mF3vKRsmVaWOteoxEAEnnCGZkT
8VM8s/dlXazrQHyhV+WJEjqZR//cN8A7ZjNMhfg3ehsDqQvWa9BDoTv4Vp57IQb9
vdh8tnmablcBkcGSsaAaLzzV/hgHofPgwxvY9ryZ/j6aVgOjPxAZM0wF5vs0RopN
KfivxwUyaxhVvin0FFl3+MTwnwztlDFbftnp/Y5ff4o08uMQ3Ukb8OugN6hnpeHZ
WLxpzrbJiZYrKR2ubPo4SzD1W5upkVPqGypdwyJZPs+jYdoKTL/V/GPdw8Efpr/L
qqf/RBck8RKqtOuxOQJh0/lI6H+OiXfPkGssZgq+izem8uni2LXuNUxx7igDZVZ4
4WhgH4vQ1uE1uMZXRh8dYENTHRLoLyM2hZLJn/6cNoLgoFEcX6Z4GydA30aSVymO
IAA2orgySThHFjZhUPmAyHQNWMUUpwLDmeB8WA0GBIzqsbqPJn4OzbaYORpmWRC5
5YaVWm9NOppwXpQlL+7KsmT1kQ3/GvRVfuWA3Mn+Qw/I1RYeHOdT6JG7lDg/irZk
MhQGKbSVNcXhDLUV8DP7hKjBaUXScXUgoARP7ms26+WWs2U946QQymLvA2HFa/ho
XA3+fc55jI2QyzJv2helwGcs+gPPuzJz7RZehNOBTbRbUTKJ5M7u6B4N66/En4wi
tgaRy6vOUmfvEq4e4MYBHTeCdW4+5+NohCNtj19+0Yh3tx6Xulj6DY3L93GvKMiA
BczqBU2vmcYdFhPp3mfB8YXpmM8QtErHr2otj21hWpuOamHn7aI6+HvhyZcCW8f5
zP0FCDstvgC+BXClqyxbwXuASDIQJ2vfVz+R6Ys0ZmRyz+X/R9sTQdHYnven/zBe
BFdb4GbRI7wwr2RjvB/nMcQrWnGG/BsfuK7szDoBzZzxGEr/V31TpTuyzlf5S+NG
xr/kslZG6WOqMZCP9z7Ma13/ziDSVKIT2DOWzp9BOG8L4Liuw0ChtiV848/iSdZs
05QXJZPtXryPHwFRMHeHKGGLquTk16Ux9zp/+SHowWq/E8o4eZBdoojUQUWiHVlo
V9znJrZLWpIfm50nKBmBYpooteOIaJ99tQpp0MFpJmSRsD8Vua/v9zjl6H04ZxR8
xZwoTTb4EJTGNrqL7ngkeSLoF1OdbFXv+WO+Z1kebll7IoCAEhh1y/bA48d+5D5L
hGGhj9HtTqIDUhoQkcumWrgt+r8arBnjo8PR0oajn2edTDwnWXNe6W8xXtLxXXON
2YBc8QLIRHVDKAC5OhORfQaRoH3sHs+DpgXGT9gKk3ahkhKwSNJWjRdhOLDRRv8u
CvuG0alNkNg9VfaJKv6Zzg+42G0Bpy1gh1KbWQaRMgCoFnleI90UDoH4XM5CzcVd
OCtI47iG8FN07XFxgNhNV9TitUjX5JUbrF+0niaNUueKejaEqdHeLXUsvq7OKGuc
cNtLnf4r+Y78IE4m4KaU/GBLaclHQA+9hTlsMrmvHOIMR9nVG5icycuQOCxvjgg3
Wd8jNGJ0biVmPF7XjMd6CUDFuCIspTR1K4OV414vXkbZhtjCk3hs8amMalEsm7vV
9CC3qDvjQC2B/dZMl4eSWN3dLi1urvY9KWjS0jrkoAssdoYcCYDAbBZTm78CeqH4
uo8IvyJ5u+csRuFon+UAkq4j3e0b+6bb0+B9rbvPPWqRpx+5MioWnBOd1drSUzv6
+1Q+2GqqfQJWQZ8X9LS7BOTi7w6D0qrsmTKx/hdAiBrJDwIwEePOe09F4qbMugCi
1S7EltX+F4aFON90TiqmQ4ghQvqKP05jpuzavz4ACVabOyz47MD5A3K9NbkYwHHS
y+2DGXJw4iVftyRdB0yPMFYvu+L4t4grw+BbdmGW54Jq7Wl4YMozeci8kxOl4VT9
bp8xOYspmxf46/g3MalFt/gSraW1ByxSYaDcHa4rYl8Hp5JZp/O+aILZMx73UAtD
4p/iNDlp7feXMp9kHP/njPxn1jfa4PFgS7snDHVusq6PTPVf/3YiVI+T6zvpdlzi
ehsmKs/yCoWlfLifPI/83QuUU/GNqZe4eUhKtAz1ERFQh7/2lwX970W8mkXUJuwa
/wxJQrdA/44N9NjG2rMWGxNChuyyeBvEXvZXKVebvHlJOzbhdjxJiL0l2WNy6zdQ
nuDVkhtVl1G+/ARbc/wgT4y0PLTn05kUz8WAKPUWYa0aGWL3vkpheATdS8unjqtt
PhMO+pJ/WYNVqJ8wdzpBh3Tu/ugHa3rqB2vR1k9pNpB0Lxj3nX5Br+LXsaWy04cX
p9y0J882hOdbvCoe6i7PwiGTONUbo66P3CGq20QL6P5EqFLVqZB42Z1kVjUbFg8B
swRPZEeyKV1fLE3RET+6dtXn6IdH712zUrWnGHX45tGXlw8YaAPBnm3JBh9M/3eD
kurOXQEyamT2fZsb8cyua3A7idz/XgaTIei6lvcZcOmStTfYIOn/RG8cG7szDFnj
1wYjh19tzYEL3T9ttuLjnDbx0lUOoUKTvGDJN91BYScW4bAtbY8T682nm5q8ti9H
WpjdKaGdJjhJXFNx7yEeNDOSVF0uypyOEw0Izo+7kjZeZSiM0GKnUudq113UJxVz
+3pCD/AZh1hUIvs0BorT5TWONg6JwagprZ1WSmBl2tDO5Ytr6BCvk+SbTlq60RYQ
w+fzADMi3dG0NNr9Si7qHL+4dCES4HO0hTxetadpY3HqExGwLSENSLm6Bgg7+v6h
vpEM+nApb0PAiU20hm1t8CxGIbPrha9VhZsEuLoUuA4qkUux+0dTzacVnphIXNHg
Fe5JK3VYoBvdTPqQf5SFGNnDuOlXfvGTUqWAULDTsTiKiDHtsdZB32hw7i3iTi/T
zui0tBoeMi83C7zEhhwr/Q6S48a8s4toa0aoSQ0eO7u97YJaK4xqmSR38+wbG9lp
66KrMTFi3gQSgZpBkIHE2IGxF5lGOlQ7occqg703+007kmexwDvC44SVadqRGrd1
x7jL9GxCg+0OR8ayUPHiPGk0bw0k1AaQEhLYveZK3WdxWiIaviXKY1jMSH/mLbV8
bJb/EyFvSWPLrIYccsxC2lE5i2Iv7S3JPpHCRU5IU+zHXeHdLdcoF3uIzisQeKvr
aaV1uhfkWmjAkgb3Bgn2t6jf5D+8cjUS/BmrQoZ7VUTS2ZCyPkdin9/TzWBUbxw7
4oU2tJ4ObC2yioNY3HhURdZizS3pANPasVC9cHm+VhabC/uipeW29GiTbexgdWI/
cBkyD/7xR1IlIIPPOx/0/nhA0l3a5uyXjleft1ZwHfdf6WrliYfaNsanphqKBCUU
hQxbyf9MlQyjYJUeCgt6iVC34NtHtN9jQudcXmYVge1ZLbRvmqdL5XiKjizkjb+q
N12ITmue727Ezi6yQKplfO1USzz4puVIEUDGJvhcPIW+XppMi2V8ShLnlr2tMe6z
u88I5TaqP//xTNo+DKFvHuU1asZudsxgXXkvQVphMfkaKegzv0llvWzQQBKxTXCK
pTthrjRinE/1pxMtUPl/qyysGaolp+qH7cc5KWRQ6vUyjyNjQZFqHgCVZJheRqKq
JJy7rqJUGN3ZE/LMq97+SBxAwSDyozjAikJn1tTdhOwm9uOJ9YcSxqcc3JeIyKAf
XME58PM+QCMSNOEWDD0jn09URZk9tMG2Zv8B9on9LE5u+peU4HzR5qJBh4yO0jgp
XqI+mzAno6UuMi08EaZ+/OiNsRcFRNBTP3/1VaHy2XwJHR53WDCdBXK3hS85eT+V
+nvwhDPM8M6MRx5/jFrH4W0F3ON+kNqQMN9+/XT+t7WvabkXr2pfmhbkHAufTAsk
6/r+QmkL8Ab6eVw5HI2iUb9K+GW8Zcxz/pHSfTdPo/wItRztv2pqUVVHg56xT0V7
AYpEytG95ofb6LZ1wJNC8/qT8o1dKGaCTZ/ZD44jF55Vm/cerwzAOApaq66mkfT5
Ti3KbzLoXoeXjEhmvpi4VXiwL8bf6QfaUkMahKS9E0eX4y2BHXs7WB7cQiGC7tvc
kUWj+vDQrbjgbjvwcG3AsfZjwth+AFZEgnkxT1NU/clKjD/YpH8t7CkeHOp8Pf1n
ABpGOBklZ3LyDV/VSX6EeRbiXOpl93AF6sIJlZkQX5ZipZZN2HEmiTC1OHcbgReF
jRfsrm4yUVtLY6Od94vR1EUO++zGd8fIqpdSVX3uNxQ/NsavRnDpuYvfXhxk73ny
bKzApaLrCCrHlsxigsx18aMnT3TwgPu6YLFW2/9RJzQnS1l0lGSwITovEyJzbjtI
VqSK8PNUEYk4SZiSJW1FG5zl4x6wn/TyW0L426oMwl2hOxLnGIpaGk79tUpODSVy
rva38vj9dWeC6GfUs1cM2qct2rV1t+vgpQrdn0bUdd+BRlM+dFtBCwYakTEUDz0e
w2M3llFnarnfwmienTWDpQUYnawPqRXH1QuvDj1p6IxAiFaiufXwSeXaUHHELHV1
HjB+fyPomMi+ulJKSvkpuW3pjdO3kTXlnp1kxS88qipp9aTLjdF+8GlFM2eU8YKl
WY8DcOSI0GPGynlxjlo88c7YcvaQPGLQfKW4uzApgZ8o965TBo0GvP/K9k02jsgH
V5anNjZzNSRk5aZng1BhQAhAH59e8mEo2bGLIzxdUbsbOp0gQKj+wwoSkWdWXntw
mPKo+7shmhgtM3kl3QZNYUa6CVIoqjKg/3rxEsVUW8Ykr/t6k5bQvkVRx0yMNJXn
hOC7GqZX4sF3drjn9momrpTz48LSp/5uazF4Wc1/Io1JBcZl76lXS0AFoYDPsQh4
V5pqdauSJlSa+iytU4QFKy0Bmo4C353gQbvLgijP+p1pSqRKKGQwEJH53qmnuBn5
XLSjpgqG36abxuMj8yYIj8zdhc57AX7cuW5JiRTZ0LpO+wG6z8bzyl3CUElzc5wk
Mnn/v5sRmm7Zb2+FG02VF6OgeSpyra9eHU60DBDziU/cZLTiGQ++UoifSkujiGif
kAphwsKazqIeZD8+7ZmZpLQTtGJoQILissmbCwo2FvEOCUr6a9n0Hs5yhzvTdXF2
2r6g6KnrRzmud8ynStSaR7b3RzSKLZhHz2a1StzWaRZPEKxu2/mr6srXCrtduKHx
UxYQjgITr8WcNgMmck18l4ZHLlaCwX4nEwj4ZmZad6OLDxKXTGrc0bckZ5L24VfU
hi40qwfLLWzZZI/8HinMGrxn0G0ySYiEI+rJaBKysJ66zKINxrE2Isl+hyM5HlJS
kfE4yhw/6/MtU+x4Zn50oOscmDgKwCAZm6E+zYYDWnBeQt/vbeuEJr5nKF76ZVOT
xjBHbm1Luvo4xQL5ri2iyqa7CbfvZt+cY6Aj1nseizFd0OcXV762tF5LVkYfegSB
NF96EKvrdO9Kyn8uq/y8no4WycqtL03WQpfiQ8AoEhfROZX649U7zoPsES8hFpr8
f++7ykgZ4Xd3vH7MhSXw7pm+qu8fdmHO74Kv3f3skAvNNGNN9Ek66aJbhwfX5hFd
c8+1OQfNIGDW5ToghZ2no19QDZbw6nvSovOxlzKpjRVaTIBZ4pMBT0FRsMSHMfqo
NjK/aZ1U+8VW8tbT5HVTCpo2pmLaS80Ubwz7ecoajwJTYJ5vjDVji7/slnTh+/OT
Xfp/Ts1gYSxWUuZiWtmpW0Z9m9PpwqoFk4YHRFR2D4md3rX1LNq22nVJFnvGfJ+v
2FJbCzv/1ImpkIEwdQy+jKi+B0i2s90OqqyHNwVXl+33tYuZBcRyBomgq6vHQQ2j
ywcVTR3j9A3NggM+yZQzBZD3N/88UNKOSMdY1BE46WKP6uyYaNCyqC83/e9xcWuh
aKpu6b4wPl9kdVG65Ak5abggLTKahACX/lUfylIFCnPf/kYasqJHQMfyfAo+7W68
4vwyfKqB9Nx9xZR1BQjyTPEAypuFSiCJPkOKQCwq0q7c7ZtGFLi0R+6328Ztqqfl
84yHvt2nMa6OUivShFPcE5LkSS3uv1mR/TGfKOkYodE3R7k1hZLRGgVDupTNjue5
WIVybtgpIQoWGWitw0Op6f5n5irhGCb3QUC8GtIppP8dgSFk2Nqffny+VkmPF0SX
w3UOV+XfT7v9nLBmNxh4ON/9lQ13iEERIZKLN90PmZ2F6SSvmXwM52vkLYN53tyi
VWYS+q7B7Dss5XzG9Rz5OCMLDxfL/3hiIQpv0P0nXnuu0e4qYBnNCmLgFUi2QL3U
ksokjF6Z5g1ZkocIIwqB10CzveL8b8JJwEW3Cq/SjDt6MtvQ/A+QmjpqffX6d9QB
kCN+Z231pQoSqVDz9DZw5iZj8x+Nh7vhKCGxEcz2NadIR0Y7vcy1p6NCFrlU9fYh
YMPK5czMMMSWXaAmAvGzl6uJo+lcLqMcGMQ6OynVAz1/vsUU3pcq6kuV/HbyQJr8
2t4GPIicryhB0+SysicIXoeos37Wl1D2dtxsqEZoCMJ5UqXYBztpcvomSX7y64Xu
ND+HlKpJA5su09dFQ/4GJC+FBENvoKZmX/BH0GmdwO2Hul2ohur2S0ms+jBIoF63
LHSMG5+pTaoW6t/agNgPTQWHV0ydHzcgQZ5sVF/dbiMvl193eUi9+nINuPEt0NYJ
2GG1+IvsENjwXwVdt0MVw54l1EQU1OLchlNnFf6il8+eUIrXWE9qEdLYqnB7/Vxy
YbhowaSAQiM61Uqt/WeYpXcEzi3rAzzL4aCW/8AbQpCXoOYb2NOYwXhxKGf2bflX
mDGdz0c9ZnQ7kUcfpLkA/6Vw50f9ZNyXbeBYtu91yEmEMlnv+Q6g8th0N3VnEOqR
mKDppqaT10o5qa2G/ESQqebt5COIH9ZLPEK4a55kBtChG18VDOwqs/2f/U4oNnEq
43DC4+8wg4eQfqBjzSS/yvf8+7X1p7hMGga13oPygoVoydeFk4GUAccn7cKtqv8V
uwqTeEOIPdm6j9FL3fZPksm35HMk73FA7l+OQknn6U10MpVULC/bMVWqLWNEGOIV
blMH9pdP6qzSgjooPNgzBg0MR5t2HMVqv3eLxvTMyyY2v7LUFPqI812veQdlcfuO
z0X18NC6/rrXxnlwMNUDk6FbgWvpim+f01TPvyzo039MHh21XUAft3TwQGewCWeL
U4UTMk6397yndBuLZY9gd94Bge0bFuYgemrVpcfXxQgmnz8p0iV/UOvaORmy0s3y
y76KKhiy6wvKHVfvJvRCux/tMTi0nw+6klW5dBKcsD2NCUV9Q+hcoI5ikNL8061J
6gGdjkLmhvHsn+6GjdVmYbK5zxaqSWNz2Xxs6bIHZV+GCu4I7g0gdlCC8OeSqDO6
SZjmpn1pBEsEzG461miJbCSIL4YdQ+/aenXEsJUr5Gjo9zoQPYUb0TXqpwgcWljn
5VDyIZaATRtEclhs2zU5/to9ATs3/OnMrVImL4YcjquWgD9Ii3aBcsqMKtvNV6by
MHRzI28vPLnKmVe2fCQWl8Uu6zId/0s7FoypI66uDJKPHQk6thAaT05P2hSs1NaX
cx1r2o2zFRDGb2l954iO9+vpQvItiBa0uqcZ9iZfZOU0Uvr5z0m9CujEOg+hXhTk
7wP/A+hnpvOE3htcfQ5p7j/P4wfQL7AWlJQ5H9+UkWRmiVX3wDWKYgK4aiKjwAKm
VGOAWhyA87ByMGL1yA7zCuHO42wNMQddZcJ74kG3HF1ST/9bNkxvebsXZra7Zens
2a77lAGZ9u1IUUw52/fPR9RRjlD/6W4FqSZe0OuRNhernsstGVtUSwDtANMRC7cF
Kj+0zwzHLYKzqyLFCbMRWUbp7UAFfMfRe5wQGKFwrtOX7HD7ubYX2eIxSZvOV1Ie
Sd/NLGzu3886dCr8Voln+KOhAwSUG4otAmYxbbfcmCZX7q1FnFyaci/zZaCrxA5j
2t6fIJwI+fgofUCIJtWzhdN9jc7YSAauq/wtxW728S46h1Pg1sbLoOgOfIcNd//M
SVupOk9PmvFRZ1pzoBM7zSWqeLG3S95rAvUzb9Yd0vF/HoPmgGSPY7QV5F4wXvuh
BND90N7adu1kn9tT43htAIVi0LxG84QkcToo+q3rY7BMCrobaiXmyzOTQhhaDjIi
dUObDR4Cl+vvGix6kzSyNuEYhwY+oIccoTjQvBbE0XjrvfRdTybbvzww8Zr/SEEP
lLx7GWHvgUBjtXGyFTNNh4XLyLq7louugx6+4Mq26O7Xh/yudtKpVWVkDkk+xhQW
VbY2mZ/w2p2RGgk4wxk5znRUDyL95Uzt8SwEdIbObSeDKClrG/3ma5zuxQz3zcP/
V4ANKUR8vfLwFVL0hbbIYBMbVQNkanO+rovIPq9cGL7b7JsXXKYeLFSoM2MHLv4W
vCIiqhlqRxDUd/8nh+2qvItX2h9HEf73aTsu1XkUm6FdqeGpdy2EBFc1oZuvx1s6
3UtW0I56OvipIJzWBV4f0SF3IjUkDD+CMEksOAjXXc3WTVMe0ezEW/6kMzO9kFd+
inFKsjhm87WSvCILIMSUFWo7TivOFFRAJP7CTjRMElpL4GAZmxG9u6Qmp3+/IHVh
p+AXi6KBJq9NqW3xsScFTT2IVteaHqTmA2Aw/iMfY3wWNC4Lo3DQgFBLAb5Yu9s/
hmOFaELeJe3GoKZ4b/CvXfADr8RuetH2pci0g1GFnKaMQk+uT3xYzlqgVmeASBi8
C+ddQery8wm+CxlZfeGcYxLw95zui108XUlhgW0umkWX8Dp1n2s2NGrSy07fyl1O
xIo3wog+zmMCfS7FqqCTiY2u3yYACJpQlW2Bw1KMyxp5htUadGppleNYWeAOPkdo
iFEU4vHVd46GxTEZ4NP2OJ3jsEmCHtBhdOieJMPaBKIa0S5WcOqw51CIuWAc/SBZ
yEkBrjklf7HnlOmGzJ5F4PHKEPSJMLqfJyYwgdSwumU2X/MDDn4OrTg+5LuEm5vP
Ydv+vrtXCRQCtpkX6T0zhD4MViqowcKJqLcIKIWKp7GJTGoTgaiNwMtjAo6u/c96
IBIzpNMKrI7wd+BxDnqWuuj5E/6HrHoY5FLpC9+FcjohqgzRLZ13EUnYLXyjDsGT
311kB2DvWxnajB49PfeQ1dER/roJXTKGhWedPkH1FxHTYVAMiqzfiXJ3gIbtuvSk
KvA7alIlzCgU5pKN0RtgIUoWVSIeGYTPc4qD3QyvGXUO95F0O0hp9ioo3aO06mmR
J3O4aLEmN9fQICkH7QubsJynT0SdsnBtgsGas+40vzV4iPaGJiKT9RT3zo+shH/N
wQzn7v0TpJw/H/WWsTrQYTpqHLUyQzSvKxZSBbDlVbm8Fr48RGlmESZxyv2D/vUT
S6q/En9bGuemqWCI8d3JXJRocSQIvbEIddHDRNx6NeadiAi71keGoW/Z7Pt/g+kD
yRKiN2KGwmShwdWmbbl6m8L11rs0FunT+RVVNgdr52a9ZYeFuyCwO7ptl5z+TEYC
jFkKe7MTScdoV51AkFNrP7Kl4+H8imlBYSOIj5y9YTc1xP6fOnhNcwp/qSh8runC
Er7UgRD34ru0PupHP7PnoTRDDcL+xGl5wmQE++t36Mh5th8PsdZcVp4ONa8slIIx
xK09rmYfbIhI9SJQAirN+9Y7GItUwC6nZxI7MQPlkqQNHPlCm8kFbCVEobSrc4mF
kG7g1DEmYXH/lGvDcpeYT8mmpBCOkdHmz+B/ewsoXLfKqJNtsluwm3NkjbHi3oFY
C2o2HJgbx0dyTyMXYot9CyF9Q7CVFURA29tqxHPHP0pooFmpcCufw7rHTPWvpKw2
Lpzkv2sH20y/eRvyLdaCKgTyjYUNKuTPnjRQ5cXBB/qxbrEmHB5n1U94C7MGBY5K
/uqdKTT2328Eq7yW4FY3AW7ynp/+t/MnxUzy40Qx+1ddSL8iQWqGmfmGaeKNBw6J

`pragma protect end_protected
