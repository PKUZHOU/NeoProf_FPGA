`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
oGqIiR86GTn9ZVEbvxL9mz+pkhpHxXOOdVCc50S/17uiSXvkE1iMrqPfrw4TXltN
AyB7CnrV4BWLoBBb41vnhGN/XeB+2Y0ufeCI/nClUZqcYt32H5X2zyWpmVgu2Fpo
EzSbCDPt/TtkxtqZ6/TggI71P9pCHexkig2ENUDp8rQ=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 7488), data_block
vIEESIWgVSzAlQ/W4n6B1Spef+AnDa+WeuBbFPMQ6MFBkASRMw04kbbnYE0AZ+uH
4LFqvRIeeCQ8IKWzvSmsw1ucqwRwSMh0l98yCoX+GlOPzcUu78bRBepd0bNcVfv4
LVg11ZOh+gEOvxWW5p7n9A4UYWusVWdtvHR//x58h0ot33356b2ivoKRuXocL6VJ
BL0nud/I4HJtTS0lvP7ZWStN8GXBFmWQCiRDFXYFoS66uvSq428HoTXMAu++nMpY
vE3rsstdcMC6PqdZNSBTVbogMlkho2VlGEXbYiJS5CBAfPoGzaLPr2HO0yuQ591s
tVi/nqsvCQubirwFJK7mdoB1EasZW4pCFgWZ7k2JIW4Xk+ScD7SErd1Y8lWKGaqi
VKIZBVjJsPJAdBTJK0kIXq071qMKuc3iyJzLjOCWIoUtrizQ5WKAzW24HCi8+miX
gsYmnsEPcWt64ujyjAjvFD7I/fQZro54q2ktvbE1Ag7Jf0Zoqqvix3VGI2S6UHYh
RSwiLgGw6tZqNsGfizWDWx0SV0SntAY9d1RDjEiVVK6Pm8M4UVn+vwF1QQ7beVfX
TlBBiHHSE3G/34hPvHdZA2yiUItiGwMx/NhVA91e2xAQLYYPsXFPQmDNtUyKWOmX
cTU1z7wmOD/MGEyM+HYOZDMcBjcM+dlMf4PQTXI9Ro9vN2Pr2pOIN/riypec5A0J
LIfmbz4AlUILD8ZG16Vq3r8jQHaAJ70oSAS7v43Aou/SyK10olAdQnu5io2gFmhn
zmRtVq3HG2hB02Z5yp/q8fHYnm48FbX+phkSlSqvR1dYVU+I2KmO/4M48HtD3bzT
nSqTcnMkTGwh2bXPoI+dmziCWFiugv33rKSj7YuHz3YCKoaWyFPy4hQ7W/jLf6Bi
w/+KFrZeL+ZSPKz+hsgXArv8ou18DHtICIw/T0zX2Ypww4rWqUbrZnOP/BY2DoPj
c6Ay82JZ18y34zCRCtwWmEoTls4zoYWY4BD7tr0rVBQAL0i6Imdv5gS0CybzoViH
WW3+KVWalRHBFb4O+j+oqL4twkJLUNi4CFxvPiybNoKSh8bl1YmaKDv5oqfhfgZv
X1YHmR3Ppx5LEveUqSPjDz1YmH9NivXL1t9f3rivfCvXh8f4s/SE69Jk0TocaYXK
7GP8U05CNM0NFpm3Mq//R+xFDazcYwdrAqR6Owa43fOcJQrRLphv87vBgwyiEBha
uAuKg1V9CCKybqQtclDHELoxKHLwvVZ2sXm2MWMlYKQdwMnEujHHBRy8T5k6Z+cg
Z3iTZ9ZlH2M+RmPu78PR86Lqp7l3wnSEKIeUEfOY0d0iYQjZQXcRbrs06DQSMryA
DXXLJUGzbNQ00zXNrSL4VT/PykwANkjvatCiRhtC/2XOrWjWw+ZgYEYDlmEDpgpz
h4qPt9/b0k/1aEGSlXe+Y+uYyS1r2bKZx9Daqevv0ZO99c2/OZoro/F8e0Y5uhbL
55xOAVUoNQyWi3+OvV555l+e5gwGJZ3hMspNf3iBofg+Yd3V0jJF6dmnBrzZVHbK
W8Wpf/vs0xRinTkry38Ekkv/Zy8poQI38m0yMsxh7ln+VoKv+KbuW1meOdDGsNke
HbET23AFeFo8XLU1Uya4636IZpvRytcSsv9rM/Vfk9c4960+sR7NsktSVaEeN1GR
RL48Nlkf1Ca6GqqebK/g63cm56f9GotyApU0tCOjEWIZpyaVi1qcrPCY7R/NcgMy
/H/unEDs8J64gDBS81E5cnT4RbsNsVMGnUuoSojUDYG7MU9c3h3v47AD9OexhBa0
JCWaQprXZxOF9JzJtvf0FhKMMwqmBsQxBCe7suGObueV58VQwGfPBtVSqnnfdyrE
LbiaUTF681eK9+cuvD1kwjwF3/FFJqQJiAv/x1hUEPGAJuGX9LVMcLZhNo1hd9iu
sfaTz2DKJrwNwMIGFMFR6KDg/qpRGtyU/ELx0VBvxC8W0X2xi+sOyRfgK/9X81Yf
0GXOuWUWyO8gsIJ6q4k56dGDSh3MCKz56+lmYa4j0sxI1eAeUQxuwT6FK7C7LMfc
VihWOxE04144434OnJMNkqa1bzDKZTFBISXnOQY0WPcI3v9ALGa/3PbpaEGaorrA
I3n+WH5jkoDOtpTQxClYfHCEMWCv3HxrpmUcHcAZBoyMAgnEmzxW0vlHBAj9g+M9
Iss0jNO2MEcgU3xMt4qJdK6MlMwsAGA4qyX1oO4lGwkS6sdyN88Rm1qnWXDuJcqR
B/uA6L/IX92mon4feTXpqYkz6yTJ8ppIUmhexpJtOTpNSGzGCtawjaPEwX2CDCiX
BMbE3tQYTxZJE6VLxG2Uek03WsKJIFi+4geqsW+iFjzGIbdPHp+ci7mZ/pLlS6VB
MO1zuJHTse02zwkf+GrRQfXGlAQqm2X2T/wWE9/eYYAXavO5a8NapmfAlkpZGxRW
OWJO8gciYp42Nf6yM5MbL64FHAt7RBdcqJQFnfG3pRWzlNFHlgYBcu0a/HlD4WFe
/bMcDVASlFk0YzNhRYdWu+8Bol02+ESDQ3m3Lhu3ofnRZ8rDg6IPrbAwfdjl1AqO
/eNb5ZW1EaBlY2RejkW5ZL++A6XqpRhUUDQ8B+odNY1Zg1Pac1Xkiijs9PsRxevu
0/y8NJqImddWy1NOonftA5apOSMBm8XxB1nDX/fCKh3Sm7T8SlKkq5bG18lBBW6j
/rAG7Mhiyqd8losWAS0rPSnN2WBsSIWKi1kZqaTrW6lrGwuIenV8mxDPdi2VI42u
vitNT455lQIidtW0gpFsgMaOq98gjQxifErf2un2kESjWU5bK4z7TyTFaCDp0ChV
7MMCq4EbtNMT+1ksnXqC4j9zXbzfYCEHHhSa4dRWsR6vquioEMfXNkivP8xM+B9E
hZexlQoPeFpR5xh8pOor3SHCExn5+uvYS2tIc1nFRuWZ4qdiBll2JDF50DaNHnwE
awlCmEZur5EXFVm+YhDOHF/Q6AO8DbDR3hQB4rDmLpl0NLcIeFAbFWrxk84f5xcD
sr7N1t8lbcVlgv1ILoL3b2KGuBt9ntwlmaBfoMey9nuo1rbOuKupYhYiEbDizNuc
YhgVgaEe9oDbxU+9dfQVaXmPk5GyJeDScLxmJrUGZg7hyb6fJZNUW2tCaSO84HS1
0tv2rutAdtms9eNubBfzC/bbMnI6hZHgvTDeBVL6jkGY2jaJY+GDEUWffUOn2cOC
vTZZwlgVKGM/MfdMX5dvawBNTbRIo6O74+RUZ/f6ioyMx2cGM60Bbn3PvmNMfclk
ihbCrS2JdRRowllMPI90ryHfArQ9V68KLfaEhJrnuo9QK1VXiNMkgbnpOC4n2kzY
Puup12uUDxKDN1vKTqLVCmrZ8ipwyfSTJOJIcT40cP8s//fBUEi8pcGIH5EDcAct
R9WPCd+hr0D0JsJMb3bd3+gbA/oUMPoEkX+4NZVy6QGTR2ZC/wPv3DnaewFaF7FW
u6XStQ/WlP/DMU2qbcQ1FJAead6g64R12loPbNuuZLBql9Tq2SmLPDKbhzpcNwG1
FbhO8eJf9Nvgr70Ki/4pxXXkCQTPiO2iCO8wksqyRx9Jqy8C0K9UVwACZbJmPz5O
v7bOwnHA1FZHqIcGmMChmGo2g2SNMcNHt5PlHPeImz1fTCNqWeytlTILpwHVn8Nd
TM0sOM5HF0IjN35YBD6QJPCog5RIeid89dnHcjHa0Qf01DqQyjt4c/WKprIsnjUP
70l3C5Wfommg9pnclpdyPwU3khUlwJJqfNQ/kvQ758GIITXhnIRPH6ixPc/7XS/f
7W3VXElfh4Zd1GCpEOZvp6eG8d12CV+6+X2bFq1Im2NppTuwIp0a138UO2MUt0aX
m7+YIQDgjWxGk+eA41zAhNjxvnA5c9MQbWJNPHb0aYteYLYm+yoMesX3GW24rEZe
VqsJT7GBu0twKxhOHVnuhYxJhDPY8MelYE4pXtKpFs+CtTkOPD+rXpeo1eEMJNZZ
RLu3F6WHUadOlK4z8NcL45akYyMPmAE/q+/BDCCG39OemPC8GHggo2BvfQ/jn5ln
fX/OX7w9UAUL5c2KXEtbXQiqqfv6qZWCsHVrDpPx8HgDF8Qs90jEOycWutTxyi/4
7KmLaKFr945fMHWpbzhe0VSm2kHu/ZskejI3bmZWi4rRUkbPh/D01EKD3f5szA1y
RHS91G1gmjzcPChANDDXCvo8VukQV2XDTbsYfdpin96LUQqRZnE7gGxmNJWmAmjG
Zt/JO3idfTTul8QdDnJOWnvt5DY1MqG+GFdHcQVl0WMqZvQU9Agme5fukmwt00AL
4WUBoO3rThDzUy3aCWXjh29QMh7h8b7Vbhs78gUp/ZKBDwwrrZZ7o2C2iWnHMJ7D
NQkiqndU0k6OdqabdNTgJJMn7Co3VnQH7jkeq0895M2fbVutH/DB6CNxQkowGddX
AapjykAwz+IQkcOAlXntygCVFZkQ3sF8/3EnAGX9o3H5s3duzrd66xHLoQHzAw3k
u+H3ruJmw13lmJCPuI6yetnC3t/WXxcMwAjBU4wvTHkj9ztH6lPmpU5y6ddIXvpl
yWvMKI3FodypxW//8/jr0tkgb6X57SbS5LMZtrO7B/oemjTcWTmpO7pcUK5shHTS
kI0fzEPlQrng9AA9npAYOKyzA+cYLo+zeNjUZSe5xSUKeDYS9vj/FSiJafM7JNk3
mkVU7mrGC1Ikqys6lEvGRVE6p+BFwpsvhKEa9hTQBQ+LRESNUZVFFvGnWwxB3eJW
jfZeeVVS2BtIK9nGp1yUADL9MfXa15LF/OyDzf3IIlwV66HkzlBLpxJt2G8jaUow
iBnQTjpRWyDmLUCVDWkKMXU1cqbAnRIHO20QFQXEDTAOrph0b9tngjQ3bTySIQls
/CmliriPB4ab3fnnZA3rDJhsSe8DEwIrmU3iH83ilt2SOWwbwBm9nd8EaulN8bUj
HGHaPmqvPweAm79QgwBUkC6geYAcAloUxdulVf2171O7m90HreiZQJ+jh3dzcIsM
ek1uqjdLRBEq8kd9tTGaGhIY4iF1LdhXu61HXvcUFS4jXrpG+2ZtUUXz3OA6uqFO
T+eBbDtywcjsFrEcyBjfSX+Mxp3u3WPd02nTtfY0AsCwreQ6Jud+G7hpi2t6qsJo
Z1cEeb/Il06IuQTglXyibmYzocJu2Kd2+Zi9IbAsE+YEiyWdGHyuL1NQn4O0rJGf
SSMuk8QtZlYYZ5b8zt44GMsDcrD1Qr1CHC8nKXaXGjUFFb/qeEhlM32NSY+cxQx9
wMmQrtoUydCWs57qX4sCHqPvu2BnQZIqU5Kw6JFxKsclwETQnrs3q7uk73iu/A7W
K81jBIyM0OCxEBOCce04Y78yXHVtxLbwS7Vn5GJ7QotFRrDxkRCufRYrRFPckSiu
Qtw80l/lHkLFcw1JQjB2C7PrWrS6/Lb7V2qvGx3LWILAFxb5W7oU+HnCtmftHE79
ckPpb013uu3qSaN5x97Rndq2IPDrCQ4Hp+Y2zm1VaSEBBaPf6A2tkAskELamsJQf
AZ13m6DXAPx/IsUjHtBt1CBX0fFrxtCFqJ9611RfwuVONid8wRYF6bejc20KsWc5
eyUVjXcOfUJS7CEbaM6DfujC93xgefq5+kzBhPQ+BB20HHy/XyTYIGkYD58QM3i+
JLFxmvzHZoVJB3mU5yYXn/ze9XvOjNKqngWrdUgWNHwM05GYXyckrbwOBconwPq7
CuSzeKwdLb/uHCGvwfaP/5b/W03nJaXntYeZNbqj6A6ieRwC+egNisqvB9cvJU7I
AjBCkanb1T7ks2zewHk9qGFHSe6ikZikzaMOsaTQ2QC/elgL5OpgzoZ7qpSXg9xK
4jvMA9MC2ctCZ0mdOHaJNn1LeB4yRGairM/xgWT29GEAwtRhS2Z7bC7ahrI4hpET
O1sEoax0C7JK7nx8XBMKcgxCnL02P4U25wMNF5sIijD7rshTnbTZm6Zk1Ksj+p2I
HIPbb1/WMdaCvv8g7mAUSWJlgdk/2VDvGHR09msTdVk2N7vTRYpYKwcCxeuRiK4X
UyU7IDYlmSAWcX1Gj76o1vjmOgY22d4qgHjdevkNX+4QGX7aDyQMko+RYEXFFMLg
RqDZ0xJgyqgaZkr/vAkMxvw1g8GkZ9GcG6ELlnqpZH0GlL0sKHSIIS1eDP0p/0GX
CTAwYO0OCCk46ZbGvCqWCj9caVPrunQ0oFNeh3Qvsh+Wu18V7azPzee3Trxbp8Xz
DkcUYPvbDQ8QOtL9Cb9OVA8cxVIjUnW1p0rwi2UynZLp+A7hGWggYIpPm+LGa5kA
wPrTb0Gq1OjH+uWEzNAVSl9e6JZ+mPTlDpq+AIEtUlDC7s6jKbFWRm5t/pWEqzmu
2H5x5cVvlb9ntNwUwzEaI0mUiAKePADIKfa3w0JBRdXVQlGlVpMWh1VbXHJIOJhB
3D7dCDYsnHUxkHtnrW4cmUzMDnY/oqtTLs9Cobu6OrwomA8eJexsEgGXuADRhSLG
ZgtVtB3B+ut/UXLbcglgRKzpIMLgBirXUNNWM80j6h/qhnBgWHa16DF/Seg4QDSu
Omf3fDa4liPbcpe8CYeedcbCvLviMUC/35Ek3oHM6iVPXTJTUIRzna7VgWlHyOeS
JAzQrkoZhlR956fRCbath63M3j6LaQRzM7413TmM6l+2ZaA1JjSoVAxyn0Cny+ol
4Hwec6Ha2TwDpzqM5mHi6na8Iu7501C4yOAtlrhQl+rJf2bHUYkPxOAOb9k5UgAh
jIsQMtBXWBivc76z+N3BgycvN0p+7ilNFW1KdkhgywgsUd1JKAZ56fDGQ0GkpwTb
vgvDC4dX0n4kGkCEMXPksz8RyYbWRIQXpGeAiC+24Gw8U/4k8HS3KGZo48GumIAI
o3UW45m6Zl752aI7JziAP6gqArrTFOFegTvx0qegWXx48HFhnp72RAmKJaFtyCBq
BZPutmpgaSHMrdRocirQu3L/7Muk1Jl7l8pVaAjH7zUTHOcb4Rjwz0t8H1s8fWks
Vlaqbj2GCm1+vVvNX5lRQAOUgBX4zyRoly7OuN0Y9ZV9DD4azKa9ISF+vadd4Z7d
PONSnH/ji0jb8d9pZjFdq5a34DWYZVXMvU/v3s5jORxah2BseQcP0jBC2khHhpR1
VoYJDoBY8bdUuhVbHC+eAvABlwduyF1qCdo5PdsuW9ypZXmSGwZ173PLjjvxTABW
qZtreF4po+ma+4VOXyrmSd0+S49uD1gkwB+QEd+v8mTvpX7Qd8Fwi6bj5puH+otV
Iy5+um8l2g1rIF6geNASzdBvSNBfhT7yBBue3dWAyOwu4u7BVcqnEOvXNzk7+4Wr
b76Jq1BVS3RdN/5gWqFh5ZVya7JpvvHSQPG/+Tu8P3l4/sWUP/qhSyMTu6R+9k+3
iUrLkn3WvR2Cu7J8b93IxuO/hU8Uhyff+w2Qi9fpQRkZykvPdTr1o4RBRiM0WdH/
B1xtQNpeCzhqT6jyVP7JH9K59uCaBuICDxAT4BJAbr4HSNCaiS4GhwSzblHqfs/T
tw7m1zqv0sAGkwO0zuRAPU+h2yAt5NmoQH002oVT8hn3wjeiBXbetpacWR4tSeij
Ka937H5J8VqEnklUOhTXre7NhiCA9HV9QDFn4n1f8f7WZ06t7vfIzgxoWXe0s+Qc
u3UwsXcuEdCAOW5SjZRgzmRRE6rIquYhJEuJigk0mQIf2/MRkTBaC4mn7ft4asFX
UW6DTSzGFjTJN11v4VlZ9f7kbJJVGMnPCfXU1UQABATHr2PUwDb6IKyd2ksxAXRS
lB8gfLZ/fsHhvopLwhfZb5vG0ntXQ+aGUaOz7CR5NTkrzJa9MJGpYpJSr6VxJ7xn
oHcX8nt1tO+C7EPskCF0E7UcmpQDndaBHb1aSrQADGh/0mW+jLkO3gkyC8Thwy27
aY5GCtR2x0oFS/Iq8G2IoVgpPRmUC3trmw47YmeFjp1JuBgOgmYxs6qCNgjiaqWW
DlMstrlLJ9AMMwZqYrZifOy9FTFK1IP4srAzhHsEUQRQA7zegO6BHbsCVr8eXnc9
U4NQ3Qf6tEG8YxxvswqLlktMxL8nLxYATyAE/sjgb3sTjvWitU1VF5oBoMD8m0+I
77jpaUJtHLLkBjD6yZCtNIUjnKCiQ8R1Ej7plnR4ESGMtUtVOGo4Y3uA8sP6Dkug
3acBvI7rzB1dzdx/cZTWthjnzSF4Y/uyRC85iBoPN5+5Np2jBVeksJxE/HSipWih
vpgRQyJ7inbizzMNOMhuTb0mBfqAW2XSzfJ7Z7tpR/zz1JLu8XmKU1iRTQaIj9IV
+n7QUnxWmpueEaNED9VWTXycMlCwnpMgOPXLt/mC+vUvYdpZp5FCSIcoAiV6ddrZ
tKSVA35xJeIO6F72IpcPTVsSGuaTb/5d0f4xzxDh/zFH27z69cy06mSbm7Dk3cA0
cX1yNExIqdsuWRjEfEUxn1CFpEncVeMSWuofhN2oPutOeDDMag3uMO2pooq06KLe
iGY2QgzxbvL06YXEmTC4M07ZQvCs6cdAoUti19AXygJlnu0MvTMMsVl+21A1z1z7
bH/pFxsiAfmoI+3Bqx2X49hkRIXNPv7dWhELg/Z79zrCLZSsJw+WRVvwRrX86WYt
juq3qZxNOmuP5LySr5kDRX9smwVrnPjs/N7a3MHQJ/oncTPt9IxPcjRWVM6F4Bk2
WCoLo9MoKbXmwNCI7+E5my5dVHuLYuNUI8D+zvmtbFn667LrSrhr2+ihepiEjFGW
IMnDSOgG0IVVY7H99qs8/Foc4yUH2IWDq4RJCibf2M4qzpvhq6+1gr4Rai1xfsl3
xALM60I9kcQNwNUqU/Y2ZB/GZpr2mrAOwGPy+pxo8hxrgOqQ+UBahyWGYisnFuTa
WuhNjsAAtVUMRmWYGCMcPUuFP/24a5ctm1VHYj9ThLDgjIusHADf2adElUP4E96r
xaO/V8kIbD1uLhn4qSM9yeMmi9O8O91DCBRxSjyO3fKf8CrhbQbXR4AtRZKkKu52
jRZP5nZSQldNGRpwIie5lrhp9ILZafTG3ddsgelFlHi/l8GJpMM6HSFUkf45OEl8
2TXLbHKLfKM9G0SID6LIrWwde27WD5yShfqvOfZHRT2Di2q/DMmH12WUBvKUdA1z
38EqF1MSchxFDkscWMbB1GrFO4GG8HMopu4qLDwVXiJCwIpg20sKuD6YLsUhAK/O
ClbEBun5pFetdyukhkstCwUhVIesAWlgFyhtJXR3haZ9vZouYxF3z6HKV4IGG16W
UfFqdhITYsQUYU+dUmMca6Sc4V1MS1B9gni84OCkfX4caJXdF2SPVcAZCK5Fsdzm
arl5dl5N70Ca4b1LkqP7Js+KR3YhYE5lV4sqWTFUsBfIxo7OMFjb1FhgmJk5I9Gk
o/YJQyP5t9Bt2KugM4gV0okdasvG/3EM8qZ7ObRVxKcqV+ZrRX08ZD3xPHm8H8pC
p6PWwKOPzZzMU1pY1+cDGY8ELVrLr46efwwc7RENQIT3PpYsVr8IUHedeniLb5fL
u4v5eAw9I8K5b2bwHu/0pQZZmS0NOqjccea4zluxyNaRKZUOGwPBanKfN7sznAzn
W8+bOGG3BlhqWS3I+7H8Y60KJockVE1JtN3d7gIlGMoTJ0PWc1BlJoHtNx3IWnqH
9ss0u/g/CDFnfkgO8+ciYYciZfyZwlFxt0WZTqHwOv91LMZqEC3B/PRwVoD1h/Hu
hbgP4zju6KZaqUFJCNIKdkPTlav57SvPDxsQ6Kd0+gT9r7nwSDgiANPcZdareUQG
w2c34836nU5N8nDLkBwrA1aaM/EYUv7NYtoqDXEtuxveAWQjO/nP0JxWBESHK+NG
48wLudN3ecrWKneAY6wPMyuCl/yIAvBqm+D9/6qUnE+F0DkjuOLnVEgAuncDnb2M
enqoiNg6dGxIckqUzJ08smVMG5pGTw17K3rd5WhUieG269m24Y4V5IImNVMFf4LE
cW9Y/upTDGQIzsj4cSJDJupyHDAwsRVBYXkCGxBt0OCvhyfiEf8gqhW37TEv5NJ7
`pragma protect end_protected
