// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
KmcGt9BtHDGjwWLsxoV/avdZzOgW3fwI96x+CB1lXhpk8xxh0qDodb3ea0FPCTOB
kbedaBmkXrQvI4RKNkgo44aKMwDYvl1MMfWs8HiaPOuzATosuX/3OfvLc2L87iPJ
6ldpRWWjW4NUoi+Tm0+qwaKb1Y7oqm2clTEVsY0ZIwI=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 3952 )
`pragma protect data_block
gKVT7yBRC+/kZQAnrw14jxm14rYOdwNU4h8uybSk7bhNtKpQmNl3gWFTpRDvXvj6
Om57zvTf8aQivX81eAUywgTzFI9q9XEx0Fjaf3zJEXOyNB+CWK59NRYGs69XwdCw
ocHOE2RXQYJpUu/5Jp7LpADum14S4s4qqQDZNnIqiyG9t/oeOOcfcYlHfYv72MNq
V+BFXAhAaWYWIcFRLhrRw6J++y8Cgg+JjQnSX7YQRkHOFvStlmNVAjQiW4L46JjP
CN+ykQTYInr9lnxtP6JtC7tmtGjqMF1X1ej9HWO0PYRgFdj1SC+eykXgL2HQ5Xkf
YADoY58aBvMmYuv1UWpxWLDeRVXIA418gs+Jv+ltOYpk4aXsDmd8/t7KHw17jtqf
mQhLcn/qSTDuKYfM0Fclc99kWuc5NC8MzZoBCGQ7n9rp2fbEZ5I2O34aMxsePQ+5
8I6RLb3qdNKd0Y6cC77pOlmoJ8kpSfzhYy1E3cTqLa6ZCHawRo3vy6ORGiGaDdSv
K7c5YXgT2zT3YRTAoDlJ58DrmY2FqyDbUH7uzS/AZE4q8j6VJRntQ4/ZNmlLeL3Q
w4ffJMSoNA0NHwu+BZv9IYvLKNzJDaugoOww8M2HtJ1hxrXfEKA3x6lONwSg8KKp
ru0ZGFfn+jMlksU46JNmomjgiVSHCb9oh8OJ8dq9IEwQcRdYc2W483TC4WrfCpXY
3/w8I9hBN1Q7W4kNBuj182RraLi8lwDk9kcJ98Y1tvNQZxC8fqyGDNLbH3AWQUgT
RPvNDPkp+BoxilOjljG2t1WSaZfusoriuXGFLJDlBkwRhTH9O36aDi3moYsRNUEf
109cikJHDOT34jgmND07E6MrYEbvWIZQFNwCgdFi7u9fbKmqMK0rcmlrPrasQbnK
xZaRuAu9K2J+3XXjdnNKD2l9VB+c3c84DVz38iLPxcCevrb8SKF/s87dvWVTHxu9
VDiS7mqd0idfDcuRLYZEfOcEneRgdod3gDvfs3CfRpjCEsNwofGFj4kT4S32TmKd
K/WeaknEhp+k+D4+KMezPv4tEIPAC+VB9wKs0o8uJxkeaoK01/2DsPXEawFeiDQf
4mfJhGGBVxWnDp5fv8Fa4EMCo8pGeSYdz688cEwm4VDLLtpStC1a3pjZiW7W5Y7a
ze4KmE+hv1ifRmFI9HxFT3ROufOd1RlGm1zWi5KcPcTDmadl4e42FMDth/jJNm5Y
oOJJ5jA0t/Z3uUTKg6yF3pM8v3cM0O+lf+DgF8tXEE5VxlpOGFe7tNpPhrMwNTfD
AVcSpG5cCYpRDRcDzyRd2Covh0gfMhr7IFUCcq3ys8dLGa8f93hGE12EPTSNVxsn
5FwgBnJ9tE8CHkhNVpHB6/QyNDzWrH8qghgFa1Vu7sQAsYmyxCtoH5o5qjJq9fhm
oVEbh/A7mfIBsPijo+7xLKVfqa33ZSr+OZqfsx6ZOsShUymmEyYhu8gvBXpPQOMB
VGCqIw33WXTdB7GyAIlb0beI8gtPNgDgB5JnKu4EvX5q2EPGLsWreUN7Mz7y37Lo
jrHpM5eEaUNLu474YD+AcJNqiCoDpBPnpgZUlr5P7RfsQJyMtqdVfYBOA0Mn1+wy
hg48PnXEC06OrmruvorzZr61tlnMDFGaWf6GRrV+qgdd7IHpNCGiT+ENsyZKGhZg
OfXcjhELke5ybvueuMLEYvTbyCjUWUqb6GlVIm4njZDXPC7ZHqr7Dm/rkc1mLh1O
wJAcKp2BgKg99usVA8k4C4IsASZ+MbEYvroA31QSpyJ9ad4VsUaxc5hLI49mBn/X
eGmjGbOc9wLk7vR02FaIBX04u5fYcZxldSNX0jkeXz0xYPS2fQI5yj2OnJfqDflL
Pho6lVhufgWvCnIiLeTdvD95Xy8bVpv+IIcjL+sbW+Qu3NfUR+1J5o8y5/T++dcJ
n0M7m0yBQmUEFdZbnCBUdLeUhsHfzLinYxtC7WPMRaP3YWRyRzMLmEd/cNMeDKED
X0mWngNJroQca0A7ql61KLElc/7uDjEYv4LZFSAJQ0Fm4eBa5ipqjFYIAt50igsW
aevlq4ipW1qhntJkUUBf3wTTmwExVLjDR7L+tpO7nKdONwQiE3ZfKAWnzl8PMZp6
c3gkmAY8f2icW9RpVl5CjgTAHkKPHdNdBiC1u58jHdb14uzoUaU7suFK4nxPIrNh
zTPskzRQC1pwOE3CwMOW34UbKCnS6SJzYgLc1cS5Lpc9OOYPBLt3Lt1o7zBVh53a
kMqCV6Hn4NdcZPWeZ4Ht5dvZ5Yl0eqV4SZIhPsO2c+2xK5E+w2HDT8hQ9qVAj4xc
7tSg0BkEeAnzK1+WeRfdnlUnc+ZhCOlP/uRITld5KNNHnZ2Y4diWLjmT8CMPPnXy
PYTwEzy6p28Fal13ghE8HFkPaWKtm7sC5eWZs96lJiitQuK1z7wc36WaOWTSaBph
zxLDjgFgagsts5ieQTPqtZVBijuCri8d1yCyMEMD754q+2ZbzfgcgZobog3c+rWl
Zz/x+zRVZ3EJFfIVInNMemTmB7j9owf3gIVD3WrQf0vV4JdyW0dJozpgUQowPaT+
/yVkk0SZQ/u689uXcHCXD4DyLew64K0g2Nsp8j8vJRhValmYwEyLKKyC3qZTkcwn
jZJsQwJDD+rDYbvQJmNReiJYezXlgcRCTSKV7PdALh8efL6P3qgIn/7JEKDvMayp
ca/QrLVr3nFU0cGxvQP4BtJFBwG14h+V1UCzC2KcKpEo23gf6xmtQcpMeOXv358G
DybPrq0Rrv7AfC41Fw+VdmkW1ZPFY1GPc3ami3WVWHUE3rQO/tGVHUAn9CDXwhZe
QWaENuwJ9omD2mO8v4rtcQUhfgrA2iqOMozQDz5I3LLSYFx4jNZQMq5BszjmAe8D
VSd+JhDIsO/CN21QjEZG4dm7hRsLDPWezf2WxKdq458kAqkqMSsrXZqdzYkWJvl9
KXrFKfulXpEuCfhvQLMqSm9uKEWVIv/9ftdfjsqEcq4pGGgx3EjkcyH9iXM3lC8F
n7WL5t2+9wM6eTyhKVedjqCQ8NGeDjq0biOFSQvlLSEyeuSI9DhU+kLJ9bwsKVNM
z52m2ONsWhz0DyZvTH2zU8E3g8oKFZjHnJGJwh+Ql0HMluBtauzke31VeeImPI2G
boxtIb8++EqxMRW5XvOW6ViSE+nYS6eJfppgsMANXyvNXdYuDBk14Gt4CFIouqke
wjOrQDaL8TcU1rwBlIy9g0H9r5kZwzAEu4KLp2UdpTa5r6dLp+qEGwQsOwQlL5/z
k4kPAR68qDbQqfgkM/2ehZN0wV2YwkppW1Gewh/i5OFJg4h5NrxByHwud9V5fcHm
faFYYcfIFdyvEdr3HDOYA0DJ9ONFgzIWrOE+kNpCHkqUZGGTvP3nlYg06CeuFXj3
vDCfs/C2jisODoSASuJkGppL2pVmsVgIDc85ePu3CdbzOe1TEU0PT5lO/xPJAYgp
WDnQFDJjVV8FyqNLHaM9+DZtYh6PEk4Qec2OUBEq2iYlmfS+GRrqv3qnZlq2M3lE
yaxDelK0oiv6DUpUVMUU1ncHdlGO+9RTD9fC0Ibq1yOy4fvkoUW4cLFvx2gcQGqX
DrvxjHMhQ7GxElq0CthoLsjYmKWbuXyRfxk9UP3yEysSIiYCBBUr553i5Z8w0ylF
bPsUjbmAenUlj8WtMBtK6iaRH3Od7pFvTw+Feicf9Idoug4HbaX9U4oiRdGGCGDg
DuNP8pn5/NaZ96wB0gYlBFQWnRaUl/mdTktrwKqwDzaxJPgQ1RCZAv1ZKpIVADAd
tJatU02rJhdPrQeY71W9N2DvZlhavma7eOaujw9SG6t6l/dbRSU4kJoJgmRTfeDE
RJkdZLL1JvV50E1yEOOTC1rRwIjnpwTWjTnHKgQkVsSOf/FXks7SkhhSLidaTB9f
0KXFxSXgrYCSKi4RdOWbCCxisH+ZkSVMXBOVbhUzTQlPGkmgOz9VVhnhkPjcVPoc
rTnK99fWYCERPp1RMoReL+JU6Id6NnHHBjxuRkA74ufVo1LzNH4FPMtSCk4L2ThC
Q6vVWUpB03mlOiRtKqkjW/ypd8azEaka1O+RloWI9pmUJfTme+uvDhEGITfwzHX1
fCevB+wmhBxk2Xoc0Be36rMlIqrCJu+tXa2JZrjX/qvFYWm0tnfVIWoGkzQ03HO6
4XzJjqrWqk9noJ5FU4gSchcsLcWv4vLVN72U8JvHWDmpTNGvx8VoulJoQXKL9Ztw
vdPrDfu3OFm1qMEU0MX0tlUYM9k0VC9fuHYoZPDMi69qh7nqCeupDulXJsiyr7z0
EBqNH1sWfuEnW0+aC8D9TdljY4et0NlA6uff2qYt4So2GuFbFj//PzocR8wX6Qqh
xCBtMTZ0uDmyJS/T/81d10MY59azU+4P2lhiFBaboPV89JEKc4OFGMFF6BMANeav
ujzg2+3mc/OrfjLkdysXGOtbBQ5tqjzmUuQ46J+BvJECsm4nP2kaA1TABn6B0Azp
XTUxqRCEwQMX8J7oDO1W2Jp1c1Q4gxLnk+IkxoIU+mImPySsJDFFt5D70QKpCNhx
1kAxEjRdPxXQzwBlw+p8acodbzu3DBrpIVF7mSpYzKhm8eJtjPQOOINVpYVbOxMW
sJwX+VJwzhLvdMMly7BZenrPSPJtP1fR3oiylQ9Id75/W4exmgt/PVQp+twOb6dV
5tbHLdPliqoboaYAIT10zqEV+4kCOPNlkfValvZcLFXM6nzJVDcSbKufXEOyGhHn
qIBbs28/SoIOu3JqLufNLbYkxbM41zIC+4vshBAFZPE00cYdzPNQmX3JEKmoAxrY
CIN4/4APVS8+2JziaLohlOd2xeNDnAmlM4T6MHNRHTIfIsIkHo59suAzp1jtvoCi
lGTnp22FjqyCAS2tW1CdnkcyxJBTYTyHe2osQpIHmb5pQzyB7i+AU02Sr4qROM/4
M7wPZGW2dbJfprbQyhbcTW+Ukw4b05wGDmWE3M4cjneJ7VovgQ5Vum5UcZSNPDhf
TJ0AhBJ62Mpd3Cg3ds4D6wj1ulU7HshjfPd82yMnt7HEmljXmb/H98FCJ+207qjB
58Fh2CuCtg8G/np20MMIgzTYFHgtZLv5PjSdcZIQV+RC22pf2o0Nuy+8ctG3iysC
KotzklZ4P7yn8lMxxcLoUPxnH8bBKmH0va8btW2DAD9JB69q94IUlT+83fvlG/qx
EzsMbE/fwPjyBWad36I6cLKqnykTUqPMeEo67ft78gyiTxLRoCJJYT/deNGaj6Ca
r9/JltbzGujY5nVZMzaNcQ==

`pragma protect end_protected
