// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
1w4c5xMdzZ49Q0njC9AZ8u7SAAaXL59PVJuBAgR03erNwGBvrIb7Q267b2cW
2/u0KTCipAP1TdJK+VVlVVYva1SdR7btwTRRii8OU8rpHhoQZwgjoDVzQhuY
ehUBqRsCuZ4GfypZD7xqbRcLI1aNaqXCN5PEjUVVKZWxfwcZl3BdTjg0vkn/
0tf6Csh+3i/2ZbKHROPUU5LmSBH/GSP/xdfPCUye3NA3bEAcbOjZwe0Zr0gu
5KXZCsdUpvPzvrwpGhigpLEA8VsX1DsPh6/tuawdrFg4lC/N0vOSX3kfZ1l8
SYmfkKIsS05bBXNRbbhsjg23FZxdbSEsDdqLRws70Q==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
AF+OOng48nlNJX5WgnYId/twDGAR5J9g+uSealpLWvChsUz4gbos3CxhIuJV
T+p24ymaGVuHIVUIvZv6OmwXhD8R7uMvPdKlIv+wsBPShuvaJrLoqxSDkYYl
hd1yMZmS6PRaRrIst1X7qk67EfDcP5LoU76KX/ERHW7QTOs9qSofFUbl2o6L
2PgueBmKsUNf+FT3emGj1xA+Kd4LXSzsupd82HDUfYpUjf0qJrrXEJCSaUxw
8AgkGj8L3aXexK31v4Zao4MJWueLTOt0HhnqYy+PZKpzmibjTdR6RLMotY4a
AawwQ8HKgBeosm6EkOfRJp1zgKUOAUvnIH3r+P2aYA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VxDWeOHNcWpK4VcLnn7HvAi4C8M6klDYy/o5QfiI7G/C5jWohr9UnZM/lY6Y
kQPVLGD+Q0MxJmSqRZJo+NSGao6GjrZPv0M+mxGkVFGjPSOeKzltD6FPlc3k
v1LR4b56Y1R3+b/C+tU+8cNjDIyqG2JWpQDvMtJzDvFAX0gpLbnpExm1rwqD
frSqz1T17K7TESzskW1nL8Kuchj296cim0Hd7L+7bg+6Ra8tRFLCBdTAUoFr
b66gBTjwd8cp5TbC/NLj87Iks1SBzt53eQKhiRT+3N0xT3dPHTMP05K0gDri
EG42cJflpj98Zk1bOyGGEzfgUNZTn1AMH5bWlYByYA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Y9tc2MBgVIY/5Dx11LFQLkmlDWG5nEKnRz7PrVvpDpCYusedw3hh4uHbz9Ek
EB88AVwG/Hkq2CpMR9s5M/DjWcO3DNLsCB4MxCbNSZqG4o7VDrfu3iHlZRJs
gYsmo2k8XTzdHU2bNcO88L7n6YVvILeq6kR1hplua/haPwoWTGo=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
pAP5jHXQozlZ02aUNKC3Eu4+/sHJ0qYCGBxeavLyv5uDgxJ4pKT0BcMhHZDf
4N15O1ML3XFrBWtcIRGDnUPaHJjo3RiCvOJ+EV3NWJ3i9s96Zc9zBEDrLNX6
NnZStHEDg0/vrHcNC8ftsNDGULn4xiUTyf9FGB+8CTJp8zBwDzzYQn0Uvab8
TQINmKWPltKgyCJydr4crczSjsVK8M0/ISovczvyF9VZ1zN6OagTpkhFPzkL
leLRB66FHGZM3DSr061bieWqrb1FFZlFEWhWYTh6HRM3GZBOhanPcd5wJ55L
z/JAbV7NDRgaB3ZWw6AWQpFQO/Am/TRx1NCGO3ZS21xDtgSaqSQIzUkl1MZG
nc+c9ZsJM6AsEFHb0rZ3oPvDhn5hl/ymt8iUAkdQp17DA8V/mWkVlsQLSNDX
yBLxYT+DiHFoZydvB6jtM4ecbKQ+gd8suWWyfogKc5t0iyu2nqepa3pBI37o
po+ZVZ+JkP0kaOTpElKyzRD1lKIOBK7d


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
N5fbrFZ2EDm4x4GRoXOj0/EPWF8ymLKG+8rxitC/Qw+G9TeJ+632vacSeRhK
JsJptc2X2x0OcESno+URJ1Vwnu4EzYYEsN1QxbuvtdSC1QO1wEygyB6uROBT
vNuKR5L4PzE4nBoljZn/ICkH+CReZBrJAwXBVwI5NMJQhKAs2Zk=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
DWjReWVJpoXuzTlj5J/sbCC42Xj3YU6Pir3bAX+jRau4JXNsy9R5MV+2Yj9z
eGj50kYBbD2CdWIeEH0fL9jD2X9RFl5MckurRzOEA+AWz4+oUhZLjOpgxv82
P9GyNHcL1ky2WTY7QQO81VdtNUiSlk4OtgyOjiJqVyqsOpdWxcY=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 5968)
`pragma protect data_block
viAElYF+W5MofPOTBMGQXfYHH95Gc7QNPDEutY0RKHgZEed+eN5EIBXGqPQg
7li/i7UgZMTRTa0o5G4CKA4Iuuh/iVwRHnYS6A4T0ItG043rjlNFmaHADiJO
Rl5ANSLP21YhcHJX0Xtxed1YHXk5rxKFRGGIOh97cd6gkxMPVLdrKZyHoCKm
WYC0gOr+9KNEqI+ZNSZV3TAyLXOb6seWWizkrS9aVIIt3mxePN1j7fCsc3bf
pSAzUxeHBOwTuh1izPILPBPGer0fknfys9sF+bPML38XEnUXu9KJCTeXnLb4
39sjzMVhquBhyUIxpKy/lShONJC1C0AD2N+5xQQHI7YtMrUiF5XRoA0yICnv
wlfDLnKZXP2SXsdtqsdp45+OqiiCBPgPmWcOQOHn7Y2zS4NiuFN6JvrsRQwK
ZjTDKlEOrx4tFye1ioSG7CfmizdVyPH05wFnaCrC2PJdTkOBaHNFJM8mTOp/
wQzkYy+SPtAAmDWVEjuDz8fN5Fqvrxxa4kcZbWJmIJtgmrAY3/C/RL3fgVKi
0/Qrk5vkmRYZVHzbp5IIL+XbKOC0M5LFT6vDzhrWCEI7I3Gs8txWtum6Vrot
R6P7D4ItBLhQz3S3x3RF4YG0rcb0i6qRHtUkTBQJAgbgVX4VxldGwMHK0Ugv
zKS05FCuzamedVFwZ4QIivr8+0WDQfzxoRtx0PNtut7WJRaqFc2zu//Cij0z
1S5E0Xv7fblwMWMqgCTJ+57ZeFLVxw5m4SCheTs/QTGddnC+xY1nu/LjxD5L
958jjZD3lvRQgmzHTnMGRxYlyhSELlQd1SyX1g218KlASJ4zKZnkNP5FX2Qi
yOCl9JhwMobgq/OwfjhoFC/I8Tf5Umu1IGdxytG67+wkAISdSYLhdrNeKD0U
CDm/qT+ogakqlLs7wawJpKaU9D9txdptj33BOOLCgQ6H49GB/9MqSroXxlvf
qonWdw7n68k5DUf3J8jFgVCTJrL40IneYw5N6IxTi19ITmfPJOmgoSkRd9Ci
7RAM8WSVvItQmR4ObUW4dWkEmoVKbWpGieqVscKIYPZg6RrOXn4lNOoVQnKq
MfTM5dVkSxFWzB4THr5I2NUR7lTgkLL0v0hiIreqkvV4eWxBsgA88vbb15gg
yz/nlQfLSpGkYhz3om8HhwL97ji9FG2hjvxmrjeGnlGDsYXISNCilBOWrAZ3
uWQtzjYgXe0vYkUq4JXgSP69rDnUYdWsiENb9I2GjXr1RNv08AfUengoIqd8
mkB0rKENEziGJrNZaBgIUKD9N9Y7gDspEAmhqOcrczT3R4qWAPtV9oGJcmhw
ivA9ihnFzeLqNCy7OYWhZEcgf0Dy9eoySW87ruDiVK0QwheCzPN4YCoMfKxI
QbBq7F1aJCy51jt4zmLqkRSCoZIhkXlvr8k2y9pA+aiCVldAWNhO8OneOSsN
b9fF8AXdEU+oI1Zw0hi0QG1lkdc6u4Sgy8O1Y8TB3LO6LtE+tmZtLgXYrleI
jApWUnxbYusG61U/XbyP6Akh2Ugwh6V/z0Fbxs/UxoVK/8/Rgn8PgsKMAIOj
qRj8J74U+MM1TwWrv/KQ2z6D2bCethKToWhNgBdsblKlBClai9l0SkHRFvVQ
sKcoe0A10wfnzUpEJu5BZZT0csG6LNGNv9hF0WIRQpkVIsNG7H/d5mXOq1yZ
N8ixR9f5Bol+0TZMLXnMCj8W0Fb71NDAT06W1K71PUbfOx79PG+N5BvNITz2
55a03UvdCJV7H8X54d974SJEUn4wU1UM/8kiGD1xVD77UsDfog/5Oac8GDXi
3x+AWhFTF3Zz23hB/3YZPSSaeq+6VBEOCC55Yl8i92GzFEerSTopp532xP87
t3kfM8RSqp9BNISA2VQiSZLydYPSy8ByaoJiO0+ppD/DjsHIJzFej1E0RDsg
eMNOmAxL6fGJ0b5EXF7SrA4ft1eojokWSBaSURJKhpTGAul5Wr70rB1JfSNI
YJDAwDwUr0oJ+KWvopeRdF4sV5GGhfowwThnvhOtPOVGlfeDOK0qxPoWHDQ8
uHGXbNFNTXdXu1vmin2IzlgdDV2nPOxGMnKRhLeKiPg6pmoqzEKcIf+Cm4pI
OxNqlkXrxmldXs4psJt8N6JqK7uY6p0wYzJ0xenzY72cIAraLcRWb6erkehk
cZKZY2ezwu3PPYXzpLOMXqI5+7PId0I/BGXBXgmYfZdtBxhsvFBrri+CJ4DU
PPdAMsDppHXoVeZKrpw/w1zWENyNHFo+V/i2lTP28edxly6rj+QlW3HiA7oJ
txr2wD//TnORyD6wwwgfHhfS/UpbJYCGI+8EhAMJ37n1KxvJJ/3c7hNHAjG/
AHZfxkL0w1FgRA6wGfLXbwIxMsj/bqtqBsiiiRPrzhT6LK2hUQJCduujXUpR
ZxHEVkXLcyIsLu9+uq/P9Ko+JNS7RPFdgWne2cxHOV+By1vZt8yHL+KGrXro
Df8/zZBcsh87VqFkZ2Anfhse6tv9nzye4HEeIr576Cuy72J/UZYANGrOo3tc
5r9be1DDGdSE9Ioij2fmh561UgiEsh6Sw7jLE60MwtZpZ9uuUetFc+kR64fQ
TJISWAWNPQm8XHY6GP/hxb1P0XBE9eLgozhJdQ6RC/WbmNX6MEN/GzBnIzh1
g+t64Z4IlohFFiuc+QYpd7h+2L+TenRaOJboWoZJQaLJtZaM9MykAQZQTuES
ZyN0qcAcVWz1gZU5bANxCUTee+ZnmfbCeEAC8MRlzXsCnqoiwE7tU3eZ2Ax9
nAJMjeUPrfziLVYlLodN4TYb2DzKL16VMan4l4aZZlTgSvHxmyL40UG22RaI
7U8CnZw4rjJf4Kx/RlxHXJqMq4ULBQHdOQiKmfiwEAcZ4GIw6X1mLL5Dtawo
KLbP1PsOeKO4JOagkllvD9j298kc5Uz0zMEW2/AWSjyKXGDLb6f/j4lkWnr4
NstzDaMIl/FfrtcDXiWg+TGX0bpZvwHNx2dNni5pHJhKYhqy8OZpJ44J2Ivn
9U1lGi+wh3eqaP/Qqv1DYPJ6yBSWsQIunUYpJVN1JsV0zsVMTMGUAazezod5
EDsfaOmK23nms22JkLfBKIosogIVvY1MoIIL/AtNH+Q9rd6Z+t4IJzxlP/XR
mH6ZWN3hqyAziFxKD/ZsGkWdTOYmapLGU6lzqVLm1iqjeQg1ELxv7xtlz+2U
2yt3iZ++OuEaEKZVNgojQ3GNeAnhe7iYELF5hMewkzTAXjBWWRBK4oAz8OAY
F1OfiPFItIXoQL/CQ9mscUyUY5e2fyJxVmWiA1m8U3RuajgeIS+hf7doi57y
0resqErjSZLxxmWa0ykwwdmhsvlRQGjLc1oclfOWUIW6a1YwVnSudKSuJpnq
2WMb+BV034cx+8wlBwQUyR3vzUrdh/hgFEB0a2tzNk01VkDDeh+MFQLivqUi
aRFGkedTbD4k8Y0qOY23jQEI2rjRrs2f0uYOcnM1VdN5TMY6cd/03fOCqMV7
vt+7aGs4/XtsWtrEgGcmIF7Spobqeac8YNdlsq5MIY9IW3w/mflSts+zEHtK
29RzuLsKoN9riKYHhhY0X8d2eZk6nPH0dC9NsPdIKmnAMj1PjPPJ5VYomfW5
LUOHkzaEcGODymZN3DxsHv2QWkSAQ44sKIqCfSIUjoujzIbAEUWxe3O4HBPG
PlbqnaV+I++aD2/Bo664jL/GrtBB+FqcpQ+NC0yadXx27/U/MlIrXhgxm6Jk
BxOZtgIElh/4wyUsNQZLEeqZJ3V2AVlPsmcWoKqY6k3vT45UoNS2M2w1u5re
VjdP7GfBlDk3+12sfYO8AvgJCYmLLCRi0Of0YBb+YBjzijHg01fCJ6KnbEGz
IjSTEA2Zcx9iAY8iW4Di3hNcrGD/KDazpmbshuPEWxLqv8Y7KIZrq8yStZu7
TC/c7Z8vLNOTTLCe356rjGFH4tlOcrjlIlqGYgATCd6vW0G358p0Vfi3A/xB
8xjCY5K50bxDiXdgWR2A6mswCy9jY1GbZnhcM4v94Bs0OAQUWJGeiB+ElCrf
N5Q3fXdX7vbDiaVJ+ABWhYT/8NhQA/rXdAuE6Y8ZlYwknAkXj+NFoTYKAaRn
5qf2PF9MUvFBIRpR9b5E6llAnIfQN+hSFsYfhb4XOncsmTfsZWIbZWdiLjqK
QeiTVc2xeYrH+Lb6wbSP4O60YPDli2GEJjMJ+XcHFOkyzJkpKww7BRtKB4Au
PR8Afpj8zQeIMGv2MDbO7cz3z3ExfYH2F6pcQ0MZfYv5gOC2kKUzHfW6VpTV
TFlNSiWSbvHaftRCHcuR+1sHRM8uSL269ujKsli5Wso+22xLcwrLq7lKEwn+
q2jcdr+/w6fcbAAIH9txE9CC3eQ7pYbz3SxD9epG41AOg6TPZVOaPurEOTDh
0TlQ+tnU+cRaU9JAEGExhfvPzd5GPu/RNjaEzngxrtqy/iBJIBDxWJ64vb5m
V3tsSlUX5EB/cm41VXGBggqGEO6LVkhk5Zt12Pt7OXFWOnoWm+YpG5WTWdmp
HC+Qa3JkKNrOAdQAjb6xjftcGwYOV4a4l1DTs89Ex7Glw4w76NkNTTUescly
Iu/XPiqCg5d75dn1RX5c2XupmwwSb8OSf9HmjPVBxQvEL/6QLz7lP+uHGzRd
P3DDMzRHzxVD6LUOj/7mc/AGFvk9ZaxJrhipD1boBDvT09N5nXg7VTbDQRp+
zeZaJPFN+FrScvDYqOAbXQC1vwhzqAs6CLLVjXamwfKrHNjkZSqQVBJdHzHA
pjNl0PHEU5WAn0g6MYFI2YKts6Lc13e95SvJFhE267/j4+nUE7rFKyayWgoL
TFiIDnOl28HAltqkJRNsWrCOIYrbt1FPx1ajJLBq9lZqLMYBl9+SSxVphMEA
XwYfW4y9Wm1fdlA2WsR2tRkMiNE8w1bqlfah1q4K1ig8julq98Ozo5qOj1h6
UUBr9Tz5kSm1dFdaiqEB8qXyPQM7fj3FOJw1PfivNC625Dj+5B4qLRfvCpqt
WpYaOaVaDQfkoy4ZsoK2dwdsX4ndTA8TEHCjtH+dduID1mhVGor87z+3WDh4
IDUJN0ZqOBFBOHstsL1ag7zNrgXgCvaAddaS60bBEbAG8Wth4tFdUm+L6GM0
MKxNs74mHlZMDrUY3j8df34pkR74lpMsQrsnCOGKqclfwpfhFvCbAyM3ytQH
MnUv9MdHWjDaKjxvdcCCkeDusrkM8HUqhmZjrZJwGpXdDi5rMHdkWAM1/UhF
vi/UrZkJJOrXKILAXIxi7y41mpAEl/XwEcxyI7vERr16CjopLr0NrGjLnpV/
I9UHx5+3DvB2mWg+6TiLzGU6fRMGLzLhty84oy0sx/qXIMf9wyxYOC5xdu27
+kcuYVqh5sxpMv7XAsCVf/KPQjQ3OdmKJzJFwDR86BR2F1EY8e4aFRIPVen/
B+EYR07AXHmnCNkCvYQJcOMIbOOkLomJ9KU7Vyt1by9Eb+5PvRq7HV2+4id/
+xtox7MIFWHHZrqH4uImBi6U0rax+Sdl2moDZcZb0e7YO01KNpvzWqn9lKDz
voVnGWdQi994k8pUy+aHiMZfqyq50YOhY3HGxmGLNTZajCUE+o3ama/48PuE
SHHFuWoOezlWMAvTSnH+7fJc73dYJSXTeHZIDqBR1DjDwYYB1noAIj/xC2cC
nXB2TOVFc582PlRV99lnx8SJCW5PS9CUgtlYM6t/jGv+6XB09KuPMp15ig7m
Dgz468GVoBmecy7OONJzD7+VCcjGG0nsXJ3tc/q6paxhGHiggwncYRhgQhQM
dwC7af6Wdl1k6gl7XJzceMG1Hk9+H0ohEyyMonfJ+picbwP9vSozGSXNVhdH
Yo9r1j9dKGs5N5r1xXMcis/8VSBGTwDbAFF1gwrcHshwbf3bKEqtAsYop0rM
6Gkqj1RetZSJWMKBGtbG3XVEeVbMnE0nXj1OhHcCzy4YiScNdT2b8WdW4ll1
p8y19Es924vfY+pVUxjvhtSv+Sw2D7pwvHuTkTlk8+d5hM9DafnVwDMlqK6D
OaUqMOrbYQ+HhcXHwDItagXgmILJllzQKRYA1tpzZ0x5uXJudu55xOjotQTx
Pu8GpdqN1hthwZZqkz0eHRkJBlxwqMO3fhwD13rDcWyLNVjv/OEbfkQgthk1
fiOKNoAnrBRr2SZGyEj5oNCZcnwPgrAR1GLQa9XPtOHEIxi04EMnChn85JT+
MDBCrjoOJNe59e9xU8P9arrvjo5L2t0ksBuKnbyNVgBI5lq6Y8wK5rmEa42c
SIISYh3H0TtoAwKmCDBfJbKn4x2yqyJ1tQBej2OVNHmzXoohyf9whV+h/7r6
KQFLevcEy8RE+rsBVZP/cEsPce/yUsuHBuNHsFEhaaM3Z6cMubOXDB71WgE8
CPq9K46tNURx8Ea5RDcqZM34xwGunSNJLMNRC8CHcXCgKTYyagB7Drth3YhU
z0BSbCGzAPg8EcL/tKdPxAYABJv9annWglBzNnhhgcAm84ILRdzVXT7MYXw+
d9CZ2Fou+gw6uTsVdHpvq7UEZaHLMYfV3fmny6z9G98/kCboG7+Lywy8BWNi
T9akO0EpB08LDkyvC3Qq5Vtxhsw+w3gnybyfyMkWghkHvSh3U3wcenLcI0XG
cCh3CK4yvZjNWZe4bW/WjN6ZPddE7sNbWqoBmNAo3Qdzf4lizKjSk1qBS/bS
qROVP6GwbvwsiA4pIVDvMm7IiuT/EbEKwZOLNfifoI2TTkEEGyNgbZM3+34z
gGCapG+LTutjtzqpZBXTBDLOfp0LrO1S3c8Ms+ltGCs38d4adunEG1erEPpL
avNRfMNw+BlT75iEo4Df3i4KLIofCYcQREzw2XSxTOjQwj+3BCRLbod9/h/u
ASV39rqzKp32mw1H7OKCbnF1ao5rDf2OThHL7gywe8Vf3JB1aZxielRxMX4j
0jmZtfZvn4ZgEEKJIQddBCczJ3PFbokRJbt2O975PL/ueUXzgyKQBSetSm2M
xj/zr3sf12+mZQIIa4quPs2thcmkBOn1LRuUdB7OY0jbAGRfhphcaUc06k8z
YZNvQE4S0JqQqpIcB5cjk7HGJA3N43cUiofe13xxtmTu9KnGrSRUJf2KoB8U
WWqncJu4mlAo9NCnxTg0FYNqxZg90M2getm82FL5l4h2Rhk3SoTfqXnbGZ5i
aKu33sGTevEEJrnDl1wkVk9Oe+cjUGHWXNVF4bjcA5MP2cPfF36UFRxefyuv
NABsblns7UyKm/6OjvPY4ov71crVacFiC+ECZs1R6ORMnUw0j7uDx/rtS6yy
veZ2DnZLOlo8aFblvgJVz1p9vcG8z/EBPijHlLKv9qEODQvLPa7a68IIJG2N
6ZjsgZNEiwTzDWfS3sVu2NjW43JKE9vMtJ3BkEvpNU5hcbLv/4H67xO7e12l
jBZmqaDgm5Sp+6FdZQWgA/lsi+G8sC2mOPRmtLEDu4uAQFw3OQlGFFIxz12s
d5d7tCD8jDNod45DdXlm05VPs2dgqsv2JByrdB9JxbiQczBiMarJK4Urpf/Q
uZZigMtQXfvz3ihGJkrAZ2XnOxG8Aoe84Musn1jO88bqXfHLVVsHzSKvhQsK
pbkaVF/4Yhs2/JgHbw8xVqIq5SgIMyVZwUuyw2IJw7dB9qviKkDwzXiI38TQ
ouOkNRw289LJ8VuNEAjIpB1xAaG+AsZ3eNwR+6dW0jE3iM+VPSUL5dFtT5B4
Ms2kOp5VwMhy/pkbtAsrxMV/3kyK4uk+Rc510STblfkJwSGKpT42zFuLC8mV
w5CrHDA9STEGBEKZyHX1O1AN+9pgCLD5QVNf7vR1PDgIKKRm9YShhAcQgBq3
z+NcxFEihxjX0EXXo4/UfJcY9mx3HpxYPzYEE+84nmUW4/wK2ZhueRmHehRq
WVC3OXdVJqhaUB2wZNrLDEfhCer/Aq3PUO/gC4pypL8wvVq/SljPc7dcPQ1b
eK68bG6Z1dsPLyFzRRVi758VfPv7DI+/AxWU2w==

`pragma protect end_protected
