// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kU4mk0oAOXB41Za9ftGm6HTJy1NcxzbbMWnCoNaMwWeEf8l9vhXPeomXOe2E
R6nDbWo1qNGB+nC562vnGeOYDXuXBlEvNkTnBNYUFSBCb615qvbO6y+odrvL
T8dZpRF79D2Ilz87G1mXJt1b721rmZStoOQHZYpwu9T13RdKBoYD2PKJRQJO
KL5C/rcV3iup6BDqhGsKAt5QCRX+Yzl4pEotPdJh2BMYoWaIDVYR1Tnp5BpJ
aONWoSztJyX18acz2dX2sBHuOfJ5YM9JnvVP9apJWkd2hnnJLvllQEbWp+Hk
Q/L5NDhRWMkpOmGQveSM3jPgt6WVL8SvJGSc0nXXSw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Fz7Iwo1OY2yqZNWJggftYY7rKget5PP11dq9QMFWJJfKCmRPlX/0MEd5hvVu
RHgeL09fgt4ZQFJ4zF1v2ZcFyO+sdQIjCaKrHBFuscGMyYIDNqcSrm/axB7/
pQAKuoIrBSQPTQ5bT+XmORZGVMYOSzuXVlHkYpMT7GRRzttoQF2U5tRJpxqd
Kru0SLjzdHw+pjMH1Std4ZNgr+22kbrfVppmFQLideX0beqIAsKzWpqOuHN8
94tGl5B3aM7UAqypcDkZhvkApXEhRT2kAXQjk8bWkbJtSC6HxN7d5tWhIiR1
cI9/mVuMz8nhn/c+wOlqRvcPrTv07ErNhY+e73Nivg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
aGa072KpmK33nJZZg3YB/8ROu6DHnbXiDMOvF76OqaXIE9I2NxlTddRgBljH
uFDpiJ+6wrtrTkmgn679EUeApSmVo1ptnpPx5cP+VzEnXWUKik0E37QbOLWa
CsxVxbDa4U5Bh9jjLG3L0rqwwhtOUhTimhTK45PP5JgjuJUCQwE7g9jHGMrK
PttEGsdMkThrAeKBQnODz3u06sKGX7pjhI2NrTTKxm/ICv2aTAsawMbo+U9H
pD5MmAeVZmqLmSTPRUEfBx1HYnHZxqlyEcFDgLQ0DgwfJsEiKIcTJBLLg3rl
PeBd78scHZOuSRKZ6uH3IYw9XrwlPVcGovnUQ3HccA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
J9imlfrBgzaBZmV7gBUfId7T+u9a4HuaY5cWikhjBwEB/8ffB016isG0hHab
MWLyYUwh0A4gpuA91ulyvyzTvqVY/XVBoMobqUnExFHeSFBRbO9T4Csh82vK
gB9OfNfj+te/dWYSiOpCi7sHQQhXHTB4xQ7IaC0Ay/087VQMYdk=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
k8ZtwyA9w2ffZamcU80CWIFEicj+tCWJ2NSt3HBDF68mouGh8dgG8266FcL4
m5/APDlA89+iWneCm4PczyfSm0gQEEYNA5S3YplLwIyv22pOEDUAnuMDMtgK
SvFBcHZjHUizDucH4iapzq3OxSr+TCfOHQmowQJLbAO0d0bU8Drp8y3pw/3s
FSTbvsJ4KyHYduJl2WWBU7dtZ4aJRlKMwk5SKBXvYdqLe4C7D/IgGSfWKIX8
tEUtHD5D5LKyHPz4fplajA6n0H4jel0Xh9AW8moF/yzr/sI8ou9LTAdDCbm9
5UyZZAaVmi90kVL09vnvUuYY7aEH23kP0QHGrcklHMbv9FHz83Q1vMtIpZu6
1NgbyYC8b4KNj2HZgarhZ/Tx1THCfTTz9szr2IFl2n4mYoetrWuX0s4sMdU5
qrfPq0m+Tj3CMBRlcY0zqa/8AnQe8kz8ZfyddBnoZzVIsp10+2NBKXYzGN+t
+zePHWxF11qTSZnMN8JUc86WrPMhTI2q


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Y8GpFhFhxN4dhj36g1uv8TAXT5MDbrbuThEcUMyT0ZK08lWmyFhnPhh9qgVa
5D4HJ+N56kytc+2e19hRm4gGzva+XAqVXTkcogG1MRl/Gcvqtad4paAw1xrQ
I6PyNoo2YZ/G1wPZx8ghdgKkhZYFPvJIzSjreX4jAOp+z8GXEnA=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
oHBlPNLNToI9P+XhlOPhoGOmCFys7hXx4SI2yWs7jcVc6zLXvd4Ac7KdSjxx
a9rfd/WlVRMoID4PJ6D/WzILEimpOkgZuEUomWP3BhBvY3OZ6+rz2DByd41y
Nl6b2TYTCKD3QjaolAYvSsEMaC/MBiHgy1csNSkORedX33fWtr4=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8784)
`pragma protect data_block
v630Mb6/8xFpl32UnTtu9HgBRRG9KEwCs87FuxyJgA5HXyPDy4xFzv8r2hsM
F4kYKI+4hsy6LnF8/AGkQnulpMh01JN1uX2+Sq+18rn2VNCqeOYq3qWGX1rz
mtPam/x5I99W88r9NNlFMbyTxKzMLpjB5Hw6uIolGOewTIPMPNVWybxSkxaa
jXsiLVdzghag9Som+bc6QK/d7lxsjQoXZzB8/GMPOK6SbK033Qvub/fe5DtQ
yR23WSpULOvyYc621JEWmwomMUb8OXxDSzYqLJcRzmvxTQOkADlWuz3IN7WQ
Z0z7pk2vhI1vp1DCK++i2jS4hDuK9qUe52esIY/7hMdo7MzArwl5jJcNtYRW
TfosxjBQUuhpgCbFOuAIhm+XHeYsfAuob9OIsSmfQH3QdB062zXAzVXrJkmU
8E7kFL35686OaXNOd/afwYq4Em5pZGrFVl08CgeKvW68jh9aDOTVKP+RDHtv
IQQy3G+gaT8rLVJ6KwZOzp88fjCNKxn3/KLwoSwKBRmnYI088OUz3HA92it+
9x2QU+J6/D407rs9XFW0spJz4HkUtUeTPWSH+scVl39V6+HaTwDgds+gvwkE
nzHTLNzPOToJjurhEsnb+9PFoGobaJqpXxMwLTDJ5JLexCjpdwWxua4ZJ04z
xJLSRZBcOMus8nZyIL5onneIlN49FImkfc9oszoUijLDu7nlkEnP/Y94PPq5
/L9hkBmzYmsmf/DX/gxkpkHrQsR62CkgcJCPNeOmuuvLBTOU5/VWkQXrsJgq
b6+jovgyejEi/uv9iLQaWyCmTIkahUJiTid+1gR/LtANPwzmvlyW4T2NkQoD
3gqEaPsXFrlU8ybJfV7f02IaUYgjX74r7LCAUZ3J9cDU9lOQsCk1+rqalLKq
mYcvDAZ6bVEHuOATjx3hWMO69wff07CoBk9lx/9TIJs5862B6Pj4KnEGC6aW
IoM+0CqJ3i/9idPqalgrbiB41YTj6wNXGSkJONGkIyO8QnX2ANfI7kPUIIVL
JgaH8QrwZ4Oy5a3+WV+HGtHXHkwiTV6LTfEHJE2KF63TnWlcQaoEME2Po9Bj
5SIJwjAEwLsJFHhsptCl+DYW7ItOXGW9ivcTMYUjj0niYzCxeEiZElrmUnPk
qmKQtgURrerxZmi8OnOzYIkC4aMgwDyBIYxjiiCucQhNYxjH+YcmprdcitjP
RU6qoldrDO3uljiOxgk42MmCCQpJSxjbXWYNxeZCEUwtj6dFvoqpJ/OfGQ3E
bVhIN/f8Y6wCCdfRcdlDskcnS8fYfLx3F5kXQwAh/fitaVrKtmhZ36RxT+Gp
9vS3DvmcfvQi7Uu37aK0IyDOLMLDfAnP/eZHwZ0mIeXhzF6/rnjaJeYiIuI6
PPbSENqCr187OsNHn1pAbRtQZNRNOgNUfFj3ktFGmpcKDGzX7bxNuvjm9M9o
1VwI/2sCKt7rjP9iY1mCpBdAtDyHv0WQLBToEoXyOO8y8idGC1W2ObdInCWe
9XRzAA0BKdt5IBurxAXensSt8fAWbgeMi+XjzU1mBL79nCxydBvLx4MBDBuh
ZzbZVip9iX8+/Z01q5gm+KAwo3airkH6QiEn459HUQZCUJ8QP/SVwmowmHb7
cCYQ66nkY2orfhcldAIp2n1CymKAVkEVfQgk0FwBZEwq8Y88tAPzfajyAl8b
brNBUkH0P/ntvXg9DxZT5+6fqVmZsjv9e27t/+NP+KHUcNiCWpeWGA/Zk46H
05wcWWgNFbtvgmy8s62rqr3+AQgxD7nakOqCpU+8McRJ4+t/A9ZqaojyWiYp
GaCMHCFAfjUOoQGHQhUqvFs23IBpRUuHrMJkalk9XCYNM8QBdlEwumEwtnjW
FAs9CwjtmU6Do/xS6AVtfqunPxC5MWUg4srcMtir8ECqa+LH6zCEC2ZdLaXn
m6KjtVQWStIW0MBPnvqf0v3g/Ty/p4vFLSdskxz8Mli75AAmlMZvxxK/j6bT
pC77vyO2Ab688SVx1krgO9okNvN+rrB4D9nfIC9m+PeAt1U83T0o4xy1gwLw
x5/PsEHo3nk6BSMNmsiHKcJesoPgq3LLTjM6NO8I1WNyc21169HuikbMNk0B
wHoX8neBSXimNFfSIw9ZthonTJh4WdCYcmhVlBeF6to/dnUVPeSx5ypYbToc
IWKxr/+9m4VHcdl4bQs4JCSJTrduItjL5AwGZtxCG0hmLBXvcviygtGpFqrm
EKXqRN7YXWPm0BFrcdmam8/TgBbDV9pjYiSKKTtNL/x3XHWfNGDsenTvoKNq
n/rd+hgsM4dKjfEY3WXhQaS+9H48dAwa9C2EYqex765MOxirsI/6Wd42ixfK
rpXqXLn4G5xKKEJ2oQL6CiQvUkKJCLs5pdcSICbK4gttNa+T0Vf2AEAhxnb7
N37TCQDQadwDdkvvrv3Xrij/hyySkLKjLN9jxxGVWktGjAr9nmSiFkv0EiIV
G5CD7CNcihqVUlZhCksYt2VQ12TA81RRqdMz24P6JSSTYPpjtf1hoW6FHpAy
G61kGUf2qV8GdEWid5/YClLzUEA99uUIpxTKVVRo3mrEbrqHRALQdn/oh/c+
zU8aKraeYz9AFPz48mxTXWHaeAxSr7jfttzoJxKLZ8QV5pytgfX6V64B9gsL
JhCdIBV7vsblMakdjgcKu/t3Q5xD0LCqyDtvl4gSPO77/R8WONXymCTZYGND
RBc1LAmCkkvRHfIPF1BuXmpGfTLRfqqYJWRYL+4Tqs8tKHwkUq9HQKRnrK27
2ifwO3Y9gPZ7Pc4QVABxrDhbSLnSt7w1MSlUH4Z679s5ZKF+mZFn4elD1oBN
9oe9TJ52n6XDAbo6Lb4TZhxVX4/qpxhmq8GzEdOB9HY7GXJe9lydeXbrLHFY
1Gpzr8SxvJRxulwl0/ZkEpfjVblUexdeD/XFoe3L2rZbovoYMuVvSDtAoZPb
QAl/puia3AKXgk4mO1EgVhnFhQvgN0km+qzSUyKxIEUknUyDHBG9MQ/ZMB6W
zYTS+qNW//5xbOI9ED6WFZNIpg27yQr5clb5iOGkUbK24an+MozY9ljC+DLD
w0ccLrUWm0QAkZgtlwIDQ6gJ2h5LDYv0CoOwKNR6zBjAWDfEekdG4MYhFRR+
FEfUA+xTZRJlBgz0HDdnyl+h1SNl5J6+TxH0XYKf2eZimdMOZYoelzeKmBnM
6h2sYvo3WcNOJuORN2jI5CWhWHxGhbfT5xtsLwWX3NELZdFefmJ2wI7heTBd
fKsnCMmCP+IJa3sPUeLa1P3VO/qQCr2iyo6JF0uNFsnp3uvaq5meUZODVOQJ
TOdIHJ3Km3EQtixOD7kJmL1oN50vJpX7DtFFucDrOm8yYFu842QnOpDUC2wO
D7hpwfPbJS7j03/kcGDMeIsGt30/dE7ct9D0aK47zKapJcGODXKlTNqvLtxc
hTfdo6LdHRl0qobZHzL8V7z9H6tx8YZl62WzbYiK0VfpuVtmeTkTSltxLNb7
d7AzIxYu3sS1PfUiORUgrHbwt824FwysfZkfEKCzOJ/oR4PIx0iNeQrmycnz
/BTVZmSZcHmWugc788jqNQBl2XLIjSCLjnZQj7UwCR/vBS9qBP+HQxA5D0Dy
yc3aWq7CogSzMCADL6cl7Pqaf0lbfC7dPyzVkQu+RaGuPKV4oYtHl+IM+Etd
wnqYc0NFaAV8Oz3ZSu2EB+Pgv/wOfalUhTiuYOR5IwLjYXMXImjhmO20hAib
gkK2jFfCwJia55jTZS9fu+2T1nQe4okAKltm18XEEGlKS4qIj07t/9iAhHuI
rP4fJJXML//XuzZsKRmKE/zy8J34XDBeFNn9PKrqpluvOqK3YV+pmrRHgopV
A7z/++bK+QRa1Sk1nrXHrFwPyu3DdVyG0a57AnG22/ufHtkS/toVcJJO85AZ
plod8rrq7QzTQyU6k8Q6fUaHkmGf/gX2zJ0+/jaKmXg40unDhqBseUwKiN3r
0Ml1fmFOGomK8FyhbA5rhaNQ3O3YqJGS4+Bc7lhbzY0gIV6M36XmJ7cWH6pE
hlhKCTgZ/yiDJmFHx3nasvTKFrAnnmfA8e0YFRGLl55oPu4sEHKEWwYaVFdh
1WblzzoHY2/IsxMLLBGi4aG2Bk0gEztrx3tRyI9SnA4v941+VqijlLvOvaGw
oKlX/7uSZ9iRx+He7B2AckcfQ0+VOInjJBPSbtm9gLbXSgIzLsSEdaHnSY3K
697S/2/GBrkrD/tgN0ea/NEyyIlJaF+bMOzD/McQIW46z7ytJPzbugnedF/1
wNjItjZWwtd0Tw7pgUky8SBBxYVLZ/qW5tVAiNQprLdmGZC5HYcYzhgZuBRx
arPPXKZGfQ8W2R9so53E1/rJLl3TfgBoqMFZCjo5+pNnXJukr8V8l3WyIBV6
RAoQL3hhdYzscgQJnoyzWLbuCaT879HCQ8i7FRZ0f1jGh2R9Cfb78mmD/3Xq
k3J5ZwQBEXMmgyIxB2m1nEevbM0eqjIW5ALDrE2vQTKRStCUBTlB/v0okzzB
xz3dKuNQLQcavBkd4v5ZT6myXttTTb/BgLHFmxh8GwJS0J/kD+ZSv6IxxcVR
QJAFX1wvsNfIl5BoErnqRHS+tR8xx/iQXPL0+FRELDPel9NCqcipmKXJIyzA
5pE2TKLN1OpXJtgMRMjMKvweqI5oBVlIANwaGyuFhLvWgvN1tn7XKJtFkBJD
ImvPLDgRU/boCYm3kueTbeeNa8MAZhhTP+aAxLZfelxYClzHTQXpDPDBqddz
cH1MjP/kSijFT1TjeUDu6E3PwrSG95iczQsW83e1p3Fpm2woWaFNgYi5W8ZU
zdydw1RotCzUmsC7iKGUi6OYtww6DrdsyFbzTHr7WoRJ91IeuZVISZiDx0bA
iAIhmhqPDclTrjd6ahbjaGGjWSN8KiFu9kpguM3kk8xSo9i0oLz4srnybAX0
QSJxGA5rGNSYNjr7vN7w9NkOm86ewDgHhDXQgNjUNFVFlN0awI5ZQf8vyzde
cba8HqfyToCOClaGw0arAZL8LWAtTePS3OFgbWbAFP7r5fcBvLtdgnErFM8N
shm1Wnzs+wSPJOmqkU/cKP90uwcbmmgm5xom7i0wK19JREQuZvKLvEE7B6mm
tesQnxSVHKs3i3uti/GCcJ80CHaiLwvB0UF4knXdD7CInr2z9wG2SaKkO2aI
OsA54vV/kJof3Nt1fx4z1Jc4oemkqqa7Oss4o4RbJhIqlsKgsyjcN6dWnp1D
xYJhx5b+zJSXzdNbEX6Pp0veLEm1NMLNxOkwWZ9wGan3O/z8ixmEaeUSWgl7
If6WI0Pt1fJXfbzINqGGTK1MlQgATxj+uAZUHBFKVmzM4m6Yf9h+A0D6Tmho
VPinYPGu/xrHSlVVaDCPFwp7zM2u8hpPQA1NLncskyn9v5ZA28dfy0Nbr81v
OIHEL/PMY2zFjL6CFlHH4HQYXrMVmUaWUYJCl6+OhRtjDXB8WstLKDcwkBte
3SWfhe2M6VNLxkrpBdukARFKiHw1A6f4/8dVB3/yfzbDdwwOnf5h5l0Yadtz
c7RvWWsm/S4U7la0iW+O4R3WZ0EdZoVPv1whvuBwsJC7dRFrBve2vdDp/wJF
t7bDcIkej/RdZwvt2GBWH6uFGwX6Z/UcC1yoeL3uGZxf0bIdE+8aW1ouFQZz
DSi7kW8t6ySAjrOXgikAs/stT+D2ee6jgQKWSIhsbeKu97JDxG44dkCAt7lN
p+aGZC/wdGghZ1EecRlg0zy/L/FyiiU2nKkI9li+256eK0Q9EpQfFguRgnhC
sTvYIMD3+jcYWQW7E1uo0DseOYO5it8R2DXF8cTbSzbiwr9hR0pky9ZKak2M
IR90LfSBu7laYScCvUqnEe9BoxAfK+sCu39kuC6Zjq+PRmcCKbKYeroDCMla
4xLAgCxDv3qXySGqdPhaHYuOcGy1cP614/hkdu/px9bFEBWppNDtF53mczKy
Bimya1YAVF+jTUYm+m+68PUHiWNlJ0T0+mS4j3HXsGhGeoQKRKaN6H8u3E/G
kbRHPfey4SkKVBqMXY7aqlvTcYC4GeiThjnSeYXK9rgnqoLQfmpFvM52RF71
fuMb9wxOrBlyoeShGvXRwZ0G/DNqgTj/yGjHiVQOxqYCQQE7Kquq8QXJs0Oq
wVD0lGJ+cHk18ooclurbbpTR8vhJYlo91D349zpnZU7RkxEeBYqjC1nqbXRM
+9+F8LzQnxiQGjKvz6MhvCbIZ5RmSwxAOfbODs1IFoy0j20+9BmA0pyXev+i
8LrwKS2PmlzsEveWI4eaqeFd7r84fqhUcuuWAigwgeR2BYxPh63cr48P87TK
nZXCrtuJ9zPxiVchX6IEF4cBnb4Q37j9E+PJEC+uYuteUqejjoOU23LkyUhs
F4Agxib1vUrFcQHDyHs06/fDbI4Q0YFnHg1dkZ1TpY6dUKfH+wiQ6Dt/zWkx
a/8paUNNWpNnoEbKiI2UE90oyrF4mIt9sUU8i60r/Dibp/OCVJddO/fR+kTa
Ix8AAtl3cYICK++q7k/fyhktI35myKxqTGn0r8ttS1ZdUwqcwvAD3LHcxwkG
/gZ58NHQ54ervsKEskUsZVUqkrE+KE6OmWuvo5WkhbgFa5CRFHVA6SORNNYt
VxnyQwTcasAs/BFXddsOMc2GJEU7CZ4gkyZkaKlYays8dXfiOgvkBwpilOUa
onYUpxOWL6OAOh+5Q04uE2Vjb849R36Vj5JWlzb8wc/LfesWM+Yq6YpJc9+Y
xdEWg/0qa10wkwjcXK37cTTGl+m0Zbb8cagQLjwexI/SH1zu6GWa84zDs5yy
GWkxsmCpOHpMummYYukkCP+2ijSz46MwRDAh29F92qPQyQRdRFrQKoZf4BSB
2PLje25R8F151Yb+QWuvwnsUTfD0Ib3KUwj5spuITGD4jqGAzCbe6uuV3iXS
mtYGejkAAINZf6kVzKD59xTlezLv0OIY/K4yB2m2A/GLZ5UAp5Yk9LpfpwS3
WSok+xCTga6zVQITiSCnsuiuBrOsG3YcTIOtiJtMu96dYVM+LLe567F1RrS2
s8lNMEoJ2euv7WXlCrO0x8fOkeLzMfnubJsn9nvYpzb05MvIBwvaaAsSN1eT
/YcSlhQkuRNn05FdN3zmhz+0FdAIzrLTgYUXdV+GF+xlZATqNn3tdsFRHe5Q
RLHTjU0LAZJp0tJh0mZVk7p2kViGbxpPvcYuQtyWPb2HbBZyKROVYDM70n5o
474XLzbyUaB/sDNiFFDoJmkBHSr1P8twxJ0eQSfY+NCaHGxn+vpoX4U85mYx
OmPTkLZUjuPF85G+yuE/8UdKApvL69dkauMgqnnSvg5kfYgI97j6lvhSnf6x
RI5ln2XZoGhqA/QvFU2LiIIkumILLe4W0IJXH8G41ABAFLsYkIs3Et/gHDuG
/SuDvI5abG+15+oJTkCvfr5iWd47H9o+kaGg8k9l5tR+ZCz6bUWNssz07kdf
00LZrrnmg/5v55QYImLs/FRgH+r77ojs8JfFF6R2stfIjbit9FTXuYQBgWJx
hzPJNl09SsdHYCr+hzTY8BzOTHS422FOWzX2ge80LfxcMyKP4I7YmsaT916U
IrJzT29w+TqLzM3Xc43tEu7GrY2K1UrF6v7SZ3+q+aTnikYI2E30+M9ib46L
ZJ7xybJTXNPVMiF3PtQU7bdGGq4Hf9v5sV4Fknc5naL+U0hN7VMYMYinyalN
BpGQfMsTlVrOi+VR+XXKXWd50B6llm1y8VXkT3alhnoVtucRZcatgICraXsK
h0QLaHPp/KQOhxDXtz+8Yq2Oiqq0pSDuQubWlYC0nUQJewFbcCT95VxLnxax
Z1YVIvZVX6Y4F5v3PPKXkBqIg4UEBBMay30UJFw5KkLdULRLk8GzI3bYAf5K
X7sjgLC1HWnfwe0s02MGPYHXLFSCQF+TK9CFrg0UMMwcMdBNB2TCVfPaA5v/
Q/D2hU9Glzen1UP+QwW9j/07JGrJAaXEuaNoePmkB/ds69wlSqtZ4pK5ZkJT
jAeb7E/W7gzrzVB6YjJg3q4Ff2dBdIUS2ChX5G0n4j90ql1Ps1fmP4rTx4D/
qDLSbqwU//+Hce0YJHkSlhk26QkrJEEzJzTzcUMRuF5MTYWdY12LlGYaKemx
anuxLAZhBtzE6OrMXwwUbwe8CG0/fIcqHbOwfdvFTGCfxqn+5nYgeA3ytj3l
xtCkic6M2/m2eNvdM8ic2YDznIDc7hxtic9CLX/2jJ5szuNjcmYgsoLel5DZ
T33M9VnXZV32yzbN/ZhaqoXdQZZmCiiVjGU31lwGgE8Ce0fewdBFlKNwVeYk
+VJ/iyghva9rLMaqeHUEQc0zdua0qlZ6ImxWvDRbIdrUTSYHC1puYyKnKqAs
nkf/JIcqtINa2joiJ0PkAY3tIPQwgaIjzMbIJ1kcL6zcTLm9frG3MKLI14Md
/CfUub4NhIgqtcCH0ow/UbTxyHD0qH5Dge94J4wFIeuujTxl3FMSKZBg7Nqv
6T5Q3sW7Akd670wfocoKKXfjhgfGGsYS4g1g9pcRC/1mzqW1ggEB25LU9KKd
3kxmnJxTeEbUu3Mj+n8Z8eeMzOgvGVxI3qbmokY8snY49N27sEA533YYx5iK
zS/rFqm37xZBTHKvCMA1qfRTO2k0ZB0z68YN/idAwH7S9pF+Y5ziKzomKCZL
/sGoDfaLLUe7ZneN+sWN99c3sBSWmGMNH+nCddGRbAEVgJcY54lB0uFXEosu
vjs2OEeXpOtSssV5yPd6U/GycZ1rNDqZ8FSpkZZ7EaTNLHKJuy1G5BgmzH6f
9KUo0MXNEl2sNvf+8pbHzvGHujIwPtFPj+H1WCNGQjL5FpXqSukhKOkcJ4yD
SF1PN8KElNIvovZp7DFffiyeFiPquICifMCTCdgBa55UxsbPzRLYMIvaX1ID
n1x2k6hV/o0L8bBDrTFbK31ng8AuSx2qNqwGaz8VVMG4H+UVVYfNlBAfR135
xi+jvtA6dJLBwoKy8w9i8tefNX8w03x9QAIvxskEBbYjsRS09p0eWQM4pH4a
b7SFURSZuOMSYbj6QODydGGLd4OuPVPGda0WuIs6X637qTLtG/QRxSMMyR9s
IeeL9h7/fS01cw6kQEfxKC6TzcUvnmI0FmKBmQKjZve++EQXSaG7kmT4B1Ss
/3rn2EW9LG7+d75UlIgOdeHXD1VJ93Npuo50mefECX+mffyAutcJ5o6n6zeq
g5fZxta1YghG82bi6f54P1pFwUcIns6SuboI0CY4GdyvJsvgff9TJG2M33f1
oRlrsg95zWyYle3/xqlU/wT43m/dfNXEA6wkdXyfGVdX9sR7IxI/tvbpsDLi
dTFpZdUC83q/RNMiTjzyD9xS0po0c4r3jirNnYC401bqbt0CpPQbe01iQ14m
WUaDTnECER4SENqKPFBIiuqq4NUIsJCmWKVVKYF1DOBJBA/Lacbx9rWTKBE0
L5pqd6rJ/lYRMkwiKJgEmIeOrXzn52nqYzT17T1jdvDefLDkS17lBSULUNGN
jvwCW87wvpfPHaJnwDXinpiTV3yMTBVb2EIoQ9bBcRjAXQu7w2iKbaH61iWl
Q3gZ+wTx/dISk5cdE4mux+G2C/cpC+UGA/CZ8CshBq1vckuTjI6ivzYyWe4D
bBCpCNe7udUpu04C1xi4WXrr2FSR2wN0K6ssoFJX3jn9nA+Qr69d6tg2XOnJ
kUGK+26No568/UzmIS1HFqfFZAsSwSOo6CVAHTZGA45nji75XxrxuwQrLAav
+VzHO29YseQQEdx2rzoQlOnOybAOWXMAFquvHJaDU8nALVxZkZbb+se8eTW5
wnpdRTMx/KyAg+2sWpehIOAMd7lKg6z3O53S5CHHT+k62ykvRdefnrUkCOlv
wa50NqYlYMtL+w7VMmeHCduvlHKI9WCTdIH6SJx4EKubnAtEFz7I9ocZKXYa
ofBjJdNaxt29I/MJUqe4q/EFo3T4YtOCe7sdybcxW5aq9fd7YrbL2WB+h3/8
wwy4mKTnXHTOejYi+ONk470y139cF/SRDNLQGJyg/uCn7M435UgjpAf7MJZ2
p1RNYvX5Z95cxtYXvY/1uJhgmhKykXSt1qREAzshzqKJMc6m2FLVB2WrJCtF
ittpPllOs7ZpoQoTe62lUmsgYgWEn+vFIgsFKIO6QcbzzbQUfUumhUgc8xix
yFlgz+88NLS9rtDPdRNvfWP4poYGL1AIXzQC5JnXu6Fu1CSq2d/LyhQ6gJXl
lkYsn4+XQ7dicb6wwOwR2/xx6KH1qPT2rHmMajEFrLwTKlzLSbotfUhPgOVa
I5niv5/ZNJYl5IDRllsB2+QC21KfDOQUcAGA1zCkzHR5QVcNkV+hjbNrd8lg
+i7tlQX7vp9TcRAVClE5/mpAJTmJ2y/C1wAOCC7oNR7cFAxjbGidcUe8soot
D6fBZpi5zJBhKvl0pX/CqBSX5PCx2FrdDwrp3ObNOzMlr57iEkkUpi/krDGQ
tp1Uwfa+P5m4VtH7nd/R5gMuOh6rq7Oo6Xs81Kzl6vY5DLvY3Y160fMv66bo
tOJFAxHcYrf9n/MmlENaVeorWQHvmbA7mS6Zru5jt+aJSKY7wgSHjkCrHWml
xm2MexXo/bWZDR4Kro8+0frlPTfvFoVLSnlilYZnzLcGzCZZde2QQdrfpRNT
tg74goNlQtJa46Z+CSa6lUcrpm46i2YGrQJX1WiODbKBrH4/tw888VF4NN+7
vw9IR79QWi8RP6gEIzlomG1Vz+3+L+ZnQB/IKRjpaWzLE3VWOP4ZpvBKZJuc
gkvDGNaU6IzMAX2Yvc2ipVTLLx+mI0Yvp3c96I6Mvs9/fnlIFpTB+EUeU2Rj
Pj29y+f7mwQ57nMwQYF7CaY0GGS+94VuFaQollk6dLYzkDdqS2hWBNx7LOX8
gVtGHG3Ur4VXngk5KP5qrzrXQQBHSk/J2bk3/d41G80OrpesBliS4wbb6EAS
qL0kQWZUV2+lsGwyfTMCOWSl8D/kVoXN1iGPtL7trVvin4jMOgmma5EL7mc7
U1SF/4FkiLSLuY0IGtGgAtZoWTR9gPnWOBQaYKMGj7lyJH4cRUznC6O5mv7M
i6k7pDsEWU/SnHDhGb5KgO7hSiZA/ujr2LRzkaQFpHyw7h6YuiZls+8gBNFS
2ujQOLYd3mnTHoUWmrUz9FQL1h97qlyi6DsfuFR6hrhVj8B2YqpnR4R9dMLX
jVvFUY6BuC3A1+2fZRCEOtg6IpF0p8VnQCGU7p/ihW3U7EUV2TvLNL09pNCi
bwi+CR7yf/fccuWEe3hdnOBdjpDZZRh0KgXJMp4AAe4WHqx8R1xLvCQ8nBZn
Sw32bh9oE6YUkcz+Y+6HantrR9/g7TrBlUbuUL04IxODnQ9PfakL3tVFchKz
Ue+BjHTlrgBVbNYHdtQGDJenZv2wOVPx8Yf5py/3jvJEQ9vCllPkphG/vVRi
GWV9XlPDu3KgvoD4Kc/qrcn5FKlcORJIQOgUQylPzICgs7qdsUjbmkhjSiDb
7J+W4xPKZsa5Qq8PGrYgBzppLwUV6IIGKue/9UAdo0ZKOIOPeOaOUVpRJV21
Uv0CHL9TH7RYTFufWOrSAqaLawLJitAnTIdp0Q/JytnVzxfgLgLCmhrXsgJ4
QaKuDdXbXElfsiJ2J7fyyKcnafx0YIu3sNYM0b/NSdFyW9Ab75qKau6+rMBB
ltvY63HIr0yJRXLKwOBGmYdKmopofK0e7OW32Hoj3owcaWduBsiprMwWAQDi
Z19WGeMysulI

`pragma protect end_protected
