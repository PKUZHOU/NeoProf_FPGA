// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
eG+nyXCYaH0dqjUY59MVjjIPFx5uk+Fj29UmMqIJJ9PU0o+RYiIXtu/8DLPzxwN3
pO+9XFEwED2Y6lsxKdxaoV7UyxX5Q4Z7z0Lw3IZbIjicH47oS//WQ1DCNprb2Pdk
05AnS4PGz2YtadoFPaY4egWNXJqsRk1yFcm2FxJY1j8=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 13008 )
`pragma protect data_block
YbFBODCda5ROrRuOkFPAqDqk+MofQ0et8r3+6ubciQnzd5PdfK7EArRi15L2Q7uj
ZYa/9OxKdG8XW9QrdqiRdpDEaTykPk1HQIoGw/djFLZ/fMEoNYa4Pnz7PiG1BUIE
PhMcgUs6h8lWKFLUXJx+zgesSHgbn2PUbrd8lCI0bR0WWRtZLKO6h3FNtBjFBUMQ
tMECuggbazODgqk+enAHPUjnZAl4Gs5p+Cm0NRl4WdzhimioKC6zmOLTQqmDI+Ho
VJrUhBosYLyLQWgnshlKWOsv3tB38fmFgdm4oevPr74kd46k5NSmmQdhGLDwI5tM
I3jawmYwP/k60TY7I5g0VhfeLiin+oMAQ2YuOWgYSi5Vw9N2nWteXioxYkRaXm5W
S239IBmYeWZql3Ht3WzWf1R2fAncu3Xp6Qcj+jqoFdGW8Q37sycVTZKI+AgSYVJI
KnQHo0Ayd8zw7TAuUTINtHvyBbtF4FHU/hklIdPbxtOhhJIG7b21njyu6elETCeC
c/7f2UhgAcnDlRmeBf3L0o2bKjUnuu+nzTGQHQNU5B1aIFzZt0kwa7daUoUdOVS/
vjeGm+YF5lfMCERcb4dXxcj5VxF7HQ04tLaxCLWTyVtruSiLl5cGNwRUtVKkDFK1
wgX7cDCwXdUwQAyN783k3Iz+k0lZbgOMgNn5HudqYmD5Kfh0xK/KOCCXL18eKdGL
Qgd9w5cS3WYIFOaPSx1hEkYh3xDFD0lSqU4kBgF5AFOcJJ40z3pnvyLitgint5Uu
gpq3hXpoxn9NgRy8G8n86xFHOOITQgWadR/hdYqdvIv19O8kMDptXUC4zKyJsUnQ
G9wT+81JHm9BM+b8nfqeHjZryuUEONU1GBwAbQwSfx9NO++stMDXzMVZde7fcmhq
6h8vP5mB5UGExy8PtJN8LUO5Br0CWF8v4ZB8dXhx5gclu9xKgx+Na+iHCvhF2+8Q
bYrJBYfU9by0gNZhbn4oq5uRX0mvs7HfPhK5dEEq6Qg6dGsSfkfXuxbV58opbq65
4aWk8gpb5da3zjAagnjWIFpgW6NnNkT1zYuHNlvMwWeIr7O/Ax/fdvbDzmrZ/vhG
Lr96y9vfOPh5NMWNPD3EbLp19giG/9PgBeWxjosS3CYl9yMtEwBw2Rfi4dCLppwL
FQA7AJoRUwEbwRlJB9k84f8fQGVoN/tU24+RCOX+PfIWNF67U2IMtclfCZv+UEKX
oUIeeyVsm86UkMPmdoTNHOWNSrdx1QTPGHJ0JHugQMbxtcM+Nv7e2R8eMHdjkD9a
Ij8p5FVyBLm9rGcTBzLWL6+yZsOKRKFNLDUsoi/AvANTriSq38tSowJ8XK2FUccx
JnBi44cIAzs4BjxRfCCHUCCHXeFPpuoCDo9668ymKjUAz5JUGg6Z0BBpr4NiXBxu
7RtOoCWTS5owntS0Qhb3PM8ebyZysncHRAYXQnYRER50ReTzI/UN2E1R+xhxMysC
nLSovQq11Yj0M/gvdA7vD9wJWHXfy51bJ8f8q8qdkvzib6qYSEh1EoFupNroOQgv
XItLNro8R0NkqJim+YQ0M0PAsyw3xYJH6jNPAFOGIlfZi2nH7hh8HX8j0YLW1iVC
DQ8uT+955e3sCca6mzEexj/yA6mcoJWDL5XtlHD3eKKEvepYNGDSXzCpPsYdRDse
XV5v7Ochg1F0Aq+buy2kBaERBh3g18vuYOGsyCTrzmx3KHRd5qDuwdn7lgGkGeby
yVDqHZswjR35KwbzJLKl27GxgHB7ZFblNjE2bUgIbQquoc0TYi3JxYNJSPAst27n
Qu8ccUfOSw/w1s7TZialzkwTSebtbIt0q5O8WLMH7Pjr3p01nKor9+alUf4h4Zw6
xk+ABEyzDq+iPVNo+Q2DSjsWA3z+FHAyOLCpWy/kRvX6zN3H6fUvnF4cMcEFYeAy
c4HQQztHZ8b0hkqbZTRi7yBuIR/60g1bKLUdZdDQrTZuZMwCuE9efACM9PfAuC5r
BNmVbQpW/X+Hw5UBJqb2DLDHYncQ/J1VDizhvSE6rKPbooaJ2jKyJHiIuqYhzniB
ZRziwWDBXglc2zlGHf+xSZvZNbV4yvvOMWA4045GLB+YRokSH9p6+4iMejcYHTyV
b0mX9pqkiY0FmoVBk/K1oPiKfkDrzeJtv5aW6Cjx9E45h7KuQmQZ2cJhkMlaSOyj
CoeyRIaIsqStQPEX5SE8d2nQQ0P9YBJSIi6cQ8iIjI/dYMzyr1Vu+2R+l+lynDA2
3g5gBaKDB4iRkxypVOkM1ILaZUqo5p50DIDA5Er3ZZ9BQPZXYo4jgRJ4ESTwu7PD
FGt6sdDu5xFBl92xoILkq+tu0OTtU4mGJfcMAhNEj9rAIR40IYXYaKbCZbvz0vh1
3/hXKX/OwDnI6sBmhlVkdoBnMvCRKxd9T1EstoQAj6nJPHK4ak/8wSKs9lbZWMLF
IDhAcabnoT+buLhbIhb1BKCu1E87kPUXxnSxVLOn6Jx3CE2/p68xVq8V5I0RFo3K
4ONYUxtM1JVioJHaHtCvmoOCIJUwgVUlQ48nd/fKByJnh4IQxIoCZ/yyAHY2DFjR
t2gD9tGOQzgzLvZK5hv+VUyQmzTkpDlF4Mtk1kIITBhDGPAaHs3K2NEkeiATone0
IKCYum/XhufJ7RJJDyiGMNbYqD5kqfVTV+zOu4tnuT/RoCckoIW3CHqmyI7IgmLF
l3s88+uXV2vWDt/b9L5T7o6KMN0gcOday5xpiKG8bQludC1tdOT5/Yrcyrhj/SxP
Ei3S7xEDh+X7dRY8ptdIQpoek9wO4xBpRDq4XwCrat/+JYppwjunm9N3ilFqBZjW
vpOjd/7yac6TtKXJaCFdSb4eS+YAlqkMsbl/d7Fe5y2MjJOauMLecQiSzeRswVlk
W/Hchw1YK/+VaeBmqdVDtAd2ZplCaHObnWzD1oVEEc7gx3L5thNoIrs2lpYl5V45
M+MdL6h1tkD2KPslIYlLjOJafttmnfoUgPGvQZcp7/vmYmcOIE/CZ9lX0/KM58x2
IFXw8B31VLjEUatGz46NlH/555cf0E91keh0ZwaKj5bTcc4JovcIMyidXSJ0tQab
2dSbzAW5g5gg4Xhy3O4V/IoL51YYvBJdIftdkxEn6TTaeNWXlnAnvZbEat9iayTD
AxmDgwX/8xg/IrPXct425tlW3wRxOqyuIdUs8o+4iWvUW3PR4J54x5coheH7agxl
d/h4IZ9gtPPesaTd3XYMow41T24l+mT+u7DcCrJlFHa5vzrc+nez1W0DpRh75wwj
ztGb51nTk1qP9lExK31c94X92wybA8YKBlOQDBndPcLEiKr4oEQialm9Cc3fagS3
OCPWw1Yvf4YGleIUpfjQPv+h1pSb1bU0GEkyaAg8lrU/1bP/3jRog1g5WExQK650
i4vpTKV9syb2wnf9gfepnBmb9eQJ3bluuKzDSIhRi5FYgCyJ8AVdGyCxuXdN7DMS
UbQo0H03lz2uq9Ad9dqfPofmrw8OQ3vEKMsHs5+Va1YeXRMTcSDGxui8dZakVsUo
nVW/eJHHHwOo3gihwf15ZMUlEUjTvqkzx97lFXp2b9E3+YzoIikcjTGUmyDpt7LG
b8wM7ZwSk/WTHvbM9nB386+fj0czfRUVoqXF54IUJKIHHkyOd7fpkQtEfL2ImeB4
UtIr9sQFbY0FBDbOhxXFVnfi/crpRR5MieVPLd6GuV82nZkr8/CHbUNNM7Gj3a78
jcp7rsVcvicuvU9hf5adBBt1nu/wXWvhyv4h5n9G4Y8BT6pwY3sWKXErlyFnSx5v
tuRQW+LU0r4cAPxJY2gx0a78WAWTI1i7Aomt9FBFCnSy/ywk9SYX8p4PzsR6Yr8t
62t0RIFytBjCZVQdcvoDfrdxyH39rHs6ayI3F6wjadUTCnPRJURKVWdBHZeTgB4R
S0LSJpyFOHF/f9hrByGxXmviC1l4ZjiLNpnfvlArgWc8wJAGWQf7R5WxnYoGKaJy
KqTNrv3tqupcqUKu+BOPpO/BfUUqanP6otkIlj3Efju2i+J0k+APro0kQ7qc5UEL
QOBVKw4cAfZDLGN791pFESjJJ8C2PS5rWIJEXEvrwfq72OdgT9jWjZMxPEUZnbSN
N8syxjJNevleGwSNi9saQSpREVqMVjs0RnuOi+I6nsBaOCmtqFrEStarkKyt/ktC
diowc9YUTp+KuK3tR+q0JdG9ewgECTeazQVZ93a1ZkKfob2maY2KWQDB2h5iEM2+
DTQXfDH2TClcujESiaohIR66HJjoPP7w1nWz32+91e90huufzBHliCVTZ24aOpw9
nMT3P7xN5Uv23kOPeYXSokQbLinya6WukTbZYL33NjLibwU0FBh1PUBEm1sLiU+I
/W0WqarVI13nFreMABlnRfy3RKRtDlAVFPKaiXoHwJKuaDYZeeQrAhV7S3zzAizs
Ly6q43V6EQ3IIFisqYDR9SPTflkcJFjcn7VTU1zqKgc06iU1UfebWS0E2fPVjPWc
JUrZopBkqsUoGVLtQgrTNdqRJrXFTvRnFn033kKpE38yADfb8+8MT3kjJe2xGTmZ
KwxlD6JEb3a97yu9ptOSA4QMNKeWRanhQWwjwUGHTNXxWm7S0ad4k3SfUSzWtEGo
x/5iBJWt1F9SwtQ5V8taxlanPcD35no91MN4IfZbT22YgMC0kNEkJ0xa9nxrgYiU
cLbMleFiqHAZRpTUk1gmFAgEEZJYJY59WymZULgLrDyid+JjffYhB+gpbdLqqVt6
eFbPSAtqN2v8fkPA9Mnfa6Q/Y8wfKQgbnTO9BaEulvI1ZDsKNb1YU5gnGC4mvdze
+7EH8qsskw5JapnGCwJo32KNII6Dyeo03qqoIv/eDFpEFwtBpmMzwigvqqeRk+Xk
T1EBZMEM95d8RxZRr/xxZyCFWQhCDyvO0EQSW6+HZIwo9Mvu3HDTa+QTxjjTfySf
DuygZZmcJmvjiwZnsVOeNXA+n2y3ygVV9rMT5ihUcifv/U/GSVY8gCTP4wXPT6g0
uCsfvHc1f54eYqQyX+drMuunmHLRZoPt/IzNFiKCBRYIglC30GK9cmGFwvpGpqaV
CQ29jpDFg+vnjWDUQlmQTQxwgTdEAaz8sXyw+PpStXpHViWMT8aBvYNNzBmdGXIF
hFpoIk4nKLf+xH3exEBJKd8/sRqR6bQBTQsIZsihQoYXRef59UmgRMzVznYVXQ/9
1d41UI/JmAlF3wMpNYgg/DZlnjjCSowea0UHRJNhPov6afSIYCaQrkvXzazc6rIZ
w9fENZv/bT75Xq5FOOMES1qwbxrTqWEPQPxBeCRgi5YPTz+QDfrRD/tZ/HB46mFj
aZaetxr580QhfoaOOi5jL77wl9nwvLIf7tQinvz8webXjW+r6wxv4XTu+jqPDbTj
rm30sXfnH0HapUOkWvhhgac25JippAiGOahopHI+6rptqW6UT6fT4ujjFpYlGWP2
2aO6eDSoBKi6vIRhyjpLS0pVg74O4UyYWti4cq1uaU1StnF7wsAXgnB/FzqVALZt
gaSGAGPwda0ZxSSIjcnYDX88GVFXZzJhW7dmCrLRT8iIkaie19v97CFhlv0SrXTi
gUhmZkHgfaTQ3Tfgje8gfoJ6IbJJobMDKsIEwJiyp+//JXRkffEhVA3d6V2Me+e1
elzX+MB74h7t9disArbVdpEh1US8AldUeIjfL+ncrFk3V6xpMfcKldhzJLJ/4Mrs
bPHBxpjaIyl3S4+G9Hzss6R5C6SRW1Sdy5Y9m+ziBGCbbfDVRcicHITLKyUHeTKS
b0UnNBXYNK0RcNQBubrd7WSD8Te8VZFoJ22tLTxl+UDo9MNHScsbD8JzDlOhC+EH
iO5q9JoX7o7O83TMVC3qhpHpfUou23vfGxAgaJjuuYMDti76PFn3m+g4vFRZ/2pE
90TIL7CRP+t1sSYAgZKzb4jz8SMoUUTHfR7Y5xcrFPxtyHC+F9eedZywY3UQ89ZG
bIIoGj4dMWBc079sfnummxGjmIZO0HqygAmcoFSRM00OwdE0zzyPAnAO6m8fuB3g
XHR3/jq4dlV+4lMfR2X8dgYFd2HKdREaBR11njTIytnPjFWJonXDgQdSr7Ow4c+o
P/DcsVy9Gw83OB+n8s2YbQSHNZdnJFQPsxCfxFYjX0JXf3upD4hVqKwdYnrTDjrE
z5tW9BkWdXA1//Foi7FgNszGCo4QkkIhasQFnv2hqutx2omOCQnBWEMB6CcFS/h1
vkQjriY+MzhfCOIGN3RZ2sPeAwVxMJrYVlIyDCjClWf5AFm8GQCGCWklmQ0AP9Iw
jyD4u729d9wCO9rKyrJr4F84nhsEAlvtmxit5OX/R3pyDN67KEE2pSxP8icv1nfh
qwSM9r4Sev5tae/xYbfMfL8m0rvoIrgELYjrsFFxspyfqtSuuYM7S/2o03VHyOj8
xSUTd69TEziV1yOPXJjMKYsHykQqS73TRqqtdtDUvo3PMTPZF7oEQfego5Ubwu/U
RccjIhQLDcq5VO0HdrKYC2NSUtw1upbCLfRgj1PdP3PobQ1vYLIUoxG6zfV+d/gg
mF2gu3yLDeG06PCdeWsBYewghBQjIQRY8l+wlkesvxK0NRZHvknxM1A0cDb94cpd
xFOOU24uxVQ70DWLmdGSdGRgq77kxJiIImiMgZg+sFOtYcd9Xamhg9FFqgUIyPQR
io27Rysfha+QPUkjhn1Yc0R3EtmqHxhh1VX+wWuL0CXon2IbLH+hh4gHZtAW6QRi
I1e+91yj0cCReEp0s3IyPiwpSv8JrchNZhiGDKr1kBRWjEQbAvGHaB2b+IKpS7HJ
SNUZwDcLQWqnmirP1/FJgP6FBIw2KUJMMPeIb4XW+i3aWms9qvBARHA6BhcUin4d
bvbRTWhECZVtES/CzAegMfMoCpacr9ViiOWV0kyAgDoJcV2jdo804dO/y+EZ1d9l
pT3PBieO+iaeT4X5ToUE3Oxy60fUAgYpeQYj9SbrIWPSO/yy35EehQ19bXBC6YpP
e1zcH+Dx80rWhsv0FsikuE8CM3Yf7532SONqrZC1P3wmpR8+c9yBMkFa92XFqJH7
/PPQrzH1TaVr8136KFZnTdInvhZ1qV8PXxFG3zPKpAYivv9a/CoEDmpcLjaZ8zG8
0eS8fD96t98VmUmuTtCcJ3iptdHwJSCGltekTKBHv2QJffxtaJYVRtXhC1FtouYf
HOoFVnt7L0BmSXsjHTIThULhVqnCzryRH+nOZxTbpaBVUNgtZt3j5V7oDdCBl8wB
o0ahRT7QWSUgWAp+O1uS9Ll09+lB2zm/g/HPyy2ESM8/x2cGp1ibV/X9phg6B3Rv
lhXOqXQr5pc3szD3k/fOPYvWcQJ01UyKGBdLDMMIEHDPhhiiRosebtfqljWH9tQE
AkQVX2lhksQoYio5cReCqhLOc5NmBh01G0GrM505DVoGqCndjItF4wB/FDo94K+q
6u9GM9lmp7PpeaFmn7CbVkcyw9tlwN0VWaJ3SxD6CFRhAzxYVeFNG9I/NtH4npNs
vlISDCjZBpBAbLGr4nVLMF32XiGCnMzWmB7UpJ6c/XkgVfGcsNlVXzR46S9Nr+oV
RIvLKMWmdo2CanW4+oIRgMBuOkAWyWtYmSzEVHXO/9UuC4b1X56xFG4UbLDuWYdR
8+U3sAEjcZdkyMqdsJ9Mat/NhSGAMF4kRLm9s607ntOmgGLu0KFPByYPaGd2aqFo
RXs/UCXaiKbWyVD1+C5nIdgOYlrD3SnxpUjIiyxBvVyGPYs7rccgc8boGKHq4zoH
C3ipQpV8bilPZz3FGjP+a6tEQMdkt7IriOCH9dPwfGGGtgEa6jm2urWg9OkIIkRq
x9H+gz3FwPHORjzkv70s5+HIMaEuamyPd3dHyLUjULelLjbpnDoZve1oAZeZ0tqX
ou2aKZZSvpyucgZWbrK7+cxQa38D0rOZWE7D8TdFKP32Mt+07qjroSr3yMi2fZSA
j4bBEgsBlCvCusyrfdCSKNk9XeUjYZLehfp+t+feRiCLZ6VaPIUVnHbiOt5/e7XC
NY1DiVYsJ4wzB4Dm3jGMMl3Cr9r/oZFLOdAmFu0hWKoFXMHo7Ll+9ffvcyo2hT6U
MZLAwW2HVz/8rwa3m5KEmamEoumFpedLIHTOUaKJ4dlxZUINU8b5JP2QtvPYilVg
Ix47C2p3kC9dSs5y6yskUs+b9pfaxvm/DIrffP+hc4Z3tjDZuEVscWZ0C2eA6m6S
Tiy7vEKQlhZuVO0d16zoxEYx/EdnhtobZ2FhkEURe/Suqph4C1WsFM6wEQO/Zs7p
/zhhSihi4Jk7W3p/dk7Wh0tlfRv+kq85FUIMKMtE4TYo29ono87gUx859PJ84vvx
5opv4ctra7C4jAdG4FI/e8nsUtKlxFwDOuzXGYxMVZmmfqnVDk4nZpDev3SAvfGl
VWy16fvAB8gUKZzzrPWhJydVlUhIAf7DTbJuYlKByleJ/oBi9rnLUx9a2b7QwuFV
DAIx41tFZRgJ1v06L/T6e+q4IPndjYESH68MtwjyC2IbHBecnZpQf3hX6zbqzpIa
78WrydyEKCn3d/1leSm5tO2a1BbC+CgDjNpbBVgy+3ESHOgwwNoX49pPAn76pFwl
DAPzEsAzw/pPMHXKimLsfs/glS7SbCyWRCI41U/mJXIj9LiQr9kZ22jUL5iCoYNI
x+tPRXH/F33k7fAnXVouBJkwsVog6mWwCXrCsdHOaoyVcdL5iEsfheXrupaelcln
Caniyur37XRoney+VrL+uBXpj+yFc7U/MfALCBIKKV2i79xHDhnwhl2dPze6eCUJ
mBSHj+kkEIIhLt2wMppgluzV5hHWbT6C6cVda6oKr3s1hLPSIwHXpUNB7/aH07y1
DDdOwTH57zYekxe3KuVe9gWqpUYRauu+qbIp3kPVJhV8usewkqyp6JL3NPkeuBM7
Gh1Lx4EvuH4IZgkDuHKVy0O4/aSLbz4nfnFBLS6emWXraitNXT4a9rc4mX7hShF5
thIni6EqK63Lp93sMDPHL5t8xBdsCRwLBdMFAdhFr9SAysEmrp10j3BFq9ljk0Y2
35K2ZIu8NEYVDIKg1ulm/SXlfNE3dsX/Mrayxw7XO3aYgwSiedOn9qyRz3fz2nQ2
74L+RQNzAhwK+m5kyi7gOoPw4VLQ/put+MuOb5Dcq/IW9ba4/jgx6q0M5IRln73g
JBY78G3xYtQqM7wnf1MeZO5DU+WBaRKnN0mVQ58V0jSBjjwYjsIjFTNCoVyjLKn3
l7ligNLv0rBztLlTWvyxGvNCB3xhHSA7BAtMjBm5BHxQLpJ9/3Kc9b79e5Fa0S+h
4CdVu3gDr6+t8Nhi9hLCWayal/PwlJ6a24U9kTiiRuKS8FtNSzwNvh3QIgwH+r4E
MA2xIMIkx/zCA0CsKRgBjZ8r/4XuJ+EizfSmc7fNl2hVhk3SWndtPqkTGsrgGb4n
l+dPtDnfcHRws+oGYQAzn9F6TDe0b2JAFX07JZujeSAzhDQODrrUTh6vIywq3t+e
P3oc5yOjL1Gn9fbXHEuSCHEuJUw7Arhs7qAKOpP6KsgtoAsNiJBlQkojgsLOEBrh
8GfWXKE61K8C8HVyuYSJMsPF74LH7So+YShviAYo5HnX65bN89S42yLceLgK7TDy
8OcZGANU6MfnqXdG6pGwTHFQFtU4VKc2eHlLok4Xy+OBvMGqSxXUK1mETgYsEVas
NVOJneBKPF3E6KRv4+aEcQuPsNBjJ1LawFEevmG6MwwPzTXN8d4lqwOCimRsfE/u
NX7LHxpKUXu0EOvUzfT5YFsqRbZxH6SqEAb+XrFgWyOzwnWEhUSdASrhFV7vfQIO
VVdG+T2XVlk/NNPaHonq9JnXDRebaU3c2DnIvpJlIgAqwvDHBbKYR7eVNv3KrZlI
Dhx5buvdKw/FRsMnS2S8mxAV7oZkBsgzRceZkLRoPV9zrDt9/PCbCKoQJdYY0P5j
ylaEjR/ckA+lBrjflev5c31aotIl1Z2387w/DBUye9mhi54rI2sTUSAhBNquSKsS
rcO3JI3ZVNShGcD2PpdsYvze7PBZPW4iBREk5oDJt6ZW6/CUwIhSvVD4LwYR+gmG
75wnRNDxj4FwbuF70ktKLXceXIh2QARQATBGsxxRpjc6tID6XTsrdaEF4OV9v4ao
WmPtRqTW/MK+4MGKy3jCRROa2iFnSoOBQqRn2IBmaqITxTK17NCn0tgEvNkM2ZoW
S1fkN4lTkRhf+NI8rnm/U0NSt3YFiTrwITMluAVHr6DPomdWVxHmflD4cB+ZatsP
TuvH3Nn0ElnfvJzXUIHau7o3dx5PgIvvUjHwJ8GSRSxMrdb0qjLXGfyGPtkW2NxW
NjFgV4a2P9HO+f/AWrrgGnUxJjq2wQG+z2qcELqxbpK1L/0hSXhvKpw4UFyoSJAK
dSXVXLmYnugIzsdlzL4hFW/3o9fwCz1gsCWKOKKZnhonBxcQ4NXi3SxWknOQMijZ
FPXTdyonTep9MYQpvt+voMcL5iRdmGUrwYRq6ECUhibfTXYkjmyieKR/xQaUfbbd
C4RwFzjTDsv7r5CdpTuPMdkU9MFydqr8ycFMC4rkC+pD+pQauO2LMqdrLiCvX7Su
6Nde7mMhai936FFBxxpQpcNi44aCUAZjaKsWtct5ReteD1N7Xo85Ml9As8WJ/RxO
KfF2KnYwCCDWUgopujXlaFjdes5SlGVNY/rjAIhq5TUVGCGDtkmsGBy2rABdXrFQ
C8OjuPcIEO62Z9TYv3LZ+TgTAssjPnP5/5VUpAhiYL/5mqz/6S/we1v0Ew5yXvaD
S94EhqcBV4v3VWOqJpy12QUMse2qesTJA3VVIaQcMYNg2tcoMbsln1qFRVcSvbmf
wKs3xRj0XvmLohNu+10tEwWXh6bywKoEE6R8MSHv/OxlPSZF4fKfMBPNtAakNv7t
zaMBySjz75Gu4osa8UNa5IQlp38O9a2FXiUez1duTq8vQEQymg15VCkj82ZU6MOn
i18rgLcM6nvU7JaQcXNJC7KkhebR+6MEsXuHYl0sJVNTZ00miaNVpqpaQaJ0CYiv
QhzE0mqQO62ERRlhxzT9ANiDBdTNe+glW7rB4j7JWwiDJQf9GFFO9P3GNfeIRgue
9lujRubQKDi61USqvPdo5k8Y/6mUKA+OR7zs19tWepZ4YGC8d2Pimzj6i+qz9J+Q
p9Y+ZsPd4abeO9Q3dbpuPuVnlAry1bGMFHnpRPeDp+nnTu/5cxm7sQ+owirqqoLi
7Vqg7rI1MxdUZCycrEInm1GK8nqN8XYqSjneRrAIz0QMW9hV+f2Uidc2ynVpSoWS
eIRaP2TiBQoY0kt+cs02BTq7CPI8YziJd5GJ04wWKJCbWhbGVkdTFyWRXwbotHpp
NO40A6ITWqIjKlmAXwPtt5ee/FW1P9+6wCXzSTzQh46eiLxgRlj7kFWvSdkix3U2
gwsggjswRCtJeoxm3dOOGKcLZrOIGooni/w0UKJ0H2ZSFoGH3ez4Vl6h5E7gTlMx
tUDJNA83kyiQNPqvVfiJobqLcWQL9mtbVhZ5JJtyv63dC5UTB+tmNLyQDd7j1bm+
ctsVlp0jl6qBU3AaJex1wyAsbl1/N+VjZQAsvn430JAgdp3wFJI3otK342qH9ulz
RdSuHG8YH+JFExt3h4yaUAFwz7QsSYVhwdnnnPCA5kZ+E8hki5zsBZVXTi84Dapk
WOzuhSAiaFv2SW0ijBl49bNW0oPvr/bQExA7g/jXhRpuLrfZA2rZPWoxTEOt+NyU
1xXRmiq7DrUxVqcSZwzG3cIXkpib4mfDNR4T2vGluF5cOozLJ0z4HgKzgAG37li5
ThhzkHu+8m5SVYqqS6pDUEZxm5Y3+s/OR986jXsgdUhPdru+9xk+vBozhwUYqvJv
tmMo3f6uNUS7W3zgP7bhaPFJSShtjWkhA9dpkwu/AORtqugLF7S2KbmLhjZh+CdA
Wl6fus5Yaz3UWZgM5FNqNHiVAj4WRYzq12Sku2wj+Tb81DVO1S8l4H3gM4AJtkCp
Mli7nTrwfCmjkxMcXJvpyOeaX0UREGmZ2Zxb8rS51jyLC2SIxWz+tXTzqxuLXgBX
dE9fs24GpcMtci6RDB+zdmDUqb2+vaEvCSnT3fqWSThJ2Q4MW0W1pv3aYCpht6Bn
1cZw7n4xH831C5Wsx/SkSR4QfExZqzivxMaUhWbrs5E5CNk0xcucJ0GmxfNr+n3B
saEU4kEXGq6TwE9BFi2SwnXkg5GtWpy94CtmJez/o5ArlfpzqqArpqKXD/aqkd+d
8lDRrYlsmAVB9dmSepf9sFZZsopdWjWyIG23nllfwhKWyq1Fh1R356Jdejdd1Phd
zobXysEz9rXry4QSFVZtz6RWWak1ptUBZq/95NVmWE7tVfojyqNSrQVdYfM/5IoB
FmalizPpjewGPLVH79DV9Y9MnH+Xl1XAtjkSL/B2es2R1yZ/zStedA1Iu74MHCWu
miSqoThlN4/hTDtAr5NM5VQSWJtcXe5kG7LCX955tp+RA2o5JO6a7KVOF8O4z5sc
Y1E67+C6PNQSpVJi3DOIEMynfi0+UJlrqX7R2h/QkVyWkbKmYI5hnk0t7sVbGTmL
MHKSey6rflQpGdONAIimHxW0fI+pgtydkLCht8PGpFGOeH9zFWOQADjLWpcIsJqV
U33QY6YHP+WO5uL/mw9ScWbLFYvR+wvmD0b1R+rRzfPGSi57R8c8hsx2vkFJohxR
TPw9rcPpWQuTqe04dCtecvCyT8Z3LHvFR90ALVntQJMBKeZVzQfbdVWKtFDXWZIa
i+VqzSUss70ppXT9JorvHCLL7VzIeOBTy0gdfHfwM/Zr5zhDNAHSiYMsLt2KXDZl
aGhrba9aAHecpn8rKkTao+f+wke34azF8Fs1BFEvzor6pCfQjyQCD89MlfEIy2ih
wMhTSVBBfJJHXRvhiQH7fH/1neDCf+pcqdeq1j4kC2rccrb17GYQkhfxTup0D2pO
cnRq1uIEKB8/pWbJVbtfliVPce91Qyi83tdhiGLRtrlYJXwrML2uf6y013r9K4ic
okrx7WFh0po1zIJ/BpiiSeqyFK26m/4uWGLJMEubE8wigzvDW1jUa9BrtASiKlfJ
gPXVF3t06rSla84dSXgzty72TbDrEQ9O6MSgUwF+61eyExkJivXsvCyYnBzPTyw5
JwpvaHrZOVTm65mXtwqtV4x4KhZvho0ESle3CWNQ2rkA2BsZcfU2OyE3fjIOhTT5
JfCw6a9vz4ujdOxPiBld0Tkm0wHYuyZPE84NBjUcQrBrmGomlEDoWqA4YjAyuGG5
yUPwq42MEEXBdrMDKL9rhYYDbjgv23lteIHDe6bP/HumxEcleTu9qpnfQ6B5TxYv
5zQ9U2CKiCPagbxk2iEeZqX6h7vYSW30GeohC/qWP7DAKSnobDuozR2gRYnGW4w8
yOSlG7FG7SmAq1PRK9s9YSIfYpupj3rpuERf4XhMQ/mndv85+5XnTkUHtKUk6Aew
rluK2p33PyO4UaL+1mlWR8vr6zX0zQnzJSDwB/p8KNSmp+dASaWo5xFfVHEwSF/c
GClWXuX792VXpEErsMLl5Wr+X4aNkX/zYsLZBmO+g2PY3uqRM2OaVRdErTUgHCD0
RyV4+pSVgYMV1K5gVLOTKTx3TY30EWq8/QdJEBPk5IbLjT2pdoh6lrdvHXIdk8iA
fLqICutmwBJtVY6xxlHHUyzK1JvBAbN6lz6BOlgT8C+DxDGzVUlu8bMi7YmpBpdT
4lZg+ptWbkoz619uQYBGIjJkjhaYnJjUG5yd96uBn3XXSRjIhi9hWw3l974A45G6
M0fL3YgWtrkGm2NIuLAFuHSvLtU+Q3xv31y4e0LhSKc8BuoqxxPjP4COx5AglSip
vckUmw7b/xb1NHJs3Iu/m2iet73eE6jLclDd5E/mjzQIyplAE7ygfY+7AUPfgPLL
DbhgrmnVy0cykfkLMVAXDYQ4sV+ohdrfC4W9UHz8eJ+DGqhz0Mf7sJIZtUc17Ci5
78Anl0JITp1XcuTPbAqBzt9JfaqozD084iQzo3KCCKbzgM3BIdo5YafK5vyDMgs+
2G5/tQ+JPPbicK2KOVoSshBUXOukc5jabRJrt0+xmmw0BIRoy4Pd62JLmHA08xdg
JctRyFTmu8yXzKt2LK0Av0PxlphEC+bHhHHpkh4IN0O19TSob7B18R+658us5VfQ
TlLmZNwg07G6PNz86vnkovubTvUp3/c+we9m5EisorX3mNlMs5F4f78EWKtVVt5G
Pi4AsP2n2bZuSIPxU7v4OyozvvqD+Jn4UP5n0zD2+lonvVNTec7wdVtJU815kuJv
l+MAckLf7sIs0Gcomu0MEM2+uKfrIFzVPLC8AQLmLug5mPl0KiprjCDA8O7bSq9v
7Mzl8xpu/dkE8X2/g8kUx7hvCqKJMH/qiSuySejgj4wdrmuWWXKIiWfhOlaJ00Bz
zb2oMhSrAHYKXyAFXGVFadL4SWZdzQKm4YfuG+R0bblXQcYV57EAYfw6m8ltecP7
MrKiN1yiDsKkeFay2fENWX25F9PTmMAicmSzQb51Nw5xogsF8UCBAHwpufmOzh+Q
D+ODX/5mXaqU+fRFTfv/MyEhzNb7P0wf7xctv1XbEixsK3BpXH0Dp2345ZZu0Jc6
EfkYkmQLL2z/Fxv4KCsyhEp14z1msOxrQ298LFZX7thUwsfsLYWeEHIKkWu3n+JM
/CocIZwKgXB5kDv0YxNTOmMrXNs5gFRard9MKckLJfib8klTsc1O1pKgAVtDi/8c
QGbJ4/t1JVvgMWCX8+QD6OPcJtvJGwLkJP6TMO/zjnHRGUe5ZEjCHMSx6amYmoO3
RJP6L6DXeG/+CRJjN6k9EqB/zVpG/Clwz59qET0gEz0V/IIYSKFLG2/taa/rbxAr
K/X5JQZ6IdhWsMnpo/d1qwr3NOU58NP2jhjH1iazUv4PrhQlYl7gzNgZlGiTE4Fa
3kMCsR2jDG1+UNvWHk2oW1By85kCd92o5PH+DgxJV2T6RsaHQFFGEOTFo/1X9RMN
DPyOmUEr2JEus9zpLqUybND+DFC8MRjyK0zRwOI6/4DKEOOntcuMPZ5+BuD3/UhJ
HCjLgWBSlWUbpGAd9+BBK0Ygt3prUbePW9vikwsnzAX4KhXju+dx/cBn6Ccc+1Ie
FcFiogxb8ACtmSSMHrrD+Rv1ckf8nJLXy8MQgMpKWpdQ5rKEdncP8ePgDvZzuujn
t/T/I1vGUSiS/jvH7ysTH0r9WAmN2BpLMIIqHaRf96RXugh3ZCJGw0e/i5fFECZR
Rrwu9id1diYk+EgLjhDL0Ss84DD8AJh9hzHO5UzqJlqpbfbTjUWVzBCdY7zcSkrZ
tPh59ZunmvChuGcxgFkIy8Og0ejb+PMeFtoc54yx9orxjlFIGKnbq4xK+GfsnMpe
YLKyUnO76PTt7WSlKXzhevAeYS0vP3wIYQo/F8twfGooZIB+fUso5Ekaofzm4/fx
YJO4EgTouYcncwQbLH9d2nFt4+dokeOCwiCR8Akq4TDzWlTWyJ1VR6vZ9MJQk52h
ZAFhEMUTUCDviKv6Ahhz/n9VeBxHCGma+ZA46URy+HmbKbnkP4T61Fh6sZkkSWtC
5vJpIewpSVSmzhaJr87YT/+tfXIkIKSxPNuIUS9QkfyJ79K95UOetx9DsX/Y8lCT
5vGVvhR5zV4Ry2rqncqwD4b111y9Xk8B9Hop7JGaVXP8NFETF2fhl9A1LszWDCj6
bQa2hZEyfHcWYqQ1vONjzsSRw0vlu9Q5xxFgHGGubbQnpvaSN/JacqH25Kiv/198
SWNHcCWzOJpvDO/wDRfRfVyMHTc5xua4hbYcURuZ8iDs4c6Z4zZCYpfdAdUiOTH6
6FF35qT5bAJpLO+PwLjH8cLpNc24vyo2eXLhDM+9V+zpHyckpYWrSPmZQ6Fog1gA
YGyWGid+yNIAmV+JxztdPJe6MQesGdu7RDTTI5SsHNXvzceiltLN8cWUXcOqJrHr
7638JUbDr79cJZh8QPPyoWTCx+v/+xSgFqqi6+KgdcAt2eUIqzzlCnUGAKX5Yqg4
B4meq2S2bmItH6sl1Qy9lN6Z/GfaOJ6iUEqgfGt/5r3l+RSi8sYSNXo+sMcJmClL
pTnGzanifGXOYfm4ENeqkIyOhxhQZELwRF0oTrZ3zKSo/RETnpI70wXINpr+qe4t
V82hrwJQLu65LyAkT+4LupDUn58NSfFGwy8OQqEP9IWUdQVYmrk0zHkOVuA4yTbN
c8bHscPp/4P1WUpd2yJz8i/RQ+MSm7ebLGdWX58CJwmLv2NIKY2XpHcuJEJJwo+x
iwPjZOVdUpmshXSxSyssXIHusIrps3yF9SCO0+LA+cYuVyshomUbCPY9ipXYcZkH
qBs3xOMoyesIbGcEatXfvbbFSGV4746cWVnTSKM7sclhL7nM1GyUG+mdTxpdOzym
CXgJdw2SyBnAzMSl54UDLif8bOKTPQtRTepSMJraWaaRpebnE63YYocmbEnqLbQr
buVVgkVqH2dF0iguxwCWaqpp2NbvqE2XtQLvN4N+mKBmMuueRE9VD4VUKtHQKRMO
LUY+JlKOLH6WFo7SeTJmr0VQ1jUWUNGGfbh1L4zGLfngADTDPj7AQginU+wbuLjz
yEwAckat+GlTmjMB5GYkFun3pP0Fh9cWxFQ7TUp2pNi//7erWKWw3Q0rf0qPl3YV
j3wUDsWHtnEq2R2FBUGfHy61gGTTTKpfOCYpyGXedJWvy71AoQ7PaGuhfpX+2lFx
z/+pmuFdxUh6dcKhXPoIL4BsQkZD4ZlNH3adgO5W5r6THqZlutA+t+5wlZKjQT+d
WAr30S5ZIkL2NBock+GFPQtgcZzNa9fH0/CyOl1X+8OFOWBA9cDXEUemilVHd3Qc
ONkbiGlnMfAbVOwpehITwy5ayTSSIDsDJN/Ft8FNYJnnOHtf65IM2ydJz9+qOcxI
RzRhRaaNsHAU0cCmEMsUJsXFA8r3vAzdeDoNULP1RMwFv5xG2HNGjYr769nuE5I3
9Z7ZtWvIurg++GN6sL2HwXdP/aLtK9BiIgrNZy+LN33BA6k3T/zjOCj/Q+OFs9AI
ApphmoIUwdou4xpj7dbENM0NyoFAu3DrUhy70ftg+GHu/a+BN9NdTXuWpx+u2eNj
XwBSw9IBGuT97SwIlucJBEwLlf7A/YHNKk52Yf+UuiATO5bOLwAmIThgTN283kfX
mQArADMxD4bJTrawmpZOkiEzPM0ijD30jv6dQo/qCWep28UNO/R5Pa0ZwTPurn99
8ydvQiqbK/Dr5bqcuz1vL/+RHSjbt48eQ8NH+hVapBW9aD27o64aEATkcfsXyYp1
sTNbpZ44WdSDAcBut4J0ez5LPGf7dDpwcJ2BRAjifnO8BIDYOD5XUMfyDUEa6eO3

`pragma protect end_protected
