`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
iuz82J5z3xXmTNL8LPx8y3ewN+jBSelQKzFQUr/Lc6qP6Rd2n0KCo+SP9stzoBBx
RRkiFbWW4wjcRkabfb4xX9P278ENtdV33GBdLdo5xPUox4gP858bRcrg6EtSgC5k
iac/anM6KvyQThBwW9r5PPlvHQrs9LhiBp0FFMJ5CS8=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 10080), data_block
CSGImvyfTUXn+AOMXdL+5Hq0t4KVKBLVrkentA5PpOEsrlCui/Oz4D9fpsBmhVNZ
by9cMQ1MB6Tyn7K1a3KEJ4fzct+ke0HSwySs2AWvDDEEVJdzoSIWGUjDeQi5KFEp
/5aW+MAgJ1w91+RC9nr+4YCFdiUqvEZZvCyLCrm0g1OGHleHWIT/qBPm3xn9yRtV
4CfI8iBV3YU9O0y1inR5D4NzavplfYe+CIU101UonRoOJiXAkYj4fWGi9wJft3Hz
tCx6zB+/J8EAdQ4qukrs6wWPfOXU8PhMmfM1O7/L5rNGsE7jVoLdiU2Y4LTz99Zt
QBv+S6kLm1JQrlFEUj+cHMFUeejsk9MIZ8qr2COfCAe7xCVG9qwuG2gr2pWx9dxo
nlcgi/HMNjip9G53uRif88Ntp4ev4LxeeAxEUyqywpaZqi4sXvECSMYyUD+Kv16R
8beJbi4NvCoK+azL68pW603rM0lEG5HD4YcrSsOkTl2jFIbuETz/3+RnlVYeHU2Q
oysT4+FcUv/8WogT9aOqGWy9mIeIDvRK/dyKR3XnJ4yiLXiJG4WayNO329b1FQIS
QZlh4p5f3COVXxYz2svo7UYtJJA9YKOIIZb2dP5nW+0xEQTbwMdUGKMY0eYOM/0Z
nXMCoKZZ1ooBmbyXe8q8fFDe2ZK31Rtx1mlKPVo++QeGOwXz+424JtOhwqAUM9Z9
T+tecC/v6mnyxr99NTrcOUe68B/LmQzRXtlmU0qqFyy2Ep4xc7HGQW2KSk4E8y11
m6c9slrT3kaAQUJu98dw9f5d2MPO8UmPnndNDxC9CqK9f/u+EekEmtXUWCcFk3yF
dskbRWr1V6n02RsIs4ecYwJZ5EKsXv6HS5gOXym7Ypdqxgofjrz9n8zIk6BiAgy6
gkJMedoZj8Z2GjF7yYAVicZjxaN5/nCz3DkkXy8c8Z95VRAtCkxjL9QZhoUqbfbj
KWHtmllAWb8JGikr306w6bTXu6lqYDDdQBS0UruMavlzVk5pw5omrVBNJfJYNVkS
lzEPTtPsVcyFh9lqCvjVNAIs1+cWJ+xhqCi4V/d03n5Ph5gDg23xZ84D15j3YJeh
nO9YuIuuOhr/evJ6DUiDktzomnyY3jOkJS6YHHjoIca+2CrVXZvwueEirCyRr1RW
vYS9hbtKUjdhkii+plE47FQ06KikHoZAf8wwgHyjFXtFNe4e+Luo+7IeangRtw8t
6kB/HYZKgxJANKKh1zXszpFjBTClLxZOv6XWxkxU+WzeqwGMwSWVA+1YUZB6X8iS
y+kCrm02oSGHJ/CGMk1wBf2E5RlZ/K3vQLkGM6L4s9r+a9/N2Hp3g4SPuNYl5tuX
enSaDsfeSDW71DTdYrJNaMBHTPkHNnWLQmH/x2ovOpwgckMeOimW8vmocr7sc3aY
1rT5npyqwuAfQPeO1vf1kZvaeakldBrWto0cyXNnTcIv6O2YlpC2fE99D9N7m9ED
NWqqz88ylV5ADyVpNeWTT9NTfs45sViulsnwT4uKcrW3lnLWpbZunIyFrxCLVDVz
ZiFRZNcVpM8+fvyzNwRp0nk+fw73aHZQ3M4IngkGPPmYi81c9XZ3jOTkycVCXjhZ
GbTZcyni8MGotZv6nyOB2XEHaix9AlRnmw3rahE6aQEBA6p3trqjmaQzOrlfFnAa
Bx6wsPRJT2Z9NCURAPBNsFAeBABVI4Mqr1nLy1SmP9iB6Mo6tsI+vch8IeQ0tqay
e8y5o11AmDdtVHqxZIvbqxpF5CL3u2CzuSIZ29VjJEWSE0sTZW9vW3Ja+qgkZ1mF
e/NVV5EghHycPnfWwY1bKXj4cVdDkYyNpm47DVw+pu2tF5pDIy6qNX72OPTs4hmN
tIQ+5BK3lA5+EbznrJrOHunjgp46XM95lIEPxtvoDuxWleUUz60G0FBsAjhUBk7a
VSwrxTLGDg2RE0edU+vGFEELeiJiz4NHIeMAxy/dj1fSolQRbRH2Xr8ytDuMYcAj
jMg8HFsX1kcKxTQZikV2R2CjnSuKx6S+liCwB1BYiOSWJ5oe5y9ds8W3mOGy4kKh
zhZlrpQjU2DdmyT0qu614EdTfidfZ/Z3EoV1zqjfn9KOFKTIQ8zskXWZGQzqLlG9
FbX9jjBw2JsJJDOZCLRG3HNv8HaeALWzjIEa1BfTwpH320ctufAlWa4VN/wLhcF5
RPjSxMSkB1BMWU2H9YHZxa4myiTB2hIVZiovAQM5r9jJEfnajxPVd5CfNyDNLFqz
rQiQr/06tGEXyv2gWkNa2mJd20PsKcFvEgv0O4bh+pMm/VTAv9YylNYultq0eru3
FarEt6iGQLx+Uz38ACwx+SNT+EgUKixwr49Q2PLXl2s39tnBpDZ5Q/rYGP7ClHa7
pHiGCKXpqEQfWahK+oZqlja/Z7651Kb1jbqhZy/vi0cLfk9hmpIJVZjn2FDskqHc
/Z64ieSylaVTBBQxg+LbTNxqwNxlczQM2crKyuKNHCUYiTybM9XvqbNpDmZ97/1/
9oz+OhrFejlMaGSw+XPtDYjX92wc+gTchFuNUYXdgZw4oYd7HNyuTTpiLCLdT6BL
LeGMFCl6j8+wQlJqoHB7qtzIFInQ7C8bfqatoW5daPqHpNV5L3aC082xPMKC+cjL
50C0ewxLb3+bg2bJ8fLMiEAbMFDYSVVkjkUhwC59EylzrLN4wP8GR26b1+bDrZsg
7bwCXwIrUjrWoPUdJd3LDI3Hitj4GQjdaZYKlX0Okmk6ADGvxayjtQQjSTGyLcsb
HVImlrzy9GD7y5wh/AbEIl5oo8geolhc5QqzPMXHukNVQfYD5Bd2NuR5NIzipney
DOsCE1/dTmk97ZlNiY1GwlHaUujVcNIA1i6J6muD/yLKqmmsIOUmnXDdHtxizYrG
vcSjUWx9GJmgaH0xdgeb2q/lQ+pCgv3P6DbopPVgqKU+rzeMSrlGHNVWbv+89Loq
omtGrUIneBJaaRQiRLOPRxFhVmFPsfwA5sQZWPmx7eqKZj3CPhGLaEVyycZh/woB
ksTWQsJf76By+aLS3nrDk6WNURDqHAdZDivvoV4usJI7PQA3xDr2xNxy0ztNvtVe
/fmdfhqy18fJbUmhHBq2XDk5VOCG7aWW4epNxCUvH5YmQwmdBV4tED9R6byrZmXO
t8g5VrDiwG5KGYGNf8QVgMNMiLghatIx0X4wT/8aZE4B6oqboAwEZqnXWAYJsduA
sCpMLQjW/i7S2O66XOTlPRCrQC4zpYXqsi+Sw8HtLFCzk5Pjosw6UYr01RaTfaDL
xXdzaBFlS/p66oBBHsNRXo2d46t6ORoTaaYmG9eDddTPiznd3cGB4OiVxuxXvA0v
mUpETeXxk4weXAhcSmv1OTRmrSryfI6z5ehMvNG+by+4bIzMg3jYfTa4vIhec7GQ
WEFqJPc3d3dmuRNPhbO4aTt9bR9vVzDveYBpTYtcvYlUCFfaGctxrdOsoBDefZ9S
0+m+AEgl9qajh98lMKvdlt1nDuon4vCP4eAQGf6kLrtruH3JJ7Wv6bFu2C+Daflg
hs1VVsJ3Y2Aq4xBY/V4fkpftQh251mGPkq0u/NbTPMQdAD/AZpitIyPKhoAVjK8D
cMBW2HTvrE9/B8bOnDeqCOMnjd9knthH4BSB8SU+a3o+lC/9HOT0dDULWbAWr7T9
chDmzX3AVrjQwhMvUXe4mIFgzxDK5cQOQnYEwvSl4fN1KPfgr2WuP1K9TOjCkY9r
jGcesXOH3eOqXPinXGcMB0CP0zkx/LmlD9EdR5wgw/wEoNtltM9jhClA/dnzEk97
tnSuPJAtrzsPdIKL4WIqaVIg4/Hp5wKjNoNDdqXRKwjb3580m4HblMu98r1EbEZA
dw8m/t+LHQALg5MexTfHfkU0WyjQ9YJ9eQoyw4KIswZ6gfLmry6NOmXuw+HLeDTS
YGrlbW+GKyKti9HsafTeyx96plYyPVJJrUNWLGydZEeSvCeoSemGJSM8nIk6M3h1
RWo4FGMHxR+jSptjina0cYjfLN6pZWMNGtNwFGW6HNZ1q7TF164dWLNCW2ALhQMo
V9QEvdY/YpMpWlnpMIwvhX0XgEFtGXNrthg9IblGSoG8bLcR8fPSxyn8a7FcD0j6
gdC/uhjwj670qtK88cd4B82XJyodlRxGU7i3YEb3MhHMCATB34Xha2ePU16/VVfj
BWcU9ReDVAAwi1gQhX0RDDvMuc/cjkiQ36HJOfQPaGeCNvGNDWcEFKKMhOubORKE
NtENr5zUxJHMWQlfRwH12Zll5uKWW2PWO29RvHR0YBrqEASmKTDsv6LAt0hAU4c8
xu8RY7swlOKujMPVoqkPb2oRTlZQDVf3XhYahmaE6w1SsZkaqBfe8BE6KM0qy73X
viGuidgUjNevE5MKuaNKur0rT3xmeIeKjPwH6FoEuD1VlCux25n0zNHFoSX6Zehy
/5ml4kJtaLEQDaiovHqMlGCKcCdUV79zPnrVzQC5gFoqRlXNl42JWsm8sJxAvUMo
2TwVQvxoPEqBCMghUuK0+mQUIZwAfTcAEfM64orkXxTHyN9FgaMUPeUZoum/+3ym
UjY/WHPkNqqKz1gTVypw6rpHkSbeBVKL80FZLOUwlCAkxQ3RTFxd25PE0+v8qXMR
M89waaDhzKWbvNI/aRy1OSUFkGBkYRbh5fkZ6Ir5DClwu0MVTMAyFPyMol4ABx0u
gdwexSlLhvnpFDjf5gnlPYlJlp7Y4ql/J3IUk/1qHrlnBXWfsL/4dHwUO0LZouJ+
2vZHew58ZLELCZ9LNtaEg6BdV79rbYgZt5tOOtizZ/kkWykvzNfk2kWPrEgOKT3M
tXJZPCgEz5+l8aClfWOiT9+78cE0wWnB7//Kga0LfCguIzdcDMOtQDIoeN0wWMPh
iKzuH3RUIoihW677N/UeJbjvweQXuN4N1/ssLZsGTaW+fVmnQP1443KxcSfZCjQ3
jp9OBQ5dINc5SP4w0wYqmRLwh4HP4vCiP6JyL75h7dyDYF3eZDz7lh4WsWEZDVSz
rvJxqaap3bn4CJ2LSonhLj5u8nisf9m5ddSzaA/+aLqxIIvqHxYp4a/dyicU4PgJ
ezI0oyHQU0KivCD2XS5sKXrxd+CptJTKpR27D+3wuIVc+4JfzmqP3BhRwDNDsgWV
Gy0HqYd1gGt35CzFYiOgtxDcENE6ID907/jJgxaSf1YEOwQJ1lX5yieqFZYaU3Cc
u0du1qNR5lpRvUL+3PbfyZYd7l7GCtB8DRTisOHOBbqKaBI4TpruwjX6YrUrB4XX
mcX2sBYx7GvtG7LVwx0vY9fxCZc9bn/XVaFryjkak/KcCHCOiDr9Z8G9jX/hCiSR
e3AM17t1iSQmWpD+aD25A7hIVH7vasn/ouDr++bMA/iitDYaAVAIn8ZsJQR4CmaE
N6nEqMOg5HQXGyFDS3tW6QszZeHTOXp5uc4buY/Uo69vVw/AlE9/n20aHcAO6acD
EX9o1rIaz/VQSOteZWYqp/NPo3t2v4OVeGsqidl1Ufigys/JdFJlL1w4Po27og3e
rmUVMQABGyZhAlXTM9MGgLYsji7UksRkzWHLl9RlNjlCR94SEFLDLJ4Q04+R4elc
jAerPgTd+2rrJTbjOFr5ZCbQx0HXM5dVq0tSzdUFmnEALxiiXGuiOu1B7d7Edzi0
WiIp6tlbhVU/+/WgOY6XOe9YokC1s3Qt5UFpUQ2syU1Lre81Fdl/QjedfXP/h33O
Vw4FNYaH/IcMi6JwL7U9+Qt89nJswFyP1hamnXcbIvoZkVZVXUh7s0NV3p4gxieN
OCopTZptO2wpvLv/xYdUNKMvW9CDelGUrfEh1EDbOBFVs/BFvz1FVz5UohEHttUU
mqQlH24ihOkoFe+GfsX5hCzIDol+F8at7EwYOKrqSSIqsrkuBVWBpriMevFkvIyW
ejajNtNd5j+uZ8nz0CRkXM6PENZ4uMXhVQC51QYahNoGPTMYY8ckYmFKw7vfXzNo
kE6fhRLuIt7QszM/8Asfn+aGI7NJgHOuJofoH2+6INvZsR8jcbUMoj5nmlaiG+mg
6tsxGbD5ysDHMU+b8+Kw/cy9vm4AfOnr2RxFycnnfgh7d15sUMKS4qMKG1+KeUt1
KFayPbXA14HjWvo/oKXnqGwQ4U4MthE+zXaQrz1gzqRj25krjSYePLDT4HnZZtV2
+hafc4LFo3FCiRw4KU6tPk0wtkJB7Y95bEMI1gGx5MshOP3J9sH0PLmExRp6BtE4
H7l7aTINjsQrwuEOiDHBLKVqKHFJpUHhhoYXd+Ws2+S91qIoamNTLFNnKzBI1zJ9
VjJhmQuGSjc61+kls/xxhRu7qPvg1oI8hU2AssOvAHK+PNS6OAc3xN4K0ET5wZv/
GMkGufma0nH+nWLriluB4mHPWWU274l5kqdOWEuE/NkCtep0gFTnEfgxxF+eDYpj
DMy9ncFNXQP+zeHCHQYNupoZH0rTNt2RjDMzLOIMy36gRveRghAkj6S657b3lbcg
x885lfAkccQuDgjJxI8kt5xY2W1TIB1QyE+Y5MW3iYIqzswrMMZ9Mtdlx7wWcw7Z
7p4xfqgS2V0HXZrBOG3ha05BAuEqs8e0FZ8BAbQUThDuqPQi1G4sM1GRv2Xp2e3L
kan6L8jERiqMoSuVcXEIyLUBnVE/JhfHrb3SqcA0TTwwLdWsZdLD424mePLJnzuX
iDJXIWhL6+OksrlP7UWJgps7cCykglJ7KQZ4wvMasYPO92LXzvl+BP0Qs2qsnTdZ
Kp9iFXkuN462X5qWwwT9JAvCWIWg/9ErjpzRvG0C3ScRMH8TUxu74c8ac17JkQKj
72BD/Ji08+mZxnJluocBq6jidpRWwcLcHKr6A9s5hdeG7DLyLQLOvu4vtnBeo7/3
bkhao7BED+NNRbjCJXjDmfTNiyJ4ms+SpyqxmU1OrT4VjiDke+FAEri9oaO4Fq2K
uo4ypyj2pkkI5KydejPIcdFoosMLZSmQoj2uNo/p4bR/EAK/yPA33Yhv7lKUZlcI
AgljbfLcxbQkySv+sJ9FlhADVwbm617CWDCu8e0VTmwaKumRONwfR1giC7SFFgND
zp5xD2g8urMOZ++BNjM6l5rxhP82al76duuYQgieb45kjuAVFKfpCRteRHJ0JFxP
VNHzZgYVR7/U3+PliJLiSEE03VHnC2oZwaYmHhlrDKSdBPy0/a76ps5YvwZBJcVa
77f/IU7pLd9jQ9XNzSD46GPdR3Z2RGIXIqYACpHp1eTc4BaZRZp/2QIufyt6fD7/
AbZPgL/F3dFUfo02uUG+gLQXuPP7+thQnmWlJ61izUNVTVXdGONNwi16yfttAqok
FFW31FLyGiGhO5p6TKblQF6+IQygslD2Uf7iT6Yf3VHrCLzPQJXtCb5aQwe52w8i
W/LKsILEXSdLKS5tppn2CIJnQil6DmgSUTUi6CvTTgEdM4LeeczDJOyL7EH7W116
SjIJxA9zfkuruiH7sSbTPxifwuv01N+KPYt0M9XhJWD+G1uGkQDuuDHsirmcskch
QgQsMcMcNpsR37d0ZzYDrFdhizqVlsggksIJdX1xqUl6vRNPwKhNpPimOf9Lo4c7
2JjCzhbBITAsDA9t4jqvdkLCkareE/VZ+dqRXAo1lFtmZNaIbecqO8P2HkpFJTzO
whf2ublEKWZRfz6qW692G+FR6BsmIwp0bUbK7lbIPt4I8r7qVa/G+TbbrjmE8NpC
fjO1Tw+16DcbQ63u/3WzSnz84UoXnAetZZVF6svOtZOh5ranrb+Cuxvu23Z9k1a/
MxlrgA7Y+stuVF27vd2SI/1bTofP6eOXp6HJZrWpvR3NrV0k0LTW/fjPsKwoxS/P
Hb8PJIFvXyNFuD8MNJoM84ETDR2WCc8R6TcYcRGKSBQA3Rgm6UiHRldXjPCIDpsL
tm2Cuq7xbe/8iqGXKg06YiqqLOK1KvNLLpQniV+OM2O+78d6cvbEQcskEGnqcJpe
y8VMcvwsKta3/Jy7OT//juAM4r5Q7w7zGhPyFZxvS65GG+Z7fJ5h+vdWujlx9rHX
Kqn2OznBkg3wQXSLsLfaqVseuPTUf1tq8QxElIPIhKVsWz9pa/gFRJPzU7RY70xv
KYGJVKehAMbWVq0xpNPK4Z8cZIL+hDOA77eIaIF+FLreb1SZ0m/Z3OQj5Yptlswg
x1Pz+ADOVtnueUZGVDrO8HEDHqGpbEzPq2tb35cnpIxK7OM1hEPIB0m0Jlj94Ha0
fNEHonMrOaBcvIzE2F9KYlaxnCrC0flfqG1e21EY3D3iNJdGj4TvZnHlvYGawd6/
8f4ZBv1HQT6O+yv6FuZc7Q9Zcrnm9rhr4usKXBV7MJib0Caxqi8NA2fLLjOh2Zei
HM6ksSmm0MpTNrvrfIDfZ1McWc2i87VfEy8/vE82swuOTL3DpT8leCvRTiZ2po5p
vYl238F0EDDlbQH9TXSXcqTTTEJYEt9SN5wvg5nNPdy8Yo7g5Wl4sCLXAfgyX9Y6
3xBLyWJeLTq2kKysiuf9iK6vdZ12Sgwr0y5viyAENpvweTFwHdWNnuUPCkeldOTo
4IgowRB6BalW57yv5SANIvHLry1J1tiV+En/8zLhjFABrCQT7GErkjYgKbn3fj2U
5+B/NvW8u3uWZ6RPS0qd+jrvNvuv96tq3RQePOxtnoJrXnQL/VjJ8l4uvVxYw8Dt
BkPfdGtty+unDjoNUzOzgTNvmrqPfCxAeVqhbnpktm66kXWuOT/nloErqPRf8C9I
sbHDMUVbjIrFuN/RP8LPK7MQ0/EYwkiV7wEGFkpxM+YY04rPmJumKo4XH4SBUhNE
vu/lyVwP9dZABkkgRSGHDt0L5p6WTOcQP+dbC8W0ViPSQF1sQvNbjS+oBQXjoMqn
NsZUCmfJz3Hf6E/Af2cph4IJAXSloeLenlJwBSdhALHQ7x93JP1ViOVfLEzSz/Yi
yjE0KnGHn0WcOEzay+9BXEe9Jj78mWrdMPGToUJ7rjsVV4kTITatQeUr1iOW7xJb
9T4VWKVcnPWqhELSTGJJXiPQrKQDftTZIc1cLgZEW+kXIhGSQ7LGZ4yCT+0Y+Vu5
U8sUzcq4tZv0nZk/UWiHaWY23sZjf+hwBh2albO8ZChzx1G6dPRhJ4B9ZO/Mbs4e
UOcRRHOUYH5cIMYVImX7Y0tNEGQq07UKhCYWKcFCgaN2/AGDUDOivl+KiYk9jxMD
HzkfRSD6FWwt+fOipw4MolF+saByPeGy0GyhNgcPA7DhOwnv0hSSNKLLcW15UiBR
g9DHQLSLpdR2my8iSvgojkqIUgdpOfo5YLMg+5iNvBJWtzQ/l1TBEFaVhuY54Ive
5n9C+N+ouHRv5tKorsWjj+1kTacrHWGFHMnd8Xaobdp+PThcw4aBmByzQWjq9L1U
UWPRfJFJGHQV9uIp0/L6KZguUEu5AiL4tqV+7cf/4LX+keuprXJqTUfZs1czuCDt
PRZtlyZtdcWjcsqwnRdT6zID94ZP7RTNS01eg1Lb/EZkISdsabrHemMkvkFmDZ4B
3ke1ATJhZBkJAQB0GaFB6043iheaePWe5flLWWsvVeXxr0fHwiAliIhItK5ctzbQ
3Ex7iI8Y4Kz/Q7+eqWmi8drqbYmAlst7nJYOounccsMTZaTN9fBogSMaOlHJZeU7
uXxxQscN8xHUiclO/HBOLsi3zoMu7BlVg+TLHI1FIOhsbt4q8cw0FU2FqNY+y1Z3
fe4p2k5DFPqeNgRFhFa6zTJzoINZ21dQ5VIqxop4qfgdvmacTiSG+FRLmYdKyooB
KEAntJr7Kv2sR1hbcldsSA5U1EFjyu95RSyuo4UhEJvDec4KxKIHNpMB5II4AtPr
O0Hplmj29GSL3PIYfDCBbY1FrGN9VszY7xZ2Cam8QFfCNcSNhGgKT4kTG1aueRWP
CuRUe4PwOxv8qK1s1vGL0P9bI5rSQmj7KWRPIYW8eaau5JNs+R4VHQF6METmY/fv
95vxhGYsSZqiKQzpDC+sIwrXYiXd5pty2Id8c1nuVZRkD3x2nlPZqSdZVdNBd4nU
pBOSs8lzmijhSFABLAsPzFem2jDibCoFQ19QEB8xi2OKPkXtDDUTTpWfAIshw3cl
gJFLs4IURCzdb2JKfu6/vKZ97wzNY9twf74K322pQ8NLJdv8u/Q4RXJVV5Ln8zU5
CScBytIp82qedEeHNiinyDmdSyufRWAMv8/Lt5lY7sDroUwZcYcbJSn9Syosb2zH
tVA0sXSoMiLTKU2HoIyZDFYnrlDqHBOTmA4C8bpLpBeBwYv/w+1miHNWc8uYwB4p
nHpt6DkkYOBsdSVRBCh1TKSfQJ8IQKIrswytoj7UJgT369N2Ddd8CiFS3jMONMgE
nm0qGqHjb6HyA/XvWJVCWCV/gyfHDcotaEM78yTWLU/6vBsPArIJk1CPGZgzPOAf
JYuaToCvhh60cFp5tsK1rgbn0lTbAOb6mi0cQzzf43p9vnRGG+H2bU9NOq1xsSxS
EzD9KZ9k5DhmDrtiJYwxXj6Iobexe5CoBSN+DTXG1zVE5WASRF0zdr/a1S3stHWS
cj6Wgl+zi2V9CT3WzSNXeVRGB+hbk3QLM6be5Y6aZhdF6+iOLTs/3UrjqHUdYOIY
mZHMA7NeKf5OUdjud6j5livlGHFL8O0lbiKh+VVzehhYHvXkC44imbxBqAV2m64g
Rjilv2Ysyw3HpFCvf9EjNcvohJFpC8y5N/Y433JyQiHy0EHV8wIuNVh3K/PyVaIx
cBLA/ktzovKVmeof6Ry71xW9qo7Cs7Dgmplur6J5SrY0AJYLijEKXbe+bkOWJUhO
MhMl9kvdEqw5ZNh/U2Uv2v+qr1uMcYbZSuUAMGA2RJToGqK7+laaI4ftozQO+m2L
YOgs/QclnVhK7SNXz3V0QiNEv79dM/nYZUK1heMou0XGQT1rrb0QwnPU7tvsdzYQ
eyj0dv8+EKxHHzsUktHZJOIlU0/2ivZpxptkvlHiOof6ehiokeqWtlmNf0q5LGZJ
A+/AQGsgCczJ+OkqBOOwHK/Hed09BPEAxmgy8k8c1GXUh7WFNUAXT7kbRQhRnmce
l6gaEGMPiBdWjKjS5s4UpfH/+VKB7c0Md22bSJo/gBdzKMZy1WJUkGuEEYLoRym4
KTStju7RAxDDnzDVLeEX1y8NsupS9dU4EY/Ni6wHgHC0RvjC4aKW30A6ruL/X4qz
gMKUsDQ17sk0OQdp4MzVh0zlSVB8MBWNQSLj09fdl1rUGlnvGQCo1CuPwj721zd/
7ildawiOPTbU3yt1AkR3nSYXsKSo+LuUmErz0PxAnjbrS90ekkwiVON1CBxxI+rj
wMWaJy3swL5miDOdgr++gIxgm5wIvOktOhcqsXD+bjAlH461RsbF+WJE5PVPwp7a
07axUZQqXNXf0uwSlg1HpWsNdv7iFOHMZmqRC6p0HX0d+ducYPwqu0U3tI8EMZNe
+nFFzWDwaT9Rl1+6T/l/zI6rWF0DjuSY+r0p7IMjbDmupIJlNJHU0KZbgFyNFwJA
8IL5xzhwIGCn4uDQf7hKXS0SmtrxbEgWWiQ0nnkiZtKvbmiM+nKxNg65Hm27YRCk
bKWcHESU2Rc/8SqdTg1yrfxC6JEcrRUJUKAMG4ovcQZ9zFHihtPTTFMUaLVntHxO
vDbdwsC82RJs4gInKs7YeXndOqY6YpwEdfFXGiqhyNSj4RREgvMYgX/z3PPmW4Aa
HrW3Rzu1Yp1bzO3QcOgKreZKEX4WCmF4TN0QHDkU6E8nSUtgWh1vbX8KP6uuBxJ9
gH8DT2dsPZasyAkhEhjgwm+qGpCryxx4I+sCAzbIzpSBcgQ4RUj+JE0TmaLwKJLj
PYTiq2wHecy0dJoxjjas6LuKcY7G74FsNgd0fNwOwIDm6aJ7Mulwcg86l4M6hhiI
f9QunSm7YnAc5M5jzB7Bm02pYdKMe1H04KZWCjW4XijS3B1YGt15V2Ef1CuZHW5Y
0yDxfPZsbHJt+Ieu3V01oj9C0na2CLDOWfL3cfkb0KS15xVXycyUa/34oq4uk90Z
GfIMjz2FfhTHaZo5fMGrWUQF2u06GkwZrgh6/ZdAcyNkA42yZBLcfnEGP4v1eluU
hv0Msn9wQFicKbw1bVOJ99XYCSQQXAgIy9RHXCdMK6Ea0IiM8grChL2uXrbQPBaj
nJR/KUYhIYbWLqg0qR0X8MT4f0+pbgFKXX+v4a45rG1CgXvDj2TzsqJt/eBinN9B
OIWWXp40Z/rEKQEG8DhQGAMSpBFSuTljMKJLpLqg+7FjvX18f7tHM3kGGhr5nsaT
QzZK+5wJfd74FBP5j8fBKqcG5ZAoKy7yVHMfnBSmavkBDn5vE7iZ0iP/o5KQd+Zv
k3HuO6FEPZtZsfQO6ArrfRfkYmQhTO3hgs4zUP6//JyZvZRcUjxF7uLHNIrOdqCr
MyeXv35LMZ+YLdTkTSNO3wFi4ogbdgU5prTP00kE6+MnIYK4VZqWE9Q/45bMnv70
xMuTe5B9UbuKr24hVJQwZYpLtr9fofUCBkDtV68yzx70yEYyKTPExmJR6mjc1uiC
JFHjnKzCKYFiAmzq7J21C9qz8WP8igxNxNemCtnwBFRJ2akXarT5r7zIwI7zAhcQ
ZnYZ3uLIf4iTyd9SsuwCQ539k5fhAWhJr6XFo/egxh8QS74HMJHY58qjzLUR2EP5
Agd9LwJwh0Up2A+80Y0GpcBlUyO5XO9elivSydS29yUzQ5wnckuFyww7lZV/uXjq
vcBZjGgLGD/FhZsGDHePeA5LYac/djLR89JBSBv0V+5iBB/u5Juqiq3E2Qgctsuw
OUbOobDq+qd3rO/VDmKIPp1CUmbuKgw6NML7A+trEtLMog/4P/1VbW7PGrP+RyB6
98z/JTw+y3qHHFjgC2vGWtbDvjPExglnMjlxyfYLdonuyhpuApEaxVkzEbiCiutJ
CAp9qlWt0+btgMtMlFO6Lv63MKHX0CtVEfP6VAf/b4DgskAbVL7kVqIFynb2Y3h2
1YjNn0UT/lbWeAXQ4NaESmp+uha8xdk/hazTNlgintE9cH6KHvYvV8wGUHSoXF/5
X9H64u4XjIyMw9mdwMO9lWjQsRMyBqhVU4A0JDw80g6HxNSAdcX26JWBYiNHc5GL
+E9bCYWXtBHt1gWNFRNfmj8xIdUE/jqqHUn6G1WUZDe9kDZyf78tbBstpB+b1ani
SFplzT+W8jFB1RZhOrsWkcucHwSKKcieQlDaZR9uZriV1XDj8bmXIaauK3jfeRhU
Vr/2WgffrpCc8MYqPZEbW2/hKh80TJMnW2UQttRYoN3a+SeHkNXWQxPo+3ld51Xj
1m2gPa3DHBoX2S+z7NNquwO54ApyH/pbCd4xw/EidRtM/w8rnzwEHcviy45+dgCg
rFbsX1wlKWObGQkcvJ/Ykp57qEZdTJHwelov01w4jxGTLEWBDAa3FUhXUfxihe5Z
z1/7EGu60ONY5OCGKrEzF+YoPQ8DuJtDVuyTSRedbIYXjZLurLeNlgf9BJJWeXiU
`pragma protect end_protected
