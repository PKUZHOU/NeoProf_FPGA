// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
ilEe+uFFyJ+NC4n/jnUrrfRJ8srIduDUdLPMwYK0kFmXoPzGmJiQD22IPEzzZjfs
llDf7A8mfDxMXEOhdzRNZv6TM7N4OcigQ9gq/Z0sT3IRNoghpVUISeg32ZCouBDa
gSnXXymrOxLg4ccq8eyab8nT5wsLcyF7CSoK4QLWVI8=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 2304 )
`pragma protect data_block
eMomaXtH4nAfCyh+WMabQthPgF3lboo5j0xiO7G5ZjV+aJjTMmD6IZI+OYY9I4ij
iUfxEwBy4if0f4hWwfr4ttmBT3kVzX8k/h5UHmbGx4UEll/NY6gijA+zuO3bJvkG
AOn7VKwBMBd86nZCiggwSFrlHZvBiks4msNbsO1qXpfq9nkOxVWGpyiv6yAMQ1mD
fk/5vh/O45OHtXd58Noj508ZQwICVzykfQOmTmQU9SAh7kN2dzCpWS9jrc8Gy264
7AKO6amquhPHD35++TO3uRO+utPl0YFSg3TJECu3OwbUrV+SqbuIV1fJ2LNMGL4E
2uBD7MWDBmFwsf8Lam2i6ybZfZnr1S4SZemqQ8C2KR+5D9g28INjd4pBmSl3Wt23
9/B9WEGoqFOSd5hF9PtutlYDcl1EBH4LyORoNeCNeRFVwQpT/hoWEubFr08GT8qn
PMZXcJg4V6fSSwIABq1PjhHyBKj4V2O61lh/GuYU+M33DfFycbeiVY8LI7ENO42h
vdN1Hv7G6ohg1d0T6nwR0U4mACpCFo0rLMR+GJNveSsmx5O8JyegNj6V00/Il6P7
wR6gCM3dOUaIcO2s4dlYyi3z9ahpjTAx2z8QjZB6pw4TJgH7oNJ+pK7cj9uU9edu
PHfaOzCtZlPnbiLtzOMJYMyyGzWr0cLv9BVmxKajkFb9y7GRdbKvczB2Xv3wsixm
TK6rYUHEXE01SFSm8pTplH/S2B++Z4W8BrDlsCBNunj2JmftWhnlW/srbdcyWZ/m
C9/MD2D5QN9CajyxEnNwHjPEMN07iwESdUUuQFQb6CCrsnefYVUjsSsBsuHHSEJM
LSytGMhYHwN6Me1YhIIHl+8DPxZaWr42AK0yezr1vXMaDE5nu+IFCA52sL6nNvYF
EdB++159Yihpzsl2VMZJtQUNa0fei04c7Hv0H7R1uQZFLJEGIoAGhHKtoxoYsxeW
E8y50CCTSV4xkH5MX0qAunI7H7FDpA2wxLoaUN+7q9kUSpx5O9jTddgK7/newvev
in4tJkDhzDVod+ScHk29+wMmU/DEq7LPOaUsF1NCpGvHmQ/NgqT+N6/C3/yZtU8t
M2hMhFyniXARyIGxqjgQBa8d1kQ8GDWL874IcUUbSXuY+9/zulyvi0zanzqWN2go
EyqKJYLTC4WvgbiQrUZql6iGuem2mSokAohCnaDb277m3sqwNQh5iFvGppo9sHay
NAr5oUUnPI+XYOjy1MCaligqWmaz0EbtoHsb61ohjh2dJlTSKPPDqGksMg45eX6l
OQSVKddqXqv2N/Cr6da6eU+GnSwgOtALX1PzTQTji5yAso9lhQJiUibUCkTPWrY7
QQavqErES6E2Ffv3c8ANUO99GpSYL6azaXaL72uWNHJuYA8om9J3NS89T0fTiFo1
1W1gl4zh9gLj/yEg4hwLT8zg0cUS6w63oknpzNiDEMMQVGcVsd3hH+ai584HvBXa
R9f46iJPp06s+9vFXdZm1IeP8cZAk0VOOapge1x/gfQHIj9N91sW+XLlkaUuv4RA
LGWaFMmTfIP1/M52MyJfj2ce3mQlQ9HC2GbHNaJ3iIvelK1prQwEnFsVvkZyPRzP
TG0GkCCUYhk4IsypehEeWYtwzHAZtLsac/vIyF/BgPcNTpj4NTc+sOnKhpkYWslp
t4v/YMCtb571UtYj0TPOZqfaXNjuRWIni9bEDLliCfExx87tEatNGvqwJgTE6wbr
m9Y+FpaGdZy+y5SqqtaHU7IFNFFMm80rfgqU6SOZNtZbPukQDxQ6EvxdK4UWUiXG
g79RabJbmIGWztG05fQ219HHPxmnuCcf3KLKmY7w4sN/8QD5VpDFqh8FyOs/YvKb
WGT09kPEMi5z47u1S0f0zPCuCUHgKNumvwzIU/oJZk++MI6T8uU0PtI0RYZkVHO0
LCO7zaa9cB7otxlpLsyUp3GyBPOUXSLBMzsu0YrWgw2zBGe91rHqwO96GPQiJNlX
MijXZ8f6ikc5Swa/2lycbQyIq1D1odFcKfFd/PNAUIufCb0gTpg2A2pL/W3LNwY2
2vWxUVC7gIJsyLMkpm7RrvJVxD5YhYVO2hPwTsgUexZ+QJNeoXsBOcB0rXGKIAZJ
8b7pXyfaljTIMLpHrkzo1CoWwEhoT9HehLest+a4PgE6ntcv2mmfv1XyWSjNUSVq
cXMVUH9iElHkdypZRHiCkxyTCuu5jOT0i3Zi735IJRF6EYjr9PL0krCvq0M8CoY3
aJKh3myyt8pE+F5TmuhUkunwYaGQhuoNplI9Mb1zrsJpuHS0wwTTbJ5e/5FqTq+5
fkC4cBQ7nvECvG7qcz2YsQLcfUrxjOoMpvQzqQgWwd2/XemWj1DLM5MxJfnTCgIc
07Drjr2T5/Zqyv63S4ZIRrT6qxKRP9ML1/AFSmcU8YofggfhI40dBgZ+dPMuPR2u
Jin37vCIQI8rIBMYcM7d6gvZMNhPVAhT06tZuW3mcJt7uH4Fu+1uDP2+bSlzUPWt
ioBfWAotE1tZr7qVv9b4hSdaIPRu5VE+fvxhXaY+6pvqv/VWkVYvtmvhoeNOqLQI
qKys6U+zl7Km3Qlue6GjvhuGoCPRRIXgk2ldQVfRBzlkHTJG1eRLJZSNcmOidu7/
iS+8t6eJpApQ+bpFF2/DOfGbGoXqb1rDbF2vf/1vS1bUr1WamZhRu3rqTg3ZWQAY
7jgLThs+V7d40HJwaTmPOxvSTDBc8PmK48AiDC+p0SPZwq8FnFWY11I+o56YkD9M
pCLpougCYRU/e0Pe96YMvZIvfFkpx3DZAh29irY6Su/blUyw6sAmbsUZ59OHVakk
9r/D8l3HY5CmxoLIno/lyetq6ZpActXO09wB+nmOwy5/JnjUrcs0M+uAH7A0JN/7
acC9B6GLT1CcK/FSCHKHn+HmVWeVp93ytokJY4BUIhWvbbgvtkWyg7cfavk+qM+u
m0v1qoYgimy/jP2mdQp7Mpu83jT9t4ZcPDp3pxHbA3jahz2dwhiF9Oljz+AznJ9+
V88Dr5stZ+sdAn84KA0HwhQCkrrO0NxxE/rrZd9Qa4vVQcrVbTuXgGwLSKqg+aOj

`pragma protect end_protected
