// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
GdXTdKDET6eAVW8K6c+EOG8P/6iTF4tEb6GJrTIphhsO4y6LkSQ5hSQ8wFO2
kgrWfoF5iFHUVWDEuo4HGBSRblqFwM1H+nZzVh4FHPwhg9K6qntCPnV+5dpN
H4EJamgsCt5us642isbSjZIhEPZh1584v3bsyF6EsE9f+srPsH98iJ0nDd51
RkWQFlmHXOQvioOCz2SvLpuMUB6EpNTelRfUxuBGua8sThUHJw5TeQRRrdG5
2GvdMfvNwPWUn4u9zR0lsDRKGClKHCBAY+LQR5Zm+3pkCNb4823SH9i03CJN
ZrVegHdrBYGUqr7MrHFyuCxsRsI9G7vFdYnDIYu+MA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
GjpxpQ2AQSwXA8oxNmp7pvhNUhY6R7ntksWVPtnEHX6hXefZSc/3DxcY6t66
JBT15CYGTncFBJNN+RMsHEC280ATl/RgrS050NkseTCFbZLYa5qO3RrMGEQv
xhxGWBWKvwuSPCjr97e+R3wXcJvLydVCZh1/0LHC+E/F8kgMSQpN2PEJu9ep
WIDJ2dmxOz1JSG+SEzGS6agoz7B5Tw03avZs33EmTEBvR9/5svZhAVmtjG2g
q7wAGv9ZxqtsGNbMGEWLdWBPZ0OwWeSMU3IKe3jTdFKvFs4E4N23hVdNnTri
2k8HGDyPggUuXWsx4xp0wW1wj5dM0LWLJSxlQP78TQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
fgottbW1pzsCTIuEAbHrZmKsswikVlroba8kaHWG36qwj8MZ8jtKIijpRsTa
KQhUw0UxvuTGDn+nkb74+BGyAELWFm0yA8tnFEwBDC8Sovei4OptiEW3Lc/E
/CcIdZ2vswqT4BsYLySHcA8362lofYehO34JrtoNJBMfAWbYfyrmkXa1ajnU
iwsywIpAa9E0V2kSEfDHa7K+hKRPaNLFPd8Ik5ytiYbZhObiMJYEVbt0xhFF
kiPEA2pXxsk713G/xZxpegqbTF6gqBPoQWaK4vqViMp0pz2yMTVF3ZCRaFPr
rIFdNRY59gF2Ah4vIfeFkGMnh9Gtz1DG5vzmBYbPGA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
RLZ0REVUKrNC4Jr8arOlrudYsj+MSi8ztYezpm4mU+85PbACtkqgf3OFkmkw
IPqqi+GwEy+c9rKMVLQMK2y8hiIDr7c4/yD8081QairwCVtnfkMuuwV4gxaM
N1DgziHBzw208GaQk/lv7jvtnkU3htZ/7wBaoYSoJL0QrcLw5Zc=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
sOaJ5PtMQmIUHzEw50jUn/ktgCmp/Pp+jodW1iXDuPNSaEAGSBZpePCizGOU
MCMeVUm+FTQicsdNV9Wpk9roMkoEzKM0f4gOgFI2wAtgbN583Szh0T/3e8fp
JlQCLiuHKBVlZxz9AxdZbr5jLuEfhgxkglh8EaiFtov8/H+Kl4gP8FQqYL1D
apWzcpxX2SwzUv1W4kyVizvlt4cf9cQkChdDBAP8YXiccZx+vE32EeV79OFA
X7vEc09CWxRnnSgFqjg4tgbqTwqv18KSUKgxiToWxF/vMtET7mjckNNtq3Au
uBaS+P6Q8OhdL8RtzF2FQRJlAGaqk3YxHiEh5bXXFMjAbuZORSUXJ2Y3ZxIM
7CnHqWo/LLHZ9IgRK5mEKoUCNFT2p2lGk0Geo2zZjCg24r0vE2IpMgMPtmJD
goiMlR6yND2eXjoOM+0P0KxvS1Ztan4np6nhW1+oTENVNlubmNfWB4tULNLV
OM6X/+wOOwEUxIgozyO1yJHtkgYX1VwT


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
J98xfOHM0JeiKhMsycNifbOV3iUGe2mpeQ1jQLgCVxHpWeoNwKY9EcBch+rI
Zexgc9Z8wfQI0eXcA69sZrfmQmn4ttz+bbq80sTWgkX0uI3lf776lCg0IFKs
KR8COulB0g/eB8iYweSt323CupsoTYqqgnBcOlPKkIfrLTnSZN0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
gBJDYLHuGFIH1DBCcTKjYJANV2axwb0zePvx1IJ1+IJouvOrHGURcfA44bKI
SRXjynTM5Gox4VrhOdHOZKa0sQT2J4K0XGo//pr0ZEBENckwNjxXxC/Vsvvy
QLyRx0YPqQhyr03FiwIIElSeTljlFzz/9Jfz1S35KO7bal7e0C4=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 36048)
`pragma protect data_block
eECKbMLe2SgTq9RQZTakk14eD/Ao95udd9Sbj2hHjy1ItJqCQg+tt9svGRGq
hzqVaWL1xvv+69mcNtdgO2XNqlGbZD9uNU9RnZMXnte/Di/uSzpDPCvL7ZOx
f3GNNNlcKBcMS+rJNJhgq7Uqi52WOeFY+gum4+c98YdaHroA7TL53IjJP6wJ
kG/HPAGWBLE7tR2qrtL+3iMX5HyzWOfzxo/cNb1v7XXqqkY7rNzqSNesKMEf
o3wYTWWNej3ne/Rsb2M8GiAHhBZwc1jCA8teq/XCSA7wlOeyKdkmd7s8JYny
/Wxy5IqJGGbvZOTBW+bRq9z36GeD6ETkK6QuBrV6/K/9vG8d0gPBYv5bSI5b
1128SLEBh7hrPz8PcwjsSHUs3YV0OgtI+Ui8zAtRThsK74/tnpQARbK1bT6M
P33chTFXMzNT5qi6h8B7gJm/0nDwbR9/gSBuy7LrmIH0//jRWWD75a7J89yt
0QUNMSzEie5WETQQv+k/hbhZ0XvdkoT17EtgB4ojf5wHPSYh6LVO9C4JcFcP
DPaB2xob8QYqQvCO+Xq+Dn0Nz1uIaoulauTfHTeRXal/OOGKc26yMiijzBjj
vQPMmAwy98VpROV5NpeUj5pHB+v7UIJrgSgqIyYY0/iHV+LwZGQ3KNKrs2ll
QlOpQAhi6hND7iuHnx9ddbF0mlvbtd43r0iK+qrdASErynl3cwdKlLAolilr
2zM/dHhxDGyPSFP80g+NhVZygliD/fbJy/afSpt/SqAoCm0dDiMopysCMRH/
kQ0HwhLeagfuy2tB0ucYZ1tw5UMzZWVPFs29WY0p2/WHRXLgi1ZnkS9wQJ9r
rcVXWQdjEyVAGTPlkvYF59oSkCXvtrOGT1DcWMM1E283uySb8Vd3q94qBJkG
seFNsmDM0JUJrJIqJ9DA5qtEbIP8+b2pk6KjxCUSlIP8aswWxn7t2bDnqXCE
5Z3+eE3emPDFOcqvS/opfW0v5HVPEiV1UUwYYojUxaZaUfZY/Tc/HBYygf+C
aAJ722qboXgbSUrMWgZjtvvcuLs6w3vr1axttveRvhBHDEwdjBgnJQCRyfTc
uifISW89PCu3I+IyXjx4bRXBhL0Gr0U9OD6B+XoDsgS+B/gTO9fXacSdfOaf
qb6ulLD+Tq2OtxToPv1hwywcqD1jQdTcRXzB0eChdiAAtil0eUwIifl1XPNw
hqzadDw6KUUtbFaceoVvoW8ehCH90o7Y97fWOb2Q+V/PNCV68fUFvQ1Nb4zG
clKHqr0L/Y4M9Brv8c+cMlvzCtgMXeZbRGz4QPs4BjtdMpY7o77B4z1jM85I
YfbGyOemRWXLD/cAkXOT5QX3iz5PT/qiQ07ZWWdNcHLgSEFRwbELCx5K37Ue
g/BNJLyXcGlpm3cL4s8pt+IDfA9rG2bKlODP+jU83QvUe+psOL0+zcvZvdE+
r2QEifNSdP0/w+PCptt5Zk/i89fapW5CtXbk+KefoBMzn+IqHI730HUxwavL
Q42yX/RsaVD+kkY0HOcqxclNF1PQUM9MQw0gPaA6NwDc4EgfvvpuC1+of1Jb
qcfW2gBq5hhrva7kg4+BTE6N4tJU4DwQeKHD4qtrk/4H/IoEyGCC48Qkn6xE
2ya8LcjYAPoCAWQH0UNeTwIIkIjyF0Age2GdxjHxWATE6b35+2hgn7uTMEqq
iJyTBdkuY40KXg80r9tSSnmTgoDNA/4t/9FCGHBY4phyTJmxSo7yjziXzVTl
vPitYu8kxDSEfdE/w6jm99hmrdaS2jeos+BLulLAIx74lAyV5LgzPhO7xRi3
FOZh/X3NGMz/mlgHJ/ARA+9SJfHChhsZ0KqPZMO3NSxb8FDGP0B6wv34jfV3
WHMBQZ10jxCFUGEN+IZWYmH6DJb34ddjZ86N74uTy95/FPxn8wzxw8Gbgd89
F60ORUB7YYoifUaca9KLSff9NrmNqipOyLQ0IjMhiWa0UHEdnZntSGi6e5sn
+4lOhLTeRGEgufhbBlJiPOMGX1SQROyCA0+EKF3T3JxpAVU9v0jw0N1lCEOQ
SCt+MgQIfzAMYnPEc55SdbgVmaYC+QIy6h+2OKnPGQsqZch2QXBGDaanY+kP
qPKIoTucpMQ21xpcichwCKGeQ0o31VH5RTFZPXjVmY+2QtEHfjWGSfdueS5J
wyVBNhTlqlQocD7OZjj1SHuovOBjLKMKYaDNMUPx1q2vMChqHAKNVqEfBBi4
XArFQ8C2gpafcQLVeM7dw0BbHz2ZDmG8ELA5nxkWUc0UuSJ9T35sX46vuVkJ
/X2VStetz1NScl/ddH1n79+mboDs1giEUPchIf5VPf6JGSOIAu6aD7IKWTY9
X5HIXx1UrnLeEVbB1a7NLh5M/Yub77OYHk5zlgiaIlkjp6SCOSLgM1ojyLKl
RBfW6gJIHg9yQ0563j5RO5O0cjqzeCJzvz+7cwEeWofDCN7O2jiYJBMjsV/7
2fEn+vIP/i+NjQKbz+6xyd5W4afb6twRrPD0TvwqLZ4Bkz/nJ+We0crr5tIj
B3YafTzsWUEiQN4szmg38qeLdlF9patpbv9fipIoL17GSh2scb2GGUGAw0oB
7guMCwa6l/5/Eoa8eiYjsKVUe5Z///pTNA4rqN3Ni5ESawc83X59NTzLMPIp
f6iW8XJwj6WoZkFRQZARNiShaYMWiRVusFZxIxuA+xNNo0UuqSyE/UfeZ+jR
BMqC/zuK2vsf12qBgGh8htUl1Ned9xr+MlXynOa2SW1rCfJVm+73qq2M+qp2
HgH9Fw4/kkRKoZShSD0jzYKTGsJ+o/CAwiZ9lwyL8y2y9g9HzwALe/Eqdmo4
/wxJotW60Wp7qconT+MZVekuz2vKmsqwb1bE91TliBGv8jvkFIdE1C+/ICEl
ou77d8ZQqGoUWk/c/O1ji8VA09Wo8ZYd5zNS36Pq+xY5oUbjZkg9ciXT6+Z1
H3NOyRJ+CLBYMWYVar642ZrvnpiJ2S3b4gdmHxTIKzakiUuRemAFCK1vzCPg
jsQXlVugD2zAFHymkI6vnbfOJWDH3HWBHJTIriWWkv2DHw/Kq9DAQtISmo8u
7KyhxnzqrV+O7uPcA0556/+Ad1+12wlfe1Dq2rxA66HWucijRLgjniVj1ZR6
BUC9CH5I7j+ogMML4/ACBAiSI/2+/El9X2MhDLKfwHovY6DyfhnfY786RQSB
UshbtFB/H9VcJdML9gnocBhLKa6xLwM+qzKnT7NvuTzMLNRNXVed0L48dI0T
jgXRgCv9Ln05SsrAOSP751mw85mn/tqpP/PPbnJS11cc5C+Sn39OrjCd4eMn
6ekV+hA6dESyapUcsrogQyhAcAvl5FL49jXD8WwU+q9zf7Q1CYrMSbctc+64
AO2QMrBWaNY1H68ZpykFseWV6KnhN9mdapNlHhRxGWsAteiqSViXey7zxH3z
19S/BEZ1nqtQ1ZZroMfbnZd/eQqg6AlPEIzY4RidPUrtHr/nZURQzdn5ivi+
Qh7vEEpclXl7e6CqnrSY+Pps4CeCQ1SMRLHky6CvxjIBRbyv4uSMl6XTctST
XFtThZigqA0EbYkO6JaDu8cjtjvE+kPhOEdq0dmmDtcHTLxkEsUzXofIjyWf
5KzVUnItl/mVVKveLF+QJtS6XTuk3Phq9GwUilhr2tI86tBiqXzkRB0HdUU7
vr/xlASe3cH1kD+1qEbaj6rGIW0LJHZRw2/gFKpUEjOaCD1oAvfduKSWoTiP
kh82hBCS+ez2PUyBsKh2ZrZM4sqEJTopQTzSlydmyxJphvonU7858ShwyFD1
6+nYp2awvlGkn/lKHktvDACXa+8F6LrGlUa3bH+SiXL33Gtgn027+bxyEi6A
myX+V7JcyVZoo0UOsOGCZfoLTYAzlMIMcyRKeGF6wYcM8O+f13XPJFqK0Jr6
WFMSeTiTzViXWGv/XvGLEJFYNXI6caN6dW8lKkKqkQdf5oa0iazpu4Y1mYO3
4B2bNTgzM7HmKAZISNoNzAwpzgmYthndjYx2tkOG7Z+QLS66zviPjM46ILue
JMCGYyk+48b0uuXwDn6f13z80oQ00/jcDqaU664vsDfNgSIdFS6p8XPe8CG/
q7n95qcz/WKryXKtkJ7tNuYWOxmpfsD8Aaymzl7qOviTuyuhHaWYml4DbdK9
n1ZW/LOKKosLuS5OiyrmP3bOwteFcT5yrbpL2zt1x7gLMd7zgYf8Bd8fFViD
rKp6IFcrhFjxeN9BuejOyU1e4FY2hGePrrIUPjbBN2hvZrQx2R76Mr+mnw8g
4huikRlSswxZdD9US3Dqyt0iI0BE1rfadwB8oKLON+NKMP9KZN8leEzQ8xva
wVjO8GZpjM7m2TSjK0nZrkW9bmFZSEP0iPW9Y8BEbVXVEaAkRFuLDFuA/mPT
JJEFswJy27KeZYPUBH3/DsIpDlRLo71TcZYLBzz5d8rQfTa3mBg64TgqFH+X
eRNt6jxdUKJAn5u3P6ABIyMZV+m4pu572M8SYXqsnxclPqgrjJIqvW2ieA1i
cAymT5c0meeUaGYr+oxbLIkIcMJdx6v2cemaRdL82mkZDXqMuCp0ZV1ADSH8
0o9Ag1Ir5z2RnlXOa8hwDrpSxCR8cHqAUSmDjewTX8T6JWgd0Yemmuam4tjU
2a54wJ9xfKxCqjlCb+cNl7TZdDAnMOfJZPux8HhQd6pm+YVvRjkegsKd5t1G
BHc6yXBy1v7D23XCix3miYUMVHLA+sL2LRNxHxphSTXn12D8hGnkwfig/wu3
JbSwyJAAu7f4VpsW7QJoGeN5wLo2MvFPQt/rsrBnualDi6+CR4AAqW1z+0Za
BDSlXj0GcMs4uKfVWNLnjwCab2m8w/t87XneSeM0p+UF6mhwhxAANj+TrTKh
VNQG94MlUfLHxbDvzr+JBq7BW59LdMuStgEerWUYMVAY9wTuyoMwuI2V7U0+
heIYnTENiDhYNUlfqGC5wAIOT/3UUFcOPnC2XHQPYi17JFPL0SmGyVG1UMxV
YGR7bk76YFbcSBwCg79TgDpn0xA/F5/ohM/hRZzg0J2MT+cWSqKPKdAD5lZr
wIYAV6QoMNQrmCIGwsgA8gmRvfJcPb5XT0scUMdLQS1GvsGXsVJTeiVssG4d
GP5rWUf6yfOqaSZ4nx1ckUcgFycUklHlniQaKyxRM3jZHGhjRIT9yreM741a
MWxzC2WmpuhkYtbpjGDsov1n/swxeSBcq/jZwaj3KY5bNvKj8k+1Ic7nupI1
HpCXIbZ3SRhT/owSOMvXM2irpQ5TasDM2Wd0FuDv16aaSxbcFfTZnXqfnq0L
k7txn2yzkdBlH3xTxZlkuLvvE74Vfpm/53VeEmk3Enqq2r6AR6uG5ek6uZSn
+K2aDlZ4Lb0L5HlT3dXUumk6XyfQ+2ufbznKyZ6FnDN/Dpz7rieEGAjdtJg3
WqY5R6aBOC8xTZjFprGfbsRbQFgei8cjDrwx6GKbGjK9GROSR/S8z3pxTb7X
X7SXEZwNaVSFRDWFWW9NdgiU0SjSCdkDoc80cPDuYwhiyQD9k6ujlgyrwboA
TM0bOB2yDY+aAHdRmGfEKm9rr4+xFMC+oQLGmG1Hw6wv6wLnqHu/Xqs0hGjN
NRb0eX8pc0CbXlUudPHgrWi+FpOyobaEEkYNyoRrJyCCVW/YgBOJN6H0T8J8
go4m28fK+0EDaxuU6/cnd3gQ3PFwzxVpxtlewR6smlNdNj7qxfv2rRhkUdm0
cmOwApoqWw+L/U0vH5fFoO7xxbCo43t59OQ131IvXDHeHJashl8idsF27hLz
C7DZ8CdR+Pe+J7ri8yBq0t9yhmkm82po1drkuYPuzDqHEfuOWX73BJnZMt/N
UZIzH2hPk0dlSX3wzK9tQN7yLHebQbVO2tdQrFTf7KT3xfOeVrrzZocI+58D
9chQtGp4vbS8WpTwNa3k3IV9KlF637alBoC8rUjWYnKZuG0LKFFVlBXUa1qi
d6U9Ik0WNwNQGR8y7EnJWn6Bz8MbiCSrv4otcLcNhyib1dzC1Duxb1aO3+e2
TT2SjkEkZ9mW6Phxs68Kv4B0cTS5alr14xnnq2hoW7Lq2C+9yqkbZElC+2xB
6SOARUCDhJJn8GqamqVm6HSZKHniktBLZUx6vvZX8ySQtQZIr0Dr7UZhEwKm
k9RGbaYvxQ86qRh+sQ2W/8NeX6LzuGh22gqOQ0q2nAUiA77mWaRIzXFQjcRY
1KiSY/6jP5lyq7TuA6CVhl3iygP81lLAngDDNlvdnsaf4EzT9XS4EH3ZD2/0
Gq6Vmtjp5Uv5wWF8smcnJ4Lc7FF8DvIfJ7lYJegWI+thCF6GHqU0KLRNiAJc
LkD8fFNuesoJ+TFHlvd6gqMq/AZpOcOSCGbGhruLAUtOqpF0Tw0PJtJfLL9s
EYX3nlBQIiMD4YaxL/D1hhOOn66HoDb7dMvVczaflHlwfB8WcxyrJ9+GgmtV
vzX0yeONbpQvqG2e59gjoPQ/dHZ/TWa0Kd1y9H5c8e8kcGmSrD7l12RajzzJ
2c/JmnyF5CAha7jvuC1yaMaKadFlODOkijG3fHZoa+FeFB4I6ij9qyAVyU74
od5hHVGiD8f8g3s5cEU5fqCkyBiqS1KDSagO0cA3vvY7agR16PZBbHpLJzgH
nJStGGdMzso6Ogl135N+8n0MRblPKiJ2vraeeb8duzoMWsyhRMkZfD5V5B2m
0durRVg/dYqSuG8NzoPggB9JIPtPFXMXbw1+mmU1sjAfVmhdPmS4HMqv3k7l
rzG3EeW93WL/urBqgO6PemTI5KMhbsxiqQ1BNQj6wuZTRaiKHln/fPvpg7hE
E2Cc197cNtTEZtRzxPWXYwvOLEfkWLl/1JJVbRg5oKtours48Da+Q/QR992k
LMiogwRpX3uG0tcY+PHHvpagu+H04n+CaWHMIbIGl210dPQHS/SL+k0W5Nxl
I06yr31SLs9VOlzY5dw0cdsPeslytcZzJ4MiEjWCS+i0qjJdkLpZq8hQqrpc
3l8oPEwQkDOAeZJp4jpPE2h2ejkYQM0lL+OhAw8bHT/ouSuNU9Eu9uHehos0
RvMwspJke/1EukKjFFW1k60Qu4XiKs81v3H/ibXnYsAToHMVK0jO/FU8norz
cEcpriPndZJwg/vZP53DM+sy2hDkObecbjlCzozumdR0p0nz3ZbdDRZb66Q3
93BQkn5GE372jz4rmOMnEQgCsjx2Q3YRjW/JGQB6kd7Ox6pY2aNgW2sL8yiR
oQqjL8N4+YCpykhd1CBMIR+OVGGLN2A6Ni5GPdBCUDoIBwx79vzLErUmgzbU
jyiG+lbYEb40TOBQ8b/mPt7X7lm9zeIJVK53W3aXUyx4Z3Pt7OYU7CkhvQpX
CY2DYd53QHq9Gax5dDo4UGNW2E4gnRNONaVmvorjKR7ugqM5otDT6Ul7IcKg
4KtpcHQiaPWB+BlWIpwFwNIEzjQVHXilfDQSor034EipWNsbXF95qT0Uypoi
HAc1Bx5A+0bjzJ3tWzRbMChMWBGjkTjTnlzi/5gUaBPDxk6CKmH0U8ZqWTic
5pTlkT+HFyho0iL764MeoAAacCOgKU9RlWj0eR5rIrk380mrO4+qe/1b+m0c
6cnuALXiFmJLhtE9yIXKLeaq0moeymKbjXWORC6cCWbVjfM/iyXC+2bduLBE
0Ly/YEdCz5tIATvtIIJ46bVwOhcXd+URBKMWT2NP+7m93mQPq3PBOREXDyNz
WGLJotHsnpzsQP/GEECdPSj8CTL4Jn9iadN80dKy2KY+jx1QmC4HAGDO99SU
jjZ3T1HAqPSgxoWlF3Ju6iIul0TRYgHuRZhFm1L0n5rDb2iscNFz3f88e++G
NQzajm/mHJ57YiS4dP7dYNesPZ3Pfb04eD/zrdivQnyxS8m4/JLDZQkMrQ+t
a/1sOi7Cjod493AV/vymA4B7rEsQCkMcrP7sZ1dZh1kxuNVazgnYFCyR5RyT
gSd6dQjgCKLR8VXPhfKR8Iogf/IfvHI66mvQos3ELJ8A4GzhHk8/Erv6qJZk
37YbPipA07EYZIPJyHOClP2CzrBRoLCLXh16ihBRPAoetm1KHrRy3M/mfeVW
Mht//ntge5KAzRo8JbGU89xQPzJRUH6w0kD64iHh84QseKmCJpQA+/RIMlCe
7dm+rR4fIouH4ay2KnQYXFroAy/O6L0jZ+Z+jaFPnbNNdaumkXCQMM/cEMoD
TxbjD9AtDx6ocfly5HnDOwA5ri0kb1KEIdV+d8R6u9assAP8rujkuD5ypEfL
VVFfASMLvTSOLR9aZzSxMuPHc6A0VCECxiKPI5PHtHqgMGdfXjrmGx8gdU+a
hrH4yd/3KFz09B10QxPB6sopBJu+lJt2+mfgqdKcL4oC+32/W62LxlWBpeBV
N9qbtZA674BZUvqcT+AScjl6rvK4JN4sc2F0y2eFqVZijIWDiuWj+pCBtAN+
X0ELdh8ECXzwjgx6QDncfD2jI/eg8R/BlvzFbtKFfC4xwPoWvvban8h904tJ
kdpxTcT1WdlDlqy+IO+O2OSOgi5/rh6wvkziQ3sGWe5YScz/QrkyQ3LOP08p
SZAXOBWnvte3QiOoFwVLtiNuQiyPXilHyymDvWIEKDwM7SRkdP7XFT3u+Z62
Z5nY6si6UUAtwBko0zw9qMs4kqyTo7xwtJqiyiugc3TUQnbgpX342WujH9Tu
u143wK30oUhK/wRZVP8dkX0yvqq+lI2LDw8rLyAyUruBkMJCYfgH5kKRWZHb
PntGx+xXLuFThEgtDdZvp/m7z7vVuGrk/ygOYS5qj4XHY3gQtskHz79PO+gj
V/GYt91nOPug8a/da5fJOl6eLcLE3s2kW7RJZ3Y5JJ4D9rHmSgJEjonz30D9
WrV/QFFaS0qCcqw4NbWBxTFjeRxrZL8bdAcD3w0Zrehc5Gx9d4tLzH/0PIRY
TRJ8q/7b1v48kHNioY8+fBAiDzwCzXEc48GqlFZtVGsQuxj2CmcTBjb45LBA
BlTlyY5OPBmSo2rh4heR9tiB9U5LP/iciU/z6wcj45GVD6f+eZ3lcsQ1+J7j
V0LazmvUMDdzb2m50WICXRiXKGxbu6U9WywwTepIFDPEIh+J/Pd53PxbkdeO
KY3gAmBQNFSBYgPr3i10rp+K6Wh9GFWzYQmtMVPERGuPpklYOam5ikJhsapR
TTc9zjq32Uia9o6L2kXQPyyldsKl7oQSiFaPrS1AaXI7qUIO53IYGBTW4XMm
f+sqgECdD3qTGOAJYGhwctp+Jp0OBc1wTbCZ6twbsojXibJo1FqbSJRTw8DT
AZSx9llU823TejUB0JMONXNG6sRsB1yLgcMq5mUX9clf1IZqTaZbZUOmOzHO
fGFK3xJi9pCMSzqjL3If8ejXURU4eckbRPTcM0vk/MWb6aJsq/SeJPNILVpj
jyOjVJOOlZgDoOFErJZfGn99cCKXdvnphaE+tQD51890tgzvs0qtkCKdcQK5
xpIJAZb4O86f3LdFWrRAdBXFcF9/Oe4pgENReGtdaO1lfp+3tp00+eccnkEU
oI/KeGBG1uagWKszBkSjqxZPBh9/RhftWILsKfs9C/Vh7bY9cF8+6PXOvUH3
iULDr9qjfPDl0sPAb7twaDYbDVy0+v3yg32t9BD4GDSpRhBVBvc7CrxhkhRd
ndPX0QGM0+NzzXSFADHYcdspEFQPzCr+vH/FXs4G6BxEw5YdpN8eFFmAY1S7
0fuEQuZf1Mq0L7rC01gTTN+Wd95wkjexG9ZXtnlf2CsM7mSaKyXCh8sc575D
M1OG54auxyqEr30kmPTCH6GrilrxPP9/8OJwv8BxAR4hr5mGUeNUGLSwToN3
Ij1VnOD7i1vlIkklNUgBexvcDjIO7SirSHIThL47GN50X+EDxd93hFe+lPrw
S+dKMrHg05LTrZNvXFhGJpLJGi0XbUuOAn7+IA4vS82tyd2xvG4coj6c1F+9
+njiZL0gZpiE2t7I84j3+m0oo24M8sF75W+g9VtU1+QJ+csLOz0FLCz8MRoU
1TAMrP9/CjfzYozHPKWJkkyfYI7T1bt37kS1pQHETc4TFP3rtBJ1/xIFlT5B
WeS0ms/q+zE5OKdvx4lvfW1eHZV9xhQZKxlam5aEQE7xwu2sjl2BpsDQ8xv2
1iB1WZT3IT7xrRPBUOqUKApHbhiwij8m6seH0rjfJCt538wOd3bGfJMye3kp
xTpcD0l9j0VC38v+YKNOCGDcwdCxwL10WYlw32+S5HZsBHYPNbo30RnFeXdz
teaA8vP0T3xd6Ulw1AbaEN/7EcI2RiZ2VyyM+j/KhqXGQtuNCLOm5rIrMyNp
JnrXtQIgGUUMXmaQYHVxrgjrb+hfJfJtKieAAq7QqQ9lwW/jAgiQvUijgFyN
3sxdQmQs0ngFvtlMVYAgU1fCv0G16HOu3ggpJAFQKyNhn50jTmW/8bnlOFTF
Gy3kZDivaThTTWd3tupZSgtU3xs3kHLt4UyCYCIAl0AfWnQ6jflDS8gPzL8s
cSBWY2TW8ppNsjyvJ866WQB+3A/RzqF6x0YMmtaN+bGVPZDqovZYmH7UtURX
JQDdZNkaujI71cqqB1ZeXAn7aLsDi2xnZdvBSSofYOWQwWo2qOEUmoyndyiu
EG+BgdqmpXvrXIQc/HDmVvEcFz3lq2E3d61IZ8h28UmTilUYPmsMxuLu001q
4FIRHaBUYvC3bLa7V84yyhBAcRngVQitbM2gddkz8tWaHjUrGfAiPUM9Grft
QRnTTv0VuZXahen45M8WG+d3JNc6X2qEympQfpucf7EmAlzn+jBoVPs8xFuY
aFBzc5rMz8SZzcSGfvEtIw9UM7SP2sOkTHEUpQKZyegVxaQo683doSh97ijj
czNjGGfYj39fXigsi/KbkgoiaoDnVJ9E43wiQx2P9MwoZC4M/5Fx6NoKkdfI
TeJ8k9qnXhqILq3DfBtdZBP3bvpRIrXz5OaPchLFr5cXR7Dl/8vr+soI0vZF
ERoKKe7qclWjtM5YPW3/ZYlhOfMyXi4zxxz5SlaBf4UBvBCD7OuA1xmkARqX
Q/pa8AAU6zuTc+MeCYXsInqsigB3pqZzMR5/BuNBGOZUC8C3qbIhqho7+2TH
3LIIs5A1MfiCx+IpoIY9x8srLu9Cwuv2WnlEOLtEZPbpitGOAIPC3zl+rgXQ
hynWxGMneHFpnEn40fBID4JyrZiu1JLlIBdSeIAoImmWYPQ1nsNfXnwTot/2
kW29rHYRSRT/QU5FzqEGpGuoB7/TkWHWYRRguyhtCxYh5Jn2cV6AO+4JPSb/
YngHz8p32aLBzlAXoi62TwDJv34E4aonhmY+4tVbN9Joea/V3UBoz2HA9ZxD
DAZ7eoNvHlYqeTpq38C+e8sdbc22iOu5mpsV30WprbH0Wond12VLsSuBUJ0u
ZrIyEmEUGmX4bKS2loUw9iOTFTp4eeePhCocTIa1qQOwEqu8KU4/PdTk6FuY
P31DkRSmk0oNL5rrRbejkBAUKDaJC7J58jE54AIXch73vxa5veRXnqAoGbwO
/Sn+QfWeF3yBslf8WHyhgRZrUPWo29R4xST/k+aJcON/UJupV69bxT6TqUkF
VY2RTRh178cFgASrhBrVIXBNG67CuH9yvfg6z3seHrwMszELNVEuaoiMQVYP
55/yQF6eT4FCJCyPHEkApt2ZbZ8bjoxDEibsT4GJpIzEU882VtrgF4O61DpP
3vfPMnUKYS7HumIxwicbJP6ChRL0/RQENrYJcaBjFlp/iVoR9y6pLji6xWy+
8RK+NWKpuvkN0Tn/eFI9uFTOs17PtUpqmzzICM8ulrFl8r1t3ewPlQ8ef8q8
1oRKlK/wlJ7ww58pG0F1LjYRX4cdAbZfkNkCCaEmgQuBNQ6Mr8ihoZuNPbhi
NGS64eiUdwfkzp2oH5FhZDRyuMOjGKuSc/BbXCxEDqXlbg8D79eS+qzpdgl3
F/fkD8Vb//nVRTshxmaHvlDnQk3zY8+0vvnnXJMcRW4fwr/v+tPmuzYV9fbY
Rr4yQGaNBZ5Mw8/bGvk+sArHv+ikJSdljjTPw6xgpDZb49b26FExm6+Y0uRj
6pu/mZofhIC94c8MPrh3Q4W+oOrLYqdG3cvGp3hj4MCnlU70PWoG4rAdSZOP
hLBVskdqZhUZfUtPGzNCtx3rSKipNFF8vwQvuMd+NE18H2oCooaLDvxiQP66
f+yRWQ1FIdRUCvouVSgIrQ+7IZQJgxdPGJ38Sd9ZXTPfFSQa5wJYfBHH35h8
ZR/K/t0POtp/1T67RMPIO822Dp9aTvNJrH0SbrgvHv3G31iLV1eQ47pbH/8G
jfRTMaGmJyxKVLMD9cj418Rz/EP+xVeAm4WMf1EDXe/e3O+WfT30CSLmL1ha
tSphICuQWHOQMEig1yRvTOgdDwmHzuALjDSE2MeCoB4DqQfTlzhr4f2nvC0r
tbhqXHou5/6MMTLL4yHLJdA6XqsjiYfkulsbvR3YLr0/tWOu2P17Se5zpu/L
G1I49QuvHVda5l/4AncOY/c93nkfoJ971KmtRGINTq2ZX1PyxynCvOm4JYTT
OqzLZMdiecFNB9Y41iRvmWG+oylZ5TifxapRzqQthIzX33CJcLPBm/A75mR2
fQpNEjZU7ivtjIqb/WMM76/dFjLteBbhnDzzRKyFxR2yz8KIusLspDzbLPj+
asLk9w7ESNJCgq78SxDZBhlim24sK89QdIccUp+uH1xyHtrsFQ9G/Szpl6Ev
vfIg9CsUERvI+369sRa7N3Y6+DgdVran+q4ULIuhvgfl44UEg/CQXti+eQ67
xRw+KMTwab8Nqh4/9SR52FC2iflUfu4x7/5+rYVWPnWXOhWODEi3yJqquRA/
6T4+AfjQEU8YDUa0aonD8CwqV4hD3AyDEdc5po4mqHQESPjZoL5YrGgSezRD
CTs3i5EXhaHq9AO+stxPdtvJ+HzNaSoIii8p0QpqCS2h5k0YGwW0lCFRkDCw
HethX/Lcesn8M8eBOnClSgUryfsCVF6WHD+26ncM1Md1PZqJFYKdT8Jr+czU
xyX21K6RhNAfnhwzNvLGPLwo33IdGbvIRloN59VJlK/EYbScvO5z49xyUsC6
AwOoSfw699Z7kVTwLvjmvqlrBtL0xJVAlTbx7sXrziegP+bCo4MsfTrD6DVK
KicFtNZ2iuJEy0JPYenuUJOvpkYw7fDx7G5GTD/gtfI3Lk64UB4m9uBgI7iK
IHUmURu8SPGV+N4/k9STu+no9wRBVhqyjI5bq9MkNb3VCvsU/2VcUTqO1If9
xphB/N4rz3m242+vjzCFojjZnlyRxeMf2kBnk3u5llECUaWk0LX9bEpIueSm
Kp6HftP1WdyseHgGtJ24BQfYa2yEeD4nkb8ERiXRwb+Ii5yr2fvA+gYzNlaX
PPjHlG9UMLe/TX7yYF8TJs5KaNbdUGQPtwn0BUbd9qze3LVR+q6ALP0pKN7E
74rnTNzQX/Ver/RnqQTq15yaG2EU2JSMd1UhjWa5BB5OvZl6J2P40y1orkLN
yKe+PUR609RK2dgbK43lkjrXO/+OZzRYDlWFSUFCpV30/F1CXBwXglGhNXzu
09Nx+aNldeHQmDuP+jo9LuFe3p2gDdpF93ISkyCHWu+gsVVqqVRBvyS6z6KG
QfNY3jiW8TpbTIxPHHjPKGEGIZLlHD/yMhgPJLM+slCBRO3jKv14wHXahE3k
r3JEaP0oZL6+eb5U2W2xSidfvhYziQqJr49spsxznmQH3U+8NmJKcIZwJ5wE
jSyUCVWmsUG/LNbbNlMrC7dKDUW2XYmWK4wf1ipcZrarnlJHT0Ob1cCAk8cx
4TozFD6d3BPO5bNiQ2UTgjRYSGlA2tiotXYiYTC/9Vv6UFJfRwdjgaTKZPhv
h9vSzkKm+xLFcoqcK/l1Fy5yfpg9gF/zeNsyWzViOthZrtIlpmq0pQTk9F5Y
w4KH41LNZBNlCXDrsXxHyN+UOZnz+HxDToeZOdiOGXvW/G0sGsDZD8JikG7T
XkJcYCB0zzglh9htpkv3JE6p5DKIL+2LJ8jeE+iedcvcPlwfFvV/MxFY/f6l
8dVrY4nLU7C1E2B+3Pj8z5ECDQI0g4ldt8m1qztsdUgza0tXRvD9qOUhvKvI
nyReiDn+mZ+EKkQbhJtXKwFsu3FML/jONWYB5hQknaMYdFWSw8b+jWwoCkOP
Rr0PDlAAssj1NYRFjbsN65/+mfex1+qyXR2LMm++NOoww46Y0U5tJKUTkI2z
nwaVyuObFhlCexRyN5x7u+JNL5oQpxO8y6ke5RjaeR56En7Q+viheiIE1n/W
8UJ2hCt8IJMitldnijWKWnAzZLNq0cdoV3zSNwGmPeGauGN/vicZSRB8BYxa
IK25Q9JJlek5laPfIO6LnOWd/1qRXDx4XJtBG6c0u6q99flQsJ5s6S9toiSJ
9E+GJs/k8wF+nKJqxkWUdC5l4qWUfTDRvc70jmUOW4eYuA78ATcIXcDPPlCT
S1aYjzd+4kuetMydfGe7TfEmSk6ZP9FjlBAE+WZ/qaCB+kBwlyd9x2t9KZ3M
o8pO9M23Zn5v09gkJ8gXbk9rbOQ4yKDhy8zohimkHatfXL5BF7SJEB4W1Nbw
wBBeIvVRTjOdzM7aav9EgRtSr8WjQNP6LW3u3X58U0seIhmTsIHUWvyinh+2
Ip9dWEwAjOHVvo8xaDtfnZXua8NdsuJuQtBvJduK1EjYODz3bbcZOgAbhNfs
2ZKMmCGlvA7B6bDRLwFmJusm+WOwUkzYne5gJeR9bqwkYssfZCA0ckuM4iUf
0uzgHbOb08K7IXlrguKDGoLWHQzMT/cUu5JYTPGZZbfxX2egTkRVYcCSxJC9
cR58DIW7FWiDw59PlQ7WM0xZxozeQj/ziPmcyUOh9ioW5VUQEx0H+TlhGU1V
GOF7xjKhnTUZ0UElaBQhyW7i5/DO3GpuuUb/zdYb5lvtgQVHggdlTpxudqS3
cngNffnbRw2qt1kmbYSMkuzKNhfZ+8uZlMywCv37OaNBqrZTfMRn6Ty8usNB
vch8fXxO0WTMxPGiTrjWRQAGDWkOH8mMjJEVaKtM8ftCdW2k+qJTATGeAKBD
2ePTQkQU10q5cxv8IBqL4zgmxK6Q6A+460vMJrNwZA51+y8Sr8/fn5nkPEBf
UxKmdjTRwAI2y91pFFB137kxIap7rcg61GYkPNmAo0Px/IQbeeYEE+ZPCvmt
nFHOqe1JFhjxMW7mOh3Emmon0TRytI5nXiTmCOt4sJAUeCwtUYa2hg1ibDAb
YclPf5xwNfTU7MCZXdelZiT2Dt/muhj1vjBYAA25Mm6vzSaZjKJ0p9wvcNgz
vMVlbhpq5E109+lQ6picNIl6rCLpcKXLTlQ7N7ALkLcP7gWayo/tI/34EtY2
qF/ARb2QWCHqXw9L+KjYGPzP16Gb7FqaE23+UEdaJ89srx5mnnFyOZbomuE0
Vw/ZS0r8ODPiVFTdx85+FjPe68N7QWPi6Wb0JujBVhERAsQG40tPCg9GtdlA
OWiqqvSy8k95/V+k9FfsgcXQWqFtsboEOVjeWrA6Mn2FMOAMyhfF8fG8vcvg
nA3pTfuxQGVFoj/AKprMiTVIvvKZUCKifBG9auUg3jEO70tCOcTzEcla56xl
1vdNWEx3doq79fzBHGtk2cUoXPH8SC5ndpeU7kid0jLM5boevTqmnjlECixX
JPqfkadQYuX1GNiVM0Sml/a4jL9KG4dGYC/IoVTEocdUnGbPa87O3KfzWTiq
Zq+MdmtIcXxHY2zivIJKGhU0lGlAznYlAlqI6vSuLSxHNta2qR6HGBnB+6hd
6cDgwTmy6s4LkD3ynabeL7zl8MfQG/kPaZLiXOkjw4UO+PZ6b014T+AXAE9D
bZYjvtO2lHNG4w6Ky7zOcsfMAjwN4XLiZm8/yR6sSkIwpTxDOCDFvxIIQgN4
baRZwcL0lCtA6dhvHc3a8DFH61flHF3lvFD63lMLUJYcdaQ/yVdXijE+nNSv
Vhpx8MKKPfiUz+cH0+6OiY70jMrFfnZH+g2PB+GZc9TiEzWtg4CdViZIKVvL
0dviWQe6i+AUFQRXHLl3xLaG2fWpPQjS8pUTs+vlilZv2UTAxHaW006a8T0i
zLi2itE468vGe6WWYrHrPOXiqG5SlgUyjY16aR+ESuH8tN5+dQZRQo/5zVIW
OiTPU7WaNbXyWoTqQzAbiTIES30FNIU1Lxv/qE0KQvq9XfI6rAA7tYvmmAw/
TFY7TSqYOp46xaV1M3eWx1Fq65fVrNy4g4fI/vaCNEf1oi39upcpW0anU5UC
3ox9x3Tmg2rZK7JctN7BkGOBDkA867fg32Tc2WfHLDFPxlpX5PcwQlZSdyT4
HkdR5i9UZSq80dqDhnSh5qlieo7hbGUhjvjDPTSFjkkrbG636I2sTFEufRGE
W0nauR+tbanAYWSqmlmKkAVbFddHEpxlJ54SIbGiWYP7cbjeI+2UAKBXkdMW
ouZLCm6WqGJGP3FtkgxF6YFlpDzXV1UYm7VUjz4cQdJOMYeMvnyiznAkufrH
1jqbBomHo4LLHIwOboU5FHvfNZG8qT+IC2geS30txm/Wu/gK/BhHUu74Kwp9
5ctveD0wuNOallZPpQgBnueGP8CVMCcHZJJS2LcVEatEOXN2KR0NypJdgRLE
L2uX3dlaHTyfq2bjwP8iVSP4nLhAS9h6F+efzKHym8fIUgQ8FhFDp7DUA+Cl
7fyc34IK1T4Pm+ZUU9s2vFJaqpsSwe0dyg/jnsVrYjBmtcu4wJvKcWqs4fxS
UDk5V2tZ2lya4Rjcf+1FgharczIlKTUoypmd4qwoWBJLEF9XKCyuzUOq+sfP
8aqx8cNH5+8+QrLDhEmU3gDj5Dju5tZMSZyUcLNhiqUpPLeDXbDPV7B9wQR+
R2308anQkvk4ECS1+YSYKRoysCSnJ1rvi7DFUvABdnjZp84SbbBV32iZyLko
I2SU8gu+LXTAZuyPST5ycqIZXMjBVcu17i8BLHRiP2mUudel5Xm+uJ/NGovU
9iKktWm8isov/WH2ZZQxvlsHVUM3iZ/XY87DzYX1ZRgFX3zWjHd1yqurhRuj
fNGBv1MDKaBC4RS3VyWuyMJhSNINSUatqyOPUGXih7aeU4uHH+sGFqk8Ri+L
8tlMalu/xDk2Ln2FmUToJwA9pF7BC9+mnbN5wHyaHHyrvXUtzlKQ1vX8ajws
WhOJxYBd3lm3HFQNpJzLrGTCgToU7wf7/SaUtRui73riyS2y+J0w1zPQ2GUC
1prtD1foNVLTf8h7X2OvdXKKIchezcEwYhWqPvmJdHom5qaYetKCiXgbVyLP
wz2ivVVT43OLyUh8z6XzK/WYzXGAwJYjLTmrjQTimBPQwlrcbcXiurYNQdqj
RmVTp6iB2vSsqz7UQkr6AaoXCwIeOApsuXlvzaajQ5cOS+VGYd27jny7A95v
DMXLheF+lwdYeDUe19VsfyQw+5QkDONGIGrpxMhrkRu7OhpPKSjKGrcTA0XX
SCXk4MA9kHR4il07YZZsLesMYqfFxCT6m5oyYs/ercyfRmAH2wKr1Vf53qGi
FvVY6MfyzlehoYYLlMScnaQwr9F/rEZ4xIKUXFCn+iv5vfsoxpbE+nGJa9i/
jb94T/B/S/WKInJjbyAFLpd89RcRJHzKmWOtPSPmwRsBVSboss1J/Kwur3dj
qtFPFmWK8U57850Glu6Soaa3N0fSRQTLTc7bL1p+kPZyXWxokeQSvGSXg7dh
2clNnzXuA4/1bhXs0O9hzq2KwMLRVR6xVMV0tNqKR3b1Y9w3wdA/HuP2A3dn
kqhlrVE/eX2Z/FJ1X9uuXHbnONJwzRz0gpKsJpQ1SKjks4RcDYuUvwxjo+7X
jo4zp5RpVLBn5i/vJMghYkR9pRBWDzZ8998UMbp3YbwUo48O3ZKuqW1SaWFH
GiuibfoWpqOUXUmRZmvw1MaRpxLN43afGbVw6SFHrD7D3IPDV/Xw+8Zeztol
6Xk2aMJdo18J4n4jJyQY1vbxjsLYFEAdW/+7+6ZJgljcBuH0+QYg7S1d76pq
/4oWWeBygOiheBcFQ+emFzNwCoWUC+MVsh32sEQEFIrt6p+ZKaHJW1+JVvei
22Rz5dge+3ZZk0xY4wPPkxTzDP926g7UJvr1H28C+KopSy4U0DXFvMfWorsX
BOs2IGj5TuidthWk/kvd/4o67DBrjIiJk9XlQ0enTIhXJcvp2rKpo9NoT+6l
toiR5cF8fgsPGSPvp4VQO1782hQyHztu6Y2TCSLKiyp2IhUCvZZlPWn+YV0D
XAF+9Y/SKKmpp35B5i+/MiD5/ho0I70bmHW/r83mxRUxm9IEkDMEMU6RNjbZ
pkLZxlmC16EG2+kYkG/CPxlSrQCHoF279b8QnSKrvlDuMztNEnU0N/Vt+h9f
PtGFZvWX+enOStZNEG9zq3J1p3Uj+PWlb6Rud+dS4+42aOZC1T01PZpAyDcB
88VBNaY8/Lbf/w9YKyai5q9tqSxQo4uZ3SRtO0rKHmjC+nz4kWrtbFJzk0HR
qLvwzimwMtj34IWcpSchfZpP7SvogEfdMK/HTQVkv7QN78GoaJDAhesaprOX
tI9OZUkOqDEIkX7/5FtJFAZpZrAMxOsh3jBsvyLixHwKIaamaV1oTT9aC8hl
RUjkYqW5EhSwZttqQm00wSDTf63VAWm1iiPZ0Ln+Q/D0R2vYQ11yNvK3/ZqX
kFFKdb526FMqzeu8WdhLvunzEKIJIvZOXL8gREpRqxaQz3yDF5+UdQ0xZsqR
WD62w7ZLTLHLKDE2DwYPWyJTajvRTYM7yfmdtE6Oe1Y/ITHaG0EVaPl8n7kw
dqUbgerayJALOJADffzyfblkKabIdtx4kN2bNW+yHn4zq1AAhsXjusgLAlsR
WIoC58TrM2cQiZvTx45+CkGNjtADKDh4e6ZeIH34fr6BFK3t1PUHl+GQ18bE
PzMDP06dIJeZROJc4q6y38APU69xcbmMfkbT58faKW6pboK+tYEwjhZDuYJM
lU5GBPcNr4nAF9LFrsTpG05DpfCuJUEQFGyple0SQxj4XXh+w6IrCHcUQ3Ul
rm0m+C6AcoL1NGyDrd62WatXI4HwPdAQtF1gnpckA4EdRs/wygdItocvbNKZ
5PZ3O0gRPN0htniYLIbVf7HGl0wjmqh8eVw7EV6wI3n9yk+b02dyTaK1qtBY
zZ1r9AMDJEwLEhxMygkTVIOLfRlTfSPfoK8yPK2Vruy23CoOVTawj61vzGo8
3O9G5anuy61TqE73kbMBxmwkkFzhSm8kTp/83F17Si0I8E5axnSOw2HzDj8t
L6mEmPzEMWdtNyPIj2m7AImyrqsrMtsuGlx2zUcFx5LZ62Ep7JQHOxAyOstW
ONIC29YD4r8mkQIS746Ylv/H4dVcXzlOcGlwMWfRHsMAGYFwVXqaZeGhMMiz
cT438H+bTn7Lj8TytBtiINCYj/GmrerX/eGuyVvVbEUv/XAS1HAQgzNU2mlX
Hd18C7bIX89q3/k1jKmcZDTObL9Bqbx6aeDNfhcnQ13CTkaIQRZQiuRA3wS1
4xfsJ7S2HvOQPtxApZ8lNiug9bUQAKCs/XcqYs8yr5XgDiFuvVDMPOUtZBcA
6yV/i5YM9TcDE73qI/gZGnExK9guP+s1sVekuKgcWJtnHMdyM9gUwvyfii2v
owiUQJwvIO0MxVB9AYviQet8EyaiwluE3mb28BR32XFTDq+O8NmYJl+KyOK/
+RTeNWE1hG0Zdl1WEVLdiYg5ARXZXN9yaSIlXwn4ng5MoKZYrGR6QRH8CnFA
8p/CdcP7beMKrO8VfcTUNkn9nOcPmV5ua05fEUV48ndCxDhbydNguLWnFF3l
M9elyQkQlioCwReV7/Xf2IRfTwJNdZ4zxCGRlE1JhYsAZSMJhJmKikCU21lL
Y3amvh30GRQy9Ig1defM3W8i38MMWD5k8Ve/gIBuMeF+MMRPkvnv5YoMXUHQ
3CO0gqHTeaz83922/JO7MOJdOKeyejUKGz1S3LEQ+LYKW6j56KsFW57pZwTY
2+yuMZZ8ee6w1EyJO6Xaigw1co4vtGIEmsX/aB+Pd4uyg3S4ctbDymaQapce
49qM4fvr4tY120SDfNMIjdH6eQDAqt1bpx8AnfsRM6cEH0hnJ1ch0E3PBahB
sGH1wnA8XoQ7MyVN1VzwxwvZoQeW4PwTwnWOQV8Yz1z0/ZiPMfERk7VnE1Jq
6XDU5qbUBq3W6w3s+FYgq7VDnAUYtEqkTRLJ0evqSL6ljsLmR/TnL+goZiyl
IDUXxF5KReCaMt2mvdkF1BowsVKgeqCA5og7DemPrAIonNEOZvSdxifnYcYZ
DX31BRiymp52SxHtw9CEtdkd8r3pTHWI8LaGEP3wVosLo/aVh2GrFwRzGqCL
ezpp+6Zqu41J6FChcDF4vC1QlrZ0Bsunw3WomLmXxZZ8eDmTFpx8q9NSOqC3
Ogl9zBzaV8mNfyxQRBsAyy9vKURZbtqv/m+INZRx1qvMJLcv0IJvDHl+TX2e
D5ih71zt2INqzXZet3XdD/JdOuf0XtuvH/kTaDxO0jluGsCFmOHjfj4I0gjJ
Gyr8AsW59ucaUSfF2HJRPH7qR1SQ5DmnYRY9BkKL7Kx+vrt+wgn/hsPavM89
cLBFB4F8VpLdl9tMPRMzv7rTVnXIbHWd1QRM/fIwKzRGMuES4+n//sqPphaU
ohNYBtlQI8Wpr87PhB6hHbWSdVwO5WNkFRXdkPqHh9nZLlvqoMxq1zNKqGlK
/7eF3y8m51UB1NSkWJIE4cG/pLn3WvqalqPYLndXCN/ca56AvHSBwdA5ttgn
4qHxnRDif0v31aEHNdM+yh9Ezh8oHjIiZu68nkmtkixcQJaa+FircpsIyEga
TLgGIWAki3jrf/NRUjm7G9o/RdRuCe9k3z0CrxWhPzh8jaATrxF1ZSQgEQb6
XlsJdMr7qrZy2RVFxb4td3TqVOmNthjM8YfGwIXOcZT34tdkmG6wk1sxmEw1
OWGESoP/2Bto87KF03vgxOIo5KNaNHmmRZTD6vXLgZetuKPAopGTAB+o/SZY
JsZUIg3amHh56ufxgpepN5VkFZMTedXcl+T0LCH89rbfQSOZkFnAhxfQYoed
OFEu+jmFcbW/cY2gfPs3eD82V4a89g5Qigfby4LnWRYBifkhi0bsh1dR8jV/
b5NATUY1tkVMQHqQpzEICDGXMJClGV8t+NT4/rDd+JdapgYbzTbj4jRODs7+
eGVK3Ggv6QkIvbv7VAjUYB1lDd3pYAZlT/hGc/gwQbpA93nFWG+QVYygZXqS
X7wxgPN4JRcvFeCRTE2LQccc4Mtx5U68krVaCaXUm+Xykvzy3eomrFbcDgvn
SUcH4HXEfVqSOMmKkIWWxYalE0Hf1fi5CiEc5YFx/bh9C2FN5R6lGQAyUPge
2XY8XDf9g/a19ZuUCTZBXHipNcElSU1OU4m8nqPvS3rgBMFgbG7z6a2fvraG
O4JUErx8FEoC24Xgs42Vcn3fTcBvBzcqX1Fsw6u3xpu1CxTB6o3uBELNygAi
ozimjfqwS6abQ6YLfa+tELOe7vYFOSRoMRJOshbl0fZr73NMMGh/pjlvGTSJ
p8iVF22JC4/a1Zesjlp91WzxwzGv7K2QN4+KcMmQT+mSwzPL0L+kR5vnyctj
1h/wTQA6Ay90PpTJ7H6ktXL95lEnKs7ZItLZpJNGQEMMWQ7ErYbIT0rQbIOG
q+vHPJD15smDcq2iM1DvS3t140HRVbZOeAEqnScnOw6cxjcdyc+7pwHtoLLO
9qypc9KLpI+XSjBVBvyrTI00Llh/GW3DQc1zxMoFAv3f6aWkIBqam8hzt+s9
goU6KigaD4zAeFoShXKJTqtdGCVlHPS0KVhH4SHZoWF9bJKnvBZkwmiAyg6K
C+AUj2LW9ANjQarteO8TGvjZBAvNEfTq5mKL77p2IjXpZXn8j4v+02jEgosg
THZcWDctyopQvg26zQ5lsRj0ay3ZIf9zdDvHWxz7/xwnDQx+nhav68lKAHw2
bQnMu2tjScw7kWByXPk7nbo+9JZs1TeBWRjudXc/hUzxt6ojOXulQuX+VfkE
jJhX7nsSLd9bkJCApPZiXoh33e+g83ElvU3ErEzlH9OPXWevwu03wqNf7JM5
hLeFXq9yhRbEJ4CoHA0ohM0GiEmMOV4mpx2JTiHFtzKT4J/J1KXbvmst/IgQ
S3LxY1MkflD0AbTKTS4rMFVirtFGDNP35D9+mgzj+vnzBPby9MMskiLurtkz
9UojA1RxEePaMzmLYze7jyjQZpzipS/It4+B4au8U7RCWvyK6CfPJn7X+1FC
X4rlm5e3Bhg/oBduRSccdD9iDPto6aoz2NzFfs/lhJNwYycOpz0ECQSDp2jy
36rFKXe3gbd//VzEDD/gVyDLgRQCDJ4oPDh1Ll4uZ+/4G+AiHqke3ijjCPtS
yu1BP3bGMa1o/D7RZ61Q6ohjBT1uUVixM8BwsrJ9AsmBBZRFJKihD6yNuQxF
C04fLFeQ+YlM3GKZ4G3/vWKhVAc8LwPlpH5la6TERzssoJZBjaGAgltT/5Q5
EqB5nAeAHMtPN5WWlzTmB5ZBN2yCzAwqHv4JzfwqewAZKGXQ9POBkmpNYn2m
68TWYkSFYXELv+XsXaxaN8HmDAXm5Y4THGy4MHduSYXPEiO400KTZGwGXOGr
8jfRHzYUvXvavZJav1MUh9eEUEYNoPxiNcFLVrfLEHcT3HF15zkfgRSldeiZ
zPgLa4w/Sp8Jzk9rTq07hflMc6QzouFo78Pya/AHLiTxpPnJ4iDs3J71WR2I
Tun9mC3OU09+/4fDTYiftw6f7j1/AC5BHfUqQ3Kjbb//UlByfB8yVuTXYy3h
aJOxat/LyngBrFK2PZv7iXpxxxnlPg84YI/npmkuMfCCc2dyPnhSvWz9r1QM
CslQeSVnbr3f8jyB8yJypecKdF1tjwfaX4gzlZB+xVCQCzd6TYZFqF2t2oID
UfS2kYyaa84XayjyXh6wFfuBKoJlULDyhhrsanzpGJHsH48ztxZCtvellbP0
eCRBH2ZPpdT4Ld+mE1Sa1vNZM8r6xTyWc1D4oMpdWHdVMFPM1Vdu2A+OGAZ6
obxhCS1Zwg4NzKjBRYFBROHsIpry3d5xBGfTcDN4THjBV1YC0ja2a3Rg18RO
mfMrrTm7SFeeNs5Nw5TK+B708dflBJHAfN00dmygcTquImDfV9h6TVqacwCW
4deUhHPpbA4pl3hTJeOve1WDnI+oJtVQOBZ2S9zTlzGQFmh7I2ryjcW3GoRU
TuFQRv1CDyJyd8xdejHC4HdnJPaELnQrFUlruwAvIKa7xH0uMRpMK9VdmJA2
gEGNHfd4af4NJLuBHDSnQDbpCgscHQ6eLJy3NFt+AHeavT1a0lf1I8m7fwRG
nCcYw9bQMpqFsp8ZjuO2etHDqUHSOKqnx1+5r8wKyMkz7j6WSFM8oE0ryCy7
wkPHeOJ1/9z815aITqwcUCe4OduTU1NILqEqe2bTyaaYQ9Iswty+iFT9c4C3
jRbkHfxi4Osp5CEhekkmITjQzJO4pKFv/QmmpWWYKql1QiQm1zn/d5ym2Yfw
Ng1qDOOGo657RibVhf1vXvL2vliznANzLdDHquG5TIPJLxbw3o04jgmP1klT
vqNFglKLPgsVDBRUloaDxa+bgqw0NO8hOp2tuIUUBbxLKLLZQLmdxEbUFpJL
sZttPWptzDVb2aqOubiBDqsnY/0xdfVUcqbOL6PII06AZCWKQTtU9XBMwQ0Y
mTwD1ybYVLw1mejgavWkTMe9bSUMHvhtXD+IP57Mf+hPij67HvddhLzy5BXb
rXdCzzNkiA93wxyXEql16IzJN6Lpr3fjugqPmud2RAWQQ1t8vnPI7iVHX6X+
otjQKMeys1o3FVS/uFYVcB2tLs1I+FJ5y8SP59DHIz7LG3sSergEsCb+xQv1
nIOmRt0Km4KdEUMKdHga/O7lpFLdZHoff7ow+559N6bED1yFg9onJmA9GIvn
NxXqzsfMTLQgWRZ4uhYLSQ/mIXGk7wiJ/1v45apK4RLTYwb8w+uJxgSIsREM
vHfZhF0EbLNf6PQJAMpruCIpkL9ef4z15ArMKMWYla0DOH0LhVsNDz2szvPn
JFVKCLfA9xQdrS6DzYbKFkfe/ZOFYzrkOKRJwoP9TmPGCPwEvXjFkCD2aviZ
8Fkc+FL3msoMxjG+/bI06Sgi+aJp9bXnTMQ67omg3A74nv0e85S48FRQWIqy
wB+smMek4HavwEFmieB+lXcp9XRtr/noGO1XcUjthA6joxQbVEzSFxhmrjpE
/w0YT/5CpgBNeHC6yDx4JwSnyvIxhOaeA3QfO/zytFnC/OJita06qcLakodV
6EHMw5pA9MG8m9SaYc9EZqsti+L9M/abSyrJx7hwJKSEABfWp/iFB9K5Hc7f
b3b72czjUHWHsSBfphq1mz2b5M5ldVamI9AYGfuzuVL1DbBmZMSxx42eO7hr
WAEAg8xpZ7WIQPo/vtgQhbGGf88FI282VxOU58kzgIYQKgGfEaI593hrAr6D
DQP9LJzkyj0q4nVsoc04JVUnjFITOBBcdBgVWhu4DZPfYorcb6hTVp8ZuZRR
1VnTIpdWwHGYLPLkSz8jCP7XACh7UiofiZuuQl9BLllkvrT/TDHqoDYyrZ6X
LTAnpGtoiuYm8w64nPR9mkQaV9BlCVCWM1kJdesHtz3C3UVEW2o4/KGT8WrC
wSl0R3YUFXYMYLIIaDudlt+/7vVcMyxaeqVQTiwzoFIBLDPKwza943MOcSBo
9fk8e3usVrL4QyybyVzYeyD3bb4fsbYQxmLPWscRoobltz9CEIkwaH1tCwVi
44a9hrcUYrAtI+t15DQdHqfwsNUzwok7TIdDA2PBU2iUiLdnHv8wreXc1/8I
APGcI3y9pTG9wuc5YWxcSYjrI80JvA8IkfMAX5pwo8s28jcEvt5QEls26P2Z
ujU77refDuRXMsl9xZvaA2F7EhQONbiP5f3wrQPW5MQS1afZeVh/PukpI30K
7NiQfpRp0Lbicg+wCSyELf/EkncJQWDgueqOHRLIFQcodG/W8kG1OjUSABcw
imr4X48yKLDOrkHhT7NtYtuVH2DG8V5ebxvxDsY07+Rs2gU5u/OR7BweEYzt
9zHMONNED6GCTu16tuiLnnYVBPo2TgYhRaqfXi1Vo3GjZecYiHSXc9apE+T6
EbYecCPqFhdV2Y20JeU4uHdmAkkOZzJPywULAZ6j5JMwwOPqIezE2+DZTRgw
VmgfpkpfBpJ/T05gO5z1OXXWxbNXdtB5ezSL/xj6vcxB6O/FOX/TWnF9J1W+
wmnqY3ptnBoprMXtyyQ3Ylw9h2fOmADLSBdo7AN/VC/sIJTnA9duRKHz8heK
htyEDnGknlR1sqjn1BVjhWnwF88FGJuuxk6QrGXKNAFEtcga5F+UdMPvKXug
hi7F89Lxg1iMUfUE/pb8pzyxxAxVsFk5Ln4aguzm6kbsLpBxb5clbsalUa1D
FPLsPSIsT8xUGXHSuhHUoq29viTXW5+T12JhVXMl3RhXjRRXQTnIu3+8jE3F
lllDWyjSlOs36wEbme7vR7ribW47FFPO0b5E4Fx8M34FmvqSmKRiyOUwpYXb
1ciFR0gxfpEBF2vWPO2iOah9YiQwuME9RevoersmxZhxYVmCH+YzDqE/MbfM
jXOZ/AU9EDs4srSFxejKyQQn/CpSe2AaH+VRldwCGHH3uR5tUJsSljWmm9pL
UjubXQZeSJHRQhMFx1upxeOGL8d0kkjPTbSLUrazl9f/alV/RbmNmMWGs6Fh
tlay+yInnaVs+a2RfYgmM3OJfsze72MFe3jveq2cPRTXJw6emIjt65w4bfPX
Fu3TTqPto2u+dbvElrGX1MQ9Q+jcIOfYHRmbcAUyU+tODCI3qMWCDvJqu1+o
9vUs1xM8ozrr4TRp1on9XaT8Yjw7hw0AKxYY3wtC9R1EfEiXpUs8mXw88IWl
95jwzo3B5BJCjE9Xit7dDBdhF0EmAecNA6FWFWQD0+zwt5lYQ8Az8zoaWa2K
1ovVKwIFe0+Wq9wvL1YaTUVEti5MRdD45/BNbh4Jz+K5JFhMh/TGwnCB+8Z9
Te5ng9ewMv5DHtY2T9H333I11nWCkmXVzij81EbHF7g8wyE2zEjGT4hikRex
gROHz8A+d04xBO05kV3P35XZqeeZ6z3YnEyKeeN3b2cj2gWk6ZQvDiMfrDb+
kpFC+QnKkVrMFqY18qkD5FZDm8O/fvnVjCRzP295tlrC6kdBMmBR6wMYnmHs
EhSMBjWiBS9VBhqxufQvJJMfLAER1of2ZRLMiStYFsXpsiOeeKMNACk/Xixp
zfkRXilWwLl4XqnDBkvPXfpU148FBbiTXFcxEEvIObjv0+7QozCRxoGbkQuX
76nej0j6PwoqlZAtLlwpD1c8fiArS/2QCf7mL0+rpbr6kCDb4+9VO3bvc6wF
WweuVkOsmjxxvMCeOsyzQqEyV3+A8LrmHCJ5FdhdBAx++x/QNdjuHnfGABph
ITkuTN8otcezJCwhwD5ZJj1tVUpGDJ2tC9FDRVr0pg8k3zmmbFSJcwedU7hm
vlsf7a4oVK6awGm2xjb4yl5ij+sxLOU9G8I6sclL4eFvDTs7hY8twZPFqrTC
CeGMQHZie9sjzZrSG1X0nOc5NjWKl/iKPIwfR15Wq37JcY/hb13hbNMrhk2Y
DdVbyu89txrl20Ig6agx3jdZD289V51wcb+Xqxt7iPUmIEOryZ/vLLRQHQbn
543s++vvrnooWmrNA6ZbzvPfmglF2e8nDvrygf4AibcYQFVkBzAYElIoNCBa
Rd/upZV4STKg8BWPhnkK9o3IH78tplL9ntAlkIBHNrUCfDRAvQF0auDOdzce
TxflSdlrxa6jFnSK76t6nGYieGYMrvD7mxTUK+zq6DuJjJCwpx/5j4fNngyv
UIHNXA+oeDERBm55qCxoaLt6s3F+Rynw73UcJGCuWBUeS3QlPl3dNjwfd4GY
sg8C+yGQLfrKPNr3Pi1CpGNIXu06tq5p+Vq0f0cmb2p11G7YzF+9bwOaov2i
JE0aey6nEqydfjRG+FvXR7tZfxagNfo75zqUSNEHfD2hqQB7XJvJpiVGl2Y+
T+CkhhGVkNem+Q0YWE5pq7vlFcQ3lXJZvHjqYes+VzVgWUEOZKuBLABh4BEJ
rHxjmTkOX/JIu11klPuxllho75owyJtSkJ1/Sx830pJDFFfGTCMc54kqP1IV
1sGaNLJitM9r0A7aqm8yljECgghES8BbBIAPT4E0FyF0mH6HOFKv1sryVub3
ZmCifgdvyVOiriVRn8obti2oFVNshLQsxaABtsdbTBbAeb+iSkyfJkwR29UG
IlEg09sGYwt7E/jyayXb3ifHlHYMkaxECfGbhoTaBid2mfUkiv/RysAri+vs
UPP4QVOW6q/auT+ki2stVbnk6f8TthjDWEAe8FPLjUnrcU9R2eM29jj4JuVN
BjhMCyUHvJmoL14edYVZEIGGET5zPHwgfI3sFwwM7qc7seQPIl0N679kDbfO
rvgxBrFQqCLJlfjlIuwI3VN3aA0uQHVUSPHuzzo/zLrC8bl+fZNJjuF/7vQJ
DufPqgFZ2fdFVpY+xjHM5C1spwwhndbHyXjAkh1ucQuv5h1agQT83QchPSb+
914CqOLsYB0EsPPh1RdwA+t/KvH0U4HX/14rAcB6wpZ/BDSa3zQ5Lxe5Zb4U
0IDtw/oqfuaUP1jwt061Mr/5jm07bPr0WWMEQJmhGfxWxMN60CUIFotZH8Fr
C0PEKkPVev472E5VplYsqEeXxMTrEAZ1DBHLdy3kJf1pMNseRlOjrmvE4g2s
s8TofPntFcwMtPcDAwFvNDy94TUcTX+KGDJGGSqeuhm6M31ujynmvY+qMWlY
5nybD7hP5HwR/sHWfnz/0mMoq9yEQmQAJVoWhVXSd/Ku3Hjk5n4EN07HE9t2
kzsZjvsGV9VesfCiHGwDUeNtgJaWsNjKOtwR8y6mjrHjuESawv1kTjWM6CWG
30K1wtNtrVC6Dmh2jEY0eX/SG6l4fR4tZebdgtpyzAWT0m2M6nMhedw5kNAx
DGPrj1XC23+rVWvrtsTeFMWBtogT7ugzCWq3EKRoEAm+VoxFzhQkgCwDQn/p
q69PBsfTTGvzfyFTNuPmvbtrouP8il2FhlUmiP5bFeHB2feL41E8U0N9myzb
gxbCt7Xq/FI+na4RgtoLiYP2+8Ze6diTUPJbpk8+f6oM/+VcFqskzjmZhG+i
mGPnp4x7xN5yFz4zVR79ze++DurdvrDqDzc/oz2A60oWKQ+8W43WW6NA54Qb
LzRPXhQJDiPeMMw98a+AUajbQVj8Gb2+DpwBray3TVSQRQzY2t6uwDzWUQK1
QJoocyhROlDNlSbPYjU1XBBH5dfBE3xQ2tbbvG8r1+coZitnlabaYiPWo7k5
9Qymcxhiy0l+lZiS2CI6zMxu7gUnAkwJvoF6Mu5BK/72f84EpAEXwpb3VF4A
LlhhYEaJGyoRUSuNDAgv63h19wXLeyusBh/uuVsru4rpORqSZAGH6QSkqaYJ
u4rCHQpFkr4h+KrJ316SpIW7RdeJzc5ir9u7kovBgxFV6uzKN8rKaRVm+ar3
Q2OTnZiWiHH+mXNr2JqsZE1C2lSRhkivYV4kf1v9fex9aiA0gUd9AJHYkFIW
dbDA3h9LhrB8HcUVwV5JT8CencYNUk0DV56A8NTOkXOVzrReXNDpgRWscWyY
PKwDA2a+Wp3eLIxYxLu3riSq37ZgPd1eJNg5xsC37xcRnPbNKJq2GMbTN1Pm
0V+hI/nfcpjYOMf1dcEx/B1XyaCmQFWQuMi2ZUdxfuExjcKKCKB6vRJnpliz
R96637kT6N60Mx01ekmicOru5CbN9iVtAsWT8bwlLYjM5wAb/v7SFKkwyPq2
fCEMeyPZ6zU3x62W6Emj6qiztIzDY20LiPXZGR0dm1GtrhZMiu2QojaeYUcD
tf98DxaJkMWdFKv+gOtUKc24wpt7PtZHMOd0X/CoawgjaCJOWSO3PPP2KTW3
oULa+4foM0RimuSY432/kH3j+KgG9YmQqyZTwOO/KY32+7f9YsB3+FI0a1HL
/8oGAaPRzWA8GlCx2J/CDsGIFGWYAZHuU1RGVglglyryn97uqwCgrOXPa15x
/YDrzoK5qI4jXHSND4gxqTyAckSl3UHj7fuAeBy6H6ss1OmTjwGVY5Vqd7Pv
Mi9EWEcnxtcqJgEmtrJFuj79vM7j4bjYl0piC7FqyHBXw+t1ibnmxBGP5CAK
nX4xdAKkPCCGvMxCgS8mumJqDO1enPHXQGQbj22V3rovHHbSOTWHVxw+vNSf
rEEaDPPwyXOc4yn+SzjH5gQmm5uMEfiNnqK2VwY6MpbtyhqJI/A6Eaarc0cf
HlEzb2QfRPdh1K6zz188e+7WQgQwbiWQo4hVDjtlJlqWNIchozizr/NByjD9
dlYdlr6PvAzCGcFXeRS2nVb8qSZaD7aiO7oJ0XibV6URGBOc++wLxRPc20dV
zptkdgmq5qx6MngYFKBO5vAXq+nWdbqpbI5U2QVhbpEuijAJubPblWuorOWx
1tEH4Tq0SoMLpzr+c3NAMJI4wH4tt6uEokcQBfzNvbmNPNomPBFiOBgGTgWd
3H+v4ZK7E5Mu983b1oZuRMtw7Nq1uu91Or01JLHxINdK4ldMpJeDZZHLG8DB
KVAAr9vyb0pzJ5UCUEWMsJhPlMPXQxgVmTnyBUrP0GCcb9N9JWbqEiW00ilT
Fp3H/1oyRk4MQoAqY6W6pHZmfOu6m9fz3HqYLAHC6aQFop9MgrVoGxTks7WP
9L/R+nf5M2IhU9APjGRwiilcrY//+GjZUY1luDBZzVDgUWUbti2bHEvy4CVd
HFOqqwXYayKaXLjMwOyRhFx6VQek0sfiPH6fBNsiwEnvL+bs0sAv0MRxEazP
Iq8EIYr6/+fa6TZ/R1z1cYSbuXtUJs4lDyP51FXaDZhctNlrDAhj9CNoV9LB
L2sBHX/LZ6A0ohPCv5x7BejcBbaOxj/oF0MS8p2W0h6vW/3nl7B+qywVMgpE
GVYWgvB4QwJaZDbF1pKolpOQ8feH/fKsL6qj6kk8A/Wn3559O5A7XS8TfgnV
83lvmlq6kAbnBWLkpNNUtaqYVPz2Jocka+qE72WIwCKv0mrlKhVsFfI2X8hu
yufXeZauXRcgkmivWE2vWGdKSDH4/Hqb+dhfNMqAQjLjujo9hyedyOdqhnaz
HNoktUN2aIPAWndlrtISaqVzW2XLflJZDHmXF4Ajj7t4ud4kiu9rX0fwW99J
oaGkHI65nmksN84rpQu7t+fUTljoD+8QjNOq8mifM8tEBQbIz8csA4CiVyMU
BSVgge02CZJpt12ev7A0IcDMB0TOOwGkABZ0ccoeblSXqJaRLejhAEWbi/3I
HWguXCstFHGVtwjcGcEUZOqLYj59F9bPWDJgQimbZZgRpe1n8h0FNpfYOn95
KRkGvKJFEVxJaQFf7fYPcGMaNjs9CEQom0pF+XJ2k2Yv9qHVFuK0T3H9ilz0
N/d9BVuf8kEGvh4wlJWOnAHdrs5b9FKABs72liUcS10E5/1rVzBeI5MmBiu6
Lr/f8wNuxJX2dXmoW9z5zsh5HrRJYQqA2W9LXQx1PS+cUG0w25uxv45fvk5O
IoR1WhqC0qpSSTGewTUj0vI0rxJihbXvaV9Jk1sP55Up7K96daXOKXAm+HwM
erDufHentjYhq5p7Cl1hPZEN5EmCmzBjfUeXSQ4d4maclCQKZZxxoF2a7+r2
hm0I/5HeZQb3rWRJo/v08SoHha2KzcpDNjbnTYSWfRnq3IZEAUuHgnlmT33P
MjYsNa37PcV3Ztgzxz0uVko5vuI5lis5lPjeFSCGc7m4+oVHeZ9Tg9Us0asz
LBFrWpiJDwiBChxZX61p119Xk7Q8xsxJST1WgeFNPjqFUo/ivtJSq7KveY2f
0soUT8lNE8xdhDrqhhtfYfE77suQYrLpxgKMBbBu6pQV50tvHifv/elBKmd5
0FS/d1l+9gETVjYAE1NEfi04xqBcDAv1yQNkYJfkStx+H87l2qjek18Grt9Y
tIaYVra1ozOMYwoFl6PZ+jF5qrvlZJwvTusngjMtYmZpjGWKr6EHigqg4ONf
TAatukK5ta9jVse1xtbcDeJia3MVWCDnirKYsOq1wODFjIqXvy93H71IfmIr
Q/7sJLZZUQhTotHMcU9GKttPQ6k8CW7vATWfHk2tyjGOhPmGaXwn8EirvbXo
g/xdo6bDhV1DfxSGpF8DrPy0R1PYZ+Px3t8F4U7KutF2UPr2QZmwNuPcHgxY
Rw1SwVyH1+tk74jZ1iLZ4BLmgap6Sca4PTCSEKweMM3hQtpkZtZGo0OzD/QZ
cw4z5WmZ18pHhSL8Tw2QEgAHWnuQPzVv/ggmelIaEw7DLbW9RU/qOjyebNNl
rGpantRa/f5DQpwLM/4AuZdlaqTkv5ptYJFd3B+j623hndUNM28SSUC4JcWG
0bk/AUvxe/gjYjHhjc2E9q7drZlMjewRLMeO8T5YyqTmOmTL4CILw/RndjDa
0kRHzRHZo9EAm+JL7PHZ3pgmykmW4P/D2ubTxsQzlfCwYbaEEVZE1tqrX7zF
ZFs9XqdaFFRTgPrt5RpT+5+BFH1QDC1QvlaRZBwXRAYzT91xGAUPrf62a/bg
zfjK2iaNfFMXiPRt4I1Ov2qid/+z5ASS+iwwPPqk10vND8+hG2gZF4i5z3Wu
VH7/vX7O88r6wb10mmn/Dh25hD411AJOBZEMQcnTDeFQ0NyB+nHMrRvctI1W
63vhDC8H1LhXld9yAIj+WoTy9x+Xv2VCJ+ChFYBNJjcgVXU18aLOQod4JqyD
wd+f3YR6ZGaft1Y2nIL57tFBKBX1VUmwLtrw2EvCC7Nkhbk/Agexwz7/wwUc
NyLYOQvRdgUJlvGuTe0cf+6MZ76qWcsmlz9bXOZ9hQZ5nv9GiH6D3E29vJct
9Y/NiJxXNpgtzQPiaWaadYaCL8n65Yt1xdYkXHJxmKSQPCUiR+/v5zDeV1Uf
1a/C27Ff18dSUXbDOHtZGU9Q6WoT4Pea9LgrM2pw4lA/EloaDaHLWe/S3bRQ
hNuaWPZVNhbXE8PnNRbjsf5Ov016r2oqT1sM52P3XLB7JA7X1YUpvKAbCECQ
YCDHD7Gdhg98vXJtIAmENYQ/TYcbKGB4D9TvqJn/Zmlz6exhk1ql4jolOYB1
s9Q78812D6j1VriRi41y6XrLYTVfSoiiq+RYx8EUZgn8U5B/uD+xHfJCTqLs
vEFb3cJF39nwRGPxzrIGSBv+uefqUGfib+uWAeNQX0XqdyTrhC+0aYcfA//K
tbGPV02lMpKtTc4hyiQSNEPqAE7Fqj9jc5IM6knkQBUo3h9IIGUd/AUHl2Xj
pd6iXTuKChVPY3Ac33ubiYxxVLquA6cQ3W2smEIhRnTQizRlP9sM87j4CPXj
fY9EP1L6nFVoaYHKg53BXEc0X8RtX1XOO7h6BJULVM9VzzgC9/3320l+a4Ke
5ckZaqIUmbONkTCVW76VItACTeL53FKRJjcG8KTAqpYKStjGf9q8n7EPNfuV
wsmrNVDcP85aEAJc0SCNv4ngSVs1iyXr9B+I0cfjIxQAmkykuyRkhzAzQ8v+
ZhnQhoqKV/tnHXOY2OP593edgGx9sidzSXDeEqNiCu9hH92XFgG+8Kv+NvlX
bVPNJQHXpuwhvGlVe8YOvOLC8Li4q+xalwmSeSwmu5Q6jlcNXL1Ss98fRILX
Nsrp4HYZEbrNTV9GB9VQdylM6ZRrqIRp+cgVrYocXsOfIRNuguz77bydOk/s
QpCqBYNOqqtbPgS0UqWIeO7PQcKdX3z4Ln4t1JlG7oUIbb9Tza7ej2VJVGtd
eZ0XamDUI73xa6f70AWis5h08tuEcQfNQg/AYy/7cCLR0jtHvbtrB2fTaWT9
f5+ahMFEBcg+cr3GYHaTm8vsIHUop3k4ldupemN4WG4cQ0OO9z/eKV7naAow
7UyprzT0Ains0L9naab1iAmC8SxKxpKezRt9v5xAwOhTjBbE50VaOmnQdjRA
wfVnDsokJc5YQOTa2S267K9slF60BCVTFhjEa62UQ5UlyCowHsmDFoHAwA9K
GPBy4TygkFWiXC72ZQ1f2gpiCUZVmYfTXplz/CWFb4Y8OSEvXmCW4thxRKBD
FDc9kkwRc4jbrX/G1DyXCJe7CTGvJQd8zU4rIY1rDr6YvcvMdV28M2cgQL47
+G4ROovvXaGAFrOV/0AYpFvDm1lkp0pxRPgYldST2vP92Z/k4vy5alnDPfnz
aixjOxf/Q832I6XSSMsbyBYbiwgQNh4ToBgY3kFkozosYuSXRa3uxCSx06K4
Nj3aCtJSeuP5FtwaFylSL6ws3RlHi9QBkYXSIhH3nlDchT01K49fkSV27LfY
ljx7Njoiu86IHKbHZJ43RbEJ+FsTZPry4h1S6yvkTC7RIfqOlilt9N0OC1R8
yueIvKNs0RvKPp95nMztueWkvSlQcdFQwpueo99mAtJzEy6OhgpDsGD1XmJC
hf3g3QHKDbhGa1CV6VqwjryxQ31TSx2DGRQeHl9x8UcwPQPdevJaoCareUQ3
DTZeBVCKCuTcwvbPbv6RK2UYaqAKSsOHls4bocIrxLqRd++kgKtPfDJjYBGw
idpCCPxjQvGCvKuFbcBoyPTKxeOh3T4GFix/VG3CT/Cm6ta7f3Fa9pJQmP66
Mytoe1lwO8nZ8sxuvpsHse8iITA2ow9SINUkIc028stfU/BLta4WhpleOAyP
YKSvyGpfPeTI+cfMick44CFsWq5W6GGgWfx8/LVTgeQ8cZb8buwdWLX13jYC
zTU/04oBEoq/MD6MW7sF8h2uVwLZWf1w9kQFvUq0qN30PWsmVRusTKAVpwib
Ew4cKCnnnlpkqIAsoq0TBPIhcWe40d8rBhmSRGazZ71+V3mXKTF/14L4O+Zd
PbNXoOYWdMOehFH5Lc3BARNb3E2M+hMUvS0QkUeIjV0TJYWbzooyRa6g2vS6
0+Y92fZVeyAwAj/ScxIMjSN9GqD6hhLtITo3J9rr4AHAQ8SytVIkdwECsdoh
/w/aYmqZgyDNRNsrCkrBU1y7YNLEsfu1QWGBOesopcg3fjUH7IuJr9ot0A8t
vgkcqJ6IvfyB4biyJCwjM+orfGjcHrLkGgk5Zh1KFnRC3Qb1eaOS9eGe/X/r
QSC8wazN+xR9ONPlRJJiGx87h8fcgOcaNaUY4vzoiFoTZ0SL5C6W+SZXWPSn
cbhBBpc3itbcDnH9QM360gQupSypRkcKCYkyu7kcic26PFl6jZI1xYyF9Mc2
X+RCKiGBpx1ZIGJ49CJtBFkRhBI4uti+X7p+TA5DhH9dpnr9K9b6ToeU75+z
XNBZ1OeWlFe3BkNheEb/snWXQ1j+oksxAqqru0cPLkP2Y5aM+jrfMRg1Vcv/
aWkMy1PCQrMdGoHQ/w/R5I5W3iiThXvLcQvvx1bnnnXnlRrRgqbMEMXs9FMj
+iIqWEjSnAe4/iPryltKU9iblj1vq/AEliaMz0UGlzxpvQoVJx+Etyqqo35i
Tez4kXDnMQ5IVGcFTNKI4JjyRKZx+bAkEeCw4S1aDdaWzrK0OpU3jObu0ZK8
R/Wav1XR5OcVYPlh+dG3FtTPC61rGI8nhrlXsC+TkVrfXFyx7Ftlje6rvo04
r3xOWeYoDedpZ7r3wxg0JrxJTkizct1uAVawowg/dURP8JotMZf+ctfk2thQ
RACUliBTrc/nM1BFmn+OSsp5ObvlgkyVkgWl9nC60jbrjhKftOCU5ZvbRhjB
sIBop6S6/6i/bUxpOIZD5eQBTyIZSA2KA060KbqY+DRzQ9c0fcYbdOxhjgj2
Zw5w98P7bV1YnE5pL/6fVhaqI031snYab3q/ymwmook+CXEH65jd2HLh2MQW
JI1kSUcM7nUErjnVnqjXea2w/E4/GNj/sLsV6Q20liOltbBZXNJoe/61PxsP
+Qvk1L9zL5KyhwCSizyJqxi1kyS0+QCMkKdP1eweJRf+6/mse/40bLlm5HNv
y0UQUVpt2vBK3oswbMh9vHOkealdjJ8ygK2oMviNchKdxakPchz4jSe85gwH
zxfFKBouNCKCgzWKabkwBXmv17ufH/4U7iMM2oAVAn0+ijI7THXFTBy5Tou1
icB8DsffHGlqSwavxSroniNV26pwUwpq8UbD6OI6KOwWrf9dSVHeZ53LtFnq
x9eyh25Jj3s0fIERZ1+Tw+5gmOyIDY5Qgqn/eYVbyP8gKrj437BBlOQQpLKM
jmkyBQm1XkkfenHSIsNNsGpBCb+ezNU8NZWZjvTosU/2/YkZ092P5HDxkqjO
60Nr02SOmeGDIdw/Xh3VhTcFdgzuXnps0TzeFWgx/d5GnvXe/QxpF4PZtNpC
gflkhIPbbbC7pWamg/bC3AKllgPpLB3fY7LtwLs7MW300GpM/8ewun9wXFCO
Z4AQPn0sB/8BOCpLAzqbeWK2z1KXyXQcDc/sg6J5RVTAdkxK6IhDMEjf+L1D
dWdYsV2GUa0VIAZAMz4A3YQo0iSM52Eda/3NouUgRMmtycB90TY3zn9UB/SE
I4TXNNuo/vZcn7TZjha+/1s8HLVtsAu4JBXr7eZ3R03/ocFWs7K32iZsxhLY
LKdwnBYHGwwBozvxkudOBWOH5VER1MXl1n2faq5Zx5Y7C17FDzNDC4CVQ7IU
nkZmFeFX2iRfKH17/v3G3JYFnJgAi02SaeJDfjYYVnrLG+sBhc/zgayZs474
r69ObXV7/w2ekYgisF3XxabLoS8dNCyxDzJz3XJaHv18vHkzSrPNxW7tSfuf
mUtbaBJztwth6K+2OwwzyRrEUm/s2xzy4jZSohlK+eiVbnPPVcxlMwfdH728
SQsdF26tT2GBT6y65wtwDJyVSvY0tf+4mDaJxmXQTZqQEa+Kfekh51sVq7cQ
8+k8x+1Ij17IHLUYIqer7zZixGYxdWQ1AmI4wNWOI8hZEYzJ80sE48TKtSGQ
4yu7ZbY7ygJRZ07/d8f0/F0B7qwN10G2MU/QWrfigJSsTTjIbdX8BKAyDttD
GJRm5WXxF+wTjt3wmC3wZ9kh4m0K3tuvALtdbElveyLDWcwOoMny8RbcUXmf
e9lDTyaUNzGH0yQIPTwyrB+5tNX7AdgUNdCtGR8LhxWLfYaTM6BwBjSk0bgr
WdXHT9hTK4xgXtwPbLpdtLOzgSm+2N6OZt3fSbw+RE1Ok9BXgMYSQ8mBpZWf
JRqcir6rmXDUW/6F91ert5Abx1V1ohFZbptVGm7llAweJlU59AiWKCJ3iGgV
b1z/rP2+dxBfEwOKKbHTSSykgW912ymR4b8rAdCTFtA/dqJNdiQrrqTmiM2S
EKj1Ft80KlaLYnHN8S2N/3mLeSKKj9KyL2G0ZUcNEYmEeR8r2AG9wCvbq+D6
foPy1wlYoJcSj06g3ZlR/JjyyaTGXnKlnsNUZvftAYZ44Fliq9LiIyxSmcqx
G6wu5QJbWqEusl0VjPXDtDvX75CFpkvugea8qllZflfCJTFMk0nX3YGZhfS2
zsyW5pxidXYCfPv427BMDP2/cdTXNN0D4D8fK19Z8jhlUiHUGyWmY3RLMGl3
xMTMjgo4osJ9V2WYpg+BGIfv3pN4bTS8y58aH6axYlL3YMYYbgznoaALibzT
dy82fqd6pNeRpkigKqch5RzaDzTirrXCuhTf3BaFdsxH4gXQJYKEjq9yjxEu
Cgt0iSFAo18iStEuPhOSudT1TpfL8vLJ2R14tTTy+LfwPWS+UXcn2izI8dRp
erxadnFqUi3AqeUzEZFUpqzXIWAdjZwdH325z+WJfjlsGpQ1btuaQi4MXfdW
PMTQfsCuwMXdyyLH2WE92rE5O0gIPIdFJSy8YGhQO2oIvvFwt0FPtilje5Rw
JG/ClQn159UiUYAdQJvH7E7kat9RrgZJdrwfRz0nAuX495WFML+ASQ6yvSBo
YRd6pcn6gNVDXwMEwi9u/O6grRkefgx79TVEIUMOTbbAGTSRlsMywGceXw5L
F5BPHP0ptfUCjpG63qOWOc5sO43ZykqbfgJV3n0IXSXcaYwSkeeqSnSNRzPI
WLeQz6Ol+v89EpqhDQaS+S5EHWfuBdhhBC8ZB0nBeN2olAWfWe+si8ouhvHU
YEmndbHWRh82glv1PAqAMwlwiz1fTVzQASQtW7I9f7xChSP7JHQT8pDxpXWz
ivvbyA1TZdGwuOmg8fj/9QEvdmVofXplG3Iikf7rtNnRBqxM3P4KWYXdv+PS
rYQbtIHGdwYLbQgH+bYzr2GvkZi1uS6GDh0AE8oxQdPJviiKmqXpGaZpB1N4
hi8bZ85XECk9wpylwWlQDt4q8eQjyf6258/mNOlRhWB21jGpqTixnpP6aeQh
vkSnsWpnMFH7G+E7v0jq42ezzZjAV8jRf21ja32Ls2AWHwXgPLnC3YgT1lp8
yeHDYk/IFR9e1xbHQSZHGJGeDca4h0W1mAGb0vOMaGVot2Z4+ZRaKQxOBIGs
b86Xe6QGVHsiOkopnbl5VZ0yGT1xOdjnccC1YjpSoXTf8gc1fLlc2+lDgEU4
4AbZo0aYujINZXNKEhdskOeNTiYNui82nHIXNWvfDQfEpHi4bO/psi80LHbx
pb6KyC4HCePi+sq9Jqhihixg9I9wHArY3pN+XL2U12GPvBxq8bd06AfSeRFl
HDVu7b/hcMu+RbDOPpo5LCI4kqIKaTwW53qF5vAVNbl2OywQInKp/Blw4r/m
7/va7xFrVbyVy/pzuTRGgo0XZGS9jxNayuogtTdyqEjhH5woA22bH/0JNJHw
vpUABc/Vj/e1ul8WT2/DXwwL2TWzljg1EdQr4wu0m4hQX+w4xxhKW+wm76iQ
FZ+JCQO7C6nZzOF91s1gBt+9k+dYRCZ0NRiOqIfbA87uy7rzAKj0F1GaSFyl
PIZuhJ3//YDFwFlN+yxpg5pgAPBMNMXQpgaJhDwMuUFOasg4Ygx81NnZ2mNg
bU8iEEcpw0kVrrCozmZgnarGqMrwMEnbsNzI+uslHazv9gCEtPVyKYij6cZr
fnkjhrBT94yX4BDdw150xUG6XsRXhJCEqwzCbv+IDYPbEuwOj+K8Ib28jAWr
jHsR4bXAsJmiu19Ik3OFY8NI3AfMTAYGA5jYl5F3M5jAWnBYIELjcSdeJdvi
/rpD1PJJmajfLgSQxqjdc0hfwUwiC98h6Z5Xt4bTHBglMASYleEvBrX7b86G
rrtE4/QaBSD0SkNGQLO6fc+S9AD5xp2p0IZl0Fyr6zAFUdAh8IcJpBJHsdYD
hct5FnOH7uYekR8mdRjCKH41St6ZfFhDJLc9NjdTQGu2u6p67O6h4G3aacPb
2bOeXXpq3HCgjOPihd1KhZJfAfpVfS4BIMoYTluiQAoY3KyE/Q9xFputCcm8
ET864CueYX0t0Ykqu2pBPzYMtFqicHi14ZB5tD5PLpJZgEQcG3ZRkHwZ4D+P
XHHHQ1xDIBjLdJGcYsNY4iNso+Qek/g3yH8QRAIl/tHegXlzXu07QBg1hCb5
2PwPCWZp2RPkeXrePOfjijNNQuG1TMRNgBYNao/hQChuWhtT6nHvMhYKsUiw
6jEGUrkkF4SJIWYqxO418kgOiLzVPevbGRn/Te9WmyRYkWoOcgNUVPvh0YUJ
BYwvZPxI8uxr1k9CkpplljtjhNYgnmTDvf5WgnLKbFPUCAkA9cA7IbsjLMeG
JePo46YZCPi2l9Xhanvr1aVOZK2c4Q/65zPKDjXKZbARnuUNAYgF4RTuJkvD
tdG/v+eYO9oDCjCt87BPyn/cs+hKIO0xTksPRfRNm2+P4iFlCte9uotfS3wP
nYwjnIrIlxGFpEnE+B4B/Lb+DV1w9crZ/7/GHpyemi17yDcab3d9L9T3fdii
fDYlPZTZ5S/g63l2x4MNAvrDIH+M7xrZFVS+mrfgG+GoXglAz1ZfHPVR3TdW
vfiSCOi8ClR6zchRj0c9eyMHRIhxz+cbxQ9d5GdEuNDs4/l1h2k+XoJL/d5R
HExfFuLKMkh2PFrztWHPtebfidEd9nsKEhVgLSBnNPSuegaouvmm+QT5zEJp
9VFs53HrD8CzqH8jwfv6WdPhUZjCB25p3oOBr+cbbTUEAs3EsLeH8a3iyPWD
ZwhQXqFc25u6Rqn/zNyS4J+OFfKE9g4vGMWrj4lJrxpaZQE0AwUAu0BU6atv
zVuBfFdeIzH3jQb4w8aLePxaQovk/NhyBGuUK6RLWLpv+ZOhYbqnjGFwMczz
hylgXyoiNfju37/PKKPffBdykbkoHEa3FkcrqH2pM0Ao0mNqhgrj/6OaDoy7
vznPd8QbeXPLcAYJSLHD6+l7OnB6T+7q4zHJXfIIpDb9H5p30uYPXMKogRQM
KxhrHDB9eIdji+urUciD1MATOzmOVnY5Bgl+EGGZFihPseKFJOSdiI4Jt6Tc
mKLUXicIbUhCt0yoLF6U0oX3Unt+VjY0erIPKZ3XTqLCJ8YwDi/kmqrKLNvj
OJ1UBHGus2nqyCfsdrHso55FzsGEbVmDJ1OejqJWyS196In+tHVCUO//7Pjz
fkcce5YXyzQUH/2mWo4yvbbb3ODa26TchykFpnkWd15qn2TZaEMuojNFGOBh
IxJgez7lmS34VwTj45KxJ69fU+X8BJQhluC0D4xZHKA4737hB4p7b5W9u7rh
uJ/AT1U9orORG8iJg7JVOqYaZ4pOLOJ5yOKVYJV0qMWygHhg2JXETZD3JsxB
6H0fXDzOEXmW7hdiGT92I/ZUGzB+jFspHiIPURFIHH4OZtpQN9wmnsL8VqWC
H4dBjJ93sXkuu6h09F/fwVLA3kkFJD1tOHKyz93nDSdBFV0WPwuhhr5tllVo
VA5qb69P8JhM3hQZpBe0b2wz1xO64bTA13zo3fsddH7FpHKcnofVIMM8Nylu
wXfFYyQSnDPLpHfDU7L0025+VBeopkDQlXZKN4gvMvr8Jh+wQGASYxmheFS+
nc41GiKeo4Ka7WzDAa38I32tOmD4wbysfLHmbsgjFaP/u4s//60ugonhAYQv
fMeB26T8rLkP/tMpwv/fCJkI3KiLEezXL3SWWLPJXGneM8MZinSalMH3MGCZ
YIZTKT97dZurXmiPVEN6K7vUZqf42+fHvVnxi2DcTNSYYjWAIWqSFdpDl//R
FYx8bwbwZEx7uF8p98vd6Kejnr3JwmdypfhXZju9z5IQQt2+rKPJxVnpSar9
UhR7vr9r7FLITZyC0qr+YIzRsBnbmLwwO9aeAXx+99ICH1Fioqs4IFbihanE
mO30CLnETkmZI8ip1QAL669ZRPC5vtDBuHVdcWZLzUmNfGQB9yRzciP6pnFE
Gtnpwef6GBtbGQPzjTScd/Hz2n16vwY3fspBYl3gytg3BV0I/QqleqwxTmFh
3Vw2l/S6xQ2dKw35QK7NLrOWfsrPjUNhLD6rVNThv1oEEH6I5+nScGf6esEF
l/6Sl3sMPa+sY2OdcGyjNgOuBOtBYqcEJLJvbHr+1tL/HbCM0fXquFrPUe66
9YaRkwijFpZMFBCq0C0LneS/Ahb/78aATj8t15LMeRSeRcdNbmQsGKnBwMzf
7Rje+AxZJud8hkcZsJeG6KbAeJPmhC8ogy0ojYLF7dBEAGKH0cBgYyfyqpNy
KMiZ+bUASw43d7Z6iTU9H14VQeC8eIQ4F184FwpBAP4/OKr5Tx5WX53/D0gG
n3xS/0nNztgDvihljLqXI7j9GfQaDMMAzuiGMuD3+KQIwBQkXShaCW3m/dcX
LOqidBCdeMVClLw4s9kRRKXi8hWeH1ixL/H0BK5zoCbcLKtmXV4VwUZGlwkx
KbPugoSHYsc0OOTz1FsWFPAsVo/0ipFp06K0t1Abv+UAwm1LUUNORKZIzFcQ
ALdsRg4TLtPkT4K/mrM7Ykjr0RvBU3LfkSDUivfXAVDIXFdlSDQe+lClkVty
raino9YP3Kse/dnPOX0gUZGAHavt7E2AE44bofjN1Jjy0Hq5Q9q8PC+hdidv
r+GeJ3Ai2v3TjgnwXA0MGXGurYvcp6UWknktllSXdSEkYfmnP9bm/Alj+0OP
u5pF83G1s8QgV0dTTWlBVYVJ5iGIvGAjLbcw/ufL2ail0Zu7raAgyRbW/Qyu
+TAB08NjSMLJd3bKyjYhY5Awku53FtWlfgJXudhFy76pdSLLQigciEj4lDpj
2KH5uPMpmABwJ1F0sXNCU0RRlrWrnU8/AyeVuLBP/0LNPmqTANg500xI7kks
ppVlsVo8gU2Y3fD1jvmT64n5LDEMSdymPEy01NubR6C6fRIoGSaLwSjrsZON
qVX/mH/9orLBJp7f2aeYa4uE/LAzVtFST7mDAE8ViAhvFE8RNkXF53nL4kAo
ET/W8fKr320tzCOh5tqs+l/Kzm5+GhCthNUtphUzroPH3DgeUS9IkfnQQFD0
9XffTTJ7uIOPorAVTL0gFKhpx1O5ppqzVEXk7Pv8TmlXMImAlRoJQUHiP0wl
Qg2fp0KNqcIBF4tatCa4qLgRiYAr2Nau88V+nr7TqpbuG+BQiWj7eUAM5EYJ
RQEU2oZZH1GX+EFCjEOqhyoDX+7Lk25mXTRHRE4RrIyYVAHeYdyy/S2h7uek
HZh88+MR2UMIvvNiQwPlnv8XEHapeystw8gVorcMiV6CxXh6ew4LyC8KTdcg
D2dzYfCxQzzlOKLwErUUR057Nf2Ylh4jJWttTErcpFlLW370QxlMf4m+Ijds
CrJShdGAMKDPpEHbTQ0jCQvUTM5wzblUyEGzbV5DUQKSPG1+/wkWmzYeRAaQ
1q5P89GbzrRKo+Nz8/ctQJobkkaZDB8jhAfKyy6xulTDNJYa2/ALMhrSSlPl
z/vUzZf0pbq3VeZxi31q2CsIHPgi+rgtcCvhWX/L4ofaw4/I+XiQRyOoCiMk
FfE3VFqW5X4YsIb030wt33s3MejxIuXpCxWxoZCjd8pk9RLP08JSSVSSve4n
xjj2RidWEUQhK9hjaFhDdLpIDevUgi938kendYJjTCswM78EynExag8kYmXr
D/0awQ1WTC7+Q1GPuma9GV+bJPx/CUuNVukfDHUZKHgzEBfdSPHBAelnQfdG
JPuAVGyJjAdlYMSNp0KMZvK6RT4HjzMZIl0IMfvC1f3sNmvZf8FxeHKPwBst
SWcr4IcoBfTpFThQcoQCU5geSJxehMNMIOJtYt2WvQGjdsOKuRIKYGyKbljx
nWrgq36EbHnEsqTpDYNAs4LJgJ6yS8WRqciDmE6awuHtKVGmKqyDWctXwg6n
4WqP7GJz6rdPZg45Enp07/+7kLHOYM7I+r1EU7o4yUwxzddOwnRfv9O4tqwT
kWvAzjtbSSBRpb60WcXv79aW+jEdWi+/GTsZFyPXsN+cQqKc/ckylwLH4dVE
UCTiFz+XrwMfFaOy4xhI/FGvAaE5fSlFZTjPETiNNVWljnKlwX/2Ap6CvRBd
GDfhY83WpQCm7Nkd7ddjLNJVgbtqqa2meVm9i8WQFZBPds07haVrPUalz1Zp
dOw0Cn+w6reEVZi69u6GYyHeP1MJ7nxAnZmPdHmBcF6M8hi0Mh/IJdVck31X
PO0lc44Jdyfr4TnCmP4X+JMyRCe2WmVZKj+rG2KbpMOb97vsUv1VWrmktnxi
WCLasj6Vf7L+pme/MA3SrGXSyKWmGz9zNxozQ7/Jc3+tmW1eL0qT4ZHkztUZ
iL0mIxsIA6Uhh3/6EdLNuVc94YIsH9wCCGaXfyRMVJmXx9spZoJ1FljMvKdl
MsLS4Ckuz4fOubSl09UjLWtX7pMXTlbXilupGc5+yZTbcH1EmWn2048nZPsA
cbUxNdRw4qygZYY7kX3xCCQxYeLUD7GPsK/r/8bXWhUyxB6l6FNfg88iYBmj
ZUveY/JWE9cV3fPCqb5MV7aO5ghCZf9d60+1W8bNEM7uuHl6MDG1SNnKst4f
J31XDiyE8HDSkt7d46pfuh1i3I7oVz8LaRgZ9lRffyAeQcwRo4lyFq+Ph53C
VnOd9OrAico77G50Ms+RxsE2crxxdiJ6tUf6VvgATavUPZYiZgMSif/b+8ar
ebXIhYM+Luc+bkbXbk9J9+uhJbDCk5faLF3thkM3BUYu0b59RRlt6K9MyfoJ
oEruox05p81tYP+89H109Pcflfn2Kzm8p078Mrf29FO1j1vdZI6EQ1ampRxx
ZGn8mSOrAi4jfThZ5olmto7fWvega92gSTY+6QemroxF7yVBS3nnKhpgAyd4
hir3f9vs00xUe8a74qeTARWUHdC0gjTVOD7x+aQJfX/6Zr/b8PNGvGVhcpWM
umtisb/ryhL7ZRtmO4M+q9mUlTAdTCwfHgIYSrep4eV4SVoP9oXz2V2yfRa4
xax3BiGlOS3HoH0bxYoMfzRUFNn/S1iWS55d0NGsCMIl34Kx+SnBC7cvNaFb
jkJ9ergaRRAt1UTaPYIFMqgOfUvUzkZPz6nrAyDX0kUrwUc/y2b2m+iy5iAj
/WgsQ2kdgUjLp8bPdeusnzFMbcbMxKk4JPwHXdn6Gn5nXgiOLerI5W391oc4
+CpV/2yiNPy/oKds2GptsW8M3tIBTmbykoNKiS7oiSbquix8r2x5RL8JU5ec
w+DRsdf3kUcfVP5rGklpS4wrrck4uDWK5nS5rdl+zcHAg7+okIvpkbAdNSS2
9/9D2Qn80GtUnY222AV47hzG/bE9fSxjcw3G/ajRZlkrEF6wWn2/VMXGvUFW
dn7A6QULafjKOzBmMCtr/cgBqHEYeG7ocxk3kRg+lAxI2svMkKGtf2Xkng7t
trD8mc42o4C+jFuU0Mm3Q4SSpPsxhI1DecnT3IoYYkt/b/CiqBDdOepTHvyN
aMzU1DJSRyhKpSqBWpK1U2fD5+Js+3ibYiBkU7OFiqIjlwzFjuAC5xNqrERA
B55UoqRw0h5KBHg1KHZS52Ij5xmPkn86mmiQwQkKkBJPKg1DAIo54By/BkLI
S56dTUkKMyG3FVz/ZwE3aSH5AT5Udb88JvZYPPsd8c3Y3TVpKzxOSQEiLqIR
oCwH2Eq1hbv5H6GycDeiJO0OwFk2fH+M7FSfE+3K5Wx0uPvOGa2p5ii2QUYT
Rs/a+y0sE6RzyPc+ohr/d20Tr2tLhREOGcZv5BS1eAmYVwh8JknWE6QufHkl
2qHGG/GiaA0fzkv5UTmhcPYZGvKHHbd/pZ/HsN8GTX6CocOhFFXwD6tQhQpy
W2BZ4zKOqia7iy0Ger96m2M6C2UAYadu0oYFZ4Zv8V46yGI27WX1o9Kw/k+t
1kPEuZAi8P5dEhxWGCvAo0SArF/NJZIZHgz+aNNiDhb4zpT96pIxS7Emfrjz
hXmqPb1yGB24J0nL50Yse2EK6xNPMAKLkSbuaDASNZHFeYFVGTsoS1S9qFnO
JBZWN57kMdXXBgnHns2jEsMeUWw8MzeBlPzTI58q1ahhHuaSiohPETcDCCXK
NvzbF3BNNXezSBrd8+YAqv6mSMTw1YGhPiaEqp1Sb/uV7dIB2XXmXpGZ7AkZ
VM3XEMbR2ozvokb7uUvBScMep+gUENr9jaNxaHUnPn8+66l7vR8yWwtZIpJ8
ln9Viejt2qgb4/GJKiatBcp0px6qLiQSUqg91Pv3iGRGQRtZ2De2CmnZKubO
8BjCF3nFnrRWZARK0hKL5ELDfUHKRriuhyXuzSrvbJc8IfAfitFeCyZ3ZL10
FghX33enowYmAb5GBZuIMM3gkPt6cdd1bpFCujb7p7QEFo7sQikRxA2aBsLy
QnMI7vuybyDzNsrwhi3IucqtvQdzb3adG1fSTdGqMhZ48X4/gpxAZxpOKHOu
Ek2GHiEg1+n7FecyTU9nJA40jbCao379RYZh2tdMF8zZ5FHTidG66pfSeiqW
3U7Cm809g62OkvHCQ9WFXtYK2I5d+cu14OQVcfaxJ+OSUor8+Q9CKJTCDh6/
wJM4ighTC/ua6IVlOgipNWS8jl1GFujSEDI/zQT4P0+avGsEFpR3X8PYse15
tN5tCzqK36t3dPmFsIspyP68Hi43pV4q183nmBZ74Rr8UQ6TKyfGl+yF9alG
3wgbvUCY6920b9AeSUhfU3Qx04HzMYmnKqdXN7MiCiGiEClOIwyEMzG5i32B
odeea14phbgO2/u8L3BTucHNoTvZ6Bq01rPS56Yx7/Wam/9KXiZC46c/fhqx
anolQP6/M0q3GV1sfStqou8ufSOVKtReV8VddSNLv5ujiUc6gY3LGDQpLPFX
ZPvsQCFMw+4xSEMF1NEd9njjwPPRiNQACOmYhocrcq2EVkjN0rbjbh2y4dFl
u0UMpGtMZxYXAgmy8tYuH9KQWABhY+BkJd4l/Kyypk2BBOpPiNlhZFMRxuUK
JjIYxm5mLtS1Hmw8jq76D/Xfmgc0JHkxK035YMb7+LB/MddUuw/43SR75x2/
twWWfx36iuWHcBFjfKAYg0fFBko5lldVHCaDijV/opUpk0B3K+AZ+BBWcWDt
Hr4M80fQ18483HdJ4jGgzotbiw7bWUN4C6KcTQLpi0ROZI1yry0Dvc6wHi6L
+dP+ncSk2xC/yLw6zMlpTBlf7g4KWZkN7IxeZYLOCKbpiCRxxUfbWXO+6x46
szcUl6odhRWlnAsCM5toSl/v8ljC4yGuoywc2qYgzi3Z42Fs9ZKVmnvK60Np
Wmc6VXC1VErLIK0W+hLBloA4y9iERs+Kok+lLEq7TkksJ2qrflJUiKL7dH3W
qxfoWa8pgNQ3yMS0xpybXzwyjfFIXpNPHWL5QIvGq6ZRI+v4rwqiYp2YLi1J
1Pr4000heql5ETkyV3QdwPjHZ/pjgpJwq6ZC/IjRhKgIxfWSEjuSPTsr6fmt
1uda+IKY/jobHipBrgDg0ssYbuMR2QR0mBRHvDOSu/36d8P/1tLQIKael7PM
y/KsrrPzh8LQV5+2+KL5Hw9TVTwNSxoIeJdqDTafi6SQBYJa47z9GYS5bRd2
ykg9v2oHHni03Ni1iCm2BWdUqRUYyA6QfINsUsdPekWZZ7H8ZVsg6oW2bbDN
Lq2kEn+Q9MjWd4tYksJH8webt+Xeu2IMrGqKgijRHV4TsPX7CiFjOFkVGWSs
DOpbCj5BZwGL8VfRpQa6JUoszPjciSk3Sc9brZ17/NtFEP0chJZf+HHKY5vF
NbHkKlvfY7mXPz0aB9f8FQ7dIS6exlpDcU2aI5PHDn7mU5Rb3nyzCXHhwIwH
M1CQJEVD3aUqYQdUcqeOnl+BlZqLOzOlBveKr5bghSeexecprKtbKWlrrYzo
g7KAiSeoWPw7tDxBw6KtvVKqM2ElJvqGv/1PTNrQMNh1TXVGHxcoLQ/O9rZd
QLuAqWNpIr6HwsnS9CM5SmVf7MHNmhoYu7sssrPwSsInmzGuv4EktPfVGC+D
XtwantJPRNlDfUkFLAWD5DlTPq6as5zzPzR42ZscIQewEXV6SHVFKwKmdYcz
F3olEo1NNxGutLdIZghTDItB8DM0jPPpSBNmnKbwnfLbWYFDoOASnu+SbGEa
D5Ig5yJkoJ0G+fKxtodXVeu1fyrYRbmvOtxYgPueFvG3XptKazSVD7jAwMXH
L2oL3YUfYehitEW0+bwT31pQWm4N6asizEnJZCB6TbvNhn+S4V5rmWH47VBI
VM1Qh2EYm+HqejZY/oUkcgMR853B4sqp/T7f5hU0Nw1u2RKtZVNpjfO/D0Zf
hv9zaW7fc5VKDvDag6fEPJ7zUvM+ZIi8uEGLlVX5Tbj1wcWoSuXmpoLoMYLn
oo38zPIIkM92o2zFUunhRSTabql/l6BTuX779ZgWlCUshgIl/SzJbx9xnRai
ae3anpys0x0bPtETlAnXtoW261ZxbJ9sY8B34bbtBOL2aVWxZ/26dFjtrjaY
FYT/hYzGPXG/S8vY+kmPfeqe1t/CCZX6B07bBlWWd+gJLH7+8GYMyZYv7Cai
c9srIPlhNkVWgKLU+8m6SohuF6zGaQniKrZQFPa7LKeNus+QKnjaPgi9qZve
fj6QxQaFGBTHg0QMQtzSo5Kk8Oy87ftG8pWTk7TFY8Y3nuP4DuAhESqwRlAh
mf6CnGJdqa9/DawvBco0pHuOstdUsPwdL/+QCyRWzV7q8NMD1sy/3b4LHRJc
CctckZ2KcOAvH6xocRVC7lamS6TF71SJkx5xyylZOJcDvi4PXfzKVwfkMAmv
v91QJjF84+63afRh7QxysHHWqBns8EhuCyiSaDafS+5FH29CN1inuhXm/RIT
UKF1DWbYLptKCvHVDJKyiC9uq3KsdssI2whKEB9nZ+KQ4dp7DHlYP/VfxMQk
oL//PI5OcTK4ijIls9lIQlNJBEMhs+uesu39XxgTcuSn3sui2zrESoEi+6zU
od5sPxqDxac3oyk4LjzSufLPFxNqP+TSPQUnE6vhjqNis68a9+Vx0p0o/idp
AVgvvozkJzzh4gBKAppr+gM6HmUNY5XUXMSdTOCRC2nMNP69zhGLOmDJNK5f
cWKk56IxTWToRG3M41AnQyg/OAXCQ/cvQSNB/luJY0GKw3ZoLDz6fRDwU0op
i2i7bpety5jni+VillOS11H/8VZoJvAnqnaEuBUo3PSOR9FPtlOLjQMEDTnl
hUtKuWKiu8Q9Bh1pTVnNdiLe5PpVTKSIYKE4+kaFHVnCqyHEaG0cxT2LsWY9
dS6Ynwzous6jXEtI5OxAbkA0Vz51sA5zLLA4m4M7dGca3llmrnirqTwE9wFJ
KRMpAn17+9oe8RRQGBVw2TNqjf3lnX3S8PPpks0DDlNd+FtkEy6kn/jkEacl
kiPgI+eBpLgWBaiVNVQUpl7ZCeHYn6QAkZJ59CihSKqzMhgbeh7JUNyC62Eo
zkUAlemipcxO4TJfSAOt19fvS9LlQUietxJ++50nI//pgN5LcdAn4MQu6+FW
YOCwDx5regt7G4Qv8Vi2UwdV+91ZqJubkyz7VxFx4x3B/689uhYvASkm7YaT
fH2RsPDiNp42SRhqvVqWMjntrDj3CxINZ4I3RMewY0VNtC5oyZSrfYadzDNA
m41bYCFvmtMEh4fknxO5ep9+LwqFVD+ubn9+T2jhRFRgcVDTEX8WM7JClVJE
zF6GKpwlkrXwW4up39U6GyqrCa6DdpSpg41QF98hmyU4Kfnezo6UOghMRUky
UdbsLoE3/8vctNDyfTZ9rolsm6atKIfgEYtQnTZ2OQalCDIHiy6/ncZJg+AO
POzRJd6Wwq6DgMZM0LTFNW9RTSercom/8xeKeL1TqMIftuaORn7Wk3no+Dx7
kmnm

`pragma protect end_protected
