`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
pszipoC5YwFY7RMq166jzq0IL18URt+ZgGNSvtyy/+eDkpwNmk1HWom5BfqDrKwQ
f/PWnEd268Pr8iSQ3UN1mogEbiLQ5PMae02i6Z+Q/vTEe4ev8sq0G3skhbQ8K2GB
Xl3tH6JHoPjxaOp+BKkFAXIzBOAN7aCJOWJuI/HQuEc=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 6000), data_block
vbmZ+NLoRXX5Xj25efO5AQ61frZLFX7WDUJvB26lpTirZzfjXWvbwUtjfvSYLA1q
YQCBNm4S+u90eyZ6yCw2BEOQ8twkt/Us86Jh+GVd2vQ5bC5s/qtHBpS48DMCXWHT
OQ9F87wdpMOX4xoxeDwGKo5ehzr6Sneifibttn+LMiFVKbePWYnKy7hJn6hRYErX
26+3PGPqKaFaeGPXEszpnTbqDpvAtw8jWs5pKgTrYrjPfJgq1GLc+5e6HOeNuHfQ
rDX+4S27l3NREXLJOPU+UX8Dn/QTiCFCqRRm6+EGhtY2bguPkxrNCoTxxbPnAhER
UW+LewcnD8fteiRMxOKUN4c1TVTFswsQZUElbupbMMvivVfVCki6/xJmpuBHz7Rx
avg4maz6OsGlBUMz78aOkpGfS43nmFHahbi+zW3hLumWAUFJPXi6TX0VShgV0dPw
pLh22mDkSVyjpMVzH8rozN6aUXEKmhDRgxddbw6C1j8AZbAz+Il0mrjMNgDkEIe5
vdcXPdKuQwD6jOcs3xVMWchqbbhn6Zqp8E6nXiZt4zcwKC/N+Xv6yUMsUAi5qSKt
aTqKzIRegUHvtM1aZQ+a2YmCboXN0W1fC0E1cmZP1MHdQXzCYfzSDnOmpopA4pw2
/sZtKwkO7vcpfujgrgBc2xdRnlHx8Qk8qWiSH4Ya7Y8TmauRS1kFYLIkq5AIVFUQ
tNzLDwfoa+8rb0bBB2WNZ0XOB71ozl77iHLX+tgrICvbvkq7yoaLu+h3QVY+F+ad
XMx2go7k2upDiWQlmCJc4EWCA6wg7TlnYwpA9XO8dyvW7+4ryrWwpl8U3mtz+T8j
iK15RaTJAVmcuTOoEVvfsjpZurzA4672xMWKbbHSqY2dMdlHRHfGBCoJNivd3wGU
j45vFRYOBbgub8a3WIFV6Ca29wLmJttgol587N652U7uVKGc2P+/VIkmMF0ZLXCx
YuqyGcvJ1d/WM5qNiu923netN0Xu8ME2jgIaxrVxXJnJU1EbeKgor3itfzt6+AJ3
5DowEYEKfsYaWnLi6W7BB9T2DhQ7kYRy6LNUOgEi8CvX2DmG6Z2PtjG4isryhV29
PkU9KfihJAg/9ecRmu9pOhOyvVgGhXyQvB387NzwmoHnoqmsZpbObXKU+/IAMh4y
RwbzpfN+7jE2/7xFRKqMSjjZbB2ZTKB1hqlPPkStfV4Whr/aWmQZ6fm+ZWyalun/
Ml1PuBYkhcAtfYSnHGxUz71ucqF6LB3tUMG7MS2wHJo96rOiQKJD9sqjeBB1h5vW
Kfzv7nef8iYAyhsd9c/BEJyOTbECsLtYP1GEnHiqIBotBGdId8bDNgZY+vkb6x5m
oP52WsTt6FflBP004n2oPYTY4JtHMXuilWc3dpgB/Vc/49pdchABuFjE4GsAXQFZ
RgiPy14qK2hHwVtnNN/vrCQMIQnv8h6zXUMI+B4DgT5qNHeIWFz3IA17/U23TTQ4
2ZYlERGEYhk4n8UIBhfp9peqCD5k1e56WO0DsM6J5LeipUCl/QR3uo5DGulkppZI
K1r2NMH5/hJ46n2SkGOcQ2/WUSJd7PwQYFPNzYc9KqkVRwGdszmJNcAVsnLmWRpH
UH65u76Yv8MVGAA1BDZ72WQKUCVipthoH+SI1wHnGXyu1LmDBVtZfdJx/R/y7Ytr
phmd4A2jXtE1MRypdaKYiHLtJ1FrsWRglCag1M33ykCH4Rq871leVIqyFCmOY1Qg
0BERLlMFVYtoYC/Ui6UaJ6mu9CcTN4UG0UsmhNJWD+bwhyonA7UmgFVxxV8HCjEX
vi3IMk5fVDFYQeNCS9d/ScF0cjpubTb3085N6Dv0wmfmTeoO8pVPez/yKUV90rXH
PBqH5jsbeXKBZ9ZGZs2EoX6kivV1/g6ioHPjU13ElZFjklW0bjaMMg9sy04DMQSD
U3F2T7vOyQa9YIV8DLflWhd+ndLnIG8nM3UkS4zY5qr/lv4DTwLt8BryvJZQoA0I
YjL50Yu7pT3MKcu/zJmxKx4HO435kTpJSolJsi2YgPpOaNnedqqp+qLSU4YoWF2e
7oGgOJ2T3RMzGMv66EbeEVCeFXq/n3D+Yink7+QtlfyN+8010eHZ0PdI4wEDZWQj
oIMv+3oxNJdhtzVukLqB+SehbjnPRsLnTcBL3Z0VybVni/PkpAvakHPHWbkbcDmW
LyRIC+px4Zvt084UcjGrRoWZzjZncKq/hSCBDKnFOQVSWXzOxY+ddid6MIdYIkFd
orWfwttHci9J+IhljCusH0FRcSiGjeXN+I2604DPX/HcER+n+dNR+RJPUkcJDoMu
Aa0ShOqgB0vCvLWNPyxdWwe7OUA00UfTMJeOoOxyLClzguV7uAzWQ8cByqoCADG5
qtnG3a+3yzBE8yMK0jw/nfxwWbVAJ0+yDqxmKHg8+vT1Y7NNw+Yx5ULhkueUYM0N
8VIK2/x4TlEppRVZZkV4+gx2ZgtUC2oVi0wA4S4VSZgSLfz4T2qVJQ6fAC4alOxc
6MBzz8lqOzsRBUFmf5s0HwNRAMnxS+t+x4vx1iBdipNdMCz02k7Ua7dVXv0g2PPX
25u2rMmrsAIcUgZs/2PnHJvOVzxaFxiWWUSiYqTDD3i/KLrUbUlnVJM1/961MXZH
q9IZztArp2/xwsdo0R+YE6CtiSbtD4cjdcLpVbGcavodlbjmeroizC/8hTq5ruwG
eaf5ZMZkX58dgR1R/aBhAWdO8N+iaX5QiUh1isdK8HBBCNdi6FOtG39BW34u2xwf
+8+XBH4Xc5WVE+jNccmJNV+mjtZVMVeEAq1GVOC+28EnW+YJxKbP/pM5KusnZTiQ
QRYteqh1bL1t97ttgaMh76gw2xZoj7R7b+rDVWg/JMx7X/BYwK9nQLHg0lpU1djj
a7UtSHBQvY5YNkOLE1fxIbcE2yOvL3ieejbqj8XdkyWksyCtJdIaJuwyVotydRA1
bOWnyvQQ1FojizXfDdLOVeRjz/RAoRRkuw773lyHRXykH9tkZJrWiTh0VwcH4Xan
IHvvhIqw4kDW7NYdsGGCjlQ9+aH5WULOBgkAFRDgYwapWQCvkx2JzcEL4wo0mwbM
Xej0SXM1bXhsPZRmm4nWVR9bP1rz9G9rBVw1BIIeKFs6ZagNiUcq0Vh4Ssa0odJG
WC0mZyAdFeOc7/YIqdp9g62CvXB5ErqduIck9j3R1KWqnEsmQ2jqh42Ed+zQhEj3
PJnme3ttVltuokQDerKES7XX0H03RPglaPF5mj2CBfGB5CBYaA6kKeitIH4ZPUgK
aaxmcAvKFJ9N+aVqFtj655kkQ3bH59BPq0mbQCUChCZiDbmVlUYP7soypsmmydxG
gO2cv7UtMhKZ3u1xOxZhs3VYoxuz+gHs9cTs2bxnrxgX+1Yjtd5zlInpw5QJN5Qa
ZZvbkMgwgOHZiYDsg0z0e/qvuV0RMbfBIT+11YgKmIYEa95GboYNt1Z35i3pB6UK
toQwc/BXrTgSjmfWEjF5ba9kGZU+vkgFMZoe20Qgi+ndVYa30swMZLqgYPAWOCrm
4MsrLr1KMxHwRNQj/K+84pBBf1wpWKbUQeGJGf+Ke0givzCLQElAGdzu8yV+XZYt
HTucazq2h4Lg9WbjFhQtHKMcMt7cRnPRY8Hg41clhp1KWACByUX/KZk5do9RAwOY
T69p99/CzF9Wio6jsSXz/sZsutGuKQ3XDHANF/byQ635lQJfkJF9FoLsdzG/6wqz
2a9JVa4A1yTtCZho+tl1vQRgt9QCDuF1ZcrVdom9YASdqrcWPnqf+rPA0YS6DbrX
SL5Kjjw7m06z8fQQI/2Dol7afIH0kGtqhgxkL3DOYi1zF3sJaPUFSuvidZlo/xn4
OZ248a9PyrsRKc5+MgnWIEXavX7VarT/B2PHdttN9heTOqBQI2jPkdpWIU2Iav6h
GOpr00dAa7NpMYUee78GQbwQ4rn1HLScudI/Bav276IDyBcWEKh4BU9+6A727dN3
dP9DvBYuXv6bpvS5jHYQNSwnklTwv8pozz5uMAShlORxmvHxLhm7ryPkWlkCCYqW
OMDkiYGmFxPZ9gyTr/Z15VN+gkIQqRgU5LbFAAviUMPOQas1x8pZDYzVFeq27+nU
NaCg+jzrQSmVtmjhEH0CztggL27Rl3nhpCcDLEOi7Hp2j8fA/1ys+LM2LKd5+hAN
2gs1akCZhK75M9IhC0H/Tw0ThuTeofPIzZ3qvh+21cvJhE+Iffk3WiIfxo85E6bh
Iiij9NZGAc0N/TTlSfw/HlZjEFgDziaWJEA7zPwIB0weaLgIkF/AS4Bt6skbt146
W/PtIEgGNVhXFN5JVuvdX5IjQ7+7NsXijJ9l+o7eZ9jel5RXRp6I/+hM2M5CIeVq
M/JZuSJRX8E/1u5xzwgEFkRLEAicUp+dQsI01d139Rym4haGITilMOraRX7YbpVj
b/6BgX7d6NFWHt/PtyZN+sRXupjl1dE7kjFZs6CwAJtv6uU90IIbW3wdOjDBe4wC
5E3TgJwDO++5RwjhVoeqLN/S3B5/VGA1LEx0LeOuwXWeIQewh/p76eXk7fSFfmDw
GuqyF6GbZ20QNac2cWAkzS1aPDJeqMTHGgN3x778FeoYkgoiPXghOuXcef0CNK08
V3CnRk5MIHLXKL1qaQBs9xrTBPwAdjmlAjSO5Dv/fODPfnRrKioJnNRcIWAJyOon
NYiLGyeQVY0Da0R8hgJiOOJverErDlL27W5DzUINl6Wj0vE6Fo8iu/6aN8NWul1+
PBp6e5Yls1PaoyvO/HCxqaIQ4bwui97U85NXSgd9zrqnKxy3aJ5iJaylVQUUGUjO
hLKjY2GkbuY5Dr3NfAZorlLTsWafI4rHdSiLgBJ0FhSP6npgdFj7vEoeTqXbJgKx
ImF5L/4aVniZyHhbIT2ktRxWWvnRzymcIrm4QTKGTWlVbasiZQ/d6f0EBd5VHwBe
zH4QZxt5kirv0Ey39A6pZEj7MEdrKcHHMrHr68IkhO5SN2gcbCk7P+zrbKVv2NiB
JRVtqaojZslOwSDbh9LY1SRiTMkDlDiBCwIZpYT8YgYaikeB/DDPd04XUAlhnXE5
N2uyx8b6BB/2MoLsiCmEp4bOdQ4216V0v7NGUkdlELlRa6kcWpv72Ya8Gj4Zu92W
tmwGWXhUjooGDmXFTmO++A1RO5INXvYNn7efDakm/s8XZdyfdoI6DEgb9LbahrhB
4BBmEyiCot29NCTNan0Lzt2hcAzL5x47Kc/+2hyBGURmBBBAapOQ21IwuIMC5Aj/
eZuwsLl2m2chnrT9+S3iapBsnHCUAdKQ7Q4+FXKoYCifIIJudPakz8LQ5OuP8hTL
Tqoqq0JidC8hzzu8phC+Ic51XG4D86AJqv4Yv4+wBm9C6MSaAqd+gJAoDZy1GwVh
OT4enGXh3zfs2skayXcfXv4v69zjw4Oi4x5lACKhrTzITNhuw+O3L5qbkyo+m5Ws
hZVYfeKeNiDU3yXPmJT0LWWL2fXGyO8FwAWxFCnZuJXGZUlWsuf5UTqQkOSkxZFg
fs0huE9JPS5ifs4Y1uumV7GyLDikDwL0Rk7FAc6fcnZWmwq5kLbEuHdLhOs3/2P4
vV7/ywNWfDlm7XBwnAjLXsBDFfG7k9BRsmtkLmfJbCXEfHHDMfAKmxPn5+DW4GQz
sXoBOvTOzxZe5V25azl1bD3XZEqkLv3y2xTvVa6osNrhG261WOxev4UE+T5Ib4Nu
m8QqMjX+jZukqzaXu5yLfrxqrqWMU2iBwz/sZEp27IhQd6FHRwnVyUy49DqI0SIi
K772b67/RS4Ac+jRh7H+t8VH481J+pG6Lr6n0pL2JsfHHrBjhGbomQ/DzDERkerV
fqaqxt6DZ1OrJZyRC47W5QmDpK7DOue3PiWjgKGeCanpqAgcXTrmvV2U0xJZGOaM
TDDDgZLMEr8jL2m1t61kt2Bc/teQBt3FhDu4EwzDsL5KZszEDbKdfzO/y/+HTLa+
RH0b/QRfQ8AAmu6kFVNzYZXLsw9xi7qQg5OsA34teoipJexB3zi0gSa8Z3CKbp4V
9ZUeVfSbgba09+DEGQf2iQK8/N7xI6+02kbolFonVRAFV4teKF4LOYqU+ya0ajsB
sFX2Xbeq2zlCJY572vLwfkNE7rfOs5ZrgBVXMMZkVrEsNPc9hrv0DZQERDFHsKG0
cPHd2IChjqXcPECCgJu5b8bpXa9AcCj7hrzESJOUzcSENJDZEGmCX435xct+2ERF
bPGyfxXyIHQwyBAhHU/zFPjBLYWzJxbQ1/IcIt4F3OEtjljjYtEWQXJiR/5Nk1Q7
1k5mW0tF58XQCga430oQz0fYfbeSHOc/8NWVgVD3u3Frk2bdzCsDFUVfZgvlf3YF
3RG4MTJnW82mFHa9an0cdvawG6OgXft/NvTRv4+6jg7pVWaedBrg9bPGDL5mPSgy
o5+n2TFYvsS17muyX6ijI1Wd6uTyfeN/G7ygccknw2GeMzzMmTR6ujD263DRE2c0
/K7B06Xr/SxAEJXiXITsHNii9LlevCGFpk8opVIkUyakcAQ/Os+EgoLT5tTpMvhD
Yq/XWxx0zPqB9kdDoTXZl9aAU2Xolr/TBH9x8K9hEctxwLonth2CvIgI5L5fM5tO
1h5Ulzp7Q0bFXGcu25aPFUsHt2vWpwVTjA0VcHgiZLA8gs+dB9qAreB0enw/qINO
UHmwDJDieDg2GhkdzFNZduRKVXRbq3NdvxtHqH73Dp6SC9GnXq6Xn3dWuANr+pRq
POO9VteaEigQYfVu1WARrN0kqaL5sGz1iPXbdfrRhpHiiVfaGucA1SbS5Py4wCDQ
Z1BY2UcJqiB9+zRrTtasw/tuBKRf74zhB6pw0JlOmyKC8LOpu+v/+SavG9wD6iyA
bjEI9YHojJVavcb4Gc7WGiRy3V1kF0CRq6eHltCIVXQQ8fdifY0AIi22cb7opVat
AK/yXyK0f0H+FbvvOB90VhVVzqfMXUtqBGQIxSHMZNLNEzR/JqXr5xuybZayzRDk
fW4ztCf5Hs31HYvzVWkcWfjosO7VXIRAZxPsBKGg7A3ojYf1p9FXEk7LU5s52FZA
RAgujrA+W9vEWuPue1bFO4aUftWBJQj9N6FPMEzFGgenhDP6PwmXmGTLEx8vlXQO
iUXC5crnJ8WekpSHAniqwTs/hxYIMEQ56NgUpwcIV2+2ngd1J8cdzDyhGD05ltJN
nCg4Q2mWOfoBg5DmdnE2L2f0dC9cTF8sMinMf8Dj7PwHzXtMGgssE0/Xtim5yGmq
IIzzPw8J/AsyJLR7n6jvlqN2Vc1RUPBiQTClEGuhuyIZR8diPc+bk1JtOcn6U7BY
0sqZO5FtPK0xLxaXQAqrreOpngLv/2Mldolv3iJ1pGh9Yda1pEyLBmltTbTrXBlQ
3iu6XRiw9fiKh5tGMDpV9qFZn6HuPXw9ff+ZGiVVOIgOekNIUv2/bmniULWeZF+n
rQM/DIhALWAz6JYC29ewVMsRfjEF1dJeVOetnAFUIkQJaqO6R2Z3ngh3pv1x2xPi
9cBWtN0Jjjidg5YtdYUrgx4fMPmPwfa0dHmTQkMz0eh8RgcdiaJjgsXuhdfVarxh
DdEms7hS5Ww7q3fxQ9V+4HW0SSHh13XAOuAsPYKfP6Lv4CDxhmXyiYiNfRQ0IP/s
vsAzXzwcRlE543kbYwfeuv62JSH0P4r6UJH5fzADDpqrSed6xL8zqDeltiUBUNHw
bzdA5rAYVEy+JMT/ZXcnfzB9s2M6/9m6DIFL3YUiaXjaXLQlqadP5TL1W1O4560f
IOYtOMHzArK7K2MoiIM25YumtuuzydNDv3/h64k7TNrkVjRG0z+ee/WJfKs8m8Qm
xY8daQ7bl5VlNSRuausF3jxIuhMTghjOogX2EgUdBXsloUdLqXbDTkuCXMin/4k6
CSNDkmBqq5r0PRngpc5dVOgcIaivp/iEG89Di3YJ2gX05vQ2kACWvAMCoqsL5MOo
+R+UIoiWxcmCGwzaKj+XW+S0wWc3aLBK6M9HLWfuUjUGvmN2nU58igQF68C7qA/a
`pragma protect end_protected
