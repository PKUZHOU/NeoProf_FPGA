// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
FuRcCwb+Cq7e6MaM1zpX+A6bvueIcDPMCAmtkV0u7F+OS0M/LNTnIARBBPXTvdBV
LXCMzS2XkWzpPli/PRF1Ago4bgQTXnjYJnTal0afn4Cwrol7C35lNdB6hHV+VCU0
NTM/LU1q/Typc+O5YCpI1EVnOnBPwDBx2ZmVAMKpzPc=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 10864 )
`pragma protect data_block
5K8ZDSILZzpV+gMPG3TZ8FX9sQ37hjyDtZSmYyqqEldnvD1oRh6FqzsMPLmP7RBx
WlKJbk4NupPBihb3jJgreVxwYtKkHwmVukuNFMk0X4T12iYubtG1rNla5AzvNQ8O
zEuw80GTJjRNEOWFVEB2RnWdo8FOeiaKNYiauorxOWCNlQw6xc1n1GWKQbPAd9/Y
GldnprsX39rXPkvbohN3CSQeIxDMvCBP/Eu3W33LiBOmzyldq7omt4kAbXATd0pN
3JgQ9zbJ0HW+YfrerVTdSJYmoRZbw1R3TyTrD9g4QPT0RuHTDCNNweXRPXaR4GA+
f0TlU+wqMBDdaNYmwBNnrnB52UwdWR2wwgvB6gZhl0cK4gYXKnrGTzcZYhf5o6Og
Rr4bew9iB/X2zukcx+Rr8EtBST0or5FiMjq0za1Pj4uNMnUuL+aejAfGdR0/1kCC
nbNLn2pWYdZ3fhRFmx/vGWLZRoW2hpbe9MkIPKoxqRZHeA/63BYTS8Rm+Ux0lP7X
ZhMc3VyemSAHlIqgCXE3nGUCgceoF7UjfqdSYVjueKe3rPNRAZZf7RQaTasirHlT
jZtLtG0bduzobRD23/yK2ZP/Ie1BhEpAIk24fLJXb5OqHH70zjOaAqK5B9/EVmTS
ZtzINbE2GI52+FE8gpl2Ph5iAsxVb2CETOITjLSxWNlN0mjY3x0JOaUh7NkZ8YCJ
GOgOydmLEmW7ERNJvxAH9T3EzXPR7LWvwRy61AhOfSjcVvLyza1kdYHQbJCRqwfk
RJkSy+kaBxCslM1iA3N/Cis6wWVv5GKs/7r/IipvG0IMYXWLmHMD6kHUy/myAalw
u+0XM+Qnn7CNyW9x7K577TwtQoi3ZBzjbTV+Hadtxxgju/ZH5XhB9q4dXbkiSdGx
BbUfhZdJkGePa3aP4RpLjbqa1MUSyU+Xuj5/PT8WJC6H1FoKFVEQGplphg0+Km5e
ooDNo+iK/kC2NP/RUV4clmqmokQc8A72YaijmXJbMJMAldpMXQ2UsJxufNIaNYF6
mJlWxWOGRCoqkEEtVeS1B4PLVUK1b2JGVAY11AwzgxiWeUJRW5+xSpjl5rkk69yk
x1RXs9MDb0YaqM0Ufwiz7/nrF18Y+TgjG3nFrVl+D56mY3oPgq2k8akLe0IIE4Mw
6wtw2t3mXfD5EB+h1V2OYwdsI0bt3t27WZYWtl1VepoR3xeMX2RRdLIn9oTNc000
PYsYTCaBy/9wZZwZ9q4zLLqAVYphqkLLZA6SfQQi6xiPRW01yuCPErD+sqHXBa1m
b7OJ/QuKaV8OswZii/Th+L3unjxj5uZS40LiePUk15FRvOPro+k3bU75mfNBXZ3a
xrAWuUhrqbeH2MFEvdXvd7dBPeTTqeReapfaOCAlPY6yiYS2PmiAb4imWqko/sEO
eASf0gQlH0gf8qYbZxJ+0niEsHETlIqzP4LylreUf/seSrycRfsUuykZw1m9OPxf
KBazW/F74rq67roQCsKU1NZbCNyo9dWar2lEJfL1+wXTDxbcHYhqQ6vAHbq61X5K
cErt2Qye/r3LR3WJq02DBKodpPoyZLKRTD20CwdjUhVlDTeOn11/7NTEgozxWP+B
CIs44OL/TDb+1AR1RIaFD3Z07AyWNpV0Ey9ltAOn2YXHPgA/HfT1tubBgknoyWjB
dQL3Arw/Yr02cahf/32MLpKg+6ZGHs+10FWhj4QKF5djqK1ind2ay+OW/UEl2HP8
KHv2Fu2EyOKNuF8FbIMGj5/NriUdT9ygPeXDj8qcxJDsLGJ5qla+dPrkOaPh9BR7
jObeXf7y/JIrzneo2T5aDMtOvGoOmOsCGAjqiuRtS3xvIhDfPY/wQcFDy8CaRm5S
FflkZFwyEMQfYPWZVfukiv+em0AWTcat/QGuiu1ngRYH+PkOTLKMY6Gpmwg69sp/
wrbADtiR2X9rQSmPdXAo/MVsVqVoh8L+2AJt/fR/BVjPUsbDejxf45nc+QEgTIW0
Lmn8aWZ8AifDmbEijciGjomm2N3u+qtV5cmpZ+IHo40nUvUcC4Y1UKisOKZppENh
tACk75PxAemzwNQrhUbdLBLEmmt5K09zZwEIBZ5VLpZ84AFOaov6Vm4Jj5d4WS+p
bwKCL/yvO8w5B66twOfAf1mcozO3mxIYPCr2L65RXoAG3LCJbS0peh9/CoaIrYzq
Gn28eHgqYKwGcswp/BLb4JBOzGwUUlG1rANUaTnxD10pP7/NHjU9vQ15QBcSl5aM
qj+4zWCmQpPbYT6lVNlikek0HaIffawL5rqQ/aREDkTwTb7YF7JjLaT9uImGZCcN
7oXkupLjW7h7zwj2WiDYgR6naHwG28+4YUkHnWweBUyn/FriX2r0uo2jqf1nUgJZ
tkbXrJhVSURZjHrWxsPafyUx8a4+QghGrMHe1vNUYN0PGuznpLkbSh+Z6f/RGqcu
Fyyhza2oG9Q9TBwf4ms22r++g1R5iUv1uoI3Q4x84VKJBrxA1ZpJhmG7M+uRcjQS
ySCxsD2/hDZRXZI5YjmxEVF6sSutBLwoARfDej01zM2OHTzwjC3MwPC/iEp+Ax4U
ZpycVw+n4jebnoveaJTJ6YQRbVLWUR4Gr7i36ly/qwMwNE0nMCBFXPTXr97hIZsX
c4LXz7LDhZLhv4widK/Wm792pW+5zIWekuazBEAKFbiAxwEbfmzv4p69THkbZMl9
5uI+MI4PDJra4DN7D+pgI3Oxmmmr9DdE57SYctNoGYScPY/9Pdg+lz4wl0e6jBq8
FZ+C/UrmuH6zWV7fI0nAAK5D/qwN55D3OWCA5PYme8jWKYyI/gFn2w31SJVzrQg2
sFkM47I7GzOPrpWMKsQ5KBV45e1hW//I/DO1LuAIzJT4hrfpjJ6rF6/vAncS3wuK
HxSmipQMon3+qb2ySowXopGRW+Qfk0gqdOYaVxcu++QQ5EvBDjflYa8jHCjXsHrz
BbxM6CkrO8Kr9jNoYEwju56Bqt/8cxTE7mQgTnBTbObOx2rBs74ro1eJQ9dsXqj2
W5o4nh+yMAq7Icnv1Uhcq78SbFyI76LrpeiF7wzhTGerd2n+T+MgnjRKKTLhGqKo
Wi9zchLIbWslEvySI+AfqX+S5cKlE3XmkeuQW8omWzC1FMmI1xqwLzYc1IRvYo4N
MjyUXcRGJKibTmymJq33Aqi1PYBPV8xWI0THcyRLAkS6IiqPzivZeOo+kAu1lDgJ
g9uBP06F7tw11sXgv0gb4cPhvi+nOmR1d08UNmmr81Dtscc/eKJLXZMrwS5+C5BI
5M7rmaCbWlld5YN2AsG967leDC7MxoK6hmpfpL0Nr3HeR8Fr2b0Et82KsrISYSUt
fT5+ITFQ+4opha2FGOTSrk3xMX4ZA+OblU94Y8mdTOa9JNQQ77DsqqtI7TQBcBzB
3QssvXsqWLdVraf0OGSu5pjUUZQpO2Nf4+UtoNYkXP5D1YMcE/IyvAawszk0krlw
T5NFDL1TGnU4oQtNo4rFsQ2NTAxkEdMEyQ/9iZEET9nZYEMI46XsRGrqCJ5hPAkQ
QXbJ7amcaM23UrZcpU9oNRtZa5uOt+AcPLwSa9Y3LjpYbhjJlfZexBFrSqAYRTsx
zL2CWo4vSunVO6mRMN1tCW2WfDtWPS0vrY4Uarjl4n3xIB++48R8MszvIJK2zySd
WVJxkbz8tLYh3TfNyqfUIu0MJ/OQ6daWaopxB6j/tss7+Kl7B/4QHWmaKxNiXkFQ
BVX1n5ck6U/ehm91QCtxYgjcy1mHzbySqnSzejHol1nnSKZAPy54/6T3rQllQmA0
3iJVO35mZ4V4WxpKPbyb+XgceG0ub3Gt8/ZLWJ77Q+rGQjlhifxctSsiroKU4HXE
K9Gd408JFjhZWQm8zwKMHTN/It2/L382kIA0GChudvH5LhWZsdhESwR56OdtItwu
kT+uHtReoWh3y3rfh09yJYhqMhIm4BSicP60u9p1RP/9wKIALnhsJN2Yw3l6V5/m
YMSQpBsiFb/FpbaefyR1lXuCTJ5Gnvz0Nlxx4Pfw0lh2RsUNa//dFYqt2qns1GLw
bQvAZ2ZLzjolY9hgAP5Iux5viSP4TE7kcUZLZFRLShaku+vG5e7YcU2MnlixFVjt
Z5TgScJtIcR2/qnU4F8nly50ywlszIdQMOp9tftxfJaeYAALeEgIVDmUeOU5iBr2
6cI3BXikTYWu/Z880ZOBTl5hw3ZyJXCYE5Ls99kUZLY2lS6haz3ijwffUpa4mKGs
wYXigZ2GhqR+dYoibNDHEpK8MTgw+Liz8+HXR+YajyKLdCj51pFGDirZUm060wG8
WXFaXxj4+BiKAOc2J4AJFIu3kFDDxWFRlCzVGuRbV/RCY4hic41dsAkkGbGhBfK5
CYjn1gCzTCx2moMENuHCjzu3tGfVy/jtJr10ilsyGh0dYiAaGa6y/8XYVn9GW8f+
6NzqBRvHfGVWoZFi1n8Lv46UYcvG3EqyZ+3iDdNqaiOTbNKHGOpBbpxQnTW8wd5l
XAulEH6zuk+G1fJRpSLWsfR4n4Wf9VuwpYXWrlyq5mWkDQuPedba+pdh41RA+ljM
kDJ6fJsnT1kGt3SkeMy9NyH9AyssUsLGBTgxueXkMp30ZIa1GnHpXj9w5JxctAEO
gg/NqmDOUTBfTiqURDll2tjva+zz+0IjbjdQSUnGBMFPcfSkh3WRGUcDWTe66qjk
gpXpSl9kvvSqtgJ9TJLHpck26BaP8PnYrqT9v/lA+wRJMiefx5VYxlhNFs/rBt+q
NP/zXBhu+SGsbBcVeF+QNv55aUHPPi51z9g2tt+YJ5C4mdtBHeZTTFI/NJj3dets
Jk242lAo4Hi0f7q8VlcGYpONczEIs47Mq/PmvaQoCWb4mBjfLhL8sj6OfIzYYMaL
vAmYUzwakBM/nj5yq2AbUP0knUEED4+VsGIpDVLnc67Zl2PywAFCCP741CSaocTp
X17Q5bpUeRT79ETm552MWAMrID7GJ6ehDHfzMczsB10BWHIfu/aEyke6AKTe55j4
1aDMqx0wstnDVy8evXwBagNk1w8TjfbgRy4j8MlwEykKyiz4LFXFrzSl5fu4C1QT
DFd7fRzWDkj+4YsoFz0wiXgJbLOdgXLeDA6RLdUF4sNWEH1rb+5mEpzPgUb9/XSc
6sHacLn5mmWo0vOQ38nyi/bIdg0itih3Tq8rMqbvM4I90wz7ytx4p0FCnrQmewjv
cSOBoQrlDRNg7w2fTy+3zosEQU1Q2Ke24jbSm/yd2bYKh9PRRNvfNwVVQtZ0KOvn
4jJ6rmUKLMoXgFKTMVTXBbPnap7hM0vx4grPQ01+YlDsl1PPJ4si2JRoODEMpyt9
4ZdkkYVOyUMOy4Qih7EXPPx1zOX7uICOyv3FiNAB2MnUDU9sSjM/jYKsfzTGbBlR
vkWmAmwd83+J6Bzk75mF57VW+1Er5NSfzKJvjNnfhvHcQBOAu+M7Vb//x2NnMSlc
qpbkzkEVcvliNrioDQmGYeEitN5wQpJXDIzlYFJ7s0BPWLAD6Vj0gadAZSsTgDwU
X/08VWIO4k5KcxoLpe3PINXbqjuvDAfkXDpwXsp5DAeEEro3cfFulCvQ3XPhYYkv
h8AWzWaBFRHXrJUiNW0LHgQ3EkeSeCpWdeaqI+7n5/2dv2vRhChD4nQSw6foUmVT
/AHlIr/5Ok4e3wZM+TP9lLB4WbaiMidXsgV4rpo1ZsRHPOUbqSNWZKJDMHZ1xquH
r5Jab27w2h7IVHMfb7NXlMyJ2KNJgJmY5BZwaOujjEhdEh8P5+cjPpuQpOgL3qhK
mu7bZuFy9UuaeoduLVDHUnZ8xTX6p9/dl78WjZX3gz0++HAGGEpdai/YBWpxlcMN
sHgpwjWarXTBPpGpcnIDnUMo8p7LaKGuPF/C3fccv8aysbuZxNuK5gVX9xTylTUP
71CtBVl2qbcT+aLeXVM9kR5bUsrsZgLyRQnUlTO71/GBF287gYMxsos9DzTKIM+a
HfBt8s9TEfGqJk3QcbnMn8mXBG7Wd5+thDijaj2pMdMkpfPr0m72VsnOmyQlnvUQ
LsKXAP6xRrTHVCqUdHhjcU7fG4qoPxdOeSvwvoPm7npjScNjXY3AZ4qIDfyJmmTR
TIwLcZhjgJIda0cg9lESj/4VdTjmL5WMuO6LbMQ8cjaD8S1xSbX2zwBE+Fxeo83G
T6ODSk0modTwOlrMqh2hSYBBU8XgYCzKEYQCAc1A6KKz5egkixhjlATEm1/e/oDw
ayPdBbl5euO+7mbOaHMFxmKCmJ7hFeYSaMqGzs/c3kakPR09GTFlN9T5apW8b/HJ
DLnRJN3L45jddiIINqVtiNoPEfByEaZ5Lr4mOprBrUdF0GPcvIwODIJS9S8Zr9XC
HBfmDEXmv0WyHlpcX/sQIvSK66ltED0Ds7IBPmBMRO8xqMRr3XLcl71bh8cKrzgF
W5BWeCLFFn/GHWfM8N8eB6yLdecOVDtYFsBKeDR33TUh8sJ8vppnCfasZyiORPPi
CY2pXQL0AeXB/5Oeq5QfQOOmOOODERfR2zqH5fhitFmDCL2cf0Ud6pPyRVOxY1c5
ROd0t+UPO3H7sTXGgXz+AwuIUV1GrncQrpT2zuHheH7TgUIM6fOj4SO5ZwN0adGN
o37D50EAClvffWdjp1/s9g+OAFozcBdJESMYK4sg9A0q8Z7Xm+sMWlT39CSfeNK0
j5jHtgaMU/SXpRTAqeNUUZsQFQ0j4YUH1w7Xd5a4/RX7ewuRoS4zB3DijaxwrgOh
hRSQbjzKwb5A8vGIcQoa0UZh5gm/X9PvUpz5xp6vSJjjwTcIQWZCfGhEdWlziObQ
VksyTanVhYwkDMG90+FsAtNjQPRvSgT2xU7t6U/dmbUPWnO3oGpTtWU6nsGT0nFG
99rV8bVvWfkm5PBIYd9OIq2rpd2NXuCUkhkthgPBynec29z2m+CQnobPvApPuiFx
AgfZ55K9y08k+t/eC2rgg/ldArPjsQxpHRSqFYEltdx1IvrYdbINWtMXroCnbO+s
wbQIsMjj+575qwyD+F2s3bFXkOb/aRy5F3gnAVfVytdNV2b9qfER6EGD+zPkSjtU
Ds2LFNZdNB5bXa2CkYLIoDNi7rbO3AJJAT0x/k0TXHeAUz5K+IXYpmGRa+iEMUwx
YZ0ewpUIQixGSMwnI37syLjPqbNgzhNOKs9CRSGD9CWiey1zIaA8gniI3oGNzf1G
R9G0I/jFNMPWW5PDvRw/kwcsyZEBfbeFCNySZl/nE5GDSBL9qY7Ks0DFVSnG+nkp
VvvHoIuyqrWGvSCq5DMAhG5S4KQLFyvuqSghZ9Z1Py7OOrPkN9NtbhStKe9/Nmkq
fB4mBw6Sc7tC0RD/UYU8OYc0HzBiw9Sbvq1Wdi/To4kElowVlg9rB2QipKOb0aFx
O99s5eQ8EAeRdwIIbTKR3aVy5YapqfYOHusoXrWQtSf9xPmqsPA8wULZQAJUkNNS
S2D64kpVNj2GPrzgRaRVbVyqSVtTmKj9RNpBZOgm0gjYBXvuoq3U4Q4BdaK9xgPD
NexnFcWkbgIn+pDslM7N9AfO0tinbYzMtwuC3eMeQAky993uvIuN+kblR/UfiZMn
kmjTRiRz98A15HZK0sL4BDo2yK1NIlM6nSjkAIfAMGH0hwBmgNirONvXjOVF6wq1
N0Jqg3V9dW5K7obIBZ/MR99pwUnjvpbF0eJmkSRCwjc6uXyyWMt9ERwdg7sLtGys
IldQZqjGNZQbdSqoocOp/9xhtwx/Nr2HddvD8RG+h7IRmvwwRbLjIZbTdA2VrbJt
9iBIPcQyj15ZN3H7SrAO5t2GjRHEjY9dduYrnmH7nU2rly1dpCIET43XfcXoqoXt
B0I6knG7vv0MqrF/s/nnAqnvVWzR4xmsG+mkrfiSsOLNP3CxlMjJpzD5CgJKIzYk
Y+P3tImdmVWI8uJ7Gb6m/QyKGbuf7Hfwmigji6XjaFruXYmnw2VGasl+qfLak1Ap
OoVcsagk9imcIEUxbT2+Rz6PdSXJX3VNTqCWNLIyCFgh2ftihKeTxTP1N1vGO9hW
/PCDRJD+JIsbIaPWWtkeDTPX2tLqGm7F1XFN+7hotUzUZV/9airrk2ZSW2gbz3n9
W6DH6Cz2Yk8JaTqPIckOmheSd5hVtMhVghROHeupGyqzZ3BnE1nHntRcCE+cn1Gv
i0hmsb8aR3D07SEcAqB1nST5x2vKuXQD9CgZrO7RnB+8AiRZyc3Cm9lF98PyiySB
SBoQI6S4f09TY1S2t7ubarRUIMwdflu0SXXqLtYMS2x33YR76FSJvCWjwSU2upMY
2l8P41x2Z5NWtOT2mXJGpVTYS0vuXW/ToyBFQe9KANErrQwA+6/IEW2HVQUgFOy7
gqgrYUKsyt8/ea7CrHkvlIle2N1JK4dmSOTTokx81rx5BjrgJSXejLP+HYU7cy68
qBwM7rT7ue1zYNSFpMuh8QgE89aSMUVf44+cRoSYivNJm3ekRGWxMm+94r6hawY2
Xz1N05G2atx0xPzx4ADNm7xX3IobTRbkfxHQz2954tPuXc+SCwD8OiS36FFswVcM
qseFq1ZCgB+3cTiEnbraFynf24FzlwQC4GYC46f3t4wftt8+t/JUdyWtuarvmm9G
53EQK3xOqj4SPu1g9rX4nM+RZEsiRsfsWcGcD3p4rl9iyx0bF3T0bhiXxmwCaDQ7
mGPWEiIyXtkjArwXy7t79YHNicNikldrvEUZumi98dZlrCL4/Dgm6Yw5iRhlagOR
mDuiZIkxg/45zZzIHajwq+I00y8teqLNcHlgMweyrAbuDfxNAAl6nqBC/IbwpOrn
OuQukqrYdMf/Qnw7Mz1NZM3w1adBjV5D7h4cRSrmv+sdO7jvG5HT11+14mivBU9p
m1Er+DfBYGV81x8Qs0Cij6G5DdHcISDMDvAKXX6UYhb96fKkSlc7xRNnQSJZ0vYZ
2fq7r9j1SCeJS7FiwbfjHshXkARUhrVIfH7hSlnE8PH/NVHkZkmobYPTFxuuwXyH
e/g9gt440LCiRzu1PgFAPRu+yQIvEl44JPmlBQmTDEd2gFB9WAaaSfu6UzbnMIDy
xFXFwntPIfOb9CbSbHm/9hVvU9qqDQ0kBsOduABx//S7B3YP/htvkNsTtSZGJ254
JD8aQ4dYB5WbRtY+GnQmBm5/Ktc/Ysv+J3JGEKnWiR1mEoflUBBUKUfHPKeMORqA
Gl944SWp5BUOelGVDZfItJ8dNqP+L79UQMzK6S15im0mmq9B7fYfVKqHymqC6P8n
4qdMO+HJq9Eh24Woj83PCYkuLr/c5Gvh+VJPHpmt7e4QCUfOtTln4rr5o5e6ofUZ
2R6b6ec9O98Z1u4h1A7/Q5gq4VW7+Wod81Ls/H4tiNsaAWq9PnXD0nxNLdlY1aFo
g9M6cvfNDIGOm/qE9IEVPnNIjol7hbSJQ14SW7u0JKj8iMSUCNXlxJwhryr1HkbJ
yUGDZNsESNlLKl36RXw+8CZaZ1S509pR2oN0FXQvanPdJ2K4YDLjBoNQV75mipCw
ae2vJSWVEVSKXjLbycP10hN4iVjVCyZAmIKR/+mS769K0NYvfPH9l/qjHbT+ylfq
sDwcA0RYbHXCSLBNhP6F5WE7WQzInaSJuXvYfO7g3SFYzA8H+WkgvPZudG2nzZjl
KY5Wro7ejP+iyHUfEtORfKnCVCjWrqHXkts4jOUGwmy/0r1mDdjlsXLUyhmQZr2l
RHH6nOKO/Yjptk58zGw1FLsV7/qLOehfW/AEo/5ha9gq8ZPMIgflBOzeu+MMaWZ4
e0/+k/iim4aQ4FtbODGKTB2Mmfr0RdSjw6Pxbrv0XTCEk2r2fbsO/1jzd9eBi4cA
QdRQ2CJERcO3K6NXVtWA8NSuSudkXjzPTz3ViDRpILZu3hehnpNZSlh/qtC5CcQM
TQFbM5ZS5PATdz2e0GJbKETA59ehNiier5vOjkAnaS9Vd4MkhunYyyOL7ujQvySx
eArviotE1QIgobvkiUriFOwZj/oZY9UTbvrCmxvE1z+Jrz9doznnPPnmEvzEt3yy
GRLe1IjE0pthQlDlOnGt/eUMn91EJU4bZJI5SERjZX0BLyFiRJx6/e960D4AiBfB
+92h48NqNctEZfXI+w/UAgwXyfsTPV7Q7B8Xm7mfdGPhUvNuBGmeUXOAIlTJIaYR
ZPS0LUT9UuNiiB7AmTUqGweJZOrpdYEPAOhgn+nEzQijwyC6cLinKWzNL26VEeg+
4LAg+C6paE6GAKZCO13a3udUXsftKulxarg71V7cI+AP9/6Vdb5d+lDbm2nS/R3G
qyzqtFyyXkjSKcZvvFr++DEACuXxDznhZJ1crEkYWh4YH+xb5+meyu3xmeAA+lPN
hv1kGWWaZ3xel9mydo8aVazce436uLJUGPbpPfv2SNtxxB93J9fV7XxTq1Gv5SKu
ZRrtgIVJr+qbbiGFavVrAC7L6zntM3M5x9J5+A9IpqcZ0RYrMW7i+nE5SVWXdLuJ
vA0aNdz2RlDS4Bi1qmhe7KJnjQ60J9x93ZtVezcrqCkmizbRwItx+B6SqVbbw7DU
qU9eQDKrUIt/eDLacV77TGp+Onhcp6KjbxvDZzIqh7Avwp2WiXoyR6IqF8TKNgGh
tqV/pXTlpIkyZyvYn5Pw5hnAqJmxgQIwogxpSN5xaRU7bIIuS6cUFYLD9E1plyZs
nBAaJtHiDpv8U9I8arl99kqChBkJDkuTXuoNeKZ1TFYHzJjJksxmnjbGsno/Qwcv
h+5/CaUyBFY/9Yp/W2jSvrYc1iqXpwh3UL4UqyZvh7UK74oPjPzFslaSopE6o12C
W+ve3UNmLnfRlKjBQPLZdjcy+qVKJEdXaNOOmANCKJuflJ/lQj4FPhhprFRSi2W4
TpqQSURW0O1wxLFBBQErQ+tHinbyHkGvbDD0cvZ0vX7tb8v44Aw0S8UDjK/IOqpI
i9/JiZ3kH1O8ue1kY31lB48k33uu/3sOWNmQqff2bjWlXruN4XzTbTs6MRDxk6yt
mBFcpN5KPQ0i3uiByrUWH9DVViFuvgMUOEApPo7cVRde+mAe4N5CRrmLkgvvFQ4t
fmq36hXw1IHLMIuwoIsi7Qdr1RY0qZ2sWXq3MpRrXei+HMyt5rJIXpXUESU/teAU
UXUYmOCMNmGsMt+3aGBAN2XelFJ7ergcm8abLztchd6krAAjTZCRhXw2/b5S2dKQ
IiUGlY1uHPKydkJjj112Tp7JEEPjA2LKTx82LGH2jmHPiTz0Ds1p/YeAg+Kgau1t
I+q0G7U3Ht0l9LF/8t3JGzAvKHYfejJGa/XhvyQkHLxHEdCOYnpofeNK4Us/Y4YS
sroRGr2RF9f80cBZxxNrwtjlAg4Lv9ul3L/h+bYn5dgWL+lKOdLrFy6nOOwfD0KD
b1JgjEaS8rhtvVR6BTdQwDpxeUC3J07aXzp2MwI2lLtNFaMT+Fq37vrMI7G/JJ9g
HkKWkF+B5cmVRcYolXaKkrWsKy2/4BvdOELNXV96wBDJrdzbQdRSfM7i4W37uu6Q
uTY3cy8UmuYDGpx82lN4fZW3Y362EydDfFnVoAtXMlluf/rMTTarCLeSXqFcWB+q
1x7gcz02euHQdTBnsy9RadvZ+A/4YYv26lWV1lmUe7OjyIYuR0DwcRLhNXUtESQP
jlMeKdAdE44rY3OlX4jkgJbB6fJylQ5HnDVUnskTGCCwWacAQoZSbmrENLddfTYu
23zO7iD7a9tNASRdeeLUhQW3ZfGkUvv/RPBA0RTck1NexFiETI4ThLbFu5aLPXba
VkThghCQTW2ED4myLC5O4rZbHj+3ReSX2iuVKKRYfYRCMtMFQI9+WSghI0tuVpol
mEZx7T8SaVGChvl6ed1uC9DJhnSwYqPhXOC7lzIonuGv1I+9hGeYRcvYjRsBv3XP
+IRblyv4/F0zcO+eFe69mdBSuMi/Po3lMjEU5nfCYpYVa4c+q+d9sTA5TdgfwWZW
W9NHzXYS7v5L2G/aIiXJ6zH7aljtZeFrRnOJi7ouDC9rFtOX/xfCuZ1U980vKgpi
GqeJNKSut3k2lNi+b/ZD+LRxpzTCktDcEXhGgmuh5i1mm6eQgjLGYR5icNjyhKhW
+etkE2jRrajKPMekFp6xaTC0RsiSUtwg+XB3wdsMOPH1FIujZDSPis85eEhISrRS
UzQDYL/EiN6rjdpv4KQ7nS+jlFyteXku6H1fhQHqVI2b2f5kCoxik4siITwa97X5
FFB+LLpRPoetHMOSDLExruwOogWK3h9N8uHR3wAzjbs3szfYKfhfyeR+jALYqVIz
YqzpcV25TvygrZfIEvPaF8QnEOoKAarKaYe/iFEP8JmV2NwkcxMMnOr3w/wTGLHN
Wox2OzQ1Oq0xQBY9BOo4zmUKROBkF2f2HRflt+ypkqDAfhsgVjXDs0YJj/rVF8up
iea/8GrUYyGPneCSDJtdC0dVIYIrFXFcKex+hZ31pyVAhIEJ2L5bGsbYuhzNFCjM
FGULtU6V7YPP/4yHxF+SEzYVd1seuYLoHnfLtlJfBKJmnkHn8xgxAM/uJuvdzXfQ
PaHQ9E2W5ir1Xo6194WxS8AcGL3ItZQrtQr+i2fZRBuhheDXT6cpkSYfX8kwCXja
3J7SR2InikDy+NZ1WBrze14beMoTbq41a5oM0fx8vWn5G6UbH5IVl6URx0GckL+H
RWdqg9rsW3d/ojpbJA8ud/BGL34EUL+M+juJwy+S5PCf6MP3atq1mqGODmNEstHG
n3DcPlAfbjkLCc9oD2Y5/tjulguekPpk77d2q7CM/gAj7lOliHgwvT1mE7h/xwsQ
v6iX1HWfA8qXd91/tSiYz0EOIpdtdpu4Th5Qcjb7IMdhgC606KpqGSOBXgQU/pd1
zHSMtN5IB27x7Y5OQyUClQfVNCzDlXSd/kFMDSFNwHxFYoDdLmAL6PH7TxrUN2eV
soJ+ogn+HZLKtgjZW9waoB38p8Oj/oaQqBogUURKR8X/fg4tY1amtq8H6/u1aHX0
P78jjQqPt7vDAYdZ13UK7SI/Hl6o0VtUgjlLdUrqHxiX6Uhyqk5Ajag/60+EeirR
9+LngSOPVJyJ20kDXL4yBP36YZl8oR0AN3gE6wl9krALQJsLZuYIFsscqJunS5P0
xpUsVhbq4yCIAqwuFcNjybGTplAM3dec7d3iN5MyRVTpOkq1AVazlZz5QwZsbCN2
cEOdGAsGNoDF7lSClsYikTsdnicQi1EPM+lvI0/XwWKgIhjAWAZqlhxmlEZYDL/D
xgnQfUpIdN+HdTTorBz2H2/JO5/S6NDcUXhozJSB17Osd0UMMuHkYU5UAGFyigHy
ydqJvuUDGkWYQgLqFavTB/W9DV31Y3gpcqzxYwRJPOjLsdwYhkS+p5nfogHexYVI
6zfePQ4gucQoaxQQEiwPisGVgZnkKgrCVljTk7xRxuKzLb5uE0cycjTouxf2NrmJ
UtsszCZpSApPCmQaeC8pTrgUemrmDPc5007cXTBpHkO7cTPcl/qicHTlnJnGwsfK
NRqyblTJTbJYJKeMXpbegYIWySb5dyZcm4POtDqtjg9Kj5rcq+HhR0y2APOozFRx
RZmmA6IA58/htoZKTJ0Ww05Wt+ScxVXSNQVzcgVKTjih/h1E/H88FG7LKCC1uhrn
0XkUIpcOpTAnoiSBqD5EWPnSNf/oj3xvPfU6R34+rWBq91AZSYs9iCoorCzVYEpi
bUBl6h13ah1wKksWaR4UsBs7C+DQlNRPYagCYp59Rv+rBJjK9SbAx/ayGZP8G5xo
APJBUjPVigpbua5+sBjFg6bIm/KFYi39FDzCW7A0mV000UJdo7pEWAsmFQJETJ0/
ftG1/qCvaVnXpxpd9U4dEfu1i8JgS8XkwRe5oC3QKyAiFIye4ETkFi2vhoUhTUnT
mNZruCH6CDua3T3GEPPwQKzDKho5GbPNl4Xkrr4Zhv94XiNzswj/CmWxgTaSehR3
FLvem6NtohI5XE38Ojtn/eduotuasxfL0peY7+QxhYnD2oIQVqyAaIq5VV/mXNcB
Pq9v2OO+XQTGcI955Pev7lSOB6JWfBExzIFtXV24N3PGiszo7Vn4uMqrRAF++43l
jaUfd/XusoSGnPyjjb/ws3cWOWgh1G8EttRfJyKDzvfn/x5DNRlIJ4b6irQReuWO
ko2RH1IvIaiiNQnr60OOO+ra/jL7133EbJH8n65NMQcaHJpTYpED+9epxbAX4kny
F0ClB1WrVBEA5Y7T4hjXvLlpb28MCKS0lgNXy9dV0tpSJplePYtHrsi2jvEN4gmY
K2nlnsl4YvR991V/p5whN9nsR6SZ9NjaYYww1fc/gt7lN+7FBGZ1UjZXXmU8X6y7
WXVXBL4QP6qiGM3aR1OBKVU534ztJDrZbsF12k6w8GWhKpXv7yzd9uDJzYwLuA/7
NXyxjtnzhHV+OBTx619YJOhnZkiGk+C02EX8j1/XprsG0bcWGVHVBc3fkkQlmiMg
Ik7wr7ChpOorg7eVpH/fkADJigNPtFbiNHv6a8KKDSxhl7eMd1ipIfa8oOVFyYBI
CdwXv9itsvpSIJ3m1V0w6g==

`pragma protect end_protected
