// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
9mo/KXynJobWS1ORqrMo9RooILLAusbA+U1eGMO6FqV/SVPwM4gZgyHNflmLvvLD
xd8TVgkVjvGgdmYmw7b7iftSVrlto98X+JUVKKdSytZIknXE+x7L6Ev3oPibAUWH
tjhqBB5i4oNeDsodCVZ3vgcAPVqCVtLF1SJugZnMCeRkL0YYTFv+2Q==
//pragma protect end_key_block
//pragma protect digest_block
zTVGR3C1Xkfp/jYglb74Ixt14aw=
//pragma protect end_digest_block
//pragma protect data_block
uIDw5MACssY64UuoC3cHyknPYgHJoSEdcrZ7o9rjKwKqbVMYq6sKzrqOLzEioTxL
HMssNvNU23mHnxWKe67+Zn0Xm8yEkUEPDTZqg6a1KMe6eGAD1U5AMSubl/yYEirF
Q3QrjnmNpWC5yr5diB/fRDxkcfx44CE7HiA0Fzj16A6UDRwdd4Ym34bofRP1n4X1
1nJwYN/HFlFx67QJReNP41srvruQWsrF3lgJtJcZAkyAyl1lLj7TIw9ygTWWmByn
uZNf5vNI3TbMXW4EFX4O0FQ0F1ebsUKeYP/NIInIRlQQYocT7bdJ4ulywDLFU04H
8DHNh192HAIZUw6NHHtHC3lv/edwgb43r8vUBaMVza5nGmlAgaQdsX9Iii1r+GVg
+9FQAc3uLyfxXEdH/orkVRhK9Aqx5jaOIMeMPEQvKVqSshWeCMJ/66wss8k0NEXc
GwYU3OhAv0Lj1tzcy67HXyZFerM59MjJGXkSTvdLD81h5OShL/phTnSTQ05hC1CH
5wO4HqBJNTiXmrm+26y67b49nvfpTpv11Y4IU/s7xxLEqxEH8Nbcb9DDSqGbfUgi
hbD022yD2xx/t+yvpCL5IDfYLPQrRHY+BEBoMo50QkHnVctytix5jle6Q/NTApwM
P8fhjuQxL8wYfQXIPIVZ54jUJyA/o0GZf1dTmhhKIFV9rAAfCGqfOmo/fOVAki2z
4ty41JEf8MF7Cegplgytxhg7Kz5pK0Ftb2iaEiO+cDoMEWXdlTzJOygLI2AHSXB4
+iKP1cWDPGs/cOts/Sqjn5Uf7q+rjvwZ/u4+R8EAiwdo71dIo4vfEyQO1O9TDBxv
3tGNhd9nAgdVUsj32ywuitl3aiCfkETkBw1VybE3MJUHaVAnq1sEMornTudmhgQu
4Txku5l6qC7lnK8Q29135EdzoE98RsDoKL0IkWT9ScaC9zv7OTUtp7vAfKvhy75Q
ntAzxRk6wLVZylAEVmHOjA0yh2lJ7dQg9sD0NgaufkxLbpdX375LLDwiCmgz6wuY
h9LTuVf5U4EXOyW9hbeVlJBtJgTL3nrAA4Fqj6nGhKyBJJ6UxxnEZESo+nzCIFZr
5BdRpaZv5lnmThhnNtxuS/1a6ZzsnEYKepVIqn5wNsk2ForHQwC7+HAXgkXnt/yY
kAr7A0DX4Z6bQw9HlTEuAYiDgOu6Ff+vPgRZC7ec3sCXlnSJ9dqipVeJJy6irm/t
hmxaNvdsSYgnpvRmifGZ8FqjAhkhlRsk3TlgZ5E5bGhne41r93nt1yRbGcPlEGQO
FbcREubh+blblM2S+3yJapuPHhX/a5mHhDtAUfU1cAWMPAB+c3yP9d/cDTXTfl3w
G0QhXJyjnPtyiFV38xMEEN6uv7qoNa0/StcE5uyYENjbhR8XShUvCLiz0vZiOfeJ
ix6NeTEj4OG/scdjioaseNW4T2BpqFVEM4++Np4A+kjKq5tG37HOmtG+AXYuiogT
0taGKWa9/H1+scaeZV5FDTViZYSJ4CZs4bi6hZvwGQZI0PJdm+LtcAQ5LSfiw9Jf
5KVQ5yzzbET6q8AVgWNg2rKRkFLHiUlyNC5J1zNIngJR1KL54TQ5QulqDGfW9Paj
SbDQXcUKSAVeRerfPaC+28Aw8I8goXPnzqfYxt2PRyrOPMkjMzrJeMkfdY6x7Dnm
BUzFJ5bwJQxVXwmPyu3Jnp9I1nN6A4NjAvyRrT8kKhQZFgu4T5pjQa7W3xu/4VYz
HQwLhzAbof1zZS2ErPMPCExprqXXSzn5AzqO0JHMADiHiuDaaiBMhYNcmRcBNaJw
wPFj7VDXV8jkjLEdN9aiPSs6K5pRN7nChWyJPXRr8vAk2gj+OusgclEAxgCFL74k
aDCA2vnYVxBeZ9wR7H6cS4sp3ZkhNY1YkuwxOv0v6X1Ghg147zvt1smpqPrl0dDq
UQtU8ncdLPuRE5RpUQcv1bbuB36CdZ+AJEIigJnHlgV7qbODpea6XN+fjST6Rt64
YFpcrVbTKlGa7CSKZlK+BOE4L96JX8DllBi0aWoZBbQbwqbwyOllJlq/4QvzzStI
ZpZdpjY/hFvHAEsKugYTLpPOIt7opbaQ72SeYYRkBu/fpEuu+ZJzErG0t7T6o/4T
nneYPx6Zbw8lRX2d2ar207DIBfmwVUjSgjeBmkBoAL+ELb9WNxuZ9CTGYmeu7fgu
a27FtHQ/PKaXFoxZ7xJJNiU9ktaxeFEPCGf6quUhrVt7gurVV7nIHyo5Oci544U/
8vHmBg3f9KuDdYI4iECYlvhvYDJT9o7fX1WiyTp5OYVwUuwFsAAVAEhoDuFSFSS5
oRSkPw4EXllCUradkujLH970gwFWLyca9go0uEsM2DKU+iNxVmTwlfREYdMEGDgW
Op1KMKeMWvTMdjzPGgFmfd22c8kYxSI5sLfdKmtGAxh4pYYZixoddtinlm+QN7Sz
G0hhTPLubmqsyWP3UsKEO+3gB0hRkk3e/O35k4qqf9yhkECy1QT5KpMGFDIGl/6a
KKcHdh3MoJZJyy924bUFsFf6x0ai4cfXtVe/VInKpXiU8rIqTNi4EPghZP9Krv3P
uYUpP2xjtc4W69xuaIXTBo3pWizTlUHUF4SxzdHGPXB9WokqD867nGvRQ1m1pb0g
C2CuYhrbbXWk/FrkoZe8iLZCw5M4M8RZOCvhIz6cgIdS6H6S2FRfetE09HEUCi1M
Dyr27LBsKa1NZvMEWKyDKLizUe6tycvkHUdoRuoGPFzu0TGsosKLh7KRnON2rkPm
WzuTDRoJCWyMByolgdLuSutQEhbS0xvweJ01+Wsy5ahXW1M25b7S/g6sYwP1JKoy
GSqM9sC/8+dX/fptFUw3LNZJ14OIP0YVK/o90N4WSVi8b1nsQKSKDY/Iczng4G4T
X9IkUMOonFqB5KiFTgTQn0eFXSsE3+B4IJeCPeEwmkkte5/24I4YIOQSlFWzDD1j
Tr76RcZKwsqSnhJZM7OhLmAujc+dBTipBnoBj6+MvhYZnJC73pXRGpg/5zEI6QdE
KXS/6JcrLicurg+DRhocxMVsgVHfE7ulWDBdoOEw8NZYeM3nUN+nnrZVqfUBWEzd
eLfxqCJePz5oM3z+0TyUDJ7/LDUCyYKZXn3xosGws7sKAk/4uKSGdGAA5y2Uzsxd
sxWBfZJ+Wded/pj2zaPUOEk73lnsXt7g836aJ3UmOBxv8AxlkvkhGbdtieasFtJI
jGsF+QWkqSebCgOCkSyqIuzxnE+yJD7QtcuYwWE0VvRHIZHG2E958QE100lzLPDh
ZTen9T/DGvpkcMBMfB7dYQ9YRy5J03Rs+pZcSCP6UCaqdWoD3M45zjidAL0zU4FE
oEAVX2zK+Yww2Pee6aKz+TCY0eN0tifN1nVmmrXhknkrjpEDhnKilAOMo1YYBdAm
WPtiFlm8+knepLJ5WchXC3bqYB4WOdb4pM5hqe4n+5f/bGAbpHAfoepta92OK8GF
wKyuiNyoaYWpM5PWRQCtopWgWRVHmq8FC0B0DfNS0kZ3EaNiNFtO2PqEnqvqRKFt
XERCktwiNoGnoZvcACHE8YrAmL/SSu2bnyzsRxcsHZbEiGIoFkCe2ae/mHO6d5Lp
Gi817beZCubirNFNmXNE2W/004U1jsTNqsrhU5ClwYRgQzwAsrBeotBQkQ56gITp
fCrmK1N8EsZYJGqG3ssjkQ3r5j4WbmNya4Jrb6gff2qpQz8xRQ80xNYOck6MgICE
8jTsMNeS2gYti+NMJb1YVfbVAQkSbwIeTpLpImu/HPq8WnQpG8WJVIw8yiWc1Zhv
JbqA7AulQO3IFiBOAkEwFOofdhH45BuuuXxGHgVktnZX4LacOGgGhI+uoDafrSBQ
BRd7ieBAaP2jKB9omIJzkgbq5mpRW/qyBK19cOArd3qoGyj4qKixmBr7zYfMPkEE
zMPlylKn7yw1iTS0jtAoZiaSgb0saBgUWCdkvx5AOOOedIJR2QNFFY6qso0Dex6H
1FKhvGrsJTAzbIB/zj4r3lJ2NEXyEit1yYa2MrZvfFSJuxiJQUcStcixY4Y6NEHd
4ADG1d03mMIZ9snmKSiCMjsYra//x8hP0HHE+PH8tLLNz5WltS7XNj38iAveyibW
Nybm6iVOW3+Y3HH7j4CAqbiBIKxHYZwe6fCTXZVQvxIrIS5kdlpENFY605mKxeaz
RvMjGT8bQa/O6Q5En4g2H49TnOjW40uSxvVkiqINKr+LX4MdrwcCi6TlIp7AfGiL
nuawIIoyJ/fxghhYmdCnTCuKSqAaCxbIySjth9TQgoxTkmE7EHYOkGJa3mj6UGTf
CPsy9liYtp/KBIMibbER5rRTU7o6Sj/NTyrXfeFSnaUVYCvrV6zxgB2A7RAPf9iV
lk0oVgJuHnPYQUxj0QYCJHO0zO74P4ryF4P/gbbGbwmiDs0u00v82IdaCYQe1b1l
u1yzkuyLjjXWy9oz4awKJjpmY/867PsqyqvViXzDgj5Furr+Oe5JktRc447z7vYQ
94pgwLxpjt7XeJuFzRhR/ENWuCzG2J8T5ENrmx6oFsJTI/mYQHImLBEXxnbxVLQ5
f32A3SNPyCY/h9ffUoRavdjuBKGU266Hx1F9FIFXVSbCDLSDDsfHD5kWYePyAegP
kS7Ml+IbcS73Y96kN0cle65o+6oyBK016pbVWJB/NxVEWCmsDt3hQG8AgLUVxkdg
wFlSiU24xPm1G55ejYd0ixOQwb+XlryZh2qhul0z1EorifEKCETHdqNQTyiCyxoP
CK56oMlr4/QHIRoo9RX4sSJtp40H1ARa2P6SBG2tF0C6HQrKfd8hOHQ++f2qajfJ
QdCtOd1CNu8QcQSFFqz+wjJOp88bW0JfWco8Hti9iKHRiKpot6a9THIzrxoVc+Wd
f9GL+BmlEOxs0QpaVO+1XopRxjMuh8N8LFE3ljcRoa38Hf4XxxajfJwJYs4FJk+I
5xGYfDCD/iaekxp1cBKB6d3/PdRGyGck0BuiuzDtnCxTWwlMw2rep9RUlHl+tPkZ
Jm1BAdPgrr0W5Urc4jRohj0O350cyHsgFQZz6Vgczsc7Pld0CLOd20XzVqMuNJDM
ojFBUvX33dfG9YEk2k0WHJt5UDSRpxageKkVhlItOpz8yB/TeQe7omvbuu3SbFGa
nPQcEmTCC6YXaXQ92AsN1+W55YlobaszRT41R34OpvFKtMF3YlfutR21rLPxQJ1M
fChql6HHL/RE8ifJaRO35JE3winhqof3y1Djqe7S9jDMHo7eWYErvX7DTNZXePET
X6dFBFBs2nm9VJT/01Q5XkWmo5HbWfsqvdOJD3PY+dQDZH6jDdC3Vf00IdBLf10R
QQtIdC+6ECpodkE395iO/RzJ9rHPJdl8FQGCamDRU+WXAG6LO7dWEp+sAgd4kP2s
ZB+kS+zB1w0kbvI9Acz4Uzj0HjGn5hBaVxVl5j6he8+ldeMWtP69wNOH09wKmMDM
rnRrRdcxG06r39qJ2dDC8j2U7UTL9MfMJDleG0WEXWVouPTkyKrHXoy21Z/Zr0Pq
N43H3z6BO2wx4iUmopkQHcR9cpYFwop4xs8P05wKhVl5Gw0VUsxD2ZIfGfmlMsD6
8Xz6SvjKG1B+Gi7oy6PbkfMv/74OzEZlP0nKFRgd2ZbcaJjAkiOiqchcwfAwpvCG
Slih6v0z7Am/wd2Ea5BGCmudP7EbAX2qzGsEpO9S73N36f+oxlKhpD6VHZ5m3GOu
zQtoTPHulBjd24EgZxIHlzG5dF54ZG09FTy94MkG9IKY5w08mzwyCe2KBeTgOIRS
/0wQZNRwt1rJL2UbMaaNaPzULXVp2pnRqcI1iPx5J7jAXeGn1tPZVgImMdJ5hYux
LshYcv9GTA7oVqTBeIHr+Ff1qMjTXruJR1cRvZBppMbZy/kEp+RPAC8SuIZZIfbw
RjaNNUiKUfhEstz0uw60eaeVYQY7Q+unf3RzZvvvunR+7uqbayFVJIDM9UW56MqR
Ghyigzbozyq41+yrThg2r/WotCFnu9pflAxC/SUxJNQZyzc2F6W0PYnj1qlwgCS2
sKNpIPUl2LhmnOytf+vucwdKKJNzuZDXdii6b53RWsDYD6yFdsbZoGHvvjjHLbCv
kF5tvbG0Qh8N9GD4H+PXrGZil72ZgnfKNyoDb9cm3VZfhfNRtuuIP8I54p1ObLI2
o6coPab9TTkXjSzZjldSnAM7o8kT+9sS7QWRzrMRQWyO0JrFiwoDQQMZl9UYKfkZ
a9QF8zpRaY5E1U3lV1/8GXNNGJ0Oe4UM0FGt6yA1Yrv7CRnguVh5NGryJ0X/heRw
S21MPFuamb/ZGW+6IrFrNKdW20obTHmv758mDclGGF0J0cwTDN17KaOyE5iM1vme
+zeJ/iOtwJzqcMl+vjKYbZ0Q16PcNsczLCENfBJ2VjAHnHFXxyGQl5NWXaVfMKvF
ZZ9bwasbfL5X+kZTrByUfSGaVvh5q5TY6MR5Ewbhn/1o3sNl/bWQYdWteDbLtlns
R1//x7wSxHI8qTBGKHxE6wDN4ZU2ZP7IN1jZbyNtBULmYMkTkFN6/pEPiv7aN9YS
c8WfIs+i9OEHoE3Y+A7zDHdW1A5aQ3x/Y2H6y0p7vdJ0sryJGaRwhTOv0JoyVoCP
1GGIA7o9lUf4hmHJSu0UM7OuA7BwdMsdc+vSPRfvPQSLoseW5PHT6dF9cXQ1y51y
/QwTBBz6ZsEIEf5DrtIGn5v7N1VGkkLyEamTnE+wqIxYFicFn5Wr9ZvXKjDWDnjd
CNrEWN2UBN2sltUT+2/cGa47P0F0xUHMX4A9wty6etiuvbZVe7rEpmntbRxR1LPf
bfDXPTjqbBFnvKxtM89e0uI68kDzIRfhoxd/U2vPPHN1lxXls3uXSd4qZLzJv7ZP
/eYDVx3H0/Y5WiCDyPM52uti1MTuLBT7ybtRNB7b0PcaNCPMKQhD/bztKh4smSFG
y4YV0eEVurmT8teGAaMthDSQ0qOLexIENESYH5RJT90gDz01XF3HI1X8EOkPQBhG
Rvm79BTaWuJ5lDOj773FtUwC217wOL3NPXJLdViWSqTJqyc/9VopSzdbAHmnLEEK
12yyJgczGMLFGR1F3bI/3Lh/fdS6emr1GS6bezKSJX2m8VGV0sR+ZNZaLMXRCmh1
yqrPyng/LNZ+YlgNenRG4PKxH+3BfnzbnGaCU34k0SRQjSYeotdByzEdq65tTVQ3
iCX8pfeMKmQf6G71sl8mpVkkFJzNbJm6vJeWyU+pz93IHQofYQKvVg8wL7T9h6W5
6pqhIXZZX4yNJe4sv4YrLZBoHHugulBC/66Y6xekrgOQLoueeuT+g+I1NyQ1wJej
XT9nz+zbar01HcuQ3bjUt4iwJ83NItH4X0YYqNq2//8tdUFZPFrpPmatkldYJwPx
VA8hDQ6ZyjISI8I8vM6c2LriC83pDdqbYOgnniYjzJEpIGKY+IML0FGeh2WhdD4O
mDr8KvFcDPRlJbytPx1PGEdvrrK1o9GeRQPFFX/69n1yyxYal1XQxcI7uTopDseg
qtfTnjfrzLP5rEhMQC9Gq4o+u7t6ax9Y80UtJSo6WYNZtzoYVMciA6DwLgsXjbgR
gpLd4kXuXqGyrr0EWsK2Omj5gVYGjZS5gk1ShYjd68tnPGZJ6ZdVDtOTpH/WDyzx
9BuMfjBjh/lLpCq4JssvV67eK19OLUm3BZLTPC6fH2yVD/CsQ9rxtV4j8dI/iXOn
MNWUPnBZumyO9fMovZeeMdg4Hdl65b1ebQOAGVP7ocIjpKFg5Wg6RbzMCSH+adiJ
pHZJlSdp22Mtk1myZPhxZ0lQBt6gNwx2rOsUap1fk4sn/JuhTEGud0StF7j7R949
bCEk3dyMAWmlmqxMNrAKuIpEy0zkb3RGP75Z2xaL0i2qvfXKcY4jI55nz+fG3VQ2
6G5JzT8ZQqXzraGqPbYP/LNNArZcLTVL9nxDVaFZxo36QzL+8q5Tu7J3YgiPL5iZ
xC9+JsMVelM0WtYDtlZ4dyc6S8c0+yRNypNzaZR53EBsQLJzyDRAV4IFBbapnkDf
n8GNrygMmJubG6VdmrHcWVwOpf/QEYezWwx8PfxvZhtGXvLbUugLYdUEht59i5E2
Flj1NE/yupOxMlzbKFE86MLXzmdm77BZuWC0ufZ3mtMvUz7RyLg0U25n/8oyPZAj
NqKnehKxcfKmAsIUARtMin526DxsoG9LEVtmgnNwSYBSgiNCztRl9ZErRXdOz6Mb
NBI3TMt5EJR65tOdtCyS0v2mg1rrhFuTirnk2MaCENHeOUk0Pt1+XBD5gaNtdJ4v
D5XbhEtwsO5qHk2O9ScSajbKNIy/lAeULfu9b/UG8cdDgk1wHo4Pge0LSy/uWLd7
5J8xP60lzy9LVs+d7fBd9zmxrDr9bSzON5FlQd8zFrePMLaXyHQ0E6P35xzsI900
7qjLdjfqLH+8zukUWyJx9QsMCr9T60lWw0hqvl2LLYcuy1fo140I0+xSvUSkT/u4
yom0NyERibs+2WGYB1533/9drsUw76eqTo85bikQwMZvk4UA4QcNHVn7YOiRBxxq
z96qq+rdl0z4oAW49hNerqtB9KiNKwTyOgKKmOCIQc0YUm6WANyQpi4rQ0cIAAo8
i2B99Xt/tfDpzzJP/c3e5zvxRabmzf4R/Gb9yS906IdimCIRcVKK+ydp0OoMvNVg
b/3JvpfIKRxqi2tE7gtm9cAeObiPAJ8Zd7QBcNu+7m5Kc+6DnE74njwEq6Qb1xEt
GCbqBQT3JZ2pN+eQxlG+UyTYGsgxwSaQoS/Tlycw0HXcSU3JZuqszr6fggaJdZ1r
rng5vmNn1k/wN08TbQz1UA3D+y19CiPJ5ruaR/aE1nsdo4aPmwm1YomC4YnywiGD
W8KLK4CiA4tu/L8+AOVPdNIQXw3P6zvymksiDKqer8hoWDckvpkjSs4ejrDcyhOw
FPwfAVCUhYdgHMn+NHaPxxhunXNUF6xG47c36pefet48G5pKQytooW3iJtoHJirF
3G4aRd4TFIk6Sj3A1qxgvJEIyHw0wySlIXJ9HjKkHCqoTkBN9C/DfGHB9Nd4b2oH
CBHCwoUU6ifW+rTOu4AZIpeML8FgcjWUqA8vIZu0DvKNaVS2LboaOkEhfh1XKHc7
p4pgO7nqWl7D544a8/n+Uz8PBfxUlBnRXx/Gq/YvKLHl+vL0ftWkX3CMfTrBn1yT
nw8SDNtV0Cx79j0TwcuMbVZX78kaWhwS19MmsKFErxCRvPMJxT4quq94R1r/77vY
6LzDj4cO+5pdGb6yPFRAQXv9rzA3WcEgMhfC5MJZCISpUH8x+tx3+xWoUFiMZogj
/TjaMJ/F6p15tmiSqSgToU1FKfsGTWX3NEqKbGSItWcfzN7YYtgWOTtJZFLMbkkx
un9uxOF2b7Lf4709VKlSiQguXZLHfBdpiIVI3LYbEoDhPL9Ql9ZldT+7etXK4Psa
Ukb7sBWf33VS/bijp8drURjmUKVQmAf+5MNYttv0alKc2tMaM/rG89myB/pZVsj9
A8RuvVSbRREIezsHlitGCoWIZ+HJhWeO62X9Gd1uXdQ+xckiP42PPlqr2RK4o+g8
EQjDuV6gFMWLj5xixl1KhwpCudO0MKQZpFKSYaOd0s2wwrzd5gnCmGj4SFuPtNjj
4J5zxRN0yUcT6zRmDzBh3fmFlxjkiQ+ybkQ6WoyDSGSYVBh8B5LaTcqkbRNh/le2
fe+gRyBziYuzBaVC7xtcNxm00VgC6eU5i2J3sMRi6SK/zN6/L+BW281eflCmKgLi
u0I3u+yzA1XNN9neif7EDHgRl/oo1apzyQL0p6cznj35bIi6dUXGebOE/cYkssGq
KUI0wxbjHT1qZgRxtwx05DxjmA6e1aYMxe0GzQQ5V2SI8DR4ucicUHm9bT/vI8WX
kQcRTLAIu3wnVNE7iDA1RNWkRt3Y67e9Ip0POQ3KRWejcmzLZOqKrEB2GIti4pkH
iOXbwtyFBxWdOZTV7DPC3vbWxP0N1QjjPtLE7vJQyBbmeY+6f5UjWY+G8s3bQdan
aSsAW8CxagxXdoeC/bJ5Vi0TGHjpKAuRmc1WkrTwWXgI4z4g0Z1IOS6LD3tHMGC+
GpZqsDgaUWUOZyTh2YWmhm/6GOAMnup7IYxqdz4Ohos7yZERwEK2YwPJ0j6uV5zF
MzytwF8liEGRhrLR6i3Fx+Lf4ub5YOQvRylsEH0hkBk11fw9c9yW2ncoVDQFcRM7
aWE/bb3NzHQgyVBNJLLc2ZptcCktSsQNMuUwpw3hbELR6LnLHja1g/rQGbJpRNcf
v6fnr8HhhSc6gaBIypSulsUDDybpP0cW2ZZaBhz4sMNXu49nPqSMV0S7eMGuZTYO
Te6Zq+8z4iU4S1XzKOmuHLeXl+PJtOsy+tfLI9aJvgi95aRF7LdS2OgF1B2RfrbD
Iv1gaHOsOLbrkwJogIl8iGgmTDxAyPARtT3G6ShVCSDm5+jH64PhcCe4sPMfm4n1
JpZQtcdkRDD1Ruq9OzWl1/2KYZ5fcbVcMs3JBhFffR77tGYK/4T8bmvCQyImepca
j+p/eVd/Y01NSdpFTnJy4+dKoTHVmR450Zni5tO5RFNLfxfDcVtT3+GRACuAM4Q6
F7pOuBpU8Q3XcStn2158iWlbg+W2MZvDNSBIb0O9FcPGOC2ZHZarjlQZn6JnO2We
UCs1qZIGB9c2cCt1KUZxiuU3T6bmtqlQ1YByt1kmidOXmRcyrV8UdNZSF8pfPxTM
9AyAWE7UzfzW+8GJ5s59WZAb9RXstZ04LodWOY2YgfM2gerCw3IYCbP8EXzSMcAc
fWcfbMCrJbOHXYBcdL/67ijNvMv4MlpQCmdBfgHpvqhrqchIAcbhtofnZRGCEYWK
YvC6YPr4r36ysaAltcpE8sDmJUGS5UsAlzCNkyzDqNmYSVfVSjJTc9U4Fmy01D7C
vO+Zh1tAx0rYp1jKRQA4UL+5qr1Nrnr79FVd5Fq8NAAflCgYG4Wv4VqSl3cBlt6b
auPoAR/NiOz6cePyie49p3jlXeWmB8KOHrYeuszDX20rKU7FJLKWXjgOPmbLX8Zr
PaGLf79BKfIL6PLZcExa3hTyNPGNwRznOJEoXLp0LLGjKzqnFnNZK9LJ0jRG0vZ3
Tr5lfBaumGiH3AKazGup0Veg+ybMKdYVBU25EEOSL+s8WH11crOtrec8es0SuJiW
oNIQALv+9p5/Ef4fJipHntXRH+CjC72HmGQ/fjuNh6P1FF759HS9tiAp32WOssqf
w/JxT79QRini0JZOaUpX28HlsEP+rzh7dU12AL5eDu15YDBRrRvnpH7Eisvj9Gen
Ds/ZGvueXbgbZ2jgIp62hexbRHzQTxAgd2+St8gKPEzJHuLyaN5EBnlZktLP6YMp
2n06GmtP9mRJhh42Og8btZ2lv1aTN+4wZPnK6AH6t04LYpNKzCaIwqREWCV9KYlq
2Bpqzt+6upYIeeMhF2GvHO9QKZySMroTlJvsjTiq4SAAY/SYqmCPDRXEpNNnng99
SfYFwedffgzgtho0fMKTATIWau+oVYhe0h/WlcvLvVDlwWrRwyvp0QAHqUe+S2Ue
pUY0//3FBu/mYHvrhhSeevpqLVADn6dkCpzmPHayqamSdnW2oEsvLO1Nt+hjYLIk
dT4g/gXXR+PLrvLkt7fkar+8xoefsLZ0IUsRqibNz/ZYo8YejCV2Ku9+4pBuR+Ol
1T21ARhm2gHoMYnfF1XE3RtSyL3pkC4eXLIVcE6u3+p6efZ/xzKvU8e+tRbLlXD1
p+/UsF5r9pDchU7GuFmcrhzAh4GRLsKN2SMV9G3x1qedSfwCXQ7CrWPDKpEkKkaC
6A40EBM2u95CMLnIcptBVVxa4hofRIq3B7cFi2oa62w6jdPudY+iIC/sjSIABeGi
E5JYut3xZBSgupg7bo9odci+gUiLc1eZIFi1TM4R9JeTUMc1ynG7i9/YBHpHZX1q
qOJOANbJysgaldB3FPzBJ8Czah9vSOPxItnilfU72f+bINXXkjzFPszYktyjAPDU
0W46mnRqHES8DQdvKJdQ2KNaR1lfhIZNlUD4XWg3chjiZaiRFCCR2wIPAUqeNEUg
KkqsJYlxiMxAVeo2r13dIZFdjLEGqGgOWcjQI+SUuM9Py3Ae1b2XOWD2IlhIXK+z
CH9gtBwrsze5rcTl/a2BFfyFaGb6F3jgha1ZCEsQwxb8WvY/BcYdvlyGGwzian+E
zPH7soAUEa25W7quE/foeZS4iTEPjMtpL1Dxar9nax/yFFjAL+9LuWO7RnPjh3EE
CFVmCyBKaDGx5cFcXiOzfQyWo+FxdtWNhh363EhrzZIkgoI++CASRZkDMyFdzvAr
kmgKcejsJ1YiN0AujNKiwb4WO875sskXl99S8NrPHcHRxafVZVf5WZ0cjwUQIqsC
C72csoFkStw2OmO5br6fje4+Qsc4nx7A1ssthBz3i33bbqr8LNUFeMyDVNkV3BNa
KqE6ZJxHl4KotUqzQDr5iw9s+GcBPqfuSG0wR2GPmlUlFn9wvEi5Prb9KhjDWJRB
jlt6sdy5lknn4GU9uEa/lgi4Y8qcc42MEcRNYY8KIBZZ+DUJbRQoTswKAV3eBabF
9Pcaw+Ji4Prpd3mVEZ050hG7iXD4TM5aNSBcvSu8eYP+fQxuPOAeCuQjtbWqth0v
2GXOPY/UyBuDXZgI51bvLpbBsw3QK3Ro/HOttP69JBBTeTrlrsUrgrmlkDcTwKKU
q4FgPr1BsLjB6nku8gaOpAUUoKVNXyG+BBGLWOAtiVIvm0assF169rjh4sTqAuCZ
JK+Fv44VzAoRdUOLFLUiqJDt8iRmsN9T0cbr7Vqgy1TBvN8wLuxMx+2neY9M1MXM
MFGjogooG2js22nNiqFQQ1ZJOg1Xp1W5T0Yooa4BKwaA9mLOiZNd8fDjpfmZA575
QuYZ1zPsWELbu9EzlwhmIep5Zzic/+joVmRniie2NCWv28TI8WkraC/3rA9augXl
S/n1oP4M0yRkjLgUC8zG4K1HRx6mHFNq3GyPTU+Cce064zyjBKIBXCLqzvEszH8b
HrsfzUuxzxHZULlHrKivcnrXNfpvL/8YhDbaolTSiBbxZNQf2El2U746Dsl7GfWI
nGhohBFhGkpjqzSylLzSADyVu1K4zxObHNCIiTZ0WVqWuQoZnwyHBGvI7eull2Ma
18lygRbozPbxvFAfkO1qzAE3EGBL02EER67m72mZInWpLpa2vXYwsAqZXCUejZ8W
Y7iq/RV5VAuAUqxeFEHO9Q7Rdt5YMg+MYggcHu57z08cglIRB9foobOn+ANKOETm
4nTZlB0y5GpB4ZuES7jDlEf0vJPXdUUhD7eUVEBDPYO6c0jSIVocAk0tUeLz9HCV
r3LSoTD9/ZPP822MS932bDdQzHdDNSHvZddje8OEAHyVvsEnzRl4KBXT7VoDXXJx
jQ9Zzup7gdoBTkZXFC5DSH/mPWWs7TB9YkJNYRzqzepEIOxdw0DHmxcxjmm5SD+B
7ze38TJ7NP4nMunUd020dY5wR8zs0ojExNLD8adUA7WYW7FndvlprhfXvyd9mtTD
P6jbIvvm5QbH0aM3xggIJTJ8Rw0l8xybldspowe7QCw26sZvEGbwUFUayyvFtEwT
GW8jvEnmZmUA0dVJkBOIuzmTCx7FniPg9Y9xP7EPXHUYeVDRUaSo+mFb2ajb/aiv
4NEcOCAcGN4v/kIjFyY71fjFnGntSwJqs/k5OTSa6BdrcnppzN+Wb5vdF2xjrGEP
d1yXvOoZSHeI1cqJBaB+TMjHL7GoNrN57lFhbpyccMdFzgHLX7i7U/LutzvTCDeD
/TuswoXCuaZIxZbx9bsV37NEBkJtOKKzAbGyWcgUeatF5MB3jsh1ldW9yXdtA1E/
+83fG775zuHgopXja377iQbcU0o+qMnI1PYHyQMRNromh470ZXa0VXDat9QxzDlM
cKeFJ77gALgWaqRggwjq+PZtxkkXu3RPYrF/Y3piHD4fhtuN238R9HkGlGvAMmGS
0xEuxDIbuvbJ0E7IfxJlfqsdRQgk7UmMjc2ycGskdNtHWofNS2+mU38ZAviqpwIM
507E7fLaMjRYdFqVENAXztgIuALKPuruE1xWK4cz8FTr7ztSr97Sjj/ufmPBfTLf
0EuSHbEM/Of99HTbpRkVzz7w0NwLZKNtCTjztQxg+0ZkYJcDDc015K3lI5MuDdAx
8R8vZ9SwKzR7LMaEQ0p1d5uCSWFVKS/B2+tCaPgFsmPnUCcaSCC5bSUTr5jHBHTt
wpjHWNclaWxysoi/pPskU1gY1P8ieJT6plmRuBj8vqablPVsst4Ukfq5djKjV+Zf
yhWC0Kkfn+WBdr4b5UMrIlkZsvA043/l0nwjC61/95o+ZefPDLje5lkLLeInDdlj
t4+prGjoDI2sL8qZrN2Glpox3qcu/F8uNPZg46261hygzSUob1fT7SBVq0OLz+Bl
3nku5U2nMBcm5Di3w5scoHTBTny0/qTVNlQQo4kSrxRN69/J35z1IV3+mOC/Xhcf
AQ5lrzzq9D++Zhk23d23/xDSK38eroxJK/J2o5sPqTqaRjl301dTeBBfhbIiAaUa
zzsHce9M45Z/F9T3PdAKf4XsLNJ8H6zl+ACExgchVxbknTZ1rOryXqNk+QPU7xwS
TKrCi/8/Lg5jkYQxqBQkufbRhtavcdzlKNu+1vyqg4lzbTML9EFfuT/Yte4L6JnZ
xwjNPToepDe8M80O4l6zNM6EivzAqjwirjYV9rk/BpnAOeCvmIcZx7ntxT0+9K+0
cAcSY+/rbNlUd/tI2mHv0mRVqHAB1F8BGBbeLRXadbUZ6PY3EwypshS4/XPYfWbB
El5xERBQWxwpNorBWIpbzHgq7ScKlRSkbAThEYbSou1rGsZwSaqmtOHFOCtLWLoQ
7pFhaHLKz3V7IB3IA2mkdKrsFrhNGt7qvrBIGG0XmQu4MkJuLziQsa9R8gPrQJ6f
X2FGWLJ+e8HWzflFV1dFb9EizkB+NIZKU67hkvw3KA5ka9e1YoDcERh6rsLLv0d1
gTasQD6RVTVHK9FGdheJPlzYvg29xzJI1JHWy2/SrQ16m8UYkHtkrh0erv+tQcr1
H27Db9vTc0X6sxjufa37BuCRBZoRjx4YOMyXuudHwilNJsqzjbmEgNAlhqJC9ciy
l30G8v168Hm72QJYISklnw75hdjxhjbQdQ8q8xMmCkhHElymOw+cwFd0TMji6Fmq
W84wzwq7mJL2Zv8aKXmao3kcBko8budRh+FibTkW8SftkCtVLoFpx+vPeNYHnWsR
0sFAM9aUVmg1ag/0vwKkRpJk0A7vlXEEkcU5ifzZUQX48Ju9hHwAV9wqKFp7Wm/p
vv35ZGF7JClYDvWYlbYenx4Gd1LAEVfG6EsaB+8mCE81a/tXKFk6UTcL0V60aSC2
c5GB/+e/+9b9H5xDmGCKq/oD/s6WkOFAq6uZy6hzmwLNt+PZE5amoDJckAaumurf
SkNH6GqBBXZQ3WNdaK7lBse+ll4ET8ZLJ5+5IxCx2mdcMf9cPba2XdUm8O+kLh6G
jr00xHSU+q4jrOjP8pMSSKaeZpq1BJ0jK7Il39AnnCAo8q8iJtM0psafEVX3g+SI
QuL3ofm/2Z6j+uoJIm6jbpGwiMty0dYs8Z0rm/yguA59+QrqLWnz/GlKEPkNdkZt
IfzSWNqsBo94H0pQm4rya+4MT98/5CqlJZvXnDuHoosKLW8atCYbVljaejsE0jU8
4KIdVdFXc7uZjs0KK8pL5dkuMqo1qMU7WcrmvhJI3IV77I+r42EsGPlF0gyos5/l
+8iu5UgFTqS3ro+DSD96/XhURad+aLMyGx07yUa0oFNO1PNxbETn7LChnj1Lk+Jr
UUUhHsBl+RggQfZnRhBHmllQxDlxpv7UIwBx9IoCy4nzzl7OZAY1X1ck4uzoO7e+
oe+G1eLnl8nNTtz2nqikWbQYUho83NEfywqP16M/UhdbpkNxfYlogMnqJOroN8kE
kRRyCsq/WQ6dHkb1U6nSt0860FiNGleyozax2ZtOmrNl2fL7uFvK/6lt2Fhb9T3C
FTKof/ziLHotcYME6x/KmGokqD5MugRY4Tjh+/zk5SIepNNRRTtyBtNFHocXX8nH
+7ZWAMZ3iEqiYogf9NyGESUQVAvw3Iz/cAWSLkt1tqTK9lMwWra0SyaUGbVjbtjL
/zE6U/qNnw/9yd8Ytw/1D/+0n35Hr/UuFai3OA1l8+ySEcsd1rab9Hk4tKl8MW8O
kgRDvCvGEEjj/aQGhMJmBtZPzaeltmE1AY42xACe5qEQUMDn4bQKm2+e8bvt8faV
K11d0Ewzq45erSQc+iLz3rrUQyAkKmdQmIMAMD8dPw+fGAD2GYSyt746RUiQ4MMx
CU5g9vMXD7JHwJnGJxMh9SqxqKs3zHgyyCylSNPUIIWIVE7THTEfbomP74NaMEpK
IaLIF546Qd1c2NQVAsuQXGQXAQI981MLUEYL0kEI/0j4fMMKZXpQO2in4/mPHQVM
Ab1tRz3bdaL3d5mFnm/gt3AwaQDSTrPLxstihLIAfPXB/bCcVaEa5DZ56ioxE6sD
6qwWPoADiL6YglQrb9hGzPKrQvuL/cj0SsyZ5R8xGDSgiZtyTFPwYGduGtUDOzei
BUrZBIZyHcWvYOFRz1apRBYl+ZeMDvjRkca5qwSIYvjP+Ud6XX6D3/JmQDD334xA
gk3Cs18WTHsnloZ8+moRmy4ix5NFbPcMGe3VY7U6EuCePRuUxVQ1imhT7+6bMN1t
Z/lj/fjNJVA1xjRPky7UMe1ucY7xBG8+G+OyqHUrn4dLWSQPOVV4aCd+yqBIJgy4
VlFBofWWQmeRUek0a0BmqOmYHd23G9mkHcqGlSzib4t/7pgaawguLv2DC5zKvW+p
Y0u+hPsYLmVyGWWpHZLPpeSOMdYdeJxYdWL1QwcBq/49Ih/kIr8tILhrLxOpTdjI
9AFPPhBaKKBrTXxgxYYSd60nFuWkIXSWo00nloIa4Z1itIrgFc6NTqeBazvM0eSM
TNyDX+ax4nWmFY8SMx3YDVgOdJ955ZTqdsX0ZlhPb0jIDx0LoZvjdB9HMVtQt2ub
vWWSE2prBINnzgw1giQsj3b+89BI1od5kjPvmBM4tIi5kESqeba9GQmTSuJn4E0T
KUGWaTY/X3r2OMYlRoLY0RoMrcLllX+oEi2g78rBskzp9z0Qxker+OO9avAI32ce
+BE7ZMpmcR5g5CYHYK1DTERQYbQtD/I/Io1WGJ/17VdF0f6is6VJ0c2Y3AV9Xz9d
JetZ3Riyd5L0hQOqe6bqeesmgua2cosTuORvc9AsepdWPRHk++d6TRNbqPXFGSrT
IdS7O0IGNiMWbYlB1axgLh4agjRhBNQQs7t2eWEMAoniKw6TF87syCsSQnp5hCY4
adogC08aa/BLpn9n5ZB+zXYbWjUwivIzJiEFVGG5nvMyD72ghnQt1MRplBd8IKVu
fepFfZ4AaLhzF4p0ir8rksTf0I3PNVVoOoJ8hXa4jwJxKMhzvk+MnFxn3PPu8g0d
lKmSZJVledPC73xpRMvFnRNHZwiiYpP9OuM44ng2/7L68Lkjf3iEUFxMy0dVIl0y
BrWnZQf/qBps0gmE7RO6eo09DRV90PPvIuxkcMbnLvD1C/Lb1wIkj5VGH/8tb0Dj
w/fkgzC0V6cyiXLD8Ji7B5vQ2uskUKR6q9nxyyp2Zx7DbwYfcU3UBDiZxdNOBarg
zaDhoBTwtNOOxO2WTI76FQZQnzzXOrjuJ1qoMOn/LcOOru8ePSJgVULw2kn/MAPg
gJca7diFUzhsFNmfmaTYuKnh72AThRpgkamxxKtEXjO0+mUng9zbUFa8+LFnTnBL
m2CdjKQTQPLzp+21xMF44N0IKguCzgkj1M7DgqRKNHjLlkSaRbcoFY6JBch/lII1
GYdds1W5zTLdEcRe/wwMrZJo2XRZjYwp1GlTZVmtvfyDfeltnCHZCXzzbPTxNw++
aqsYc5b4c1biIUzC/Wm11Fh7dTFZ+SO7H30J0Sis/3AmDGAl20Ctl1padebB57aK
HgByW8af7b0mLcYln++Yr4CaZ0c9AywhyclSHQl661lQ6+//98yp3ESGcSmdYYzd
S8yeedMi2fZhYXxCyqh3bFrup0tIkWGqU+BmuRzb9Z0xfIyXL+woAkXRPyzRzU/M
s2u53y/VGantPeCHgiiFoK6q/vCRJ92iRH9PtE/+CaBnCSa5S/NYfbPFrne7gyNc
u0mjczPyYFDi5cn1I1Odl3lFnYgd6PqWTfU4fhCB2Gu7f2j3DFJDtjv5B54PgvXF
UEr1Z830kwwsueI1J1wBUoFtbWYXRdPozMsmanbDDZnDbOhKsM6++hPe35kNAhGp
eh8wN8MaBFCbnBH+wyfDg+FhG33tj2pyoNZfqLUuK8A/eg8b83go6roDX+BPwupp
NTkPCvo9x5/K5X4u1gEn9dvpB0kycGVrTxIrTwKWZo1SjX0+NVjBYnwVxi2VP5K7
dSc6Q56fiBIaCH6hT//S/gVeLHp8NgNXhqWkacM9vT0/OZzyZdhxXT0Y7eZ5QhJ6
ABVXeU/Bn+eU1WJqtyzlnDF5xPzJAGSMoZ/0nFq/VzpPLaAJrqwoQX2akHFDLHGI
vXKqYldk1gwFVaDk4xUO+/dQ54X75q3tkFEJNTEHqyKRYxToRSN2ZWdh3NMkFG8W
aCUm/qdauLGRn/sNCdTbWXJoF7zmWoFgQzgvCTaw4Y+3xDmrwlgjBvlATJB8NAXj
Q6Jrk/FVTQ8Q8P1SjRPbM/u6Pr1CLb0yjQA+RR38cJyhMgUhPL8B7Bwj50ctJKjI
991MppSxVItCIkPuj+43Tvw7lw/fyvezHAms7tPMI/xRpB3n9xGcghskN+khRG0l
F63YQQClnD7lgoBeRk6ltl0WUdCQ1SPhPxV98P36oE9cdpHpaDzpswrtoVqdRWQp
eU94TaLpKYgpp99qA5t7NB+hKNBjCanJ9H2V2GeE3KgSWQt8rsuOZgF1b9xNblnu
1gzAwsSxJgHiMIxpG/5Il1ytgAywYQ9SdbU2KdegRsSFYkOMPT2xdOAXmOzFbxND
6MKzN7BH1Em8jjZczojIg7kgHOWII6dhnzveIfuaBjZEZZYHKPSByq2FC46i1SNB
Gt3rd4A9OySq6KJD+st5sreD80Lu43P5by0n9dbdk1+rog5PTtmpjmR1Tqm228Li
Lc8an9S5xSzVETcjF3u1EsiFuKxmp71KcaCNNC9tOpWeRxMtFgqJBbB2E10CQiH0
2mhGENZ9I3Rg/uMHM3jKce1hFCSC4luLolTV9XKvf+xRdc3bzBK/aFTtYNwXm1nu
qjzcBf2ipBe5nnkNwa6lOXGR0kOd2nlesT5gr+F59b+LairGmEFHjNql00oCitEM
gAECStoCUZWr0mFUSuXjvKevXOZG40iJmf/e5RRxph5wTEmF35+7LgsqWRQrLSDE
9MVV/ORWAWlOJF2E+Z4UyFaUAXxc1TwUlSDfjRobR0SoP9d0fJix597Wn+AL5847
sr2rY1BzdS51MF9emNf/uVRTkFVTJJsIpwanr2hzmRcBBWCj8db+5gOEjmc4Ywfz
gdUCoIKooe987IJkrmTDjWgRTf2S/SBvARwPh3qSkiYCJc3lIUaYmhEAxOxJ8gQA
UcV3/VO8wSkTsLsOqQ2lcCX3qJPGPp9k779cvLRtaLyeB91KE+kaWlf/u+8mY9G5
BJDkJs04K4MOLdxA09gBjET6Q2rr9gd5yBxq0KFVnpFcGIuonhoR+3aJnqk2yl4u
U/zgh+0/K66VbYcjzayXF8n2cjVzge7RGA664PSEmOMcZ/TVAzpBjD8FfHANctU3
QuiFXMyIsbj+QQ1dF2aDlNXQf9n+CYzPkLJLqPDLiB0nuZqXfBswBh56wCBAcIeh
5Z/kCmEvY5FiZkY2W/wRu+c1U+x+pXA3248KlzUW39+s4YS4Od3YuhQL+01x0gG1
Cd2vdScjBYHbZgTOPd14lXa6LvSGRn1ViEgKPieAQDkP9HXgECS9uhfKbcLsr6Vg
YyK+iMrD7pQbUPtKRcicrBA2ya1z+NCgwcEqd0twvUMb45pgNoe3JYdn8gvp7VQ3
Gj51U9Rtn4W7Wf/N96WW8/hGCKbvsvUjiCNbVvYvXnC5GxES5iQqNu1FmZmfjw9u
hkZvZVjrg3st8Tba4zHmX4RV/BTKy/OhF3YGyewh2CZsvVbkHgKhHzYDwYYsYdnc
/wtlq5Qxj56uoI6pozTORlt4icVRv4u8mKi3n0Pi2Oxu4ar4yqHmtLIvs7hP5z6D
K7BYzGQ27JY9d0ICaSYd4LYIauqWx1oGRIDXdoRPGuAiWKa+EHJMYGdLXE39FGMk
G3x40/FOemMnuS5aHxghOyKfKkLs2Gupwh4l2hSm4fwUPzCzQ9N+XlajYf5FHblt
LR+m3/06wnceMmd3CUXDdk81aLoLc0B+QSNF/DxzpJqSyza74ErNoj0gfVmZ4PDC
zYTzIt3CHDX5EnbOj4ar4eAlXDYXC1imkyjCJCwXcdAH7FsTI9FBTqfVGHTOtW1x
yaOZDu2t9NaGn37fjrPzH5LwjBM1/mBNSG+CgW6ZIhxM9VhaROehvPSP/o7XFU4L
yjc+PjNDeMqyv3u+8dJ4C6QU3KAhZ1kKP+FA9qZoqgo+22SOvTyLijdBxcuYKB8r
L460fwNUYcMHlBS4gdbHnSOFnqiFwMdqeVnSG96AO6Ww8tsM7eKNrw5+Q6yGPwJb
U9J7XjjAV52hVVMQQKGxGboio5GWISUlbhpSAGZTZfDuxTXImFIQZljz9iM6lJH3
H3ovEacyUYRFODodjPEqEznUbx2530ks6RBwG1IIfndJyn86FBjqJDOQSlCsaGFq
HngiUTKM7i2Jr05gNM1yNpqU89lUrWTtlsV3rG36D9t2crllZ5Rm4D7uz4EjBH7F
cMg7cLz5TW9EmR9fY0PaHSlZvMGn+bQSSY1Z9Y4dVGh4s+enVtd/EcSrq/N8ZxXg
VQRqSmRftt2FPgtb2I98gectzYiM7dkYmKRGsL+x+QyJJeQZo87FqP+K9/N27luC
xd4LqFbSNGb5D9vsqUntL2Gx38S79wA0U8VKkdJhcANwiDx/bs648qbHeUWTSZaf
WsQf8wcTLwA9wkSuulzTHwrSUGsGeq/TM0V2iVlDRMlb9z3o/fLs+7YPh3nKfmgD
a1irESe8i/fm+wwol468iGDFp9RpTysspZehreYcfwjGo1hkqkMrGrjvNW3za77v
i+2Bdi2irBT6i3xoI4edZ12inmkQE0+JR6W/rCRw8j1KTEqe7ArLhOQwLzN8srv7
9TlJM8J7UZJh9H4azZxiUlBLeJF5GPvp0822tDFNNkDYEgSzrMIrdZC+7yxkdGTk
hNqtHVSTnOAh5nBEU97AazOZadGXdsAJ0AfTNz5D++vT/N66YJr18Qz6XL0/D1EU
v3SU8LPEX4ll1GYFJaj4ZXsdRwE/ryBTXCuHd5lQz9NqaqVKpDDo2vPrRaLU7Mpu
xQnj08yeNO8Ixzs8W2CxINPumgkYlts8Abm+KBclNPm/imLxGMxC1SVma/EpHvpq
MgssszG39MLOZz07OglG2on1EYPcC1qafzUIteKuEN4LZZaFHuRd7Fh5wIb4ptYa
OLk2M36wzRSjIkLZxm+NNazKHYekA3adBKrn/mg3bSOuCPBZEOzBVa1sYAHmnL1Z
H0uxXdBgSFyrlWCh3FbBl3i93QGuOKG4NoflqZWXRVZlLH3ecmb0nIl1e2STBCzJ
o52nGP9nO7d8qzCtpWSoznJXU9V/AWJHMLW4a1ilF3shYs3R/rM9gxlgV0nHSSKx
XC7vb01l/eqw7+uZg6oxrV80BsuFTSG4Bpx1CCDyxM0QA0yMVfyjMJiD6KmDl0Dd
0H/IPYfzIV9fImsZLl8YbPG+xEuYPCALNfplVPavMrO0IWloiKOcgn7zgtXrWWzS
Xsdmm/p9wcNhWZFzLY7VCUzVAT8aNb7YG5uN+d8VBlALOKeLbP2E72QXjMGB4ICU
qB33efcuVa1Vl9UMqutClXOz13QNsfGZiS+h0MvTzlBkkype3R3vI3q6P38imvml
ffI+BqQKrZxdSWWsXhSXCK11JmHNuWXNUBKkJgyTBQTR4xmIpmdSR8QsUzVQzGBt
CWacXNzxk3s3QL0xt3xYrpnyB6R0BldXBFI2d406AZ7ilrWTyKk+v8QMCc9Rj0NM
0UtxlNFkW7v4SGp0MEpTy+Zcw74FObPqkTN5kyr188Qk4Se7E9DJwtxYopL5WFZN
SNDCRJOgOpPUaVAgRqvZ5QX0AzF+RZsbLEEbTUWR9zYd7gUEo7jPmh7p8/9HKrZ7
JXTjm05FR5ATWo/GnRcJHRqgt5osSaTguGPQfa6RuExzs6Trgvb6G+lwXg6eKT/G
CnYQ2FYQeRncWd6hU1kfuvucHshT4Mf4kIckTb8WFos0/oUxTAVYZJES685oRZAa
5Rn5mrb1qJvU4o+VGJbSSsq8UjwPpCyyVkvlHckzWmt8VlT4SyQjKmoX/n0G2vt7
yIG3Plc1HCyNeOPW2dN7NAXNMChLezW7SHT359YC8Te9qoADDiMsAr6CZkGMHwpR
9ErGUBuwGOdaQ2qIkHx33Dx300aA5qFTy4lkxUY7t1HCYnKI1Kcnkb3RXRxymJkc
HtCuteyoZRlUlZ9qoDtsKiqcbI7KzrAMVEC8Hg4BfrZPB1tWSC/B5WF9nD0OWUmV
TC6wJ05fhq4ytbJksfmxcz+U+OslJAEAc2FZ9KGyXyWJtg7dUD+2WiuyyIJss67X
myMxJ7dwPxwxMObv4xWjWZwacLZjfOncmIsJMaZ7xlbUo4tZBofd87INhDvc9zZX
W9bHwn7e85/hKiVCMQytrNuPM9RRu3TOM2nqEEjFalX8N6tMC+NiRygICSE4Ohzl
AWpad23G5LDQIaafaXLHIWcUpwLD+rc/4Lk9qSqitVgzZI/a2Vg6nBB93/WYoL78
zy8Tl6LLVL28nsVVrwPuHAM4Rnqm5lxWHecyQnDUgFp2+c1+sO+DSXfWJEpkENBG
XQiNWb5iXGZAbrA+Wuha77el9oWNs0b6ZrTpkMsXw+ZPLuLvowLREbj90eI/NP1a
DyI/H/SnPyO4hc3dqsl8cFZ9HtrjgcZSmxfwcelLNiT0sxD93YxvhpFK+4XtnPhi
VMqJDjdxdo+TqPVKOZqzCX4k3u+CylQeMFoNHz3b6QJJDdz+EZwqF//71UF4mCJN
/Q8dWPmK5KKitOwpIbjJ3TyAEoain3i74lGOY4ZHvm35TnVnI0Sl7kOeISkAhVIB
ieCQkIzY52xniLXQArlItlghSg40M7valM1mnACDp52L5v+qNDHa54FX0D80KVUc
tYuYl5LyCaadXbkPvXCNkAx2qmoxSPDk1clG7ZMN0yWSGF4s0kfYn0OKzEjuzSnU
MSzd9CwJ8dH9nk2cpuGIGVhBFaHH7fMtFaaydxNdU3xiGzU7Yft4vMasjNNGRFEF
j5bUd2RVcDvWCglVqna9aFoalouA1+zdMv3p4nPeS26r0jcR0OLpAMs0EvfT4Dtu
xGa5bfF+ovleAAtCmdHBbxu37Gj0BUAG6kbUd+AnNNb3sx3SJgNDv8BjNuaC/Q8c
s1QkIwLT4qEGM9sf0/p6mGfpCmMi2JFnP0BW5seILLXUkIOweM+ZPr/IQT3DKxfm
Z2F2lq52VjtCntlpT+Dy6vK0+O1I7y4De3dH98+cHZrszAnet6fgCr7kIu79zxzg
rCcAOJBbyanSY08cJzF8flPvCShybogOSEJANx/VyVDbpK0PguImDiZbUi2xK2NR
NuegnUIcNT7AJkqqvLqEJKLvNjvdNOMHeLiT8q4JkQwoOvfed6Qn3WjK0/m3NgjJ
oyNnkW6IyVWA/3deaeCBvBXDOpWCq1gOq5eV9qrttklyU3xc0UB73d+I5VTM2Ex4
NTAmzgXy6BtoSdkFOxw/sLaPcRCrCRvPZ7RxhFTJLsFOIOP4QspD/OVDNCsxNAmt
H5x9ZlC4y0XSqnIiB9LHhFGPCR360rPhBW/kQXaqD6sR24dPhqK6buq48XAUv/gW
HAuQYjCYQhSGoalRoWISeGlwWR/kXMKE2WvCHHv5AxwEutgtydQC7qfeCaltolcs
AuN63U33mb5mBwpYs49rK3boLUxzUtRSOcqSnIPXbvZ+2MsfT6grIt3vQ4tBT4r6
bv+uYCziJngCB5nUuPUZfGUFZvi4k9wIP2XMqCdoKE29sliIgwVTLDWvOAYprcXf
d9fLnTLRYEYJS7vmKJgUBRhF697TC9bqH2wBIGNO6j9PobtxdJKciVrNQ6SMnQhT
29+6IVClcum0rtxd50mMIldAzdNSrdGAKRuj8w+Qj/Yd44kHue6HiC3k3XYCYnv+
73Mg9ZAwdcDRBhMIE3L472u42kU0W5iIBOciGGMFxbyNpxa+4W4HbA3UQSxr2XEG
mT5RU7s0ShavPeiNd3PHdTkr0Lm52B+BQht+80E40djcQxHNlXBm1KOMCai30rkM
KJgWHbo3FuPds3zJb/j+b7AWg4iEUfVPuspz/Y9qYNKfgy9MsCuJpOOyA8CFATBC
sRa1p115DfKK8T33oOn3i7RC4u12J3htmBLaQ5zNf5CcnZGJL9kjpRSqc0nE3NfX
hCINUS+wa/j66bwqGjloqDhDHDuVBOVpGBOWSt07RrFY5n2MOe4V3I/2T4OQGoUI
Iw3DvXkb+3E2/wb1NWkBlusgsL+18uL/APrWnngGor2oU0K6MENJlITgiCJmK0dK
2gbZiafIfHasTVOVNvqcxa+MFFwIfLLRVdkGLSUjeCOL8ksZ2AdTkKNMcf4ffrmF
PpT4O340UdritdljcZRV8+6a/nu7BJbDrFdcT090sD1+uZgD5yJxebS+p1bNfIft
EdE9XpoyzsjOvOuzVxgkjgWVVH+C4Z083ydo5pnQ81ldmvBAoDW7U30RxCkSzytc
IfpfSsDL9mHwnBnhkcp/jw/yAx5zwcbzUlTvyiPR3nOBi7Rb2rRXWgTZdu3arq1k
SW+Ins/OXdRGc6hL49RUjVr1HUPkvKuAkuajhSQ9ha2KGcW3tDy+b+4SaFOvEx31
yLgg8VQF9omch40TQTDVQlDUJfmngXmTwRXGcGk4SdPPefwOQ5CaSrbETy2c+wOv
aZ/7Btu05XUxv+2fJ+VgXwo1iGvyq7TG3IeakQ2OJ/lhPgUn2x3E9BVLMQymamGq
n3ldDGA3pEVUjM/w8N/Twu7vLLPmKKk+miV4jcJzIwXIOJjO/l419ZvoowL/qQNU
5zPbddaJjPrRlaPyC0AeGSNoSUpABwAAFTnasqZuaB2iCizacq8CugF6Rwe5pV8I
gbwU6JseDLVv90Y2+WXmlg7V8dNnIGKnwWl2ex4Jt5GqCK6sm+HB0+Fg2TDBGlOM
b1FTp113blhkmQz4HPxUTeu5vocj5mL4oKNpBfknKeypQlKzKyt6UwnwkdK7Moas
PboTHE/PxZniWF12CV3VhqKPxjb+771P/WtvncurNhxMZjKi1OIh1jBlhi2O144G
fkEl7YjhUZ+5tDvsLsydyvagbmpeWuQ0RN/Ty1t61LMptDiiChsA1mWh0RdNykoj
pdF2CTb6Tvqnmd/Wk05T7Qr1TKqrUC/CLIdyRAqAmj7ysMLJU+z+oxzJBSWLm+hq
JDj16GvU4d75bUYVLMc+TCV9HVENHpD1scF5herMTGGr0WO5uc07THjyn3WRkeo1
0HQGkrjmujuG7Bhx/01Bvxxc9BHruRUZYvKevJRpxwtRcAnoOFDmdGcYZrER7DvE
cLAZyxe468f+UljPdg0jFpe2k618GG8sP9A7/4z/Xg4rhqVJ5ThMsji8cwtLOLbf
FFRdHVteGjAhCoo0PykaZMA4DvGKdElETE8tGkK5GJ5uFC+8fsTnULxx2rjx4dHw
JNq9QjF2jg8DSgFTJDKraq7krgZcwGZMcSTkCC1l7I1xo2+HMsqmkX+xq/8AQ7Wj
/1kwe+eKysCQtA4rbgCG6aRanBZE7Pov9FAu7dAMOsnro6Q7xuqb6MAg0Vbg8x/e
iBSLBeE0ncw306Mhn6EC4KsiNlP0ePSTtkTv9F8TBbzCPCpB1p8jvfvhxfX057HP
dkcRj/WAl1ojVQeN3IGLxQhDh2HDA4idHCblXIGEiULh1sMKxjz6inJEsbAWZuOs
LAazSza6kOkj13gWPZ0VUWvJVDvAu0JM4QywNHMQk78nYkdk5XltqqDaS5UuvEPC
Sc1YJCRBRDC/J0BWIj8kqQkZJOOD6msoUM+xoz02FjJZ7dk4kL7Gtxh2kUd6+EAQ
IahkDmKNTLFhWl2IvX3wXMKcA/0HJ5rgRICqwu14/gI25u3Jv3Yl84vpsMfekJTF
/O2tBXpFQ5MLeuk1m9LXetf/+ndz9ImQNuVmN7lXGvBrJtmU4R5EUZgwSg+uLjHf
WjY7zrpAiy3neKYI7ScNIhcAeQweIWC3ZK4RbxQ6RYYjOyGZfmBTyp8E5hdN6kwa
1pngOC1QB5cR6IwkyH4K/udCXe4CvoymaEi3bkwq7z0Egll+kpB2R617HytqMOez
JlGkvKBX97npR9DX6LAh7HkOh/hgMMW+AIAja0QA0Jh8UrsRwaJHTW2rvFO3Owgu
MfiYPnLh0yLkAu0a5cnhD66GeJF9uPjpxto/LtTpmoo/oRm4ARDWiYOHjBMhJUQ6
D+YHpEFOztYuZK0TUvLPk5g8/x80MAtQDt4aUO0uy5nvQmAjC0uOqSO+4wt9+3Rp
Ln0i+H606WSbZMqcmYPPO2V9R/en36cyYejVzvPaZdyhQZdU3peY1DEiW1yzzt30
3VfGXtxmUD8hxyV6fEfAq/O1vLU+fEI4EZThtO50AqXc8+HyM4n35cMAkt1ojAmc
+osf6SCFlehEjBUaz5DuVb8UXG4nBhKtOxbhzBaBaRmOBTw5o0Ap9bruQTBUmRw7
dpYi9nhNKm5nMNPt7SOCQYB5TW24to1Bls96Jfl0iPB1BPusAV13kIQ2HQl9wYTY
uHqnM+KP2EWlOT9cvJUhLWgMAY82O6K/0IAPtgIDpSPxO3U10vYQScWJjcHB5uEU
ErIRGFKyC+O3x8JPStpTXnOUJjiq2mSejvWfyHihuKf+7FPK65BMrgUE9j2S+5iU
BlDW+dLxXtiK03cOnR53huiNaHWz/O0Auh3/KoFIx1I2wP3nat93o/o7SbKxGC8Q
K+bdTg08dMoBkxiin5/+/J9whZoFjh8vgWhh9DY0xPvC2cSbDsopYUCVKgKuih3D
tvdHD7/wUrsD1gndGS8BUMQgbXuDWzdTtTR0ixlh/elGv8/yl/1lohSYTKzdQE1b
DeJpR35XJhBswyj8HTEqaax1HohOvs8H/5gO48i0uxFi2DP09y36Yz+GI+8xSEr+
5LVrPivEdV/QZN37B3yQYU576iOsAlbF6FCbo8xn1czWNQgEDwQtbSF6E09dozak
qjK7my2cm4Ks0942H501F84N1MLq7SwNvQVk+o+ww1Wt1i/dDDAEQKhcSvAfPw2n
yGywzV2m1IP1PdYVp1uj+r3xkNsc8e7hd8k5wQsdmYKC5uFFw/SPoimrE3fhDtdu
mdsaqMCtNdrqTHiGTqNOMjCoeiSuwGgjgYNG775Z0k8PGrELu0iFQwoDPIbLNmVM
dfTA7aJS9JL19ZIV5YD1yIBVdamoNES6MJe6trw/7xX85Z9Wocuo+FG6yuKiwMps
QipspEl8z5XbAqJnExBxfd9UX0dUOFZKPK6WwHkrcCPDNRmyZ7NTy2RSJfZaBv80
Wiwn8J103XmRWt0Xu9gZmDJtvnrl4FKeGkNM6/FuNzTe4b31XWSSDEIAWEwwm23i
udal5ApnirGbqtwIxn8FoDtw5p7QT3EGS6SpJsXg932KP+N0xCALiycZDI1O77K2
Ro6WIacJIhMEwRHk5hU5ccloL6dOTQDmcsB7hBHonaAL+pwyI8jNUnO+GjKmhWn4
s1C7Tcvp5D5EIyUW30F3dxs42UeR27EhYZpq42JQbMbSr0GJ+1gEqBozBjOLow6t
WxRpVuX6cfCWhlVY4RlXcN2MAo1W7whhqniKWVZ+vXNGZKYGYIViMkgg2G/3S4FO
/UTO+2V7DdPOMs9C5SCRPb/7DyoWoeMVmCG4+3dcmDh4Ii0ShKF3xMd3SJG0js8U
OnnPwZKYch+S1NpU2Khtpm96mdrv0q4pmsN6e56J+DMS7fVD3kZPOwhQFY/aaMtg
AgjvVgrRMSiUB8ryizS2XJYTfmEuHprRLC2luXl2b3GbdMZPRRMNtdyIv4ERUu4/
VZ3GtJFXoYbwaMFaxcydNcrUw69TBAkXwRE2oHT1HhxPCX4vfgmCGhugXPp+v3nl
nhU9swFialiAHS4IA9y0OMEk8SCG4OTmmwu5vc50atYNLW8/M1Fr2qUlqcEB5GZd
8EQPynvjRO+hOKC4VBP/de6Vb2sUeJ0r+r0O05C6kOjUHlcUqN7COtJRyrEXhybl
tXMW9TZ6EU0QN5p1tZqJZxL8EXIiJfV7CZg/146YIJTdGluDsLGE1mkxksP8z9Vp
oF5Cy7Q6ZNK/lv6DQjLA8kQGASnsApezrqKDvYYRTzmjljN8jNUmDK4etpeJvXcv
y9TjHHCr92EVGbseTsMMolVL3TtAsH2V7zbYL6qGQCv+QN0QynP8zGtK4TC84vdi
BhB5Yz49bdSJoHyoR3LWLJNsazbpM17yvgVpq42sHq3B8hjZB7EFaEJyCJYcyJjk
GnDgz6Dmwv4kuveMBtP7Z7h+0dNr3oKWBNTT7dZM8zmYe5XepClTl5sAEVlgtuj8
oUSImloRIbNfuVSs9Dg/jtjWPR1gYhAuGJfK3UiTPD0kSQzJLqSYjAWJQPtYNgwM
X7ca02eOeIGprZMxo5z84h2ETokWkDVERfrxaYYcGyd6C5BTVCgYZP0SgeirHpt4
UCjsMv+I+FMpT0Tnn2LAbQ7Zp36TItO9nZoo8mWtTZ2sm746aLFrwKpe8dtI/U/Q
6V9zJka0aOlnVIDqMEHTqu8zwzR91c4pLSAtbAYQwmx/kCPVQ+uOeNOGc9rJsRhh
8/3zabF7oOn1SAfyj5hsNLRfQgB/r2Q0tFPozI5gPbO60RuBjwTkxnShmmzJWS3e
0p4IVX/s6GNHFrI1lWUiz5wFCM8Tb6bYCz9qMiFAhstk9NM+Wq+wLAZS65BMGnhF
AFNsBifYaOO/XHjUxaYS8W2tdqZ+A+LjA4an+t1DhxPQZqsLDhTPc1uHFegcOdG7
s/1RPWvdyY9GMsm0HtVxCzj79VjlRCCeIMN2yGLXX+cAdoryQLcpCY75RySuekhB
7UTOXILTfISCopkrFzQYNJmqkCxbnnp5jiQ8Ol2n3LKmvXFHUXA30ZWg+PrlECWc
+a+Fbq1GdcHTPKGUaZMQHU61A0LKeueDFh/c7ViLSIFdVl0u53dP98pF9uxBbZOE
jhFGxb2JKlvlIrbdxrag+tP1uDrrb75N4/k/GvQ5OscTcZ+IZl/nKYMbeXwHtvMP
tB47H1g9sEErjCCIN+ME4plU0C1UrUT+KB3sDJd4fX8C0tutSUuGCmhOR8kTnDhY
azarvVaXzKL7Lo1AV8Fzerb7dD791BS3/TxgXWa0s/Wyg0MObRHmrh0hxMTOwnpy
nuCBWte/whZf8grBYvxEKXCmZpxZYGckLOlkG6CZYaHxam6s86PJXVr1no7jElnT
lZ7FV5CMJGF3+SBcN+qUBiT4ETPr4EvOBHOUB1qBx/33+O1mdjUIfnhxq2SNW2mM
wG4Yownz12io7nTvg2fhoyf3nmdvM3Al3xG/qVeUEjOWnKuuW+lpvdXIGx0qmS6K
EYQRLin4qPwlzln2uo3SVLPvSPFxb7nplXK5eiJNn3YzTeKrz5ptQTd/o0mwBtF2
iDEwuBTUaZurd/wIBrOm5YDs2AQ2HqTMbMtVDe43roqMO/owKmkPexTu2Mc+wcyq
nnlFEskaRl3dsvMALn05tSvRRmqmLYrhvyrMqsrf10U0+8A7dQIMXnW/jCrPoQsP
w8io/wO12UrYSPRHjWxbUodPoNFvZMQ6cX5MXqYsaPPQN8DGAMVR34M+04exMDws
GTXmQFQKWTTnZhq+P7c+aRR79IczM4n9leGPC78vNhrWovdeAF4J62EEDWKRzmrR
fLh57V4YCEf9rmfnsxM0kOx8uxCNrY2ru5fEbtFNw4jmLz1Y0ecbmlhPFbaKRQOR
AA64pNWDTchgk2/QbFr93/6gTvUtzY/Y4r8kPDBg5Ga71/ilEB7wJPNHgC0KYba6
37lMpIArZ2J+jAxX8lUKME+qnyURq6tPQEcYJjIzRAUK+vLwRJNrQz6Ig2pEAq08
5j+wCPTG2heer4OeMdOjvvI6vJTi3g48FjMEKiWS6dUXj+V0VzZivZPLrXxMGgUx
Cq/6CcvwXhLY2ozw/CocB7vMpYMgOt5ajLtQqsn9cTIblRdyjWi+AjcIC3oxB+Ks
LOYGrQGZvxN0ORCU0HvWrcIMICplNfcxuDeYi1z/oLwydEiGhUkJPyfu6sicqUqs
aZ1Qd3M/D/VaVKUTDL/a81ykTTZl7Vrk6oAsp5seeqUYtZMTI6ZUE2+eeIZJfpkx
H2qf9Wz0I8Aqf+egP9Bfvmb3U9j5cVYXU/f/hADeOtnB3Xejrh1bn324iLY+h3c1
q2pTIy2wic3ltYdaJGXtUzt4rSomVt4ChLnZhD2ZodLSwLPWdmsmoDnomyA+qxN2
Yp3333qIKN8pvWZ8h44jFQshCsaqc0K9hSSuUo/r+Uo5vIkCtnvJK//f1iJDURpP
p4ZW93C/XNbvulcRUkRyG3R6nsNbCCrTWovuApKOyCvVA3+ksOR7br7UdUjabNLH
iJtrVIX3bj/w5ArLCSBOKYyapGQaBLdxFA9k2AmdPpjFZn7sTKm0f0SEWfRQqOTD
Lix8v8yTadXkCzey+kN7guuz2XUzOKHg1nyPF5LrXVfQgkb44lvY1TT01CAs/Ho8
V/S2B9A2+7+P+DkIkA8fmZYL3KK0glTLqDXilFHLICAi7RxqLAwZ72GY7asylu6T
W57UurYyRG5eKTtqDPlOWQl517HwhSn16UkJyVoLgXXfDUtF0aVMhLYLbgCbIlV9
QJzhV/Z6JW09Iuyo91IvbgjvqhUdUH/8F2pWJz0kogBJEmjXMgBI0MVDnj3BdPBH
A8nRY+XykZMijqo86cC5iN5E9pa5BEtVqVavX5jPHla2JyEYMlPkvqWmNWtq1HFt
nR5SElW4ai790iUfbup9AZGWbay3CIB3ZGt+s+CXC7rvOhGBeepmMCZoimLZleYF
Y6ngnus6Q3Fk9eNmNlE/aEGhNPhqRxO2IoAN8l1Pr2ZCNH8V/vAFcGlw4VOTWQRP
mcMYMe55fzCE1l6luBVuj6XU5lFrIcblqU0srrphA5eGUybt5UA5FdOypKVkGrPO
dXR1Gqxk9PyYIJDXCRd5zTYYXbv/dpIQ+hjYvYVZyMSSzP8asvWgC5s+N6Hqki1B
4/w1/lyF01W/+NnJ7QZuGRmu/ioY+Nn7pHGzTdwnlVtv90r6dKgaI2GMn6c5Tob4
v59UCueZwosEJORCrLtFLkPUcQSvMxhvjEHUffyFMonDTEs+seTLTUFs+n9LVLgV
GyC9+xIM/hZ2x6ShvLMxy619pJn30QmAHzFNt0RvL5GaTYhLqtv+ENsJnc0whw+R
pYGpDyNmwHd2VXyudyK3qJPtwheAvCulbfAiEoHMNZrMyR93vH2yK+DClfoodgVv
drvPWv3YYXkaS7waKlB+71PuVzbFOLcZI4KK5pEkor4beRjJbamxH2G0+vxeKCGZ
4/+JhugIZPkpeYz0tyD2Y3vGsd2mzN+GLxG74rO+YgpdjdqrporGom5TMBrhnGeO
5MZj/x0l6iOHlkI/kIHRQlteZk5DXk+MDbvAIKz9zacYuu8H0BgTdRXRkmoIV9To
wHYgTKEn6BQuRrt0K4uCOC2zDOR3hqMWWibMGziQ+E8qlXW+ZrkLgOTTzxa+jJoH
tGAg1KMv7XBGNzoT/o1XpLKyuSfuMarw8/01NkICyMEvHJmXOzPxGyePZ8lxa64c
snzQ9CF0mB9ScdtvmX8Q4/i/1zihq45iHQZvcIObNJitd6RHpmu97IR1qY44duc2
Cq2AbJSOy48Qev+a0xsY+ss0ssDjHI2BwhCrHnEzM22oXP0ZYcGslmJ83mZycPCp
vhXYG/RYh2X7iccK+IcK8RA5pKCeOH/WiluI17FXHTkn6I88ARN9AR9jHE7bKOa5
KMAihqQqUNNmpe8dGwDmyIY8gu+MO82fRFNxXkN9KZcOxKKFO4f/W17uOHS7vc/p
4HVpT3JyvXU8L2WfkNbuCubVBqJWkKuvdX0EhSeaDd5DRkl2T6vAH6PabTYpN/+1
J9BOkxF5gikDgWJn/rklVmUIzPNniMGW58RvUUXtkWeLMrCoNBiGiM9x7n36S5cl
PYbNA0Kk6OrgZuZ2yCLxyVl3zqwS0jyGBa0n3bx11qO49i8NblXqW5m0sPi9Ww9A
JuMI/7MNUgrE2vLTpptYdXpyaZeI+mfG+URp4Q+QR/tdvzwYuEL2bi71uezhDanO
Y7Yq3POMVaAWRAw+dLKCcc0fFDP2osIcsSc95CqFp6KcNYwJyRr5RudMqIzDcGhF
tHIW2Gb50p7HBx4rlry6vsELtDJV2Yr6PLDkb9BEzrwQBrWDJuAWi0OZL1AcUubJ
1P1Vl2i4+G1UO05G4eBlh8DeOEzcbOgGFoJJMqIpcuvaCC8F22C/jHnTsXDydXJu
xRnGVXtluTni2ZxorIlb8SShpcrO5J8+MVg86C3LSXPN1QR0e4urwrgXOzmhQk0s
IuXLbo61/Qp1izGCc4MB3Y2IJpmbAvGoq0azeoLt52WF4YRHXblhPwzWBZVCzA0J
karzzgvr64676KjVdJEag4qlxTMldYqspEzPNQM/rxO+iyK5gEOdbSz+Sqs1tgWF
mpMop7Zzp4ybvg4SGWNCDLZkPrhUSx69zexpiTETW2VGYiRZzTdDHOy4U/0Zfhza
HcTDkGH1mVLiiRfZ57aHZLuSMHzMCUSVD4p1rUFziL5gYgi5Er3W7yAPeakLJK+M
vuOKZbOAYQHEibhcJRmic28Jp/xZCgdb6CtjxI/px9YNKRE0EWtzrQNykJhH/Olh
Rc5U4JnrCSug3sas+7o4T/F4NCYVv1o1Ar2Q4pNTQxTWtugFG0OOPIdXMF3tPg4d
+k6zQRyDoD8ip8zQGNI/I6vQPW8b+a1tqc1qEJGwtI70Tdr4Cw/yx5r+VI3NDF1Z
zFVpi+gr3XOaTII3252Um6Se+k8KvZwF/ISKaQOkRz+8aUq0hI8k8easqxw578Wy
3JEvw8LmFSloA28HTUdCCP5ItKoQJnpdz+iK/x2jYrQORvRdxWBFrFTQMaRQ/Dxa
6FTzdzFaAb5JOT23udKQIPC6VQX1PibYp0Z1PrOXwtOp7u2OlcfbBqk7EV/DaWIY
b+leblKRJIDnUvKKay52Zm6GtBkupoPvP0aynAw3sPuC+4BA4biS3WySU+hvqDzj
pFjHnSb7b1Z6MQLS4BeTQIINwM3Nl68CYYiCRxgI6B4kVPe+HQn1cSgSnlUe7Tr3
amPyitMq+7FIIWcMGv1H7AyzjmxATbO9mIC2rze/T7Efbmjrr1dzocvuouF0AVOJ
710IqYRm5aQS2y1EGTbEXg6GFbtbYT031MUz0jVxCyrIwWDjHgEEqzFO27zfPvA0
ic6Qzm2OglLEteUqbCqB3AFzo17SNNRLDuWqoT2yEPlQpjbGDFg/ERKUw2GMcSaW
71KtT2lA7wgluXbhV/p9fLHjd/wrfSjVokaqKajM7yC6sE14Zdcbxy16RUcSfCcn
yhORhZYMQkixePTMjbWxbtVraNnMyrobhKL0r69ip4uAbD479PPYphW9KpOTL3y7
O+YlT6Qu0J6zQl7t4LUuuF+7HLbOAvMHwJFiAo6Hiqd68xv4dIYELHqqd+6zX+Ti
E5YZUw8FHnGh1L95te6BRKnSq+sDU9b2FhY/ijF2oiIWAP8FUp6qOIOrfYFJcPaO
90YMdMvapGM+8hwTQ9LJnjx+8mLNnO93QQGnQkM4wRFZf84MB0i7mS8chGk5UOe8
coA1hWd1Kc2pdta+fot5wO878aHkPhpf7UETyCraCQDNPqOnvRGIs0Hg+6WzIYWy
cPRbNtN1EOBEKCVja4KZ/IdvD9tHa7oeXSymLAUZIM5noxhN0dMVk+Fqn9NTRSR5
w52yyp0110lJKUk8YjNhFaWecFxnWz1hRTaY3hFvEMdRrm0R3fNFHtPdpvNQzzxT
BzvfwcCIMVfmzSFBHX+sKC54P5+CqPGCsJCqJ5rTEadVZGzjcUhOnM5kghD7p97N
TjpvGcpayxhMqqrx2ymnWLL9FX1DgLsF6aLApdjurJmarevTX55La4jeWYOurdqm
/fCUyVvfNqbiFlWcDu0p8CpQfhxu8aP7NXqLoIrMcVztHQnBKqg+M/bHDoy/OuHz
bDZNe7irRcobibEIGjyLd+/FgwTcShetuEPxZjnhO0JkdCUGgzFdo09PEjiMJsy9
IsKYP2JJcrs7CoFFyK1dKthRVxCVEWd9Xp09ZL0IgLx3ltWSw9cH8gs8a/VkLKm5
XxZk9iy38DUwSSKm/6oomD36BhN1A8Nb+b/z7+IOp20Y/O0wo9KfHDHOSSZDW32N
rJzLXmIMu8GXi2UpKeMMINI7bXe1pe/8b9AEiOV+oen83/0KtAupViPy3+2QPWX4
QGD5uOmoI+uMyyomg9ExJQjzLU0hxBf5pQWCfe9FfKOIXXwWxGIPLwqWmJDNDGjW
aLgUM9KTmlXdSSuK/NRW8p/0FpYfeepwXwSJIDh/b1t0G08rfKMEVIec/Da7tJgq
NsSHEyiHzugomGxsxDw7oC8Lbz/IjUQAqz0ffvpCPegEplWeDnT2Qq4gP9Sa5Ima
z62ktpFf+1L3WOv1zSqLYMOPfAqC/B2q+9FMDDSqhw8L4wvHdz3paMZTTozDbkpB
iLyFwstlqhAsHT1D1DKf2KTuRuHgSRNYqGSYZqskb2kV7r+oXoUncCQpIVyOsjMs
wMWhqvyqHz+MPxzenqUb20jIW+9EWQUVjq0YRGeEf5dCSMwEykd15A0saGVamuE4
r8B2Cei8tfSU0H74aE1UGYtl6YFsK4t7ZnIHPtBXMl/1x8lFEwmRpkyNzatqQNbl
z2y/qQ3cpqXPbCCGuAmqgBlAuJSlUzORmvpf0eK2jBd6M5lulbz1kyvubUejD42J
DaKOGHhlMU1OnYLQN8cg5N5f46OgqzludjnJEpHuVEUGos2kPZKCNrg6kI/MEHyr
jecJQIjxiGvevdpRZWBEY1CaDcXvbpC2AE6N5yZLdlLlVTK2g5jhu/cT1MhiHR7j
s2lrmvdy8Y/QEZSezipZSyMwkyjHbViNO2aYMXxq3pCQyYYSDVsTjWEkoQm8lwrZ
CFzFJSmrKb/BS7jL+LB9CloPUwz8v0jO6TMtn68yMOJE+qYrdTAN5bQxrQVkvTxs
//GSr/9+6nE1/20IfTfc6AsdroLUCoEfsQlpUeMIZAa6vYC4YEnzV9mVUVzlIcyr
1sSHLkm1kokjGD8nbaI/AH29DI/uS0D7IyJbUVKne03G3dYwDhAFUr4XW/jFhtrz
KPIS6cVzw40KJqQhhqO3N+wSPyJDBkyGi2s1GyBd6slbWNiVL1Ps/z7ei2cXLOUH
3y7dB3KGUe35nqLNvdhPwrV/AYYxtfzIDDJ9QGeDzqw46HMhuPK9B5rFMpJmlHeM
AznBQzDoSFf2E8O8F01YvbKgtDVLsmqBuD5QFMrEa30bOZdWfPNs7bP7SeQc0tp3
ONdjg1CagRlK9rVSQDusdqoNiW2RcU1FnFJFFvqavVcfLkFd+TgOGTkf6QN80oTn
beZq3FU6J9bMZJ2CO3biywga/uDm5kEUT4XZ4T8e/Gth+jwriA3mi0YKQaepHnUE
tLIv0gt5Mu/It53kjSMQsLjdaWmF/X/Vh2YnAmSKnRRdGBhag+LAzP3ItZFP8aJY
wfpNImWlpCtBTwaa3UFBRjkHKPRWHrJQgahxXUyZcIAwtI/CVUE4WlZB+Nt7pmo2
USIMVQk3Pca3j63zwersfFnmrFQkDgSC4FA3pJjN+mhXogQc1m0mAdJ19loxFMGR
1ItqAMyOUjoMcaFdvbS7k1zOZ2mZH6Gap1ALV48P577wJ+suiqkU+VFyaWS0bTqY
G+RwmjuVstG6750nKlrUb3K7FunGn31k7v0mMmTiGkecRAl4Na/fImtHm6NQMQ4C
IZcsAZ4s3i2K/MrruQ9j8nvp4V3BF6MMbJr+3G6BngvdjFOD5UEeBpDp33tGkDj2
XmduXUi64i4FYpxnj3odRVLb0nK1rynGgPGd5qs6PXm+JuZtfbPC6tUXyHJv7INq
pJ5dBMN64PKRBH1/4OEfJLuXizdfCXCfVWZHzNE+KVBBtbSFfmd7V6j3SDWXW67L
lb/Ji+T+C3TejHgad+0JBmGsYurlCR9DqSnoiilTE2WuHoYmOcSrGz/dvWxjZvni
Zre1s7hxJ5cYcjKA/wxHkCLc9JDns2hPw68LZN1Qk2TGhtTIc/klhKNEqspiS0zn
fHq3Ok3KiSGgiXOW9yrFcWBdaeUCtBADl8tY3sSUlQ+tF4EPbk0ELsmxFTs4FVPA
yjdyKN9dn+lhAkTgXsZfzmxkqYV8awQA6cRQ0GfE4IdcmKKgBroOu1RRr0K66bw3
TK9qSNhktgT1LpB3DJR1ZbUfcDJemkv2Bs61MII1nFVe56yUtFVi6SIvZwTbu1qm
ReK7Pb+gKQD3VYAlPKAdbEmq9/V6lUj5GlG/F1D3lWWeG72zHXnFvbCzavx+ekB7
4uyMtwCWSSFBqi5HprE+4EuFYN6sQvEu98SF51z4sBVAWpcOHnJfNEt/j5VKa7pp
p8O3K8S2wNEYpGc4pWysfMETDux57j/hhtD8j8Ep+zaBgPREKbQpKPqG2+G/HH+a
sCHgUpLVG3P29pMdWtRbWKbQovO+ObNL6mtI8236AnJf/T7/eb5GUDXRsCDtS7Nq
hQ8W0zZqHl4Cd0/0GNHOf+ENOSSKvO8oJ83IvJsCra1lEBva5xTnfjTZAmovu2N3
1qGAgsguVbTdwwylzA0OVHe6MmIIF2ggX8FR1vtdWYW5qPpXUEh9fZPHPteAgeig
59UjsOR7evG9a0V3aKCTq7dQYeBTmdPMgJyJ/iIE7mNTsPxTYGIkJTS0O7OTohHe
PxctnK0Q+YBtGlx1/LgQHdIbkPPmEB/vW1lXG0BptTEnOtSKyw0IrIDehpp6MxPx
EjftpYlSs1YjWlPBC70yhszkv97yiyDayUlBHlFPrFU9sA3MOjk2/jsRbfvng5e1
YCFLcUr5tm3Dp+mivvsMjFoid0kqEz2LGqSCuGow/OvHQdE7eqNbfUE4k2nDKQhJ
mEbK+QegObyoImWiQTJ1BCMZM8lXp+JsQx4iCdSIPIAqYZKkAJJyDOFjx9yyn+wk
2nRoIoHcIWwTdY6Pt0jNvfQFKJjQnubyY34Kc5pTQj4xDt471K3vpMSPwOwz6Quh
omyathFglNgDds4SKps7XEAZEYibO9Br/EytXgLsHwmGo7xs0qJBgnbs49oeNTnK
Z3k6rgHexnZWkfjzPT5LYHLqLE3KfTRuoJK9GiVldriamezK2q7deG+/99Y+gSCj
Bw1KPdk8uRjMVx7qGwt1nvPdwtrdRx6x82QuNnqbTEGmxKMycDy5B+8wxiAWymPb
Jlh8+7PtzzdNuL3WZ8Czz8Y3KGjUWAYdW1QU5vel5vkfvtkgQ1/nyC9J1XfVV8+e
7nDBe3kG5BVUJDITYF4qqgXzT8n4oIqX3dleRhw3eVAUNtQ0SYH6a8OA0/SPCxbe
AFONq0kp2r+XwgMsHbbk2pcIlzVdi/Nh1jUKENdFyQaYfsuMFzVTnbGYNh9XFwEc
4MNiyAfLjuW3ensKDOOn6CjXFeEMZ0OFE4OzM4T8zk/MjRqb+31Nzb4L6q8HQUAo
mH5uDyXxBgYjdA5/NghXikAXh4D3Tyj4WeD/6cVzM8D/EApBlfYvYRpJU1+qobJS
C6v6EINmAO43Sv5Wd2bUP/tIVPT5PddpR4yTI7pgLlbBsjNpmA2gEXtQY52JLnYO
9heCVqijcsGrDXg0zZXkmuru0vdZrYLQFhmvhy2x+kKK5UqWvuZzAu5xcg9sKcSY
yBN49ITsPEZVuzuqGhEVx8qPcdw2g7ZGpTkfUITEeFBclOc5xs2Ws27BL8XosQ5q
4O307ah0lxsEKdoY8qTmf4Ul4BnEU8GQnZhegYjBmtA5nwc/NlTbi1jQpEpj4ThU
8Au8I4QCpNUACrFl68RijfRcKL38zl8A7L0wfwrQdhMfZ/v7H43sRHGZYr7G8fIR
CqLiIwYomo3me2pnH25+7HS07K9kVKuF1+4FvEbml2U/fHyUSy3AtZdl563nyhTQ
VQpGKRc2xM7gipa5DKLvJcKJd0uqkxO5ENn0zpw9zohbuerl1asrN4TspolMUdoZ
yo1RQskzEtywv9p1Lk0LyIDgU/rpP5hq0F4uQ8uEgW92/fYtLHIVQHxXYgyl9ul5
16ZPtJ8vrL132erCzWrz7ubbIU/g4mFrfPzb7XA/mKktNQkUFKtcXum4jTvtQdLo
NktKrQDZtX8Jybz9+xoWOI2c8Vayfbbu6OykyW91joqCG7dNrR3BiN1oiUOpbbBf
JaOV6NSnvTzsuHqqt8juyQZ69VDqHC3dC1arq9TVUQ85FOMkgz8vBviXbbbq9atd
OCtC+bXkFoxEeIWeCOp2yEDQERnXfal+wuUNoOUTvY8krEzSjHa9qzkSfA0xamGn
uh+DPP4PoMDLA9UCLKamdBva3ROWUMRZPLBnyPpx5jsbmh2/djZ0U0/17qIcxYBY
FhXqXLhMQEKZ61j6492pIrwHGbuhXXFBOsh+GdYZmnMTgWY+H4VehYz9RnAP6nAd
yoKDeXMVelF4dMkJGowG+C53o4BX6ioNo0B1LtHanX3VFapIHu25tg4Er6xMYZor
ALMPtQEu+N5nKFkY3Ksi4YNi/HhEHktskbLzbdMxlJp0M17sUe0dCZGae/H6Adi0
tw0cSJcoD+vMgnM3NTXfRMf+42Y6RctbUjSveEANGhfWoBqVFeEuu7ZWdzlJf2FA
/PXl0jpFF7aOSn0Hu3HoGsumkWlU/UBDJMuaB26iB2Z/shjpoTq2N7VLXXW9VuHa
JNyNAglOZeQxNGJXzPbzOC6hI7viKac55JPoRflT/lQ8YYpkyE6vW8/kZADMmC4p
8tlrncy1VZiIPgUjDduBRyxmBT699TyNE1cvBPVXAuNrFwmcHD5QmA21ZSLDVR5I
dNWVM1I37S2BCAuMRlrCdbaHD6mhsxY8NWAECyuHTW+hXQQQVYPELootzCJNGWtK
eIlW1YoUSxhw8UEjR8EYnhS7Vo1GBkzrNdrD+k7Yhq+1JoAsWNRqdJeIXBb28dWZ
F3Hi7SU6Eg/SE5+ncVXFpjFpQoP4r07hRMDGviuM7ztO4sliMOdbad1Wed2VZ7sp
a35w4GNNmA0x+y5smEKrEq7Fq9yTbw7N6d5PC/La1l9eCz89S4JE89wo3bzZZY7L
ed9LzTkNamgZt7ppTL69rdyGTBEWtBKB6CDsUn67CbMRzZIQgmCxRiReCnluQdD2
2lBMsPNn1cObSggZSL1W78A1/4NGXWi7SIsx51GyP0gB4yBVvwW96jXGyGsHzzPK
vSeX4QC4vbuhF7pVysb2VwWP4AGV3TIoiUBcsHmHZOA3nKdGcEzVbsNX1ZQAjhJE
Y7PetzorNhePWIORnKQVHbq37h7jhkNJU87UBAQUDOvEJTChF6cP+m4p5lBZ/sWb
BbSuyKE7aBryvPk4zoCloXUw9zkX0YzLqKb9bF0/BjR2QG+TzfYvJR6Q8HU+gccD
YXA2n4jJ0bD2HHNlXSc2kgX8P30RCvfvXvMEV45+hld/GNtS5muFKr3DPsFlX+gP
A0rXXgQx0N18LZ/maQ1czYVNS4NeC6HIGhTMO4C1QWEUmsjwLqveit3hFYgTP9J9
r5Lj6cXv6lR4rXmqQs9arUWJn0zLvVr59hc54fsFsxtovqGXSL2rRRfEs7CpHada
nJ7dk82MMUHTSgpapogxbp0DEn0g00rKpQf7xJ5Jx43GjFkIPKHhC8YPmqQrKs0x
u+MtopPKjmLYQsQ+d/Ep5gDVnjsrIlLfPM/b9AxR7sBd+toMqMUcTaNtSw0Prdpa
gCoGDDVqXIG+efc2kcjJRLgs/W0JOORMSqTYxZBZpNSA0buVXUg6bT9xv4DJLHx6
zQJaMmqkyJsVfpxE3b81JNP+ZBJ673zVvGgQ0XlKrtA1iW1pBPsT0wZyw+SnSJmN
nfjzv/FxMsubmzdLjbryi+G4R3xIuIPeLFcuhO5v9q0BHg4X0M+hRewJBw3IGw7x
ZHt8yD0pJcXM1GpIEE9Jx/w2Pgd0sosgzULtL49IMJhD6AZdVz+sjqfeJh+C2i/T
H7Q1biOAnEf9Ju9wWrjCMHMbFEKmYKTq1EmwtvxVldq13kC1vHt85jo3hqPvpBL1
83SyL2VPL6R+RAg55GlBzkWWgkpDm7DGMhMe0lbNzNaMxsNhF5qJ3rckm2SxWDVd
J9RB1OOi0A0zZ132CjZn8X40ccbmYPmSdA0e9mKsc1VDOEj/azfsCsUzWGFlo7GS
WiUWhfpstvF1XTaC4wWx9XZu3ikJ97vkAAbEUd3t/GR6Jrk81yD7f9YO83X84X5r
82qAxAXVNGVrHdnIqpPi/ZU0KQcVkQB52yNK7nbCS2ugCHHW2u00rXhCazMBIsDI
8MCbD4r96xuz10SoqBS1M17ALNBN5yeVoj0MTiRjhQLU7zJGdiK7adAlKoJNxABL
Aig1rxWTGYpRzGkYXgxsSqtUNemH8tCtKcE4bHu8Mo5yceBBj448FRtGkOsQLE8b
yJFh13Ia81ZZGa8TZDbp0F+cpOWzgMyzYyFoItDzDhjqVD+HOtmAiJBvBJrifk2q
oj0WLdzcMRKW9Nu7OIGiPPulmzZjeN12lLiiayFuZKXhXC/Td0iIlpB2ij1ht8+G
TaETQ6xbopbVLHKs32KZCVCqYGEY8ScXXYVjTSeHa+uI+MWSmHa4iN0+VujkQAtv
0XDmlyZwp9Za96CIKv7buEOE0UiOY0H9vC69Xh4mscQ3kWEiiH9Q5+0NhhxpPblA
W/AaKaU/06baL5r2ZPE3oYA1XdyzlxCOwVxCjCwKLBm8a4wx1n8chbxd99OjIZXE
jHmjxravyyhOTKb8xNF9/0+sBWHxsuCaFBZM+/EpLuq4QgLPT++qaPqX0xuIldtc
2LVd84OrmpLO5+Gr9XXhI6TX0AhihJxrNQo8lUYMfxJ4fs84AXns9nVOVtEs6nEw
S2LRiJc7xY2uVt+/ObMdgZRbUtI/62JOLVcmPp2nNqCY4xWF1DCR2Mtnsuu7JLhA
ONOf3kdo7W1QF2Xkhi0gJgfpAywnTLU2YO0BKCJ8gzekzCiYjRFmaXeVXWH2tpbS
Zb/7KNcKfwHAF0K3UXoVM2E4qAr/INN1Hz58U/WcC+gExyEwI08Q1PWpvYuBIvsk
vyaXF8zF/WDw2D8FtOrj9uGEWXeHYHoT+LQ+gM7glXNc7zhtvMg8o0EC87KgE6oI
efltaP/H5z2wnPC1IAAPQbogY7jxPL4xisa2IIUbHhdc+l9PS+uiBJzSc/qhrFDt
+3EZyWvswa5r8lfG+FOyjji3MBZh7N2lxNN6FWS/WnaSpK65wkA1QERN8fuLQBLB
XXmG/2RAS/WPuF2gnvUSs5igkwVvdrMR48QCn0Tw/cDzGE5MjngR1n1Vav3EKCaI
MNbNYb3BG0iltPFnKXY0ZJeFK2sc6Fg3z0l+lQ5D4FENPhGKz9STma1ujidLcNvS
mEcbFQRDGtptJie8jr+HdMklPkuT4kErkrdVXQAwnrDqiw6OzJLnf4Unfmjkv51r
8aXJD3aB2Ss6FigQttorIKGyvB1Gd1mgPGY94Dgz5Rke6KIU+V23iZ8Uz6GVOTFm
MtJ+KXfI9rtAsiJDFTQIx0FocKurBXCkm0aIb6lC1b5KrP/5qMmThhXlgMGrmjp+
5tHBrO2erix+Kz5T9gaVIsMzSz+CSfT7YyGXCUxWEnnjUnn8eyWiEYDY4k8KhFka
jK3DOOlhxQX0FVz2FgcFLE9gL0EPMjFdE0YUZzg+LLeQy8o+OGPzb6N9dYkV+TX6
UTwKF4iX+YJNP7pcbUdAtZBmxS/QsRY1sTyO+ZaxEL1LGLoM+b14XghVIyyC1c/A
/1mvOaW8eHt5lJH7GlO/TfLBaQZLGcGzjXkoPw/1Qb6sJAXTVxinelGhEiPvYg3W
ejDiTpYKHRXXqNA7JL5rywIYcJYCS5ZPEW1GH/4gtTjfeoSmxiorCnQISyu8jlc4
VgbLmg9dbx8gKyCtMnAR3tKRotjp0CBdgXFp3dcXJS8ZLREz9Qf69alFkgWmMOMo
Wtn7k/X+RTXn3OcrIjE8VBHWQH6Ykv4txlnTUPjwAgj7+J0sqRh1xXZNFPLQ/lJh
XL+JDNGbntZmOi+IuSev3wIKGQP5cxCSkQkD4BftNo+FAXDjn4A+uvlnlk3hEddQ
qhbFV7nyYCvOQc83RHIuoQGTSfXDFqKBtykZ2SZ4ob1NeTeDGoGNXAQ32/wRAJXe
9DFuu/wOlMEj8UddXoZI9K69W/pqUVCSRdg+UBeDnQxNCbjrd9ZPBNvjR/hrCdVV
wJ4L6KSa3p78iNAPSvQePibvjYkBUrF37GxXFvgoR9CVvjjlxIXl+TYG1q7YItnh
OWnFASEjD0aD+pwCTrZu9Ur7LjY4HKWBoe56kjvUE/3KP9my4fPXcu1pcERHFLG7
T6APKZ2Yv5T2dEZtd8yQxU2KQKSmiP3ha1tC4Y0unZQ/J9lqrmga4NLUJeIiEj9s
xPvsIHrTMZJy2zRJ2FrNySBIJf5ydWd4txZJg1qvm9Ny2uBOgPMXqMTz3sGvzBF/
6Xgs6NjHoYHAu1sJaFLDHltdBYpJN1HxUQB0g/y5gqRtW6F6i5VVtVCSoqNOtUOC
0tqxHu94o7Hmauw+adu0rARdNuYF35Hwt6F0qDh84lSJXlL1PUKLEP16nYrTZStz
3qs+WupJOuvJK+J+d0tczkTpCBOMdhpMvCRjaUmoNUE6NFhq29xtsI95JmU0iVag
bHyrOnFymryP/Gi15A4+SVxRZij0r8I1u4HhVcT8+vZyrtRXXdhQeC38Q0lU3Zm7
aBN5oJ6HvNHg5iv8aZXrX7sd774SKPch9SU4JK7C8bz2AWO8r7Z8SIXBBuFchm86
wZRnFfKBY6q3MawgvNCdmqNj899fR2APlgGjr9mXZTJRyKhg2icICjyJL7uWGHVs
ayPcZ1JuD/xs+tKBVxtBPw==
//pragma protect end_data_block
//pragma protect digest_block
YusVbbCAzlB6aQ4klWb5iBMl2bo=
//pragma protect end_digest_block
//pragma protect end_protected
