// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
qP3aAqeZyZA7DfLvr1jR2Kc7o+Y76uygEmYfxnnIDxVdVW9tyKioOUVMkbW074Yd
Gh5u2qRJc/AyHOWkqy+GEivYts8ewtZXsC48Qqj+/ql/6jeAEN8klpihqnx9hqtr
lDx+ISVhl7Qd5yr5WGOTZnS5kMV7hNtsi8R4ydzn7q8=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 50208 )
`pragma protect data_block
Q8XrvxSf12y8lm3AZFJ0c96ROp++DJRaviUhmEjIAL4KB59fh/3Y3TWyTmyRLqVw
yLmAlYhBIF2zX2Rb+O1BgmKd8b3Oh2tt1GxxHWbhE1BmdEWLM5lv4OBb21V72LXo
ICRwhql6rOT9m9WDys9f2rE+W4eqIT/OuPYCFZJ+4EcYWwxRpbzd0CSyNMsKFSF5
RABMWQ7nz/zObBlzAuPWu2wcgY5G6dzn63Exk2wnqGyEcYmenUnHX1dnXrWJSZ05
v/FKbYy3cobp2JGU3C/NdKc+zDgUGtFnbFu7/xOFyROOs1arLwFiqlY3pcwPRDS0
AJz/wICIgqOIHtyEFSVtXUs4A7aXPDLjaBWjgNEsn4UzJVxUWSrV5P79evbRQqCu
LkClAv4ZV7w8K5gpigDH6oXFLggvfFWMgkNJqjvH3gDmQQR8N7lFkYG+z+P9EGV2
ebUstJv5ZE8HAMWU4PcS1/GGQCv9QanXQO2jm79ymCACJLIbdfJXiZ5ZIHYYtNPM
6/v4vLJjbEzKylhULlUzILYjZQeWvfw2Ix6V/WYPRevLouWd/LRv5BYDQHCd3cJf
8AbXYz1wm0NhSThfW4LrBO1c/X1gHn4WAPElXmqfm47JQagC9M9I33NcVtHr1ht2
D5jB+F8T4RkjMz7PHSTQZSec+5YoB1h3XmadquIZMj4JcyoW843AsCaxeyGbiRKg
efYxfKa+MR4Zw29JmbRQOCY7onxfQRTZwd8ut3+/Ne3oZxDE6CguTwrvmL7paoY8
dKnyKZNzlP8lX3XXLVdnmOsDTylr/QU3JrZdOSi+y0SJ6/vi20UF7326+e7UkjrV
NfuYcK3/LLwEgoSJnhF2VPD2NUFiHDuaLNW6oJCyyR1apb9DH6tCnL8ErkP+Shtn
e+dqjNOoaykw9VGZf9bIUrH5TfriMeAj0C/hM32Ug6MeCad/w43g29nJpl+MR52f
Eub0XHZVMzzVhxBiuR9b8u4BrRA/UUwPcQTtJtis91VMpcbw9CSMEcWlZPK3Gck1
GgghcOdo/jIXE9yxlkwdfuyFmB9/WAxqJz7Hz9SIU3iY7OCTtxWnM8F6aJuiIc8x
0AUdHy5LvB8w60x4jmm36bmrGFwjjSy0CNv/iPaLhONnwmsZ5JNKHV56CcRNMeuV
q/8876JWem5eg5h6AhfuTMjlPGdfFaiD3YzCclDaqfGNJxkz1zjIK+qaLGwbRLrQ
PJ+mvrcSBQqF9SC4x0DLH4m5EP/yyQe6JkSEtjVeQXdNPsXoyajbEIxepdwk6WAJ
JRNX31Y8SZr2mtjHfYy/d6kluh9qMtovzEHZBAMRMMrYefSN8RxrFeoKpUg40O4o
gULm1ceqUs8TuzF1RHH8XVurJj8+hr74qvoMMgcDelUuIFbuqeaR2qda9YXG23rF
IAM09wdF8f6ZYcULx+em/UJMU2XpzUXQnDdi+wHTEmYv+uo0d8TTsBH5RUvWgAHz
lI/xqMyT+WY/FTUn35Ww7DlciRWdn8WSSaEZyjSf0pglXRn2tP8NOgOop/QSu7Ew
qXjx7L/h4sg6XXVoa8pqKOp/qAONf0382J/BsCDOqkgSHALVNHtUaIL9GUsHAD93
0Rs28MpqtTiGp57e8CBjEo4AsxyDJiJKfSWU6tVncwy9KV4WNKpS+8FM7JYTEhVl
16F17pCINYnEnW6y/qiC/z45glZZaj3T4uMQDC856/63vXGev2Dn7dbUEtpyx57+
jTiodJE6wGOpbmOuSfYSZZ0ZOIok6zRvbsjNcP9lgNzYxAO9s14pkHdTB7dXjD8M
VjcObuK+6So1nj3YE8xAU2InhmXavz0IcWzb7w1PDjcZ3Po/7oAbIG2gR67sLwwx
5PfSWn7Gzs5A0wOSyIYgWmeLIaakB3AGKO1xMrM9XK6jrwHTv5xkLEu7j/ikzbCn
pNvriJLXs+AeRLBISuAN0QTWMy15EptPLVkjSkk66IIcbPCNZa/HMqeHpxP6ctik
YeaI+1W1U1UFv0fuQHmzIJ4nYTPG9LKaSx39fsbLMgIw6oj1chV1oDiVKEXT0x09
OKXWvsPF26OQ5PW9arT67AheUCfjBnSajL86iPkLqKDj3bduvbbflQznZYjcqZJm
lbqcy3cUcQ80w0XNBqGs7kVwzR2k7DVo29WZhxyPrtaHWSLkTYlgwqAIM+syse9M
C+G3K/r9fjpTVQAimyxrEiYSAqVRnHMtvachjg0BsnROTulOMTNp6LoH3X+4GD7c
qvWblKtRMda2TNHoaxE2IuAblC81am8kxahPGDpgWiT9PeqG3Rfq9TPVlEGqVfdq
NUQxPx/7YENCe9NBpzdQz7Wsf+6EeKhHuESQaumKYdAf2zZJ0WfPepTNEenIsBu/
zKmLTeDsnWUu7+S9owAEf9G6HjHd1EHNZ9WaQ/qZTPwF5HnkTKEa8kV5Pr+iJBwA
sau1a0JWbp1UUhl0DZLAE25AmdQ9ZLFFJq4Tn78zawL1wlxB55gDy9Lins3q3I5G
HWuFDZSE032mIWkZoafayqi3ijeVoUxbP4cAmGKeeVmg64funFA1Hgsyii7MNcc9
ZXWRSP9iXj1pRvivHqamB01EfTrCkmpkoPlrswjT+5dZrGa6Y0cc6XhgO2WYCXGK
l6pc894EMa/x5NfjYXpATFSv8Bg9X2fJ9jNoa4YZMOmMq/HMChhpUEDfWOvpCerk
oUWFrNUg5IarpBL3AbW7gtIcU7CmQxhhekwVqybE3NKtBfeepdzg1CylLU+D7rYk
A8RnAa1jJP/+SmG7Iwu3nyr8XX+nQvAmG51w1viigVBKmUNHmg3aBokgRCMUSzlB
pM1knUAF8w58wlOPglhm9U1tWbkkXVUghEEtZwDdGofp8wP4uvsV+0MggW7wFzOy
qkzXAbazkAhD2i1QTD4I9qzCURdyqwqbNMv0K/wNeKvvvBMgHY2N2qrSWsgky9if
M121Ks5gMfCCjHaFOC9CXVM0DXmcy5KhvPmF05MQTh2HRmgMtKIrkiN+IE0ts4d3
LpXEJXA0nyqCNS7l9zjccipsfpvAMJ7QOa7zURGGaEuWwFgUuGwryUvkn34LmwNo
z3688eaK+Q1vmliNNXLCUtBnDZ2fYjsLWFrQCRDcStaSlSx1IfcOjtQ0KFDPfXMx
B6Qhf0QfqIHmvg54WAZs/OfTV6vMK4XD96Pbi5MA+NEpBw017URlJKLAna2z7KTv
j+SXM1vma3Oee6gVxLkDEzz1T+tNbrYiFhOs7rmlv5k3Q77y5ZBWyG7xkMyKMZcc
4X4h3tBBz6kklYVN738jtQr/FAaqeea8FWecka02IGgnHdpT6g1jCOW4ZAMzOAsY
MbSGHKxPG0EkHVrXSuWXvKWMcn2V6OrfB0pNzkixunwGUnBomOOQk4QLF7Y0G6Hr
ZLrEAGISG/qEnangzNS5qiWHDcnLonXv0tVSIYzFrqsYr6IZMIS0hwld2bk8gvSK
64WrwG2vYOLZ+/4UaMkBmOOl1yu6yBKcp6aJNJRWYvo8fw7hJrQ+TuUNQJfQs1Qp
Ts1bCtrYG0I0fUCVnlUUYp+9K3xBCTjGeMUYKeob0GbfkEWj5ClPuycaU9uhN72U
t170hqbi4jYTFbc/zPwBXJvHjb3cjMwTmk60VU0sWtzgpspC+5jT8Q5rtxdKyWet
s298NLRE9ZYhwX1Z3KD+Di+I4MtI8X0IjZeGHrFco6+/j57Naf1vHaqD2A7J1dQi
PIWaRfiqp+YxJQOhiYZ7E++uDyUlR8EAtqyC7HEiUlclotxVbecCdKgXtnGHAfRx
NnuezTHcqj3pLwFjMSt1pmWXDJ41ve6lNtLzrtbpNO9aycD+NFRLIVBefkxewfxL
QfNGD5SlCzVn4K6/c5LtWxASjkYcX+ExBYTGBNA6ZZtymSINVhu1C2aI0MeF1HzP
8hcJihWbHZ1b1JOUSGfUmpCnLxnxchNA7dKC3o3Ve0CGwZvTFHxMGAVl/RIN4kZK
TusTTnxwX7EWSSgoiEpwbKTROKSTlgJM6j5/lwERWTgD7DBNFkaijWvdHJQBBpaY
ntopQslk1P3qwOnogox4HtMIkLhZdgjK6Mr0YRjOHIXU8qr5GGLaCUxtb4C4h4kU
O6OrdTCLLIbz12SPNgvSnVM9oim1oqxoGn8VTdkMtguRrTgMp3ZMfk/RPG2Mo7ex
zgBAd5fYlOuST5eM6rc+qrnrxsPwriTNTePft3Syycag8Sbl1gAuUV3abLav8/iL
HK5Lal+YJoDnluxSsu2m80wJkTA18zBGjHw8yFr7jWFvZMPscquWk35xJ5CgcgPT
EcFnCLEb7gR9v3wJ6G5mDMv4Q6/gGjjDjaK8P5TBMdFRte0COlmYEkyxJNEVU4i3
1MN4f+WVkVcwy5vwCALEAkiVRsSK1uCDO75/Ubd8tsu5zywQPN4NPzgQHCXNWRL5
32ohYPt9eStPZDWvtNlGCta1gciRzKteCn5Xq1m6WGBWLpGz7iZL8Htg0YGbdHzH
JNLxhV7uVdsGffgeYc5Zek0oTq/mlXsWJS6+Y/N0sRHMYLRUwHLfhutwO1FbeYte
aL5tZItorORXC1PpiCO+0vLmQGWEkfqtzNWc313bO7JKYRNYPp1TOiGhHwnvOYvM
uOsAa9U9mi52zlVw0OYRjiam31cAKDEwa/OH22GXDW0htB83k49thMLItT7N+Bzf
ow3VyQonkUDT8UJG7HlfHc1vcdF1CBSTY4xPjfQQKPO1WkqzRocy1OsUXA9nIUHs
fAiwC8RZilci5c5rarNL2+ajjtkipu4zP2qFqeh9tVGi6NsOfsbWO5vbCC39Wu6v
+lHFoZO18iVkJDcttb5DCSKXyr2PdSrhkb88vTx3lRpzxsm0XRq2xz4OIdDSvTk4
E4e+JqXv7sYcTboj9betcqgSC31jl4kWr1ShYSepmlM6s12zOxwmBNLSNlcTrXZ0
iPGPyFjhhVkwSh1P6wC0ppoek8/OqWuudhmvLgMf6Ch3gzOIXJGkesTd0OcQR4fh
DZK3WC7gGJDKG2pH9DFwG2OcYS9hjD7EJLfBmZZ4Xa78Z4g4wX1eEb/EEK7MnBOH
gh5nmYvgLSMyAmi4nDzIVvwgxi4yrubij59m+NYIY2fc8Nb00OO0SI3pMY9jmilv
hv00RC9+ovnyvrVIe+ir1sn3iKNssPtgrhfZdQkF1F7NotLJu8cMJtN+bFoXgP7i
mOb/4Si7gHRrYr5qZqf44/lNjPkVbjhy4nzdFp/ux8eVGSAxcV/senVHZY+Z+kgl
pAwDC19a/MwOUcqICiyYABY/vHnl87E2LkaUBC10O4LL0x5pKyUSM3xGB7c63fYa
C+PlYLfeaQxXwC+pLDRsAcJaacVdWMOiVijsvBbcNZLIJvTkOJrle8cjIiyWfCKV
C5VgRb6gKjlwOjc8ZFs7cKo/ik1MUpo02vtKRFv8EFS8NDn8jtXYPI9zezZfIC8H
d0c7igL/6l7NEBhq1D0IqANqh0SgG3/yAoZc/BCaE1yWpwpFUjW9B7Wu3cGeznGZ
H6SXFTU/v7BN7o0BIEBbnbIBLJ9Y7lJipXDfBZRzvkRcOiO0IbCg0MwSstrPXMO2
zO3VvJ4tnObYKJwDzk0frEXGd5tFMCKrevWb7icTqt3JNGLQrVG2aOlmoUGFi9I9
4BTwpyrVt1dMUMvmt3vYRPWe9waCjxjCgeNFKUDvL/uLH4Kair7SMdWClZza7Z/k
31HeEUXeDF07aKA6e6zi0hIpEaBvQ/zF7WX4gT2A8DvzMY0wZv+bzCviYasFKfmQ
YwvGn+pxjLNFeayep8WYHeM3K3/FDMoRpBUxXiorlyxeqIXwXiAiLzkfTLGnnWi1
wOIHDl+vRo/pykVbFmLPieE2uBGyRCC5QH8zszbeA95PlfuP91kfatu5vwNvve11
FktC7ctPE/zavXUSsFvNTlZcVSMUEs/OzazRNCYUN12vD476OAoLtOLlARKRFG/h
uTa09Ib+kVADSxWq8JuKYg4rErC9hwDm6pEwBpexUG65QNu4NINhhgQbUzBpfWOY
nrPVhs4xJDHLgqaLf6QeFh7nvTx72UnW6nS9Hb2ysETC2qOFvxIgMFQ3OkWfKFjV
cR01hmoZeLnvDuyTpIyCdgdRrfaURM5fOyF9z3PMG2azW73ctje3KkDRR31Vt2To
3NeTBxyDVlBCi6jj7gY/Mxd99INK6GpQhFMbL9oKhHRfx1Hq1Sce5oVgcqu+fPdI
OrV+f3HzwG5k73HbSFElMNu7xYClS7o4UmEFJzkErRtr3xuOp4nig+dBR7T5vUs6
Fe1QSrKTZiAVIBHxPGah7WNqqYuEs7bTdP2g0DnNvLCNgj2O4zOA5NmY4/Rw2yhX
2a1vQ956ylhSNi053AW/WQ5BaM9yz2kVBW0O5us56ETWnbpjAAuTjmZYI9h8i3W/
oiN6XpdqNUN/3bCz0dhlvaRtiTqBn4emolqnP2oq+ccxnxYIEkR4rKsA+FT2Dqh2
iSYfPjrique6hJgvNmn0Zij7DHV5DcUDZ7uSWtXothtXertQ2Cs0vRvC0DcGtesA
ZTgKGwbmPDE7PAUtgP7uLRp6ws4uToI8cfBtOLr7E+zLPgivphm6w20hEVbV45ty
miFF2RZjuAKsA5mw9D5rKoCnF5twTmdivJnE4MWXdyFeaA92P1JxNte9jB3OBekv
lmni6uQfYtRbimCbBTQOsRstKaMuLxoOLbn9qYOD0njK0z5X6i1snkA620a1Yd2L
7W6W0uofYLY51gLydYHcIXfGRKndX+8C8zrmxRlVAf4P7NCnVW8ypSuyCGHEkXCr
oJ976AeaNx8Gq/koUICdQKjXB4dBu/y6lhWE5haUtL1zM0V0ISLqDFJIJuvq5s2l
3r2VbsAVIF2/jcp6HW7fQeIP9G7yQbzb0dvFt6VUxHgQUocV+mYHDN7FTMlUOOlq
E9e1eQmijaNXhup2/Xvui0grMj3y8I3vVRonurZBDAICBYc2zzwjb3xnQJsavmAM
5zfaf8QTy+wKPnCI+SW61Vf1NNHG82rlLf6FWkQxeCe36gyKwepscFUwIQQfMuSI
rIgQjcOjH49ruKof6laD2t+7+zacDN2qn7CnmPqzzniMXrSxVgkvrOJQc/CAP/ZP
Mf8bLrDQEARgrV1BX37PaAG/HrcN4vfCEqIInLLJhLGe0s5ONH9va77rCt/UnstF
oEMLUXrC14KJy99Mz0QOQGr9K1dKbdKw7LhjN/wHLnel0s4MN1sT/ssJ/vZfkQYn
bPcgP48c/voN4Bvr3C3xlkX8N0QZrxrZzQSIyMW2Dku62cAbFTAlVDv0cdtZo2+p
f7BqwPVmUkaCOD8xAER7UMa/wCLyAArDUT+Fprtm2Nbss0UKzFnnzGt2kKSW89Oi
jrCVZVzwpqIetmf8UaV3Ebdnhcf4R+cLF5LUsl8tqDqiQ5YBZOGIoPSeJDPKIib+
vMPiDU6X5+nYPhDakYuaN4svQdCigI9YVt9+joF6gPcfhHGreJ/vkqgIEyaznbKf
9/0habnNkdwOQyv9EbT6umtqMlP87FXOGLLthtPRCkPiTbm47FbS31moSzfwIyFV
6O4gBFx3gmHFcADtL/zxWYkugb5SLhPFXqj5yQqyObx0yY0m47vWjr+5sYJ7RPQU
LcOXwWdnUCE7zfnT2SPF01J7sC8xMK9D6uOubjECNLrs7/JGIrfpC8+/6cK6ITX2
TgZhy1g3qNID/80nFsKXoOqA7lzUO/HGmWhL8qhZARaY2j2YHLFU9dIsGnM4qBF1
fiwZozEuiyX9QW5s7XJsq7DMsa2/+FMNJkKv0wc6MHNvR9D+T2yjBpZ0evRKuNZk
FSRU19zsoF+GyC1wSpfrbQg/mkTXAScjXXRmJ6PYbA2TDy4DRRk6rtXUAHfxrhWZ
zzhMJSwBzTB+5kNoAcSIfCRVToRmZcdyA7cLNQGHJf1w9ToQQG0CSJcbqQX8CqTG
HTA5PuH5U96dpYaXj1bH+XqpJId2fIA1h/JfipFvJjEcuQo+O4y//Emw0UBgabXu
1lXW5o08/THzwofoImntMhHq3j43zudeYq9B8QjUVZRRcJYCeqJ+Dn6xQ+Xk3bPR
YHqVBVUXPiYEDLtPjzw32zIwkSVSkIYwqy97aSQAa4FQ8UnvDUVTtfQW0rTgyJtV
hfFVbGjcNWiJlRi0ZWIDPBpBOKB5zrRJlVos+J6RayywSF5Ijwp+HOPzb2o/ZobB
A8Y1o0k19QF4gIv8SKbh/wZoqxlf7kPYYuBdQH2+51H+5qRZd7TLfsSX0eQ9+Jce
1VJb085q96i4F0vH28xamrDoAFmURCJ4svAYFo+n1XsP6+XtCvrzWqtrZ1bxrpim
VQMT806PF/Cox8mbFp2FV4dPugzw8XFn/102fgd5JNL7o8V1J42snIryLtn+S5HB
+AVDQr+4yQCWFq2JgAvNxxp+wGXiiUjsFJNiBA5UEf4tVu21R2Fj+Kd3KXz4ZESC
pj9WhC58Wx8ztDm6ErD9DhsgoTXuVCbdaEXrfzf3SmI3JOFOyzd/uXLBZg+7eBuD
EfZzOiEPjxzSXw6ngrf030C8lYjS8Is+vf0dTRvDmwjBicZSFWYlJW9VsTFJBubt
V44xJ5N/k+m/LdHsUwXkMbKacGp/ckHdY79BdEaf2duSNKQdfujz9uW5YGUDzCIs
nagiuiIcFi+eQgW/7DsqprA7lPkE5QL4ifgzf9Eu9AbN2c23tSOmnKYkRG6xjeXh
GjqQPHi++vNJ2OAMMluyjDv5v+W4llu1XpgeHyWuUbKzwLkrevNWWusaYY/yYv08
Lux30h3y59W5oqOCIeurrFBp4CotabY2eKsAU5k1X4cVEJG8vYvWD1K6t9qUaahe
wVRf+EgrVigqylVTKt1fNd6NB1qtU+sQL/LYLdpbHYac/8RtSyzYCP/Oo/syqHVE
24+ygeqfo55mdkzUrEamYx4yjYZk7u3SgZ/CpCXqx5cb5Zq9Dwmvf3nU1prGc8ES
BLAfU7oDl2PznoogPISaDkHRqYDzzMb3m3JnEMQ+C50Y+Qr0qIlGtFGkxbWZynLY
0umUJM7JZk5o/ZUZ4ebfWAc1+m6bjckf4xIh9C3F42oeCmZG4SFsgZskkGs2BxTj
Z8zdDbUsLDP7URBDCz7hPtRegSH12QoR6pZ0NI7SR0L4AG5HnyRihVyQjSN7inqQ
pTqadSjQGgK7RD56sshBf5nFPkXrhByYBaFBjEaFwkhWzHxwQYFYUMWtmiycKuZz
7PFtitFmzZ0XADhrKuuPSlqG6sxlB16fo442WFvBC9XOBmq9Hp97k5f5iXKGu7lk
s1DBKKJsmCf09MTkNrhCbSlAJuAyaqK33cAXWHA6FQdohF0fft1fuNog5ml07XP7
yAm8P136/7lCiBBPfDjI2rUl6SkjxPt3Ct0r+SD77IYxbQt3cPzVvPXw3+OYNWL6
PF2atnX+x0FOQtbTf6nSJuZN1LdwTO2cNCT5FCRCA1GKuieQ4/y1D6UNsyMRdIgQ
Jli4NiL7Wnln0s5KO6X0M0K6+168bujaUhJNmefGs6D2nUe8zpb8WduQt6i/PgGB
rW0cPo/jot1MiApKRY7gV3XIICVOVRINn+7z5tYJrJstzvhWN0LCgLx2k+glkejj
qPf5At63H+b3RenDexl+t+dIDoTQUFp7kfhqQnQ1gY95AUhlCP9uBeYvEf8wYUSv
rJa6WTJ3wJsXkkD/vo+WPOeEzz74PK3snBqSQCRLXHd+hHfM2s2nBzibUz5cojeC
4pF64KQh+Y5Y7EIOrzo4D3krxdNETehUP6XgKg7RYvRQGTozzs2NSTeaK0ZBO59O
Rhjyt1NdkZIOc6vRPzStBcR9i7cYRCufyM4mwbCxuYlpK/wJq7ca7ffYoGhuLJUe
48kJBblYdRhllKXeEfkuR785THZtaZpg0p7GEuWWwVw76rTyOgvUUjmScLUiMMZg
EmmZLEPrGvzSuZ55vxp8ZU4tgNXMhrGQWCaX2pofQ/qqj/1NOvgYxPOCGPdJCgr9
+eSSGLJo93IYwY4rRNScGlV69PDo2QmwaTIpdCE9m1wit3eHfQgjeZCOqgvfZBTg
o1txrb37Z3OI38xZ7zhj34lm2xpekMOp0QIe+6679FXh7aG9QlI/0LPVlWn2RYx8
dJawXUzsvwHwjYtEq741rjhyHAg57jSUIcOonwqLRCZhNyD0lRM1UI6uIIxtcltL
y/WNa+6zLXndbZG1O4iQdTs7dUSYFhkOMsddYsLuLwuLJGZH0pfs+CTcvQob9aiX
ruNyokwwesJQ1WZoTxODWe7GlwxNVyvE0tmcCOk+6GTpuTNswWO5QGo2yEO3rKU9
VJ7hqZTb7Y0/PRjhrlhqlkvZpMcYtXtBxTXtERoriyGIgzBok35CpKGC5j6pzVa3
BMGtuWAI/p9KZNhnW5ubNzGSUhdhCycFs1kRdz3v6v0LvhLyxzZrVBlzPctzdWmh
I2NS/feAKMCSmt3IA4O5SP7mSa0+nWJlXwTN/Yu7PiRxjAKb+g951qsFnmzLpdIV
gy8HTfttvwfc2jJmBJJoYr7xN3mznx2Fm/oQNhuGw+0NbKby3LAEg4xslJoeExaq
opFY2tUC0O6dtEuCcD4S+hh7D4P2hjsGUQdkCZvUGbuAYpYfnItB5zs9QLdFZ990
XNqFCZOP8JkuPIrV23kEo6oDqMk3mI+L30Cku2lMrVltiEeSzNBqgf+Zsq1pczRC
ilPQGNWxIDpDxjUA4efqv3yJC060aQby25Z7uXxeLRcuvv1lxMzLVybVRuyJgyTT
HjodUJh22+VPx7zyZ5lwqTawJaKsT7PHgBq0sB3W0Z4rK2vpOftmWitXZnE215Os
9kwrqGlZ7E0enaZDI4yfs4e27wMppHW162reL9uuk1EEXbritAvAbQMURqgydiub
C97wf48wCJHr/b8eOwTZZ278QvGDvlJ497/XWmcXceXiYfC21PvJ3pwL8DYKr4ZB
7X62rmXhF0NY0WbCqp8bDk8/MZX9Y/7FFBhaU1m45FgP2X3bSlJf8qxWAEPc/3di
0b0kkE3FBLQvbXYwuQyvjwUn2nbJyHQeXRX7OFDrZH12C1gE0yX5R9wxP/WjnBif
FEqYU4tRuIKLhkCLvvZZKEUDPr5bq/sByzsHOe0GFMTLpHXTqJlpnwMdDcfrur3W
wa73ubGyBAfLlZG39TuVgxiJlemW10vv4tRRDZtgns4vrc7CMW/065pVxVfjbP8H
sQ5gJ5d8PVjZrdEDXMxDMoOmLU1flumK9WeeVGeCWUm647REyvdo/9cmVB9sqemF
b6m1WDsRSmhKuvj1kfaGfa/p/UapGT7gs1sLm5tFglu9fskCx0iqveYEpAQThPf+
ilY20BmQ1/IJdqJYgGDGrHt5Nej8/Rxyu419xGW+SSjkcsnCbpuhYAUcZQH6JX2u
4FfNSunGBWsPssMNfbxnUXldpaSxJxGWRX/AZKfnERxB+MJxOXFvrF5xIb7dZFjs
wM0XsEcHefDA1AGQLN9h1NXvQY8RgzQhIvdqgVnmQcW54M3X0U5DrgIz34PwuBT2
z1yu8Ft9P/3Dp6HaQat8FFeisySDnLorD9NVWaHvAiKqXeTxqOqmu5zIYvsTFYgE
efGs0xk0d8W6qrkGkNfGu9i3t81FCVpExZ+yR4wbL5oCY39PQljm2a5H2TOJbOyt
3tOmB5CJWK34rjA0L29a0KcUTMllyMlrGwmuPkQLZxX+yinrUzgDwQMajLykdrRJ
Ho5gPisNbdEnD4WKPtsfmEkWVu0aSEXWw5+g7csd19fzCDpz8r9n7U0fdHYa57m2
WZRmStEkTIZNx7o+hTBhUeK6lipoBO3NBbkHD8Xx/FCHQfEEpGlfb+e4S+9sAgkK
ZCQSTQU5bDHSv4oWzgtuv4oEc0G4AF/SiIV6S7ggqbm5ud+/BZhMrbJ0PgyPuN3Q
LjbpmXnJPfRrWbGRLtFspEiWK+6mT4WCklOhbCXEoBu7vXEf40kQTXc9AglUiY04
zwLhS79WLyh89/gjpS/veuuV1U4quxJ2yNTeyZubEqB1/VdLldS+2xUHHaTiwkHz
n6zFbEcIZ7gAq3refXz03xXtEIb/UvLG0jJTJXVSfG7WJAuPaPGbeTVjGWwwrlwZ
yNkOU6BkYzqHFQCq9rXDpyCj8ndUMyk3KlPzzzbOp2a77a32xDZUiqy9DI9k1t07
aX+VyC2bJOuO8lL0xS32Yw8ZsV4Fsj9TcKL1QCR4xNgzdOPP0/oly24G9rEfDU1k
JHLqJyPWh93y6WbLgr4/UuHi6PVhQ6rOsHrP9R1UA4ZnaUNWQBI0y1mp+IT/BshA
6ldIpjZzBSkCKOGdrYRyf1Y1hg9Vwh700+xjPZjQYyQkRiZwtmePUEXuSOzaYP4Y
sewkRx/jdhVIM4PuJHPwo1ENccRuPcLcjXncKIk77QyyJAFqEFoljIQQmyyAhveP
XEVFkomubs7/m+qdqJF7tU86wRa69MF2e4WoR+hgfhkpvsJuSnV8BEevnGLWQRVA
M38qsi48V+OcZamPP2cq2nTkgEIe77R7s3sQLKA6lW0Bk+aIp8b1/S842e9xnLMI
uRU9qTdILyEmq/yafxRHZra9v2cVMjUohKK072aGltag7moUONk86lMgikZK70pL
qlVbuzF5YOuiXNBc9IeivQuKfh9cZ60Za1zArXecbMsOddbD37xDtKpWRsM56BBH
/GFj0mJnH0eh4MukBxTFbCV9qNh2lavvbL2ehjF5u3e3WbjW3qYp/7r23uD6rDtZ
5a0m0D5McVJVF+JL0Ze9rT2lni31Zl+uh7HEugKKYT4vbqP5rGKwIc0aaMHdEbaE
CPxRAf6PQkpLcNSLYnYLy0PRhjOAYmoKdBqBqOHCOG+iYpEnDm3WWh+rXzi68FSq
lI+hqpLMgt5Pij+PnLCAa//6w2Tjz/ZYqsd14SibV8gteKUMRYjx1vg9YZ4HLVxe
cXdOIG+zWIqPCeyRAqN3K0OV8ck21cbhBXqSUFtSpqJcrT/UNcBa7QuWIf1aHgae
4xv6TDv5sX5KOf99MDtdCzI7dmFQowCvTX0c8xwRKwVOldmsx9koYwRihNFt+nEF
OUIsVQw3GhMtbLBXpUvQEpICixsxG7sNfmUtLRnKE88l39fnap48uO+O8OITpngc
/aeXirJr1VnDHXwI8nMSSWw8EV3Kg+2IMPkMou+m+fgwiHXRc4Vpa+/mCo3Q2HUQ
Xkc8KrgzofFwo7CHFcQLNX4S8d+VRmRVnX+ynGZ9zxY5w81OlcmADLZuTCVPv1Ll
vAbofsACl7nOyVApTztGap/1w6wZHXVewTbX+mY3x9ekTHQMIlFZ/CjQshJzQbPS
Pn3bQZygDj9hzvBbwGZss9Wh4E6WKSDxBcKYnayRuOT3ns7gC5a1cAMWtmubMkVK
r7/6nxGnIazB2iUcaaCIDrzazoy64jgjyc8FIfa9NAzMG6IhjljuokrZkzM1RvJI
qXEETIzakQfn0AkaZsNtxaJ1+SUNeMP/8wKZjqXBPdPMpUr9fj6ylBo7ccmjMJ0t
0lM6uLaaHkfdY0xodo3IkhjZuPmXj8VRe57r1QY6AeKpiIKtYSvWvbZShNjDNaIl
kOBF+FgzwmoYY4DDE9rmP/j64XWyZSJFqEKOCFb1dYdAFktC5OPAmMxeqqRq1t7L
SBCNHq2zhu2YONJfntovCzpd8eayESGZwhpaupa1oxeiIKU5NMGbtHRNCv+CoFUB
2i05pP8wk7aLieF8EZi8NPPG5Wii+iOFDc8YIb+/HhY4xjWC1YJO6B+L305LAA7E
SnSS5tU7WgHbepmTYwrhrkqoEhJIABJsmeiFz4tVVB1jUIVZKVNot4uLRm598ARx
KEuK1wAuSSu1HNKiVDrr6cbMspr8QGKztsz1fCXDjY+Gtvdgv/VzFwsJ3mosQkb5
ws9q54H5ajZGJKPILKh05VNH1n+XQGyVid8pk50oMovE6qZUrmLUHWMBkgmzVBER
ks15U4R1lhFOiu8gkzo3z02X96jxvLrlANHB4kZZdzexlaNPTU1ot8hDkUy/36Dc
y7z0oQ8lUWtP5QyB4JDQp3uo2sz+7OBrshgYcD+g/Auj+sWOlYjlxPfhWYR0PuvD
EViIBNXDFcQZMOSawRKMgIikbpjESrtbTKycpD37UI4WRMwtdGDU/jSfrk4dcXdx
QfBbO8Vf3PjA8ZKSV0aez7KnGFofMilDJw+CRdc+AAjN1hNYNLGaF/0/itZeWhYA
pg+xxqvo00dTogBhkOfHiXtZa8IWw3EthOUIka7J3Ffb6qX3HEPYt1TZKTGX7N2K
0Mtyjp1tYGKYzmerBYmcqNiWDPxr6kfv7mQA3h4tu6KaFhWx2Sw1Es5uGxWBJ1kP
0EG7JkSXp8z4B1iHZ8i+pt6Pd4H3iETAUUYWvoNh+sAMuvZC246uZIB4sdRFWNy6
x7bO+FFpm+ttSs2o/+NYVJ8lu8p8MP7yzrF5qpdq/w6LY6yWFzE4B2IJe36YDUEB
FuS87/zxd2WRtBZs4wLMP9FqZlxvr0TSRjdgZGWuFyiA7WCyFSc0o22sADggW8W3
ZPcZthvXVC4ZO/IXoWNqOk9cOjsmRkmlDz8eEepTPZdUb0CkW/bTPZQR9reIZWkK
SgKIaz/LcXnQUa34roQHZvsvQpHCyz2Z4hDLRE3paNxd+sSZcgCL4QohY36PogzJ
4712fCBWJvxyCKkFMnTfzKBu2m2p73aLCi1VL5BoDgYrxMYRNCIjTQiMuv3FhRg6
zxGuYaCSzLHlzrs/AT8jrnJ8BvQnHy5oCHmcR2Wq8quWzrg1LEK+CEHWRow0O1mU
EL1LGrDh5DTAfgbdtHUOk6dt7JUgS+3B6IVr60yGrTzQJl1U5aBF1acXVxWX/bua
Wt0+Fx0rnOrnxB19a3BOvCsfDLKF4H4RT5wOdtSn9zRezvSmZZD5m6Di7q8tAF+7
ALwwT1jecO6R5u42N/jj9kLqqfwNkx/9A4t9HNCWdCW10u+WpdvHMHip8ZmQYaBh
jriUSlGwjjdiPiyspqU3Br3QpO/EsLfjZ3Szncxpnfzojmwq8kewoD4BeJ2w52YI
+Aruh+jbtuONRw66RbFk4cUbBB3h2vQp1w2hjVYvQ5BU+2VHPmRnCenxpKuDA7RO
aL+U2y+xAZMYcK0EtB5Z1utcQgsNtbjs8kMzZo+LgiHqmmteLfNYmsEptkDWhpsN
QrR4QUFaa6PmyBQ6zs42y+M3fuc3H121msckIpEDlAaXCFiqgAO0yajh2XVis6cC
Pnh6tPXVoPtQ+zAeEpDw3fvgkhy37/VT+VrlA7oxxcaHcrcqUUIUfUuUPpBahiBt
MN+NyL+FzG1y40MzKGKXhXnS7A167aQe9ynl6gONFSNrfG2P7WzrJ2lT2yg4Hi0h
rK0izonZxxXh0dI96A9FkLzYZKHl1MBk3trdJSGNqyICT7wjoW03pnw22TfjcAi3
vnUDGNRX6NSlQE9I1v3OGzjc8ZANTr0tvsemDWmREvQfVi9LmflHDxDGvEO+pLtT
OwVYg55RG2hSvLIrBfZhJAtsi79bNoqXgxh4TWBE2jH5KIq6afmJxSgXw0yyw+ha
Q4Ww55Sa2sZpQiwwvIYiP6KhTZSFCKoehdNOw6xU44AX3wndE/giKcwfqmv9PqpU
bH4JjWiq5Fov1OwAavxRt4Vo1HWuXaIp4y6Y8N7Yt+nKMEg4uFBwakBxaAaf3m1R
YYl6iNcYGE9J+ozT+7S8Kc2PjfPaOPyzIQPTC988lW2n1Dvo07ItkF3NAxZBLz9C
Vtayjlds1eCTGrX7D6jOZj8m/CvgtqzLu4jg+vsYYCIFAPVEljVRY9H7WBzMu0GD
2U34sipd90xKiirYQzHl5/ISyEsVzuTPzDH8WYUZg2PH4cs8xu7SzoObmZIlkh8u
g9vUTghNzflyPdbi1jYf46g2Lw94Me25PeM9Eqw7Z8EM5GlhQ95wDMfX2UqD8LbS
dVbEkV0mSl6coPYAN8NVBZDh/XEEqt9bsbE2/HfKnQdOUMUAql0Me2GqVP3/pEFD
VBz1vtsWzKCHuM58yKDYXVgymKw+IB5n62RsPUlpnb3R2L4cDhquVukiJDlLA+VJ
NRIU6hRx82VX248Wa6xA6pPI03hIe0O8AgbDaAO0djTK7NQHWkexW0NLP0ZcDhhB
KgtTiN5T0kBSfoXnjLqk9goYLLBLHy7GBjwoQxV9yv6yADKMQ5ooJEArZ7nlETyd
D75scpYixVrrAETBf2qaHwPd01aQds8YRWz4l6CUn6fGMD8WuUGYxuBFg861sRh2
uQNn1xNCdq5PW4E3qLQQtjyBsW7p8gvp+ggrbx3ElnysP9VDtbWAXiNIEKGePkrQ
mizqSSDAI86mNCk2jTuihaKz9XtZXxfiMn3iQCd8aB9BzlvZ33ZjWBdkVM7vVA8A
L2lbZlkI770UmTilUwFD1r0Pg29/cv53jD4cZ3XvyXalTrVAxgvu2Mde//igRNzD
eNgpnXNfXehPvKr2cTUfij1WSzlMJeXNvR4FVqBdP1GcDyE/xVZuCXfCwyHxabFO
KT/LIUdLSQGSYD6sTAzKFw8zA3g09YUfLH/n9W3wxqhiOAtjf5Kxhgtn64LK2UFs
5uX2d+E+FCuPc6cvPN3oJfw7F/G2eS4+EHhrBDQlDHQ3kIwKy9GyQ8zrQ4cEultO
dxKNuvTxcNKA5bX4s2wSYxxU4EGbqEKLNe4d+q6dXDWYZfTSNKawDtpXjv3s5cCi
vbUkRCsdF7ru+f/i4hDzObqrSAqkKB0eZu8jqz7n9kOdC1WuSswt7UygDWIl/GAD
/rDX1IigvflVYX8LvZGI+kINMMvSf3DePqT6f2tKc5/QWQ3GxmUVJ257Q99Yr2Pr
NwjT6c84LdGMJj/+VkZKxVZTBTkAihbaU55q2vsZYfPIvyX1CHGM1gBJ9lkrHo84
OdACeEtOBKf9BYvqxG/9XbURynu/b1CxInzockU6avKoawI5XNraJh05rgl7xOee
N17Brj1kOF9rm5TuZhwr1ddRDpMNMTNu2aCkitVyyaxpc1MZC5HJgeJBEfzS3/W9
MAHbFMHymEf34PxXKxZIDuJ/YLIjh0SPBeLpVl5hm7k1z90vAM1X2xIzKnO8NvuW
q66ZbXCBmx5l5WWIj4h+MTr3cjAqwz+aGwj8erqxSm6itngaiwT04Q72VugqJILZ
Ar9qtzL8iM0gT52OFBA+OR7nh7O+EQei/3Q8HaV3dB2+/aqLCvtHprFbmJJ3eqHW
6BQ+Idtt1jUAyqMRpVCDwsnsyi8eMv7kxJjobbSgolQcBi0KImBL3rw1SvqxUvx0
lPva2bY3Sc2tfCQRD+0CYrVXs+YFTIsZ+nwTeWYmV8Vm248boWTDdMZkQgfXUQwp
ieqTyNnwtReG7ccLEGphl60RICsAbzCfGa7GZtZKNM4HQ/ICTP7RkHA6GkW8iYEq
2bEGWlukBWps9tmOBiUk3MZSYkR32cK5ly73l5cydUVIHYYw8MbaRoTHmsqPqmee
jwhNxobcAjcQKPTIPTBCOP/7BjWNAODF/r43E0gdSDmzQdlb0uVybnMh3RC0qg58
n0UG504n4KUrWwZQl1gwofYpqT0bjD6+Uted6DQFpadTokJcXL4iXVGM5FGzgbnu
GxIvsnpSa8oesgtuxH1ArNTz8yN4wGnr4K3wbZsCZNd9GHAPr/S2AidpVlM46CKO
jeCUMdE56nY+VGZqj7Ub+LRlp6x049SUAGnZYtdcy0uPSyYI8MMfzESVCvKnWhzY
A1RNHXXJFzuP0S9YPNZ0hsoUCQ183ON7X3RuKvKiUgk8DM0wvZvvSi6fdnfovhsd
JexuRDxl9BpL+EueGMU02YBz02zHMdOi8jb9ywBj26/B5ocFsItpRMsQ1deUHJxd
MZ2K3+x+TiP7lzCrkYXdj/feF7A5pV7dS2K5IzIwaN5CCltQdBA87vJPHrRJvwki
yJLCq3xGsDlyRDJMq2EFnT0XoqUf6UeY0w/BQPkQnVYqxDzEGjuMhYkpwZXz319y
gmpLyx5KdCcr4Ek9MiZ5Jl2ZtDtEreI10oZiZYJguWhzBNOFnUCpMHUBU7Cznl5R
F3DMfukkvo6rr7Yr499ckCGHyXo0ae+mZHWisDSU3rfpB05sHGjiQtD6EL/Ynll9
FC6CoOTNXlyzMDU1eyE15T3uTlpIHZfcdoFubn8BW/35peOu8LREO50U+WgUuUWj
bw6ZBSjDhyfn/MQJapzBc/wiZPUFbLICakSkD4I0cbhcGSZ0zFE5mJAX1yixCPS+
UhS7pX1kJJwzIQ4Skcw9sSo02iIsjg6HTRQtqtzXtcv7wvP60zcahrgUXIxfCeNG
BMOF2MVZ6bj/2m4qBWL+x0QeR9aA22r6wyyhcjCL376t1RA/BUZOiAs4EeDHhUfn
e0ni1QbCyzN2za/6p8KJ2MWvHPbqNqKA35vqq5eOhQUd1SvVdw3SH32FLTbRjNR2
5HSBmwYy6jjCyBm7610fjKz7Fzy3K9fZ5LGXYR4bEJiOC3Hs6QJUn/EvUjwT3k/N
mziSz37/bcAy3N5DpzUdqF8EiCJ4Yvdl6lQo6JRpP3XjLo0kSwx7TXVWQmbGorHQ
PSYWB60wsi8J42HqAR75mZrMApqChh+3RYl+oxta5/hSHrye9eEv1FzxFFKJ+8xp
0lHrcPVD5//NyeOV/JHf/A+lCuy+yHTh1her1oYYGf6AufCl1Lr53L/GIWkjMNr2
K0NA33Xfp5DlgyhpSA/W1AeYC7DzYZieFadsZ4vuN8mJJKcTztR1puH5ESf1IAm4
6/8XX+pFlkDEJO8IpTZeAsb2v2HCU0jvhXchqYFBgEUVcImwcFrPjKcAcA1UdpJ1
kuQ+de4E3xkrNhLkHhPWsFuO4OOBtomCUyjSpNOixZ5RGJjfDoR21ryrf7ASWYU9
3nkXxiFGytZ2PHRTG/97sO+kGwTJHZDgbxA8ssOh10QfPdSlz7ZVIpEEKV+RKH86
NKvAIJUc77B2hced5WJntvQYZKY5U/5qRFNGnOwfJuMhp0XtiC8QtrVXBOsFj3Xj
x+M/G8N/y36aUnVDBdzoz0WNt4yUUKsRZ1wXlU1+PZFNirC3PukK3/yllbjRp77t
eyhFvxcrSjnP4qF9owzAoXQiLe2LKp5XaLnksLRJy4Au2CyXt9LuwFtJhlC2FetF
54DNqPYfLsAcUv6Ug6cTUhrQx/+tEs1RS1EpLQVGsMXHehqbqe0BOVaDrLDp860x
rXhLKSynr0t0ZBTUcumoowwWBc1HsOW8ZJTB0qHCnxeCqPwGD5nGpxQ5QBv3te1W
ZHORt0z/Y0VB6mMvvvBsBOOtxadU3/g4QrdRs3qOWzaB3hKsuOT71PV8TketSXVj
TA6ZbFgW8QqrXVKpPVtJIRm0nC+omOPuD20y7kREbLhY337qHP0byp+fDq/m4YQV
teKw37B2dv/fTpaVqTcYubBwdDm84fx9E95NieC6+6taMW3IezvJ1rPoH2je9Put
1Q0QpuwpCO4GEtfgkTQ8Wy9sbpjj6eXAtPpgT/pMzOUkcocNoxjaaNu058lNzscg
X8qEAXHzgB2s1TQOJoOb+JYVxynFVFI+fyoAjYRznvk8XkOahWOPDHpUhykqENd6
3Iye3g/XG71u/GdupvpRYbHHy1fxDDxDdAOx0dVH7k32sdLriARylergxSHzWYY9
kdHxXJk5bz8YeetKg96KOeHMYo5ERLFzVS9oo+U8zdnBpiD21jv9pt8Ui2UV2rj9
wvAnN9bVc5uDPBpQfEhX2lOMpCHXnjWybpIYsOuDtBqfE7M363gNKNr3TVSVlXyb
kRIUZEZuUJRQlY98mx/147qoOaSKBLOoFMK1/OoFDjIshwEU0ru7TvdtX6qxlpXe
z3BV4QGRXwuxqFrtI9kgfyNjm1a9xEQ7ZqRCSLb9cnvrG31ZDjS8/UKHiw62suSc
cP11oEOOL9qpufzIHJteJ71vpAWUbe3dGbe79mDSJ7/tSVi5QBl8IW/2vrcSYW6S
ft6OyegebUXWI00P5E1Ow151IqT4d+a/ppWuVTmUMY9WaLFUr3nc7ZalILqfyoyF
GksjAXnPO0zi8FZZYiId27XItXolxD8SK3TaWBYV62YsfkljYU0jfjM4lzLOF8XS
CBzrSCUK6KKs6vKw/xpgZS3bRsxcrFC1JgqeXsJPhGeMe8TPwMhFaO8GBdYuD9bk
17iWseHe9Wn9ma0lYkvM52402lBD1BTmDR5FG2PkClJ52yeWNb0wc+nIPDto3+8Y
+9BlG/eAYCa1K56WRriJET/FUU3MeHIMYaEWSb0y2NJ45yXmB5Gu2ZP4hfWncsWW
GvWkuSHKG9hxOc2RLOv0kTDZRfRYxhcmypYDYdqCXulsDVrUe4yvuOpZQx2NVhlv
AKAmlGlWOD4gxZB19GOp8LV0hNrDa1vxRR524gDvr3UeBCq0BUgoTxTkytxr2exS
YozlWkWBW6RMpbuUAt4zxQXaSHyfXKqRBkLhLgweNrBbJ8uVBc6JNYVuowUSAnnd
a7vl7OaLkvxkiiLmEQxuE154KMNFFJGhz+wqPJsUhdaZ5vt42IzDub/rSp7nfC0J
G0D6oqog2OG1xJFIHu7BzRe2n6daHE4cqrhuT3363bfwrVi8nWre/a8iMm7ZvhDL
FdR5bjEVb2ue0XgjyJ+sNeVQ6JMxBefWLYQ6mW9a8G9XC3FjglhwBJWkO996F8Au
p0auV+Fi1n72OhtOsii4S+r0Mjkb4OM5uHPPzjHA9928++0FRlaieh4IbTvCiq3S
lRN/lGYXmfV8FjXTg+1OGmTRyLTOyEIUdA1Rf+095/pZ0ZVK2+apdaSBBuU5PkIV
A5bDBBbQF3BnNGbZ4MZlbb31yL880dRDxhz1uTUab7ZQ6OQFr5r86+OjP8CGzUr+
xsBWoqyBtYS7RXehoutcWmF16mRVM1VzU+Bl1wrIfFglMtk7vcAwhzPaTKgxvu3F
Vf+fVja1Q2Yag05doIyyGZ32SOwk3uvkBFlUpZKsszooa4rc1vDT2g3gm0fTZP+c
+zON9OWWWBj74MA4x1Di3v1JTIfmBPD9n8LqHpS3ED9gr9OACjRI+w6DWxLJs2HB
Y5r7FAoUcjkgreqgJp0/kuE+5zImiFxE3u37xMilsEzld9bbp5XEUn8XqcneRyZR
kr2Lr+Z5fpPsnBLwj8h7zGt7h7oef3SYlbAsoruluiBGy0gg9dAPdnmTezyYeajv
yaDr5zSJ/XUYWDlc11PpV0bShNXWeob1g6PlwdJ4gJk9sz+OMOXrbokrFtsI1JAi
ys8npyHK40+qE5uIn7z0ezfBF01ToQisvDd83XYc8Zc+Rrknozkd17z8FKwIdvCj
yIbKuYqY0eowHxjJS7CDblMD1fvfCTIqeLt3DpGNwdS7Cpov0CHl/I14acs1reG2
1wDdb6WIHc7eTryl0RNtBsWbD/D7jAuuqQnMHuPbIbO63qBRs9Cf9B6/kPhqSpRp
H4X8gJEf0M4xE3JRjdYHB04F3INlFKmfIjD5du+fpmIs2Pkqt1vuKYyTWef6jsq6
N6LXtHkuQGL1b1tdF8pzoMH01tvbcIUdz0fFRUKKwPWog1sJhcFfbnDcHOicWf3s
4w8GEWtE+aBaObktl7CoqhAknRqtyI89fTYHwDqQC4K5JU9pFXwbtmB+b+gKzoTq
AsKYprs6LI9ruwQXmXDcO/N1sqnLDRHZvaEFp8pE63RS/aPSg9wgScY/lo054Rmi
QxdF44MGxFjGwkNej8ZA53U/Ue9K/K5XmVqPTaJRjgom44EKFQOm80TnEvLD1cx9
7uVYnDZXWv/txy7TJFrxurQqcTW7PuwFaoWNfN2GLZ2f1B2CAAnLmW7y0QYUIr2q
1SxDa9uXoyxpwz8w0rKCLjR9mkV7QmrBCyToZL+Ovz5yj4gkJR1HdpZr87JWD336
+LSHU+Md9eeptbK7xJ6wjGztiZBvCjr+djo1QozCcsSkgcMiOvO1TVSolRYiOFHg
xnvORjReuCp8qx+dmEMXQvcx+mR67LUogoKxsfcJvXcd7pYnepGVRsRnZEVHmsJQ
H+BN4R6H5qsWfFaH5m2FHbSWDRenvgY+Kzn7MNo2t5UqShybSyc9qh+gdzfGQoTD
aGdaGZj6BduTcf/BxLGdezjffQ9ftHcWqWdehnKYjR+o7lcz/s34aIN3N/scZ8e4
yjgiFso7um8g0+cOGqGRdMQLyiVJvUnucTECctZGNToPoZu1mqrQoAtuOJM02sMn
PNpSbzeNZdYXkzpKIJ8UXDPK71ycvmuUrw7m2StkUZ/bIo3+5Hc+K/0lZ593yuBd
JtSw+D54LMdiLZLh3FHdYvKkjNol00QvvZnyS8AdnuwC++SAPZeGFOQb8x7QyuXD
IPAY0BRe81zOT5gdub8QwwnOkddiWMN236WxL1mMCPxArWLXVTZi9vREnQMOr9sl
+DRDtYP3cxlm7Y0XxrHjxTI9Nc1rlYyk/JSHtyiBQlHwEmYMpt05pIZ9csfTU+yY
j6YsQXGdOv9Eq5Y/MnPrKLp1uUuxZMQgU6KUDCygRIzPCPY91x/D/rj/MtxgDRO0
dml+OCFq2VOCnUsqwFpHKOuOAlcFLT7pzscdH2O9LCVzhIwQZkKPG2PeHU+AcpSR
fdZzL/7Hd+6uNflbDqzlRu/6Zyx8riqQBUeFVSbqFVoB2sFsRYlQKF3x3na5U02h
8VucwnhYTJgpcwbq4o4XbDPR5w/hhMC2KaH3GWyqKJHhFY1nuXOO1gVFR8BOhVld
RK5lKGZu/SpiDLOGBsu3RGOdKIRPcpyJzysC3P1n1XxaZllDTce5FEUnyli5XXYu
z3Fzw+sZjUjFj164jSEXHuvIIPMMXaSRvQaKNs4tR0olmmlpN5co5SzAXn6oMCCP
d+IOqq1Q2kmwDvROUhP8Jg5R+VH49LTSpowdJswXvg+j78eJY6mVNLT+pVB/GmLF
yK3x76OUFcpfEJMVBWzNdOERKLfpneUW2QSIFKZ+c2NQG9IDlw/CBYO6713HPxId
AyDHsXkhuvsU03VAXcuOZmc0Dysm91QAW87xEkhyqwJxP9Lw+S+is07TcpVika2l
0FVXIG20Ry/13/Y5FNdwE5eohsTngTy3tlPAOq0VibcpSxlSzGKhs2/Dt98Mps4x
7tdAkQdC1wkAPd/aZRpT6OFmIbsEDdy00Ch2P6MbwDujKM3FQf5oF7NakzCbsTsy
UhOSYrWYDOTMMAQRTPeuLRMYfJwwjG3DhCwkZ5KYkRmngfc+WnPg7PlZDAQM7MmI
bvUyAA2jsmx9RPPCtV1jdEqk3SIt/mxP26mz1ROUxKlc7VqL7hcN9T8mLChSDCHU
4c3zbX/0BuD4zoVLimJavcep+21I0QS38vvUrbC5aBkTq/Ew1G6f20Z/MqWeJ/Yd
/1B/uTSfe12bbUSdjwBgDMBIA+BvHE1Fh24M4jYGqNcawC6HMoVXhfNJ8Iw/6HUi
y0flR8Ch6GP2nJznBrvn455T5cQo7eBTuSJHrk1MQYIjhWpz4NlOZSjARwHb1jE3
Mu28Dz0xUuauqVpMQKAOLGomO4FWnKKbJKJzy6G8XxL7uzdA4xPTmRjHYbWx0DKE
dPln5jQKZSfWfpTXtM3iwcaU8ik9YXAaRyaIEvgyjBOvkE/8v4WhX/fL8OdslM8D
1+UvVxY748W/e146H9seSNv34TbM3XJB/c6wJGbTAPq/sWCSgaYRbICiB4XFwTu9
4pdsC5AU3ZwvREG5aOwl/vqXd7VVMXD8vydWZl5qtKe7NWqAJKQz/ckC84VspDyc
Gz4A5PgtQa9JRVXg4o7MEUde8qY208+bPzN8GuaYy6BhVzUnKzRUCOML/8Hqtxq6
Zs+2jgv40O5V9eGWyYJZicDbFxOlPby4bPXcHxbpbKjhZxsC5Xe5z2o6hkgWv7pb
kan30MebejMudmv1GeqEVp85pjjSs/GVLsyR2wQBiyObgmdfrhqwCHRqtNw5g2Cc
qozJscaKWmkD99rOGGEmw2/vhUCK3lLNs4HyxxBXEXZXNZGYt68YOJTr+EnJRdCd
6Tk9l5/E91B6wOJoPSQp1SzrjKjReH93+vFnEu8skr2tOdnIQm+cTyoquW85hdH8
LOf07DbnGgpVUCqZgh0te7ua6FxafyBRcmwRMwqDd/1Tj57TjhdExjPnxhe0w86T
vj8T5mnrTAUumNyxqlKRIXHCc2szokJOxfTALL+TWqgtgJw5VkVwblO966UObFVz
hDJ8z5udWuipKfTfaZP94X3lAwa0q1lqN5P4vAfh8ye2yON1eulLxU3G33UFIcpW
02T43wW1b8XZRRWI3qrE2ry8T2rcBbuNp/Ka+U6MNdK0+OTz4QrFPegl6XlD0BcC
54bnuTuOqDNZozwkQUZzMkk4BXx5EDL1G+jchmps6QyV0PqDjklp5BIlRGr/IE78
uZQHUJzY2WGjLlUN29AhKsZ+rxR2XevculoHMt6LBLei3PA3vSyTt4Y8eP8mZ17w
6ThNohadFRDEDnFY6lvF9yf+C+NWQYy6/znOiM2OmE1tj0Z5NP/vtwiDzizvXdck
f3WtQLEBAJtCOkE0a5qpoQs7DLi7yaG+pekpPS/JjzUuwnyUbfxD+4Q3U8RkBBuo
rO+3Psio9ESj11KEbC59KNcCPAZRdGBg8nsxzfa91qLDvQh1WCKadcgsjsVxAGdc
LTaiTB6mO5uv4nVtFNbLOaPK/mb7JdR1uRWRwzStYwRAs9cucc0NT4RFqcuo1E1U
4NM32lrfCbeaR//uHvYptUluoUp2RltlhtFsSePS3JqYX7HmFpHjkTer4LXkgcVa
Z+wIzaELi6cNqpzyMksbu/4BOnac7r0vNsFXzwAXwCAxK86CKVbGPf67JhrbtdBP
mWiS14Uh9N3spFh77m5RlN/nA/mcyX77Wa2WRMVrBaZKEAk3WbBIGwTHGVE4Onkn
xBPZLwf41hz38gqiSgB/tG+C3zUfpqNLDbdmoGV/mJZpunKys7XV297ryYriCA86
HqkmirWt+yBCTMQdvpMPP9l2BsIj1egUSCQNWz8nAbB3WiL8S9VrrjJqusIQopey
k1s5zSovRKAkRVV/EiWZu2ji9kixMuW72ttY6whmz+CPQp8D8LfxbmKcKUXMSjkq
+56D2et0kEgBg6wixxglEfp4oB6G0d4kH7LhZuLnkf+AfHD0NlnQhBX2D+Rsn83S
h70miTqrm9WWOTy8JZSRbf2xbJhzPBUHJlMhEfb45HEMF/HWAS/DmNguKhpBH9zT
ZcYJkU0FKeECWQtj80VSdI4k9TurHItaTUEd9gxK3FTM5JqKvCkgcW/0ZHUjb4Cj
EVjeoK4Wx/Br+RGzIwY4q5VGoK5ukXYz1Dj03BGFjxyQY/x9liddwtHjuu87JgDg
ZFYW8lhdQYKq3HFQXNBachujBJv6QUKQwg7FrzZUWhmPetwarY31m7fbBipzFU+v
AfU5AZDaio7aHwi5OKtdpib/BFSVMMPrM8t8Fd5rUqR70D1vA5yg2IZ5GXMeycsl
dMZGwIvy9CK6uidrDGrN1EVg27ur89/ioE5XdoovHJngNLfncL97C/Ri/GVBmV6V
pkHB7h/Bi5TT8PBHpMVsOo3EaMeaXTwpydvihN56WvZUzlpxDIFHKIL/fR5684wp
X5c0s4oKATA9PQO2y+QAn3MHpP3qcpYv30NmfFyVqtuHWlEHsZkIOMNEpO25MB1z
wB8twPx5gY9SEPLsVOslTGZbJqCW/BDvRW1Wyo7hy72jZ3KIbAMKkcBlP/BJrFHE
QwoTVbbxMMWict+lLPCPncBZk0SRX+XiGgzEzyJplY1mqAUxki/nVeuax5yGrmCq
k9NOA/8f0hpuk7x6wGKu8nMifNaXySeNp9OLQ+aacRKDw7pcsuFPHOU5bjU9y5mu
kXlReXpxmxex/PeX++TvU7gINHelzOIJ3CHo3dmxhogiNYQ11kE5C98AjKjjeHIM
GCly0EEXB68AX+1yiiMo+/MQaGyrBqzsYo348gj87HtbHWeGRW/sg5xpupcF+oKx
zvyPk1mO7LyknxJKsoOF4SSVzLDoko43z+0wTNC+6e6TdTiIIxLmW7dMSyEnJWMF
mJefedt7jUZnLxfKdVrLi2BaF5KvWoRqnbT9vVi4eGLn7lmZlT1BBSIk0PU2USJh
TmzTUiC1EX3GMqFl0jJM6fgrAigJERmHFEJF2sgFi8bZS1ZWHNOPXRY9/4NzlXNX
EZyEHGwlGVlBCPA4YpmiImES1XlDrPMzGFFML1LMxFsGroS9LyTMhKQ5fGfGhpiU
BYinJlQMndcLyth7u5IVKsVcpeij+DZisgPCS6t5HWCb1G0ru+dCFt5oO5kAfLnL
krQzQPEV8kLolRuuX/T7+/mJBclHww2q2HIsHsLKwGf1oaXKv6hYdOrsEumT6r1e
kbC7FnzAlhfAO6gu7EnolQYfzBmMI2UempytKYB5TpREFnW7vTgQ/S3AepmAe3tH
vWmb/pgsYZK5VpBSkzHd1vmIuJYias28HDN3T2b3J+vmekTDoZ9cWzVHPwo8t7uR
O6Agrjrxxlem2KNd6WHk5CmD/+SMtfroNgkdfMCkcZnCWieKvLk7UrEhIddmkR7l
GC0o4aZFpnx+etqN5/FOw8dOt4zqmV3mzN0WBPBlagY9dktxt41Z1poT0EE6Mz2D
HhOX+zQN+/Tfix3TKAmCGEOb/KxDj7BkHzmHU8sJRwd7RPRNI4gudMqI6VUOtsQ9
57g9uy1xtdE+cAqnhiRGgrus3Tr9erm4ocNuIrnfnel+N355WlTLl5C2DVUvdFgy
wEhDbrFAaLBIORJIGtsVNyEPtgZhUeYzG6uowCR50c5Zyy0Q4Cssy6A0txrVtNR5
94Je/HuewqO9WdqWUIeMBs4RH7gUlnoRHwIZrveWtuPXDHhoLIbNX6XARWVb/kYx
MkySqj6DTCfJdm/3y0Ba6k6CHKZDo1NiLd4qMnjANYtLr/h7ITTfMDR48z48Sjji
37BrnLJn5DBehpb4V315aUdChjmf9gJtCY4ZN/QwE63NpNLwZDpQ3+4Ytnrl+1i6
MEZ766TOps8S/Gz7eAqPBRI9vORpbrtTgM0yPJ58gzhMRuE7/nQxkn7jGOZIzqp8
B/o6ZP0FSh0TRFx9CHegiIOmt4G/lZBDHuL1NUiGYPAnyGrHF7dRUgE/NZOnS92a
2EjQ1gY4xNfDKULboPxwOI3yUWQONseq0vO7VzZif0AIyPcKEQeGmteWAah4Tj4V
c9AaqGRf3HvY4q0jqWotvRdBo+bdJkhl+eiKEjSyQr5mMIWTpBJsmWR+HH/irfVT
663fe1cYSg4lZjSpvwnfzG34Q5/aJ5cetiBzv1SgWXEi3RW2g5nV21t+9YpdNuqT
Bwz+WvMuHiRdQ+J+V6Qg39K68Z6CrHX3p8U9xklTpIWy8Ccn3Sw8IIsV2Xj42RXc
geArlxwHV0E7jnqNbizZoo8mGaoIyFwgfXLys2uGsAhO1I15XlzLyWAirYFZeUlQ
xswTHFjeyF3E73hXoeJImqA3hxnQQUBWN83umnPVuln32jVDXHNpQv2WYkSBMHAx
2iBq/Ko49CMAL0PdZ51zGu84dvtUZwudkA9oLDny0V4lqlftbTRdb01hymfuUgQx
afX5VnUB+0TIPjwNujYaq3Rso6xgCYQQplrVdgpetkDodwFeJWNZ2OcegTpSwojl
Cr3HWuiCn5574AdTIeUe8zgFOho01iL/DXNLnr+y/6ytghirlO5qY2RHeeIWSuSB
2qnBOEPnbCsjjraBYDCOif7CD6P+0zuI0Dodhg+OJr9LK/4w3tJH6Re8cpcv0mni
ifJzUGFX3URJ+fGv0QRBWGMZSzLfo502KdbYLAhIVxIQye9welB0CDPSOFPJhwXz
tj4Eh6wJIA9Kc4alvnnCOc5vSxKwfuNGzy7dQVGzoUX1jFKrvHXgWWWPj7r6eI0H
8igCrqv5h8NKCIMBl7u6RLZe/D3uIB1MmiKsIjbdLuJUB8kSwgCe9KwQuWw8duPy
EI7tc/hAjFEzwRBZwDBDS1Nq4OqNcmz5tzbivSNC3rnH+r7HxSO/sAg28KjT+/fx
FjTK81R384z/lN2n1m0u2PJzPhxGricMh+p118NgMYKi8MZypi6ArdOgkYp3LfQ2
fQXeEf1Sy+YeknGYS8Y1x0NuRkPV5qApURPbb7CF5uABwDxDcvgkiqqnVJNv3GAL
yfWQWPzMXDKrGEBrt8Vvrol7Tby1UR2m7UbdUFqTZNKaQ+nyRq7G8JyBra6S1Eej
eyqeJDTbsKhG7QHxYDBCJZwo2XPVmObLC40lYTiVr06xF0XnFEOqWPwsCJ+df2Ji
nkTUskRkE9NdcNtuPxSki67+vQEmzw+A6gyLDtqLHeGB8zrLU7yS9yXUeOkokgDj
Rvb/ip0TYG4Lm8e+KBMAR26YmP0C5/2xcEnnlKUsfkT+A/WjdOvAgZDs1C/XUMbC
OlR86m8tRGWqq2BRMToR6SgBZzZ0ZxwZuemBSXvLsKuWFSuiotbWWJVhJt6GxBqr
g9btaRTRhP2glZo8Dzm6MtBAFyJpDxlp623cMXtSdcUmKRGKk8QhOluBXRh0UwSP
HC9jGppuprjgZrT49efLYWDj9EdDLnLl2uImOZrIDDJNvo4kdx975BdvFQEzwPdA
xDro7bNGSHeVa7CjvMVSeBv1RykOQxV3D/xb2p2l1JHfY9SEWEwJY8WQWvIyNg4G
4g7XNFgAzxggm3ess5tjcm2PsflZOv12zmUZ3Gn6MSqvHG88COWD21PfSc6YOtUI
Xjng+TN0oE466J5XozGIZiJYpdogDIxw7qiEqfSFblKcvTgVFU6TD2aBatp2hNzz
gdBUhDNd2kNXRi/QIfA4jd9Izk3jf+hT22hoYI1eufhgxmOYoNjRR5zQtft1Lzpc
rEKbzxLWZLX+/bf+qtLyilud6v49fVU+zY9uIFPaFso/zLtLr80nnr/F8BeaeyZ7
9Kl5Tj3kIhY7G6nkFTlAD8ZCkfBpLmVYOnSyGECyV0uTRD9OlXvABnjJ9uZAfXF0
XlO2tfKwjMbFp6f3pJSMdBKZUyCdVYkkmuB9928KeK81nDYq9E5cX7lzHL1hEjGu
asAVOt+vSNsA/01DOzl38WCcquntc924QG81izQgBGzRRFuhwK1FKb8dKX5j40Il
YQoLU7iGqpUwh0xS4je5G5BIk6zOHjGZEok3wk/sganyLeRlrZCuxWpFIZgQYUS9
/bHgNSZVD1ahJI8JfXpSUuVFOE7Y/o5BYxINvmuME4irhOE1eHDv9bOH65yX5Rou
PibfxjkgLks9dEu056YG7Ko7MrENjmW8nlpHIVAAQ3+6pw3oMVFv199ORnJQaRTI
YWCI7dhqXFryAjd+AFeawe82GjZ0v+p6je38ccV/aFMwVWHR+U/rMWORSh0QCekP
tXFo/lFXA8XkWjDxFR6GAxS6jBvCWr/+I4EI6com7/OrbFnCAlvo2Zt0UIljgjIc
9Ddj92/3tjf+sD28iyRYs2mmAjazsYawms60xyFMMvfx4XhBZyjVnQfpaocOy5Q8
n2yAP+ZCC0/c2u/A//txsR6ABA1WEnutx0yKhZZI0bIyWFRHG4fyunw+we5l1qug
bB203hNjkzz+O/Q8maV18W0z08jRHFGgmLQjidOOJPxsHZStG9ozE9vuydTQxf7Q
RQR2exXykT4NCBNWrNJqZNF6QCOISuaz2ojatzi/Z0Z8Rwg8WrGDV0B6/r6MXP8P
cWyXO1IOb+UvPzTXe2wk52fOUz9+Ew6iP4AnvIrnrsjds4PvB17hExFkUCoFcuvm
9IAXDZCZ0Jx18My9dYGydGJ1BYwIiqcbfK8EFHnD+Py2g2srKuR5oef2jW1/10w1
WzL3DwVLg6YIl/VbUqtcc4qIQ4Mmce8I22fp2Br9LRwuR/ocdYi0w8iDD4UutEXv
vVroSph++86eM64tyXmVE87xtQ/rDBqi4P13wiXlTuCL+rT65gw65xbKqxOS1F6i
mc2RsT5paB+jGOOszfNkb+I3fRr2pR8LrtBYHrUU6tmzNfer4EmfkTYnz/fsKgWd
RqFw0U2Oly9LWEDp/DoyGObY5wG6p7aGmR4rBYO1WcI57nEqV8JQZDBpMo6J12Rc
pelxK/CiPxWpuT4iCQYMZVwbEYRWg8j1tCotnXsK9KuJSEKNDS/91Hdt+cADUZbk
uONKsuj4EVLUXi8jUK/9ZNOgIUzqFjlwu+qUr+IealDrPeJdEOv5XEribpyCw7w2
3X0PbbKIVKRp9PHUl9+BhNcKkU8UgNy68St0lPKonWEvh4nOSmKcNUeGFQUp932b
MiXU+MzaAxMIoEjaXTOWYZj3i4UjQIyLPYxhb9RcmYIAhXcRKNuWGuTUyjCK2Npg
SF89eqYwOeEvlE5A/ZPd2Bomo+UrEsHXocqI6UVQDXMtjOF7WS9rabM8W8x5SXcC
MaL4OyFnq3dxz+sU8YVR19V88kdJSnT64Pus6fBrc3biKCtM6DKJO7Ukz3M14nJb
IsLMet0GjZ3Xuts/hK6rXnZMcO5LcZZgnDaVjxdMFQMNnBIXFcWLbLj1WkhJeOpd
he8ESFC3Q1zoQMPkZXL1EVKZZZaMYkfWPbXvqYMy++32CnTkuLlMg2oLIjz1rAnZ
vPfaMsLzsHjSL3/h2LcUg0QnhNIcr/RaIv33PDVIAf2QRYReUv3bYJtVC2BpHtt4
g511weEA97CvkxnIkjl3ttaCgJl6TEzOt9hdGe5BihHjBVoOCASZJQ3xBDHpp/Qa
jdZWYvgIgkwDs+AyP0iwirD0bOdVFnElNkqsp3Hl/dn5aEoG5RhqB/uZXLcODgw4
ywaixdjDqJ7yuoDwPGC86Lm2Mk45nHb70a8wR+VKSiYfAG5XHzihy6ndpq3YoI4e
TejX+pF6+LbP7ta/fl57ZSEWnwtb860aWtU9HyFQ/uudHmnVKze4st5HjKwrszCc
b4QDTITtN0aVrQSIUkWbC+uJmeIxVQJsWILU/b5N+J84UDrhc34DBrOxlRlYVCYz
7+uEuqPSlD6y7+MVF7w99T175RVgB38WB0cznOn7c6igy2T2W4deEqVlT/msqrYF
XHLAiyBDQ1B7d4106gjBp0AXbNpxaxKwTh1yMjmB+gWB4fPhIg9ZZKZN/3VdDY5a
sqBIS8FcYw59jOGj6e6OdLw0nXFRuYNK2Wj+KS5NmYFwubgPjgqjCFuihYu8cKyM
5XLHzwxA/bGf2H7yu6xQd+AAb/IJP4wQHG5I4BPMjVzD47+Quzpi4uMcnW1NPJby
Qr9qmhkuoHILydCKl4oHWsVywNPhZYkaE0eiqN+5KmTxTRJOrfCQAdSALHWG0nb1
/Jd5TEB66MwOcKFoEQtAdRg+ZK5I3ZOpCi22gi7Y5qwCzBdS8TrJu0fSRbzzfRdo
8VSeE8XNC/772+HYd05lQmTxRqzgcpTnaPfRdayonhl+ABUBEVE8zj7NUMYYgAzt
6rPTSkXIOrux491QMg4T48cNOO3a14oiRFPloRP7SL52cQHOq/oTMkExCtNI5xNW
JqxcgpPUx4kSmV35L37uEJbyTT2Jy88FMbssFAIlmVqr+vk9rhcKvb/PNXOj+T9U
PSfb5RMqsAAc7y/LEgX14gKlagvx69sMbTiFSNVXjCuYbYkVrlaCt62XStysNkzC
ST+lFrhnrKxKBVMzujSQIZQzPOAPL9Rh9czQNUTZOAAPCcAiAYxMgqHAsTCNbSiW
wQBNcRUIKPRKWuUD20eEp9QBA7j1VIHKwCoHGjEQGdBp1NJE1KBWqyDqE6mPxF3/
JndpP57z3RKeOpvctiJzZ8Vz55hAxWodoobvd8JLrpLMgLsLJ/lua3nKs+0p5ZRi
sVUdwcKiCMvWfVeOCDFqYjur3iVIxs1xkmGKEQgAiI9IqhQ8PMJCWDbSY43jKVBy
JVJVm37oY6f15RwguSalYJNbu2IqK9T5EAfiomPk3fNqSR7s8iIPnRwaQvqvZQaC
RE0VCOIdfjG0VRC3CQJYayZrFNBKqXYmBWnPDxs+LE6dQ5S7W8T27Y0035gXdRXF
3eMnkWsT35qmlMJA02KzAhAAzZmeGmQ9DXWSWIqudv9ta0EESXUuCqaPNUIiM/FR
DLJ9UztquKWz/WL/QuT5/jPZPgJXGpzfYujiFSwBmzBjMaeMuzM6ooqz6Y/aeO61
MD+eHzjM28OzAXsh1DYs0n60ax14555l2Y9DVTD8hUmxHhI6e7l/2fU7mTsUuWFx
AYc3Ak/VRCsoHHWVyetxJ5vwIy5fyhB/xaKQbj0p80Ccczv/YLRRmq00F0BD+dwH
Qg3oaZOoX9Sy5/YVzXdubF1g3nj6h4uEGuX1lE1VsbeYK2ptPNsw1JSjB44gYiLk
Qf4kCsoaIZn9HFocOOd9Lb2Katj9YXjibrRd6lF8L1+BVetwNUhIN4NrHZC1QP2e
yI7X0reXJAdNqnO2FrI2pZ0AV4tAuj1p8P5zZbRo4ul/LF1DG93qB1+eFluxUW+t
EnWvVv1lqDIssGCqldeha8Wq8Cg/l9jbyK3pdvG4JKkY8nRKfMdEnIHgfe1OzK16
Q1G6dxvvC5YFJHtoWxrGi3ppB01I4vsTg4sF8s3WedrFOKTC8BKvhxZrCjsLJrGY
r40uP8nXsjlZ+FHil75LWuiI1LS8oja4nkVJBZBmSFV9D9/+hGVn9mFAuUiY7oN4
EPYWffANQMhnFVR9ZbI2yT37g2QvI7fZmDHM7uyPjVJh7kDVcGPMkHxF+CSVd2C0
X/YKQqmnLDrb73hbP7V7d4XkylhVHcGj5TH9jUSSLtxQ8q7qiNF1b0dwrUd8rynH
eqnrD+a+GJ28DJUHMf8Wbk0W1uylEbZYL3NidYympQfmedC9nbNtny4RztnGXoxz
gBah4T2V0EZm84JZLp6RTIM+QjMezrU/kUm9RcSdAN4CNQHRtnSf6+Oke4a8O9xW
Q+mieQu351c+61cTeu6v1DP+0OORaWn47iZvJPnfujTJlwMpiiKZGyTeGVDdkmIg
pK5mWT2LNYFT3Bq0Fl+pyZHxzKnKnrTtHnYyV8V7HRN73ze7QqHIn03N4Bb6QY58
5M0g6v2iVw0ci8qcLmTyGaN8RkeSqjioNz3Ak2rP4EiWq03jVI/Tl43G+SMMa4Nc
QKEO+MB6i98KU6U5YhYAzhf8oGY4i4ye17cyboH+yhZjd5LK+1ckdHISOmr7YFn7
8ppznq5hD4xzN2/iw1jbCKr8nRUiGnxEHy+govD2dhQeyIXJk4MRnlxlku3RWof6
zVs8fxy1fIzJHFpqvol4t8kO5UCGNKp+GUIocfHf965iehhmlJ+ByNUilnM9ALig
i4+ZeUzAHeXmKoy/QHDTwJRDMufLnoqSop6A7HT3PzT6qSE4E77DeBCi9DsfYs/o
FlINIg+bj+CaePLII6WxCojtzP3nvnXxla42AZqFQldPYO8hhvnPG6ivWHPbRA+6
FD3aX3R4YFfu8hLDlemifnKgvA+EAXsm9hIduR05qO5V0CSVsDHUq1geNY3iSUiv
56xX9QXA3LV8KGSjEGfRuR/jNJJbunmCHnqhTlzm9TmiO249TvcgDrKmevpi2jNa
WWdbDDZYRwVJPPGCfmnECVfGaEjsYAb36MjiN21sdoKFa4IEoN5z6KUNzRHGKsOX
URGiemsD0Ih8KyD008J58a/poLjW7ZSRb9Cw2tcwXzaFxAisI3d89bKVhlbmddzN
QDnhdRwU12aQ8wwsW9Kb7e6oCyHGNeQzGquOEQmap8kocBb6pnR7wi7KBzApwjno
3uzr9sTGTgZ4rFvnuYuuKTucf+Qhpp7S3vcZOU8fn6dqCV5IaXpy9JJVqH2JCf1q
JALrtEWOai3PADGf40gej2Pt3yzjK3C3OssAblTPhkmI1adVDNt3s/4lNCcFG1Xb
cHn/yL5K+7jkeJXkSiZp6b26vGcSAzK4thUSgjHK9jOKQj10bzEIMSY/iTZ/yE3q
WXfVJoUfQxnmtdmB3GWX6grZ+I5FOR4ikDLzu+ZjRyu2Iq44SoflsXBCHizWhiYQ
3cITiji74u0Hbeo4A7xiwLA9tTdBJULbkPX1gIJ6JVadPkL04Q45baxncowurBY/
bP3SKcE3jzdBgRwZZKRmLbIV6a0RACEw8IxIUEhzCpeVcw7pARcG6qmEKCVQHG6h
GDtptVJfOSFn+6qyK1Sca/omb3tLJ8BEQW1gUWqmJNRnyBV5wjgUBrBfRSEhD16W
onHu/46Fk04vcmc+VUOz6+R/krMX5+bwl4sbYaoaijnP8RXlv75B/iai8pDz69NB
MH2W7/wo6O7asFDDkw5r6ZHPF73axr/Ieoym4pWrDKeQ12x+JpU6HQtXH27hUO4V
eCUiHEt8BMTfDvcizi8OJv2qS3SbXHUjjCMw+Y1+syVeq6N5ptO3NzXxgjcFXqak
xzoqGWm/sfefF/I3dU7S+8zzpbudvpddMUqFq+uT/5U/3nWqkRxYdQi3LvU6Fzty
xe9DedxGyyXiKmFS7VEcmm+qiSHb1ltL65eNuJz6/gDVfMoDAIPb/IrgnRUPaoH1
llmKs+kwrRMPx+kVf7IUHCMImhZ4z1rkvbZgTL2gvA4gcR0uf36amIbGtMtnHT23
ueIarXSx5apB1N3uOAc+YJpSfxAUvpJN1TQWPtSX5RU+kMAXZ3LWEbe8HKGsTrGI
kH/BU5JcIrkQxNPyLKXRXuhBOPSC2nypu/csgSwLg45m7FdbtJ4BwrJCQRoIje4+
fR2Ocg/s3ryniFZf84Eo1nnsouG74KPQJh2jMCv2UaDGeqr6nZkizr8ZsHSD4dPQ
8eWPnc7hIWlm/rqjWliwSCte16yg+7/7Y+o1nWKsH3CZ7aKtIwBxU+rYtlG2Uaea
uXlb+cgYh4BuEL7tX/UJbmyR1vcowti8K8vQDRYOFUkj0aPaqnv4C6H6gB+kj39u
5D2islJmoUX8ODxoP0wKvLSqXCt98MZNvvqDxH3TvECJRs97AkHKQvcjgNp/lBL9
hORrte4nC0Q8w7Rp6BYtPr6xmxfjdMvri2kFpORkGoYxkyJHhIsFN91AI/gwkjXp
ZyhbFNpu/hFKEiswYFpPSkLLl/sR0r3ZWAC2+8YJxUgQ9DzPCw+yaj9ojECVhwub
ZgYd0VmSIjpfKBc/Oml5LpAmmUDCwT2RLI8JFeP6Ct3Gw4DU4DioSdZtahDqLlee
yFY/bBKMAz+uq/LdCNFxvgbRf35uBfgdiFGLz4Zmnk/HpJ92QjtIqP0gTfOgIMvX
YUFls0OcVFLqq01bMzDQNCsx0hcXDKurGdXXZy+AV3DXC+H5P4bzRIa7oTnGbw/j
KFg8R9C1pkyXWb9zqzmBH1hd6JqWgEelKOt70udmeQU6yfv6seLtd5K/cy7HQfM7
Mr0aHOm9ILKi/S0gWrj39ILJ9I0twr99uoJ1oNPK//0OuhJzZNDbNiY2d6pFoPaG
IOJHeF2FE+UNT+vqVJtqaLZZSu2WTdfR1CT6Wh6edqD0CofoB9PkVBX3V2HERyFu
c8pUouTftarPS050IGsOZVMeCHMGrn2ywcNnHQg+mIc5sO86tOLD0dKVW4w7Zrm0
nAHlMZE4DEf0OBmbGAZmmYajlif0WySCAXqL3Y3rQyaUQO+obD+f5wdMQ5CFUj/5
9vBODduPVqozCGmf0IxdDSVRVGcZuQoDDszfWGZ1lTXEfw1zxj7ni2YR7DRhTfjv
A+P89THVEziqZZDcb6fcV4TbX186Od0wE9O58XGx5T2gcNJ8MEOywCUvZTeuN9Sh
v8/JYHHZ6aPT1PLXamGfBJ+5azKVNBwls7n9DNf7NpsGYB1o9iDHBc/FbR7r5dEs
m3mRvstmPdLTyU7e6+fFfpcSM59k38ulO/QuhOx9xvDvlYAK3P/koG98tqXtc58c
0uUHIaoLEiX+yAlUYzYz1ySMXY+SW3L9pwzfbGzzs68y+ruPmU9jicYztd9mLn97
bA9HZrBSLebJLtCh7CbMVOAPKmqnQWNwgqbFi8ps0227P8h5YCkbqIG6wLlXTf+8
nVRMzstuYdNUPT096m0g+0ZbyQ2cDdzLSppQqSkUpKeM25fe5jKRirfyLYZH/+62
v3k84UV5v0UmDeu6VCpgPdMfmAMJHgj0JSoKHEvqg8dD4jbPTDanpbDlrZJLX1Re
S9GGuCKW8URLIlEw8f8yIJQ6xVVCsfWmMzVlUyag6Uz+OdG4ISBSV0qHuG6eOWaC
l2r7niBICz5Xtp098xOsxY3Zh9CHaHFbJon6XiTkt1iBpRmX7Vt0ajXP3pWAM9Rl
K8IKyys/tr3qjsTfRmigrAe5Le0+Ie/nU5aS+O+fbadjeW9DA4EeRuxVQlP+2SOt
4eyYlRygScqDmvlM2OraIGo+T7ULLSqe8uE2BrCvDx21hZx4nzp6nqqmMkbOBJja
bvSP3ftnPpRbq1KNC3xEgjSmqJwVShp8uXRBOx/RW7q1dJHXpMgMxTxZIDxxA90w
CxcGik12CUolBUoJli10VyReG18IRJ88N/ez/KcaHVnQ66Wwg870fhVS5q5c99B2
Lioa/onUJscTEeOyDjjrXCBovDhoYnOtQBUuc3NAPKdY/h6esYkTHjKF2FpAFvs8
xRa2jvXHVzh85uagm/CFzabrOixXz2Y3vinj8nxiNYklM9JLJSTzDKoKbzNmpJM1
s4Udew0JdK8jbVcu5ukMrZfMqsR3M/+9CSqZgugIyTNWclg8GNA0JOOBzengaOhM
xmdz347OuvTRtHUPEFhuNh2eOunv8ul1h8A+L/v0aojRhDJdBk37bnt/QPdNff8x
GTBbNGW5E9NzjgAP+9vCaQhYviE/Eq9MF/iA5D0MfBV33sb/24VrbSrvMarxHgLt
56Zt9GzGNaDE1TGKoloGU1MdVXJ5mA31HmCafY2egUhfz1gUc2gqvOXBnHgpGs8B
YMBFRNXzJqSITqyvZPWu7Gtq5L2q78VnLuREXArVatCcvp4i63nHr9E1DizkLQ6U
DiQYytQw9PAvZGzJJCvqLD6OpNo6P0eZob483OgI+lURlqMdU67XMx1Xe7wvFA6x
2Ic34XhY74j722yB2+nsr9s/8sQLakRbkUavazpsZcU0AndacDpqCP3yXligJPEa
gtExVRAtozUO8DApCDGNlqD+6vnCpzS4dmaO2fi9Uf9xZkeIUDt9mZLTTSxKKOxi
vD7K6Fgy+Q0bj4UlnsYlBL7qBScFpObsy167kMS7OmljEwSMUMCRdmf7kMAK5vio
V9a5y7qbO7fPjFodG/Y61uubjSghcJMO28Yb+iXJCJUL5eKhOuEDeFNslMiq6khs
gb8LRnydd+pl8EHK0Jmzra8+alxZMVKbPTQc3U2dY0MxVm+E0FtTwktb3uEzNM76
tHw0FC5Y3sTWyWE76bU7blQnkQUhWqoe0Y1MrsRq2D/+RzUEfkwQDKaLaMnklmo7
raEPokSPoLvH8UVweR/fC78lRlEWsiwZepDWSFPkGPXkDVE7vyduied4ttWlHaUp
RVR8NCAAyKqjXsmEQOXoETSD2nCcfKMdtUWTiPU1YlVt3Tvx9mrfZSRBffD6gBjN
tTPK2Zv0GrIupu3k7KjMBpj7Aa15X2sxYtiRrfzE+F2zUeIsLJHoyuRSyKAJ1wj1
LSegBoFZcY5veH8AgWFRXtOYWsziOyhCZdzeYvyBmojFyk/kQ0fMItHQz/pM/nqH
mSQ+tUWgMKzwh1x4nl7PRPN1NRLc09+n5/hnsIxFeZ2GJLRfNBdKL868EfA1NGx2
0KDqxeAHb6CWieUpBmRrDl0cDE0E0ocxdG3KZCRtwJVENPdNneZcTsuQ6qkNlL6q
Yu6gXOFMjTwV94wQjMLrwDk4c0pXcMYu9Nl2m7E1J9L/C2xJ1dIBS0knjyA0Cq1v
HZmz8LXxo7M//9cAFkomV6mNc0EDL4b3mWplN4EfFGSh7zOYIFuji5AXCvigl5O5
XhUPjZV0YRg4lmLb4a0vUbUjtqeGC3NT/jv8j9kl07Ams3CEntbFnj/xhlc0u0QS
N2gEOzOeE2Cxo9Mky9VXUNVM9JYbmXxLRozO1e4K/OLiT3QQwfCZK+239Q+8yvEN
T7K/FI9L6SQyiVKPp5eBVpcis+8X7lCnrGt5kdWV6NAFs3sDMb97rDj6sMv5ExPR
tJ1cweJg6/Qzhje1y9QKIFUxFayzJVnOS4tY7PXYwBSmm0738OAjI3N7ha8ohvKd
ge0NaECGOVey2/HuPr4qRQhWOLG4I4pM6iiTwzIBXepzT51CSd016+5xnpWahlL1
I2WYIWEEaj/oCYCNNeAMhDgT3noVzSLmFbV40Q+Jpqn1CMFnCmlqLy3GpC7tqceY
ermb7V/vFdoIej2RyHsHEyg2i1LcHzf24zc/RTQ/ehq6V0Sk3gExs/xa8m6dhUx8
QxjCZ+7RrdBcBDs7MbV/RsPqplWRwPkdicraFxJD961kDzH/ATDhxRyE2IYW0hHO
vHqSTP3bfgH543ErAhzQk8ZBNApOhkIULBmDotxIoz4aJY7p7tk5nDJxtFqv79rd
j19/a90HmdxWxVHKV5I5+KY1agVpkF/pDpC1XCxOe4FhwHHPrlHwv//6vYfHiThU
qJ1xu2PNAZwNVUv8Y35o9GD0Gb7vbosKOxODKmZaDzx943vFvVzYRG37HA6U6Zx9
yUPA1YnHErfzp9ppP9sdt7ubC3+M4y2R4r9aBBqgENvePHHMX2TcN6b1I1wOEhyu
bv7fxX0Xy7U1gQ/RlU5ndfHfZx6wcU2PIm8Qr6QYzcs87C8G425A5oOEuoZLlWdi
zTprWlMQOKk8M0PMSiEQzqbs8IJjrHusctVE2HoOCnEoH/hFwBjgfmmjxDThBXI6
UGf/+w058KnWYx9uYYLpwEiLMRiwm5CYK+W8OSFqCW/erG2323Il1I9eDjyxicnN
qHXX0Eor8UFruAc1im0ZW7IlfS4Nr4rX7rS2cz9PsF57wZrgg/1IagoTAV4ypafH
Gyx4ckOhhiw2az+VURF2VsekJPClDbuaRjQ7OG82MnGIj5oskxw0+JyFraxvVA7H
LkVG3Fox/tyAavrHPbVhoOq4RSMsYRsIWz0tSTLBbWexyk5QKX5jsiWo2sw83nyd
gu5RoMlXQSrj8PoCYQMhMyRc8fQgvA4bTXOXI4dnmBDWvg3OhQ+HquzF2L71aldC
ELxflWUSHNn6PaRENx/6uZ8slpK/xZbu/RbFt9+KBJciX0VXcWlvYlw2VDqAHgiS
uPDh+nrLsikt0kajQC3S5fFyRblD/1Bjo+sVqN+lrwDYQo3h8vq0iyci3Wh3wcXA
OjJ24DLWJ7c26V+Lj0KmZL7eovzAnm3e9LAJHPEMABEozLQPCFcDefgCONe7okE2
aiyJ5A/qjy+qdPPVV6u9Y9CQU4RVPnOMOZb/7SxgdERdjC+n1fEq76t9Q45a938t
Oyhn78JzJiRuOyeBrrWhRurGgKqHZ9TfV0t+8TwS676mt/GNmh/5FYOlUuqnF41F
QPf7o0KDVgc6pLhNBSjC+DCVCFKYGlukCiZfmp+aoosBgW4N2akZ8z+h5qsYRzzx
G+qZjn93p06sWPedUeQ3ZUrMNi5uakrnfF80np4hi/chYhCGHFh8bDVnht6xBYcu
F04VeknNlaDN/4kkPyWth5o0BlSsmbqXeY8ALjKcfGoTS+nDsEZ0eS7E6Cc6y/AP
nRlsXAdcgotac1e8+sW36kUFvhrTmCfQwuXfKNi2A7PMs5olZU7n6xhKI83IzzQZ
ztJ0cGexRtjNAuzZ1+pzrn+fUndZ1gR0+d2WIqhEJv4w+o5rF1IAIANFoUIujYUa
HtX5O0j3iU+mmEmaiWUTS8VBMlLy0bTR3Ob4ts+S/Xtn/8pItewNjSB7g9zPRWTb
zKgjV+N+cwxrygHjTszCKL5TuVUmp/BQxbOMJZhJYEMQJYpA3lUMubGQdmGizCJk
t1Wvst3bc+rjVX2LjMp7o02Q+pQLkGXhhq/n4DLV/4CNX9gjqZF0kATmYrjQN8eB
s1D5rabDPfEnRk1LXdTwCPa6p7k47CyucX2HhGvs1XKsi4F0TnvNnFchgImWlDM7
F/eTNBcE+IfsmNwwqN/wu7bNDspeOJ6AyOa3IUgHeXvOGubrluxyVym8/mrPUrTS
v7y6lylzW6skFO72uTNeY/w+tvH4+kdgkGX2V5eR4Gal0GObTrf3t57So5HaxFD4
Enwf+vS47W437q0Jlpig93l52oBnrrCQ9He9FkBwDOsSQ5m9QxsNhZgGZ42omlFJ
biNgzy1aMuiD5JJzL6iAZ3tMYjqFeAAn2XpB3juO9T8u+7UPIgRLYoz2VSV04hTX
DNvjSFjBB/v23Y1XoGE9gCf2rBoLjfO9H5XGNToM7FMVm4njKG4gCatmrMdUvNQR
bdn3rl7RNwQYjC30gZvflFg8oJOVgOMXZJbi4RQRjAKFGq32w/uyquJ3UpXBeEfb
HhrTQs5bccTfHthoOvBqK0P8qnwkDbavDrYEZYRPw7PGUdmg1Ha0IXjgFOcKnhW6
Zhokd/Dq8Am8uT2J8DijqTR7DrDZEkF6pkjWzWTXl0kPCtI86d84QYAqsnG1VSWv
cnWU2Mzk4uoTN8X0KFevgcJtZc14RjhfAm8gyit59kw2/6jIU5geFc5Xn3z6Dtlj
7zyWt+un6kHNPx25en1pIV9A+vE9pzjfe1Y6+sEcdsl3HPii/kI3bRApTqMRo+v8
cGV3d5cPygcKXBDZCHxXp+XMsG8UILrNf+b7fmyq7DOMnZxOHKHEPW0wsISBbLz+
CZOXEd+lnEZY/BfcfYNgJ1++PUkt8mVZBMTX8z8W0CvzQtFr/l10T9AmdXklJKHM
JDUg3vhHz8Y+LYRyunCkb3RASykBro51qoIPa8mSJKHQOORCqArW5gNbVOUXFqIr
TZO2cwLqeBGMsKN5FVnMvia6d48pzAAtHNZ9rkl9Nc2/RRGipaLzQfTj/X8yX+nr
ZmFd3c5Z6Y823OsUAScJvieyUHsjKe1FrTv583ADBFRBF9LvltW4GpESN8z6GTRo
ItLcfe1He5GAFQwqAtJaGSl2jXV0y8JG0UW/vGMr64Hw8LHH8uKJTTbAA94uv3fA
ewbwKPCYVz6QjVwoIlBJ9TdBxlTpmKUsTLiKS9hgV/83S6+G/aDPL0bIZNeU29r+
ImtPGPpMXnxVYPwunE4+21WsBu0e6nawInwlDZrHNjgar450ndyXJL4qMIFaAx6r
RtPvbyqhk/9XaVqJR7GSmx8BX0oiKSpXSohD2ca2I3yU5xmQjScNe+rcPiunX0EZ
PmGO0ZezQiwqsp1wwL3+iB+9bLIdxbJMpSJx0pk2MLy9EwrBeT6d8jJLFEMRAMYF
volDwbDRjDH+9vosceyhOz/x/HyW5A9A2xXAiP6sDwLYB/KAvqpS06kUPRtvPiqi
r56dlOKPvUph439MYc+Tn44LZTmh9uw9ymyuHqKxj3tZCjebN0J+rJIawIPQIxNs
6MxJROp2aWGCeCmeRwdoC3cBUW9oaM4Euip28/oHfYxHttkKSH8/3I7OeolM8BmH
myQEdqFK8uyXEO88L96HAUs08TWDAMC5/WIsbW9aJrkIJJbKRdkW+3/sXyZexcHn
oFzzRS1+c5kFD30mhsXaKl0a6zWr8nPjRxMrRg07h7YHziBc2yDAZJ8f3rX75XAM
PtvCBwz5pUB0GjaOgxMnmXW9M5PoD3x8zVuLq4PgLBjskv2O/gHeNW1tz0TOh/uN
T0zl1kbgStiijf30ZTupSpA4tDDejjR8r60jFYFc0DLZgB4al60swrCG4YwSV3lI
ck1LE+O5S6v23bSfVjoUJGsQGGJNpK/EhHOBk19sZH35XYVsjyTtftbtOQT13Szd
RrP6AIs0UWqtRRmxz+EA+UcRLAkoqUk2Jj3Hz6aFZEQE0KlgjsLPVgCzo/loqKpO
l8eN/ELhRBbrDIJCPhcR92n2B2/ZzKD7KCd7S6AZGV7EtyDIyoxxQ56PAzCfupQM
b+/4B4Z2M7re/HMA5TDV0wnWMBAZrIHZBpjuQzGkslM2xAZX5H8ism6bWMsldAci
3MNM4BOrocQMAVWUm4h0FnjO9zC9kFzFKbEii33DD5GaeNSUTCGVJfFl3/4mecEI
woRxD3io7xPjnheVXrT6RsbrsPlRAUacANri/DUQGu2lg1PiDYsWf170QZqBBfoF
pVayCGLc/8lop22ctG7oYoCvs0T96v7jmvcbwTMNkjwl33DdOllGmDoDC0Zddrjh
IGpGN+nBSYnxeEAoiJJHRgU7ydd8+JuHbM2W1r5cGoI3k+m4AM/NqGLATdeI7ffd
adEIHv9fCCBSHG6VwK2GdfBSlM1pdo71RUDaiObBOJdoAktRhSfBR9KyWRCvmewj
KNb7totTNGmzr5Zn+PyO6Ob5FvgG6CygfZC1WDrA5EYY/G/d/mQzsN5MWB3Q2C2i
0Fp9rZIH992HJIXXIBaN1rMOURbxQp1WwI34pUPX5mVqi1w6bjxPdv2dlwPX/7nl
wEbY2dI+A4RKNKiZwsMTMp1GM/uvKHtVxMEGKw/XUdL2ApHLdOXDPFeuQXUn50rn
dr2IlH30EIAzry2tEMfkESbV5d0xM5G6ilIurwJr/gC/fx8Bf+VlqgR7P0z4PvXb
A1NZcyhoa/yJNrD2RzV9YmKVrO845wo1g+ZNKC6F6z15c9JkKB1qdpZbTUGGcw6k
d5plLYKhCDqLgsqB4MxHigsPsG8GGKZ8Tmyp7GqBhMHV+CJAZxAplahCqd+0/q69
rHQOam59FqsP8PKxVIuSxxmOAxsQwhLwvzzFig6wpr9kwm6wPJm54wFbXzYZgpGE
1ouY720dqccN/K9NSw4bMtOlC6CmcwTf1u7AxxUdLIC9zAk8qcBODNw+o6VLJfNb
NUg3r7Wj7zTF8PbyiB+gQqEe2Krtaiz3/EDgSkW035E6dVi0jgO/jBkp6o2o2PGb
UGAaTz0RehiXYuuHZJTdISqF/mgnFj1CE6rXmuo6pwK6c5qnR19+LtF9NBzvJVoo
sGnekxsLhL4F0PBTXFPbcsHjA6d7lk62FEdhv7mRnbkm7fwXjLbYekhxEpHcArf5
Fu/IhZ3wBxf1TbUQqH7IsIlir6WuOJ2GLrvPSPXlIgp3qy0QK1LA2ABWsOCI15W1
zLR36DZEXuAsbkqqfA4pX1/OlHkvD8OAAw1qrO3GlOSFX5pauP39/GNzDK5baXrR
dQMga8xWxV949BtTWnL/bTx2Z5nUl43D5qLR50N6PZaO1+gdEimi2nmvCKpB5j3l
v9zPmSZLPw755c3g6imqNnOvuFx/k+BCV/GIoM6fR3wuL3TaVzQTf0Bg/iudtXnQ
8Kbo2i1H0aTJEMLAMuMid9hMoqmy0hiA19QECFMyOJs9preWBg4e9XyP0oU9LzmX
/cY8WlHMy2timkeqh5PBcdgaNCLo2GDMTjaN5TgV6oLJIYH8a+hawyOgt17fm2yj
fGPAMU/eNcL9fn5AiL45gXEVc1TSAiCVjwIUTXtJif/SsbZXb6K5q+Y3K2Q6SJd0
aDOFHw9Rgb+mPLng8WmesBQbW/eEceigW1f3VVVow7TsNKOvS3cAIVIBs1NYo1ZZ
OtyMP4Tlkokp5050eb/Dovq1ox4n/+tAT0T50kxvZOlkgddX0k5CZfqAooJR/Dtp
iOwRC1/IuleTrUsnFPvkNwCQBbSGMKpVHKg3zsUCszSrP4AicR4uZzk9rEst9aVf
uV7gov6ljQBHwBTTRNo2dBbpgF/2WMzUFttk2gKVrKJHHF53iYsDFn02WT+8z37A
Wca2EPhSe5r3KRvxVqwjncaHtDNU9UTwqktBuFSDr2qiMTDYoogjQPhGQW65arg2
6B/efbbt5Fi2Ls1ryP/D9FqwYzvaUWVU2HqQG72Em/J/KV4fWU7kp1z76Dh/pR5o
u+Do++lNyIbfFNcN/kVrEidMustAQkx1tiZMJsYTrvy8AsIP3izTcpj8/GVs6x5a
bNmdlTkbH4jd2HSwzHVG0xVEu1znDzvVe6bfFWYVP0E9scdH5kzW7D2MFSqgzAt0
HKL4JYWAJm5P4553//0HTnFMrfNe15fkE18oUdVIjGEZDtiRSml84Ai3mNIiUJPu
U8HJZW7lbokWjy/9MA5QXo9wn6RzRQouIhb9eUV11LSvHH1ZIBud9eMNH2CEctgr
RLfwwErL0pNEXkq8P4wDcqiW430TJjYv10RJtldpaL8zDztCMgzeMBGUM5A2TT5A
9ZDrdb6kqW+9vQEtKac2/1FAu9wWjdamc9Hvl9Ns270V83inlHzanJ6ojN83QQnq
rZPDts6AiGO1rwp4+DVQSy3cKr17/dwSxy/PhsYuWfVtQvhQFQh+7soKYe7Ysnnw
a6fiimY5gke56zKkkh3+agKFWu5AnKGh2yOUhOdE/2TY1GX7R6r7TuSy1y+BVtsM
nsyfLptrRJ63g2V2waf1VElok5Kb1D/dlxWsnacD9X4vCcRfoUYLlq3p0hlEgwbb
R/ty/obRrcHmpB3Ojn+iwO02DBm8lQhmdX9gPIPbF2mR87OT1NY0FO2P/4px0ixQ
k4Sv5JYYT6HPOtejztuiGeODK+7Y2b2T21NsuPsiTMyLdtc9lznNSkT7dnTFe1fr
p5VHvVglcYRWXV84ivzCzXPS5gbNcYLd36cIJXMUEkcsq4RndtTcFRUR+bzXETrP
8nyaUK8+ZFKcK39XqaoimoxiP1Ia4xVrGgwhCpemu+kc6eewirq/9gkJx27+FChr
cAuu+yCHwX8CGhk43WmIcQk+KrNvjyS+QlYTm21mog6o/sunjdL3SJ3fu9C4sv8E
AGsHpGAMCmY0oxqQKHVYrVFxD/snqrahlB+fM8D6sae0yvhcWKhbWbhiPMNeX+HB
LdIbZQICoCZ/o9AjmuzDsyXxcnjAxYxqALifhDl//qZplWKvRU9jk5Jhk1C3D084
VYYURJgh/0aybBJwQvk3in0Vfh4RHWAKlPa8U4lejXCUWJjaHhIsNTD9h4TNm+zI
gj6/Gh9Hn1ohGBemXNUEdVCc6pYRaXOtancGTKHU8IXjGd8ZkcBBIZMecf/gcaTR
IK0Mvldpnff83gRNZ7NFJBFYuTTUq4F+8M1ZGxlWNdDSmuMCMNp4t7hXYJQ1WxGn
mbTgMb30Zt6HZV/fZzboEWo+pFjrbRYvMeeEC/rUT41inMrWUEwZS7cEBkMMaPjE
2xgUpIVH7E3gx9YSoC9u2psdmi06Vay8PENQayMBUzOaME++oTNF3Ho6MATV7vqQ
TgsRQF2bPWjBRsnHH6JvCXT2rTUk0L2+yr9jSWYrtYweF0hNgTHpbR8Htqh0cNY2
Q948DvrR5wpfhkoF2ptqE3xvz13rymHZkwoyp6bNBSVmoZf6wClx9q+WzY/cKS9A
/fXCIUNNfH3ldvv1M9aWzQOpN4xWiq5x2OBtWre/OlrdUfajFqOzf+5vc/lbMKEr
HLAaL7g40jysS7iCYN6d83DyMNVwk23DM6NEur+j5bQwEMHvjLfjHQvzhwvltDtb
sI+pDXtwh86A0FykYhh6e4UIqoCw4holr5H9cIMHY5jzrpqwI3mXFbqoarJxD5mZ
dE0c0rsqf7upeHDdjrili6SIruLnI662LoT8PCY5WkQM8hf7gnUb/x4aK+3HrPZ5
CEhna7uGiU5qDJl09mNKKWmLIA+ecPbodPSF2lyJKY9xhWi2Wsz3r3ZOBy+CpjNP
BM17IBvjfU2T1oHxHfGnOupQjiBNQxRhB+7M/oXIEddxRQjOjLMQ3+b85FalI/tw
ctC8ZEOAVN1UPh7m6A1rjmfn6J4e2tvt6Ap5tT9wGWN++Cs6dUXcB+KY2g7WnWzr
FP/OLQeICbALKEO+F9ETjwRlw9yZldzC1M+Biukt4BC52l/ulU1G7M9YAb5uB+0x
OTqHD+GQNxwjJCA0zZEgrclMiz+/+mltOavN94lg0gzAs1GZ9QujNbw6oKIykdAF
gH9FgXJq+/eA3306EhhdSyGm9dqN3SI7SHjbDg+WpDqfcBV48kJzqnM6EsaZL1sx
IMfBEi/Rq0/f2RfI++1OvG9DPco8OKjQJPuDjC3gvKyCcO5ppv8KJ2wS55YrkckD
Q2xgKC34htQzqiMPbJDt4ReH3uTpsbDJNP2KJU8BKe1h7N/Q7EfhFgf4rzMARQ5w
Y7Nu7z6G1XOvkSxdLouO7h4ZzHLV1dq71HZ4f8hmQ63DdrRhsKDFLCfTTFMZBW8q
v9Ypl7rZwUl97BwlWjwv4mByv+S8TmPVszn1J3YpxGN50SJjMcdaaeC6UMZkvdK4
jukQ571yINgttl2S+4skkweEPVYDvP/dqKi0l2dBkAAacRxFvhaMkVvJV1QGEbWN
zAhj7rybgPQnlUErytUb00zSth7hjX/l/CwM4kEUgKZ0uMMgqqlKTCLWBZ1pWmQ9
K2UOkqwv6WoZvpt9tKfwr/OZ82Q0X71Y2A+xw1gMQKl71cwBx9ed/kXx1H1M8W3V
oErcSnR9ilUTf8heAPThtWN0R6N1eiO25FHA4eVUvPvfwHYFBCDY2EAWXEg3h4N3
dUHvoEXZexbR9x1FmcQhkBAnvV1D7s8Ob8dhz/KpxrTnw1WFuXAuTCAIPjOqsknm
JIAMQlrYAHY1noHzW2+kTHhV+vR1s2rbdaHTiSX+ELMmhyqd07RANos9MenzknMe
doJCoRwmkrcLhEh6aUrkqKSMURfnsMXRdOD+Q6r/7fHs4003Art8/N7CGvgB7CM5
oJGBDaAyqw6d1B0oEtU0p0oeiIuTpJJBhwDNLwMctVtebWnW9GcHlLHGLcuyAxP+
t9+z6s8F9/Vk0bbmrluw1yN99PA6zCHQS4L2Fmq0K0O2K8wQEatOeiUjJb8b7+tX
i6CbU4yRyakLHEufcPg/7/uDfw3UJygFrT5RfBKZ5c+e2unZLce58TPoxBD7DX0W
oQx2bcXEwUtqMbGCWzWjyFHQSvRYCPOPUYg9rczT4H426XgWBJbtAcGUyegTS0Kk
7d5C2DsDM2EgLjIDcWkpvqGKbynKkX3ISUbnB0gCW4gZGNvNKEXsmA6RhM6BaYhM
QomrchfI05v/vp9biiE6H+D40jETKg0aPv2oJf+eZf0RxlCaaSEJx6iKPn9hCrqu
vqlBsvRL4cBMsTWStaQNXwCaR1X3KRlXNuIjOgFawGo037suw+7kD3UUPcNyy/yh
UdQHmwtai3wad5+5qIoU9k+X8SL055r5AzH9wsGgsMy4rV9voz8W1PaBGBzcSXzs
3dZFUHf7loVsqa+lf/l3mynXyzwzzLBME7pk0wHValILAxgbeGM0AWMWUpuFuFdt
LrifAA6WHCLHRUXcgvmJWRTfwLcUcIPV+0ES/5U6kf5PzRH6hw8LjMoAYqKLgyY6
yuNACZMj8kx7PBNs4Ny6fUdwUFklej7dIaQu4pLkMeNaHhgWeE1OZIYKVF6FRfIy
/ywXr+xXq3D0nLZhtvBWUN/GpYzhUyiOsyeW7uynL5M3x0EdIF5e7ZjWWfcbSNV3
z2dOenVuIcXaBJe3Kh1MajjdH6jdPgqLJKqCYDGG6eG0uy+aRYobizlEJwagm5Fm
BG3G0J27yf+BJNyqADD9wNPkOlC1QJN/ONisNSE0i3KNV3FEOWyzvsxGaeqz2m+V
XdiEC6AGj4CHbntWonDEXI4cpXnYEmEkD7x/mtJqYyIA922mBv67oIbvNTM0g+hs
0/r84oWAxdDysugI/FMnQ3nTAUqpjW9InqfvcuqkC/ufeWOPC1GS17VeCXLVRUpy
9IMrswx5pRD2JfDRroyJxMeX1wtaq+xR6/Osu+SPIirZeteeG+VEJItRhOMX0OJp
rABd3see/D1uiUZkkwFPaU6EBu5hkxpPzHmCFkeQ0l/UNZD0/wRmzUIoWoXb3l2u
COznErmpuCgW1i7cusdX1EcUTEYrjjCXj4m/6HIk/zGQYGjDffBmqkLsXL5BvUGl
Hv2NyTDvg9sIYzo2vMtrT7Vj3udilJdMG5Qv3wvkD/mXUGQxaD03jE7tq41I69WE
3t/gC7dP1vNJqXuGf/VS5ft8F/qNYRIeq+Ry11jk/XuGVIkKM6VJ/Wt+CyD06IC5
eLVPKf39EbKfIgfvzS/To0rqMNg7rFgpST5gm3m5spvuUZOd4bGHaTwD43zd12Yr
Ybf22mRHx0bON6n+O1PDsJyBVPwDNyKENuRey2WvszwfjwtTNJWL6ZJc3SvzfFIO
PLKA51P/cF7oO1Z6Os6H/eEbfjZ0p5lrNK0qDa5viLd8f9MHu9H1nYuPLkZoIRuE
tQKBbEeCu560L13J7sGGetYFIQgxEUBu8BXb3kFc2VTZtDfUG2WuKU7xTgL6NpJf
+s9JNrPYe0uYI9GgzkgJVx+Ux53MJqVSGvuk1fTSIFY5FhEpJlMXJ+BkVl80DXKl
IlJ4E3RCyKEzgEUoVFyQcvCPPMWkPBYT2jHndRTW2KoXl+jLoc2GZbXqJpAUotMM
05vTXd2+hJgvSaC9obEZdpJ/4IC/BAtCEiSB1Sdndhj6ABG00kIBLJTdSrpDLsh8
hGD4I5brCV9JRds9GF3PNm6buFBLSiMk5seKfpyqMoF7FGu6S+9qnxVtajX0qD1a
SHiq1Sb1IvhJYJU+36KqZyozah48Z5OF5n2swHVCSqm3ib5oZadAO+6Es9uJImUu
M33+xmCn/RaGerSoCM8qLBe08kn4KBAjWmDAs0VbWthYjpa4Qdf859T/UNJUpDjg
UKe6RA/yVIFINt3MUw8BssaGu4KhC7q2UDNPaW/URBMyEigrK/+hB0I8wq3p8vM8
8PUyOK2iw9Bmg7P2UnqjIWh5yTZ6GsK3HVRptrjR64uUEiDAuJl7LD3UVLhl7QyT
1AchnbVv4gZ2nHcoCfQCvC8IRr8PF7lJDaeQ263lqgPv3sOfpnO6VK9i0esTNvzn
P4ebBMXWXkg6fS5Ao031Yan3rqcssOEY3H/Flp8BpyR7D3wFS5Pk+jhVx9SJrsW7
3GsEOrt0HfCCJFUwnRQPVPi3Pp8Ul2sAJ60rDd1CcEoMwK9vZzNadkjr+IKoW0yW
V3WngQ5RJgXlx2ekwkdNzyuq5hrHEeueL9zlA70H6b+NQS1p6Ms6JgpRgth2STm3
8S6M8Zaf9cSASWlBPolSvlhB6IEEPSooUeM2lAONhoiuniehzujj/TMwMeEst4ZS
7EYaWHkxk93SV3fF++fNkBsfx0pel1EL6fN5VKWazV45aJrpCnOigs5w0hZd+2S7
Tltcn4Wr3ImOyV+Yhrfnp3Ej+EI9BS6J4B+d0OAcA9M5CNpcqSoOiv9f6O7IzRww
rp/NbYPqbDAHNuF0mk8d75iwBjWwR3irQfzo83VytrPte3x8hN8bGJ4MIKyvT4am
9siCcn094RTsmOqCIkynPLeUTD5MXW2rKyCDbVYwLl79F/4DrJT0dp5M1JNbqvxs
wxjo3+jtybvo4bjeRKsT4SgVdBqtKG+t2Pv3/mSpTjzpPKv9OYKzgJAwawqaC3VP
TOcfpkrFrWqoXeRveNFMtWIlVabScA17EB3VBUl8M2OLEwwu11NJ4hgAJ4gSd8gs
5vId5JOD8eUllkmweteWeB+ML33GnAEKrUx5zD2uOiaEqID0cRlGLxYHihNJtTww
63RMUiEeVTRCfELwWt5ru89iz3wvsHSCQ1XwCjIYCSH2VHig+lpUzC71OpVbf7bn
y4DRXi1JJYJVDaYynXNg3tdgRsPSwHZcM7EmpTu38FQAIr9KZZoSVz8LfwE4sUVM
wAW3P8BgaYVOcMZ4vulENRqA5vfMh83uMItguHElVnRWWUI4mNgG+u2i3qndSlN2
7eGjzj5fp9sertqey3K0+DYM2stAlMgIc0rDKmMwb3x/dlkOp581hFQ+fxXLE1KA
1RxAHjKH8uOycmKyW20UJ3DMvdVwRnL4XH/+7fwVDUQDh1h7NL98Zf9RDGyIb5h+
xFCnd/Z3aPjX6kylmbjFZY4fFCwp5gQGsQj1gbDZ4HUioWUP4zJ1Gtw9wy6Hmv5W
xLmSQcqt7MMU1uSxMXi7i2W1wVBvvCWBXpAnRlCWJbYcLkb93izEPPvBzpYXzL5b
kH19+jfumPwdwLkjXLwDbnPkiacQ6j+yodY/lnqjf9uqbps/mdMMJQFKVY45lLxQ
vvCzVpBeHjkYQQN2zY88uT0pP+472R8NQg2KT03WpT2BRgM+m/V5blGNqN2mmyaR
c0FTwqUqJAcpEkJt3Rjc5Nd0NVxOpn93AT4vxJvaL3/pSD086NGhm9uCA4S4Dx9l
lpw8kZWiTSzS+WvtrpuLYqL8chHWBjPAOBTklWiEa9P3fIoLTrTEh73VE17/3fjv
gmM+qqGzOKE8D/QoGOr2EGzy82CXyeD0qb3w7j7nC8/Xq1PlXsxFLamKF3VVaw8h
YF0r85esBB5k0qEFyR9Y1HK2OtCNfGby9dK1D5hAvg+KrB0njpKD/JlY6pUgqaq2
W+v2y+9J5v0GKIvqhoVLTzGHQnYLxuSSdAiK505dsYDT4HvhjttDwKJj+ICQQs4+
achBMmQWakmjsUupZ+nDl2XbtvgzHp7Qgz2sliI79pDG8pp/co6KiBHGah5X67kY
nanIxBpoEsv8C8M++dvqHRJ6hf3z0SriNvstMoogTPLb3ERURAfl4wnSxubS3gXV
g8GYnApRoM47lm8s4o6CQOOxjM0e5RAHAEG6L9/dEC5YYloOCIyntDWaHn7CJUR3
28+VlCZYbo+R4ePlhTaJVxQcPObxfPGd4z8kMKYNPY9czmQM2hhryA8iBYzcNd/Y
R6K3VoXRbOsrxpMovEh99/McgNMtQPxPcvVa+J/0sUcDNYim7/7ACqmXt6gxOzxx
rRzxJUW98rhmlbmkQxb6s8iPdGBYkSILGnIZB+eWROc3MdUitXv+nzkPf5RTCMV5
4eJxQTxCdAwZLnH/FyxEbgU4FofWjXu0P1+P/OHALdE0S3RSakJYuBeyZy25xutY
Q+NuTI7Ye5rj/OPssdU3fpIlfGO1g79JhoBis1uGUAfu5wu/TD/YliLefuSm83U5
HgNoG+cJUbDRURw4Sa2WVPIb9UnLlcOp2w4ujnvN6bvuZJ1Vy9A79Vcg6DunxZD8
zmhrGenrNgKDtCtbeOSQGsF2XSMoHVj0s46DXkQ6/gDQxPUMOclddVbgtbpMAAgZ
TPcmYDozGvd5fRYZ+W6EfJCPFPia6IqW84xaZCswy9oEv8VDurKdYjXopTTV914c
BHusfGrdh8ZkQKb7yiHz9+IpxNMunQCuycIg94Ta7NNmOpymQfF8UIGU0SiK/pbd
o1tfL77vfwrlThpvZtmTmrbRU72X0ml5L5Ra4ywkJSfaeOuN6Zhn3lF06QfdgBmG
4EBU2Qq0F/88AmjYusLMUoSiiFvDGZvVZzWmRrIoIhk4za469/lKE34XXIagRiuP
ND3LwCfpGclnsZb6ehYwVyJh7wdsyZU0egUl65l6eMnFNa8i6AjJslzKnpjSRhBw
e0h/2ioHEgQVaBvxQXgCM1H4Ft2q/AQrKgyzdcuWxcpo+UvcaI94Jte2mwTPgw2Z
NVOWl9xIxSF63D90UQZOIoetzU3Y0hk85StQ+swEEtgETSzJn0bw5HzCjhLByVFT
JyH36DWIZYfTGDe2HYzZSKPrtvbPcPCY67Cr2hQTCTQjt2BXbAkCwzG2RDaD9OBF
jUfcC3kiTN8CNFHpgDtXnaFaiaTBw6vBairb+ROF1Ch4TMNpZ43Zajvk17u9Og/g
AUzwui+FotknRNPcM4EyZW6+zAINKkI0vMCjimy2nMDY8YA3hUgEGXoL18Jp9xxK
JgIq5UioWkHdBs3Ww8IYrFlW8kyunYnVDmqqckmql7NJCtvu6u/jA6QvomjcXvYe
kd48akdRghTlG+mZCiKwd1AYZagyovPgJOptBjNkvL4C78fi0H6jfo+eEi8KlPTY
N5RPFBbCYb+GtgSb6Ocm33FrTYPTYMbwE7BREOaI0KJ7ZGUuOvqDEagEXPzA5ExO
PBsBQRNsfQ0ofWCAujyUyBJsnUy8/yX+5mD1nLDy9Hc0WflZRhzn6rrpC9YPlP83
ziDlNAC1wNZA7Uzv/HUfqyLpa79g+3J+Bnlo0n8NUmZ21VQCka0meIatRlVdQFaj
vfdQxglIALenE1496E6OL5rocjYRgLNOsKbytZ19O2GGBqnWMB0xlgkj7/jMo0qC
vCW7Nc1l2m51GIomkzo8dWV14MdG+oYnld0Yzc0Unv0H32g+0yTgeez0bFqG08WU
RDerVF+MCo54dQA24RF0cnMwXpgeByDX+CH2f+4LYWRcwT814STdpQ7groZP6yNa
gv0BbPOoXae+Zq1uSLhW8shC7/gxVlbUusZxfW49Er+p9hFP1r9wARWt/RLKf33H
1bQXSC1Qxl9oOY9Dv8toQ/zOBcyJhIWGvmKmQ3FdxPH9HPFGTqXBPlusLZrk5fyM
Ilyyvgh5Y7tzUh7Y0NgfLMMhNYkIXL5rR3qD4OKD0syCvmq9pWdzMpRiZkZhDu2n
ldCl+vfuZK8VTIFEQeoIKf6QcJRqWEgfagh6TfBjOIvRQV8MG1WXv032eR6dF3i1
p46vFq4brw4OEy4B0Q+46C6XLQabVNZj/PR190prejlt9ZW+nzEVGlCmXvYMATGB
HtELwEGBdhe0KJzEJOvXdi9Xb7AleKxtJUvcF+fGZl3vvEGtYEbeQ1y4ZSRZHvWq
aKkbj1rXxZKRL1k0IX3qQ1epZKqJjiYeXaRiGogUcXSP3DsaHkjHvEIgy2dBp9x+
zBXE3ygomZ4NKTWUX1QZdqRWjaQ9p3NhxIpO2RAXMYLXfrBQb5h0L+4i6Vj8gfg9
okL4HWlMMDGlYWyvJGfUbP/wl71R4Vr1Zdd8hZWpYjQf0+xm51Pud6Dr/97QmY+n
CdXXjY5u6MmdGEEdNz/u8Zy77nurwUAMQ3zeDY5nzOggFiHimjcgtNVdrq7q4Nm9
EMW0rqqijJ4ihi8ieBL0Gk11Klo++nS/ZpUylMbnf9Uh29ohfWFdmes7QSJsWiB2
xvq09qtoFUPxa7av1CUnExSZHKg74MrcNarQUCCCRyrR+UDaQv9rn/nJuX9GZy0H
a45QOwDTBYlgZvI9UOIS9abMmnaZ13uVhNCCjZ/Vi3DKIjqlTSCm6ZLEIPEEp1Ao
YfDH09nlIBzBarq3sp95gopPul5Ft2/o7omXHyQfEdY/cb2ChQ+Cb1WyJI+lgxZe
7UBnip9+GZ++7YEZDtBbXClH1GJFZRUm1COERmOXRj5m4WqVRa1OVd60l3p/QJVa
RKtizsVlS4Z4YL5MlpHeUSfl0fYPlzEXqlcGU3Zjnxt446OXiZHxSVQQFewbfT0k
I3veK+qqYpLnuaxNRYyNn4R/VJo86hJf0WKmFS1RKyK7fO4LIqWRf7/BEVdOb0C+
spWnh5PfxyxrEpyHV4UWgrAf15fYT1oNe+goS6HyHRFDxn/2OgYT5mTg8YXgM5X0
SMZtXZ4+MNUf+1yZkagGXHe8beerSxkyLv1e5p4vMiUHB5eJ+CkExUzfNkbMqOsQ
SpJY8YmQHNXT7T4ky07tPAdj0Sot8lE4xB8hndHDr4+1GQeYXyMsJ4WICvcgs+oV
K5hIljNcW8/CJYFl8+UxZvhvySnDnLtJ1elty5EOrSoUxgCA4i1BpT3iS2T1Cm6L
6CmSvUSwGtupHxDMXALtrMlfbfE9CUKu6qFKd0w1xyzi/w/O5DUKY4ZWWsgk0+T2
b2QdJxOwTHBgI53FVXhbe0blIkbQA7kJS7wi31kNl1fAQ5b8EuQSG/e0voJBGG1B
wGnVdi4NMdDOxJlbOiG0YHUPHc3GNRDa0I50WkIHEnCAeKwy253/QjVm+K9xprut
MkjyiFHwevLKzAX4/WbbsS3cvh2rNu7jeKaln9o+PpblKbYmwJuc5XqvHqevQ7BH
pmpYrNzxaKS0sMf9TVUwDD/UWfgF5axsSGC6dem+KvIJ3EaWl2ccFSPe4daFg8RH
R5KSMSznrQsrRpA3aO5ZfFbcdDRr6Nlg5ucXY3KBWCG8V+OGHcnVQvqvhlSRQwq9
RR/7ANXHU00ch6Uy99sqAmVbb4rnU30z2pI1uAl54Nc8TLeidyop7oNmPk9aNFCY
EZ4zmdVqUEDF1vhZp6JUcgh0m7yH9QXZG1zDMVoH7aPsnDE0PXl0ECV/VBtfSgWs
TSBzgKybt3JgK9L63kwOIptCCWeeOPy18OvyYlWqNYEUZF0tAEAK2KslpI4ZbRlG
vwnZtBe6+V4ZQX2lhoC0opv+U9YyLn/JDOdfUp3UcBZG/q2qB3RCviP+CZGs2tW8
gf6/caJvQpk9CjdU4pp1JIFdtEsPyNSYnE1NmhXvLWwEMgPxQq0GdOHSSAMpudvU
NMednTMVoJEdeJI+MuZIuts2R3j/+j3QLVSaN8gLe3LAedSkx8CQvtlDY5mYWtuP
Oo9gDXccP2Wvxx3Lg+cBfmEvCUuYFEMW+FWK4ce6W44dKawlXkp6gcHR9D3qNGeu
o8icHNFuRAjF6svuGQ4ae+cCUzl0Nz0GeiVczebzPit/VUd8TZ+o4eH5VFcLQXKX
gqytr2JcmzaRMpWPGqE6wq/lwXv7lEuYa6X4mhrf4TZeVtGV2qmzkZpnAraJG+OW
dPM0d8L1eSlOXHiNNRsl7qYnTdR9wcKm0GCOBgH+7AawLNZQ9un9EE8nRBNdMxX3
6aNvVECRoM0J3jfGQW/tLEGhfgY8WGZHyARnEJj/y7XJ79Q/WLESL/9gEBIixllG
v1mKIhHi9hu9eAP3wplFYpZaknZzcLDpKVLDhQyiA1FG0iIj+iH8AOaAMMB1NlUA
t37qHwKJLrLJTGuYk05P+U9cjG2/3OROdigYRVDiUITvEnIKbYbzZY+iHZu78guz
j5f2FBJQyERBtELpMDEwmOPdb1uq6Xa3B7ugb5wpNQPWRy5SCrI0dX13PJwQxsz7
uGa2fpwx4AcQxy6REKP05A4XaejYE30yoXzXMrPqFbpnPhbsk9n7O8rV7R/NIggI
0k1ypp/7vj5JQoeuy/+EkO5qKXenmnfzO+icYxrxMcFfnuj0Df0g9AcufHrbuYZC
L0aefOWSEHFFC/R9Cv3InyAh06q6XPsCrXP/MF9Z5hYq0B7KBiK+fQKJ2tzbaiNw
vqh619I0GtSKn/QnCseDEuyzU+2Jxotv8dwa9+c4qpUC/ccU720P0dNe03yaCnvk
QZktAq6nIdSay7SKvG4k5SFEfugxNppkuyBb++vcHlvs7rTX34RHFQGd69zqzMJg
1dDk5XnpNsgx48b2pMwA22d/HDeZ5wFiqxiYsbvy6uLpA87WX7afepFUzRtse1sc
3Ydv/ti+e3+RgxcWcIiAeAfP8qCS5/w+0OkM5qpm/LQtENYswDV9kpvcDxNy5sQu
8qxZEigFW9UGFImiMDmri8XjCbfjXoZRDho1kgAKUc1gAW9JyR0B3I9QjDvyYANo
KAmOpJRkLJWCWLI4Bz1plGNNkLOycSD08tx2iV7PO672iQEiN/zo6ZC1vfLMCl5Z
ILJwrCjg3xncft3y/4+oFomhxX1CZ+CipsxaZw/wO5SQ9x04iSp1hLa1T7UP7UDp
NiJHnjGyPzwTogYm4AxdvOOe1mRR5dVE3s0F2chuuYpQ7qa8Q2NrRT6sOx3GgfSE
U9FzxXjLSFn8SAod5KS9H2XKivXo6BMJA/dzJN8+KEXB0wZ3WSmh7qhOETFGuXHe
z9k4gbLfSESvsbxxvl2Tko21L+Kl/7x2X3Tb+d7twKSL0Huf97h4IUd1ojMKK3In
3MhW1VJv+iaDYS8xUfmUlFq+BBsy7Taa2g/sgfbf4kzSyFAM2JsF4ppw/HLGCXJh
OijuEPzBhbjS/B63CICBIA/l5jI3FKPF4tT+cS18Yea0LM8TL9S+2B+YbDsPSk4E
IbNZ228UerIgT0dpLUZwbJIRRgbmd95RRNk9Lnsz8Lj/Y1PGgEw3thXyJJSPe0B/
P2uC9q8dxw3oTyUKBtaNNZM+N/RyaG0ENwBVghgtcwL+vgGvCyFfga24Dt1C/ns4
Sc1WXRgqYvUEwMTA4WSS0H5rKUKLVYx55lXbHEsCxrOPsMbIyGTS6AedtvwAxk+w
I5dqn+afwFAEgXVrcXHQsBWMaI+NQ0UJV0e/MZgTt6ucuxDdAa8sFxKDR/CPI+Sj
ws+3yaDmL15np+iVNywuX7gmi0+zQcvxbvn7UkyW6kqxKkAfVG5HOPggNRVumI+5
PurtcMAD+0GKeqxyDuTiJn/ffVutNA8Lki51sWVNqDRtiCkfx0/a8b1PYcUWDhnq
4mwOj3+5lhuA6wp4yT8UT4XbFk79x/8cCXsdZ7r5DS/HBA2XyrLdc3aRyemlt8ln
RuqN1onEgiEfPslGyCbelN96B61NJ0ZqV3ehsVY9ESCFHasDF4HhEGH5GJntmb4I
tNYZWpRkM7QzfST15604J1JiSWWkNa0pgdL2poIAdm26jDzW4UMoylwzDZEV+7jf
E/LyP/0br4d19qt6eGGkSE8Ag90+m0JlJb5WoVEN+1x32MKV+4yno5XxdL6E/hk0
fRE2zVbjm7mbbMDFqRYeoC7eQldd8Qd/dtGhuAbWoPMxG2G2JBK9qxOOi38VUAXx
/eYbiy61YZ91H9bAZev7QTZP8ZmvoRp7XrBZEsiMhxn8p5O+9Y75FRcB1VCXcdE0
/kmLbjYKIfLtOcSFauQFZ9vNKu8Q8uLsGXNahpBoPRWYAlgKpFkQRfZRSKzE2hID
1rjE1K9pewVuuxwA1ja0qiNlz/t1x42YvtPmOGu1B9SGmCWXvwKA9CrU7Wwx7P8K
zYM4RVZBw5HxktuX4bO3epsjR/gf73jmCKRnWHHg7YICSaYfY0gXG76mUVLXGXpY
79Cu+bLHJ6uS+eNL12jWu8p4erpA1cOzDnyE9Gc9Xzr7GuJGJcdDHpNv8OqN4Gzi
uDlJ7ioul3Dkm1qgvrwc6/BGTGxVorN3tkjptORwbhbLkXpIRv5FsmlqTSl5b4X7
UlBwF52O/3X+x+WfQfKMu4GT0+yZuEX2GuEAD6AT2Db6i/evD5HXNBFauIXNuzOp
UmXJ7+BNDZum2UM4OBx/+5MR5wLRu+IYdbW+WDWU+K0p1be7fpPudlrBvv/5raKs
/kvoQ29zUdCKnyQJFLSi7AkwmPKF9HGHN25BNUE4DODDu1QFCfTGHPCDUHm5NmMe
TR1HZcIplsFzejdIat+yl8ufg16DDGsoXDH0SSYyMIwbCLYk3AhYjKd13KCmrl6W
JeaxAxuidSpFSwEI0sjrtxOZx5Ox6V8VqJAWdSi4qIrgqNgiU0hWaBNFlnQVnLXm
GJgXBBGCn5f4tKv/DobtWsVMxP49HawPy109S0eItT38vZUf8DXA2Q8rEb1+v9eY
eBo3XN6T6TYOCC/EcSkqqF/jhGI8H2UBHRadKacZ7+cRikQdlV7Syz/kyG2Grq1x
Xxn23HuVj3t5P/dgJ4IJg17vXlB/KAPSK343lBBSVF+WA5TdGiLWYgfRYJs9J89/
r+bmK3AW346Y04KdnM6ABQIK4tQ0SsZjnSmvgSBsk3qQS4q5uRD10tnq6NImCWMx
1LMrwteHSwI432O8UQM4AfBa+gC2a1BJTHEz5AHws7nv5AyyJzhivnXPuxS8g33F
qt9KGojWH1YVM/nnGNAVAWJ5klKICJ89TqHzXPyWY/M7Q46Q7SruLlcqS9G3Mlfo
5OjACMPowhdob3UeHUfaVrgXmZS+KLJLFuCztPOb7TD/SnPTZltIImQmbHt3TtVk
o54XLGwMreYL7oKbJ912MVFLpzSUTZfO44+dHpvuzRrdCR/uh2m303L2qi6q+o1I
6fNRntw/64YS9cvm7zgRivyYHPAZrUJIWC9CwVT2sXREm0n0vKxDJdUEz/9bqOwi
7dbZ2ZcHs5SwaLQDmhxDzKznKOWxOsNzPn/2vrKKSmf7TJfFo8IFIc1gvA2E7EPm
8vSGxqUO57pMpIUIlEBQjEnGKwS+EnEFz07hyY4/KTeeFyueeMiPMNRrPGfKU3PK
YeFe+87egfTrU1lH2d6e2iLqIwnv3dAsGL1uXlDFabqtGXSy6C3xSQM1bQ3nPGpD
+sUq6bhK4hieTmNFmH79gH0aKaaM7la0TjAVQ2567j2AUP7mEU6ZUuTQz8biw27c
3P7rUStkZHIjy3huMI6u0KnR9CjAENd882XtO4QAAZHQMXjGxiQNpLx6cvhII+Yt
rQScsh8Dmt2TjtHSECwUmYe8zqXFJEbfKZuqoyhhyNeSmntPWA8FnRdZp70fdh9N
29EAdhZgvXLELBJ9YkQXuLq1qrWhAer8Bi/vvWPEi8giC+qk1cBclT9bR8wFPD8T
lx8BbCyLbDzZNADAUQ/ohg3uKMHhUNuNOEnOO/06DHXPDmhcokBqvrAo+WBqxeeR
Ll5wesZMjaQngHV15s4y+7pZaqQwlTuGzA5dAWr4qzEWYCdQQhRW8iyNVPE6S/nF
1+Y/EwB5snWZl1hDqgeE3TsqaLefSg39o1SLXwNIkhT0Kh6R0zC13eMCacLaGaY1
M9pXKJg+ZjtNjR15hL3CYUb0Xmc6WxtAnjFKCsPTSgJWkKZT5LoMMrewJfd8Omh8
MtvPVIja6WjSUc6ChiMiiTGuGO8qGfFPsDPRVJ/8V2S7pAbjL03oppAoShihrn4N
WMcMt0UfTJFH5tGgUtTdruRQnHmkIMYCXsFkXem9V+bcl00TJq4loN/SFFanMIl3
7O8jz3DuXgYoWHgv7RTBocnyi/nHLWZFnm3Dad1XRWV564JtX05v2AniCpaFdt8u
C4EknNd8JCGKz2mATBTE1e/Fxm7oOSGeDuSr6Zz7WmhEf6VlK6uMBeJwUMfWZ4Xt
+QH9MFAKV/J/f2xXM3SFAKtMa9brKGz/frv+AiLcqowJiAM48V5hr/YJwluLex/c
TrNsOkWuhR7peXSBibXB9phpR070QkvnuhzjOkVxcU6k8SNqlPCqA7gNjjkaUpJO
sZI1Z5B4an31SFHlRvDioHg6Z9yzURbqdMHvyNEErSymnnSr4HxwQeexxfQXYHVP
/R1xSuba8ES+fbTR+BFdO6asJUVRC6z5GOhGO1R54l8spC7lHWrE5Si5WuP1kV4d
crIjtkP4AQ9nsdx1Z98lVus9PfWrpXcIFGtcR/ZCR/yjULdiLzbP/J3tN+5QGFew
ju9Z8ZHVzguZETOQXT++phtf2IkhwCQyiFWw6H206qEWnNsQ2OCHo10lsTQNJ7lY
b9hMYF/7ld/7rsXrvVMkdphClHLgBpNqvnkbSwFI3B279PUB0yA1CDuWKcooPvxp
w6CC/AernVgXiAp8jl47kpBBdXELZRNPZlkfVnQyLUmHlNIujFOhFp1rnhCYveyJ
RfTZxcXuPSA5r3ntB1zCbxGhAU79vF/H8GQ7ZbQ6keq0Lrmq5Mi9qePxASRzH8kw
fBLYxBj9mVxLSMhdQLH3DLYNirOwo82wAAxptEe8RycljWaI2OyH3VT6ZZvl1gkv
BZFRvx1iwxACfFvXVzSgTNTvspoBhRhOKrWNPclTJyvId8jUIn9pVMYdxJQRUqUZ
iYs2oR6u5kUXRtU+dIk+VXd925nkKycz+ySX4LNjAb5tBvFBB8jAuQgcaQy+VSdz
NHUcuigy8Jog2HqJKozcosCOAwHH1mRgXNcHZfyZ1n7AQqs5TfcWCBYOfWx3/t6Y
Yt+RhKYNmbqNahYgIUgl5UQ1BVQK/xmYcY73nW5Jrz8nva3q1e2GeoIS8nn/T/IG
uFFA9e3fdPm6y602GifTzzuOZ+1VlM2B1rbS8ClDr3mlts/lOiGpw700HY54+0Dl
zYQMRTY2UsVGjHYYfBijiL05BnuZGnfXG70rFqMTPGMJdhdv3sZ8XqrE32CYUSAq
wO2ZTK0/EliRjJv5dEeiFUd0a56e625xVGiifhIOY+L3smIqlQ09qdRoVjtr3YTk
olLtUGjSqSpD43OsKT0EUc/jK9xlDsLYjZXvmJUuXHV+r73BYdBWI0tP+LjVFiCg
yKIH/u1dRLGWakwTPi7uUeTFbUhAYcp+YFlSai6xushQEmRKYIv/Py5LepDGL3Rv
sRlqO2NYrWT6o3FMSG/Kh6FRRmIIMPdNcwp7h7hR9Y9N5Uz4NbM/QBr5YnT5a95n
MbsP3nOCQCKh5OAKsoiK7ScNl6lYZ8Z9mKcf5yq7SDqz6prSqoQibHMOJbNFr+wL
EzeZCV001Wz4QNEFNGUsVtXDd17zfzA1fkvGnQEKHHzdv5ULMUytfv11fPPcssFQ
CZ3R+D7ltzC4U+qTbNFzY2TURlvmwaX5vt88H9m9kf3iTAUeljdwpIlLA+9PmnUR
zUaA428rf8rquSqS/DvDJiZNxHKyBtULsFQMo9+jxCn941DcXYSN3UbiwqFqbHes
JBtFNWXO9mm59Dl5ILXaDBLqsT+tJ8bOSwPezGv+0kCFklmnpSLFvZ7/dy4ALiXm
Qrh6Qrg5Nap9mNbzsZKt2yX+LTx0z1Bhnpe74df/nPB3hebthP6TEg2kQxWZUaV4
w0i1z2laP0tbwnWy5wcAQDQPrGIK33cCWPCt+I4U3bUMk13Ctyp0TEfUzhksbvIL
yKwWkmy/HopflWBOyE18aTpBEAZGArMviCXMJWriavhQhwcnB0A6+d9x4gbhRHvb
SeJLQsmRd3sgAIqw+hRlBkgCI1dBUL3EqdKt5fl8iGhul1SAm2Ilr78QFvvtv/sg
mMnZJLjPpUH24Q7nN5V4Nxab3yx4YmHTkTlX2zwHkrSxLVk3kmBYQu4DA8ZXpHoP
1FuiizJcyFuAVte0YCyNTf5z4FqriecM/Nel+Ha2TLeKAYjVhlL+mCejrGfrGbnC
gNTBAvRNPD73LIu0YMCIBitZqfnjfmkgW/L67S6VQJ1GU6OyDWA7gBK0etey8rO1
gWygu5ZxDUKqwgXemBk4YoLAOh6R5AD7RUJ5go6sWwYmCM90C1X1bhqTp2lG3gPD
eAvm37cwBZIfDBI3r52W+E+/HrHXzSifLZwGS30iX4q8Tckjgd7OivAUs3ZF8VMo
FNXcTlTthxe/xwNBaLqGodoqG74layt1DvsrS+jiZyn1mV47hSA5TpYvUqszEDl5
ojaAppbnJDqBbe8q1jbhxgsl9/nI6uTG5Uhg8QBeXfqkO8+F3DI18D42ORdIj5r9
CNVf0ffSBCze5CENHHgwgurkeoLLXNTtqRQthqmtE2bgmznoQlr2eHsPLGsxFuBk
QfrtdnVhPXaoIq3JdOdL/f7oisi1+UEbucm9OR90u6FTt2jPG0vmN/wfb+Oj2z/j
Q43RF1I+USl8JY2eV+ozOjUufiZFB9PyPJh2zCT7Y3sJ/TL5Zef/zDsqg5/ClJ3q
fsqOlnHW989PsAoKhBZwtPyDHegeHP68Pg45CnpKXmvjuGRhiXhDyaI1NOBRq4oi
SksdG0345ax0IIArm+8ekJWJ3mIplbbwIEVvj0MmczoPe3ajD2sgewZT0QOj8+c5
H/UzWCWA+AAOu9yW9u51VQf7cP8XVyNFVjZRKpDQi6YmAdvo09unFBJ+bmfiOFdq
rfxP+d6vsDfxedzfuKNQFjnVVnjfjIDyexq4iutz2kuB+NxF0gCfS0yXGp8gRgIB
hstOQcbtK5GLxpQhvMM1M1y72SBa2tTaz8dMP3ZSjcwCsNbSffwQsOEECrhEpgDv
nKODbTwfvcz4r85XkHxUx8mQW6WRqDupNY/9pj11bp9oNaUPxkljkZE9ArxyUaoS
ugwp23ESEyvfWjGmhj07oh0IGXjGbpgsK658kzWMd/P6RKXsnXj1Z6ORlYEKUJC9
B8zI8SaToBSsgVK9bAHRNOWFbsDlqh97joVtn+IWJ7TlImY7KpSgUvmt8w7pS0/R
BimGPGn5e9z63RvAu+7Sdfesv0o0wA1OXtBa1xBcRHhm3tvL90VKW+HJXzKumgXJ
KymEK7c1MUyy0yw3fe7dCUzWNoF3EauStbFCCs6Zq5dYq13DKB9lPfIBKABxdBy/
bph3wkLssS2gfpE8rRDHSuF60RmHgxBmwfzIiDmgwvLn/Lxkwif9Jexy4FS5+Ts2
iG6kDqNt9aXK0dzKbhJTHSQoCQ0k0HDpG6dqOnx9E8t/R4R+ao2HlevmxrcdSx9o
/TjZ99d+ERAY2L5AmB6tfTBfG5NRFniuuowrQq0BB5XlsgrKf6gl8H/QqeX4C3Pn
4sfqD0EGLopGERPmXIjTFrPufiPZxU2Au+YgMwKQXNdurFBeU8oOW0UPjx37kiGH
pa/GD1w8Mg8PullwkTMIc+XOV9P1ADv2a8dP+/eeJQmXKAmkAqqsr3xtA8t2pylK
ykJcYyW7sLnb6xEcO1A/+c6GhPfqYv0FyplzK9EFTM1v6axjl1+EQ9SYTyiTQSyS
gbJgYcPbxkbgVzdz+0z4DR3D6il5NDMppUa6O6eP+Eas/0zh3DNG+ge3qhK8ycp+
q/kCAFD7NQYxQAGf9EdqnWRhs5XrZRYXWdR5BAQY4aoJs4VChZ4a0idYffNNZnak
4MBHBJXSj8fdhibC4cmc/vLJyMjxpwRhut8W+w7tUL+Xq5w9sYJ+6TSOFHix5jvN
ettuhIOFwmRM4NEOatL1C8HDFy4MzFcfN8Pc2LzRKxFl/KkklaIS1t0HGp6HSrKd
EHSFyztSC52i+ELAfJhvKVCAOEfcJKVQGgOzSzozFlnBUw+72PtKnunOYOAC3Mh9
sUEsucXgwRt9q/OKS9ajoUuf4FYt/bMl58Jn1fJjE20XobK3k3yZoGyeyFZLy42X
kh/ZItATtUTjbd1YT7m1yvIAlW64R/WzoxzEu2GRsdeK1HR7eqxsesWLVDwFMjbR
kj6j1773gj1zjIE+BcA333ul9zN67LXGZBNl30YN/VTO9yaXmVtquRvgYuYQbesh
WOzUhfLXqmclvOV9wwixf+X02CqkFzvZ5a72yhAGRaMJG+LzeHwYcYwM80i2JbCo
nDyUxW1gU7SnfFN7zK+YNXeKgaz6+8uvMuN358BTBiSVkdUc2V8YNi6tIjbVRXkf
0aLRfk2H8M8Xdll4hlKoQYsrdA1lCDbasstJvTDF8W35ywSb8zEzeCUV0bqhqfVK
Yl/HHcTjXIJUaWdM4NKvNMHLgrGUYO70g3xg/R4mnCb1kVDTW86C5D9oOhyfAlQ8
qzd6RPYi5xAhLgrzLS6PfZ2eQqe+NY4vFmnH8rlc2gfFcnCsIoo64B1iXTcBzqdw
VjDMOoo8+s5qmRpi04c6fSpKYSy0+dRirf4xajT5vjJyUm0fvC82MkaNu3hvYc4y
7jPXIezFRV3YKwPgW1bRd8rJeMwenvFkUA00EkmgVjy4aSCuHD2sAjNTZepPXstM
l4w/qmspVqGARLNXXC25rWVYYVzoIHjINw9w6/k1dgkeEdZmim9sIYpTXO4DyP00
e9GfA5MT25a3QByDaYWwAN/32NwKyQ2ZrNeFZUvvL3dAQZd+4fq80GEi8NKChHs9
niLWhkV8AWd1tpKPcrf0HnYNlKgtItcx5tTxoHUS4ZHIQF+rr5yNHI3xtu7gTUeZ
kPcLHieJAE1AV2YcmhviSfus1qKs5NVcLP6mMC0Cc9/9rMCXieDaNh0nNKD8tLBC
6WJoFaJGg8Wbj1MJ07hg0gjYKi180zCv7Q43sgGwZkpTdjlEyMlZUafoyp9nA2s6
2jCpoYZmqzRiXaOovhbEiMmXSRi2VzGjKC3sEtVhgUF/NouCLSqy3m8GCFS9nxB0
XhEOu/oG0Oy3sFcJe1pOpw6PorO9qSn+u6RjnmJprPrZAHfGFNDRGft9tD8c39tm
sRigDCtsN+MB+UFfsGPdB+MAi1BKUgVyVlqUCeFlo96rtLIUgTvkMdlsPXOswMp7
d1GMmI05pOPCKUvcmg+6xg8m4huhy03g8rWGcjOLa4DJPpmoXDqZNX7DEXEZFnBo
k29O/+F7GRbwlLsscCC3d8pQ65Hx1XCF1962I0XTmkNX9JlJa087tRHgYXALenRa
s1b4E/Pm3YlKqTDDnmi/g2Z9o6DGId7Lzo3nBT1GfZVzS9bD96h60h9XQtgBL+W2
lcVez0n57X4Y46/e/A4i2d9GhAcw9mizyez4pFZXupP0oLYPAbQHWjKda3YfiG8s
5IwnxedNlodJy7GqFDLAXE9z5pKBLq5E6C50dMI2DDdQr6Lj79qlybTz/T///Tuy
z5BEeyo4wfqDRpVm8hAqP3X82Oo2I9LuFPZRimLtsKIK/h3h/HXzE+N9f68JTQpD
6WdNc8a0dzbuajqTATXbmZrZUDBmjvpUUAqmHEwjOXgQQ+O8ktbVgvKEyNDGDyWJ
g6rPB67ImFBW77bGb3SxjIz1/HwujuQOr6+Ek0JRAHCVXbNpfDf/1HeFw0s9e8RK
m1lV1y1AgIWgWgGedyia6WlLYgkG6rVQdgXlCxszxtWg4FJzVQLI86XhosBMjDUK
xCkIyHp0miEMH1Dgv4jDSVSvejBlqwll/M5wBAtmtmk1zgklCY+sEPaGExsgg45K
pBDOz99wVan6QhoFRYUicdD+ACeq+C1QyK1V3K8ivsB2pDU/H83ySUzgUqAPDA63
wSrLlSMcNcenXKQuHEJL1DIq2BDN/lNqZ3h97BFnj7ekvJVIqzy6xZZGK2d4Q8mK
kDzxrzoRDKCVNVTsslRYvtCLI6XfUT+oaJC059v4q29uW1VvIu0jOxkuUPVKBhym
Pss3iwq8nFEivymC1eQCLHfCt73yWmOmI+nLyhAlYZNCemmqSJQVU5T78oNkiEXD
NU86ewSRcTXWg6sz0S5kO71Lh5yRoupEDnh4flYhZtUvzKsir6m1raNJ0tHe6Wln
AGCuD+3lsCK/dGLRrD7f+b757nH53xFWpa6/nFNX+R1ooM8jqtb6zHKWMyxKYQ7U
CcFOqOcWnL8U8cnFBifFNxq/+qLYmthK7DV0qtF1WGjiHUwNEQk8sVtF+LWWzRHq
OkQjPNbylQetdHH/9oKaSwo6TXu+RSnQULfe4qzkoo6fl2L6gQLgOsS1UluYGQX1
U81UFkvlt7Wb7kctGirgseqabnVy8fAs2B+iIS4L2d0NXuhx/u7V27S3F1mL0yh/
XsGeC8rzx6u4PDVfDQtAoLAU8lXULc19Gl80nwbwUVEItlgIpZgv4fiiU0ZQ5h1b
4lAzbXmVSSaG7ALjHVSnD1wv1UDBDvA3UNr/xWoOAk8mR7Lbw6Ml4FvoZEH9Iu/j
rRXi0IvvpzTqTmn6t30Gjqs5Ozcvg8fqktmn82hNkfYuVk9ZMme07FwV/u7uf8ms
dEEbCRLVCOBf66ZyO57hopx0qG/4osvPgkWDF2WdMP2M8iL5jgCP/kk7keAEVZEq
o86qDyTPteMKp+1AE5SIfb+5w/XWLOWwEWQ0oXhi/GAaGI5fW7v1RA35EeHmPADe
zDtk3KnPvUP37FeeJpy583SpkvUtTtclJnFKZLEyRbHn/t/4UdGiXcCXYJCCGdX7
JJZbIq7Lj4tdd0y19i5PZURPzlDHn5GaGBNWyRUC9GKHPERRhfarAuLSUJM2jRFM
+L2dPW5muKzegrAfhj4yZWwfT9am6U61YD/fA3rNvEUXCRgeV+x8TCfmvpw8mEq8
XmjntlhkqyLDDPxoklcAFzGYjQMHhIYU+kgtY/IStonwywpKWwo5cnmgFIqFupmC
yMB94mlhpCm+RYa3cPTYYZFL9UZbDpeZX45JHCtus2bfy2pgKrVCpGvZCgEj30fV
6EuKqsHHS0smayJEJiKugQ6JWDkQCrWhcpyDv+HV7ANfaOzYtYfMliJvKoID/tiO
bqjKOlYdh5tYw8d1AQn3vliyykE4+moskAfHwHPfi+CtMf/sOHavNrCT7F0Yefq0
aTqKxZSbKbb6kX8kNhJkxso42ndmeAc4p5JA2wKOtmU9NcwESHhsFsa6h3VKfmXP
G0diu3lXp6krzS0qDrhJ5nOzBu7O60jTA5hkPONs1E8t3S0mZKgLNSL7aq6fUp8d
fgUeQfgYMMsUbXavcXBCUfQZOY4zwkkNkfDMSM7lQ4LgT3isgtuGwF511dVwcn06
I2EIM/2hfqZz5+LfCZDM5pmhHlrX1vIoCUt/2emdNYuKvIzU/6gfg0PgShMF4qRD
1uH4rERHxLoB/AuEzIoz9QylcLaSY3Vx6FN+R36EpVhOxb1MM8vx8PTLsdaI07SQ
JkIpGyrFnkE8XEpfHmC24hcdv1LDR0TfADursiBYs6kyrU4lhYd/lJHT/RXQQTJT
V2kxY9j3LWgas3l+S0U+74BB3MokVdJUsHJso6V+511UftdqDQers4hxJE9LLrtc
VC+0+msDEbIbNUOUsR2vhqSWWT72GuFEolsSU7eqIoE2WB6uJjBLlyVXkFIg56gR
W3uBWwEYNDvNtRz5z+Bw6MH0uR6LoreDOkdZxmCBKBWBGhXENszmPUJn1JJDvVXh
+DC4Rc7Ki3ksgUEvON4fHpYFfsaKn2Xrj8BIXuWR+hIg8JnWZRn1GdRYQsKxEGAl
t3qkiQJy93HbqnuVz8TSX6CsUu2slbpm3eSlUydq1aWiqAMsbgh6Bw1zCxoGkolS
LMDuQuaaWvYjAiLzVJ6VGOqCLgfBhnh0s6wOLI9LFEKesAd+kKbzzwpBv86KR0Re
QXcNqvnV4GQYToYSoZlLBoszrFbHpbUqLbeEf+b6sFrMVjqWWU2FZqUNCvEFLfTl
kmrz4AfTF1wjEgN07jWlVGgEX9dh5L4fU1+26E+0CeLK3dxZXOZq0nFmNO2WRLjp
+w+qs8zSzpdCVEDDiKKDh+2BMQghOmvz34k14RRnJv2a75h6eaUkNqJildWDF9DZ
px4Ix7z38GLWPadt0Bz+FijIbNn5de42fk9NDzRZEqrInzud+1DqemU7nIfnMjYe
4wwWO7v6jKaaFdcBOkBkAa/NUDCPOoTVDHflt4AFLbK/fN8k9sSw8nL+86Vhz+iz
VlvHKjMPfqVR/3KHvIBLuJ1rZEvSiIXtlYVljhQ7CvcnTsiPpRV5ufy+iWuyeCh7
zux6ktyGRfSWrcujWbCAis677dYjx0vrXImpflZXMWqqWKoAPRHVK6/PshBSLhKq

`pragma protect end_protected
