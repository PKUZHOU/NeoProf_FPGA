// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kJ+q/zWFtQWyJwu0Gg1l4QV6dDePYyPBSHZGpnHjV9J/Pon1fAObjwmJ1Eqe
x6hf5VhwWnq6Symj7PGWqKF2B2c62jbjb8q2hS0dx7+00FLj5q3FmbF9/3Tn
MJUqtD+Gsn49rTDzLYXqjQ79+3GYsrXYfxVnnFtZpKACg6hCq+eGlRXAV0Y/
tI4FNII4vYim3Yzt/YRRpOVNAiVTTxs/baBqk+pZre0OUdRU2F8AN8oq61rP
k68eSs3h7LnYayS3BM11rW77qh7TPDBDjgT+hC+5a+f//BXtnqhgGUI406Zl
6xAhOiSnd9xw4BpzQE+2Jo46/P4hD8raxr9AHpPTaw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
A4EZeVMiTPUw/vhO1pmGMNIOf03UmayPWVkQBMYGLV9yU6lC76O9+0onIj7Q
lB1TsxXP12LAOiGUljxmpoxNgcIscMjCBbnB1C0301MNOlb9+uUjPAkc1Bxn
f7FAwpfI7vjzBwvjP454SS8ZSkppAGszx5EiGPtpK3rXo6kmf2u06SCAk1Ay
yOSRnYmnyWQxFKXKoaDqsEDLcJEomfTyKkPvnkgJLjhcLW4Z9jr5xtkb4rkv
WkV3IFFV9DnI3gZppuvDI0jTAsPFPTvq+5MepJkRdxR3RGkZ5XymiA+CMD5D
xvZ6e+eMZduYefilDR/kpqNOkPhzr+Bz2BhfSKXlQg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bDJLSDkrcewSKUYKtaeG9us7xqoCdzKE/U4ih82wCHvizK3Vi2xEO9pugtjq
N1jObWHj2teY1XwqyOY0Ge5uDNUshVSB0S4DDTK2wqUKO49sH/RXeWfyAnVz
Qaftt6h5Gv8Jr3Tol8d/NamOnrW7z5rMv39Qq0rsSlBMkNorpfzAVjAbK0Cy
6Hye4VwhHT0OhjVLrxXRsMaafMf5Tmdl+8j07cU8PZAlsz1nsP+Tf7sKbiH8
oEml8WqTxo+ZGfqdvL3Vug5wQORh69SxGKa+CW4pfkUBOzeM9MfF/7qby+yT
Tj4gx6loj6k/7Y1Oc1QDaE7jJ/zUvQWVWIuQN7jiZg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
H4JtPXkvgSNk82uhF+9dt9s2IzxFHLeNb/6mS5qkXdUJ01q431llGi+s5a92
PNYAnGlhflzPVD3y1ieEfmAo7Dyw6D24y/wpZeFv4tCe72GI2dVeHtDKrXa7
sQjF0B+bMaKfUEdGTo+FwtBWOjU04CQQRI9IEZJshBnUA8kAqRQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
T13PpCDif5FwNrDWZ2NDPjK0vAieXDY0u4GgfczHneG9Ckcbvzwkj94CYFo1
+dMwyA+hfRF32mo2SBQvgNFKCROkRIAJEL0OY0JK4uXxj3yfiqPPAF4r1XLJ
cRiJUiQFwBVWWbjy5R//ey4fcJDa/fx56q8DjSHHfKEjDPCS3QM+A8RZNxpT
bY8+95zuFqE7CeW4V6sXdm42Lwd0rRPizLkgiWUW6k2tGZ1zqLjmuWrDNfJJ
+EPFO2Rr6dBza1KrTGiM78z+oiOkGCW0c7KqDguPL641qorWe/he0Maoj39j
Eb7Cnmv2/lbVMzc1iwz9NNBU86sOB+8GmCZLhQgfD/Wi9N28B+XNVMbcrTCq
98tcU+4h8wrPwp9HJvxpU1O5M6uGEbWpfo6uVbtcxN5YCdHotnn9vDVZ/KDs
/f5WgQW2j3lfhCyypbhgSBz0o8NgQebDnBx3+wyUkv2G7k8+sOM16Y+t3Mwo
9BaF91DAppoM0HwD5h2Rz3KqcxEtqPXD


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
NnCZViQ6ootg0tupEK5odhmaLO/1hKNINUb3oT1hzzv2Jkl0VwMO2vArH0Ie
phZl31TLHkUuhTt+lm/lCSeRL+Ay7RWc2wpIAaOoJIgN0aMhTZ+/pZfgR9Qd
aFi6eEKqw2Hj4bcxe/003DC3j3Q18/v0MqYb1oQCvbe5Ajwm8kg=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
oNVf4Wy/S7Z3D9h0GQ3EQTQytK9A36Xa6o9r0qsRqD+pRT4OHGcsXEaiOC3y
oclv5aXNeOBETYMqTkX3+Bd65JNMnkL/pbjQMWuHwJJ+MzajYokzkQ4rBjMQ
SiZdvVPDjICoJJPC8N5V/uXp+Yw+V7ws9Yj065kLoA8VSWTvIJw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 17552)
`pragma protect data_block
igdsG+nX1jibN7ONbjfs5Qo3+oUdnVzeVVIX8qGgPJjrB6kZoV+HbGl2bkDt
g9Fl9l4mLzQFPHY4kemP7Vv2fHlMXU6Qnn6l7mMsOa/NRl6ldRjL3er1chC/
75W1Kj0suABgjXlnmkCSqtqBD29gGturEyFDL89KgsgQ5B0vd9kpPHfs5kd3
BO4Z+4Xmk4E8PA0Cvv0dFgQ03+nTW43ZR5V9ZWS58pRniE3n857sAwZsFCiq
qwiAB1xX1VAYAqq3x7Gh4oY9HB5JA3GvJ4zDDNIjLdfwBfeS84Mv9RHFNJk/
J88AFhoGq36YrH374J0LQHZ03YTdPBgg01FjlmH4Wa6qlFFA0x5A92Y+VQw4
GV1nuNqZZs+BSENh+LYYuA0qYazCBC7cyfaQns9AeV1z/HslXCG68A2yZppQ
GGhmyzBKvfHk5ZOzdF75ImXUMZjGwllo7ywjRv0ndIxBltbuQ7mSMRaIKTxE
yLYZbNuEySUFjx2mBW38iwvFnlA7T3MhRiiFEFN5gf685nzoOhPLk15jS+IJ
ukibCwteHuZSujUw4pkeqRI5L0kabAq//mm58CuV+4qtpmdLmygy8W8TdyD6
LrynlTzMwDRfmpwAelhmc+dNNTiYjn8h/zdU0Qa8ibCy9Gwjdy078H3O7/Ft
/0DNcq+wTMCOE/GTIcK0vA5ICclPy8sWVj0VSbkThqUJvbeuSm/EaDrNxzVr
fTat3eQSc8vxs2+DASyIyOeoow1FeGVPKNT5ggQSicaCfBFrC9WjkXLWkjdU
fTbCmVBRl7pFijWJZ5UPBsRby/k/M03g+F4KE70mzTWLb/S79I9nQ2NhzNS3
MwtYwb611d2sUwYPAVcIj9FV7F1Uwu0ewWSywTdNwyY/XpwT/+H3SgDV7/FI
MS1v3bV3NhZH1R0e7A5ZJATDhZtuTYo1w64wzf3BG4hj4lXG3FkekjQzBLDB
1HxefsZvr/Uo4+JMWd8nvPpMqOCjGYu2DMIi12vgN7b1hY4cjBXJDazxjzWs
j+yibeT5jANCBH/BVFYsT4++V2XqOE6PREuIFzyQ65duUWmFWbBb2DzYz4sG
UBn2IixtaszcBEVgQ2TxfPOtV/7JL9UxIhEV1Ae/TrQcJ2S/bB0yfSGuhkZz
bdNIx5s1CbzmXmV8DtqQtX+i+QgBD1ywRjPIeNmC0qeJTzndtLaY4BU60BSX
hiHFggT4UKZ8qZh4ifm2IMXl+FRZJGZhhQIKHGLB5F17Q61LIlzM4JB3b2YV
+ahR5ILiyqm46AKkMUCeCfN93nMXAWShxoNZOXzRmsFzqaquCs8fL0L7mZNE
fsvBPry/RSpne39cx82j4M7+jXPMJytOgMtbYjbkwUMKO7cSO7Fh63mBXHX6
YzR88HV01CEBG4L2BeLvqhnjARdXYeEgbnpqFXRYlbZxINpYOW4BNUbfdjio
gHLem4Tlyc6Q3j66GMXNpDqMkAdbKECmitz2q/Gxnd+/TTG5Bd/X5ME9VfW7
ceqZkvgmDvcBVYobMdKqiqPOL3V6WZxO0UGu99um6kmd2UcpBMBa6GztaUdi
weMO8q/h7hWVP0/UGWZOpwEy2ANfhv+L0u0hJlOi/m1UFQIa5vvjQ3GOKxke
g/q6bY0ZtQQCTBNzAblZ8DR4kfqlqvWccC8py7iHNLFudaXX4UbGtSuevUiw
h9EkZrpLxOjORKNg4799hrkPARLGCd7SHDHb5LO4+koTRpiWBUU1geKHF94X
AwjWe06ZdT+MqyRWhyIbE6gPMCRNmRkidLZLuFLNF+Ny88X30AHQpE/AXaX9
ISiMBAaHOcDtCg0vWSinJJqkmk8pRBZ7jIaE/dm3zHJFJzfqq2I/4aNh284E
xeiGcnZwHJDdP4rF+cuSYBPeVCMLPrNx8FwS/2bRyl3hKmqTlp/T2uSGUYNT
/Q3P2LOF3mKogKEUNN5pMIKcsYAtr5HBcYeXTIlJa0GkY4Nkdyd71mS02ybh
4fhKLU4QiXxmem4lH0ygD852kU4F2id9rvyaaA4oseii1J+XwzM+EeO33qS2
EczgaqNUoMoboWp/oSJ/aH/LNAgw8kmklcP87kzaW5gJwx2LOklbf/5Ab5f4
zS57av8iik0MHmh03nlqNogUaC86wX65QbaxGeB0mvHTbTl5yNQaZtKTDMrn
PXBCNjrG1t4R5KKD1omi7+3GI2j9A5rboznn46pttZg8EDLXPkYjls6H28xC
5t1v8MjZeflwITQ1QsdOX6k1690DxKibVXJui3Ny+Q/QRTAskGdch+5SGnzG
BkvyhFuJX4JyHSTTmSKSAjQbDfyIGVpAbikZPQTtBd0J8f9JcQTk40cv2+bg
5FtCzfMZu+Kp0GI6AqB1xRzr0i6fynnQc8T/qL6zRfFcaYuphfsBzXDKuOMH
lLbzDzXO5wgau2XE6qwgxN5YSHJ3GlRVm/rQ/bYw3xvqhscxI6h3Z8aJllbu
Q3knAX1iYfuqqKOYwRNrDfyxcPSdLmv3NjEqWLtRQ3GtL6eqZkWJ7x+wGpsA
H9wH9Q7MJX+gNwF48WfeNtwZSmb4tcOTOPxabWZBFMN3HomPUA4M7Yl/d0u8
DppBlOWrchcrqGI2lmyn3xq3GK/REXfBxwosXxS6rGhDKNtyfrbeyrhYGZkW
Hit6gCwgZZsunox3/h80jzw74FnSHfOLlY23cm2jBFX3G0Hy4fkCZfU4dd4i
nABJn9jcyCdQvJ7ZO/pcCnKSHZDQ4Ot5Na9oUKHFAIamGPPbdO1JJbCLfo31
pUqjNRILTF7WVgn5dADQ/UBnMne80Oq/1OG6gSCGeinPb4xf7SsRBWA0ReRo
RQzsAia7CZ6YG/yptbNAFrV+SUyD04z4BhRx74BEOW6QlT30lJGef6EYhlij
JCUuWidC1h9+T/ZiNw0An/9MlAqhrdwougcRkyjkRnFMZH5BBkpwh2OyCDRa
Mh7PAJY7nAIXVma1WAYCEqD5hqc0TnzVr5jti60jtD55wL5YmZKqYF/U8v4W
sp/b0sIZ0/Krbibh6CohI8BNMhVjNpXNM2m/jCBWqnBAcO4rNvoGPQRgt9t0
IoaL+0otJjCm1YBWQUp6RIYPkl3HJFCz5Rr9z1NBU9Bf00YPkd/Mow92QOpn
eZIz0AkBeK3wzz9QZS48bmOJzJ+hk8py7MFa0uclmPRUTciSS4vSX1XVLyVK
FPi+Wxu1LjoD42JJY+KZBA43/EsgNrNPs+QdXpubsGMxDAfT02FVNiOLCV/0
vxsvGjG0ygNNsN6LX8G5/aoNLLK5ImXczkDBDpxw4n427XgcH++84UbSgQIS
YlnsohWFN1dNMUSa8IZyInTAu+tqw1TPwM/EChHIhuKBvnszSs7emv5MomwD
H8GfIQC8XB2864u7xGRZ5WSEW9Mc1wudgwBRlgEZ5NDe/dk+z6IaD+MWCM2x
4rkHmOPgoa+rCtyc4lyjZFJROfe8GQtuU2vCOGgLJBI69IJjL7m2Og/CWrTH
vrVoWN3XUqvU57qthBarcXVpBm1d9KFG4u3AKs373BkdgD9fMrWLYJhYxUgO
FCePCWeOh1QjRoSqbeM5RFGCMV9ZLiZVEdv5BFfrHeZhxe/ckIWBq6m3XR8p
BFeaxwOeb5rwn/2Y3V1DwsqPFEjFk/ebMBwtrEg4bXd0kz7zhozkWuBgy4zn
MU+O3gTHxUqSwwyMYyQztpCvq5rugKln69BN3393PQ0bjXzcjUK4eqLlAU4w
HgnEsBMVJfQ/tYBuWQkU0cs+7N4dgZuZXopDaEMnryvmtmHNmWkWXz+Xj7u6
M5SlcOIOoryFmPxvBa/U8CzZOrfMw9SNV0AAm6bGGsjb1zXqFN0Q6VAZ6daI
8fL3azX4UnrPEqg3LiY2KwwuCX1U0SyNCDNZS1HCL2xS6a6l8QYrbrdzD54d
fcQo5Ddy3EULS000fmzXrWoNpvNJP9lQ4p1Is4f30dhlZoXf0LnHvsuD7Ri6
asepWNa1mpaoKM0Tps6gz+ONiQ10TD1Yd2nUPa3qT1xypnMQ6qCZ8d3vMXtl
pDQABEzBPejW97qm0ETf0NdNCI2AAkNO/AC9SF+9+Y294WJj9jQGrZit1QPP
a5PnyoqIs+NtRqfZ0mcMcfLM7C/ksQ3FJHJsqeP8nD4+NrOnwBFqZGejkbkd
rBwEsi7JssF5Sg9rx8brriN+VGgm89CeI/DHvTJnXPcSJ7n3c3TzXqozSUTh
RG8oy14ee6VEOK1mkIBruGo1Yv+xp1EbvTEuOeTG6/lEVMVckJC/wrgi7Xv8
6zAJ2T5idwz765UQc0O8g6B8VFXtfQ5oJqLOghO2UEE110xLqUJjKnXgio4r
0ICo+K6Vo4c2meIcXCV8oeWIvjLVf6Fz6/FI9aHBTFvysoXaEm4iCWcU74Nj
DFTN+ZJa5HzJVpuNuXE3ejqAOgAqfSUDYYxoB+PJLG8YbWOJl61D8W2PsSwY
Swqk+cMj78oRCQMYOe8j4w7fyqRqrGEZ+hiyoyfdZw45wMY/9GNAUQ97wZmZ
KhKxQCG65KYNJvY+ZL3K1UmF4HMj3ROkth171K1U+VYgg0icY2TC1PJ3QMOW
QI9bQOjkMuEsVvoUCr6GP2tg2CHXuvn++D3Ls1/ARZpefaSFHZkVPGpVZ/kx
jVvfgXAExdu0KyPIdIiAFOWKcxkseVDfIilg8pbrqskF0fs5NaVaxq5d/oJn
fXfCmlD3Yl3Ugl9N2TSKAwLK2KXK2R/kaj2KN8brQFy3osJKC7LS8ncFxf9X
PHu3qWXDAXcPUBKeQ7QFtkkagNdaK+PGmYDnikGWXvPfYexJg5jrf9wB/4M2
+bAL2ZHz3/GQGM37Sh+uEPlPWbL47fWCjUu0mpxOox4i5Jz0N/O9ubVCcwRq
3av5jbCUpe7AcbpSkbMiPy0I1WQiNMl4ucMa5cWOGULgX3+OkCURbnqJb7nU
mTCWh6Uz4BvsD4L0PGBOtU2I/Z8+te74tJz7GofVC5bQPb4EzMalmmUL9Cx6
bZS1C2ADKWHeBqkImTjFY0C+BZmU3Qr8AwO5rfvUQpIOLLMevu2bN5Pk2rOc
16407FToudOgWUE3/GTRGhLBHH1ZBAxCJM7Tx5xM246Y/Cw10+YkAcA6H10A
dBdyhZk17FjQYmHEh4PzhNv2v2IrBRnZMjneL8AaLUxPY6sVv6js9YodSct2
RuO9WlMDIgfpkvaYjByCE3eW2vDFkR7e/2K3AjETAHAeloM+DiScqz81ckaD
B6M5tZrFpWwUY0aY1QLWERDR61U8V7v6pP8B1FO5SZFMH3ksQjFP6Ke+hplw
yd+rl/LRsm/NKqwZspPe5bycmSfRGoMz6gyGYDHtsKIQUqRhxlim0qEnGwd6
M1NgQZjeeO/biMYqi937nEmMfr1NdJetNEU4gD1k7sD0CIrEDMRtoCzX5tjr
Doxzoxrl9k4xGPKDAQEiptr6bqQhv7QF3uomrX7Clfvf8x0ABYue/VDJYXtk
ddK8oZqoM9sjzEETwB2QV11XvZ5Hv9XcnrxQFA/hBP636dWm6CAxpNbtoqiC
amaz9o4zwG3qOW53X+TcR7XIg1sKNu1C4f/Uxp/YmjA3eIfT3qVW5G4r8LNO
btFjlwnyT0OQgCex8l0OaIsofsZrBCMr59INGZCxWr1z/tTVHn2jLqlXCUGx
Oc0gdZLL9dwflJ7s9hVVizs6ZYv292KpoSBUwc43GV6EenVmt5XxaceuZ4sI
LQfvoI0CpHCUjL//4Pssk3fMvMaotZ/gJTzr05K4aXjkJxwThH8x7XldGTYA
WZ1oYipEWFFU/BG9TuK/2QfjwDzHwxJfXTdolqlGyg1Byru0GAlCnSB8O2St
JCfv1WvzfKwy+OFx5vPI1v9n6g85Ta+ZiSPCt02dR9Q8p1PITCRyks4EH6yu
FqEoAzEZBlTvsiJrlo49tvbSvGnCQZVzMlSwkRjrZJVqqj8c72PFB6FRo6kt
QLORdP7kNNQTQVwFpJMYYOdsJahtjz5j3YgFckZTcoK2UMY76PKUcQr5wOXj
y9QPkB9LHbt/e6euoSQMcAFV8a47j/UffvJ7GG1kUn2hodQE/EoJKMlXiDOJ
Z1e6jQYG/ys5brdqRC2MHNo5dA7hK2D9Lc1lXswqEYcXFqiIua0pqWJSkw9D
dwzb/wrgC9MClh7cMNV5XEOU4PYUHWb99bovPjYgi+41IvEILXXDCm51KWLP
VyopImduLYNAuWFI/Y/ecVrmiGq/epav4GecZMxpwtH6AsnOos2okBU2cPa3
VNIGOLaZE4tQ2qY7/RifWyU1DZcqY3COfHm0vtJhTQnyUYnIE5rc1e9td2xZ
A0bRjVRhNNrqapYnLkrcvevJneoWlEaLBatR/fbg1Bpn7dj15WiFHo1ueeX3
8HGOZQyNeIZJvf7zZK45AL6/3Or552P61ARAhkNygrit1uXWLVM92g6BK5b2
heT58Jg+1FpaWMh/BxVBdyRmFCAm7FqYJuUEnc1Rj1jj2TUTanNzXpPvlcvo
Jfm5H7/Z8pz7NS/ZbXIg/S9tnIZ2mWhcuMu0YUNAXgHl8W7Dq3FXCyFzyKy1
QBMgeDVUIvhTpjf5bSMCO58mMLpSJAzpDQmd5jok+KSpHxD103GXrgDgR1CS
i8ErYQyLTP9qlRfyKSJnXPM4iMDs9LRjBrpl7LW0pgdOcjEgUFfNzoNhdLA+
GqLeau8dzCKy58EAPN5XMDJlrnZ2C3LhqcE9AUj02REEZHcDYvRPnHMBmf0K
lZDiPZ6tGqWTW63Hz30kSIz3TZ6j3C+tyn6hJQe23iowLFBmtOf5/zwjB6Et
sG5M3Jj8yRdFBnGMG33ZSRC9Q0osJYxbs4FMH1aJOZCzEDwG4fYyL2apof+/
dQ57x8pCSMhx2EQE+1VomfX//gJYXfV5JdfUPZZGjs5RxUDd9kbmh1kGOQ4a
QIIe1X6YbYQ5Tg8g3xLypErUaM+3vwLKWmG+kmSVUff6zPvQWhp7YdU0xtau
LcXBhfQADgfurC189c1uUYELTIxJxvJdi8vhH4RAWgNpJ9G/TP4UC17qQaHw
iEZVeiH2m+LmEab8yW/o4vtiYl/jMT2H0mQWVmETdMZGsb5R5e78NIO+V5Op
VvuzGIJCHUyr07nIOOzFagG93AiBjQk/11Tpb19F9Ui1fKuxD4bZ4ceQU96V
yPWr3G6wcefLsN4Bo0HPf9uAab93Nso2KUXNhoq3Mc5g9uYkn8akbmSjggq8
lRGGh8cSjY52NO31nT4vVrOOPR62XyThhsrWVxbAWEJmWwJ5qdnwfqRj8HE1
CckxhnHRZoWz00ZLoVQPZzoRCTj5F9hbNnyPMqakaZESi50w+rlVoWSmzbdh
ltxG5mkbCRWk2MQiqmySAb0fEooRDF+tQlyFPn3mr/56eJ38t+S8UWNcE2z9
gEZ5N/1hWL0+r4cOFt3oKfvdaX1dyAqWbKqurZJkFr3OT+LP7YXIeN/ntG5j
g0xEVQQ6xwNlWVlpQg969q5kZ9K4OazjHyjwxMcakyr5hsxBZkNuxd898T3O
BeBj20Q9TU9EOloh9svDTRtu10n3Ehd3CqK3UEtaM/KesMxOjOzy0HbyUKn9
oGGEhsEN/42Dm5XPcZibA7xfjTV0N/uhcGa5dDHePiDMFldHSmhfUHlDkh8P
+yxtw40W2K1g35gmDRXdGY+kGFZBRd7pycP7BrZ4YszG88tHCZ/SXEGFs4Gu
xXvtzVJDy2loHXkzQlHxpntxRbdVPZmKTanR2TIChnA8b8wKx2J7zzwYyxrj
YN/5vER1julJ2PYc7l6pGJY7jxYcln4es39LvhlWDAa8E9ZZuwKFOWqiLlFp
Z1qnb1++fT9MbtUS3Ttwn83b0s+nRWjOEyJvvLLAe3lZSwyBhMjju6vgeeLr
fiLo/3eaCJua5knhUs/OkZtOwo3f/M+zzSALanNEf60JnUrFqog2xw03QlmG
pN2vXj9S5awEqCjxYGcBgTpvz2dspn6+0kdWlyW+13S7pMJG9XYkvNokizqQ
ZkIsILyhuuqVEsCqm5nqKgxF50wP50mJC2drAafPYe10mby1r+eJZByuYXvP
JuE/aH0q8adCqm0YKnB7v7JuO3O8WQWp6gAHFSKO+1FXdrQfCI15BlVJkl5O
pB7KJtWDtaadCURjSqW5rbvOc+tV3rXsFwDrAOS+OnCOMCIsdJNM57JWmF51
6gA3wLD6w3zDiCWBJMtXPhudzjTqhQ/DQoTw5w8c4AbcG4E/fbP/16rjfWC6
2Cl9eCshnlYjjjfNJThrFd4MOxgfheUSTSBk8WoECKxPDrtZWdHyWhWngNMX
RzPOtiA5R7+DZIGoSjKLzePl87GKa/MmqI9Sd1vw7xlBpiWNh4Ae5ceqaROR
YrACEAofy1XUGkHb/jb/G93W6diL5K3acHAW10OfcKjRzKIfjIF0k/hka3F+
WUrFJKYib41pLcluxUK53EoZ9f31ysjMWwNFb+1+b2twWaRGbCH0JhUivL9o
5oQtxH1g6qmI7GQVYNNdVJYgjjL2aHcNj5ctVqnqACjNGb4I+bhlo+AacmD4
BIkVH6kOPns2ktfULkk448ebgIGqgO23SB0PjSDFuNKEFdqlVjizFVnY+bXU
FIqsS8ww4QJxbyq/RIY4wE/R+YhinKyp8rcm/hocfjV4UjyEDjAKa6MJ5W1H
SFLtK5BvPSQWloimH5aCPKnQ66+xwH/BioemRHS4e19CSUHNTTd1TQqtf2ix
LiC1IQPMOljO9aLgWLQaOwI6Oqki9x0rX7vr/WSXqKlqRJZyt7+C3flrF3D6
cSZ2ikrEjY/xQuUHn6q3ZPQpJ8vBgCWZpY9uRwgTAdXilOsA4S6UACMKetvA
RdUSrFlt+hayFXjRjTktCUlDzrX89Ujg6Bye27YRZS8N0M8VS6//s6UkAYFM
A9gKsdfmhOymGrSgU+RdRFMryk4jzsHVlVdAzMidZo5emduHD5oftFfGEDtT
ioS1n97k6O3G75B7J2sYSPRDi6Ww3lEJqByl5F8LHi5DCtk3ZA9GhP7gDjx4
vCZVSDewnYOH817eFfOgNe/l3RsW0YIlmzzNt+dhtfLT1DAf8uQn3hfRs5D1
BiFCQA+ok1Xxb8S1h3uc2uNWH2dZr4J3StT/Sxr/k9Zn9x95flNTwRgulWEu
FB5Fr/XZO3w5HXBEvsjnkZhFT6syzU+LKoSM0E8noulYUvkPrvzb+i0oVTcz
hr/4N6DWIGgwtsWRlZF5pM8sKJOgzQYf7p0kQZZd9SVmAO7VfiGZzqA/FlUz
vUarhxp0peyxpeHH7iQQAjIUWKPcrqwuCWAIq8oe89RdBVJtbHTQ+XhpjfID
z5y7YzVFDekPjGezULem5FDvF8jXQl2TljUogcChippjyVJe5CM3CcF6r6ui
P5vwuJLmFDGwBWszun6Q2F+/3aAhZUCZXgAbQc29pnulrcPQYHZA1OCcqGsJ
d/a/2P6xuZiMkuWwdEz/+l9Wz/QdKeb4WeUNEOCslm3YKqWP17N5DX5ujGit
7XLUN6vcIgf0b6AlrZAKX1UsbN7jRsGL4rIVD3EZpeZ/1tWh3b0+l2P7a/XD
7ph0TlnU59HVBusXoTtjETpZhB4zC8AvaIegitjYfj5OgAnFiEFCGsvOMQzI
W/1w+FpQjZvroRUBPWNRv5X40GcXpLEHLmAdrvIgcyhycelGHmTLWs6XzPyw
XBSvuzFtS7V3Puj1oHH1SCNitGd+YIsTKqqf1SioUnGkk0AQQESzlCaeS2Kl
mQUw5Xqztuk4VF69RSk+bFfaLJEzfgttZ7oUOjkLlGHM++QRGKATkPa6pCJD
2fFrisBMcgL8EcjFH2YfJdimG8zFoFPlJEsCMVmQuwIg3AziSlC01oO4fNfP
535OsHdJQ6SKaWpmVnh7AAvknp9ATO/zFkE3X95vQA/E13gXtKlkTvccbnKy
zWTA01lr3du0zkSnFbYf5Vbb1a/s6W0KaBVw0YfxwSyj/AMr15EG6Y//A5M7
b+lSQ/R++0jCk6ZCHczac/2lxvzMy1+J+Y3uNrg2qxfRHmYipr4RQdL/z9BX
8qsr5At0rnKoPV9Q8TI5uthz1k69bWgBnX9O8szJ0ZcqChVWp1fGJXR/DpQ0
BftwDbCd/loD0NPlI2mfC/NLiQ2g1kZRgK70FEsJE+5EpzLMKFitetNMBtHq
wAzmtwXLMQELms+Z5xYy8rFzYVNp7/2ZYTeBfH4eo/K0pxG5JibjUeaDkRYy
keGHoBN3EeGA9Xtv61SZ9uaJiA2GlEEby+dxcYDp9gMd4HYaIPYIOgLaVpCM
KhNc5IHW7VumELNwDuc4lCIgqrvlD1dsXw0MbYC90te2wTEYAR/YVsi5aLbo
DY00EyjvdrT9cseMeBhSW16euaC6l3eKlqr5+JaMez1uexRLrgPB6ZYky6wN
pLbEbzS9xnlEWKrTtrQf/w/TTRIubANbjswB0wzcjGHfzUQPue3iA7Xxfbkt
9Aocn8O1a2dPVUxOyAEn899pc0XPIztnmK/9a+A84v1+ZGm3W8KVS4X0oh+O
HscpF/rj1dzBMUalyp3Rk7TLRZ7X+TW7zn7cfGgQQ+AEubbRZ7sSrJa3ZUDW
p9omxlgziBtlmTfVPuiSTniE1tfuz+Uu+ZwjtKrBlW4zYV3RuBt/dt6qgPI9
yH3/vbdBg14BLE2YItVKD+iD1ppj38oxxak7bHQivhZb7SQcfv380HduXH/T
nDYaXgke2hxhH2ccpt64pJZapN3OJ0xu7gYug0fFUtjiWSDozqvDTZ4/xCBB
rJNvndmOrDIO81YaDUTW6qcNa8FFrY+p4OntX410rL/51m8z7FO6wfUpd5uD
ZkgMUSdF8Q300orE0EgGjF8s4S8wU/1aXKEVMyjjL/8KOy5Y0DD8Gcp2LAEH
FeZxrih1fDrWzaCc4bDPUoBT+TJdBKQoHAz0T67ynXTJ/469q7b5190vyQu8
P1yxvrDkcOD8KYP1OQPN3nCUO+kVzpl+pz56zl5uKutfz3vmI0cwteEh4Nqj
HYdOiKQmk5bUXcyVKcWu/1cOc/f4Eattnu3gXSgRCfrkPy7lpXDNLTNovtyw
QEnLKtmzKyhyniioR6fEQSa7JbJhgfyfJnlvvaXq4NX6pN49//YK8kCedQuJ
EYbQZaxKkFcYALYxBDssVRgQ5icZsos+AIMppI8Cq7UeoY8uaFvHWZtUpm4g
zs6adz4kwYMd9eEvMCQwpWysxsIM8VSOFRNYfKtebSVWnOI9u3B/4gJxixn4
NhtOh0Wld/0P5+aDvj1Iz03hjquIz8I3gGg7BoYl30e8f8wbxkmMl23aTX/y
qozqx9hTWRKd53E+2g1UQH0tSa5DmVze3BpPUGcEzUvBV0cq+COdfC2lNLow
R2dPvkAFRyH1VXMrKEvELbr/MuJ170sqpbaBK2xrruBpYjjJOsEFygOQhMV+
GdqDGo/g93qk6CK/SSNbvV5XWaI8g0cFJk2U8aWMtjcLkvq2fuH5coKQ7R5T
l6mNtnNiY1iqL/buUYKH591r8NRU1JSJlvh5CVWthBtYa0LJshR+Z6SNdfrc
aP5B93JpxOXatziVW7+kSue6kjWQtHxmqKHCNvObwgv4Zgb8ZZGYnIGfTBzx
yfY2h+HqEHfpayhPyiCexF5i/sZqjlQilrN1XdUFFmSVblrF305C2i9VM4f8
MIvk9ygMnc3hyQxnmkY8C++DKmLKXyf4vU7OgjSBi1P3+pxO/8WUbs880aG1
5Wz+qd6gIrvJFwPXcHOQojt+qy9Nay+yj9XMooD2OiaD4sfsNTVxowqjWAUz
QAAo2s8JAVQ+Alet2CHaEvLfzo//o+hsIzOwG6GvYq/HRj0zmwIj5XQx9H/t
vSAtbiOBiitKv/60xJSD7PjjBFE2Hr2q8oj4Fe452Ol66a5axQJeIoVx0rej
/vajMifuKm8/D59bSm+UzC4+xMe2X2b+1Vve1H0NPkv+tdcj12BR8uvh0l/+
RcS8bCDylWDdTTq6olfh2UkdaIpzc3ipP2WtuGEwLvGykQ0LBj5rpKV7WF67
i66prIf9siICt15FCNuNOwtGtcAZtDT25Wy2Jn8I/wVKBhVOfwujqUVMIOkH
S/yE5fLd2vN/cC6aLarPRMRfQ/NCNtzcJwBRFEg+tOy4WzKjO2gxblXbyXf/
BNmTiYVKQKdCJNc/ORvwiOP0yGwdqmBk4cX4+0zNlf6ssUaR/AB3sJ/S1qRR
5jBbimFZojM7+H/a7PbjRjFfCm3uY6/WdzyLhvQnoZp+DDpwZ6/yYiGvm+ST
Qyugu5rBBRXHh2Lg/3RjqhKLdB/3I/RGVlcWuN8wwfLHH33KMnQ+QBVNUouE
+GdqVBBDd9P5jxlQ6pkYKzZQY6601i37tmD5rN1vUEQirpHCBbab0rJk+wCD
C3++MCfLkdF0vIoQ2jAk0nCBSE3DTLEkavo4ProA1TvMrsV06uqC6CG6hMRH
+u7FY0eGPXp+R87CmmykluW6tV0ZwnVhzIOyuuWKoQ9524P2mhe01QvgKcAa
C4YKKc3Rg9tBspZiurLVMgTpbcMTi+u75ZWZgLHVaLpMNT6sUYSjb5lWa5He
mrC9K4hwIbUa74/2BXgket4MrvZyYMPgJHHQC3ZHP+Dds/Cet4ziBjX0h7hu
GhUAwQu4y59g+NumH4Ymt35jbRe4NiKJLy3HVBL0qNosyPde8nIw1XMQ0V4U
cFM5Le5QbAaBdvJisD2RSdJpuxP+xz3338/Fqt3YjLEH8qKpYFXtB+RoydFI
nE/Pqin84SWidCHupfL5EZ1SYuIAHfzdKrCulA1OiVCg1TtEO1cFym2aEvMy
VUAeOZqTh8Yb2bIRE5uQaOZIxl7WXMulc71nNlz4eTpT+AtmyuyA8AWu5g3m
RSZVmSAAp5AC2u3Zp397pOJ6zMlVH9eh761SxlwCwbhxHNWknrPgZODALbn6
UstNKE88qFIBzJPCSbEmwutmC3IBhM8XQXu8L9uVgGu6o2O7x0KCGZ9iUH40
qoSVcKnNbkNaTgAPqNDfo5U+etJw7WWbp5Tgn28v1JRrVXtkakwKcrHWechG
1dUjarM7DFTyyOOrMhD9LiP4TOFbdeOjCIihxvvCL7Ka5lEj0K9/07XtCVLh
44eECmWKz9YEX3WKucuZxC56NQXCytKMZjj/z2Ac/Vgf34AnAa0TtMjOqzBv
Xfh9HckA9ha4Wg6PAJ23/5825bTkutAnph3Mpv/KyrnrUaVdX43IQHrKA0t/
GrgQ9DSpYiAI7694Y83O6kgzqtMMPPROYNihC2ZNb+GIWHMMbXGQ5IMHfTSh
FZS3/7cFv0MLBOgr8A57oPpijIhvD4OjxxIR7bs0Xu7o8+aMBLqt4K31wlH4
b0Ov5xFsM5nfCKi0L9ulcOzV7NrcfZfNX4+lyAZ6LayuRu0VCXk69dvdh98K
kcqzHpy+Dg/hGxWqcHNJJVZoiPbzXuODzAMg4lXJl4QGUqv9KR5OaP1fbDa/
VownDoUjIR5rZ4d1x1L90OJFvH0HZGjByd7rZVhgH6/M4uexjVVki2Icol1L
XA3su9yR1QVAh6wVRBHTAByjn0tQiUA278yTQmbkjkNtUOUXLi2in9bjFt4c
SWCGryhyqrrLHpfwjrZBciN8ZAUHzbxaob137ajQUxJeCVq/u7GyWOcEwo8y
4ThZ+uWmjv1FkIkubnpJYmr4ofBtiyN8PYLTQwEZ/XhynxQFNwI35+Ks+7et
nqx7Kpkq9wJb8mdVgnk+wsp0ctBZgJL4ir60MR4lTfKu9lbyXASRQXhJUfCA
Qedka4gvIZBPHXRacLyGNqZfYV0wV/ftoamU/qU4SUsEDhlGYok2hqYNQcYu
cL6qwEyFe5Jh/rH+B/ZcdW/1Anj5TZwC+TfGHkCgpcEr6hltuhF2CwVXvBAO
38cCEVCUnxtWLqG9ms1MujYJplMWS9h2rprMeuIHEVXs/qrvLBRxRudrrbPS
uL4qEF7NV61imIpMMtWCrqYYoFF8KtRsvCcLrzRZVKP+AnXHICn6jQAaW/0A
LkM9w6cCRGj3UAP8hd6QtAbg2v1RhtqCKvx27jU0+fJM6/UeM0pRZmR0rYVO
fbMwW2Wrm6dtMAhEIO+NUVBYswwXYIXErQpTBK3fEIrArwgGFnOkXVCokwRt
XgyMv8IyfR+j1ihHe/P4YMe4gvxphszDbBEbMfpKdteo4LoOxzvJ13XPNe4Y
vB5pDiaPeDq2IfzswMjRGFEIfxiT3ELJugKcOQuMiSBwOD9CZ09Qh1kx/FFE
+apRINXwcXCQZWy5MBCmUaouOue3ItZ2q694DUOgEIfxfqdUoBIhprGSyu+P
EZzCyA0efxHaSOPlFGq5/XKoc9aSJYeYDQZVnTFi6gGhnQG/in+SbRIepdJ8
+MqPKm2NZve8U0LYP5Yy6GR09uP++56PaM5Aq+kGBpDlsNppriKqE7ZhDZai
wkzylWKAam7wm7o43K/EEKZs9DUGp0wXnOraA3esC1ERK2fFbR6sqskbRbIP
irhrQrbJ/Dw/YtkwCoWAjvtLYt0u1txaA+Z5zDV+VjfTCHPsYKrcOZD0F/Lb
AZmQT+23Hxj9WdCD6YsFS/Eym8z1IyGCxSRB9f0o14GYPPhPeUOhacywA76A
HrYL5jQzzyIZj1ip3OUDBbuBpd8x0PG8pPbq/8H/WPxW2a3Ag134KWkBlh2u
DMZT4ZvuomqQYm+4etNNWwnZDinhxKYP3Kgcvuk2efiGaHl6TuNCDBBRovlF
oNTnJICdhVc3y/N7Ald7SISq8flyIi+iLTZwvjxNcMtFpr7d2h30OUYMDsKt
/JPXiClySZ/ZdYioTDzbZpt13zORtzlvCT9nA6LpfdBzP75/MrcF2iDpKr4f
gcb0Jdj0wtXVimdyNmbhDL+n347dFqulmBUO9VV0P/4XQPsYIU3AJab3YWgz
1aQvSloyYUIkJ883BO+mjFFxXBShkvy+9ckF5n+LgvKxZEFeOQ/yHCBJkihg
0uK+42jKAqCW9u01BxHLqlazF9inGik5JVNwuQrkT4R4oHHIDLGa/0F8oP+j
eqdn4BTLUJ1JKmGUwnoTcoo5m8ah2E3ifQ4PsNIHk99XK278HMfjGyzj5ldn
2O7trEiqWeJcmlJwcIa9Jt/ZfGAEZnn2x4BYXLFKYd5VxXN+KhgxwQ0ZvPIs
+6Pyus0RJbIX6wdI8fR2k/840P4q3aPOUm2jNApaA5NFXN0fhYvn44DKa/ap
OpEnQo6tIhtFoIIEFs9crlAeT92XKurRmea8TcEcK0nccDEeJ2vwepW3IIqr
Zy7WeFjDXC/rJUTRbEb9tuDSYPRLcVgiO8qMRc9dIVfibfoMYu7lwQJrXG3B
Tjlhjcq2vVavkHDoECbpvXnCBo8Epd3/0trns7iISebj9bcN6jMr0fy//+t8
8rsVdARHlmUpgByj753DthM6M3ZCx6MbKxNG3JDUqirUnfLrsV9/KhKMJUmB
1HvIbuPZXhjwqyJ2ZawNgC5Iz0BxUhJrpztvKlW5+1II+GrDIWV/ZQBMfpiI
TZyD0SppXQm4ICVddfW8901XvObnz75nZqJeKX/lbSvyo0mcvjRTu2bHmiLY
PsekLvY1FAsGXwtHfgiHtIOUY1eGxisxJ5OZiPZo6+4nd+xKfZwAqOkxTjCH
zJephBDvHSM6FhYstzJxU4LVoFdvWrW92VmoXphKfOpnYAeMR3tQ4Fpm8XOz
Jv+ZdteWJrHjGA0K9Ie/z16oNvdDzmss/WlrMTX7iyYvBmsmW6lb5j7Z7Qqm
EQvfzILlL0uwLgHZlgum3JLKMEOllka8f8V64YCLV6X22hYIcafG/aTV2L2f
+KE6PQvqGmcbAV0YJHPS5kaTbjePvAQh4TzAffR2sNoT6/941MUpk7L6xJAf
yC9+Ynrz+PmgyFt+hFTfgqT3G3vhC44wUpgHaQtVQUgb0WLkl/1JEDqAnxxu
vuusYcwmwnyWjS9sKEWhgqFO63r3fzLhbn64HR5lE7rkHRbVME8+tRgYxRjf
2qBV/5KA0wc0rKVPjLXrxS8Q4orKdpBhg8/egJ1ikgNu9uI2w9hhZGxE2KdY
DapLEWKYEoJD/yyGvQeP8BLeGoSMjx54tF/VspzQ5YAliz4pKxVSMWwpIPRG
ATLghq1et1e8aaMCUfeVqBCbHSVAPxXmgZVsiYhSmQ+HPf+5UI6PXwH8oSJz
nojaatl6wEFOcJPu9FUmTdmweqBGF1eut6ppcLQRZYP7wf1zPphFx+prOsFs
RiV+D39naEXAwvNRxd8ehaigy+9OtwyU+eiGg2fDJzrC2ZYV2YfdVhXcPtaf
P0SbwJ6UyEl+wQB/TkGtRDQpe4TwlKlta73FE641i8zN871YQMs9Qa4VgoCJ
+F8wo0c04LTSIYieNnd2AIYTXf1hw53bAOJ7w3gSX+rjqdIXr4/k9043JRtL
j0zaaVFpjIOvXoCgutZV7t5d90ePgsSROm8NVCo+uYMiJxrp+dLJcDDjscCZ
QNoLO/695j1DgFF2i7UNbqWHthzCm4ZrbGxq4Cl8rWyG1z8JZwEmNGbaO78R
nPL09bopUpRhHKMQSY/zDG8cJrWZSpeAjLmbxxcLml7CmOfwuEMrtTNjBRFm
mvJCcXvIIOCN3dWTJT8dv8DYLdj7KhVU1NLZ9lW40/FqPuq2ig7mfZQ8eQzH
80eBoKIDCIV9A9eu4aDhYYdN8Pfxmoxygpqk2kW7OVL2zseOwS7L0z9yAiHH
hjCgDyUhenZiE+7A9svrL4JYepmcLRJy5KZ2yjWv8y1ihXX1LytlUili+bKz
SHocCygusGpbqjWvF+C1Wc7OjFZ886c9doMltNSWudjEcBTIgW64VykauC7Y
Vlm719z3XYa+5HGKYaOpYc+vo7+sv+sTUMZVR6BkPT0FyvTRG0zxmcHwEsui
2JMCoXddXsENc0fklnj3cJYws2mCGRcIaiYVC/Aa4nOp5V+RvtthiLHVYen0
jqc2m6XFMvs74TMqejIRCU2du9Ldj+KUAyEWH/KLqxYX7GlFyYD2BA32QuXv
ujR5sON5mqVh8UcoxyO0bJXNZGMEdRLFhfdX9VmlgSZJlIuyFYx7Jz1TTq5B
QFvjAg2rs0ajsCTdIJk4XJ+R/xGe98sFm/s+4BAJF8tECWHBKY8CsN7N+0to
ReyjK2gDn8xhXC8aGzfcFICTwrTd0kFq6hSCY/PT3aK4jhdwoSn5BnLnU5kn
Hs1HsxXz/v1E37TVC1Iflh80QqyT7oESy9DiWFhrjUZ3Xdbh89+uBwBeZrkX
2kTa37GJQqzP1vJzOLUFlRjolsAbTMiL+wPCTopuXda+0fP9dNHojR7Cts1z
ObVeRG3yZJAJjXp13zLbclXSZe3nvG0u+fkjUNc+j+d6yvRRK6HildRxKPw1
+Nu+X7oR+Hh9Pd7yfZuZsXfhvfQBemav1JEQ4+Z3gYhAmn+QKhJgsYiXU8j1
Pqv2hn0Re4KnnVjOVGQdPO2mx0F5BRLNSVZPoeJrfylBVSmy4v5Pm+gUjy3t
Zkb+ivUJeBBjNFpiF7CZ9I/aON0svLJFgcbBkXw3IPsogropdWddAwGpHJu5
qUCqfrBOhsirA26mbj80DPhxjJ0Y+y7EVT0b3HKtl6tTW990QoqT/Ahvsld5
pwq+6/eP7QJWcHd/zHeMGzE7E7uWJX0gSVfEro2Txy2XZqM5D7TaD3/wpFgP
gBKRpOe7JD9z29pXggXug7prfL4gUUSBfDQAsklsBud/IFLOcb/9slXbyUq8
7GcRcU4Bwe494+TDZIJmPdhp5RoOixpAg3QtkEK0xi0428PKClqqJ9WYaL7u
OYsChfWUqpWcNODYbBembfo340N1SFn0PkungpSeDpGFUUkYOtc7U767IeSD
XlYnJOP98Z4noxigCEwYNMlWCgHSb0NdiBjTWVZMJPYU281So16gNcqs6aiZ
7RjaUVrEOWJqyqMcXG6hgN/wg8yg5WtvD7gEvElkx3dRRQQTH6IyvxL+yOgy
THY6sGE7kIa4bXKKsQ4gOtTvMFwjQvoXqL8VMVJJ77YI9wii/vb+QrmgDXG5
CELgHsynyxyfLnvHMKl+R4BoTJRl4o9Y4Mzwty3KnLX/vE9sMeyTYSw6KemZ
CbL5ySONlL8OVTh4yDxSzA19M/1YGfgZ47am4o0EMC2mo08Iv3KEUvA04xx9
Sy4loatq6qLA0QnwD/P8I6lOPsWaU4IB4/ESJKYH9A44f23Sik1TcY4H0Sdu
6tVzzAaHN2hWsOy6b/jeaRb4TMP8w0scK2djpY4UTvRUDQRjukYrHlNhB/uL
UDLrcL8TrGmlVkpTYEFeBPiuZcIr2n/V2UJwS17mpNdN1ft+mRQUAotVgiCa
fn4SAkcnUwRT7d9JT/iiwszWBRu581H9H20To3FwQBUsSxWqLmkcoXYWdq9i
vlT4nETkSBKNGG1Wpn4QvdjrPYseDDPkUUuJP+8HEPtUlzqZjKWxif1wMLqT
7u9U9nPf9GWfb0TWK+pLem0uRFXCWVzn9AbQjPb4W+xxRfxUIE4jh/uQbWvX
Hw8lJZvo24dvOeUlxYEjCfWtgoM8HZqSl9v8aH43sXJQBZRA2H0efRwkzWlK
tAcCfWNo7deSemnLpa2HwpkR5uQBYfyXf6NbADRYAWjnPyPJYu4ge+v7rPeW
Kgzp7xHlPKtOnr7QtXUF8fB1lgq2X3CNu3c1AsXyalBKYraGo2xJmxBzsE7c
n9/yQxSeKDu9nMCslL2PaXYt53s5NA5LgB88L7TNoBQbnSObShzdfFHE0MjL
79IiHE8bpa5Q+DzzXs7byeCWU2nXdXKc7BOhwSsvVROEtgTx4zpRxb/ny8YX
VUh8N4AtgI39irR/DbfiiYFk3Fx8hwFq0ltnDW4T4CU0HUBdytfMcTl2OQCh
SGuUvtXqLg6ISk5vX/3ipoyUUOT3GQSUGPMbGQAMKJUkhHBgLrCI+8ZHWbE7
HUx1Ci5zkbU1DUa7Zg1X2f7DoqokFdyeVZjBOKMvU1Cd3s5IHoxHB+DacFIq
ZRGRgtvfpWtdF3ptJ46is+w2bJm4gLwhykfHrS3Y0tI8Re48xTJdgZfQvF24
WiMXCLzqbpbboBoHpg3oTUHeXQ8jpdtYb8jPSgviZBThnWOBO3BQTxEaega+
lMzc+MO79HCoeVZgpNONbq/LhlFUQobv1dnxZq5vimv8Z8+mRGP88IVExCGD
nFrRjP1sSgIjOHdd4MbWz7/DfrJXQfd+tFV3zrVVU7mxkA6eFoN8bZZC2hTz
ln2H06y8IClUbBi6KR+V9bNvg8S00/8UlT7u2wc0hSn3sap56VQ1UJH+TVSw
xm+BFp2WBrsxKh2WDF92rAgNHmFZSu2g///LD4QmSN8IlamL77JC8Mmq+IW0
yR53mlt35U2eAE55SstFu8VJSv2sFuRLctqsXpcNDFKbFDebQDG9AbtJ+yzo
UIXk8pAlidC3ckaeTtIuPPByye4ZOZI87/BfW4y8EBkl+Aykc4KjLp8RoJpj
9KcF+BHCOaDtH+9b+thxYpJCaehWrCsK+sKc+bhMrSr2ehl7Ph/pFvoiHWwe
Zmd+w66vF8Jvk/LTCL52nZbiGMHcvzMYZH/n2FZZUfQmMjJkWbC8I8uqY1+3
greXZq0xlpv7Rrip+OMZA0n8iIV4vxqqVUyh93KhwQ69+80sRl/hgELFwmBJ
D2Z8h43WP6ZHaJMRu/V/DND4fH14WyeEgIAlIqf5rTFzT3bD9JALy37fqt/C
ScjL/nvPtHhuIssBp/zzOY2w/5fhE4Ci+Qo5oD0ua6NV9BjB/gTAH2bEhWvV
UONmhXNhFJJ0XDBWku8pFNxhvarUraeIfXGVA9iB/fycwsvdLBWi7B0fg1RH
GTv++yekl2gusr0cX33JXPCP5g48hScvGkdmv4YtRVAIZfwghrn7YpwgCzcn
m4+gKhlNczRShJobEtOIrYh7iwCKp83oV9Vxzm91b7q79yX0wjeIrTbV8Buq
7xWdfOtUHjjCOKbvykBAAsVdso1aBejJXy1Szcsu2B8Qrzv/OrwNSso2TO2J
kI74ZTBcMGwfy/bm15TWRvRE4u4N209Knd2i1eK5M0i2SL5IJ87mow7410H5
ST+GTs4shF3IqhvrCvqtDuLDZFahSv2pB53l3BGhveLrYYXu9RNJTcNFzb32
zRWmuaAggFNAD6CxiRdLjcW6eDOWq7uh4ZG1lAm/UJvjGFh/dMsSX+qg+OWY
tRjt12YE9kG2HCZSXFrtUwj9qvbZsCKccSPcYidrJ1gweKEWz9PCos3TNj7R
CQkn0jFjhNqbd8IyQIQMTNZ1Iakunmjlvy6UWQ1Xba4nhLiOIJ10qTOZZ+vj
Hw8AuZtLPNTCEyJAeK5RNLN6rg+5wb2kINBeOB55eiV9sjmV/Y8Po0FlmpV7
y/mpbq5XWokwipNaeGzHn7HMxbhTbGSfYVWtOL/apqaML8/smLA9QOlCNpqa
eXpFkbVQq+TdCid0cNKrd+TsyOLqcDTjvgIMyaJ9zEyVM91bG4Q3HHBJxCoE
2uEwGJT9iTxFHHg5ZPOBNwFQktbXDlnrlqeInM+G1Bnhsw7tIu0JTo1SeMNg
I/Jixwal+tKB0Il+5qlJFBGLtYK6K3rdCZX7QDFiU/o0NG/XYkYKQs9CwjPZ
BOcEOS9BJLJlTWcPRoDY3L3TCLpL4WzCWW6NQMoZwsreZif4tSe748zwfcNd
iufkd8ktl3tzhjV4l7/wkgArjyLwVJmdeHEXRR+TOS5zsPh+Kn4TEUXHAfkJ
LAmrPlftiNEy2ZIIBRF2t7k3JGIhX5gm+eDcpCQRi0fiIK6NzjLlGb2bmLxG
g0xsP/nXN6yNs9RpYAjXIMCG43rErm+yM9tozU7b0KPBGCMx31ydGr6kkHbC
EVOIj+6CebfQg0bx04EnLhBSMfDPc8ETowFl3qiLbjIWZuFl7PBGyltXth7+
rUwhY79nIa97f1gGcLQgJu7fCHKetSxLFo8jMktjk3j8rua+G6MHBjOFhfx0
rVyrdTJQbGZXpVOi7ZsYsi9XcIJQthYsnJcFeG9kmFdZtm+JwjiGA1QveY+Z
i8euj0cO7WkHhPrqqfP70M5Zmh+AlpwCVsJmUKUC0THnolUFH7Vd2/tI1GIJ
lWaj342+TF+ah5sPVAlOOznXmLniEehOatrZPWKMCj4hXxDsCF1oUcrWc+tg
C4DP10A+FOPzjLODVcuEoM5COTRgq8//yOodPyOJrQd0nQW9NUwx1idn6W7f
pvZ8mZlrAnB/FOxdSG8mVU9pqpjjmPSYF4yiZf1nOJKEV/mkLKEMXnAGHlR/
WMrKwO3RO29HjoMH7PClvgEsxAn0HeJn8tz2V8eoOSdveQF0a20sYT3hltpK
rxVqCoeWQLpWqiQnCf5rR22P6qrQfc84NxAeUzJo/xsgL1MJtt/sP6KMPyAv
scho8OmVCHp76uR6i7wl8AmLLPN1A98G17W+n+gcdk8d2NI6e5B3TocFGVzy
lV+YOi29kqutthpMdHuhYFnrTqOZexSfzS3fsoYdDEUl+AaL2dD21b3HCFV4
pRiBG4h1fxuIW6pGhURRfswADpw2hY7vuj/HexMrmSh0tYTsfcuxT7oAGRQK
nWQMRVkxZjqDsAT3u3RAiOTRhCwjqPcoTzUlb/6p73vXaXTOUqO50xFQbJ+o
bc4iZCaracSUs4Enr26NpHxKn4i1ZajkyfeuUQQVYIebIna+8Wausm8uAtoy
MXTJkTx/fRGhqRvbrfHM4KEBj2HLCmH/Kr95DgaE4/C7hbldsxdQ36mPfCke
ZJt44l7WNepSaai7cDkKZ147QUdj8LS9Ce/SJxLhL6MAdkPNAxGoWwJUYlJa
PF6TzpxAgNKLuBK8kjnuYOp8Ia6A+Cf8Rm+lTRN5cNPgOg8iWEYSChd/f2jR
47x0i6QXng4tYjWgVfvFgckMiOBKXMrfLj3bfOKvuBoDKHyqt4APzmsu2Icd
e+q+lIZv3bCDbRJf1WhUZnep237e6YQXTAV2zrRoolOZPYyIPZcc6jN7ruco
RIRAU+J+PmvbyspkLr4nHMq83+A6K8Jn5uwFlOBL5Ys3wSHd5s1EbdeRpQzy
c2GZodnVOrnHFC3yChwkwTnsxZ/qvH47+WbWJdIUu26tmde/eKyND6ZCm4wX
k+rV6VwKqSC97J03TUdKfE5ijgwA514tc7NoqTZF1ylNhJdpLczql8/e5Ahj
yfDH5mYgzFBC+eEVxZmusSmX+1nDOoSDo8KjPb5cwcEDC7lFy6FFzbYB9s88
lgtGn5wG4N3lvCLehB3R7Ht3m4ph0CIQ/3ZEEmiX3wuWHR3zZGsz4eOyuJPN
u/Y4E4WUbHDnIC581DeeKtpOZJUdlVqNNV6TsGPYkiXgKm6jszX1A6C2Kzpj
wRxc6zh8TE7dNtMqRShliyrKRYNMQ70wkfr3KJwgMKrcUidpGU1qAZvc1n1r
GEjzw3+SkoXEEncugSWQxMbJZkKOLV03b6pXqnfotCn9bV/FElVkN4U0K664
c6Uea7TFn8x7ondk0oeNFTFFkyZDGJghxpMRRhUj8ooH5rCUzvfIjxn4yW9y
BZJZpVB1OuXhPzXkmU2Xbl6SjkKNnlbQIYokRWpeALfNplUcuu9SC42gLlyo
w5+1wk26gkPaf1kZrlEeFaJeBMnr5pnvEolQgwWkXFN6swKqZ1qlkCv4d8/q
S+/wPpYn2b6Fhjz+Ux1XZVUCb/U4mLgDfjmq5cPh7dYarXoNnNfWzhJzj7aK
0/OPWUf17H2xWxZtaSzwL99ukd8lZ3qUaAJMscepghlkALm83F4hWEko+6I+
9IQBYM15BVw4Fkgcxir+yAcQsHuJ8EUplN8See1V7RI62kNU2X3YhOGGRFhZ
iBV3mkaRt8/SDpeCt8il6rGF2w4MnEqo/egAKRUhqHA0hi0XJxVklzovFBbb
tRMexO6yE32ecg3L7NXyGAPwxqxet/FMKVgWxGvpjk2I9qakNAo/Hw9UKI2h
qch/4RGqpbth2gergy2tBCi5Nym3ujfgi6VgnBCvGCkyk6jb9FseEu8S03D8
yY6qhCoBwBXzYWm/6396wWYk2cCmdGTvPk/FJkGk4lln9yXBAhpMBGN+j0dV
PZptxTR+P1SnYze8CRyXfHdysKajq9up1AC1+NJrDmMgbHzhpTqnYeqBt1Hh
I2rjFRcVwWJJCui+SJ+u/q9IrpqcCFSH6Oz6QGq2jKc2NvlBYk2aZyoHR3Xw
E04a43FYol5K/REkROJrQm4I8t/9znInJt/FH3L8GkNJ8UGW/COcZ5x4E5gK
dm0R8rW+x4FD3T3UZyf39hmSX7p7uBIAowJsgOIF8PThb4asq66Av0ac85hM
rfHyk0bYYIno+gc7zPTNWfyFcZaj0+5Q9TZVr3xQU45E5T0OB4fsx0WAhZRK
msz7axec0ztbm6eHw3FpWvsXfaC9g+JbS+tusFpSX5C6meijr8rulb/1W6N3
Gqk=

`pragma protect end_protected
