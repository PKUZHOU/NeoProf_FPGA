`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
N0dfsLdLjRqNBp3M0O+H+ypf5vUTswyJDhvuRgHW4gK8gXX9tIQIVNAkR2oSbiyh
R0mZ+OlL9i4mVBeQGlkFBjDWh04/rSND9YQv8ldXEjddfBuDwdYxTScjcbrjDgFl
3qPOwlMurNBEvT4aGE6JKEj0A58Vdg2oeTaejmCM9dY=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 76960), data_block
xNdkgpXDu06UWOCICN6kRd/zyUaQ9dDLA7KHOHx7B0CLYgG+lXnqG3L+jTSPZz/O
uNF7wQqL2+6Bu21cNDRWP1JFDxhZEq3bQaeSInSVjnjc/vE1RBrpeiJh2iUDRbuz
aR1qfUoGyqNcds0hW6t37roYQv+1CfpNweQQiJBdsmr/NC7uDcT8s4X1ZDdoo2bD
QkNhwYSgiPVqUHiVtuOZMUzF0JGrujKnynk+3lb0rFuPGS3UWbmq8SWUejduMRdq
wNGr0nORu/jHXXC5ZsGPP30bnF0N5L2rrBX077Rs/yysu7AxHWrN0pG5QXY56xay
8lpAxu6T+/xhl0d1hQpGfsT1W3Qv4bIUp+13SgGZiEmUlwVNk0akN3ZNL5usq7AQ
MYGZJPuUzAiIVxxvkw1gl1rMAXi51lIRmyn//JMXs4QAiC5jTAkn3PG7jWpB6b8i
Ih9tcYduNW3pv7Hq2k1jiall56uf1f3EakQTiEmyCTMoMeC2rXP0CoQu5AVrpidz
LaGcUqk7yRkBCTjfub9bBMmkMwK1BXNxK5GhLT4PWYxmkP3bMFikK9NwvOmrVNKG
WZa9XagNUMvvZ8KSqJtlLTOVNcjXOxRozpC0RottNYnJBuTbgyXKn08rWVQrgylX
1qaa+BcoNdAq9M6fD08DOPeDfnLMZvl2fOGe5I5irJmeJgR/2II/RsGNqnayo2gH
H53CKoUAWrbCBu89slT5lkozreAApuWHxosk52/EcSRU8bvc+2NrhChncTCrT1c7
bcfVt8m8ci/qVJRsi8Y/XY4eNkI5rdn9+62iZu1iEmBQH/MRXYcLzjqQ2/cY70F2
h/cxuW4UAyEEfYigcybIlyYnI6AGmoCt3fcNDM8nSexJCR6mvQa30k/bJ6K/200H
aKVs3APpp9EUNkKAnC+sbYOteXjbIPZHXkDm9ypakX+KkTedu344oXAmyCp1twv8
OZCfdt/4VZ0PldO5Pxfbl/lkTxPTeHMiqARm5r+t3hEi7wYtK5zXexmhF8UUl9S2
q7K0tXmx5C3jbsMlKiQkpzCLnYtcxrhERWcvgtRfZxpab2i6f3y1yBu2EFn3j4TS
ZV4epUGtPMHMwGr2yOHWA17P6nPx5qUM/TkJxD6ll0BCoIzlBW5P7Q7z+y8rSmPO
jW4BdtmkNNjr62PMqoaoW9yRUDung90Xit/V324Mn5fhgotFo06Okk6Q73Dx7WNJ
mdr273BFyQHUJrIe1a2SqY4qpGEuys7WE/wBdyo4U4FuyT8j6Wun1QvTR+zMjJHl
BiA7ytDqR4nF8ZjY7M0goMjVR8wo6lLhrdqsMR+hDhB6M/RRGy35lXBUNjTFJ2bM
QAe1csdG465HZUpNdcA/V7kt3zYqNZNaKuyyfXD8qIHmOeMJyHkBn3VbkSIk5+EG
/Hyw/OJfeLfJCWaBKRtzIiw/nUNYUBRFLQ+i1+4IcMSMEiO7FZT8aBwjJdmXalm0
kUcXp+tpU9AF269PsjiyxbuxwkwBjbNEVEnCty+y0Co2bsYJ2VZUILz8zsHiHuhL
Mu5DzDjCLRvmrIY1d22ZJa8KIquEbu+n9vKCN3u4qKoNdXGItjkdt8Y+c6dplIta
NzyEfw6FkpZ7MpiKEHUhaehkC9yQBka1EFdaLFEOSTXPibE2m0tXdWU441+1xc9d
kEkkUh3wB3ixru2denFZ3MtJBAxwGcyrCZ8sDDOhuaD+TGRfhsSuB9yECVTlbtLF
F0rQqdPETDSYhSD06dPEDBjHvv06Mo59N5+mfEhP81VDQ1EDrDc7EdWtMOnFcJRY
q1WhMyyF1twQsb7vWERSY89gwYj6bPF1Donle7CW6j2c50z94l9N/nLCnjee4wDw
3J6uWI21/ShzVk2xSQ4n2Fvx1KLxw/fCBPQawg0gnEXur6MjT4QdltPtFJDMFYnH
rPZFVfQdznIjtDm6DUm2Txe3dEhbyrGYe+PPlwUkhw6gvuVtYe+lUvjWsBwN/0UB
8ziizuQO2rbXuwePhp8GmpCPR5jAy0Efoatd5tH1xK9qgRbxS2WK4/gSrAFl5qmI
2AN/7xtGaMMCbUtL4IKN3w1z0FVomC2JR1FNfyhRpe9HFE6pZNyjPk+fIIE6cI7d
YQAjKSo6d3VTG3eZp80LmaXyLjXa5XNfCuFaxdzSnspcn89kuv0Ropr2z5qlHdXV
RxfWW81izsLEN1k9FovRKx66wxzCASpWcVAQnsJjgz1i8FmwsjnkZ0HMwwuhdzZ2
FiAHNhm+hlH9beV+UeYgqdE4nnjfuJMVD7KBr5FgKRCs3KBi3EbQE9EuwVsUxVEe
AE3rzy7MWhE/z58UH+cYItgE0wzPhWbVSpj+gc9HUm/9IITV8856w5fNUwicp5Uz
8bPPR9W5lA2/WWNmR6CZmS2AmAdtfWxppmtSauf/CA2XgPAVf2Qa8h9cxXEJyFIp
URGbQQU9wwxmlwsNWZZqCGwNZFvi+i+GWXpoDSzVST9qWJveyic86XwHjWRbUYou
ceqjEWEuLy+ZsaqUOHZjwHZcqlg7/rbEOE03ib/HRdxWb7xK9N97pa8A0Jnuxvg6
NLfd/UYe/Mk81HAVpZTn7VJ2OEkUs8EwfdZ6ZgfHaydUddrbmoYC9tks7d4DY7Ut
uQF5OBpsavZAO8tGM6t570o28TeEpBk/ed8hFw244wLuDeKwQoW4Bx7dJ1PHF3/A
YH7rZ9MaDTcuEvvk1TtgDifMg5FnkPt000hnijhaOZ7VC6OhZt//HmVH//LjrdSj
P+rhbSjNmy9ZTNB+oztTRSulZtkryStbKOISySK0LlNhm7Zt6CZY4T8X5zu+YFvT
jGSRcNUnJjoK/g+KnELXph4/uK57iPUcd+i8A1fBJmKMFgLL382Bxm7md2Q0hZJq
GBiTj8sZ39aDuO4Pr1AktgMAAxi5dM71XinSH1D66eK13ib+Z14buhNDf8B6MZPj
bebgipadagu+SA3R4BTMcQPDtnOdCf49v38fetMPbVXAjUX1UwVGCV69U10JrISc
3Olk2rG9Kou/8YPnNtmCbhTsOHdO5nn9Rh0nl00zLC2LUU/qfXKbC9y3gf7q4umC
IiRY28cLLDLoArMzxILoQlqwwXMZJ5haiDqFHRu9+4l54lYrR/0uPFgBk+eaFKPj
94n9r+V8I6bIlB8/CBksZnWvAlnlmA+C+HJCslaz/khZrpNVi7PlMgTr2glw2Q/7
HYJdUEDWS9woXQz1gXSvGWUuOefqGEpPLnZAJpFKpL+H8CgS0Sj/E6EWnz3HVNDp
Zft1le6JnM8/LB4W4T9OeUV5fcH+YbNBNJfau++MFU6bDJL09XmlAxwT5yHWhKk9
+Bwlu31joAdZjEIBVICUBdaytahvE1V0d8TPm1ylr1VAGj5D+jwCmcFF/9xcBH9B
gmrHaIv7BwPj4uHcj6/L5GX0AuOv3398JJbRbf8mFH086G2jgQoVahxCbZn3KeRT
1Wg9f2l7zq04GmtFTLDD023z0adlge1oYzEFcGuoBtLJTpCXfFOLJAvQKQPC/V6B
IuHCV8jrEYLDDNvm1oBeWMywreKj97ZhaAIHou1eMGJD706JdffR01U3YZWl/6JX
bLGv9h5JoWxAhb2CEORvyl+XmNYYunmiZHtBdtyVAyzOstMqMA+jBhi3dbA7+G5U
n/aGL+h2LpmLwWOxI6Cs+s1fFLYSJY3bY6/BbMPLv3cj5j/+bVABcl9M9unJSj1o
cPuB8ajFfLV700+3lKguFlNq/k+1qjDbkkTyeLwTY5v55koXEo7aIOcEDulG0+F0
ChbwXh6sUyj7ULtCcXsg23RsAQ5tu5qIeIqvOH6tZbZYvSwqd0X907Wk9PrrFC6H
mjy/iKBh/tdT3jMBhECQgarNHyxWA+vaC9BI9BV3MAcS6GDDUQduaZC4K6Gzllnq
opbQIR9uBAmIX1qpuRS4AB7ILyB4VVuAgltRDvsMN++Y8V1FwLaEqUdy0H/RHxTk
FgOjAW0mscnqrKmD8Tsr54oYh+xZOwWPU3g4LHB+qT99H3if8c+DTh1VVH1rDdk6
3lQscUC2GmD6dk8s/VKqv5/YI5zkRXmozSI/iEskbBczLpU8w7SU9/FpD1Vs1Mi+
JtfbsTus/yJ29HNwTakyfqUhIqv80bVQmj6is1llqW8Nlx4BGiFeg6XUsXZ8HD+h
hNJSeGNvUOJt7DVAJgeVcDavL79H7f3V8zZysKYWHxBXErGxFnR5hbEjzFdbZj0X
ucRnBw82uvqhqp+ef2mEHE7INKmAB5xtiiwr/3dTXQpONK4a8Q1UxCiyzOJRpz+I
MwEjb1LuiYmMdIC6kn40BFBXEDV7/i5QI0JT+3t1/FpmMPIBAjfSYjlu0wz+usf/
gMlSW7QiKgb/BXUdim/7U0QK5kcrRaT2D9hX1Ispgq0G6Lcepw9nTkwiu1PiE3Z3
eCxPwxmiYrWK8MMobR+MRqvBQqERBd3R1Q/oletyIeQrrCiv+SwcADRa7aoOEBOp
yhAUGjzAKizZhbGYG+xQ2o4iTNhRv51Ql52bgjCId+f0l6fo2Cl7E5k81wCJ7Ozc
WbxTmUk24iNmFdGiSBf7nqEh+YhPWmR3DuaLLMATgviW/yM+Phu4gKBWCXDGl7kx
635qckepjij6OUPcKRLt/+3ij9D0urqBG2HvHDdyoqs//zByibZ+Lr3mHUlbGMtj
0zXbK5MGUR/89XePKcVl0AAgZTPaayisqYEmQAI/lRCZ+opLob4jQF2GKtzi62QT
+zYUiPfbc/9LDQK1xW7w05fQ77bNhdivm13pnIKBxHmukXLbFcEuEr/w1a1pY9jm
vUcmc0CDmKS6kcJpT1ux8aGHaKkgw44uaXEXZNQPjK+hNJZyb8MYOlJ0DMtz8TkZ
nnL7x9Fsrzp2oEmy5lcLanNt0M+x5JeumWuAmz6qMQ2Pt1CotizcK1vDHsuT6fcp
h6RYYjm1D2BaSzjyGyebvrSy6ajSb3iKxwdCL0hJKlAokyVyq7epEI74xUX6wOtx
S5TTxtjOEDbpkcilcCVauNMqWKfklCfdoWl0/UEcMDqX44EDqjKsPnc3ABMVNRfH
lSHbxAzw2MlJCC9IVdKSEBwryEY2tSVD61z6Fb2EXh+q0S+jkV0z7HHyxJsm1psa
99WnMKFt2t4XXjT7x1FOoPe74fU0pPnAcAvz5dED9oDZyyFZlxkEudl73gJOF3GT
dAbuUsusulcsGKQYtSOgCkIbC0cocWhbH7jbhdf03Bq4S7vnjt43qqOyHQsRPxKI
/KdN7bMw/fgOk9x9b5mSXycy4MwCdOL8kKgpELNGNNNx+5FKZYhrk2zdA8pYJIju
YNGMRA5nycti3/JDfyc4gCUiFXUnW3fQ2obM7WCf4OunqKq6sH16RiGReWRkhN7I
w+4vAnAyX7kiohOJVKZV/Vdk5KzLSNs3Ui9GZl7yh25R6rGlL0FWcDdzJKAC8sS8
nOg5XtIZJNBq4QTjvLcdRO2Ztov4i3nbK/GAB57H4XGtf2eMVR5hPO4r6FnIN8Jt
6yFGze+Utz+NVSkJXBtdYMdnnw/tGy+F+Hc5MmN0mvCvCaM2be08KwUkJ/NQVHPz
f0hqNIGS5Pmi3qhQdbZtE7sX2YUuW0u2+e78NYJ4pHgBKsW+TiHtlmIncAUBtqZv
WxxDdyolgQdnvuaRLc4lYgaUUnA7ZGi/rzBSalObwc2lkdT4trsg1aUjUivtIHal
3fqA+WTFlTSNBSdH/RUh3pmezmJ6OjAp3J3+loEHlY+L9PPj5hUc0tyHJiQBFPbF
tqyZMQt9DQp7rpHrx9MkwsegcrzblSiiBMGg03r4BGULCG5iYvOYC04CQoXpgrYk
nVvOiAXQP2G5q8gerh1SXX+6hb8fpLAjrh85aSVBAbfKALmJPRwRXbk2lad8PbKD
Eo+gU7aPlqxhudKoDIpVXFtYxqjnjEUg4bxtMpkR7MXoWsEg6SYaBuzb5okJEbxA
RTNNyFWYjWdKlTXHH4eYKJo2chjP0pB2azvL+45D+VFMuA+/gaxjiReHHCQFv+tz
uucW4kFPtQM0kWa0bj4b5D4sKVlovbPMsgGMLsAkygesnS+WS8jkeXqHmM2kpkzx
oFqK8mmZ7pcMojBTcCVYstyfu5v3b87j5oUU8Ld2QnhGZRjebGC4SU/1fPfsXsEN
W2yIwZ20DoRrWqihVD1CzH0+LDl2gXzRwxlo7zxu1tkVEQsEanXe2T+I45wo7xDW
P7hFRrLkA0UG6WbVsdqNqrVBGaa4yQ9jthf7wJWiBeIrqsGnxK2/ZSllT1aQTgWE
5leTZl787amyyol2mv4KJWiOYPxRHZSTjeKjG+Q/bIZ9d7MT/gD4B9Gpfo8D/1+X
NM41foLsl45qoipE3ixh1Wu9FaYYchb30mPXmJHYmqatwErP/YTjHy/uH4ekux9b
KDByh+DaldO9r9IDcHEnJPOaDw0gIcpxKZaKYBNX68QuNAWIhX9Z1ubj8c7GU1wl
b9XcE/gwMDqpap2ojcKERYx0r/w1Dv5zpsQ5rEDv0Td8Mv/qJXFO8ejXfjqGD5X1
w0+c28VnN7sOQ2FaQAkdpP42zNkhfKhJwvg/wMtsuEkFFwbKfqtCu7bw/78m1nB2
sdohobkxP+fTrNWOF1u6triHbnhaNEWFbjitQ+BZuUNfhzr2ZcFdVWg0lrg8/vUM
G6O+ntix0/Wnc9TGHi84baiauBmWoV7xISS7GhuIk25Ier+gQoSrzQhTShIGP7Jn
Z84GSQjbXORh/0S9C9k4HxiWoIFU5jeDVgohkPTrEh6MNTU3rGZLFvjLoWCmMjDT
UxHp+/gb03XtDOtcnQWz8CFcDgLBMN7CYFc+3OGForu9wGB84+kFS/41BEhtijy3
KhahHWBgM8dgfuZw5NGS9QJOvWyZNtSdusFVbPDusMIPM1J9ztFzlr0ff0mwAiuZ
Y/XSUX1C8veCTOpp7ZaNeVaLmJnVtHu2NT9qt59x4xW6cldoTWcGWHm/Rp0TCfom
gTDd3zgJ02WF1Wx5g3yeMdHbp+Ckr/0pkB2v/LJ5btQBKU8P+UDyf6WReRlV3AU3
g1E5In7IrIrmLCbcGSb0NRCbe3aWLk5yKVbNZZtc7jnl/2XnC6qHlLogxalpow1b
2CHIyPZlI9mbb+mbtXxc+z6NuztvQBMU7y1i4LmzyHQNHokBwdjm6EXgYsGXgwfE
hDDdWD9USOFkRvbJmg6rrJV92hk0oYCu6C7ImmiSRrnEQV4RJd4E+q7Gs3A2u2G2
6HwI0xcK7Z/XJPxUAJGHqXFfVGu7GTKHXJDKlsvHgZextDty4TsLgKRHajDLgEn4
h/SZNVpoL6KWeu9S9XWtx8vktbVZ4pXBPalrA3YT58cqZMxT0JPxGx10TWtsoi4P
R9hv3jk8X3oQmrz/DilYYU4F0TWjjrSiugpaaSEp0KWk/2mCC+nY2IvxwVWEhIHu
FnPx2wN4OCgvb1IXxS743lffVgnSDNXKEm3DKmvPRY0APB+hnWjRD3jHPLNEwEOL
ukLnraxJKcNyTbEIExrMAw3PBh4ZXzARmFxfafokUkpt1YXUpwfe+zp3A/g+SrzP
lxl7NGiqYQJ53A44usn77QDR11VhOJXu5QMNLjIUqg0boet+aw2Cb9Ik62og+QJd
Ud0FliY5mq5Ee/eOgVMov3uZjij6rZDYaO8s49KrHYJ0d5b13zASflk78vjM4o6T
NYsZPhOcDKrEWgtLMs2VctDIR+4tiyyIIWdkINAzQheurDyZlRzk7V/Ktqdct2a9
6wWzA+Ne3hnfDMcVVshjs75QhuGJiVL6YoaJXjZufNVXlDiyx38Wt7jxPzxynWAs
n1DjHUw9g+GVR5VmIYf/EMV8fBHCLiFi7/tcKXYPHy3vYWlFxwV4F2lVfhFZ/cNJ
Z2BpdTqZZ/jPMjYczZBNC8CnCqd7k32L+HqwrZufucPVuBuo1jF0LTUfW0lt+hls
bg0J1pln4rHHh/1Xw5ZbtQmkG/ExPLCEu4Gng54p/vveLLmkD2/eJ2vM6GU7isTp
CCldtSCtnF//+hDJ2yHG51vnYFWPjX3NSZp3aXYw02X7mu1Ld4Ogp7M1/as/Dj7R
R3oVsLuUBl7QJ3FpBCc/ny2Bz2mf5W4F4WKdFx5+ZU9EioRaoynGCgx8gw2hdQMG
lEkOG4pnMUUQ7T0W5o5ujziLAegIrHFjKHszR6rOhRI1Kn7dJIePTiTBi+Ch9HOf
uwbyZevUZ+JHeKoRKNjApLZTY+h+ppUX/u9kfwxsFL/sqpkKlQ1QjbwcOgdwbtfL
K8M+MIl8j00754Tn2Zjw73jg7ZbRLfhPCEP2RiFELIIQxz6np+SXjY3Mb6NULqma
ywS98xNYTtBhtg29fkgFhblQ0wkJ5LHV2SM1uRBplUZX/u+qBCXATndc/ioqrHox
udtN7tFurpQgr5SjlbHcw1+zYeuKrc72g4caiTZB4sUCkJMY6kpXC7uxvLDaHoXY
pRQMYvTlfLxlWb9jI+qpt4BqRU/mNKzA4Kit6khH/wFhHD0dJoVU5jRbiiwN0UvN
H0xmnVamPCBVG9ba+m3gEDwyFymgsLuaXIr5FcpcCzylSvMAQa4hNBkKa+KxOaZa
MDvY+ITGhruWfLuLVsBNhDfrTO199Na6DS8bd8MmZVOv715T0oA5C7DbRSri+fQz
Hkx4kiU41VqQ/5KKokI2rB+38hOX9/hOfNadu9u7NOQ+x8fBwoB11Xztpam3MNVp
2ARUW2FKKu1xwates31Vdd5pYP6tB42DuUvegg+rUHCMVnKxof0dxF0fQFmaVNF5
VyKaKosbzr+8UpxbQ94ExmnluxddweH9sdnTB5nU5BAwpaNLEgUhF9oB7kmmyXDx
DXIyZi18s8mmeKOBdSycLMm28s2sBd610iLVAt3tb1jD5jr3NYyVAQAukLDw6epZ
oK+PG7uY4GW9PoEBKce3VSJPkiWsalR3CdPh26kOOFOI7Vzm/B+pvTeuhOJ8LXoK
RrpOZ8qIgIB9WJlxwBqPDGuKtcF988ypI6tvTjr/t9nYdL5e33Lv45KLtP8ZLV74
RXc5xezYVc7Y1IKqxEKoS/n8CJ0PgQ9UauwYo0RH05u0DnAragSeDyEQGPniCgbn
O/iIRBred1TKkwX4cgk+5cRuDBhYx/apLMaXqJFptNLwIPI2XkVhFRXTQIvZs/ny
eLh7M8Au7LxxTNOIQWcylKK/g3Kogi6VUzcmJgK/i5kh2yF9cFSspdNJv1fg5l5E
rz0p/1t/pTnhhqV29WnykXVuyTD/+ybwjrZV10wx/KYQ04eK3En8ujUJh78o1qRs
Yzh/SjSVD6NmSzkkmans34X3uNiQnMlZHObT489LpOtX49khfoFQ6RTZ06ztHSPT
AZ56lQsK3TPKhHjccbjEc1Sm2Iv2tICzhrBe3/M3MpfL4SXFQxqHDa9rHxup74YI
Xbjb/MgnjzrxyxRAoDY4kj2So/Jqh1egcsrFAa0D5xGJQzH39viYntyxumLRioZR
bvt7j/7U0jUP0bq2SyfIRhio+I55YoNV4vztpV15BLy3xj4upr5NUxb3VXehP3ec
7UAmRqdjF3tPScq8Jmkuxn6oLEzkNF4rEYYMht0UKTG5Q9if2Vpbe8Y3pikyLf4m
sNmJTABzBEKq36ijAIcbjM/T8/wVIvfqzppesQupZDohR8Crf8l2gW7oO3tiPczA
6FZt9HWiqRNPWEb1JPXJR9DH6ovv+2A4OzUr5YlhgydQXVYYhPQA/zexuNgVodnw
Q2VquuQGXh+lG/3jN88lmUn2dneEsNQyq0rtL6oX/ypz9TUFy0qRsnfR889AHC4o
xoKcS9CgOSGaCIc0STAjxmb/viwys3wTPTByw1bBOnrVF7RuYRfO0qkJsGmJWI8U
bjlcHsAnropSUWMSvfyGGUMmEp6XGlr2FzpKIS4/1PZbnB6A1ZwB79MdDiEZFvjC
d+cUWLGefRHENzZfAjYFC8xtKYVfFdzXx3XJgJqhdEpc2tGvx4zyCw3KreUXtDtN
cjCWot9EWX2Y/KsbTTD8d3/UnJDtDjVO8t7FB0TzVKlPFFuGb9Vrw7/BAeK0xRAj
7p25xtGIvkUeOH3YH/jboR1nSS0wgz9yzCpClTnO5/PkfvmYxJrrSBbA3S/trWci
yyIE8VRCxnbnsomyffZjKNf810NqRL1WYYnnvwDpGvqrpRaG7SijSisQH57s+8Yw
ue9x5ukC3ODwfTQSGGqy+dLbj+ZrOGNngaTMw4zmkGAlyf+vkecS4MWlAXoKTRVj
RCNT/VLSZ5YSsDNeDzgiWJP3sJym11tVXSKB2cpBsuM3xUZBwrgT22p32vPpcAwt
6iDOeapkdmZv6ilu9ZnjBHAm+K3FtHKQNbNzqL6n76ghoJj+KDLTk7UcaToFmjGX
cQ4t1mgMG+5Z5cAYAZOmUgqty2e1SP9NFPiHSdBM8uUD9zeX7CuSzQB5/2njiIt/
cVHI4t6uK1mwPOpw1IChDmEy0ahxL3EPgsVh/QR1xvwCkJyjprEa9NXkzwZSNLY1
VBHV1VVnj1wJwUSPruGSjp8AOTY3KUdk0u72pptNbyUeuUiAsCOsmoswBJS2wcXg
uat+e0S/Euly8uUke9OFAVOr+WZsGD2YZ3EK3VhLjaOauy5oZmBmKYmBVjByqLrW
cQc359FBOvYtIqqFswtK6Pe/azK853Odm9zk3K8rmzc3T7y/dapUdaev1gV27gar
xqL11EL44VBe/LY1iFZHcX3jRRmX2LIVioYhaUP12Luq1n6PNX6vLUpyyjzQdG91
RlzL2OANkLIxmyOf2XsHRp0Eo+i9Md7+PU83sThm+mq8B6lUryBC6tdbtjJPI52x
SLzNSMlbKqsm2xkIIbQn3tjAJJtJrlaeEQIAm0bm/jDXaOOLVH2d3IlNctoE9PCq
lh94cVsP5Phb17sOJE9DVmhT+fJgZiljanB2mT1FYaHA3RPvMhHVUXoITIv8jf2Y
1fBmhOCrnyPlH5ug/yc21kzOLufYS/9f1wb/V//ar2YvjQ5UiVlhE0ZL0kVsc95t
PjAvyV/aUKkJ20mf7LGm5lqnb0HinjZdQJu5Sl1/k7wQk44MxxUyOCmLxO5RUT6d
S3IOr6ookNu65wQN0J7pTJTkdP35PPT1chjgRJfJk/IiXIn87RNw50vzNScvyMiH
/iz7Wrl4lJZp5/5atbwsPWAd+n7WUccEQeJc1CdVEMlWrHIZIIvd55/ql1dT2ncT
BJ7DnmXuTzGjKlBEimcc7MjYYdq/dN/qyFyUTNJ+U+QpoxrjOMpPLvKpZz4W5zzC
hJ2ZYsLOz5frGZM5yCB47elew6IHeHuWWDKF+DCAFVuEpfXA6b8NU2dnKD3hJTFg
GTegqCwUnTPp7K8+lzxiH4vG70ki/344nU4KZK96ca2oWkckCsW7Jmp40m9OrnW/
7i/TyyBUf4C6tJKpgSTVxZBiqR8H6hww9/bs9KzUM5bTJ6z3w9w4EnaGBXBVO3Z+
DBd2MSeimbIO+hskwP48RCOX/6i268KzpuW9T6167cAvvxpqSWy42+AWw7B4gmwU
9Tpl06cLkecS3s3o/n/d3vm21Vzoe826uFwEQGrP4CYwEiiXiQI5TOXue/AVxcIB
TnpVu5Z2S6M0/mU1bs+C5H9Cy7wsuPemZjXGHrqIXS7qcpSFOBWVDvfw4urnSSXt
NXvtaMgYe94+XvBrFlyGv2//v7R9gX/RWG4dl/qejCp0iE/tjdqpfxU6HPraiA+x
QMhzsadNCPLmIk+8xR0Ij6i3VPU5d1mbxKC9Pnq9WtguDRlpdWCb/0XsX5NpgMc9
mbH8YW8ucMcjeUUy1bcg0xABxmXG6Z2eqbiUhzoORhBIcF9gFPzc0KzGaf54q9FU
gRDFPU7yjEPcuwrUsVqyQYFBbvN1t03l7ypRuCBY2ktPUUpKELl8nQ5juPWjorpy
C4X6Jni3lMjpMQxVIp+F6XaHj94ALvG/8LJi6S0uzaSq98t5J1k6aHlOInVZ9LvB
8a8qXVJtFDNJbngrX/Yv8LH50oAQKvHQPi7cwQjAuSNhvhMlW2etaGwid5A8LsJw
z+QUDU4afFHhru6TXv8/LoEx3rc2klhn/1oZaQs4pEW+eE3zpSK6vIMauTPVPFSc
c0eTAe219kk3RDHVbswJuYN9WB9cdjZnaVt/5nMZc9M6OHYdRt2WPesfR3+nO7Hj
NcRT+qrHG+z6waa/1YZPRW29joIjPAxA/pkJHb+Ylk78bTyeHtC8KucfzmITpXOp
ZQyx2GoKZ/qrThdY6gcU66zX6PLkJiQZsFB6qdabHRHj9d+eD04gqKVm6kgZ85NI
HDcgbw4uC2bFP70PjEeLBsyulT+owPwHUO/jjZkeWmzVPtfBvRDeCdq+KvrLZz8Z
IgxTiIsF96SJzDpkrongaFCTyTi6CnlF8lj92r7+tp0FsZsv7JfO088lyJrIslsN
zCyMrn7Si27NoNTf7IRtoONtJTEuZ65cRX7d2K8xGJu8vA6XvgsI2gi1ULlF994Z
cDIvFdFtlOKj00evdXYVvFBjp/E2ih1GXsJ1JWDS+fA0CxdhXbMO72cKKXLg8S6K
Bcn31Ap/yC5+/9bF/1x3rKpHLmHvWDpBHjBBaPSwv3LMunBqtrW529KLnA9HPvTv
qMuO1pktuNGtSjDSRwCepM48DiaDm2jKUVRfBmosI2VSp1uNdIO/5gUH1gCCG52h
/orlRW7W2S0I44toBxxKdwTMNwvpqoGErlgwd7JbW6sBC/QmeFfkFDbQwVilaZ7/
p0m/G0KUnp2nFFomd78FV4ssTGp8x5KB2l52uEi0aEP3k9yiqT8pD+giDZQYx+9c
5UB3APUKa4OmQ1cITqZtFCo/XxBDF1bedIf6VL1HDofpufREJ5Wi6C2IlVD/Ci2V
yvT6s2Kqsxqs/VLX7OUdubgdwMcVDnrevP3dGb9eJh41xKIh3T5UmcZctmUxP3Ro
Kz8kGUSBJTJo6CUb2SBLpVud4YroOsIMuPC9FaA0Z5c83E2OoHq+TTH48PUnyb3Q
73Lm6rlC7CqPcH8cIo818iNThQHvdLlsqQ+f3CWKSG/8f+F4UDWOEF2lws2gby5E
SEZ7pIhQoowogyuCTZO9LR/78+Ke1iOGcprMAADIq9M4qY4IjKUMO84R2oA1IdoX
YMhOzMvz4Rd+IEBK/8PeuOJQRLvj+1jfSHvWIYsXIV4EfImMOgIKOnCr7LJrSql1
PP6A6GmrmE9aoQ9+9tGJ151nbqS+QUhnHuELyY2m8u37FttI8R4p1Q7NmETMfH0F
oLbB08o5p6ijfhb6qIM43rDcdW8Wuqza/Si7lXrmbWzKaUqa5nD2Mf08RKPlrLR6
Zod1fYxjzftEXF1KxNn2RXNwtJ3HVcisyAC81OIqcvVL50j/4QYrbcBm5yWq3dqF
KjA8ZIe4TcUIcPGHhAjQxv+lG9fBHDOsfI3eSxLC9gvMMDis/AIfKcD9IzuRxxSp
r9i3RbNCUyWBaa0krNnVFgPFlFTvMFcgC1BpTQva86y/urINOynMAHQkTstdxykc
BX+7yj7iTCnUYs9PiihyXatJQNm8SV2v0/8fNDvakSVv0CviVQgbtH6TtFllzogK
d6y7+fgWLH6MLdcd6KW0ctbyljYMvsLQKo0W7HKkAXKQkLcKLUuJUoye/KYLgTcS
kL3uH+u/rfItYbsSn7GhNuCd+NLrb988Ld4H9JSZBvLTcaWHx55CiYNg6B/ThRXC
cREBKhdznGHFYDcENFT2P8blF0vi0/RF8WaFYkPnHGGals+ZwvMpFi3VDVq0Zscd
eRHlVhFCDAALBvWDVXPcIxL7Dc2xP8svBIDEGmgUCPUI1wIlo/ca9hM2H+L96bbO
TzHah1DzhXgdFjq4v30oqdHfGEgNy2qZERiGSceKkmjrKnG7vfOMrgGCFHgRzmPA
O6YvM+qexWLh/sD5JTtT7cNqtfYf3e3AOWHU1oYk0iKURjRBD7iaQTDyN7faYOPT
bhLfJuKwnGOTUx6cGMjM4IRkKiEPNEHPcoaGhWOb0c0slo5PD/xyd63fJ2RKtV1g
cXu8quKybjb0Y6zvJw3wKr/i3ExUqDuTv2+rCRuQdNiBEFflnBRnpBoslwEPsLVf
9TYXHP9tpbD9hkgEMrt8+He4cmyUzM3PCgPcp3NI58f2XUe4gxIrTIhmSywJM+uk
69CbkTha2HqZU+mYYqkpatxp05Sxl07Xxir0GKpcs6f8kSPD5KQevff45sXuSiyi
k/9qLQUBzcDyIsKcVJ093j5Wj7LR+Lnhj/lRcpb2uOfa3eOAooz/9A3a9sYBqyWb
Y+2sTdsU0HPRAOEIDELLMUDin0/16yflasxYgmpvrDUdZfhR9+dT/bp6lNGTttMg
yc9XXPy6G9uEKWvoeCtwa4c2uBmN4QN4YZszPUVp5VDpYC5pMO4zGIwWUMGO+14x
52paPaDsW1taO8Cw4orhRsDSh3+Na9ZVebaf9XqdnQchY5Mro7NAWrL20DcWqEJk
PBsLXzXIlAyHJ1E6aMLYX4UZuYr9OxcZbJOFOeCRvb14HzyIM1RKn8w7kGoRIqVW
XjcLtsfCIwIgl4yNCxSmOup3nTgodrcLa9OaD0oQF//6IGDslI3CmJvroBGSWJca
OxjxR87ZAhhwxhGO/S5Yu9mCW4K6zHJKWjRo1n9tmF51kJKsZWx0kmvXwby8vAsU
hFfXZDQoW/OAGt4q9e6EsbeAPDEfDy2l/53XImYqflDcrak20Ru2j0v9SkLeyHf5
M72GairoWddXpEYdL7cfo8dlbp3Mxc9EXDta6AqfJEFWvCFtgAcwyZNovXPpMq0G
lkmTfMksXXPgW+iLJPoSRt8vTT7Fmxko1Mm4PB9AMvm2fqY3FwO2BJ2lf0s4CJnJ
E3BS9usVJkBNvrw6P48oDK3potfedLsHyjBxMTWPpWVUo7MjxI99DktBsS/+PA4d
CbuhxzJJoAP0oWQZ3c2oYWSImAjdP6wL4UUoS4CbbAbymm150aga6qXz9kd0H/h7
zkGIFJB+EZiFbQ1OCZb3KpaThNzz/4scBQ9FzQGbmlqF/4AZOv0tjFLGcVYzxmKk
MbGThl0lIcyLNjNfZhomfTFCzmg1BBoeC8jEvL3xkdnEfCPTeE9yKS7rRpA1SkKk
ONbmqKEdkB0VN1X1LexU8wkZuhkM2t6cn01bsH05C7fiYjG0lTAnFTn5CWLVrrqI
wBMwA+O7QKQnyAixCM+sL5gmEg4EkUFtDOmtM1B5RZEi6/r028TaaNLrlYOawRgo
qj08iWZEIUSjwqrBLOZNHAtZ+u63O9l05cDQz9ixNZ+LRbnQLCifHaYkMi6FLvC6
SV/E2qOxoONsrclz/5rzv7PMiG/OgePQkXu1uCkwSlySIgSuY+4h1t+UknpcFTVT
k00fBQvbDyTCzho1mO9zsGwzqNk/TftoOJFLhsRmxpx6uI4joxmHxta3N7XADVY6
J0LckJtfqgWw/RaIq8BlTzmxVFlLTX67Qeb+LV7phanYxLAawdBwFLx5Tgh2CXEb
3/SdlCs5xVxhJcn31/PFkM6HPNp2u3L/Qo/keeoJ+w/g2YQ/Q9mcOuRjo7I2GjOS
o0u6JPGpwRE+vbn7otJKhvt5bF1mXDPTCQOeP2ErsE7mt10LfXZecR6BWEtiTiKs
vBIRXZzBMPe4rrrW3Y4YMuJIWMAvdZkqDGqcpqsXEvzrt+QMnqE/C7g70/Afb2PC
5dfGqVV251dAZOnpWBNl+q0TXgH5nuk7g3gk7olVsjttbl7qCBPK8X4/sXmFI/YP
dflR4foTRiWlUkD1Np1MP2ldmFmgbOpISKezZqF0hdfkO9iX65O3EizSG7MTfJCm
NyW5VcUZrVnM8/1y5o8F5GbBGnVWEz7uIDcHw+jjaO4gYjPsCR5WD10sEQWxDLPC
5A/r5v+MEs6PlvVY6Mkl+g/11wl/F4N3XxqOG1XS8VbU6qZptqZM7v6NdIR/sw9s
lbWxca8Em/TCkHovknmscV2uLTsx3DroVP1a4k439YGHaQYzDUNEFj8bc/efR0oJ
FR7V7ZYnbvEQjNr4p7C/oAoybBc0a7Ao6FqnMZxscyMYaBIyL16VF1n4AXYBDXNL
3Owl0NnP5lM6SwGQ6L/eF7lSxDQjJdD6oNFs9uK0K8KCYhNLAt/I54Nocz+Wkm/W
2JIDx49vpqXmBCO/ZSk2UN3uWImEtJz1BQzolJHeQeicr2Bi88QJtzSOIZ3mb/W4
Fts4Th/GI+d41n+nxzHI4B1+dh93ooPol8KkYRMalu7E78aceiawdA1Zuwjz8Jex
b5+nwDwC0Z0bs5T7M58eozvoO7b66O5eLRUoDa8RCv0DLanrkOXwlE1YJGzgMOaM
vW9th0f3Cx/rw1wqenf9rQu3ACvsm2Kv1BIghPWiv61Hl4IS/FAaQO5YHWT/dMt/
iJC4uPSyAq8xsAhpXW11n1z5PoD0NRLETUWBk/yk+G1PKuPkQtm/86aFnHe+X2t/
uwxxsZ+IsF3XeYEGyXhXVDW0hiek7f6af/vkc1QPklzZ6UOXbfRp2y4ZDZFIcCB7
2noT9te0U/Va6Ns86ZZq7VCeHF7P0azsLP4WO345goLBM+kQGHTscP/0uiDXlF6k
HxPq/jenYxmKrdVRmkLDHradWIJ/Btx10I8Xt7ziLscvqRsoT0iumLHlduchjQ9b
OHxqq0UjqI6xba1r1+Nu6UZmJRE5MSEcnp90yDZI7lW1rHTl0XWwk68nvidgErOi
km8olvO/iP7JPQu+8IsQEfjHGV08DKOD5kRNTf6QnTl6p7ra4dujx8BPGBJ/yGr9
KELAlTwYvEINFLLbV11ATjPueSGDJdBibciKx7FV+7hGxlhqzx9ZDPomUzgT2ROQ
eO7IoumqAj3Tn4ldAfqJnXffu6b4b2OnjZHe6nfDcU0ciBxdNm/4UizIowtKJPgj
hZVcqCzF2b+sgxRKIvD8Go8VxIcmHwMHoNJYosSdaPq8X+KWDMak87WbM51QWc1N
AgsHM1I+v0cNT0+D8XyRhs7I6qjG0aDfdAB4MMVSVmgY8C2EnfG/l7+DCDpchlZS
Z+jYw/dH5UTnOUY/vrMUOdvFB31WFadSsRGJ3ALs9jHnbp55MI3zKrwSAETIOTln
nVbHd194YqBcKH7PAsZ0OO0XmOfOxlu8L8i7+3Ffci4G+gKzYUcOCrCEHNpMCNqm
rrc3/pry63UqppLwQ+ucaAcPViTfnZHOH2bZk/G3Cnp7d1u0eYcIZ80knbPULmlD
hriEm9jcgfCgQ8jkUGO/P1OzbKPb7gdt1jY+qRfjMkanWcHttn42VrPGGrEEeNwz
InzX9Rts5mrpkChnvIISLGpmNaifdIoVX7I+aMLHAk1SXPduwWAcG4so14agcwoS
LDWInevHcEFU8c6NZgrfBBEoxAIEb20gKnOYSAF6en7hm85N127d0xCGTkoXu+1f
elEpiJpnAOh748Bd9ip7aSH9NjyTWYvfKvi5BuFm9BEywuUHe2a4VcwqgazmVoRe
RTM1OlXyepdFD1b6ecePcmt1K4JcmQqjUfkGL2xznIimOhd0XgTpeuKW6e86F56i
Kc9gP9IayTeDkZsfLOVDX7RbWaqlO+TZf+ecHx7VYwlAr+ntwXsZzpgHGuRQ3wHE
jQfiAdHklbbFT9cIo6Ni0ZVwvhQl8LN6Rh7JieYHJ1gPxXMedg4IX6t30B3Bnr3a
fTDWmNpoXuvKcYvXVe+xeT60S72BuELd1IX8rXPyD0duN0OUfnu23hYv5uqfoBtx
soknGXqGnpQ+C8MFTcUG8AsTeyP4oTrWMqzbBWbA26EXQHJn3O7SDTR0cnwdNcoc
3ZZ6UEMzbHS/b1p7ucgTElniK2eBNhmhnZE/XdKwcedW3xywChRpcL841vZlHdPN
sDQ8sdmf0wOJw7/WTHOKzwlGiwBtEbg1XUYpKsj2zBCGxxYvS2tnvxldPqWbJJgU
SwdZmeBjDLtCuu5s0NL98V7rwuj0lexVPBTkGNZbSNk+RCu9fp5whVae/eQ/pioA
Hi6SV+W39il38IpyC/Fb/Fdw2wOS+Ub0UPtufgG/pUtCu6TVidy9dUwIwezKtbZ7
GtSr7KOouiUMgZfi/5GO7yEXmMK311gsvAE5jWscTsXGo/Rx37WPyqiV6VKnCsgz
nrSruSVZrhtbYb9mFoziz2Ku2qioPsm2EA84SNwZ6NPmKbvNQohiPNWz1UkJbJq8
ud+14/dyf+97vp+xlUo65mTJQicDsfBRVXJXUtSG73sp4hfhHdKvYxAECM70p1Ik
vDgBobu7n9ccf2lxtDWEAIhSKDj7dwG251yxUKn7jCL0SyzaJEtUR1PnsnfApk6m
oHXFQScpPAQs82l3l3hUkIrhG1DJw3N1s6jwyTPKg2Pmn19yv+xX6Vv7f2GE13ZX
vulP8YsISf7rv27sERFchAEyx+ULZrfONZpUvrE/xkFbW1+DMN0NPn2s080cFvTf
al9jmYiK4jCpyRIdkiGiByJj5BKDcKlMTb+2xIQ1C14p59sduDZeBNZa0JGfCO+f
qztyBbSAKE5i/Tmd9QFlfvnV3cPiKYs8+84yHicPN9+G5gMse3/aD4tEpT2XvcGZ
91HxTxazIxtTBi4w0kBfF33J/0COtYyasAMt5IFNOdK/DLFSTxkHzov3jzNNHbtU
6dyUBXkESRuqr1mv/H7mF/ISDDjzZQSiMjyCkLtBvpojlotoORJWdPBEumd7M1Jm
1nYkE4ROAdfE27DaPCNkliB2H4DMytQNW0W27cZtCZeWhXQCi52nmt5Cfhg98wU3
L5IBAB2PVodgR7wK46DbZGixghjHbgXLxvJ7Zps6RBPcLCuqud/abBnEADxABadj
BLQmU8uxbV6RjnZpWB55UKlQG6umckvFTVyFzJgdRU/+TrJ/tpXI5x702DwzNyxa
CQyES/K1n4pY4T98dfs9gxdVt6TeZ4ECV/LVwHjppN30KOIV/H2YZBWFjz728iw+
sP/OH5aRGOPgfzLDMGIizYlZyyj843qkEuHOfg/XLcK9RayqXpcd+KKxy28zFwqb
pANnoIZ/UsWu0+d5H+JEk9aFPiSMQia2O4iU1QpkIC0x57GmP0sEVqZOU7kt6CLb
k8sgggXu/slESeoGPveigOYy6ukob28OJh7LMrspJ4Zxo0rWPH/WcwxQE2DEKXZ/
rzt+WIL7B1FvR7Cl1XqqYw78S9pqDL3p2uBRYOahkSMXrf46In6OkX7cJ/NmTk89
yx/W/fYVTblwUnIQq+AtBxtd6veox/cj0pLQERPmdhnrGJUiUJa8ezDRbxvYEQ5Z
7YM1h0dn84RCt+Nk58qALIZn4jWhD8LvpnUVqxlnpNfk1Aw+E4PDWVC6K9NG3rLn
DsNyPyNO16ConpO7fNOUDwANznh213ND0Sp3kTEdpWgthXhTVcis04h2V9C+/bVN
xrD+CW3hiCOXQda7phfJ4IwBJIxGTgfGVYIXQPBGwm+mEul7zoIJmr4Sv1jxmSAx
IptcjCAsx3Ds5MWDz3IRnooc5n5lBikS3CmvDiu1/HydZFLyemBaqkjJ+rea8o4Y
uLd/CKatGIMWXuN9fXyj1JHPDszkaRTkS/wk+6B+JokO5+rVkC8tQvzbvZDCApfN
9ZNav7ryRtSmYcjdDsx1864PzWE9uQ8y+Chgo2Qo5XRLG6mv15AnOd+6zNbywaYw
AUPfCuZTotzZapFjQdct822BKxKZUWleVwCfkJRHGr2NvBHi16ikPA5fcd04DK3G
SLJkwhIelfDziov3K+wbRcWqveaJBRsQc6KuLs/N0zVSIWLf4i+Wgd5rccJxv/DO
+pCvqVrdFfPUW0DKp8M7O8V7lXXo+t1/xoWaju6vMh+TjdvEo5Miqs4KtAYV3z6o
o0z6O17gX7VLunykH+PdF2MeK0WxTziRNpB5vFyTPsK5e4PACBDQ9HIA6BYIfOSt
N34SghRzUcI+22TAQrXWfMO2FxdcspVOM7yTonnlZiWniwCxBmQIzar/QVYLMwmr
vcd8fmjW9MxevmzzOcxV5rfhFakDx8piMMRow0iBdMGPL6zLrE/jlfs5dZDjRbna
DGakC19T1LJWIcUa9HqrHyICsGUYu4IAPnCA4D0VP1dsLeeGK51GUVimS36i7jOs
hzJmEFXa3cw+trM/ztkqyOKbzCrT+oLjEMHwD6G+/ZQxKu69GojCQY28pgaSnVNq
tV+HfetsM7msk7BgV0ZnezDhpg4nGUdtyOPhd+xJCKx5SU+q4TApe9sH1bvrTQR+
mYdckeDxSeyvVD5EnthcXzKBAsuvw1PLEcFfF4aEpRKUN7CP1TH2zK/Q0UDVmXgK
ozRHkGCDxdYlodOQTIdHfZG+ceLqAXsDXvmj317uiPQJzYA0j0VAAU21B7TkTZyB
t9rbXLkZYJO0OYyzfDRBjQH2b59RnMsuPcNy7fuFqaHUyiDqfWUd1C9YeOR0rOhB
p6oy+7n9RYFe2/MHq/jthXkiPKWXPe3rckv4pD1R/7RMEz/MwsfCgU3e/2DQOWbH
OhKWFjuIB+jWT75sBP0JVLPspVBw91RIamDPsqiwmk+sdhOjOq5DcpXx3q3CtAkQ
FlfvlmixbEeinKnV7tsUNTvJ6W8ZT33Pk8q0BOixVFaUle+30iujvkQi8wzVFnYK
+VwZT5q9T7zFia65y9jkSycbLbWzCP8lFeVdBKO2G9PUZRnFstxTTELNyvZagwdi
cTNPNjP6ASgPUVZ4Ebv9Ua8pSQW0YXjCl7Gyaj/KxSqjvWqE5BfhUUroC9abErnu
Rnk5C8a7A2BLNOGHMYyQEVMfKZSfLQ+tkTKuawfTP/8bkHKMXKAqLBv2epKFzW+I
ojnwBIlfGbS4v4EKQyUJlwCLwSKcoJAPKT4JJmmmqPx2VcDx1hLjKJZF4815IA/V
BfFSC5kQ8zM56bkdYLaZ/uqkivut3BgyZjD+hXqN6uXwKhbMLyvFjjM1JkYcpLCS
JpRmaJK8nxijnf2MSwQeQ8IqyzUdAoxMRsmgYdEzNQeAmKLZUnGhBI4tix+QArI3
wZYoHw5UDY8Kzg2O0C12aYTfXIM6xuiTnsutRWrvGluLb+dPxJ/UDHBzgXi1rEag
Hmq0o2A3kav+ebWq6VYzcD5AnWeygbXe4s7zatZqwIQgVWvCLMnp4OJhQ1OD/mTY
CP6Xux936ZyYOs1DtuFWA8dITAh3ZfdsvmAvb0ii6wkbIsfHtHa0Y/qWe3geNB7R
X+ReRzusbDsxzqoO4P7AWkLd5xmhlCnQguEwwbNKS63TDQC5uQWlMgGg7cNLdqQn
AxofDfWekb5nojZM4Umci6RBP3SGVZEAHylFTzd63hx/NNATfbFBLaYn52wHxpWe
9NkAGTnHRsgb0A3426TFOJmJs8X0iNplSU2p38QHNWJNdunmhp7ExV5PHuQjrnOP
2bFSGWylmJLeDii/0tUQRXyXH7aZNUv2R0h1nYYM/nWDCj4M0YQpaurLFBVW2Hj9
t5b/jCLxKLWOs2h6X40m1RMwjdjiWA+0uMDohCr8zivKd9ApsVZOx4FcVulcazMv
ICQNlfVThN3EORQ97dyrFiLCfilsLQP3yzAxv3efCO/OjSvsKDa0MFV+8qS9NNyC
Po7NIZktSIQhlLe/Yan6DeiRn4R/hXIxpgeHtZyHSDooI6Yf9kaNK2f+PwsDONq2
r74IaPPkiHGmn2XSFYDXPdXpHos6PhCTgGE4wcHq/bQNGITAE4G7KlhPBoJ0J7j7
Oh1H5MlumIJwF+5uqtRKsxVqSO+d8hZxGHV0GdHQfPssb1m4g4iSLdO+Fw3+M/mZ
6e9wZWoRS/KzTOpVsEwCj73rHgeiQarUZ9to2IOhRFxVNZjrUjS6BKSnP27I7+3p
BF1ugy+1RK3OQ/WAJnKxmWcFSv5/TPNeht/SZrfKA9vsuDB4FMD/ltOBhiLkyFnP
XbaCOn0Pz7yedwt/UrYrzY036il6iycBARwT+eFxpOQfBdXgQv8Y0bFMVoRp6mPC
wPJTJQFuv6m6PaDXcDcRSRX5ZZlN2aJtdNaxEWoDml39G1WkpmBHRVvhtWX5SnfF
VgWxo+8LVYe15NVMw4YccDDSJeLMTg0JYGxV8j7o21CIN2DBcLD0g4LUXhogxOSc
GnDZw8sZG+psoFh6CUhaHfFDyoG6q3pCi6ymLcxHIIGtOUnZxWylqvl92ps3tGfr
IAA5S7+tedOtSbE+xvItv3kFBUuPBgSY4lj3QeQb5zVroORwW7RnCc2h/6oFxhtT
l2m76zyCGS6p4COkCOaq9EoM0eqodob5w8iEYE/9es80Wvkq4zKf3eAbRhBBbSeV
LunkBRNbhB885Wih9HDKzW/s7PoLTejOHKnWAM3aSJ6EzHsSJkJ0aGesURKHJki/
ue1/SRPSEKF//LgFc4pD5o97nT/HnflrMaPX/XwzLd1FuUxC+oFFXFR9UTOmaDku
pfjpykQIZLCu9JBdej+DVsMak6ghzJ+byAIbmV4JuSBnWyutovdLUMHaAwF6qkfS
JZGntzuZMcllhQ3b0eCPoQ6xy2Ni7XoFMIYU612EI9BwfOhuNUoKZk82XR0E3svz
UeemeRferm8wuYtpgrGEWqQIheXlYcm98R7uYlO8bqYowillri0gdOA4SukH2Jah
brM7AxGZVIjghRtm8ujcwy2tnHpQ51XOMyxKTj1eNQDXDVDv4q8cHwDGgHjdSCdq
fVSzpC6vcyY3yi64U3wxPScCTAJnbJyrcVdY6wGliGuwiSu0j4Xg+S+8bBjawDRD
Y9K4OYiDJNVMMzQdyS8jZkbGEDvupdiBXELQjrHvrMGzvGe87qv0LdqHUR+JLT+3
n7+6rVeVA8BoZXFaNnc8afF0Km/3XM4eyebNiwp/9YxLPqdzEmf89AlsnZA0RYyf
vbCEh5y6YzQ6HXauI1zsOUPI3FFbwIXQthv6Uj4g35OKpQIlsH0XyPhpE6oIQF3b
YmrkyXrvWsyA83yUno5sojv9gUZ809T9VI4yiEDw+7TenZ/6kxxE37dQCqFUAC+x
d4K6V0N7JAHYg9d658rY17BSeLe+plMemmPOU0xcOD7Krlr3sRsQbSYuU0Jw172z
fjq9uEzIaYJY1YyLgPNJQNYdbFHHEmbQ5W/fipFEEMxFnvC6+MEMreZrHES55nEl
Xtcw47DoPPdjUX5CZNSfjweYWbEuZi6h7uF8cWW7r0znac4bpdlGgmtB+2e7LiC3
SZOno7S3kTCHyT8GZ541lHjgFHAVXuDZqsdzy6ASdtJsXgraIgFWDVFY1PdGCMpi
QTadLSil0/di5DHSFRW7wVFLEmj2kqvpijmJq1irnRi1X7ma6+8wCaiKHupDHJEU
946BRKyFZadjW5FbowZeH6WsxOAHNFP72m2IphLnCxwSvQYPSUdBpPIC68AmfiiN
fWHdvmrceTx397g37T5N9Wn7teFgN46vYoTsn+FuEpFr/EDelrYj7rI1N4w4ukVA
jTjHMMch4XBqZwirl9ElLo1z/GT7QCn9bbW2bGn8h2/jB62vWmpqMXTMOgGYMlAB
dZnj9Zj8bx+BXqcqK9Btr+KI74EllJPF/pRqBBZ7/sAY606rJ9sDVHisSh28HvXt
k7GTramLc01D11c+2tU01guQT01sNhtTZ8Wx6wVVFwGfuoPucuZF9/uPOfvk0Oms
MCnwnGZg7UHMSp607rJEk9ufQv/klo5UHkz9Z3iCoca5ddQ6bsSs+5yxSQLBReTN
7HvG1oiXP95Wd51ATrWEtkPbJkRSrVzVC6FW7E3DzGD0qhCEBHU3i4QmXMRtzsn+
R0xQ3FhC5944BMsWhcRlQXAKeYFrgJWrmuiWtlq0H54IwAFDa32uT3Hl9SbYpDuE
baJMMC7RFQ2fWklu16p/WCWMBWDhSeXoW2CupH+6GaItG2p/7Hi8NITKOeoPteyy
nXmFwHfvE0t2NYEaG5ubJTrwnEj0U8h1vOOPNAwGvcAc0suUEfNhHD6wtEUS4wuW
uAIeZcwMe8dez9Q9Ht+rx/YB/C4qMAydxODJh5G9OMq2N/lI7ui0b4BQnLjnudUg
dgXlPsSMKB6Dfm9eVIa7K7MckWTtsBs0W2VNV/up31HtCq8JaIuFCRlqvs8slNQS
kdAKEEsLfVYpz01ckDvQ68vct2uSxFd6+tEgpIA+TRVliew0lXCafC0n/UHVvZqm
4rtshcqRUaaaB/RkGkeC4PMJkopWTQRW+bszE5ztx/d9XQbkOjCc8ClvJ4b+h5f+
oah27qsh2SWSHZFoXaNQSH1ah71ok8/VC+g3RU48wT/HbRAGEmGTCctD07MQZaT1
OBVeQIZqzyj9PQi6JJ9vu1JD7gGLY39kF0tFISvCBtdSm9kjxysETc88ARqtdiOk
J+bxoSYH+MydPM4s7INA9ZcotfoWrOBDIQhTDlrAv5hyCxodAfQTepLDLzw8qZuf
tTNGyZEj+ZX/nAh69cf437SGgjkU1Y8bp98yow90TWwaztSe9t4Y7or+YBRBNn78
xKLCTfl+yxTBL8HDwmgcx9E1OSAX3ndOfQYQHkE6z4mjucfjTU78Sx0bi2yVyDDv
oFn4/G/2Ab4Nf2J7DyPxMctS/HWb5LcTydJ8ipKUKNLDG/zXq00ZRQk7RRivKQ6E
k/Tu+8NWm/SRi+a+RCfpvhKpiaz6Pjm9nQS5gpCPatSFiyOVWO34H9hlEksgCVNF
AOl7gaXn5jE0PZVSO+8z/q1aez7ogKjPsIrfB1rOgzup4cILxACJQSBUGO9fQw3x
ebC6ckbLlakzN+CppUouvAtMBZqUTuOlnRd6nMXUrfqD/zWd15s1zSSwNKcFGdFL
dLMtsTtrVKqOK9/1S92DVlI+6XAqVTTtjuk7MezkBxV3gF2Xb6/CKZCSEaoGVfiJ
n2kbu78fMdGXzEhwawoQk62h4r7RalFq9nd7f1iZi1IYvktN+kQUTEqjtELbaVxi
fqv/g31RhV3IEdgRqHSOKDB7TxDaFt7nPOqoRqQ2T7Py/ZUeW0+ELI7nKkyCAqy9
3JMD/nRymHinhKdWkZUv+LbmY5UDO2Bs6tbhw9Bm8vcUhENz6AlCVAG5vB6kwHOo
R6SzP0AlA7YojhLyp/z4dIHkr7GGu76aoqKTGmzeddTYTGU7kSgVLVlq4qh5fv6G
HKIknaRKQxGRxA+IIDY9UqLmPCY5E352kIUWsPQ7sauLInZxG077ac3SzMK+ziWz
g/CR6KbWC9psubx86nAF9SUpQPfIqS76oghy74g4BuXyK54Pa3FKMTbLBs/PQLq6
wjSisSeanvXZU9TYTKoAbo5faPnH7jyN1kysdA5O0KGU0CSMCvg919fc/ldPm1ll
tiXnLX5Y4N5Sjm3cj0naTjYsQkZrD7AJKkfRZ5VI9Jc+xZw0X7tyYwp8R8xafReo
Rr6TT0JD5/s16jDJC293wi0Ja1w1nRyiIUnBAZZuAvFs4ctI5AnlGYi9KjL4cEp6
DYNAuu0yHiL0lHXOQxbzTkscn2HjN8Pzsl4ygz0rgOCJNpaLqmcOT1aZj3xS/0uO
fZJtovelEAWj64xXmXlCp5ckSsddTpTUqbfoEGVYJfduiarxMi13I1AaG0A0gID7
+OuL7Iso8hbl1iVfbZ1p+/tJgZATdMz81o7sILaBn3On5jlXLm87yrGB+zxYAwx2
vmPu9GY2xryJwdmcGYRYZoEMgWi7V6ZRobBrys7Sdm7Ybu2chnNkYbfPQX326MB+
GGmOnrdnrP8cTQe4+kutZjvYTDpZ8McKZJHD5rum5O29pidWLMmyB9253wwB9Ibv
e9L4guC6vAnDocJUTSNMGciRv6cTHQbnmpLPp3ZkxB1ACmAJiGhYhjEJGAzM8SZs
9vvrq0f6rRYjUFxuv4ZVyNxd5F3Z0Q15EdkxuGWAVZScZ3DvAhfA/SyHWvy8MS8Y
rSg0kedK0bihMzamw0N/XXRTzmafTDFwlSRNM7PdyfkZYrZnSTQ/wb24O6lFuydk
+NRCfffAHa6QB1nAN413BBQ+rOeHCQnSa9XZSxKVkrTsVBFkdfXUg/7ZWI0UstnO
wiHQbcdyX5+R1a/4tIs6ebTjIa5Ac6CZ3cNjQGvg7ok8cQ38e2Y7FtbecuWgG3Js
j6B3qUja9B4tb8hdG7I/oTIWVn13hyKouzBLD1aK56Tr+Lv4OxkCbmgKCzpbGhGE
IZdYRqeNi/TmtBPCYfAvhvjsxmrfqipQ06zqFE6h2eb91AE1PC3OiYAW3DQZypeR
xt1YuozcC0VKFRiTQQlVsDgOYZjKGZ0O0xBJR+aTL6iMYaaT+rT1mCBEC61vTbDD
K2sM0IUAZVAPw556kgvgCISq6Ec7U8ah7+TFO3sRBNAH9NJRed7NyuN6I3wYOgFw
r7EKmoLFczzqA5VGhO+f9p9lJHPkzeDb5pdHtvxp4qne+PWtfvHPeWMrTFqCOEj6
vgMm4UwaiAntfaybO7BPLwImUiaYuOgSXvEkcCSVHtAnXher6he0LlXmXJwluici
Ovvi6o9I/llMh9KRTQsq/JwA4/IU2XFzb1kgwLjlKSZJ/5GkVHZXVmtqaWFIpsNq
yU8D4GUHtjkeG8PvzHkt7GxeYbAJQuy6JFVuXsP0Ksx7lvNm1GiSQhV66aAYK0Yy
EQxwkdDsK09r0COlDSoMOob66p7FNRkCIBSnlFcmiieZoGFuAmq17jIikmJp8hlo
VpDF/d6LU1uM8MibeNCAST8zxucBLa9kl2IVWWje+RkYK/2u+ePesvLxI2haJIVK
QKbxprYk9c1Wi2NUvJMQ5oniYrGg6AQQmS7AzYN35P/ly649XCZS/ZcD5yubZgTb
TV93Qm6Q4IAZUQ8UpexpXyj+KXudLLumBpaKMKjqjO3doyL19F+UgNaPYTirdteo
4glTm04iiasjxcqEGKnJs6xA/6fbcn7YeBdJew/JuOwExEQSJtuVc24rmKqlSvmH
hTYana6DwoUGbrM+mgG/lICYHhFrvy4WdELkczY3Bn5n3MG6iHeWFX9vSfHJPKqX
tn277jA1S9HAWqeaLbc8qoh3E6+UKEt7MfttHUXrTd4yz+A5wLpD1rwW9Sv5TpzY
9eA7zy9JC2b4dglc+4Cc6wo2MjJj1iBl0P5AnIWlFuAJDzjKJisFDc9I3cqsA3NU
ePtKLAdDXqkDI1S6ONV+/kfgd/ZeKnztSaxFL/RrASAAo3eHWZh9JP8GtSZ81a+f
xymBAj+Qc4npltkTNrzobffwFrhSWzn2+0q8xA0358CHGXyc89ZJsq4PSHlxgrjb
jrs0BKC80aDfpceBkPDB9YCT0ntWFnDWvVspl9XZKMgWNQ6cUXHuGWt1lcVa+bnD
W6vpQyXgOf2CxJUtWMj6PXIyWhvEZL6RuqZ5NTYDODMjeF7F6nHxbvt9geX0JOlN
hTJnrqLmaoYR/fwVCuSN7cSNOEEupyQFz50PSxOnOBK0mf84L+lfZ1ijgui/L3En
pSwj5vYL4VwbxMpOjOFEdTkKpSZ3qp7EEishkEAdnBjtzZ9/ZLbNLUisP/9UDh1y
hHRcZf7XIIHwp0MC4J4J4JQxEN3c4hclulAbghXb5dBpswU2U+9BAPKgJzL8qbsL
Kxjrsul54iEae1b26swPiNWefBL+bbEfr4RY0llESLVCJXD98Cjs8oeWd27H3N5x
sSOcfu3jtArySJnhZI3F0GlSO4/fDzBA0aD8qmpDXW7CfUit/PhTQ5oG2qh/Wx0r
vu1/RZ6g8JqP2/gq3EFiZZHEsUv8WwAGbczZH198gBMIQqkhh5z4llOXN+BTAGvX
+Sp/lS4fGqQo3mWnCdgHJtbiQtxxZA8kIA0mRSn2YynmnJ0WqwVzXTJfiqCGilZl
MNazolrHbCY+Pdge8mFboTyXboQPIRh75loVXLTIjk2eM56zGXHo7bUcNW2YHIWU
OR9fdiOoDJt9kwztXnTuEvVBQWRiC49ib14l1LV0L0QZcZ/GMsZpbLluo4El59dy
z89NjqQlPwOTI3wwMJ47RQrxLH74FvvqlBo9sgHvw/apKptZ5cEZtIJMiy3hNvBZ
cfE0s5YKuSDpkGGSR5xZWwhphWXvbE2DRslDkzAS+JA+WryXvdY2yY3WTvjUIvdh
oGCkTZQ12kQBCRueN4JPxBhqfVx3I7RvTr9PrBupaMm5WVnLm/kgY3ogERGN8Fw7
x2pZ89Fyq0JEAyxG7o63532Fe/rvLa+BbSTI/uiLktxUsqxKR3SWLVO9i73k0fcG
WxYAUsWyWw3Z3/E3jdHW5PA3dFpzprZyhHLQvPoYEUSrnmY2L9qoPScbx3AicgQ9
tQaVQxeY7jFInSk3RLlvrg2v9P+n9tLwQUSxFqJugqPE59zbczvXDiHt4YR07KFo
odnvIc2/yHGhCHiyj1tDYyp3vnnTs1Qwh0dl7rbHI/3Ich26SR77GUtelhoY4/IH
7TF9xrt+xRrAf59gDvBx7jrLpTGFBwNZYZbpFG/Ct+oQYBjSAxO7ZQaMbFphlAZc
wfwOFboR3pDv8E9xnVBUHEor9q85Dmi56yX0KWVy+X44xJftmwaW4kex4zMHji83
QCF+o7zKNkRmH6Rw4CfFcolK1nMM0sx4a8SxkbvaZjVvH9oNjRFfu+ideOVroye3
V5QQxH74yTNS+V/ckMy2VQ9tDHkZMJuUxrnAUOIA9/SNs1a2OIDLubXxrBIXBx1f
dJvi0NWrLgksMs6gE0s3mNA0eOmp4ox7tcdu5hNWO3LKXzSV63wCOSYpu7SYiiNa
frrVAgeTTJgcmVWZzmOQS9ndKwTTvUZtmdEwnyt/+TqjiUxFmeu3GXNsCTuu94pC
fTbv2q4ifCnJIkARiRpmejKi+lkCS25mETkyIT9RpuAjW8WAIO3z7aU6Hn/hBgyS
7h44xgl/fVT1VBZlFm3HIemals3hIe88g4LKG9p/0u3CYCkPVUgSJd05/IerC6ao
pHEqRabDMtQWLxz95JfGOBS0MDNVkkbN2mZMzTtW98I7VTyHCydKbqKwYdGVclfT
bp0cKPNFc6ghInVWhahBElLp+x/asAJBNHij/+cdM6V08hnkV5YLf/rcB2swG8/P
5UrB9FL/IkKCThCbO4Qn+z5NqhOBSMc2y5vFlrKDV+Z3cy/lIy/DAY2BLe4KUlc+
u3zEx23eh72xYdUCWylaQ4/liRZDOoLXeAezBLj9xUG7tz2F2XIRnqa8ohovfTx4
WHGw4j5/WaRJkSAM4Q6f0vQZFefl2qN2Iw+w8R01jtvszBSy3QIXILIZ7qmDOK9z
5fUc3rbVL0o4EYtDq7PJFGAzgmqn3IXoawGov87xDIBBJIZDBfxogmk6HBXVIl2U
pUXteKWdA/pitFy2s9eoRZVUCDoarti4mEkqECKQtk/V0umbDaWFshuyBbFs10eM
OYGCGlilYThNLrJqgRR8Y5Q09MJWherYMfcV1Lv6P037yGU2kGeXSaLxklVJzbGK
2BEGJFXM6Xv5UB1IdCtfBn2qNaZihR3BFpMEkCEEzgNY8In2ntlu7VTsejhRHKEh
f2si1zTAsxBGyxvMzNHgqzWbZOSOrdMCfEAmA4uSw7BbqzCbjmdZ0nJLgWqq3VWC
jDZJgRALSCDypR2vVv1j4BDIZoUeO3wKgvR0sekeVMnbIzIv/2paGfCnTTycEdpT
SxVUUdhVeyWQozh2FHKFKKXsPfcGEQ+uQZkVStTQl3tYBremLlYukNivZNIt6lBX
VlkJorLCznlKTJp9S1ktaTJWJmE2zoruN49qiPPFGjFrKYq7ZPnCJttkJ0MvDRR6
HxREg1AvZTmM3/UJt4epoVz2e0y4pmFMYCQSEX2dmeDMk47xHOZsWAn8ahLk/aMo
UZlsV0DYf9hMCjFDOzLRk+nSu+PvDRhrcOkuM1Z/uJyYb1R/i/aHh38nnfo0j6Ce
DumDCTUPT5gDOWATaG3lTMlRPBdU74O2RbAGxmk/ylcO2eEOnoQxrMJ3xQBd55w4
bMVw7AT0irXuQ7SjqTk/mqfeFYk8dhIiyEl0stfN2glakplatxUNKYaMrtVClpmP
jBGOR4jJz1QrXL8ZVDzzWr0MFcZ2L/7rbZu/+WT8FZOTkUkW4fhvouUUSEiDu3rc
C2HwO2SJ9AXUK9vObbk5z8/1FdCECLCRvUO4Of5RkkPCwSWspp2T6OmRU40ALd2s
d/2sG0MX47Ns3EatOGXydqOLSzHnGv8/5kS38rMUhQUfzqWll00YFCvXDMBUxpdN
ZGMSDXgyXHICX8BW4ctx7wDLoPcd4LqdwlBYHih+irwZPYe6kHYug0CRFpbeL7/F
PAppAGLaXd7viUCIk4X1B4aGj1hnNCHSXCE0UQY1h2eL1B9qteLp5aIYJ8gluh94
yJC+wzv1zrMnb22Rqe/LjNkjk2txrv7nIq83WDk17V59N49cpG8DF/7IHAGeZODX
ZG0wcW8OoAQmcoRW2OFRka/lzJpI/6ElHvi9ieWRtZxV/C53nbGs80+lrDGYWWEg
PJ6XQBZMHG6QvHjZ33iS1ZLz4FUsZNw6Uw2e/oiblyNgQPh5LeckvtWVHzteSGgr
6yM7G0Wax3eT1vYiroAoi7wsTfkwemNZpCXX4zDK5jCR6yVqkF88gERCcmeNiM1h
MDid0ywDNWNmURqMRwglVfNVo5pauRLouiMd+fIsSsFXt5Oxw5F0LSnQeEf+ObUR
oSX69LBQO0N9ckCXBK7Zh8Mfx8zWr37Gm+2Xxs8DIbatJAY+8FI7EwKtyDa1ugzI
I2KnwhCJUE1hNCyQtObIyuaLVhceUaT+bjP9qoM23BY/oWGQhfVoI1Wxf6FDQMGh
gN4DBUhyZqf59myi3L7stvQWljAk834qy21/NaVaU+HnN58c8tAshSoSO9gJhfKU
dMhDco1So4cPtd+yFveuOS7SRkkFPgGV+6QK9QErb6YvTJBAW3FFpG3fFL5cEOAX
zBNMqOT7lvg0PeeJx4wFnFQx8Lzr81Y52/MiTVhm1WBgHZLAkCHqleOx08x2b4s+
5CkQWriVLCoEm3bEuoYsE/T6MYDzRgj9RDLac87kEDgrZE1DCCjeTtDJVYbdSozl
B4IrtwlqDujx4dHDyW2i/CxAsua7F8UgtUJYx4SkcWrJCWcR7Lqmb0GshZq9quRK
cRryo4priJIIVgys94RaWYodgim+TQEm9cQUFFCR8K/kFbvRCrauUT8hG6iGwwdR
fraNVvkPJtSPWpK1pqKlF7vuADYVKDv2EplAXJ5Z+8ZvTCFvx0B+Q2vcHboJIs4S
kXyK7/lJJR8Wy8wI/UUXBJygWNTtYOY2sRZ8tJa2ST6fNNONKvXAFdEw+Xhuucao
HY3p9KetBYap7HD6lUI+jOtDA8TPeojqOayPt4ZyU3gyI8KMGIN15O9TxCelaO/Z
15e2fMCY3ECPm+KJdxZu3+DxYJ+9n3DGuWVLGWj1NnmiRomZF3XAd5A1w07jWY8g
B2D0hH+BIzb+S/DxqwhntZbaDhFGgTIB0I9c9D0zZxe/7k/hhfky7AOdWP7z2mYz
28QTkRaGdx8lnQhRFJHV23+JShYV0qAIsxJPRnyHFrxqv1TJP+zULuBinhldsq5E
l2Hsw+esencQGQ7BXsHN6WNxENP0Rw9sT17ad108UvX5gXTKFMwHkNNOdNfrnFuT
YTsKVX43UTEcxtEtoKoEqYxtiGwatFfMejUDcnZKsRhTYdp/spzRlxcwMFubJtU2
zEicLvr6xVa0cg8erJcMhJ1L1ndKGhsf7dKhkE+9jUzeo//GoK/6djIv6apvb9Jq
x4AME9Vr/5Oa5gyh/UOwiDgU+dSk4ZXzMf9F4eSd63E8FXmFI4owFTdr1TnXHD6/
OfARrJERo6rChIQzXZIwnWRHaZYR/Z0LBsaBM9QLjHQo1LUy9BlLxHuFBap4scvA
sVobRqnr7B9pWZApWI9o1ufg/UHb8Aq5o7hZC/En5G0QUZff5Ta7tuT2b8+XHu7i
VdxPnZ3yKJeN1+HnQBEtYljNn+CPUhCTRHIBO304Ym8TILYTATg8MtIKeurdCWQH
AfNkAAM9/WS5CCLR+FpmMNgIhIg26pJfwIuH4vVjJb/HEsakq82EKmrNHCXuQea8
Ij41jPErjlGPOvfwnTpi9stBfpEZ5s0/TtsLdDYyTgTb3xrvx+20FT0Mn3/oFPUO
WX0f4JKLpDGtjNzY+Uw9DV+5hnQVUaf6i4YZsyCtcWyiD+rIjes9F26tP2JgdJn3
16vo/JX4jPX2wPrRgcwKIclhUpDrOslnRWMrEEw9i1dQkR+Lj5mOqs0xnzTH0nBq
yEIcjFF+9zQEN/+yzQwJCEfoTLJPFUZ/nZrorEeeOUWoXeWkJ5ppuoIfKRpbCliQ
a6S8CG5cfnbL9H8wWxED/ggBo4VsUfdNdCkE+2aF9RhKZlxG1OYTvxPQ0IityoDN
TT94UVWW5NmqOyQbjNBNd1bQ/1aLI4QVPe2nbnSaVaar348Gn/+Nf2zN2jSNlIKA
etAJkCSbGN3UKHZOxJMjkgzQySlmUz0fh1YRqec5i6ukfef1A2lV3LrsKMnrR4t1
LpBprx3h+k9vSDDXeDMIKk9cc7zjEs4KFyiFvBf0cN1sTTHOkn/6RlZ0ByOr4Xur
BZhy6KBF2Z6x9KG9PPrjtZz3R/6UZsfSdYrZI0uzpomUpdPZAUr7H9ed6frWrigu
Fe3Ycs1nwxGG7T9aNCqdq7fmEA32e5ryi1srs/BGk3h/X0tdEcGfbJ7sgZSI8z2Y
6yYAgTxhKssyQr1+RSAhPXvvxLEBvErECvQe78riDQ5uF20bMfLRYxMsx5aAFm0V
MXJPPn+COs9CPrMs5EEMSH2sAeHSBqnzdWTjUoy9sBnW+7SNyw7Bsd4uJWRIsdl+
cxp4PUVtpKYp8HlaXzmQfBCahFA4MXuy8qNv8OGdI9bouHp4nghwcFYjfAr2CpO4
HzEteSy9N0oykgVRcBSDMALsccAQf4LQpaV3z7m8vRD8/upCd4dDYj9h00LtJhwD
QT+/Nq/kC0Jw3iMexXqYivXro7lWH5ehlYMdcdodbI6tk4hZEiH1nYYaLLQeJ8Gk
KGdEddYCRAk1ZAPVJQVNntX7sCm7+1PdZhuFmYUXSrfMn5kW3iNC95k0tj0xQgZK
Do7PKGLDI4MgUWhitGArXwLXo+8Kfc2CwvUio1ikRa62CCC7tDZ0UMETB7uQBu9T
51tsGmqKlbqhK83LQW73UJeuaWf6Ba8S62NxDXGh+7K604uS3o6VKJX+tcrK0/pi
PYBRqY6/24RIsv369LoIU/SOt7cW1rKkNJjl2OboNq0Il7uQGUxmq2A3HuLqmMNf
NDtgXJ7+Un6SUOOZq/A3Cgyr8G3HgNbJ1nv8vJd6daVe/lFSF7Aj84orfr1SzS+m
+Fuzn+msce0Yex2OUacgDxZh6GW5FVGVjX1O87xipAgYDdV7B5E7ovQ2pBYSZZ57
Pb/AJWppNyrrjP7jd11HhCcAD1YCH3TSsJoBf3yb2+w90mY5uASJf/9KfMdeA+t1
sXBebj4S5mw53PEhv4ykc3UaCLpdMcK0TrkK5vEksBdafIfI24T4nlUNvbXlh0le
FB2jN/qr2jPpcOBHegZjXUnj5YCw9qiWMfpTo6mEt+ZlG+mzICB2RaX2hm947Koa
Sngw+0kSAxaZ5XYDZAFyVN5WEW8J4ygedmyXIEN/PHBDGR4pUYgok1cFGNA5DAsS
GdmBqjncxSPgTULnF9Emt1FoPRRuCnn5xEqu5vx7HY3Se15OSHztsQ7slxEpJKLr
7kJtmEnQ4h3BwQVWpynFTAsBrUVgE663W5z4uYZiApGAcrN1D9FTHDsLuk4pcO6q
YTOO9iYfsniAjN4IVem0x22Ix/0+iWUo0LFY7j/CREKWphwK7SXsen91l6yr7G7C
Ywa4UQJmqpBDsvTHivLiN0FWi08PIWnw39VEivsDflikQQkk9G6dnamRpEUNoegc
kD+tfDLjJb2Jp450mIfyDoRuSSqAmOm4E9xwDLPAhmC5/ORPq/pq9iw2OnyftL6P
5pHRfNipI2Dy9+bMM2XRWvgzTcwICnxNj5Zxqxdm5yhGTXgQQsMpJQ9apKELlQ+Y
sr0lMAkskvz4evdoCViyJgT/e/TKax0yAcCnp8WXrRj0a5SryeMio3Sm28jthvDP
70Ddch7t2ic6NoPSRQ+bxn/UPxXXRN86tO15uyXV9eHtTsPlzz4ePYwXQD5G4KZZ
Fkwmk5Gh/68PtenMj9sYxkefQY6WrlYoKR5KkhHHjTjNM/UTRXwSmBGevEnXZ1PO
YUqv3RblH3PYBUR4msQwlYpAZmITj5/LqEtsvFiS7DsWd3lg1Iv2klgRmasAwAp6
YcJJv86Cl1JiG9jp4UIetDhiqt0Zb+vHhrQlR2OG5VKVfOGdHz1NQWbIXS0pFJlb
hz+/8d7qbuDdWxrmPSM9/X6iKShVH48+9mN1IQV25Lnl4uT5K03kQkI93at8WAlq
qeCHokLoXGhQwA4citElc7EvUMHXKvdGPX4hp1heP0hldU+ynUD4dTRliBp4L/Zr
u5VQ5DJtS0k0+cRpSPaULU47MqcfZ56UIXIFk+9IpSNZvBy0eA/1obbo8xxHXfkj
ssv43vRUy4BwEz0uWSsXwTiL7I0qh/HSQC0Y9i9L3DnvdPfKDchs4UfAOZzVkQDT
FLUTIS3BqURHfGJIHL5GgvObk5a9LLnHbOOLRrvZiIW53rmOsjgm6ouVmtiAiY8o
7v4bCoNaRDdi1j0AY2bsp4Mtg4vvhsYW9tI+n5ONzptmmdzRWR7YGvQzP73ynh6S
ufXyofICIIJNR3oo6TkRKLqNMDERHLhlBXAZzmK7B9xB6EdNTSkTyMK0OCVoYMF8
36TRAac+DaKSrDYANMerN2BTZv4J80TF1GU9Ogt66x4EHLVdIclXW70NgyJweS04
JpktnJyTtbU08vc4zWcDjJxw/d46sUUxlNdGeOovQ5M9i+9vHaRG9DaTb5Xv8/o/
0zmDOlWZ/si3oUsIluFqp8re5Au8H+eZ+oF3xF2k6yx8KTQr/mtDykJzdP8OkwmI
qN3ErrXtkIYKnw6TF+dhnPB1Q5rMRFOjf/s6erNkZZogBH+tmzgEevG+jSXpXKGr
zGEXIkRpOrYfpa5PhevdtUb+10l+th0anN9RHiR2ZhMp0vDzmKZAbZIgNf+SNBkt
/QVCjnJtDTTtZFWg5I7PBVeRjOhd6XsusR9jSqQfU80rMvStZGIbXVVRLTMjVJ+C
UzvZ4KbPT8lFx5sfKsF+e4vJbXC8ZmUKBhWlVgH3+Vxd4UPZTCfGnQL87WJBeN4h
kdk+2Oj/b+CjLTv5MptEPh2cQI559LxoqLHF/4mFrfURE6pp0DlBotWDsTNmPlCS
+ALK6g3HF9RYbvayH6A6tfJMhe+bZjyHANN5auvEONm3s28dFnXzPbWCR8mMaQ6o
56WroCY28N8DNVC8YtaoeJWUv2PvJTVDyUqT1eD9ZrEVIZGiG3l+CQhUlm63eonH
ezL3PFZAtpetU6nTfYzhYpaUIJZDn5HEoRVAFRvmHT8m5RjnjfhbTGuwFBGjJ2hm
nLNJqgrbrkEVQZDt7quRijnaUlUq25UWY4nGlPwjLDBz8SmOKX3HYFP/E9MVitkk
gEGevqVH6LV/fPwNljW0oEds4osHLy/pLalSAnwyIiFTxBm+CeIGRe8psrQek1iE
s6/aAfCG7p/Pc11Pb2F36Bcs/w3op9oscXezmh9VXVd3ID2e0YOJQYqVVFlYMUwa
sZpibsyP35sCx70TUZx367IRycUvF6WXjGKcTPBkolWaEEyocli67M9Z15mshXHC
04kQuP2s3wdSH/kWnwLS2FbTzdW2Obo+J9JxKY1R7220JWme7x1XK91710BK0pyu
q6topvx/riJyYDqdqXSdX7qHvlNk3F1svVIDkzQ2muFY4ERwXIoo5RuDs3zVnsdL
aYbLI5ND58WMFL1eMjpEBIQGx5gIS3wGShfZKwS+NYSpwgcZUr1UGq1oBVfhSat6
h8D8TJxHTq+1XbbT2oDYsY9l4G5JkEuDP2JmCfAUbvT11TI5LxpbpfjKV32Kcan/
C2JT/hitwZsX1YuMu3HzOBLFuSqClzxFihjNDXfLsK8eu3bNB1wi/ACRvVXA3AmH
b3bvqOqX899BHSnva7j3ilyRU2F+2clo726PlZ68cIhMcx7VknJdCt61ipzrUYhu
FheRE/GOw5E393jPIyIv3QnFSx2fY5EufZ+BMozU6CKF75SYdBXvqZ8DgPzXG6H1
iSGWgT9vv+mLPYlUqnh9hk8Z61qXu9wqaRxqSUPGa+Go2j/gdlpCpmgWObVjLTSs
XxgGwSRW5JV0O+oQ4lTXUttrqsH5lU5RFZKH9SKAzEBHXCHTFaSSK+/n1ztrJ0Lz
zbyGs6fDqNYT7uRhyPl/hYxm4KfpOZqQb1eXYdZPcfCAd128ZAOK2TgVnic8i9kD
1IpQ+IwufvNTjAj7RULzj89xBl6rebhrsZVXB9odhMhoJf7zcK1d8EkjrtsD+3Ls
kmy3PE0qb17EeLwl2QF2CNV706vzmBh2RLiyqh1OL266JYLWy13RZ6lr9dp6l3dv
vLNBV6op922mlWWf/zGGJG1fh/n3zaTrraOaFEAH7xdj8AN6IJN3M5/GPsNc77z0
uKJQ/As5G00x16sm2GKKIRwOjQGdxldfkJkUVDPg2VKqVa1F7ox/eyo+Ew8Hl38a
O/vABqgZCqJxE6XIFtNB1tuv43NE41p6JDYORdN5iHHgOOEmgZ72MaTsibBrqAJK
/sYBv6Tx0jQFVInYcD2phGs0Ch6obHp7YG3ZVy2ZvD6d4HwrqaRQZ9FHzXis9Pin
hvIS3UUWO/4oP0hk5UPV8UXfs5khIbJwHdxeg1EyBFLmkHgRRAzN8LNpAX/MZ6ji
dvpS4l0FJJ5BZsPQXkw8gfyC4fW2SxhHSfLNDe6gbm1GXB7ZtO2GM4TZirh+BlO3
e5s0SsOuK2uGruTREu4RwY0yF761KgPumCNVHPbD8v5cpJFzn9ORaPz+EU4JakhV
hK9rZSO4DQcUGcmzkVmEceXvdsJ3fxvhekKM2C0P1n6m45SP98E/XCs4DcW8ulNS
ox89JT/Tktde4Tdq8qmYAlqyzRHBEy8s6kq+k8SWlP6Ln2ZIjw2RTOuhgrF5DIYh
wDE9AEBle4wQx3e6+aPl0foWUICQzhLZSuPfqpah4EwOYY8vgLE+P9uZNa9Zzbd1
6RfE7lz3WNCl+AIpUBMezWbiu//qEoSpnP3VfqFIRdRRpWszIBFT7FnA4SWBKqAV
NxMGO741JrLN+DHMdHWu+lT5rhWBgoRS3FKxiMKFHcAbcGe5jxpgXoCMgcIOyeKh
JbFoz+OUwQl4RGc8p+WIonbdUjynEq9UpOCKuevA6bly1eI3VTzWKc07yMH9zq+7
51Kg8FsdciC8i6Jx57A26vpk7RGsS5zZ1Bw2PkIcD6BZjhk60Osxe3wWRpfEbdZf
sXsW05tB6iGbRJ8Jzxd9Ly/bJg6jkxlMedl+14kL/eqjrKW+Ms5qSkMYPRxGnnb1
QI/00goHxtMsr4calmBuueoyZWJWTIXOxKbOMVqTgJ13Uj3CY0I0FEzYvKtANn2Y
3aEPWZbCfnntb7ZTpcI4fUxZHh/S4d4FwCfjd4o24kyZui++fWsVUPLl8piqSGoL
tvyJ+PnbMqMKniT4gAuZRhLn7pcusMZmKHNq23Vq23Z6FrdHM+Gv/VtrYetpeILa
IdahYK+Kovd5YPrFbF+UtQKGr8nk3kBFcf4QXVVH653CDOBkDc3VPqQTDJaeUCqC
mbvlVqh4UggRdNQ/pigVMefhHaaGoCam2XuWuvq53TuR90TAG9E7YrP6SK/8Ezf1
V+KM61ZLojYpp6U6bMhkh3TtNZr9LV3PRi6+1/jU2muJvorqWFhlayPPs7N/cI8I
9GJvJ5U5yRUbBELZST0KrI0S2tQp4EWAqiukuAEnXKF8f3H50M7XrPJ6G1qJN98y
L/knaV90dqp3Ne1cXmX3BzLMPVaIVF7RKkNFrVQ1TzFR2Neq3T/v4egPwkUBTwt6
sv9RdbxSXxa63CkHSx2pEPETg2FCfW6EYMULed85cRZRwgsGA5zSk1GEsI0BJMCr
RDUiuo09ttlmjDn5shxJwSXlSvpUYmM0B/kl3hFOrgPddZhG/RllbGEucoZbJeU+
HHtHJ1xsRAjcc0DEHjkQexBmhk4j/SGLNzPzd/wvDmKvBiKb8cVp+bhkkJO2JqFr
GSc8PVb2TwojHhqLVx5LDs6OSiNdY+y6kR8yY8XccaOgcYa+V0rTZWZ83ehNSSG1
3PjMCi3/nwJsodknvG+WM9/TuJ3eMgJFIFttB9/lMFIll9Fh2VObjMmYEYLLDYu4
Gwa9bq4rGUmjRMcYbDGhCI0YEkutp6dLngGAVdV3TZhOQ/m4VQypoPoLZyNkPMLN
77EGKDmCc9TyP3U7a6EtaArueUNRJvsPz+j+pugdeJEWOKRdewzsF4OyPPTLNC1/
22O3Q+/elHKuvn9jupADnoaNCurjD+7TMy7TI9v7kUtrgfL3ESWiWHs0EtM/tE9m
bVjLh2RUvM7XKhf6fGlJ/kXJn6p2ijYi0cgSzNNFtCGDE8MiKa4i+0kanO2yBgRY
D0mCdw7/2kd/aFOpVva/LwHcn5GQfnsPIZdmTdbEFyWc9V0ORIN5L1XsNYlUJmqM
QiclsVe+P6ZQAKZxWr1iypyrZaA0b4MfTExL7Pep5AmFiqeYI3DSZxjbd6SLa/5W
QwlNZm9pkaBNYAr5zQGIudmJykfuaNO0YI/KSHuTdpoNr8nlnDd47eDk8ZIG/E0r
7eqjk3obbJLLRTJ0WsF+mo0Ut0y7xCjEGb4LuOwLiYg4IlckCaRlI9L2lN9ikz1q
xRZ6nwo5nh14sGw2qVGCJi+2eeVF2aNTN3UEHFfMaLHTDnAxN+GdD4xFNlbdKqfX
hI5rbrNWQhWit5EenaowGz/EtTnxJ3CZFfUous7Mf7HIKpBoDaJvEYNjzz4fkeDg
3MtLWMx3Fr/kLrlgWKhVe2gU5XJpv6ZO40cj67oRqerqRu/ekPILgmEo03crz42c
qJg3amuzW6rM/oS/XtMyM1QW+0sGLj1SFWKn3BszJy7Qui9sbOn86Ss6LMSjtZMR
+y29CA6R45qy2CBCrBefSLNtTkW+NTEUzAapRhEY+gMiDbSr3czTyHePIDpIqvfg
GgmNeLVUQKKcS2ZqQKPQvU3Ga4xhsUqsCemhfsllE+IfVN6IzwXlCOP5l6hWCRAZ
2McUz2uzI4RguvjIX8gba+XiThUmHqJfTceSB/7WGZoF9CuJ6R0miJWGvOuFbYbr
4+A3p3XmjvIUyGVyhuOTALCyGpmVKWZ+P8ZESV3whdY/ZNnJV63LjibiLsxDeX8G
cwu3rdR7iAsxY9rkFZFmRQl7VBg4wRFN34dISjB6jgKnISnqJCS42HPdnoZDMcEc
3xM2nIOQI1HMy4CaPqswtHjTgMyQJLSVWeYauVchVan5o85So19JSv5IsYOpOPwL
zgF6akoRQZhNXVt8ttAxxjVpjLMp3qToWBclER6osNf2cbysS4Mu5xGXJOw2Yvx9
b0BEv99+JBUtBI9xHS4r0RXvsLai4MBI2sc0Z4ZCxwcK3tWq10afnNGVjZ6oujvN
awyggVpezn1S5ySUEAJixsdTeKVkfJKqV/sFYbljShg2MO6Q/bDtsG8yG1rw7KR2
ZcvrWRuS3qPu/xQu6EPqi2GNT5XCGNTK8WpURAUDFNjiw/6dTt7arDCOWGxDwceN
ls7/oWTrSqHeZJeFXME0AsefbMeDW5FPDi8TTmgwaKMktcd/AFnr0nI5ahCZ73VN
Fviktu9fd5L0M+LihNyKw+k4RMllZwPxGeJFEyCzKfWSFT+ywS95fEjMofOrl5XV
knzqaoa0jYiHQgxXQgAK6WjW2ym2YbS2AgGiDP90V7rHXxRY142IuPSX6Lx/1wGt
+CWHTRQ09n9rSL/7d99UbOGLDyHGPk6/rs9jpOYkKIwyhtXDFaRH6+5447acdVq7
FvTv2Z8u0t40iHQPa6GFkL7JiVJGBYYsHgDujmYGBuX1oHyOGG6MIQlsENITMN56
BYodoqc7F4BWe7EQuhKfQO4QQ13jvhWVWDfPh6GXTOVTsMzSJpgW9MI0j1/C0C4G
WfPZfVMlHyuYdlT2Yn25tJk5b9LfAqROM03V6EaR7dMrKlmLwANopzQYhTHp7Ofz
gu86jQMJkTJ9o0cS4Wws+E5s95aZywbEjRw7RqW0/VdVzy2C5Kb7fSLoRTYlPEE0
SP1xZHg4dNwATL9lt+56v7pKEfFc8q+jmDkz6kgIzpwwhyJvWTLAe4/ipVuolTU5
kKWR1V6ff6QgSyPxF0cZTtnnW3/C7YJjJjCgvguT1v8aJqG3S097ZHmy+kdAy5jp
DbWNM/SP7guZ2MAXdWx2LZJ8T7jzexJ0lw12DHSFp7uRup6G+nR3FHXGFbDKxb1Z
65xMONuEHVCwB4CX2iTAwrj4xkKu9rIcSCPg1D+ik5KOelJeIORGYYzIb3fhJSzO
YSdhvpsF5Aj8jkwKYgDn3os55p9h8riE5pZ4bjlkD/LcahWwCgFWP/llDpHW/5Wh
Ohgf6Ped3MkNpam7hfEK3N10B5zukqi9s8EqehMreAudLu5LtqtXFykMH+jIhrSI
biZJebfN5bAen+UJuB0vkk26ELPrHtcJxAGslR2nWGf5Urjx4djY/A1ut5lzGtkM
KTZlBNTnm7ZepECyYC9pGl7KoEmR4oxXVzPia9pMGAGos6ClOLKSv872JJl0D0rn
PVKKVh71mbY6sxwN0rCrFAfMG1hG9eblqoxc+vtXGtbl5/4goDzzQlCBBhF1hzBQ
3Ee3bmuhpOi4wimCHx/O6xJ9fcyJWy1L9ZUOH4jQ1+CnDaqSdSFTtDvYbrvymDH1
OFj5lqd/yQL40Jjiew4BbxtD20l5xZo1ji+DP8LGHKUlgjSzKyPCozn7JWUL627C
rOWoUmhCnSLAvgDr9K/bSquKIbSuDAOCXqBuNnv4T04geWAPWTqNFlCRrJOYd9C6
vKhzMAwY5UNRPTWtfvOltjihVgVh5s3/+hJqSH1Hqbh9UKeN79Zm6fsHaHcyzQZt
EqcaTSdK+3OMKljsgG5P59/PnxJm5Bw+dBzNBdZTXnjSpmw3sqqTQmpqqL7LifL8
Zp/c1TuKjL4/R5HazKHyDyIrQ8+Tli60I4cc2yqnqrowL1k8HdS7y2Ts5uMw8l5V
DVqb5vcjg+4VxcGqwdvkOmw+whZ1W+8FEjFxDv5q4E35lE8RuD/qTqw+mU8GqGk1
oEdIuS2Y7/MFOJ+SyQn1ByCnoIwrpRSY6XNjABzG/v00M1N2oyPZ8rPEuWhWw0px
1L5ZX8S4JhlhcSLvXnRUQiTkZJuf4swir1QwdNR1Mh4abg+3Yms8ZJp816sy4SPz
wQCiXiI4q+vNQXG/6c1dM/H7p42j0f/GrEy0QbTKYNTjuIlLY0x3Kbowwo2JWvqd
SQXIqQwsMAbf20EK45UZikJIKx5JvKzAbk19p58V9KXAa37yI0v+iqLkG8rW1ENg
R2Fu6Q5yBV4jRp8nkdtWQkmLzEEhPEyzcr9huTYE/qRq2WjZjKd+srLk83DipPTX
LL1L1IU44au4eHhSKzwsmWYnP7g+6uLRL4t6TvaIEdMzJ/g97phc+u13gJzrLaS3
1D+Ikio2gzziLWD9/jklZOAyOdp2n2+8O2nuIpXZOrlzFCZxsm9ywt98RKqN3Q1I
5Gx6x1AJR6Qzq2k+uA3VwLAMpi9vxF/doc1Ht5JtAXR4UlXXh9z8nM4liSUm3an8
O6A2DmYrVir0VCGPwWHagRoUwKNgl2BULYMa16+w09t3JULuAXzQPbosXnpjVjIF
Xeb18T1E1VDMdRa13HLTRhAvgt/fs9pi7TZruroNz6TpgbKIFXdD/4swUiWK6i85
yen7F3n1OZfS9X7FJVc6Ftfjy+n6kegrMn5I06OHV2492Ajhk7XZ3SEAf77Lwy5c
/NEYbapeSyhuhwD/fxrRAHAj87Gcqi2utazXqL2en9VMVInnzLYUAdQDFuPzbMqe
oasKqoK3I6dKLcpRxdPABsIh0uvym0Lv9Glp61g0eruAVG7NPEPldz7E6/TaCgW+
RF0zS05uqLmQtalo5JqWFHO5ryV0qvZdr+OGmQMvlh+N6NYdpMNqQMcwwumeXNTb
1NnA2oE+WTQ9B7c1Y3xelQJJFaFHB787yF4TYfMljXOLetcNMltAVB1iz5uOiMnC
gZVoW2iIlMUwskJUVv30sjzCoCDxP4CwLfqvaR4m+4mgqx4+GmNgUgi3L//HXxUY
pVRfZRNJRI5Isks1/OsG2EEIE26OsAnWOBUm2D/2la7pUQ9yuMqLbUreHaVPdMlb
naKMhTHRFS93P68VZotFIFGUNcHf1NGItIq/jXUzvhZ9eac3H0xMEHc6tNrQ6KA5
AXAzuoJV62dTEGfi/iDQIG+7uhCdBgf+08hQcNIvNqm/N5iw6CZJEjDWFPGaZdKr
yL1SNka0BQWEDeIka+mcMiL1tvVFdnLC3B6hBINcXqLVyL5HWx+yrvfCnkSzOqFG
y0eiakCUIjLetmwwR2kJlV47LdXwqJAFrAq6BJX6EEXB1incbt1wknTYI8SIg3zR
QeaS5OeKrV/QpGPRsfJwcRrSd9vg5EJTfs/q44JJ9QIp1D88aCZqNPqpqefchVKu
G7EcmUPkBy9qoturNUtmL+D7uHYOZne8jpbD1AZElrCLkvbBtYxPH9B5S9A1o2W9
RyeP7gbmGGIsA194vA+NjY896l3DfkMxjl2Y+PVASznx0EhufHI7eCXF/vXO9F0G
8xIoaIsnQcZSUKj4c+bhrUiE3CBql/EEd6Rq5xWlO7javo/wdrIPJBAaQHy2BHeY
dh0MmmTgRdQKB0lzg0XxsT36HUmv4eE7C9JToYIkMvwYsmE6spcAkDysG2ZB5F2C
Xkfa3C1Y5LbJozvHkxhL9mEgOCvh70Z87Zfso+WxQ5CP9y4yOSQK1ONEDX5Bj+o6
5Kj6Uqg53sfY+ZeHHWvv0iNs4UeMh4A58DJJnCVBvn9+v56Egx2Zc/M5BW5dGHhS
eRQLtXy9Op52nqn8wcZS84HGRzZm4eg6QaL1VLO35nJBDSS70gI9m9iLzW5l7Oa/
kfj9Jl8g/9HrP17ceKhD0+yZi0cvYTT6DZDE9xIxV5NceTwknG3csYs/HpB7mbhn
gh6+oCqzbSMdeRGgUITQ40Zc9o1JykrbrNDxt6Ux7QegwkK5+eCBwgstcGN8Tx3O
kVWd6CGIRz3cjurBaYMi4ivGy+hI3/Bkk7cAhLpVCkiEPn+m5Yo6GcfLy1VjAnHW
1XgsqMOupxLd2nfw/8AJa9mO3QOz5TtB4jFsIAU4knJjIFMT/I2chLrOqLwNuODb
+EapUTiJavAVyaBxdmK/m83ZSlZCeJpbLsz6zaTDVDVeyK7Xfk+Y1NPu+4ZbZTaW
2zv3DyU/QoCCm26M3uR5MBTrSLouvbxP1fhiQEwj96nzkOJB4awiSHiC3YNeZrIG
TH7MmavNjabPm1dmKYmYRbja1oq47NkGl/k/SIfrZdt04/2RxSwB63PKWNzSxk/Z
ADd3cRNnhhRxrI5YWLoB5yMl5NQ4trT/wucPt3Ym5qBY1k2dEsoKWDvNts46RXvp
ddyFPXCThKBqZ9on45XrtZEuKYQqOQ/dCfRxRMbyN3SJNG7uxI7KcVujkCl7efwT
uCQyYCQsepqotB9X5K2dH+yG+2ES/uZxDpjRJozqQiUuHq2Fune/kmPkJLwIRl5l
ntAvlsLmML58ZZRq28dxPSDYg5X4FJztPX/4mrJRlYgslse/8zRibC2AD3n4LAG5
HY2mlOsJWPUOQjwg0YR3978poxfOxfaHF4MzJaizkiJKDMradDTkO323aw6cjnYh
aWFqBGPYZuOyKbA+O3TC8tUOjTWYbnEvhOPZJpbYZaD2LDIOQcKjR1eak6xeCNXY
H8Jl2LKwcS4cd+FKbIxG2t6bBcvfR4oqVkRaBcoNbLa7aNiQj6svv9hnlz2SPztK
WiOhVDTe+Z5TxgBCcbWg903WArQqGXLAlhAWSfc/eUke6qH5D9jhPkCUkgdHsHfn
fLRQDLic1g0RRNmlCc25kKk80KGbGqWuDvnhDeStNSbG3U4f0exj2QFOafB8bdf1
XGEuu0ijHUZcecFOaH2gUavT0FRbxFG2AD6wO8jROYRR3jykj1kfmC1+vqorGCrP
8H1autv0x7gSL3QBK9oUgxOKneJnQwLJrr6NwnB4zLuL4L/h1FaM9WJHATvwrBGt
dUkxCug7m0TctSi7XhoIQ6nstMGTSB036e59UziSIftb8oSEap8PsmuEo7kYPccu
Q/go8WicPRg6wafV9ywb3yOADpqY8QgyOUuAJjooRgBTPPqPZjjVb3iIncOa3Ry7
V1p+vDCEyplzHW/FHAgxvvtCa5c7cI0TKfjQ3PLoQ55ZBbmz469WLX8bFIeC7Ndo
7C2mDsWFHF2EE3+VCzNFcGFY49nQujbuqT+hRWiSOJcMaA774gZq59PbYrgeF8+z
4hXLVC/zxycYdoBU08zumWSk0EBN1ojOmRKTJeXtFDVR0R4+ixdgZaSdPHYqfCxU
cs5/i+HASBijNba5WckK9v869djTNZGNPSS9Tbo88BRNGqZ3VHvgrSL8uqDuOKAD
QlQY49M0gjdHVRm97xrYk/QizBnjwO9JBhdiVem6fqAg2GOaSSdLSDi9qKKO1ys8
VeNSA7sr1Veq7RMdLnw4peieAx4pQj1oBgvUYwaoTRM0QktzG46gmCeX8kq7ZAwL
leRbhCOb+N0i0Dt+czC3KUD/XVUBwy86kRVZ7Fb7XXrM0rE6rRNmDDsIkbyBBnhZ
JhP+KYDFMX0ORMmQGxlyYGFkVF1OW1uq8NehMatTnnZLolcnbqGwFrD95peStxSS
QZSozWUddMP+1kaf/SbRLWtYNHBFudjuMhJfmAUVptVb2vofnQUIno1leVCzqIY4
ztNO8eq0Y3tZKbOA9ovum1CcK8iuXavbR/bKWe/YuZ0TAfVOc1Aesq/ki0dN9q+t
UU/aG1gy+E+SgIz1rddNuArs0etFv948ZxtqfwVQ0t6Ur75CXbQw37DvnC+PgfE0
MMpEbBTXszwkLyU8imWS1bimjS//JqCL6XSReuSQFb0D+01wslxJJIJcN99fUTL5
9rja5HXSv+NfJgcUBr0GAKGCMk9yFj4Vmj+5bySyLtKgyRDswcg2juALt2TQ6Hd9
j1pd46ynWBfu7UwOdWp3ELwyH1Hi6m5+87xjTDAZ0LlvUpIYqp4MUqQzTqx0Ocle
4j/HXS+VfyF1Wsk9vX93ObDoLsU8V735WDy9onDDc4YFe+GGeRdcWroC65r6dvmK
YVPOz+aPj/8ANrAoDDQEOsnUlvVmaDPGTHDuKcj7/QKmD9gKFEwdJ88BF2EUYUrI
YLhPuQozqsizf0PXUcBegNy+y6nWKEug69e3WNNiG+yhwwYvpLlOmZah1Yfy2bxy
ogTLG6DURCw8JNBHVGYi8HOsmyFdAnucmmNQxwyiY2wEwGJNyX94zCC/M1MXh1IY
Y5i0v2rwnPjS98bJehuVVoxJckGFcG28nQtNq7JnNR2vzXNGo/8QopBL41mpLMf1
1FP+Hs8DjJUKdNnhzBCyvC5LQO2sCwFNgxDZBOcdLhZkcwf+eDcxWhBn/Ypk9Jfc
obwt6dn+N7B1vPVs1UqPh2+p/Le8j17ey820Ds0W75gNIIihl3XdkFIuTE1D4rbe
kehMYYOQ3kpadfDLV42vg8eZ34b8HssagL1FU13qMxPTrz6XxwRrrvBrZ3UhYZEI
8JjHfoADEgtAkS6um0k/8+Hn1yuiDoyjgqyJ5BDMUVd4DzYzwFcBf+EctZFM9Jj9
eD0pqPb9y5SJqAFLdZalxO+zLZk0BVl5G0mItHyIFaBqPPtcLlTKDnRd5WKYY7kQ
Rz3oQ+DPzusfsQUHXL0RRjuyJOBOysNBW/4x7GcCY8smdOiaYomaEehXuRDJczdy
ql6gFz1EPgAZCmE+MZKS5GWmuKJQFKDNW08ZTFo9cE0IczmumARiBIAc+bwJ7gsI
jt8HFlN+2j7Wwwk3b4nijWGqOEPjHQcZEGHczmGyvHMKU4FmZ/s7zHVT+PJn0MaC
5S32qmoKRP00yaUofKx2blNb586X/r8FqqlXI+67XzYFRWktcX59fjp0K4Xm4EmL
vUmSU0utVoUT3xLm6A0iinKWUBkW+fyPv2RbEimFsfEQi31M+1n2Jr2UH36WnfuO
UtVata6mF3wiAdV5WcGee/EfAEnJGWHPgZs78ZXK++0APvofF5n168bmaxaS9oG8
+87RqukmtgTVnecBmWkdD7k7626aZtReZN3O40J0wbaHUpbdd//t2KicELm5gTTh
sHXYeFc3wgzhLYonKW8O90+ozVIkzN++ivZj4+DirDDwzPkVr3sV35WDzlLO8/ka
R85stf/ygJS98jYk3cS7LEEWrtoXGaRwRYB2wxRcOzRVvIwluve3IcISAltAPozf
WZcjWgJzUtcR2VcCf6kZv8SJr7qr3RSGcWRJR9XxnM0BJ6hbBQ6Euu82VZ4c//i9
s40nNy2ZKdPncx62oBJbjNjcvZtyCrCzZBPpgmybwT/64LKDACjNcX7lLNU79ncL
Zbf8cF5Coi9uZPu7/gtd6eIFhEkEsoB3e8SbFdjo5pcu/MH7pTAXwWWB6SMOYxY9
A1+FQbdsmpdVvcUVhbf56CZFXGsTjHqL6ZD9oRL+9EMaWVlqrdktz9kNgEOhWecW
jqqpaN23V1r7mXovG/En424iH4Pyfbc8uMRfwkcR8Ghzy7PwQJI37bO2fTry+PN5
d/aIwv33OBW0HYvfEGT3YPbdN2bkvfXkdj1p4SA40GPaZ0hWI84SxsiVrgTsf5Sd
QlN+8OY2RR0nLjQV3p2mmiejcRrlJdU7IF4bRMPl0jdnm1HZnRaOHByr65JIi1Kd
ADbR5pP5/unPfdNRiMrKvi3njJTZeQx9FsPW3MoUIFanwthVPwihL7s+YUznT6V4
BXxj385DW379d97STxVNg+v06PLOSEVNgQ2MOQxvh7A3fpWags3y+dMyZ69ZcwPn
RRe6V7JGCcAbDtxhOlJAiJP6DxovC0dEkX3FRJItQTl2uJtbBBQefpyc7nRFqT67
1aeI3ap1ObJkB3nqDeEBiLgm1Pwvu9iUdDOg3fhx8YLdYD6nazn7SfcTB+AJt+ll
oHMutYTU5VUvJcgup8NPP0h5iu6WEASd3aJkwveu4NTBGXp+Ob68LbbWfen5Q6yE
MsKefyPJx0YapctvJ5iWu4BAO10w61dTK0tXm7xHpqFygfMGZPsDKyJNpLfsoPNh
cv82zyE2WySLZ9IInfZnQHGZ5w7glDO+0HVmG3b3aRK7kQ/cR0Fj/+ubpaAWgj96
o1QgZ+ua3mHCkzJ9Q9PwceItLf1mE0+Fuw7460b6jTQLcnZ2V/uvJ7ql2te8C+Kc
WszKCNJBTVi9cEXShCFL25b2YOQrROpGSWIaHT2LpmI2+/GOvl66xLA/taDKqm/U
Nl2mAh1xtQFbGH9DFzu/N76J2UwNL5gctk1N4n3d+sDkHU40mnp3FH1fpK03XN+k
5lCqWuV3ewqZ/rhY+r57m/9hu9epafmywBjFIcs79Bmwv4DWQ7CMinu1+hiREU48
oSXYIehYiWM77ttsxdzhrzDElMHnTAfoHEminnwRDTiqx9e9ybYoqEGOXWq9u+A3
dUbQi4fFsaxl6E3BOikH81UxLjLsF8xQatfdoaQnMd5OWP5qp3Hy7WEnXfr32B95
FnCGkXjpgijC52I/dlayTF4INBG1oD9QOB1A6iqXsy90QrkM1+8qpNtWU4siKzvH
xOTRWDghwFXxSWp890mT8o19gROOUdreuQWEoeRGmNSjpswMsLcMzgFQfq/eLMH/
JRKmAH9tAaoIeRpUxBmuVkJCg4i0iby/mdWHV5NdpRd6vW0PkIhSLiC7VrTY1rfi
ziN+5uySAp0r/ACNHAJTHrFXgOFWJmU2JZATNLz4q5LsYCx02uB5I1rW7Xm2DWWk
dlI4HJPmftS9MIfiLBlpshgbRRxSHTo7DMwYau3Y23nRYtWJqAr3UziTRrHHPMnG
XmJYUfwbCZkfUVrFBmD+xTJOUXPJkAwpneC6a00SmneLoBqEC1N309axti3RFRjz
qYTxHrXvWJdDKHO8hLDDV9qy2r3S8ZTUtDnlLhmCfYZdfkmNHdjDWjSd5Mgt/AXv
T0A3296yeQFPDKaZQniC3VxAu8vd4yMko6h5Cnhj6vWpexFH5nikA7siEmBi6jhR
uoty3KY84fVGOwj/EiB1LKJpHd0Za12+wmQhP9cwPylUVxCO1yPv48Kh2FbJuK0S
TBtEOTnPLyts/9/Zlep1JHKJApR8ICRqAh6ipN6DcHXx09rBKLMTvV9Ohfjongv/
Wt/aLuwsamn06FDrHiLIIbVGly7BL9eNvjg9vBaH8afsP8w0jsnFVxGQKEdQT0vD
sb/CiMWhfJ5Y0i/AkEWrVR4nIqb6wwa9Ll9O3EsxYCkCONljI12okmSxanTr371d
Hux0s5MY/3PAgSY9TZSTOmqjB6kRncDIaDGAhX8yRU8wFD6KeUoBDdGOeTk4W6Jf
+CgXMRtt9LfFItnZSJmt5HrPTQ29I8e3yI2y3H8hJfn0xFiMgvj+1GUrczVajL8a
RYz/STrFOgDxDh7nmDdQzO0PuTe+ftQfaZ41Pt9YY3tOLjc+uFSLu6C3swewPk5y
iYbtFbhfT41yCHzVHJ9sn8VOiP/xKyT/Z2xjxveQdA5cqIqYk221laXX9B7wQeWJ
y4JlDtlzrLWGTwVqubD3ELWjrO4qeHiNvByD448WxWtrbTpW0L/MJZwSUn3jyZt1
Sg/hC3q68nV362itELmThOEfLzTk6T0GE3sWtXBRGb7B6saIO0p3srLVVgPfR8GN
hIpAZQW5/mp0WY46kFXB2gucLi8KP2MGGvmM2xDBl+XfybneOMOsiIAwOXjSIU1i
hiFIF0pG0vQzpaRhDRN7o0gi7Uzb700wAM/t8yQYjyRy3igntILc9d61FUs9MVhM
TkqitPsH1xfMvk+55Fk6+f8lCuFxU7ftKg8UCrYnh/5s0KdYBY/vpABd6Vb1ez/1
mDFCZTKhBcZPoCOOhwzIh/Tt/h+MfReJL3+OUhcjXbVgHunpWCvUXVYYxudtfv9v
4Zmd4EntseGenOwKdLd3b5iHht/0K3iqVAFCO7L3db30E1nNJ0HBjP6nW7J1xwcE
MDC5FncePtY12ZtbxPGwA3H+3ro3lvzagBrbe8KMzqMp0PmnHp7eRj9WiTgEnL/R
UGKWAlwdy/WlR39mYsHMTdOQokypTYn2Hhz5wNjZHWt1CP+goJphCPIu+sSiISSg
NbBKJVmngGxRMLmHAReeywAx3JNoeE/SH6Tx5y57W0A1xZxuxplXNU/O3N8xoav6
lk+d95+Pd48tD08UnWJNP+Z8AHzJlxNVxjnPa966y74zCpn+sQwOQ+BVLrKaiwzT
f7wIJptfIPJeTcT80HW8CMyOUnQ4xTRlh6F/VP9oomTFqefu0A4CIIGtxxztHM8k
X7m8Ewp0ffR4YJokIrgwvTprs1pdTRJ22X7uK9LHHtRCMdWMHyOqaFtfaHb8Xz3i
dMUt8xBvWovHCc2lUL+M7Z1ppI1+5RXRMRsYbR2DzFao9cm+ySsgtKSNYTvotXka
OE9AJNRJX7f98l+b5iGfS3fFQOge0AClW9+1luMRGJDVPc0hivBKnWQ+jaQ+omlJ
zFWy3/G0O+9LlXmpvk6AgxHs1aB7VVkhgIenATFRCjNC4g8EoRjZGL63rnzF/KJt
UinpIbkxhOHK7NslQC4tHDErPrQLn/GQeSDhCbDJ0l6UnoWLZ0kifm6MNXv6Nw9y
VNrCwHyep9CzZvDLRLsv6yrt1tpS0H2NOGGJPy97kUzzVUMo8dF/BLOZm6L+aRnt
YqbVsI5JLEwTo71DtxzE7Ea8X0Kd1k4xvVloT+WrhRHPh8UwqfkbJ3D7mzgs2bmA
c6DuEb7XTQrWTisF2/h33XTaqZ1aSOT7GXODJqDnB18eD4oglAOzAU/b8NmD9zoV
4b0/9GT8BkOayxOep5pwQy+8rMsZxZBdDLxHW537xBN/CaP77CfDIfl5n8kuWP7s
yW+bxt0f2QQDIJCylgyCX9qRSK7ONfVy/GDKUvjfV+v4qyPQLw+ExhRn8EOHZgny
Skfj4i+IuJdzYz+YyLeqbRBuTOYavoF53LiJNHg/V0UcSLMvoW0pO3XjAHxV6IyM
XFf3hQdw/hMLc9tKbzIp9cx78RXwzvZVCKfR97HGNhLNlXrsZtTnm3pcBGAf8Pdb
Gc2jSewmN6RnbUeWOsdsYueW+yxRRbX7UJu9gwkYIdShYodAWfzS+QJvdAit5tHg
UPFhewn2dIyQBNnGj+S/TdaC/uDmhC8XeXYQIoWcio1SISliVwwbagtHinxXKIdd
/8AZ5woGDOPXuzR8uFuvXsX6EG76XYz0gWTMHjruGe4IuUPb50dljvSIFJwcKa5T
3JUZthZYaxjGvqQzFNARgFW38tuNlC5zkigDcvHZWIWRVlX0MmZFCEl7zi3Cjz7D
aP4Wir8SUQc4nRFIuMHHafZhp2cUMGF+a19hE+KWlihrxPvvwVnvwwynj7ZlT/uE
CfARh2MK1UXO0y0XFa5+qsKchtHwfqzcy0O/cpD1x4gjHYYr7upnhU8TvwndDS3l
S5RarNa4Eoqsc10fanIbAzbZTdE6PN/JGKINLLZFLwP8hvIgdPXdJL0NXcejy/Xk
+UPA4Yek4uE0d82jy/Sc5WXMpUIt1itpSwJKkQrcUjUp5PSaagePOUx4nyxPG4wV
mQYUFTCSKRlLUsE+f2oOZSzC195AxpoORyGkPHxpDLmB1FWlN0dkKkS3wA8dNHkY
3yhB3MIn/fYqnjmpu7LejsRzZQbqJnzhz2x2ITU23r2gOzEP+Rr6Drsn4fhNqx8C
sR75pX78DBnzrwn0Q1xyjdn5Cky7ZlhJkqDC9aAxosvcmjX9fRYIc15nYz0Q1NyQ
w/vz5Pn0+pRE1nAt8bnXtLyEc73oiqzHIm0+B+Tyjc73H+MA+GTkT3q1bqRwT9X9
Ttz14Dmn5OdRthTzvKltBrgIOdzIkYwsfx/PNhanwjQ+pvrCluWlTzrtdgLqqPEs
9vFE8szo8igRk6oBtxroKge+gihfeqa8sHZgrabAlX7/fTG2pB1U61YzaYljJC3O
2GsYxUp2SES062651+M3lL1yfg10llCRFvOsDq8o+A9C4f7jJ7oFjsb9GdbYd1AL
K3GKFhy2b3TTjwxYIKnZqLYnXsvg397aEmwYAZOFNeOZLWdHMPLBjX5lX/D2CZsP
Wq/EskvFWlxr/XKarPVfs6qmffebXRHgVO6vToZydcAgl3tLkOjZwSuHiqip6tZF
q3baBhv3XstDNayrhJNiCFx3GUAjBFTDqwrlzCOH9zDDNhTOAQQaK/afZ0qJaIT+
Bxw+/dC9a8LCFzA9UsrwWSnRV7gs1O0i/1jisp0a1sju4gklpFTbg0dxCmp4xDWt
cSTL0OaInhGd6K3F+SbfWUSivMNPOVBP7YivKwYLZaSAB9yQwd0FEnbNPe5512Ep
fq1NlDat1p5rCYPMiRNYp/tTNXHXCSbJZ3Pzj3eqXFMdRkRFZl51hH15Wn4w2QPa
dDKfm+AHqfFrXX6QKpyVI7G98o9esGrX1Q+ewgvvIbRnqilJX5kUKtwk7v1hMNQN
cpMqGKLQKanvH3hfLcH4e2Vy0PnGjaADmddU1m9FTjDQS1+568Z0o0COBAk1MGDl
ztDUysS94MTnSRMsDopR12+dxXLLk9X6bPBUuVBk0J8T40TTd/6m18V5snMNyjs+
HpNHTHy2QIPJVy6Xviho0A5Bhf4BlJgN+j0r+uCc+PzUbGVql1GObEg0XI8a+r8I
e+dUITply1wQyjw6NoFiONYHVBcSB6d6GiWH0gziVkoKHs2wP95+zH+fPkJN3V2R
YiiMH1E+KbjY42kKBRsFTScXT6+y+s8RizUMLfJ+NRKPkQyw5YZ/7isqbDcqNB4y
YnmzpfS57vBA2ZbbcJvU+o42uQ0cjVIl3xeS0NwkX+s3yVzk97c86LzajXd6AcRG
CUgZpKRFZJGE7uQAo+8/b5V30w4ix8xlFUX6yEaeM3KgxthyVhr7esklugMEoYcr
1KjoAPXlNH/vNTsAp0f7J2cuZHFqAHjVkbdxjXSvWVRGE6AOUro4sx/yPx5DKzNt
pX+Qzd6mqoU06aAJwimBO+JcvmzGL+hd/E1Y/sGc6IFtKI/5zDfqdtvGkeIlYroG
gPEw2eMIl05m4EpUsgPptSvHYNrgLqseNuDMHWlg29HOT9joI/VMcDlvRis8YO+x
I6pUXhNGkX7KBGaz4DicR36TTrOV6dA1k8dAtIDYTPjnnhULEyVMg2DvlEvemC52
LfM5QUVENuzfimFSPh/NGbfIkbAux4v4+qkzf8fXHogbJeCinwrPdGRrCIuPAeQp
f+HlWmg2HY/vYUGqicp4txQR1e2SPyq32K5eUcQSHFguCdTerpdlb2iCyrAVKofn
0eg7sgCNCthXIiqP1M+zDfhhBRhzcnfDZvuSr4BJK5u2f8hMOAYnLTcrjNH8yMP4
CRbf1hG6sxNIWThB46SjU89S34jr8kf9VwRq0WRV72bKY7j92rJNFoyMcDnRp9Rv
Elmg1/TbUCLAjrl1rZa7pGaV8XJnkGFB5fuJkjIA2SsUOKInFwD0WoQPxnamumgV
SD5PKu5RbRPJ9go/hjp33qW7VMBzMIpVDupZA+2Qtv0YuQx9QUkyVpEmjiI05oki
yzetpz8InbbXdCIU65BAwEs8ouHEI2VaAEcK5onoPU2SMt5o4XsM0kOs00cIDMrb
1FLX+lSI5pTA+SMe8tWP0qOjOax5S4C8Drf1vzEEBlrM9TQUOQ3mbwy79hOG7xoT
0ydbNH1EDN5PDoy6LzoCrZ+RdD4LphwNHg3AJK41siuNLGqrNDd/KB+kuveL9rr1
67BoQ0NfqFjcCxas6hdwEUW/Dr6LmlfLzFQJd7IIfypXLWYDv/EmWMgj0dcit/BD
4gDgWzl3WkMvsheHKnUam6oPmrXN3RiwKnOzTFlvSWdF7YVTlJqx0SMoBF/ZjDc7
iUClC2yf7Ytitwb37Zyv/XUHHdkwS/fPlhUKmPxrPS6kBW0r2vYnBjOyk5ANI5eI
SPn8Rf7S1XK3vm2ED/RYGfNkWmtfvP9Q1zccvvqGr8tzgehYqrxilPLDb6pelEz3
TC1TLsjPoTGFndc5l6Wxzerun+C4sW5XK0kw7bsS0/+7UtP3GXPbnCPUWpRQdPBA
9uU/5EfvAzIOJ4f12XKOVJVreCVpPgGCZenckZcgZ5+3V1/4MyUoa6Co36CDMVT+
jw/20pqsfxhSUIwLeAsSA/o1SOhxcl/l0Wk0plCRwyPzfL0JUQLuUmmldPmAQ3ea
LKum2JyvjKSZtdrd5RHfnlDt8YRlKJqO1usZLe9yF5Tlrcfjzx4HrGf0UUCYteyb
zQBsHZDX5y0pZgQbpF3rvF45HF+BHFfTRNWDKdrbIC4v+jU5zafdYmCnzc0cipxR
sMmPzAu1RkudnCOF7ixAc8E4RZhyStbXgkw9yBcVf/DyhwTnYpMS7EIDVLJ+hYOr
7/WcV6HccraqPnuep/OlpDbpvlSoIjPAEpDbhC296F4T9NIVhw5haqjw7ATuaMJW
CNLiXn1MfwldWTwU3fHQXKIsX9xLznLaYbKsCdb6ajLpDszLfGr+EYW24QYPUZ72
l0t4FTJIEG+HKz3JARl915WrYeiF73tSQx/sosl14GJ5fWqwpJq3kAh8uMdDnWFS
G4VdcAq+/5sgYy6Kq1Edb4lurjN4QXOvldRD7zDiuyrsrXVvOEVenilCshTo+T8r
cmAkhgVn2atgUW62ReoROlvwkvgtUDjqHdrFIxtvKDGeuWrF95rHEQRoSFeJmG8l
3QT95lBFF2hx+Ryx3erNZP5EekfitSIKzQMKSpHf0x/YpUwpX6mzvUyzwK3/1+4n
FtMgug0dFGPeMBUvTO/nQu8ohB+JkJRjpCnieP79IxsrLMgOXTJcOlAU0Rp2FHiB
SXgieXLW9VAw4uMLvLHkcStSUnv7b1ZG9ZY4IsfF132z+emSalF66XkWookqHtRH
S5cw0ZuME4Awvk6FM2PMZda0GkGTkMOFLHmzespumA/drLHoWGLYJIHyKlcq4S7a
HN7LXlqKSomLxD2aWkE5pdbk4cnE8aarqgJuSfMVwN+A4JvbyV1T0DIVUzs5CbOp
kKlB1adjRvUcW8CmdkN5VzdR0JTfzONhU2HjTb5DkEI6UXQoZIA7O2MUmVzt6lZx
d5kEp3uoszy/yCbIyJ+D29oV0AScJmU/qwEPYAYSZCXlT2WsIT41DDdr/YjvN0cm
vjkt1NFahy19avmPsrQ6dR06311mbuEUltHG5vlSXEPClug+dabS7AFTMIEE3wGx
4naZP6/4RShKqBm6t+nu72m5547mAMkwAfxq2Q2zzNtCNTPFAiK6yNC0mEdspa0Y
b2PQJcz/JmawrNNYztqqQxjJvdctUa+f95oVFJNxnN4OgDUcsrVB5vLOLGL455w0
Syv7DS6xkdSrrULTCilXJ2tPijx7yXxsCq+ZNi3iioYbAU40ts4zIQCzqz6DosKy
AP1eRPgMs9Pxvzo4HyjoLv16NW4tBU8YwbLMA+Qurdv+Hly2AgkWLhV0w0/Uc9vd
D1OFW/wRUwZ/FclwKF4DTKu2eL85bEaqjZlMISLQXdrmBB0yRBCJ8FkUjyJ73NCt
MXCQ6XoxSj9pf+iQr5OudN8KtZtyssRaiXXPEOv0SORLHbNqKkndaRXBmxsxOjUK
4qi2eJnjPAlp+wK8FGNid2I907iic84Nz0HBvCjDH0W8Y0lCVYlzj3A1GeGqsuXO
GUzH/8DZfiZwGOxTmpV+miI4kHChnOU9PIYvPQE17MP8BM+ldZauDZJlyvbfHuYc
Lohp++D1YXO+UmrYn7eATJIEuJs9jyy3ZqrViV+qMIydpyWqW1caloEb3eoGRFNP
49FqA5cmUW1mnxwIFsr+9FjyoKSWj+r98d6mx2yyAKl3xisSkgWbkdNqivAFZZJB
bXap+dQ0nMC8SqvqVcl3cUQhyo2Ob3xk/tZFeEWWdxhd+Mj0M5o3wFs1ViyZyIU6
RJwm+1I+vqRrmWWbXuqpZjUAQdp5pCB49Gt96C26R0nm5RvUA5gFDnvhdrlhtBRj
FCAkVf9w4qreov/YJAEiefoGPpVQEwggGOHGlIxJ7Hf2udNde7PqhGkhvngdXjNX
VCP772okUGCd17bpip7eGu/VRFcB469pSXOcHxFd4uld+YzU/Rakq7Ike9w1F7U7
LzUYMnpOiA9KL9BChlPCLXEbdLIJMYFxr2Ob5AYrVdhv4p86t+HQww8cvQPNUPae
W2ngICBds2cbMij5qr3dSqEJ7aq4d1TLC0lWc9fj399Dz2zr0Lh+edHKhbC4vOT3
Vo5tqFwpKnZxsvYXUQIiftc1wwjF/9XTjH/dTwTokDiMT3qC3LPrtOi7F5VaRjkS
5otaAyTNg7LcEQ5uTAcHW4PSlBftRH68PkGvtZx5WjPMYqmhynPbMl5nN9kjWEEk
/niwIxJ86aNTcT5/ms3OXLW3r+a0vEWlw0/4maCtd7bCD9VlmFvozVMdPF8rRhuq
iaFudz9fyXlPbRD2HqxtMOSUMSIgRevLfnOqF/C81Y4Tdk6IhsTOhD26H7Gpt25g
IaePwasQAj+jV/wtJdPxFdFenhtrP5soHgTgCU6Z6iLhXJl4lDsjduKn+UcaaBji
FKRFefzzXsOs3mOgVMFFeB1GZyh30Bi0stXslg6/CXakkONntuGO1CF9Hz7knXFx
vjfs5OpJCpMYwDt8BCUKPQ+4TWHZIkki0HceiuhE0SF8KGUEIpvZTM9RR2tD/8oI
gweVlp68GCUyPIjDH5871qlEM2BHlSLU6fnAjJ0eRFAlTAyJZ/klV9mpZef+1z7j
YE/haxlagKboRfB5QF+wLJFm60lhqZGqK9WeyFxTRUaJ7TBXoyJ3NzcfDDAl6hMb
SKBR3lBp89w7gFIPKFzUi7Ao0dJ0vspkvfFZilfsX5S4kY1qMPBZ3qDewHuSrAMb
I1Z0ZThyylVeo8NnWK7DvEIA+Kl/AfS/L48x5pdmVnq3H3Uf5WtFvQ2JOhF8GwRy
VsTaA0mnOc9IGjNMxEV07iZxwMGLF4ZksSM87n4PQJQK/1OjDguhBbW7ClK2Itmc
ow6/wJBeN5SeR3HyNNhArAOcmE0DKHmP1D7BQJ76KDcNNCwV1F72sk4tj9Jgxpqp
0MYeNkUoX0gvLZraad2FiXTfdAZsz2OJPNsnAbRnhYi8ick+GEXK+KsmG7Gf0+0T
2fBCxWn48jQIbJTTL2ACU9IAL1O0Kmzc/bYqf3/nPkUmDLpFQ+02xX5N3YpvrvoA
/jMCoat/v422u7n/mroEFhPhRlZghVABWYDHahCq3S+2c6wL19frQ7SJj1lodW/t
IorMnGWBlF9Ar7VI3phxJX4HPwRH+i+GFypqVLnpMYyZaKlGffMRZ3HhxY64zKSB
1txRg02uk+9JNQmpbzHHyLGd2BvTk1BhgL6eDgjA/xcOEvXZxjyss11nZwjtcS5U
nQwweDsCUn2QXq5pMOYoKQx4O71bhlyXIp6DEFi0h8WsgnVo0v8+WQPfquXh0nZP
q6mzo6SzFwtL7A1QpcBmEaBv5ygA/Fb838iwAN+GzdR7Pnt79xSYQEW9TRWwSjsI
GwQK1TLc4iX3GJNXWsiDIBM6HMIVMxJl59Ng/f9uNAuuEPn/iLIvf+T2KWy0iobA
qXrMZYIZWqcQUat8mbG347d8H/YF0YuJ/GypPXhHjz3n5wYFyi/QZ0SzfWAv6BMm
XRMgcM3gXse8/Y0IhMQZHwqLWIsVsSFxTeESRiBGEbLFNrf56I6fWiBcUTJL8tZM
xNvFT6cv05vX6arO3nYdxXspxKkcpJ7/goc/QfiX2lWL04rfl88vc6Y8gqJSKI+X
aFwU6Kq8f1NY7OfgFkElLrws1JLfJYF2g4Fbshs3xpxDMVSxAuTL5JD7OVTdJIzG
FHiVSPuTPlaXRd8vPaooke81ENm5cKQSn5JMjbXO4d+3LAlaRNymatVoWKqOnu9e
ZsJc0xmnisP45IgRPkODtobcxj0f6n+ycjY5gv5ul4Zehsl4ikyI45onAlFgvkL7
YG6oHzqzqADQ9zQmt1rm0VZwOYSSbEFpEnSzPno6Wmgum8ym+WXDOti1lI7UkBjM
ozf8TmmbyKfQETBXRaBY00zAAH6FFPCl87F6c/0L/MwM+1q5ZaCXW+l5/xOLk2FR
1OC3k6216ERjnuPtrBggZRqCksXJ20Lin5gefAjQ5sbVdPn42nsKUdcab4TFSCdp
4oI9giAVPP3bzU62Y+EUnFTnFn0EZaxJcbbiy+j3HbnNTFWooY/3vkZg6bsjGP2G
G4dt5H/gtp9D2wZWJjcOzTE8C2td5JJ+nLeJaWAp8Ye0zGm+QT3IfLKXGAuYmOCv
1ZHicN3cewZcDv/SWRklj5A/PbGaSSgxoaVF5kjmZjtH+ZTQ9qvvzYAWdKJN7UUh
Q1gDny196yS+/VStfVuz7LUsXDrs63cmIq0OZCZHUa5DrnVeVMwSu+jXqRqKNKHO
uXagKBmxHQV/SHebE2yLIIuNFm3d/asM/Nc+c97NuBoDnkDLgQFiCr/52z412/qI
/pOEJi6dOVxtsDr1j4/3nxNNZvhlgBSGy897xSeEE2RgheCPjNGAgG1IVtpdV9AY
D1M/PqfcpBY+yEHyh7Z523R2JgBxJzklWPmfudiojgamzTNU/DSVh1mf4WpNouR9
M2hvInQQPKKfToex0Jb9S4gTAwgcBp7edZK8It1mk/3CXJvlvGRc6uLeL/PEq6CP
xi2T1HVWYd/lDCxdewQJX74cr7jqchvFHbc30TIWDCkwWh3id7QKJz6J7vYnMVzq
O577M4EOqNDLm9VwMn6UV7xFBh+DPMlYbNALVd2nrketijXgAiIEKURUx3kJv4la
jSRvW0LX4o698B4JjAwKacfcMdY4wYaSILYwsrq+pAfoFo6n3KqQ82u+jokwSJQ5
BTaUSPwtxul8cxCuJx0O8OpvUBAzLSWEwDUDo05NfBTKrnKPMUSXgD5HcuEEw+Dw
TF7x2p114xrnf3t6JimEoW+r0sdTfqa0R5CQURTNYc9yGK/hWts3QFYEjKTOIxhV
QnFK0nDriLevE3JTL19QrQNPMzek4ZzO2M5WCNYgOgqMmKEhP1awF32xfJlXyMfL
zC1nSkVCmxBcaJ1DqwtsljJUxFvKt9URaloJ77lGR1+hHVD6Z7c2LVqnwEZRJg7t
4gMQpXYFVimIf0OZollG3kjMA0U10KPyBRywiXtFcr9Ru/ChZCF/mQQBRCyNwxRx
SJHvlRD9QaSZOIJikbnQdKygUzFB7mvAN0czEfIQZw0/CYyKJ2uxdI3DQhrskwLV
V/mbSXKl6M+msC7quNvr5hLME1VmqzjlLrfRd+FnZ+7C6qXfOjwUVIYiFzsETzls
l9mhR0MirqwvLBRvd4PU15MZBvvoZ9T3TKNCVI+f+3FMRSalhRc6ARe/LXqpqblG
pRlONlAN6j3OV0+egy/jo8K0mKNGqF0VQ1UL8fmENCW47NhFilaDWBLh+QCbpIwE
XufQI6zPe0fsKzK/GyfZV1ZVkEZJuzWLt2G5WE5dR40xwVnOseTCa24K7rnkjjX+
3jQzStIm6V+JwlSsllQGn0/YyzI9g7N26USoKnSthAgXhiWhyTcFJZBiuRaIW54k
zaIKOT2Ht0CDegfb2vMjt6A+GccL0FQmrANNHOu4yw1Z8uHdgmoSfOQzdt2bDee3
7/vD7FQRyEm6vYezLwCMSlDp/RTefuRzUluCC0aWJx55QgPJ6SHiJaNHjwBBv0OC
B2ayJW8gWzAEsWGI1WnHscBMwm40UrK2K85loWByhL7rJ8CVI98KQvFHdetHrTL/
1tTK6LimliPIKFnLzyC+SumK4xFEdD4txLn69hPOmbDlh6NosK4xLRzm2FQQKYqn
oWRFiUVEzqGY4Kkswnomtmr9z8ULu8BkrFUSOxvPjh+ItP1PSqh+I+h36GFcnzhf
HOTQoUF8k8WBEyMMMlacXOpiTtncnSMywRzmlm+f0XpAR0Xe1Sf00w7AUYCBufag
+kfezEDlANJ5fltDNet4gSmJ0BhMvQkP35vKah0BdkA3OYMknHhAl6truHzt/d/E
OnooGwk5hLaz9I1aR13vdKURWWn/BALZIE8PHRzmipbtY9JI9EvMpdMrWQ5PAMDt
6nte1qcoszFGiWAyBdPQU2sT3WX5aEejuJ/Uqrc42c94aY4RINBBE0F0IBiaU58v
lIT9tkVuh34lTlV5bgjb2zM0Ti5S3uJlv7dw5wz7YqQ8T3XN9ufUb9M2zrAQmX45
YMrGq4XXrf96Oq1J2bn/7xU/d4THuVz3KPd//FMm+Y55oxvunqekAnOa0hp9hoZj
/Xo5LAmCivklzrVOVpZpj1O5VOPUOR7/9CmJQhVAixWt67NEs2S50dgtnnKOR4bj
IK3DBCFTZ+O4QrInJwTl28WrRldEmBSkkYDPh7bSfcxPHYwY6PAG2aXVpXnKcprG
ULwJri/0fUiz8iEFHtvv9+65IvpKOdDpCAPvYDJ+/9Kx1bd3xZH8JLpF0+RuzaLv
Rl0D2dc99ha8E6kF4xUOrderpxcvEKvtwcP3KmkyeZ835xsx/XOLhXpioFzbkVfm
7VhzDqzzv3hEYULr0xVobAzD0sgm6TzcRa7ftiez9mjNf86fFSlfvgEIA2x9z6MK
Ew92p7KwsnZtp3fDUKCQ3ZYXTLXNW/CdWNOvW1Dyg8HavkXRShst0rzZU/TTndrq
mSdhktSNHoSRTbx18NHfdYgekPEx54HlHg3pdv9NRLPEVUDzMwhXlElOjK09y0Pa
JG9nuYxoXsGbP32XtTNzngKYSNcaVu3gCpBmLje7lBw+j0qt4rLP5eIvQo3BGdlL
gd4MTIDhc4bCki2X/VTCqwpLBN8elUlEKiQiM5dg7XThWFepWEPc7FWKAKHtPxmq
UzPxprjUeAnJvpVUvEtn4rQr1HPKdo1Kqazz2jQzbMDB+IP61TCcEfWTAXXP4sTk
Ae9Mri1CsEtmGzJBPwHlrd97pOpvKrRrzAfjZkiZS9SEhwnSFeaSlngU9skWOVrx
k5r1Q4tRR4jmvpOQta2kCepnjPDRP5oy6XFk687nu4LHjMsJKwmmsxH0jMm7Z02s
8+s/qJ2I/GzH1nPSU7uT2VX7KgFbA8LuU6yInREH9SG8ZUOwHbNspkVY86rcqvyh
kTIdIS8bKlBjea9USSRL3UOoz7ORxH4bTisSDSYqrVcN1twedRHeur8QGwYMk/cw
8sBb2BlEgN6zXnAukyF969xWrgDvsHoSJOxsZPw38sfzVCSaLPOml582bmxbdeY8
TqjwsMw7zXPVgY1TBo1GHWy23qv3DSevyQxFhPv0v9XN95q/Dui4QaHS5ixlF01z
dgH9DUWsqkpD8uHF99cE5RNgFavGtJx1wY80MGAiUikEuU1UIpq22AP1IVqCKypo
Rvjanhz+PIjyt3TZ8x+deBCYWGbZBo0tMEHWJ3PZkAqry0DrvTGiNJp1PiRIFf+P
AIUDmdRdESz+oWmzF9QfNi/CLo+R2dAtu95b1d5tKgxD/JefQxzZfoUvQLEjZvg1
8euTw5S9uk2GOhL61/tp2uQ43dNcpFMFVZ+RcVbpT2tQ5AYKtJZ/MSBtKIqNDSUw
ckTho69AycVlQ1WG1lWMwxwuKU1Cp3RG8c6TeuYpHgC7uAq72uWTNgvv3N4sfHYi
lBb96zdLG7rrOf22n0MCWK+mYDOzr5obhd0Njb4sZHLPpcyfgFTJnu/sQMilB4yo
BR9tYXjlzBGCyPWYCxPs7yF2Nc47/JqY5TWgK0QLJXfB/t9KR0rZTL5JOcrmqI1/
+VGpJ7H8HYq+c3kNxCxFUKzIPae4PecgZxOz03vGm/pafhP1ZeOt4hyxrmsvn6cG
I2EUXgV0SMY+MwGC4btIo9iaVPI0eG8YE5L5ncpY2Diy8d8CsfI/zauncXL5aUDI
LFcM1eZRAM1TsCwe0kXfpygw9z6mc8CPaijM6LZjBsdrB9AlXeZNjIVJQ8Ty7IMo
R2802gLhOBtUr9gnQfus7+fWzjKXsnO2eDxa223hbawJtDYQk7f9f0pxTvQdc5Qu
uGUdJ1tL1wecfp/s/BBZk5HvUvPU504+beReVlfLMXozXwpqG5EurocNp2CRH/O4
Ro4fmxjlVgpcwjvI2+yeF4oVnDq6yQiSbxe8CW68nTNNElIh4MHI0roGtPHEvP2K
Hk6pfhSwocDC/i20VOj2vVqJkMyvST+9af62TbBFao0GmPJxH2+202gHdUD3Hpfm
NJp8FfxZ+mPuwUFQmp3KiecPGlAC+AiJk3mzpSQgMJKAznvn0cMANPZv9KRTVqZQ
/udHILQssnTRmWdRodJaVH4ocQCk2GooK86J5yFmcaG16SchCPsyCLg+FJ2vp7dM
6h08B+acQWe8YDtst95mJJx7LN3yuiGHrkMI6JwLO4TwRrzoMl2HZZoBLwTr2fLR
z2PyyGQvC+7ADuZHRX5tg76ceGZ506Qj2OoBiuEgAiPjYilIimVi7hElHtAfvA/U
xhly0Yp4gfggEkCrismTFYufsVljMI0e02KQImy+1QQUIaBhyRea2+zZwo4wkQyD
BDqH45k69KSGg18w+9G17c6fdm4qn3hhkpyzHQnfIiW9R8GaF8zrazT0AlgAd0pk
eSjUw34pXUWf0D15p0vbpYewTf2HhTLQbSXhRbjigbFoDcCmLzvMgkF4drzZSi3s
/BDYZXMReOU75SeHfZZdlchfp7oxs9S1qUaxvkNftFD0W/vrwBMvIcXgLOYNQfI/
5dE1JgCNyssLAxVfgNCrvzTwTRRtubW+XRvaYhnx3rqX9TNrfaVBREl+nIgUt6e9
yo+d/rTVTBaPiN5h+DaKVsZ8GfQyzQINAyAf886vPALwhYwxVAUMtzqDlDgtL74J
tDGujhf9hD1GdApU2NB68u2xxBB1kohjw52OoLd6RquPH3WY6eiOVLks9oyyCZez
zPuCP49sSgZDlGK7/uFHMYmaNbMy3rnsr+Ey72vLtOA1WF/eP4eofmF9/pu71Mur
9oUAire0tPH6NV67vkBR+dP48uiaPmjHkdwTfazYGpXNS/SaGnOob8tpY7ib+e55
efcpt4jDj/T/8WZ34ghh04s0ieqwyPPse+KX5CL7ouGDK9JSwmW6ZDLb49TPhcxk
PRnToh32UhAh+b2MKRboCLsgcTaT6xsl2R996Y9xkuUIStdWesSB/oiXFxi8hVhS
w2Kag2Hf8jU8X7nxxJL3gmejrvMc8iimCNOXidVLAf4eR4YXkJug6cop8rEP9sw/
TK5PgWXCuG9ArOYxzqGvQ3Z0j2+gZAiU1pf9WOTlTV1E5ur/SSPGDj+/I9d8LW/n
lLhPIBhZLohT5NOlkSMFaky52gms2rFmjn9156JRULgwGE+0jM8LXvmy507gUOvW
2s6Q2Zf7j3YO/DSC70GF61iRXX3EeBBEk1BGUDHbpGl/Gvvj5yIUBj1RDQYr3bgh
QF06xmimdzrGURifm/3qspSOnlJ9yFZEYlWqzqshwuhY1FUljq/QyqowulDyvFFB
qa6igGkJ/8AWQeDjbai8F5uYp5ddOMheIA7AaAkpInVmmhfnXCoj8HZCMZ7jRoMp
KMejtM4GrrAFI1+n7Wwuh+6WgL781lAgllRDtwMsHcJzoGRAcx/LqubDYttqYfF2
fgpIUVTo4y1wAGavEZq5h7gNPBuGFTLckqnylZ84xWXI8Rxo3NG6LxJq9/dumxrm
R2ahDvx9AeEpCUT3g/lpsI34wg7PFq04riO14YzCwhr3R6cDLLY+uP74DkgZ927L
7a1GE/RcM0sAkyZS6acVksH3dErwCSub+Pm8ib3W037oDZpCP+jJC8rlo/SPJ3qj
4okWpRFvd40JrNhVcxLOjQSFV8ADHhobjEQBmZicqkDLlfwbFtcMJjFMAN8lcd3D
A6jKIUAnzbKOJjYPUrPxcY6AnG725MmfnpW1gWFmqj5hViJBaa6PZYr6uH5BPPSI
XAskjbjqtFq5wFgxRZWe3t4Ya2tqwnkNbBWDxQAEXPtz6LwHiwSJtiOdksZW4PfF
om6fwnRX5WcGa++F3VHl0puJN2WaiV/uQnP1fQ2wdRwvPSarcXg2DnbkoEm0zadn
brIf6Y8N9R5W/1IllpWgHqoxOq4LrEjG5VNHjP0rqzZEjYpnV0iHqDAXMWpoLwPv
G+J05O55kQoe4uOpZhoY+pqTvFnGfOUFzV+++RxQpDTPO+vtUG8GHpX0ZlDBs65f
JSf0E7q7tui7Zo8d346A+L9P5rhdPlLd+XfTsouQFE0iI8vEOPGu9siDBugx1+lr
OIUzcm9tXGnhE0L2m0lIEdTyIQ2eg2Zf6OlRqIUfxZrfgUdIgbyzADpZbxeTwTTu
Pl/oeKbIgHdpX0tdvNexeQ6UEE2sWNHt8+mqtJhcThNIWLdkVoA6JWZgVNNYVQ5e
pLBtCMaXDWCafvVVQZtLrBeqZq2JIicDwf5CwsRI8JJV0izKDaQpeK2iswrv9mly
JLAsv07I7ZKynzxlNqWeO30Q3ycJS83tLbATWuMprqwuo/6EbKfUpMiiEC+5FgJZ
p9bW/hwzHxhASiKK99QMMVFidBN4E3Zud9W3pYU+bcyz+tJQ+obNgVk79DnttJoG
aCoD36elSIQTvQeasL8QyeYg6mYF2VTOjT0LenCK5tABYzN2VSrgZg4q3cthFNQR
KnGQvo8HLkNxDSMnNXO0kipu+9OnNXR0MrTasEGIpUP4+C8H6uwPTTKGt+46/r0F
4AlbBY4DG/GEkqOnl6JDgnnUgHAh+NxAysM3YhuEIrTBXDIB/oJvQpskFxe4R40T
iNLcpBJl7ullt73wGmGTdI0CaXO+7mYDvor2GfvNNEeHHUxATy34qHKt65H1wm+t
Byypsq5l1qH4sH8nmo02gaWgSWtu8wnnntEcGBGIkHE9Xr1ZvNkXxwQJoD86WmRN
eEbM0xeKPLP3aXoOk8/c3joYVzPRnmltuof7CpJI/l8wecaePFeTCVJvD+FGxNXj
E0u0G4LSi0zlhLgirb9jrB/WhAwGfmdGZFzU2MvTIM9eJKAh6Ad4pA1HmuQbmZ+N
3fDAitc5pcVzOB7e6rpUWZQeAcsDTOmCmve4mUZRjWAGexxJTEgboRDlCPTpuSzS
C6IkkYkTkX++eVlGj1rqbg9fw7u2yCY0Su7r3IICVLNaE26F+rtyrpfxcJN6bKIt
1SdklPeR4KfPHpUwwaydIuyK0PNJN9oPLKR1qO6QiCbSu4kvswXuTT+9gEKJoIya
rOMleaIaXqIuGpQfmfiTt45x1knrco6xMNX+6keRzRLeoKAbP9n1UWsxaajEFBF6
BRjY7+OCLoDdXrj2De+7fu0o13TgXEzU1mL8U88ezd8W+tkwnoSF4EWhVzrMq5h8
1b3Pw5cJmdB9XnOOe2Uu/cmXLSpoxbgqhg8Nfv2oHcpaoMOfYupNsynjRN6zWvhC
UPf+NVD5KZiY/TiBzuoeQF0prgx3x/A6f/lpYnTe4OqCp7N0GKLHvJTFiW7KkO+H
Bh8Wst4VDDoZ7c4Uzv1k2OKOBzWpcrHkFfrkMxhCyogG5NeKfbQNEUYGpcg19a3r
5oyaRKDbJpP1NhwFp6zAO294GmRZ/Cq6gusbj1Zu1+yf9cuiJ/lozxn7/8LaeQVm
GxfasmZJToFbOkVZvRPr3bm9pDnfHunYfeEiEvv+0sfn/pecQp92T+couXjrgnNg
A3YPgPzQpNXlu6lo4DA96+AK8k6+wG6WpDiPwyU2IY3b8f9vrXWQjKOJ3PqGEIyb
WK4BPmFWryi2o93675r7ODdW/GG2mPm+8wuVEqdWuevT5mc3ZLuTxypCGM1Gp2Px
7PLWaUBhGqXStY7KPOvM0C4hdcYSS3AEXbngBnntymCqcRlRgi5ZxHS0VcPkwp8k
VefCuDLlAg2Yh+ukU1PTAAyf3VxkgBkQlzGnzAGNSGT2MlFKV2Z288f1ZwsYKpwd
k1vKbjFB1eF1/xWsgPllQffukxDBXUz8GghWeT5jrG1NJfGoqIbM10K+pKb7OmkI
XShTwBlVwzJc7tbrig2PaziPZOofkkBNE5jtNr5jlBwKcXZrnfqJBiyLgGjOIzN6
cD4SuTRnxmtr8/XlZFD1dPZFSYd4hXYTLIn1UjQnSJDnLmkv8YFKdWLj3MHwkMNI
A6SupjvrJNQWI7xlxU845PD6r81cbZ7Z6n/5+zu0YXiKHHXngs04HpwkTJiDt/9p
mtYjampA/YnBOA29CupGVQS6+4piv/ZsLGRXpOIngt847obbrfFiyjyfoMlKnmWt
0s8Jp2ax7thmDKjdeclSrooVx02kHnhWpjdReCH7gMjIeCIYOsY6pMGhfUQGsSBd
lZ203XPFAs00n+P7dGQvcDYDOhxET1VFWteijVFl9noa3NEyzqwqaV3nSKZq9bqz
ZYbA6e9DyTVGeEo1/hOLBpFtPUW6+SslzZSs+ZRxPz7PmU2gsouGTscwewjBSwPT
qHs3GPf9QX1CNzWxC5/igGOQerKO6lvt+UCm+MZZDMu4MVZyhXpfCTr0MeIH9SXm
sH+nvRw2JDb46lCgZNGmDg9Qs0gN2mcnE4dVqcPpBDLatQxdztR93qqq6tmiHgAt
QsP7/njcktqYygfNB9jJc38PP+nd0V9Hn+pL5759eumoEhAG0+c8F7CcLsamfsZi
2Qa+lF1ayQ/qSUGUWIYwTlnByQnPJrtwOoMoeSOdmE2mGEOHYOssLgYZuDF/r4Wp
uSKYchva/t+pThMpvS91onRblPug1MNSna0cGfYvyW8oltw7jmfIfmRGqleeXgmQ
zXnrCdkxUryagsftULMfzvOfduN1TTEdqTF1JsgiFS3bDdAdqhViGjjNL1JfYK2h
yNIngNZ2Z7R4IxIOCN+VPKmBWM24dvTkml63O4S0omEA35CQtLzVN43cE/0r+x54
p4URvGTsMoAJltnuH9vPZeJVZa24kRyJN56bX8Ia2Dc2IKmppZ7hR/PrRSltUws4
yZ/mPu6YDa0EI2l4UKv6DhJ0e2ZH5/4+A+5EZxUT455UZ5JO34TLWQCpVK2rxURm
TuR6NzFxTJeAbGZ6XdcsWExajoE4cdwG9G0HwtCffQQ1/m9i3il4HOnFRq0nzLD5
aBPQtWsZNdv5OVx0wRbOjpw8+J9J6OXiwwT6Gl22Uim3ezSKoEFWEdOhRD1yXCfS
DZSun3oGurPfnX7FJOcE72zTiYfayrd57Aq0sFTo9VxJuVkZabx4JNgYL7xat4CK
cm8RD7tychupneVtMqmP8nxtegW8UpEBVwvAbr1vw6hlTvWSoOLfL/DH/YEillx7
NPAPOkeVk9mLWOJ/bfw81nEXHvHpler5bYGEmtrPrcyiGQ2lBDGFAn0stLrRiZ/f
lFM0k1rnZz2NeLXcHCJVo5og8lLhJ630+cQpWUkb1CEJH+dTyn5oNUYgRc7usWt6
xTgVahz5mXV0cKLZ77dsztfsCvnbA73IRYbM+yVdeNb0EZujQgoYfgxZ1mp1fXCq
3yTOd4fHDN4lIpx0MK1SFsj5WvCDv79bC4HMbQ/pebAEbf9vSoorXLBOsUy+YhdE
U5q7Y2+GCfKuRA/iJmcZEQfEkImbumWrog/ZJA8p2Djt3aUDOUTWROQInPManNZM
0uKkS+iYTQAIVFUy2QOuv1HjgC4UMIpFiXkC0BLWDTylq7OR4wcMM7Qfd+zHFKoS
3/oLjCiZcn5twOQfcd8n2EVWyuAjIenThXW2Jfh2/CBopV2UicttPbqzT+U06laU
OOFDyC4jMgfzlLVJGoSoEnRT52ep1MXsTeDe4lYX+abdg1zP0nGrWZkSwQznUV1m
88AITJHcmM1vid2dt4xlogEg4wY8dDYdWlIf0Y6u3bqhiIox1YAIai27p5fg7ksD
B/DFRS4/xW9uNoi86mVAcLtdOJGSL1+GGGpy1Lui74mfyomcZGvwjGYhdwFw7EGy
5IwVh7m5MHveW+aiZVnzi1L2A0ysX3KttdIghoo97oWVEvRkajchnSMyxZZDpwQX
ODqbMjuWPjPF5vUkKr9eGhtHR8Rif6PnEwZ9LB7QxMYuRrIgJWb8b6l87Ba3n4A1
fkC0/LAspts0+C2XBnKUowza2/FIR+t3nGRQOdNHO0e2IonvA8fMTaQz+Ovvuzpz
AysxiRzivRj6NidW79JyMcfgtZYjmmwVFyANpJ5IVxsaBGLZUlv50Ejfvk+pP9wt
JlstWo/LwX65ODQxF0SC8DbnFOF1YCQoLwdQA6hIA/T9BfZSfvze5YSlz3SodVzD
LnQPS08IU7b7v6KJ3ntrHEm/cp05QQvVXeis0L4O3siOvUH8bFw/vzXoUl4GDRYs
DU18unC8rTevxCBGRghstxr8qFyafcVWP+y/CD8I3pIazQPhqLWu8MTJYvvgcJVG
5fCQ1ceR46kEVUk9ZCVO7LBTWeVlZfRYksyxmP2IwbmgWgjsBkofEYpMV/yLzM4T
K8mPQTik1MgEJPtsI94fDhzAA7A+qcXqNfUx56yLjuMPGRwNhW6g4OmLK5sPcn2G
wtpR+C1TZrdhI2RrsBT3h42imyTais3mbrxdXYIGuETd3hUjgWRLcY7w38YYtQzt
apl840yz/z+yXhyjcK4rUS0FGaiZbHxP9iTO8xKCFZmCQd8tInW+c7n/9SSvu/HO
gHGaN0WtVFV6lTTimGx7jF9TR37+w+65z4Nj4BV+GwOgejZ4b2Z2dKxHePE6dfCR
lV+obSunP4vvnq3OGy3X8666pQ7R9U4waBoX+nXOV1WrMzUfqiylgnWwuWjoCeXC
KwojnVFZah6vVGppyG+pvWCRUqFXW0Lp74/WUKX/j2gb2VPXFYw4VWGWMEsLUJ2Q
6ek5BxC0BpZmleqVKqklHrEaWbAxNF+M3xVQyUuPF03NOAkLfOpdiXnt/gbmR24Z
IwSiTv7sFDj2WOPyHKs10N8OuQF2lIOiQOu2Npmg263ovkeqPF0QH83c41agenzO
leDa+LSqdlcPJ9j/xz1U7K1W0SOxgOs2P4lhp/p3JuWYvt4fa8yFa9vfNlmxe7bp
btij6BTjwidm0LOLlhxc6EJWHcST0sFE1LiRTpgaZg15bw84RfAe/VLLrHRL2ALt
6Hl8s35Mrjq6RYnCJV7eC4sjsIoqQZTWs4sT/uzA/w/a8UYaAAh/BDV//SaJqDdh
Nf1NqM0o9o147m24AThJWX0kHbmL++Mp5SGgaro4+Tox0qMnN4W0m+UGA4Jf6G4p
HvwtV2VJAWIF6rUHmBZrcA1O7yD4QOW+/yyRZ6RRVZ0byl136EZo9g0JBuDCuFuM
t8kmZKSST4BzxjVLIaolmZ4uf74WDxS/xqd7XnC09uP0Z+hPSgb5rB2274AEsYYg
JJjDrJ1qTUkUO2tqqO70UIRpG+sJe8J1gK2KgF61bYu10IfN55tfRav1/sBa5WvD
26aqfnSkTYjZpBE78V8aSSQueU1I/9i2HssiTQpMZK4+pZ9WD5G4s8xBAiVr3YNn
0/8RTjGEfMCAcX/w3Ij9Pd1emAENFTUF62DglpxK8HN2VENl5hTokFGWoprBD3w5
/4M1bD+dN/eycf1GPLiaYytoA1wigL7afDVsj9kGd0iQGXTM3Z4S8KOkLi7vamIA
FyZMcc/C/VmZc5dN8mLPfwHncaG9zsQmvHvYJvT1Vhq3utccIg58fhktEsn76UrA
ux8NNRMCL4k1SPKI3uY/S8bLZLXjcClr/3uamNDQ1jXD/DZ02V5u0Y8Pey2Wk5T0
+6lJ9uArYjt8DBtJAPi4mleNt0gt3T2evHXfgKG5I3k+hFGB+8ZTS4pTEE7w3aur
bnPTZ0/jbtfE5X6eyUZDoT2ncjiaMuP2Z9GiBdD8L4XmS1PvVFfe8D/LUT5/yucw
83vuy7wts3sc+CKrvKpbjknSPjH41c3vcMqIU1HRO2/HKPf8mr9ffzJRjbWv55js
LRlw1sIg1t+H7U8wCfJew9e0xremXcUks+v/cyhPLJv8Q4Omm9N3nLMZiDiu4HgN
lgcrdwJBnJ9JGXaD/v8lhCYp69/JRgkLzq6LUg+7p4rK+nvTSzgFD+SYHsZeoCfb
71hxy2a6pcahV2MSraPRgbRIiHxPuMdb8+IL++Y49TV5CvBxCmhB8L/M8+uBuv4M
YQnT+gcSW6SyieFzXwwqfzqI5lQ59nvwUSFVNHG/VNdlFiOtfthwuBLrpf+MWW8W
BiiXFcSzcHjhq1uxezzWo7KRa65IsL3fF30NAZ28MbQ0JJ6VUoowMUpS4dIpTUC9
3kfilVgBcDe/WRCevYvFNclRcu38JTK3irZA61jJKKrE1aQwzEp12hvGOc+ZaIUP
+i+c4VMWd2YAbVlnhfpzB5KGnBtWPlaNcatqavJtrDJIJyrFS9yXr4CfdJ2Ro32M
RsRTATB6i67XqWpwgmZNYpH7GV7KrWmdGYX63sTAZdr0k0cYzke8w5iG5vB37dbJ
l1bVZnhah3+7QnibbJbR9CwcnYtF0MkHHij35NSIR8H4t0T1SauCJy8zgzZElpZz
64CAjvF/sPC4zYnclnHPmpryTr9uZRxj/iLeJAM/hYcSV7NvTCv17Qj1b4ROy4XN
L5Kq2Ebq46aID9aChXIzYlg4uAJImLKMDKRCmc4Bfx1BiZZiMUAQpnGKk/KNW89U
Xv1M41ibTfwdN+ZHhIoKxnipcYPQca9U59899t/Z43+DEpWeywG9zqBcnsgFVAq8
BYcvLYlBrnfPLcNWRpInYcD3CVwedqwawo9s8bJQW5f6fWoXT+zYUMr3OsR92k5X
QJZp6IOMWCcDudXwlZw9yxmI7Br+rtQ/+lQaJaCkQJDpvjyKJXsaMTWdbi7A/H06
Tnlicu1MiGfMJ1uSVm2YPJlsQ5t6JDMwShfHXgq0n4BfIYjfiFx6bBMvrCuQQrLj
ooZI7EutbwdFhTckIWZngw7nUKh28rcFIoby2N84UcixkTjcFAc3It4X+5PvHd7h
wl2qvmFL4NbA4h5DBqqSlwo9bJ2bkaQBYZ7Q1u1FVwTeSBnLOlJaGJlK3hs5+9UK
qvgGYn6kMwiU+BYRrcvT7yUUrBaFhxqEE7cBPGZgIhXrRIEDUGJFcMluqBrwnKGW
RQiKZ/FzogAhYU8W5EOBpc843ELKdxCU/uWsA7gawNEaodmgAjofAthvIqDn8CRv
Y5XTiJcZuByW1otCXRKywMDgWGzD5HTcs5EKSkxfWE705l2kKVFttgsN4ubhfvjo
5m8P9iwFoFpyNz7CsgnN22F6kBaZHVDP2m2MUv1JUzmGcvYOyrZ0NIK4O6YLjqX/
gB1Krw7B7g6I2wrj/N86mtMu+seD9r7eht9xoUw/fMjNqhPhuMxtwDSqH/3651ig
AFIInoTkFXLn/ggg5RRPxT6armQR7KqAnGRfUgrBu5XCndFkoT0YYV6bAsRFA7g/
nUSkmogLZU0vY1WHpnlHHxvFUwJQwYGEaBTyJFCX+QqiemAJWS72uu+RWed9YRFo
HioxRzrhZli7wtzDScmbFo4YyGLc3sWyF4unvTVNnRHjosseZ9q3w49Nt1R4S01k
ejxO+Z2CzWXXRQuTnYAFMcc6T0Hu15IZbkuT6fhAO/hRxU0Qxv9j2J/2WcOpVQ4f
vLAOUjgEGSbhaLZ4Wm1AH8MzNRbqcsEGy+e8t8vn3gWi5jP36jICRv88eA+nxyoq
Qfe+bHsDArf3U00stNXwFIgPfYvSeVMnrPteQGfoQCyehmBtl1vvnUcoNd2Pa03p
YFC1vQKx3vL4WMHGKB/jhjwOrWRuahtcFdl3EgbbD43Zcsz933eYObctRj5PTpIk
mdu6oKlka2nOBIZheNg9h6e7cwOXzoEmXwrrvO168LufHzUvQZHjya7QhTNF1/vy
LlTpmSp5118B7lWC1nZ2tdHknUcQXvjkqzphwAyC4p5VPgFBwb3HamUyu91pU6ZV
BrljGzQJOZ0sdfLmfw3QNpxBK1IY3f/V+KCTZ9WO81qUXW6XVW5wjjIazyM1fh5m
o4yTYoyi6EqS9bzzwS8bJ7Sn2coq8KHxmgFXcqyrrJUtDEhMrtRLPO6DRUSux8uL
bzle2ThY1w5Dw8ekSSRIROoQ7PQrBnQZXqjiYsx7WBcHV7/YG0fLZNUTMJFv2k3p
9YKQfQ2irroLVN63O/ik5YYCQb4ZXbrTouAiHMK4D8V8N/3FIdtGG4LbbRkSXmc1
X/8zvCeoYN2lxpX+W3P0iO1FFe1lcXAqQZcG21n+NaATIzv6r3rwdMdibkBHR2Ru
M8LjYsZQJx/wDhIUO0Gj37czUkQ0iLW7zA0LuYzlG3x4Hpobpj9rhcTgnDl9Yxmh
huOpe/MlfcChX5cHqijs5r5vmAx1hoimH8Djo3v8mFC6t9l78oohssNcyeC4aMD9
TgzAzsh/aRknIP32uFtpVMQbTxsds1dU7zzknPSYF9n9MP1WwWSg+pW07kp5S95J
9o8fc4eIsPjJMomdPEBUxC7OgkTl4noC+AjBKTbYz3S6CaJXSkFBJeEn3QHtAxEb
mJ21ulnpUu9qkpRMR7iMFUpcjXJvhzyRBsDqTd660TYEMqk3dW56We/lb0AyLQqB
Kwea44vs1f/0uh3rchnqha7b8IDxISkOw45kkFOku1wv2Sf1Tw8TTrscdYWS1r4h
oGMxv+obDXt5Pt47B6LQ+3JRACGps66U9jfBw2YqYcDhbeqSosItfqsZgfia0R7r
+xNRAzZ3JfRlPUa46Sa7JJJ4o/LkJOIyzWc4lNTVJC7BQIacwUiiSf4TNLRGtSNR
8HcKcPJdFDW9eDjFqKLihtguu7bFvt2p9CUe2EX4xHYEeurfJqU9u69OTSMb8aAW
wDndPljIqirjZYxP0iSt5owfkZIlwmBWtI71FGcvEAut5+Wmox125+VuPRC6IPOw
0QmSmdrz4f7sCU4R514Nv0Y4dq/t8kpPkM0JDtH3Dxh6zOPSM6+Z0+3jUvad2Ncx
hLW3RhZWqS3JjPxukpKIvF/XN33sNa1he2MtPuGeJusfvcTu0l3tPOBI/OhKHyL9
NmbdYSBbHq9lZXYZfRtYhiP5UqbBzo3fibQNI6/8UzD2WvYUBZi8ZA7iSW9kNMf1
2UzBVoshmYbAu8egTREy2vIjlSMfUylxmwh6VbZ6ywLjyhDPvnFaoRtZesjwxvSv
UN777FNuNtFBgFQFh3Sc6/d0xObbp0+cESfW65oc2t+fQUMCKS+syqNyWZECZUp/
T/w/dtLrgWjiKnzPeVxul++YjPbyfapE3Z98CU4KpCF7BP7iPTwISIYpa03Ov8M4
u3h9GkVdagfE3tack6dVnT/1iQS0FoeYRijaaj+OezH3bZynWDX6v2CA/SAXGfhs
N+6OtwnGi8NZ1EYOfmqOTYYvyAcELCcT780hEDzKVZDlxRLM5WnPHbW+Y7CVamWH
/jgccvCtF3Y42aLH5C5tfGQEDBtixRX7ZpAAxNVpFAvPJMTPhlpqXiSBLEKjnC2h
PebQVlNaqgM/HWIl345hN3SSTI/ylbvCEBCq33KqJMlylWsrIpN2TKPX6sgAEuF6
1E5P9vlEu1Qc9UJrWjOpESqH0mAhiyAX7CnNepvulZNob6BOk3uQnDqyx26EHwyl
MEDcyHrdP+1pVgLCjV8OVSjLjJPg7Y5vgULyZSZfD+WXY6efc6oBulmBgfk+g0Ti
fc5Y75Fim9XR/SKuiB4PR6uJbaj2JkNeJ9UxZuS4Wvf6nxFDbfC06gxGDdBvPvFr
bKMX2v9S75r42kbM6G0KMmHonQ8r9R6kXkAZHIdTUUJCM1hh2DtZLdkxmqKDkfos
MF+ZaSXHpJa/OzbCEfZDQnAWJHtPs8/WAtUf1wnwHUMy+aGeFDv3xnO7E5JY4l9c
j78qrd6TXps32jQjTR1KrMlmp4L1FtZvIH9VaHgbRLzhfRHfK6qa9XoBo4NdNyWz
Ewj7N+2/AuuNDXPZP4ytmhi5KK/v+Oghdd9g4akZbOy/e/U3BywJ9LMBLJTb0qpu
5JP/I5w0c92/4TBqyU8t7X5xj4q9Cf95kinvNdjf2JhmfZmaRbO7a6JvaJI8OSQe
0RenUzRtU/Lpe0vtjOWKlvIPq4AD3A6NNhCEYdTZDj3eWoSojdjZtIPRnhaM9C2N
QkJLH6K8eb8CpGuX9VtAcOoTRrZM19XssGllvaP33Ph/ipSFDIcumA1URIJk/6UM
CqNKd0LBG8xVvC5y7yBf6vwbujmTRJdp1Z/NVZ22XWIMKzD8u/UeqzPwzcxavXK3
+rRm65yk/LtTq14iCRv1KwiQ/5/06m6Iu3FYMlO4SL8cxtI411IGq2+nYtIt4w4K
cACyVejNk4l8KCdeiw0Z6EY9sVV8UDzg4IUkjpIgZqs3uGXeMwZRtGQah6XfQJOe
yWvtJQxbcFZVfGgvRq70d2sSa8nyiOabZenUfpqMPeLvv6/tkKSKel+QnWrT8T2v
gKCCpM6fTitJ2i1qSImWBXXgMB38H91PmdUN/fDlgjNvIwLLcS3bwBWTVnym27Pz
C3Q9Gu/VNVDTlCm0T+Xa6yNuA5BulcHNrNZNkJrz8GH8rGVmRJNkI5U33//tmb3p
ObcDTpKel671g9NysAZ3HA1HjIGn4kAHIZyBk8x4Zh1KnDgzh5zAEM6aFkCGNL0E
j954eRbkmjr+MjYq58X384xjPD+IYJkqwfBT5baBZIY9b5+hDDU0LmlapXz/Sb3a
K4sUOWk2MzP7xq2amilGsSWDmj/xwhxP5dJAETQzo5HiPm4L4NCpaRWqbUda2PYa
gvK1QecLgfUKqbxMt519SFOw3PDdq0ZCgI/ys4JKgB0g5SA6ji83YkS2kPyueMzY
0D6jLzzvpKNZ0C2ao+gp9TA5IpBxvBhEtKWvx0evWWzs11cYvu6ZvMFUBv4CwU3L
KISBCL2CGYBM98KkCOAaPCMDu8+AeyWHsyua7mSCDEISOBj7xPpOVv7wrYRciOQg
Wrf8DwzFxK3gahUaLWevwDTcesxSJaVO1lTZU2OuCYwgvYHdNciHhxGHg98wO1wl
vvMs/ybw8StRboohvwJPO94+Ibz7CxBVHgPKFCPSHLMv2O71EfB2jEWI72mcuArM
WN1TvSEI/y37d8T7Ex6igXaMzjroB797RmgT2LcOMcY3AHn6qyOARx0tdwg00HPD
ktwZC0HXqeTI0VAj5/pyO82GxbQFSADWw8eS8tWj9DCSlqMh/kCUvEs4p5oALiCR
TemSZfqa0fFsq+coJXFSnVhNdCDMoLCTzBC51xx3VTNbQN35pLdYnNEM8INhDn1S
h4KWXmsCzRUGdHVPouRkHz35gle4/ad6RYn2jcx2H09ooqov7bOa6yJm+CQt4WIG
hQ0BAabevvbXnlIk1fg35MxHhoxAdkksuJPhsiAR6AcuJMTK9EBM790OP3wmoM11
l7ZQn51cnGVQC8RbNtZUFApRglfKss7T2CUCjj4mXvqN8K2YERaD7N9zM4dUGYSK
TrnmXmAsa/888ot9Hvwm9T30ySSTQs5A831OtGkxc0CBm3JcHUy2v3sDokcGvqRp
AYnD9Qq3o68JdHvR4kf5VV14N4vQwkQUwF3FIw0uoHPJWEPAOG5NiPruullZUmxf
2+J15qBG5U5pN1mPILFaXelNOZMliuweYmG5bC79GqSqrDMAnKJrQMZDpnzgFECL
ADkO1Q8b+l98Pj7EskWz7ysjRRUaOPTgWAGTLKaIT3PlWt3S4pfSEFZu5iKNiGLX
exqfqEaA6W/qPpi98Q3W/rKFVoneN5cywBG8r2svxzCPrwyZ57MWTafVcAUx4HGz
kWTwKWLaJ3Dl27D+gtqIa1aDW6FzGUnKOp+G6Re5Cg20JkVvHDIhpMupUOkkeVMD
uaCLcugKPMDgOXZI+VgtwsXGy9kjvM0qj2wMPwj/QyIMMvfy7B7i4OaOZcyEnD2m
yhmpOnbTWlQv6lIy+stgw0hgFyymBN5PeXOSHEebBu/gyjtuwZA76OoHghCvbqOM
nO+Ra/GDE3jGzyrzYlRWkfJgRZDURPCN4y9dE5orkXSIKI1Y2DFnZT8sA7T/VfxY
v1si+Ge59s3d73Q7atb9g1tUdg4m4vIn9SFxSzyrGpPEFtvHw/15mg6GOqxj9DuZ
OF4rj7u4qO+Et7ft2CnYqSZc35/1sZsEu9na1eWjMvf2S5dUnLqjQ4o45RN6UoJg
eAF4/VXtp6vAxn6agcE8DNL+lpyMVfnbd2E9Dlg66Ws+Uh2Rv4jTG+eQdAFkgjLD
gLYGRjPR5DOl1GfftoPqkgZPcImvppv6S83nfN6bnm9IgGD1UDND3PyFtfLF6RvT
opdo2ZYXY/oEH+oOJCf7YWYrNx/Op2uvP4P720XSRYFuQnG0UzdJU2haYzrChfs7
pfsq7p35r7uz8fdSf+ZRUt8i9u26MZBMIZ4NcFYL/TwkVWVLkgF8R/iCsxuDiLsz
M4SOSvq4thR0ylQyuelljSGD6cVyGDn+PHtBj66H+zPX2QROwewl5J0w+daX62S3
k5jy31G2TylpoKJbBsNxnt0OZZTb22/ZRVQl7xnF/kXCF4szg+FwAlxkC5uop7ww
2KPMavI6vt4OLApjWCehFx2q5MFO8Z33ZLQzneSgcVpBjph4oHkM/NrMPg3ktfxo
ais/ZVnpk7/mxe7A8bGNW+j9Pr9YO3yf83pKs4OqX0Y3R+houw1tojD7s+5CgcYu
fJSDIhumMK/+BZRDRdTe7ZhKsbG/CDAxUrAEJaf6d+XJ/HDE07ZWPFTix8kp4Qvt
zemUUtQ32HPyPLXFGgDKnsHjUpjnHxE3HarYuOyMP/sgQzp0QexY6vCrK0ttMxuV
HYpLD20lJ0azPURh9sdws02yZdYHqB+NaOaCEGAVWmk470OBu5XUrXDWK82YJEbQ
xHOJf1LPY04lVeNiuIv68LAD3unvcpICw+p/e1VyeiQLVHyuo6SLG+pk9R9nW+iW
DGuEbyueujJC95W8wfPTcZAooHRe5TDkCWbO97LSPDf+k0pqtjNe238FQGMQfoFj
9GUtMWXACUw8RY/c4y65G6w5KC+kY6SXqSXCbeFDBAoLOmoK/tUfp5e1gQJ7mxRp
APpw134HeZQhRRivZBgUylqsFiGdpxWDDzi0vqWdcNefsrBRWm2LFjM9hj0vv337
RVv8/4XJRwK6Oo/1HFYJHB934cA4a6u5/AnlHflbDFSHLVR9E+17gFXNZHuVi+Q1
TQt6SRFJb9b9xIGtBHhz6I5gS/Ew1vvhl4+anOCh1zg8wJojjEfD0Z/vrfFxp230
5RT2re/AOJZnJqhJG+8E/1pmPcO65Xamj5tCdGvzZ6mqlXOnVojL6+TQXIgpu2L0
VMEe9yyTmyiYzdiTJuGs7VPUZLoibKz3TK0LoRVHmjp5E8vaZGXu+JOWLnn1ouFB
DNxyKR2tzQlIs6fFNpupCXYWoMzPCLnEOr7r8KbH/xL8NdHh/UBVblh21V6Jgtqz
u6IHAcqasLJWmMKrvjiq/53v0zoFX/VYc3z3OaXJP7YFMPqK09afYKgUuxWsf8lY
5e6RvSnpIFnKlVXJ69s8Nta78dgvRAP0R5T3jr47H/+hUvCd2oZK0k08kvZ1Qijj
JutplDdIXupB8KNra70wNwKKdqKCWyUhbwRgMbdy4wwm054bzXa/0OWNqiJKkpZM
hwtaj6LkrqZhbnOfDq2Rz/d4iF9Tt4R2pyDdhOmorpkStYzp0fIOHCgPS0CGx9qd
9bzx3g1NvQ1j2XjMp02DAOQKas0cjJhfZSoxZEYZuiwfAKR8hS+wDuD3RTEOc1q3
9h03tbsy5tjPhdxbcAqKV94nYqJBhGYDXdkaUpcB41f27x6D29wulr87H31TH3O6
A610yrDJ1KyB3oTe+0l4uaz+7PEzz7JS/QbAA1dNox65+wgxQ8wTRI6MuS1RmFNg
iYa3mcc1VnjZJ1zQOkaf5HvkCbojZ90s8q8s9lB+xtFMNQHFkFdTvQKDHDMCsO3w
3ixJdDBCtUE7TfBKN4Hued1s5aH+IOzkv8cfvP6jkdX98dktPi7bibBEPnnMJNf2
57bYRRw7e1ThhK1j7MQVYwxi5TuigqI53foEmnhuzjL4LTiryB0yDSRZ1EzQC2y+
2UiTk2L/K33ba5KKUbLpAMzVGLNYf3gqm7V4ISb/x9TfQdcEzw+bDVrw0QsZRucC
eHu3uZ/DLiuUF6ZgDvnTnbu3nTTMDYxINoIhhvnOMUfOXym400yoN2TMbtUZksxU
CbdFhcOFcpE5NTVWVIgMigK9uI0k84CyKIUC+2z3dWmXLr6SlaQ4C+pK0Y8Pwg/9
A3bp6UDNXbWGMx0U7/qvUGxUGSZZ3pT7AbGJ+FXOgFpMQxrQ0P5cW1BY/obXXytG
gHwuyMrErXmk0PSlf+K198RbT4di4kJvjW6jqZmm63P720ELaBvHVvDRXJnrSE2a
qQ091Ri2Ynp+1vh0q6Qlz2K2A74Aaf4jnVuhF6CllSFbZdna93uEDEwmD8W9jv9t
50LJCMOpSuOwduObi6RdfdQPN5Xe78I8K9Tv4BGqS1MCeOGdPsiMHnc7UEle1els
c+Oh8StrpnCJ80qzxnaXCCxa9OZ6vX9OJ1g6EKJZqoXq5PY6yQGDoA9VEbwwOOjL
8TX4Qxx/DbqnivPLzPRoiULGgxZu2Dm2+P5o5i/n2ACScUPsBjJ69KF1DsTYxhql
ldlK3GZaMAiaxffeiHfQAY6iNYohNlnqprdSSe06aB0AmdhH6MCxfJdEW14m1m3m
DsLsGiimRu27CRvt4PvcUEPIqcOp/ziVzRcn86Yx/r8amY2mNMn90+oQPErtuc73
36+9IXgliGev3zHF/SFbQ+0n35BkEmBwtkHabR8dKzvM0ET767eUpOYWKWQzfajR
dfFbm4QuuUKGMAa5nIm6QM6snppmETC5ZIgXiAO87TbB7aRaexMkz7LrHpDkGbNW
GE7J6O1B09SNCXDTH11WVM8i96SP8teasgc0pUcjzprE8jt3LfqsN21bKqjj/ZqW
pBpEkBAMzje7GQIYvlJBAMC0t279527xcill1qF5GnpaJMPI2jbhPLMGyyS1SWpU
h6UDjw7KAwSDOFWZzBTmB26VfMA+AO4orHysNOAR+mTElVAJlJpbS/A48EOK0G5T
4EUlxtZuZv21Webofc+xYJY3i0LmHPb+xnZeTmYyXrsgB2Oi4omI3klgIaWji6oy
+KdPkw9xTrO9Bxa34G3eADiQB9hjvWQco0cJg+QJdOLqzHDp9L83D2VjNpR8kHYE
rA0ugEWFKsBoBNJoOXa50cfvIEzi5AjzUGijaJPN3n99RV4PzGiC7/yy3r3MrbTY
2WtdOVdZOTQGXfxiITf55Nsdc/np/AM8W2OUHW39KXQ9SCa8hmgsf1erc69R/X0D
CfDh6PMj8bm1rIxkvZVgZstKfXMmL56mZXwEzxIRx48fIgOg4Fd+OGmkC0rtVXkN
N8GXpim58CI3hG+iSHaujfDB/qKR+xK5hIh2ObXupOYG+hLmN8QVWTC6Ik2OH5lZ
o0e+g7OPCowDXtglSlRJ5MktmO0mT/NAomxjL7LAwlHXVdo23aKGvTO7WFr7CaRC
ZJYcXpGmq+MSwQvvnmQtR1yMVPMRferLBk1SsNGgOGISL5Cs6Jkxx0p9LWDH50d6
KRE1OhR3V+WW/Z3+QX6/OIhgDn2ULugmg79LhCtSPO1SsX+Az2fyumCmffXaNIcI
W5EtLaEt/F5fPlFFRuvNIkAyOTgZxxlRL3AbVLLO3V+20jdzr25EWAAlNPxWlYeE
3e5wCer8Njhb5vzib7tU4be/kK9NxB1e3EgBNZcenilM/N0DcRCCPP0ytRHeEfw6
YfBbHvq5uMXghhj2cCmLrSTvK+OSXCFihjvOrROyAewP9fIQ8XSu+6PNA4YdqZES
IKRJ+E5ZEoLMYd6HCUdc5RPju5CC8YErk9fhEFJusFduSUOo1Led3XvPSATmjPFH
09KflhWY3ZZGkhPPeLaOp5/vzatfGp8eE3fycOOrJOAG8aAOKji3ne2fAPr+Vd65
4oujwdfp0pB0sx9whXBk3ZZivKkoxXApBkv3kQCKj2TPZc1c5HSxpbm1Hq2utm4x
otM9h/TZGWC+eTOhcUrOQsSZNIOo7R+BAvp/uhZktGcZo+DRCmqPtYU6LQdaBy8B
/w6I5bFi1zEMGPf0apE2dyciwluoPuxFsYhlRkjq/sUhrW/qIm8sxuW0jdGjQILL
OHtJUzTrXnziqCB4yFbAOJm7+l3dCR8T7n79FDsWcUPfyRZ5GTFOoYIZ9afNkkrq
CGqyILv6IPkltKfilVRr6BEVvYuVA4u++/HaxRSzLNFdwEfNX8tU16eM/vkUyzOE
tpHbuTT7IqY8XMOfT/W+D9J2hi445SAMFdjkwS+wSsdyCd3XvQ3mDqF53XeSx7MH
8wXvQ6Uc1spXbEmDttjqQlK/yEqGKijQ6ic7HzDltn0WOuUEACU4sVgDKa9Yx2mu
XkNNrEMP3tMZjNUtpAxYp0FZuA2vdrlCzEPtlKePZ81zWZ6VAANKKT1UrfMoUgrP
U6YlKCvd9GwgfWxE5NlvGpntpDskYbNqBd8wn4e7StJCjadjnRyczIDMctBP6a4l
l4SgQBrGI8A7eUrCokJhlw1ucYnYlSfk70uBo9T6QIo23RMRjr6jc56QtXGD7KWx
OWx1/rARncAfXaqHtOsYqqpZwxQaqLOQigcFo5u3kpQLK252gf0WYTPeEnOLxeKI
3j41bRvhoazyiTqgmqi8kFQEtsTrI8Cq1RPmGESXmDO0WFWaIuXF94AnaBY2EWCj
YdhDZiLDVEO99/CJaOMdWeoLfgB7slSzTTQ2XlRRXDc36cO2fa0hjpFEzVjOX/P8
V2Y7aWjPj39HzOhZACaPJpaGh7VAoJUpEQzxNiYWPrbV8G8vF1Owte+PwVoMbTDr
l5+2EIYxbFiTbx1cne/DSarOd7ytpEMOMZZs3itVKd2I1oK/ExsylBhp7FUh4KjH
/v8SRDL4Hb97vFcN9EVIkbw9FR5eoDPd8HXvM+APr/2NwJF+o3mxHaj7COd1kEaN
UVfU6R7gILXa23G+uO90l4Lsy8V5BwMli9r3YLGpopYyqrSXoQxivpBFZsHFpqix
drdJn3gKaxJXF8RKsWxOYUVBpuLTSY66j1lBfO80cifL6QpO+4sD1aVb+phC87r8
Mj33rJTLOpWmCjbnS1qdQ5yd/TWXPKCSaFa8i8lqENgAvE1vognA7LMAwQOB+9vP
30jF5DjWun8x26rkXXypl1ezfsCC5FaRW8NPuAC9jc8olLrjuw9FjifIkEVxaLoN
2Tp7FRzg95o3u6KWJ/a9KOu/Sa+8AXAg6aYp7WGNv4qpIXTBG/E9YYISCzshtBwl
JKOjgo3HUorvhOElvzdpC/S/ddee+HoCkoXcs28gCLqt/jtWnzmcWiq8FhjONe8A
LA+nGf5NFAn0Emkl906D2fJttQ8Pw6kd99l8HO/rz+YmXIbIZIKSMX42QRv2wNDL
sS4xQOL3soNuzi73md1HPEPgpVTMg48QG9wj6+IGiOfcmKUXxDiFynvrskWV7fmI
LDnoAPoqqPlCzvzgJrcAOPq07YvcXjq12Gii6dCxQ+jr1K5DBln8EMx0U88zNyVp
MyHETCBCNFPDkJFQ1i5Yq9DvIA5SNcLdQf0gZHjv5uGHOIWzBKPTsB8kQKpdgX1J
QYdD5J1vJuFFiYYLhvegBJC9X9U2HfbKRAbSl7Gh9AjOaaxd7MXbyYTaPCBl2guo
AFg6EQjCd0tpKAu+5FE7Xk2lxWvkGrthWWeyPVyQH9Dq2ySwzZxBgF3Xe+O/wJvH
pYBS/iIUIEV79ZKaNxhczpwVyXVGVh1KwP62Ms+e/pbvhhEzNpkMNDE/lk7QpX/E
c27c6mg0NlQg3kZ+zCNSE+R3pwo8S6BDU33X3kf7kye4Y+LskGSlUsELhufwMRW4
brguur+pV/H8QJe/yN5iwL0VkygZIJkHyUhn8wOJs/3RiOR/o2N8PbdubI/aXiut
5NCtJPssUfim7og97i8aWCWfGKb5MUlQIM4tCyCxPGlAbTFyE0htGKChUEpT8e0v
2AOATcisrbDQqGy4hWSOEmrfcZf3nQxgxfCt5AurDooG6b4czp/35mQ7vLMz+76p
nf6xGgYifwC3evvA2P/dMT9sBUuMNK2wshdLKcdto0cM6nCVT/1/kZYHWRmQBkG0
RT8Znjlo1jgc+vEB3QafBQphxf9AyoPHvPfG9uXu9s75oxT6JpLQneVMTHPegNSJ
TgBmLaJBiPHbOkoBjlQ7CCuyiAuRizQy55CgnBooDliZJOYViMaEQqtOs2KhKaP4
+61I3E+ixGLV4JtMITvT9OcBejrJpmzBa/YOx91opv5j8v+LtgAZQkFzlogT05JK
MYJj31MtMVONLmdJdnwszotSEwu3wQffLCFwX/OPx1pNwOSu8yngVy3itk7CqdbD
GjeBhhtDGYCuzLdHgBPlrQTxy3SmGIkwPdi+AlDM9q1oGafCzT0XHYxJAIvsHeHB
4mtFtDSBfGL2gThJ1KbhMXNxkPfe1i5DQYPNG/fFeq2ow9namoO/1PHp2AFKjCNZ
72MDMGhIE95hus/3WyDGn81AMW5fh43ZgsoBJtsIK3V56n7G6lIbiHF8CGLK52S9
st9MbmoQjBaso4H0QYqawDluSOaEiOv1xpBVDGvme25s7M5wgmw1RqxDLoPIuoog
5WtEzKU0kszQbjGzii183Jafuq8/YjyGaOhfxRQShunSCRpMym89re6BZqXW5h4P
WFKZmzdMaTpW4HnUOVYKBsu7bASLg6+dtKSIbhOc5CG3vNm8hpvcxqfbI9Yx/W9B
s9sYisy5w6czeFDnLA8Yfb+I3AsCpLDDQSHVeNxMQxqUJ3/cFfoyRYaxMdL0l/3p
sYlO6qp8fpTx7gqzW36O/IFou4oYfA8RtYbA9z0zYrWSpwFqZgR67zGPYGIeK0FW
uvSwXA5RN4q2ycAB+vtXNz5CsYeAjFs0+4t8FF82rFwc+z+UPqmugSt9j4OpwPVZ
J2EzggYTTjNj6QNlETANy18xzvhOabs8nIjsFGzcWErlI3oNSDHJojza7B4gTal/
0nO5ZQ43SIODp9CPS74j2UMZDIPxsda+/DlH6o56hOt5kvvJrtVPvDK9mDENJYTN
qEE88IioA8rubo+fCpLzRJBbppHoDyzpR0Vtr6TdBUFnru7iU5cugTordCX01/RK
TYYP24t1VLcZbjdCHja+C6IgdyMJ0EsYgMOYJE5Hw5sBVCyKaWxXIJSJAdyMisS9
Wdpm8eNDeUt0mNqXoI9ECuXNCEwapkS+zhBUUT5YjkHb6P2EBJtcXQ3QZZebOFy3
yZj4l5XHgL9DaUTgEG1Fyr7R4d9MnrPysUghJdKqtIBwbGuA0pDgs7IQywJRvtuA
JXjA+6vDFD+m8fUb2eANFcmbPhRsjWgNhanPnz56uY0g1v77Ml/j9DpTM306i0MB
vP233zWgy0nrarf/oqI8Ut1lFEbJw25EdsrQGBWiRnqqkPf9EqgUtA0i0PgteI/2
/g0uCaZj/xuScfRUxHOA3obNrmzL4hW5WAAiD6ThTCREh6U0K5zRDfFr0Tb1FP9z
buLZFlNj2pclK1vrOLVfQLWfkb+4DYi8n8RHe5zoJzzvLxARiFoTG6bAResZDIso
5SddKHB06jFtJN349Qr30z1K1vv/u5Qif1SIPBmsUiibiPayopm2h9wZfgmCkdfN
ymstru6mbcOKU/sOwN8MRcltDMWXd02pvHvotbRb/F/TqBWe4hcrto0EH6EEXIHh
BTHie8ym1dd92RnVyxoHzLnin9LqmR8Uv0ghtdxMIKG1ZBc7TlCkG9tKznLgz+5m
pCXArBR0EJhEwBbl+A9bxPI7CZHBeA7MaQ/vignW/tT/EpYoxyiKzvnCrAkjJ8E6
UuDyUYsLZLSho5qb9CVCMh6b6YB+edIYQt8sd82wS3UiexPOD89UTWcS6GkTaADk
fhw95FFWpZPNCXQmZfP2EpRkjIoYS/UBHLqT4yxfdO1GTvFUC6c6y0QxvXZHcwOt
hV5YJK/e5Vfh9FGBfwPnJ47MHi09B2cRQGNx7zWinOOs1tWC5uXkqdk9pbm+M+pu
7aOS+Hr5XhKQODbu35+rVLW7s1QpMoK1HW/0VLJ0GhirWFvsRAPp2g1vNiiP8g+i
mQCotlHgwxLZykqC1iL2c+1FOEaHbm72PtW8aer8HfWDvlkqwfHtEC/iKzGxd0L5
cDD2SHnSH+6UfJ0iavNi+qlr/KdQkyFDQo1XFiJxp5e7CbhuOpY7WOjDaSSy8/Q6
P88w2MEIWMKShXb6zHDeg+QQbfO0yJKsoxvJQfaYOklDHf+HZmWjpYn0wlA++OgN
EzBmYsbDrUKD8qDGxXojoJh0tefJSpIH8zCFN9/QFzdZhaN++ycz0mQy8S8u6Lci
ICh4qHAyYYKUS7zVkuoZThu+cyrXrIIJsP71PDMd9CnDhwPRBpxZPOD6lQrVdbG+
O2FO3KgxZDJQsuH9vGf7LScRJmfe6b1gyl7Y1X+tXvdc2F+GJf+n5DcYyC4F2AMP
5U2Pe8sp+2/xA3u9HwXvSwYMuGAl1CTVwDgySAhRta38gJrvfocwRqrAwl4Olk4g
k4fUsI6hAwXOJ2QEyR9wydj6d+hXjkZ0020R+RvhPSfqpZwUGls8QYx2I0LIwsrj
4drslg71Gyu9WJGgR+NVeRfksaxfpM+e0FltKRMMVkFVppHv2GJhsbIqYxTYyAYG
u6Ka3Ly3NXtKTq9nD/tPkZisSlvUZmaOSln/f4gBrkRK/vDJb8nN6qsKx3bPIr2y
lMvx+ENn7mnZyRrL0dtYwhqWjLZieCfVsgmc+ZBUr0mYU1bwUv8bX4Nr4yEVP+X/
scvuffvPow80Mxn3izJvAcPf9uUHK6urSUg/rB9nwyZR3sgSDCiAHg4TAQ4ZyfA5
9zTZBIhHBYxg0wtHHEGZA1nUDCf7cjCCOkc2epttG6HEdvYQdNqvfljmsBHkCSHf
L6WBxCSAemN913WPIKYuC1aK/ClVAfuhI680Er1iuiDIdDYWiBSKVgyo7Yhmi/6/
2iPUfTOhu3BFJRDFIyxLkZ+UXianvjtiS3ltRr9GRH6QjVGwMkXmnvUjQ1Ny+LlJ
zSQd23h9chW2QPeehmmanFndLuYbEazmcisjPh3xIHMjD7aqw2NuCQYx6VvgCU4F
ylsD1oe1lOZmogUo1gk2OSh3iwmerAJDjiBypLfjkwb5nCZeyiRoOuvIonx+WPLR
fOVxdVbn/nBALL0p40jcvj0hp2Yp8KZ4YNfSYgaznk/Hh1ekFPnAi4aFVHYiU2SC
tErtc3NwJs2qm98zPe1iC/yrPJ1SsOnChS9O7Ug3WCdBdGVwbzylWChTbiIIuCt6
mdmfJhHqrByVwydckdqtOYUn0DidACxRwx5qpIQgPZDbmxOifCx0KVfXQb7ofnqz
OA+ZfDccLmLTkRV+YAZ7+Fok11+Uxaimfe6nrvV43amT00vo2rpeGJfsTUTnR9U6
xcvrOgo1W3f03xMepdglUHieuPHUAeNGTl7klBZs5yMMRkbYwkAUomhE9Rmmngbq
SXFs/9Fs3LzPV5odigWSyhw5ndoca2LmpcmsuvcNxVvcN4/90btnmnsZzUHo58g9
ywfQr+y9QIpYiR+h1rd1Dj3JNxpiyT6rvYWzulL3ik75a+OjEuA+8KHPJc3odaS4
UGILQY4S94DywL9IZ2Oi34OuuH7uu9/LovxWak9/xTn9heCKa5uTU10ED45MjCLd
f2xZ9mAwJ/REn6ZoJ/SUI7/4/Ga6DTR4qlUOu868KhbtnUHpQnDd2vbZXVSkLcSk
68UfhuuHHN45ApNFaUuaVflzteMHvgp6t2q4+fQ/Etq43F0hwGZc+4TqohZuXz4m
lDt9alC+ZgOqeDv3UkmbhaCl0mGmIQBEG8+y/1ylvd/+t3NfnvXZiqamitVRsiHv
hrswvDGlAgLc+M3H19DgpIzce9eC1h2iKdJ2QodW3I+09GJVboOXMySPFNe3mJp0
H3kmRXgV7z2l8JCQ+1IL7fntAFtnf4H2hgGQ6rqTfIxWtlTe/WYlh+HD6XKwtlBR
+kqtwMvQbPwqbvCc2J7rZXPynaDR9kU2dTANVLYegeRhOXk6AGB9tjLDFRU2im2u
PiwDEkM0I6yCLcMclG75UOymH3RvhvgWVlt0Jz49aigbzbhje8WxTpd8PAJWdfED
h7FX5tyzh9GYjDryou2+C84X4Oy8GI+ury3A2tVa5HuHE5Fpr1BqEZbAAQs+cixW
mMwJcVD9UivTIuS+TG+Dm0FUvLLRKp/F5cMrRaWEz8+8CsQ+lpMz6plRSjP9kX23
ub0eiL0oLaHdbnm1ng8dyd1Fr+g9Bd4y9/GVQuksup5zV/f+WimRWfwTvb5X+Plx
i4YQYtClyPn5nfx5cmeuWII7pdmn93wn672LuLU05ehgeINW+At3FGTwe/c/LAZv
g3LDfi29IsuYqm362M8OpQWuiGcU/DvL1z2d4WGLrepyJwnTxrJzbut2gcIyMDyV
rO5VWxpQ80tKXxe1vgfD/G2eEFTEhm6EG3ozagmZMIuKlk15G9+ibte2IhaJX9ZV
h0LPacPPMYz8BIskmLmV6mkopWdJ8Ar4yUIy2/XeuZBS7iODxlxzzZC23qXGLhQy
nFar3kBX4eF0ShuqhKnWnPyLP+7WXfePlJWRCj6t9ogtDIWA5iih653fXOxsQqgy
FV9+eNxT3wJevYWKApis1TOTKcTajIEAE7/YKGdBc9TvqpZHKhsLdOCqWIqACQmI
/Qku48b2zfKjWA9ImckGV752E+Mzx3Z6jk60MWpwskzr/4YmZDofFsLN0DYao37/
rlxAwIZJz+t3/IqvRoD1jutGtJg/EVXh2rl2IRSrycv7V9GxM1BXFm0pF1cEHx2y
aCEDvhCu3pDAjaJJiZVADsSJgRIU9u56bhftKMFU2075aMBFR9srZn/zT4x8bnxa
4XgjL4chAAXEHi1Q3O0D0zNCgDBQftBAPkRgovoYNAb0ODFJ6q0eDWSO91Y7pfQ5
4arMXSpIeHHW+rcjOEM1srC2WQ7yYMjoWUGSxXVabZ8ISgRKx53qqurwqaFVFc1i
wXpJPUNWFmpiut0rXlpm8IF4tc1cGIRX+WQeyJwTYvqeUn7/ES06fXetOvKZJke7
OvyJm+ZGZZCju0BjIT3hS0SAc2pTwjbSb/RuqJ9g0ry5coi7KATE1tXXdhOpQa1h
IKh2gb9ZeiiQWR8pQgfYx3vRFzLCD/o+OuO6eeH0w97b/9O994ck5XNzhhhod61x
TgWkgzgELPiPtA1P9tuMGhTaDZYItvh25eTLxgjdB+h7x4ESBTyMSWOBMOhutfLh
Uho6WE4Y9mIB1KTF5euHCGEckDvw2Y4XMwJKz1Pc8spQeNUJIdqbfuYQJchQmApT
KUqw51EEoBEc6Gm938dVMUet1TdkaWB5tZgc58Wyr4gLsfxv0rghIxnNSkLSkRR+
ipPQcg4W3aBMsMNAskHrHO/tvpNIBoIrpRBfs5NxNNf4r/351SfnJgiy0Rj1t28+
1BLipx5MhK/qe2sA28jJbAU3YXD8MK1sFi2wjGkHpsDg/N+0k40WvIkN5jJQaVDK
07BRKbmbL/YZGoiA9lCfAWYaLrDIe251ArMBPSDM/v9lNIACv5bucklcmr/nZjIf
AZQJPrdIRqETLtzHVaFpD9sdj/lEINH3HsxvnS0g4Lfl47oAoRdzg/0dNgql0xYM
gdA1nzR0WQI01U1uc0vwmnv1ZGO44t7rlNaTtOK8KNfeAbm5/zjArP0OtPOE3/Lm
+Eb0Px/bDnIZtQG2Lnu65O7Hp8emoJGLOsxLQsZM/ths7+virQSRSuxzlLPqamVf
W+oN5TpMVNcEx64N50R4R2oHO6fe7JrN7CQXzQJhQ9q6xruOynXib5ZCLsz3Afj9
8YTl64GZI9cyhyta2w1CYQaMED2hBOz3gc3uTHKh1P8W2CvHxg49p3nOfYWe31R3
7ghl1zhtHLg+hI8yWmQHgDdTLzaLqnb6sy5nfLwNc7n5GrPsWHC2QjO3wrTPXXzI
RSusynbziHoHFqjKsgeZNTypGHKv4y0BRZVdvWBeU096HTVYzcNvRPufg6Kn9b2O
PbicDvorf9uQQN7eKwOBA5TomcLgoq2srX8M6bHXQfQ5t+9WNdbrccTXstaQU1/H
g8phr6+hpe6zVwAeZf/qeDN1T3DvLv65JX8t+IZgeq0/0jzipD0oNrmg69CIzqCs
xSn9JNWpqDxg+/DGyi6gDfeGEPcadEkz5W6pRrcu2hvJ5T9jJXQ24MO3y0AQEKCo
9rpTCoJnHUynlWbUn3BvZv5We4LQvlIDQHdmqggKecODv5MwMBIkt7SVtn/nqeg/
7hrwuO2etAhZ5dL98+OClKNCDq/L4k+Y0CbBoQBQaU9LgDrRnd1SYFIQkOb3aU6d
Hk4QVI8HLB0H/0qDGxzIP20wUWRidWCGwMjay1JqkKsIp5EgrlygSEcmv/VQejsc
+3+Z/mpKRC5nr0sVQLEDCB3J4YQ9xP1vF4OPDwL/Q7KK/lLLm2Od6x9r8nM7zmA5
zDcEaXDdv3AWvMUeu+pHJy0ifUN8CPbf8NSW1Ux09z3uaKJ+Mc3ZzuTWsBMIGmkx
ynTkVUXKOMYX1zrb+qaNFfxl1U5F/3CliTV9giKeSwzOWZ4TAlpr5hD+kzMHEzj/
EnXF6Cmc1uiVHjYeEVVlNMCzH+EX8ssSujF3loqfLsIfA0Xw/2rt8lrMwVzQ016T
f/MAonvByccFltuSOYx9uDrhrmi6vOd+Lu5buBE/+wgkh11I+AX51nqOfQnHZeIu
PlJCkOmKzrzJ/IpftSWP9oRyYV3cFJn+AxAa1L/O4UwWjCGhJqYDpoIe3FTS/pLW
BU8jHKUxF3oje2G4bK6qiRg57GKZmnqpmmRDlVQ4NrrFirXh95hw/7KFsYZ9Y5D6
7bHFKZHPDibusZGnuaxNxG4vjUh+8X/2BO8nfRLW475lxPcWTDhFg3tX7HW0HzLm
vbLWn4bdkSPetc2vgba9ajssbZvFS6E+sVPAiy9dVcvGi5W/4Fe519y+KkAF4fAz
PtPbLum+TC2f2a/B/WdDCsUnExZr046xG46rIX++/BcRQeuhQC4bU80jHKOoWEUx
IyN0fDWbnh48kNAY31PxqTyJNMbsc0HDkqP/sw1R3CWN6/M1CWcJf8v5KNHgwoFJ
dNugbY1qmemlOIoWVF7KCB/0n5NeOQJHb8+lSpCTWo6iEV5vSVg2GSp6igPEYP+w
DqCmU/XwrOm7+iZtJBUEGmG8Z04J7WHACZToXjRFzgmAvpMMKK5i3faY3o/OKMEH
K0VFjYqWbSuhmxNG1QovFW1zAYqmu9DPd3/+zL10MQPu1qIE1gcsxDal06T9HlaE
6judWMcsIpld00olqCgPQGRLXE19Q6IX7RdsCeKDHdxpneQjnn9hxp9erSAE6JY0
cKxQdSjUEhi/rJIwDih87lj0TmWu2uiv6kegR/bTTyi3cf9IfbOt+5WIbQ7D51C+
6qSblCG3849iUsr5tU1q5v8oi65PuELebd2MVSniHT/9FNU8rjZDNwEe9Q5vGqDm
7iFBJD7JHGxID12E/7Y+tsrhNaob0O89FDo1NUEIfrFtSVx0MkNkNjB6Ax06q/bM
wg+3LmENE4xmnEFETcS6fNLxIj6eoDZwLTraUN8egv+r/034tsueBBeLE2UjAWL/
ZZYa1Hk6M4QspE8K50n75qLf2WI0uQgoyXYhvPEaODYyMioMX8YCzxof8gTfmqgH
2WI/SGPN0Qu33TZVEw/ySGDg+P2HfuTSy7P15VaCzUzOwumZK2WkzNalS19uY8rR
X9DbIjm3CMxtAPtkQ2p9Uj9NoVwaRl12u9Qw/SlEE6paV7x8Pj424P+R1RL+ARIW
MsYUKnUR0UlnQ5xx3NmSTVSK7IqP01HfDysFU80R6YLTFKAxJwWR85MFnInnrr6Y
sHUTXW5cd7tNIJ+eJ2sxfPjRk4cO1DmsDhr8XHtXBFQaGeCHifXQNj2USOJIFSRy
DeMmG780VuOJ4A0XPA+fVHXItdBhtR3xQ7+cz2Jmx2twP8TfYb21G0zJLinZXQfD
xZGamw/OSIx3s9/0E4N2mtQkaBqKPe3mzzKqAqwffyxGfyuxzZdTcXtj8Aoj9jdp
d8ROUBAsBRsBTsVoJKvo8FE26Pr5IJUUs3NE7YlJJHPnXt1AQsonXeSOJQpZ+9qO
CK6DFlvndz3MpB0gTbmmtiSZZaS0WmDeqgqaDmKtZgJvkaJy2sxApFAWTCBE5H9b
6v5nPxHMH9d95YdT8nBXMm/vY0kbZR/6L9qk5KPLeJJinG0DD2zgjqrnB2+tRH2f
pk5V9DUTd/IUZZSSpW2akIsVcqTz3g6w2lPPtUENvt8QfIEgIlQ1+bjntDRgRhTa
fpIlLFWsKc3hkLOj7ZaKwe62bMPF3lAXLIYHPbsI5eQlnMmT+EiqwAwWABm8cDv4
AxrEOQSEMpb7EwIBHL8cZP0qMXAU3UvRgDe1vaEa5czWdrEBVhYD6dmw1XKkXDoT
FjFT6TLRFc4RkKOZvVqeQUW0LH9k40q99MKwYtL8BTfNZBZhO87OwkGP026ubJLO
P6/QGKJmmyr4EOjtblPDh9Rk5+iixNIcXzC0d7LzibascKZuAI2xaq+Vw7d97Epi
7MXh2c7w75uVBFLfUmR0sbSkqkAz5n3KyzJs1gNI8iMFN9rEqDb1jVVffSpaDjOt
aOSYsU/J9iDguCCplkKlZfWVO0gvMhRVw/BGgWiKSsSG/RcWcZ1JL0/0xevdiTi4
iglmccwgpbMpekBNRvxVzW4SyJWXQnqBD3G3rrK9sNROKFvQOtNMdNa47jaN927x
GxVSD+QbkfDa6snXtnjm73I66yd0bmddF1OJvOwh1PzXlZ1ZnIg3ZroKkXlD3HXv
WzJXDC7bCF1rdiC0LQWoot4OUWazegF5sEXgJEGgUMEhRbkb9mluXijtygo16Ozo
bULYLzS+3WJOsiTrsT0dVoi+lkZ6ZMpJ7H+RDDiOVsrIHMey24GWdfdTCkAB6ULs
SiVx1YBQNxrg53J5037RSgHUxtL9Uf8T1WzacKxz9OWSiMKhkTTPy1f1sUO3DjQv
/IKJlLn53HMo9vBw5ybH9f7NDG2UH0l3Fvc8cw9nw2w5oSWWsWEMNRLKAtPc77kx
H+LlS79ew04mbgRFZcpUV0A+WlY3fHtK8zYpWHA8Xj0pmfJoLbGEJVMA8oOvKLhJ
uriUrk5xPza5SEzYu2ZzwkrAdQlddn7il61nTIfbRIzULR3RwwVZzu0XxdfKxm/y
unSK2TTrQb0P70Z9A/Ie5XYZ50W9ixHUA3xwzQVr7XnR21FvJVYDA2Y8WA5ajGM3
pFWU9tGMoijktZSBrXAZ4kt8nFBf9rg22AFMRQ47mh/H/0V8pNtwJKN4aFL4Uy6V
jSEJqbS4oUzf9SK0n+UpZB8UQeu5vWYnuREA0kflWBASyH32wdmRKinETAh4VSUX
uu0VQr+qCpsZnDrUsvrMSG2Om1DUXZXwMUlc1fYGofMy93uBQ6uBCNPvkceAV0w8
5S5ZL3NjSi9Jt45tv3vsJKjYcft+11te7m1C8YV7S+OJDEYLQDsQ7/WhNt/ctjWG
y9WgO1RFTES3qPVrjoq9vttt0T2I6R8SlUDHKX/FDu/pZdSrD3wRP/pRuLlxalh5
93n7XOXcfqz7He0wsaoSBo7wWUg5nf3/M7iBCquYZvse8A23AI6DW+4Cihbm36Qa
O+C/79VOIHgOng2xb75OrfeL2EFy0d2odHWQQ6c8G2wGgyrw/B+RB8APTUVRUZLz
SbmCvCtaEWxtrpEdfFNdFMkl1BL7kxTiKrAx2FIJtlwOkQluwFSDkwbGa98Oy2PZ
eba3KxXp5rv3NVxkCv1GsV/ggr+UVPguB/U1w0YaNsZrfybuBCnmsFM/4bArrwL3
AQZZCEAg7ZqmVWcZW95IHSQ+hdQHnWS3/eJhYGZflwYP3DwsP8q+2dyoATcVNN4s
j4a7R5VaqJJy5ogRORYIiU40ksaYYzOEJJu1N3tAzlklL82R5by6QxzPymzuSQfk
Cemof7nWnRhb354rz12w77/lQUAgEROPEcqTKHi+Z36lPHIY05HG9ExzIeT9Z51F
WVFB0vLt7q/EIr95x4cv0yqes790v5uUNpVLd+p55/Q+NxdjzNsZAWOcZ1mgmHVl
XcTt5kCKWnuqBw0XSOOQx17/Pow7XycodrC8PvVWOq0Yy8dx6IYHsVsmvWPC+NoT
c7BSjOAfSoVod6kbXML7d4VoTwCAPeEgygm/p2w+QhR6V0Q1gUxJ62Hzkyf9tsla
64cBk5x8+CccrMGb9j90MZqNyXpMAuVcJGD9gzbVnZWFydoNc3Fi7EzhNMJTALNu
baF1QJEQw0Z89SntUmX2XEZ2cMZPbpi3LyFmZk9IAyfpzSFBqtzEvWwBTaHykHJY
pNbuBF7FZwy4vtMHlZpZ9RGiPUXPyMjoaBeV698y7W/ZtzKQvBNvTS4h/dS1eDhN
vJTujfTl9FJYfL1PhaC5T5MqjtWYyxWVPo8T2cgr+DOVIpUUTs2dU6UB/LPh/+o4
dSVyhggvFGo9FQy5NOnS0QZbmN/+TR4bt7WGfS8jY5rWihbokKpGFZtY3Ao4Lz7t
Kr+mKM39Gm8xlZk3KnKzWGlNSI0Aw+PWN9D2oF2bGXvjE8MPSWMWrvfMSg7BFPal
o3D/HmffZEnrc2h0ZzwvX7zapZN0IrKn8e2nKqAFx71EEm3eIguX4WMFXndwr0vj
4d5wr39uCwE44hd2We9PYmVkeSvSlBqfb9Q1CldujdNTkR4MK9RJLufBoe/6W8kd
RkrqJ9cBsaR5gVKuekOJtwtDZcHGcJmGW+KXPUQoYE0lNKe8aXZXNfBt6qq8+iB3
87omMY5rxQBfZfwx9yDLVS4YzBMl9XbnUsei3xL+ddwXeWJh6FeEQN9/kezAOGlS
aKdu4bv0RE8IiAlUrqwQRkY6JafuTuPOWoA7pCRsAeNTnMAbaFDP7esNldaA0jAS
cZUGn+ax5ma6ZkwpIBLCQLo9QVrzVRNVwW2T/JGXSFYgEiBWEUQ9JRZ4PCwxulci
pcybcwhs/eyvouzjx9dFasajzWRdmdezIkhVenXJdmsuYS47Fo+2abYz1I5jKToj
t7Fvs62oR06XQ8ypQ01/AvNGOyZsE9gLe9f+8eaCMATY6Lodeo3zn/E06a2JJ58B
4gzPuzbsZXhx/XPr3C+9On2GErdgOVwUcWFcZOuh7vnMMrkMSvuTsaSUScXa4WWr
GZUyYVf9Uifemz05zZbcbg48Qr8BJ/vVc29/sHAEcVoka/z68ZtmbY7drwH3Wtak
ayLDv8FPUFLtbNpUy/KXqbczJxYl6ZmXZWeXBEyEbYT/6WW+bnSAjLmnMhPZ8NYb
UDT4eOlF42A+BV7gBth0UkFvPI39hrxJMSmNq1vBtrctLOTZRvFwYSrbNEjNhB7S
hTRDYIDjQPMCcwSFuiTx1qz2SbdeEq3dsHecvd9bwwojFoLy5BhLqcF6wnfAYzta
PhZIOVJ3NEly5ajCcpTFxZ1Vd+k17aTHv1925dBNAsAefx7V+21oZx6UFduTU4kC
sxxqjV14GVL+IhhL/GIkM9GC54oOkP90Vm5BSGl/ijM3t8Q8jSXeVPyL1gGuPwUw
Yrr8g6tFVYMfK9D89aOhw5tgTXV6BDs1age/2ituq2txU+3I+62JnSxdXef2NBhX
+ShR7tmkoA+3fuFE1jzsPzohkntyEYtcz1Qt4hnucjsm5L4P2n4aT0G2AYIjr6kB
5lxACMMXFD6wwq4kljohft0hL30KygOJJibW0pLcprjz6m8YAHp3K6LR1hz2uHVm
xdhcSlf0ozym0TnhoE0g17slMznnMqdU+laJfvYL9VcFLP3rcQNDAWX57kKvj72i
fUjBb9Cn8gYy0s4xbSaTiGyDaJ870zLKsoMOdgw5B2xfiJt1vLA3aEFSUEr4i0qx
mhK+ChJKPpfS/J1UXS3aSx2ScRMmKp8c+9NhmsYzobOKuhUhzYQr3FV/R65NGF0/
Dc9Ya2djbmVNPPHSRCv0Sg62rympn+WPZV+Fp1SXQyaoQwv/X+PV+OLgUXk2c+nE
vQwrCEMuHW0lJgPZbB3tTiNEjGlUoa29gjR8rqZRJzSiHDbyc7suL5DS72Sn1DPU
wIY9wMNb79y8MFs2gjszgWsWCp/q7srZJnTZvr94wTRH2kEGjjOfVczeaH/vLu/V
NEsCq3cUdMimv26WZxkFcXbxwKyHO89Ty8ZnH8av+i04giCGpM77cRLeGXwk0JHD
49/hl0b/7Qv5q4epvTtiM0o0+HG6pcRKN1VDrRfIBFISQyESrdFGaP9Xa4eT247G
Gk4pAWdHuehW0LU8bWP79Btff0iIEOSSUOMosYhKzdt6bmOlklnBOzcta4wdv/kI
HPQcuyppr+42QhjqPYWmzQ2KX9MLVAHoFbKS7V6SUR+f1CeslscGNI4PBrLacTvn
XMSl21UySCHhEPgfvSOAc9PyVIrBZC1Wy8YcOl6YEC+WXLE448xbgDVpUi8QbkoM
EFbIDZCChCNIDP8z5aZbOGwh+DJg57oiAzAXDFdCHdMzTkndzvfnr4fjWvZ8L6Dz
FOeByyhIbkG0Gm/NR0SJqlI9zP/L4WwPdxDxEIwSwFI6Ms4XWTVo7qpC9v3JodPg
DCMhTlOl5qaXdrNJIh2zGHep8sCV6bhVyQWD3zrf0doU3PeHW7XnvdSd3zgD1xx9
fx0odMsmohZGn828uN+70f4rDh9QfRzSKI3PBCeKV/yGLPhFSb6bBk7OmO07vbWc
boK6wSwwCDGdQOsyFLB6FSvgskeu3YNVD5ZEtQhxw+ImA6FyUMo/sZSGPVtKDrOL
+x3kHM1jhb1BqMrmDdiKtjahN7uGD+lyJsgKCfmNKSFc68UvItQYFfbySRG/a1wt
Mk5NFlDcwYvDuasZdt4bhqY9qcbDLkQj2ZEnLQLyge8HlWWbNiqCJ5bsHVkq4S1k
Zhl0wAWix51wcP+TvdLPOxY/SwI9LEH7qBn3uHiLsso97w6B9RHdByf4HpEj+tVQ
1pRac9xAla5LntMEEPmRc5Xh5J9SRUaov+WN6VX5FtrKTbozTaiOpg+hwbWYA0cC
PtmIawm2jY89oh6dfc9AkvS5jS8n4f4nn9nMyO87T38aAATHQfO4GspFXV58GP3q
z/ymzMbLbOZdIjUXO7Zf+KP3MEYp8PlCEY2FpwD+p/77X+D+QrfzUjsblAEKzdT4
f5JhuRXbpnfmOAhvmixlV770rGlIbUanjN79pE82yjmHRtNd0mGIwNCHXH+FSBoF
vNcdiYelkNGhUoKcAADFmpCoFEmCGMb9E4NOFK0dhXgfojyUV+0QEt3Ar8qird1y
adcWsFrSpYpqFkZ9PeyEIIwigDX2T+NpMPMUCdb1IaEUCHukEueEy6FdlbeGB762
CdV+SsMCfmP8uyN9+Dq4BGLRHimnAzEFVyPV0wKzJB1ZIHP4YkFc2mvIy+zf5pHl
9DnlkpJP4msOYxDiKKGr4btHCsVKkkN8PZP+NSW0YaoPrBKsGo/qyYS8sj8ITiB0
WVBsPCWVwjaavpXsF7s7E2pVjRMlrU9VPYyV26N4Hh1Trl/AWY0IMFeb8FpbyLAg
EiZ12vJFSeKkMyUPfuL5GqYi92BRHKcpB+NZ1VgAqLvv9oiYRvTNhiL+3jbNYQcT
hcyLUii2784OTxQxuseFKfwYAdJVXSNErB/DcMskSLGnY6cdMvmLIrQxsW+d3+5V
Uk0eW6uoRF/00o16X7DzepvQ3BuIwWGCVvbEc3oOnWYVuKX27SBL6mPfrAeGb4/M
+eFSFCWBkp9mNBDVZRSwWC00zPLXEc3Y3K9DlDt0KdGtX4Qc4KTv8pbtUdNBLMb2
rXV4zd/tkL0b9mRsZuzycNXHDHTaEicZmwPqOHNqFBTR2WUUjAP8zhBZNwntBajh
iNOD5/NrovNt5MsydJqLz8+aomVQQybl/HYs0g2ygJNLf4+W6WNV3Tq92Vcw691w
60WzubOfBEaiEOU6rOWpdMmxgvFqs3xhyLXfXqNvWy5QOIlSZfX3qCLDFvteND7F
d0NpiQurcJ2hFGhwbc/A3uIBYFk9oivSUU5xE02SyvtmFmBFfD3WGZd30GoPX3hk
COt0km7QmBJkSO7cx92coF85Egf8qA1rkjTwQhwiJj7L4noxWZLO2F5CV2Ug4pTk
zDBLqezTV5KN5l8dK0ebnmoKVfiIPzuS16WtLPN1XXSQgwyVIEXfqehqTB+O52Sz
8dQMTMV4xIpIhFtjAxJgL3DbeqHvzsAOF41SDI6IUQj9BL61cF4yjEjNSBGHlCoj
ZmpGoeSZxGmpOY3B3zFwCIOv6vka/5lm2j1MynSoCan7UsTTPrMLkjzmKs+ZMlWU
TcU+qJbF710+yx7CjU6kd0soJTOPuou13aEEjyp9h6rYqjZz9KkkiQDo4tNuz3vc
2ZLooXTzHAbkSLDQNeJon4fDA4w8c7qb7WZ/m8giE9auytVtJxaxrhBW6ox238cn
+g3wGZ1zJB55sp/g3gu+anX1d0SR2CyBk3DiQYSAcgqKFrAoAg6MPM9tT/3DHWTx
U88meM4ijPYpLD0rgEENCOdmRVcEU8W9Xw+VzuFEV/Jo2VlXzZRJJlAY/gJl4HtM
lx8zoa2+/nNNtFnOq/HTqo3rCLqC5JlISoNCZqtndHXBngy0T8E+L/GAjVEwWE84
wnsI5UeOj6YkIg11JYEB0vzYp/i3iVYjO5OSL9r1RGiW4jNwH3vErWThHwUo1wau
bUIZYI098AcSuD3xq+xrGf2v5vMzLuPPq58WbEqYfveIfJHk50NFVnCPk1gNAF6i
rqsaJPIbuPKPP9Ivz153bFuUn5wijqqEiItJhFg92LixfN+sA+KFGYR1w1Jk5O/a
eThdJbWD24IVco34aM/UN6vU8yxwp48mvDu+SGKeKvaKjOctDaaqSTwxBFRZtYmc
5L1xgvs6Z/ocZeRNWuJJ/mTXqJc5zdE07Byf3/4/KCKj22qt7zdMMSJvT7jTTm8a
sAH3uCxg9/8ECdLV1ob1MzCWVT33o5QPBd04T8ArXTwtC94KTHovVC6ynUJ9JGTa
4bljG1k1taBM7T05ZOc8vajSZChLLgJMVC90hqRLVXVdEH1ZSP38yUtz8SzRnQzp
22VRC/1EmC2hRKNn2+GAHD9UqhulteXvFuQMLzYITj51EZHX+H15byl45Ez7Gk/W
zJh3AySpCKvwGiu55J5fx94J5ym1wx6Zq/vKpYkVoH7xuAL6n5tE5ICZdFWexDaC
sIKIoXLa3JHKIfgwOVx9z0lw+vz0NORCbKB26YZFxEqbhmu8lBSXgi1xs/NjKvhs
6yLcGgp8F6wx5Gm9KtpDr9UjbjUQE2tLAz68LyqAsZW3U09SOuKtd1LQS1Ca821B
hav7QraNY7GOKj42EdYgHo00eUYG9GPRffC8csA1yhee+hmV7Hp2Z3takBy0T7SX
z2Kljle64BUrsTBNQzS/lvVl0f8KBdt8slpcaMfe49wshgnijBwzjlqodp4TYooF
DHH/QlDrJL/NLJWfOyCwdsKCQCaKA4yVexSFPRDdcu0rPYuOkt0eyq0kfa346mpT
EBgcaQl6DYjy49ClG/gmd/sTDeRDASeIQ3Wv8j/14oR53YAbXp4WTtYqxJqMxIWG
kVu19Kl6badRlqlsQ5RKyu30EvFsJJGiCoZbGM+E148KHVCUevV2Q99wM2bJmlZt
rsG7GgvYZhWHTjBdkUefjn6LyAJUlTFHq/hv8eOgWdb3CKFb3g9iVJSXVCjIo9OG
rx5ZWVcHrOxrkr1XxvQJSwydLtHcBdi2aAnGvHc+Lo6HNHe/89IED/Wx66yG2aSl
o8l9RjDQ23jublWz22Rhw1iYecXOJMwf6H0hTknzl7mYEqmiPIl8CwB5dpna3sD+
gH6YkcXz0nqN5xLQDk/AZNzWg5QqOgRof+hyriize8GDeu+mT56c5vQKBjanosjY
n25iDko3/479OuNCQPPAMqY74smo4vPn9cwaU8ujVJU+DMH7ycP3pu2dmI73joPL
g1ihsCaqwD8OPwbyiYFZA+VEZf5pYRpZxoVveYFMcnkl7jo2RxmCjOf9hH7323hS
B5ODi3md1IzPq6Lj6CxUAjWKOOyRfNvSpTzd/MJPcibECzoQ03A0EgFDYObmN1ZT
DFy6UyCZen5rdX2ZZpXsR5PmIrORQjXEgbSMLX5tQW+XxBrmHSGorYcHoFNF/K57
fWrpzsTgut/gP1CS51+INsMUxByZS9gUdCgf4McHFw+hVGJqvLaYde/J8/7hBeCm
MAbGyVYXeMMlmaAFrjuv8KiMo9E1qpqoMR1HKEMna+0Lo02k50ag5UQLcVdL5nQe
j1aSUTTdJasbFIaCuDY6l5bmVm8s6Y5ukxi8091wzD0D//9W+3V7Yvv3p7S3dFkb
3VL4v/Zlymj3UXW7Z/6VdvKzaZTqvQh31n/WstgVQOSnORN+XT2n47Hlztz2fq0w
0O4ktR3N3FtoBnhdeOmoyu+j7jFZc9j6qOc32k6TUUS3dh4bE7EMfLEID/d81OGL
mFEHRsvQ33INMyGxi+93bUcC3hd4PriNCg5CEoW7rV1eQBs5WTbZSDxxY5A5785+
fOA0Jm//1hULixljYGiVvC7QSnvZriyKj6ksfQpSpMyFBxsa3ptH5K689iKPP3Ab
Exy27NeihFLDNhpXefuT+Mr2bgndkutZQFVr+adyzt3gTOO/XyFcmwt0DougW0pr
mauvq39Iwn1HwKoZMUfrHk44Ls6c5n7JHipbPf5rbEosnhDXshdJcsBplxfMWkw2
EKEGcxLhyYFl89qPS7jDT0piN3udRqTfNWJ7ejF8BP2zZrMiJqYkV0rIHGtnUQXI
pPp++fql7UVLsvN92DZRkLPSTPEy5CB6uFOdrRrDl/Iq86hrkYx9uG2rXHzeohi1
Rcmv6liPm6UkduLnf3OuC1opZHNpI1V9eXE74Foxk3bjXfLDFNdhc/cQVwgWi2Yg
t3LEoSG3mnygCC4YGzm/C9g5pwmq7OVQ83v3ATKprteToeT7cQA2L6cChSHakxRm
ve/RV4OCVtYwEIJpH7aQuUJa5GGYH4ulog6Jqt52C9UllBKNZ6ujy+xOTjXPzQ57
LiHzySP9XU4UdJoEYNw+rwO4rH0LaGrz+oQPALwjWNJUkz4q6Za2DbiRm/kZEGjo
HKoYZbcSaMdaLruS4LNqwjqPWwvRd47L/H76li0BqnbDfXqApWqKtn59OuwHffxe
MQRmGwp/+DwdJL+ouS0KAT3HS5QtPCw0DG4pG2czL9KwAf7yi1Nk/tQWPlY462Ag
Tca0gyXPa14QWT+0GN0Z+NpKWisK9Pz5ORjnU+ekAwgj8TnbegVvIWF3AVGV6G+/
dhT2WenChuQ+2Y1wUHC5z2AQzJzb4i71odUE69afeCcgCoyo1S7Cnw7Lq+R1PgLh
ltBVbsVl9N5grNYNSpnZCjB2uYwmHwJQxMVrYCsFQZBtcCDlJQcpBuTnXNXjghxs
Clo9ISefecfI9DXZRc3VBYW6IcplzQTTe5A7pI9/pdk4iYIky9NbpdhiCTgJIBRA
CjtkPztB4By8pPDiGYD+M2uO3D3dsEGGiexyuc6TmJ7J4TnY9PKJ3KPaeaa/usSz
PWPXoTNKPXXDNNSREgNRVQmNgdcFaagSJlmL4vtHn7ph9dsoRz3blw+OOMFPt+3I
rThBAaSaNfUCasO6zgv1daU8BWGuFUxnM95LyKt4QbM6/f2EpjB39JttqPVvpD+a
yFb3htbWxOF2BOs69W8KodG25BZJ1Pfe8HR7wT4Xk9iV6yS0Izd/Qphoih2Sb8Na
AUnmms7Vl0Poc00ibK1SFej8rQONOvRgvKgqh6H1U0vuvSRnfCuSd//PyGw0T9uq
8GMFUY7sf/dGyXKadRtXBBJoGOnGp0dulHxeJ2KUsRMwt6v408VTmsQXX5fxu9wJ
Uqw++fjxii84qo7XLmKD/Ga7KsUzytK0+hksrHu04tBCkB4zugMCX1aQV0iL5Wlb
l0303dNWmeNWCivNRjlUAa1sSYEil014vNAOZnTlwXAJUhutogS4msTl/nclC8KH
96rfbhSKDBlVXgC42k/EblBOTEhwa9bO6EkaUd5s3LmGkRx9tBKlwEgcvRd4Nfi5
DknBMSbTlsHdZSxvbYFK7zxTjexuk8WG5qWsB8S1qE3fe9zLBCIR7N8/hsf1COuJ
ULLHm5R8/f+xNoerrtz+hHaxrVumoA3GKR7NUJZEv/0cHxxKk8kFtCGN19OXmV7k
eamg5PJ8+7oawb5Hu0l0dl+O9mgFCSMvyQ0JKiziPZg+ySaC3DTGWNZ1OcYsHwWZ
nsHtCRBSHUqTdZYDjqdHgX8+QI6BNTUnR1CeF5CzHpN4/nt7He54Gi7qlOeCJz1O
f+ALbQuEF29aW1icEN4l6YHmxfYK8QQZEqiz4KZ8MYVCK93oTY8V1TStDowmw1Ne
httOoIK/1TURjMcQSnWaIaqQ2G6OOg/AZozkgPWgx/07LJm6wn6TptvA/bzk//Sk
vbLwDnCxmin+iav7CimUDqJIpD8ES2s6Ny6fauaQLYbkLTkqdl5Wo7Wu0Ky8AxyP
tPjTZHSLJnGumPPKlWad0edmlJevyPmefZwYAi5DWLy4T1pn1h4hshbKbp++bIB5
9Gz8nFxw5ZafjtUMdvQqoZrN85lxlWtaHtU+o1vHFaoCVzc3yp4+8zz4OGaGcMPE
7wZmBbGR3DBwrp06YNC/xQdvmFBQGHHpiUR4LzuGD1y3QqR67aKgZidRhyBZOqBp
GaYmhINYh4u+7aOnva6DJXRt85lrsHM0CJYuEAWmqi8aFmJpT9v/DNfAaiE4NOKH
ujcsux0SvsFxSa+N2EGwv1B8Chi9g3pdbPlyoKrXSaPMOja0lvCZU2ByF23dP/xG
nv7Ga/91Bc2lM2czIkUTEMjAgMnvdC9V69ILZUfWYquucLyfvrFTulkbK/aXe7KM
nfYhpK+B0z+3mYsz5rDHuml6QhKV33g1AIm+wlKmCahC+XsIJpEnDCIgDm8ZORBw
mztqIGf3K+RUS231SfdSU4fdiRX6ncpS6PgSa3MoTPR4uC4Ejs/KvCc82xudzoTV
UvUnyoHsQtJzvXEAspRUDiWF+ZU8A/vjaeoZQn6g4mbZpKuAIj2bMsa6vd5YBM6h
G9d8PZ0oGXzNYPzBK1gr4POxkiB4DBSKaRuif6xi02LvR9p6qWaBgH+eKfzipxHQ
Spef1hD/KYsY+VrVxqgo6hvTOWi3x1eId8U9OEFd7E2nxcKDT5VRI8PjuFLsmf7e
VFQQSXn6l/GjVMizqDDbmi4uzmOYKa+wZw3DAootlcwFsMySef3ELde5nUXKpuls
rE2Y8cLF6lxd/sjDqqSW9zEALqdbijfC3vksKgctJSAwA9mNmqtAZQifz8ojhVZ5
BoaNvNZUFzrQs6uhMkImPQJWvgJlmg8Zqa2Sgq5mmFe0Y9LNCy6EbyMix95/+Klp
mG7wlUWn3zeagOUgdnae413Pi5rHKVApv5nv6DiEUwq5BPqNt7DOAhvHzNzqd/FF
Mwzy/XKbM3Uoa0Kk+HkorF2cPTb6Cily40yXGX4i2FVp7EfzlFX+2w/bH2UfrV1A
5SJdD9MMPADVMwNuzYlap0qOhtGRQHVHuHPAb2/bgKI40wPJsmsUE+Tzjmk0mC2a
OMlyFF1gQWs64+RMbk90tPxoNVu/5aovOleKvMAPC55rcgvDVf5X2NsRCA/t9R+E
q9c/NFiaWOsiNwdxwjpeapVaY36IZSkdJ71dPwSV6cWEJfmwnnTTJB2Jdmon+Tw8
sZQfZBnWQevdvzg2iiCFGl/8pNi9CVhzb7jP5M6g7SzDV/spggovyKwbERECHE9d
3R1Scd13pc8+76kA5l4G5G6896kr66q0PHe16+Ymf6iZQqMEbdE/fA0ed1/W3TJY
L8A1unbcnLOn71hrj+bTuxgKkRLWwA6A5fNln8vAOgy9s0repaRfZYSkamhujByg
K++Ddb95ebCMoFIjPygXFk1iyHU8rOiLuH8yChFRtiUwxm8F6OYd0rFBReT/Fsvc
4sdPwJxok18KjDxKDbo24h91DcJp52AohnfxVtykU0a2wM3CbZtpH0B738gB2r6I
LCG5SMTPYld7Gpd6wvNWdoOAHphwfVlVWIAehIPNHagvWYiB4+wyj1BzumNVa9fe
ndamPoZO22HT0H03Dw+iX9ZkXTMuYvhG/yedZ5d1C99Bos5dji8NeGHZHWaPekeF
GYJEuBfD6QRd/TPud/XuZBQRyjS2v4Afp/Q8HNGXpH5loQAxuZDBrIdlc/7aKPm5
X3jgpZfActAOHZ95Xqv9LpdTTXCnHw3/1vJh8FC/EJwaG4z6dj2iSBkboy/m3ORr
Wt7fHHjFrmJPJFGXBLzdhWigL0cdfLurz2rpwgg8AoUre8OEXFXS8a8iFbEtD35B
eyBZFBHWSU4UAoIRlbOqRdwr9ZJ7DxDgX+zjOw2TKbrLUWWPTEviYXZtZ1Eg2HFp
OganeqC3Z2sdw7MwzLRxvs1LhHelmtp3bL5ObbPFBMeGsF87xMPd4Uk6nkBNWK+r
zgMox9N84th4J6suMhCzmnUEtZpwAp+tQxiwKu19SXFQov1WcGr+3UXUwrl7+32g
o08VG8qW0KEzTiSXR538tGfLDc8Exy3yG5xXQw4FHToxfAI2NVXMpC1mS8jj8IPU
74iB5jjsjaCkuo2FCBsnOb1jwSlFKiA3rpjd7e8f+H0Fe3luzAdadX8ahHae3o/X
q2udG3EA+O8lQbiAb1Y1ivQHeR1Uu/xygLiq1pRLrZeQnjBSYeFUrsRNYzFQpo+j
Ak7+2s5ZI8JgJQwBloAKVygCJ2EV4fJlZiczl5k/IkGHxwp61bi52I054fYpLwAx
RyHEzvg4WaU/40J1ZGCdlyvR+BMzFmf3mnUiiP4dvbl4RipIenklaRerZ1JjPvcd
3amrqKolTiXPmOCVwfzPKFntjMBKpR2H/IED3rEpTM2pel0zoUP6sDKUMb4c6JXv
fwM0upkvFgkjJeeLGPqyHVoxtQYSLWtBcASqBmFWAGahbbWvhM3cxITPQ5BpHKL3
Jwyv/7Z4ntuik0LnpTBjSYCELXKhKivXI5AhUsFF5nVvfbZbEweknFaInr8kXgqb
q62rY+CeYeRXQ2vy/xzNuggnk9cSH70X0TsaJPpf4DcunJznYr2MI7Z27WSkMalB
XQwWeur6PiYJ0QM3dxFXk3UOB1oIAVtZcFlpEaC7E/QLMrU65kNhltN5jkmfzDL6
WkDKCMeGQ5eeLPgJ6Mk8n3cJC0bI3WBYHmeuLNm4dQWI4RANKnePX6jnHSdnRu1w
2bQKz7nL5o9UjkWX2ReD7w==
`pragma protect end_protected
