// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
diPvNF8COa273cZRi2PEwG1yseMOigrohk18pVC0BkHI0yzRNrZplCVz1ESuge7TE+i9JfO+/gi4
EITuPsKkrV4TySjYzqtm+gLJK7ujdTrD4bRtLOub8Fh57481bl5A7oU6B6eiaGGwn1uO8mDpmrRS
6Y/OyGqp52rvJsdp6wYr/3ew1zE9u2cn7d4mnAty6I02wd9jLr+ctjJvDvtdfO4TM6I/ErPJl0Ks
/Z5EelysLFMTUpBg4uL6LjojPxSQ/3nBgBrRVcSNwrDgrN81lzJs/S/NVk6UrbkfAtWT+M7bu/SC
GDeeSiQg4WoTqMnxREi2Q/XS1MM53Wwlb9POEg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 2272)
viMsrQgYYYzd94i45pAIWHv6jWfxBQGda6VGdl1IO9cKz/Hve68VA0uoHaNsrm9iurYVkA/NUsTU
twwmDaX6Bc+tHjhcYj9n2oYAlnnVSdvR3dR6MX+xRHakbnX+Yk0f2uu2mxQ9EdMQZf4Um+tsy/9a
EVbTK0WzuKf8r2uIdoR0rJtr5DcGcMiF0RLFh8dLledwwo3Q4BS7VQz6LJ2B+vfjvbOvTic7l008
IPOoSWgekC15KU0su9yI5HaGjj/9d8ei4qDw9sAX7pl2TzlKWG2Ys2uOMo5lHEY4cZ40Sbn09MQD
NHg2wdW0PmR9l66IwK4V4mt5GGdnvQi2qUZEPo5uFg9MYNJUH6XQnT9gkwQ44zDjxWYbpvh6BeeZ
n2kgaDOjnSCxA1byOM4kfe0TWk5YeiOUVJ2vck3L6mExk+xDuphfV4FWXXwd5uOSqD06ZQsX8lW4
W3tDmtlmIcOKTuNx+CemRZEpB63s9M3tGGkp4KWBEKxC4/2MyLbffz4GDmnW5I1OLilweNsxk77f
oIQJy7obEGIGBwghFTKcB2dIxd53yHic1xrzWQfATtvtbG68BiBUV460pbSFkGgDvpp1v7MBOAlT
YPD5z6o+o9m/4YnIfj6c/OBmZAr/EUTyJhryjBZDCv4AcXN98Eex9EmPJEOiZsyxDaqoedjAUsKp
0O8L1MVHJPKD3mClv6xHCl1OKiokUQdeao7k4lTeCGtOjgRCYPrceHQ1ci0brCJVQha1seWHElzg
JVfcC0qIGR+YScxN9lPIdzVMMGRk64giSCXafYs1MWo+SpiWKIV0tZYdnJw6mK25C5uTyUgpsF/+
eHSLvFF3NeTlOijRdoiVHWNPGli7OM7LX8jDTdMxEzu/U0uJD3oC0TbP7fDddO/7bo+uOgwWfLDy
jrSi3/ZIoe+GLyRi0c9fE4fUbehnUOYRIO+M5n7egObq0FRQjK2dEPsK/y15tizNQzUUxHMvJMy9
a/e2trahHAKHPNKZ70PnP/wRYncfbtSYZQbL4mh1IC2LSSbD7gnbRDAwUbbhIDwP9Yks8qaYv+f4
8jOD2R9vqqrtHeYdy+skzfxHKAMLhn1RrnxlMMF62qDFxaFq0Dmwxll8D6GMG9Eg8FJcug0tZnBk
OAFuJUsv6RJ/uueGf2G1tJZeZ00OMUhJnI3spOm/6/AX5ZUqrR4jGT+ZnxXhXUsYVf9zgq+Nn6sM
qr63cQOAV/NAdmKNXXm78Wh1M3wuzvgtIn+W+aayuKBA8JdAVTbr6PkPpflApVQwYPBBDsJIkWC/
wz+cqkW4Q2LN9Bk7aws6heY+DnCrsuIByLCmDQ5gmnfIw6PF2khCDW8/AddxJyRVftvjZFLfegHY
x1WKtT9Sw2uWrqCawvRLsh7CZ9ssK8mDvbpkk0v7g50Xy/D0o21RB8oyEboo9z34DDio8d/WX2Eh
1VsIBBkIJaiX8tsQ1/vxaPWL89l701RsI4YguKMBLQ6XbQvbH55ScjC5+ObUL3VgnXWnaNeW4ljG
0JKzvGMVYGo9wUUaVyL7zFJkbp5N+DDWuY9invakN+S5wc7vAO4Bntn4VyBH8Nwt/nr9UllCmG7i
D/Ab80rXjmyM9WF0jxsWQTZxSArfe546hvIJ9Qf0cW6WtSC88sZ4LJ7kvsb+afwmatjnO6c0oRbp
S+7LkexDJmOGFid53k3mCK3SHRiE0D1VQpAlk2imGM1iwMokxUY5rALzTVepaVnTXdSeiDaLz9lj
K2v9NJ0jERjiPlYO6miTapGGggoK2giIanEhRkCvus56L8ginnIjZyeExtSz+wm7q8WLJhE8wfHx
yKLMLosSq33ZJif/7mDH6ymqiG6dNX9sD8dWLXmz1LEkylTwHe+OEe0aeD/ZtTSRj8sw8Y4yg4Pi
PYzJ0ljD+L1BDPph3PYM+PUArMM6F+BvPHD5AwWN59mrq5BtK7BL2ot9A477OQlmN4UXTGpYMaCD
qOGRPr/3b2g2nsn++cjjT5Ek+EyjN+yDKAIaxnd+nklgJAa2ho3luMwOwJoN36LQKFpJkq27I5X5
7hqxEykoftZSzv6HiPXNQGNqiQ4XKtNqi8DNtjtYj2OqNhgMxZPjJ1JhWZvnUY9J6wcbdKB0lzP7
u9mMbbY9qtJDn8j1Li6J3VIUhkR3iaoss2d2I+SEZF3R4um4BUvoMLO1Ku2pOcLx+3RXYZsbZurq
u7Pv62zxsXj/7/ZM/6PLOqYGPm8Johwuuk53kNg6APm9nclMFk90Gmm5pNfpgMERwiY0GOQF+xll
araYzcJzpNArOD/fLjXfohAj7qExZsDWQ7FyAtAiqLHEjq/ryFtptlsV40KelGLY06Ct0JOm8idz
LREKbFDuFkllzDD8cxnylJPmymDZRGW+hGCcqzz42ZB5zWYRh8UZLug3PJUSJBxtLtWFoDqvcCCv
5bcEtjGniLd2XgBS0kCqi9vVBrI73fXO5h5p3eBL5waZTFearDaSOpFhFxL5bV+A0fjBfbMm+iBv
anZlwF1Jnqj9iKNAnjTr++51nHivK6xzF88FTAqFV3PCtYEXsPmythuV/p4J68FhFq3aUzHd9FAf
Du56X5Z9pyYmiux7G8BhadrKh9e1t309DcQj/M5xP9fPln5UXznbTij8SnvxQ4BgCm/jQXwL8jOt
4FTKBSRFQw9pYiAaVVgxfKGLncZuqnbF2Bwdgk7sZgDO24bPoqm3GkgbauVVCPDY/QbWfgb6AM1V
wGW/n8P1a19EN+CLW/v8ShxVbRlZ9A/Ml45OrVyG+MWCvWpgl5LXewwxUE7mV6E5SB/BhChDQNb1
+e8aBHUDI5AK34acJikYyb88h1UzL46eqvb9CuWm0LixHcSkwWD0RC0TQ1SHxg8TobITmqGWH/ho
8u0dE8p3l/z71zD+4e2XzNm5gPfqKLGTf+/TVuC6OTarhTfHw3Y2H4RD81OcJQNeVgjpWfscRpx4
fykFfhFdUkni66HpJR5aHkK1yky3TdvA/uHthrpNONoyeGhy09hKpRuSWm4sasz6vQ==
`pragma protect end_protected
