// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
BjU/afLy6awQGx7AIoEWPTuLHtfKBT933jCOUw0nf05MW0OBobRVkOfwRHCir3tF
OVJjAUIZL8LzfMiIJ/jc+GzLZGGT1TJGabZy/iqzSXdBRZnYiVlVmWqOA4oBgYGj
j4/m8WK6y2Bx9TfJrK1l+s71IBYpD9BaSHEOFHYbsss=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 7408 )
`pragma protect data_block
sXv+pz/WQQ+jtmwXeAPQSKthDlivFA+12Wx6fz96oEOGnzl38sp9P3q9VcJbtXgB
FiRS/CuyOZ3ARniKtCi1ct+XXCAMIRyv8VpHxStBs5NY7CHVCRrRnT/S+Y5W992Z
7ssFBLlhzUOQU4BR0455K1wbRd5u77NqmZT5Pv06/rBCQNSlLkgj9ZhVQ6E0EjyN
5Iy63jJd5uhE5QfH25DkhOD+TGZmFWi46Q3q1vykr1wFwEYOFOf+QeETPNFsCmat
ljLtM3P5hGdsmibWJ23DozkFFmV0V9iyXaGN2lfVrlZaEa079qEPp1F/+mXyIkKI
FmW45f1CeArbR26uRcYeBV+Nu5ise+8IUcv282wr9jGFYIbwrh8Bf8rABiUsq3DR
XtX8ajoM8wpLc6Kin6u9OaWlJQlRuCXxRc5NZqrf9bmTX+Dov5iwszQVTNfWwwNQ
kVxkTIdtPcD2e6s2+1AX7gjcOZALEo5VQs4jF7dKR64brzfEZNAFjw33ztvafNSU
sIx1tnsRzcvjCobCF2iIntX6o27GVK5dymkmxkN+LuQ8mSOUgPMLVBnOLlQ+CqFl
GKyI5O8Xo5FUx2CsouZTT7Y6BJpLJKxJ13jrnZyeaYSA4GWNF3vxwJZ6/kdUG1tq
agkBZpUwz38YLlB+7lql4VVgmxPteIAQeZUhoRdCujcjFjpimcJGfR+mjuDPCb2U
JXAxV8QszdvpF4l859BrVV/czGeNO1BVAh8IGWbj0VxEhX/2eovIyiHlGLO7Tdm7
4c072WkXV1OVMNycebdkqjhc99Ki+/blUcyAAMtK6xxW987AZTBHGMBloPTq4/oA
JWY9W2P1nPFdoUFm5cnqrTytp30hrwmSMELe30CcHrs05xVMDkItWcx5bNxJUxPl
VjPax+Of3BidbkJMjUwsC8Rb2K+W06nQQvbvqVVfVkVXPMoVkiSV6NFg1p7GoSNj
bk7EpCiVea5pZ5WWti7muwiw1Yw8RHh5OlzqICTRf38N50nb2qs7ETlMqsC7TAf1
7VfZ70z7TRjVUYEym6ADJ/udeH6+RYM6BkM3yqXUsyWkvHG+MKKjgj2g7nv/Jn5/
64zNR8fheQSDpsPOL42ckFqNQvqkmWExykKWeXk/9v7pF97T/fxqhkbhlqcf1mLi
Tt4zpXQIxYs4prBhGQO5eLj2bEM7z8nZaLXydipoUG3EPYwuqH5vZ2oTxFQYLvnq
D55xQHrkJrmI90zQZEx0oNsBM2V7V87KZnYMUu3X6iRiJCJxPTjVRu7VCTRkkwH2
0cBhfzCPdQWVXGr/8SmEa6kTocsBYJKl45p+kzDBnb+QD8go3WEVQ5IaCWg6XAmW
61J8Xx0rDiiyCwyQv4rGTV0aP4UvRHAQ4J+h3kE6lG7sZa6fW4Xv7rD/Q8Vm3J1j
5MGN/A0YKBsz4yYS9YxT1Aqim7p5AVb3yegg/cpt/AgGsvGxGxAptE0F/O0DKtXW
Pr/uyaD80l563WGoEAFXb8kPKhF3Ntx/5hLYf4Ou09tApZQUViOuFa39atdn4m4i
ibocm7c5SRk65g9EKjXZhnllz4oBy/eZsqNnicX4xe8Q5v5beNGLz3IVW4zewKPa
eG9TO0mjTbvZmEnmH/fqmuCZs05dWcq/8nGQB66seNb+QBsBK3CNCavJuqLWAa/V
9sLP4CqZAvhTa0a4P18wOaye8CJpuAhaSwUHRjB9lS+eoSKbNjfZ0VWLVBVj8HUS
3d8sh/bfjVfjVqSoQoRXGJ+LqGgq7jtvjUrVF03heEZviV0vgZ9TFcUEcfkgMGhB
78Yicq40U1DvMEh2Qr5xk2/hue67LkmSkblOTISyx4wWS35K4cs9fT8TyC69/b5s
MX+NF5ykE/cvE814F5j+7v1J0TBSdb+zpWjt2mMBwlpYHnFtC6jTKWDJrB9xJS/j
YGlnQ4H76F/2XEAg7sf9xHX/3ZGExk8/f38sL7payL57SoTLCRJAVlL2aRdERIXz
qFr4Hh+i0S1Z2gBgRva7JskyrNjGZ0ocZHEc/kbCYe3UrlheXGLYwGDA+OOT2kEq
tsWLstbnnYeDmNFiPIYqIo2gblGJ70utShBVIhPeCQVk+Qog1TjVkOgOalWko95l
91JTWyYMskfhpD1s8fUgOHO95Bzi8H+a82yK/EB79nCBnEgr1sjtpELxKJlgNaLo
xpS3zc/SUlcXZapdQH9I37N/ZYeX1jQXJtti339s6kneXAF8UVHYWjnE9TbNsq3A
WHa1n/z3Kq9oMRtNaHP6FRhsOKtLMV0rWG7R9BLwtNBNIuDC+OK1++vm5GhG2Ygv
xYCuicEPDQdaWYeFCR9aCJsiVvOcr5Fds8nCLcaQ/AcONxEQ8hrwBhNzLEiXczEw
YoQ/qwqzgFhZjW9Xj5SJi/UfPSTK70A6tRZvhFZKpM+BWsAocMCQ8JUxLGXMwO2m
DRtQ7oqJczTrWqmexNSFBaEA63rZHJ3jqN06vb7+RH7qBUtyLEYeUu/wZ7tHOXoZ
ikujtv3PbvdwjDLXGkTnKzd2vaJAn0G2vZ6z/GoXgrpgeWPnIypeTCv/24S/5fyR
HnsJuDyQQo/VAnTzaIDTmFa0sBTDusIxT5DyoH/y5C1wMUcWqxUuyBn/A8TZ7/0+
qdfubeeO0TXsiBhKb4N1Rcdh2XAc6bzCRfWdGIQt05DXSSQUuk/YY6CDO3FtMh4r
9hnbsbKsH0dOdy1w7QzzesncDd7Qj1opnn/4UZ5AWciJrbuXX5p7hvkw9C+Hwiup
Wevpj/5eD4lGGXii2xLi2tJQWVH+S3vSdNJOAyl/dnRzlveQcY6+r8ekSIugT8qG
ol2gOub5nIjqyyWNWw/uJ1/y+6P6QPMRLVPft+628EaqUsuIOZ7vIXk4cptXml4e
Khh8EtBbvUKsP2a7n1XlrJZgcYNVrIKGVRhpjrHOVeBk4v3ZPQWccxk8mnohVpPD
0TC0cUfijcJX75YwNl++5ak4JwULtrjqG7UfjJJzy8yCVrXJZAdrBR7B8QEBXKU4
IWAGCFcppt8SxDtqcc5U1vzaOybtZsrkQL8gT15S3D5KyQ6EzoeysSu3w+TRzTwv
IOJ2WsGSYfSL7Ga9U4CCCyxu+Z+1SIJZcU728AYA2qMEb08dPWi++88W680KsvhV
Kv+KYdNGAyfEsyvkU9GVWIOyBo1LomNj8f3sufpVU8vCZ1+9BVoqjOIy7KXrHpP8
OJB09779BTDFQTypABDLCVM/3wwoVqWSGdsxUiZQpFunCj+Cx/YEGRCA4jlIDigh
F2lNJwMVPCoKE0OIgxmjUvzXh9MHm3vQuGTBHm3Iyp7YhdCeToHE5vnVeGAFsyzs
Zhyy1L/LMQSQf+kOiUZhmVu8NA57STWoYBnzvlDBVHRiUcVToPEypQm0wW1K8oKy
GJqqbr2lZL0I8dv9Nh5a/+svQ/3awArkPTiNXldFFPLfdcEufYzH22cSYa/2MQXp
CRkTDoKO1/vXhzSD4Wdg5OwNOgm4RbFCzU2aITDf0KPgZJBKfxJFCptzjaLgej1N
IVOFJ+Vo10PkXlFEFeQfLfA1kE7WDBVhLIVE0Kz41nezKtUxEUdFz54DgGBLhE1L
bPdtlhI1SCZzs4WbfEilTNPUeHwHoN49FGAEB3DFoa1s85U2xGXmmEmAszFzno82
aRQTl8E1CIBvkzrrQwLPMmoadO4/rnnV8NZl1S2Lwmur59L9LSworQwrwnI86i6i
geZ9iGPt0/x7MGJ3JekCNrAVKjb36OO3lzt8FsoHzfgMH9MQKecFSx+aAofzCU4P
52F7jlTzGvDkr5HJ7WOcZ59UGertrNymQ+gU74j3mOzhqewEnlBKKYocMTZKIb6I
uKBrWNBLaa8deOVdxM0ZswpUcyO8Fp6Boclyox3z14YT3HDt394/8F8tw3S5PAod
LtwmAPFx2gHBpuJNXMn8RyX5TCMhB9M3OhSQsyWsjaGSXd4BmMZho2cpBbIfd8bh
xKVky9H6RRWGSpQwOEo6MyK9fd22G177/rTv70fiXP8OT+zTF12F78krxsq0ToD7
Bce/oU0QW+7x5BL/foFlopSb4XH90iNlXHQy4vVeJd8Dx00pmnWxCoDHo4sxzlkT
Kl4t7DLZMOonYRiAze6jM1P/cC0qOgkG51ITedQRA9X6vVSuvXa7vejwG0sTxZbh
gEi6y+6Rrja3e8nGTDUY3+RQQ7NXvSGgydl6DShVVi0tfvDePpR7AXJFjmOpd3L2
aAZjIa0CoMSQY2WWCg+hX/aQ7DxZ+QKjAzfSA62XMS5rAqUwM8VplFDFElln0Pd3
J0pLpmff3KtfteM1jgoBQBvA0CMytO5rzhc/iLS30f++i1PjzfJyZlU0MJwto8Sd
/HSQxYGi3f/G1Kx1aHKbMs3Cq6efR1QjwDuzq3Ft/8rbo0TDCdvEXI//P+00XGxg
uYF+hA4o+j6Zfx1jeSkgukG+CXE1KWfqTok1n3BRAjg0RwFaH+mCaQiUgPDSj9TT
4464RZllPWTIOwEkaLtzOmCmxFwAy0BRI1QTxnHqfUUr43KaqhZSadi9Zz5+vC44
152W6mBYh72Elae9XeAEzpZ2S0OC+yWsvVH4uBBNzt99Im2JrbSEQFeH0moTqFJv
n3JvZsK6yl7msTfev/yu1dG+2kRz9p3C0ZGc3FRrCd8wsSW4iqfnMZw08P5oNh8M
kl2TkfPCIFAAj9O+o3nAmHGCCleYwIqZq2ZeG8LbQW5VdtmL+g3B+NDhopP4UMYi
QRHlSo0fP+C9LrBBasf7BAtUgUkjW0pxAzZHNWsB7tdvySnhNZ3arG3bQiHLOgNL
rstT15oHkeKBYhfCFUgzeEhR/tEr+9NNTdQq0CuXo5MroVFedAVHAZdU82vcIEI3
RVC0q/7EMEQF2HL9MPIYkrHr7zVZoU/gBLv4rz55MehuKDPwptKUwqiXb1zBpfbV
LWSF7YWxWjgNDoqccify9KWg38zte+ikdKEuhdgIMlCLMIDqpTrpzwT9ZT/Re3pI
L7ZWDFKRDiUDRF0Qfsb8+d40HyYVhypxzhX6Y3Rky9SrGo6j/1oO+grDVF6V7PdF
8WdoZYNYgP4iLyryucKK3/+Ql9SkwB1lTdQlPMnVmAAEPTrByyrWxnRKh0uICLJG
Xo9qd5OYIqYQf6pIpXzWhgqKxxkT1gkZk0IzpvSUMWgPVc01awA0mhsQ0Uo2VOGK
DxmfaBcxQOdcSDtrsPYFu9KAAdHlrbAJT+Ow591Z3hjjABi91Db02/Ejda2GtfWv
RXP3CwDaZ9Ft237lWMjy/ckOhVmDZMVdiImm/b+/Q+ZxATgYBVHwE5Vc9ueSHAlh
1BsUxmSIhmgTuMShNUOY2zhqZVV3qW1fYrnM5hzAS8Fs+GlT/bP67MKK+F8TsHBH
OQIXsrj5QHuna4hK0mNNLZLi6KsWegDSx3incCOi4xe/iB7Gr60yubFlW2gWk4KI
bbtvgCBRG+jvtUnkTvFhgjAzgPmJZ7nLyRxek7PICAfO9RRz2Y1OYzHB6cRctLyC
cngaLq2iEkotxKSHDuMXuQV98t07Ka+BiiXIrdadLuKKn7Q2iX9OU9OIdS0p+73c
8aIKD7LNWSbM7oUv3jl4O5p+E85fTpHbHgKfFNPkJGH26XvcocNOdJ2Wct5PKDEP
RqBLUB3bSJZBQaq41++ld0ndA+KBGWwTWkAgh7/h0hcevL5owyGpNovM6aaAr0Ro
H8MftB9UW1y6FODCaIhCL0OHbTf+VuiMA4Uzj+15hHLd4wuLqUVN4Fl2S3SmnIrT
iIfggj9+VPr0Ck4nQGwRr+pTbbLhKuXCRVjaG3yAqHRPDV9Sf6UhghTfH1mf7kUg
EjpHP8JLgHUWJ2qEAwxtABem/O9G9wZ9jy54sPkYBxjwr6ynFQirlTxkCWAjRFiJ
3OhppTW82I4Bu2OUOn0IziVX7+S8UEzjFC29X6FQK5Au1PqXMqHS4cwBQ0vilZfC
H48DcEtc4tlSqug+lMNddG/9L/G4XpcdwUgEgPzux/hWd8O1w4JhbSKWfoIzm3mg
poEnk6GKeuSUDsdxXykaLIom9wCPkwprhkVG+8ue8+aaFoEizBi8wRQi1Dd9NRTK
rgi9Hb6C458O4omy6NaC1ZQQdR9sX1L9Rq6Z7izJk2SPjZLwyuYEAf+aVKliHzg9
nsZ7lw0pIslXugBerK6+6NNoJtY4d3oPHzlvIv2Rwq94mzTO6HUzz8s5QFQTg9Vy
NTXCkxN2X7npuyFwrzvw4hXZX+BgUChmUu05y03dwIaQDITe/C9IJPBX8o12OrX8
HJ/3OE+OxRyYNcTaSsJqoX/YR2krCsIyk4fyzqtPvEPdvjvaJd6ofDoEWMiu2T6D
V4aTFWImDzFQl7NFNEfAplSb+YzyT0jaI75iK5JOQSDWPcvGJA9bwYl+mVl3MgD0
Kg3Zbv5rUVsF08Pb/Ad/RSE7RSGcgDZYRfr5D24pfY3NsD2KauTMKGUnqNnCjTdt
CU6EbSd09ya+SVaMRBUgcrSZ0ppeT9IO21FBIIYujS8L2MX+yvSVcGNeZoBlHpRK
epNxDDMM9+rP4PMRGmt/ic3JtopgVu5F8CpDUNiK91m1ggngdf8eesIdHV8SlqnH
OkhK+VLABf+CHYANEIYckliK5LC8GltABEx1O2/pcjrm9WkPcvdi6EuqbM25knm2
Wc0JJ3YBhpP78KJsm6RSjVKHDE4qwTVRoIUgr4MA9gGEY8UsrBd+xFi7feV3J29f
lLRTIL6lVvtTrEy1qN07FfLiv5/vEVrcGZG4hTdDc1uOKreahBRcTTfohKISCbOU
cisyIZHDi2wFtMmsX7oUpfVXawVbttawEdNakD2kFqPR+sFOEIsq39gCpazRYLTj
zQD91iymv0N1VRPDZ5Sltq3h4l/MrZ1aAiyYEyNXQsQhC5rwCYtgmX1816NDzmnO
hacvyCSATeM43E10ekYNwP9XI81X1/QaBL6KjyD5bKRfrZ4PGYNlxm/5AHxDpGjn
A0upYFBxIgYR8JBOUiKGero/h84+Zv8CrS99icBmCmapIRhe41byZkZDuYucV8GJ
fmyJYYyKLS6JkEmkS1X2vq51mZZ7dBMHcb67WXnoHPtSyVbO5NnSrbs47bXn9rb/
sWV35Oczq+mv549e1BE0BSm9MyxfnGzpg989iCS4oYfGFaFUd6wT8i7av8IY54wa
q5EzlTBNFMy4GgAy7wgpJ2puODneRsDh48a0/kDsNfvHQAcsPgRGgk4UsoF7eobi
putEg8Z0R2mlivUVJwZsKCnWZOWbB1dP3y/DGGrXgUtolYjGshL3NtbFCmYZHoDj
cppC1tgWlpgpV5HPjf319+vYy1sIYrLZl+a9lLBBNtA2NY3S8WHsgFWzG4ypmI/M
+YfAjqY/lSAg7tWnw5wK7nczEM2dRaUE4bCLrdSYu/coaqlY7bqAzupKJMdxem1Q
58HNe4MvqUiv4c8LEVoSmTWrA7gH5gw3xgjMqwkXRmUDsB1ox9hT2slvggPWEnSb
xd2f9/4R3GD3SspOmVHwIu0DkuU6dBApGXbHG7RkAzd8QPllY+IcG1lKwOiSZ+CK
GbFL1wxIzAye+5DUxKlWb+AllmoDwbna/FohuKYv3cE87IJlh/0Mx2drPNZZjmou
7g/BmzvtwjnW87FUKUO7gbjgUTEAmdfwHTdE4ACzV0r9zdhmlxnWDJ21l3qBSAd9
fsjiPQlJawHfm0CzTam45lF8PG+9lJvu/k1qGWiIJfLBeubXjJsv7VZYnbYXMgfQ
m8nXTZsunzzKkAczr+sjH3DK1x67mthbIw950YpJzE+3H4qiCM2wWsWns0aJBBxq
EP5Df0sB1tM1eN0IIRxX/MjAtsPZZCG33P/fp22UtNBycmTcsZ/c0/h6LzYulS2F
WyjigfnGJFhnmBnxuZI/9J//sT6sqMzAsDRqSEhzhS3sYT3OUP1yeKd62sgY2dQQ
jt5M5I+5RSaxiZd/ADKd4veni94+y6ZpfsMRptfT+G05LneVb6QRdIFe8rcQG/+0
XFBo5O7fDsYhfs0YDcYcG+S1ZaPJVfQE4V5PDVmT+zd5n+NCaiE07D8cZSl0+LV/
s069+45WB0UKMy7SFj4FfSxqVZiU4eLyiBTwWwCeXfXfoen7miRr28gjgFrQ8jbI
p2R9q+hVApeDDcE7tC7PG8Qw6GDOGdPzeIS3UYtGCCH03LQKtSdhSuLKPw2eHuTv
TNqgOU3gFQcLmLs+w9VHdY6s5pCeNRc1TqdvEEHaANTkitpLYEjVi2fKlXM3B96I
BxQHByQ7yANFk/Cd4MR4VOSRyvsSvH3RB3/pRDFtEZ6BkXr21/dQnd8v/Xom5UXs
2eLmZa4Nh3FLkmA9HrALZaCosnp1FR2Z3rY/gs/hEE6dqmsVYUyFiz9m20yLl6J7
onUU2uUPVGNz7AeYlVGt41tJXfXT9/xnkjapmmmN5zM4XFlperxlgpknK064/W2M
95muKYRvwhfR30frNGTaJKJOb7Xzat6tGodm2GNTN2zgzyusRrSZVo/H4TOAepE5
JryC1478/Z2Nirj1TapbK0wXdJPkh2F2Ak6pk/elOeHa1ireid1jTIj4D61b/lCD
1F2CWRDhgq5gP3HEXKZTEJyIz4y7re0bY5qKmsedU0kZth2qmLEdG86xYAVw6yRL
THFmdFJ8uf+mpuifQu6uBNz0sF67PhrHSWbNEiFwJ2NN6UCBpqzdV+tlTckHF+Ul
3GXOVgz/jVEEnKjaPoT+Ni/9vIg7w+/t9kyodU3tn+RwLlHxGmz9j/YQVvHr4UQr
3iqdSJAQAa9eygaQtbpXr9GFKqrKHxReVUrx+dYYdqioaRYTPIe0r/Ie6TK5mDGt
SPoQzaGfqbsli4zwnWErQC6IfPmKp31EQWWL71RTqP5KUPDu1dVw/PcKR9adg8nP
no9Bcp7fKr0HiQjsiEQlUhKIo1Vlm7IFS4NOcx+RVQ/4wcYJyt/M+mdzqOqieBSn
2f/Xn06DQ0Rtil7CwKbHysYtCPTkQ/mo4DJY8rjcgs7rYfCfI0O38EQE+p5RF77Y
FD19RIkAZbK9XHBGYU0DWHuU5KilIHhh6ujy05VF2xKm++drseG0m1+VBjpvcQKi
aTKYiHhR5/C2bCpQdFEvmT9CHuB/XiaVK+bR8eDOCkThfq9q1piAxiXspDf8i+o0
AUajZ+UuVCJ0iP1A3C0za3tUNx1TOC6Rv/T+9tV8ZJ6CUYn4unnf//IL5aV51rBi
vUkRFnZuxU96IwGnI0kU8qDlIrD9i/10NutCEwcvUkwNnwEJu/D9lIUagXvQsykV
rm8W20YbE262oUy0wVKszkZetxcKYAcStlDJraSywqm8TEKDfPqnksQb1BO/BDn5
v6HPgbPB8rCzPP4oRp6tUfyO3vA63HElcC7syryUKepJECQZKelqdZWIqHHqobKW
oJ5BotscCsh3fxoysJIkEhPRy+aITStajo0O18dpEDTThefXC91JodfFCw8ZDb/T
A7Lgpk06qjjHNuSNqxMD2/WGbkveGGGIqd/FCaDxADNWLCOxavFG3ErEFA5Vsb+Y
gCbD4+lZ1joHuMjQtGq+LOkd/prGoMcxhGncaH9Ryig9yBSWnb/kzRNDA6aTCble
B9Xyfn+1XEB6PyoYspFq3iUfHUL6zBjAe+VPyWQt/h0+eOmN6bY5xvaZ74MlnLsr
QMI71yKJQsTJ7mBBrbCRGxaa8aSY3FEo+B9LUNxfFjXVet9ZdpecRUA6GQ0EUP16
ttCuc1dIh5Ukaqqa8TMGFwpL4luDBHDqlv0ZUeS2GB/6Pp2FdpKOPng8/9dEibpL
DbkvGkdL2y2aTKYYoZc9rs1ycYeFyNO5GKLkeKrgWEwIsdhuq5Oy426iQAXILGnd
kb9bXSXhvZuAuUsVjgMH/g==

`pragma protect end_protected
