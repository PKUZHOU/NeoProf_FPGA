// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
WoSOytLnsp1ZYmQLh8soZLqosDbEaCSKo28IfTS8jhU6t3nBj8nHjuP4ibe/tkQ6
ot9OyV9/DyvCcmNu0AuSdFlOu4NHDqLnRJwRr6yIis6eWdR967RAmHl0Q8Hyh3RS
WbCxJX3RHluiUhmSJ/ZxJA8rb2Nom3P6uDoE82qdxsg=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 93024 )
`pragma protect data_block
9cj31HSZLrA8APbu9JimBfTFaApqYKVzvUlY82DL3BrhjfBjVr1hYSWIMxOG8EjP
f17JQ+CcAFFfOgiLpiv6Ym/sjg5iaRi1UCRweZNgBso9Sj7OVU4wa28jf8VHIqgR
xxL5Gdm7dYF9xiBZhqlhxTPL+AXYZolf6vkxZm+7qzwR8eYVXo4JVK/ypHzrZTl5
UE90DQ4fg9rW1ch+RauY6r4ct6CX9VyrCF8spiyqjWdaQoIiNFNSfzUjeKA9oPxe
Byrl0AYyZgW9bM5fDK6WlyjyNTLuAEgSi4Oz/T0HBK3xITKuraqRLs5nJGeE294d
JSKLkUeLGrOEjio/lT0u7e75JvjQ/Ekw0yER09UvOHGzexZPCXZbKUMtlLhceWoe
4NyU+9yqRm1nwfl7iBOnc+IH7w0t7DxnMUU7dlp/eGJnQVufbqUMhNyBE3X1JSTz
KBe1rsVKRzfRLbZGEhHyLARZzpbR0s4xEX4/arkpQY6+V2KTARtS3DeAWQtFekir
1IwvjPUbyg2xzHi3S6kW1rNh0dcg0uFOJ5lPGW2B8rQMW4Fi0UtX1E32Jbt82kNP
25cR9NiS20a7dBes0TCnmIqxjPpZhqo6gorTu8ic0Yoa7WuOn/COVuLQUT0YajIO
ZiTyMYWJ3hqxqpHs+ckZFw6nZwUkuz9+zcrSlIsmi00diaqn+0IszMxBn15lGMXX
NAB0rVjmfXoDChfvXqApx52/YByq/FTfFXce5dEIPXlsIMfRTlSKXu+C0Y0D/LVt
1DrB+dLPhp1JFw6LMy66yv3tlfqg/AEE3SwDDNpLirisOoT+bvldz+JuQWMtp9Au
+Bf+XxsJfCtqF/ogfbFzYQ/LuKgEN9cyl8qOrVWc5ghpiBXhqz8T0hRlUmNzEocq
r96nridEJrArnR5XWGN/KnAdqA7wCDIbrQbagT5ek23Dr9idJaGXsfhsfBY4xklS
dk0o2B8gmwv1YLGVt3xHpOVKvEewNyvoxEkGAh9U0ctszFyyeX4aklqRPgZBTSJv
cTFqHAhvhEg6rLXSgS39wcc4xsM3LyBJfF5f+Ot8tbra1M7/51fvFyn8nWsneYmr
mNysmg5bOsTdRgfeccbisw5J7aaNXQyAiaVOfs4gWiCD8T9zA/CR9QonP9IWNN6p
8lxiruwYZOLe9Krmp+6zdrkohphjzj9mMNf5bNAyvWb1rd/b49VIG6rtDkr/jOLJ
YH7dCDSB0D71s+QtV/d4l0EZUk3QpnFEgprGKQR4D89d3Wo/xDAgPRgAp3sh0+Au
v1bKlRzLuKdg0GVG+xHv8Mph3E9rRLn9UCOV5u8cFIJkSYxqp8SlwipxE+HgYduE
98RNWkk7sesiNQWIMrLY4tEpm/rtulSfn+MKQ78cXMKLQ35ZWNIMB6Sc2ZghIR/u
1sI9+7+2Ar5tHUAayoJAcNgnjEz1r2iei2KLy07x8m/Bfw9bxbtFXwlnFBQCVGRx
o2kZMhmUYEb/bPHNjPilkyz470z9CTzsJccXVc2ARRfWJfair24nLtqJz7UPZCr8
vp18asKuP41U4ykcJL7gSL9kn6SOxWJWvqlK+JQNxvFpUWEEYml2duOF0EcGvJr8
Dk2lT59/NoychRVQyFV9qFwdWv6WVJJM8sMIXJjJ8ZAJYylFWn8os4ivsFyneWCj
e3Ts4sZLygV5AB0Cdu3Uex1k410fJ6PhGUcqeQITLY/JEhNwTF7EZFtO/KNXbpNd
F8UZss8YpEOr4PPheATjodbJ/TtlM9RI2TPRCPMTBqzSXXDpUsXeJCubZ/PeY+9z
79rrp0lvxwcFhMCkzmBps5Ml+fuzWzwCuB970mEPvZyhQfwHs85Wmskj9kveLdsR
WDL7DnU4zw4wtT01f1hwm4rG+KMxU8Pq8uAy3ZnFLt9fgitHwmFrasttDAzmZOog
sjzwj2KIfSJyWlrTaGmOqWYYtXNH7SkR2w5mtyMEvpOZT2nge26xNUrSGVWRHkv8
w2Mf4ogAwyFwIvrA4Yam76yAioGXwb+d5IgD5Tfzt7skxBKOub/3rNdkLovJKENd
wvyFkDQ6eKCP1iJvMkVrksFMpaV1d0wPOpmyFmqMza9lvoUxjcewNRebfcLz1M13
PC50IZ0jN6dylELb7nYotcCt51lqmtb/0cgx/PBD7i4oQ13uBQhvG9nlo/jfcsZ7
XtLFG3OaM1rG6tSIo3RAjKTEQEDbeanR9wb7tak/Qd5qM54MQEKtNRwuTXsXv8sG
lsA3RRc1FuGBY3XVNfAEMQRPfXvc5A/xARQ7EWogFQ6lpwmXno9XQ8v+BjWE7WU8
iVHc4slguhyToVn++xQ7AVbCGZqQ2rqjEDAHVQ2EExew3YD2S+NIdRqDJykhp++n
kehyY3tm1OGb4i2X58/J010O3DxwmmMzaeR3cd6P1AGDjSlcRC8px5+XMwtonFdT
TFh5LfNef/fP1MWoFs4pTdmLo0sF1vdr2KgRz5BwYc9uBULs/KounPOqi6xGa0Ld
+qqZa5fTUUU/fV3tDlzOMZzAddvWL+L8soSK4OzTGAmGYmxAN/u4X4+TQ4qEh3RK
XX7VfbN409HUyiLnj0XcCBFZp3NP2j+KZmHrKTb+8u1mZjtQ4JwwFn5bK0jB5Sxb
ihZ+KJiDo+zVp44b7Y2uF+3oRBppK3+4ddNxrRrw5Kz4MgBEdOL0GhRJWeuozNfm
OYcObu6IaiXwpXgoaDV8hQwnbHxZT7IYC4985+R/yBGVw/Vq2rl5K2lFlH93Iw06
ooKP80ySD7P6gtuTzKO7//qEmu7CJdSHSZlAbgptWVTt/xMGacUEE+yonthfgaAV
Ud8iiH4HnOjrSJzOg1M+Wpc9ugrwb6lRc7hhmaxhkVIYaKbpKg9GEC4+3GOp0O9P
OMmtKaA//tSHGvzWVaNiRwoA/hcPPdjCy7VrpxWmPaOgg82JIH3por0GdmMWtJKA
uNWAaQKuVaAoY3swUIi5SmfBpz1z6OMQURRA5M2ixScS70+X9jgz5dsAazVZmtL2
kfIhuBxDDJT9ojBvHGglr8fLzh8zDb65WJK6REV1w76M4EmyL9rbmwJUuF4Aw0Ee
Xxk06CW+vkJYIyijpqFmCN0PRZJi67qyu0cS5S/kIQlnMNRZVAESnqCMmhoTKeA5
10jpA7JUZ5rhQTlwIaP5pz4O4d+SsV7vSVsUkVnStBWEmp5WqbwkN8dwdn3EYd93
QDzn66ZJa52x6/5gjQ2Reh2qlvtK9uqKGg/2edl6Yd0q4sm3AbgzGBRBVnFgzXxC
TL6uckmEbW7PBvI43Vg/KBlShKvIZe5pidI0U1cGE2dNj74BtLOHOGOVyA2MI0d0
R6+KMfa2b14/Zu5i6qm6YDjPfxqLbpJ0akgt0H5afK+EK0qIA3SFUcT6akTRT1BL
C/ZIv4ng+TLUkhvCOqFe7tRd9WU9gndb4wRnYo/Zvldrz55l9P9mLW5UvwT0G19o
XEtpMVzbpKDphCmC1t2qWcis+FrLwFfvA1LJtAxB/PLsLMcdNMh91xBd8b5+uXHu
QHX5aQGEI86YHzF/j76HJHEJkzJX2rYi1ioXGKjGR3dOzt+ikChAMEWTe14jhvwb
JAQB1oMKfDPo+6whOWLKHM/P/b3bsSZd1cw0QFpGeD1e4LuenYh50o3V/6k7mPBJ
qCY3BNSC1DvymQi5lpElp+h8UHC/VAejK5naWmhKWMGHXtPEwp0Ja/bB95kqQzAB
lk7enPOWFJ2gtLZE8JboJ634isLscTtroneXvwfl7sQ1Uo5eprmytwmOYlvo6wni
5UcC1/tCqD+42fUz0399XFF8NPAdvBvlXsiMJiO9T72m34A1XRdKaxcFZp3P2KJE
E0h83NHDKuorCqKpL869dMP96D3KrDYLHvRPPq0uEQb8O0pnUTMT77zaVopHi0RC
Ph+xgUMHbDTycFUnlEMB7U387ID5ncV6PM8ZxhO16GEgydR0qmo3oiOlrjjnYZvz
zFZknyf8TZjkiUopEdMfwVytWstajzZQ8xmFrJUuQt/XX/JT+kKJkQTo37PPmjF7
8cz25tFdlz6SLjTjXvAcIUMfgqoWZ+3Vy9OeWtcAAodRfD0yW0tYd+9P/tFLUG4S
aPVtt6kAifzg+PMsa7c87SOt1k8RaE9Da+GRqIBkhbrxv/+61LAa6ZLEjilrQqvM
FLcXvPgl70BE5OLo1eO7ZEV3Cdo9yQ9eOr7kr7k/RgChs7h2GSQs38iIFzL++C45
T+liImAA2J1x4Pibp/c4JL0881jmOC6QP1tdG1yBazLqIHtfOJdBOqJkAu9OIepg
Qse3SoOypuveabUpNIQED9xTZGc4pgUTBrWavBO8gTFZl/0qrDT6e54c9DcwMLOV
lsjj4u74Bn8CKWqbt+PdSojEkIaE3Bb1jttGHoDzavXr9bjxJSzyPv8P+v+LIpWh
uzt9VRKlM4+qXhaz83QmBlvlsJ8aqXi2DHmRwAUBlQvkhlD2ZrCGjK0zY/l4BRZH
nGJ2tPGjPYL3U9gTS1lqj0ApJUa38YowvANbEzDjJe4wYD4ymhGcNyviwdNhFq4L
2QIjJtQyUFrXB3yMyQs22KrnJyFdRFbvOat/Srfc6PhdEQb+w2eurchEYVLI1+xl
afixIXlWxypAMl3DRbZ/x+AU8vzTIghT2XjLCsIzNx86b4S5g0qfVmrf8S1EDt/z
EF6Q81mOd0QwRL02DwFLdjx5QswKbC7XMTMOj1AsliFea5FNa4k5KQqNVf20NyXt
hSgh7xxolI0K7a4gTe2Atle+Om8B/dUOTnM7qfpSfpIswqaEWEb3WFpHDU2BzU0/
bQdYT3tNmwGADau8PluB02Pz5CMSJjvpyHkwctvRoaBRap4ZT2NVczWwpmeVv5wP
qfA50bdokOoNCNIa/koi2rC4NHThkbFYzT1q7Bx4mPTbzgx06f74uwayrpf5ADrv
E3rVHZhc+WdeUCnNNQPcSR/bhOGFkFQgaSYAQEVsFjzdfwq50GAcn/UwKKBUr78K
7FFb4fi+t5rjCAWnEyIbMnTV0eEUdtE6FAs4oHvtMTjdCZToeFbyuzEakujQpR7r
tTuF1BDFJmkZn8+nT19asU6pGNsb4dSSzqvJqETC+2zSlYliig1iDgXMjiE7RrQy
7gyDjuDWqQ705i67bsonNVn3+7bglL458Cy7rqyAT0qxMIHz5T9Jg88UCGA112Ah
+WVG41+a+x7ZdMuHgzqE3rkOVMkJZgcNQxqDjvp/1uU329d+/Xfv+HdoQM2vUG3v
fyFmaq61duetyBo+teycQ5OZb/8lXWB95FWGuEdQ0/SCW65U/tA3R0/MNgtC7GwF
sskj9AwtZwcxwzSNmCXsKqN3iejVMhwBsHAel3vXPVerSw+mBvJs2/18ocUnYI0R
98MneioAL0RG309whhRVIb1R5AFFFzCQ3kgBymkuk6CFbbqK+44WzW+TYGGseX3O
xCbHYk2NAXLr6gm/MEfRqBcdDRU9D2xxrur1nYhsUV4X3sr2f0Io09w8VRN0vnlD
2I6ip3YuPQHkZh88kVra99fxXHNgBTm1jDD72V70PCyggp08+QFc3h8ozs/+0aaf
eVcvnEZdUREnnKQ8rPZYDxUuG9qe6pk1X1qq6aH1EHKY5r3w1JIB2yjoj4sVOVfz
6+A/Kx3ZomDmfNabq7jVWt21+e4228y6YkoWc3pyoWDT7qbeYpTtwWB6bPuGzjxt
gXTayGfodCpSPX+YKt/Q9YLuFQL74mgjP40uVUsEM+3cLIEbfA6Wl0RsfT2BjOkG
+XUakct7gYKhkmQH/9o/sbfQuKWJUEZy5pqEke12MG6FuoJZtGBxAFBpXY9zCZC8
VTPTuFqCSE8EzS25+Nxha4KFtBsA/uj+4NaqWlxfkOAMVudAZVQf91hdGbI1tFDo
9uZ964qVqMClw5u8hxmwvcl5jtkSIroVSd3yGVZvC6iriwsfVlBFNbFwgsQXQOUd
qgZqOrHp3yiZqWtk/6Q7gaP5Y8Dug7my3eC2jCzli6OBNhC1MUgV9sgr0XTwi6LN
3hm+rDKSad3RNjPs4A5jtmk2YzcldYTKN4DqvQGxaJYx7JxsQpn7I3bxmgFIwD8j
esJPq2Qrt+xMPZnBvLEoB9vQibTfLWmL3Of8Wo8lAN9qgRNPNFne10EN4J4w0TeL
ifpfWDlhof0vI2sAdlu38MSMcOVAFkl1tqo53MDKWCylzSDCglHhj0Ih4JRLtZt2
C7+mt2bDJAWAa3NTbpgRReyJXBQba4gnE+eAq8ly3wXSLJzkNGo6UsBFHk0/yZLF
+OWXOdtlYjdAdlJw7Xv/AkYh9l5hlT6C5X3uc2iYzheF/po/x7mw8T+Cys1IYP2j
edJBNJozcdLsWXNFx52yxCo6mW+ZHJ2n8QsVz+MpfuoDBEYYRIM83rjSHjWCqlWF
xJ10TnQ8uifvx9Qx7Wy/0+olhFFoUAQmEi9QN5zcumHxn8JBgjollvHvSuuUe7Q3
tv2jQGUK9avwS8Cg9LK1RMHyalB75pyFK3D/35PeBhjWd9e2U4Zui3/zW7TtwLYT
eXq3Iqz9rnuEO5HEY/sg5DlZCVMjL1/Q8LtPzK4WtfzxDRaKsnDU+PXUa+jnxSvE
hez/LSgk7jJS+zEWpa7HYeFLfywyxIXHx0YaQG0hm4aOsUK1wc8AVmkkZVlQtBec
scloWEcZp2FLNndNql0XH9brehbPvDCDdbHdNQEx5VtSXGSssxZZkmWpPL80otnN
NDJ9fyK04cUitWmXedCxVzaM8pAIP7FpMpe9qjy5f8cxAhhRcvcUeh8EBHaYUM5Q
5fd4TrfTRVpQZDiXA44fn76ouZ35WzZJ1ZqvZlURzB/ajjGEa4rHCZ7beT82uJ0l
u6gDyMfVjCVdAzJEX/svnW9FbD3tjzaynqbTpyqyVuSG0Y0dSPod5H2QNiVUIdn2
Lk/pp6QbjTk6LtM3K7Jv2MeH7qA6m3wYgmVGVZRv/G7BzcaocJPFedEek+/s71Cy
1dQlHBECAr1pCiG97qn21jqpYjAopaPnzMpeR1jefQOQ8m5okl7TNsP6vjUXMUSw
4zBe6lmiw2+5AlwAX2NCkBYZDAIkIXSa2wwQAG5l5fIw8m3Cf6Ya8UeJv05ipcOR
ooslr7T2br3xcM09sGRunDxETh/B+bT7o5/NSSKraOExcFhc4hYEe59rzpeAtNQi
3h2cJAtq7lAlJDRt9FdTwSuY6gIivZis0mEygygmm98UJxwMvReRsV7OVV250mh7
cya8yjKKMJ2VRqUl5pirzhI8W1KlAg0l5APg8mbmJ0+waL3v0qNKlHeiUOktukh2
IMMrfswWaC3uA12FuGswbkUQlBqDbRX1YkoZilb2ADa+dqUxmnwvPa9gNu5Nh2n0
5BNcGmd1iHYrYGiNrtHbdgdUvitUPc9m8aP9sxhQZeS7Yb/bN8M7TTmDTZ6Dmk2N
K6CcWxDGYXd1sINF9N5v7XoJi5+TDocHF7Kfz2RlIWRuSHf89+mtgGx6GsTeQ3LK
DePY+yVXVIJ1PNBb1NjyinXC3+B9K/cEpYp3EUhgkfQmlebDgJYQXgqDOubZKfCX
V3Y7hXcSMk0RiYogsW4SE+pH6oNRXQlqFoDU6UwLUvV3nDkWa1+ZmDfOx1akIALZ
0WuxzhZm70NX2BKb4LeB9fZbwvdkL3nJdmQ43V0IOmK/ZwArsqH/ok6Pe28MxtI4
Mb+lFdK+kATvfd9cLwISVQEi26Q/gUa0W8HtYPVKgXod3rFzajMntiQkR5d8OouR
yqJaDROErqH2Bb6sIeoSX6Ld/RUJiztt5NypBm00G2LKDqYmAlEPWB+sj2EpwYaR
XE5687TYT4L9/UEQW/IxwJgARLQjN0gq80xqpukST7O3RT0F0Sx9IZuulaoyCuI7
9NYlbOFTc2VS8o4hnjFNNnf+jRVMfCPoPWV635Dqr4sjPUk5WFM0hjeTnAFhgn9f
fy1tSnukNz6ahTkojxBb87qtFf/U85T2wBfCh9HCuW4U5ioG5CH19HLRCTJz7ISe
ySIsEtqaDzuh8M0qgnIKy4q4ti/ayj4OifKxTkMUDX4uP7xH1GIRANB7NO3UIzuH
f/MBwTfyeR3jR82io43TX4nATuOT22Fy2q6Tp6WkrD7fpBnoS9u17miC2UfkBukK
GrTowE4Gr8QUyMbIwZA8LKPz9IyeSdbrBr8T+KOsctTG9Krn9xoDmpdt6knOMQCo
Hog1+y78Lk4XpBSHgw8upZE0EnRFWHe20PvLhxY4fImw0zmGM2B1qs4e0YSAbkPb
3FMRB2HuPIj/G/Jb2uYSyGfqeoSc3HXDGQgg0UHh00uSIzSQ09AYikTKPUEGiBNl
+rF97vHHHsDPNMu3ZpitNVsNWulfEwt9H89lY9OA48784MCrdiRmBfQ12SWi+L1k
vCX2Fn7Kp5VE7N0hSFpnXPlJ6GKc2UI2ZxuB8WPcRi5SzEm2a4YxGAiCGxepAPJc
uzrHg05hYUeCs/NoS+Q+2fn1k/J6IKCSgJDk/XcbOczBuSHpcigkkz/wiX2FZYJU
rb+CPusw4YUmXL/kd+AxONjpD/SVJpLdnjz8ZXuB67JU5j6+YEwVJ6blLmvzgQhf
/oo29jkb0peF6F7woaJtPgKubbPoP4yGs0GayxtMt5/v66yZuCbCMWvOuB80rDkR
Ye8I4HMgIz618jsKRNfDkOrzfg6zJuVVFpt6OEIeyfsX+J1AIjQraru/kFPaSJZm
/+heJPhrdZ1JtOWnhklRW0B0hoZlWkloXkiwzVlP/JC/c+HPqO9viZl1JFSwnaqg
wGq4vkGJhdGoi1wUflKOuww9ZcNYseb9iOq9Q/uy280C1Sb91tINZxQBFHXU2ZN5
puFvJlvIZ6xFmCNrN36BwosBZMm/nP63yaGrm1CYAW3cxqtzhpeGXY/TPevyy+mR
KBAUZWojgRlqaHfQmdFUJfg0H2C3frkogw2vFSgcuAM81M2t0as+BtwnRt2Fey80
oqL8Bx9LzAHmvtMooZZOJDM3ywto2XXchY9z3xOyRMUd33WtqhhM9umiuRGI91h/
xsV1iaIOj8GMnPvB1WyN66D9/nsXr8gfjIXtisfcTK3LtWkwZlh/cmzUjowM3ive
MH626ZbEtYA5D6Dtrwnv/MoT/1SUBOx5Kl3FQlSAcx67M3ZAgpUtYE/YsMAV/8uv
FfetaBrgk2WjY9EaZM5yf+cKdk0L/QSE+mJdOpPgwOGCgw+7NA/rVoDQMMY4k47v
qPl8GGZ2tM4uQxw6Clorc7v/MOt4RkaMOCMu5GrRVyNC0an3D+cztXrXP640bgSR
q7RSBekFTBxQu6PBQlckWNez8KdPjgPYYXTCTuxFYcMkcSBNXsoTMlIFypq/8SaO
PhlBXJ1+R0vVx2l8awyXrk/KyRcAdW+M+XelGUWWE/Q6YsjW2MiizvhWO54iAzg0
zxC2i6IxmuRmesDA99YGfYVamAwERONdk/EfB4iB3hUOU+YWLz6JUwGlFkN7BsnN
25PkIVh1bP9UWbGgxJd/w783d/yv1FeWnqA3W4iShqfQEf+lNpbz+B/4TSMhRWiq
jZGBMvg/ucgJliMYcabeNYkM4ep5gElgslgiQhaAnRCG2/6JBFNFv9rAhEs4MtJd
T5nnDNtyHknMZz3kbCXZp8bfybuNTbVNN0bbi3S498p96yf70FDVWtExyoziqT7u
h9Y6vxWPYiGrblXKMoXtpHWsAOQS6wpsKfLPPF59/AlPDCnq70nw4zWFMSFSF48r
mYDaltCnxLwR5eiMv1HD+AR3XwGGwF6evnS1Bww/0OKRSMeYER2EKC043bsoOLrR
r6fSutc+sZLsMvZLtxszlODQxnIp9deFTTiKCywqNr4231+KIlcgNaQsZvO2UU1M
914u6iE5htAsSx3YSzseYjDnNneZPG1xoFNVmW0X6meu29DpbFj9r5KhFQkpzat+
yV2EhXE3W7ZFjVBkXdC3vqGjQMLo3m9MXDaCHqzT1mPFd1TO9/2MFW7DRu+iAsy/
ukPYvbLneGi6jeev9mVxGuGvxBvmVH5szBJZugkc1A5w/Q5/OeTIvaFpluloEdfP
oRY/1RiJuV1WNowQnmGgz7Y0tmfLahZpXWJHv1n06t3WkavzEJoRYhniC21wt5FN
k9ohYeLkVFqEBZd0BvFoq1JAs8wLAVSa523o6TQMgwOZwnPLvqp9yrfKmqR+BWVV
28Rw5jy1PWsdTnGK13nhggaNvBYnrjk3+Impt6oKW0+EInR5im3zeYl5qDcB4p+/
4eZzjTAR9560IBj78CXVVQLyNlsKdI4mNfBVzGNNWSvZfP7E+hzIJo0oraM7KNql
04zc1ubV+LYrp/uqiJ+GVVBUq1wZwQNQipqGAvzgQjOj3v7KTnch72L1Mvr/rdL6
2de/WhCAUHUqvwzy2b4KzN6QbXWuKaDs3xxFTYRlgSwgNmsyUtCdWdCOFL1+w+Lz
gDtAkEbgeanuQHVBw8Rt8Vfoc189KjP+NMP/YXnXabXTlVV1TqmtDx9HLsq1v5oh
3olStiVB4ijBrglPHTS7i7+qlIQORKO2QArWdZVAQx+SqvefwLvLOpkHujA3ZGg5
UexjAHCxGOfDyXkqTrapHu0iDksmJp7Yl1VAOkQtw/A6UfzTR3q6v0fr2shgNaGP
+i1ta04JKQNVkvieN3Sc445jc2uB/n6rtquUvaDVqPzMKeLfkP5sEjJ5fXZhBKcJ
VTYLkt+T3dWrWU2py60R/oU4n6EvpSihG7etoVwf8zGHtpNo2hufjZMeV1a5OeAz
8wSAm4ab3JoNAjbIpwihULXnVQGwQlDxsjW4jSfw7z9lsDMmpC9sF3e8xXI9HCQf
4cGNf+5+AaZ2QV2yltoxwIRnRfOywBfhm926Mg6xP1DQ2NV5k9boLvYN7vQ7MYYP
hAjZIvpvFBGCPW2JgsnHxy9FGXUT49aiNr/3kjKH81slvgDQ6yju3sTsChNlFWir
v2NDu+W8HhTqy/tzh0+Z4SLlnqZ8XvxnowiPKAHzcaUs+zKFbh20zvPONnevKfJ2
N4KAccvaILLmZcDcpbxhHUjfLQJBcO6Kv717gdJfBmS7VGcYMIGjOcOMWWUmGmoY
Dbd8VHW5LTP348cXjK5F7Pv+xNOM7v7tnxRVlV5iiitFaqAZF/FQ1+jvxbemZUto
hjyKNIaoi+C1vOizilL2xhI2fLC6nZM6vUcv/TkN6nraSK+mvLGAxdTRZ4VmTn5l
EbwLHh9uX5QvJTeH+KagsU2b1ovIGYJazTGdpqR1Mk8rgFWftvmOwDh372eCgbBu
aHho4G+u9pGgQ2n65qNjrQTdZFOwMu0euOEKM0Jt4KAA8DVWo2d7OFwtyGdGxE6T
YSBTiFSTaWKdPd0OvJFmelZmPSvpZmuBxQHHa/RkxEO+hoNB7/qailsDN5MKbr0q
iyM8AC/4DMzhIuMRdWBwVLeExtznqTEVaxMo66ZtH5gCbJcBy0AT4drwKeAcu8RZ
233GS0J5nPV6SImhhPeGwBUOXbej+KaBYdH3bBaTu6/guj3cK1vrfuWtSLtsS80M
qIsmOepY+ef0f6gm5y4p/hit8tDXJUfcU587+gwKAZEtF5rR3I5eJRxj3xUbRWi7
0TemT5z6tVuMAZX7AwKrPEzP40lQ49zoRGis5B+8YohpaULybsHrU81sZ/3Gi4DM
SJJiDhSKEW+NczJzftvMO8UOvT1Eb5pXT5OoF1BySOpZ2HfK6efNoazpgIxELKgs
UwvV2P/p99rxqLpfG9mO2nK5/8JAypDev+IoPZKPAyxl3DOAkA1GHJXx+nSB8DPz
AVYzZPV9CkHfyFBYd8iSymdp60sry8pB//3VLsPsks6PZW4siubUok4qS2cMjQfW
k6QJE6nnsHcnxshLklpk2M/wdhdA/4lG0DPHTWJgD5uT9YiCQjJzRvojsMGKFJHc
S3nvozW8s7MZayloeVcZA+myUGX1AQfjxnSWkuKlVt2ecVmxtRe4c1zl9RoghNjA
rm30YWcL5BNpW78H4i/CKjAoyT9ELw5BJ2pqeWrnHRl3DwsYcNyjisdenMF0B/7d
EnSAjj1BPrctBWgr7OrSjOA6G3+1w29JsSxvlLuJYkpdteGVRDwxpylTnYYsf1Nr
GeiXK/okR+jalUD0++4OyBNn6Y24Iy4GlaX0V70npfMVAo5xBk1BCUsxUo8TQOHL
ukwb+zipNF+bImXJAZK1FUQJbEi6iwLMQdtUFIVesZfkZJIWCMIFUE4351wreROI
gpTu8r8LY9iRbI8YYioSe7rMY5d1YrPQtIF5l/aKr2EWiFYP/781zu99/Ax6xrVq
LNUFEJCrxYaUDao7HDQgXzBdryhiNL3/5Ly12hPHDUtYv1ZWd0zu9OrjZADlHxwB
/e0QmND0ass4FzouLkbsUhgZUgbagJWUQyOa+9gESVDjn/n3o2DV57+EPg28zJIx
aVvZSWOoVudGQ3/uKH+mwDHuMFdNy+/KhuEutvMy6WpPBDCBRgVuIkhFoX2cg3oP
iVLpGEBOnoFudKemGjngtTRM3Xj3WI4jGmZNiAY20//UsVfv+XPravJqTfkhNHWQ
Xj5FegQmiQXfXc9mWuSyBYAz1J2qOD9iXWjbqZFg7dszHXigtVkg3ussm1iZz7ft
ee4nO46i6NyfpW4ygUcGMjPcEh/CHjOwmLsPKPDXje0ERGCpqJKuq1kD7e8YyNJ4
//Dn7VcqRLPow+rukUvrAKrC4EVWKD6wLeRyIh43F6giRfpd2Yc0VoSaA9qESxbd
OZSf1PeAykxDlsMCGatXcCB4/cZ8W+R4BZy5U/hPtiZ4sdMkX8+1oaSfppNWOdYM
UbiEAGhFKxe0oqkVPLO+LCrfFBcwRONd442flYuE2WiwpEANY6NwWhphC4LbKPyJ
ANb9WXFjcluTKdpWlRShFpT9X8KnURFZAp0uis00AcxCNkIJzCUavXczWj0AFgvH
1pDDMRppP3flROS2bKMviXCW4Zv6wv+gbAbf+6f7jwVWONUzd64HP1njUyHB09vE
4Mk7D1KNQwxZrJbDMsLIzgJ4J2TGQEHpTVXVKtL+ToRKdd+sgjhR/PaRSHixv/Zg
A3xaX+ZPZPUH5VEAgSHOIKEHvt3OpvzrmgDRb5a0liAJudMs2ROSTHiA52AbJIXC
Z08yk7INff09gFwmH6JL9XSqfo9hY4PAAI71XkZ1o4/c7y3fbmeqG4vKaXawfuJp
Mxt1yeocemZj0kcDJklyEJJRFzFHjgeNruedFWs085buJrK2wc/24V7Vp4XgkrUp
ToxP4kc5XeccxtwODv+O5PpNisr+f91HfmTe9CRCTObnDGOIS9WoN7GNfZIZiBx3
2CtjBhodVD58Tt3z4cUxMQIpNKa4Mc5T2KqJnjDvqkKGxhZolcLi5kjrUVlIFZB5
MB/yZpiy25Gf3LkMIdlH07xJJvvlmgraaBkoAflZoayqcfILAaeiwPjSQzE7r4oT
IjNzC5dqDWYgdVN08eyQawHmVghQ1kdC9mQZpFcMhJWBBiL1H7zVHjmVfKtlO5Ig
Go1ReP1nvt3WkeH5bXUfz5iNnYAsTps+Kp6TOiPXG/isUjeMrtWGdJgGGTcFQqQm
NyAzC9UmVJZyJ5Jcl1asAu6RaOUBXYLt8hG80uOTM3smb1xUY94iud90y4s2lRyM
/aaIL6gIdpQnx92Npk/79s3PMYb8VYB+0a15+e3/5C5fFxT4opjqO6UbtLupqhAd
OG7JShG/HEvxoaI8VhmwduiLMTTtIjSqpdBE68FvigXnSa2jPyonPtz4DljmwvPT
OB6Z8aWDv+0I/jIaffRgd4jcxr34Ne34fUK+fpjWxwzTwLocpqj7dCo9J9DoyUz6
2TGwHFFRcGVe61GxIZVNI5dPcm/dQpyKSDfP+qja1C0JBD8/fkPWrsu9dtbb7Sl6
ZcKtLGIngKqbjhjRkGX+4ytPJDLV+lHBIENdq9dB7TPXvMkB2q9jatDFrd/VvLdj
o4LVK/uFRKfU94fieBB4lbLiWuJwC+9jenRSNYg55vhwwSq6eMrDScer/sHRz4XL
p57BXu5q7hnVY3rosmyNdCbxowZIQBBa+VBmVnjfSprcuRJZR1vzeSlfNie9TDT9
rbkOP5IMvHBwowGE3Uybyq/xtomz4gc/ZfEFI/y7oac3x9xH1t4n/yrYD+p7xcm4
3iCvFq2OXEOEIH5PwZ/BoBSRFvEv7ibRXlwwwXkMSvWhOjEzhBUvTRjCKP0r9T8D
G71JVLDTOnMUBx0DDo/oe4F5lxARCD429VY1M3pM/t9VmiFZ1CQJqlcKfGRwLM+M
rJmxCTTONbt9rIbgh8lDoLgFwZ7TbnW3OKx3m/iLJi5dR/5blZm7Ecx48K+ISjOg
Wqyi2zCldHTEhvAwsNu49MUIcaLidXZK4NrWlKf0NuIT7StCyJTsb1/qWIh5JL8z
STveLDIRysctSudBjk0oe5BcSlmT5oK7fTtEexD2lN8TaMjDihZxhtjDkoXxY9Hs
kM29OkKGl1HQDVHlzqFksargEAUCIGRzmd13tobAFUlTkW7rRsJnRZaA3vUmsWK9
+1PvL2KAArTzF+O2yTAl1W7uZyTjdy+THGgj0KcfiKVVckE/bQxqlwOJSgP6cytc
SUZr6Mpq7h7cfkWTiCWnOYQKuwsM5yadTMqAByS8jzdPsHqEG+ez2whU00xb0ptr
jRmuSlHSZgvk1THbSYY49nUaVch05e7EctpBWKawnSfGJV1Nufymc96TkP1HENn2
no4dH8D9x0R9Pmjk4THqJ/uZ1XuSHhFSbQz3M3EAk+H2QF1PhnPYvWTMwxHKj820
Zy9n240YmWH7zMfH5DwvnYN+9wMoIQSVpe5iXq3aefmIciqbCl/ijsfNUEHi0Pdb
XzpKfwPXArMXJuoH7OOWsFMgh+ouqF7HeZ1AIeZNkDr1CEf59zfuZnIj29TvhJ8I
R8ZYppNyIAMLs/m3wg64B9DV9PIDBxUxa5GHZL7tgPkJBfeRzKSUznfr+FzllLLq
rGsq8yMwsx0UdmkVYGLifTokNwmR9PUO7GryIU0kIYABi3EaeQBb9zr16iUKGyrp
Ew/TVG8BiAFqOgW8265zBO4o2H0LlXLnGrsVdE9QCj1k1IgAeVbxUnigZckuUUju
3cQmnya9cGSnyrAtWOhR/3p/+aS0YZBQVp1pQF3NuprpzcpunxIr/ScgpRBizaNi
4jfMv6ZrCCAu5uj14b7OfQEdiw7jVLvNODrUgmAz1/LSVTQ3TxFIaUEs1gAXdlVD
KZQUpM7iOqsFp8pkqudP+lhZVjFovu4ZCGrgvKad0oo9CVBSvwnpuKRz4XXNETv8
Wua/jyR3WaHdkqLZ0Qf6nJGZoBGQ4W3rW3Gaym1lrcr/Nl29+3rwgLMsgrkEoM2O
X6ISv8Sg/0eNeaZbaP9yMFYEZYJq7HIZQdsS7gZpSvlMo26kVtzrcpCk/TIY+eO8
0zeTIcrvkiwwgp9A2x6TGlCJnBI2EdMi5uJowfLSt3ZedFuw2zQzdXQfp2588/zE
LxUYby44OrlajokbvPXEztvvPIoJQi7eeHW4GKLi2Ewd+RrQjL+naBpCqgelW9CR
0x460QkC80PeAeYCjlbr2q08RgUyyt70knQ0B8ZY/mCtYMCDbZEhSWHpqKISItNh
V55pwbyLx9wVT7fRMIpa3SCStL1De+aRadPBQJeHOG0kPZI6Mh8I/qDA7IqdIqgO
MWSW7u8+Wj4AQEqjzTnWWJJ3H2h3JTlV9E7zCraezm/T//XR6fYAHEggmE51TGQ7
P53nVGqGNn13vOuDwChkhVueNRsizLIW5koaLtqI7OMV2VkOO6Q+aCOMdBAtNp6h
VI6fJdDlTwwX1MhRQfMe6e0jkcW0rdJgCRwo38UjT6OVi7jyvXlqqdrTNNaD1S6q
UrouaTJwTdbVfXmD/I5lQHbJfxOsFO6POdIrg03R5yUauSbsl1DOBQ7CizP28D+x
bx0N6fPApEjlob6hZ7BPFfwBXIe/v8oPp3EyoIvG9r7vNKMp6U8HoFml5F+z6DnX
tl07ZJv3yW2USgF1Qm+Yhdy+fc1jX6kFj1TbTvCOmRkiev08pV8ZLOp1C+7TkqM+
pLNF0E4ksoMw460qSbGRuURBy20NePghjOBYh4MuZoXcVBri6U20mD1jJ8vgn0FY
tP1Df3EgjVRGc8TmmCoIRBaTtOqBkfJ/EgGoCjZL39SFyC3bE4420emBMQctj74E
XgdawisUTAu06e9ixh7KXt57OWR+gFAskSHQQe7IaO21e9kvn2ZYOYUSZ4bP5Qbe
NiSIPEgJECmNAnE2jfN7crFENhhOT84uX2Nqvbkq8EPgjSK4wIyngr9cCq8RFRcT
abCiaDIGEooec2OWx2wmGiL4osLSijwgtC/Btf9Y+Ckz4oy9ULCMCqKwCSO9sRiB
GXGoXSXjNZu0wrk/OIijVLtlQV9apR+zRmDrzVkoA8tlwh8x7UsKzgL9iWUML6jd
bXBjkLy4rw3lJmwfE0WAeM/duU5WBbHZFA3HjPBAZTcejc7crVAPGAj/wO/UpKCn
N9cJO4NXJRERIwBhrcNdO7UaT7olW/9cB55VwoRdeI9ZsEQxLOyBBDS+FAnNXW72
P3W+NJY9LZRRVjF4SVLxwGh9jQ2NqitLR2CsV576B5QCDoiNu1qB1CAOikg4EXdU
BJ60EDV3GiZjWPm9xMfO/MW9d2mJqNsUbfiiuuesp/2Qx3waCMEJwEquPIfgFpgq
TPuAclmKZtxWpLHbwIeeyzL+oDiMd80CqjPQimt25YwqApss2OHvHAvciMDOWdXy
dTcWn+q7JcQbgwNY4MBKALN5UyYaTJHWvEfCnYetg44kG2+o3MtS/4jp2CX1F9ex
WCwxXEu1L3CKcGD/hsJ5m4bLIgrLVz+1B8arG1zDQ6vAdykvc+1y+6SZv5eR1hen
YMbkCM2+8fydrDUZB8nw7keDNQB3EzdcuuSlYsJvVxcM3oF7qcFmAq3fRUVW/5U9
0SD4bbPqVSHJiQU7WP+YrgWWznrTpK7fUQJfaRRL+bBDmJl4G50WKnasetpWOPql
d1z6x+OCTeY/piouDXNWGLE5gr9EfpzYRqjtqGalgPD/8oe75gvxTT1yQNEUOTVT
4rzXd1YDNIOHI75AWlDCdVNfYezxswDP4enY5YlX2tSBqHYsyBdrozFYokBReYso
K7rVb5M0UWBqS+FCxIC9DhsB1gtwqbzUb5DOKXDPuyZW0p+F5HXRTL8i3hb4Z63L
62nhaeMeZcZ49rkEhuHs8y3VjfcG4LQtJixODHYicOCiLjPkyo8h+b++Wx5DxKAt
mtZxudjHnwGKoXmIwcDeNNpMAqI16RRzDzpOAl0/lNpoxIUP/BUfCx4k7T0Dq8AZ
dh9rUCr2o6/DrVKg5HhBhdmYh0X/U98eFkEH2I5x4qXiSSmKsPOV1X0rDbvpY+gR
nmcHu6t5ELFe3GYi2J/xw/TnHDg3jY9gx3P9dv884eNLLeAp13PJ8XyymR8diTh6
xeKxMqSYg45lv9Wph5np3P8pfaGt/az7hvXtVeuxORaQilNZzmvjoJ41FAPrfdda
iD2lRpPzeJ1y9fLB+T49E6KIoXiV0sUL1EHRG8pyfxnDvVZKM4BRyfOpj8J5x3MT
Thx8UxwIo+NQ712bDprRVSMAHm4R7G8Nx8cHVjI/HNMrJLtv+S3q6zw0RuRgbkru
cx+7A12SicKziDpZzUA76+LzXsKzXhmb+fNPPj48fE/R0EY+c+B1A6uDOmBcmoGo
n3Z3UsEc/5t8GTTaNXIjJg+gzJ6HMyWauyBQMtM2NNhH6W7W60inttT4bU7T0kTy
jb4PP+6McNQaozPCFWBMaS40k0j6srRnMST6tXZJ6G6EWwsazxXDSN+7SBMDWxTa
8OzYV3H7N41oU0UZ6GdT6T4qAUkd/M1x7f0l7cChE9KCUTejSkoR9gKuD8DsVWsG
oLB9GmU8pIVze7IjdnY/0rmVREJW35CQjA/DN5uW21XViLnbeQePVC2kO+MlO921
yGJOcNvE4AyOc78z3N8ECoPNPZ29qamIqNvSZC86ZUXAdiAzgzZ3uorpAvrYEKDb
6b9oRu++46ky7RJnWTG8YjtnLQorq1I5QAA1d1JWvE9JGYjdlyD4HlNgymqx02T2
kEWCsemdnyFqJgD84SSFsnMiVoLWOzFXIgJOppOnfqFaB2+Nsjv5lhO9JXxMmI9+
fn6sxRhmHVrtaA4I1u3YVxAwsoeriFvPGn2Q2eT+EYv0qOoY8MrN+nNHhOpfmo3s
D3YEjpc6bmP0V+Wgo2pT1vFV7dkfiQkYt/CraOlzjKJpvrmSDWNXCM7NULDyTeXm
9Z1qPeZ//WK+lDlDfzmxTxVbxWozmjdRi6UMWb0RivMKEDd+tNuklcz/teCpouuE
VSg13NkQqRG4b+apBA6Z57xx1/eUOMiP8Pgnm4wzv3r64tANT1tl7u6YXMJxWnmO
h6cO5+EPrVsNGF/HijgYVcr1+xSYBJWNrGjoQTiCV2j0TpOccYA/poIHnrgD2smK
3M8V/MwrsMEMmfjACtq/gYkct0oFHMeJGqR61Lg7PbpTEGzUxOHQ/bv+sBWQsWlp
QMiC2Ek4maR3IVs9xADj9cUnWs6QrNui0IJSkngkHjTYzt6g/Oj2OtgFnqQqv1x9
3cFAeUTNVxzXEGBTkHBfyoh6hpqrgkXRShrxukeS15YvzcrwjP1Jx6LaOVMBYG0T
U6Lay1UmZcQSvTvMeAZx7RirRAUk0qkYUK0zoWwKzArbrvcvQ09a3SttaYtQwtKw
fWFUJOZyhzjV742XswRS106PJ1GraVtHWcfjG0BZo0pnF4gYYWGGVBW4SvDgO6wG
FHyalRV7A8wX+DKpmo37In7uMkL2T1jqtgNTHab6uhSPNMFO3D8AghqMn0Z/kbGM
K6N0tTaMZBW073UIDsj0J/PfqZL1RwFV+PrloS0TBXZ486dT2SJeT24pj1VWDEpj
6+zdDFYjFpO/MmGfu9WWtJ76qLiiVWLaY2dJ3lAiUJpo2snj5TSw5Uu2kwrRMen6
Xjpp0r8q92YPR5p5dc/kWhQ77s64W6dM+XDjh8rMhGl481f2EBxiuYuupppJoarJ
GjwUEYK8IES7jonQazpi6igZ/PiyNVEhbZkRIfgFIkFwlAdyHFx4APGCrkTjD9Og
XvXasARoGWDe0jsWQi6DxlmBudXEu57eVp/vETTWzRvXrp2M2qEYFtspxWMuab9Q
kZDUEHZmvL85fm5k0HILPeF4LLcjEanVOs2bTG8Nddilb/+TJmS5mDHTSHkQ9X1K
TFMabl8IScpJk10p/oOks5S2Kvsfem1m2zDbrP12RuA4JFcNEtIpgKPTdr3fp8he
yrmC/Wz+OmUcG5Rtqqztds90F7NWYnSlGOSu8vLYoMiINr/XHt7My7jZcQmH1v15
Y5nzA/jKDDfGCfwKzgqiMhWN1cBy52Cy3r/8dyEzDqy7pzAIky7aeNSm0mbawuKM
yXee56L4JHe0ItqafIyKsY90FQMZiBzR1SxvXnTzTPbOVoaDoe+nxgNTUq3i+qP9
eiLQdPuKd0CH06Weqhq+v1HUrpITInYkAqRLO/Ih5J51XL9QQ4pLdCoZ+TnPlG41
KVhWyz/KOXHvQeIT3zZp0VfzKbiyulGATbAjhe+QDKW+miHcrPlof7fyM5d7fcGm
3PELFJtigEZKVfsqBdjK0Rtv3jsncX883pELiEpYtDZPXA6/KPPqBAA7xSVhQMO4
Ew36I5L2p9LHL0GqJ4IYCpCRvRcLnE+ywRy4HuQ1hc5Fk4f05MIjTsb9QZ+mSKWT
D5X2Dtw0KCkazdbYcTpTucZfyYAjwLAVD5z2louKkdjU1i7DpgkncdqOS6oximgc
RQaEGfqHYFqzJ5wW21ofKa30UiJjMysWsDppO7SC5GlD9BPWGtPDxCrt6Pq25ZtI
uVlkeLhGC5Y6namEEUuukJAilnRSwtpwbbARwvWb2JvtNCvzlKSctm6n9rVgvUDJ
pxU0Lyhci7+HNriFlzD0Kik/7sX0TOvJf8yDgsnq6fFSVkpcUcLPJOLXCx0W59Le
8UeRZvmb1RDtkDOSEPMyXS6vVJ5FIC9GSjHF0nX6WbM5owoojHMoEbjWtGwxiN+e
JejHQLcVyk0NQHt8KtbbtZneoXHUj91hPVHl6y+bXLDeL/Zd3F5Lx83CidroAA5h
K1a1hgbWHKdzlm/vqs0VibpIvCXoTZZNHbMXmml8+J+9B2G3oM/PSjTcU5oN0ET3
66OIKAcGQ/BPDEzYtK0587hMAfw+VZvWPedpYEqLCl9LCRuSsYkiDtZRaqbjozrE
94qX0H86wDbPTiR3gBwXGcW+fRG3rv1mWA1wAWrAid7iWUBPRvW7lsj0yJO7XExr
xzeNzi8I95Q95T1g5yofA2HDVxMsiuPCUFkXSrYchoqEUFHGlM9mFbqMFxUIFsF0
F4pq2MxB/aar6Tkic47c85igr+0NP+CNnmgMUIftID9lu4XMgIMnYBqorAbi0dQ2
qQi3TAFF3RZqlu5oTNGFg3lgBAihZvnED/yfrkN3uXhaGR1SmdsGpnvC+Ut83rQ3
kstGQATanHnIJhyARQwFn/Lq2584dE2aiMGybHBh1xZCCymOcla/yM4aMpyE91ps
VkaGi4OPROo5hcFlYWWMx/mc3CqJLPLViK3aDVN08z8E4SWBWW+gjz1FzgCzyW3u
bj0tViAFQcRlgGSCVV7KIVZIYzcwDuD/1qSrJMHx7H/HzIm5/pXXloKD8qxCZ5Ds
aSrktPk3p/rZOHOpQ7gaJ/YI/Dw6HLjlXGwavVKxXLLx8CHacbccJod60lYhQ0o0
oJoVLccVFfXIdaouptkvYC3TK7tDNHlMeMBeNQaXF4wckolATUqzUX/N4bC199Kf
kwliVLDzzMjBdcaAJcJY42KPexO/N6X34tA6L+U2er2w25N+v+adZWXUTopWrfZc
3n4a9TNHuoLu22cUTao7c06TfwpNIRXUAH01M39CHjbPQH5NE/GiVGKBim+fH742
HsxReik2KT9/goTYb+7hqK+Vv6NbuME+tj2xC3qZnYjQeFY49PJtjI85f3oPmsJP
HbV3gq2A1jp5/gbkN6MykOJRWyTOOv1CxkId4WD4MyxWMddXT7K/9AO8/uW3nhf7
IV2vVfCiKS/ykek1/0TFZVAs44VEwkQOWZFNBF0QI6ddejk0HNdOyLgnE5jSCHgt
SJBQkJkmc+yZ9tQeCt5dkCFIqYhsbWaigXUnW6eV6n5xhuRpxSWRMoUJLWA9q7aK
BmyLrTMykr69xUBtg/8NTk268alTV26xvUx3/3koqXiwN7EGmaZYmEuk2OG2ShWh
nbke1RN+0SzF/zvzU/BcQ9vP/jxRqpIPCHoC8xaVpYVlMFOLcD6Vb7Yc/sKh5y16
TaguVU1ehPE/QOTT2D9xJSa+4+OmkUjHlfETBrk0F7irBh335zHV2XPz4WOGgDn3
yIwaiGbqWHPe7bQDv1zf0e8psBQQQNFWLdXuLeFXfo6jZd8A+HWrafECejHC89l1
Lzs4SqVIO67HandnwgUMt5Ys+NmZiYGk3ppGoi7/E272P/eoZOzQawreX8tBlmYv
3/S+6r1zWZN3z70wUD1mRLkf2OlZE0bhkKHIwD/257G+t/YfY7mjAxmIvAjW+6QX
EKH/CbKC0OdHkAPcBomsMNc5agigGeFxDkc1Smy5ah/ilwIKO2smIxKsxqVx9+Ta
yPA6umeE8l8pF6VzTVSvyFU9cT+BRkQNqVxzkP4Ub9qVSE/1uX3XE9VCTucZDcDR
uLwN5wXBZruU9IWrS3bEDzly7LmYCcCIjpazTSfmqZkAZPLtZVdwKMcL73aMaPN4
8JIrebvdRNal9VdHXVljVyYGzKGZAlAyVl8vK1B8RkiN1Nxb25sXb2qwSOzmmcy0
tAJcLiroA6plpNQ0Lv78KdP1L6r5YeFvXiQzh0MCxxU2YEXiD1D5htJ5CK3Kc9aI
WMzmmzzHT3iLdAO3IWA7/EQGrtY7OSOxwbAPgiZ4oJnqkWNL260yhPSrfWczBKyA
I+aXORMqfQ8kgGM2xtEEB/Gj14zLMxFZzfBwTpHHVHQPA9o02nY2yd96+8WMRqxy
xJDAE2PSTdbnZkCuF/ZRb+s31vsEbvpFuvuFcRWeuK8ZVxhDFm82YQF3Gd2iH85i
3Yj+zOhbfE2yjUAT+dG2oCCYrDkk5N/0TDQL5R6HHazXWoM52+ZkK5Ul8QxelmmI
vN/4mbvid8gXD91D3FLIDWNUa2mIvOffwti5KxaoKHyGov7BywXFoviqsDrpZlTj
BUJMug4MPEzb56cwDKyQ6BfiVh4mk25R63OBv4XS5la7uNfp6z+Q+Lcnd8ufUy9p
jUrRjWwfBoyas/P+9LzTUCix2oaGe8hAZaYhsk/FgJrG8Xc9f9i7Ip+IdJJRdg6n
9gdnPKkveWKEeZh4BeoxiZN2XVePQS38UDozySnWculLz6zidDLPh79HDYzFSLUg
SAvDAnQWyCtZsdjoONFZzzsFgGrAV+Q5lO33w/cW1I4jYGubNargwbL0hE99a9gy
v4CB/xS4/7F9u1pDrPGq29Nu1D6mjNrzA2oFvRzbgqwskwMu4o0o5JSHwFCftihV
syPlhO0ab5NDyIEzqPrrFDCtuJQ2iCdG/4+yoQpWVSwZFAqbOEHZZuixlxzdOuLS
UWf+A3GGSk2zXbo1fgoMPXLF82ZLcfhF74UFIHKBmjXJVZsgtvRHQDEf67hkEoJk
7VkegskCM7X+SS3Z6BzyotGNiIzzIzikn4i3Q9QqwoF8qFROqrt0RksjPoZ7mDnP
ul5slY8rkXHgXbhKkGjeAWABhTmSiCsJLlDiQ3cxdJ3zbsUJBMLmxlioVehHvjzt
q5DqnadUoGBXb9W9mFNfs9OubuFvron31aUTr96ABoaF4BASUu4VOyojLlf1K9bS
P+4G+4OJBXlnSYOCUlbhgzqmOZYkR7qOSkybv4jZylr+s5L4BF4PhftM5AbMlV9Q
4+wLmBjQSF9CGz6bIs9CEgP5USmnOGByyQh9GYa4PBp/8ulC2YBs5gSehmaM1PCj
waH00HOIagnx1lCgVAxgG7Knphu1oe2hNgNE4FANqa6zf0KiGoNXEvR1FLhBkm50
8lqNQK4Mh19b6gDOk9ckSy0Gb7IuHjEzx3kqLQB1m0dODfYFlYkZOFVYF37MtPbR
fD1c+iua9uqyoV2Vi1D2pnqnS2lgs0WraQukZJmhaQ/v+FTVFC5cvg+Y8UquyIH5
zyJKUN191/RhhFIA3n1bIhdkV0IRWnip8LpGiSqvUQQc8a4RH25pBcfZVehVQ7so
u51+Q57Mk1MKwxdx9+YrYBKcwwkI6AnasMkDV14KQl7Vg5LYmlgO70dDeyGFWbiZ
3fRZAGjgrFXjvRat7lqs84QUWt8YbufzXUjgjstuviM0aewxqRO9LZ5Ojd7ENona
T2izKpAa1MaWpsWp7OhjKBdDlpUOXKGUbxIyubf4+WuP75lg0HYDobxYwB896RaG
yN20fgAdBIzS2VUfHMY6Z6GtBtuPqqBzx8N8ULjPHutOsGy233dTESGVWA/3RTkT
cLDPXQ0ua3GuZi71FTmt/oqQBHdxBbMuRQhQvy8GpYjk1E2ZbjkipAjMx+CZ2+B3
KgQu3eDlbBROomWPWME9mRjWS5dnaT+u8Wnm0cUzh/5uNxLUhlqwfs1o+fd4ZY0i
eeQ4Qnt7v3XRwTqKg/RgUY98TTPPtOyVI1IjntRY4LePh+k2u52ZB+O+zgzeo4QN
TYfXLCkNrGMkt4jWE+xAAUTlowx6X2hYfBqaBy0B28cLhnKYkreyCH/K5697+FU7
D+6nx/V2S3A4xyvEtMRKcyrcusDnW8FvUKQJxW+XLp19awkg7i0+dVvQm5rJZs30
7zhXbjxArH4YxbJOLolvcElIy5+WWXcAetvwN6btSOQvuSxjwKyQbm3ygn7vlh1x
XEvPZfAlQf9FHrtom6exOLGmv8y5tZpDyaviXHjLsAaOzwv/8U8QgUtzZT6KeAc6
DuuhYZq71y1au8ia88SKPwvmQs00WazVZqHmVEvOm58zNuWBBrvXZlBgbo/3YjUl
yWjbgwHyS1duJzMjL65S3qwqErwor1pJ3JQNcOaOW911wDyNx2Iy3BpwULsJGD9x
go3HxoS1A68bfBvwTsmDW4Qgu5JDxJ/YOs+CQ1Fbdy0IqpJP0c5widYvj3q5HUF0
CaI8mjmcKy1vrR/xnF5LxpDZQjYzyqFvLBuYRq4+mn+4KRVfpJtGAzLngRqvmNfD
S1XhXemOzXkLOqvJY94/zzSiE6T4OWj6tzPh17WIXKTluXzzFQxSU8rVSANjf38o
sX8jlm9olwWq2wukP3V1gkFKTQN+XZIc7nD638Z0vRurIUwiXh8uiICOplwlnSw1
wuUbwj+Wwz/u+/OrOwgb85YiSy2lh+EDS+jUxmbdxvjnNq/a0Q/eov+UiKafo2Y5
kJcmSgO+djSlMmY5C0je0tnj8nuBN3nXGvZFQ31ymilwEsOReUfhNezelcDcakS5
5I+w1nSdaGkF9lAywJ0ews0prJbJrc/dTTVuLzrjU1HSx7WwPJh0cFZQD+OsWP15
Qha6O/BIKZ3bcsUfP98G75cEGyRSM/bwz6CLfk51VOJG0lxStBOCg/izewaGxw7R
zFPyVQrLyvwC1jL+3nvJVm6k/RwGvhqS8ZBSr6YIvGnF6npW2mpsg1PJIXvnqIwB
G0zqhzTHUSlXctcaKssrR+7pDxblKT5Phd9xoiHwf9fU3ZWu3todj9yVP1OJV6Z4
9UPGEcrpfixXQxOL/gjDcZ3aSGFkUALlr5kLM89VC41C2aRInJRmwnStiGEPFt7O
cZ9PHf8JVOnvo8/5zDMcYWfJJY/wEPW2wf+utAxdprcj6eBWicLh/X2kbroQ/Afy
vgso5YEG7whqbMit+Ua9fo4Hl7S95CcM5JJSpMa6rOYcEMxtcJPZFYIuT++FWAQK
afuINziaRpDuI6BN3ialgj85JovkKx56kXTbxTdWDhB2XgmjwTiashjJV6ATyMbh
2qBgF/4PQkEw2+forimBeahTf/DFp4ysv0y0lmbfsw9Tp6uBX0W2nyNYBzvbLm2I
oduBBDh7bWr00IbQWJK61EARtmJg7ukK/5WBa8vUGioRSM74dwhGD2kmVOjl+6cQ
fM+ptpti3JIYqzDM712QTn8e5afs+8Pn9kqewm5TZCF+i8d91CCVvrdQe2kAyUB1
EaMJRh3dx0CInvh7KtelE2ZcMzXENcwEmXZMVOnOSa+5eXh7lI2W/0fNSKh5Z8wr
JsF8b8mZQUaG+IxbBvpFIyTyXqcfr7pEWdC4jgf+w1oLKxOxEjXJPytV9Jzt2Pav
YOQGHf4XOqNer9HqPlcbEtbUKEP4H1Fa5NxKLusKPjl3KbNr4+REoa98PBT7bfWq
Tl7qL1e0qDKB/khC3EP8GBO5SS0o9mh9rDE1rk7HUxQTYA0RiC5MW45c3vRycGzr
4j0E9IOnio9Yag5odfeUSuaZd3ooPvCzc/1gQiA8lmn/tX8RzGzbNTOhfjcQOKXi
W04c3C1OTcRiBHpryv3ue49K8VaGSEYermdkJM5rurKPYibs+/1MlpYsUqYypPNA
9TWDTfguZxzaG3kdlPe2I+/4G38CZYZ5Rk/ZhqsoU5y/rrt3uRQZZzvXpdnagsPQ
ZxpJOCqAWzUG8FeTBqa8o6epTOfHtsGyGtXNUHFrjG1DH4riCcwvgwHmUDEIw1NJ
dP7LLUGFYkt+QpbLNqhj9am/gmGdHJCZHRazRIvykzAhu8M+I7lhJP0P8LKFcJ6X
+yhLoUGBnuo55/Ya3COkxbC8sw25fpeFn8xf5sneMF741hQ3ET8d6zDa4SdB2XfZ
T+RAM4SlRHMKxfw2zCnk3Bm9XrPmBFHeLsaAw29ipWcacn+X2jBzbqsYkmXjnJ3K
l4gvMqJdiX+zxr8n/qOUeJoHjQic8/mRVD7yf+G4YUUGuN/0Ly0Fr3xkFkiUB5L0
Qi5bP6pxzzo2XRe8u7DtfF8ZMksnYOzDR9dp0NJRCevYUowR2cryFZHloi4aAsWy
B42bNhCXpTICQUcsaUok9HYSqKHc2Aeg6LDYP//BQAHLY0+qylFcbkzuq7xlLcAN
sLEevuLsUyESg+dWOthz4zAhLXEHsmJtvmL78HlkoY27hZMmJ5UFts9/og5jQyIL
qfeKIIYhZB6ycWzcuCPL99kugndaRai8r2GvWkf/6NyKBjhVrcnrzeJMYlHfgVj8
OLf/2ExDTV+11EjAQJyIwuG1prUSHRDdDi+qccpseaQY3tv0ySzA0+Fi+WdJhUKa
LPBgHxOS6l6b4CeehybgIcI73bjzSmEf+bZGIdCZrvjn9WFNYwAQDPq8xkHo/Zoq
fuLZyApZq2wCsKMNol27zYnCau6W6X2wWqlhzH9KRakJzJfVCbJ6oa3YNGn19G4U
UjYAmbCXp0wk92ZVeOr+ExwVzOE0FuEnlumSonUX6EHYDYwd+UVjdy1kqWYFd9Tp
mamiP4UCg47UZzuxrIigJubt42YyeGNGPAM98DKNFuCvK5ud6g+XKfpUxfYdRUTh
XDQGULJBPQ2UDa0WGe31dKF5R8D+WiaN4qSwgDox4Nr9dgN2bpUi8nKB0yjEf3gI
p4mrF2LoSATdHUjdIzPBMvtQsUFbAiTdidhUpvDRoTdVdUHqGH8NZnNaba9BmCVC
EhEuGbOZTpMVXylOiSnMSnoTLMq5w1ROKb44BmRZAvK/nMICM1qj1S+nflP1ysPa
Ra3IVVrQc7NTYNAKNIOfa3ZkDD++aR2IYGFAMkkdyOM9YerABlch5kvUPvosq8l6
kyV95l5cCbbpLPsFIIGunOKo5wDOEQv+kWyEMRVNhQKIErntyXd+v9GunpH1p3vh
9MtXcnu238Qg5QdcucHir1+6mjMNQTsfyYbi8Dzd2vePDenlVvRyr1Gr5TwBqNIt
HQ6l/pDJ0tOpj7QDhxz5wdj1nbteq3auRLW9FwUePpKhk9x3j+/y4gLxqwKBMUui
ZAupjI58mW8jbNRi6lhvUnl0nBeK89MGK8jqU82FOb2VakxdzJ04VQvM/NhSLLUY
xIBFuWVnfcqrNH2ktK+W3IYUb/lIleWNGF02xvS/v6+Ll86ztfyv7r7j4ItPjnRO
kxjog/qgqx6ihfjYCxWsu8O0NYGyVCpoEBqIsiRJvMqEZmKcFfUTxLnfYFFwz50q
vJDF47yWBiAqC61mQXXMBjHwmCuQwg48dlgecHs0IPoXINgfw37QJbQDgOw6oDDA
txr8B7RQ3cmMZO/5AqTM/2GlAzxhuOXEmmB3dWOqhl/2D7a1TWgi8T2BypVLIHWm
h0DhsZGL/Ij8c7pXENqVYe/oEnGYsTa5yrpKfdpMFmc2oLf279SfmsJXnJtblhg4
YkoMIquboCP5r+bgTW5XKEbyQ6dI6tPQrBW9e/MjmpC6xTIJwv9hMtwmiP8i9IMZ
cz8uz7JbL0mE99ApAor+UW3yBRc34w/43jknuxPcXvphW+4HMWEAzp+g+wc2xub4
8CpWCzenIJH8RFkKC3ToaSoFl1vUjwXFbe9rnaQkZrN3AEdqWfSW528Lh+2Herwd
E+6hWNBBONVtT28JFMRXdqX71b3X20IJdxU8T/9cm83cKSYCWYQYo0EbA9rS+4lb
P4S3Xl4zD6ZBs8vbFIs0snqtm/V4Orv37MINw4TBFyz0oER++3S1pTx9UwCVtDNM
oe1Y+bESGG2exRmMiTQR8173cbgKIo7PTHwwEqOkDNC1zz50O75CEa8bt3ejnQBV
jZdGNDQ7WZ71zo5zPZFvSgdmVOWq1uzI30zGNY8JG5wUub9mIAoj+oEpcxEsoYbN
6vjAZL8fzjaDMKiQhqFsYTy6bMrah0mn45jYz3AiLTVZnJEtsvBo0A4ECPP7Gqjg
v7nyHc0VQVWX8UPlRop9bfApd7LvXXkcq41cYEiuqRrtY0fIMgIHmra2n1GT+w2K
mhiT+zes9W5Mpa5gANHY8+7FviCcgctACTabF6vY6YiUhzLRUuhsiek6U3nq39Rb
+PI62Q8Nbj1zGEdEuBd06twvFG3u0zI+dLcNCOt3fVYQnDmS8amqY13W7jlL2s75
SWxysE2jKxJucIAdPIN5MWjpg5a/hnm3icvYadZlPwMMYNS3IF9eSA/yzRC2os9M
vfpJn7pbwMic7DdtNmQZHBSkbNUL4siVS5FMZA1OtrlMFJC7i1u3jIsXmaqwxceO
9iYnryNF+Z5QYx9oKZARKYxj6XinNNFFyLgRgR2bCQfVnTyQ5Q2Wm7C0aCq+t2Hr
MhW/yinY/HsOw0H7fvdpKay52N1k7KQxMkxOOb2OGO2B4A4ox8nP7HKknqvxOuJD
ER4PZdofJIJAoGf/mIBXTvPNINiAHwt81IVmHQeKbmxetkAVQGUcCPVpeX0ma3cw
B609roQoB4gnYROH3DNy4xqURkZVSFFGA+cDY7dQjGiX2FkP1MXqEenkIL9WSeeI
dyHl8pGBc9NVT+I1Ah8ew02kf8VV4NtFyXnrMEuR4J0qtr/4xwiaIaUfWiJiYxl3
Sjh3lNa7rVot/gal2LDcF2zbTMeYIBUr5l1wI3V134I6Olf4+vuEXWWALTTCL1mv
JXW9WduNED6bslsMVA0ivsdja0u8smci2YKQWhzYQKWcrZuD10Gxkqlov9dkBfsA
gKtvfdAFqxjGnbYDy+tnUq7nLVxTYokHhYe42BQlWIM2J5dfWmyGloNSJ7rar3NL
M3uRR6pHip+F3VgUIxTQQcCwWm+PLBy5lizEj3/UZLdWAOVgmtDTvmnK6bU/+l06
W9wPc/vYUdyAeVCjbYq5awlFdRJGfIKqrofz8O3xkG0Pz0SvsR+MYDmise0xvLR7
dzRb47R/MGs0ZoCTdQNNdBLOuI5unuwutywQS4Vmh4LB2GBpCMeXMZknwd5ueTkZ
WoMVLobCPOi3eRPsrz4QcnO2FtINnn4gfLuTdiEbHvLHhZsCXZBX7KQpbOOQnVFT
UsCsihOEnNHQUpw85YlTVmvup2JFZi4Tz2cFuQXJtLkFkKXmRHyCKjhRprWJTFPi
GKnpP9784NNXh0hijqsBotm63tiTYAhcSveblxv4rZE3hb6wD6zWiY2Kdm51uqhD
RjcQbOtXbgzirE18OYpmwv2oUS5zJKYeUn3tVDhhRLduQlMkYCoB6PM4pEG9dxh2
ipsm67OwU1gm6QzeSbFhsjz5futmQKs4oTIVqDCji1GSyq5d6YDdvLFplZ+2+0D2
NJRnTzUGSMKk2UVegcN3Vri1uPhBUnco8ph3k3P+vKPIUNcVRrMPxSSRwENLcVpG
NjBNOdipKfVnMz6Ai14ZwaSXoxL8DIt1m0dOfz/VmeluzwZrezxYx3cAZtc8AQUs
J1dq+Tvi8CGkzFem/FhXUpF9ZnhJl5wPD1nPqIx4GSX1qlRYvIMVulonqVlHr0mG
DoCeu/1IFZLf0bBjfXbmLbwsk6QQJfjmo7rBuO9NsVSpLbSyBlKjRoI8UK4QVPLV
cxadHWg1PRqaWP7QrUoRr0nVdvAjlooKT9uityKfpeVNCJDqhVBtynKPHcPA/ycR
x1RgpGwEDriCKdW7tltuBq4OwpciZx0BNW6lAp2g0EUKp2sqwZL+5Ebh4vzG3xgT
9kerTXr3kZ7ktIZcN6xImLSAWFvOpnnPtfNhGPzUftmbmpkcB1hRiJf+POK6pxTh
gfGs/O9AN4t+BobgiuZAPTgbaSH6rsRI4UKDWAw4H1IYtrffBk4MGPqxAR/N/kZq
O4M38PnqX/pnyiA3/L3e+lHN+yT2Ho/y1pVZW9gKj7MWa37idU228FjdohCzFJBd
5EvtJPQmpcrHLs4GQHPKXKfMyyxG7MUyo42+hhVaQzHxsR/iIQ1+yII+MZfnF8FB
tmoXsbhVDAautNmR0buQV4CvLoAsmZZBTnvAEQyy9/lckjSmXMZVBj7Zl7aU/6dY
3PsmK3q+TIWqp6iJRXgHoFVgAPPhQdUrRQGjYFW2kZUI0ixUQ4w4PlVEj0dd0hwd
7gEZdj2hHJvRfcOVkXUWrPwVAJSUUE2YipWQe+gFhHQrxDM4Mnr5FulmuSuCU7q6
jw+J3tBtkyRs+akxmWuAQ38QCEFMrBoPsmASc6q7ORGnMZcYICiza0JbG4BnobYk
CXFOgmI6MnxRPW56u9JZK/9erjmYvS/gxjXVPZ/OcOUQxBZisKK7XOXs15zVIMIK
Ceszgf/uTm8SWqVWp7kU+FRldL+U62yRW8+SRVRwM8k/sjm+BesmmcEwWHvcmtW7
C5S2ITHylHRXCDq5jPneJykB0C7eynf6I57lqOZg7SfqibIiztEkf2Fz4LDIVAN4
vx2CkronirdsVWmFvZRgV7vgL1Nn+I5iaAOU2vVob/FUeE8Ghxcf2CKk3cg474oG
vS8MSqOz2+ms9eBOLnjEi0zmIcCeQ3hJqGi80jVB2CifU4DhvAGmP5tmzNt/QVOd
wOjaMoiTP5f2xKNKEiP5Bi00KwxNltvagDj9NO9b1bbIcn0wgwsADI4YU3fe10z4
MYuj+L8zQNDuqRLtm2+Mno9ZOHCavUOh8f7k5tvmUZQmmJ2+W2bbKcHEEcoq4k4v
e7uxG1B07pj3+e+599nYFbkslggp9+3EA7c2AjsqunvyT2NmI7feI0gWyNgH93CL
iDhmcKf3SsV2l9523lt1hGw+dNMEU0kpGCHvhdAW55cr7Vfcd1/Z0IoepGqFEARm
7bGY0fHNTMpMY43rXW/HECj4+V6sEx4QM/RcyT+BUIkeYM2sdasClNPDy5pkPIDx
mRhhhHv9QEi9kqeqoKjxdS7xdJzuB/5gbPu/f9lX8J1gffncG7LmYT5923tn2GHl
WagqO7Hra1/+vgOt113jRXVm1GNQ9MlUpj67+TR67wodPrH/wy7e67QBAGDxSacV
v4wvESnvzZcij92p2dAF+WFb2sQ+QdK0HQ0/fptBlEF6YblnndN5oBjBjLtngP0d
BXu7aeQk9KcdTAMZetGOeiAXBY+Q839tRh7A9MzdGQZcvXB0uvAlSj6hUfPX6xt4
n2Fm8rQW2Ztv6TR38y4zoHiYQlCls1tqercIP43iz5GJmr1/xMifsbKMc5BCN8L5
JNwx5KJtFkaHXOozvO6ouvO2kYRjkhVFPex5GwfcGX1WHZyDX+RIeJkd774tI1Cu
n0JuYjBjbFgLYvU9S/PpPpBwyH3Aj7N76bNEkFFVKomt1Vt8iZ/BxwR+hF9sFer4
V+u2C3+UcQjAgrD80ScLeDMsHynENpXeZe/dS/zPeJjv2uPO2aTDC6yK7Rf9VIL9
zBoyyDYYyVyKYhgFu6pbLLRIKbM+N9t1g1yTfsW4wSgEmSb/B7bZuUI5x790Ev3a
yGY4hklFITNgoddg0eBFJK3AKpWJATK6KSwyUgqDSrBAEKbbkij/yrYO5k0Hfhg2
Bl8w15chgFVrM1Ko1qNCrTRAGOXQsl6+5ezBAIRsgoIUN2cpyVfLXoZi2S0I/mWa
31npIWPsWq+mGNRmJpZYGjhw/AF4ZzCctLiDHDZ3yzp3PKvt/hLbZVlI46bX7K5n
yBTxx0vaBFifTdedj43HPBIWjI0I8xyQ9yEOoeglYBaklU65YwIMlt3PlhBN68gy
bk6IEqOVG2yL17Qp8p/BC5gYiq+pkzD8yZPi3AptsMZ9rAWcCzu2W+Aa+Yo3d/r4
UoXaaBF+D5Jn646qBIbHqw2+s/equ/H6FJV1Ngg/FAhHFNfRAtGu0SA8LYn+19Io
ofhrJpuA5HZwd07bchjNCAjQLwTOqtYem8R28ChrqMjCxpBkKcvBpMELIfFCa1MH
PUghIgL4AdZNApdDx36gGfHn41rEZiWKaT2J5UX5mXNb/G1zi6RyEwNAxySc2Mee
nM3tgSpQu0FMTMozjy9ay6Y41lPT5uQou2YTWTrFpdBcdg5XVFsLh6ZOaHGBpAha
Ctshdk+qKMmrUjQO5AMAkB+MNp8/ZE54rKOAolvA8fnF+ssqe3cvIoPBmsNITqpJ
fCllPrv7tgxL13zBRds6z96uc3FgcvUni0ooQ3fGsk9KtXkeJHIVfB6n9qNIQ512
sCbrUVmHNxg2rqBO3pPdplaxNEWGacwaLVtr9Ej7RP5ttQ8TvkdtMl3kE7fGREi7
dMRt6/CphJAG4ya58DeUIpCZClj6SNFBNqkjc3Ygkdu2xqyLcFvCWTY2D7PK/pF4
gfjAJT23IGCJYrckV7oLn295n1avuOvu/2NB77p1D715LnRs395BestyuaGIeTz3
HQjo7GsiHi2qzZqeZcHmcdDp+IAqjtKP+xZX/Q31zEcifCdu1rotm/Jy1rBuC1Et
CZ+d73JtorIs5vIRSkvj6wr97bPkjQ9qNZ+1poYXxMMjt4lae22QPFR8HfVMOzuN
7RzEv0pr/1n13A4IULWqwrkAhKW+fmQtCrbNbhLo+A1zb/U+lmLxJPzFWlD3er3e
+eWksJ5Urle8lV40s4qKsJSV6eZ4pKqhcOnjoFop+J1ZUDdcMXblSySQ0hSc23a8
zPu1+WNIe/Syu3S4QdgDgrBSQJAcdwJXUvxWRyjS2FMleio8rin5Js0z5W2hJ28B
rJPn8wEjLcZll15Qol48aQt7qO+6o9mm8SioxB82j2cSq9kslq4u12Intw15M2p/
G+87uyqfWEFNmF+QMNyi5FwDX5jfQycxRWmBW7S+lh/J0s61nK7OHuhnrpMfPi/S
0dirHRqAUVqEtyn+zl8+KFHGPmMRBSYxYLTtvMEyu9s6b1zBPZ8HU1jq/3neEfdf
k7+Wt0IcOkJerKTQ3hTQag0+jEme/fgLOvaEKgHn+ouMd2dqvE7wu6ZHLcnZISnC
Mizb79qa7Fvau0pBi/9l8qM9IQLN563vArxdZ2h4oVWTmUsk5Wywm9KHhfnB9ChI
qHEM1fn73VWrY26AyPbj/nrhdWLAW8zqHt2cEsxkNn+ej7IGRfRloGjpfugK+iBM
4CrdCKkPlQ/fVi+KJ2DeFrf3VH2/evbRjWc5LYUVmR4vl1NS9dzuPTZa2GeiMyGO
p+3HO6eYJjwNr62qtJ3RXxrii9BF8/Zc9ajp1kO+UtFAzXy4sYuycAcdJZbdN3q3
I0e0/UAoWVlgmb46coJmTF1pxpUOpJUzu3j0C67z44efTWbX+xb4J3aiGrIazYFZ
XRVdSphIhk2a+vLfv5ABQgA/Saw0QY7l3fs0lznjGDvHfql0NG8v4PkGG67AHA3O
DnQi3N4nGO+ELq0E2In77SCYmn9A86eCfhadlsRAL60tI28mlMJM0moQljVi3dgE
QA5YL2KuGLz6KNBWsy4xsoNMEpqgWFIvUPxoSAKv3Lx7XkxxwblrTu2uN8Zm02Xn
2xCh29RnldQZQ9YnYQdCzeZukwOAu+NInpZftM3erxkfO7KB5YhdQMoWGw3BiiIq
vALX/Z2DpT1089623B+jxCdhWdYtbZWypmnl6WK8dVn2AbVeMnMfbEmOmhOxAQb+
XZDR/TOvk2ZnQ+tNjfDGEnUQoyg+TrMQvWMh55bmAOo4ninlTntJwDnVayS2RHWE
TIxCVZXa2SKKW6UI9g9MFYfdW1EPgap5ipdGA9x/3GwaT/KFKlO0g707NyBJSZP8
VyqawvEf6lVc6LFzwaTQTN1VgMto8aL+7P9hZIr9F+UvryXDJRUnolNMU6sqkKE0
I7NFK/J2/PytOYZCRRd93qzMRs8yJztbX/r34VjW33myjzB5+usxTO6yUA5f50qd
i7bZpnDpMEFNaq9xHwbGTON3/8e3zafo/q8ypwesPeaEarCYgO6szP4pbzsuVijB
0uUgf/r52Flm8RFhgHxMc7QumIn8J8IWMt3HDNZZSJvduYrTtb/9BLU5aQXt7noE
u7iPAfITKEQQBLP0BsRB6+CavqH7htZnDoAKtx8nhTkNLYupmL0/er3WGl0sW9XD
gvt/HY4qMIxyNkM4Myw3nG+tLGmzjx4rfWrrS+2g0ibuxL/jLL0uN1QYgBGKeIy4
qznbXyduJINW0speshrmjrAFu3L6nFJXnIXEk3Hv/zzzL64sSjie/tLPalntMVbK
ujew9ecRmZPIAyjv93AD0IVpssNqrasSj0J3R19ciDDFfImSv2cwhOb+ozTosOSc
r1HXvxSM3T1NoXK8JDQ6MnS/yH4y5L7hRdq0Lq572SGkQB9EuLd+WCut59PJZuDo
kdDXdK4cV2a0Oh3rODkOeBSJ0n/TGNVc22RWfNKLkA3zVLZzUhJ6wWmIG1qtrrvW
j5HuuucLzz6Z/f+tytRH3uAm2ZSEEjMFxLnkz4XIF0yHvG/5EdLD/I8l+bNcl3Em
7lQXhQF302kN3iQqsl89xYknUTSNx9oIxyKAbU/a/Ib+ZPbkcBrmY1Li16uLsh/n
+o9dCFINpAsi7n+nn5KmuJp98XJrlLMFX5et/VeEorLT293fkroz7kIRC4QYMHub
qA1mqpHVV61z+l7vEk5DLO5/p3mQX7fGD/DhPsm25cdLrhWtL3dbxeEZgFpuRAtj
M71jmsyjOPrip7m0cI7er5sMWmm42W2uSt65+SYt82CWW+kSRNKkXCBmMbcBr+Kq
rBugU89pZRMSCl6H/V7ljfZZ0etuaMV9BZUeMHVlttRe2XCg1HPx+CeXA9MOHAF1
f6ngFw9X+vvLlzgPYpIOwdNzdaqWxnrmc5WkrUA1cTmlTuk3kccAnjXcHon6ZUat
mXFVvfG0DZoPtEsESmXkfzsK84FnfKr/ifHGv3d4c3ciPHTo0GgkiOHjqNsDZG4Y
I+du+ivMYhovPa9qTYuJ3EpOZIDn4ymzIHQQVr20mxbyQlrsunWNllitcZ/7XBMt
uWtiBrDWymoX4VG5UCqdOwOBvMRiQaFv93NEGFK7fLM6SmmI6egESJOgSwjRVQkq
cCxM6NfP+YPd9GXZNxRWm84UWL1rQwL3AVtcUIa3EdD2QRcRQwITx/3qQTVuiZb+
ooNUCU4CPbE/4SzwuAZHZwDmR92CbjTsmcmha1CFlyWd9pbiG671J9C1AFomZx4L
n9QB11MtGyk9AgGc5hhV1c+Ib2jaTWJu5wtvQzEuUICxHMx65mrZMwqOdhwHUIH9
/7zoSywaAtFPCfRhgTf1lrXt/Dj1zPzkhFRGsGpFD46PiEZU5d1ogvPvJ502IIml
8h+XEOzChhaqeJpVE/hqMJ62L2EMklt8GDbY2aGgjL1h8HjPxjXB26W8wNmctwuD
fGw3i/OCIvd/vYPS+0hSO7CzunE9JmUgBOpe/0qyYWC+P5KfJS0aVI3M0665ftG4
DTVv19x/totjPoTq8/aSTfbEfZBs2HOy5x8BHXKmESNT9XofWaNEaZ2Q8makxKwm
vAJ8Yyf4U54Pw4s6uG3lQlYgtwvfFwIPlXtL3mrSdONyqzp5Q9A4uk46z4TzdYf+
wGDuitu3iszIyPU3/LNwxnLjGZ32FyLPVfGa62PY2H+jkdYSwsDjMeZbH3z52qfL
ZmcrCyboiJB0Hha/D78fbzoW8DjSuSuol0+VeIoKDvKaceXDQvIkqVS+97UWbzdF
RYagc+IYjB0PTLfsmq6XBkQ0iMjTtYJCQCPEtHrcVHuKeABTpAosBkojm43ay0U8
gRGVTFdgYcFLF/ridpgSj85vjl5T3eDgVaZ0F0prxGQ9+UaRU0YEkhTnUQ6XGRuk
GQAO1XMLgsBRpSAfRRt/e1yBP6w9Za/iMHNyIwgKeT1CA5M79KQBA5Q08jCI4KqC
CifC5ffzZJZ1Q98VwC0Kfide01pkzTIys5i7rNFhiRuyIP6kaEm6YtyUTi3QgrmH
M8ZCt+sUckIObBUcyNrVJme88lX7pLJT3Ffs14ODefV8krlqjtPtfHCo3I+y559v
57jPZJyz8JoEVEQlbFnYozifi8dgykOjHFOJhx+Is/j2ovJyT2ZtNcHxwtwlld7r
YEZyl6uRWkN2ZbkLOujDt66MKktOWBNIuWqAfAty3GwSMQyiy2aUcf3nFE3crJCD
GD7Kg8FHUMWkX4gcQKVB50ZVAfTOV7jpCfKuZL30jH1UhlV9RvWWsu88aWvkI1zK
ptY8hj5isx8/A37mc5GHY8txAShg/+xBp0KG5XWUve40ZG9Ly2KGTvl4ZFbdthkL
cZL3TRjv/PgvDAPUixzMnfO+y5FzeZI55Qpw9wy/K0nN0GeKPVFa/vIjGck7F2NH
214I3K9rGks05V1sp4ijx48xO2gIMDXRIHCBC3WhLbU/Uw8J2dNU5NPbIPR3EXXP
k9I3gCNmfetrM7tGRpVzEjvk/ZK//gQrkblVTxj9ex2nY8gu5GUBrAyQIdn7WIKR
ed+l+1VSxIvw/BvCcoggmEyiOTmGvDmkF4HdmSramzbxpIQDUN7cnTt3jzm6rlav
w6AKYqSiIwgVm1mohHtnOd+zQFOhgQHVebig5I+056BBhIguF3f4J8X0QO9bHBTw
DDV/H4BpDlkXuBlb9Dp30SsntvKDvgiBT2sJEUIT8C0MfWFFLr1K3cu2H7LzlHdd
Ajd79lqTtWmM62P7iK4u541pCFeciWc1tMc2hj5IZ7Lg5l5OGjInfXOyNs7QsO7X
nnS/DOPsEUac4KURt/O5wb3qA6kwd7O4Vuq4ESR20WB/ilmidw8LwhVJO83wtoHe
evaO8noINdIvEO/20HKOYzbR9CgUtcR2aQfyM+I+iSbP4AT08OYgKbkOvQ47nMRh
+rtz0HN9LBXKwTecustTOQ5IBg1ADHZ2brH78AJJ1dpRseJhDeF01CrTFT6qTtvQ
qNXd4vV93imvDpWp3JHJcAHjVJkLkHSX/3AEzGmqHkzCc7xSf0Zx9QdEnWp8WEp5
MEer2qfXTyKUqx+ci1MF6UNXZ2VsrVFFuWe4U1aVfs/5xtVC8OukvJzlkyZWtWMb
ajIM6M5dWuipYdrCOhTwFmNXBEDVPr4Mql5v5mI5nq1aFNPCQ25SSslxOqK8dKwB
4tEOv6YVJ0EntoDEdbEyIX42vP9j7CKl85r2IEfo1Xlq9XhrHcUZ0cLg+FjCnZE6
Y1qfhMKXIt1JmIEkt6LALjCgHHkTnBJm/cpRiRfPFApNxJvuzzRYsBK8AkDY1/CF
Iu6PysAvVgw4NNPRzx6sW55Fb+Cawx6iytRp7byBzRXUoXi6pT5AnYON286XiKls
fBJkZF93q0A96KHJweh+ZVtjO86iz/vksEQte+sJmOux++wu841o1pc1rFcivxjX
g2lQgePbpvWR6USaDrTQ2LS3gNQuht2Kn9SEDR0ugR4LvGVVFvj6hG3T0vpjyz2w
aNoAQs3548+eI36J8WiZ+1Yjp+3ZxhmlvTPI9Eg8Tosi/Kzgo2RC4a+KuosFIhZ0
KJL+4+VG6CRBz6ms5p2vMupxSZ0EUA/2dDFr4PdHtXVzxWoQw4ae3fQRgoSlobNJ
MqQGwOIXr4Xloq7Wi6W1IIah6Hkr0tCTNu7SjsOQegcoZafPMasdNK31Sas70V7/
TZQ1NR/wgPfGIfccwDfciJcRkVRamI6smUltDgB8tUH6QNWF1y0RiVVAX4e6OlvB
LMSuixstY3igSGhv9bQG00JQbVwlp62rvMyh2a1b25h4/R7Ok5J2OUMXITq9Z7Ul
UhgxxV0IGbku7sLA4G0UfjOIYQdFh/X76AVX/ny/UOY6HEwuKkrmzX0fyMapmc5t
PwpK3G4iyOw3CD5R4aTKoIpJhug/4PjNYXwouqljkoywXP+Lp4zu4tjwUeAvXvPr
onL21nATGfTeijVPduLBIgQhjqTccXySPaHnrNMvmMpmXPcmmVGZg07IyQx411JT
fGctiN19ME9KtnEimfPHYRDMfiZ0Ix67pAg/1nq3EE9YHYfclcATugSEVsAh1Dxq
C0jaJkQ0/aClr40rvL6eqzUO/yTNGN3a9IuH29nEet9CIONp2cjcPJXMH7H2cTsZ
dbtNMn1e1O4xHtLYtK4MfYQP7x4or4HjVdptRkWaWIYpu0CwNEIq45GhgRQKjSNe
kL//oCQpAp7thNd4NBt7IOnusT0otMPixwXcLaGAGWuMUcQ2yPdjOD82Jzb6ueaJ
Mu1Glgj66PTGfgZBPnGWlIR8MB7hKdGYgHAJ7//ig5Up73CN0Fvfzzza8jGYHDaN
EBPhZAmcqf2b257Qupxl85k8QOK0o7Ja31zsycuzN5weRnWgBM1qGwLPt/QRjlsI
hpN9DfEFb5ShguFl89LPD0NyE3HyCwsTRo/tcz6HPCiYL4YC+VYOsBPW4HMsm72n
lEpol+UmxoJwBjBThOJVGDaKIe3PzrHXqe4IkNCDrbC6Cqi8jf+LLAu5+UkA+lFh
Y5gF5QUtxXvwwoONqWP6zH2QwPQ76YS++enGTilrQpdZ3JNi+8/9zED7Npisso+e
o1O0+m0B0cW8KLM5JOPbFFjoKRi/UQkI2P7h2P1/JvvmZ1AJDPwRGh5p7++pSHNv
Wp5DhQpHP3IFy0DCmV7w/WPqN06i2O/zy/Cf75f8RKMsksB4qDznapojxvok0pTF
ENvTUChUf0OaV77chcnwCUb52h1sC5Fq+OWwLj72PGmZk5OkyPTIai4jw9stXA3u
WWhg0d4xqQf1kxaWBWe7ba6wlHb2fUrWcEba/wUrFRyZdxMclyZoXi2WdOZ3Qzt+
qaIi4Z9usT+6jelf4rQCL02NvrbNnwljMTTVOlI/CFXfeEnjKvh1gCoPWzkWoWuv
weO4lcIxmY8RFsRWOJZgh2mLxfH5aDoVtVuThvZDAKqPkUhwLR6Ao+LI6qfRu+PR
jK14LYQnbAd7YPNLFzFQ7dpw6zPNAT9dWaX46DyEEXD9I3uGV2Wxywj1HrogB0Nn
dNEFwqjVn7vFWYE+JOTpQX1pg8UGSKJmkb8F+7ywS+3ZdCTBhUb0XrV+kCIVlOcl
p5uUb1LRjmkpWPrwzy4+FUcK8y9hM/XiWj0a7Kiz9bO4sDNmJ9LMAN9mE8RHfGo2
AO6bR6h4xMojKFQEKBGVis7qxNIjBIGNSmHhYSrv1ki5GLg5j5euHSRqJvrpGQx8
F+riehdoyeds34E7lMYUb1E7MyHPgHCgAYW+D0FSgAF7B7UDpPRxd+NRiMd93Xp1
AedyKYLx8MSJrBDs0P0M7xRk6w+SC/k+Y4Arq24rmn0QRbTMr/PbnOgqGYm2WpXC
JdIXdUMs6rvtx+3N/i8U5mDVmjGrWQcdkMgwY2aEZlYvgKLEeAWz672G22iaCSBv
s9dUx/Yz0JxjCPgpRCKTsbK2qS6IInRjsNidFnmqSQIadJ8HigfwU6xhy3XCVvP4
M2mLEP62LhtQIQ7cjqZ+HeoxebP9x3/vuSpE6d6etLRu4HPJdX5+4wYMHDCBd8Rt
vQMGIUhxQrb8RGk2L7SedZWzE9+KCG2RyVYxZt7oBBxgx4VKOBBYMrd/kOxcEwLC
o2RSi4AsncZDR6Cf/cM8jzo3CJLNPnvDiMGI4k4dZwnZGzB2vqE4uZAljpfUaJLX
lHOIb4bf8o9Xl94Kg1I5Uh8e55e/npHmdwfDLvBhcPDVZxCeBmDDb0kmuQWhmzrH
YpcL5T5qHR6w8uQD0SORRwF63hDuZkGwnKlYQcdd0YI7pj8cy8tHLNSHqVklJm6w
m//di0a8ToOrr1GU5c+4XUU0llyEaNvywmB1HZRZI1UjBliZZA1xD+07YtjTAboU
lfggLka6+8sSCd7HRIb7ABTvIN58SeGOJvJN0DOoimbLzBaLvtpzau4ZivOrX6EA
3lPU0isHmvu3eqDmNaMVbKNL3ruyeOiXhmNoUwRM5Oyf/fXrBQROSnb7ciGa2Myp
o5cvZVBHblqApjIS5LOTe2dVKtB/3nGTKW85LQCeuZXjyaQERIDcfzu5Oj0pJMVp
1D6G8QHrII7swXCMvbW/x6BO95+YZnVVgIN3Tm/zG91CAc9uwhZmoxT69hIkAIii
HYz+iiVuULjEjUdgHC/AW2kwB8tI4ThHJQnspbLAw2cII6tbd7Ddb37xOt1QQxI/
qMqHYashl4YszeSTxfPBIEuA7vqNZoK/4nOdgMLzEHEMU/WjiClBVYr3lXXSSuD+
i7oT9Ii9up78Zk+DPdXshgIFCDRcC3ifiQ8NcBCs+VeZDGxUEDyILED92OH6Rccn
oltL1KnLalwN6zIBshQxLTkBEf5ZXce3AMCGJ5geDwrkrQFdFeZDGJiTdelUSpri
jp3SB8CPsXw6IuoxN/fk9aMKqCH5XQ3aAuO49wLsaHtg7AJBwlczS3Y3ksYO78E+
qu4j6TpetZVLrak6ryjXg1AYRz3HNpq7VeFpzD+hTcXWrMmr0mkkIqUvkKNbBiZ7
Vst4QSgy8YGr436IcB59+TxhYCdIJZAkAB361zm4K4Ifya3e7cqgfe5TNF+lehw+
mBixFAzu3DqdOph2e5NEddLPmWqEzDJH51exevMZ293V5Ww0vSSUCVmXgN6f8B+d
SCGXGXpsO2Tk9896CbS0vXUICtUSq4TwSF3wgla5Xlo0pxJbKg5H+6rrguRMsc46
c7BoG086ZdmRnp2Q0PbTPJs9xbTzwhmol4NjYMaGCFHs7PojiEm0KD06eV87ZAJQ
pOm2T+8nYjQcVA7yJ4uDe5ajBYmg8/Pd/4AZ1p+kHQQ0PqM5KGGL7VoPZGuinJ1h
5tqBrfDgmz0ruGPXBtEDM2S9BM0+J1OkLqGIjo7bPCLpQxB0k1A3f2FLFms1rgzb
Hn5wzLSLaQrH6ecZKSxYXOU79Mv3nV3EnDv6ArWqIundWO3XV7onqPSeYdWqJBxb
G85806jXUpRcPmqZS4hB5yhqTGbAkO6SSi508n9YBHpGP2TJFAqdzCYbVWbx8wXs
uV2kpSpc0R1n0hSTaqNo4FuABqxM6kj/cHNrhbc/yZkonAKa2KGw/51qQ31mJGCw
lNiDSCWDGhXHUhK3xSZVqMp+cKTzcqcubabuE9L92dwJ6zLWEYZC1mfLz09gTygq
ETkb3eyzoeWk2bDIxjE9qTY8W/kTRwHEiNBLKvLHsIFb/jzFXTDgUGCnBGrj5r0i
Tbx5Oxn6D4DqXiX9fNlavSswql6+zOm9CCTvsoCaIuTha2N9kE/wL2piEXgr4Li6
E+IMGD8nR+6Spe5em+/DO+bumkD5j2boexYpK95Hf183RnxZJioHF0JwpZbFQmAR
rbenhu7XfL2LyANUt0DM51P/5uSO7wo82cy2psMjGsdlt3MtQnELOR08JDGkJxSl
VeUhpDIvripoP5+FVgdfWxPEwtL+PCzh/ndXYDkYn1IHGB+gwVqIf6Swx/XnKHOt
rX3tnyUtpPrdd0aQGX8LL6OuOOt9kZu2BusqIeHFMM79xIGWzljC6uEjzMPtq3vo
8w1qV48QjrcSYHCV7mWrWBe2g6Qdd63/yHXcdGCLa6pqmDborLknINTbJPbaAarN
QWYQJtRfGipmCEKXI0g9A4B+OxcApmmg3kmBx2Ut+uAS0saCqROjT98isFkjEpxh
hj2VaMND/wBgHxqRBMqAuTLRO9uHd4t+7FcFA+JD1CHCsjWFPJCS7RI2NSGuFGrU
VmbfzmyXHYSTeVHmOOMxZDOXh4GNA/owpP77ZiIMSrTaLM8u9uPuXk6iFHJjZlFE
QLTEd5WHRSa3n9H4BZeHIxQtL86RPgoFbv95Md9OyB+NynSA4BmPf/TvOg/ewssx
oeASCGLdZOqDdh/aSpnsQzgsdJsXSm83YGGETVY6Bo+Jm7Tuo+Wv0AIkr7DzgpAG
JRquoTXAq6rrT/vDcSIp/AHipkd3eanMVymWwUzhWWRxHHkw7ZQSIkneC/zrtZIh
W3nog9gXGPWy3F29cwwn6dBHo7tBPRoyHDtL2mDOrWQw5S9IT9HzlSp9pY9UB3qX
hxKODGoncf/J6Fhvri+hvAYlNeEAwPyAywI0B+TtCnIqokKJVHK1PEFJFYFH+A6Z
EZ7vzz4M2UCiWSy7UvFQ7ysdPqzrJeFJqzwaNEj5wgUiIQgeIDzPxslUnPqzN3kj
dABoYAX8BtHdaVhpu09g2v1i3QtUx+ADer3+nMxKaMoU5vHaifCBdWqY/BP0S9FU
j45ItgaOF+7K9+67t8Nb+UYCWQEAWdu5bsf/a8Grx+XDo01dj8lzg4wgCdLOs3VD
N6ugQa0EOPrwUDy4Q1WBWkLevvsy+2zfsEs4/3G8/93p/MAFMVQcv9s5wzjgYlvu
Fe7SAaFoMmem7pt3vetn/MR5m6gsJX47OsHNAOD8KUj3otW2IPFGrOVaHee8AHAh
3Vp97NRil7+8NWpyanNz/y2TbVuNgXk3ApeCfOEPsohb22V58JRAgm3yuzvQVaoB
0DVU3W4JxFeyMMAQETYvXSjoFVtC/XNPmj7nph+sn5ZjHcmq1W3YTW5y+82Q5ZZF
UxLKHzX4n0TLcCMLjV3z1BVRe5Vd37RXwrFEV57vePFsZAWP9nRwW95baUn5bwI6
f3gGql0EjtDhfjBWaCO4DgzMTYNBmkflrjonhW2Pa1L8i21Hy019HV3t0J2l3Y1E
vykCLQahASkBkbJvqsMgTmbNgaCzQnthVo0DvfAkyRl6t7uK8CrJe6w0YtBc2mcM
SaVzE3Gxs9bFGni0nz6JKF80KPLBLJ0/2yvWKVOUI6ofjqAvik6EdXkl81O33G4H
QwKMGH+e8G9ZJIuPTTLjtkZQjJVf765/+xlpv1t7SB2l+PlW8iaAmAXpmGroPPAq
Wh6hBmR9UZO7QCSbltFz36Q35LmYG18Yo8b5l6yTYERqx++kaNsCHn4kuF/u5uw9
0cmCCQkAUtimqRD2YRfBDvx1pEKwOZHTd4hvYgYJsujv2blyIG8kTtPsJjjRskjr
5fnS8MekQCkjy+jZr7EDcxWswqZcANCBT7S97c2vDqHWPqPVoxlXIcfdBArPMRoi
pkedTLXjhUoWGEUrYLXEZTlhE9tHOvU7jOxf4kf18ig1PrVFjaUTAgbLMkDxppBe
1vGiZXCTIEIRo/yNfOoIfgwNa9GshU9RoEozNGBR+eiBrCAhe52ElgJmtir46HCe
QP1x5IzvzCrFmfbYwTHqtEQDICz6VdPDaAhHJKud1/vjAZ2jR3FWtjgc0UaL2Jhg
q19XdIaHXNg40HvuaNZIrOjmSlIoM4E4QGebn3cJ1dyXNUEIutXmvzzGEbAWrm1T
v+L3LlCijKXvkreDh/WuLev5Jlr1PtVSeeht5cBffvwa7s2ygQ4rmtdmhaakEm4T
UpWw3z1e7wSUjjRjvUhxrJbmYsP39TKFPFj1degCM6xIKrMO0MlYx3dQYzh7UVlY
pz4yrIQjPWCV2o4crMl6w1TG7O/aA0mFHohGy+LgpqIuICsv542WwKAemFv/2QtC
x+ZVsOjcVpaO67CfqGJLV9NLOoGBxQQy7+Vy1k0/KpEj1cB9LICTKuMZwfZo9sD5
IjHFzxdBeZNZ7dyE24R5a2xBs6nH1W4H17pbJPGkcshYzdiYOUXuE9bdyxXyTau9
MKE6shSX3fN74LjJaUUIvimysBmVDdRaNusHiwajpHBcY9rMaWo3ibo2/M3OtZT5
8UUvCbiQxMwRp8WM2LWnSxlIWB86YhdFBGKT0S+qjVEY09hgQ8+9Zf8Hi457T+M3
dEPEYHQoG1Chg72ib2xy+k7TKn0aeIAlde7oCvYjCy0nu/xYIIIRs+uQr2Rnq6QF
s7HjtCsotFrTcmYgA3lkpZSAXWBg8P7ItZG5w9bpYsnb8kt1dIxtuJsxxf8l9PGI
Wtq3Jrks8R0N0c9lYSjgSS69NwjS6S6lQmzuwOytiJpyZxkgDF7FY5x0O5tqzWQB
SU40++iyynBC5sZdCTpawRJ3BN30q+VQercHIRiqr2YdihwsQ/D+7Ex9QFG5yScw
EgqdqiLGQZ/tx80QFgQVJEihYYqe3WIe+5UesAd6uqcV8ViWEpK4ATwwTuDZDaVQ
tx/sesJXzRelUGsAKPkMFhvDAjBvKXZGHj3AObmWQauuukKVPYtxpKbCMzrY7/5v
Mxy8McKtfWWPSd9lDXwJSPEytJrmLEI3MM/ezriJGldUvtHjzP3nKR51IsyxsRTd
8yd3/AidkCxcgQ6X+SKV334d00hXaHjLPMiBjTTAJ+fM9Tdy91NBJ4UWR57I6k+y
CgqRdCkDBbC53Zr6k44Pj5tO0zmJn3+a9KY+W2nxlvg8tTKJV+GSOZh0eSWEQfZd
jtMkDANPhVGR0z9MFAaLCA3O1CMZBpdy/nPl0py38WG2dkgXKHFCI27ZguCHSjuQ
EU/1JZ73DRKllsVsu83QApqxzYcl1Xwrbu7yakTUdN0t9goRPmvnJE14wHRZSmX3
QQ147kS8rpNaIVPvHYVV0apbtXjjvw7y8TMObGQk+YHijguePdn5HpjtG3oSTpj8
JHfOoj409moXPgaRxij2FQtn+C++mAkP+hMPGKACgDS8XUR9Ow3T/JorBTh0dxBL
+NNfJJbdjas4jRaj3dCLdoQvEBinpKCvGMcyJGzrjqc+agXLXoEhVYQ7hqPmYtz+
/DMbb96P0d/60pgSh4Qeb4JbA4hCFcYSrtgRHH6JEbKb9km1WzTE7aq3wpJTav/Z
tjp6TvJNiSZhynvnXYEs8qpUFXn9Cehx12u45pLQedR4PSbnAIJZJtKtrbRZQBlF
cWfP/67vvswsG6e8381r8UiTtk82iMJiKZClh1Fy5d+d2za74Yjc75ITGJ2X+uoP
0cjuM2MhDF9Sqxc6qO5FP+5XKLf7DWM9OvovqwcFhnnHXAS8f82kQBUki/5xkbjy
qz7kVb6mi31DqLRkNLkw56grymumG8+0qoRlwmE9Td1YvIFuNwMqFx3Fy/nQMEwS
Ps0JdD6I+5vM4nOZ7auW1sg+eza33k5tCNYFe964XKsDqOi342avsGpbrKdXIW01
UwM7e0OVmdHaxwDwmYECJHhetvJXdlZ1lQO9sy36cx4TY5cP1TqC/Q0K36K2r4Q5
omDCbTnrKjsyzXrlpwFSUc0FfeIMJMrs7ZJwCNTK/e2u6t3Ekfag0aI6OXPMTdwn
iDqM90pjW9LRtdCVpL9o93bgWluUh758FdCsQxTmmY0N8fMwFBvR+uoZ83aMinsm
3xKbX+OypQlB4ZMSCgDEPajBdiDMlETlIZuCnCVCCP5Rv18SZDbM3z0JcbM60eiN
zhIHmDthhxxppberWIa73k8i8yYc3Fsn4wDBCZbtf/hEDntkeMYOM86+Hnclzd8p
wUGNcJEcFsFpopvpzFkDYarmj0m9C/anfbMuKw90vKWCTQrQv5xYRKD2cFQcqLu5
/7gPw1xz7oeWCvu6/kGyi0qsVAYG3B4DSxUzSsRnqaUJb1SS+k8wWXOTnu20usDG
NzDNKVwi2t6Jd1/I3pt3UaFHpk/TWIb6D9RR+9/MMpv/QncZc1S/lPzhLzNOnddW
ORYbk5lGfKi7TUiR35/kGa6CYO5lwpW9T+FmmN1cNe5qO1YtCThW65i5LV85D50/
yCbCMiEHqR8yoJk5rntRRoyDjDPSw+0GWeGtybl3qYQDEGnfirJbc+FpYJ63hNsu
hax849Ze+fC1JQTGZ/bDvP/Z95FZWMau8Blq5t/bJSSCZ8HPw3ejnxwXBtt6gkCy
2NHeNn5jsphns0i6yBXVBmgGZFWWtqMCZcdKmQUDFQ8bH+CwglmJdmQ+wc1HB1pn
U8R+ujFWyLj+5xV/E5fkCKAW4b+kk5X9+DZSe5ecDTOI/sj9eHWPZCfVlksW2/gX
kGHH2sZtirSr0lAAwgeHZ5tTONLs5dTlR9x9LlW5v8Eer+G0yZBa7gBECc6uOoQj
Wti4zMQCmKqJXs8gvNVoU0wq7Vy6VsO7avxRbgJbNrDEEbI+jyvkZfY48eshCDi6
MDWgQRSeVfvpLjbK4ryEZTX4gUQXK2cfCJSNKnHRxTumwVJW0TF/7meHO8bhYo8u
jO3K20tIXy9olrYWx8jb0zzlXJkYhS4C8C24GSAZ0fdIGQpRao0gwQXmEBGp073U
ecYd5gQXShorxSHybuFFh4BsTPW20wjYlzAPZfb+P9L7oCH2BfusF4KIjPcnQZQ2
hynmVvpkUmOdONbCBS9ctR5bBJlnY84Eb2o5lv75QbtkG2eJInoQXvCLEVxvbMtM
U3NSrUtbMp8mTCV41PdQnfu9DGh/n/YFUZ8jUI1p8ZV2jrIKoaAKm1OX9VQu9XGO
+HLw3s3YFYvTZpFrEED4Ad7jNVo///tUDqYNJoxTlvPuXAIelS8UuPIRy17XsdMH
/XGGMYg7Eu07MJwRdfbc0JQXbBad324prlXE9HRx+dX0d1/RFENT19uRDzv3SMz6
jJGA2b626ScydjkxfUxnBmAshX88MyV61qMraoCKUwKVhl7ZRWya8ekl7irMosSt
/LjIkoXNK+8BuSuApKQP0hQGw5aRN/RBbjKEa2Px6bdNR/LoQw/+mCe1GXpQXGYn
5UU5VNw7Gek1osB+RzwVRtL/ZP8MSeDeNXYe33M9rbF9PWbjNIWglzK3nJl2m6XF
m4vD/y5+d7rqsgb/UvECUUAAoM+g1Co8OXht6/mLlVGBKigDSEBAovSG4YGNqkxy
StC+YofvwkXqRtXXiP9NaPBDoefqWWyvrCjW1wvYTwdePDbJ1t270A0E5k1i5YRm
NdFVZHxk7HaLM6Ws8qzbdLNCSpjrhCcp44gLCe7f1DUasaY7TvhT80ALXVPKOf75
KEqaDzmDnPAnqFkCqgxuspj5iBhZra9b/bA0aW5fQalMdchZvkwgWOVhXhSVY1NV
5OEK2aZrDerFAKreyY8RlWQWvWvuG6Q/AoNv2ijaUJkHEsEqdAlwc9Ka9wGbUivb
BAjMdrCylrp77xVs2t0MoYoye1JqhZLnKBIt0lfcVpvUMfQfaOHY+Khhq1xA6wI5
Ao+Cbw3EiXrSTvyB95Hl0NbhQ/NFHT44EqK0FjP39pxfiFuNz/2AQpEF7GQlcAtm
OcGPAPu/E344uJ8KmzdmavmHeE7YKmxysbFMhDQcvvHea5hCiZy5z6P64AiCEVJW
6D9VRN2dnK+sEPNQuaZ7C+nRsYDuDOD0kkfHjgJXvEFV0uFwj+7eFghaN7pQmSNC
84ReNqRCfGOiYLP+hhOgE6+tni7RQWeUFYCwCfFLosC6Ag/sROJtvohNZdAhn04Q
R5+J2mx6Hy+pmqeBVXw9SLADDKNNPGAUTILb7FZR5FiT7S5f9QbW82RF4cGEWHzl
frGSgkVMaPbv5el546JZFlTmxdg9kcH0BdV4ODRtTKg7BwDVm+nNOetwUME9GlN6
xqF1gq5fJkNcv+FHlmRhKkVpIEOw+Klf0rRkQ82zV0moE02kUyxbCNZ75s8IUYqh
Wqv7XSekIEhAC3o+LYvTcXAUwa1cyL+gIcdLHA7PGjbk4lF42T3oN+xvfo4biiaP
MD0MI0KlleaXGsZPKjKww4whwffYgqXSu/V0PuqAgD8H60hqiiqEM884pGSYOMT2
iTYlEl/eZdpJlwtGkgZS25ke4QFXZwcWBFmKjL0LRb/2tAXuxmn8Q7dhGb30P2xf
zTh6AkA4IIQUn1ncIPTJJYm0zTqNopRJso9e+hA26YGm6QkyEib7CqVaCTj8kkuA
gZitSwEGare7BM+i7DiPDT+x0klQaQsNMWzqGLEn4geabmYhwYmeP3ndmIN49phO
lvLm/Pw+vjqabNGmUi5GmWHPrqUYhgkhWanmlpomxd0uDQi87ewB0EdK/oq+4zAo
2QYJ1HSUc25jneec8J5f5VmFnU0rFGuB04VdDuOb9uV5h9MlMO+wseCL7Y2EstYO
XZyH7CBUzujqgSIva6VEm0MAodAMSEQZhvZED4Eeo0xubOiFkYROB6rW3VtZplRM
NF6ukQQmJC1+SsB+cWns22q5JLKTtgXeqjDYi7VRTHeq4AKJvukM2frgoQ9wWa4J
22R0KOzhJ/eNqluDmOj1pMOmCPJLvOIZgYTP9ZVfPr4AwZWL36UTEFR/De+cma9j
yHEvGk2KegDgOxmoj6HuMy0+u/9sIym/Cil574yngqriQsy3pMQjhHRMvNaIY6zI
wgwTKp8vHRkdU9uaPOweeF02gSCxlzCFeevBpkNC+NwAan5t0BepLmIUCJljyFSv
+cc3YiVcWSLSreXmZ6W1Dp8w/Bd57PDlWwehvXwbG0LjBynsY07hAm/xFNwAFzh+
tYUBKwn1gfCW9CCZYz2oxpW2+UzOqTYOn8waJnElyESnWxHbK8Y/M/OCjKRyy7XF
p77Pcq/lXbzZT50rNVUxnccZbJz2EHDJsX6ng6Ay+GTQoLbsdRXcWDfCBUOvs6KZ
pvVCB6vf8HjaRsL8dRjYnPrWkX0UOsMgtfvGeAxmLRtBfv1Gz+eS/X2wsz+hFmB6
bSF6LyyEEs3o/VZLLbGvvcp1gPokqXzV7Xp45KPDDTrpH52GWU41JbDmhWr55ui0
UbVZ6zr3bxT7PJAsOV4UMsmQ2XLhLOXYsa6FsD6Vz0L2PpWg+TykxtQMB4M7yoN3
T2SYAZzyAxI3uN1QQbtN0I0kacPWxLiL+MgxqhJsvcAjNE41D9dMIjh8rvglhiMV
75s1T/+maJ0r5s25pVc5sBgEOOfShnJsIZZ1X0Yyl2klN6EqxLu4x+uolL6H/I8I
AxlKEvcxujj6jWfRpD91LL7cJ/vIpJpEEnH3BaDiT6F5ny07gKpaDv8Kh8aD8bNX
72tIAO7fkjbYA5LvjH8dLgRt3LQrsHZ4X44KUQWxYXPu+kpEbHuxEMhYx4Vr7lFz
muw+ade0WBcrkcY00yH1B7TEHNXi2lmLAyBhwaXvwE8pwfT9r4IwdzMMUlAhy0R4
f5LkvsiTHH+B4fYW903vtfGh/Jk8X3Ejn90BFa7ti0Em6UpCrTd/9NHzPTjw67H+
MWfTbfyhypCJQfPoAa1EV37dIwZQ6xzYSXpUSzePOs7H6lx0RyUYRAmm0J+DeVvO
8jSWC+Zgo66b5Fe6VIDzrPlcbpGnXS5clpcjBH4V2uEJnS0lCMHkL4m0KBQT2TVl
+sbR3VXNgvzvQ1/xsgfkB1Dk2oW9larThj3CG7JzNjeel5NKy44HoACZwz+EnMP3
hA07NoEmRFo8HbO9kEgTnUZkIJ+gI/npMO8h1eia/FcniP5arnxKTgvdVyOzkQDo
fw1hpJJAld3s4Guct97oMtxnhQgL3VkDf3DKLIJDhZEmTQmg3SboneN0jkMQIc+j
U/iWg9s3q3z8WGrYL9ITErIWzIN3nu+r8FEQ3HsluEKqYRuLvFk+k5tgk/AZsXUb
lILxPzSpsLgbRClL3OjOEvIzzQsBAEMNid/eqYGp84CEXBwNidhkPvMuePzGihbh
zAwmdTbIM8s1o0PvvOY3u0pN/rdK5GyhCNUSlzZOzGzlvPr86XospwzRwWHudF36
eWaNN3tD5+j8JOwDI52ZUJoEaMGFTbV+B7gI1yzt/LANuW1vjCFlrGybGeFNiT7w
n/CrICnIzNi2Uwgl2VElFNP0d13jZOB7P/HNYHkl57tcg+bkqyRF6e9XbDhNr5K6
e3uudSWrpybaMnWyk/XkZ/3JU9dim0JtT5w44kxLbmXWdGHc0ljMDMXsFHqa++JG
CM3m4OCEyY0tM3M0sxS21lzrbAQNgUR8eG5Is7qvQc9aCdNC7JPBt8UDspxYRbN5
zDn5jRZunvqEd+/gf3Crr/1v2UmT8PWB6ATu4S5UcFksEnMZ4rtrZ1HGjgFmrr61
YPygce21Rm0GzIhaosjcltGSbaNPdLBwY+LjFrVFwfB4chzm7J9gwBtvGjKJhw7p
P9w5co51iJZ+qPAXHj+UMURe0Q3he6l7hTaq+S8Nxc+Ks4YJvKtLnGfuPLLjaQU6
RIQX9msMXXrxF52fOo3NhL7njzOLKehiWM58dlwZdcWadfzc+a221SvxzrUj5I1B
oLF0FzRoATpGh0BaPqLc9LxDhn76mlQnnPucPOjTvz7HlKxCgfFq8Xi6V1hXA7ZV
0K+aKl+hEBdbVcc2Xk81cpMqQFjGzLD1unjhfh7Yk7cwSd/09TnWJmArtuUys6RJ
v/1izOAMB4VhHXrgPvGRMXjJPUvsZuwqWt91Xlm/wfBW0rvS3M6CGTJMObj2yDMF
MufwCxIBN/SlR+X9Sj1vh6OgT5EuHoovYYoRe9GR5BY8kb5nkgG/FQ57Z0PE6dTp
xZQGtK7ZoAc6CgFjSRje+SCLNN+6+RAQP3NiX7yn56eQeMrMuP+N60VGLzIkJ0QT
wiFlbEmyuoBahrw4BitQtZdN6Y/6wwFxFQiSOf3SP3TCx6fYR2Xd/LsswMs1Wp7Z
aaeo2r8bsvnmiKTA0+ZkUZstfMGl6WvZXEJLOHcrGAwOb7h24pB2XCXGJ6xRfYjD
/HG2St4r4TpfQcI3a5EcNSfMuIZVVl6Xea0ZdTTwafzsOLhFADaYjmyIJ/YV+kLW
m1sQ6qjYTzJUiiAPI5aJBryUehwOhPIym25CfpB4N0IJHSZJaqb73FRWohUhy9Td
JUrH1xsz8vlpUO18RCDAefh1qNGPR0AuLU6cllmYmDjENM2mG0cxTqWoRQDoyBuU
sBPakS28fLNXjjS3qVZGyS+S6wmGGSwrGWe8jOz5b1pMt/LrirRoTtprxWzCM6jO
rDBDXAqOeXq0Jn2s/7mwsOpyfd7Xypttf/ud6XWfujypmwnJ5mapLD6N/E7tXYkY
xpJzxvj1iNc3guU+R4ce9mhi+mvTxHxTkPGb1GzNFkEq7CD8oJTl/8pPEvtKZqU1
ZZpEl32dqVG8QLXw/oYpoKyniE8My+DjfOIVJxZmI1Y9Qcomu4/p6ECiS3Noe6x8
z8C4pyOzWoJtxkv8w8SgrI5dWGWaEbyoZdOCeRFpHal6CO7Y+g9vykrGU0yqrpGD
iwcxHK3f0QFxJtp9sgpNGiD3HPEnvcJ9U2KXO7j1NFAlJtNfZ75bo3Q6tyL2WCOL
0qCYWrfHh7IEjGPkEOnxTAzaPokq6jIkFzkEnPz2qxoeyUsmMsJDwUDcWt/Ibdl7
gAWbxYDvmrFq2IgARDxhsQdJvVOrxAPuMIxbf32wJ6uC6FzAzuoxNNGhgCJ8aezo
4KkclCbeFxidu15bzwJ93nFcaAhsHWn/xxzj39aDc4njOLxzAt2ipulgTyzk39Uc
OO5WrP5HzPw6b7OKgZ3QVeonED65dXFG3m8UFfaZMvITOLeXEY876gmpsO18YX1Z
FOdPy2rMyJAF7dMDavRC1ttkp4DT/LniHjdPGpPyp6mDv6I8JBzG/Uw/PrsVrZ6v
YVf/GqFRlGHwuRuDm/0Afqh992tMtKu+mIcc7AjPS/7h4DjhXRNfazU2X9iXYAEh
Wjf1Dhj2rrdlC+gzonruq4W02q/WBPvi8PIepBKlglzqClTYi0Vm+1V1VWqxMe6f
qfvkv8HDtgh3loRYNq5n8YmNvQ/4xceGElzAxlU1X+uxoskwWZIpk7Ty7SfqSdHD
WeXELZXIzAll2zLWbmulNVEHm8bQsDfxCtEXZFu8GcsGUE9Kl6PMHj1Grr7LQ9Mi
vUKjqq1ZpwW52JP3/4gwBqCi6t6kBaL7IFqjwhAaII1LcShAXBFVVzdRPrnr5WQX
WeOpDXSiTDR+pfuaFsx87BzF2/dNY4pWTkj+qJW5V3XdIpxYssjuFlhl98VASpWB
RS18mXbbHa/nagdZAVdq2iBhPgSmdJkxW1JBIWLFZV7NURzn3uXsAwXzO1h8gmYN
1x45CWoSM9UqxfDQdAs+aafJSztBIpdCfQgj1qPdJPXThgfQkW990JilPBEAfrBN
9v5WnSCGNfgebw25jDxysvyStCBjv7T1qiz9JoJlkVYfsE9xqpOWpPgzQRiWqrgX
GEcqNmUHP6tNy7VhqK/pNbMJpd1DPzUkPwWnkN8dikyrMe4pnjgTgA3Ie4SxEx8s
szLK/ePFmZnwbXd5zoO6RnYTBIKeHLUYh3uCVcoRe5BPLUHdBc8LHxHRS7TvOTYW
LaCahZaJs5miLBF7TmzoD+SlfTEgvJYoTXkGvz2iYiTtSeb6JtiFPZgMQPH1txTN
pEpY3SwMzgAnAUc2YhMYjrJUzDpGUTjVj4K1G2xtfzhQ5YtWT1l8VZ5q1KRwLqJE
yZrYW7c3SbvxSWnaCv0Pd+XgkMFMjsrcuNGMsHedxBx4Z2rv2Dxa8n2YevMHzwYU
2W1r2ZzUX+HEIoGZUuwvHOT022zagzbp9mlqyfTkCC7Zx7TZBZmp0PVRKBrLiqjo
GzPADU12+uCWsnSk2u4cfk5VR3o6iP7w4uzv7iKrnqz81YDDxY84wrf7nrSnT0yQ
WD3JR5572ZTz2a/N2m06t56iR0asSQ2EsrhA5NBHfFylr0lr6sofz9veKU+N6dmm
4DaJOCQvV3qaR7WK12Cdv9m5/gCyvUPuCRcjc/avgfudzOLEnn6N4AQfoaQeBtCg
EFHZXWjIqDBa+7LQN0SOuGsau69xeL4OXYiKHOmGThNad4PWUK8PLg4lD2HXKipr
YcG/1IF5kVGmHv+zb/KgTrwxZVtSVGqEar4JkF3UYCbJ2He0U5WlXEoFsWhYIC9+
tN1ilOhRp8b4K2rUgeI1zI9apLb4Eem4kyFS+Jih0aWJWwfJatDj1sDMh+uoCJ5D
al8hza/HBvFb9PLtbT9bL/SbzdFwFxxxbqLz5851t0JUdl4uWNvEPtr4LKmVdoLm
S3VAA+3eHIw3jchvAcs9/AW9Ji1tdvGxpHZCQU9YA0PF0Q0hEjr+JwAAhRm2wLdh
pFgRE5bTANWStAzsNXEcPaA0Eg8/b0nmu5tjZC1Fr3/ZtqE6eokyTkFpAvFvVOKE
laY5rOTh9mHAExMB10+QxfNiDxghogIcL8KTeQOjABI2TRtXwZo62PXx1bRa0aFZ
092BtstUEVObfAqv3py3slWBqXcwzwQet95FkA9WxrwZc26oAXgfMxsyPCde1byJ
B/tR35beM45L1oDQFI7ny5ffQfFKNVsRKdFp4ia7vIOhrH+5aXStY/B5xg40XLAb
8pEyxtTrHuAn1grh4JcmMbSfuy/S4oQealssWcJ1Gm5Oh9VvoB1jSy+PS4/VEXJw
pajPdDpwYacTv7cRhPvCXJ0RVKboffiS4ngmoKGPK227vopjwS5L8PIOzb4ufQby
2KQ2KyWjGr8ZepWxXFuYp42HZ3NFUuJpHyzMNcncJUnrMDyHNm7f8gDmLGIen0I8
6VbN+S1jmNw7juu5erf2Fw1IwyIRZcP6GwhROHZG2rH7h8C672AiMSgSS8gxUve8
mXlJdnqBv9CYG+qH4KTWVz5Xb2GrYp6MhjacH94ptEAx13bpY3pxzCm6NyB5WXzQ
W/u3UqVYlB3HiUR3/6/Qk2P4ZtLMjVAgc7lPMY54Lfkmj6JVOUdusVIDm36E4Hd+
O7OFDRlszg9YpXiJuggwJ/LpP+247RstaN3lg5mFFuAz5CHJTp0uzXk//quw0sYY
R0DNZQWAlk3coRckd4oEehcvUP4kvpG4NH+fcBG6A+PPbPgI70SN23qLP5cmpsWs
gsCen69xz2FbeMz8vYE+Kzzcjuf6mtRnRDGbnxdpwcnFa2mmMUczIYwNyl3Wb47X
KE0hAUTRiCcuqE+fUsD7j73F6eJhnmIOOTfyGaSnyYFOQj+iEfhCsXcBQTSrz1Q4
DMBhDXdFQyEES1gDH34L83ik/+odP4gv+XQFe6qUAIeRNpJMt0+2W1rdAyzJGZjQ
if9YF/1fiQuh/1kTB7e/BNqS9+hkayFta5GDJLjnPhXPWl14jZCsN0IFH9Yr1GzN
W5yXXlHeiR/D2hb8XLLwGrqNs9nz7flDBlK4Uoy4GWe5GIGywSyPpFn1MRqjzoEW
lbIG9rwX/b/c2ihc/qQK7pT2X85bvQUhz7nziefHG23I7xM0MgF7XNu5DlisWfGH
StamZYroJkqfpUDRtc7njMar5Lp5N/OPoD5NFMdLDGMCysYs0AwkQq2bjN1n3FmC
HLx6n12wQoOR5czGfY3/1CMe1LNpfpWWq8NTVwupnvgeE1XzVwV2Plumw7sKWdDi
2i6cBcrCPop4Jj6Z9te/EulzBfVVznNwDECPuoEMcma7w7TeHmAFgAQFrMoYzDoL
WthC52ivJtyYrsrsbFRFDV+fmG/vKTNGUyxalIDc3HxPdeHfj8m0hKHb8QIOuKAS
pUhgty9RwJIckPIkR2DxSSCKMlukhWI+Pnj25s0fjPkx3W/95g0tC0yt7ZRz+uKm
j29iLk2Hc9oG+FZayAsTzeNJisZCyItAjVZxiXK70UxyW2Ht/G6WSJsWU+DEI6W7
t65i6k9PvW0OEZlViiTQIHrdpN2/05iGMEw10iepKYtqYZ1/MUW38idDbcn7utnA
pFUjEx0SmYBuPjA10VnIRF8gtAMt9car0gvMsspY2ftyNIoPuym3S9zsHk/Xp/ec
1AL0xUZbm0l43sk9uOoHCpll3Tt4TkU280ZXiojtz2NkykXpubg8J4cVAodoSqbH
hd04qTNyBilMW5HiYugfoSSYZwg8qpUSpRnWcvj+tkYcP9EU5DiQOVRE2khOXnig
pfdlqR4DTAXEsMWtiqypXe+egigYcYUatyc73f33M7cKtIdVI07ig7EV2LtQ2J4E
ov7ILa5V131InPnNgtXhGyVoLwSEhqbh/rcaIf5wod20JWzgoX/Ur/6EkpFJPy8D
mCU4ulxcFWX/DpoYH28RB5MLRXzr9hhPA9M/H4J2RmbEm8Sh5OUvMA2GaPaaxpXG
IUUeigse/gm+0rxKfgZMLwzOPekewBXyEOQPSrjaQk1fcQEjWTd7+h5OjzR99ccC
b0/pCaujsfSwaCNRv0Ykfty7i1a8aAgHJR4CzwF0TlspmtPFkBPtsN7cLM0XKwLT
Qzq7/Bx122KZWFHdZ5N/gPcbpwnehY318I3uXPlIzhwG8LocqUHdd/MTJC0mCUSJ
c+xhKP5ZveoH44TCeU79Vf3SJCLSE0SziLcZmzx21bzio0GuDRyuEHW3ynSFn1KB
rCZVsirKXc68Pwzb1dFRe4CJN/YHcc2OCyUZFDo2MT+hQbmdr65oyjkjDsDaPK3m
5V5PYAmzK+Ism/tdNhZK5Gh9+dP4XXm72dwIasX1ItGe9dbK+AtRr1C1Vkb64iDF
tyESBXzAnOghVH/Ec1nOSlvYtzJyrfDck3W6tYsrQ/9CQKkM6odxugQIkqRVvZO+
mlGhY2VwAi4Kq47qLmKFyF8eyTZYKXKzaQd6znF5tbIHP51oIwBbZ4lydu3RrL3a
7JMvmIpT8WKfoCP5Yeue1YHyOsKXOGF32zonlQY2NBCW7EUg92pUSHDM3dcqevOf
SiRwdTXPOe1RkK8cAlFWGTB3FXEg0MTNuYPOZSvyGwnm6Qc6pXofsXPQWcyBAV7I
25SPAOeHaJnde8y3juJZ4u4cDCe0TmRU8kAI5IGk10cR1ce2bYlCFBUjVJfG47Bm
Kf7cEaM6Rgh1suPW1s8iuKJHYTSD/R797nQyTMZYPupCdkMyNdtWKBLqWGJc+Bpy
jabKBhse6YM+4VBrooQSt1YlCPwiMBH+WolA6Ac+8RiNfp0078n2+M+8HKkgTLwX
yIAd/9ZJU+O6udIlHgtFDXxRn2MrWFa1oQJRakRUcswDZrqfytjQsVM3jfOuErCe
eCnCM3APgYV43bbYDZOc3103BOdIlIIr75G7kWlpOaOAqAk857mpe1UpmNp220cF
JLjBVjzf9vwj6RZ5K73ciGVxCVrfFaz0QET09XWGZqL/lWCzB2/7hHIoxsCU29PL
FSijD1G1cIFrjgwMqd1bV7GUZYY9crF2r3QZW81EdLvDQ0a8xyOyAUCFSgUPbt8j
KHk8jfVi/anozqAnr7ddW+kA4LmYuACiHdmwKPHLSIdPI5omyMvrjGWTBAIluBHT
xV9UlGp36uumKLYtiCY8gj8lzy8nYDbwJuljWzk2f0+pCEdKPTbsI8gf1JVWoQez
os8MShusTTc8ielEyVKKG3PmohnJYiRqglMT1cu8nRtp1zsUg+pjJt6zcJXujyPc
qrhig4j/EtdaTqqO/fGKAs+n5uMwYSD+1PZeykTXkHNBSllyathPlC1vDpAKWFTi
W/HeDv2rRgZktdJmlCSLusKggg+rCdT16MiwiKKL+XAcxGM3o3ifGGgP1dpmwtzW
dKIq7SLmSJAQRl9dCDGB6w9P5kvpHLMJYyR8q6cuwZqwNypKS+koAlZXZS0CnIYd
51npYMf4sN4gBJz+s1fYrbYYB8mI3ESl00J9PxbXmyiRgY1YbTJXba8IYkPOh3s5
azm4cFrvTn8TOUyMhGzc1SjaE5F7uDRyo9QAQdzgShVRjm4J5Kj9U+CGQBU9ceWg
9hmcrKEzfsXvIXpITP72QTVdEP+jXdU0SSsBTLpV+BmH+xapLe7nsNQVRv2+SWtl
xTpLHlYXAS9a6uVhjH5ez8g5w9UPUuKPviItbu0Svwb05IPVLtSwj10WEaful6wp
cSyChHdT9iez+vfQWvj1aBT9ZBqKG8/MZe/y8vDDpc/GyEGjqqqmrZyZWEfztAVv
x17H2BlMzqNxXIFTcDh/pesQtB4AgmhYz/U7Gt1fUpXZipbogwCPsMu78ueRzLQz
UFIZKO5BT/YQmLz9bAsYoh/59tVw15/ecBi93YeiprybxCXlojvjNg38X+PpTNzH
SGyEw5yUVgGJ4vacQ67vDF8h27E4O94x31WD0ImAoZ1d40ZYAVI/usu1/ghVfWLd
7/oqCbcdCaspXZ7/F8wahJUal/MsD//DCxBcFflyNq2iRjDRaLMV6XeuCICd7VJo
UfKN7mvZ+ulmlm12NFZ/YkZsDbyCBYHqnJhNZWdvJUn+qyepUCF39l2UHrRFnAgp
Qmgtu/ZOlxo/mLJ6zrrpg+YCspbwNMO7gs+ZwL6X9kSrVYhRwQayxpFG6Xte64z2
SMCTBuFA0Gbyj9+UNwi7md2uqGYmY0JxrZWf3vcrJw8/9aeBtfELPJZ5Fgibtv6b
ME38mTRoKWxUkMVgu9ISGt3u3SpkfX1yWcrSbsZ07dmpdobBOkSIQRri7ahB9FJi
qG2BWvvSGlr85btuPjIUJqec434TIZ9kfx6qu3S6NOrNDAOJ9vXa6IyYnTP1SPOD
pmFU0lqMoQR66yhrAqBSJOqL+8KDi1hlNusY9KDT4hBSII/On2SJIqH58Q8pMG8D
Ff00QqIWm4b6Wpr8HAvXoZoMXMUrw5BXHUC4pXyJDQ+QIBoXSd82MQCnGnhStsjN
dL5oqqwi7mUjExQIIE3kQW97WbfjN0GeevCLUV/lGUpnuqU8aR7Js00LOE1oiDki
pJ00d1PqxtLgpi8xlboGXR36HGYtHGtL3e1vK4W/aKmxqSyExvTeT8jio/Sn5eXW
4N7rkFwcaOoL4xDDae4hr3EAX88BqmSWUIaHqHH1jR23e047YzoA3VaBYqDsgsj+
7cBzX2G6x2wMcrgvY3GfxQ20MyqetZa4ngiq8hcE/ljmUuRB6zW9bT4E13K7dBsh
z4LH2/9k918OE95aOreZm5KICBfpzsWXBsjPVItU0VBYfungnWDrXxbOxXufLqWs
n3WMX49uBIK+OHf1wgwbChQyclo8G5zjTRPTXdl8lyZXy8w9EwO1b1VrY7rKmqOq
qX/31DRBdsEh6tLn7Mvwa8qy659sg640XQKnf40Uq2TGB4jab/FUvR8+QL9S86bV
zAuz6Nl9fgsDuZYZVZuCGrS3GbIia1ll2IkezwQYZXtTnwgbjyCWknaBi7fnafpL
9NOizOAjYemw74fkkEOc6LLS/rzLWPwoAwnrxs2aZyf5dKjeD6/iMZ5RIody4QR3
MjvkKAt/R6kUJHlJeGdIHwSlAIGraPpJ0VnjaqV0RcadnCqJis7C9xlVtlUALGqo
D7Z6+lz6MQnCreKIj6ZW60l4HfGl6btHYnyBQxBXqlqfx4VHeSBCsqC47ebyVOKf
oDoqkOgDq77H2prVvr+RymW42+jOYZiHOE3FtaJofNlfXNg9BlTSLt/5PM6f+Dlu
kthEB+Z5PIC2PU2itVBUetXH17pGmhw+3bxP91lp0W/Ub80pl541FDE6S6/OLfLB
CuLkvd0d1fmoJ86DVPpj+OKf5AKZBB13FJRgeBlW8u3PEwH2BO3+SgF8hfqY6O7r
fWKKJlk3Qo2jwqMfVGODHzcw+poxCEC7ne5fbbVCHEnKG6vhbRUYVp0E19gJesBs
rNv1AxP3KANHzDoWthNF+F820s1Bl/60MaRS4ZiBYdOVHGuNZgMnOUHVJSEG2srG
6AMjy/YEjCIPR0tftflIgIiY/A1ChAEl2P8WvAVOYtMyTWoBrx+PJ/65NBOR9wtQ
1KwjUrPUInURwmzPpRs+cGLkve3yVG9H/LS8mbi+OwKoEPW+iFRt3v+PNrCqIWme
eK6QAWd3RZKJ+EWZer75bV9jK/ahFBn86LlS6te9Vfm7jHkrxemP43jKOFwEnxwY
gB5lSvhymeDnOhf7EvZVZJDRAQngLykNR+uIVFnXtr2bBK0amqoXEMxqbfD29eSo
TYK3Sho3cPsfmxJhljIxm4pSUMfZF4TKhCJrFLQDocExW0SZYKpINbsuRko0DOGT
yX67L6ixjxbP4RJNOZoX0yS7uzyn4zzjhlruEu7W6ROw7kXG9aDjgRVbzte7CNF2
8SlSKhEU7mIxj5+jiyrFBaNYkFC1JWqiya88yYIP2pSlCme7cgWWOTC5bTHisBDE
M9hF/Jxi4uXRKmffWPNkrXQcKHaUBkLZb9MkAJjjb37NMlRC8w6LUklbil3oyHjx
g52zSx2OrWPrsjscxV9JkIdtbDSfvpO6k+RIBRHKuYzbAUUuw78OO08FEWEaCLAZ
QhA+PssbcIyAYNnffcU//rpG2EgPSdqmPkxo3s3J0SvQrwFaI+B7y31XrJd1vJVg
uGmcl3BkOnVoYgDekbXrvmXYC5b69BIhu5Rjaizzi5V1nIIFwTZZd9iH/XOhDgSN
q7OgtC+XofGz21idWbKxYo2vYQmUJG+ylbfQY9IdK+BHu9XlgIhZCN8F8thnIgZ0
U5+17Tj920L8bI3c8O6YI+ebB/h3rLCVTQvDIqa9ypWNSreKDUZEopRNnlwvwdew
muZWpslk0Nuj3aB0xGRgMNz/OuVCuCCe9skrJsTiKLZMMOQnCSP6c3Rsu7aZLo6Y
yFA+VVcDQvU2tmeJJyy9z5RrojDxZGXJxQqmJNOlFrzQnGKQZ/Qu4v3pkLdqTXzU
+rDLMBP0CVGKEUhJP0/LtvPv4jMNu1w2htgvRGUrsRQeAeq/NY/fBrxeesKVQiVN
intzB60y5L0SLQ0jPD6tjEvn+AWoPzQtp4zBv9cCZlYOL6XyNV3XUZmgti6BVnO7
4skLi98/1iYuoZRQgYa4n3G682x8b5c+d3EjdPa0k7iAz0grzT2SU8pNkYnQNRhl
pci8/IersPUfvP5i765JOUXzuGmkfqRLT7dKT4aMKUCfWRQ2e4G/KtLrMbsHxKCJ
ikprCsKIHPXI3zGtaODo9zaoMBInQFY9LyD8BSTI/XKc0pLOhhM3bkFeSNr+TrKS
YvUymRaC7dQ+Ih9PZXuIV1A9xhXjVOKmG9/uiYEJ40NzOSM2+cJlTh2znitQHQDe
nPSneV2QUYnI6KumaGpO8Nc/afijW/iVhsy6lbuAOXk7WaqriZrIwDoUVGpXiJ0i
LpW/AQOzwgQS6Ai/cSxjwdIyVtORyx2GMM8vb8BCdAXh9n36CE2/TdM73jP3t83N
Yq4n0mp6rY82GPINQWFAtnDZpq99tfj5XSJtHr67k50F2OvfZDzbGfY2kKfX7ioK
yqlvC9qS0t11T96hy9eqA/di3NDCF71vTSfUn5OXPKqCrlGvLFFioN45kHsUxiVN
0+EPUkwDtZW5vPocccftFgtXI//MVI7bebMvjSZtzX/k/oM5vZIM2zrr0XDHJCCQ
VeAc8bizbsdO4xE09c8G7ZeXhucrv+usR2TXZrhRhuO/JubhnmXlSwXxLqCBTl5g
LML6nGymNkX/LTFWuTc2q7uio2pxVwwYkls5TKWnn2Ocq2oW1u7Wjp6jIyMIiHrM
dsrhg9U0OSILqgxZA1mIG5XYBK/aRXMAiG47rVr+6b9wspk6ndYr0AuyZgyfriQe
RNo4TcdjgCZsrrwZrzuBFkqFVk4Ls1Yt8EbtXik/kdwhBgV6QgN0WV1u+ttwfG/p
CtWp1zY0anzcFO64/8bAdLVm5GrXVaKS2gBcv3y62wKERIknW+aw2LSRp3oN4gbL
lpnii3dq7iyYPxX7UqqDNKJIVF8fm8F0BR5lx0jgKPnmXgcIoxug+MDQjxszCb2X
bAAYgMvQ+HWwCEIeh60DACO6jFesdKlq4OBL6hWiHlRuXoEKOunNuDTEnOauRqHB
41PlzJqGL/z76B5YZq82fSdJnbltqwzBWnAq80qs1PfZ4hmzBIxbnz/6fnxyNz5m
A4eSlZPCwK63vVY7MSyEvLOla0sbdS7vZcBVlWS/Gti3X6HRBQko5gG5uMHmMPDR
9K/RMj8o7K8fe/1xk9uqbBnEfoSsQNJx3Y1Tc3L16si7UEOT5n1N5eeYuFXSJEgo
VFWWUI97DtjEzOn6dkKVeN0T271YhYdcQk/1AvFE3Xl62WHtoeaIK2dq6sGa5Apz
fJlX624qY2isIgf6nUl978FZ4StBVgcplFfQ3afZK5DwuSGaHlvoOJ2/KzmzelJb
yk4hvDdq3rpuC89TpMk/KxzNqItq0eMcK1cW3nIKdZdyhBWrQ/XEbKpBqoplhkq4
feiiV0k46u3NIIr+2T+mYLi9w4cvrtEGTo+SzUc8V4NFpar7U3HMwb5sJehxnKd3
eDNyrM+zGNofNT0TyTqVbe5ahCVQPYOzBgq9Ntgb7MTZ4kY1p8+MR2LwTyPUUihY
q5eHSuO7x6edpO8IfVFDeAdtsYyD0HU2GYvM+JdhHe0rzsn4jnUiaMEPqT+Nyc6Q
ZjbXodtW5drlctdqYQrMwbqJ/kmXYdt76NPS96wjhdINPsR/St/yLBz3lo/HN+B/
njOBkIONPk/AWNV17i3aQRW/rV3fkqV8a/sANtXb6FAcUOoexIKLBAXgVReWG8Fr
sRpkOsxSV5k6ThTDGPJ/s+BJZi1Rm+faCj3c6MPYlVGXJz48bn+6o6/SUM7YXVgl
VcZbb3KtohtOZsOYmW/7D/HXa2uoto6zARK1E8RHWq5xC5gX6te70ZlopjdWrWR1
sHQJtlTnDB4y7uVv+Tr3l/3/DUagWDIzmyPpZl3opMA/NmtmDpP7VpG/Zou4d9X9
62toe+VvKLp8XuOXHdyzd48CC8CE2uc1OdDdpVGnOlgTsv0z5xb72WG+aBQks4FM
62IFxahknHiZvBKL5d+a4QiChejbEnFv09jETXqc5Hpg0V6aP0jC0PxPXkeFbKEN
6nizNDmgyG/GPCJzLsjLqnGRV3iJfydbyxHHtw2t5z8OOuAg2/S98o7u+7DkS28i
b99Dy5pHZcM+xFb66hYX0TxmrlAye/dkuyV7xX63mk196vIlJzaXF12cov1e4Fn9
DFUOZi05TtbNbktsUMxPz/QQuzoStVPPKTyTio6Bs8ET+Z1PHQEyjBzw0lsQ/ZBz
hOnGgjtW0KPnZkKzojdI6jPZDjVsYmk7fiOOJYOQhwzEY/rT8LwKI1+9k0VEi+kB
4+ZItqI09TXX6Oa7X8F9/IKdPPKYANCIl2gMNWpEL4TKno+42dc7JtxPhXph5ldf
imXIKMl+tf4RBNPV6s0UiRtL7i08jDqHYs/yZbdOfwvs6G9Jr1YdYHGSRp8PyjbH
fdtkPmvP4fUKXSRb2qbRKvSGstMEk3rRbwsLJ44dpP5JoRkKRRTzbYQaaYTSjgqO
LvPWNjQHxLHb2GT6MRS42MwcUSskK3+/z8WGPESKRIPMRpCbcaHsQsTMb3LGsDco
bkpmck4S0X9UOixAIEqcw6QAAYp6bgcjC8cJyf1od0Ec5Z4ZXhpx8t466NReKueR
uKaP3Nl/bl2aRiLbv0n8WyB3eVowibnb8Zzi+qJ7qOWAH3lQ8e1T/vralEQpODvA
//+n3NE2ugIxXl0X4YJ7V1gtzmrhoUaEs4CmVfx2n8UP14vydumu1SYL86vmXKET
2Ik8+N1v4plzN+CLh2Pe0JM4AfUrUu4z2GI9WhJWD9K4BXjGtc3cQbtfmB3xue6U
bE/dw367mYFAgq/UTyK0ZvySEGCkwk8XIT2LA9nW/taqGkWdGSBTLwdExtx5KBXQ
DABP1LRLGvNAcZV5VHI+0lQJOXLuCSP29JD5R4PnKDZblpUm/AGDR7ha/Q2toZ+p
Vt+DgrnRE7dFZ3N/3I+gc6l9m0OA8KeU4AHEhhoqJgOjZeFSFFxC1R5+AJ793Kjk
xWPCLYej6Fr+JBu914Miz+JU/EIyW2fMkKk3O7AabFgzqbSar9Zr6x42pOMVhzW2
Nek9oPHHrIO4/9euBlCoYodFefS0op/syeQgu9JJJuD+hQCsmp+gVE4GPbClWQV4
Q9xO+1mW3iJeoWOEBu5i7GtwFQ1Ohd8d2G8+wDdfL3HZ8C5daLdnTn8Qn/+rAO0E
i30VM/k43iL4lDpuVWsPft66NmsTikM/UPd1Ke+QcIn6rAy4/dN1m2ChGL0hT57a
3xa5EZMz34dgfX+If6zm7fQgSOBSHO0HRDRKplkdLLeduTfa1BbM0vU+NcfWmzyZ
6IQxOxIz6vOLQYVUU6Ix/7rR8b0oAHRXWkaFIyrXmWDu0g3y6L9TuD+I7Q0yiDrW
zv6DtLwWByVOUeOXF9xj4zjwWNTD0aF2LC1lQnP4tfm8P+AYOXmOs8kk2UTo6TZo
Q4sXjsdPHOMaGY2HS0/t4bcUTDIxNrHNw4TLUtyFjJJvD2jh8BUtWtJx20PJGCPz
Wa8eFSajRGtFHuutNEfi/XlZPlXIWgd4558S5Y7JC+y5HjCNuyZWmtwLXkixbPur
Mwi6D5eIkrhsWY9Ip8GeSf8VWozpv+H9WVE/UsoBuYjOLvgSWNzSIEj8Z8amJ7fF
frxqzowfITnjcnWuNR54NZV/WgrqhZ0LvcGih1dMrLVNhO345Q8D4nztw7muGkxl
k/16sShKmn7c1QwunlNCPN9LhIGVziWBIqECypGFwbkTWUFSBFGlhFp5BQYBkNEb
tZ9LpbJVbqtzPqdVkHRfVyA1SrxDai+dZnwXobV3E6L+1zz16kDwRda7JRaNsfqK
u/7XZaNZX1cDR8mMdCKNvEMTsvvml8/qzQdfsmPx2arso5EIQonLW6AIMTTErMVd
CMbxoBdyj8kAaGslZRzjG+kNPFp+0ym1wGjcfyFWDmxY+ZN04KTCN20pHcZgNJAA
jEu8FWn3GnnweZqpe4GN3jjHP5gLHCBNPNFQxHmgHZaadd6+FsUANccO412q4pDa
MhrssuKEy+2EM7g8ldbXZrOpUBqNu1XZW+nRoNwdq5CJddyqOx5+xnTop2kIt/KA
qZQ/4HQd4bq8/wmLaS24Bf4omoyu5LSBH1kCqk41mVC/LcJebxHZZ6Y14O3oyG0u
J6SJdnMi+viBA7Lvmk9De7Ghi7Bec0gOE4NJxrz9l3zZ4fa2yOH/I5p14RiDr0Kc
wsBPc87TOxlQytDjDbegdfxaqal4Uub80DANW57n9nRUMPLKCAzfoejZcd5xfcOP
WHs8DaP9dEQLh4Yr6CZSKn0Pn/ChYnuEkFALbwF9n9fP1Wd67XJ0lcgc9et5B1ao
NIcUWgEdhiaMPgzAN8/4RS6WTCdGZsJleD+BgQq3g5tI1dkzJup6ka4i1nlVW4vu
NaNNRIHDtTLZtaXxWnAtnxkUl0XJgGcqHA11Qr0jDMxDqVP1AKLAwX512PzMEvfn
pADyemONw2ie+1KjRiEfSa1qaFqODRYZhtxA4n38RjKn06yLlgSzCmEflyZ0gzuQ
f8jt3cd4AsUuqvGcyfU2VVvyETx/iMEcGvjxtsMwuZOT/R108fwL1l8YZWnYkXAF
70VZMSi+7FvEQW2mgTR+P1RepwQb0gvMUFuXR/cYHaUjmNkoZpgLE+7ZUnHMc+iN
XEdQujsULQ+B41hlSG0yB31cALAvtkb6vjY0Hh+yn77MJqB+0pgEKH0ssZ/9MeS/
TSXa2CWTlQSSemCYIAkQ/VEnPll52s1VS0lr7Wxghx6J7Yljr7Lh3amHx0XQLdCn
pQa9vWJAwHgtH2W69ZRHSQV52tuNNAAjuF031rOvl5JKcRacd4S64yeQ9OKB71wA
PgTu6DfiknyD3DgMN6Vz5103OSJaZA9KNFswjc3goFxNncFUtTiK2n4a4LwZWSC/
fl+k7BpPZ+Oa0imD8Yf23EWfHXv8rVV+hseWAmyecOTz7OtD/1jnWbqoqES+vjmm
dOblVeRCfA9yfDZqNdLWjghqDhEiJxHYpxp6Pyod+gyCMk3/bvarcJ+D7pxEIQmy
SnP7AtX5HXqQPPOfEK+sxSYdxXLdkrEYsQWooqADCLpJOfTmWaqevndugGUCYklo
0TCAMHH3jZFrbfNGVxUHB9IDIH3ZhboBB6HqRjL22erlmCfVIf/A9nFnqPZMjalx
2tkCr6lZt0ihIjcbU8wLP7rpfJVkF9p8pMWF7cz0l2klMv+JewwJrKjS4Dx9q17W
DpZVAe3f4Ueg9w0Mdu9Et7ZhUQZj2YplaP9yR2Nyjng0m3zDMdU7boyGk/SRGvct
Mbl/m2i4xgKo08EcJkI/QYp9ejWronn1sSGXeU+mtHxU2Ueh/TcZyGkv8cREM7a1
xGOAIqaalGgEA0Y/iESYrSHONLIqZ1aKas6otFT8E78h0iczrUXauYMdapoTQ2wI
OpOMB5VtH1tdxXHfaiFE1ZrWlVK2UGH1LVCQfNmipdu5QaD8eR0D/WJNA8dMKVt3
4IfkTEwdOSN6hv8WzWejljGXNPcgf3yRBQ9x2qTMSYX3zDCaRkkeNJa+y5kzPKq0
+91oTBdkdjjt6rOTNPDbwtf5ZSmJ/ELYTdmMQdsvN9ncZFnr+IPjp8Vr7dGTMPCq
x16AwuNHr350jtQxZyUEnyWBYHirDCchnKLOoy3AFJIzEOKSBlptoFDH1lw5RmfH
70kWUtBReDeN3HZEfuwI+TAxlKqPi8nvebiITooa6OlzZWWHCy2RWNSC/Dq1tG5j
JRNDpbqXq59d7iatCa/ZaphtKGhaxmv9mA+9dyUGTJP9LDPqYTGZvKOmbMreZQiQ
Tse4PupAhCqbTRajrrgO5GuYVVtCS4Ud7zggmXYSiFvED2O0Bk4jcIQqE65AS6Z5
jkF3OrCYu8SI3Nq/M8A1wnOIMjJtvnBDmIxd7JDVE6evSxyias9t3SuB+z1hn0Ls
nNJ3lUbc4nkhLuH+W/3xSnYRgYZudHdsNYWvZBmpFGyYysy8WYbvHzUa2fpVyuHv
p2RU2V2FAhUkOzd7HYgp+SzJpBJ2I6Q7pCWq1xHvOj61j/9ILgA+HCEcKWqFaNoF
ZBB3fi6yIVrjXDsDWTdrlkgmnKapMURKuvPBqrwHmHzsgVAmVPzGGLwuoHDjeIbJ
wGtY2d6gD1vCC+LAtiuNYoN4UkTaDDrhfy/7T04TPJHza054PjpLhz2K7LH55oZC
UWL4ZrxNm6lJfEplW0x8PAaotdrbyQ+Fhsk0ZKoTGLCdRUH+OI0HMf2ZxOAi5doK
5ZZIw+l1krhVW+OwdtzZ/5O2hQFAPqXe8Ay687JtujnxuLM41X1QW3cr0DGxkRX9
b0CtRLlNM+wrXd/7/0N7oy/UbDr3Ses0HSLOW73NFxyg9RQ8BGAGBKwzp+Rv1iwS
79ahqcWNsjnMJHDBh7MdjpfY+MLqtuYj9CRS4q47ANnrv/QP5jrJiGRTJFlxI0B0
dSMEHkAAlw9gRSC/iP83zGQEmmL/COVIAYLD8VHxWAYozGLk6d6mr4VDTMAoKp4m
1CLO5fLNGhcBxNzRJM/9YyiLhbYwWD1zYxcP8u7+YHNLi5m6rFhwJ6ZtIpGTmS6N
qXkPaQQK6dYihgs2d8ASRmi/6kE3XbkxbijQmhtdqh3B8r+B+wvpL6TnHiSt9A/w
NFb7M2nE4kjPwP0Lp5PrUkzdK3b0vH5I+EXbYy5QyCv8zc0Ptp1jDJrejRmc5QfA
vDbvTpzdU6sdbT+L8x8dy6dg/iPw7bG3J/E2CvRFpjhZ8x2ZrpnyWnssVPKTlJP/
tLE3Ij7qKEvM5s0hQHSVyOuwoDbDFaujEFKcjPTp3H6BYmcfbX2F+gOFl6+y4x3W
0CpL3WOage3ma0N9Ojj7MaNSFbrNLTvvdxGTBt3Wk74SFwE6WNDuoz7+Snz4m430
IMRhcx1ZXV30VyxLMx+Wm5ee58Q4HAZO7wDg/jAwVTuaUJeo6UwMITBbl9Nn+5JB
Zq4DY55PpoIuxUSfcUn4lg8W9s02vOgxlwHCCVnkWbmf15lbOFZzBLHuJ+c00M9c
1rQGXP1cYkT9EVs1asQTJX/o3vAnwJXrDmQZBzMhpxDDoxCuLBlSgXY6SwcJPX7d
ORsC2008i5vTBT89nxzVedmf51vhpb2oE09BqQOv3V8t+8zIi9wSWEPURrIXTVs1
tzlDNmAzr2iucBcmxO3R1NzOHyOMFaveiuIeSdCZL8a6GjqZXmHuq4oSu99eL+w8
Cgw5+PzoKglaXafOGLKD7GmDKec8hPmxM69++OI2J0iecs0kBuwtv13AlItpa09K
Ugtvmzp+5aooiuLG0JTc4XUQkIMlTSJaMBlDIO50ipUsnzFHkOeIWibB35tUoK6I
9RvihchZ554knPMavIaiJM+39lg7Wria7y6PO+85EDwAH36ENwxTux75Bb1qXIQu
tIw/CrE494rHuhjXj9BanVogA7aKkzNC+jahrvFBAno1UJYtRwhK4Hu0AQzwDvaA
pPaz3Aej7lJLiJXrDmEe5wO2fX9YdYB8JRb4Us/Sg8UjnIH8AuQBzbsFmQ3eyYIW
CtC9yrILv+ct/1s/Ij6+GeyCXJq3pDfXc7pkSY+jDRQoJDM+maBxhqGGkYU+//e6
hgKLBV1Qai+elCyvieDAwMwnu9+zG78NMWyVKBYPRChZCI8CgSjox2MEkcWFGu0a
/62TeDJdO0bfHRY9hWng0AQPMkGDHaeO71g4eF2LIUMCR1O7sJM7m1QevN0zN1lI
RbZQ+u4X3uCFB0zCfwcLSvbamcBAkJbGWb2CfjhuwkJzjflFRE6+JRTtZpgrmREH
PM/n/g0c/Ff0FMO5v8FXa5W1QGQIXdpwQzQ/4hT8v2Tbub/VuX02uYvI6WY230Rm
98eLi/sJgvESHC2Y5d88x6KfSNY9VgAymzbED/sYUPQbkLeWbMFdb5m+1UBhQ7TF
o38DwApz2adH6V9hgG96Tawj7xeEtwfpAJACP3v+aKetKheZz2C8IDhNDgwvO1zf
QkKt/70If7hC/owvWPynY3RuhQSNOi63DMg1fNjNaGV5uooAhs4h2KOOsX147nuy
RStqOPqxlgQP0Dd9kEPjc7Am8wAo4Bc7QCUSAhYnTKyaxiI9ykMoTUjK86fxIRPg
2wMK1YHuTnAcOvE12EzRkCDR2r/awncmCnpB2dw0dOVhI6LTuXRYA/lz+HSTfrV4
AH+iFrF7liWmUevOBuQQznhdOdkFN+rOpWfhr9DfLAG/dij0g5vZNwORsXK1AQcF
2s8yqXZ2yd597DwrSw/exgDDHCcs1y7vYHFsmHkY2UdqwhrwCjl54/et1bPXOjgM
c4cySv42pL+WBf7FWObxs1BICjLdRwQEnIWBFDp1Q+VWlNIFvm/WHXJdgvo5gDby
xPDMZ17jizS3zH5CEl66RIvjLGMUCcVG93xzcHijXn3bsxa/5/YOIFV3M8J9Mx3k
EBU7gCrquHqVUR5W14zC7Z+FLKDXOwl1FGQDE2mFle122hS9AXbWpHQlMx+aBa3e
uTImqBpgDWeiZ49ORmXsQI4J//uS17gk4D/iaUZhQFmwbykpmTWLFD4K/sBWbSFS
qBYbmVDqlZluXiX+hK1/qacwWlj3AtS4N5z3J/wogPgIz9XIlR0btjg915J8gAqE
ZtAfu1aAgntxhJdL8ZIr/mT8TJdmRMLLiOMaYjLZdEYsLDyIxKLdQi+D8dszHN+7
V1wBbZYC4SckN6oYMd/STZ1W080vGt+UO7Xk17ds3C6JcdOd7W4TGFHl1Ps9Y2G/
vRNdm6n87SeQmGxJc/7/kY8zm52s2FHdIeP5jaG3iaazNEosxubK2ioo/Z7rrQNX
gFmtvxAT360kznNsUsRNYQdBjXo2TQbMw97JdlWcNs+PVCDdRHiZGzkF3zS9qFO2
uR+E9Au2Na1l6r738zL0bcpyEZ6si9IgNzd8/OL59JLjrCQkgXt/JKwUrGcByUyd
9x8PfG+T1c/jKlyEgxvFph71M6sR3r+86TctA8vIicdWHXhN+63OyEcsxzDpA5Z5
FNBieZXDO+XPtrEb33P7FbbpetiU8Fwl24+wOREGpCJJ8dFMkWU428QRqvtN66P4
NHEt1f3iTUQK22Ha84LHjhzfZhZ/K7Wz9fUsIHUtZR1y/AlfgglcEHvklCfT78Vz
nPrPPDBFoWQadrvwUt0ZejJlYUCb89Issm0X2u5WaRMPEc2ry5vpNAKjB9jKx26p
GOzMs+eKhSnywr0mf6EXfy7VNDn5Sak92IVlyLpdc4fXqiL+7F43KI6GYHMVszx9
mfyLpPUmuGXj+EiZwcPqkjsmBUoLUCElcL3H8G111lwRL6k0JvG+vJj1eWiWH6jD
/XVAdtQwsh45jwTYWbPAMLpxL0/pI/s8JQlYu/QFUz5imC/Rnn9yF6zbbwTpKhrg
ZdXLbHP+N4Bp34oYL89zKUE+QxapTQb4HapRvR/S4XaojMD1ExZLwapwIu6QQne5
mji380dYn6zXnnpCdAUIe1eGqzYQDgV0Wesz51QNjag753TPrXfFOr3pI2/Yu4ZX
KD3sslMEycQHqLbV73QkIXz//tFQWDY7iMa/ZED9mIcTJqjddpShbwB9IE5SnMMs
sIQVaTQz0y+aX3K0u97LdXooWPwsgxHS1DVxPWhHlkSdcgA2hP6ogzjTICi2eg4C
GZ8H2PL/MYTxBGN91JZIvFOds450283m7U58xhBWaBUO91ymU5EVDCYT1zUyiWqR
IZmIXC2kB4G7Lt65/MlZejkOHzG8BaK3HUtLyRG58aclRks3qb9GAwpAbumIEVrV
NceY45OkrgfK+TQ55Ho+VnKJuVc+M4ItGilUvbFVpzrSUy5weu7PvnlUbyRTDeGz
ezgFgxcFZTKMt0sqp9V+G5JK4W15pyVvqDcebZ5wAd2R6RykSk9Zg/wzPdTB9jh/
BFZrjJ3RW4seAp5tOyWk1e+1Jo3KgZXia9/F8wyFeL427gyz7HUvhuDT5EcbTzFR
PvHrBmJDeYplAv6BDe3YIDBB0wFxVQgS/chrEVULQu6NR2YvGqnyne1DIijIypVF
L8z5R8WWFB2xTuRxJDK873Legt+oR3rJEE3AnrYSwa4dK6IOAtDdZwI0BXSwWr6b
7TIo57GKW0+fQfuT2pcUi3auoRxp6ONhn6pKqey6idRt+Sep/lnN5xejE4gDMJk9
L4Y9/QIclNoW6OJFc5uQ0BXlqxv3GB0kQBlpeNe4iPtXGEti2MECk+MGuyVWhilC
ytavslPByNtuPM2+b2g8JYw1caNJ0SzAoJhDjuEs7NOiY3zAAVyljvHyr+Xxwutp
yyRfbX0njwDczYG4eVRovB4ELq32gzFmLFMhnNd5INFVGl1cUvG384z5Y+yLIFPU
j4K2cz5kZG70k5GJ2M2sBmn6dYSkJ805mo5YqRfb9+g7SnJbMKVSZ+z01cWKlUgi
8yXmih0YucCaUgb6K/nfW2vXZOOmdcyV5/lNKYgGZKZBSZCseV5/AEhbEBjktSvr
Xy/mVocsto2U/ERU4lWTEVJEHLLH/tX7bu389VicUWOLN03Pn882oOvwtJ9nu9p3
foS4L7kAv5MLn5BGd3R8DLIK0yXOvk15Xi1ffyjQdyakuit8v4EyMyajhsmgfRTC
0/1k2Rn2ZcIA0qAhx+woXAUCObseDwCWSw4U50QJDnJ4eS+tV8ZWFJmqoni3keDT
zjW8Wf0PxlpweXJk//PtivDwSgWPQr6rntYcmnkUJR9AkWGYiC5pkKB4M2XHPT9z
eTHIr0wbcg+e6EHrUETftH3kAvvCHVAgKcBBQ25LtVHJ1g6IxUw0l2DVJH2DRRne
UR4rRhB+gV9sRnII4KeXD+twUh15nb4Dy/8/nGDvZl13ftr6i8qCJ41EO8YT7nYk
fgCnh8fL+vxAM6vzMJgrKkUPQcM16tjpnDVRdowEKcAmwaapSYwEZMeEgkpQiZ6S
Jm3xQct2/BtJhocq/dopeVtLG/57jH1/S6E7BUHolCe1u270rtrDX+18hkUbuJ4Y
QP3zeJn6zjFVMRSxYq1RGmic7nq9tQRy9MznJAyGxJQRYVLX2G0K+AUzCAlgPHPK
U4PO95KV9o1UqWeyNZAlu6iEgSUvZzaNvsSjbMdjtjzwRQUvdiiEl3iEV2VKqTmp
GXQ4t5qVI7C/GJnvpdD4HbtVwIRk6DC+jOxJGlcjPQiEcLxkZVEXbHs4WndM8Wdk
UMdPCNu6MT8gekHzgxtZY8+XhDy8cJD+TMCDl5rqsC3MYGKsaHi0JRz3tLndxrA3
Pc3nq6c8KHRUfroVHL6AlCPnomW96b8IKeAqk7h8zUweGKJbXL4GAOQYUCSERoe7
jgJN1qyZWeMazrSTY58N7aRqZuyi6RTRYEZvan0bfyBjnH4h4mGWjiO5vp0fj4wm
yffHVCxn6x5ZNB1jLVT6KWUJKG7GE87eq1gYK5t109A3qdc3uWr7dluO+QDzgjNI
DeFz+7enGYf0ILXI1XkAJRmGkE5SDNfSgZMIYLfCJpfV7Zlc5b1RdgNF1/sS/vbJ
yKD9xKMmDJj6tFqXx1AlRZ/88ENMTTD7CJ1mbSx7yxYY2XFO8SMCNVcBD0qQVqoR
TsOUxpuIqpsNGVAaah3zGjmjbTQDlF/+jRxnx+0ubCnS6PEwiJbk6G3oQqutxvOQ
I2PEWZVfpxsPY31ih2KJ336BzrYzfCslu3nelJ55DtyZ1VuqhCJXEfpQD+ApHPyK
/i83AsXlmD+rDr2s1l7Lo8KhNMxuRJ6lUeByXObimARo55/YKQywOy3/DBuJgC2R
RDYC7QBLk4uZZAAEzkMEWMdIW5Hk+ehPanpTn9V4aJd2WYEgnFgUXG1Kkvwmb4b8
a03PhgL+UA+Mn6PhfcAQuYS8e/XF84KODk8tqaKuMYWsS76fTbJe7PHPUdiQe+gi
3647DhzIBBb2tSZAfCGHX1KVwaVunJGcuSafjXaowHxwuoVFgpLhynFJg72jbNST
ATBx2oyoOQvQYPUz7C8CrtWCzkFUkHVt3s4LQTjr+xebw/kqhL9592hrsAhBcCJD
t7sifRPwEVbDpeLfe460LdgSxfngS0SOaN3C6ttPkA8TqzIgG1wlEjtA65eoKyY6
VGtVnNGFFd8P0Rq1zOsp3224KfG/Xiflkd4Ly1BP6codsKNdO3GDhnGVgpqAwT3c
Q2hKf987+0Ksfik7+r1ICuI6KKjxHIIwT0DytcOfchq23vgDmd3+YHTVHhGrx1G2
vSw7PJNavAvv0ET8a1gPkx5q8bHNROTh1HKRKbIydWP0a/AFiQHK+ESDzZUL/coK
/FiGvwvsxOWBqtiSKbtvysbbrsccrrLrCtCiTegGbcyU4HulMvJCDFhWrFXrCsvm
2WNMFLfAyBQ2f5TVUroejW+38wbWomVmLfZIdva9Ud5Mx2hZkWhguCk5/ipB8/E5
3njBcxgT3ZksMaInvYvR1v4AGCd42n6DIc7IqXKj7tv7PfsOKsrUQKRhrMRbFfYh
Nt4uh0HfTwRPhSyzfJQCugCl/aEGgejUEjtn6R3cK2jroKbJ6AN6SccEjLRpsjM0
JOEO4zHVT8Ft8L39V8/EYJzMai2o/yHH3U+mdbfcpz9V70gu2ObhIMxOxS7NbD/y
PIqnRluVQYWB1Z8wfwBvKtSptFUBcShLiEmPoTo36kreDUY0bvf3peWdTmxb6QuQ
sj+JlSXO/In0Sr4Z6dcgtBfIPR6YLwHZpQzhhj04cI14Tj5OEhBtG6ZUKfj7MUvE
xD05xzSGPovgJ7GKj0CMGhSTNkU3xhXLjJu1cuaDSavKTRdEpDlOEWjQbu+Lm0Mj
2HEmW7KaoifC3mJDt2xZ26ky8SrKlm1QnfXgxmd5/IP0BY/P29hDyojcWEholPpc
7Cw3RZwbEBEyOMchzZB3zixWBFqunjHByB0Gt2Ffa2IOLxGCxgnhJr0Vq4Zqesfu
INURr1LmPCVt9jzxOVamLkkr9u1jMt613DgwqPc+WGgHTMGNY01ga9Ftz4dwrhok
P6TNkg4OySW9DmjKULbDyUGoxH7rR3Lxkkn11MeaFiWGnCau0q4jtVdWWVJMdXhE
jwfp+jfh+1NMMgtkXmwcAVgwBb66OXWuVjKozCpdamKLsSHf3XfMJcMLkCoF164S
1XXu9MiLI4yqbX3kRD5dUmhCivDQioTN3GQb0WdnvYUQXlrQeRuZjcowyjZWDgUg
eolmVSoxoHU550u7xETcvvsyU0mQWJg9/PiGvvZX0A+XbRNk9Yn5FUhsVRFi6o8O
JtsdSqUIMu+hfPDt0IgsjRbEVg2YQ0rXCRL+FNkRWaxBWX0IZL773YQ4Gwun2pp8
Rznwwo3yDOb+NfaIsdlRm9eSwFrhjGEyZq4iNx7c7ksC3mQPoHz4e2mqj1AruJDv
9yniML4Va4gzy3t+9ny4TFpxEw2Djun/IYurMTn6q3AtlHIHmlSW/pnQzbjjhz0O
374kYWTRANL+q6EvozOp3Ah0hRK0mxGvLb35zJCdF9sy5e9m/HJ+/uiQnS5zJHwz
UJw3xgTMUj8UEUqDA3txmYoGAJJHlj2DIVqbO6PPYtmRxkwxGFsTDIIVycakJOPN
VQFydgxIlxxFE4CLBuRYuzm3Mj7u7krBzsYgQaq6kT5GPdeuS+9bOCYKvWLsJzJL
kPC1zuWp4brk8iinNqeob86VuZDadg6mdmdRtCCrW1q7D7AXBM1lKuLFRnqbf7IH
5nUX6+51J/mEPQkmWCO0s/M21afGBD6yGueS+xNsqzkXASuE1+35UDWxf8SrVBKY
FYFLCLcX60bAvtJ6qGJwjfCWA8FAfGL/RDqWLp4Xdc+gZW4riazfphwewrWirIiK
J0QFAdTGX55LMKOSfBVuwhma4xhynbcGvKgjRdkPYcmPBUpaEhs0QYCVEANyWB1q
f8uxjqIevb6G/DpdFqLjLQvzihVKbz3SIYGGl/Qrf0Ie884UdQp7zZhKoyQWS19w
EmizdYlPIxjfn64WiYrczdWAGOHeM9cLgd1PldWYlgtPwBv+fTXBuIXn7jfFKyh4
PyJdcX3GtE74xkUluaKn2N4XDQ2Iovs19H77ykuf6UuBKbEcTbkIbmc3gTeMXQ/s
EkyNkiiHJUpGYmzT0u0oQOAHGOeYDyVf74YlvHIoh5bbim7bAGqpZg5SSAB64KxX
0FEKbZl2xqCHZQKLJ3wFSVumFxvEx/FfGQsnFn2ZJBynC1LP0pLt9yovRjnCmuQ/
3/t2MT0I9xAkFaED1SCBIXUOr6yCEQNtei5MHUXP9VuBXHbU9BzQMWT2rgJaqBMK
oVvoYQZiAv8bQxQjtHns0O+AnRxKJZDZhTBgeTOtXf4Yco9l//IV69rBecXhUbyx
rlaOPdC0+3lWEbQjcB5938MHz5ymAy6EQ6sPjH5Xo0ZTr7jnmi8NfUTbpVtwO0vk
GiLG/yBqOlOPxRVlBNfJ9ND2HEmTZNbyheY1BWcQBAZqICfMsoUiRoDEputvu2k5
xers9gfBd3uvuwdz76zu4KGJeK+r770Uj1OglXRe5FA9F9bUvoSzPHPq7aRatVrH
zsXNpWM9kXc1SoOfIzdF9BGh2qXrH+uTNa4BPhIWfNJUGPkGKfBun3jrtDYZ6x//
YNpwnSVdZ+gD9jFegw79M4Sxqj/OK9bc5kwGr+J3yDJdi7KPLVtfkgu1+zNKEYNF
a9m+0RPVtSKXqMZoa5wfH+f1T4VgdKwmzLYngThvzqGCOqgfYbwYTBu0w5+TF7hi
uzEZY2eSUgI5HmpexsU5Jy78tnr1Oh5nl22Rd/xzNv7Jg5B94vrglbQQ8EUNdxTH
Ye0YyhWVq+dQeGBjJVjxrtFG4x9Nl1wdpiFlMlNDiBSAbNu142bJ7RERr1rk3pK7
ZBA7HiVpw0r5GCPInfKv5TKDHm+UsE3aM8/gxRdjBVF5KKgBYvSqBgr1tr/rE1kS
ASEcnuAcE+t8UzIIemoB+F6wUlP4Pr3JZjftYg2fpEdoCAUNxWTVkRBiosHUznoP
54h1+bFk/IwPq5oqz0vihQyETPN81ujPqlO3OrS5KATd7ycpvqBFPJSpFF6ZYgz1
H/QuW+obv6YWmx5RQA6TCDfwkzBXPTdLMxLvi6Wg0utkiWKOWm2oO2b4ZxJHFjbd
gDQLWO+4bhE5u2Z9vlvBOkEN0s8gzLF1nd3dV8prtldPQG6v6qzr58qgFczMsJmh
9eg24ZwXkof2x+CO3EqPiHa7Xh6l2OAsh9pLwgkygw9fFZLS0nCM3Rl+IetXuD2C
WmYSI117AgRDY88rTFK770mf0k+oRyOeptsTxYR+oGgNk43yUbr7kzXEF5jfeUK/
Cln2zPJ9m4Pmz0MuBduiiVLosII8mwgypASYSD2KaBl39g4u7CiwcAluJoCQYAQU
WRc9gfPzTLS4rQjZ00stsM9s7zwp2MJB9MZrI02QYvV7HXQR5lziRiKaqlnkYO4t
kXcLSzYbmGlJhUl6h17fLEcu7w+AcYf6MDlpy6qdS9/pF9CGHEWLb+m4dP3m8m6C
gaEYGMgGHTXXwwKDniCIjrcdTqOHgBEB5A6nmUqVymrqzfayhEpraHOigfvGb5h+
B5v96jgqDiOcrRCi3trI31UDFaXi/Ur8JnQQweTDL8/N1w/Ca81oj+ZZqXkVMmmL
nKqePXi/HBfyJbQLEHOjsEghUdEptJktoRpwLJI27aznLiqbYQ9oARq62T7i5GBF
AOXy11MABaF6CRRNt1ITpGD6mX8kyyDvC/hRJQJgRE7trZ/0deu8mD7QA6C7h4DC
liIsf8dm5ooQnRos6ESo+fB1+oSFyhgOe4NCYwzybupiXMLPtEezjXvqRxYDNu6i
1f6rmAYqUwFF+BarKW96ri2eawWatmmv0ACgrmjvmRmsQUz3opB2X5/0gZgUfIFX
Tjnfcow8GVSvi7S/Ws4dbhzwqkYelP1eXNgQJcVyAmlP6e+U2XKOMKIWO6G74RBw
X4c4k0hgTN4TG20V4eOUcHX0jueuXxRPQXXAkZPPxTvhO+C0yMKkAoMK1RuTC0up
4FtMr9OY16RFpiS49ziEc8M0T2OrLKU93ZkgC9t/+RUvivSMRDoXBPq3GHaYNLrv
qFfQ+9YSkldkAfx7Zvlce2ymXsCyy8cuT+cEFFYvg3OEiYw9CpxKZHcIzCkAVrW9
Xt/KAskDFs10KSx5VjnBmZVCgnhSnb/5BsDQ7i8T4uraefptG895yJtaPmKbFsKv
qBIgr7+SbJV0i9fix7QWa3QNxGv6P2C/csFfaVQs/2HCjlsVM0t454a2kN4gC7zC
8OhPg3844mPK09OR6X6LUb0W++bvzS0kRmNu9QrzY/dtgQFfnlipaEux3opu4ntm
w1ZWyY7ffTaqKS9Ku5v/BzMBJyNTiADr24nJWhVSwKQEx9u2zalC77d8sYmGUAfU
GZ5ttuo37WbJWyAGwXmKHN93Nu2i2qQLDW82Bau0GdD3xOqns1MiBljrAvmDQB0y
81+nVACL5OjAzy70allEWT4TdHErcAhgT8UBaB2E/cdRTOlSbk3xyYPrnakjz7pt
298l/+iPO0DLWhjobE52AyNOt92z073d/b+7OjcUOsYzQ/wLCpnWcXh7eurd22Zj
KNh+NtDb2R/oUAeBmx79sPkcgGemBUMQvrpLhCq+uGcnqolZPYE3CSeffGYriVPS
IwdFlybsMaz9uYdn9keyWF4V/AThGorBjj2fuDU9WdXohQptsQAXH+uf0o/RkG6b
kQbEFdA4wcVxIY9HxwEO8KBhwk7fC6lBV9FEnxcejlZ0woMk3e519FBxukOPUdSU
0d/YX5CNzClrEY7tmbCBdjaW9yb43Ki63t6QvzoW3ZOGw/9t3KKpm1Yf4I+GGeM6
syDrfUAEaSWOH75eXtplyinL/PlPR+SSgpwrOxroS2DBj1km6h/ZsH35gFIhHg5s
Uq0ISomkS9tX96BJ3B+WuyXxpKY9Agyb0oDRVVq24b7mvM+hCvx+M9QrXUaDU/id
sjBOtIT/BjPV5ynqmvwZ9RG2NOpEm1mOL46GGEgnROqJWOqo8cpSznrV7Pfr6dF/
A5CrUqhwlb11c4rw1hJGEvfk5q64HQpOq9aeHI/LCwwhz7p3QNVnwc853mZdDNTG
V0/Vg2WEMf85zXrHPM0S0xZUrh0wjp1QrF4iMr2SKVkqT57Mvl32Ko0eCgEkz0lY
iuZLeE4njKF28pAW+TWlrKBOz9F87KQpr/DKvCUs7eZbExogG9edL9kk/PDPYE89
kFUtj/v3dTgKtuJZZ9QKpPV+kxJwn3RA3yC3DBiYCiFaAe49JZH04LyzyTxX7O8y
1QLxol5ZVVIrrlz832N2V4hC4ogwwmojyw8r9xu0qxD3ldXj/5E5GA2BTiYmCNfu
SgaJFTxPU+YMF4XynhuQLt3i3Co7jZ20zujgktqd8K5GLW12QLzGrNzj6oNsIXvg
VhU/BKdGgAihRNZkUOYEJJanpIv+UUIU1vU8Hoj6AGp5k5lZGhkO2NkZv1jmT7/k
JpkMYeCTwfthfThmB19+XEMAxojn3ARy5tfzxVRLnC5yjMhj+mPegYSzHvPJvAS5
xrjo4DOklzCpUi4OS6cEfmBBhmYX0enh6HEtzmoTJZ9cL+HAN4VecmvbKJvugMgq
E6stRTNaMFGbg+bk0tx5+UhbsqQWGwfmoitJ/+8F6Qp3asthzxO/7qT/pPR65hJe
UajzHyKhw79x/1XPwASF+p160GtZFALrYJjcLMawIj7siV6vJ2HlnFcmLInM0/Ot
vKgvJGImqtjRIlDAFjBchG366jegC+YUoIOpF28IxN9U+5p0sPSREZ3pz1NetBao
7oC69attHlxZsICmBse1RO5Opf/5R5DUyV9I7WyNxNTuI/zfgRoV+7QklzfptqzB
YcbBZnqHvtea5AUQEckqN+5kGEBhrYy8CIkayA0mautTVrxcxSPqoguI7aAYeT6S
lTnpnmdjBzYjdHLExORRmFtsyHyosIrr2/vUOL8OKvR8yS5USId4yZ6/ITF5tYHT
PLB/Tf7U3/kDCKYZj2daiD36p6JeaQ2kaAgWRtjYDsOlLeHdB/xcp3feLNZ+w/Nl
2Zog1cHfxhhZC3LH/kthCvsXjghObf2WujRmai4ixFxBgpZwDPLDAA0RCH4nYyUq
0SdV1Sdz+fVwSRchtU6BScBoXs0xN5T0O1+to+JBDDy/bXC+l25CVn/fT2j0wrHo
r0dhInMGT0HsHFXtWFe00OJQyxCMai7gEZA/2FEg8vhMr/QUlNAfyHPNI5ZceapA
+LEGgNNgbkL5TUMMunA4ujpXxb0RZajWp7gtteSu5WvfBEEBNj8veIgP5PSN1QFr
HlPwv4zDVtT3iZDwMr+12bGVxUW+8Cbqy61bRpD0sVrQwUrWVT+0EQwYLHxfECDX
cPQi4PSors20FggwfytaasocGobBkQZl+aei9RpMXBJ0HJ4okjLKcqmf5qD1z8qm
gAWSGheEGcL03zEpJPZ1NHX49ieHvU/zg+uKeXcBxklyzAitOypX+5A3XatsmBvh
4KSiSTMScwVPyLWyDQpDfsDuImTX69P6ZmlPh1znDzlGU/GHuYGU95ru4F7OvS+q
g15qYXddwKNJXACfG6KGRNRakWVKKQm84pepbGEy2adgm2V6ujPdudad1YqHQ6my
qkuOx0pxZe9L1Ji76F96UBHYwazB9Mxwi211Z0c3FGtYPRD+hiRHvlbAgFaiW3NW
MfH6nOvORyxL6z/VN0AZoKVllLuD7r5oQt3KmhRZFBR7SOZBju2R0H3ZvLpf06C6
N2j668wBdmB5IkXZXzrGFG7zSZ1qzHICOLl/oenpJ3jvT8fZX5W11EpTLXJTw7UT
i8zpRIRZOGUB1bgXIWukheUC8Esg6ZPQl1e224GCbC2bFlvbAkSySkpDApYcTNHP
e4rFIMfcuRD0gigOLbhUlDFK6L0yL6EXkTyCdsR8CWSNr8qMZRGsNz4kMnAtDEQQ
YgwQSTRVUC2OwvGBhPwt0rljf6X6jSMVwSJ2BvQ+qDLVxRb3ajofRCute1l4yARQ
f+sHgrduPESTKEBqDQV0hZdkJOgBYvSRfu3QSZQd5Ht9IMNGxc4rgSoMXSQvWc5x
WWw354/lrpOaOYS0c39Y893tyAjOCTpx3AKzOcTybjAnwYWjPx9P9sRnGWkdzq3f
wo51hPPF/NJqnxePZlWWtffmY2YIS7CmfAeGsZCWJFdXQvtxHbawN0gKqaMAS81I
99BZk1UbvazL8EAYI61pAv7IV8NJntMIm5FVSIcO2QT91m+mRmC38zaB5a6tQn6v
Tx/HjqF4gkj+7FnUF34XvjwjtHYclCuEpmadxuZf9IC4Se+6Rkctx62ty59revIr
7nd0j3Hki61OPt/JIKq++325wqxQaxz+tdLk8Dt3dteM5JFrUlMeKty6MWEyNn2H
PL1TaSqqedLjImPzPY/Tz/s9aVQWT15mLgb9mYhf8E1yPSZIMrD70YzGKNdRg4r1
OtGj5rrEX5TskpogL4/6gTT5LygXm6LEVE8Ol7SSVoz5fOg0v+JiG/Jsq5uCQM58
4Z7THxai9Sd04dCpu3JUItJi1SqXNVpV9qXDzANg1ATdMBh1g0eBYUAafK/w33m3
kT/fLqin8gmj2tqKU4RCGQncfbyTQcn2YJZFTzyW1ObyycuOHij6WR6vmilWa24Y
cKt/R418nyPHaTU3uepxVDnimCMesCZS27XHTwzXhB/7CM5sa97cpKJSf5v4mUMv
5rxpKBim+UQ/PbWpKyTOKLAiL3HYjMkp6MdYG0bX/GgAbJWID+EIVcfmRieCJzNS
KI04py2xqZ1q1VXGW8jGxTySWXdYmgvAVQVIEWpp/RusuB0QiS7xXDNtqSIAy+pR
IYX2dS3/BmDgHKZEpUiQ4oAGRwyKVklAia0D1yDIHJWisi2r+bTp7vLtAooIAVYK
eWeSmuZMk7H4w5Fcd7pOo3zeTqHtsZRTPjLut56GHAgnQ1nxskQNmU+PnXu6q87Z
IYkZ12w3WQ3z/9IuuYqtl79+QxjCv93Lp471IBdmr8raado/0u/vaBTfTJeV0zX5
Hr+9w2VnDYIHmSTMhhaHqfdPtBFRTp+w/a3gNFKwUTrjMDaY4lQjFn3tf6gYC+th
Vm217GXevL00V+s6EvaZ7tp+k3Cwn3fK/lfP/9dkZwkn0bPEV/aKbyB7OO5G31Qq
I4Gt+HVRcdXBq89Asdse7M2cAr04nY9LsEDoAD0r5xBRoCbLZBVmh/2zB/Qn2gCS
54xyyc/9qKWsbcCXObfwtYZVjDA71VRYbvzV5yls78VKPKCBP7N2dXHY/FQKBelU
KRoF4Tk44eFV3hBgIIvXG/iUOvrVjxoesgo1wZ8Cq/zjN3/8D41g0Nzvn1fzylQE
tl9L3JhR60zCk9+tQuhZEQesCXo5pwcaNg3jT78Otyb4jgaaK2UjgMNtTh7s6wQg
tRvQODxuKBvNXGJNGv3P3CLOYutjXNxTicsBwklr6oToERxktl2rK30BWzyM88qB
UZ4HiU3UYq+pzUjQtqdayMrFJYtWTGhmcuK4ncV+eUAhFrU/cFZxL5f4WrvVJAe0
TSdiNViDK4jr1xRwU4VNyWIcMNIa06MvE8/2pm97CC4xpXkZ8J9Laungf0lR5jea
9RNYzEUZigcAtykX5CvRaMDCV35YStX+2YXFRAOYLOZvc5FetLfuFXJSOTiUXC95
OcYZR7erFvguibL9Zadbd5j1HaapYAF9XB5pqbmQZrmcdtavfY6l6QumB5VHkn9n
lGQnMkcMls82s5Hwu96NchHqmSxN8tv/vmL6/E7/KOqDmKisU+YY4CnvjoUFzxuk
7G3MejbygrzRK8xRwmhQIW8rZFqofPB44uJgw7r3CEucgqhJS12pl5hQhSxDwRlA
fRH7FxMd3Ls7sVzZUCmU3Bt1ed+fSh9oQl2fLiY7ngqXRMwJMtrzMK27W/B8cN7c
z89n7U5pti3utLIj+vSoheoIGPo1CMOqHz0XKrG9M96qAi2pcFnqVjlqMlBabR3d
QV01k31Q59R+f/n//zwSjporoLhsyqtUBTG87snLN0o/q5Qj8hMQlkoGFnFcpPw3
gfFkQqui63e2dCL3o9h94lJp+nMIAyvKaFssKwffcRpKQ09/7mPCiyCUZ+FJjwfu
osG15tmwnFxv7rLYkVex0a1Ta4RdmUJDwcLQoDTa4UUCVdufnk4bOweLiD9qLGQL
jPPs3jrON9/JV5dqBCt2qKt1JBKRgJF6ksrIfubuACWAV7Rz3XPe5sGTZ/mgMjOo
aq693roU4CbYeprUUgMJXukFfoRwRTzOUYq5GZZsG1vr1O2Jg2e2sUPHJ63AOSs6
T88DMOwZVY+SIBOcEcLAY26BvvfU/Vw4Rh9JUhva5ftEzjSWst65/RnAKQVA/jBK
Y292IIY33oiaGCTWm1BUph5tQGzUswrX+lTvScmCcqL0/lhN/Y9XI49UsJ6yU5BF
yDNlR4+ZHh+xd+PkGhhU+gXh9oxUfuhyPcu7Dl3jLCLOuQsQr6iXjw+pYXFTFK1i
vi2SH4sh4Pf49Fk8Xa7i3ig/pyixDMfzYPgyJ5wYiCM/2V9pz5h6581+uS8cUpzd
tOj0L4/sGp4LsaDrQnzZ2jgeOJ8HKPGSEOL/7uSmIor7vQU9PJV+9kSphMk3dkd6
neiH0WOZF+TyHXTiS0at6iCOXfBIR9OyuLYSikraNjoszQvJcNL2TKNchJhNsipb
8WvYhAq8jpNpxPS16VKi49vx7pnWN4XZgAJX7B6gHQh7Wh0v5s7f56nSg5c3kaxv
caaJVhBPz1R6vCpl9MaPcxZWFEJD+dkBED3X8yCsMkc5jeyWZ92WxXxlZyrZ16pl
kxpJQ1z2Z0scEz4FzmrgJo0lYOFbqlwwbTjLSZaOd5VyWZWSmLBtTrGmkEB64zq+
7/FsQ30RxVL4PdsPZCFh9MTTckoe3Z0WWUazaLTP2IqHXePlHX4PYgSWgm89kPds
CZslaJy+pOfAxLKY/Sh2639UBa/sZ1h1nLZs4R0mZlO+Wte29x9iP2ra2PYkJklM
6GMmCT2lzDhXHAlorFSv6nt58RmoAwQLL3YKaV8O2gWV65pe9ykH+VEYPGWX0vIt
c/GHKXj/1ybGuL/35Ag9BRLb1fpkGIa4cGE6zUVFO+jmlbDnHgRVE6I+35UR8HEL
rDeulU2r3xF+4LEkD6dgyabHy5+KxlWYM8j7N7qfd/qNYyOANjbACooJHOdx3T9Z
fPXfuWMAXosMbYgQfQSz3AhTKj+dmeTtoaaqEzClGckYyLuOk5GDA2xH3cQD4PPF
ObXJT+2OeVwL2oT960melHlARh5q7VC8jbJ6jvuCADRNE+fhqmdZV8M8dYeXP49Q
5aT0NLNsdyiXRIBFzZa6+/IKPvrzlgenN18f6Qew1hhj7CdHTSPfNBbEGsC6xGxy
rK9a1dNwFtAi0swITCWYzo0h7+WZNT1u6jv3GGkW8wmm+x/ekiGGKweFp5xMzY33
2N4Q4OEewsLk7/n4fyABuJKa6aw/xM6Fl/D8M+TTRHnqEwIjr6Kjg4qL7f2koWaM
wdh35rbV8XECdAjJymvV76tGMZgbOV81Q68TsdK8U8CTs5B3ldFE948DwUzKOJBm
h3Lf7tXPpc1Ex8bfQ7z8FVEgclEloGdWho/fx2plu2oBrXCZY1q3se3B2oUieXwp
zbaQZQqHeMlyxJoiO+xuABOQlYduuL6nxDkTjr1q1/xKHUQVVrqVogVQ9TQFTnb+
8wTEnBxVjMxf6fzgaHIhhHvspNKCGm9ndqjdbOJdq+9OQkCScjcu8ZVi/tFj3mZ8
giGh0DfxW/ETE2DPn4hTd76oJa8/WRECE6el7mljo7moYMfeIgqggCFSLgolbeGj
rUBuYaTZR5K71gUTydpgTv8iQPadMKW82LLhElTu7gJPP2f4Bp4jrUlT2waBTvbQ
oPK9tcjUmKhLUOPYt5fvmXDlrLELFDLmpTHaDoRmnanvPlNIeSLAlK0m//iXnQvH
0E51zKifrE7UzuJ0LaPg4SoNm7G+W2keMU0AH8UIwkHpZRYxD/BOdGot89s0+BH7
CEHvT4EcYFTmwTRVqN1jAL+/69qEHMHAk2XjLHtNpdKYD69ipwCGys0XV3AOiEa/
fWubDNzTLR6TR4NFckUkCFGzcwPudV5a6AggpTfL+j6NoS5+4z0bPWzIX5+eOtNS
95YiYJp4xUH5fLaggOOtiiKldyekhqjJvP4SO+3XUkBJUz2aLYfPcH/sBj8qN364
FbSrDjrak/ynFLGAT3ZVh7knDV7wBpSi7SxJzb3+X7m0wgOy36ecmpdiKrn3DEF3
jpuE0Mk1PJRAMaR7i7TeusThMnd/rN8TojgVZT6ZsVZ+kUF3iWPRAX+K+HyWLZ+f
JDBzFHfA0B7es3BBY0M3FTmLZBdv5wcKWsBx94sXQoFfSSv2zfIeBJHJg6EstfJQ
EKtK3HQCeu2gz4a51cfuK8kA4gfXNrul8vBVDStlttxnmhvOv4qkXgoptS0SsD3/
IyCbUhXoTBpQN5BZoyNPFyiNqyLgDSyL5LXNv3FwfYhMurlJ8T/3koRXWAWCndh+
q3XpSqbQPOc1PoZ7oPIplA9/csrO4urUMMLXG5tGWnl+a/pP9BV6yq3TPefHsrO3
MxHXFbudsLztoRPqotsKUfvBo7N4xeEZD6dssoZ9UwVs4BcIMPg0kQ4FqWlN3vV8
au6yEo8VpTRZQD6t+s2LZRAM6LYYepy4bdw/WLSf/rHv2KNhINjIBuYJkuDFtSvD
ScJ5OO9J/rtSxY0FMJJghjce1g1VsmTN903VqmXfjpTFV1WhCtf0IQvYOo9Led9S
PCuaEvlvtv0VAgfMNiDmdmtEtQetX+NUR+b1sfrlkFQ4pdz8v+CZKVKdPtwyg6X5
lH5iK500EXHGkdwEQQ15O9IIPl2M81i0F94KsswayTOaHzPxl9cFdioTcEd3MoAo
eI9hMGBJUDrwMhCwedDDIvtsvjAEfyvAD9w0OG33A2ynepv44zPSQyIsSSQ6Y0dw
55L1ym3X8Ty/GQHEWlT+UqDAPISDLwqgA39PkNLhp7owp3HJqa1U+2p7btiMe/u4
UlyI0dVC+9Y6wCHW3m7R6FRpsR7BoqRSN7xXV42gs/qZoA2zD8PkFmQnAmCwU7YN
zq8ULGB1ULkzSvRGDbOqeRZ/Ijuu+0Zqbb35dD2fpEjMfYxHKoLQStIhgD4gtKHU
TblIOO20miAAgsUK68q7QSJhwyuIQb+pYfOwV3Tg5kc8YImVQWsuT2LHGc3DHgE9
wJAdxnVEnrhnu1W/R7/e0GuMLiBQEPaDp1Q5o9juv7O3icnzp1ktwDWCjYdmoOOq
fywThQ6YnBBmvYnNWjf7l1y91ErkG3kwifcjgUhQ7BdLoPINe5J/lKFKFCaJ1AJd
J1TTdlu5bPXDXkxqnk5TmD4wrA4qS1CUQH6WaMaREGjTXcL97DSU9sC1PAFXSufv
SXSilO0b4v2tkNa+6pA2bo7hbqXO6dc6wBKNNBYSV/IlgyVVHJdgzzB6O8Z1mQDM
M4rP22KfceJ1CUh2CYNuaKNv3JMwDUEXwCX/8KuGhY+QaLi6Niv7mhTHYi83MnKS
pbxQUWrjE/CUwpqOd33d1jffKouKK5SxH6CkO7uTUDb6pwxVcT8M40EFtV1bDG1N
i9ZG/2+S88Xd8lLkEhJp9qjgq4Rt/J11MZy5YmdVvtCT3a54i5ErIC4sgf6wpbBQ
jJj+sp8zPB5bFWUNXi+PqWjlMxdUSZWLPE1FOPHZUnTmB6AOXt87B1kx2YmHFpcO
sWKpUUCle097gLd+LFpHWqpXXknTuLHr3itxBH9v2xosc0+z48ZkC5nSgWtPvbWS
TetmmxkroYij7ycAj4I+ZhY4gOcsgpvTjNp8wluNb4CfKmTsYxHWx4yeI3Mhbmcl
3vBfXhrdN6jTtleG5FFUB7QoEk3nI645b1S2tVP4/cub37ms1F45ziOIx3mjSmze
ryezfvnrBEdjP4049uPTU7BkTCQUo26RYIkLpyyOleHOcAFbYdz4xMFBk2JbWcFL
axLBWWmaNc0Xdmsc1O8NsCpuopVtx/0bufmi4t43Gk9fhNTLts+mSSix36jv57hn
kpmXq1BemX9nOFnRgmNYgSgpkCSW84jeRzH5driiXr+WvVWk/vPPPaVEYravYwj5
NwGvDlax8S2r5yYL8/dwwWKNor6VsEQwqHqW/ZqkGGrqpmHaBbHgFt0j/glASQbf
g9ZecNyvsEpE7NkFRBEPlEYyStE21qlUm63asJdKhEZ3ZIqVy1tt/6IPRsH4Jx87
pTK1SdqMutTTQmYguxo+0sL2TgDnoU/grl6F4zkqkZ4MMIaGnJtNBsZuvZe7MeSd
TJtGyh8CxIB0XBMJ0FTICQpahHkANJk/3c4uGsZ5eOP/a+GnkQCv9uKgwEu0QEKH
Lfh8X66GTRyz7w3LINNzjAai3CIxEpXawXVrxF+sLP+xpy0Aze034Gnyutaom4GY
l4/j/y9/MSqoDLKzS8bgQlj8+mdDa8SyuZHT2yG1Oe1kJ5bWx5vD161hKteiz5d9
zrbWvtGKxeUK9zS7pK3J1WRuSlOfXK8/e4QE5gX2YZMCkaWB5FjsaC+WbOD7NAiz
/N0+Gn+bJ8949Qk7pNvh7zMr+in9tu7km5Lo1UzhbDHQ0GlqHVuFTHEqbw8fEeMJ
DW8EY4YFDiCZKVHX5Ge0VSm3ndHdHDLY2TWY8+vokMCxq7/yR0miO6YeZdMepnbW
ETgb+SnPt6Pc0bZnKJFzMjc8Zoz3MgA3eVA+iDuOOHfnRY0l4HUhb+MjiBhQQfYQ
FJRuoLNmnrmk7Cun0g9B6Ofna9IoB9z5iZv3iOrFPd/mueMcOkStoZp2BBtawm/E
KmLNt7dvmwvk9D1lMEVNiZsXjzy+eRjy+Qugbr1/xjhUhaF3jip1Pst50k8EUIFd
HDBhI6Cmh4MsikEb0O9X8aU6aB6yy4CfvWJmjRZ/BC1upze/+RoOrdE6bve0dYc/
sjskld6TFvnrtfyuJy/kqrElRvo2i+WaAo2+abFBJYb1CxuDHjRpMs9Ae3OfHi5U
xDdR2QfDBCX/4md4qWEyZEwMpTNafY9YGz3lgyqS2FKhGrZ6FdYvZkxx61mkKeG4
GUNoMEKRCjT0qX251p6v+kTX47JIZqq22l7LnAC8hzXfy5r7URSpqVHoNYFzZH4b
hHSHujJ1nACSY20s9fYcTg8yOvaIXFUgSIwnZmty23oTa/TfZISlqmffnO6N14Df
GRQnBqSWFwvz1n9IGxeZwx2dXm7+4cb3A/XIsAlV1ldNU7SsILk4Bv5Q9Kg8PRNB
MrAgzxNP2yPbEh4Pto+OAwWH2g+g3YVEfmozdjAJFRRP4A+q6m9b4iJHqBJOEzO4
fNxQaN2IhXAsA5V9a15xzYRLoGPIrIKGzk+XaWrKuY39RHky2Bj4JfafLTCh+PVY
EtjIpuNGJv13aFGthV/7K9EfgD1TjiRhRpoTofzgQxZndA5GsQeAKjtn4V25hge1
KSuzu8EwRRZ2MbkF3A8Y278nPDBwN+dtKghIvU7Wn1Wv8s5EvssQEnKaYZLYTa3k
NlbT17bD3P/t+nDS47bpcNxQ2ApFc2Lr4KXYLlWLrrjuAgpCWs54Vkv1H6Ld87ID
9qsD7FUtQxBt0y0cP/XFPOB5VDChArD51rVz/hDLRc7RVipIhNaCf59VGO3+f0wI
lnKhSZgITPd2lKjYhOgyJQpdFx3YCht5qW3O6s8GA2VYaDnneD/MiZ0qGOGZvFeT
rReCLl9pbRPfqOHfiuK/XNFLyrdQ980EKRqzm+uMRYnYT5jmlqeUs/ERUToRisBf
2hKi9f4e1Bgd67t/Ck41RoYqhVrVQBQ82FHw/u1X0zGnEKsDy5pvEzmZ9d4m5JwB
tq/eraFPVh+xTNUIomS723tgzjL3le04N+sHbOs42UrEulsLYZEodkyxBq/6tOSd
HScnjm7gxUTBJ//dcSMSpjTX9wPlsZER1ojlVQlvxPldV/15SBgRb9fgW2AACK3T
b6SrofkYlLsmMDTe78W/yZ97OSYxe6DUU/V/obcxfJpd+9KJ0V3zqw4BSBNizAiN
e5qaj5bBRtWkEiHoKiE/+7g0Wt5tnVxkEQFh4ZMWrPg9TX1+j69pBJvTDnEqqcLR
pQCba3FuXly0i4VNCLra9xC+R9FDsGJXbHm3SXxjDoVikmFsWjZCzXfNQLi4t5Ps
8LhRrPIEH1E15voVstBPNC1wvxKvxZx2kMnYXSzDRDgs1S8j2RxIhgRJNeeV6Mzg
T7Ixb2y7z6qk8fKXo2c1QBahJJpZ0iAYij4+QKz3skyyk0TYT9nEWUi4LfU3xgMr
Dd52HNWlednVwvKc8vQbRBajO2rVsLQXErVECfYYfRKqWYdn8DP01HfTU5exbI9t
NbhUBGz4mXR1mfRX/C5/XUDHAnTdOOdHE71UO6Kry8kOEVlx/INuK+C3bP689O/k
oTq4o2tZ5w7AjSUXNKYLQqrxHpaoQdBrbVswLsUbMYa0iMFlQ+xFRH2VnylPB52w
wDuejLsXbLef70/mUzD6XBm8anYJTXK4KgQC5a0I0CSCNOFAqcQqSZ+fWj+q1/j3
jJoDsSZLBnt1kpJ/CzpkzjzgyfGWs7PsAo0ElTH0J+i/taNHXpj3zhPNzD/pPoLG
U2Fie++011lf1xuUUB0IwY0W7cBxkRxEzd8KtBzk3YMVOCsnUyw3EEx+TGxphMCY
b7zTYAfbsbpEelwB26FWAx9iWphPKIZOgd/nlN1DOZIYVQHRnX3xEkoz9QPieqFE
YB5Je0KWyIBC3BunBdDjqZD77F+IxatU1H2P4UtCM3bva3ALk7mRp25tvA/6g/N8
0DghYDBOzce1dd3EWAI53SR/lrVqvfF4XaV8De4JTOFlg2cNIBaFucZLBbOS/xMw
fq4id0TizxY48BtcjLqpKtcFMD3WZw3vn07G16Mol1IDVaPgIohbguokKpC/tamA
EwhbkqoalJTtce5jnvtmKtHOED42TcMnCUlGslh3pW6QFfdrHz17pvRuUFahSMcZ
G4n5v3IOPH+kB8m1TklPsGz2Gf0hMtDFBJc3ec6UlEy2QXoM+irx+UOvM9jz8nNI
uy6NuuQmlSadUt3Ww+DsE1eSRTPU2LJXqH8Dj8BYrdtoY1bY/puVqSS1/lw14Ysy
yMEEaOlcKWrBeR1bMSYkBLUfoG2evvYPgKzJYyYsvh+4Do38/M6WZRypMMIJayBY
VsoIZBDc8ptcUENnTdUGvLkBeSgG1fBX8vgKAGhHb6Myb6TDemmg9YBUMrugPzIL
TjGljT9EfTl05TjQUFU1Pen6JzgWN5Jy6RmuueBNEEM0lOhIqwg+y15chMwaXaBu
glohwEnCyv738CvWp3esPV6BGA5pwSByN6uBEBfUWJ40Cws3XkjobUJqX9lGZG3v
4P3a9jm5XL1+6GF8V82Erj7VhwVSedbQS4o0dMyKlC/4FXc3cOqa8LYsr0rEswas
0fZRCzkQGPEWDNrUQbzjIaZCbyMlIJZI8jZiObNGWR/yCwVGipg3KMx4+PJ2EaWT
QztGiasCAoU7E/hoNjvPga7Jrxoqutj9Pku8yRBSfwtnMSRS0EGptMuyGmAxRo1Q
BxD0MWGqTpqn0Vdh0FCfYZ/6Sb5wCAVeZGfGlHG28FfZWCruNJY3QyHrp5SqTrs3
bkbMicadd8K+OqxcdIm2gKML3PGaP8RYYD7hPFRdtYZJQAuscyJIsld5izIgTnUo
FeKn1xOe8id4B5Ouk/ATwyiC+6O80v4sHWLrJ/L/UJD50rGaO/Ig/NIoBMNSRH7/
g5COsjCGrA+S1IGecHoYCRnW2dAr0uHwZDm9sd5XcjyP+kcaZe3YzF48HmLQ4tw8
VaEcWHkZDJFf+kLUU+HkoGEgvReb/2wZ2GZUD0PpN5zlc55TRZHaJV4bmHWZJxHC
2FdDIRvEYNbsub11CrlGj+HojSmdPG/4/dtVtiQ6jHKuVhBVFTkEyNW0ePkUmZcG
bQ2GH8i+Gf9aN+AIQEXtVoym8AySYRO3EAOHzUBC6k7vDZYF3BWi+z5ROIjnbMnJ
EzLW1Jm2xdeU3QsZyodhNurW8BbsNNUP/7GdJOMOnAAnKXdMpEf03At9WPqu2RfY
XMnm4wLFXt+hGELIztC4RyCZSxtA8Uja8ReU3LPpdrkicP/bLjzjLIifQifYIOPo
rlIfcaPi1KfANrSXwZ5ApG9kFijqe9hl/pBlWsk9a+6e5SKnLHFR5z/rIbPzY1/G
aAfm6tZAL1XHn19xyRNSEthMbT8+XtU/wbkyrlYnWv8X1aflxLhVOFe+iQyfljLG
N8zDEmZXO56hzGfrMdY2Q9yf5Z8zytVO1ka+3kXfSqWjBvw/MBZxmAgkqWHfPjRH
LXwPRD+YQdR9gLTRjlZ7Q+LO/tdTrA3N5+juirO/54ADM4mtP7aK5IN2pfIVdnrX
2dHFaNSsnlpm+3Sc7rR+AYBv3Xh2THQK6E7l1Fi45Oer4uOJ7wTk/lhcdke8Bwsu
1JG3o6HL58bLhXGgsj9KZIVXLtk5fs06cZ+fbygpbhe63H4Djy6/582u/BI1mOIF
YmxHpVTCnWqibX/kdqu9eMXuHOZeSvzLniUPoqQkSI4ABMvwxDS1QiOMbDwsWcfa
avAStiUrsCcVhyuNmlST2cGKGT+xekLktWSirGx3hU/NZSK6tebQwyqraMBbp2Xi
jxt7+21IvlXIQUsRTSMLh5lKVCf0GeaGozAZJacxc7JqXKsZRMymWI/RpttFk85y
Kfk2ARABUwdHgLNDseeUES8Nvq8to/p05U7ByzssrzfGC9UMjGhVcZXo8Ds7hBBd
1nrR/GUkAQr+3kZWDBmQvtuTajyjYQdsQnPrVq+j/3LKEOUnM6XZXvwGhQPHGzMh
WYDgLy6xWPk6XTZYYSSlwe/QHZsLFofr9IawvYZJ3MurbCSGINKJqAtoPbwVHPrD
e/QJpZdlyW72qvo8GMDtSIvu+Bimj/JZQybj13QxxUgwr9O2tLyCAiHDCIPHi0pi
hyu+Ndo2QH7rZwf0pCD/yHPfk0UZS0dsqRecyZRnQorIbCX5hYodATQbia2SRqne
iVSwvdv/rJOnH+JZvVgWFNAzorz2WH293DJPulk3dc0bLwCH7FhDka+fmgSN7VDi
oDX64PmDkOh2h8SZtwyGn8bAaLDt/bDfKT9suBc33JX/fltn8kxzTY2yUCihCUjL
G7BOu7D7+lAeppSRpzoo52ZzRHeCGZrZeZpBzZ1W838QxAlgJ8EerYgcmZWeUAzD
crE44atdpN9Gjwq6YS11ZJ/sz7V0xfEsNxTXHkFyPwgfseuuHjHw934nedtqxZou
CX4E88ncCl/bRUPHy5+cL96AD00Rvu43lqsFHHr+ioKymsOUBu45joICfYKMjxX6
FitYJAxQdFN6uB+ufvGxSyhK0tnV4KpurCRBeuFKw4g0wXEZUAILbQCkIM85w57I
rx8u1cBuT1oIDc5xfq2BTW4Q7OFQm6Z2eQn4nzhF6iBACk+DMwQdiwhPSnVb4KAw
al1hPaq6yfH969tmat0NQ9AW0QlQEvr3nQqOpRD5m0tQItqgNMhaT0Y6toD9KPEw
d8qoY2dQTH24GKZQdVFHK2w/+SF2TiniAwiX0G+XTNULynLohsc+Xv7zwJoBLz5t
OMNRK+v/ReIqPGcF35rtRHgpxH4V2c43G5K9n/pSZ94EEhP10BCiDqNDv07Pnf6N
PDiGR2GALkqwj1Bk6sQ26Eel/IHKj05i4/uqHOlKRwH+QVC2p2RML545plGDjnsi
yIKGiXFU/Qlvn/WFRskjcQI45hzUT1xfaYbMv9D/gkEFB4p7HvrKsbf4TbNhz2BL
2O8GlMRTNAAaPJmon/YqFR4fEXXLvz6Y3L72FydrlP1WXiwroPHGv1vCve0cQXD8
lilsv8dICQlalFx+0XH4u3O6SB5JvDJcDoZLQYttfM3QC+GssbKGqYL+OAmjnX0f
/7zBdkNOKrt1vQgkcNI9U+BWsuhNgsxdplawPxjhGmQ4BT+dmF1VSDN4v+wx3SYj
jz0pmHh2Yn8+r5kbEimIIyK6P1HcreLzU9MSNzrpbshdv4gZIQvwp3V2vNL2Jl+H
6mCQRnJaT0eFeyT8AYGwsHxkYGnxEUWM6z7bFvZ5Nnim5GAZ3LndZFDoSWbAcvGc
dkPUT59VBGbUc6J7owVxl+lw3cVN7jajEjSgaNhczBSIfbdSau/3aOCHqzi+xDJ3
wHbCu3qiHPs5R0q4LqbFX1IYr1crEoU3tDSIKLH6Ght/RweLdHFX1lhCZUHKTrS1
t7vVPKxehgGXOBbH9+2rycoD/wHGT69VtEda15Q9DkfE68P4LpCBMYsmu6gaF7Jw
u3aoaSOtYsWQkb5M8X5YWt7q1qqa+zev6AzeI/MXDU3l+XKeg1/CLuKgGWfNndxL
S82t6rUHqUDnkP7tNZju5Z/rYdKI0xyL+LtQ+aRUm+y59OBG0Jp5lfI3AyLrfVwB
0wml1hwIjei3lV4pGSoMBFAA30Deyco/qjBJs2p5VjZ26Z8AefC5uT5jYNR+1uwz
k282eBWKt3USpfcg0PfTgXhNMKD0hYLheDrHhWt3wUb1GXd5OkW57d9JbkTbDYaQ
PkZi9MMuohzq09hcMp+wIhXFNFH1dyNghtpDrU4ULPEDAFhils7huKNl73zcsf5B
YXsZPkSMJs5K4uZ400R0EZwFbxz1q2yuIMv/4quxm0ylUPSWi8TDpzjwF63M7/BG
tQGRNnZfb69xL1Ep20cqVN+hFFkipdnyJs1vhiRFFIkFnzCib+ZNaoBInJ3Lz8dF
64sh8ZP7zAqR1DwC9NUxyuvUCjnTZI7bYb5d11oWbPHsSd0HeyB4WDXAAcBYLcto
SJpUAJB5GKbEYB6KUJgpSsBSLm2Pp6jNOJ9vw5+KPTVVpxOj6cf124mePXM6jTjR
S4lUu4NsWW8P4LOJF+s1kKOrrwTNRvNRmn/YiL1KBHoxOIcTkm/WTZwTdM53RmqK
ym1CpkC4UmOsx799YndtLeJTghjqRSpJlRFg7swwV27VydjcIPMuE2t2+d4lRW7W
EQTsQxjV0vSL2igibRHDSeWwy6zoP+FD24v4+6sqx0W/rLKE1lm0vcgIsoJl8ydj
whgsK95l5Sp7VWXLOCp5Dkgabi7W938PV3a4N79/2sL9aGvCqJVN5g6fdSfe1qkJ
PAx3hDbJjSO4jOI5bz8dRcX3yzyiUNW1ig/WMQN7dd4d6MSwM8Ji/LrjWoQlDLgz
k8VBUG8bUOSVfFp4JPfQs2aPOzBDWUztx0QTZ5vNhjI2jYCFYnCcKsgdiX14dMu9
lvd7O4WamR3HMhczHp0V2QCEwxm6MSE81CRo2wqY9hNRsib53OH/sQikjDXrtjAN
OGqro+MI21eztrP7XETFbKy7Nn8KoGIaxlWZouwFsvR/HfMudiH+TIwAhd+T0wpV
q775/ZA7jy4JLHr00EPIIts1CTaCvBd9JqtCYbaCDZS86GbW4S1831NOsu7da23r
oiPZzz/zjiTdAVaFredE2S5zLp98eByyLHjvDeflEpOACiDboL5NaK7WVaiAD7cF
eGFEPvr9vS9wUbtCmnDY0LSzH5IaD0BS0s1+Wu6RKipz5b1LM7mnsp2hRGLTDJBA
BF0joCFTxy09YyXl41Ntml2N1pBEeMLM1EfJdDv+pY8s/ofyTwLlSJRl/Rr+lzLx
WSg2huDtXA0vnkIRqnVw5GnH9CkxNHLA+2cYvpVCxMJOQXvhkwLG6+qBi54EYKaN
Mmy29uuv+6YnAb1l7KRA6k8++EyIwzqh34DBkpLAC72XElZnVH5jCSKAef0Gm9ZW
YEl0iK0fSHt/nOTYkqu6bK9SMR1vqyHTUeLECP+SijsP6MkLIlKuHjz5H9SDVdh0
fNhSuWujDhedUImtoBdKr70fsdZb/vfZ/l/Dms7JWkBEY9ftGnl9j2py9sy6R3Pb
bxxwfkfEplLPQHMF2ma7h1kRS2sxmp29onqEScI8uvXReklJ4+T4P6xhsyGGgf4m
w9oauaoRPKvMI6d7ivu9A8s8Es9HNTzqCuxXF+XuRpbHyszWbJmePZApcfUgIK56
re4trTlBu9yiy+nbQbdwk+Yp2OjgwQRbXQ2t/MgsTaguTeT1XuD8IL0pq/ICu5Dh
Ne18wM+ULoUrDMEkPh2YtPyb+gaNLQ/3+tg4T+gKBlP1JfF5JiEti2QpCuc9nkuR
p5kx+RP383dObupDxFYT5n9qswZe6u7dFJgZl5w4RDXuNoMhCOhsxyqk6nH7xDlq
3om2D402zwXvlftm/FR1lmoJtBlAkR9qcfKQz7C7XoWOYfEz+uEz4nKNuFv9g0cb
4Q+odcXc1iP8kwt2CETDTIW6ooY4ZHe5CG+5vI3cdGeVFlOqYf++PS7NHC5kY95e
byR4zT0iMZr8PgMuPnBBPklMY7m4djwvXjOJnn/HQ/4B70Oje/exNDH87M2/j9x2
+A+UHjl4CtGwdixAw/ramt3FO5Mr2fyDlnI6rrVQhV0NtBTAtpRFqUTuCCAarfE5
+A+bGzr7Zuli2XaspUHS7pnvoe6ni+kffjj0/Gi6tSauHf4mumscGNBtidxb9M2r
YxYjGozy9lOyPs1WdlevlAOM92ZON4O1t9HM+VvrK+7QdOOTjm8vdtf3b/yB1+b/
6sJSVOeFGT5CF6fLm6bPj0otJv5v2W8BbhikHSXlFFsuANgBI88yA+r2E2ehKpNR
NDwn+DUendjyJ9a4s1Hq7XNFWaptA5Xm4k+5OiL2XWi1pIldsppZ4mx10u65MOx+
oS1jzFsxexI/W2eKbg/lKMXrpy0I+nF7gNBgKMUaTBSfuUJ9Selj9ci1+WGGg5oz
EOyXCi35Dr+Uupi5BTX3RKHzygu+l+1daFXCXyHeexyCijrCX9SshD5/XpkPGa/5
5ZX+/ODvkuMAZd9jKRXB81V7tTJTloNw24mp1h4WodgOUqrazbBKUYGRoKl5UGkN
y50TzGqlXS7vHf1dXuRPQyev94iixMbREGyojP44WJP1s68ggMtLimvdjsDnTiz5
ymB9ml6hXU5KSDmE71O7+c9/6vZ6sSgcLC/Rz0Z4B9PJ9o+QCFh1QlB/LdmgpgsN
+s/8t+OfhANoeIwFbpyXuOYKsVCC0IeT+3FddZj6Fe8EdRWg2wlcpwkS+t1iq4zs
4PIbF2zZgQLlhJrvZ30rW8s5HdjGDUChLrz1idz01IslfzmJcHOBNLxkng29hpOi
QC0l4v4pdE4lscsmyw9+Ifw+il9slLf5s6eGC1/XhimsgJJq9AT0ZN+LVDNamMXT
F0ZPtD3TZ27aKwqkCngZ3kenPMkt3Mri97Jyq3lZXmbrshXRMLtYaYBaGr8ceFAH
nxhCAyzVVQLVB5t1Ofo2tUXXf2GTlQ0INcn0tryOuzdChNo865DyqYsFX5GdUxYy
9gUid4TQaAVTUAb+EczuUqtWW6X8Ico9Ek+5QaZ6B03YoLqJjSIELrB+HKxOa2hj
anCUGeLcQ+19eZtnvBYunbxxoVJpioTPvtAedHae0qvGrWPPFReTNVjWjdcZ1zbO
0p6LXa/ZZ2t2kF1uUGpn3fPVle3tfh3DlABHZpmrTrpVEOKHm4sNZUCk3W8HaVD1
rm8Z7ACC2RrOk7YwxVVyncURmYNUz0mwJGrZL0SHIstyaNx/EVbzqBStuF3+gOlo
iTGAgHLlfWXO/BO+IH9jjSX8a7YXp1mxUJSRl/VJq4SYIBfchzb4IknxF/psrSQE
LlL8Pz2v0obEmSGvrazh5EcDsiWaJK7N7fY8TTmc1m4TzGgd0BnY49S3mhCEUZob
ExOFlZlIbg5gMxK57a1OeMoS/+SbRA1uK6PTQ6PTtlaOvVDJRvQAN9VfltOrUZIB
zEG8sAqqWAeYdAtlcnEAvXsW8rGa0W0rWle2yi50mbBHYIp5HgBLB+aZzltLJ3gg
ZRW9+NtwA1XEGAkWdO2UF1eZobtKoQc4T78uFpTFzYREj+ubBwA6QStf+BV9asWC
9K+e+uk5tE8gM8MDOVev6B6pEp7fRVH/KvUSCP2btM8VwcBk0yNWSNO39HU2QVCW
ShMXGl8Z0+ji5mIKBycgPSgol7+A6095ZiGGOLYTEc0TblrnPjhufSbdy978DNXo
UIjE+KVApmWvILMbK99UbCxaOQ9tMayjCmz6dnSKwFhteiauLQQrlDKkSJJRMeLu
gZHM/jBIViolZ5O0t9AiZ4iWqOI3vA6ryGEj51qNZou4spHPozuOfASO7HvEg2eu
ZqqKN8tifOkcFiFAUW+IQj9v5VNhv3QaWMC98T5L/ff4MimMRjImgx8MglK7qDRk
k0d33HBerAIvdRjm67xuIuCM3u2BlD3gdqw5czDSAWA35Wp2pC1KdWKbAC4LQWE3
oIRMp+aOx37E1q/1CMpOd8cAADLXXgL2acqyiSlkm2fgvyd+gy8wK4lhj3JmF89/
SUKwgWcoMOQ2xlfnSUN6cd6kyoW8XwgWRaHLGIeP2I+hAWvXzUUePIDV7m6h6ZiI
c+J7QjslkBi/s/rfnwI6tNJJce+paklQog57BbRurlkOYXlW2/pdbbVW2TIsL028
LfAaaA4cTjr5ph/53mENkSpcG2xRqjcA8wQ0MtfH4dH5GZB81vWc8MvnjGRK0BpC
bvg4h/mFIhNe/uwG+vCy9fFaquhjtpNiTjknNwaCxvL+owxvo7ZT4G+aF3Zf9VmO
5pawCHxli2sk3B1diVi+OFdzY+bu+jUGEZV+DTSm6U7i43yA/QFGkqJbhqbgAV6j
2HtBApWGwfYVa3S10bbVEPY12YLFc0wpnOy4KWH86gyMs+SxT/3XhcaBnNJ8aN+O
5+vcLUYRTSEe91djVfJk7aBztJZalhvEvVWd7IoUCUTYwur67KvHbpdV2CSlqz3K
qrPaqKkEXvmk3ayobTsglRN4QtyGEpuPYbEnwWg2PZAk3DeSMgkJGYqEAaKkxbIP
QVGQoxxMVSR5ZiEJ1VOl1YQf3UGWVreQYLMFfT+ccWioZwBm2yqglv0Nsrq7XfJJ
NpR9H6peqTlXRLDDwxxQ04l2uIHVbO3ic3ITkP04HIglh0idv4hw0iWlxsMaqUiF
KQ+BM9JpoNO8Gr4jwHiPJGqXIuOYi2t3rLrPZ3MU+Nl1LyD/PvMpYEEsmFXe05+W
ktkPqFpYyTkuE8cZnSO6hwcldAEmTiL9NspopvH3PqBCBo5qlHIJPYUSBVM9VtKz
MuRdcZeOX9ZfcEES9S0SPYCNXyWFw+/nTj+2p38Clfz8PQ3NJpQFftBpFz94XWCo
yyjXfMvKoXBiHYrG09rAwvSPXnQLAG/cgozXj8RVx19oTcZMewrG+SiEwjERxAwp
aRyuWKjhZBDXVXSbiIl1d6JJmKgtGUc3HGj1tE9iugbO8ELK7znWQgd6Zc7CUE8Q
2EzKdYgwl51I34TiG5XxoruaK7nMk9ORYxPlh65tqaWq/a6z8tePzBFwmufoAmLV
Quuz2PF80sA0MkTXlvKLdXEAhDYGvnPOybI43GMyzW3TrwI0vXU9xBnZHgV6gNlC
w67yhmAWIvn6Mso0CSvjfuyI7Guu5xe9p4MLHKPAIAs6i8icW2jRN33Q3JpKAVIL
wQSFc5bdagwOUWt6tOkpTUtbYlf5sudLUurxlNmbiGF00IfagoiHMkFgkhLOYaXe
5P65JoGjA81QPDwkmGLHwrJ8HucamoOIriobzhA8/jBdysmMU5TKgwP5FKB7raL9
H8ZCZawK1JHaF8MB5L0VA86/Z0aw3ZiAvrwFmgs8DnVXOKCllSX/1YoUrz7I+vrZ
w9pWIarrgXrGURf0efx0t+d0id7YD2rdAgL5eunux1WeJj/YUj+BhJBR42yRS5jC
rJ2k779R8TdXGLpPSAMgZEvZiyjBRGY5O/JT3PqE/rheRlszsAcm+cpX85VyM9ns
Ac/lWKL3XAyGPtauDz+wsAipS+dwDtXCuhna6N3V+Pt6emue3MHxu4ZWi0eT2Fea
sF32scMgIlIQf08CPee4qljMhpZOzEYQg/s4k7i5jtFh6Bm4EPb44LSz37r/wexi
CEQgSPGSlcq458VX6BhoJwNHC1ET66KKx/p87HpEmBRhqJDfttLQKD3f8l2tmTqT
CjxSugE1Mx7eG63QshaWmTQg5JXJs4ThkCYiIly7S6boSSLfelTChwmyBvM5SGQo
xu4zpe/f04mIcBgwAJI9hix/qwwiPZu7K8Z6CVD6p68sEOTPTdXoU51PXtD+7UQ1
NUOIy9/3LfXyNjum3gEsV9z2mTD1RdPGMJ4sBfpwV/8TWAbtc+zDBUtnJ4A61pDj
yEpY4B9beRPUSAcwYs9HM9Hacqj6AXRWsXm39JaSMi7kkAQn7dd0M8trgHmpKCpn
/aWEYN7vI/o6ShppcT2slk3F3bNdJOb3E0PEs8fM8evAZpGYGN8mzpmxNNCbTnHK
h76JaUSfZhb45TVoapO2mskbQS83zdfyIIMm4Dj1VxxDHv/kuupQlgJw2f31iXj7
hirlY9tiNPMlCemAhCjXwpoERz/GsMnirJeM8cdnekN6hjpOC88s6FZluV1BhSlR
xrdrZmL01KrhFni3nVHp7uYdkzXYs8Ey16RlgeOKVfa8dkaiWd6BrPmdFsbHaN0e
KSzggOUQbLlufxAb8NOHvrxWdAcT3IuabC7qm3dLaS2Ycid+NaKAqJMTI7OQw1Yw
fPIFSUKm2giL2wKAE+HPGetvlhYx+Jdoft303mSfFjDCpIod31d5Npb1ON4LFydW
N+9xzvdfP1tfBUKXPzWua7QVmyAFIvITLaQe1Cj+EtXFb+pQArxAT2h/2qBKsok6
grXg21P6anIAiAjyP5FzdZN7xZODCO5mL28nLV0Z1pSLXFdmkrNVyNSqj5fPgUgn
vVttmcBTC2KV6ygRdamWLH/I+tyip2O+WGg3ZlLff5n9n/IS3wz43zGvXfZsGuAL
QQzm8x00YWM0W36Rm+KE6YKqIUUfZ5/ACWgo4vxJmVTz+eyxcmKnr6s8oyfii+Og
hjPOhFVuX5S1TOI+XPsDgqwSP8Ig5xUPVMMOEuSCcKzw/X217b2HQjj+PsapK9I/
xoEFTgrMCQezwkig99MdViLpheDKpqseCFgfKuGvKiexzZAp/CE2PEHAX6w8Cvh0
zTIa+PWUhOoaAGXJ3BGNc8JEKGHx1mzDdcIbE8dsaMedw1Ezx9+fRPEd5i3Arn+W
gN8WtdlixKh+hyvsOSourJPqpmYy03TOcp1y95AzhqcMEAMLwi42trNTovLNY++2
IF4AtFiMiNnojKIfltEkSmAD2phWHYqXJCeEseg1c+Z3mFJiID42DOCWbTwY2nRy
NlIRLcmwU1RWbFtzIRZTcEz93Y74I6m9fAzXbMhiWW6ti1oU32sKdgJGzsLtsTsz
Ba7WSyoLaR2pTFLAt4cS4EVf+lmRBmrvjCIEVN5mH1JysoXyhJLC2dTq+az1tezh
n4eb3eBofPMZ5qYolW7d2jh98qOq2FHLjHsps3CpDkx18O1S1yreX1d5gCEHm5x3
L98PR5+DDQSJkp9aLgP6yVer/u8IC8TDHmW7nfKBCqOCrNInGmuqbXq2mcnWpU+a
wARWBFkDXTSIa95t9w7rCQAYJFeV7SXbt/0F/7Gzhzf9ev3cIn+MbqM1gBm1A+6h
Z6lUv0Cn/z+HwJ+2I2Jg6tegRz/44iA8IHq1Nc+jNye4gKyFQv0fzWzbssYIwBsG
xu4sI75vSJeLC6dTYZhZDlb+xNra8NYCH3cQmJ8GnAaHOd8BZ5jPTQ35GJzyPAOe
DybI+HPZdS77JqDZitFOLCHLskMTtIVIRi/C0MIZZmrWy6Tm7tx76TKlNuDeWcnh
NFgWgNUo2npUt2upJuxiCQOBfvAXl+ADryBZAjEFz2pu7ZfvB0ByqZ28NcfDy01G
H8/Tgki/oZkeE6GWJdCIQyqj8N9QJPehmY+1Igo4R3XWQ5JM0DqlIu14Ed7j5/EY
wXX3d/zBu0rDdwLWx0JvNqfibGJWRiwbnlQCRn4U0tqEh7tZAu8gkwHyHqaz9UaQ
6w6EjSEk6EKfqWREjumk0HX4g3Xv3noYuu50n/izEJpAR/WqWX2/BaJCaQZo39WZ
V1GuJ74EUhi4kxG3Bdec7tu0cAKyFDJZ0/c2SHKMF3/7SlKv7qmpuHGZtHIa/lQT
foqwUhuWhrACuWmd1/nALaufM47nz91NekcZYmm2IIlRiF3M9Va5mjIX/u+d3/E/
mEfa/HNVX2BdcYz8nIChPQVD1eJaQCiOM4C3QWhT3KfbGhTLzqWolQLs5sgIoAyK
KgcH2T/hMjF4C66uD7OtOquV2FXk7qJ4lxbE3tOnw8AoIvmjyKr6aK1qvXZEsy5n
3WxRvSom8cZsd8rxxoyJsEOlK/RC0jYCxyypUOmS+4xhX2xnrUKfSJbK+zgXps7N
6QaLqjNnt0fDHSKu1IEoQpXSjj9qgI6G3saLPrh1tQE4/XjGVWF0/UpTBUPYLdlR
kdz4iXmAZljUbDE95g5dOY/J3HAAlF59AUs8375YjGeUiLEJrIvf1o9SmAEwEOy4
Q5/MkHLy83xk7hpkq2rHvD5logmwyBK5P8TftTT5WMf9OE5Qk1SoWkMywDlGL7B3
tFbXkn+R5zb7/oabmfCvvlnWRB8Gx94UhL6sAzsehjekAKo2+VkDNdDgIGmm23AG
VkIFA4oYxEYhESWlHYBxc7rgRVtZbVkaL6Mx0cdn7r4msymBq8jcPid6s0wpELc3
76jt4mAZhGMlwBCt46/v4vhCwNAO+C6UVnfmksc67bLm7yvA41EGRgkxX9zByHFd
IRiBFQukTjAYE+rctc1vq3gidWZ7D8wvR6ZGW75gqbV8i2CqNLWo3/NdwItCGi0J
WLQP5y38y2TV8l5lD5jYAh/2AR9rLf32MKM1g22bKPlNwsBjohtV1vEa8udAmZns
MmWJzlJ+10CE74bTUE6xwTgWdzjAaJYRRmcbAWFd01GRvsV2VxJyWW4yEcmUW+t1
TA80RkKWrU0WchPQHK4cabpAlUthWe25bhCNWJk8raSpkFguPinw44clDWd1BQN0
VbOPCj3x4ht78Nv4MWYIXcZ7CkGrxS61wACeb4uGJiNXBVuK0EufFcZwOr5ET+Co
YtM4BJHiWe0OYGvVs+YjqGxzJU/X/2APhpySkAmfhpgLdVwbegf4ljMXTbAo4FAX
vL6Uza2m0QE7lhfxTnstge6sDLpcQU8y98sxJTg+NxZ8/Cq/+FJKmk70RwAatxqz
eNGSP2KH4SRhR1VNxH5+ROkUc5rvbnlTyXiwZQc5KzqHM/QcwPpUMhmyjyWo5RkL
f4FR+6GcOAwdwRrMNkUG4z7ZAPcXaEcqv1ZKnqJ0HrfRmAHeUD5FT6oYr/6s01kR
ywVfaIw6WATfY+3Tkkzqbd8CUpdJuDo9sp0GMJ7YyX1KJXnGlRP7orjxSMh7n2hX
hlaAcxOIdXHz3sP+LumwKx3rFtb216+mUVWXCNmox49hEm37qGKtmOnfXH6h99HU
d8fKsaEL/c/hl9te+kvt4buDofcY3ohKmyeYOX3dhSmN8I+Jikx4cZhq8hEMikh8
h3wHyC5TvW/842Or24iGBZfJ3QmHRgF1zBkWMeMh4hIeJWNjuhHWd57coWEklPYp
rKmNKw8sl/oXxApwcs6/ZdCaQDgcZ/VUlNp97Ehi3z5cDNt7wgMAbm5f9Oz/akrw
rX7vYSeeRYZhZmsAX+sOU2zL+eE8rWEwjozrZgqcK4tPrc+afONo1rnexn+CfpoW
YNKydJ6hnLmbodWXaMclrj9dsoGna5YfqA9mk6Cim64ndbjDXqvGJtuf1NERkmoH
Pg1KANZMAW3eXo1LfXA1l+FZ4IUW/jItRZvY+BQWxHps1yogqVhRZsUrR4aP47OH
Ji6JBfIyUFfvtUj2IPC3DdREYKh7iVofuZVc07Xu0BAjKq4KD4kVNqT3TIUlgu2J
DZZHWexi2z4juxCSdwqJJTZJsvv05PVcwOPf3Qm2FJbUlbldtKRSTemlsfxSh5pU
GKxrp0q+mUJM87ZyOUI65pWa3AKC9pN7g4GmHS/k2dsQIwsCIXqA5WpNmvzL1I0S
3GKpN5Ac3aJCqRsIk+IMbCAhsrEdwOM/D8W2QdEuGiAX3zo1mU9TD4Lxg/vi5wbk
T3hR7YOZGJZc1rNJvmJjWUSkFw1LlR6ycTHYdXFr2DIf8RFpR3cABbZuftwh+1Ug
eScgJysTbgANy6hlK/DQznHsI5K4xA07Xuw+koMq9g7IpxfeolkYLC+FIY2rDPFi
YOUMXmotmQgg0lKrVewNa9vcWQkh3eXLLiiq+t2zz9yz9foX8+8lgCYjZdh06XU3
2Uc5rf3s6LnceXFI7CcXJmL0yKFrKmRSjz/V7vFkJEEIH8ims54D4FMXGis8ZFbI
eWQFYeBwslnAqWJo2YmTHL2za7tiXjg0XXX4Zha8T6FMhPjrW55T402Td/J2ebEk
o1FDj0ECVsYTqjpZ6QnefT0q7S7+eEMSF4+llcMcMxRnjfb5hS+3Sr2yMijzguUt
ZlaaIz0B2eDskyCPuUO7Jw9lAeff7QBLKNAwOk5cXJvy+hgoJfcg7wNGhzxreB7S
/8cdq8qNs2HzUtJQNbp3pkxKbxGUaSZh0Gd551I5sbJiCSYQYFh1Ef60rdajerN4
jDOjVRrTja5/gBdOqLdBPuD2F4ZYX2d5UC42C8vtGNIMbj1p4kK8KlPBTe548o+H
m4bmIbrpyJKc5+0U4xBe/KcRTtsMs/QsWSuZRa9ooqbXa1csKvOHSzRPlXCWbkCq
nOkQEpbSBCvB9tv0wg0iftKev7ZSv57KmxSrvWolNsRVhjT98qrwCSam6N5VrZ5K
HA1wP40cJ0Zt4ANrkuj3D+kNs+XO9aQsj6Pb08U13vU8Oa+zoGseWi6WRJ7nmMbc
7Enhc7nAtT/hGtI0OGT0lAxHgcv3THLmlVx9MCgEuE+K71HNs2F5Y/EIQgi7IHMm
TkfN6n1vNRohZyJQm3SeVqMUX2hv5T/CF38Vf+AjQCiJVKmfTBaNkBjVeQ97KLkW
uGuqiWypZTNcFqoN+pkjRGv93d/YhwO9ESxtLMLNgXTqqRfn9c6uydOmvjEMpfsM
SNtdNzSlvAa7aOQkPEhqGCuJJ7SSIvw9V/DHN5Aj05UJI1lSWoNiRRcb1v5k5MKd
dXdr1x82X3bKyKB1Pma/v108FXjYA+8//RneJDxUV+KbvrOodz5SNOj6sltZhYzG
aACZFbrVhDwGFzdQIVYVxZcAAkDDBzKeGS+xNa+Ak8BECS30OnZY3DulnaY91HYS
DHMXrmRpmPSZk29dMZW2aUkWvcPWcl/dQKzZWazgOV0/ulsKovlFGgm6QFTsIsmB
06OXrMdVXzhFeWczzlocPszwtx1uRUD3rWLGUVQZbLyC+RGs1n01Hgh14Sdeu7mi
pbsy8P3BnLx5eEZJpDcpxBSCBup+OZtvlLqaQ8MC9iNq6uUYQDjKEVdNZF5Rc7e8
dYvTRWPBtm1r+/HXr6Wi745iWGKCxuxFUnVMVc3dpchBXZyMEN6k7yoJ9+YVLdMK
32XwF+jUBTNwleswpgd2QOu+aWKhFK6k2mbEAJqTcfKGl/AP9SularFZfArYqaWY
diN91lq/WoNhy4KuM4g2r1+OoN9rHal+nfg8s0/eKGer12CdGR54DdgPEDBCBp2+
0OrYk8bHMbsJD7XJKsaAkHAcfFQ6Q/+NsRY3ZPO6ZGS4j1w65DQ4sHEp2kqNrueQ
bmSr6YLlRzqbV5tLvXkaSyhAckxZSbZtwmKB7bn3c1tQA0LoUMso44MhhC1uzEoh
XMWbW8y1e5LPp1jwt+h9S6nndqWkdbTR6x09QCflbepSeK4ipA+y9CdckmOWMhvS
8oVpDHjDiY+7hzbBBdD8fm7lsV/JYx2TvDs6OW+vqicL1n82YAB06f7JujDH8lRG
g0HZiw2vOOUUUztO5eK8WHt//Jhpds0tNxiCbECAWPEQzdYDan6H9OXdfeqchN8i
DETpcGlU9RcoFWDW4i+Ys11xPIp+OCRjeZJWbv+Dht4tvjUfjgsY+ziHgmJLoLzd
/mnCMWXLGaAwqTUrOuYtXzzqvioayIpvKYlwoqFj1vbNaYXd1lXK8q4IgFMotMvQ
caRQv4tkCh4f2AhLeDQ3ibvMvTwNPmtPSXL4MPNNLUesDUSBNKKkuw50KRAn4is0
AKczuac0KnZCF5z+G7gQq0UEw6jXt11ENnCxO5C3qPeESA4U2P90xfKVeVYmfS7a
aiRNDOTEcKqT4sn2XdcfGbTdXIAFifnPjusGZEHvxV6xQ9Li1J42kRlxuYSmuVOS
Yfm24s8JCf4+JJru5E5JU/9ur8RcafNgvPDHPNhNi+8kD3qbFvFPbXP6o53kQual
6rGPl7ypwgu9Y5IPH+CRivkbVtyKadYPIUh2/fcN78ZMSUlsOjWmOxVHtkazDIQD
EAte1MzsF9tysBpNScpqYyIWA7NNmBVhKorOBva0NL2R54LQxS7rITnOWgxamtwu
2HtcNmTxNx/G+mhfB5HzXzr+gsbsJarrja0aPPKs/l9wlker2fYS5hrD9G82o2zx
/wvcoD4p4uhY3AYYNaue80DgeMhJBoTTgR/zWcxZ4eOFrdC1n89qZahIZ5DcKVAd
PNwr50u9a9gEwteXQueWyxi/+ZARlignIZu0dpWcond6F6pgKfNd9mgdEJNGgdBs
3hvu0hXRcApjsd8+FvrQP7xGKqScvQE/a9g1BXD2DR0dKKO6uicv2gRocP01gNYf
SzjQQjm5CRT6pK1GrC5Z0ZoUv3Q18MerFSUzMMc2wdAyVuWIlp5oUOtWyiT/YESJ
L5JJp7IZAvMBJXHVxKuJpVQjp7o2efzVc9mq+Tv/YwnZtrhtKTKDJJGCTzPchbFq
7FYKZyLTpFbPI/DVr6fQqex1OqbSkLIG04n6Odoqb9WaxwYlxY1noAigHp4374Sq
OFgf+eFgHhNo2YmoY53vilWjUbK4NzZT1zgdwZ3mCKXHeN/PBZQ4dLuB8riyNla4
LJsYJNrA/6t0a2W5UTc7KzPdcvW6EgRHcPEp0j0BUflT6hD183urT8jwI5Ot7RZC
wCOTUbb8DGqBzw2x36eZJ0D4m8kvnYqBkK+2vKIpZ00O8Q3KS2F8+KSbRQF3CeMI
nNuGvjBOn3k2gBXT8eDDS0py5jiZWkJnQMl9QGDR9r7lleT596R5aYuCXfe2h7M9
qcNvK3b9eg8oimMmi/qUDrZ1W6Ot8lh6Ai/ZTRzyjU75+nYAKaTLW95LJKhxjhqb
MS8zsQvu/dfxCIcYMdVtAZczVLW9isCDEZL0/KxrqZyBfk4Pg1PW/Cn+i2fT7wRG
wivCx6lapyPowyHIHDicuA/e57jiykrFaNyJKlSGwEj8ZHZmlJcu27UV0E2cwNEc
huq/vlxqliwmnnn38e3RfphHChWcE6//Vw8lYN++KMAWeeu5F9Ogh1Z4mJzqKaSc
Kg8IkUlMHq1AZPD3Qey2JwXhg8cFYXlXTEbTDZZ7HHhYbJeO2I+tLdha8nBUDC64
f2bG5axdRaojLY/6pay7VehDQ8OUSc+jolwx8ZVMtq0lM/EO+NIihFePx5o/JYik
awZqM5tr8h7/Q9EzzZOBWmTNVv2X7pvSnH3frXWNrJBjyDuXAiMYAVLHjMu0iV9d
2by6p4LPEO4/Yh6W92Ptt115xWRej2Mw0f/tpkAYSubLQmaQVjMGcFvikBnS8F9w
oYvL1fA0YkXdZlFJF7ojX+CdiwHqVcZ1VAZefhOqNI3//SP87lEVUeLMPzZDXxWd
Ex6Y2Ki4XFwxxecsr95l4UHFpIXc9VnJ8MQe1jRYWaqplzC7RCPP18cMoWjNn/4p
twqwpcN57iqedi8d09mjdZXfIfqrwccNmv7NsJWR+e94UWYaw7YUV7kXoEs93uFu
pz+zeZssuhY4XY60nx+oZPqySbqFEB3J/Sb/1S0Z2fmCWzgratVAvseeSSNBdDkP
PLUSIflVLVrzHUAlx7XbHLrIQjoiSHJOQ9CWGkt54LxhoYgdecGeWJ4V0FMF0qpJ
Pqx+yt8MNJZg+z/tbbD9pyi2bIyft+i5HOGUEPV2yBWFVwYLtMsZ8Sq6iTqxazLV
gXSoQ4iLLyMh4UfkaZBqdczhWA/pf8jtSc5J4DuVkvCxWU3RaUBvDRJVWXvSKpA0
ggfsqwKZ/T3p7/5UW17cGPsi8VENA19pGdRMw8AG2kCfKs+2bHtWsaCaqFYI7a7l
9aaohZ76bdLwkpvTt1vV+iZIXl8KolqEM5uc0jqIoa21gXNXHpGbRLOGdoCX3WhK
0lgoQ5HtQazpRHDqFPVCuf8xm4dTzX5F20ua00u1LpAaKBZ3IHHqH8C/POqbAZZp
enPDRGOBRYFO83ZzgTgGzTtf/MIPDVFg3pLg04iLTCGtXKU/a2uFZobshROxBuRm
bc17RSGOxS21VL1QPs580EbEXfkmRB7guiLqWunkwIuXsBqos/hKjC1WvvyPz0eS
L69VN8lLNuiPzflww5fzlkBeyURz1W6PbjKkGWBuEVMSh+ymHqaPoSt6zWwBjeaL
Y/ZsVPVMVjeaD3ExtxqSFdcjr3BmZwBu7y9v9RX+BYeziGZJTWkBXM2t273C7hah
26yufUEkA9Kv1ko/cENl2z3R5RkDtTkIy/ConHd5OfMt4iZC3P3SGcz3aSB02Iua
G7gFyEsdZNAeEAqMIMV/wsDsohgr3r6uBbypa2vn8g19Vmev1fkoOiuaB5OJBq5B
cE1E+0H2JIdxXz/MYqMMaNa5jhA1KJ3uRzKHZhIW1dMniJjagThUDoVT977dJq/M
BesxwrSsK+pwJanVB8ZqH9MiCVHMYVxK2T3yn2/AejfqYf4KJ8Ux6346C6U+tK8H
BD+bOahBD4SzKvKQ5uTDVQFHPU8t4iXd6DFh8YFRs9WMdVChCVC96jJkTQQkVoLJ
8PF8bm+Ww/21wZVM0DtbAxVK9ZjTkAGAvsPZ8Zfim3dBrOtISI+o5agXgQlt8pQ/
3j/y6hdd7su+8EZGfpLb38u6uAHTTYd8eWvlr9ibdzjWMEK/xsjZbCY9uYebCBOM
DBIXUgyJz925yUop+zMHEuSfWvFzoy2v9Vo6yN91tXhZKhvqT117LjxgV1F9td9t
juA+QhDStp1w+vFP89SXTCzvkBlcETKD968kU7cuX7qGxhvAPhUr8+ykO2/Ti3sO
lN1Rpno9Yr9UEU+9oNTiW5m1T/6FKzHN3c+c9nqT1JswV9MFS6SmnvJGGgwoQzwU
17iyYPXTBTMpl7/1CEaKeWDoUMHEGLO1XK8S0xswKUOoUU2KGhzbeZ3RsZB0R8JS
/JqxEHdDfW2JZbdprtTwcyaTVbe7vabUC0QVui0MYz/DB0nUbIPRKEVZGrkpdk0q
2EFZAK4QoZzqQBDSyRNh/SsWsTtj+FJuk5seISkABjW+LBWRLFXy+3oP+QD6jR3w
8rik7+6cl6T8YmDjqdfRiqVCB3NKHr/22VxffDjdxA51DtIGPxTW3z/aSEf1Q0pn
yy/X4uBOSb+ql1oM5LJA8snLJ6UwPUNRda+xk2hQOXnigCIJ1jIBe2T7tl7Oh3JY
yGU3HvmUBQmv6GWjpD4kdZkE0HxxLAhdQLA4Cu16ZbJrwesl7IXoBM4uZ3h5A/c6
qcO+F6EtuNFvffQxnN5WeyBjhQnCSIqkJvEGIjlh5LEFWxS3IsOmvH6nMuZJZ/Gg
xD5wcsXsMs4O5hjYgvBvqBRrhzPbz2KcVFsf9TFAuFmEJr+jF0xjTNicxmlQbIfx
Aik/IRjMXAXBN8n/nnRWBnF0ZUdxo8SIAWaW5nSLDnFYPKD0YmJ/Xjzpdss5IOPp
Vks+aiCCMP96wzfpEWfxMjbfVa3NspsiWGVc/7bwDaXOFms84+bnOFu2loNHw5+l
WFmDlTh7v3pFA8G7UQt9+nS77zSs9vguKUZV/jwT2CldILBI2+18+tCAyrfJXFh7
ULqQfGc6+23ILCUomPOyQdpNRapJ982ZfxoavRF4mF9ElkdtOvcHrnX5V4qNIDFl
4Ph/5m8XXdiuXO5kxjbrc7rPSJiZYGUio7Ct3borTM+lbGCAWNfxyi9P6VCr/QKD
Tvd++AbC0J6S//xGOAvZdhcLr91aDQ08V0OqBHY89cDqrEr5p+GojtxX7qt8Jo2a
MyZOkQcC6uFMrJfkiSeQ1GuEhlvJgyO7Tcbst+4hcQXWfJKZaAVP30gk+nqc26cS
IvZ99XheBrBTsTNN8echyL6yJ+j3V6lJqbtc6zxBo3PQqc1rAyHbHOnnctHHehlm
9detpl4i56F26s7+2/q8+Zr9Sv0eEiX5N78sguVi/J1gRc55ZF7uBDcwgeUOJM2y
xN8xTXmRtGFvDz5WThjsXhTo7Yah50/0Re3IUSfL6mI0X4IEoDHElVgub0PSwe46
o2OI6uYvvGzyTpd81ns9ql9sFGYBBGqFRSiPL9FPR1tIvmp93es4R4XOxcRJHXok
4if5xSgW5tztjqcbmCwUvvqc8u11lbppUjgo3npQe0KE7VFwYU/VaI0L73C7+T+p
FsPIcyjsdhH4x8+U9ql6wn+pcy+IQ0SJw9QnbgZlg+SovF0pYwYjh8+cJSOanE5p
HHR9CKw8BkM9ZJYwhUvZI2AH3YfY5IF9wGVuKnlzK65qWIpIjdIk0iDuwtjNx7bL
erHkI666DR2HBBpmWIm74tjhXDFX748q3SR2nggIwdL+iEwiR3yVTASjGbkET2KB
FuSgOI043NT6BJxCOW/crqU97mOc8Zu3M3CNRXzMY3o9UxuaMcMmr5EVNORQ9fAb
viK/nlnDMLF6vWPHtB23dqgbcMqRpH1iVaVOTA6QfvCpv6JJ1R+4w83fztp1btBL
cKslKpFLWTD6Bppo8GWjcPPdK2orbINP7SVEMc1qhYq1bm9ueraqrlebXK0wyV93
6KoPLNNzO4uKiRNizGUYWRbChVOXNlq20MeoracvUirrSbQ3S98lfh0qX/0Qs239
IWxiLutDnQw55lbOGFr0CEi97r7y5B6d7QSfRsVzkVm3xRkC2ONGnrh/O/enh7nf
/xHAwzFJ4Gz+2o0xmgJTTBVNiTMPejah0ji1WyOv6bF5ieQscQZvY5nrxvNBzQ7Y
aOQfSkBaGonAE0tCoqBpLLqhKV8aklZGj5UkyRhyza0Lv8ywiAN1uCjcaW/vT8t4
1L1PodjTNa9wluB62xgbn86F+YouDoP0755pP58WS+7TqoNx17vsC/TiYQMG8ucq
sLwVY7JmSJ6LKyoFfjjORYJDltfhIVhCBEqdLyZUUg+mX3OMMH7HnAFPmZAS4Fvm
ShnPHGd1jTqpW3JcwQFSCIViGPUhMulDVnoO0aYUPWB+xpIppX1NAgTB08xr7Jw5
HffFcVoTarhgZ26kOusI/RaO7nvfJb/H1xtKlrziOK479yK6Rzs8vnFHXyFFCF+y
+XfZfQGRFMahaXv8tq1AoaZls4JW4OGuli3JzEPbq07JtyreYOwH8GYLUqtGadkN
QDMTZnkf13t1Lvl/u9Lb8meHkw25eYHtgpd5HyVg6VEl8rVW2JtDobly8fQ1q2Uv
BHS4/AXmwxtBQG7sOgTmty6lXfnOr8wK1K81ufejAW9jUqEPx27Zg3osNpTe9vHL
LK6YMzRSFIZn7KFxMuYQ6JyoMDLkPAY/Vn6RWyKtJ5CQAHDwapGTSh18DxOl4uve
iK3F/QPFCTXuPyQN4+s+HnlbfS8sNBeO0O4UiFH8FOlcnPa7XJcwCKjGdDF0FEMh
2nggEvLU6YGWXuwLSCZsjypShyH8R4fikjpAtvxA4sGCblhYYPY7CaLrWcoQZhKF
QKtfygKaS9TQeKH3vK9cGOc6KfGDSUNWvIHAf0TSUK2Nl8G3Ewm+mJ9e6s83baI7
JomH9ow6nPCr6drGLPUBwpy6eEDcBFTrMvlm1ZtxPeSDU0CO+bVfPbQMP3hDZHqZ
WsECzmmwrSTweYICstW7oFP0DxPS0XbSJlj6oPXlLwUqQ7kj5BHPg8Fb8Mx/wRae
8vvOm+Rn4R1VfhkkaWFMJLg2pC34KBcDBpi8tD/sTR/JW8+EZrknSbUAZXOC1vjf
Mr709lu69w1Oht5H8Tq0JmYR0GKifQCsypBW6erjHTxoHbPAqvbG+VoBYt9xWCje
iMnoSr8V6c3/sxUB/DDhlRlLtjOr6qrLDqtVc0/m2YykSt+j94uAMK5pj6jzZIK8
fwfFfvsR+zhb9gn0QUPy3m4Onu7aABzmPKXsYNYgokrw5d2orliFHDfJ3tP5hWZ9
z+qeAoQR5nnej7Vax1hbE6VLzJlyHlnoBYdFZv1SqGl9HE+L1rTeqFJd40RIIlbp
DD0j5zSlW/E52eZ4QosrACcRZuamX87RMQ6p8w3LdjpArI4wlZDoiU+7Gh821qlu
QqfwPltztJQ0MtmioMyQoZxfDWSTN0CH2Z/YnZqlk4CnaRdOye5JMmzbqjozYPYv
caBbtGryXX5Ly98rpTP30sxyl6QByYYFGRR1C+hWlxUtK4ugoa/QqoZKA84yjaCI
tqaDh3cguuwBO0D59e/A2abDSEcWlSQ5F63F5mhR5CHoBabYkLFTbQXe7ph4ZlZb
MeZRIlWUL2W2Mq2dpO/mw5yotkEQdk/vcZ9eJVtmSVkqVUtC6KvEcqOIr6oCYce8
yyfn3uH4bGZXYGFWLu1O6stRvOgYk+uLhnRdLHu89PuKF5aSD/8MMC4rq+Ia8R56
QDOuOS3LyadrygTRnppX3QEopU9f8K0C0CQpxJxJOTf/MOSH8JjuAZ4UgTws1jaY
RWOnkS+i/qmGvKbvsucVYcZ9kAm/JtP+b01+4HETy9B0mVhMP3jX2hNAuafoiiyy
whF63i68ieiL8VLJEUM0YKfktn/2VyH9BizqkX5IesBxB8Ux64lwFp3RcKY2D/pc
CQQ17kRWnirPRZpaneu1sA0wJwpshz0Pei7jglqxG556Zewau3ei892trjXydbQ7
4/sqi9Aa3DrZRvMvkkLBzthBH9skZ6yFBL4QiK+I210MNgz2IM6UwkQPz5sorLhb
p9dneD4mhcceYxOo8a0zl8XWOGn1bObFMdO9TLK1K6JRr5eLpHmkoZ1uXZ8xtocc
f17dCVd2FZ0Ij+12VFU0lh6qGMVuIBoJHrsH8JQhvmGfaMtPvCb8+UNxqBKvfKqX
YgixijOrmmfSH+f/E1ou9XY2YtHwJ+wAs4FuLhs4/jc8mbBqCxMRhMR2rJH2FZDp
RbTlPIrCKdXYHXvK3BODh2otqT5MMJpFw/kMoRU3rz4J2b5F0k0F9fHk5XPtG7Tq
B26tyBfD9sc4+W0r7eWovL5Za9xuW/OjA7048lz8h9o+LOvGlrjw4oYWl61qAt9I
oMw6E9NtPtn7SWmY/zwsW3mmFZwVbZT6ztoldCIjzrWdnQcAv5bVY+8NIp/CTJk8
rCP40Ey1x7xRsp7sIVr1WM8PJPsTRyo/lCac1S4WxNdf2WvXwP05ebpkhVKh2QTp
U2Bym9YWityBSKmS3zHWzjI/eFfQpX+qwqLWN65rjVtww8RDfViJABVjTi4VEuwN
XIyPJHM9zdp5CYxZ8nHQxYE/xpIV70Julwy0V54HxCvJlSXlfPnlMjg+3Quzl7xM
QaBpeP3Ue4IhXzEptExJF/MjGl6+spWe4ViG1JjFErXhKI9lJJp0UkAERKFLit1N
eQBbbp697uT8eay2TFvD4uLupMHebQE8gcbWh79GXjFCC12JGj4R2sIbm92iCOxS
7nEwQ7ZXFqncxUVwOIpHfvxsWrarEp2SKVtA5WGKCvaG1hB1j6m764m59B0jwFHI
LnZGtUtzk3+eBpDbqQHlodGE9wqHxLPzptaYEzSfSBPuEP1fWfpTkMrnFec0QUKJ
69J7i7oHK1ZKnLQEbarXbAVkrvn4m0xcv3md85AWTa/LGnNNyYYEOb/kEQusbskZ
UbGlZOyIiyXYIfDF4quSku4ssMcKc4TwNslkeOfziM67YIX9RFDVliHUZUuPEU7+
aL3e6u8qLK5xaqEr14U0mzSGRwfRBRE2exFFiF4n/B6bEc8Jm+vDdfXqOH8CX7v5
xDIAZemdLKr09WEnZbZjEDLWGqt6drxe/6WYWE0hGyhmG77bPe/vbc0RRMwnpHzg
/h4i8rtud6kHoihsyWtXFMerY5r/uWVAKtSz8ZuU2qGXe6TfQ/gpCfoMClwE29Rd
8SposDlA9aoyfrS3nfZV78uczTc5EHZZWVOtvImLZaXeXhD5P0OJifPKnXUG/ZMj
+GryBmQ9DrZY6OadTFy6Qps6AF3ICoEKwdS3iG5uG9hB9b9IzkFazOEDWdDQOeRK
xXuQlp+m3fBig+BPRTbuP076Fpkr2w+skMa19en1r0zSFfHZsUV/8jBmRs+dhPaH
3ZaPEersSxDhcEOYeTznp/vP26ZNFseZDywchtoBuavwOXFI5cAjvv13P5UMVvhC
B5xpe282K+Z1ccfvxg4I/giVyjH6U9YCPeHgSAoKnl1fedPNOyXcI5lQkmoL/5tp
6IWrmlyPG+YWKfrB6nfbx3iOjPX1Ikp78XhwLp4nJId9xgM+1UCYwGM9xbj8wui3
LBaYMZG0bfR8l2p1O7zPsiupQkXk11GTtMYxxdxbLOqOr4DUqKMb3Q0GE7pGIRVp
KXhBt/D3YvcOMauLtKlEaPe3bz3pvI7zc0rGKn6MBTNL0WEwGh1jlXUPys9nOY31
Skc9+RX3l2RG4qzrv7owYDy8RCDmTK+YMHTBkY9ohZSIB+sEWWrl2yUwJ1eDqyOU
A3KXZY+eLAm6iInEt7SCSF0Vb0uL48PCk6CRg/zHHG6TbAy8AR32AzG+/yMUlREP
SPXWNGAnX2h2lFNoPiGNH82y08HhIpvmiHZpC5iH1D3LLjnWUTOi/OGsJCXNh3Z2
JYNGRd22zn6vnY9uKKGsKObHD/1uLs6yRrXbF1O22RFfbX5VYCGExjqfQ5Ziezoe
Ruek+SAP6FDwEMkAD5t5RVECa4jU8SCGgtO4GyPxRBkjHG5SNe94g31NQb5jaixJ
F9ciXZnnJLK/Dt62/ZgXixAPgWg4X7Ew8Fa5GmJaz89BS4QH4oGe78fv+YTXRx9z
SBhrWVJGfkMOv/9/B6N9H/Aic/VpcWMWmxsdjXz2P5EQMJ/Pu8giXJU4TakkApOC
iOej63WkuUGfiL/gUrplWa6yNXqw6df7D3yanIarimdrwx5pHdV17J9cZc789WaJ
vAQqamaZ8cvbvZv3OtcVs1hsGJ/f11DYAJFSh7gMcGl5efZbj6TLc4TE2iGGYhWs
+tZMj2aefpD1fEW7zcU2cfrNhvWSWsGSLUH7BjPvsVK+sITeQg22Wv+O/lM9ZgDi
2a1yaQJP/IjpJtWF91X/z7kbFJOjdSGoI9ctSMX7bI0iAvNYIk9pj5K4bozF8YHv
vyd/4xEIWfw3wtIeYu1pv4tv68VQ7XsvxDArmDlzyBdWzA3Zd1QMTBdb0ceS0C30
aYSrNw2UgaEakCMj2lavCf+cPA35iYhMzyK5BGtRHwbnU0EUdZsvtur64pMhVmUt
ddxZH6IZ+gPPQSHqGPLwQPqS0IB9T6aBP9h0SQiFtSPcFHn7iiytVdHaZ5FKM0UH
tszsQApEMTKZBlS5P3dTE6jQY2aUrz/8WwHshloVaZu05DWzH6083R7ZGNyl940C
C513ukXNEihFvTTdWEWwXIUQLC9ohS2jqh6yQCI09p7TFcBzFZfR7u5o/pxVFdXV
ZvMynwmMJpQTBiNB7dTKs6lPY6lvRxXT7G+MaS2DQlFsohYESk6d/zbnf7sFhwQW
Ae1S3nrK09hirkXU7dDlRqp9PmcuKnWZE9un4922BdQSuxdhpOQ3SRGbMCYoUyNF
F5jq6damJk7tPb7fDZ5FsD+LR14taL+Nnn1g04YKz140nPTzSsoVQCO8QKyDZ6Rc
QCEOfbJ1b+xybY/13ppW3S2nmuaVzD6vpBpavgqbZnjzoKXQzfpvtkKhA44NOdiE
kdsZT0BYc88uClQXMhAvfWiErUWV7lWIPeQJOAq//i5kTlmnVccNrWmJL4F/EDyA
0BzE3rOTIg058gs4j2YLfl4TPpNqENaHCVHzvozSFLxTZuXExWJbjKAqHW0Wgupt
cpBctXo5uN0cedIClOHN+WVEP6PIhWRRNwUxLNwGy//0/rFqTsUOcocZFRXsp3zV
8Mxt7P2MYeJ6xDNTFDqZbMPDTx0yEqckBtWv+Z899yklGVo8SSQNFOYnKZY6D70U
HvFZv2iXZV0Llz+ujD1leDOczD+qNIN3Ivf2Jea3WQDjAhRdqUqSjTn1IEoQ8arM
cSsU/eR6Xcz9KcVRlALsVcXJ24h1CsvJ0il6Z4nyeXbnobps6FjFrhXlIsNoDGMB
aKhQjQ1ZhUjXw+ZNkZ2jn3zi1a3lo5+/UXdHEaNzuojXKTQO41goATML3M+7OhBG
xPWV0KDOVddsOQu2UEZS3/8gJB3dUT+FwjgTzxi5NueCiq6Ui35FN2Xm2Dw6BIMx
6vwzFW7fGgdxl6tR0trRLaNKIzlXelQUToJMUPdRVoJ1Yc/yaT7R5/hQ5e8RO2Lr
zLCJOx3500k00EK8LNvr+mUaC6lHL/g3MI9pSfeZMS4Ks3eiJTpihjBj0Dn08NOh
fomczEMZDMv1qD7Qhi2VEw8Ykuw357xSPwzWmc9n+647zv95i2W5SPBp4/WccpES
ecUO1PfgtRu1uaY0QDHQdFzGaIvgvlm+vZc6eUng4uJmliPdVwPKe690valktxrx
fP/FG3DYT7rWVnVihrA4r3Y9qcH+MU3zuuJrEGiMJ9PbVOL8cVeF6rrKqG7Rqgbf
He4GIKiB/xWlY3Cf9iiRlIBHfiIPxWmZ+cTUriPfUKshrwcawCFVXusItvA9Nd+w
0V/CYbeYUgL6rGMUoy9t22CivMoZ4Vs0X2IhD+kW8rIqxH4mHqVAtnbWcepFEMcO
3tc2yo7aIfDlPeth7O6XDIKAqjviTLX5SCjvx0Wxy4AWK4UybooOyxAMTQvuDV1D
zIpTEWSmMO/Qt7KmBixkwDgVhxF32K7X1G7D8vLardxvKzQR+oEH309k25dJw40k
+HQ1wqd0Ewnr9BZi9NaZp4iSgcu4LqRMIBZsiefojTp3ciDa0Jjqz8WUoKZfiOpZ
hKcLHd0ZFy/lCToOcYa7CIFnrVf5zkKRPP7MnWpbT6yLsJVAgw7vk/NsqWYni3C7
eE8NTdsj7dwiw7F5ns9E5mlspCr+kbO5ZzwswS5i8zOwrD89i5x2ZUwvzZWAwivR
yI/hDdwzqPCIhoEZZpA/BiNl9eH4cEAPhD3HrobKKqOyCOZ29u412cUTsCZpgFfL
yJ9i6pSAD3Tnid/AvdSnu69t/VHfcFqJuEQN++kVWwws9dE8qP4TKaSQV6V565IS
7Oc5Tw9WiRCDoO3B5uXhVhwK7FB1mz9MGtljXIx8IulBrLU2TqnjQyzv2G7IfjMR
M2EagHgxMKihB0T7CDzDw89Po0mkYf9b1VIgzBDVOm/HO9gKdLtWARB2hW7GndKp
JBf/Lfz2OGynCW/fD/ZbRY3HHxr+f5QzfqjcVZ7yITo4jLUJpBJVa3STVHs4Sz7L
zYHuwv6+Qz68baGXvrZWLOVylVnV7KF/EvSGxAyvUl0qiF43HC/Z+tTvDgNpuaEi
LuS57k+10gZq+1Ow/KtgvKssrdU+ctdKBy+ClDq4BjcAbtCOwQyEBQYzLewrQ+Wj
jd/lAR4ZNP79S4jrlZfjAiUoD+KpiBDumQ6C2dtY2ZLm21mU8LXs59xofNhLOUYO
qUZopC5+j14mziwxAsDKD6yjvCHENSX9N0nP2DKFrnnNHvERmkEMXJ+PUGx1w00P
+K73oG5+9d77xr0jj52QYJeGjYHEwBiPl7kqNSD4q1YyqPSTq6+S1s56mL1WAX8A
qHJlOFOiT9J24DpM7ISzjgt+M0ryIEt9p9IyNhTWmESMsGxxNuJgwIvscIp3J/+y
lSCB1kCdYV/MgsUmytEInGdk5UmUx6QXcUlIte+WoMQ+jJ3pGAw+Do8EB0isU8ku
8h4NybH8KB7wLN28S4/6ybiXigVNlPRIQNhR8CyCUOGPscE+8pcMs2yjSRMXar4I
IelUWFYXZpiaOfiYioyn4YzztHyhhmAwRDNthJ0MKkcQsxNMlNT5yTiINO7rP57a
yYdDS557/O9VrNfOx7L11IuLSpOZwlMfI02SebOP8Gs+pdy4ZhWF6X5+KsFQAyy3
jJyxGInWfJoJm3M4NJEBlRJAyiam7s9weJ2ewPJ59yTzIyrr03CEALX0rnVfe3rS
RHa/4++JlOw3QIkuJMDH3klOCqlfg0fofU0Oht9Osnj5VQeeDu329x6OBtjq17qQ
iTZug1utVcHYkadaa7iRZyMcW+vnCisX3EskKILueAgD5vJeIGrm1EBmFUqiYxwC
ymAckW9e+jJ519rysX+7fkiIlzGp1oEpQBPN1Pf4eYiQr6hMB2S5da3fIjz9l1Gf
LozJ2td5moAptmBuwTnOXVi3ngXWBtEjYmKQHjjbqo5eZfDelajVyGWIUrZ7SSYa
uD3MIGhrBSlbHK+KIJaOEQbj+ajVKZVrHrM9acCZtMah2h9wjcFPLA2TxcVkTWis
W6HDCijbSeVK5frTnG+udW7Af5FUOqsZ4I88MRYfvt8QQNYlFMQ41+kvWmSE9YCg
uXUwf3CQeMp3p0ITHNxrVogns96hMt/TK+h2V/akWbBeyMcqdFSIjF3nLyYdPDX1
X939E2/IRVgWjoVhnrHZia8ReorKYQd4BHOZLLGB4TS9UZWY+3Daj2PW1OA6aO8Z
FrQ92Of/79kR5sajTsCLqax263jsdzA9xDg44a3tyzajLDQu5LUiqvKH7FADiNf8
m6bDTZmB9fHWmitNdEzxlmMDk4j7I8JSrMJslCvLgDAoo/rTEmHDHWqPZay6ZpUE
G2e4Jdp93cQBYGDDGqjmtr1Q4e4Dbm9/Y5eN2GPOgCilyHm458r8Ps7QnLYvIs4p
fRxnaU0j0cECKQD2dF9m9rnDHq2pvbdMWWL+8qglI6ZUwe+F0Cn2rRjOMQnMF1DO
uY3p0b3FfscfqRyffZKbFFp1k88KV/zlqvX0AQcbJ8vihQn4R7OYqaPeLK7GuRho
vKUyzIxJ5eX9TjxNjw7xMvbysrAavrjMqw+0jXQaJr+LGAWJQY2LAza5zGl083GG
Q6K2DKzmQ1jUYXlCdx3eUqgN5/5g3PcQGgmNm/ifM4t30lpFRxyBEGW+UDrSK7k6
qqd7HO4Ogp6igzLnA8RQa8klmn/AMuwC+k0uU7+2ROwS8vL8R6vd3UJE2X4TPJBc
pWzECaQCCRQfH6nOtm0gPKseqyAmsI2z64Wq+eyuxJxU4dVTzzF5TC12n0hPs1JH
jY9RTpyYGq/4o43mVcOFvGwEflIl2OjTYajmygOq242K4nOo7UP7yNAXxl3M6p+W
Z68oXr/yl++D5LABmS0KfwiksieV9WQw5dVJz/n+nXx0oSrTbwRxuOlROlIUt/a4
vNvT07retIKkItLW/LAYzmC5GlBm5CeB4WJD4fAwuQ3OA2uMhfY8g85WOIRO4WT1
shNIZJKs1++WJCblEHEoyKO0uSpV1zxHfCWBmXSd8Ruhzm1YRvtGHmio1GIvTkAb
VQwLzo0ouCYWCvLB5ev9VOJjgF0PNBrJVYyc0pe/5m/XJpmfIh+92z21Bq9zfR7L
zXbsuN3rHv1McO02nSxaULpKhq+yekJCk/Kmw8oUqKaxyMIvJEgtpxgd6Siqi0em
tmq/If6DfZ86m65LbXQu8ZtMa/fEdaFt6Tr9bPiTqpa0c8dfPQ3DNRqlzuCagLYq
fsvKmBNBu2CsyqPc24IZx0jYr4w41IJoicx3X1HWQS2Mk+bNa1HUFNxzluxsIg5i
7O1WyU0dQIHQ+BXHgEdnM68ijdJqNJrW884BZf7HSKYlkFEDJI5cgSI9YI1XnQ9G
qHMuhKo1ZhgtHXzESQOED2eT3a7SsZS8rBMPrAGbXR5BFsKSsZzVA4SVmcqIZjiK
xcsfZPG+5116gGoxnl3/YxKbgsM/03TmIcfzr9O3BYXP2fYBgZWeZ1bhatEarBho
/5nl4KYxRBh+LEZQ5ajeEPXWFhmCEfe/fHdXnac9JVcrMdbrW9uMRKjBz2K+xHCU
MPDNCUnDkZI0GXEP2tdyM4opyPdC3Wh8fKWvYX5BINF/XpSLz5GT8WhZwuNrjZtv
wVr7/IIzGCXuGLZjkKQ/hS/nEp68YZl33PTKzMwDG5Ly8uxALP8d97MMMHLLDCEF
L+1NcHy53krTKhv/vM+0Mr4DyJujqCKLmo1DN8VV1F6vnOC6BDEbyE+oxi4/5SQx
67f0P+ziLrw2zI5/pp/4Jztan7Az1oGBK5Vq1xpgMBE9pBZGH/8LemQPQizmi+tf
3Qydnj9AeWufREY/yIjBUP/EBEYRcDUB7bkTw5Cr9oYHxDVicNuhH5Mdrz4GWt0p
GqUzLWwzcN3ZmYDbdWPoUwKe3ZcsoSL3yDpg1Dv4LPeURKrQCdsRYURzMd9X9Vvd
cm0thp1l5XvgkHuuRszEDRcJ38Vz/6XgQnHTawP8wiM0jxufTkuLEoLmbx17eoQZ
vOzz/Kso4yMNohhNVdzGbCE78TZnIWq+ObucWTbbrQu7qYNEB0tOouBZi+IWBiyx
rELacEoi3X6m3f2Y312dngNUafPc8Ti9WXNEMblYXz7ZQs5o1sU1xVjdp+gUqi8E
o3nq8pIRujrmN9fHbJSNHV8B8EwWwrv/loXMKi0Yi7fGTp30LIb33x0gXru/GkDV
gnPHiWL1eHfn8fjjXW1Nthdc59Ae5j2ivex/vKNdvtXHEZKzgmsvHeLuozp/K3bj
1hADEM+zu3cjgYiovIHXWlLee/o+T1/bEuSPfH1a5AW9tkeLiiTXvjlFCXPB3NAO
E57bXuHMgRLEVs/ZrOZe8voXdd+KjIF6/l6MfrjcLSMMmP9U2noxpY6qQ7QSctb3
ewOMwdMb0aMiFrd8R9A2Rgy7kgZsZjwdn5vHRXBULMgPGUPFf6lqyHbpdaMYle8y
zGfx3NxF0wm4arfXKUIEO9fBuqISN3J8sEyjDEU2PCm6+ZP/jWYjxYqxEqeCrxtt
Q53rc9BpOEBgoosfCCu7IhtdvNEDDhCjmrU593zSn+4sueChXbC8UTNza2KGdYnE
xtiEEcQlhiXGwcXgmLZ4cqGi1H1VR4kOjGykdy9bCHEaABH4ODItTwEa+4HVWYTr
fCY6YCPVObvXjYtjLarpaoh+Qz/SbLBbzGKX1gpE+5VInz3PFtuIpRBVC2MHsoWh
cakITajUf1CjBMYKbWjoCO5mj41EPSozU19E27sMsAXNs5iB041hHL2GGtYQKN2k
bx70Y8j2BPnF3/8MVrHhYSO9f1DopZzq2A/g0hJCgHDwKaQZ5E3EoSl+wuyNKOxu
6aPPsgqUCi+dWaC40QvMQj92aowI/ykQw5M5seiRqrt9x5cf761c4UhGyt5U++5P
8lQ+s8/DT0nzLJR1/vLCga3QE4QtAYvOxik1CgBzgBukLIGaYUmFxVcSWql0fQY/
N7e4vUBPcG89aJ1ZONxD99Y9aCvPx5mjxkazwgJOfImQTqqsR7k1XSBnHL3zA09Z
b0qEf+3KoXwLBKJ5KGyKwq7Ml7PwWGNfkIoIUAn+ZmMM3bN5agqMo4kmtvmz659b
YLcbYD2UOBprUTB+ZLlMVDfKoq/NV3LVQ9oAsyIyhrrdKtXKkDLXDpIS16WcBewb
Da59zeskrBTqJAXnkgpvTgnC45iEljWAparWuyyAXeO4lxjDJsaFfWDyvTV4cbwv
kLRuJPmDaf+rev+I1ylC3q7e5QmzLpcgfHDQX/YHP1CMeSu9y0w4k+sDOWHO4ImG
88O1a3dI46MjXicyv4verm8wf8f8kK9iX9oE2cxNxn1XqyBeoA8SMeCJNV7lx/Tj
OkICBFXVkxRxLf7E6U/UCDPB2Z5RVdsF93kfLwFhB3MJ9R/lADbMtQKvkRI6VkMC
mYqtL5YMHdCFdBOCK/WNo0+XC4/WfysYmPySlv5kWPBDOZISfvF3inY6PlVDx9Su
yWxBzjs6QM+J7AsWaCF2FLUsPqVWNuLvnPsAPjraokFD++hb1GIkSaGt8quZx48i
rWtzyRtu613FR59v2SIBYKflotu+06Bd7x1zbF8+LjY1NefzvEbWZMao6isXp15c
YEf+BTf2kS2JUUSj1gQ3VvKpPsWcTbxEXPZq1zWbRL6stOZ788S6OjNyMa2//WJA
hYSAHFmI8GGiSRXocw1OS2y+tJpX4L5G/f+yr0Ug7slbg0B1L8bkxezNIWxs5H7Z
vZhbSi4iNz82Y0kMqCy1SMH+K3KUZgewRYP7Th2KH8t6qlwcuK9rZaklkSjVlSdc
9xh/MX4ilCpajdO8KA+kWBWqvx/sUTGElIvmYbq91aoDN+pG7iOPq7YWx7dzZO11
VG0SyvVRC94jcopkRjdlIO8QR8ysmpd3B8xcReFtRo4uVOfwLrjoa2CO9ZtVNmjf
gkT7l27jlm/un9otHT+qyXGOKZNTXqljxdnPjKNJoILkMuVpSnUmROIECl1Sgc86
C7W8Iz96lAbG0sl0s/IG8nTwnZzdJNPnit8kenXO3P8VpZoljdgIfQaffUgyTkWS
zhcVh16AddveCwlg98saBVrrB1djwlWdfqz5xWhgWUIg3qB21Cw7dmXmLDY3jGd+
2TQa5PHbvBKNsedNtifyc++AqY/elfdaV1v8n88jFJOh92gcDbWG/v9VIFkbtl0m
ks5ZW7nM76mljcPwMmEKdG/kz3JrUBWCpDZc/edsBpBobQ4dbOylouvVW4HNg2Ct
NqvYsJVnXbt9Z5z6KSdlglxpsRGV0u4hUzrJ+ESO/wofZrp1lS9FWjvw08RGCrio
0rXbYTdfnYkNJ9ilai/yQAJX2HYhYwPAWgDYr7p1mfAKf5kUmdJZchPcy+tun7Qy
UPK3q0mSPVjG4FNG+IT5sMFgv0Kl0sC2f4t7DfKIO1H2cCK6qOgeKznZj+jv62Hi
Rjr4HkTU5MuDmTZObmtm7iceqVJLhLdK2uss97U0toYAi14m6kdoGupI8MxjMwos
f2AJ++lr2I6vTJ8jl5fRFmEutG6VW3gRrPFafeXqAK7djsjEFL0goBcAaMZANHnH
B37XCozrQVbxDtAL0g8dG/59mS+ZhpWIoBdeHI/UOzuMpe8WJTZuQhjEHHDasC3s
+1EAP3c/AVcqH7ixOt87TK9au8ZNkWLXzz0rcT5BmofaCG3hspO1kvbKYsjwT+Oj
1OkapcyuW6V03u8NWYUdvGvWYGULINz0Z9yte1MiU3/WDNzKPrXSkXYSuawogxYY
vgYb6Qx177cpbr/8zDdZgajAD30urrPyOxJr66BnVWS9z3RdV+jghxuq8MPYhO1Q
r/fEIWbCLrZahnSDdu74QAkgu6Y3AnJ/0xNbO6n/ZJN9+CKVIYKuHGesFkli2UhT
egPcVrRWA7jx1TJqCZARrs6P2Pc6LzX1h2ZOje0qG5V+B0dBsgUwj+DQ2DtV1Lze
uqBZXBxWXQWzgFSzylLTrTu2EkXdqweXbd2mpVD/C38+HpWCg9KQeJgxC7f66yMi
iGXlhJW8BY0g/jy0Q/k2nbbxi0j+gluDNJ1D63jHr5flDM/j1hQKTHGrm0VPPajZ
0OdfnVZr0SCC9jptrCT6fruXwhwZWjfT2rk2gI2fV/DBqHIwJL3nJqSM75gflOax
K9lJLFRpfbbLg7mVtYoGCzC2hu1Zx87lOVO/c9mhBZVS4ha7qZ6nqDpcZfA76z3T
mU/OT37WzoPDXotPvMewAgjDQVri6Po6iD5Ek8d11+nW1SxZ2U5lgWChDbRcZHk8
96Zf/OwBWC1AvEIMEFQ92A1ritn+u5hDx1X0JMe6IwEvJ711Uqkb30P3AGjklKmZ
rndhDm6gzxEonaiRYvpmrSwYT4Fahk8MQeaQ8nLF5SiszMrmem0sTHohRmEO1GWC
xPU0+xMai6plaVoUHg032XTKPMzEDV7VSifPMYYhZnPjURPdG3HgRyW5Nsd/Zhv5
xa+uGLPkbld0JPAWitr3XeBOC/YqK7TPgj/xzLCGJYeN7KMg12tAlA2mWxwUCnaN
QQBwAK0jy7sQN9AhxoF0FQifD2G/OKIuziAGlRjJ8nfAWawcNSfAo8DU46xvmGdW
UQT4EgZQIoqE0FkV+3WCCheaSDke0yBNO/H5c0lFOBS3VcGArWVB1Zd+KVvNJAKW
lo2hJ8V2fctNalfMQOI7EiBKAFpnq0wMYrKtNGOZ2YkyVAs9+Lt6of4owikknJgN
MF//NsQcxjRxOK3MoUIvRq2WwdIhCu37gQ3P2M2sYb5lcwN8I9MaPjoG0N4iGHCM
wnLzFudt7C6XbcYj7X+mlXMAxlDx0hlSZRKysMujgRBTlz1+t15JVMkTOPtaq4oa
Gys0mnxbhWnVCV+wpyhh0vyQAqkYowf3FcyBFhHoo5gy4YROf0Q3ObgoufxpCJnB
QhLoJAiL/yqzA7tUCMSzqONCjtt63u13EmkTPVr/c8qQcrDEgmPpjnq2F1x/uJfD
xfdA5QQc7yDxi0BCv+uc26NoiXoK326e+DDPgORlTmv9d2bbo50rbxrHIWQLLzli
uN2IqA8hdhn6sRHt6IX9zVatlsxHlyMc1/JNPfH1iG4Bm4IQvSpDzpQ9wj41Fg/S
bdMbVp7biABL8NVdY/n5hFm5nGcpQoYu7jV4nwCCX/I0HGKX3LwdlV3rcfNOrDiH
csUEZVv4wA02ZmuqApXXTgPO6/6c7t8m9RYl6ET0DLYFbVq6yUIEHzrP0iB6LYRd
jZ9GuFzU0IkE9MePFpFGh5AEMp5pO2Y1bWTsm5m1bYF4v+HbC0W55AN+v1wKIDpR
9Gv0FWBrdmFwVgFKQylkCWhOo+6h1r7AvzY9+Hwx0fNFh+hajWPfceuaJvtcqAQ7
cgnr/vwLc6z+IB8HCEbM8Sp+OXHLLhuam9HUipW4kr+3vweMAmuuCbwiaHETcuHZ
WHAiNYn89/vuedvmnuYiEsM1zguYi+zPJHpZdvcrIWWIlkDA9ecb2YncOZnZVe/M
n4Ha8qEPgoaT2xaRgz9XmYGcQ/GywxluXXMJ011gnNYjPYhURYILmxqwCJwjn60p
AyxCcKJxF/AROcHrQYt3Rvi3n+5FRG7lFATrMXH1DdRngrF7kJirIXB0ntGdPjs7
+/iTaqVf2tcDRs31xjILaYkq0DwKapptzeTaENMTYOaGrJJXn7x3tl0RgEDO5ngS
uwpMafBhGjJobbYsoR0eXR2i61Ck1attHKbdaauKCofAlBLCZepzy0T8Caf4l9Bv
xHjj2lj75C5dNpzQQCI90Nbehqz9nYCj9YLl4UPWOMk3GeaRymy+k9X/wdrC0h4o
Stju75voWC1JnnoOnxD7LAv9xUqG13JqXrlNq3uZmbwQV0f9d6caQBRGvo92FHS9
KrrNsmhXXxFim+VcyHl4s9Re7YcqY4ea4chFa2sBJMYBs0Lye2UdaxuxBdqZbdZ8
C6X54IOKhuol0IVgv5RFpvPxbVPf0w7yyKQAayTJ3PQyIgQX5mq6fGsiePOeF0hg
JctP+vOIy8djj7Z7YHpDOg8onVsqA9kztsvjsKQddgurPfZYlAatcR3hcaYOAJEX
ke9T6GmkmRehofmlF5n4tCnB8ay4SIrh8llnFOejWoTrrTlPh6kzGvjU0P2SFcPE
MtiGwpyBJ0Nm91kLO/WCbgDda/sVtUIOYweOZQeQ5iTafCrAv/P3gGNz4fb77hDT
gEMDBtEOcliRotBf8130RdKRH+mx40YtQXOTOwCMtOxqNkUWb9LwZx+Zps3KGpwY
+rNhDOSDrvFBBxwtJboCoHuzd0A4dXjQi68ooXQUWy/jSWPAxxr2u/9zfHNXlpTa
c9D+2P6/n+mHJiOBb8cUIHinPf/r6EXVhz91XwX4vmI1hslXxfGt9Lz3pYda6j8U
ycsRoLJ7L+ztigBfJgwaY1TmteRoWdHdEBvSNdviVqtGlPlUvpp+5jzDAcOlixFf
YPp7hvNq10U6lVqf3OgWxWQ5v8Xn+z7D3aQKTIqdEpC/9JGtb+Ac66SvVPQcmAd7
QB1Q93xjBtq20LDx5BvRFOYECjo1lRVDRgAUHLwKxaNkZ+X4iPFff2KyvDp0ZWZe
oCIWnM4fqLu0KmRdo8tFcb1sk9oVF7dkHvBiX18t3cWF0F9QrzCzaMGLX9Kc40SF
zXDjeZxEMjhdXh1vkpU1Ve/2tX9GZ0+WjGsEzh+iPo5/LoM1ilZfUtgLwc84nRJN
LCtQ8blIjMntDVTGXlHmMJKK8FX3+T83mK2cTlWYXpe7maJcaHXo4AvKx+chs1cP
Ygoh83oVV3YmTaX9cQuisH5EekC1NLuG06fx9FgT5lWpTBGjwQvVsCBjYW+1Ohdb
uJ/o8lBSsN+rRgikvdxefyw160In3VozYOEyKwKoZA/7FcW3K9Uu+dCH9XSMsK+p
YQmGyyOTlSR1mew2C2e8dQr0CQQFdVCiDXh2T12IYpSFU1u+D9tiQwFVMwh3YCOv
IY4LqZFk/mTqOiexb3GUVRfhp8SBfBuzEOiNTUIDW6J1AQX7c/3f9YWk+HLqbM4B
p1pgqJF/AGe3n8dqnG8i32NjTFEBCZtpI0ImvnuYannQhs34ZRk6SdaT42Sj3UAq
okMmbQbSnQ5QLdt4B5vBn6HJVq4BmCmyhnNqY/jyFQ8n4It4ln3GoUswjJWKHEd3
uFFjVqKBvJ6NMcREQJzMKAxt6twEiia6vjhW81PWONIJizA9baaFqxtBCXxS85+c
5aGDEs+G7RxstlYNtb1i7jUxFRi9KNLiPcyYh02E/lAXgdQWlxSG15QEKMvppbUC
BeMqqvPPSEXSU7zISqHFRRH7YLLbQPbFLgtGIIFqQXhedSpdvh4CDBBKt5/BNdTC
9QiM6qFEdD4EH7EWIB8E/E7vtbWZXSLnFubJWshZCVcjh7JYo7Va0umAyBAHq+2e
dga1JMRVRb9zZ9oSoTlpBxdw8zS3HNkrhR/SRVdNy+Z15A2pxvfHt7w4Cj5pnVYi
OvfSnMoe2F97LtPmsQTeKT3IUj8EquIOYnRh/5tsOKj0KS7aWGkl0K0w1S+Gw/Dw
pPuZyEtL6VtdM9Cbaoi2ZCPkqmIzTFFLysZVu9OKMbfU41YdfIagdSnrastK2sDl
E07Baa0izqcR6wkL6kQRnfcBzFUVsie2W1cT8ed8LVbz2lBNpCP8AzyGITdioViF
8BoD1VEzpgaW/7fe5mZN9bxULEX5nyDSMXXmsmr9OF6eSUZklQN1ekKBoXxKDe8e
0dVJxHtd7Z257SSSO43vkESbNUtwBqBMNhwwhXKsboCnDB3bsZ2Qt98tlS5RVpRG
dbl6RUAa+UKYBV4fVt0by8N+Wr5vgQk8JpPOORop14yvjee701vzOqrZlgFimR8k
6kiVZZGM7lzKGxGglLqXnDGCxl6d4w6tJId7B5PbhzVLVzhfBufOlGxyY+lsuWqo
beQf1qrxq7Mr5GXPdh9H33W5S77cwcHcYeOoTPxuVLWwMRB+4Xt3niMqX/Pz07og
kUoqcaG6Kcc+4/6Xa+r/KA82kI4lEDAT+gs9FN8kB9MYkiTvbkMKm3J2C+8/tAUL
zIWTddK/eWX6e2RWfD37MNrsNhzapsUtswbZXlE4GcAR+x6Mge/F6I6bi5ES/uEn
uT9EuK52Hls/IMaD1G3Q8nxhgRJ35r82ZWCdEGtWFIHtGIMdGvss4ELiUvtjwBPj
+AFWJbTNMSwm90gDZ1lrjP3RYCCi7+Dltdlf6wW3Mr3ktVByg5U94nfGPMtYQW7F

`pragma protect end_protected
