// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Qg2VcyI6PEbDctq1pu47SO4OwOk2w4eEQceG5LKCB+dDaSPxCbSXG9ok4Ecg
uca6r4YAO0vVkbJPLtTJH5UUk62L8Pz/F3h+FTrqIom4QhXHNwSOGtUq/JNv
YRlNi/Jld9bH/KYRFFYGfBB24M3t3K48/YP1ovSi1pLnm+jwBRLVyu6LQh5B
YtBZzs+tL//DpBhT9Ry1xnf8KOfGPtfq2mFMzzmTNi7C8lRU5AeuQMI1tsal
d4UwL4YegkXT+w3dfkrjDv26j/yR7UJFRo1QmS9z9fLSVbz/zFrl4agq9TzA
2EKo3MTj8AYhzwjDgVmQmajrtgMd/C4Ow58VwUz1Vw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
CB7SgdkbtwdcWlgsR0ZQA1qp1aBNjdh/Vdu1TLn6fVQaRQXpyWjxhhpaD3GS
HU1iD/GqClbrl8NzPro7uw10mJyFPsfSMkIm0KzNx6dVqMOHmHMp8F0aQxhI
MuASZHpoFq8NiBR6LSwSFH6b67POQCT9XX987As9TyW+YccxXxBxngnpgqP4
T4t3jQ+KEP/L56rp3w4HeQ9JzJudnLNdBlp795t9vUKcCjsfy4h+0BFX0YYd
cEFNYW6LrHxoFh0Q8SrBzOhvtn0dkkeJEsyfCXFhvZPkVpoOVfzRDWhVoLYC
Onqx/1lP81plgmhpa/CuwA5/0Hj9AWd1BPQt9lGiow==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KxY2lvIrHloOAo4yTS3+SAP1L3/01Y1h3nPvvaolUrwxGOJYGQ9OdQF8SuP0
v0fWOQknEB6efhsupSfBX5P1Mdd91F8vFa2oWwHsGwYfducrIb8qdp5qoXTZ
BLMOxIdo/RWbEQ8jks+6BhVlTgBS8AlPAo7seqIv0QFiXbf5U7LUbJTSF0NW
CoQy7sNQMDFgwblIxI5LX/QfCKSmAaZ+pvJTRlrOd71CX7njnEEtSyuCXt/Z
cu4hYuzg4dgTl2ZThs3m6s6ElDyWke5rQemAiacdBIEgml2k4zhSOEbBfQoi
ZdsFRgiYul/bahgEWKz48KyAE9JvNTtdeYWjuqAA9g==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ZSXCItVbc3h2uKX1xaxBOYaGSBC4SWHfsA61OHHtbMOob7GVIsznGoUUhdsN
Dx3f36p/X9CzwWhGm/+p8Jmqpf6CleB4F2/BlhrIDkj4pvR1Ia/8vgB3XYQX
HsKkekoolIyeuGfQhmUeD+/UjC27v2/7KpOV8Zbf87RooO/3eVo=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
XBPhN5cQao7h0xAvrMrYl5Ba638B99Dyfr8LwBKmRIR/ftKl/Re7/BOTnZ5F
BymR7l0YRXJ9TC9H3U2rBf1QSjhssdABUv7/n2ggOoNuJ0W8flz+CiRs6EKR
wh8FvOLGoZ7gOxmFdbnNFhL1Zw7lvYkQ/oW0VcQkgZ2V31hD5PMt1UCxm0Y6
z1vevq6fFrpY034bgDGLoDEBA5kFpo5IFq8+SpIJokoCFPDyBTBxreDtl/aT
dGlucubx6WGHHYvwfqUr3LDCgqFsQYOZvZrvRS5130fHISWLtlYnunara4xy
7D9CeaLSYRt8aSRQ4n6ogVhMNVu+u0wUMYG+tIRl3Uu2qmCkrwquD6bB799U
aRw1bHQBqzU2awbXlaW/TkT2PYaFbBo53DfOxfz49YoF03d6rwKMxL24I+6R
/CSgdM12iteP3MCmKNVSbeyRuQuxrympUpsMR4jUox/ridecv/ypkil1e9uE
XHw5VOhJe/RSr7KtvsLDoyHxNcsCkpuy


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
iszsuSYiio+04qsH59Iiizs25LxtKmp97eES82/SoVCecJ4DaUjX6jQ/TzF2
QeS1jjgnxSlfPljHXlYLRZTPbZ+q3r9NgN26YQzGYB5CQoRG1/gdJq36eBdi
EmUKiOx0q5oh6PArUsLzFGqqE+ItdEQ309+QgJqVX0i1eWSzFpI=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
p8+gc70z8Twoe/yJxhRXyeO2+eTMzAPrD9yzTPiMJ9uH58nmI/doGQYdCMdG
zDpTI8n1auS998Ge5gW35fED8pJDzv21UWB/ihmXa/teEtEn+FaEKn0QUnTv
CeAn0eGqHIQoNKCRJU4iDqrgqSQnKN5D1fV65bxab5Wwy+rK+pQ=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 93744)
`pragma protect data_block
HM40wu7LQuSuMXZ/vahhZ4PJW+Bp7cuBTyLwj1jwQnv5U4Xm6Qelk+v4HvBF
7eXCoTHCkw6sKbnfMHrgROZ6ZcFxU3+SeuE0JJ6pDX27KO1+IVomEfSf9t63
onJXYtMW8wH6egAx7B2wKmDQBfluclycBW898ZcK8vC1jYWf3Udt4INelRE7
vAsa5+meHzk2yTRzNKOuT+eJ7r9geuFqRrSVV4S6l5DNPZwrzNC0M4T66ism
VjMosO/qvieA2SIqyDBmo27k3L3EpJppIAneKiUijRYYCX8dwkCUwYyN/Cz6
bovtPMe/Y9jzgJ41IE0HqFp3IQ94dnKIw2Rexzw5beWkzi58AnkuXtWpUjlW
B4kdlIC7xnoa4R7sJymFsQNcNBbxLwQLwPpcOIdkw7W8mX4uwINh8hr0vv+0
WXVfbH4TqOVXtItIUltOZMuUg1M+JrzjVlhmFeh9+/8jS0ZySz00bWwlmUqG
XsabioFovdQTMb24L4AmF1fw/gwmJ/pngPeZ7UtMCngkQUiQhG8SgGMml9y6
Zf8P42763sH87i6pt1nevYE4Y3QaTIrJc7qW9yncXNyyiBDL9PVF9/VsJjUQ
bWaIxIpoIb/ldGL7Gl7IHKlEPAxCFl4KBGsMsLaF/IxzlMm3e0mHX7bTVmpj
5+leFp8h8r+AumZpvxVWxSIRNM9f3zvnrKILq3494IakElFRpUNyxvRvZfby
97sHfsHkjMnyGR7Hgzy1JyoAnrBrgfo/GkPllXcCVYSmIMgg5htff+PAHtg2
XHq/O49LPJo7n6D4LPO0BcNs0HQoE4s8u5CQB1WGnnJESBPrX6LNEuGXhu2+
R8pWEVC19uBFimewP3GKYDRqJY7kpxrQ1ZmkikdYQxEVPZpTSeT4qF/LxOPq
BLcYuE5O2yOkWh5upJbpcKGEiYw+diV8O9eYS6PF9MsqrNO4duG2kLefrpyR
QWVRYUw/HQTnwpgQO1fQQLNt+4CX4e4jPpLvRsb0cUIPxfeGdXpVJo+72pO0
vyvDvWnKGYHYumPkOR9pKBbYBE1kLRMXugAlN5Odm5z58vfWWzxUg0EUaOTR
IcTbIYTtwPj2vKVbPk6vk+TKIkCRgyqo3sTcOmdjAbVdW8WkpRhEVNUR35Ad
5P4PR0eVBsTR2PwXVwQO0atWQHLTATi0YF3AEXg0BdBhKMRVI9CfoyEgzs0a
Iv7BTx62cEi1SRqNELPZhv1aFBia/wNYTSJZiI6d7aOjgyZqBZr+U/1pTu8S
xYJYeqpldi2b/HuWE8TxunBsxenPRl3sOdGhpcC3A/RJOfuc8/loRU0UkuR9
xk7WKTnqBcACZ9KOT0L5nkjX+FQqpTczGoWbzudY3Rvrqe+d6i+SQtapsnsA
EihAScekropWv7Fx9O7InaRYEky7sKFDfRWF/3kJO1AVbCglOaffWC+9C9i9
Q3cdeLo1rz+yacHilVu+711td+w2z1cizsrWUJf/fWQw0WdLIc5pEvHgNhPn
3VgglHQ/cSL0t2QbaPUCmzdP/y2tLddbLQwZZ9FJlg2nLkFjxruvz5LbTGep
xbde9PuEtCOhV4LDilmGxUqVirwj7vOpZZUlrCZBRmHXL5B7FA3o1fz8PN7Y
47bgas9ncKFUCTeCGF72Y7O6A+1m70E9ZZXjViz8tulIXWLUm/FNw4EII97u
mtge2g0hDN8WP+G1sfJEVuVQmXHxBroPxb5rEPVD6g6cb4tsjqP8eVNUUbbz
r/r0hBdoB5er8wMyXSs68IxqvSmGU2blzNranKltYSadMhxS7EbpniTSxemU
A9ShiE08ukT8OE5ODh1YE562UDU6V/P3mmkVe7o4bkBs1NffBjw0JzQ64uz4
kZ2TwS1RlgWdlVfZ/fk3T0PD1k7IH8k/5QUTcLIbTCLH6s6wIAzMkrX11zUI
x/D8A5Lh2Ygg2mxNs7lDduVppLMPdpXAvK0sYC/2P8j8QuI1a/extMyH9XJ5
1bfuUwmdchBwtQdMOiBNE0xQIA+M6/WAzc7e5Csda0YyF2S8X0ixDc+P7xz0
5lhA/kGwKRTBjW1VnTLQvr+2Jhcl7Pl1VsHJ1EWt/CNdanQG8xGFvjSBW4A7
wHz/Xpwlrsf7VmkO6U6uMIE8QbXfgGa7o5rdaQ03tzAkPwkdCbhWLheto7Pc
0OFM1/DeZHlBJ0JthjeuQ99RG7gvjWpmXd5OoaBhHm7nRw7WszfTBrmVko01
KSTdPTM0knKNPpztpXlbwn06rGcd8ldYGCIX8jrvjiLJYdbG4YtuMqD3vI1G
JD4q0skifR41KWvVmg3THstTbhMUjnfoxXABWTQoVFQdwZLBtnMF9Y4xHk3O
njWGhfWg3+XR2PU6FDOucoQP3/pZP3rn9z6JJnHarq25lWEg4dUeS5Ctm61V
1lZBnMLpV2RV7GI+qQLYP1JaSFwpapAL48mE9GBPi3kwdY8HluV7aqZMC/Xi
WX5gdThmPy/hTieHnriuqvSAd4/sJ6A1k7tw8AQJo9nn7XqwrEB/IgyGQ3OA
q8p+EX4hu7N9XXpLJ032i74neC/Qi/ES8eU7KNdomsMmquzc6R+bf44WwgcB
X7muCd79BVkPGiUyXFKYh4pQcQ9MRXby3VIUpRPsIRS9dF6RrYznEbglymf4
9Zbu/HtAhE9NUOWGlk+FwFCZJPolfVoV3YreuSukWnEiMlC8MAZSojJ+eQ9F
C19e2LxugSFuV/PsSZLcy+SzeHOB6dpCnrl+5Yp1oR599w8jNIpbBsJ6w5aq
B7DNU3Raaeh9afwUP3XkZQqrk4yN5moSgy8DTdC+BA38V9TCEUTuDQI3kzjD
SpS5bOXqARnN0urxM3HJYm47aIgSwC+mPqj3rlaxkSGx/HSA30ySA/46H/hE
hCU/JdcLhW+5fCSpspmfZOuWMjIq01FR45uxX13aYdqEVNddTQk8lqsaJ1q7
t7muwak5/GlUNLLAqowv+NAJh9OBJZXSfQwrZMEDjCgrF++J/5vwRgU+3ta9
3RgqmaWRRWq4elBBbkn+62n18eX2rhVisLcoIUmNw23S16FHAJokMnb7I6Nk
h0ChUGD7FICTeHpJ9UKRzeHOguj7JO09tFI9bSLQeWgHGzj0cdEMUGnTKMi1
ZZRcVSNk+XTXQbG98yB5oSVqgBjp52JA1UeaCOSxf8TfxhsMYU5ijjrjSx+r
LXwf0g7ghfBi7nx16FQqSBa9ihDxPkTOTnJnL155CI+rN74XbmYqdH5pdwVD
KHuZeIipLQOI3ulpLRScxzsE3ZhrvfND8hmxA+sul656IFFZdtP88zEXpvgF
aaWzMne6lDkP+3SjxrKJSad/Uk5OCVMhgYWVej4/e6N8tBtl9ILSifufuy2y
RspRCNpEgk7A6aR7yoS4f7nm+E71pzElATsN0hBm9P2loga6dyjqsCl1Ulmi
Rj0dn+FKnA3H818HYK/XtGoFQoi9YQWYnVsn/717tj9OvHXu+bx68SOIdln6
hoHrZ3cmv1vxCftQMVI+gEAi/Qz22WZ1bE4IJoudn4W7pRhErq1oQG0XibsG
OiPat2ucQzcC6RFZ3TtVa5fejfzVSCPVUmv8dRky+68lR1xq5XGWMQFv186+
sIIWQw9wTM8AW8FlqKnKJ1OGJXArOztarQt5X8srrz5JSwdWcX58azRb05Uf
4NdwUNsxcd9JraiJyDgHQ80EzIUIKg0pjJXKOlVyO4R4yZTD679BIcnZyK0L
OP14gl0DzNswIbGQ9veQZzGQH0StTfkN+jsh0J3CcAsRh2buXUPBFDOW7CVz
yFP+ESP+97n86Yd9Waq6Fjp5obQk3UKsp72/lnPyPLJp6PAvtbeleGCoOyQ2
jsy+bpzcRlx1EO4h4SEQVVMW/EhQO7vMxj/LwFGMs+1Mn1LSeaedjC23D2lu
36IZQbz6BL+i7HOWVMMEalL49NCqZp34mDq/GNbU7m8FBL/0xCfa/C3EmuCt
V7tGsR1o5qkOvVYzR7V5kB9EhPz1uDj7CjhsssAh1icrW8APwMZ7GgD9Q0wY
kyh1H39WC+VA8GAcpEJPIWe+qGE2n+4USu8+LfeuLZnNkSGoK3lLstnLGSvs
yr4CwE/i85fB5yucizYZAlLLo+6eLjgv1IBWWBYFOQYbFC32iHv6kTL3ArzH
36WCQcZAeYCHpYS7W3ud0/AZr0dvLIylyYqtp8j309CH3SltPiRp9cAG1USZ
PkQfVklAIS1NTAPmuzrES3jeLUcktx70Oxu89PWAw32zmXZ4Phnj6mD8M/OK
uY9fRUvJdgL7kWtzzPLjivY1syhThUoru2ZsXEHo679dUHkrtP1/GZgZLtQW
JwjN7PNJfPffG+A672oy4tfmluMWLe4rqEXCL5IY1qr5qnQUEg6va4D0S+fI
kP1GME38PabXG2hZp3MvJbXtKb06vOgH8gLnvy8t/kf/FZk7fbNrzNAAxh6M
dSrUVOIqx3tJERMUgN7cAAa95F1IbSedWCaNl8TfERwtfghjhPfQU+l8owSL
9aADQJ2af+PSZmlInMZT0I3JsrhjKtMWj+5MJHqLq0qazvMhFp1YNCvKjLux
WwRSgAka1onO+p4t+llUDhaNW5vexouylbeSvHmKJsx83mhDlgvDQbbizYii
vTX+RmsQi5ocvduysy7eoqzbLWspt0A07AQLAMBWABx9FIA70TqhXTYdgvYW
eeYEgHAkCF+nxQEXO2qYxhmXIBSseC4nkdOPsrEhArj6bSXAcW6uUs248gRY
vsM8tXTHH/zn/WSdqTNEiqoCzgjQxlSTkEhSBSDmn/MDfF9sOX0Ep/phjsS2
9pk7XwWH45wBi11tSqnPvfM2uvtqIhxeubv86mQvlgSI4IyrZEbFoykJ7Yvg
tTmpxGF3qXl8ff9SbROxpp/IF91K3ENk602MHWlqSDwRwAx4N4OpuIg7JNbg
8XXSaeT7brbQUQhI5QdkVH00SwGgVkzUMKaqZ98+fBh0AQOU+qQ1UgLeM3k2
8Deqa6r6nlsVrgS8/HWsqxyxaxB8sH2OlK8VGwcVGu6LMwKbf5V4UF3yfWFA
f3dmFaB9bmMc/tELffKWiT/pPVMyjWw2RHYA/B4LiEvUfcG8yQ/99Cd9dc69
ruuxTmoV2KZyibihAHoo+H86kh7R4StUqn8+3J+cGYOZxUJecZfmPeZsPs1d
J7s+PBwAOSNo95HdJ5rzbj4Ga1AOwiAfEU3yIVfFfzhC7J4wx1rEnvz31caF
iArxu0RFhb6umrs7idq4gny8IIsvtIf7HyjuUAPoEYSdxOVFU6cS62k1V4L8
wE+ARI5NuNMjjJxsT34WKZmSazjj9eWcPL+u30/yU9yWDIx7abzfaIv2JVOM
PPah0AV2dwO4W95ww2+RrjLHGpn9vGezd31pfyHVy9XIr9JLHbrilv6M8zr4
fGM3GG3G36TNqv0+nkm7GXpzgW8LrGHt1wbbGzOpbiNOmWYvQ2lm36Oht6tF
T/aqm4ebRYZFrp25WjcITCNwFCaCojPjF+CF3mSyFLyvPOhSNRI+Ff/eS3o9
qneb3jND9mXf7hJiNUaJqxJNIgb4cVJvsOnQNSuapnStQRcEG6AkyQ2b8mz7
3uXL3lRyaEC/BDAmpSs6yFfrxZoz4NZQxqomPTJRsOs79TrNhdRBqvqSG21e
OVC1DSp8T79Qm6ftVRDgyL2DtTD/AXZ/GbbI5wu3Rtr/Q+yL0Qjsv5Ad4CMA
Usjjuh3P7+TloKBmwk4QLAktNg+0lJNNMfaiyhgcOzlL5ZXB7OImNHFKruel
QWkXha2qgpFtmanJA2pJDpOO66bbaVWkqP3VDMvrjs2/lEfYrsibpvfSwXN7
N4BK83xGj64BfxXpCL8tDahQnea8eD4vJKi8ao7sxJ1YPOxS3QOmlKDe0FTm
yMwYXHMqGIVCnbuwUTGXHFesbPdx0iXLJM4uj/dsselvLHVs9YLKgNOiQytY
u7Zt1Jk5C5VS+El875Uq0e9I/mSJQsejafDg9w6EAqjdOLM5oFFqqDCNKm/3
uLx2tFwAjOyQJ58Tw/BDmCYtdmKTAlIlrnpO7fBaSYyyX/qYXZtWVdEX0U9b
wGGM7xVJtb1TFaXEIaHpypAnV2/+E3ZVcgv99O0l87f8hXUfs4PtqgKqeg0v
juzpx1ico0I2cnXg4wq4eAbHrZh/59I0b01P83w7cRR8uQabWJrEOeSVhPFh
oavs8zxSJSXrHJzfOkv+NFQ2aZE0xjZp5jn2rV9bKjAsQcJTZ9zXME9TN1tY
TTS2Flcg8ZmUNgm9sBdhxHnn13OY5sqwkMSqDYjj2nllpJSBKXwylqxjH2T7
2xapn2DVVUWjPoaGcJkYUQZP0xyU0CBUfYalHhDfW8/aT59ez2wEzyyxGtT5
/b+zw4XT8WzYiB01WKvdCfdd1Dp8uqA6n/fooLciG0qSmbaGT7fm3yG6Mo6+
8cQP8tTb0tEfkeP6IWfHA6JEQsRvBv5T0BzDHGwX+E893VgylDEZ1tHrUvD4
tDLulVoorfA2l1flTCgvD+9TOa9HrCyA357MGxrDBIhKfVxHJPHRXrMy5zzK
fbQ6w5DeG8BO2OPFqRQF8bK2fYlrXelFORfTFvTYD0wnidMxhbWWJH7Ao5Sf
HRDnukJHjAmp48zAcrIOh/DCkCLwd52UUDeuKjt81DYMgXraFzaD4tnbYYxm
V97FFRHmurvtpizIYOcGwNsRe7DDQwfKRMexm6c5uXaKG6S2W6jMyEI8zEJu
k6v+dAESqKVycl8wOtcntX7gny+p/HPov7zOtO0Yw3FKqvsapvHtDHqgjoBv
U2To72rUx+63d631R/xz7xwlyircv2ImvuWGOlg1C0fH55wRBz6VV5kJoyQL
/FEKw+WZ6GnvPw+epYtiAkJ8ZEOPJ4MxNSZrcAItvpJXqY2CyHjT1gotbasQ
nZA2wT1P08d2AUl/T7uAVqy5//q1zrYyoMRLvOyulhq2CCvHLIHJrmR95aXz
1GhuKgqXHIZv0bA3O+cB7SV+BBNhKVdQNSKBTgyYKI/9ZW/YJ8AYgAvmvxEy
S/KdxBx+zpEaimBGcoKKiRiCK1H1e+K0x8sHtMyZKzg0B+KGQRqg830RM3pF
zfOTZya8xocGUrVz/q3fOpeu63lJJfgjE9ekROQnNyt8BTWLhbmVKC8VOhvM
8dZe5Dq7ZoXA4NbyecidQucaCwg8Jb5DdjG+wH8Ha6+5LeC5yO/NsKaTfAIF
MCpwNT3JCI7CefOB3TnZAYK1awb63LLWVnuLaDB8cO4vOEu+2gTIeYjriqY5
PjVpeoS+AmeYGQy0uHJ21Yxvug1+whkR+iMzCsPowLc235+RLvmTm96zRAra
TXZDIvKWy3VlUMpismdGTqLqe0WTV5oLnLzybolVIvVVwNsGvFSkGfbKEQey
83Jfs9TsVY6GN80lqfF2Fwh7eic3yEk19hCEHFByaNsjHSrPzs6lz3JTXhLU
p3QtatfnhnWhCpz2KQdKacoDXRv5BxIKmiy+Sa6ODKJU8hRdx/9aihBY83th
JgF+cGT0kXd6oz3x/xTscSHPnLKGEAWR/n/QVbtMuCyCT+YIf/Z2kxu/Lijb
IjsqfRXRPrTYX4a5RDFgRNo75umnZ1FZFStsh4Bq4q/GEKsPocj5N/cQKYjk
Lra9T3EP4xPoXv6LJU8buSMS2zarjMB783jcWfjeC8sH4AS5mQ9xZQyoE7X8
PrIfwaQAIvyesrWBvbb25gHqmOdzDJcgkOZyFoahZ7E1tnGTNzd7SF7jb+9q
bL8FX4A3jNuokVIDvJmXRGXICJxBX+N+q4kn0B4j3tW0BVDUil3U6S3Y4CNJ
EKGTVZ7mmPvyMi0uQIVC383qzM6cYrLYiTLdFht2lIXWJodrlAmonOvpRVoQ
TzxXSwjD+r0UOV7Gp6wslsGzBDiXmGsueEPVIMkMfHXqvHvi9B4XRZtUmPQa
g9nDmVew4X/JuVUr6D0MhVxd0G5Nn8VGOuz59vPGURgSgWBFlC0i1jUNa8HX
e+dTWqPIAUmxBs1BIQWbS8ghDTkHVI+BZgpyO/pelP28YVP0jne2qtochsym
clOlkT5YWMl26aWlmd+kgMHAKopSGw/NlDZlJ/MdhcJWCw1rHdgpoEs0AZpk
i5AkLEK0veJpBKaqV5cu56DPEkLA6lRd7bSCNa172i8hPqYf2yEFtB3CY67r
dZZ9MQfZlDMh3Cb4kwV4ZF1rPP9s/vspzz6VsFjgtCvlD/WDgupp6NNgiElo
zDe8optqtFnb3chkTnlHuVGRY1Q1bSez2IPtZdOk8Pezl1YN8r7uEp7phmQ3
i9MPQZaKzcSFCJmhPn8neHiHrzXpjZahMpNa2G9uzlA17CLuJaX4Z3x05OAE
IyO8uS2GBoxWzsiOqFdeACJ8nMb01xkTkx5Q+tlG3lcKmSiuAPNoIi9J5zpc
4s5/+gtGVWRb+AZslwI9VY+Za9U0Q3d9EMdmWqkbnZIBmlb4gHb/hTqMQtR4
Uloj5gnliZBX3q1+xqqwJUrckZDGSmm9vLeGxctbGJrdfeaciBbn/1Wlx0ac
VsMl9TuDg+vh6ZtWuH1ZowLAr1oLHHOQkVXvJmqpZ7qzqDst2dVcueT87z+O
DaQj9BPX8ec7ntJn0LP3gfGGVd2SlNGYBYmuBBYVAjxCf0eaM7eOpHb89M20
EC/cTCw9TKv/HOd0NRamn7SjYe9XNOADUOBSguRy64oHFZPNMVJkN3/AZ5/E
Ra2lfGWTz+MJjhl1Ek2/stEKfb+7r0USUBsNdlmi4ttFWIt2rVrakY6jC6n6
vBeFOHegrdJZDyNAqWlkHBG54sY5Dww+kRvWuYcIATO7Lx39nXP722eTm+h0
neTo9fE5TohtlIyyKHsf+D5Svfk9lG0heUoe1GkeXo/puDk0BSH2ZyOrrDAm
qJdnfhFKXVcMDT83ibK52XU9n738+9WYcKfyA97wa5OWJpvFFpoaHjirLRp7
MlkTJAImGQsEe09Xdkc/QACf3TNbTWORXkyUGXMrxJiCy/hZ0ggs4rKIpeR5
cXb9sUHkVrRRRrh5qEbRz1i9CUXPl1S9rLegr39Xh6OMcs9qqq4hCCiNGDiy
KZsPrlL9wZ12Hr9SsgUKPXSf9pI1HF3FtazUfp9QlF3ef6VfYvuxzuVJEV1i
rEIugCbYkYU0xe5Dq9anQpnrLNWZprTw6XkMvlxJA1p/8/wZzBcAw3qHcjbl
B7iC5xJmNFsdaX3R1JmF8MHWZ5kS328KhaEhFKPTJ8v9UFKpvRR8cTqLyRJ3
njxUlZhFHiHs3ibtHgzCN+q1VDRq2QEpbbnvsqv0PjeX6l8izVPOYK94ARPf
p74olc56511ZIrXYPUP1GzpIvCaVenenkLNNXxwiV3HxiddG+YoTYHQj0zyo
OEeqzgSfNIsYbej5dhKXuMtxyYxTdyYFjEjd0PIzr5hOBO64K8gvgMryFhkw
z1VgVd3KI0yPakfdMEdPvhi7eB0aI7coCL0t2pHbFJBaBJLE99yLJ/AU7j1/
YAkC/WEoscHrps0Gu16azyuAF4+x3+C09YLyPaJTNCjERr8IP9q7oxXdO5XG
OqQbl1Ghm/lN9cCly2Pr9SbpQulIlaK+dSUzszWXJhVNMlRqNwxlbHOrkSWI
DuvGdy0E6EklpdJjcjDpNrSECgS8ud4UFM/zehx4BG8jPKPPr3rMffFFac1s
vzWSGByllnAEwp+s9/3WBSioiLvqbHvECz5jcS/LMbtLoCtHE+3kHSNjaiMG
X0enBN/ReSsINn4CI3Xf4F5IQYpB7ZgVG1Ln7JAggVx6T6KKCI68K5uQpF2l
r4JtCQgPwktey6CCkD1WuhEtgxZ0G9E5PoRVXvZxIEJlJnMLdgCAadvrc+zi
sTQE5HwghiOC7s8VQnjGBESXG72lcNE56dYNMdco919fBxiI1XyQoxNNc3+P
Gmeucuuz8j9hCuL0VPlGrRg7IG63OQolD/aZWv7Y7y+ba5B2noQPVcYUu+jo
Lcs5mi4z5BZtBExlX/hfpcGjKPwAqBkUmW4x5DIt/FHdC9e8aAngD9XAMBa0
tFUjUkuQ0G2/cNvVcwpw1Tc1pIBxwuYU64TKdI9SsZ82uLGAeVdVjC14uLI8
8SgoBUOpLFs+34y1bkPwvdlK4+BeGK2SWouIDLE+BtbVeeqVBmozrQNPjrjb
nj7W+rRNol16Caafp/4V4iKZNR4fmork/QLuI3iCJXD8mXP6GXnRlMbZRN70
qyuS5zKCcIUIHcZAp6vQMh7PLm6o4OLmsvzM7/U5s5PhCmEjfOXNPaEYnQSz
l/CkHoZ8KqPsKuvJuR6EbZlLZK0rCnf9qkgErhY0vPgelfw80WrrDBkylzdU
D3PxPMVMrMziF7OE4r7K+tUdI2hNjCTU3v08WOzbs34WuY55K4w5unqKZRqS
cJnaDEpnLQqg5NI8WSqkOCvaBqa+nUlaZ7OrN+Ig2B1CZNJXtbg6F3YmA0zF
i4yOIKeswLTdqfQzc+dwlfq6tLBptm+RRtw4QiBxO1LvocWLNKtQiIK1Yagj
N0HxdNyn56UPnX7WX1n85zn2mgWH3o9WQqmhWsc9kjH9RrXDZ1CbJKjq8V+l
pIZbD/mtiKRo4/TYxOYuK17fDJSsNDKn0vQVVbfgSU+m980zYQeBMudqfhj7
Zm+BAky745IX2WZ0xH6u828uWENLl/29Y9P+2nvw70AoLYZAhQA/Cun2NPrh
M/snCarDXCda9c9F6SeBZg58xgsu5JDiZgrIpdEDFplKtN4H+lOpEq5X52U6
12NwkrQRRvb3zERRFKgToG6k124uHGeh6bB+eAruLI8f0x0lpgqHFuQ/iq1R
gMD3Fg/9Dh/s1rmVW1QAMgRt48Gnfqadjm2C4YBVmI+cLzGMchBSXjM0y9uT
ww6J1LW37uQycNhgZ0YZkzAthvOy5cU10AsW1pCNtCstzXR/R8XhM1a+QxWw
zvXH7BERBN+OdOrr9tGwMcIdzFKIuEFa22Tw6cZ8KwOV4Ya4WTQeP/xzIoT0
9yuqJ5m4FcZNLbnB8w77EjQj5FZK0gll79ACsiaDQmzsegMVob0KAMH8DyFL
ybG+aPUXcY1vW9m6fBqzxrK/b/y26OTArxK4i9oPjbGjoOdJISNXb1UVyZn7
oikCrSWs+cq2m39delHACFUKxwzyFR1mqk/qikaKkp2f13iCVZLyIv99Kkl2
hAI9X4ZTkgfmm9hVg+nBFdzpvm4bHhmi6CKMqzs2cS6hMNhevMRQp4hnizMr
CT+Hoxe5YPWfzjvQdVwuNIrWzvqUrfNXPPYcJMG1EYILlt+QN6XSgutXhnXJ
yDaLOe0pVHcceYt6eOjwTXPF1jFPgsib1u8IGSS9wd1kAoKCF4sETCU7yG4P
6fpK5rGCACmSJHv9n3wz1JhG2a4iwIjdVNZEQQRXP/xAp0+9UxJr/A+EeeG5
B7UxTGP1Apg6ivS0spDXEN9/bnww+BPm5wgWa5HM3Hwui2nP7As33Mxt+Jgo
7Zxu+9Tlk3zMPPsJum9c0ILZxJZ0sLuncmB1mhWHbk9LQxovXmSpiNS491oq
naCsHEfpu44KhT2nJ2Ze8maAZZOsIbJXNiJ1/IdhRW1/lXjhoSTZIgZOXVqV
MWTNhY9/wItsaOMd0L2nYRNCdXiDf4bCzb2u7+uwyf+MWwZjLubT05lrN9wI
LsX/3dd9VI4jG97BNeBSQ4spN0bZ+5sc7q5I3XWEKAibCKg1SX2HCLwIWNkP
BhzIyoRZQeljHRjW25IDb4bQ0vX4m4DgtEeVq0eJ5e7Y6AhzWnbu4u5IK+Yu
c2SqcuL+lW5jClgm9P3aD8GEQxmH44i0E9/g27o8RxmfSoAGZd7UoahPwXM2
ZPKfrXN9Erwsfe38+ASuPpLjLsS3mqcwU54aMcnOeY4gZFsBimVeRvksYM7u
SEkHG3r89UmPLwKVrhBFYr9pwG/hqUx64bR66OCCUgMWcC34goBhvHPhho7p
8rPFp3eKik/Kowk/L++1NHZtd5fETa12CrSn7f2uYW3SwzROhdiVqQe1xp4L
ZjS++aE541+aql9vhq5C4oL2WZvYq8GHZqH0mvGh8HTRSXH+fp9IkVVhE51c
EQ4bcVECt1vspLWJB5azs41LJAkdWtJ7yt09uorbzk1lQ1LUBcLd+XVsHoZ9
jLPAXXUi4q4q+RvYSAoooyYh/r9KRRh8QcAjCPZGgLxl8Z5m3jfAuBFfZLgu
fKQXVCl50YeNKdlzLU2sC4Eqd8gqZF3BU/BB+aZLfVavh+B/Uxm5Gdbd+f9k
An3iNSR86wMjeAtJCghGFF1+Z0e3VFTxOp70Iey3iiS/9tGI6ToH3zXzuMXD
aVotvkcXki0NSY0jC29Y4+NvqzUch44g07gMu+fCP03ABR1jSvojJ6O/qVdE
0GIobRfOYsfGyWi2XTug/SJiXWu/ikY2zR3FHA6CkTjGDK85aVEo7/2k8aje
TMrM2/LAVNC+WWo/5dbCG0LaG2yGCqLhYJON5pnLVJH93c9Xn9vckNGBpiHH
BkIBf43pPKjmvDou4x5JusRTK8+5NqWdlIR75tCDZuf2uiKX7PLswcn8iyO9
XWAUqB/bYf/z1KDvUmP57rIVeAQfMQsko3TTAxJz6JXr+JMpGEn6fkdruMVT
7cCVCuyEwTL9SUCGxXcsO54uzhIeWkglRazszvfbeJ+YKnguunUkUtOT4/zp
6R2yu2wI29kIKSQ2Ca7PbON3x/IeRMKErd8m2qSKFcWQaAkKI0O4a7M7s3N+
wPOmXj63LdplnPTDdNhKS2k7i3laD7XOR4ULKIE5gkGoGg6Z3P5Ourt2CcB/
NJI/H2TE3p6FN6uVPRlTmlT4mpPJJD0vqpwojuGuhJeU0TMFDMqI5A8BD5Mc
gwdRXyYmnhFCviqZcpCTiqAx70s60Jiq7zEJ5HX3OPpNQopO5lw4J+imIYtb
geW9k/XV1DKH4HFIRXG6YjFVW3mjszJi0fNT81GGDqCXTyHw2XsksCs6b+Fv
cNKv+MU0oIb2tcOxZo7+rYKUcmu3EpaQLuoxWpPnsJs9CAU3NYIXk6nXqfMU
dO18uKh1cZ/iqXpbxmx1vI3Day1DZkFaHwM3hh2SAcgk5iUD329kh6w/amm6
uLyiXU8mm0HXoFpbShZKm0/FAiXx8R5c3P2UTB0jO2YlN2sT211nJxB8NmKK
pj9QBpWVvvlzJFtytp1K0ziPY/sTuhlBKVh8zInwvI6Cob/BbykyFYlTl2GH
7Bo244tB0nqItu9ckX3XOKuXrZ1Db8fhi9kulvIl6XYtuAqm9b7SXYGIsISf
wkN2dvwnE4mRHfvOA3+RFCr+EDGZOxdTKn/G3/PS6fe7+Pqw2Gwz/C8SgyAf
/P0R1CH/zTTmrqnOMV6LX9LwpCqJYZzNmUi7ywWEWf+T6Ze9/Y+CLgjEjBYW
I+JnnCEBBP5nFgGIT7mPw7sv/QFk/7VTip0LvbdobwV3fxQci1d7PjC18MJ2
3FAk3ASRjTTRUAVBPT7AO4KC4IQR92RIKKAQptiA7x8e4Tp8m3V/HbMxRB4C
d8E0KNG7ENAYlCwVy9dlzwxax9Lg3CCE1XUxWLGoTwa7yFGM7e71qc2aRRk3
v80HFlO606o5zY3vEETxP3Qs3maJ/mivVoLxlzs/ay2LNSOt2cir4hWUhT8w
hpzJwZKGVnqjqH8O7pVdOpvIgSvVvvR4rGcy52vkSHvfOwFmOu702ZtLC5UL
+CsibDpz2fILcllohE+Md+J3uKRpSNPAmmSuYYxVRN4Ayge16e3J9wzCwiyO
ffSOoTPdTmr9+Ql5BDthDeTqNQQUAiKTg9NK4DZJQVQF4Q8x5iuQPOTXj/pd
gm4fpvEP6tzoA7Tma6nQozB6+jIogoawng9xb15GgEq1CKomwNoNNuhw6Bn3
ICY8JJA1KUWdtdBfVCjexSYIzfqnC4zQjKSR0LzNxEZGgy1008rYGX2PpM1K
hanEmHHrHl9ePJY05ynzfE49xNP9zN/PKEyGUO10bQdLCgoe6M4QgEFeHo5c
qvUghnLR/AsRqpqVm+2GyCH5tOMSd81xz8TgSML+UU8X1/PtItrQispJYRSF
JxByPMTn60S0QiHv/44B4ZT6rn1M1qZ9orr3rgQSSj6xbxmvB+KnWd6fXSjD
/C0TjoHI6LaBbdM0dQq41P92vm4Sd3qIPdzpfxwWTGZ4AL+rD5xGfO2ilOf6
nZ7dYIz8fRYpNbZx5ahp7vn5YuKjoeklKabVrzP+Qjp5keK8rxhl4xDZoS6a
GSnASchhuQqcSJV7Adh/CB27vakxHFSfDdggZdtrq/kGGykiI21I3k1c9Vzs
20YqHy27JWZfN832e1CBWIykXmLlppkdduIQzLjP+CkD46u70ZoXOStFPui8
eIW6Ok/HcgPgFDYyaIpt/282IqKTqFzNBM3utAV70t4e/tlktov3r4YPF+yy
LDLZEB1X5K6N9ixG1n3IxKZBbwfWlQFu/wtfwrgfZRwe0OZ2+n+Y2QexIqJ7
b+3CLslcPYOWnl3N5eEjfGI1IzHu0CLTR0/8v+//hwuNER1fD7HdB426Tweg
FTB+BUL6o03dgfi6mrlJTzWdUXpOXGu0/cO6+OW35ysEmatNbaPID6S6ysYc
7wmDvmEROyvrtm9ExEfBjVFKVmLPHUz7eiSlkcbZqsRF9evOXNoc4tjkrauI
k3ExCeA8ERJOqddqQ+XY0mx8TNeGCpzooN2EWOCG8BywBxf0zC2EkayEzzoN
dlpLoxDZtxKM94W1qhbH4AjrM6MO8C5tktNXtLAPeOAXZtX7rYGiBqtnr6MH
H7fhjVNWIwoXf14RVQ0JQZ/TzbuoMYKHTmoz9Kb4fCgkeZKftXsNJBc2pLQD
aP234m3LGy9qrKuR/RNBZuOeRMFibEZOrljAnapCmu5+cMFw0b1sLdSsLNae
Ap4wwljGjfFpPISeZkK9cUSKay1dbL34RYF8NLCloDesHPez5ibgzxFoQIbQ
wWkBa2b0lhsJPCIjUMqf9HayxrFR6ZP/H2bnrspbKCsKGdukX6hMa0zwF6Bb
WZwUWMNU8k9thfE1vtbqT8RZUSv5fLumNHkFkqcIFLhY7vdetAoHMxGZr/FR
9CbReNRbRpnZYy1hs4Alc5LQwFqHZGURtBh11i7SJrrcfFQtY9bbubMI4V80
+LM0w4OTxm/XhFxwjJt7i9/qhIjeUoXfWk7rGS63F+7dqNQB56x0R1ikSXHV
QeZvt8rqEIL+HKf6XmGB8Qkg/jk7hsN59SkMH4LFILawe04XvwByggj+Uc1Q
mcrUcxYy/i4psj/rOHp49ai9zGzpiAYdbAdz/qNANA53LLkt0jvLlTR6lfeq
NoMA/dQ6N4W6iBmeMy9DI035gckQHtuJcZugduxPX6nxlQl7D3ywzX0L4e4i
FAF3c/YHl1LDeWmx6si7jdfV/E2p8z87rs1THhUuAdJZrTccQkbiQ/OyEhsS
KTGyoU9712L5Lw238Hq5QLr/dxHkMD1CFpFhwIBQFDkKIVpPitgSgjsYcHa+
X+sISfftuicvH0LtCnZhDGYeROIROQv6dx/2fBdL0JlhNuidoqzX3Vbun0gC
P7DKjWp2ayNy/EV8hH0ExIYZrEnATN5swwhtUDrWOFAg4opNQPpc6NzrE5jH
TVbIRSVh3ZAltHGL43bEksrZDiR7LuUrgWMRrVrygitqCs7azZpY96yXU7Sa
ckJhE7zu7NuT76v8zZBNlgGI45zEnMDnUmX4H1sGLgQebTq1Kkx3lvfeS1Bh
eeOU8+Rd+Wu3zMdOLA4SfVVE47q34/R8DAPwkBZndPcfNBQWB+x4Lqkbxlht
4tXqmmCRsRuy1tO28MdbZ+hw8ATga/xLLZimUEauB8YJLJ+sq1Fvra38OfgZ
bfZkMoMJCRnc0ykdRlFc15hSoD3kXvY+p5+N2zHULMzTvl4KUUSbsydD+09e
rDeqoVJyZ8/X6eXQqc55rliMRXpb+JNHEznrcjraxn6gXcwxR5fExoDMEud3
5z5YhbNyi0Q2ilB8ayxyUasF547XCrvLcpiTluKj5HN4iXtXwTbd0G2QvVak
nUXN7Fa+G6XRLWuD2Mz9dGq4RATqukV085nhAHvvi0kd7YsITc1b6vpKlPIN
zePuyyVx2kQNHNCAodOf27AEK5IId/LA/MFaeorkgeD3guUf2dLSmHOj4w0O
FJJSyKsp5uFXshJe5UCG7CEeXRuHtnMbYMRAb/vpoFreT73N9zHukEHTV7/7
x1YjvrtBvONt8JPFCySn3EBaFjEjxNa+mDzTX9zFhBatxV65s9kB56QsR23g
mz+cG4JKA6iVOLuHPe87dbl1XuAGhVhSVNf+IL4QmZPPgSRzwHKE3d1Prwul
LFkyKj5xDVunVCQZFFZ43B1743u1U79FdJTJsmiYV0U8MTTWUqbIS6tTd6+i
j9GQcXBhXTg4hoMoPhCz7n55XwFdV8CTLD7Le8JW6DHVsxKyQtprukpZrDUp
3Uf2UySnucf+9XT4yqVJT4J4LaoZOjd177UOSQMfeQqzmtnOVfIAb2jcuIDf
SCLMU90sQnrjjP8OudIq6cG34po1ccHBWjFqaxFqE2be/FP7/XiT11um0Ls9
2Rrpi6FRdlWXLzvGEBXr334aXA2EFtxQkyOqezwGMSJJHVOmoQ8MVi/FX6Gm
6qXJVAQ+5d/VbUyTzXEpHxGhB87BsiOd/qcoUU0JsyAXu/+BnWVJXOE9uEiP
MBBNmiNVaW8bXR85XPvjZVNXBKg5huc1ryXORM9cfrvk1SV+6eyGpilImbU9
5tLIsRfCXvMd3Ge0A6AhFtXSCw2HDXhaozuLsnnjUnABlcC74d6ANX9ZZx1Y
PtegcMz0gaq8Jb/9OPBoh+ChhThgGFL/a286mFrFGF6C4yndJCIu5GJe6th2
2xZZfa41J5AaJ3qHEY5qN7HEgnH58h5MySYBpFcew8lIGrCAmuH79jr06lUi
6IZxNslCfep+UcjFmxFvhPwYSOmBIUMMrlk41bUxl1ccwktsULZ0vHhTmpbg
gz6MPA8isCmII5YHN6JnkYdk4L57WQ8qVzMoUNJXuQ9Hyz6vcacv+JXMKeJW
EI0B3uY28yKujskeUG4Uy707Un7Qar/uPx/iyaml6ieqq4/bsyLrJsGL34oR
wLaFAMiIbACn2FL7/1INthUtaXjIqjNf9AzM4/BBgEsUIIpi2EimMI9/bY0N
RxKNzj+PCpR11s4bw6uFXpvLM9BicHbyWs5ZaQlRpYYv+o6/gJj1+FqB/sLs
4SDLvAzW8nRe1Uyx1aSGjkgnwMNeuZxPSvSijue0fuH6zTDgIDmdntaCcxxx
vGgdv4HkFxv634QSc5Vh2m10ApDVWwAp3d2+T1BgfH9WGdJFbZJc6T/a8g24
dOxZkP+m3aG1SQ6U1mK9CxDxNcM9o0hn2zntxFcySmFPnfC9p+nGnerlaSvY
m29DptOQ43Ak6T97Rg4sS4w4Atv9DklJZlp4sAR0aT1vzikfl2A4DjzyNs6U
RQbV96TrL8CvqUb68TlWr3+MPMGTGLbfisBQeHepCPPq8ViHygbZfuoQgoz4
6h8jUR6ZTD7h+dfRuwWDxjM4TAPIBsMwntEAqzkEkBCZRphSYJDHLwZiq9Df
PtSBU9c+22N8F2wz7WszZwC0bi6t8L9/leYumGvEqcJhPjLY0ew60IBl9y4n
iPeuvdu2wlazWQfkeXz07awQIWA2TCaTz2Vx8YPc1Wv2cAuwWEiUXSg/JBIV
DoeA1sDXhH/geWJAIGPaSdjuUwPuScAsFWWWCKYsa/AI4dH9q6ncblo1nFWv
4VidPi23ipAAzp/a+7+rTcsCv7FIwaX5n2mGxI6toLHQP5+tcR3ne4brsJdg
BhaADVOvr7UBHya0QAUvAkDuJ9+MGKRUca7DD0JFrZrIE58vfEPBLyiX01Er
W1WAV6bJub53u3DB4l5rKc+Sk/TizN6z7kBlzdQTbWpDGm+/v7CwUNJKH+WU
hBz6xGXb/GxvxOQ3vj6mnFN8olkC8z4a3sAYDFxhVLOk21c3DLu1wuE1iiwR
o52i2BJPu9/XAewdBMND+vLOqxy+ae+p1LOQUkaGBP4TvJeKYVScO+o+oPYr
LWm/cusWaxhZHbjXUdBZvNAH2QcuCIUceQwWp/enszqWhJul/xuABFYqj1Nr
eMiZaIqZFXLzGyLFvmTAs/Z+HBxB2wFyBOHwaTvpHoB0rqBB4DLYfH7oH32K
2409khTUlQS2g+/Ou+ZazfsfVtvkB3fwNu8gga+NgvM/vBs4JM64Pnje5Tg0
sofpP5MrJMlUlNiy9nf95sR1iwcjFWOmWgzaFZr6M0H2gVTJ+NiEVtSVcBTr
gkfkyRvEgZ9Cm272YOo6hDhQ+cat6dbWu6BWLMHVbsAA7CFb5cLjzbF9GE8D
6zqGnk50miYL9MuZeLO2GPdL1EImAaqsfZ3pl+GYnSBiLw/MpEK0nWAYplQG
uGvWXhwSTMijYpg18YiDO5sGe4N4q7+cLLKXgiA5tkAniyYLQ5Qg6COjp/vh
FPZFmmwW+2YDSpfOEOWY42SaZ+H3cv9afrIjSyEWtr4N9gh7GY3gvAP4zPHC
kOPw/37Mo1gG8siMbNtUUlx9t48xtD8fvwiqR43ueyoZomA3rgDhmKt+mPrb
MIuEsFSGcfB/GQ62P1yIFG6c9gckNAETOxveEnQCgHWpJhRmtNsmfBK6vuj5
4bfnB273w+dZs+dFYbewiwOKaCdZUOMP9WbvSrX/arOUO5sjh9iTK6QtxCe4
wSBjsBthIxWDydBZ0MlLc7lOswO88aSh8uR/L3DOh1Hb0QaC1uGogBo/gEt7
IyjRAlVavTIRLKI0jMJ/UzYOHfRRb+9QdrFZP+KoudBf7bx2QslcPqXa6o13
P0SqNmRLJ/dzMhCw8KwwWFvkVV8RpBfbpWD0AsUtJXuG+wE0FU+wgP9BWOu8
h9wWS0Du5koKez81Oi+Bu9ag+3KrLdpt2bEV+0xGaWe92hqpVpwQrIIHlE33
+Lro639jQKCIJ9bg+t0zoteF4/FcsGr5cu+TXi8nDC61LyxdShFxN2l5recy
w2k75q6SShx9UxbUX+sF8rgd5YpmdthL/uT5ToaeOc3B+zt55wP9uht66DHO
n8bfK2I5JbZhR9GQJBkM9qkzRf92vlsgJLJnsTgMiZD3mhHYacgtXuWndgMw
9Q8KCTEnOQhT6ZwJWwxHaTpfWMfpILimxhvFIzvqUfjZsPzaGX9VC484Y42y
0v/1nPKcvnmfutVLC0fgaDAHEEcz/D0PALyg9p7+/xAXaNN/Mh9kE2EPfF7D
BMtQ0kFZMlk14i3eneyz8IvKQ/v/SUv1yQACcTU9DWkgRSR2vGLaiRxLwbk6
QEIn06S2gUYluxtQ+KcxuzW0vzeWk8U1LmCHQ9pfkQ+7U23qpMq5yIM/AXSj
Lsr5uu65ebSUaroKyZCzD6+1leLJwrGiVcm83tF53I7+QFQb/UOZsfHCbcp3
X3ixt9jaBK6UUrnClGBgJs/CBRzuzVMYJgHqVxBDeD1A2RJ1ezsUnqMdv+HQ
99/0KG0LVlnGAccy9L7+e+zu4gN3yrUpsUhuVVT2d8VX6A/3oHtIlawGUOgl
ujNHyBzDrXVXjvi8asGvsXjRaS1nn7iriivM2oTsi1UiJH/tShLu9wGs3Wc9
NIH7TrOZnfkzNJqneUGv/RCqxKXqSAYV2w3CAmu1Vqv7p9OZNd02D2XDaQrH
L8uPvKWVAYgeNLkmvTdoGiGUj4oAfvK2e07Y/YNhAAw0u6soisFTgRWyhtwi
oGt4X3Z0p6geDPmQFOtOKI+taFDRqC22VoO8Kt+BOgCXxLvuggeZ2LQxZI9G
BDTjYmcin3QMrx4f/iKuibzbdwizkOxi9rVdR531K4Yh0tzGSE4SCdhYb6DI
tExwzZ9XSdJNrwxmJSSQeKvIhK9leSEm8Y5JLJ1xzded90KePocLk7MVZzeJ
mnc2coLLgdUWDAnAsT//ZR9LfNb2lHyNfIUk37CKx9wMlYwI2jpI/+uWUaM9
6pY44ehLBdcVem3yjKX3ggFSnBV/IJq7GVPbHycNu7+fEetozoPMh0Wurbsp
JHV/xGJmU6RkjaZCG8OtnGXvW7H7KX2vIMUvxKyTNYgsLWWE2bTQz9AZO3ES
mC+Erin6f2/cv/SPzie+o/xQO0QM1RuCnX62t8vZiyy1+nvWwhtUJ0Sr/a3Z
1xdv7sXe0uyhrnB0Ba6kGpC0noEWe/dZsG2HT4qLsBeELD6pNe8XbYvCTV7J
4rflhfUF/Gcafzpo+f+2qNVyxtwhz+yMoroIeE5e2MbrkbHL8wPM1jS5WKNB
ek9nCo6/yCERtCqkreLgV+IzrfmoN0u41rqTNMG7qxGtPs4Q14gisPUE7t5Q
rx+KSzpYjlqssd81PlTjNo1UT1JgklRXt1R0I1p+l+tOFDRO6CqT8xH+xZkZ
T/AuOolfUx78917oBnKAicf+e11G3xRg46efgW47nWeqtt9c0q4c78Fyiw9X
wXKJ8XbKLyHeTzqMzMeJLlnHbUU8TnrAfIKN4wXY9x3TQnO1EDCxzSyrC1QS
z+N7Fxeyyyf/7N2wICdGWNv9j3rtJbBw9FuDYzb+AhBfCUwdu4OA9WVcHO0L
0/Ya41xdiSkh4FjIZxFsAL7Lx/23awDFdQY5BGjwMTlljUz5CYpKrNHo+uIE
H1lB0QG3mpL1H5B/jeY1r/YpI9gV55EBUQss/rSUW5jDbjborwiIojuGO95N
PCieiG7ZAXrrgUA5IrDGfYDqjxQdqS8ySGc0S3EpaYvuDtbetmCOYKl3vXDY
W3GAlNj0yFqgiKdK/kCemqrcSUIsLYcSNJma+xzo2Ml+LB2WlbyLKfyZz616
upsVUDyFvMJDnX+lgTdFuRbfo8o+2mkslT6w4GY84YfJcQqKGm8GQiAxoXgr
AWVtwGuF/fTQWwRZiiBg5jOKHjNyBIV71zAgZBucY4K+/5TGyIBZjW+iIAJ3
lw7TNkw872U5di6KPL9ZvFNThx32pFWiOleD8+nYwsT6VxPpwH1L1e72sIpA
giZjAAP39+hpoZ0t4ECZzZVE65y6jML0aRrJBP+yIbnGpVRUL82geTbOZiVA
EzfmrdTDAc7z74bRGjtueUVCS0l1cs6/2HrCazKgUKFu9Yute03aSJIO7juY
glV4xVSCaXoIVxvdNt0gElXxZ2NDraxcQvgeiFuvp1P+hVw0/NwI3E3/MHne
s5kLXK+z8R5eA1IqmwqDE3cr+sSMpsoM8BXc+6iCda+/KtgxpTLDSHjuciZ5
yHD6KHJX2tQUL38siLvpobc5dCaamcPc4Bhi6V85gdLrP/S4LM8dDvvTuApN
WoR+5U+/SvnrwLnZ7KmsXh2Vf7WcZYCKwP18px60UZprNUcPIrWMuZUNdGH8
pUlZTl9uTutY4Lefb6uvS16wKyQXM2rL3WHQNaVJvyFEaU8r6DM4O3/Uz3T5
T6JdOu+K1TjWReV9uXvjFnkZ+Yo4IbGmukjQjW1sujhOT6SoBbKdV4vUO+7a
SJ+xAVmjLSo9LVR4VCpMOGtV28KuqMbSq9gdPOA5WGu/ggcVwiYorXW+EfxG
CVi8HTnkVgcgzP/e6DcW1ecVAUaI0TA2WHffbjncJNLn0ORmJGaHhdxp2roh
Jq9Aw37iSSVuKH8GEpW7r3ImjdIut1K7Jo16eQ+9B9OcvIKD7Qlf+tiC9rHo
tVVKSUubNK2oAiTa7ZAwcOSmxm4lVKc3AdpFc9Ib9KvukRWt9oVjH1TLdmP3
aeZOd0ozn5JLmjChmSVtwZxlxHx6jn0+O3IQvQCTpFKmwjU6ZcgVZxEtabdS
D44v12QvHFAQAF0paED/ipmw+bLT1MUr04dQJZToxxwJMcY6BPNir+CkpCIt
GH78Xr9FgPgbKmy0STafpvlDZuVQIiUi9NqL68JOxVvyZEI+fbsaQbfv/5hy
pA8SVrYSdGrFwaDSXHxC9BC5dzDHi/QB5xakWIozBopzXdu+2RlyX3qgTkgQ
3O1oaM32JSA1oekq4F70ah6zA/MufgZ+BvMgpe5UgmfePCYvvbTayATabEgB
HDKX2y5B7aiHmHXCGcHSWAc6On9GR3SZ0ireXCYJJM0SbCSa34lvc56EcDLS
yu5teKAR+vLW6EHwOKyzXOnN+EGZhhL2zoJjSEtLGU57MZXvAmMuSqRvz81f
MmYxxi5ujuKxxB7+BIzfSKUsqk3i5+zmNNPd5WDEE1hr7YdKKyaLxvZcC/ER
lCdy0mKMXNEdZKFJQUoheqC7Kb85Fv9v+JsyCoMGcQGXGEGCK19nG2sD+7PF
7ivitplf3U1LnH4wOiZJr3br0fbg4NSDSDGm5a5qhTDH358fAi7n/gi+LsQp
XLsAHjbilQC74QNw9IRPkjEty3JYkzAsh1c330YkGs9iOH6pMZfqex5L7oDX
PJ8nTVhYRnCnGqg+b2ufshr19bLOC2EGU2DDaKUK0ocRU+HB4+4JCIBk+vEF
ZMYrPPpsuhOXmhAVZQUDGPOMoZHNC0MB88XvcWv/4HfYwxDalWVaf2OdoEfm
CQLddlzx/e2w42rlONwjPb12fGqZiYyjalCC+fhF/CHURgthrVP2UX140wE9
4ev7KkONmK49vDyZuU6GmgGz9IZ+FrejXAXjiu4Qm+VTQ6C5jUjrW5Hx2f7F
GxIDoVRKI3pOXXUUNu6lC0yKN5e38zxCljN98c9mI4IMS+lcTY85M456/8q2
G1cZ00UcFu50lnFk9Dxy0VfjMTbFrlfy0MoADbWOjK75teCQoF++riswJloz
5zMLFLQYPpF1l7GaL2Ms/pDY5b8ba2rhnHoXU3u4mHN0FBF+dLQduR0iA/Sm
BSFmnm5yw7MVpE8+FxkZivle2QkmDENECOGL3VtMNLplLws3S2MOn/RqCLUU
x32I4+sEcEsjqT1ojknSGJvspxiajNvoPrmMgQ/Slk4o7TLCnsxo97QnJcOP
7DaVrs8Sz+YeAna0AFCDvRSAxkvAhGzBwcA76rdEYI2RkgDw6AF+IxsYmVCl
k6AOHKb3MNDTys02V3TLrwv4BpvpIKxIKslspYPJDRmCHmKsttnrXPCVX4Dk
vKExIfATjyvQ0zyPHAoW09ou9u1cwOWXaansHc9KXBuE3gu4HmZhTcuO0j4T
tl0xtc+FhDVGHYjT2UYopRsTK67Nm/L8KyywH276lENXFLboSnItsgzC4Lo9
6+FiXmNlha8jkOZ9s3ItXMUk/EoQzgzWbLWabk1FiG8CMp5/lSB1dDWlrYzq
JqTP7qBoBunmnEy3QX3mI7/nwwHndeWFZIRrKjp3RE717kOXIzIr4HBojG2T
neC2gcksZBaJ4UNHVr/BCmkvwZJBOy6yG4O0Bho+0T/Ddp6OWXaUtnXsIwSi
jBHjG1jdPlLUV+38fr57YrkPJL1Yh1HN2TGICF7WHLHUPTAf2od82UhvlKri
9r4BSAyePAUWQod+gVEV0fW7L7iD6VX2/3gNxuSHtswL21BR4jqAC5Mm0trJ
m3+y+Etsj2ltkZco2XMq+VYdA6uRwgQBpI6KWeHzZfeOSATclZ0TR0TRVh6W
TXbcmCz9qf8n2NEmD+ropRys46bOuioHXa1IkZa8vRkH/VtM5Zzg5sdM1sjf
VXoGIXiAYar3ZsHhKo19zMnwVUSv/kMWzVqLUoqsPlccb3J7vBpjHyoWf9I7
FVkfo0LO6HFSXgIm+wgA1dEDrvg/NJ5VI7TNp9FQPgrQ0MBgvd2LZQmjxqFe
8BM9fpTDPIbobmVsSfNuI/fveZFC45RuLoENxZFY8yEk6aS5IG+l4PZkQTN2
GGwHh5WAxXoINarZf5aZWkH40DORu2uxDl9T9VyG+rcxehgOprEPTkWvDPoa
4RTdpvMLJBs1oVs89CE2+12S1zGV8cLuHG0oWf4AIbBm2ncU2Pv/myc/XmLV
F4WnnkG9KRcbwDEpTsx9SEEySAY2ArI60eAJM5mFGHJ8pM/Q3hWsdC6rpEJI
mdVEL10ksXIUtPyAftQxenntRJ9olduKHboOMGLow7Ljx0RAvCRPAejXD4r8
3gMXSoYOm8nSmHU1OkIz6wsYrYTVi+tcrWpO79ShdO1g6r/4uUCtmgw4CEVT
albcuGjl/OfNkECLmjkodzccJmueNXqRVOUlNHZJogc9N6Dyu7W7NAIh2NW/
8p+KeVNhLM/lBm3U/WzScQBWLIBcYDWKtkuXEAQVYL91RQaSoDtiTwV2j2FA
tLlujWhOWQT9W41NLDhzFqHyvilvTToCwET/qzo6uSulvsbBUZ0zXa8Ry5eQ
Uafjo/VEqQiTv8Pwf0w1VyGWefkqayyp83YKalT4K7DhQn4KtE+WcF+RqGzC
Mr16PfyQdIr9/KR1rgc97TlKflbnrmLGtUgkzF86jlVxV+EtK8T9xOmFXD+k
HLOS3Jj3UKH+/uLVoge1JY7Y651hBZczcY8wbkC/ylyBuQG3g0giQn0LcK7m
+KMvnyPg5xFUVRyRV6oBk+vlDlVcc9YmRm8DA9WOWHtf9CXfOxVhDhcdqZW2
4F6wdAjcM43nq05bpxlsekBryXi7XYkrCzqazvnIaX9SChtAXLLb6tPS67z5
+3j1YUq8v9LIu5PGUEEjuNK4vjPfCqqtkeGCl0BTA4/RImlUpd6Tc1PuTPI4
/M15DbuVpQiEXZTmOBjiDK1uo6LWzO/2hF23s8A0boMyfaK6GSjFUTmIFpfA
uitYWNnCb53Vqcgs+1wfF2W87jFKkYEC3ws2R6YS3f3CT/tEBbLIYXHvnruC
NAZKSBD9N4hwucoALAeRSRU7F23N1LCltm/pd23mCdb4gDhzKRzgIPW55aon
nixvQSP/9FNjMauWp8KJ4tf6m/dSNrLFKbQ5TVkrOD+UqxnbOKnpDKrXwQCa
myZq+V/v8LtnsXhqGO+aGK8M7Pe9RdgtUpHvMyzJ1te/BIb82SlfBV4Folgp
Hut+ApBdJPb0fk0X/E1pLY/uvXusL+Expq9pruWE3gw7McaK5hzWHLJUtbwd
hMN7Q9HHuUwxRTgtRb3GLNMsxzNc8Vomu557i0Dg3jhFugYc1cSHuj/eG5a3
yA/y8pR01VFWR+XowZw5KOEZEmI+rVm84WCnUVuuBCBVhKewJOkOERrnEV4w
xcQbHGxM0qY8Qul7vN83UFamygU40q4wOwTUmwlv30mqJItGRaa3B/22T6Al
0fzWkn1kVXtzzt4D/EOR4t+qBLaMqFdao+5qtILtQPYdRnZrOPEQiajYb+FD
Seg8bBPJLjhq9+AbGtHbeyXxsrtRxi/AuWcLcEQQXgyI9WNYsX18msujhIxW
90LUdCA96XYLgUAVrD+5LGgLoW5qFRNF4CD6VW+1msMIzUD5+VEzWwtH6URk
oUwbVn8NJee13sndxBm5dJsZEr3Oxa9MQ80EaLaIMFKzz4zcVsmA0SB+ePdZ
93bJijt5FPI0+Nb9kfFk32FrxGDTjxfahTqvIBTc5NjjddecXNjSO1AquXCX
MvvMgJQNt7fvSq3ovKmW82EdUUDCiM+QTZWELua0QSajWmTQrTBUaqAQyYt9
R7dNwogqYWAewqG5LLo2JsN9M/1Z4KgFEYymtCoytkNHEsPDkbiwxXZ62O4i
c9+7rLQ4HzBesFlsVPi5YoPyehiHMrJ1f/W5BSvH9ZpxbiUF5NAOcvrbyuci
hxNyIlMCnOLG6eh6/xtiKcrUQN1mhYB23FOiR/shydrWQsq2N2kkpw6+rSHO
lDU+rCH3XLbsErFt0j0GYt9mRfYmOcZbBWcCAGRNWboYmDpSguN6LSCh5QHp
gnQIb2LFCoV6qVT+npTdil5VBxJNGj3n3UdebNxNTGn6URwolxNeKwykIGqd
MHFQye6hDSBglkqepBLY7dOG4J6RQ0Ah69I+RX7/QyCAwCvHi8ncYmasxrCA
GlKs/W8rde6X6fByCa1OrxiYBq0Rhsc/yEUHg27p4WdIx7xWZ9kA5SMZxN1O
zVvR1wHuyF/DCM3GIGLLr3JMtuJ9//IDLzKVeAqsZjFIZyLI3NwzTQmpmgaN
5sNgzfvL7qVoRIPWVgeLpAs1YAapBoE60H40I36BaylQH2+AJPvI8/T88wHb
JLsBQeRWbDJHIaDznd4Q7pvy9ggOIR520tvv0byXm9O2q4ilVJH2ouJU9+sE
RDpl1cyu5l8a7XmOCxjCRhpA2zmmuuaVQTNHRDm8nQPivok2hBXCXAYkGnix
yd1Kqz9RHCy/oepWfdMzYko5xeg244qlntzLdtFOzk+UraTJgwy64o9C+1+9
QJVl5Ym+TbT7sUjh1AJ4O8MecbjVBapxAINMjWhGbHtRi0VQm7rBXEMRb6Ex
eDbU6ycGa6oUHCdhszZsJ1LwcqdugTcU9kTAuySAqiJgELUPvP388Lw1q4ml
gDQJtcBfE2iA1kbx50Kx5KkTOVN/11CA3wYcZhiNLkKRz+A8Mw2Z8XTR9Ne0
/E0a13u6le2vFZW3FgKOv5cRJsY+uWqu0bFp0HkKcz9yNkLGe5WPdvVNz5p6
oLYj9Y/SKrl0K85ulrBWphyKwD0Tc0ZplqaQAMNEU5Ye4XbIt9JcGqxZXvSG
w/hLCr5eW1F2lBfDsTueZDijv6jcp3gLT5pLMJKRNhnBQNU97oOw0cWh5Km9
qe3wcrwEjk/iHOUhUwMWsbnPsBR7kTMwF+wMagA8RJm2qOXoRUF7QSU05GO0
AQ6y2uE4A29KSPVyFjzc8b1bi+rHBbqEAlV9ywUa0HznOEU/Q3IsnaSll0/J
A+IJaRBjcCYbAN0cWM0NwUWxNPMT/e99jiJGS3J3somXVEjufRnsrolTeAFr
xXkb9HhSQzA0PXA2sydrqhR7X7nAV8NE/1IZ13RZCLb8jvd6NH3Hf/qCTP+e
4/bkMPel/+baCw5vK3JTFCKcxYxes20i8YY5n+R3ro4uRX4jfBMcLwdh5fEf
YDZSWcPXu5WYJgWouAYuZp99l1xCx92HjIPa+vqjGXBV6m6OuB8qGTBfnLmI
1x0Eh3fG8QcSezKykH2ePhv9xn5At2NeAxmtOKVA9a13OwyZb8dKChPdulvK
BJLrK+NliWw6M7KQAZFOhG2yMfQKsmoM0oEYkjm42QgasFPDwwfpd9aPgHCk
7jghQp1IvPpAJRTSHTZY/U3QTvqcrTkPV5vNNCNTlyJGAI//TB5ZXRe2Bdlr
3cwC44ieR8JfjLMaH/RmFMwymJHZSMZEBU7F55d78uDEJcGGwE9XMLQSaDsG
dd8niOGLHRz4z3MbSK58rcb9BQwPpw8IOi3slldFlUsT1gdgzWPISrb0Wz9g
Z2ov1jjvKZYuDjvkMDuu8I3VtX1fa0mB9ZMHwiVByv1AA0trS7rvNJRCa4DN
W6t8OPK1LA0sORh7L+f4uPF/LUHj4sIc7j1w4bIKOS06Dov2VWpHBTImBddf
NriA7huuFMt5bNGEmNNDcNWkMrjObJzQJVEimn281y1IYFGW0VtOFDGmM2Tl
2PR65Uq1/knnCE7Zs2C0ndEWN0EtTPNP2MeJ3K/R0CbYwT/BAjF4/mORh0C6
7U41RY3xwlZnNfNlZD0jiLA1SRbCm1M91Ctu7TlSJwA1TX6Dfe0WUGHIqntQ
4MhCCvI/85g0RtMY1JA84NIy7A7WNoqo6KqLUnheJYS3FsT0zYyJ6C5HPndU
S2l+Lb2sL+yfrT9sU0Ruh4eDsJdf5htLhRS8zU1+ZpJk5dmM82B0XTP72/RW
tkKIb/fdpy8JjoF2fQCx0StttiZFE5WzBNqVo9iVghZk3CvPyUXNRG75j7WA
4CRMYYBX/Nuiw2XvcjNTFuIzl46u4Yjuu4E+lEisMANt03uJ7YEDWadnFO8Q
MNaktrqzmj1gxPhNlihxAz9Y/S0sYQOtqz9zizwnxFPRjye2Nu7Gz37llpCD
sJDWjJi+tZ1qYX8ako7OSXeQpMyQwPHf++kZd0O1ctcIJjleUdnJNEignkrF
KbEhPnJ+du96+REaFwB0CzuO4auvcUmZgdfG3blr71fAUcdKHKsOOAPNCbuF
1NKPveRFDj2v1EvJj6tk+enprMUU2RlT7Y32/RggJUf5M5FxNjD8MvtkgaNb
nBtf4jfQqpfq6/l4/j5U3GKGUvPd2GWuL+8WFHsfj0zRYLP8VvMQRzNEzgzU
px/xDziyEJD8GTysmuKu9UNmSKPsO5rz0MyYrsdQdS/FaHZ9GVlpej3bXdWY
1/0lR+JWWqaYhCcXxCSto1D4CtS0/kdwOF+UZFHJ/emKPrqNN3zTpbQ5xH6l
Hqo6LCA+67JQiwmhdPKY/1UJ6k2Al9X3e4/a/2wyyYCLtw2Exdw8ne5wD7Fp
dFiAC1uFQbKGK1SFBQ4T7l+LkbkWZ4mwL0NqiTve+PPUj+NAyNyEhvJgMvqT
3B+Qk6jQ3Ij5MY1T33LsMmdQMtzK+UEwgEkHh4jV7yUMGI6uui+wj7MC9DOx
py1A3Ix2lfO+FMUT3SZ/3qbdUghLfyXluC1uVH9LwzbFXoCTd4rljchZmgfR
dFrWSCceHQ81BWKrJVBpjs5wGX7P9aiVy/LOEN9z9+ZGV07Usgh+kxXdKXC7
EHsEIkio2WZq4gTZ3HJvnYrBKOvkZRoUvPGBAcf+hdK2hhiGitXoMgdMfLRk
LqWM7hBCbwkWSKrMcwy9hmFxhcdtaSdLEdq9qAHT8Q/8oMzd/VFVsAUw/6Zs
JTtN6pqn2QJbd0Bqp1zdfZPW680JH8VrdMjw0w3LqM2Hjm7qkzTUl6VY+fTW
9Yw9pnCFkL/ntus/kFbMt5/W033jM+XvBn6fSGyjJYIZ8YgiXjncEC643EpY
pcxy98AiSDIEgR5fTOK3qb0+GMGEtSSOcIhSacR1fxs9OZ0aH+431uwRUDlt
Wns3PltvriBaKb1Rm1ioO3evPk2SeFFdltstgx8Izy5qCs5/GVwpkxvhtLo+
RtuDaQR81ybKzG0X9zosx6mzIOhEuXYghIr7Zy0r0gHjgjqRhWkczXfLhhr6
k/wmONW6Mv0WYXt6Vxhdp5daTyZT1VyfMOUcZB450XhJb3WkJVW0iBwQzso8
frDFSkNDQ1kbdXpypCqkFXVB1nqwUPFl/EG9JqOsB6h/vdPLPvDaDPBYu9PA
7u4IumRQaHjWMvh/qoqIOzgV6kEk9tqAqegDpHB7QtNYHVjGH3h03AgLB6z9
17sGLDlVIqZwybuvExXR5inccoydZNPzRk9RAAQ8PZIUA2p6pLy0Pp2A2yI+
LuheB0lY3JWfIO+9CZo7c2fhBhNSt0UhYVqSrPWpimEObtSVgxU4vRXi3lOi
UeY4K5c86HwS0hlX0Tdo1ddOeJRCtAfV9fkExTXXN1ePMZnFQfAbSXWwV5DH
IFVZRt6pYpD2jeFgCReJ+18eLT30uahA0Kq8Rf/Fk3hVjOu4wA5bo+wxDqq1
kXN3mQk4LtVbzRQHzlvndh/5GEK1Hylloep/ucBBTbSXlJKF5yDWIdf5Yrfd
mf8tTKwL0E4iEvxmVTOHoWopRctteFc1SaqFufRHpDoe003AlUmIwMPz5T4p
eIL2/Ufn8VxpvmJrrssjEYHuSUUUKGdZHF4vKMQdIFYbNMIvNfpM+EvUO6jw
/EccZcb912Yi52qifgmP7uLMugPieOVgSxO7eU/9o5XId92A3xiyX2CPmR6p
v3OiCCEiNDiNx2L+zgPsv99LuIFrCMgGDyqhgl3ElXGftlTut2rtDEgia5zk
C70BeEp9bNmBLTEIr7/G1OrDlH0J7YaTg8Nl6lASIb1jVn94OrN9AaKNmDo8
IGWrVgasAZhUvImwCmJx+50M1zVl8wVtdaw19gKD5gr9FvD7ivmmFlktaauF
RdPhwPWEnL06/8dK2r8+97ZEA5yU86av/SatE8iMK+Be96Oa9YfD133L4UO7
e9MT2OoRixoZtdlYc6esZRNjds8Gmr/MuP36AI6cNdhOpQYZco1WOvaBLGgf
Nm3YdLGws8VA70mwwCQlZ9Bu/WxW0G9J+EnCItYqWu20ABvMgXxlZVD0kETY
eildCkrDhvTuCXNhqiSgfAKOt/yR+MSygwZhTVb/7kom7IxOaULGP4dl/Eub
qcq7c0KEJOL0sNddlxrqUNwwxMl8lINpzWoeH/rtIBSKRG5bm9uB+w6fKB8g
fiTAON0cJGitCYup2MVGUv2lXZxby3NQ+Jar2tODjLQ9jZ/N1PrmkRTHWDh7
fsJDKTKuLwIKiOuuL6m7Onj28ytEut93cespbh2NhRTB5PoOcBxdhRZkpzlJ
eFjhI2h16z2WaOIeTYr2pX7n8uhdbA1c8jxmp3TBXoxc29CR+RdayB6I8FKw
WHi8SbBQ6gKcm5VOsz31TCEAqbqV2HVqFDedE48PfkvK8O0wj3PvqGWomnwi
P5AcSmolkXZhirGZ619TrtdskfqbFHJYDy5YKFk08ReORy1yDFTb6f1Tyl4x
qorut6Ac09Jn5g6uVPRvnlQyTtc7wTeVtxs/9XhixAxVHpDgTbD5L8wxWk4F
DY0eTLiLkUuIGsZHx9/oC4lZGeSVt6bLRUp2qMQxFXzqML6D6sNO72tvFu58
PKpNS0yNf1i5Xs86jav/TUVJsu8YGU5z7gtpi8ugsTXRe6KI3/2zFyp9jvY9
CRX84OUsaqNpOCUcKvL1nRqHn89bJDwVPSyv8bdKNQSh9qas5zqnYzjjwxtj
750Wj47Z8TuyTSPJaYHwCHtZSOKTABEigBfliB5M7beDujvunXNibifOszJ/
uVbprtseW51N1cNQ6q4ORN4fTfsOZnDsSvj4HmZ16HhctMbKoAzUd612xmof
ebWYSNTgh0ZpEaPhZYh0+9zqTiCrzUEbb6V748SWw9Tgg0wGi+SXz9LfnhJx
wMlP1S2bFarTbw6DCDfrRJ3+90Y9yDOjly5rhpalTwYLca4ocrNsQI1v4Ufy
jKNFqYzGa5nWt/0LDYa4aCAzjvai9FohJpCUZSpMVejwU9Kxfpp7wbl39Ls3
dRCJ6U+/Qocy1d5ZgnedRUXoQ70AkPJgCW8BnH48bep3ir7Bw5BO843Z28Gn
IApI54uKuuLtU5ELJC9Vxwk8Py8GThNNBkUdDt5GXU1vJhRXRCZDOscGoqn7
t7cyoS2SjHIA0zDkmFgq8yxXkTNhYLvpMNtWNjK3ncVv70Nn3MjCt6n0t4xf
VVOpDeWcMyVacu6+Zybvjyw9yf5G1YWsrk++FNWw4qeERp/THz8iCjxGN957
VAYc6deBmGjB5Dwyyb3MnqbULOhwt9+CLN2zVZAKYt1jAng5fCZAy23aetLl
11Rf74f4rC+IcV1Y3E4BnwmnpmGQblot6gJXmjz7nkoZl6qmpGrp54pPQtiW
4huzqYeVgvbO+ocUUpjyswijDEIU2ITO+Wlmtm91RWcyEN0NqzAbHsZKV5vK
A374AYVgOI0PxuO2mB5KjYe1zWKMqh8zZRW3ZSCkMzt62CYjUt8KnTcCpQxG
XHm0kDBuoFfrzTXpawZBOmRJXU/uky+n2lGXV6EBtf1fgC+VdaNx+msmyu69
r8acE4kAks6utACebSB8tZ+DOBKkTOBlsDaJ7yKG1MzRQYSa8E7tdM7HPTBT
IrO3qbO6j7Y6Sbhx/kD+cGSkJMuqRIj7ZnsVFDKP8Rk95seBil6vMNlrEZSS
D1oonhUUyxBriS56LiBv12FNHwNmyb42ELAM5ziWLQ+H3FHsW+wp/3/5sBev
0G6+vQ/vLfb8fQRxgAtbDSlY2q9whtSOT84uYx9aqQZL1W7dWPJqH2LOWjqE
4ac91a1KfUOU3WKge75Ac9VD1NQnLiIx5mAQMncgSw7PCUllBwv3Y+qsvWhx
WoTN3YG2X8+wRwIv+YEgw8FQbDLYTEa52XI0zvyfACAzOp87wm069WDz24qo
ysljWe3Kj8tZzYD2IpIRLqqqvwkwjiJ9K5zGxn1o5jhE1rF4YNkausPF6zG1
lvhSQOHu97agTrsjBBa6/xU0dGixZ1E7PNIc4XPsLFvntDhhiXgzri/iSsq6
qubKbjvg8m6FO5xu8x39HcSS/NMdhuknO1OK/aegCFA6p0/up/qtGLZtJ5Uq
LA31Uc9SVFUrtge6kkcf+eqbBBK8if9aQvicZ6wYHUu6MAJ5UkHcUdW8E4cc
QkuPe/viK1ecyw1mX4QCIjGZF6KJvtgnSBDiyUCYJC4bJ8cu4NtjPBOnb7NY
5BZ0e0b7rmutbvyvCn9pIRwTDYbQ7MY0cBFP37oWf55LicUGEez7qgNJ6O9/
4fEWlyAB40jwBqeIsRs+d+/AD7eg0K61qo1/DCvzaH1ThKXKqFTyLGMDK0yV
lvrv2zct3mAAv829GDDUruwI3xsYqzk5slAOwl7dxojoO1U+zoMRFby+/AcS
Rf/IFFozFa+xXaZ5/5tMYLg1VPpxek0r9e05r2jZS7wAf2JAhudySnOy6UQ7
R3dOsxZWHmei+dtmWInUwS+/DyqeZK6LmJH90RxdRP6DyhRfnTRWBMvVgEAA
ujZbS7jGEYJ6fJxAssIIS46DQSoNEL88kF0UB1N6FMH03lU6ALnZwK5EFlaA
wNuc+HoM2PQ4wbhY4j2fKicfFKIpZi02voZy/wPg0Xoklrf+jn0ei9FCnQML
51AGCPse4BQ65tepfZEc74B42ILz4hWq+ZZYhon7sURiLzUuIC2BK/abmIkW
JgGQYnIIn6yudck0jW7DIw+54/6a5fr9j7wqPZYhUyKfMhxT6mluHf04uTAY
WQCB39F2DzBBg124T2HHxHgkAe5hI5bt9WHbZ0ghJb/gAIRPur+I52AZJjCK
N3BqHfKfEip8dtjFZWJh9TgC8qY1NNZ0n8/HTStlxubH+N50ekuY3+oVYQdE
glvL1S5kDAeHsj6mM4pJZloQjc7DQSOtoY0hWtgwY91Ej+/H206PUhzENE6q
53W4Wc7mlC34iinN95T6GNOH08PUMiiGTzVahc4+Z8c/CnrtpG3yKHre89zI
W4h/RUjKrcs5eE+I1Y1g78Rr66batHaWiYKqUxX/AX1G2Mpj4CNYXrAlo6KY
8rsLnhsi/9Br8agfNE302iTMt6fVqSu+QkUAnQnmB2++Nx4vBtgfBZf9LXcu
B2N5dWFoS0as6yZU8lI7KcqMXEB8ey5EWHAX+P1/ktbd+LSTr2x/x7rXxjvw
uDINXnNTQurcMSEMFJNhxFioWC6F9CMFldRr759sUXqECCVzYatAsk+vmSYT
XbAAfjAcHDr5wMPB73LALSDCY6OFdNWMHdzEuQU0Tye7CVBYi4scrwwnp6+X
UKNkuoyQs291bwQAddDWkFD/uyX1oQBURKRMNZ0Kjyusq+xhO7X+QfZnyZvj
9m4TeHzHPN1ZvbE4NwjuulTZLC9B+2oOvyVtQnR3qKTMyV0/rH0DQ9I11mQ+
Sa+A12AYXbRyHjWSu2m+eUURkxqGUrLHgRKqB65gCfUyMOzD1Ik6BumU1PF+
MYK/Cg+b4v8aWl2EmFMBeRqZzUloH/rhc3iyWbd8Fe3o1WN7i1cCZNVSpq+P
fHN/qKSONttMqd3WXNVg6OxVpzVecFLAyX7HAZjLfIGgVZYaHtkd9WdFDCDa
8wlN6UrX4ABq0a6aEId06mMI+bVqVXGkzLw5HP1X3nPmPZ3s2U4wohzzD2VG
I6Dt61tx381Zcsq0coGlkGy4aCZfcEa+ccNVnx5TdNcNjYHeRtgy3Tw941cs
dSTHXHkmLR+ziwYIxEuhmwir6wxSAeGBIfQaAtJATKMDhPemcLTeImKM3EKx
+/DQwL4bV66o3KUJXEsYMU6tmlmE29LB9imPRVupeQRXIc/eJeH+D5KKYfkr
bWS6w0MoyiHLgBBRJTvu3gFivpGYm6iDU7p3bSazrA8OrJbGpTUOjGOKvAXu
i+l6N8biTNrL+HRcvZ8jtyvBRWcDMIoxVrDtraMfEfitYigYtfZVTJVRLwFx
ssAUwcQ/xgMn2Ph/k+KlCRXHoGviKDxZiGmfhpHpAwFqBT366aOe9FyOPH4N
K83YeZhGlWz6GafRRsx3//r+y4oKC2YYbs5Rlbk0xYiAmkOWsWK4MG1VYhiJ
hvqpBazzJ5TpvGy4X3uc64sZwlu0PcAqcvFfFv4YvlShETuhXbP+Fn2IE1Y/
3CVyucj9Sn/ciXvaRlNBKHeEQUM+leOkw4wiSQKP8KXPE3FywexmgC1gnyoR
eu7h1n4U2zidrFGIXTYNsJwcrtdwk/22FJCBmcWcrn+6d8SUi2v9vSkDulSA
uTY4G6UfaGA5G3Fdwrc7RCYU29V5l07BGXOV0jki5S14lZXc1Rb2uFwRd7bz
+jz+LmLngkJyAhNz4JGkz1q8fORqqrX4cvDcYk+55wna89ZAy5f9P9nBv//0
gKHw3SWKokyxO0Y6vGq3dCEd/uIFJes3y2Jchc2YwR9i7BaSqu6ULiThlO7n
CmuUMF9OCWNKr6kZ5SHmv/N13iBsJdy7mp4pEJDmwiPiUDM7TDhPMzn0MJME
wUiglNgwI3cGgtN4L7wTupl1vDtx3fcIX5pbs9X+p2rVAiAm2jZxdyFz13Jo
WBK28PwjAckuMLxbK3c6M1v2v6Kd9T19NI+kbS2QLWw/HvQrEIprop8vl8AS
iLUbmElsn9u7bKuijtWKkjHjiKGP+2dqFMqqXUM+Lz8Jw6vVD7bO0wySI6Z4
aNRFfbQlBKWxgetGUZ1KYWnAW9M8v2FHj8V0c1LitCTX1wJSVE7t2nxNZrnp
ZzZFp1L6AZa7T6L6z66Bhdtg9u6YfSfTFNAb8tgx7wIzm/IzBcV+mr7MNNKM
6LqUbg/Pr+KtF8OOvskvG64o7ZYx72sffDbkvVU3QsGZTYFAH+jX1pnOxe/K
HEfLEylDXvFrcyUd11LOiRczGxR0ZC4nUBSRlS/wyC9chuPIu7bd3oge3tdW
sfv4dXrKjKqbDkfVK+jqepQKkPlcmtiGZhzWu7pEIbS4daAJJ57T5lpIsAIz
E9CQvvnZ90fStrtD7RakWJkRsDovIaj7Fm127zIWdObzZdDl3JNKcoBMSiC+
W9Bs6DgBJaACP6Cdkl+cl2UIUMCrLH/4ricuzWLpZ8dzefyP2CGJoNP0oITA
e6zSJkX4BxPGmXSnUPotmvNHzyfy0HT8T4heIqOL/aRz/0OMOSxM0udiqQiZ
tkGVy3qm3BeA1jlO3jB3ch8HuTUNOKZ4sOVxCEiI84ncRSx4LzZFOBkPBqnP
0PCsfl1SxcalNjkoIX9VZ0T7kPFgwMCkQv0o0Y1YZIx1qIzRROO8v/ur7fOJ
e6ySLsbHOt8tkdQ7DoK9goW0kvdxx/1g0BDfqXZ6Oa2JUoqNryrvxkRdudBI
YDEgrcbgZwAASwUDWWQvCCInF5rS92fLF5tntqtMCDgJLVziMtX1IaG1x0Hv
lQS+OisR5bbZoOoZiYpTIVbMLPhH5idwh2sP9hhzXnzoAzzTl1eN6oZex7Kh
T5CIfzfoukrdhvww7jlDxojbgMMKTWMIr2mFW5YGssWqz0XmBRm1qVHWdYkv
NE6tJnCnsdOj7QWfGAaX/ihfSd2DX/ovcg8+qqTUi+3kcOLVSwRf/pat4/k7
XnUdoIDsc+ZDh1zM6ySzm5WIsnC8qElfKmErTI8NBKqm0pr+pKD1Kofkp3kY
GGUF3l0hyLvRQMER6pv9D7H2Vq5HHTCt8QaRoIkxEQd0H+LD/XDs77lepskZ
wZxt0uDCll19UL8v0ryTJj+23Qgyn2iyXZPsw1+SKS323EfbAczS4yLJBnHn
u4sf5nojS3tsAnuMeIYv3C96y5iMg4xEfCyYhGlZgNs7kLqnVdRc9aV0hurG
JHWaUs6qzV5mf+cpJzaVfUZ0Jp4T/Rmrfzv796CTlcczyLcfpWi0VOQP+c6Q
+NI3FSXY4gPHZk/D7Bo+DKCMruKWJ6fOoqaqAYSnMWj2YxQhmEGKGIZnIoqQ
B3skFvcuLQwKPf6KgglrnR9Ybn3OqQrswXnugnLqvOn0oR+z3Meu7oaFd5Jn
y2f+nrcGvoDsQqvgBapvg7w3Pte6Jaszlnr/drPXvfB4iQIsMHw367kGylg9
rXrVHTp5VhMYR0uqMnRNVwUVLfkRaNAEioGiX/68mDvvXe3NIg9Co0K+zt8s
TkkFrhVKTLg/q5jWznQSVCT52EoOqZwVjoVH7uNwch5N0WqAeTfvfZ6RHgEI
lxqqUVct1qwvQrKFRLxF9lnU93OBvpkthd7PxpYhE1E16dHNZ30n6haE1pSu
pyOgD97iHqJCneXU/qJX3Axovr3UzhRWKs5gln0eH6CBJ3/vk6iceIfWpGL9
9VLAWJOcTS5MgzkTYv5641NXFnuapZNTIIo51kt1FiU++rQHgS1utyMYwNu/
2hpOUggec6YQVwa/oAm3iiXq6+kbA2JXlLH/Vn+CqlWExhSn0eg4LA713i+B
GYpoYXkx7FzzW/NfMgov1LQobXCZr9+QB868DG/M1529EYnISXtkbdowQaDs
NolhVcPf1njCAUSTLPJQR7+BxdbP/hZve0UjEfrWATMIbCKdDoopZj7t+hv7
K1a3q7eiTqD8TWwPrxun2ym8CY+5BebBIHD4NsSXFtTkXQNS2QxpzrRoxlfU
JAcmjy+zlhvhlPxlOvJ7JfUy/xFYQnB7+/8JgGR6XF6Y7upV9XWn4+dsK/TL
XrixtWS+0T8NDs5z41jSV2f5zP/j/fDTvRztJ5EmzvRPcVWH4qZ+GRq+13x3
AsivoGi18ja4pyxrbVcrCDRUnbm56YIEsd4cD0Cv0DdU05fNXzzLMsXNZGea
TqKKTCK2Fk4n4eGAKCYAt4JJHWTjrt1YIzvDXjYqt2PIA11TGXogfLpO0CGV
mp2gQUc5JlcB9c28curXa551xZZPIZZeMawrpy+LenCFJVr4WjcxfnJ3GsdR
HJj8LwxrSZjzIxhJ9Ats1diGwhJ/6Qikua/kQDif/tmShDVcXkaZ20f6V//o
i6NqCVML6USRZMZ/p7dc1mbbVXAZOwoL+nOlQzM9sbxWmXAIfH9LYB0p0ydu
Mfc7JyPFpArQTt0+AWRGjGhUOgc7QU4T7fvS41jy/7x24JiTiESVuOmCSpar
fN1YGYa6qR+DqMLebzCY1nGbEt37ap5mkLlwIFWnSLToe4e+OtxkcHVQfZQi
svXGXRekgnvE1lg9fW1e9lTaP/PC06SYdmRw1NN4Pq1IaUlXnJQCdpZLhs+c
VdWnazsrREzGWJuUKbLSdtFdcxZx9JFdjZaPW5GO3pWqKXvUmQEtOcTDJnBy
tf1HjiUGtrZ3+zt98x6rnTsEg+IhEjD+19fh3mh5RQ+wiY0geN1uTV5OlqFu
tCw6o0icdTl6+3tpzJLUuU6EookQHvJhpPr6SAui+sPBxXNcq9eYWWOr8RUg
3kyWEctdkLZoHDIgKHBlM/sELCptFVs0o9lgC6XafDZ6Mo+3UyYDUQXKMEML
K4BvdCmZ1yI3Vpwef45Z1cA6uFLlOrRUEACiapXHR4/+8QuaUnUvNb0LPIEM
QlCvX+jZSeUIkIRn59UQ9paXMPhbxYWvdP7Fy5KejeBM9tbQNILYDoOJjSfW
52VNifSERolwFJL2vHDi9gYcLkTvS/3aZeikMM3YozU0aPGbC1HzBXXI4dPs
KMegxDJf6KDFE+bqlSl2PzY6pgt4EUjnkhYlFFBSJi4WgoyJK2xSD+SVXN1+
Pc/JmLyIsRIH7mtmcADRb+wyIdKG1DmlJ2YmLU3SVU1R26fzHK+8SxsIMCGO
ujJbN4VAvqdd+PYYmvU2tGQnHMPEmXLGl0Ilj1NjKyslMSUjvSY9pKCVV/tg
8IwIYr/FyNA0JfuDqndnQrcqLnDEhLmFs4Hdx1r3U/SlFuYta6fNra5w0Hl5
+R43fWPSmVjd/sku2dYh4Ktt36GpXsl2a39+96usgUN/rlVkYM0IEkjFVALR
zh8/JOftykRUOttZjjiNonwNMB2x6hz5p2PTBj86zOZI+EhkwhAyKCx+Fgz6
gIblh0w1BG+0zQyGdWIQLVUgADVJQOFhnsLy8RkqbQZMMGPqJI3H9ceTCYBU
+mudFIw7qUZC6MQoj7neSUP8+86qRKfcVUE7nbz257z1d/eVSBy1jcSPyW4G
1J7eWNz4n2DzCG3fi5EB9ecawmjGnClT0R7eiPoykq85p4RaEesaO2PS0ZHl
4fvwS0ljp096eI+HwrLU7fAUmUI/xcHY1mIeDBhA5OQpufW8hfy3h3J6ZftK
Nqqq8hz2OxC3V80ai5huguBxuROlbRqvEzuGzJ23YVRpbsznaCd5ApQKwXZ5
sBVMEzFO6lonbMy/jd35EWwLJkY/Wzuuc0pHgRlKv/IpjgynOmqO9Uo8XxRy
VtB0wPV1yR0RgRDMhs9JMKyQJhoTos/rBSvsgvZ0tZ7f9Jly98nT+utdkKhp
vkxH5EU4a+8UqvAD/tsIKJKqWCR8H5+mrpMlIdZUEgMV09/+rWO/JlNjp8xd
4SHsEWl6wc2hXeB/WkSQyV81hLBS+5UFndTSBGvS3iCcONHdf1KDykkraIRy
aZtOO1rzoWjlBfD8VXy5ZEubJ1yZ18Lqz58U7iqgJuPLGNdUGGhyURqTji5O
Stu7KFh4tt1raNrBZi7cKAqgDtQN3FpEHVGgl1ChK6VxeRzCWmRN8GFkb3sl
xyaDI3EX+bx4tVRYnabX7ZtJQK1IpB+A0JdcLh5uRyrYUm0vrgvtQLuuKacM
AyfMIk0bngP/tx1+8PKe2V+CMa1xUxVMxIWSxoyCdmek+az3UDtCxXuctNqz
o+Ps1mcOKa7zkm3ljkIIutgOamI9CQ5D5NvNTpMOVpj+JJjZfiuJ9RY6F4gI
fj2HnDBm8/ViuOqHlFBskB+VumgrNGMBFt+zwDv7b6AfMy2vAqzMJOHq1vbr
xrdRHCqvBwuc3uNezpLDmRw4Qcaw9zwlefCTQ7igVtfqqEM8/CJ6W1RpqK3a
Ndk+yxT7QMJxtu6/knGuL+HYph1sCgqIwHFpHB56rtWaARDqIOBLNsgMU+2u
KtHnD7Qd7EhC1Fhb1d05PDqyBirFgwNoxCnmfHdzOG5LOz8GdzAxo+kHGt6B
SNMgJ49o6o57EoS7hTlTFji0SMvnTrsqgAR0RhGeS/Rfv0QFSswJGX95H9YJ
ui/G/wU7OYZd+5QcCUl02cyhgdAcrrhAt1y1C3obufr7gGEX2ig0vYNDli4E
O5hQuHpI56HYdHn+TEX+rSmYjVL40lmjMWPjGgCfCgez5Acw+iTLAhsPX3rq
tt9bNheJPP6yEJQ8MtG9ofSpHuGSw0m9DGpfI0fangi5lc9aT4i7goRw6+z/
uoG0a74tM31hvu8fF5eDAq/wHGJG87hr9ScU4hn4eHw7rngGJmmk39MlTMwr
BMqgfNdNGvicebTMq3IGQyp/H7KEDQZxbQufoaJBETq37e2r9tKdQDFhBhNS
cSFwfSI8Ks9iNQRKglaF96LytQmmQN+Zgs5NklkoU4ILzWiS1yUgtdswR7gQ
14Js8P2oQQTiI+gN1kL/P5FlGNMcx+atYTRmM1K2YxI+BxOOyv8zw/bKmBHq
t9pazo31vy34jbw96ja2ix5kQRhYeoPyBTRkun+vzC4diPLoT8z2D+HNMTIv
Ul1PJj2aokL2qf3GbYGiK4LUGBybvXDFC6tdtX209dP4vacOuoSFCfKA3dd2
53PNpYDznP+2KtfYy3dXJaM1SZTBR1uTxyhiYCLoagu5kyO4MCY1PgMdFucc
+L+jaZM21TwGll8m7X/7OhHGVNTJ4arY6uFI0GTGlhHkGO0UilOxXs3Kii+A
oDZyoDO8ivSU87joYXKdEfOl7got5IZ6uMc6Fh1RRf1Nc+nF9TW0YtiOWJt1
3AdNOFIO0Eua/VofsqcEGqZQ3d5tDMH4yXDLYkoBayvhbYtHPtFmeEpIVsTo
r7xSf6N3Dp4soUrj8d8riYrw6Z+ncdlvKCv4eBXFn0CScKACrzHcnqFCGNbB
B1B7086vLEUdWhTkN3iKZ7BG+llMoLJT7BMzCKwuPHXuZLSFB/Dk7ji7dqht
v0AH+ZTnBphMyVtZJa37kNbUv01NBysRUgtXZ35rzL2ic6KTEvDoU5+DA2bK
SybSAsWzzQIy4PgmSqmK5vBB079RPJmdT1osIm5QzuZcnBI6ddbCp5Km10Vg
f2KX5xUSLpJjpAxu9Ngau1POjkShP9n9whevpinWkhCWjbGNU0Jac4/rohfx
5ZNs8400ixKnoSbG7sZJRP/az3raQgp/9IARX8icI8zK/lAyOhBevNtRbGPa
1LT1m8DhmVyQ/Eu5ltYIyZ056vSjVpjbrp6AWZedjfMx/5l/jpXXUSFE+uwJ
751bEv+EYIvEdiGQD49D+PHkDT+xg8aUA1eLFCJ9YT2doXK7oFs6tEKJiCLs
EM+xuCXYPLSnYsTexWzpJRviPKc9d3DwNz+qJ6d3aHfVA1QETamimkOnRazh
zDE4DGzDzVDia4ktpJYpFCinRKpwMb17Ml2Z2TILelczM/1dsYnJTi6AZ4Pl
fnZOvXxBn8ygT3FDSAjnX17Kl1hBTwwDWuCL3oJ1JRDAv5W+ysJ/DiOvdX8Y
6UfA3jNCTx67Gy9MQRF22NKo+ktdz8t5x85QbTMfROjPEWbbbwV3r7mWboai
Ixqeq+qzKj38hiW7GHMD5YDGxZBi3N1zapRihzyrGbC7aF3AIBvA0nkZoFbN
t4NbJoHZoGE+oWUm0bgvsJAYo4QEHA8ZbAgtg42ApMjCttXLBX1Qkeqzp2rz
g6ZW4noi7PM7UXtEcBW6XmzXRlXduCYHipC0ofxn2Kl6Kh3O7CLqfNNyH1Gu
cZg8Y9MzkSvGx2ntp86qBh8r2uRsuAQGEi6rR2ch7OsKN0HJZa+yPamI7KcA
8MKSN/dcwy4AVVfNivhoNCEjkKvkKqHYYZ/baQVyvB67Fl5JW9pvPaNCn5I+
EQZQNxALAJXhKI35mlnOR6gL/3grGfY3ppKs4Zpg/aAiSCayar+sj15QluRZ
M7b2eNg4h2AcDpOyHUqVK5NfaAPyGiYJ99T8flP1PGsqYg0mVW+aZ09XSL7q
7ykD0Aq+JkAn1HIRn5nHVx8odMB0Kjkrof6sprWEYFG8jDloo1NUUaWEHULl
1b8t8nRAY3pL3S0WXVX3z8fe5q24lukmxe7qNoOSTd/GewjqRCxzFlXP5sMx
5obxz0UO1AaUJrJdwl/7j60Opepw0Wx1V+J2N0fd5R8auXoN35AE+AmJY20i
bjH7NS9oaEfMlxFYWmPXrwEo7u9YESibyWMc8ZIT17YKkAEjLPduxtH93+PJ
CkFjmzKSoioVGUZ29+Ci5RUYGhoCEkkwYQZh3h+gsaK6Y45TPU9A4iFxxoRY
sgpqRmwjrruZ1udo1XlkrrhuKpGF9IPPi3/v/F6MZKoAaFoSVo4cvf05+s5v
xuRgcexR+Qud75GjWhn2fYDMymKVDMnhVo26zYelWEXJRzhayJ31mng05XZ0
ePss4lpl/8uf0hfyM9zjFAKt+GdFeJoXgO8ilGoczX2IP0e8TXSXbGY5fX1n
9boAShhFEV5wuvE7dvvQXDqnAbzcg1yZvlowt0F641p1a7OdLZV6+P/unDv6
J6DRmN/qvrfY2fpn9s2m7/X7ylzwSwj3qNHO5bBYuhWm3/F27Zbxg7H4uKHR
RJJQ7xZZMv/0jvUtjvBC/FPeZG8nKz+0BwipE/PuEsprYZEfE9cVPqzy6Wfl
8PY7eEUKv0suYVWehdLyBLSid6oTYhn9/zyUr3+HEdwL1X0OBLkqZvaU/yen
3dVX2MA33rab81qEfneEgUqlcEinY9yrNlRUz/V0GryXWDdmuibRsQvYSd9+
UwD7ZwR53uDYlq0m8WRnAazyjCt3lLnjVYyrzMNzX5L3Yx8lNOh6HxwxLA8P
VqGskp/w+b2mjGPOHpWa+/OdrvY17qsU7tIptVr1dj9Ua/sn1YSeifWb0MJY
7hvB5D0EtQzNU7vH4LRTUXyxE3ltUjTgovESejkbPzwIO0u05qn8swa5k6IR
KcwZNp1YmhefhqdqNwl6MZ76k3W2zKnMFYM0pxVJYv0bgjijiVzOnc6DZC9R
WIM2GvEEWuAjDoa+OdXtHKTSYTsy7QgOULsq+vrJE9GvjishzaMqtEpAnF9T
Q037KPlfV5AVn8Jlphhr28deTBX+DUJpUXddwL/1LADBDXTJieZ3EJirDTHm
/LYET/wOYi2n/BdDDYqMPSGcCk1afp+8IvXi5LMpcneOmoOne4TLfIlVImLb
Puszq7go29lG2Iexr3Ffyiebw2kTifxjc5ZXm5I7gcdSYbrnGvqLd0D4LBlA
OMA4c3tEMyL427WUEmJN5IwiPEY3UzsQUPfR09GdBf28X/EuDVmIaP9l+13s
gZVj9IbLdmroFSvLUCQ6+ZK/qHRqUbeVVVHzS5B+o5Hanc6xsA9H6Uj/C0aM
aOUqtpC1WsssHZhul6Wbi0kDPVuwNzzUuErB78k9doG1XyNpjrkGHUTDuMjG
lGv+i76nrxQOGysJLGfWWYb9x5FhIo1KEv0lKziHI0Hz87XcPrNJe9VgjuA5
MrafI+WLN+9lBeNdGNL6tkKMYFbg8sB8UTmUNBaiXT3RRCyFQzvqztWCEh9V
aSv08+btQUXhSqep8oX9KP02IJpovbAHDVpgNypoxC/Hx+US3zCIN5P5iwnK
lxw05xB1oQouJhDwIAyR7CFpEX+6s3fC64r84zUQ7NOblh/kwoiW0n+ko02n
MpyIY5DDJ6pWi1o86/5NemGNtPiC0cNhaZF3z1EGIDRqi+khKwyKl+5Gci6T
ob2z2x7ekel5qRrb5ZzeIfIXUHI/QaSS71L4nHSHNQnk/hE1FEzStaFL+PNO
98YhUmSDft5sK06HzgCUfpR/8RXVb0l6RnNs4MmrQAr5HQ8OxJ/3T2w7MmG4
uX4VXwRYRmP1HhNfrcvNftx3EaSFrqbvGFNL3LHslvqA8gc02mZXjQF5TAo1
viFNO5//+YY03x/MZ+iOAsk2PonVQw6tfimLIWw0+okhPS1p64HDtYmUTaDw
M7sKMzwvvMxtRughubKj8II8tnNLFUUheuyCEt+UQTcuFQca8Eb579R4zIJf
G9KtsqMjqVBCNcRn3qQZDu/nvT6RKVzDidq7zOgJzXRPhZZVMngmKav34SAB
FGfoVg7zx+XhX/Q+R3yWG01R1fElSuHAEY5vkVibXbugH+1sGIWcBt/G5a7X
hO4RI44MZGQILtvCGJJgq0HoBzfqDaRDw4E0zfalAwWTAH22ooydJoYFrvvX
zUiuOS8nM/nPWSxPFu5kxxNvY6gVJpKZ/ql1kNL09DB9W99/hJumHdOkoRp1
cEkxGcIDM+SvlAcI8HtPNPYECbMnWOyhv/Straoo3HyHJU1um8fN9ip8t3XP
n1EiS8PZK1mx8/g2sNtrcBH0pyH74F5fcIInk1B8HfabadCQK2NxTY38hyqv
LLuiMbd9toQYTmp6Ij9Q4kVu7dzmxNBmFgIojZcNaUhkvw7WnqBOfq/8CsqJ
UynnkvNG+6XGHHXCnk0Gd52BLEdo22Ze/6ja9bFMChWlZB6oY0hzQs4Rh6h6
BXDs2hBiQqEaEJhXaOorjLQF3EM7bXxzggeO00nczuKiZEiQSHHNXpgYwLmQ
ZvzTiYTYPqiCE2LkWckVyP8SW/SOPDCAQ3iVNh01zRT2o25hTUrcxiXu8Q3k
ZAEGL98mcfTH/cqC0r5gNKbwA5fvG/4bjA62/HUkW1aEbXYHCepRPjeth4dS
zsvzsk9mifMPQhb55Dp9ypCBljCFgUIwTJh+PtQX0hR02yiy8H4PhyGOT0uZ
X0mmBbAjQmPjdLr/3IqzBBmXrzX19xGBgUGkWGAVI8U7xchUB7uXa4uu1qKh
Pg+pGs4qRbyFUdxpz5tWihp9X/ENP0SLjLmUuD/QQBrWft8PUbUxTSr6IqBQ
hKQd9tsc2yQpMrp3rQL4Nsllil8NsTY9l7rw8TKyfMKVIu/HqjSXgM2s+QfN
Slj7APCiJROnqGZJy4G6fMFSqkNA0xL8g6179IGKTBC5yVOLtxka3mLJ+o4e
De1+UiB3H4IgQAWpDbhXuHh5MTWH2F49Q+KBmD4ZtYaaqE4ClFaE77JvmfSA
zhvoQIE+Lhro4C3InhPicCusNRH5cutfpttyUWttIm+GEo4OIK2mNC/gi23+
m2WdNVDkrlGUsxfPo1+WCjejT/2WARy09cYH30335L6GW6XVBh8+598AeOeB
Cwow/d5miTzoYlEbYIKABnncf6kot3jAsBdM9S+Ou9tAr1B330fYjdI9LTiG
nKVoEjeAG9XakdnN0wvxOnxDpoqpwELAmnlTp5h5Jty7UeMgfsntJx7dWxMV
fx+Jir7HQFj2T445oAYCvXmUtS+6M918IEWMEP3DO8JAozuo9HV/xSD40wF+
C4rkqHhMo8Y2xVJ9oV2yKnaFR+MEUTXZBuI3zjiNtDnvjYF3a6Dl/W5jFy3l
8CV2U1Civ3LU9uwGqfWqQvirfQ0K/4tWLktnz3VLoMtPVp6kA5n/uGotllTO
3n3ayLgBsayRXU4Meyh1UYuzbEZ2FWJNj3hSO1tsuyZJL8fpqTbvY7Cc2RtR
hFaT0tNqm0p04BYU/sWf3nYjNCaxy91siI5qHzRm+73paaVu1ocTAP8x6tCC
rXef2CZ9m8zDufrekkZI7s/1n+vqKvgO4fxpS6eTzNDGuYwtLh31jI0vHlBO
sGRuXljZPm8zQFbMseu7G+GWanVwJILVDNw2XtecDAAD3GrnhCogCABzurtx
uA6K9eoLDxe9B2azavH+oc7cKOgsyRPS4viAaVTm9ZY/RTuPg9dbDc9gUqGB
QmCHS8EolyBlt2wzcBdm3KHf/7VibO722QEVMyQOXiUd7/4S5M88w6QZ0rvY
tX/r9Md/o0A0JLot84CqaSk4lVdB0+CdMnI1TUJUtdEVkp/qWy0uF1xqUf2W
JPdGO8RWMfZ4gpgtIUoVls1hqD2m7+Hc4cYZf2DWOMbztXQrS34508CgDRC6
53bEHlIGA95mRai7XI+oYkMJfwtcx1pwu0ypzOdaPryDKmVrOlyLrE3z4tSd
Z2WTO7PURaw01LRq/aZ8URETRzmLBT2B8Sx3BtX4oVwid/4ySqyt5w9c9pwS
oIm5ccG9K2bEsP+MCGVGamhBCmKhHwtP+RvwSFPIHxU7uVb0AW30xfQMq/x9
JSe9q1Rb+D4sCylGkIWbBUBLjUxMtlT0MDZfMMNECLnbHIi1gW/Cv5RYiiiN
WudiU0tSzszGrTE3dnVGxmaYnQRZqKsJObKHF8BB184Bt3ti9nKBMSU+eDfo
3WFYJchQQYHQsY9a8xa1KnWRBqTJIWFiF8SAsXpGOos2l2+T47qnQ0OnICtH
I2ehlk3V7t4WGOk+lbc7c9siQpmFugHgwnOYCYaWFdFR0Qhc5fg5gkR/Ft6I
Suy9TscM7Om5oRzej8RezDXPKN0kS1+LG7NuYTRYRBkBeiokjV2UaT873Eal
W0b5agoGQDcXG5of4IolqFk0iShuyIJ8WGFIREEkddFfg6qZW2UYjQYBmJ7b
dlTcUWypVvSPe12NgCa5rX0/EyOYqt+KN5AdiDxaO0MuqSkM94IfpPo2KVXg
s8zJOckdrErdYEqP1JaLawOctfkx1M0nQHP8MD880zSvDj0t/mMPf3r7Npol
0LqAv8xaggeRNfPypv8ruGb5q3B4jDv0g6OcUAYH+bVDAE2DknD5KB04VXRJ
XXPqpC7a3XjQh0Uui8uN09PT9SDOuqDNmkjTdVM39FIbwS5IxiyD0+CQ//F2
s3T0eOAQg6IDD8GUdEhQ44zOod5EPw/Hp5YQqA2KDEgXOIgI8jv5BvD2AJar
jye39WZdpl10qITcfMUSlkGHj6Yc3AQFO5p3inMvyQL5Ut9if+fmN/zTErvV
B9btHtPl1BK+AnKXyz7MHZ8XPlXc/2XTOMwv+IlxZTLiC92uWUFh2MGVGmFe
zNQQWNsmPt0c5OJhxTIL+o7Ni6LzDgKUsk52yd+Ap0SMMAph7gB5kJ0+609I
9o5LTvk025vyitaefXPKp3BFyn2FJxovWyJqLKLFObmwpUPtEPW60DdEw1rM
QPLP2btuScqJZ5YNjeyEbHmhm4Y6bYGKHQDxdQtN29S0VCxyePNiXRkZ0mZH
8oN3YyEOH4KT21BSDPRQNa2M2ocd730AMQdOzLIaCOIjQJGKUbKB6Rew6qOF
HRkCssU3Qxgc9TUPI2zhJmZA83CdF0CL/6fs3GY1sdjSH9B03VqzE3fMPAaI
4fRW1nzboB/8oLAei3qHI13Cuc0CETZuUE96MrutZOGj7mlxgP2odj0ox2mx
ESLT1PDE3Vke6kSF/aiedjgsoDk6XNvnWcNg5rZbuo3ByIVLDVZKUkyc64t8
phw6yEN5/5x7bkRzoU7Ozg5MqlZaJUBdtIlB7oYIZHbp2hZgqRWGa83sr1UU
b4j3kJWaXkmQFZ+XCpP8eoWE2VSOPON6ZTivahVoQ1Fx03WqyXK4o984gp+6
6yjHrXIq4Ej/RThnSzvI9wEUAFoe9yqxeJst8KhHaQ+uah/zu0jvAJDAf1xl
V/9mAtf8ursAcGm5CuaFY7AkldngarHjeOecKsgbDQkGmqqLpuis/XJFp/zh
gqz1IUlCxP5bgDhMuqtWsLjuLcCcl9IybbCDgjBLzBLaG1Hxz7yxQ9BLSNRm
i3/Nh7MUShtK9EjWVyFJqVDSm7R2vc0hkg/3dkPc8N/AWA8zhno84IwIyT6C
96qG3Ofq0loYCYz1BekBaSI/NB2GABXg5JJrKWHSV1AE9Fr0dR8P7l312Qk2
cTIX0SCVNrbnku2MEo/B3Pr+yjlu4YD7+8gV68EoauPM9gKbAC3wNUeOEJZ8
fJt6MfKUmpH1mxwEeV1AalJzXX2xMJeO396AozEfXsIDLRI0SkA5e0nMFF9b
0owM5+jn0wuxSKw4pq7qjYrSZE1R9ZpQcRgdPXzfA/TqyyK69MnIZnURkR+V
Jk0UrvjsAO7lrfCfYxIs1Q6nuGxPi1b6pe2N7uXqlVG8Ba6u6Ymrf6HE8L63
ACK9V0IaJn8wHcfFp4B+FWiyc7gV4LIpJXHDZo+NG65rrsroe1giq/HxtblP
qUph7g1nIHTsxxK1ng+hGTrVxUZrZZoivmvxSLBIcFtUkIi+5A8rfkwVL+1D
60Y1wRiv2UrU4ckjFkDtEq1eLOq62Tnl1wkZFyhbEAqqnxuE6QRxwLZYRw7q
s50YJRrk1EBeggCSAH39mPuZHoSfUz+BaahAAPLCC+tA1IQZSPrZfKrfFJF1
CWBbd5iUclyKzQkF5OTxY38B8pbZkhlzTi5O5KxsRAWPPCwejSUn7s8guGE/
XXVx5rqEsSstVoVK9GNMAJWsczKSQ3WIWbYiY2bGtl0NQrz9qiZ4BgQyKQFc
+R+yeI4THhkj2TDTva1NQ6IHaxUTaJo9HB2o/y7sklip+j/Cb8Hq9h5xbs/Q
w7xECLGnsSiu9CGU2NaHvBzEgC0V4L0p5dxvF/Yp/BgNAV43BsnT6qbD6n+3
vM+xreoTvk3WGgbimUrM3a1U3QDiPI6VEizxnmw/HG5MBHUZtQvrh0uhuDDO
SRU956oSRWu18ZiYwAIr4yNdX63SZm0m0OjgdbYbf8KMv+CBHnqFf14u90sS
c4TsnV9mOpfT1LiZ2oAGu00ogIPu0UzjtSJes/Ng3n80FTL+jv+mP2H1IHJn
Asc3MHbjLFs5fCx9bX6BqrNf1tI+mlr4QjoDBtwdvign8BVd4Hou+b75UtaI
pHMPmmczRalGcxL1i2kPZViq/MFhd46A+gNy3OcADvcyTSa3mOVezUNL+Zc/
t1Y6fai6am30TBu6vNaDOig5BJ6fhXRLGur415i3CRa812MWs0zuXLpPRsIP
Sa6GiAT07HBMKuFMf2uY7IgFVH2QixVfzr1U2HkuUIWbe4V8t4sT7W2knntu
fCcBR+Z67rww9LeksqqRjjBBB73y0V2ShEI9Hgl7J5SVw4F/sTYzHZz7K/71
bUaAV4fJMVUSC/88TUhhX0pgOT7aV68rH9p/DCH2ogvFKEUqK0oAP+Uxk0b/
QDAXf6navPWW26FVs3Qb3qugIGsN+yinLFHkcfZSRuqFIR8OSkF9xV29YxLX
ZrmQHhDJYGkKRZtMjP5+qKNxm1qyaKdbCd5iEDjXyQYLJAOMWM13dK7BBqwz
DXHVz1cZLslMrfcuJ3wAsZ4nf7oQjEuTLPGu/tA/lXCsA+ggxgd3vT54TRfY
oxZDjH/Q5hcroJZ2WupSmYlaKGG98f0EOwHXHazvMPPsy7/BBAU4YfS2kjpN
4Adsh0P9pQQ566aVq+AbqtPQA6Ovh2CerO+D+NDPohzQWwNI6xacJ5wyEI+7
+oYqzcAJc9+PTJfB1dnsLDQgDctI9PQW1iZStBbRtecwAGK4GSiGySbM2/kv
/np1fp8cDMPpnVj46azUm4envVnCn2NNNboDIU87GP39DQn/7ApsDO6QHA6U
3v2deOO0xJJN5lcxEfcB4F7MiJVnVgD/L+E0X/s4blm0hjCWFSi2yn20nL8Q
suELb2TGPhhE4ZFTgIBzgC5tUaG8xfUn8fpu2Laaw0eXudoSc/ONdotOOxlk
q8p8/+rv4pJhODww9/jUv/6mtDmxh1LbKf1hsCyTQIjHRDbfXmzL7SGv8qZb
Iiwsqo296tVBA+DSScFQG2YYNciZgLEiUu7zn/tlV+oFydonbXLyEo5iYSLd
RxIyk7k7os0IOsxfw46nz+waI/qZOXp1JLxscR0OVWFlNsG3v67qBH5QluV6
yWESV4+H9QheiSkmqxd//vRxREf+dqZ/S4NImJy2qNurRgVJRhoUGwjKKQSY
DxxNJ7KC/MEJhCzHoQcVadbLa4Sih0WiReTgpb6fmzuaIg3k/TMjjVHtXDbA
5oWcTy54lwhjsx6fupOyK0S9hTMJc54g02QmtEQc/hE59IkNwx9BOIoEvm4S
qVpUgXNGKs5nbsJtOG7Hyc2YsI0sfBbdtEHpGwXhIQGiuszrHCPU1FyzGLC8
VMbVluYlQ0tz0DDo3p57HuIvo1dwVvy3PRSVvKOgeSxF7PJ3jMwIn1mMsy98
DGW2ZOWI4+YqSkIWuHmo229eL5p56RruCF6ZR0b33yNOUHFsTRj9n07JcfIF
sP4nOsxMaRwFyCycXs1KIc0B0jDiAEesvPfNZiX48D5XmefROiNb/Qykd2GU
Qy+jMI5AQYkNrz3ejs93UXELsmTMoG2iS6fezx3vaPfy1t4EHp3PihtV3A+7
eRjz/hZcoPd78FYXkEWsR8fcrnB3ZlHY26dJovQElTAPqlPwOIgeCag5ghi0
e8hh1oaNcxIz0sfswtXc5FF8g3WCqVvK09VknyLIoPTiTr6ET6BbkU3khWkF
hsKgChajqvEsW0BOWzWeEBI29JdqylTQJugVdupKgVYCePOI17cJFK3uplM7
bYvzVul7+HB7TMkTE/XcK+uEnB4PGQccSjvI9aJzh91qMDZTj/Mw+Th3aST2
twhTN/Co/K2dBzbO0s+zkyxX+ziA6ofX0+6ur3kRFDYL9lbdpQVcpVnhtD+k
lgq0B4qE3knTq9spGMkctwlCKddotqNGHy5QRwdqvtvInR9zOKmPp8taZ0FW
VC5UsSQAE5/DnWQ17U3B0ctmpV4T9iifN6PUWd1GcDyvK9wRBZQLHsLEsyIg
IT/G9/3F3EePWmrKWHzG2jnYKFZh4kNKLyyJHBSyfbyWU3wTyA5vSgTHwzEm
3GkCgHN4CWM7dp2tL8TUZ7Nhu1KR5s3cVBVsZqKxrIzK4BLyrx6nBgEa7O/4
WR1Aiyi4yJNgPsGFWIVWw6DfJ1LfJ+ML9QoRk7/Xi3jSurEWEgbEulWJEoGa
P+SD7Kb2/TiwVzAUfqzpsJdD3qBOBd9yH5So/shLa77O5IsM3tLmBRUZVyyL
M6aFYm+dCgRGk1xs6TGfDMCeHOgg5+IO4UNu1gGcFh30bZjwRr4Ioj3cKsl4
13JkC7AEoIMwmeG3TTyMiGWYQdZjZBesZVdCUzL7zgUgjvuDUQp0W8Ec6wXA
NRTS6MenpE0ZOqmdX/mgMOXStO97cYi6Xku2DDec6Gjh1jRQbjkTGJsoBkif
mhznSRvjIfLvkLs2NKQJEdqYw5yWl+YggGLn21xCR4qdNeLS9GVTJ7y4C+U7
X8epDSPH5UFOqGEM5empLeETJ1wYnowSrDs1MdYVVVekuXw+Emfuagydy8UO
CmZFc+SffjAsQr6GzGxtRRQUZGyRWuYxEmdtcDV7wIcGVpuq2BQeUTTGjVeY
KiVQ7dY2qymHlqa+tlCZqgfDlNFfdSw0VrknlGnRJ7jYCClBawwgMwlD0QPC
N4/ZRNVDiq9NuyUQQqIFKv3o1Lv4P4JKUjf4uUbk05cCh5kfw+5pivEFqDNo
4tb9O1b4Ml2iniIckzE+f1QisymjfqG5VY2uAO++NElVr4jzg2h7pM4HduKm
Xqeaf7Rc7d0fCtX/IEh4ONZOfRUuLE6edzKsRQHeagzTc35kGisBxIGgnYKp
NSvVXHrWp6h36IZAaUNor3oMIt4BDoAAc5NI7I7q6KFzs+zG9xhLDQU1V6jn
eRGGTywTcvLlFaQXDySIaeRIbcjcBpirh7MXyOLCW9hYZVzmldhmRq7raHWD
5TghLqH1snl7hmgcwYs/eVAiLojHv+6L1JxPq2RQShsjQBmXqKYdAuaiZQDB
w6HxleyRAGjjR3RYcKVSfPKgMC3nJ8thU1eCYaeiarwj7L4iU66z2b2Ai6eo
I8u1+DkAD49I6tjN4wzNqj58I6ru8G7y2q+bihhea6n8i3tzMCEeItu5NDZh
bYNgE2SNOixK6mx86FmrWpxj0XZSORqCMX57oxLH6GXyP1nVaVCjzs0+qrCT
/kpcODhagee+FTONupKJ8t27PO7rY014TMswbb3Dqi4oFVsK5lU8oTuDX8gy
D7pfObEy0R7q2LYQSOu83AYTOxDreN5n1bZh+Cf8B+Ig7IyyhKHavhotc01W
WficoRMZEBf+4wvG5zUOlRMavdzyCLupXs71/X7HHNDJzFwGmawSBg19Zf5E
nBg5fS73LA75qmfl9J0DDqnVCMwqfeTVPFze60skgfEy4MZXvGxU2gT+tpc/
r4CiSRhuqtuY3/+QJJcCm3sk8/3AuQtgNaGmvCDjUMPP+qXZWHK7LsBT8808
STEvZloqIfD0PEC0jn1HZnyrN59dcmOERi33CHriZQgnnlNVXvmKg5Q+i82K
qOy5GDcR209kjgelFEGbP6B3fdXl49pv/rLEw9Y9W3rvq+HkuTF5gSHeIneR
RCjp6rIUFc8wt0ZtmYXM/uBDn2A8EpVo9xqt9NvuwuFLsKo8Y8qnP00kyohA
Gh15bQGdqt9wLGH6e1bGyILGBx5m0gXcJotRTGTBU/Bg7N/4teKusp31dp7Z
s/bkIqi45aekDP2HDrhZ8/NdnBgz3D6GXggyniojm2up+UBdQ0A3RdYbvHMo
/lZcA3wsRsoCSeJ4hRGK5Dd1jacG+1INlO6cy0wS32ACNdOncXMkkir7p2TB
o95+vpPKzK2h1aEVB0H5s6YHhWnyte96kxVXOQTCytEz8mTT4ASM2zHaxhdl
5zGFNi1EiQxJkZWkZpfEtvaqDqV1nBXumHouex3WNonPrnQtBER25Xc4ZS3G
9y8PhekFTJG2QisdVbPPvhjCoJe/VUCKj1rGM1DByHJgZUFBLAYsY8EWh3So
yr3PqzRobnPmEW3F75q4ethmSXfinTQuw2HwUbsXx59GZvzEdlVZUUspALTI
sAr0elpGVrTaf+wJ93cFsbkmZkT5j+rxSTeGWsPHJqIk+cpusLZ1Yu0GP7YM
qTNDTU/N3aXQHtSnucgRbixkDO7UYebWREsnf0jpNd6y+kGynW9wbr2JyjM5
CsOSsrAwrf8kcdBJNFHMbsApzghvfTdOrTxjNGjXOrDb4ge7Eehvuq0p857M
Yg6Z+/AUj7PffOD3VrigJuJENYtGGslSxVaOOWzppZ/g+7weIMbjJ2OigjHL
ggM8KbFHOk3Y/QojxcDl/QOT//HqyDK3bIX6QMOdr9wKdGvqOss5DeKnCQ1J
mATW+oMp5RYkGuoQ6Ypki/h5Gwacw1gDhDGDLAWA9G4Uv/BhlHcRmj3YKXLj
24HI4tbtwrVkWvW/g4JjTUSzg+m2cTsZ6MWAuiVwtd1niXEp7mYcgSL5qzCK
wHozsGSn9VdxXf+Btdr3hDiEAkQxI+SbGLaJ31JJ6Ks0tV1upLBUDVlyJ0Aj
2jT73V0oXj7bwDsX1h0cLJdnmrpbfR2+6vz3u0bF/9jhcuJ7n7PDX3ymwoKF
RCg3tP8vvjY/2cYGHctMCTuFssFEuc3Aq+p+B1dqxT3hVU+WddOF5JYlW77W
Uwdr/7T+VO5xFOAUmgg1HGDXAHVHV+eTfz2xS5OT8f8jWhPy34AI2IJbFwSx
+et8t5sjKv9JT8ksCTqSiv+hely5F5Ala6/oyCMjIdQvDFB9CRTqTfVKRY9z
K/yN8bX/GGOzLgwWlhi1yRivafLNVTVXu8t2A35Z/wY04L0TlARFo9rDT2tU
HtsXrQfY9hmRD2UOHusvfh9Lt2GLIyj50Uj+S9vqeqGlDESxNzUTP0qgz94u
jNMjpgdX3fTlZ4zuxP6mgcrnTjQLTwUndAB2IkVkl66FmymatXKlffFMt0H1
1WUKQbl2piPbmsmpWtyJyjE2tHzIb+b/Z+K/oAASj4XKx9RkjQ1bLkOTdmCM
5KVYx4kaBlPRbkCYL+YeNgXO8KcRvcDNJ944mWpY+7nz/fepVSY/+QJRlP7t
tUtp3d8MMfxzj9hJerw1B9ITBLsm5gGR8vQAToGRHXCLGCAE3JT7YaKswBlj
DR4Bnm+dbfRHe+IKKUsealNjdNyhAIyoV30wHK9Wlej97vavQC4TPYOrCPHQ
LPDl4HFSezHPzkxvzOiOmgpp/mdqX3shNo0h5rfK2gevFwqTdDLbC/bdhiBQ
Z59Sa9L4d+slMCjY56FJzBSHoaDR5Prq6joV0nmWLPfdjCQYSdEV06uwwyUl
whcekAVC4sSOAcVT+9odZYjrTGAlIybvlq0qDyzkK29wgLRqLBRoRR7BBz2S
QkoUehgz98ASUDJfb3vkWInl7JS/nImNeWP0C/ec5FiCgQTiHDwBydT4yT74
N88iOsUyBmDbtjv+7kiInZdiN9l+erVJFC1n1/3EZmAwqZk1Bi+e+uKmpu5g
RrVAbpA3sgObHsxRSsDGorco2e3pzL/1bL8HjfU/2vyaSB27vjyaJJUsWAK8
x2sbCt0n03LZ52zYQtkHnNMjW2RkaTudURlo5Ey3pDYXhohP3iAVAZixl1Zx
uF1wYwDZaU8tPHRoOOJrTxJbuZ95ZMgO55xPP+XTrYJYMxIgBnpO4jNn+ZR6
rHhnhBdjFG1/CiinN3E7hD7GFOm/jiNfy/URNBXgudmzQYyP/4dsslOzH+If
Ewhi74rtrADcT4JjJdY4wV4DOngGS1Yv89GEfhJa3pfH9mEev8tDuwr4RCGt
Z7oKdw5FQRAZS/kCZ0BE3txwsNxozE/ghAmSxCHa3LYIWUGRR4gxZUtH6E0g
F5D64gC7rR9ebca8nLuotPUC6u/c9BtKPetCz4yAKbfvCLYbcdeGlUKQNtWw
JQypZZb+uCmTxorMztIf3YKzzCrt+XZP6Al4X7Apo4F2sNJRADCmlCypLHAI
4hVwpRx/gZNwCNze0DPtKBAc8pCiEqJMigoau5nr4VCL0NazJpOupjinPwyW
WEOxnT7T9P6nUOk/bVP84AeZEnkTfZJvssrExK6n0/IKuX56WJ8J6ENCa/G+
mApMM1kemUv4BPahkJ1O9uAWq0gm2iaQYIvmjT7ChLWgUD7zc5318hW+zfYM
5BdipDBHE1crU9GUylhqM46fwcVEzf0F6Th8dRN/YbKwvHN/pqjndccY7z9d
bczQ/qhQWsP1r1qrkko9qbtaTH7FRTKs2Zl9H1XrWEbwgS3kEYrFtRj20Gvz
qpWdhV2ULwMPVNi2QIRtXz6rT9vsb0Or13BFkLay89jI40UniltvZIDcUnA1
cM3RBCywbxjkLyticltxAtkYKIkSEE1ZzqG7khj3XVYdt3c2xat8GA23j2ur
ulOMi+1KGzJeinSkT/HROJfrB1LrGMavBqXub65+PJAgLD8uD5npsKBWR2Ul
p/LeOls+R0mqkEVX1jwBVrrivzWOxgAnBFwlcEtIRlhzBfSrErYkOQxJan1u
AqO7UItd9Hi1I5l1CTsQ5RGYTbqhsIq7njcCCuoShjNM2hOGulZWB9u669tu
Mt9pm2goaQ1H0ESYH029mpfVoGNgz0uwgBG5VTJe5W381PMgcbH7+soXXMA0
AETr0F6ba8x61zK1Xw3XoGTftVLRkVuMFpAynayv1sLO0HjAkI+mRcJwguA9
vYR07M2sDjxm2O5/TkAj5BK9ofw6l9pzruN5Sd9TQ9eTOxAp2NEoUvnIJNhq
rWu8gqUoF/Mg+78jgBjm/tFL+AEqOsBooXsKijs6kEp2al1n4/ZSjLAFSmlV
zh+xta7lkkmIuT9R2E5oCY6cavxdy5ZJxsGHt8AqnT89BPGLjdQ1jZTa8UWU
qbs22R9KI35A4qQnt8PLaDLvsFXHkBEVdxelC98HpITNjgfy3GdRiUJZ4qK/
AId9t+qYWHXN+5JyWs9xe50DTqw+nR7zaAzec0ev8Wbco/thOT+soLD0Ao+v
PeusiSCuOjsJbu5/t3clFKK+O5SryjMnwsF88QPcQm8QYds1VtNhSiEvzw8o
d2ZdLyLawv3Ng6+rKhin7ATFlOH7Rn/BR3OyGGdZevPpbkx2phJ9P7chONzm
yjIcxuOiYfIfxWN3Ku5qXACOgfIZi8S6b/oqht12Z9y+pSGt8VCldrhF52ce
5sqHHxZbuSci3CbgLbmr2CYSIvlmeylygLg/nQ3ZwJ4ZK4zWR3wSleKHTRRm
MCP8Xe6aDRL2DI2vW7G8NKXgD+uSzYEftWEXcEsVDfOAwRi//Qx2TyGVuIS2
+lvYBrdEL0ZDveUIP7370BFD8QTCxaAT2NWOvAeSInPaMDXvbAFLh0aTv/Y3
3IfCLS/Q2B2QrpUppH9bUw2+G95GenHyG/uB+pZDVqiy7IPsFXItPYa1BCH/
TJflfOOB9ePK9KRb3pQnJvx6pf/kctuSkfG5BdOULA54AKyIuxdEayPzoJtz
pLdBHCNKJk4I1ecAquDMI+tnQbd8EYOr3e3qv1jsj01Rzixg6e/cAu1m0Q4x
c/Z3lypsT9X0GvbkN17vXrSXJ4GXF5GZFfVWa0Fgp+TDfYQutbeAw1CiykKa
bw25iNEBz4Sun5zqkVg6HmaK+lMrF56HDPO8MwdNr+eNmEAKQ4ESJUNsWj4G
GH7hllAxDZCBfeGpuhbgvZPgmKC/uvGyLqrPkNLBQZxFZw/gJNvNVi32mGVF
8JgADl7/aYLH9sxkuCQpkXtTaY3u2pjc39yA8q1FLWWVRTGSCqKZLEN3jzGk
zrmP4E4Z6pmAe2Rwcb/0+oombuezbbpisCTnOBtfxkT2h6ktpj8WrbGAYhwb
uV59ImEZAZCH5wV2QfxOjmYt4Rpdxtxo47abOGswdAGi4qTdqbXRVYcG6aEZ
EaKF28kLK7u5kQVt73Z5ETvlq+GF0nUBWG7RDh7APE6UiiLvEYMCJolfwolM
MmnHNB8O5M7tjBOAl6IrBEMBo1mcHBul77JPsnJeqlQ2D7RzduFBfSWbOMEr
Lfb6XwQHMwvR2RMvSCKY7wEZ/TIBUTpuod8Do2xVdet0YVo8StLZLlJ63CPm
3u35WiT+LZS4cRUOKF3b7qwfE0DPA/+SQIOGqv+KoEi2C7PfobpIWZtFLbtk
6tSE2PhmfBA2RPrvGDEjmY0EG1j2z2yqZEXJtU/AQHVPXSNSD8z1TzpmZgWN
eRypQzVLX5CdOKSkrYKuE3xrWIF9Gjzw4p5Oikeh9xhNZJ80BJ8N6M8+iyP5
CJUx+Wl6aX7dZcQPlyGpDItrgu4cmmXUwjzWXOl2eR1w4Tc9RjSwAypbowd5
vuwfto0FJvIn8cWdsCZvH0TfQKFo2DljYVtSOZirhScbhcqLsfij2M0E/p5q
Lyan8KHdUaqLjuGj9U5F0b6f7GKsdbXT0jBRZ2AQEbgfXXy837Ita58Qs/Jq
a6xk5nqJSXkZ9Mnqe+No4O2d7qFHFPr7u8QMtIjgbEcguWOKiilYj9iOsJjL
p5+j8lM7Nu8SYXoW4GduvOxqwRimTpaED4Z2lSfDzMci2xwUAx5c5f0VD7Gg
p8WZ5FBXxzZcR7T0tRcCi5gVgDm2XhF/f2kDcrzXZN01i7Pc0GjkLthkRgsq
mkZfXHOXlAGvqZqcir75RqSm8cDH3b9AydmqD33otNvgxEsCw1kpAzVowFXG
vgxXwLzFBXaq57w+4M9yeTaSCXe/208zIhIErNlXD4CZeUmYFvXkARDIrxqd
i4clMCA1XvyZfjmwvdxe/BN/oITRlaIR/0AGBd/Ss4LtK+/DuPnGsGK3DDB5
MELn+1S4oD/tUaKZnNtzujPu4cy0hCz2DtNqsMIvL32bcUEW0v8eJdANcMQB
ag/IzVMMofi61jFZXtahXTWZqd6wNE9mYfrvI+jTVBeOl2I1B8jUDZb6rYcR
dMP+B+c1L4f8mf3CkIIpLkmjf0SnbleZyMUPqGKCf74f+4JHhEGPYbEM/wP/
A3RvnD+yCYcPKzgg2yCfnSaLM+9PGk/LZ9OX/D12Vr+ZU1F+5mC6vRo4BRdT
FXpL0tpzKhEiLqvkdnm5+dYsECJXqwNVaimO5UIK/B6dLOqLaDISJQzClyX5
JHNibejMcnhBoI8OdoTg5Pp+GYiZltSKav5eIFWqBF0Kfoizy/2K1qJA/OUT
IoB+u83F2w3xwb4NsXXGvZIKedaYIwn3i/PwFW8NWRO2o+VLmHq6gIndPwiD
ZyA89g7ci+gwnHR/K4kWeoWPL/lqYs39B8p67U9KQvPe54xNrQSF4d1hWA+X
0BtPfwnO00q3kz9P9j9UYZjS3VR0qod0My8D49EEuwFnUmkuEVUp2LxPzlQG
VggM8bXj/vb+YtWJOwBRaqbYaHrCCpwXlq41KqjhjUlXfkivaPqxVwNIY1tS
8DTn86Y7x22RWH/Sva4qh8nTr4GXnv/n3z2w3YaFKlaFugS3oQfEfLNV2OkE
bVk+FNTmfzWbgowDBZHnSLWgVLdCa3Pc8dZ6wZNwQQ8ykFADLmXFR2tDQQnE
6LmHhhrTZXGu6rM59+dlNeaLskyBuHNr8Eb7GVTBMkMoFsJZBgYt9TbFfYQT
jSf9eiEBS5JOa0tWD5eerHsy6qbJHaSC2Wro+9Wo/ztPI4JLB+vT8rxPSis/
zsfxmxepe78MY+QnS2oPAfniNmvpJpix7O4h2DOUZjbk/4vEc1MmiSlNT4wp
hNS1iz7ZDgMtOLx+RAUwf1s9lMc84iwSX1+4a2a/gRZ1wi8Mqymhv37Sz6lB
4hHmCJTa0pL1M/DqvpO1pmVabPRg5KOCW5U/1a2ZLjPUIvN3zfG0OENFhGRv
oloj7WlmxxRMVbUenj7l5cgmSiC90bjYk+bx2kyr1pkauM7GcNyBbHUFLDsV
6XTTmHTCg4/PAb2E/s6CRfPCA1HOetnnnhIbYfcdQ34NcPMrhw3UZnkYdJUn
dl7TMu6mOJfImSejtMY5k/ZljGqM5stlAn2nJgnS/X4MiNv9MxUXy/GZVJdx
/WiiU30bGNT3IHsHT4eK2pU25Qq0UueSnRh43nNXy7Mps931GHiSBd71o0b8
XK566+PVJkLQ2xR5xWedcb49404Y35IG8V6/uF8uHiLSBt51B8AD4vmn1zA0
y+uDhXlS0FWBL4ce+GEJGFLZd6IqxO6cyX3kmKo+xMdoO1k5K+g0P2NA60Eb
LTiiZSIbb6JA7gA2yq+TjPRmvnBnvtg/+mE9Tov3s5xUO0ZshDlBH9sbOLYw
m7a4m3pSJJDXG/M34pC/2q3MTuHcXvHUxieAhXvfEbxvwI4yIgavtKnS8q2D
Rwq2BXDied8hjjoORZ+O4pEhQhAwLRT7K8nHqVOAHs2zMnpJ3Tlnqk+2x8uO
JPj2HunxTIlda5G3TPHC8H+C6mvpFg/VObDtBN4bnWNEG38KxrBRNL/jltDf
KWBosfvnV3EiYCoREIu4lXVRO+87cVr/qemYl6sVkYZILK2g8jV7T24y+f6S
J2RLTmYLz7gRjoz1tefrlMth0EaYlGkkKqELZpsFBaidJkIL/NVj5NdtDYgu
FB+/12Q/Rmyb0GfS1Pk+dWrMLQWdCKF4eB9bmOJKYYHX5zFlEP66YgaVSw6A
Ktwo31XMUIyT8M8jAVda77hS0dwj3LJiWBLhcoSnBHGQulYjGK1XuO/SMQ5y
yKL/5r1njGzeNpA0ddYzZZ2B74w/99nHbilrqrYI/56gZFaPdVYFKNrnmp6T
ItSEaJg7anBM3ZIxHruKQoiqNbDsrur8u7J/dBPLyGxkODjbJJaCpier2/S9
VaX/wBXJAfumQQu1rARKIwUpjIce/AxuINJl7kM8a7mrUyFLPTyen1kefgP0
NIrkcfScLe4SpTQU0n6Y9cELj4yy/wWd6JdjCLasOEACLwjvU6ogKy8K3Ktt
U4d1MoEB0597C7NHWO3NHiQ19KwO953Wz4nlK02Z25+E7ZLnEOeQbh2jG+HG
SsWMxX1GR4qRHfpU68Ovo4SX0Qv+LNg1dPkOuQo1ltZDenh+10UTzh9Bi5Q8
0hBaH9Ebg/0F6Mda30YT7gz80Wwf2NThN7t0cyCvSUlltasWxHthAmhh5hwx
l0ZnuB9nCGcWRyWWORwCEBneyx86T/1HR26CxsStlUK/QJQeAfcRYjpWOO7C
1UN0m8qN9bXpdvRp/0/4wTeVaRPr3G4SKg2uNjRkqWgWOom0Y3yM36GgJ92Y
P9xoa5QAqXSDEgJ0bvRsNKHcQ/uqMqIDRhcHIuQ6Na9CoX7Pvb7Z2hzV4haC
v6JA9oqlfsyyt7V69GRJ8HGb9TG6wYTvFsRsMpURANp8TnBTzI2HVk5/wFAG
q78Q01ZzXI1EPIeD8qpVsTlaWIhvilrEMtxYLW3Yi7QcYKAQAc9+ArR6Cf+p
Gjw9Tamwm2dBoP2OsqmYDVPuP8B16ryGsdIqg1c/HqVXyJ842gSqLoaLAolw
DyvKXsPkdop+03AgzTr7VfGD71VnfPrvelCxA0MdJxtYHAc7aoSfI/UoB/+a
2gVn0nBsRnm1aiytsgQkNlY6KNZB7/1FOVjlrRkxlBK6DKnRxyvXu1YKCG1a
RKE0YmzhNlxZf3UdJK0+sSwwa2yOjJjKWjQLi7KjXQ0LMzKsKmmbGxd53qIx
wxMx4U3HjTHovx3Lum4TL+z+U5I/RyBAWgQzawkzrZirA593RMLJpB46iOzv
sgNlal9GHpth6jGrY3CH3gs0HmzSQBVZEIYQkXOflqEQLTC5Wgbv6uinSnld
36ESCYBxYz5jlRMF8pIIxfKimmVLvllDfXpj7LzRW0oap0E2MI0qKVPFao1U
9vy0jkZNcGNe0j81IL0uKAC5fnZLmJ2m+t/0itWt/NcR5yNmfH8F98eexWIf
HkqyagbprMfzOUSiTnQ0epjQxCyrga8QiuPC8SZszu/RLwhGRL8ka5bJ5LRo
XEqOSSkVCOgETx9xGwS5tAdw3T7Hkxe8B16kiTd/Pxt0mNmdKp/3RSu0Nby5
LiRZSvYUSH3cUmJhDjiSCxCv5GxGW+kBLeKQbDVkJCYd/4dFYGrCWxQD1yeX
fh2lhBh0RZjN0xZNI8T7uOJPy179XEzLms+hmoun1XXAzXXDdmnTHc3kGnQJ
z63reMeogwLfvqb34P0kUZlxqWC6hr2PjNHVzTJISg8tfyKh9ZiXNXmIg25b
N7iMGPqB9ycNuY12mxWSBDwpaKvvXHFj4Xe4OeBQXtE9jzGaP+EpcQqPv/cQ
YidtwT/ZLlyNuGdCz/tHEKDPHP4cq6G/2FGNDVzMDxIjVQyG1jBqL1A86/NI
ZG7nytRwZsGg1y8r/QX/WG/LHjYHXagvAsc2jTgbJHmsh1Yy4w5fnFXTgh9f
0xIt+0uFKwVR2sGQm9CZ3KxJS873lFueVj1x/3E1qYDOMnBejTkJKPHWgF0i
ewgkS9mnqfA97LWVZNQHDmUgArBkYZY5nmEJ+3cfOAffHpcDjMOyn+rXpfxK
SYPDBrTQ9mb1aVRjxydmDIp4pXiL5ACAWzRNfYu2Rr2NN7S1t4QunGdR03uH
tm9mEDl7xZMkWpV9JCo1yw/pbDVJwwNKT3lrI6/L01VkOH/Qi0P5ig22dGeo
34y4qUTnA65VPzKZVcT7kjnLnTr8xATNckolDtdTYcDV0Pwiwqy2ZUR8A2KG
9kogeCMjmE3Yls7v9/wQK5VjDaKYenNW4WxFV9XqXkdcZYjaIvmOWbLGSZaw
9DNLNb+6EnG5CAb34ZK5PZpZbSWADkCMJlxC89KFXbieUC9iMyvCmlFabhhU
AVmqbTRYK4rfjcA8qVB4SBw+iscZ4dUGhFt5ehlN/iHARsfrhQyR2ZSFR6Gr
W3xdhOFiqmFR+2b9Fq0A+aao95eRqk7asAuEkvGmsVikVRktj0+Do26Vs4N1
zXDTv267FhjdNJQmNjML+Va5l3JWDMwDRKsE8gWVDswXJMvfqwZGwiIpT/XQ
SneqBQiPiZAo9YKFxM4DhD2uldlEun9lc9ZrGOYrhh+NxibTaNqDYx+Km3MT
CHJWdSKQTdZ7R97kI/rxvJb4kLnxqSCPqrXmznMLZyZcfDkySRwZIYgrvgJs
TdWzf77NwzkHerhLkVX/57skBq5sabELX9qolckK0yd2Drbfl0gXfYEwv1HG
MPFks/AqA5TQ8V+LrkB6N1/zdo+d98SfqlcSLudVlZEHPUR6wR/GY+1HXze1
nadHiQc3C/+x5/EVb2znOT2WxlW8EKRyEIRZhpp+to9bZXoLgB4b7d62tY+9
7+sLdnwg6JKnJKhtQG5HGbUOEKAFjiDD6gh8z6X+MuZCPPsIOeK7oW2qdz1J
8dQjcg3kUyqAM6pRHGF78m0H4lPhbwIOfZDDrJiHcMR9dd2XQyWQSJ90UHE5
Jgl0DlzbhfCa0+xwhuQqH7n5Eei/h8J0wEMRxmRDPsKio1gOxuImAzTq+anG
9oaR5dIy9RV5nuOHkBcuycK8OoOiAxbLvlZU5cH6p759FWRVjcImu+mT5hSX
ElIMYOJFR3Hhv2fMh25NzKroOKBEJhhgfW+G2JOfBlQnQ/SYqYTtF3C+Erjs
IG2elfCKGj429V9Pw0QJ3yMizFx34RFEFEP5/kulM5c5Ilh6XEMIiqttHFCQ
shPMrEO/2xfipKYAV335WszmWR8qVL4DNmzate71n61jn8zjzFTKJ7B1aBYQ
/+zCnqSO71xgjYBKs+Bg8EyjM8BpgA/2UgftjFVqpQjGeeTwXvAelltP7EEz
lKpVN0yOrC/BAbClZvRrwSdb1RDV+E2dRgFrl0wnK1BiuWjbH6riOUlUGOf5
eq8BCqxIPlONZCJweES6JUNlmSyR186CrQSNiVVCq2F2ueNe4QeTgnzfepEy
urnkJZnVdPRdu9xMOGlOjBiX5/KuUYUkVRJ0eSWXYN2S0Km5KHOrmQ7cSoW/
JksQDeLDdRHAZtgTNd6uabHABAtk9JmMkh9AaG7BByvMEkiP32ayflaf3nRm
uwLIxKTFLEknk9P510GFC0qUUIQYpUHGRnnFYcBngoa5crscYxEEo3636v/8
GkMLVoJlpym7MYLwwa8TGPjYSuHliaj3g4d9DwRQQoTvO5E5GZltkI4b82Ry
UCQKA6jj+atmxdaCOtlelc82KtF+oLFfl3skY4kev+tghUXd/cre5kAHYl2/
WPPwktIHiTBGamG68w6waCmTtR2tWroVJnSad2WVHEAmP/YzlO4kkfxEp7Te
ienZihCCN5fR0gOYalUhXsrJ4doN9F3CH77EQV2CnevsN8v8Rl5W/2SBxwza
W3pLm5BBjOM5Rt55vzx6u5KfJ7GSPefhERmDkiQu2vismLWMosfFqQ6MoT7d
bg3qb+NfANzghsbDP90z0PWUZgesKZM+hG/7ZKe+b21c448WlIPk5TG8Uh/R
Zb/uHVdQI8CTjI8wbaI04i2hvqYwkTPMBy8LCqR2h4AitgxnFoOQk3zNN9Xz
sI5vce9nUKezPlv3iQ5En7hqiJYcnMgjwFLlChbVQhc8sMkISMw6+CODlsUm
C3Z7D5VpnFMVyWTAkFfz7GTUAlc/TEoPHy7WE9VIJ9xbAXX9+T/k7xS6hGPl
FkbykPJt3VTkM/dQCM4fP9Dsea5JT2TAHk/KS49zR9aKxIipBBfDfjZjGar5
PXkyfhPZT6Gt2odWdNKjQJNOjnVHvbDxicKJmB4uycHzsmp8gjo93wIYaSDB
uehAfvJ44iIWwxuBFBR69jFyDtu46eg8OuRcjDBRWTNWhSKad3HZ7YtP9ZfB
AvlamCs9KbMSolx8B4YdICgZXFS9sH1KsRFgZZh0i9D/7UCQwgK35aHOAEdL
5FFw33kzwe95WNT7KL4OuDzGOWM4xVAHLj+PHP/TAo1ga5FIYWpQRrq0joPV
32CgV02/4kkpzI+rY8KE98yoE6bPXEB18tZBuLRMlFVT0KDU/r8wHYSlhx2U
UJpC2iNbU45+0C3rBqdF7PZ+WrVoZzqr7dgijayHwIFhAmjJ/DMO1ncUzPRv
jHfqUllQtvsdIA+93itIf1gEJWbJPPQV4HnhH2ZRkAUF/jBANNX4+jjuo/Fn
l3pHPOeAsP30z4BnLrLxiNHN+HeaAmD7vbypop0KIZ8a6g+8RKQcOS5TwgPi
u/rKTrPgmb3qj16rv2gMt1jHJhPkwOi8lRBmIP+ihcF4W0qPY5v24i7RFguX
NhD0gHo8F0CQOx6mM18ISBqiQQdMICqdrvYbfC14509mdbppbUV+ryks41ti
2MmWaebUiSUeskwPwK18F23ezMFJuwUn3mM3iM0ZZOP4EFRfp2/y27PMWO8j
Baa/BBZJABTcE7VLz0Aseb5ctVJ+diOLbAcWelb0gun8ACceL+Fc5TgUqJUj
0mcz9FxVdvr4MKqG18pLxLcZknL3x+Tk+J7OYb9bYKk1POO4BjHCbMvapd48
PCRKYD580D/nhTC8l12HmVOu1QXxmPDxb9jJ/YONGZasm7pz6x6Wb6aLhyDx
Ejc8bPhuXwhS9LQCOCcGP7QHfBrAln544XVEQOUS3LxLO4w1CX9wmALh0+Xc
TDifnNtgc0uUk/ofg7oM4Hw/IupyOKKivT5RwFY2BNTxrzi0E5mDZNOIKxHX
yay+AtluSPT7TZThHS6pH+Mlpt1i8DtLELuVtpSDhuCKeAmx6oebKhVn1Jvb
fN1dQ2o0MOmZojAMnMft5knAOWm4opZtjo5X90OaeQ/4ewPrSO5CsORahasf
c4ECOmUeZmP9ytcTw3shofar+7ZuQ7YUhlAwW4KJ4ip1GhwomX58P+hdQmR9
mw/0nrVuxHry36v1S1mldP2loE4PWOdbXDl/kkxR+TAFQXuHnsJHm28CJTNj
XTjWMOzxOtIWfmiMqOwesGjpnYCxP2UR8klIpO+O9gy+sthowDOVwQx/kCCe
jZPHZvpKW2Dg4M7G5xMPMLEF+hydeRpfVpOW4xxqaW0v0qNmwyLWeIY4FhwQ
qNRtfwUWifQROL/Wx1m5D4sQAFHqe2fbii0lDc0IqYwwGokFPhMY5Rd/frNv
3v4ZMH9xgJmpVF+mNOq9HHGZANsbbMMIMAtrrDMiflehIgrvwauVPydTatC9
Pk/s4Alzt5ZraO8hbaibk+mRYmIV6OqY2W/IMs1JBeFo55UIGo9Pth2GcTQQ
muosncSi/8ZsjLAHjb9ORAaYl/wbEougYHhMz2YJuogs18AgWHaWNSEndL0T
m9NRxcM15RxCVidmDDK84DdYkhNluMuyksHaafXhxYUFlptjkn1uGcDEKaKI
q3JIgHxAaHib0N3gxqsKZc5EANNdcPauK9ilXPdiq+Dny97JaUUfjLNB0V07
5jLLE/pWs073WziYPjypY4T6lIbyH84qC74lYmThApKtxDVcdIRew08MdJTi
aDX+LS2h8MprQV72v3iXZlcqbS2q8gphr6l25C5pkQHshfcRSVMUAsv3PCda
b5kvb2nOAR5gSI1D7+LSal3QWiU/X5fjFpagD/eHwHN11y59t+AGGaAY4aeg
u1ch5QCW2QJFJHeVCQVU638/mQ2+0rzz14pvUVtjeH5jhwE/oNTnBa3Jsc+N
jMKedBNl7vhUwmb7V89gLAnFiQ4iCcLkVF+ovHsktYKg20NHUm9Ie8J2Vtmg
T9OapKwsozzwA4F5NL+QYdATQcKS0ZFK1vWiu4iJOTmddZczZUmBA7QW2jeh
okxsybGHRxF5sfA1mDxv/rzc8/H5GrOPhIv22ESmRtQviKdP1AbDWXDqkhC1
OXfe1J1aNzmGqVPr7OYqX0lxNYZ92GtD1Bsmsb5Qhl3MkZHC1dFBQn2pqfkN
3ZPgZEyK3W2T9aRcDZUPrdqGM+KJu5e80yfBDpSWs3mrztvGgIgazzzW7WfM
ap4kTY6e63DrG+fS+Z0x2PnPePvsboN/u+KQXaWNVil+jkxegq1IN7tVtv4R
b3xjM6nvO/RJ2eQ50D8xqleLNwL7a5SKYR6Xj6C+1gvOFS4vE70lX/uK2WFU
qKPj4Wz/I0+NrPp9yHY46tkXYhIowv13TzqJGyvo5ikiRYnAttTtvbAhZFgu
8cc4iDVsitnHE2jzOI+onXRU1HGiCyFLsWnrvK7bsru5CbjSokEHA2KFbsC3
mVc3PwS0ZcSiFHxn4P0t39ReOCSj4CGwgya3OFVJGRy08R5/lts/emJzAVJ9
A9IhBHJT/k59tcHaFxxU47cNEf3pbI2BskRUoANei3Xrt2nSTV8b/QowHYzM
++k7KyYced5k5lufaKY/I+nY3ngfe4juzvHkFps5tsem6IvtxcAlD0+F0dov
+tjp9SyoAZVSacc4lv4DEKJl5jx/eJOrk4ceU8DHA2ucuFSwXlBOz8v8quuh
USPY4PUFHXhuM1Fndyhv9/OC6KJo8zM3dvLNQiZPtqtj7NIrlGl+Kd3Nx3g3
ToAESvO+6MSBf9FH1apGAXWBLGAjVrovSYRN+R/weqEiRMWBqfYI7PNK9ZrM
EPbMzaD5cT3IZTPgLtR7iOk+8l0QDF4YGrrQJW7lZFqQ0/9U2afJ6UQq24hv
/Fzu4OQoYyOq6bNlfVadEVkPwn2mLq8dxej6D1IwNWw1VKOZ8wGOkrVJ6Maj
Y8QpaJBjOxJpurkFhh1b/G9EGI+mcKwn9W5AhyJiHdJy/rcTf2nXbf62QazC
oVCNn1fgcxFhxXRMnvMgUYTjA5ekBBeK/NPBEMlR49ZLX1BEYQcCfbNsIVoH
E2b1SFkK1ZetdhlWawAYod+NAeN5i6M8Y8MQmYFyrGjaNQlySCOCVLoiJD0c
9StHnRtDmxyzv4NS9q1jPWzIbSwXIWKPkbHlG3vvA827Zh/mIXHAwiXDh0yh
i3r9wBSu8WOPU/iOyt4gypULY9RsVG9Ppu8AcxoRCmqiTlE4odgUJ8dACmz4
BQ0sE9I0ES8jcH63hsMYLV70DaX6VBS5Yn505DX9dIfkcUvGxbixSZQEb9T0
WyhbHNrW1+X4DqiJu1Z57bnIcFlR5I0B6LtvuZtDIBjm+7rj3EoOQWohprQ1
zG50+FHiO0fQusdZCE0p1HEOCLszFucv0j0eVZWwN7oWYIgH8ThXRNbUpHgU
8Zt5zHDLjvxS2otzKEN3EIH1BwCp5haWQUsOI+pD2kj/yfXCNu41+MvZC8Hp
CyAxNe72SkABC8ijirdOhQOvoF1mwV18dXgfrEmpFFvi7QnL11KSxkcNd94w
WqAjdv66WKPAro893klOrRbh12DJYv+Jt63OCRRHFS4QLTlQ9VmPp2dUs4eG
8JW+reOFv61er1XGWA9vZjVxY4iomvKrpboo69xTJhpTMY8ymLWRbm/70odw
nH3iAzYUJxXr4wuwsi7fgsPk/ipoFO4t1z2ec3O67Ew2dbF9rJ46Nh0dS5Dj
aaccPHlJHRb1cbFOu+fI8NNE7rsaj9OXnxpogIFzgfTZsltRFcVeIsyJivg0
IzMv1ofAG8GPs9utdj1sizJCS+pU9Mm2L1EvWIhaE37KhUuI6PJJarbymCAH
XgK+goHKNchokGz4WD7viJQaEvqrOeZ62CavUUw3jJgAOUzdhbVWyKkan/bm
DyJpDeL4waBOwu1g7Czz+Qz/AfD5DOkqEPxIxkMDmfYPmeSBysBp45r0R8xw
BkSYfwKaCxNb0XkhNdRlA8LdmI2MP6pfPmTgAjXRgYNjx0JWjxnHiBDq8ZcP
dzrDUpxLCiaDsrzC/kKpyVsRQdTwYGTSDvk+mkAW7bE7iRBDqx54DPfunJxL
grzRCGeA2UFfQF/J+3/hnq7spNq/+sBargdDqpz679mRP5NSZfocAnXEikki
Sgzf/SKejsxCRgYB3Q4i/T4JgFv3aGKJjh9e1SXEpXzK/pamRJOzOrWekWZu
t5No43EyHcP8UwVkQdj/XNRdsGUJeNUAX6NI8+5ZBVzMDC+gofnF5JHzv0k0
Y+CNNiYwGgr/Y1BNAC0hbPwPqOX/ZlwWVj9OLwdeTILLQGFFa+URz/A57ItN
zE5D8uvVoD6bgDs9sh6EVyJmBk4bmvZV2t9HhQfThhOvu0vkRA+7Dx150MoW
x779HdooRktt+DmidaKhCVwEDj43rx83GkRNWgpJ0xmDAFgy4sP/Sy82er3O
n+jPCk44F5Q7LTi5h5/6MEDE5LrWcdHt2CuhruMgO0SUueZ+16Re2F7LPnZg
vvwo3GzAvwKHzAnYSrZn+Vqj4Mzd/ZUxuJuSqdckdxsPCzThJtUkknYLkDXk
xJnYiYAuww7EjofAsQYUHhxVHzxzQvMHiBDpX4r7XR/8vViYxigd/ixNYcq0
dCTWvRnq8bW0jYH9zxF/JIBgKOj8qgo6qJt6PGjN20tD0BlxphVu9QoHhzGw
GHqDFyUKt6fYEKyLmJPphNsPrOJ/SZKsiaNGtowdFuTfTgZa0QLc8KD+jHO+
MKGnu52fFihTzNHj8C/34n+rnMwXqXW+vdA3vsLnUL8/c7sWJDDV451Y49Lf
xLO7KVOL8i1Rc4CiAmclFUrCOa8K+LHwwp63RwxE3QKhNZi9NhHrcxO2XSOh
04T4JP2p4Kf5wB/AyMvfjh1sscBexKGFdSnY+Agjc9jwEp/Z5PwS8jrPtR5m
8UtGyE6klmalkr2/3dQ6MyF1Y1nZltGiqPz05piLFDcCwO5s0OwgD2Krpqqy
9hxMBmzW2nSsSAPy8zdwTmlJpca3RP8y7nXe3TyiHtRwwIf9KXn29aeZmqIP
aYfv1kiVoBYhdHyyxrHyL44gus5xLaP4Xa6SZeCopAQxhQwA3FmeID348uA4
6c960hIKw2i0GmZt3MiFZfXiFCD3gOGsvs7LA5qM6F4Jbu99d8XljuDtnFEQ
Rsn+3SMWZ9PtN1oY71UrTFX7kZCl3cCluYky+1NpHFTXRolwEzROlE8LIpDh
xqS3jj58R6HCaXVvxiQWNEUlVEADjpFxfDc+QP1wjlI36AJDUdIxAp+WceMX
D++VtXdXs2id4wjM1gmPdLDeL7WkR4yC0gEBvOag4cbOs9j2ClTTubSLntvD
+ci2/xgfuFKXZXLGTojDGS3Jhn4BcS3A9gdNlegydxP89U6nMV5RBoruEwKU
Q7ZtF7w8poh2jA1PJeZLIF1Bd6I/kzUQ5VYYYoktIIkCRY4jbXPKY3Uot7B3
28ZiXoNs0QoXbeUjLzeRFaqMVQguL5L81b0QddxQ3TtPEaI4rNmumNpsobr9
B3GwubJ0x0lnlY7OEwpEIw3Sb4S8xKtYVVtveVnH8c6jIEhJ/mdbb+F9Rm9j
zw4+doFOyTGszGV7We5IIHLSe0CzmWLLq8ib33Qc0yhVz6I1SQIB4O3SmT+Q
X4cOntyCSq2R1XjJx42JM1WpMbqkoUUa52LzPT4vrrzRg+HE7EDrejSvn/Bf
aMfngd9oyWpTnH5nqtLxYti6I0Lf4D+elLnEJF5pY/RqCF9kt5qWZDVMY6DU
MyKMrq8MaM7+AWjOkbtdAeK3pP0I3K8b+ELGe5oDnmodz3TlVcnnH0wy0494
mMfbkL8Meg5O0XaXLqwxT7NK3ZpnuGpwjtBBhZSzT/CM4x3rGdT+VclCXUiB
3AxNOXrz30rj20wPhG9vR3mkkah0Z+YCc4Nl4TYrOkFuZyd0n+o4ifEF8W1w
jqF6WLFb6yLf3CjdjheaTnWtoOlz6vS/KHTNZT1UKMcCnjDn+sxETWGMUbVl
Ik4qdtwzpmj2ejF1Za13JlwA3tLmSz7XrbPPyKF7ZDaYjkoA4nAplVGS/h94
DzSvC8J6hlgd/RzK77Aja/MmNzj3kyk2iVd0HN9SQGaHpN0nh/x2TfkmQOxJ
YfV9XYs1fgWphGg9CF2ylF8lLxkbpGijsUJxQBvHz3E2V6Sy2GFrULMgOh0t
5CAs/RWSxMbYvkpX4P1CmWXwwnzfgdPEuCct40UoXfdtCQvVMNi5XdGEVB+w
3On1NgJgYdqvoaVPNCEfXOz7z8AYgpdz91qMMATKg9UBNs0kHQYlF6NLXVVx
Vc1qb77N5ghCVhXR1ObZUMEvIDDOsbfKl7R+beTY3UtOzX15O2ooamYTy7vr
d8UmrYIxOChQUetqPdbcKSuBOdQS4ePdCIlc0IKvAFLQSh3nOKAwJacDxdrV
6v4LekvBC9s6HFYCJh57VAtVzDLhSo3npRn6CkIKNj9682xRObfxlbAUJO5x
0QAvMCSEmYcUPhx61Y823QF//yt10LO071SsE3ayPvlx526Y5nAzg0DcqSiV
gtSud9t42ZQPdao3Skki8HSh8xbc6MfXIGiJzlz7UM6RPCYDH6MUQiusgVFd
cDaGY55bROq81D96McQ1936zNJ6auV717AIXPxSGS7Dkq0mG5rtnrqdFkkZI
sd22KU24gUKz6XP/gIQYvH0iIV5qLemX90c+TL8VOXleCaOd/29dRWo2ou77
Fhf8Fy2GptRbT0ZQrGC4nXW9r5MpV6YQ9RkUks7Mx7F1uQ1oZ/fX9XmW3gty
2Ie8T1ZVPJDStsoqsGzARzbcD0ci5krSmJAEuMeDgHJty9YwAWCVT26Ut4tK
TBwlkdxPx+KjAjDGT3nO//hYdrNkR9dCrHkuUsZsNzoavO+MZ1k6wi0yHQMh
B+sWTn91M0jCcPiXTlUbegmzk1V4wZbLQCkFtbEy4C1W1dfW6lsmbZkCtiGM
sy3Kss++qgvaO9sXA0O0N9lElMSi2ASY8vw/pXW4rT9qyQHbJt/3GJ5j2uLG
4TiVeDKPzQd/BxfYrkSZ6wfTla0MRIDAKcQyDnxKeoCDkXVZ/Ws+oeqmSQqh
Cp9ztzePQ148zJ3zsHw3U46hwhC2HDT5erEfKVzVOILVTdKMXB6dr9yzSqUd
+a/72voQxaQVk8lfudnb6erQzzoXoBrXPgEafLa6VE2YtQmic2rY/vJCPLxn
nJeh34UdjVbvz/y3piVd35RtS+DnRTRCPTdO9IG8gEFduKvy84mbAQbMxGxM
B5/b2NhMyjVwMTDqHSUPQGCxzCwCCPiktY/oIHWCtjsig2fwzGSFL38J/NxJ
R9nY+Kmwww8j2KlK9QbKIqaZF6nEmKxjWJWgDVDuzt5lNR1Gjc0hcZba1nJQ
aBVZj0Cg6GcrctB7O0WNRi7rcI9RHVVENPuHjWQgvkYhHWbH2ol/N1fGokGm
QUd7R+FyOTEJW2vjEvlS2BqoNsP/duUzUZwTmuW8ZZlHdtng2D2Ftm4pfYkm
E/Y6rEUgr4H5rgXATYYLQlleIZ9SbKdWcegHHOfSer5dZhlq48bJb6eIHxfe
43MQzLkVHpE8+4Zc+Ox5BZAkFp4JyNLZTj3QhAVxQrJJ7T04d7R99FwcVZ4Z
242O2meakC6St2L2jJGBML/bKFp5Bfb6QuC2fiSCFHEWzDtkWT0Ld07IzqKe
y3ZoK7qNjk2DAPw9zzhVQwEKCX3IxdfyPc6bZepE1mvRm1moJUFbZ2aS7M8y
T7FSPtBlDOACKJynmEGKAifergezbeox1upBSrvB1vq1ydyZGgf9rgyPXape
7Y5+jPjh10nv1qedQi0afpRDd5OLTAgiQcThopOqVdSWZczUR7xFC0yNgOwx
PG988vIwHYdnvdz+OE/xNyzOSrjsC+rdX3QrRMLiAmxlZvXnH+XmvIZ5qYz2
pv0h8zMenw8+WrCaN0ixM5bBkQ4x/iYKiigoFZ2JDPASdEQGNRuS9JLPw4FY
NWGdGe5cf1WPQ889mxr6AUpoixyIy2brcYAfJPkULfrSkZJ4SP5poocTYCG2
jKC2Edw4sJAvl+/iNt5Y2r9c4rKnPdxCcrmVw1EDnrSQEglInI8vDclKeskO
dMeKEeYk7OD0+HjvH1jcZcE50UbRuSf57OUrnJdINKT7tuGuPYecJDeLJbXp
r1bcnfKjzA8+1HCO3K6xptx8nCg/zB0OE4Rm4UxphwK60vXGbHnZRQFzdHut
fAHaeMS2zTL0d5p1UK6mnbBsv/cUia8aoVYgN152vQ/LMIw1Fetr29rOrqeD
+Se9jr1KkkaBntp9YmRRvqega3QQBe1wRVESP8dwmGcX97SWcETjedEtnaSv
4UdST7ywOAqb25NV1E/6JZujTUcj2YQdUZKG4ewbBLQSc8WiIf+ZRAA5CM8g
KlGVNG7AG25U48sqd7TG8PunnLNlKZgWbP2NbO8zugpv1bje88RBraKUl+SG
eAJ1VIckiVN3d4xMYl+RVCJP51qB06Bzp33Kj5fyjhwvs35K5EGkPhQkRuqt
IAaZnTJbtZFPSMx6bicYhgC65zqx0WnK/mt9/YrY0EiEIxHUyxV7oo7i8OqI
WUsGwLpACQrPIsyhuL+SbguUqqC4p1EW2vZJAoPr2DS28ORx+TJObLV+pZah
noSwHVQLaLo3UXA7xOX3txdZkdL+1WqCt/2WobMn1oRfNkrujFWfo6NueNHA
aSR/JpeXyINhWNQY8O6ouiMyFfSQ5JweeYy9BHstPlmFGw0gyrzYBV8zHX8X
pzfyCapqrIJppWveKwZ8Y2of8GK8CPmKv4Pt75HnBgq+jydKb/xt2lSyZaCi
g2BDFOs9fRX6NWlOtrOSaFayt8bOr93p5/eSWOb15zgGrHPa8h1OwV/JB3p+
Yrqgn8VrQ+qjICLpN4pIaUgWbeOohCaRWtJ0fQIYaDWKwmq7WF0RUCBOBZ14
T5U1albcenZBhhlYPQOcjKbvI1Cwqir70UQhnTC9PEkNYNOkJ7cA74DtlGXk
RoI+kCOqceF264+DyhN/QttSqPXd4zKPsj2N3pmwCLxLdDRYVRQQYZ58RdR8
SJX1KlA14lD8EmpX1F3Cn8SphH/54C/Y+x1sbL1WVb0lWU0Q0dwjYuX32ezB
TVeDXYWDxdxSPG7bfzoT95jyVGy9gPfT1KSf1G01/pzd8v9PGgbKlTmP9iKe
+mrsMzQUesL1XM/lEeeM0dOEgDVbzb/2X9vaT4OfpfCPRWzdzYxC4jCBhW/r
elBPhFG9TH1CRL5Y5+ifI1VmSYIjLGt/xq5xGPldUQwkYQd85qtX5vwRblga
QKmE9D0T76qpzpxowvR3eGyomHD161ANZ0xLxukKR/73JlLJdXe7FRl9idcH
hFwY7iFdr9a6zxfPZDEVjPhbjK1cSRmOJmHxR1hVi6CK7C1SMiR7Fm9UmUE0
zTg5nGy6Br6keWVZ01UWyrrO5rGzFv/hAct+7hO2Vs3Id/AY89R5jMtiJSqX
ui46Hi6+7oEMAMwKFUeytP89LELBbD+T18lAPInk5PFqjIzOEJYPbCkPBHXH
10yfDEi2PJnWn9Lssw1mNt3UJhwt6yz7K49MC5bO4e45GTSopRQu2V8ZI5ir
olVwi5QRz3iwCcyl8BmaSvb7MgBvud+Fb/rguDWGLhur5uouJIdCQFhMXve7
iT+d+Aml02wEZrJ8w3xVnfPn3rXi3mNF5KBOLgOdOi4mnhYEboebVXfx1Jjj
Vw9eV0MUnM9h8tmLXxBEPnqfk34ln3mWmay4xI2/wZm0fO2NkySnjI4lqDtQ
Sw0AvqqMzxjXoCg7hDLV6AoYli4Zuw9An+xT7rtdQCyW7nRpi9Co2Zkpxeei
1jyinRe6fQXOVpxufA7ofGYAQVkWzc+JpmJ6CJMchFnbx7BK1BF40bMMjPLb
EmpxPPS5qLnoWe+GpevIeeAheMs07Fy4cwfwCDVb+M0DO8fIhEv7amFPGY2G
wLaFtrS1qhwJQm6sEBHbBtzaJC4R5eZuu1ab+UP8Wz3bBqFwb3rwxuq04wo4
cWgVkvVGTGs9/ruxtBE9qVSxrewtzc1GfAAjBPbi97q8CCffrkEPS7IXlEgU
fGF2HauxTt5YY8vEyVWeFbMqgp8kRmdPmnF1vFuYx8hPsqRtjIGF4iUkB3Jg
06P/LArLDu/GW24cmd/6t8Na6aQLdFuLVfLKb9Z4ZQxxSPT7n2CaszphTtK6
QdnMGzxO+EwpE1wTOC3GAK2kbShucYi7/zjlM9CV1HnX6y0MVBcX0Skgmu2q
eDVC4fJVnj2lvo8T5t35PSm1YTk+wjkRdJXJkxRuDCYU6s7eMNIXL0KLrjd5
kDFymwdwSTHXekXgLLn5Nl1lIVf/gWVyIwHtibeV3/j6/LsYHuXoL3TRD28H
BqfxvJo00HrwcbMTPNjGlr1ap64KeplRRspmrcmFdlpnlqh6zTnpRgngUsWc
+26wx8J4vRibPwSOO52vsTKtR5oXKWfxUEXadsLDWxDFgbIa4xXL4o1jIPY4
+KZ3+kgwhvifXTFMh8fDikOOQWd2E7O5yCU2VEa4Vai8HjhCDvhSAXbfMFXD
DA2Gm4P1E/hRwbFLfaB2C6nDRr7kjhyD0EwgvaJhu/hM0uN7eBlDgyKT88hU
SX+z7Lmq26juDM7RlBAntv2heNij22OENYnLww7KaCtqxP+s/fEWz1T1re6W
v/Vc/LilTewdnIhibh0UzcZDVr8RDCQc9pXBcDRtbNFf9Bbe24/G+Jsoe+qd
BcKyXoYcIPsixMe09Dbum0IMixvASAn/IjuBnr/wwlWraqVy3Totwy/h+VyY
eASj41AQvxzSvBXqVPXoOGBywXAnZENHlnyeeqrguBQuv0F+3daii0ojABRd
yWKyUiClrg7eQZXLxwaVvi90tb+XMXRK1ECyq4esqV+P6uYJEy6e5ovu6WIc
snqYeOKump8BbPmMc8CiNL+glNA5zPHykcX/1oTXqNk94JJnfk3CbNJPq3aC
xt64odTFhi2AgxhCBjyrxrAqz8lKppMHm6okK+IT08XRvIZ4U0ONqj1tAhvc
iOMX5qy23LKnEqWpKL2Uy8DWkDEEAzywekgzlhaOjUN62pWxZJwN7697VqrJ
dK0Zw/Ava7sQfQWZj+yeO2haDfGl45abB8oScm7+7VtLSLecI8kadL6Bj4ns
UWaCiMGpEcnZHWrpm/T+wjp8CkQbPGIx6FiKVCBhK5ADZ/pl7hxiEpBCjuBV
KRHvE5LieqQAQHeeWktj82x8esM14elSeqFQBgx69i8I++ObbWJAXsMeJVTc
9PDxzoSaM0apnIkC6OL8/WIT8Pd3gtttNkMw8wVS2Ze5qctx+FRlCqJxJHGt
JjZIYP/8mxF+1AB+TDscf/OwazDCQsp8/zTqmdptTCXSQUnKfIOCEivPc01/
VhlJQBERoJ+nw/gjW9Q8GOeQoZi6yUQn1qmogbgyvSWrSg1ihx0jwHNoUCjU
cUBsCQffsX1eqRcehK3ynMXZcx1vN68aC/Cenr4IwN/jMAJcIDtpZ1NapziW
PIZp9TDscmc+0Pb2/LgZrO093yuprTMx/EIzMUeH+sxelfAIsDk/hhVKqOiA
W81NWsQy4FhyMxGUEuNYojX3BL1ZySbFCCUZOnzSriunPNG2wm00Rzd0fGio
UXOqY//Znmp1w0gXvtyFS2ZEXGNJnAL4VuHW9AgZavNw4Mkc3BLLwbfIIwbK
Jpp6QQ5gSRC7cJfgGxYPP6XVhqWM+GhicwcCKVj1Me2aHXG4SBO7QWwVJrpQ
lKt+SkLjbLVIfzIq251pkDiJOCp+yI/oKWFHpIwSgWylOQxu7M5RtEFyIo/N
uIXcOxgtvOug0qphiIMTE9nUamCe85GBxriPP7LT8ew9sqX/t6JCaU6dU6LV
mhXgZZkaEum6OdIiqzNKaQ5LYHFm9HFsOoB/B/M7wBIDHxuG/GcievkLwyMS
U9SWh0C5ZKDW5uW7ozm32sNxKvDU2bzg/nWH31CSMT0F54B8g48yCpON6bgG
hSjr8xb43nZt578jo5x1CylFXCKOfw2n1kp1BL5xt0EympzP/GCj52RMjNf+
KvRaplJESxM4YrdmHChuf0u3rHaPsOAx4OzIAH4VXNJbgtEL+uDg4E2D9np/
8YfdLop7iYdL1TWPBralamWTXWTT0xXGp638DyPSeZB5/YwnNK0rrMOn9e7E
qSYhQ5f9/qRk6iObf56nBNMYQpIWDaBmLTgq7DF+RxKmHB7yaTq0eLdZsR7Z
rZ38Gkx19zX60QMIs4KPP5eyuFNmG1cGH8kJSIomAeQcpE2J6JkIKR8socAO
B27hou5IELQBQlnicMNn1Tvl4yOwFXvLbpy31u9JSlc6C4/DJfJ8KzKuAKVA
QtbFFHgEkdQxhDzybfY+ilUgbieV+kctbteHI8fNWJpeCRyrq8vpl/VTI2V3
t3DKhP3b6Cz3t+Z4RtM8b2opRRRuJtTLYhjLSdtM2J2/GMBnRMh6DEQSkjNW
EbiRdZvgPdyx2s/NnnsKmGq0b64ctEgEa9PBqTnb8xz7QdBpXD6ql/odzUia
J2eOvFsqy84Qvku8tJWMN7nVNACmKtxyi7ivMGaZAZLbXWgSNuQt433D3wMc
bidOZDbejG9r2a9jQGpUgnf/CgrNbKHZw1yOF9KBoGJNZq37JORZ90sERGge
Fw+bBUsWJEwxUknnJCBM1VC3ysd908aCVmdeNsG0prP5ROKPOOqTuNGwnYYU
ES5Z4+SxyAhIDRMQfWGJkV3jXamv23iKrjlkWPUR2afeE8qt8OiVFVnOgg0W
k/o6kGGCH/MPYTE/Q81siK1HJkB4WsucHSp5vZJhPDjrjzxbz7X1l9eRnjgM
K4tfdfkC0YzzAGGtMrXkJeBoMdODYFXOxJs25Ujp8xesGx6X3a2hNPnoArpd
rEyUzECZflxZs5d8bRpmrOHGrPt8YsFyep1qF0OFOY7VpFX70WPpj9qAmchV
/y22WxXHmGgbu7RTS668eYXMlk6xiBSgNR+oomtavkwQvik4ZmiwTS1WWuJP
VGwK59qIlYfdAF31t/XNdg3T7BPVRNtokOG9G6szbT6GSjd+2EuQUYolwZu+
YgEG6wQESGNq2uTqow3iD6h/SqT1QXpR50uyiR7Ni8CYhtGFsJrSU7rmf8wu
9sHELmtoYDHvYq2+6FjzE14otKYCPHDlJr+uGms1FsPfJfTp++oQQtWGEdbc
vY2WaVHGpeYeLJZzDD/gheGW1sIuTw+xhxqwh/vqMKeqUKS5GwunR+xZFNYc
W2c8WYsakRhrE8+oqNOMffMVtUs6yfjgYfesBPGGVU0rYJrKgVePxPuAlDou
wV0PJ7Azd/NsoKZmciC41lX8fXhyzktu3z62ENe/KrkVDY/aFKQLYDpVXH9f
X1TXKeIy3iq+fQdts1q9px3vqZ5BJgVbDZ3uzWAyW9SYQaYwkFjGd3pu0c/N
AE9XBkMwqu0kFqpwC/ffhyqfnfNdhCfNa6UMxR07RVB15UX/lzONRo5SCbBv
Z+tHmntGvXl3NHqsvdFsYS6EERNUUXlDxGNULDArSZf6FlQ9qZ2oR5ojDAtf
bXSvCmlEmRUxAawxj8GFqQmKtMAaIjOkhbI/bXojuV2BO4nP6Y2Qkct48W1v
MwXTTydbjQLf5rE4oymXT87NsOkG1rE1ylRFDM0YN/SVZPHioFC6RkBw5Xyw
5KKpMZtymXU7qySAUUp2zWmSa9Mxc6+FTliAB0oItM9j23wAtKv7ulcgCBBp
MSPLkfSuzYuHku/4jVAG8ATGWvkUOprCSWrK70PuDKJz9VCUiiud3nnofKM1
6szl7TZjVA/ko9O9tI0OHQcnHY08w99Y70VeH7lSunBWIty8hgO0lkmCOq49
KjG748vntKFIoj/J8hZAS4l7EXJlw10E/FIl7shlI7aWgF6LJjENtX3B+x6B
dGyD1i1QapKyndjWW1kiDIdCAq8vkRW/doFw7mCNkvRm3wINuJtY3MYongoC
v6+gIqpQwo7+RKnmQDZZBiaRVWMm6c9nbAUElZaO4nzG2VxQqC6FecCH9m6p
8nUUywgjYkdGEz0q6IQMGCLbHU51dKBWzG25GgSE8yq6OTndIihiZRC5Jtu3
8GQ3/2v5rNcZZmgCTluQphXMtwOJiz+FARYfXt1YfHxAV3H4nh6Af/OUG9+Y
9A0Zzq9hcUv25Gcy0Fby2H1W/eQPDC/kH/hWikq0jfcWhclXYJUVBcOfqK5R
ag6oWe5MlwOZHlc81PlrrBXKI2pivBk2fGtW5Up92vZfwaSbw2vJDuea6Sdo
JfxSNxGDOvVeZnfQPIsp2a31JPivCC3BguQKxxV/Iw0n/qD+1NWwnBs9Mow9
81wPx7w3VdC4Q1BoqayKYdIHN+A/8COAtJaDptUm4b9UuWtKSWtQ6jEW3efQ
Fl7AYXa9JWCRbhsNmdfhX96IsaoaucCjlypSpwzfO63Cq6nMe/NyO9f4FfJc
nGOD9uoExuRXPiMm7CWhN/KqKZP0RxP1OUxSzPoMHMCYYUR/BgKUV+aC3gwI
KggSLuKLhMbLozwo+K6EGD5y/ZeDhGlysVLWal0bojcZheWRMjeBBPKwVSEz
8oaW74HWaUhCsjNpoY+J+DTEtiDbM9CYqAtnsCRfC3EB+xuWY3vlXl7zHQZT
P5VngwpyVmPjXCr0Qq0/TmOqu8VwR4OhrvQF5EkQeZvuN46W7mC9LvUK+mFq
aYd2oeu+BGRUuzUlKiTL2jVMcAF59w1w+lLBQC4GZhr/MZqTwdePU8Sa1CPs
/YBZZH5q7BPxWtmeP+8LMyUG7YTV6DzJrBGI9nNb8vHzSqt/FYezu6csLvhc
wLbbQ6xVnZuFAUwdamw8KGACL2A/sm/Yg8Xvxl0VanZpvJZSLwaDNv+YBJGN
FXj5w+eDfvLzldqFpYB+JWWJT55nq6x+cp2zDMbOR6SBI2MCsKcdLWUQ6KP7
jC3LfZQiUMfOY/nw7BmNEhg6dr/vrAszwpQl+tgUGqjUKr9tlHb8iR5n1TmM
B2BiBWoWudtBUoFO91dleZJilgGO+DwQ2+cWuhNz8xAgBCR2OHVBLXXDCQHl
RCKyYyKhozIR9/94IjLi58yRJ7qn7yMwSuaSpTio7K47ohZ5+u6XJFQjebgY
kwSyFB3TLUOwkwLZLeyzOUTXfUwth/R7teckI/lvhVe9pEZUkweo8+BwPINE
QjwvcKkjXsmyj6F2zhkuYcEsMeflfqtGofKMcapi7DlBBQlRReQeIqq7sFNJ
fXuWKM8gsJhcYX1wy9n7UK4tUYzgpp2Nel8txabk6pUIPEbdBt+dIjG455I6
gVdbdEqoXK1SxR9DHjMMMTuZGtJB/vrO3FGb+Bps51/SwATP7f74/CyD051x
8l79RSHhGCv/emzuJFvguN0mvRAR/I+xKdUm/Nh691SsqJZKPvVtdqcpnI5t
h+jqVitHzgYSyGBWwBfJXSoBw+6NhOR+bYI2ULj5ixHn7RbVUZi3knLkPfj/
wgGfj1xHdQ5ivKx6EMDxeqp6uDFbIGeNiYBnB2HhkFeJbXj3YKAXq7rh770i
1qNqPMXVCpIRfSrFz1fDldGhvp4rya4Cecq5n4CCpem/HRz0TC2ZY7aehH3T
sT7atpy76BQP4n8ttye9sjQt+t+ZFzZ1l6f0n0kyXpDnkwnlhLpb1ZvAE49B
hRi4LCBqMsp3wJLHIUiJwGeuMKTNzt1YqkkfVxhN5dw3WPgCU0A10aePLlOZ
mkIabadtvxcAuls/60nxv5IfAq1uq9RjtsDRnj/CpIzw9K27YidQDtG2DVMx
PFPoZr2J0pzIoHGyFVEPVEVUdce0p0O+gV3/U2PKyrsPImO7LQgoJ0D6VRKh
TGogNW8rKUyGxYNhNxPDY4/7EpSiBPAmnx868ZIoOMyvczqGg/SSVceRykDF
sDpIuwg33t5vnJmx0S0Wxi7gFrTtlCvTrihgepsWfcRpjPbzQ4mWDFfCh0oO
a7ylf0ahN40KL/9RJdUU8teLxGRZdLSBq230pWWbI/rbtADug4yZJWYd9Muq
WEdhQF1x0Hqggvx2Ksh+ENDVQGn+jXPSv0pLsD5Ex1Ps1z0D60ZAhbpMX2uk
UONUaT9kcSeB+WaDgBOMLx9bpvK0iuxBKfniYAD+jTS75oqQbvL049LGyqNd
PuKZaBhZrbvwqJhM0VWfjhL8WtZgCtjdeYQJftV4Kdmc04OfdZQk/owTZdss
EgnEBgC12AsuqRTywlMdSiqCT8XG7uB/KCJL13UYSxvVlRrjfiZX+e/N6kMn
a7WVrfxXko3agWHTvvQVItwsu7Mg5qX4fP0KWf2Wn6zNQO8PJc1jBLp6lWBl
H56+VHkS85VPlHHVlbWomAwsgfNHAVgklclMmUW53Sc5Ssr103lmEwacCAzu
3x3uKyCacWIwqMoTerAd5v8rf+ldDSaKknczbjrBY1MHGdlzXG4cedMFBEKC
dOiJwDNwfhkAXzf5J6tGCaJk/Sv0NgQ1uLYtfb9mDkjH3VT6sdKaRtWfOgU8
8siRxSfTwpCbtvYceLMfDghN8TNjw7ea2WkcuoXTBaUcwCj/fhW1zhxDeVxU
dnwfjneF9dcbaGqJ9WxaICvSSGxKmIG3HMuScnG8WXWmS2xlaWVC4cpfTW65
el9mSV6p+0NjR61G+caWkH7aeR+QTiydcVewK8Jvu1evqdUl+U03AFchEfqx
W9Ez2UwX9L1AxobKSY99Xo7ff3SittqYjgluGggEPUrwpWP3UGlQXGJzg2j1
VeEXH55v3Wa7YOE/sshVjbWnV8gUF9FQh5FGjm/VdB6pW6J+432IliBN1vLR
XqPU7TohjgfQrt8cpTdRLwTABDyY7kkBjaaJdvvb5vbD6hoULNxRa0BD2Oma
7fH5XLrTVkdfx1dZdURTSxNtk/oPZKUEEowmESRHCAl79T6DVKuBnAYo1wTH
2HNrfX0ZNbynWsQgwbgPmCsHj+xIBDh46aQxwqjZQeDc8UdsrKEt12GN0EIr
Gtq3/WzcyRUfkk43NRLTQjg94Cn/Yapbi4iYtVUZ63Q445Hm+TPVjmQT37/M
XlLiy1kSctrZcOSTzYiibm+mV4htifqZRUWdHVhJ3O+zECvbyNcgbpQFKhwT
+3WjIFX12FPNqgpG127WraDe4NIZCEqZSBHpjNmzKtV6piaRjY2xG1pU6ImR
xQETWUhXfy3QfQAxYZNm4+eiutE5LWbAsQ9Wg1aG3cP6YYsF0+A0uVrf+5Go
9aU02mlelHVv5Jd2jLfGUqFG++uZMf/z+0LaKpdgpF8rjBA/vuw0ToVdHq9v
TfBYfeB0pc2zfbGN+KdoCis5ycUVZo3GfiGxgoFUx6XrpnemJHBNPd3xAoVW
BPHBW/GAOenw66mcqi6c/sBAOTEN78Vzk5lC6l8KEErVWm1swN4LYrXGHO92
osDZDl3y3TrAWCyqBjAr4kUY65S+MV9SG5qcNsnLSctbs5jISObgQXegRyPm
CBKQBPtyr3aF1l2pNgtawX0XRpbDVZfu+bDdOwD3s928L+vwYqz8LJBYb3mu
BnXQbmxFj7EeBunS4H27hlW5+unIjDOlwVFlD+SwCc94AEWGHH43XLV6ty4i
c1/6zBdoAbix9CGJa4HTCGqaGkl7fKl0XlIWCJLNqgJIjFBCzEpMzwrwtccR
DY5illPl41rxgFZniT3diHreP39xdr2vgXFAiqsPKkCLS8YFkh4z2cS0zj8n
WXnJpII69r+LgaMi1IOkqyVkLtc+apWiR8mBnvDmKbuPa7pQMSHR/RJpBeFu
Zmao1AL6HCOtrKz9dMThbu45vg9n6PVo6/yJgvzD1JDB+p/39XuVAHLcul5M
7rJWCipQrX6OxIJ+wHpgZ5s4WveJ9k4/iUqNBRz4AOsMM1I35ir/eG2YO+eo
D4azodkPvCmhHLQ+Ehfh4cRJwUXs2hNhEWKhXv12A4LPqQwd7wb8t4TZ/gEL
OV2TK5q3T3LS7zKORX0F8T/K6WB5IuoJebDFk8EmNadu//FzPvHnb0ZEibSb
fFvv17TCdMukP7xIF/LUEox7eU4kUTVgcWXODCxggasa/H3pKTjwYvgdl9um
b3s6oln0nQlSF/UAuKC5DzuvqlNsbMh5b+Supudhy9pxSGRBgrSt+ktwOXpY
x+7RzGvkKIi0PGp8/U4jKmeJM9e+Pbb5N3LPb2qElxftlBoRgp1QDimqOZ7b
6LHflmmmbBJ71D6DbqBb2dsl9Ah5skYgEeF1a/IrW9ut2AfIO/1vxtlgtFIG
oTUUHWOKxI53LjpfN2Rn3ftaXgyqKMhgaeJm1MvLlL15HaKQhyt1fZSgPqeA
L1YppkfHZlP8yNjzYlw8XDrS1ixqY5TNUsYzTgcCjB/D0llIBGd2vNkEZ6du
Tai+PIsL72l0ZJENRORoJnTLScVE4Lm3y53I0z5p9r3COzFTn6J5LZHE0Xy4
SgzDseVu4yjIDq/bbLld9ONLRNSb5fFEywcCcNLzw49wHKJPPDS/uIHLMwES
3f1ce5b2+6wIIsi4HfAip2aeJNnY1Rq9dAi9T6cFdalXkwZiz3l/P/lVsRq+
ySSMbuz5F3Pqb+b7uGNd5Nw1f1r/t1rXZHKbOy0Fkk6XIY0Bv8jaXlYBOx9H
AeF67HuiA6KK3YexsqKYGxZy0qtqE4OzDBO0LY+XwWSlLye/7E6C2RAZa6r1
74PxRFQJln6syrOKMY648Ml8mY84NIUoriwBc49NWlJicabJJ8BnktWB0X9O
djI07nqhvhAV9Wn6Qam/lY2lKt+Zv6dlHHsoFylWkxnpfGcnQLiDXMMJixte
ZnpBjK0iCHA8saqgR0ldQfH6qqp91El88QNQD4h68WhvHNqFLw7OqI/9MIdQ
MOkj5y3DELa0KfE8/ES6C1JaDoM5mqtHlfNf6bRyKfHdeXmc7bNT/I36RJFk
rkI1MuaokRH45zZxvF5g4qw2RtFChSzZnLFSQErr8WAVta0C9AtMN7f8+vN1
Dn1CqxahwpnZ7ayvnr9g6pD/cmbpGfDiq722DqtFNzBIKyft5NDCJfUhtxlf
PiZ1lWRxGV6gX4egOv0bxbmZc28qCxQ3iu2yfBv2yQ3Z0dUGvYyLuclsDR9m
V7TDjB1pxJip25l4Iyd7NvySnA7GAJ9NLvM08Nu7S9y1ylIzk05XSQ/ubUyh
WSWccDRW+CrJlTiSfhiWTKWC8zlyL7q993Nt9FPkSewlYypK8eMcU5AqucEh
i+kbqplkLuAf/3v/I2/Gpd4gerWcY/+qn4+TiLSN6GrRCppZ6DxMNwWdHJcg
uZtfhepvxTosRZ4jZmOC08He17dKwwMuV1Hq1lIFJB5gaD8+0iGAkxYJx+us
obvApO5A0ONtTRE++YK8e2L3T/8xQrqgt45z/GI42GVoYaNC7GupRkCVVX7+
u4w+6JpLdnPjH9v+1c1tCXzMwpgwZx0o7KUnF9xnrZ8/lAeFHHD577LRLr/2
7xllfhaJe6PwYhvZol9FWYsNxfp9ggxVoTDRT9xSWXvmhtaMcis+TzPzKq2E
9ML4ZzBvq/ugNcmz1iJ69jh3DoS4PPcqi+wnJlXVGmorwFKyoEGhjEcKYJTt
nry7D5oKo9desw9/YH3AFgUccDPwCWI7WYh7OfikZJnl3XW5HzFjxCxQ4n45
tmyOPhgMUbxhMkJp1pmqV7qS9Dp3McDk4eLPvtVm10SyVAz6/Di6oPmfdXsa
0Qb0/QL0QQ2cgsCCdyN4X3XnEbB8z3/93aWOhhpi2pvfRZq21JGhgZX83syj
yZADGtBDN0DbIJHKeW86sayejdGrjATa0g/uUJbBw4Sx2KiKYDdJOVhXFVws
p8Vqs8JdIjKFLdn/Oba3yOmnIo4TCV/Tkj05rq/LWjJOBUObg7Ybzf1ZfbMr
nVHOfGFMn3iJY2rio//6TKeQIoWaaRYp+WHT4d4ujvHaj0VWQIfqPgquPgUm
X87RN16EMUrNwUoqrvlKZ7zzQLaF2i0ziLB1G02a27+xthTz1/n1Y2B8HQKe
fwwe60Cs1JIVgFuC5VjrKMcXBFkfh3RCwyAdqHcXb0S1l/Apf1acBgM5cQRR
d7pbux6POQd/WI8q4cd+hXndgtTNBqv/CejhfQYpX0nCphkVtRNhfJof7qhO
UhfatWrzKTrQVpdZFKxd7Hh1YA0rCDaLegwHILGYiPuYBH5/tOYY+tWY2aKQ
rlhhk8WhemkhB3ihlID9Y6Ti4lTIMmugCAae5llpUn+5fI7JjCZp6EB9j4VZ
Ea3Uzcs0Kl59c18fnfabHZsmOTGo63bjYX1xsttKcZ+CymMhf0Se99Z9tfH/
T7BXlSDq85hylYQae6XXVuspIntyN0dPCYZyZzoTLZ7QZA2p02uT4S26qo9S
ZC4pFITZVQHNkYntwGeX9KnFXkUwrZFi2KbvSM2QsGNi3s+ctai/TqgCrD1n
ETT9vnteBsUs0javYR/BNu2ZbCv9BWDFvRqsb1vznba3nKlm0tIFOdxE9Tgw
cPNOu5HD7zAUbYnmPc7jSVOKR+Iq7sXsoB+2TocnnwNmV6/iPau9rfs2zEh9
0bgWzy296InUhCbr8Evj9nSHtrrfE3G8EugzCRJTWZjjzCbewspaW1LvyMI1
eKPSMW2nGYMv38rA7MRt6U+T211Usf/oRCiWj0Up132kpkxQOsOy3B1D1pBY
o5B0W/89J5+PlQ7ibwhEJnrxqn4k9elspnhZmcdvKs2QCuPgfYJXj00UWfGt
EyGlhDqaG4PS1pe6xyzrJh2plQzkuWzJaDTsy8c/CL0IhQFfb5EVoCPcnyIo
s8LvIx6C1HMxdPMm1xOypvoELzGDMMWYsohswJArBfajtDqJLcnarRUDfuj+
ZVIaFsGc0WZvBD08eVfP7msU7i2Kx32ZwvqIhr+HW3yVfQz66jbJYK6eJ2K7
1osH7Ml36JNrImQAs2+xjrKrWxIkXd9NYTok1VIMz2X+RGicoU9eWUlFjRcq
w3FJ/MLXxIor+yh1z4mnZfk59hmUt4l+i0zAcCdsj1hQ+0a1ElEOglsLK6Oo
pT69ce2fc3im1j1KBbayO9ewMjH4J8af//UrcWznIf/sTUgowN9wpzTJraRJ
DwGe7eStn0r5bF03H9mh2J1tJimrjlFRsEMIXbDVSM2DX4f4G+UqR55RK3x8
Hkdzbn0d8MJior25Jg6sF0bqVQCv2DgEmracQGIkw0sesdpH8fg7q5j4LuKc
oeblcxlyr8xgB5T+kGX5uV4jm0Owbc1kfgG3Nt2M8LRu6MCeN7rK20cDGXyf
zERUt4XWKxbx98Jb15tzXkFOoZyjuhFmYogzL0eDlTXzkqARZ1gNjzcNrm7i
/mSxCIO9sCYEHehu4HmBTLjPCkO9ssRDop8u4JMHpaP1shTJd0X5mVGyAjYs
RAGnrRbe/Dl9+zVSX3vIa8qmMPg5H0uhYhr2dzEQThIqO6eM6No5Unsz1w9S
8tZWF3Wbh0CSN7Dj9BrTInrhjGolrBTqZZqPVvFMvrEgnqQnbymSQTyewCKJ
C+cdKuo37j60yYq3aygKNA49dPRJvoNpruac/eFcj1zyORWTGZlMmEEunbog
pzPArg7RfK5QoeBVKSeoWdhZQtnaEx3/9QMurnUirWYia/R9EN88gmDG7638
fSUJGiDOpGN7JNWMNI3pdFATmFSHHBa0JqXbP3Jct7wjs2S+f4r00QFy4Bx2
KF8tULfNatpXk3drMRtpEDDC81L6adtVhG3F027KuTkKY+jn3yJFy5qaVK3E
ZQLa4b5RNkA75aTI8o2z0B+iZ/v5lGkkrD9ZxivrLbHbHPOWwNpgM5K+WKEp
fJmHRtRLmqe4IL5I9j6nccHO2/pQ/bz4tp6zb/l5vcjYSX5TfTthobvD86f8
5cbSy/HU8laonCd/qzu0Dtw+yye/iFLt9r2tHhe3AXcDhDYF205ZXCnjoS7x
rliOV9VRu9iQCWbNSHOtPWgCKSns1H/Jy9Vt5lr0j9fURcIKt0edhiPePfWa
0JlGW8t3GMk9opxrrNueaAiBBnyIs97VMVq6cCsAqKFueEL6Z5gD3y3LKskd
JwG+Qu4qw8t0d9Ho/SKx2LrNgdJO3sdoUg1eAaxEKk3tTTVjTlQ7WLcOGf+c
yYL9gEa3/xns62h+SSUsEriK4E57afiVpcSzDJ4GH83EgN+1UuWP2pL1uFsY
kfgwg7/x5sEC80N/ffcqueQVsIgzzWPWDRlz5OYl7jQdolv2/YqYb/FcSspq
hiBHXm3JDLDs0V599wRiSkKZv/DA5VpPm9p7ea8a2ZDwFBIn3F6tKg/9SfZJ
O8NjUZC+nIYO9fJLNCTUlzWW117sqDNzXpUwy7PprbSYehrm75Z9tD7IWPJd
E1Ym+pryzdwfVy5UbmyciBv35mzcODEYcmmnHyXwjJIbuiQNNBjN4g1OhTPN
EZrbSgqg53ux4QbYuuAInc80xJHuGCi7wLdZbKuTMouFXHIq8EawwMwHgF4x
B9louv9Kq88ukSs/lSTYTA4hsHihj5cnKPuOIVgnlUZkrt1qa6QBP+rFk5AR
LwcOgQJ5vxWEVUBJyCBqE72YoZR/+in7WUevRoJpvroBW5spsj2jbREJ8SDc
pPAZLBqQzkC7Z+27EML0WOMiCNip1D0hu5gN4eV+8aCeMTBLhySL5pTGXnYJ
ZWrDbI+gRBG5aly/JeZHl5KJsujv0AMYzucxBj3PhGEvhquSBV1sEsiEUVlL
eR9wISTWa1Jge+xpuk2Ca+v6At8CP59/kEQj7/Z2TNEDKJjcXPBtU1fI/6H4
wxuBFbVoZ/e0JqbTs/TKd2Kng5pb1Ep8kKQydKk+eYXrDeBtTKWl9fhoYTXq
z57e1fZj/FYwSYQsDy5FPmlKLy0jNe7h/brbUMCXcWf5pS/Nk+5a9TFpqsZE
OtRlS61rt7cdldRHFHC1I53zPrLNqmwtehr1UkbsqeY49buuX31myu9tyakt
d3UzFleJbHou+8bfyTWTMq448EehC9boVSo/XLIDwn49Es/tfAogOB+FQJX1
pz1kpZRMYMupmmsnILnGgX2Pl73qk42IZcNaWt8TlCTFAsAHuy56Zz+wtFxF
xZ2k+rMBTKkLEUb3TKgoqg+qhVQ7b4db3ZoMJJ6XUUB3vWo76kxQi+dZz/od
RbOHzaKTcDaQOtwFME9J/YI8gFlCbdEgq9czNfJzNTAyGZDc8zq0dLdDiIrf
aPL0EOdUVLY2WJtAncgWgoLFOLawOoNsUpztCwBgkHu4J6YYht6PmkF9MGCt
jBqSyR3cRi66tVrXPpt1qqwqyADrAUJUX8WDU2bf1pIl3ngoTcSsIautaL6d
7QrZGTSlL2YFGqAdmeW+v4/WGLNSRxwL6ycEGCL7v+sSuAeK2T/PUNvRsvpf
bcPmY8QcF/E0FJSsdMVL5fnDpTKskjq2z4wYpKku/tYjR6up/QXEO9ibtQEk
+g7vL5fuWLBpdPcWHlVQ5B/J9BcsRHY6XPpb9qFkhzcngbJoRizxc9Mtww1o
WySr9vZLQn5xya3Lqirx/WzdkH/vKMLRWnsJKt4tc8qEiwD4T0oAys665ZcE
0SAOU7ft8XCCauWsgZcmFKvg1DE+4/zb7Ls3YwLASRq9z2JfqHqo9Vhm8wgI
8YhBPay3IjCYqJun5oc23lPhx9VQsQUXpzhkudTqZ+A4mM7O93hvyG33qJcD
T4M2PCle6c4Lx3bvazpGADBJUKevgCIKh6ew/o5iYCNYMAYTJsv+4j7wdFOC
fb/3wZ/VPiJ9s7d1iwGp0Y7reAw70U9neRmS5Jdgvb844WtBsrfhIL8E8/pY
TW/pviaKjSA3ray/H2Q/LCbEk3HbP+sKnD88f9M1T7YUEDljNRI2O9rVcJHF
xz/dvYV9Pojus7h8r4ptVaEoRO/b8pxLCNTSqo9BI9ZfnwuzuD7biuM1I5oQ
AFK96Bx13rf5vSDEX5usMLHYopO60QRw6BYm89Qc46rY0USX4NUE6nBZZxvd
FRgf9wRFsvez9IbfT7OUcSOg7x0Gpe4GyvVgmRLcAhpJir9eT4Utrg/4CClK
bUD9SVFNd5cxiVO+UL3gGiWLk6TG3iJlJuPabypRyZlUPyR8LkOowFF//CMh
//F1bLv133VavjDaa79dW3bJ8FkI77lncX4cf43trNo4Vjur3ksW7soTY5/7
iwzfzaz0xGbAkvauIyCc5T4sPUOPG12pElSH4b4kQ8KP/ghlqNtMx+DFgV66
v1hE/Hanfds/rVQzXHtqXra832NCEzUuegmrQOTZb+m1PhCaHJbVmrOHKitN
TRuYXpV9BNoeaRi+wywFzlwVOrCOpVOUEmhXnTA8AnQYv0t3zsuIzhrUUB6t
IrQy569SCtmT3peRLbrrFXmzBV+yDOGgho9aWwyima8LRC9z269MsYtwxn9o
YYlyV0tuM+MD2lGaVFDDi+NeFilen0qUAk+e0qmtRLDnk2fm/9bMBOmCefbQ
gH3QdQ6P5mxgFl2yNxh4s5oA0YKInOjEOXqag8kgawJ2qKmsEdTUHRPVP+2/
rrCEa08cHqDdL/Y6IrGsdamURJ/i3eTwNLIweMnFQ7jQqVOTkBD5nBFgfTMt
3U2gZOvgJWfpdSDc/ur5M/R9b6mCO/iWeaUvRvuX/OUD6JYt5weaad+SZkeD
7gsBH/rnP03no30cePVml2wKcw/jR3zHSy8YPH6wMTq6fQyWFLtai1PnvpVB
MWHOHjWoESQrga5cmu34GR9x4tmb1HCRM8oRtS2mLjNltstTLAQ1jAkeDP3+
duHC6NsO1XbRfie9FTB4FGzWGIlxD3GKh4ySnNLYzVMEigs3030Nr0q4G64g
t6AQguGeo/d6vMGPAEV8dH7XZmtOBb9Q8Qs/7P5VdKi2f2ymJVSZiqmikjDJ
cD8LbLO034hhw4/AG9HegA2XjKd1SbsdG8BKJzjYj2m7PQne4cp8mCW0Q/HP
0br3KB1h67lF94lZruUSqgJF6q8vmOx7HbrF5RCvqCJQq9RIgLV2EI1Cl6Ht
33j1SswzTnqYo4uuGE388g3JVg+cW+yktJzMTY0UL6owGE+FNF1J53OdWqSs
ZMs3RXESQVFSyc1YivB0ED/CjzodHmTRpRb8KRp4vLTk/KychkI1FsnXIpvr
4wgtaOmHL5nK29QkF2PDd+nUXP0bqtdf5hw4chZR8L1eFG73gDOKrDjwxXsB
WWj2hJ1ChAItx5WYmE4TtlwRLTKXbGBo8pj+4UJLlCdqOVF+SVqLIEmi8XPG
QQnl812pT8k4n5iLFenzecSsvOp7VNWzbJC5UOAU6LMeuSdKl9RCb66Q6r5t
XWosd4FeELxybWK0k8Y+XRgu633jprMTVekoiR/7/NMU2o57EJbU+3FljSSn
ZJ/eV/pIbXXxAdrZVblF4rOT8c3paO1LgdsmXIdnmNFGQUyMdQCd/NDnnbtN
88wtUqJWrw2h1Kx8AiP3TGvFITuQnjwAdwjSE9QD/Jxe7pySp9j3eviaTcVb
wQ9ftabtRILE1fpdLE/KANicizL/S5bwSQ7OwhL+/YufKoodvYkKN1iKyn3o
tXwtCJO7Fndeaz90U5pmRnj07V8zpfk7yfNfalMrUSXtrLP5ls9mp3hFN3vN
DmBUBohxNQSa4G48+Q7BAbysLuItcCKr87U6qEKIJMfKZ3J/5aY5Hiew1y3M
SA9YRtossFNVH/DmaaMZazC/AKl7mAKdwDjugvwAkjDjAjL8tX93wxne1J8k
BQ/CZBTm/GMgfMFfr4w6SCc9dkAN9Md7pQdbm8yRLM6Hx0Sgg4XtQfIwZ0FY
gXD+uDoCK5SoHb07BkrZ6kktEjhM4Sitnr4/Mhc1DvkEyuF0w+Tk8PudfmS1
yZGZIvgYjQxXI6XUGJ5CnWFH1xc12rxKMJQ+QHmkisaiW711y1MUSqvB9yY4
pacu5HsFIpaiPVzG+7Y1vkrokuKESpYL4IZDlS+mXHIZIVH7UvANS1nOwU/Q
R6LqhcFW1xKBaP8Fo3qwrQZj12CscmjRlB8XzI0JHzb7TWRTrEJPnFwXXB2q
0OpECBUK3f62QHgXNbt9g4ToGWfmwWeuweHOnF9XIFRN2RZiWpikC+hhNZlR
z9W1iFzhkSZq7jrXBvr2UPsmzC7LMX/RUEHG6R6UtoUyWuI9mZp0u2EwvOFR
Un8ied2n7olIjMwTQ8NGYYnAA06QogrWHRtVe7EpL6TtbAik5yDyKcm6teyp
VhSB/SFlZpWWzDu/EeKolPImFOi47eh43Kz6eHt4iZIebwJvC9NrWrTKFlM4
fBhroqcR1tq3JPZ2yz5q7RJwxKDWX+dULbhezWALjyknlg5gKigymuvyIzA9
hVaqLPNhjqof9pTNbRw9fNuAUuzWlUMBrvTYIwnAJdi6bVYatFOSeuRzb6EM
X0DuKQZ+3aCXZCCjX81/tiV8/JYDQHkk3QVvRFSBgwH/MudBzlugmA8il6fz
918KBF19BeFWhlKPWHA9Mlmtj9CSxTbp5WZIgenvllRVmUUDGXtOPj2U+W40
I4PTV/Ih/Q5yPuZoiX4Go5k9p6SPCvPhCIyuCIf9uhtiDxwlz1VMmuELzt1w
xKhpdVYOgPixNEkW9mzodmbE18u8tNdNNK8/Dz1N07IkwkL154AVlxmyIyyQ
E8cR43BWktE/3FEH8dPghioINT+98OdMxwVT1ubBg+8GXhPwavCIgvbTGs8m
Nkss/nk8LejgrIs00jNuttkwK/6vvv+xL7aOzr6JILX6hFKBm8zYZpud2CFs
eKOjKQXNblkBPw9+eiikLT3rhHXEOwaRqXWx9XLprbr56citfUqDmi/LWKak
Ao21iiFmDyWuzbxC5GHZZOFu7Kq8NmdciZx6S7FABnVPcLjBqEdIx+Rf5pm0
+1J3LaSKP/RdajUDIRMRH8TVU7s6X27Kp7VWfqKGcCkejOpc9fJ9TTAEA8n+
g60RLXR5/A1G/WvUd2W+GUqcC0CYXKnCa5ZPz9DSsIT0zLQmCL70BoYzOjq5
bkDuSjQ9E9IJluv4Ie75TJtHslJjd+mU3RfjtDMrnkBga8DWpT+0SArWAk09
CMR/9JMSxxTevwVEZhb4wHdYAsYZWyjChnQLgUig/LnO1d3rrKcPwu8C+fHg
T+C9bAs44D3BE9ZcyEO47SFQ0oZZ87VZy3MNZqH0Sd0ea6S8h5z03fvS9bMU
egRgqhAPOzlskus/TAxO3BimP5u3LXJR0/oT+AoRCB7GtqXYHfX3wgikn3US
UpPO+rDckdOREsWrtEkcN6PbyZAbW9r3N0K+SKaot4mQBJW0/pwCqTKPCnuz
xWNlNHv/VUwBZVh+GbheLbBb6aoBen+ie8pNw24k2ikgwAUjKGuxkPCWMV7+
toaK+yRKOjBKo3j8A5aaq0uO0pvg10Q/E8daO7oeIQC4pXSBj91mtezvIS7z
TC5d7ooO4RFytTgT8QnsVJ896Rm7QbdUID0d96VORKoJJPWxAB/zgGUVy/Qt
8Fd8ECpOrgaM5FOubUft24NIDYJf+LnbWWQ75q8jSopSma6MV9dY82jQ5IKh
btPwEEkTg3NoWqxtB02181rKn+jx+SB7H+l2hnKd+opJpM5MKGef85XrXCTe
4Uzwi/aaX25oDMjLqFowk3LjNajvL18PQYEOi+bjP2Jca7jRLMZgYuNh4TS2
Ka7tr+h8V7MpLsDxMhSzk5wb3zoB7KQohkRnbvYbHzEnoiE6zrfQJlJIK4zk
WIYflTY9qRbgpSdXZYC7vGdGpNWkWVASbRjoaWAr8AY+tRkEBbaAieX+/QwT
xHJJOIEtGYroIJ2sJefjs65BFY90y10pzWP6t3VY3/Ufz2CCTAk62qX4KV0w
A7LpYvlZUG25O2G1JLuPkxeKpD3wQteCFLSKc6hf2lFkkupBvjbaZy6844jH
3pt/ROMEpQw/XmNtXpK29Y0Qq5z2K1WJMfvnMvn3KWlCdRKQAV18fJ0cY3r7
6cDRLR9CmoE/Un3zXE2/QbBQZ7bdj+gKQa0Y7ctSDjivdeKgd0/L4GSX50yz
QFvliNBnzD4FS2SQ5fK9kaY2t/kM42+1vA539zr4n/HmZnVsGPBWXmouHhlh
yc68vGiWzLbcEaow7qFbcQUN3R+e9VRwvi71vSmLcRu2x6uJpmfppOz/oOVP
dry7SwdjdKCS0oBCDgizJRgAacdp8p/pe86ZNvCdB0ply/Ni5v/h8DkawQHg
/h0n3mZTCP466AVf6xf4dXkOuWrQ0EZJFuYM13S5CJZhk7MlEF9OodJcAVgU
aHpjukrTVLiHx2jYAA8JhmJhzGi+t5JHavdsuLRZropg8CpVNClp/kVXc4Wl
SvV2dFh3aAUzOzHyVHTOR/WZ3ggIYdQphlPeOS6uy79opgVAqMG2dymsqhj4
/lxgDi7ez39wKYxkmNPL7xjR9TwSwaRDDpopAjqYnA0voLp1naFMY6Fos1Hw
hjTtdP2iEERduYTBiubDET/rl2iDUGsu7tzYpiCc3AgtT0p2DoXZ/ZZQ+zn4
bHKTEEMOtOPEVMEQzFxIMEqYXSPKnvNUuHqcb9bYlp+hxtuVEmD+p6dBLH+X
wWqlnXWvU4rcooMJhE8uwc3XatENtDASBTf2j2VHbgEGcvsgW0vT9m2uykfJ
PSBR1w+nwlK60OzuaSZ+C139l4fLtR2jNIXsMX5UYUHSOtEI3Mx2h2EWCIrt
JG5Pd521N7QkpHxpy3L1N1Qm2UwlLNLqlNqK4gPK491gFEeqkS+AfzTPDhgt
zidTbrnCK+b0qIPZa7+IjMBX2EjUYCgn8VUnUWylZvBo5s4LcU8jPwzrw3TF
BYJvbn/cxTn1s/LVXiUrsYOdyyk1skM+p/+DDPgqSreDGU6AU2jxhzL4am18
XeCcqZggAPdy/8Hn+Tq7YrQr9malEHlkt2hOhHkyE8I5SW07UzmDEyHewSwG
4GhhOdEyCqqIAe+rfu9o30dNcAbqTLDEiW4ETV9xWXmmFuR5Xowqb9K3N+CA
F4firdhHyfi5Td7W6WPGjNA9jmt5crlvnzbvv0bXi/neSZaq/Zx2wluf06Bs
zGqqvgSRuTa+xV44+MrsI0ND1Hj5o5yMd8FhRn7L6CaUdlpE03ckuXn9mw7K
AsxKCEYUStLgeNVCn2mMIobNaDoXefUKtueirF28J/5pQU/loH6GFh22by/r
5LnQDarI8UAODsJ7jM1sTX2xu3AmjSyidq6RrjVm7/+ENSyxChNcBV4zAJBw
PfITnLXHg+s7sq6R+ZI8fEyl4PIz8zXT+FnKScWJ5qvDIn/jaHzOzPBwPWV3
FNMJQYRAGpZgLzaqzuTbRd4BanhhMwGzZvpxvhL/UtL53Qg1VHi8cwJi/Csf
eK9pJTvrBRlNMi6ISNMpKIqgERLpwfWlDCqjFs/BOa2m6lwOV+52hx3IBjHo
wJTdKsemY1v/yroqXFVCAXIA2gYRROH4c2gxcP3YdAQ0jVnu0wyyy0OmNM9P
h1hj3b+RrYPh83snV9huMgpnbdiOD4D1NpGMvstVqph5rXRvcyfjgXjQwe0i
2woQfPI5IcC4P2XfEhpoQTweVzLkfpVTNOZr37U1iqaqgtovW5EcxkdWuIYJ
lPGs89skvkHOUIvphl9ETIR2EUt8Y+7hAw3AQXoEgIjJGW26ECXLRKaawiM9
vV+XuKnx8Rx7FPL8Ve16LwG7+yOZ6Hweli1Nfwe4uiPGCcVRhLySmNP3znPF
K5liayE89djZFm7aONLd3yQSbIR2xM0sSVI52m9U83CQJ+wsg6XnyI2gIZAD
uKnVZBbkyUDq87OaOms8Y0gQEAGAfu67a++KSVl8RQNLI5JoNSit/8Wjjwz5
hOZdzfuDF7xx2fJWLml8dI7717KsfhD2fOpN7yGQGUJ2HGZgai8CHQL631kM
DhjR+2qZh0czK5x9qp4nUiyoeqa9etUch3nOCaON0CRurvZpvqGcc0u+rO0Z
oAZWo9xVjSkRVEsVtUXMnZignoYBFCjio1si6qMtzvMpWaGUEvszwoJKI4vN
eimwNeydoyZ0Tgqf3Xn5ITnzkawUzBP/VBodWRfDu94MB4CWUk6FLPAGa2Ay
2/FF0kFVW37GvY21MBCcbF5ictH+7x+pHtEU6qAnEUkWR1Ym+PAwTqWWoOag
r3lcv0iZ322Xh98rIsMJZ312SSO+b2mLFp3j8T8RVytgnvEMHrIaSJwdwxn1
g/3pCClGbaFYIhMsWmZWrSfff8ZU1+gjM8tIIkr2w2hxRz2mjsbt9pmyThFP
jqg6gQP+Gr2Uvz2/CN2p2dHf8pXQkmKLyJgCbvDKfjlIfx42WhMeHvgO5Aeq
ubGzHMLm6Be6gv6PruddBAED184RRsjTujnWZbMkUhANdKUCpBttLnsFTm23
QfiefGapJW+aXytmzbgd8lILXsrV0+s3Pt6lh/clo32+5eBcV6Tu/S3BsKjb
fI3DAejM3QBU2fSxCJbaVX6VpZNjJ2OYCARNrNg3ezT/obayOr4lRD135FBG
zFFSe5QgfJHoLe8iMAEwQH6P+tinqKAGH/W1C7pyTDRbD0kzf4Ge3bu6s6iE
dQ+yzfcfZePUpMvtMKQm1ZW5eUIslcRU8PFRLSVgRQfghuVTgmlYxtG+DbT9
gKh8lnC2fRkj+0RuwxR9PATeXbQQ0A9Xzt97QV4rCd5ybfUUeB+t0ITYMt+R
/jsmraww9Y9ufKHDq0RsgseK5ANcEGYtud2kYMI5D3XpUO1+ga2jwtcBIL4s
PScspqLrC9T4Uevr+yGUQa7xfcPN8/NH2wOU+ojSsnzcYziGFYpszBsX3uZ6
dW07RCtrbGi2HcHe+9l19iqDX39qMLF47psT26IF/2tLYBDHdEnPsKb9xKY+
QTZyimKJRNKU5Eq/AEP6Z23v126GXsDiUf9uyoWjV8NIjsbfCpa6HnFnBJZI
bzIlJLHbCnIoUFjrA4mM6MTN9sZtzk0yvSBasm9V9cfU0bSQCpF3qdFK42sS
WxiHySpohxXzMOoAeCi54Qi/oNLpqCjz5wz0noql/UCEOUq9HxfmSsp/gA56
jldHUcsWuTQeI2Cym9zUEXpbbuu9JkGVAbWAYKAMgdokiyP9LzlTg+KKm5do
B2JR3MjbQo3+b+Yh/xWgsgjkSJhkoh3o+SYH9opV6dtZROsWKdN1ZYwIOY8L
DhX1to2fErKN9mPb1x+ueVytu8bUnRmUO9/on7CnyDjDxAbInwMpHrPvqOwQ
Ia7tU60gUMIYBOw2b4nUjdg76i/ssF5hI1AG0hNd8gd/WE81JE9IwDCv002f
uDG3tn8ku+Tbf+C5B/updBpgHHOViGyT6fXOEamc3QTnFRbbz7EfCYmApxzP
uytSVAVKIZBmQ5bzZdeGFHK/NnVlPQ25FL8HRdGrVK4Y34DHRzVzcv0KpG8g
le3TqhzdlsOfoHkkwfqrYtFR8cPeFkfps9Q4dlLm8T7vAAWLQiAEdyv2BYrP
za07EMK+FVYJ0QrKlF28BdENHr+5LsMMfc9xjgt5tuF7K+7CgHvg9KacOuwg
zz9MeDuCeOFqFi7zJRuV/LQshWdBgOtri8wMIf39TU1uA5U02LmyNNlVGJid
wnaJizI/FfHx7f+rVW5+Or3Ammi40nmRtjgqOylC+jCaDVSjQoXWQ+C/cCC5
t0lKZSfRxJKWZ0+ZwznLPNl23vlmHSQIS1JcxJpW0PJ6hq/FHoo7ypmS07O/
LdpL8yl3eLq6ikbQGr5Apg+FRsZGT1W44m66iR6mvSdbMciJDR0Fjjyc1IDM
E3VXub20WfK+YOxf+2QDJU4BMsO4p538DKzUKZEmLnbVqdi7mG3OjwJsJ/Xn
tHNpykxTO7v87X1qRSYzYIItoLc1dXlP3h72M/dbBHsO0MIcCKemY/llb7o6
CyDRsVVtWX1anT0+pnQT9Abs1YIFT3Kknkk8Qs9UXcwcPLO9R1bj1/B1WvhZ
7J4M0r9OPhuVgUvN9CYOSj7OzG/B2/x/NAnsvdSf9XDW9eixwkqlJlW3R1Bo
NlS8xCB+l7aHWijj9uNGR7nzf8yKeDbvFmICykvdTOW0l1Npg9hxr0SXFFV1
bVssemkJXr7obhJOFvlNgGeB1pytTRi3oik/wU0bkeaI+kZD6w88RJ5rtZmB
uVmTPaumAWtTcd8+3YBOQOBq6KMdiqcj9ZLhl11phwxPysOFi0bNZspmyYE6
SfW7YXpbskAiQtFxRHqew3q7pP/VDbE/HBL5mzT7eEAb0qQd39ZVBLyUbPm7
CUvmMzuTaySrB9ci5AdJb1JOOmU+ERUTPOemaDOwnt2c8O8pHLKij76ZF6Db
aimyInDia3ECdHFNm5pwT0OAHB1b6WFnWksuA3AFyOLSHYQK6ZP7NWXPLCGJ
jCj6edj2Cqp/QIK+c+2lKAMXr1SjPh81NHpUndwxDJoGijh+sRdC6xqc8gc6
he9E5g+YGkPin15MOWMVOu8pewt+eUr+bXrctugFdgfUfH2K5iiHQV1clT39
BNXuxH/Sxa4bTnPEs0F43oIqTuEINesPlbU4mnLvlhJlIE9dYtWCE5rEeZ4I
dGFDGrwNTt5ANUynWIAGh2ZmCnvs2zGzZifLnLuqSnp7Qm6HwJ81f7Cb16xq
ogiRKBtwu3jGkX9GE2EYxol3bDC0brdJrN/bDlQHdFgQU894NNNw8qNpWksl
Cs+CPtLDfyLJsRDhvmjDIED5vr+zDxRPulm9NpOl3itT0ko0NcFbXF+mEGGs
2owahg9Lpv82OTH9tB4nIkGh/y4TEVLwoIGLH/1Cxbyl8zharln9TNs1cNYS
PS2ZuvQ+uGLaweHld5KJUXaTm/kbHKxwbslcY6dtfXS2xKZ+dD9P/2FUDKyt
Pbll3+m1lBT58kV5hzW901xJ99mu4JbpwuerwWfyrflMJzHVoFAjwgdmUF3o
hBhtk8vDHToUEBHN0uprXe4ftXtX0j3eLA8H8/SpuOva8pZnGjy8DeGWbnts
3Rw7uxM5VbXwjt+slMGEzH/COZtXRDvC++yxeqTAemQED7IXJvWa+WSCWrum
i0W/MvhFFRvyE3C3PeXFG5WH+JcSMaWYZkn0Ell/LKxag9+DNopSF8MkiJ6j
OuegulT2WfFJI0hse7pzkVtlm/IswpCdF0caoSJ9IeVScn5sXfsoT7YG69aV
9ltJvI+XtO3EfGSdvtwrhX1OTrfA+Dna48WNw20Vb5rsphLB6XjJQ6CuV15w
F3Sikpio46I6DbGGXCbWAxOVO1FC9bDtX1MPKaY446r/VBWDyeNDsTdvzIhZ
Z48neXtWUawD+1Ij94T1UScuaryXY/uEPp1i/Oh9f/2svw1FweYmQCbohNUW
ZEN2mE/CpXTQ2RKrNSLzzYHltI2yTKOVpeVPOTVEAeH+9NBkQlXrGZeSbgS7
+BPTpd+fOky8YnClTcYn1mwD2Ow/BgB12vZrvaS3tA5VVMCaGfcHDrzdPvzU
JREPl/+g0p6vW151QV3KZOuFlfs6YK2Q/L/zPBlOKfPpphkeRWsThWE+p8HH
pjzbHfxwZc/RTZFhAmyrJS2pB+3iTFnM6iXN4asvaEq1QhDTrNe9T9FqLhgO
K1Z/cLKc8ZjQSnEECxdhFw3W5/1tNysaotb4vwg/tLp/j0QME6yOTTMyqk2w
RXJoE2zAzeI2I98RJXPWQO/QnTALkMH0qQUB78xnaqEPyAMXAiAOyGkr5BaZ
xqtc2pNt6aM8oHVye8TBT722w4WXe/CBnN9UJXlxr3RE8Is0Ucsc2mxJKhCL
NsXjHHMSGNMvZSa9v/3hx3oIsG9QDziYHuzH1R44wdQq80vK+LGx0eqQHwBy
JM4wYDnir38bCRh+ydvY366jjFrSwq4IWEknNo0M44XorHrBK4MgWsA96k3h
5wVUp1sxaOJKVxOeU5iOgHLsZNonsILqlOIZBqSyVqtx0OJYk31UnObB5Bv1
r/uc1rJS8J7RqC7JXb/VcWbOVxgF468P+kgj+5Rr3BZUzU9oERT/XNTqv8dG
S/MqJGOUDoIzvnbAixw2hPp64FM2SjRXDEvZU3PMcU6F6gH99mS4B1k2lda5
zXquG/cXKAju5oQU09lFFnXUqqj/KeJq4vQUBxJz51dwFwJlUoMXvSRh5GTh
6hZToA1gP96mfFm9qk46Lhj8sLDuOaICE8ELdc3PuyY9H4ibSqbwlBPDUIgv
rOjx33pSeGK9RhySdpue1gAZvbV1SuDBsTXVye3awzyLAaoXBNMkm/J0mAaX
z9UTfmPbjweJD6mhoa0ol2zTQyCwXGjlKYUHKBRw3Tzd5a2bsiNTSQ4UFBky
uFNL+hK9baUUav8BxCvxaiHePqNg7umba4LELYmaUP1Kp+DJ9axHdEfv7h/h
93SJBLWF9iZu5IyDY1GshcKWWrZuavGZJFcTcj20JPwx5FmdhOlwBBAmUEf5
QOvv/NFh3OdCAs2Arr6gpXzhRbu4LRqzsw0nJhb6KtTh0Su5JV6sYeLZqMpb
KNgrbxB3ilGYdaADfHQXvfdlSzCcIHJmCoyNp6KDziVvAf2Y4miKKhXs9c1B
IDXrzAcrY9/Sq3vPaFKdUc0bp7RKNkz9zqKuXexoO2uvWeCj44V+ZUupW3iZ
AK4KwoSHJMub7HZjhZhoTrGOr6K7s5sbzULNzvsRwqHqMWrrKQlaSFQ4CdK+
oT5DxHyllzPcDPzfIHlJ7py8pmhZdCz65MEkTmiEa2SCLCQ9RVVYXePfzzBX
hdkTvRkoZtTrzSAsw1h+tPah3Z9DJXDyfca32k4tK6aEu7LkanUXkwPLIeqe
ehCV1Ab00uhyMJZBkB6qJzlOGLk09uvbuXiJ80cEVbxTJIyWvnflFLUTRz2U
0uYWnDSVa7l5Ac5g9yMzOtFK0T5Ue+lfk5z79D8cJvhk/l7xp7p5pe4VJffq
zivnukay2fICkt9N48hym9vkks2gEDqOHrKBKS8RvZsVGintlhr6IcW7hP4v
1fpMiUMBKLBptr8304ek6TtZOW4guVTtb+KrujUxmIvCrAsOHRaABlTMaoGf
3+/RvMFQrLwdP4JecZ/I9DUGhN3+F5yY73oXJscoQOO5XWQ8eCeha85wVDxf
mfxQ1wGaMo+xWDKfKz3ygFgGNI6JHBTwPcNGYkWMRlvB3sau4RnIS/f3g24R
TBvz7wRNDeKIX/aMhjp8BV1tsoAFr4El/rGiT7Db/2fzSVDb5JC4QfdN1J2Z
CvcEnNB7EM8LMbuXDywvXqjzqM4Nm/6Ncaye7R/6vPRZQAKUWQqvBfdpzZie
dI+Cp2vToo0iJqL4vfQckgoMINYuk/luylF62ThefgXfMpRh6ZlYktJUjaZ4
t7HY6pNod6NMUDBQJ9QNB50pch99kU+o9xtxcT+tzTGVf5Ptg/6qbq9UedyK
RL0w5ymzF6HMK919S6aPPE0qIqzZgt8zOaZezZX/6gBrAhPbowK/3ADD9Jsk
9aM5vGqu+aOLS6cshoUv36/J9faAZH3taEgxFpkcXja+AbXNhD37gGaLCZ6v
nl+OA7NjVvOysLMmSv17qPMiJPGNW3ijZqk15CiE5oEwDro9JMqGtJy4AkJZ
FtfjoLWZC3X+dQoAbOmg2XCxOTOVEWVjpbmUyT0s9CckDs1Nj+kn0ulN5hrv
+sbbrKMrwUJTtHZ2tmnTSPtHGcIaD4BbZze4dg2W4OsUquvzdigUHuWy89VV
UYizs7dMl6ZfkaySRuIUMCxxhujw9UynruJQBOD7LHhjvI26S2gWsLJODl7z
bAXG09i67HinvU1fFzC/G/bYWWNvmuH8FmzyQKUKJutriTLUjOHDTF5LtHEH
bYdc7F/beEFaQu0xNkF9NeyjazTbpOFG0yxlDmNnpO3n3GflocItf2lKkpHQ
coJ9WlhVu+O98H/as6ZDiOq5sGOGFBmHSQuTRZLuqhJnmiAweDAdy8yn9Kaj
ZDeqciyGBzNrMl5xtQs++2wBxOKIzDo5o1sy4nD7FTsiTc+1NKXR4Ad47NQ2
3cf70kOSnKrJXiJu93W2dxL00mhAyqyPdI7kI0+BLY40+n9Me+SSeNRULhxN
s3CjMwx37oZ9tmsherPLoCp+wcM/NiQwjogWZBpENTjf/bnRDM4VOIvNhteC
7KzmgGIbgc9NfuCuiDhNwVxo4ZVubVkFNltozLRB9LDjGyN9KM+iJDU0PUzF
4kfYOBDUWHaNwOmK0q1nFbQStYTqKmZNUlrP4iqd7GSQQJnl/xS3hkLepdOW
THCp7qL74oJP7LDtDCYvuhGCIJB3am47UX2EXzn6gIDM3nWSCbrzfASEvLQ/
hyWRc5gq4g6AdPq7pz4lev4tVWx26hKrqkFhet19Fi1YSK+mSV1BxFN5jiRG
S4HQRMxx/WK/DS/ZAjDTOxHuvDShdm0wv08P9eVUAcvSQmsjr/2Z9W/oUX5y
cy5q3GCH07jDDfZBmC567I7H+8a93sv2PuBcUqz+ECUwH82PRzHg2+lcdqKi
NFSMVN0s13PxPD1yh47KH9zkbjnh8PvGNgHafnC6rfhC00XIG6ZNZD/9GufR
Fzii4DqE8/mSveNUugFqTI5cj3waoDpYQ/78bNXtWGYJdo3RdXnoBn+vbGUb
fn5+KkSoqPpKsKDF53iCCYtm+ro1FfVASAg9OZcvG9JRPSfNMn0huXg+oNbu
pDI7rdOjRoq0pB9qtJn24ofpLoeu/smZErVUqslUCKdLsz47aq6CRoWyaSiC
I8Y3S+ypGhfIO2ApsY/FbbKqzulYwDjiOGZXhZebIFvPoMVRE3n38liunQ4u
L5oUPahwPpL4IYiUjmRhEXBlgnCliPupEhuhF9cyZPdszO6cQh0HDlnovQOP
feVnYGJKBQpSZOHjjWb6dumH7HQUuU2ZXXyFGFpc92uelAbKezlDHp2Vz4wI
3RY9j1PlQpxOCorkGp0GcRbxfqsWt2BDrSSnsiH93OQYk4SJC5FFD33jNIju
dj/8hiCUdWnu86LX2THhhNVDezwuhLuTOq+p/VzntbajQKqSIxseKxsEaOrZ
V+opGhdwJuiN58yatlacMC5Yb+l/p0qD4Iuvvc2VZtLFt2R0Ssw9GhdQ4hyi
Q41xSwRe5Hp+hcdTv1cMHJRRh3xjEd8W2pmlV/w9iw5jcaCEwv/fELetj4+p
kdR6Kze70uAHzAUxqvvRPAW65tMJagWN8arHofaPuu9+w3rzbVEdDuEShpyC
SAD2hpADYJ7rQErVKM6GzuTJn5BvJhYzACu1WUqSnNbGQxCptKX9JVy7ET5v
rGm6DCVMDFCUp6ONXRllkncNYz1zZrLIoxg3Ns+iw0+lujWqAAd75oQhTTji
4vk8os3wng8qY2sLZf+oAG6YHVGPkCxu8gQmdP9hsT41zfVnBLLdQ1ZcMdG8
4vKMOkLY6TodK1+MltDLqjWYiEIBaoSy4oaj87B4uHML4OI90nHrrz2TdU5N
UcXfWb3nJa/0jIY7pPs7tjRYVZRduyDbwnl0Y35v2ItscsBqUJ9y3zjNrXT4
oPgGuH9RB6CUqGEGCRi2bozPrEkXA5tcwLuefmRhS7Kggq/IPjwncMA6w6wY
mHtcPfj9sr7pjsR9c/6yqdvnr4STXl1wqJ9eLMpwBhmmVE2rH7XpmTpj4QF+
x3Jvu1tbFQBJaGA9W0aV5QzI87DEm270K8ZkOGeuG3t5kcm5JfvcZm0hbuGe
bSOrCCEGKVzKBcpenlalTg+ia2gPx3F+jpCP9MJviLN2fit8SHpvECExcOMt
nB9Pjl17ABOJk31/gUX83AllP7Mvwa/i7bxKq23IpNp4xrFEin9FdMeH4HDk
xK6z7dJdzvmR4THeHaaURoGkzAdJml40Gj9s6ipKjdzg+ncJJjiVEmXSSsnk
4alYxy6tkY7aBjp6KPbVW4hghif6NPhEvAXmfc8LalG2fqL4JyWnTpRIImyg
LlGX4dT9FMtKgUU3GsVt5mwiPNAQdFBx8E4Z0XrziRGjUoiGCH4dOBBfd9/K
R3XtB8Aphk6aVq5O4y4fFCp+aG5skf7Gx3NzYLVsSs2XtRf/x8Iw9tdwJoAX
H3G4AjIqhe5oTngbJXTYOF5+Z0zbgYxWQQCv36+k0plRETkBWH9xwXZ485B3
0xGlNQ+NYCkAoe1qlC9RvRglhnzUVPhCNLxNvCm5LBbgPTa+37w7kQCQdIBd
4BXlafg4TQwKce5tDhZuKWqvJ0rBppnaE4U3Pu8j/NuBMZAQJH9T4VmUwoNx
3xEASAWKd671IwJt8kpqi2GmkXboJTCwoKFCUQ7KgQwwrlLIXuJAcYEm6a0n
7Wp2Z0SsdbTICsAFgPtrDwYAozIMxRfDqRGu3cpp3V5A5f6IkXMUMOTfVJTJ
bCVO8PsCPuXeIZ6Su4Y8EtbWYi3NKz9vc7he9RuM+3DDpJuuIsj6ieVWi4pl
UqFPahrQjBJrNmoj96M4zNNIX2XvSXyhmW5lDrLp3+Jt85LnhhT2TQJFUfyK
cUk3rOUqZD4c5EYDC4zw36adFooEg9p1DizcC4Tnbo4T9pYldxeMV5CMaHAK
ea3BWey/yVgopFc5+uuH5ChrgP5opw4kWPR4xD0Nj5UPZY/ZQCtUmiLbAieW
H4FjiGbmp0JFg6FIl5Z/rse5FK8tK5sv4De913ZMlpHv0ms4VKQMXcTBY4+O
+ac7k9jROugazVq35AKWL0G3NxPhFlEO5H+m9vAmxrJBqtfcPcEuCI/Ddoay
34OVzZVTtyKoHc3shYP0hIW7NT+XmBCVRT+R0YUe8uFxZXL6LyWu2lKT07oM
9kdJ1nvqdjUGSM6PJQaFTwKrSRujchG1dnS+UOqoTjkFoJoCLEgXy0Pu4/FP
1ERjHhzzMWu/pSBb09TyW4fJyCDg3nUzyc20ywVFmezb9GR9Iv5OvstQeQK4
XpVBoUxaCVy+XH/Z9svhY8aBzEh/Pnj1NztTd8TMgIS7FOvrNInnOClSVKcB
Cfn9Eb3dXTYDqJlmtDq8PTyEee4hi9R6SyVtqyaI7c8PF7j1sYtiNLsb18Co
p+iKLBsbW9jk2wTZOj5fod3T9iB3ut9iSo17Jsn9+5i7eyIbDsc3/8Sg7eV+
l3bxyeWPRUrrgZvduKsN1oTxaMebA4fLkt6VrrrirsHR35iUBE0NHB4isEM2
fPUgjISAkO1OYWZ3SEYVcSMh0vV3UVpy/fNAczMRLmCy/TtplV6ITmKKoSI9
9S04cMRFZlHTl2BhcA+R2C7jZzoLVA0hdwWO9dXox8Cu5YPpxGt0qLTJw36m
MPjwwYqcBD6DWKNRevSZ8nVgHVoft4wxYaIzXbUZn4xFHvekn+vbi5lw4g/l
+JucLQdbin4nI0BjftaOoitXkIeMRPt1co7Xi+NXTGUtyAZ38+hxfRIuj48E
eTOsIll0WS62nDgIz0dS1U165Pt1mURwev0OpOmDuX+zJUGA68GbdjPNCNmD
U8xzuZ3Ub0vy3AQWHO5A7b9VtiDuuZFyHwC+nnqwbxG4Do691ANG2eVErENQ
/FgrTjNV1ukHRBfCH4ZOMBWbVMmiZKVzBfrZ1BS/QsaZ2KvsYbs3dfHoyMLS
lrUCR1oNnle8g0auj9AB9yttB3zFKDdLZ+khsGEWwdZW/FRmCp6qF+T37R96
DQE1CFQmsp3g66KyyT8VpJyYq9DRJKbYYfva6xpCHEJhQLm96NKKvXRudWnV
l9PQVgBpZE7zlH6IIAQr43x+ZOIOunyZ5OpxnGVe0gjwM2x9SC2LUlbiixsa
5HCpjO/z/aP6JalQHbGxUNq/nxmjd4ma7uccFfno6XvSvG/GMG8Jf4shk5TO
OztoQJH46a5XEro1agPj19pVkuWhiSHl339Ly4yfbnmCieA1ZZ0hX4X1s9Mu
a1QLbNYWjo6Zxdc/yLu0sydMD0s9RE5BaO3i4pJmrpsERCcCnZ6YGZnkiTKc
OPAMbiQY6gKTxDf4fQT75gAW7cXiyT6us9Eg9qudRds4ND5KF5Xc/2XPRFJl
97wkFdyZB54Qu5ARneKW7GHXbXNlqzFzpnU1ohr+O6QIw4eCRbDkPzm9nfOf
KWIq2YJWJ9Fqzkt2KXTlaHANIcJ9pYLjzOrE5qjc54WfKbYIkORvAQTt2HdO
uUrIm1x9T3h5PRsu3zJJj9ekEzwwtaIWwAq+zQhT8ZhKQUhJhkfeRcVS9+ln
GPgDBdILzkOWCXmGVCBnbdE9lzGXZftW/3YBpI3tEGO9EsgojApwA+NBDhHE
Ot2n3DOCfrFR9Tq11OFkIe3235FixOl4CS/y2Xq6vS22IXNJM2HyXusUwEc+
B0LA0yJQvWuPlajkQ11NOTTNw0DZJtcEXBSBIof2gK0x4cr6NygrICA1rZdM
Acl17Vv6nx05ww6ppZM6y1zIhCGZngAgjEVPK8nBsOIl9Z6LGmh3oSh1sD7H
Kswbjftzy57fuNqPOdPiej+0Dc94Z/mmJPLY+5LNZnhQNNI6POUhV2wJa2yx
kovpmQ9iVNnlzALtZOPzEvFOXGAlVbqeWZqOYyR7hA+YQafZp0/BtdWTn819
c+6Z1RPo668l03NP6lhCKieXhNzyLJB3bXfNG9iDyDvISuTXXNyPWqix5Nr9
Q27becLFjZEt4VQKGqeMKw+WvuU7fYLEu6/y8TjczyZ5K8iXR+FtiJG3F+MD
ueVyiSXU+1DEeTkszkTz637YIlb+bPqwnjFoGbM4RrGec6LLf/HTnwYEQGVn
YgWEjGzNQueTrVigf2VTL5/1ras9n8Que6pHj7kF0h013ulfgvhLIIKSub75
8tc3YswSo4GhtGCuYiUtMkCykSZgTfnDzMXRxUsMtKK8NvPMgSpk2Yt9Cie8
Z44LarASmfrZ85gXezJFPYrW3ZOT0uIkavcTGvClbWNUPjHOX4KXlUK9k9Xh
2BS4Js5aqxmOXGCzA/LVRxOPWzy0EEZEu+rFSAKFJkUJGnw/40Dz1/cJDCZN
d4gz2z5ecA6MyZu2mQr5JwXOdD2qIqWTM6K+JkRiltw03wxbYiPBfwLV0H6n
bVP3UtU/+egQuniQpVq9oc+qFsG+C2H2ZWnVeQtiMVGSMiS3bFFqrxKWhaCQ
kK7zXrR/5NKiEt+gUikNjycE0/tODGm6GEKLBCKYsMVYJ1h7UcCkSaTVoOQp
0KWGVNoyYwhUe/FYljc3Hpv7VKCcAjs6HH9aFk5kAlwb25V8QqS6B2gw46TS
TrPcIPdzKdWJNWbJQinPVaTsPpB7LtdKqhSbHqdrP4k0GgiCqKyJqWRb6cOf
qketQS/pJP+2rfb+KEzzXKUdRgfjVLN2/yXI1sHWrVbqciZiuy18OvIBb0HJ
L9edJ+TWmuR1leI5bnjz8AopDblsbOExWcI0MwvisxOiJX7OQEKYMDnkHlOl
K7uYZcgQ5yQ0lu3965vqJaD5PxkTOEWfoxWppbPrRu0HxZGlAYXJyBkPnMRO
ft5RQuPoXd0w8xZNpf97MKZcnJeoV5/mCz3AiSTSSU+GF8exDOUPsoSz4wDD
q3+Q/cNhMTjFH+OMsS578NTN2f8QEK5uSuq5w5sdYtt2UE0bpBjuBIPkx3I6
B0O8ufLrnVHxGVRiSL43zV3CXMIPYyLBELch5yX3kq162M105DH0m3q4agCQ
PsvmIwEVHQxajkI653vs/bIeV62nRJ18suCC6BsJouYM4J/w1DDgMEbV6p7i
sGs2j8+mP42FKqQRMrVqQD+Pudnfwk2Ycjiy4ZYxNKp5BZ5bjf09NzDI5V/O
1yzFLnD1bSrZPk/ezCxwHCOrO6x7G7fW23L6/8/tJFxmabIrwAPEOUQpnNdl
HhuyIxAsHwv1LsCQgKgb39n4I22PysbDyX12EDHxcqVpokL9yd9QOXxkVk0t
kqBMC6+Cnzqu/FHo92fML53wk4JtvygAmrg/9fVhuWAyYts5UORN6o3KwLl3
0+TeAcGOp/5em+Lr5WhbTNJK1VYTo/+Lty5lrQUk6j7WK3iLPyqPPXhO4x69
bKD4Wi7yJ/SEDJ2uygTw+NDpiRxV4Ae050UfATp35qExHWgO38Y19YeOcgC5
jQida0TptuQ2dLSycLG22tXMMGF3N+f8n5aWT1Nx9zBxENTPLczlk3nFn7nc
2zbI0gONXhhzBYiO5bYjan82a5vG4q9AX/WpMGIejnjZM2nEAuu5KuTKf54X
yalQ7jqkbc1BpUljk3vOwfxm9AN4UAKzYnBQWAWT15LqkNzPsyOO2TUtBS0x
xFDdyUmb1mEemMs2LQRxlQo3kZq9uT4WKuR3i8bV2hJwrOZYTZSQAQeblYUf
XCgksJO9L+SKmPrXYdCYicv0oQHAzKQ0gMWj55vTLQIa40IF6pgi+PtRQGEh
jjX54kf3O19WSlwuICxXEtSf18kUEMV5n+cjxwutMmVGn6ki7Fp86s249YOr
DkIvkvj6JPTmMiM4NimwvhfHTgP4VtTk+QxCXYB37fwwb0FDn+i62EdQyoLo
B9sqjUEyEK2tZnA1zoB/Vwbj6RMeHNV9GcQJ0IFZYuN25gKiw5c51MvX2UGC
/nh5YDi29vO9DkH2iTJ0dKFRVpMJYV7JcnnQo5F3CDof+25e/ueBmq6uk8NQ
xTVjnwbkG0lSq5QEel6OKOBq+fa9rPqkXdfaW4kQxsZPe3QX4SIFmwvixJuV
O0qdiFL/kSMS1kjHRAr5ITe0m1J85Ux/rxIX3dbHdHeXVr5TsLI4NLYibIcy
wi9P4drEGGslfxpB96iEKgQqQqmc1C+mmz/NS0aDWsV/XBOPJ61P7zveDNjq
i5gUmilb+0ObUNiHGXEdgHlYWlt6E3aXG7Llktnd1eRtuildYUlLFlA4vj3O
ncTNqF6QNzTtF1WqVkGAnG9pSZkOdw8tYsWg9NiXRDrxP9Pn/pYbH+H0YELp
3qrD1zbzBSlgSDAjEaV6t3+RQK5N6bLwbNoxG0TnxFOyNHPzGyUCPt0bMxna
oN8RbEQp6LlK7tpPIWU1AS/Z6kVEvF76iFin240XQ+m8M9k8rnmc/pkafJdj
Uxg9y6fpXlxOTR+DDPQs9gqXqI9BXRKHXgtwDEEakBQysJQUREcshFYhzJFj
chsG3zgsP48w2XkEjMMnS+YQkhWGAUZZeouveXltB9HEPF7+CRUZ+YGPmgLt
RNfbCu67zclzPERK63exRTERmQTeFT/WjdT+D/XQLl48xRS61nWkyLZp4s64
8FBmRN/V9FFTbmAZqFy0UyJs/5eBUfoARCB9kT9uLZE2/sYAO/wgKYsllQ+r
NKCxIxhXeP8p3QfSop3oC/5t6iJgW7dlZwWcvvy7tWILSRMNPbJfCNeqcl82
y22rdO3pZzkVEL8VeSp824NfC0tQJkH0TdT/XVvrI5WvYQ7zmgHi3sqlglaM
vysbX4pPVDNzDIb902h0xkbvMavZ4ALjDl0kirV8lctM7HjOtBX9yTT3cuJ6
mosL+eqCkB2eus/W1EDQfjkyvfgRNxnHA1gfdERjHDFvMVt/+7PWLLG279iN
6PbkzfsWf+XzJVj5aOvVVkYFE6talHBG92mY13l3RKiwyupDMFhEm6b47z7H
Hq5Z4IvZl7sRGwMSkaXQCssVF0gC4jVeFJoj4MsOW9GUZGvDu+XudipwmNJj
Vjn+0qbPQjPHyd/B3Izxcm63hSrTIgbGdpYfe3f27yMy6ck6tMVLkr3VD6p1
vjsIq9JEzpbGH/GEPN1Pps04ySsnBf8CQtrFugNVPnmdZ+5BsPD0t9qao79i
MK9HyK8zY7iAkyIriLdEO6zZdbtic35GO2mJJ9V0LTq8anrFRusrQ0IhNT8x
LMmCEm622n1+caA63Q695f6/2Q9V+xZSqk50rhj9zQEepymteKpQG0fcfbJ3
OwcBo4E3oyruN8tCWYrFGcg78J91S7ytCjHgFN5q7Gbudrub7uF1pqw4sRx6
jg8xqUmEX7h/uIw4A8b38jWRKKY3tgQgEgv3ZFiblhSfsNe72weVZCw2R24q
B7UjUq+s3perTBWI9EusLQdKUSgriHSSvFI9ZfqV7l1AnqiCnUrYHErfV+9J
Sl7EyNSyzF3gjveYUpdMzfmLDLW2iMcGFDdFCZucyxOYb16oxr7YcqmT2zlZ
v9Q4WI+dqhxdh7uqNlew4fHW4nsV2KYisOfWospSkGgDKsCIA9LoSFhLUGao
PSS1P9GjFRL61XVPuHgTqx2o9WggRhozTFCBu+YQb3U/tfcrnt5XWvoMkGPk
a/Tq8CZDLKS5wm4HSegRTARXSSvyWtg0kAu/ykK6+nIB/Vv6yHPOopDFWwbN
RkQPFo7mW8nOdbt7Nsa1wNdpmsT2aZLVCBSwKFaDybtYXj2sl7J29+nvmV7g
rGwQaF3mnxCx/LEFinnXBKhOCo1HxmLoWXbh49gSj7mUA49hnyNVwIr2LTWi
ddY2ePfkNO8pT3fMCnNYlvSPXmkUFeoYP6eThGUDG0buQIazim/cxy4GMeTA
+Il62QsJarUzFVBqct1rFRMGniLfRXCPm9OGEcDDwBmkMKhs/N5svvj9f3TV
bp2UxduCZczTnsJp5QpzUmoFi7gJbY8GIOFmzSX2gTeUNvD2MwME9xVcXSBm
UVax95PyFcUV/QS7A87kCdp9j96xg+CMTSSf5TGSYJfkbPfilUz+s67u+JuP
XMKijeF2SLg8PWwG1yANJDamiQKy+L8+uoXcdtMh8HcgfVvvacIPt4P+6CsN
jOzfph9/FgqhlZKZfgrorC/chMDm61hsfokSSqjGnmwSTIwwQDfTPbbw/J/J
lGFnXPX4lmrcmcwNQk+uDlZXCXOQplVRxt3lYLquBMJfjvkyA9UDF7whM7yE
xrbIFNH/V9UlHWr8n9qHuRrWFF9niDpZsDUrmz2tg3kjV7K4SKp4LWKG6W6z
z6bxrNxuZKV1lx42mHHAiqNVLA1OXqpOE/D20e3tw+N0C4K/qWXIXdCfblj6
/6OZ2GoH+jJ4YpWbI5UD6PjpW9wLNkndRJ1U5Mw9yFbHmTWIsK1KDPNp6i3l
tbXiIOlQEFRy1+NRpfQzK0JVpTONpBosdNNUuLynNz+WZx47Q0AI02gv3kJJ
dEKR9NpngR81U3O8BN932GsUKue7XtsGC5W6AcuBSpvvoW0fQyHS6flxB8i/
050filwpkUEmx/qw/yGAanQbBf2MGF1csLSeBuG5I7rGP00DplxtoAufe1te
Ezsd/fJ2X+4ghQtY3w5tHvU0fm8a7Vm3WSwq1kYRity6lPM+BVTRurgaGhQQ
r2a8PEhw2sE2Dw2gXf+uSjiVQCmOVBGjZaDDrfOAGnaO5b96LHZXRmYet8sN
t6Le8jR4MS1XNZvOYEpqj12A0oBZ/2M2TpvdMBD8a3pydiJvCQXFa6shCNXb
sbUqP0VEaBYQ1+xF43dloSo+diXTORjZZtGdW6ZEQiMRD57/kexuLw33X/Rn
yXcrIABfaojBjpjrKgjYlBlt9rxZt/JQ1bK1gO2NaKCj5FIo7NI4eiVAOau4
j2g/SHfctK9isqB8xvvcArkAPo8f0XVr6IVVxFgPB6iqxOaBZT3XSz5AQ3mW
XZHTTevGDwmfOI3iWVD2Xw5FfqJWHhcrXiyw6zUSQ7Nv6edkpapptceoJh9n
nT6r2JOCL/9VGMxZhMWovJvJO4okzsktyQEwtiRsquPVsN3l0N38cm7Sv4PR
ADBhjkX/WWvFn9sin0Ruu6cTs0JnXDPKjACx84L7b77g/vwXBH7aYKH8vxRg
pB1ZsdFhu84v1QAHUDwnGwxrk5XbkJ65DyktsV1zJBPUHD2kyqei3AqjiRkz
7QU3+fIiRrVZ7/PLhFRmnGt9DkguY4WZdTQMI4pBikFWmDNSiPbL35bihtW7
cbxXrBrcDByyCWayEhR0M6hkq8Pw3ROkFjIq6P9D/KLipGeGhxPsW19UHIQX
YvTNh67zo3TS6B1TvPF+A6fNLpMmz8g1jPFBl2VlTugM3uIbf4shRJccaZy7
qmJG5SFNKgZelEeXaAaAPXZqOd/kGjmTS5w+SOsHJUkv0G6FKOzVaqvmbb0j
aU1CVFJJyWntjavYf7M+4ZAqSyVa+SJ5e3qaYO4ZgTXgzBg3C5qi/KqCCd73
U1SQf/UkxtP+5AysaNEBI4XkgZWnscbyc5JZsaB5sACnQEGW97xgm4ttoBUe
Gp6IA8an3Az6AWpDGH965KcGZ0HSHwlvdEC+MYJEjCgXqXJkdZOsOcjZoGzB
dgguO4d5g3FiR8cRLxv70Pp3boJZePYRNjYOMFlcpvBUeb5emkDp4t8Vw2pi
hc0/E2JNEkN2ZZ/Xvqevq6EqTgVCZAwh8xKzzQ48HieWLV9gVNSrSaAgfXCR
yD7xpSOr6HiDz3hPWIh3b6+4sZNbaEU9pqPFWW4cw4/bm4LWMyUrufa6nPIa
GqKHPg+ARmA0EC2lA2vOJAWfghIoguGK8zntOFfM3iK5YpCW+lucq9w+tN93
uPPXdGuNS29T7F5mAPxZMgx+gBBjIPnBnfIhnKcSKfOK35t19zug12yE8xun
McxrHmm3DSxs+LYM6GvUcXRMN45SCdpQ8ci/aCrthrRii77iVXKbgX9jpRAv
b0jSoHgPwXuOS+ABzlLzoVBJcoMjVCX7NBli1W6ytcyDbjzarAQF4Kho82QB
9/OixepETydLyJSShYyl91RXn/MJbAodWiiQy+dPHvRaC2cGbMyXjMH02By0
dB0XAUdBhcjWpBSVIYXm5uTSosiPxQh7lS+jVkZyRbmAoTz9YbcDt3Ljss5W
lc5uGdbbjjX6pdqy5oMHEm+UvKj8AkT3vORS4YLmVamyga7d4PM+m37kf7XM
PcorUQtPaFR736v8gQKHnAt3VMjFYjC07fLufJXPdQCe9BoAYa2QpewKpVLZ
cqX27CD9Rr0MkAdtcmNSbjjTWLfi2Z74H7Gts2kctbwvoDFARt8407p91Gir
fHrq/XTnJS3C0f821fx3ymd7R2Dci6PkGUrgZMvS9JYBEjlxiYZ41hf329c2
GYV+63zodLnpRiOCG/ayi8KJojjyG5/rKsxt4IyVvZz26rQ0gvEbJyeMtmYT
m6X3YdIaEEjF9/eb2wYRPBH8PKdFrZAIzcXOnm5IpcPl1R5gdH0hyoit0emx
W5Wj9hR8GBwnaUmyFd4KcxnV5WabjI2ITiF1mcSCHpKFXzeHFyEvleNKB5hg
SLosjX2NnFcpojKUemej64Csc5b+m1JsS8nmqYvYvOsXammHbDkp8GRpV3JY
lml/CBKwNf5BYxDJ1sXqsVHO2DRY+U91t2vZrZEWGS00ATYNTVzXklfVFVD0
QBeZLkof/dtMxO6oCM4QkAFZ9jAKHHRjGObAvIRE7cbWbQFfu/6VulCVKc+9
F37ZY4CtbxIeEvbuUoReomnTVOv5VdyHSks8nZ6dZGRp/aw1MlVb3xWlirKb
ZxkJCdbZKppU/AchVIgP8onAYQIPqVIx1ayMNsa/R5CZ7G1QwFTauiZ1ksQw
W7QYRz0+uplRQn7NSzCkng16g8TAZy4W7gruZ5cf1KPvrTsXZ+eOQ4xtVLTU
W63f76hNRSMjCgCY7apxSUsuiJ9OFliwxhvKwBs09XOCzmNIvGZ9c+ldKCje
VywmSau5DbABaITYckLjWjK6OT2qvA2+EuCCOmtReXFO7jh53C5T8PPzAyyS
Z9qqKbapJyAn/ngxEKVz6pLXOucV61a/OBwcbBLq7IN35bMECC1B9RPg8Un7
UNU8RaiQgdRtmNT4d43w1ol1GrlE74xAHirJW2mzJGnpOG10rvizMrkBF5Lw
65xhf64CDa6Cm+wJfTnuvNtSEcc4udXrxmAUOjS8QbtzGD9bb3q0+6xeijUH
dYGDDA2nsVSwmBvyMqW63PaS70HO99a4mnoLkZ0/7B8YMAKlAcBt9dEiJ+Fd
LgTISF+Rvg+gxtSL371z7Mf+J04Rcujw9LjsKqJXSi9d5Ax/0bMKo6mqHvPw
JmwbekJ6u194LetjCLyJYBbZ3filPsDc7XrqUy+O5VSesbsG5mdLF3H7HY/U
zWtaFEJJksnSm+AK1FDjprmPaXRyd0umSqpZbYuKmOt7F4m4o1HGZr9enzHh
1fxgQ3vfjKQTdLia7S2ohTdp1FaJNi78MnY8QAtZzmiktsYZyt5wUfQZAGvr
+N4x6xJI98RLRuFMD1P+59lSw0AclPga5Bp7hNsiKeZT1Vnm+YFFbfbbwgnG
hGv+AIzFzvV15B7NNOZIk9MFkq2E14auocRkEdOzGmTiqkoNqHXrAuvLqqpD
edR0GuyUU44aPgv4zanFKpxLRWFZjH83HUNcRWfDWZiAOVtsmJ8bFj3jzbdf
RvvivpjCCgO1rf1ltdN0KZ8+dznZbH6pNElg8EQLxjTb/rcU3Pt6ruLWHkzJ
AS7eGcE+fgLYdbrNlt5dxtstu+2bplF3DWjG/2Gzg5goKy+FDGiDYGTIQpJt
v7u6hR/YmWzrziWQ5EHzlyl4tW2CfnfYCPYOsCWn6BUlZ3mZp6YLBUojXm0B
1bMyqBq4jeHhRvdTS6oL6c+uZ2lOeYj7CtEsASwPnmq4XIz5ZOtKhji9PVnu
d4eCRojQAMdVDG5i7b/coKEIG3NJbUkikrd65vm8V4Ohi1qdqrzUHDoJ2PNZ
X8Dc8AH/JPYqc8Dxu/VeeKC+KopznlLMf9qt9lIr1z67r064hnKvavJ9+YEX
URw4XrnpM90mKPtEEpdElQqiKI9mhOMNhFNq33QLtjeECX1i2rGbKXbkU5cj
hvkugn3DJ0/YpMIXwrES4z7Ialbq2MizUk9O686cERSm9kxF0/q6lEW5xSIw
qr2+dW+f+ifQO1Ql0I4mNqdZpYbGCjxTjpdKlmzwUmp7zUl0WLQU/6RsxcK9
ZOw/HifR9sgnBpNps7Y9yNLFLJdVNmRe3QTWDwsDQlWk6S2Ih6+OzjWHcNS/
EL7hJPeCNVl9e5WTYKDvA08DSKdXRuKqUhesJ+iv+VAYbS+tJ6FSDQHcD7nl
W/LU4347tFC6FS51yfZ3jnNxyN1caJ4WKaN5uMWberfMQ+zxffIVC+nvn+w7
Wjn0+sbcqTNfnxprGOMXr4oPEFtyVKtukItSlQ6XxwANFtK+KsDH5irK1mPE
0aIs+5hjsGAXbNZ8m7RMMKNAaQ5jpTbgyPYZ2thc6SGuPNNQdqgYRb8v8RAz
oIa8ECOyzknbuC1M9Jz7zDCa4IhFqHn1IItcNtxR1g7uQcbWTjA+f+datVyt
kIGZ/1iX23oBJGm+b+QntzyQF5qg0gmFTqMqyrtCSlfGaCP//NmJBMR256uK
1km/Ee4xfBeWopXIPFbv5ZOI+MtNNOWA+H8QKOC3/StnP8GePCk6aESyM45d
jNl0ze/Vr4UHanMhCps8Rj20VtLxe61FUQ+/LlKm+y+W9pMvOxfAQKYgIF42
m/ddXSCZkjo+7fYPSPvtEiQA5VfcIvNfNDKaoVHpGco7qQEDU4NU7ljxq6W+
KvkZgOf0sET/MvX4O/zXVSmdzwXCNUBHNwIlJ66h4A3RMRLppPs6KcYcB6WA
6jA2zEM12SHP/fkj7JK6Q6mqyDuf3i6uYiju4dGkCzesDE9hsRVKYWl8vkng
kpLDsVyH5C6uD8R1K0J4vKH1wA8gd6ZXXCebywvm/8bLr4NnWwk/O1jLT5pO
UJuHwz0zFL2Bz+WhvxqmqqHB/dDeFPz73JGhPSRttjinZvSizQhGmG98+6Zj
t42W+4sGxPX9NlgXTZRy5PYR1B8PErR2H6J9EzgT9snRwaNjQHlf7UWIHuGM
acQAajmuqBCAtXyKFzV5LcBB7W69nBm5kpOLlN96DHJIgN11/8QxbJGG8czY
cwkfI11SYUD+qTb3YWysVSP9H/YBsS0S+FA3TrbPC1Y9cYqqQ4elbsuViZ0z
Wd6Ar5MAhEGk4sXlTHJISD7G5U1fGG3Amv9KF9DHV586JWZaRU49RKKrd3d7
s5uHD2kQIUG7cWx7LBzjIP1NqzEODh03N4pPGIlpLyMCou+rC0PvxiFFuyGt
kIXDqnA3oW4cExOzATbAPNKIDf/JQ/YlWxueLcgHRnlUDg420dw0D2SkwWXJ
xilkgGuPVcAlVu/6GfOjiKEehVUdjyeJ+4IjbkO2e2G7VObrVd7AyBAqgDfy
Ys4JTdPyBWehS8NwD8XtltwPrP+hosc/RC9XNEOExqMjDjrIU9BMgEDKMKT/
JmzcW9YHV7/QqEYMXICONsxuISyyMTKZ2Hp9s8jMCY1P09gfp7PXciQdlhhz
g+R5dinyMqWHXs9zLAQd5yz4TZVHj94COOYz+FM6H7Sf4MshOgU0VWiu2nsZ
eliQs3NFGBmUtqI5vauibTFWSkHcqjXQ4rc0ot2VqZ49tBNG8IaEozMLOitl
0w4HLa8a5ZU+BXO2gvkxDPs2Z3XIQijtyLtXLOTRjY6Xr0NQ8MZcGjWy7e28
m6iH48IGtFOlnxj1kOibbuYCFpPu0AT/xlga7GanqznRLKPE7Y/0gIukc0C+
NoJQYBC82DNFXYyjHIksJpe4uHrZSu00vjqggy3k/dl0J7u1S55WI2M1d1zu
FKZ71CaBnHNQ1++bt42uqvRcqqpi2jL+Fg/yiR6fLpfmOpzr3BRIMMc9C+xB
RtQwFAobFq0CqP3Id1QXyyiJB+kFPqE9rSQeVC+aRci/sC6Wj7gFkMF0Ykd+
QUZKQ58xN3OabqmLo5pP9jwenWjNPDJRd+Q3IDYw5MWdh+vvNmmLscshR1Zj
I1NSbtpuc1ax2CCFkIhEiUyCZzrOHnN9X1rGqKJerbchE6Z1XCf7SMdWz+LU
RcG7aLvLCqXSd1ggj/edPMD1CPh3Agu6pxyBkHWFjrVUPLPMnWZoYnriAEIS
Hz9rAOxcvOM6PoOOXsoh5qlRvbqioO3vMGCq9asP5fMnll4zfFI4sPzAOAJB
N5SNKGBP9BGqL+LuWTYL3Bn858EYf7BXsfO0SU5iZxrHuXx8r0NRAvx+19+n
Ohb7nQwqs17T+lbTZNXgHrrQHXMuZrnikGJo9PBCu1nIx+BQJPAiDD+hk8RU
mqJYQqXBOm9pF1SwfIweyb/HMiOkJaP/oX3sOm2C60EeJxH2gbOp7cLQysBt
AyCBToNylIanvlFZixcfKjAVUSc1/X8wfBEHDuu/N8LK4L9HS08jVLlNVfSm
ldownAFnjf+itsG9IgFSIqX4eR6W3FrsnEH+3cvJ6FwSaxxncDg2TYvOtSlC
zyQClWcEd9kqr9OoKVOVDjp7zp3CHK7jAcyiXTtlz/chKgTvfeOAGEa6iF+T
EXRh7AlPPUFRRKiFcyPhMFOD+C4akK9B66K1T0WLCxYj5xHcIWi1YHSvFLXw
xhZtiVXIvUCs8hdCXTZrTS0Cknqizc+XLy2Jc8MHAvXl83ADYTZe36I3Rujg
MqMfB0Mpqir+jY+oKYnv+Habq+NIjCTS0Y8+765OqNkPUkxIReeaga9oOk/+
MKU/CGFS5iPR3okCjG4nj85+xRcKRvvrUBlCkG7Y0fJZ7kYZvOzWqJU1siTD
eENYgeFCfrAeoOgVmAL18We9HPfbguEyaUBLA8CAx+WDO4re6CGwROdI2Gb3
5EcDfmSoZVZm1EKt7X3mmxHyrH1tvAckk5OkAvADanJ/U1PPu30u0uk+El59
F0OBsKd7Uogs6lG6gH1/hjgJimHOWkPhpOe9fKEVMnx23nLdBJmjUPWbxKqR
seKL8XqIZlOK6pDjYmsOidWD9LkJwfxVEtEFOfLTY0kdqRP65plL+wWq+5Cu
/00oltWB/+mfnBepeVpczsisfq9+x7ecKnchtfzX5qcYtEmjEZpueOu97jov
XhgGj8pYAiTqTFbFAQmHemkflelg10Kp4LpNv2sRQlkirt5F1azecVlu22aI
HioTI7Vz+atLqXip+vggBa0woOT4AOgr+Uk8DpeZ+JRs7jCjl5MunNJoaOvE
PBhwGfcf+LRI2KFqcJqMjO+srpiFBjyUkM8t7gSakSBV+XOKKdr9e6Bs1sfK
20OpG+9Zj9gBcFWEMpQ6cRjea21oj4kVwaUlxwSl4LTrujUHj63+8/Dlumm2
tvOwr7cqMqq4VLjra/BgGvUClAf1M2ob48i/BYQbDRCQD6gWaQMAq5gGq/D7
OH9Ph5qdqfVK5GUcbRRGkyMMYaw3VvQy5ksSAcs2UNC7StYrGv3QtP0KUleD
hcYsbQO//00HWC0etqDUeqzn5I8i36LDgAGctjAVafXWLR5Ek4OqTkKaoRaf
EdTndaNULiom54Y2OMPs3zreQ7TVRbjTbhArTn/qMXzdKwqBZMhpbil3vL/b
qh/F9Xdj25MmpYBuI+pivMXQ1uHptxZfEFCyZWa6t50cqwtidWPY/8MFrH6h
kst9XB0vcg94TE8LvVcmZmchiqHvsdaNx6FMq7NBSkjWM0ODaV2eG7OHJP6z
F6PA7pJbPCeEseJ/N7mxuEUIBZAp3t18FJEnGEO855wZnQ2urBRwLXzII6FQ
HNAGU4zCR6izTsqINpR8/5mq38uZFjLKnq9Kwi3ZUz8uRoyzzKSpPonDC8KP
qgc0izAwnn+LLrg2KHRnN5AEHAbxXG+7vNInYaKfdn1darb4TLK8OyxG269e
Ntsm9ARBcAY4fnVQB2M9cz0yLbiEOJ4vCfQOFoM9eLsXbmy03+IY0PjFh1ul
scMx4+0KIyxc6zo2kWNL6BCklcA6RPAMwsRNgX0TVEPwHE6+HHE9137LLtbQ
1WXT4zjU6PTW66eRQGi1iTTTS1AZOXm3g6RixBuQGoZiSs0h6zeFLE/sR4il
EodDXjsrfXLp6d9u4DcmGxsMxj/TLU3B39YhRhZl2LxL3xxVXVYZkE6bd3GK
PyIswg6F6VNfsZ9SxRGDs7BzviFqhsuJmp5peLRRxWQxBS3ugIAHu3B4UOMm
/S3AubDvDVLygVpkM86T1CLPJKsIFNCVhDBXCF4C+gyWIG0HSFzbSTMD35Lc
ZgXfnwGBNLirzuM7OOFUKHQoo+SDzozqyBm852KmLVnGBXhbXGoQCMjR3OGr
JermKXYYBlqqR4+XHniNNY3H7CfpCuR7/i07LITXC3vjDkVsHim7PewMim7p
5rUi5IQqbFCy2zyj6DBYncYdKVChLL++gO6KJW+Vk5chCO7mPmw176R6qIYt
/1uPP1WQh39AHPLoaSQ3ZRRgifHHz9qI5hrmw+tGrS9jLKtnw7Bb46zcXVJb
xLcNDc0QFOPPHz1mGqY0Sc5nlfnhmp+ZL2bNNXQesKKTK7KuIALBS8OtW0El
uCNlTaxEIZAD+0Kd3yCJdPKGw5dmMemqf4Cb2+OD2nmCtx2dtnF596MTiWMm
DP8VzKE0WSsDewffq1K5S0bhd3FBG4TiI4jEPBaQfVZMXo8UCXlRMgg1808l
Ide96v+XShM8SVYhCRxP/39QsTcUiWvRvEjbYd5ynMcutFo9mJyyGhc0m4yp
VHryZEHVB3KWlCKtsz5X9VL66G4SNbcpcKKE2OFTp5z4mRJ02hdZCm+Kafoc
21/Gahduwb8LiISD8q88odwS3if+5ayl7aXi9+JOrA4ZeiMTHBcbv3BhgNJg
UmIHhtmpfM089CRRrCuDj/wx4kfqon+kfAomRqzhH6cAsw1m91su10Kd+tQ4
Vi6yKX8kRffu6TPIucGhdQETfcGp9DCBAqFIP3hwri5YM8GygLuFaQDGbdS/
Q6GXrjx/O2EEur/ZkRyWnD2QelxPTmflDvNL405UVJcs7M7vHo4/jrs9hNzL
Iw8zi2/sPVI20zd4NNXmND4Wik6VeVCRZ1rRyhMg6OocdQ22NEQoveCxK7xG
U/5gVbyG2qsZrH5iXd6AhfdH2CJKNMyJLuLoGlDChuJOGKVu3SNF5cGr3aGt
8VJG+JcG4GepGT+SdP0rEzc3SG3K0BXLJ68V4CeKpvPWC4Sm1luT/gstUUcD
BGQsVUYvewgKe9NeRkQ8h7cr3sl/Im13EcjMneqwOp2GNikebosU/c5EYXus
I1zDz04JX4DT3W5f6BGfpJNYPpLTzXlqONkL9JIB1vK1AjDc1X83/7qIlyy6
BU5PmiBrNyR0qCF8W8jFqEw0Bxz0PUuCwc/A6ZyuHL6amuuFu7v2jPzzTeuV
wgLKiv8QxRLn1rFaZvCKigM4pDpM2q6nULXSwfAljUYoD/d+qobZ5OMOe8Vd
VyGQZEDz8rtCSasyLfAS/gQoiLbecHrDraoJIGvg7u8pwB/fUxhhr3ODWQ0G
Ut8Jjd/3Kb2Nf/FZkZR1CGE1YN9w20Ah0KblBgnxLEV5o7qnByFrXhvKeg0s
OUkRIaRk24ZLXm2pBMQOTnBAPM+uDn9du7vZbtp7YenVcrRq6ul8Yp7TbDtO
IpIlehONwQ8RAxhC55DXWyQjCGi2TFrooAUWti2wG9uCvgrinPMEyxUhDseD
7KIvTDqzwUkZztYYGV4Zkr9PNJcqbzsaYnsWcBCN62jAmbZzGJCikDgHfFwT
zpAr1KxS5XNYaaLaN239IlDBeWFPS/bX9eCPSq0h/0wWLnDpLS9qS99AoQeo
Ky3m6/HXIyI+KyaAebtprRO8d4tU4SzRCza8t6xSaDMRPy/OTgd1s6e3jwHi
QdpZfkk1XNSwaV9nYP871xzR0VBv7gv4Rp40pjH3YQd6NmRcZkQScsISe4fU
XcbdijBTG0PfDpWF63HeGZ+Ug9p8N20laHlJZ2DLb8SntUrFDVXil4apSgky
tMaAB88mzr0Ab1SmhLrk4XOxG11PeluOu4P2XobdlEA5Bty1zvNaw15Hbq8w
H3r9i0wB4dt55vJcPipmtgIOEx+d0JikAJ9EXHegUuEPDcJzM6YsvDkaC57E
2+kxM5OgR/QWUJsy8EzOOJiOxgTVZiNZ4qhEBFxs80Gjzt7op5FU8UudhAyt
RkHr/pp6z8F3VqU9WNWwo7iKl39w+08OnmQt90Hn9Emo0v9rM+VIaqqx/qQ/
mLLaaWC9hDUMeA334G5EB6WuJ+mjyZP+bX/pUua8nCX0D9wtsPvzmMj7Qx7c
SngqXUiOm4e9XWh/GaZv8c41t7LCXzsRfgPR0D5EmilOx0i+4YAXR8AH7Z8i
J5x2vIZ7+FQMcpBFrTCmbFWfG2zYdqF7XAfuIh8C+R5ZtvZdl2QMqRizmope
wHjy3k+serc7DTCPCwpT5BIH96xX3qTCQFNHXNOb1v0WPUUePsMb4Xj0Pq0T
16leinqXDxfTZp8/PKxTpZIErlrJZSTmaktyEffYTIFoJ54AvTxkxNrAqChu
RESpco9wNBxfa4fajcooQcrvm2NeaFoUGs8f01kvNfQ6GTx1G4z2g701V1ja
dysA3lxRbidjepXVKzPrGkumVnzMtVl5okkPAz98mxnq6smkTj7A/tDsmLPG
6v9sm+2kFf+RX4CDgCnnX8rKUI4N9OoRMi/YLtUU64x4q7NaLlF/pz1Vga1i
QIdjavSo2Q3KtSMPt5frvbj2pHR3CEHivNm59yssS7dLQBSl5WYrQMvKbnxs
pC/XgvVISkRXbaqaNB3QZj6b0miA8tdWivTgeekv/J4eg76HAR2PbaVN+0PN
u/3s2YsKuRvtEa1x81XO62sQNL3u4/plf2HqnFxL0J/rbAlM6h3YJ9rr4BMS
Z9pXQ9TYK7u8l9twwoeid1CwCqszaCelHMqCKt/gJgy/UwO6pXOd4sjXlESw
1Jm6sivCze7UlvcnUBWocw6TNexFz36CpJOb+6EL1YdSebpPn7F3lt1vBG4k
jL2csc/3By092Dep/T8i8YgAQs9dRogeCxNOa2MAvyTfwAKVMWBLepg95KgX
91G6nMkA5N/IE5pdyyixdF/Hwgl0ptbNdHvUTYd9tOEnM8AzStbyeQbc8Ws7
HeW6CREN4puAcl5D8ycPFD9vO5yZxCUkFxqa1DtGaVSb942D+LVpo7WuJskb
f10bLtNVFVILTyieyN0psXRA5yVrMvR521sUp+OdY7qpoHPTlbxRPIMU9nf/
dY0e9pKBt+C1ttvFBujgl/Oe5AYCBtKvfXgPqZVvCroOKdN9fk9yvMYdXaqU
uyNyWU292Kl+yyNPH1vrHYd9JLT0A4ze+P3psjwg4iPH9tiqf056VTLnesBZ
MWyyX1nQQgk44v+bxW4wdyyGdLYC7z6f24xN2Ocyp2Q6vdXw3Q4eYeoDZUO4
Sa05dZ0lvZkvtDT4qzS7mqSKfAJLWNbm3PS9HSDKlf9ZMsL3QHB+MSqs+F5A
BnNw1f7fVGIE2fkyk87nt+Nic2dNFnwI77A8WX0DxrcZsobU0aBjPsH53ak/
uNYI/Q4D/3IHnpTGWTgWZdeatRP9ye3457WPr0o+ZwG/vUK0NTHs5DWST/Bj
AP6QJA75vTJVT4kJznNAL4HQQLJGbZNulO17McqkL+ixau0tXagEfcOb3rPH
hOxZuQt8GNiUYg7NaDgkEIBJSOzJ1/3DcgWClKtMWF6uxXQIFeb+WFquUBch
I5Ddm2lrr3GxiMHV9u1XkxvLPCCBvEQM9+bME/8s8JdjLXzVBsmW3NMmk2de
9Wn9DTka8pDv8gMtLsSA6yHy19yQuzFwEzbstwiKux9zMCk3mIoYWJfr1DfG
NGX4ejfYk8/9ejBKVsQ7k5/kLEf9Y07e8g+h108ME0OcmUEZ7DESoEWEFXz3
k7iVYHfivYHzW/Qqb9HoAQPUYvWKigVvPfOyGfsBfquhf1aoTei/bpHujQXS
fnvrmVYcd5QCC9X919GOec3IL++zBV8HIAiejMwP9aWLuAxGggAn+oBIRMJ5
SoWqOGAzJuSJ/ChljN+n3awV2e4kjM5MYPlEJfoO5eBOT4ASJp2d6eUy1Cnc
KrCguvu6cLBUBNgmcpk3EMAxLGWFsM58aToKdG0xu4ICUUd+NwCbSpQcn74k
56k0+HK33bSkP4eMQGSY/kpU+YivLKgZriV1yNUlh0sDATCxQqs2kTuIvTDr
TjLzqLABLdxyS1XPM5Dt0d+9A3646TXw6/S0EUf/pJAnTDb9q6ILvAq/Fa3a
ae+npy02pQPdEPem8009lsMbTzp4P9JmcdwGmbcJ1jIEu43MMkgCfOEqAlAb
qgWeZBM2t15E2YsVHFJdTLMb/p8Pm1HMBQTt1svJKCaGLMejQz+VCk3rmoVW
onBpVGrZRztUyC3AakES5TCsNPaU04toNizpdv9ND5EolNh7JV2NNtRXqAAd
SxUIhC3NSQaaXcVvcNqDaGRP/L+YfP2PngrqwHNOP7olJOvsUv9jMHjoXC1k
iTRiJ7AyJwixGTB47zKnJJVWQ5XT+kPJTQXP4VVGYsZvMz5gtL+mmsX8E+R6
kK5yNpWAxPl85TCAVXwiGosV3qF9FtOO2IYn19R5DkSuzzIAEiQXY8l8Lbt+
57OEaaODenlkCe+5B0xKfDdWz43mvF4v4+qi8mFv6lSzBs1ilDulrEsKfNlD
o4kmmpSs+9/23BEMhXauAO/7rRMjV1dy5xIMUMGGOZy2jFEk4+/YFjzrl73V
8wkTpnIZDnToh03FmQh7A909m05UKjKUs2HlinmYiXXouZTycBTLadz4jsL9
PM4JMOszmDAKfRMhndTcdeED8+G7fDZRHYdtIiSP9h0wHeWxdFM7u+TUPnWn
FpLRP/I+3M7mosKXYU53ssCYsH/hTfeEgHSeKNxhLHyf5SRTNMx9rgul8kOe
xlxYQWtFuxiHCHU/smOoA2HMcGihEoxlhsmpStRjCRRWEOLNaQN9fKZeSfzR
/ZxSug7bgb8w5wdzwL8ssMcemUVqom8FLRYtUCshoIRWlbmxcGvQ2HscJ5LW
JTwfgrtF2P1R3V4az04Uu0vQv8g7W7n2Uy1PeQ8UxKIcBIVsdOaPlvQEJGHZ
+N9oG8vHiEaPNqS5F/ycq6ogA3Ynsnan56RDOJIA98tsGAn6Fs1eBRykKevZ
zrxbaAhjrVQuobH3qS5WxI/EVjI23Yrldf2DhIiqwYaNNMdkwZAOKsl42u/F
SLXtAvdr5uEbF1A31yoTbUV3+FmJD7OLb3GkKomKSsYlOeqXWDE5WuRw7TjK
Xqd+KCOeqlxv9vcFKxdzUCJRmVh6b3R1Z1DRI2wXvpyx2EjL6b282ESOcKkK
iEUfGoQUu9cMMXXR3FglaaGqG7lUwyHzyHfa3JR4h+pjjdxSVwwYN01CrHCN
/SijXmoGeo5a8rLExGKGmoJEujlhol0IoIpTUaoh4mwXaurfIOtx/RXObuCQ
hjsIZ9J6+PTGp4/Q7V6UGdDtMIMC+IH0F2LMOFEc5M3QuttFGTeeCug2j+pH
6G1gTsjHSWzQlv21sdqTnRgVbNQQBPpnIBc9gEXVP8jt1BaacN+6+LHvHjbH
Vkr1/GuvVtHNtc7PGcbyCsb696Gxdt3RvinE0L+wg7RCr7AFdHJx/xAuZEwp
hkQr3uHanXomJCPCeXWTvT+auvWlOj55zz7z9O7+3npv9JNxjqY4J04q/1+2
YB4GbUps3uXkdY9YJ/UgtfI0tgnn5oD8gNBI//QazDXkuivkG781BT5h4T7u
8RL3GhqnbnbHGphfTSDRJykFzpeRwplnQrvNewmcXTKqYbwZXSYxIopCGkjg
Nt+dUiBYyUahFO29cYo+8PqVJhtrIJFkM8Y+aKYGv5QzKSXOqC6w5fQDlaqP
fIz4233FvhvVzHd199tl4io9j/R0H2a+URQFfgEpIcjW7a985HqWphZM39G7
EBHQMcoge+4rA8n5zrYpdRJb63hZqmQ6fXs+WqJ/xR/TdKn8q4L3NQdLtPmf
H7ivtK0sboA8FkGQUywyKD95LpoJjQxqwIBUIg60h4ezsj7GS03Y9jgeqKx8
0mmJB+kX/qziysi88wWig2/43ohQIZapkinNm5CUo6I+/Dhu0tJDyryMpwk5
y9mjXizkVGwHPF6mB2KmStUkZEBzzEFjEaF6pygd1QGM503cnRtYDYs83LY7
9bMvwayJdcBIivFOx0o1Ttrw8SysoUAZQ9EsqDG1lsAu/X01OQHmMojHnEsi
5KiLzOVsyKwkYKy8MblxrNZM59EOogaOwuyq0oPeUDtE6AMMEQn9GyNmLkEC
9RcksVdtZBU/F5GZ9pruWh3REg3j48JvtsLXlMFz69MuhOBnx4uxH1/GpbBF
UIvX0NsJnI+nfOkcbgk/15y9gazUyWVG1CfEz7YE7iH8k//xmOqT5j0aGsZu
5+mkf5+UoHVDMcwhSzyGV+jgeajRhdH+dS4eYRsFgW4M/IKI6464WL+yw24c
Epqeqtq12QehEegfM6fKmYpqTEDvJfe43rv32fMn4lqJCS/psAQeZf5qIz4H
DskR5OCgyWhkrJEF9HivB8mrjcfN4wFJNilI9bT6S1T99kp/Zxt0vAIoMxuK
cM6Pdoz2t1TJBU0ydNe3nzTtUaEGAy4t9wq/VNXlgaOaqL8rIkbgIx1kJMuy
J2y7Q6E5i5Z/1BPGrSe0IyUDzbh5pAtxO7gNNr4U/rcQ4zi7E0v8c+QCOFQH
Rh7o8UrN4Kg2QANE3DYjcH0uKenzcmkykJjz/GgH6ZaG1TQRQTkyqIgHNXVl
KyWYDumNU2RVqcgzcf+lCJOzRKGTZiVr6dbgP9A6PvO81TqjQckgVrPAES4+
qVtGziyLFuzCtXtgjztHojAs+vAnvbAeXstrczwR2BRPcP4tjxAREa2cWLei
y+bmecGUYZaa95/qdUMOHkgy0PClmjw0a8yunCpBFcbkUfVtGFkylKM9JtTo
FH9KEVKzuei//X/l+Ortv6gDbVXpvFpKIQmCdViFlK3+xRrH3NhHx2GBjYrj
YqzaUDd0wuBKIbj6Hu5m3jzQukhZ+aFH0kD8xqgQ1T3kYKxywxIRthvTo3j1
37m+4zCozxEPfJnZtRA5OqvJZ18bJVQWrFPGEiC/Fc1VCblM9HShixE4wCFG
yPHvqDRLjL7gF/qumDgmSchwt0+gYiaBDuB4m1V//EcT6asaI/HrHS6hv3qD
4s1vL4YSARWIpInvY7XjlRWBsTU0k6DPB/O0VffCxHEEQiCt7Frwa3pq8Y0Q
LmwyygQnQVJef6ZMqVQjRywXrMbaIobZGtazKJJCHgU23NU/0mz+2M2KD4Fe
uAUr6Hpry9eNIJQhFv93QxfAsm8ajlChdf7yWcxeg9+coOM532m7cY4P2cAL
/1EgfCOgzZAIItV2IO30onbIy0uGMgxzcWTjoh4Mfja6Dwl9oO8EolmhGLCn
sTT08/74vQ4jqHX/APg8+O11jBhG+FLnYiy/k4ldfxpddhiikbJMUGjc1qa1
IH3zH/K5ukAxi5TD66/2/meV/CYIw72XbkX+VuQOuHJnjr4GLulc67cfrZ0S
bfw0A3yGldGhpLr/nSrD8c40/xUKwnF9tjj3BLK5kaE1ULuu+yC2ZiBDsbwd
ToTERZtsMJeMRrRtM3TLATUXE0PxXbTnV53nJ1mfuBi9UrEiTQLI0n+S15Ho
XV2oqmxOD0bX6jx/Cy7yG5v1G5LQdscfFtOL5PoAh+VnsUD3k4ftj/OGyYKE
JRYpDdu84fYt/GSUTQQMlIavkKn97wseosa9y/M/zHo8l3wYvJLK9GU5ebE+
4ha9QJ3RmCUMCxDyoznKcsl8sezNq9Z0I1mDnF0SCA85uoEK74kDxX5h2YCz
CBgIDvurQn+kBE3Fp1AcdD2x3xCvbYU8NNXQ1f3wdJcm11ksXq4tpewBKQPH
Tdq4POkOo2DtSWWrnoQYJ1XaMd3x+c3B2ekc+ZfL8uTgfRfiEq6PFIdjohib
jjxPSlLgsdfduRV66yAbeoVANixWVDrnFedu+E3iDtL0JSYsRmRoIXnIf1kF
Fz3xmuzo/ECo568fqi8kf9KEAweppjdPerKwAnGV3tkUvif+XtZPnDMrNIyX
NeoTixOECGP/4hAr5Qj1jPGsC1hAz9mPs44QGy0FNbykWU3n5leAhDNaV6QX
9bxSrghoMdQxYAVdLssPFEfheYax5CdqVMyz24YUU6CBepTeESapBRWv2p1G
n9i/GhXvNOKI25P8rOVmbOSEqX80pG4ZaeozBGNXhFbHaw2GOf3wa0AejQIa
iiBVkW9pnlHvlIjhOVd/pbZ7x5peZxJAgYG+k4fYJsYlYai9LRCgEo88wXdb
C5YSFZUsyRWBs+sBCIZgl6AgMYsV9lJBhkn7o2ol8vwyz8Ltg8+C+aOyUph7
LfywEBf6m2eWsYNJyPV9HGE2qh+zx98jJIy/gkT92gJeTT/a8dFEpA4QUcBk
AZE1U7J1eKdzWxJ+7Ubjw4hUekFLIbS8QEtqm8x26wMcmOhW4i0Ir2cRum6W
vzVFgFwLReF+cqUva1uLgncPBGO/IGqlo+O7IoAnIaA2QKJoTGweaYxJYzqN
+Xi9zqO+oP9HA08wNjY3ce25cR3LBdDvaEbju6y5O9HtAse17n71jhUjo7+S
HTA8CNd3/ElMn/lVydpBHJUlPmyG/nSbOVYpPsIScAxuSpa1nQ9ZY+Ym8B/6
Vwf+RIkdWnP008G/ux1gEg7pvSzMrgIgP1QvI0K89bbYbfS2W/mOn2qwCWJ0
3s/rk7x6++lxEYgkNBcgkZGGmP4jp6uvxVf0vZwrIWzBLqphQc+2NVfctREs
gU53Dt9T8xzNZRiQy5nEJ2OIo9+N/JFBj6ttBHVHuvMAxTRm92hzL6gTEEw0
9YrW1pthNLDAiO3Wnwxlo7hdxJKH9tCkl1/SfzaNZW/lUSCkMlKZApqLCaDJ
bAzJLpDbILJgsxcrM/Dw2W7bFIQp9aX6O0diQ4DeesgXSF9OnDzQORXToN05
fK4hLNh3flJ6DUokvygy78AqXazSnr3Y/n+jjpfwOOk8cH/zFLNddM8/RGlJ
gDdy63fdtVRYHqeNv0CR+n8lk5E5g2Ul7wQ/21nO6rTx3v5ekEW4jLgB66Nx
lQ4/4av5PlbUf7bLQIK3kHfnOFO+xebSkPMs6M6VhxWb6UqR0n5OYcA4T3wo
WmD9f1WtsLvRD0JoSFco/Hz620xjAwFysEyPkY8WnfUbQLmIXbhlvBI/eAK5
oZyC40yDwB38tJAK1ooCaStmEi4mZOL4QGFzF83D5XRJ0jDP0cR8B03fKxie
S3lPBL7iI0LUxmynQnyN0sZJ5utM+5fkkFicauXdNb0Gj0t2JLq6aFLCe1En
GNrSSVavyDnSJD1p03VflKHq7331St/3q3Yv+XMNNv6LQRPYV0kJp60ZtEqf
IuofLbaZh7LN48tWsoT23s5gEqSR0XJQrWtaAqHv+7JxEb4mduysnTf6/Iw6
6daGIdGQTqIZT7igC8wpHOageNr80IN4L240c8EfoaEJBXqXd+xHqJuXuJvH
MPGvDEbbDD5WxPjJVpf7OW6kXh73Ps5mJQopYLrVB/DuPNBtW0btnoh2ni5s
gjCEGhtkXKSC2e/9JBunTwp8Pkjtz+CaknhQFV9ruwvZ6yIgA+7vrsVSDXSq
QRx6FG/yQd7QdQV7SaAB5k5jehx83Lb8+2yeCLyY1gFW9cuiF1MHk09oJiye
UbGuakpEWm8xeKTGfaAGRGVvO/phpw2iyweERS2IbYcPVpPutpTP0+EenomW
mbWcB/oizJegw6jkWFxgZ7CLMxZRlrO1F3lAsA9+sE7E6gN3gJLZ/Y8XmkDM
Q/8tyCQEL55y6Vrn7iOgIgKDCaV1dylIx6WzRCVhVEO0WSnUZwxPQ+5BfZlY
RCKd4mHkv544IoWhauNayvViJXWJ+gchqG7Y95V4foN+e67dNfXsUYlQ9AoO
EVU8Ipdzema0WOgg0j6/PCecMNZBenUfh0BbFuyBUAi3/0rE2RqcRkKgg6j3
q8/4mca2Wk7UDhqVmoJuUtd3qF61Nv0vJI57FM9N+NjQR6clNYt41Pkve27e
rtocbqhYfdUrUbYhoJ95oaeHAd1C2CZ1FtxpkkWCd0QoxSqUGHPrvDNh7BTI
kCH1WZARcCdQ2lyEqGk9KYnymF1F1Xt3huxELkMdVg9HVx8QZzWP4dqZOEZS
OLHQRC2ieRS5c7I9cmNKIRKqMdRiLdMdbuSLf9LeWDoUjAZjaeia0Wu1PSUM
XJJmWImX1419

`pragma protect end_protected
