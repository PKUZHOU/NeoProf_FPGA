// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
brOlx0bUYw7EExeOaMioDhux4dxvbK4XkQykzugA+Gl7P+vutvva4YJGl3LKXxNF
fjmsOmSpKGbkaNoBzfGjppnGejaABJ+mjbDBV5sv1ZrGQbgYLPD6kOpXyy2E0ezE
07QpOdAwNN48y725TWXwTVKor4ixW7g+AOiJVjZ2oO/1HyNK8xtpog==
//pragma protect end_key_block
//pragma protect digest_block
FvgTygtnAwN61zXf0V3VzVNtIOI=
//pragma protect end_digest_block
//pragma protect data_block
+/y21kC6LUfMUDbg6Tmkoa8sVdEtdZ2SqvSwYIxNltehStFZPQRIzkAaXgf+3L7g
J9INRjqmCxDbQGYaL1DjLNi7PtneIpcI2nqTsATy5i71Hu+Iv+kbsiDKn9B5D7CI
6xP5Rul1sw1khRsbNwx4/of/jMoRWSapjAI5hvp5P7Pr0KeUxZ6vCbBB6DJww0y2
gXUPBHsWHBhN+fFMsonanCf/ciFznZE5AnvVsHe+auSnClkbzeK3hH5hzmehManN
Hgq1QP/ic4zvwBpOCYzEYjcMSMrijMAZYnzj4Waymcb+nKOwB7j2HkcT7QpdvQAr
92dszti2zzNJ+WTnVJ9ObK6MExnCbiy55QGQjCMy+2tcNsVjzS9aJncHhLvpuxCs
+cTFyNIpoygdihhyHNX9cY0EuozzaXJfUPlX/K5SQg1HW9JmzZvUnm3qPHJLUVbe
0omVhcmcLV0M8JuaikgfXSQ0veTn1qSF55Rc8ch91lpVWR8xHS3V+ScBOLBqmrWX
CxwuPYNPUQiwl5NbihwysA5iFsyYQLEl+kTvE9c/RhLSAKZCYQ3b8Fjbo/O0F4ux
QnZK22S+ozV/ERNGkZSdJvdDrMHVBhT0UM236/XrYDBkZ5sBWNHezvMByY4DCver
Lc1b09atKtkSZ4tDad5VpmJiUmryrRnvNAMywJik/rHzkEKaXpOnWABNq8i2wFYM
Dl/C3hmeZkaB81Nws2C7TJTFBQJzamB82N8cIJf7agShTWgSweVraaLlf4wqmwwk
bWGWngOiuD14D1cN0hMFZOqCtPSYQIcuFWeuWABlhvPUZvhAFmkuYUdunctMCPcJ
8GEcFgK8OcJ2LrjTbA2wKzwtl3CMvS8eFlPjr/93R6xex8CI1mGZ7FmulEY3Kbx2
9wvp1ffVikIXUkuuuCEjbXyKSQonlUg1ZtA0OBxXyBmLzItt4HGJkhRDUXpPeAcL
TtBN/8zzSE3v5UAwmqMBTrIEUJyJzKatMNpx9gLAlLAwnl+hhOH6Qjdbzvs+ZIiY
258IJotS4ge8cA6XvGEC389+eFvEgKHeS4Z78FmxDTP2Ls9YYqiamt2tbwO29W7i
kH8Hvu8C5lW+YqplQCcYcQ0lDjp1ZF+/IEZDRsxcC9jd3ilLvv1QPHc8q9R1TwKE
Lyap5Z8bOJeq85he99WkPJ11RUL0QrcSfsxF0Kx3KAwCC2+SWUUUWCygTYpDBPDH
ouoEavzEUmu6TvuWM7kfFeVR/2aLcLOMyFfDzQ8Me+lWR4M2QeAe5H0Hx1FG5HQS
ZzLSMcTvhTnkQQVQPMeJdNk2mEKI+pg+VB2q+t/y5LcgxepxYFKaszQRPBjn8fuU
V1SDzVJwBBtFf2eiPRgY9CNBd8G3y2pyEEC3YVSB75bagsSIDkSlJNpFzl4WJSVr
ZchQkPpaMYBz9Dj4fwXVgQx7dzLG9bEWZAcT+O53ziO2h2fgI7zFb0t70U8iY3C0
UJq7t1mpG51eVhrSWCIKSyn82EzoyraNZ8ECiFCEPVRxP0TEzGhv1yQrGDd3I9NW
tW4SnoTkMUGY3A+p7djC2dbwv49BUwL4vuV5M7K8qotx2cg+wlpfEJ1ATcPqhOOJ
M2fU36mqE89QlfN/R0Zn4WjXAIesojCfm6Ivz8KXBpnQu+UGWa4zEj+RryEjyb0A
vSxLoXvC6cRtcPLyx3WXrFNAenmxtu7cJJvBMNoFVOXrCy4jXIukgYXwZHaMpQH2
oqNKGaDJxFxO26EmwsUTex8D5zOslbFacxgK3uPcsAKia6OL9zdy79gGxtAxGotG
B9GOdu87dltw80sjOpNO+o8sks7qn5o1GD6E7vcUOtuDD7VBEPom5xyQxEZvRABi
g+70j+whj1/1WbdHD8JDhjVP5i/6WRxXyhsGXZ9pwUe/SOiEy/OKwrOb8YhSIVB2
Di+edHvAnPKYBOXzzNBlq2hCMWh5s6TEoVggcf7moEfe3ni4hfDj8O0Ck1+H26DE
8mP8Ra17McdkTiP2mgLPRi83A3KkXe3dcVfWE4fvyLx9C/r2ArVBjFvFaHg2jTzZ
3TE1vJnBX/rF80a3AeHd4Edf58fV/j+0YfoMbQSS6SQVkwvsktQEbkUafqdoNmMf
taZncgW0NKihJEqOVkyLUEvr3iEpCbvH5VWQGzaboBLUnkTLaE2n45jkBAJM3dNT
4PCZcKfBe+/TzhcWze6dPSDwD1+Gmq1fH4SOXGEO3XRhVc9vt3RohFVd34DOckDt
+/6SD1+BCVyg7cypRywJtaqRe2s1KkyRu+xBHdO90CJXf4BhNYyzww04tMT6tiM9
0i5KHkHkWT8wfyv0v6t+r/w1iXLf2klbVbb+52UBpBildX4NhYZG1+DvmMNOMb5b
PMWoGPjQtiF1KTjfWiEKnfOieAWJPznYHEydXyT+HdaGef81OAF8ZGXcR1wkNnMQ
qyrUc9eSL+MlccBh8oiyx+ZwHxCsdrg55ZDvc/EGFpzq5NgYLF8KQetw/Xo+L2Wf
DbJ23hE6L44iIdeJgw0r03Ys+s3ReSw4FEmTXiI2sWe80xZ2763ImuJ8wNDVBimx
chr+DPMNZHYi/dzJNu8TVM8nC31S2grWUdRqWCmGui+GhfiFMCIR0RxHm1wQK7eA
IlFAQxLTEssceIqFrkoWhZyLpe0L4nkPmz1zOBLUK0RdytjnFAUn4kCS9H08cb5G
jcSQlaQ4AvJF+CZ7j8b2u5w+iKSupFAHewXGddaLrWuozrXaTC1PYHrlIAXlTqvA
CMvdChT8mrISTub/g+qPl1aLygihGgV2Ub91FXJjuRoXeZSuXBBL2uH/lN0arSs5
kNEa20wYmr77HhliZCtsvpIZ6iFT1DJSN/QxYqFMb6T2902Ki1BZyT5x/w9k2blA
DUH6wYg1BxStgfWg/pIVHSxhJzpHjLqJ2G1HxJagkMgyjlWBDX45Nh+lCKRWUMVP
PWKWRV9nndNSp89kFEQ9c/cozEB3fke0F6B33ZPcMGabXwtZkarpLM4JuryQMrzQ
mG68+UsLTRuEtwM5RaZqvw7JLYye+Y78hgOSavtSbcpSUTGv23eQ8VEV5bzfEzNp
4dMnmUHR9M6NmZowIlBpqgz4QIOUvpVXIwRA+lb1o8wOTNkcavmubh3HJydCUcSw
xVrWRjZMHsDjETJzn9zTDRPUAqSB65FUEg8ZKWifgEyA3jJr6DSFd+sXzPsGMvcz
mlRqiPLL09NCmwtRNDgTrCmWnBxmbiKDkABP2WiE1+uZ0uSYW2H5qawwGXfyK5Hl
1YUA1Q6PBwAlXDG7OGIgYNLRLfTcdiseCl6bgPwnZxJOq4v6F5h8b+pybXse0Euj
26EWqyCtAckk1OVGX1t6PHWpgylq9VukEttjJYIryFwYPB1kbFQHNzpb/Ev6BiF4
WQO9gJKODy3+u3m3EJa0ckCSoG14G28b2HJECMhaRsIctjf89B5rGLAXy6Ge7ARt
e2o68hsGV6JUHVLcWOtE2lEVAm/rximAmInQ0cO03SMpaiElysHb14Bx6HBpNcb5
Hph9tHJFOYtwPZA6ugzke+6r98VwB93sdPrG0cgBzohipL1QhXpdq22gfJ0MfJcz
Ea/fhgvJQBOHhTW2KN6JSXbWJvVglLeQhBMV+/olNVmJbTsIFa8WjlMVHPrybEoL
7w8ZEls4b/lP94NOPuYY8U4MFGlu0Sb4tHMEsCgsisj86c7BG0wiX0cnmfDzuzVi
vLbWTFTbQG+YMERZp/A0vkDS+Ck+gjokA26lhPPiaAqtcXvqRku+9NhlQdLBFNru
ZKmYfaeHa9FaE7/VzAiq5Tee4LX0HJmCMjSVJyVv6I0cFaKyyoS3qNI5ksLxcdyy
DaHWos2gKrBMaZKDXh6BXoshU5x3FtzID39sKRUioZsOOYk7AxOVbIiDX6bZ7PFm
2TxHHrWl3sIc+W9dp+QFcX66UbGCK4lq7Zlx92Q+9UtUvwKC/7D++5NUYt+N3c7e
vhTzKiYhJCrg63JgeJxt7MCj+oNCEYIzASqfQodxCF6rUb8UUUnxhKWAPkj8dOHp
uQh7JbNC785L6/uHDplybyYqTK5uVUpCBP/fF2F2F0SIYdKgE6nXQYC6avh+oCoX
T/dlzKF3isV/iRbC5BnENlX8wzahqz/HypQo59vm01XXXuoJkNUAAY13PPXa44lp
1ieRzR7wlxYLVbH9qdU0+D/Py5uWlpAHzYvjdeZl1dWu1SELktYUAXRBIi5tOqjN
9tSCQ3kfcCTbyCmTaisJGuWMvGJ3kMXtHRbpmKYKaBPDgL6B23FtAsfzMZg5eFRv
/kuEAkCFFC/LkAnQy1sxYAj9XhNzLiMjOKeatBKCNAXSUzSMtSvoDTdRLUGu1M7H
jXgzPkxCgJK0iKRA6z3wyvW+edVyST197JRxQzZByfma+nxW1QTwYiciuj29duCO
VTNHFxOpSWOsZTVZV4nGiUFElIf9euyebgZ64lHQ6xY/uHpqwgEfHoACx2+1PN8D
6m8bygg3sXaUF1zWrL6Tc1yWQ2BG+TV9QvkJ4mgIwennckAyPVRVsKX6jX9e6UgK
OIYqpgfiRdBS1+85oTEqZxfPd2N1Yjbw/9CT5O+4YqOwGrrBP2K2M2ztn9yAM/KT
PnEDHVIXcU2gZv/aDAqh1kdNyCjPi3hpHJyMDD4j/uQg9BQ2A00IOi20mA+j9rtJ
bliJCyMwpAaOnvuRHiSQSdMOogzESN/JTWLwBFz3HjqLK8z2Tqh/Z7iZAf4wfR/4
bMsTYAxaBQPckC3QCLtcbkea8Idgp0tqzma66JgbjAiXzuMzigVfPXuAL+qQE6B4
llnAtkTVa1L0BtvbaUxuPRks0Oopv0b+aOP0dR9mEwwjmDRiYCG4Q7xZVn2sdDvr
LIG2PH76dfm1s2q1n98vDp1ELRf04I6rW2hYNPZP2TsZjFaesua73T09L9YRFI5h
YqAaJ4FGWB0GvU2erpnjUSPTLplnSaBis2tKBVUUoAfCBrb2U40GHpOvrzZo7z/X
nm7mrIQaR/FScC3GvICkrOrUSaQIax+Uzg8twsUFFOafqoS8vUGS/ZtjX7H/4hzc
oIZwDgjbBC4mH3+UIjJhFZ4XF/4FiF5nwoHv8+1NkKsLE4DfT1ceJhlGMssriDrJ
tRXJsnYC84yPuZiLHtdSAZ05TYZUlZP2LhMtsKVlgIwptc4vg1S1pQZbprXD7xnp
GchDIe+Xd7JDnQON3OVf/VdTX4v6oKp/WsjHS/YX2+64pzNm+kDOT97CBtnUmRzl
rpHQufa8RxHSj5kRgg9iRXtPshP4KHYQiNsuxhj66xkZ+QEGLPXebYWVGmACKbz0
DZzmpwEZu5YvctBd/sWW9oWoQoJ/egiyDQKOo/CFBQx+m2e4OiEm2Zj9m4Mpmqi8
nqATAc2ZcNIXL+NYF1PtANwr3O6N7b4GXn1jKwPG2YzrcqvqK7hnGqHhAkFnTxzj
O0dfWhlwGp+Bhf+ZVV4NzaZjKOf/sqcy9OQcDQDG/aEOo1bdkGxgaGIlI2/d67jG
CtooYTrGNESsrEXUGXqB2aJaim56YKC+WdMdo/N3g2WaIUcFniDnCQpZ30eVMaue
m6GMzwbSFThQ1e+ZD0J4OsRrwNQNrJoK7D0pS/2xIDKrmiwI+bjeSOeGAdEcUVFA
C5rC4KNSyNHbhFqTSoj2tA==
//pragma protect end_data_block
//pragma protect digest_block
/+eOs71rK05e69GtPn9R5LA5sVg=
//pragma protect end_digest_block
//pragma protect end_protected
