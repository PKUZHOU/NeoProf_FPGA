// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qDSucYWIjIOaewV19AZpAGbJdBsAscPCurxJIXJC+WBZ6BL1UevSKiaFZM2T
MS6LEn78AoBaBLb2faLVv8NgwlvhrHckHojdArFpX7sZDxahr1irb8MhNaLS
sg0OnAXNq28KrW7ziwPLkYEeI1onw2EnBBCvezov4jMCtYcuWVR6lSD4BAyI
pb/DpQhQVBeJAAy+uyolkELjqePSn1yqZxhN7Sg1cmsVfOzTyJDvAp775Fri
BR2kUER7GBmHe4JRmDLE9wsDaEjtciGSX6aIRlmwL5phnjopUejaQj9bxhwq
NNY2QKo1xpn5ZHWQgoy2Y018tqcOYtd1LRUYOkfHag==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZtQVZfNyZC8hX8zg9lhyh+xQ1evFXcymcdwnWR/nNy+Gpt+xY0Q2at9OXvlZ
AaZXi/1vDopHKb4rdo9EdI3t6y69Qvxsq4mAjwJlqO+D45O1Spbvxf+vzHBy
15CdknYJK+cusOYgHejLisoi59RFK8RkSt0F15dK9ZNZj1CG1rzsNzW6dobn
PGsUy9mCdrUxnfCSlvuS+FSGh/Wwkj3zkFWPnTJ7iYYaQAfIJRwO1alZ2SFp
cj+KeCl+oQ2hFSfdYlITyGU6dTjyR6R/H318QvumKvxf9cYHbzyX5DESvxqM
iyVNGTFIAGIXMRcxeBulxqVdL+mKfWT7ErCa02puyA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VRTJmKwAVx+ITCwAcbXndcIkrB4dfRWdzbQjlKyo3Im4LG790S+E4AmHy6of
kj3WvuEJPz++SXrsuAm5Io2CsUY0V3wQd5Gi6QIvnRlkkMGwdSVknNZUL1bS
trSY29WCXny4HCQAjkd5KIgaWsiQdCUELEo4XWx4UW+4+9/IX+i0YAv/0n36
1raLht7KNFZed4MNwEHsdVGHMYvBQ+2ZdCuiOOJrK64tzgop+VGakZXeK9Kx
O0Fu762kN33i0kqFO4wTj3AA87/1JzS4t7sxdFMEfhgbRJUVAlsLX7qjQ2GW
QkQooOpg7RuGvicd3bh3hJq4gR9Chl7Tpc4ddOY4gg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
gSdmY472nFYaC0NGeRpfGjASqX18oSiP04yXbJ3ZDlnol5GNN0hm9EBWAPDa
iDNA14jYHnhkUNgfWHgl827qRqMWSuNE8emhlVvyMlYgS7bKnad5a7kigiDN
QMWtSX0SvywPdGrsiVGYHNmQzdTOyOrEhIq/NO1xi2D7AcLDbIE=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
NvXjiSoLFHdTj0jlDV79shJtxpA9CiZgpnZJiqud0EimZabWBGl3RmL5vkPl
uQFohaA6hXcRXbfpadfr+O6GVv/JJwSjbccu4y8PCfWyna3DvHvmNh/nbG9h
krc879mOR9rklYX8jDJ4FX/G0c8M8wa8HJ1IqRxBFTwrnK4LyXRfLQo90CYW
XnrsldhRSvQXoCuxsDo2X6AUhc5l+gTIfBfyiq5goS0GjGVly6iS+1+a0u9k
pFfBQkJqiGg/52ZlnJtbSqDyFaDtigWF3Zo28bPuq51rPhSFVClVQoZ8nG9H
SYSk5E12N5xAuAtj9FFzkF2oh8SWRjaIAn8AQmMLMtq3Lus4AowNJ32hs0Nj
DVyGQtMtKwS7PX0lf2duRoZE4Oa2LvKs85U+aHcBgUPX88arcDSXeOGTgnBU
MQSmqLKEH7ho2i3bvj0GiUX8VjMfMSxUbLYy3QaNjFTnMjzHUvnAjOXUCBZq
fruExIDNO82b922y7KsycxIr8kRouqrO


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
fVJINVS3TqMB9SFg5n6SxFEGIlQWE3z02o0Ny2AzLwaqUJPQsFnuIdEfLfHy
PkKZkVwJz+p712bTJoZmgJxnka/GbDm0Zyr0Vja4bKCN6SXDuJ+ssFOKxgQZ
YREmw1Piszjpr5KP9r9W+xYwR3JBP7tnGOhHbtNJo8M2NT3XIq4=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
K2Ub5YmKhRWe7tFfdPST2tHSBkbFRzUKMKCoO4mFdS96HgEvBn70bmHMlVU4
Mh8n2Sqjeq2m5EFIzeMtkcSY9gnUcVVAVW5Fh3//PVxd9YOXZIS7DAVIh6FH
yfupjNpVKh6ULmfUuMjGNQfjR7jwI2RGFkrrY+6bM8If+XusBgM=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 50608)
`pragma protect data_block
Xxfszw5AmF6IhVshOLb6YedZ9sJSQ6PqJiC3OOK3iLDJbBMO+wZby7ND/F+O
K+D2JtjdbrSGxUDE0Dt2AuRN6O6UDuU8sDhXU2vmKxzMXMnRKUFfbAwDqnjU
b2r+/uk4ht1rFmWiwwLH9tqMHfXGxuHNfTpM3Dpg/EcVRSmCnhllApL4TWnh
fGBqXJNrHi9dpMavdvtFXP29+fuopXWh6t0PHj5EAQRFdP2kmJUPLCMJ8+Td
5o7nwRF4KhH+nrevm9+UARj7MsMDdqFKBFNDfOm9nl4BJKQ5iIMILU349M3N
wKysbmiIKcEKYr1avOv45swoqnQjGbFYNm/wkb5f2K/lh/lpd8OGNgpYURvi
whBtvvGfcA2oTijmtvzHfM145mAmfMdKkP2WmMQYZLeApdOd+Ngob38L7iU7
rEwdV5SnC4++hD631yQBaxxIiuey3gd5Hg4Xf4QGAkWR/x60rTWY7KacdK2J
uQt+camBYtzxgCQr0xe2TZo4HZ6VPNAW8N82c8PcfUDAzD8l3+GZhEfeWItM
tEibVvNYhDvWf6Jjz+XD9fHejHsPVsZFFHK1PDksRLKmMLJ+9FrY6AtCIc+C
mqOvbf5WeIyiRcx3tpZgKPCeKCtSKvWieokc4R7T+NCW4/P0dc0sT9ZG1PCH
XRuTdnyf5LksKxt3F89NccIgGqLURXIHAQ+KMn297GxvuH830Law2cHbn9tE
ZZGFrJ8TApe+pclVmhL3ul2NND1BVt6n/KyPMCaQkBTo3h8H303DyhZudZo+
a7g8tI/H2ZzxFTmUHcbTK6habc4+BBYLi3feh6WlV04gFIu6nRfQnW45HgY1
XQNql/glAHID6LCEQfPGVJNTjxJWmD07y35wDChyR+CuiU68JSoNTAlAYm/j
O9QcKm8s9+PiUxOBHBgwSBkiQEOqnRg+Moehj4uXyiOe0db61RvBULNexKVu
TWhqkJTXflpzeB+766Os3aqwzxqXfncQRM7guFdJLOTqmZjS1oCChU1HDzeH
tKmh7KmUN6VIQPIBttHGkX+2MVyfxaQxnp9W8TwSsezqYI14U/cqKbmr1ZN4
qMYxo1JP1k0cm5Gm3JR9a4uhKHECY3/TQeL9bppnVVYwX0Fg+Rz+LsGvhxnQ
u8dfn1dinXK5V2T2V6g7/dI5oK38Sm7jrvNx0P1fzDCGcd8sFA7LNOqVyENy
/6V1USaIkR9j2XHaCvpUe+sp2qJaXRFjYNvUzIFn767VeXAMZ0cKxCYmCl2s
uJd928RNLBBlPGRodpk2ovbiSpn7tf1aGdFMcgAfTEEIEw3e1ydt432/O3hp
RxIoCh+kp27OPHjfO75kNIzUk+LeEaOQOuzXsxF99nVNF5DFlqFdaC2PYjLa
ahgbPxUMiXCdtOmJviTW8SVYGrqCUfIqD0cfevXgWmtnbAfI7OGA4I9Fx/o0
5H/GrGZGsrOPjA7pmmNWKgruHdWFSfNzEmQ7t0ETuHIkAb1JI2Khv5XRL4vD
SS11dfsDl7+816+ahaCP9cdjHUcMHZ2gI/t2wd8i6h8Hcq5DNvMKIVEfeWDM
nHR04uRoHTFAOq/4NHwiBPTcPnTGqAQNp6wgGBWPrhRKhiUNipivXgXO1XwQ
+EVd24f2kfRrOX0SmFdEeqidQKGXGr0r1zqgBkt//bWo2o/H2iWnSA6lzYoV
HwSieyiahYkoSrMR5LQkvUbgOT9PTx3ynkjZczCYR0wkXKeHwnuioPiWQecn
MbeXO5+wxUvTjynpHyGidenIsk/9WCBlqjj2vSb5GhUYY4bLbY+9uY9V4wJl
F5WYlpm1JyF9LOKQtFGmdAOaofy+o97AxAJzgPD0PHBCPBhAZx2BzycfEAYD
L5Zi+SHY22vEqMzdfE+6it5xBYdeD1Psn1ehM8Hl7ajhkZkoivjUE3/qxzCU
EsPRibePxFqtQGdCI3uwQvq9ojBXvy+2q6j2ltLTm7WPOgzxE9Cby7YY3bo+
mQqwN9l7TcL9yjQr3m+/KyJG3WQGk8cXNd+sLsInurVoj/e3cXkuCo6CcHli
499LUUfsQarkHRdrloi1J5YmUsiFepo+efMkcEGa3+uMOcEQIDoCAP2J1lWr
lH8Zs6+eUqFIPwXy2uEZQeCtWGOCc+2HWLOMEdvYQuxjNAJHSVutnLRrCjAy
3cFwuJbdgyIJperKo4wO+EIR8VfIKk4LhPl9tFsHw6xah+LNiWn3HBKbpTiU
f9rUHHQGJ1JCnoN3jX1pvRwPtJXVd9lVNnea1TVoPgvPGWE4e13dkVFkLr+j
mBuJ7lf7t60VJzn4+C4FXfAh3knJUfYU0939xyrFOJU5QxRbamr7zgzdlMo7
7PtIn27dXZ6UnIaZJK/KeRmElmt9Cz/qOFdjC0YfB03PiioyT5TTugW7M4gA
VzIwEgZAivPgMLB9qg1dxv/zcapUKBC9xUt7WUfUr0TUDfZlt0SysNuby+uD
RThflWVPVKgXhqRmWzkcKD0L4M3/j2M+fPLuqMks8ZXzdMkpp9aXyPPvuJqP
QQFjxyrN9KVgnBluksmuqJ4uvGv4i7I4qNazEDLm3yZ2mb4d29oeiluP/hdH
EHdxZNUtcwYxELtbWL/XIEYcvrCHJJPEgItP3q4e+ebfG3l5wNhHB7GNuc/C
Db6dCbP/SlHORbZeRbDBYl2n2XHGn49RZjlCUvnJ2nVWrVMoresEUnV1WdLP
yFdJhnvHNFBhoCg2gAnVINggUmFlJBYbW/ligDpI50Lq9+5U5K30RhAy81Vj
THM3BudsnrYEWaN3ZmRA+n2GPPmMArrL3SdQ0OSieQqZQJvkFO1cyJfnWpQM
PSpCfQti3aZCq6uA7JZqCJX3NMsiaS/p5uNoiI4N4PowiZWmArfCrNIYHR3y
QuFQw+B3fhkhGgEh/o3Jjyp95Myt2aAENUUqryPRv6LzXKo+MisUCns3zt5Q
OKGpPoIiCQp1wfHN3dQ3E/E4sIRdldXHuv4/x3rNan3G14cq0rQAm04L/Hht
XylvB81TSB0Qq4eBN/Y9AkewU0m1nbnCYlO3tEw72hKl5VndNllG0lWAwAqF
fa6n2Ad3LE4VzIX4dgKuE4mJVuzbPdGoEvGaVOuPWEHZpMsH6E3j55xDrKQz
uWwk5ZkNbMcceTtMSdqhQ331KuK5IPhybzuo/aKLgklVasdURH3isX6LNq7T
YMx2jCPz+6Vn78UdkO3yVXLJGKczK2M7w29fJFb7cKns4H2IFQ+xs0Gfl2lg
w2Kd/TBcpyAkzRSW9g+XxU0JbIeYvSkZkEKuSxQR6bKp5UwhhXQGjWwH9dbZ
PEJCjv4b4WS2d0WEenZCmjLvq5TJ+edIAM00CqbSBXT1b3si64gHbxsQkHZt
H1mVayalePlagaOb2ZCdH6nxKqydUkbF5O3qsSuQgT4vhiOD+erT9cokBGcZ
sDN+GX0iZIArshzxRwdojEmVY6Abs7JRHBqCFB3yyYenlm33ZOlgA5B9QDC8
B49Cf7DW9sYE1AWt7GUvdm5LB7o5YA6Dg+5oDzlPquP7oL+ZQixGauEmW/67
OVKgrg+2YXUNKS9OG1xWiajwzRTesVY3trJDYpkyw7puYx34kGf4A+0RH1UC
bNnRptL2a4H+276wnFKazPo7U7tXTuNk8roRFXqy9PVS/6YfvzXfRkDqDvWF
yRdikiDNtD3FAIqHn3UMlTOgGdKiQAjw974yXnW2n8nwCkFn3qviLwy2AM62
/Vm+qWdEJbpYT4meRxH7IAUHzbvCTmZg1/B1osPk+BZ+V6d+VmpWC51F5ihD
D8yFycfh9PX3Y+jtlRHcApSn04UzcROY6DzaNCAhsZUYOvNxUyzgoZpqWbj/
75Ehk/aGIVR/SU09baAqn6XkoLmnMi4EbtTZDw1xIel3Yoe/a0gUPYOkQBqP
sYGGgxHVErBU6hZSnaT6WJOpF6PEfLvjJdQrn/ZxG35cQB+vLCME4EvaG2N/
Saccz3TfY+7PSracXJ1047re/FdiOC9U7OsSl3DeqwjIvlvvBgnLuddi6SgA
2LCEA1MozFP4cXT8L1OSh7sS/7xvdb+DkF21MV1Gzqbdsxqny+dF0eiMkCUU
cPrQs32ETEPvYrtwcre9r6xPFjLBmJwOlXVIPx7/6e22IXcDLWFSRULBB3z4
IfZya1SROsGnjscbT+qnTDGPCqFA+R/UUEmKAD6YCQfWN6mjVCngIcp7g2G6
5hPNEDMV14cOPXRjSEWDwB2C1sDhwXpwLlLYj3OvL+VCuTqzqD4rJJkduo+I
DlS+b9v0pQsWyUTN7Fr8loztut59I91htmB0/HRAwgwk0/qlncqUjzXAKZxo
fTDhBhsGLTdRmvbWTsDS0oTzXy9Mj/JT/BODjLC7X6iJh5dbqqvohsjARPLv
OdyuHJDB/v0T/nj8I9X9dvlJSjA9tvM6ihvfct9wb9koaQ7BpVKpys/3KPKX
SrNmcP36yp9QycOfvvoQ88YTF0BHUfvjgLy3zixInGtQpl7m5n5Qrer5Unw9
kRuYR6R/gnMSk2zLi5B+RyiwW5MYa/SCI4+tI18Oza1AVygGposHTmM8JUFV
Vpef7erDvdrNBuh0xgEn8rULR5Bl7HJOUU7gZD/TAz96w7j4fJ5RsyPwiW54
iphLwMHIhONn5r5B6eG6/1EG/Fg50ZFIbifeekqjEfSlmy7w0k92ierad55q
WP6HbEGv/bm0N3sYJFZNlgUVOXDQh9eOrE+pw1ukcb4nMf0tJidnM9fvaRTy
PIz6RA+Pn8vWWRy5RijY6cVEe2jJL7Ax/fldSQKIhFEVmEAg8slDmSXSrcCq
ecVKixPtBq/j5b8hbGXgqVTgFJ6xu1MfKbI4dZxoATwuvadsBydesU18IlX+
EiHZMtTThb0WKR3nBpIPNOBvBb+zORicsLf6uS6/bX0JnctDWH4avscqfwJg
CjcJ3FUMfAHok109+AaV9dYe2/YGqT557SMY4tpVReDn1clIyAWGNXELZl7J
6dPSUvA9cNfYXAfiUVsv/v0QEshPvDmePqxnezd9w8kqsYwiwb9rkQOwoLzX
v3qe7VjAuXB+cRTb4fOuMtA1xmtkvuK58DSdZyxY/QOcJjnNq916fFV+T4Rw
PXEdlQlsXzpzMi+sBvmXvo7byNdolp+QF/MylNmv5RZ8b0o1sRXLw9MY8ocv
SttnyHkMujKwxtUONVlEeCjjEJsr9kj0d5nuQj6VW2aPzf0NtR4L9sz0IEUe
CCOSWPi5ZFeNcZUN0nsxrWpsnMs1lF2XIjiGpoDYUfm9KRXyCouzQCbYUsmS
cpEbRpw/NNGxc6/GbajDJZPTAz9+s5XAAh/u5hVcCR2UZzmb5nJlnIcUxL/V
zz2vvuwVVXYGm75pb8RZ9XUJvr9Worldmpl1mfX/fQ5muB/BIlqu+r2wy/o5
wK7pYmWEtHHmq+huiI7bl8MZYmqw2hlmYY4Z8n2EeIPGnnqnokFjuQBtJP4I
uNNSBe7fdriL+uwrscF+RKe54AKjrOzvM5W+i9QE8Qwnbn5/TBDwRkttvTyM
anDXijm+KQJ+jLygmkBFt3/v+TdS+0oWu3eChh84b3cRkR4niRRFc/+mjRJr
CYrLNNf2El8r7lAd47yJQVcvxyvS448Yc9GwywdR6KYeXeCZ6kj8QUDfJPyJ
7XuN6trrhNpcNYcFNykLDpWo4VDcC4XeN21GjB5MrRinh+A6i1xkXhbL/wDv
GCJnmhPhMGmyzDM6gk92Gh2ne9R/fGCOoSUgP1Uxc3CDcQSgB1OCp+SOjJPX
ItSvsfjmN/EObBtY0eh4AJzhY65AN8TXQK25gmNXRstw8zIeAqGhDf9Pqgxj
Of1vYn/5rh/3fPrxwbLXUh1/wW3x0824gpZWzmxJtBjY+TSqR2OjliafEyj5
VxXse8pwVp8MgngYrWe/U4h4yTX0hh+HIta0cmTsJoINq+XfdfUoqj/PoGPy
o0VzTWreLvHWsIAKBN7zKFcBTP0dV2OKRanJ8kkvHpwLbcuu3ev7Bq07oOM6
3KJVdGQO3yKgX0fVUBg/yVOjIDxmea+hO7uq/ih27Ws7mQwg53Y6oQE018uZ
K4dFc35o7PdEsbR9U8cfCgtm6LtlSXHS9L8B/4/zueo98qQr8XAvQFfUPjDh
jWm1t4uWLO+in3fopkQAsNt3XdPC8/VtZfKiBlwB0P9xmuedqJWyIxQOZ35/
ikObUlDaHLDt4DqDd1lhi4Li3JeTeXr/dONhuQETEyTD99KCvWM+FsLqn0ZQ
+1eRkMhVwTn4koiQ9goKHwCDvwhWcHZ3rIrQ6GPsrmxwHzPX32URI4UJFLes
zr42ybwcl0v1wSFfFLj+qJ/Zw2NfNC6fGFGHNlThgtGU01tEihToOOVCACc1
V/A2VDP7F8thBZd6DdbJz10U+74Nu5kg0ym26BWflulwAXLw4Ku8KP5YMRIm
qYURaQij71MMvXLfVvEmdHJUQpe9iktSs+luRiaWIl7yPpiOufBZDnd3ieia
9GLYkx6jJWSUv4eOtaMLHT5RHVsvu5b2LTZAvoL/luOvmUAkFH1N0xyqWVRU
QpWSEQ2jMIzoFgcPkxddHBxjTB4ca1C87eBEy5fyGE8pGxGzPe8KmHhJi2pC
F2X38yWgnGTvKMbqSJBu6ntFp32EM22oUuUbuLNRAD/Y6uUBcCqeles+gubu
2K2bqEMjuYrepkG0apAUG+DGnrGBf7kwsloRX17Y/2V9EBtVYbNpaeoFhXJM
dCETE3CGSzODaktDwIE0U4Fh1BmeE2zbuggoSz8J2hpJ0r9mNZjNGO7MEEn5
6M/noYU8EgWc10TuM+vMMvFi1am4l12Sr3+3YqbFjupbhlpCP/J3OdTgznBP
SP+UMZiJUjPsqu6NocitK4VSZxenCI09akH+LQD2Tg9Ls7H1Ybf/s6OYBAAZ
wu6nIhqxwXYXv0tS6ercuoYRve/BEEGOdpw7JLkzWmC8rM216iewgxCLbqCm
2+eBrSy4aGek2tXKWYpeSgqs3ZQtJBN/xd2t9jmpe8elrAdz5rVkHakPMlsA
QQ8/uCPn5fSBR6S4fuUHZXx25h4Ygl5RHZlhdS5hHO8mZQOsYSTcNx9Jke7I
s4GXDW/LfwZuwqGQ9Jtc3vlMEbZEnoEJfZszq5Thv9us7i7DKnfkrtp6Zpoo
FWOm5cYEZau3b0JkYlsXs2ifuGJw0s8aiTocjJ23+fBeIVNbXN1RiJJFMdAz
hx10xR6FAmXhSQXET2jIfyCMym3aZkMcJ3m8EWRvptqTOANZsR6XIleoRpzD
5I00DDf1KB8wNZ2dyRUMHCJX1xwhGwwCeE93N48IQijtUj8Mx1wqgvGO4TJt
VOEWpFkm6wDwpFQOI7c5s3cZMR7dG9szm1cFGCNXWPXIYyANYQoc1yCWv/AC
HKR6doJYlpa44omXRzXXoujL8asqF4dZACHSDD9eOsNeebj8BCP/7yX4tk6a
LEQkZH40/QvSW1uDI3xOBtG2tWux41DcRKO7oveFxtcG4eUxmeLnSZ3+Nhz+
xreON9LsBjFeFJwZ4sjBzePjrZVpa/Yad9Z/xz6WD54u8bY+a+e3KWfNw6k4
xtkYjOXn0twC6g/IonNtsUUjlvsKPLO5r//5f1MQV1yECL5vL4Iu2SyExV9n
zCfMKO+onAzpms/JdZJcILBxLARee2R3IHm16xtRRmY3YEyjH5uptjj/yOdK
dywJ2MEOvOgGErcaG6WF3ch7LCDOkRfSVwfa960ObuFhzLUf+fQkwpHtkvVT
RmeO0XZsPE6rzI0WN/Q0BGe0WQrNRWK7AMMYILTgVgimtSt2S5orfovcPGUG
hkrDDk7TBtSf1/d5OvXGOLlgVk4fV4vrNzEqV0WHj7eNt7VM8IrqeIv6PTXN
P+APKyV6U8GLwxqYHgDwljCm3lbjpVeUdF1g/oZJhIiCvmIYNjttGiNE2A6C
/rUxQxzc42lDIEB5WOh+lyuMc9kZZfGtLuxSuiMhJqwFntmrKrV5bHos2CXg
Ku4rQCOCgoD0uOiQ+sqSsZJkZ0m5Hc2YLb4l+pyyUiV/VhVDhIKWsr6O401D
Cipjk2piq3AA0z3qcFf+htYJhj9SKKbPIcGJ0R/eFzgjR0c+Holko0DJ3ZID
aLrhx7fc28/egd97KFASUaLkwfPoYJEwuM6LrQ1VWkDMYjFVnXhn9lTr0XBG
FnniNR3bmTb57YT+HOoaMl38AbpNEy/cMj7J99hNIplN0WeJqcG0QtBzW+0R
eI0WfVXhvJblrCy/dm0secEJCHie6a9oQEnNhS/a96A9dt+itdEV34EvODIN
BW46qg04qAwXJ2lhgKGRynuQLLg3CU8TCJGBGujY8JFs7KjRzJzccyeFqb0M
12SRcYAbGyIz19LoSwku4eMgweK7TTZWdhlJgbhvCA9WX+IjsWwkmQvB+5Nz
W4FJW82BcQ8At/sM1FjJug2RgCaPVd+EeWFb+QdUFJ5IWbO7Su6bP0FexsGJ
ORvY35j+wJEABcNtMdZTFpPhntLhGbA/fKHqUQLdeDAC5keqsXDU2A+8YPMf
qKb+tG8S6kTBt+fB2qDkR3tIT+C6DnjIgeXct9pA3tpu0kjS6BxdaOkbXpP7
i0MYntYo55YvnwKgToiU8rvyuPm7uSl8FW33eVyQLB5t1fwzsYbcKt8B98uC
fYPitAppt9rh5oK0cukGgOfP+2dnehrVVbB0Cmh3ZU4YLqUGDDnpM8+FX86f
Q6RQwYmPgswRXfQggy5U817hdmXvqbTqgv0Svrl6HP/0UIJFajic65Lyw+GK
8lLDuVTE5w1cPhG78DKQVfzWA7nw1i8IAP7DClbWm0XM5yyXXJulUqqCL63H
57cWbo+I24E400ShfiF9fFV+TTqFtaaXoFIEVvWi8ADIiCvi2uhbsplhTtWQ
qWq4VG8ZH5+anbxd7qkus9aj+xDwLevdmxgPdp6CkmHGNzrkIbivbvNKWr/R
t0XBEG7Bb7PEPJqMn/lx2+A2/GLAY66PiE0xEEerJ5nafP2KM8y3+TxTgRkv
qPMOqtk2PD9uLdG0h/h6ZN+xGFdAOQVWafTgrNbuzaOYhY6Fd3E6OjBBtVq2
6yJXCWWfkNnQpSKMnFPGnXWQcb6ke8Y27CkL3GpCbCqqnC+l6ptqS1ghxyu5
ZQpPYYgRYGhWU9zFMDNsmF7QN4qhxDRGb/Uq2EoZD5XKgev94XlWm8bRElCc
eqUbpPEL09KL88LoIKiHNX9OE7cEj4yO/e/dnfUWQ7kTfOpVQuwF7A7oicrB
fJQeGOgfC2g9ePGuY6Q3EsV295UIWRYIpa9gzJirttn0QotQXkb8/HiNxzwv
OaOovZhoNsnGUPlGqZtDsXJkQSN1OGtlux8zi/CsjTkkQDPOVB0q5F6FhOYC
oNMU2yPmIV4SWc2bSxFJOpJ1mtRS7T3BJs8sb3/E/nhmWBkh4DOD2W7CfGlT
eq8VTmcShAYRAf2Vpc7PNcWNYpmIHo4/n0jf7yU/FNWnW7L5Ua9PINB1fqVI
52x1Rr00v/EsA+g6auZjE6kIS2IQlDAO6KZFp+f+TEAU32GumhBzmFMWpUSe
xj62IFin98CHZH6ERd8CG1WukZ4QIIpAuNeQ1lMiWj6oKt+AFt2JrvkRguwO
r6umtrYIY0Q6Lj/+BGwCHna9QyNHHr5qfAD72M4Q4Z98lLIcU//D//+ECN6k
Kq6qAWQCOGXfJcSZlB8lhGndV/eDtMUcG81mm7gsXYf7HgKO9XoZqkUoy/SL
4tct0GXVQbt4psoR3q1MRd9JURDfsKAMmqcEItEz+I2+q6ORMnM+I5xdnwZN
ca5c80kKHu6CixbBpx9Bs3zCTz+aSTK01PDSWF8QNratN51YOry3KCvKpkhp
27iK4U0WzKtAGE1KC8i0FnKdyvWzYhsolP6zKsL9vfZXj7vVsDt1xDg517PR
bt6KL654KDU+JAD0WugmvH8XBxEsskVyzNrjKnvQSCzMl4unyPItrYJpLlV/
+P1eR7hrCjJfNG5jNCT5JcWniniII2u+5FasXmv8Kk3fF7EXVEZTQgQSBBp5
3WpRpX0hm4hCgDMBwFUOjKgobmEUBOd8KIncMPG1Bd6CuP9PuzrogQLOcBLy
f3CA6iKAOrmt6i5x8TR5myqfGw/08HL7r67v/x+GXxno5prnHi05j4KVAz0l
3H+wJ5kH1zkXx3EvOIc4OPbjg8Eos3j2BptTxav1iJsqTNtXX/xJKjcS8Rxz
NOun4Tu6c01rhLE+teIID6DS5p/OmKOccl6yOJ2drX3n7tAVTHHsYZHUP5I3
eOGiK9sVATgOGl1YCgxFCPv+oRjo8npoV3r4WlAKvdpg5sVImSrnsvfOy9Ay
T3IV4Cm8xo9SFbV37LzIBfI2+LmCML0qsuKYwWx3EcmX3yQk6/vkAPTgGS+Q
qnWw0Xkt7mEiWx7Ekh2w7qgNaDP09T9HU+UlSwtlD9LnVEwMdqQ9CkhU+IBE
9alwNLWVyPrmribwtxl16xN5VGUBLWCoDJ1HuXBie080tZvPm6JiOIAt4gaa
nNMXZFtDfblTUac35+mRQ3KqWV721FOsnM4lHrnf2I1vdGc4sxukQxIfXx3V
FArMlge42TApFqdh42J41+/QBIAz8dGqw0REUFJlrLnA/Nohf+k+b6tkFt7/
oXV/1JyNUFw9oMI06U1OC8uQBM7sIeo/YWRVj064L6DRoR3r+a4I3EqMfWxc
E0TREkckQqNuviG187b7yIhLmz9a6n3zm3beiXBlCkkHsoIonkI2wdrL4vnu
r0DRuNytmh/tmLBhsyliwUmCeJf7hFx7JTIAybz76cKci2sK3FlxpPUVmdUl
WZ1jpOh5ytxvSOR478A5MsUBmaRPIN4+nFiETpvBVo/nuIXFjBrOtFQrh8sw
N/TPkC4H1t1LidM5rp0d8K4N3c2ye4hUov8s8c65p7lDS9sPBcpZuwnxcAH0
dzgVhKyu0begnxDHI3Ib/jM4jAaDwdDIqrMDr6aIimKXNt7e9/Bg19yQu+au
134lknWMgpNVIKaELkzxJEKRDuykgL+VLArLt5hLxaebcXGdlbU4pHkvy3RW
7/xQHeBMRurRAclt+FOTirkd6RhFgKCtTluOoY52fgYBczXBt3hG2XLFcoz6
hp8fQuMutkMHcGibQZjaSdWWw+qlXRK5qALmyEDxY+VZIKDVNmFKPKaPgCe2
d9NTU54FhoJdpeyJzvwD4psgFBwg4uIaxdzC0n9HI/z+SxOxwAM7gZPVPMWn
zekLddySBQhgXPJ6MCRlaIre5AQxBitcS6Dzb0Fk50nxuLhzrltNmfnzDqjY
hgnNIFg+cIZKF6+1HRnP/X4JJeKyGzVWCrINBbiCWrAXoecGfi+S2D6++aMJ
jBZ83Ekf8zLeyPUeAjCtS+fFBfazA1h4SJTgBQQwPRp49yh173pqGUzqGO4C
11pM3p2eO/NeDp8Wv3wgENKbbc3oBbjCzkGRHqEIpVeh1pRafUpsdK3bQBbh
YSv2e1lPeLX1LE5HAcSVADsnmMIQTXEyyqpXN11SeYO43/ebnOWpycYz5ZKl
8KBSkN7r3vPhOiDGk5ECKicagbeohavWxtS1QZNz0H3jVMf8NRvSRIGvbLMX
94VkD6KvmwDNvnufgQfhnZYn6fvocMPrBPbahcM002HL4YM39PSGUBPWvxjV
bDjxQ7w1Ss5fGp8IoInj/pkhmEt3zv21WOxHvtrnEZfFOU/R+iDgkRxlwjBw
fGYyqwpK4N55l13mXStmyrPo201jjt7WRBQL6STeLx9SSsJ/Sy+sMEyOUYL2
qwtisKrbBYEjYxAS+EtOpPGXwOg1GdfepRuBxEWrHk8KKhI1TLYsPle6hJmB
YHW0qPH3KENYMtqXy5UIsQEZTrk+pV3fnjb2Zt2VqOW/TpEo8/KFG2a46zRR
yBB+OPF0kMtEctwU8pDCZe0WMz+jkVcVvkfjwVNH+HUHXeRgblG2+W/ZgSmT
1kMqXiu/UfaHVBrA2YsnF7GvSxcEj5GcGI6wTVtRfQW2VvrYHGp6CHpTUmwf
UgxzkpJaFgG7JHsnH5I3Uo9Bep0h3+6+fh2cPhgO+PbpVUszwDq+6ANMIoQ4
9v4l7faCKdQJXbxL2bgKqVY1qf1EyqwPIrZGZQB9U46yP7WlPtFzJLjiVY20
wCXWX2Hx4JqDYtdtN7Nqc1UKoILFxHUyFc6x79ZTfwXvISG7fNNUwssMrlP2
6J5+Rqn+U85MxJVRZxlwYDfsSJ9zZR/kYZtNUYX+h1p7o7gQVRCPuOoVjI9Z
MT5kGGQBKJjnbwP6BjmOI8EwqppULu50Rcs8S20hexH8T1KN3gDyWcrRatI0
Pv3/fExohEoakVXq/0PYNuvHe3RH4zV/BZQpu11ScjUVsB84V/ENTT9TWYnO
e+PWqpSBHYLHn8ktDqSOcATvDig+nXigHNIybizpBJxVK1EdXFex36Bb8spD
T3C895Bybp6Y41mHg+iQkbnbBR7b1xcEZKp8rZQuwqnnfjZeQVPvrHeX4zPY
3aOxg1RRBP9/U0dAiLcs7T70vnOSpc1fCdO6ctYB+Zo2/rtHifTyivirfOHK
7nL2/VYxCIEwoTfLBc9M4eS4REEUvyo0hlBy5lvK+5ouKO6By1g4+Je1cBgC
QHws4UhzuBg9DVpDQYMUC91laAL3+rUYa8NnO7FCqUbkTyZm/A2MEeS+rVCQ
38gr+PpzRT+L8LT7yx/HdTiQxuqlhWQR7ChrUFkv2QMnm191zFDkHPUKO6Dv
MrmoEdEUsS10ygMbe80UMnn2mItVIwrx+6B0nhfmgiVdoOomfYe7UUEEMd4T
Cpla96ZveJjWbLZOLuAMD2HUfNTmXxjIs2ATO0aBTElLkJXj0rJu/CJXb8Zv
6NBAo17JYCdOPzR6LwCWPyojnPl+7zODnJ1p84DLgmHW09UHq6xJ1zbzVFnE
JZ1g+vw+Gdxeh0rpBZvFx+WweiFRhFzOxAAmwhLuQ4d5/jteDQGdYgthZuMN
rZNGTiR/OckHS/cf3esUUd4H5CVfEFHW8J5ZmPMSYuHS4pp7fwU689b1eaYz
FPHwdLjWSATPNr3ycD3zXgolBIpSc+edOmfLvPY2nbEtOmfkG24dj2c+zHg/
VMeDXskO8RYLUjdNU5Hza68tojzRc7mW84jlcwfEbDxgjXqENmYwgk8FoRMo
fNiYmCofENsMtm8fPghPsJSPyNPhlFEOpum2SZYph1IxbHrp0WkJuRXSWSvU
tePIBjVRgvqeGw7Nscblrm+YlqidGBMKZv7TQQLHUNNAmjfDODOADS4TrjK0
BrZs7v4gW9EACNufFWrtnD1KHlQp9rXccK10v4OA7L6hQdoaNco9CQ8yNeFf
+tx8ThSAMIsM9sJmrwZBQ41A1RuvI//1r8F/pMSlFCk9SFMBRjLz/it68ZoS
jjiRQGOpVvDUVAijgUhZmyzRw5BI4ULk0NnP72+ceg1+upkixxTVTtHnuahk
2uEsu9dfKPqXejC6KcNA9E4XAsi5xTeCKQLQP8CqP+sz1ug1LyZ8Zs8tjnBt
i1MVldJhPnB1q+viaWdNX3UR1HqYCQGXlYtKIkJkvxHv9kVFxKbYQVXEbhBz
BoExlbcfun1nw+RkPeb+yxs4Mu38LesVhCCrjn7IXAOENSkn0/L4DhlHXO6l
HOPhX6tzTzvdIhaqRzzJQqlubBmhXDfzDhg5uTWWm9nl/1WNeOcYKq5Lw23S
4m8GbDI3oFAJ2nsvdHAN5aa6IItEW0mrwXnqWvP0R+FouhVRUbkgmY0CGDjQ
n4lxoZKyJ95qiL69WErejngPCtSNIEkA1tEuCZ/kiEne9Oa1oh6xVjmp+e1q
ex6Ay2+boqAncMedkvLp91G/NADNFpitlACN1iS462SH2LZUD/eGi18AfQUX
knI2R4TVYkXjd+MSQ/uNYizh6DcicPowEdtFaUiIRMmgd3yU/1IxeKrdL6vV
/48FwSm6pY2yxtwNAhaJBCP6YsumQpQJVA/hmjw5dNzz0GJOJzm2rSNqkLRg
ml5v2Q1pDTQEYpgGNi7fvWJbzkwOEHkpFaUZOlvT3IWvTbx7Pn1rFptXDtCg
pBjJmx37P6zPT6OqZxh1025KyF/yLHR8qJ9+ymnBhuTIy2/ihIlkBnA8RJ4Q
QzL2NDEBve0rbJyzfLiI1y3ZvqlN1ByZsyIRH9X9auwBe8V3qUC2aa4a69jn
irRrqXLCg83RGwmrTWGgAZIpxiOlZqt/FKDUacmygY6VdcEFGlfLOPPPfS+R
5feyuQ+PeCi1hnfXr60xhsLkI4PVxE7qrW1KKsb3b2D4biptKYNDXtTSdpzY
PKzfvWvKmApR1iZG20V36LQyXXnV8KBGu1fGyaw+5fIl2NFWRRiveNcOvTtD
pQPhknWMIBNcZkDUld4bIL6J1wHr0DeYJgQA8qCoJUYLcb3R/DS1a2Cx9MMB
EjddAjgJ7VieZktzrwph+/mZsyVezwQMdvfSDSzW5VoyIyHzgvAcERYvnbzM
OdiT/WClNAdROUG8+r60SysasQmyhIBbe3hYmvAJSpMYtOOlo8gG3ouKzdJU
BaYfUZJzLxpVIdLeB1XA1EosAVCxdRQQmjDwvzo6WCxGjHR5IIyEzKblqYw3
6RYtjjbzxFjvvr2DQf76zshS99woATEEKJqK9A/rDuyQ+rv4aKKQGKktRdUN
Pely40o/cySrQ8Bn9f/AxkxlrvpdR/EsNhwoA9R/w3tzZtSBtjk3ye12gxOK
ADRduuhof4l0IIgLoziUy3cGH9k50PnXXla6vEWbQg9JoSuPhETUKsZlHAJp
vhSgFQmjC57bzV9K8Gqx/rI0tilrFsBWKQ18sUBBaQh5NgG7UroZA+C3VSpB
KUS4QRrT4ZDYyMXqFELLj1INTdgQsn6Ve6Wog+RrlWdwZZIov1psdRrV3D/c
S8JdsgmdXq4IzVJ+mXWKWQ8Tct0mfr4ramg0fb6xqp9wq+4W/zXti27Dbd11
flwNPDL3oJZjM52ww/6wcVtvv4+DW5ufA7W8LoQeuutD9RfS2eCX4tuLGglL
XRlE/xIcP4ZE6asm6VhkVr/NVHOEhYXZLQC55+OAWBRNGHaQq5MCYl5zOuv1
XX6ZvCRFpVE6IOx7NM/QRqjwjyA96BhqA4IhAxWhwb3LqfzF56yq+mUOkj5W
T3i6oZFRllavwxc9U65mEAysZO7idZ3xr360uFj6IrqN4rV+d6+HmqLSPz3h
Uke+xahALeL374fpthDASF19WHykcGO23WVo84fedPZntCI7ej79P7pzeN2k
ZqGCanWZPhYg/XSU/YJHY7HpragrGzc2XTT05qKj+OSrC0VTOevRJMRCog2m
Fk3/zOLNbdIAU5lgXUR71f0U6My4pn7tQY2Y8n3BORI1vhOtAnguOPXEjQVE
R6EWE+KbNLWMoRCP+tUiRErcMij36b98vqpA9B7RnRj97/wZHYEFulPKnhFt
FHo6v7wdbgUQF4E6QBYLiSexBGJ1m0uN+bK4wU2w5sF/yQNs/iXvI0scOZGA
tNyQUgbHmvHkZHGQyn1899ETWV1dY8gyx+PiliRmCE31laP+qyll0N/fDGbb
gNcmc6COiQSEW1rIk5VZ6vx2kzKKTwbY751AmNV+2SnvwrVHT0TO5fBH/K9C
a0AEmMztlGynIMKkQ7OL5KJycdgSrwbXsVreb70fnm2inMW9az6coQF6fda8
BAmFZ5MhOdR5T15SIvy4ZabjuzJ2GSD6W8lAV5gLJUBlfTgxhjR+qC4DityG
SZSlq8R6rBKF0JKx2vgGFg/pzV9OEmC1swqnZTwskZFVl2BRfqz3sLlFTC5N
hwwxwnXgdwwymHH1BPnTnd6spSldnaPa4BEhAoG2zMVgwpRR9FijCXpIxyAS
nD17ToXFRPcg2x/TzPbe9ie/gBc9hJjxKiNmCsbpFLdTwVbdNHiXWx9AO5ob
3xlQkaRqpXWCTCqPfCghX6P4StJXgvCRVeA4NgV8EDR2X00BCq4W9KQr4JGD
K/Y0V/cxA8Yvs0HLmdlRfDE87BXc9ZLAVRy0xhD/b9B8bkB0x6OZ5YHFXkwH
C1iVrTWDdsJ9cQ659PMy4BIDue/VHYpUGY6IIeEk7m9zaZYVykA4SGkY6db7
Wqsq7HDlGSmqrZO+IL2SZCMP69gCLYRedZFOuLOACek7Q9NAG2cQ9DIi315j
/iN51xv8g8HCDuwlJ5blsuo/Yw/xNlkFR2Z5+qyzwVgaif4HzFY4pSUwyaCC
E4e1TljJIb6d4ifwEpccqIu7dJewyAEGlc6mxcL6iJxMAsCOOJDhgmAjK1I4
ds8+E5lqpjH8TWBzZEgKYe7+OYlOT6U4UhjSfUzrnREitUzBZJCnrmQlZSYZ
OrUUHDNzDzg42ijC7m3YqjA9uqjMgP+qtEFzAoIgbQGklFXPjPLxNex3WVNn
HphZRI50d1gwiNsBDgXBLdG6B8V84rcGlBeu3t+WOWgIuJDGoWlq3WduuXEm
cexT2sZuE+8vcl2iMDVBEMMNi2vnMp01RKeCEWS97fq2YVaifWhFgd8HrUeV
paj6/VO2R4kGaFvkRX9vhFK2Tfu98CT9lIWokI4SryunNCrzRECg05/yegiG
rYXWcGiFBVNqhCvjuCqcoqJ1jD/6OK88/rqcpcJQmn7FZ7X4IVrfD23Bl6qZ
Tb1llNVakyTSRC1IVudqz81Wz2Qdg2aA5ozBciZ8v12Mp48ibwCNXVBIt8I8
xVhxjXZN0Es0OGCY4vUDoT/+Ae4WrGf2T04W/s9Bftlc73rivWagPDJQzaby
smBUl/5Lxuz0Y1zMm+3/U/TLlnpiwLRXy5+UCOYGkBApvgtAxB48WEfQhZ7L
O6qIjP/PM4FOf2nEojZNKtCdDoFXzw/rP3NFoYX/zX320GhJUylouV/phrEB
zX0iXHQueiKCpRFRsOoz9P4LaH+1k/OZahxlmjfiV3l8t/cxMBJucWTKAYW7
E5Mg4tVTx5aAiQHPFk+CDrKvMVSBoHFeJyXjYLSqEYByTEI+rUT71nxZoTI5
5jw0ae9aZJg0yTfGUI5FNaLUt2ZcWgtGnQsfdMRnwsCXWBrB+PswUAVWb47l
LnetjO2C+UljbvIIQKis6Ji4hHbmYpb87gege7oV2jGQKYbaW33RKUM864T7
Q3GRckoY/KOYrR9aFlqsuKTRoagFTScmrk3zpvGFPElQXVDNo24s5EbfjKVj
O/hAQ8Tesf3aDKvYTsHuqnhxvCDNVbG7kX/kJADREAMMG07uOmiZADzFAeDb
7LmL1wLpemCkadN4hjkSCZilndED/p4hZRMg57tbKIpHgydG31DX9pGjLF9H
J1xvBUsyYJh7t1FrKpvwNfn469MKMka7233RsMXswhyz8Z6fdw1flUVnVIkb
bgPJOTU+t/R9Uubv1Pyrf+gvmiEkKLV1dVXMaEvuXb2KKNtwpaE3hqt7w8Xg
nxnSY46St4NUvZSZPWHmMICIJ2EIQkN4d8zNtwrZjDKeMSCjZFcpnvLdeNJ4
byVoXmLnwNia2k7IWabkcy2XfbrDZbSGchw/g5M0yQU/LytM4JokeQQegs5g
5DMHgRuSi1r/qaycb2oBXUUwoqj6VVu/Z8GkCxi/EQlyKKmr5B1d7wNnmfui
SlKJls1wtNBbl8yTeG0EF4yAmznKxwhcp1hO+QrhF0DmVg1f67MPsy5eRzoC
Tr5uXdOI7w6/q0WIFEqur+WPeVVwy3gSujL+bHwJMIAGkU63aijz3cpHuf5T
v6M2u9mRwkPSqOjsKkyGXwYnqpEnC7pRhpkhhdDdTCI2IlyzhTT/w54e2V6O
+FNZoW+WqPx8Ggf+FLXTlLJZ8ERTnYwtEzAH2KiynNF7sN9fK/mRnV5zrNQy
kMooa8vFLXfsvNZU9/xurv1PxUGy+EqHtVdhrqtZ7O2NVEii+XO3HMwZmPJc
r4Q45VtW/LnrcTTI/BKtcry/AC/SNRZxu6axJmMKFI5LfRbU4Mu+ONJMEdSS
+ixuBi+Mjszm+2v4ApcOCJSQ1Kps7W1UZ54iBbkl9V06GPuzMFPE0Cbwc126
nuGe8AmrEPMK4f+CLsBPgDyg5DTY2S+NQZ3Akd5+QJXsbH24L8MhOX6B1WBG
bJYBQ3B6AnxdChEb6bdl9BoDAUaioP386MZggBBZ/hNnHxPyyaxpvxQYFjlB
9r5aytUCqMYn+NM+c6xRkU8pZ/VRvv7B8kM5lrmkGZ/Ra/UeCc6CU32WjbQa
EZeAnXXLAMSglwM1U1oMT0olcXivgTiZi+TDZsueTg4PxLAmyjU1fIS/VR3p
fiJbRQL9MKAm600Ux76iYSp2ak37hKiClw+rBC8hk5/vm/MmDRLS91UqKRQv
vaqmQxN/9FGEtLvzBqVbR4q2bTQmFmabBJ7Z30fmDkm2EEon6S97a3Od2fpB
csYEWxsTUeksPJIlteapuW2OWcuyeR0OZ/mwOGmKnMlOq4ls9vD6HwAObmTz
G0Fa1BdHpHrWcHjVdIUSfwBdM4+mi9yv7vFniHfoD8AInKtF96QgIEgN56eE
/6c1E1nZRC31vLsj39xOnqTve3Vrr04YS/cyAVJW18lAf64TksSgp48V/Ds/
5oDR0pykNz5wQBHMguyX1s7Y/jMPCSxu2jkCJ1WEGXzwKOlXX8H9ZrhuDobC
he4Bp5MqAJQ7gwr1i8WPaPiov4ixLwair8vU6JAnWQlK60pYnReKq/CQ9Xtj
dF/jBcBk0cuNJec/zX4GrN+OozPc0F4cFsrNy1OA4t1E7mArKu+fjymnQ1qE
0HWJaphswNN538nGY8lhWwF9M/kevliVTC5CDKE1rl7gYlp61sEFygbnv9m6
B9Dcxn7KbnJhqJRkL90jYzoQnPLXeuX9OpzzfCs37SV/3rUy4GTiWRK8hWkt
yzctnTjT/Y4Gc4TEBdJ8PBEVX+7bJl9XAQEO1h2qAIHuyl5s6VxqJGnzA/V6
Pv8tOeqFtPdZ9j0hvH0SGDqUh+HcYZS6oWJ+EltPS6iPiFNkwv8bNVajiI8f
NuApWfan0fxxmksKyUfLAOMtSZ0tdewCsWiA1uIe1ckIXDDx29xszm80t75m
crmCIl3eeizFX676CKyMmFcCxzGolsImVLacaJ2JRmmFjp9geEYn6hLWyZSE
R96UYqMYaokYrrnsmtFBVk54r81/eAag8prMRpe33LZPgqhblPLK9fBhOz65
vaq75eMrZkCK8SNiqee1w5kaV8FcoHf4HC+t7R+cdQpHjauDpG8aQYVDDadT
0B7dyDkSDm8eNoAt6+v/VufMLbH09bFl1VP8rqjJl4hG5hLtm7g1YB5T1Eu4
/J625jwm3BT0o3R24GNXhIsOcxe3enRPB3xFXqcRcXjhLf/KaLKrkoUdS8jF
MfYib6kY8a/N+GL6YPrWIaHPR3FequBQ1PsrxT8KQTYHqw7XbtrfS1n1dk8S
Sv8XT2OkwlZL2CwvvKFO02s/FhZHtdMOaNmbGecAishVMEat3PMsiLEqV3jr
uyr0ENV+Yw4ZfPf49337oB3E3MwmxwAD0JUsHP8bLCZE2YQgigFasgd0CJZM
K6RVkHsmMNT5VZoD38ysagop40R8ZCKg2+R6yUb+pc7vEm0s/oBgLRR3swBC
Kk6HbrAvcCu/P2P/nFlr1FZYiHkvciJq0YdUqV869bi+8iiUzks/8hUHrrWQ
Zio/NwmzsNtvWtDZsy7nPQ/tj0Q0TP5CgSBzkPQ85Eju8LCsm4WFwRToV3Oz
bOaMtJcRCi2dEQHDh7V3DDxC0Nj7V9mn5V/l7vlfsgGkGUXB7weK8H+aXVSG
0OMNzVj/cv+p2LX0IYQit8Lc1MMELZH8PCpH688yEyhFmccyulbSJy7mTIef
VrYCjjSfeZxfXm9cdmgaQ11MqmmRlnMtyc84M4dMaz3f1W/ZYDUKwzbrNfEZ
Ruq4kKTgrMdfcmB+2XXbefm/oZhFJPXTYV6B8DOZgD8dGzp9raLyTVYr2jcr
l1LqkU/yZLkkB75zioLc9+28fJGKNbqKIypwv3gEgR4KCQBbmod0oKEkjQp5
ZhjX2yikTFvHVIM88ZLU8j66iMi6iwS0+LElnc+8iMqdng037uOWWiN1oBgV
5Ze28ZOJ13Pkubzi8qKuHk1XYq9gJNi/Hh5O113MkbPXb4mZvuXUCtTVZHHs
MFfH+XSm27+a1cZavUd20cEQROhd/H8voNXZD2bVElXN8zxv7MrKziyIc7eA
AjIXBR5Tz3ebQkxn9wUInyhVRNKK9uIBseflRZmllh/uzwLW9ro7t8tpLPTg
xVEeA3MYRylvtSPal6kn53NhbPSbeZ9/a5BAhhICaxMId81odJQrXOTbQFR6
+IkqZhefa/fSy2ZtU4eKrTUEl6jKVvxHEVS0p7lBI98uD00ZAiEOgPyEqMFa
VL6qtuYDdHglV0EGOuFTcYC6qY5nvRx+X4CH6LvyQuq0ieKCHwG6A3E9MphJ
7jrwEaetu2C03LOY2TBeJ0EP1Imjg9acq6iwH/QV1lcrHP+rEhnhaIk0AjfJ
wf/rH5bWCl6aZWkp5EY40HTTV/gi6K0xn7sJXpbxB70flIT0FXx27sFI17yB
kO6K/1L6ToNv3hSM+DfyOVjbwEy5GzYia+9r77c35F+5BZ+nL2twblxN2YLN
nD4zpxoQJbgqBBQ/1zKja7KkSnRGzIHDDDSnAgz9K7/6E50HB9UuPwCJ5oXf
sbpQCNI0NTniVGRGtfv0gr6nOe0aK9P3Q+oBaTBABogT0aRHYIxxvlB9Dg5u
ZnsxN9PWkbx4R07KB97tnwc2SEnxXPHg5GxCQGizCMc/em3D0fAjtipkjzD5
rH5vkuiz5UicGzIqxmR9PrmiB4kuBIiKg+lzKAJEMFMXqaw1rje1fy+i+jfq
JzIQiDoHiNbOUOVHZPRGxB3A9ej06PZFEOh3Mj8AVSYpmRFYJxO4UxoJyDzs
XIp7dci82euMOj059IOgks9L4t03sHU5mIlrkHt26CTSVKlHhBME2ck9qhew
goNrMf8Oz/AQhoEwbSGqqCBshYijJEWcd5syXHFcT7pwaRdH2A+hCRdJhZHl
ihNPa8tiSkJqRUweD1xidfJkupJPPprC1FM+kLjjVQcmzbg694bYVcDU+bFO
HQJ1BKSaJQogroYKfGYpvmdJpfNqj48U620GnN+deylnyKscIHl7O+9LGgdH
2btWS0FOH99O6rMixF9R5SPo6UFeEXollyxWzk9jc2zJqvWDGmHYIS+6h3Ts
2tRs7QXnuQNIABEVv4iY2tiNkdcEYNSmkFdSPLjAcTvhS1yZ1hbwpYC3lSrd
phaZ6Q4sh1Izq0T3ODMb8BqlPv7gHeY1ZMdUFfCuEoff6+5rkaRNwlu2u78f
VLJ0oCakccT0R0szdTkdhMppDRZ1o23/S47RAl055/yRzuwPpkcgZs1o5jj9
z7+3RZiUjtazbBGE7IxuIA+BsZjiiokNBsUHG736QCAjobViKjyyF2CHz/iC
56nmoPIVq55Ck7ydby/MV8Yj53S1jufoGcPGwBqeEs0VKb6eqKW1Aqo0i3Nc
IvEy/VG8Wfyd78Yccnm6/uS8uM1NhHZtgXkX0X2Gu9tMYQXSevzKKNlJ5sqA
uaNgecuMsl29HYxeuq5y4J2/XcBIx5weXJrev4GqSjBXMJfEmGA+Xp5IXz4t
xqBzBbOi1FR0rMYJb2ef5pGHFca8v4c7UBGng2T/GVUQXKfIPb/pW6HQseEd
SdH4NsUAS95zoJ0SdSIZoWxiGK4rXqRJ3kyT7CzJ+7BxZXKQVIGHfyg5GsVB
4QL0RaoQuY43zryz6TYP6X1xzcrSj5Jzm+cK0WUe42wCrreIfEZuYLjaWA0p
5Jf13fFogxeoPHfVSkVlPsnV+UwUHPsBO6sSh6r/z+kdFmQVdueWmGO55Mls
LnaxQlKjU0YjZyNT+ppml5HLfQp843QYTljLBsfxldE+2l/AuCAAPxgNxv3b
d0NBFc6cTAiymKZnSV6/tkLdpqfHD5Cq1hUUx1fn+0g3G9U8YaGttAAGdjye
c+WAuLO4gbIXZBS94LgF1Cw1DOBGcNPjK0OrnIL3zyLyjl6zzPcPc1mtxQcs
ATwsB6Khl2oiQmKOYoLYCG95kPS2O1jwn1LDtz0lRhtN+yVlG0sEKVFT+LhG
qTTEsgd64UQ5YYQODTaqKsoVKk7H2JAP6sisRJA2boGnXmkAztxLlXe91PLz
16Ti/qzZwuIHCl7RxQPBc21mn7YUR32REEnQ2sfqIiJXNTkxEchorRmg7ri9
F8NVp+IOYPJWFz4By1l+zAFcvcKy6lz9PpiLg5ss+r9zKGIkmYmLuIxaXFIZ
JSpl38StAACQi77iFJL0uniUvM9OE8fn+McKoiXN2QGvwzc3ckmB4y51si01
qRVglYZeCCcGDlacKhfoMkFuqrU/1/gXTP1bYGvq7YGafHM3wkvQwkj6bfQm
pbAwG63Kld/R8nPj4oddpWmeTCI3wiu2rLG4Mt8ZKajyR9OmPJ4ZOEcuIMcQ
2MoSwPMg/IDy4P4m00X8JHFteu/oq4AXQaa8IXmRI2vWq4GScbYy4Q4pNgMm
pSYMKkVwmjt1rbSww33EYi7lq5wp3qk3NV7puqZdV+vO4cKsPToIGnlqpMXn
xygcmf0DRzKG7io1d7cviuVlKV37ykB85sOMJILPHBVhn7uRJBM+X+GFHzYl
csNdmrnkj+WMlri5p9CvUTCY6mh8Jb2e9tILZAP9FNv24yBVqEoIqpIjTCUe
LFaTn6qwKFvKRR5L1qrtUMjWRaHW13U6WDhwzz4EKrQtlkuxNgOeaMiXI/Ld
tDF3TWAS7gPj/d00HsapoZh9BXSu2hksBI6OUnppOsx0Xiicdlh2klU9DthQ
qecXqmnElO5YjVL0uGAFGPOud4jQvkTUAygnGdhSettuuqRbOd5Yt8+ipH1S
fI6OOsLVsqDZKUcDL2tSjgY0GmF422zqa51p+vLVyn1EIVIUiyHvZft8/MQ0
KiIrKdxAkJg5tDYX5cIvRsQSApguDZ0d8Vfx6pDK8EZQ2h0wVp4EoAoGvVwd
s5CNBkQWYt5F8pdvCyluEMlRzI2048LCmQihKpF1PnbvGzSTr3FjlH37QPNc
8riJJnnPBzs/+8UcADVfwmlfeXJkZnk91BmtcAjoqeHMe5mYJDBYeDCrc514
DH6a/+6lbPXgDxw2ZC3+GEFPByrVyeBgGAu2ZYcP4tfTngBXIfoJY2Kq19cW
/nBmc07JXXxduyeJIt8FB05Z6tAlnnuSOBY+l0Fw4U5lNRirFGDWmytS7A18
OViuihMa4DQubdWc5fXQJMXbRmLwyxokzILEWHwmMlDuVwANz2LJg1XDrqJl
mNb0y2EbMUw74eRlaVxxCR/BCTASSEzRjMyoa1+iCMDFzHnxtkQwHKJL8jt0
zevvjD8/pqz9ENZBAgF/R5wKivGweJA2wxflct7V0gCOHp7cJnz//14NqTGP
Y+qyRu1COUEhVMfYrNrHXlJrsvWTTz2eNYWwdnTDHQhzdpIoE4aLXxQTg4/2
WDsLFzj4P3Iz2/dIPGNL7Iyyshzt7XLAzg3yob5ontvoKB0MZAwkRJ5AvEw9
a9YtrsWTlUwWfQsfZ5Pu6XwxuTFmKtUnYSl8bhvlwQiXlaSLwV+jIm4sT2Rp
rBBGmmm6fLoVFZrW1Lr8JezyN7+AUu4khNHETtL4hDCXAL4Ex1lr0+ul4+VJ
z3MAbMwSbrqQ6DerADy0Anxu5ZB/B3zWZ0me+7PlydUjOvUXjbU3GG1mAQhv
e18f/5wjl8982JCmwzey19+saJaVmbQmkJRWnKn2cYcmssjgp8uTuihIVpsz
zsqBK5NL5jaZ17gQB0bc0ie/4jFGZ5C0SKnpDMgIW/lmWrae3JG6rGZo3AgB
QJ3hjkfQRXBFGxVwUFCk9ZxDoEl8y4SP6SA5aK3vbkVm9J3YdsgJ8hDGd2zS
UQD6sWSogdZdVkCennYucpszNMnFMHN7tOXe58Ln74vpOpBFxRuMZiFNFtNv
l7/DApjrtnN0HQ4jkOSECH2vWLpSPOl/YSgDl2oieNS9OTwZ9vAWEFCFTqTA
LlRo3WE+m+jbZhDi4o6EFTY70FVbQUxByqqi9JKkhMh7J/dFRobO4wEKo4bO
4zm5rTbwWZx2ux28gKOY9XEqfH8nFKRyxH2n1XE/LG9DKmXfZUg+nvvg3Jfl
yUS6R52g1A1A3C6ZUKsRlwoGNtKQciEV5l+RHX9ETM44fRh5LKVuXXuWU/Qe
bBsdv4SqFxo8iTUIqK0CFj2C5Qvd6oxmHg2QHtaHfoh/17y+wbsTYQmqEM0/
H3l6PrnTU9apK8D1shlZu1z0M4GlrdP9Ij1XZ3LCAnW0if0qTuyddIo3Hmo0
mqsaIDSf5lIpPebarjJhbIujdgloJD9iUSDqkiZ+bnkIBSqDDweKc2KuyR4r
VQ3jMRoo35T+x3ud5zzMovfYwXlJhBCi6sxay02zfViIOtgnPsSKt9wPxgkq
EBu0r+mt/c6NM6uys+iXQUvccKO+h9cCZkj6UiiwrdWnOakFz1LfbswHpU6b
TevazXfKoBm6/+cWCcTkltFOHRB8Fds4eyg36O5Ezu3IZfTCcsUWF3hGMbC/
v74pmaljiadndvA8+IDVNZNicoM4CC7LNis7LYQqlxOxnnU2OhHpoBT3BMUU
JlTfnzShwAiylI+SM3RCNH+yExU6JtiQ9E9dlI4K/DNkMTYGxTFR4Jky57ev
LfXSBtdFafF7QiTpaGJsDbhBFCwzQaEG9nC3lgBI45nDbn6uDC8+JxdQAm79
nH8oOhdRx8mShUNtB9pXERT1ximEkAqgZZm7lTn1HVHeU8TlQY7+EBsGR7w8
JgONjYyIy/wXlyPWnQziaJZxjgG3/nVqWz1NZByUP9QHuT0Ck7m9P58VxKSE
HRZPUTnQa/CyYFCgRb5qZLVsDMmGRhSnewc5qygWqXQBLjeUvHgdv10Dqd7t
oaBHpltQr+Pwy72+pLFk4L1So9Blh1DPcePuKeEH4gFUCx/eFipOlHqHYS7B
nyo46O94KZIGjdG/fpEr8uC0Fx4Vb0xs9IfVh36nfZWLaz4Sz6vB1U0BZ6Lg
tAwcFgCjLDw6F016nB0LXCAIv+vmkzjO/+sKPlQotGvvTFvqifhLGKZxBm3N
ba99QifktRTpVY1j5/xX9mlAyXU48YlcKqz/IB6nieTqPGQcwMKO7YP5izgy
wXiSa3JuT54rmSkOKjmen47CoX0uySgyOWngIMDtmbE5TKSir7Yt45QbRZWy
tQaxZFKYYCYqc6JIZDqezLR3T5qjoOR52KudaSUd6YM0dXZCMZ5NqF9AMbV+
Lf6RvrWuUx8LadQjxRib3gFH7kXanSKTpUZgwmtQEIIm6sYYEalhvEWizZ9E
ePuwDohmP5f4wTI5wv9L2tXqsIHQ8spdh1S4vqwfgKvUOAfvF0l0ceKpAVuw
QAsfpjh2tEh1Bg8P0iPx1vSDqgJ+uBPFOYX2Dr3ttnvaG0oDpT10ekMdlNeH
NWdy/dVXL4MlyQ1EbPPFvQNjJn9F2yIDJcG6wCn0E3SDzlzmYPKdweWtNe5N
n5ZoH41fr7nd3ZAbKMQlgioZgkxlb4aQ1Zub/lBvkxxneyyDdHtJXFRKO2k7
lDIzwkZcgWH/e6TXYwTOqNCpMTP+rhK+LGUi4PATbnowOi8eZ3IaTyf12S/B
iUjD0aY/qma7ugP8Akn6/iB+MGAkQXyFWifAOLGmHmK5a5oILb6HNMtHh78l
vt2OCW7TEf7NTUsLsP0bNg6egvKgzh1NyKpfF0uK9UCcj8Ber5nZeBhSnbXm
spWKM5sZNFLgIRn9cueEfKWZpLsWNHG1yJ2m+HHvlVrW1Qk7hAJHFTOOSlU0
JhfEpBcwptNNmBMLOylg8bALFfIWUTr7zNxBzEO0cKnrEdxsVnGZ59AFcnEQ
Sz6U2rp+wMOM23rJPOOm+UIem/K0cuXwX4MHtRwrj+FUk+6Kh+Qpb3Z5hTBy
S48JPoHan/eUWURQ5diHWyvfnY+H/nvdqtlYrV352fFZKHOxzel5YRK48LH4
F7ZaE2rkCVYOsudI/SA5g0F7yXXkaULTmn1ou6CEN4SnUS0fahLd0sutx4rX
Nh+qeqWZR5JCSh570X1bmiAWx2tS0V0MftUoFhN/cVgsDAH1ibk4lShYqzq4
Bme9ZfSfYksAwInLSBwArtmEeJmEK7ctrVIyNGk6lf/3rckltLYhIXnsRJYE
wPKSULYrGS5xkbg0YRp6R64QD29f/nJA/I4oUzBnPOHSP7Z8uKMiG8jx5ulG
ChD+7A+Zk3Zb4i0qkcdC0XsfiTZLMpbnlsThSi0LtuTGV5cQ9jHpRfDLlgH2
jt01Mm+kL3DChBoGG3kKpFG9NER5oYohovrV7grO4v+cMsa76RxR9USQc3Do
jvIYvnxNWsAwGjXsg4+499VnRV8hyngQ7OIAKKQI4UtBJyVnaTqe/YQWXO/K
DDzkS/4f6wa4QOFfjCIdZfBFAqlflrdfJ+4mqbvz/NGlbo2j5Pd2gYVGMxmS
LUGaRzMa/AihtTbl7C504oGJdezIrP8xJYlQrtRZ0LUtzcdkzCOS8JbcBAXq
JrhYV2kyuhNvQ3ipEOj/0ZKcK2h5vhNErsK/qOorkuO7f5BvSfEhuP794gWi
PJT71wBZa2CUp/uB9hLalvjUgvMn8BqN2z3jYP7AMJBiA5vaM2xh1afNjLh6
f7bNXxxbsymPImLFALlj9+sVz+NN9UmBb+yFMZnuj6TEkBAAsJa0c7K6EHMR
0i5adQp0H8rCnTrcrl1wpeTv2Oa118+DtKoa17sN5wpxuaYwgSgZttsrn/hN
Uri8TfH+nU3EfTN1/2he663SgNtY+r7ZNg3xyZyYsFltYhh7YI7IpJ3n4OJo
zhjaZbRknAX21RUpu1nU5GcyCHjX+oYd+BKWz4uTu2Nse7cUSCAJQZL9pg57
fGnJ8QM7nrXtS5ITNrDHCcTRxCqq2s7X/jz4DlXfRYlLElnBi3jtzeqLcqY2
3bwDP3BUKmzTHhvAYLiUV/IiJZkiVyCpVM/7rgQwUKDi6NakLEzoLVYMW90K
ypF3lL9pCnaaA353Xt4gfrc3HxvGiqg8GVDdZnVtgSKuXeNb8I1gnOGzEruZ
flQcEAUVCYXXNTG6PnwJK2e2y2cIFCpnIYCS4IFQW4v0y8c/jVhAplZrEMc7
oGRQOR0NkJKqtg/WJTM62WZFN89ggcPr0vH08H/gelbJLZ5EGB3xdymip52O
DSih7tUQTUPZmffPU5l+lXuNWp+YbJCfJ07ywJO10Qyv+zXUV4zNabJBQ+Kv
4bzirI9SVCFQBaPOhgezcHeVaenJbWJCMesDrY71JDj5xh5RrYZSl+7Wfi0r
qMX831fAXJadQmceQ00LHQWWdyj0fFHjwJEOq9aWAyDY8R4zlZ/rf4S3jUMx
IjNxry/eD1Dsmywqn+zqWs9GlZg+Yw1X/O0mzF4JvZUvWHJ4ikit6PmgAiX9
Xb/vBCPzowqDadD2L+Y2uqzKuiAYHhjBPEttk5EHQSbbV0QAV2nNmUNmF8WH
zwNB2SpwJUtWUkWqoypiQIC+9NP0XI3NTvh7PF13ZGrpH/5muHX86ZteCVXD
ocLW5WhXRBExbSaORiIIOBV0SauYNBgLPyJ6eZT2c22jH0T5rX698DzYj3gJ
QoB8prKdy0k/44KPL7mQ/qaB1X2XRdjENF+O/+KV9cT1k7CSU68jvG1W41AA
AcpzUTg909sacwotMWnnM7/jkxPaBviFV8huZ6AwJshNCTTSn4Op9lmcvyS9
bI53MNQc8pzB49aRUvxX7x6XbX3tHrR5H0tVQnhntY0+fYk23Q4x60axLtL5
gaHzbf8Ov+1bA5U4AvRVWxzKvFdWVnwrRwg1K3Al5jFUQrchLndwX5xI27sR
Lgt8bbnYNCfrFRntDJ8U3GmMkRBG4QcZENT3Pw8mMUipBW1GIIBwgmVBxJdu
4oXisk1AvjATrrnCEyZoWO52F4n/dlQFm/jee3Irt70+YVsrhUYATvFajT+8
1AL5H2aW/m7TOSdytOQ4yEUsIVCeYnDKxM00U4i37TceD9qR06P9ieAc4JLB
5JBInN3cbF+5nuN0QvhctU66OTow15+NM/Iqig83SYAvvvoJlV+b1wE4wQ+Q
GZXLemsPFLSn/nOslXPfUW1cMUTH5AdHeUXzI5RqMd8Ih2Cwro2VHQF/ZgXe
QoLXY2wghfMYROzGa/Z4vzbnyM6K9frOsVJiNfWeagXZ/yAhCPXcF4OOOf1I
IlhGhr4ckNh0c5MZoRpHM/k67c3k+I9rh7moQsIYuFpFdcwfvW1Ry/Swg7nL
AVrbqXm00BSFIksMV7NL/baYC/4/0YWRe75vORkHD0l3ebBwqZHwPNTcKo/a
0wZjOmmt0RgrIsQfADHm0wjNxCkpArxjou1XNMvzxKNiUqTxMivfGnnpQzQ/
XdMNocGCCapn69XWEjgbaLndAd2u0dxa5ItRjurSVudh5/F7TmYDeiJdYbTO
p2BeJ6jncKq9WCALVkMbfJfVv5zC6s76+3AC09mZgRhwIphrznJu/9Wi53VZ
NoRx3Dajl2/hSUtrujlKkqnILAWl+p0a0WcW9GNQHY9l4vvrQ2vt2J9045kn
6y+mZ02M/nf6yS52ua4KbVgMWA1QIiKw3ohK55vxJfJGEAcFhv1pGOlBhcFb
ctYAzW/yT0++ZUJW9YRT9L7RjE6FjOmcO9n7bs1B2BrRIUgaNAzvzcA7OlBp
LtEqTkcF0L6dw0zkEmDlayDX2yexALWv6SQTBeiKz1Mwd7SK9E+jTRcb5buE
sPiNCveybCJm/AQHHDock8DA6JBaoAFS6gHHliuNnhvIyBlmXyvQ08sKN2oE
EjsoicNnTTrd91fZyA0fIiA9wt4YEnHuiT4HyKYFlW/xbKkFMsxTdeJ7+YOE
QBcoWYpbrwoUOQ134hwYoaRIdVsW3OwM8UB09F1LXsqQd+S7CLPH3kgJ70Rb
qJNagJSVxCs3N3Wv3OuuLuoAx0RomKFXgqm5d2O/Kf1nSUhPD9o7z2I8Ia3e
jEIinjX99doz4GKuj/BdDxT2e8lqvHh18wJEx2WTG6U674ZLSai2K0SCVy1p
0l320ZZQ9CJuhmhH7nsGqDACY/uZLfvYf2G1s2uxa1A3ru/yiqggxdOliXRR
pJyv4S1J30TQwplmEicA6OBU5g39YhjZmR8Dplzk6aeGZgaN5Hbv6GnFQZpe
poT1KdGx/H2qSW2odVGLvRiHr09pGwuIsoS3ZsH1fFmTOMpbaNKbBrOneNs0
dc67uifsw4Km6FPJ1GXzBV69M9Dog71lpZ/CmlFAasKQilDNgNISez+0rdDT
qilBQFSliW2jJlQ9mNNi3rRLyP+SHor7tzjLiE6ibNqdkScSWRlcDIDXWBx6
tFp7bYuKyK2fssoI/jCFbmMui0uEZDNIxxyuWZBTZgj1aoRsO2GDmBIfk11H
HKLHp2E9zlFHZinPRBPfsiMbVYD6OxzUEDJeE+9wox+WSFIHa6W7VP/O7xCe
rw0AEbgB1rrU+P7pqO1VHJrQUGRaOKLzTtzWk0zcEktUIart1DXo2M0wHDnc
1UvCHxbaXvFCCx2nTAS7e9JxilvjK4fH5YU7JDhPjRPaKA1s1OEqwbYERQZx
QKuntVR7rlF9ha9H/ED0AEtb7bYe49AeWPRc44vBqL7oVKI/JMCgebs6h7Pm
8Mb/gF3aUjfpHyep58tKXsxx/1I0gWacXnuLQnGkNPxXHu/ojQTMap2Q0Is0
2RAiqLuXQ0uI6zKcGZE/sBn5kdIt+17ndwwAhEVy5froR0qMHhq7S16ala67
Vrr1FQKRTeXxMD5SuXJT3eyj/2FjjfzwlSnI7mBeABPbMzcNsswTw5NNjQCp
hwHTBNz0qRgHPaBS9GnWvMUFpbmbojQfQi/kg70P3RYvuRBVEl4GRlm2YWOx
JaOawMN1air2Xk+LtOy/KFgoTaAkxrf51TGjgqJDMZUHXN0TeF7rVtRLg3NN
x6AqBLSnadE4wQvOuGKtvdOALFUf6gh5ERflzeyitL4alEkf0vN/70KLmxMU
21s6npzpnivG2g9Feqflqaf2wmXcZ6juYEKqKaLeG1NVKopP4Dd61d0Fq7/b
NxgQfqwCi2klviV3Icg1Y8g2Dki3ciyayYQD+uY8P+23SB055P3HliC0O6kS
D9lSCmUWKmT+vE+aGKv+wmmpqGcZtVtNYp8wurjS4k9bUpToi27PGA4D0bCh
Qr+eEKUYlFjdGjyrL4wS1rEgocMh0f3PFo9DJYv93YtHRsUe4XfXOUs0Wqul
xqUHh/K41bwJZsqSRIG7apPej7dlocczyO4RK4jnJ21KWZh6WNwi8x+bux8u
YZbxBhahL6SunVmjOtgzE4Z/aTzB72Ecqvm0yhq0rVhO9VtPrvzZitYqCwG6
iWjTx+Bc/aPZBEIj6HpitpzDQftvcAr3bVy0SkifHjqMxjax2J3hsOvYxO6R
8jiIQwNDwRoPO/X1TQxVdcK3FWkxjANwwZ24pZdXwO4OTOgBBo746bU8+XnY
9IVXQG6zzk2n1PtwoZMKOztn46kAbnFhXOBOdPSzGxHJjBSD8XWyeb5PiTRv
quUuygyaqyCn8C0cabBkk+HS2LpOWsC5bVqHWQm0TWNl8XNVRTtEhUk8gIcb
p13m7J1uywRE+9CFs6pJn35mhyiqgq+NoVwBOgm4LeDyFNW6mEmjnvEPGhho
Zrx1gaXdPVn5UKnIi4AyJUtNk9qM8zYfhv9hsXv/KvVopWJGpEq65pJTXTGl
iVv8JqXxSwHuxHpSGkkl6U54gDQRNh6AQN+u4taOjxTfAM5JK/LYrOczT+1+
5KV21DXKDiR/g0DF+2BCy8NIpouvPnS5UtQqMFFKr1wBQCHDY7kZqpS+Pjja
lPKjCK9giLtZxH3qJGCOtN5tYRa5LLoHd6eeORQ39voaYIG3aXIOcJnWgTOt
nWQSHgMlj8/W+4bifA+9sjzd1g75N30jes17FQyHzZw5lXDCxhs8XqKgonrX
0yhhFCQ7kUJUlMcAL2QUqDhPlvwjOXw6txxcY1Lb/Wmvgb/LCTiXRFDPQ/w7
qmaZbzr1qVmAeqdt9qYlEEqm8oUofCFyHXEsQZBxLYAncQfoWw+QeDV5PIoX
YVaU97V29fa3ybkeRrNCUIbkmcKgx/q7HcfmktQbTrETTGddsXeZ7TmwirFH
HAtUxUSGnvRbdCh4mxnKhze9c87AoS7ixh9kaZfcXKqLFYxMJJRp3SJZp5HJ
tLbjb7kBsrF0pJ226UjPrj/jDHGxxmP0Qc3L67YVQ99l/o910ldOcz/Ps5af
JPe7fjxhpnwL+8rDDzG1aSAXgiYMi60cvdnj8ObIH6s+XiAkJiH50o7XxCSf
nEz+ZIw881ogOK/pABnKej1bT9I2bMwd4E225jJaKOCVRc2IzUN1GmW5Wjo0
YmyuXgadTtZ1Vm2WYt02JWtQphB8oR9zwvf48XRLAIXxuZWVW5ZSFwaGD64I
hVwsVIwKPBplgVeGxbl11MQVTg603w/UjoHL8ZcYkAFe/Qv1pL/jKf4Kip0V
rl8V3xrPwf65xfimioAiEl+mpbtFXC0iqUMbBGT9b2R/JiOpYx9sfJ5AcDKi
er4gOXPV1woRX0LF0Vp6dMZeuvT6VIYEETtoSkdkUWHUfHfZr2vPKjHZF2Wp
DhW6BY/NIi/jhmKEl23H7ZH+vPsUCuT583MfU9k0LREed/QCT051ljQ+mRVO
MVG/IDtePkDVkYZdqunF8ADKXDsKjGheNmjhNR4q4CIemsp8NAj+/nV+fTFl
/AlDcqZ97qGUOpQ+NnAG4l+o1B4HwwcYEfzUylBgW0+4lKFNd0O3vx/qy9wG
Bk3SHfx5J41vEKG/uC2jJ4gco0oI/RYGzXqmpFPOTE0bgtdHXCfUVFsplloC
YqWyHVx0v8US8ffaMpiNW3lvxNJsJEuOWTU0s86cR8ix4T1J1vsSp9OU3F5Z
y1jWW9+vEJttCZABrX/75/x/uLu/nHd3O7O0nBgRSdCe/fGxipWYfRkuDymJ
83Yrt0coRC77DtODlfjCsF57LZFNlPO9YDb3xNBQrdQ9iaAV7gEfqrMNGVn+
KgxhnYqJD9BBnndbHDq8u2G1vNix+LGiUvimmnSqCferL08dotvgNxIwdfht
kuIdEk7EFNeGGWn2RmI/YfAuz6H2hQn8q5wQ2s1jti6qjPMvAiJfpxneqREn
QfoRUs6poZm2SU7c6P5jGpu+XK04BWAwE2jrYXz3U/zb/fsvcN1ywW2975cy
2bo/XgkaA9jARpMkXaUo95GDhwKjHq1yZ98HBtda0f5hRxiJT78Y6OG41acX
JhpHON8YMVKw5BROESdZlyZBdGlWVa2ToB+5ph7TTRAe8ejSdu+6JUJUdrEW
lifjva2epDPZR1/g8wM9AiqNw3bfssHR8rCxvq8dAZLtihnxMqHV3KlVCmyD
7oI7rNlAArnZh2Nh6Xzee/wHint4LIkjce+W7IwWoVxCVtKgg52ePMcI4UB5
pirD/OZFb7UG5MKk/fvNO6J63ogX3HvvLCx/0Gp0b9f1dw0WAVSumVPgC+39
eZI0KPMj6gBt89PtWP0Wld5EEGz87hVZnRN9OhxSuGA1Ct3CE4RZEIGvd0Fh
g2iyXhQW97lGByFAqiMtnCmLWYaCjY4uS9YpjT3Z6PNxKmodzfNHz/Es59+H
jL7yi5tyNOqi2+61tJmphPQxZqxvcPi/DdWdpz/6H++8RRAXyaC5yQdyqLU4
R96r3ayY5TLVyyW+2qnhvbzbkELm8iR9OX+KfHFEvTTdAHG4qCt377iwi6Ya
zbfRW2qAXJMceF2yr+ts2WOqS9Jyy7BdoLAzS6caTpC27uVUT3Yh5G6XEMZ9
3Te/fxi3txlogucq+O0K8wFNEGE+ff3BEgn52H6KUgC7t5Nq7LBMk4pztpEw
zKQDBomdQKTR8U4mMBrTw0TXg2euOP03ZZ18f7H8Q9B/u/E4Mmu8WC7O/yR7
tRfPb2T86uJS8kUupH0y66je+IRDpWtPm9HOfuUs5IbHAWvfMaLvHLsyVleZ
mU9Nd8QdNyXTvzry4BOtbtwLd3/qJXA7wrPOYNxQuvfO04HguyU7Ysadi2zL
fn+TzIAQXjILDfFNEBk1+OINmezr9hgsWV6VXQUVbAHLXXkQ0O4lbfRl56us
jgkNunBuJTc238iOs6rpWEGZoSIeKsgwQjkKc9cEmLVYin4bAjt0yxZroy0x
DFR/5MyIXWsVRkyCr0Ep9Sx6aq0HMlUmjnEtwcjUYCWlAOhRux16xu6LvHQF
of7wjh5eufVbzHblvC5QDJXPh9HdU72tl5PsmPUuqKYwDkqFGsHxAK21Mc7B
jOqKjRBTVvtHT9ewGFzRX+yY/lIqhfxoJuZfd6gGj23kfMSJ8ijNXxATg5Hh
eO8nHnL+ODS5N6IQ6+iKrDMZPoSL3wsV1mKbvKE1s4dR/9O+yyVbQ9UqmJhb
u9dm3U3W47Ti/SmesdRcqWG7EKQ/8Q/WG9A2OazmC3/eEn3LI7tDRrwRC3oe
ozxE3fGulJhUYAHA2ax9JG3bNpu+KTHE3J3qfTQzN0y/FsDZQtwCspV12aOl
9PCPHAeod6V85FKBQUS09ExtkOn9n3gq7Prq30siKPPqmrS4aSkmSOmL3of5
/CM2RDZaZ8onqwWfFmWjClKufsHOdhpPL6NXbtHNH52L0N5J8oAFuHXMXTNQ
2HVBNAf9tNBGgmYsz6Cdtn1E9WPzfmpl2sXdF5hNUK2wtZEpZgdp0ABQSkPu
0hYbG6z6AbfuAHgSEafK1TEs1xy22PjOxMLZay1gxRNJ1Ar5+e128ING5drb
MM0kKRWtJUtBCXnjvreO6Gm7Osn3z8doql3OIfgrzNjRwJqgJwqFnCrrhtwW
OAa9BijNKixRpjmGhn1UbZX89gq22VfAYnipza8gI4MyyclAmUbPgpTpL7I0
fpA4expMEl6Yaxz6WW5/fgIHwVApLhgTFw9Zr3WnHZA7V826yMC8XR12YJjG
8Er3sZ0ERtS0q+OOq6IlOI/xSBBx7284UdhLzaUUQbplhvvKZ+goO7s+5RFY
7OcPsSJHU5T/P1VMCWHpIW4cRq/A7USzBgxZbg3Cw0M4HdF7tPtLXWxKzn+4
o8MxaKguklmj6Jmn8Wx5MSEN88exaAJEMl3RL4kYKuDOutsKdxRwGqhrfNBl
R9RlfzCM7yrHvXuMwlRVdZOCkDM4ZnM/t1aPwjoHRnmlLuukqw+dc7ZrmiRT
pifI151PAEG1YBLZtfUQtI0RvnIg2/q95n2/jJU9TxUp2rE+L40ITVSRZp2m
fr5144qkIgsD3iV7pqLN1wEtZ77miISwuyG00GlZXGW/lgiRKSMrcRZ7BG07
HJleU6Gs3NoQdEPdgYoO4TcPWYTKx6Fp7Qvr9XDPm2y6kidJ7X0ODSHUwntt
a+61PwFP0SS9rEhttzfvHtEI8YotCWwZQXjC7TkEJxJUYQBDv561I35pZ0bY
Wt9OuVApMhe+Wrl6f2rKD6WRtkXinfi7/aeneYzLLWN21bdOpurm4JKkAiJn
k4dCDQuTig6YHMH/7nq0wR1wCAm/It4ILU7kF5M9btSGFO5z8qWNdaQZYh8B
9Ot8CHIfra4XiXivU+nbcxp7aPd6gBW5oIsLDl/AIvAlQ9E1BFfTvyExHAB8
Ld2rPY4mt7ar6MaiXIx9X7C5cHo0iLRnW6l0zAaBbQdm9RamJh+hkqcGVz9I
jUARnMDSR0xfjxAfzfPvV2G2rSQ6voEOuG+mJonShOO6J34GdGM8D4YORNPI
SMhAY6MjLdzZ+VNVXXjcj2pXdrsDkjgIB26SLvfJe1tBq3xfJM4hyKmqfrCv
58qv1ILI5C6Pi3h65zGTgLdrcgi8oyntoHIu/WL1C+xqe4tnQk0Ox9hObjg/
bqBrlGHtHeeY7H05H+VrjW82vYEz3Tx1wEm0Y34T7rjJwF/uWcmr6Us+jjB3
P14equCjln1UcPdO442AgXfNFsCGLbgy9UZdlxrXfqWuDAlwdautln0HPYpr
iOgOMl15YI0cp8Jinz/TJumbJwrhngrFh6drFU/xHKG0RGVvxWW1q8F4w/J4
2GugLGzlH1plLauD+MSohKHC5bNbZOLB6mdljoDrxykDvMz84iQWlPhPxcsV
R3ajA9bG3DpR18dk7vAP1NApeS7WWl6shgUOCGlMh9mD36D2+u6em7AfPxqm
QuPjuxy+rrybJYgOhZfwyf5COLYgl550Q/RRxew7mRkcMcdP6BJoTAOZbCAn
+QkTmAeTICmlIM6iA8juaONCp5pVO8NzuNAv3PcgUaNb22JCB+xynz0vslCJ
GQAQDRHRdP0BhQlZr755d+DarHeStakcH1lsSb/xIeatRomCIsQyw2viuBlZ
zB07fZpR5qBMekSG1kQg2G2amPIXgpwU5yJ0BfI8ciE8yIXGXk2gIdSuntaD
3b+DIU1OiCq6E7Pyas+kHgdxByyvINp0ZM4JZXp9gnhA275/RmUrlfBuSopI
G7eDAHFPxxP6T2E4nqn3Kmuj1Va2ov900edujGRoNrpj0fOTuZVipSW0Uwsk
8W4jlQkAfRDkpaxLCPlqVPC0vmOOE0Grl7qWHy4PFupon6skVsgSsRWYqBBV
HbGm089B8OSggDeZVqV4qx0qOm0cJnoMIsfHIBshhFAMuLmbnWgLrg5nXNEV
93761QUocJ0Z0IfGvNgHtNcN2BQzmv082Ws+LE8iltBoLwaDcZ+l4ker7k/s
xjZ4LDKMKq/3NVP5yfvOOtJ10YQat3eQJVrWoIPL0AzIHQbzxnHFxx7JOKVq
GVDYQl5aD7r7b0MMDwqCHQ2qztmL897/p3NhBNoSiDOqbM4ayuAJrek8yS1d
YsPJng9GJmM8kOA931jNcjrjZu2b5CoCNlhYeeUOuy3VJkftf+xP4nH6v/xS
jsRWniQZsCch+K2qAGcyW/rlQNyC2U0EB6mLX0r5CT53bjL0trhbQXRUQb0O
r1Avoki6pNrseSB1UQbnS7C1r+b5WY6XvO4UTUnWy/8xbB6T8uvcBUrvTQAY
oXbvWs+PkfDvnc+nfoK/3r6ki79GSgInyqaXab1WWopHeelmCn1rywGGWfqH
anCIzFmtEynEd2Cl8TjypaBUzF10BxXQYAyQnnCNV0qMG2QKkI/MnCVUd0KZ
1XufeMypPgfQbF3+QXYXqk1L2XURt32PVBgCapoicpKaXVEcnSJ8aOg13rEd
G12zVxYOG1ADD4Kj1InWHvMqrjgIKtVUDUT22Ux7WUkVY/etQn9lUlhnYMzg
LLmw/iBijfQwRslP1q4msu+OXMfLtra0weDt6O8Kn5H1JIH5/FGgczTxaSQa
Jo8tQtpIj5ISOAOLa1ymqKrmyoqPLdwiJVBCs7uiU4QCWfHD/8+O79t7nCsb
gqm/ibvnlGBtVMZT4m5iWE3T6c5s/vZ8HsGV2DWJNHmI8xdEyVxYeka6UXrH
kcKwiKBRHHV/6A27NJaDzTgOKkwGSXv2cnoLqnNH2TYIeQS58qOuzy1hcErW
m7HkSY6Fhtg90ixn8urOxP42NThmmUC15C/4BqY4nddC2zZmirQ+y4XPI3ET
LgNTwmeWJeWcDE8o/ezagHMFBpJBD+4fPGUdVj2tXbregwyNU+MILIMhxODc
bqC2UgVQLIsCxE1pFT3Zhy2L36w2mju+1vMbSaCjPhJuHhqNubAp1abcRp++
veskYBdSZP/FxWA7KT7Bar+Vn2//T7oVyxrXGqljwcZdCHeVhXGiiQDOpS9v
crS4/Mr8AU4fU+qWt4MZTMEZg9JVs+Uk9uz9LMW2fJKmNQRk4UdHlD0Gs7IK
TH80WCwScr+RfA2EteBaOErMHaadq2KwyYFXpPfa25mcXX3+8Gl84XLtZlMa
6Wxg+PgiKlO6Xr0S645zCY6XLDbnR4f8fqCEDf4kBE5K9qpc9Sxxzgl4fN23
WYeyQOnoiPjc5fi8mOI7jm/hzFbpLF9kuX6OJ3DPOTsEf3DeylROiXaBnWVg
9EDadXM3wPtrHlTOF0GHLy4bLgEmj7Abv+VNPTz7woP/Xd0M+jQYZxodE8uD
13dllpaIMHc1LwmFMwnvLRp8J22ZSW5kMtbiyhddd+ylmeUI016ZCYyKdfAf
WanW6mmV+u8dyb21vCcI0QNpgaM2/ms53loPLssRmsD/e4ZABMHqranZj7VZ
VZySivYQNiV4S8pZD3jKf792VUqOY2LX9m8lkLbHHkLZi7X49qH02D2oW3yr
7nGWVjdHEKdiOfuinvvFFffmGSY+J6GhWyXguRqi4Uc9rmiM23k9GyaVy8Vx
96MJuz/Ph9YsjItjalntStZXHX519SrJbLqmvKU3b+2acLb2pnCSNj/FuB8F
fIWnvb3dmllUQxXKoawUROcFerF37gjmWT7Q9/k4Awi6d8NGBqn1HUoIs03B
aF6xI+56oSldJ6QNWYwvXzK7jz+CY6JxwTlC6ldo4Tb61T8OdYEsjVUzun0+
mxj9zxzS51cHi/ddKnxQZ/3YVeuRTLQLkD2XYLEaiP/eXzo0eSTc4PAFhPTC
WSUcU78lbD62A9Q9vU3wPqWTkPMaqntmAg84aYNY3bw/Bd/9zjIAuLR5zbXE
62+wwZl/B4iTBoeytGkvzCgfbGN33lImiQDmII/B9Kozg2zYzWkFsPX3Wne2
Eo0NZQNkWU0DuV/5u9Be2G21PhClX3XR6YxB1HtTZaBY0gG472F1RgO6XH0H
XjjAitu3S2R+b1mTXqo7AxC1IBRTlRJednW62IccTAGt0f4zT/uVnFKNM3Pb
duR5ZUe+Tabu8lDPsW8n9F7bIVI5SbL70KZOU3etFHNARjNFKmyAznK08QxA
QDpuc3StRvPVR72hJI9Rkn6JrLNsXzPvmEzUut1h2LA1MSR0pJp/QFRUhBwk
2Z4UpO88KmCMHWyQl9F5V+mZZs0ildv9V9KhQn6d1YXOtBhR7ZF3FeyqzcBC
tcqz1b9tnx6CxcpLkUoNMl9AeLvYQhfcihPo1P+oVYrw/OsonDfkwu38iLtK
g52moah1Fp0Z5Lx6RCPD/Bkz7KU1LKxvh8pMLOJwgIDQhkE8wBo26wzd1lzR
UzgN/KXHAihTn+G8c5/SV2IUa5MsOqW9OooE5iPdT5MKgBWOFn2YN1KloySB
u1XlCl1xOX0Y9w0mw+I3qePd81ChXRkWyTBlIOHR7buVEFEEmxAMInXMW1/M
sZ1+fNZRJxkvMympUd/Pt36vfcsijoij/I2L0Xpo+5ZqjAsgozEJVVw90z/+
vuQe2d2sXu/Z/gX4UCj9ixJI+u3QtnrMrTs3l4rPFoaEH0NxD1vW9b3KBq7P
/W7E0zVHIeoQbHSa3Gfa/czedqSjPW5TyIVcbSd35GY3HLNiyACqaWNGLIuE
VihjJzmZE+CsN/ageuj2LUcAFqfW2R40rhAzL+rbm/Mbhd7rsQA0esFvuolX
+K6qjCPtAmkttWuaWUT5E/GUWKOkqBbGCZ9t+nnk7bvqyXKKB09FOjGLDA9q
1VT9sLcyHGSjMyskR/zxYOrr2Tki7Sucqww0g2BatsBirCGm5GCjzp5apWJO
EgqERDGdtUPrvRaxAylfjPNM7v06uRuB/PBsOsEuONPFA4M/8u5URgGLT3vf
S4pUhQp02E1WfZO+FGbWBykvo7X7mk1GX9Evs/PY1PcnGzO22smerwvP/quC
qOsHh3yAUv7J+7XjMyeMdUWi25Pbvqds9pX6N6KzT8Y5XqbAab6muT05io9K
/bOHm6iY1QFwYtzeC8braMpuZGUoFAnlevGoaMZ0/ZVIkeIA7fLibkw8u2G2
8SLf1LTGAg7zG411VPy0EbNZAHWvQo6CpSWh65vgN4PCZvHotNVimg77tdo1
Bmc+0JnuMP5q6qd4xjAXE3Tk8HA1MSeMzJ9fYffjxrsglHgRhcZ8LtqnTbiq
dhUegtdNnMVGWmUvIl6cbLNkSio7aCGNEMNyXj8EubeHSeFNkkr3luyDyNRq
ZLLBrJVmsIgRk787VZF9DLRl3WG5eZ3qNoixG3UglXV1zD/pE5zid01/0+2A
xdJPxuduJ4e2gxBxgg+CUvKuzKZEXvYyiv362cuQ0Ld5kR3jaNxT/43R9r3a
Vw1GjL5cmYgIDRQd4jKMWbmEW/NwpmTTqomrHWiIwKHI97V6pftzDdGJ8UzB
YN4xyPacU0r+q8D93tQxO9QRd5J9XVlMyNdKfCPqgEmsfXZoEERdQz9wzbag
Jn03cScx9NKEUEvFJUXly/fYBGYKkdvbedQZbqUatuPuDYfxSmxA1YFmwbth
00nfJip3o7Ac53lJ21O1+ijkI27eIPESqzBwq9dRJJw+ptstuaYqdLueu0bI
fxxDD+sHPJan33KQjsMuxF5cuoGit8DDU6TkDupZgih/68Vhh8JherIDcMvO
zBLWZ5CHl2UeQPK1UywcvLcghgo+Nwjfb76bglzRnmBRanhsmgkkKqug29uj
PxkmkkrEJWO5yhgU7//rnBHU7ef1LjreUPMYXJWe6Z2vc92QPVMLAqj0pPsw
MPcPM9RYrH8d4LRYYVn1fzztm6Z/z56vP/wklcZvnZxfiLHgd+zp7mIfR9F2
rAlLDuUwFucjzkSAJ2foi2zgH0Yws152yxXq2I2FhlDZq20iEyCxbbmdAEZr
WTeIU+I0mztcUnzZOUlOYVLPLHEbkw96oHwzWaqBdAlqOhoU7iDpoOsQpNGl
d8Z1TMZf8rNqZiWz8+q4vFgemYY5e3qbjESkYJVZ1k8Ur3aLSd8h6p1nYI1O
6V9vAJVzEgOpuNSTuq/kBEenID1dLbZNa4vuUN3qTL8HZA+0nGm4Z+DKb3Gp
k52h9+xsy+P1qzpDeHbBdM9eDobZA7j60HoP6jH5o2f6NpvQWTgAUeaYt2Os
sL7eOdcKqbtBblqbbsp9f1lE4U7A7+VWHzQZRS7Ch5I9Zll5vC7tJBKFbqRx
HA69BDUUvJKvxsNlKzCj6cRm+zP1H447zajUBH/CEIYKTCDK1g4Qec9hN+nw
65vC6vle/0dd87ZzUv1/W+fDN+tuV8SMi0xLvDONYjrwwHlWZ90BeGWpHTlp
f7aw9xgM3PM8u3b/UoAeD9vee10l0X4ZXf01yw39wdMuUGIu9nOjbd4UNGbg
v0UJa2GiYPMrCwdY3n1dzmap9inGFLMo9rrQuTiCDsjFYdPkNtFLl8OVZF6R
xWz5Ye6N3pHl+/qq41k2YouDuX0TgxWV3wDlGoBLsmY1dqqZH+z7cg0AJdNd
yJjvz5ibixlEocM+ZlhZrUuZy9Mg80HpmMNYzWqxQz2QfLDWqyl7dVJvN/YU
rzgMgCmnyDyw6G7tTHwDwaalaZSN0FP5Ip5nAyuz/pJau42/vtAKX53P47tP
+R1kNHXJyJvIliqTdhZtiWilrVD3hp1zsDGYEK5hYh+73SMMrEQqAmVPu8dQ
a4Uqx8OHVjKrk+19Re6LP/cBLTsF+qGKpMyMDTe/sFWrlhbvN6+oBHPSbHaS
pOtEuPcHQva+GRKsyEDs+cGrCyOTniNi0yNi7/Qolaiw4zvN10auEQLRIILK
l3q8D6Ua/4dmw49BAr0zOlwU+CBVcW3YQN3MosLmcuERMMqS2IBFK+iQNii2
YQoR7J8sjv+Ozw+XAjvxb4IF2bH7SkplquCL+oJjDfD1GLk1/IRRM0hVnxPp
paU2KmOytsDTPH00mleqMUPrVOZap5J6YwVoxG4y5dsbC+1udyLN0CLoG66w
3e95jqecidcjTDPYiGSo/GEaReS6G7wBnHyj/AlaUIrYo0xCNxXgJf3Z7VHJ
SexQUHXC3mXCpq/v3w+j8qAk4VPD24o1f5slTt2rdDNvkiUI2NKVcUQF1bBI
whR0IX1V7pYTMufrk2bRBB6r0s1lvVN5AtJ7lmHAGgAT5utjASeC3hOo7n3R
OYUNSfUpYF1RvFqdmZrpdQ9U/Ze6oaUWWx/743ByjcrmlNz4sJmWc9LXRrWN
jMCQ2oLBLB2G0HiUp4Xao3m0cx4pg3LtCCVYCZfziYTSPOeEAfNDBpXyPkS0
PAvz+6jnrES3nwIzMQ98PHwLFsHkJXIG/kz4P5YyVgK/lDFplF8WXql30+YX
oKvGzndRsECrpEOg2M+1GClVO8tRBL6fVoQ1XGRfFzqmo3oyNNAJGRTXsSlB
1GajrhtTHxzdlW8nSD36OIoIUgAA07VUE+8Y1A41mBDSM5aim/9zivp9nZBK
EYJutsXoicrKhyJNIP4gGxocoR3z9atiC8d4fCV2SWXrc+rutz6CzRVPAjmG
BDJhjA9vf5CI5MW3nM4746Y4UxDXVuQ9DC8fZHWiLHG7bSWIXtHKoDmY7Pxl
wxEoBML56KJZBlRaS44AnitYx79RRjGNGgAYct5DDG1DQNq7ZD/bcNM9k2bo
30ayITi1oRyJGHXXAHVv6FvfXI6cP2uZ5+QQs7Yfn4kwcwJBzHoWaEqA0m/2
NsmilK2ihA2YL02WY1FaFEShYk8MNxZakP5PNI6Sd6QXdueue7nl/Tei5s0F
x8zp4EvrOlI8+YMJMUls/hI8HPb+l+Jmb80pUustHr9W4eXnXwRkfIzTvoD6
1O2d6H6Pc70ei7/BEFX3iPWe+XFegK3+AKDSMntmzPAHDP9kDMwQ816UZzCH
iQGylaPL0quAe760bh9mG7PoBUWFBp4DJuc12r9YwhN08jUX/g0f4rhOjuwX
qcmKeLx0p4jF6vGB5k8H+8rqz+loer9LkOnvz2tYm+Td7zQx44pH0dupNNGx
QJxEJOWSgvx42FlyckV9i9ESuTLoxIu0fbTWfhSfnBeDgBzoqmt/1jpPpcsM
yWjZyNG5BG3uSZ3eGLvYSX1aoczQWGn1ELBBMHMci+vTra3Zlu9DHhnAcc4P
C/1v1ieYzCCqvw0BDxvaTaj2XuOq3rBDcjDcUjoUCdvwrrbeCv5qBJJiTMep
JnEWplqmLyTmT5FlWH8oPjQprkN8b+4iT+amDmfamhCJiZ3hKibvyvdP9mix
X+vM226RjepGkRwd2FqcjTHamprb7uqNFyjyYdQ6IKFilt4pC95Pt1Gn73E1
u+b8JYdSZRY4VzK/9XR9AHYBm+ZbxsuWVXAPJQizPYF2g4vQbGjcB+Qxm7xa
w7/HV8M89UksjzdLPpkt4lC1BqWR+Pu+PBVsmfwKgBWVIGSkzf5aVwKxSAgV
GxawEaWHJDxaxk2KbljyScHzj4oAHXCdlUKMCodBnPurdjL51BVayj3aQG3C
NFAMHjv/4Se+eSY/x11IcNG/XND66JuZKAUfknnQ1AyKftzxxfd6X37/tQF7
D6Z1kn3trr/BoRr1UhHc4Ry3CfWB1Q0Hf4WchUqQSPdICXLRHWnIHvwANpS9
gtvkHgWKWQqXO9v68R6fxwJiqBD4OQGmpYXikUjJ4eZeEVepZBnGqgIgm3HS
8ZpQH7NmLJ2AUiBp7aINp9NkLBAvgRUbf7Jx0mvbUWwUqhwJdvx7bkxYCK1o
bb6KD5C+v4kNx3seUgUeXT2aUwTve/hzqsVzg6giiRjUcidilYbGTq4gsBbt
GuE77XS9wD0wi8z9RLHiX5rPEItHqUxzIisGdQ+DbLd4PKI4orPLA4w3S5yw
qn+GC/fLmynzR0xmIKDPH9+M22J+8RcN0rga1eta5Wg+GHmVKlkoQKQzfVkW
IBgpLQXL3i7Cxke0gknPp+7OPcOWPo7KW8vNtd5LykNffMTANm8jLRGnGwKE
/ngY4kM2g0bMf4mKbOy70kVqGBoAwwE1mUpYGljLeMUdexhc+jjuki7TK0Ks
Uu0YYYpUO/oxt+acic6Jb93hWgzpxc4+WUU+SWkzMb1/W+yvtDVIPJy268w7
MKOfaEBo1kHdc/SwWi0yhuj3sNQBZf4iJlLsknlnts2Ur8BZu1HczUja/uAl
UuvmiDOyxOzz32xexER1u3dAGsZRRh04GjlR1chlk3r4CcSj5X7iAFP3td0Z
3y5eNGs0Fp7uvipQVy0XHabLogMQIq9pskUpe0sF79KQe5wbqApuv4B+N8J7
6OsjEzrFKO2JnXdFsi5DwHhqxyjFGZqkhalgqdunGN21aPFVJSuCkDnWOWHe
qIY4DTgoax9YF9MoRXLExL9sdi/AMUens7FmPgdj6otTDWFy+G0j31pARK1r
ATJQlg/+GVybB7gpuw2Y703y5A+vIb4EgGbcPQAVFLkpnLsd8sFj13cnAa/l
ZLVyREOEK/t7g8bYKprQOvA0Q8BLglUdUVFyP1wuXfInmSKePlvEDqT+BydH
4zkb45mMSC0JQMyID3jt7tkqnttP/Y/clM1ir5/SyJYiqWpFuQLIaHaYmpd+
Y+unYnU6VY1KNmSVxgCKC1I+n8jI+DMtCo/GhDkg+HrKzy+zzI42dRxpbgB5
th5MUYk6i9jAVSr5O9X0Uly4NR2GcpCACrSX0JBvN8/Gj3Ln6A9yXQtrBc6i
r4R8Q1CYtQtxQK4R345ebWxBlTO4PqSGZVMHD9090RfFWYkhlU47D0k5zYg0
hJcv0T/o2KoCvFWWx3WxpC5HWwnghchH7cjSw0Ab5TtQedTho+vlWaOh0bVD
uCQeAiECmKtnhF6JZ9lKVObc74vjnQVEQw6ugF2VbBopJZe6inCiDnj9eZxn
FxLwCLOb6aVhwCfMDJ4/gk9n2qdE1FJKZlltso00BOlM31MTI+X1dwc9skDI
KJ7t5vN7W+G4C5Nv8rSH7jCXKvDTuklCFv5sRIlsJHN9JGBs2f9w7Mj7QhUb
Psls0jO3T6+8ls5P27e4GfrgPK2pnXCV5oLAY3uLrSmyHMnjVptZnlntI/gn
HLQswgmHhHBVCJ808D06SO35WwEnpmFxMO8NQON5a6ZLXNqcLCy5z3ax/iir
ceCHpod/UBhTV9nRkgtQ8sJFgIFYgTucIJLG73k+SFXo5dyzqiC1244xvkuS
792MQNvNSr5bSn3dqzyOlifH6VNBGcLt4X05FsxDYWTfrYS3Eyso9r1tjZo3
rHmCYxlAIaWGYyIzOH7aB6Jvr1A5kWrZVqt/cx05aB+K/Vh5dNe88kaoiiUS
LV58ZT5+AY7ogu/nIdsMcsogYePjv+CNzHUgaBuMGb+MaykbuCRBQ6A1icNV
i0edTEUrRS0LbiuqNWyNKZfhKT3or1wpYZ6h0HHP5NZiy9273Ch9DboKTTcx
4l48m4eaEHlZ0W0TOHrjGpl0kRc4V+dhNvxpRjMjO+olsIUY2RV60vFxAcst
Eoj2fWqFXkXMCHaktQ7zVguiL0BCx3JFjKlMHFqqUeRMUWbIETyBD4zU/UBi
NS83n+3vTPE+5yeLlWvNnMCNUBZxYtauAMguGfGJxr08oP/qhyVu2pv74j4a
qkLB8UMBda9vkw4lO0+Q3qcqKYrrpn4JhtviwbHu6uKvPjGmdqxbvOUIsJse
F1sAq/EVvScR7JsBByacwNaB3c7lWiSGO8bSTnLigBpj7b2c2P5ndiBFNFwO
RVTxUXMD4xYzWXn+dJddoPexH+4hUOMln5PM6bQqfzryjqbHaMdnqjdSxz/7
rdmNMyjYdr0BKl7ef9zX+2qm1UQkBNCaAB29IlxOruyRn4DjbQZoReNAFHfI
wRG2sLWqoVHccmuhvbr3b/kPA1PhNV5TpKL0eIuEIkd7B5oBEuUH5GAMw/B4
LjvT8X6aa3XykCMTG5IKTRwiuaEld7x7DiYrmjLkLQz5lRqIsoxn6JJriiqR
mGvOxYKrZGtBQUEYG4BZhJSk1CFkEcJgU7Se1aySImcg0WwVaNgRxPNkh29K
XqlnsI6yUpVxHobTak2zsPCLr2JsAKSE03WiPeIJTA7ALC7MF0amJcMiG7dQ
0RkCT03IXOvDOLxYQmx+uHna0RvTkrsuCTgWCWPdkLoTC5umvNQZhMIEAaCN
dzXJMOb1YKKZ8rEfzvx1Rd0BLf5ndmMKOVwfDBNgYdanIclVOLvQR6D3aF8f
FORfKicZWt8vAf90fsxi2A7T5QZRLa+7UHyIcke+CFG0oqxnECdDJqdNzHqm
QysdPzIxZkIf+sg2B+Zhp51unwLwvDQo7saOy+HWzb54Bf2TwQYqCLUy8el6
UUNsd7soX4AMMzufmOHqtSZYLaEngbHa5bNBf29SNQtYVGTlJQ5/4CpJmya5
CP4hgWCNJjM/db51DhHm1GXFiPI44XgL3Q7IzFD5k5FCHdptug0+dHahUw8H
rJ0G1CLjf6OOf04lblHdwI+BG08Ql5mVuvTkPKSjRkeMOLFmzxxb3AZ+7mZ2
YGCrqlStuQNOWsREOx4Rc89uPZ62dPB54YfKqENk/6tbDXAGP1NAQRlO9NYq
jLMtz1nNn4YEpTcF7om0vRXRxoph2TFzLRIQQN9A4TH9SXDxg6xmguqgfiMb
6gN1xRuKVHso1fLlxSce2AdeWapqgL6La3PVFRZ4iGuLUMa3OXCU8NAwCARX
p3pfGp6JQS/A5c0/kHGy/EC+Ir1qBvAGPjL0vYDATSF9PQzYA9sgGVNeOAvz
ApDqMmC93JjsMh5HWPfVHsUTcDz+K3JbQGp05sR80S5hA4z5G/BDogiEFKp7
rB0D7TLxJBpR0+8G+bNZ+uDctwHZ9OHWuBZdXKX9s+pHDnvkAUUUfVyidln5
oni2j1JJuv22L+dHRain3LhitSGB5eteDsb4qya1pE6nyfdEy8dicR1vplVP
Sh0w/sYY16YDzmZoky6gGJr+R9v/jO5tbXN9TD6UhSmdM8iLWh8dy80g50XV
sgnn7PjJgmY54gfyXz83NV+2hezYWPCkBErLbKHgTw62IH58yob8omYnQEkZ
Br71TnimEwfL+jwa5KXUav/egHUuAueWVSv1SujjJ6VOxNPj5/ES1p2rC+qb
WLHQCPZK1KlRE6IzOSTl2vYl/B6ZzA5tz593TG303rt9UjPW7wwRZLupaPV3
e9T9i7pu44EdOh/q2kYY2SlkpTIKnLBv1Rsg+Ine+NN6GCRn0FGcWF4A10Ys
n8l7GCqsjOUl3KONVaQ+rcQ6+wHOR2DWafk0Tp0I+7jz+uhWEbym6rmNrmVA
5urxoVJWTlRbNlP7mUPeEmA/mfsIlmo/HmiTbOUjAnbV5VL81O8gphs3jSbT
oDD/HXbWpvCa7niT5rclAAYAwTXX4NISyLWKlNuTqyfafcTgJRloM7X09A1O
qjy3xMiLWNNgontHL1/058W2cuFOEXxzK81G1fusD6C/Q8f+kBmnP0vsV4lR
hd8WbmKOXoNA9ijDpngi21MALlJwXURXVxwOSIUCi/4172AAxgUNcDtdyCh+
sFa/UKosHDTEXqwRcl5pwdTdzD6FV0Ij44OeGEOX5tSlzbUJ6TigVgfMMfvZ
3YGwtP0KLzAd+Eynehab0VkuMvvMCazwlVpIjoCak23KQjl1VhfBEsyuvr7b
izpQ4TQc+DPDRE9Tr85plxYTfvZpO6K6uMV1SrmImUi1OhsIGUcQYjrq8fTq
DezM8Dm697AhxEP/OOCIDB9bhtSVI6/hvlxAvm7jHXkUt9AUCWWs+0nwdN90
VpVLW7Pu4hx+12NRC4Pb4uIzOQcEBFZKGchIfBDN5Nnkq99vycKdj3XnJio5
J8D30l6hbGIGkIurce7EB0qQxAtqdrYaMAjDy6Jk1YiGzroSB1y6FjmCSo81
KRo+T4eNL9j+tLefDEYhRkb9df53mL2E80hCRIN7OzIEbmJXQVMyROLoi1Yo
WG94Kw96NN+Bs7M0cAF+CEFOeMHw794ZVJoBJ8HN86NOP85vrFbzhbDO1MVn
vj1GTFkSh2Svqh/v6FTvIG5pnxyzrsuOm3CqROW5P6UvuiPeYNaD0Sj3shiH
WAZRsaFbyVV1B2T2EaP6aYqGRImkOHeFnxPGUdsC2vIZ0QjcUbVGRXXwo1rB
e2/j88u09MSIQ5zlrSiuuGlmyKy1by43rM+NUJ+uBXy1uGWlhEKF8gKhqVYP
yJm7TzpLdLGav55b2aytHRmZYtj4qKxEI2BE1OU1M0NM2lQFR9zqqD5P8ts7
76FBWRYgtVJk5anRRArC8tyfaQQm6pgIVY5aKRMW3pjg3zyY+kf/erCNLkqj
lfgArjWIuo633g5EkU1z1ttll6565RomI0x3zkO31DoyPVJzi1TFlF9UayZc
nw2LovScv+WvbnPy7WiPdSfp73WCMgnd383ssDs/I9iqzS+e8B0X8O7tKWrK
XFPrKiF5V69UF4FBxkStZcV4AhC/Mh+fX1YN43W77OVsb7WoImVdmRNX4Q+Y
Co+jwkjyceklHux38cZC9cKplJSR6wtleMgt4Z5PnLVdiWU71W54rtvxyr49
l02WW1+WErs8eE+qRJsJfF9/mwucnf1E2YjkOZgJhjV9o54enFyFyMW77Wgs
COU/9nJxjrR8v3ktPEHcwS/vx4IcCfc0DDd+zifjIgcKQpRf8y8DuzEQv58U
LZCaH1rq8ZWq8bfumram+jJIYheGDxwZyKfEYSMXUY3HrgSE4nEA+W+S4Zlb
EI2iRInsWjpE3bgBElrL8Jp8+s6TxiKMuS/XIa7h9bF24kY5BLs6lq3W5tUG
FW5214NJjuPdJ9Fz7ljR0o3z4pA6kdzZOc+mQkqSDh02SL7NZC+2BlHIUL7D
eD8RdP9ej+mcuj11YZf2QqqReoePVCi987xzFHOGFu4d1etBjVt9CJ0fmJFj
Rbub1OxNfNA7x+0TdiwP9C18YzKzA5IOH8rUTP2EBnVjJfHfaHsUK7cCiNSA
bVbpMCrabgT1vIlouJVEymsFayycbr5dZUCPpiMlvHn3GlICr6rG0dLl68n0
lWT/IvKzydo70RxuSTM4c64X5kG8Z/xGUXISYwC+gy7hxwzYOaReTSYp1BcF
R/9yF9fTCoVxxYvJDsyV4xadLFNCIfm0LkCTcPIR26Oa3koCt/0wDoUTk1+s
B2Jm1GHL+PHSPGZgPoHAYr0TBSGJCM9FEjBCLr7DyskoAcMpI5246utKC+yp
FdrY3/11EYKvew6DPidNhQ0+asYXueUnXXTiJHCSjrZPiiMmUDnprhR8pyHL
U7qJpnYOAjmmiMKoOhkU2nblQGrzYhYOtqSkjG/da1cqA/MYgfa7PnHQ31gi
0L8mQGPpoopJaSk7X4Qvb3Fnvvh/Ajk9RDwrjxIFblnZOXzk+BvFDtKYwzcw
ONtGDwCYCVPRmPuF5JoRg9hU3lVsPC0FOBxn+zRvqjz+gK48yVi/H9SdKT4I
Od3bMSvupEZsus+CDl7xigEkMAkibl9mhaxymvyGt8/kApgVZPBYnx+CdvN7
oShsRl6KT53DfpE6CPHeUs2lbFU+gA/x8mu8BucPQ8ZPCsBRQ4AWmmNsEQj9
K4PhQAS9wNqa6A6iRHzqdIgU4IbwBQj6nNr4LkXo27FQhvJFgDifJECIuyrq
jMBZieU6Kx384XOsnWW6c3B8jf+JXb1Qgs8wOBF5IcnyBu+ybdAbQkI2v4rY
axGWOy/QQ3hFCUSKBUvaqnzKMkXFKtaqnTNthHpyL3ArEJMTcKiSvlMdaheg
phh+siHUfczw0SSDVGvm0gkDMtKlJHu+pfoNEENKodRhdfQMscWAlOooG+3E
J098jaeHKAON5QOKnEzO4w99ZCd03lKnEzagvT7yp3kUySHzQHYhXjvEbd99
CebRtlgF/Evd0ujUvjKu0p3noX320zNQUFY3vr7Jz8W9b21IWDoqyGYPdKel
u1dmjE3/FtkeeqSaTWBSuSro1eKO5giiOwm7aRXc8w+z39zE7M2DhmE4PfDl
w3ZG1vsFcrvBTt0OcCOMSdMkfQo+IU/ESaAvYrtsA6ZJ5Y0o2tFrcpL8DAqE
mbXjVFoUrrtpwvuV+w9UpKHEKNDvYzYZ6jzhzjkgYrhMw2WDv165fKsUZREy
No0nEGUxsaZonUaZOBxY7KKA/+snoZ9SYh2rIXUrLSwMPa1IeYWyxXhNNwrV
RP3xVIMYIcAdJEngOQIWSG0TxS0kOjmoV7RBHtB7FRuRhE6bbsP2TzVqecY5
xECsB88jyhIslCbQUpFJOlPEwLhtPk6OBQmZ5RdcPHd5o/XWpwejNK9Jovym
72dEwuCZZSiwHqp7aiMjBrmHyTQBmqqjGRGoxOijDbz3Frw/w8jHXlAomPLZ
+1fXeIArj1029Ik5yJxxeSEX/8YnaoqMhokV/6sEOPS8wvp9+l8kGX0kk3Q0
4fsGL3de+XsAP8Y0bu8FjFMrm7Be36DiWhHFdmXFjIhG7aGK7dHKYu9vEfYX
73AoxWLpusZBWz7tvQu/R0H+If3VjXbU/ODtXBIuW2JnO9GEQ0WjsedjtiMq
jeegdfhgQz/9XizxyxhIILwpjx5v5cTLAsnhxF4FuAj8vkasCSYSjE2ZKNn2
TxNtmt9r6IBrCzh2xDDm6lR8g7NacyA+asSITznzbUAvuJZPRGnhUK/MDnWg
JvrmHYjliPALNMYcV1qEAVCcJChUZnWH6l0lZlrOg2aCG7X8qdg5A2rGoiYH
tjkgwFSHOFgJSOCC90geE/Go2ZTeKRaCjvDpSxOZuDxII+yJYh5tjEqpYt3s
9M2jh0M8S2kImAaWKUaooqgG3VvP2NiEx+v7bVpHVuEAW23CdKxjBmfFrJRQ
bi2Oh46rhmHyGB0A6UGR2zTpsoNPfQlb+EN/PgysM9lHbETNpghlI98DV16R
Aivb1C0UgE1Zg7hcNXpL9xkZUy1rEbZvvwKbtKJIGfVOzGJh4GTO9igXLsqA
RYqGP4B4N+ksPQs4dd9RY0tCictDLThO0xUCru+f8rB7I8+0JsrJabQVdUjv
CrQTqygYzsJPdrIe4cdenNIg5Hf/pFrhj+rpLnyC2bxV7/k7bCGR34wsvKLy
kPhLY3yfqTBC/dHnjO1hZsNejE8Sz+B9u51vDKk63Z7rwC/oAPclxpNV/HtU
FUyyId0PNDgSUEZso+RQyjz7Ym1/XaXE0/dapMGAUzPxqkRGuRtGnR2NUOS5
p5YRcT36283BLIyVtWUxD/7V6HiXPsqiu+19U0cgnbjmtXdNJkPvMtp6h9z3
Ji6BgedGQnODGCJyGzf7eqfIm/789rrWwZoMzGXnhb9LEmq/40CPjlfflCb0
BEIe8sseMbD2iHvZMnZ9CZFpUYx1KRMwxeCAYlfNl7sU6MtZrdonaTriVL/k
gH4lRP1YTqfN0WUvbchdS7CenqGZDDUM1iLHmfre1Fizfq5ZYE63weAjGixy
scje0HerfLc270P9ct8a6HBorad3vLdNZUdh3F0fwviSSJFkkT+OA4KvhwnN
5wJfJxqQKb1y1tWPiRCUvr4U68qlAnYyRb2jX7OotX4Tn6E25veNMn6pSscD
uD/j9I8vk+jTvkl1IsApJR5/4s3pPDSthcZxkCnvYxORhbpqibcrM/o/yPZA
fDOhUhmQztjxsKeAt52S1xBQI8W13lLtKrh8es/MSr8vwZUnJHckWEBcqgo+
Z7JPjUmuuXMoeVXrNCJcTBIlCkskHalA2nyDE9fCYJZzFofWZPrVk64MncGg
W1eE1uUkeaRAyHMvGZyzwRYbOneRoRiULBTemrCrXX3SWvgcun83dyUzhDZU
g8Rk0t0yLfSuFVRKSMTLVJVt28Nu5R57Ljx/a1QcdIqve1XH6VCWXhaXHv41
Y9RH8en6DfTAypFjN4NT7BuKIOvzc927BHbLItFDsrUod9d/6Njv0TxjkLiZ
MEzYG8VvFKx7n9W/OZmnEz8t3DOAkxD/DONcuKFReYiHf6iFzWOksdG8cxXo
5/Vw1w83LLhZV9zw0djKnFKnD0qubeZPGxb9QXyfYBAT8SJw+Tty8naajBEg
2Qcteha+zWipdlTzSeUHcz2mLlvvyvDWMk7E0VAr6f2C4vydg6H7+ZTKvkxT
K5KCqox9qJVaHgpci0Zb6TnqLegy4I8HkSsJcUa/mSxfik8Fdsm6hikeZa93
QasPO3/9PlFTZsAOJHbdqA3OQc0RLdMvMN6qDmBPltuTDJKpvs1+bsIAKwy9
Ijuw0n1DnHb5eXeQx3h67c5czX8we92YrJXecsR0v82ysYe7aZDJrWCXjWuB
r3ryWlQ7VhM50ko6Co63N5ngZuvXIDFQdXSc+9/V6+7GTPyEylKugAt8fvcc
GpiT6qVNN1Q8afi+TyQSNIiTI2SpPAV0riItwHZRSwyg83wn8IHo/T7hgeI5
87UUrq3E8VTcnfS5Q3nifWBkCTWNBumqxpmqdy/qKiW+vBTWpwkRZkE+CGUq
z/DcAsc4Aqi5+RW5oOyvQBT+tboH2x+I2assL9iioOwAyQgq1lIi1pMLQHdm
cQmCD4wm4fdBNjCpTT7/YgUzJWJx6ykxDTSJ/5K0LtDBTT668EqKuI4ZClyS
ezHsgUPNZ4mS8nhFfKY6gwx6AenHoO6abm3rWEvMHziTbZay3RhZ3tCAVQrR
5Yd3o3q29u+rt5zTGv9OK4qGHMJJI1QNVv6sFUoi7SuxFa6vUSoQT0aQ84uN
LAV+j8DCYSj81lE154ZGjT823GMV9WwGZYqQL5vjLq5jDTaDTYaK5rHQfuCZ
f8z0YL9m6cokABj8ALLLHtiddZYeGWoTEGuVdMgFENtAOrH4Mc6nPQmeXnwq
S4laANZevlDTtml0jjrzM/tHwJTI/KsNQtZ2LgtfVNMfXxZiPqnfOo3tFmpV
K1/M7krt6KuWLGVpn7DMq+F7jWonv/KyBJWPCaZLr/VfTvkk8Oyx9OL6ztFb
ePz/6YCG5kVCh5HAjmx79GZAFfVXZZHrpGUcdFX8nmaflpby/x7F2ks7ICY6
LPYu3OcmnFX5pWGggyvUvlAcuczOZycqpUQc0Z4MvKO2aXImSBxgyipP6swb
uVIOjfkWw7XQGhFT8TrzEoF13SntIJSqv/PAiobbjNWYyUi4gzdX8tfc6owy
lVQz26hpeJlwU3a8MOWExM1kxDKV7OWxA1TNKtDP8xlsK4lgtRri5CSKDk+L
YrXMZMtbmWPuC7RU6sX+jvljSNNeJgtiE+c+n4H6Rlqu9cI2KV2H71BA9oUM
B0pC0UpGZ5hnblWLFkFuDZ2KEPSbWv1bFxkt/CrvFSqBpqR8rplmZqhSwRjt
SdiWNb+FBmbnFSPPnzZmR6pNYkkjSrQk6ulDVr13UdMugwiTzpLWe31Oh3go
MwAhwt5l/tFwPLGMSnRnF6T8D4zfCkcM8QXd7Qv4Ff6Y3U7mAiUYnpgiFDfj
hgBM335trJv4J0Ie6gJIkFCosqAgUV9HkR6NRNzCP48XH6brDsMjA8kj0S1u
01O1rmAowI1TWdQL3SKfklCKB4HRwYFt1tPV7png6SP8dcnKeRZZ0F42LH2g
FxK2hOdAjB5i8C/KCSUGSIXxOr8ce20V7oBHhw6kiUdZWyfTY/JwPAG2OL2U
tFMCCobU2zRvFeE7EdTrKcJzim6r8SpiPc3KDZuqt7m0eso52Paxf9SM7Evb
bWn7MF7Z8ZhLgoYX4w0M3srJrU9I6nTYCnpPQxLZtAtgv/pZp7i3J+9IMaRH
RXM70jNMJISV3HGgwlx7smuoDXwyLy9k9pGe8INBrpkybpOi7ZYAnQ6D84MZ
FBdRyqw6KXC29f1+uWhhfmGRz6JwWDA9TBBLdgxuJpWTiKwnWWOuXHSPLveW
IM84tCk/T532Xu/UwEnyco+Hk9h0MgAgRUTLfF8cmiyZuub0a6Hx/v/w4/W/
2af3IlQiCeeRrozAJL8xCKUJ9oe8DU5k/J6Jwnm56hwqLvIv+5/zKxE//3CW
Zhedz9ecs+6BYoBiDtVFZUGuycabfrQi05wE8HC7OI5isb+A086B5138TVMX
3ML/lNfsjTHvugDU4HVO110aRxuxTxFILKbwfTJPkiR7rCr/J+tT31T0mlXm
gk1Lkt6Djy7bZ9kEmRlByshP1ivf4FXE2825n/QzBYlyyNv71UUWy661NnxJ
t+MTfyPFJ4Cqg9IokHPpdcyrCZmJsC647AvmT/THGGtHjD1k0zAvtjG+ObUG
CwWZwMbjRZzwBvuU6u+b5R1OC4BzdzNTaWCN9BcuJIBkwuzR247nYcH+pTjV
heAojGawtAfmPth/zxYXKVe+KhWF0Tr6oi4Kq50ozB7J3H1gRhzse2yixNvi
VhqQXAT33lxFKf0ffN9Nqazs3GGJORzJYs9qWh5kM77J/SvfofFA+8EbCf1U
Rub1k6Z8gnCQu4wgpSOn9spkU1AsHXRLHS5FyxyOnCqsS1O5qSqLfpkVtl5t
GGNx2u3URNu+VeIkOR7W2OXAnjq7tLHLQo1n1eG6JHCjz5NfUY6WRRzhL1sz
w6OK0x4ak2Ns9qCze30X8ygkm3NH2C1wNXA3y6GpHAqC/RhNYH0+m/SYZPad
9EjaGDTH48tW8CO2Gz4PW9/LSNfY1O8LzdHIP9yLNRVuNygSMLT4EPkNNquQ
S/UBmQfQv2XwqFAEyPvVyaAxY9AAPXqFEWpEXVj5dTO1lCrNFFhiNlep6gxC
wCjdiqNkGG2hKqns4jcvJcNRuCvIq4s8QGxchslKDVfHs6Q6DGKmxL9uVmFz
piX2MYEB+Xzn7m699FVWNPYgyp/LiKbSm/9IOQ0bRs6xdHsxCYojJ5yuxRR/
CZ8nQ6hCQ0FgXynj4wvhUiShcnaVEQWxc8DcFfGzjldV+cyUorcDolUFYbdN
wD2txd4jlic4iPJeZSBFvoTgSl7fVo9Z5QK4fek9PyIqPO0Yhnur3k7hoA4l
/YkrTaBXY24Msfy5w5Zpj1B5eEfpg96ignE3aT9+iwa1dhlTnoiKYD3lWFvY
1hf9UbThwVFOUDXB7a85etYEp/XZ6E3aJg5BzNm+v0tyT4BBQyTxJMrXuJcM
OI8/20ZtpIN+TW2fDeoWQIpvI26JvrT0y3aOZzaWKV/qvIbYv+rejmVpAt+e
rr3PYVEededC3+yj6je9ddVtSN900EYClIaiMQv1X4KYok3A7fRAjBmuUxuk
c11RXrZxhzNRKaUoaHGPeg6ttFQgwafTP9JvEYMr5fucUPkH18h/sn7kwAGh
vhb7fuQaDnQhyYvAe2Js3T+qubDXm41DXZKQK99Vir7XY/1M7+oMn1X3x/pM
D/skTyA4e2or6Ha8NJ/UiJJbAbfnSSnk4XehxDWG5Du78ch0S3gZFhC+Op3x
6YOuuJuCX822TLM2COOPg7mMQINp3esgZcyvwAwbfnqRHErk/e4DcYgLRTPM
nhmj6um94VNLjg4+cElOBWnO/fBKp5bqkJbQzgMcYlJlI6a+2L8ayM6N1Gtl
qUbU28Zhwmd3lPHm4xYtyLWPkwP9NA6lZZx68Q5ssCR1IJechTeFyntGHEaZ
ssNNGRjRD6slK8HgqW+r+GQ2N0krytBDkapH2L/z1sE//Oa3ZODCvx/agbX6
bPHmWHJP1qmCZnPmQl09wiYScn+dkmVL7wnCt0PqKXVHbFX0y9l2xJymUEYe
Jpb6obH/8/b63mmztK3hmPK+Fa3A3D56DkU7/K1//5bSrJmomr3dIWliMk8C
/c/WQtJHwjIY3BrCbqX0NDQ1R0q0UEm+/eo4an5fG2ZGlm/lBJMLdrOCytdR
fU+oRwmgsLEayzq+RJuHfJteZsVLcNSMKL3ad7cMyMukwOcF+g31fSWQ0jah
aZPwX3rE0h95hjYf+uMa4nyx3nLrDNcU0aLc7GEkpIahyQnQMV/dX9Yt1Pn1
P6brHet7hQlQOHPk+rTwz9gBZOJdF28jO8E0qc7MKOa7boamiTjp3S2jQ/VB
XPMvcSXqQceFS64vKKbuIyQTWxMZczlmZz5wygobrWzCqpx0dWxz+oe/0Lv/
mjuWVpISFnMBP8k9r7pwTfz5PBTvBszf1d9gWSvHO4PW5yWLaE/rvEguEwOw
+H3osLA8gl345WpaRXYDVYCph0uRQmQr8YqMFMc+chnMQhsVDO+cJ5iEdGHG
dV2Tkl2f8zuXZH5AgvZ8mlNF5U/KcysX8p0m42UlU/j5RchoUHdW0k4A1xil
xyGwqqsv9XY4oNVPda5DLo8M431Yo/E/860qWUvhL8yHVWsaRvMTOkxiXV+c
1ku0Td0XHjg6crlYVuEpALgmc4UVljP2D3YGGC1y7Wy8vpZ65xtvC6AYqwQT
MF2afW3iTcM0UBJfxpDrOxGu+SeS7n2ZU/gpG7jrWIKInQMjpzVyvfpbpSSD
c1HDDF8bvFPbCFTo8KhE+7bFupGvGBfae6xYIf7padb7nIFp2Io+t3GO2WTK
nlNCW2s2cFV6EAwzr8PGNUUyluDUM2v352ezSuEnCgr7KuVbp53jac0H1AVc
eFE24yzLowYrApZmT7wg3Bvamg2PXECgG3WOGj04QXi+iYfYZtThBaK9i0nl
gP8vX2tG6K9LwzhzzBiqOtzVBzennnvOibGaZxxW7SeUb6PICnWkXNASGdxP
bmNFfnN1B0Bt6XQ+2QnotdAoiQq92dJA4dkv13lGC8XA68bLaeqBTaggSlgL
cnnRkJDHqyWpWUic3sNfe/vgengqrpmrXYjBEz0G/RhMoD+wwC9zcFBqcShm
PjmSZONTqm6fFF3lOflQYmYDEyOX3U3qjT8iZMe+pWHbMM42kqNMHq59V8y4
bqeV1jvwQ27ZKvBsafZC/FWekXDiHXYcllvpAIy7L9FM6Hvk5yZ0svJqeQim
OHAgHvxUeE5A9NTFuRZymn9Jm6czKfPcmvKqURw6vcPqerPK6wFna/u3ZAzF
eZ63KZ1lJWH9XpmdSHv2qTwL3xt/F9QT4kHeQggorupSkxhPJ7BIdX4c98kh
ZY6ZW5gWI4gbh8bsj3o3gfpBn6IGdHRTPd1mbDSfkY0x1r29IHJjWz+t3aTr
xmy4m2xaF+75gTDs+wNByHHS8qFes70JJFNTnTYxaYNePfaICfdz38RZ+55z
WDsg2skYZGRkTMBdUEUZ45wL+TKdrHf+Q22zl0+X5NiyucPr085zHTw9FDPn
XV+4NknaVOFj4gz0/mUJUvswx8F/KdawSsw/oojMJPZ6FKuBD8VUVnX6dbJ8
OVz+CNYNtZClKZvowTaFH+jNlPNBBacXmxI4bxAklmTUDBprWbycRXckVqGf
03Js0hRR4FrVULu3RAsxjKE8pAi42nE/eilMfuvYlBzZmljPcC3pgPaMjk9I
DIeqzp3jfBo6okdRecA3VMjN730IafDs6QkLzNNzTE9hpBcMDyT8gwoVEq6G
ZUmiq4i88ZZms1aKLjxBvUIxRO/IS3F6aqREvkDv59KHQ4mmY8Jbl36yGCWi
6++A2AxrYPqVGXYg0b97hh73pEH1fOGbGSx3/xCmSe0Z6r3T7y3Y/buW08Bv
Yc2JQZXBQIbW7jzVzTtqPwke3YPuk+oqeVb2d9nvsvHNTxaMTGR+AxF9AVyH
naI61GMrB59XWlCFsmJYUftvY1YjYLgoCCTa/NEmGFN9PNpk2c0ZKTARfYh7
9vssPi04c1CCwPJ7k1wCQjTP4pzihEj/X9DoZ6l7z4c/Z+BBvP+lYDSneP+D
agpJieziuTn3d5J8NGMOknwO3iRex5s8ryOOPXeiD+6wuTULX2gqWIXB7Ks2
vsC70zXgwU72xVS1NP0/cXmE66OweD1AZWYauJHnSTlVZkFH23suCf0hkjnR
8iftJEOUTwILVsIF38mA2ukeuk4+ThWAAgpxe0d8G4xXtNfioV3+Ev+9JPTl
E4lLN9f/Rm6tdycgqH7SMrAA3gBA9STgNZ6nBPfuC0ab7NWA0APlOZu9+LAh
wWZ0heHy6FHGjap4FRGE1V++EngQrTYZqVrpZ62QE6pu+AU7fjYsWNsLgPZk
5LBqmoKBxNdXeSquD5u4zWVo/doDsn8/zBlQW8QCTWVbyDZQunnBQgZ3Jyty
BhEJheRi1wnMAvBUjQTk7mZ9OGQSLy/zowaAXRqoc7sBDp870U/+i4+5pkX6
odDNFd6N2b3g68V9IKwBhXCrJ/W/dHN37tKAXnp90xmnSJh2NUZ9Xj2Rxj/8
J313npL/uo7RRO07NM7YetPIvU2ZIfUi12m4bNThbJG/MHlAf0zsW6d8mIMm
IO8xqfFmHtrkyHPIKv8R6gvH0BKp1HIHLY9mekpaUN9GtA1pOsRL1bjJcHRF
bQ2fXHwIfpXbTtTsx12kP5ajz57hHrkLIXQgYDxGbxWmxFReQlWmEp/ja7rk
0/XRcowblP3siwb5IVPckRKArn0Ev+iewpVDmCpG7L2202bEJgdov4XiUA/A
9lEgZdn96eauXHHmxF6q5+b6EnZqbqLaN1tW3F1FBaxvjQt/HNZOIANDhy2S
MdOCJ13GFVWybqnhjhzw++OChK+wUvl7hzHUl1oAyFqxdPQ0pc/m166Yl9SN
zMEQaQFAvUWfThSWM0URtFw3g4Y5wnHDmeVj0fEoxetlB2n3a0Tk/GyqgFUU
rffZKuLbjo+/F65GBwqMGubSE12TLZLpfu+gosNLQ38a/maozuBLsjGtkBqS
b7YAUsSnYXmrJ8kXXVryYwQwCD6bKhQPlDwiomBXEvODQ07Z2Q1w1Gh/en4n
UyPxmZCkAZl3AfHPQ/jVPvX0XbTM7m49Lim2UPmPtDGqZ2Tb8aesP1TxphlF
3bvhm7HLDI+x8+WhO91xYeO07HpojR244n30QTnrFq3x3/Z2VI7/sND1FOxC
4C0dPDxxAt+7QNxDXwHW2z4nf010fZffAMrshipHDX+1BKvSCTCvj+Fuy57M
uGkfCAi4WIAho5YUcjH9qpIdW/D9o8AqyPiRAl+kzx6KBqJ7bO2DDGN9wCJ7
/Y2ELzt35XMFV6i2h44/u6AiDO0IqTdbJbvOyRDWHtJCZtsZAAb8LIPmEMwP
8aSOniDztNd2ebcan+KtoIOqnuZ+DWhn7fiJrVzea0whXYCZ1DgMk567mik7
CjIk84Gq7s2tSrsHLLm0ou/mBwi5h3p/0nUUQ7CvSM9o1cddqNR2Lov1TSKH
IrI0jhEW5+zsLl7ciKkKcm8cfhhvt0hdnDqCsn0JcaTzsrtauU5k49qdcRnj
aJqvHPGBnTsNGtSEfVtcSGxRiiZaFCUlxvaUmSYLwClTg6v5XkkW2zdekLd0
vZ4XFXY+mDA0JZ7Ba8kn8eqv2mnd/ik6gANND6r93ihrAf/G0QDywBE8E1sg
/V6Ew1oibT7MfadjBTawZ3kz3EfOzgkD7BkHDU1HhzeJ/CGn1MgcBhUGTwl5
w1TFi4sc4gTcWchI3z38rYMpfD1PqBQCeJU+8UisXtcZ2IG2eu9qhhULM03N
fkTZPIwYEK92XHaz6DZsKpXp+XzzyL28qw3CGj7Gxi+vUjlAlfZN0bDDINgv
LFSIh97TIEYROa0sH4iUgDaglG3ctIy4TG+4CA3FJME1Pd7TTwuA9Ib3Wo9G
5nnPfHxxG6t90lleYOO5pGbZRD0bfe6Fnfw7j+0U0mKFFktcnBmj/cQTbhJJ
GpUIYgaEdkfsTlENk2RgruB33WU1Eb5weoRSaG6dAxXQ45QRTxwpA7CANOtq
uqRwlUKEhDB4RnstUCuGxLIXDxfTF4Q+63bYy6puYViYaLMIJbZc0vvvcgpu
j2JoF2RlAZuBV2Eusz6N4XzCujxExohN/kgdt/wtzZZrtNDRZnPhhWEX5FnF
DXyyOLOEvx9dzxNzctiL1BgHGYFXy+zoObkxt3xC6EnKr+BRrDohGOZAezKA
3HDI2PmKCBYMnI8GmnnHUba1FK0uEggZsmhwhC5veY9tQ4Oz8azQxdozICgZ
w7KpkHeWsDHi3mnv8dorli0w8wrvKrZGDVhmKwirQYW9CI4dJZ/2l3V33Mdo
o8PGz1a1MP4tIvSEIeqbXt/Tb8Q9SGs9csd3143PqKKS2MEhMYjBacJWNubC
fSYu+/CSas12MbZYucGW6NgjIsOJqREpTHOK3IA4mMIwmrw+2XudVDyuykKr
HGOZhlq61wozsn4N5pbu/TSsJyOGDSU/sD5R657gJuwzBWGM/gKZy7YgoePk
AZaJMtGAaJR87GiByEg/vbwrrPdYG4YrvWiUJZYB2Ros7nUFacNBPeCBlTLW
XWTR/s9RlOyvCYpGdPltPQuggbrgZu1+IMlOJNJ8BMA4sGqWpjgMUag4HLxE
lbjWAjsU9Q4hIPBq6zp4T2+nATrE0A2BxDlzlAnBWsnQkXNNh49GMmRJomjh
xKx4CFemrYmMp93XeaEHnnf6jB5EJVtpF4VaFGCcZpmHPiNVjy5BWI71Zy9T
144RC6K05KsWGdPPBnBssUL97r5wudyZyWVVloiMsjLaGtyjPNblbE42n+jl
IASmsZJqDDjmsJGy1OWkpp3nP/6Pal2sR9wWGhreB96R1ELs9Oh3Ou3pB1XS
p4NO9w+PeR31//a5rnmEy3Z9TKRVnLVizzx56DFjiGNR/Iik/mkusdBgT2Fb
F0TxKsePbVJgIaZsNkoc2G0aJwSa9e1YbO0uv8m9ZtlBYO73LA4Vq+oIl53i
ZP8KOk8+qMZIa2J496isyGnnrtRZxtO93O+LSODfkNKKFZ6xyVUgrPjdMmn6
3GRKWdcb1msH45Ehiqx+CGbkUtYDxBPe9xe/PakDlv5PwsW3jNJuVh+tLMO1
g6sQAA55u+Xw29kzWTl8xZf2sXgl1VJfN4zBOy8hDWc/jOmB1WDaQYau/RL5
qLWCmFR+5lK9+pucc74CzLa9GIiI6dUM+twH/A0c7l8fJ3i16ZUueMdKxxGt
5Mankyzt7Vo7f8wqrAJe2le5S6hWBZOM927HO3ANn2N2+L86TusE0GCVlQaX
2K9N2I4D104XscSxUDMMI207ENLxOePFe8vzpZr6O5tZwkBFuWw92V7hqpLy
E/1tGCV4NR/BFqabtvvFDfdZ8d89tQl3ar/6Fu/I9s1Ko06PP/bjBh2DefVH
r/G6oDiwgB4q3aA7wl3YdRJFw+Ff4yks/FazuJU8/WIZCkKUNtohqtrsrCeL
N1Ug/9LutgmRWAv0qc6VXrpO/YUdhgyQUMu1d9RdgAqXA5m89bTopIwT/iVW
fDrsFCuxoH1PMFjtE/6V0qQtV8bkihCWBEP9u4aLxoM/eUdqqyjYJBaTrkRq
CsAHVwVKBMl2OoV2xIkS9EErYMOF5sijREwjVbynjhbJhi5mEG5GmVmRIBCu
rCHw7t2zIoz7GSX265urj4ssNt5qi9wEn3NZXCT34E2PtcCp2CWjHIkXuSud
C9RLf62JMwBJY7sem0zSkz1LOT/3CL+88xUDWS25Ktp+N+4By8vLbkEhNvGs
AkhCoFzwIL3nxVUw3gdRHaMTq/bS5zi8AwugNCZAqPCjLxJvRvsvpJMNHELL
eGdQvCkN5tRheCK3kApSElkHGV3WO2OqYoSMDHYl3I1/0csEGAJqlz8e4gSo
S5DFOzIz98ebnrDKuU8nWH9Lf3T1g+6cTT7/ncfiwpZaV6NAEG43HrN/W2j5
KFziHHDTV4Eog5BBluww9JBYxNRbxykodnMkeI9DZlzMZFgKhqKnTJHOo4rU
z8043SgpzFt14nKegueJ8jqs9lM7hz7bV6wlZbRJKEAv/G+RcOa7t6ZDHt/U
TpodSeGtyA1D9PSD4cYaUsoIqOcZ72evOomD28AS5U6sMnnPCpX1zMr+7Z9/
WGICoX2r6Ca+WVLdEAyS0pwGXEFwJIo2mB1Z964V//jJDHiKLMeqnedoPLKY
aD653qcGJAdgf+xHbzoNccaJkZ/1dYT89nYCUa6Ad5JNbH5+brHzqhcWwIts
jwV637rbrW98x6vRYdLOyr8wDzDw31vAcSLIxhXU2j8CMrMABLYprOIsueBs
4TLBOCUe/cwBnDuoNBzzWvxWtYM/BBp12NLmNtL50VX8q3JHNTu2svrX1oT3
gB1xuyGtJLvYXiMN4lx5G2KxfCL1urzjXST5r13gosJyDAa0vd+Jo1+P3ixX
MyLDyonvFYT52FWH6TJGb+UkoJEtJumwad16iDJQRHgXCUqXz5EhVHqVzSBZ
0okWUEy4dRJndF5I5jNeabg6ey0i2/1mdqzWLcDrL4agfS2tn0W+YZkDPZCJ
XK0ii/y351KO+hDZgYz+ORi+zZStydFQvm3s/oLwlbK1dSSRnY521LQ0qEBK
ivokNskmWclapJchvPWVMv4nYvBzjnLUmZDKOC75BuVvkRrz01Tw5aDAtAfQ
g84MFfh9SZGZ0JOIC/+/WOrUoxGff/dLVm4+uPQW/XIRL5LQN7HNB01B1aHD
SVW+GQYoLd8fJw3og/QrjsddZT/I5sWnV4PQahJtK+Rm8h70/PdTaxieCrae
WW/uozEp96eTA+IxQjIwv0K+Q+qJ+3P4aqLvOSmkv1MywTHY4p780ACKa5e0
2X+ssBN9X6I0ITuARIvWzMKHROaVa1ZLpTxOW0GuZM480epfDrmZtM2BTZdE
KzRijTGl6eXwTxmDcKNtJ2EMREC9aoT1vtWoWfYHN2Gj4kzcOi34OLDkDEy3
FrzpWNBnaySu/vY4J8jrS6in9TzSwtwBCpsy+eNWmkBJisYbJVZsVC+zQd2B
NwhZmCjD+GeWYdTmb2JuPbnPJG2Qc/uPrtUjNMDLMv6Nr1rNdUrvZ7n+UYPr
eN6iMyS2XlXwcndxbq5x0LKNCpLNGNOODy0CQNDwSj3BymnktIl8aTZOd8dy
j0P1T71z8OLwnnuTNNy2Sy5LbA62bish05wisGOmXgQxDsG9YI3j4EaA59sN
bbVapmuQp8g8o7A7lpP9qEzFwvH2sggNLXP9sG138SFU1BcY6xsWC8vymF/c
sz6luG1o4eyUkuzvLYOt8suUzo6QQK+VpUMakl36yxLE5n3nJVTy1kMkxfRq
4Wsi3kGvBFrbniQb+Bj5hBkAq/DBtdZwxe9pJfkoKcSVYK5Dhbh8fmKNrYgw
IAIJ4ICbvBN5cqGSyO3PmGce+0JB7vpB3nqyGS9vhZxcbascJtmSXfb+gXIk
3jL8F+9s3QKEGlGWOzVyhjlf5ZBEOQt4b+Jw9Te47AWG0iG8BjDpCPnT/aI7
NJLCmqrGamIhZqt5LyXmn/4iHIYkxqVyP21At7JPnGrdiRZndUakKgZyNdyZ
//fpFTzCCsVoNJxe20qYOv9jjIIpzv2Bn9NUNncSSKmDXjYy+dm8IfvsTrwk
vrkHBK/n1iOAdDQQTWr08z+0TsHchwL0Cenkn9W5NremU4j+smCasJZk8d/z
ejmjQc/cKcdxHl0yhGgljJcy7DwcgTDBzvX/y3ARXu6tgqjSMv8xPEtLpyrW
x1gYA8WhffqM7ZzAX0lwwpzY+cO9I9IkmvmJFpwrz5P4bsY51f6sPcgqgZbG
HHNEoKpKEkFnp51kr75GrbEiHX9mQQm76JNwuFtgPkvirZ5d6/ILLGPnnc4R
5tndBYSF40Mn2SZNnRqnWp3EuLLcRD6pnp8+czfwPrNTK9SuRx2uZJU2UgU2
qdaj9n37Iv/oVPyhXSjnfTgtI/5Wd4pqe+cNejk2ExFLHfJPbNpFqEvHBy8J
SFzVj3X2oOuuwriuS8Ni6O0wHX4SVhRcbJnYQIbfq1qcbESysAcGJQjZlUJ+
uOOgWwlM8RGCqCWm+rqm0KdvhCJURQWIxHjisnZx0rWdQd42NhV16AFSt5BB
C5XjUp3DfzWCLxdxklIkj7Oelm0QJwy4KGsN/BUKZ6XITKuWb9RTzluthrVz
eC/7jLUSx0teMJpPQ5tWN9KS3tfiWxbv4phhSkCBJKTP3IINV2iV6x1s2Bng
YTWn3/ZmZFyRKq0avlR2jTnG4tHp57gzwX2PIOJRH0TNKvEkCHNHnJ9inpqq
M7bCKWNmD7n7XPyL+4T9+VKByDCRVrMggaYVm5dNDr6KnfCidcnDc0LW2FAz
jw8k6Hcgwxfq2Dokyz8mPtPYEsK5c2PMa8qrtdO2QZ3/JWJFeuwF6Djt7Zr6
YRtwuFkCf12uDLBp9F7niaKuWSgf6wdNkUVRFFOs48TOMW3aRxb88vr67go2
svA/bWRtnPurzCugxj+wfC9LzMZSL/dGtsoktuAdcfmpYeR7811lUW6ugZes
DjkBMOOSmGmkOgodUF9XnavwDlfGXZpM6h1lOZ7Ygo4Q9XfGhYTWfTUuuuah
c7FlBhM4WZXdx99n6BXbl3Dxe2EgQDIpL8zB5NbGyfySW5kkqt6LjWsON7Aj
XEc8Z1MEjtZGl5LBQcingGausa6VKSuX8AlRWKQ2/6yQXZHJzo9+ozhhBGBS
Nzh6oM3HdKTbWzAdtL6KmCLnALrNzmK8MnF4VQXowepcNfKr2YrETO0hnrLW
KcjUA5PKC+7xUNu8dGoejN/0YtMB/VrV46YqaLwdMl7aWeyhPr1kRhMs29cu
kYl/yWDPPdB3mBjK0lgU3ZKFTFdzo43Cd6oT+gBkdKZQJXsrIaZgQyT85oms
Ep8VNOH0vE9056cHNLCdFc4hJa2X2ym5VJmnaD0de82lSfyEFhHePRmajUP4
e3fUDN5pNIOO1Wax5eCbRUKlhl472rCKq+tRuX1joePdcxLOiZ9oZ/MYiUk0
z1vQn+WGy5W26FhVjXU/rA2aYz2n7awnGodl0pGAOPklTPgius/O9+OU+kHe
T/jy+LgP7JX6mppzbEbHfcwlf+oOaR3X1//VfK3AGRbCIsLhgJX+TGU712Cw
Kkxbi/8xiNSoJNzCMTcDEEcaI+YrH2OpJCiqM/5YREw+pxTOxzY9DDwhVozG
r1g4SP6Ze6UEhysgT+dA9DRrgQm/cIRYR0Et28ib270GvQcA+EKLK6Id3GHY
BKuVP0/oHjUVJzwjpD249+SLfSTBi/1dXRLKfXgNcaQG4y7cJSjQL6pl2c5X
OkluU92kTSA4J9/f6lZV0ldoADbAvxMk/LdzzTJhJJ4ivwn+jICoY/ddp+6M
p/33QQe1xTBk//WyqfUv47eiQzhbIp/e51ybsqrnvB9DCrhu/ScmakrgzWWJ
cSo/JqM2wEowc3PbYoeSL6+HNxRySw4rKOQ+mgaX3SXM8VyGhi+5xjjWIQJa
/OwIizCjQB9b779JqNR4mFwZVkMlYI/HoTv3INQf/d4s4iQH72aTxhglcNxI
pjQ9I4Pobo19DB7+7nkb3nyirO5fPPzVXkbFUmzw7zay9ipGdn7sZLApCwdl
wj+cRXP76sH15bYynKru/LS/wOLpyuozEwG8kUBQj2s+FICBMGPhp/V1qjQu
ziSXDTdLZCedsF+PIXAEkJeWFXf1MRAz0uY9lXKfokxajaLol27J7Af3CYZa
m9+oopZ0gJe+Z4ST/EO7b6a6rxZKAkmasRdK+728BrU/8Bz06e3wHTwDrKxm
EJJqWfm6XetHinWZfJ6IAP6mX5Q8EdY8kxjKZKHIMpAfLfQduTJ0oiDNiF/s
wSNs6xeAGCzKCEg9eR8JDQO7PkpnKZFroLUvLx82uAZ5CfuzpxZsBNm5dYV0
CpnekIDYn1CNFy1YTDHqiROk1bQwUCSjsAVG0GiDPvdns6ApgMnfnlvGo3yc
VBlgw/kCg7aSspU2t2CHAbv0FJ/HoUm9j/JpKXAm9shsfNnCAPBVpUUhqEeO
++1b+8sBwfFtyyTkDF61lIfOO40DjCp2YdC6rk5HVCEsy0+AlFY11Xmnq2C1
G9bcPK+7jUbEz3DA3UABazqvgieAT9okxgiyBqt9Q2YWssHUVtt8/0D7NZqZ
r47b0DMap/CFtvPCHj4sLJaG/s3frLkOHorDUDEXNEqZCyRR02NEQIU2hLPN
A5iOpu0piLN/2neEajUq5md6Qt3BhlXRuNQ2MlNqOCUGKLN6+uY4Eh9UwqYf
7GoOE+kweK8UXDJ8Nlphe1JR7ug5cFCn3VPD/gu2nJm8LUF8TZMAVhs3CsRj
WVNCzJ1yxqhWC9tJQ7kOpbukoKUfN+cgF4hWNvmfqG/OeB6cWbzwPM83BwTh
kY4vwBOZHI7ms27aUxCkcZzxSIQD/yjA3no2gjBF79GZcUz51daiej4BI2Dp
TDB/flJfIjMtiFgSvRMawYjKFULBMWclovOr7hlo8dyMKF1c6e0kjFuiSGPa
h+q4JY5/H8LQzy2kcdeCZjHL6eQk5GjORT4StZri+ytoyB3wy296ldyk6zBS
CzlwJlEOJ7jHfPFNb4GvZKlyuTvAvvSyVkNfInJ18t2GpUVBsFvWJTC+B1r3
eUybTsTrBgEn+d99FUmmnzY3LrolZKqK42M0VyhhvkYXzpXTK6jdTzhUi4bo
8436sWKRtJhmzXWn7xulCqoq+BwsDsgBHxvX8gxLuLbXPl3PL5tackLhRiLS
ERif3BtC69HBU0JP9oXvvdRHnlJTChuIvydfTvdCfhgNOGoK7lNoKKWTKUhR
QeRgunUQs5ls5K/sAVfMDlryTxOZpYOSGlj8TeSnxULhYkwCuOjzKDZW+UmU
GDpmhwwvzoxdQqoMTBirTqxn8BRt6vluhvrX0gv8KuIzFGDTLLqXMT8cK3lr
H+bldeG1df0RMM8q043BWEhNMtuuummDvEJzIaD7DTK5lsOrnAp9BAhgacpY
1zSyujiYApzfc2f4v+taXYKB8qCKqoaaoC+PLx552fZJ54iH05mQC1dGwT3b
zPtfha05Y9Wsq7DWOkebCsy4tboWhVBCOMTQNMp6WroVJvcNmljP61nvPmpo
xxkQRpDNE12x+WiJUsuNGMjH3Sbh+ocYZatY+6wxLyka3tbUTek6TCwA7+uc
vN6uZLXz3VhQUXZePc+Y0mS2dAmsX5EImuBDEKJI3JMBWOdtnPN80Fh6KBbg
gTvEn4akirGraUBBztOaVixZFDfYfOduTf/B6V6YpNDAD76HlkobLc151L7R
krpTSUAB+ystJSMh/EaY3r4QO19R/92Fw2keS85LZo2VnOPE1qP2X6ZlIJBA
WWseQjiqCdtTUBmogQlsqElwH9Tp4sDNtsI5NgiMx7l2AkupkR5+YUilVIHD
MVUau96aIAFW2bvWKq/+HxVfj9Ms51XDpIkUuiTREsqHn7cXkqt2fM49MLS7
1Msy0KjqGu1Fwo4isJddYVguWM/SvMf+NDkYTdcPWPsiqN3mMBIabIkm+PjG
FMDWcY4dmu843bxPQ0u8j74naauGueHXUIrxhQvL3bz/KDGwBB0MVCqdrmun
QJ6RH/Bg/A78Ke1K+HeGfIyeeJjb3DAzUSvnznN9mLA4CZrilhXCVk1NMBIL
W3gKD5FzMxZ0jeOS/nM/aOdiPbCe/YUuHQR40B3ETN1Wezzp+Beo0iyk9f/2
P1/SqZWr965IaX55d14V5XZSquOLWN4QRnwJ15nLrC+4MklR+QpsmM0jt7on
nXPkZyrPjERM19sGb6dY3i/ZgK73ULmNYeBMk87wcei4fCvnIQPFScziI/bn
7Dx8XDHaIQJcGkuV87+j3oGnxSve2dkicUx5BUHhoOKG9wcDZbXTcVRTfkoL
/pi3U/zvAs5hfVCFAhvElBkxOdpsLboj7URv+BCS9koWkdFcbCDNK34Pmw30
AbqpeY/emsGD+ULI1l0AHEEVcag31wzKWV4SvDkEi08ZKBfeQ5g8FZq3ROSO
3htcUMsoa/QVOgWgRYLHmA1KqEx4D2HTQ1O4BJm3g2sotAeCWa0gqqpZ7xC3
tcqNenLIWXYVrJwkiptS/YwLCZO8lR/M3jqhJ0/vs4juc7hMA2LhaG7f1mOL
heylcIIzpdNN+iq65tnZ96KrfMCIVEfvINZVY8BH/1IUmC8zN75DLr/AcJUv
azpv9CqRWqUjB9AGwwxvdBLT4EA1aNhpTTscSMMzkqiUfSxDnlc/zbcl9Vl+
CnD7key/yfKf7UbDb2Iw4tP4u5VBaikPMcmq45TOhEQSgoBO6SsKV/HRu37N
5L89C1WidfdsobL/sqLkxpqBCFq8sMdiBXcKTQZIo9t6WgPhkRxQ+stpwa6e
c0TNUFPnUAS81Yt/3IENbRM7WmM6j2IEQB7o0h1rSaeD5dFE+tozBmrIGapP
EYxLjBevfL3XUTzyBfho/wg7TfuTxdBpFldU1jc3AJwVEh/3RcAXnfTX2wJW
ceT/NDQEbhvyaJJd1amY6xbXDnT3v5f9HEfUoRKC7Ji0B3zpju7kF6NCm3Gl
F+wXSOMedMNOI5UDaHlnDkhagv6jN7E6xHEcmY9laMO/UyGDdK2c6NuVrwzK
0eaWuLZjRzoEep90tmGhdEG49l6aFcG/kGMTmf/+zHwKnQEhYcN2icPj7vkA
n7t2VPSGO1L70ykce3TugEyo4XH/yPHLnF8VfDYse/bBK5wtqxbSRhICk2nq
yfmAev2YUMx+bQ/kGxNkcYLdDov368EeMIvV44FJC9vAyn7CZl7a6/rvh2zh
lgqf3mjWeRvangbJEbAz3sZmzfMZYhcK6h/ya1IN2X3oRDiW23Ej77R0yFou
fxIbKEgHk5xL2W+NHnT6zr3thERC8uqd4Y7GKxV8E1DjpYGC+I9PCfRdJNGZ
yKhLX5c4Yt6uR01ImikbWb2ZnhR51rEDqFqUXI58x0OTdxXteDXvk389rmMU
tIu+ykgyh/KM2M5qu2eiu7gCiAy+ieVMVooBkEVibR9t8yJd/A1Mn1fyEKVG
iYghJ04PftshmNITcrtU4SjZfyO8M8K9HtKS23RZAdZ2mOGpoPW3JL6Bd/PR
AUjxrEClb9BUOpSg1mMgUfCxLNIwZ5moB74ytB7FLtbrHH6OzpRCmFaVNSFi
veFrEWK/rNi/CKbnKB0uSWr2t/WGDO8DZFAikg==

`pragma protect end_protected
