// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
2lv6sKFFhmAffLWTxXiQ204s1UgHtvOWPaIjBJSqGfmF3fBgVwYV8FlGGx8lJZXI
HnQGUj51hjjXurn6k6VZO2Vg4xk9pJCM1ZTpIy0OML62lVMRz2CVuvFFPJmRSRec
WehPQeJva77hUMwm8XQ2Ge9sr1yuS/CATbG+GpFyJ2E=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 1328 )
`pragma protect data_block
ndJ7l/5ofKQ4A5RVs2P3UanJqlZtAAVzOKttMlA8ZdUbgx06A5umw97f44ulk8ff
a/so1GQrDWXVXz0ZTizdd7aa2eXOcIbZSrpetkTDoESwKAZpPuYaz85t7AFnQrAX
e1vEvgbzcJ0W8Rbuh9/mwHnicdfP/GVdDFPs8kUs6CADl/ZUYZflduxMq0H7MQoq
erPpgKM+V0p6p9UlgKN0kH5kMZOZDe37GbXbCj10WkkMmk4Dwzklhyt9gIfDySU3
sWadY/7JVJfUZS308Ecn3pOJorHzyUZJVnkuqZjjH5vzJpuMMvmwPRQ58sJU0bEi
meUwg6RNUEBq/h7SKXQYM+hacvHxv9iTQkkLj8ZfTooYMTeMUdgjIqBlmzdcx7lR
Xh7CuRjqXjKxmr1QvaiVUhNbt3y8yKtQf2wK/+Z2BGHkmobfxXdBHv6s5vq4zZ2j
bxU1z/brKasyuHmGc1WbuagDGpKXfWud8gZMlq0WqILDzAyOY8IO5CPBT68KHqhe
2p+9L7emyX0gOlmZ3wRKLJVvmynGcRSGwToCHG8wxWddf/h6fEnOXZGu1OLF5I8s
ITzZy81iZ4wK5UG4xEliaVgM+SBhq2KBgsqa3J72qFIYwAQ64ku4AiAt4aPArqbu
rxVHWiAdJ43XAG4rLoYSvkhy6G4S79+eJk8Vq4VGXC9dYS8GetCKQIjKZ81z1FPN
+zEl3BGNF+u5cOgonJGso3oguaHsDoWw9eXvQhMfDg8jLyryWZaKpx63045AD6Wo
eF3BSDUd3s0Gq/B+/oKARcuuok089LLoFeX+Ko/7mxHxA8jGghnloGFoIU7okver
nGRf9Y4I+anZkXnM5lp2+Brj7YxAIZ5e7UEd/V/bCBcYmDureMU10behGTHI6I1k
UMnND9eMURgARlm97Oc0oa/ZQ+r/rjtnoVLdKZVWIXkjt6iOpbFXikHBhbp848M4
05IVoeerOIz1EwAvFc3BZVhFzL4eFkVoqArqHPIj302WknwyZq1J1+zm3+0auXKb
cWilG5I+cAl8gZCmjTBuE+kwrN6pKhqH1QMlS1F1JW4E3aoNH7S/BmC/Bxz0HB6I
uI4wu5C4Ift0P4739TQe8M/c2FPYyLll2hz5A3D2DH2WFBeNTMYPNHQ6RPcpTcNm
aB6cSXp48IVKEzBSeoWeKpiM3Ihj2sQPomtF0kQZLlCrNGWqaaftuanKJVKO3/11
XAXMtVuw5+7GZS46FFQH7cIKb52dpc6ogO/BSQ48uY6PIh3EWrJohfUTRc2dLG5u
6wGenonB80I9ckOyar0FZfULVj57r5fiLR+LQJO/PDVnwJTvwqsSBJON+kyWIBRh
G99VREZWgm5+e9nVVfiOtB13e4mMeOx8cQ9FtDPLgvwN5No4CEtZl9Ucl4ILAIWc
XbR0jMn7uWEknLM2zvLgRhcSqJyIoKAKg0VRNLRbTsizBotSekI4l1QNy6DzCpsd
a704OxTFNe2Lx3DrzuBVy2jlr9Jln3ip57ZXZ8UhtMMwvLORBQv9PWeTxmXYih8H
7j5cCei0by9scYC2sjK0Cqfh/P0r1EPBJZwBdGpj77rA3lipIY9nw6hL0vmosE+k
BY2q3t3BxJfSJS1hnqzzos94ihM7xAyBhAsJsfdyrkxv/lzUiLxdq5rCyXQDm031
qXVuyCsEfapbtee9eoJc1xJsZsapHb2X0jfq8Epas0ZbD1Et4K3NaBPEDOzmlJMn
uzeqg1dEgIpnemlbw9gyfiRvBd2Lw3DJnWZdrXUhyWg=

`pragma protect end_protected
