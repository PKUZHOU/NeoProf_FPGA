// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
Mx/teGTdZ7U6bnjTz4Q2GqnUFV/g2wyXM1Huzmb1H++WLaATk9+JYr4CECOJKhAH
qKceaw0dSZvPNI4knKK3xmoi+fDWJEX5UvO/9MgeG6Z5TXAmvkU4w19pXxBAPGA5
L+tI4gL1Z+CKZRAlnjmqTQjUHgS+8ZqIe6IfLggZcjA=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 26592 )
`pragma protect data_block
HmAAcvS9K2F7L7XxHO/LN0Y/PLW0Ahw/3hdM311Ko8K1WT/q/YE+K+JQO7PvwsZS
uGSaQoqmoIGUvF93oNZEhQu9DBRRhaKxTbtJcZn/UywPoRFIS3Vql53W7llQ+8qm
vQ64k6p81327wWs+Ge86gD8MRxnqT8Qeo6Y3KE5ackYhUdtJmy7AnhU8oqhvcpew
xV35Fk6NJ3yhB85VdyPkB8UdfNBgpOPGK10z3zJUZ+oy0CFvyJQlCfA6904ffoAp
9J+hGlHfXqqa55izwMh1m2OVLM/z9geaVb+mnm7vA9ntccdLV+k7t0nLftZ0J9uC
9nRqKcFJfuQaaKn6y3W1kKrfEPIduRGAjk9FQ+q4/g433dtAQjCgnHzN3rVZglib
wJDJmSSBfM49whdnXxAUFMxBOjeg+oEdX9UbUM0DoBKlRYXZNy2eodlHsBuaztRI
RuT5r5hSAMdjz1cwnEh44CjSsB1B7BsfalEed/7MGPEf/UxIos/bCHmpvUDMbA9s
KW/M8UdMj1RrjJPQ+43OvFNn1+EtbIafHWo+Uu8dX/JtNxrpK0aAwZ2Iq91cURaC
p9MW5FLh+0yNzLsYUI3/icYk9LOrLYQJ8lYDf5q17o4y0dH3k80tPlQ/75WjBtRM
Z/wyEvkGpGzn9vOEM81rpJMy3dpEbO2vnCU5P9Koss6UaCFra5r+I3y1TiJwheRf
ddaIGAQMhnGvT4OIQTX86zZBv3iQjv0Jx4LQx92ZgiQDaMayVAWySgG0yEjR5WyC
9/wYfDGSY/rCS9/V4HUEW+TqVncLKbH9KuWXkR7lsBUGRsFU+8PTA9opLIEsysAh
ZOf2RyaSWR9miDXkj9tyuouA19IJPS4dQKRSuCxH9I9Eu7Wm6jy37mtcFx93bkOZ
mTuzakVBUNIz7Zxmvwbec4GXG5J4BWXY2QGcN0I2of6UK8ybJNSwYARnLcAAY4Ca
hoRI6yPRy53iupN93iyOczXt2KaG3VIjpa+xq4WjeJ+R5GzqO3JyzyAQaiWwxHj9
tz227AdltGnRDZ/srDGWsRHgOEKeL8thf/BqRhms2mDZnZkZaJanj3F1jSTj8tdy
QdnCxTMt5oMD97F4dDkpYESll2vlo406jJLtBpnR3qH1yYJGbhiv4kCzyG0aVyGq
g1UmGAE8g70BxIufx/rXX04PyXWAERGQ5MwAJG8KFZcqGQXdIxsh9EcIFMaqL+Dy
C7ZUlxNsSAouSnveS93bsyb8CykXKRt7j4ySMDjqFWa4yKEwNGsq/mb10XcqEbkn
z8Md3CpOEPaBiKfkd9pYTI1Irow1dotjCO4okGE3cge1L7OLU3lgGikjdRiVZ+7+
4Ol/cwOUfU19LVtC84/B5QdhO6c/OlMenVoFiP4Dt11ThO2KYpRwsOhUinJS4CnC
dAKa3pWU24EEICkI8dWBsXYPDkk/tRbRx8RqsxA61UHlPcjDmHYslX7AWjxAxe3A
ijVYjfwQOn9wJ5DhHeMYiJ3yfzRMd71hZefUBi/nRkO/VeVZEc85aeojK+sv6HbF
S8t7o+II8hwSl09yjtEJ1bDpXIPRURGQ1JkggQ7mbxf6N3XmAG5K4d/AN8uS3Ipr
wjzgUWUDWeCzdwldpyNAg5oWNsdEwGdAWhKjTGU+1I7KXZPMqYszfZkFFkZ1W+vs
zi9hqt4RK4XAXiIIyNJiMFTqACfnUR31ybhquhYN2Yoe5r2Qcb0qv/2Vqi4+g0c9
vc6MNyhLxQoj64jo6eagTGbwGDkjmxZOGGhQzTRsbOZIMhTBxFgYDbb1aqSgVB0C
wsKo4LxXeksq1ta8FFDV1JbRTOeIoHeJYQ0+Qzby8gp/5ZWUCOO2sSraIfh3jeER
2cIrSqbaiQVbdKjGsiNRnvpFasE/1VXLhaF5Kxb9IA+yNiQzKdDiLxTAZ1S/6yTI
mGLtvyKkQjlvt9HS3B+TCdBOoeF6nGvs5OOBFqaoPIq3dN8rp3ryn241lWogp0P9
z4MgJZ/4MJWf9sziIOQTn2UigqpjZP3fsaP7I4j0B8xeUb2S2w/2XOopj76ZjxZ9
dgyfK84+WBAAUkKVRcA8m+vQicEjcitAyWRBY/ueHH3/73mr9hYm8LI3T8AfxvrL
VtSpXZANfoRCs63NgPL+Yff00pk327cmDXyqSqlCVurt2n+sd7NOJvQrXgQiyIDu
wPu4m1PPV5sigEGpSJlLO0MwzUVUuM67cA9oIvZGmYZBKVnVsHTg18dy68ITq3EY
4os3f/0L1hsvF+r9VwwH6pPvZ+eprG5ps2IIcpkLR/vOGtPPlbl7H+p1auXdaREK
iJk3CaIrCzj0tVuf/S7fG13itSuf+cskwid8WFoGNWdIxlhVICXVI0doWOqB4yxb
sb/+Kql1KmEqSFsMJ+FoJznh/fCD/Nentc/yW+lfqdRpZVVZSOumBYJlgV45PRoO
IlONrDnOyUzS4Po0TQR6mogKLALa3LBMZ0ck+5G87O4WMIacs6i2p4+YlIU7qpCd
6IbFn6KP0atufRRaWqxDstKc2qLHy3FmgSnUmQ8u4vdJkoSfC8U2Hpwhh4X5Efq6
v4A0Jj5zFS7Ukg40a7H6Yr7LnUMdu9YXnKNKg+nAvIG1ickHnQcDTCyQuXHD7p/e
rMG1hBXulzJcFuOnyzqDkLyfOAXxMMARcOQCp32o7UScdk6LEoSzxstF1LCedznZ
jUxjOI5zoxrcMOExOc8uQpPV7QSkRbcKm7FYx8Uuki3tQNKk2BvwXySiI4SKntgz
fan/6XrcFjQcuDdwfGEpz8HJKAp/A1AKyW5PjjTEqfmS46LqaBMkvZ1479RukT6S
icWjsJ9QOtGVQDZt0J0tbO+/zqoOTK72nq5WFuAUGSHYK80FFx6YzRAhUVNZn+MY
jjgmh9NGdxl5ceKfbVPAYR86GK2ZkYBekPi80Sv3yLDjpxFWfcLQsLaBUEj/+NVD
TpGgbjusu3TqWbWQyF+HjkOMGgpBGvKyuZDVFNHU5P+vp6W5VwXQEiqYtew2ji0z
85lZ6CA2G3mRYSBg1DKxGf1xmDMy4+nx1I+49u1UHiX920LoGGnJZv1783qlDUsJ
buLP/oTJABKBI/djP9bF2Gdg7YLUZRrOb6+gG36Qt4spZYMUz0yuSw54JJE7YsDH
E6MubXHgoRvkJJM/mnJwic6rVzi792S87/gsoNBGR1M2c0DTcG1zuvplyMbwx/7p
MviBD7BGMPWEoCdo73nEZXLjr9KM6EA4397p1bsfg3WecJJw7Kd6+qoGcE3iylXG
O8OghO//7G8mRZtbFuzyZ6bvs+HInCmGNhC9NXw5QsBySQzNW1tqVsUEdLmc0BWM
Qrh1iLF8gL5r5msA53auhR9LIywFCUbI80HV0eUJSMd57iiyeS8ZPx3iZvEkwJKu
tyRgFURUgyyfYcDCQ/HU8dHCZ50HTzqhO617I5tkOBpeUvKh7qSakNkcWAuD9LgN
YwYc+S0/ABjWkF5FvCOtdUXqzfWcqhASQt3R5XtxOdGEynzoSg0BWf4ufAVoSPwM
opvtO9Ze0chcPAR1+MY0pz6D/XJP9+Alvgslvo/vaS/UzbkkwyUsz0W7uOp6zs8/
r1MvOH5jsebIZZTye6xFivjvvjnOv+N5VTPfYeEraMcd8Ekwf5MZ1LEt3WqKR+JD
fkncBQksCyFS/4ZIdXWwBRv45aUZySzq7FxYEmsZ2pVtaOEYVnQJvVvhHZGxFygq
52IRncwJoGQOKIaMefQFihAS77BMftJUtUUKIhoDOf/IBle5Im7DrqZutok8n0+d
BxwXAPivOg+7FgY+R507YQBpu8AL3AUVWUeWSJ1KdxXEnNWlhmt1DaBlB7BC6T9P
EzAWZm6pxtLp+AWw2mbJOHfE5QWz+IY6TtB4ooRrbyjJjDmPdEYRVQKZy6JMmCSO
h5wE5q1O76ck8c8w+hsdHB0kFJF77ECm9Kwc3CnaUCysw4ytqLhBKLyaxxCyQC76
utNzdKuGrmv/k+Je9airkFuXUyXmRR0BR++JL5GDH4YkABiBVGg3LCSTvBGJospu
fpPZHsijz9xNfFsf5ZRClAApRDcETrvl3PsTVmWfxkEk1DrnyjIATVWJ2Y3POUn2
YKnZ4G4IHPpSuE9BRkKKx3kz+6TEN8chOPI5e0gEbPip/yM7Y5gNdk568IFszsFU
OIUfN/igxTKrrelozN8674SPQmwfYfgiD05vR5IjhvwVuPweV4+/US00QH2mVO14
nTORjg2yAe2WgJjAkpDFARvoWkTnUSlss2lo2s3uFz/8wuj463yqM1YubCFB7xIk
vvNmHGUrPW4o8RpunUYdD5Lm1CVgCc+7zRFzgEc28vi0smXzeSrKwJ9Q9d9o5R5g
jr0oi5p0d5Qfm7O30ahhL605F5HT+r0ZoLgW07c4jeXQik1QlvwVXJVWBlOAXy4u
YyHa0XgmndazVwQYe4rFxCSNRyTjHjO+VlzO/OO7K7KAP0eZQrogjR8CwRdQ2sxM
M0qQ/FxWGPFg3atPajtNaCYpl2PZ6CC/j1mwigr+GDQTAucNY+Xyw7+afshKa8kN
RqYColJUzCPeuxwpfHOr3/LVdXJE+GHdRqr3/eYcGLskN7WEnbu45Gm3WsjGQLGC
nIsou31pKYVRSRU8a/YQZfAviDMc8MASUX5QPV/m7Hk+5ZSi5xmQfa6uZiUVIhm7
c7Yw9tNHSXGFhK7uoCkrROhbv8AwYY4Ygv27Qfqd7CGqnEMOf/xAz8AI8axRKIVr
tcQCwpCPQeDoxTR9nT79dhNqCsDAxXq6t3VcEHHOblTGuPNyyyWaGWC/19sQp1+P
uyDYVREfbF0d7mEq1B3hoeqzcYXcdBKZFzFwkfSghKWhQU/IsUEHphkY9pvXChgb
nZLeqFcRnVwmsQZFwRFSyxxjATAG16QAZvkl1B+4vsWMmcNMzr2Qe7AGiqWm3pXS
2kOb2e4YyQr3fwSq0R5GHYCkzsuuTFXY+x3jh12NdyBYYmUXc3UK3hQyEqfpeJA2
hHdjGNehl+YYdShGCbrc0xoVpw0sZSCYfnV8udizrTvxaKdcWDgcnECNcOOgvonS
UCLGp+ljpSDKnhCITb1ZsMKke3eIGXErp7CyKChOuydHky0+aspxgtFBSzvkR5ip
de1lF480eA4Ra95XVN6wLbkOiAu9rPNB0rQ9q2+oJPo1p7yaObXJKtKISr91Snxi
XA+kOuIV0YNyeYGIbiG97iuqlUUcHQhV8Pl1NzLwff+ET696C7ctgj3zXRaVRhTp
cMlCCxwa4EoxR/FWyaaWfI88MFdOCmCW+DHJZoI+o7Cdj809ADCfN8LGLrwX7QlJ
akKq7whNI873ZGGfUINfSW4OAwfDteLZtapAL39Qjpi46JA/pMIQf1xWrfxOCdaV
LttTbSu30xEnrB1dB0Xa874LOzDoWf0/lQ1ZqdMbuqXTC9VRCjUKIx034POnh22x
OK++BbgusmT5hGaNYb9zefT/nTuAnKn+505czwOBrCGs2AwuqKPPM17d8WkEdvnS
OyC0J9Q3w+M3ERn+3ArDF3yUROBVPow5p0VxdhSOmTHKJyI191KMbCJ7d6+ZpzBE
RtYhN6RbdFaQV/t2oPWqCWfGu98gNPNnOZQ64N8PyPxD1SsPGiHXzG4lllAqdORr
cy0pTNpJtqnki0HQyWUxP1T1Y6kEskH403N44Ns7UdEXw3V4N1uSsgys64aoZtOB
HVhkjSBOFyWMNkQZLOgvsw/GUZnfmgS1kiG+stVO1tKIpanQOUSf7DjRX3Gbymxr
0Lx3su1OsXJP0WSRl+KpoDG1OmLKgjyMJEeGAz9mzMJjujuzEjNF5ImaN9XoBV8r
8xDHljMJT6h7nwkckB196e8m2dqs5A61gT8bhGo1j2W/Gdkdt4lIA2n7USJXBRfZ
sb16QjyUrYFYNhkPvHzU731pDy5kRpz8PtyQa/YCArHEPusJJpFuyEN6j3AZfBDL
ZycyEf9ZqoQKa6wTQ17HQLZWP0ZYQPCVfw/CrJkZIPZamFKxqFxSHyQnZA4NB147
cmP/DkpWsDPtfSsiUnPQTjyU50jZF89riTWTRWvfjd5FzXBK65NATRdEXGFCS958
UBNvs1UTL4GkHqcWbmcBpUYP1r9m5/9N6s/Sf+IeKv78odP8WWWpW9UM1W56NUC7
th8zcX1IDeD3Xs+Nj7cuODdbfl/uPRrXnb11kOi8Gjsfhb1YipNyAnpRudDorgGs
hEAxGHJodl2RoJwb8JNrZAHYFOJs0FpIPpgmMlR0dWIWqm1w9+BQ5cRukcWUAQJU
CFLKWQ4zx/CyhJMyJGxk4MRPqyBGlWLiMbFVOjQ3kZhyVXEzlmk3d286rJda9pKX
5apFwNGDtVlZTP5gQ68ethlPNRGXdAipTP04oSEptCXhscpa7iQ8//C1UlkJ/vhI
oT+wnh1P7O4yevd1HRLsa1KzDn1io5gNDxc+wJ8kY1OLgBAxyTquaZkI9YXRWNoL
rCWj5V05PUeXfkGaUAGzw7Uz/cQW8FW/2vTEmryY/frIK925vVudJFeQwlkeFfFT
7TiQu3rvvbe6jxaw6a/RyvguvSjXbAw3Ll3Kv15PlMo33hDW/dtDUf0CoRB6SiBE
/2ytNFzO5syXMCri4hafC1HPeHxSlV0ERm3+2mS44gYCE3u8rjvAJX95hhIpmxJA
8SDa/bFTnPcSkxIEcLThWLWlRE24tJy3bhocynNbMQAHGQBmGTOdxyyN/p9apTx+
sQEaNz7oR+uAY3JmpnwWa8prFryCLhFgsQ9D7G62hqTKlwN+jFNKzguFBW+AhyU1
Jr3teFLTqMCthp83zZ69eidM7q+ozlrWJU1HPTDsnrpagyIwpEsg4wp1zXOTMUlZ
ssesSZzslugKKBpAQDv4PzBP7MOjEB5v2wtPfGtzmty5Eo1DVkk/QXPJwxkwdTbY
Q/A2f0nE3Crh/bPq3LVyN2EBLQTVdcLqXJ2shCfK/ieOAQTcKIO7UU2DhE7YwB7u
46OCLhSzt6vdJmdtUe42BS7XnkdAtuDEHtpQp0nQipTVcUNAaC/ThlJyIaMALYqE
SzaIfKT3YVEiYtjm0dwdm+Cf54o0Gndj/iFlmNHkDG29/Fb82LmlnEFhDnXcPN4C
qT8+pje+YuElXrpODWgBblP9Zj71EkdovsLgRUvuJxpnQ0eICo9cpM67E3f2DcGb
MlMD27calVHtKM7f9eLebcIoxL+pqlvIYkhg2kl4tEWKmsvFj6EY2c6NUkTPm/zE
cuMcK7zPAzP2ZIiJuVDzlRP9qREq25XQNWlOV1GcUxLpvpTLcaQL9FlGRwdFhAPl
F0P/MOF59yTm+b7tIXhaNJVShdp1g5pAG1zR7J/QGkgCQvhRVNAcQwo6b+STrKuo
bLYtSsKZL0DuUr9TC8vJYCy0nrmdn+Z9BoN4GZLCxjRvHC/ovDSMWtMn5bVAGNVH
OD0EJiTPkMTppjrwUV+pcWS4G+QlPigKB+ZBAVsfUXfZXSyanj194vfJgc6vxjrg
xmLtEHycZhWEUqJu5aYVzrXlBZWjhO5tf83SQUL4LhK82LwXZLjkB5qVrmc8SAUL
L5Qt0Ifxqc+9pIuDHktkYXTHD/bA9gh0kBwyHzJNBwIU++FVauemC91UnhF06fRr
nQjYloFlooDD8KIZwrwN4mjTHhVu/ZMmhukMhvizrKORWchN9dnDmIc68/98B3hh
6PZFqC92QDBe6jBEGtnygUuiol+yUxbfG+/DZiNNUAUFME1gPitED1YuW6sxVk9y
U526Hemsx/RZVxHekWAXKpMl2O2Fs50/puWBYiEisFyWpOAWb8dbHQPY8CuC0baG
LJDO8H5DXjZdjvPM1Y0whV5h9+MI4BkezZPtNpmZgf6vnogqDpiOf82zAJ+gXWmQ
XtmKYAcesaHqyM1pddP22M+H/zdn2EzDvxTkyw9aC4xzK04+7X/7qDd6JvF6CTHi
V6ZWGCUt4BfKE36TzlSOJiPkHZQItaEzsSb8n5cqyw5SAYRiGrngV1mlUnTCC1Me
JzRDs2b1BQCsk/p9KMmIS5NhYQdlRPhp2GyQ188LqSlwwxZyXuPlT/EZZY/iBCYi
Tl9xIpQAG04PiwH+MLt8qZfl1PDgcEi28ywaYQEqIsNQ4U8ELc73ygChs/wEddHU
SX3jtYna3ISFxNoDjBZK1b6Qgiao+ComTWFUDC3nk+5F21SttQubkBb8Zww6SIbF
YE2HTlllk9BVHhFaWnhMhoo+tlyDzUtR2uuE+Fg8ivxvM4hs6rZXbhfKRoF7ZuIn
NqrSRSRkmz54ADsN7sKiQaF2y+QIbJjoPi9yCLTeeUsFE8twP9bOiMXlHxAhcOHT
FaKigYoe+PU2UWVvFqjYEcRMShqbisirqeoWO8pBrnMlVbsFGveO81rXz5ekfW6c
WIJQ9aE18tjstgw5MnFdo4a+GSbncOIrKiafKFpy+teXEWytARXujJ/BPZ8t0fAx
4MsZ/Iy/gcbRFEKhfemH1VXIdum8PjPlQCErw2TX8AsZvQ8D0oT5tee9CdztevDz
ZG2An2zKVw2bGpmq+cOA6kiaxoF4ajjBzwdjifgfb12BfrwUsj+u+Me7ox2HmeXv
i4HH9Ua0Wil6FwPscP9jrvMoBkSAd+Mtutsp29ZL9vpGb9WFBk4AbV3gfoZNeHms
8RzdTQlXMJJpddY6q0VF0sRHSb4QnuDK30iDALhaR5KMiB5e1O5EizkUStwF/3x/
4iCrPJOVzLsGx1bucf5sOPHZxqKxcimZED5Y0+jCYRFNxj5/gd1idJ0ot0PD5CDs
iQ746G6BzsPUKUYU6KAyaGHmD0WnLSDd7s4NINjkRACLyiqHcjbRbEHKiZpPcaIK
1ZZlzHYzUcx9nZjo1OLa+wfrCUTIBPdq0hoFBZOXmO329A4bXvg60a7nj2SXEPK9
ytRkMO9U8haqvKoVRaM6cIiwfHyPVpcQaWt9Y2asGdvA6jx2sOR4G3ZUoczF9K93
CSPyWo1Hml6957rvnePMiEsqcG48NHkJth9whITWS7RJOrpT5ksTlHBu/KuYwMv7
stYIkr04RpTegcUsHMGf6V1J05GW0zibLj1lYktZVApRltIZvq+kjtq84dsq+4Vb
Lle/EQXQ4xACuQIQcBqI7CtVOUtCwuVoXGl229yRF02Y7O8nfREw2hR+UtBD97aP
EvfpmJ/UJ/a2GDCopGOS3NJJT1gRZZQv6tI7tU06ZdFZDm8XMiVoUUt2O7BBOCZJ
QQqxiipXVI9ITfoKqWi5qxQ/kA7XoYnB+OoqZaXzNMGdAT7AsYwVd3GMiv6iQTeV
an7Xpy4c6kQ6GOJyoiJ7jejy377xLIOc/VcwpwTeDjE5OxfrFe+2EGjTLAE0HLF4
4r8LvFK3sumK/h7S1UQoGr0JfggNXpNcHN5JAI3I/fD03HCEgn9psmIQCNvLvAJT
qHUf0F6aG98TN53gCwvHC+JZJ2OKAQIXq5wN1WjVilx1DqzLMNYm9tRaM5VOWzbl
EcmQCf9QbNcG73Pr21ljH27qvVqvigm+1wLe+0cxly/LTnwsJ3RmHRjcqvSW40hc
GeRHYQleYZow0sofJA2bofY0D7XjqIyin29wRys/ISFgOOdm9IJ/5NByX6fNIbnq
eF1USJF/bxjhJ4//rlR36enkeIVEY6VwF1K+Wz29MceRBF8aDn9GBgJUad9U7fLN
sPOWN9xqrH+g0Qlr9oVXnCPHVsegzKWhmyL8VgmKhemon4R+/Mgfan/JIbfx47so
Hs+Ox0vUT9ejz8LHNouRP1//VMZVkEKwEv0QJFvj1tUDRMGpGHCYNbo8T0vNhif2
PWJGfwAtyhQZfTbrKa1Fq5CKHqL6KO1Ub/XSa42UHLFNKslXi8LaByJUiB4UPpdR
mZkv4QKauKwXyJoObWdOxDpLvQcjywjlOx3g2Bjh/xPtA0G3uQTzG19IehqzdYex
hTgKwxpV4KH3T7I0tP1KBNfwrWnQRw9zOvPZoMT37MqU30WWPGhGQNWyKrc78/9P
4RDAgKWAFyg7C8TLw5uNV2sYX09WYFFltvtbH9NMsIt215VTK6AYfufCdvYNFVUS
kUWcW2xZQ0mGLcKfJvJYZSeB8684CkE508WrTBifCu6pTZeF6VSZWFYS3zO+OdtS
ahWIZakrerdbFSISt3wbqhaaRMAYBr9bQ1M1WwBJt5AdpwEvKSsXBNwvDO7EXDu3
F3i/pKURAmLBSX9VMgiGML/zezuvDTw/z8Z2wzzYu02nxVKU1+lRKXQl0zH34PTj
8yuinVaLT4FKIjKxg8U9Pq3vy0Mk4Cs/xGiU7P1BFXKpsCWVqALcJ7uqXPefuFE+
GCmj+dbP9HxTRMnGSXVnTQZfM0w7oOsISLPCCakWs4iRl71kkuDYdCpBvRKNQVKh
c7t38UX39jNm0gkP7d843p7tQQGVVQsLbPDPr+7Ym4zbh94usfXTqRP0dU0EyLW3
xC0ScsA4WuJsad60Gs8eXVIMkFrQjO5WgB7PVTrD+0Q4qJ+tYIgfiqux21TcGjKw
newPMAyURNuFpKdRjFsLQHpOYpJV5G9qf53A/bIMfps2lwL4SMnsVrTo9+8Ed02q
A+h0SQcq351o6EJ11A12t6Dic+BQCfgSwHF5CCSNOYXRgsUFpNilQrPEDbqX0YnI
weQInMdndfdnnvOXvsOFD5p31GEgff0O6pQAM4oA25LxIHVwAXEPOIJXlQDoZCuR
w3mqgFSE1iiulmzj+DdLqSOIB3B3vhHXIBEHG3HeUnYDc8cIcct4nnYMys7+l99e
ukFYI1cX2y1hJFJ1IhnrlbT4la61ektX1omdLO/OBSD+JNVLmxhYTWdtIAnDSj9o
KTDM8aFpzgXX8Nxs7G0vglgM5093dDRPslRrhRBY1jzkQAWIB+bhWaSoLqjBGoOO
gLuGGZ7lQQjF4XcPzCZ2CFMp3Ds/ByPVj4imRrZzbyn+ioaJN0a7FDYjShV0mnoV
lhi8anxv7CF5ptOIyXNzZpr6GyoSPXdoJnV0nQfCW90bRYxEQ3yFWhv4fjas6rzd
mY10ejn9U8mk8LMPBsWQBmA5EKWx1eIGhTCo+lu592Dg0sIh+o3pQdjGU8+Yqt2G
DhfCIlaX2LWvRsqYAxA9A7/hLEToSHBI9g3ayydZVTvv1soPBGFPrEYLCg8Onv8F
HGLjZY+3yHjAjClJmbjgSlUSbOPFZ7WecyWDCexLsPs2n6zyH6NJ9HB+Q+j5fMqN
QYmoMZSGnrPZFuO+801z/xM0vL83EfmzoAPtWcRoc91E2jTEz5jFwh0yGwR+dBfk
ngjbmQM+uP+mb07k8lXIGpwkO47tDyKTc1ibuX5OzotVYVa43ooXvW3GNlUTCOLp
ulTVxY0FnhhKXMzALavRXHuV0jEyZMXci10FhJe1qym9Xwmu5Uz8Hi/qZylPXSfA
3HrzjMdS5Bww0CL94Zfy9y/j6cBrEvsFV4J59RWXbDbc/OZBF+JNppW0ZnxjA7yR
Q6jvX8YyQA5UNA76BAStb1vwBKMsc30K0h3Oao/4Mq818YQ0XWb9ByGHy87hAfZA
sgWLKlsKSO53P8LiThJSjojM0Uk7iPkYVpj0AVYLTvuywaQ7P5iuzojVRTBcXSpa
WbZRb3pk+lS2SF1yB4jVtdXEkUoD8sKHjXfwICiQqqji/JQO1TLxAv8PpEIkxEAo
D63/W8lS71Qq8K3EGA9pM1Wmg5aDU93kpPFhb7lT6m0Jy1FFZynpTwVoGsvnsm/R
FZXrPLzBe4BW+wTzsU49Xhipwu5q4uUEiv3KUH5ef+PvmJpLoq0JIQXQ3x/+c8y8
iwn1aGSp2RyWEA/zgYA0Aq3CVJJDEyvz3WVGPAdPVoTQ1vO/Cxm6t6G0srPwvAYu
Fk8AXfeKGuOtYKxT1u/Ep2OH+bSbXSpj4rOaaSeW4jjDTkhDp2V/l1+hTo2fJCJZ
mexzoKeYecL4i8UXWrtNIQcNzARYFEQnRa2RFFw/8+NIJmG0Gb/Q5NtJ6QLK8aAU
7oXEZlKw474SlSFd4EY9HusOD8pS0ksyQ1Tnh3UJ2IN3VcW/v8Gp96YZAcLOPH/B
J/h7LquKIFkQGU5c7U/rqak8RH6TnfITFUsYp9OhaAFOAT5JHyvjArP5mH0OzMY4
rZ7JtpKTN2MYSbDy+7sl9k6qhtbT848g3ymKBnPk1moI1Bn+HJhI0e9U3IjzfBwu
ZbKlBF+6YYnxYyqqulKRnhuyBJd7OUpAlpdUYWpS6U1tUVOfkplA2lSk7RqeOo3+
g63LtizQVjoID9TtZlmC1Q3WTK9mssphpjfOJ51JngWcJYiJrj7KiBwIreEo/VIw
68c3xREQJLn9PV0XO9YO/vlClBAp2Ica6cG4+GONNhM5ATVmZ/gzqIWRtsx/I8my
IqW9AArr/dBIH4dGjL2VgVLt8qJHp/KtcjrWxqytqYq52fdG94mTWbNJZQdFql8U
/ypSfWlAzXxWiFbXqI99HVMBXpVCWJTH9nwbRWsXrFLutDh6jbTFSYuvxGiDi2pt
aA/4Ad825xpJ9zuNs6Z3ApP38E6m523Is9xsXh2Lflq4HdRQ6vrk6LWfDAfSSLtn
Gaa1wPcyJK8GtDR4Wu13cQhzU4DyMCQ0ZIxkcJCLWzx/w8yhnu0GMzQC0CmXBquH
3lKulhzxoIz7qu+k3QaTi1blcyrbKwm9xHBSaBBVsh6H0H8CpK6Za2QuLC4ktBqH
h9/GTmnQujt5SKrDdxoIpyla7F4uLY+pLmnR5J3KXdULaNncoquIOSB5yCSEk4v5
fcY3dRp50AEQmmEpotIPJy6HTSBofB0nvFn9D28VNS/nUBWTXZbvQnV4m4Se6eEH
xtPFDZTW49iH6xFdZQ4iE22q6hHoOULfo283mzibAbzwVJAlDs8hfmixUvOOil/R
92AKEYNXPH2MQnnL+Fu5zYL61Ck19G+yrbBslkKM0HJH8C5D253h8lGb7SAcyVmG
ltQJIvasnf+Tz7wVWspBxG58BWAfxddL/UmGzjLfTACayMa6M6IU+5IvlmJfv0RG
DgIvPZuQUkO8V0Lu+AUVXXxtlKPqfsJBVbooHXaq6baeyL/ycUPUUjByIwX38lEx
De98mkyQdqXQct6OLJDVRrtMF1lPoyuB84dcQh2nmAijWWpJavC9XEIo6DZ17goO
mFC5QaLsshtaEjcTo9KTHYe5H2jwaBb87paoOVjm5vr/jwSlv6aF+v+oyDmEF/as
ITv2jjsQNpHpM0ettMGgnr2aLF+JRv35+fLbrf/3GN2An8WZbfVHNmurKsXe7HGF
PUTGYZCqmABNbrll2dD74p8hCh7ocoF0oSv3hmWwp1LftLbd36Y351nk6GBXDMn9
e/PAlEgJR66V/UIT290jhY02dSJuA48PvbolFC6lw+OOeX9NCICBBpztPTV4qTf2
BVGZ7fxiZuWORcG9tI7fK+b/vkZ4kA/kInOsUYfO8pETnC1D1UVOsw33MzUrTBLN
uejim76G9jBV/UpVDhkFsRB5jsfsfad+lHuxGASLzh85GdPY8kDnzXhKD1dqholM
x5cWAMfXIIJcek5t463ih9yJDXqHXXhKU0PMdePhWfobjJtI15QoCOXA9twGvFYV
EA2VqrT91AxaFWNHfJJYEh8NIQHy57SwnZZaLbblT+hw4qWi+8u5TbqiaEnj2wZk
5kYmbZfH0+7PfqD3aPoSIwJA153t7ZQbpFhtLdhhySVOiTL0Mm04LJnaXlu93/RH
n94mHgaAE3BFpAk9TBjFKw6ySxWGzNgobG7NR41M1Or+49yxs8BhFpacCbRtfWYA
g2gcEPS8po82yQxIVvPusFz1vXJAmzGwK5Nrro9/goPT+8Ypj7zCpwKHeZxPKNlV
w7pqStuS9+UYuOangV9biI67jO80Jwz9m3B9fjLb/DNYN3EKU60rmnEV0eU9YdOl
yY6u8iwsdo2su9Jlm4iddjR0npzU7IxyaTOhqbZafxjls1/CaW6j+WJcCE6/C+ir
pHV2wAcm/PXXHvYPlXjT4v+jV27i0/bLx7eZRKNughJi8n3Mom1b9jV6yVB3tyqF
WhHzbZCg3183lHuWGAzi5K1B9Yi91aFQ3Ov7lxlFgsMSbK9MzB5JmIRpgAZsLUGc
DTWeiTAXAhnDZJzyzM74OBQ5pW62ff8RyzB+kRS2OjL1+su/00z76cWJ12Cphk0L
ZaR/TIbhdRLPvzfnca1ucsdD690K72X9Lq4T3m2RFRyUdXDaQICixtBKsAMD9Zut
GhHrEmZB3C2lytyCDBqiteDmXr0ADGavwdUmVT4xhN1wTwBeNcZBvXiHEblzPpAP
+dBVHvy1Plb2gLDtYNwqnI8AXOFB+eDD0J6rQz+zJneOpo/DfjZHF1HohUTp5Guu
hK7use4MXvOaasz7xcTbFunRkzfYcnsEzNZ8o/9h94d102dG1qQW66b8r9+zMML5
DB3tpKT2ytV004U8JTxpagGn0XI2PeOxbRRXjrRb29YUGVUWz9FI1mpj3SU11jSu
61rS8/6HOeY5KiPWcCOK8pAWWj+jyt4vxQoiFMh9NXcI3hFUiP+vgCp1LTeovaCg
TDFjRRouyskCi9CXBY4rzajkI65tTgtsdcnzMaW1qt3Nram99K9P16BPnk0oe/2X
0GJU5f+u1DnzCWQLBomy3+Zg4VY6G0VZI9xEBOq4Zp9INtg30U+bYgicH48qjVW0
yXz3p/Diup6U9m4K8M/6QVjdYc94kqOszjj/vu7Yx6MEHWERMN6Xp5viOQFT2Kwq
8tqRR5PMTaXyajjfCgr4SrSH7lLoD8wovn0E/oHMtnZyxfgJU80yFpSqnUs/Keqj
mBCM4mkzLB0f/cpcSdK7T4ZKHT5RZsr0g9h8yTjwGQIZLIOAxUczwscnunKeZCfL
o6HdvpADDMlakBz/095pyWPRZOZU2RYf3E6jVfz1VLa6k/ER6oUfHABFPI0uMgKb
FJXTcNNQMZbCnZa4Crjm/VtAFe+aULCcf40Ue0sdaKu9Wggj6QSk751KRTV+Zro7
WfOo+mvDYX5vt03ooqpdlbAyRIX9CfkFoviknn42AhXpuFDo4LyNcF+LZK1ayoHv
KZWpssfGjuaHo4V0SKB6ruTWE/1F9JjC4yj5odoqzp7UE0sI1Kn8pTvit8kXlsR2
wglJCCcC9Bk8XVArpu+ZwuuJVG5tx2vBbe4xeZxI/gBNva2eoCKfhQWMTJEbSaMc
SU+MBGMvFah4jcjbeQYP+D/gPnF29t0K30zQ/XKlAcGNaZ4Zn750aGs2No/0WugP
o0YTeQs9JulhgoC2srMzZuherhO6YvF10CY4A3bmXOfENLq7TqG4ODNmB+x64D3z
x106p8fj2RwKEDMEEy+5fC54hh04FN2zWQL9sjCAjUh7gG5RP2FgspbgIye5199G
GW4FNOrtpa4FZ4Q1KnSTBizhxAiGEs6SBxod2NagWZFIP6GPjQ4guwmLRTA8yQMf
XV9XZh/ZMAi9ihbbL+E8pw4IF7H25dSQjxyTayaFviFQ9gtjHPi+I1edcrg9gT23
oNPpDrWQQA/rbA1QGUD6ZKmZ2fxvEyTUmOQrYinGFeXvpnx2hL6q/5l+crSq9/Yg
MP+rtXw0XXbQ1+tNvRiv5dS6WrIihgB94LBAfCG3FMqCmB7DvibcjDyPQx0cHI/A
YX52DMQ+QOCQh3740Ldxef4mmjHIAiAr7ECSjrSAIoWzKKod6d0L8PxQkUsAIBcN
MLLZ83FL4v6He/gsaLYImELyJ5M644NZgAgzodvDC1/J4b69FjBxeMzb1XvCdyYK
vDXPhqbTHfnabp13gfV3w0nb4iYEn08r0fViU+8ogONOqvJ71HN/1TfJ475H1Nmp
frvZ1GqCel0Fx+jm5VhhbixrorDw0jM9r8YVPl/C+Qw65+zdyEzSMwvbBaEVfuoh
q0cCI8/YX30hE+r/neKqWLH+8FqolCddgD1JOLgUU/GSvBSokRVGdJIrp0tMtj5y
VVfJVnf+VWEmj/54//ilL+YVcJ0tWakjEYHJLKYyOBkS5viVatk6jpr6+EQHWvhV
EbZ3Wsf/qWEdvdB7GZz76pzBIA2z2PGwoew9SapiFdJSrOL/QbzzIyRaxKNLHiOk
0G/cAzfcdswWYf92/v7yMWPO2LtQVcL1eC4n5yK7qhkoAPvF4hF5F5GiXDCrVnoC
l9XEwTpjFHXElNe2IM6utBvtiVf3wpjpiKacqJXHavs1JVbzU7ay1+1Ut3vvSPIZ
8IO7au+/wOtl29Q8N+LZ98JLZT/b12dIzwPvDyNf3Dp8XGPzK3rAndMhwXL/rzWQ
p19rwSuOoHk1b2Tef0ZX8lpSgyAKJFYteJf4ifA90+4zgbsPXl2NHKE9kLvw8Ank
BICCypwqN+osPkI/vQy7Fswt03c36I/2h5Ranhqm6l1Fg14Jp7zuOk9+OcOWppZa
4kzQtlGP15RZghjWltD+stXGkpqU803UmGzlI1xG441o3NcD04tXfIg8vSnBPvMo
X2Zqv6xY2z7YnELbBw92PxN+qrRSH8lMmFo60364mWuQgx1pbsjb4cUare5T2e+L
PVxlu42zRNmWU+2v1qV3L+9lpfyrvjEYCZJntMMx2LrLfTtbCN0/qa9yWuMF8mPP
QTRwgZ8/fSpLFqykpA6EWYPPI12D9/waiQcG9DJWiEl6BWPNeK/2lF/CFMuhrPLt
paD2G4EA4X0UPEQDJw7EIWlGFzN5oalVZIEwSquNBkyBaolWWS8H68rgFjsezgMC
I/3Vr0HKGbk0DKUcydL1G6tdSxf5t8bvkWE1s0YjqYXlsGwSm8Qyl7QTHC+1WhOA
qMudd28uzZRwDJ3CrkD6LMXOb5N6H41VKHeaGxzQ8WnazbDtJ8gY+oWfMpTcx2t+
mMrk02wkX0NME8HNjVWVApKZLlsYgIhCqxZdrLWn5fB2v+SAPCN93TJ7YiZhLy4y
m/WOq7s3B5netzzCYXtb7+mAl7NFYFmaqO1FkDKSjKXYXlpe+US3lmM12dzJPf3+
Q8OJn/H0uLBfVjOO9o7ins/gI6owfFY0IG6XN4dqtw10OZ7dntre1U5fwEkbU8LE
uO08w3hLoQ8LGj6cHLbbf14R9p1p7kacZ0dBrA7FFBpBostLOquuNntv6KxRbsgd
u4jtr77BpRiHVeJ1Gap0WMdD+ku9VstoIEGHdxZXJMUvbSAUsv8NyRgT+aLb5kHM
uh6KxmWG+1e9bjlXg+c9zHVJZIMIrpoCRmKnwO+bduLkKcedZYZnW3lkAlzpOtSw
PKF5LPlj92fRfB+Kl38L6ZPd3DVZ+ZNvhAzO4kNtD4aKur72lBq6AyQY/ui5mHc9
S9/3SA0U6971fRz57jv0t2obKuoy7F2qSIaLAGl2190lzPzgI6T+wSOlgYJL53pu
CKZMmRUfKSgJy6H95Ly4U7YH+/kF3szZ1aYVBXuOghQgCPKWV4W8RqvQcwpD4s2Z
KjAiHW035NFnUMW1ff+bCTiNLNR5ftYL/LT3pNRUdrW6VvFPbncvkG16m0rG+U1v
VGYUxQtwIubVNLTQ1phjAAelvNX110TcyEKhPmduva/lhTAcYTaL2B4uVPmaI20e
4rHJrYmHYKHPG03KXERXjLDmXty5JGSYpECy5UN4dBqmufAtn2NPIVYO0zahozAF
WwN61OF63C/thjyy3x0VX0GOLj6BlMgZmd+xqRig5pwwSD/hRUvAMwpfy6EAueVl
3A4rqwCiu0I9jegNpijef7pPKuI+kFaHr35c0Ge/Rych+8wYpZZNUyPTUDAaiF/K
kylPtine3wK7cks7dJO1W2bQcVzlWIS62pYYl2p+Jq/7JTGnuT/YIik5PiOGgLOJ
eQXBaJYfLYudiCbkWYSW8dABWOHb+NNOV858O6aqXrTgnfAMm0aC/9IvTgonRocc
4PL4YAeC+FYnupakuitlQe9rsXPnjvAZY2nBw0Z3E/HhbU1KZhlE1MD1VYRlmfhA
zdSFtHg8N3JMPBnfewtthF0MdNMC0a+LonENZYRebMdwKdNvMy94eOTMMH+bkMkk
CFK/YUd8LL4/+UwqLEAKr8u21fnYg9yayV26RSigbGUngMDL1G9iiAz05Sg2knEj
ckao58dZISXYqAkQO0nCIZp1pqrOb4ZUGRYTsHPWSU1pO+UlCsSVZwfUyGGnJB8W
8vXVOJ79y3cHhhgsSnlvpVPYnDgAqiQkVI6MTT4lqQkdEW3CiCfH/QMf4J48sTQN
JTCV1XsEz6H44Wz/amPiHeOvlUODV1ANamQPlbF+3fS8q8plG4INlsvyfNMoNcd4
6OaNvcoTjq2elohr0Op89gbTSa62JQZoEWTNGdpmgUArmDQexc9b8311HpCnxP1d
fz0Qu4sJwzhabH10z/CZnRq+TQX33RQu4gJucCY2XwMZ88Ss+mYVUVTGp5rGlf6E
4uFOip8fxirHygDgFGL24PH4/KhhKvWLhaOELSi2x6WtyU+BlwbQ3KOyXQhPv39R
IGekGEamzFyx+ePI4VYW2cfi1BMQXnxoe3HNa5kSXkLjxn68OM1M+ciZlfiAGamd
SS4sXsYm95+M/h/DwDE1aAqldYEwhWHjH+ittdGNLWQsEF6aeWeDkA5/L/9jZC0r
p4usE7w4YngkrkECc1TDAhRIT6eZRhPZKSC8OXQ/qQcNrtPgdOLizQxMoIaX1xVO
u3He1vVQ2PfPZ/zLY8A3TmNyt7mZSmbMlRnqxX2zmLKak8662HzEJ4Wk5wLDAefO
5wEV4bgWlsdFAsAISvlPD28rJGLGRmYQmkv6E8IlJVMTIeY3+FoM+8YbR33lXAHf
SattYQ5XaijfC+Fc1wj7/Ww8svkXHLunlC0dgwr6JdX3p+9WHu0PLmnev0/Wma+E
KTZW4/zP63GbUQvkzlQGf6O6Spbegma0erfluE1Y51c8okYpbjzml59R4yJRkmqo
7/HQl+TkTOZqeDRFVoooi6RSf5CBucA2rVpLjv8K/u9/3QDGj1sXykahV+Cu63OF
6LAHIK7xDdsdRfIpC8xuvfr5PIMdCBp74iLscwwkqiaKTnMXVAc/++paGoGJH/hk
GV0+xIi4qr1+F10Gg87et1lgAKZnGXInKZykg0RgPur9eaO4wWLBvBXXgloKhOdQ
DDM0ZOBYsSFiPgxsXvduqgp1t7FMTnjWYvL9OqDog54LxnQxxGkX3FJrV26M70Ex
RyZqnBXsNGYx5KOlOn0th+VvOvQugDhtvyjYZHzmV+Pos2krmYm2oKFKNo4s0llt
EM9kDhVBkWtSfssWFEO09/sdrnGcdO9syOIx9PKuxk15lmEzgOUitUoaWVUR2saD
6PjnqYvqfrAT8VXJmCtAX+xrrl0YuQXs4smt1fCwaVwwtdX4fvg5MyM+1H+r00tE
Fa0HgyKfN+k0LoGgh0O49MkyuLqkNRcSef0Yzc7TEQttE7wzrI8aS5YVZZ1NO3qy
emizo57nzEIRjN60/H8gzN8qYpefEDH+fu6SR3j/yBhxd8mAlpMJ63y4jgccwfK4
1sZF0JmQHUdAp3Om9j68+R32KCxVU3+qA0Y3QE+yIrZcNOphB3Kh8EBS4ldlezA3
QS5wONf7mbVkQdacCtgOo794DuFFRYY7oEUf27umX4SnQOuBoQiPE9YtoTdVKwzn
mMfCD4Sw8XoDGfp5Xc8o5PZkc/ozl1kK7G5gie1k+CcCU5/L/QA2+QM88QT2SsTN
skn5KO8dMV/q21yWPKngWZBcTfMYd8ur2nsU+D15HCRFF8lFCAvT+/DEgfzxrM3r
aOsWLH5gDk8ZEjXoYAjtsaI1MgpbrSIS4Aw8N4csCQrhgNidY6whCZzHm35mLQZY
/bfcm47mow+1yBjGPw1INI+meuMNS8EyVMSdOli05RoHp8DP42tTQR+JVe7ac+Ze
Sih3mecO+woQ3pd31BF8R/X97Qack0B8RILh3F7XX2B4SGoPXQHlb3EFcD1pPgPb
g0ZnJFY11o7EQjYj7GrXFGATzp1ySeEMVPlIyf9D4QldRVRJeRQcNYtfgRif+pwU
dfRt1rzwn3iSBDIvFcBuqI0AuXkNFdtg6OCL3NOon5N7lkoKvSKdmP0eBwVG8e8X
Z3NL/7wFLn81gfPQ2pEowTn0chzxeDSZnk8lBq1M3mCVaee2jsjUTtaa5V99J+Ym
zDAVks0gvNjQtAaQwbALL8/Fij30/L8NB59y0QCHC11Zcgo8ETlWSuRaXOeiUiaV
S6eTnTNkbBVanw7zQIOwagWyHaSC8yGvr0MKVGd+CKpGpa7/Nkh5XVC2tW+YjEHY
iin60J5AitVy3KMyMyJtPzDfRALHRFTfR2wQ3kxUVZz3GANy9l94VwXsPqRiWD8S
xyRx9iazdqrD5BcPhofPf09nTYThzyvmaR0dFdqP0agaNjuQRQcXTF9Yh5SsTODd
nixDf9ydJKMgCVcy43Pc6W6rJb4oPvs7ycRhHvKIKhy5SOn6I3uUnJ8fMVWwAp/Y
jP7FK+23gftq1AbbN9m975Moahk74JThoWhbTx2sm1L0Dm69h2O5Wf3jeJYxhDxQ
RxZt/md0ZZ5BHj4o7FKDau8Drx/fFwqXd4p2EQOUfo1NTaHhbKE5uP4TxjYL5iPV
VDZt2BheyQeB2mTBz54+BORC+3tGmyCpuJESiSkJ+ib1YCs5ZK7kjhgbRsACOuVa
QUU4ifojPgfQ89cX1Evvs9tMOPTBJ4WW6LVG7WrhWDpbN1sDI2Qe+BkpWwnvD3QE
NyrJGeES2Y+URVtQB5Onvhdmr/ZQ33KZr66iDsJFLKXDgmDwab5/wtFTBtllyOdo
j6tLv41wev+h5XqKbVCHqDgMZaLyPDjV199bZZaTzyC2BUy2KYlv/0upt49OuKnZ
6RL3fCk4dgBnHUCeIwgG9QVV6mr19343r2lmTlHffc+gLyuU7Wxi3oEcYtWoUpMo
x+ZQRIC62JW0oo8lOwnAh1/5MBkqQnR5aPldEw3J0/WhDa/MhFKyesG0PhLGNEWC
+54qaRwmpiX5XV/POBZBrgoxosfjGD0ubu8/MPAyozOZtvNzMS00+4N1r1ZyP6RF
TPiegN3A+0howd0Po3m2zM6yLq/FaYfjukOt8pc/iZI3bUsMLXamdm7C6xsKjoMI
xiSIgxsk1+uTJPByn2b6PC6IDMR78wXyXO0qoCUI5C92Aq8/82Q5TtjC3vGnXCDB
vORKKuOIxJblqT0N+q5hBgntSVzwktCw/mZU657aV/0/aTvBoJdWtWidVH7w/kOd
coZhP634FdZ3mYhHGHjFcCalLBfr6XSLJ+e4lwW1sLVYsj+j2FleokzuCYqLD+Bi
cIrY6Vqgq4RQcJL/MrpGU1r9qgEPObBoSUqRSBSbTjDBWvVwhnIrDYNJutYZiFzN
fDgkOiCsEtKp5Hb+LsIsESLG5wSTaxtoiZZuWf72U6khAEeFlk+F31aEjtzt/Gh7
n3NZnZCeOVkH9S8cJNHNS9j/ElunzRVQqmD5eSptiZCrXOefKQR4GGoDzF1nGsIO
71KtANXqVWo7DqnSvLkafNRWL09KsmwIll45Nl9XvN2SUN44louyrBRd3l/DAOL0
sUZwtGoy95hE65QXHVU5fLMWy8WqJF+Hy/Z93hdVVNt43PmlV/9dZX3V9Vvg20u9
61x0hmCZa5YdrbymVqKN1WNKY+NthGvyopBqyEC11CBhBTGigVNLT00EJnZ7boGl
H6Os1ELVw05T7V0lgCyGhNnOmx1RBDbqjQ9JO5ZqHNOrrF0U7wXLoO4Ez8KRVJRC
Ccl+JPkQbP6I8zv5/QJyFFapqMMv2oKBJgVj4W3Dt1T+ABc+OnICaI+W2e4e9Y1W
C0ScBDx6sn0YM+BbPCjI1fKO4ZKjCdMF9QeT/XdiF/aGQTKApw7fYogmxeFIgTNV
THYUmK6LS52rK3jluZUEfI8mwAsQjEWgrqiTP+hLK4f8iodNzlQu+MzFCSkrD34V
g0PLBrUhSyL0DKrx4kHE7ZuvhlZ7+HldzllPJpWjiQrp/DfcVxAMjHo+IuholbcY
CbrYIR2IHlJhKTc8KWVzuUMWWGK9frwKsCfQh1nzJUR7Sv0KvAGZm1gsn/MtAUY4
8mp/t8Eo1HDB3OzZFgNHpunIIcvUxa34El7vrLlB2uQw/qyeghScAqkjYgGyhRdG
tmps2WUAK95qmP0ISTljaUiYzo4p6Fv4mQb7PxpqyA13gsvcTOfCLsUyN4xe/sbq
S2Vks+FWIZcgU4t7BfHfTm6zLdrqCT1ngm8a2qZAmm8dUrg+1qFEFIdXA527mNoM
ckU3A61/ktbGfU1xR7pmennv+EY37lFMZ9sagLqg6zebUEUX67hDznuRl2q4Bphy
iDiTF2jGTcBHpSXRhVhP+D0gCbX+R/nxCcKkMTVYg35AKO2tnn63HqsxzL2kQZLL
ZnpS0zaUnIVTVFTaddqwY4h9090NIoa9c4eT+5RnmIw+F7jHMhHARyaEzeOJXbM0
XpYsUr3zQ+Fpe6lRSkfyoVK2/OsZoKrhItg/l6re72kYuW/SQMPABZILC2K2MS1h
LDOmzE6gnHKsDHKhYJQ8P9Av9oiDezSTDJrmmvlk56F+Z0FaSyKOdVJgl1TPdJ53
6/VGjG/9mZFghbJLOxQL0V2D9AT1L2pC3bZOIhRrwdX3CGdrkg0dUWJQzxawFRFL
6n7PMP0VOQHl+4t0ewRApjBPGJWWxFirqRzWfipEyzLv1b5MECs8UqNJIkj0l5pa
axU5zxo+4ss6sc390C2MH3KPTn/QcN67BI4JoQG42V2ZYanD3Jpc8S3DdD3eSkyh
jibPm2PuUjF2+jCsWg9t970bOkXuo5OYvHNMA6uG2qbma3tD824Th2fsxxA5p6bV
/enfb2Me9T3yjPOP1GuDbhdPVk2CDDTbvjBga/brX/U5YyTcuUjPzx5icltHGbvj
3hO9ZOVKy6kRFhXUQXnpa7Rxieo/Kz9Osv3BLsP7BVGU+VXsZbD0yLW/0nCwDORD
Zuia+8B6BA/2lPYi6NhRUi4GlXnUnDsHD2uo47N3qSrNbacwXCJSQsBLdRu3AvZj
BNADv80YxmjdzGM7GgZ0er/Hz3zShbJFKJuoCSu2leqjLZ/SLWicElGK3AcWKltq
eTn1ufkI1vEBanAIgkYsWtLfoS86teJikw6VD+beIWBfqR1MVieaSgk+xuKr64Xe
pgCdjwtNIxTpeYYkwQdSZpFSmdepKQTP35IolymqVH9yC//4ybUZeGn5j42mfmNY
7zyIjR7fAOGfWqaSkKPZ1dwpQ8tzJPQdTkKl6OSoSBMTcRnola++5pLr/7s8FxI0
Zdx9Lbs8NsdsvD5rR+k7eWofB6p2QMwwS/o2xRe7SI4cjnN1KO8rjd2yp3fDiMzG
qwdYm8b+TzcRwIAsDC9GVJQJaxSJzhzcgCc/twuzKHoCLsUzSiLApyXGOgzO44ex
ZLTdIYot5oo7jCVuHNG78oEKvrfyVgzwG/E/aAH2+QZxCgNBvuUxuZJgWNVCTe7a
5mCkCFS9sP2dkKgpDco6ZpQlDDbY1j7tYZPw4Ea3DAzcJoHX3TVTd/SxWyqePzHE
0Gqsa1OR1kCnTmjhQsbOelcsBi1i6lY8DWxmI/RlvK7Sq41x1ZPvIuJA4/p7Fsgp
kx7wmR7152ptAxN7lqGac6RZgy/vIRxJ9LDHdL6u0wvSp7eJicFkqPMNGmgl4OYh
5CL9YXjM6Jc4r1RWFIxXgsY6JiFLKk6StWzqhnIhLTootvevxiuByHSBJEAJ3h8F
2pKeFNx3v2h/MFF7xD4j6m35Ub34Y2mZNlVYwteXBqeiuTTHkX+Po63ThO8cjVmC
5J04zQmfM1WJEMQrOa1bMb7g2tZ5I4uNfR0IUqB8azoxSY5+BGE7rikY4alqz+oF
XA2AvFRgwES5baydmUhRFSaxcJeldHVbNk4J8VXqcgt/ygV9QVL5nsyQbMyG3Eps
cRgSd2qhSXkNEzImvfpjMYoYHte9mctCmH3l8jnrAyCiH4f0pGt1nnEArbt/VBgI
oUKYNSIlweL5vn26JjahAFzZIpB4jmu9ob9cUSHEI7AEZFuEjiL+dAOWYWXQe6Yv
WmmRp/oG6WtJNu44LmYYer+0T49YMXemcWuj0wi0ZODzOb75qQ2ogwg6289b2YmZ
K5D1XG6/ytV0JBTWRzIaJ8/pRIIImOAyLTSZ3AV+/xblMpyGBIl/g4kSVUyoNakf
RST+qEZbCH4nfPuQQzXr201zbuqw8gGkzWjHgvgTsNQVKnP2NwFgYxG6vXcN6CLk
6MlfxDlV1PBDuh6UqnaZXuNI2bz9aC1E3JkxsgZTy80aTuY1/hgWl21urvWZg8Eb
E/9rxH/EADVES/85kQmcAmtrWkdZfevLdxI5FpoLK6yegWCPPS8CzooitLa4OwMk
gU0naavt0FQBa0qIE/4odSUvoXOOpyHC/VjeNNOTOf6nHRCMToHxz7dtlq3cjcT2
zae7pOeuulnj31O83EqiUCaCFxK+7+ym6x7d54QIyYPUlEQYlh8n3X3LHoFaibzZ
l2qCMSAnG2uAhO+d46pGuN6JMgqyQevx3n60ufPGGsRLUZmRRIvPbowDixc8L/FO
NZRiSbhA35CtP3ze0mc7lChOYNd23un384T7Da/pjwbjQDVn/Fs9e4AVgKxqKZ8q
PowOS2hFOWwgYW5qCpoK+3YxveiyVG5a5zU2fBSukWR4EbQApan0910s30Ui+Sdg
cF/s7CIe4gPm/Ybr9xG7qVg/Wr7xDru8uIfxxLeJB+EG/q62HcpbADUNRtFwJYxm
3zIEvcCFyQZUB1i9Q3tv2X9pBQnWNx7S5s5cvimRSvMTetU8O0lVZ7VlcBvzZEga
JtUTOJ+BnkjNKzrDcsc1EwrpLHR4bB/n3AI+SowKSHvG9jzSt84qu6beGsFzmd23
wbKTdqJl3mgWDyZCeFzakBLdsk9igc3XpuyEvNlYT4KXoO3ZZFpqvg9Avp8spq6W
3PNxLTu3JkucfVEX4zSH5xT8y1kzw0odfainpanlWdJmSV+WF+QpieaQ6qRfAlQq
jzUn//mmZE/3evcqXMiafbl5Y/er6E8qoP+KKVNedTk19OjbMyGYAhH2pla+6mDJ
53T/aFmAqbVxYSwk3FuaGZvfiaw2lDCrr8OzrlJLMsv5wHoF79vxf398hbrz2iTG
uvbJOE+SOwzJNR2sYInJnH9wAfsiNp44gyzXl0XUtOY4yVf/lZeMpZi1BSlVnpuH
U6yIPiniNRwWDcYv5smv19/7LTTT8JrgBUX8e+begVj8D3KR63eSv1fHI8vvuRMG
NFHGlu67JSLRwwxM7RIzy7AqH+U20MpK3lXKDHZsGeUpjeT5H1P2V109hg8Udgfn
uCT8OXd/WAKulwtYdOZkacpBznRHz08Li+CBSif2pfEs7hOpA0GeYfwEx/hgxdJ2
XxpFy+k3h3ZPqgIWpbedYv3uckDmgAWuUwCIQiAbG1sLZuc2N0QvCN2kUlY0nblf
al3mdjzxIqQMiZi98kQoc73zKEvTaU9zSItdtuxGXJzmA7pgbzdxGwsWkohxNZlj
a69n2UaOyOds5qIu1T5YqB5xm4SGsC0tEzymIuAu3UyejXy4h3R31IYd0gYjNbWk
tiPj6U+bc2uJsxpLr7jr0wmkOH6H2FodHc3BDWF4b+4qlw3ElA5Kq7IbKLXzK8B8
ulTaVXirpbr4uBzbmcAyzHIjifE3DFnR/5wqB+jxWuZ2nMWTOtyBFzOE2s/24B5b
gJXbhLp7hTqs8CC6Z7xzvLDyi3OmIvaMjmrSGy917nclT8bT8OQdHcZbeawGO096
jWsAqkjM4b1FXcpU3AtphkXqxrJXA1yA0LR5RASI01MLPrRQVgTf9dnBX0MvhB6z
MQ7o0SQQtq54EGdPO4mEYB/g5FkUFgrXux/O1NeZ2mduHC6UDOF0HSi2wY3uTEyK
cP2pxrKEz3Cug/yvxz6GH0JP37vStXp6rVB6PRyJC7SfJqckkwzluOY+MQ6j89b+
zTwgybrKpSNR1JS89P6PXiUQCByT8yVrZsZdAxGwQMP2vtWbtL4L0IP3fmMXq1Bd
VVWEU+Wksw63pr4bH/5o8Z7N4k69HS56imCgEU3aFXOUsQOvat3lUbX5KwFv3Teh
H/+bS3K5mZWZbNdpXso3wM/B8ypjQGu2MJqBGgJtVe0HomPBXZdcKY3qE3rxZPMa
0F7w0I1dG2Ih+AIZYHjCtPVoMPWXgEZc50+jRE4IVgbC8u6qh5IDap+rkZSIsVhb
QQyhLsAqQW7UnzEku/PiNXYM2w/rvTNQyT70/gd3sUUfhHuBIg5ktlvZ/efGvIUy
mLKIT6mPfOXuO2YzBM3SBRyb13AXhU0hD9VSKnvl4nCNrn+5a5tMEQvYyEOva/xr
pT7rHfy8VoydUqZLazlKVsNuwUm2dLV3fI39crDOihHQH/z/H7CkUGYDLgP6GuoC
vVaO7otJkC9oP55HGTXXvd0OtAauwvsWjBREuYvPZQgbyOOECtTMZpB7dyFgDfgf
3u6KkFYFaSjnRRgu+fXW4HYAdUUzLM0oesiqC9rhLy24CHAxeMxczZNe5nN2IPz+
QOYs6xlsHc7ej29W8j4pAwXpc6+PWIRvX+fraKjonJuJmSV3Om8eisG+WL0uVTpr
QOnQhcY9oifzOqrjV3a566rw3wU+TvSv4SATWkalPpsUWPCM0OMITETLEjt3Ldrs
w0tO5bG4Txdrbb5/G66rXm97BhYwlOFZxZ8TyAAhFmySmDWQ6doV+3AIdxeq6oiY
ZTCuT4llFyqEMakeJEk1yomMZRutiDiWRSz3Be9OoRYcI2riGCXDwATeuZY5DCg/
5iHE6Z/6Zztyn5Rd15HgzPNFLDN3Mv6Ur3DbdQQyc0O80FDKxRDVaLgMWmZjNWy1
MeLc/Qrt/XI94r9LEbltfZiU77YCz4ckwi2B9g9yAr+pDyiVKEH9ZAaHolfnIqQz
zGN442M0toerfJ8HAKP5RAjFfk7VPZM++cpC3Mgp7p8KKHiFCwIfxvPdoWG8obGa
Z9FZmuoyJhsHdXaKD/gGWOT8VuXwr5qdL/z0LlvLyl/zCNVJ1pm8IndedxIP60qP
XyCM9YeAoOKQoSv0U1vWwSW7gf+TezZ0DJGhUbjvnEaYzm+7Mvf9wlRATOY1Li7b
EY67+kDOWjX4M9t0Ax19WJdIZLTcFV3mP3YoOuqmZ5NtCnNa+NVP86vAVrwtMqnu
GTErM+xnxoEELJ5Ee4an/ZpkVLshyAQNuAULUk1p/Wb9k1BSr5yh6MfH7C5+rqpS
L3UkOe3G3/fZaGeMTeXBIXMmmQMJwIAn0oxnsly74rFuBzmI7EdnvRYKt6vn39Tz
NENf/CwZamtbJvta85XcEtg8JwXrAHy9/oe9oFkIeqSP+w1zH8RnxkchrUQ4b3z1
iIEXvJdumqjr6LH7aGszh4Lw2+P1nTCob3/E81Gb82G6SeDOkHN+U8O934rkaS/u
9QkoKl6G1bR4+cOLET0RzU9iGnScZqYeHLSTXGdiiCDwWaac18xunUepgX6jI9vy
fW2a3bjwBMfzoxwhO45y0lgX1aUIEuGO8SXfPGwyFuhwXGsrrKwcOFkkqOtmNbnj
soWr5iIbWNjWZ8dWywlMfoL9jxxIuEaBabysX4Rac4Y8E9u8fkMX5Jcr68xPhNbF
3bZFPm34jUvIjWKcYlHdcosfsleweSnP60icwFeVacHNluVCGCtjff4/8cehchlD
XZ5whHjbxzAHCZ9QTkAZnN6b7kR+vBF3c6tQ+bmXhykU0M2KROCxyZ/yJSJDjGjJ
PNTeT3Mo7BuWqu63sPnih4ufkS0fd1rRSdmhLqVQHm9NwLl+w18rHSZm8/643qZP
tiCqsgfSZ99PmRR1y8XfefWPJm4NEFP2gkxeAFQ/XurHuZqyT/cxatxLjKZFBM7+
wtSj8GffvPBhXkVtToRxJdpQhbcRY9H5ATJAKFz/3DMmid2i9m9Nm/2TnVGE1aVe
ZT+I9psvi/PWBTLUKwaCb6qxIxu+GkaTn2pZhPGENoRHRE/zvu+j5If/81vfrn49
f/ZFa7HxDUEnOgw/dlo+mvnUNqhDMtGvLwte1RreiVpm7BtZlRnsJE5K0y+JxUnF
qQ8PmGj9FocSsByJep0AylcKY4/uNhZWTIXyOYRkvJBicIzJ7XI9MMFRgTGDd2E4
puRvotCSrDFWzZkTXoUlkJYDczfA9mV5D8XAjF1dnnEhnpyH1iXmsJYfbN7o8RQJ
csGtfm9ntsZDxY2mro4rSrgkOytxqaul/gmmZog507oiPwGo/Ea2aDp1SqTQ8/9g
GYHlrVXpeIVHEKlAaME3p3lXkh2KXCjEMljGPKgintmPCxsf9cKUgGUJVNGRGIke
h26Ze5VS1kF3w8P9nFUhktOfxZv68rsnyWivE1I4quftLFhdDLa5cDa58W3beE7b
a7NOpAc0HbbklNKS8+yystb4TxUftgvjb6LS9ZxYZvajMrgA0zmDBPoGl0fVcV1X
q+Fgmb9ZKsMC0uhiOcJBcpzpC+TTltXRw6W7tIwzZw0FBFqm+SXEWtdoHeFmWT5X
g5lpGdS8oyGH5pDMDwcxphoDqXR9P77x0TXyVhdhUv6SUbtP2/4R2Yuvb/lK2F6s
FhXTk+9aUmey1kkDdw5+5KnFLCf4rEB+0ZCuyDz2avMEq3RBW/04/kmh/qraP3YQ
J4NcEUCQsDuvhzAQl8wEmNa3OwbxuyqB/Jqz3s8gZNvGrMNAqqf6Fjy+9fxm6WcU
05duUnT8rvt8fTTl6mwtbutNfTPb86pE7a8hI2W0hX1ZeYpJg8UIbgg9q+Ks+Fb3
Xb10yFbPWpUMa3GzioiIUN+MTkVg7keZ3KOIzhiKRCMur42totTfJ64jLkGuWPyq
ttwoIKYxrFOYtOdPLN4WFuBgM8NCUJo977eQb6kH/A5R/42uqfVbJAtnELKF3nz7
4lAUCZwa50NKPwXQ/RNnNZDnhgoFhDi9oOMqvHrqoFL0ut45jZJXeXmjG1lfpT+X
IhCpI/YiRLjYbkVa0eizjAaK4wTSVgvrPTqI1pZu4P1/u3GXPEpYQi7rMpae0MZr
Q/AT/d12Wy0u5RNJKqrwkWXIPe8sWpK/vzsvar3sPp9gMWU3X9JV590xO1KiLOZF
lt0feFE2O8jZE71Ax65V3RUZnOKsSUsESPC1K5Dj0d9VDgZD6TErtlBxzXhLtmWX
20w9+m9fiZstgVVhYWMggpvt76OpZS5rVJ6MrizUMoj33EF2Erhej+Qg4GtZNURg
osDxp1KkgRER/H9//DxZhfjJGaDyteYhgGLJUdL5H8Cfca7X5KZ11oDb5LcQ0jB5
GQp/Und8JwytZvhXNBZ/TUoEM3IfTqwcciHJebt8+j4Y+I26c7vkOHNVdZ2iyStP
CQsmKPcFcbxPhHLWd8yuHQfT6GPNfDopI4GshVUgGPJ90pMNvRVyPOdTDDxiySYc
UUTGd8JuegHP6AWXPP6ir+VSIxPo9dGAQtoki2qfn45XBClD4NnJofoN4usnfbdZ
6xKT3vFYQ0sc7kBUiVtcpPSj+GNTi7kpbwp0oYCyHS8PifvioTovwZEmV5yzoIUL
XWbR99SxgNztHrQDbG0jABCGJAvlYVMLpZEWPI3jJpx41ckp0Mv3BTe/avqySb3R
Rr3SoDPzV2ccXuYJIPJSTb4RFDZsYh3+1xPt4IMltPrscn7syn7b2C48l9Hve1A3
lFzVBmgiCXnsYP0QtX52BYge6Nwr8y3FkhA6oYJW54p0ZYM7XAQEhwxmxWGlezQN
5YfSCpqY4cPQ9QDt71IuCyBtEEBoOKUWAcTtYoeKgY105R2Gq4T5XPVuu8bCaTh6
BJn+fVBhbOczDK4cuoBhFZlgU632knPwqwSwVMnzWaSr0S5GMvGSkaVOq4PfS8lU
Bwb6h3OTubZajKPAAr7buqlKBswTpb+56IabeZo5TBo6qmU5Qaua++kr7y/xmqxE
PbynECbpG1JY6k7Wo4hvQt4dMLKBi0bIq0fYXaK3hLByi2mdjJsgtfkSv1n6Fp3o
bZ2gu/GSDpUWg1kUc+TdMYejMJbii4BrGitExJuTOxjsFtBuMyPSmNi5VQSOsEB5
Ln3eR0dAmKF6lSuvHvjC3rf2hGTqKF7mWfGRJZ9HL3MekX7IIe+Ebi8EqSz7D39s
owciGo61TUlMWnxlyWikTRaGJp8lGmkSS74A15O7fqSzxy4Yqo0OyVNUNbfpR5kh
H+H2KjhLqnnL3POV9c4dZ6IZOAoLjmeVKV2ac/QzE16cPuZ9wZpk2nsVVzsjirWp
nXYECGWRqMcFYwILgV+Jo3Mjen6SHiShsBBz9uVEyXzhC5hMX6KMT+5btNdjOGYn
Oe0AjD8BCH3VnNg2P78KQdt9ftN7jPeyJ32BScATJImO18HlK61l3h2nB2zNkvW6
q4/NE41ldxfbLMxqp+BvLln/jzpVLtWQTnVpbd1IOE+84SXU1ewVYyKUY7S6NjZF
MfcFfbBiI9I1gD+zGe6a8C7a5xeIXWAU0OAz0ficvyeWWr7/RwSSLPN4rhetOe7s
Ql5GTquJ/TbRsGAhUQwPCOOA60RBTh/jjGfCowVx8fhR8r5fbusSjxPgJt5e4E7M
7HUlnAhatry9Y9epP8fA2sBi2WFw8J5qlfyGdrDVJhjOris2zLekAxMJBE2QTeO2
0KaLUDhvzXc8TSYLGel7UnqWQ6H/pIRHZCxQYe4FaHvJwfNjJFAmC3m6dYALI2Rx
z0SKJClC0CI0J0lJesQR4A+PcHZCy8mUK/7M+otyNzARgHRzvrJvuQy6dV8QrCgI
b6Cxyn8zmaoR+DJhBZGJVNbCURlV8mEy2JI2WSnsDC+PJnhwX3DgCws9t5u7FAIP
wmVEl9yUpeLk9tBnlXLxFxlDjH8wKyeLtkmvSnhsv6Ipuiw3wGQpRLuYfr1obrzJ
z8EdRCewVBgfPK316tuJss1bPqUfaGzLRImwDP1shwNoMkYlmpyL8nPJ2W2nMZqx
6yaa6I944cUGCZ2kNDy7UIGeai4S93s7YTVGfVltfwRmzYi6wDSbzox7L5KuXh/F
JQ4EJ3d8ex93nXDZIVhS1PbaHmMk9CcKfGmKubVRdhoxOrNkQhpUzYh9slh+SsXi
wfnvgNG9ITzVrXUHV2f4QQw7Gb0XVs29YzIzeJSGymzmfvzY1A9mQ+7nUOBnoQnd
pCuYQxFThndqYyL199mwFZexd/Yy3joEVBk0p01OAsMrLnQkhPA4adh5njtyAeL1
BSwFOAWI49nTVFfYGHaOuKEKaayEmq6dqujuOGvPVUVeFBHViI6LeQmfQxepm/gM
Q/LcYOoRl6cpZIdGfs3iVuX8rZVFkmgzruJmpv7Q0KNxLmXK8rqoSGyME4/via5g
MyFlPvF59uLD9spLPO0JP3foOehi4C8kyYfJUkv48trAHqFmQA45sFjzkqkEgCja
k+kd6iL42cWZ2iB6eReCefiJFHsoOrxkTDY4krKQ3rdixyEOYh0J6sHrLnmSqPh+
zArDk/TVKsKBJecrHGIV+q5fW4xrHCMMrqpqdjP4rE0MYQtXYo2UUqglNz37mks0
iOPDfWcEQsfEjxR0zHk/3X48HQLlOwScCfJ19NVLG7Z/tXLA6z58FsdIlaAKCzYX
nlZzmVhCniSVNZ0JDBQ4A935yfunP36k7VFjqYWqOHXdqwhBl1aFN6fQ+Lvb5e3T
MU/7oHd29hDn5lXDrh2XoBUOR9k59kTB4tj8VnFJD6gEVhRj6p/eGK05JdXrRdJ1
ktdhdzdVMWySzVCXuWOYJ9TS+S01I0RBp8BVnihMrWvYMjlCzqkdSP6obH7M7U7z
oAfOA6hchYouBLo2IAAqftYv5hWW1zilddVtuS8J1Or/ruV0yJOKHMBouEpkzkOD
d1F+qxsXO3uPJ/hePPLyzYBhjJ73oZbGb8DWgUlxHvUGupqXltw53NULD/Vj61nd
1+xdCuDBuK1Rqm0ZXBAMqg4XvsXaac9Ddk2cQZ5ANz56UciSmAO9QdE8/oFuol8w
6uQ4qqNdcht7hgurgpHHNd+ZKL58cOHMt07PCgSrjiRPY6txogwG28LuYDyK4gZw
bLFKd0RgzlrER91OKARtXxkFuaMcjDsOQpzAnRTP08VK6pLbS8J5qi0uxjQ+HZUM
Nj1RD3Ux6cmpVGHO+dfCf4AqYx9Xot2c/fgXKFxMXWSfZNM2X/4uRwYnmkFh0KOg
yM4mPIOk6+bT9T2nqG6B1yoHWr3AAgWqK3ea94aG1u52Fz+H3heMnOb5K4Kw13FV
yos1Ed90i6qGBcJ+T8bhDPdcB2oKmCl78Evk1egsj63Mt6sllz1c48hptnicUVgk
uKcGxb3YcJNsfHpjzT4Fg4pFqCRnXZjmys3swgsdG0tQpdoclFDRd8yNQeCvPS6w
di7S1i/qjEtLdbkN0/ySi/SI6dg5sDYKKQf+4qPb4hd3DbO6bo7X05szFLHmUGwn
5+hhu8Vv0YtRdyBPKpUrwTfgMDbJQeqWfFaUyrFDzTHTAt0pYHw9/JMNUr8mCqab
5bXDvgUkVsj6HZ8L8QF2smwV2/r7bvOTwmLB3PWLC40u14wM3zW85cxq6ztKPThZ
4jhf0y5Ia2ffaS3hLMlWvm5JY7kLSlDiL/enDJuhA06vYjzGSPEmmQylAGuic84Q
35j/pA4tgzC7gxr4wpt0ZqoqAMjU9QO5uKrIC2mjkzBXGb50C38JlWfEFDNYguxA
ID99DnNJMZn2PE9fPV9sLBzTx21RaMV+90sYaTbEGFg6K1M+qZyzREWVSqlYCL1v
uGNnlsV24w4DDSIel3WOw9z4SfoIS13ygQvlWZ8MaKSswkRc9BsUTO5toHV5Bl++
oQnq4F+aFKoden+trqMtMjBmt08tsDX+RczbmUiLSU1L31HxtPiEsGefJ7Uw1h4H
mjB4V8I9LN4f/BCuRUOidGctU9ChMhYbiICp+alDIED4Urturcu/x14O9qRlye/H
KPJaOrvo6ooUbem1vltDPnp/c9aHNqn91g5P5b/7dh/rp/Mur1Bo1KkCxIwZC0B3
MUGVxrvXvIAt597eYSe+FFPqE2lMH2scVLHNtzV+JPn7jEzEPHJEVC0FEvksx5A1
kiioQzeTIKnvO4ZyUjyis42LoVRGFZGZDBQZsx7By0yWXEJqPu29dPYooXApNNQS
s10UfP4K+lCWaTzixc7exASGm7KOkssPfXX1/Mwnpfldt6J3id+whIL1HMBCdFjh
FC/RgZxFzfJKgXaQrcvkR1yBnmrXQhvyh81NSYqQ9C9eW3uXZ7ptDeO+yntAI+NA
V2X/2g5TbNYNu1lbgZ8hwQWF0DWDr+2UCpnFpTwEKXxrTjsRm5cz28Q6BRnci38q
7yehhMHNM4QYozf5z1k04GCgjHXpRrdfRdYCunkJhmsjBjx3wKRvOtQaD+E4CIKt
WcgXKoD4Hay24hCyCpcJfcaCsZcA0TGik7keQoP6VadutyfXinrnQokTwBkJ6aN+
O7ikkwpHrW+lsdThCmVVSLUUjKJC0lG7hi0vQ1+iO2nRj+d09ptPfJossVbsaQUA
xXYHv1DUvD/8NsE+8nLo+udmE58kWzjDDTyCaC6n/+WyAbUo9f0Gfb1+Ee5NFBp2
gfBwBbZteIYTXSDpZ3qQmBi/29FA7nHfV9G0JPCrKFVwSrdmqivGHoYyNZ4QEhDV
L6r7kYmjNju/Sh61nijshPbMlEJKB19idCqLddiPV3r5gY5v+/c+qsKjfjzAbWcI
9ZZy6tsJZ3TGxfgVfl2DYBo/9GQUMo2NqIDIHft/qSvl5GpiVAJhRjsmPa38wBA4
8p3RHiII1XyRHyLwbKgF1WtysnzueRZmwfzMBx17q1xSnTMEE6RK+f6AMvUOCOG7
jHh254i8j/P0DKrXeFyadtAPLypM372Chd+vRUCQd/MDBtjBKCelwuAqAwamVTee
k8x1n44ZuBrmDuYPm8LQXHuR61QZSChqlRDHv8TWPC7ynQXuo6dSODK0rv2RAOio
zWAX4Di5b96Z8RPgdAQ/T8dyOkx5VSodjwjTkcetRNDLEXy9c2dV/9sAkbig2vfD
eHSFueD2ei3y8mj3DfJAnjTR4w99yq9kwgs5ZTHEna+h4XNCTIajwngu2LShIptt
6hB8rw7qbUXNaZrwAgEZ2+aofOV5KgMhDCOAMFRWXHxBsitVg16QHbYwrrZigS3j
NTfNw3iwasBiQNvHnYa2IRKiO4yETtKuT6T/rat5YxtYloPBd4IMCh/k0rmpmpce
pPD//L8NsVYgI1p6RAzX8YDxZivsWvmY/iCE0trDAApBR4zY76soRzX7IZw5Sm/x
AwoIzrtqJpH7OSZWfcCoIdSjo1/+V4nbDTYcM8FYyKEayL99KT8RSggv3aD9eIre
fqUVqQuH+FGTgIR6tTH6VDghTV6YC7XwgqnhWDBl0UoI9ykFDMJ7cjCis+dqVlm3
srPWYkLRfLO7AGhZE9f3dibRFixbsbrxw4tZhBWoxrLB00KbljtR0mNW7Kkyos2V
a8GfqsTxDchDkkrtDLUapy5NhlVoQX98qE7I0MkPKphH0LxKtuhciuWfqFRzldpP
xvnMiU51x4tQgsURHL1ZviPv8/x2uzb96GQ0E6DiOc6A9Xj1RHJ95/jld47owrg0
yeGrrhaC4UWOW7qDrkpb1lWm4t7gE3WrhppKvMNf5YN/BlKqfE149kUwWKNXI0YT
rCS7/Zxw5aA7SQFO5yIz0OqbL5uFzLKQ+V6YUs3269g1dkTUWvvhB0mdO4qg/XJk
7oFeLrAWqnvbJ+erXlMkkhS+Uz9C5sAFQOO6A6j4YuGbBfZlpkstsetU100uCVOK
CIJXPbUvLgMk07a/Igwgj2ofZBxg9P7FVSmWXkw/dinI0N7EiBQgCPez3Cbm5PPv
Lmt0xJ7OP9j88hraDWMkkGID1Lq1lrzK/mFMdyqwsQQzExmWns/FsobzQtsGBbX+
WihpsiPEPS9lw6sN8IxU3gkFYdxuaWyJL2SM7wmOoHdzg2LiqJljG5cZ6EwFu7my
ey4ddfmgYrVtKYYu8l7d3RkzHD7zUVjvn90m/ymfEmEujpQ81Jr42wa/OusDJ/Os
V7IXfUWt5zYJhN/I6WuvU3R5qBzM6UGikXjk0zJsHKlIXj9nV+VlEZlCmmksg2Nf
+4dH6D/on1at1kFpdp+SVceuX7ghsFBH2JuDyqULddk9hFItg0WMeuyy3bkKHYjQ
L2BGzqO0Zs8chE8TmawL/A0hPSkw6YqHhccJpZLbhZmQ8lQEjEH8spkUOvyJ95ig
li1lNXW9TgFoM3dxoU0AQcdVIDj0WFtzyTnGhJpbj7xA+AkpK/JaBC3g5BX1RL08
JQyFiLk1xDHBfmaonaf8rw3laz62C5rDymQ/0VVzhM1V4JqgrqloKzNmk76GHfbN
2JtVOEEGBvj+NK6gvv2dRuANgCGKCPK5UUzrR1P0V9k0bXJTRum3oQ9qoIkBAkzG
JK4oOeTVV0//z2Us8kVLm2apB2IImp1Fu4zmzbnxOvd4u4/IjRtk85E+uZXH7Bu6

`pragma protect end_protected
