// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
L2xouLi18Px2NS8QLAeXdpJi5wIGjiIzS7+jTaL1sYVKMVBR+QvgmmAZzmPsANN9
4zd5Cj8dEzUuiyyimrn9Y4RZfxXJIamXdISYILkPZ1YZeZc2HYBFaIomtUrA7G32
oExoOtsEfAdYIHycB3NS9CEL3gZpX1JuYb2NkNw8dmU=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 57664 )
`pragma protect data_block
xg/nIYG97j2XVtL272uL2P+W9IK4881n3+7DTnIJTm6rI9KNvZ1ZRI+Wd+6yv5CE
SdZe51whlRb76Y19oth25qtaAFc9qoX2Gy52m7hJsaijm1/CxwDqFvOq/oWB7oUa
5pSMO6eowh2UxnyESgcN2U4plsaKf0QqSag3Y/DwbHV3XV9yd5Di+3Jvfl8j1kJI
WmLSLLy9Sqf6ptGE9ocQHUH8V2JWcHLYfEOZ3bXkso6kAI9o3oniEPwAklFAJvhy
ut6dFFTnGwjntrxbQD0mL5yMkKbK65XnwGKk/JYS/wUShkOZ1Ey5Z+YM/o27RomG
+a6JToRC0cWTVPJOFQaK4Z07jCAYpu/5pBbGMb+rvrlItsguQCs7evUaM9B7bDJr
uoMTHMtZS5eua4WKi8J7GgDzChEGT6WPvtEgiEPtVBpS30Poa9WBbV3ysOfs5pK4
lNtb1XyKscK6UBpqbtHy3GmfeR+yAbrudP5Rs3OyafEjYC8rdqc6znxW657W5HpM
fs+wF3vRDabrWnSPWMFIzlZl7jtMGs+pyZ55vStlqsFkROwE8JmTgJzNtADGMuCX
mtvXXKJGOBnwq2LJ28LbFG+Mg5vl/28XJ1yKyLKEK17Z30zuWJ5itnUl11ulggrp
+4sE/xT+apWhKpsoPjMtQ0iH44mY3ovCI19sKeNUKKx386xUhdGhKn7bWjyutqON
uXcNoSOTT2TctzDDVMObAnnXpMRZSUnDrN+YdLh3l3nZaHeEm/X7IFMhZCnGqJui
MEWai56BdaEUFUvDik5m12uLCWa9n1gnJdABpyu+NWmb0KoNvomJodDDtn1a22w6
eGRTkv76iN3ptULwEKfAaBNYuEpMvGap8R2TNIjnnSqAlOESLFre9XM+NAFT9ABe
IkNMCnFrWkxasETxuafKHh9EaRHn9icOACxvJ88Y1Iciz+inhemQETW0dfgjX/6U
vvSd4wugdceAAcQEy7wIKRSaeaCoSdpVTevC3To+5497YnaM4HPfEh3KEzQZd5AM
IR2gNDarm2FdUNgjGGhVnvRIHgvWD+fmBnqh83TkkapHgdYJjWWdr3utGZ8AxbNn
HhthOmIp8FK6JR48c/3r79mhkQt75JNSuF++f22u2/zyVLf1k6RWlDmVPDhFkLVI
t/gEXzPDRQ73d8kP7CM7tJC0WKKwer45gqDqlTbP8a1YRwJr0gzZcuvVeeASH77f
hD4kD14RkEwWR1P5ALVuUK8eLJ1qi0sLgFq0I2UPuOtSLxh0+GfDQtj22u0MgV2P
AnTFtZQDMMvw5cd243kCcMmJz4CUSX2FyZjkr2pJMj8sH1ez3bWN11fyQ8A0b1dF
2VLzHdC3DQGVl4aRQkc0LHblS8ufoFSlpoAUv5PJfK0jv1ZKcRhup4jQVctbr05w
hxBxAZsPIcRfaLuPveaCF6h4Dpgq1wzhpeizgYlaCoA5sl4zhrqaJtrH1tK8o1g0
q3e0c5uobYPwkPFJleK9F8LffIHrnkfPML+gv6axaXxID+7U+DqrKIbvRp27+2hV
/3K6iXIFfDkDVeQfJ94jfqXLgaPrrLqDx6Tj+qVj8FR9XSVCHWuN5D4ROAnyWQKN
El0ZqF450jr5pYAZC1RmmoruRmOI21L7nKAlX8/GonYvno+XGPYsBWSUsBoduEZX
aEmgkjQ2gR6rqDc/cV3n0H26ITfktVZVrNpAlGIEZeIFblUoXwoLDM4iq4zz/gJo
wrYUrzaO5JduqrAHTb0HvN3wkXNQawFv9X4WRmgYd8WQARTBLx9vQgLdOcWkNEAn
sP1MhsixO7Nh9wTrOBi5xa+js8CM3sckj4xO0t9dDTnbIx/KFWAYM72lfovQ6TJL
hl+8Y6nw6d4Q9hmt6vAUeZ/W4F11NqGXQ43bwqXU7UWI1LyhAOs2QRFGhcB34p7H
HQ+CmNrRgI2WB/F2TfwOKwPTF0wXaaHE9844+WVs+N5opXiUJ2tyRMlJD6mUriN2
3Th7LQaebtDRskyjOvr4X00yCZpt/GWrkeic5LjzhAPvPcge9h9Sggmrj/egedLY
64ONTduoQvxfqkhc0blfwH0md4qdIW2BLUkM7Wif/sJH5uA/lH4RVFt9qcQbTKr1
fA5+WMyeo/1+7X+KPQ+AncXazKUGuV6P+M8pWD7vLGHbd6D7jJdmZtZxOAMowfpB
5aPyxjYTrahD+En6MrW9mIc3JjTIKO/hUI78da1epibrg2QYhLTlVdpuG10yUcu4
hSr+s0W2zHW3wrMFru29NMqaztnsnJdBdWDfKmBp8KwABgVQ+h/zjjZXgbIgGHFd
FOKwmd3SSPWGDdfWW6BlJjEvhDq2KWjLj9srRNFQbFPv2djlod5JNJ7Z49k99iTu
0godwlMUcBVnV972ttQQPm+L6PIJrDNHdphwthNdnKVJR/UYHpTtOtwCR5PUR1DW
dSvFR1ifhQ0P41ekIGiLvua6hz/HGSirqdBM8a10p7My2ILkszfqMOJ+766W1wui
qpeus+XrBGfjSFSiXqvebYkrpkkUfSPCvZcLu/lczQod7ai6l4xw0tkL94eZq1jy
RzXeoI16kPEHpRgApovZq3ckWVxyUxM4MXzDFytoVR4JybsrQDhniIevGnwlm0Le
KuXDzXgVUhn5iH905RG63PDhBg6x3DA3F/CHUIGoyvUM92i8I3FffXU2jELgjQq5
sNu9WULVyirr5+cowLceOoqczM/fLfmkJazIlz0wsMlUI7Lw+r+6/qhJPE41VcTY
OUlYWMixdoznV4rlHThM37Gar1lpdJtD1u/C3TyiqTvLAT9i8sx+pm4KLmfw7P6r
UrSZqRAgFKYjeYlqrqhIw3PVeFvmV/HYPJyfvPmyG+X5f+JCg/tHU7++LhDE8/wc
eSr5d2fCVxm7Y+JCF+ePbd/rxAFFlK42Toub8J/rJjbUtEFgWuejjFHeIpBa8qYh
tXYSzpYjOCJuZU8lWHIKiUBiKxYXLtKvrGJcnsmjd4TIFH0hGUQF1jK+WvYpStst
1GSlzO8Y9Y9mMan+O0+yl+4XybSwWKF6SbyX+bSWASmepJTjkYyXPtRKOMPQK6KP
0JpJww133MLPe3ZcGUQrAR9PBASruk2aIsqA1+/bm5knlp+L8zpo6fxgZM4pmv/L
TnwvLXZr6utixEwkRHJjBTdIr0Qtn7A5IquCm94NGNgwZADUrV4vIC51nUrPmlCe
wzjgXeeeypXImOazZcioPDQgb8MBWCXm2bhiiPIhT8f4aRtoNkzntWNHqeQ6UP5l
Irqr37S/99VOEDzh/EUbEKm5v+4L7lj15MDgCLV8zhuCVytHPspXGpxgj0bRytwB
7yr3+MVKLDi7fD8FXUXXpVsQMdUFR7CQLnfCVwQf/mzu2K9VhDCBaJAP0USv0Iad
H7yTmvEM6rXb2r/Pw9g2RXklGZG8PeOAiFE3OFQbnsuWNlKAlGObKGbvOjqO68OI
m5NH5K1y37NjRCgfZkDHjAmozBTHNqPwDmJidp6F0j1StXUuS60+8ArnoDfP2cp8
1yV6p+Ur/sD7Dlxq3khFPrlHo71HSKUbu/3wipKT4yY3aGnn/Whh86YZ92LfmPZx
fv2TiHyiVNfdI04kfdhDHoRbmeO57qVdM5QAYoqra8mkH6i6yAFjgaqJqIEFGBzv
klgPcOgWAjqA4YYMpWpfxmuhYgaGXNLRQBMYk7QebPm6u0WGQD8lRed+TZZiahiW
k8WZWfUj5bdrg5qOBZ0mQx2og+XotrrFMIzog5jUZBbKtTPCi7OBE/fQHQDWUyHq
1UiiQrxfgWV9wutxJB0zjlduuDyIYDs/q4I6WEuJfXX9fI4jn44QKc1oRwKy/rMa
0qsbEeDfnHq+rSkqwsD0C/55c7OBeZwiE+lWYPJOeogfLqrksWc1klDQtox/bAge
1OTVNKNmS21snBUUYsYgWDlJuE/XamcwgK5rh4g1LHIu5f+ZLW5SNPc6yFHhDUV4
bfoVH60EgvdszM2jOzl4dZ/vO/M1kpS5JhzvM6nG5SZ5PAdMrOtnuig7L3c3I3pG
nQhYYCiec/OI00bq4oJkkcxQQExEz7d+ZNFIl+QclAaOW9GBu3dmBb2CDd4VGehw
3KGmQlzeJoyCoHBiFrSqPVq3ERcUrQDivAyQ/oN5fHeq9OTUelnHZ9fHcv4TRWpn
2g9MShMKJ/V4a+oQway5MNG/3wuOFusLYpoaQxTXg9s+MztfZi/Z89jga761xpkC
+hIGK6u8iHtH02eQCTywyaj5vlmY4vEHnWRg/XIV8GpsS/6jp0pEp0MzjaK53TDx
aXjawoF3DjlZknUp2pRZ8BSJZG7cZMWGnjsBvcAjRfa8vZJf97N2O1ep6ir9jzVG
8z5o93Sldt1qchLGvfBgp7+XJkmQmeFp1WQgNnGtcDZOPRxtBeh4MfOG6Xv2E36G
LQkXLSW1hPLZc2YBu6TIBZpOgoOV3KCEa01BiRmJOfE5Cj1KKx6wSb2LXVa3Tc3z
2mQ0hyKIZvYFglQHFDiN4cjeUOvrxwjx+vp8hWLh9PhZ82ZNlbnRWpY8SjCpHT57
28F0kqeAPlzSVGUmMfHX5qly5qGfwjoOKaQnbue/FOWX6IrHyOj5xitEGLzBTB/j
jEuVvsku9ks1tnp5ZsDUjw4PiK0bKRy0GbCcjPgNDj4XlxrJ6SC9YMHaUlvzVXu1
08NjaaD7/tsSTCLqxM9dr+bUYUXGRrJxAbpaa697xycaBXnDX/sKQ9j/F5A/ps/8
4LC3CsHyIbwdK/mDbwCqqZLRPEf87/d0p5FSutyydehLS5EI7jQdX2X/6yXvRqcS
efB4QA7hgNPqwbM4wMhgncTCam8/nwldXNjPJZwn31Ud+fNAJ/ISertyxD0eQkH9
aWvwV/rz6S9tE/VG0oUgFtDqtB+AYyldcXgpacBMsJkOaUZHxCnXCva+cRFZfIni
ny8oxjC8pJI9SASC6AOrIP8Tf/1/vE4UMjubWsl4HhSKuQh9n9x8D2J+YqYQo3dF
tVuVpMCb4rP3lOVXdHKfeEoOxjv4YG8JmwG6YtmibJgnqx1BxaKpF5E4KKbHlDjr
5MacmSxRvcTIo7s/8YFZHllGtcCwMYHqhfKrVWJdsP0vJB+XMfHSoaR/Ykum0h06
2G1zwOCbcCHlQN7nhKyOH6SUeCHbkshs39m6tY+4lDphwX8nh4et+M3cjx0c9s3V
AyKDlC8qRd11q9mwYbrW23N+G3lrjK/JrOam40emEvjsOpy1MGstuLNQ9Fd4KxIf
5/yu8NTO/IbWjDh8dFvWC250n1fE99YksaDU8uNcRMuyLFwU7rVFI2miMoFYnY43
s3tv2Rsy7fZmKcWmjB9o8yUvuhpouijtEJgpqh9q6UR9gF5v6URwj+4eAYUpH7Z/
3vD7vzJAoBkjlW4YJPfzgrTnizAIgSJLic1FlEIqcfKIfRtfupEKJy5RGNZy8B0/
hC+2yaSpECHB5/jeihfkAG8RqxNG65x2WjUU7rG0+XC/MVgvBGWaOPB3a1FzcKOY
ETQXspUZO1ACS6guv8a/Jk++u1mXZSxdqRLu/3rjL2wX85XK7CpX8rLjbm0ro50I
O7QvWhzinV5qXFQYOWS+CcqQhKJK9O2cTc+ML4KMo59ZGcXSH49L6eJiAv99TeO+
V7A1jpF4R4LivObnQv1VY9sSzhFBRes3WHWiHWYYz1Pfbk6WhQBRboDw+N9Cwx9G
x1X71ZptZOP3ZgJm68OWUsZtE5byyxR/dbd/RInI9hK6rLjQ5u6Q+HdwheOZg4hD
S2AVqjg+v832XhFenav3aZByZU90UvIc3GESex7LOP4yKu0zQ8xgbHS8zQCHVf97
U+E5xFIHuOyrzC8lPQbua6GBk9limWQh9V96C+VwcZp0sSkeF0jv1Ny7bQIKXYmD
xw1XXkFaBBHx7j/EYNYFGun3Y2ppagox0Kgljwgn8X35pmmupekjlYxC3ZPasakf
luA3/jfxVIGK1+UA5wLzJFDm5ESW01yTQZyU5C4OVXUnem4kkxx0qINHss7i8qaU
cbKlpZNZGSco1dDpbFl5uD7Ua/AjqzKqN5z3VdrClBDWoD/bROh/dF3HEozQcI4n
pfca9ih+4hgDMKRFWOYWOiW56lhFnY2vEsHcZsM0BifGdQUCZFGa7Enqbhjkwdej
HCHpF6lIXWFkY6ghlzgEIakzKyCXywGJIPR4PybcBMmcbuot14B1d+p9qx7VE3fv
X4Fg5ZGof/U8W9q1K+A24ExbxGcrNwk46ecD24u1QDrQDxSquTn4RtneprbIM8qv
ZyhpWqDOuzWLsaQxM2zyDFKmdsEMOrSssycryWec007MATxQGYPNxs8DL9wH40Il
euuh/GJL3UTlpMJAIL6Du2X5d9/KmWHBoRYc1T4c4qgMRF0QPYGK26mzbiKFcJ5f
RXLgVvwOrFhi8eeYf9dVCwEwRPtTiBEM7OAhOs9Jxwj0dhXNb+97dMW8iRqJ2Oyc
twfuBy1AFUB0NOR59rFonFysZ1pjtlOsrxb1yVDTKh1KvSH9BJvJ4mlDEcXeelsF
xEv4Na49RVutUOS2eFS1a+W5b5FAz7JrP4KJ+kdwwljkpB0VbddnBbEnaWfKkClM
XpU2T23XRyaWPgdKd8DutK6Q7DrDZdTAtPjeUe62DqunjA4KCaFvlyM9mnqjR7CL
r7sbiZTglH137ScZB2LB/J9xDvmXx+fBSD3LPJmY+wIleifuGzKpucimQY7L+QjW
kU46ZEKOuvQ1vCvUT92LrJ5DKPpXmPLoD8Z5BWqa9fj1S/8q+N9kjbdhSA62YrnK
JiTpBPjcg0OLSTLu86u9Bc7itqAbzlOZo/d1Vdy2rceRwMgz5J5AuNtpC4IQFM+s
oguqwHfF9e74b29pPsSaQh8HvYndFbfOXSc6hOC8Z4rVm5BT2im1xQy1eFCuMgCU
k2BVUKnfItyAPlC9tHihq00FIb92xwam/zNns/R0Eq5GFLqVyNfnGY1yhpxjnUWt
Rug9Dv39/x73v4pNEjf3IQS+6JkM/XJq5qEZHdAX3PGJIOB+UKnmbOxCMHqeYDF/
6el+seCxffMGyBDK3Segc5inZ7k+Ot5lxWJeiHxXNv9nuioA/hS/yCVa2Z4lmJ+U
m+nologjH80G9d3aN3sdH473uEBX9Ncc8b9CYxrFwZ7q9GMhuRkrv6XZZoM5kSU2
LA9MQgg9S+fFcyFcS0zIuAA6bTIBj6djzPtUP8Tn36ZB1L0y8M9J0etL+8maDY/h
gf2NusePbbxC+LeoPtMiQLq+DkwiJK8thWld+Op73RA9a0lMcNhsjEJIQDpGaUeQ
7JOf7GukakBnoWbknVvHqEkc/tiBs2dhxFWEuifkC+WUKFaYOPZXicUsQLv49VKb
Dt+BOCml3hGXttU4qBSzmNmv/Ju4ojkLCOb4iA48JSQTUL8bI26f5+NtOF+wNlCr
0P+2rwmL2hBamM30CaBHHNIh8mP8N5T9R6S1zNKE9fOGxfX04fBo5+Pht7iQBtPN
ZuK74csQ8q1o2bWGfyppXyX9jHUpCjNlrGTFnVTsH16kOrilMrL8adYpkT9o/W6P
cVo9/AkPrwT+xxqz8IUIX3/c1VZUFzkiCrLhrPBw8gaFA3DjYlexvHlOg+RU5H49
XErdDzFBWFvwo7hV+5FK+b6muuhm/RVZvyK6O3gNXDu6JCMb1vOQhD9oK05gwns/
z0xQGbqJAnKhEBIj9sb+/4SBW4ZYBQwH0fPIUlXeQe6ePkANwtvDshwY4MSS1nFe
MeQ3498WjlrnvGFz/ELzrtgiDWzlr/EQJrRY4qw+ouCLxp9nOhMooNIeLmyPXjP+
qiRDumWs6F+7mATNZ1ePsRgDPAcn0/zhCz47HssVa5122ycfO9Ipl0WoCfZXDRLg
z4seAKG1/zQo7a0ZDk9DWqABi1wNTTcqrwnvjRhFryfyZuHY4rhMlEDEx1KA+zx0
IcrYeIUOoxAcEqxdIv3tIjjY9wV9rK6jAr2jSxNI8TIlD3sxJC7KzcflbnDypEHu
hqaWkMXDTvZQJ34xvK0Gzjj+9cHNUgvG2dTO8KD4mkRtCJT1GzQoecuUdVH1H42D
Z/wvhWgwp+W7PZiuUhjkaMHmiNpK1/Ni3FshTanb/n6Y9HVDzxS7rGR98iXpqDzC
kAk8bnkODMCBisJEPDtLHeC6YeWraKe8SrGcDtWZd10rux+zq1tnvcusQw6G3wfU
yBPjMWWl4CxnoBjSiOpg+zFfD3jpSUcPOKghDdOFXQKk6k3p/DN07FcMWepSBXk4
gVRE/qR7+inaHTo2QxSHY1qgC+KKNRGgkrB53f59WrRCKwCKt3T89UxTK83WF0p1
3tvkDP9XTmtGYWKnuR5ZmdGuyRgLqlHbYFmT7hkA1zd76PuI8PX7+3NPDTbCEhDH
osFQSNOpehIh759OBqh7j+LqkVi1pq3gMRN0qrtJPpj4/IZj9yNgqfQqt9xLT/KE
JzpcN1xsI/5HptZ3/iZTcQ0m4ez7b6RKIWPI4630P62j09vtYjcKEqcQD+q47OsV
jj7QinRYhla0yUogkqoZeiTjhgE4LqKQtJCnNT96EvuBl2NfMDr/BzsEr3aGTOCM
Ce8v3IwKLr7V/o0fxl8Or+X5xNsOgyD+a4o6sAzMYQyMrLsithnGKfEDQXWTfPTS
tRM/IQN3iLlrUznsPVnYSI+1jHHegDqUGaFMKJqwf8o753ljwFaF56fItPySNO6d
lIUSrvdVg1Yx/iUEwo112jxTWw0N63hLPgs18Y7BFUZD3vUvc8dG6bo7kqAO9Mvl
XvG8mvzxm+KbRPipQevMOIIQ46aB0RG4yGJDWHDa6MqI8afk012FseofU7kojvyg
7mwwWkRqqVfTq2ODk6igFgsGlyMlGj0sdTfW9fXIHP0XYR1RPhtYDFCxeHhdyBlo
s5MrdfKzHlC4wO70hpd4EAyyngBqoSp4uyTQrwHAck1XHUjsGhgqWoVnLAuCPuxB
9xgbQzEaMENxnf/X26ChcLp0mDbycAGahMOBhH+YsYLzBgqHhoPLy5N/bJXCZwMA
FGtxljfwWY4t0axl9UeeGDhoBJRgl5YGgOSu8TJnBq7gtf9lX23J9mDj7d1RY8vV
1Duxo7PVUmBcxuH5iDLUm2r7Rf/pGqwNrsQMMXks14JyWrBnTocrYR/DcGbTtkB2
zvO0q8lEJWatFZ7D4Cr+B3xRVXPxb6WLAu+x05RslIxmWwfu96B1U8vj+tNPND08
TX4ySYWFWw+X4/HCnBf8HRPuVL3JyLXcEKB7yT8xtjYmDr8+mBvtMY3834UWniMT
WXDlRdKEJn7Bc+ofaNivgz1fwkgsLEbi08xIrxVDLwYOS4r7c0j6ssw2fLsgB7kf
Bfg6zVndrrTiX0XWyTzNav2GJ6pLp7KXXi2bH8Z5TlxHQkHgEtk5JH0x03KCjr2l
UqdhVh9xpEGdd5jdIqfxJJQR9rQFQK1ytAqqvUEKv2Zd/qDfZnQcOhRkRb2KQGJv
JJHTlZo+ZndITLdwp9JvpZtZsYtnIzGAzw10d1eioLTxcui3N6c7s9jTm+e19pMK
XLwe1eZ8vlBGGbkJBUbYO8I/DFH+QCXKRPCui0bzzjv3t4d08at40hD6jaJ0rVk0
OTDdWDzdJ4nnhiVvlV8J+EzKCBEzg1gmPM3bit/2rtEH/FST3h/jEJFc8xed+qvX
TwUQnlUAnHFo0oRFEmP+NrwFz/wbTQJ23REtbQHYZ4YtXwveXZX1ieR0NT99YS2w
wukZ0Sbz+x3ZapBBKF4eKfjp68QTjqfmNDWyPioe1j5oLJQ3+e/khVpjBMuZbqCt
/PEfsLSHm6h1IYMG5pfzlFufFTW/bebyNA7iNlRG7sb05PTZhfE89dCoJFlPjJeM
ASJD/aP9xxBhC7MGJmL493ZVn90MeiGMRJh3xzt7No6N7tHFG7GOjlcGkc9E432l
B6320UtwRgH9neFQQIAIGDo9B/9V1hQrARRdnt61pyc57TvM9uy7hOhgARKZ+vyB
0nKXItfmoRP85vkt7eeRB1bzyYjIj9YGTYRo6XIQPn3sODcfqRuf2ouHxAZlFWlp
hSmj8cf6yPoPfFDiBpnwe8g6wG6KKykJxN7U8mcovc3cnL9t0kfB2J1MnIiH08OU
P6/JNrg1gE/63xbdJeR1/v1vVPLqe8k6LoSl1z7R2ZdvFcBtvVgjlbbEPfFSm3Gw
WWrkh7glUu27n/0rVr9/FrdLynAYYvEhq2lhHHlgRcB3c4YXxekP0USm9JGJ4mLJ
mjrMwLsko8jABjUXZLU7JE3BjkVJYctbSwA1mmqFFZ+izpWxlIXzHLH0fkooAijS
sYkOAX85aqBm28ekM3vowLLo6PAH76ndgPDSAAJwCyAd13HctCO/t8wmbyAf5SBT
WJGAsFaW3NdByV2HB+Mtou+zaFdX3LG+2/xL20rhbpHWADQhcN5dgDXLN+/l4tKA
47lGNQslJyouY9cSasfSzx8hXAcg+1/91pYSAHsEm/+m+FAMHPiLwcBAIDVAWye3
QN3m6854lNhc8NtgGrBq8gt0TZzOc/hoB/Sdwq/dO98yrA5A/BAwArMP7G/jNKrC
ljT4TbXSl7Oc8hSrvKqXP1DcrAAftTNSu1kRXoP9hevKvD5I8KLdzaQEfvxZULs3
msEXQPZDq3iL9qLsBjpiARWwc7Kprrwb0JbzwGdamH8gqMwpt1l3SsEE5D5wGIs4
vbF8bKiG8GpZ/jyI4uKSxT7iUD0zlRsbXUuLhOCVxLClJPWg4GedDFEfnEkvib2I
BO0F6eiZOi0YFPUhO6fajyjRrujZYFiqFX7NrT5wZ86pv/JvWZePRHa2rqp/iJZb
Iv1Oto3Ruz6YTCjDFNsVjGWqJz+JW1ozkZynT8ePt48QDVKevyJUHY5Qk0OWjm72
VxKwtrYQPMn4gdijwwEoXVIpmCG5PeNPEkFRc8L5ZNgQLw2IS5EyuxN+VhexjLBW
YTyBivvbycLgHJUs29aBDfiHAxkdCvzoGVomiDOsaAY5xBDjVgvp0G3+JqG5EmYh
OsK+unsV+JEqScMawX+7kXGbmZbVrPHFnuRzZ1voFln+DNawoL7VjIDwQ/IPguV4
cfoT6lO4M/nTsprc8mVaCH/wVT13VnvWbnRk/K09bIgC11Bj2yjpRoaZy4+yB2K4
8md8oempCgRNswIaPuRyMEkWXAhdkmxBPjJTUhox8wxgB2NyYBw2nIo/nGnALT+k
NxNFVBdj6a0gt0gyW824gCp6VYmpQJwSidufTAuRIwKIiXUj0jOIDk57M4TTgDIf
UyydtRMzFIgFX7qfrOkfy/ydQX7OE+8GRAIYRmKiKzI66eMTRPZfXj3hKTjfyvDD
ElDLXnCmxBX3Dco+AihpmACS0Us8MWoOh0W+wswiVw1243IkeIB13zsztriR2aXy
AY6WqXFGLTfTmWvCTEmAYLYMqnpl+1Ccz3FOxR6ten75/AxhxnWy8mCnChI1A6j+
k2CPnSO/9VIqCO0mjGaPXukomT+XUG5p1H4kvCnrmuJqr/MvlDMqv0ZEzK+fhML6
HSfxID4JEzgsfQdSMp8hLkQ3wZyJqqQgV/vkZRtMJeHV2Wwzg4M+1ELbK4CseVqq
oXWrIv0ux9956s1X1A7OdX353a3pq+FG2OqzwBYH0Sfb5srkuL4KXxZ6LaNPnYbs
SAKl7oCbP+IVAqcICepjuE+kF4dgRW/UGkqUO7dGzATCET7FnjcClmRCc82s3w1P
DmxGAmKYj9mLnAd831E6l8gVxUx491+KnFf+bJKQUB4AH27DvhJnJuiuR8NdRMVF
TilBZhmKbiiyHqTUkZPmVCgBC+teCo49e989rAU8nSh9DE6G9qmPgI+mBNAQcoIG
nrbNpO53gQ2CHmCC7CC4LRla4TteqrXTEDM0Ko23+zcry+L1fsQyffzu9vL5qa7O
AiS0kQpeQCouqJ/3IJDrovavecmY3Wzrl8EBPZlr19CxNpmQhqlali1gA4E4I17u
/4JRLlBjlbIxnPW2Tn9tEywNmpZ6djZWaLi+s2zcyTKMtFeFj7rN/4uNlZV1AC+v
U0NeSJBbP6OqYgG9JIwnfneyi9+vrBHa0wwFIBcrSJBn2x3OZPiw97nkmf0BKmR1
rKTVyZk+DZGMeOhlr9T6795QUA54bSOjuxjfh3pEJxe3PNvBiBIHlbKN7WSF4Qd/
G4njQuMWAn40DT5NVO7beatNkTtKVBnw14bMnDEjyylCbXNJCIzzF7zIhYPEWucx
adiWJmQg2pJ1KPmAi51VJgK6tpavL55wrYrXCQA119FUDrmJ34Dh6jHVZrPPBf84
mcdjwHdU/3YfIwv1EQQBAgzP/KGTVwOodG6FU8UI8fhWQwglaysapTrh2+hP222X
p09GXlNh1x/QP/xNt3N5T/tVDJHjLr3fAHH2H1oVIUnyULR1fodI3HWnHYn80iub
EBa75T6BA3dqAWo4jAvaMzDpAkJ/LYjoJDl0PxPaPuxFW3Xb0IrToPcJTg2DaB+m
vzDyfB8eZoAZSKX6MFjLhd+mvngHxq7isoH9K6ofbOaStSYdqKYum0lnjxmMl+ab
yNeTPlYHk2Qv9RgRm/eWJnzKDDNfoY82MygbaTS9YtMq60DZI14mOK7WDPRkzWOm
jow2OR2Joi1tRlw7BHCfJrvL3vFcam6aE8ZW+s58ZWlPgU5WChvjchP8jueqmm0Z
hW7vE8xQIVJZPG2RpNagM6xrlFiobjiDNojerXHmJKGdc9OLzYojku0YYFIGwv1G
lGYdtID5camSPvV+ch3NosLMAod5uDnfcpeK7F7VproULP0s6j6tpvfF76U1uFrJ
4ssSZ9bUxt79FSI51fPHbaPo40PC0KQLk1ysqeiflTyLQgZv5X2lnKuKFhIQOwwg
sD2G3JXtBnzEFsLlYVPVi8MXWb2Re+E6lle+1cTw2wsQqp0i6dF3WsVe+DvHb7uQ
c7pldL75Gl/xQl8CPUhj+J+mfDAPakGTohCyZQ/A7Kovk8FQ0eel3cthkIgpuSxM
vBA1nFtA+oBKQ/t5kKBa9nNI8Dl2/QwCojDdI08Rstx2pYFsENtPxrj9QwDSMWSf
DilY647ir5p6Q+M+jubomQUYa4f1RbgUwrbbVreyFyBbM/2y0FsDWh9aZv6Zggpr
zwUIiAGj3fPxKU7bNjWdU6ynlYRtFQojZkFvXeUw4UbCCnEN7GADIbZzi2b0O9EE
qpYw/boiHzViiPXkTQ3YBx5LxTVwB1DrjbhZtSZq+vSM46i/TcZZAKTyGD0ce+TH
KqFHdzEn8i31Gmr0O386981C0IIVtL+uqaBqoXkRojnLoqnVv4uPSrE61HhZWXLe
nTEsAcbR5lghsqu9YVTUVdAevGwLDn9KxaMFhDEUc/JdV9pFmwb9a4tgYElGlHak
JDdEVFN2SnYXCa1C4pLGBOb8RNQj+rd7XHkFjIuYOD1pM5jvyfoXmpXbkN8xVCdY
XzmKB7G1Ocb3OcB4DucxBYJPW72svNip4XP9IKSCInytMRGPKnLhYWtyLZ+Mkzr1
hoi8fyJ8kMmGPm8x0VGkcN75iYLqQWMQFFUOJvGWSsaX+QI+3iZpY4m8wnC//Avj
wm0rxj9Hx8PXWdHRJtPvwKHfkiuSBm+YG/b6pQnZz2/rNNNpGySk352CaMp5xTGb
01gAAxIvMyUKiZWoqo8QQh2c4pv8PuNrgLi98KSbDmQSh+x55UMTi2UMpva3AZ82
Mdi4bXAKWq8Ja2aE8KmwEsXZchfnFmyPw9J9uXxsLQiRS1Nw/h6+DYJ/jBJrw4lz
5Mr3SXU12V14DwxvKq4BxpCGFuow/yzq3K9QKvdwIkwFOnuOTXI44T/4PJxli9lU
rRKkHKkXLfGCaC5vWvWI9EkJ8cKbVvUHyj6jXjz+jKNkA2yM6Z300VVNIgVQ703w
XIt9/IbioDp2egGLQPFYT+9dWlDYoSt0vEQipjAh3Mt8w/vA987MwKWlrV5lGOtO
XD/XMeH0lfaKPbZZ6HTghtfcJ2RMF8KA/pq8IT7Xb/3+xJregk/zbieyMXr9Hcgr
EwP34PhHhDAFqFohmm3Mf2yQUB1Y9c1bbiptDHQSwAqhJq2Dle6GNbVWhkEmhKBt
qfRo3OygFyoafUut5ryp74PC7GIuXAK5PD24GslBk6L92AL//39uY4/amW5o6KBA
eQjaYOOaDNhtypSfY6+a/onXunLSGwP1SA86YB1HBCV+tUSdxhotF8360CYzf6XH
DkSARaLZ4gR2W32MFw8fH2k4wuFRVnLmN12sWucm6A+1ns0+DNEdb8rsFzJlrmoc
STUBNQNQ0AVHMuDMnS9g7VOGFlYI/sD9THC92t9HY78BmiTZNYgETGqN/0v9IjH9
5ZlAXeMedVZ2slRAcbX2n0zoZCS6zEymgdEnl9+dCl5NB5O/VfKkL3UU06HnYRHO
e0mkrQZV1qELNafymykmQHw1vh1M0OOTlA7dLkeWy4bWwCrIreJNeALZb8bL8Sgw
cYXSNTbjyyWQSIED+sTcxXMLhNdXZFM1EO9vA5tCj5gl68YqmGXCiRmw/TTg5Lfh
l+bkjUFgIJdPazQkeOTeS0FmbX/SN5N3OqkfeJWz/PexTNoxqdVfF5lJRYtYVJ9D
cVbh4VtVt1aLuTKW4TNTQkjdQmuX5nX+X7Aks8b9xQsf5DtYigTXyOQzK1G6Gcii
K0Kcs/MwYJByl5lh8aej/8NhKsBYTyNnse538oaTOnpQ6GhnC4LJeM4MnvP05ZXD
WRvWFe4SfMSqxEfgXIrrs6dsKeP46D5MgzZ3eXukbDlZDm8Y5eXzzgSASSyE/+4S
4GNp/neEsAmCDgdtiI1AuiSKForOYkpEVoL+aFdoqutyd3uLqZc+ci7wr5F+5hxE
SIXwfybm5mJ9s0+9BauYUTHb7vV8HsBQbRyJXF03INkUbdM/YyQg2fKpfM3pz44K
XmSwH2FmdMsBguwFnhgOnoY1n8deDQzmHSfm2efCG2k+VqAndJWWpeNudP1Lo9EV
mH/9ZMAmuJPsPfzqrFni+eKELd9PBDWuR5IHSVZoZFA46lLkMdhnhtrmy5jWP5F0
mFExmtXpbEs+xPQH2QLE01eQZgVYT1buySrE6u6XQfoHe7RC3rgeTQppbXbB5U8r
KjWEu6GaYqAHc2NJRxqQ2b6kb4yCRvnbhHhm6EEzUMOFGAUmO6UJCk80VNilM9vH
PQaDBs5m/dgCejUDcx6qiPc0qHtiuWhzGp6LeX2/zCyRDDRg/G48nizaWsFiLDTq
fVIf0jDPJb9StSuxVGtEV5KR0UHfvAO7q+wTnXmGL+2F+Fo05Gn7PkJKNg5kuEh7
b9ZO4JkwBcKRBaU7xmA2p5iBOBBtbL86fk9q18YmddiM4uktTV7onzgHg/8cutA3
yILwh9o7cFpZKewbRwuBT9NqJllvoFIu62taqY+eweWafOWNd37080i+NdshP8Kt
LjfKseScWVJXru8rbWeUTqEZP9vkSLDhSGYeXo5ADhMGYBPTvUsSMfluiRhFgHjR
SG4wekGk3MaAYa4dPbpkiCISVBmmwClq9eoJ2dNosQdPO0I0LKzDj9LV6juSbN9r
9yCcfnY98lW47QeC05zE0AirPx1S8OdnBcJJ4HdQctFMpCnjrL5VFR/dxi9aIV6X
HattTVZYlMF2iHgtHNRrUex4jumymqfupISv5V/TktOt8szOA8ZQDEmEzdNMNqFd
ggLbAhPV0ZArjqtu5HCidNVxf1C9w5Ja/86BQFOJOq2ofLqXOS7OCvbJtjd3C4Pq
TToscJma9vEJ/uEOAAZfxyppfjHPUzQQyjvUeiKa7tVEQBIllmi648/FKBLK1PRj
HIFR8JrUEygPgclr+gn5X8mReQGH2jzDak5B5MEVAKA+QXV4f95hUzcGAW3RA80R
BrBZdru5obcCmon1Q4Wptl35Jn2vsbEpA75D81duLnOh0+ko9SHDbd9JDsYopwFJ
4n8yeQPIyXTGLTQsNe/QDQPgJlWcTw0t6YMUIODGyo1M6YwA6d7oX6aaUrSFRLtJ
CCM5dRq1oV7V0iaYSs5teeuHXnf2JjyDHLayVpkFjkSliOSz3zDuVmSs41owlRKo
QZqzjVrDdchWKzwmEAH5WBzVcQwG8NYDAH5w+iosVso+xd2m6OxgctRQaaj8msEI
UuP0XzGgrE03n74BkHymhfjb57gev4vRlHSWjmYfltmSYcEKwOL6A5npqHGBZCK0
AfvSSKI9E+SJbb/+TAmuPxKS2LYzS+BkLx9WVFLXEtS04Xas2IcLzUpQj6X32j0+
Z0M1JwDdk53RAf6w8FJOCkj76l5HT7FdVPne4hPz8q93yyEUVa1X5ElQTcf4vlDV
Ae3SmwsWY6gQomnxkkVOjC7uuUSNxd2eqC9M7mTYzNdO5A+ZRJtNa35UE6E+fnLf
CWg0FTY21Yhq8kbs4Mz9mc7PyMl7uls4FRPC2yi78hf/O3ky5y1jHmtL81ER4o6y
Y4vKfBWMJ3mLpGAMNRIZBErY75oS7dBhRthSJCV3fFOBura+vZpRC09f7AXZuxvz
kTSnWspOShthLXLxVsAugtek7HpWDZebiVIn+PaC6MVttuXYKp5WL/pznvxiaQu5
qTJohc2MjX4+Yr1QaIBByNHftAwpdx0YDCepyYnEOTm4YLT4LjgzBopJPYOTZHdv
LetvPgmHoISqjFsEPObAbwbRw/QnMwDTyCzXh1gS2dqu7Az7kaJi/NT4FUIGYdAa
ZKL1tmG7eKJ4jZhkO7c+4D58v4gY5G/lVb54SdxFu6NioH0LHhdvtW/k1wFawGUx
VnixB/AqrJTNdp61FuAkVAEdUDzLUkTHw6kxGugLsgJgN2PfPw6YGxeBb5WjePxi
DdvUgr0sbeW0brDqXFF1JAwDOiI8YqDAQtlaReLSYnM48JD0Etltt+KgvzRbZlWY
Jj8n4XFyEZLTmHK+jt4DmV5XhnWLFXZ+6vsEzTtcaYUcH00jMqxZaZluHe0fgaLY
rnqseMZpAA5wrASYXSoLPyxryvN6Lr/w9XWMA0HduZfC+pR2UaY2qBN/STeErhj6
BmRXPK0w/GlWQbrlCeO9fxzbLEDr8hnkYPQkgP1NDq6FOoTIJ/xiJ7L0egI+mLzm
1QRP3lzqebMMJN11idzqTTMK9wqbdmKPjMa41KUN7tLi4x8r3qP9EyuFuMVzj9o0
Vb99JKB9NuD6a5rCPkdI1VJ+/s3wv76Xxe/PXgu8++6x/ERS/MKUEmq5cxJ1bHGm
epgNaqL+lpgdwAxMuTRNSQKoPaiZ3QRNZRXoK2Ph2XqyhNBIIopTn9qq3OFmFqWy
USfLJADj+gBlfwUqQQt5lKnSKzEZDnuoP4NgdIlqnQFJ0nJ8HuetfOr37jDzjlLN
JL93BYJZcM59Mv78+M5bHUJsa7rQ7Ob309qCdVPv1YjjLSYMizEVXh3nvhg3Hp+c
1ozGL/gqSWrHvS1HlvhJcD0a7hZ+74YowA2hvbg5N6vQRrngpdl8AEsPB6Hg0m0G
1Or66iibH4Ni8fnTQbmzqwV4aHvYbFK0X5pCkmA/NNvQYiYt5lpNjVVwEFu2/ZLe
G3ft+zzQiZW/JCknAmKmym5k+O8vct0SNIwErOoUd9qrwIwq160n0pKEEeShcegA
ZeH+5IfaZYEzT8W14Pwv38oimxzXM1c8x27Zbq9kn8WcIeW7FFjUiFKfY1BnomDP
gq13+lUUQuD6MDWXtFVVcLX5yyUmEk/PbMvN4mlpgws3LPnqv5AawHvSNQO8DnDj
lnmYzqErGewi9nVDhmjYq2eQv9aW22W02KVsBwaFIkN06k9w2CB+X0U149Xr2brV
ggENR0As3J3RmvV76hxxaEsolNeUq8fQ4cjZf87bZL39z6LTErH10RFVCPjrw+QM
fFrijKuSNMYuvqCrk9fymyxfLutISZqcnRs5JOu2ZYvu8osmvg4HbnnYPEIP8osV
U8z97xdFTZM1MClcP7e2DXhBCXtAZSOeQbyAyB3YUB4vChqQPoKxvJlSzM3EfqaR
0kwPn7slpvDpm3CWOO2t8KijM545bB058FWa11koC4f/mTjOwu6sDK63uRDr1NAr
vxylZPsf0rudeCnHbT4lAM0YQmmGwFfadYsgAzn3QcAnUv8P6bQw1Hg1FXV5OrOq
pHFzg1/rvd6HgCWYlVtac4s805n8/MMJK5ZuWRnf/0xgJCV+rviP1e/pGjoZnODo
L4JlIwTy+hkThHs1BdpFHYZvXKU2ljTwawO8mJl/8VQriMkcbc4xmsUIbrbyopxl
oYPAmAiFKc82nq9Vmevzdk8Z63HJNxLbu27iVdjs6hn+0wqCgYNLy8EKHsGES0+d
0DZyx7Kgtjy23peaPop77Vhw2RIyn9eclLnfkMV3JpOAn+iiDORZkPzn36yqp/BD
EesMpL01WfaWnAZczu5LRcD4/Q4GJQw2sCREt2Z//x+J0msmVfTzFO2W84F4PBxd
Omd8mmPDanrG5QDjIgG2kIX10WAuh0fTiI4kZuIwcP94nrE1E16ye/RaBZv1dMxm
t7xLr351pOywpc1yderA8F3qZuOrWHzydIRhtx8gc96wdAFlgI5KXN4gH7mn3/Zs
4C0YvoQpBMGMm3say0oBIfkblwwd2aA6K/QxztZdOGVTKh9VH2JuZesWLHLxLBwU
+BCdvcjYG6Nz+IBinurRjzwOzuFnOYYBtqu7ZKxtvkXAnh735gZmPd8VcljQe3c2
IvSuc2cA2dgE7F0rXpesHRp0CU8vrd8nBLrIzg+ihMJmjXjhhprCG0SVCNTm9UmQ
w5YXku7XLiYsuxGQ581FNt33XGgenPnpu39FwkfG4vRyL2UTqukIg7ns20bY9l+q
X5jXVHJAZh8Iu5wgtjvH3z/tZSZkp3OzwC90qiOgFcJU4p5lBWHzSHecrfFPB8+M
Y9dDo5d9jX/kMcOoSjlvDCIVC/0u5s68BoU1gKCmiITcvV4dTIbGJahSB+0K07Fe
X2UGeKttLUekNvoBcJG9KHniAKuYo2fGSzEZ7A/IEBIwbjt5mmkvQrPGiua+So8j
WL/V8315ac9xXRJ2uG0ArMTFJwPCbXu0vXCYkhnJXzt2qx9ERsN3lZpiGQzgvAG7
fDPAXuM502o4vRabOMyuDwc3Rgaij3nwHE2F1HeF9+zphEvtFp+rcbEX3btnVeL3
OrTFln44++G4c2Uowcjb2zNWBCZPBD39hM5O1fllRdHdsecu/B5iBFE3msb9+bpL
sAaM8La7Xj7WLz/YXjrURYf7bSLO0ogH4lBIptKebCHD9r3Bl1RVxDMGevsY26SW
p+RJGKH7vdf2SQkx8DKbOPFkrysdDSLupTQEVt4eT1ISh07LtNlJZ+R7nASssjOt
Pt+6+0LRNi+D17aukHmJEvUEzzWAob4wbozb9pf6TJC/YDgjpdjpg0Vd+Br2FQTT
CIwaZCCp3339HjsLUSnwy+SVp3s1Ed0Vf3Wc5X9gxWLh8UNi7yv17uXflgxlSJ6x
UG2w9Fxl/wkOhIWHqTSqnlv9AwtGQu4LXZEOapkQwrrzwhnIldyRw/zADhAt1iNV
de35uePb5cU4TNrlWarCJQvxAatIhD/R/VXtmlGaYOXpi5tN9pARP6TeZ/q8t4gi
wEP4iL84ynoWEO1jnGimIX2Mcu55KTEwouUPQ7YWxw28Zakv/FTaZ9Kg8UEYimJr
N5CXfhUEKtTp2dgo8wZwH4uMCPke0cfi7Yp2FuFhx+AC2Ipawg2vStXbXnxrQIt0
aJUU+pMkFcuc1mjfWvFGCI5WdBdv3DTeueIQnpNfL1Ag2Xx2O+4sNDIpXy/UbQ/y
QgIs1b4BB4vFhgD72TQ5ZQv4xCAjpzlsCT+eLstHt9zzNZ0bff0KFYTwyGDHHBwV
36WT/n0/Vw3DlULZ6ylAsDs2f2cKGOQTpCJgPHBIbQ80LavsNvsfWHJdUTv1uJ0b
nVwoGMQz7soI0GHGdiMqqHV1SNpbhyC7RiwiLoTKlkl8eU8WYRC+RD4HRsxaStfQ
5pp/7bX9mF16Jx6Q1osnwV8e357/Gtm+iGm1Y4K895mDig22bLHARcV7fw6a6Ybd
XFNAIb+l/AZQhQn6LLB62BIbj3Awoem/9b2oA0+HHpnM/B2A7TwrEB85N5HgsWBV
5Ln4XXUKI4v8+m7FrcIBnrGL7/qci27hgrZvp7rk+gpYBmkE3DKYeujCJvsRIo/w
+HRA38dHUZ1pnzbu+sOebjs9FK4eUr/xG3srAmKAORO1LMzCuVMCiWUTH5EsEDTL
9lW0p7gFA9icwh9Ci8iQN7OC5n4ECyhj8im4Q1N1UC3vF+qZ8NspedYG6Xgk5l0Q
Ezcm9ejBF27ZVJv74WUL6PxlHrxMYgsGxSh8TQAnXuOcu7RPcj7N6gL4+gMJRLwU
9U95ewWb0q5Z39Yo6tEOCOkNT+ChJHgyl3q8XS/J/N+d8ibRFXitME+2/OjkeSPy
elAFutN7WWl5DQXnJXKytg3RlFQwNn4uNbl9Flz4ycA54PMHmToZVvMXV1ueWT5I
cXSI303ST3GBr99f7pKaqg0unjuKhHW8vrYQYaNfNISFV2hdN29Cr53v9jHVR16C
HQlLbGfLs44xKTSnddyTru1Q5aP6kuEVUvjJl5HxzZbV5vz/O5eLprcfWvjjTPcH
2czHPPoH/tPykZ2mcWkwwqio4kRBlLjAqO/B6VzKkmDFxZCiteBeTUU1KZXAcCu9
7DSnTg+6aLBgRMxYtx1I5+aTiEl1g3E008V9ZdMlkpuYJLxXYBFKrpNhnFu9rENO
UjYAbaS5geCXLUh6vnEmPC6fpqN6HzZDOw/TU6ydtieNhikZpkYf9x+kmZS7+hZL
fUWqdzG4W/oTDhjf2AVOdiAofPzij4MytC3oIj3iLgaH3Gjf67O8TcJ9j1HXaCoD
0C/2ScGdbNxlckcOTbJxPpH9p40DdAmg8sPbYNkPAFVUdIsbadLPShaRbJLF03uw
JSUdT9F2v+/qe3LLzY2fxRl7JYA1OAx9CY/XspOc2g+uexHN1K5vkFIfhqejqgy8
kaNXP4rQ1h1lMBgnCh9J7BR20B+Yb42+cyxveZOTaI6Ppr8MkLym7hqjl7ihIlTO
Fc3467zY5sF1WOh9nk5wz61ob/b/WbjqvS41Ku1JxIqDwKo1lH489jPJDAzgW4xv
xaNtnycbPsZzS2j09B+oCYV+VRjwwpdnPRE/HXYxATMcb/fJq1UFOTnQiErPF8Bt
9xWOZNZ7RBb0IhhuwiyHG/lGb+K11QuGBderHLE7CoX1Ha2mhZnZ1Z2JojYwso3j
wLrnmGMOmg4AQdlbUX0m48Vf/hOv0iqbZwLlQ22pgD1QByEEDkwwx9ra5ORmJrLG
60++AGFD/E5o2Gl5SClqbzf5sgm9FMX4WVqGpRWIvBZSMc+ypbqcmBZZ9rFW0Olu
9ZZYw80hIA3tVtXdkDIUXDFmGVCCn3UrzT7P8Bxlp8it905Y2J7Z+FbxbQDYpAKA
nwy1BCkf4QwwDg8ZpAZFamL/Gt4S1YM+mGDXVk5I2bYcetp4mlsq2Ks1JcVAcwKN
xIRaljg5jFoxIhqrybq70DjJzEH3v34NV+TZhWvRREPVzM+8TT8ZMUqZr9kDnfgy
WdCwNuGHfPMtSPgI0G4hB2KKuTKngfVKU4wVyiA7zGAAkg22RMttWvRBzvctpW28
VQz5wlzK9hzAag9yAT2aXBGa2K+DUpWPVPUszaYqE+dUEJg5ko/JVRCC+EwA+1cL
O9GPuUwjyX284ukfXrEEs1eGVEtyyMyomnaux27B4lYHmbSc4sVo9QoXb6+ok8F0
EIbPqreCjosectvp1Yt4ptNOax8qAYfe1u0MMrBBd0UZFH6gj8KrJ1xAcoYHO2TZ
EPx3khb4hwvpatl8CVbuk79ZMfuH1PVaXn0i6tJaJ85YcZWkyBwF8/bvMxBDLdE3
pnO3JOKBDo/8++Pa1jh3Uy2yhPMY1cgcnRoNCXz8RgNdxoOZaoZp6o0vPzeDSa+H
li72PTO1VX+Z73eKpE0dUG+2rvBJaLzv2oQsfdk2E0CYp3vZ8Xlqsp4VwPaOQid0
UFimtAS9hLr0UBgQPElxhrnnjpu2pSH1fF4K/lqfU2oxJnp7qmUtWjhZuntJik3z
SyopJwLnviqYLJHv4uIPvjvFOluBFstrYiOPiEwtSscM/O8UtzWeQ4Tjg7KgaWW7
OgKCNaQrXBdNAtWW/CTY7+mnxLC/K7YbbfkIl9NITXwXNmNSJrmDFCmWBJgoQtGg
KZ1MlhdYoiz8RQvWVFG7vG8zlAILrOFqQt+GIQm3dU3v6275b8GlsjopeAYD8HIU
0pdED9dJKy7q2r7LtDq7KnlZ1twpSl09cKL3GCLTOx4ShwCVcxlJbCPG5Ltc+UEn
DNHtNiG2zvgMPSCUXcQ47DNitLpkO/zFo2G1QeW93XxpHjRhXXUMwQ3pqH9XG4Sl
qbQ4R48K/C2lvknqruGkycHjkuiPfMBRVFexLSlXLCos4qPJeDIBMqqd4wxFXhOQ
SZS/LvYb6x+JrkyB5gh7+s3o8YruwVa6PsLZ+YQRSa7gt8Oidmrfpmqh8OY2XQ9o
XmO/hQoj0JWztCKUzu0++6/eVG3PUfCIvvVDRx2eiaZ7KK3+D94+MNB4qBF/GIfV
jlPt8K5gxCJ9KXct48pe/JNygrfcWAcs2pbS3DgJ8Zo5bP0PePmoYV/+y/YNhvDO
pmKjHz/48d8lPH9dFzNr8UjyZnped6Gd0xQRjChJsYWfpPc/apCV8Bl4L9LyfzWj
HJlgF8yy2F7uTHuPiv/RjznSGzgQZm7UHpAmk5Pc26/zQVvPIZTWyEYmk12k7Pen
GHoFrQZ5/CiYb3w9mle80euX9YTdqVX6ybMbvbvWJkvPFuZshMYVeI1VcAdF8aKw
FTLtNCPpqV5wGfstoHzI8CVYk9Mnk+wCIOfsakrfPtRJp7haf4OApkCZD38Inac7
63q8cG0r7U8Xz6n69o3jJ0xrT0WUww1/DFbvz6nRYq2PtM4sErSUvkDtkqBIXIUz
vKGEV2XDVojeUZN3RxAmp1jk9ZhtVCWS/wh34DV0QRj3VLYj6V6krBPRQAArVLNP
rz1nT8bVNcw7OH1dvXZE45HNtWc0XvacCVhvmV/CIMQ8lDeNc3FvaFikyIBmaV3T
hSmE/EnyJqMdU1iHVO352KkzfPTOF0EeVQz6oKLNegn2xdi4xuW5bJFMUbbiTWsQ
MPYHqxq/pcsG/v6AWVdG/DKuPCAc5dehQEO7YGM6SaYYMuuNFpXohapuaSM2cfnq
y669eVauJuSnju6W3SvLmxAyyszoJfd6OIpirG7oTBdUz3r8aiqDtm1XGQwDNBG3
lyhulalbPI2BHsXztbDGTug7BJPK38T1LA8rw2FPy9AGbPzXH2TaglSefEJILx22
HtF+B2526SYqMQ8edNQ7jbJm3L3eINf3liRwt0RJCSEMWpuuntQlzrLg1JeOX2OX
Qk8I+6colsQAha0QKVa4BHZ7cV4r+s2877hY72JzI0OaD7ueCyEJgdOnjcX7uOcA
06AXMGmVszfiSNpmykM2rFcLS/2WCIiJWAcU+ZTz2uTWTn43HFwehhXZ1GOQem62
8M3is22w0ci4KQeuWf+AJOl91U2wEU6j013BqAjwaYIf1oipn1EPfymmp4NlLr7e
zbAJpgui+1T1lh+Y2eu7P0OvLax8h+FF6vR1De+bEy+yOHJLQVEAYsIHEAO5U0+6
KzZxG9+OcfItCL4n5YF0llac+tC2mTHDWfGgSp3vJcJo4YhR32UtJSta0W3Z0oja
XazXmwT3LrH/i6Sn2ImP4npAV2a5NyRcXTnuSs3pZbvRAnLh9FUYQZVyQobc8PQP
KEwkdLTf80bOsbbWQq8MJYzDXa7ekFs7leEnsJKWwTutSlQc6tLqt36x7UtdL6e2
aPnRCo0PdXAxZ4XDaduWG6F0Ual/F0il9gtokQ2To/NCWp59PvqyjIBv9h+4ovrj
NuPc4mxKq8FMyz0ij5v466jDT29xveY8gU3iw3FYlqd5cN9P45wBXEf2x8OamF8p
xsNyLGgdh2g4iCrrsod0UOHEi+ljMKqKpjbudb+cv1VgsCffUZu53STWaAYyijMv
CkfOpcBVUodrCIPaT+zPo+D67Va81hs4jezFgTBTDAH92296lu80l2uWQ9woX35M
RwqRhqoaz436ARVR47KJS8LGsitF/lZADZLg70CR6g7X1vn6lx/U9Bn2PcXZyY8m
4z3A5kOe5xW0kbVT34OcKxRwHyKlZzfN6hv+cPsAhVYFuxlqClbRaEwgxTeeqZlu
UmLLH915G83N7B7MgEdC1MapCdXFeQOwgJXOUK7H1GUOA6wtZXyApzkY6zS4AR9T
ITtId6Jh9B0/l7i/+k9BbBjolJlHc1S9ZArMCWOWnX+GsR5tiqI7m1CfHtzSWQY0
u7ADZBrQZOCk+bU4hsAiH5Sy6jt63IA1rAvdKm8w+xC1ZwxH/VGfUaotqzVz8txc
yWXJN8u7j+sU8y4G3Hi8G7sSdTqsGZrrcvmwMMcriT6sRBBCoWQpciCZsDsjJDvL
8KM3/QPdtIaRy4wShC5W+kqE0bKbTuqfhdL0wWXWBSHxQt9yFQvWSn0xEQ7rdoUO
meI4W/Psftlh1Op22AMYcZv0oBkdQa3YnDFPJ+5GF82d4yWD9QpTaR8EDiVErGak
Iv3P97rrrkpaSke9N/NySHru3CKGFJjM0L3RU3w/0WAlpbaPL1P3VNyFzJZUJSzX
omj4W1NeK6WceMpaEZxEnOB7Cg1QBbuloPNbLXM5F7fBg6S3dR5mRcGYBTkMMhoM
soQ/2SHAbOrCCl2wzrw/NjmT2RpsFN0XhSdQ6CFruvjGGb9VeeraMy+7N3QdRVWp
tk4VhbNBryTHCR4krSGJ7IfwmKtuC7YFwAklpyirADMkLy9fohPSZZk/+ZEfoslI
A8T8AByibgwSgQKcBZX+7gzDTQqCiLX45AnVchWO8EnZO+P2tuIQqLdttm32jANa
yhY+qb7NdhB15HMqG5mpHd1+y3s4KykdGDAW4/wCXBdKBlcbfQiiAEjRtFgyX11s
Kj2XXrYOyNO3tEZ9zqhIsmp9+hCVs5x2zmD8s36rhplKu//UoKJEX0aHr/0XJZf2
NncZaQWvlSe1YYZ4hsam23A1UFntzrkXkwQ8HPyChF6wuzJ9aIUcqkKkEg5ZXJUa
dHa5OysFShY0h7XN9s767lfKvV+HAF1huNSFmXGWewG3cTq/Y2iD5X4jtuPnZgx7
8WRJNBV9gRpJsVnVo8MWd5SXwQc+vpfQTZQqfiYr0vbUYViFgfnBlyYPq93QxzbS
7U2Y36ScRDt+2k7MLI+jIHHvcSXciWg90Ryu+CBWdEcMiIbTyJANc0mA2DeWA4rj
UeUAPQQdvwUw4yobL1C894NE8okwjlYEgdPC2yTVj7LJvVS5isz0TGKyPjMWNq1V
236e2fFhr4AdjTlgTdhNu4MHWDvNUaTzpzjVL7GSxARJgCbbolUIdkd6ONQKIdpt
0vTQ6maWHu1qh1x5eeiLMhniFyypsLxVDWEg0C/hR2q2q76bJBdRFGWQeD9hoSal
s7xmsUdh0NJrBNGHV7kXO0HaMsJ3DNq3YjTlntz5X+tw3FvRav8ycAuVcpq9xNkY
ZHbVm1h2hG3Y9Kv9tchFy5DK5aHWopW3y6p0Y+ei1mlBcZeMMG0rvV6VPh3xCRfD
91ZYYZQNY87Ui+lKtCU2/EGr/aa4jRpHqH24yhtFIq1aNi0FTqjykOgH/dJ5syFG
p4Uzrm/OTon6YsWbULENJJCJrE+eXbXk2VxN4yCSOCNNdxxGLTRAGhokDO0oQaQP
WsSJAPuVPdjUCsk0D6CvGJX3n6N2h+BnpsSRVBBgh6Qi0BrtEmUY1J6pJ0Rn3XYi
DJb9CLYUwZLM9U9t8bNTQv6PWRN61W48snVyZ1AJc0dNPF7BRf1Xbq13t22vWTeY
GigPSZzTv0r4alssuhlPkzrdfI/3rvSmhwswm6p6nKCyeQEX1T3qUpGRZd8epWg1
DivTsNTFcurknTrNg7zP2uqlsoSEawEWGl1mN5mccM3bq5hbExHAVq0ElJthwxzk
B5buZwkzjb6JcO72tuRJ2afpAeP/y8OgeCXoEeWPz7nqgBPsLgoFbBM4T0DNoSxU
j06IUITSzvSrY0hT0n9sF06hXEIjTPKVCMwEhriTySKnu23EUTVkqPvf7XcQkWG4
IBitCa/dFNcvmdWSk/wWYwXFBJEI5rNXZA5VESu6fxdxpFD2t/R4U5ZC9VssaTud
VPxTHhKuW1kaJnG4zzVTPfTCtSf25rYDCzGFiLR6JH07ZcLKAmQLygzJ5oc6t8op
PAe5rQ7g1MZgMB3xpmPXzkf0PjVSOiImdLL51KlPaaCu8YFTnBDTBnVNZGUgbLa2
R96pyAJeIV0KuYBMY6rWinNdRoWH10qO//fYltVY2x9p2joDI5ir8aR5lm7AV109
jQvQ1Xja8cZEQn3++bw3LujpsYJQ+TW4PbO9+qOULLeFUFVpI5abtIllfG2SefYV
IYi3o/XYd9ysoI3xPrsySgovQUM5JqTbm5892RFYTn+0kkS140WDVhaTKLAV54Rt
G1Lp349mm30kzwwEDysbfCtJ0JRDPcV+b5sgXpRGAVyyjqA7m+FEi3LAENutfKEU
NDoMKDkBNDXzsUpH3EJyNbXqKsObkzB6cBNUEO7dl/WZQjyCP0PVq0kjMjo5t9j1
GeWSPFmnfeyiv2DeEsBJqlYilyf9r+xFlfKF/6VtJQZTlAD9P88IVLoIFte+IeZ+
PPdW2UBOMzGaVPTBHa6ZRx0YEoAaOwOSnx0w96H2YmnKRrMl8nrDXocnHY/ZWM39
y6HeMtziEA2LljPQWH9CH4aoP3Jc7W/g9EFMedyMICLumK3rW2ci/rTGPtNSNuYV
BB/kJuRABN1X+5/KKuXlEskt3Z5ZoYv2zssFmDUuTlCzVne4YYNAZwKsq8tsRNeI
AYy04b2/OsCmlaOJLW2XmJkdzOdSfyySskPv6PAtuBPhXXK6m0BV5QbCIX9Pm7Vp
ijh7sD9Vd8zx5QLX9FgeXZjcPZ8TAAkcTSX/MQVtozW6ioh5Y2DoTI75woVjYF+x
l21SNcwdlzsjyfBtGycU+uvMiiLzRzWL3OxmyzwpkMywORJDKcqr4h66p54P3Vsf
xhSf38EX3G9tNA4YhR/V041iV40TFVFWeLRWBuJXFIl4iO6P1q9zYMvet7TxR0vT
jYplhLS8lpCLvPS7a+sd1tjc9mPTqVnTpftzrnCZxbedfLt3kwKFrWf5HnIwDz+r
IJGJucNPO2o2xmUR554Z3fn6YxejVjze9zgZVpmyBpT5U2BXkIUVf3CDySr3el+Y
NphIW6tl8s4Vlv5oJpnqfnK52qoPc9KBZaT4ZB4tDURut1QrXdmRkDrI288AdsI/
CC3oTuIjb8o8gFAk4sojLT0drpUUrqrL+7ygHOFCO2c01QlvYJ5wrLaGwz+SgYbP
x2wsJRNzpkOdU84zlNl5gcAdEBqLlB33hgd1PWxJbflpuj2erns0LxzwXYoF5TjY
20WefHciEwkWyMnOj8Z2nHSymWnfX4UqXgNYCOXUwmZE0KZR/SeSBIA9pE7qrh3C
e61ksSmSTgcBeaHJ2F5QhOROxDoWfxtLkNYr2dd1pRa5KoHcJSyDtJzxOWdCECJW
6TU+LsW22SngMlRyimIyHv/TnzfNaOfb6vk2aLBfoxCAgseeziA1gRm6DPng6VTj
vGtCSXjCyG1O2yEX7BwJW4ntqOxWo0LugWUlQqnWf49YkFK7F+MNgp2yzgE0TCyD
hM2Hl4b2obIIGDsQC77ib2ctODRnjfIot8tooFZDEQq9AaooEQCRS7/mBK6msXTB
p9jebbNi/KttjWxZJwHdiCIzzS9iA/Nnb3Qyl8U2Y9Q8SBewTgmgT0RjOkAV0fBp
ozdm+aZqbCbt60Iom+UlpfhwXQ7DkdQcy5XjarXBSLYgjGL+wRurrN9m+7FlVFxI
F9sd/7C573gO8YSxFbcZYd1JwlLoNpO8x1xzHXRasgQQYLBPFfvtK7a6QJcG3xdI
5F+Xqqhux3F70kzA5TsBCns/+HvBQ55GLOv/4NWszPr2gRUwIbH8JCLNfyUIeX5d
fPoHk/fr/qhvU1dkTDOaAlVq7QKqoysifg8+ssemSV5t59gQdFFCKBShws9p4lfs
20OUq/cpi64eOpxK7jZ6KCyq8qOeAY625gYFGZOABx4u5YUR4iCDe9Ok9EtLhrhc
lnFkKYSjj6CvAE2Ekdf+RBQ/AuKLKq1IOAj3CIdpPYs7rHeETBpXXLty3daEHH06
VjDPils2FdYeiHrZ8wrbyjcJgvupItzwO36h+T3EmteNwxZABr8Faq5MSGMoTN8Q
cYhLq9Le/Tw7Zjb9uIchEDm6qYdmZ2u32TSd/N3bNPMRvz3KMawH6KS3RUdFfbrV
4WgsuelkJ5xiG9+BjlJ1bPwcnk9MxmQBSJSbxMLSLC+TKY8R5espkZ+8T1SHrA6f
He1kcCP2gDndy84EaLQxIkHN8m86fBHx7epki05hdTe9XZ/IJA4XVsFN78C/AvuY
B0dnpo1ocRHWlanGXi0nRKl0xJovnP2WC+bPj/BxrhrcXeRdBHK+Upmld9HMCP5L
UW+M9KmN9OkQfhUX56oW3FpelpE0gePS/LfH7fJdftwYo1J3okMFFc7iYLQk4mYY
Psq6VIxt2ZG4csvtPPgYbF0qeoSPDIe64ov5oMaaZBYddECQonSPLU9LRBklpXmH
hS7T7rPt8CKiKvR/xaabJCxfj80vE+CuMUdeLHOzzL/U49DmPVFZSeBziLsMPQaV
fk/gAHtSSyNQxT3OmJhLBe6L+caoZrRhrl/xIhK4+vzbc6iKIl6cVrehldoRaDjR
nhXtcBeAeC4O6O819lQBhvtMPPDmnG4pTpDv4TfjfCvntCkLJKeKi7N4urLZg0Fq
mMPHmfc55Tr3WmH9tgaiHHkLuGflLHGKgTe3tLoXPxJOLYQseLy3ZOtBdrHXG2q7
61mdLPNNBA5UdlLee5JMZc3dR87r74BWPVZBBQ7IPQDe5IBoP2SuB+yJ6bE03y+K
R1ALfhebW9WL9iiUwOLWyx8FJDbH5fqdlWq1xd+mZ2PNkwMyjXUj9IuYcMEts5uB
gKw7HiGpAtX/lsgolDtpKoi7DNZSIJl4Af91NG/14+yS6LD4YIo1HwdGs4dLkV+s
mXTZwcFiBiYokRKrjhrm6yzL7kxIqEJ+vc22OLQfTLrdXJMY+LOi3e+5xgAsu1xM
feEi3uKO5DuN1s1XCzBcEFKn+rLbrDQIbC1yYaq5wB4adOa/5pDpzHTXlxV/ztYc
ISVCyZEfJxL7JEQqP2XbVXWmy8k6NQk2Nafc60OtLARiV6jJPgZcqBpN7X4GNhK5
3WvyOVTzRJoyQlycrWyJyo1zN5zwd/4cdNRe/lGBJjpDpEcEaVYfEbaJ/pQJSvHm
vMqGuB6dWI5nMrL/b52pX3XEvXFLLCH8Pbfg8Nvud1J2aCTNpTFcYBLx9P7KcnoX
SUq/HNx5qElodUQtoI5uAU5RT6waLKNynQGpKkbJzNswgfYZLO7QO7hwEFLZtw0T
70UpBwkYU9GcJm1f52MQYe0twZb/yxEVm2iA/8805IYpMiowv8skfPxt1G2Uxtg1
hIo/N817kEM+yfM5taCdi4EdouQJMNbJEDhqi3SLzqIKmi0DGeAqSVSHim95tdE6
hOuK3d7CR/qU+VpHstJrkakV7JLhZwe60W1yrH64ab/ySeuO5h3hpnaw9RN5Sb9P
Q8xx8AZfjq1xxyX2Xx6GlBEpy6s6pvHfn5sfYSszRqFmRb3Nz36Z1+5R1hpoyj4z
lH+nAaqszO5FxPM67XB0+xAIwNq6GBKk4PRKE8d31ICq58y+rSIRstXoppjxGAvE
halgbJHbG0HQFXL+vGvqoxh7d0ZntWNC9vGMaXs0OgaKWcJHVsz1iVO9s5F5Y/27
NcQA2ydzn8OdpN3OpaPl4wxkvuTemwQWOtGra4iZUWtjJYiFiltH4FFoQ6dAy/PC
/NwB8vNtz3I+m4j7dqGqqgTg+M+MeGVzzzL/vKk7S8RdxORnM3frz/k6NWuuY59A
lgMTFmV2AdPSniDHpZu+6FZE7LTe2Y6ODs+Gb1+Ph8d4KsI+udrefmqm8mcOT/0k
3u64xvjarvgQ7J6BrE3cAoytLNgi1lHNx2nYWVN5lYtu4gQ8Fdp6DbhmX6SKIGu9
quKkO07EMxVB9LYEV3459lZL/g99Vl5pYz2ZjWbxfOmBJU5ZqjvHk4hM1qIyw+l/
M1WWzEQq3Dywht8BsxSzfMAewyprONviulpn4tWflmByHISJnVyM8/9tJPVjpWa7
8Q4v86ndAAcZgWHF+E4vXjvIxaBKVtXdN4kDjmEb6i2cbZ1crVXa+bk8Lk5yMkNJ
ei6tGviM2pDlJAcF9eJNIh4xuGIKOJaHa6vM/iUwZFI2qWqbHubXM3HERY1yEF4L
yX+jUmHm3cFFEt2ndTEQoPZ3Ehx8rA16D3bpkUz1C+Sx7ilApFoEB6PNMeNoNjRZ
FTAWTz3vjSO944Ap0yKsb+dJU2yC6u3ohNb4IpIN6tFyZuBFwy61h5sZGBB3FDgJ
Qv4GmIxpcrcCj4XWAsvNw3HJOJCpBHmvTNcRECApclk3hgqsFu1r+nNxR3xMDCGw
IOdB261A59ITi/UqqCvssNQGwwqJir0TT38B+fuHHsELA2yQaYgstN7SxkHK8inw
cp953rbfNU8KPMRyliR3utlZ6gom0GnGkP4Lut1smw/5mQ3s3+mkdlrkAcfz3sn4
2sce02mNyn48BlLtq4uAT6g83GDwqiLlsFOWcMPlqTH6br/H7lYIZ5KZ2Yqc/0Mm
aW4RumUmVKKm/Do4Mpne1QkgaMI5MQQ1aCw5nw1p3ur+75X4HsjYawLUliYFYxPm
MDZFfV2h6kHIX5LjTBbYzbjIHDF3KJpZ5VKBLWI5WE2ou5VZ7htefPI/rHiCPnNy
Flm2xYPsdihMy+QupD2dwHqXSkR79kIc423Ruen+pxalaaYwXaVS8/zoLuoQK2rV
mxv9L234tQZNIcFCoZETFtugz5XvU/f4EBKJ8wxZRwmbOatzVBKlolf60EbSdbXs
qQI2Wg0Qz1kFGK6yzGh9pi6thUBVe8wpJUz3+a+lavZg9h+WxiVvn1lwg1NMa2ed
nljrUm/z+CZ1iLU9xujt09fE4VY6W9/Fh1pd9ozUvqCRPmjkxbV+KTrs1YWy5ZY9
STpvL5H8RwfyQMcZSgtw7DCgIMyZUn36mpn6Fv6bvzDBMfNjji3rgwJ/3s69gcAQ
x52/1jTOXKPLFyK+MUqcFy8rN00rrqHLMmcBe2ajEnvrz15C3Zt/kWpBbrNGmekt
azd8lGeoy6XKYvgqpyZsIACUoebvoC/Xliz65e3zbnHRL6twtLOX9Cc9CsTaC/FZ
6nQtaMti5fLbUjNcbod2lD1FIq4fcV8B19hzDCo2WQvb86BuVtLaxfrA5hmJG6IW
hIIcr2Kg1hH4Eo5jSgRlmf3hh2HIFE88cZonOKWi1onj2UfkJ6lj28tcyO1q//ab
OWXKPNfd8kiQhgIQ3o3jEXp8Bipu87E+W3Rr66/hVkQ8aRQPoqgZ3b1qJbD8dGwc
cC5r3fmt8UZS0VUscXwnKI9t51SVbX4iFc3vOvjHXLCPm/Q8BmWFlsTzoISEAlPQ
kJoRzO5DylQNI+QbAHBArkg2VRuMl6R/5TMC/jnkWv6Agpoo/bmPuOTIBNr0vlmq
c+qtoNpMTC27zkWvuOkDEUDOkq77tVMMQOL87EhgTaQgSYrHmiGtuEw2dMoZNpfC
t/cpletWycdww1llD/dhkNRxgR/f3IwDDfPH6Taqo4zD6H5CqK4+NHEr4x5a8QGX
28o6Q0REKerqRG0g0ssjsARjmhsfHu13UfNccoO/7tO3jtEg8UKVzs+1e1R5kh4S
na0b5EalemtsgclDygV23imk7gscIW/uHHvlqRsrw39tJhw3kmreljSitnvuiyVJ
Bi73/B8ae+pIWvbAL+iDoH3Px2oKO5797KWXplPArcpe6NUUsUb9nddJGwY30CP9
4U27Er8jvgGR8tZiG/0B3RuUEmd7jBsz2CcVIduu9y1tlMJgxMlTsnfdqTE/oJ72
+mijkgDl+Dx5hk8g7mWnbz7fsEkfRdIBa9rfY0zbbOGU+3CBw9IH5HfI0shaFOZa
TNXe5hJTbGwLMRU82z/DBZsz7oHLT0MyNZrRSgeE0llrQj24zX2C9iWA7qo8pAk+
wPXLF1GmQezhZ6HPlMhRDBEvZ/jEcw9i8ScC/pY/wetzgN1GkpHDZL7OL2MFyIrp
B2XmVgDbpd9HLAjE0zdWbM8EzkXGg1+zibYM2OfCKEk72yBrE48VfkvMBHojrR+h
xojLD/uxK7a4e9olNkuaRjnisPMg6j888NJnCLkQhusVtMkiPCg891RJ4xrP9t3c
RwLswBV75IdYuAOnuPviCo+WDxI4LkAw8aIMfgJYH5KlE7szK1koLXNXznhMMFPc
Rn8N8+0KopZ0SUMesdzjVAI/x1ZjY8/jer4ON691tu5Ljfyxh3pphiDih1wyjDVO
tGLrZmJuHaMtClgASpg+daFVWlPg3jTi4rUajFRQn8mGBXDKdzKwjIirlB9Z7o1s
553cRBuVMgMEwryyeA9RjewHOkWseiFIQhb5EtTlr7/tffgF5QbYtBTjKw9MH9rP
mUHfCTXtwdTXwp0OIohoFmMphWFJtT5aaxX2tGz6YXa1KOdv3jFm2vh24Z5/dXdn
u6vJLs9StseybMbFcIpzmqbnLf9NOXmNhpYJ9cRMCqtsvvwDs1VVr+E1ptrKoc+f
ebSxDKMHUzgYbltWZTRwmr4TKwxhwgs0CA+7QYPc6xEteoWYZrQiOM22Az/VxCN1
c9jwWe+4L7O+dJJNlOBloQ8lmDEEA+RBKGyP7xyvj0A4SOKd7qUfr0q6WCTb3Yon
WnYLgNhAkfqD8ks0b5QAQEsLtn4LIkxO4uLm20U0xNN3VqD7K7Qmr1WxH7tHpRrZ
eiZ1A37JfVI9+3pCocgCF/rqDV0Xw+s9wJ6/5+YUK1TzS11S5sZfA4zzy6Ad41XQ
vMkbDTrzolQ/Rsgj4tYueYO3sAcUwLvYFPFEnjVlCX2ESf70u05kbjv4UiQ05LkC
rZWlRRRrhUsmq9y13JemEeJ4tVVaKgNHqJMQu+Fc98amwNAk7UiWBXOw0xUa2qK4
G6nk/PwRebk2GEeooHfTZ+3sF1c1qNkQIhS3gJVC0u7scO0g+M6Qrx1cY3PnzFaA
zIGuM8ljvaLiQCdxecwgDEKDGuJ2WfqqaJ+RZyIrKDmq8oKYj76USb5RZ9p2xzNS
RoZDmX4//3aZlFkkzltL3yuxfWZM7lxPCRJzjRK75z8UmkfKKymzzvRECu1IxR92
2Mspo6zn780n1SNcPYgK+JvMciWNUfWgsYcDb8hPcq3H79EwMNfTD/u8t4v002Xc
jBqtNQ7M8Uk9tkkL6wJUBi8L0Mlh3vEpYKtQixrzqKg8cxV7wdCYK5OWeSE/a8YL
obsqX20gW77fpXwbcLldyLrmf1kmzCPQnb1z53WyPlRpWRf4Zgg0PTzNO7XIPju2
04ByqQlIeVovaCNyzhI55dIrn/a4ycFGATdjePOy1XlyhbkEvvFgjNcfS8onP+SU
wuT5smStqpULC46weLCt53btRPUgl62Fx5iYeFCwuxxXuXWfmY+x94+MYZtk6Dpz
P4mM7nhiz8yJ4GtPJi/PfX37CEGIf/7sFygy+2VSYPnNZUsG5lJzBwOyxSLtuY1L
mhAKx82ijsH0Bk2JKp0h5r4OykKqoXFtrwHilKcuHkBvuAQjkbpPuAVrS3bArGPv
kYI1IFDdxcb6YbAPoEF7cy5ngdIAAjloBjR7M6tgA/LjCBcsAiWLJGPhrX1ZZ/lH
ZyRdZtVL4mIRfAJbibjQ2CfdTDFxJD9IKyLVC6S6lvFRKE0xm8hHoj7UaSnF2d8a
6/9OQJ30mn+9uPysfds1WlETAWPTqehOKtDPS73zGzE9FQppBxz9/O60xE+IHd+Y
HZVafDLUBjO87bBQe3FCYWH7vd9OUIc3a/5HuH3fjn8FfvmM48tFgEo6IF4y/01J
KGQCSOE2Css5N/kGSWhBLLnm5Xj+Sp31khWJ0kZISjYdrY9efdbRnMvrQYDOTq+N
iYnfmso46VKEM1kKGSDj14VjZ7qCfPi8NnWxez9bYYrMy2/HBVRvbO1MctI2OLIa
ot9tt6jJ/IiGqhf+CBRKmZk10vn1/s8TiOb99ZIPQis+flAwF9czaxtAK7me52J3
Bb0ujal0vUSdBYyhfLoknWO4S0+XGqawr7NU7jWczHokbSyRfUqISnmYeQDOnX/q
zgPEmVXu2XOi6/qb4mZeSzG4sKc2GDcvZOYynoiPpffNOdQaJn68pLLVTDNw6veK
vJ/rfxiuO04WpLeqTmZyK9MytbaCWMT0WcHZrMRbuuMflpw1B0heFsLTCMc7qK8h
fsFnyLXaeqGtcDml+gZa/fzGLkMRJmg4Um5BuujM4D+BmrGLMgubWzU1nOf2sjAV
mH8Kez9KOH6VWblh/fOqXK2DYTndpFBgaxFxB/KvLqRne20v7Y3gWwCUcJs0Hopq
eRsdvAPjwS4XVH9KyINOtA/bzgumh7Efd2pWhQ8WpQXCqV9n1KsCva/v3SsRW1fk
AO2a58J+UwwrDvllRcjvBypb7w7nFL+Dl8p391ihgczgkHXmwIJVWrMAUwQuXCkt
wLvNx517JMkVpb7IdpINZJv7pI9a5vVrnIcgTSY6+/SQTmHv8WFHgSwrCj71w18q
eTMzxRVy/t9t3Lm7bQ09DX/dFV4eGk15hUIstpbHgCH3JvIw90Jsh92pITFmNWd4
67MY03XRoHoQqSzAqU+TgNZ14AHIlkKnb/CjPuHHmOQn28hhicIdV9EPSPUU34Rp
5M55/Qc0Fbyp7CcuYFdA1MkR9vvZj1DEFSvZyHsrZwhNbTuvK1PoR3n8D1Vx1boj
JJgnKaQnxGe0WY00TpPz54k8f/lzPaRXCkvM2YvBZjKX3Co+99t8YyXM7W6W23/t
fFPAjvQWi1PHmRtCb4Zr//zoqbGsylyykIqUxpm5crsjI+iaSpIbFU+if/FjyTCt
7OKCSJYc6O7+LsM29hQOFRAmFw558yEHWTq3HwjfplaYlVFX8opEZ/hujKzmy00m
QZBUOszY43k5KdG/1GOqP1+rnSG4Sd8vCEA3rkUSCbctYbX7w9BI3fZqkEhIGsip
aleTVlsCP9eWrgtMcN8o3PeIicwmgGfd1P3+AxpHTucXzRFRSueTE1LMQvkk752I
+VIIOInC2oLv1EgzoN9Jre1OMdtQMhdOSQLzvdsSwr2Sn9JNVvVpi6flHsvMfh5Q
Yo9fRY9zv1kol/nuLPeq/YaV7yrmERaN3gNxsBDhACUdmkF4EnDTCw+jJpPs5Yjz
OuYM9ymiRM3qSpvqsJ52KITvWmAtoGLuiNi+2AXfqTBZI84DHz38S8Ib2rzrGyAn
rmfIYWGHJFPl+ab3c0ZJsAj9zBGLg2fBTbwlMv4BJX136tOqpE8UAQummhc+dXkW
WmsdvqI3eM4/ttKIRd9bl9fBKta+15r83YhQFTaKFdfN7HgxtbYEUqSfJt1i6dhX
30Qt7Be2CluHiehRgB2nmvFUflbF+EMEoQfLa120badxSlyrSOKOJhXU/AqZCWlr
EyBYx1WmfISrr2ruFBnqDltgUa3WerJnpUtJkY68xG8kKv8dqZOM32IP6XB0M2fH
gnz31PAlKzO5LdvmjLeMwNnREpk2WevU0b67FlRD+jO5M8Em4//ZKJZRA9ddUuaN
a4Ksh3qyMrDx1dzvp9bSKJ0w0RVpM5prMUgQKcxDzOfMgqcOERNSwR6W/VRrngR0
AwxWVqUJnfvD6tAXPVQxHly4Lh7Gg7Uz/wQN1bf7OWsWoO+K2h8BtMrrfW0Hzmt0
2aLofI0ip5NrA8LA8Tx9AS7Q+QLegZihZ73v0jkFTKQSF5mdfxQaDN6DNhbKCoEn
DnDgj9b9C1bR9JeWPSpLUZwI0QpmjQqUZ/Fs9Uj5sdhk613akcsZWYSTY+jIY+8N
5wWjUUxT75PM1mlYzRe5RrwEa5wm4wRryrU5ZiE2gUCcR9Kmm06IQ9tcldD76Hd0
uZ1kY/hr/pImlYp5spMXCFzWYgWK+7qYvVIWGVoDdnURBv8GfoHRsZO6d8uVnceB
hpioRIlHx10OSAAOwt94/C7IE1D3byKXxydwqPJzIkKPsXs9zQMZd4o6DRW7urm+
Itv8i1iLm70Q2Y3z6juDtVhV5IQCWfpSx89hk8GzH85D1zZmm1u3LzBiprWKhseu
PAtIish5D5k3gvKKfB7Qwi2fRxvHTfuCNIaTEmI5aO5osvcekwRv8ru80ord2SlK
F8B7+Uv3sG6TpciaGsHcv5mLW/egmkiMrfG3zPS26L08Ep7C+O1F6e2vWtSCXSwh
KOB9bOs+8ZnEDzFu+/os3a+yjrpiZ+amfhsy1ktoQraM+vA/pY2BH/P5ke9zZOt/
v4Fixif958jtPXc4VcIg6PvYUfM09WM+YemkOdHndSGv2nVVY7BRS61/FbUjEy/w
PYaN70AD8sD1R1Cm/iFjbWCBeuIMktqTzqR8YCh2AIHVcFymHjGdqjdXhtKfmmep
vnI8PQxipH7gKAxV1W+3+V+F6gyu/BudkOhoGCTC4YzuoBXQNvP8ZIbgcKIIUs/M
pzX7e+m9ZzIvOenIvxJEL+v/Q2/JXO+FnSZv6uu4ERQwXv7otvDnRntcE4QdQCTj
fHDC+FC6WVCVZBG52yZh7fkmxy0lICekfReCXpqSQajta1Ifuy6y8CMdJUGGld9s
wKBDEPIvlkjJhMWBygkjhUfmpvuLxdtoytczqHdCyrVNDkENMVCK3n8Xdx/R2/qv
HGnLlNZ4X0lkZ9WyixMYJ5xJ4EKNqJjiYaPT1Q1ei0B5vWVc9+CP72G1bOgaY5md
IDM+Hdq9O9gZcSmqXakc1dsIDdgGIIIP+chP7TRWcSAFwvWEMoimmW12nMfGbx+2
vg+CQxCNcN9hguV3M7+DStGCgeSfeT45dHrGcvsQyZlClPUZVpxFCOvSTNmKA848
L/6kTVzO04oE2J9UQ7mwXOcb8IuCjp/I75YDSEvgf39hKJ4b72RKMxSLejKQaLDp
YQ5M3cIJ23Izsk48UIdZNbFZdZE2fY6TM2sjhamLlXO66ehEDOdcAOUiHJO4hFL3
UoctBAO6+d7Fsay6F/YaUMaJqrE3vlJBoX/e1vi9mWTGM1flpsqLsahXe4YS6Ks9
jMhEmubOr+DgRDgV1NY+UtRtIZ6wlhJr8t1HcerFe9dR05j1AwmCQQhO9Bn27PzI
0qvVZXdGpZgWMAJS7GdiujIs9dw4D1goG+sn11w/zVKJtnMWIj00VowFvdIZ2m6R
rC8cc9H/SpgvR5SXcwW+DF/oxIB1aZEvRAnOqFS6lHli0qeD2wZe7GyNHPFJasLy
DPRiBOY4EInoTxP7rvTQObdFaevnlirUyMcSx69dJjXO6VinSS7gzxW45D36pEKr
oJgT8SvxGeB/vgSejMxPdZPGL4wYsNTVe2Vz36k2vIcoyY7Nf9eAoh4FDFErWdvA
zgGQxxJ3vgdFRv0D3O8CEnJewOY2xsBjzLDQMlZCUVpc7tOINsN41KOHPLjD/I3M
c720rElkpDbuyEAJpMRMZkepwQnk5XOBmsUqzalE3U2A20VmYv6Olk/ZEh2H/oVB
QPEKOVuykHZg1pbvAxWAmxZq0Qrw31OQRJ94AQKICThsV2fLXy4KqWErLgyTCJkK
RhNj7MLZj/oXMW0yzaxZuXXq1mc34q06TuAHpX4nafuq+BRkokAyastp9xhHIc3Y
9Rf3A9hFGm+xRBByhtV6FAN14ikUd/OfBKeFfFO4WrsfGEUbnHqa+47c8B85w4Al
CGFrkfjJsYJFfUUJTlwWmST59AtF40Yris5MLdXNVdMH8lf35oysCSpWl/FUNO9f
Oipsk3paW2jOuW3pr+hluWPc3GvEehRaC2hmv317XVfliHHWKyvPqcgRJPvr0eIO
X3S5eLu2zqyhcyFTDqeEZfghdlekP03JOTwaUArUwl+T0rPcjc2iNTQ/aTo2+ihz
GgZUuk4yfhuccovqbiCHMmJE3DybtCwLghuo0eJGu85eaOMmrXFwVKWCLwuTd9V2
dWee9qSY3Smb9WoU3gmv7hFfqlwiCts0pjGWw0t0qX9iuSvVkIQOcPjSSJodNOnM
HR5dq9y1C9CSnpvXBogUMfwWJ1/8T2dTlWZcDVJZotvv+I33lOmEVCbblW1QkDw2
gMnD2ZQF0B9WUA6kn6K4OQ9jNLXfw7SdbJ1O+78N1u+feB1se0isPxVQbwn/ZzV8
v+QKkfal6iu9CPLW5pxiSj4BoiE38L/zOK09rFn3BJ9U8OCI+RW5XSvlYVb/NEH3
XFSkV4OqAFoQdCOX4eyWNKsH33WRZNn+6zzFBVFAN26C4Q9PAMdabdF2/MwV0HcE
Y5bCMRRhY0cIgB5a4pelEBrkRNJywGGgfcllm6nDucECSt5UuO6v9/nyhfv9vYhF
hz1uD9zKiNyUs44Az1U7qCQgY1M05Vl9dFqpDhR3GNdtaALLHeWNWAJ3NLxvaGNf
AS2tEGN5/rpWq/6lokhQDKfu37SXQm+jHqkRcbn+k8aYq8IlEcEMmdRQUydl5pW+
jvNeLujpwNtYqhhrtkf9ZgY+wUf9vfPL2IzpHMUAS5v84notvEAHf431b5ltX5PM
FIwtB2qFestDfgigY1grQzQrXBNpQH21DEigOKH6TepG4OdODcxlQ3WSuhwYO9Ud
TLKXo5jF0+RWHUrdkHdpQ/q9r90s6JIik+ALJQLuy1Igygr1vMXFHv9dLZG3x3P7
tP1T4b0C6ZNXwx/askwtV2n9/9NQBSWj7yF472cp39RLH+pIacTL6mYKiibIH7aA
N7fqithzZD4cWCk/BziHahGXGJuZymh16iTqTMOCu/0o6kQ7bu6rbesg75JBn4uG
StlKu6F31tLBkFOnCU1cBOlF+dqq41jUerdR9Dwp6zYEmy87SiV4mIl9I7q1CsBk
v4asRvkONBYdfjh7if51Uhyrle78ixFAmiFe5wfH1JaR7o63MqbQi/JeiCe3TpGw
BqD9RRdeFAJEb5RvOTBMnPYQO7r1Olrb1PMhn4oSim5hU/fZ7QAEeVA3QIgC0Ztz
OTWuHBr/FvieSMb+Sg0iyFKTKbK8awB7hdjOlvb1DQEDFEdUxmWfYjGK3FVHlGCY
wdIerjvDYqHor6wuC4jjldPXRn0FLm4/6S5s+D2H+Jv8+G6jZyznEOkqcgvQzuTa
LJdezlKHAbswYZPuuDUN3BTt2rF9Fqk4KnV8foPfKVdinogWCCaTRwEj9RTEos5j
XueM6th8ZWFdLbgrrt3Kzn8nAIZA8dHl9WnzPp46jraTS/C3TI8dCt9ynZldhryK
6Aw6Ym9R3iZAwKhyqT2rz0x04+fRltu/Q9RvIAt6FkUyIV8QVBpcXhhIJT6EyKJs
p9HmSu/vfxTq+w0JSf1oQnIchfkGw/pnrAl8N6FEz6ckBBAKMHUWvXuIcYQWIjOf
B+AEFyhFJ7Rytdx3wxUxN5ZTd4bj3tCB1KvY4YYX21HzRTBKYVTYHO4R7v12EUZv
x6Z8UnudMYPwYwlDB7EYa4epaPWBocrnDZ8aU/sag9VRh09FBuzjhW8fgreuzgkL
e4hbZpX3Am+Sjc/yjqulLAgywpUOCaTNBJcK4cySyP+SyG9dE80PR9y6Dy3GDjfj
ZVuQ73NlRN4i+q1iQDGWBMhH/r08zLMvYDvZgLVuGGeoen4U+oMWr3QNG6wcjnNU
C+pNtEQwG+Ngve6yzTMWEnu9SSV55pUA5dMl0Ycy5Hdc3o3+UyFpJUS4Qx88fDq0
aAUSN4ymkmg2r2SDf5lCqddEmN9P8nXgMr7DNeVEaPQs48Yq3sRTKpfPqkZ3Wzei
33yI/DqMzrJbMrOIQrQ49Am4rF0EIm3AM34ORbk1pEbBtCYcTT8f3rxR2nIWdq+q
iOWdSN6uLsw673ObCpHAinvMWn58eL8Ty7zVcDsqsCV+KYOXSCYexUhFM2PDN1Yw
whsol+wNxEPWbg9FYCe1WIsJ5WSp9M9aC+k+kAifiNx5mSAQpfHtdKHXtPSvkdYC
zmVde1zVV/3OmBA28PzLLN59ysERTkVno8r3EZuMY8f65u0KRw73Newb9SyzxVE4
BOjJgHbCYwS1SYDr8Zb0ouAk9DcSkLWDQEsQk1N3V5jI7fv+TqrOr71gBr3tP7LM
wgOO/OuSOaKlFzSjUZ8ro+RgZlqLeX1hOlXSYVS8EcihAmqc/gQ49yYPjQFX7tYK
A6IQmE8vm5ope/SPcYdILAhd36etJ6b29eognoNuUgdHhXLgHrfghP8i3dOFvjob
+B/C7sXisuaWogDv4CiGDh30nu+ry0nHFrPrHAZXrKKvSvWwUdNJV/rAhdCUBi/2
5hFlt9ASTfJQ15XW7j4FJ35V+b/BI+muc0E+ddlc5/gHHaZpG3cVu9rOBB3+XuEb
d423Fv4yhD5ykKI6NQjNyaLKc0kTTBxyv0bg/GGwyise+UBDSzWhs/gCfhBKGtc5
WSanEYrMhEwQwPEWWiWbiGvm5vwlDmZER5VLNWc1czzBvKchwldF64C45ACpvT/S
m9zYBl2p4PYJpuHCrzAk9SVMarqlIt5caRy2V/Yi+ccCgLcVghuYlLQBuZ8z91/x
GeY/iDUk0UP4m5QH/WxbtdPyYPpu7NtlCD0rT45FtCYMwvJiDmcFU25VZwqZlRpG
DBqrjP9kMgVE53ViSUrwdNBOPyQ4KaICEdihUzuY3WW268XGYVE+dm+qyBLvNKgF
Uz1V62iYsPDShkbzunrngaFMy3Rd3Qd7RERowDGSuUhG8pIjK9g7ED34S+sKBY4E
HhwDv8JAu5yHedfJ+xhk0WpZ+wNDXIoK6Sw/X4sJbUOf1dnEeeRpjsBlNO83sCWK
W9nKEm9md2l3khFkyXLheyqpgioy/2QuXmcj1P3kV3dSa5E/JtAiMkBsZ2w9Xn46
RWiXntIu/eYjDeAiPNPu07lX9fd6DHcQMhzSdkTdC50YnBkVz7omS5Vjd/yHfYB4
MehIv2236jw2UdnCSbBkmJE6MxxJX7BD2Ogh/sCPjufoZvOmOVjBN/NYRcU/TfUO
bZwHs7fQ918y2BrdQCfQ/v3ZMyc+46nUtZhyqogfLn+ynglyPuyhmxyE970U2r2Y
tw+5fmdOTA+hiIwEcqzcYug8eYX6aKNzdR/R/cNE/eilAsF9mE7jCjuGqoZyOiK6
QSpUUjdGAA+TMCmK5D1COISkwTSDQelgmC0JHTOuZyv8G3mto8jfbOOmpK30OhfO
gshHz3Oum1ag6BIslncK5aCyXc5E5d66agt9MqKSZpx1nRd2MS80qhtBVX8lDOZz
HSprxwisWuU0CHvfMymzRfZI2yyTdCtQxl10Yckc8lRLdRhzOXWmiGnEewPHvOBX
CLMYVTDJPRcstpXTIUKO3HxvKajVqz7OnqIvALqD3bJbDEINEnqJ/V24JJFwW2hO
hBVC0/gT8yeZpFs700lJvmAGN1Vml9jfQwzEHjqJVOdCRMKdwj72a0Dkg32f1YdH
H0ggshm9v9oTlwmPmBLMljwXJe+8JD7LR6oIDp7zzQCaq7pTCRiTX2uvl3pufymQ
PyM2DXB7rszFdnN+6G5rL9iy6i/+WcB4aE4abqd99aybyB2S5WhyIFrHYXnZJDcq
lndRO0YRpdMCVcq3zWIKwIQIMMDQuPLCNFICfA3x2fxn4SL+S748snh7AgTOS7Lo
HoR4ocyyOu9cg2JGuW5m9uMUG5/imZvVYHj4Jm9JO+fMoYeOUA2MDLQJWqL2Uq2R
T1cjbc8KnMeZoS5N2jZQiyl3xPRfLrskNmcKyCDLzJVFKLZT9KPVlG9FubULMny9
Ha4q/lX6VFNMca7piOgCQtzUkgG6dvQRkxLRomMyYzP7D4RikTEchd9/9OP1FYu+
CCYHFsLQ5tdLWexINDtTnn/cMimEaywUXUM02idNqKFCg3m0vOxV+52N/J+tUFGc
ovOc93QgHqTSD0O+s8d6fYCYcRxAITv3qsYjQJjhMjxqbkwIFND8Kx5Cp802FfVE
PVlqvhHNmyadOcRUKF8wpIpefb21PbxRXywgfpDzrj6SzBFKZRnoOjjinLIz6jOV
v37n6JfUol+Icr3Cxz5KZXbXb6urzVuI0H15brD5e2DJncZcvLwPA0VuLb2eyNDA
gOsW5R0Mg4JcTATlAXRiIT5h1+KNX14THlbjI/Ftlh6wZnWZAsB3OBAkK2yMBn+g
1FRRAQwbXXIK82WAGf8hmsBuJi002RlR25LS6Dbfj3pJc1E6lEnRR64i3w05B6s2
4eXcxqWZbc4DUt6tNACaycZwzOkGP/Y1OFqf59oc0ri/fAwHSdT/hw5cRWhfEW65
agdINVW6Lf8fMzkLCs+QyQhdUuHVd2M0ZxmksLyQwNhq34TbnwjJwYDrBvKvvjyr
f26aV/wq9icx9VWfcWS2Ay7Ppk0sqiyzna9EuAX4zaSp1mNrAddLciEWmacKgk1C
HY0/aPITnftVS0giOhZrvhBbXNjKIbZZCDnhUDSqJhZMamOfsXq02/PBb+JCr79G
ICm6S3M+mXLfMfTwI0/uC++SOVGSeDZRPpnDByY72MmrqZecsNCssEEuNLnlVNAv
CCMH31HM9bgee1AbAMn75WZbhP2oxyr5Onh9Ug7XsfU9YVahCChYWNPXstZo9dht
b7csS3xFWH7XA8lMT6PkTdBiX/DaV1+E6bRY31HgC0jTnzDZo0/99TXY+MSESFgg
qtyowcz2WwGH0zqdTCNHVoo5+EYlDdRsZbMBoRGnDY2e8qZaGMKrxSylad96/t+X
Yz1cg3Hm3njxP/nEbb60kAcv44GZdJ1HbiSc1ZELEGtDmj63o6NZAFSavedr8PBi
0ImtqQdND/JMJmUFrYEnovCfIJjHgP6XfS2463yAO+RpqPfB6K/9Cz2Yr3UdG8JA
u2F2vyfAXrflsWLZFxqdmZdjfXRZISyNZZ1tHZuFI0LcMDhyb4/097UrM4TiOOKT
16XiHQh798Y7UFUqUf/qsLU3iLNJJMJzb0fjVQ8QFz0oMX1AL4HdTC+3ZwO9HAEE
fAO28SbvhJraI2a1KoX2EXnebHl31q3RpiQ1mb0CaqjgO5a3Fow9OHVlfQ+wPCxg
YBJrcOahha8S2P5qxz7Ot62zlJEnbg7hVstr+XMLZ83WNvEE9eHH7CSAhN4HwW1C
IqRWEclcv2pn8J95L82QT+1aedVQRAiaFD/Z9HcUEKnYq/lUtvHEQYBms+Cp2toX
v5jUCvk/KQvMY2cFphy4BFFFrQaYsjp3kVY9gMI14d1xdWvnjPveKO0q1Q0CdMdq
+iAmPZK0+4YJkH+oOH2I9GjhvUw1M0stYVRLOfOKdZbkmw2CtPS2vTPhKjrPjc+Y
28/Ok8/eNN8tUz3oC6RVH5U4L9JeJKpgjdSMFwGYMbussHMA9E13+hGbWTEGirXQ
UlHUAklbC8yOL1vTSlsU1o+bg6Bb3WOUJKamykVx0afcSx6wcRv1O7x+MaPBJ/NQ
iLnyUyCbTWqf2DCpn3W2LG4d2JHc6TdEL+t5TO4yMOvKDoX4DrJAFERzjIOpCGcW
h8m5qLhqIotbbiMHXkjR3nAdJzZigJKfWauKZyBwFDZbBj0v3+PZ/9NtHQjw6LxL
FuvVrpvKT2p/4PfPUccQp06Q4+u/s8MGdlh2F2YK82ZiRViz1yuEGISx4FljnKgn
pYmQV56KYOiqGnl/PLJ7y2zrxqwsV2i6wWEc0kRepqrLAJkVAFixfJl6QvgzEs+m
NifAEj7OjjiKdq1W1lZ9Ek3eMKfSFlqlqiKcrWeR9FDKULkImCAda/KsWcOAIywy
D6W+klYWUI4QiPLsvr24xuu2PG0TcG7KFFcDnDi+q8MkIuxhbK4fUlqDpI5zXnhS
ntqm9++nFq5b7ux0AxWtqlC6AjmTb0nYplojY8TqVITw35XZo60kwbVYycfI6UhC
UqhVO6AhGc4oTs+phcmpl6DG4gt/ktfePqTB/rCTTT1933PVDWNR//fOEK7hRwXI
f1XckhmF1ZYETwmSWIJSFE78z3s6AHYNQ0nJwtp/N6B808ev25FsrgdJzmr45U+z
AYXXxJye3aLsVSeIe1aoa80KesgVeX83hsTDTvjQLxWyweZIG16cVfZkA07uCVKP
8YZxzg5mSMr+L6CQT3FNlO66KHwob3eGRkxXvBR5l+UFi96iQKXqZ1JU21Wph7D0
QDvaqgY6PCBb7E7QuyAizVoUkuwDXnYGZOaBhXZB5GnnrlLMKTNHnZUUTZcYh6nU
4kXYrGc/KJ1OhBriFzy23wD/dPSQuUs4w+J53BCwdRciD7+b/grFca6C4YS3DpRP
hc/5CJvUJ04nwZ+4+1Z/mDVs7dYPjINFDktxq8oMlzQv1y+Sg55D/yiGV1PZHNHb
I4IyA+WlIokvWlocAfpgmLaS2jCoqzeWQLik6T+Ad099Z+Wza7BXBOiICRlkwuBb
72M+CCNHbfE6to4m+iDKjgOXIlVJsTMRruNEWYsOYYaQdqq0VKUUUINeoaawfEL1
li4ixhiGcqRYVnCRw/WxJ6bdQ+A6ssb4kLTkaxfsjgC/lvkmLWcstWkL4XOLlO+Q
LGgnb35IcjvU/QK5Bv2R0AZcIqcHb8if/W2KBz08CT8eODAxH9JZCXa/ID/+d8Kb
AnXQpLeVFFvfQ96CcUY/QZdtSRtyBFLpqJ2VPDT2nq9aB3BvXocTXOxqrZHV3Gbl
fs3Wy9DBY2stFZug3fCLQGHMraIh/B8cnLZFUwTxm/OKACUhPjCJM+1OpvLAyIhX
DctslRy+WPD1tR69HeFbcYc9t4ZfCwM+3DoZ+XA03phztNzc97Qtpyf+6YWWJNDK
TsaObIhXctsLllvv8MXoGk9JhJ8LaN83AEIkFWv9tCMuI/1AyupZ2INKF/gxQ1UC
6+vKx+mp2WQJAT0aj5POxhhWqpmQtdDzbn5HOOw5yEkZXrmRClpXkQXuftlq7r02
Ao8+75YxHoQ3nowJdkDuinExDQIsUiHNB7AMonkjy9PzYqY1f8PY5knaTD4IPw7x
QqPTgAxah+URH2W7UrHDq68kzvAmpYF7mIu9wAjzMl0SgP8fX+/dGQHdtgLsz/2T
UmbYqPpwAJKExlJHbbBt7o2ZeoKr6K4GxBwjfsBEzWzMyz3S9nZde4Fz9uRGm+Lp
lPgxqIMdZuAymGoErueJL9sItNOiXTRdC/i/FJm/FpoJbUaRvGkiIpkqQJhOboFW
0aoA7FVTUsj4EuyRZQU+niF7yvhYxARAYGbCurIirhRtwXYH7GG14wlcE4gQJ6u+
ofDYT2/Ql2fC7W0no2m7xXxCAFlffQXXwczazLT83N/FncVGaJngb8HjvKIakwPx
mB7mPaSKNkxxXE4/zTkfGr75upIrO/+dd50T/L8G41RGy107AgwFDwni3rqPa+tE
yIF25Y0L4zGGf9NTUcJRNyIwp1f95dFMz6YXgyu3Y04akuRLgD542c9QStBTmBBM
TeuJyUeWR6XCX1ZAcbsrQx6tnZb+bvmKqgskqH9GBXamn9V9XusIAtfhL9B+Z5Pg
fuxeUsydjwfMXftAh1KA+/6dr2ZduspOBy+98jA54t5cltQJfWAvSRD1ZS++D7Hf
zahOTXOg9ENvI3oErBzYMtF8PfwYql/szysLMEHs4O8/PaRMSV9H5TentPiMQlM0
e5VXGio85VZA9LP4adjZBiqomlf3HwaLhNwTdaH0qE6gO9TF2AFv9SRoI05Zlqbn
TOnCZFlZBtFC1ozEsxcIMUxtQPSPCsy270XabRzdt3akS7IG6GBfkLtaVnvHx5EK
tN4Kt6Oy4nqIh5QXVZ7cyPIwFdm/tQysVAa197lrGNFhYV8TPHyjGJc9d3xJrkXY
0d5z0nTd+q8gR3EWTCQTYfsuupmItqeiIRReBEVFeuIZiTludApby+uYN/lLsTRf
mC3U/5UgCD7lOvJleQEfQZH6WcVtXR2Uh/LXrf+zK6ICVes8bMiZcRx0L6htNpox
+E5Eef4hEyJzkMWkPWR5gm+g80FOFeH2ZDwltrjqN0mz9+Oo1NSDIsMMo7ZB4LLG
EzSVbLLy895YkTTftYC/gtxDUF6lanQYP7hdNhQzLwwD62aNHrtUwcdevrXGZOT6
a27aKTv2FF7VMF85Cl7mULxm6jKnGd3kvJhpMwBQT8vC8+gt0pmC5o16aGsEJzq/
6k6Sn5kwAIi38WgdogHO1rDuo6roiP0OIa+KeAi9j1uegHu6+S1RavVHnRAGVROu
2jNWrtHoDcZ6IqcluqLry/JSCK2z/okIYqvggPjsUb/2Rm9rJxVhD2aDqR7zcTQ7
bwGhOvrHqEIBiDeF0rTyIyaA5jQq+f9ar7BIZ7AqKiOEFeUE9RJ43VeTloiERun3
BU3yqkglwaeIGbL6VIuAKv+mMNKxYfWqoYs2MQj2619qyLYkjUNvuAOj3/gvretC
OZ8uUsEeXpuss+ti9PrBuNbMew/U2YbiEvobdBYCcQ1dKOzsrJWUoHQa0WvRN/Dz
NiDnDIP5DyTc6J/BZOt/Y4IJ5oKrNxvWypTYz917HwiPhCvQ9jiZp+Y3h7Iqm/UZ
uHuLKiH2arOHdQUKTOkbOJD1X57VZH4IwFykcSVdYpS1pD0c/WzVx7M9l1QdB1AA
vrfNXaPFaN4rPNwCu+WzUk+G6f59BngzVW+A2BcwU9OXJevtDtr9gxqHSODie/vG
W5GYB8KYACFlPenFDNMiQn1OsmVk92D2oDJJL0HdgQ16toCl9QmZA2+/buBJJoGR
7VS81+NJxKkcgiz3MM6JpO1obPl1Fd4TD5jbH4IQgEb0Kb4bz3n6Sw0p6zK2kO1g
cQ6SMVUQ59g+BFT8XpqJNhjUcxYbJHwMsSE1OpFrJa8IVRMjPlmzGe8BsnAslxSJ
Ck81W8ig1tO18WG0NLeJ8hpmhG4mRg9DMnqWzLl9u87gMYvojnfqa5DlAHWo1fkW
XtTXiZjs8IHeK7MCybQSuy4QEkxnIEwkVyCObOAu5JPQgPf6Xhukvz2FIN63n0hW
zGPUSFKG4PAiyM+iciGb4vmi9ZBklBoKQR6VpaQYiLdM3aX9x2pIUNT1ptQlV9Rt
hd4Bqiysgp+VqD/Fi+8xtk0rhBil9VOFfCCcX8pG+eJFZqnrLHi9umGMehTHxz4S
Ve7uSfq/rkkbGph703n8Cr593e/XpBnBSU3b6d0tZLb0gPBHE5H1FGACceYi04NS
zv+zshrrNcgLei1unIoS7lp8uKGmu1UM84DjWNlqoGgsj6HgfHhnsglpK+TNIv0a
f9k3H7TJA13Y8vRDTGP29fDWLUW3Ubkihh/QDJCqG2KNGChUACz/BSPrzRajchhl
Os75JgmfzxGNPVqftoWnVJKJelynUIUQm2Q2gJPoy2dvJnsk46zxPjNYzIxJqHtq
Gs9djx4uliGeE9IhiLxITdOTpvDej4ckcsuaVvYhVp8gf6UVVO+A4vhVWPuQYYBk
ot3g6W/PQEJgChuynBqKZWsUT+ML++axdxrTP4A07d1tZMh9ITLPBfyQ9vsKwAh8
Ap3WqfAxnVBmwlTwU6S5JDdH4VxHjpVv30CWfQtcbEqI8/NiULG2+se8HKEzNtYj
1CLMPwAPmcuPRWwEB6uD3yM0qHJjno2MioV9j/Ya6DI6KnMtuddZUGTqgaLKMvaF
TXe3B033POmsj0vqfZSlDgNnEbcdZgXOPFabKOkhnMfK3oj7jczXG3NXx8WNkDZs
VbptHZRZ3QEDHrP35h6XoqvchKxhp623ckHlOpp6N0YvzinPCI56yhun+Eq3SPmf
CRpe9agqJnDbh+PTB8soXZyK+JOnXry0Z1MAnwHAJuDTTftQuD6w7IZmNeHL3LPy
hEIyoU2FrQX5kSXDHpr9WoE3Q2g/iMpLRJUjFvk0NfopU2DR8p76oyedb4rCPhkT
aho8kSn8AdDXxuOzgR6cVqRH6BHzBnnvCZv5I/Q3jDulC6x9Cx6GD1qVXJcAtMfV
iot45H6Nr5BxjxEx/I5j6fom70Fsej94X00GdLguYlCxreN4H1baAMLQIBg+AKN+
5IELEZvoFaFU5gESP3QDm428c0xNv7WWfI9shbvsOMQPDgwF6VbLEc0DW3NkuLSu
ZorZj4SI990AEeu6x15dCmedQggcNTjqeq5ImaHoVKrhD7O3D7nB4dQutCHQXF52
W5AEZ7mQ4k6aso2sA90zQ0QHn8E9dW1RzPlIyzKz1EWwJ4rA5xA3bitk578cC88N
PJhllm3kp9cy10Jncewk4/GYUbr2KLD7yaKMgmPrVdP7X5qEmxgF13nFAWPjN/5A
JAerYtA/nZQ9n3qPZ79W9dB0CYdeUwatwB3Ts5StSOXBs6T7AkaJQNH2OjR4tWmp
O/Dl/a3KyJ6jC33XiHKou5lq+Bv8umbhq2fQ+/CJGCZq3Lh5TA1MaSvbrmWJ5dvg
EUeee8Gb0UTtw8/vpo16PRKXF6XzjlWLyqoCpbK1jHLDB31Gz6vLNNMNsbxkdBdI
uT+0dq0BQYyT8MskX7uE9KKL3a5jfJRK+cKJ/SCvfyR086myYiFljL9mTLI7/7iN
4IXND6ZSvHhZHYKAO9GXxuksNj0h4Mqn70qO2yLfY3wU+t3oIYHxr7dg0zKjMVsE
IcEVGnzYL4HSETP33/UFg460H2FhKeSNqoMMroCmDCRq8TJF3SpRaRMtRqQo8DZ7
3W3ehkymXI62SuaL3CKLFum4lefTJMd/mUqjgj18HmVaGWe+I3yuKzw5joIW0G2l
nvT24XTu6B48dwcuzEP3c4RgijqmZHokagv4pUQzjvj5hWlhu5Py3OLPo7cnUbl3
S61oKhyMr3pFWV/G7vL5Hj7Q/WLyfJnTDT1I35nwY5kgO7iRfd1zxMGf9h0FuTv/
qlVznSJigtQGXJlYL+kVtoQyJS4A9AMEEyE4Nt1A3iJpg76m41qI/pLLyFrJf7kz
ZWBkgNaVt0eklhsH3sHDZ7RTolA5XUZQqWrrm/A6R6xRMRzqEfynG5UhN0pWlsuY
HVmK8UDZPz74TrNhbCxz2jiRToUMhBu8NoKODAQp/BfWNxz6AzFFDTM6B/CLJGP8
xjgu3HiQ3ll/+DyKPuwcxJM92lvMAx727Ll4CT8fj8GOg8d1cBvNyzf32lFWuIQM
MXRfviD0N4y9mtW7UH1rW4m1xVNMyoiOzSNpHhZ/uNWk/4yGfc2LVnxX1mkl6h2E
uk6HnmEX2yI8ypnKyIxQPPBOol2zfh5EkQZLan6hAC8+FCtzYyPsLHy1Iqavh7Nm
JvuQLU7jQDK3RoJEzccw9u/VKj6f/SryYXc+q2pbdlpE4ZuZoVXZzuVUEervciAE
55Qbc/vP5M43jSWVO9d9ObhfVnNuG+U3CWGs/AgN+dimro8+dwCPYPR//0UbLzzG
7MYIg/yXoI3H55yY65vI1wIkWVy2+vwoDAYinOp+LxbXVK5Buizi6413NlozOAOs
S9ueSr43B9SEfIBPglitN2I/47fFBU3dLPOJKzNvcjwXj0PCyetj5CCQpOu9crv+
1SC3Syev5rzZIeV8bbJe6FPSlLmPt6JqvMeimGi4j3CK33osXNmCYfs8j34rzPI0
Ooe2P1HtOIZTIH+51slkgVzhvWnleLV/Y/qX/BFD+9jJxzv2Gk0oRDAru53i+ENL
FG83U5WGwdV1Hlj9oEgluBTd4D5sNe9p4UzlQMMuxMlEodCkMCSI/QktQSC97BRh
v/B7um3ExKuTeinxtGwKZa+/g8/xlQXVuZTu4U8FrI3ZX63g1wgqdLoa1JFMIE+U
FfkHRBrSuwcu/at/N4xRM/XfdUGjIiZK3PzN2Dmq3vmpka0RvLAZjnG3XLhahsnK
B66j/2N+/NsccD7sbxolPd3TQflDYAXy8PV51/1WzVgz/S6uJ9DwOoFg+hVzNx5I
gBV3IdFszBNRCLHu+KdTuvZvm2pEggF0DMX2Q2fjfPlLQw+K3Erd+ST69tg+VzDx
x0aZliNNIxUFHKRPWzJHnUgHQ36Ia3KppV2GyJZkbB0Bwe39Bk0aLF2svFwOGxZ0
ccIvH4QxcSSk/BcvAT9sBuWsq3Czec01FS7APMt6x68ozlXMudoaDaw5Sb9Qiw1C
kYPPZsJLCrZftLrgdRUwdlZKyqbBgRhqjhIjZsh+NHveQAhg4mVgMS+wDOQT/l2w
fO0CBP1gfSsTcZeDMR22OZ0gTGr+g8TnB8oTjj+cU640q8K2Uknsa23/xm21xsfs
0eUFyMBgPcMl8a8BpwEfwlxXgumsJ4XP99AN7og+YZsF9kftZVpr1aVqWr53Mdqf
s297qm7sQMdiFQ54BVNIde6z0uScfFDcgbQlg3rIPM4aBJlEYChkwGHnMIiML+Xk
koH+CvAvCB6qRI9yweoOBwbaTLr27e8Rfzb2Z8RVD6e4kt0UbJs5QOdvMWfwAZUK
uEqP7GPwT3Mb2riSZRTzqDEvtP3kzj2ALaMh9MIbNPEm0BrJuKMdES0QGsc+BrnN
sstvbFA/ZqZv4RjbZlQKxm2vhW+Z57e1TQ3VM16+jN6HrVLIN3HZCzFeFYQ2cUkr
FfEJPQE0BL4+lst2GwTx9e9F90eEk+sjvzqyJwdGQ14dFfcHX2Gx2/hbm9xSDNrC
Si5+FWoekDhbeeXax/VH6euGFC0e+4hS5T9TXqA2JH82uzo0mqM6qm4KmFtlFZIT
qXgIp3E0chKCFkrP37jdej+c3go/5N81xA+yaFB1xER27be8NUJ8pJ2UQCnmepUB
Vod1q0TTgezivFzJjsX3S/GbjJqDLOSc5zElzkaXjs/Cic26Yc6WzCKKXmHsrfRM
XC1fvq76Ncr8/PSklPoTbTdWvoEhVOIZhihUkLA8eCuiACAAhTJn/4jLV2pvkKGE
wEq7FSAyncLQWsgMZHvoeU1P6qHjp2khAk+0TovKJeHkXr8Z2OWcJlfhVic47QHV
qp4eByUsDDlToImeuw/3dk32VcCXKZNQTC6pY4a6HDS8EGKEZ+c81wVzSLWMl1E5
UXcfrG18w9yCPOsKTtOFx8zxQ8b+bcRjsPaJNtuohdqXtrFkyAD9vqy7kVuHGE6O
n0DPl4tTKgxQ1QCtZ1aQsaS5FhpsNuSeu90tFkJxAwxADKtC5SIR/5/A6araAeKb
AhbpbmfHGh3ebvkqLV1c+L5fOwumRL/tUwiztZ7b66nwbkTr8LIkYUEFYaslWWcX
fRpNSeYhY7YiI9HpQhhnS0IH8RHca90xoAyPxCBpT+Wg/w+a6GVypKWQNg2smGL3
IY7j9En8TfhY6AOPpvP/YghAvW7xTvW8FRgiS//sbCAAjig+GrjmX0fOOEfZraTO
N+DlZHQuwpbOoUR3D9RYguk50KW2hV989m2TnK1hAy9H/tNMrln/6CZiUfpxyATo
BwgBnDR5oHC0OtRG/hteX5fODSdfWa+S25ImhK957i6Fzy3VCW1MA28B3u6BkMlY
NYNoJDvypCd8M+wBJ+VTXdUinkgXyWKSvIIIAwWpfYecfQsDPlY8HIBuQmhZz0/3
KTbeOWBpaZgBpGxlLm5bY5NLXqp8stVux16+2FN+v6Nm9BJccDXxulM1Jb/ZhyuR
Uj2V7R9+eboS5p0/4frY109tOlsCLwNzxdBAPh7zAZUgpHn3yFCkutKHGbMdp/zm
Be04Slwx3QebslUIhbfHO/A+2W6rnKMmkAXuDs0f9rOkzItQuHqnJLoSY7BsOMvN
KGd6LW60JxrPhiAoavsn+FAt4lLhUFtX/GmGPAk6g/fPXSaMrgJFqnvnuykgoRzb
FI9BD28PPg8gV8izFgtVBr1pZxQA/RuIgJy+kNg4mFY1KSnKBQmBmsuce5uhHBjh
75cXBtXTCeky946QdVY/5bprjB3lbAQ/Il//CiSlNOfDTLfcASBDUCNYXPPrGqDG
gTzNelbEm+s6dEe+ziHuznFxLU6uBO5mFAI+lXbab69mln3o2Z8rMWEYgLsmU9T6
89nRe2vroC/gRNQ9dL1reCtKELh8RYm8bUgJ5PNZqvHKBL6QmDhqFNIusL5MZzfb
ldC3962NdDezv359Q+yGLefweBEleEbo4JcI1IoshyausMMjUImyiop4RT9b+Jbt
kZK1kESuQXmHL8ei1M59YGPyRdWsMckiZFoPIPUQDMLuEYLiBag+kOaHJHllMifL
BLs3FoBIJFSg/UmZ60giA2YXo++hf0XCgS2TS6kDGPNHLncFx6EQ2MD21ElFX90m
SgkzM5djOFH+yrhnwqKPNQ238wcNa8hSySn113ABJG4HoaaeDEBjwWjJeZzt4PFw
UT2izkzXShCc9p72jjHREXh63k+j3ZqiEQc7nra5qANM8IGFajGOxsZasqolnFNa
/kl81ySq4nM04xx24HMVK8Ag2rDklKhSrlxyG82F9NA6yiVG6vVzCu/8hnxKR//5
jGJJf2x+GePqCdVwB5gZrvPRFgco796QRBLcle7oLE3xaLbWbM+HJaCucqmj3kIr
q+FCAZQZRv6mfLCnNRbU0AzvCV0uz02qKrEQv1T0DR4AXYKrMna1Y7Am1zNR4WLW
LFM4HLobLVGNoigOvWCPj5CyIepyVHj7uQQlOQRS/YYUG4B6zLPSCZueFWldk+xR
UDVzdfwSdaMEusOk77BaZhB4sFgl2+Zi1QT8SVRN5Wv5kjfMpbHK0qJNFySuEN9Z
4P6lLcEQv4aLQiPGrPGf9B9Ame6uc9AcmLoQd5F9t7I3Iq6TYWnxW9WYPHmgA/79
LGULQKLHW/uWqOqq8jcEgao6ZeCfSpzi9rrtxPTd8dcVObsunf3LrhvhKrSWT3du
CvfiHsOmCeGYVFvXXi1TvWFd5wdfiQjldt2fuBiGPKuHdcw3EvyJI7SeMItjKthF
ODmt0nRZFuvayvnwOy1vFumDAbBeUam/GUdTl7QcuIXueN/0M3Fuca0G2QAN8gEA
HhHHc9VHI8fcnljAMMkQHMPnYUX5EhYidrvEyBktsn+EvTNW32uGgCuoN1GB/NNv
VotthKL5KMKMCf5g0/ub5hKTVTE/POggbwwZr6F6Tyyt8DzdnH0n8Ahi8gIk4B8c
HEcxSo4ksM6cGVPgDf7VekYGiCEEeNqHSToc9B0PHClRQe4t1y0WpoC3x8e5WTFP
ElUp/uBFZN4TWqS13a3bGrPz7bR4Q/7k58u88eJMWfiiqMGadjx5+GmIsd1czgss
B0yvr3zQQlDDZR7F6tFuk919auo6oKD0QmZcvrGnhYfwh8OYFRDc/tF56Od0QuLa
5BdMaARqCcJ3ce2hiLM8CsS2oAMXfgTjehmPYLjYYql65ll47zFOkZnqlTBHvvL8
kG6dfaO5GdnXqZTG9nIgfo5FEAaVcHzSZxJxVTrlGDpMVpdDsGHXcJIQ5bFr/S17
61PIGhyHDM9vpwnR+FL7nnSC1eybHMhpZYPX6uBeM44cJELTD3ohXgEe004ltJ2u
Suz1uVQNNJrZyCcbzf6VxgcFZ0c9yo8npuX7AuM2/2Wc5KwVeatTJPEMDgZS7jPg
JpnjJSU9dR2hye8FwSzUzUnfetWQlnok6xtpGcJ4ExJiFPyz3YAMVtT7V2W39Zk+
m/XGQT+1AcBYq24BU+U1jiBzS/n+FEODSco/u2kq8BWVOlso0SToEgJ1RNS4pzEm
oIamLO1e4gI7vistvwrGD9UebJ9B6TKjvC+0HViuTjhoe+zUmmGkKfIHoA0G08Nv
yflOp4EoJVlV9ARtGg7GCiRx4sELSw3MpDgZpXOiEACUPPCZjDJC9Kn01lo/x4Mz
hjBBhmToC62UaVVkb0tPrOqA1276r6qN/3mfUxpxJ5YuoRhONHYOI+8NCyrsDyrR
R2TZwxnEUV9zq0shARkbUv1vun5/SdBzXyq+3hNQxdynphTqUhlqWfbxttKD7WG4
aR4P1kEklEHQBE7P7Eq3T+UP2flgdD+H1Vv+NmyMMe7uNHRDFoOFOnq0x0pc7Gk5
tuwsNdmmJdyenN3v2QsUccojgfQZH/iFunWkZSzaEC+G3YneEcZy8KFoaHtsEYBq
H9Vx+3Srd1RWM1aJzlNxDePA9qfR5rLrDDzWDhdMME76zDwz1TPhWezKgVxlSiQl
iZ7DvLXUcU6AtQ8t14maBkgIH3UO8YUYkP000b8r1eZavXJhykqJ23iRgAWqEHvd
/QyfbHlgd+glJy9Hxz9CZU2jDD8v5Y2/hjVECNBpWhQASKGVLt7VGc7Iu/vWoPlk
ySYBn/FuGUHP300fBSu58rpU52q8Wae0aL+JSZn7llFaAGVEb0udGrjCcxexJy8r
i3sHmVZMwHzTxghj1rnLipKF2CjTYE0l+lOoVqOzRny9uI+BxYOCa5YUNzYCv27u
C1FH9Z+KBw+Ryc6qI4NkuR/01qYLQafgWDZ8+yyn2NVDrQg6kBAeqSsiroXVbuCr
DNctFRBXY0ObrjAYH2XL5xjPQdKNM6qdKR084J+ZMNqNJhsS+ezHco3c9K1n+XZH
tt/2MScwVRBNqrDOOME6ze3VYn44MBFlPFSyas7nPyoPMzEKKiCnmS4TvppCA+M1
w9x4ga0hJEA0dBaFdsNaXy5t7pKlBcqO0IlWMyLU8RynWv5NP8xxRwynvCwg8Hcx
iAkvvomm1ffTzTCZ7XNY8QDmHzEELt90GO1MXBEigL30G6x7pxMLs/vYFq0FGbnU
vycNX0pgKhFuTpXpnnPZHlvqZkI1lE2CX8gPFBkpAooO5D9wQacb4Fn2egggY7oE
2gt1R9Tk0T1LpUqGSC4IPNO7+cFogIlpsuCd9tQFMS7V1VQQ5i4B51sQVxyLUtlm
gC8Q73WLZORk4eSemvwLdl2KZ58Ag6wRvFGh9qSJ89/h3OXlrXZiDQ0fkFR4f6nw
vPThIj+iRpZ7DsM23i2w7wEtxLW3cSsgCG+8fIYuTIP9U60yVDhqoDPOJUCFs6Je
UzSa8KbdJriPWADW0AWimVlMnuwjUwA02Gbqiu6wxrpZOx9yHxjr5fqysNztKYdX
6iTjEBzeP6Z2hsVysndW53jgykeevmdH2lEAI2hqLvRB1J+CxcOdqo+UuEsk9O0y
5Cca+GhSOyZSGzaCxrRV0iKEpApsDWHoJCX8uYCBoWlwtrXdr/fNoVY2F7yxwegV
cbXhKo8j2epi1CNQ8i/VNXXPcQ7OuVM5+v98GL0oeyE5NbfAx3Gddhok8rls3h8i
bci7BsBHq7YTmCKS8AFwJgBJzSLKSEM0N/dRxUPK2oR0Qa1OHl/JqesLhghIXHUw
QSEL6KjqraPpBWw0almMYEBPKSk8TV2GGoQolgwNJ6qydFRkyAxHLEDyr2VnBgOG
ovy5OFIYsozY+gyton1Uqx2YkIzXCx3gA8NiVRn2Iqw+j6kQXXqKSgKD5jDwKF0E
d/OIL8y6PU1AKUbtxA3v1GhOPflX87DTBSsACWo3l+TmoZNWiEK2NyiZlbcqyquo
wcGiaun/FhOfHdNPtIGnfEJzXrNARXDCgUFDX84xKiJkp4og3K8ObUNSoRSLQiP7
YT6r7VG81nttrA2qNjb9MIOkHeFtNvGtPt02XXtuqoTJ32qIuSG8sg/yn7AsKxnR
Zqc78+29fzRbxDl7pyqbdLja8NDNN55TxcBp8OgTX4A3UdQY89BpZQK4G88pLHVj
wpp0KWFgLUei2v47J6v+PByG7VZs/kObvZ/5f+i/3nEhWsEDLS2s1VAa572ZFMna
RxL2yBwUgy5XzmLIaKqNBWXy2GzwRGws75mbnYUx7m9s/L3hKnbd7AcBNtECHy+v
BA69OnkjJp5tsU9qeAkQMrt35+8SrEtsh0fdfqn0LMIdPyKkY4gps5OEn4qS7XDZ
/TlShnwrRqKJnCNddgnVYcHA6XyEMYdyqr21DMmSk/Sb6qGRJn5InRhKz/d2niYj
O4/7CpEXfooPzb4JEBOtIH2Jt95gZ//TELvegKRH+JvGSqmnkmPFK6qs2O2PILhs
jM/xRh/MBfBsObNW/YZiZ3+teijACKEx/KPfqQv8YWiqcMXD5gupQ8mx42bknN1P
wV3sB6AWid/7XeUeq6/uhG7AJVrPoxSkOT3liCcTjTlzq1Nwo0FawqZ3l/OYRVxd
nx3h3w6lxFR9DOJG1j0ks1s/0rxUg01nm1LaEOhOM0ZG4Kf8hBUgyxBut+F31T0c
w6T3owo7sIqO58ixSy8lqBvJ4i7BWpfgZgPqVPJHEgEeCgBO/LwaVkfbNdRGPxxR
U/E9Q0eOOObkuCOG/dQdsKh0wMKusCPvYng8s/XpuwBU6gPGA74by80GvblDS76W
bSNWP7Xy/xSK38scLrlNoRE6LJr6UVKRKKJms/Z5D1plCUsX183ctnSZhQZ8vKUO
uj8lf5EhAVqDhDwFhMbNMrCEywwfzt+SoH07/zP+4/4r1SROV/mGFhpKgodgC8Sa
TCW8rJl8iYzB39dxQvbwykkQC1PNGzAwZ7QNbGFJoVD8FssdumHxkgwgj5NYOJAT
O8nsK/6NIM7DjVN1cycoegnJhWBAkRJfuVmd7Ot9ce1jladsbnBo1h4JToRxjdmV
bfvb4rI+Gvz7lMTk5nuxMFls8SQol+4ZkKuxOoyt1BK3XfnonTnvF4up/PhEbIBb
q33DmCmCNs7djO/QU8uCbGRGR7ATx+QuBDxwk4ljSDZgPOCNWKkzKs0Oj11xKeX1
VKSO792svlQ5qJ7Minu+1yOnreWRebScfmXWxStxA3g/hOU4+OfQ/nuY0un+UwOA
/etESyTPC3yA878mq9D/WPMrBOHTpCXwxjpujzu1lMStt3k144Z8xTdYRczx/P/P
mY6yGkJlnUZflEtc5dThmCLSGSXtCT0ckbov3cLLhptTHJbRPrdMXA6pfSrZ+OpG
1IrZlTfjAqv2QAFDHlqX20j4ix0nsLqb0kkwrVckIsTjqtO2apylwFJjk91iC6ea
PXtBgf6Wn+3uTtNXX7uYCm1l/OR73JVuBN8IO8m78BipFktm6NqfHVKiQWBNcu9i
WDnm6Kyvr92m028G3Hi+2X2beQOJPwCLfnXPYKRcrEg/pUGAGiPYz+l6JOMYf1hs
krCXDnOeJTX2aR2pQBKfznwIv9KWj5WJdWiaX89mpT6JlSxSmFVxx6EuUaL+bkph
VGOJHt79sbaTD2iqmUR5LnQ2B3OizCVA5TrsvFF8z2Cye41j8KRoWDDxyviAlUf7
+710nwkO/8dfYodpI5e1BM9PxzZe+ufJ29u695OaOvgsMTViBXg/7PYBRadCBSaW
t5deSnM8E1lpOYs7WdARIhrbMsV4/xwgXcDYGC3srgR43SSH87zp2BRwqrzZkC+o
Y2ty+xvWZLTsQSMLWxvJ/0O2x0IJtUwugqG1GoQqDt1DqrGICgS1yG9TYJIJUd+/
WgvxOTtauVeN4Awg6PrQyuR+BAcF6SFnuS4ag72Fpf8FnGNSyGemKlmeP0G4V5H4
YRJW5tkkh23sfHpMk81bnsrWk9E6h6Ztj/+euGtDq78/Hc19xo8WR8oRKkXJdO5D
BSKrAd4o4Tp+bt+IsjddN1/HoKRxjHHcFQaEdyUXqxQR4+bd/leTw4SRJ566FtB4
T0enjUQjorAK344gEgmErlnDXNXbA1TRVtIwYCzkzbXY12QghtqxKS+exiO4E3PO
OV63Az6DgkDibGHc7L8+6DUpy7eIyCSvukdmM85gW1z0I/pSRtPuWo1SYS8Oft5G
Zvg+fxWlO/TXkUOIF5w6iuBfKS8PNzJNjsdMJ57nGtww/+mpQl28O7XiSqn3XOWg
ZNfU09B6XM6eZWqKaFqUeQQz+0CjzUjkHvfFtCEr8oQTS2oN342xp5zgeTGpXqSD
R/sY7Pf5xO/ZvknCSn0CUV3Zu0GtUDJgsdxYn1inQB3vyw1SvmaU1Wo8j02po2Kj
K7x9XQDpcOzRD39RAU4Kg45Fug+sJKzdkMPvJyVs1B2Y4zbfk0VV4cdJJ2BIWFXx
7uOFrZBN2bsQuUZ2vjjakMOAfYfktellbDgS3d0AbDLG7+9PeRp4+r8xY7zlB/Mc
POmSFYEsppwKd/nu8bYoB9ZqfRMXWD5Ox0tFK+zarhPgm253HdqQ7DMWeH9DY7yO
nYnTU9yw8uFW+9QLVxvqmbplvPXPWp2iTj86SGxwjZKmclam3qYxE2hU/XOBbqGa
Ky88uGlYOuzg3ANFD28eRqll4a42XssE7ckJPKC/SYBW8AySbxq3mlxAHaMWCNgN
sNyl0G+yaYumkssQ5VCnhCbNEh7VU+ccRJ9u3vG9h2rmGPlaIUBi178AqDnMmWfH
LfZCyNdYRP1xUO1n4owsTF/zcMJoMs5GBPL0etm2CKTci57OZdhSIqoCvZ1LHplK
6xzkktIr4JUlF7iMGbMTsKkibIRHIUNbaufx/XuR212TOgDOiJOHlA8v50JVEZ/z
nnBm1onRisezVFYlJKLyMs3/m8BTtovrNPKW9KoDoyDVs6FMkbChzyy1JrJlGMSu
YnkZhN/egoOO3l4NGCgXyy8GvMkCGuDMqjwRDQPw+4rHsjO5a4hWrIol+iL3vu2P
VKslBdaabkuCBcq2V4l8uGwUVxdtEWdGtA0hYdIN8SXupfl7q2npSn1TrJROpzrp
tbFIdnBLPnKHMYokKMwaFw7Qp+GUDqG8jCmGKlE+eJAYLU9g0Pq43xIbH5GYLYTn
ZLsSB0P7MoAu0/QzJ888NIWGRJMmdWSNkS1oFeIujdDkpFIJfRTBGMe/T8R86JI0
CREv6XSzWj/F6owUdKWod6AP4Mt6DaQnCrqKjUz3stwD3qjQ+Gp/bevU8UIXYkX0
0ibvhAcOgyCIqDJtrhizJKO7b8d57OsZv3YuMp2QlP02fHB+/pxvfr2Y4+msCybM
rdBdAA5beVvcEMiw3Y27MVZCRUI0LzVyOP4GvNroPZsHx2mlqUSeJtNa7e/tFtfO
qvJRH9zx2/yz9bVWtrUMJvL5P+aCCg3dlIK6SitxfOGyrctxeoeGZswAlHC/RlAS
j1qbWYIhqJXKcZ+oCsgV79Dx/269ZcP5dvJmkZpf+snz9PXScKZFlqceu9ZKWAUU
1mxhhiDBz9INPDbytnaxOhYo4v8v51mZOxWROIMWTVccnu5OWV473jXUk7M9dNwb
IQg03Iu7m/dh70+EgUffrfDaIA472X4oBzZTRUkUiD/Slam/R3CLIqlOY4wItup2
F5qU7pX9DrcH1pG8whsZtKSX1UiLbRpHpQLl9++NYN7hbaozT5ki/Qxm8NZnxWSB
CC/cp5cAE7wMagaVOu7l+AJ5OJ9tlaVJRGMeGaVv/ETH3/RnIDTtYwPkIiHBQjQZ
2uhfJn5bcwgmhIeU+WHl6mPjGW2nykM3GoC2dqPvJ1OjKBWiFVjsoAD5BHpCXuhD
POR4lHSk1T5GjiNl5dv5wWt5FPwM613rVAZAY5EGlv7eaajh96FX+Fq7zPTJQWis
qrfioJpW4rIXbu2NquRRNItzZwfooiotf2hkh+ugu2uz0bzYcJPXVe5grwJNhZGz
m3Kz5ELDAVarm5TqSeekCpERlan4Bp3vQMXRETo7liPshXpw/bHuUWLWMUyP7SF+
1L/m1szIXS3AQWcV332KN/qmz523COQeo3rlPtyz8liWCQI2n+0zRfLYJ+DrSpTp
GqpLQx2i6xFEpxRU4kWeWaYYSxm1qgXkqNGkMJK0HK9ky9hp3+Vyf3XnMreLf43y
s/6SlPLiBVsTpKmIxX4//JMtNfYeTFKoeUIKUATwXKM/Pv+5TNdVjWbauUL4U/9x
9rvmWkH4JMvR1jcTXk4fMgKNxyErgTNEe8n6RlOFKUdeEJ1czXvnFsEr62M94JRm
QDhEPTJBd5u7oah4O4g9SvTBHBECH+PB6o3OiSKuFfJ53iRAVLjXdQvpKDLDGD+B
kvOTUsxsik41HrhJkSARlM7698XE9q0CL1U3QtBdxqmFVsD1cUdRzLl74vhJCMuG
jH15liPwsT4kdPTuDU5k/ZbNc6rMj/C6r05lwgvKutEZAzcCBD256hWozXyspVsa
xgsTlYe+pMiKs1nbeNqjEMYiSgV3IfNIpKBCYVC1gFkyTrSactv+2jEGBmC+HWT6
83rkymfniFYGcEptSEbnq/HKmnWY7OKdWlr+x+yrqWmpb8irCN+q/mvB6QdTKl/+
+JHrbHC1c07P1mrNGaIU1MV4paQSz9MQsW6pH81AWbbEDu//MuZsssGp21ZNrUQs
NgPaxLh50QwJDYvHfa4Umq9x/rdNalIH+5NGWa95YbubUJ6rzjpmaIoMTeCmNfWR
qwAwcJJi4OnOC0nv/XLEx9sf7z9zVxzGfaHMiq3xH04UzzoOg9BiETv8WVKu87DS
9/dre3WMOJzFq4zeaPHPFnaC5AVaX3YolH1njE5+KYVCS1MulCPmXb+Hs3LCjMG/
GpVoGY527xEMIFTuId5KCarQGW6i4ckAdjy4QRvYywIKASwuiEqpXvmQREdYSueD
AngTIqdpXJhXgMzXzyO00cpB5Lmn9uUW6Od0j8gi/GGmoJc3i4dU5IljY3se0933
i85eXWIaOM4cR8OEe25+lyhylEmP+/yFQfhVNVxj9YLt76fC3pgs0kU4o3yg/86U
Zi6EUdw34uuC8kCE2uSocBtJ9VNRTClEwbxh51ni783BXyB0vnfGNh0l6HTwGzTe
czL6A2C+W+3tyy8gnxXFpH7DI/KKyps/wLgGY7KKw0n04n49vxlpvaJjrfrBVr2b
+Lca48Y/SyEktU6+cEn5B9u/vaE7NFdiiSjBkX0ro+iMjCNDW3BwW30c6OIjcYiT
kPjEVoKQR2Snr7ozKlTbdSuonLCHHR7XxjbILQCdcAG5LJsIHazryCvkgAcNi2DC
0oZEjF8ltABU1GCHwpB8HCuDlQhTCdek4+FwXRX0Ph7PCiP0YnS+/b6uCF0XN6lN
TUNJnbe2n0MUFqsBOQwSPRSYP2oe+oXlH+uglwVbRtSAJvC0xkrYy+rBuMlykkJW
frbpurFulkVBFSJY+KaKadnsncxTncBPkH4plijPXeqgBvg8ImVdJTjlLLEWlc9c
XDJlzLMwbYBBG778RaY/693NYRjaqL0m8zX/AZGdU7yOszrPHRao3WhA5l4I/7eq
E18tMh2v41E9YJ1CM3VexRr+JSzX3whH3iFZC/xIoAtMoqrK/iHTQk1RRidKtBwp
Cb/BcsC8HsZrRAy+ky4+Ej+7IMM+QBxKmD10r0WQGMCnjfJSkTYE/8vVpvXwHq1d
Xj8zuInSDgygAUMja/K+c7O07mzPA2qiLRpCl1dT1DfYMdwHK1fvh8Mc41YbBUpg
KGDxJ2QglMIftDxb/oZAa0bDBuWexyNWZhaRFC8p5Pa5wI3bOPbJPP8mVddTq9tC
EPSLOhPs92k/OMqIDzMwRB3QgZLuH8Yb0EoSLJn8D9OyWw2OQjUxB/Xl3BLgi12C
kHmTW/mbbbuk4NO81B9eo5+ol4to9X+f5VQPJLfjvURt/deKl2xOoW21gQW2jYqL
gmdp7RMGr3q2o6Pn4EX1KNqlkrUyJh/xLK6TQ+7r2h4kxQyFQlns/GIe+0hJbqcQ
GpBURr0wqBWO425TsORknZIFJpoGDauiCwDodQ4JowMLbEbx81aPlrv6OGSTQqKu
/n6aktwu0RB0m30uePk5fvmWtLWLDM58JHgJ1+lRX1NhTTvk0wHj/cDXdohLFSP8
h6xDmZGOfduB8HILXEAbGgBzbNtFsPtOR/XKQuWfwCdSo1/29AFC78vfyXPHloOj
y/OJlpzFt7xmGUY3K/3qxyYOeMaP0sEq0zu5qMcJ2o+YNs7EdDyChMgtXLlzkrg7
H57oY/vRYi7p/rFo47HbGPfyrstBU+6IJy5hazFVHJlI4cv7rfx31N8vjpGzmt5t
W2rRSZY0nnA6q9gDO1uJBIyduxhI3hCswJ7WJktQi5yjdz0u2UgHopVkc3R/LMX9
uTx3u0WNemQHwB/hiHElyHdTNRO166TtSxlrSMRlKygLJfJCFvdtL10TUbTuyQor
2g9X27LyS32pfnENNsmoxLPc+5yYLe27hcB0b+VsCW45s98nEMDxn5RfUs+Kw+qv
6056POq8NlVA4IsmhNMHHD/6mxq0UyosTLXVk1q+BVr5WHXb0W1O+m/0nvd13idV
aanG5IPqYsAVcmOrAqs2SD4iGVu/G11KNy6ohRnY8Ixmg96sLoEtbSLfA6AM/tdn
zmy3Y9rbiDpyT2L8PZYr82AWdkAP0APjxWCGRlmtjPOGeQA/ggRBthbCLED9DC4K
e4cJeJ/P8FV1/uRpjCVg9eBWigxWHahSHLvUcdgB//Cj9OYehpnPGmAzonY+lzOj
RFTGfdInSkv21zsSJ34G05EnFdYE041LWu04d1wrANhi8LlmwksnKJFtkDCk4YW5
TQdBQkw/h3Eag4Y1GtqHiec3xltdJ0zIXhZQEQGNAMMKmyVIxePwuvpMRSvVdagP
vZ2hMazTcRMvtuyCazWTgABGH14pAd1SKZ/aTEILkNi3m2r6BYVe6CxwlkjfEn3P
Pg4khfOIuShY/dwgW6/K8gR2RoED6qf7l82TUVaKYAe3gY1gyi69NkMp/uokASrA
BBsIZv5jY5CcTRRIeZMKbpmwBDfyZVIIckJhODEgAKTTaiuBZVJqfcsjVJTDTQTD
wNWgmnwZkKz/mSDmhri0GqqHUGNqgdHn+ip8eAl7ftVCG+zhV96BwqU2I1CIytJm
Sd6EPEsRKxir8so25BJNyT7Bn9OLlA0u3wOY9xojC7Fuv0Tvn5MJvltqrdAbd8Ei
j0ZViz1lE+NNUbEog2XuL6EjBDNpSjmUF3c80ktd/rWXP0R15T5UWYNoWQUM0mWz
M11IBZ9B1u9aYeGqGIJ2GVVo3zrRzsTKU/yIRL9/WkyzepL/mJcrJiG4bpuvDGU+
7/p/4nnLqHNl8rTrhI1+WSZCen/kF0/Q0y9iHRqD6WjBxSjs0hLhd6DW+8AlP441
0mUlWY8Bgdah1Aw+stb9MjJfAw55Gfi/DwSdIu+DJ6UaTTtkxFNlgKtajBSIZKkP
A0JJl7O03cfpdRDeHZ2tGhkDnZxFmSaIc71O1f2l7dMLLIc0oKVtL8vWWtNh0+fF
Vvn90Uu0Sy/mHZnt4onF5EeehRJGScDGry7J/JN62D3sraaH5yrk2kY5YhkMSLv/
TWUNEogivjZQSL1KqIBzcN/x5GS0euQYs7xpARCNwgIvm247ktfdcDUhPO43n11S
lvuo29ybbaExBTpitZq7OnNq/B9BW80ncm0ac/YXCz6ylrbAyiNb9Z9fj3srDGjI
DaMQ+M2Oad60eNTHnhYP9vvk6arXaa6zWubz95pMfO9NYrQceNE6DB1JcHxkznYj
f9dKl4pcDJUcoPx7mi9NiNwmi5xjMx7aIA0eAKEMfXIQiVWqLdL5PzXlLBd8HXnv
p5/q5pMWnDsXrsnn0f5hQpMGNyt6S2XC+gAqLpn/A4kJogCrIEvtKbV/KzCRAo8T
uSejCnUx2r3q/J572E4Ot5Bh12gplWtsbuyEf6yvEHLyBK2rRKAj788hTnvDvYNf
h/RT04N0hvYKkEZ0DuDouq3rspWngqx2H2vZfpQZ8rZa2bq0N+ESi3lZaCYCamjC
TdIhzJQ/eX74gkEFVHegBdqdJ6u5XarM55FYV1CR3YlMVUDOKS/VyrrLCMW58V+9
lw2piEAzJ28loa16iHVeihKH01/oowuClGDSGHQup6iIUXOgvWyAtmTx8SKAMC7g
U6zXEVtEj8RedrfJTlATBBHA6Wb8hfLGphJUU9NkWfxChhUNOzAEPubMmvek9pGh
qrqeNVxwl7WcJvJ9IJCRcUT3xCCa1EU4fLDD5+5xTuOPXK8Ful1NwvMVJp4oh25o
e5ByjfcOlcEYYH/u/7dumVQi4AOx3yazRGQ2+A+P9Oys2S/4HFbiRr+ZSKFbLOHL
fT3SDXVhXM0czwApmR6L5cmz8+pc7H3hzVuJb5k74LiigGUaTQ1xdyjpn7oELOTw
xuGpYOn2G+Utpmqg/a8it/QayxPHaTuWIslTAUI8r9QeClqlDk0pxdv+JGEiJXrA
vI7itBlsO/ONlGsCdC0Xki2Me5TdtjoTCw9bKB3lnSTOfQZJ/SWgQZQq/G6KTHJN
HAEscF8lJgdvz/ueiaCZsZWW2kj6l6ko0rsSGsKGH+MktjzYa3tfhaahsA1/g6h9
m4XHhqiulunbADk2rbHGWDDus4wfkXQZrrZRf1E2DqrJfjon4cFVAJqj0RQWPEsv
GGy4Os783TJ4NO5VHoJ/fyI7VyGKv34RoNAjz25WA+pD8B4xf/fpp703F8Sxt4uA
XD8aQUGPQPeEeYj/ifqNMwcoteJJ5G6ztLWyqF78eiQBxFXJv9CnOiSvjNYPx5A8
j+BUIdUH02rqaExJpY5bdTNyd+hcodi/qqci+iHjlyyA2mPYRhvIIiSFcpzKjC34
/TFwgBEoowrk8EE/Jy8Pezv4TbnGYFTd416WN2EzM4ZWQ/MGjgOuNuSYkWp2j1Wc
JYWNoK/N98xeCCCdtqvBkjUoT3E0XYK7QEh2OPaBi7ARDPTKBw5MZx/jrr7W5ltS
gLXRY4C/Jgtwis/XSbXF7eGgDIpxjB0iYwnztrwU/QDwYCgMCTcahCMJILil4pWx
o3sppphhORk36Y6ZM5gvMeWaszZPqzSDbFlg7oLRFgq6TZQ7ooX7YSU0sfS0B9mL
C0E2wiTF6cBT2wbxR4kabT74ugg8A4/b204cC4GksvURckLHGV0i9FP3ZSEtMavn
RIfXzewmiJ76x2u/N28H0pIR0+dsf77pg2ZfbwjPF9rjbReIs26Wd4wyHkf/KTF7
fUiGxid1sKmbcXwxWcL28beLh9cP4qQ217x47E86X1NDK83alx0VeCGF939jwi0Z
YlgI505AZWKdXOZm4SXQORaxIE4JVBhsjFOO71uOlmqQ2K4rcgUyu6kGwsDx1crh
DGhxShS9Fx9XGuwrI5ufSrQh7LhnHyJdgcXCH9g1FeoxYANlSMIAPXuHvOFwEaxz
TKdxIMxw6ijtzxFbeMStyUUWA2fSkj7EUOp1i05QTsUbRg7L5yZ/ZUqrBIUS+t0k
xKfEzMAmcMU2VRcgQUes/SW81LjZsK0Qp6Sn7RG+5YyoeZlEUlPcZvBhz2mjWn2C
2g1QbtKScPDL79n4tnfQtbGBxO2ZlQbOfEjApqNUARPCQuHEQi2CPMvkZRI9C+CP
OsqrPic5Ltad1mHF+tdc5KI5UjJveWz6/g7FTAI0XLWW8jEoLZN825sdFvgdOO8y
59WNHQ9ZROw0W3wjEV+w+uV8mn74VYu/eMlvcBowprUis4ls98HrmzITo7qjzcpQ
j8aEVV4Oy4e7F5YXR3EJpE5KyRgtFZuQYzNL2ThQE/IoDOq0RBJqIlCt6oaG3QtJ
1bbSgPQGoBb45QhU7NRQzfSearP2wuVMN8BJ3acEBCRHgZyUUPqCr9k5SxfHeokL
agL9kbx6hicoGplyKtjGtrUWJq5SaNkly8HL9/wpM9C1vUyzbsMSxq9JtWLJIZn7
DVrIgSh0e8sKxzc72NeuViCP1fmJq1Rlshal/CtURM8NFCZ6jDpPhqW6Ow01O1w8
IUVZ6kMXNmdBN7bzzjC3E8pA08XyE1HzDCADJ61QGG3fPvnsppuyAQU0JBoHzzPi
prIaDbtv3Xz4fE4SOz7fbU5FORTVEri2x0pkhkmF70tLWybLWfM8xfujSvvagFI5
YIN/DK60mgqiGivJH5CST2gpTKigJ3bCGpNGzgXA7SnEWbiU+4jELXSJiMk4RUkg
8ZYLRbEnlGRH574bPyEoUeClmZmaXhMhpURGrXeUZFBFU1J6yGsJFPuku39OoPcF
RJ2En5Gj5xMcROJ0tDRI8l7/lYCiAmLuldv796u00V9NmLZeaWXZzXBlUNEmuzRe
4sRQ6nXuO4VKgUxzOLsdk33Qbsd6LLtVqgZVPvZzhPCb2PbnLiiZMaKGW/nKUcVF
e3t75+1u91Zk6KKbyOei1c06s9TwY/aHSIg+sUaFfCh8/jRbG1TleXlQ/3isOLGV
19YPY1Ej5ORTWWfoSXgi6z5+mZcZlc5dtdNjUlx9rY5qjwDpKMiqksT9uAGO8tjj
BP9Gs8keB8Lo+0wCGJ3kd+DcCuKJNqp0puLTo3uWkcxe2QIoBsb3N0ICQ8+1oSuO
94vl5Lj4vVU0zb0QYH5BSJ4RTFzmTMYp1kOwEEnNo9skQFg4qO30xpkDBX2KcmFx
uTieL7jbEzYAHGcvIx4RcXtRjwl7oolVsIZzQiltG4OQw34P7sFmbaC6gU4OPhFi
lCbvRgbgk5nuNHm86bzB19DJQ13T6YPd8AoL+DO7/zRvHAPnQjgLzKnRTMi0TYRS
OcYlVhY9Bagbyjx8axO8Y8XA6I8EVRsnZ1OL6u4/DV76q4JpTHlW41sbt2qU/ZtL
yOSSuNa1OeP49slxfdRWPqWVM6HjBSNPYezbDWcf94zUMb5ja/uqezEsDTEMWi/A
utIoYf9Wxks7YMxBDVT18jC11FD0a55+GV0dHb5r5vmAq2fm+GKO921xldrPje+o
/1VIzZxN9SQa2+ytUIGRGEt5pgC0di3BOpeWNimMsFtUg5KbQ4DGu79oIFTrHIhm
pen7xwfqKQnVhty/gI8OIGn8hekBReXmAQFPJkkCNZd1V6u+y1BaqIO/SKKRx5lP
Fr4CLItq8CipnCpj48UuM22UiHPZd51EHPtZWBaqyIRNTEyuQrxR5XHOGcW+Tokr
Zpjs6fNrg7FUIKHRslHueQIy4SYWuhCxSiRzC1Ox3gc1eS1Eyi5dw7FigM7oBZ9a
kemcSELGZcoULQWwIkAwlgWXtrD8buHq9rozi95M/Uc+yCIdBTg/dVidBgs3VG73
+Qmr0zR5KbPGD43zq6E2wbPPT17i6ZCfvJQw0IbG1rMDU6jwlcMrZt1Ieoq2YRKv
wPWQ594Ir8n02zmnsmt2P59jRxCzoM+aIjsbiWUu/VmQN2XKaht+Cw25iy+Nxca1
DLETGoPJv0OZil5B1kjXzujxxjZ3NkTIvZ1ouorRllZmdgtGg4lut2AJTOj3Rg2w
64CNLheF8Mds6/sc8cRL75Lua/t0AV/iJ3FIED/+qlbr/Q6WRyzI35PSj6plLYfn
JLlieAXSvWUTS1oAAC+eTqjl5DYifpo56SdUXO73aj7m4N9OfpfNSk8xLQfMsoXP
41v12sD31fqLVoeBkyBS6c8BwW2vqTOav2g9FAXZoCaSmiBX5kWATfWNqHqAl43K
yjYNfGYEe9t2xTKGvfpHG6i5IIaesL0aNt9WJbDu0JljEX+U4DwI/5LM1ipCHzfv
DWMM7653okZuD4XlS+/NzHInHwOHwhUE0JdXXc4GLbX4nsxxBzE4WjeLFccYxCq9
d/N82bYscN4P5f7fefTJ7aQLMuI0rDNN7xA+O3Emn3g533FMFxNGC82/HBFust+K
/f0Y+25WfZuDERVMvsK/b3MLCd2FGjF7SBDtftNMyiP9224UCb1UbGgJ2SPMtgTM
a+Nx/br/2nrx7T9eyPuyv5FPcPjkiWZYnr5qgeejGNikng4ZY2PtGWB8SnksZKxf
Gfuciyw55p4ZyinVQSQWIaXp+u8pgi+d422KZaj3zvlzoD05w0lOd8neunfqSxlb
cjAqvTJu2yt82OAN4pqt3w4aF8wxzeSTkOCAGIDTvGJVWAUNqxdvRbxqp0X25lmZ
U8v+nzMTk5jkQgXMZiXjNIPI06B96x+1HXgUtpRP6jiy9BFonGz6g3ERu2W5spau
KIEiHpur5QuFd1hEtM/6/TldtvjJM05fnmwGCwaBbSKF2ljdLHRL53qEAizaCq/n
WgdZvU8tOB/b3N3AJ08rR2m7ZbCdCl+d0q8tsANSmPbK9jULkKnkaKbZGIgg5bZ+
3l0sCP6eL0wMHLqh+4peqxSVbA7qPcIRYppU69Rk3sBydLaRwp6S1mTquo1SSQSs
p/nSKgXxN0fEFbg5eZDTg50i9PZ/cXa+AOgd3l+7WWKJkdV8Xm9Au9ryq5K4CQte
6jZBtzA3ics2HNZavCznhBWHZVzwu2V0NVYzp2lyfcvi6HOEQHTGwZMR2CYRB4rY
/lu6wymr3tks8WyWgIC22hW9XDvkOW/OxJd5y4gS8wQMJpXCb9w08hCIuA921I0x
HL1qXnNI7j31qIH/aj8c5LedU2BSojqyTNZeSMZeMO359Ud1/Y1NwuNSCvjUq2am
VqFBag68/DsYnezmQHQY4KEwT29CHoDBdIVk4rUuPDOr/ALZD4y5v6ZeXZ+5XuAv
ge1Ojf8ihzGhMcj+isqo01GoKW67RZrYkiCFNULO2XC9muittmMor6yrkPoOeoTl
Qkdxi6uBlUF1uYWXZJuBMcM9UWTZthtcKM4n1s/dnwa5KC3cu6KQLV10/zl/Wg87
jShM+mjPtSu/MxYF3wiKiJw0x/Ydo2wWR+AJ6HHy3f0PMzlvdu7yIyCxK9ZwNbxA
TdKCk7hnMvHzZOTGP9Ln2Ox4loIo9dA50v9Snq9hOPBdjfBSxRxMEOQ6Bvidu6c1
HOhAZYXFv24t1X43m/Vi4xL6+4jMcAc8UTw68inzuUNKkaiJiU63Ssiej+d+fr6L
NWBCl3QagtlKKA8EevqnbyxjDEM8O/2EE+shZioyaBRN25qc1WArvCmnR8VmXkSJ
WNImAtvdaZfAeFh9EwrKk1uri9KObRMJECBg9DvXCkyzK6w1qxQlg661yHAp/AzO
DDHkFSm7csR3sB3rg7WJZDfwLVz2B3NxYrFL3TA978KYDxCq0diAy8ohB3koFktZ
hQqY9aji+PiONNb17Hm19RLNv63B/yv2UxZmFg7OyFgcfenaCpwfmeG45brdV8FI
8492oh75ZHkPGWwmZKyG+N5UST7Q2SPc3aa7qJzuKzISeCi3JQG5ao+xtvqEB1C8
VymNFG5XYc8Y2q8DZxkQlrDVYSX6c9jwLx9W8abO7UDFsnM6OWcSFpqnL0qGsnCr
W2fnPTdE/ceprJJ77EQhNz4lJQ0W1QWQaTx8NfFtXfhM86CwCPrVATJk2sTWvNUa
7euIpntTviPmwSOEV6Vu71a5w2psaPaimAG1qRACJdvmqHbLiCHVNtz5kf8l5gr5
6R7vhHly3cWU+GhYEhrMbvBQxqMD+SJgEuailp4M7B+TseOfysEKQ6FybWSAb76k
dLC5rrzkgbAMfzuu+wQq+LHnA5n17U1wP6RUNPRXoPuuFj2HyPwNQUIUL13IVcHS
QjP4xrNfsiimM7KTmrDxX4b7YH0kxa8LKPsPFFeo/rtNdGVIBCzGWbuE2Nmwup0L
8aWHiMWgyJjdBWLKWzs0C1W7n7BgN2VczyzHhBbjTm84t1vUZ779N9UceJylei65
mMy7quEmwrWglZQA6QNVua21xxcEDkQ+Gd8u2vEpP+e2BJDifFDzo2nEaSzihQEU
kCm6xylqaAYEUc4yyYbDVCyhKHNai6m+LohCIvPd8k1z9VLpXBeZieovD9aUP//J
lxyfR4CcFmex7KolQEuyQ0mBLwphWnhOUBePW8ZDPRJgEUoQIPfMoxFw0c0Mv0av
3UJVcrk/zaNv+g2X7veEKZKo5YyZqEOePiGZtilBcsDmGJ5mB+cWVCa/kJ8D0aMM
I+gOJpVJX2ZRrFUgc2D8dobdMgvO7LqK8H2F7CGg7D3DA6mT8D97WbW1LWD6tlGO
395hM9KDRxeyN0gow/sXAzOrIEBWBW/oOB9Wt/jp8sMd3TMo2/54w5c7+84SCYQN
sMgZgX2VioSQoqZwv1oDvw7R4Xkik8++WziaAE+WXv0XkeX9J043zrS8AARq4InT
iedIuLYZ4gaidYk4uYFMUfpKCy6WrjJVxGjc8kWXUXQiXuA7TuE19I0KbdwY9LIY
GffV1MNKYO6liyo+eb537IbDsxnlv7/pNprXBDKpCA2DTTWYtPEhlKVqGNGmtAae
/3x8ht6Umipgt0tff+3X0CLkhx2XyHeajuc7X2pnquH+fEAmGRgHEXSfmevoPuJd
DWbJekCu3RKaAjFx6YArvxV6F3YYEC8iUUvD7aMVSG7MQR2nuLgrITs3HUpUBU7P
2zsULhZiyhS5taQcLkEG4bXObYj0fNlqmIjPgYED49HRSjYF+euXESB25s6wGAYL
ZdGUlWMZwTJwwHmHSCsV2nM/tXQZq1neETYVJuWMqkOLbgM500cKL9ctCTcjgQV7
hyjZeha/B7BDIkzhE0HLJI7W/YLPbRaEeZRfNR2Y9M/wM5GruPCpA1sVsPpmQOos
fiFZ5WXGtjybpUElg73lfT/P3u2A9TdNHjOL/2oCow8vLqKrFCv+brOzWWIa0k1q
Z+0LqFkVd7FsDiyV9Ie2Ksmkf8Jq5yP5oVY7XBEerneMAQn5vkQnEob4SIT4Lx+p
UwNc8seaR2HzwmW3CeOEkZUQIku/Ykh8HUaj8SPgnrio3dRI9edO7dxPRB4q6Jyf
9x5JFhaIMGMprHa1BmmIsfqrPF5b760YH5WaSuU76RMjtZmHopHm1rR+1oAIFkHf
hSM5ItQeD4Whj54bF51/9BVTLHZDj6Hqs4dWcH3qpmTaNb37kj64BYk6GB9aJ3xZ
l64IAMsprNaEpKjuGZ7+wsbW4dxYD0yGnNvRhlXmj6WLJCZqjpbz+esKFkcLh3QK
s3Ec7ZkB5cDLh8mhk+rL09sz9SRsg17N2l3Lw21v/uIJYj9Xg+mkK+Q/S3+HUgly
ajNlFENPMbc/3mEt0UIoZ/JpueAiCWNBMR4NzV0YF6PyQ+WuUGtNgdWSQF8+nhY8
ezJg2/qwf+9Kx3stTnFJz7tbstHXqRXVAhAM70vELlwlLlPMJwzBLGUQfOsg2CQK
9FoPpE8CB3634pzAIAEdPM+dlT3NX+kALnEPAToH6s+PPODNzTYcAvdDsscaK1YC
imowik8Qwkhe4Te8gWZYoNufr++9LQsKuljRKLqqGTaaqTGIMpghCoQ+roa+RrBy
zSzIe4LxVHL35XVRpY91M/xf000o5DLVxWRRyCroPGjlkq3hUCE3rvFwOM7BFWOp
/5t7mZVtb3KY5APeLMLLz1PKI+5Td99JGpmGdZUkcuS/A4gPl8nBDV4Ny6KEoPJw
nuTFgT7un80xbNgSZKnsIoaqITAbjangqTI6zynoonFj+F4igvto1OPY/kD5+k6G
woPZtrW6rjHLMid6SiPA50XqoX84ESkmrtGAD7RGzw1hanjvaV8+5zLhIyEWB58x
te16fFFaay9Cr+opvsKGQYZEXLIl9qKpdotJ2cU5irqWsEsaNdhFsRklC83QeSaP
8j2+s0FLdyeWP5KaptOBQGz/4NPud1LsWZ/6nOQuwhFAbde/ohw/wzGVyYBSzeHA
0XptcZ7PL9TJqAttRpz1MLpP1E4dcaYajbdtjp9VQfhj6sztmgQYWoYfWmA9j79j
NoaZ5L6HvJPiKGnK9H0THcxfm8fr9bObPDRIzT/HIz5qClNKthx3QGpCwo4zQVXu
0ycQ+RywmoXvSASICHdN+54Wgo4xPRUdsaQCjq//9OMyS94wdrhSlTwfh963b8fQ
w3ZQ3keLh/Ue1NATeWqaWvghwIT7EVvhwx6XrViWTa85DHL05+z6pGy/EtQwOLR4
LTuawGXyqmARDG7spwZBPNCfnUP/dXee1JatKv8FbfBcXwLn8znS9Y/WLUVsPbCH
JRWvsk4tneISeKH80wj/3TcYO28GuvRMxUC3JlW3as30Z+Ag99l66s7lsNMYagMr
KO23GjYhXoITgF4CbxKdYHhiYTXIiCEiia/CD5zl4YQN0Vr98OU9Df7rJWt0rqHw
q+6tZIHdMPonY1gcUzXjAO7+QbHJT34rpxt6nIiOHNMQe26OhjhhqVgdGKqpE3pb
JMXroFz5satO4dxAJW9gXlzuCxuNA7yKbOEYtoCfFnNTFz6bOG1BCJzi1B+7cx8M
CdquauMEBdvMK96o/0ICxwqkvQrqgkN14DYemx7BOtPq1SHpOR2/70Qa7Xt0bYk9
76dmpznXmjZUS6jJgWUNgV9YPHz6Jv6kxXTzq8UJ6oJZ+KO7nyK4V4m5gpcPhG1T
DBIo7IYdVJmP/96AeEUJT4TRbLowWaQ01it0r+VqPx92irY+6oGsdeZTvasRwcrP
H+fAzksk5bvVWk8UARjbPtzq0EBBNeDB3DxWcOnZwGm5PhZpCDLTcCmxmJxILp5M
KmTt/7yyHhtOoqQpmEsGI//pAENU+cI+K4RVyKP+l/oK1OQvNTEhpH181deSGQdg
BsmkkXgrnjmCzqvcIyu+e3AwYeqyC/tDzmNCuS6lrqWZeqtnflhVRrIlmjxUWWf5
AXFF2mR+7bPfiesBgbG6zX7CD0yKlvKQDAvF0YXctNOSQLjChBJvMAbl9IUZSeYy
SqD0AEYqhnHe37k/Y4xuDclFLeDLf3GIeVVUIYcvF86D4F+weF38x9WamCnizoUg
KVn6ERgFQdlM/dHNlzr63F5rGiNOa1S1nKr6iL2TsYsWJySvgWijGNG25rQhuZcv
thtEXQMRnn3krMwvkgHF3MFVtc21MWNcTONsxLOAIqLpPpjcHwQUxewE8yZGhpBo
D8eEkkKmUh7hwSerlTFKXgpyOwLejk+U8eSLvHrIIQXQr7x01PnMUqfTMQBiSZvn
kkkxu9mSTqQYh1E0vpWe8bMX/Qucr8M5H+9bLyFrByRWTbx79yTH+ibY6dWgdwnC
EFOGUt6QeMeNRMH1x4gn8z6LLCtiVEcs4iE+WIaJA+LANxVLYXgHZ6O6Jj5fzRWC
yw3AXNIEBbNVs3L5lcBbaKqEFd7aIYkHzSeh9kQXwqbnMaxYlnPrCb68Kq1f4Oud
ANfmoAJQDxGKzsf5Qynziq7qM/dOTCQUFrMbBrGFRGLrdbXEurOeyuzY1iUTkjL4
eKtEAc3mM76v5rs7AqwTvPkvus1bteicfmZzZZwsjM9SoNPTUD44zLBXt5Z64rLI
xY4PmS3ewzPYt3J5KnCjWj+bwWaSV0QnVnXfAsMUNoKm36aJDbdNH1ODmhmGXaA0
KNtXuPjyjriu1h6Fyp0f2oyNOvQ5DCsE/kfdK3rKHwfR98cczV+Z1o4ogg1bXOQO
QCKEcXxxmNfNfeYiKRsby/5t4Zrj/G9k1RV5KFcjSsUpS3KCqZ3Hdp7JlrdkXsMN
Gffz3tYgVZBwKFl4uZgBFwl+K2fWDGsx30/LBD+JzGtgm5kw8DIlPmSw7Ys/Z3At
Cv666xScndftrCPuAm0Jww00or81b2d/3IrnAjDTvuNqoxDOrFyfkJk7hn0j07Hb
TLbYMyK/0cW5gFEGV4dHYLVJoIjqsIJaElcvr8uN5qzCClsZP4PflLwUELCyyV9T
nulGPjIiNVBSwtCL0/0Hh5DAFSC+HRkeURXYsiydWLlaR5F/GtbWM/KW548Xr3m2
DraMzo9Wmj4EoQs3B5HJiddecIsZXZDiO5i2p8iMXNfYCxumogDw7keIsMbqz2KP
cUyckOPEg9HG7z9fnKJmGfJeL09zLdigF2Zuy40+R6KEX/msY+hkoZae5Ud4iVyB
JuX7zoYY5Ruee+gAwqlGSuRX1dnrvR2inibIK7FAtTm/08AJEccsg9DmeiA1preS
GlqA30v69rdInUv9LQbkQgeUmuXB3B2cffurKgfUU6jT6H5txPiH5Hr1RzWGyXf8
Gr6uB8nXkfYpMeGoVxM5xN0kTA6zCn9Kow1xu7/1X58NXLmx8wI4Xy4qnI1fXR68
PMzT0bEaVWYjrPEWlC4BQDVCsgixKPAMOtjMuVQrSpF4mbOrv/sm6rn+iDNaFpx4
4RNrQenI8vBL3pT2ZGBob2Ow3dHuhF2hS+HnH9ChrvgplIqB5K/xUXDaEvpjEOOC
J+7Jn3cumNGp+nWpbysepm7Wgd5BRJZTh213ikRp/uXnfu+niOGbWViGq7OuIM1O
dFMbT/FxvKOfu5QtVhcUYHCW7aTHzohSr3Yz5V9/fGPD/spRWAnbZiA9ynTVsNPF
yPyoylbUqsZ/QHrzDZpc9MtKF9+mCiN7PNwmoRBWYIC1qflNT5H13qeh2JKhqFX2
kwBrUfmrUz4DMwHY3mbmNJCtNv/Fg9GG36ZzUm7GcksYdbaylENhpQYwPib4M/dE
ezyx9LRlLZuamj/DlAy49TKU+kKRzoJNd+65/WvrqVWMTRQLp7Nu7ChAJbDEqn2I
VDL6aArf/8uwJ//e74wkCrKwxGu+ZVXIDMRD8H6JT2S9c85IRLyXg90ul8+uNieX
XZ9n7HanKD4I4cRFp9oPoUD4nSrrpEZHZCQ8MkY+q1EpgzsL0sd/bLt/VwWrKuvB
vWYKRQOPR7YuFaN2iZUpmrOIamLuLYMCpgvv8oj8PnDltPth0G7PESe2aXNY5erI
qJL8aMF9FRRxiT8Ig/1aqMK4ulERzHSj6ixV8/1doq0fE4mHaWZsgxvcB76Jsx1U
kgI+JLKQSw7J2yo4a1CJRwgOzJmvkPzImJWcOyraHHsW8rHYMEuknkQ6Ao2BVSpU
p7DF0SbKfMSs2abTAF9eJWty1VHRsfz0sww+bRmwu2BvezR20bUFeuHpwZagPP9i
NDtkX3tdkTwql5SY5VHIo01zilh1MR3gkvSbKddrarueXlLeLGy6gD80fLi1WSvT
DrJA/Omp78jjNgK/+ldB+JRMMgheznB4I//ck/yYhMOF9CskM26SPnF7olBOwgMn
iQHm/AHksmW5S5/kZl5xaNrByJ1l/yrsV8pMyhidZaZMQ6G96SWKu+D8xFUCk1mp
1G+lDxsc2eYpfetnfNHEYTvoBq09+tCOEGY3U84LFt66yAI3ggVj9Ixuzehx+YVy
q4GSq3/9+6xYcqsDXwWWmxjGAMV8C3QxZxZA/Ha9rNy4/aoMW74H144Qbk/V3qma
jzatMWnrIfsIFXE3KKsrl1ooM/Ft3S7n0CzCAqkTl5oArPTSZ2kzK5khv1CBFyRC
PidqV5KIKMDB61ZB218BnFUSuYYNq3kEKC9Y9JFgF/CW1hDj4YRVt2d3YYALrBoO
WxggS/ERaM3LsgjAaOXTM7ftoWeA0b4ATu4Tg5M0J3X2WhfA0pSnucHuzlaMlw7I
7g9/BIy4iOXfS3qFAbIZso7rKWiWD3zEYC2LwfxAhh718PdVxE8MOwpfClAbW00E
XoW/Ga27KFJBCi+2SrI6jX/sG2YixrrycJ/VmmoGIp8NbOhNHkQnSejqV03rREta
yfCJ9FCQYgt5ZWKbHSaF67slG8AcjoUoaHZ88pGqEx76u5dE+Kfign00r23g37+t
Lrk0NTClSazIWYxc3jaIas6xH2QA1Fh7RMEAzqgMTAODMz3SDP941S3TImr10B9p
0+BLjmeA+TUjg/GJeJKAP5VAGwRNDIKOnJDU9VIjrcPLwcerhv5u+2eXxCD22BPg
21n6B+uUXyA2TQuuTyyAbFcdpHPQ1OJ2BBrthsZusD2k1UKSB+Lpp9bj949vrvB6
K9qp2PjwAyx373QpqZX6Gx17JGJRe67NbNHimymPVlgKN1FD3wi+Cq92Lfqji1E7
JE5DiwXZrueyjImMxTZ7QVc+xAQb6td/rHWn19STDgZLRgUndsHCeqb7JyPdUo7q
UzTC5xWuKFHkNaQ1gSoab271/5pd3w5i3VGf0r8WETD+Z5S5Uq85pROZ9Dvzow9A
lhKI63nQG37zGOW1c2x6qj3zF50GOLyK4/2nsCjb+Py6CfxgdWyb9Y0L66MNC0s4
4aJerjbJY/Y+gPCco+9GwiFL9UqD+JFDWS3WX473wkZi+xrLSf+BoGT6Y7Avw4Vr
HAri41ks/sMctF9AZS77OYnSN2s86JkAI6U557bMeFdavLvoylxVgXWXC4MzuVtl
9pWyrQEkYnLRNUuxL41ksYqxwsPkKfo7H+pX6HpSGzKP2ghb3vZb/KeKDvcwv1iB
rDtvQXhbSAB46bVIpicGgUJ5qem/VcIwAFoSpey/Zumr86PIAKUZOXCk/Zq7vgep
L5/6E7Egsua3E5lpyOCv7U9LoQm7bFDtdU1bsm/UzSWxTWjMJCW+PE+KcMdWnneN
jVcWBwFMZ+yPRop+4o8yzOAoewsZQM6KO7stYIre3uexAW/N/p2rcNodQkKivZou
x7cz3QMguI4Z+VgT3+iW1A9SufNObe7c/UIVI2VxOw5El8Y6epB1Ga4ZLuUH60ub
wvbwuextlY5g1ytsdOHBmJPwpBCqYk8kPQrdGTIsubzKEq/gimnnGE8ns7g2VCJU
7s1INDJApYm4Qfhk0TFnABfuXNDq6b/CWYiQI2bW9tAqT85BxYLsKCDgkxXeC9L8
5ld9jrm0r+ww4xaqxzMObC+ovwmFVnQqBSSpFn1h4ggER8xfo7Me4NEfUMqrGN0o
aDdREbok89ydz7nvDfBQ+sVg9WSVzxNMW+urhlfZE0EJetPD2ZkjVSSFiO2d/G2S
rzlpjYfwBthuwk99mzSZohkZFla/qBsr1ZwZdUIM715t8Sg55+QjlZtGle1ahO4j
OgWtn1ESL+cR9wyOzKMUh8wCJVRivSlzW0KJPDp31Kv9rniKkTYm5Z5q1B9W2qMJ
iMVvxV9ZzFSCvDZWaKb1tRjJGPrKNIWQ3BeVQ9cr5ATUB4y/9aqGJL8kZ/vWclpl
jIN7bG6hev6wyBClvVF9d7yiOYqt1xZOK9M5Hata2zyrBZkxW6I7ehOhs7zAqdtE
29e5yHXJn6y/ib2e0adhZ+cDSljm4rOFPYJswWyNc2k4JYSAyi6ixMMMwAN5m0hp
wS1E+oAFKoyay+SlE5OM2VRYTNqxTK1rkZEpLBi9mCxwpsXjgNsnfCdv6tWxOt/L
O1H5hs0oIKxLf0xNAluDgw==

`pragma protect end_protected
