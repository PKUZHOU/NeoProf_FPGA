// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
AfTKyMlD6Uq4KaEq3VXbch6x/PFWEQ9l3RDXvYJGSiEPsSkCW8B5Sc9qcFy+2s5z
3ufxCY3nvF+lSK5wIq97RkAHMNkx+elIahNS5ToautsKga9NVyQm43pVbtd+9NiQ
qK6hxqP5twwB2W/3NCUqhHFCWiFzVGnTXYsQAaMqxKE=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 8496 )
`pragma protect data_block
oWVhz3d7mvWdAagxT710qdttgdZHiKMy/70Jr+G3nRttNzho+j84zu4+TG69Co0q
EDNWH1gFALiH4WDkz8lToY5U5uMAMFaJx9NcvLkxHmXh88k3j6Il+9zrlY7Bw8SS
GVAXgIFfj0iZvq6zWYimqzGIy8YZyflXb9E3JDtPXHLpD9ADOCFD5pEZkVVRHzLP
osl7E1NAR227OgsYjDzeAYZJGvkNGSsy7w1Xyxqimsg2n4xerBIte6/pG9NhkoCP
4fNNJ9VJAKMB4zEKhUQIt88SlzjXiiOvcOLzq455vR2xrG5qdL3RWoW0yJ2Mk8To
flwMXe8Y4JWv1gwmsRG9oYypBAo1JgBV7sGjxTs9nauxUcrB9FZ4+0TMd712Bxdz
1tHu8EuOalYb27GsvlysHATl4Ydlrj1UKzsXgIGpl3zKJloolNIKgM6hkl50XUIR
7bblN8j3QRdwUtB9N4RZkvHINSc1Fa3v1yLNkdFSKs9BeWhS+vJnP7mjANjVrcVe
TU289/CUZ6t2DdR9eZ3XGKii0nKtuLwwVIRgFM/f81D8Lj4bfoUurfS/VlJVK3os
zRz8FHnlhoKUiS26lE/L9P7Fvs4SRXFQULFwGSQktP0lOxdmLnk9fYSZ3HzwjRy3
CbCipwYqlpoInJWSXoL2exv/Gf/VDZwGHvdMHlUYPG6tAnM3JssaVXBxyX+kS5BC
CgIVUwL80+eS8cuDkRWI+yIAOMDmliB1KESTb3sx1ZPwV5wsnpM7DkrWb4FExj4G
m9XhZI3OQTwgFR/PiB2or9Hosg5XtMyqealwZNiUAnORXZXGmgVoRPIu+2gWbmk3
lxLJDg9kSeCsXrGVPsAuIF1PBQe6KSJihNTPf1+heZKt7dMKXqcX7bfFowLWQU0O
eQ67Y2ug3aUQ/weBVvlxtYP0Om6Es/XVjNoz24ignaqKu2tzjZHjtljhy/L/Qqqc
KvfBPUdzzpTl/ItJQosxi5b4hb/4Fpl2j4CI9mt5GDU3LvPMzdf8l4kJ2F9Gp9lo
1To4S21QjdgIzPKa2uA9/yqILsApbie7rcal2z0HjzCOX+V8tkzmSJdY9DixlXrY
j6c6S0r6bJuJjQc0Tds38ghjpmbTqCnGKttjzwARni/uYW3R687dCp0yCE3/vaWw
6ueSY2pqmtOa8RokeVwh2grmSAyzQTNX0YcipIn6DYqZ9Rb3yB0BclS4EGEYt6GM
tNJp0XVR/i3bCIhexjLH8U/WPOAcPWJXgNzOajv9zpoboNOBjOFq0/Nnna7+sNnL
JS4p9AkzYgpQruvxvgfeJhMg8Fv1N9EZwUUbYQCmDqhFvSZqi+kzNG5cG1QXT9lO
Sqq5OndlDEvGA+IL8xP+6kfSBCX+Hzi2fTQbyou4RLVxyopr4b01uDCvkEUKPyfA
5HiO0BL4RugQSPwfsQho/LLgKvIHvRwKa32QaAmw0Xbl291f6EoCEdEM442Qk+fA
1EENx/pT5wos9cvC8H0ci4Ckp+FXWlUG6L17h3J5YdgLZKl6BsZjgf+1MYIGjQ0M
52zJ6F0srxuVCKhj0g5fbyerm9ttcN1HdIJpfagqwoqHVXkI36SVvpokicQn5EIH
z1XSBtoFP1vdEV0ohZbOM8H8zF2Aee7/eSiWAP5l8UxSuUXqZrW9BhKrsr3xV87n
ireKw8FWNiUEwtQL1IYTVC19Q6HKkzYFWMdYJRm2Y5oltcsPZSfoZ1bn8UtFPGNE
/5jJ3lGO0BXLpXtrGrexXdRpX06AJOqnHF2bmpvedyyufVNYjv+aJDR/X3PZrohO
XQZ74toFBS/ziyED8DfeuQS322v+ojsfaNS8RPVN8hg8N7zowTb1inVNaEohhY/B
hielGFV6/dDa/eeC8Os8YUM5i5rxtDpnLCBLkz+kM3A38dy2MBAZ1lb4f9Aeluky
iiA8Rpttbh1jmFJsSMXL8j4GHUjwwzUraEtKOoQpIOGx02qu+VwcQS1YEmAR3/7e
e08S8vuhpt32qaLir9YeD66lU9bJ31igjtw11Qr2mKD2GyAi8IaZLT13KC0S5xup
1vHdjWpr2eChKSaa8Zu8J7KSuU+wzMhwW9QotuaTsrOUESV/5wFPqFBeUxJDOx/w
TCvjHQlDVOmfswqzXWWQ3HutxfQ6vKGTOdtS4gcg3xGWgD7zhCWL5xfgDMonQbIp
RCCkeszXFqG/MiSSzpBzBnhcEBImqRh+mtL2tyEHpA/pLZ5jQls6xbT/tgYAJ01A
sRsGpS/Skgcnu4s5+M/VG4ljy7nrxYgertCgLCCRFS5DQG0jHJZrMbfCiSDRXYK0
74QA16Mr3nO+8XLd2ZtzseaGhzCQFO+vG6vdZFJRfKhTeszegt52yXztZd6svTQZ
gjVuLpm4Dfi7+yRivKZKZWSjqFDJ/WZDPmqaqQtUMeiWhWFMXwnKHL5qllRbcvaf
XTSIqAhT89MKGUEC17Xwu9h1GipD0ZqOpGSL0DyNSSywkjsR6am2MKwk5etHlayJ
JvI5lLazUZ/Vouvry1YUCzpebSTrQ/iAElhkUynAKpU5NCsowHce4SO8QNXM05rQ
u645/LwAQcYHdmAEZORk8uVO5y0fWSylwUc2baFMHBt4bBbeubonDEKwfr8RDks9
edfWquuD3PtAqYHPTvIfC5RKrhPhj+NunOeuGm2Ko8Xv3zOGsD/36PWbyOP2Odwq
Vk15ZvCDsT7lK8JI+44o7yLn9MjDe7n1+WUcSK4YuxnFRvO/RUP15d2LlJDQF3jV
iRtFYlbYLWP6PAlkjExMi7Najw9moQvwQ3zEn8mlm/0a27qdgRnrqEfYZmSwVscF
MvPepZ2SCj0U6TSkBOqXltU/JM1kWd3vQ7Iu3S09Kd+ni/xspzOslL3VEYC9V/6U
d89zJ8LUvKoYg2g+9RsmVhFDjQ15c5+KtmaDHJBOwdy/3NaeDNcohakvT/Fxv/Z8
bcRklpUNLLcksZSlIIYmExqjlFFifA1riOqz5mznmPiTgEYzYPako/EDOctdCAAX
na9GwZrhdA59AJf6KpqecIReuVt5qUpmzLTWyKUvydkc7B4PfqJb97i+OOiMSpEc
kZ9/B0BVPbiBZ/18v55fYDqjlSB45VpDzLxMzeZJei613dMyePfK8DvKlSjsFkR7
kULFJDUem72Ix1H/KoCirEKDF0CjCzqLUMMmIOHEFtt5xaL5R8iV6ZNuppb4Tego
8HJEn2+gb722+zOWC2cr57O/Qz/NjtgW1BS29lsqjdfhP/ufxlxJL5K3CRsBrKYE
F6ywdmut6sO/UuMsNzsc5q5cyNi7R5+dDN598EUZF7pejNQRZTf7TRM2AlE7yotL
D+jdZlY+53+Z0u31eIn8RNaVVGrvNa9BWoll6PaGp2LoPosmbVDDNSy/hRLgkFMA
wHX6huRz/PWmAePN92lJ5OFZDr8iguATBwWZY/OlpkMYwLqY7ve0HQQHzgpCtORY
rYUQG4hFMutel0OuZZkXPplj7i7vHiEMqvbuCsYA/W2sEoQE1uIh7nXFrPR8tWU+
VRueNhNiC8PYBuvc5iA8WVc5B77GNGTQxoocD94wt8eh+uRz1tzC89fK1XYqd7zn
oSlZCGevZLlnuPJuAGUXXAejrPBiE3kADM8ggJLv/DbhgEMmxf1ti980gTy2mAxp
IpAgYLaB0nPES7jD9odTTV7MSufoZ7jwSlDNLSYuGOqgTNzNjJG3K43QFGCaB4nw
7EseDUtPnRxyZ1+8awJDzHoWjX5RsEC1xtguzXJzrAVbX4Lta2c8kFzfQTOW+8q8
eY2ZXLEXgVLNxW/76nVsM5/N1mipioynNlAevKpsQL5oiAbuepToYuOxIUWt4ubW
p1w4M4iSKNJX/EZt1LreMnfjqRdl2oIHg3vAOhLoCdhWERvu1Zj4HKxuLDdw+M+3
Ez/bansFviuqzFWf6jmtr/eL4+kt1jTf45G0OGwnMk9vKZlU41snU5vy3+g5AqQj
gjPilIb7Mmd3GKbu5ez4DKW35QtpSKTc1yvY45pDk30ud5P+KPsiSiahl4dAWj6n
aV6JAJp2Al3Owx9qz56dlZ7h+Jl1i7gYNGuAnuFnxb3UYP5QInnrHc0bYz16fQNn
Nz7QmIAvHUzjAttsuCvJMhDCeY2XEEJml7KVpIczSAekxZhG6YDT+CxhqBrfFNQp
eRKto2jm3CSeZmSS8yTQ+HefsS3MwOU9rwFZjkuguQsa5ywXyA8nTf8XqkebYvqR
ZuDR2QrnwllqCaI8Yn2B3caL8uQxmpTYU642wuwF3RVz5jolSX+xgGUShxCtZH8K
vAWhPGAh1sy8Spx/xaabiFadDXYOAslpHCb8NP+qWVLKAtsAaKn4+YYiw2HY74zV
XZWYygLOlLGuLAD79ORLWz0y5ekUbQdS9Vh/bAhoq8rpA5U62RMy+3GVZYnnzhaV
SmcZ1W9R5QJlUhD3gq2qQORoTgSOowzWmUCET1r1EDGclfyjn/Z4f0q1OWUG0fcp
Ba9vz/PlApSIrvlcnhx6OXBkIpM4cbnxpE5y2MBau1KHOY6X0frCTaD3kxdL2lKr
mqIEn45Wpfh0ORw8C8LkXQ/Sgb88gQv/+9gf9mWjX2BG5Ez7w8ZSyM93cQ1vgeUZ
yIgmOF+InfLIcNZ618M2oEwYAaIuoOlgzm+Fxs1jbyt3AwkJMAoBpahZ0qKrfIX/
4ZPEGcEKWM0Do15kyxHPKNd8uVKT0u9iSmfgeR80NpA5RjiXytepJwi6TEcdcznN
SkPmt+oOeLPRxumurNpcaKy8IBUaO7h7JWrJfqCngp37W4SWXCfa4kkybomKKjEz
tI/h9taS9p43jmFWK8LqxBFwhvUJEW+qLeFqK2LDj4yBJyudXtpdKu8UywU3JD5B
ns36x24TuBG0wNBhfL3ZxdSP9a5qPZv0xR7A3WYmdWkWHRp12PzieGxgr4Mh6GG1
U4rE/uuOjti7gS/SbNH/qsf5fU+6ow51JWYuxVRF7ZSLhiQb0G5aL51MWe18mxBd
WkvjWuzLpR0G1Rycrh8StQrwWRAl83YqKfz3ogKmAfIh2AHcfTN6xaGUvav2dbT2
IYU44ofrsO8mzqVqbtSSmaKKw96PCi7T167BUccbYYQ46XV7IlhLA5rLM0lQO8Vd
yaIBdTgvVjuqOYbrxm/2lII/M2gDOz6XZ4JVmYECscGMG2oz53nOQROvkQv3y5Fx
udH8T/pM148gbfqx52z9mh4pH2IyG/QipLMhMHt0bihMuNXt/9WrCPjvuL/98oyV
dLfNfoOdRT3rjDN201e1s+39ekEI31sG/HIJm3lOflhY3SEu3vbXpY2hdjJZCz18
qzpvlgtztvVt+bg9ApA+3Fjw5bPYb83krQDuoUZ9ckc3qua0Tnx6pVCBCnJjyA5x
frt243jOIyOvKK0vxHPuDuFpwUnXCHFzOiht2iOerbxuXyhpjCydLtOvwXV2QvAB
DmwQ/AG6hIphharf7Fa4OTlVcMyHwz0ooc76Ccj9Mcimsf2c/O0Zm+9doxg4MEUq
7UxVgSMx5NE9akKhoLogBdbfrsEEGQL9XqdxWKKBK8tVmhu3jRSZEPHeopDBxJo2
mieIkdqSo8V9QCCUk8TrzoWnazDhXny+/oSGa5Six+rrxfKQuQbjg0tUnoW75LjQ
ShoSz9aikXVBEj0f5ELeEB4mb++EveM4PgT/wJPPK5oUs+YezLOm4PwOiYE/IrTh
37UDjjYKLr54VBMU86DT5pQgs/U8MTeTKuH5Ae0m5J9xjs70ST8G4HrkT9H4QCQi
JBECDTSk9vWDXwb9h9Vp7W9tZ7f1K7Z8/YoxY/wXe4BdOFeheR3cmS+7Ojxu1J53
w8QvJXnz6R5Z829vyo25cvesAfCjbEQgWtNUekcVYYxyVC8MdSV8wF99U/bhTb/I
Ecm94vK3VbP253PubmavgxG0ERdS6V4doZozND5Vi6c7Fh79crg2YXnZK0DoYP3S
q6alI4bBGV7L0+Yt6rXvSQfN5h2pupv2lq5Gw7+hHJKV1SyT9b2+gb32dor/JKPY
U5cHpWmUu9gQKCZLTmlrsKIt6Mc812cSUZApQvQmJthk70zoK8v3JQz+/Pp380Me
D2aVGFGagkAbm1DGr84vvMRVtq8kVfN9PJxVeY19TCrp4Z7Ojdus2nVvkhM0aNJT
yGE4N/BS2cOaXFajdEf9TBgSr322ztGigH794ewpQjQwoCl4snwovjoIcGdoa/sr
E6WPfaAbCa7tT3ypPAXxdZNFKIjlLQCB9HrtH8WsOrkgUlO5en3C7YXP3NG1d8+h
qOHBJijaT0x6MLOW9h/ijzps+ag5Q7O0+KZLCOyb7xkbkGonljf/1r0hlZNy/zGA
C17rHeLsVgsivZD4kUpjFU0bZPCXx4xHPrlYA+/MpgSsCpGt9Lg8Tko3/B42B4HG
GUzwm1x02cmxIcYbBwcXuIbgRLjnEWJEZPAghEUmKhuymWChd7d2tSQRd0IAHE4m
vOE9BJ3b4fxa0bgKcF/nNQPgtbsYM3FRrjL87/FQtDP9+EmS2bIHIXF7/BPsgC/T
XmKPT2pn/2fphSW6AjLku3Z2cW4VT0e4pjnPqh9Gulhz5RzDgr8qI14eOmgwRCfg
RU2ZBgEWW/rLCd7UHZFS4maQg9sbA8/pIeEP3bQ13isja/YWrbkamf/8mnsAYx5J
MlHhL3WNF+wpeX81Iqb3cqWp+kVRipFUueGp0x5872CxxFCVOIbg2fVySQMh5BBh
ovOxed2PZrd1QR6Et92W3WgpFhcwQx/Gw3fuHtyt6VVgRiK/fyoZDOcOW5DW/TBg
LLkJ0m9d1N9tJdgyWVCAJWX59KMzOyvgQXFYOMu04EUdso75ExLYy7Gzj/KWGOAO
3lPDLdywifngb2M/bC0/BG/ODi9NI/l91payv9O9YansmughWIL2pr7jJkojPYYq
cnarrGrSWMkodKA2DZUFBJW0SPL258mrt0aGxEvpdoXKRJEMmUXkQk1TJIyE0gBR
mI6QUBylbekX49w+AOWuRUnM4CP/rs7omdxkp46QAVY4kAQozr0K7M1OW6OVN+zr
nP9DFoC5LcOyToFj/5lUxYok29TvOPKK2tn8xVRGVw3cped2lfq95d5ZFv6u5auB
GSvrfNyAwK2uibZe0Zig0lCbf85AA3WhGdLxT/Vh1wvETQGJBNJ+eoye163BDvyA
IqkSmAa87ThoZCOLHIz3akuaWOLvC5bc91PBRIv/I+TzJRM47poNhI3R9ru6PxCC
lhs8R/j9c62q7iOwaUl/cYrWV+f5hCxawYGTppi4Z10WIaPtEw+kTSJlUTcrbeH1
SWSiz370QC3KLp4vrwQLt6mxtZRMKEf8bv/6vswr8usjBjmjGXDNrrdrODEHOgpj
mPTeUG1oXfAEqv0fJydXFhceaHKQHUfUWd4R2NwnCt4HDuu2JmBYH6XC3qbRTLtv
vfZjr6UA9Ry688Jswn7vMp42dS2kFv2D9Zzdai4+sfFJ7NpDlW2pswIUH6k+gNUO
xFEBoWGVBWqj5R/fFPrDo9J2DFhapIWRinDdGjxoIAF8eDBKEjkdPE3kWxV0Li1u
BtY8+p5zqucrSBUutRikm2U2dlm1QHj8GqvphBJ9911mzy1AxzPCklUXR5uIjdbw
ZpwnL6+LGFohIA7/TAypRf0TeD1wQIcFBavanO79YKuptbSqEWUpUKOK0QlVeX2a
u77g4h5iEgAnen/dkHK8hNsufVDc09q3kjuYFBC92jkgmN33zZaJ1IY5XXwta0B7
/mXjaPVV44HKzHWl5zZK3fLey/5riJKkBCDTglaww/9azQiLKjnISjBQpfV/lfLt
6AQCbZ8rHtuEjMEGLGAhPJ1E0rgBdV1fdl/oAKmyiHi2KcmGL9FfkiEootKhGAYF
EgQJFHLWIjjokFpTYsshhhThXbuW3O0J6/T/hUu9BZ6ohL/+yLHji2XT2Ix/k/1h
acYdn2u4DmTM4zegAkxlQZiHoQ6cMStZCRF+AtRv8Be8xdCqdZKR6WujIpYseJXy
Ezpf1fk1+HaOljLX57B8beqxsAXfbUoOvFo73uCWKNc1ydmWtASKtPTbSxuilqde
2HLSGMuz+y6YzJV1LHrMYnPlYIyrsc7MauqLeWKSrFowcPoKigP88DEcYIsck53D
eWP8HeJZuGI3emyi2ETniS9FWoUCAeetGQ2nVg6uEPuaXJ/rqDYsc/nwFPJshHQw
OrWgvxnn6/qBeKSrvoZbSLfusZJwbDZTuEW0RuZuIoXVTJD/XwpRipwV1r44ZWS8
DiCFmxS5Se8+5jXjpBce+vveEH0RtvOE/m+DLo5ulcfZnWyBfCxKFWmyIZt5hd/s
OPcdCUC+mIFSxHUclSv+huaDi0CFsVcIZouvOqit286aWLr5lf3y0vv/6Tc9W38c
wR4uIJNLx5EdJuRFnEBzeHNHWQftTSFqhfZ12XESnFKfySDclPVqpy+I8Je9tXsG
J52UqxOADy+1OC+AJ65pBdP+xPHI0/uhrOWshdG4A2KTtTprSsJlxJ6wAG4/NEgF
OwS7tHRLfh+qn5LV9Y+8xoHB4qhIBoLp7AZWa/wtr43oF3WKHcV2LdYrnV8IiAhO
15mbMizCSpMIKBga9TcOAxKvji46y/iYEoveKnOrsswuW48VigaFxJLpGM9aID3k
lUHx6MipqF5hs0e4ML+QyBQIoFzXc8w6J80S37iMZcyBX5VkslV7Rz9VDSsedoIi
EkIDvXeLcMKiKljVCzrOgCFpGoeOrF3N29Nei/85SqVWfFoG+yo0Os0hSwa0VUrR
OauLVh5TyK/nZTYaqIkAUdXBQoq+1gFkeTCa3EwbKyDGpROiYBOWInkhpK0y61vu
yC/f5+PsDlmejdFsMwlQwdG6nzZiBBLqQLTeOItuDquKI47ODG7IfOlQ2RfTm7DD
nBw+RG+weo47LtZevC9fG7O2qH0UvTDdyMnv8e+fjBU7CwLU12zmWbvO7E9ZpjED
7h9WXDCeCeEsQpusFGw13CSpgseRHjvXZ3KJAQVJle+YnCkMgjwacje4rIXfAx3K
h5CTylXMhNJ7BfQJRW4HDTf3gxoiZ2oC5uCaMweiGxJNPBtVTO0kHUKqwMv/xJ3H
NYUPwwYZaE2xtwSTadtbnZpF5uvJ64EpiGMITgcBqP2OqeDxY1eRcnOrAN0qidf6
IP/VdcedwP9W1/k36BHHuYtbAJCBie+5vl/06WFW2mY9gusp2IH+BG2dCN4Xa/t1
Owf9DUosooBkJG/VWNZOxEBno8vPYNDG24QFTOGVJQZML9nG5oz3oGuixYL+ubIe
syBqk/9S57Za21GH7gruPlpQV1Qy+dzaEk/kVBK5YblbmmQMX5+EqOfX8W52t/3J
XqZDJM41pPbFw5VXWhteYV4PrP5uM65vwN2+dYPw646O/2SQMUuvSwxllxbjH6n6
0n/SY0jDp600C9kq6seIv8YMMn3JrgKWNq59qnRQFqpY0g85KD9Pbh755DxKobfl
rltPnJRK5iuGoPdnWLkudSseW5CQwFIz8mCgVqc4bfL3FiNRc0b4WWuKrSTAs2H1
B/YZ7RfbSsd2qkRvoqBaxf+6rmFx7pIniRjVeqWJuUySQx3+c7rWWWD6AKUlnziX
6zOVdR4EHCppGLss1FgZ8OLA2WVPxaG1j2O8XHoIKwhAEuDbi8ZBh6YP9T7wFQXP
NZfYts/zxkfsD9QcrzD3PYmvqatwrUiMD5ZXLgy+L/sDscalm7/hmS8f8SJ+jIZb
Y5zW7futNnb1QbBCbgg1mxa5MVNkUWiP/vVwAtTg/4ywGE9jQlmkwPVBmgRQxJBp
zhdCGbfRYP/5G+xxuf20eQyVdSPX0lMaddi7CSm6zoQGaDX8lc0/Txx74eoOWz8/
Z6DPFNen9pjBLKCxgjbdBBYTvxetZbL0wCYreK3EHbURQxPyDzYE5v/FIxnzGYtw
mM4DD6KgKnPB2078mDuVTfVDxzqJuXiKtKniE42ixZAmfjy/y1hCDjvbBOJERE9m
PvRdVQ7X3Sk2UhMht0YV7HxZQJ8tZDPJ0UZoNFWKfPS6GhR2hkQKTmYIR+Tv4WNU
JxidYyh+0QvKpoAoBCpu6aHQKwzRDWv9mOR4kxtlnhN0XgTY2eceaTbghtip3myp
ZM/EjFdBTxTgxkaMlV4lM3YGWa35BxKLWi0PvCild60V+2KKowyObmDdRL8OcQyx
6tEpE7sJuBK918QbOu97RTwJiBHv0rQc7QJIOr6iHAykDIItF4K/ZuQ5/1mYE5KC
+EzDurxZZRNBoG+2nb3CkqAslKnO3qs8ADOj1IfaeuvU4SI4frS9fy1JY163BzvF
BtmcCl+I0bqvKlOW9iiNjhTATSI6SZBgupJPOM2ogIIknjK8Qxk+vDQYhViAtt74
rBcAtF2pP6dPyQOseOeo0aJWKRxwwigjEoF4YI/qVkfb3ijsi1SXp12YifLNjzAG
kO8NjFovv04GipwE9q63avoD75O6VIzYMgjjBQf0fBx+G4SoIj3WGrKuagPCHDPT
2/q1qdU71bdYmRpcVstiblTdG0V9nK/GeAd18ZzACz85XcItRWGLeCYslsO6v821
BGNvKqOvbioT52qceX/0O4ozicVP7mKNQEOqk+2oFJUMLkGC8APcmDdwBXxWIEBt
tadD/oIrGa+wUgk7DiZK9UytV0NcQ1DwUkAWEgzCalT5dFzFvix9SSgSPuMWN/aP
SsZd+NCht2r5hul2mfVBIykH4GuIpB0RKfy7C7rE/n7rvI25ZjKG6d3r+tkrcekd
w8U/fZqRRqfAVZxVtnSpsqX8PnNGGFYxFlbq5juewPUFGrRa0QhHyeNpOkA8poOV
5pKuo6aVVeG1UJ+VIi9o+/vu6NljHx4T3C/tpV8pTPIR8MkukU22ga/Mjef/7oAe
umM9dfkXuGpZ3pIWmkQK9oKdOfAYFRmj/ZulCZ0Zdc0Hggx2xlUHCo7LlZuLJOrl
Tjq2bf+ultLlk/iXEKg9o2fuqnGZvfy6OIN0JZGAfB+qJjPiE1kdM0zVqqMuvKpu
OUjwBAAOFLASspXvpT8oV53+HHXPzd98ryp65YzJB0SN3fmKscqrOqaEXEO6J858
xyi3CRCEyg6zY7PzSXj2Lf5vNiHOpZ98IM+E0Zso/VmIuw+708FKHUeV56POZoXx
iJOvC3Yi9QtG0hqsdWtE+icn8LQMXkA3eVOi42tRPWcYP+odGyVqK1nXIt72JrGf
uMWSoDZqtxwGYBL9aWlNlEeAnlKKjOg8jbQtBt5TEZ+zwp/RgnSe3ei902PRb7gO
gNnK3IbhLZI1uKUrEdxfVsf2CosVMdNqOliZB4pdHp/dVsXltv4cJydEwDL9E4Vj

`pragma protect end_protected
