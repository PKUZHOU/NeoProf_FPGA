// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
io4dcHVPc9Ug4cEEJblSXTVRUk4olGYQDa1XQjXwSFz0EbHNpF3CMneUjTvUIFkf
JAixSYDCFp87Ccseu90Up77rLVsW4LZgAfhBheUUecNRcX13Qr3Ft6cQKI6dn1cY
1691LFbkgaLG72Ebw3h9+oYQ+ULM6SoTSBpDHmm61R0=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 8768 )
`pragma protect data_block
hD1S3e1OygrdMYrjnHpK/3/K3WxTrHsf6/BcuZOjX7dZjlx/ZAJhH+0ZWSwtyVmf
SiIFPDkV5kwQ/mDfKfRZpXMswpwSRF5nvPB6uJ4BmQbX+kF++R/UTJYDcPCaDE09
GYZaG+l7y8WIOS8g8d/xhHNLYvGsdM2g6P5IrXIlNri+QdMrva3UrBDVQ2ZPPyyV
bIEBbyXN+tc2mlm/WjhBy+LdGY171RbmKwMBixxOiDtxh3yZQguB/tyaXXeuY1St
LyIHEhW1dfOZCMlEz4UmoTqTz3TB9owII3+nvT1WFyC3AKrD7mc6uHXJe49nc5jM
H71ANkwe1fvrs51VgmRYK8GO6/XP9QfPy4Al6TL3Sg4yWqJ1q3mJt5GmddccT/2s
6jfSMcTvPJieFQ0UtZfLj0m0mXDYYb+ig+4MULbXlJin4zQUKx8a4gCUvrsEY4mG
eK3OMkmxx9LwilfX6GT5J1QnmdwIZkdctqBG2MZYZh1Fj34QHfzcAWqf1WcknSmY
8Cwj8wuOs0e/+IlBQMsn9dvJxySYkwYOxWGGEBUaa4kvBrocA8o13idBSF3q0i1Y
dVfdYwbFgUtOOVWb7gouNGwQ8NpJuL9KciVkK2pt7bAU66UGTpHqFhNG4yq/mPy2
ve4Tdkr/uWOlZ4idM5OxSc1oUWpcbxYyaDGV2d0XPwfsfIIpKM5KXaa5BfiEVC72
vkFcC0QkDW/1HRLrkR7OA16oEumCs9N1XwDHJ4it82qmpcnwwScAbzkPGeZAR3Ds
sZ3ucGvzZaBQoNEELhhpSiaJVZ7uWn7IKJmAvUSdo7K4XQAYpVXiROYGtsEFXurv
HROQDHcOIvdgGBvjvW0hXyVKICoIw8uizYT/9lnItSvVwbx0QP9MqRwTcyyRkSbF
/INYlIP7GY2Wdvlg7eJIS6EE1VChO5IkZQIBTpvGxSBOqq9fHUBVwHI05SJ4gr6s
yw6bzipQkH5wieUQLTrueMEdXehJRo4LR5rHDOSRy5L7lqAX1nfQhU9BNzmRAdXo
p/3rGzbaV1illmgjZxvPeA873K2v//rlQhiCsGhGoMkRK402mo1Fos5SfW7I5OpM
USH+6dXseULF8wImL3e/f7nRjGyqkmiqXxQDpoYGlAwkTm3RuP8lUxpiSErA1B0F
9LAJ3PYv146+auruI5/El/mXQD2OktOrGV5emqkQQmSul42JBP5gZY4I9jaUBGnx
mLPXIbOvSKV1LdHpnhnwZB63WwrBdHQ4VKtaMLDTTXlqKetG7YvyZCZyLWNW/zZr
HMMgAAutcWxGccNyo5a7fDVrms4m5JUrGtq2u4E80IOLW70IktumPqw496mfzBw2
xcC785kf2Fv5Q73IJnVf2orYT/sTjCm2afSwTUn713X1iqxxyKujh2HhtKbYTzHg
U+2u3mm2cfDzuArRs9NGnNAIZMBi3oqH75uP8QuVfB5/4sL9UX8vArzi3800rBlO
luxnn6fYKhBkUn1tsVPkRxc5RlD666HUQ8iAOusqnJF0RZ/JNRVlPS18pzYZLzwt
6Li5kJgaik2hcsVVAsKxGhF6TDJHp7fsPc9xh9XaKUDtIFjYk9/3jUP0sfrmZIb5
lxQY3nIsR8DElK4m2Oxw4fM0yJZc0INjo1PGNLF52dsp0XNmmfz5HiZSSLUStWSv
x45FnwkfraNuAZ0VQcsqjk4WrdA/IhBKdgw8fMG2Y8fcgVBIWqxbzqv4oL3IynCA
9QJ6j2qhHzUxUFSpLBCLh2pwYWSF4VCfQ28cFPrOaXHBtyfYCeRKiLw8XazZ7CKV
F0FnonV0n19qDpyWjhnjFNx17gQ1+y9XbnqIIJ/mpDPgMKYN4OfMaiNV4dTXs3WM
WELRjndNX4hajZI90cJ/FplE+uqr+YvRrGMG9SGH3YTTL8vbecsycJo9PY2QhaJj
SwRrDkICYyNTLIFEtEdPpiW9Bg1nhYThSNkxtVhR1tGqHJQseUnXJMrbETIQzV3F
1i76h3OniTzL6hpMIa5BgDAUeXmstw0Jqv7lOGk1iQvq83SucTdK9kLsQ97YObdJ
AYmqVaZ2eJFOWA6O8gKsRM9kiD3KGqIfqVgDaDePnq0anB0KuL3kH5UO6VALiSe6
Uw0QW6UDZOMQWMk+D2M+rC/n4TTRzXwDS6Z2yaoQR4wMxjoq2+m6UgnQV17dV1D5
TsSJdUVbSQVSYbX3ES2SGWESK5pqLonXIkSHQkYk7drC///Zt7M+i7LkHT+J+m3X
GqtnlYmhiyutfDJ55SHRWmgB6obYhEbMGU0XqgoeRBXgv5VTcL9t6OWftaBsnxvq
UdUyiSnz1vJVQPBM+9UHcaD9kZVeqv5GfyOAWYFAVa0FdYTfvd5Y9Ez54MIsseBF
pVPSyqWSVzc3kuhBdk3WmUjtdlAVZ2yOkmmZh4ewqdbvj2E+U2yy552T2wmY1gbl
vxHYlsiRtDgRMmjUCw9WNUwqjZT12KOat60lVXVyyde8EgVr+kwnyoKUFkdb3II/
3ETnmK6k5nIXN9Z03tl4YZwpke99zlGyndpHyO7NfkB4V8/N6apakVrHW9+up/z3
3pDcOr9dmpq0+dQqfwytJn9uloWnljJoNBC/z5TpKZHrZqkWfvTBCAeBkX99vgo4
dAtKm4rXuSNhrFX+2glK3Ed6bsX/f0XUQTJEpQza33cS5+QLO8FwqrId43BvJkw5
aIY+3mdndb4PJZq3FTf+VYk0kOvGhrswhdxHt2C27U+5vHUIn1r/cofFOlPbj0dR
SeBKX51y7aiWL70gpFY7UejZt6haRLhnzn9FAeddjJt68f1JUjVnGerMChpuOJWy
EPe6YZduAXy5/8wi1n7DErjluE0uegLTXPGEouveHrginXurTpTl418Bpa1TGjlY
YAPJjNFQBhn7dI7WZlOWDbDEA2vpcnWqao2dkDS7BI9PwF+KpmuBUumiytOwtWW4
XGxl38v7XK624bCs2/CFb2ZYCUgNYggnYdZMsG7L7zl/WwBjo3rsX7sjY3QnmPpg
j/AtoC5zXGK2idSewCf6tTxPYyzKACBMPNj05N4rZiVIV97zyzqysb+9NtFcgXG+
/+2T3a0VKWw/EjbnwuVGAxG961R1YaASeg9k7PUB7rr9cjUxUlsnSaX/HkErqEVH
SVgPed/MfnfoxcUqJCkKqk3uKrTtBTSDXfj3HT79Ea0r+dVyOo/lf2KCilhtOOT9
fWI3YHcYVHxR4f1zc7tznoMLxsxkNSihjLntEQHDa2g0lelecRIxymY1M1LttQlJ
YfJnBOwznFl5KkoIpI7xmbqkEiMHTfOQLyppyNkhejgulM6d2yvkBrxynuvYxK9g
/SDW2JSyYplZMVTgo2sTCvQwZBV0qBTJfKpjWSzsX53grB5THDiaqC2Me1QYEipT
ML9iFEsdk2hagKssaZOiajUQYkPmFS68hwPESQDFDjZIbPjGo8+y/vaD4NU6jlmJ
Bl3bLpHXuFfpGVz23SqdCYIkyMLzq9AnN9tp3fquQOlhOgls3YhB5JYmoHh9q3p9
glT9fWxLAG3Lhu3VlcBWCjgNu1s2tYK+OwnUYn0xfM9GhTR1GInCoFyBbzuSH+4e
e0OIsllJCMftGEIvA3ZUEmi+toG9m3u5KBQ41N6pWraca6evXMRJGU1nsSJGgoO8
k03IhlpnBd/R+ALfWwJ4zlI+g0axGi6SWt31NLgTaFetAjbQcmhRZYajlpTFcYDr
xWqD4zmEc93uLAP5dx6CMz3vkZ17O2OL1e1LiHtUYhaVYAQMtWh+fCTaQS6tg0uU
u19rY86Hdzr1onc3sOapvzDyw1XLw+IvO0zYovxgBW/dddgsWDJKvLmAi/AQGDEE
cI/SZyl4YnIF4v+uOOimFsEixLFht91GLAh//bMgSHx3L7M6h2rZtjMiI/9/yAgF
qyS6U+tFilRlolr+Mn4OhtANbQyfuCfEf0mAeRLNpXsW9XAzUKqyWth9sPhl16RB
ekm9BZF5Q00Oek8ab/B1gDT322mBE5ZhJWDQn0jp35iKC77A61Bf+st1d13TK4FG
I+KgrmQj8B+JbZTA3xGS8N6Quvqgq8SRkx3jfR2Im2rwxfbs1ZKPHXiAXZct52Q+
GRFs2nxSsgnRehVpb99XvuxKlDp3qm8/81kLgQXzaduo3t8b3MjsGPhImyv9/fRT
NvHfFn2ar1Pp3bMbvf5Qi0clO4ttBdKk/ELbUaSvLh2e98UM+XXvvlubv6838Wie
nV1/XRnlde5wkv/uRbunYtcFn3DYi73jVXVu2T0lsUdepKkYsiNEtFzIrNbuacEN
lfY9gzwL0mp3Zp99VqkM0QSlCyoTNZMKLMg7zYKJyBeTz5XJCDPAI5G/fADk8DQ+
78r70Fe8JCZi90SqFpft1Ae8XVB7TVK9HQrZx88wuR2gw5Lyz28KdQTjlNbvk2AO
dLsDivJH08Dt4KtuoPzVj7RZt5XV6HiQ7LhyFpyQk+mGSbfYHjrs7iL9TnmbGkyr
SoXixoVe4fYjeyMABqt7hA9LeCMtMEKTBO+9/1vK+oERN1TPTcbg8dW8+z3Gx+hd
0O9EkCv2cnTxfNiwl89MccTvjvC2Gx7v4aytwopYvUReA/TdPZ/lA8KRRzutTiDD
sMnhJz8owXTFk9UM0/3dE6w7LpyVoXydHdiyXHC/dy+D/HgQuTpIn7PicWK3O83e
zI7N/bII04KNiGRArFMdMeK0/EZWYb7LDcIzP6yCJw+J9oc0bw//JAaidzssFE7s
FAkCOY110LNX/4HWSAnqxMo/e45zQedDp0qFaKh9lePMhnNzZhUspF5pm3hJOdj3
egOcGAlNZeGRmwaamKKkAmOBrIFOp3qFMvFXvtRnNl9s6Ji85fheQzinOhdoOgYs
2B1neD0pmtGTDiy2hXRZ+mnZI6gZRSgcfgj9H6Mv4dc+hYAk8roDXdPw+xZ5wsX4
p8jX4vu0vFrmCsJHXaOsePKJ7WedflVLvuylYN0sXMSbyjGfMFnRiO3T0Y0GOQHn
jpL9fTj8gW7bC9qSsF+bBA+po4t6Izm+x1WjqBdL39XzKyQG6VW4+ilhCcjtDc/M
dWQIknF1mfT4Xmb6PAvYehbKWG+9P+c5eIiU1KWkcJWBFS5k/20wTkPnVnzjlac/
hKyyTV5sJZwRhWpPmeYMIsQttvXHx+8ixBpWTqJCobCr64ZIyctcaWgOtdoIsHjS
BK68xhODLkBf0xQB8dui0waVLX8tuVP78xE32Y5kNZ3gdz9eUpgdTwO2vUlAPqqt
X39KOXE9ciz4bPSeuCJn8S03AJO+ef3MpVbN4UsbEdTZPdqovCQyRoWfm5uzV6Oc
VhqkflwdP0Erdt2tZntxdLck2FPK2AC55d3fmdkA9LSbRnfQOk7DA9Ng6bvv0NxW
si5EDAsq0J+7H7ZFK+9UymTbWdN+iCaG3ZttPrBLuL03L2JcOSFsQHZIsDA5BeJ3
6CloP+p5B2Tn4rUC23toBrQ51xpb5dUGWP67UjVmiwlqNuH+Cn8Lrap/zj+p1yZD
qnbExqsKhg99xoEWBxJRoyN/bG0aVL98+3+mN4gLMdU0HLLZfPYI64m2D+TJ7Pi9
m9LjVqaFThnsLeUtPRHRmDw0jdn1zVB9a0gbCKOvqVFpsejSSvflorobJQuOAndP
JQ1WzmxJ6yO3BS4p3VIJvgYlCBQtKuZbwTMWn4gT3QiSr6Ak6gfJSefDAIl0rhF8
WQI+jnH623FMQhRu0a3F604d316xFe1pEW7eFNcVZ+Vcfo+exfUEpvB55PuZJQ5T
BrcyPDNFusuFhQpSfQek6zRRtPpn+MiWMAum9oALt/l0y2oUzt4KR1Ni2uoxfvv1
H65cdnrHuZD7b7vMU2KNEjrPkdnmc2sbYPwK2ujGuMbaG71unNHq+eDSB9lYhJDS
MQn7JRbRa48uz6RtGz1wUgCZU9nn5Ma4sSzKLDLZRwYNfsGkLKN172OLihBeze0c
+9pst/chjyVAnBPY5Uyb8TL9NJ2I25Ryt1krxk2TIzL9sginvE7ihBAi0TH6ZLxu
9GCRVHK7a13+0Y6s3cAXzfy/qFKSxqQBpxJpzb3+M5D5gErAQYEn3cwbmOL4mulB
ugzVUtVeJ9S+kQKxJ8DDRKGDfkwfSCCAfXCLEntWJxh2ftUuSv50FGHrEV1RBGIf
j06J1zCNS4aUCICSzSQsfMA3xaFwrpJqUhbB9JmbhNCpEmHSX1DM7nljOpdvs8LJ
V0lY2/060Z56+J71oGEJjz7ZewCz2201qCozhCd1EVUuAakC+7xtesNWDivtzEqi
qntqZvWu/gIiqJlAbNAln73xRY+SwTjNxAd+cFEmD8gaJfObkqXptZe75q2nzcu+
BCsAfLya1/EfzOgbW9uiPDw8+CyUhQmV9K1q6jLfClJvkIW/0Vc9zdvTIbDuTT6F
UT34MYDuaZg96bjGou8GhZuWxiiaAuHSA4BUfCoTGdmPxdBWbP5mMKO1MkBX11yG
r7EaOwel0wToTZWwmOIKXsCExMRqk1ty+90YVo8QS7rX1Perz8pO0No4ZZP8xwX7
GvY0rpFp5WP1flyNgkbFKideeMUiXl13ZoRS1MbskL5nkbtXf02jqoPhShecUs4O
Eq04j5PNK/LRAEtKFjwGbb6o1nw8p7S1n+GBqaM6CJBRvtv763El+QacdvPjoWnA
xRNloAM7v70xIYu10hV518o1Y0RmZqsMON7bwKxgeYmBfRSJnXymXd9xWSMkEPsa
IkyjujTctgQOlQslQ9sU7hEii7hG1ahdBPOGmIlZu9cHuTLiHMZDvmfKpNJ1cB/I
43qQVL2nWflzGzZ/L0Rx+OQ2cAwKvWtJzJtoCfKssXfEJ1gc7y3Aa0I503pLmw7S
nTjy7uo4xLZXbKm1bgsqtMCKMuRzlgC3ZQwh9Czv7QPqTnfwGArxFKK9jAt4P8ej
V57zc07vxNgcHcfpL8CO4TSSkpTvSJFc3NlTPEv5o2S5pmOhu+Z9+VX028PwULrz
fFhbSJqpmWgnFm6dQwG1d8rbOI/ZY/FWQMvctbs4n1z5PXg4ipzsdNWToBt5kQCL
lmXxiS3TFymSyzEr3Nta3Rk3L4Rj8xzJngHnQyU0VdLefaA7k7wbm1WvFDLUkvHv
8l7O21iPjdcok+IzP9iMjO3MX4xTFCFIYbWP//EK1r+5eMhhdVOsLTIOkORzkqkO
Qkr5k73QUEFUMpyM7N0gXAPBCSnrSsy5xc380yUb0xd2UWJAiLTMpd0MDwo8Y841
bAuXBUtF0rK0Nh84j2x6imWTSbE7XQTxsiOAl13TdbWR6il4fQBdBoVI3XIhhDc/
KD/ePSbga1ABk1vTRYLibYow0nOUcpP7ELnQbOG4IzWmUURg3Ht1G91r+XzRoQfh
W6gP/cIVAxqYSGBdTOEEI/q4Y1PJKe45TUpjtYksy4zPLBM0i99lXEcbKIPK6Z+g
lITCEXqlasQtW3IBfLCY5gsrIacxIiOgQ9eVVXifaFtSf1oLYP5yRcAKU2oB/UwQ
Khc6dza/zqYq5mTcp161klVKmyXBIys0HfTgLSpaWm/o85Wl4+h6K9gR1ColO1y4
JrGemnaYDJPYOn+llFOb5IuC3B47ab+ph7YFv0KLXvn5WLSUU+Anoe/kjCz7kzR8
SnN02hYwbSzhgNsPfhephsjnRq2WJ7V9PA4VOuEjo9nN0eNMkfLNazOAdvSHebvN
68H2lOxIfQwnHYdOThTAzU127JMzHBoU3xfJ3IU9zpCX61jt2PSOXtObAhzUIANu
b/IdbTgiXGT21lHKEadU/zhqTtwjI29Yv3zeG+ckTFaM8aT7Gn6OLgyRPvhLtz+9
em6zBLrDQRC7Tu4Hjv1XVVqE+QNnBu8E/6X+Ldbcqas/M4alk5ix3mOv7688AEfp
lMxOJMk5/is8kBUrGWUvh7g02oEtq4qEdkmzhkpRdTLmjOtyBuNoINz+TMKMuwD3
42MbkK9JXsP0U/XqUT11sxPDsskENM+Iy0KYz1VzAa+h+LLxMwpbiCo5Dt+EqpDD
nA+AULrWNEEg3zVpKeAxlpcVxKKQV/17JOstPrCKYqhuI76ibxGAeqAn2W6mPPyi
+CE1SgteC4UH09NT8Rtc9D4aMjnI8lEWAQ284VWysVu9wzItapPyVLB/JyRoac9D
EU/WMvDyUqCU9DaaAMNcTi1aOFNk6uGvQBuzJ6H8uvvBEjFz3MDQwjaytpSbL16K
27sF+RW7aE+SsyjH/L+nK31bHhD+V19QxnGoWGRO7TW7+y/V5ScM5Ei1BNkVBkjD
pSPS1rijPhVqFk+MY4ghDHPXD8KB7hm7nhy6Nx8o7lChmj10brw/Mj6zBJ8631yN
MrUpWEyjAj0FlEcy60mK6uzzWH4H2/kyN+GoTI79N3cZ8k+2wJiLO443NNCmaz9t
naYIFi9kPcRLgOEP8HU/z+g+aKVZ6bXieKezxYrQZoaVlHek1g9A8LJT89bXm4iA
2QTVMxIsR+xe1y0nfcETAEuw7PvpcrJrdEQGn6MnTOeFYZRYPkbMf0IOks2hy+Nd
TrDh0Mhj5lgozGfCtdLNzGD5qS9tBAtUguUAphP1mMOAHZRClBFDJaA4WrqEnVXI
YNZ2jcyLPQgIbo95dU/IOd2rcArY43a9EpVNI7SyQkO/5mMriXz7N2mYXjhvLlFf
azCtKJtxilzNUz0d0DE6rcDyFSHQ048W4U+BMJCT5FToeaM7S0U8EEEps7FE+b2Z
+dXdzmBp7EygByWrUwfy/g043C18G8CCrZdwDrmI9k/TTYRoYoh1N63M/RKVVVBz
6PMFHlAwVNFuWr5Hr/4XBSCPtm6kZLtkWmUDM+SBQK96FkS8jEVUr9XXt9YDUQC5
0NaWuNzhLmD/HWFq0/Me68rwBHNt7O3hXfn1KguSfZgUi1iQK9w9W53jKkrB/4Wg
jcksxnN4q2t68l9/XC3C8F+5u8bsCos3CpX3aHZIR1aKSTydYTqNqOS47j8OX3zH
cnXKuoEgGLE52YEO57JsEkYNrXJ/zqu1pXJK22ACzriwHMv1t3phvyix9UJUEmXH
1grTrKg4JPiZ3t7tmBJgNpubcV1tO33J5AKC+Cs6Ed/GPF4kUX0NWWvDARhl/O2i
PScQxIMCw+wSMEQs0kcZn2RpvZrC5fQXOHeyuxgGv/7zU/6uXcu+flNiZjsxMMWQ
+KoOnZysdW7QuX/3GCy+belcs8+lCcy8IStkpZlfvlaQMwQv1C+GPDRYI1oxzTfb
zMnAMu6GfKewLHgB2tN2IxfkepkrLBiw2/t4RRYXMk4g4sfEMMkGiBOhkiR7nDTA
dHH9TDQV67VSwNOIgCZq22mzz5wurB/BctAfsBIAw1/SRjzsqCxUq+HqhYQ/FrQ7
uHdhJOp83hYGvoT6w848y4aOVxqzoXO3556nIYTDq/Py+hf7pDrf0HinbqLNR0+f
hC3DXfqSHNcm/SZEBev17OGj90yMhauVFIkkjZgXN8hYgyy72dRhPzAazJegwgm3
nOXJtMRuu/IxRLJa8yu3ixCWMCWjc0EpEMC1QQ9Wm7tYMyWh0XuNvUxj+7HGWY+b
NtbVNf2cV65TTTQy1YFp+delGPpP+G+XlwBeq3CrWTq3uXTF6kp1UA42X4Zw4pSi
I3DKQh9nSaA+BYuBuSrmQA2AOLQhStRd0rf03pBxtnOH0xoeCyOHf93fcmq2VK+h
hYjfI/fXOycdqiEmnxk6uhU3J7hJNcNHlKZ3gbk6EWcqVJ7TME25MckavB1x3a4J
ekKFVAZ93v7RnfIQhgHXxS8MCxYhDhMcA+dFWIV55sW+xXiS+QWxwWlTJhOO1NlP
ZzqjPaqrTGKsCgzqsfOK8MNg0CDEnHu3c8boTHHYn+TA7CjeaW0q6Rf3PphaEh6F
uTUr/FgC41Or2ok9laBF+DE5vJgD0jlm0OMZOwTjYRe4n3pv2TizyWN9AijqehPA
qwEF4NDxA3L857V4CGqwpGcfHg7onHaP1dWHq398Hc7ANgaDaFVxm2el4toAWUyp
ChUhmZZBEAZQi9iNqCmTSt1sgi4+EjpbSG4TNOW3qAlfzvE3h+ep3pDooe+EqY+9
iM6e/M0nnHBrRyESrdbzDXmOAfUQuJUS208GyGqTE1E7/D96LO5eOa1juQPz2WI8
W3pnF/PWvKlVPlYp62Q2UvDWhKP53sbcQmWwBmL8qUqZr+o8YKMJ0G1/f4Cm1LYB
V41/z+kAN+284dOOMCKioEVeZzs89/8XfBdNy4+B6NuGHvYpDqJzGpdKtQEGRlNH
9KtjsEgm8zlB3/EYQ6JC11pXLgjqC6mmqw9lmtlCXc/KToQMMNtm10EaXTU+lb5f
cfmJWCbx/Rhhk5X0OGy/4QxQQwAxCQOGuJgIs2RhXK0J0byJhnN6dNwYEHa8VY49
CG1bxe7YRbDFZ0MuSrdqbAep5hboGUzt+DHTW6s+fiAis72TsbKNKLe+kKj0uOav
z0VDPu5JS2xXpW7vwVQyFaj/tjbUPwvFL+WSDduUTa+ltn5dIdzraIdJd3ObjTOb
Vk8A5rRbfBmx6kd3lOKWvMk4HlinNyk1b8o9dnUTc7GshFwCYRR4QTaDOae+oeyT
FBuvz7hLi7F6N0YGOHzqqAgJ1NxK5exgqd0nUAqg5cIWmeKVp5DV/5LjyxmpINVs
MoFj+qZwWFZFX/hCF4MOYg6Gi2IUwW5OeYWsY/+xGXWC+uFGLh5vD2wHI1O+SvYm
4UA4dAfF5/z/fJk6IaB2ZHxtDGOMggX/gHuVfWNLSpkEX0X6cHlIZWxhyIbWC0gf
s0X88PFV1zLqcn/degFmWDcGumJojngX3wKKBNPl55FYAPh8rye+qDWYAU3DtVaF
8YQMZh04lmI2M8I85Ur3gIttVrIrfylxTuKga5n5YfUnwrSKjIid4T+/VU1F0l0X
niUr9oezc5gKdEArZ1NeXWdtVYOKoQ8qiEJBF+0Hi3HSLugPlTaqrxNO2FciMKHu
fM2xHPh0ytiUartoaXazaYbvmnMIeYLUztl8TAKQkZ0ycGBjFmuK5nAgejUAai08
WeT7ktpqa/u5A1Ig3s2qfTmrnWWi8/0uAbZjTzSD5U75YlUdX9DxD6Y/b/Ut75Nm
Yl6KNJzEXQeE3vkugUUyNHSrnxJYSnIzUsi50OCTMxBPiAXWSjyrxEhhZDXINUu+
MitFdnIALz/LK3vIyNfbodNEmwYgsuUwW+tnYITVfi72gg+T8ZzNO4cBbYTqiihY
UiyBjIkahXudLB6DU+ZjArqTDJyEYsinSQQNFqX7NafmmUjBVXvZrd9dBqpgRLZA
ECtDnngqIdAPqWXb4sBpIHmrGk7zyt2mx+C2twuOce3Z8EYGlRjtMjighxbs1CmU
1K4NTI9qPmb44Lz3QBSIPrLY7ghIiC20qxI7XSMFl6C+17GB5nQKygkJCoxpYb0v
y1vFcGIV+VBgSRPKzB/0nkA/LrZDGbOavgjYAXjdI5t1M6myPlaCYsQwhdPdtlo+
pUNcsE8k5Wu1fsrY7aP30rkgsMZ3tzEaLN7YciOER3FL0mTN3lVU3YEwFdy8jCjM
zxYJyzqRK9QaDmfo0dHU6cY2J8ur/bHZdddTFXkMTqu+mMM07mi8mc96dDHngtor
+xRvrAU9pL/SAXlk5qGbtOgBCoY+GMe12sMrmL8ZtaA+h2d05PMFpiRIufW1B9To
gDWAF0De7Qc+K1DmYNgohdl403ElFSZYcU1SsR4LYtk=

`pragma protect end_protected
