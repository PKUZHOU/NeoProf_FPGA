// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
DMPQ/U/RchbcsSqcB/RcYwbX9Zksy/2PBwLynB8espcm2ziKNFTBGzmZuU/96Bjp
bw8OQ9bA8/0QZtrJcY88dLwCaNhxe3Fxe7pCocmSPiRWdFDdfBZWoRdqdAAU5rrG
PP5yhVGp05n06Exv9BICsGzpuwgzkVYYRpgeUsvSfns=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 10560 )
`pragma protect data_block
uHq13S67oKVWhSybCgk7i85m6d76vUggZF5drAP58JC0zk+VgA4oyPD5G5Ax7lG9
6DNvVgqwN4PPKrgBmj6mwTWFc0KJpZpNLJZ7HZjPbsDDi/4qVxxuSCeWxSVttLX0
ATlOa31VeMifnEr+Eoc0G7GXGANhr054MjmvmzgwIBicP8e3VHNg20BNGhMswW9M
OUzxfS2i9/c0I4Cjnc0UdzCksUeJMNfVFnyVXnuOA/Nscpcot/Ab+l5RObB/6FTM
8NU1Y1fxbAM0zeOeagRc9A52g0j01JBsfS/FLmhOgi3lhA9jwtzDxtn//5ral2aZ
hhkx6m1bLAoD5mwmzLKCioLHNFmRSmB8xpgKN9gMSIhA/YJDzXUgD32h4qzzIrwC
eVaX7m6zfiw0Aw1wpj1Sy3RXblnupyShcHv1oX0WVCL5aayTP6CCOK2MbkwUUaSi
xlS/sWUHLNVnglY8lCyg1WrAYjStAzhSf0qSq1Xib+XQo5bDqhX6f+djaJNjdgsy
CMfzWCc0GV4VmVOa3MhQgp4VZQmxjgjQpJePVZplFeBsBRG3i2TN3w6TxZzMomRs
ZQ02R0u9XWTERjbL8Cy88YRlrvylNEoahdJtmy0tutYszMfNg8KEi8sdgvs1kp4p
0F+RU7yiMfFGdQA50Rzpo2cMDOSA86Pvq8Av6uaupz5GcanVYGMMauRt5fKXZBFt
4MKLvOQRJRK3o4b0QMYELT/6+01t4HPHLXYGbW+j78RcyDM6VaoeGDqO/1EC1oEB
7zjLMLY8Jt1HE0Rd4kE7Y5Cs27nrJvyZxbiCXuxeKNyps3HccUipKD4CcDIlz6vQ
jh3cU2lZxzRukcL4FaxLYFW+XE0pMosnERP9hZaBwDRpiyxDO1NB9CbTcsbrBKna
t71oaNpSp/Axy9rQ4N1pF6FUmsTn8277htzFTcLcXcrq5ywWgfqUBDJHd//wCijV
p/q+NUVDyegsJiBqCftK1KQPLsDeZ9T7T7ErJ3fGY1ETrwLD1Y0VukdyTB+4zM7R
LsJZ7hCmjraJ6V/xM0LvDXbyxg6nmPLZpoWMsIfzetH6v5GH4WV1T3sNMZ7VdQTJ
Kmg89rR5eHKKaTuAuf7RAXPdPpAnCu3/kCqbIuwXEvEJ0lFHlOluTkjcpQgscKp7
DWd/hBS07Yg9Je+k9QQezk/TdzwLHWEHiboy1f1Oeqe12Nw2pAkSam/kUsCn/7fu
jPrsE99CTB2UjPBxbEw1qghWVuQdxyfT4nOlq3yFevys5l+ovg1Eroo2qFSBr96n
tJ4S7C4AL7uBWFaXnZWUKdNzQ3WMh9HafTiSS6juJwaFUMku3/Iu31z0o17ZZ7ws
Bpv5BwrxfvJhGKPrtd/OJXrwn583HLq3QuA6hN1w5S+KoD/ajCjYanGaK0Ei5V6k
qAjlJtmjSUc24gIbLA9GfVpai6lO4n8OzpJtPnIHdzvZm0Izm59MC6fDZRie2Ewk
2/PhaTZOEwdW3fh7nVmuc6EPe/MrGcrt/0aNCpXJe4Y2w6jcJM85I8+LnScqMg2J
BN2Pr74lRjWp1qmWUUIqsPaoL4DL3GL98AaZcYCoOBL4Qwj/ZKXlW/UorOHq2md7
f06nlKNtgSQgrtDv1+20KWwRFQZzdwkfnIP0IOpVB7vi9GRg1EeKpKhspOwlVSiI
6vkwzCdUSE8uhOZ6i8mvmNAwOTJJDfxOKTxnrKbOaWEL0neTpWvWSvHT7LrTAgga
lxO2I46MWqn9zQwP65C1csOqNnfvKTRFOP/qPTcJax8Ibei9DhNfeCD9+eHb5gDp
B3wiPB5ExzsHOUt4qbq8j+W27VPHolc3gecn+OIjWJ81fMx0V0v+vZQJLVVx5xRG
UlaESJqKXFX7k+LL9xqtjB4SWe2zMV8siVrryOcg5dMGAisTocP0EY3bkHKk6c6Y
NffAErosEHKNjH8sGAAaw5VXNwgLrqPDjoZZ5km/7i7+WaWiL0wo7uSzUcWDk4SM
BluHa1Nkm5L1S5XLp8q2Tf+p9HNHySDtMaiwQ2vODGzp3sfay8vudMj0perUMRJh
AueN0+muSq9ed4wfOH+tuOBgtnu5RnfjO4sGZhxAT13qfqay8716p0lKsnnpzVp0
MvCPjisbNefNM3BtFXhTkh3/Sl2yDSnT7+j3DBih7hUzOKxyXTyfNIwCsGYltv/t
JWuh1Ueh7KyD87GKjtpezno4O7zoFFSe3dcX+iYdrpgWOqyEJ/GOp+G1fvb2UX/j
JfQNbSBu2SV9ir+JeGSCqgH6j01iZkGSX75tVudjRKSA58i+6uzC7E9z1QhoLTSu
9KFtrCHe0UjcIisuuuceedjA3dMqdEe9o9/Hb3Q+VkxeyIgF9wF05jzuEl0ds+M0
ykMfAMpTgwnRjF9kfKBcOHQg8xCmTyqv1Jk6PRgZB4i8WMaNgmJz31tmuBK8tZeH
WPTltNRAC/lRZmt0P8ep9yLhfJdT5Dpp6AoaaXAQOf8ri/I51PpBDr9UuHGyMSUq
J7laLTIanZAoj7GHeSxwxFLqquNUOcDoaRji4bDszVDqCizPoOiy6CERRPtZxGaB
wRjyy6IfIMOFU5tMVJN92iKrNp24Rfe9my9x6Hb9AnxAWmlk6/KCkV2gvOlAXbgK
XA5B+KmCp9AcePCKv6oW1DXiijyRDB4vB5Oh1Mqei/SrXB17s9UwQQtn+OecE0L7
SjHpBMRCQRr7OAornZjO/n1/5OFx5gXWvbtu3qBc/x/uayKvgWFV0m2jhuhaCIOb
b5jRFp2+/tZEIDuDeBxwhXuNbPHaRRT0coG5XFX7ubeffxUoDJDtQDPxkwOOKb5j
B9JI6Br+u6cQnI15UWo63g022O8KmtiqCOSrCKtbj+zRl/7MhWytIRLdcieEAkUx
mSbXRSuNPd5SHWvXbyWdqX4nYfutrRug5wuMFUuVtD5m9Ga5xiTiLe8hKXIdNPE3
SYjJT3q3HaWJLybFDsTUmQGnBhL8/Hgy1UE1hzif2wjSYdTSjx1DQ1oaxrJxR3uL
+vtI/vO1T/magnjmKsGRQRrnNpOPyaMLfyvADuJwxyEby0nkoVAXFbx1+Qirhvwe
2JMqnNhAqtqFLPxV5afYxjMvvjS5K0GjQMymPD1oClNtl88ybVn6Z96OwHjLkVPn
dvm3eW29pqY4GhExAIdX5Dvjupe63za5gJyWOP8jmzViDUK5P93/GlogB9ovx7rF
zKO68ui7GZi4cCIw1dxZm8ZKQjeEprtcup+MOgk8M8kxMAtSgaFfmMyv0oXEVMF1
EeW9O/fj0oSFk2CmpzqA5py0oXEQ17NqpRyAinVsdRA1tk0e2+JpzsCC365HcrOt
yGdtbf3TQ2IWBoyLQyxK+cGqH++m+DrSrXV8hfj3VYJS6T/C6NTTguXsx736PrOe
xougcHp/XIq3FkorHA+ZvPfrq5tjOwl/Rdo3tIl1uNTcUCtQCz368DjweCrKTTwY
GEuDK/A2R+oLp85XoCShjCpCK021pcGc2hU3fc3lIjrYpnMFJU+eUcLS94P9wZcT
suR7pQMXcIVN8VfS0hof8CXU2TDwloxADDJzNAk/9DHtjzfjKxj68oV6vCYOmYJd
F+kbf9mfHf/nb3gFwIPXnIFOL0pp/qW6/ecn0ETFX5une4Hzo2pubflDktQ2Lp06
IpZdVs8eRrldBNIutQaCjA1SuJA9H5g95WNpfQY4UXfYazv+lNh+GFWogjh4U7/G
ede8rPU7uaP7myrp0I9zmyOVlMcAb/VCdBSvLS3qzkzxe9wg0IMECdVZowAUJaQI
WiXTX5zr8JB5RitdlCOcXbLIXAPplXcdkEl2PAmIhmoLJLQmSVTLqo5XE+GcYtcg
gbrbpzJboT48mlNGRa598V+A5h01zQSZQP1M5IJsnjL9lsKvQg/QcwohC4vR4ozl
6iNRng2LmcbEVP7fQsF2zRVaQyzMgc77EqtHsKagJzNipMLtt85+IhMO7xXiBw7W
4zxzniMjR7eD876pTkZnQNj+Z1JZEsehJXukYJrlpOyqykRY5Hfy16UkSW4VjUaX
x+uZMPbyzKL0HywDcHKlsJsC9ZVBAW+NdVpBejzWEr99abwtl5rY1xsvGQUvH0kt
gqEIwr0y6PnaDtpHdJQ3cfWEk2vkodUq/ptoTb82J9xi++FWSRZTS6teAIIMYlZV
QI9dOd4GlRMjgzqMEdV8XG5ntbnbfJC3OX2LYW46DLh/QQqylwumDTBWmRavjDw9
6zlRVhGX7zTLrK89UXgraYWxz7VE0Rcqnn8Hamf1RePyi8NVCD6INg+W+fU5lvM+
Alah9FseqQd13K297fg4hxg72HoulKAu7ymCn9M9/9Agpittp72mi1qwRkyn1lz8
FqPufQOY/sdoCXFBKIHKq5h1yk44sOe3m2XVPZGti9MTo9yUZT+nXGnZBQxV1QDY
25dE2keKct9MzZpZoVZpr+iy0bF7REWOBqcpMzTfKK/nHvMnRNFITtKvkAXu+i+G
vWGqHOFcydJP9tkByFagkwOqE449VwJavQ3Hm9KL/S1JYjPa6HrIG2tUfmX0Ix3+
Gh7EjsxfZbNK2xqQfYMuhBng8I/pKgJ9suj1dBLQ86j0D4g4BRG50o8NEQC9PSdp
VoVeh/V4vqUPhpelaOcrlnZZswpoa2k/yEU2nyzy4TNMHUhuy1TFfHgOr1TsnvwW
44d9eBhsvFyYI5mrCgEnZPSrVHI77wz/qMjLILJLEcod7+o0MCIpOJy7hwVSofLF
T/C+t0W2WbmkT3VVpywKME+2s9QSFG8A63Po2HK6h9mH4wJrsSYEomDk1s8BcpPZ
+1TXd9s8EC0xBygOa2zendqtnxTqCgYNbsuk2YiyVIXYVCtKEy1Q1EuTa+GI9nDY
lEqI1+6knnW7bo76jXYgLsZZqydb03PjxdJbOevrqk2/RVYSfw3WrtLHIpEMTE4e
x5tqU/PfCB00WGkIlrivBqvhc/ZH5fwLSSk2ixpZT8sr19vOn4mRazYz8tIdpzp+
zSIRikMqlyjIcLor/CTTzTvjhQpNggOBEVRRq06GAFjktkTu1iwKW5Dpb8ddWadF
gkV564anZtZ/Wz6z7UAzs2AdfhzKa6VAbW4S0lwEDHY+MXZob1Sv9VEgV7paj56m
nmdf98pLzZ/xVK5dQ1Yf1t7ThxDVVRVzgmgOoQE9Tu6cH7v6KfaJJRnPTin1jd8H
b92VYW97loSd8teX+9VRn9fvPlaIFRGCgqmbO/VETXvr0RYExWPfSQy5cm5Vl0bt
v0N2yy+T+BQ9mfcF6VT7J5RWMC86VnIKDFj3YroUzK4XQOTzF8O5t9H71UomDXST
KWBYaH3OHtD/XnmiHMJJXtjkdvZfl7kDiNyO7WFNcwmn5g9sBEiLGua9moTomw0t
e/joj2XZSM2sHaaxVZZvjv0j0r4Urh++9IKA4+btZ+SbhWSUkRwB8urCcyFo5mtX
L5eDdimZNGLWmbnN5FFACj4Z7qhWQYZwCkV37vz8tp+LRkaB2AdynaDceSsUnbUz
ZiBzcgq+Bf8mJBW9YukMIYwocSw21V/vFLIOmi1ZQ3KXhb/MK+y/9XaQlP23nC+A
qjogkG5D+OooscY8ssP0VDcWj+dAASnD5hrL5us6jl9dAQqVdBUz+1UyhzNSwQ89
JWJG0n3ZjSdNZJ4z8J/uXgJUUxgnTJeRWRiRL03eeii+VsJYDJZImi8g0P+lRdp6
OZMis3xC4ISSY/HHTol5ombkweQm5DSh2iyJD0zO1IPqa6ekNPrv8Eso6Bf2yFnW
e5+5oPMUAgXnDc2WWdGUN7nWnMBXAHRMknmw7tlebzEtL2XZQ+BglowGyjlLbbxG
3I0CqX6e99BkQir7QzDufJ3j8BPXRFxm4R5fjysdWtELliecVf5s1iOS0aF0xkCu
sIG0jK8YLWLiqNIhrZq8l52R1HHtUwYd+zqFcxBRbxZABV7Gs6myiPA6ReapeANO
BuT3LSUNhqG7PntpJFU6IffKhlNmZdllsT7Hs22xr3K6OADmJvLxBpMB04ld3e7y
ToGwImSk+HTnuuLBxkwJO3KwKiTjhLE125i9ms4IXO7M5pWVx5KUagGiLzHmXcVR
6rWK3cdjtiFREcF5TjhEaQHJCvcmka22Pzzl2sEOULtDl0lCJKdNmiHSHaFUhkPY
A9Ye87TBYUZ7VZ5JMu0NWN1LtdX7jCRm2TBN77lNV+22YzxM/7qU8kF8/PjDsBPm
sRhG8NOt/uwbVQNLFfGrPdHv5WrqHTJJavxvmqKUr85+RU0GJPCrcWe5w8qudK0/
nDqEL6IZHqCLeMRVn9T/xw8CKqasHBU70nRQI6NsAPIFq6+xVHZuNTwcDHqVNycR
beqx+bFl15AJuOmgDM7FXpc2AwIqy8iuG7NLtDFoL4AoxGee0i3bdcUWBuW2f+AL
VwFmmUlDRWdW49ausAogG88ftHrPmc5L/H/Mm5Ec8xeBdxlVnkknpRDmCqr07CkB
elIot9PITTphmpq5T5MiZx6IP77Kja/xW/d25Sqs58x+bABxfUJ9rewDYU414V5w
9tvrXcj/S5aS61Xlzz0d3DJ/nDgQKHTJ4l5s0YUD/TlZ42kr77OiTiMNGLQMc8d1
9SVtnn8fxLAuNBQd8W4ZQuCYPFTrr/HcmK83RPgzME9zEiikAGB2VryqcQWt7c1E
PPUsVQcJ+Dsrd7993oE7J/fmzbmGPSSQxF2tKa/E5bmxK4Ycaid2diNy8UfDoTCJ
J/kfbf5bsNA7MABv5+TvMmI0iygo9vjjVfTCqi2uNitmRD4AvQJDa4PEdQM3f4ka
2V1FYbfaokIkZl4fsFa25OMyYue+g1qGuuIJnQjAMJQJ4Ft5MYuQEIVtjv5grSw5
eH1/qylaSOOQOBSL4nVs9msfdL0QXZMH/FqbPtAhQjeLnfxa/0l4ermpb0+XMQXa
gcWPbMDfae+3cLweaVx1B5MXrypAK2UmngMuV/7/RpG59H906a52dhf4Hn3Q6SQa
DLCQ1PZ/kid52nalCfdF1wRy2QSZL//rFaD+PlwtDK75BJQ0jUBX/xPB+p8+y3O8
0hrDlovq9gUG7GkaH6excT6dzZl3+vPKr/CTeOI9VIwZvQMRjAUAPscFxIqey3vM
+jfD0RXd1eEClprqggX7uRR8g0k5Vfi7qMZ8xGHPX42VsKC1+yzDrrvUc1iXoPaP
OJVVjkU/CndUrRUMDHzGq8aSouSCgEy79pSizKuTpcCtfPaCzhOs1bucu4nnRiAv
iBXuSu5GA+x1NgoXoK57VcfzJTr7Xp8t5Ukw2rMUTiDcmwGc+ho3P/aHuDx4IwGW
lHdhfd7rRgylgzaBz+HmxKpjXa5dwLPX+DYB9u4MpcT80Ax5+aMBa3AIbY3aGaK9
cVdsjCtck1vGXQc45KlggZVdV4WkY7x/+J9AAwTiXDN245xggWGOO56QVNu2snxH
/wiKV7H/IljbH5unbsYffMr2o+LMEZJKTXE1/wfH1FHx75SfFUBxAOpjPmWkU6HD
2R6J+8E7j+DMW9D5aVSE8hrqSMFG+qMCeVz398dhPZ9kqLJVv4m/1suJjbnjptD6
lyQXc9XXw4212dIyEqt3Ww+S3yf4gd9he/JDO+R4tXfa8937mub69YgZRh+OIXbg
uLWnPgadkVnmA+Iy0FwM9IVtNkf5hPHZMtB1b1tqj0Z+NdXF8eELo76Hw5kUan8W
mTDZsD8lgxrE1uqSAG/MlFeT5N/t8mVBGCeah876wyCxsBsS3cD0WJCEbmOH47pB
bUuQuVxufgLVjInVTdvyRJIusVVpuaHFQuOkwehOvXo+zryxv930fMI1hVIh1XTq
z5Znvxc2dpswOESWI95d6P1uwL0AVT62ZFRmMFlxS+zOvwikmNDvytxaGhuujx/a
D6Ji/XzaK3Jei2F9gvFsV57FBEBeDtNWrD0pGgFfGI2Pk7ZFY6wCQWnO7odBUYUJ
CujSUfEMrkrv+xufzn3EJftRYFaHzVBR2KBkIu6TuOcyRRQnz/ieQ/47V+fn2vDd
81b2VCeoFakhl3q3wNAgX2YqGFo7mi5iDEgVqaSCesBqRWqiDh5aW2kNx7iNTeil
K9kTJoNPe60bdYh9QdqJiES0li3bvIGXr0slSIYrXrpYM4CjjNQqr8YINoMtL6po
5tjFJucL4R0qWrvqwUavg+xRzdaaYiQZ0w4k/CwQ27+LSp3if/lkWPkE/r1VEk41
z2e0xrhlLbLs9tL+1LTdYzMLUENq1xudwxOYR8bMmPOUIbZcsWo/Gd62z5CEUhqI
PqGxNKa85TVUVIa4mElaO1g2XERCXOU+PsLEJ+3OkUOds4GfYieh4J1bq1HiZ2Bp
/4EneTuKjuhXyVnPBcwu+wCu4NWqiai/N0trQLIq8yZsG80S15fBpqP0ZeWLPQSw
uCMRodB4qfelnkr5IGGjyqDwy066XlIZUhaZ9tXYqNl08LZRWGNQtRUDaIq3/0sK
JJueJkivwj3ySy9jpz3JpHyE8Rw++mOcZcS5V652l0RUz77fvvasLUUReAzG/9fJ
ly0+lWvcs3ZxiYjHh+01Mo8dH5BAlh5vcnmvanacqpJzlk5do6UYfnf+8I7PNnVX
Zvkw/5qIzMzQLG9/zYUdyDui3uwl5anQPMwtdYVv3YnGm/6YAb8AqWxmkM83XdEI
ifjZJ54joTfczAkf2v9V0NwvoDNiwZ2dbpMWyq5bqCZB5/OQFFUCnN6NcGi5Xhsw
VYP3d9hoX/CoBGxEjxrK2xlE7A2KrzCkKMoUyNMLuywzsIot8etBXSxdueZ0CpWt
+GuQ1eeciynlqGq37nNkHIUUU0lMDxm0qHXYCoXNmnUtzNrb9/Zkbo2qkiPQTUWB
ARobbu3hB6iP0dCMnTZfRx2awNq8s/wsFT3S+SA2D51zBL5J8AJkVpTz5T0daIO2
YlwAuQ0omagRv7+b8WeLdzEEtvJKMvMmLaOdRbAYHxyZ2zzQ316p6oqB6W8vaomy
eTnAqVxeN8cfeU+ZRWzehEWtJZQjsuMM3NOQlRBqPRpjWZM7aBz52IlnBjrmAHYM
4WU2LwBJeOP4GOwO6VZpKXDwQ8ieS+zRjJdrEhkuW5G9O9HwaNM7XUe1qhmWiD3X
SLw7LWDJB4KKxzt/BxrdwiAXsTksz9YqbsahUcd1VY9f/EVvISfiDOFINrmZKT+4
7l5GBMoWlqCWecZPwKV0BPXoDq6WoFYN/Yl6CskQ8JeUbS7f60M4pSatrnzEcOOW
Y9BIkVZ8C0Jw4WuZTv9A50CV14QWmAvduReW8iR+ygstXC3EprmYUEWF3QPb6mgK
EUi77NM4PJ1QMWtJAjcFgNYeoe5RXJ8A1PSjJRPGVJve/9PIMHzjuJ00m6Dmpdrt
kjFKH3oevRFwTeZJh3rkplXJzNcaV54VEtUb6dEgXbpYC+6ESpPRnaU6TxsbumW4
o03rfGctVFwo55lWCs3RGCmnlI13ZwMTYgEI6yr1F+CiscyMDIUxRLmmZ79yYDq4
spkfzHhO5rDo57CmWbJRv+EURwQIbpZZktO5ZD0m7PRyNBFKkOUc5z+hDntYPoi3
yxQv967ons7d8qBFScTsvBSkz18h/K9C5cEFyfn3jcnZpRnZO0IXIKRLVnrHhfVD
uND4j22/Gny3wkmXxyRbBtHigmgSmLyR86T5n/dTIOhmEqO57eNDohQx/Pkdi4LP
vI8x7d9iNuDVpuF4NoaREAqguocJDF72hh2sVnO2mXavWUNjOtxn5LRS2e7TZzKK
GSfuCdAbjQ8DyamFr7dYc1AQm81cPbgHjqPGlAh7uJAb7ea/bjneuoUkgRj47+TW
L8hVgi+0fuuuLiGo20lPMMo6HknY50vAs12rp9GDatl14fo8zs6DF9dNL5PFCQe0
OZhmy6+Iw1KFuIEOAxh808mtdZS/8zfNBTeEvHa9xnv1B+hglajVi3i5UgRgkwtz
1TVpz+HUIOX1sJssPnbtY61yqS0YclXUqb31nv2qKoyyOepB4/EiWEbzpIROpzRp
9q++r2oNDFUtB1DGWnsHOffkM9BRHwGbTAr2sKyDEacfYq/KxoqTwXJOMWcatZ1W
clSxo+THBSS/Wv6+01KqHQgjTFQePWiH/WSTjHz8ibU+00NBY1Lm2Gamooc2bBJV
Hbe2zwL/ZkXtCtRObcFtJ/8puOgDAuF0zzbAQ91vFKHZxgWLhwJSJJZxyDVklkRU
Mia8EZPPdtXy/88eKM2sX2+l6NN6Ley6GTvXb2LRxNgMdnZrQRWsXpTU0OlpUbZR
HVkJik5bDOFJUTW2fkoak/nx63v32kSEKTm3psNgEjeYfSg9uVGuKlM/K6f03e/n
SYDXvUKxbBmCTxRGSXL9sdunonaO8KdBD53xpXreokbDvBYLEaaly2f0YwQR0p/O
KXFCLFaH6/CQxtWj3efn55xwYpBqxbr7p2Lqfk/fYDGgb5a+j7A/8LVMth7VLFCP
mGy+qUqiii0P9pZ478RCa7aU4REdulZ72+4oaW/Hej2FKPcu7SVtDIoNM+kBi4G9
1EMx5p1WpwE9hcpTvHMxgDLjoCh0NbYMB1liRNEjoYMv37kW7i4A055r+EltUWEG
onl5zuKOCNFYhBGAFksrgeEjPYqUGVHWCz60KwQTfPn8FQfQ0Z6MrKNtBJiTlnyO
n9r9wlQ/Sp65OZHluYsD24ApVcH91e3s+zhQJwGezmsZiV9R3JmxtnEPOF8DIJB0
cBjl6HeyRKgc/nDgEosaeTXRIThkqiIjLptuAJ+7g1Vxu8izxeJ/g5S+23EEpHwW
K/80aGVOvyhfIv6DMo1IIAQFdQ4bCzjbUc7VRWT3LWrm0h67G5QDM9xmDd0TnI/x
8X3s2SQ8yVrEODHU3RPosbVAWlJwOfIsL12098alB3GjXoZJsucztREbLlP4z4YI
dyBgLd0L2rhgmTZoiXjELR/geilwuulQEIX/ovum4fF0annN/eF//dTsxYpZUpwP
YqeUpYycmLIhNTRXYof3QnlC0LwYoeP8bCOtw6WQjiilVICtzHP/KIaN9eOx0BXv
mArWprgXcRSEIkrerwf8CDw3C0H2Y7JDNAjJjNSXREptaoS5QeuV+iomUtW73Mwl
7BwRuT2ZRgzxxQuNsV3jFnoY+hF3xj/XAUR75lnZ+RKtt13Hr6mbuLayKIAsnoaE
4FHsibDVTQ3s1s8yAZlBlxLSq2zGYi2ji8ExT1FCezrZ3hRpQ0gGFQKAhDu3MuLS
YndVvg3FWjq/A0fIa6DykJclkVLHZPjNspiBHver4jtv+iHheYcRy5Wr7v0gYujb
i2MiO7YpWIXVdz0GCTAXK4qTHfC0sVZS7gt1tYsF3gg3QzNGx4KiCP1H+CHYGT2u
64mD+tm4/lVseBC2GIc2wpGwVVSve3tAbziYLmmzWaqMc4LGzVM/X7zEtXvrxowd
QHCBtH3Y8JmHOJS9t8vgJnKvRA6MC5ha9nkZUZdYEiFYEuiU7nM/hhpR23dtbNRn
dM/9POdYM9IQX+DW+bG190Ow4heCtNZ5H9aSKNQtu4k3EC8ifM7svIZ7qys7gqlZ
tbZ8p2TgX0nY/PjunoEOb/9uXM5AYhf1qHSXUZdDsd9k41xxmooHYni0m+SkYBQK
FZ45iZI+Xnse2n+BPjisomucr2i1u6iVzF+16wR+jxKwNXIPO23wxIvlaTVODQ0k
qoWw0d4izvlNZ8sX/8RmtrpNSyqzxj2toWbK2Q6bx9IcPCsYLpuUAbGIIHreLjAa
foabDbqV1fbSu+y9cZFdpP/sScv/81KqLXr9a30xPrgoVC8lJA8MMfxp5cfnO/V2
q5XZr9ldcF2Vc3d+734STGG0TrUtyJUWYgH6t/BeD+hxgdErg1YdIyxJjUQcyA++
ecqEA7/qRjDTm3pBniw4V2R0s5IcXnvEZ+IJceEIUe1bXvxCSHG/xfkRc2rfBY6t
pQK/HH62yvMMgTDEO91QkHbgZfdkMesBk3US2g+gWP8DP1Gwgce2U3ddxVy4mESP
Tq2exhoBa2iPGsB3M1cJxQUkGAoJcH2rvIOzsABnQwYvjYoRqlIIKytyGCOQhpqu
wMqm2y1ZElM8hC2mnWLZWJODtMcHfgeVITxUgo/BwlRtgkcUIyqBmvjeApWdWVkt
rHMSzL5Mw0Mlz8H3DFo/7eAnxTG1PKkHRdhpseJfw6hzpFe8cs9AiSHdXHB9nmFJ
n7q+s7I7yZjvYddu+EdZX6aP0x/CAd6S0cUaJcyrMcqTcB9vXgeq4QkdUlmc7v6w
3ym9m+niNBABWtfkzjPft3ahJMaGFBetp5FsqheGLDmHrCqSjS2w77KdCMKcUbb/
WQ5ijSB8c/ZS/yeoZpmYfuD0+aSyv+OZx/T1Dlq11MBspLg9e9t0QuMR0nZ0BSVg
NEbJSi5+/5wZ41sM7KCYvQ8zv4pwhaZTbbZubcGo7QEh77AfBlWEjhsc9kJonJ5b
18kAJCmQNjxWpGQAkSoZo7SFOo2I1AIbdkxLq4QG2cVbqWXV3PKmjbJhac/uI8ou
AS8SynFXNt8r08H/8VgPjIcL4dJHjxdBYdxGA94jdk2MFf1jo324yFQVeJdyyrhd
SvRvemFPm82Mya3nHQPu6pDJT4t4Zne33vtqCsdQZ873qfjuJ8qwEf8pYKVQvZgp
jluE6jT/2+5RHuKPFxQCOn1GSyzGwfkwAV0SnZm80aUzeJ5BVE60DntP5VZM2y5/
EWVlOpF5UXEEepmzwEygGq8KLvHhbZ1zVDhfxfNUzXhsMBY0zexQj2Zdb/R1tLq5
zCnBVY/Jy1aJOa1U3kCs2GJh+4YBq1ofwTUXMgvX4WG/N1w1BE3RfMdce0yw3yb3
F+kmgwwkT6rIMq5Vd/VZ2pyjoHRg/BAhWp8VRBt4J4KhplbYboelcZJgIUzMkW3z
Cpjnt0XhTCF1+fI2W+K8UfvXWm+F6y4LltAvMKLpSN++kpMS/3NyhzlWJS1sODlG
NeZ/IG4YhGcpxGuUNzzd0EV1nrC/zp72iVP6F2pkD32+rHx12zCqZXWWF7OJuuHt
SMLxsx1ssYbul7N7PLYJq7DueF5UCRLoQI9owQU5IloAaCeWlyJhYJeDDcEdUjBO
XpcYtU8plIMgVBaQT8p+e2AcncIj/bwlaRdL4BYZDURP4yEnqNeRLqJRoJSufugz
i2GqANmq3VWMtS4tWn7C3an1/cUXdsDcJRZJrSUoZPjfAUPC/di/PRcm/jSHi3UC
f7YeZLNox+CclsByjSVlvkPNZYXzV27xdcY9oMV8D8sGHonB+fU62TCNMlCSlU3N
S1czFgIHioFzMnHBDcbkHYQpjHLekq/qe8HSkCfLohdnl+IhQSUO03bs6gIgM4zu
LWBhm3h3RP6K7ZBI+UHU4Zb/kNaZvIpiUMOoLSe+HcAoe2Ufn8hfoD/b2sVW1rth
6lpfCUNh3Hm9Y6VPhFpmNbhDZYNmoUq486ajwwK08/WXmzBqFoPtVEd5i05afgFG
mJ7SmxFGy9EAcn5LmrCp11UvZiI3RDoldGdofry1yUp5FquEsy0XlKNgidKmKF4Z
iO/J8Gz89NE0dMk2JbV3cF3Rvqm+UcW0rOavEY5izrm7Ugh8x/2418r4cQEF+ZnS
GLnWSkjyKbw5bSTzGmUSkVnuoc0LnpI6J85WhMf16juOcxVoEkUH9RS192UsY7Dv
ui7KSU+r4csuN4Qnh9JIS8AxnzzOZltugvLQSLWvk6h5lx6NlwPefmTzh/97DdSE
5OG0dEUpXlZpZkCjNqTf1JGxaxbxkiUSTuk77bAUbOjdSNRox6wfMd/6pumOnn+r
+QCos2L18rQoKZk89T3Lsp9wHCrhFKwgzf+q9dFCz7JSwbEzDf3oPrnq8ih8wkwo
3/X+gSRzVAJOYQ/iCzkk/E/QW6lx6Q5wBj3xzPtjHIsyBWIQUJAGuhALujTjLAwl
ej6pQWtL6nE865BPpIgz63J0LXUAU3EtiJ617rJ6bc7znyNOL+ffOgtfWphnt9Uw
x2JXK7hNYqRmb14i6IwvQORmw4pZCy3/UzHdmKWVWZifoMkR0wpxRGvIF7uSeUyx
BSsgmBSQqWYaSoa6T7heFn6sH5Bej6gmE2nxCndEJ7eb8+scoM+kQcvRIqOiPtNo

`pragma protect end_protected
