// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
STmBYx1+mGHf0V4yl8Vrhl8YG9C8a6KyikpYokQaqBP+IxXR5sH6pKwtvtrgtgN4vrY7vA7Qi38w
1NsJUdJVfcRwM8xWoo3WpafFVfxZpdI08jRiAHhsV1zZFVcakCvuyB8N6hmtYKYb9zc4M6zPu0xv
82sb9wJH4ITo3YUf4z+YlyeApUsbSD+nHuAVR9ikN2EXefa4dPE0eKG5wfcJ9WETAQiwnjq1/pvS
Oe4odMcbeRN0cEaQMrSy6W3doaBmGaHcPuSkRIZLUkdodAr+G2YmAy1xXKAm7M94UTsW1RnsVTj2
xQ8z8rNciyCUzcwVy08rOBIrJxoUxeAAHGzm0Q==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 8496)
4Ui4Pqm5b/hxT4pAuoMLG/wRqtniDxB9HKql5jUS6TQlQksR49aRTHBZa4M7cq7J5OkIbODN7DIC
/hvpuM+EbnWvizzqnGWrfXgXt9PaYI2Xt9W+OLN/nMw2rTyzzVtD9IMqYoecu3Z9hmwtZDSgzE76
iTgwGLr/u28by6yJuG0aMYeMIp4ZnB/mZZFNS7tyGL+WJeogoFpQ9zGel5rIDlaT9ueQ9qp8sRJV
JWhQHdof9oxIm6uVwOjSc96LyTJ07dMEkACpU15wBAPPajVKqBmEB796s/xTys/mM8/M2rAV9M4O
nyMd0hxfvpWrH2hac5ydggUKcURd5k1RBHp8CzoXo5A0naGp5HjpzjBrJ7tqS9t+dwVAyUwa0RTB
hh5JBBtlreZi71WYVJy7ioAElR3O3IAQxJxOOTV54r18Q+Rb/i2jGYs1JZ/+/tcQLMUzJ4tOW6LB
ukQYMmpsBKkWF74C2qVO3iCTtcnfLxqePG/y5oW65UPlQ+wfRcGmvsFEA/SvrC5v9JXGoOlf0Sd8
OLEYWCb1T4sqpI8JY79z67jMU9avDS+FrI/xBYcN8lzGu4bDXQzZEHTaueXAQIApHUExSBvr33Ko
9343ALbMq40SS0OF9IjSQMTkYAmRvlifVZ5+5Qyg3BBueNa+eiu9cA0UHl34k5sOecwz5P+FxnnL
8kQK5VNNUdp5B3bcjUaqDBlZL+ldnBl9TgU+DHRl80s1RgbspZtvfgAE+r9HbJEPVVsl6IvI/aON
B1wjcpiBOuQflt4fOlBNM0sy5k+9dKG7lKf+HtCdh/F2rYT+Fsq+XDl2qlxm2K4kUXqtvAz1K4Nh
qLIrtnCJsZtr0Spw3Npy4ZvtXAGxN3d4ONpYolOgp+Jq3Or6KiyacgktPa6o2dCkCJOyyTo3rul7
wlY1KpAkWZ0pMFvMcX7eKp6yZ+zBIG+xarPwwzvutkZHptYwSQFB4WJ/BtEiN6LnxL4e0XrJdKxY
zGFWC2HJjTYBtvtHB4eUQ1qt2nOLqouAPs+Oh2Qpt7Y4WeoFAj2L1eakGGiO8AXtn8YyjQHBdaYD
wglysh/nmY3axo2zSWXDwxoYDttPfKY8VdRjJkrSZ2P8KxaU4EfvrflOklmXqnosx6geSWRmOhcr
/Cz5VXxfpvUgDoQ5gy+kSj+zxwe0tPbvl3N+GGWibg0a298XoQ+h+062Lvr8o1nW5wVuiUkQ+P3U
pstDcdsfKBfpZu2iRtM7TzaYxFaeXI8wdsGFf7pPPcsNSjY/I9qHOpR9tEx8rNEsNhmEaly5OE9C
Zg9omUyyJJU170+OsMUvN/ojnRlG+oQGIqab/HMP/QbWruh4ayC/CjSrm4YwIlR+xoQOSZRITpbS
rgxryTjkSxdfljnS29mZ2xB5BZRlGjU5Y1HYo5HWtwToXle9uSHj2OBf7kC1itrlWjfraRLTgE5i
YH1/rMXZdU6oWYM6+yN2rO5eU00+rjH+59Rbco53T6+h0yuB8LNONIgSi4W74TV88T/7gGKSfTst
VqXBW97xeJSYcoCH6voDvqiSIUgXVH6P/N5nab0wGr0gRKRbwGkBPYBTwsqCO5IyR5XyVWUry7fx
SHtBAe6c9iBqOIsIE4zI+93Cqwwhs9kzI1RImRdm7g+eLnOSUwiAi06KocMBnFT2GydlOhfiFfJB
lt+qwTVDmLlm62tnRWTCz8ZyvE46CuooM6lH0oVR1Nl6kS+QkzfVBlViT+GE5BGyADITitZtbTC0
GY1N7/3/vdh4rIfx+Gk1G5/xDfoPbYggbdgFhcwVPJYcod3CMJrjEp+6AnUh7s3NG0wHdunxCFCS
TpcvSzSCKVmh94b9kUPhFapG2JzoGd1qLDAOdrvlrlyYdQ3nLoc1saqe7zdpJscG4BRJVSYDbnk5
HKTQim8UaFBUZT0hoRwpYZfpLdAZoQA4W5GjD04p+hup9A77E7zKbWQ1SbxvW3rjZRDpBa/au3OX
hrE9j2CWp+kq0OR3jtEJa6lSSGLSm9NfNaQQ2M0OrqtkEHbK5eFKDuLFWsFM342WmM8WAg8a1Z/X
+wMFUVpxSjMXFQ9RVxLYXZ6WOTsOXuTRSzMeLbEhquGGhr9nIclFtZOXpV781YmoRByza2S0C1/w
27+7fjMnh22P0GtjuRl1YyorbyGdowAnvsZUwdUIUt+Tnq+1XU3XhwbHwQ19oLbPQYrtQLociWS8
S+mkxFbRzHeT0WVgz5bGJVm+UqwuW4Ck+3O5GKdQB/eVBpU5Lkhse4D9WVDGFqQIjWQWBit4O05g
eIYBRsLQoYBgrgCbUqlH+PweSW77tRhR2rVHXvptsLKSSQdz9kxsMdGnUkWIZrX/M5nHsugqX6tr
EiN4mSLLAuucIzZuXAiq/ADCfWwmM+W3jlzRfbb1+xfD2sUEg0xCR0e1l5UP91byypj4MFY3nn6l
LjYdpCd6B0JM55pEXazTCf4Oq+qlMk0RpYt6h3BgNu+x50jeMmfXrIjoPzPoNSq9kDsuDfW91j68
yN3JOK5NLj/ixAWFK5TUH9IHcQ71MvaBdXWfYWmMdgtCog0j4NPtQx+8Ap8jeyTs6I6/ErHz//sW
vGtGXqN14MnxDYb+IOluWf63ALny3fUUvH/8O5tFsEY5XijnYFukhYcYHOo0RCZdarxuBEUD5/7b
JtMXvGjbhYPbh9cNp2Gq49GGE0EK2APrEvbuOGxzXcjBVcoYkKhJX5Npl5QgLLMKKYOZSMSzk+tz
DdF6ivevdmQdGeHtJLIhg6tfKRGgwZTgGemvqbXKMI++swV7cZckt49A6B4lb0CkGk6Hqu2DZ9jr
A0BVgZz+slwPFVi8QdOBi2sgqKaJelyqScGLxqsh7Byl9gf4vHFRg872oKwTU5Qkb2fMGkzlgW96
l8JmsGtzmz4qnrlrL8P7Nh8sMdCIOpRRf8U65FcVuwZgYKaZKuc8Y4dvaYRIqks2wZR1FOj15uDI
knUzJIdykuO89TuSPIPY12xkassynGROF9uE7A53A1U4yt5Jsl2iLRqo+H49yT2R3LKnmWImqS//
+uneCAFGk9odQln2oExF0+uXE3DS2VYcJe5jKVHtUwfVK6049W8vL2RVjzfYHE3uRHQvMD7ZsoQR
JQ6sflLImOUCD9BUE9aKzzClOyAVagpo9Tt2uwclBxGQKmFOd1uYVGV7tfyd2y+wI8ZTO0kERvM9
c9cd1pArGs9yQw4HhJlQuAUyTFBJVMSX5rbHBM1Wi9RIYswmWjuqrkjk0/uT7Y/tBPR2FmCc11mh
sCtpwPbp0Jr9qcWbQ/fa4NWD1K0EBz6jguHAEGbY+hxjf/wm1nn7DJZVQJPosmc6ZxBnKqCWSZpy
5l6Sp+H8bHtzIiSqoR1Tb+Nr5cGueeDFPKNwQ2wIh1UNph7g92CsVojUUXiZxwgdawtlb+26SNqC
YPn1PEj16MEVAIVNOZjyUNu/jCDRtM0gWqTi2dEbKE1ctSAlqbtKt/F/sAf8kyGL1fqF3MP2qQEI
m83c6/23v9xnjtlniAIGQe5O9kck+lFo5MNWlvcEccRwFLMHq/Ht/SneeQaI5i2vV4RlMOnosNr4
JW8HSFNEretaEiG7aAp4A4gGIJph8seb8CLbgQeFhXUO7moZSe3Lw5nDBlxqWGhpZksIJeeEkJf+
aBbTV7ZnnxVP4301CNSdHY6F05HXeFejp61xKdS6Np6G5yEK+FP//Ovp2wouTiRzheQwKKO7TS0P
kydN0uXccj7Ruz68rOHDfNrc25DeNq94II2UpcjaLJU298Ilhcshk2LdjMCxkYXKxcSSdSP5Pt41
XLEuCYC89XT4qbv1i0nvLDV0gqCX8rC0W7awY0Qj++R3oiP6o3MGgLujhxtDsDLwWykr+NQDzncs
tTs1QxMJUe6hYMCWFruBhhqfOjTtoA7tcWH5u1yTFFt7cEzW+Lg9nQQhFNxUuIkDvy/pKWoLwc14
02/vwIJiEigZFkicD8eZFgzV1uYyWKzdN/+CwJtcnsF5XzdvzCa0I+fAmhqV+BT8dWAyyMCed1dJ
ktlYrXXfFsDDFI2nSy5AWXE2MEVxqncEqzLwAI0oMIVR7EzgPNYyWry2o7+5Vr18XTsAuBTRRRbA
cLh/4LQJH2V19n+Mn518Rcvzb3/Xv3dwNY9+rrkR5r5Xq78sBEIgrpCmtV4BNgOHXedaLeGWk+1X
RW3fgco/wVUFRs8eGASjnHjlrZGWSPjC0igU5YbPHwwAxAxPSYm4tRwTxhUbyrcVLiBctpdqs4cu
X4Fkm0IYdStNRuim83Aibw22SzG8FrXfpIIZ8ZT3EE6wg0/NwvZPkQj6AoHr7hqZWB0Xhb+3VAcW
ZAmhHXvgouLbzVgckZiSvRFOAbpYQ9tatAvm3H9+xyO16kv2BFTMnLPbEA3vq9o862WE67ABg2vl
hrtrhStE2PQgcfbKhuStoeziSKxJsBczZtjb6cX6sy0YdbU9kLSjgKiEhpVTcwdNKGou9bwuNeY9
XI7ZLFi1aCeegNATrGbvaHSDbb9dqL0wm7NYisplCPn/HV9Nbh3QupZTBkCsLB67bCuWHdLPG7Kv
9cf/AvU4VT6e5N4R0TtElhXWwW5FYbOFako7BjXvyqeXP2xjBBY5Pa2oDe9fqM5JR/0A5qEM3EKJ
fvNVW3dJE/GMdjwFWpQdjvYDXVcErxlOYsfQC90s/UICUypND2z3T7pU7ZCjFC7Cmmv9bDy3k84o
X5YWfylKmeoOhW1Kn4fCsiUj9/BqEtfQQuQ/nHPemRcQNokQOkF8yROzsRrwV76d7l/jo2p+TjcG
eGsYGJNKUxV+/p3UAHOPEB9Y1OS5bWeLcEgSXB3boekA7K32mpgqrJmTWL2kF9gnQe2alBgn2lJo
R9uNK3Rkwmt3y6hnDCWFXJ5G4yj2y14IZyP0eotb15MAexA3/F02nWm2Jh20L7dUNBkVrbHgknqD
foUeYkUbb4kfMqliaFXqM7H7kU/lA5Hl5i5QCONYDnIh1nmgydmkIVNfbEp6iSk1P2DHMeA2ySeO
lcZUZIEVie8J6Eh7wrELUNdBeFjfkwq/fVfdmjjVIChtXIKH03WlxEt5xjaOUguWbwIxoTJz1FlP
K933o1tuQjvX9udpRirzoTUJGK8BEYFO+qaElvbN2jaLIuUiJY0LvAJUkYlN+tJM0qu+vchgwrS6
q8QIT/qwpu8YDCfH6sLtcLzy8zqOYBrF2mMRm/wAqq5rIWhiV6Nq3VWm7cWL0RrTDbj1JJ7IGrfB
Q3UzgMDI+vkVrbw5/20R70PeQkbp7hA60C1nx+qRXDXJz2z+1RO3c9oEXS+5RC3OOl3NIPI2Bw7l
w99BkmmW847JqknPZZRUPErv8SFs5LZ9l8fTGRTrK4ZBN8mS1vRtpWlNej89kkBlIMASO+aaAr7o
Xd/qJobEhm4Su/rxmK+8rasS75HNtJJz4h9H5TFSGqKBdPOQOvRuMmVbu1HCthv8H8DiuaPLZDZN
8zVl7U/kubYJypIq/y5zYWPJXuJ4/5unavD6kRbW6weuHAv+kGW3v4ZE5SoG1WbikxNNWwJQZ7jJ
zAOkqzHLQ6bcZaUAthDQoNSPSshuBOvZFqJVSebBTLPB2QSeOwCtco0cF5i3YFGzgx65edy0dhAC
Ca+SiTg+zXi4ILPshTuqO1nWhPNCAppJbGqNjxzNsvp4Gy0Zfw7FAikn2hiDi/022WXa6tAOJkzu
EqUS+ICUp3UUTMj3xhZ019Qf4Ze/Rid4vlgTBu9FShxGqhavuYrbPeqdDmzXaRmwtzVuaJct2Cia
EzL9xTJlnsYTGmuW+fA9GagODEtYum/9zkyDkYiVPG8LPDdziXWXToYH4FTJemON5C3dVjsEn0yQ
suBqt6MaTk09Ptj6hMmdQ7MH58Dj1W3hMSkl+2EqusBj2ePCGb1WmPwlMjcgRKrk/nmnRVoHzRz+
UojjOgL7oDhkTm1xnSeL/eL4W0gzpl/N9kXC+XQdt6tYvi6XO4yY68IKV1YGJIktPxEVB2LSDi4O
D7wKzkg19lZJ4xsBV2BmJCE9Yw4yoQLa0LTTIki9MaGWr5QvFakzCdDenhv669xV6F9xQrk4l4uD
dSJZXGgPt7h6lIwNoYlVP5Hx4/fza1SZ7JGXYaPXX5HnmGseFJnLpO4y/HKr0ZF3lawsozJHmNYh
Hhug6IBzDAZ4B5Op4eK41h6tJoub74mDiFCeMYtuDbvoGaSdRO0nEdX5weir+y0BvUnxJhMZaBxF
L8Cln5P0XdelIEWkcg6+R7WFfUIHMFUdISEjZA6h0rwLBE0nBxlWdTgRHuJT3Y6Il+3hv0QZtusC
dj5G84E9ZmX6UI7DSArVBTmewWhaTtXz71V8rSr8mKxcRxYNiEzFs51UyktmNr3W8kkPJpvn6R/+
SxBhgEvL65tdAd72QK3PZeLs1Qo1oXy489mnOBvvObWW41kMc5xqZQeWjqpGtZlnI7d5yYTdpi9C
HrOOnukzPbdA+ndAhzrgpuXFXFQfyi3HGALs9HGjm3kP+Scb9s3gvMbdg3Uq2bban2vaJhWsjUix
6YlHiHI3pXcHc2rQOFgYapHFsipHlM7b1I+QRJ3WDFabN1Mpu+gV7b2PZLcBDl67Ed6lbeN5FVEK
r5tU/2G8odTvDCvddcw/WrXM4OWrmJX2wt8pKNJpys/GfwOnr8tWGXeBzka8hisxvH3EJilAw+8G
y99pRG7kIm5hyJwHhwNiDaIw9OVOkxzIbVluvZ9d/phGGqP5UjbVdeX4TR7cCb+AXt5SS60G5BGV
owzHakxDY+e4Qc1SlGvzddJvrlzexxxsiPg3KTFj/1LGhvYj6VrOR2oCwdmSypBY3LEfcYcvomWf
BXOcz4pGr1zYfAB1WU7nogXku4DisvgbGldNZAxyUn6vwpNYfOXA15GkUL3x5Ajz93LRewlAdRg3
rL2CA9+O2C72qQtxA3C7NSqPeEbiZc01+s1QV6ght7nJe/E8osnP+DX5zu7RQ4SzioLHEJTKbUwl
KT0IVdp5fWS6pIEyz1ALXk2KnSz6m9SLMPzCjDfCXuR36WXgeaVahwUegQRjoRYz5VLfcSOSyNwV
bOfBFfC6vc0zqM6RwtqV2P1VA6rtvz0mjNAjeJ8DmBMWRswt2zBQZIrSUx3+55eVESkBCF/LMRmR
Gr3r7OkUkEmwWAThYET+2Dirxu7HZy+6+YE+ISRKe2sJOpP0Fp9Bww83+wAsYye0El49pfWGZhWY
KK71cCG20TiNnmJUYPPx3+my+jKL+hfv1dG4uwcpAVztJHqca4SQH/S3maR/XZNtSHBthVTtb1tt
v+Br8vYOGu6O2pbKqFewT9jurIZCH5QWujzyJhLo3iBc267vAB/SWbR2f/ZUPkeSH2jCFTiPob1S
f+XeBDhAs5vYzBznchfJ/KiZKUAtGp5sbSqvh50jH519GJwuN6dAl9mGq5+aplIDv9flYyPC0AYz
sTaDCcEqwXSnfw6xHeyknxpNmOgu5Z72ZQ1vZbWMHqIzzX4ZjXpZDOnfEb3dAZRdp7I9z4/r1nhB
xjyO/OIHRaljHockuH0H18EZ9e3Amuv3uHTM5I2WfGg0CdV+USPxvm8PpX0F/4B8LLN2+ylr1ApX
pKTrG/SWsEX67ZQB5Gzil8KJXcQU6KIf6aKgUeBffDoiFUP5G6/yBVTc4j5/VH1IvnhmwS0aHuUr
GYKqKv14P1+ZqOFnbK1NCrQpP3A88VeDrYZpaCuEEHx67/RleKidGY0a7jENpNIO7XH1AiptngpN
3IYtsIslVTxwm1CphfkjeE6EQeACz355nTQwc7ufoB64GA5x/EXwJJ9tXjWrkMTaKoifKzncMw8w
ex6Uym+g7Rq//arpmaza6EvvVup9Gr0COvVzXbtuSOZA0IVew6Q2tClJxUlLoVrKWJ2RM0xf0jga
un2fiCsiaYmrCGRKm49K5D2Dcd8Z4VU3h+z88K/jnx9RIhFzA4KbpB/oysR3+b211kkkdTyD4yjb
+X0P2K6k7OCZ5KmRTDU/Rlri8EwihH1B+GS/t9mcYFMkKGVVMkitvxTqSuTH74cUQC8PlR4Yo9MD
bHM/OFN6MbJnvE60RyAaH+PGERXidT7MhS1vrKyb0/NOWORYkLOj3BiwOMyKVd/sAIlN0EXAKqp9
21slqi1dbOR57PuqXf16AE8We5XC3X72Jo0VgO1TGhqP1YDMtQSPFSaIklvSpYJ3qhilDfgZgQfr
S/SwR/7lczrICNAvapeyGlAKCfHHkyE/VKm2yXFimwhgrllHpXpRls3snjMpn5gH7KLQ7aWwiOh7
arBde7bctnnzIh/Fw6WVi88Sg3QtBTBVrO31Z6qcERGy6QBRKK6jMou+H1G9EdFM/il1dPo9mm8d
nYUJYTeYB4mZEjmDdeSq6Dj2DwEM7uurslItTukSMQhF2NZR+4ZyXJonUwNUHBjaOGdsPsBKIzrU
SdkRJxK/qyeekvhcHvKJqQADhFFfuBkq34a9Mpqm8bZxLh7ktJrLupsTpcI0tn8JSWifKSS/b14W
qw7xsNuNgGacHAR7japsL2dslAvqhjqBPCQeUcRD94S/INwrF1LUIicv11V0CmsPGIflQQNKJmnX
ROyXAYjB2xQOCXnCh0lHU9Ka6I2Jw/JgcYWUNgWU7QceLThezv2QQrlxe+H/JwNYnwkM7ckuudJZ
ituEcHqkBdPBcy9BX6PB0bD9AsyKqT02nZySyGW3tYy6DbpNywEWc1xS5uC7dyUOzSW9Hli+4SMB
5gsMh0q2K/mnknq5LQ8F6zm6SG02v3OEVLLsNphWXelAEN7YuCZ+ZURMz9Mjzq+TTABCDYHCTCKK
np55Wwjm9uABkEwZ1IvoxFOYWa9MC17O9nAfIOvSfaaoWclwpgNDci2xFoad8ChoODQBid8e9wcD
mZNvLChZjDgjIwotB4bche17xfKMftXs5aasENG6KneEz7AbpKE5hR1d8ExDsL130LPzI+Pm52M5
VyLCcaFe2tRafISHMpsVz1Qae1PpMMLJbhHQDsPDjdxufcwwPKyRaMGhMI2btnjk7Qha84CR05D4
g/93YNzKKXEJFK69hS1+HxbiHqa5iHn52c46UzzzBXBarL11VdHMmzNFxiQKoCPnxrWCRUj2F7Dw
I9TP06b1VSpXHQA63frSY0GNelpR0MdafafHeyN2FVqn2pr049St1f3wkHCRUb9Lq8gHe6yDcTFY
M8vHSAIkr8MmcmLzHziFaV8omsk9lIFh5zJre3dJdvZg1EWCOVziEDoZTccl+Q1NyDQc/dHiPH/b
ftPR1kc9h8nqQ6txpHf1hTLrFbDipuZRXHPZYMPf73D+r7lqi2NVG3G1nm2sbIZghm+QfuHCJpCC
ufUaxh4SOYX5HwsxtYRAqKvvDaSWz1E00Y9XcB9Bx47XsWc7lm3uTgV+oRGGLHqYQ8IgbX/sOF7I
dgMPv0VSDGeGltNYkdD79reuRf2khv3GyNqG66fdmlzFRABh2qlRNT1CnG4hhaHexXWGEyI2/DTB
uhaEIdSxtR0DDUpi42xbIN77y+sOiGrR0cT67qNb4udLDzm1bkMQKlw9eYTPMIXLZ5X6rvBXPZvd
lO0YjIk8lm6c/tCJaYWQ2orsJa5IoFUYMGZM0ioFxGZ7i7Bfu3MUvSLt6OtMz20vECbxfFwFLx2+
PTl2sY6Vat1rojnQZJSU3PvVe6ekc31oWTi4mc8m0upkI9F7xxTEgyMTVELMNwH8AR3VABQa8UWJ
tmp2Dedfx97TybITF9NtY5ohU++ZxOTMu2TR6+APhRaIr42I2suNEgC4xewwgvD6uWMdrkJzaFil
G02QfkoC8PC55ELuNkpmYsX1BT+PZyNddLaoK36u8dtmR8Y44uJDWjuuPkrK9jxKxfEHzCu6PtuS
2hErAQh8FiEI1u3QLdi8Ufjv/pdqQqbDbiNyk60PgZN8IugG4misBxyAp5n4sfazgxgLF1MQ8XJs
oOix0nEWGvS1D569wwhgqlZVoL+Nu3OSCGjADUDTYZjquLC1seOoySxwGeVyVREfJjmq1RvRG6PU
9ng1WYQmE/8E4cG3V7hKEeV82vesWP2eV5RDUwrbOdmvf5ve/Yls7F2sDFRkdhHtdFTfj2kXG2dj
FH2pfu1uVdFwRqlujYix8TZq7+SsmdbbrwSkqn0Ywo3ZfpFzxuIWxMd+wjjCSdGacJKvTUBh78iO
YvSQxct0gneOkdQYEpiJgbV9psz/bUXuOVaPv7ZagUNC/WHF6nKXc1w1kf8RpI9LDjjw251DyXOh
tJhlYbLUYj6XgCm6CA5bIU/gFICOljOWUUJ0u+itBhgjiSEiTlxfUU4BNelZ2RBgonNW5fUwG5Mw
3Gmr23PAmUXJdxKjnliG9NhDu2s5eqJUKgxCvMMVE+16XUE4E5kWptnxkP3xp/z2PC/HGFU4v+w5
WCOFpPUceEu6JZq232hRUXMquZbbgqTuvOKcwmYAKcKbpQjadpfT1qvUPJURw7QzGC7l8YmzZDZr
DfTlZl0O3F5Q55grCwChxzbqG2TuKvCaOG9+tJQbZCW/MLEhzg5y/u7YgX7ayUoZgkaobZXVZH4C
PEUcrbMRmKh9GktkPCAx0ysspOvXqLOtUZMQNp3J72CUDGxeMzet2Mg4Wrt4LxHMLBNrw7K+GFK/
m/c+7F7CDSjCsxNNqBoCEqiODEXFKlY9GeoGGfUgijXTZ4EwhMWFpAYRSim9QGrIOg7wVkRfnkL6
JWSRgSM92yy1NCJidNylVLQZ0FnMUaYBUm3qLHoBoCQsJoEj0tTSO1VcKYphbuzp7sa4TPa6w0Ri
m4c8dsmA9jxOUeq+ikIcvHjDfYQFYksIRaj6FMANT8tM14JfqJydQEf5/Sa6T8fiH2IYttj9CLr/
wB2mFthNkaiCdW4dpMESoP2pPXb/g8LgESURpGUPMU0j4FkiVXD1L4GzNpdzWzlKui/5MdnnkAUS
i6UUxXY/pCkXlpV5a+AGVwf1sWndNFjKsbHPj2zUgWVBm7nniCkqJH5EfIVUCH9l0XPp7yK5L+6S
gJJZ2Eb767phtpbxRSp+zL99YXzKPTs0wbsAGnYsP6iT+zDqDZ72YtIPtPcTgLe5+jaZEcBdVy1y
gazYZdsjOhvfEMDNizuzkMd51nT5jfmYhftQsCzHBHyUEa4NNCzVZShZqYYf7qjaPXeBQoXOuXXH
l/oOS820bHW6dR/s8gNZw+fXc0fQ9WJmIQYrSuuVQgk+TEWQISifTet9RGKG2/tdGCXFS+aQMion
tT8JtWX6v0N3Sy0wmsTowTRRFGB8sqzlHFNGLMnkBfZg8OObQ7F9m80+WiLxpyZfRg0++Ezr4vZX
7kVf
`pragma protect end_protected
