// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WnIGOjAcHvI+6LyNPR75490wAAd5dfkTjKhsNL26FOUB7eevVW/hV27VM9fX
wLoraq5y+WnOJyH3exrv/bDo98iylMqt+RBw6hZ+MzR+Hjeaas4CyHsfgsa4
zhlo2q8TsAQ/gkRG+l+SD4CzsPfI95HQIK3/9TioEXwW4dQBcLL95Szsv1Jb
d4BbK48QWuQzCRcmA7H5hNkbzzQWkUCdOFGlpGIcaVudL3RiH2E4JYwGD2R9
ejE90T+Igdnj4DyWJYgig7IWLS86tBBlRjXNw5SwWWuFe6PvriDdX16AtIg7
eViekKSbx3pagud7N/1EaZinuWUdtzgVi59oQ37Ctw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kp7yjUf++rBejsX02YLxEIexBz0stI4eXmlowHVPc4R6KzaaZ0VeLJffoogs
+b8pHyJwavcPMLw4vcyaaDOB5Y9x1OtD0J0tGxAOhR3wVn3Yc94yvzFuB0ij
4tPNs+sPeI1hHKUuF2sv1E7yueVhUxtDJIzGQMz1EV4Oafd+oJo7k3Gn9dqk
HGqDus2S2ZXzcwkWwK/zcpbW39aMt/AOXJduwHH6l1/MsYd7y1v+YiJdK+Cx
ia+t46dLACnfu9DW5BN5mnefNEnJ38C2hC0Lm89dIzW327f8bW6rA9ALpLtG
kv0Nx6pD3LO+WdTLurMl1W3md7l6Vl5XlhQ5J+78hQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
P3JFT3jty6aMi3HQcaRMLfcXaCKpeip67Px+ELou58toqcrRlZ1IDLMYLxnW
AdvNWcQhYLFJS1ZJFxdpAYZ8aqrcwqbdgMD0pusungZdLhfX+99nJJ+yYML5
4lW25Hv4FH+Ng+UxUoo4w4W0othq3321ls7fZevf/BjpE2J+F7kql+qTXVXM
KlIutQ6AQB+6z4W/r0ewHw+6Cfj959SFSLpyld9E51KUESCDytCDpldj2T6E
ETLmAZLQFiYh/0OfFjFbsXxQ/kR03589ifQzbYCWmSiSiZFGLqNAmi5NnoTu
6wst8Z/d02/UlaEwQBIQAJaSshpj21DYS6LDmc2F9Q==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ogIYDf32PJXAo10nS2Zf4RmzZ2cIjEC0UVXhDideZplNI2Y3ATl1j6XJymt8
xp0Lsck1rWspS0vlDsu6apN8dIzMCQlsQyRZOsyJFWHOZXxlWgYqbBvTNKnz
5Tk7X/AGfH7v7PXEqwyaULaYkbw1UXx39cAVPMcaNRwPcFVOaz8=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
DuWs/P7cMjQGIR9PkGX5HBYaAxM4YQNpV/7zu82TSrVWN3WB0OYLY9lZvHfY
d7CRcx16i7XVR75ZESM+M0Qv756aTYxVj8XCGmUH/cUgMYL2tUWmklP5fWnY
IcftZMS8a6jxU9Vey71P8TGksxJUKVcL4ON2Caih6z4uwuqISsKkW0+FLDxA
Sn76K1qw9vCyLLqWmLPg1Vm0LlISd9WVyb7NcCGAOK9X9U085K30jqIxC5jw
PtzvKi1eT+ATIBNnh7QLfrTEOzGzJ0SP6LvfIyREgktbIOaUZz1krT2zoLZQ
3jL1DBlg2hU0DZfxKaCfvmxTlBo5lduwA47mrg98D4s1OaVwizzu0fHLQWiT
lpcoez4nAkNu1uAMtANk+NRFc2j1M7xHj6UdZ9eMzn0+hjvk2Xy4W9uIFTy7
oTfuBe+qG3i6cvFhRHg4ts4EEjbPkTqYUeGg30N35wJ3Q67Bg0WeTtXqu0GV
hkSZ6TvR8vntxbLvPTj9DuBcXBOcZ0IF


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
aZQF5MFLzwQXEi2YRmIczG8Kf5Uv446DaqI8zaxinuTPHJTdOGtMbOewv7cu
mpXxDGMWvZEwRvgbfPBIjCqX4mgXaclOJZ7ZTp4OSRt4BNKA4XANrUFfruf5
sYajn2fQCPu1B5u0yWgp53Ra9K7pqqchXZPzwoFpws8gbOXBbIc=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
tj2HN6r86n3zngTwco2q0YAL9kfJL/H/goEjPflA71x0yGgCTNn3kitLwUfc
JMxe6lBSNdqKMXCDQe3R4dZDt2mvM42PD+wcxlwYilINNTbB76QFYVRlR6+i
XrhohGr5FkCnvfsMKP4KXh70qCOJazVdhGGRTV/MHK/Kqx1lJOU=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 618960)
`pragma protect data_block
dEJBLBLWWryoLH2WRnzdDrUwQa27dBQYqf7KeqlI1zYmj0wRfthUkDW5Zfp1
zpBEYOJdbFaVKA14nuvqTy0EebuE4nI1CCI7fen35sFgkMKUbnzg+HcHDtQ+
kSy+bKdMg/CNBWU+Yqauxa5wAOWbcnzfnv1cnIzLGwpoHHVUAhf1jpYcutew
K+i6oPmx6pwvq6ksZZTw2TV71hh/gPVSWb7WnTwRUZKWyACCbhJfijBb7uWg
dkRurXeCdQJzeqcs9DR9hfVmv4+BMi5XLIQTx7Rp57W5sc/LP8wiGkNrDUo0
WaXlgyx5KySmT4IaAEFz7lt75tztOwyjxE9auVEJjTz4TC2cGxzulHT1WtCC
6L6H6B5iws/Y1dM7ptFw5giTj4Z+3mlNvGNMmdY8pGdChkQKlqtZkBcSJ786
VarwSUP2A1F50y+NTiklUnMNC4VTdZ2NXvXXOY+J2Dx6g9040aZK+4p2s4oI
P/RAT+FVLRURmIkrqm1WXnn94HmxVDgZnCpL0yoVpOLagtrGjh6nZpkXCcNi
k0fvAoF0i7U9qUwYb82ybw5h2N7O/DaQ7mHCORILOA8Dv9R3nqxsAb8FwqTC
KER/dcHDu+oQKRSZFaUpD/TO35erUsK4a5Q50i1ljIrFRxYYV+zkwuABF2wa
b2e1gm73m64alXxAMCwF4Qe9oqQPiS21l386vMUA7QYRjVlBlldvVJnMHRUK
1B3eSKMLGlDbavr/+CDqmIydRxyKcsCFFnO3TB0gEPEEw8W+L43mnC8q0CWr
2p1VYdOjmv1iRFrgX6Cs9OhdmhFCQppYLRFHQdruG9gBYQpDu5cLROBX6fbN
0ic0OXuprggUDE4x4nQ6Gqmj+LrSDdC1LevLn4wTwAp53Tc42LBL6+7UW5sP
iKwrDRH4yyFyVGeOJaQXye3DIpQXmX2/9P6yNrvD5jocZuGtb4XibV7JeAdO
wOf0E1S0xWvETwn46qNx9NdzDHvNyaqlMaQymUoSpj7xLukQk4nS5lqUOeR9
WLtFWjIwnzQjiKQ1lcVXQifQziaANWRo96B5dTdl4Qk3WCTyk5UD0Sr2sKPn
tve4sagoAfGZ34LwCrPPCXwgghG4R5k0KQlyJXnwgiBo6fsIaBlq41Xxmrmi
QTcNoSVrP2WeeUK+gJWm7Yex1d4m2Sy49n+dWJcv9kLJ+goAm7gaB7NccCzb
aUDo9pcJ7TbTYL51uQzCkTxSwagzSEccj8/Z9fqEC1+pz8TMV92YRP5D3uoO
AuKUakpNT//YOaVW1RMMgoO2kYjXb/B13rkftxZFKP/gMp6gbiIDDW4AJaJc
3ERnytJ+RUf1MK/qle2GOINYpv05iq7yRBbZWkrRb4HtHz1zo9lr/2fjCN5c
QPYxJpcqziWI9mPdSNdU8s+5ln40Men3l+/QSOHCJ5EqN2klcpzwnnna6lm5
vt2cTN4UnLNE9jZXx/vsqjcD0BgD0L8yzYsTLX2Azw99VR0Ru7Ly/mUYikQ0
yfHb/WivBQaEgTSCFLq+NX1hDDZLB8+WCOEaoPw1bBWbDr+d+2HTIGHGvdyO
c3ees+0xKldinP3vdVVTAOBL+VZlxEsvbYQq9f2POrCHhppP6JwPxAd5Znm+
yH4qy6v5htVqaXTd+RCBnQZSkCA0jmCjE0eJSQuHxo506x19QI7XSpdwRgV6
8B7UuyLB6i+o+AFCTYIs73OJPMXkyK+2BhuUrYtPqTGH264EnS4DaHK0anM3
e8wABrapi4RewDLyMzsroUy3YWmCMdwPTiWqvFIy+qw+JuLBhnI4j4NEyQRF
ThF6/PsnoVT6mdiApYJOVlCKxHmrh6JSZ3NAtXtCLBicWkktnH3aXEpTqdWA
62EWqMAnaaEH3H+5c1GHin+N1filxzK4EQ57etlfBRHcBtdxZiaFXx0WCzwt
79D29XPiyhvoDWPJyaU3yxMCd3NtmiVyPCyjts9TW2JCLw+TN03PLUgZBGqf
twKxLzPdHJkpdq2VsvEejFH5ZChOSkGIbgwR4mPBqh/ii3+XZ4fUMJ8jEFq0
qhTGlC/D76UFGFXX8d1zQ4oEWRIvQ91AG+qR71Ma/aKc+5Go7nrBAxdHgop3
kuMk+zbqXO+hiLbmKAyv4eD0E4uCP9fYhjhgYb+kkNQRerrvndSM1S0bRt6Q
1glzZuciQi96uu10b9JQpyGdXvfAfLEblaTm9WlXZ43m6C7pT/SBiH21H36Y
UHx4UrohiQKU7lPvFMMtrAIv/2gJQejn/RE7hql5hpboD2sWFP2U+HZYvj87
wZONB8SFuEu46rGwuguI07BziqrXc3lc+BI9IVQsEcwO2Z8WCqHZaM0IB03J
8MGd5qycErfDi3BIapo5scJ2g8Btgb4bmZkBXq8oLfLMoeiZXrfSf/8oCSKW
XM0cyySDdKa1T2ZoYmU26sGEpemUCDL41o+SmJxmP62tDpCfiT8PQZY7azSK
PezPyhF+ZK/7j835F+GsAUTUyULzsHt1CbnTXtru3OGWnr8kAuKEqfl7Ps6D
NK5L3eWTbBC5EZ6yIFfIH22RjETDZ5iIpr5fBzdYAXyrHtjlYi6t+KoK108e
iiH1Ly5RqOSRI8HHqduw73TSUImlgVDWXAF3P0943dfr7pImAgy4LFWXQD3X
20polh0ibR13UwKppLuKjPipGoNs1csJe7rK8NI7u9/GvLBEWMD4BzLBV1xZ
pyR/YEhLhIJlisk277ArgAh2owGrjWsF3dfEpv9VZ32aSkyGT97R5V6zu6J8
UG6Ofb4rrvG7Vpyv/CvlTM0tM6qlerCRbkgsZxiPrLyOHSChBiVkaIpqEDYu
eIcNlnb+V2r4rA3bNFfufVB4s8IxRHepUTcZeO3GAZBs3rmbdznVBEyr0WVy
pI0zC0bFVJ0r7TAQrj5LX4mppELQo57Q7ySI/KfgAx2xXi/zqs5W/XuYDirh
QJMwBme8nDJ6hJqBIXoZyinZDv0dl877yEylqysAEav/B2YNOnnpNSuxwhK8
Uy5MgVNdEZ3HYs2/dnNToXdEQf/Ih8VDEWm56qCTB5nzv909iJBY5bKIVqy9
Wq/+CC7L8nAp0hMzoNzQEhCuOfIMPg431zziJUjpEITtBlR3J4O1YOv7q4ZS
Rt/iUXYZjmOoo6nZyx2loCqzBSJIrO8FeasN7r1Q2h7scH7DL6BHfMFa5zW1
KfbmgF0v6nAz3eZ/srR0QysG2GJnZ0GBKOuN9RMV0bbO8UMyWu2DJRGmRhsy
D/P5m9u6ExDHYpVacftn4ySMaolvXte+Json4Qa91Dqk8m9mnVoZUEDJK4y7
L4JnTV4OheCfwfwiZjuOy5++AEATbnmqWVU80aCxYZSTnKdfyl6Aogg2gyiQ
IF618qkx2quc3mjmDGrG4Wyb5wtHImEGPb7NRGHbmaeHPNvJi9mZl6JsT4TD
Gi2r/t9QftzfZDLAikdPwntK4X9QMfLEdXHa10yv062/FkL83wVq5ZbsEHEj
8/03faMO59wx6eWdCFInipeAn33BFSqEp9I/3/qzS1UvlrNEoyFSOgJCNwEv
oiv0mLMKZAbsuCCFr7382bIGG3xsEbDbWvJiJJBzBGwjOJT/cDRB4BYpFWkM
0XtBXIi3+4/buSK61sPUH69fOmIqk/bXMUqMGxX7dAREb1s9L15PvXzvguvN
KYOxruIUhSZzpXqBp4nrS6WW+DXSB8wJvDC4cNTcsYSV8Pa2vyh255GDZ2Ax
DkCA/gKkxpkWwdHeJhRdY5zYp3mnmk8cJLvAAtUr/B8Xh9K4O8JBZrMhMbMa
XxwQiPtxgO/ksqYYJLEgCG0D1s3bDZJjt4MIcIlTWVpwLCFHsKD9GztLOYKl
0SYtMS7C5wTL18w8RRj3yFpmxnrsF4oCPq80vx76C7H+P4Db5W+cXflEnjqq
ymRAZgFLUXN7nBXo3gFI/SPJrRZVT5wzRz5s6UAyXGW6J+IPfemRbOY1l0XD
PAtbCGmcjW5FXc4Rn+g0D9Cwl8uZUsW7GSI/zKcPxxFccEjGpKCIAjBP47TV
lTI8BTABWIuiaR1Saz/ZJybFQQkw5NZ4hxWCL6EtURD5VMuMb6MuCMX1d/rX
r//bG6zgd5EBut7tdJPkb5x3wN4XCxCQbTeE3ABqm6wT0hug4NSfXLLXMWAM
puA4AE46uAAq/kZWzH9+AgIsMR4A9n2CQB94KZH8R0Ro1dx4KyCLQdzsuGhf
qlcytDjYL/3hgcTzfaaGuFQqKnm44Nv+hGxBL9ld+Fph0B9bMbIHjKCdJ/75
SMLKcf/zAmagQVS+OrvFAyi0gd2j6gUkdXcK2vhxus8s4ADbfBgBaTmM6ZH+
5Uz2SdeR2G9XKGrp5fxTfWXxcGZDDzCWpYlo8Dhvbkl/2g2MuYzDPxxGVcQ5
mz9KjTk7dFfbrWFex/1v01t3ZN1ztmBTuqgdElkf+GtopDvalFnz1U0X9StJ
9viX5v4ICX3ibKK8P4CD819034SHGZdZYN8Lwg6bjeHTBffeILcGZvBAq5Wo
VZdE/wvaMz9VhFeFrtm8XjFKeNtc2eI0vQnzxe+LVhj/XVuxevdz+oFxrBmK
TfdWqeZHc2wKkgmhN2WbGi4YflsLWxchx647kBu3Va/ZRwT0xCSfR9JqSRpe
XBLP5Xt5XKk2SnfGaTrGP37tCvG2hX4iDgqD8NhkG6kSIP5YUN4elQ7X8Ayw
xZsxAbc0FTOC1L6uRRgwuIit8qhPpPL2892DSj7yy/2qxhsq0/EpveJIEJqB
iAr+SKZuxXo+MzIchl+pS6qD3jcHyYkKeuAPD/tlaf+xEYjyfP27ssjJbWgb
2hhYJ3ftmaFLLnbOnsTmymKFsQuk0UzUauW0TVMLGsbLra1yZ6MLnbssQhkT
ssAaPgsyH3zpUXxs2cxlQJuT9UXC3LaIJdWY5jJ/wqgnPNm8JZxHosjRyfyg
e1WH6bY7ytXRtDqcARUEGI3TWpJ1rnnKV2gcq9S+8Hkxl/7J9awfWW5Nn5ei
ogTvAkeMA9KpJCLuWVoWiUs0aQBF/E0drUq7HC9QhCwQrvRsDHyuoO4P+anL
/8GDiPSKrs+7VXrtYxkgBPx6CtUencI7mpXavCC2IpXrFKdToDH8Aqu51bRW
SoAXK/2KOCddNc2YLsK7z98AAAWGpjneY/UYJB9Kl8P4LGWQVkm9oheqq3DT
fvsYuC7la4HAMBxb1gQwKXv5LTEAisX6nHkrwTK71A3RkQ1hgnIdzbGjNpxv
M9Y/Ag/OluvcaPLXXaTUZpzkcolZ0MDBRX0S7LwwaMt0YpzLu0SjX7c68erk
umSbsM1N0CNT0XOStP0orck3q7e+/X7Yyt0uK8CcRxwcH1X9h4mmWazgh/Kg
eLA19lC3qn28UrMoZ2LmCnhoVAxChh7NBq6re0h1j7hPpNhNnG/rv4LQqvpR
dQjnJxf21eQ//siSaf9BO7oR1ZsbVfF2G11x7oAvM44G+2Dc76DFxgYTA0C4
s0du2X9EsTDoCYDE8Zrw7pXG33IW2HtZRMIneIMncnWRtE40aD63a6XRPNmK
oyJfy0nAQ/cPUJ4jPONtLBgh6G1mbhfqMH9/O7zVn/iX6DtPDkARfBAa2mIR
pewkUE2v4I4wrM7MYQ3Q0220I+k+p3YYVOjPyhASRHpaM4ZNiMaOQ9spJ/qP
5HIUBN04pG1aWD3XmYs2m32DRoPMjQp6ytq0L6pbSswXUTwcR+8IuMey2I3X
iidM+hQdX99cHFQE/Kvlzgu50d04sbhIq7h+snJtY1+y3sn7VCDZXJI2fDHV
XRl4dOZGcNnigTzeCehAj8JuNHWx5Sg1AzIXtG6TvP2PFa7isqYS7jaFZlu7
HtFjIfCTP4Uk5G28+NPPxyU6eLAPD9Si431KBEdvG4Ug2/0/RuUVXOW8tl94
2yL04wpUce8qJuZnV5xFigY36ZtJLAnmLiE1h2folPt4/loewZZawfP1tL1m
zpYg8m1A6GsvF0iRCOteFiodyenZEpQ+ZFXMb3KMDyjpfSdlcKJ4FQ/1fIfj
6u7m3ZQS7SttwggcgurmkH49AeXbi8Ncb/CBIXBVXqvsy94laMvaarM//40B
1tccXum1G1b00vSCK+h5z/z68hk2f3YfAxEP4KuJotW7VyXCvxttI174jezr
C1UwhvK2i91qt9lgKYficFV0GQN5jxs88S3+abkanUyXQGR9ilLfoBy2WJ47
AqMZrvA9WJLZ7rjMnyPxJa10IDKUYIwbT1L3lXkbsutEFio1E5X/8+bxFKzh
rhAShnh9Bpa9DtIIsFLg0UDmf7pg28efmjTrdO+QnTI5pQwn+TcOGM18aymn
Bq201qYVLDwmBMM1emzhT6/1ZJ1s3BTTzONHuXhtEWwawrPtCustLY+0ID9Z
wGZFJSEYZ8dzuUZLF6Pdkd01NQLFSLXII8VsH62jwXreDkwyEn2dZbugi2Fg
XtwiHk5Xqjap+X1PEpj08MLAIjU7xoPZg5bOQBACAfqm3m3F8FVIy/OAyuo+
RnVamsL7sc9jpsdxd9onX0kuSnmSYA+3cWNhU/VpooZcZpRTiuj1KM0h2rs4
sRDB21SBIciruMCPEWs676LTuZsOw254PE+47Y1BnffUb4kzqNJ6bPg/RCic
F3hwbBlDgwgHretYraLmzKg3km8V/vs7zZ7BmfFQQTuZyylpaKsxzP56bwdj
idQb4veaDbBpI4I9U20qw4vEqckI9rOl1V2TogOAdxx7ZZ4pHTKjHUrkWYDQ
wPlBp/hR3Km+LD7+eHBnm4nnctsg8S75+XbSBQTJNH2MRyFkQF8hyPkvSNdY
2SwcxcYqcv6J2X/uFWiVqJDT0ME/75GS6vtvSySo+RwXiWCz524QZIISHu4y
7eCtNSCC7t6MQLEb3UYZVhxXjK8jJAKXA+qtv0heP+6IfLVUj1oWeUPCoKFx
EKx+eL+WALyiMxlGgQK1oFdx2VVWQINoT6F6SkbMMiZ2fqeAPu5aPCype4g9
DrfYRp3Sl3Gh8RRzVynqQ+ltlqhqSvd06qUrU5GjktycbUxC6mj6jyPprE7Z
p+OCTGsnsPyzOEvrRZdBAsdedBXymfzlQyDFNvqpSFomJiu2EMxfVA6HJWil
KPclviNKpiRnoMm5Qho45tuNQA/gIDbO8vWLgNoNZeG0hocNOeuW/DPFsm0J
dIVg/ThTEX0Tuuy6hvtY3ZSBhW8+L7ZLe26mCogMm+xsJXmQq7onMPPWb3Zx
KN4ghfDp1B/6lSYVn+eZFyQHDh0MmJ+tKfWfGljOJH8LlDIPjoK0PM1GuPid
PJYFwddLieID4U49kfbCUWLRLuywI3X8I6r1Ekm6KLsGXR/Kz4C4ezfutqR9
huOJ5CnhRH66H2cQSyqU0Ruk6qK/p8QcB+Go34LVNTlaowUwWEhlkMF+86Ka
fd9nOkp4APVGrQu9wlOD4APJlPFf+1+WaKwknsYrSxk9CaGepyvAFCN2qw1o
F2Xj8Qt6SrdDSnP/GDtOZWzCHIrTrXsgJzQL2vUdF8fjBcdQMGbhhKlU+Zhr
DJbkaCLb8idTyVdleS1L6j0zG5+pcUmVzwzozGxSRTHV9BC0Au5teMGP15Dk
NpaHzgd59ySfVJqV5v/i4u8giRlXPwdrIQz5E4OY9zse9EqWzDiWYvMzaq+q
3Z7+F0qa6dQ6MGokytKQv/3kVW7VVg+5ImgA3OLc3D9pVynrurRO5IoJeACF
GpCQlpKrBH85NW601B5S5w8NhX+1kHlXVmEQu3pUpTsYqslbf5Z2glUpFvSR
A4l8vlOj11mhMGNXAUNqSKtfM8amfmDCQ56XXkTqGwRMdyzbyCIZMFF3d024
NIT/zj2d/HAjchPcYo8/Gldc/qQI7Veo+IJJZFn2LecL867BXbDbIIfefyYf
RVVTwIn5S8CCYjLbNuwrTwuIzwb7QMIKdxM8DARC7uvQU8/RakjGSxLHjjdp
FfPR+E58yxnclKyFNdib/w8L+8lj07Q4a44XpqOuypgy8xtbmQ7TWlLYFule
zmO9WG+e3yj9ZgC6Yg6xWn1nNNR3/uFDzl9zD3fqZEBBNJaYgsmtUlJ0qz8t
+Pt7lpeJwJaUbf9+GEe7v8CEoIDscwapbNdSmAueRmv5gvtH0R81jEIvYgrH
nFXNFinBnMvfDIoGH5XEb8jDuPrVoLvT1KICN+sqNqAP23bx4My+al/0zIdC
tb14XOXhdghE+hYqgeLJFiFV90/6HQCybWHcUMlPqs4JmGtWVmKNWNxTybXD
qi5Ob5MAOfNf6lwZ5rFVFAG+M0xDGXGG0793f5+X3h+fW8CDvYLgMTNYO5wT
kORrXU0jo6Yq7EW6/2WnP6sun2rYT1u+V+eL06PvUynozBhd8CpvTfGIf55I
ylSveQQODhEI5PwVtqjBOSg7OWvDlauNJOWdHNkqcH4yOZ5lleYzrK/c4UbC
B+KFIuOcdnuBfz+RDSEyoZo3rit0lBNAiNPQreb+fJp1t90MlT0e8fXOqKfE
3s720Rk+MBZsgv4gOGW7icK2ovJ/o87Ut7jTnS8kPw43OQ1NBvlzaJ5NRdd8
H9D+2jDyl4A9hJcmOQ4jqu9qecqI66Q5NqFxelMiCK7MIkviRoSFfVqv+943
d///2jwn9tYWlur5pioUBhA9N2InMzPQeB35CFE1Z2mhN/f2ZA75hzoIk9lJ
w7r8AlHZb3wczmbaRmEFShUb5++bCpnLBYxOorDLuCvakDaXmBJpkpgprNRL
Pcn5tUTcPGK+2bwW1f6VopI/HOI2gTXZGlxzVYgHDABw7dWfurC8F3uSDfsX
NV0HvUafSdudHurjtkI+uHC8BHHDYyNDIPMaRRBLGnOrWhxTpVlh/TNQgiM5
r4jmEMgzu5UBwCpeRDT92jwNsPoe9Ia6nXL6m8voIPqD5Yw0GY8scf4de5L/
bE9JtQfgX7eOizT68XhUfmQQZvwO8b0VHy3CvLNfpPN/6DVyD6Otgkz2ngkb
aC/WoJYuETq2BWmKHxRlbcgWlqjKhj11y4BTceD2Gl6/0CwZZ1YYoYZgoPf4
XtDVpEfBycn6ZMLndfGkcTlsQUPQmBb+K9PfA/qGm+7xwq8dGqLAcUeqB0ER
xDGKkR5JkMCMelcIFfanw3QCrUpBriM7KmhKTGQjmuICaJMqvQlMTtH5kqkN
Vw6wDk92g3ybRQ4DrSyRjabNNHzpQHmGmUcG+zVgboyenYneFHJ0mUh8vmzz
ZmnV3y0esWPlabpk3Nv3uMBvNdQcDsAVwEth8LxYqiXir3Kp4AXYPHKPZqdz
kIWoTzMIQsxG2FLY+gRcBzrmjuKouUPORiYJYDyg9coDFi+9v0XW+yvz/Ym6
pny31TjxJF+2MXbdaNHumTykIdVl72HGKBIqiWfOV9OYY+R5GVpPCDW93u7o
hQNUQajMLHwNcIxKKtt2c4Tev2vZCQExWHO1pHme8OPNrUijNNaaBR96zCU7
c6AOTGb2Ocw9FNB9kFF12BGGb3/fnAWm6euYhdszy+kT+l8Hm8MLIMdg4e5r
d7NaReGjfPEPqJz16ig/Fayn7knBlpPIM6VNdPN49lIQpr2aXO+dKllu/Ti4
LuJoESLwL7ZTkkYt2epwXI8rcJrbDQIEKc6DoswvC5rnxxKvrIGZcn35N+Qi
i+IWxrzEyUiXXGdSStnlvttWAd28hqvjIqBPASMteJMIrqLGyjStr0Img+33
2kZtA8c7D4pjYfBiZDIr01fD9xM0jbuYLtQWSL7MWT3fZx91e9gYhrbDag5I
MsdDQgf6tyHE4nQ2gxLi9WRLXCeKYEGcUbbtWDoqP3nETfH1Ob2jB8Gbohq5
+QUViqAVfqzjNZ8W222B5dNYSnkK97PD3hl3GJ0KxG4qkPY30dYGDetE0I9h
dcqZWaAEOeBpWnGitz9Jt/DfENeoXOvxq3H3wa9IQgaPOgITgShtNCyGvQ6L
YcQ3hLwPbZuq+XWSiepnrgNoI5Jyu1zrYaY62d9sNUhmTmMPBaACz+G+1L5d
EQO+3A+xgH+qRmDopPcF9lXde+BLbnihTo/FVyr2xNuAfRb1YJNKqT1vDq5A
uw9Su8UIKncbV0COyfy7LlL7sZHrg1sLubdNv+sb8RtfDSLn8hXjMEDDDsP6
orXoWnInTPoEFxnsqOK8EWenayRrZA0abJPQCP+MzmzZ6AFxDtG/qYLrHpww
/5j1uCWmqpoKGUqBMZE7EgjUDplrimwPNiNLzKcoVmhvd1psvJD13AJH3ULP
7L2DmHMWNbFqoKrYJ6iycXmFoJklLiR8CHjukE/aO4lvFKpinKOhwHYS8i+s
iSh0zBqEw1zDY94557iMvqQRMGOAp47exhLKGGYROnJgiJzSsgqO9Ml8TnGa
WKpJjEmkXlipuqDRiP/jVvKETXOkga7zAOKwsVXRlnNBIrzsMP6ETKofyALG
sfM1NRhrW4DWWwXlpTwquTNfr+Sr5NDW7AQXZDLaNRuQ2Ba+7CIlCtGB8WS/
o5xTLMORJ+PDXTliVMNFdYh7/rTz+aEdzslaBfTxiDXj+QJJPrk7fx+JYxnJ
sIarS7FkHxnvud5ZDfU8h06uVvC07jpvCP2rES6H8QK35zGjlHfEZS38dfuQ
2nar+hbL3S9KShFdKEniLfxXQ7BUT/NozgtmItLgOPWl1HpCLE3W7n3dzDZy
JssrGDS6yVfHfD3CdNq3FE+c2fvIIWA+jX//6ZAFFXm6/y/OIkAHJyILkAdJ
uUAdSms21jn4RlCjnR83s0rLSmAaSLfqRqvB9ixTnmwnbYBxfQ+KTcuB9kmn
qIFmDNJNJPiAlUKzfh1Rz4RtPtIZBQHC/Eria+RTE66uqCNAj3CcUxuC47fH
zTX7YTdxuwvwyP3HMMZWaoXM+vOOATU1WG2SW7YNcHBvvvsqU21FkyivZOqf
5QbJJCHJZ4M5jxSJNGVoObcl3GT6BdJ80Iu4DqwArha46HhG4ox0WvEQaFhe
Ite1hHm996qEtmHaOmp/mIjFLpnDUi01jjWOV6yGzvudnpjI9EpDIObGyOfX
jNz6hcJ+uBMCIIaf5UCaKJ7zcCUuwlB4d0SyiLVn4yJ57HOHaB5Go5ZAjZJE
HWlXEbjR9Xp8cPMDaCwQ1zPFZVkJTNYX6QzKbhj8Svedcrq4TGjA1QYnnui0
kT4Kdqb7+tkv7e+NODECH+UXguaqKjn7pJlZpw05x336YcyaSz6cSKVZMwAB
hMe2rNUNLHDftEmjQJZ8N0lNd570luINf6rKi9R7pL3HRCKMvEceANmz2wHC
4Ew9ilc7zsO4Xj/xkbErLUDRnP5yQSD9E3A/iv2kUVAgeMjZ1XJvgMVMCPoX
7lqEh1D1F9roMZZnXTgrmA6B6ovN6zzH6jGE7/VjyfW2OqZbH8nIdxEvkl3o
SA66wKjsvuYG6ZxjCu8m3nK774W3ShBWdaonq/uk6+TDDDGt+GwloH7xPNXq
ukTVdfnVywSncmf/1wLtgh/g3wMKSrd5xy9hqKqrB2PcxprmUTxCt1DSqtMY
3xKlHYj7ANGYjSfF+FpJwbnF6k4KXJ/JtO1WWl2a6cem5tT9tN73vtuM0/l7
yd761mbOopuUCzzBzN1wfT7HYpyrxR8yGdiopL2GnmhpQkOOD5bnavoYJVF6
r5PYO2gbeljG/0rEyojfU6LiuKoJe+ldgfoVVN4eHUKVlS2iq4Sw+lre2C3s
XMx+i5rGZ5DZcGRvq7lO1TnWT1jj2Q6DASJMGdVyyX6e0wuCw7nB7bI9y4dO
UEybE9ud52iSwuqDHwhnrL8vG4bcTCPsXDEdH/MSmNDhldRJ1rnD44s807cU
M4mEyI4tY8pZMHnM/+rCWXUEt7sEPyZfvlZcsmaA1W7tVtSBqka/vGvdN811
lPvE2CjDKKXGLrnJIU41wwhxF8nUlGd32tlD9kWD4v5uUK5uHW8zDRwOEDHQ
m+B99dhZD88Wtn8QbXCByx3RaHAZI3dpmjHhTYsHCuYezq+7k7Lkpke+xFJV
YhVNdn/H58d+LRS34GXeGkDMuASp1TZu+KFy9gzv4MLLlokoligngpI+4wyL
lTZlAEZmmTNBmwtefUz9a9aY5LCKuDL4ZcoyI4QQKQuGacGWQftLAPGRHscX
dQgXphk9PcHQ5WS7IVc4DXgsI6+phpOPzytWtK8zzeNSg6QPWIxpfFgulnPD
tikqrOrjsKIL7//OJCu1DRe+QadSJ9F4JEHp5zKPLW9g7QITPAmcX80FFpun
1R+G5f1BzUZpQgZZHgrntogBVTL5H5dyhbJzeKFOdvVx2qqI/qTjJc5YV2Jm
iYjujAr1SiJDhB95aHFhVdko+hWvNpXgPuFEJtEd0I7FOfSCJPYcT//fsBq5
3dteGTU87pCMIzLP8JxaFmww+tXRpVE3c+4W8wLzbFm3xf05XHvfCJqLLe8W
Tn6e4fKO+Bcv/v2kQCzf52kFYpZZMWMTc/WhFt/0EErvpyES2lwQ4pJTr3P/
032IOAh6HLYg1s6OarWycCxaUYPKs+Jzq2Hw3O9lS+55XzllOWWQ5g0p71U5
U7NFwBPEjkZ2yFAx+jIdSNN+PAjxXAjP1g9G/DPwnFq9N1f7qfxWtyKkTEEK
mD1MUtXK7WSJgYfiEhXSu7+larrzLub6JBRkd2pQ4kPqi6X9SVwcXBmyCLS8
PsPo90G74gD7bQjLweiAkdXCIijh6kvhhcEQiITuhooxEdJQKi1XoX9N9wip
WEvMTkV2nj3sdjv92AiCR0zl+y+SMb+dVGI3Vm8P4g0LwGyYpKkwwGmv8zir
gynLnBhWE2RQo+BkosoSQmyU8eB0H1FJi8fUUQXlL9uLT0LISepja7N/c3WD
o4DHrhe0U+iyjUgqc7xBR01sk/wjWNUB1XIyvX+uEJVHsVUS5pHAKHgOZNuM
yiysQd3++0bxu79O6muMApe3YV/SlsPPysj5I2KrSIpAljO8Yj11eLUlBM73
0bwWUpLrF0rAO7ha/9EcyarU39gtSLLdX+cjgvpxcFQOcZ7/rcCRoppsOkSo
gGFrT02TucOO3MwHiVkMG7wMFBUqbiJCK0gETdPJs5Qy2AbEla1yWeTJkSUz
zaorzSJvgU4WiRfgM0aVaErjfbnCEatYXsgyuyWCFU+RENjnvzHpSZQvfyHd
hq0q36Ny0ly4CXRTM45n5XfDEODy0k7ge3AYdMdeP/koqdeAMO01PkJgi37E
DGtpr5zW3LJSZB7OlzBeADD/3R4nxhs6WWoYclORWm3iBNK6v4CsHDT58WN5
+KLfLtvFTM9pikVoEkYnIHfb8k2oL85QuRNBgfKmmaLV5XlAnyt/zITtJU9L
DUa6nRBjVnCU0d56t3T0M3zcm/UAjvj//DmMJurVoa9QhuS1iKaf1aIBPB8F
SNWagEG69WUf4NY1riqi5/fkfzq5RAGQaxeRzaiHgTKmVNix/9tXp1pHvqAz
Y/S7JFYpP4MP2AXa+UivPVdakOVeD6i0gNosZF7OXUZQK0EU6AY5xHxItxx9
gTyYT0obNmxFoGLC+RXnLwXh6skbbDv2wfsG1rxeG+gkgrVujW4c5S1prJM6
nPO5Vd1r51zSpuHjPn+sb69lv0B7uvOC+g38v190iPzHU5B4QJGrWZfPBLMs
kwxYv2EUbpgIPGBYvj3f/HGGGGeeKI7Mgjq0HYDpx1saYxyLTjk/EIv+mCWp
hsoYtXemlcz304+9Gs+aWQWofet3ddcv90NH/v4UGsns1SwXCgOkUQGN1z9O
9HTCvb88GwRCPCOdSgeY+5AAV1waaVo7+igtkq5U0KSKugk+uKayukuy1/Gk
4s2B3l0juJkIgMPeuUvo2uvhrgdf9B4ZeqT1uszIO4Uz/DbLE1V0tg8g1n+g
rIitbAeTYRQKctAs9LljufegjDI5PVXkfej6nD/xLt7C1/sjYvl86rmG4RxR
43UIb1uh5zcabq4TqSJCnEMUIBf0oQI2YVV9RALcCAtmjuZcTyQn9ckCSbIH
eLQpNIkRNpnXNvCizVx1pdLnDSqdIkYKe9/i84eG2Ij7jg4ux8Yeq87WPeaP
sB5jduqillI8qrZPrPZXOnwuyQmDXHLm7jpWN64UktaF0y9bbZcnZRhWtAhr
Ir31g3jBGBXApxVphX6DihJaVRyh5A6YVBgxy9oD51LjRztjY2abNQKzsHw6
OyUBSqqF4XVT59Lej4pqD2OwaAylttzTIwcT1VxaC9tWgZcpA9B1pdN8qiO8
dJX9IK7racUkkPaksFBAQCmzS9C1y/zOmYjYib3AAvd2XuMr7P45h6P7JLy+
HM3tEiF2TffEpImfdioAs6CktqDFfSvPbZaSutBtM/Z3UJZz95JsCVgXqDvB
OF4c65ny2Wx2noOvhgf6TItpkYy5YpprXFSN5S5xZq3aM2VmsXmB+wwy8Kfm
31SqfxpVVc8PurcM2iCQiSNtxsYGQ55rRc3c6lIRO7WyhgXAuV9t/hXpgvlt
P0JJ05/fexNwwjMDa2L1nNZPgHbnFTrsLC3ogQhhaFt3648ZTZFZ+neR/gQz
DXSZRNcjgNbiCNMXBrQQprmlNF9M9u4bAGQ1Ce5X/rIQool4Rgtb1CVDRc2o
NSVKGZA3MsB9zvJfSFIEkeuAYyPA5NvVyVkJvJyypGyGmwomMqh4RXoOtLr0
zpNOV8K7jJRFZ7Sp07Wb4rJ7cnyyq2jbwkkPU7GqZYRnx4fUwp+Gz+W9cYNL
YvYfn9QHmRYkDgckIBFa5mX+q3CDHFafVVa1MKZsf5fG0Ub0vQLtVh1hrzDD
VxTFhvDTqOKNOfEp/3ebvLfNu7an0PhzQHzkxtqeS2Fxb/MpTPZvnxrD4yfn
YwMOz33zE10vkf7zOGABk7EoNC1Y8beeSjPlbFWs/AJtH1zYd2F+zeRqjrYp
+mDijdi7/6L/eLXVqM0npwlYD84b+rde2y4ardIzJy5AiTZWanvf7CDVrFRa
Tpz4U/4rLrIDEb1BT4eKCTKiQgQxtcdAcCmiC6++nsqtYW7xzaxNL21Mr6Yt
44AvlTnUXF5atX5nFZXiPNBGok77yxZ8C580/4FKGsPXjdOh3cXbireIy2fO
ZIslJ7Z1aQU9px4hvA9CuaStQIiqj+VsZmx7oAqOvpkatUMJOSb07faLvdnX
QmcrRvcne2ypyFd1uUxUOJ0bhHjLTSGIHO8tTr3+78LlLyPdEaokPnxGh6ie
5meu4pMYQbnHTKK/BSaTydd96odxo0c8lbbzDGphpTu0pb3R0fPAscerQDy6
uTan52TJiGOn6db8hEB0Hom5lfPYnjCl0OiVucFMe8MhZ1TB7MjF+L4EdowY
MQ6MgaT60kOosoYhGC0N4zyQXZ7xUfy3C5xjjJ32MYx5gI3CNGL0OQcwg9h4
b472FXB0ciIRsHtNJK3T8eWPsAAmytLpfzCE5aRk1ZdZ0y+jNt6R9nniHzFj
gNIUkOlZ3hpOzPFDJUoRvgEwdjXgCmsC83NbmIKw9OLq3tdzrPFXdo7Q8DKi
FR1QOrVjIGgnA/4FC4QBPG6MoHqWPOLWIV5Knj/DyJSSM8XwV7QA36p3qfxq
HWRnFevowU+DgyDQMoNI6hJNoV1piIW+YlG6UOmjW3JP3aWemNbfglgD6j4y
jsovgAVQu1u8FVPLdsHVJ3ralzT5kdXZB3icd5NApB6bcHMufRbhTu9/qqiS
R+jfT2gK922XrBijT1UHJH0hhfgdRNeuoIFaBZFgRWUfB+aUiv5z1eID0McG
Rt8wD2AxbvOcaQc7NRohkzvATBzixKYUkQGFPGHcDC1Z413Zzx910/GIwHvs
zF0S5o63yPpfVV42S/tj5aV1RsfZmdkct2aDmhSXfLLpzS1FTzkSDnAq+qdB
A3gwHc0XdyiFeIEHJ/dzkT4TlZeAm+tHE5NRbT3JPssbRCUZCX7FOa9ASvbC
+hOW56UBJ3PDOQQHITPkDVOFHoT+rLa5zDDuvkKkRXj52/4kOaWOmA7B9OLC
tpOpdHVCUV1+G+4HQWbj/QypSzSqTRwXAba2h4hP8q/Oc6wsLEmrNdvSilk/
8gGL9yM8+8z7cpOe8Fo/mBKn8u9N913T8GYkEnJ70zqz76A+nRj9CN6X/KCw
l256qnMih2RlBHhel4BiEZCAyZcWFujTsXylS/8lLorOF57tZjneoQFv02g1
vyhcQfTSM9er6zbHBpCXqQWXTHAbZV25rHgkqPnhtO+yvlaSTCWumZFh2dcx
JVgYzgWsmocMSTRnk5hJd3wCnHVtahcGhYXj2wY0n6Y0nTmKt39vVgBFKvFH
FN0Hy+DFagCF+KK7J1VfOScE5sXtrpL0EwmNB/RhVcT+CCu56h1nCYyeHypW
R+P3q4RdJuJOjBYwRLDzmfzBM8idyyae7NTWC8sIg6S/6iWQT32eX1Qivctm
X/s2/ZcyxcSIIXi4AjgnGXuDdWrvfZXB9IZ3srN0i5fZeXrcril5RKb1LRyR
yIz2Bch2wYsm2+xan0fjjydohvPjRYhWQZ9886FSefAG40imt5dpQdg8Fk4h
3zgcB+eZ7cnEOzxGRhdxG14+WqX2tlawJdy7IpYd5QdK5II2konq9gbVYfMV
3+wh/WfGcrjnZfZAq9Vc7jfg7nY9Tvq0wcJWMJUshpIdrT3qQBN2nfejNUw2
sWhdQjqpmvvxVFo9oGl61TcORir8de4gRcTNCq7wVvMA0vM6+/8h9wh25p70
JZNQDuoaGIMAEU2rlMbi7Z23h3SvseGRjtlr8/c6/P1d/sHyqDMsnTRFAR9f
VLFaV17PopwQkJhMySh6t9lpNsGjt9j5fQDRpbN+72W/OQTmldFeGlUPt2Xt
Uf5U5C0LrfvISBvjBh92JgZVq1JoqVRLXhopHuW2hevQTELH4vV09kx2rEJq
Jve9dFH9wUYKzAZkz2erGEbuT+i/JhsDznaY80IG+e4zziKho6Ie7EGVKh1C
H07d+4g7tvE1jPJGraL+miX38S+kfHoSvtzTYLJZMPGl6NG+D+MCRWMiNsNT
cVdFxt6UkBZe+bPpJPxP9o9m5xD8a7YJvpPFcqy1ugFevcbwpEvunJVvnQG1
flCNecimeLLrNf9c1h9/onpvc+b/gjSq0KSyc88JSbVEZi2cN49DE2D2ZkVS
wap21+43bs0w4ou49qiZZzdiD/q+v/FG3joIE7jk0wCFHtY38zznhd3oJj3T
PZbddpwMEJ0YV7c/q3De1dEJ6cQo2jKWViVtYRmxjdQFt4VTIxYDQt/qwu1+
aP3sgx+cxC9UwX/Od8QX9E46rzKBl9lmqp20R311R5eOD67BVBpSgkQfa5y5
XfCxOCctubtTCP+1UPyO/cOq9odTkNvL8FYGYcUREv5Clo2Mwf7jNVFcFLr3
dv0zAYLY54F/W0CxUOwgs+ga+0dcyWzq7ni4EXqgbnIHj9NKnOCdpYesOf3G
wr5/T6LUSZqi6CPwIndMLOQv9zYj1YaSOxwnc2yuiNiunL8dfUPedZlMXMY4
ywzbN7dvALnJ1xu7kJN+GUTZlZ9u4T2BZyhJV1Zr1d6P92O1SFkvWmORVT1E
jRD+ukgw6p3L6ZyBNC9N0vMQkvZbuZxJ8hbUJr+qFtOqvzU+xlAHmjO+yS8t
GZYm1kwgIlmztdDIkODjHwvGbY4hI93CinoMJtjDwojjOU2dQziFyatxkN8F
erpvy/9ZbMxgt+nUVkSHzsjDmPIB8knznP7k7NuAyLkBNDfrpJRpj3GYO6bP
4WIdfEyttDgm4s0pLudESZ2FPBtdD5YO/kSfUzyAAOIkjjcN2SGJRZ1z6jrt
2Mysivy9IK+126M3Vu7lus5xLgQ2rWU8Hd3HR5vGxA8GEosEwOa8eE335e2Y
yH2cbvNsZgHcuRp4p73xRiHM318n6EUPwYsLIi1Iq3j9cV9/e2lzFSDGcMjX
huft+cjuSVNMvBTmtaA9+yE9bGtlyPoVkQzHX3I+5kGFB5MDkGJgGKkM8Cbr
gFHSS53F/QsDZ2uF58F9mP/pD0klkW5/7zRcQQTFbx4Eh0/dD+IqGobGi7QB
ZeqUE0MnD+GNMhXYluiiFig6NEB+kertY9N8GCkp+uh5e6hgNjBpl2uPNUPT
sADZ6RxesQQwM3+ijPu1QWt4wlfOFrJqdlF1RCELgWp8GQaRKdpqcrwSYxGA
sp/9xXYVUnlWLdNRm7++qSMRQxbuv92f8V2xm00oryfawZjx7A3UcW3ba5Vt
1hV1bfmV44DJQYFPK2EGvZU1M8yxRs86gXBdx0DBRc0fjtwJG1hwJRy3LBC1
FgZp97FSarBFZ4aAyDnIiLqsqdnPQ4aCATtJ8nR/ypKgq6gmYxvizDTHYnwk
Dt/VuEvAmvz1VffMUjfR69HXFT2tiHOcdFc0bsWdaebaBMsgPxkTQXp40d+Y
DB6r+aqPhYsaAcWo4Rvm/M2XJM1rbq2/RzwMm3/QqF2ZxKVIbBWJtWkUHzaD
jdXtc3dKM8jfLkZs9K0vumINdWgeZhqCAglhhscC4vEj+Wvhk29Sc14yVwjf
GSr7rCZOIwmABzJqC/+UOOC8V1bB4ZE1GU3WUe+uj1FXE0GMeLxZ3FP0uq6W
zgn82+UhQ6Jr7D30BPgDFXNdrwR1II8Gg1V70waSlMxbjt25In6wvD1Cdi0J
5pDrvTj0xktUeLIc5aoYSWeQ3t396ox2T/iv2quB8ZFL0KbDUoHS85c9j4TA
IprJrm21aauig/O3NtdNGZyB75K/CFPWXThKkzAcUeBa5TvFsSZhxu+CGpd7
hqmBmlYkpvMOkCSlQWTC8BB3hMdS62vMFor7PYOEUPRxQ+Vxkeq7RnG3/s3o
q0B1HLWqkWROM06704aZSixJyqitB4SNdt9EphQTpxPBxdZJm2LWNQSobkih
TErhEWJKc4gVx7YBXk7wT5pewWyCY14Ii/x6RdqkiR/2F58KGy0ubuZjzUPv
TBPrJGMW9zNb057Ardt+/qbe4T7mx8s4C7ZRR7Wjm2NZ1eyQiP/X11+v46Aa
70obf76/qjXUUvHyMjnoIO+KcKPMME6LnAwkJl61VskIZjTLR17nOdN/lnvX
2OzaSXVlqJZogk1Iv5n38G7F3N7tLSzSip0ie/fHamM9wpYc6u9GuIJPflN9
8yqK1OUwJeI2gcCrLMWdd/mKSs6UkwIV5eXCrJTgWqGiS94c+Il0tucSX/VL
3JgaNhGT5+EuWJQNGMA+KyOT6RrdRLy6gK4KCsdtCcjvczrIhMnugDJmJxZP
6J1diej6M8Dg+UDm+6m+HcKgxrXAernXqAF+uTEBo5LoGLemcLeJNPySNFhS
aPfbcn4ktTc/M0TmBFR0kPY+2EFRFWUMuTbeCvqV4Pg6sbR4IC77MviQlCt7
N+rTqiJcglKVHPDwLt//tA8lmoiQFt6wASfsm7ntSjSFTTaokY4LmmBk9/AM
4V2fnfy8sel1FmBfSqtbeDCu02uOlAZRe2Rithy9Lml5HOlIsO2b1sX6KEla
8Sau7JGWxuUvmOPI+wJsefxSZm5ezSSST2SuVM8rMbV1duHCMZ6IqLHX5o+e
NGlmuJ9XUhnFnY7Hp3DqyKj+Xxqmij1sBbXzDYeQ3s4qNhW5s9legbL7TihV
nEeTjOhpOq41C/SAZ12QLrTlRg86UtLeEBY7bWVpHMyRi+DbqQoqWIK6aP1R
4X4c35dnf3ZxcTMX7TNlZJlTcGhgrsIcv33sSBajmQFvo40ecb8EEDpN0rJ6
F9D4p8l7+bC9wr/CZwtFVYL8gt9A7+xJPxhPSYDkr2uBqQp7UoYB09dTYJ8Y
Iod1f3Yd2X/i0euJ/ABiQxkoIp0Zoc9MDYXpNM4PS1wbYphccjZv/WvetwEK
lXRDa/pHvMADTNTYADaGvtekdp3uxFsNt1yAWVg1vhSOiRAGSuRhegp9zi4t
mgaaevXODqiPMGfDB3IfvDE1Uq8qJNMaFhzw3lCl7IUptIvnbgALhmYZSGXD
brGODzsZPrYL+uulCMGWz9SGZ68o9V2f1hIrcAcDZmO2IspYkkeMcRQ71Xz8
fB0MepfOmbBkQe/9AE0XhaQ7tyVcPKtN5F+xgOHfNAJROeZretFQNwcf0fXt
BuHCSWWQXjma0H5Br0vpvEbknYsEM13agquLQiXFgqf3boPXoheOnd2PFOE6
IA6OGh6VgYhG6UWdIW1cV6YHwJdNA7fNZJqjmoZ72l6/iQf1eCKNoZFH5lQR
mtONwePta33McFrZvVAH2Onk3CCTT4sblZHU6+e6rQj+KyUXJwSNy9S2O0mk
DeBi2otRgvGh9hSO+yOimz8Yh1sME0L2Id/vTgik7jdWWWp3MiSFWSUTk77p
0LWeUqjDFdY00MGmYIsdsqAP0+obZgLWlHGv2hi9GCoQRcox7knAlHIKQXoC
NhCxEjN+zuh9dHg1GiUkVGJmyBSQIH58NqJ5VRG9qHavGNHo10UpVBlGvI0/
tVyLWYdSHmAf8bnznVV0gwx36fZJQQX4TeXHI4CM7F/fAxXBkEyabsS+A5o7
gnuFD5w7kR3cvnOQAtTBmcLTaEjlXD5i06wwTViVWlIja3YyaUrtkg1U/3yi
c66Dg6cP14+Zf2jEbTnuA4s95vfD2Xf10gHhH4gH4jhwYHWfQ4RFpRGue+L1
q1CjutIw+6I063JUl2z3Nm5R4qe6x06JS5JD7eajo6u/0/yWpczTdcLX5/KF
VFuqsArRP0BIqKiTGGN++0H3ch3Ku3TYUvqngoDd4Kfr8F88ZASv45SUII7o
H0dB98GX+QZh1BE1YkcO0QqpHAEqG1t+TFLk0TJVdkWTF50QKHLwWXvmbJ38
uZOsMvatY+AA1nvl6RKLh67LT+NQNlar7D+AoFb5anhEMHh/WKcpEan+KN0M
nigCR9W05J/PdzNgymaHkpVCqhd93bECg4NQ3GGxjOKX3I1EfVVXlcmWtRRz
yiJHi6/Tj9wGV06ezzVoCKoKThr2NXzv8iHFXO39UTyK+m4d7TTGKJVfWjVx
iPwiXYnCUiDXmsVm8Q1YG4r7dcMOYcUpvKfEeewFjYrkSr/4mXoZ8hUri7pi
JKxtBFCCvIwcJDv3DR/sTpUs11CRgJ9uUzLIomr0clGfXnSZRdnpyhKZzL43
n7Je+/i55x1jkd04GkTz/N99gbixY+3WnymMYqwu1w2DByQXfc5IGzNeeWQL
SZtxLleAYNXHhVDhJwb8waEilqmAY+tc6V35ZHRjb2v8SPaxum8e1+EP/SdF
26x8XAsgX92fFq9o7U4oys19VUH8BlBWvdWVAdCitBJqlmXTui/Y4c6LBFkf
vRu/SazvOoOaglvZil8Lu27INbcWA2cqSKqSSWXHWjGNv+CZBr/O6B/ry08i
R7Ri3n7Usnx49ADZOwbat1XM2rDtjgILO8E+NCQDYCODLhiYI1+2D/P2WNrh
ay5/Qf7Kb86eHEJfmb3k7k2X9MPX3IA/Dag2r+zB7u3UzDtHlT2JykqYwPID
stGhsH1eUufJzLARNYBr/NsHOs1D1Z7o4aVN5n6cmPx0L4sUEnwFsgPwqgd8
Qhn9Zn/TDLCdE/msRVx5ijz8CG6X3+cbDXHRGd7sJ6db5nMm4AMwqnhthnKt
8LsMJOLW2C7FiWX66lI5rcJqhExu7vaCNredGLGr3gTCkknxHfXcxDmeOn7n
UmA7a0/mQpn4lfkDan/qLT2JTlefb/ybYsiFvDanxLfPTeCh32aVvQvL3axq
qNPCiW8BBpKwm1zEnX5TcwdlpUbpR3iNsNn896LDzXKaKHUGWKS0PAAICVAV
LV2CTfs6KsbAxTHQDw8QxtvcY3u6ywxQqzw6z9jSaoucIaHwStKEZ96vojR1
S0fYz5iN8W4Va4D9iyrb5BucXAMFJYWLe+PIOoIRy+Nh0PrmALXA7cwiaGOS
Yb1/P6MiXyPVAEVN5xz5r6gIHDgJe3tswV7W77+FVK0dm5Pxvwx1Ux0tN54t
ADkjvPMlFTcIVrsllmZd7ljZ2QQnDqMBdSfC/QiQFYSYrc5n8uV27JGkoV9+
7YIOVyDyQ49ag1QRpTBksN03PusjRK7LaQjs7AsvKH9aZqQQZqjl6HIslk7m
GY+yJlAxlWkPoH/E++/Igtf9B+lgnhAOl0lkt+eW3U/5yhAti39daUm6DKVr
rRqIB9iiXSXWRLM8V5pzpB/SmmnUlqAhFDhUmfbS7pKmAkdY49A9vCGgWRVu
DtpNAk5wxHr0TYr3V2tIkXpBm3XVvIM6m5aKWyWRt3umgPq22vFPop+Cu2no
On9IbuBNhEM4DMhedIDvwITCo4fkrDB4Nwzfh2KZ/9I9IJb025yf3hbeadlu
KpkldN356wqyij7Fmr3hrE5RkJAB4h/oQJyHbNFOJCqWa9ENSSKAW2g85aqn
K5oDOOSzYvLqwhraLn09JGY3wvM/Na/SPw3slGJEA9FWsB3q7vWgJdZIZaZV
9b495DJP940Codf1RdS8Sl6sPws/9OA9c/yjzp8Xm2LKeXd5uO4CoCnMbDgV
9q8dcZ2VSNlmWFFF81KmNSMw96neWf3Jpc3bbHlbsW2zN9t1WbVybfPB0rw0
etWm32bFE/JyS2ElNc+jqQ/qFDZ0J83BX3vvHG7DSsBlKlo+gWbJEzMWffOr
nFwORRWri5rElBz+GS9EtWTFIOqTOatrZ5DnC32w6qVbfvHT8OqssunoktWD
DkDXpJ6dU4ngWB6HjU46RpdNJNPnVzYczK0tNWrocleN/PLVWJD8Fe3JT2ug
a9Owv5Tml4JvD4zGF+jMICVTjxkUoY7s+YCgRC1c3x2kYUB6bqgKJ7azEIAh
AlG671kriJzsu/CyxSVoqy65ke/ESJcSaD0cz1btpqE73BgGPn5HUIQGK/7T
FPmDiSJDLv3yM5YuDdXGndSow1Hj1mC2zp5xv1qkXErbzSwY4eXTmQN6cKdx
EiK74hk1e4lncrMhagzFdIJXTTJNQirgJQ2tUHSL3tniDHe9g69CjMkJ/kz4
zFpzoaT/q3Pj/K0FP0XI10dSDSbIILRD/Q/2eiZnQnXHfnzIgrZEkoRvqNJN
pvBLp9BSMQIgkOVozbu2ViDBLPfNt0ejO+zGQ5jOZRZGdm/qUCkLaFDGB6I+
BNKwgMKpOD812YfJkLunc5VlQz1mfZV0ohphZvCk1mDI9n2pmuKxYVh1dgRv
NH26MgulpZULakeNXwS5UEnM49IbUWrFjAWYmhNuM46Z48r5lg8Jzvvrt3zb
+2YonbyKrmuhy3CoLz9B7LLRL+B0SQbeBZb0JnRO9S9h2ys+aLctthTODAK1
6ex4sBlVdUvgG97oblvrfH31/Rg+/+EoadGLjIr4GhEUGQoV3QXjgrhx+sQb
k3e7Q+mtk8njd7F5W43IUYRbpzAkLKNpVZSBB/NGk3WE8bF+Ob1wmLOyavuL
oSSCCarUG1N2w0xx1coE+dNj6dyPRNQQkY18kqGIk9PEP/tZmXWwMGLORm5Y
S4jbCtBmfDU02QS3W9AveiCupKcOB5wHmoUS+cVXG1W+pIuiygsSvsEAGD8L
fEFfBx64iOQGY7OpIT223Xl6KXb2//gmWueTi3hYGDuqahC4hmONAPgRV2TN
RYDSFjoiqBLLE8ALEPsusvPH9Z0cNtPed+GusPaK5PjyspHAx6aSYx3dq44J
3fLT0gHYtNvzW2N9zretXEF+iQPr3RboJKy9vM7lJbH7wSyRH+eB3sjL4OAc
YFcyQYyL4bNoLfheaGE2n18hY1nHni9z/T1Qhyr0HhfCezXeGKhYizERcyBq
xYgKSKBfwl41QoPP4r1TgBgVcvY98Z0QvN3JxhT3clUun9sLSWUf2usm2zhJ
b/rwef3d0w8nVp7Cl4HcbUMknZP3Gx6mAx904WdmNkJB774zONEtLN+3yncJ
BtdV6t7xvpNZfkjfOaVyhfWxg0HNjpS9oMYtQzfxUo/9AVYGbx6A3VJBZFxo
F6LggFVSBOVHDAv1Hf9sb6GLQWTzX7LCdw550QCqW6Kt258w5/TMho6dBdnp
2vFUO/h0FQQi/L4nobJLGaZjamd9p0abYp53be7tAm46mFeheyN7JtC+x9qL
yhmX6OGQtH4S7CwBH0GxTy/i6d5tCLaQdxjdoRi3Qo+QGWypL6K4sVaY90p3
HH4Rke2S1BOgG0ttYpAHHnv578XbcnxwjcvR6p42oLRb5Ofy3j9nzWm70+K/
FULcw/VCr7lA7Rcj96kHUVzsNA/AoWWQ3Z/fx99cMTtGKRZaFSBmxYxi2X7e
hMzdpDs7cPBY+yadq3rSS8h2Zmy7KoTddIHc75By5cIFQGWP1Q+9q1C7dxbm
ZW8yaA3V2CDNMrhrMQdIDLzituxduvbFZGnezZ4rsr0KFRQQUKvL+W+rrVtb
d8IyZ9z3M6AsVyL7tj/dJep3NL1FHsvJH2WQOfO93xY0D7L6Rstabh6gD5Ps
3DWou2QNcmAB/Zymj4LMcr/uOx1Jo7cKzgxkcBmVh3+zSkr7x3fqVvpxz15p
2uiErntDqJToGB6Kh+HNY45uV6LgrhttarjPshGmR/TX5iDbkOytH8UOS7ro
AGbvh8jyPkTD6wxSSPYuEJpd8Y4JOosgbHtbqFmZvtRwPL6QDoyKMvQDWF52
K7sPggoFdV29SEp6g5fZt+oC6/e5kTFa6RF761eaa3SrUOvo0dn5nHZYxrJK
Wz+7a2O0nqve0sdYyNGXzDs36E+HqDq5j1mF6Ql9A0VcFgVGcr4aDM21l2EM
vnKnU+ASMFuBG3pxdnUkbCo1MrHX74jDsfiT7zctTC749fT27GS19f7wTMs3
M95o5xVG/pmDVV9yAOyXNQNq7eWPqm2pPxEI4+fsiy/cE72VpSaYs+asqinw
D/lfuMRxVkv8L6Dmh8yRoprD6pNUbFrFwvmoaarqWnikWD/ImGDQsZstPnAb
yKWptXN6DMeYTffyla1IIR/XVXMkU5tgtfF5SrM0gsxMxnVPpUkV8OeyKFoE
eyzM8k8Xssi9kZMQXtbIJEMhbdsyW7ev0YjKjbzb0IolTizl5mvIX7jkA/2f
NSgS557QlV4RknnShc1KURMH2NLv37KeGtoSYfr9SL7YSoMMSgKNbpFtXqKs
8rPf3cxf0z5V5/ePQlbgttzyZ6k9NqMJB8VXTSQdWcRYWlA2Xd19OB2Fkddv
GrPidsS3haLFw19RJPBbeLuiP++DlkNYKeTq1XaTeVi35zcYyC7f7G03X5sj
Ym0gy7PicH3eJtO7gDKmMPBdg+Kn6+nMV834A1O438hpEtIa0ZKSxlHcuko6
MjtJMhCA3pg3qW30wV5h7jFFRI/Fmt23dhDyTbR3i41AzRDwBOEwCnYFShm4
zfdgFQViu/NESFEoF5DlQ0d7ni7JP2xjq3YYrtawB2kOHLwVIhG/8ZOomZob
0agH0qmfyJIxjZUS179CIwX9AQKSp9OlWTqQ7ACrUvabhg1d22nWx1dCEsLj
lY+sfOVqnTjX4C8ugkwd4Ga58eyWh8MfNO/1pVkXoHtJKtKYjH1BN/kAk92u
yORg5fAMuk9v5CCbPhOlzZbv4uJkTGgBWCuRBLtdLER5yGcoge8ERLQ7SYNu
tIsCjrMyWyIumDU/gvw8kvkvzhAXqF7NgEiQCF+DactYWmkoUpEm9v15stXz
6eSN3Y2LIJCL41XGpgeONiQMNdGT9F1c6IYb5FMpZu7ZbhbdDh/B8eq/p1fH
J4IRupuTx9p11u8dorSp80H/YRTOGHavDbyp9I56dtjIPeom3nQBlKott8zg
zCmsZAPF/IbBsYTPiBjDebUJpvQwvf9g5XDk76QVdsXs57oE17G7FHaL5t25
G4b1aE3guGI8yyWlEuc+vR637AYyvP7IMOxZsV0RbuvOrtJ5RiPTusML0DOA
NzAZBkwU7KOPWr73N+L2gefw8x3k4AzmWENFk1t0n307kpCntxsI2t4PI3Mn
KEwOogwUCqVmdwRlArcf6DNcX5iuQVL2AGyX4bSfchTSXE+vV4GLleTmO2YN
lw1MErFpKhUbFNPf2ekp2SyQt0K4Z+MuUU9fxp8MwiOUI3r/7CYAJiC6qRZu
ri7McYb6kc6UZREu8kuKvNV1G4b9jB1bODdwOwMkUszgiXYbBzB0K6qbxCvn
esTMTjTBuWtEaw5DvaLJ9fwWJdaQd3/4aAE6ZicBf36x1iLmMNdds3700GHy
r2h0zybX6FUlv8Lo2Qi5JsApK8VPQZeQ/FrHJ155HrND0hiESdHuAzbDp7WF
bek+xCRoaZm+wfCJ+QRXmNbcE9//N8Kv+zKPwxasXpAmrdcqBWw7ICrpcJX4
mvHOBeH9OIKp8GTjZwabVQnO5mh0EEWMneZTMhSH0RGXlwEyfTUKIHElc6/5
X5ZF5HvhoyCXSCwAO+4khF34NmgNQJ5TSYky1wq7mKSe+PAVSW/8QsEmvlbA
mVguSGt+2sjykxdpgCmx29Vz1CypO0tLZYK/EPNsVy5jPzoyOVeULKEfPkjL
aWai0kkONWVVkagMQYlC8ZX3FuWcl7sUmplOFeBw9wjJ6Hgsj2ugw4frdeeF
3tQvb6DINPyi07jR1jwDNYQM7mjRuwWoVB2kXe62FE/UpTs/5JDLQu63ehOQ
RmOybhXN7LeqjfAvYBJcitfqxxCwGsveihUmyVSqeKlZdz050Q8XffAeUOgK
H8D11e8Gy4u55rwAfQEavSJgJvUHyyUkVzYyV46kLSDHQgoknwKvGBHj/8dz
QGy5TloRAe1BwYrAhdilqhGgRiUZMrEQ2QrzUoMEo2AmkEr828BJ5UnQ8JT0
nf7J8VcBNa0MoPJuLrJYDW2nNR9P19/nek49b2qLo0nHih69O5HWsMDf+Bkf
i8JQev1IYY712d7o/jBWkNI4wCTK7hLChW5J6t0ZgWdNC0Rmh0hJssRtRtzL
w4wMNGRHj0en8lEyAV15ek3pJFWGK7iAW5FGWukzw1A9iSk/fjA6ZzADCVFt
oiQcepjWJchmKqQKcCYuBcwZt7hgSB5WxaZlEO0d96CjhvvSJBRPpOOdl/QG
7zGpaylnS1828BSgx1t1YG+u1ROZVCy+vVDa42BeZlAsLZOV4Lc9D4LYug28
llHCVVd3ZHEbBYb3wWgd9yz9KIaoeD2pBv7t3GTJk7hnIpbIdkQb2W++Wkis
pKls8QtOLj80QkjEPCwM72p+Z/JmkOHZK1UTLSeJuV8sUs7DxSZm8nnqZ6O/
4DsbEbeukWA19LLAzDjQqw/v5k4AaMKeMGWlJY7oU8VswVvid2iXAd6VYQtY
dXvWFYWIO72k+vjrsM08qAiqGahuh0tpw4sVm8Ald/4TyCca6iDHIBetKzPP
0M7HjYYVmFXcYbnF+A8X9jWHePIuNk87n0If4Tkg3w9yShhFvzlNrs12pjmX
4htPpnaE+ZQ9fN3W0UxNXHGswd1rW+6hMTRT1fJbR19tfwuNGou4YMoFh4OZ
km904C2CTX/eqFa1dJq18CUQ6w61kDF1Aru0ETk/Lp82BsYiMY/cDpwvvCqz
AGY2bLLoJiYZTwupG3yBQa2Ok8FeWwlHEpzpzXPiLd7Dny6bTYibO2vpzs2d
UCsbW3cdVbAlO7g3nTPI9Tb4OmJ2+uFa/VEbDbmmEY+RcpjhBu99n29EAdht
QVx1wy968p7bc/vf7JVOYEr8Tv3LLntBQUM9WzkBLiTwy+oDH8K7a71MHN0j
tkpQilGmmYOeqbRLqkmMq8BnpjN7IZ8QkGBH4lPgrngDwdP8q6FJDYjzK/zF
0Qc0qIiCHzQcaDol+VY28Yg3CFviYRd6Fr2GHPm/d/SVdyt3y/Aas/1w/6qa
ggW5xs2KdrhkfvodbG6EORcu5qqxXCAQNmHhgEKzZ5IWx0Fn834umsGfBw+y
cR52iliTmtOUBTbmfFsH/d7+pFfiA1sutSulXn7hgIZu/kbURs1HRA2fPUCq
L1Hb4zv1bbJz6dNJ8gmeNL4OWZ2aziJfIUj/k4bJLRNAfNyX9p7qVHVeiDe5
7AzNjcwJSzmz2L9SpRpYGxGmFHI9IXiQs0k1/CCU4COUy7SvjVxAfm692V93
Gn4vcdudbBGbSIf64AncWV0+6zVSz1CQNsST4IMP4RvzKrVfl3fwLftIvezJ
fBZE+0OHLEJgHkT5b+tCz1LeoMYcH3JaEQEBCJXVxnHfuw6Zr2Gd0bYB14/K
rkbEgU3/UGVaqTj+0NTm2rqI+ri8Q/I9KlRv8/1oWI38hBi77fEa5NKi/WWn
W662Hu6Kij9cprb6EN3j6DTu7XbdefM6j4jNVpVc5U26bGP82yYXpkGJkPx1
Yy1VhCSQLrfTnNNUlNCsbcaFc9nq9qyFF2ape4XplAoeOPj9nSelPnUJxV1N
kdAx3Weoa3VQKAnaegzJURoZsQ0NjKyKkEhfddODmorKUOcF/84RSAvB/SQK
nJ6Ya291yIPjC+SxHu9rBwaB5x1ZK+98DuC7SaqgqIbma8aFFS/h0yJ2FuIe
NXeeNss/D6hWeEg1vsUWlBDWJStPPvKrQdkBTCT36MjgffwYx07v0DblxJ54
VxGeIA/7Hy/sQFevWQqc7shzUxZD8KAOcoNLckI37Dzy+3aUG2hE3F01Xl+0
WMMPuTttR9LNyFUrUJVTfbasB186NvfGE+NLhaSs5EPkyq5kmOpkxra/Dmbn
otZG6x3MA2x/A4ULZvrnlMwP+8+3waDoH1tT98dilcGAH/f6dQGf6IgfE4/i
aDypejGRtIMJsKW4tfZEgx3nWVAN5cu1Gr2x2q0ONdITStZzoL1GfABtoBY6
tT2fKpyWe3fkr2hHJql1hQxbKIS4C1jKWyg0TSFAWI/vqNe3RNLI3aWTFYDo
tOdR5j0TJmTeiAlIoj5wwluOG0Cte6ebExPjsNN7AR9mXGCJXlldXfZz5DVK
xK4sP97NE+tlTsbOFfe73gL2bmRSo5N3hJBxPUxQbDIlk1giJDWKTQ7GrzgS
BNCYi1prhrzy9/Q6d0ERkHYXd0CmRF2UJC0RhJX2Ntj9A2Mq8ygUIiSj6aoW
xNLVESolfkGttxiou1//2rpx5HqzV4fZltXSUQHGnlfdf105eziMDlHEjXGf
g3R/aSrVe2hGYP+SDiqMXGtSpsqehldFLb0i+glV7TW3RUgjo797fPSrDgJ/
d/uWL4Cq/zIESYXNUl/MJPmOU+opOUogfxNYcOn3ChVQfIi7+SoIZ/DJiL8Z
bS1Pt7Zs5ITr//CfKkfahZUfb9Sx+qqwsFkrNr2DT/hGW5n6dUitBNQBIOjY
K/vopPjs560lt8fqX8TOs+qexzMWmXwUDgbZ5s3lbnxZ7MrFfT7oxl7Y1wfK
jy0IlthjArMrprppbuAv8aUkcyvk9tBnBkKMNxsfahI9OwZxW3v4hgEm4GLs
JY3OttTHXVG8bwd2oy2SJ3E/AP+YMTVocC3zX0hYeavSRWIdV74RwSeYV4tw
JJCeTxjH23YzXgHJ2uY02i6qdHvMUwEf+Sr3+VbCrkbq8ObAbEho4XAhzlJl
jFFj0EFriZX+8RrWvdtsoh9sLIajR6Rr04d9DM4bk9v7gPKbzYvkMdpsvMW9
ryORSVMXh9U4qaybJCZprk+qukdCsYCvrz87AZggQXLGfsmjm2CIQ7WsudOc
smhHIGEc9hBRnCQd/d0hNwXlDhUlRUHHQALEAegXpNU0xTcwbZe7936MyWgW
oHdLol6jFZP53Z+8qk6Z/K1ThZMfUBTd4jv57btCanPwlkhPUIpffSSvM1KK
zaR6p9lHXutP/WgkW+0hyXQIIneqqnbJ9lIEPXq4rSNeiqBlYDRgM0GJEyFV
G7O+yrr50f6KRm9aiCGZ9qFTsEP0FsoWAQK18rTmRvV+og/KF2TvjruUj1Ps
HZTnZSUEaUZt8SZS7rfA8188t0x0Fw7JWEFPvLHiZbPuwjRN3/HBtSL7zks6
XcrbFJBbiWGC6XNK+a4kSl/2Q6NJVb6DoOn7Mko8wtQKsA5Zay2g1YPOaqjH
8SIgPJP6haUPFkowtOWNj7Mn/qR54fvtnS9jZ8oK0yW2taFVEdHseXGV2/JQ
iHM+QxYkFqJUhC3r3J+v6igdCelxgok1g9WMJGv0LSYSamM9UhZndzMjwRyz
deGsPJAhGH10EFzyp+rnMnFWPOY3GiVoFvnlh2L+FEQZ7eT6Tt+78ZT/PxF3
SBLndmc5OfQUKgM7lE1gr7OGhC+nmnc9k2jlLde/PAGe6BYQY3Ep7Tg6rpQa
wRgqzg9BNfBiCZ6aO9XKdXTwZu6cusk+h9vM+K4DIhn7kySSOJ1sjIos+QxZ
QCwhkl4kTMrIzY+bE8lBcf3oGnpPpJvagL1iYi24iLGuHd2SXBnKnyFmdmvk
WKVSflGcG9Ms5ejwP1ZmdyaHPchqqXJfu+jHDPUETQAKDJQXHLZN5sGPJXVj
ngYI/oFCfXywSsVEwJDx1fmr5Xr+jtiBWs/8aev5+Sobw23p1akUV3GxQm3V
/3IwuYj9YonJ+/PCFmNXmeKqU9EI6NgAdu4iGBgoJWFykpy+F4bCzncaxfob
59jxKQHOp4Y6/34YSOOPT4EtPVxCyuJ9Wh26MfjsqNDLQJgvgERR59LWGskt
daNngLA0UnFIYUWKvA64ESFSh9OLTjDTtawSpwh61fUBn/fAWqXoSC2MrZKD
FoA0UtXwpjmm5Z6FiSY91su2UGm/lKyWPVbq5GMmjt/5ODCC+JTZU1EGe87g
xMXqw7yuRg4ISCcE+hl1wuVEzpIEGwPLz79D+RWVixTULRzkHzwG3/ZLNFsN
FgqrUnDg+JQNfoclnMripHCogSTPZ/QsJcUivFS1LYPMll2Ln1u0x3U/T6Cv
5OVBCPhB3N8iEoSYGzDSmbumzjMZaBiEhKX6a/mPCAQO7xeyfMXn+VOxA1Y/
LEJBvu0+YCOYh0kWu/LExFq5GjbUbV9ckJJdAuNe5pcFwN2KjJuCFB1yWH05
z91PnnPE54gtNipdYmWPVHlnGwIJfr3vhvpEsBpMFLG9xmoi3mrhFsgg5JOu
OLvW1EvG/4sqqp/0eu8Cn5WKxWLghh6NZKnw9Rr2Q5ZwJXJgFz80NTdGWAt1
fsGwo7xIaWpLY9eJ9fBN8X6TifFI8Ppw6SkHUz2vE57XQdWFHlb2MRfrnZ5X
CSlPaQLCjXc91ORCioSs3p2CxsPbDL0wl2Jkfb9kIHsWtpnHe36FF0hSP8tf
3ICLxbvCEvZWDfK1fzmAY2NDJ56BiRYbcSGGIp/wN0gLY1AJ5Ku7bVz6Jmwh
rEkwPjdxHoGBH0bNaDLHBrtw0U6MLBe8qvzup1NRG0PAVhtwim1EavgIYU0e
JVf5OON99tW1jcyqLWn7W25NaF2iFuGVxr5eJ5529OzgeX9dgW5rGRnAKD1n
lNUmvJGwnffoC66sV4V44Tfd05Wz1ErG4jlAN2JKQG2GdnjynDY0GRj5o2aY
vKDrzfAGUek6cdkffUVSLbUSY1/7nCqeDkYGQtMlqfxL6B9C9v8aWASV+s6o
RbD9ZG1aJnGGOQOCrm8arY2EBlbTSuAg4YZCcIvPq1V5i9l4NYZ3MLbbRQLC
rzqVKT4gyVhLT9MjakoaJrFF6IVivUwR7Vf3QNC/L+1o9TdE2LbfRX+sjXWi
U3tzX6Mv8I5eu6l5rvvcEPtsFDXz4ULwNgCNNhFofN/C1RdZvC8BGyJyMiX4
QQkk5Eb8ZjPXdL79B5XmkYe35bpGh1vSb1pTJixRLuF7K9DmwtMobhrTBSbo
wkU+blbxonxwWi4LeqSZaXRos8Y7yWh2w/BEMcn7VXQ4kv340SBZB8Q751n9
uHIJ6qeHqYqXFlFTR3t4QlsRx9masrrR2F5lqUY3nt9Ec4KQlk61vVRkT4DH
QXuVPB9Uq5eXEg4NBO/C+jCkiJHdWTJEO8fILt9DhZG7HqYEhhl/FooC/f18
9dOsaF6Bnj+tUmAxoOzW7YLiLfWf8yXuKtDwhP1GD8NNNtI2YVGj33xNX/Yo
XmSIUnuc5GigLHjTIthVEDrKP66cjaKwgPikPp1IvfMhiP/okUbOPvAUSZsM
CY/3RWQ7ngy5WlJgRwtVERknq1HdUz8/js3oJJgupvaFe7H5LAihdCLue99a
U8x7zcoMkoEJy0IIGNJIctxBA5PAeBJJj1RU0gtV6xMeL60biMBNkCA+kaPt
JaZB6iB872B2nBEE8QWwTvQjhcuKAPg4KhMilEfWOxi3kPUhr/6Xu9jTuFZh
3M5bMhdJC/vkN+VRc8l7vTGcIlkj9+MWHVQ9WPFEfWhYPnKTep2QqJwb2PnN
Gv513ZQHVahIBg8XDekISL/dgfCb98agRX25BVaADOzxq3FXOVMLzaRFlKxc
o9TF4U7wcv1gWMI3GKnXV17ejbd6IvyRd//bXAznWUpAsrv8eAROiUhIFHhV
vghDt/F/q/N2Ajbe+C7ZNm5Jo8WhFO97Yc5/mqfGw5scat3KhDEHATytWj4H
Itftl6RrywyYVeiKRqhEk1IYLuo1aejpNsC6i4j/mP8nCDSg0S+1B1NpOQDy
PPBTEy3FH/dVbjRZeEODsxXevuKkCwiOL2TxziUJMVRP2Qe5ifbeeSzeiH8Q
EhITYJgOe2AjQsj9DKP0M2mjbfNQYbmwPZ4erKDwzLzTw+Lyq5NHgLI2XSXt
a4eIq8Ozm5hsGbEFvdEUG5UTE5npTQ/zaeVco1JjMORmuHMxI100fuDOXQ8X
Fp3D1mxifS3mKh790qvrbkV4OEkepisTGXHVjWPmXsKLdh9Vbkp4O3Qvqm/n
eGv07IZnirH4gI4ZXBd8NlpbdiGzTnqHnwTWR46a57dVXkH3Ua5qyeidGMlo
oIT4hikVA1A1f+MZ9w2D8XpONhc6iceO/oORUDCXBXdqhuxVsKyhCXiHr702
PhvVfHDgbNLlImsy+OSwEvcX/YGyzjOI3JcVyslfFMjjKSUiw9CxV01NR/36
I/9mFflvjX3XQB1lWjQCfqFhLQ9Dz/d258yKhcpKqCvHxTXOCaV2cvmicsJd
Si8pKLtApz/bFiwA7eyYpuOyxHrs6zFG+qzkkkrMqQKNhzdZW7EdCZhZAVLz
XwkSnxBvbzvgHfugpQel7oHrnwobiFonIkZYFcJxO6mTFplFvsQPh6rSswzq
DrFrdZ/5GB+ImcbvAvEJjKrj83R/D1lxKNmdZHEmvICdEqatzS8msAU6RUQR
sVkV815bmOzII+bm9UyYrWfXqgAn4zNvlTg5DEJkCOrs976srs4RDd3zsIpd
pjMP6wprCFj2iLkkNZ939EEOkN2w9eqMwfVT1/ijBP4UsThDvyl96M904dYe
EZDMOkA8Nc1H7BdTuMfO21IyaHM0OIezpJmrssVjXx0JRaqzg56K5VHPqr5T
0UtIFtA55H5A+Xa9wPOtnklW4L7IDSr4WitDdK4pdn/qHv0G+ffY9WzbAg84
YHG95B+lgabcHs2lZUDzW04UUF9cI3DYZSjNCmpiyvE/lEwv2r9Fq29qgwv/
+qzg9mI7jA3L8JNn+NDeGnPH+exj2FxarxC3i7ZwmZWdlrudEWxEbWLmvnX5
VMW9oxfsfTe+A4tzfU+y8z7nSU/LMxr/OK+Sp2bztzwLZVqcGpiO/12Z7PuL
m//ICH2CxtD5HQ0yyho1KZlY25i/pkhFGCagFBEy9GSBd2kWTzNhtenAXhc1
/kc9wGKENa+TB3rC6x5Dv8B2mthBi0ZxeRU5kEswXhzoMdnea2e5qEGItyUK
l4/GsM7FNXqjkmrQ+0BrAE4TsnyL7+CJRB9E8JMbEzQGwTY2ZHutjj/OfZ4T
uRq4KO/Ylll4vXDwjEJwtp5R/WmgmjlOOgjn4Q4Qo8Hmt2TtVnz9Nsygm+n3
rIYIMvMt+1NI0tOGiEO1eCvyEo9NiI9DrZ77xVDV6TMhuPgJ/Z3keWZIOKkg
egzcZ1ac3fVJVoz7ldBWIyegbkyluaKW7B/3CqDMtCe9HMJozY5JPsQmSAJh
ewdriBLanh1/Sp1DLYU0yI1QDesFxfnfshfFp+zEDgBYFcK6Z5oZ2BVAiO9B
lOsqDv6g0UltJ+zRuNn02LHWl4NRiJkwoiPbMIQ8ArVmL1NMGEcWLemNYJ0d
TAsMcgXgr5iH8UeXP3QJUpixWHq3Implrq9pDf6RaQtYT4DtEbxwsntACbXT
y5m6oDwaGcbm0N4iEtWTAz2ZfWZisJw8aHycAxbcrFYcp8aSa/0NYscKusHA
1eGwtqgwpZ+X3ytBb+/dsfuLwY1wgoDjxOqB2kyOO4Qopn1l2sl7ATVhPqHq
d7N7kmv/HsLaK7BU5bFSPz4SufZIB624wnY28WgNr9mmYgo9hRwpQ7xnpApx
vaYu/gVr/TUUD9AN3dKjx3+BhNll4yG4DcbzaEF7FNjsl+EYP2Cacw6TmfVW
IXtk8hbqZcqhpsAG6KO2NuETVnIJkvO92kEtIk+5PKT3UDxHt8SmQ5O7+fkq
G2pcp3OvqnbqGJHbq5AzM3oqP8FyN0a/BICpcUNX8KiL9SxXh1U2GdhqX+sl
Yv7ZfOnQSCtD3F9OHSH4mmNYgm7NZMoeKlOTCIN/Dejw3YaO8fB9dn+MxELt
n6jQeu5HmgbJPOFVuKyv+qRCpH5RoHRrnKXatzWA6lbeJtEnnTUEdMwudoXE
O50mtjNNyNgRMbqXcl4PCE4MwkD2DnzX3yxc3QBMtQiIODtdDZMuV8/DxFqJ
dJUDt1NLyPnP6IBw8OXXjDVRB07N5jtQEDK8fuAJhXnNAa1wPd1u4MofBCVs
V9sHCWydJnrG5UH5lzJ7SGP/ryz9czdGHQKiMuie+TIHLtKwnlO7JXXm53iJ
KqogeFYreHVL71bllnFGvrPop5DI2NB5rqRvIXThZhfNQS/63+JUzB8qpbt2
A39k3BmiHDqQSOUZGQo7087aYOYTjJeNzhb9/HkPVCGA5WSh8cpUuu4FnWgb
d4ZHbKtOn8E6d4cyeo07mEKmjDzNUnrn9B90W3lyzEm2zWQglZqMB7+gez4a
IR4DaPTfkU0OJH3Dw1fR2rfEOIVvy+VxHySwo1ABj+w1abywQzYZMt2ZD8RL
Jhi+61fCWAnepgJz1cZ7bwolY8ediK86am5+/ggY46ftGvtilO1v0R/xASk8
KavZN6UIB4thIb0ItnqorIu/0btz5/6B5EViyjjD4JlN6n7fr43Vv0lVOdHe
vX7hPt8/VmIauuBbzz620tZp2AxnderSQc/nTR9er8w1OIE7ZhnxS5I6Wa+u
H2WcwsgMw0dkBr001NSeQi585MI5a63FkwfqKhHf7m316esiurG7H/LRdaNt
cZUanUHZzDZ/1lWnHi2dLXUYvCRdzFBV7S2n73Ux5Nm2QwfO1EYziV4Qv2wn
xrc/ENRPKMQbqNLbU6c9uvhXBmrYtbqb4b8nPc17+UmN0/b0zD//EZQeKwOU
bbB5uFwk1Oj/QnhNh/Hoi2449jQsQso/W3VH2VOEAvLnCFbONQqs3uB3P+Lw
LJcZ42iVOM9+EAPqjdT3a28Bw8cLkRI5kaJ7Itr7q/XvjMbEZzw4mbGXxU3f
m4Q3JKevV+PV5eC99U91vYgmUGGwn9bzaoTKn2tSELfb0K4iLhtU9zrCyTAP
Xdub2I3AljpA2UCo5fooeHY1UpldkD/C997ExV9BMyJRyXbNjuD3tMluD/ZI
vTZb0bFjEP9ynGeJO61pfJxo/oK7O/dGvTUFRLWLX9hqpba+BzOs/FzmEA8h
3+kcftc741q288nHn61C5nw1zdFP+m9nDOELCjxMEDN6SVmn0ljkXOQKMAjm
A/J7q9f41JKPB/kdrPaSwKLxKduxfhOm2LLfKUuZ7M7FLjY3d0dI0MMG1Tk+
be71fQm0rvz32O5mg1JU4/nMIbsB4qAWjPu6lV7mk7ia0ZEtaEGte04k9IZg
QTN3rSqqG13hLaNDrWXL/H0e9W2S2SGVY0/UHsGWKNAKLZF4wFiimizTqMFd
+deR16JEvk/5bqjMmhSQCZLO0qcVr/PHMcJn9NguBLrAfRoyuNhehy/ymu97
7gQRN8CMMz+3TMCkyJkQH3OfBll5EMMBafs6Hp5x3vd2MRhlstEezFdqaZCS
npvSVRurGoK+3pFcKbMithZSM6vDF1hlNDARmeAX0NKBUiH56J0CMr0gph9r
Bm7QAARVfV5cONpVrkuVQ9hBzVezF9e/KrLXYMBpTXMsO6mK6xXtVTqWUNZq
5WvOF4RVaio4IYNfTfsH3kmhBatEoQMeqTn8ADZqQe5/YclOtNbEBWkLFiKo
DcUT5zFC6TLNI5r5v/8hfrKBBktBprY3bmuIZ9E0WoEne/535of/T2cVLzIM
1GXepJqX/3VsG5x2dB0034PMj9f71AvtKFgSsQMqcwF/GUFBPW2s/WsPaXZ0
FG8p5osJG1AYXHS+0mm3GFNrBXLKSBWfc4nhj7vVQf6PXODBGf3nY0r1Na9J
SF1xS7Aw99mNPd93mOSWRXsJfLQ1nYDVVWYlqMVETJi4fqxp8iJCEptdRM8D
ygn7RtU5u5BWWegK8gMpF4BssPHLc8JR/HMiZpFSl1ZWYJf1b+ECOozMTyFK
0+2anXR+MNveTilvYd1teH1+dodV4xLF3UCc5hbJgXuwpm2K96eyo7c6shl9
fVl8wVrNCF9C0/i6Td8/bInFpuTbRtMjjvlLYaAUlEB07l23443vVmJJ7xOu
xI0loi5nE6TW7sFesvvoyj12NexyY7K5NwkH3/S7WA/wN4Zlfm0IfdlXG+FK
RKEDf9AhgSllayLmUAREphUOOJ+kRU8KEyFtMbSXGvt2DgByZZ/qpP3VNhUI
kGC8eTXDUEaCKUgmQtwpdCcl5Q8pL1lKhgqfhk9iGOxCY6nZI02j14blmr+c
/ujZmR3DJJ7bu50v90BZLQyi3+q+2cathIs3NypRHl19eoE3QPXxpk3RPMSs
3YWr8x1Zday9e4GaGJ9erJuHiV6pph2LDvZ6snCseHQV4tPL734Kpz8DjG/Y
oKmCYg2fF69ghA1PAG8JCNDTRv2P88AHUrgseYLI7Sn7MdXeqO574dhXBgbB
CgvHcqp2Spgd9zGb/Qb848yhCfsC3gV4NmK+8yuRuU1OSoLBU/hDn6B+1C1E
P1FEy3n+A2e/Ww4+XhUMS8WJerfCahPJVfPuuY3jRCEyRpaLREi1DdFf3EeE
5rgQqLfNcs3Yh07D7wj71a7z3WLivjAojAjtg9XbpaWB9fVtMynG5tSU9Lcz
5ocToytrHOepGAsmgeW/kDOQaSdnGrH18sBeMTIeGScDkwvALY5O1uVq9Egt
75/0cCpmgW5/b0I69mqr9fete0uJ8X6EAA9iP7jbedF2+F30bOAypkj7R9aS
R6m+ipufpC+vkkbn1hSn00HT8tEN/4A/6sTZR7JVWKTqB9b3vpGACwM4p3UY
ewtOoUeXxKfAiG6ChDb9JieXdH3ZL2Xwrxlc+6YUz98wiayOfFi3svMLmkOQ
vHQmbBCVTliUVytpzwibh4QVc1t+AIuy46lEssE0OiRJljNS/BOXVx55vMWv
ub4n5Gu6KZxqtdac5qr4QwdFkPBWDEqhJhJAvS2guMGzFyTUTmjxUxOhYk9S
39zfpjAfAGLRbJhnA1+1uMsakvJQB2rXVSQtu5nPQzzKoNboUaGFKkBu3jrq
U4iitceEJebdHA+6TxAHzAFKVyXEYOlIIK59Lv0f6HO3Tm2Bmn7NvVI6YQ+a
/ce/h4V8cvSJaGMDISjEcmgy2K+vIPGIEtqBMmoqELb2hKgtbbFPKvqxJ+Y/
qHyVhrXwAop4GhrFijliSIytpf6HCAt4dgmkxqtRxp7ThAkORVM1df0+N49Y
XUpEG9gcHG2Ad1XEO0ygbJGPo+y1i7/y9p5HazqaN5QSAjkVBOdyP1lzYa9k
Bsi0m22nPjSDt/IMH3oiLRSfK9Qp5myDyL7YUaMVz+mZ6UBCnpLgu3TYb+xJ
HiAq4C4YyV1ZPe9LsWGdB5IcyQKv/4i9srT0r3+Tx5xDB/7KpTjWcki3e42o
rIK5fbfoWXY+PpBlSNAMlSQazF8tkx9H86sRORQu6hB259W8nJ3TovYwjGTH
XB/PNFCcDTtvAnY2YKwhK8jHexPuVdV7Xk3Z0wyQlRAmuGQRO41bH+rgSZmY
jAivk8sEmNbASsMqjbHI0seKgtaNPBM7fRcoWRLIIgjwrKyq8iGAE3ryL5r+
RByWw5bcfXtJvN0tjokbm5LKs4eE4Y9fykk4Wlxt8gLwO3S9q5klN0aJrrMS
10LRWK7Mhh8DyooRE1/42NYmcpztCHKoshB8g5LClLddHO3w87mpdjAq+9/f
OkER8uUxGIN2xF/1r6wgPJX0BKxwnGzv+KVuv62dgBcLdPN8TaOD7WQzJA6Z
1DubbijxNg0KzXwJlHE+QyE0F7OzfplX/37HTvRrYvPvwjE2f9dPjCKHUSIy
5KHduAncFxvSaQJGgsEnzgr8rt1AAWfQX6fkenjY3DtdvYD/ImGRldHF5dk5
+H76A34z7YtSDbp50t0P+Ktt2c/+erBV37uvqYMCKzPICOmFLW+vU7h8Q9mS
tB5FOsi+tltAQGBmPqfaF2K946jT//529rRNGV7tfgIXcdbOwY6k7r17RLU8
ZMoFu6brUc6t1SEZNYZpCkdUV0XjzzHmnKipF4n0Imj6mdsAJaao1K92un1L
63Ve8agxw7CagzGH3E3tD3WDzpBb6aOcA5xyaRBva94ds7ouW9P35rL3BSWZ
G00TGQhY53gQKwFnAp61ADliDDOXIZ5FBz2v3Na3o3Tg5GENWb8lQFMHcU2o
sbzyqua9vjC9UgX2k76SKAzEI98rRu8V252A5ZCuvDTIuSPyLxoJTe72Pbhv
2KoI/4rwsT00Y1X+/L0PV+z0xIgKeNUEG5gy7jTv6llOWuvfOr0baGwjHpC9
VFVSUSvboM0e5/+WzRbaP+oQMhme1Lpq7IGQ16d43dgf4lRnlFXDE/K0qe7+
+u5/7TY6QoSP01BD7mwuo+MJclC1IG4SH1KJp+1mofPfX0PE2j0RJtPkJv9a
qJkW5YNfWLi5esss3nylWUocReC42QisMXpLHkFGQZ04xPwEAUwR2MsRJJiz
QBVRLNGsQJyaFcu0y8Ag31g4u6bmRgD4u4/5tBJQoOgFl4ze0SS+4XXjtQQw
4l//QL0gsrk6ErrhkSR6MsyTu7zy3oSmj72+zai07+Lh++xdorx1qryyfzTi
MoLiQ0aGuRa6Q7NyvMjww6U9MnFdkyZ2dhZ2jbO8i7jaB0HKQcIMygR+6fvu
aHjvun5Dt01Tiq6/QevRSlmmNFiiBFxMPGccextczp6wX2nPuUiyKkYasHs+
Qe07emUmNDTuCIMibj+8+OKdcSb/c+iWVYwNq+l66BbIugHTRg+oUeVhJov7
j9LepjrRRoig5pvsI+4dtfmg2cBYKSNEtHk44I1SIyzQ2y4nFlzja2CJSFl9
jfuY39OPJbIiqdS9yJgg/M0d8M3qFMkXCxuq3qWeb+5jewKfbmJ+wBlXfk5B
2OrZVGAPWmHtPaew7GuoFQwW9mMhOAo7R4VocW7weFtN0NtqQBqCLZ7YfiVF
S3g3zD2qnYyfgZ/aTGBmWQTqGBfgqeld/Iui0laC8tUl9eMjA2QCQ4bMUqkA
P2PPmmun161n4NHVvoDyy8C5BXghS+Fi29bfYee0r7xbx1hcxC5hRPaZgyGp
gW27Ii9d7MjPlhMkIQAZ7jPp+wNY6xU0Ggh+Ew/0i+iz8kDh4hvLJJMIJ/1b
g8MLkkvrXl9CKer8SEx5jL7xFtCsHDTnyIrfLEDvf7cJVTjD9WUi8i6QaZCK
djI7m0KMipAa8+4XMUQJQoLubOvs35CicVJfxsmtGpikHJa4kTaJS4rhHm/V
H0kocegudi1C2ybFIAdHR3JjUBVji/9ithsV2l6ICgMzYD1Jnz6jEklIz14T
NH3i8TscmUr/I/p8IT4dKdIhJeod9IfUqKzggrc4B/2BFTyxE86fLrF6uZUm
EjjPsrfr7ONaAuJBrazV8Jol7bSQNwXKd5fR2yNur8bZrsQJThs2gh0D6HAw
5rVyysJiBfdTUngfwJVLLMhBcUUGRmaQP8As7rB9msk/IeLmOJoSSHYgFWBF
xTWf1dH9V07CLUEzt89oZqLQ/t/G1oguuEEbtAwr49OqqFHv7xBma26q/Kue
5EpZ2QET6aS6wDYAhnH5MryMFWeeHibLE8TZPkmootISMTWtUlNrmGUxuyOi
k95lFlfZqo5QBW6LCweOrB2XAohEHyDDzvucZ/EKf28laI1X/JRFYIoZvn4q
QaC7H1fyCmSAsu5uTWscnQfI31rkXK1oVIY57M+eKFcLXAPPuUwDgJ/rM9cH
fHduXYIWZd/bNTiU+tPml4lxIITS1WQ3chBSy3rAXVPqwx7Hn4tsMlCwHY0e
X6E/1TsBeiDS4eaJ3ttlVVvGW8rl3rJDJQ6VXdUEtWXqijPNu8pcwcZcW6tT
lOB52T5xfEuMhLW6Af8L6S8A3JRf5PeXSUnyylxquwB2G+fDWj3y2z9+Sfvn
p2nc2hOTwCjKb0qwbU/BHKmCayK0vdcVCsf4JFKmC/qZ6Igk7yqK+99AEkTP
/6pLV1A4LaSc0eQBowIjT6LdRq3E9mJW+UhXumlw8vWKR8bRwBV0p7l8khec
9aL+tdUqAz93AKOOyJzbzvWxBLBqjDXRL+yCh7WgCKh7JyPJLpm42PnjUNuK
r/SCiPtCwg+AJt59LSdVrAhOnXe/ShMXZLIbWzAj/5XzzEuX+kxaEryu9gWU
64F7SEZ5FD2XmF4H48/HghpUJeVmedBKt6+Iq9br64d+6pZCgjHwzt6WcXqj
DokN35UkZrDwftjOeAK2jEJ7JLY8G3AFGaXPBH7+QDh1hDWD5H24sfSQa+tc
kNoeIuobGVDGzQZFW5GUzsozmLX8bHYlXRXll2BIhd/xeQRaBb8MOXu4pWHk
XhNIfbyQ/htLa5GVGI8yrPT46+1d3cjlvouYy3gDY1zyx40BNOS9KX30Hv7z
TKbXCCibFEgv2GTmEXHhqA6UBfCRlZTQov9UzRv4Num0JyI+saorsO8s4BaA
FWZlbE0zRmc9Zq+IsBoQjbM5IXbJ7xab4fd99Jx3h5cUgEYSqhyAkdO8fgUg
p0ZZfmDdtjotd9wm9m03Z+uFgoyzx35JRl0xfNWyFyZjlGiYsYgUky//gG9m
fQFL+v62eustimcvOikHU734C4PRetRldHqirRdsfWoAZykzD34uMnTMnMmE
fwOanLFmxjG2qGXPfWnK7TN8+zwX6udkVDLfpBLHKbl15dnMJCVXzR8Ij7Fw
pkC9ruM5u5TcdqtyUgB80rEayPPay9914z6HE8/pvIzW1sozPvRp4+mCzp62
Hyi354rB5ldjKhLjt6KO2r1a5VkDV23kic2Tu7h/XprN1GyBDyLItrQuLYN9
4ebjueHc37EAYO/J92SJdYWrnV7pqb2bJbvPaMauId8SqW9UvP53ccCrLkpq
6MrGtt8vyCrCrnvh4ACgIIi9r0HOzTVUIvEh67QfYmtWr8FyRwxYivJ0Cgwy
Bb4K1nZ4g/Upm41Ge7i1BnDHi2HEAl98DdQdI9WTnG8BK7dyKp5Id0Y5fufR
Wv2d+0UjuytGgWhXFlZNBgzSIhKinSoC6IEGdu/qktCwIUjqS6nD2sZK+6/E
5aYCAzd4HHkGQXCEqSXcfeoY0Srjtj/c/a4GHg1fn0j+GRkShxPOU5+KgBd9
ktIMK++bEco6KxF0mFZ4O1tN3X8DWBxCvkaUxc3eOBmCvnLgYkQ6ZT+or+BS
WUQpT1aMoW7EzZLHcdKMoYSwPRMr44kPuB/Pe3z6+FHV3IaUW2Sqo4yx/i9Z
t3ncEeLEvyAT76hUBqXMGBDsMAdfMHQUwdrFJpLKz9wtkb2+uFzmxFRIZDn5
Jqg8w2bDMrfbwhy04ZOvke4GLKRw72+j9wzhxrTR2mXO0Vlt7gRHH+LGsq2S
CohCBdnuxMHKpoRqBUJC0Z0NGppHwcSv/GRa1pSknjdkHJV5Ru/fvKGDv2lJ
coCvFFRdyES7S28WOQUhSesM4mNcJ6IQ9qkrC3YBWMmGfbKEEbHeJqQk1mAK
nWfvsCVAXfmQYVUoAxiss9p6P5sbTF720OCleB1mkuidbOEJjRnsvUIeVOZ+
GwgwzXtYQo0uGrkTpsetiGL0uA45HPWJifKbNXJSZSgMM0wU7DBwWNR9l9gQ
J9TgiJU+NrnGuTanNRgw7h5TvmVHX8Dyf75l0y5pzB652SFHRK3D0lewcERZ
fFlAnMGnT6rnp+sGCw74sGK17B/aOi5uo2mrCui6hqb5rLTatu9j3ST/hSmr
dWmyUlgukWmKheRwFy8XiwY3UiKMeXb7C20tIiBVZSEptFubkPAcsBYb+MbV
cmaKOv+bI1U89WKoPMzT8MTa0aVcVhnYApazcVpHLPnjai9fhNuEuHNtQYg+
6Fw+xVKt7sBrHRbZ1gf2oGGfZb6JrYvjow+u/JTBp9ANxmpD5j+ytC6QbEUj
LrvBmUI8mbF9hvhy7m83fyLDILUtWjC95O+l5Pwc/oSzqA+tGsXUOpZbCQBv
IYjbJ+qjjQb8lG97atzM0fqh9LGffzoeZEbSs1DrXsH30qjZCBBac1qY4KM9
FAfsTPJCXvwRO5dN5RkGJJ7HR04C9LGzjiSmKFEswC120+8CtY706aGmkdFK
4G+JEiWHz1RoL3xk83eU+1fmBftUFKkDmSX5FGdNxBz5rZHWgskm3IOWg32K
0dRTZKYll1hDACt+lYVTEklVVanPWj3DpJr9geLrujUm/UA/m7qm/JtlVIVM
RWNo/Yw66oJzasL2Aw/+AWrH7Z33In5XXnhv5yOml/X0F3fe19M9W64bQL41
zkzc2xQC/p5go63H2yvrWXjtPPlOBqUO27FqVXk21uQcS/fDz3brNaaH0QXn
daFOWY8P3V7S13sAj+GtmvL6eE5H5kYtilX3XJVQL/jvFyDV7z5E8IPBjQa2
UZy5toVj9ryDb85E2lLrQIeaoDwjMYPMjBP5L3T2JKBZEDTjmYXZh1bA5q9Q
BZcMabw3Hv/rsq13LGbqK7kou1C7TN/uSKXtapdE4tCKLLZ1Qh0M8Maa//SD
BHXCc1kfxpVIF4x3UMs7ulTSAIGKWl7ZZBqPqkZsJ/UAcF5mTquBH9SII+dd
a0Hu34SzS8gJ9opSpZTeSk/snwcldACsFKsKBvtPQ6Z2/GVkjhygSONAw3d1
hCXu/xaV4AS6SxOwanoi7aqZfQdLUJlYrQD1MgG705UcAIVdJkMdvpDF7ksU
Za2wMs58JUqW/qESf39O4kR9rDGm5z1CpVhqxqfv2lzQ0XL5pOKQEdc8UwFD
jUsEgQ+c+mYRMBMPd9i7gyiFv+NMBWFTkoxk20Z5V7PC6YiUhXMr0K95B99C
D4egNVgdFdTrEzSJ0C+XvQFcMvGLWvoP+Q0VMBx3TtYEHqmQ2FqtTrYIDJT3
ui60LubhgTNlKu7WbzFGLVOHZvzk8lRU3k3d9Dy9no7GkN9asWu0i6GJN81s
Gkj7fvR98R8kC429IDrAA/9LG0oGPznGLV7n4xzzO5eiJRr7o9+rJ/OgZscw
8yJJ89XwwzlqcvR4F4baXtNynSvSXj9C6UfYBfdqC0sOgkvGSvf8hMJcdAus
9iZZiF4r33Qk2vdWahwICS4Cx3vCreTLwrrvF7dFjhO51JAx6gHGq9g0melw
/svkIqJHn5WBQqVEDxQbWAWsh4knd0e6hlhd3Rb/ZoevUgpEcJ4yG/DUMWhi
hE4VhYOj9oFl4iyDZqgDFJOOpRGcKUyq+e/Q18weGaGE9qrwe6b1jhzm9aU+
VchkvP/8vHtPlhnmZUHvhikGf6pcK5giqmMu4+7L86ehirYt993cFg23t51W
DoOBupWaRorH14xdpZgXJq3yhPLCtq2QY5gz+KG4MiQYQQiMBPB2kySmxM3G
fe2zVmpcBT0aZYLbTvrtgQoZu52QOcjHmUGfn1Dcnp9QxTIl3XuXMHxKkehs
b2e2qguXOEaWDkql1Xrjy9kmfNW7zevZSsE3hMlkPznOqBFmEFXzgeYtzFfc
bK+H+y+AGailhRw4zQfwNX/hOhj8f95/20VwYTV5f0AZgGEw32ig1khcpnN7
33hZYOq2/r8XlLc+9TYKYZnfmLDzRYIua036G+RK4Gqxhwdb9CAlikUgNBvt
+YshSK1klkSR2VgW5rmPsp4hGZgNBmLYgD/E0UPUpxixBuidhj0zc0eM3efP
2NPSqLxBcgZPPgB3F12EFcy8sKcv2dx9XteWUMxJOohYE9K+sYSZ5ijZ1VL1
VVCu77jA8ebVlm016Lu4EWioJ2NQhXsCZ6wwm0OrcHT4B6bD6O71Q44rkFhM
HdKgsyLfvJRjv6+iumTB/yUsflYJpT1ZPoa47zfa6LSXE48JZtNPJ+0fu3Ri
t5YiXfla50pSmtl8dJ9PfBXBSaWwA+B6NwHDd8+qP+xl/y/iIcrNHoyS3oQq
70TkLxbW1+Vbl82lOJFoHYxuHJdkfWvssSYsmjPrJyd7H4Ev4zsmgKeMPjei
ND6cwFSGeVf/4UWnEzfA3VGHFN9rhYe74fNMbyb6aNg21zO9lNMQdwfDNiJQ
OHAjZd5vSOaFDuwVG0+26Wj4Bms+1KHWC17NCEIcCQ4hQ54BvLFWILtMjcr4
x8ZDHsTsJuzgv1teu9s7zcevAzmhuWj20j3gRWy2eu+DI29irJIQAZsTCQOd
bpGHO+jFqBVI6iA1pIjKE15zC9KBnt9mNgdDFA7GQehHSrqpRjo7eytEX3nR
K7EwsqiWvQh/lJ+HL5cUb0uYt6pyR3dlxl5XKWsTuqcXv8c/9DvU5rN0fUqi
wFP2Jr+6OlwF3WnMIvmyyAnVKik3IA+TrVXLD6NNjSRFa6rHxpl25RNUeWvp
ZHgcz/j3yO2FDswCHaZNwsSdg7zdGugC1qa3xVZI+Wc+5AKUa9ZbE6LNUeVO
RMyr2BMQkeEqo/FwTTFS/EtKIehG9YMMlRWQkYr92+Y+QS8xoNwI7Eg02tUB
pZaCel9mi5ZUcAngGfN/2k5qVmuw9QsrH5wBfzKWjVG3bQIyklcH46E5SbX1
PhDdF4rjX5ayrZREpZVq0hj+S8nbPtNXi7hRdgFxhFwwVMCEKy36sLSOkOKm
aV6MMDOGtFXYqaty8q72YVJWjtpAOB3yG+qID4NiwA0317RSRkgMSA/06Wnb
5tKbh9RIq3ym2ZSs7dm3RJc+z6Qs8jXn6Y8QzMGohWekL/04nQIyjxHOUE4O
QqG9fArLraTGbU5UbBd4vxc+r+vLWoKjo7/i91CsTeei4Q8cHTBUueDkDSy9
2jpILv4vTZPRnjvGdkPvYM2UQJyOreexDsLpH2l9mqPR2m/cwcRYcvMa8blW
y9/1BfYKn3rj6t3LtRUPRlNjUtj/BXPX77slvMmGvzf557xH5U/WGucfPvlB
nBaMtGvRq7hgoVTUXxmHVQA6Lb4cjB55pSWemBSOEz76EkiSrFHa9rLpeg2x
QS0y+gI+UYX/y5Fg81ZkdypW7XFGRwgsWZ1MCAPGY1Thx2K5c+u7wNGXAgY2
KZw4pOPy7YayOvwNMp8pqN5UmPKwInCb7YHrKQhOvwLV1JbWIT5v2HlWDTOZ
qV3WvqwDYZr1w7U9YnKVrwtZgoHQJ7xDUWCfA9ykVmDguM/AhhmQfXDrJbZp
YghgfZKSHdPT6KUOCmgeDt7Wlg2JjJiHvaPnsep/XnM59Uz7m69XzkUv833T
G7pS7NKHKnKltZ5C70jsFMClvjDVQOrVnk1D3mBpUgFtQp6Ix9BH7C3jx12B
ITsxPrBe64gN0VP7PMQOvmc2ODUeTmpx1++DNAQ/sRVtXQBr0ZRJxUXooogW
fgCHUFrFiM9SALdGINwU6acCTI7Eit/O7zYNu9GUilH9DWDjLizpcrUm2RHd
qr/DVj7qtf00mEFGngR9DS9a+4W7C0HFBaYd4RR3VfTnfL340twFuZf8QDtS
T1mK+IlRhQYFBjO6MxO3gSwFcRK8/l09NRkkAz2DoWUI0F/Pnia7p1vbXUqg
2K4G36lYN8Q3ul8bKt8pE50/lS92e+dMHrfExONoyodiaB8ny3Br/RdeAw5r
dbkKA7l/UMc+cugMt+KHHu6WmEwp7vRxH3IC2e0QXeEaol3tES0TlQmEkMg1
HcToyDwY080yBpDa2ejitcBBqxbxO2Z/KA8x+WHF1V0Ky6x7lsx6/8Clqh/5
X4XdoH3MLoSqBJ8fsZvKP6z4QuIvHcswVt1hG5lklm6nxLtv63Q5WNQXUsdb
Jk5LxTQRkfLPw341MxhXgE36S6g7DdlmVqQ8Q+P8NcE19nNu9CAWnRAudPzg
dXlbXjv3je9FwsyuW70tlMwIuI+GJIhC8AFjs0ihcnW0sxjprwSQK06tHo2r
s1ZNO6P53ylfoHTs2fUofTn6LwfOu81uOOD5qzQpu/RubVC7Son4VjVcVSu/
HE5rwl/B+LkoosOK2IqweE+8Ah4ga5zofJ0Ub/qEdfcNXCWWpBS3c3c+O6dZ
SQcQdSI0kJ2OkutslM9eHUcNN5Y1YSnJceShnT6AzJ/LfNqn7xYdvm/2djTC
ApIi3PeTIW0TNaIrGUVxvsuiiQ/t0YG6VcudszPqeNVXb/k+JTLK1+uVsRzm
uNLNCpVXYnwIIsURBW4Ko9gWovNQoXej0qaXEK+wufsLGnACkRInFdOZ768T
mwfmwe8Py8nY2fvJuBBgo8rY5s/kmREBLPLI6j8adbSJH8ZrIVnOpzjgxMHU
+3CogzDIGknTlJOL1wdzpZR90aRQJRFihBAKTBSjnhY/KZgBHmfsLIdDt6sP
E87/3mzT0IT0izq/8lr8RDEibzC/k5fuPJ4Z/YvxOonoIALgat5Ij5uXgeR3
7zkIGE7Y/sP2m6TRJY3cvjn/iW09xai2EfrXj6I9N5TLp2X3aZrCrSNBHUoF
RBX9E68m99SlIntUmVi1VvQA4Ig8V2BuPPxnsR+tvMSIkUBmqljIt2yxUE8U
FFvMqXDVU9D40vAfUZRJyrN1CtOuWbJBvbMvnXXpJnZiUZHNIz4YrciKzw48
07pvJkLBGSS10HAOF5hYmrqlnuLMh5bzn2HYLvLD+r3KGzMlS6qeo+3ObkHa
TfRAvbjDtqoldkJtAPl2r/qEkcZ/7c03R9H/Q58iwmIjnMVHEniBKUU5VyrA
OtjNQlUWHVttuZN6opS6HAz8nR+V0zPWUY4u+qUDTUXZ1hu6pdR3OE1AlsKK
LyvGuCg3eCGK3nTUjFj1tZh5Hpi2sO8ByvKkP/c9N78/hc42wrqmsn9zdgI0
7XJ8XNWsCE/vi2s46kLsmjuxYe3DYxLibqk79MlZuWFXYG4vxC+oLSc3J5/C
+jtIdSeDTytxRvLVCVFWUT3Tu3GmQNW6Bo5cB8vX4OTEdbSewRTHLX+p4udc
k7Rn5BXk0rwpDJqOlOAWdQRrXLBbSdIAWPcHZcjMlu0YnPlF7kXw89yGqetU
3gbcxKyrfGNUIy+mL7xP0pHVB9mt/QybE57nXgvLcj4oeN9s1MgyrZh4QDMj
CtjeyKE9Uv5i4BQv6WK1Vp2RGl5lyzwZyDOzVt/ZnsNOdYYB0yZqN6YCODpq
jTnr8DUvn0oRYIhcbn9vDucu+YGFwmW0q9WZetgnrh/uUuIOLbQj8epSiW6E
QMoFkqdrW545kMdOC7uocueMPRisYXbvbCgz129l3XIFvknUDJyfnfRXKERx
Qv7eTieF0h2JGkzoXfYHv8qCMvLPCernonnErYljXKoNEEtwQCzW4vmFjD4i
hev2D0vy1UCy6A2qNjkl9rJHVn5nG/6GciRM9d0we68F36xQz+9Ju1rzZUGd
6UVcA6EE69DZ/onkILcQwk0ZespWGjtfEdlAGWvimJ+dMxI4F8HbMNErqJjy
QAixtGYvJtAVGSJFTuX1S+iczPEVeZ6vhZd7pIh+qFi24WsbxjM9OeEVXCQ1
ojz6+qxkOnunAmr3HgVhm/RZ8L4fGrZPZtr6T8mgaBhZk1CD2cye5mEe6CRV
FmyEFZ4TpqnFLj0de1UvEG7PHY51yPBTXkyJkvt08y9X77AjIKfY8w+yXvUw
tz2XM+2xeKw9RLEah2990ZiwUCGsqzKiAv0PV99A6C1wb7t5NxWgtWK2sNlO
GPWBoNyWMARDEk0W3JAJ8OiYPbr7+bzAH/FS1CIfgj1/1UIHrvahX6igdQAa
MwyqRrU5Hl0JyHE/9ZiBANhQxFhRrSvtcQNyuonXBrQTJHOUaBgdh8S0CEI2
Lp4fT9S4myUKdr4Q9tqjOndP4ZSH3zTqiiTd2aIYN/5RRyaBud1BYaS/j6jF
GiYqjHYCP0U3JXZW2Um5hi51wH1Fflbmj977q054aOaqoEr4zH0Cqkjj/1Ig
UrUqGOXAQwcdF48ocaGdXcjOlni/Z7tPcvEjKRhr82bOL0LWokkSxC20XraY
BKvRspyRyFIPUHTLSULqF0btBvz3VPGSoXt6GHllV0N4BExv5FPo4Arj2Ika
Tj+tGSyXMNsbk5af6Jmm3rJR4rO1Lse6L9JYwBUEaqcnnjGUeWbB7QSBCbuy
NNSg2JbovNGP8pJSeA7b28Ir2sQOCqWIdyJrRsGOeXtjdI8+cAA4LnRhVXT1
bfGpfwzPVqvKyuuCglKWu59GfMebhVc4NpqQ3v0GajB0O9ALmciEiSq7mIti
hHGxx53TQiF/pbbu4F6da+mgH/5BKSqy9I8CgFb5wc5LTarwOqrfLBZFLHNC
WwYsrfnLRzC/X9jVW3gI1zt6QYl0P1d1w3LGHdQxe49EcFr75tu21Ps0aMpU
gDAPr8M57FlXCVOOiEGZ0gArf0A1hd40w2U17mMovb8Oq77Mz+69Pc+GJP46
71AQzXrVya7/iAiO4R5RuPL2jPcu0TMBbUF7sgtn568v0fEkAY5BKA10JDaO
xLrXCPdDmeZv/h6XHqA07dSHE474LK75QKYnpVQEBmVig7cjmGkITCxzm4LI
7Jsz0lXWBP50x+ERBWVzaGZeKPyv6FFCmgy0c173vbM8pvSO1F/y4TmzjAJs
AcEY/AFUbG7lXZJLdhY+U7BjqA4/8cJM08OeG2oaKDNt9t06Fu4/qL3bknnN
dpntsQIS3iVY8+tUm1JvCB8agsOdYAJqFe90/Elycrx5D7nYjZ9U//c8XQHz
W6Uq2rag7a3fW2Ooaa7eZRrqiFctmsCWMDg7GKjqmB5xk5SV2xBid0Z+cKYL
hCnsRNBUAH1xzrortcCkuGKUhlmguj7kPwCbBnm7+nNh9sbLeqz+ZrtMQy3W
ofIPZwvqhpQefJSmpv7kUI4KfKwPrI8RNcPWnHSMFo9cB8wFvydgrsH9iWRY
hr7m0iriLczgj4oEX6zwIObIYW3RXFZQvxlzm6AT3G5Ghwoz/ffzEVmrIf9N
bUuUTwhC3YwWhDE4YUJVf75/Mnx1HObMqpYC5z3EnappwPOx9TSlPnUUk89s
OyZfqkrHAY51btt/adEtnO2CzziixLl0RyopgQyXxStffTW/37VGycxE//4D
bAKyECuvnY9hLYNsaE2p5mx3pPBURtnoYU93Qzj+MxgAIU2ET4MvuLX3EFQ9
6BxdiPkeYS1TgpF19hBcJqGfhMz5MXZclpiOwENjUILv3+Kqy5NnYs9LIYqF
lgpPbLP4rluNW09acT4ylBuRWpC5RB40D1n/en0AMN/XXAHiqcB1bHeTGHAa
zoZ7cMJRyCH+DqXwl408N2qjQfTd5MIt/GY7rFR7vtzDR1AUnfY71gYz5Q2k
2/hz1rZLoPT9nTlYHo26/uLYET5YfMnkTtnQ2d9T4zRvkL3M1mBaF6iflRqg
bYFavcI6wljY1CX4Ah58hA8bDnlG+HLQq5jAXLSHidcgeLxNp3M3DormsQsT
muFCO12izDi9QWkMfZBAO2iZBS8P9wD4hxQWtf/wHXrTG+RIi8REfhuadGK5
CeUO87wUW6AD21G9A0WU7WMJEkEaW2het6WKzWumoc32UhpI2ph0LjEHILxt
XSPm+aJX2kcHWbWH7UDOlkw01QDDlkpkrxOuIq9MoAwFuN2Yiei3VWEWUY1q
35qFqf70SBMdyQaKZ7IDvzLH/V3QtQ5tbNSKJs3woCmwI2ekiJsqijjf5IvO
mrnzO5wuz9q4EOVmvBCCAznMNbD7ZUElMrh5esf7Mgtuc95Nod/pZ0ug5Y4Q
/UFHk4YhL9SxD7BIHoR1k8I1is8yAYweG1B+94d4twQIOFlzi6toPX65Dtms
dDndnAlx5Sn1oIAd1DNY5YHVMBisNAlRCKOJ1saPkC0hW2pCoerNMF54XJf3
a2o3tD2qgLLPzAZoPAs/oLU4B5s2j2CvjZE2+CQ/EkA3fDThYf9s6Xr/SJOJ
OZbyLa62F0yt6jf/0ax+T+cGJbKZgnD84lycJFMPjRIh9hAUVwzCPED7NjIU
4Y081Bhu4jmAVgGWUM1KuUuaCbYOOj/BHk+7kdWHwDcnHhjRUWZ7ucSeYUL4
huSy2yOnp5oHen/S4c0IcwMO+rR3qAPqCM0JewgoT/u66OGi9SQrnh155UN5
DvF1/jzONvwIXBEiD3DQzgxMBfaIPnDGVHe5Xvzl5xs3GOXBprTal3ER8IMO
QwFmSf3z0lHRl3SNALYmqQm+SlkeNpWDdTcjxJtJ92PtZBjGw+MyKZG4z9Jy
Tt7cXtzLXjbsgyUMXxECoq4SmCEPrB+gcDydXZ9R5k9JjWbGNxJrptiOSc+h
tFzgs6x3HkP3Fws+5d8ouTVoNj6LZUEEIyPdUT3XXjY8LL4UzlRs6YSFDxD6
b+8+nYBgD6ZrywK0zBVsq4Iy33sfV6eOtNKHW9HEkS9EveGDo/t9j6YXZqn4
IBTkfPaEPpau/Q9e41y/SJ7aG5Q+dTp4qBstQ5OvvBz1XLMrhpkpYQeZsWOY
OeKxCEz6gbol2tvpFvuQuTjW8cur9ttHc7+RqPexVBsZ+cFsCC+dmAshLiPw
4UfCpyRmTsx+DQgfmGqUKCVMcOdz/SvIrchM0UXvk1H8+7ilQoZP5drc69F6
6+atDrWrcGCEFGg3fvosBugtDhGLrTP7GUtLydsdZGHIFA/LJ+xUo8JmBAB3
KwoodfSMKlI0+7EVcmUaBDBHr1ryf593eJ2ksDUU3yAdWxHSsYRZt/+XRIy4
Jmnuj3AwfUBCjRUTx6L3HYXZm5hiBj/mGVM7QBBhpbFnDvx/A3+plDZEtmWv
opKn6EIaPHtCfxhQ7915iIOsRiSW4AVH4z3IPo4tI3V4HZvdA9EU8I5dqPaw
2KpLYKqCaVWryb8qqlogUoXvV630VD2H39RBSmY0vaJsoaYKRaC4ZYed8qey
S0teOu14T06V0mxdFikAtZFf731H57aXVfwzfErcjpB7MphBELkkdzbv0gGR
9c5a00lRu1i56NTzqMlDwlwAqR9/byNzGNDAYge0VqYaHZCMIa5zdH0lqsO6
SzFt01Ng+d0euTkZZcY4XLY1QJ87fTVovE8Ks/5WoMenURCh+x7sxznUsG36
wuWv3Oo4EVqB1B7XNAP+WdRD8a3WriSwJncBcGCCwt2mDZKj9dYxZK4YMiKf
kCUFz8G0ZcRe1ZczWDbGYtkk6P2BTje4KmzrYIcjJL1YVhQLKkKriv0sTKqu
9NJTldPCyfWbmb5E6kA3WisYp7/JGZfhb09smZ7cqwtUvF9A4I2NrD3rWM0e
wJQXsowo3YchsJFIhn3mvi8OwGgH8phU8HTOpDEt+sCgIJCm9Iw3H+S4ZBui
2Gou0O7IxamYDdMXY2nh2YF3GWp5l/v6D2JG4fYIB0mROgfyV4KqCHxEiLKO
IGCD6QCGq2WBnTZcsbJirVhdYzqJtIU0BroaQR8KBrdiGORi1i3wRnUC7WqU
KO8sbggI5gfmZ0bTGZ0hWRcOy9XrIxaUUEWxneQjI++T19LJebsEvcc+32XX
BkucF8H6ft3g081L5TCCX09Wau0Mc/6futKIW5EZOLvAbBAYtZB84RHFGJ6K
MKjknfWlQkXIUD4ApE7P42K0CaLgQ0vXs2kC/zyunbJpRqVpRRlf36AhFei1
BeNr/wxfJnm5Yke0B0QttlbHujSN2D4CDDcZFwW6pSuL4USBSuwRcM0srL0f
GPDy134M/RVV0iZB+V+LYZq2tgdqrtrlawWcjtnkYIHYLcRhh7A3v6/SpH8+
Vc9CJtvVqvElrwyxS//ePCvg2okCvEFC/SZUuNDvlesmxAmJCBHZ9A/ASjGf
CBT6QIeGPXfCcKASdP4lmiIs+q6g0rpfYGCnl4NmYgNnPLIHSOvB7MGUVyU2
MpAcAujsr1ncQ7jjqaNsXVWppnjgv4+fdqxAy2TErJI0R6gsBkqXGLujqitq
WWH3l+gOTV54vw8foCJtrwDWA+PCA/+SszWlb0dTyy9FvOm8p9oRj2xZrTHx
hQWTUFp/ryQk978zAr6UmML9XuB6QPB+U769fKIEPnAbhWFvxbPBZLVUF0qq
IFWHSqaIpLv3pPD3cCivxHinqa2D52vccMbwQ9y+NM1+ZL8Rttt+I8IC6+oz
0NVQD4RAQHG/GhWuRTE4t/U3VQgqPXqxJ+wRm/fjcSRkc8g92FRpHPYYGCTU
bAidNGzVi2Q42b3ZaPRn1MMDoPpUmKTYZz3shKBzF2YW77sejhU/q8v1vtxL
evmojtIO4s2b4oduL3E1rr+ntM8KJqeJ1LQ7UeXTVPgo5GIwo1krT04dqBYW
bMvxY8iCo8jHEB5vfplIwy7FTnA0nrhk2ZOkfpNLjvTbVIKCLNQDk6Klfbmn
wBZdslwyx0ushrdSokibErIpIaOfEB+jj46Q46H3TRhiW6hm9V2CKo5iZGXR
Ja0Bw3bo2+QUzrHB8GJa40b9B+fbaMiPQhqzN5IvEBmdaWG/9mzYmY1etXfx
QubBkX383WrmmVcTrB90137Al1h+qTmmB99QBVl9aEfEYuPMCT5slkqn/yQL
0VamSfzZ8dkDrjj8H4OSwueIQAFMZgrPsgcNSr0ylD5+R+Mdkme9NtWXUXNX
/bZ67Ey8jVhgvGow9QQuzPGMhDU5MWPOc5W487rmDvVbjJbYAdpIFhEgSH/S
CkEsNoiUsmuOztiuYUb9462gPtbkgxEuL3sQK4oTnQZUvV+n1k14FmiibLBN
CB6aUBVRykkymUdiGeVl/6AOCaY3TwkwmJZh3n46oYLc2qMuJEqInuyd2Wrf
tlJnU5vm77KaWahLhWmgvBGUTFxfNsJEVSPDZBXYxQm4m/nPGgwaZQei7p78
JqOrbySTpM09hI7S6+nF6rEGpEmVw2wbKHYxAWTj+DoOgoTKtd+m/4cM9wMP
qzbD99kb24wkspMggNhD/fipEbBzGPX3IBUU6COanPsPD8OlSq0w6egljExx
7VwaHYtLlhK2dlz6X/pQVcjySot4TnetUcDj/U1e6mX3aHLNgcckXvR9T3jP
VO/VcC0oXVtJre/QP/2ja9jkMGkrXMNT0h7HVF3XGVLEpCZNTGs1E/gbFSsq
6xLL1GF4NVH8W+ezLdNNc2QoLMIFZQoQKcysaKBVT2Xq9DtCptCde4b0Ui08
eDIrJU+fmb8QWhAxoDZ2ni5BN0GJg5Udhg4szaeVOz4ACFfxnfsh0uk8BY0g
Hpw11P0c9PwZg/7rO4DIOcaq1yI6T6XeRVqyCxP6yJVDhUXbeqsVdw1GLC4f
XY44vEL3EzP55A0R1V1/8ZGILnlldfEgIcqpD8n/mTsjZLeVuITC5ThEBnzX
oe1HXl//LZs0ChLMyz7IIwzOr5GUPGE6Sq7xVJ85ux/5Vrgh91BTDyfkQ9jX
sLt6ZJz4Z1j4WQWodcFVHI1g7ktG5XCi1dstTdJBr5VAuYGjbiOCKAOmIiM4
XnMgEFKQGdwtvDYGe2igXRkYsuwgAGsNaupEvTHJFFsF7IVLC3MMrSQXK1xR
YWKJTxWKnwdvmN0C5Y9gaGjZ0f0f/K0y9ztTjyEmKYaCHJeQR95faSb0AEoE
cEazaJjZbCFezaIXcCicdhWxywOiaQmfbQAlu+jZU5jGe8ON4eH16VDypO6C
ozunmQ4fYN3aOM/kqtwmNKaxl/RpDqMKHUUuiOGWCp7gDhw/LEQL2ZlrjvOc
ajSQ3Z4iiAmnVihq6ktVCnGC/0PNXPOqXmMCfDbZlDOaS3X1izMABWboRy3f
tsBCFO0/sspokXx1b37aSxUtjlqvc3Y4JZXnl4Y1LvgE+zNcvrAXHwnEsFVw
9Lklc9ORyGda4IksgzwFgNXJFFx6GAgEAd6k6Mzhra+MMqgTJ8QoHB7kkSES
fijyEronZKw3ktzdkEA8Uf4FNRgfgm5qp6rSicNf1o/wy8u3mFLQ1hI0tR1f
mwPD1OVwPwWkONZw6mORkBrUdhIKNRLpQjuV+VFvlebqvxWbssqbgJM/GRh7
cl5cbDs/lx4g+bMzkFqOY6efvz5tes32uuFHBtynLb8b7Lf6xx+GUIn3uMSD
b9Bwjm5w44bXWlFJVFVl6JowrBP7PlqugTYQrgIR/DFmxTpqJfGeKYPhGAjx
pqd7eF5y3Ye/PJDBnkE0bOyYpO9I59WKQhQ2S1j/9MRKGx2JYhN407/ams5b
W8mHvV27rhKO3mjDxMeVvuncxBXOaXIQIlyQ/vFCEUvb+4O034tu6JqP8zp0
s0m8wW3jzNS/eLgDIIq3005kg+ASJ3tcB9o8aK+AF7d6AV+4sxmioIkZWu+y
XoTGJISDHrEko0yxsIYO70pzn5nnL1seI/9VwgdrU3XCeXG/4IvaeUQO8EdF
sHKGEILGupMqrztRJohz53MP0XWKrlNaM890eQUFZ4peLvrGe3gPK+Vtulvh
XRMNpCFKNgVlLYRTK0zGc+C0AxoMp71hSgPtbVc6F5da6jlh0K+ox/COkIh7
IEP1rsp8SGIv1B6E81KCFA2QaAhVZisI34ZZnf9hwPpZajp40W5t4Uzmb5om
By/v1rbgzpEwpqctFQi3+qPSGYlRjyeX6+NhSqS70tkSem/V94HD5q2V8Onv
v+PZXjLLANPKdbb21ok/XV0AtZQbgxkmfXdGwnb/Y03xDORH0uwAdE6gkw/d
Rr1AkoJeaKMc28ZGYYQD/ussfN17OgwV0qsONdOx60+9HKbjWjcOsf7R6xS3
LWdhIJj312G1dUDYRpW+6x4hLla9CtTjRlxqYsSx7cY2c3uGRnQ9qDWe8cjs
avxnbWTmh+mb/iSCyR2WQ7d6/jOeLkYyVo1LkCeeKwqeautZYZrIUblQ0CI5
x5h2D0DBcxMNzOP3sVSC0fh1xmR1Z0gZCoct0tgcvGScNtBwhLfqe/JSBwOI
042sRoH00A8BZ3EC2qNLxCg9aWvpoORQq3asSnDKKlmqJJHN8fPiUyGLXT3t
nSZmcrY5Tl6hl2URgggBNSmGVVZAzruV9jjz09uVw6oH9LouT/qARhIrVChR
AwtYaE5Cio/xYKnSVPtOrgdNj5wB1EVfNSZYQBoBnnZuoxaKxa507hdXW9CA
YF2AssMZ8JvG/IbAIpx4solZbTL8KJ6AiVyRUfyI8rbeoE/Z8slPEI8Y++4j
3Ib1cfJXad/TZPR+zpEzoFK+GEy8IORGjswEbA9/5zQIceMZ24ITpBWrzCDi
uE3rRFVa3j2x4iHPEeHCqjCfTActzw4q2aAUcwcUSVIegFpvOTkwIerDgUx5
et663pgFIsVudRiRxsz8nEuaDseOvh7DvvND6CXQ7bzy6O2BWVEE+gnXOaJt
/ZXHlua5qOSoEt5Qzt9ukSiWAbBdEN1hLr7XDerqygC7YmbIAhK8oLxnbXon
I0KITXv38hkJxXYmmqJFbRkH2ibz9ZxO5sO48omM0ZCsbcHVYxsDOwqijzwZ
S7uCDtGVXkbgI2576yXIJtdaSwEgDh3UV1recl52qZgqv8mtBv9sNl6bkP2s
9F9RMlvk4qpAxR0UaP7OFk71gYOsvSsPOI+mtasD0TBKYvejpVxwD9WQSy2l
4rwnfCSdn+4cSn7Y4azUgKDeA26YN26vgLYjmHQt/CBwTgTmOl/NwhvIEAFy
nXMBq4Zkjwm1C9lPm+UzBjsHcnBxZ2kIKeq2BJCIvYNnNqyUOoM7sDG+Ndio
iJn7f5AQL1At8fGMqAcU2ISZ5A8W8UqBoYJe6ZXGXCpezQCs06D8woPBgEjL
hSc/uFvAHRySSQdz1VcnwFx0gsq08gnUkchBJXYgnIHi4jc74oAYXveWEyhN
QrKvZkT2VMDWnXMCHuVshpy4xJBZRk07oOudGO9UYn8+M310RIQy7cjEGtLW
AnyJacIRasoYEYSxN0mPinFQFtDkYn+hvuJ0m1M5gei52op2lgxjumCl18DW
ssnzG5GoVzdiHULCs1iS71RzApe/Y1xKWOoAZiuIVuE4Cyh+r6gVKmZtn4gY
IN3jVpmxSw1OikBFkM7e5ydGELvaD3bY4n4HNPOs63yqNLMxGugOtxsVq/BL
NIcivOHpoPwbCg8zXIatfr7Rh0+ek6Nea6+RakzlV7+lN6ZrABga0Qw++h1L
3/qgrT1M3a3gc8LrCHOrdBcioaBfzhC0z8fnLWKSSayMdDxz9g84NGkt2xtK
XjbOluJxGeCYZyTlrGJeb/++C9dmDbUh3zB8L6ypKaBXJ/qo/XvOEnBys+8D
JXf/lrHr/AS039kXVQCEOKta6aYZ7BPuAPLyAp4x6WQNQg3B18ZSM5iT7SQp
GXesdvGgvj2NbIGqclrmCIv75/XyZdF425mA3kjHHid+kQOG4IXwduiudo6F
ozjeHckIQesH/EkIczVBuls5sLLqx1AH1J6Xvn2ePNWeK0Ib3IthNzWlMw2r
uvL/WUMxLrzvM+m8i0TBeTsiS8aESOFNbRYiX7vRGJq6v72iYUA1BW2mNndI
LhWG9LhCZhgVxIlZ8q5oWlIIf8EnTJs+2dTI2Tt7Wnfla5y5nq2X1Bbcxftd
pcpACIxK8nPNInNAUEOWjDxoYRyOPbWJbTf8hENnxnSg6MkmAh+GqBH7nbiJ
zaPzOceRnk02xUYFz8dN8iuG8d79jyh2IOFBz7E7Z+uVB9ToZUWI41H+xfY8
fuQKY/bZA+Dk9b6x7GUD1Zr8HkeaB5ZkIpXLMh2GK1fg6X2zNFyLAQ1V7X1r
Abaw9bnrAneqJHhf/OKQnmsqH4IOSl9iwXG7PQlVxUJwZXtAZGN3EjmmbrkI
dZNvo3DiReU4L7uHFGWAzOGSlgiYtA9JeVsGPPd4c3p/uEuAIFEyrYKjly43
r4fIHfCEqkPwAfuwKmO6wnYf/OViI77vzzJfFyWiVhgFOJSgitrxMnsK8ckS
2XCWSRmJeOzAGwfXoXOrXvMEi4SZaSw1C+xsKnZw4/BzCmQFozPCO+wxt0Sa
BnI2cIWjbgqTGiRM70UL6oDqr7qWPxYyg+F7zDtrV+DJt9C9Naa6NXlaFFTP
J/Gqu5jis/76DKM3eCrDAxJJgUpNmeZRq/5aRFC7vssYW2tOuz3NDzGwG+CQ
GpTXchY2X/yA8rr5ogzFdmm1T2IGovu99hBXkVejngkguvSTPMSIqo2+AO/n
48+CZxnW+UBUFByqSpmGzTQsfpf3szvZIbAGieAfT7yTmDROQH8rULoRBp8C
FZ7igrb/hfrN9Kbm5Ojk3kNiK7JpO3ywfxUa67EofUZ4HOrsCG1+y2Z6qsXm
txW/uudEFnMk881fqKDIkao+jkclIrFqpNnMJ+c8u+soQN3aNNXFeITdgzkp
76K3jq1lf0t0hVbvtQmWkLdLr0UwTBKQnbLIfijkYd+43go8qoD5D6PP9FWC
7qyuWqGPMMAJAMtjFfiEieddlBDcgOIcOdeXz7a5dURKiaiQVuTZB0ptynIY
1yNnyBC3tRvo0M4heU6l9ee9eexePROjL8rZkZPk2lejJ6tOR2EcVWNKQPV4
a96vKz2O++wF73ehaeGuqRj0WtRDMbbW+li4bz0Kw4r9FWnbf2NWV75c9VPY
GtHN5NA3teDf2Y86VItVuVFgGpnwYqXM2j4vGMGWIss4An9poOBY6sUslSVL
r+GTAWjfRijddqCtb4ULtR4Q9jabbLBJRp3cEcV5Ag617aFpRRSbRVN0mQ3B
yuJ65M0F31WKyjhP1AoZTwjVNF7WCS4iQbOet1x4jFaUOL2y5sO2shy/Yfw9
k5tZi9zwwTBBPNbUA5LiFFhli+yNgaN71QAFpUywPbt6hoPexDbJHMH7pG+Q
nyM8lhOjGDXny9FtxC5fjWK0tqJpCxQxeCS8IrVw6H3KYGq53fWv9j6MGOqx
yXqRwjjK0atP9GgpT85iXMuzqJb3k33ksE53k12affn1CyYALXinXJYmA8RD
qVq3rIdZil35VfC5hY965EbehH10B68xrW8maDLnLBZmnOLyuPgydBAb71i/
s1aIJdvceZzSSUFs4C/iZQ6HKHegzb/BrtZTtvHO39Qa7Hkr8e/DAkDeIXeO
oviOq0K/0eO8/pYEyrKOIxHqK3ZkDLaqoLE2iA7GFf2nIa/pH5sVVe3c90ko
ml8EvjFW77puX1R5Jq31gbX4ylNvAQV+vrNSBMS1L+hI0d4803fly+66vbnb
72TETHkUiM6ZxX8WiLw+DRAb29bEcmpgLh5F4Cr4hAOoP9C8p3dobjaRkFjT
LKukixVTmXWUtGo01nLljzaE7gogOM4dieIEN6rUb0uhacY88uQrVw7zaV2M
om0aQLRITZGi6gPF/wpoSuWVJ67TYYODP9/507SL+2PuPbJoYDXaL62DktRM
EwtbHQ16+pnhRcypE94WoxFR32CgbdLdSGQoGo/rXjUBuaDT4lh9We8zRtwW
XkOzFRQk47dDkWuWPFQ0HUG+2L8uneT7VrthIcl1QqmyzWVjzR++bHfVPpCA
rHcv5ahP5gMLol78QSAQP+YVrUMuAH44q71pZNKhPo1LZpCNrDd3YKRqYYdJ
u04TQpWAkffgKFYZk3CaiMXbBAHk1qHMxWM6KKE+3UUE8MNp54S8WrcPREqA
cQAlX4UE39Ai0aYNf85kZ6cQZQvrlbRe6JdaNDWiNclUpE1Xm6d0mA+aalir
HyzPiqLLW/Hq+1Ieg2DB0JWvM53kemvYCeEVR24zyhFsGqv6RW1U4FZxa+3+
f6FOwxGqYEkubwIfWx2JkwVLWlutEJkeH2wZ9rEfCYlnzduzMCOHVqiV3pD1
Z8DZZbHUowG+L1zKpuQXecPKsFXLGqlMb+TyShRrTTJE40EekZ6Jo0Mlwh+C
QMy5h8nV1PQSOO/DaoVkCBxEr61uQ2tz2jlKfcU12b7mgjohCltFa5fC6Bhm
JNl8U+VR8Phsvdp41VFMo8cX7ewC7cCwZVp5tc/6XsflubWwViQC192LHruc
T/MUjDPaI5ohIEAdHJPeALgtYqtDUZ5r9nLtgs8aIBis2/Uv8lXHbT2G+6Wq
sSF4EFrGGoRJVX9aWVbDr7KLFRrSYn9Lbt8xyqhylKmC29145u4T5Iss8c7t
+cJMI13GcRKXmmrcolwA7wHwK0W5b5QFkLhLzHPKTlZ62/zLCRANQF2ziI4a
G9DjHNSJR1L7D0MKx35Osd1XkgkceHTQZsR++S2hIJWwkLaFJlrRSDBTlRv8
NVs3N5DvLGD+mv2Tm79wtZ7dv3BM+CBfFqTqniocIIEd0hGp0dp/yKxTnd20
8Wvj2DK+jbPkhB++VSAYyWZ5HE4awQW3rJLQXtCDLfGpFlNSAKhGz0Lba2aV
wShAiyKnWVC4pxBnVVfgIPSJYnuskUauzhMxdhBHizKlTbtDxOda5RYTPYo1
88FhF7QK0+/VPw02lw7YKAtcu9RLDEA8TCt5tsX9Kuwd62xmZ0yU+v6Q9Ez9
hcJgFjZeTIZHBa24Obo7uuUCU5pJ1f+iLeec78Dhnmo9RIwFX1sFQCNEC6OY
3fAjqd63oVqhBzuc8hnajIiXC6KeaStS6CAlC1ZDFKb2qzYd24ko7LxH0aCj
h+zj2lAnLWJAu4yDUMlhBEEuRfQ04CuMo/N1lS5HrAYjaMNaGHeTVim7mkbL
HXGaxrc1mR1cmdR2ZgsefGVoTAdvK2j6pK3UD07DXaWjxlfSoIQ49yFQEwbl
zPp04jYqSPmxUJiHDG/ELxdRLTUcbz2slsTBVmcE5+CnOKEUXgEspLa4o3io
WRf+0Em7XquK6p/pKsRLPs5s+TwO+zjqHYC8QquCbsH9szdPWkivAmDvMT5Q
98CvPz3bhr1OzOuxCksPPpQDRkWvHWmR+RCQaUyC68zSH6VhZ7KzaGEoTooG
v8r0KJGbFmkG/vCEp74ofCR8BIMXIKZv/0MrprH/601Tqm5uaiavqZTM4ccD
2jef9rdAvWAZYpoMEOO9lDt2hRvsNpQVevIcHxaVuog/PSW1kLiZzbjYpWpc
rSWKKdVwHqqOj8DXSumsC/d7bHqRhC9rH7ewdZhTi9mpiwszjLNxcOqUakIu
ublWG6xe4cOiK4F5b6TMjOansZFuY4fDpCBrwMZv2cN3JuaFpDXG/yjXZQlf
KQlDjAVJeJDzAvTBRs8XiLwnUz34utAGXG5Rt5y1IAOAZDCUa2J4g2G8evjF
QNK6lDPHTq66OpisLezYuofTHsv5zqGFYzMpo8piOIV3ygrCx/QtFzz1rZaE
Eit76ViUBfCJjRrmUZHfs/SFr9C/h3GwAZecRbSC6LQGOKa2bkiYsZl6b73r
wPEozm06kZQ40p/vz+jwFWTQgyooUWLezDOFyWjyP9izh6ghmxCaBvfeTS2a
4oLIkr3YhTIAUPpJHLYgZwF1eRFQO7++xOBLmOegT2wR2w8r7IdrnkwPPkga
PkMrn4Y5Q/pxL07ZFxyQfQs3klCLkSBDiRT5azZ/FQuGUNEEYl0ndoUGGqwK
WUYhAysuhHtLoldWMh8ZAfjYXEkQxm7dIvq2KtwQQyMEPOtv2+52aq3GU2Wz
mkNWXGytjwAi5cReHiW9Du3WORvAwJngbGTto7Abcni63aw5/dXT3IAt+S6I
49Bdmhstpgth4+ijiGN7JcZAnNGPh9g0TNohpX5NG3mL/RdVAPqyiOB0a3Fq
nNzAc4uoJMOcltgeb32x1NpCeTmZeak7mfVUTqQ1Hb523EycTVqj1iFEJcW9
1pp934wJjZRWSuYt35fTi20off5zR18eg4LuSaV2MtfnCM9OxXCcytR7uXuz
cCAgyRDDs2OESbivxCzcrP5SPOzB2d/vbAT5fYme66m4kFUQyJqPLr/BqXHM
aWpl01v+Q3kJWJx3IzyR3o+xHhUkZT3S7AF8zcgg4ACa38GNRrck+i+czYSe
mWI222a3jYkvD7nmx4lfaXK0SBPwx4lq34BpuozJafQSxxu5yNPeaNFsRz6L
MqzMxIgB7tN93/A9+wVrlrqWeINkiV79Ob4fk4qNWIQDTfi+xFqXvr6D1Lps
zJKJwXJHZ9XWR2v4X3czys7YJ9FhpSUIP2RKmGTIVzv4Q4zcNKb1/ZNPVKW/
aAMLzOIMxmjxDXtDGt8PW55oeRLTZsPdsJ+pGW6kiD5aet5I1EU3Fa9uWK2q
79HIb/79K9OuKmFYcTBBoaW52CDYQRdtj83N6bPayalYyslx8JypsGTdGOhz
8ju2o4VVHvUsgzaLM8GK5CMpE0yROrfMl6MOxol4X+9ElZteyLn7mBsjp4gf
9wCHzTvxYqqQoo2QwNjfwV0LxDEkw64v+T3Fuh+4XG6kryrPI28facxhNR06
7QWINQyjVZEqx4XsVRSPj08I0Zewg8bGZhh4h5c6eYcqzezruCTiIqBXC6p9
LHDTm6Zd1l0f+jW3LoBzCXWNHmQNMjnFC6ckuYLstoOt2mYvOZdijHSCXX0d
SxChjUbAYNusVoyXJ5p1T6wOEl5mNal+RkvdlALcFZavWQLuQCSoR71AU9bA
6PWW6DJD71dfX7FFdmPmomzGCc7I+0szcXyxY+TogeouQ5X//fkaNuS1lOZG
/3HEs92loprEz+OGRf0M6GDSW1LHoCvK3nQTfXx781RVfZGiiE5J0Uxmr/K7
lIepNT1GbMDkmoJLBJpQtxxAezdII/w6DgI4j2m/8oVGJ8/Hg6mz+wnaRuiJ
qo5hHCizUK/ex+cGIV4QnE1NNZgSkQsydg0TCp7mjST0NflkpdJIua2t79JS
U0dWwNfb090x19WnnM0LlMwJasoQDw9I243n5IYbDH0gUUIfmRw2+8ITQU8m
yyqaLSMnwAoevISYy0jcLXry6wK+SEBzuL1ciO0L+gpJ3wxwi2gBnWqBc/I+
SWaenHDDNgfmrFY137WSp3qG5yTgBuM+h8u5mskWowcfZYTioNHAC73yWHaq
YOP7v65iiDLoIq5w1IEouSFW4+5ZJzNKuczrv9/eRKj9IjsSyDW42wKZ348z
hICPxxkeiAzu8C76Ls1+Lu1b8touX17Bjz5/Q1INxtCfa8+dPlEyQ32eceY/
KRBugw/2ZvuNrze9csHIPEfwtJj84HQxutSzpE4z+rNAHfhJZAHzdkRBdjc1
wGDO2vI03z24K2xNKGxrLaXuOaWh57s8CTeHdcUpM9o/Pe+mhYloEHgW3LaT
zNlC/gYTNS3HTggmqw9n9ijoekx72oNmzlWY3wz7uxEdNDVJJOQv5mZ7jopK
hQUS3kHTuGpX4E0RzhkjG3YakFbHRqMaLZdQ4ZSeWILpRhdWIKn0TebcIjBZ
oSQeIEDWM+fJytQtB8tRxv1kocJW+SBgjQxkJJnuG1YAwujhtyE12NPUI6Es
NlMUGgM6PFHj4Cy60cIeqax1ogVWpdOkO/IqJyt5SVQYus1IuoHQ0ZEjBkwj
u/bi/vEw1ifwmx4+TlR+rYVqqUS7Ssy5WX9PpDgwbao8Z4BuktPnr2mI3Pyq
HWoFjpVa3uRgsE7D3gULY1eQetF49Tj/Z4NGMIa9AtqPsQyGs5SAoISYrDbi
8XiFDi0a/ddcfJLAEaqeYGlUbUYjM7L7N9Ne4iHRI6HhSqnaK89GTE8KvGgU
x9KH3c9/0WF4Mhsn4C+cQ4TQdfSu+HA6QKFRF4DtZ9KWTBgfAOi5271VhwsJ
8TpkFKegsrAhXOb9H4LbDqX6Vqs5F7ZBp3t+4MPCA1OzBMVxLPK53vYr09ZQ
hPkIMviSJYJoiTv4ImVICGRUfY7M6jVv8t7EDGu0YWwRwUdBO4t7zj6Ywlb6
EdEM7ENhr57NOqj0YgOdgnsl9v2swkPR4t/Q4BYjSMdpmXplTGR8AMve45FP
LDrjuEz/DnVWewy2ESYDZL59yu3CPHAcDlN2/K5Cu07sOZmjHOT65LynaUFy
taoKIxNvXCkcqCH1WJaCSNtSfcHe9k+bP8erowUCBLlKZJj7TrA7qZpUlXao
yHQRu2lkKoMEKJaSVYNC4aKCztLjTC0loHW+7OBZYTM/W+riwDtGUI3TCjkC
vgR/zpe7WSuehmhm/IrHWwm5UECaqYFD3TP0V1ltky90CmGIKzOKPS4DzaW2
JD1vimH08a5EF7qoRXLZ9xKEvnOHMcP6BM1ElSx0Hx2UxOBVrTjTa5MV1IXK
21Q55ub6+JIE978lDl54zPopHL5xU+RwkXVXaFLH1HSG7Tl9JyDPiCkedXZd
5lc/ASTo7IwQ7cfh6Trbou1ArFu33fyzTClauhZ3oYKkEdqJOtN07mxfRws0
p9wsgq65vXb6TbGWQa6u+vaQOLzVTHksF+OF5a/tmTv/cnQOcCaBz3aUNke7
ZnUAB8zrI9sVDzq8Hcv1LxaCYHztr8nYyaCBr88MqffHn6uM5zcNq0UmWgd5
cYwQ1FuSK9l0ko/V3LradYkJFuBqKGWTLLTbGrC0CGhAcfw8V5RiJc1kGrwE
RRbmVwiiUxtrFloblN2qprvNu3AQdjL2SrV7I3Izffx31EJ2or1NLifD7VjL
HptrUiB8y5sgW+E2TfPWKVu3+0x70xmXPP6NKL9GMgjGvpQTqDlACM+C52oy
VUznknPXFyCGyfcHhKSptAIz2VRTiF1KUqEdTGpK43QXWx0zshQ5yiMEFFEX
JqIcg0xcnOgMCrb4w1N0/sc/eTG2Pl76PNTQVxv2tO1kFJ9pDY6yb2asCm9m
WNxGIk1VcAC+Uoqiu2CXQ4TqcWDq8z569s8q7DdC9KnRQ89c35eg3qnYOmHA
DKuIBgTsnh9nNj6iuPMjUOJTf9JZN/wfXboCs0dTy6MLt9RPQG/0GjHCdmev
n8aASpbd/g7B54NQnKCZedaqV+zZaXPJTmgRUlqKLY8GBG+XvuDLrfswzqjM
VvNRlNAIe0mF7xuZTSbwx3lIOQQbizKpU2RXoEiFRLHDviOIyYp1Tz8mXy5L
w4jJGJF07MByZHkJW4GCKGKec0IKIM44on/e8xADxoT/POwBY2lIBAl6vOZN
kWl478flbaIWmup69/D4NirRETM8eRGZzHsSjkYK91ukf1fTrExE7JPj4ixQ
QZbcKOipaTXXRRsMxtbmuRk0WlG1m+LDNLQYSc3rhhcb1XbUr+rWlQWwqYCd
z8KBXXS5dZSeqEOkq00+sujVruG9wWDJ79GREKOnZtANrFbjv5yDgkmT1jtc
6MYz+DmDoYJseVzapbpya9ADq0SXajWlphpmdz3FahUPn1Kpvqa+Of3aRsd1
GfDbZLDE6ch68uv/8ZrWFTRJYOOFvXwLe+GUeG4SHD3g2dp1d3WHH9iuFjCz
rtWsKO7XttuuET8NLDwDFY1Z9/iW6oHlwaCAxFlNQ4bVi3mWXhqcrl0PWoVJ
d6OgojA32rGEZLxI0HlzyZZTCVaoxJlRzoL3J7mGW+p956WkGCteb8nurnJD
MyYXtY2Z1MiUO9LKrQoiIN/Q//kauohpAYcPUHepxbAdDBSLMkyPnxlB9vYw
CphTsmYR76zytJFtzJ/PSyWQqRciqpdWCw0x2e8rjOd3Qc+RIe8HpeLJpQ9s
V5oGhe//MeV25M5rXTsKC6Tw1XxEr/MthXzbknTMiaWhyTB6ylLio2gO6xq/
NjNb1K9s2PEWE2Nhf57DTO0F9HQGzHeR0XTrw9gUYtWPPdDmrZpOqhhXQ/4h
LCAqKHafR40+jl9wB4Nwv316pVrT0WUmcT7wV366bXuPLdWYnBg6arYDSgsw
OX0gKlaAOH/24+Hvs2uDgyHEjkSkgZiwRKG1CWA24Zo6gRpwTliuMNgps78a
aghnk3dq9lbcCvVIbsMj6KrdeY63cpwZNpE08VcUfLl4wTGKPCjEhMuK3fxJ
D9R4KI0ZwVYv02H9Sguk+uFawT1C2+9x6OuiHevbD2ZcpinXBI3V/HdxEpjL
Yl4P4IEToclbGVlfXAsVeB8MWUOv+CLE7RfbH4UlQVB6UNZyl7sKjrKj3PCk
3aoWARGb0et7JQJYWGluE66vB4vt/IF2jHMic0USBsgwvNbDLFt2b6D5/Y71
tPKBfWdsAxDloBnt5S/W9L3eRtKpc+xov1n8QtjsFqeTkx/nZsvk1uQWGZ5M
rv/Hngmam5upcFLl7lvZT+wumettoT+tOnVmb646oCG8bZW18E8Ra5nEniTz
uy70bqWxLJuauKz0dujztiOT+RihzJlBgeo0wKa1gASR7pyJN8B4iybJ7mZz
WmQE9vTGLU75BMxYlxaPFUHFSKEAeknFiAHwtluRfroOKrCLpMe/WGT+alu4
oxpe5BK73K4hr5uIPmPYAiNG4QXTtDvnXMBF35KxJac7smK/7yd5HsmEH78R
3CMvOtOL8xfEv3uBgvWDmzveRtJXnJ80D/hZT1taFt6MsOw8fGtRLzdk1C6w
lQVA93PKXYb2MlX3cnspm1Ga0v1Ogdp63ZktbSvpmfUj65wa15r7ejFrZkrR
r2FQAhvsN41B0f2kPF0rWHqbQAOYrlPO/6oBEoJKhZoBIn41wQcbs+EZfQp0
JheYlFbEFvlm5dhSUzjX/xHGcpGq0YTYye2Q9VoVdRdZzVmIQxb9Z1l39vP5
4NOmPLzgupleslSzPyRuyv1CjEI8g5JloPlC9wOxqedRKE+qA/tSSFvzBVY2
qr7aXMRn15gA2TcdXwVOuCDd65vV9BOYuEoFoEY8//bnAuDSAMQuhD2iEnpK
/DPLv4g8GfgEC8hFHNrui2AlyikZbtIktQJRFpmj0/C9Q3U2SU7GpgYLVg/F
1JdbkSs0oBxstiB+qSOrHJKWopbP2D4x+rWR2fudYR/KnbjziJFsrfWxS33W
m4dAsNSUybCf4XgfXmYQZAPekWN0WexW1E+1IULl6C94a1dwdouFe0cv4nED
Sr9WUQjADpT82vYaMBnnLvX+w1ytG46Mn1AsgQQdB1GXeHrzsXxBmcFDwNso
71pK+tZEi7Y5XDSpHin9TKFOeqiz2s+mCybUJyqV//gAoeE6ll2UW2igBhyx
SlnLottnHFhISug+thOWiXflTFHMJ8QdQgEYHXK0QxtCnAn23Lt+n6lOkggs
sDqGJbDEASa8lTcjMFsVzc3t1Ul0OQlpKgq4cMrCzc2weFRNLaAFcvo5nFS7
Z21aXXxUjLz4sr9M70T0DrMofrO60u6qYE26xzFhO9iasyDY4p6J0bXJ9bZM
EmcaLDhyE8O0R4dLGYFgdkx+JGrA7nBugF8jkVaFs/TeBDbDpsTn2hxQDkSQ
rTz2qPz3ZV49VQ//FGnrOPQkVpaQ0gdBEb4UNa5p5I4Nh3iODxOe1amU4PWW
2ZZ0oPqD3X+QEC+98jE+VKvT/31MAMHZgsywAyQl8Fomi2yKHLQlc36ueBMj
EX0gRS5Fb+l2rFMWscKT11qyzPmM0c7ScDXUpQ0IChbwPAoqKBoIkAM4HfDX
1dn7y6BQZz2GVDRrzfu0qbKAnqHXPZpgVR/lL+AY1nw2zMWjEWp+ToxUF0UA
GOQrdnV9YRJ019oXqfs6maAJAr+zFDjd7Y1+3WPtcYS+b3kti01zex/r5qmw
C76Im/eV6Y9Y7NWC6/8A+rBgdFQc9WsuNczh7+B+DiVKYiEfuyd5wCch6+6R
H7X027cBg2OnD/GM/WRvIfOsma9A0FZkUyXlve9QXdULyZZS20FqTaUBmluX
S39p5E4+J8J+UIe0sg+eBZeZO5VO28Qm8cxgHAzYzu/v9trqQjzZ5Amd+Vx/
lOo6SvGhn7Rcv7XIcaB8Slwu7LBevl4pWk3SZW1QncQKf1Y42vHs/t3omfdf
TnrKcMP1NJqA8Z4ddPOFZR1+dFYCLACr3FUsB7GPlmQxEHk5i58TvYNoPVS+
sDV6aTMU4TFv1sL+k/QnrMI0f+SF2fT11VJqjWbZLfvdND4s1Q+DBHlCxB9/
jtF9u126eUypq/1Ivlgv6w+Ne1hipGTPsKiHqh+7uZL7beNhyhdW9V6AHyw9
DIMP38MO8CT7WqJ09fZyKNI09KTZ4a4s9TDR4e8Uve4DpqCAMW5soDcg9B4k
M8jhzI16GLhuOEAi2aZgfb9rIK1MEcw60Qb9vEsjvAduuGIvE6riLtmYzmFF
vqJRHclB8Xn97PDiHMkmyfBoXNZcAiawckwpzUgNYACzAJkCG8grGTkgF3ON
O1DdIrWdGnjODy73e552sBgvPkyy3Aas/aIeG5tlR6mihTKHXGYqo6U3BzEK
oI4tcQa66e7OojizJWKI6NwGulWuw6jyWLA/B6xxul5uJzbM3q9OiA9kArdO
DoQC4x5hOUuqjEPz78IsGQ9WMQg+dGz2uytJus2Hp2rTH7pT8pk5uR85rCuE
P9258XLV6qIGCbxDKkCjTK6mgtod08uo1y/MUChQE4f3z6eMr/Oij//D4HN5
QrvEVn4MNuqlVk/pjPXdrvBkLAXotsgxHbxgStBbEhljOwC0hMZy7Nelm5pq
hNlZnRwKd+POfLqE8yOtFK9W/Lj2gPjYET8aId7C32oi8eTZ/NbOxDJ1YVmm
/wLplpukGa+BOK+aovuAfCieVjJQfUvkUmR0aqzLunICfWfmJ1XmyEk/KGiY
6JAYlO/LEscEVmVE1A6U+b2xDq7TKmQfGctkmbKPNxqyrbbbrHYbZ5fHehWm
Goe89wjSVsye4uDQJtTWybvt8c8zhzCjVgKMwxkW1AM8E1uIMQyXFbwlx1U+
VaYVk802IKo03Qt5yjEHNCXVecuKdVtMmdj4OshowhqSZz9c7SyoYoInNUKD
TssZnhqVennAEtYPmR+EMPL2dBTZvJd1MVnOHYIBWBgYLoEOIi053tx40vOH
FJXemXyPu2f5tkLtHG+vPLWgvR0hEnsbRTUhXxGvOVMLAj0t4KNSS7PygD5A
SZ+7p2DBXRDzB0+CEAs6NfQPUqdmCPRtEEnvjeI9YyogJSWslpixH6aOShfe
bXWHSfUSHNbz8k/VpxMQjVWzXkntFvHCFjX3Utb83A+LGzdHA57Y7knu6FVo
6GPVZGG5/W/HgqT45KzLZke+7c4UfjltKpopG5u9TBg3nWpvvpwKL9sE9JPA
zNDpUNrYdnE9km4Nsz12+Ts/BZEMTjwdbP1h1gto5vpfcJNU77+/BbQ1ORlo
5ufWKSIl+waFGWohwCGh22TKtvZcb8LlHEwKJOl9rh9TatUwAo5j2dhFx/0O
BAyDWdnLT57/5BLciBSARWchK2SE7L6MI8PuJdr1hWtKva9EQeKIadcobzUQ
vxXs4qPRA5uCQwPyJ7runcjbcc+WEOmURpIXTufogSOHRkRUUma+oFg9zqN3
h9IVZsScFE2ZkOkBPKW4pTPz4hJtZG2Oxy3VEN0v4PmlgD2jTqLSkp1KdG9L
W2NqpPFlkUpjKfTXrv/ve+9cuWj7EWl0QdHuPj0MESEkFhYKF/hCusYrwKc4
S8IQ8jaXMSEnyDlAfcEXlQcKRATxfNCQCNbbmGhTcdPxYEpra8b+AU+Vh7LN
i+9Cz9+QnfIJxcYVGti5AowkhqwsHto9Hnj67RVaC06jaA5O3e/EO4/dwLsu
+EV5qrq1LavF15ZL85B4W9eGj1k0Qa6PRuVn4yJuTZiLjMxBmbB60Td2ZENX
Xy/uT6hrPiTC1rqOXSG0CYbzV3zvkWax1MwA3XCND0khsdBJ0Wxrdaiqa79E
G/6XlCutBhr0jaI9gUsqTMUXN9PDSuZJe0qlHSgkLvtjDS0gPU7dXx9IjtSx
KB4UXMhsxIpVtkhN8kNQKLhhrFNr49TZyl7oQ/abBQKuMsZop0tRiXoHLhZ4
Arha6QJg8cvJQbEcGnoWOyx43ppwTz4tskWhfWRIpJT5Uqxr83GkXOVMveg4
sJVsvWMOjmdtcOZFd/jU//MCr+NSLX3DI2WfAdF2tbEeZ4mlJ4tEshFo4N+l
rLocOhP40DlW+xYKaE2qyAHlSrcxdMvV3L1Euot3K8TS6ik5ho4Z9IHHRa+p
UCZT392fYNPGQXLc697248Ay48tuLicERrHdzxTuAKg++6AzjQ+3bFZE1QbX
D8q0hbC7LVYWJ84DCAapTovDl//2a7W0v9r3lmeM8R1eYtLIqKdp3kmCHwz5
terJgrfuxqV5IaA1S39D1oppCsiTMcNhwQKKitUug8y6IrWDBQqJ+vESZTjg
gG4NtHl0JzfbEe/VAM6jwxi728DgsmNuBekRFneC3oQSIiZpk1yOa494X3PI
CDzVpCQKqr/ilQSxE1Eb9HTvl1gHqQsYNH4Qhg85MaW2k/BK8DZ2UpY8NFuK
y5hFZHvmtU2y0TPY3qqxjEj9cuVLCLzfS7D31k9ED92yplYTbd0Bi34RMYmO
KK8OHolW1Kc8c4ZEZD2ssY8NGsByzgT/OoOk9hoXyf5wzv1/Pa6xhGpTko5d
J/Ub0HDc6Q75niKAQuk0/ozH24c1m3tz/HZa+ZJ8JJHXHnJHI0krkj0WU4Zc
ZCRYRjn+EQdMAVGPCLk3pw6A6ecgWjHE5FAM2aTmTbAOr6FbZ8fEYx6wVDMT
xGbzbmLfDtGbNELLYszZXqQMuOwnc33AAKxQwdSt2kA+tt/nhApE7Ah2YtS/
LzUgKtciA6QWlD1/0x0N/uS5DOD8s37iKLZOPup1OpsgkuusObAxZLew1TSf
UlWavzUu1hqg4rFADfdObvvuZ83cpd3IAMTwPY7PYYSurkIjig4UB9MSt0RT
ZYgKEls7JS4S/z6cpmFUznXHMDh0Akalc/eODZ9JcF8l3QiII3WtaE7GwAqB
Cg4RutNIULaF3/LTzuPelCTXcPOeKLPsvpqmmO/hrZZNRCbwj34AfGNEZXYC
JJs+W/34cEiAhPRcB8LFMoUQZBeHlwZ/WNoIb+cUuMTY8tQLOuxAZ+iKJeni
oMFZJQeLdDfaAc/m+i3P1bfYVFWaSovn2+yor5xnyU1VnVNsXG87vpkTcuIN
IUaWWr3utn718kUsBTcfznnY9Qk7Z1JOkoZw20dHuBjNHPMSq96jnLUj9sGA
bQ3KRbJjH/m0D112o2Xh3XyncqqxCeGyzVbvlrkGKmjmvv8aD/4fxYSWaMec
0qUcVka3eFq3xOuRBTH1/f6wjeRMR73segSzt5+ilhg7SzHPUovzSWzrR17F
CTAoV8hjTq84bSsY4+dyBl6CVHaMiAx2duUexhnfse+jnDeoQLEmzkEqRddi
BuGZU6IY4KIrlsC5IRj4Uf151Hj02rji9zVpN3CwYTgPCV0yYfw18tLfKfCA
11gRjryZYdfkn81UkrZZofW9S1zIIdPQPfwSxkATms9Ynf2gNkTGQzPSSAL2
PKTJD8L6K4NG2uUNgfxn2DwdI57Tr3HEI/815Dpz6EsqJxhtSmd+pYd1JgV8
ldmknV38FnvFKpML2lo+U+PZvBjyzu5EIXtFP8K1J5admtTwwLql59wJMJJE
3NoUgmF9vmBpyLgxNz4bjQdv/j3BJoCcGkzW5OjMF6zR77Rz2a9DFmFuSyWO
cGgrVRRyBDLuRRRS5p7WVo55POn3mMYGTfSX2sZC94zqu/1Tsl+xGEsnETfj
ZvoeLRksH/6x8Mi4nuEbvcIdD++BHqPhOcebKCW14bxSi93UFCvsCc4wFRth
OkCp8tbjwNP6ec50IE+ZKQAIuGhopqrtNdByM9UHXNl5cKgQ5KlQ43T0fEeF
DJsYGmUveA+0cxUR3pZIhuwtARxq759ms6qs+YOJtrk4mUvbrS3JQiWUbyke
c/a7A/uBFlOhtl8mfqsx2ErzITbGrfgdrDf+J//UGfeKPPI1rt3lQIXSQRAy
VEjH5UHDMi/8+o3Z4GA/JPZoztfAOMpUrbCqpGzsBeBLAbnoQYNRyTJiE+gr
iHef/C1xCMhBYFrHfSyWwWFk4YgfFZKadem4r6fxQ3eHFQBXMj5SEy0AufWO
xiQLtztvj89PCEFf+NbpddP5y7l4I8RargkOS+YabyT4OkT5/rmoAjqpRLRh
31yKnYrhQZc2bj7sY2d5e2A9g4foTT/OoWeWbKZi/ip9u247WRc7LhUhSoYz
5kpZIXdeKS/AhqS6Q9Qc4EdNHX4Ya7zxQ8GeVJ6eXEnptTBLXVlu5IC2MJuD
+zXlFAL9MngXWX4u8JdRaH72yzFraxAPkWVlUUCkbPWJdeGcRHP49yG2R7QY
w6fpZf3V2W/3bXVWG52laeMDYKh7xbK73C4iBs0U2EW9fXgvAGTji0gDOW/h
24OaH8T7Ua+rDEA5DtqFlW+6HcP49jwzK7lD5OAuHrWUlF6kM8aOj/q24Ijn
Cqj5FeIGdjp9uQVdle7j4I39UE5t8vmTqaaiEzmjoj2EOZA5Me1UsLrT0+qs
il1/9eGmvzdKbGzAiWRnBpgGi0bVzygEPOS4ho11JV+Z5RDAikNJ1KIA9k3W
eOWonFqmODfrkBJutx+a1FssWbW6cy7QaCk1NXQfE9+ZJ/5VcjrmCQFFjqYw
l9ckv9cKB/dkK4PCCFQ7iO69wE/7LNbIaYhVDslG5UEcw8qx7Qb4v+J1borV
Q4w9vwXQ1b9hUgi0zTfxVoF1lwTYxYSurTu1sXcRxvOUr8NU/U07iJFlyFvX
23fvU06j/HLCxW7CfLfeRg5p1AGp5zr8g3JF7Z2zQkV2h+Fgk6bMqERsLAV4
qYw5FWxY+iRQFE3zn8OwA0YTVBxNEnauVkafTAG/U2JxAm6GIHSwxhp943Tq
CtDkyE2bHfkJM01pkdUEBXMlYEXTerIGpczZuoeo0ad3wHbxZeKybClTY1VZ
GtKrjUUyvTOAjqeeQzsy/Y2/rhfnWtB+Kezpe6aQq75nc7udIAhxNtoTIS0i
uhUvX5i6GmRRafBlE+8rHHbOUs/pKh9jzYrBZ2qqkkbQTq3rCZq52DiY5tdO
4cJscYOJVvH3Idbx4BoEJRsBycN+6PG3b8W+PCCKi7MYO2OE5MiB7/sOM9/r
FUQUfnWa5C79+o6ilxJMyj8LhrlieBr6njyVC8SyatOnG0SF0Cjc+zVJXc0t
t936xejA6dHWmX/YZXv2uIatArijPgP/9IKOZo1uWacK52+nPlldgxbBkvZT
mLYiVoRpNTm6JG7/FJCy4xRLNN08U95Y1vA4L5njEF7gliOTHLcF8TcENaJn
C0RnnfBq/plzyNGRMhIvEv9v1DxO63mp/SdJ1bRhqptP1j73baFPNaVFzItY
DmmxVZ6RvD/RCjrLkfTYFKRz7uLcyH5FyDjqnUZZ+teJSBODao4JEJjH9+RM
W8mPGA3lHUBvt1KYuKBFoodWfeZN/sc0XglWxV8mWuCUggOcDvbpzIvea+ak
a2NfKe3Fmvvn2+bKKzbHBe4vJjeEgzOy4k7+qzJ/yzNC2XGc08gIKNMpMSU4
fqZyOPrtijnjjruiMhGAz5w+JLhrBkkUOWdQ5Nc8+v2mjKHe3Skx9dXstd0e
4Duy3QCFqzUAKJuHRZb4vTr55qE674KUoFMLMY6z0NWSiTOO78ehgN9dUE1A
N6J+m5cCHkhQYOOv5HdA7Td8JaaEdCrbSXSH0U93sJwr7pKVTgc6Kof+JIeq
Xa1wRPCY1uGLBLp5khzS/yS+N2gtMt13rY4IAm/o44zprY3bP5Uc1lLjXCxC
mRGx0LnKnYLl/gcp6KRHOMFEIvCgR1X74Xjdt/bTSlCsFa2+iMnIb99S9iu1
RBYp9ADF1tWaFkxyon2YGM0oDm7d1M/ub1rObPKHqgU7n7JgjcP6g5t56HRV
DTT3ME7jh6WwhQBvmb+b0tKKxu4IU+jvSApJsTNwALNA9VUrI9VACJT/3kxx
SJWe6mswTwjPXder3fnHQxUcaX+34E+a1jvJXH0xNBPy0E3loyL5YZtC5eZj
Kw6zkbP9uIA6DOLZLdaJbE75jOXxf5NzjRmohdfqFDokHrbXJx2UwPK4F8PN
uf6Ea59r2cqWA796Tep370m/+noKSbgvfoY1zjob/dJmqYa9aiVBSwMHzJvG
a2oGmwdTTb92uG9xFcIWIS4toHEpNhipBJdxczU/tzuGRQSwqVlFuyaFdR13
a8s3ouJiEKfTclHTwH+RsxSrlfpL4+6mUruTSDqwCEa12cpAorqHDI+IhTeI
usZp9bQ0mo+W9VWfeKR3SbAuTe4G6orWn8AJGgIt6c7bnXo5szUlDqA4VWsA
8In7VO5M8wIUAWi5hR25Sq2NkYI1bopIDzH/HwWAqFHuvSGtgV9eagoLF1oQ
RzvAqVYM6o8Fh5kBEB7Pv2Ebf5vczLwmQ0NqsVcjfRQORy2Baegf1xByCLcm
jZsU9IQTYrfDSaGVU1S/jvaordtG8EqXaofyk6v9/Qi9/DTH+Ce2Zb5TXJsz
yFYlj7sujrzVP9AHvz4O5zrjIZHqiI1vASWpr2bx7aXUQgbMMI7S3rRGdBTy
gvwuY59X7ydK5K9WJYy+Uyb3nkPjMVmzsnlZcf7wD8EfT5dYV8RKqP+vITq0
/FzsQnepMlWlNzwa0n4EEpM92Mpy0j09hL/K2VEfrSJhRO+PYCo0MgD4bMCM
FoklDxWDFQhhDx38DwFmUozlrsrenSodUUr4NfKA85Vc0t+Cx6J5Kcy/d3tg
Ob3Ovd+pKzdW4mA0AuMhGtc9G/yPBk5LHUCiKIa0NC5E8EpJCJ+3aPhleyRD
2Z2nOKGwTySnt4YmGn1QU1EScD+GIaYHd0va5qlKx+dqSQZq2OBx3cDo3KNH
OA6e6n1wOMtN5s8DLzgJDbP1Ab/LA1oWQjSGQPSzKNlGk6X9xiMw+w/ouIny
pmZAx2WArhvUb13c12XtzM3/y47PCFODO9wd1qgJB7n5UKuUHdC2BASXvmeo
ULP7OqXd6HhC/RCaUDEIRwwzuPR4yEUySI97tddeuwphb1rJnZWMJfLzu6D3
MWoY7pm8RUKSGaNTXga7PFNGD7cQxj8WJ9j4ONOThLfKDKEIYzAJZS+XKIlt
4SeHYhHX38Nk8/PNeBOroCpBvmBFX2HakQhykIm5ql0JEQT5QtrwprXpGfXP
ueC3DQEdEm7JeoxEdQPshdzH0Wkx3W07PuBqbq2PGzT4HM0SpkpeKmw3qgKI
jbKyQiUbTX+qeZf43DqzxlhP3ejgkBe1fmaPTYggwlxzCpNhOU5gIYrZt31i
k6rJ0K/EWVEHwWZ8PaVq1BNFT39TGTHWRKIweMq4gGSQWe5PlB9r5gXH/yY9
Lxbsj0H2YaonksBMZigPhvQq9+i+LlTSrExVOl2V6so0DkwuNiXRWvSId7EW
4Ga3Et2Fj2015Tyju/ojlURCwnmGKHpLUnB2m7fMzafMa76/B1cqGqHnLdTK
RmWBHaNLqTXyk3krJdANfHR2k23mtuu7xrjjac0g/dR1sgbqwkxPigM7vVyy
VFstDAliiiLo+uf6CbE0ayI9TOLHao11xYZsPiM5PpCMmy0Y9sMCJjg/Y4o/
ahpvU7iXBjUkcp6puyI8RmHKB8U0ZVwxA29/VKrqjij6dNf50ER3OdFg0lKx
bBwd+ghnOYMZrLIaeCO4Pp4+NmhYbWy40nVBjoSwefCpkyzj7ONn5Q2UHAEP
WWFeWMyR8UJRd46zoyXO4JkMNjfpjNqwasfMYbwrMBirhM5t+G+VvvUni6CZ
3Ug16GdilB893jXeWk4HOXB7wN+6GLgWaGU+Ts+lX6qq6GrRTYofK3QWTN9H
XjssUGEgUlj19eXY/OsbXNjb0TJASFP6PAUFyUE0LFNdbVI50xZanCm5PFTb
e+VJCiYBahgv4QYVwx0Ju6s+BKr2guHG1CajdF/JnB0+tVQhapCZ2uDLovxF
HpE0vjhY+tUcAGqadJI03XnLLSE9uGbMuUK3p1SxK+bG4u9BK72YSoIS+gzW
IAt5na/UZy3U58484uzUAOVKm7v03LRIz2vhSaxzDiIoY1hvGDgCYlTKdSRu
+mhaJ/UKY2+GZthzpU6XNyWtFFNxgTvDMwXeehfn3rV4Bbt+Xp8EL/q6xYxn
kwYjl/rDFwAk5bHQgYHDzDf1E9+HvVur0Fe+i2o/6yNzJfNhqG2cAEvyGFqH
8e9tFxA10DYBTiW2gsN+35FN6g7LIrdSeXk5CzFJade98ofoEjjPRVUir2QG
0Nri75Lolibgn7E+Pp2TRHNAK1fvA7Je1ka7wLukY2750RPJL0H8q+5NCr1k
fRe7ysi8xmb5s8z62edG7Dk32GFwciajbb9kSyOYiukBlqu+CKWdekMhSuez
dI631lgkn8/iCatLkmTcyWcd8PwTXMRQvwK/vXmnDwG62kZCkhXqnCUVmnzj
j+Tzq3ItDvksYRJKv8nVKRr4UVuUx3jFiOZiMtY6oFjL72t5P6O89CxpHb35
+mWdC3KgAAE55j8ulNA0yTgYHB60p9R327ouLiX4o0RlkdolOYVoTuozTk4f
10cKlVOLpEoFywx/by+cG9Pi7OxTQust5p8WNKLh7Fnw2CcerMH7YG3h2mS1
K88V0R4Xcee0EBmMhd5fbKKkkSB/rrGCc6Jv8wCwCs/bo9GY+yjQnRMWdC2U
Uo05Bm3dSMJvhFIDNdbV+klaI2yr3XnFyqfKjJd7NUKKFJpR7IfZOeg1mkVv
E8bsyoC1RifmVQS3vPV6dCdfiafsjMmqCwIl+ONbDeR6+na6IkmpXFMG69hR
4lxMe7ohyzaespVrE9pv9+6pFRu+IETvS/U4e87J6HxRN8R18t8fuXB0yH2q
72s9cvZJeJROwFDgu+in0Rifv2w4cMtHOm2FJUvc/bNH5Ux2z/bT8gAPFTdz
BtIVqUbhnP6ezIqKLc0Cp4Rb1eHvSBeVV0gSfY1k7EcP5yeSSjqYpgw0l1fD
jOPOzTDCzqeCAE6EoXzobKYHBMe2VJwUviFjAZ6JpFuBm7Bpwl7T8S9TXcei
0BfttBjpRMFuTsDPiHlYT+d0daPiR90BV7A4qNIzCkCnbN6MyNTF8Krzt4ZK
UJvN/Q80ZoEuE1+dzO8SpWo6GUoYN0tf7gZ0rwlzmsCYF7LadBnHu4pGXPRg
XMshuIqwHWkRqgm61LkhVMwNQI1sbfAs+3zEdH1mZmjtHeC4H1jQWzhOIoqI
kb8lEqnr8P2xZ34jL1+haE3IEvYm3nrnLo5iZr4StT8NFkr0q7DMDqnbfLKx
8mpEQvC8Eg1Lvj9LURptNY+AGIszLP4oASc4j7r71mF/yRbq9cMIVmPVkujN
o7xleJXS4dHTzk9n669+snIeAkbPq7WvtQ7RypBvl0HT0nl5HebPyoZwD1nr
z1uilQFTsITc0bg3/8oP7+H7CSBg+E/nizrwt0x/RUzDpLOg3MQ6KuNd/rtZ
ajMnlUjtQ23UQHGdXLXiRd4seGlQjiliQst3qGeoXmBanjpgiBCrG9SkCKCw
hHLgmCX2sbMFBfJbmvhMv8ko04fy3jNm85FLI1EDL4OM56lUpQ9UDHyB0YwI
L+t5Fstlz+wUBoGylJvInylPf8o9bVdp6jiH7+gp7nRkVpywEoIiJ1cpOc58
ncPWs6soDdIVd3hrHs3hTkZp7TAZMzM4Q5WFfAVeQGF77rg8KC2xugdM65nk
MZv2qjbWoWgx4p8FOl26Jf6M3EyEHi9mK6vQbOx9puJn/yqTm0bsf/2l9qRu
SL1N2OY+UlIkw96JwbUGOwfep/nNLVqHAySav73amJtWdPSSDVkZJv5QxEL1
rh6Hg6eLEYbvCKoj+XpYrGg560ly3oSN64OtjHGDuXvaNBf5sB+aTElGLlVK
qPhhaCGq0T2O74JbVLURLleo8JfWjPR4Vqeb0dnhkqZI6MVoDA2X6ub5j6pv
YAS5EGOLfQUgTPvenEyOai4lGiEe2/wMX7I0kwx4lPWrY98BXVxnnxBWtccQ
J0+pHc7qnEHGdRX/rYIkcwUGVMCMswEnjEqcWi+WY7HzLtXBHKEimHss1aYl
q4/QkIisEAnUF+LpsIQhTUVN2BcQMUK8mzCITNoihPzY76yFcn4RY8VSV5yK
zKiFp66iRF+T69dgYGaREmn6z4ADj2pRTswIeuxLjKhtSU09LJfmOARezOSJ
+TFeqk8niwJRHXcZjDFQM+0avJNxAOgPeZ+OqHFpnAVZt5C/IxvhsZDVqX7o
17dKWFu/tZC12oPj9BcaL8iEZiSYerab1Wl4rqIDYIqsfsUL30dQnRcnJhZv
rw7cKz45nq8jxJaGT8x8so+Ih8wAeRMvYsLtsDy9XRdzK1YQQQu71kEh0I88
IJrJtKMSn6AjaH9TyGNEt5VgC3DxmbkekH+ty/M/chrrCcdWBzlQ3e/FOuUD
IvvP/NxijtNZ9FYt2vSP8dwnpTPGuEsQ39g4Tyg3efXPSMcWiGNhrOp0DxAT
ky44Y50ZmtsM7CnY5SJLba0JTHDtZ0Zl14is+N+CFdTQgEyxjlDkgAJBnwne
r3u/zpahQ4HK7UREkYjXFHNe3yw/HHwnj3fDg3gl2Xxf7VXiRfsLjR68rGey
aJlN2uUZxkslVqfi8Kr1V3Snp1RJXVw7N1M9XBH6K7D21h7QTVxIGrfp6l7q
5djiXsOP81tHLbnTGfyHLIK2oLsoQhJh2z/trR9gjCxSIK+6Jtc1w2XT28XR
052qrIUHgEgmfxJPCOpFZ+iJqYSMXm6u+zY/e6U42oLZMqKGNLoyjQF2Ctuq
UqH/FnKarmuMVztIeNGkWBTbBChebkpDYNOJxr5SylcIRy8gSuBWjIrAX89d
CoZ3UUTDI+n/HcGY49C47DmOMxT73xT0qtvAJYQjZKVfyU2Mue7ZWI2+BVU/
WVDACZ6LnX5pWvPfHC5Modg2uaCnvjP5mOlvLeecTjXHdIh1259ECx39UgMc
5zA7u0ZY3f1F/2jPYjW4D5S9Tz7WjusAadVtmaV1OMVdiUtuVWXOFxM1RIeY
IIBKTbEiHH0Q8Dtxm3EsiG2IX7vqOp/HkTEm8aHEcw8eoAxvHhaFzy11fZCj
vWxif0tickYRvDkR3+eo+Io0vtuRDYIckr1RvaEcbDlx8XGc95CcdP3n+gVx
Ub8piWeick1NSTiQ91RSkDVEEv2ycQ1baSZ2r9xsSd4Qkml3j4sRoSOoWLHL
aXKcSw8u1abv3K3tLEyT305EK3bM0Y7FVZsp7vYyJgvIgNLLTyCEkEygWTam
L+KWA2g3W7dfmzTdY+zeKw3gQeiPOr3tz3wabMQ0KiqmfwcIxckmnqblDLwa
RF1OZqXbb2OeYgteG/MKstMDYoFXji4qlgXhP4saaQeDz2WsLVlKJvvtyaE0
+mf9XHRv6cFSaV6EKnOkC117o6YoHqRnhZ9RhRpNxRyy7CBLA4fzgTVm2usC
Lamse3b3Uh5tUumXeXsMq4vcI4ylYAAxToYRyxPLJ4Zl4CYOaiwCLuiguOFN
JF1D5fQ2FfEWYmmhRS20CcfBhsRC/l/xpWGZwUs8v7xfDsSFlCru1xHvEFuM
b43fekxNYLnWNdF/ke0QohzAtPgwu3avQTF7i7d/BVH+fLULHbeqaHG25NTt
pIkbZ3SwFA9J8zFSCplesadII8CwioLfB6XVBAiDgd6ExCVMFEJdGOlITdMY
YdWzj7eHUTu8RtA4M8fzxZQ4HNNi/5sRoI0aHkZoTK6S6zzuwFl0u87E6m5z
Ne6VkL5i3hptLMZ1Is4GPS57sdjgLB9YRONrFykx13H86tWTun/66h/pSpK3
efPJGBRWEVuhrR3d7zZELSCjXJYXnIxi9NwucFiPwexvSQTXfhgCooGkMZgt
7YCOD1ZxEuQ4SOCpN56YDeulyTDqi5/+Rx0c4qeg2gAOYX+pPofpZwYi13R6
/6PGoeQr9QK3XHWhp3UG4flRN9Ct8wgt1c9UeiWGarv5jAvyCAAPzkdjBbBl
LKWz9F7Vx6hzRwg8hb7REu9nhvgqqPHALXePNrYbrj19lRDzgEWPuPsW025w
0wFW9Br5cg+WvL/GMgBLYNU62heEDXUYlSz8s3TkoopgBj6Pq6MmB4Nb3Qh+
+UTJpQQZr7xNxb65VsilTa36/DQ5SuhqZ4Prx+QAS5zlqxq7XwOiZ3oD7hRt
qKWbkwsjGIFh21Jq8D3bIcE4PSAYM9SLQiTGVMPTL2Vgn5J2mmeHimy5hCXU
/4nQ3MKrBL17Znix001trV91jR5FDm7ly+vbS1l7Q8dx4g+xA/KXvToL1uMj
7QbzfQoMCx2OY36iri5Z5hL0laxCzZ5M718EEb4TH2nJc0TbYwVgU7ANOBrX
1OD4I4rlMlFKEphqQFZasHECg+bXmtHKghtyJNN2fNgTOrd0NIKQlycsuOqT
M9DOO/b/n6A+nkskquGAcqlZepb7dliYXcV1ZiaeMHS1qFrSGV2cy0sCCuIY
P51Shp+Ewe8V2VpOi8qXKzChy3C1Tq8Km4RN5gxbvRGFUHJ1XVn6cTet/EP+
TclDJdEdA/tTf/2fqmBCmLwZ13aC5ZRvwGtjl7aG2ViVukjcvvcHRRo/ia5a
MjWgybFG50mecavwEWEvJ4uv2jXeN1+96PZwH+Fc6SjvMhK+ZGjDH/em7a7I
l97RBq28IY4J1pTQqC7dEhhtdwKKaRWvD4G8l3N14VOkEzeSAnponwyIQjRh
SDV6i/fGSWU45VWmqs7yo01fbGA+fK9SOLM/Hrmzc0ZVQDeVMYycHaCiFunD
PqWFY/CbIhDbJOPV0OtwDFw4bU3/Jgnd7LhYQ96BOJLDWb+25465kY8qjMeO
UA6bf6AmP6hJONVxBcA/Z7hr1j/xqSPQbsgolR2Z9FapEn+WyQqglDpXX2Cy
vq0+OvRjpMHfbjF3OsH7zDriag3Bxe/Gg2rYQWSmlqpodEpURQdJG1XlwkV3
2QujMAJ+d8l1zQqzYH9jRBUNl7sauzucIO+vkYEFugrs4oRHoe8NqzsYWV9W
8AQELfSjlozhqFu5FRJFJJCH6ETUaosyy0e7gXs2Y5fCCGjxZDC5ge2zYSZt
vPkWF+OIQzytBuH+f+IVfUs4Mc0JXYjK9agouU4MqpGEkgRgbuGOIn8BLYLn
TDRW/k4iAYJi9htzN+IJz28jCfMUTdThgJREJI9GqOFAsI2bt9tLmJ5YkbOC
aD0iCqRfmqfs756Mj7uU4GlSj+Po2VfaLTg6QVcQ/P2k16RmK4honZ7RI9i5
RVQwUFOEmMu0PBbdXHK2RNDFCiJ0n8BX9pl94hJK3ccc61BsaFov5GqkIGzw
/AkUiBFhx1r1vI4vH/lktL++GAaYCtRvCCo04dav9JCsjU8vytVE5hOFT/BK
/0hMCPA8hafqmAOMJDWeU+dDjxUozpXB6lTrevyROY4LuVXEPuIIxbAk+Owy
YB/4+usmzDyZbYB4R34vB6SR7V+qwtbY8c91yFgYnCe7pEALX0aPu53osWoy
0N3sMUqN8z58tnxGMaBBEOUWkU1bON5pjfmNLlS1GEKbHRy2Ph1Z5h2FvoJU
w6C5cMfKX1KdjRTDg/IVOAD1N48xBdU6emCOnJNw7ZCuUbOIz6At2YnVIKPP
GkruRF1OV9rkaFKBE4efgyAaaTdM3oCnWUTP+OLLqyhwwDEq6ldi4G+K4orF
MUFwm1o6GByhq4Tal3YQI8vpQ0Mez9kT/PIWjWlrG+i+K4ZpOpPVjba96H1d
dK83b1ZHcqwXN4zTb/DKiVTstMwL4JgC5eGHfp6qSjBLZHavsY/A4WL7xKml
TQMxnFNodiiAcobtzsaA0EiJBLVN5XdhKJ6X4Yf7IB9QRNizsxYiMkcKSfn9
GlgEMDt4kTkQKxGx5lrduq3p+7e073AacZ68hkJPeV2FULGYuQsQuO2k85vG
ZJ6yeDlCSObBEEfD2a3uWK9xpsRhfJckWjIWqX7HrIxrC70Qc6kpFC5PMlZ5
8lgv75ScJhjlswuxB+EYBgoo8C2zSQFXTfw7T36vUTCdBC6aTHcVeE2li0gz
tBAwSXS+VCS8X4r34dZI3ezEuO5FliCb0ZIP+h44FB8zy/yqi4FndnMqC1lZ
vXu9MiqQaB4Aqc9W04OCgH6acZ9apQ0dwqUmBP13iU0wE1o0vC7sQeNC1CBQ
1hSyu6tvCA9XUMI8raBTYAx9YOW0GOXiU/XnD89fvL6sZdMXDtX3oKUBTDB1
1wKV6Btz5S+os8yyFlA7FSWnpWGQJcF7mkLPM+kSt72m63dOPDIHsqhvIreB
DzCScdKF++UFbIGDGoy9CetQSTZtM0SMqOYLaLaJXJ4VO6R/e8kyVkeJkg5D
ks02P60O3x5NwXrAjIfH06N0D8s2EVUM37zwNEwbIprOUARsA2Z0F3b3OnI5
twJ2yoZVpHomgYywonEeS/oRjlKo9CxiPw117z2MH6QUEJ/KynFNTi6Xt/w+
4K1yze/RMEOp6Ret7rA/esxXlcaNPW+IIG7iarHl9imKfzwXFC3Sn9ug8rhz
v3AII44gPaRaXJajr1KhvrGS24bzrz3wHEpOTdqHRZwpG1BsyRgxFwAwipEI
XhkX8Sll92SP/NXoB1P0+9TpzJwGe5hXpvRLXmktusyQQnJ/ex3R5zlr41hD
HmvSEBDc033cmcO27KnaNb4la40MJ1Jqai3UsMATCXtctOrrPr1iuF6tOtBi
G7PrnqzLFEjTJiWiuZAhCOqclDGxuN9/gAQaAOQBZ63GpWlV2/6tm8fNe7NT
WyTvOIlYVcLtvEiiK7Fgn2M8cALfdoS4eM+4in2+VHRXInB01E6LrlJ63g8c
ASc/iljBEdRaX+O/vo8wb7vbq9fiMJ8DRmJ1BnsukvGEnvFUon68L2JdWCxN
cEgRubYjHqRUjJZkZz4wpV72ousK50rffg8yaxxzADtfM1j8EtRoOcrscuGV
hrN0oP3/9Hve+eK+SAmrgJSTWklokgpBHh2uvikWVORqfGOc8mVm8XJB13JU
Uf4D+A2MEDbf3EmGmk6W6cONhIn9kz+aJnv8WvMc15oubKkQaQV3KrPk+SwY
RyNg6VWSNywQMZkV4DO5f8AaAcZicdNBTOXzeT8Kp3LvX1XyDwDBMF4jXahD
T3QIoiK3D6Eyu7ZvR4evJN8MbAJeFZGcIHGctZQZhaPwwnRGlR5b6zmYiJPk
WCxziG0zu7VtaMdIAAf94SX86tAnfeWvvVXITHZwkt3d/xMXzztY047w0f2B
l4j81IaqNXGlp5njJ+vH0EIMYfd7Es5SwoxK14lyg2jpJyHZ1w5NmE9qAfsf
/ig3IsM2EXmoTm4Hwbps4tjs3SHM1G13GNHXEA2py8HHHbkbgBIsm9tbdvle
Kc36lXDzF0GOPrSTc7xSt1diOW7iLfjD/nv+33LLBr4vgfMISCykpx6qmLp1
Ja3WGYs9O2/HInDHmX7bqJPV0Bp2Y2Xh6cg+XXVvrRx02MeV9KJBRfMt0DHd
ct4sI748DQEHLaCPXICjIY7dEApjyHBCHWUE9J7A5CCZWG9HVnQE5jwQBu8l
tq8P+v48aaSOk0gR8P5e2Hd+SAu/WVctHNKJjC3/iU7Vq/vzmI/NUXPfQJZK
DIe7J39ko5ik9OJyWpMk+wlMlj6QwjPXMERBKSmIXXXr6AH46+E8rFTqhHZP
NixlYsSJ/73ci08BlxjmicyAg3XhtXAFdxRYDZyQLW8w9ezab3jNavyZvjsE
QpDpiaZ9LhpJQ/nUAqP9sQIQUwd4QAuvTS4mAVCn4FfgvU5xsVSeh45vLMyR
r109GpMlM0yEk+HDyIqQIWIQfTWC2DP6WfDTETiRW0F09sAYof8q8kLcurZR
zbla+nCKRnEfyUYpAHbiSHoXy4M8aBgg1c+jWjZUz5lrpEgzoe+QfPzD/ZhN
yIU35T+WkXCcMDuGV2U5bWqm6809krVfKE8+st3yIGEDuY1XqG757ipuPQtM
39KSXM53OPJVHSj0x5Bw9atxWRnVKyhZJcGiBmUXHsjYKCRVYOW5rBonIMdL
V/2pbqBF7jnI+dtiL/YScb024Ue5DEAVWw/JBZSJazrKsjN654CvIC02j+qW
1RISxpqutmX+hqhpUWGzDhJb/+QOue/UwakvQOV1Hcx1Z6labBfrlRyZYCcR
UpBGIb6OvStJk9UVak27dMmIBZ9sUMVcC5uhZHK+zsB2QD3fPdyaw0A8f5fp
p7Y64s/alrRCSA9LgEzWooNryy4hhYnw94jv4V0DSiroHyDM/VoaMvi+kWN9
/5gUkpI7xY6ANXignZIqBukp5MRrXbaT2XyNMiucmQEYAmz/qlfIsxt/2+UG
debiu2aspNcMdWkgLHT7yqMYbQVKF/Ixwf4XA+sxeie93D9/FR+HYtDgdtq2
umywRE5SB3qfknf1ThJaSSq+22in5ItCS5zPfEt/SIFMw9daSglpETzVQi4l
KWwMM2dL2jrvJALD5q/tcBZ+FQFpgN0QVMJbQtlaPfU0muULBrahVfbAuvU6
M4zaCJZgWjBuLlX5AuDps8gHPAjRkgfvIxXZxdUYKCl3S1MTtqNeBtiHk8LW
4PBQPtJgRitwEE8xx2kg4C/nb+nTrAeK2SVbP7QJdiSS3urPPvbL1UCBK8/p
E5eWDmh1YyYkkkhpGFr8ATOSYqJQjxnk9d7ZBX6xKLzWfKv6pnp4iETAb1zb
BGUqyDeYnwgG/Kcm02T/8yQkBA8clSu/UPUhWxvWLgs5rT29lDxwqFfTt95q
0+tq50z0vaE1kd8zBRqR3UGktXvQ+qjnEGGAW72Oqz2s5eS7r+ZmKnu0WQNc
fAhviDnFZ6KEJ4YELf9fAVemjpMt23vA6tGvb1LIl64HxKo6FnTY5ihfSa5P
mYHccsiKB9Xc3IuENGKBpKpTvg57pp1PcR9tNcmizYn0CxFt/XhapNGcvTW5
jM6O7xjyjSy7/5PNw+oyKEenDqjz7B+SSh/Ii+zqFN3zL2UnVcr3vGMyZ5J4
pGXb+KI0QvVlBIseC8BZ3AWLkStazafuiQXZsXiPt1mGeY0JSjPuEAHJrNAJ
AzgzSOnS2JEhpJ5NbvR5flRT1mXekIn59ySHDBbJJ6NJLRqc3d7L9dcIo+hO
RnJ7K8rUSCiJywfj346tcKa3vxHXPZ/ndOd/A+ReSU/uSFuQHB+IKpYAvz++
ru/gs4bqhSJt3e/HTEkiJWuY5TNicdoKZOE1H0oGH0cpexWiI0sMW7eVUWs3
gMQVvNTMyTQi3AwJkuoLwukXOaQTb6K+o9c3SSQMr+EXQObXI5DE6nh4qdU3
7gZYj2apjb+DaE6RPimAwaeIyYFv95ylw3Ds2MDmhU0BXoNoa7T9vGEhXwab
bmYzIIRGAjEDCXS822CtzyxSOGV9gmXBxWxbbIG6IYfTuv77LEhfXb4xeMv2
pO49AoITds6pUqK2Ev6mlnhN52Sj39CixsyJng5OfYgBmeO3OV/mxaE/EtwY
iE6iT3anm1AxMmBVrxtUWzZoiWlR1jO0JV/OEuyYF4nZueWMfB6udbI0mXVR
CWOSc6FR2qVwvAqEzORDzpFTfVraUOX0zTX23Y6M3K06Ffilx5y+mvltFtbl
v9LS2EXxm8emzYmSBtabbiWudB4gTCWO1w0nAMozN+GSqxb8ltk2CYE+GSCr
FHbrJE2Ac8Dr6GGJNt2ZViO2MYEA7XpCOtLsbMBv7EPKhWrwnooIRIL2tEL/
x7RLeAoOz+Um7wR0a+RCdRn74GcTcxL2BHiPMAXLWsOAHpIvzok66bir4/9B
JWcDkKY2vKYuOvmx+BPPgYfWW+gpU74KtnUgWZmW/yvxXIcmFiP9PpPIVahr
3VhYj5MkcTMCiXiSIL+2SHC9PjtUd2y05+ag6q7RNq7AGWIH56tqI8d91BQI
OI60yIuzE5UaLvbOvBf+ke02DBcS+ptT6iyvkrHFvBE8EQoG2+ipxbogMMvU
wf7grt2N+fKR21dzAGEps+xhSUUi9TWeFzJlFAQZKQvY+6RmGBE8v1RrDYek
zPt5j6BBba7qMfgzRLkRtGS8Jy+7NsTR3B96sGu5nqpn9rl0eg/9fFQHmGSf
pos/7sajwY5Bs52eBPTuxDetUdnX00JhKYng4BRxb6Y5tPoB9OteqKj/nrWo
jCYpZkkKrcgDvfi4tGwcfLe7PMpxrAUIC6j6h0oPLpqevGlpIKvbC9uNQkRC
Pz6aOJOBQkl7+OWl6ZHLVSyxKeVAIkyQtG7Jc62G0Cn6hRWwkKqCF2f6sGki
m7ZiJMCNoB2mY88awb+/DLGgxE85M1cjVweBnhL7ZVnBXX2Kb1V5Cnx2ZPiR
veQfueLzuElOP/5vS9t3jxv+VHBD7LYobkEjD4maESdRZX32fNLS6yJUxO3Z
1qbjZiOKfykFS2jVna+p1WQiWulcgQYmDp7QNV52yzbMlOm+BJOz3Ke7GyjI
YzW1saNz+u5bWX3H62FDyEpcfEGCBpstLbIOjz/MRcvRjx1YpAJIRwojP34b
9GgXUC0mlHKQpI47yeGxDS+ZlNNYA4L4tOAS2aDc1QdRTKkN2zYOVIfbmAR1
340dMSo52Cm8jhsZs/C+oQZn6LyNQTyq7lPOewaT8wVglR/Fln9HHu6zWEay
ptoU+UzYiLClq4e+w7iEWfJuYW7oOYJSYyrnzqUiafqz8Rcq01/OZ8h47ETt
DyqKOAy9nS2FYW61NZCY9kXo0VRW/l7qc3IRhsCXp625s4t3TvziUss+tLSb
KBbz0PoV0Rdw8qcOKSfEDEoKci/BYZVHToSzuTKH0CFlcImhW04TJ1L+HSuN
qDJN2PmjGUMWDXwJqUR2Sqpy/K37RuIhhonJ4lE8mJHB7HNAG23fVhhvHJ9D
2ubJDSUoSKu3+2n58kcyrOZrnyouo2az7OnpCOLcmWIElY9R5krrErcOCih7
TsN02J/kNUFghWXUAa+prdNAUyaZn90fEsT8ZFcQDasR6P+JpFUM5S3F4qik
4CVcS/4sHx6+zcoOukV/cFro0PleKItZb6e72Y30HcI+R+BcnG+lY/UBVWyw
ipEfJTTbYY4nP8yzzI7p4X3sSh3JK0mh0RfaERcjwSFzs31oZFAEbBymJmMF
ag/2a7fG09FGpWYaYJXAMCyojp1zqBGcCLPbYX0VslE/mzsCCSI13kHijKqy
zLIGEgudLm+sJIrax87ERNxYjizORHBO5rgMoLm3WK091CPKix+nzeIp9F2R
/i+j+mIzno6foPuzIe9fldCBNrxEEpkOCweRocVgScMbxv4YdpDPJuJYI044
dby5/WpqvVqjiPVRb8JYLPdW8NEhEZiIqEJazhQ1ikuK5P5s4KMwQdLaAGon
ykxDr+sQEtC26+NPxhwGWFZJ3JlLWXjG3DYK/FWgSLBisEi1fIrAbWeE4UeC
JG3ak35gTH2jmupwPEJnKeBdFGIhCDDMSh5nahsTGr7e2HF+7hsAZt/GQU/R
KXQSv4HQurJ6AM8WYpwmRXERvNnlEuNEEp5H+nFIGcxL2IawzY97VtiYeBRN
kv4tTB7mDQiylH1WBA4bAKjArVx84mqX0MUIAWNAL0uDdwXPaGQ77dDju1Nz
sosvQ/XRcxlFO5yb6eTxDBOOSkXCxCEOn+GnQlC4iFFV/0bL2niTFRI782pp
EXegf4eo323ure8hVX+X7/9zz8wWPM40lRj/HxjvselWBK/PKptCqDQzb9e8
kbpAkSRbfaBa9pbgURrLJNv5A0EOvI4O8mb1HOiGhgal9WEl96v1E3nxEGGt
u3hCOhtZj8cn4sYhab4H4YDYLVuRcJAAr3RF4nbpWlSNbTu3JmqRjLZwRSpm
CHyHjb4ZJV5d/rEDmwsFOGEFJ9Vk42c9HgqvFJ3GLA4ob4eCLgEMg0dS4GvF
vzQIXMK/6p35ENoAyVXnjvcUFfIb8DsybVLGyOQW21pTptFE1Z4HUZN0jKpu
VXmmvq2l5R1Dkl7gEDgYxRWydUBIXqMRFzbTjB7fvPTu8j52+TjK7XPX/pHI
jq/0+cQAJXUeTYQJ5pMfe66BAefMGqsFYABMTLBbbBSbG/+5aM1DJfvxmFRd
u59WFGKCC5h8dzYlsi/2aWGZS9tSoDoHBXFCGTx05v6VNlhrSdnZmF7w/8Oe
atxy3pqZr4eQlIyZcWaWwkWVa6tySktPW4SKeW3XL4WXk4RjG+ylYMCxfKON
7zeWY4xxCEbPZOS4FP1EEsED077ASCCYw/HI7tQhvJxmecvO09nxpU6Y9Ul/
W/McVx887y6/sfVxH9UpRKFuHo+POoUgEzqZ0vSBp+LxTBW9qMuHYEyDQVSA
NQcUFT3fJ+TQpzbq2Ooc/g0iaOCCS/Xc2d5oAmi6Wv41Erk2q/L3gUF7pOgm
DIcxC+tT2datxrFXzF+Meywi4jUZt4dNd2oFXC6M4gsXTBNY0ReI1Jip1yyT
84bwTLdqGfG7jEHozLF00Vijx+clzmlmDUE3FqsGHuw5qHb8E6oPQY3iuXvM
M8qmElCv/9nrWNJdqmtwkUgn6jJE5BwKYpeR89MYQK+wi5JWXneD+O2x3Y36
HUgCw5MSUs1VGIhK06gNtXb2uk/l1YYKh9LORUw6in7vzdEpPTO/0wMfZZ1F
CkCM7QGA/suQUASZ+99OfkKchbx8r5Gmksl9D3Wi0Teu00RpgCr8mwgPplIL
0OanTuJ8+vf7j0QD+J7tNBTpPHsaUstCD8RYplm5hA6BL7s39J5cUlsMGrPH
WLnfWrqhPM1hxI8MIpec/s98oSauMKayi4+QWRfUG9JjPLx+v52QrpuyaCvb
wteU59yGlZUdav7rFVYvBTDreop4otSqtCTaxjxbhc5OmOYMe+h1Bw7cS/vj
y+GIxfP49uKhCykYB0Rm+UhTDv3ug8GGd/Kpt7TjoXZDoYRYCtxvhvryrU1x
VmZDVVLsMZ88Mm8coQHg5MBmIBbMSDTYPg+juclyXBd3jYZAqeKrl/AWAs7S
VBbJ+HTXMv7jRwf/f+4WnhT5LhgMieq2R+PXFWtH+SmSSngOqXaJ3m41Wytu
DyKPpbxJZ7lLpUs2gPdyRLnFlr6HC+z81IGlN5wy1MUQ+o8sHBCBQ/g+qAdP
85AqcyHoVasdq/Gf7TLumY8A/u4jSawsJ73/D0dTRuEWnasqlRb2QXrfIT2l
cJp4woqCwGeJHmSPC2qvgN+Ihe4qmN1AwYweQIsh71b0X5scjrDhggfFCLEd
GIHedGd5PYEappTY3zu3KzbKDIg2cPOLc33eJCgCqVpWLGnKoi5HDIBEVCJi
1EE6ME547yq8GijtZmp0j9gMghFDmihv2+e0HESNhB7JpzKncMFfmzowbWoi
HXz15rWTyK0941SBAIGeboaLYgjZW03FTlF0Yf646uGZeIgKsynfhHgDmN//
pf+eoKFurraY1JMqx7DHezlaEa+GBKJH10N6PMJq7fqMtZHY9np1N+0Kc6lo
pVik7DAfz1kB7Fc6TUmj5578uFtf+f4DI6I3jsKhVEpqlOHbQVcZmWmhUcL2
54bQnPVWY80SV/mDj+f4xuTy+ErNp63hpU8M6sE4ULq6MUgO6Af8FLGD4JJf
JjvMW9reYtwaTCPkApqn2vQVMFeDMadcyEFLRfrlHgbx6LozN31cEW4se5aP
IyFc8K3FgAPWfLt6LweSQtQSUnaWqV/4MsW7/1siuvaDOcUO22UpXh2aRFpx
VVshqbShdgeIkTii642khLCuh4ceQZkIY3+Asn+7Rh5AT+FBGU0eiGCyQpH4
++KN3ZWvdOg9sq3AcJe5rJ4HwbLOLohwzHBoCeP6VGRiFgpeMTZp2FIbwHYi
W+ElBRHnuh5TafzpTw/HhABjtP/P8cUJhiCM/DtTTZ6JXzcFBhsKKr3XpF7+
uUd3Qo5hMIlLmLHPmtwMav1dww99B4qvZC6CXH4nfK6vH5nGJWFNellrs0em
NwPjcSAvH6QBvM5Do3i5lOoL2fiRJ1nzqqZLwUPvSrXUrn0RRkz1KgTY3tyb
Wlcd6wrhOm7mOKaEysKtCJKn4BqNOF2ju30YI71t4n1Yut8XGrYj8AXr/JLO
3cxKkSXiL53aFGvBD3Y7VStxUlX+Iaw3Vt2/G64chGb8REh0/HPZDo3ZIGQZ
VqNEGn8Yq8zkniZNwXzlfzNqTgxj/KNTupRydqjxHYHuA/NPs0R90LDEWsBW
W6e7plegEy3meBy+XI6Xk47GVtdnEn39y8aUxvmKZPyJi+IVZxovtHgryBJk
mTzyEIw9pHGqNYeRgXdcm5nShiWF7V4oklhiGHH8kvjQ2xd8yzQarExGNbKe
UeFgu7MXb4d0hp/GdWAAL5ICF09OF5vjhmjSdtpEtoChQhbr8tX7ZaUaezFf
obNcJASqPk8xGRhVpUgi/Ro4MF9GQuqHjfpwtT79nRzNhkMtXKAl+pdHzgk2
xNY/5qMwSf3rkZ3grQIwZtxsliqDXEHO09LrK+FIx9IzxdZ/w2duZWJ8qr6V
7wA1P2iBegJaLyS28mn31VTZ/nhRoB0Zj7e9XLHVVNFUrsn9Y/FkshzZowdE
9LpzVeKQEHMDeNhp9+uwsTmx7ZaExRUgsnZ60Ar9fhB0YGi1iz9RarpjSu5I
o3rPmpZ9hUqDrGwndRzDUeV3VlaFXaiCk1fuIpMaWQM6HusGmmnC3gcNtNU6
MlMf38nVNmlN4TAPPTCgHdRu85djXdXceN81JczXDneovm4iYFi7KQPRIPH0
c3Pzpsh5sq2ONcnMo25/2PY+TRw5vyOgwMnh0bpMo0rVQzWjuBHB61stSFjI
Q00gKWms0+/EK3N2t+FRWGdj2xgGVQTyXq31IV/o1ndEWM/3wIgmBGcVEUMj
W8jCwWn4645vPJBH1EkLy9g5oT7KR6f+uBRNuqoPvIOIz/HXDo8VwJZBTI62
bBaX2BDCG1DW25ysNTHf4hNlo0M9EBVxiLtRy5dDZSz076OdvgoKtSAz1jCB
VSOH9o4OCkRTjSmiJ/MoKlQ02yNLWjUE5waCRq+vumJ0OSis2myKfC8HRJ/g
ttEXi+ee/8TnGfsCZVgCsF9i77huxvfBZVIa21Ud7d3/qhUsfpUt8EIId2C8
zTWxC6J9sU8oTb4c2WssQE2IXwbXDlbxx9I+EI7Msm6SSAPfwnajKuVMgKde
fActE9g+ehjaFN01QmpkHGWK2K1puSHvI1o/+1Sula89xMF1ylvklSf4HE49
AFiIWc84VrU1hjT+EyK33HecFpLBIPIcyGXqU11Eu7wK7A5PADQplU5Om9tk
M49JAvtGT9k3NUEu+4t/ZSwKArgANCLfEURDYkdqk8ph8EiDhnpo1z8aYDBH
YaQU2tzryIG5cF5d3Hj4J1i0B4/89fBogiUFaQUxC0GpKwLUSl+ge5Jtqn7A
LEx6m+2lOYM18Tv3p11HFPFe+goJ6le2j/jyE23E1Tp8OG4yzluajV5ObbD+
SsRBfSOp7PZ0xbvfG6U02/4euhjetEr6KF/BXRnYMfmjj/ynSgeayZWmfhS2
h0kXau8P/MwQNBBfK5v3avZ9cRig9fgL0c9i1fi3ys++mfOZaYXxM859RRAy
W/DydXMFcfWOPyKK2lrC+AHdGuBfWorerBOfIHiF2Z3HpK7MR7eTueuefCcA
kqoOkDgm0MVywG0ZjyaXkFOc7qKNW87bBEy6lPNRXZjVOqkZK7iLX1QdZJFx
FeLN6t8QyOy0R2PkaX6daVQg3TaTspWDitsdEIcs9WpR8NIj60BVNjlnjuWK
Ek6DRJxb1T5LTvh1WGDUZTiSwZNDMLDnlLkRArDG9/KNKJvqCnhjf4gi3vKC
ALuBK25gu5QHYALY70AutQh0NTfEd5Tg5wWdXud+ZQQAIlILwujj/pHdBH06
3kwTTUHpA5PKGtOK1EpSAbN1uqNUDhVa28svdhmqBF9zvQOHg3eVFwPXM4TK
Ak0fpUbWGHFZHX59gozxjRepG/3ckSijSz1o1HfxtqvAAMU3ZAPzT+tHB9IS
jAzKoNBUcGMn39NnaUom8ltfirbv5fHQlExR9XS02nwn5U4vaO/MKO3Ca1yO
kPd/WmHhaCpInwgSZnVpYjnND2q41ghSEqKFaExkD/LX5qq4PHEi4Wc9tNf/
ZE1yvlmx+kdq9X1zhIuKbGyeqwOpn8uNlvoeXIr74/FmgvotjZysihoYqhDR
Gd41SXseRZWA3gonPD31Cym7z6qXARUOj4yYeZkadYPkkfSbmwOopIt7VaWd
FVSUXnRpyFcb8m0DarRLzKpSFlnH7sJxu8xcEzaRiPOJ7aRacm9x++LNEjlZ
2F5d6+50bvZZy6ksZXMVF2m7lN25MsXaFg5zWbkB+QOo1XAG432LYoJKroDx
/fY3n8nyUbaoznZq7YfjVL9oVhm534/A2vqZzCA/TRpyTUVnGEZLy1SxoSM0
fQD5O2J3tdiLWZyE8L36hwUleE2z8GhXyjUA3Ac0uzES23iQVHTDWuHOw5As
AP+ZRce4NYeQCFD8nGd84f2CQhgtH7XrIX5MXIalnggXrTZ/N/rl0RTyrQu5
4kKhkEe/rg5m86BOv3XoDXgJ2csu88lWUYum/Q27Fgx7/oaPfymbHbJNLbbE
D4SxEQzmEnSHqP3JcmPDrgcqmhPtCdWRoCtHlQMANqzS6O251XW3Scu5+kUK
Xxh3k6Y/9SqcDtZ1+4ViQFrPTYSr74d7aLeqyzTvLHGGmFqLJ4FSCXYUYhI4
t0kGjVvBxfz5dlkE35B4SXWLFP4Mfsj1OO362wFfPM5uauNtTFY6YhrLRf+A
tXBri864xfOKh0QEtagd2Qk3hrKir3jdLHcCCdXFyYbWZD6FwSysUdp0ZZkf
YqsXCvEBiquowWHKAu2oKbJRXrO3C/YTUlRohEkYvqZoHRv3fcFEr9ULQyro
NBik8/S97kAGFrv3icrgUiqIqSd574LpfD0tCcDHpOdGWEt6XydZViSGIdTI
2IKA+Tl9p9poiLhV1OGmkBULZ1mCh7RMgVMAJ2BinY0svBaxe/4fME1IZge2
MrYYQZCZcMkgTjtYI53F5tL+W1syJQPhzDcN+uLPIyXz+gDEI8k5Zp4gl/wu
C8Q1bRfzq8SfMWhQOeEJmlUhv3NOmFBuSwruzK++dqRB+qH84MaZhIOmFt/2
MHvfEYuG4+Ud8FCdfVbM8rWPP2enCsfCFyJRftz6wL9Gj60W/BckRR2SsE4g
ITWx/agDGWwVduUsoFmU0Cfm68JnZuJgTu4frxKNA0Qj46Ycah6yNitLjq1V
AZZyvdOeNkBUbk/vijvrr5Tqn38NEHrmS4lPZ5fVWXryhdBcv+v23nSpIYLp
rL0rqGTdM5J7HxCYFDuiGmyJyR1Ms8pqWhdCQuldQLjw6Tl1ZCbrlwLc0Ny1
qrzAvD5LOOD1tSnP9C+9+QHBlmem6Rp4KADlUFozG15AmS/2yOFKkKRFAxTU
zZ0UgvAC8X0rIlk86mwjlrnYWmp6cqFZen4I6TIwmimItRQC0Hnw5O2kW4ad
3cpHcYZVsLJ08RtviyWrVLOqPy5dB5+GWvzb3PYP3w5Um9O7O1/J+v9mbsO0
M8hL7AhSx5U6ZHqjQfD5YpEzrFnzqzTAaD5eYxdAJMKLmj8jTUUX5lb7H3qV
drCqod+1VOmX+vMHz9R0DxbvdzeOfiM3qYiUzvZu12gF+L7cB4YvyWCz1b0H
2jm9uw5F2X/4MrYVwAXZBN1W+/S7ckJNRzkxbc/CVyNsu3i9Uxd1mwOysSoJ
hSlmTDLoo9YN8L7Zf8YLtdFn9Wx7asKcFcaCnf0wwwsMCk/2JuMkzLuw1PfG
ZuuH1XTD4zlmqZFHJnhbcM8L8LeRj6Ivz9E6caoDcFdz04XgLfMyStzkzHNR
drwLKAX3Ecw6ehde93p9C9qDvICrMg5uQLneVYC4I4lF510pXAS/7zRXz6H4
qIuii5rxHntsS/v713Ug/a1Z+5rkTL40M6lGE6sF81S2ujsoAJFgf18P8xj0
tFXkT6EvUe1xDEPO07iJQOWht5qNHlGiwWJEozOUfesNWyUaoypY/xUBqyPo
A9SH/OU7kylnRgZqXxJSygP81dtgHOh5ayH3eJ1wPKm4Yg8LZRhghrMCCNTw
J1lxZJKXkPnK00KqcK8kq0nEpy/EQMzAelgEZAYYqwOCUa8e8EPxOqBBJOp6
8E7GI79twD4xwmm+DxNAXOTaSnNSAV3sa0JJ95znHrLvdibuoujqf117hCwf
1lk9USytSRpJmGm1wZ6NEVZOPVIMwZSgipiDnHR8GrOkMYPrq885WH5i3OPe
AT+4LW46cT1SF9x6GZFuvSXH1xEEAvDzTp4SWhfF9UHmyUPNfROfC574ILoy
XFvIxUYc9W8aLPLK0WA6ZkPo63m+3eveP3gRgP8brBhHR4l9pQqEXj17B4XW
YP/9qpBeQiZZJAWmVxlBwpiCa9IBBi1hBE6bf3BpDxfrvcGOVEHxDZ/uDjHi
8ISnCi6mIzyoGjqChczeowDGs3oNqGWwEmB2kuMoh5+Dwl7JF+qPkSD02QHc
tMChP176mzKjT0SvW+QG2P24RAucU4uDbOQMQ1VdiAJGZJTCmkiFdFwXHRHv
GwouC5VPNCp6TltvurtT+0skUdJszOaF4VVeL+KgfSvryhZCqsoDeBc5js90
QC1X0OPesPZ6wpyyuzdP3EboOxv3czmTERo3O/IYxmFhiSoIzEahX4Ck7odW
uAJiB3A7ixeWzQagK4DaxWdDML1b18o3sXgsVEI5nHFkj7TGCh9cecjyrMne
07H9MEJlxZZFTVjJlmhCNtUu+ah/m/lCBOKpVXLa0Sv9+T7bDusMOCYrTSWS
67lYh12uSjOYPXmS6v1BCRC5E0XNpFdG49rLS2ML5ebC13AJhG4d94q4yb0q
zSGwz+upgHmfig0LOvHsHlDGB5eiyTJfprEy+F3iEHYWmxfISAtlvEu6bkxo
0nqVpEH8sNLUHd2sfaU+AS6F4lStFCqrBRN9UGuMfXbCH2yWh5xq/kR9597u
iMHm93KKumnyR8SMIVq2DO3T6fXaYxCta6XnrGscvUiqgZZZLs2rixUCCxJu
SiDLHpCaoAzpvtRUSCPFjDogiJed8//exPVxbUspynNWpFODrV5znV4fSrvt
QiTlGzQr5ypknzcmdv+f14qVF8F9eGAs43k5/xCzyEd+FqPi2Pkhxgb4yILe
3YAWYKauKQAEe9qEUo9t/aX2udSy9v45l5UNl2E6Ip1xukSjLmoZ1VOQlltk
T+0HHieukr/Erm0udeDAG6S+30gq96wx50/W59agoEIz5CBnVvL4h7RNSqgJ
+TsIpbVgUVq8PEjAO+fFJ6a1gx5lkRaUYQOud1K0zeNcTwT1U0IxzPV0KKNS
laAxbxYRl3F9XEwN1RV3OrAPnlK62zol8DYaNrWAaIZUtbgtMpoxu7iE/oUT
UJtMzDEkjUHW7OcbdNKFBna124qNZDMm3Asz6g6Qu8BZg88mxIdpCBITpbio
FuHMhFmzUDAY4DYnPkKr4k+rgd+0E5QGf0qwtPgCof06uInCldLlvbSJxi6M
WqMJmKyeCtVWaswBc9BEPUUz8Db8OKMu/ffsmkqZxVNAGUC1U+QST364wXRZ
5AFy9of0fOZ2SqpFKtfpOGJ5dOoS9aGI6DyReV4J43G4jJDKt7/6vrqJmWc/
SPZ3y8v8tjEERfe5EUC7vOitwqOFqh6m0vuSIRvS9owW8cQT1fGlCaoeCNSp
4XixuQpo7DbwGrYr5gqbfVc+C4fgVXQRfUQDOXl5q+SAbULRVWjBrfxItMFc
8ukbNDxGZ4xcjsYTiGSHvZR29v36Pf35Xg/EvcCA6TbmfXfsu7zjvyTGzShI
nLynOxQeG6W/MqhqPPqh/zAs5vVIN0iX+Jh4BmHn6JD5OUC5MYfGsnDpkPAk
wzEEr8jnJHpFb9TZjFy+RfvhQDlVAWd5qirU26bdR8qLuf0HMcL2xay0n0ip
eUKVDqL2ilXjUOY2zDg0AasFqfvl2BQCW1gUdoSTMGPwW8bFsFMb5s4so+qr
9LOM/6NAMjNFrHWrXi/h3L5EUbohoGTiHQ/d0lTqVptjq85JXkYrtBghtSwy
PopWqMc4CXBSJcqYXIKZ1EqSk2nHDunHeElr+yLb6ryv6a0oI5e6VcDINYEU
QkK16A7z3oKzZ44mRCu07vCmk9AF1lkbUjHmklUAGlCfslxgLTKViFmN5z9Z
/hp5XPh+QcMqMzvfW6BfRXW+mfsfxTxd1YLg6tvjGCQ+pAr06n8U/bycNir5
AEK371U1tAqjtatjlG6rZPwDfgj1Q5qMLUIoXV9kydNbq03b2uPzT2Vv09qz
UrTqHtOsQ98d5iowsJCvgCJbrU+jrPFA1Rv5YpRPRTAU5Y0dXytyfpxOqhU0
Np/CkpfT7P4GmIiMWXOujrlqV1s0U/cXnJHywhDVD1UhXLZJ6GPP48gUOqYO
wh9BWUYQo8Mtf//lzyGuEKkaiX5ommPB93LdfuN49vid0nNp5yGPX6scKWqn
0XhgNCAr5zRRu2PtKtNUgBacYwC1qQ3Jsu4x0PmhxCzAme8rZnz0a4QP811a
2dyygGaK/j7dSbsVt+Vh7Be1ZdQLAOUq76gpQRlMMBtmw2vMsnkOxGoDmrCP
ZdJUPyaWt2sgEQrPt3+H/R2AY3P2FPmqOTyzbqJ/ABVElzZ10bs8494bikjI
4PvmyfN5wy6aqidD4dEoxb+nYf6g5byQHxebfmQZHd80bymsgcAkfl6KtFzS
ky42OE6X4eUbYoigoeURpeFjQpbHVgQl6RG3JwcXpYF49khdnnHvHKDBPBd0
JgHzxq+n/0pqpmJaPP+GEOOT5ShzaqSlMziOL6e2aJkm0KTNGBVw4Njx7dU2
h+W8o6R1d+mYfaIKhrO/SFSUgYoulzKYxfv7O7QS4ndMXtEePVHkh1k7uc90
VrK7JkNMRcbyO7SBV38mkqYnZsiVJt9IuE6g8xdvbolUb8HraAriRazjef0Q
6/wtbi5coGga0nPe1XPTxUXD6MBB3hHdlPjVcLnIr9DJJw4R+p2HHGrjL80e
TbJU65zntEm3oZSn/mmfzoROjSV1OhM2r5Vrq5KIzZsusY/0Stda+UFIsyl8
svnUPmF+2vAWaus4yosoO5pHjgzv3GW+g250nko9+AnpKdCJTWxTl6eilNUu
lpzux/Kt5kNaJfRuKkSVuwfv/QpBfLa+GDkBIySlbOqcZNSy85h6NXyZx/8i
2bRgV6EKZm1kox4NTO+xzqQPuM1tTgn+Ik9Ub2VSKMeePYfw5VPMS/HULaiI
lSJRtzOKPKzMOt1iE6LFFoitGoBkKU9/JvvYoXrOESv+Aevv5AYoIUTun0mt
EzYyRl/W1B4yFkz1ukEIGUm7MUywtarK2fVpkl0Mxjb4ZrxwyFTVi26bdMfq
JhTsw/faWN5a2otLZZvs7NR5KVFYbm5bSAXbMH9r0vVG1/L8AGvo//KvFKX+
K/mUB3dLQTUyvJsMdzHV4emnutnFNA+1zO+y9FVmnwybVNjEw+QM6uoqnDJS
76+drTXLAu4MEYkRNy07LOmIYmkRTQtktGjJx84oa4YbZL8vdnffuTi7YGmK
ESXBntIO/Kg+8AUfS6W1Hxf5ZmLryZ9iAqfFAgG2qtG9jG+tYJIxrTH5Q2PF
E/9lKNoFi7nqeUWGoHsms+p3SPdedMrl6zTmNknUu1WmTSr2DNyUHrCJ2siQ
V1Cxv39ghw53Dr64lCs1K5mq9NSGyo3MWc+NUNy+bcnAxgVQyR4WD1QTRHWv
/cA3CViJzLuC67Jh4qdgACcSxuyd7vdA1lNc0+VSS9fgi7TF5UP9pd1e/nC9
izgRARSCOCrnxhbrDy5zx92OMYJuSyNVw0z1dAD+99sG7tbcnIApyd5rR1j1
L9G3HWNSnhlzOww/33EDnl7/Lei2rBjXXHgLat2Lw5Ow0A9JYhnrbpeNDxCC
oDTyH4aX5DXPV+PLMHExBYlVtk4Cmf4WOysont5Myjth9jqmCklfS4qcEnKo
FockPaaQCCIJZqS8YdaExcaJz1f00AfiM8Ds68VckJ0Sdf20/n+swi2nAjOp
X95fB8zZAM0J+Rzym7YSxlq9WPy8qL7WEFWSOG7n49KngLYVeC/67pl0vvrs
sr+UnTbsI8QLO0BdeDv/7S6rTEwuHklUgGAZOS0pt2FhByfZZu+1dzmXTdu+
n2TjHEf6yviBIbNQNsrkReT57e0auF4EGoine5tC+MUoPU1ChSDzOVnuGG4P
grpBK8n/DWALnItbrKq3IIeWtsM6BtlLJO4uHPgZwQlElQ9rof3Fx/+4EHee
IOAWEukU7Y9w7mDpx7Myw2DFFwF2ITI/+7T0SaBe6sGMexbAKBi34DRFNrjv
f1D38ileB5jghoV0E4GvChx0guyF9Hc9A+L9cnMbw8seJj8GCwuSS/OBOScQ
RyAI1wx24DF42fH9M3E6j2FxLfTyNBQl7TmP70saDa39+qyDiGWcXKYx4HWv
SkLFn1Dcb43ieAsoPXYkY3YDY4K7VAr697UnGs0yFIrAvyf/wG0B41cCsMr/
Qm3QwZTihXnahj2N0rt6tl9KIvsZ+bLf9fJNEFnjHKicnH4UrGCRBXDiflgu
msltb5gLqFTGOhUOy2CMonEjS73XuhX5CQ5WxM/AFp139KppcQr3nEceCEPn
iVCuFmlAD6uy6sKw3MH2+7s4KADRw1Oez7lX+yxuvtUx6RwpdnGYtWUkUFt3
U1Qo9XZhoRGF+mfhBQ3g0iS12izlS6B7bhM8PhsNBkZ3QqcxQ3TE7YFQDQOe
GF9cFNzdWQrZPibCLUMSMChjc/lNO+HSvvi+WKZ9g36rD0IwW5hXDybuJ1dN
DJS2Lly+KvMEraAmO0vdILmQLXxSoK0xUzWLGMoqbdjD1JdowYKPug+x1TMW
v6mFsf48KvOBbD8gozC8wgTIteYAOhwItZ/mHLi1yDkM4u6pBg6xYAca+nKo
CIl7VheZ6Ne496Tlmcm52/Wn9upc8ZTpofpxqkUXB0yqXnNYVRlFeqT45isW
K/bfNuGqGplYGasAsxYach9dAkuwFvycYmFKbcKOKc/odt+8xYJzUP6PuqEM
i/tJ5wNbj21q7sC6rWvfDh2FoilTjArGESagjA5sxE39865auG0IRCqxcCl6
AnLyDvI/Y/tVel/fmhF3Uk/OJt9K9o+3rnP386XUCDSSL11Q9ChNNS/Mp/LC
jlAEv4zCBAxsrzisRGDL+8SNj21cOGo7pNMwx+VT5LmiRGafCXH+D0agR/DL
IkRPcjdMx+0lPG9B4D6Ffwj8FeueY/PmV4Qx6C9VBX26flCElD2SupY83LEi
wzHYM3boTd3MBflFc0D87rHg8eD3DSQprQCSc+cntdU4USIr28/SLHlvbpbA
jG3AX/bLJ3uJv9VnP74W2HT5V1LD5w+So0e1kyV8MhjscsatOZhTsXIJx+Ds
YqidTW9WtWaGOTBPg6uVuwXN9sNuAmgFje+kRyF1hbe5XerzVhDJZUTcfldD
7tWUvYivvVLeUW+Lldhr5EpbSew5CC0IGv9mmsbBcYoZKyfWykL0pRy9KNJO
pfP/6vwOeMsdi7KlC+2W4RrAQLVlNVVLYeoamsPNNQemh/fTM2E3c+/+yXbB
mpnDtQ013+n1qWVNDzzBUW5aTb2kHivBDmwnbalLGLEMUOZ8koIngKns6dQY
DabDR2+p08SmDyBEkTIWHqevk3YAdrBe7Nn9n0HM1P6uKHE/UBmtL5rv68A5
c9s2jqFjnFspwpg5i71hdIVuxsaei0ohVFKGXNjl5W1amg0EZe3XbMohxut3
MfN5NgO2ZcKis85086nGgSV/4DPf1WYVP/qtjyoQBfEwXmCwrFzE0YSGJw3Q
p3jdplri9F7cTwdKwYmNMKyJ3lKJNkgAcYbOLzPi2jOR4b2RW0Y8Qomy/ey/
jk7eBQCLLPWsxkCHoaTzZQVaySDImb6OFp7kF1WNS8r7JhGZdXic+frSUg7d
XBefeCLLkPzW9U7Oc8fDSu6Z0laLq3hKiwKdJrJwiSfhonWh10TZrgFTxeYx
jXVxCH+PUFLeaTb7rraoXcHufwZiIjAiXgXy6+B9kgebFx4lQhJUhTE4g5v0
6SmbOjFuxVtATNLmPUUzKbTpxqT6xVo0Zfg+L5c1LbKAsTHqrbFYHMWRutcR
U4VfKxPL4Wxt8QdeAMhQoiNKlDtL9FYcnrhc2ffN9FoA/HZeRiB2huaj+sxN
W2MEbdRDfFn9TKh4pANK57X4WswKLzzGGd3yvwfya0ghxCzU8RIeTSZwRmRa
tkJNJ5Pfb7Ok5NjrSPFPfKe/dNl8OSqu1hALeV9OCuvNXZY0urhcnWOUtdOP
KdiOdvy9vpTwWpqJHafNBF2/CwClvftgxsDLtNcrwQL9ZK3kcBZKFZKYQkdV
0d9bPeM6xRRLxkhYF+9oqPPGwA4L0Oy4dqiQsZFjAVQZG2uGP50y1wFTlr4U
1ASt8iK1CpwC0QH81ZAlwBxWNMYTpr1GyY0kx559XgzTRk/71Dbe9/BNoEI4
lhfLQNbKhzAdOyOqkXi+TYoPKYwPVwP7uTvdV1xCReZdLwrH2G4NALU/9Pr/
/cUGErwtV7gbmWgXhPZx4C4Zh4Fwcbl/NLdEC1ifMn9i2S054xFpaMSzofNF
dGRDnqkTe0ofqO3ryZekMgc1snYyujbnV1clRNmSEho3QjLkY5lNoeo+nmua
+HQm0XMOgABioj5HyfiWnHuJeLtxKC1pP8+cb3tD2eFGDKmjfzSBXsBqVit2
7dutVOHHhMEvvJIWYKWQ/0EPj0cNddBE7/AbrEXK2Wn93hsONdR7snsy2viW
KvMvq45aUr8Og8jWN/U8HyQC5zbqLCaebgIbQ/HSiTLuvmkqajd0h5ZnxTke
JR7LM8TScCrHHsWP2dH9g/+BysGvPl4Q+IlI1SDWKklDfHbpOUJcEZofibtA
Z6+J7V8z1HEmh4y/FfRfsOV1+fCeBO+Dl6H/1JuEKNVI4J46C3dabPv+xU2x
ZxPvdh6nzvyYIL/EdjEjwiK/iNyknAce+JtS/vCJ/mtz6G6gKtZXFRGgWctv
i9yl8IyjS3fcgb2asaSm/e5wfVp6/sEzlT3jCI2Tyv0aypksJhkpXLp9ETOt
JzQpY5jncYusl12G55u+gjz0oVIcAIieEIKkO8tNqozSgt9sGlpjGtE8hMdH
dLywNMEojnaFzmPxUk2Ei2/UB7s8JxCDd9S91hGV+5jIre3GEyWdLG5zuapL
E+3S+fBehbPGJxj3sZ/8Y13m7aS+ghoYFMsWL3NG4UkSabKT+TuFt8DITQHl
qxxULWTTij++cxhEn43+3HL22w4EDvxeILuYG8GmuATjk+BBAgpuPDG+gZEM
/wNXlWQBrtuiJo4TbqWzOZlZVwh57w0lA+4cmDSJ5LN2ZsoE+s6d6AdEnyNv
wD+WuDwkLx0KWq0tmN4aLydzmENGL8bVbFXhUt5qcKralERRJJzZR6kNw78A
7H8RgtK7wN53TaAgz8r7oGpEdJYi8HWinnaIaHMJADYqqoOek7v1y3jk3R4V
dJnOCeZ+h2tSkezN7bU56kWxipkXA28zXVbxMUYVLMsS+ek2IFEwRwbm1aej
pgjwYwAkU/+M+k+laVzEINdMbZuwZFzZGlCodswdOu5of81tAuN/gfyllM9X
bG9+B9YQLUiGrBmqLXr/dCgkKOKhWI10lJ37NatNVOYVEX1PbhK7+Kmw7mqY
dcWVLuOYXyXiqT3LCDMp77HTm0H4Q0h8KDVZBud9cp4pSuMGR2BWrBYg4DBu
3RKI4NzExzX9dtSM6LGHYO0r5FX+f3Z58rfLl4p/eileSVGex/SbKfBMUA/e
NRKg1Fia503uy89ZzgKQ6zUKFae78c0k3WGCgMrvDzVrQyLNJu6EnxkDC5Zy
a0rcdOoy1ZlfHeoucQ3bvIMx13qTTLo0yJIAU6+bff9SEyLvRlA7pTuCslAw
acskIjZvUfAKumDsNl1sV9NJOlO6S5sw0vDXyzeXE/hy6AqQyOOzAMPBYAUG
P2D+dC+fGpA0oPaMlX2RcmY62PeaVoHSg6XCAaFCAG8Aayptf3uqZ+RIcBrP
669yoCpM8XU0ecVYyj/WwNgpwmLmaxvHBiBVAn+7QoW77gfqge/4tbXZF6Uv
ZT24HEqb+KwC8PFFu5u+PNZWZXV6la8P0zvhDSWb+cQKOSWgaMw8oZM1dmRV
fCqsZwtTEV7YLVB3hzeHsvAgFPOQjJe5ECoLp+etbFy1Q2PS0eaLj/y2R+qi
PC/pdFlIdn2Zyv2LcaWqefg+/HpbXVkrIA9kxQwXcvaAbtI4HSMF2gXdaXUm
yDE7Cb5g/mH5lImbUlLNDBv+ld5lEpH5IENH7baMA/6KaSuD4M1U+aL/pb1w
/ppLDioK9scvfoSuliIYl3ANbr6hTowHljhljAM8zVBNyYPeJNDYydVairwL
T5b9xqsaHUVCIeYqEEkm5Eyu5nmGu4KOgplKoIDk8kajLgNDVZVOKW4TFcu8
UwtkxoIsxzwWtNDqjXBMj3KdfHVGBreKpUgkaExdJPGuMX1UUPtL19PxL+6H
bwFV3fFkT2J1xXhPYpNvXB4mpwdnudtkWkNm+KQom7c2PGle2oR7buygAJJ9
DkAl1Hhjzl5nkdzCxDk9bNLzTFXRiTZzRAdcZU6yqmeuhPDcGPYYThmEg1sF
5HU2riuswjtCYcfPeU4+2zKCgx+7Y9QeITm//w9cbtWp8KD0TJXsmsxGCcEv
EBggn4AdBwiGwRCCiKVLMD9ssWhfwbNNHAXW9dn/Xgaow7HGkNuj+JJ8og79
EVJ7Rhg/KjaSj9p9ZfzS2ou3qkH/QQrg860S8JmUqkwqmnc/LFZsCferW3Zk
BafZJWyEPm4yohV9PetpWh3iR/R1ZyIy+Un+xVvOjmCvGK+yujDtE1qEJ99G
i96E05GC0CO64Xf7Dv8xs02WsXxbVoNmrn77p4mkbslsykOzjqeYiEF/HmVv
Nhfy48Ge1lR8b/ofBo6Q08ttPEOB+uO4386T+tpCUNNqRlZ/OisqezQKTv1O
5yqpb5gVbOjmab2TUSt6YRHVbdnqg0V5oOyPdUiU0x73vhs1uKmleIgPcVUo
jK8bPNQbfH0YlknL/0af4DFmr1sa45dlfXkyihJ3u6Kfb+fn668LPzVfHm1W
Nsdjbl1v+f6O8UhIud0D1JEfBh1GuGLwoM/cj8F9SmT0BcDDR5vQ4xyqk4lj
5N9DQRo+ClLJKsUsZj/rYjHqggkFl4QXgTJXONKtJrJ5fctR81nRXHvpXodx
3Gao4hJjWB/8hDnm+4C/Nlkt4AG4WuK/jkX/4ubsOBRJ/zVPXRlG+dB3e4/p
eBFBYIRYqlLAl7+itIcKqFDxAyfe69MInSyz2d/qitU6gqawaSJ/HWnaNqqf
8MUsJmMOM2iuV5ks1PPM/T+ypJOOj6gHeABQYaKvdfWvkH04EE7lscks8+q0
lap3VNXPNFOZPtMA2MDxsIz9aOaaL8PzkBlLf9OG+JkQJ09mM4RQS8v/olBZ
1C0SuAwWE5w4E9s1n5S98nIrzvioAsSHdoiUC4oMkiUVA1CKH1Zii/F600Xy
EYXRWd/Cu7XesLjRkJ+EBf0l0xQNwrWH36102LkUvHwCQodEH5eiiBz+2nxg
zhLNG12x2QCvt8fuqS/uQ6CtKarIiQual9dVEwc/o29ynuC4ngODsPR7lO3T
JZWrIyW+RnQEM9g3hBI79UrLlJkDac9JT8ci2u4lQy9XJRITdro1CYWV5gd4
MvAPScHoHfKerWVhzTU9MZGbb7jlSAXa8CYa6JMMrOxoxT73sMwubQtLx6BP
NnKErf+kKp/7nX/DUa2URW3foqJ+6Ism3GPTrPT7osnRvYtQi4UfmWS6YPiP
A018qqJzchgCyCqCl01CvlZnUyb+KewMULtyTqKQDPACJTj17QmpDuy151ck
gzPQ1H07VGDfOS5OX5gNToCcJ0h6PfLKM48HdWHS15HoMw/1W3VeJo3fZ9+q
OTqszjFNARFilNU9aikhXfZYVlB6Jcr5HEDHcsCxyEYXf6NHo4S9Q270Fbj0
EA00gr1L4hKTztmPQ7ZXvj4v9HlobtQL1MPGsjhiDSAE2+jIGuWtPtFPVJMq
mEyT0wH6dVcYCGRKycgX8g8K8CJjTsURBj/gQCiWOePRCX8bs7/jFSQQ1Tvu
2af1Ohrf1ezIEY1/G3q0pngwxF5xG+j54wgyf+MdwWJqg97wvAV57XOnu4Jh
7irnzRJOA4ulXJglJylQj8FC7cvHmSCESQ49AehDlvTwbE4tCLm2Tok9x4ZN
nrS2k/Yv5eX8RvqYZUGn4sqG0PsEfSK0zEgIrBpJljQti6r9K8vtyxgB7Zq/
EPqAnVxoE0je8HVMfLhuGURe/yhQCZJyBU7hNljaTRbk6eAhizPXL6EZUjx9
2WWKr2a2XzNzdwK8CFnIfTouVijJOTufsySJiCRrLqxQ5vsKq0VHNx4UqGVq
cYJaM2pXSxv+l4b0EEoCN4ax7EsDLxGjy4Evg3Vefs4ap5SExA8TBCy1Suzm
XvaT0pG1IlRt8CA362IVlqYgzPlO/Q9kTllBqfaAZIdJqsgiv8k55O8W0gy7
bJjfrOlqBilNLOoritDNrjU1O40+5D4Xm+Vb2kpEsgzo7mgAJxsNFtGlnlmT
pldqvuU1gnA+qgZavsf8dGN+bGVMw1tbA5LRfYvqHqkTk+sr0lR8rNVa6/3C
UYpmrtkDlPc9DSPleoFVZSCVqsezdztXm6Qfmiudchouh4urUg49G4ZQJTdi
9kXS4U6cGlH1BojC78/VVCDG6MelnCQLEUx3mJfXwKdD2gookaoEhiXN4qc1
ObF68aqDIIBmnEUGCvdrvIR+B1tUEAfg8DrqiOwOc3AhH6+qRRGCiRoWAYsS
Sa0jI4w34vF404V/dyOq/6OrUTRuzcY8gtzxTZFpkP/ttkguJhQv49wVU2CL
LGTT2CQCvYhbH/emOIFLXZ637x1ZtKhRdCdC0btho1BiBnlSLXGt541B1G1r
tR/LY2srGMs3QrdNXVLzu+nDTCR5SLJ28czpRiXIyMJUZt/cUvTo51zTOCWn
0hjCcZiLHVx8JVZp2bBrbm8PZFh3eOfEu4XTm9xxrhzjGvmu80kIXuhXAB5N
onjAcD5/RH+8MCSXze/VJykQrcgnYtOSoyyV9y4vBQNXTGDS39KTV0O9iZ33
c1n30eMbGzNL2l+h7CikRD2H6XXN4vDR45gQvYmJPKB9HSjjizZNY5TCe5Li
Uh6IkPqV4iFvNBEz+Mm+iS2NJBCcIahlTvlYKtxMpuOrw4fR63ZHgyvTzNhb
OKrcRL0sJEITUqO8UJTug4CwBCoc8dtPwrAFyITgEPeDrQX1uf46sJHORw/7
0TSQ6dsBING/zhFelUSzMdrsYsAf9ap4lIrkw9cvUL+jY1HX1DWvZf1/MFNn
YRcB6MUIu451er0MhYHEQXXL8MWc4n2Udj/Iu/Cz0PN1i3Q9hubKzE184BgL
TuPJ+67vXQQDdby3T8ximhvh+ymGCCMQU37CbCoe9WvNPc/y9vvrdjuTR3Ws
hHfBnvvqrJ06aFShXAwDVlKuY/rAWRQp/09FZFJbDe3gcVckkvQ+mZ9nEQUQ
T1QYOg8BRNq001KmQQJD9ycTtidu0SXhvXTUfFORXhzGCev37h/AFrAZYxRd
yAJzZoXVSzTkGIXBQEsZhql8SFnEqkc62qdRGqSm4h0NyvKYRNz+EbbAEGIE
0MhumjiwxXJtCB8NNCS1v1s5l4PrFhbAg3G2InaeTzJZZQZcjRlJb/CBhOv1
/keik+nQvNfyVrcYQPr/6LcDHyFlfGoHKMiKyykhQ0l5dxCWSxkX2Tiufkom
08yzWaZvzFy4477OivOIBDvfjlBQgLvXqfMR9CHl2MAJX+4ql9VRxgNXBAYb
DRHgNqPR7PenJJn+gKF8wUXuSSH5GZUi2JgdoeommXbaSZc+UM7T0/PXn4DH
SKxP8lGIjxHT7/6PNXkxr5xkZq79dkCwjbnhc83GVLN5JdlVdCUr66R6lLbG
d2/fH4gJPFePKheV5T/JuLB7XmsVsLI59H/pTeGedY1PfHqlkTir6Q4WPT4I
LiEWUTU/wabuJP/MoMXABAKtwl1XdW3o5BoOrlvs5XhILVeZVEfpsj6yQaGS
ASjNo31CTf6PJnKj9c1MEm/n1sYI+SbfQEPsrunQLdqHNzSvHerx/ejsGJsD
u/eHB34SlAIi58qCF5/IfNxN3DfAlZ9De9kyMS5NxMHhcghdqtd336yTQU+d
y6mphrEkK0J3K3PD09ktkjFO1WrW9iIR7D3+4ONgS4c7XHGwZspcT8/ugLqK
Q9PxB2rvTBugVZ3x6K36bcmgtgPVY5pjSyuiHWSfb3pwSWExU9DyTjAdLBHK
PDRVbzBV4OnjmMlQVjgaX7QI1M8MDRemBN0CXaNxqu/Wgw3f3ypdkRMSQcxd
dyBAPks8n+Br9T2HEDJLHkLkr5M3VJg926wacDLXBp44ek3PLryL61fbdGxc
64JBjTxfFJqHs4nOuS9lZ6boe9I0ZFOYmO0fayUZMNcK5ehyELPtU6y8BPoF
i0nfby+0lEPoacueBNbDvvMLNRF/HEwX5WKpM/DI58DFJ57eaqn1w7fSti9m
FG/HG1vVGGpWEY4I4ZpX68qM2fZmhWnIJEZ58rJbxo6AkKD/hCWSheTHGbkb
Q1gPqrADUx54YSJanIphBFg/Ub1W8vw2QG/KwGhYdmiULzkHvWDw77GX9CYG
4wpUfhyM9yNQPR0JvmGn2/8RAK4YntkaeDEs57e/5XzjHqfJspjpdWlxN2wG
v3Pd3pNo7j39H7NWhd1qQl6LgfXgj/608kh9GvWaOYwT2HPy8Y39Nt/4buQN
N17LVEvhmDgfW4MY+h+c/AmRoFWsMT7LADHa9Nxv7yo9qTPe25FQeGtTYj2X
jRGiGmdx6Q62Ox/OijmNmVKt239T0VUxD8FQ5Rg+XhtfcIeoqeSBkw7mODou
XwiP81Drsx30532syvgm0pt2e1Z7xUFT/Di4ruMpaa44T5ezYEr2hGP5Nll2
tHzoOP2lMFTcaWkgPjSQ7WjZn1bfD1zLK7FvwbT+S/C07zXnOX3IPEqgGVGF
d9PiLXqGcXL/QKlKTrJ3hZgwn+bM7xQgXUlYFOTVWrDJC5ilAqFxoxaU3hJ5
zV5J5+YYpqNPWl8VunYSPwacLOzqIRkKUornSozSyoPjT4A8N0X8cgsq0O9x
uFe6+UNuV75rHXDYeIrr0hQb3zZ25Y18iYQI7bNW59VXlhViZgom8uZvV9Rj
z8U+UAAdOx/bVpSXkFAd7/ut9boPZ+JnrLvmXAyHvAYXkscTRINoPoKoeuPm
Phc3YqZs9NPL8vWoMTLxwK2MLduQvt9Sa1ZbbreyI0manhhtub23Icak4dxq
xBMGo5qWx4TNu3F0aCMiUwlQ/DlzNu6YW1q9weh8MzCgqcGP4NlDxUytWxzH
eYLRINfbXb3r/tnzNsGtA9Gaddg7KqiCyUnV9K5BXaZH4s5CTNQvkbzEaYf0
1fGmXPnz/F9meeLC9Hf76Y+3u30cob1px+pKNAW3T3BltlwItSddnYgPi/dH
HhBdOtEeQoL19ZSvSrN8FBXMdzPlqushj09XVMPOSJlu2NmDSQ4Me4btgGMz
NldpuKJGDBZUxs7BP1PakkRnhnfc5LmvHvli0JBt4QRbVbCPNdo4b09dJxD1
1emltu4KRAQJZIXqXkj4fBMRc/F9jL2DcOuLlt+qLWfiV/Du9Npr+u0Kd4SQ
Yj2q4Q0+m79Cq//sKTJtPLo//diBRFcJWZp0X3NhI0TjoNy2ErAQc0+jYlIe
EJDda90ChLCzXZ/pvLYKXXrj6sQbh9umjgTj2mQSoT/sjJNZ4+yOuFLOVfbw
vVEAvKPWZ4znfjhWNIsUeF0ZA16y4Tmf1oH2xQAUXYVpQWy87dBXJ1GrGSjL
EAfwtlx+xLennRgCTvE4XACwOr7P9SGn8S9FBBmYWFK9Qnonm57Qkl7gSO8/
J8p59VDheoH5bZGmpQjTop20BDvGbU/kK54crYhTomlhu79doHmcLT+i12dE
KRZBWCFfhqKh5ku9XsIgOWn7BZWnYWEnCKTeS6Jo0FPhtOlLuGAQ6G/tSIMI
JM7lUeM1hCi/bgMs/yTERrq/Ra0PAq5hy9WSMuQQOCFs0M0ZeI/B6S83XLi8
3U0QPp2xqI4tKPDtiSOH1NuuKvJ8z9ttf0nykUK+pev56Tbr6Ea6U+BWjeN6
x4HHRceCa2k0U/j5v0nhwfAhDFH1uGdtjjKHuneY5fv1O5Wy6EBlYeHvSLQz
2ARSbinSb3iLlfl4H1prXqoKDTF5/5N7CVF6z4FMZVWeOD76PkVHhY9FlCln
cuFz/yfXuOniE5zfXyP0tWWE2JI9EC/jZCmVfrvi9yZ9/ScpsQQO6gQAueXv
vwUM1To/p4k3yRR8IHqKFywODTrn2diuqF9OoDiFIdWosMo/sjj8tqCipTVI
cDGMXePvSV9SQD9BE7hQaKkjy1/jyFyCGzKjVaHF+APXlPr3xSK/VSNYDSQA
v9xM1H4I3DdSK1t/GVsao3BHl93fMDKKN9lf76eW2yId26LCWLmhLL4+4zzI
TA1hJOWfKwt2bRvkoCCE81e6aVtymKrsUW6ZpUhUWws+5Q8oCqCUbCxXjOaD
GQOd6cjCjWNE0a6oLh4W+ZdHl4AfU94IN9BRT2JYZSQZYF1gGZvZhGCINGoK
rzHiB7co2BSsICrtGXIwiK8Dtv38jl54dERD/M1og1J5AwMt1NWbAFve9q/U
rFaFMVio7IEFXFk/pylOy+7pXwwYf36cElfl11Hu+yPRAWivG8ejJkZADZlA
qxcyqA1uNKCP36RFc2Ol20vu0HC+V1RZBytCrAV4JIOLqaLeRyBVEyzVAa/j
TL9c2uX+xh+zdRe+Alze1KKisLoIilnivXwzYJDMc17m9BRPA5pfQyBnqRj+
9n8SmqeF+m8gg9hEsdQnLlDQkK+2DS7OZW1H1Cme5I2rF2oliL8XvMZIdXa2
n/FxQeR1kGcDZbrPIAPS4LOj43Xm9PvhLCNuCudQECeXmFvk29ycwbMqvjKC
PdmqNzLq/ptzzlXPjJyyFPGuUtsQ7WL6SgUQfPcOC90FEEug8uu6ylEjViJW
TTKBPVpybWIjOZd9YPmRF/1mGj3MDFueyfz8HREKA/o6PjgfWFF63TFbdcN3
3Dc6qp1lsZ2iAM8h6D4RTsqI1ky12DgzyUzYI52L/GZv0PYoJ8jz2kw9MA3g
y5n7PICJnzeEb4cwawZGquncW8+zXQPbKGKYG9iBOdtoL79XbOFgDAtUc9cR
hYkGyIC51Cz6eqBaQ28MXFmCkxvjRRNXnsDjzMDctBCR/IfQitAyQZr6GXz2
CuvxQQVhn3iMvk6EUzCSuxAtW0ed71JIQVZSgFOkJlbiN5NHKblkRnznPspZ
c4+eS+RnUiIZaqz3/VA05Hx65Gj+wObEiRn83ZtYhRSfN4PipfO9+oScs/jZ
GYiI15HHRb+5xWDe5opPAHoLsNGIX6/WiWEjy3+cD+IxNfWdNbcYX2+xhCmJ
uNujpqzfzNydDOJrXh4N4vQZL6YPgWMdi27b2dVBjnshnoKlBTk6EqniZcKh
/Xn57Efzq1tzsKWToD9t0bCQ6ppjmfYcy84nKmv+yajhm4EQsMBTz7LldL1P
6b7xpG12KEIwCkU0cgqLPR74KmPXkJ54qVW6V60Alg8ttI1CDZbjV/ugFeT5
/zmQ7jIPS1sRaV4tfvab1qGhCnlosTZkJY197G5zO1WEjHDY4gjQA/0t/HmA
9n+AY7emgPXhkacvzNpKmsogrTMyzadHL00pg2VcYASZVO/bmyaw3kz5cMCJ
A6Ef19mPSeXNPDCC4K0wHkUqN7mMzjQwujlSOMMGH4+q9rVTgHGkWLGe1Q4p
+urU0AHIQs3K71v6NM5Ht8d58K8PydndAVcNWKamfiDAfdQVeQwxTXT53AyC
jgjP73t7wcpmAdABOov9VmJ8ZbxQ6WIO16o4IFCzVhrzhPeEUCFv1hRfJ5Wz
zF2oVFYC79KhO85/dP1mXVFKYadgHh70TX2BBqJtebSgevOjrftuV8bgHD6b
siBpzhx5jETWXNe8Cdc2g+NaJQ2RTK+cKdxHlEaxYYaowYdcWcOzWoxo5BvM
WaTJNtONnVAs2XZz4gDnq7DEOJAk9qUpqGBC3KCYqyJSs6jtwWPAth+zOUfZ
hquEuJF170MshL+Xvv8QmdAWysF52QMTBWZxC2gzTK8TpfInzQhCByhdT6V8
VUoRT+5rqI9TCiWRm1H3WV17Bag1aczwDlPkexmhOEkqowKND5DlsMRz3eok
eVCM1WzbJYL9Ic23h8oVZGwrA8EAdiD6ym1oa3mEDbl3ip70MW+kZYmA6N5g
m6wBlIGailzF+96RDImFXUILPAgGTQ5yF6zEtGH/L7m2MeRUOsg1GskEQYrJ
HbSHwsB7ol8v86LXq8bswrAbp2BtzCvYCpS8tOg36npwIh0kQsYI7mEpCyDi
5w9ORUdzlsEKHI576iyEUgETex5SlrXdFjkhBlPPKI7LWvp+pAttxgzlRFSi
/0mXVINHwUg4Cpvooe7/HF4oz7WxeCKq4amv8b6hcQOVqzmv60zOeQLzFRIA
trz0wLBzjQMlNiOz8MT3BYAj86qDvHueRQSfzD/x6YXgDr5/eVui5PfD6W7Y
8aBa41VCzQO8LC30bxEtRstBTBnvyGezfkx6+//rb9yihpadFd18L1pn0UI/
9UoVMTOs7bIgFcD31F4RvZkV/cXgbqKfHXdB4QbqoepP2fBoD5Orz+hfVQnX
1Qur19UzkJITjF15LFsjdxGP8lnrlTmiu46KlFYOtD6FZQbEE5VLG3uewx5f
O+a2cBIvz8QOKD9f9E7ZlpMHzwWvlz4YLF+opWyiDCyeXL4KI1+3RJ9J6fdP
tvTn+hqNX6fUhAfTEg9s2sS9QQIK9oA9R7TJVDGRIS3APk1gg9fEbWNz9J3o
0qcCF00+6l0QBkKTDzMsWS8XCRdoCGOTaFvpIASXJzQllFWEw+8hggDAVvPY
Ps4xqDUCX0a8svTcTGIMfPBtFCJMkusRflnEYHs2DzO3p+f8lMHUXURcNdxk
xO1w2ldSjc0gXdM2JOscsVS7nyuPSWc4aeLvBYFfMoJPp4kv/zW39BGoPxVW
110P6C5B6jox8rpYvsRYUNvr/dsSDgXGCfNMkwRMKuY9D3uKns8+lIZbYDsD
JPDru2gA4OnJiKSKyQ1IiI09FZ+E0WhyFqjh3WVQbj/+TsyxMz5MLx3gIsuM
4zsxS2dUhoocDsCwQf/G4Pms+HvEUJbG+rpFJmue5lYhwSBMiXGNEQ1s+olo
abRCDLmgFsN/rMZTGSyp3qUhuSVxkoub9LopuOuot0O53Q2S2Amft97abLUG
HxXQcM8VTqY3b7N3ldB48bZAgR8K8UVKI3zOFQGba0eIfE3s6N+EXjmGzmff
RxrwBUU12Bp77xAW1oYtoAns9GFmmuQI70tAyTnVyvjGR/yRBQvHhZws22TU
hkBYrnWq4sXcWebALuoXzfBQ/Wqgu0Pmfc8WkJ2EzI8z9RHnBtvXmHDVbb4e
Zil5ds+VSv7RlFiGmiujbKchkTnxDHrsWqvAZeHTB7uKUPflAD45zWL0xCbk
gm5kMAOcLG/x04KPUnajkZGM+6wr2p1GNN9pNRaZZzt0NHwrFLx1P0hHEGR7
niF/Q5KeQw7hRD1ccSjbkdalwIgON305Xvga3FHLhk52ntl2vpRYVjGq0H+2
i19bSsWntpFK+SZO3qUokubB5pt+lqfGtHdYVtAAGGqGtfoiFaSAUiPjM+LH
npbqWSj5OY0exieTNWU3Uxyj+asl5sLo726Rm1Khaw94gYAhV1DN3QtLK8SK
glawKS60mJVIO7/WvhEr8LE2STzi78qwOp8DwziatuH0wtGuXW3zDdb1o1BC
Jy25N7SdKApIvVENkYVQhsGI0H2aIvqODKcicg3r8vyND6mpA0uR1tNf9kNb
BnuqVcSgxiFjhHo0ugSiwjiX35HC/KO7pRegkP2t5VZVo3RjG93h7tZud1JC
i2O2ug48gjwE9oXu3WjjrDCVygUAYViXJHFe2eJIWUaopNUfXPyQ2jlBNJTa
OovkGtJNSQ8NH0uPCxCcuaRxP2Wq+8d833hnEMwJhCMSTyFaCsve583GfV8C
k7R6JDttc2EKBaDhIhdnmHlPywUbIR18HDiKD2aI7DyhGzQL1TWeDJx4LXD3
BFhjWKbAmeQr4CBski0Ql63Y1/sZcga/JCPjQ98RwMa7WVefQ7QCIo7V2ZH2
uSXkLWw6o6waTQFKRcHkXT7c5AYE1n1pRab19zkfX8E7i9NuMXnnNJLJni7V
ab23PtT7aga7/QoihCdSm4tOXMN731ceARq/4nqe99yZTGbZdBuqvEkibkXp
vBzDiiqYh+7INWlG29VkelgonDDhCfo6mvRz005RZ2N9rgkj8Nx0EoBu1y7A
CHPalnM5rlKMm55PvbNnK2XpIWbf9Xu/vYREct6k+Vut7cdza2UgKBfj/KSj
aPKPf8w0njt4nPgJGBkrArQ4qtuZPz152dRkj+hQsHVjRQDaTn3HkNPro2p2
GNIHM8IT+BS1vksviqJ1VRmu8Vu6Auar1W8mU/Q/5XLxJGlo8MSdFf5VLLuX
JyXzCiMnmyBMWnleh6fmevGXlIxsa6b+q4hNcAuarvOIIuDSvL0QGbXaErdP
ddoAmpkN1cucEvMSkLQDU8aQP+RuW0MmDrkN+KX782NJYuDl9Lxjv46G/nF8
sFYJ/wySIHtDIcyOPW4OS4Ic266vPv1+3IV3ZL+JQoO2hjBSg4/FwQTBbBbe
EKuXCgtCn0r0vEFc3iTz4oTz7skD1ECYN2kvs0nJ9BOCBuhefvVvgv0FQp40
KCf87ESTUVsn02iks17J2ShIJueoaliFomHuZz28V0C5HSbcvRl0NgU0lFFe
58L/BiO3My+kk0Te2IFyEGG+pDoyBVEHHuOTh5n2ZMRZSJ51g3k3UMl7at0L
I0sDkL3GyS0+brbXQCxOlwqNqeZwObHRYE4TwkqFVsXx5zNad15QXm1Ohnt2
qpCp08SRw9XqyYRImBYQgwp/PE83l+mu2n9X2aCcLMgp0PFlInRo6U549ZhX
d4/bIwg9vFxejNG3DDKXgCZxCC7yTOFo1eBYcgzegTKHUYH1ZFy/iorjE41N
SWk72z8mLeo7ONxzgLqmbYfkj1RDq3K9cO8Ow4TdCtLegOKT40pVjQyjQYHQ
NNhOCNkBSsgfdxTiqfuM2TshNJnLj3qzLfLqgmKeAjk2/BoY8I1Z/ch93L2K
1AOxhaKKjEr3ldQ11+JVJ3XBf9H7DSYlolJqdEflJnirpMihGy/LaXXW7uqZ
K47Yd3DymQEiZI6GbclemxKW6L81MsN6hfV0cncU2dVeeNmgzS65eGF7IfPa
PYWzg3Mp4if71COihU7WKtP95DkFHaKoadc+k5KL6g2EJUt66VkJ22janQDT
Sp0M2njHqFgkBYwM9bzKvTFheUup6JGHjh0QNFgy7RExwrYd2m7rt3BTJAlh
MH31k/K0u6DPgBb1p1V/ILZX0EmpQ5/+BdxhUacsRHZGzeiCn3cVaCFDA6jR
aDFYnJIMcyMukSxvLn51TmRpfCxycANurnRhT6VhHNGaO75xYagvQHns/1l8
moh8zcPkO22tAxDjwT/C3/6NfLmScy6XPQLkvlWGr+bMLzqbGNpwZrgNaJv4
tN46eCKkhTN/lFx4G9MNKMx6Xn1ltbLhEyhueZPqbDNjWThuC1faJzx/BOG0
S3TRgHThL8cl7fPsn8puoCFGKVYN2j7tswMa4dluiQ6n7KaqaSc8+bX4dOEu
eoEe7jHsANWkvlMOVAMnQtcjjtb4J0EJXzwWR3HByN+GLwaMxK40eXohpZx6
3PJix0/40+LwV4zKL6eUzJyLsUPmUacpZNtGMeADOPEBE66NMP+szcKAvMZG
BwNi8xyZiMrmrNEW7BD7TPIUuyGppxSk7jXb/exEAe/+1apctytlgVXf2mTq
yBEA9Fr7v904a5VDj4iQUfZ7QRA9tQBI2vuY7Z5v2sCYfdcMUZz7ZT1wBo7t
uRplxtMWAUIicU/XfYDETIG/uaAfaw0o0ZRWV/ukvDRR6qmgICSOzyXxAQw2
PGkXInF8sIKKwelZpHYW0mx7uU0eFoO2genCCZ3xPNB2nquw1tXkcNLa852g
DDwmFp3MnpSN6YN+LqvcIcHkApO59tUfS4LTYzmuMBUZA6iz9MejX56/hzLL
1LHtd18xqtQ+7qMmZumJnc/bSAdh6RtLqXZxzd/sx32opqzSlfSkyW30RYKw
Ke1Waqzkjnk+FqOVR3BChdudFPy3TPolkRmJRrXlLUKrzQgFg7Mnl72aNZO8
lHyOkSfi2R46viHDcIyfumWzmnYnWVtxyyb0hTMNAjPYwXqPnkbc5+HxlGYo
+M5u2b9SX8/mlwGQPjy4iTbGwUmKCJ73+tcVa2ws5H+asLnzWXVVK0ReweEq
DCAWCUKbqXoFZoJfsUKupRUsY1HWAehR9AkIaFlX5RCqRa2rziPVwq6NrSA3
7wD8zfxpM8MR/ERm41D213fkdzZvyK90zKCSgrfsZDFjnS6U3wB4kMHVHcwN
kpkhqr3IwWVsSsOrylutgkmakIOMAMuqE5NzLVyE5QyLg9A19y9WwiiRYNrT
N2TC1HJMP4mcEg7SdVf+KCJI4TM/fX4AorhSUAbfqzj3FYtzy8Mpv862Sl3c
vojP21BcYmSjfWVYpkDkbk7z1bBzrxcB6OS+0F24G+g1KxpwFNu/dqpXbm8Y
fGwIRo+RDHsfgkb7C+WoxGpJ2Xm+mJmuqcdFy+i32VYS6jK18Wm5CGD4u/II
sINpmQ5ZM0zUgUAMPxF9kilsk675QwmH4U6QSn+MaoffHe4otaY2+ztABueK
dioqonXFgZP8MSzVRcBLuHfh+7M0v6qTHiYjxx/dwUxLVLZmV37S/yXj9xcf
8vhCbLEZUSsGIGC/kubPyKMXtSFddsGGkDK2Kq4szbwQFJE4cAWpJ8yHpLfJ
nirB5TqEVOM4fepZuslujKkphJTcYAFCmR0+M93ZnYuwVVI4fsue/B85Tbid
6l05GECcO7s5N8rbRTihvhJp066tn2m0Z0tIW3u9uv2AfNAnJsnfGz2K/fpX
EQXQ/Lf5Y+aZ5J3wyglsOJ71m7yATPtCWZ1+4uT4+70WY16RZp7ER7hvC779
scQWuhn7f/ztOsJJ9q6t4mmlMiSsg1byefwGZ76HaEIQvG9QWtGIhaNqALL4
c3o1qBIAg9WzGSjP4zrQxRSHWIHix4ZZRYK2K2THiVJVFwhpmTCAi3yO2fB/
LQ0NFnV8lHH37iVQEDJUiJLG4WQNRRvp2TuMAzxy1SnnVR0UMyjPg21HJJeY
A2paYHuAmgeU1yiJXwxbmvNJmcSZqPxZJHF34fku5MKVR4OcLsbVyYUIIRPP
t45Z6lANGFQMqqTBncon04Xl8MgLWwToS+4cO855KKkiNyr5HhbNcyHTjzEB
9r32djUr0nkJ0Z4ytpMyxa6zr6IkUMoo+VdRGJiOvXk724CGiTDgt6Dzjuqg
WJ6gTkO7CRNsDuDJfm5QLKGLpnHhW/lXhH08lO0op4H/iJo9+K9QQXIBPPQp
UrDNzCCCQFb0SQAjZPzL9WfdxMUGclK3SBjs2twJcZvN25zv3dYS01bjhFPk
XA2xRBv+J5FVDUNkaR90y2+oAZmpCFRlFWQPWlI9hIcGzlP35f76YTSn2ZmG
t+LYTstv6u82dHPETNLbtlu5evuuvCSQaZOYNJTp619W2d3EogvXbbM08lm7
ZBfEdX/+bgQUh+3kg/ULykqX0sgbWpWsGvu52mkrVduRYIfXaw93gLBSKf8K
rZl+sz6xiKvj5ghjw+yFJexx0qo0ItKlWp76RoBUPSf9+feoGeQYqfbJK2+c
7jzlfMyIiJSVc7xqLlv1YVrJBEZ5/7u7VVBDDxgNI7GVSyRYL8macabMti1g
3OMIg9tnyHfaQwbJvz59nEo5SanSKj5VpoP5H+09YhFtmbhEcACMwf9EWvMC
cfvSHOAn0BibAkpZURqhpRc8hl2dxnGphfGKHvfuod/MQFY+blxkaSMYa6YG
MV3hTdxGbF4Qim6cl7DZvtuM5mwdE8CAij8mARBlDnesFGQwVpc8iFFBBWfK
co0xkEcX0CqVELcJB+AgQRr2yn3m/HTe5sFKv6Ro/XwsDfKEIEJAPmHZqUIf
9OjyYZWX1WlBAFXrBW1z9qMhHNYAV/iJnTOlIAt268EAlnhXZNoUJiDjy7fM
4Qp28gTatEcfo/mtODiJcoSCyauDrtN2m0bPRYZr4iXLADGg5ICLNHCF0hnM
3jXOc9OHrLEqxaOLRJbVP8z+qguA0ZCV1pEB8CQO8mySJH8IAe5BCwa+tpUG
fR/xpIV7iSPHs5MJbQoKdHDh9ntPAwjza7bPLyE4GXZTzDUuXC8Iwmvd8LCS
eAmekgGsf7Mi7A+p4GEpW93uNSg0nm9R8tl81S+EsEx/Pa+4IWDlKsWDyRSF
bkFpz5xhLpt64AoE9psRSmZQ5kyrFP7G/7bgvaD2uuhAQ2e+X/7Ee+7vXItS
WuNKwFpvBpdmbTxr7zBqYk5V9PAOSw6NNrF/FgntssAgqTlR9o2/glsHx1G7
5T5OYnbXUsZRhK4+L1YHjDdRbJZ02KjbrQwIvlJQneD+EuBJZhNmE2wWvXww
v5XbTaqjN3HZeTaQ2eTlahuoTA8algwB8fURbT1g0L/n6ofycbHcqTkUKSv8
EyKl148onnglYDvAuJ0q/+NLLDdx1KqXZ3nTQiuwtw16YT+G5TxbX2RYt2JK
ukUB509Is3q7C/mVq3ebsbyR2k9Zh/FEBhTTQO9mYQFgzrg1aAJ1h/robg6p
b+D6YtPfVwTjdXSNRap7S3qiGjBOdcY1wWibcACINjv9SSqQq2bgT6HA+jni
NVO+lYuditjy4/WSDh5UKYqtXCYoTzem8bhJ6yCJzvkKx3FbLsPNqtMAjOj6
FgDrgUAgpredTaknZQIdnPYJhNpXqp1N38AXXMK8RLYDxRfj8YN7qiw9Wu5M
0AJXbkQYRpCKdIs1Bs3e6U2mGMaehFHdWL21LM1E7JmwFk+smbJbYYaWiknC
aGde1lO5Jf27UrQFShm6052wnA8wYPtFDCMOQ1eVpMdKLkiUgsr4n68x7Dtu
F8Dn9d8CEqxjuCN7lqTobQJpqr7IasicECgMQZfnh1x5uDXVck5kOv9ZPYCb
SSiIoCt/ZwGY92I4vm0fhKe9wRytq30s/gRIPZb8zwpy7wWOJPLYZ2CLTlP7
GgJFe9/+dL0uH7CkeyBwUqwyyyilffuFfalnPJwq/BfiTBGH0qRj+QOw9M+s
P+jh1VFU/wavTaS53C7OPulNDHb3aKaeeH7T8LhDtSxNAsHbqxUUuJd4nrT7
mRTtnjSdiK+IApw6voGK2dFAwH/sSMPUlL2GQmAE/7Hw0QQVAZeIYR/OcRXn
RkV412ZDxDMTVpzZvK9XzumHNkZ3zd8cnxlFwgNcaLqqUCYVvPtByJjMfbPR
OkCgNHcMeuKpgQhPwq4/ap/BTm3JbBC+KCeKyUsyNwaHbGOfsURBOWTfUA45
Uv7LTpvOVQvpwq9r3W6h4S0ibkQvmULbvb/UZTJ5WwB8zHGv7egk2W9O+YfV
3RULEl/nzxNYRMuwgQrIWZLS/0cOkFi6EICUNZRjKocjVW8UKW2f14OuR//v
THzMc9dFUr8DuBQ9Rv22Odz1OvOyG90wmewxAraGHn6f6O/ZUKHSix5mMcRB
taJCjhMCP/xAPAau5jxIzzryQ3NU63e6X/sPNWTpzd5KFARMjRwmMIXv02NB
C9Y7+IziaJ0s3QlXmnFG8XHWmokWimCjW2jgHdo/y8q6yrxnsu8exwQDx6Qd
MgWxBuampwwmYxm+IbC5MgiO/i+Nhgln2WZ1SDCzKe8j2dgbOAhK/Np9Aa0A
QocITBKPsb8J8LF2zz7YL3A3RFmML9sYS/bLVAHOlDBBsUzT6SsccFi84sUs
VZRvkazFHicDJ52pSRaedGT1dNoH5mNAWtCJvgxw9RhBIr5C2Zz9FuHDvsZY
AfYrTewxbY0pW8slATtI6KkDrCJ65bYLj15eT7QSV75qij+t7HQms46ExDwV
+3FSbd3m0pkGG3GAgTGyCfT9CtRsVaMxVTjtqPo73e+p78kaEfpB8cwnb2n3
mTLP6KZkuJOcmRw/Yd8s930C9tEDYwzkrKXOqcFMVbE0Hijm8kECB+ocE/wV
a5bKsRFM0v4N6vLl4lO3p6ElyCJi8Xy7dWQuAB52Qlx4+fNybul1/R3pRiZJ
xaZTuq/PkEddmDKfQ4WbLc6BajMTkWITjyk5dUva8MvHaXNO6KArqax0j5Gm
5I3l+e+B5VZBkWmm2F5TwpWyH+Vw+Bq4w+2zCyQpECYJwvDfHE5US4vOUp2J
RpmwGal4PbHeJinFq0Q0ewYvGKqfkuWizP72hpCgXTYwW/W4Uv0kn5+UT7wH
NoYBOWcfsZdJBWrpvqogCspC62pdxJ7QKyHjVpz34UnKb8oo4E6GvI5mvsy3
jBZ62oZs99zXIP6MgQMKVJH0bspAsbIeVMEcgXi6dvhuf4LkVMHxBatVVU+K
s+TLf74raMQJkbzfVJqsKEOH5MvOuNeKUoncUK6mKVMtmJtBF3wxXJ0Cea+9
WD4uZQotiFOK2sq0nvPuAOvklg+SysTOPVXvS9kggHhska7YiZvtMl5Bpu/w
xjeaUQHyyDDIzZNPV3G3scob4b7T9eWlzxHM6OEMB7/ZalQv6l0l5JMf3Nql
BDas6Qcq0HaCDEmPtA4OzzolLrSyqnf8pIqqV8q/ZdT16QFKn3HeP4EFRZPP
vX2ggEiG0RcdphD/kafTq5mECtVPSGqjLN74mLYuW31+BEOxwa03Wrx1bfWp
f/3DqTvemzNO7QoPgqNXxVcR8lTHh2yeOy/IhZIjfLE3k4E9j6O78rDpVB6f
nDXKsV9HYR/gyfvjToh5ZmsHOBaBu7pYmaSgJn2vbpt/gLO2/WuKqxR1GKQH
9dYDoRLa9EAvfXP6JAFyrM9e4FyKta9WWiMurJV5EjTAS4BL3ScgRCQr8G8c
oA2VPSzVnhaxLH02uKw2IVSMBIb3iJbTPICGk6SxDsZOJ6xvW1rP/dhPQX7I
SjQWApLRyDo94XLuCoICk6Ex/ciNj8CmSyasFZHFFN0O6aRAxvYm3a8pGO6B
3nOWXz4WJwm01cRyGauILV2psVqTvg7UQpflLd7BFaRRyLLnEs50lMyX+Lrc
v/Sb5cx/SxPrk9DfZrKsPMdO8PRPRLKlKZxxVP1zBO5ipBs0kVQhakbOv9uj
86frhH7HdAKbYYlV0GTJCIJ9QcaZXSYJ1trFLL4eyX7V9nnq1vp03RHg2oft
iimnXhu99EctQRqzGO6vHQ2wjHjX1WpDosglqfwB04ufgLSOGlqVm2pnYjFE
rdA1mDgwslvsMoaor9DmvNRyNyQzkZamWXC/1d+62utErGQ6GVHiCctVO/tn
UO6v0wTOa2eDegAhaBFVp79SzF7A0DEiZMTOJZBesrubj9UGSpgE75eEz9E3
00urXEhaar46IPoTPD+fiMEvqmNkG/eS0JMd//ZjJwKBj3x7B6lOSnu6O2G1
v3BPSlyudLV8RoEUZlGLGRNuUsPDEgl0Y9q94y8nZdfdMy0Yz0+YTbwJwu3m
0jVygI8/2etTNgsektslPpPi5whG4ZP5LGqyp1w5dD8pv5fTAU/DwL5zkCim
UmblRqD/YfnbY5oZsP2bSJGZzfAtkzRRtAroB8kDdkUvhJLOH7l1EX4zqKX9
kuA+RRlc528/umc2p2NUTPqiocJnn40d8FhJA9H48ffbFolckw+w9qCZgO/p
tpTWKerLLbhJvC0gAnUPfKLoZrjTp+XBYQbtnLTLbHyFNrCD3ViUX6A8XHu9
ora2LlsD1LFhoQejs8idtW92VklqGLuB7E6hHktiSB/6dTyE8zaDwqMs7ISV
U9OK6cBxVR4F1eeVUGf7s+zJbikwXnoiDlVixQolqQdq7yqP4SWZhPdErpdL
uYy8y3r36jVRwEudBnSbYCnRDkSnzIbPZVXljHr8RQn3G+DH7bFrhyBT9f4U
AqnvpFwoefu2pXsvpf4HdLcEyCd/5ktZM56q6DVYEzxqKW5x9wufggfr64KG
x/ICjWPot6DaTcOczgeRJC5vYLSJWaSDWKCRGnQPYMBrqRCHX7HqLO5oSwnP
4q6wFhA4a2ntEVi8jkf1oh5DP4mOK4pSxzjlFQXZW1pVKP0hMl50yLjFSHed
CoBIIIvq2tv9YXK5XUVB/0PFgrcX9h9hKfPwd8Re8OgK0d8l1qHMzvjeA5Xb
Whz+MuwSC+JYmiEouHzN5wm53KWCwCcDZOw4e+QSw+RwfYyZt4Pm60ox9um4
fGl7zThSeWw905Tl/zDFo9pbZqTnST6rkLQNGnS2NTirVMDcf+FCVpnlpS2r
tWG+fXkkiqF3zyq1w+D9s338fPRA7MNOaBtclEuyy0KUI/IVL6C4PdkrAjNx
DWBs2Td+DoQU6XoBXyYe/LO54VrwUbfhPDa4sJP/fFeHkYo3iRLSxFe96yLp
xAjC/kLY9CgWXdAJsYCNl2+dPuX9d4nN2zqKRbP5rFZMHp8fq1aI1Pq0x2MD
kzVpUbfTCeb5MgxGZwyuXNNGPTCI/+Clt0HOUme8t0ju1mSA1u6MJZxmjbQ4
AiztaYdzrIm9ZIFI6eH4AyQ2/UnEQK1nhEFe3m/AScoy2VN5dhWdTCrGGPMY
Y5N+Wodrh/hykKUsP9uu9czD07v3MWbjeCf68JSfR1Swg/kbP8FuopeQWQzw
DjSnJkT68980qOR3y15DHIZPj+GpOuzuh/sovvV6UQaSn867cvAv2SjKMXEJ
eC0UvA+V/2QrSXKqBve5KVaHSzp7kelCAKiPdBJ/pzh5wZE/lXrdwpDKRNG6
X5PvDrIsiO6kiuZCJ4mArTw3juGfKl76wSH8zCimHYeFmGYUUZmcu8g1TNLA
8a6NmihhJLuC01vazPH0Bd2vriebu1usrYVX9iCj6aK3Werblaiu12B8HnXF
0BgrvZWOaNp5DLes/AYq2yQFPSZ3+uR4DK3EE/nlW4rZTxzl29L3hxnOGGJ0
VbYmq6xZxA+92d8QADG8URbRklxhycBKE8s+ykRv3K0CKwlwsIqKtbMxA0ZE
dvDQgTRwQ7jt4ygxKdMhLkEoIyCNtJZLW8MjGBJtdUBnx0xLaQwQRN6ut49y
BMugzg0PYHinBZZ+WPovXcx3GVyQ8PvKGEe6WAsTn9JzIQDYZ3+m9aIdbGny
r7p0bFfabsx+lusFs0F6EualSbNcnt/E9qGsDt+d+X6oN7oXOnkldy32YRmL
HuKroFxYdJanYXxCyt2lVDa+6ykU6h7lhHutyqpAukDbkJ/yXGJqlaaXBxQI
0HEvKuBTEbOl6/eSh8mL++ZzneKx7akqmSobcvz7x7CBZa3aOWrX+Ye9AIA6
3Pff6HhdRW2MkoFNiUt42Y5Euo/3YD5PLGt0DO3cOFurAm6Nv4GtCjHHXdCh
ALPWfCsqcdLQuWw8lwxcj2l56tyhrMcUF/mvi5F7OvHUepzMUdNaFTfI4tj+
nPv4YWTRezyCBA02F3AoTbfTA3ptIpQyijVRqV9Vv2fyBweGe2+vrW11/KI7
eKuXt+hYQPs7SH/hudaXFqFxNvvAsCiZwiyIM8tk2dROMSsUaUQHHaN2BuRM
sbV5mQjAPC8sIjSCqBiac3iPvfnQqioPrruryLWH0bi/r3iLIYPpUehFse1h
ObiCgx4Q4DCMGhdK0A/E3hbRPO4XxgCVSlyiJUM0iIaHV7GzBBIjYbM4rKEy
WlaKCnKZLDO0urCMUUmFxMnIVEG+NY11tuhIbB4FRLN2bp5zKdtKIu9Ice4Y
mn4niFFmp9r6fbNerfqf+wjsRI1GTAQm4UkNa7FTATicXtqyQhuhjqqB7UpB
s/JSkFi8FkfK0fYH6OlkhbNCQ1qz45LNnSqQJAf75+bGYEAFRIS9yOBKh3sX
9WNZ9V1PX+9l+BNhlytmV2xO/+IQsyvkN0tUsLUdA4qkWgEJo/X82BL0QQfa
TZoHFOYr11/5I/JXj6rPLZL816AlBM/1qUa5j9Ac1Bcmd2r65/ZosrU1Pp2F
cU2tOOQNigx9ZWfCdPyv1jBHqY1rGCm5IaRBbQ1niebLWFagcXkYdZqFDhgd
etqcj42L25RpmMXroXxdll/6PEOA4Wz/Tz85dJCQzeKHqYK1+OG0DFGsWpjf
EJar0KJL6hzCwZAu0/gdoK+JZCf5Z3AWHnZmwIBQJNw7l21G40tOGnTjMkF3
uafLdwUiG1UX3AMiKoqXU1b+n/dK5Xu87lu3YKaHZNgDjBgjVXFMTSFdD6UE
Mqscs1SLTiZReJLc36+SnoYN+/XB4fARf4X9Xj617MNDt4wCg+nO4+g7/Uml
zmEkfDxhisoaJZ1sEBe/7iijVXoNufuQGkPW4lrvnS81TBX1igjAXR0ed8+9
6CcQRDvhn0BOSa2DYRF8n0KbrEzLYQJ+us/qqwwWsotbUtPED5+kP+POTbM3
BwFqCNuHYEvzBBpK0cH9eu2ZfX2oA2E3NI1aKBcpcJ1l7KQ9StoeqfBR8/cw
3DjC5iJOZBKC0dfSV3j76ZnZ2dik96yKvx7SpnG60xUhOp5veAPqwmuozwDB
PP51o9vvMAYaTi1QwTrzLSUB1opesv4qyMp+ReyUyGIoy+7UqTiNadpzhgZb
9FCxWS3J5NbcTm+XC1ff6YwnIBY8u8xl5mpcLvFu6uqjngVRzE/5wsGfX0h5
soTtRt1R76fV+yfMKl8sFUrvTMktrjbeEY71Q7PyTNljWpsh13Or79T8XNF3
iUrx+E5J6DQjs3XmUDg+EHCzhLSgMl3o64gp8HBXERL/fI6n5UaukJtxcVRl
lK5CU8bD+wAgV5331vlVIFwl6SA2biVy/5bDGuMTRDlqhjgQ+DsclNebiuKI
Q0ybiN11icS+ZOiztuJW6t3KyZovu3AfjYo6Fw3ZYC1kM6k6BzyEM4MbIo2F
eA5MTfiG7UKwZyyW90beMYX4s/0F/waKQhT82Hl8uNfDDvEwjgHDGBBacg+/
OooWZN5pSsLqbSawnUL6HKM1QMqQDVLM1Xt6cJWVom9uUC0vO6fHW1n2h8My
aa90IOtMJ/bZanTOl1c6olPoj1oUmR/HSqT+KkALn8rvLhg5EWraLyWkZJZC
6PAgMUUJRyP+FgtewZASxWYoI/xx/H2KKL2eRKqsYGbhyZPxlieUcTkMLqnr
5v/h0+F1fGce3hY4ccXVUk28x1r8fT5dW8alwqG23R+TJKp0N85pnXzXHGDR
6F+pUeaiK/WOODr+NIFUqRuUwpsVUdW1WojW5w0mW0dj45OfpykmjoW2kgPJ
Af5BzMkLiz97Qqmp/VphM+7w+g6gyPXoYuYh09p2QW5GX0Ek03Up8uZf31Am
WL38j8+B0UTY4AdtILaQIDmAyxui7DfRrfxSZF+n61YjnDO2Cx8SUQP+RdoS
SguclnGg5pE/uyy3a8R1NnN6TXMj6gETSz2qo+CMcG43puC2E6HAvnsn76+E
/k61dFuIIFApy7kUG2fsSTLUtgyzvan8E2L053Mzz6OVYnpEN9IMkS/eTgOc
P4Iv7FK1qvM+ZspXP+6QhT7/g2N1gUiIh0rlwHUYBx4kHMn2E1Vp5u9VytTw
gA88eONITu7eUGfS7OFVoyoLbPvO1F6sq9O40qnH/r9Nb6e0yWSx+JvSLgtI
vapKXOsvf0+fN75p3dgnHerqZlTllnE8/d7Xf+u9PiLsiKR4H0ZXx6Q6QTd+
dqUWXS65N6pUpBFtt4BozxO5BOUGfCvscf3cfvCvgbp6EouEUIdqHZlf80vS
OcaJ2fCjZ7is/0J+b4FuDr1qhKkhPQ+yNrpapNt38LjkDuMI5Rr/dZswPeRw
AW+0rtAgj2XcGgYK2Wx3XKKCNbW+JAIS7WG3auEREnPOLCJLNlBrlyNQOSza
zwGQXUqHpcF1bmDO1DSptlgg9GYxCg8brsovlRDcQcPCpCvpwq+pDvk84DsX
n1mZGIAskw5xzEpvbTyU7qgZTk6lhVNSpkDY7qDMTdTqsXxi70DwGINS5XiK
HV7ZojEiRGkaGbyy5PyMmvlz0DG7Vx/YjgjNC7/hRLS0JW+Zil/+ppHfvmcS
uBz7e+uuNoxnI7YDMKOUuir11EKQ0dMfz4lV0dl4LUBEm+XFLXLTdcev4sh7
ltGHv2WBkPoJvhAs9HvkNLfpC45GdZC03Xeb4GaVoaLcxyK0I7Bom4GX/svz
rIx4ploekf8FZbp8Pem5K62Wiruyv7KMhxQ0EBfeEraKGrBg/CHLVOjiFx43
5/E9YRc0rJkGgK4e0SVrC1V1t67ieYrEesOkP60PMSWxHMRd+gD1d44cEii5
0Z11zFw2veiq4+aKFS41L9UwRb6WimyKUyVRUuWKX838PBRrLyU+1eMzoO3H
l9p8jm2G29vlJoDEbetiVq31ALCcpNT3NrvoX8chBuKfKtkrg1qwpOogxWqP
eIPkdHvH41Eu1XkebFhkecoSV68Sz8JYOjYUQPKP8VzVVDKwi8qFDlBfWBMl
JhYftXqE4PC5ATZLsmaAOkB4gKCs8j24OOpZ8oph6XX/kJ+2wG83xEvc21u/
XmW+MTSyUAZ+fhfLoBSavBLXNURxUp1EITzhjzQAOZs3rDrbTsFZAM46DkQw
yotCV6aGR8SAnDctI26JOOMc68po7kEuCyT8B2GnhxCEmwrwydseHhSyqjxC
3J+2qfuKER0p+V1hM75a+mYe2lNqHbdGx9501NpSYtWdQO9p3K0fFh0ksrIR
aguJC4p4fYARa6z8TtgN3OaTqJbPHHZrZYGQTfQDrM0+TsjPZH7j1Y5FPcc+
8wPb08cEFN0iIKDQU7X/t6toMdWwU3RE+4fVjZE3zufxKEiXPuQlh2Dc1/Md
pKt7wAhevluGzNA6R2mQCmVKj7DVRq3Kpa5GXrYezv2KVvRtum5+HTFvzXui
ZqVtkkNlovgxnqFn1+Gsg5M7RXy695FVMQ5AZc2BOkf6J3z4IAXwQbUQ5Q18
wPc+1Dh/OWc6ePcjHOReUTtJqASve7J+QEx4ZMbmJEJCjEfzL5NyvDFFXmru
bWmBJ85hgJLwy8TJsli5XPnTWsDF5yokNUjy/0NYPAKzWLkdRU5G1ohVzyDv
0WGF0Y4bBeAMNClQspDkqK7CAD8o1HRL0HCxJNx9y0NsqhYVkC8oz6J4QIi0
TCaCHncxoMmN32T++H58JMh7WVcD2tBuPBnW4AW507irX88EYqnsUaLPdl+U
xGc5GQMacoreTACBAhXRUW5tCQXHul5unJGhdaCv/M3vfuihGJvkwjAcVVpR
4lX6Xt2grxwOEdzUsQmg2VdMvvHYgdOx59kQZ4oPBBiV1e17iKerol4VbahM
YmKgf/TehZzxWBN1UkzIj1soEnnGjl3g5qyiGYx2bnXNHmg2R4K/6Qjm95Z8
cHUersOWHcI4YPpmnVY0ZR4DqYMxmnxhL5xir9D8vQCJydNv3on00/kTkcMM
JVcXAPPmJ42cJ6oJxFZqJ5DiY7uweaUrmybKdB85HgR629qFQYlmMBJWbik8
OvgLiAC5E1l5aKXc7OLVQEQz6DWVfqoCCNKBGdBRR4mMYtiP7zo68hKhwq/x
pHgByIxQ10vQFwSS0FYcehvnIB/OTV6g/pT6J5uwypkMQHtCLro2V2fNChJx
+xe1ybrPdiI5bCkT0ulOJBTtq3bGXo56siZS9amFyojzPRc+xGACMNizWkR3
tx+Cza+RDYSu0XspVB/1Qo44I8CG0xv+YQPJx+Gv7yrSeOgp+58uQdZjRlMx
o7pPI7Jb74cuwP6GSMEdEBYT9k48GSZlIw7fPSb3FoOMekog462luUDv2tTo
z5WVSPmC1LHNtJQQO8R9XiVBlQp+rhYEib1ExbQkrJqDfrnlqFTyDh2DCC4g
2AnADksJeaONI8be0fXYelJj7UiyexKB54EBlKRtkqJ6p7fahnjHtKfoyZ29
Lwe4ZPyVbQis7jMsXurD1SEITN/hEsvB6757FHemJ2EcNP++xdVxS7o9pizU
LPBO4HbQcqwuUXxhaqB5QSMh/2DxkjYcDyHQWCv3SO/60MQFo3CvrqA/ToVr
gORuh2tREH4rzVfC9kWFgqWlM4NsGnuVjI5cK9iC3BWuClgL04lxxmeFDCF0
D2cB9O3ZhszznGkJqpXhILlNDu07GIeh3B4em1h4CMRWj3bxmoNsbFH2rIgE
bsP1hWNeHxF4aSM20T4O7zsStQ7h2ttdHuB2s/Ge6s5c9Hquag0xkND7Ap9s
kvVnuE/71KTsfNDX5Zp+exzY7Zo2EalrxGJScErDlOBiFZ4fKIAPjK83mQLL
H+Xc77WyVhdYMs/Ekwe5ifYfIJ51BVteHVDb8K5Xh4m7PIhuHa8Fm022i1BP
/aoiE1qB2BLcoHnJ3xMkruS8V+ubHO6nYTIqBF3AcXagrhOvqkUVYiuHITDK
7gykQwAC9lt9u7jmB++fBf/+sRHSQ3z40V5KmLaJda70RiE1CCuW/VhG/T2z
Chi36NswW81Y3u+oisDWJ24YYTPkt3l8eNhxpdm8KKzxrTutcd66FSGpTVpr
nhc+5XGCTBcglbMql11XDlkiCwWrTljeb/1ZA8iA1dRRl5lre/mDY7yd1d22
htC3syFIXYzmTg8g3xjQPjZskgBGVlbm7QMLHQyddFJeJnhNSMKcNHhxNJ2d
BJv7zIWX+PI73kEikq1YI0MZxVkHfZ7YYhap51maVamCUlIXy/BgQWygi1zf
TNUekFPbElw3OPiUmPv+QKe7HVV/kpcpTWFTSo8PZxpcHG/jYWMJpqGD8afT
PzN4rTLLeDv0bmamZVIOK28XOArHbxJwUiEfuBP9AGzvGYjMe4s9S/44oIvr
cgV/9MJMhkrSI4GkJurkpcNdvG9AMHEjUIXfzwggBn+Sz8v3vTPEmHlfkCuu
GfZxe0yUKJb8QAvw32wPrg4GAhgoNDgR0n7L8lIq4lmdCflGYQZ28LaLe8A+
HIrFZ1PVFggy+8p9V0EpizKUMs6rT4BzeEWltcLH6G+WCBxtviuTB3epmdxD
RoTv/PLfv9jJT0BcH1/ECTfqMoxbEqezazTVTSz4t2/r2yE87BZcWx3Yv+v9
gWORbvYWwLujmDWOCx4SeuMQsH1GuTgfbsNIVDVIfh8/rcKJh0DSCooM3dyu
jvqbeH+yqC/yEXm1JYizDO5Ef8X1DQw75i+smVeaH01S5iHNW7Fr+QqHnK3f
pKYr2qoEsbAymlj4Bjq8Z6O0tvSqNdQ2j0I7iUyKE+rGFr7veOYwILfAfH/6
3JDccdNl0W4jEsC0oHkSHkNQnlw8S6VkQfDuDcUqYc7JX/1BrZZ8RsYlnkul
HJkYw57EC7NnNYzDHO916WLH5YlEIRzyI00/LuNIoMYRb6iBoSsefHfvW3w1
e51rbROw6te7CIpvVGJawe+ZjvjFiJAe9+PrJJo/2gxevoPeqOL+0y5g6RhP
qVoO0r0VxcJAnhXmzAGCbp9S42oYurkdpwNmeu4gBtrcTY3mnoKjqDUekHC4
gTgRCcROFI5hbfnrO0VTrGB1evVS1kFFdxtFj0GJ3q6TIT5QqfBddkvWmMdL
vdKImfZjf/IgOFHq7zLQLSsgAdRDIT7YJdXUMSNXT1g82z/NdyRZqI6QGeoo
aESaMmUVSqgyN6Q5XtE6XrTK99oZ80lluu6xhs3zfelVS11Hr9MX+fFSmP0T
+CH4nPKbvIOg8BNvJLVXG7SagHQEOShbg3KqYUrtFaNgL9YjiWDFgaclCn9M
lpiSEVnnnSnO5dIG4j12G/z+N4PINmkhSR09yw2mbTYoA1V7pVTukOrVfwA9
mEBX/ttLqdtPh5KTPGboWkmYm4IYPQ1xH0m9sv4BhDy4t1g/ZWJmVSVsFdwI
elJz1+gv+IZ0fGnq+gcNcyzR3JXpNanedYJyddQm9bArk9p352JDPlbsgxVt
5ucAISGywjH0qjK9nuSYNSjy+kaZJAUKhu7W4dshWPl0Xl+98NQTQ+/mfx+0
iq1bYXrk8vc38HTlCk8NUqCiQ2V1uxzOAxSBosBu+y/Vov3nT3OVIexvTztU
0YPSbabeqHikkUeApYuNUSKVLUI3D1eKaa/CixoyowYrrGxhqESG8JqIUJQs
uH3VLGFXxtV6s80uMjUcnYuNkiSoPWPwJYFvI7G3RVfgOEdCEXgCLAPVyQOA
8iJ+qoId3ptewVo/thsgMea2MCEqmIC+Jz3gmjw/dtAp2Uol8WoxasdiJ2Rw
0/5BfOw9j9cIRXqD9PPmewOAOxBjuLTZEl+DEk4bbIxhuGzE7PS4WAJaXtQc
+StllaqwX3q/Cw4u/+bmwx4cNaxBHkJYSJTP2zjjlBPrqYN13dbvE++WKgSM
7ZEa8oMsjxlk8a3LGkAmUP/nhtkeRjEowcgrACaRxIgfcfbhoX4A5vRa2gio
oZ5c9lJlXllTj1C2ncmGeNn3/IZGfncmoZm63+Boc49GZqxdl9v3LuWBCf9O
gPKNwZyqZH7raXETuMstGdF9AsFxYrg6FfxzGiMOO9GESbgl9oRyZRT3CuCi
EMIFAtOInIxxlS8cbrZyvwItY1F1s1LbQ+QExq/rYiI6M9iqOVKnQHVbNC4u
IIca/zHYCUuvXippJv8YgDc8oWEOkGaL9cRBOZBvV+7CAaNsVnVdDwVkDDbn
9J9obsrv/X/eFvNGbqJ+Ii2KqmFFGnHl18T3copzPpv8NDygcFgbQxBuo04e
EH1pTTDjnkmiKctrVM8GD4WuJZrwbw23Bv6x/4M/2KxP1h+7fFXlQ2O46Nzg
TEMcBBE4gHlnXSYFe+T9zdlxJliSN/zbu3u3v8flbw+UHr9N3CKzgUaRKlAj
EngF+oYtDHmcAGXdYJZjpNrr2BW3IOCz7nwhrNSeToa/8up3o9+9z5jlI8r/
mBydlHZuQvt5kBMG/elEEwwgAIbXjbMRacxKmrV/GBzNhjZjf+GRMtQlZvju
w9a4qrDp7tx772Ewn0bwjQSSTGlnst/QfYpqfcVAeEODV40eeoBwjSHWOKS6
ptIGSujVmOGgC4hOqyjmjGKNfNutyrfWVFmuIx9EeZmuBmsesIxYa1JVWZxG
FdxxWWENf43klVlXTrg9yLSyq6dYMQCOdPiX6juumJ3qIwpfE0fuRj7EJymW
uGd0mF0tfjxjQSsjvb51X3yRSxRYepB1VKvyr7AujaRXU9zYEwqO4FgJzbow
y81t8WxknrK74hBX/hU6GbtP0RpHs57jCJ1v7nueTMMGt/UFLG1aGN39AFK4
e9Gc1d46n8wnHWsCiOedV68EBZ3/9/IjwsKjHN4ipm5skijgSyGdtMyn1htA
V883axw1AggqitdzTMsmbwddmuNf6SC54pOD2kfdpwFlbjFPJ+AP6yHYXZNX
CXp10eId/gcEZGlccoadzFFiTJWgBVN2tvhRxOp1oH73ol/VAdzjPS2gFrG0
dea+2do2WnPk/rdJA9M8L8kmxdiAneIsYyFEf+rcrU0HVQqED/zuRdZkZ79g
LkmydwJ53Bge7hhpqJCfi2tGw/zIuaNgc8kkeLBYd9cmhW8BhU6hzGtMPDUg
fyqwV1DkA065oyPBT2QeawA2aMKwzng8M+CVG0zo7wK52buDO6jZStnzG+Vv
xSAuP0SOQ7qneIH+QmixafYuYAmDt5MdYTosTkGjxEHJ8ge7TRMi+Em4Fedv
/q/VdmOTo8B8areL5nAwtPgCex2T++Rk0sTLEq4Lk5fgyToEHJVw8bYICwK/
GvS6Dq4xcCM7IJhoFXQn5OVLmegEAvNg6AWIn5ayZeysuA92Cy3WNzcFd7by
Hg2Jd7XytHpu5kelwwvMIKzTqdqKz9w30MvOoyXS3hYGAYqaY5TJ/4BM+QOG
yZlNgWYPQJ//M9mFpbwK8MY0MFxmlyjrpgM8y6ioi6SN3l3rPasTe0cKMIFf
5/pPne11NCQaWyEVfJfrewtKjLk8YfjgAMcQd1UAKI0tlXhve5Dt0G0JclZr
xXv3TnpjjadilkJvAO3WRqlBynfUlij6HpL9zZLpNWw4dzLvdnAG/vvgoY5i
6894s6XX6zstqRyhI/ClD+vbLSzTzSs1mjh7Je58BFQfDG0MmZCoLu9ZyxgD
mVZ+XCpV1y25Z2QZL1GfooBG3dsNSOQ0nx/94pXtuX9oNkC4UkWhEKHb1vcO
oEzHHB3kkUWlT2Eo7SEYOhpSSxUWOSLp89YfTLkTSW4T2RTgLTwUWE7xFuzL
WEoFpeD4N+QA2xjCdjbHrrmoQqYUXjXvPYUw1T/NRCz2ycEBspE+BW6y4zLA
2K7xuPGDTOrR5xvREj4+ZMgXyGDSwhGfbE7e3QlhDbWx02pNYD9x4b+Zcfxe
sKvxsqVw393HrRFeZIIXfbEFIMVPOEUeYZfL4GYxU7/SwB710vM/qAVVMjHD
dFz8H6Iufu559fpB1nWdqlDjO4NhEZwwhyRdy38B1m7WjUelgtpgZS3lFLsv
2bU9WqBvEOPixEoaDkzPVAfNzjiF/hQfI+vtWAtu1vePVTYBFgUDYyhF+Ojw
O4lf0jgth5v4vYh5E94VgEnmVO7WKgEfQz8WhA8UsBZoex3BQ8msfCwzeDvy
87EoiPeN1b/mQQZLVy04Jy32cCV4ltvzWFfRxvQtBYvZJ+S6/l73N4QIGOip
DISe0pwPpcOQY16eHmOmEQ7DZVmrcy6tQ+SKt2tkSigKcXPXHlAkoQK/yr9C
KIcz4sxL4yWC3Xxl2k9kLEGCEs2RSmmUzJGnccvZNXG+pwjHABpDF5iJNVc9
1AFItk7hDGqcEDP020qTIc3+Wftjyh8NKsFhCgqQuHwXVUB8SRSKJyEAVaoY
u8a+GbeBZRexStuPiop0hjikGs189te7mRygnk4YPzJR+aKQAu9WGn5nlu7k
vBdeXfE5z4sunEZ/oFteLcJMG9OfnLkB/ITf0HHRZRuoeW3O0BsereUgCr7w
uD52b94RZiJebNnTV8OuXmCFM0WvWoXVp1l+Y2Oc6g+0ipvDCJL3xCmmlQQx
3Ft+s19y/lHPDhG809KR29NxmH0T7iNQRXqX6qSeMNTG5Lv8kf184hXpQq4o
2OwtqAEFE3OZAOmlxlQd1B/qCziUHN0WyQIxfsoPXTp7iyPMc94QiKHG/OHu
tF14BxQQ7NXqUpbf0i0PT3Ng+CQA3v1s++0z8jLnuaTwsay0rJ9UVyUyV/sT
kLNZMU7jd7S/GwgikkB9FJwyyB5TAwRWeBHCnsTpb4j+f4U5ygNK6QTVYqr+
KzAhq2ZlRRxE0xVN0MEsD4MPSIyy2YBCmJIXO6KpTlC03JQ8H4GSYIJIebJy
5VCQI67SJR0s0CXEOD0ApbeLXAGOXCPI7l4IigYT+evIBVhMxlMj2319gyl1
VWbDwlQEexI53xI5sqEfL8c1JLhcgvmGX/bfOtky/O3UCS+rLgN/vO7qqRML
56JDfLtnpVz917bbLkvu2Qi5KUm8IJudIwRcIGXkGJ9hliwlFqzdCBmWXVSf
s62Wavz1gl2vRHTeif97qsELPm0bUVUpwHBcxUdmhHRC7BL00wm+40I2nnf3
9VYFaiGtVFMyrLIplVkut2Yacgo+V7ujPkZ6RZ+tk9JzkNj0S0qMby7Da4Q2
7BpNzx0UN6c8Aw+cyidDQ7J3aFHPsZGwsH0lXg+RAAG1LL4dD+eeERGFVDRy
PAyFAotjRSVbQ1T+5R549whH2f1xbOaEUSTKcIYl8JFpjAWFXFQ4lRw2C6Sp
DiInZgJMZz3HzCkgSRMg0UdIJcVo6zKbh6maT0U+4e1b2JbLWxlFQ9cj7Ub5
e/kvE+EVSUXldzai8C0GTUvDKpNu4yAE0tLenWog+MgkAlxiIrd3DBEJAzLi
lLKgsX1p7I7VwR7P3v95hX+BwQmdCmpTBx5Fttkod2GlH2sufypQ7pBYGw3M
SLl1H2KPMeopIKZtMH7EFHZ5HzLILY2WN4u/o0+Q/LROexfTGSoknYGZUcGO
MDeZPmUBzq8ApYDd3oSGspNfoWwhytTnckdewXJtek5zZIxW3++WlpWl/VAh
TwCeQJRreuQwwBQ6jqOyHCObn8TAlMd08fYkT0K3Hr+AXxWh71U1mrvL7Jks
dLHsr+ig7RcD3RP60uDJLn/tX4jfmWDiteBCvSkV4EPyntDtAXbRxZL18qzf
rDY5ylFZ1GPKNyCuKV/awJO9GpEmMDT9Sce8r4kB5tz9ncsdi7rZAES2gMOS
aqbCob6hYyQa902uWERKzdbkpNHASQwc2RhPqWZj5skuMPE4pKdzphHitAg8
D4apEdGztS4nUfPusTGymxgKeLCqm4V7HboZN6ITqXGYEErWsIA3c8qmt7oG
iITewYf8bqahaNbbGA2kEt8RklnIhRyyN2KEYLCwHfr4MSuAy4XDq5mCNdSW
iiFdwIkuhI9V+obga6cJkVtaJ/72jqvmtOtrOA0JCszy1jwmTZBso813ZYGC
oQMc/GRYrL7MLTsSrA8ENfsdCRlCRok19m7esrySy4tlarozeHn4rXb7UtWE
vstJ5aafrliKcF4pJhK7sn5U+Fc5Eaelqh7msTC/wg2wOxwcidfeYciTXAzq
4wjt3jffYdQvBgX/3ly8n26ugjP5uVyCHmIQWHIRVstuJCj9UJPzuor4AEL1
1YVli4OwHufRTMOsN6L4tzm6LsRp6VXLXG3o+I63dHpueUWccIf08KtaJ3L3
loyT6Oc7gaLV98W2DRR/i9tX8K2a4hzGwvilcESQ7k+AxilPGhaEZHluKQuH
k/mqxV/XBQpX2jQcjRZ0j+RGIqwV8O+8NlZqagLYLHCd3NSZ8ulAq/9Z+bfN
8z1h+GcrZonQ33Ry+MKc3IlCznKmZkwJAk+tVPxA+IWKsxx5w+OD1tk8oxst
UE1RoCcbW/K96oF4oT/SU67d1OGgStapYxc7AE2wZcOWab/Arr2ao3zEJME6
FsXpbgoI8B8nvGwwvf3UIVJXlYqREnQrLg78NaQTsi7qOVhBQzHNH84HwEyn
TSW055/NU7/NcsPWFZXzSoMxN2TVs1kWmid781HafDo+Od8rMo20k154JbwK
sAJRpX1CJCljqbHP4/Sah8+J9yRzpPkXvesFI1eDI6ExSLnDUuUQj/G5+FU9
HEOMsu4m+U/SFuD/53PptmSscArFHRhvcYotBb+s2xoxUV2pGdyC7JvaO8wa
hB5kbZ+jG1P1GVPGyjD3iERujG6sFB83Lh39OL01KKKsoX+VWkjbaAVSOwV1
t/FVtCwvXRdLbOEp9uZNEA/ZYmRGTbbdVGiF7bi6LSmfOMFFmq7lIrTuKYre
8xBEEvY3nHOONu/KxKwKEGnvSNQ+oVsUROIvSee75cwaU0K1eV1eqqz4y6Cx
fqUsLIE9OoyVS4UCGtoyxXsgUyok6WuOliPl0nwzzK5oTZxG2IKEKzps7JZB
a7lPQm5YMTo2bNypOx0D8FH0m0XAdi99irm7ws3g/I6wYW2bO8Xm4lW0SPUP
1BIAjYXdb8v3nuAjz/hiBna+J8sbTvL6VjEx/iuc7kml0DuSj9lzJcZ6Nq6E
tlKAI/qNfXEgcVpzlYy8iEYuV1ePy9LyN7Rme5omuCl4Ay50T90MeE4SikE9
qbaftIf369v2DmUXnxWqKqEVBAEkHFvnE2FJaGBI1rldzqrH7JTVqNMPakFG
Vyahxu6231HGRj7LeA9euf5Uk77Oy6zmwtUZ/g0P8wUTAZRB9SqKKyGGlUsr
/NQ5i9OcCkYLFMypBu91c/W3dGwh2YWjybTCC5DFtVh5ITibQW728fgzB8Dp
13n3JmGqUiYjEkKjyG7FeM00iwCT5I0uMlStcjAnafhT594uqn3HL+5nb5Na
NRiQHeChQEujFnVnkoKM1IV/gXXWSP4LiLn3hHXg2yz0WEtvICr5gYaeySvE
Gs1vUpTazrsucE9XsPuq2GdMnl/uiOEti5suMEHLf5RhkTiJTdgvWbHI6zX1
iKDbweBAJEghSDWv6WTkbKkxEcBsf+lnGT3yOigc9BpQfcK/Iy3XIHaKKpD0
T5t/pdEYJdNeLH5J+VROvRAYN+DBcFCuQRX2K26Zg5i+FsgiRYL9gff4mv2Q
L76eMK6m4gx/xd+jcPvYqhB29r50ao33D2qKl55RhCEXxZ+ZKgblrOMN6s80
HyZrL6KnZxJfsd4198sAEcc6FfRg4adDC5Rp3Lm6bVXRNLCbh6aQZ6fSFW9x
5RxnE8PO5WEx1RaZGcp2jcQoBeQ0mxQSEt6JAQX7tGBTwv8soAZ9qIOT0bRv
8q5uypUrvB5eJbcVAiC0dwlc7srLkBoR4uHMU+BfNA8nu2reHhPiQX+UsmCt
TosEQm17LBI3MwwLF6OeZCPqb6vUhZp0yS1NhL7/Qm3s632EHq5wYx1rCr3A
MqqAHHu4cdjUgJrt9M3vMsuhJqERbIXF5mwpVqIpXtMqrsfUlIodylChWK6p
/3z8WHUFc8axiUzlfxVzNfUvWlGW6T/uEOSoz0q0dr09BI8NdrKwj+SIW3oE
0c84qJTP4vLave6VW6t6rTlqe2ITue/qUlw8z9XFgiJaCm+ODEDwoNvdPaOI
0oHWO5qASlCVR/e0tD5YxSNayV9rifgq83S1XNU9Qcvl/x9wLblyruFjSu/o
oXnHrU/KYB7yn1bgfHVVSQ1XNP9t6S+UsCt/d3E1FWMdCiM9U9TihVv6De3u
rSThfIgSZofQtreHYjYVFiILOMI5rep2/IRdVcXK1I60t1FS3zCCnBsnn8FI
usnEWriIzxj5lCSqbYbAVXujARwJ1kFFBtfmeaaepAg+hmYTc5u7W7PnYNo4
NJZKS6QgdFiwjYx4xg9zxcu46MoJBTNi1aGWiaSHjZyiuRI6fKQ44m08TLSQ
iD7HXHCeySOwTUaTNbSWGbKu4wlaE+u9PJIEIK+kBSVPxITQ/ebv1amt+lhf
nWmD45wYD23ciJaFvHAMW2Dajd0nK3iod+2EchbAdcAoW20adlfWLRwM3ykL
KT4Ghy4IJyZoqweUO6Rr9qYjF5shy9QkBizq+WvMFRzYK9s8TUQrScqbeoP2
034+zrui4YOs++44r68eHenBUgAhh4uXSgpUzBIl8+860HalVvpKypYAKVU0
jIuP//CgkKAkQoxOM9yMPXtfYD9A/IehCRw/SdWXRrdIMP1TiccFJyQQYueO
3l0hemlhbxy93Safto4iUR8UnmawzX2qjqB3PkshzfWMj5jPBQf95FNncvzo
yBs8SjuFYWpkjaZtAAzQ4ltE7Gg+a6XEesyqk+HIqgKiir5CACfbhJ/76UM9
/eAAJRmv+UyC6JExh+SpV6xu+mkIKmsWmuhhiCHQ1/fNwQKyskM17nV6bxi1
7S9ywRgbK5MUZEHjJUTNIJ0jc77EjjCnj0pJTb2BDIeFpk9UXAaiMTN6dI4i
InyFydj6dpKBT2VIumtl3ApWBjCZoq1EsSmJsSX7ItgzCMB7eLEmraHqHGfD
7s7EeDNCrgnMWoPprOLOmfEf/hoTTaaPDzFYjdHovoOX6vHtYxGt2zWZe57q
AU0gprQ0122QXGFu3yI6Gpn5AQRSvmovHa5YKm9RBd/0xFqii9Y/iNRoxMjq
sexYcfo7DHSQ7cYS65Z6DUS3/2mUKm6CSkWtshn+pstHLpnkX52Bhhl1LqZp
87X/z2Bz5neuPobl8yY9mxdgmJbafL4dbAty7L0M0jpsTxYE6yL9Sflm8qlT
LNh5facup2a5PYQR1ggCZ9IcXoj4oF5jxb3I1MTNUKmlPvh5S4jxNgf8iLla
oCvz81Mjru+O0KmR/abykq7r4z69PkmFYWEQAsBd0cuSKYXffWsTlieH6teT
qnl0n/fCiRPd/kpqdDJUBcVqc3tHQfjEVPCqi8qtej5g9RMpMkNszwsT9OKP
ET//laK8CxoVj2V799wiwrgaqoAg0oFCs957vXQdSNPKf2C7rUVhsbObvA2u
FV1uA8K7zLJtrDFyZB4lGyUbO8rmQCumPW6c3hNovHOoFYko1DqpSaj0d5be
Pbre/iUECobOK1IrcvBgp181X5dmXurcKRHCufU0uXbsaDfr7t8PVynhQYXp
nBabnDQr/p//i4TM218TmZXdqECvkot27dr50/hH9QKb3VpR1JOcgLCfhjsN
djS7hsFTmOxb3pWJlrXRHRi044AnRzrMByT6TdH+T08s50NU23m4JNlKUAvP
7uG+CTER1nM54kDu0rVmJhe4YOPlyLbunuGFJn3vlO5VDpA+l7WMmGFH5ZsN
wMer3XwXyDqxBkKp2/5Z4PvL3kjx3/UOm08vNglUNThRwqMUXJ+2tF2k+unw
Ts68cOKHPhHVaQLKg/ScC6F5cmlrtM5CrJs7dyvi9qhB4e+J29yvclagc1D7
oVVLXVwiW78fLaUGwfW+JMqrTkDdczRHDpILy55BW0oyBuNgCWiTir9ApxHX
3I/yCuky2d2d98pLn4MQm7cHlsXrZBV3cb42+Q6ks4gJbVvbAWv2SaC+JnxV
fqax7a+gs23++6HS+y0Km0fbGYXJREOuEbZX2vjMFsd01A5uUbfT99jFT10I
ZwS0PZcnS5yGinL/DUv7dZeHDveY4tfksnSyj8P1iL5boW7NcR08DXP0bb3z
ZFHcy2KNrHc4SdbdiEqBrCc4hQ9Q8ODeydnoHCqjY/z4y/qJ+qBsMjeadIZJ
pIdshz/rLUcAhe1wbuoP6ZpIO925OqU6pAyxcqMOtr1cB0Cnr/Emq2dyjJ3z
d+Xe7SYxgdqKDE3bfEDMQhB2A04E4czXXS80nPVIGqayy6DgE3uKqTu/SHV0
qgK/ltXwGfaMdc7bAUxme1qHPIWUO0CMwnGex9XTVkixTIsaOyrPnSye4feI
6T9YOjoCS1CIq5G43y+FWgHmpocSMsZYVGrSKN1rk7GeI3ISIZbzo4PGKGyJ
hkTK1GlJOBtWoK4LTMMSmWFSvpSrTcvqdgCASt81x9qz4M8W0Rsgyx/mHWs0
B+advHJxx2HvRK6I5K5/TjM66Gclzy7fws1p+IwYaEI5qxe7cKCflcXDFMc9
ykFMg4a1WOwGPOnAkkVIjkIJvMnAv32OMC67zVS7NgtughObdu+RM5UiisEg
tNWHuJ3S3QvshmpKtRrt1gb1u9VNCpDnhFazkbQk49aGhBynnQVldcSVhNm+
H+atGhIY40EwoBCtPOGkjr9LwD1nqrInWsALnLKaKpdhoy6h+Ncbynv0vwoW
dx8s7QC0XQsMeAW5T6PK3eOXD7CxY/D+h5XuCQXQioDzcoEzevNneFDZ2jeU
vQOiINWljBx9pOYhn9+zXccFyAo+XRpfnkdLprJBYyonR2K2BVQBJ/9uCaPc
50Zm4VWZuZHBbhHUSeQ/Id0F1pAPzy8CUPLI9FoN0FOyGhD2PNNGNsoGpCg1
4Ub1He0uY95QmeuyV/Bfb6QUNkekzxZC99IOHtUQWhTOrZl92E9qtYL7TcvM
YJalbgIsRxkuoX0aHaKt+t25JacD2w4BEEZbhOJp1Y9oiTWjy9LPwIWQ3txF
SeAHDuJMK5HKNe/TXzprgD0IxPZzFqZpsVZsb6F/VXGKmsWiZtmThA5VZpKj
zZHktpoTbBsTZg/9E8YckIQcPoCqa+xQBnyyeP5/tmjEFZaiOVuUHsVqz+2h
EJwGIeB5SUojivTi7RIXU4k+SNicN9nklTfwZjz4368cS3wi9XDuh4+oUvTu
CNVSaH+2dOYq7iDg/pVEXxvocahu/8Av9+7gZSWouF/2JCk41RUy+o98KLDB
/UcR1NLJAS3FMs1e6uMAMmVhJ2qDKtDdu4oiAjIn4wjSVaF50tumrsXcrYuX
o4+rNTvkMyYzlO7LygjRGEnValB/PeGogKVyafWbcAlEh0YGlOk820O7Ok4z
2rZR99BROKwyokjdvQ0pZs5oqi7H++RquGQ/4IL4QZZ3uK3v4okAJRmOlFKA
Ze5Wo6rQmpqrD6Md9gDdKjw2SOK3mxwV6pY2Iaxwd8Vum/QuKAB6tqr7oJbO
oY5o072fnO51iaDx9o6j3Q8pkyj+3Wk03YDk8JwjPKl0v3u6BQQuy4P68f5g
7yLVCsiBEoLbXNzx+co1HjnHzNSt9YOFlwSCHD7CIdRAAB//+ohUM18Q0FPu
oP7uiwxNZDO4ywOie+cnt+NozEifrvi5TGg5Xz4OBH++ZJvJ30VDJ7XyuCAd
is0bXzU0r1L/g2qoRZQCsdxLS0+hOtsXbIpTL4RvytgOAEJDOQnhtR12bF0M
gJT55AgAezOT03JHX8ab98052uiz5AhBzfMtu26Itp9tEB63ceCgFC4/egZy
1xXJ4n4VveVKxTL2COnJ1G2nopLPojMyY6EvFAUOWLztZ/LDKJLbqAUma/Hx
bWhvWcliOhwCZk2TcSCcpozpyCqkkqbxWHbeAzu5hEpDyoqhdPUbXcf8RxQa
Bi5tGEOdPnIBdB8IyBpr/TSZam8BtC+WV/eakA6G5doqms2+ZA0tJVUL7vP5
HK9+QZm+6M6vQASKPCb2vTiXk9r3AlzyRT9O+eUbt1VBKabGDz+MUps+ISm5
Ubv3KK8ZKGVL65Bt/+sUkBgYwtZNGjud1nPi8hzfwGT7SK+UE8lKaKV8nbtb
LOThKUH/Pc1OS6DM/cb5fxkaivbenFfOABCUa6ZdmiP+enry90tkLdC4eP3o
c+Y56nzuy4ufcQ5lScPrZYwxc1ua64SiiRvXgmjdDOqkDl1S5Jdaw2wh4zhd
HsgAkwmvUednwA9LswVayFS4PZ0PbF00s12XJay+cU8/RMZBWzD672R54Fm+
eem04f1KZ2P+oEGlw12d/Zs+zhBpYNDfI3i2JNFfBgpNHwFmRjD1VQqQPoO8
Pj3wlfqyvPVJ0wv+r4/BN6M+GdZ1KJHOagxreji7FISFu5GghS6FbNPhCM0q
7vqw5AR3s0X0qVQpKZGMVmi4lKFupiyrqBVQqMOzIpJ9FY+PivjcfY66mOTr
qXsYbQHbCJa5YmU4eKpKP86+EMi1UmQlToPycelrhvZ2R1RIB6kaV/XTNSlZ
Am2x6p3l2rsNF8W4V6+be+Kst8cQTlxLhUxRyrmMFnS+IokOTIzPth+cipmP
d/CPBkEf/B8DoL35LxeGX2zyKALcOflwkhLtugkJ/NN7RSywY1HK2Tisufwv
ZXpNKIHNqFOI4n2co6lUoezTFttUtGQy4n8UvbgqUDyq9//J7ugX+Zway878
gG6pFo+jDu1Mlys1vl5t/99clHedhQofVAJg5EWGBOii7ewdT2w08J3j/Qci
11ZBH02K6QPGX5M1kxGeYFFGvIIPUDkXI+wupeURPjX0HnJSvwoRWKowBMAt
ja6Bgv3FNYyEg1rTMiGskTmCcBfxqls4vv29h4UCNqbp8UfW2tA/fyh7Tr5V
heH0rJFvXv5uLXnXk5DVKqNPnxsQOkM8cqxYlpWz4mJkLLRSkS5qDwrapxi6
uXjo9WuVDnDIKGUBesQDwm1etXc6jgfEAGvRMOqCLVYxGWNHEmLzl6xj2BDo
pLvmgiWg/CRUJYltpjuR5e0ZX3iRFwy5xIgy1AXPY/POnoZvEUKn7HPbdgP9
+s/NjacVIHYmC8RFYSJ8rQxF2Y923SnkTIvEA3VoZxeb51ojCvLsiSK6pSJh
w+qeEYYf5h6a/FD1MA860hMl3dVv636l7oSyUqnS4+0+iDK0gmAEEAUhSMlR
5o5+ZF44UUBORVWeKNXD5E15n9vK9Fsmb0JttWwa7YuXXbBC8IEr4z4lHIGI
/tNYlzHSA6HqBfcVg7qvcWdCvReDX7E8WWatfPotX+8rSzPWbNYvxrdzq/3j
KMEoOjJckglis3jjywbUuKljp99u+5rdGH98H9NE34LNzN+tvPpQEeUNWtzj
u1uZ7N64A9BA/lma/D5JSZK7NPcyMOUwgB+9HW0Sf73NBP5hCDO2lucCTRDA
pKBipvnn58U0sHT/G0jwujTIWtB9OR+rWL0qN2nSYBHI5cw/YexNnqBxOVii
WT4FB/Ow5WbP5C9lzUvpX0uBa9McKxXntDH9NCakQbOwMUyKFAgDp5IQIKb3
ybursLgXy0q6Z4Dw7vloe1Uk5jQ3yqJSkhimJ8X7Is8RbAWiv0GjVc9qknFW
euXjd7ZQK8uwzSv/VnXfB06nOXv+rpDAnpCUIdJPWeMDKI+3XXJ+dC/psWml
GnziFd1Q0CLYsk5a+OdEiXyJKMg98miRUuYEpycfE4XMuDBsHS/aYDLMwOKV
yQhSAOpPdry2jx6dZFSTGoq7JIRucZgzr1NEQu27d+vKDTvpftgwwjuIWCpY
iU/thxw2KCCylkXjZmglG5bCGHw5gA0WjnoKE+V1RLOK3yFBwpWFFzCgym0R
v+P5XPpAS8zcq9e0UgKr4JlI4EslIDm1LUny+j63mD3/Z/YJtz0Ah0MApxBk
6PFppSdOz/ghsWlqpPA46BeM1irSW+w1PV6YMRKNFYo64xhIT5brPWNDWOOA
oy9Mp4+SE9Fk9ghbELaSrgd1GOoG4BIpf6owuyAeFtO3Gc/oP+gdwrG7ZQxB
KemWQdlVjRNH+KQZOS58SfXpyRTb9yG9Hy9zOoQCgiBVJQbwjJDGbXncdJNn
n6ZQXkdu7C2nKHaTOvlmEtKiw8qwR9IXz11r+Vv6RbOv2oyqghkiFxATYM4Z
tvbCSDdGApCpVSGSo0s95IsAUJyIAQ1OX5Oo0OTyJPxLAXx7BvIuPLPNz+rB
jB7+X7lf7Mww8EdHNPxpK89wcDJxwJTPCmFG24iK960z5f4p7AV0643JhekE
M1xHUrfejg3E6xy5oSt3t2ATS4a9Lv8QMPGY+hbBZrbTD6DOtXwJ8gFDZjIS
DuSPD8u9/Cknwm8BS2P4pa03xwKCMAIpxQQOF2bzf3VQnp5masaz0LMF5o5E
RYv7p1qip3YiVx1xK41Ebrx+qzQ0cDpFJhYDyxdd01yte45QZ56AULNSgypt
wY0jqDmsAhMEZ78/4UpsZ6hscViOC1HNVKqfU61C0AT0XTtfd/8VQnBk4YyY
jKxzGj914NeaQqYntzhvWc1EEVFDjwsLVuFHtB8tfDyKive6QNMj/29VTVUX
SsR64nL6tae1zrYsLWM4lE+tPLlw6y44t40KX4Lv3k1G3ylaZupRUPQs7qXE
fLUny0H/p1K270LcWQDYTk9xpD9NN4DNmZ5a8WJjYPJGdguBJMx9ixcGZghy
Q0EM3X7ZNXgFi/n5W/AfxiZ3mQ/AgWrX+FRDfFWJ2F/2qlPomTLkAegY79AR
VFOE1m9sMhJgFJ6AsSHD4AbRfDr5LD6Lu0/hjAb2mquDwZ4VmWqMC2YecwoB
xPe5fbFEBvKcvQ1EkBeS5HKW3G0USpKe1uRWiUp+txdR6B2uAyhytQieT2dX
CsOF/YNOF2RCfOXKC2WwH3H67UK3e6jdrQfp/u27EY2CGTn5FuiaF3FJziAV
Yh1ZQgmOyDkt8Sibv6xNDE0PF2mnJVH040GWgXpOd7aBhIIPMtesJpy5wxAO
8ZN2p4tnyZvFUh3gtgCy7XYSeBMw9PqpqU1ugA6IVnbeJEFmuy20LAWEsQbv
6sHE89AGBR5mQfO1ZzGjvfzt8FqvH2anlGPO5WO+fIuDR/c3BfuZnSdfGvLd
MwDW9JSCwoy8W4+98j+Y6+xO5qgVF1bCOX9bWBzdYiStvcp3riaejphcs9+x
04tCsnDSisLbTt55atYuvGRHApnNpfu1wjLmgy6tfmSKpgWi2hC9bA6/5R4+
VoUppySTXZF4OnwBrqetiaQK+6uxiDVogIBFsZw5Vx0bhg1UH6XQPfm3RbAM
s8YwOiALMDf0QUOhkl8/J5RmL+J/9/KPyAv2c8WPTkYKAaBDBHjiRWdjhWjS
ShAB+fQTwF5Gx6hHP/XJRZHT4MwsugBb4s4M82emR9Vh5XrKR3djxWIepxOY
j4tqAJCCKOsu+9oIK6j80yDsoUKNJQD77yEzgt5aHrYJ+Pgp8R2+z2Zpp2RH
nyjn0pAFLnIMz9+8NHJz1bXOSax0jP3dk0jt3oN6NzNl4a/NSX1tn0rccLsX
hQeaw/si3Cv98MngQY/y9tMoVT2cluAK1UXXF+r3LhqLQyAGrMj/unP87T0Q
z2pDgSeMsY7xQXf/bQ/eEuZZrQdxByJT3s3VVliq1aLe+IWqHfc7at0u+Ccn
6NFTwyFMLSllHOaBHfPkno96DQLftqzBV8vxkyJXn0gVEOQFTOvRmYcOXwj5
BUUUKHbuodI+X6m75rIID9GbIuZhhS+i2/IlWCH3kmeMN+5x5vK3XgowDgKm
dPptxnntrGA5L/eWhi+mmUmRRg8EXgVibraSA+gXmfacudY2hb65SU6BBmTK
5ZsxX1nB30oAN3gyCyVw+UZGPZ8vWf1qxF82e2pN0kISICD4XYowmtbxHSo2
kOL4A2VG5ulTmNmSOAGF7nlrJvmM2zoZfrSkmYQLZACFieyZ7a6k1MSmE52v
kaAOBk07/5IvtqZj9+Y70LtJztY3CEO3hrR9Y4Gwxt7F0WsHR+DTuqUkzh3Y
51xBioDWOpNBUOKnJiV3bdIEdozX7LkgqxnAftDDL25UOujrTcfHAl0bZKZ1
z2hCebv8m+6kHOhg2LKGY0aiWQxDune1FjZsUxC1mFdmdV1TTZ345EWVTHph
hZPJc6EuEYuPzJmS83/RkcVZrcD7gVQf86FY455RalguRpJL4bHhkj9XjJ+G
NcQDGEPXevPv01FD15JNut0Nikuosdlxz7mpDJqoYEbUkFgDeM27ag1ynsiB
yEjjGyo250w/pYvtLjQBCT867eVjuTuzxa4QZ5QbJg3twA+ZNxKhzZ1NrpHn
XvWJE/BYLEypYsOkVi0yXmkjLjxuvXxmsTPdXuAKdcl5PGh009EODpmX4QVG
3V8YUOY18sZtDye82pvq6TLSo+eOLwUg0lItQocXPC8yum1wLJMUqmsT51dn
MgguCl7gzCZaUJGmM4FYNVTPbhDyiy5uzmjDJRGlmj6QxsuvcyYJWd+Pijuv
AaH/aAsSx7Llr7jn2Tnd6PuJxxrlukUQDENtaT8Ct2ZeBwTVC4oJmZn2/D7d
4/WEok224JK2j+w6Gr49o/Z4TEprqBreq35Z8UnQDldAkYGUxW+LNZzl113l
jWVQ+401EpeyTGnC8UApYBpPJQumkzaWCC6YHo/Td2/CAjKtZAowFA2KAwBi
Xwc3Xxn2l3Szh4MiYQHU8ywfXIF6c03UTwYjZJucsz4sHtIuMznvH6KBa2Mx
lLQr12QSTQPSQY5g516NSY9FltsOtGnQ6yHwH6b7D8MnZ0JtatAojnvoef1Z
o7uxP3sZ0GlKDD2iX+s5izkyj3ETNC2lE0wevce6zPJg0T198WPOYZ+jLZd+
xx/X+5av711RNHzFl80WZ9kvjqxHZM8DgPK8OQFyvg7NGZuSU7yJULL8QhRZ
hQcRZNwt3Zxxu3fkjM/7lXhp7NuyDrzT0RvDcMVDwNFWyK7IOouQc2QMQ2Om
swB6yYcbrGuQICY19+NxDjXRkBiRlH6DDyv4ebd0N3YQ6cRRN17UCKLcior3
duORUbcHjgtkewaN0fy87ZBO7lB88CfUsp5ts464xgHkl0+2cxXjPNWf777Q
5EMEIsL4OwuHE6uPB4k2FwO4xt0W16hab3XycuRvqoIj/NK2lJWQ/7Ziu0n3
utiAUw+xGAHrrDCKTPtZmYiVZOMn/5EvmIpr6ZfJ9yee75ZOeO+eEe8T5bMt
zXOGMe2PG2TIdqX7h1M56UpSVgBXBuMyhCxzXSKX64ELrHoB2bNOO/8TQRVn
JCc11kVqpC/xZ0aV1MwMt/jyBcJKTmcvIcvX3ZWBY3bF7G0LhKiGOjTom8Pv
b2WGhDfhlrp6h93WZdVVtB7Ye2+clW+WXk4BljGuZ2xbZwEAn+LPHWsOcooZ
g/RW1UHeUO46kBdOEiw7qEjLoNA64RbQaK7I4iKBdX+BBbImeRIQiqiKWuSW
gAbMAc01kg6liUSwR0rw9kP8ugyV45fkAfDoz2V4Aswho/yvVA+Z/Vn8yzoR
h8J8dG+k2TgWLt2Bl44ZXtRlwtZ34RYjwBSZLBg1TCgkJlsq6+iZ5L59DZia
F1kflta+rvwvTBlAtCS4lgd0mtkIRoIQrZP9aorD2mhchtEPeuSnzfy814lT
8/ZWZOYP3XT9NEgvu4rB7ahadp+Rk3/6nLLBbf0jUr/fjkCbG3X3hCzH5K9t
bXbHre6nGXOpmr5Cdb2848fZiXKXs+wHEX4WTNRBgxrrMAy3IXluQl+i1BHJ
vMEeu1zVJvP9vNdq3bvDQ4nTtttzmB+cjbyOw+YJp72lCcel3K/CjB7LZ7hK
ZyGCd15plWR1nZkPxUOpOXf7yVWMC1fuTlpUUh1iPtJGP3k75klW0plC9SiE
iOAD6rL7EKDnx6RWMuOp9j4AZzXBmJ6WqYEd6PDg5uuNovOlViRL5ZtsrDII
8tVRJ+wdcc0HX25EN4hbD4Wyyjt+hhGoapJ/B44hjEvWkvL3GqafnlpL3RaU
8yn7ShtxCgg6tWBUgB3NbvTT2iOgGUNoN7GoclIAqSQT5SADenp24TazLGUw
ewxuO6lMzXUyUImkShVlT7JhSLIG/1PudOieHz7XOGCAlyutrknQKIkJ/GsA
lEs/wE6FEeO9JueXW1s4Eip/1VV0BDnwRq2Ku+HgHGxn3IepIyidWEpEjcch
tIDftvPyAvYFClNy0It/41L0vJMQlGG5UXk5vBwHn5zcQGnsHscWkwDdA0d4
ZSODeMLZnnG54QuyJ5BQ+yH4s02alKADfZB4Tk8XQnTVibEcgQOTq9LVx1av
k9U8S0NGZF7JkKXcDkUdQNWA/6pirLfVjeatvtrYPukQO32dgnbjwod2Ze2n
l2l3AKjlz22H0K3gcg8cX9MSvKNR39GU2nZ/+xYPTq7aESx28iOaX+DdSlcI
Dp0cXfroPTn0UpzJTTqly8CJRs5Fcf0yjfwI+knlwa3C/AWrxEV/akoUQxBt
aVj2v9JzZN9TMb0QwgE4LHgg3jjLKNdprnV3j06OnKEzwZN1fi9ipwLNKzEX
EAhTF7E9hLDb5H7h9IkBEGZ5kpq6ePASdxFCX6sCpC1ozhC09bG8b6d+Is1p
0v/DmEn6kZViO/qduXH5akmSwfEsgQkLEMNbEOZQtub786m85YMXZeeBj2qs
eEsyogqHEwA4v1TgyCAND6H14JX3sTeQnHk2nfGaPwGr7pIi3hvZVHwfZvL+
D2SyBfFjVrUgrNEl4wKfLzFHiWPsAomnivB5d6sAk2kRJerAN6QJiypTA3YP
nSOBXSzqxEnLMfCvvcQA5R8eMEf9WVLuiugGsK/Ii6KsBZVGTbIFNcNAZCQv
Yj4LHaqVeJNuP06s6lCozbm/Rzi56dAZegzkXaDn+QdhsnxARiYaU3cTt8Zm
/58vSWlWf84b31ca5pxga6d8PXPIl2SRFch1n/5Pq4QaYMFtxF/KtDafaDXz
1kWbflAi/OrltiPBAXHLhMOHDQQOB/8+fzmSeu0ROOFvTQ6fxBu4pM2FEfr0
NFvhaWDbeoKwOf+fvmoACfyU9//D9pV2k5PMVz7NSpYCZdHKesiP/3kt/z7a
kpXzWQTMQnH/RNnCvj8pLzAl2oJTH0LJxVcDXa+UV6d9S1MJM1ymBCYp4NcU
8vaA0/UwzZinXTmweCC7OyuUb7KW/N7VDW48pHez/aAPjY0OrVZOD7NRBXJj
6kwY5ZfBcgSHE7PvRKrU1WwSONs4aaoZ+Hc8gGvnx4uMnSlIyDB6MCSnq42i
d/FCRieQ11FT1TLTEnZG2bZYUBw+eEa1Wse1rclmjK6ZiEFRrA0kWlOAyGkz
Q/Cj+HDw8bt/+09qZTrAkuBZo9Q5vrOyunACmbWfAXAqEtec+h6XusEEjUPN
mftQvDxCy8nKe0G6wYLw0JPJ1g5T54Ial7yXREeBG3dJN64xZpFgXGy67ep9
xtJIvyfn9uyfBq0XEmyMM2XLs8WwTpZZTy1AJVd9DGDJcUpS8TGI3Zn7zvp9
yH4+67Z1gRTB9YD+Ayw3yQ/WnmxzZLuWlLAVTL5i0GmfguxUTHEk1WahPtG9
VgroORA0wWr6yI36kcnmo6M08ZB7KADcmLXx1s4Q20BatEGZnD8wxTl7UdD2
NkbBp31ySbPts1pnD3PdtT8ZDbHvtn8t0syp79S2Pu5T+4Nzsi0I5nMBhPom
GXWYkR5a/shGxup5+1UHxpRzEh4h/kucuIsF6tWzJxPklUDnbdlsGbOLNMlv
X7mbYaf6/8ax+v58GmpT/iWCqifU/9jxijbRgVYCUBAxBG1QflLYeYPzdtjF
hx42JCGSjHkgPijCOmmHuccdZeRMXkRacZJ+1VVRD7FCd7I/LHTyiUj+wt3e
Ti0qRVkTu0KHZvpp2GS0T7t94GtdtHT0GX1nWbec2rpFqDYa0UNqMNcFuBbZ
p75Uu8AaahBbUxkT7PvFL6plKw4KrG+6YtSzVDrmhcmmbNogcktb3dB/1WLz
IuadIgJLdOeJdZa42rOmI7wFUfhg0gYEvEoMn2xERO5sOC9KvtNkLkdN5aBo
gOwm6CC9K/cAXmi9vXnd9GLhYhAU7lEmhHy8m8v03gmyDkGi0hekmECanqXv
gCWdV1pj/aKMN3wWHqIU4Fsh0D8CezFF1XdTKJILKVgcy890StEhjKswrWR/
CvtMa3D0CIngaci2dC8oxbhpdYFnU3ui8hac4E4kqvDy37XTE2KeqU2iwlus
9aMhH+AXW58gFczt0zan2mRLdqfz+heSj6E+lqdRKZXtXINkneVyVDazTWgH
pIx1DjqCAOUTifgSxMR2XhD26IsoaJ3TQwb4y190M2iipcj0gSgYytcHAMdY
gJQ5g3es2yMeJyyWuIt7Wqp/4KiN6lZl8KQ49OM4Fham9O3QML1YKM/f0XBF
Lri78az5P9R7PJN6jcOjrI4Ex52xjpxdbKGtiev4c0VEjLupwBXE+PC+gPYU
3ktQjz36mIk9VfPReQArz/4jLWX9q/bueS0c7re2Ctqg8tW4dGr1IG7abNAI
SCeda4uEFIYdZSknx/kST8zDMyQAiJnejQVnT4liSeMOawZbMz6JZJEXlNdZ
nxtafk2KLUZRTOdLBrLCzfOKRwQexxgwi5DuvqWgzOjUiyoOTu9ysG8rHW2g
W5zL7iKqu4N+IxrhOiB1AVSJDizGJUcihhLmT3E6DTUGZMn3OQX890muQa/e
oJJiRxvOaiTtPsaedjkmEjM8TFpenl472lLSAEmblm/X5nN76SBMB62TXezi
gF5LX2ZQTmEvuHZ7a6168ffos2TAfzRnta1UXhFhyZfiToovultlAKUq0yCM
FKmpumfFGiU/vD95O0gDZ3/SyrWn89AaOOTnAJegNuXhjZDiiph95hDF+SmS
y+0NOar6wFz6FrzqfxRp9X+2qyBC9Rw0X4Rjg3/aZPN6AARFk0XcjKHYMNgE
RBUEPfPJOhwNATyfc1ksUjPaj3vTAogLLUf4B6EI31raMuQqFnmEDfCX0ep5
UPihHG+QKSh8Q84L7BmqwJr9p0i0MfUbb0pWaWFWxtK0z9zSD29BTm/gMKz9
ZgyoMSJ5y+lWx2wwt9H7gfqjTrm7/+kNpLPZ9sKzQCb4PUbn2UakNtYFqU2g
WQCGFmq4aGJXBfVZZUkay3TvjqqFpNJ2r7MR73xatBnFLnEx6Ixt7dGIMD14
SzA7pUtOmS0cwsfMgh5SOj5xHji906mvorbD9iyh7BA+EXUASesajjDPzNPn
xD2VjJH5KmI3CS7yOy1hjD8qthmLPp7//lY/EOD05B6D+U113YzF2v5YoN0J
Ttt4nvzulGkDur/WkFkPMwXeR7/oHPd3E6Urjby+imtKfYZaCsEDTwOKRHz0
CP80ga0+uGaBRUUN1qtPDS/tFWSELaSjwtaKoLvlqjT6Q7MHifCWPYStwwUF
xlEG77u8sdl0gyj/Kr2lgEz/VcfEIVXLlOMUWQds5ADzq3VntPR9bLX7JqSx
2MYbY1bIzwR+iZ1ffINVacg9CeAFvjsbDJ64Qjb16uF6WJpSsW66+NnBxYn2
uCJSLfe15dXfxC0GtJh3W1ZRf1f1bI4Iqbae5/ZYI5tpq/2SVW2XDg95jJSl
RW11d/J22Arv3MTUuU3VhIiuOK7k1Ix0jLvpMIkyknGaBEhiX25WMWmw0q4a
wL3SP6lelKcGJyy7kw4zOGd6CMlmR6da9vmM6k2Hg3YdUOnyI16bUN/uR+bs
ZFwSrAwu+0SXckRfdYQTlu6T0IXxfUEB1t9JK7Is9Z9cvhev7CAqU/HFW5As
BbWuwTzx1SNSkiaY2Zd7M+5vEBXg66j8eHYlMtCi3ccXQd98YnUO/qlVYPsg
5OX7nPK0lABYzTu7AEBt069IoG6nzYp20JnmfOukCPKO29wxcmF8nJUuDIaD
0gsfhXtgYUUqarGWpgDK6PhSrhVo1YnHEKFlGAV5HPMQKWtI2BHjUDzF7ctw
bxrNKzGFv2awwVnRRkEChrSwya30fPBrAFQOiQL8QK4sCtIwsrNK02g3yJ/H
yXpUcyY/ExbmPCPE4EpHXBDZyCJu5v6tZzcYkpWONztV/dFHrPy5kVCWOE+n
Rackk1fO7Mie3tcG5mu62EyehE5FSSPyKW6NpJbYs9x5aVCQ/PpeMTXcnEg1
FnuFpFZf8auTV0JvxH3UCLItjjc1uDQG797RjYYLhTW+16NBqgkNRyF5q6Il
0Qo+ZpoABE0ukBIAvPLrlFIEWuKd3aIcMUNgliIZ0OZVmf072dxVe8zQ/uxq
JNX0yHUXHBNP9dUVT5y9gBs2UXSHF7RCPnRRULlxlVdtkEs1BBrHw6FN4XYH
JA4qq9oyTNkcxb6T7uRcGvuicz0JoR+i+hut7Wc8k1cz57ymKUvg0ZV0oYr5
zrpAYr516VAx5ZikiocK0io/tnqipIc8iUAebl/bTrOsWE3elNecx/4Ogwn3
KF77iKeo1ZviBGuTEAwm9/Kw8BIZ0TPLTTTheNSyg5MLYfHvnXzDBSdiNC+V
nO9Y1gmmWi059GKpF5tT6F8CapKTRjEA7fZl1ZNvNrlWTgijcHPJmfnaXyBX
x+vadkFo5FH4P3Pz6MyIbSwXEhx4cC/XmiP83NT2DpC7qFUbbi5niuR9yqkp
oYl1rY+WLSR07pZFMHUIt5n5H6dwtQt12m4JhVrrnDJUBAFxWpRnfNbbdEUV
mKYfuQzvNKb2/RBgiVthqoaLae251LYXAxsiHT8XEqAC5lrKhMbkjAogQ3GK
Rcx0mBQwhbF50zCuw1A8DKJvQLK6aMS4aQfydwDBGRHfaORGax84FiXBTib9
RXgW7gn6sWELOsYlW9I0OkP+4l6doCS0tOR0Frsu02mCpneoMuZR0iTThR+p
gPfMH7SJWIGgt0DLur5plmR6ouVPB6nbfVttSE/E1iyFCSH/aKdOI0lyqVmV
jQ4uCJtEEBd1KlISBqQ4TBQ+S4whly0ozmHyp4CRd5M/c4eV7kaigysjonQ9
mPNQgej/8PtxIZ0V+ohbQKKAuDnqEOwSP3CEaaqrZQjoXLyFOtBcRlQt36Iz
5LsNxELU+J0Mxu10oVg/3h7mNghlJWwihYFwIuj+5WJ7hAJ2AgJbKxGWJQM7
ScHEnTqIHMqKctW42OGe48xhBhU912iTqKSTmsnTOkCtXeBRN896ChyJwU2o
j9e2auch+CkK46TNI7BGk91BEQu9hy9u1AGzpTf+KfupY9nwYPiXVFpPvFzV
eRA8WZxhH+q8HqNn5ciUB1YLFSw+e4MVlxGXSgshKRYbxEW3vB0yTqwAjtc5
kUTopkIxP/SRy6giCqLkxQaIg2dWe/bOj23Vlh90Q/KdYHrfg3S/MRmXbt6O
WG3oL4pzbcslRZy/0jngaLWNfZzJNBlxa6RaQfzXU2DA6RRt4huJYzTW8UxU
YBDO89U7vJa9thPGD97P8uL2nlwAHewVrA4W9Y6GKWfYpCv5rk7wXzQFoJk8
x8HmlMhL+YCpAQxMDXo9Ho6Aq/gt9vsTZpZ/hxTMVROvWoqOP5TEBBCf0Abf
ms0THQuv8Bsa9chx1qje7wSVhCsRsl6ZxmmkGszXxDSctazjfaebJjXubD7p
XQ4rN07jJXij9SOJGU2fjWAs0nm8O+qNfa7IoHyYYzlamBVl3Ii06jvRAVbk
QmUqvIsU0URUk+nhIPf2R3lvqfpA2wxZTzhw0tk+Jm2gpQh85mEFqWNutcnu
QddDSLO7Obo9ZChRB3RrYcVe36BQ/eAv0+TxGQCC15JZKRXtoIo2CbuK11iS
gX5SVhnKvsIvy68YY/EFWOhyKrH3DY8wmj3ufowGxhUkCtIlEhu/mnztVBZ9
qPFHFBqWpT0xRVE1AjedRAi/cLK+uCX1AdjOxiQZyaSrjiiPFZzO6U5V2hin
CxPzjTA3wmFadyrf15POWNjnXbK62FekVp2iHckaTX7+iemciZatBezTk4Uu
A9JRsJ8qBZsnrGY/oX9QdeJJcRhvYGrVnlwemcjWoHCQrBe3DB6WyzmV4biH
hap6mskXc27n8VtfjHwwCrYLlUx47n0lIEtreJ0quWiFimV+JwtcRey+EF1k
O6Is/oonVtG3e7/LzTEp6Ve58HlksOC9NLdR4otlLCVlAkNqrGmiSa9ZiQBX
JUHIOhhjftHQAN4BvhVm38tZduUMfTsMM78DMsL4A/azkkckW4QNnh1B8cub
dMUsfaHBGhQvrOw7ZtShxmABSN6w3hvXsBKRDzWXw6ZdMYira3BiiFbTtbwF
GI2LiaqOU1Dnr0rVmGLJT//i3hGkz47Xlf3tsPTDQeyImxef4t8faRNLuZl2
NTfbAEFyGshwPOd+UNk5hHX5qTdJ/mFTl9U+QowkzkSgsn9nGE1ku5BsgXhp
4lSjDENYu5qSQh3qhhz9mFWsYSPEYcWWgiU2rj/DfayJs04Dsy+779ooRXoZ
32o8dmYSaBYfSWzaG3Zj3dT6i32WmrTFTxTxjNrG9eKZfOlFUDLJbhShTRRe
oGB4TOgk/CaYdVbpTAwcG0zfrDra5uFVxUjAaxhdIHxkMXT7RtQhBk+xHIzw
CPhEAw1Q7TIJlAbotv5RTGiT5maAn6iNLE61S0Q/pZZCyyK3uEBwKanMNbt+
XEJ5aRYfH9vCZ8cUn9hVukR+n9NqxPRTXhBKQWFSGW33cVl6U/72w1bFl4Sd
iPhw0yD+JodXv5C1Il6a8zus0jAiVki6TMFAZkXpSwxTmcFZ1LioIUwu8kEF
JzYNaKItoIxt1L87Rg0mV4pCLAhXS5DV9NcLZmONa+tvs1yqBT27P96RjFcv
WdtCQ3IU0sThChp7cxl7Y+6fh9p/c9sFzzTd2krZtZYDhi8jPCL8EFMpcuNt
gjT6VB1uuytwSQV/diTc5DRgYxmKOdPlOH85BbswjCrpEM2snkON+cXmyWZQ
006n+SPZIbyV1iTuoDw/qhvE8LWCtZ7C39FzDI//3ObOvaEIVG4EhNyaaBmR
/IiLVjwdiK596XSmG3bbS4G6xzZ4pyEKyyjs0eJoQOHbTYPjKHqs6BSgdtl4
ZYvFtaL3swiJqIFDCv75+eohkwxA1iG5oVkefkPV6eKbindU0n5SYmqchUb7
7JHsReuQSrJRCBr0uNc46ig/XBprPxqYBDPpEed8x5sGdFITMjaUUBZk2S1R
X6tXLVByP6iQPRlbSYLnBR4UvE0lFOHEwKMX6AV0OPEo7ikAYW8KDjmsaRPZ
wVte9uigVLV3VrEIAh7xHFaX+/nm2PXzr4UwWEvPSnqFpdiO/Gme/JDgfCRP
JN1p4+1f6R5VrWoSv8crFfGz1FzvlTWJfB+w5RBaEj/PKJ64OMEWgrx2WcYp
/VqW+sOegcG/YxVAyrOA2N+58PCmlsE9MdFkJeK3+PrgXAValtQU7EqouqGV
iYS577hstQwLWHtq72XVi8TG+IwA7wXtKuMvC1mD6cApjCa0yQF7T7hRmcTD
pSmHZPz7gLRgN9paFwLvCq1jF2ddyF4tgKE/Nm7StPkfZBn4XiTZiEYU44oS
ysGeOx3yP5Ram+xFwf6yojVtgI75pPGjAbg0dFKAW9q0ostL+CE6Zv+dhddG
VruWQ4tqLtLaHyYEHV4hftyccJt+a+3FL1IiutuSRtJ3uRpR0iRBmLmc91NX
9Fg/vshpXb+/qMUOgV+FmW/nBTCWkTBe1quPNyN3yXwvUZzHTX7Q7+8LRPyo
QzWQWgqK/EqwxF8tzUMGEqztP6BFAqRlZpwchPEQCQd2/FzFyZ7nbBWMKLHy
XoPfe/ElkoKAhVDCTk3gKuXn/JUtihTHsaT8dzG3x5Bg9Ch3OZAQxvzrkO+m
EwqYkYIGnP0HSVm02McptmIzd6IDyZUt2BiyPVqSJwl3q4A1A3/09Wugfr+s
l7045UgCv/ylPCFYf+o4jvb5YPlvDleTSmm9qXPDjk29PHMUVOEfZ9xm262k
pPz8FFSdzFMYadMyOFnx47ug9Y9MNGJuD0AIgVGsgC7+UycTGTmvPqfhsL7q
t+bAZHYj3WPXvMZLxm8EJsN/F8z9pcFOdBWNmOFwiorjnjxHBaUXykk82F+t
9HxxG/22m/gqzddYbug0w7RXYoB4kWA03Do0sYsbW6QIEYAEM5ZmZ/uvJ79e
2PO2DkhCsJ6tswUXeV91oZEFcg2PPr/+1TNL/5heipLHlNnOwGlwHH/H2CZ+
5s0bz7ifShKMtZY5GM18nDK0cGrX5qlkyIY+fcGD2uBrkdq6uK8AI8Z0Dr6d
0vnyp7NZ9W82bsZi+uCyegaY0nJbjeX7XbyWY216rHq1UJI611SRMjjCnptN
iqU78www5spIfI2yjOowaT0H7GhsaiAC2iZilDl4jRO54KT/m9xzT8ENCgrt
6xs3Aiw5HErJ142cDU4LotFpeJe/ZtkGBla0TwY6Hy2lJmtZics8l8vPE8c5
q0DBe8rV+K4CDVDit7sJ/7i+r2NtGf27dFrPK3OqY6s3JMQJRpUn5rm+erv8
rfyxSK+Vb82k2uDrr1+ZLdsBxqPCIQRTyJcTJNRnKgi61rlfg7bIe4uaZ+bC
BoCMOk+sTbMcuw6cfe8+/dU5LHnkkwQVPBrlTpJK3u5u38ty5MWgbKGA4t9y
NWSPuvR5E5pP1hlcKKHdkVRB7kKekend7eznOgCulPARprqUv1UKbNd49cql
8QzwHJyBEmNedqYfpn1aYw6zYgjMcI4dXrSEirqNN0u3y52LopcWkhFTJHlB
WPlG4tkWaHcbNnsE3bk8wAlhJkTuxBW67KDPg8+MWyvJfXearXjloL/nboGy
29zlZonQ0KGYxfK2iZtZv0DSQtPp3+vbW86sfF+7gKv7+14I7kuUC/erJPWJ
tXOVUnlydOWofsLSs20vNNqmvu0pctgHa8W0bnCuC5MsblPtqUaR5JpkQfWc
z5bDulMUVxfVOszEXXMYkTPljjkpveXDBdCrffL3x/mWjeN82enwRUKG03Yb
DXbn1VFrGra2tnN3kUFdJt/Hqem9FNwfiaStk+rynewzZ6YZa/KyrT6HQIjg
UuCHN6e7+LspKdtkR3axkVNdBgIZC0Khl19cqsYCKl9EIv7DwBYlUIQMJunv
NfXtvrxI/4r2LqYQpoMaNFkx2MkhTfQfrDL//ZxQ1SHb0BnkZKXAgGiUmKuJ
GaGAhM02d9PYUk6UuUy8k/o04wP3s+eyMJluFPXEyNpVAHV9bib41JH2/W7e
7g3TkTpfWQ9QjHlmsVNVPnwjOX4FXdPWKLEzl9mjbEhQA6MsbKN92eSkZyYt
Uzya45JruniqKfKim6zvmKRnu52FwUdupyoXzjDtfUKZWQWClQT0xXeQTld0
4u+910bf75KqUFYTiuj2r/MaSClb4yGjoHzNdd6YyqgQDWamvcK67dvSHBRo
hQc74hjrSm1Ix4LL8ENJ0KoWRueeyXQHOFlu1PVHKHTZQWa4lc+/8NprzxYo
c8vnwcPs2iB0pixkZ9nXsrL1kE1HcelR3MJwa+akPeCmeJ5OmdmbTbp5UBru
8WwrYlB/1EjDu/4b6LJSmD4FMOE/bxTOPyXhX9cktk94tcSI7ZT0EO0L4M/M
pvMyLcj3PETanPgSgzIr0R8nMbR58BW7kI1Bx95xM1U5XE0vg0YlHV1FvU8I
gVORHJmJgzFukIsHgXx06u3roqYZdrTdlMiI0HwbhfJD5ut45ZAgcZAlu/z3
OmlhZNpar/FOwqaQk8bwgAnssEro+NAUiFyXJprx98+0OBTR1g/IM3/7zA6b
Zb8MZM3saZQEiTdKHRCoFDG+iyIgKtL846kAcDglAZHeKjIoVeWI/xG35QDi
mynGkKGDoBjeRbJjSR5UyU0c/ieKGNPwR6dMGQ2MKsLXMW9tEr+FVJg6swxj
zQ7cGe9/sWZfNr1bYeQxvElbjUUpFuVmYBzw9SpLr8ApujxbemRs/dTbRDKE
9rtMfdetzzitdos829W0vMyoUeStllFS8hV17axpK3In5x471vPRpjk8Dm2m
Opb4HCxl3kIsLJjqvX4aySxM12UVChjV00Qqtv4OWQQmh3XLjDqPTTrnEgWa
bWc1EzotOPmBqZF6tNfQfL/ExagKGqk4rlVYkYMezr9xuq+pWwtkCsfO2aSE
bBinQjL66jhj8J1yGOwCGdokgVXQ4M3GTE3x/A48qN97M62uSqOMMquUz7k7
nFVZjjc8i6JLIKHd3HYuD4Izekf1lNC729ZuXKoBG4ZwvAorPi9u40wvQxQ4
VTyxpg/IXY8uxZfFpPLay3uDNDKChl8jpo3t5M7Rj9cNZEYpqUNlu2csxsxn
WzljX3heS13Y1QaYIyWH5izGGQF2Z1nO0Hq5PM31AXbquqXTHPpfWC+HgJxR
o8+BNXBoT43I/kZdY8FRs1oF3vAhFGIuXWWFFZ6CEjWHrYce7nfymVy6oOs7
O5OV+TrQURGRy8PPD4fXuU3y9WTWB6TXBe/6sMGhXntAXpuDvPZth2ZgJ7Ww
u/fuj6JQGe+uyF1daxgq83Zdco/FWIqJ8ikURGUSL1M/0HA9eZ5kVT1QZCV7
O5F2/SdCT6GShMf4tRGbQ5X3uL2UF1N8y1x3SbbY6mL4MfxZAbGtefvKmnVo
lp7j1KUZi+7QY0Z1qZlgYAOrwSt2ZheBY7qIoxQTabGwZfDRI5Te/D/R6Pv5
d0sIYoJ+9r/YDBibwfYrevR1wnPE5APmZMJKs2hwOgzRt+WoWEYJgjrno3gc
/y5ejczGSm31kGWvCUYhi4wQN7phw70UfyZscsdw/RTsYh1kHSP3pS/86Ezd
ODA9ydJPsIdT2Rz4J8fkB3/YFtauifaouGOzMmEmUhoOaBG7TM7Y4Hz3eYle
RzCsy6w6/IMOtRUQ1lcLgzHhrzYNXwJ1PYxkh94kWby753Zx9Xj3e0Qsu7Py
hG6CV1XkpUqcJ99hLSXFjSN6IjprHP9edRnDmlMyiGZCZnXCUJN/y/kAxBbo
Fg6rq5+dOta4GCj5xyCX4W0qpZ6Ps03llt194dhgp7DNBDQLGjR8/Ynxy6e9
uDo+zAWYxhZ6Gz2zQHw1bwrf1AAjY7nhgyf47AKQ1oOR6FEHebhoxCc2LY7f
kMgdRFUEAhUnvQJAjq5hhRzOEATVK2jUQdculMyAH6QxKC716HtzJnXqBBw9
GYw+PMWpsoYYeC/UmpPowXHYVUl/63muLsBklBBC8002p2J7N1rMXqb3eNdB
ogqEUAEfn6rhoQ83QqDiMZJta35AKgJFPTPy2vl/ieni9e5s6vVKWnIxvyzZ
cj2Ft9afiYxpFds/a11NLuMl8e+1WTMyS/SQzygLRPtBx2urbypRqNpSYLcg
H7bk4Op7Vd67gBJweqiUwjFHRnZ4oem2jw+6raciwptG6j7YgeO63dZhR1fE
fwWOL2U/y2FQN9NFDVBm58QWPyX3kymOJ5Jim+RUJqLyyHPu8f4tJ+2nwWaB
7bA+hzMugZ2pkbz1dmDzQg7IFdM9lMHxCCgX3LuRPQLJWNj1HveP466XCr36
JB3/qiIw84iXscqJt0W4B5CqpsjubBv8YmCXATrDtAp6PmMczBPcjBeRNmAM
jezMiUFVamJOamjEdT7vidcGx7cGOOAQi4rD1U+eZrOBUqZExRvqTtnu8fEm
754l9930fThsueocIUxgulpJsvE24igsJIttSJ/2ati+N7nfXY1IKPJ0Bo7f
xYOkOIvk+6kRCNrbdES83gRvLO84nfJKnmK/CGw60f+SskUZXY2eG5VHKEZc
CY5Zzixrlp5fQ7YMkXbENSCHi+7MtMe1pAm9jle2Pohi1opxy5/5kIZa7qR4
tlE6gzwB7C1QzTu7ZFhipsY7L6YVg+MijUpinvReu3tkQDv8nwiGRzgl6I/7
PxGONIKGNcGyWAkRE6woJOnHYtQSZfPLKS32/XM8tqE1HWa4BLM12PxG7Oyx
i9Ub38cpFXU1dH+ir+dKg+kzm2AjmWgqwd9d7Fk+hjPIfNJDAMh2LFu+rMSl
1NJBfICOiDqkOFP5SMiTiiiQXKHNlDPrTpS5TFNdCHlG6qkAu4PiL3Wkvel/
K4z5bIKOT3apdbsJjuhY/DVKaUsVtZ4T106NMQ55WImrlD9yva790D4yEcga
Q1VRT3f87bc4M/mXIQOhT1JOKDg9IQyhHdD+FkHV+yL4ZvedxVT38sv98vK1
hAQbd8dmyD0JTaQ0qzAaoIdQw73/boPhaF2cegzHyeaXn9Dd4qJz+EkdSqk/
5ll4QEHAPBGfckpnw3X2qhWEvFMV0JICvuiCct1BYSaG6Q6ARKSGhQlbK+Vw
QVmKzVvfunVJOX6gcnAsL56TM9/JX+tKLzx8G51T7RjS8jwo2SIOP1JMUiNt
9wdCUpTJpkyM6igQUqF+2vZiNmO0KMuMi6BYiiW93JFUAB0Ub9+7CWMyz2Xs
WAnAgVL1T2rK59+THrzJ1t7pZr7bP9u4KoaC7J6/aaaBMn8EOgV2EwLzUBz8
EgGTh+NwrF69kac1f87hdz8s0EtlC4G28gLTCmsnJCm8fgCf9k3sVOeSSq+4
zcZIPxkhcT9D+conHbLOonNJteJN8XvriLoaOgGhutr0DTnFEFILJ3s/zH10
/+7gDtvenmINAYJTh8XRCEDJXrCFkgHxYBlacTdUihLPwgdAiDg7PlY7vxsl
w2uZJ3vZnczA6rFRlKGJUaV5ARCCpoOxf5PzEIPN4hyTeMJJBL2gK1ANSqp0
IcRutOwAtsFs9xSlifxPtV9Vz5AtOR0++C1ZBGl3jSN20V5+anv5VGZa+0Hh
bmmio5fXpLAztmiMuLLal2zvzpMqULh5ss9HDyVUy5OTl7IPnNZvl/pzsIyw
XAgGYVoGIDnsnTp5afV+43Q5UFv4Sv0YVfg5jxTF2jtkifLhIJkMSWUdnNNE
zgyN5OVKvkgHdDKFlcTbvPxILIU7aBO2QAMvKieiuE/gCE5u40A7+Hlh8bcy
aMDm2bvXxXy/V8q/KS7U5fyEDJSU0VBAiaSJ/agnaBQBZaa4D9QyV3xhJ4dF
KS+Kqm/ImfleLs0R4ntu8F0sQkwUpWNl0sPRDCpy6SpMaCUr0elmZnf1bI+G
CuO6RV99U8ZYe0oS66p9BiRDSUGMSFMEIXL+B+LsjzI1YzvB/k5AZ/2ELKnt
n09AAwKgU0mwaXZhOGS6yaZdssjx2BxUC5Pb2+ww/XlNGj5c77Endz24wt4I
QvdN8NQrjNutyRwH9+BniG5gmQG12777MWT2wl6RckmxmtPwh/TjQz/zjDJB
0AFQh3MdQBvO+ra2/28bwoAqpmNEVl3IADI49/AsUc3FobnUVqNiR94dscrR
quxEpYT1i59Rmggv8dvBbvSqvzxwbS9aM5e9wUhzfUABICMnU14BpaSk4ESV
MCdgw8skvfSwWCwLue8A64o9Di1MP0Kp/7JYc/Am2hiYfxFqLsBcBiWHv28u
mkVjkr/ZIF16c42HDew8w0L+E+WRevaxR9Gk1OrNlVPWIaI1ZHlAtcV6xN0Y
3d4+qMzXpofLYWNLdGkeyKBtl2P2J+mi+YKTG5xfwHIU0Le959BpO2w6OTAP
ys7MlZ9TNJEuSAuVr3kecTSqBOpWXTIsV8dbc6N355ArQZEu0RW9ECv8xQgh
MVcZH6uKy32H/9p2NyluZLwVoEVWiH7i/6rCGS53ErX0SyQTvVe57TcWX+xj
f2Mg3m3X8EDx+TVBtq6AyhVoEYfS5xjCqoFxq57RTZU2K6BcB4K2bMKj3Ozi
kz/KffwqnMfKhNjh7gh74zMIldSuFq+VSUuicbrUVg45UsENdPD1rhTARGOU
/L2XFdA7beUXVbbvn17LC+yXfnsddc//RIO63RQ9p4lWCMzB1Ba4EbSMB7J9
gE+xMyJzgik5daQMEq1VRWRzr0w3FjZfrPjxUmeoBxpiYUPIQTzT2cR9vYgK
n7KpLhlU47YmvcN86FkyfMNSjggyv0jsOPJqhLbVMU4UzZCS1Ox9Hq38Sfqw
QAQwf0zW8hGPpyn+YWPXKrGJynHkyywTf4bd9PqeZzuZPTcpJDDEEqXAZvQ9
U71WkMbc/G5EJ4+bD6VITEQfgKh/sFbImQ9AjGxG+9rtQK97ouMEn5zIiuqC
TpW+sLfoOkulUuBQabazCPmNi1lR4fR3xmZUGE5TNJ0rdSsd1kLC02FcLmGE
Z/xUxltsYnI6uu+4lV+ezCaAxzbnsCj+KD7d9tPBMJF3zDhG3Kxz4nyjoRd7
uX1uvigTk7NLWU7yn/3m9+zEA4mzlLQtWp3tjV8G63Cgq3Cp2vYMkI7sxw7a
9o72cePmAjB+jPHuMW7dePVDQbLZFHbpnELD+Cw0IdhL5gmhh1V8B18Ggx3E
H2WMcWHPFYlpZQ1/MzoxRnSI/qyb5OelnItNZQK5rVeku12aD95TlI+UgtxP
6j1dRN0ZWr0k1B6ayROrZZVQF3GkN15khhiUV3GKVjb6xNv4+360fPjHEJWz
il+NejV9YeBxC1KQTffsP/TEhuQGqB5lyprgiNkMrhIh8TP7g6iyHEaVtZU0
IZ4x+HXvNia7WhtEida6K7zxY6seZ5MDs+L7gQmqI/t0bcSJoBmWoNoS6a9s
LOHPTA49ltRihhn0pqtT0JAcc5SME3yXUwAw013WUNG/0YQqrNHYKbFKNp8J
KUDrNHU4xqXbWH6i7bH6dPk4/4/dckYEItNO7TsQ/zv/UVg+84UhIfBubuNM
J3EkDg03gGHs1ptWxPMarfwWRWMAh+g+VF68Ii0l7IZi1PkCOt4YMo+B9+HG
Oci5mvW/lB/nepD4MHUKC+13f9Szrgs/0XsMlF0EkKnjz2VDH4phUZXMWZdy
CWxsdeTcQxFqg1z4UZkEOvXjqLqdTz2vDWGddtDBt/iAUUyvSZNYOqVYzAsh
mC80B62lYxxasMGhgCzNQ5wznpndJczoJ4I1iAsmJIAyTTwZ4CovNSFkOXvA
sNIJGzWK5UBaWLfldX0xY18Jym1GUM00SA7BRiOGjtcasu6CZM/CYkXvpi3M
ZT7n7Li3fJCe6EYkqfhfdnJXOUD4kDPI+z+KdMYiOxne7y0nYtWbZdfqqgjp
i8lfx22HAWDzh1uKI/Ez3Bibl02PrlYd8GC1vOU3CdngCOKp2iIWU0MWpQUb
A3/Jtbytuh7gZLAAQK1nmp4OXw7Usbe38r0B5cfiE8HiptSkKO2t8HTqv8g8
5c6MEaJj8GanpSGrFdiESrEVrGb6OUSUBv6yJNOES2AM5qutd2YovwdKteCt
Uogb3l7hMyhszRoNExnFZYEWGY2iifCapBqGknwbufXt0XIxXVjUqTQE0893
Bd6jBQMOL5FGmCLcVqgJLik2/ufnyfqPFglCCzQI6rY3g+KM7kMvXHHZhDV2
vr9EmF3x2s9GtKH4LCeOJKPWHu2DrdbkKqPjWALFXjZ7chJ7FWPiD2N0Krn3
Z04yQufqbT9q1JPXNUG89zSnfq/CuZ3cuZacKtb5IEv40Cy8DVDmDor86Jy6
89G8jY2AOApLZRfYtkaAhcm6xKBaiFXjHWFzTkck/8n2s+7dYMKO5vZPS6Ex
CJ1E0Us60hXiU7zuwOTS9whT2opcyypHd87f6sbPx7/JTcyTKXMeyVq6rgGD
GoBTIXuFj1WTYAs4ZPqNdzXDB8hzR/AgyufjeUzeQQjnyk5xAq/DKWE99FNW
aXT/tNp1G7CrXEqIicRGuoXRoX5DLoK9dB/e3CICm9Nm8IB4BJLKy1+w4WI/
NCx7I5ENAmWVONsY9ZVv48UWdo82NW2xx1QPK16OuijMbvihTb+pyaQ0tu5S
l1xbe4Xuyyw8cSdjq5zxZgGMn/WR2aKiqwouK3D8qYlgQX67h9halOb31x+A
2YD+/DU7YsPcQ+ll/J/yEaER18SHDM2J3in6d1eIfilT1JigcQICYXp6+wL9
u/qSd+JrTIwJFoTz5hmFIeozgbJWQgEBpKAG7lxTjffFOqEbsUE9jQKIz+z+
2v8GGlSNlr2TUtL4nOxw3PWd5YLdVv259EvQcyEF8aV9IGpVFAYgbYrMYv5d
rD7a9xlm7COObk63nkYFdQI4dx6scxBP4ZUWkIXgeQLS6BEuLhmY7eC40v8c
1DuG9T4o0svsCcJZI9/KxFD/CLBYAjTpesyQ4Y/52XGd2mV9XmhdnJIlUzvt
zr2TaA3rOkUTLi8lCYEb++fw1N86/QyaQx906/a+ZhI+HBVATG9T5OGZnaZU
/6XD6guxG6CGhGxcGMO4a4B0xL1NpnvfnqSPt85uDoPJgcLlEwtSyk+1hLV8
CK5FNVHNa5SCbv21xOsKgarzMf8BECnj02F12A02iwav9s8XNCLJ5CAJVZvi
ICQjseZVnOsSaPeTNPObsQf3wcenU2PQABAhKPOBaaK3ZxFxlhJGrmRFEDbD
i6fNPARsji/onHVrHwsoAkkEWQebbPr5anz8ehU8Dly2qVl8e+dzP1UrfwxG
FTF8LlyIEgEgg2HwcnD2RafpSrE/QOZMYQSxLcdKqsvQfDdK82EF41xdhU1Z
FSCiD5T2gso2xShWUNdd3tnkP7FEeSKPxtuP7ocoSi05L3tpetd0+V6s811c
LvaWFV6AjLvHI5dXRhwgz2GGqZm5Jm4DiGDrdVHdPMursg9VHB2Ma9J1RE1L
hc5BMyE2nsZyi8D6J1d8VeMQOGMvYUqmFIFC2S32iOOX3LiDch9YI1QTIjBQ
mlOqDBxi1rqta3gz4ajxJ5vRVZ0RwnOhurKQR5qPu2umSu2g9azKscSVqMkm
st0EyuIwETkLzfXst9xO5xqt0WnljmyQU44M7vDE8sii9cghhp+r4/g0tTy+
N4rSDO8psWaqkA4oRpEsGjTOa5w7KQi20lPlfcDiD6tE0KM7k1XSYAo5QT7m
JojV/ChXWL7gg9K0npi7UIwb1u0onj3CoeaVifoRN24nMeX1ofsN1GsKm1HR
HY4QUUXLHiOAfvCRYDNy3XWhqMoWIvD9Z+ULV7Xd9eA3AAOqjZy0M1vZRstU
9EUp4rqJpCQwxghsxsH1euTVXVcnlkNj1ERCEJbwq26WJAYalxTR92jbyxUh
fS0N0aW1VZamh66RrDnt9PJ5wso/fd3hdBJ6aRRJOp7MXjgABsWlJDshGSse
m35MatcEwS0mRI+lGZrSYmwnvoof+m6hkvth9AXz/sGXFN31v02bL0VGgNpE
3nh0OXG5GMB+1uaHhevaIaUFblcDr6qf4AUHLbdArHyDE65owm1H9lqhzQ9o
gctmxkPLM1sGOqbeZu6yMvM1xQW+Gxk3wovkkXOaF2xd+4EvN1kQjdUqnLvZ
agwxdwvHGzkxOCNcR8sufw1a5v12UgBaM6U5ugsQCz65kQwDN/fayMLzR5yh
dSCPeT0JLbQyBHnrQVKvsGiuOoHm5CiLxMCV9pEckyEuvszGxHH5cp5Sz4QF
bciULB3r/62fGmdYO0vpGs2qF4MsPccVRuE0QmLSzdKUp1Y7CLooxLMXbNyL
LqqtESlFuPcCnRIwYSEJ4AnYvP8xrsWyjnpE7+PbsG8ib8kvPX58lb3cnGDV
qdu3tXJlwIYvjLqVgrZP6HRYemNtPoGT3dD39RARMU66LZfNPdiYddcMSuSo
eyrnfy+A5E9hcBonPu3EIjjRid6FLYvIfFnumaXAVWezBikUHc8kg85eb/1U
TYYx1Pbvnml7mHbOSOawqcJ4oUCqE24f6VJc2ckDJmtjXoTHJ3rzaKzy/rKz
CxuZe9AM0ujIhNK/x8YkrPDSGnJCjR1jX0x+4sCuKPqJMOxuYNW6o+DYl0w7
fVDVUzdVQ06hfvzJ0eDzs5h/wR08qHM2Yb6gClluLXXUNg2IQR65EbWCOKSI
Y4GSjnbWUO3mULl/f/nCWIWjm2Q7z8XATJCPrH5rF6H4+2NQAoxnjM8t9Sfl
G7eb4WAsOg/5MHEtsUQZsuGQ925rB28qAg7ybVFEjIBj1WhAEWBOXnXBooBC
rUTDIednTVbzu7WLwMxdjfZtms+e75Xhvpt6KNsM5FFGGGOBrRbEXSJ5UkCr
U9uLd8rIE0yTb8beg0HNAXwzdEyNUcINw1nQhBi/MMGkUwv4a00ozysx//5v
DZOg8UyGGGj4JqhxlSQ4VMj9JnGiRGy24a9U65Tu9XWrKanspRgUxC9/k/+7
1aC3bR2gMeNQHS0aV1I3/l59H8lJ6hmaSn+0EfsZmH3I57zc+m5UTNuZUBlq
4knpW0lRfHh+mJIDWCkseazBL4sd0FpJJ58fGOk1Lua2gcFycSEOtIGQxIIZ
G3AYwaDXnODaOk/zCChTq3xrUadn8Sq2vPuJCtcF7RO0roi8E5796ZtGvMq2
k0R/SQkFhlQeCMht2tq3VUSsnxDu9QnGJd8RCZ9tj0yX8lOyrDc3FtuEEML4
9oqWSUUVSvehNcZ+JlFBSh91DFn5b42jB9erWE4bwyqPRjn7d70fvLLSHOcT
fBDK/6FFZSajF4l9q8WbJitFPrnaTyt/HIIkcE9/+ha2LL4y00RZk4PDMk4g
MICEVDdkwbzY5oAQBPHrcNPHqWtKgcMvyTzrOHJEtWRh+uGYkAkjqUwi89J2
wz9o4j2GUcHoqGMEiK39+M7R2l2n92AdXrJjA6TJHU8chYsm72V2l6RqLXXV
ptPmPxHvpqJzLS9Lkcgwkg42v++fLStTmbEAA0zpnmu4zYLZQj82VcwKOTLS
HQCgdUPqJsOUM1W8yAEleHmmzZ6yy0j59fW1DIix2AegysZvRFxfbhBzCk48
X1UVYZ3TmkPJRYYYoVoj9YQ879xlMMzcgo4sv5o6ogsowdzjckjydhDOFuSl
ptRClX/Ebwz/0OFoD6co7jRy8h+/IctEjqOFETNA6w6xcKQh7heA44oY1zQ9
L6vIh53swAclr9Mzr9eQIP3wrkv+RGxr3HyoeJFgpy3ZX/WRQYfZRfCJGRKE
Js5up5fsFvtxr1lrCp9HTmnm36W3TsjOWUB4Hun34lJQnC1hAKj3QlbEn6iw
X4hegVrsAjrceM5SXDPAKh464T2gwMe8kIo9wazWZLo5S0hMDw+uieFiC8wd
GGg/WZ/2rqt+YpXeemGKG+tbFRXXHn8EX6xtpYF+6ztJiQcP7rdnXtzHQIAC
eQ15jbW79SfCXoJURYOVNJL5GLnpbMF0qHc5tok3sC+LjDEsH16k2d0qOfQZ
vLFy9FHk8TjsBLVqJjnKhh1FHJWcxSgL719sWMDlJCPHuZJTURS9zXAk5X53
YORq6t0YTtDOaOrFQVWyJkXlAP/mUKVg5lYu53ysEhw0iwffFl+xOMCQtvsa
ZisDfJQbmT5ifncjucB84GeYjfJvK9fLkN5y2mYpgw8qBN8xCnrdbuVy2/Pv
bM5cQrWa6TOr5gEqop7zeHus1AWwYiYA21993rYwLf0IWGXTzML++AQN3TMg
O32sfVv5mheibgdF21yXXBfvWaoJUnIGPwBMMynLxpWn2nAxZ/LLQUy62OTF
KotbG5/GDtNgjlDkOTIuRRxLkydBsmo50mMaB6STLPdv4vAbGw7Jx77poH+o
rhIMeJ3Y14TV7uZFenC0Ike2X7gAwpkq0ARZFWHlcCSynNHVDedh3Smp1Dm1
3oz4rbx9Xnj307eXDIBpYuE+U6iEx72vxE9SjHl67pFFlhMbZMAe60fHzePZ
ZTlnYXEMVSBFQARVFmraV1ayvt8/3Qly6w7bmOqEMuxESlNYqvCiLVnjUABB
MSQWd6rbz8MNpUdOSHO9q/HUiIrwx/jmM9pwStBadBmYPF4eumNWI3Y9UpGq
Hrd5C178qmP0j6c+cFhMo5b4989nOax/P/kAkE6peoovRTvuPiQt2cdPzHqs
trR7iyUJQ1d+1r3xH6qaYCaLCOW+4OKVVgH+kTdBkpsNeaAkWMo/TQAWcBx6
+w1cce6dw3WlWo4EkkCBygo5op7ubrYPuioKKHt+QPVY7XztB+DpvzUwqMa9
F15+pk0JFI9YLiA79ESDmwU7GC8ZARme8PTnO2g7rr+qRZJLJZ8qRYOdCiJQ
ECrDLWPgE0gKwUE8/j+qNJQB2JH4ilBEP3XuNmpGDZ3u13OkOWEWIKDiFYiA
FINRA+eJ11ND6UC95NdQpAzh2pUanL2i6uW1qQ0ufh6cbnXRJ9g3szmjXH3N
1i2Tb/4anm3Ze4yi2SNCG+SleZubWMzjgGCP1YZrgORckdsCxZSY1RHCuHH5
6gbbhaYVcPsj0DFZwzeV/NJV3R6XkL5q4iPgpmRWjbNe+t5i+V8nsci3u+QQ
6rR+LQrI7GDwSGg5/yI7FhdCMmsDSYqOebWRrZFhoPWlJMmCtxVsuSFalNEd
IpJ7fqdV2ryiDrIPzGl7UJl59GAT9FzPodLFgGAXC474QUbJI01NQvcHHjty
wIwZrMBSiV3uLrSXqbNsBux+H1d3cxCn8JAVQAEe/wy+xDsOLczsK6Wm0KZ1
MHCec3sAkJpKzvRkZm+oV+L3IDppjkfar/ZwT1gW6xcbaHO5a2lkKf65UotL
xYYVEIdvseDCpLsuC/ILnrd7yRD4Aj1ID8drJI72VvEhmlVXBXQerGlOQ9IJ
SB2jcNahGYiJIXTn3G5xFC0UUSRkzZMdlf2r2gzx2zcVaLc7WYPT3u1FVj6z
FP/ehFvM68vR7/hh4g73+8D9QuhnXY9CuSekhIF6hlf0mSsqurTxNrvuGF1d
2Eu+EklMD40pNJyhFZ3Ra6d2ha1YjC8eAnTzPaY8j2gpOmSwjVjUBT+WxU5j
blM9J2ivQQrmgcaCBQ9TMQPwz9n44WgfhXNFf8xnI4vhXB4WVceebP/8yoyV
G8dpTYSkkeucwPRSFywCzNUkuJgzvbCVqQ4rOA0XTn9FyCGmGfWMPzNRQ8km
PHp7tMLR5kdxdTxmkbMC+yC5DRfJgoYb2+O6hY5MzdOUeXKsdlqBXI7yV4AU
HMu7Q747/g/deJrkLomfVA89IIIdx/nrwIrTOfikm38PSYfTzqeBWk7pOPJc
Np1WdnjM9OHiIVQvVyh9UcRYwAmm0v6pAUnMEeoXlvjcjah4stsJusdM0TYh
DcalhvBcekszWVw0bNlpdrKK+R4nB8gusVNczuHeA6T3XMX/GXLEVLq8cuxs
cRJoqdeWMTvGlzgHhw01ShrrtV3Zy4KY0BiGeRtBADjaObSA/pjBBC82EtOT
s0AHfFywIcp7AB4CxJDC+jHZQPeRrnovP4oeNgjKKkHltVi5BOjWUJRWgNcp
otH0PFoX4szERaYvK2+5XeeMCOrSQyhx1j1At80VFxIWZ4/K1f19OMkzcSUJ
K5uXBewYFPZ3t5SOmpy+mxm67z6880sXCNPC2o0G8wDia/XMHRt2eM2iYzmH
uGQEHRvSXFzdRVVphe5zDXSZW235LHL3aL9O6szr0UaSd7zWerm86+H0J41x
7N0G3dpqLY7P3+uWhlaDKMv1WU5sjxFoXFK7FcaGiRCH+DQUfB+W2WUPrIkx
TJf3OZ27QRHPWAlJH5/+gMhzk7EvSdi5huzJy7A+memJwqHMnt72A9NZfU/y
mTqJuGg0XnkxvN1A3QrWcN1dlpyKPLV+SkDVJTgptDrQvD5ZffCr7du8Kkvk
JbYvjs/O6NQGjZWjbekrb2git9414Ur1olJSZpmpWiPtNgFEVrbG137XP38P
ogtUkbv/1rAvJ/4pFslBhVA/8Sh0RNEQzo1ZNoCGqh2w5vibNyWf+6e4/pbo
nHmQEVYzssPPRirKbWQehQZwAFpmTLGLRnU7sENlabnZ16w0Nbz433aEU6Je
4kjRXF/aUdw9pIDgEzYbvbXVFDmqCAXvLPUTcbRQLACOeCEyMoZAMvyOxmdb
RV0SDCOIdSdUZykvfvy1Ks9dj/G4qVhnZ3ARnTYA6QTfIHrXBZCYBTKtXaM9
Y/gyuyJqQbveSrNpvsIATP+kccaubWF2pgcNUHSGCneHkIb9sMr+gzrrjB2U
A+jBeBWdSmvboO1MFQCvcMxKmB0A2zujaq7Au8pF6aOaD8KUGs6d2pEjGg7/
I1waeUD0uif+cXzUwrjWHsWY4NLhG2OPZoVNR6Ng8PG9dVOvvnsVxTItdxqr
M6WtPGE+igc4a59/ymUY4cEk1saiLx2upEWYSObmE15AiJjopeHaMUp6CZEo
2sP5qzLLrqbrKOZDjaOKNfkq/n6ktUdtWFpd+GItKmPcc1um86l3ZWjqTDvt
YDU2Cz51D9WHtajiOS5O+iX34qU8to0W0Tg7OGF3isPkOKCOpIzdWoN0Ec5y
uMJdJfJB+agM4svF01yTlyXbzeEXIavWJ91m684prvfufchtXs2PHTgjlCDB
1wFagUQAwTcfNMUiaqZaa2InQFWPQfu0H6hfmTpM/REqomwppmGj/eTT6evW
Bd+n38y9WFKmPWCI7aqQbazraS1XwtzSW60bQI9dLEV8oFVgHH7K1iF3mccp
DlzxPYQEncidhYr2soRy2AgSKFoJL19nq7qIGfiyPOSFbWXAIZ80ZETaLl9x
6lqrhSVh9ZiDkfenQF7H1g1cox2sKMxT9OLo4t+xKxAPpVyetFNyvF8QgOD/
h8jpFZCus6uzynNzHY2ouYwSXhAjL531Hh6HqrjmNPDmcwdrV0SqbnRgrioQ
2NtwPteDxDiRkYV5oAMU00B2ggOsjDT3wYB+Knmuj/v7/zhbXOvzzuyJbmZV
A/ZCzc7KlpGbjs4dJ6NGDjFfeastleJ928uzPWl1J+5t+TDxtQM8d+mopMkN
3ONdyMebNsqBAP+wjcgYdzPFesKsTq9I93jXDKng8bK4YXtY2ADwuwZiRkAA
kJfEfuYwMJjN7iNma/x23QkfxU2BMsgBvYwV+JdCOacIwKHSoX2/noQq7s57
l2TmHs5EwuuwWKARTmKn2Ty061DlGSu5tPtU5VXtlkLi68i3IvZH5fEl8lzR
Azb+3np9dQHEH0DaerxkzpKdcIXoQmL61qL50t3sjzydEQjpgIf4H7BMGDAX
08zl28A68RyoJF6Kwq/jKYMLG6zldXE+NgbltTdRthwa/naHm5ZFaq4qYsao
XmUiychXhx8D16dt0cdl2G4P2cu69XSokWPMcGVaJzIODkmJ3WgKQn4oH+nb
GYtpjlAnsnNgbEMSBFDZwr6tNgTEok8OCLENdlrnZhdFY2/JOpG7UrZWqF5+
FiEK2NZ0dhlrQnvHwh2J5lI+6HRAmZSN+Kn8w9kfj3KjLy8cSgwN0OACzhsZ
AM5TBdyCn41GjigXVN6Hnf4WBHUBKeg6IoiTXsHNyFe6MPfr73ttdln6DOOb
yvFAj6GFgJZPW+rBSaMaZkT4NaPpWTVStIpz9ZhKSH80ssLK2eMEdrzRc6H8
bQbo8dlkdxE3dRIvhQ53otN7PkJZ5xO65ayz8byxWmwM1caccWCvM2m3aPYW
GS27qsQJD+kJWzA2rsz1laQZJH//sOkSjYx/1x9+AlBF+zKf/FikGUXIgKxe
HVce0YOLXzvdmLBrxMRev1JKSyvs2zOQ2Cjt1t65/d2bY5S0Eh26o+8I3ZGA
L9WnKSOdvQNKrZXYv1friHktvYMaZfQdIHnM7igi5bpn5aWd9xWsBor+KT0I
zN7QpY/gE76GRVlq465fDm1ZpeP+jng2yI/8JFJGK2Fv8Ee88rX/UgHtZYer
wkAhlYFHM2jSrkj+IxLLyZGX9ne0/9vrYBQ7jXHDGKHWG22QV4+E/hM0lokG
PPVKcbIbExcJMjkfb/kqGDLTkd1MDmcdmHgNgsPsQnct+CXYdpNrjqveLMXd
kXKLWAxwmsnUX1jB242gHgH5/SiJgaRQwG065wVS6GXVOrRBjXRKcEl1Ao9p
WjteA1oJHo9cU9OU2B2yWdDmqa/VSjk7NiY6kxQ3DbEMVwreryeeUK93JUqL
sv4IanLz5XwsHeUvKPx9S5quGJGttVOqx0XFoM/4VQkQH1zOUUGrlKrH4MB0
U0i0emK8sTVkz9l+CWbq5w3L39z9s3srWMn2LZUv9/AKTkY8cufSb6N37Kg3
8eHsRFuKgdACwtJ8Ylv2tSCjXiHYKq3A+zKKSwkBoDxDaWqqZvfIRaTfJhAf
rfw8VvIkJM6dRyQMRS1zb0hKE8ugibVhh3L0kRAghO/s25WUZm7H7YMlD/ij
sU6/ac+mg3S0ZaGqQ8E57YB9vc8/Wqia6vYgmoiTgXuyRxrXO9jsrXfNsn90
t2vpSEZXZUzdsouzZjTebgC7eiGwXKi44wR4+4Jy+P5LpLR4SxyWPqDaUoIH
3YyH+LfeJXl1MlGoRkQmDSNf2oz8DmbGlnnr8TxnwrFB9qSP5onKhdKK+vDj
AXsbNNGHI3iNtZt2dz6DyYbA97JChF69v/uCV01ThFQZru38PDkgbTnI7o+5
iH96lk63nNopioXQ0p2eiMW95+k1U8iVS05WaDk5VRwoL8IlnyKQzHCXuYEA
j83lFrKs1fZcbvQHDB8NsP1CJOGg2jxE7tB2SB0IsvbMplPq5YMVnGS1XoKd
/saZ7HjPjWaPyAt0WOEwI0OXgjf/jmARWFUd36eiQHCNS1chQxdiEJr6EZJU
xYwOfxHgGmAInYaOFQE3PhSKTtxiofmaeFEnTD3+WgWnO17023sZtOrsJTvJ
3e5V26LFybfSy1ku8QvfPHfsWM4soJJeM7IMqhbYwClHZaoficOzpo16Gy//
5Kh/v7YfNqMiQ9NektlPpjeBiCS31bnCQu3sQY94qtkgixpg+lq9oC25wg8+
g/lCwEga+fbcnYKfKyqXwTUNOJ+uFizmBG5TxIfyfocWzAXKqBx1EIhYAiXj
RwMrpFkTy9JCjPlukPrt2y44ohLztRuasO5/0RD7OhEHMmJnp+lRq5YZw5w5
6uYOEkw7DYXl7H02HCw2YubdXNieGy5iBWmN1TufOjwcuVPfvvCyr6Pqcspw
f+Euc3j2hH7u65vBQRjlSK0nZAY40+spz3kLVTJFXQuGP06jMn8JvRDanEt0
yKqCeYNZjeP49qb0qep7Uyx58pg8LH0BNVztsbIc8r8Z1quJ31CqykNjmp8i
4rqUeCanYasZvL6HKtn9Vec8MLQU4IrqxZ5vIiK4d/b+W/bHpRTMHAIhUtq0
xMlw4+CNPWZDTxZY2RleEV+7McqERyjVPo86ZR57n5v1Ja8kQ+VOAqKuMRFB
3RcpmbeWFEqqE5I08i9w14PwjRUie7OUfBUwgI+yyoZABH1bTjOPuOMH+up3
nC70MWdZcnSdAfS5lqrbiVCCOfgfob7y4bvI7hPe5bLNiio3sQUtX1HsRlvc
IiraBR6yvKoVsy/PR8oYyl24O4PgwjiDTjvPat81vfypHueyiBlV7E2XCSeY
JrCNyJsr74kwuSvWwCAFWjfSVfrFxjyi8L+IXLQeGjRg263hOwDifkXP1Ua5
B5rH2VBpArYOGkfLwIsIpOAs3n17hkmK4VlcxjQ29Uh7qIbWybtft4smusFR
jRjcxkzQ7TEX7NEDz13EaTtrLKiwUX0VoRHbP8+BAVij7J3lq1MzgL4bC/cy
k4FBFUzC5DnyhK91AQMArT7dsyMRXVDL664S8ZF5H0SyAzYFW50HW3RFpAdX
TLsaz2erHM5wSo1BaxBbzVjVuVxmClA4T9VeFoSXfXtQ3syEGF4NzxrYMQLH
X/p4Ez9aQ+B5aJAqHAVxERc/20AlK/PrQnfFwSpUKUaVoiTeP2SVuTPAa1w9
OjM8IKxTwbEFRQCmC57c+V/Ky/Dz4tGwRiDcukXTw88xK359/CUll/KeSyUN
9m+Qr9/avAXmWWKDXsNCXvmqFN+gt9BcS9l2L5/ZgROXv0tC4VgC0w0IE99K
SQ1sRud/mk3j4bKaB96zt2xMGu2CoVLmpsWsLS1/Pwk8V3N6JN4OX1nb3tIJ
BWiAenivWrZPCpiyNw4+Lukqjod5ZbqxHH4fzwwqIl4fD21P6W066khIcyjp
bF58vIdDDapOYIjT4ZovhXtAM14FKBosOYr6rQZuCMFoZjtKoKZGHb2PGwwU
zmAMzwBM4RgPkFmJ8qokWlvDOPv/9WbZyqrspNabw0tnvRvkk013fcFTztnH
DsByIcKDyXDzvB7iU8iox7lC8hdnF9f4LCIL4KSX6UHitZnfQdGnv8F9aOxD
KqO/unYYn5iWErQRDJv4NFVErKfWa/1qheo16Tp6IHoZIg4FSfg++GWixrqA
kdH93T+n1zBkjcND6HfsE9UWD/BlscDdEgBmpA4PmBT43iJ9PaRt9j3b/3Ya
gtchteLMwwnNRiccrsflMnYgapsb74kISuN3aLfUm7K3fQbUrX/ucupAX3ch
HYXNlO2vMoYslph8APCM1O0IBP/syM+rtrssVsuHTQMLpdpfSprIKNekO4gq
Y1R022zhHMh4i0sizAhgD5vy7fSffGrNFprUUMJn4c9GAyEffS3cCsHQ/L4/
aUiciSW1oeZda+rA48OiOzqJfVI3mjcs/1MD5Inh7Doh6U+fNJRqqjYw6zHe
ho6+A4nb0VvYoGC0Eiv/ufCFLiRjmNa91iP8oaKUh4bCgxjmD/vfo30Ry/zR
9k37hEtQ8TgVr6ov8VjEaeHh7fw/O1xf8NiRtQ88gjLDLmHJl49yTlRqbubC
Dfta8wwReLzhH2qvNEqDr83JZ34EsTpv8GATGhErIfE4C9sqGo5erZB18mfl
C5vlzUdToBfhCoTbj1NazNmsOsB/X/UvBFH8I0B+Uh9JF+vdin4xguqv7Fh5
U2XPJ+Idpt3esbJMcWM5kwZ+ps9Fk/7Eh+Casp1Rjq1E3E2nmKisOkyJq9pn
NFydMhfXbrxXdZLUwzqvSg6f9g/8g/j/zOb0YIpkv6QOZWOK3oRMXckfVpcn
tXanRP2/3RiWxOCZPg+Q3mGYXOQdLYzFfmAmsO1v7PevOZh6kR/I0XKbZ3I/
U48KaCNZW+mI96i24vvDXT++AZBVwc1Nk9Xly/0GUNDYBoF/OfzK5CivCADY
8B0iBqDW4rAi38ZHkKrfZDOMbFzOpWz0oMOjf0mPLn9RMv4wwmrM/KQGGrG9
9k0xKt8EgxcUy2yP7WeWYwGqMCLT3lXdJeUrAbeUUKJFOCkpusa8m/ccQX1z
vmRuxo9VXSBkrTbRIQr+c/Qlbyx25gFD1Rrq49VRsmmgX6ZdhqU0twC0ST7o
GuePI0ls/63xJgil8KqBBYB3Sh5ZCR1wlc1P0Mr01odWMaMHLkNg1k0BifYf
CyWOhjRwDD74rQgBDEqiPzrCtANtVWRN8m1LTIFpWEEaqtZ7qVGLW6AjXt6K
sN3wugAnCar8Noc107jvRdOauyc2HW6SsvaayX3RMPRTxe07HO8P8sTsBNCc
VEBrtRcbbc5T5mR9SouYAWU0pX40RS79afONiwANk3O2cKiq5/tQFl80P2cA
kFQ4H2JTPMXu6IXtpHBjHv+pd3yhIly0YhPgkNoEr5xvxJ+xRHR3tlWvPM+y
WdnvwuEMZgq3/ryI+PXhIkAtxjc4RWTFDAJ+XjtzSAezQfPfUxRxHCY6tWsB
bU3hkYbtY+kdNlBFMZLRPOXZa1jwdUwl1NzpG682aQrRxnKhym99JE0JWXB4
BaPK0eWQUWW5XIveQWxB3ImIpn+upgSYovNeig8kGqvFeV3DOAmdB1Ge02Os
QvOxh4hAOdMTNXiBjrC77mA7ct030s83Ic9YKYDt93J9h/AG3he1atpBD+Zp
uHeYnQpa1EQ5IIP4EtUL242jOGFgjjMkkOZC9Du5xmKNyXm4S7/bGahNbwTs
gpJ4phD0nAxlxqvE6Hg2rPjosxmlDAbvkFY7THCh5DIm60aEIHELS9tem//Q
dT8qtjnIJMYAV1GYEpkAaRE56QBCVfDSigveo6DdLanFCxno5dPaYydHbr+J
pEbAQWQ9ItXIJ2PEz4bZjobTp5ll9hZp/1tlzdney/8Qn8p+IyLyaRl8EAut
3w9QUFwknE3+j2lAh4sKJJ0SF6Rc1KfrOhuFJR5F4qCJSYoIvZbCYc6X5aIF
e/wpCLyBv4lqsbMfaP+sYbgC0fUa/kaey8yXZAYLeqthjK1OA44hJ8yJtGT6
OqWrpZkShrSphT8sxLY0E7sATCDwKcyZvn2EkTzksl2T6RKqCcRdgeCBCa6G
g93s53uHxEhGgDBs87/1L8WBeSccty83qawi3yUPeuGXUJSM9ZcICvWoFYZQ
zfZkmknPpSkk6p28MOdZwR00APcqmi1oXLSSlvYnL0wQkj/ogTjxSmLTBxYf
8pWM5SuTh6Bc05dbVk7WhRca1BsuvnL0xNxK6qOi73pPysOwH1cSxrp4U9MC
PNptVZBFaz5knXz1SP50xvC17FgjjZs/z5rf3YhSGs+wQPgLUX4FOJmLwqiL
zunCCjIeOIHsUKm0J1DsXpDDBsILefbYdD2QhapXa2msa6p7ZsuH2Kch+en6
CC1/s3iHRXwPTKgy0HUB3s/PsdYNHUOOLn+rnXf9QZSfspqXvvH7Advaxjew
WdIeNVEczjz1DRMPPgztd7e3n2KCLSucJOXLl0IOifVZYXeb2B6UJ0ZB1V5O
sj4LCRGAI6xEz5BsyFW2VJgvxVpa6HSXEV5SyMgISP6LlDIOMdxGvmvn5zBu
O9vKjCffz1yl5afOEnZiI+jb3pbYOyXHbjtNWOTe4JlQrVtqppfCj2QHZbth
BLf5EvjeYB8s4JDGLTMJ7H4K8Wn0/253d05OmobNSuen9wKTJoDhfY0fD0oC
E03i/JJlfm1BU6hDzwuZGuUw5Wgdy/Fr4OC7LngWrJ07mDJrgSVHzFPf2Rrp
6/GwIq+IqbPBsRMZ+VE9vNnIOtEkZhAmKry3kue7Jb8nVF9tEtJPtaWZuIcs
uHFcyr6TBi4Ww+Er6TVGetsDlGUiiPPJTiyYa0HsCfXFZdkfDHjAAMGEJZ7R
gNkPfz+2PaC78YlKhqriBrCs2nl6wDLK9V5/HylJ+19NmiTHCiT4Sv9XxmJd
slzvAXw0IurVRSv/tRAwpzld7BzqYbU+IZHCXaan8z4sXGQh08UKVtM3Rlig
tuQKfmMnmCOrhG+QV7dgrctEY5CWb70A6W3E564mRu73Nmsaa9qN/xEeWkcG
QDRvOZcuyMbFKps3Dg9y/UJo6qQ44CDkTQI6X1h1k9MytDuzOa3Ok69dRc/P
WXy3Ayf30B+Vx20qSdQB28/74T8aSQfJoSWwf0hsLR2g2F+6LdN+cz43N+DS
gF+vjg3pxL4vac9JC5liFtVLDtAZs6+tfAKqw1AA7kxWUnAwoY7Ngw+1caNE
wT/Jbejk8AKQdTIoo5f4ODFlJMrmQVHGauRCSi7tj0zCZQtWcTBjHciMqScU
CkFBxdPTSLzeAeAQR8nXru0mXk310THvejXcMSTVY9Z2riakHjtkH9XgP+SP
cqRIEWRymfvwCQLdMmYqU4E2rVk5HAn6Iqz1chDNt0NlBLBcoYm/esfBUU0m
ydEiq/OIL/rclH2Y0kgcBqd1cG95knEqK8Bw62fjmON92VD6pU8YXu1VoxFC
pGyCVKr1SoXpqDY9ZdMMh0x7fL43XZj1DuGqQLXU3oqbCo40n5K6mjn/UYaK
o4F9MSEE5tK8leWVLv5zTzDendSaqGH+55ZIrS/FwDRffPeaCCwFcQ+gsLN+
4g8K8Z4X6OLxsZpRQh1PYc5++SGzCwIvhdqbxSjB35orcFsJ1xo3AiVxmrPH
JkMR8pWv8wEnBuSYwjzjZwbrXeszv9oU/cb/6SYmxPWWZOjh3vuO3SyqlkuA
FurWIl/dthvKdvTa/k6EXN39R4GQ0pshUsr+vvZUX3uDrF8maAEl3kme7Fz+
qIlyoacsllMNxKt3VabVEN9oxR5DUtnMg0OHsWGk0YxSGgLmDymdmZeanlKB
QL0itajIaIMwyHgntPu/sYC2aVKXkDotHVVy4vHHjPTi+MIKJO0IiYgTzOHM
DToX5w22rSt8zW2kAFm3zgexu0b/DtK4B+qvze438rV9uVZoGPqMGBieiIFP
WuN/Gfpnon3EpBnBgnEj8XZXKbSZqnV3lhxMbAsGYCMGmds9d0KU6GLm4cC1
THmkTdzXiq+MnZF/dncJShEESbXEJwvIy8gVZ3QnlXdtOVcmCtNeNlJkN8Rc
O4dlOXsT2aXRXxfwO4FiZaaQLBXCuVvTkYkUJzuLkm41AC/AswGa9rIGRqT3
WK6/76Wvw0ailpKrLpH424AWbIJN6PmCSbpaB70FMFj4/yDO0Bwt9LVGiXvL
dNUK2Y6LlNtwdfnyMr75praDwF7fwNtysBrHGXM+N3tXnewsigdu+WYzuP2q
LTuNe9l7Aen0WDJX3/U1yDcTVvyVWED2p0O3+GYmHDRJuvELvQ7xlZ8ewL9y
z9wZS7JKwtsH7MpcIAVv2Tk30VQpQs5SSyhbcP/2BMx+a3jijScEWEmm/cuB
aTW1fzD1yizaxF24VLNnDcVsU+LHi1eW8D0XIKMRaQmMHc0aHNvjxxML1OfU
S/8nhc/4ZWISzKfAo0igORY7WA7xaZlnjI36OdRMK3kOzsuVzSaox8gouLRQ
vbxkp6P2dbWvs3+azji1arJUyFx2ewWF8uv4DI9xR8osOBSHkpUAijwM0P9E
LtnssVqsundERTJIOck8ekbxT6e2M2ayZjLOuEb/ZqV6BXwT6A8wbgzUrtXb
pEQXEnjDVt/r2+Hb/69SylrI5DDak/gewiadU/luW+2pUZvwgur45cp8llC/
cKrN/0OqF8XaKmgoDuv7nGnVyTpru4tO2XBexpnzw31ofAuiXutecG99OClL
qadLfAO2BfEpVe1EN2UeD7CAGJPtbeeKkyfuH/YfNxx8VgXR/aTTc0T+3psx
dFPQ8f3P16lCelEg1aTj/4+mUHfxfj5N6e+vJDaykjVAhQy1YJx1wJA4das9
q6imo0jg3Qr6OaiUu3G/MNPXds1sLUoq0ksibWbtPKZRDcKftfvBkiI31ro8
JBl549qNnAKFQcGaaLUG22lplZ8LBVKF/mNvZ7JGdyN5dVSvlZ8591NliD6f
4/KpDO5dlUKel+oV1iEhqWmpBBUu8srlDDH6M71VpXgUtrDul9OKd1eAVUGj
TeSX9PuARLZ/f/qPlrNOMw5uupeEbpUq7A+yMihYefwQZWQ6nFFq5t6M+giq
ehr5QkNJSUFVSX3lJBWPYLtlpokcasJGAm2HI4PynB+DoKnWTpX+kkOyPEO6
TJ/fG9DSAitRfN7JDRNtndNTlQxT07dNTMEdbgS2sE7Z9tXQh0x4tSWw4/F9
TaLdbtmQpELLo4x72yThChYPSDqWfhEWkxadaysfjfp2Am1diPCTvvjyBbme
/46dTLxDXnErKmVpvNX3iSv0XbTxHTMZXgiiqmJ4Ginz9xoPQsWPB8CLVVtf
zuQDkW3Gyldwl9DHCM1nG4GfI2xtEJpWcuWG5G3nMvB4ui+6+SFzcQVYnaGV
ExyWlyNSp19AKKfuFABgDrpafCCldnX5xKkNWiRxoqfpg3vEOIihJ7dLWZWi
Wyu4xQkj075S2GfmorydDcewU53JExO+x0KrkPA+RqNqhFIC4vL+qp+R0dTJ
L5yFa0pp4INKDDXBioOMUp66WBf+zy78y+g5VyvIUSjQikulm3s1Qi1RrLYf
fTLkggdAQouiwwwATb+SFJwH4pIXUUqT7v5/OEVGG75waWNnkAWcmIKEfloW
ryhvFnktKSfON6m6KVGU12uO6O1cK/SLZt5aRt6+j0gVa/ODm9VRXXq/brgg
BM9kmScdiRkSGXUJe3JU3K4T6FI1aNTDzCbsKAgI28GaKVeqTDUmcoIlOgWU
u6jGixln1+fsbqetShxrMnFTSaGgU9paIbXzDVoLjYdoG7JTXkii1K/7tkCV
b0uDsuVcKCeo88g8xyrdtBE0N6hzNoURRwROaobMdUPaWvvCdPKHljYEZG2X
aPp8P4Orc6BCpTfzNlhEu+ytcws7Dfm7CuDDDvR2Fy1cDMbLkQWjI1kLc6lw
kXUvIyd9dCHCscsMeXGlZL0+St4e1RSGasKkSwb51I+uLfFbZaC63RfYZAwd
+XErERXFrLHh0vhTHROcnUtrO0uP9ojI/96Jb8gV8+ROdnWpFiU/QRyMc8s1
fCQ0eMhb2iOnM0vUy/7KWTAKR1ePG5uPw9euZg5nMO2J3OSDwr0Zgl591nYW
PBx3RSl2QhSmt09nOLVQotI9ntMp3ftsIafpbEy3uffYqHpdYuARHzb9gUXV
dBU0qO/BBfaCkyzbsQvcRcmL6nK6FQexdbUGUkgQQRrJIsyETIMMJJTvTriM
xq1SNqJrd5z3+/wCRq0QwCwWWmjRkQWPwmvAp2qSd9rlcwmiT+TJY/hQZ9rk
Yu2xqU5KW7m4baKhAn7eKDfAaNQ1q8W6WgWn/QdmRZzZ5nsmewsrlYTke8aN
S/iPqimtUnJK1eBqr07y9ZsWaGrVUtn6MtUxgqUf+BmstI6db67PLLuqj4s/
mBP4yHQfI8VqQBy18KsWtVaJhndmScAj1C71dIjebIprVTxJZS5hhgwFQScm
8LJbCogCiNxkQkk32VqX3R+j9k8mhvQ9VZBeNz2P1x9qo2VPVr0tgQOfIR4T
gIEMCKCYz0IOznjTXC/HZe64fxylNuHdhMVUthOoXUtMRRH9G93lKG6iIKQQ
zMP7MfaqdOBchMRbr3GS+naD8sVM4PIbDuU0wb9w2uMfT1CS7hdBDEWcX/d8
6m55YLtJD1kF4umluuZTLoTKQzDNXmXBxr87nqLkA+M9eUdQPaRxAQPcBVCY
S4iQZEhrC6cjAgBYBzGDXOQXy7lCN5tnVGyiekNr2D9xt9b88ZK2pEr67t8W
VgKHsmVjeNh+uqXvH4lAjmr5yiQgzHq3YiB99MyHDaVV+IIavvbt9jyZKD7W
omZ38QeR9gMQbci19/qopf93HoWsI+C86wCLSa6ur6qDGetFuXdMWP8uGLfR
cNZQDVSG7DY8lyYYUWka0hRgJY0H8+gpdVmpTBAbKJ1ygEfbYQhm8fne81E0
GSkERrtnkT5mc94yjBF8/C0FX1bKn74aBdETR2tDOnjlTttc1GLZwsQx/4Mm
vzWFievmL70EhvYvkz3mz4PuHof/StkVp4mJDYKLNTAE7VCzACQtZsz+rFKw
A4Q33DF1A+65CKh7TLtGNnx7PFYoRHnB/OcbffFTqdqnsIJmT4alfAaim8C7
+bpnNAjxusX6Zr41bJP6UPNWwVxlgk9JJlIEPNz9SNLpSpftvQbMFwVi+Kga
LLq+HFdu2y/8sM5H/a9Cn0PRiqHPVYZymCyXCJAaEgcig2DbSI9B36MfBly6
x0pDVmrucCXxsJ3TOV2UwJgqAYbOqljqt6vNgrNW9ZmBFSyjWU4k4laVorev
U/WaHTmznyv4M+ojNJiPhxUGmP1bxFKb7sZebu5WmHE4X0JxpdYoPYlTSgTu
ZpyRG69QUYxM3KUxZnaQjZ+fdQKmfTZjCI4GEwEBlih5h5IfjGGypFdK7Ovp
5Yz4kpKqbxeVwEPXOMKz5t2doSkHrItSsqrNTNRafTrUwbQ9Fba1dYRwiRl6
04mAOpKzUT0zust89EXdGtAYIjNOsOiCHWK9H5s2v/TsHnKBmi9MUNQkXJz8
5lsg76vzDSCBiGr2dAHCOWnpy1MvB8i9ARuMCjpswu/8ovFuqtXMYP7w2PTq
PI9/oNXcvPpCxYCfCYzK6FJyqktI9koeS5bAgX01afhm09ZieBriDk8oda6u
37L6LMSd6d/HAoBB3+dMKX0ppNC6jLlSmzVvE8LwYZwRbm5+L7BJq0QWScWY
jzJBotahQUHCI7XJ+AYM2DThLI2P1u03OBsXQlVo+ucvLXhY6wey8etKssNB
HPTTIeK5mOYXUaPY53dR5nsRyMoFNUi7TKEUV9YwxxVHo/GkCAunINudgqJW
TRPNILrWNucvDLabnMW8019utd9UfpC0KnSderWnMN2Yry07txePMRwcxGgq
swCq9oDauSHxeTk018vfdTAbmj5//Zcar0rUS9zzUt/NW4OKB1r4XIZDjFiC
bkSGjPJmUlhCuQu/uoX+kIUreZk5GxpmCCwIH3mHVy/hNyXCRXUaVF/xBJXp
TOu4/a5tTom8tm/IHRXHyyNURNnTZaJKcq88xx+x6XFk6n2mVMaakZDhe2QH
N3kB5Yh8st/4zqmkfRJuedweh/oX73UPCqcXVw5vlOoxpO730sExdGgkOzba
JPrimH9vWf6jumDdatqK7bLkUF9UrrtqdLRnVQOAlGg8yldlhPVCVY3O9lCx
GzJ3+z0VGx6SXXhI9g/d0swerYQy+Fq4h5kLSFcVnaFAynwfFqz1rnoOEYVN
pgWysyHGs5cEYmgE3tkUv0N/RLtrzwtjcWUb+sdnWIEHfm0hKB0GuivyjsyG
X7XkfIuoWwrvBO0KOH3UFl7hadVhgBXD4yFk58XzI0CHob57R8UbCqnU//Bl
OEJYG7hOZnSGuCIYoF0f5ZsN9Ino/GrHBaM4kO3vuPp1wzbMYc1OMempOqNo
eL7Ze6vgNvYSuDNOkTi1d5UYwsj6e9MmDZdkHd31ZRaFKE1Ue3zEgceap7Vb
BR+0OFhq6e1QR9ruy5LTGkR4K8sVHsXJMd5BYvr2A3OcuYfVxbeTn8kIWFiv
L3LtEzeBOwfAYcmP5Ea9Y0pFh8hqA1XGwKN3GKfoFD6Vfo0ciFYL1/9EgDXt
QOQDLB0qqPIBYjk7Tw6rmoIQcd280FG/aHaVuwfIWGwTeWe5Z2+nbSaNeQJX
kNVEbjjYw3x1bGluNBj+LQ68b36lb51W1CnoPQ6FnNJNXZo/QMB4fokQVBXJ
fvSefZTngEx4T2BI+nxr/SmRhNqnom/zaVxNmm0+kPYAd/TA7F3+3paoO6TG
XtmhjHjjPjHByNoU1VKxLK7T/uEpNaNpiSE3cQypaPOj6LHwiumDOB0mCIPC
bW0x2ftOz9MX2FKhkMOKpjf5mr6Eu+WieK5e2Lp3qnhJCyL/APr61dPh9o25
aSlIlaka218WpN7Nt2jX5AnaJtXKy2yWBAKpqEAtJsypKOG2VyHxYRCdM5Dl
cnHwk3HoGrWVMn9t2GHBDv2qDmY69zlSL0svPYt+jBBjvydSuGjlmPy6ncWU
sbFTRahInrmVGsKRXTva4tKIO/EdNIZZk1EFyACI+EdeUM3+tLp415i+Cjob
Yy/UzLaa72f9hobfN7xxxZHk7JN+v8IKIuw2oOeRHH/v7MoWn1JObouCrz8t
7rcloYegaSbgxn50cQZMAKuynIghfF1FGBTbUNcpXH021uiwuxhEQsIHWORr
qu8FUCVipYfsq9Edabm2aGpA3Rkqbk7FeHclEd/NnsFsAw1UXbNYRGZK1Jgk
UCF0eV/NYBudHylUhx8SjwMqLNVSgQKutPT45W7ed44YotaxDowlzXlbFC6i
W0CRHiFXHZqW9NYJHhtOqJzp4OvpGI0a67EuiyHSNOa66kJgW1MvtFPvmg+N
AKN7/n8IyfoR7rvRoPs9vJ7K+F34ebBmuMaKQApICKC2WFwtylrlFys1zksQ
XnxGZrgy9iviJLqh837T/gTwD3Zav+3XAeLmntZbWxWopcMopgF5IMaGACFH
lDLWsTm0kTFPIJF9GIiPQvFmbS43KDpRlViBe/Uc+L+V8CKpnu/InqNd33ov
hUDkMLFy3/7loXtgTAin09yAdZhKfww/cJL24TC8fOUm/2rB8FFr1YfKxzEI
s9ac52/VCr0g+mwzKV6BZWOoPBQogZgmJCXeY8fz7ZnEZzjTicEhCg1b0MoZ
ljRYok5VeenNN1K2QueOXfob6E9ws8ilg7uQFfUU9pcAviEdj+5wbxC6qVJC
/INXCBzt0gaYb2kjbshOSGxZa7+/xpneOaYOrnmZ44gr7h8yQLrGj+uxK+01
wSFRJfQKGZfJcImczMQDBxTkHnIYahGlGPV5FpIj7U7Xvum5WGkfDtfRr2Da
QlJcSsELKKQwsZJIA98VU2YVaE5r4S1D2NIugdBWNYekgWfLk+NSQ8Nr2ES0
Zld4ID63XXwM/D21LCjBcwWhCWkB2LhUhN55lPdmgJuGZ0Ot3ijkjbcknfKY
3lyuXeSY9Z2aTu52sqzsv/JUFqahcGntYMIR1mjxQE3bJ8umFu5hvnj8CWYQ
ZIlyIvmDmEvRbAnEGe2CQppiqyfOZChi8eVrCIU7awEpjaBf5HN7NTrTGpyW
ZBK1uIFLSpQAFxz4HKuAR6235poCdfz6JrE/k2lnxjGq4qlV81yk86AxCS6o
B/lFCwGd3C2PuvEoAtFWvaQmoH7z71vZBNDs2y1wznqV8EaH9m7kpuNLBnox
wFvKGTwunbIzXIKnHItX3EJJgqVcgg3Lv+SVX6/TNsAWIVOQ3i4pv2wpWSV3
R1VwWDje85NIZtZwu+0Vx+M7FUr75oB7hhe3ih4xGf/iHRu3TtUzp1ZXQZP0
7E9gj/x95IbEDY6EnKWtMPvLQrTMAzg3p8MyEoDwBigStWIs2Wl4LJXjbAOQ
D9kCfhbd0BbT1+Bd1OAIjtXYyDeZ4r/RH/8bhiWsQtR/vNyqhXLH0EjGx27D
+kTZJLAgEFdWZ2WZov8RlEVnw5UoeMNPxxQZaSdpePMAolGy5wX/DEj3r0lR
YbpU7Epxdjw+aO1IBYM/MqDQIdwQhKNjRyPbrp3AtEXdmCvv9Yt7JEeJueWm
DC4Ga4YdXiXT9gR6nvSLD1I6xai4Tl/WVxG3Mqj728qPHAdLXsmAP0ak1GzT
7jzwG2555xiNOhjSINcOnW3c+Kr+zeFa9R6KhQm2vMNkYEeHTMvdBwL4ihvj
mxa/PQzc3Lmpl0Rd45PnBtiHFIR0li0VALajNVX4xlFJKYv6r58reEHsZ+oi
TjnhNCivKL10u8nQGNaT/62NJV1iC/jH8Zfh7gjpAP8j/Xu4xRl17WP8GphZ
xz9CzASGqq6hBLn2eA58fsMd2nm5zMAjeQ0Azz3LOzNVRO7pmGUE2LBs5fUk
b+qsvKodAyV/Y2doEGHTHrf0fmJtpgvYMaVjwnBSKT0Yzf3XK4Yx3zDtlHSp
aTJ9qytgmRQKtPggRNXLj5o+0+qBqUOoMeOBS/UV3AyBLYGKyIhYWzuWrkYF
h3Tb/FLGQYVG+5viObISVhKLNcmz2NRKZY+rkXdAJziuvRYH2ZWNlUMEmk9M
18nA3Kkd1LdoApdPIQxOs7dQpSqyThp47L0U0K3NFChDD8f8ASKD7tJk1nE1
lwR/hMb8OQxXIB6YfV9sJMQ+sgqwlpQbln+aTee7N8l7mHgxtXCTrioaTxi5
2Tn71OraqN04AAWlzZq/wALlKGN3vupeow4U+YUKfr31T5fWNJ1lLcfQPIeN
eUBl4Qi3KDTQsscjMrybCiSBSoDulbkjmQxDBWxhfzuqN/6nSGTOldVpAp4o
ZNdSHgGVXw/OW71Jb3MjWwmuwOZ6TNpmVss9c4BC0eNPXhphtUcBIXoOzyC+
pJsfXapXslkvirYQ5qHikuRgiVn73u0n84nx/yDqrN8AC/EvqWz0SnXLuEhb
Qje9YqKQAh5Sb4cpxQxG4WuM5UzR1dNVn8SICMB5YSgJntCbKnGRG/r2QTFo
tEcr9Jnj/gbGsUR/cdalbUrCf4C5k7RoVzIML1w7oR5nunZo9AxErBiuvxAA
mVL+eOaCz3luNpAOLVmL2pajAKESbr1GIRnDcceCkJL/blAnZIcGJEMsjofO
Dh+A2Ya6h6koSuHMqlBMxvFeiIj8DQThMbeRJLqdO4gT/fLRKFZ0YPFmy89I
gaLBnTBljQQPFsWFXVbvs2TwdOTrBFnLTLJJTo5LI5Y798NuEJHrUdo/BMJh
QxRyUbXCRFsU5PReKOPtcWq/LmahsS2gzyTp++SQ/EzfkzPSS1841TQZ4wtY
pAciPANqfhArczVp2uqGlzZR0tUiLg7TYgJ19z8dBNZazhM1EgPHJFkSZ5tp
Rs6IGAYeZ6RQvk96gQ5r2/BKZeqZe4giCJ7AozObyw4gFqOiPh2e5OoOJWJg
45kwhUI6WYljkSAwsQ2tLcvjEi3yks87UebuxB60KrVXRkz1zj80cI+7RAHa
dmY4PWD31rZLN8zloYnJfgQDalcxweMmMsres78zEuFvnlxGLsBk3W6yJXkg
VHy4rzL0shlTiPTBmPlGYVztLSlMtLhq/6wNjq3Z21wWKuQJWI3g8KTnuCZ6
/BX3ikvwzh2p99aCF4WE4S9B6gtsp8lOyvL5h78+fzfDvvmWm7VuWtcYXLj6
DMJgLdOQnjC6DPnCwPNH87OdM8qy/XU4IF0/W+5gBWVOOxWRPRvEVCQdjLUk
bMPMHU6HilXLtlGpSHbtDQsGnoSVat5kBb7ik6/waoEWcbw03wVDaG2uWXRB
t1ZhvfZr1t4qnO3jdNE1LuusRzpX8XLrFcAwJBT3NcCmwsBeQ3Pq9yWNpKbH
ZEgoLr7tMsNoKx6Q0Da/yFVCjJtPuAtjzFoxZdrOV8u8o/OWfACaaN4CAhjQ
iygRMVWx3xdge77IAMwKH7r/QongccH/XnJrS9/XcI6645i5ShvdiKJIHSm2
GxCXaAxtKhz0kzc4hP66kA9YlRJDkmNt15d95ywb9D1TiWCupKby8XaBoPwa
Nd3ZC9077Vt6jUBCve7Pj2aPDb21YbncCzQWwNSFf70tVYP3nwdbff3JMkLV
rnyIHCC4v79yPk3438+cxiyjNfLY9OY8Mhoz5e/Fwp7PJalB6XHuMvxLIBob
clkGoQk8rTzItZGdEuiBDqUVgI9Cp4pBmEwowszt4Jz9jBAmLXEOUhpKHVOb
LRiYmL45ZGq0TFj0c9ComaDdBNliu0nx3snGp5jZMn6Iz2BNsPOxM0MG3NX3
pmwV+b/pLgfRzG/07kU4t4wcJbXFWAQv1JDgBhsk9PnuC3i0qovTmT8Zd8aU
jFh5mbPNwPi2S3RH5DnMVx0rNWJXEZMG7W/5ldjnnLqW0GzK61O/7kyh19zi
3YbAkwxZzRt1ktpjjvRUoMpSVKZmV3dwfGKCyCoadB0pRBceOzXrFbm9ZeD0
hDCHPRTSrkMUvjVWiy8TQKnzXg4eMvgdaWKCqJhJtVQZyO9D9RcKKr3TwRTs
fgN2Gng0o/xtW4E5AHPOB8zUfElh0ZKnss1hr/th3fvmY5P0GECDpccHmiBF
VNFoFrlZlfh+KrTm1q/jxwoyHd4u+6cOZUBDDiwI4Jalj6Y/EjeijPD14XGu
OcA6OEdCUc3HJyfCAn7O6YJEjye6YZw1gaMEF1X5uFBzvMSlzdXnMscThxyk
yA4/l9DDmb0APD01X7bGBBFLDtF4Oz8pTIncLFMwmblYSUbqdKh+v3rbaWd/
pDyL4ucBf5VUF6lIjrnzSoEEI0LQz9ZULdgJT9beggEw45uMXo5cjddyL6uH
CuA0P17kC9wmo0V+yerBOC3uvyQdFIpgMtYpRtSPsQpcn+HGYWW+edrdvYsF
Lt6Bu1Tauhm+yCwA6nJIfDKqEDlIstkqN+TBNvvCbfYL5FMw7hnqWm4C2Xwo
Hm3WWGIo9Y+FC6eXvOsxMWZB9a0ZUPLyQw7caHn1zmshyKrIrjvExfxInMQe
JxgPX/rYvjkPASwmC7B9Dj1FxAgUokjCjRYJ4uuyJU7/KruHwjgWYyIvutVg
oUdBeP95Cj1qHOUOxXl+8oYw5TNfXH8ezKB+A2LglVAzhGpXkFFRneMYnskm
VQNLEM8HnIWRyFUIWAbNaPp2GaQkK76u6+PRTaBhE8VF+EjytBIox41puass
/seILnVGhPiqtaGJ3iqXdjId/cItlZGleu7yHurA7gzml0D9UVeFdve81ZVd
GTHMRzd6P5SYu3LL7RvrhRvFBFzisqcTbrtmiRFOeOrbvOC4py/lhGPJ3VsM
x7CAZdGWeY3tltbz1EdW1AFzOPDIMblIegW0ZdqhwRh3EOeKYDdQ6PKJNG7/
P29/WeJDq2IQ8kzANvwGjc2YG2WDy+H4IE/KFv5Tpils2OSEu1MXgnyqctBt
syCv23NolrYZbwjz5TxZ2qKA2hIaiGK6j3Yf/a6IhrLOYTuS0lGHVNwWMNqf
O79W8lAxLM6YW04mMqTTPTYJe1cAQoLYiZMa1Y9bNrIql+hjeIlTtZrlpB2z
qPIS7JncbAdQIcSjIG7095b6V0hXS6VSkziLNVIsPLnUxbe/HXwlXke+HKBL
2+vpD0BC5dbM2s35y+EWR9IShvP5Ph9kaU2iVUjtn/jQ5/GvTuUNsVSoft6f
OP4n+J/OjJN6NYcBumkCEqDuEMNaL2XyWUtb3Zi8EB4k1cupnaQOU9sDVQX3
eoi6HPZ0LvoujGSXKXmXhxBgnWk5jQin0O5VLlJ7qZURpadXGD6TGAPNp3Wf
lMH0vb6wigl1vsLhoEBacr2hTtKq6sROFl+fy1dHWylirhij4c0pI/KPK4fZ
vGqnHq/EpIZoONQ7W64KUhtfLkc8xYoHaPivAvZwSg9w7tzwPAwXtQnMtI3n
fl4XHyBgvar2T24GPGueabW/WmsPE/vMZ4c6qAl1FtMOLwgZdl/rZTt7x45A
cBSOQQFJlkYE2ykHXwvEK8JBXmjTmZ7RWCk3Jtg6Oaci5HH5X5vWYPt4WPFs
II8fZ+nD+VR12drjAKTucjO7eQPgMOCoe7s77BOs0LT6hFDVfXMOdn2qYKDH
ixNEdrK0gv1MO/+E208Vp9rKWBKfHM0YH3KtKsZRK8E7q7bX5mQCysCznHQP
Y8E7GxtaSq0/+ybqnfJf624HbKxcolpUwT4bZ/j1R5SF5+mVSJGCjyA8M9L0
oVDmUuf9oNoX6Ayo8qVx4ezFpxQfFkEgNOLqNeMLdHv+zNaR3u74uUmvKnLQ
bKUvtPLAJG8zXRuTbF6dQjgNYHVDKBPh56vHazCH6DxGWds4AMsRdMbkDFfL
yDHaVAEOURdwA4Ni9FrW35tbBMUrOQf8AukVtkjJPuF7GSCdHC92FGC0E7g6
NN+BpA1dDhRSzTfgHYKFF+jVzvREHAAb6xls2zEW8Yy6QkhECzzJZNYTlQ7v
EbHQ+Qp+PyJOBaCotd/ZlEfYwMrmuGgPz1iy38reFDAOpyXubtN5824PKruo
Zo4OwrxYT0111OiJOS29q6EB7hXTNYhrTt4J3SeZNRsKe++Xnx3U2VHbP/KP
82+tVWlyqjGndVFxtD/as6nmcfO8dH/YYMOtpHdBOm+EVpUH1bs9mscTFGJf
wsilxwJlWRlTuB9qWYp5SlPmV+PU1dlaSATqFdPTnjediiefF1giAt5Wua0T
SAlwtQwai0qfANgUhKuCBNcjHurS3Abs+mtI6T38snsNqHU/Po44C5fLdOqm
wjNKFsy67An0pNS54fLhdC6DhnuoD3/wOXl1Yovkr3/lioMwXKh8ezMp6FBQ
LSTXSCKXXwMz1o7nMYfSvNmSn+WppEg2ZLplz39Q7VAK8E44XNKkdtgDXrVW
D2iGWceThlDonnmbPvQUnEjfXy8jGTwFxrcbYmg23jZ+79ajOla6xPtqgtp6
l7q0ElQadVSWKw4FqA3vnq9BFumX2BA1ozf52Pv6Nm5HyECFJSwISrBaMTB1
sW5VcdDO+92wLTxHF2JIQTnCjv/5Vv7FNCh+PCSJK5/wUm6EXubqeJuoSw/e
4kaOeucJF+UnW8+5+oaOOGxtf+cdsuqW+7M+1kN9cNkfi/c5vnDhwTmVzU+X
lA9UMbDSLJDpSRa38aTZCP/1EcE5qkD4Gl7d7vdqWQqCWfQP/7zevoxFs7ge
nLb2p+DfGAGZw4QvQqkn0ZbfDBpdu3lmlJn2EuIq8hw8153M9IdLz6nnpvyz
MJ1wcYlbWVzUOXbfA4bhCo3rAHi8hKMzyiXwitHnx7J6T/yIessR/XfwcqDH
oXPWgMycde/6gLzshrySgrTbeBvhoNFMO+BKMGIXP/fnR9US3S1SQv8+V8fG
vOVMilvn4gw+zWQvJyabfc1m1Ljo/sU8+nh2FTl00BZQEPMuDo8/VXLAgJhH
ahmumd0QphdsBJjw289AsfH9wEZ2zW8ihrECfBVmUQSvDUcpzoEiYOvdi4vW
yx4/KOKiu6wWFaOnD+DhU6Ua4DJjL7wiWKfXHpYzI6tOSp522KyKrmF1E5Y+
wP1PrilisDYljOkyYGmFIcVgkR/SXeav6+pnui3NXdjrIX5DWwFtkm/9SpfZ
AJVfDkoK9k294OH9V0U+sRrJSaLaphOv9vThREenanr0F6DbCgbK+M2Kopzp
vkdgS7rzra0/MSBEiBcrok6MdBxYZhraximupCac3NLr5LfMC5Ojs6CsDymp
RchEeQvBn2W7vBTPxWZDdl3uv6ItA5VGpnMDiywENG2qsro5eGUwipx4aVlJ
ynuJ6tzDCSW4paFpucYF2+E7HA1h23zEW+Rv/5PRZqlqWU9nKIuLz3BMaNHO
07bjeTijfA/WaEnwpmgBygYy+M97egZEYi5c85HlOOvpr5iw+lE/YQfNxj/l
pp9QN4EeqBpI9XYxATxEuTIMuScyG+0RgG3kz0WJIsZu+kIqyVmUqOdzWQMs
f0mGMBAbecuchm3WLwI6UidwzJZS0BPoQZ7OMg3evUvFeIsHHhM4/WAPPZl8
ZPUvwc+c4sB10kISfq1xw0hlg4YpWst0N7eq98a7IQo5ISKYXeCx2dWPdLRq
AzUO5lYc0I89/mC+YaqSYzgLOJrZcv0368K87mSpbyCmZg3ms2ZtdElhIlir
Ssm+kk42RtVEB81O9+DyfmauJNUfd22tGUEoIytLk3uahv6AvMFhGyMrHoor
TuTfSLMQpA3AyP3d2wOtCXj9VQawP/F4VdzAn2dN/pgQfs4zQ0QrdeSHj9mC
bAzRhWTdw+PpI8+0k7yrfZimTEYM5A8zeB85uToGaYpDHsAZR+wDcv3ud2G0
QFD5VnD+v9E8Nb/HYN7dOgvhgcHujumwgjFCx3lo0w5ddlcckDoLFWQtWu89
cJaIuRezzm6EPC2Wqipt+0Jl9Sd6L9LzwgxoZGgPQ0uok4Nvnkhl97GnAzZe
XKP5ZDFRHmUPI3sOX2TZzAGcvPWNAXdtaJ8HWPzqaS3OrGj7u7xzc2vT5e7U
jDkeEkXcKjYixJAKFZJ1dgxjJBK8MsPPcmiLPAEQUd86oGMZcin3LlVaAVOI
w09kgy8KZRG+AQRw8rhXR1wlAbeHlXtbI3aS1W7e/UCjw1YkIrjJq0GwRBDZ
Jd6n7DFTlTS50gKc1+T64Xs7i+0jfOaJDzCec9PBdLeYct43bXB/5mdkGytO
PsD+iPlz5FjrmsKiSTt6KDDr2vh5KuDBGRPU7+5BlhfB3XwP2WXBmvOU6k5t
PDOgo9LsRBTT3r1kgtBMqRNSKO7TRGzAP4dyt+6oAnRV60avm+EedC/anjrm
+3xYFzqItUV0VOisDXK6cQ+zKaXc4CuaVac3GACn+9wQ9xbnhuL7LhkzXu+m
9V/+ZkkNSu4a1nJEAS+eAt4oaMTSZYsZMXN5IYxgrPhELeZVf5UvEQkDySqH
C7JXytVRDJb/SqkSoVIjDtMTTNeoE5RtOwuZDmg9Szy6is34yy/FN45++lch
DvHAlKpCOxDdouc4U2QYQUcqLkQvWMBKrVBdPjeY707Scr3IA/Y3o8W8NSWP
4scnV7lU4p+v7xfo6b8mCvoYrvFD1A7X/UgchCy8ShguSV9Q6BmRXJzNGiVO
yWgdILH+Syr8BNcspBvEce1GhmD4P9WG3IRg5b1R/rKuHPSg85q0kO9kfked
OVUm9I9Xd+FUqDXtQeqVzF0TnODlxJClee5nCBuGmcF7njUWbu75tEXmpsNY
KHfBlOmpTBw7jfTwiBynAXXj37ej0QHhIBgPGvpQjTqyrpBvYp2D8rG4JOep
OYyEhWpC09iNGcRYIvB0ZNlyi1QguX/iU5Vgsqngfg2yyHrT6aZmC3sA78eK
t88g5522ujIdWUjEPU8PkbXMioUPw8NJo//IKCshTBpdW1SFbN4/SD6Dh5kP
uwUd6vXuln9+TmY9hY7xhPfGqqPxPgiNg04FvmDwrr8qafsTdOd/UOxjAf7Y
NOtzIJS4sZoMcFDtyVi6wsJ85qb2k1i7ykHbtG8usq6f8hY58UHrUZD+51Pa
R2OQVPta813m2vg68V9esdKBLaUepCe73I0/a8OU0ktkQ/1ORFsxzUuxxtAc
qEVaENasR7E3Xs2LeslSk4jpPiGj5OgdIEbr3oSw9zlVvx4Eq5QoikEMaWgJ
BxudZ8h3Z+AWc3KocQFwxqVGHYpcFAh+HkUQH6IvUxYg0MdTZ9ISwEwXfmCk
qT9RQ1RGtzOE2omeVMB+juaIhi9pqjPCcjk79hTanJptpDVjnGgI2IgCGysM
sInRQN9xs03y5O/r1CFeVYw4u2FfFK6Ac6fyM4tqZKjA6iG/XNTKsud/J1SP
9LKC+vEPPKoaaGFzEicumrtt75cGpkb1J+JnuoAWiZ4wfVl7OfwN5Bjs/G+5
phY9GMFPGDwJr8gfbs6SV06QfruyoTUfDghokgyQpJK5DyCAJnElO+KkYtAS
Iq5rxfAcvomirEgQ5urWpWHo19iU4u1R5z5zGEMlrAHOzaaWsbwQU/DHPNbZ
Ts8UQ0CQoUt8e0tLmfLW2bavKAXUzhcyKIckWLH/dUnUzrTkWH0S3SIXmY6A
yy48mbLXfaJ5Wur+ZfdVOimQ6e9JN35YRoLYlWEgpkinSEKbce2WwACBaNTY
Z/GO2DPXKJFrLkz/lpmIUw6SiFA7G4TrkYnYel3C4gizKMuC1oc5QSi2x1te
y11KqarnNgrn0v/j9iQjZhLC3bhfRFbMV1fprr/ZJx+7K7zZhhA1m9WYg7Ja
pOEi6YTwmXI3aALQ694PXJTo5Cn59b/9Wz23ywe17l2BDvBpLHd1A8W+TXve
v5eT51Jjo6gLd0z0qmeVZmI0C7loaWll28PQ6Mptcr66EH0zPv6hbhgT5zTc
m8KLHKwEaxo+chBfdafJSp1hq4vQtFMIJ05sDxaQ7cWr5bhV2iZL8mdBxwK2
GPPyQfWgxKgqxZi13r+XCi2Xvd4jflpSw6gPOp4GH6c6FN2HIpFaYgJMEjXb
We+G4LeN67MMCVq7j1f/ebhbB1Nk4cGCYtGq9Uq2IsZivxrcjGwKQ6V6VIl8
SgoNwu+QcbTlUcYh5YDvHW/sWqpAANNpfnnNrkKuHiq40+HmA5Rk6UlKspqn
KnFobyzVBB0FSkNM2MEavDxgNYVA7XYswdsovdIucbTs67/YsYS9iIHyYKuZ
gzZ99fkLmarVCHQHqHdBcnIOFbFeOThzp6uUMMzWKmhGW/itLkQXqLA39BLQ
S6EzHC5MyzQPj/3xZwD/GMM/FObhykCFNNnWCrZdCFoy9V981McyyumF8SNF
b4Bn0iHMyP+7VCb4lN2lVC+eOWobWfzw8I7PLx3ZvSwEtAMBr6StxkaxS5YG
WpobfkAiHZF6YO70p2/DbRgekQRyiPb6PCJUFLmvdiKDQ8zemGAtoG5rue+M
qG+PWnGL9Jo/VRDqYTpHLV8bzaAd0gpNdWMIiP9MMC8X3lV2rTa5VMHF2A8D
nP3KOqHc1aMhqFj27YnCMq+JiyoAeeOptsWIMREej9xAzcK+kLa/t+DoxwLL
BlqDEDPcknz+wO1FKFf0mR/cvAda5eh313H3yHa2r/7gYCySAszDalsvf3SQ
jlSPtcBOUmdxFDyO4fDi2VimqxQwTKD/WIhgBdsKVAOR23ZzMMJsXEPJv4qd
FjgrhIFszjR5tM9+5vZHylqal9kB2Ax9zDUkIPEhtJWsGs2edh1utfBONjQB
aHm83bPPDfFMY8oC0FptiusyNPctatJqtpm16wnKagxi3yBNJHiH6/qW1tIx
7zus3t+kfkHllKgrvNfmKYFPiNIDkhrynpxWhXugRd8sXhnxJgloOcCGCj/B
E7Y4ylFNBOO76jUmNffXRHPgHII2QKnVqTKEySg+tmyL/0vzz3cZ0tcs/lAm
H3700DEjqTaB7ZHi4g50LCVFtpD7J65lG2UQydo8SchWGQA2z9W4hFpduo8C
A5CnEkDboQOTj5tftt4jp7xwwuIKkO4zva4VU6vloVH7mDqXbuVo0Z9Fyin7
4jxHQA4kRBTTpsn4O5IX67qunepOvE+Ai7kXD8UVDfKQQdLvXxTxC1sML0XC
k5dpLOTmyKZba5bP6hEXAZzxmerIIMaUALorIKCZUdZ/+wlzXJlsHHdQ9xhC
84NAQE5LcZt1s+NQVpsfd+uyKhCc+JMQXK95Q27ksGtzUICE+N7grE4Cds2B
mgs4Z4Ef5hcsmTA4ztTb1AyawHYEcxrZjD2IUbezRXFGyhsXs0hk5qlsYysb
cMrqYdV3WRKYYtAJmFThdBQqF4bIpC8s/pScfPRbkyDgwf4VAzJAZG2Gxddj
BMGeSzGZJohGKuHNuQxz/ryHdqctzGU4XGZi5CiJ/+tPAWKRryNE3nHqww/s
XOFTf18wNB83/22cJjDrSaSlfZB450uuWw/eDQiSdqxIA/aKSvxex/J7LvFr
3dIgMCh7UAbOk4DmiRqqc1eYWYQSzplclNKnKf1rzGSl+VW1ADzcApDMXdiv
UedUFdptQQ43jNiwCxQngfWMIAeiUB1GCL6C48H41jnCHNgYexjUPGp0KQM5
byIAQRttkkpS0Ad+eoh7NoR0bhxXyrUJvIMj+GcDBHLmyOQ7i2uhHPkaBbmv
Ks9+dPBSLqfzvwkC9ZJwlf5LE5p5upigQK0V3vTWJN51yXL+G2+TmKoARwve
3UbDtKSPrLOTHR4B5ViHAECgHoiSfWi4hf2OXq9S+Oin8kmJ69/s7bhw99F/
mCouXF1F3hBluoNuX+JCZ/oRzh+Zny6Szi8vfU216mJl4VzTJ5PqKCfmX14o
wBlF8M1CqsIxGBE1ZijKtGOigioKrrr0yB2LgBr+qipMAYfrnM7YmMRuxT6n
EPsmAxmUlYpe2FLkbRDexId5wbc949oMFGdhBQUgSpRyeLp1j0DZjYuwO3gk
ow3lEXEZOAkvMiMmfLyqeWJjdx4hDwrWRgkJLrQQfwxxzwVBhFFHGUgj6W17
Orhx8sGKmmNM/RGbBsFJhOmvbuA9DvaX2pfT4O3z9O7+9dCWGFQSH12ffHHX
Ye1T1C3uTZnEfJliHgl1a0M6gD3H0wSnvC32wTqcQzdj48coHhxJ/M7qeU5v
Mi8vjcWQSy5CGGwbrzoYo/8lMZENwm6m2PTK6CJLgx/Q51DtI+VDbaMV9rX+
Ty7y3lb2gd7/1K4mRZRieAYaA/FJmd72i3k/9HhVmDpFlipDXUNrmeyohAZq
HeE/ayYc5L/gi3etdoif1s6KB0Cum8S+2e0EF6EsMogtyzxnSp5vaxW192sl
k0WkFe9Lof7mDpEjx9I7nJKLKyLHx9E3xnyuOwfLqMgJdEtwjyyogwQV9FnD
Orh5NbpRzLu0Zi+5iCDYr80rPKuJXb4MOHeCGAJI3Rfk513K0jiBNirtUAwS
zN48wXBsa1K/TaRd3ZsDgZn/42+1qYPg50YknIffGAAQkFucFt3WjHFPV8/9
rX3kW7mAjJtHFY/FBVYIF8CL4Q8Mt6Pafe6VAjG2u2r0tWWEmzYe9r67PunA
JAiGqs9+IBqzmO1/mkrT/PHsL1TNGDZpapBqBmIX7Yn91wcIPwhk4yIP+Iy2
H52zgk7fSGLxVwCTXJHMdf2+dTAAO1UGek8bpdydGv4MB+wbhTRmepMoVxDF
fSy1fIapM7f3203KqMHjC7QZosUBtUQLNM65Mj++zie8IpvckN39Fe6HNfOd
LFDXwcv9oQwW0GAc5txJp1JVDBZdZXaS8YeJt5grmL1TfOxpkPM6dSVrQLLw
36VJuqI2D7YYPoMpR2a5jlmFQ/MOOxhL4lxgboO2hWubdgUX9XPL4oBokPU5
R7XLRwa9NQzVAnixm1joA7kvurcU2J3dFzwjvwM14frZjnfqgVZgy500B1Ne
VyjXILVsmVNSiGkq1aUkPzQVgH7YbuBFU2sgjOINDj6X0Yz8XI5Vr7HZVtFt
o6xgKEaO31a/yl8HoSs/YaixogiPEhj6tuU75zK5+wPtegnLJfs2nieOgdB5
tPLRUvjElVJITde5tlV9LQ9laBEM+MKJT4XCHAbYPXNpyKL9KscBY0JaDI2p
sO5yewzynwFjdLp7qYM18ltoYGuxtibCNy8RUy243JZ9ELUNDyZoSShyd9mB
o1rW3i4509kxNI1ugCEZxgYbligq+ZKCZXjUZN0v7/YARAIUm92MjJZCrKq4
MvqZbpaHiHDt7R9I/5DduimbAnVpDqrGRSz4XtP1eV8alBr1YjCK2v8omya8
apCXgbK+0wgivjZfNmTkt+tBk4K5l/qecNjDIaP55CU/JDc3euvksiGCuTOb
79edA2Y5WsqG6lt2GIA1LjRnDmHQlQehbkrrUDHxSaGWZ4mEOyPizt3Mpx5U
WJVgLXe8PkeGuOhW2nifJQNUVSspKheI3ytmxRIzRBOvRs1O5GWcGQxomYcx
HLmQJwDQFTvseCOtyihxYHAhuXioZf1WaIvN98i/ZsYgSHUSutZXCvWgBAeo
BZ1VE68LfiKdbgdKzjpLeYnF3FJvVGQMFpUbJRsznyNM+XO2nPLJbxu3DGa2
SwjyR2PtLXOXxhqfMafPD0hMMQfpBFQBbd8DYZkpXy250tkwQp7NrX+QImOa
30Xst026+zUryIKuq3bc6VO4pz+qq+noFDGHf9ItYWfVvPj5yH3rlMKhQ4hT
07H31us0GbAOLZjx4yBEPEJknXav48QsCcY3rilZZoBMg7oLF0toVJSYDTym
0Go0yL8v9+n14lLGqH+6IRcCHeUlvFFPHjVpOQTUe3o3JzPtSRj3Tf+8YZyA
RxkMXtFYOTvZ8uKqc6Y8ePWLI12OJ0fydkoxlES44K5S8UCw0YXAPyUujGyy
4nfTjoY4tVU9jr67WiqNkyy1hIpBIylYgVy2Sq2uE7Kxi8Y0ezulzRfrCaR/
UOV4+bcr2P+g1snbZklf0gyCvs6B6IViOJnmYZvSDqv/klHAoOG5DIXEFnoS
YRNyGC9AaEccqQ3Qtg2lcGdFNcaA94Dh+Z5zjYle2ykiCE6sTGzXidpPDQJj
aRPg4amN9DjsTgv2vdKItxFiqrmthlNlkxfy4umN9TtjbX5FUPrOidcqcrzD
yx9E3i9LhPLKzYu/i+c27gHcK3QxVROTj3jSZdXiAB1X9MciHxv54E4JZhmW
IBQKwf4s6M4fzWrvMRbwaKfw5JeSOKthx40m2+B+NXyGsRHLqyxoqDX3Qhj4
OjXBoVPGReRS5a39wW/vxKd+zzmmSN4paiOh6IztbW2NLu4XAKBfUGiWE+3R
zu28SzZ+Tsb73qCbBfKfuY/xYbFTqSVodqfUeuxzPhAHs1iFL0jY+bgochqu
cNSobn+00Ee7Lp1tiEd6s8RN6AC6jpcXoaPTxmAo8PRX3GKydKpNvULO1/LZ
CzidRWoocjrWtYKCwkidlQv3J5JDfwe0cBDIEoVWxiR89rdWdX1e8MBnDX2r
DWaRE4iGIoRh8wNxPhYnpK3J9+B2p6qqSn2lpxVgoXfNkkjEQuNYQ/kZxmYm
PrAHv4iDiKBMfkDOi4aB4N7KHXdYMQ0bnyDkMPGFMikNI12PKKTpVav1mQYl
uEUgmUq1y8E1NiVj5+6aVYvNiVSDxJnyUu0/IaPAr3efXkPQ8HmADH0HKb49
guUoSArk+LbnA2zcHeG9Z+/MMerOpivYrGMAaH/3udcxp1adWmJIlCPXtKvn
zrLa8gsiy24rjXjUYTcaIRJ8qay4HGQdyDIkqSLCJTK/gDS/TOt4OI/OD63E
u0RKlSe7TE+OlMpnAaD/yHca5CobIln4eDwE8OvcgtNWmLbYrOHrQgFz/iQn
S8dyET7ovTSRSkMONys9gCr/d1yo1Or2ND7pzfGKz6H9vpgPnCXFaRNZVB31
qsYAIsdLH5NiwVG98lLdBpq/ZgxT+CPcbDBSDoCeFBwdqXr+fh5LUp8AsjiV
RAWhYODJUmaCTlwYxPV8jUkY57ZwUnkkWe+NOeFKHzdPLryeBLOMWDFRqEw5
JTcBIsvCg4TRDzYB+zcbsMrRMiyHcnakpH6z6L04R+1R3uoToGzq9yCcHqoW
GeteAI29gBGWa710ymny21qM7/f1XBvJoQoL+lRkaDD265/qLpCIAsGiUXzx
h3QACP9/VRr0N/UAZrODOhenA0eWBXsOSZJ9WVZfaSDOAaXYTGQiIQ8YXh+f
FecKQj16r5SPYqIdLzdMv1Y/+iq1md1UoBMm0W1E0Gl0DKoKDnu1pxoqvwTX
lqfssyNzThAg7smLvB0RnvIkTQ+yIoYw3edB8yNSmhEwvEwFfH0QFmtMhurX
Layyz/teTWt9V0K6OwJ6TO5TGfYQZnRn07x7NEkfPXo0wnnz3yOx35ndRp9m
AMO34Ab+Ic9fPyNknWWGz+kT7LicsCnPGzFAGeOYYJGUpX2/F39TYYpY6QgS
e5fjbJDyvWLrOa9vkOg2k41u2OVXCkRydDKQREERgdAAiR3sqvRfzMfLREq2
NeJtZ50O9B94sJCFb/CAJnKO8VWT1pAYOCrGX3neAu6H/ez1miQ2F958PcjK
VTsF31o5rVJ/gJ14VjT+bOswGipWENaitcc0Hqv0b/wOojAbKB2JBZ+p9UVT
U9nZtGGuKKlKSAYip+AtcWkwh2SJe7Bpqv6da+JsH7efp2n+dhR/DL/gAxiU
WNuhr9lGNI6NO6bBkaVTy0zZIsPOKVFw45YpjL6A3W0dwdxJUukHYyNHN2sg
+DN0MfvpOBDisqeciB56ZoA5Jc/+i4299zqVlmSRwPJQO1g1OI22usONihb9
uEjcuJqAnbsKVcZQmqylU+TsBBkXMOcP6xJfW26+/93QMfi0jOEUKP+9aSIV
2WD519eeiZdPmQ3eEc4F6v3Bv2QclAS1ATvQgaWfdXW1DzKb1/W9EurmX/6+
grgHLSmCmZa82T1U8kBABXyX7SzlRgfwsC5xYys0vtbluaDlezGXFOEee/K0
DlLtKuZgShzxM74SHu+DnaIpqceCRVmcRLyxSfFw+AtB56Ca3aMTqoQy0MIZ
wce9di0828brrsHFr8P6C7jeL7gnMbc3qjSrlmFKoMm8D0wOt6Yflli18Mx9
OlNZ/1djFDU0l6P2LMkv+KMD6zr5iTCEc/GGzwRRTHAVWDTsgFZBCFSg4pGg
ODwep5IQ2TUws9M9jkvDLO2rsuesaAzL2YgzB3z6W2awfrk6EjayP/9gGXh6
AIaP1vAl8IssAybjI0zo4+CR46FzrUCztdyliO79Gb5yCEeSdEJTQBvLo2q/
Bfyv1sjlCFx/ywK4jARbArHRiMRgRhoRAosf8PY5GAfYc1S4lMPBJ+i5BNyI
/HQ4QtOm29p/V4awQZkkpTZjQRZz5oLM2CpFyt+qmRQ9UG9TDouTntupkSy8
D/tpIVQzfhNhPXNzJTCxoFmuZApgJo/QP9cf4WVFW5MbYFrYvUG499V5T9ch
eO9lRQXil83HSMoPvFSirQeEbHW3SqrIWanPGRdSEb/GdzQUL8lZRYwSFu3H
bz5UrzyRf6ML172tEC32r17wtEwLBBYdqNmWIqxSz+UebKcJgVUFTejwdmXR
YiGs7Ow9F7aa93ryLhcxT6zwAtyamHD0JQsDSGrplyx2bTWLu8pjzAe7Q+Eo
XNEpj9smgNbhZFP+NLhWDgLhqF2Hzu8d8GofGOg9hUdhTr3I/9pVKyy/zUjr
r5mpYxgU+SX2sHB5i8SVx8bFj3vJTBE1Oj21YgoIdJOhcqvVA6J7VQHdVzH7
LOs1zjzR7LOKBgpmx2gI//nyO0tMugV3GxolSyqxGK62OjYfM+ugEaqbEUPq
V7f6HJVquLC1Pkcomue0uL47WmK5IIUr8Mt8UUBXvhg7PBCtwqQL6Zf2wbxH
bYHhqF+3Ff0+IV9zcgQ+cpkwUvmOrC7eHQTvAhHfWSX66cXliXsT+a/f8GWT
qcVMyJcQw+mnGwnuPn9rSfYA5mUJtiebundNmBgmS98+uAV/KwXGcU/ulj1R
abQIZTwn+5QTFdzhkiOv4cdYt2G/fMxV0M1tpT4z+XJEesUxTlN+Adv42Z7k
AJRnNwWF12jBDgTwvBTGflkeQRxPPzE6GXfcVsUQMQatAs9l++2pr+gIivl3
KlxpCPBAR8E4UKoccWDuqsiYYWo20KV5s9xCs754OkuX0C8sZmDDXOQ3vE3+
j2Ui80uv93Syx0mYmgLuf0l8y2Nx0mZiRuiSz5BKye6rUuo1tSJJxY6kqGHE
6j8LdZSKpMvJyl4uA5Gu5E3XInPZL/b1lNHsD5fpglaekLdp04X/f8qUnBrJ
QrdXdofCEfQ8S6cj2cTzmUPwea4UE9wvvFdxDzurHvAVawFFgxjZDjFKqBNm
xFsiJeILGUe73MGgLLQRiAp94lkla6sW8lpMwJmJGHlI5hYi41E/y7b150xX
BcmKBpRHyHKGde0zh03D3zkMuNca9ORY8WvYRWmwbrq8rmENzf+XzAKEN9Fs
Rxu98jhtb0cayPzMCckYd41JoTtomPZZyEOzCgM6OkiBI9/58bXyyoFApBdP
wJ3+uajhzvzJp0BobkIs/GBblQPU5NlfNN2j5FTpx2fEOXcIIE0/VzNTfkI7
JE3onMhHjDzQysQ4r8iD9n1W/7wO3kLFQGKrrjZMzkHI4RZv1SAzO67OisaS
jIRE76gk6JljhFxyDUh0DnjRysMTRKEDTZqbG3lTiYIMhasVj5AhKRg2RUgT
hFlxrRNcM/HGDcqNbtWKod8Yfd62tXsOZUKBwEyGLyW8KN9lG5HFAhZhXH2Z
rsaFZuqUeFObX0mgmZtoFwA/xsZ6V8hnuyxbWzFkFXChbxY2btdkRcqYLvyi
ZF5XILyg25A1L0E17w5VLed/+HC/hLjS/jWAN6+Qd02tBDnazwGKYNa5e/Rk
SC/DLABQ8ZIli95Hs84Tx0BuM+5KvOlYLE+ZcpyXZUShlnJU01fgO3CSJX1o
fzu8YKtyU/PmF2POSh+vjQzWDfckpXCxd29+OX9wqWTB5OQ3pE2Q+if6RKDp
Y+Ebd34ItpDyovxKr12zE1qc6v2Yp9SbZeoN8F09oMvZjIb7YD9Bp9oxZSAQ
KISTRm3qbRPZxoQN1gvu4r+Hw/H93tFzTy2OdGwB2qM9InO3r5pYHgGoeERA
MkUiaXtAmUEFxjd08c2MF9lapnn+FRiPBD9g55yrQdrVBryY1tJHTsVK64y+
EHNcyjgD60afRxCsaVzdhm/ELJFcE1NWX6X75g7wr7uohyeGGRdDMblaJNty
R0ABt6fBfQMUBsvUN1AxO4ykGLevNsVS/2sdmUb0wBDe/WkkLgsjhnWwnOnn
BcjWNaLH+iMxT+6CTJUhOZg7qnrJWH7Tx4XSvCg3Fjms7W1SKi9OVGQGBxjQ
tt5HFuzAWrCvB2L/LHrRiY4o5zUFz05nuDJHxiJ/RRn6J2rzbekhoR5Q4zrv
4UhAfVE7GUHabDYssOy+khVIRXW/ilm4ntjrdbhPDnXaJWLz1ycXWlqvEhq+
PIyA7VtckysTZX3P5Iq6h64AmTL/FBsm7hSHLEhbM48e+zpeVZaRMxzDxaPl
kotwsMS6byJ38x7uTQJcNEo3rv0C9S7j2xpngaEun3qeqTtpaAS8b9gbJeYy
Sq9vfOkmsVFHkKiD4E1NwzgBmEiXaqdauadUSU5wD6zykd7vJv6ffNEHtK5f
VK0tbmEKNrA6zAp52FPBF7551AfzIq/BJxo09VnB1VpyfresmHfI1ZxYUjwj
x4bRUH7UkHbPitI6IcFQEluH1oHlgjUNg/tlyKHjzyWrsFbN5PG1t0NE0nfd
OHpJGq9xJcF3KKYl8ChBBJAYfKSYhTSNvXXbQsqHTIMCuj7w5g7s5HA+6QYl
9ZixX6fbNeHH5ixX2FE28pZjXNTmMuAZM/LLghFhviB6dgt2PrnD36WuzM8V
B/iQ99GUL7tjqRTI7OV/+aUkBp0/YcwNZoTmbbs3w+gck0tNUHtgzng9VVCo
edX5i7+boOupBYGdGiulU5w7C5KOjmq+rOzxKFseoCrXWMhvjKwGAFFq4AkM
w3px/8KYCXduHV5FMBd2uYbqRpxNvuQIZA+JPqd+Poycg10otfpnpCZKCbKW
x9IOz7r8alYT8ed3ACcjq2yOkwEIo+Icw3YSMENyiaIM+o55eAnz0GybAMgB
Wm6kcnHkMUW6PzqK48kH0y8vFOn4Ytk3DLA0yxDPGGyxb2ddMMSN4sXidGjl
D1kKQdBEuafLva7T3TfoEQEltUHNtJf2ubHvj91981nUbbWpNtmunAAHdSJt
LNgsgDwVPwcpUg6VHdA2W18YKDPqfWZREFnICQIHa5xEmkFaoOytDHAk8RMg
+xXZasN4m4BGcofIA64ST4NdavuyO1mD2K4GNK5tie6uTW/ysB8ck5RLZ2Hb
wpU6WM2U3e5j76V6a8Nu2RfaLFwK3+U8hhONzafZ4Honz+3etp5BxNcqPw75
hNErqviaCidXrlxwNuLhysQJX73N24w8dP0eu8JSmnQSBSVrQxH2WmI6xdok
OrEHWFZ2/gi8TURnqkjO5/RIC2FkZ87jWnmVWzYTtB4bcSc+bEj9ObKndsCQ
vLQXD4rSOpijVi8H/QaZJQiJGb6pd3RuEGSL5r1W/ZLXQDDz779VHoCNNAsd
n4/m48fDPv+htE3v6HuJW2sBwzajGA+C2mmkuHcsfSCl5vXZRuRJABdhiyu/
1QjzliLA10k9T9IhJLJuHuSWQdG+mGX5p/FDDWjD9OXp2pHMrXKAslVxQdy9
XHWdsDjhr28LLehzW9IvQGpQOqQ7LdHokf+UVfOYYoE5SX4TPC45ctxbSHF5
/B9uvcWr5kC65x+gPUEm9j6ZmUqdA4i8i0Rp1sAyg8y13Qtn4MWc8cgK6Hrf
g7WB197fzni/Fur6I+b478ZNddvS11kmnElnBtICA0XvolhFP1BIEsw/jmxb
+XUpzZH3dmd1pSkhz5cZwPEryet05HR3aOMZ9N5w46cmWlWT5xz2LZ/X1Cpi
CYJri2k+0Ww34Q6+he0IfETb3QTAATGVEkBOi8Nf0vcqPIYmTEYhWH0hhkc7
Ugm6JlEtdf7xY9GXtqtA9MEf+3/i7M+DQQzoVHLCrDfpoHMrnQjhwmnBA73a
28Zi85gjl19K131FZ9r/wjKwIVH/qtZ4suRYEBLqFD9+3LJiHms77h0+s/tN
zMioXuoXcVnPa0ZIjn0Xrnvhskp3DV0zGKqFr5JvHCL9tQWSc5Io+H6xXBC1
yGhp9UOpNpMFh1301S+iVUXPqbxO0dMmA3cAesowzBPhlQHLcCGsRDiD10cM
/5LfbLOEyyqvFS8N4kkfLoWygt3s20wBJq5wzch9ktpxYgSfoWiyJgaobUOK
eLjEKnYxw8AFQCIABnrk+AQXiO0zrpSqa9Yj433HAF6EcaqWKI+hxniHe3W6
m5rdoaa9hA1SUvD5wUv4GxuwGRjSdXrkWSpHtHrHTnTblwsM9yFaAeN7EU45
McIrAFZ3tcx3wUKaZuHAexdN4EQs+U5W/dz+QgI+IeNyXIq/64TseS0OYac/
d1QAedQoRY6UN37ZgvuUVCOUY8UNC7Ll5EAlYev0yIbjrNbU2DBVE300YnML
8OBdAMoa8xNoqQgd+Awj3u9jvENROUh8a+7Eor5zaEj9+aWZ/4zxXNQcab/1
WbR2pAleLfG7qBE3qq3j/yfTjxcfdPv+eliphS5QnHi3ZRLLFnG8vUPEa5UV
YbS1yApvNUKpIum3zK8AXIwjVKRy9cRh8N0Y+MNPjJ//1m8swRzABlBcbgsz
Yd1c+Z2eNAW0yVXB0jk/0EEGg/jddjcONOJ8ICOUf4Dicq28jshm8v+3T1pN
sofYCPOFUwplrmDxI7VkXNt4Es6+Wu1dCWb8h71zTH2l0mzIqOWOAI5Hq1Qe
JTdmQMANxhzl8VGLLLA9YjwnckGGB7jJj18ESqrL5mDMYCzVvbyLKvlzFdwC
9pKD3i/mEDlb/F5xkQhpFkhHdt3rG/pQjoTBHbdHnkj/02On8UdLsI42UR2C
MesBTxRDew908FiY3CN7S9HgEp9ImzbYJJg6AeCv0MA7CI2/RZKK5eiH9BOW
iWmP9M0g5KLwaVKjmSQ4dQnVAoNfp5KMDQSVnEMSqaFUaYgVSlRj6MEyk+ym
FEZfiPHfTehjSYhR1XoHRM9yz5BCEEi6qiGb3qoBXYld2lpKZCqhot6KGhlM
5bT2mVYJotcPIyOEiJ6bQSbbRT7u/3WOsILUhUrAILrYcUQHiDCZOILWXSJf
TkUXWL9M9oQZHqZEhjydKouJOcE7Z2PAFBT3dOQeYfuBM7tNznjVzgxV1Vi+
SCcHaVjOsWerStBig7XzSKkCZq5S1A6KU6S5pQbKHmajDB7jVu/mgX4D+f0R
pklInp1l+ZF3tr6H6MeR+oCAbGjC8bEyn0hcWmolShCeYswoNb3IeHZxL/Ym
4nKRn05yx3dPxNZgub610Eedfgo0Euf4X5nk7I3rK8ygetSi5h0ASj0jaKN6
uaKW9kbHUmghyRKxB4IpOI//xTI4Iyxy+9+EgIdkEvYkrCYksk5Dt3cB9lE3
yrlSaui5SEK8tcm8VXTPEgeiMa4WwTilRAgMbZIPtQjGWbIbXrmESZbthTRV
ZzpEGoHB8Vh5iz8+gDeEq+2Rfm4mmkGlOdiYwE/RqQCLROXuWX3Ngl7owAhy
QkMlbP9YEX7yMeGTzq1V7ZkB0IwHukaA4cNG2lEyDkfR1syQuzhbvBXl2uP/
Eg3eJvnYCr4gPVH5vmDEru+UUvO2WjM+006bQxZdp1M/l76FLLhuypNJaMRs
tvkPa4xOPSs/OnwN8OhpR2P+1sZRizrUwiwasr2AsQIxYw4dhOUMeXXD7FD2
B861MUMgk+pC+AgKdSwXJoytRBsqGhbR5N/fBDEhp3oPuGSRVMzMF+vAyk5t
RpCv0CJV0VUgl5Y3K7tEpmTEQzVQywk87jyC51z0cv6+Ftx5AXFwblRb7as0
FshAm2fGa4biNarUQKlftFXTLw2nclJ08hNchpbaa89SeYYxdJ5W3/+kZ6Kf
owJ0jXRc59uCtuzj7bwEeaGMxhwZUcjWiO7LSzfeqXr0Abb8aV+zwEwOUJZ2
M30A26sb4xBN06ErY+zfALDakS5tZjv91uf3EDsEpWVekdsH4jzHZAvSJeaE
PBeckA8fvb12AmBTyrqi6op+Lvqj26MwiEaP7KYwtsiJI0ULBb7d1mqGjY0R
aKD8f4ntva7Pu50kg4RbhJVfEH5TRGzq/D213obMyl6q5eq2znghJJhWFtS3
HAwvje8QOGYwsOraDAhOrAuPM/ZLe8L7hJqCPFWvavrYJ3e/MYmuE1aGlimU
Cb65a1dhoS8drrKy7fPsd4T2fHbObNQm5+4RDSpzDjrxKSjmC+LFBmi0uUTH
zrvnT0ejrCceAYBxB0b0lqSFXKcHF4StJsO1U6w2V2UrFG6uevMS/9q4ZXjx
02lHfMVT6MUlZAJFPXWFm2hrXjLweaD63xXRAp57PEJVThfGEVxA7w2HnDo1
Nwj3Ms6nWfAc9nBZwhYFUrtzcjnug5Q75QpUeyL/04yDnLQXW+2Qgb3ni94L
JQVwBe3onXDpiytM/9td9cD7PI23tpWeQPteZHQRaFfCdLTAnB32LqIYnjln
0zl7paQHkKP1chjb9ho41DrqB1jIbvdS3x2ZoIyPMsfW5kHNuaUlbESq3BqF
Sn6BqEwjZpDeiIuK/SQjB8cNffm+ioS/+FkYDE11qL6n7I5XhmUU+iBsl135
R58QRRr04qOovU5D2Nn7FBfPu5E1tbHGstFToKFF8yOYHawrvyEHH9pJOVSN
AdsrCB0/yFMOOyN/uf5XzLD+XbaVfuP3uLFCR9uOg8105CYSUga2XulJ1NAp
Y3TDnVj6c0nd4cQZLStJ+T80Byie2Qu9Il41+yX4SkpU7eHEdA2ZnavB5YIw
Us3hVU21YU2ts+SDrTVnUDDeBrL5HHWBMe+6vVwr+Fqjav7Gpk3adWkI6I1p
UgP/vbNphiz0hi4VlR2STupopMsglveBw91TW/731nxhpISmlJjjtHjoXsOW
eME90fVejJVLqOwA5TNLmOEiG+SMTKy9ZtBVQg2K5iVYiqZpiKcU1mv98YGt
voellf4wIBw4IKFCrf8BnOAnnVgNglSLpSgAnqKDCwIrYJ9wUAKi+EfoK/6E
YOAjDmsARgxj7o0BEwnPLlq4VzBQepQXPvRKWDXUY3tvWZRwOa4SCxvPh5tX
up4Tq20HXynwUVzQxqrHWumXtZGBeIEELCvSaCYWmUwdp/vYYgkxzvYAjvDB
24995nIP+4YeKgCCzXtCuGXMtHIfN7kD9tFiHyoF2caG8tnMJEWv5yal6LTf
YRln5M6BZ4yIylAcK+lci397slC1DzDJo4WALWMKAhyXP+V3pZJ3IBfkPTH0
M6QonlGZ2KUNCwvQdThDClI+hPZ2nqKi6+GTROwuhY04flpmJzshT8Xl8UZK
ep3F1wZKDSnVPKmCIGMiKfi9CABY8DPiVuyiJpXlgzMaozqXKxkXrMOnn7MF
0MJ9rj8HDxdRbOq3xA+YZm9ST0dWlF7+4F5MbzVBute/14xpVJhtYCExupAg
EeK+YvCmQUWZDydYEeb4KEOLvtMlozFgmHPcxK6YnCG9OVQ7VikWLFMySqK/
Ozsq4VJgiHcf7kjTth2yTIncQRxaPTdQQdQOi7smqEVwNeNp1ncqdQW5Z1qm
hafxcSYAlF7nflj7vzkdX2XNXOhEqT+Y9pVIHhE/vYnHNGqSe95m04cVopE4
vVXM4YkSrTLUamdxMmlBmdesA795+AvJg41pLXNsHsYa8kNzNK3rl0u0MVjE
5WU74x0VkLdWTw7JZNJIhhOuy2TZgfRJAJ0PnKErglFxdqkcOs6eQeYPCGfy
+wh+zG9a9JtCBEHOIhFqbZpk9H1iv71e1hIi7omiv5PPFBqnxkLjZbw3X3hD
0wOXuVJo+qcJ1uLkfZDIWIJnGVmIoqH29poYyIjx6AADGs/XNSTsJpL6bvVj
1/sOAgKwFjMhnTyUg/mLbnIdrFHK9CTB4NdoLnhG5vTQ2JQpjZ8JYbAVIiqV
8tWs6J9ohn+1c+F/bkoXiFMbCRk+MEWU2001yiUluwSRRk83QQ7wOyQYRanV
eABTFGBhJ5Rno/hiV2B+DKG0DJCbWO7wCPRYTAFsLslq8t6Pw2XZfK0aBBjJ
ba1QCQJXM/V2c0xn4J9+l42wle+rXm0MKn+dE2eIX/D57nLR5Tl4fSbHdmFW
blb2jR7t6dIhBOZqgFNTQx+tQCZWJB8Vv9qJVIso/YsEiyLvrUUolJ6Xs1Us
WAZG7XiBgPtjYfd2+vubY6Z7Ut6LYpPn8wCOpkj7asjW3DcPHE1AXd52Al/X
nTnezv5VJX2rI5307v5GCh1ew1XR3XKGW/xLBjsz8icekRbk3apw3ryyNFC2
8yuM3RAJHUamqQ1n1O4I/p2/NJOanuX7/GhQ2kFn5HANl+XbLJBcGtC5cNx6
ah34PUNrpCiCdTznrA0XMWts10rkpMY8imeKxl6wSp+IuRGrP3DV0ZlJtDlf
9CxO4cxJ1OMTXeLioJ7tncU7PI8eZMbNaqWNkLX51Cn7dQ6p1gzB33PLuRvv
9t/d3A1DpddQbfMzShiubMsGiWz8VP8Nmkeg79+kqIQV5XdW9s0BzLTzyhQ6
/A0a4sE5TcULsc5zZvKouCweJ7mqAaHmiWQwAwpIoFwReMe+Hp5pN/urkQoh
BP5vwkh7ggWQ8TSjYrlFqZ5+vA1SAcYv9JbMQtdbGxWbvCmZ5WO9+rWUCNEg
A5oArL863lKhEwB2+ts8csK68FwWaqpoC71aJm2pzhVZcpRsIq6ERZpOfZok
8ss9nM+kJM+NCKKFRfNK5vJk6KbeeMMdSRqFjCHNrk4nUPtmjksSPtdAT6xz
0q4WB3IoPvNQG4lBfBY5JIBMyZ3LCXONlN+HDn7My3tKFhobZyk1bqONUQ9n
j7NwgYRxPIP9kjbtpo73Qid1I+UzlilkU/4NImqBPoc7ldwHHpt4fWg8Pxzl
atwebBStCW+Tgz6UkK214w0th8PzBz6fPhInuKjQgFQf/IU+twnRLzvC8Xsx
WIQKZLUb5DYZWUXTBSmNH3WzTTrjU6JEEFzbxDGp8trMQtddjIuelMNRctEX
z1b21NPFqvL2kiJaZv+TdzwRriq6oGWdTlo+tgkl7dj9jSrwU5z7iCvpersn
SACmBfA2Z1QFW0kWhHqOWZCV4UKWs+bSq76Y5gJ4NGOje1DJkCjgaOPSn5Io
K+BwLkqWhGa0Yj+PnnsP+B/oQ93iHrEpSh0ugXbDdFysnOEAypGuLmc5kiIh
ns3PKNblBxD0Ux3ecomoY1rR2w4FzsV4VEQU4NYky4Jq5UtIaHNqvqqb5tRm
wmhvoCpMfKX/NFC8dEOtAZY7yBSN1SPbcVlSLnuFjf2TaCY47PF6Kh2Q29jw
aGPLzBeSHlGeMZWJtZQqDylo1PrN60DzHzBMmst1fvWAH2fLYqlE0vrpLjqG
5ecXvTBnGrUrxBkuVGxU2wNizEU697X+KQLzf8Uiq9ysieJ7ehyy3u8fy+pg
nKPg6vdhXaAaFKmR0l1/hMrPoX2OQIVtQE1dpkC3RQfX6G1fkdP3DYa+A5A7
9X6a4rs771UI00zGMDg7wa9jmB8I4ic4w4z5CnTdgMABjC9TRBrWHVyv7iC+
ZfF+49ENGRFQ+NISCnuHb3IcbU9axaZBodplrmY5F6xlkeFeYIbNxDbQBEe+
lu0JW9tO5bO9CZqhgVTBfq51XDWyVEOUqLQ6hbNYFU+U6QBp+XSSGVlnz4FB
p/gyHDHUiLiIJrOHnyeknznDYbCa3jWIohW00SxrmXbTQdDzwdauJ+bkhCs4
OeRm3rS2w7TTJ9FnnnLpOgJvXzOgwwFRhwZhRRYPo332ARWUVhq3mJhdDnyG
GRI7ClFRIUuPD+2WhrYyKLMjFzbPpSjO2Y6t6N/gxc0ykgZjQWLQgEh6j3fj
Z22boi60gq6SZW0LtXgslwm+ZDDzojZOEcBD7v330GCCiHuHqtm+Ajvbol0+
ELbG9qzfaMDpoBvYAvNI++b06e6N30zenyeUU9c/HfqoxG8q/jCQuUZJTJTv
lDvaxVrieoZ9AT7Q14E66JLvaAM6s6Le+8aFy48hI5Xo1+Y4ZIXPCtIit1rF
CaHOtSWeaIR7Hvsfy9MHvC5TJ91iM5HnN+/FgwyfERSvSwCsgkCSqbD10ruX
KGCp1Sj3b618nryvAQlpj1JrAjnNJvkODnJgKOnTq3YIQ9N6VRUwglYNU8jN
b1f5Aus6t4XsrtjP+ThOV+bIQRjyGfaDZSj19k0n7VAA5BERVsLaEBq6ypLA
ZvmeYWjO5OZT54QljoBv2zIZHmv64rYX7BJJcaBvxPRwP83c5BSJkrj123Dp
aREQB+7spOfZAKAikFGi2Rp4dDu/LfIaHpK/Z+G4MxmrOpHksz0JWpFt/FSA
Ppau/ekeR8zdEIAk1Wz5LqvCP8WKJblRfhT/57hO+CD1VF6nFWxQ+bJzCP1P
Bpxjc6VMPpKdRoFYeIZeWOQsztfpaMbmymsIrd+2smxEPIvMVTShLBCczYYC
XewvgqsjbhKBKw5xKlO2BR8ouFvBKp9vcdEqPixox5FLaGEuMqNNqKmnf/ld
mF991Rw6aOTQ5ENU0LwpzOZKIprf4Crj6ErjXlDzU23aWiQjJrwX7sZujZt8
tKHa4XEMdie9ZEhLtMirY5lZcFC6lrU7lSzbK1sE7Ot69P+Ql7SG6RCoopFN
/ahwPMZgtxuOIlpxN/WOOw3SGtLOn8mvlRlr9WfaWpfZTsncubVGyRetKQHP
x3DUAma2la2ancesq9wj/V2JpZMMnE0ACT90iwvntNHRDj93D07xQwmuRtrx
3gBcPOSOj5b3CvDsALgWBlDcdB6kGzdQkuEydnh3MdVVbI/DJtkZQioDTdpz
12N125wEX+MjqFr0RVszVLL8GkqPVOUixlWWF9BM7bVS2qKHQyp0ef/JXEv5
QVIAlw75pCi+QoknHfgMoCwr5aaQJOJVwvOTkhtE0sorz0TY9VxdhhaqrHWT
L1TcdkINIaM8WKH1JWPVB7uV7CuV2B4u12RNuXRuPO6lEAIhEnaWQ0TlSqIG
S0+aUxlyJwhtD3i/weVfEjS6T7ozt/V5dUmwgCTx59p/uf84rLD5OwSCnYxS
+lIL2jQhD4GuDmo0/DAQcveeEP/iot7zgwXfS0Xh+B85VphJNXr/R8WEqi0K
p6wsOhzwEOKF8XItwi/shx8Bg61k7qtNZpDthW8s/7G03gOJ72n1Obex86jQ
lFatLIuZUQtc7z85PojFkVwt8lygA1HxqUMmNdJhqbGPNC1oZNe1bXiKL4+H
I/2kxWP4qckLlqGB/WsVx0uESmsLcfQpdh8AIx3VkOldkHtMneksOBwGcr5U
uoJKcxwv20243mFjiv+uVZ+xwPCdCNbKM/rD2qUNdbra8yClF0jw1ngJjdWc
OYTWwDgoyl7JjPT77qfVzyQKKI9uF+Mms2DTjA1ijf5zRKq6JxytPpqqhMEt
5xCmrEIj/NZYqB7r5vuuXvtKZt0hVcdKXweGG4txhImC9ANWZq89StzwkmiP
C0QT4fpSupc0WyxNFD2Pwq60vH082eGt744R4ep6t9VE7l4NTWrlZBv8psej
v9aLDDALEBq3Hqxpe9reDxIEu5bYwsToX7+2ev7BTQRekP2Ov0ee5iUIeJ7L
cuNTmQVRr9qMgsMdcvLfVyCI09mjakChvCvLQol2LPxfB2GKKcQocBI83jtS
jkApeRYDXAhYyOfFp/Mt8D2DI/BIjV2X9uf1DZmP9PXIwvwKOGHItiyyotrS
Ao4JH207ZRzeDslxEncgf2V6zNzMDE+3sn8/uFNTlxh0WdnXeJq3L7v352+s
gX4MMDoohf+2/bH6XBb6g9dpJFiidmyPg1BoSrHISpmcxu4bTug5K5GD9BkH
fN2DRGEhqv7Y2uynRN++5hisc8wTx72SNN3KycsWxFsChVcxjRLNHXwwJbSP
iM0X0I/UQvpThktbRjciSPT+lhy3yVho4XHaCKh7RJBg1/sxPTHFN5ig5XJj
W2IyYxTVaHDOxSMTu6Cg8TRGxjJ8GAK0QTpslSzQsdXoaPEOAEg7Vz0vsnvD
rBJu4MuzFnISNb/zPfFzstoRVl7W+afyzgnku6Z06/QhEu3QhQ5y4ljCKR56
OTFpteoeDS6HOz4xNfxgxItg37G5TiaAuCYWCSb1/b8OjngI0kD9YRsHOt5o
eZEu/JFsmsGZ4/35cH8Gj/ipEzhzMK80Rkjzn9FEB765gqoSsx3Nslzusi2H
j/Qbl3HCntNOlpn1hwmDyxH1DWbsb9pX2UCiKILtRw3mns1sDudfVqifApB6
uIFkF53wjTN5HP9x7p5JQMpIStVLTVBx9KujSP9JCQYHCwZDKDP95uBA6+WL
doAeLrhc3BOz7Y68Q9o7Cc4K42VWevJ4HSFlPyEp71wAmXqu15vBeymUhDoS
fnKSolowy97t7lFmM54Xf1Q1QP31v9sMUz1Tyg58S4D9COQ5H/CzES3Smm9C
+iiaAVMGyjYSwSsv45BiMrBkiI80LDe+TR3aHDexsRrqsf8kVu6UvA/osGWj
bk9pGNWmluadMpFMxgufMogSylIJIFDOuIiAS/ii3Gdg1tcVLRBg1bvYxCZd
/lCDz4MS/UXsyOzWsbb4avzfOUp59CMtc4WIZGpheJsPi6OGwGl27VqKjzER
YALZMDCiiDiQao9BdbO7NGREQ2oqPZYmPu7NBXl3gw6k9MGFbIy3A9Nd0SvB
CgU67jQTxc7NHK6jbWAqYCKecUZ59pkApggxhKH2Pe0CT+K4cF+XSleW82Lp
Kt0Udierri+SDKEFkWz3+cgDqyeNpcq6n1wl6qHwhkNVMs/1+K7JZQcWGzme
aIArfEuz2h1lUFjSYfAOfpvQsftLumUv4K9RsHxgWVBPOaLAbgI9n1z3vp2I
+xYMXCmtk9zJvQpAhKh5YTbpEc8Hiqg3bE0vopx4uNS7+gYAxcg7sr/+jskn
E7KCVujhfYF9Hjv+iUv+pi45lsJ40YoZLrgHX5GzlYl7Z0ziKo1FvF2dLyNb
HZ2hwMsIwwRS0YNvLDmAtD4Vg0kwYj38zf8SQfIMyvDKaC682kILPoVjame4
dGxrYhp/uYJOScWBrw06lMOJRsKGSnObrr2YBq+K/Ahop01lHAs+Q7vZW2bW
fxsEH10mX80xJwaCBbdqahdZoziTuXtx5dCNQBrnjGOn9dO7avfT2K5Upt68
p6d9R1NX5UXBe5xZQGMJhqSN/wJLMYpWdAvkE9SxKpSqCypji+HC0udpEult
J5+i+z7X+dzSvP/WU7rCKC1jWrMr2SWha1I6QrP6674iQWIEroT9abxTuZP7
I9DHY+RC+Wqw3A0INlcbJUS1foLjYk3dnUN/vPQBGz8CIN2w6yynpL8ldaIt
cxsU7rcOrGe0gBHGoljLDILO7ODHSVzCj/Qdlm4q2/fXJ44+hC1wwC36C7nQ
Rz4hNg3eh4EnyYQJ7FeSKY5NnqkBWxlB0R1nM8fAYEkVLcjzpYaykvn1TtMb
/x47yvLVd2eznk0PQh8Cf3FZhCCi3NHyEDT9Y0przgVzaWzBepRhCK2Kobac
1lhmmNdVzERvfsTyUwwi+ZluquIpjrvMOyTBULQcf/XLsIvYUq2qjdz1uaxX
aJNYR56VfSXboyzxjJejmmTFn7WtVtOghnRSPky7ZIJ8ydQXhJcOsUG6JATr
H6uAt6kqXF5tJ4I5i7HujrSadA/kq1DErsjV9+k6TSwPAKtTG2inrY/Ln4nO
OjPuY8dMxCs/bBRhIf/wDtS+XcM7KUpsa47Yy5nhhAddQaervtTuqYFgsyB2
gYE7gKXsQj8EUBQq66oy2fPEweD9pYyW0su0N2J7SXz+v0fEh+pX5dXlf6ct
kAB8D6mOcwK/VD+CCOHUAov99eRljvQgvYUQ4K/iUYUqhF5Jn1TvEJ28uTxR
WBz+5wh0MT52sIAuyLhSl3jz4QXIUVDoUO8Y0zlbEGEFKvk6V9WcIvxdpYeR
YQA/c445H4egdV5DflTK/MfiKpr4QRAxDkGwUtNkHY4ljAxWWpfuoHX1Donp
xt6ldAYMB8lrn4BU/svRkrjx+AUEyJ3ylt9A8g46WaOu5jWQDGMgy4rCfmJ5
42QHd68E8FZCOuRZ0jHPww57fuvzgZ2QakNFO5D2zLLI2LgmFAZRJ8ZYNmnm
4gheCiK/6rygNqcJTEloR0mTh2UuOGNFYSautejYLsuzg+HVrzEmt+WNNfta
pZk/BApA+Zv35I8Ayy4NN83otZj8dL4zrB43TYFArq6G4pi8Pd05PHYmwsxG
7EKu9uGMQ3vQzpkZY/SYIbWKZ4/xNEi0B8iAfD8Dx+pgLjeW1JJMDlHkkVqs
XCy1Hcx4BYS9wsn/fw99jwkEB6UQVX2nHMsydKN2PFaHnk5zcDQavPebMmKF
sBc0wPTY1f1q38mebqKGNxPMIFgcMjWsElUF20X04Ta1vblCTHUfGK0Ww9lm
qD8ttqt45Sv4F+x7msg0r0YhpLeyoF50UkJoyPeUPKVZIESrqgqzUywpz4Nx
eboVnzM7Bt7+M4cZUcShChBMFdqq6isCPbgGpuswV8QtMkwAga3StLRKtz0J
QbLg8PletHJwH30M3qhJCejhDZaeQOqoPtlP1hfyeD/JN+NDbd4ndocoQCFw
w229kB3EOc0nCq2c3PUnRm9sDGJzlPndSHO1oqEJtuWPKfCILYl3j/IZZD5S
1cCqmuTzIfrot34IJE8zeiqem1dVrIuWIQAhg3q2jIDQhftb2WLRzHgZovZP
H44Qu9fvALw3S2a6hZnOJjmxe6T+xUE4RQGHfK39z2TzM4PzodR6vQWsKFwC
o5eQ5ZSL5HrnODp3849NQvj1H1p3jFwA82ezTw1OvOVEj2mW9A2FRPBT8bUm
vxqLBtjTiBliB2fGSJWEh9y9+6KNHy7ctD3mWh8UocrfTGGw1YAyC7Oau5eR
iiit5I+cr1NVAuAOd6XopYVcxqPAOJFA7ngiI0GzWgt75S66zIwQxd6nMvR2
+pQ3bhUUQk0wMrbeK6ebhR6xKnE8lT3u1AGx8klF106IohE6dZMFB9hYrOXq
gwqq0A4FBGo/lUUHy25HUBmaGZ/uG49exdMY7LD/7lrWOvrfX5pE7EbvRFxL
jejsERSVuywqPWPO+rsHgu4JVCEfzyhh3P2EL09+5EPUAamsXvWy33ikvGzj
4tDDnGR8YJoKXxayYiKE90kwACZbYpWHuX8Q/QfcX8tHzFUprGlUzFPgpH4l
awzDbvR4aAp/vSsX11Oacy4oZa8NqfE2Clbh9XYkUQZ6IhHmzxpyK1P+qUzQ
mYfDLR80721HIbCTuZa9pXyD65Y1ubujIrz3Iu/VzuNpzWsWQhnBSDjbvqqC
99f0OKSweUd8q827UNU+rCJpUGEvEf83IsFnWj/n34BAlwOuZ4BiClXYB+Ce
ry9tHcXYH4AjRcmoB04FF0DuaHGgUmf0oRGt40Yl0NkZ/1rSTIsvNqWO1q/3
P7OGqmAwmrLrS4eos+Wm8MJPxT8uN7igT+M+H6ubLpVQaYqEzn0CwN1I583t
994+mMXMjnZgiyAKl7IFRkRat/4x99tWjYiQAzP/VCAIPR9VXKsoa2tcgf1b
19VSbLF23XBZk45leVKH8ErXGziBw1M9zXeLw+9drYKyk3Vrt7fwlh+t99Zw
o8G7hO7Q0VFxscRaCqOyLHLhQ5BKdXmrHBsfGW2CHF92AN2SteUz20dEXMmu
/xZNImQQlUZmH4AmhmzkNSsMOpo2jOW4akDe2AwgVex9+fr3aopYZd66x4e+
Vpoejtrw92YBuTF1t9dSt6NUjYKwNV+Ow9sWzqg5MqZeBFg3aT5j8WjZ2ED+
gEwU1vv4Km9rh/GpfiPXPM2M0D5cZhXB24an2ZuIGyUHnB0qjnvDc8GFq2VO
IQEc1x+2+AaJ3+VJDYSAlV5vMYaxIDjuHcZWtiRWpXNelUsqC0fqH9DUuEqc
xy9BZxQsn7+w8qLIUpxBOAiSMpEofbzeJKJTROpuWIrGSco3cfC5c8BAdPMV
tcO3Uk3hZ0d4Npq4rPYeoqnlL0nS8UilblZu1kgAi+YBdYIiTbtLefF1jSCA
FMHLXanL3T6HXcvWzyLkilKjGpCCko+qNR5n+LzaSj648uJIPqbXvUdUCjKf
tiuMd3QLFk7wdBd2HB2d8LHZ4Lm5LSX2oAx9lp7Lwa08wqK6NQGkgk5Cqx3j
QJzb0Yj0UUT7h1y9JnN8xwqVvpfldFrnoc/PfyxFYpvG5/iylX0zcS4RfECT
xZPzHYK9P+U1MN/f9VjAXuomYh97BXSG+XIyK2g3DzShBwOv0MjYxEEA9Yei
TY1RgnH0UFJfAbE22AN6Yom1JvTwGT4+R4mMXtkN6aV4rkTI+TRGvnbwFDV2
MtCVz+W50YzY1m4Ksw0W9HCOrxGWgLMaZte+cN9XPteiCtLbqWotMaWA7FM3
S0LBC5C6i//i/Cd83iH9tVhIzHojjXqUTIE2HgK3ZjnpgDBwoP6CToGyzq2b
IQK9E+VPjvZwsRdtT8CuC0TtZSurKDzK50Q7IC/lhAJ5hduKu155sQVXdPP3
j5jk3nJRI4+yUuVcktVb8Uhk9qgavH3DW4afBMZKXU5t3mHEz0KaXFXe6IIQ
DC/R7vDPmaGJgExOCke03pZskvarNscdjAqZlT9e10C7eaVK6EKWBPR0Mj0V
gjg2dT3qZw9Tx9xPcqN6alKtkivsq8cDhz9ry0uEkq2v8R+LzrOwIdRFHsVN
uiQPp8hAQyg/ifpk5LH7UT5a8ub4qOhPH/DpQNlhGR4ZcEo70WsWmkrZ9j5y
s9rHacCkhiggMhYE+NHuKunoPnFouiEBieanRmwSysVTetREheSQIPXe9PxD
hEUEYBCI1s9ysucStfNYmVIxQdD4GCGyU2wEQttYv2oHJ48lO6fudw97Z3zb
FNS1T11PRYgUMpY9r1KQVmZAM/DlzwAwlYjLcG1C6J92oiUZ6Zf80w2+FfPs
bb2t5SRpse2KPQpvbP9e7BUqVHQScy3ALcv+ebv4EudX0EvP4jKJHVPdjSjT
Z1IAxpBmDHSdZUs8tmBCmoy7DPcdnc2R6FdRweNMM3sxGmW7+y3R8N9wlr2s
bdAklBFrTCJRAr+Q9Z3FK7luLS3xoN+GS+E2cds1k0RuoRveP66UAQInDrF3
4+GIUdwBrNc3W+FHuqZ3qHQcwRQC6Qol7Tr220pAAH9sRi8899LsluiZfDgE
9Z05oN7zzH2t66tyx0A7IvbWjc99uAHchA35rwsWydE7361jjdqaipTWA2d4
mm6p9pF+u3L3LNxZHNqjF2m4QYmzk0/aje1InTQjtXqNt3as8VSb3+0KMuut
N42oaFGYDkFvcz9MDEvMg3ozJKVakJfIpNCp1DiiQQjxaZmsX9NlmJuYlKP2
AZNcbJHK18jpMH6rDL/8Jhfr1w5zH4eT3Bf3vNWoqrdvii3CzjEpYlUdC0BL
SrcF8ezSzAsDJXqL3CeHe4C2F+uPSKL9VE2b0xe+Yn/7a/uhnqY8mFHD3frf
5YPfC39kb+uDbnm5lNrw9exodS9OyFGYZTRjEvDrDoKMQZZxhbFAMkr09CbA
EKXWiA+DCRjExZsaS+0lF1Xm8RVcCBTncU9zDVUk1EwhbEFwBDQT327Hz8IU
jG2U/MZ2zL4k4/jGd2kC1XHsTRfulW0bIpxryGa+oG9ScCZVC9FHeK9aK+7M
KmeAIeSbiYRuAeBsJgdS1q2QYTjrR3rMRg6HQM9R8N/dKyp8WSdtW3lqlSKD
oa4NMrzu/iA1IWyk4WwSxWrJkMzHt2oxxCJkW98pn6TRKewMF55Mxwg10fxK
WeDWREKbqIlBAdeh8OUGJembii8mVZp/MhXmBzucWUE6khU0MsZFlZGLUTWN
+ZjwYNxyBZOcJmoy41+zZoEyCYATAhO7v4nlF6L5pcFiYnkwaPNAgIIq6TOH
EHQIoacviBkKk0O4uPSIxIi34RTAlGoecVBXVQnifQzl1sqac753JI55i+sv
VzjAm6JfiuyMu60Qegb1EEmd52Z/2H5osn60vPv1wkxLXHGGDwyYGZcRQPq1
nXRIkb4CZsCgenQxZUryvbzZkySa76ajBSaMJVZwohf1G5X/rCbWT+BglkUL
NB9/UW4PN/h3WUzAiaxI6Bf0ITMferLOlkI8tSMEmCmuJ0yDIYyND/ZBnJKF
z4yP+VVFiGKkXVzGJstrM+cjt4qJoOq5F0f0n8xCjHleIMhtTpeuckl6a9m5
//9HTJqwP9YrMjnksi/3rA1R75FXIWfgdVJvMZZ53/hZLwsfRORe2tZcN+Lj
kxu9TIWdQFhsRmNL1KPqtBUobnFJPF1pMg/eBOQqzLbHxfic3BcON8/8nFdk
x62srUNRKmezcJomg/Cczp2kerGyLcjixDze0vLTr9sb5kZxsMYI/p7b2QEe
mrqq+gltUFCz1uBP8PPeOX8yUXJ7lYPqcbwPa9u/qkq+4UcvKN6rghWbltaY
sC8X/f00aWRo/MBLjTJV0uPz8wCrzzWJ2PW17Fu27aHZ/liG1077da8oabDM
mVoMxXTWIXpKw9Bo/9PRA0mLfPW7TMEGMtN7U+5YIO1YYzLunfvFctDZzE2f
5nA5DDPqWCLUA3BEYnPrzDsyJiKdHJoDRSEQKVC2qPq+PojTQLNWY2YmfUGD
hbZlDhu9+ol7M5jZXK5FA84XpwQH5eSQKVeBLMHP6E6zMHK5QA83LED1fEM8
/3D2E2psHqeNfATxrcdtXJK5Gfjt8AriV+zO/BKXzYzQM5YSm9qc5vYv7X6d
3GuC1LwRnOfjVYK6+gb9PSyd2j9hH1JasC0IU2X6I1oWyL1bwbhREH5VWV71
A+OdCxUoG2mx4VXgsQlM0C3jnCfddvW05PY2T8YG0n/3Ft6X6X0Qu+IQeW4N
YufQAZGP8ABydjYc6pOQDzI9CQXPWz0Wg2I7R3f+bauP+lyPfPgVj8NZVtpq
/YkeE7FqSUrZjQAIe/7KCaks9ygQfbaNGh07VLRbTKZZtNBd/IM2oAJi2O3A
ioxSNV4oP9IQtz5FNU5I6Dse4Ywr2VeZ4L09bJtEGePEwsK6VdDamniCs5o1
UTNpYSoH+LbqK56M3yVCEqlxQnx5qHEUxfQlMXXkEZ0iI7TO3n/6xKwPoyHg
a0F2VggXkb3mdeWNtpwMhVvEyHzVmPE+2ZNdP5pM3Jt5Ejq3H4pU7Yp9ka0U
k+pDU8+CRS9qNJf9YeTNkpMTbyN5BxUfiPmajrfB9Ogquh/qPuwObllK0t+H
0sEnv3s1W+dPKhElOmDMGZtOBwimLgnH+hjugFugGBvrZTStJuKD4nApiUuB
fDmI7JqzIeGLUIHyFo7q5D+bDKtyBoTLj+gUjy5Bl9MxgAPeWX8/jVi6RkU2
j4RQSsMnOVGW9b2LhK2T5745k/2XI/VnAKB8x2ujnEWaajZ75Q4OeY4aUbe3
X8NWVl8OakI13Az5/Ze7BQYYtmQI5t/gUudBK07urYq7cF5A4kwtWkTPAnmP
r5gOnx1snSC4/kfyovAhOflqZ58xfMy+sTOlwPPow+dYVu2+ADwFi7Zc+H9M
coSUdy82Gih9IYnTUY8wup9/z6vVUBqEOxNLWrnYuK3zjP+7yBAMhGwec3Jq
/J8pE73mhxUwJAL/LsLDDa8no0z66Y0iI8Nizh6SJbfOhN2hrdmMimY7ZAP1
TLBLJehIk4yHu6paGW+tzroa03BRAgikpOMJCMXxIqewnTMDbiH5GsfWjHPO
WPYZ6HxqINnDPJSHCY7CxeJv5zPDgJW1ne1o3ymsZ3pSHkMRgTN7HMqUC//b
ppENyf3RVsKFvBKThqi1aQpZlkQS/C0lPE7p/wI34ximqkNk73NZlLGhJFQx
fi+T/IujNqP//Mm6fypKNrR3bJtmoV+jWOxqq3JWM7ZfOmW6AJcrgUso/Gmi
p6nAtEbgJQAlaE7vjRl8mUjoK3jCLNX+eSub5Tmjri69Bc6QWPGxzNdmIF4v
kzsXpxMg3i9j6VllQnet0Heei88Kc+Kpd5R7ScpAK+Damsxrb9zrm7MP6q/E
mVsw/UwxUtMAi2V192CR+b0t2X7U0KH9C8OEGPrhVWC/mXDGsbj6JA+avXab
k+5EmE9WmJJBH2n5Ay3+JNa+FnEtJZrCFdcjLYAv8VShLs5vn5tCrWYiTwxU
q9GDrgVK1U0yMwKpSxCrYukVmTdoz9rtLbVyaTwrr9O9lvbdMWuylVb2XXS+
iQNtoHdlA7npgK4Ex2bcj/2R750UxQoe4C9MSgKqKSo6qr4EGt7t0RI5ZFn0
KGQpQw4aBtI7U7ZrbRKIWfvfeXFZf5tWxjB0UIQj0WUp9tmzXHPFSl1JPBHx
DARBP6Mc+zzpIlNCp7ZDBTuzf1rua1Diqq5pwSTJR5Q/vHg5KGhHOgdk1TVs
3IzBvVN9RTWtZ97MgFACggxco9u1oaGs/tChVvVc1G+WKy25Plh5LSeMTEwN
0oUBoh9S5d7Evtzv7xzda2zrC3nc5QuwsDmZWATD0I/uNz3CHQjXeajhylon
7tFZNL93RsLVpaTZylixKRiPgiVsv8jHzDEYFWZ4dIRCv0SIrv0E6MAsSdU4
phjg4sdHyegaJgA4XIkZniasE+q1EhQfnqclFwwt0ARoPkC2JMRTvPKNK9Ri
ZQee8uOwGI88r2h/cxy4tVoRqB+CjY+enEKKh1n9QrsIcQwrLqrzIqDR6eH3
oCVnrdS2tK/qjf1PDhlosphKgFtB0tlFsrsgk7se+dgrGwntwaF8pGptaQsB
Kz41gvu0CSDl8w0DeQa8N6I4oeJsfW/FUkBV1aSAkHyP+572As76KP8N1HcD
bhtr8fC8zMYaVPjCwlgjhGjHdMRBXAGTD3NfDn0xeTdAQ2Qn9YAEzNEptJyc
6mSYoKoDwJLVEJVKLYfnqbtf57y2Ec/BmgM7EIskSAi6FNENbTbBGp/9HRir
7O3XJNR5esEPIJdWZEW4eB+Zy2Yg7muHxTP7PIZXdq1jSTU+OEwiJZFSV0ho
zdcF3msVKk2dJ0cAImtdWNaUo/sh9XrtE4ikyrLzoOXHIq6GLiY0fjBNUDIJ
aAY4mgL/hgOWbCLZCh1/dv+rtIlnRt9cyKjXq+MM1Tf93ZCt9bBOBjB5/Jie
JQDScaW2SYQnBePe4gZy6h+q6AVP2uOfUFRqr2k9OJ5DQqg1JUXJHdV56PLb
C/ROj6UwC20dq7iOWDGEJRM5cXmDRG+jFTItsEwfasyhYWRgg5nW5wSLM6Zp
j9E91nYOWHuhcrmyzou74HEXpQIvmRbhYZBNnJzAO+N2Zjb6s4M64tCvSrMT
Pkv2P80xq93oVkMrKnds8ItWMNXzdBsP8++Q0oLU6U1eJRZ3UhV8Ox4rt5KW
vV419rzj0P3s8vgN+2ur11ETuDCyZCd0Jo8ul2ThKkAeqSV9tsyWuqT/HKcq
k4gvwLB4cpdBLRowY6ANVE03v0YmEaAMCxk8Bxg4iwtTxTi6XzpnOLNQ34Os
ZqSln/KTKI8Zx5sthEuw/v43CwFzgp7X0no6aqIKaZlR/oxWRYJCNltfbneQ
iBP2UqraEbNC3zQFor5yRPukpV7yExvCIjf/LHjimYvIZwdAsngngX57nMbn
rtNK1pUgPsasnUBbDRPN8rYX6qEtOCKBspd+J4k611mGu8sDeyW1yjRv21M7
snOwrPe2dog6czi1LUBQ/f4NwvzRFV/OF/wfv1NK8c+Eb045kGKAhlvHNENr
0kuD2PnT52hCBjKK9NgYFVgdHW2rw4xrwc9SxADdcjHSmWYRx0KK9sYYAAjH
xTX3IQ5Hp/qj28FWMUPoTw6WrqIA6OvpoVyzhmImEFd0YmwCs4eFHRZLH+dq
AGomgL4PS8j0eVKQbdWL74TJ8ILL9pSM3KYcJhP7MFkml/gvPT+IUemAxUrt
5LKT+QMq7lN3J0FnxpUNFfkI3qnNVKehRv9GSTqkXe2u7fbQruaxAV9lQV/+
ZHsYdvw37mMzgjQqf3lEHkJuz16F1OWyS3/sn75sITNw0WEJa6oXCvloRTQ8
SSnLb40l/ETArOUsFPdJEVQSenB9s+s8iFfbLeoVo3DB9S4aHxVpYSeZYdSi
1ZrVA1+XR8LwL5GzhaBBJi4s+cnx5rVtg5ySxkKLmRUQO3lala5txzb07H6J
CwbLTJI33/SgyXJjAlER+rXXidtRhKWuiZM1qr4qkymnn7A9BJtoGyqe4cOi
9s5lItCEq8Qh8CVwhorY9JVm3ROdv+hkuZxJlA1DEBmtO/F9efC+WQoYndQ/
2jymDwBSr9sdJvz2tp2c5P5lWkL61Z/408aZGkqg9fY/8GOPEpQLgu6Z8apr
DKortxMts2mhWlPZpfeScKQV6RiFoGWykiyVnWJrowA/7a8DQXW7D7cYWrg+
lk029sShMh8K+3h7S0elQMUfOu4breBcMuikpiQD+Zt8YcyhVX6wjLUOmVfI
LexwC4UPglEzguy0201RDQxkiRdaxkhJuOD22IFgC0TEga3ULu8LMAruxFdL
vwOt4mrfSXXItICSzSDPyXK6DA8xOgDQXkoTe5d1No/bkaTqE3tw9XsC/IkN
OJloRaK1KfwzONNSgdsNwGrKLE5G/Bh7UQf7+vkaA8EF9xwv+q2THDQPCI5z
Rxn6jVDsPjZ7qbd+QL3k9lK1Zu72xHJ+fnhej8mPQkBCmyMTCHhgv7Mywd60
sf/ACl8ny38O1wsPp1o0tAeqeDpetnbiaEF34/hoZxQOy3UCsakg1dUJSIMH
zbTHcBWdmNMUsCVTNp/Bst8ASHDcX3B/MN8bb9u30+XuM6qsoGMGFh7+k/sf
4Jcc+b2CaYc2mURGuMkHbjWIs0WE2qh5RQS+4/YOUilhkE+x/Q0LX5Bp7yo6
ciAIxyRuwKThl6wTwH/0ozMvt2OdaXJ/SsX/EFYbhHFe4A6Uch+PGjxLbtVw
KnzY1u+LdNqdM39idF5IRjcwQdwqIjdmM6oOdeGr9uHk5bulfmtT9fTKvApj
g4WHhwWlYPZDILCpSy0RaNnmh/dEYCOCDhy9VQkviZZkO3ncOrfjIznPIFe0
OhP7kLqXo79wyZd4uslwjI9MTSr286u8JApEBQmQ4aAKasaFN9wjYSrLS54I
tflSJ/XcvRw4Pq9mLImwSJMhwwm276JWlztmSjNQ29pX5FchbbwBoClLPaTL
DXV+MK8zwi5DCwNTuNHZ/cxeBTA57Vcz2ZKu8cZGp4NTO1uvC71Kb2DY7yBB
LmChQ5xDMVRNGRd6sBS/ZMfGl3kJQhZf3F78jfcn37YE4Q6CQ3ED9Q4Ek7AL
cSXAfLhA4K4+Mg5DRH3rjuQLkmCfwDxcT+HDshmraZf5JxLzXB+vDZyCcNEj
0/25bCcuVgQ4RUJXufo56zy5MzC1pV6WMMxYXpvI3SwBhQ6kFfCVQ2JOtD0l
pR0WYgevU++PT9mTWRjPp+NygY2mut/8zMk8M48yXh6gtm6cw2Bx2RjQCLeN
E9+woYlaBCLEVvvdq4M8Sh5P+xrV6zfj/4fNIFL4UdVEfhOVBJ6OQZ4fW93H
MVcvEdsKa8kuDRLVo9wO6NjBw2fpkQOiNJCdl3tYNYsmTNqsTxuONj1fUlN4
SpM0/GMNNZAj3/qiLsR1/6BA8OLUQl47YL1OJBh+kDHvqDVYcvik5csy2qQw
UDqUcVn6LOn+Y4fOi2EE3QqzDWEc/u8wPWHjvwjLkxf5dYWaehd6WqZzxxTi
mwagV7DEGF+L60YQuTb0dQx6Cj8TngDHsd2KW9nss2UW1U82+jkwT1wAuYwJ
aZXGCRovW+sYBYIF0bhyolb8lw49mRYkUMLky5ZilqFFI/Nwb9Y3EHJ8hRtI
WNzJsw0jeL4YVunKUCVhEppNmDNGAD5Irjz/fNaGYB5gge715q1FNCKEe5+p
mMSqRifUSdxw+ObZi3rxsJAiz2zbHekSALoLnkmr/rlJcnjeh6wyrVQUsua1
BXz8FBw30z0aTSeYoCKlkWDmi6036f2IabUHiuyXh2WefoNjWACUOHE16n86
9U4rHvGcANQRrMAyQvclcWLMVwlY+hpwl4gJZDQCcUbMOMPKqu9mm2fG+mOu
J/eukhplFPoAuQiqcf0yJk+CtyoLKUu3A7YY6Zbc4bGNAeRFN+2xZXnjwjFw
/4NQHFlN4TYEgl0ttQ6+ZU4+SkwOlKAud9c+LT68NJ/PdXe++dR5UUR55hW1
HG+VY0fR9wFy6h+3twuqPA0LDpYdc8diznouGIZOF6k0svIin0Bezr0+Xhtc
0n8m8mU3tHGznG6K0uAoH3RJ/tQQIYzcAxuy+8wVh4+6QSPFIn5kU0f+/0Hd
n+FPb0q8vJY6J6MBJ/t6PbR/mLwldVf9LhLwBoBqBUHuaK/kmABpXNYpIUte
bBNVibfJB7/ydhZgS5fJzf2vnI2jSCkQiQ/OcKqW4neK+ax3XthUpIEGfurA
ng7DRExe5ttD1V7YDLdulEMZJb4ZFz8BlUhivLOzc98olzxqfXW00OtjlzCN
8aZ14sOLNAVouq1ulHYKXJY5/YfhQY9fGGzcfljwjyXGD9lK2rIyB5kcQgZ/
wxf/uA9qVJbwKf3yB/D1r5oT0bTnyB++Z1vKOUuckkPZDfPoOvwwMOhc6zUP
d0vQ2R33Y2EoXDGqYCRBFcbKrF9xxGDc3/3tRDgZqeIdkHXjFmYziUKvCsxF
VqT6D0mX8RwSQE/msutfrkf5swlU2HXdYwLMacZoHp2/GaJVswjvQE4ox7uP
kEsCLKVaJLw/LsAtrU0ZDb9qhN0kd0NtdmoZ0jGQjXJwREszY7iDZZyiMnjV
ZkUBHC15KLUqWchwXNOk01QLZImn5WVFvUFUIgK60hepwNvmSg5dwbVJUo9r
WMBjlzaNJjMJZqcAQlZH/MmKqvGtzUnLdp9jHnRNQAaU8/fSayV9bgRsM0YP
muBs2pEkdn+qZXL1XbOnVDRi0kn+BNKfmYVi1d0QD4sLQNFvLMjUmWAp4MXb
KZDxcTdEO/w+Ni3lfrx+y+aUwZ0pubDlL5aV55VnLI9wR/bI6cgSwRyrSuGF
1v4VJDtnUCfQvvSPNL+u9xCuyyTxj6NlDAZaX7xVaappguvQkz/yd0BLSdMK
p9mL43C30GeLpCq3P9wgbuNO8g170JKrKNgYqRjklb370whre1mjysy3kxh4
l8ZxG4CXk8iFIFCRZuJo5+olnW8WRUs+ukAgFAhzhFTBKyeoGdXNYMuJhKt+
QUS1kCCXYUN86s6OMFM6RTfP8NKEELxcjvK0g2N+F6UggiJl5jjQhC30X4w0
WSbY5JpXnTaddGJEue6IhNjgaaNNwXjiktcQpLGFDlpcLPewJ4lJFf9bED0w
uWKwS14/pL+GiHb+XdCGannPvCV8PtVSrKiQgHvF81uOGY2s3OmGmSCFRo55
fdkEAqqFQN6jkvB97Fyd514jVF2VUUDPvzGd3kFEJYcZncRTrvutXiKlFAqS
M+28JebonFt/GIpPidC8Chm4PnWVjxXli8lA5GyhCQytBrnJQP844Qacaj+K
mN7NzFL1yoIMrvTNQrTPuZ4JvNpXnUSvNRfrsSUGlCu76utKegbADgN7R/Pq
wAB6G523XKU8vIWVIs+oDzHIS7bQ86pv379gHUolUWnWSp08hHh0rpbvQkDP
6d3h/Zn1Sr/ys10bkD4VVgLLUcitDVeld34bsR+DtksKNq2O5V4NJxLVWUl1
6g2rHKawiAiUFWNCzjljdIgVCKF0FLqkQVpZGPhUXm8ucKKFrTTonCJZpHJn
fDOIEV3tHLoG0974ipwAJnqPzCX9M3Y4AxdS2xSU674nZe9u0fAfgZhOEd9L
CwjjI/KXpZnSWi+VVQ3zfi0BEohDQndf8Uk66QxKi9+qVZfkh9T865TNQNQG
2jVDRKNMaJ2ufAa3f7BptJAQMh5WB7QCmeZtvGDLHoDCi/qmgGBqi0My87hN
doQpaUu2Tl+GM6AZFSyKJgMAsoIsjAHSVLyCnTJnImJRKJxvVZw3qNBlE8HK
Nx5ldVBn4mik90mLwpoJCt4Kfq35X1RynubU1V+ERN4zoK9ePfj8T2A6Oczy
BiaHwRxU6Rh6BouGWbLtR6OFY3l01lzD7imiuEIXdvt2vzBOVUxyIohOcQyX
k6gLrLMH3xJ/ZkXqy2W5PeFxH77kn3/n8lHG3AieRYKYonx5dnsWgsI6P0Jf
NPQvj6gluRhWQ1LpGXguW4TPTJf6Mc7Zaq0iyAMQi//IfRo+P9Gusn7ISAVI
UdLqclQ2xlNFa8zKyqE2/yyaYvpHJrs3gDZIG9anbAwvdt8jVjwyUVwFG8qu
/ssW7qrGMyX9eCXKdIUvriZ4OpZyXQ4QE31udA6OTeZ2DNBZ6gvRWofeYXfd
+YzdGnorZXDLIm5Jqh6skirF/syRyUgqkLDebkT6L8iiXOx6zV7YwSmVmIde
8YJwNESu4MZLAt9e/5dDVh4IiwI2gai+H2lLT4tZpr6Iss1tycR0wmWdazn2
pw/bYlzAodBJVgj8QF4rzL/88xq4LVWU7VnodGVFawzwBB7xuwnKTjCKMvJw
zTQZ6W8Alz33rTLm+2WpqWsuavC209YHCV7pG2rMqAa/5ut2KO5EQRKvtYdp
7OvMGvwi693ild16UVpBrHK4ibA/aXhZZD7/blNYBDSIMpTXRURpUc7IjhV7
IPKtVdF7FK1HHitDAgkK3XgJnRfJdlrFyfZ/scMbVA7EUkfU3ymOzuNiAkop
0AyTB/DRvHf30zX2IOwtQOntj8EUDCC+4ZvsfwN6y6WZlJ8xnZTTBLnUgcZb
BJc6ZACiFyS1ccwAMhUSdvegxfgs4GcsML/E23Dz96bxMAZyjNvazTEiSiY9
/AxUQ0kEQd7E6HkRWOwd+awMkyo+7/5THFTMkQ/RqHzC2hwdAwuSLkXz2hMg
Db9VOAnc0cbmsPJtPL/nEJk2OcGGJ2/hCsm5G1B8OVk54FQcVcwyBdb9V7/5
YXHdlkHcAytNo6HnaWcyZo7TCo+6Qy8ibHqxvp8jQbVmdzgZqw1epzy9rwm6
bQ23Zfbav4p25TVIhxcbgMqcmoizhsEU1JY9oUCRxMXjIhAbbAhFhQZ0zLtQ
zBlkPKKjNlXoHIUCQyUUZoRfhEtmWFXBBvMxDT2/z9kbGp2yCSuSwFXEg6Ml
R8KZ5b7S8ibjlgPX6MIRGm6ZOxvn07iv/ZOHv4gb8fkfxH1f33FsxNwYClO4
rFnz267rsL1pv/9yzKMBCu2yN7vrhQgGMrIig+2fKbfJy12j5KZEaK5Unujm
RlLdJFSF5iDN6Yf+MqdYVApn2/4IiVXJ4Ib818DtlgprI/xceMbeo51Nk8em
AZo4YmMWuz4dxfyzwCBtzGz6Dkr1EEAjIWmU2090N29nTZ4gcP+J5YXUDmDD
0H5XL69yftJWfoGOcfxMI/zto4/zfUKhaklq3BlHAfILBQjWojRbZc4bMySh
6cJeQVllUQh8fbiGkkOri15p6oh0uS7BiFAEj0VNpwgZPyM50d1vvKDr3f0/
r9UFBwDBnlHwAibpSHG4HtCw3dglWjp1VkNTs6puEWcM5aB+jhSHlCL+/cpG
8pXWqEynXMLBcqeR7gWyxF//s88PQsx+m2ZQAcEX8jPwYSO65jYaE4ZHAIlg
ypOxWjWgVBG57n5520ERQuB1yRHmN1KLhTW40Qj3WXl74KrpMhBmKL5sBH6N
rFlfbf2hLpukI2Hagv3U53Z6YRh/UbNLJ855d5i9nN9+t5hDZGk+enUvqvjJ
m2565fYxMgrGH4Wdq62hwEY/6e04di51kAxvmAJ8xiWqAkRX9fCHKuNKVKrs
1k84HR2pUeGUpZC4BejVxiNRDNQAgBhXFWJiN1iTX7JJsmleTkrsr2QtqOKi
vlxWHKkOd8QvwA7xOaHpKFz7djOYbOOHUu/K4cbT+E94wXCsoVmKexks/cRw
O6OQ38kNCJu7DRk+S8QbP7jJy3TDD5xRlSbbklhN9vYBZTuUpM9m8DfOh6UQ
+SiCIPn2r+Qy94XgODKXdXyxIxMJxvmYOItBDpDVUSyPjmaCNU8qM+m2Ct5D
BxqNzs53y7Azi6SuwOGirrO8kcsMNtNHKjOc+Rsz5flwvUsJsmoVespr5pig
VNttlUObLeA1NgoJR0/qegDTRT2/Tld3nu9aAHROM4vZTZvltyFxnD5O2NL3
ncst0RuYdZIsDaqgMdw2D6xmjkNE2CL/tiMv+cRt8gEIRxSis3VapukzfGup
qAbOUqtaelLPZtUjwCC+R2uCm2jalXm0Mb13qyYVlzUPyB+yJt7Z2JDyfz+z
Xx/Y32iLbmDcUS3lSgoL0XQNQVX0wgsbgDws2EUZO25ICuTIcenmzJSP6cuj
AP+wbZGmHAEzDEsySz6PsDgGbActYQxgBfi/JJV4mnpXSTARCXNtLETjXi6M
ov/xXt+qYPZCC3H58S4ym9aSJQj4KMhI6BAkDFUQ5L+m/mX/ZvH2tYRp+hIc
DA4FWkPoW7WWCiRKydhnvicB5VwcJgJrlmO4CiTMZpfw4X0wwKo6GZMJ8uV3
pjK3YYaAkymVq8sCv7LbFY+BuCffhk+MsAVBhIN/32+Ygo7AD6dzWfwI6JwA
+CgQU6c0bVfCrsj/DLxYQN3TUz+fMMwCyuSeS11d0dQQxWycETRniEY+xIHE
f2QJZh+Dhi65Ek/NhNYJBj7G8MXirCh/xveIHSFurhoG0bLO7DhYcWqV8Tol
guUvcL9ZNYKmCwjco5O8LlSJY3OfC5i/BjFEr33ge7N5ws1AI9V73mpwLyuI
+gMKkykcGwqSExVajH6fk+sovWRQ7+hrtY4w98hxYeYJ69DSlfVbu7ClScuf
VSzokxsyv3cxDkVc0WF34eD08Jr5QDOYo4TdioLBJoru4mhRAGmywQSWTe8R
jbqekvY6qABBYFPGUOE3dunH/TvkrkQbDjXbjC3f3Ftn+6iXJSscsHuYNn53
n8BjXdTbfdJxq3OUFyGj086Th5Fdm6bTHNXxjGtiU+585aq40GboOnZtQ6Ok
inxV1uN6F6MTy62GzzoYfTXqT8MBGCKPrHdwu1oaxYA9n2YJ6LOpj3qfWIos
0B5h7rnwTE4jDCBuVXkaMD6z7JTKzHPfOgAza7HzNGTancSCcvlwclwVkTZT
znRls0BiXsZmQ58nmFypvkBh+qk+avXEZ2fyyytOtANxuK2K+0QbzUl4RT9E
IOTrfRqZHAwpoA9fuobk6HkwD6wkWD6lJt4QsjjRd0YcGTo6l4j4bU2BEePZ
gDYCttYsp7GQrip84hrcB4k1a34rNad2j0oC1iFkNHsSBSeF9YM416EMCiHD
UCAb6joef+g3IiDPb8JOLedPdf0nlUx8QshnTTsgz6M6KiOPRVaQVccxc9//
w7voeJEQPo76uWbF7z5CeLltQ0GjTwn3CChgFitywJ+/ZEo4tyfkpAZ+yltx
EHlBZ2uUfOAw6upchieIdR/NvhWyrY4vaikC+riF5+rOM1lBsdlfALbkG+Ql
QCCt7rU5tQ65e5J7S8KNq6kOTjP3YXxaU4Hm+/Mmdr7yjTM3qMLvl+M42yLL
7fu86/NKfAzcWN2+1qn41BArq7muZjDn1bh/8jfI6nx2gA/l76aJyDIsaL4f
J3Avm25iYrobjCTIlvip8lww056zZhddH6u3mFvieiYY7vKYQKHdR3BRpqfr
QyTz/3JhIC3O97ODUWLZw3ABf0DM/eyCT4KrYSU/JZAr46W6USkX7cfBiDTQ
bJ89Nv91AafnpjjZ+eozw7m+b/3Ifg7NE7frU6ukOXLsKFZGnk+wIAPGU8Qe
aIHaaLoVKdv89aI6/4hznF7bOr0exU80edyPsr5HlesYA/gpzyRrGA9MpO6+
0hsY00t7yWwwxLVFK5PCiyXPGGreKPMgUfo1lgV26vG8O8T3sCXNnrxlYF/F
F0Ya9qERGi95slRfPqw4yDvFKe+vgTdgrZ4b7GBQLtRv8nzXJ+05W1aaWPQ2
HaLd5qJ8HjD86Qu6sEQ7sHoO12hTNNqPkigwL+dp36si4+HvhTY7iaDEyofP
KnLhrZNIJlLK7QYoQiFhs81tJk0ZUhf/daUQ4RfpeagkwT36OX+yDzqwEcl+
I3yKI2HD8heLc78d1Vi/W6G3zLxkK4tVzdoHhRSTKmQZ94apIgVuTZgylBUe
q5OAYy47JqAL2NqozDPdz/F+pXu0k0GTIHbxunPptqtvBay/ydAiXenncvoA
2jEKVPpL0zpxKjGAa+cRGbi6O6a5DDBQMn6fauLxsSKS2A1KK/WTjarIXXhB
pLsacMM615ol3N7yMdsnpbQS1kL5VqP2pZUd8Z5Gda1U8RwUCUADyBFOrS05
Ndimyjh1VzYzpALAo11kNBLK4SL2FRAx0cLPI0BhjUjjOGKHqFJOzOs1tj8B
aQTQOd0lbJ9kNAYAnJsI15DR6detRNph3EVfV5cPFymnQGcMJwTr3eno+l9+
b/yPdby34KIqLklML6FaKdi/9cHM9jXHI6RMd3nLNZbVJLkF4HZQ81oO5j4V
KHRUaUSRDRmVSTUy9tX2E3vrk5f0u6LxP+nhELCMSMUM1M76XQvxGIUEtSFU
57g/Z24QyLdoPY1pr5IdWm6uRKbfYqHR3ok1ig2Y5arFyPHGDQP5LZ/k5xU9
RSHwDOKdVz4vkelOdrI9b9yP93HxIcTPgWbZ8OKESK4XmrKR/U47tXC+WdhX
DMKuTe/xR2IgtO9+ZUV/jIJG2PduWVqeM1mxm6d1vuA91koGhyruN+KM8s9j
0rM5fBbDO/L0xnrEdEQ0yZ8B5iC7mwbSryAF/511MMZMFvWOIrDIX+3tfAGF
gC5wKRpz626/Un+o5H8gkPD0jdWeNtnYIJnHNqElAuSYYEl4a2C1NihcnG8G
iM5UA+onoCnz3gndjHx+YbM5IN+PTlVS08n8orC+InPv+zhpdfe0iW6MxT3A
XCFiTgWwM7/t8VaRR+1tH4GTEMYjelEEhJIGH/Ftb4iTgQhG0tD+X6zmMXc8
lera3bjay0aAfIzaAq+Siow06prUyFxzw4w0p/x24eh8dQEhrflG+xgnyv5E
KHmG45JzAg8UohtOnXhZomoO0VV0y09oz7uJ+X94UUUce/NPqtrpaA2xSbxi
/hDIB2bcwqycNt5FGzDMgaKkqMnHymqqaROomkCEXgR6sZWTTUAn/5cqkSKa
ADwl/DSl45dMMuCxdiYquVVuF7+fpl75ANc7focLnhVcSzwuhPS8SzEzUxt6
i7J0rxcD7i4Dyfg5AAaIlz54nL/x5D7xeDdV9arRxMhyfZRwTOYfJj4wrbGR
4wkDWO1IHY45Z/9uNUMok5FghcvabXwLcHnb8YN+asnd+BDZ5nb9+VB1IKmX
CGVmy20NWhnonEijoK6Tx3ej3n5CeQUJTUFb0bdphL6HJja6E9V2OI1aAKmP
6ejBi/+n8gZurCQ/pM3T5yzuBoyJu9vfjWlAkn5/POEjRqN6lcRIL1HGXOxi
EKAK8eU/sRFVPt9txdTjrH0JaVLkoI7aUWpeJqSkueUCJNTHFDuqVXCRujGF
ZyorchOSDKF6ZgeQRn/OsvGfj0lIUYCSDoPtgXAqb0sxKzxcBXpZBYTdjCSf
VlgTMbJ0PYlqHGMNXmGzikEYR5qTF7LRg0/kUwJDzkuq0FFlSoF43KzPS7hH
hvZaiW9IP5g2FaqIk9WiO5mTx43WT/oteP4eE4j2R4qxU+1zRi4RIQztfu+/
nLRvt/NG5zYoFBrI3mEfeo9AQJUzgnGSzpQcNaxhVVzak1lGg6XI/cuNWdlY
6mTRu+3PIWXoNfgEBTK79XgQa+cqVuOsyEE24M9UYjDFF/2pLVltRK2BOoln
drsu88BoCJkA5sz4aa6G/jxKK5he2rOc63ZhHxXYvVbhMkka++8uKm8YToCz
0BvVddAdco93TQ4sd7GWLcbe6Ul6NqidPH+F+py3pfiDqhco8Q0EKV3gd9vI
jYzUFxDAFX33sXTIoHJiodytu6kgct6Jaqr625MRoK56oSgh86XI+GJwRfVG
rAYf85XvcT0yEzbCAe3rvSP5qqytTxKVW0EUcOYweHoIOwF3ue++O5sYQyLQ
uSEHdTwezlmiV/q160qztd8Du2w5KHMB94yglqm7JLzUoFB8i+EADc+dijzq
9QF1KGH8J60CvNCbULDdDdZWNaqZyhtt8COjlM0S+XKsiQ9DRDeKbrFkqilc
EMnHUJO+0ibvXNhmVRYT53A7k8BE7PQxP5hxifoMj7y683ZMdlimra10+hFr
UH3ghxV6NI8EhcWWuK5i3P3Pz7Ov4oDmEg4+dYZwBdnGlTuqwhdUSaO52gE8
Eg4mEMZWstIzAD6bpRv0VQVSC8SSjm/RvjJHefZYlfnM1uTDP5ZpeA1kr/yw
w2dnO32TeZrfvi0FFjH154E1s0MngmCt0ZlMVi3C4lhbH7ZR89mVCFUY1521
ltGfZVXdAZblZdEw+z8dagk4AWKRRUDewWPfKbjlAuJEApqhhe0hRcW0xK30
HWzRNr64sc59jIdGFZvVSv90kcdxHnlEh788LrV87WZbvGGe85Ko2m7cvPAy
VSoQmo8uHGFuG5+whC+4ioEnYzb8gr2RcLEK3KuKII9b/O+kYESG8+KpUyPn
Q+u2y4i6YaPymtKVzruNqVc2VRXrEBcMoeL0KvTh1XCLUl1rW0iaSAU//7FF
QITSquHzu535ErEUr50WYsEWOOxv74LJwz+tg/yOX96l1rZxLM2dHHt2PSIJ
rbQhBzCwQlLDceN+lEDjQ9F5dFtKZq/yRPqgPdxLzwn9Qaj/CqssTdu7kG0L
JI3EjqkXnMB/wSu5vsFQgeC/AXdEZXUq7xiiOKNAiz0UW14NZ8G5JJG7hUpt
kYErQ2WcyrG8Wav62obkiyV0PDfZc2hLkK5TnlF1ZK+oVyNSfG4fWFP0w6Rs
BbiXQrC9BpbpZFhwZ99TUt2E0kRw3dbRB4l8Rhg3jBZk+acDJw78Qyx8H953
Wrs092i1kS5nlhH//CLEV5cOlK3Bk0bVyMiUhmc6oW0D27j536C6Y/Qw8Q5g
SErKlB03XcAw2dSd/a5ISR68O6yNTBCmimIo4Jzimrjsqn5nfhLF65h4sJa5
m5+tR/X9Zc7vzonQcEFyPV6F91Yhm0SjRqacqVAp4nEKmKEZNMApX18lUIZD
728aOTBvRJQLTbs6JRoSjgKw/tCx7IZZxcfrgf01ILeaOPHhXmPq5U3Lf5ds
70lX56T5t6O3zHQqy1eeJXnTDrnto6xfgW5i11dZPNS8g/ALwIhvKcx0laJh
PgIi7K137MV7mItLrBmCwYRz0zoxRwRuLYFdJU6NPY0DVwIxuQYMUwSqCPv4
XeptAei39PKU4gWc1irT9ZPvG9aUDrSgwBW1kJfDEZhi18hWCDNBEkVOaI/W
R86iUzfqc8TZExUsaJVzL7sFRESdOxaO7upLXqoErvBuv2arr3AWdniKn2ib
DPZQS3bflIFaHOmEuydgj3/0bYrwb+wAE2DvO5q4F0A69DJz4GGid0EFhoxg
DoeLrMphOcUsvYpTBrOQJ9P5fMh8mM9eOi5lwUAyttZY9BogxsOO/kPXg3Jq
PGyl67RNhKVJWhsEwBFn5+SkN946koBYYZUn0Bz+jCnde1HIpHu51+89h3Dd
vToD66PZJqsSsboa8T4Aj/ZpfoVapcd4FQlcjKmcKp5rQCgbslit4MSUisZS
r/heH8nrzPh8yElh8aoWXSiIQB+YOVlcXKfi3xU+lnpoG1KN6QZoSlvQjHq4
TcBZQW5L5IyYRpXebM5qhS1w5kLJRBZbc0cl1GN8kalBnWNHLj+fhv0TgeSR
GjQZUqk+LUSxNf7Xzq/VZTlgGV+eZwQ3y9fU6kOLvTgf2qIhxQHtL/HzwsPv
YxcWSBrcwynM6zZLULvumzOEdmKvY9zbSweGCAagB6UiBWSWJ3VczXnw2vRo
qDqMlyTG+UnqPrPZJHVVzjCGuLkJwc8Mhf4GEPRVIlr75IldrP+mPeX7vzV3
W//2JzMOtqrA0hcKpxmLgbUk3EQOePxNkdqv3wDicT12LTEPJl7pcwGOe/5P
OOHgxnmwTUp+LRxLF8scJa4hBdcVw+bcVQ9uuNc4HbKbRLqyUG47dN6/5N9H
ykRSbx14d7IM4STAxRVbIe7RWJlxI0Zxm67kgIuYBUHHdww4VQqRz/+K3H1m
cL8EUDd0lMQpfXc5GenzdcZFVNWaxZvyeCoph8B+UucLp5A3a29be1FCrfxR
jyTMFmshvVG2CQpKHOf8kYL63H9WWUB6NRHBLW31d9t77n+jDA1hnrRNXh/6
l3I5RQUNx1uYMhf8zV5p2YpweST0jXm+NM/3uM8OopbwxRigMLvvBfcgobX/
fH5nJrF5k1Zs1Id4E0j6cZZiIEMO0xxa/nSVdksZaKOzPFLljwEJ6mkYX9sR
f+4x6+N4/cHmYB+tvVIQF21z8jHbecY/8rOVK1BWaUA76tOEf2UEUyAzwCkc
ABFEanQnZiNY769zLLxYjvgnRQPqCQzm7KR0luZ6e7Z4NLY8M8YEb2+Zq+n3
/Fpw89PAmxhpF5zt4qSqalInx1bkjOtaGSIJqiD1V8mvZ7qrvIP4Wv/utUm8
ZFJMDcTEPblxtKdp3Q+wiBiL8m3RDWiNwBb9UK1F3PUpZeiUvjwK271n/+tj
PiTzghxIgf6CA2hbgKr/huOX/vu+N+D2DDZ5RJTbywx5QMeg2goXsPjYP+05
k+Pq6D85iZKwQ5HSW4f1ostD3rdD9Vr3gQalAG9IO57MWt6+cVniWvn5HSIg
6X9SHNwcIG8O3pll9RVvw2vmgPW7Oh/VV0G6EZ20I5EGxEB7CsWKb5nAeWst
6PU/E6IXSpaKsJoynLRVuU4UTV/TrfaSj5yOcBwEy44NWW0p08cOUeX1pjAl
jaBtTFYsKG5v4a1Ie0xjfDDA0e7JaGjgHXzAKvSTcUrSawvarSuFE8Bvv3ZT
Z4zomRHu/z29iw+2M/Z/FlI1CG9E7H9oxBMdJxwnYbXBK1jFnwYmcGja0yRG
JU9ZSreI5+35uz1m+aF6NQtW5rkw7bbHeQ/1mtDf+cqqWxGxdFnUrc17vjr6
RcXPvLiXPcUcJrrC94v9KqW4vTQGkJ6E95+8m0Hkr6CSZv7HSM+G1D9REKDK
ztJTFk23ZZm4uO5rS52+o7Yf916+rn75qdxEnJSLWxAwVBDyC35F5X4nEbBr
hcdrpl0Xxvf2/wNIuMr6mk9ttdu4N9xfb9nLzjafp/9k0WoNwmu6lu6xRckP
n5h1vcA+WNpY6q7j8BFUjB1EYS0KHYUmJ8fioDKj3W+KYG8sXz49koxjnWV1
HLWTRwARB7ob/FPbCWQTxV10O492YK8sxysGtIyh0yhLMXXislEPVui2CAB9
OSgQudXgr+0JsJRZYUsCy5/vRVmrpYflOCc6q2QCprQ/FMy+Emv5asd7OIO3
Bw/QklEhCcpi3+suhAb3wG4qwRrYuZbMF3x56TDDfggM+QCSWAZr/pSH1LES
FsfbZLwqD0kDd2n3WjHmM5w2g7iuGG6KjpKjuosSrsP1TdQvAXionA3MXSt2
YlDzrV9FrG2jROTNZDRSW+pqcMu+EnctAGs2T69XljPJT9EoDo7BTIadkoh4
pdMYmy5m1Ey87T+QmATbmvAQFHC9KPMxGDSC7uKK7L4Rj0HBrfqcmNwK4LvJ
0bsCkWaD8Cs+lSXAPd3Qy6+Q3QDv5MqDqmj5/gTX5pRtLCWJtjsBqiXwXTH/
t1wI2X7qxsXml2bE1V6iSt48KHsP6rhMseOccU1QWk5ctM3lSx7Hic2uP1rz
KUSYXnK7MeDhBfCft9Je0xsQqV19FLzfWi9V+iF6oPEUzDjPQZevtgLfebMb
otTwt4UCQ9TLbslexB7nli/0jS37AObWSm9vZMHVaEfA3si1x35QOfbQ8Vb5
nvRDu96vi+omLl9Zw5xam5VVvh9jBcD1lmUur43mibFkcPnb0jEhlGo/cJ3a
46Nb90lkynUPyXWo9FG2aoh2/4tWuxhcxRzU4SvDUK5Eek0KIwZn4qwwWz6M
JKzg8m++E8k0RQUNwhfq5UYIGXffhXGM+b3pU+U3P6TmoA3YkCNlcVLSwcmw
cAuROYoaiSrh5kbrbMXHi27nNbg1Q2hS+Ow96UCGzXIrnYrtYpvTZ4+329IA
Em5edMvlA22KT1Icu4LYlsKoOOcIiB14mITheQScXFTMr7XYfa9pZh6uNsRh
UeWBvjOtSUK7Zs5Y1OjAhqXAtA50JHosv2NbRXovayZKiv/YQpP85JSZEL2g
MDzhWtuSDdmGDoy3pTjtCbBGSNntVCMyvacXgCXJYAQdzGBpZZtsylsM6EAw
gyDz2fFOOLL55lwjPqFZVgGRllYknRbNGXGhrRriMmx2cl2WA4iVyfpNjjZb
G6gz1nr6GXWiCLXM/taKttpzJRsxTM5Gc3xCs5VGE6+P7aJOe0FnurCHmKgo
tLgihHDNx1gQyWbtZsI1SjuKQEz7Ug+TZsff4Zio0F+7ZyCHaRPDOiLDZJKN
DuZci5NStnFo6DWLsIfAjaEJnWDoBD8kWI5nhrxQpdL9Chv/9PLdMUVBGBip
egvRKsmmOWvoW3mYlizeBGY8T5Q8I54SrEGWoRjLJSHL/Z36PY7kTds4KW3B
B1XtSX/9AlaYScv1kdVd8Yel9JI/VnVjdeBhgE3vV6A7F3zVTnMlPZO2wady
zk/SIURgpoe3tZmzon6GLCNaVbjJhjNYzgwqzICHGjzrXBw6O6fSZEV+OqkY
bcAl3MYG6VsMdsHy8E6Ar1jRl6Im9Dbampb82UVIub8ATjT2sAS2y+eTBt54
3B+zxRPHgtyjXv8oUNfty9HKVO5smxecn6TmAAr5qv6ru4soexHOjB+Zcrhh
+ynx5O3c+IpU61GllcYvKquxVtotknE21C5I0EVbDbUNUd1nGEVMehkPwZsE
UgCPY2p9fjGFh4KNT7M+NseFa7Np30Jk4Z1lvisDYTSuXzVIMi7wc0bKN/88
ENpSeQjLSbCrFjmHBnc940smvGXpXZAv9419TRoM3xgPUqwSu4pNFXpytiep
AnOZBpXShV0nnED/JnYQ/xb1fyEVbYkFX3p2Z2VhLOnq3OXRIA/9KMJuP1fB
gP++cwyq4RAIOvLWAzNIhc6/4swRcOpaM0/oNC4LtEOC0fUaR/+EqqrxZ1qO
0JR5DB1zPCjABiyd2PRoMANuS0WJ2M+rXMpa4yy4dsjHDByugroxlnUAo+q0
9JtCkD2EQm46xbc86gaixf+Yyat128fjhDYJjBrWUw/AccURd/bDBn/lU+wz
sfDY2Nn6h4x8dbosuVc+QsboIj98vWStrlPHC3bHaHFCc5r3JyqCCvwccUzr
OQIdTb10xltBeUdlhNsCRq9gkAiN+9bOJcftRpZ6jsy1PcOVwlnYj4m5yBTf
4Ff1AmMh93SOJJBTtCimuDiI1AuyO/8wS4rsOp31oFECCO434WI6zuNrKgT/
hTUXwmGQhfaZXd1srLYQGZucpJy5vPfco+agiHpY6CaaE0qCCmv+A69LChTH
Zw2+V51BPuHlsGbJa1NGpxFxUP2uSg2Z3Q6VZFNzAOUW8400q8o2L10sFs2F
1duzg/Z708Qau4ajNoPsfW2ngSkfpJocxwqKHvp3utyYLrJmmz83lgSlJlbW
d4/dGTG7i66WtYdXRJt1nHOGzni/hknSTz4KitGHipDhug42Ik5F+kyvrJ4D
JsA369lwe4ojleoJFXkxutPv407j4aBJFiKHoh8Fy2u7ZsGuZMRTA6qfLlZK
F2kCBNReXFCWFylbtLAkiAwsUnPJgHWJDK1cdIiW6R4nXIZDyTkGOliAt3KC
wi30Woz9HGRgfF7p6mo8DFb8anGxMvaX0A0NyYjR6vbqv2EQMdA9Xlm05DbK
ghHPgoXj9DeaKWutYvlJEkl58SCIYfT5EMA8+J/6wCfN7e46WVU8TyDumVRw
GUD6N14nszdt57fnUHffo+x51a8zH0zUAKZF8Dc9sH2zdUrUfNBU32JSzSW3
SZcdPmchSoK4vi5FCiHS6cEgM7sVZz0FqlkLBs7O1TOUHqthjJ3co4aXLFMW
q6opBgVH/CLnUz8cLh9Mu/FrnmFvWYIcvHECKbO3f1h0tjLf3V5TUnQApRgZ
+vSKbd7JZ+9uyZ5qFFR4LUeRK8kBGCvLpPuqPxTBXPhoGGTVqP6fjCLjrvtr
HrjsRzlGMD67SQeDPSzGiUdZu+jr8qXnPbuZAmWt1cKQYdMDj5cS+BkYB56d
9RH1eSmzFajPVcHgh+7Z0KVl1/GjGQOX4WGOG9fWF7OrTJeLVz+bKBt+dOvr
N4d3A2i96UDw2O+/GKV2FQrzbPn4TKANaY/uqFKBXG9SoGMqjw/TcVZSNgdq
8NxpUcCn7u+xUQXBs6pa+bFgyQ99G55SaCcMg3kBQG7mo9ehAeg8cvMPLn3L
6EYfyi8j92LNorTAyy5fX764BSocw/JOg0Ws427v/PNjBms+QgmhaOacK4dN
NFD0J+pedMkTopl5OZAzGCYe6aDOiGgYk7nQiioGYHSMVH1TxrrXKJ0oEhZi
YZXVWFOcUJNl638QFdt5n0MjqS+upRJUnTSwk5p32r5jH394n6J40eadz0Re
K2xuUwjwhbAZzXYd25kxyh50e5/GKawGuWp275vnIcGf8BCXmfApHL2A/Dsh
zK8BaSrHC9Sptdga9zT5wFysac/9ssRY4aqRn7MKv1fCQUDFIZPcGmFrZON5
aIncU5rmD8U5Hhw3B1wkQ1VAOFPTDQGAuuEtQVLPqwwMHomrTSmkrxsMDEs0
B/G0I9jqJrI9IP44My72h+ifVI0EoagDKAw+Inha/eosRlU4eb3vMsxb7ZDt
cXUGyuDPiZZnYZgDHqwSHbmHqDpRS25qP4M+G/HLnwuEfm21o3gVk+26MUcq
usyBzwTk9GfU3c0XGKYsbN7hYH9z0B94JK88k0TqIvWNZ2Z76HDET1eW/pGE
Pqwv7ujfZKA9zx7AK+pMiRbuqi1iXr+/sliYHcgXNKfunh8GG2nWiSmGRaUg
yaeywYekSZxtkaVbnoLScc9LpiUAYx1hJvP1UECs2bwt1lkZjcOsxQ11xBy8
g79PBGl5RTbi99lnmdO5WY1/nXx028m5yDa9aQTWHqmlJfJeLw0TXoJ+tu66
Ua1TIwyv67D4Xb3xNsiiYFiGUPYsXIS3zNg3QQ6mxLo/F9acD1XxDIqqi0Ak
cPfnQ+R4MeheYxow5ry20CjrY4PJzy6D4wg/wjeJM/kNKh75jYeUDpNku6FP
71XoFze7qgyxfiFrphjtjnPBwVJ7Fmi+vxxuzxsTBLddTIy3BAxbdwBeiAor
rgOZO+opMljbL224h3m0GOX7b6d39H9Rwce335hFsaBmbZzV0bmVPsJw1UJR
Lbus+TKMxOaCxRG30c4vHOzJmi3XG8kPgv7NlqRBwg515uQ5+K1UJo+EEPec
+sMQ+eTpQhem3+h03I2SORYCkdCpQBvmuS/OcIS+Kxij39ZIziB3zjfOPQo2
a1kbYs4Xktk+GdvllVpIlgODEQrHIJlATlrQl0FoxrEVWDFliAo+kOHdr0dd
G07WbVCz2iw06eUpdbZq9BNkeoGhplmj8sAZ5qvEExfIi9OLyItqh4LFvrri
Rj6Ju1o3DuULhsor2lYoFQRcbOui7TA97fiOIF4VRPiZlpPAKHXLCpPuAiEf
uIBqA7J3vT5OsS85anT7FJ7LAG7ErfqUBB3TezXKBgVbgCNioo+oDcCWnWr9
vtzOgOnsMUdEkj2fMVbHHn2IoQEc2UBCbJwiuTvEhxluq/zahFlWE5DcT+Z0
gfDBp9Deip1wwdYLeSvDe3/a1fv9Er+QrhFmOxs7bLA+qeeL23GrQ0Deol+N
r37q7fnPv8An4q8x79n+Nw7GPvhyUEmeJfpSfU5KvjshG3oWYLx6cDtm8pKP
mEuqLYtLNRUDNkOgANInGEUiG1+nZZ+Bs7oyCOnWZ0qAJj9skLNEOI0Hv383
MwrxWm1DnoBedr88hfiIqtBTLeAIEA6yFNFVWiXh4OcyVWhgBfFgNwBfxXFH
Mq5NswjslTvoxUZF+shJqKEX5VvToPsIXGkeh2ZDkvqP5iPWTtNl63q63pFa
jUWuma8VrWSU94ZcvR73j79dXyqF0Am100Sgw769ns5DZWFrLVr9G+Ve1WyU
O4RdrWtTRkPxTgjEBOvj5flVQh9G6/MN8EiOqJQ7KZp8POfIYQ2i+9zvecXl
3dKxgTgic/43Vder1+JCDrjj1wsfriIn0XOAxvZ4l9Qv8Rh2pI3ijJrVEt8/
VWQwPDbpZ/Jzx4OSLkSgtbvNDd+2O9UMV1j6EzQrsGoZIOnLl8S++oUSwkC/
rLUcOFasPZLHUwAh9suz4T8dgGaxEvs7VlfevQjIKvLZCu9qIv13uQ9rO04p
CNaTzgePgyWVQhsR2MRC7IH7zFhufSFwSWTWSYxwWSQvRo/PayMVOjsFSlrd
UPjbOD+sJBU5JTFYyuwFocKL0CJ9VRy8WT6dTbC8XaKo46iqiYQ8IPGsPLUX
HzMMTTGUCrpxhRYIeA15LkfK9igan+Ou9q+xSbF4cRmIhS2JfVeKk1w7lPVT
JUeim8922MY/hhuTMO/SKaU1zhrMD8kQnFkot8ib7QcEqwrwmw1ckWkzit+k
eyYChXUYdkC5RStLyqOiG/ipbcyP2oJmNU5D3RtebZwIzo9YlkkB5PV4KBzS
jfalzXoeh0zFt06XDi70mBQIrdJ3FmsWUgMv/9//hJ+0A2hk7iLjUq3o8MW6
/IHyIXsJ8VDGnzj4tHiSfDIz+r/C/vMZ5ePbAbFl7mCBpNTEmaGTUt0zxKFM
OClIh5ICxXZpCZ93OvPIKrd3gw0/m5eIIjmNgxVhNdHGekiAtAR6YH/q6fL7
fqR2GHYZi/gUr6BkFwzgm0gxuaND+DXiHgCgyHHe/39p5XYdQGFokPsv30XX
eMKzRZ1D8KjLhTE1fQHHiCPRFcLILYzVA0GwVjtuyKyfteYpES+SM7EVlODJ
ZBYl18eVloKe+yYdMDu3861x6LQ8GYN3woAQWR8391EQY5OmQ+OrpqLODhjS
OgICP+iqA279rq9+mvQRHpTFr3SN3Xlhyz+DFvZ7qBWiFP1JUjbbaCGwzjI9
2DMoNOoim59P7M0FqSVO7IWdjN5zlFWTsYEehcdPGhwgYGLz+UydQEZ0am0M
pzzGSfWs/K7XE6YuWz9W2JmwXs1BFSZY+y1HwlPnTUJdk8VQPDo76noP6/nZ
mI3EXgqWzY9Oled+r97d5HsD8dO3tSylWG/SLCzdMDrnHF8pXEJZI9IrgGnV
p09y8s6U32A9++xQSNF+ijP53Q2ry5znogXWErs8Rr2OrPyuUmS75k5nNQG/
CPKH0429HAJ/9xZHemu2oIZc2NsIiGCDdRgBuRLyli29uXv4eQv0CadjHODk
qb/u/gj/JHvh2rPyt1gcoQIEiF0T55bd19wgEb7N6e0ymcSgT0kAAmXLQEht
LiSckfWHK8lBgKluWhZqIpqb+IGx7uDrF2Ua03pZag5IZPNBBE8x5/22LG9d
Ra2DDPeKT0/sOtc0myND4z0sNH6RkVFCx8b1fwGh19Fs09B8u04S++k2Xqi7
COWrCoaVP9uNvTn8K9cZ2++wMbjcrtLVh0ZIhOAuV8BWFf5Gtssr1EKmwB73
cp0kqtUeZurS80Ilcy/DkrjN/wN4uwd/JjXqYvj8PxYvozuPMmI69/Vb8Ueh
EyamSe82b/mYa2KhQ+1dHo1H+i/0Heq6kpYKWmRGKYM5oUDBIDOT/0+3R6fC
PCgstpyJD4dZYy7Yo7tzLXu9962jZFENl93HsljGeg3KONJLVu9G2sBIzDYY
gkYU7bybcCr2Fu8EjcvTsGvQcPJutzptOVrgi4g5GxTUHsS2mMTcjJhxNB/3
sL6kF7PJmUvEf29M7mY7v1WxzKLA5/MWt0BtM0UMTnPGUrdjYzEclDO4Kby5
wbcTHn+4cTM2li3WE1WaFzt/kEgVj9khQZHmmJAZnXqoWDvmHwiOPEKTM25g
mXo1sNYkEsh6HHhYc/iHVxdeQ0NFQuHIa75hVPN5QBwPfrzzB+w6uT8lmnb6
rHjx5QF3nij6n/+XhYsShuT0ErsL0rPuochF3xQuCOLASBCA1EovIl0R/AON
Eu2lhqGTcD+jCHepPCTR/gs8ydNbXbpDprsQXqKd+0SRGhoFlK81lPWRQMME
g8idv8tIpGmOq/5nniu4mIiDwiFG6a3DMsqiLmWf36jtyk4FakcCSBgn2mND
/WxFEbHEBGGG2pmUjaPzmypEfEWq408yHIxM7tKYssYljBApUSLNPxsFDw9b
l7ZFAVsuuHX1vBCbNDEVF8bAuRiZfsJ/9hoSW3RbimGVYxVxvCyffKKqOu5F
lK41VS/8LcwaWhMyE03gQ1hWUlwNQ9bho0dCtjlPSzzS/KSlamfYvYiaZ3wU
hVBV5OpCv0PVla6J5oz2mhPWgx2GuE6LnyP2FErJCEA5zxGQHKHTKfF+xQCk
lm0qMtafgEi/af+sg2WZdq8X6Dmc9HKK37s1hRaPfd7kClxPWHM9CMaMu1qz
wvQoNFKnEUA20KQWyhcH/HDagGDz4NDAoknYrZXBu7gGpcNo8A/askj0TEd2
iIHrC1SGAJKKl5iwNkhhieBdr7PTWa3/kAU9Z1kaFKVCJkrt9gTB/FSBYcau
w77mfk+yRXK8H2lb94xy3TO8XkT/38HtXlBW8WjhAAfckZ73yQXsYStkuN7h
qy6vE54wa6xIBRBPRiFtWFyfCFJfGDoZJdNJexVhRZq9UEGLUmjG2maSRf3l
lSM02OdSgxrVVsi7OCdpLaRXBsBcKujuFz1udLSokm7ar4OjIjROpS5R4CGa
QUSBf6EgGacOB6kbY2JRc8MKjemxGoh9CVHpMiVh5nvHzgXQDztB6zklQk01
lxturWYVDueB4DhOgVE+SyR2CAF4PGCngM/4Dxk8BukTpEYpc9JBUasH3wi5
es2V6u7hszszRMZvDEHNSqcFUurQVH9F3cNSv/J0lRMwRo0A8+4Mj/rCRD3n
MhU1AEIgnbdIRsCXq6gskX1iqe0YVOleyR3I1mOrQk/LEDjg2Zrz01FD4WKx
99R4sOhg/keauZ61jMSQLpB3A5aZHYp0qMJGutt5vsmlCekaBN4ta2flwkbW
NsLFX4pEldYWfMvET0QXZi+InCoj6r6x73Pb+W6nairM1T0DhfEkTpHsm50+
1XQbSOf8UWx7fe3ZBRYTFNRKpf+jPvVVMSX7ak5IZErc9+tvJag4RqI7op+l
2JNRSFdIW/l9gBpVOPsddrBAAciHSoIQ89jRBUoaLylKlF6rfLgzc8QCMvpa
VAIQWIYkXvyxUs7+T8/fTEuhOs1j/6QIt4jtPg4aFk861WYlsYUxhH49fQat
EM6sw1oTJqJSX5pwvICyqGD6mdZqI950tq76KB6Nv4BLRoXcO8NDb8B7B361
I4EEJ57v2zBOOUw0NQ9gm+B3keYLKKdU/1uH8mbVqECgqSnufYxzKnlcrDU9
T6u3E9p1cQB5Sfe6IQySI23qBT35FWyudYWrt2aPtLKtc2JMI9oE5teTBavw
nvL+a/zKEd+G/zfgHlIaz+WBsWtUKeDIrg/waU9V3tv6MeVpwfKb49ZJX4aV
BHaB1p1DPBqJiQtfs1Ksq9MRmXZYp6FGTQbSbrg4FP9dLc6wBPyOCczhYPpp
+TEfgOsbB8qJ5YoweO/6uJ0C+JMKz50k7YnWrI+uOImp6cT9XzgjC//LB8B0
cYVLRDjFgyFuHoyUNQVpe/6kLsj5u5+o4pReP9/QTm+P+6qlC36CdhTL2BSl
2y3SZC3g6mTQauDzbMEJwRbRgx3htPCdWxbL+By+lHXJJLdOeW9I8+xJNF0r
Co99oZziCjz2UPdnUAWGYGu+R0gx/lSVOMYSabsbL63/DToFpCHzT90TO17Y
tj+1QXcpa8BLu2EEsW6AJVTeA+VFESgcWxPgMiH+cWO2DSqhsbwBAbOIQ0fJ
IRtY7LdDwrF4Sm8xbJpmPfobpicxEhkKxWW+Y1wMsU2XUfOb6bkkN3g6LZmT
DpfN0VbhdiWtGuFb45NzjwH3/EG2OeKGHKpjbe1YsN1Wo5qBHJQI2VtiiLUe
xgER39WawLDC5zFrxXdQ24VKBHKSCW68YwqSrrwiZUkEHZjoeHv3jCRoTGsx
/M4Pqxn1fIreAxpvwVPjhL0NFSDVrOwmGMsShPWxAsW46H1NukERT250jKmE
tSJYGp5uv+PFHxHMr/H9yor9XNCwKhgzfjGi6gQTQhXNsz5jqJEieQglzzV4
rhBoxOuVvegi2hAUPu+mcMNhUyJywyRQcb4yuEdaQEi1n17RWv/qvnlcey2E
IQBe1VxWhvdt7pQD9ZaSFhduq4Q9TDJP3Un6IIFDaAIqu7mH8YONmhI2VdUS
f/7ltb4jO+i/2wIspK+Wt5c6BynmUH0qbGNx/VFEbCDIJGpkrJfOrxEwwsu+
jOJqzsiMdR5RLmDSIKhYetpH6tp6RZwJiAEzRTswWhPbEL9azAPzqeJ1ZlZH
ATaMPSysY8vjivEhXtur1INzxxAD22KMt9XYT1UNsd6zNXgFBDHVbtN0xq2o
LZJoYxHZWuXxj8nlSzZzFUTS/Hj4wHzCZOjVWL0kfy+sAS6xdrsMhuHrpZ96
Npug7gjcNGZwq1jo7thmeVzCyQjJ5eLSbqx8/Ks7S8XTK0sSMGHl6HNd2pWy
Vi9ALhZTbhk8oylDKrh2W/7NJMd0hhS5x7wtegKRpy3nQoPyuGLbYjoGBLzD
oee2nb1YGSpW29mvIsjPb2o9rqpHKf/hFpLU4pKRtzdPQasXr9tH1yH/30aI
q6h/V6fXughfGDmnqNNtKQbJj3zNIGB0zwbiw0lj1C43KcVNxMO3JqhxxUIF
/5hMkNhAsaDtHO3xCNfNrwPFDAB6ah3Kyz5HRF4HGN1aOvhVVPDHGBUuJXw5
lToiQm/U06LOjGir/NYZ8JMrxI6VLVT/lkBCiGyE69MWp/pcutrmRkp0Zmup
e9yx+nJlI07HJGdyKBTyqArx2j40Dl1NKnQEg5vrmeSY0fOiswLf4K/qltBD
KvVWoP7N0HQIY1jtW5iIhaun0Qb4wl1Je6+E2qF+W408dM/uH8Y2TfvMUx8t
JbH55iwpOLQCpWAhuyyMQ0zxWqx5clAc9G/UfepuWdvEgI2dA8D7VkfIDL+S
bdBuT6c4sazH0rQEBbp6+hrm7KQgY6brN34WnYa0ASMM4Fd9QgQ9leiziD5W
9PM1kf8AN76jIlnxkG+6rmhHpI76DqiQthntEJpHuz6E6t/udgYEKBRlvNzQ
5be6N2Gw0AWXlR0uauuEgoeTmRHDzG5+syAwcSEZTm0ez8L4uB2rKxOF09pD
7dbw0oUQ83MxeHKU3dvQalhNCoAPZC2Y8pqxnIWhlPIJWFo1dONMZ6moOlKn
Ywk+QsFIGIdpXFzOSPJ5RdMonc/4bBohOT3GSb49wBbbfFqkmVk6InecIbaG
u2DXmPXAr7n64bvE5Xgrr/gxRAq7pV4HT0D13D3jEyax9LuV0d1L11FSKVRk
rLYkKPBH1DO5awTB+69TX4JVOUqF4J6b7Wv1PIolsQL+5KWsnvE/gCVEcJj/
V+XCR8M6PiCSmkGrc8WJ4cWGH0lGjPc5MX+brS+2PS9f3aFQzSOb61DpHcLJ
+mMEcpbpe+tURaxy3WesVU6Mp6aS6dJ7uxJCTDYgjkoZJZwmrKgBOx4nlP9d
EZJpOvEHe9DOVCOelphuh1W9M3hZEgl2QFOTByWe8idzO6vJwAgmbTsmy9vv
V9kRQ6M3WIi5LnAOhIb1131odvMnd6Oo0w2aLxf6pZwfjF5P+/qO7nFFAl4V
HR/mnDgmB/o7HhU4fB9gev8gKftus/ctcI/HYCFRQjI1uKVsxqOtdP5dxIOL
otirSgkL3Okb8s0ROQq0WSjCYNZJfmqPL9kSP6dBnt/tEqHAqxwZ+X60KBrP
jPjEashy6YzXHP93gcN8epRX428H3g9K9BjnZ4gRAe/Ueoym62xqgEPAgxCH
rO4nfueXGZUNPdJ0Ht786E4bPeyGwhceDOUBONufIaeySYDlmAiS2gmqnJ7k
gM9xem1rLYNw8atU0sxUjg2r1MXmhsdPrrpE0L0eHOGw0JbWnmfo7uJUGwjt
2PYcfazxhFU++NzAwUeybVjgy87TLwVgOZChuGqk4u4Uv7eUjBMVl+NsWIkZ
JPkek0v95GCsrRzwiur3flN5qkc1ibvVgeBnLp3wYpFL9v7G4WVo1SUHVoUm
i3QrKLstILDhvI9G24cmzkPj6kLU1TL3DzT06ybxi3a6taE6X0jChV1cdxOD
vtPdDRswd+Oiqk0e18OKF5aY0+ti5O4DjCtUTn+rY9vzKrnXuwibN6HEqfGd
HhlIfs1KhSWe9yPUCXiTB3iZOWhIzGNBW+CVcerQywiGw6IpJ+AAazZ4BRx7
yYzQNflT4k+yNwUhK/4+R0T6/j4hhuGhN61AXLcJ2sTWJeGBZ+YVDdM5ukxk
x+39V/isStNm2j3vQJEuqr1X6oa9jF9VeUs6ORk5RixiqJvO4H1H52CSobGn
Hiv+OzuaUAlYgsAvfCS0UXy0MhDRiLOp2p3FQ55zoLHDQZqaGhMuraVpmifH
9NJoI1tEDQ+1X0kXOmrrkFdKezMH76OheX3WMqHuSzJPUxM4XzthA2f2L5Vr
G29MRVuIFSG2G2AKzgE2M4aSGQepKUGTnzgET5cpxc2n/9IjgVXrxRP/MbaH
TXNm1tOyaz3/ZyL/xFBY9AIDVhsvxkZFnJPKru4RTOhXXs9I3MCYaVVATkk0
i/4faXa6KDpFbtougaAJCSuukZ8YDvbquY2HRrhQA1Jv+VsqWkGPZbEwMKcM
OTXl8czaPIk8nSZ9HyUOyxFBYyG/qy1vVU8FTBAwiwPoyosUXDyviL/1QlHq
+5wAqKG8oWQe73tCtRUAyzwMmAYfBT/wGb3zBUwMSTBv8TiVKedmTrP3uLY+
J26EMJ1utkA4ORpOGXNQpLiwF/WKiHUnDXBnlO0Sq8Zj9L4H1sGEvrnS1tcT
En47yw+Q1uODyHBoJO/xrNdp5oWhUo0/tNVCM3FtIb3mUhUSSUR6EpeRbaMD
cWV4wpb7Z7qjsQGxTYrnYWs3jmdyBCnw57PHb3x1/TsYfYi84ReYU46Vyop1
RVMfYI/Fz2Sn+kL1hc7IXeicsquieG/RhAbR4tf6+rPOywAizIznR1JmZa7Y
WGg/x11CkCnp0RLuoiSwsZRH/zjB3EP7SsCNMYWTWit4N+WaAPfABveVCKn4
a2BOClMfmO4tinsDUCfneooeF32fMW9yyt34pF2zKOtXj0XrU7TADPTpxv9c
MesXGiriq8ZcFCA5pXwZCcw/WzGpt3Q06OZzWqfvECd9YxDm3Aa9Hfh6tHHj
p6f+RGcrbPnXnaxg7nCBg1KParWgZsXAO4Qxcv0phcozgZs2E9nv1HXZJLU6
6UL2b5cmDt8ZHH+kUEvLxVfJJ6yGiFWMdhhKxK5C3rJ4sq7bCl+QaWT1YkUK
NEbBiDVm0/YPjaUD8NgLJwoe+bZWiaDg4j7iHWv0xXrIDZ/twITefhkU2n49
+1Iv8ezaQ2GDIirlJMatTVA77Eg4qbadO0AEnUj1I/iYTvg5kRAHZqkphum/
TrIQVNLkxYL2h3ur1cmzgIUI1WlUZqUF3wLA8TRwQlEn+q8ERyfCokx55Ep6
10cpVjsnsGprsi6rUDjsMUFdPt535JvlEty1JIP2NXnwY2Txof+QBHIEP/Zo
f0CJCXA+Yu1mRrMagpPiaIIkYWiRpIkp0GwA09nIaAo0CnNisCfAcvxdfy3l
oKF7Z2oRpbF+do+Ruup8ZHMgDqkxFykqCAm5j8kJsSlLpnNjq5aOxN49sCfI
z7Vnc0Ui1e2QhExYsEvkNeDYY+oPkaJjIPNpAEkibfhCzuvmt2CoUS8cncbj
S/lnt1trMXUNQavHCsH7lWfw4YJ4heg5/hP3JJ/uTA/9eahGcQtHv2/B2l5Y
BGVGCScO81wOuws35dLwftVRZzwlDN8NxBpwNOmz31vIafXKs5M2xqf4+KUH
6UuX/WTsuKYsTWuwp4Tcdt+YFOe5hg+OH/KiGPZ32x7CweepTx6U+L2Wu4Gx
JT1KEc4HfhBBYnyLu4uy2SgZJB9XGhC1xFaYERooLA3b0s7YblOQcoXtAH1y
CU/CB1u4t5t/Na/sqcmOZVt2jjMTWOXUShvN6S3PVvluI5K70UHLZYEoKlDU
bZ1N6ExgUPkHWM7jeq8k3Y0MsW5bBXI6QN+FBisJ0r9c9qeVXrvINrdveBD6
97uzRlxNKvpzJGeqKoAOd+u7wovAr0eOmLKeoEYfopdE6mZLVTlRzemd9l3V
xwinArkX8WDXMpV1LUCL3Br45Cuip7bhiX7If4fJ0Je8zqEsXSI6SYzF0vU+
EzJSpIQzq7XagZrRLIGBVwYx04TkQTPc/gu/asABkInPfcnQ8ZNKcIPFXuUS
9u213jVplH9wYxngr2UIt50cJ2QGkUoWws/vLleVU+FW4mayDiJUe+u0/sjq
ZIN6K3VkWRuH/HycA7QxHEw2GrSuAJSe6tRokSvAfao+xQR5e0wsvwVQCE9o
ApTDBOk88/S2j7nRSbmkiwTP48JeRwrYHK+o2Wv/kS9nqhVoMiA1DhZhmSZv
ZXeMbSWV1JufLQX889A0f0vh8BBKNY0atEx+1SezT9bVkvwxhLIB/GO+RxUD
4sXXIQuCMUefBRo8c0ZCe4d5up8tr2+2QJwzJZdCdS9BPW3Zyw6v9mU8syBM
iuREszNNwzNDdfoLUVJQeQ4h988DkVxfLs0k4qXSOrOi3RF/LmvQqHdSH4bN
xDDCZlqcELm45VS5brB5vHQO8kecCWCccA7yMs2R+SHL8pCcNrSSQhL/n+4o
uj+SPrZo3Q0qbywB8cZ+IQAoB4oap08wM4+oPMt9ZsB8YdUVEixwS/dH9Q3e
gYBXRyVPkU71L37kMtxjJbMrb7noeVfglpTvvFjBBPjoRNUNY84egWre4TvI
lo6QAhgYqvY0ZHTotk8+Nj9pqAjA66qCJoHK7GcU5kDZ4v24l1lyjyZQAzLy
CqlFJdFpsexlUqzGTRKYdXJR+wveo9pc+kbMcPVf6B04V2eU1j8Lax4R9s0J
0ZRfO/lk47y4Vw7z3CfdeI6TMantYqVHcEWAfK0pEQ10vxFQ75xYOa4Bqow9
YgjwU/x7cn+pkhAWC9aCUElZ+oeCyrVQg+sT1W/Bolo4De9inHqRxNwFJt1r
cOyHL04GQf9zdbNhzl+ecPCAwZTVZ45JmeIcjIGP19SFIKvdRbrUnwqi0D9f
Pt374cfOdyNjh0P3UbmC7l91EWChgy1y/IVQnsI34Uj+O+CwNpzJfmL8D5bO
4H3+6xn+V/n4fJtbzGMBVSFPepueQnJ+6nNgAIYgVtyMFQlTmRBZvRjko0j+
js7aoMJJdsZe7loQRfgygFK8c1rA0jrUNY3koEx6Vd4nXlw1IvyMjuHLLQl/
My0ZcSp3Iu76WxIY6KF55zexAVGxFNopzrFXCDYVX8QIrJcuaa8WzySjP3Pa
UihQYpMCmYpD9u37x6qlVMNYg1l0BQBUPSvBWnfO3CefQzszWBFi8fPSZN0A
Ia03CoL1rmBTmuBxfOWOhUuIJwJvtj/DAmpT0atJVVZvacnqncMRGQx/xHH8
bQRIIh3zx1YtC28aD6elotqxGbp/dfIE1GpnAHBunBboSHq8/+gXEZEbypcG
w1RRrxM3e8R+cOxMjJ/f9P68hBXxYIkNEW96bbaZgbEFU7S9x+s+o/tNJk5W
u4Z/9U63eaiI8ERf61d4LY38kMwCVvrQCpgQHnXOlLd5eEcSr7nB+BA0kRnO
95q6eNVPM8OqriXRfp3zVRpqXkPnI98sSjZSzG/dZhc/lHWL918cGrTQLusF
eoKlg4kvKHQ9qFzvYDCOXI04+ADzCEOKmn1j8iNWDYVg8zhKOqWfJFi4O4XA
EUPesiJNKXM3iszzGC7Y0JeyEjUD0gfLsvd4ggwCS8bAukh8iSpuVgVxFG5h
7y/CdgEjHqOLeWJkCfZLafHBszxgZ3IT2AGpj8D3jlM2QI13m39T5gvunjvX
XaZRNTu18+0qwNT4QM1y/uvkw2xX/c7nxsAWPTh1ihBNHsfQKJBFEuSyDCox
bHFT8HNN5KYxwCe68GrJkGc3LpHmZSE3h0LU3OrAgqmU+cjaYELLN78r2/+D
ElkyXVAJsc04PkuhY2bJwiL3lp9TcY0SYv0gYkHcgfBXaRhlKHs9mFuTvcRL
H46DYbeSQjn6ee3FO3/L4MZaXKwOJM8xiTZOmUiLMbli3fNXMeEyEysfV+2Y
JhpMoOKFP23RrZMLHwowx+UoEBVE7f5dJOjJSEy7uh5CjdYNLe6/1yMFdFMO
dkkBXsyGC8RijJvIQAwZv7IdfDOfAYF3d07IQI2B0bMbpiwGWuLcYgI0qXAo
PceKq6Fy5fiMnkTGiWD7Mtg7xcJS5htorfavSt8kx2zOP2BiJulW3l98OJ6U
xFKun9nQPktoCzHZdrgSEAjwid2RMfVzPxs1jav3KOdFj3MD+ZakHOsdrcDx
tk1PUoVm8NZbIeYqWzgStGg1PLBJbyWPoVsxQbzUQy+O87sqJDAC8l5GcHAd
NJUeJb3NhYVxivYV1Y0yBYOZ8UoMrRVRGZEHQCTx72rY+xRfRVytbC8jUuZe
XZEWP6aJT17Y1m/qpHRZMbgWScNDHGuhH57gXXSHa546Tw183MQrhDv458/z
/YUzDnBiptyJgP5zsmCsatyyRrmHO1A86QesvGPBgZrrJDPQIkLrqg2b/N/w
MIb+p0OY3MoZZGRlzQzA6Wb1M/T6ZKo42v01O9K/nIQEiZ9r0ejnLBkrf0Mn
oGBwKAyhwIDokxn1vbQrzGgA15fMln9Mj40MgylWxQKDl+JgptAvpfeRzLgE
Oc7P0YndseAfW3dpa8cuzJC2bWrxOdhEUFNkJVInOfAJERwiw8KIE04TqOBz
WrIwKf4VDlI0Iufk+dOET8Jbc1a3KDgjjDkgL+wgJ6irv4vqX2KpCAs0o2h+
juc1WmeHvfABomCrprJnfYWuAQLznjNJLve/asOGNIWYhxq4uI6sBpK3J03L
mBeFxFFfSLWVrngaNSxRyvOJ0tOLnMRjI9EC31cnCKbqXi/X+BVLGU7FnPPX
s6nMo7R39gWqSIm9Uy4bKW7A/NyPVV3+HHl35thlSU1K7Z7nU3iBQHw4e8BH
r26IsMR7sgOXbB9wuZQ60t8jiB9BX+IG5r81liMJE3fu+niqV+zP+HeA41bM
HzZFCiCtrnLjgFgmoIYIVKalhJMNcDgtuCoYfPGuzIZJBx61dEe5L7BU9oj2
uIFHvIYUujJA0qQZZY35PJmLiJb3AjTwAdb2z0eNRE5ck9fVmDQwyIhGC+3O
QwPGpIHRLGlJnOAgnOODu4gf6qOoCs/HaApU0+c382EfhsVIHnLcRn9Yi3tT
/1QgN4JJA1ME1o26M7va9FCYXfzV2FYa7Lj730pt0Yqiy/BvYlHOQhslYpA3
F3483qUKsLqx0GcwHy3mzAsUUZCEp7LE2H1ksT79esG5EUdBI8tOvv7uNUeC
r5APdEB4zByG/Id1RU0s4jhfLYKPxLr8bmagKfluDU5k2k+Haodu6P8Ih63r
pIVZOA2G1RMBnnyXYe7X4/NEVz9M4nEQr5K89upjU8/B6YtAzZiVHofyRTlX
T1IZmrkqMIiG0BXioqt2pMMwvKof29+oeyEzg2ghZHh7VnbFbGeGu4zWIkGv
IVoFEGqxrt4AttMOFaboYpxMHD6ZLBxEG1cQKwHK68MgSFo20ivQ/+LhciQs
MrwYAbEoXxRq8yS2a5qTop80eFGQ6XJ0Kmq5NGFI9FGcpJ2vpH/hdnM3Dche
WqjYiW5X/rcA4R2LyudjghMaXhMhFJ3/omauyH835UjJWxrlFJyTFBQtWdO2
o8uvqptsL8jSi9pGoB/RU8T5ypfTi4cC6t2PJinX2TbR6WS4wUmTBjvMlV3S
JlbEjLo1ils0XzZd1bs/WATbctUXmqo5NlM2GPGktoxleBPeWiX9fns15+MF
53VycDiyHFw/ImS7y1lIhFUpXYNGBWLv+t0tByEACssESGBtBqH6R0CaEacP
dTnSL+yKUhc5CqV53h7pn7b0E+tRI1SgaWiNk3v9TkmQnRtQxw9J7li5j8V4
6SUhNNTncFtc9cjislRJz9MzeRAzpqSA02ciA5YyUJmtn7Kvi/l4/CpVByaq
1kaHUCMjWYMwdRbNo77B9ziwoqLVKKQWU3oLjo7+XhaVlOitMw0IDvBIqzCt
nc3q545r5QytR+hlgOKBDJjKcADrNJY7WiGE3/Dd+kLJpM0f4oUvKxQy3y8E
6uqrCBTo4bQMgH+trhhJzKKzJ/MSqxNvai4/Ni5A/TWOO8Vfi7w0NKZoZp38
hhT73GWGJUjjlesUkrRSERnJzMJbGXNahVszceIc0+44YWv6+1Z5C34abLZZ
6weLzvbsxyXPpGScTlUkOocropscwavQ5mfGh/ytmRaF6YYRQnOqHRTJSuZ0
J4CBXCNEtO6VpQZe16SduH04MjrAJngYY3l2U5duh1//D+1DJGOp/JsxUgEG
lI2ZdbUWM5F6HNDxYVCQRPbpnLegCau/NlBvVNs+Ued2RScXqX5QSsbQgFVB
6V52tqZv9bsDcAX3OFG4zOg5wb0/FSr2kT1iiu4smQHC78z53PH2iScvUM3k
fhnLZsNrexSV/lWuoLm4ehcFZhU1yQWVJD3iGjC0fJPxKdyKUtGryDG4PSE3
oMl6UKChI3GoGjiqSMjjvO2ZVwcYC/KzbbFpQ3nkvzVo++mUC7Bxq3JRHiHD
dni/FLEhwbSSO9KPhQmTV7xpWFesZluQZ1cDQL0A+ER3ADsiNfH3PPNtnowO
IVRqQMTi7mSlMf7sAJgeNCqefPshSXfMaX+9bykGy9jSBwCCBnzdj/z1Nh5a
PPC+D+brvcqDX07hep5P4+5S+dLgiisfxnm/GobTZ4fSfkFjgfCIhj725OWh
4o0CoRwv2MBhWxz4bSVSYO+hSkEdQ6F5fASSc3jrpzSSNCkRLv8/BnTJWNRH
bMDPAopgsCbbshxuJguRqYzKn080V3smBePjG6nlxmIvbO/eb0x4Frw+zI8x
uMRVJBkTdKvJCfZixPLq04wZPozr03ZQkP7hEtfsqh19LctpUYwT811JiSzr
G8NjouDUVtPQmHlV6KUTmlllN97KEeJ2j7++yy/ty9+cUVjNuWE0rurzXaEj
Dpy6nCnybZYb1v8iZVGP6xpWZE+4+WtVWiciVe4+/K8PDGxuV/O828NAVW5c
oLMhTzc3GALGwBQ3TX4gp6Tczrck5KTBQfbChCb6EeqAgD6ShyCDRsXqFB1H
MS0OYxwiGa/G+CcCIBu5ScHOJ8fCV+MDFmNDykSyFiWx4yj6I1/V5TcNjOkb
7Qb5dRah9bkY8Tajsv6xt/2oa++xePWgaSdVcQ0eobuw9ZzaJZEISODOQPPM
RowQwHNLhPIu/r/8J0rajuaTFlVTeoIr+AIaXBkkPmlbH6n2WZ1iRnhqhv8T
oZid1crzFq5SR9ytCkBCmmkM6pMn44UfuKP7lwMTXqJJhLWgR2gCKXrzXEYF
qdLGDszvVdkCenX/E1L/5Bfxi/dQ3lWEDJCRbxsL5JGgjdApYcKSHE7zk2sc
yMYaheVOWI1d10gcD+wsqgOJ1x4ev6z3SfiUtjX9CEH3/Sbkznba70lYG1IW
WcsDBlbQUIEu+CvP8uA3PjsEIxagbAz94ASXaNXVZgci/awa+4RlbiOWhdxU
cM2H+bZEcnKPaOSDS6yamhCAGK4vlTULxW6WHmnSlngYdDysk8EadiHjjVdD
F/CYEfvqYHqcMiCY1fq6NclvXabOGR3BY0QAvakjlFIrOj1ubTkmflaQcE/D
85WgW71OQdaN5buRuzBNaI3YZEeSr3KTZ89yJuI3soXWpUoEFyrqbIYo/BtK
pdmRTVPperZWpsLLkgshY4SLlchHUafnusvJDzoDufFoZu1rFfgr9TKZrcr+
MsscnFNBD+0D5YL8zRyRF9jMk0ttFR+PEtwd5AL+jJBmyMrkhwcy1i43Myq9
4uwKmd9VX7djfWFlg70qRP/dnVkPZodgyowfI4Nh4Zt8IDIeCOSsT4pQgR8+
ZfRk913/ufqE7kHZwoH3qJAPuoEjLz2cee0hlC2wWfb3mSkbCS5C3FGEAlnZ
w+5Y1dLXZI5ATNi93C4h9jT4IUsqG7ZZ5Re6/0mu7n3Qst9XDBTv1E+WZ6dF
CJBYC29wLkftBpOiGAGHNXkhdkQ4QUcwau1jpiYuL9CU7QyTTZxuig51O8TY
T4iBOrGj5qNj2Bn9pj3TwhoxjyBekI24tX+Va279ImRuKg5QQLq2TJ2HhlHe
7YZ3DmF6nGF9gq0lO8kGLcswqBeKCIfcsxsc2hVIx+U6pFA6ZXzZrTJWSHlO
dz2LeELMfpHano8Mnt7n4GGAUXy3wclcQMyB6TDn59iJDkNPC9pKEX4elcnB
riVCKnxR/QxsBIOu+u5u1Pp2x+VlMS8LCIEKbjWlFG1ddLtVPdY+gSntGrk1
A3GVHkB5HkKXWaNGhTwtFPnyce+Ppmi4YGmDPnbTrDzA2MOCJm/wOLTq2o/a
zEe32NP9jU/xnBtuQ6ebeniqZuiC1+eNRI15/TK2wfdmGJD8U2Y8n3T4z9pp
V4RjXJI5CxFn30x2tnoBXKC2lyjZmt3j7qGAOe7OGv0WmmJ10SYmYIs99wYp
gOKVh/FB0yOzzBAsZ7O6qyG3EGH8k90DFUI3UEIJ9HAIFUtUL+HHixc3Uiz5
uH0XOgKWmy6m6Vn/W/RO98zQrgBw846K38w8ns4S1B4iT9z7u6pPmAjiBSBD
8Y+7hvshlF5oyzVjLNASHixMpWtePLSS4/pWg5nQAbPlzfntZgxgIx1jAxb7
2GcNW6p68yIUKQMs8ki/R1SG/khJ6h3YX2Fb8dwKArqHXC9t3GdDZ/5KuoOD
Uq87z/CUcrvCRHm150DIkkDKV0C8hm4Fs5o9U+VMTSNFxy3f9q6U8kW4be//
LTyMy7wL3Zdy8BU0RNF+HMEzgPtQ46PlFK45/8/EV6WlM/fu39qWGzjQOnI2
nT5666UptezmzWv/Dx3eAGjOfo6D/xvDgUTwTNUoxcrlIVD3Fh5fPGgwVrrz
Zoa87Ua5KsYeaMgz44CfJYxaj+Z7aeb3BcvHN31XE9S+Ze8PaLi9LWwBVHgQ
0wl6IgM8B6L/M2sFwRNdDlrc9rMsfPpQufjHUFrT1ymufnEgeh8syP52yCOd
+cVan/iqfW1L47iU/80D+Woz2TeY+QHVxVPDLca7G2vgkObBiDz4F/NyVQ2B
kEKT5CZB862IkvAAP/dD87WYWFjKeZF4X2365crcf4Drc+Ihqz4HOJge1NGu
mMhjiqxrtbmdK7dX262cT9jyzfS5wlmUsD3FyLLUhWjVH23SaVo63TOdd6WV
z0HQeuWt7Yi+JcNfvwd2wOeuo1Ze7D014WIXDWAV4Fqts0ngTKecxmAIPT4Y
Oxy1utGkii100wWidwWCndAZAXuC4TiaolZZ6msdvE0HI08bfcL/WUMZnlHv
aRZw8YMNLKuxD4G+W8ymg4ITnt1WpaQ9PrXlunvPcrgvobqbbFcctfuKqf9p
RteDTnZuhfWEsjAdMmy4GAOs+z8HpmJR6FvtZ61r+BSOrQnx7OFc5MO4ya7o
0Jx3GcagsEG9lF8bgnVbFB0ebl7iSeO9KED1Wc6Wbde+e+yj5cGJY2kF6wJA
corz8HDRWgDAdJxhTlF7HsGmONY7Sq5aDoQKiXtNQt2DVjVFkFjKNs7PmjsF
rLOZigXYLtO26Zwi2o5w4MKF3yaHjZfkqMdDiIcts+aTt6dTMs+9CP6b9NSV
PtabkP3OjsMPhZ5lAwcQxbOZhWr8gTjeYgbg8sE8tai21qPURQdHStz9XGsP
MhKPUAnu3JVntqS75TFKrkfLhFqBl/T/dg26QKR7mFLNxRSBjvIlzcIVAIPj
e6cwjYJjY7zivOunxGQ0LvxU4alRnd4s9Hkf5kiOZgrr9A/tUE3hLbx5siTZ
iMUw2oV8Uk3YfxdSl2YpNxa8ipEo48wYN2Skrn/mK9ZAHPGRpgkfmEwLuI/+
k0huZ2gFm6UublfMQyC+HZS+ATXaR8E37DI0BzM0eaH+mCqtxgiIO0raBne3
3I+iPVEZj2wPbHB/ZMw7KkArJ9XnZMgItRZGL16Z9FQvUwOrcKaqd4ISafY5
7DXdqYGKW56YVETIfAN16NbLmwBZAc8Uz2bjKtVBouwG6GADlXl88toOU4qZ
XWSOTe+HYfKh7pYQdqX9s/HulYl4Dj8IzUV0FUQHBxAfrlEaTEei/Rdr3a5u
evObbMk9t4Sa+IlNu73W93qReGd6wZhVYkp339fZd8KO9SO08szRGApIpcwt
7Wo1FHS3Qjy72kDamxcWOZw0sHSa/YYj0HL4AU7fKYMXVbACDRBKlDqslygh
UBMTlTEt2Tfn6nlr18pM8Yued6nGzjvWDTFAPM2+NMw5wuBDSeuT9v0DBmtT
yFUeP1NNNxbvpDMZ8aXepYTqbS8q0oofE4M218mXYZd1TqVTtgAVk2MIxv1R
S1il6VhX3vtE8Is44AfJtvWtrY2VuCUqN4z2D5bPSqNUqyCNltLZjntxbWRy
+YtKgUcgwKwdQoco/OHlodK7vBIUOplkNYs+DOkUdmY7omh6MMNtXrJDfg3N
baveEjz3PmFh3KnJlBqnnlVgn0pn8TSuHJgp2a3BOEbDK8Zle4GTOhba5WJc
ilkyBaqUq4KRy88RohRQS/57qgIj87c00u7Iqu6uGa6NJYjxvxg+0YlRiZW6
g+IeLCr5igM/qAyJ3hBn1AIZazXruJP4VeGNPxd1hnokwwbk1H+EGmcQJiO5
pbMrYxuLqsMOmpXwT4pLZCjRsGjNEVHsu1SaxGRb1DZGsHVJWYdegePzYfhE
lsjHBmPox2iKbI35Axk0KqZkmnv+/x08dO4W+ZzBuOy5603AZW5O5VEABOK8
NozF6aHBiqdcUO5ogv23j8n+fOdZB/C5JRrYalSOn9nd0f0CzgrqDePHMcdn
CihZ4IYvUWk40ZBhtGUFzbHBkHtxJP7nwLrtNtyhvPxV2xgUjxke0BNRX+Y9
jcJvY1i+7ssVJ/tRlxLcn+wxic0IcMMFhOV6XVT/Jbw+XBcEhtuptD6IBFBw
B4ndZAZX96CedYxl2g3TSofy9Dc0Px0EqKvfX+obG2JC/c/iyvLcaaJQSFRH
aycy1Kw1mFAE3wkj1AFbDQtRjQn4PS35eKRPNx76JQP1uLIzY702gldhO9f6
qPFgPynpT5UuFJ7//B3uUtlqPFNerUz2ZYcV+XKW764qLV413m+tUSY8NJ2v
n7eamu4m7yNLDRczXMCVZPf4zlUBFvwnk1R5Kgf0NiSYn9SYEPJ299riex7q
AcosbXstuNsbyfdIlMorfXW09u4QKQBty2/ea4B/ZmyCGQ59VYicHyrzEhQ+
qw7BcKiW15vih5YTAqMOMA5w6CpuAKGbH0o4YjHho7a91pT950PmodOXCdZk
EZTNaAHe3TIfmi6kZVuO7o4hYI1CgpgblhABdqdJxLg4I2JEYOzhuWqNmqHl
BJMgIVu+JfvEMGd6bEwmRAfVO/RWdo6+5yoAPVpdtFc/aDGnzfpkw76cww9/
49qsBacznLPRcEhnvrjOJyXSukikRqAXAC6iv6NPRVAELmfgN0a9RK6rsNlj
r0zDV0sNfQzOOxLwDaewc7YKlcKiXpOwO2sdUGNgvY+umVmHzW7nRY31Bgu2
PBVV0CIK0mkXpeFzWdtq/6yQYr5p2kf+8yUAAUgcopWiPUk/0NB2aaOeRdsq
fnUpDoFK/uM5slDGJ7vBf/deiTiPYGFMwDejaxZ4zocLWjrOTGbl8pF4ELfz
CUhwDaHxBC8OqgGibR7ur31MJNYxYqw9bTTfB4yKNKzUyYaClgs1OvMeRnkT
n+b2EszVvjT1+UERiTc4CRDvaBuD7KKg89IXre6SbX699U9c7OUMl37pS/X8
I5hdLtavWBGolIVqwSgPddmDYkWmgEPjUGFrZ2ZDUCu0tEEBWjLqIC1yZ9iU
bQEIouJcVXgHgxLOc3et02aMUdUkTN6O9CS4YaKOdjGSGByOoPCajCtzPEu9
JzU1DH6cfBJ3Ex4ANofwfJuCwOlxJOFhM8sbm3HLlUxPvOPkrCEDNgahuBZM
vNZ2fch60Y8m+wrDefMrlKWkDW6clWY8i5hUr6udy+i6UeLu1tFQh3rY5nU4
GYgBvplHKKtGoFXbyc4mp+YF6t55TfLUC7vHCancu19QGWID++KqCXyaruY3
jOeQOzXe5eUhd9UfADXKWXqJ4pepltSj6M//iNgdfVNcYSdfK+zC83abb6iC
OFl+XDWT0bw4sjUI7NIk/mh4Mk3za44+Rcs3DcbKzGUgYkuQj3/CfAi/fIFw
Xu0uoLd/vuNppmXmuepRjVP1A5GnStJ5oiO8Bi7FQOhzBdSxtxF0U0l//Nhd
KqxoAbIQQ1+X3wQrh4EWZINuhnCMRER1jC4g/GM3QXHmTJAFld7AB3IUHG6z
QHBPynEI+jllPqybF8yxHj0dhIy7fLz2TwhKfuLkNK1p3tHMF4uanEIUhkGW
IfgF3PQ+yJCoZrbiLZfnvQLRO1tQKBnMrgZDvgxgblfPfLya8UlS+MRMoC5c
GlVrH3EvtPQhjqrdD0u+WFja4RLVwY3GElox3DZRAfUNTcRRtErZ/vEmWMi8
kvpWkYKtYWrNtlXCa4RTXAiKg88ArJDYXNHacxgnXYq3CDfO3Js6tsaz0pEK
9bIsE18+RERBACiObbF61gd7ZCEtG7gE795GZfRfczwdGOFc0xLpWdQzHxp+
AnLIhA1aDdttCv56an50xFTG99FKWkHy0B2Q508GOcRNHow3BcN+564DHo15
7L1W+MKzn7nRnipNP8Q9sYBNmnjM6D/HVBf4w4+fHphKRWxo8iHbnpcOhQw2
Dx5f1l6haKPu1k++hJhwpHs2v2IbFS9rZDnAGqkkn2PcXfWsOoB1VKiVZLRX
KoCvHeA/bNvm2tobwCjwF5S9CXoRMK1Hf/8ucWc0bkmauvk17lhLGpNeK7r0
tG427+1p9Et1XlUSr4GV9B/SacSY+KBmFibdTlW/NNh+uQdeYcs+zySDGsA0
2m4PwE+LMRaXev/XnmjqnTXN6q3anClZ5sJpTEyN3nh9nRAQ8kqkaqX1hI6G
1q6GQiZRrpKgW5FkcSgUBXCiar+i1B/o+G3RbxKyhuFtAJZA+w3wdegWKooA
yYO/dYsqNaTQXxgnMBz/hvvuBYNUjk0LE2DpXwn5Mqj0q7m4sgHdsdyZNTjB
iNautgTrun+dZPhhUPTU86uhHHhwPckfxHtrLD0stMDDn1rlWnzxv2hj0tky
yr0HPITky4s8mMmYi4tHEZ2tzLuSxYhXS1yf3LiBfKI0QffAbMMsYLQU/16S
BCbWQDRx9OoVCS+l4MG8z+eRrpadwhJv5EM6hL2LMHfChgGHTM8RIhHjjQ8I
Pnsc3fpsLTB/rJctMXYkKRIUzKbnf64tbQvTBB9k3YHcydNuNXBJpIetqcgY
x5V6aoC+RfQ55G3DYgqrJ62SOMNzWXQ6el0BmUXRTcE3L1ERlX2uqgahdpkU
qjrqLgGXJqMI4/FBk3qjM36AFunCxn1qUxmjayXVufc2uwwYH2NZr1dm/8Z9
EsMkJr9NQvL8tbk70MCfZy0FVQsU/NiQ1GajvoUT3R54kvxb+PNAOkNbjiM0
+YQUWQRIrVbZ4Gn8fEjlMcY80tJ+ut1KjBkFNCEzWZiTrrOe+Yp0QBZXgoob
4VQdDmHu0PqHXOd4E2iHnvnOWHqybS7fHl1g2Eq05ZVR0KjkKxsQTe9CEtBq
T0uyV7JGwOfRvXFpHqLwbpPn2znQSegLUmE5q5KGEoa2uvIrvtjmuW0jWjD5
z5aZYChoiJBGFs1fzTxRyAeNpOOSZMdhJHZQaCqx84HkegkVPgp3apDvg8/W
PkNSWZGWYHwv45Waw40JwY4zqWbxtGlWnfYJW8ilvgbxOEJF9nurxntudqLj
n9Bb8DGbhU5SnFbVY1lH23nXPApmmGQ+v53IzWqng9v8miIa1jlkGnFshqjf
RbyESu5lrLNTbKXik5AFzCXXyHkWAfJV+0RxxrsJEKJ0dqgAFm887Y75ZqL5
MlHhZ+7shyyQ0qMdsrurgn/r3uvEhxPz+qs0g+jVYc5JbDwQHaKSFezOQwxP
50yLEiDpqEmZ5U5HgjIj9H3JyOKg5HDIJ0LBKf1iv4TBogM2/o3/ZOTmkShx
UTg0wLHt7uQOtorOCAD0vImWtniT9er1Ld1q1GCw61eTm94Hw9ey+DazFkbR
AkE3QaVER5muUDSgRZRbNwGesL4k2KcjdJ/OAlSOFC4ejNhB7UcsCNW/5wcy
kgSj7M1R1WA4FSxELXJ4QT9xy6mdUu6D9Xb5uaSeg+rSnF4gpumC+BhJCyW2
3bxIpHkkU6OGZ7bGl3Z2MpeKSjut9Ck6vgkod7S9e1LSHa+xs5WGO3CNeR4b
VOR7ss3TZXnte9wGZMTKCLuUjnXIpyriYP4hvJ5/41VUClSqnh6lRrOWjgsI
vbh4lY4NbxB1MVE5JERfPo/xtrHM9uJJ9+e/mfJljTAGzfSfW7LNXtXK711D
DXpkCcopfXuTILAC0B/OXUE9gDz0t6vgz0903K1O97/loauqP+Tmt2eP7V4E
o4OiV7uymTAVbjXV3vvGFv/0C/3ZIbTT3P+Jt+Tx6T+em3v8871xNDEhBk5l
WuWTodpERi2B6Kqd9Jl4+DVj9k7g+tfn0JA4lqkSq9DnI6nXY4GC4DfRL09V
dun6NftOYJ+P3SsHMqsaKACr3Q+9ZS5HPRMjsXih6CTAA4KxvC9o+bDosB53
+VH2sVlmk/UAP4G8djMs+Pjs2w/BmXlTtTDj2ETITgNhjTxRROfIVrMWHY6L
Eom0uxsjh5B1pyZRyY88be1Z2iFM1Dbf6kzJbW967Ul8j0JlyV2NbDNuhU2E
R7iGUmjOG+46nDk5lalhoBDVDZczzifIxyh0mq4clb6CZ/2NJqvp8bsu/eKe
YkimKks2lSPgZK0dPOLGy3EZNfnYd+1EtoIAEc1+ln/hvsN24pgcacAj2Meg
Rn11vYmyrNd9FSsFN+fXeVBjPAndTPBrd6BCCDo4IVotTon0t+BqgkDk+yLL
mkalSJ75Copefk7sc3xFl7FRrR2lBBxdERNet3MjXffEAaYiwXVnAwjUt0YZ
+x83QRuIQQiy5CZ9MkVisK0xnYtdGlWCC4ng3y0T8ZseO7p9vyvKbVlDQQ19
NstmIcMh3t9iOV0VFuHX5vngse1pUpQZ/Fa73KGtaIoJEBTaT7v7sBLpcWUL
Vc2xKr9B3VpUdQSzcJkJSKEGAGOoUavkG9vhEEqW2byogpg/Zdbd2Y0Pf4my
KBKsxQoUsqHyWX9uqxt+bL2Uf8sz7KcWGxBMUdeYfx5568i/9z2GgZ49F0H/
484uq5EEvqB+5TTHqHQ9dNFBDTCMPAJKM6Hv3kLrBwiA0lIU8bzWsyBYlj3v
pS/GqZs7LTK4fjh8tEzPtRfcmOHsVF5YGln/HmQYI92e9vYRGjirn65Yiug7
nD5oj5RWx7yYXxtvyTiae2DkIUcHJdBKdjH5fRnLJnuhWeqU4XUcie9NtmIX
z4fnIV732XpK8MG8p/LL/Syc9SJazLxMjOtlAplM1DVRl+/yjx5XpPtEdplu
cpiZrI5dUe1IgfC+/OoboiUwR28Qkdp8xlVvPR9nk98hCLp/riYTiXpaA5BB
vqd+z8xvkY7z0PRL3Lco7oC/OlrKwDdM9e3L3GmJBHYNQZYZ56gMeHgHDFVw
RZeh/fthme6CkHkFZLQiXuncmW/7mhqbLohinu1k7bV60loHIiiOrnbj+2je
n13mMUO5BfjyWppAKKab7AKCmw9fKDLeYZ5oMD/oy4x9lrleNfrQZqESa3iQ
/F6ME69XZ3+Xm1VhT8ELH5dk3OWPf83F3ypWjdMkPmzvJkge4Yt0Zou4bZxq
XoeYo1+3bUO9QmxdM57nBZETATvVW+ZzOLk341hGh6u2/hoGANMoyd0i/3Tr
fCMviveqXBZywjaxO683z8AXlRph32pbOT+D0zBPbR0qAQWpfG+2JGu0ZOU5
ncdjANZCLMHRQc53RdzYKgSoQUyITiXa1qi82yK1RuGaFzmsCucm/GDbprBR
2cOQtsQ6SJZgq8ZeyrKFsItfNNfjun05gIIKC+tkEJa+WkiMA6qyi3uBb9DN
uHUGTlBwGK+qBRclGzXNLOaZnvbXO+LynIV+IPPJEZ/IIejxfGwz1x9nnXni
KzsvaA3o6Ekin97itG//5OtZf3OVIczyO89+H1MpPTBXsZeC9r8kOIO496A4
jfQwzCWa9neqhnFHX46BiyW6JosmzinAzMPWsCV1uX/jyXDASvd3+V7a/MHo
L6A/dwt1AWiQqmG8kk/o5bV9u+Bn4WL8ZZqHmlFryQxQvdqezUQFUUxrogSE
sKecKwegiQG+X8k2XQIxDWeKg3LbjLTKIcgCwW++Q2SebWf2HEQdoDC7rPYZ
4STFrY/VGnUmxA27BGlKM/ij1TkX9evcmGxHRSAFfTL8gTfIQKFci7RbaaQk
z4H29l198f+DvEou4xN5GMOYCpVmbCVMWPrlhXZwRsGVBZbV8uMERTjFDoxw
iGtyz35LlRGU1nqdNYspHLJkqjI4iBSTHdR7Uyu+CLBRdYSXXAJR63QWYdHI
8OLFE1BuODE/xoAK8tZ7hgxBuyKsqt2nye+Glru5WmhFQY7njnl+AkuJMMxA
bMBAL7lmX2TaK/z7o1vRZasH33h4FiJONiITMFrN3UuVMg89dABlEu0Lkl2R
jtEHNma6e3YTwz5ckmnGhEIRicV0k+ldFAiTerHrK5oL5YKaBYa2EhFKO2+W
XA4XsaZC5BKNJgT2Vrwy7mxQqUg+TXLErpQoD8Gj5pfD7UWuOjaDZMZ/16dr
Suy3ZakdAyxC068xgxGtM8XGRhnCqh06QNWgkmggvGPZgcguIKKswuPKgIqW
WKb0te3Wp9oAk8VrlmZrMgNhbvRXiF6l3z8Y02Ym4ZJTSC8QjDiAloeYmrq6
EdjpCPu8wOml1aJpIGrYiE5acwbhc8epYd8fN/8k6NJTH5D43w8qmuS8mx49
mXwsSJXXB1YmlLCCjBJ4suMV05dDeRLyfWoj6vYctfKHmd0OEJ7LY31vGzif
st4TBZJLSsscW56vsIfWdV5p9TfMrXGbZlEElHt28Mlt/el4e19Vzw/9MVcs
L5Xif6bwAm4TzzOyH0S3E485ROQJgitGWABjEHFurULYR1ci6f5RBtSkFLlH
9bK+DKyOJZidcmMttmw/LKENUNLgrXI5p1Gbh8Ax4Ydq9Pfmq90FDIQ9oYiE
Yc6oB0qciFNA+6kabsDjk5pwO2YK1lEOTpS0iQpf3++Grxi27L/TEHsbZL6d
M05uFKU9+emEhfvecyucub/FxfnARL1c/Fmnkvp70WmXokSYZzsu9Iql5dBx
SegXFYK0O47pksA0S90aC+QYOqZwFCL3OGC1WcTzM1NcPmpnrI/WYZkkcm29
efAQZqr7Dvgt4Iv/DPdJACRKf/FnTDKX/TyPNcApp4+lwYpcMlHYZ5CCJOfN
EhOyhf8dhgM8zG3r+Rr6n57ILqzR8mx1lhXdI2lFiyN55LaNe7BQyaF9KmJd
3tmQKyInw32oRWqyBdYIaZPehbvu9iDzc4p8Bl4/eF5KyD5G2+VYGAtwPT10
HDhsIPQ6zsshEl1ncIHBzwuBykxfO/epd1YaXxd581mxHFxPzDapPKZ22lWS
acidVrjTXfXlZ++prbvBPUDTViCfIDrmc+TKV+5hXzFrkHc1Ne2vXDm0LTA0
0bmkrjiGXq18eIUQ20qgtx4+6uOlcizOTemifTOngb6U33jzsiAS0eOhsoUQ
SGj9upSgxg+DrtwZIna1t5jFpnWXvlzMicvubm9C+uQZsKiKet1tMhyiSwTZ
6zu3jEfs4hkMLrzGwgBCqAfmiijo/XrzxGqDXtYh0d2tjXmekT2K8lH35j9I
Mo2ZCvxm7ev9O0dVZ7sXYlMY6ryEG2LI3HWR1VB/u+MhbSugvkE1doZPg9Q5
QMJvk/RcOCdxMFg11ZHMozDePLEvpIbmp+zqUY1dFCEjd/1I5KlYMkSU0AYm
KJfj/NRHkcKeU+hc8TzhM+5T6UN6fR4152n2oz/U21FQsSPagjKHZugnzOxL
x3+4Uo7HHLZ7yzxvvAN9PAqff4cHPp7/e5MElzLL7E4L13CabkXgNFJRIO9i
9g/xTaLaYq2qU1DTzr0nKMg94lf4zcrpvdblAP01FB61OspLknmGI+q8xWVf
sB9R4f3t7AKx/tIjjUQsqaDBa3088Md/FjeSEfCTHMghEeDzGBme6wZMqCpK
urWk7RPh0m3hbHw2+FZXJhiu+v2c9w/1BLJnaLXhfBAGUt3hFxtbOfWRxsOO
wU1ZtWla9La362i+4pkRYZYkIznWb+yK6zdfybzPA2NH/cmi//OaanjAQIAo
JyWorlfxb+LcyZaDUPtgwO4ILYatz+gPoyDhEQKKFZOFsDC5UP8Hb7/ek6Md
3q7Q60akqNttp8lJQEe2UL0QjW/BTUIJh50EGmEDGEJqxWq78osFNoXo+DA0
MeSY3H2Y6UO5HB9Afdv7WrPYdO+EhzWP9+QBXHKix4cPEM5AFbAQCr7jDJok
1BnZUVa0aMdahJI2ChWQljh2shFTRLsBCzYuQ+QWKhilVa+R3e2t1eUcD6Hr
u5DaLJY1xchX/Ul08svkXtlE+yb3YsVB+B/H5VBC1SpNExURccssdeY6ouPp
/9FM1meaTO6kmBOUiqRFcq4t9nzmodD3QPD/aNsczlG+ZFePSTnO/QcQVowV
PC+HO35dPco4Mc1ekuk48UMQsYbels+0ec8a8gg+USQD3C0wRB5YkM/mZi8/
DiBIDiVUdDUljYYIJ6DylQezpb8EC1chRYShc6l6oXg9eDz6p0Un4elg2Xbt
ulml3hGoiPQ8ALCUVLi7ZkAnhTngefsruoStV+VMDFX+2fJEQM7CyuaPqR8k
c3Ka40i1wihufJsqZDXvh38e0YWwErhZFzEctFOqCaIOzbUpwXUbjIPjVq8m
nXZgvyPXu74YFBlq43gwYpbxj+sjztOfhYqxVFDJ9LFWfiJGRAklz7w1zbVs
QTOjeDc5SRqGk8e1OKyOq2zKQpfMR5PCtIRF4O+nVkZXAliQf2CMYQTjAGq3
D9yEoqu6LWobU1lgw3aqxvmSYIb7z7Xfx+RK1tLMhF+iScAhQZ51kqmhr2mi
WGmOHeXjf2hcSeonF3xTK5rb/mWscjVidsZ5Hv1ODKkAH0sTTIIdSq9IM78i
fgL9wueg77zS4qDMSFukKbreIjNDSoLwdnD4q3s6vpeFtdfezMRte0W5/6+o
zqRsq9PBcoipYjS7SlMvJY5PmKsaZkQ+oFPCVn/I5tg1WfeZEeB/30RRPwiC
WZcIMWIWnsdyZ56uT9/TnWUX4HQriPjMkw5KZe5nlSVom1ckktNBbwUvkGK1
uZZXAKLpNBtSPEEbARjO2g7FHRjqBvU2HY5kZZOHWOOukVdZitR62RnSmTD5
5EC0WMFX23UZyucnYI9oxAw6XfbFoe6ZbP7KAXyT9ox48VOp1qzAZZw9gMwU
uuBzuK7mhMEllgeyDoJL76tl40rHCMHlW4LPX3NL6VSJQrgPbqjuRxGLPVCq
1poK5SDugSTKgsI3cXdxsY07LkpPGNw8PTA5gP8ul2zXN7T/dg21/3/RXvKx
xuVKZBsZG+ixDC+qc8w1os93RTqogOGLD7QrAOSnkM5b00WAN5qRYM037A+m
M32FAoLAwMFZ1dmu65pi1EMyfMBf0EfN/R8GF88xFvwm4Tap2KSL9xQlEwG4
U0n1/uVYblqVS96par/6uE6e/adomnl+Twmac5PXesLJcvc2x1XRWJ9sAVnu
+eAMxoXZduOaZSa2b8XHHvTupsfbYCKN/WhVEtBS0Aa7NSZl9Ye4500i9KG+
BjRbUfQE/Vdhnr/5zfo61RFp02rEaIF7KOjSKuNYwJ5rm2DSDNNBTLvWc1+A
rm4EBRJXzzQmYIASjVOB1sDHdDa0EW8qfE0QSu43jO++SlzoH3TA/4xletQ1
gQqrEb/Usdo5liO8A8c0dCYY4SPNUgLhvdz2D2EnrTblwtzBMxcRa8NKnp+G
AJwH6zS6q/DVXJwGB4+eGuMvU7CGE9+b5aY6ahirNNag7Qs4/1e4j+dtm2SK
uLzjuv+Xkp2PF0M8m8Pa+u0ZH3dUfdg+LmIlpbXMsC2TItEOQyHKKb1as7Xb
3Us8McoZkAh5vmulcCkTM1LD2HKJ+wbhl3WwR9YxN9aW0aepeYk0E0YFwNpa
x64HKc/ZaXBUPTnPJpXLbHu6iLGvse8bWkNr0w76bdEZ5clDUcN5ULc4BuzD
cNsAcg4amxPbtj3nDWbyyRAr/7wmg+hrzUAN6JNmWmiKbm99RkUNazQ5Xsmh
On6HqgrqF5A621DgBPZ5j4ZPVZUZoRMyBS6dGQnMXYbeAj28ry5ZCCopDIIU
m6dO5tY1dM6TYIPWrI78ALegMott67Kl9q7duvKvnjPNrL/Wj61f4Qi/coZM
Z+vmxuK/MlyKLApoTLaqlYdxH5bgKp4q/idHVju25CdteBRN3Aynu+rVtCh1
1MOWChaPzL0DqX7N610MtxGBeDEomjZhkteDkRNwcHEjdkx8wE9RTyjYwC4N
aVrreaWrVKhqYFs+wCyhLAlGMorqSfdHjgghD+bQ1TshjKcmz5KAISGM2r95
6wYfEGrVBGGSKZyWuvQvdfL+yjty3kYvh1N67ur6b5whDj/ZlY445OQ0D0Be
n9OFGBwIWcRGIUJbUyMoYibx/3LuiUMllBbXrkNtu3XeuaRBYPVIYS+GbvaE
+dHnFM4qQMmqw3Dh+8RZNfrxnAaAR9UYrRPUKKGyKnoumK0RDYwwApmbiz8M
pqkPPr3KT8g97wiCnqFx61O8nH+pRKs88kmse/6pJ+FdcoNolJB7Wh6FtqkX
REO+N5GAfyGMi8XIUgaMyd5zgIQDAQoTg6BG6HkmiPyiAXT0lPHZlEviCJ+8
thiuQ5zc6Sy4PleyGzf4kV5W1nzrmu7qcGYNxIN8r0pGbqeMAsdr97/8szMx
uIOT4iFOpM3sEv6mWbnM6VZHZybN8k04VHJaITaDllDT9xquOKoepWGQhp6a
DDNNFuGDKGDL4/JMO3fBBYRrvDs1wLXBxlx3g/YWXDkCSlgd/Jp5Qr5blyJ6
jXWFMTbr7r5bEgudE+PUQ19clQ96LVOVxHNd22fcUXz2aijtgJVVb2CQnihe
NKGiXfYAQPECFcPX0zKNr5DETcsehOrKLDt3W3tLiTpdGiH2ue0QQ9riMviD
kUogup7hNIsc6FBVJTXWvJHw8Qszudc9JTvVkPwnsU+c4neio7GMpnWIevdZ
UQtKhrSQk55oCt8aoTW+2lOspdqr59LT5/pFZtWBrVvOhkBkgG5gWTlb8tg7
u33GmjtQZCHpfG4rP0P+92bfiViVaPu5PQCfsy5BtgMd3c7k+IUGw0DMfmWr
g4HR/UxtXyl1qruSdmQk1vBnEJVAwlD9kAbnSmkM/TzV4DLva8k7kref4Cji
974LK8zbS+SjORTCMTLJ5rpXHVfOUrNozHKaWXrKILwmaTAfQ4vJpheJHBq5
1m1cO/Qk0sfwInF6QwwK5/x32NA/hFTVNWRmyInrYXWFOcmiWyQczq/n26JI
BZ0e5DQ8mjpSv+MmmeH22M+tX8pkAIKYWRthCX/rs6gGHC66IRe2iiYxzKA8
G1eZEEsX0DH5aikal5bKeeZMEGdw/WLHVI9vgKHavTvY1Yj7aEUO0mmKvNeD
2k7BPcsdDRx1+RU9eAnlYTzesmBsE1Ry7Kc7ijsqDJ3cU/T14UUsstToTjqp
wropqcQfGt0e0kqrl2W4S8wP4YKXdmkHiuZ/s50H4nu0fsviKFg4xvK431gX
emQiYMGcUyvDJLcbWzR/1OlYILE/7hDGcbEc068LL9cnC/xg0kVhi541jmeT
ujjSHfiQDQY8KWV6heAVEwdPDDRnhpdottSB0tB2xGMVAN3+niVTJTidCQzw
4HLALH5S0mp0pXgs4vazmz8kN3/rvYu2PE6iP3RZeJmYQUMpfMjLtbDUYl42
qbPYY/uiE8IDG5SYUIcNWe1KppL4wC92HN7kSBWRN5LeLKgn/LGH45GRWC1e
9bMLFMdBHQitVMHh4ibN5AYTi+KZ/Fxoy0mlw36ZGEAAaxnQq3CS+u14gSA0
Fu6g3QA1PdKZwr+VMaJ9zSCX/wsWEJhSJHoWKxZlOHoBa7LlaomwWjNNH8Ij
V41Hqjw5xL7+dnTQk+YWqiPEboLCClpEbD7pI9kwoK7gzoUV2M9OysDQYtj1
MxIyxp4ZGN5FV1clbHzbSi6ftmTaItqPNhKPz2iiJNVGOhs0Mwprb306BVe3
Zqxe4+JHvHkZwlXJaVJ4hr/TSGmqQD6KGUiM/lTA01qaBv7VXyITYslzLYRC
YEDGp8FZq3/NqJV6W6hL25zCuC8fRCa4ifu2V12gv7tA45HgFyST+EQl/rdV
k88YaT6ulzMRXai0sVPsPbN6nm0xrRDaKNWgIyjzPDVhzVFrl4t56Uzj9Y6O
CILS/TDxT/qvDE1J9phPd203QjGuimKkAxh3J/JkbKcx3IFIFO92NIPtsnTt
+Bx4W08o7/4NW13AaXv62XrxTYP9hHpMDGhlX4DG1LGPQvdWK83KgytFhO4Y
VYTrQ3jr0rtta1Hn5rCvbwD5p+qAxMcqJv98RjHs++2+V3iy693V5LsEA5BR
+8ipFi7fk3duZDUQCzU4LJ6h+J8RNyWGeMCJ3KPrUuCRIKnlzQi+xoPgoyEe
1N+kXJcS/FI0084Z7X4mKbkU2PeJgit3AR6sygxy25x+uTGfcZWYix7Awhp6
pgz5g0fJieOXuG6u969ThMl5WAySd0zIVjMQy4kAEyKbPzz0Qau5tnHgU1hF
fyAuAzPoyvIYHQ+qlEVJa5qcmcRanUJpIMRpuZ5SC8JdPNptUbx5bvqhG5Xz
POxtTrWZ8PHfS05FXicGMgr9V75vkTHmqbc7h7PLtbrs+RSthknZNuCL6zW3
zVP/i6qXhQzIF+V8ZfEP2CFsYQL3Cj0yQwjlEp3qoCbzqbLzv2DMRd8OyQmN
cKyQxk8XjrHqpZJ+a9jjpy4juW/VHxB4vhor+/qZIXQdNv4Wo83IWzzgLtTz
VWGl9G4etc9JollZxelzS/OflkAM+kaUpRcdornxNlSE0fEuTHsrMx3SHura
AZiU4uh68XF6iXLX/CNWRncUjmBp8kfWY01B841TAVvcVpgyO0Pjbw3wp5qz
/pNieroIGXVHW52gkxbhR/7J+FPhnrXEalvbS6+NerpUOD51oMYWiKEJLhAB
g453+923NP0KhuAfXbZ+XjIYdNKAYJMSNRuEEKcauJge/32yJQm40Mh58mpv
YRN13ohG7DitiAYAKiPmQlRtQQCZe5AgOyzARplj7dupaImBicdpAESi1tQz
1FQhYbMx43DwvWSVwy/H81bRCUobMsGlzFccVya4fIFJ9XfGF/VATA3HfgUp
y3QLOauCSpgur5gK7gYr9CSVh/UHOC1nJuLXRy1o9sINNTnAFodSMbHoOPsQ
PDCVAGJChcKQspxEHr81IPlPG7RJtpGrRdycQJqa4fe2J9ZSMtb8UGkVrdZi
3BQfjKTh7k7d5g4hQv6Q6pdETLVnuA8zxx9jEjFK2B9dKdLKbfbXlaD9pz9V
pbTYop2jlJZW1UdbD+v2bEprw7eRYZl/O8kaeRnGO1ZtXlkHqe9l0JabDAZ6
BgHJNesbMQU5pGnfnaLHE1XTgCu/Cq6mB+JmenZeGqspCvjGDwCldgfqk1M8
c/BBEu7MMSve6tJBFCTjlrDuG4fzmLNWtGUa0+1i2y5RDk2OG7peCkwf9Ui2
XXm7FBJWU9sXx6GWDzZIQUk6fL019Laiq9VZr83VV3nEHH5o9WYuCsxjw0DF
oDECvro53D2JgCy5l+vU/wRKuUU9LQ/Js+5EKBIMXbtyCqFlJuyPyZCgPRpf
JpXXZ6Jcv60wmdgQdoCF8oe07Y/UC44V9mILntD4aZHyOfZRtBI6dkmmZp4F
UUuqY4+yN41nx67CxQ7vBUcrIdvZ28roZxBO+wyeqqmdi/9yOInbyFBrUTsw
21Nr/G2GsnDNPXWUAAYNehAdPpMRp/z0TmPUuXSc2YcfSUxhlpL8SLwAplKz
hzp+QHF+YnVE+OqbNMVtubUGYcdIjoZke6OiKrpiz9rwS9Ab5HvmZmCi5jyO
HX1gwdrRuqXutMIqbZyl0ZmS5vp+O/r3gNkmr+x7G0Ykm5sjHw7vf4GPnLT0
kmodWNYX4f58F+zphXmpuI9wNkArljMuyyoxaOjdVbijJe79bj5YTDLRzLvb
5/q8WPEozQoeCnSRjtc3pVsPLHVTBdPoWwkBhP4tL18jhOOjdIfBSDaH0qsA
3xdkAEzl2cWB0foCYuM6dES0/2AVRg5kjt88ZpiLJQig5AVF4EwZ3aj4jrgm
Syn5HsSRNKL3Fhc7O7nxzV7+M/8I5EYdLrIS15oSKKAPXxfAPLYo9XzAsTKt
AVFpidb2ky/lBfzbcWml2tgUXyLUVmN/Zigywc68BK+jj4YEHsKOa7eHBDeF
i/Y9XA0j7VpY5tWH8ry1TPMSLmCQT5kdK7yOnAkFnf28qKKqUuVn75Ez0zu/
PtbbyHJ6tP+JIK6Pf2FXw/i8pKl8V1SHlVhZQALHIENPgZkKkraDBYxajqvw
Vl/guPg9dJeMrYIs8tlrThNR3NNYim/vjZYg68Xr+yHd9tjuJ6FXSHo/23My
5NTgaHuwlHmVzBnnj7HpxW82Xs0h7O085f9X76FT751kA+qclZ85n0slqxxh
RXTLbFeJGGV+kKMF+z7cy+R7eHVzzeOZ0pRrVjmAMe+TqVnlDz53TluRYspS
XkPT6Uch3ft1vjg3iJJiwgUeQP+n1srI2AUuq8Lv9sj8cPFXb4yOEiXO2Yua
55B1gGcPxfDTiGpiNeulsEwuukr+BWZ1X/gWvPiWh1Dw70WDVVptUWWH/P/P
+j4LhuphR9l9XaN+JhhteCARZB0YLEv+LjMIw+SjQ2HGRXVy370j+3+ezRjo
jWgt88g/BB+uabYXueczjbEm9+1/Q3jO2p8Xz4uxeFhEasClybVNji8VPPkj
co9nzWlW1Kz1xqWtP2g70HPmeVErjVPcKKy8Yx3g710/MGxAlVE+rK5uy6bx
+AaqUDuMvKO1JBmTrrjiHlikRgI1kpOKaxPu8UTY3dpCj5HdKgiJHfTI0f/6
2CpsQ/ez8tbE7cGjt3tzab5y5ar6X6Lt63QlRm3f17tJV0k0wRK7OumBCm3c
24QYqo3YPZ84PQlwKvi0YoPsLp5koMH4nqeoJSMZdtwqk+FdtVjD3y214n4y
Jl2g/6/OfIwTmvSarkKHyJJfg1Ri3OeFyI+FkxntjwY4zKXQiMBIcGChzc1L
b3Xgm8/J4tI7mPqsuIV0uMbOvxaUKUcgJz5ZRcSYthzZuxgNabHdaOnjLEPG
X9FN4ZFi69ZLHgJ/yvaKzXPPlUJo/4Qa993urjAm88bTDQRC3uLdNDauC4Jw
zxaBvkpcVNtt4cocnkWEfuAvLLL1vnEe2uqf505qQX/nO0TRFgU8NBz5zCtV
/v54OYXr68czvdNvCBTD0/RDDwItqkRKCXiYbjXgX+5i7t/WkwohoDO39HKz
PIfQs14zw0ebQlvqOAauikMh7KF9530nIm0RON4wx6WBYOJvPu5DmDdM/F3b
vsA7+dkhdr+uUkprVD1vzVG7Wo9jGydDKh1nwzVRuZTAaZumIEFA9oImZXZL
G+pBH16rkr1c2RI/yLKYnwbhrs5KYHBlAx1Xs99IOCjxucYLs9tfSoavd2gN
EI/Cd4S1IMs24t6K65E2CDdbhdm6nYlNYkt2BwJux691ruwmUmLTVFMW9GMb
+PNaitbf5/Ux6quU5tzB0WEtMzY9gdhPFpSQbPFPZ29HXlGFpd6AsX3GeelK
YZBCvaNp/LUltIIc27W0wtYxlEEL3WahWmFdoEVVZGZpe08+mfsHGZYwAOI/
3vbYbgHAm1IZDt3e/g+xgPRCf6ekhPFaTh5CujEpnwD/rxrWAG9HFO0Ohu/c
lbHiI2Jg2L/xf2syKXc2Q5fdi3L8wsMUzEGxfds6RH6aRFAoPdq6Fg7BA21d
h8A9BxgkGxlb6MMgwBgutKo5XCP2082XfV3fUAROBxxn7BEz9xwRF3sNwwIo
oaMlPvlRToclruHjC6vP4lDUX7d1u2B5oLizUri+6IQKu/oL4q8IpDEHNy9W
rxyD0vbU27sPGLGmdTvi84Tyec+R9mgoG3Rw0deCzL7hp6M8hqXn1Or5kxQW
4Gwy3LBQPqpFevUdwBt06IWCmQDSERZvm53g+2j959rahGJyG8vTpQuyi9Zb
b4shv+0LLz8ghVP/7hwfZ6+12uqAmWPIslFWAKzA0TV2orsYKFKWHkyvbmOB
e0w70+/F9F6u637xaWq6wPNhxumE8tWebarTIxs+3KWIwj+O0giXR1wg4+mW
PKf3QLICIurVJ+qo3rp6f2fZX0V64rx1ZWeMvvtBVgtQIIPrd2V6Ne8hiIOQ
dnozDTLWIKBpt2Ftvpa5AE/Enato9xH80ezak949qi2cKi7ZdhCR4vmatHSt
JjB1ic4ZcGY+ElkjByVtKl9lALWegmdQNo6sm6WJ0NKN/CuqSNMxY8idHZ8g
8r2T9FScZVSAYONtIbqukdAkZiWUZcbC+hAUK1w2eIvuqWGB5imjdiHszm8p
DT7YtOxdwYoxw1PdvTpxobJ+ylR1QMCnwyURl7nHxZ++zIT2K/sdweYsZw7i
7udL2sbpwOkSVUL4IhMjtQo+FKeDMA2BEvdWXGDZ5CkURj79nGSnEGd4Kywa
lyFoAkAgicZdoBKUP3CGi31qWhUK73JWfjx4w/SViw2VCC7efdtOAvCOXzly
WB85pgGd9oBq6ZDlk6PbVhvjU3FPsr7KQQ7iOSu6man7CbilMaFZ3/C1lRpp
F3h2uZ9wkBtGNDB1B4aQLDwV9SmKzqDe9motLtSeVbUzLDcYtrMn/6QH0sFR
FJ8mZoc4bJwtQgIAwTCywCg/Wd557/Jki0B4cHURTpJ6FlWd6sELmOcM0Ida
G52+nY+U5ifhuCJndvU/O/LREuNA5Cmv1l5Qo4ema4r1k3kBCEQhZcG/2XXn
u6N9WJflRb4PUHHGcFXAhtk5C6wh3uVY+oNoLNsmKUuOHMAGRHOJU+g+ItOw
yWyZADXr9fUTkg15iv1eSbnr9VjL5IDNUNoOcc/D5XYSWC52rFCMDzvRBScA
sHLWY1D9GJurz5LWu9CK+VG9OZx4pinqLZfJAovPlUJXVcBaOIWSK5Ggt+yw
ZgspcXk5RVPaWQv4359Apd3W8X9KKhXGIim+ZzSoNwM+er5NpVDfoeukFhYA
GKDpx4GMJQQJ7QevrMuwUdNHImlbLd72AM1VKNfzAQF9Jxzl43S+FKz/9Uzg
cuOIHKRzy5uA/oOsTF9b6aZ9pm0PCLMnZIPzBlsPsCcoJRkPfZWogWZzMjCN
u2eX1A91sU3RLRv5y1E6e6/WwdNrNTl6ZHTbDqMJxzAHj2LdaeZvROdE+oon
JvEt+91cocbsfkqywhQtt0FcZt/ZnJ7CuTgMmKtnoP+/APSeuKldGlU5GEYY
K13N2MCvIZhQ5LKobke7K5nGCja01y749G0m7s5NvR+4PGBWK674mfRsQDlt
KIpl2FuY78hhdE0UiiNDJOo0TdwTxHBHOUqDjjqg+F6JeXX/8EIgTbC9ZDk6
R/e54GXLjFf17Oo0jYL+nh+OcENh1Vwt5JCZOo+vLkbSSpgqQt5e3m5whESs
rD9N6U76Y7BR3WdiDNt3+F3vRtbEgJwFIdY2llANCAH4kCuhnZGwzNf2wzk0
/O7LyHtcrSzhkA3SgOS8qnryjSAOHT0mOfUICLUBt65zE+lcE2m7hAvxlvGz
rfQcNu0Xgjsj2s0F2gXMYeMFlGreooGQL+xwwVQqhD6MlvjqgCRfe5DF82T3
I87Cp8vIxLCmEoWxukxhdgBDBZybtYwQbzBnsGMnMLCc91DaSlaQBvLgu4c/
KfhproL9kzkUpV+M4HtvulcJ8rMf3zopVYBYCoTO3ThJOR8j92WM7gkQfKSM
xjAjWCc8rj11l0NgUZEDHAHfkZJzVqlzGU8aeFlGqVddvmdvDFVBMQx1f+I4
iwcEw5uFP2dn2yTX9pyaksUXfUNvXmOUXvk3fW3jEIJVGm3UUFzygqfkWjIR
3bh/1YYPYT7Cjins+EtRwFHatbFo/oZN8ab8cXixciXMT1zFBZG4HwrgytKl
NANoa/i9yOC399a1uUV+aLpt1jvqsSiYGsZlhALrqgGFxyy+Tn7fbCqXZIEZ
IUe1XkIN4vpORdqpRzRFMBMi9k2KTrHFvgTkOuHVqEpvG8ueZzatpy9iLXXw
T5gHdUFrTD35Te4AYsu3J20t14ZjPjYW30+2ieYeC43WVXEWyx0ziEralJER
M0jAXPVrWmQ9z31vPtfFqiMFsOdX+x/EBKvoarLGWODSVO92W9rIc5a4qqXp
4hqgCB20+vudyIYZAX4/fzHhcGrc9WRXl4fEIrAOdFS9EtaPRni2dPFigGCn
oEizONn0tXfUDOUWZoqv4X+END5dHAA2zwKJhIw7AZ1gyVzI+S7hzVYfHjP5
gif6ePrUa+BxNxjSxUFkV6xLF3edBXo1HhzePffu97e3bN27w5t0MveCsBSM
y6M1xtJPzJ05BHMlLhIGPDlbQsGR9o/u92QPvMyB8lhix/3ZxlocTRVowAkZ
JjMp+3/aHrzK/qQZsWXnG2Q5KSN85sna1jXw1YN9o6X9Y6sM9vshZLUFiCXs
SkdN7d3K2g+dHPLeim3fjBq13DVD58XrN9C6mnrWQyd1tDMEQ2VqlfaE1GIu
B5/Ov/N9LtsSdYrEk4MzVELa9T30JQjFy7/mnFncYAAM/UH831jKy8/wUosg
ZpJJQreEWnbMYHaB/To4o1CYTziljT5Mf4iCqoZDBx65Cd++2ZmpbYQE8aoP
zABRjGmBIOQ0+YSZbhBe4KIinqFYIl2vFgOWCfybtNmRzXFTd+q0eou9h0rm
a7NZBA1pFQIcl0lekaiuYhIlH0QpxpF0oWGdoa73Vx3JF7S6Hzm+odAi9VbF
jxHxb07wJ9KLbpzGwCz2hONTgo9iIHrijVoJDW1YOuCoRZRu5ocQWKelko5y
HdAyjoRhuHcJOuIlVSdD0pIg2m9YKWy7kuUouiqRxzTqFJ/t6QoaxiOVN75u
RhZ5MXMtlc95zPWORJShzWzhRlQt3bfjtn+VSq19U0aoU/57d9yFVmroPaWv
9fsY3FlwICW1wqiF8IpyyCppjHz8RzZXqY5sUltywJr5FfOvT4dSlnhLUvqN
ZYhX+GN9wzjt5Nowq9gBkqv4yqPOfiUWE8tAC558kot8b2PGF/p4iAtsjIMS
eXVEO4SIrJigjzdaJ2UdMgl3HP7OzNXvXSW9G9OlUims8/tldqY24g6rTGbK
jfnQngjXg4gw+Sm2yl8gxKR6Z2jOXHQdV8tH37PF2KX7fzWmRDBuHQeB1mb/
IwyhQJj0U2pboLuGsjUxCa6YQe8WxpP3G+K3XV1LFeS1kAZnexW/4s+biQcX
8CSirwCQQ+eqhBRio0diRgKPUCjAooY5NKarut+i8hLKwZiYyO1arwni+mO2
PvZ5Q9mUi86akU9ikk8z8RMSV1nOQR3oo3qMrZ/YtDhPd7NfQiRcx5uom14R
G5Vn0UuV7Gmc505erXI0KNeK3hkb4qiCSaKBdEjAzOEF5UcOfLtig8Ru02Sc
g/eFydkXjrib2+IAByw1gY9GxmX4rUV+K65f8kcx5/Bkd8Fpfqi8LrAzY5hh
v/Bc9WjfgvAOiILpltAEb4I/xoFSUHIUJS70JdGHiMLXJuydWm+0mSywnqzw
/xi3/efBloyXO2OFL3R5m2yjOv9wQyg3TGa7nCtjuVMmVR/FExaLs34JqhTj
Y0taN9FyBRn8w5zN9x8RCPJO4JL1CDer2eQ+bXiC9NX/1FcJ3Lw03Kn0Unhy
LfuoiQ/zRTh8rqGY3G40M3QpcO1cHYVLxevjXJutoKcy0gdOyj8g0uccIaBd
dBcLhJkYUlrQzluGbQYxcpnmOMpGY6HEVTY7MA3Aeh2UMlyJUvq1qZP0fpSH
enJy0UGEayEV9jH08qW1xEfqtfLUagScuAgtwWYeeMH2A5Kxi2LznKSatteL
iJHhhYMMquU2nxoBGjPWNI/ST9cCnTN/Jb60De6gx1RhdNHDpPLqISBloful
0pSEgzXA8uRlYLdY/ujQeB4gg/XBARL1RDxX1wFWxI/2ohJxc9DBoR6gb3vX
dQJQLKi7jbYLAapTQDnyEWqsvMqhd5PoCvIBnkZugergx7iJVc247HYG77eG
pzdlBgDKW51w458ZILBdi2ga+b4W2t5ZBY/Xtyavjhu2U7jkzuy/CVYnuPm6
UkargRe6/slGjAImqd+v9N7Vxabzmt8GPniCvFLxY37v7JCuL1EbmG8OAuf8
tf4ICK5fIHlOGCPama5vca86jFwrmg+Pt5l6BBnXpajhpiCbgHn9mmD85j7b
XTeAqNBlIN2SmaxQybEa/vtYbst/YXn70MnfqJjnYhQutNtYv3mu4YFBQIOU
IbxeOcJoRN14uvMWhYpffrshLolQOeaSKuLv5JYPv6AKcpMle0TaPtU0pGF2
VTdCimJvAz9e5hqOa6Ab6U2T45yathtDSCLlh5YcMswICfuxukahtwadJQgv
XDjLJUGqXmLtHJCfJCUFALvRN4Caa7LA7ClTtiKyjsfncCuAvC8PRK1scdhM
T0Nfv58OcWHb7ZCyKKJncLpQg/uUcwpqux+6XlwoY1uD7WlrwML5yOqLhr6W
YZB8OZOVy9BAuCxMF/M+56FySNK4Jqd4PdfnHfbAkqr8uc9jDX6ZDXX/HDJW
34xejOfxOfCwFC90dCB+QCgichPVVodboa6xNyFbXeIIH4s/PirPjPRHJbyC
96hLnlAofdYcKkiqtybutwSt1QEeF7cAcTc6PAewielD9Zyp3zXObj53gdbQ
EL6fXD4Q/VgX6Cs2xo+CpyExeMnx9cuVeMREgXD89P/jBWXCP41h1PyMx4Cw
gKu+oXBDqgrfourRqPV5Sv7bEz2IlPWyjme41toV2xBG+VskjnDSKrxMfzO/
FapbfVX16H/tiEPZUdsVBA2T+CgIoRCn/hHrYOVYvT5jiNK5aODp0FDBLkMc
rw7Wyl/3gGAZMT8Qo+rYyh2hmBvdji4lsHxsCAXoho0B1xcIvVnpNCMVkGq7
+ItduXKiHdv9q3E6Hp6hgiakmpxwbpB6LA8hxbVrWy74rpKA7Gz98r8s50AD
omVenySczoBnv0kFKKfQrfM45lObhk1fTYUF48TTuduaf6ejQmeuhwm69GSu
kTYZ9yZbascaw+v3TmLngffnYsKvQyu2F7YovXrLswI501qEsKXwSWwM8w2M
ZZJaT3vQH5huxNRGxBy5tdxP2Hs0s6o6G+cuZmtvNxCJ2VyS/ll/DzAGe4/z
5o7gRpFt5kEybk9YvovDPFpRuJQnIv/GkDx7hJHKl2tH9dpZlwsiO9Dk5c8s
ycltFv1DVeyKUne4g753Rag85+mxEFuWOzwPt3DtI8vjyjE6Gx29005vtEeo
9o1rmwad0/jKiMaad7mRzDJaBNxHHgIZPjX6m0p8oxIC5DnwJD8KLcLILueW
k0etzDJ7EdDZNLQimuYU/iJh+etcq8PEgM7IlaUrPW+xHRMqohvAUREMmvvS
2Q389HXCjowFi5jgc2L412cYs3f7g1g3JIMW+0i9eJngoMNDPDA+6rX5WI7t
ct684UTNmJcsIpwjK86LIZtDVZ0R4L2D8S2plOs3QZNikJkPqM46YxQsnirC
RuZYgHXaerEztwFkBqE/j/yilfhny/SMj3nggo2XBr2C/N7DgjDSP+52Jk5B
G+TpGUx18e1KQOuS6/KFHO6aIeq3LtsNwE7j+KzTnicbvEYEr0meMkDEIQD0
MUXCgl3RJ7z6OE0M0pVieWG+DqV7F47hYlN3hy8ejcMBJhXiupRVIQ41sGrc
kGNTW16Cjaiw54WxeuO4bzaShhVT/bicqeAJ8d5OLw3DCMYNecBeCtIEAXQd
WQzTObTXHFOXhu/gRfjQjSUFWv+udny5mELAaDSDRAyFiR08MFWIQdCkxWQI
uryELtexaLeY7BBdzaPNexQv22cg7TOoIaHYHz47UMVkiDJ/Av9hYgQCc/Is
NId48u5hfqP1XTMsDtgtVKJToHrvAz1amXPUf78bC9N3aq+84yM2PXfImQZS
JjM9mX37fME4Dt1r1AIReGpK25wLTYuUOFYG9PwGS96KeKkpaCgE9WPslft/
T/fj9R9NwTdj7p3M3mwIf/U+VaMZK2UApfBj1Ape3bv5P2OOw+/xInSadImu
22L53gnIBOfdpoGtBeVMWElg8RtWd+ReFsNEi7anJKGYfjtw0K+UZkYWCkyY
VTqfJTqkDLu8rEg88Ns1m7oAZ5998Wv76oRxbmPPXzu2OauHSoYTPqNB3prr
E84Vd9MPjlVaznB8KLxwtttbETKW/A0eYr/FvSn6VMAw4nHv31yxpPrIe89U
fMGmkRN7USts8iN2uyxDrtCvCu3Uj/2c1LBFxwzFbsOEfsDtqOhXK8/d7qlx
hY66bl8w6vCxO+3OITd2+yTkyPFsAIl/7ApUYSVLqls1Y/DSSsDhI1uVeLrD
KuH4U6SQ/T4Ea3hmWRMYHiYLTziFSbX3SW0s5DCD7ZRWzzNaDHlwItD242OH
5lUaN/qnl6+3TDeDMQ+Ca8akTr0ForbOpLavWCB7SvKLhafl1Qy3MmFP118d
4+NhVLoBSZbaqRIfnPHZ1y+ZeeCX/vV2yxVHU9ZO8S4LQB92FzfH/mkCcmfm
Bn6Akw9qD589noBFDK7BQjz4Kb7M3+GSvVt9GbtsSY334Wyj7b7A7+ZYO5h7
wf6/Im1s5ndmHLOIrlvobFg5Lg+g1llP/+gg0lMPR52zOYqmXByFVNgfUjX3
KPeJWYjs/sOmYnNPXivTxMUE/+Kz7JK3QDtC68WxD3L1x7wWxTj2ccQRh8mJ
KVH+7jBYU/xpayYMXr5AVo6azkYyIrZaAVn8qf0AIXaP2agbvQXa4tF1if7U
hLvWcWwK9llxcClyMpJQF8QKAHlADNNtRqCWw1/2IcVWkxMwYcX/VN4yg/9N
Acuqq4dkreB4i8P17X8FE9PPtUjlFbp8SdXLP5H6DMNAj6xFDkzEo4tYl8Qp
uHZ5BbKwSzaC0fxqEB4E02ondKsz7C6mNM7Na5Wpn64Oyrq5vSaSFdzqPpk4
m2KBAekjJFrfqJXjzJlNbqyeHaT3eah/wDICm4yNtmJ2fYdazdzhYJ+Z/Qo9
oTBPa184jn12GtEu656IYclUQEX3rfVZ0/0YI5wI4HElKnyF5Kx2ztRESnia
TtXcJrQHblcF/Lr5L+i7tws+DpPiTh5zR9/Aq+nMrHRwfMrhLvPxbid9Vig9
ZGnAKPqf0fMYOD/wsjdZ1Ydt+HzpvN4raA21w/1X6zWAWkBHAqA63ieWoe6f
9+Gt/YF2kO8MK6PEw+KeQRsj5h9AWQbp3Ezz0BnI445tV8T+BXufUbvnn701
h0Qc32YKtkCKlHxrqhXoyqc2YBW3pzHdLnYJC8uPEnLyK2Axdzc0DHjnxFcb
L4WQJzTBCp9ANqGQDfLAJDB1KaCwdiAjekTJJ76aMQl4yRrxCnd7uQGB+3pc
+MM+/uIS+WbD11p4uALiKup+kzPoo/2f5WURMBTkOU79VvgcjQXyRwEakF3d
xprfex3ZvepJIfXVnPvuZGkoGwd/IDTHY8Qi4KnGlU4AiGAAukUMPHzr+pK9
lR3TGIJGskqRD2MeDM0fOml9wHPMW+2q3X3z4y25fMv8qMnLWCuo2zdGPakC
N5VN4zTaJ4hdIy+FDf27hA93GIwJ6rV232xWUxK4yjtq73G0Col0M0p14rjq
dp0iUWf7+K/6pad15vJIr2w7mjy9GqvUbCRbzHzld16T8nTdLxb9hoCXJ/Si
u6DXVchsLPRvzw6Hc7cwLgJVkdGqaStf0r8gyOkHbwHxbkIKuzNLNN4RckQk
AHM+6f0TtZE3SBA1UzjArIl9Lu+R2iG4OED0CBDya7iHHBLmspYpndlZRTvU
wQgqeWsloBzLIErOvPpDngsCH9e5nHUJ+//YmW97ood2fv1jBnqp9iMJ1L0I
R0IfLnNuooKxfSx6iOYMnCXHDLAqvxjncMDv9MNw9HfXnpLChOznbVkAIKeC
P3YwcXjfJTZDUxQ5n9ZKhA5j3NAhZDSajfIxk9DzReZlBRwthOQFv2vKDQiN
fzIZBqJeDBxdpTzh98/B3U18vywS0bXseT2jB3bBClK7hQQTv761jxqimBa0
ZPwexLJNzmfdhrcS27DFdhV/xVjea8zOjT02U7Er6EQhL2pfXxDkKUDMZbG9
978ZJSZXGZpa7wlCI8dHiUKHOktfd+UadcqNxwP0gr4SrzXmydUcuvFoiiOJ
ZEsiETyFklZW08EgGwKP6G2jC5vPtQAgyioZia5KTXoJA7v26OMBK6VTHpB/
AqGLyYKEkNsCLxzZi91UcG8DUAXSivRW8WYsc6spxnjjCJEAwXcz4W9UX+Ls
BwPE99zXz5n/3Q8lPOPZOsCqM1jDkBcLQNJYtF2t0L1KtKCBDCjruR8Q9819
gFhdrDamX3qSbIxNQK2PKoJFrLKzLUXrst3B+gT1QVslzLLBtktH18pK6KRq
rGlfGtknZh2mP4ZXBawFZ5IXeufC4F/ScT3T5Fql7Ok6LJd5UMypnMHQXRWB
3bx/GrV6+Q05b58IoCLzRsiA4GVgPX2FDsWEBdziqV+ZRKlsp58LxO+N5D+/
oQNnfcVE497jbus6ZunrAi5B4ig9de4eDHpOhznZVFqjzzkMXpO6WmwKhXcK
1WaFMM4N/X4qlyjoIagWmKW6Z2COtRppJ9HISGYjQXNhQKrFu3auoCusx8KA
DINN3qS47O085dFJRVna4YizqtFsSpOVkYDZQe98QrZu/yxcAhP4hZyKizLQ
3vQXRUh/8O0Wvc9aOoRXx3ApVK1s8P2k/QxldlBvEF5tyAGWo+D+uyimK9/f
3IvKN3siVXGSWdPHmslpE4sqCXHPXqQj1Z+R1n2zJ3RKIfWDxbe2Uoo6IcvO
e2kku4X9o15buI2eroPIs7Clnc8gXcJRHoM8cofHi7YVy8ZrOz9jrFzwBdGt
KpIR3Q6FjfctD/9NvG9zpXxXex4wXoyA/b0mc9ctGb8qPb+EQjHkZDlyrasA
9FZHHIFVS+BycQtpZwWf9avDwDenQdLimmIqtm/g7+zcs/vmW8jRjLKrpJjL
4FvWU0Z6IYM47MEzytxCEDDxZf7CENhKGBt8l+pkyVCSy0JswSOGEnoV6YPA
VyuXS3QAWi760vJlZxVOcGGBj8a/T0x27bCXhe9e0qz7O743CinBb5Y6AeEa
rIZtsO4FHde1zO2b6N/8dQ5HCMt6KMaXrHg+b2J1sVeRKaTqHktO66fDL5k8
HEGgJH+7K98dd2fOHy84Sc9TZjbvGwOxrKWobW6s5MeE1zISGNzh38sCkO7R
iRnl2F5Imirzpl8oprwXxlIJ1OJa1y37oxoPvxbMqqUpxjoLk8CaLedhMuWx
Se295bPU3sIBpcAQK7QoWWw0/4A2bLHDghQ9XYWVEuJhw54KavcJbRKB1GSh
UB3ZyqmlxuXsjDjyQMiXNbkjaK89QqCmsmvMN7HGOKiPr8XXsqC4pn2Qps3y
NggguljWHtcRpu78a0MBLUjOlHohri0FZR3xZrTxAaTS/zhWKQwlahBVe7Nz
g0MPDB9AgrOue/Vk6PInACdHK6ljE+Y5fDlGblnOj1nzgmLcafZycUM8RtYv
yAdgR1YwLDz+CCXYwlCPetJeUn6WcYisLIehFMB6BwWps3Nk4xlmH/uWuN+g
OmhgBCpvCM9JqP40OwvybNA6wPpMf4h7SamOJErryzrZR+NNbxkstFJaX2cy
3/rOaBGEZjKCS9be2X+jFFVUoRrSFXOONyrlohM20XXm17JvaiOkjeFwHgtU
sSBCrmTz1kW0Z106BMlDuFXXhLS9tVXXiLFbtFpN5iafucufjT2adR+y7uKL
6RqpwmCYZ3SOzuUn7iWxB4T1ueg84Odt2EKG+j03J9gUMEiBILMP+SQl8dIn
QE8sOZcUtJPEUFkh4InbQujHU95yIV63BRe4UEQWhG7ec55SbdlLz9yJThCK
1ov0yyZvoNMMQej7OCYB9acwcmIukB6CAHm15KxN2w31BjwW8wfollM4OAYE
ecTT1Xp3f708+KRCvZCOs0H8r2g4t+MVVQhj3/8OaW8XcCPOa46d8D+UgR0a
kj4zVKGDT5dbA2ssUJmG+dteqvKcHVVGSnLibNWmqIyum2QwyHoV3+egL21I
GNsl8YgkvxFmm+zI4D6jtNZypmRmo5GOgNUW4EiH7WqzaiEWhNWiiUtb1vfu
H+NwkOzaoUB8NI/eipqqTBEmm0FErw08/aihP2xS+AFDjhxUsZyDZQ0vKGPk
cFl8oseCDaD9zS1gkt4qwybE6ZIaMQ6C6DPordzYG4fii582PRRsFuU740+w
wcDFDZ+QeydCS6EitdLgy2VQRJkB3y2lBkwpnWa23xiMaJYBUEF4DbjIN9zV
xFT4qpuwVRxBylpDxERG48TJKBvrWiKWjdVm5nqoHCT28V/w4U2eXXy/H4E3
hECsMcGaDFZQgbwyVHCWbFdw1CcBh/7tP+rSx3IWJ6h1nobNenIIqWnACPD2
9BFPF3lVR1bSF+REhzuH9xNsl45ECuie6Z47Cl1jT1GAVzjQBEssUrsXuDb+
yXfULwq9gvJQhs5nA+Drq0YoOgfDWujRyyecpkCUrfM9B9z8Qsy4FJdd8hFw
oSBjjMQhpOK+4dRKHZVh5x4l3AKBXBvfOd5VrBA7pv2in+A8PbNv5Zvca+K4
/tvUI7YB2XZzwpVTbldofcGJLjwyVeAP9efkZBboN+lpG/Ov4E6UlBF6plc6
ec7eS67R33YTG7m8OhSyzjaiS+z6FzS/+1pBwFG3451iSveCjq7kjRJlRkP4
UPotVbksjGmwp1QeEhurjiTsm95LXRrYzmmm5uNvEwxKEqlSFNLY2iK5YW6T
zQsq98PrENFVRM+JonleNvPppzj7SL9UN1gAHDjndlJJh1Tvy3Em7IjSxNKX
HPIwpB0v5ZrmbSHOVKyUk/t9QjH5vJDQJiyy9i7P+0L5lqVRhaWThxvjLSeG
DHvaPcVSe8dRGBWQrYDINcgM4EeU9b1b8a0h0t5mupe0cRtYSqNKyvJQTIr3
2mjBIPYYs/Tkj8T2pACD8q8Zwx0OqNYp9PCR8I0TmD7HByFV49zdkI/uvs4n
kj9jFZC6TLM2ZXOYHcsDLXknmuDSFOZVnuP8VLbbNVArBqAFG99BxLI2ULdP
2OtHg3AcQxB3HPKHXsVEo1nVp+EYL+LuCrkmjuriONYPmbOKkRAiP6l8/03V
S+gk8AmHsUKKnbSWjDIbS8j8DjTuGn/pVyl5/marwwiGkiYOWqhKeM6bH+Jn
ItkSLjnIE3MtxOCHv3Nry1lME6i40aIlRdBlyPcYreQxcNs7aH1gYVH1bEkT
8+OFYulcCagQTKtmdnEG5AA/IQumZau4a32AgY0LrZIh5CzU2yk5Os8rDkR9
E+P1DroyGtyyHLQo7KJZSZV7UlqbPnkklSJ8ZwrOLpp37GAdjihxNj5wpUh3
DMvdG/bHYfkvb8BEsHKjV6yBGBmi9sJdnhGKhp2dAtN3A3zZE/ps3SMnTIFF
zf7WA2flqwnp/Gg8mrQgQ9T+SyaXGOPY0O4IA7F50jDlWeuuhUcV8ikXlQ51
DqRN1B/uamhWtPPYJ+5ig6088gAAMRNSZw+npqK9CDNAshoPnoU2/9PeC1h8
iOd01JHHW7+c1+38iUEtxYFWeaMBbDBZZyiGWpoI7rdGcWO7URIEq1S3X6Da
/ckXeR1wqvDsh/TrrgXpDYozblq1BLlr2r5ljKtDoFIqfDoZYr8NX6wNyLvH
gF8X2Vx/SEkPRUUqpBKqTIg/uDU+2BSG9rBVTsub6wa2p6PWHwhsXJgq7yhS
eY65y8wSnTIB8kWlX92PcDRuZdn6jhMG/zGtJvh+Xl3x0P5/tzHoFhjrCGYV
IAxnuu6FoLDsT1T0UjU9jgNNQkskSWGbpef/N7sgvVBkFQUlEmHZ1BSqyPEH
SZ8CY/Y9fDdzNNiFU9sRsDkq3XNFlxUnMepEHtGzd/H4lEf84BfW5LNiWlM0
GwKidTVhG7f16NJ1ODf25/E+v8tMMrBlHBdQfYx688nzUdFwi+KyMbW7LjYr
n9Yl4PW2ucOw4931R5C6oMqELxB6xkEh+j+UJojnKvYBL835ADfqUo7h4xLA
rN2kaQrlcRU5LT+aVp0/0NUdkYhVtz/j5aZlKm0Ni91FaIQSe8BDYDKmXAzI
AkHL7vAjQwNiPPrjarykvjbV+GgRoHvyn2pLS2jW8HGeLUAWavNDyYkk7znl
GVinphka2rZvwCT5k594RKAPfHMAcEXmcl7Rc7/KeYgCyhA8Eiz9KA4yccQL
gSGlYd2f6LZ38OgCjswlkz8l+WGy3/zaK6cIL0z96C5QbgyBrAar2B69Te95
yY6wCE/YIsBDAJ35c9Prn8sA13OkSIT9YmBs+5UJdw5cbPJhEYyres8Jn0lP
cDT/GVIEYBOGzQNkB7CNwyyrRkZWC4jCn6kHoAt63c/9dQdcvFl+HePc0LO9
lj/GuIFUOJC82wyKujSTsQi4wTT/vuxou9eBEw4mX1544tMQdBTRxWIZU+K8
g/gyuMkWlI15fnOYvMYgs3Fm88wjgYmyqC7O+D7HMLTGreXu55buyWCT3ZAl
gvbKhl3uE3K4Tj171II3hMD5Bs425LU/LJ70XlWATnATu6uo7pCu2fodAY+L
TXwepqWXuMeLFoB3ra1xjCxTu2PRdMCPXkSf1g7sbCm2PXVWbBq2HjPJcXm5
cm6FG9XF+C2Mz0RyC0mFqp9w8DBvJkfslsNmK32uvi9Gd4cvGK+5w3q4VkGh
pOxOMB2DJkrnPMuFQMAwnE9wdg/UpGXa9sj6SwiMSE6W2QxXuam4Zf9K85JP
CRU/npuxWuvufKaiDmowPpivhiwDTVhL/SnDUv52pdfP8ZCERuakrjXHDq0n
TQeSCll/2qzU3KjMNrzc5DDry49w2fc00G83cqfucze8pGv2ndK2+hl9mNGU
RZ9SR8h4M0T3bsTJM2Z2OcwLujupg9zzjDXJHKmB5OKZYetWVpN+6S4sGvvP
UBD+XuuTuWgltuqRDZSTW8H0REPK5Nb4U2FpYDtqqnFOOSEyntYM7eTp+Eap
guAsMCidW2ID/j1i63D0A1a7MCvUDVCFxr8gpLAgO4ZsiaP4xgE/cDt6budX
6ZFRRr3YcjFxRJuJMJp35SQ3fz++FT1vUxsPp6nAk9KT/5RqrDXM2DTPrziH
N5Fg9R9xXkEcmp4CwnjEjvQc1HrInDMyI5p9wRfp7PkOE0ydQMZUyM/NjRuK
GDUavbCYu/6R6U1de0IBEDypUJMO+Jeko29KHS/1rrROoXF/jClNqcIqZQqq
NC3cREbpRho/HV/DxBCY7ewivD+s8JOfsUVWMYvlNvrlvGiSqboEW/Mu+Lti
9bO4rKzggvI8sprGZHzpPi63rLzmrS3BNih7A3kCs6a0U/Eq9tGEJ7eUG2fe
VW7Nz+x3s3fplJQnQYjEzAGXYMBWwhWx7x1c5R7uvRwdRLbzmjG1gnVEqi5x
k85efWVQbL/lO6VMFjgxfdZTbIH7FXEDsEPstT8lmILqyIjptb/kHDT85z99
lxuXOGnrlCDf7f1e8XuFLDnNIffN/XwBlXuA4658M2ZXKzOXGfgNtvhisi7a
ZxgkpFjZ+M4tv0im/KwePVL03BgYovkW7oNos1Bqm3QSQhVamJa5JmUhnDZu
dhX/jphTrq2tDRAkYYrqh2pB7ts2uyP35AQgI1hD2T/+Es3cUArQZUEXyF0h
B6APUPPQoiYzvIGvwAs6/xX3ecmv/RLmrXd82OvDGGckjRmEpxcmT2IyBQRq
hXqmWdMx0ATPhbBlU6pRtiNKwDULc/rh8SjlC1gux4CCgI6mTWkmlZzsQ8d4
J1vBXHji3XXZDphKmJL1muBZ7qoWZX3yENLO+IAQRI5W/TKICySurptZYJh7
jxbNj6TVWKJkrx4+KgEwlKkbZ25ykjlSoHZBX1XKfXM1voBNfdTCCXsMbAhX
5ahno5HT4HPwO+cUoRAV7VGnetrJ+gD6/Za+81E2pXYYrFKxtgVipFiKJdar
oWBKnKEcB5iVL+HzL3xbcABD57czdvmjqMwuu/l8IRY2fMqBCMQ5vGSr/zNh
iRIbdZWmNay2Vs6KeiBdlq6ljfiYqdmV2hjvBTFjW6mMENA7E7KNOlrAGYiT
tC5d+ipsywbB5SDOt3AMquAtckFKraVxZjj4BignV05I7uhjkERyPw+G+D1L
2pzHL/Q4wfZjrW4vVR3LE6WD9V9rjeUKTm104qjXDqy+dNu4HmCOEGuVDwPi
fcuS56PHgRyPMEokhWvVZDbOr1aXBZiq+M32flntfxh0ab+IwYh5YyPi0bgr
txKyCcXITft87SK7ydryJZPdaDdqaSFdfB4xRyP6O7qmM5vb6T+gXytVDkoS
q1n+KJ445L9/E+jZd+msgqiJfBemkDx3fJ/eks4Rk+/GGhermNcBIp6d4xd2
zE/RoPLWHAgYl+gTIp2F2wpCCtZzQmHCip+Ix/RwEBVUd4M2VcLSq/v1LYv7
jyUbfGg79L6addwLwESKivldFiEA4gSoMKxAnz9alUxkhhPqDKM2/31p8rFd
BX7zLfFBuCNBidqcUkdgMKC6utFm4TgvVqNcEDVAmh0uUWU2pUwCIscECQVq
HcL4Ob1RM7OvHxYBV5dqT44vRixoncC3/190V6cJ60/AdRcB3V2F3swL8+j3
j2vgZbnj/kn+mAC8W50hsIZODfbyZfH2aqu6OuWPBLAL3HWw+uNIyp+/ityX
EQhx+bUtOjnBL3HGjE5gYW4ydfD5ABMzodzLUwbDSOqNOaXPOboFM9O9LbJA
Mud+s7qO8Hf97DyM3pGwKAfNWtJUwU7tK/AzVKrqZxd9L92/ufNTxM7QKQk3
9Cz+b9K375UBh+tOlw71MRqgzTsqH/REm+YmAwFu0CNU7eZAwbLbn50HOgZm
WGC3SUFuj4HGKzSD5JFrImOj9WE2MeeaKate2NFRAwea8hx7iYrk/GJjNIEy
ALkgPwbXWq1BDKOdZL2b+4g+fonaeuy534TFfNwI/ZPzA9ukX8HeCSkqwaTv
LFob+gAK0+nrFwwlZ7pFrbtwOx0KfEk0Sbl56kcSiDyKHxRwJFgG+2rug0qN
dPKZA/Ri6gFWcH84pFzbgNn9rPJ4pTLzTQTttosLirhCzN9BvVhU+HkfA6GE
JrCzBMPpptvVul50ofrHTXcZQu4bLaayotPjmVcN+mcdgwAgsfqlm28UT/DB
vY3v3gEA3lbl/L2PlWQUulgTf8216prho8VWUiGPMStjpjfnJl//5Kyi+soP
HQIbmyKdhI5/90c7iAPzFHex7ZUxQ0ugJAZKO5TPExGbYA3fwQlfjuKuQvIa
fN3PSqDPZ/0jqP4zKyWpOBzTuaiYB3FMdVj+dz90WLiTKZ5k0PiO3/b/dML9
wm5+FWqi+vP9A0c9cR0lGPXvcilTXuRUghTZbjhSQEpOeF/WZPGQ3n5hkKdr
wspRxAx/m2q5UhcGQfc8YEBf9wZXlyp6dLvKgxTEGPIQeH6HXwam3kqUVZLI
x6iAesURj8BoJ/palY5bA/5/PhL5b9ek8WS+fciV1vfanTncvNK8evvyLYoK
apbMWPqX9Ji5pXbL0u2I0reWGjGMjrsQlvv6O+spkPSoYWlaChpElLBcEGjP
kk1N/0wdNLvyiwRu/zkS8E4sSzmWLO0Ppql/9ow4PC9QeS87HCwdGXT27NTm
ISFZkACCpyLpx2BUTukWrQIoDM2exiTnRpwN+vDuyPbNu8WJHu3Hb9IMbLOx
H/dNTbhflpNokwrY/NL9bIgiB7rASP0Uyu147coyCsMZwQqMn1HH8DkkYPZj
7wrFrkGmoNRM6Wxrvf9qJQDSuy4ZfV7e879QeZcZK1y9MM7VTgHpm8jirrqZ
NRx1rvvsvqONpfVSKULsuUwOotVewnOZ1HHf4mY6RQo7dXgb7cBJnRJ/bxGH
j/l8WBtvxmUXMr6d3Vxis5SK3FuLbkFZNBr9GN6Ad6vYdnS5y2+LDbnnKW7O
lywyLCA4eHGghKNryKvbkui0vQ5bRIw1Xj/HwoRlUckdTCkBj50YuGyo+Yjd
VLHxQy/N1R1zY7fCpVb2qGnR11HIrNpdLX0T3J5bSdl0+oWoTed6p9TXYAaQ
jL9BLgIhef+091MIIFAmI1PAuSsXAhA4wRoLEcp+Nm940YrPZTCMtbCk/cyq
EDaMvDBr++VifAk77YZORbJB3VpMAKnK525hcz2O/OcKg8BrVx0/ziVQnriF
u+mdqnrJ0tYv7Fcyq5btTEJ4ktI9hFxcmR2Z1kCyl4lIRHp7EpqyqvwORMIO
6bw2iOiPoiQ0N/PbMlRjDKEZImi30NAXcdzNAw0qfA7K6YGbpW71PE9dtmCb
MxF37wwTsef9inEbqHks3/+MsssdB1LTA3uooeVUfKd/vzTZ4BrXCp7pPjTS
Kr+9+usLe9/wHg8q9wbk/SI+H+C7swmbIHiw8WbrpXOsr90v0sbhxIqyBiAu
VEmGgyVGtHJvok0VgIH4JTIbCkOOzDjJocymbJKBymVOG50g6Bmv1Q6ROSNa
eXf5j7c2U4zzrhyYAF+k3kRUDjvtxnc0ugGdQVHTpm7h5U/PDBWcnst/s/LG
HoXzmfPDOHsQlsliN1F2HFB8LV1F+cZNGL5qNlrtcVdcW8d933TlGUj5aAdn
YSWeUnC0C9Vz1446oy39Hs3qxF04gmJXr+Cu6fRvwwRFTFICfaJyA4x2rf33
zs6+RIatNBoqlx5jVGfwJyrIzR/lvhezv3vt4NjRxPcp+TGaDdWZ1budwboM
DMjNmEIhvKOs4Zd4Js++KjekdVRtbBTNBApUbujS9fN8VHjUu38mIgfw11hZ
aEpYIMm0PHnQw4zgn9CpSRjVPysP4ZhXO5vQzLe3ysj9cR/upqzGeMczN6xO
WxXvoy+lMh5cy3VaDB3M4/EQjqjSJrJPtkFbB1Ue/HGZN/4Rb9m7PJckaH4T
x+Qxqvc/4xqvrYjKmrGYo1EcOE96+33VvQiA9gaY8jwjnUOiylDj4LwfIP34
9XWZ7dYUxaiTejXLe7wbvv9Ag8UNYOqOLaP+n7w4gMzAjEKWUOrhsU/I/CvH
QyPHlj6hsmRB47v7lszWVmC8MTffT4NRorB615k0k3bSgEH2J97M+3SVOezE
bJRONxcOgN71Vh3Mmb/Smh9OFiumSKOdgmP3Lp9gaaP9PajjOqyXnVjBxWwU
LhtayfqexnqA6uejUbu2RjoPlM6YXBSL/tGILfWjF6jmdeo9KfG+z0J0771n
o6B879KLSz3zAcwM/KqVB3iwM8VcsIqheZUwsAVjAoOmZWLLbKNIMcM9jyUh
a5kselN7xhIKJ83/9gbZenskyYwfLGGbYfhP0+Dyz/YpjUipW3R775V+VpEr
nI1NzL6WTLFkakg5EyMgTajPgJD472eI+XDQ4NRrRHibGm5XlkYh27UBoOyI
OlebR7pFFCM5Zz9tOjE11+9cXddjq0SOCo6PMa02x2mEVqu3vWStZSssAAGc
KtIgMNxpdTCNll+9KPpOfGbPCde23M94P5AfwI6xgdk3rxFqswxVcqNLdJ7s
0Ba3HHxrL3bMVS5YvE/3Xxx3sepbDbFNWdptsvWRmLfVbV/BRlaElSBmwUXb
IEoksPibqlOqxOPMCMwoTmICCbCLXZfVmDwTiPj37KFyM3JRobZbCnxtybjQ
yeZdxAM3Bm3BmFK0UbMqkVSmRxaMyZrtb7cYMFvT/LPASUr76ZvKgLwIFlOT
O3ok9ewY69/59UuAH7DQjlhBShLlH1OGvAXW7Fpx/Uq/QHiTo9ySu1lh+E+t
XP6f0frsqocPLuewp4u3EzMzZivhbYDsmwqZoOPMj9bD3vV68BFMAsR1DCdx
0fW+0TxQliff61OxYLWW5AFpboPNFm4KF9G5jJPQ7UI+FCJuONFlC/SSXsBX
cDBQmMJ2ViOnbX96+KIIGtbVJErKqsrEsB1CzwHT7/bZpq2U8gkONtaoFMub
aHGqq+ATzOz+wfaRqA2+6eQJVixcGJHac5Jz2+1TW2cB5T6K5/IFRnUjjTah
RhcOpdxB3rnzm9Ljf5SpyOepOTfhYbWD8gKRaf7IZCv2NzxVvltDX11LREEm
OJmjoV92BzgMyOJctFHQL8ZcV7pE0ez+wj+fnxMPo2EaXz/aCGHqnTE7Xps6
UhzPT1rAA/HXrEakl41B2fuLNkT1OgtyQqrFw4gekHsWAI4XSB1bWjG8FZOw
oEABxHbB8gmM/aI0PzzavK8FZVWWdXQ6D/ACBi0ZuH1ya/XyMHP4/5tbMW6O
x+kUYlopuly1ORjXceRpVUVyX9KHw32Mg+fIvTVc9zaJmbBueiqujOMHa3CR
6XUjOFLxAqFi7VB9o0F9a/dQDgrxTaN7Wpa4PZXcoO562FYKa7j3U/sQ/y1P
JNP/7zMm/m3GUN0cjcfdkCX4PvNq6TQXqvuCM8QR9wrpwYUWNKMqITPOLbm3
ytcGWn4jwCmE14j8f60enBNTlt93GYeBersH0AaRSxNRXiSD0CvUz6STVYls
gX3hw72bgWNWjWVa2JQlgOwLT4q4nCMPcmBHSOZqxCvzsnyjtOj8oImkt9eO
ugKvnnuIBx6THXevR9gpNe9uczWjJRm+GaLcmUyzuvOyuy0NN3FTOeY86WTv
cOjXK+0nRebvbBOaWCRFq9PM6Pgh3iOoZDT5JV46+ts8l/D/dKzFnMCSaOKD
jAnqykBXvneahTP2KvK6GSotMEX8kl7bIlUqnA7pgD1sFeoayXgvJ6mjTZMW
4IQjxUAHc/WsB6oSY9UzyuJ2uMNqe6HL+Sa9MDvu/cp94BwBxpl4CYysGF3n
O9pufglUXsDyHECrs7VCX18HUSBfeZczb+tImwnzotV6FSoHNuQvYgstZOF9
v1+aRDdmRDfJg/eYAyTa+b6RaY9icdjhcMKyD2w/1SzO4wnVkqdeJOEW5c73
6+GxJOxBVEoXWkJcGceNxaONU6ueRgkU5VAOO9TQgD5nu47EksnKzFofxs7a
HCTBPUl0QKLBp7yj7imoRODeQqE/14MFbjNIj+Yy3lRWjVwCdU5xlhyWqaWV
kOatu+noDaTYaAl7veKM5gWN8RHubGOo/YGrlO27j3hf22tOU0dSnL3fr5MK
ZNE4MnHxpcYv2mnugNNvcQeFMxMmwovG6qW20QHRv2oNm53qcDwhlmnyv+IA
vIEnU0LqIynlb4mPSQJACMurvqcuvKRrZeWv9F2p1pBsyVZit5nHXqCFb0qb
mt4XmGjgcHRrCVKziETzTUtjJMR5c7WVvzg8upzllsdavnlNpc620HB725K+
Oy1PvxbrHoXNnhqg+7kWZpnNTj/D5V8FP+lgU91eiROCg7NL1EjAYILjqzL4
g10QscXkn8SJBLUEq0xqGNQ8pKzOOVn88n6pt/5EA4VWzgacx7NtSdxU7dcU
huXdVcksIMXuQktPWWqFJTA2zLpOSFQHUa1MDH6VWT1gm9nscBIikDauaSO6
RHMonN42DB8wbxPvsOWRhb+Gb2cP9Lyex5uCWxF6KVFDakeN4Wm4X2DC2tfu
b0Mbjg3wL58lmV9Imsxjzo4IYRGD8TQqBcNJMfLVmpDW7341ThVICgrEFAqJ
r2jJFMPjjNX35//efrtPOvL6Pz8+rKVLicAz2GgWLbKWvGAJHRCLOQ1pRdyf
VDn+SIG4tzR1XNljbVQV9qI7BC4MWYPXoy0DvMj/AGEVlmPRXdnYkVJvHuvi
FzVfXjleDUurQktm8TO/ogfXu3WrAX10mEctUuq19NOBpBd1TdljounRP29A
pL05fOgBNktsPlJEaJhmOoSoB2cDE5+Kb/Bo3FTRv4gSZKDZbQCpBEaW24sw
IJOO+isaE4iw1Ud2zGBIHGipQcKnlM0F0EL4rPZdCXdZN9whsQwYlJA2ajel
XDpcwDL9RSAV9BM9kWVy31Ly0ozybqUcjdRNrrbaU/jutbUO+CKqwwFBKAJm
ZX6ciMu/V6CO/4VIMOqQta4HfjT0pejewOWnbXbx8SvDTeFSJparO7cfkUUm
l9dP+G/LvYJYpPQXogTbDswlJh8FIcyOu5C+DRtR7+sODGCvwYfIc7KNbsCp
4EDM5xn0SJUdh71rhX28rfwb2s7zKRhhq95A3oo4UP88CZSvO8uQaJJOSwRG
N3gunLlHj4nsU9pz2PGHwk99OU3/QB63QqK7OFEM/3j90hQqwHhAjCdRRBj0
YGH4R4GUZtAlbERWutrEERBigtAPdyoMnYa2WNl36psFldhJ7dPKnSlzS/11
N19hjvqIEiwQvfZeEq1ZMBs/Ygczcx2cS5QZpcU9P0Vt1rVic5XoEiJzWnw0
DLBlPHTdepBwWkkQjKdZU6k+eTCyiYewRsatjxj2zybQgnsgR4P99SAgswdq
b/jefMroOx9yfD96YKdMlI+Qh9kPhke5AkydeIf7Qy3pd+9alqxMo2phG/sJ
TrqZnGwOAuDzhpF/mPMK1EwLQDZ7qpS+3fEWMg7Q1bpZOtSFkHve1XfyEmbe
d5MlaGue7j1EIIrn9A04nxCkfea2YOuxwBr0Zt3GvSxSg5gVGJqOT5PIGuLY
3iASHocsyijWlPb9B+NDETlcZU9bRa7JKR9mAB6afPDOA8RXViTPUpfILfNi
OLkWAD5d2FAHXQtDKyZBWPdP/CrM4w3qmh2XH6ArgB2PTeBiSoMP2TkHlF4Y
OVQJSdl4LW9lGvPXVNPV5fMbl43twZuS5DEoHjdy3Y4O6q+7otGaLTsiL+PT
L7v9w58UJ48dYdx5GQbisrmmu6htJPKgb0JPqgGpWPMaeL/9r4Kbt3SBefQI
LgauuIjxhcCdZzJYBwQ0XIEbUhCrm9SMtRprrwH1v9l7dM8fL06bQSWw3n4z
DroKcThsnW5DN9cWA/mdwBB5sEGwPA6qBl3fqTbnv7sLwuOLMrxps/nWAnnd
1YevEVMCUNlr2NeWxSFTCb9wftAPNHnVkrYzxv9vflQiAhLiLJygeliWt5Ui
FrqWkmIFh52zpFT0NMRGJRYWy1bbnhbx8D2hxNWGK42k88l9cgDtlCjQJfWQ
8N3ZoOHKYJscaTcXiNXRh+eB27oa2NMKQftZSwung6NAznj256bia5/ikdXY
HkScS++hQqvBUnlrHj4sAuULxi5N21flnLzkgUOrIbdta5NkzwoCXKA5ZF/4
q55SyCIL03sVIUAsMdgeL3XreDh4M7Naudls0CCCDemIgarQtiSCv5UspifS
tsaBf+Zghm4EURdfX3EW2c3C7B5CDUKMf8n1qUxRhI0OJT/DBE0UpzvDEqMM
9sZhRkel44J/UffF1WY0wF4yPZWgZkv2/awx48lHIndZMtSNmvw3lD7kOjlt
nHXjxFR+ScPmVJQ0VrZH42BUAQXPaiRRjsMhT0krvsC0hcQvqB+66twUgg7g
vMP0nlUejMcdjuVjYcF6KTzj+UCeIUfIoXuZ/bhdd76QwAl3fD1HT4PmQ9TE
YB9+aE7rtjc/c1hBGjRZTeBRbw/ApbDJFEkbnrgcdrJ5WllXqkcE0JziWIGb
Nq3EWW729mH0pTIkQHG03PQ7Xw0+vw3443RsMSHdMvnX5H0S5WUIZ7Zb/H3B
6TIsdXdRJXLgxwTKc3rpDtCMSpA7yaOOV7c2GllGqD1xGQcq9VIz2oe2+icq
Vv/aacA9m+LyUBlfpc+5gima9mJtpfXbXOtYrUVPtudy+2kW5vDilc7Er0uQ
CyMq2dSQBFSmWRVeecRdesB98IMeGZnSKTfMg53oJ237XJfKvo+wGQMJ3Pam
cFwRkQk3mTGNiEGQxBu5C3ZNTYNuZJKdwElq5MY8YleDgaII6J9kLLZAs40y
IxuR8Q5lbWBDMPk4AXMG9BB0C1nXywTlocV/S4aybBPUwwaub2xqt9saKAOZ
bKzCVHlFgiimTIvXsDcX6867HCUotUJw3iDoXJxHx9TmvkTzNbc0pMwBrY4U
oqGXSdQFUVml5XgffkkaLKHUimtbxjnEfIhXzsHUCo5hgHtxr1+9aNx9fHd/
P3h8tpViNPs1FVpID1zvB5ABIZKhElFpavYOYuCXcJQ5hs8892NX0PcEg/TH
Lvgl+TCw57e7qXtcjzo3TscCJMzKdv9ARncxSg5YmRn0iOoWlYLLp4dx6Okk
1HDa2dF1ahGJJYpy3b3NcOg1afomqh5F6G2jJ11R/4jjEWK13gP5NdEGqqZZ
g4IUuAjX5Qmgpiu3Uba5GL+RlQBbT2+mQ2mzVaiiVHwQrRAKSbsVTJxHJB5J
Hgf8xauUEKWI0HF5wxpO0k2Bdu7rJevchP0DQ9ueZhOmN6S8SR0DigkEEIl0
b57xrLC9OOwA+AQu/cbmvl3UvCu7NShufrsTQbFaoMJKBvHfDtdy+4jPmUly
DYHPqkdKg6K+BsKvGTs1FMYCwPm5AZFswGLHzLY9eltYATJYUdloVIMyHo62
rI53TuoskTaDlRcEHv0WmwQTorELVQGpcwZvOqXJQMX3q1G4S/UFKmMdc8ae
98CIcyOS23cRHnkzBVn3LN8LZmwf0QO0aO+rjjtQc1IJpBAyVaQgwMCzeoOA
EkSpwWXb4dP+D5K8hlGbQkUuwWOPfcw1A9ukxCXU4mSX0uTvvN6vgIOQoxoX
snBTX+dZjI4SDA8SmdAChe4ZqJkZIsidSNZbJJWtQXdl6C649KDzscHuGE05
wx9PyYDYWiH3D5q++eLYNXjwGsjUcrepfuTkJjlNPLG8Sas7Vv1Ly1e1B4tn
6gCx6CAo2CB8TCtUEn0uZruTivH778oV5kylvbTL6VEcxIZaxOTEXf71z9T+
jbKxnQA0YeAnrVNjLiytlZMgEPf7S35k7xGjZEjE5EuEd0x4s8ilRJ28Ho7a
VjaVMauqFtbGAnmmkJ84jxc4eGJVm0x8DZ84CfJEsirIBJCyrAOMVhSBgXMg
SuHoWJdGDgtfa1BCgimzOIRuQOR9xx4D6/zI7CCOWuK4JBti4dj25Bp0Xk7K
gRpjeVbp8r5J8p6rPoodBtY29A5z5UgBn0gxUf4p+z7qynGEge9RAb7slki+
mlWSWJDkTdaRgu8EaAGpJo6Xeajn4LE5GZDddMU86wq/AQpxfY7Yw4oaSQIM
r/gr4XTvdQj3RJF4tICYVPUxIdBjS2Aqz7zhM1vV4HBv72/Mw7FUNq/gBt7m
T0GwJK71PIbFgBAg7YT21vSz2ZBeU4F9mEgEPGvxQoqZhwznImB2ey9ce5v6
jJ5JYmNaMwzRhgK7Sq4HarI4WWceZx4EphfNfsqsuWxl/HtgtRv7e4AlUlVK
MgTQx4eYULABxaiD/vo++RWXKae+iaMUbwci+kI5q0Ox/17q0EBw6uYD+sLe
tmGxA17ANkU1XQHOdhPNoypQIxmKDjuFFtD7LW5e03wovKEJqCcX48MbHX+N
CDqYp+Uux49Poke6gOiPXzgENhJBM2R/oa3r3agQN5OlZUtY6o1zWFNho4+N
aOpya5lHHlap5JrSkXaty4eeeFAReiUvZFEIWcnyoW4ATFHlXJj8mt/Pj1qY
8z+p17tFsY+tLCAWgxRoF+8O6KEnrSwiaMJChkMxrhu+g+cOvlYRDyfRyayv
SZ986trYcEpEFcPmFiHqPeEbbdl7ube/TvH/0ed+oFeu1eY11ELRxHvhLIvT
qZGDbqqICrdgj83dpnxsleWpnxgi5R5HTYMvHfAIe3VPioJTchElWE/v0ZvF
dmgVIdLDXSv1eo+lc8RCsU7svdyiJZLL6WKfqMpqfR95Mir2RpeymsFQn/zV
RHUT2++rlKaYiWr87IMJV8agHW8jSURh3jEXtkV9pk+YqZs80DSbiTStKfBO
sv4s/G3Ip0j7X0qxFAEakXeNiCHWYpYN8UVSF5aO1h6eInePnvzesK4+ADdk
93Os/xrh5vh1OxFb8L3u5PXJjJ4xuQDZW795vMIMK7/i/VrgpZHSHHbCIdjE
eYl25uPnhOcc8a6eMfrEXfxdk6bEyTaGrztqADI+UPO2O/e5eaNqHeO3BT7a
NE0nlJevvn4J/Yt2bb9XCjVWIvTTzxkVsj+zGCRiW0X95CBL+n1plRp/DSkH
B96PEjmYNJklTEhXDMhL1ITvr8MJxUG3fidX0yg2BmkvF3QjeDpaC3/EQv6O
dM7wDzqeEcEID2TH6CRz1BiuhhvyIkuWjjBfdIEgKwdHimcjJ+/GtbucMSty
TNPCHfBxS29d3afpq0XhqoH8Gr0KMJZTOlAMuKsuWlV5+bgaAuI6qRnYVKZl
qlHNlGTWhP0dOWwYlfD+Id6oxHLFDukwVG1Nw1bk6pMNdhHU8ysgsGPIolSQ
W9Uk/i8r142459fG2ZlefReMc7RwrNkvfB7Yd6EKib4mE8BIn6FfSerEgCB3
wcp0x4JZvRfQ0+e4S/zghNUxZmKUeYhbGFgwMqVyN6Sx74HtawV8jCk3zGKx
16soR7tK9+YIBsNgE6CuMgz8/2fTtsIzsaUZrx34X+UJLdVVFeS65CiHcvyu
Rd3yVOi3lkwx1h9y5x5RvXSHAB/9LcxcrG8vDwv8s4NfzsN2qu7fA69PGqd+
eknFFUwtunBC+9ywpBa7f9Rbvlvk2LOD76SuyHgGq2RlucMzBPfuu/FnhJ0l
V4pHpLOS573vT4K9fplgZudoTfuV2+ivCCUggVSfHxWV1j1REC0H5fZGrWV+
raEytNJk36/5OFx8k5L0n/77CTcdMtXUln3M3JmUIUTK7SBSwjooH5iscndP
PXk0+DR1aXUcOV1/HkfCxVFaQ98G3wQeKQhGwJLIf+/n6pdqfkCd9PLPRAcS
kjVBIGxaLMs404dkbLbBYimvg6E55bW/l6P4NLBhEryK99fJjgmOSOWEhqFv
0PkQaXeP5nc22ehUlPcEexogFMR3qFTsApueJB4PiBuuN1bcFx/z+ge1lsiv
5M3Oo31YgBQvC7+NCariGXkRJMXwU56a6Rm/M+01mq9T2mUiRhQav8eb+kV5
Kd+dHx/93xfYkCs/HL1QpysloZi+Pr7eT0GmiwMRNRxbJV4Kyo7hoWaJRDsy
JI1NcRbrstB4gQvNSh5/1R6bn6Eq3cfS0Mru5EswLlIgsA3jpbrLwIN6PQnI
7UispCK8Yt5WTuQdyyom0kmA0PGlieSk1VdGWmLYaGdUgOoDD9UPZh69GdG4
SgsN0lopPYVoKtENeaPKrZbf9TPOGvtsfChKV6gnHb51d0yir2dizrPHYGag
HX5AL44SQFcNNdHMrISM3Sd4GpkcHptC6qBG7XkOb7L+BoPSPehSy/rCcVcY
jVjizyINWOOkSMyqScxgYXeekGq4ecLlCGE8lg+MO3L76MS4GoRHDd/esFHH
VYAG0JkyVAZ9MtQV78u09eg8kzwd+WAL9+208zf12f/wCOUicHoKYzfE15+A
KCgXi9MQcfBUODm7vXSCBW2gQrSpZZ43xHXG8mvpc0bBV/8INUJpXAzkd69u
Yrtpm6tu6eXZ5XBeIM46SJW4lrmtgWZszovHwewmm44cdbg6LE+OmPWOsJnB
THxQI+OEc1yRaKHmSslFbz7zPzzDRDTW7BkCUHzPTxdtNO7r/19LSq9bpBX7
kV6/Ezzun7U2IC0pWMoqXKvAfMNpTegXIfXPSu7kKsGyOwcw4/IesFbleZjZ
PBYa4njY3uCGH43g0Oq5VidtM7dUU+llLBIGa2eN3A5qA+Nhj3nfPy+6XB1Y
hvAThKFIQzFy48OzmiEtCsnr8iX2FBjQn6FQY7mnfyv2MWg34fYJBWPZXpgK
oJzA2CcoJZ90JXjdP4q/hufpsr2ac3xacsjXjTf7zEVWhA+d/rfweI7Wb+Vm
AKnWk9jOZBNYTRGbs5fiFvitF1ShkQy2vA/Md3GEY3Iz3wqrkodkZxy+Tljr
P5V8L3TEIJugtWXNpobJCrdEgBbEBo/LXDJdH5BSUBcZM2RiWG2bYlcf1kGk
eBrXoGKylf/91SCfvtjfTt0q4505UMJx3hW7lnu/01AYuUaJBGSH0Igk/D7W
h1mEb+lrZbHEFz/Ax4mG+mJ4ooXXRgSJw2z76vonPsmaF2Smi5orGecVvhrQ
ttetZG6+66Zlqb207vDdqeF3/rxZUkr7C+XUs3lq5+iuu9IvbuJ2pC1H3XHD
tSRJWQF8RQvOGX4V88kvupwYet+uD6CrHYEm/Oy7Iaf5rrSO34wka3q5yHlr
Ut3yqTeSOF5uTVdDfIkdWWce1o7CsCKdM4s9whWhTqs8lESqA/jT9fb7sfTT
JzNKN68mdriqxPpoINWztB1oLpgHDxwdktfp1DAByavu6XYmmHg//pBVi0tB
JM/9CYHgdA+HkDk+WtWJJC5JIVmfQD0uxW5OsS8CVsG2GfFUtVWkBox7w9sh
tfKGBup0eoJiZ3tAoZBFUczAZYXCLo9GKbQiPz8pmufh9E7L7vBg4HpivrNj
ZMMKAn32LB4/X0f6LrsGvJKuG8a+Z12y8Z0odiIBLclBhDi82Jji7whthsNm
sugR3iIX7wiTBAEhL4m5hvHIob13sZaMuMcmIBTN1h9pSYn8GEQVGU5M2oFh
zWnLfLBg80E4ZS1Gwf/4oMXCmK+ks9IUWabFYtg8xzDvRUldw8+fabVI00V7
ueReEPIkndGlLz8ZKPNbnllsGmiL73MHAXjXerfEfBYb8ILP0Z6QU1xs5xLN
NHZeIg0kVqgMuDqpvTrNwwhvQQvplTlyyPwX1xeDvf6H6vXfZocGaL9azrPn
EytjrGZgDcAYGXUBx34j1g70wKWKZsP3jyYeCSBrchOmjfCyINQqsxigG3SF
E9xMOuW71boHDauRw2IwGmU+AbIU6f/POb6vRBGidrNMo13pqcffnHGIpsq3
yhi7ZCfwPTiZ+P4rDusb+7fcJwC6i7N1ajSec0P5EwpN7e4eDhgpR2H/9cG7
klpKrUs0awkjkVtSBqeddksIF7qUoW0VCtlZ+ZIaD4ZS/U7Va/Jqa2+lJxNN
04rCxBC+3gTBZy3QhkJEV5ddUMMQi8z6ACE+QYCYoHIEViqRiTi8az+Egijf
puVI3P8/+mOII8v7j9ct1sb86NUDLYuHX0+CnTMRqrgz/pDCFYFo39R0RhqW
imtI1EP+qv3rUbCHGaSwpMsXVqCz51S2ewbpVHdg17IFOpBUx7p++kEmIHdf
B8SHI3UjvTeywlprqPqFpY2grw9ThrwE+mNpI25BPOmF7YqKbO+/GxpZNCvo
nts2W33561GvtBlhTlUm79+KIL6optRoW0Q+HlanwgX7Y3d1svdn3PpVMcUU
NSeBsPVhc2+WfmGxlyv9syrueQQSbGrWHNTM4+E8gyvLsZ/Eeyzei2Y4TuA7
DCx4+u5PFtnLw4323c4tliGX36oMh7BJRg+kMnpWn/gpAUqL1ytvJeoWdHKb
ZW+oc0gNtVrFjTMESHOVmD2lwhGQtITbtFIVqFGsylom5P+bHOJJzUDZrOTs
L+L0mxQj1hG/iJg+xFvfxfD0hOHznGW6MEefk9QJ5HaECP3q8fBYYcDdZt+S
+BSib4Sl403QDoLOaB1Al6ZJSSP8iiezxe2VYrg28k4tzUfi+l4wYB6VIk3j
wTUKNgu5QqjDnD+ucxk3GZuOkpF6Aa80Cehz/yCBKywdooWcyQgt4C0ldv4y
AeHtD0TslixHYNG+p8Ykq/VKqf8cAeNWERyXwElwURS+c57vrPWZMcxxFaBD
8vMpAWoWH8kbSr2MOHqv9S+vmR1SSbwoWB1zi1anPjx/IoWsnmvTXBu5o9lu
nhwjrIIfcCgcRxcTS12hLz9rUviJjrGILZ1TVMvEBZ+BD3pXbIMRK276j7Px
sJM2mqLdHYmz993jvmYCVUCGS9uf/OD0gwZABeaFPFAXqVleIM4CoZ/0fu9q
x7LHGXTqXCPpur8vv0FG3+NiHK5KJUCe87B9Tn7iNaVKmBLsgJSyU7p0XQDk
5J0G2tpNY9/saoRMfY/2Cqq0BgsI0DdCqSQ3uUY8hRwKfTj1dRJk/0WevLto
qcEeFtk2nEer3WpgWe7PMSG+fXEQg/ktys4F1TYtlhK5oO5dsCkUrbmxLKDL
x1KFGMjn8K/PnK/227cgDzG408SVpgQp6zC1Mx6844vyCqpBXxJIg8OWv5aA
qreUCP5INJhZ8bgA0S3+wtz6ahSluNp/vjCsRPJ6zTBFU0QKLyceK7bdA5Fq
5zbcYH/jtJ8Y/bJmDwvCqz2MBdL6dFHpKcroenUH5+54Qt5tS5B5GXvrZg5J
ma42qaqS28EeQfw5F3OxBrDRyUpVaWMfKMu+8DGyKg0iIk/zCSx4cDtPkG3t
oSE4oqXG8/v9U15q+2PepO7Ka1kIkVXxSzXTycnKB06ScGFy67qbk96fUqum
9hBur0D9ZW+d2rZknV2qSgqGtcROlxzCuv0zsoJfohpFdTOdngSSXWtuWQfz
DJ/aSeL4NEtXLPH7l/mEAWnFBzsZsEyA3BaELrrI+qHPb7+Ow54chGhtk225
XGt+SPKs70wm+AmTnDvd5TD4cWvVBBIesvP4KzkRF5+AAvwSO4hUpgbs0zOg
ThzLlgNKZW+Vcpmipz/ydrlMeuRL7F18gCcx+257fArlXFSw6h31tG8zjJaS
E0u2DBBxVHs64Ddpj0I/v26cPYWdTJ5DcWO0vLfaAc9g6MEGq/cNPRqMkFAx
/YJ2nPDwIkA+QJWzzLOnYlPVm5eOlphQNprik+8wsAt43JEsCGK34velxjVY
t39KxFugxTG+DDgTYsvWymM4RnoXQGyGyDrlrfqElGu/B5ZgN9PEhM/Y8sjW
A2GZMKMsQt1QBLt8CopWCkUu931yMCAqDs+X4MvCJwtGFW/edcJH93942WY/
F10NbGbx726daslZR4IXzZlWO6AFS+i0T+mG60ptTnYJyVsTraL7xbHR+w/e
OdunjR4IKNFhKt6ouvsB7LU1Dros2Q205+Osdcb7+NqGzJ6ujlI7+XN859Rt
lvgxmDx0pjqomETdJQt8AEaZ/1ysUzn95UEZDrw9bFdB6Sn3wdBLUJa/bRgK
/hSNecvI2ykri2PgaTEarIfo7fRRA0+FEKivHLX0S9S1sAQ9yTpeLxsaD/D8
MXj7brhbXL4gi/glAuUK6+QTfCWBGlNBosaKWKDAxv7gc5YuNO/s8q/eDzML
G9err5i1KdowWxc8HXZ1/S53vBjDpK2Y2vmryOq3+NVTgQH6R17LjiOzSMbk
KViH3oDaVg1uL4CdW+vg195T+QaVpC6W0F764WkYA8MO6kzaVyUH53rSbGvE
JhM8EnIrz02gLQbneQgIdolHnWA26Zq+shojCuazFCaitEbLLui/mC8NYhF9
QrVpGun0XJ9n2GzFfdsUg+QBfzlQ2RVN75Y8EXxzOt7hGOxBGBRPGdYMsaqS
mmmw1WWEtNQonF6OGc3vDD5k7p+uCtF622sbWNzfX0cw37Uqz07oeiKhV9ur
l7hMZVPme7Wb40PIOhbTa7qeJwa9S+B6BfxzVD/u8wfkat+49kj2xVgWiyk5
MyugB0WIPI6zLmhS8nAkbh6Xuopkax/0jBa1CLaA2YOjB0PLi7E1B3t66GeS
C2lmRJM3xA1MEpElv1Fu/aVbNv36b19JntjjwjWgDZaSE7NGII5AZihfFFxK
j/IyTkUI4e6SsUTeBRZdRbYhTdCmiFzqUyQzorBZ4QCZRj0KoJcMT4LrB80h
UcRjmSeinp21etDQFMzNvzd8S1AyOq8IVj7Bx69KVz2uK0PLxsjETXJCnZ1W
zP/Z5T+e21xxftvVRBVDhTO9HME3lgL+wFxW3yAxm4ID9SPe1chO2kJ9qWD3
d+GqIvC2NU0DnpyQE7RLk2uAxEl4tRp7zZgB73UYsqBbSAUHOrwUSw3wAjeM
mIH9igbySwyhHssH5KYQ0czdGoVHIMMRPCDRAHzrtmRtHKO5c/XVjfFZaC0m
E+PXw0mlklF09JR05P4ak4Vq6Zr7C1HZx9SmExcc9vr2WQM8fy81+eGh0oFA
JYOwc1giJXz/ZOwMsrRmhE5Nm80FZKAOHLNaOe5JwEwtdOxU5eBtVlZ3BpER
ggwst2XdLz5ou44si8u3eafiHEKOveHu5VTV9PF5KiHEtXpIKDGhLUzi/MXD
IHAkaQri8vf98L9/shbvtlzPMwK5bVbOusGgxvLXMokc+T250EoLYCf00qNA
XUVGnIoyMh9r+f6rbqF/Dt4oCrQ5HgvZhK0X1pTZ2R6jcFr0iI15rarYR+RF
7rA6OmSGKLUr9HRLNNzppG/di54d91EmcxAQAbX3xGcDU54av43Udbfum+LK
qpEbjBWv/7JoPb44ExuXZkTLwp9PsxBy++omD+dSxxFAvSaWa3T07hbG2Ut6
UdBgiUPcrnhXiYPCqiuI5I4/qEoUGnoa1F6xlG1aI1yOadLdiC+7KtVncfL+
G5thZxau0pq1h4NZD4/cXsJyWEvWvqHNJPLpruGtOCOIatd+1PbUk9TwZHla
Pg1Op+/TcfZYMugmpnTZ24zIy9YWv5ilqNo8gsMt+6I0SxIu4lU3oU3AqSSJ
XWw+vF9lLvD9Bd4i+eAfR84CrtIKW9JNnNvv4/9gigTO0N6BBNOGlOKwoBqK
xem68DEVm5R4VREY8R1wAj0Pu9kt+mdRct3iTBv8dziMtITOxECT+Ddk1mSd
IR5NuCNBJrSmeILDs+4DtrXXMDtLFtB5LoxokLeiFjqknR09PLVfFGU8TIbF
dICddOC+cdexJuQkpkXzrwMGy+VuXAG70WZdrZDjzCBFeFJ32xBIvqciSJ2v
xJQ4hciKI84OqBELfpAwrIuN7Igql+lpbiTQTQmMMYUJknDvZX2iYzbDPAO6
LLb5YbUtlXw9eTwD7giTxHZ4lCWT5TErqAL8tbmFkZxloqzG5olOURZtYTxC
TJyFhAPjPRcFVa2s40eUhJL/dr+hgOVj/VaXixHvZNG5dOPzFtcYH/T/fwSK
gtR/SDdyxzOZyVNIj3eoufKpnmUiIotLlmBFPHnhhtHB1PVvi9cUMLcifHps
wfBGBI2ZhoP/cYVEclWxQcusqu2pAJP9DLJAy8xxgN13jy7VONh3t/B+/Tot
BfAzqqbQNgOe3wbM2TyUjAwyBf0Wik0C1Ag4AuUYezp4CR6hLxw2PoWWwEVq
NLveScKwqzmoldjA5hM31f4pV60YF4iNHggxNj9cv542l3FTNFNxjwaTMOmB
zexzKDqo65InS8DjEnR/7srLWNUQjsklJ2fK4a+NuS12UrVRBgxn8CxUOe3D
XvcZAz/5TBPuSJxD4J/IY78HEM/bXt4q8ONpeNCJ3un+5cCPB8ZY+bIXJm0W
WH9UgGeq11zL5ePtxQiMkNRTrkIMGakcynHvweG8FeDQKr8x/tocA7mA+TqJ
0VwJ/jZPdoFjLERK7BkgBbKq5VmldiJXCDmuU4I+kCXdYuFsn9tJzBomTWND
LIpp4YTBTk0UVesMQiNpddMfFgTCzu4GXmgbKqxbqBzsRzMnsSIrV7TvD2qo
wshRseYBnRBkbrTFK7JHmSZMY0nqbev8DeiIrDTq2AQ4OuTARoJ3O5G1yCJ2
AzWEgjEljfChTDK4H2ksfK8Ru1mSOGlM9unSBAgRPXHGu3EDTpdvY+6bTKJa
kCoFKXYo1EEuaJGFfRRr2dSprw/v5S5BFn++k56n2sZXy/ujxYYsvaXCG/1i
Xi4KIrHnrb763B6yvaaCv+yN+gSh6h8jgyTnDupTs/1IuxPFUeJhJCpKuwKW
2DdkOzjIY0RluOjdNbgxvefjdhy0Pf4Y0g8N/5zICN47iejPziodv9T8EPoe
BudSs40neP9kXJTxIn9xSv7jSJu/mYRPTiPhZPEtfPY0Ot3fDxK1tmZ3NCwG
Qc7lR/AR22ThysflWkpcVSqsX/6rtc+WA/AiqyzOL8opYkdros9Aq4gAAxw8
7Ev9kHum4wj7jpe/hf1+8w60UuacfAtpoZQIJ7L96zVArC6qSDlTSbu4v3ye
VhbPwZ6n56TwJ0ks3C2GU+y5ZuUwSENTzxM8DVNj2mOo/TKeGz8uCn41PW1g
5k64rmzn0xCTMRy2LWGjYnGJkiO3gx4N4R1pNjp2bUFTFbGZrqxMv4HaapTA
DYUYkDieC2XIrNZlWhYrXtsv+H6nggRe+vi4QCp96sSJAXHXPy/2Yb0CbuI1
8Ivv/xwUSK41/lTBMIAei67JJJmRDi/nzONOk0fEY/bbhCEc9F1Kcs1I0Jr0
dzTjiUKcv3olGsx43lpOwR7TS1MyOAmEBY3qOqdyGtVKSHcU2/QZZ4Q+mDWo
+ziottR5KaXl1yWCRGWUDz2HVMv66lBBIfdb/9mQ19lWUV83tWb2luCt2I5B
EPDdZaTMnxoPMSOHw28gYzB+DLttENeMwW2iIPsIOz9N4zgVwj6N+FvFhCRO
dnRniR0FXaHio+boCj2p5BpXlWyLB/Jr4b51VSvrB6iyKnyVveqUrl2ipaLC
hUQp0pbzvMePl1JgH2Ka7bKtZYF8RA1oKnzzBLt/x5ZGdk+xBjTI5N2nn+1X
OsRhyEsGDluemFwBjW+f8KVGau8HVr6tfgMvZlNLQtv/rBLOGeqypEidwzjI
s0+SpprOUNMtWFR4Oczv9lAIXyuLDT58rmjhnb3aJmC/YqQiptEvyxGkKZ9m
2kdAgt/Pqus1GEEhv/Ljjzcf4/qkTvlZK8+qi9kdZmu+BLbGAp+wFABcyCDg
L/LCRKZ9PcjklwIuLFgPGhirk0VHF0YWuo5iUVnag3+kNBWIqoSJ6iH9tNED
UNl6KKl3h+ck23FucgTr8gTLlge7ZPFVsFeo9bgZNDNAW8ktF1WB31XL4ZNe
AX2bwBHTqqRnoHqgkQeLp2eUsyDRWtQmH9vgVohW6jqFr/E4zZX5XY6Iw+yF
5ukXyu3WN46bLraoYmq8gVrwu/yPABixtJVNISA8ZSEVYdOlPFm3P3wvjV6Y
XFYROaEPA8w8zSMyZVCUqd6qRf0/mwoBVkxM+6Hu4ctnjNPtb6qK83E0fvar
PzQK/YEHM1oUAT6mxrlgUF/GUuDjztx3CRTdw4Oc+mlozxW3xIKPzfrtynlZ
hFozz8m3BCIC1uNnbFI2muad29o126EX7f0HQzttNaKXfZ+JVPugOzwdHO2Z
LhQR1+hFsuYWTmzm96HVYj1hq0NfutMo9ZFckUAObbv7DCoK6c2PnbHaS/6x
aL2cYWRIX3EhEKhiOuyOe3G1QnAF6ZXJU2JLRDz+TgFd4YMs7TcEutk3B7uW
VBbi9ipwzMsOc19PEmgSZJ1pv7VKyYvMNXpbAMayI8RFoUe0UQDH314ORFoW
ROoHB98cMLgPGIzcFwZ6HsXwy/fH9xE3T6KZpl/1WW56iIYLyZ0OGmGSkPnn
Pv3S2V/qOf5v2f+vrK+SzyXC8cFDH0k4toalGViYz7gdEavIRfhNDVlaTNiM
H0IRrxlmvePDpx8PDrT31WKkeN9F/7kmwy3BnQDqhiwuhGJzlWSPGJQZjhoV
AeqNAUuNySrSVwfnHF55K8iMvxd8UeMzsdF7Zq0RXHYePQXpjDEkB13rSOCu
G0uWFy+i1jOlV7VvyIrYbOY/CTI1PdExL2nKnnljUIh1vCZqUjvmP6rbXzDu
sKl6jceyZV4CpsiYLUf+00r++8n5FiyWtpI+ta06fSWL7tBd+vrUgsuGS8zS
YqhjirilKOadI+B/WUEUTHbFDV/dclzp11RmmHBZgLFEhd+/hVwudnKhumol
7O1MS6Y9JXK6ZYlhWQv1TqmF6d+vMZqHcZgJsRNyoDXOIfrNK0/o4PB2dHB5
8O5PqsLp8cOsSuOFKjxG/JLr6rEq7B/Egdq20x7rj1S+1GduBJxMXMv1pD8B
tZzr2AEk8CJrP6zAq0L8ofZ1akdg7Ktj+9OcZqI6oRo7mixMpgAhK29S5EwW
j872VHofMV9zT5qUcmKRXKpQUM7A6xHIPV0j7NKwU7YueHEf1a8UENO7Q8+s
sWetXc9GYD0yKUyPp+pZCvyZHZEgnT1qBNnHoK74ZkI5vz+2ny2fI/EUtyMG
SAWmA0DYLWMpxsLsYeAJTZUEs6kwEDfbq11UaDWVp1lX9oxRazSMBQKnYPMw
UfQNxmxtph5ZPnVMRKMKkTJLl+evOzZmbT+JXPIsFATKG6e3NqkfC41s3MW7
yggLSnGbmyW3tRoALCiOp9JIZUia8vINieALMcu+QT/xU8R00QX4WGkdKkd6
4NYzUqGP9rmDS9AvCWbzZ+ZcikEQW9SK4DIGOdSCOdVzAJkdp02kHR7Wcrka
Dgw+tNKlspWhPzN8GyxcAD7ULOrB1zp2+qczIPcrVX4ajf1oKlxdvh8Eueve
MEw3q4vD0GQWA42j8T0HgyWK5ZOiOASP34Acx/afIrgKT54rPY0Lzct5L81m
lD1Yn7X53mn6dC6MQdK+q+mIDZpbV3LEPBvYYr+izYAT2B2r09EPIE4lYo7V
ODHQBwUKjkRuecUjlM1Y6SCNiALi2RWGxZhg+/fVwYNhAMUcLc+nlFS9DDDU
xvOr/0TFzSs6GZ4bQrco/1QC6qBC6qMurB0LEIGd1Qu//e/qjyaHC91ijd9K
fuTdZ4I22O54m7O1ZFEVHnPclp5JyNSRzaleOfpDtnR31klojSIhA6W7Vgln
TAYQuAXvxDt0HTpNE4/fmpfSeKDJijHV1+lDI60vFKASdQuS96yi6WIOS+EG
so/7kqlQtrjF+nVr2v1iLSyTZi9wW5HJPRf/7P6oKJ8dO6ibwbE5HPGJdqir
CIp701BjdcMJJbeRRUTE799hlQ5bw76IXaC8UiFoha/T/ZFUDvVSMRqIWyzg
4mkRCBLDdBy75rcor6nujmZRaf0+Lfh6mctsekKJu6FDO1THQkzPV1dQqDdm
t8S54ZEDMIltZOpzWw8g/TrQeqd/EgXAOn4F3x8jahXwESz0I17UDOEANOq4
g+0Rr+UMH4IlvJNL0P7ShtPOX9m5cQJzRyi0afwGcQKDCP2HqYB7jWUjgjaC
L9b+voqOr6LHffYXRbT8SfNxX0ZHkVrWc7YI1DdVDrqUjuKVKcrmlsBp1akt
71ZJF869ktTD+NMLsJrCu3YO6Cza8+fjUmu/iVYEkq6QdAEaDzckzGACGgqN
Wc1WMkjfPOJoRLz2PKt2m1KgfKdW1eTmFcsjJXzdWBpqcttSovumxmqaiieM
jDEWS5Au7l7rEhk8GIlT5kefIMebj6lVMZybAmwV6r8Zyq7GT3rmd8SBDDvh
58AwzTmgOsXdJZYRADG+hryeLAvMvnEPf+anhozBLpYozvXfYd2CiGqDiGJh
07d/7bthH7dTIJnBUzsjzFIUECVJJCAgvnDecfRH0lmSM0aq6wLNGN8k7kKG
8sucPHEJlKbUiHhLUix9kRU1uk1qbKJsNkFvW+Xjfawrfzr0oyoWQmRNwfka
O9oTlKx7hr5VxedICxPxx8Y8z/ssXQzVLjSI+DQPdwzSgmtKZ3ZiRlwL/n1X
Re6RukDC/izjFUxrhQmQ+MhzXOooHEQQOPFtLfciKW05BIHQ09EKAde1VYzP
PLwE0yU15zJ7aPQEruxSJwnd+Me6b5Aks/Fz/BoEveuTJkn6Yr30CcMczWMc
8Bd+mxGkCGSzCHCUZggj2M87ce2ZJ+uPMkWQqorB8FVUijg8fJyQctRLHuOm
e9QfIawnryahswW9VvCwNJ0MAEJ5MqDsX6cvDOj5nCUbiFS1ErG5qynvORRh
mHvMR9hQWvG26MXdUpDRNEBoTpKguATzCidjdKWSe01KhGBgShkD/oP/y070
mK9/eYsNLBNXMqmtMQ8OOCDRvTKJ+DKCqV0zx6uubC+V+NZzx5eCs3je338M
KXb3TR0KHEUL7ZgAv3TTZasd1Q8vGehuTkl7eIfukwoBFQkFBPV6/XzR8YBT
8FTxHbdkYxwkO25nyJk71v+T/t0xdpIMWLgItJWir4vak9B+5NZZpYFFIZJt
jDGrEUgGrLTCbpBE6kSkiZ7zfS3Mo2d6QF/CkaIrJnnZy5JKizDo/qKnbox9
6nNGz1b+n13WF1RjnLBi8Jwy537mD+xVRA/GEXYafTiDp3oVEFCAntRYR2lB
0WgEMPmSbsvo2wSbnwd1HMAxvY7vQa9GZcpgBDa+nZQvIpREGHuaxxj/1ZOb
kRuuZEGcNbMYPFpOb+6QGXyXAM5aldC8kTD55s87340Wpw8C41Ny1mucQPYC
+oNX17TCKMauncNF5V1ELRPey2DEhwgCF45RdEtdySAKS8badlxeG0br80Jl
dmrNaGMDprwrLjj5pMSg9HmFC1c0LMUxdN1ExfO01Z/ilu3lDC+uGSkTahge
FYgNrY2y+yRZ7CgVSwr+Fd38vhZOCcnyjeohRRdLsEc6DhiW7BPpg5svLvAl
15z/LI8pCEtKJxJInbjg/QQXURBKxxMKEYAADpv2yLcQZ7oNClXZrq06QyO8
cWthW8ZegpI93ID20bvZ2Sk8bnyjvs1DHA1aqKPlIBA6Xg8ur3mCIr4tWin2
08raXYMDIQY1XsG4eh/OhrxuO/OUVRvkqAyE6MmSpeeEhrwdjIVpoYQUsAzB
GSdxVCWXymxvU9Xje+ir0etRhyHz1WYPzCcc4+XV5vOQ14dEVwwgx0CpE0l6
Pr7ZCTQVquojKi+Qo1TNRx4gZv5KR6M8EXTMUUPw2pGMevFGE9vWd4y2YMI5
/Jp2GUFFUQHFhWjXK/ZqjkyQyHG4KjrMB00pXJEZg2zy5gx1DqA0E6fHsRy0
Ms6rG7mQOH7WkkstJb8H9/fFHMzDhylsidNBXoQ5AB+WT1JLUC6iLUN+xujg
9aiViEkqD2iOAqF7pJVUyt5Me7hg7jzatbCMjdVTu1mcO/CnPDZ7wz/hhSV+
8TBTg8yHe+A3FLKTtlPgp7aohq3+M9vxP6hv2V2BpugJn9489JOJVYQx5VH9
ssv+8d30rwc4xMbIaCTwb6abGrMawlWiiHatrZDSvFt5gdjWE+k0UuT30avc
QL4LGA73D8L0YLwUSAZALfJCAh6ergZXpuEA+ED+BI393tQoACZw6dyRHHUZ
/uxGNhWr3gry5L5o5UjaTJ8ZCPiXgLNH5ca19so4bp6LsyabcZUs+pKLIrSt
4JpoE7vZLxpxCcUmfJEzMjWguIg3Ck0wH+9DAKbxajNQQVpGDA5cSQwA6gpi
AzVfbTBh+GVtY07ObOxtqJwEyTsI6Lm6KUHWgOtUaVfZWKeBqyWe05j8qrOW
roaZPQoyNcF9RZIcRmXAgwTHEcsLp4I3Okr9+E03lj1cwcqLawsUXbZPhqDV
bmKggyd525PUy18NuyPSnw9fVQNZxfpqpI2dXxWP/VyJxI/pWxN6whE/pvNp
s9FMG5GUTcIvYsHOOyuPFdxKekOPn8GlbYDnk+mM1R2MhzoNc6h/xLWPTs+J
YupoH9OQowYVLvzEU/s6zkS0zWT0OWXaRkFFboavG4aDMhd1yFFRHw0s7weq
XL5YXcuZEN1TAnxj5Vns/NAMslqa/iWYE4PqiiMigunfGGWd+5SZZhephkJp
kFM+wv0avshuAig0w1BTJOnRJl/lXf0PUVXACmOEYBOEWMPanEij096vxy6q
bcf0OzbQMeppie8cEOmjVoQeb3EFL7NW7jvFdl0ArA9glAO5TaaHFw0wCnVt
WxTMUpRzIqfJL5nwTLLFya0JzQgGwi5LS0PNBb5iBXZ+jNLfdne4jH+W1tFG
zIezJchgymjdWmE8nHOZfgFagPs18ekw+rpIZhwF8Qk88fBP3pyqRaefLMhr
PbqD4gta7h/4SDoNxGuKUb/dr3ZKBd9a5/Yyus+9Iu2G2Brvj7e9WcVH4OBT
DACAErMhoc5oC8/oS8XenB0apljV9BcUcToFDljktWdTeWpLn22X3VFrdjKO
Pu9zPaot74phljvmC2KxVnu5yQVJANKtcmLESvPuwAxLIDB9Pvlx0a8EpLqI
beM5TA/rLbBX2RqkgzMeCevggmJfWimtkyNqMeRO6YI7XusnyCOigl4ANJ0W
embXwaoeTac2S8lyd9ulp6TPi7jlByHTXC5Ri9u795eYnwXwFl3LrIeF2+Hy
NgrKE6uVlfRfv/dsnrTSXhsmaHk4aE0lRLESCYUNiMiEwPcSxSIBQkGUN47t
PNhqK2fUTlkWXpphYKFa54DNMlP+6lRToaAblgBT0XBK4GutBtynr39lThuH
CSzavbZdWoQLf7wKlneJQDFUfqACuMuCbH78v55IW6P1gOILub4AGvZf6bh8
wE3Wgxl0JEEW1wLspgAQVIfC9O4rpdloRAJ7+h8ZeiHqur+CqKdvtsBhuBtk
ntKBvvhWJYkZQPYmxvT+fcNEr9kqz36X5IXljq591MXqfIIu2hXWIqJm3c6q
oNyFB0H8cgTPE8r3QxkDOeCFpFYFun/NnJrD35iGBnXTMYdocYG7fj9wvh+I
0rE9f2yufGEHa6WI1Lb4PHmm4bMvu7EmbjoPqLZaZ1q8Gs0dO7Lw2/Gy+6BE
2XorWMYVjktbvgym0iHa4L+QO45g4pMkUzEXlWqPDdsss3heroposCve1Jd4
b2XIShAJWfPzy878O2DTnkwbaHrRjCrfKVgPqrwHnADTbQgc4ViBkWIOhfFC
kkNnXH5Pdl1AlOzgM/dQDSDKV8ZCPPUDp7noTj3seDS0hhUQ6Crzz4iq6gzf
nwXdHlXZnaCirzVJaADbIGqp8t0CyLUCp7sc0JlxSJwksCw6bOFsudwEo5km
58wywxP+f7/96OPM/WZB0ccGhXtdaqIN6HoOUJQwOtuwRX5MeJhdBRKWlMQw
7REkueJEM4Xa1zw/7p5+gPz5zNrnRPuLa+GrEG5RqKKv+S7PIDao6LnUKQ6Y
sH+kQ4jzV4drNvQxQtraN3/ePssedOgzQzJXaeM+yKl0cj9LTtWfA3qrXHDD
gFU7pHJwhVB5pZsykZsjiCT5eqrxgUlcLolt8x7Q492h4EgUgtAw/OrgIe1/
5xhbUvfaR2DFRyMXHa0qiyMeZcBdrE0g8g6tP3AF08XqPJloj7s7H3Jerk3T
LmGV0EBeR9KKo7m/SJxKPcpSDqCbw2qMEQMLFdFZhZjv66ZFZlvtkNuy+1jD
gRdobNkcC9ISE2d42uPxSvB5F/29YJte9zCu8/aJ0hhkk12YuQe1ELYz4HT5
shjibbcRtk3AJjS3Jc4M/BPXwFKKB59h/cU2RCwAob32+hnQTZ+U0yVSik8v
S4f8L11pUeB900r523xJ696yKNA5+bALR4r1iWzhctiEPkhgGy2/qGywG/VM
Z88ZLOzRs4BSzB59W4lxUC87Qtos6u+oTZ3eu0iE/Ujg+5KCZdOBMBnao46D
uJt693hHHkW9S2IqxR+rOO6Mi0X6Z8r8MVGOI6Dw9S5jepN3VORljTc2O6kG
VMG5wsHUQn0Le0ers/qr8l043N7+DJxsEkVgmreJOIpHSPK3Xpt/Ns2btx6g
OJ5KMuBnI0lPMgOGNg660uvTVB/BHymPt6hRlHCX5OUobMIqymPgK2nPjMCI
pHrCmXku0z38uK0k9jZ/pUGKQtM/GxXutJUQnWIacm8uQ37/8byAXB5mfNMs
Fim6mxSbfZFejAGOcXa2jwRHSRqiKZ+N1UlOnSmjqb/60Mob6Zd4oNm3PK2l
/t046hB8eFDHcBQXmOL7GwO6iSy92oo7j57uDVGifXQ3iEwrRnPPJLHHHGqF
S26iq8CLGh8JpaPciQU26xLOUqI27hsbvo2mmvN3/1u/w6bGcF0Adp0z888a
HoneQLb5eZ7kWckMsCtjgntQyZWG6e/rBvtO1HS73aExnSBbG/+vNrvxc7yH
Q9TyU+es81pdVfHtlPrqzv1yUB+6sMJx0fkAi3XCiZJxAgzmRTZc/jLw1oQw
SyPTDfnYl6W6TF44fzCCuL3FZTvcImPESQdR86eHu/Czs6T4+5yaXQKHxbbk
Lm/JcaJX1l3YJ6nqyeX5jpEnT6qSEMXV7EaIyPkdh2gfi9Jn3FongNAHZSTs
4elExyDuvutl71MFFV9/jOP3XgI/lyN2hxealvPRG41sSGJfxBM5pWA6GSxI
Wqe3GCVSIh0rAmdrLluOLum4GPgfho6Fywgwl82rbNRsCi4FYPW8QPF9zTWY
Uv4s45IptMWP8IBO1aWWBAPCtiYO8clc8GcA9YcBJGdo4UTJk1vkmNIgxapn
8Hagbo6cFfU2E65r4HTjNsNSMJo1yMyumpOgeXEmTBv34xrQ/RkNin5Qe6RY
aI/uAFzYmLM0eoXV6AvBLApM2Tl2DbYjihDIIHxhmEccewhtJk25CXQ7DZRS
VQBddc42xAemRTc3hwj99vG7zwXS56frhffWhkxl3NPd4SrSZjA431Q5DEom
i7cuJUp2MjXyK36zkNxC1O5iZY4zGQe4TaCh+8SxP/ZetYGgj2sTmVemOs+J
e4Bcvtk8VDHLvEFBQQjetIDk4UsHQgD1cUMYgzqRZkxptRgJihtRbFp/kE1L
j/7wFXIOz057e6Y1IDdjojfklqLeieAirK8lhgMIqc4kTn6D/2Nm1S+r4ywV
HyurL+uf0rszl/hayglbJk2C528UMA7GSLFJWq7JqDWwK3YTd2Irh5P5N0Lo
6UgN+S0tWzru2kUr3wTwVIcFQDdykP1GlJDkiIpHjxTJcP311bNJv3Y5Nxnk
DL3RMFIpxs0l0XH6G/LaLa5QiVS3KGzjrEfpGaURd217CAKgYg4agwIhncn6
QSBf2+oNZDLlP4dh6Fv88EbO36D9K7FhuiglG4/2xeAab/sVAr/WVbvAxdJf
CGrBvkf6/04ATbaceixP3FWh8ojgoUAQ8VKe1DVCLjYU6yrOzKPIHQfn3LNq
H4arB1aUdHNCxMgIwS+eIH0LQNp41JxXteaxiFm2/PeCBaK7fFtEea0s1h2b
1WtJDgh6P8NVobSdvrkLT+vLzjq3/0wGPovbebBEHTj6gx0bTVCNf59if9Q3
i410n3GgK/dmz38mPBK/GHpY8LmgxLQfP4Kfua25zP0N6sSa3ecX/Vx3J/pc
fr7m+Q2QteIh0PBTd6jtE1PBM+qLmZx1mE7wk++hptw4eCbTFHApT4yzyEcP
6F6wtu12mQkXCRSjKTsr7I4MbdS4hBp2kxDIYv5+NEbbZaX0Cr4jUqnknEgp
b422FR5xMbASjCqDV6g6nFElfUTJkGx3kEeksuBoepct6vm+6pWVx+1EGY/x
gS9/nWtMTQTppJKCOEgjkob64fSA3Lt+uogSf4x6Y95VZnKJVhIDKcoCxy5y
d2cTQ+U9jwi/6rXrs5gHJKNy6BG8bQN71MPMrXlJc3VeG0qId3nXdkixELVf
uA+ICCxdQGkEgkAoeTyNYrn4dv+bdMNK3cAot02uTb0a27kR1W27en4IaSE+
jCvleGV+G5j2FX/wFSjEsZzMj/g60gYA+OJVftA8VylcQhW4rDwRhw2F9ywX
Opt5/gDdTRMQjzMwQHhc5to5khLo4fA4p0vrZR5kWZxMg+J9oYOIjTlZ3+gY
FMN58eaJdUY/JggtzV+p8nlCfHu8GJatISomENjO/ZXXSgkpsyPudvwgTsbu
w2OrvE1J9AivC0LoBwavsIt54yh3vvyeR+h50J/O4x30K5OTtK8CfUU6DJDB
Xw+aVFOuF82bYRfi8HH2h5bZEKN+u0VaGztqwDNN6JTt587PT2fjHxxfPsIr
eYEO+EcWFDnH47MhhaGM/HIxFcXgIehD8y4h02a0t/2c7KVSc+E7Oxz3/h6a
svSacnXjZT0n+o+KgeAdlJDQD5W5sqpmcj0d61AXWDX0/BcMtuKCSjIh/XCD
avjYrrteUxZFDQ2KTRGXlvRdbTkqB517iWOH7rf2jRIiIc6+14qngC1isFaH
7+kpTCNdkL5m7j7QOfMqMOQxgwYG4fnGJnMa4QHJcHBEWtNWaBsXf+7CkBrO
pPp9J1HpZKamicqERsXjDONCrayi0GPEytiTff8s26Bha7cZ/GUnoDf8+hJU
r/lpbnyTxTpFDns6AaXBQ4Z0sfgnhvtVfGP8zDb7YsWqU9bZmkrzr9pbtL1M
Bzf0DvLprupP3bB6iLh1Komt01WyEPns8c5YDo6q+4gofyehgN6Sm2fieIqI
2Xi+gHkSH4pgrej3NHKguFPe5JBGOAp7o0EbjjfExt94WPV/I04AYg4RcFaY
AQeE1f0cLjvxcqcjXCkGs38CSEO1gD1Q96A4oDiHi4V+Js1KPE7+vA1akQcH
9XYtsWX+ybNVuaZ4fRDlEBy2DmG5f2SZ+kH9NFfkkfaLoxPPCsFWsOPFAhaF
jxVJ3NSpgaYUeWod12umgI4lBHDYdvBNyqtdHbs1uVXZheFIo2ddG2JPrM7Q
5H8YMauKmZfTq9FrlsSqzvKvTaJNZ1OMirH0bkI3zJObjcoEvdiffXD2YAu6
AC+S5zYQ1hZNBn7t9Jjp5AA+GSg4MalNmCwXn38kJjkwjxYt/hYyUKGW9JEw
ZXdxvH9kWN1BhK00CI6pvx0gTXEPcYTY03+FIUwmVO78C/9WDE+br6BiPz2P
zvwMWxRko4MXp/F/rz/CwwoxVC4/tSvslC/wsqw4djaxnj7gy9mmaJ0b66OU
yyMCksRZZD3UublBopNi5bStpUI4mKkvhLeqTbAWjYXCdAFAFmW+gK0hgZZG
zCiaIlLdnjt+E7OQZn01SMODBomLUXz3gM1J+dLdscN+5JkLdokUtA1Ydqt5
kU3LJ4fyY62qMHZ08BbdDXMJf9TtSzwqVxoeyI6npBel4iXjWdc11Nxz3vVV
WLNV7let635KaE5/BjaeyT8s3wl5gOSdZ+3YPiQktd2y6gLGfyCgFSsUVrSw
dnbEZI5E+Z/v5Mciao/Fwc6s02N2A1UfQFsL+MLz1/V0tXRLC0Jxb1JbIaiB
V/YnOm+5M8JB74mxCcHvGyWwcniogf4OZcmuzzkFKfEech+qij4dDlCIcZeQ
VjjdgX1J2LOHl9y5+9Nne4l27AdJcrDdaqnhYiQaNOJpry9knQf4xJeiWIVL
HoIeAzYYlaElIWYEd2vCbCWYgOWirx0TBDtY9CALT1MrIvkFW6BsngCFea6C
yRDXkyMIIxk9icXhRDQKAUu8wc4bCF3ZKLklYvTCtPRo+FogKnObXKVVR/E2
zPW4GZLJutIRImI/JE5NUiBG6gY3XzofbnAgAsl3A62CNRBYO0ovU/Stlxdq
vr7PcbvU/F1+rC2AHXVSjJKfOkHTNe4OXux1o8oUhG22O/ju982zEzdcwbt7
qGOJMDD1gpcHP0iwHxKQNMl7VHgv91qjHq33XKNFORKCqsdSAvGNFNE1IUfe
FlfPhEueVjMRyCe3io8Vhya/x45ZOs2lVbrba38e32xEA46qI6X52aMMDKhU
TkThGJ65iYRwXGwdr6voPBBqEvZ2pOxzHYhftshTpOLtCr2/CSt/5lP8lkDq
cqNptH/jQE8+gCz40F3hzOSlMLno9f2vilQ6CAdQubiSQ739N9/96GaJuhp+
FL1yQVcf+JBLAS6xwwWi3/DvfuNWaYU3VLzJYEzjX/AF7xGFpQLJu2OsLyPI
GWAUPO3DgvMaemNNoXuoQeSezjTRFcwAt28kL4IQwNHgh2+foUnuz7xMsmG1
ps0516cqbpcqjgldJrHDiJGiL8figJHIVpOWv6app7LtuJYveuZOu1BdjAqH
tjmsEV21EF8WgGl+HIbqyPWshz9xIg0DdlqePRLWN6umT8A69/8xkLts20hO
DEbDMWXuJ7knqSuS+Yhso/su+zVEq24qRnojewaCMZyNSZMRkec55Npwja8q
IxFzJAGLEMmZkV5eIkpdQUQ48zzVBOX1EkCv31fIOCcBNQYB0jGKvmE8fat/
esYSprAiF3OWVCzHDc7+UB+R2tOuWm55XSnOt15hG8PKMBkWqPyU7hlVUmZW
RYG1+6+V/6ZY2fPbELLkit28BAeJY3O0Qi+HoBUDd9yY48sFKdbsZ6+Tpvqf
VKvAIuqvQ1rf6c3ZKcXf9FoH7PnYMiOSPQ2OJtWIqIy7XmZj1J9GGXJiuhUY
QCNjQ6ogkC6XaoRHQkTDQXQR93WT65+d49eaSCvRktjtn8gv3kF3eIHXIXz3
6FcZK9W8A8yCX5CTb+MwfvkrCdt54R/nATdjmcM7VJjMLVU+vHPvJvVI66Gi
oskfTBlj6Q0IsetFfXOijT3+Uf38Y+B8rkktJeDDUuAi1ID2fEqcLbIMJrYg
fZk+4w0VL7HH/XyGIRXvSM3PG9SMXGHsiJVFGeBSEpqcFHig1aeYR7uBD7pY
w2kAjBBs4r2gZ+0lBEin0oMNMi3ElEtQlrhuXkf8Fx5R/306meTyhtBJXTiN
2fh8YWS3tMRsMZW3hKhH52LEEvKZzHq2jhcR5Np+XqhdNOCqREj04zplubsR
opxm5XUBwVUPkhfqdtkJY/0D8E38JaBZ5IOaC/7bWxz90+X823OkoGfrodhi
wrEb0g3rhfX1voqUBXdi/ifIyvgnJ+33mPWTbI0sU4VqLawpGxhYzj/baQRi
HmdUWUJjIqcuPQ/SsraJdaQA1kajsuDDLmWi/Xxakmbg2XxiNgaxHNc4tnao
3s8/EOzfsGgYLeyy4RLkuGmXtxKe/dZBGsyiFSIsA7bDBd91Ob06VAjSq/sX
efSBIPDNdRhJl45IQl/PLeUzBYCmv+d3UFcw0cd0R6BWoDc5hlt5vOAE9BWw
nnzOhsnbhR8B0mjLNdYyyv3Ri+dKLuXI7mIr1ztEwSTdHn8JpgJrJ1sECitR
7ZUoxcN2ug+WI9pt3+5pf2MDoZgtn3XnGBgAj+hWSb2JUxV6ixMXUI4YZT1d
NBQApTxHcq3CHztka46ip9+BnQP1eyMyuWBR0oDG9y21mk6jk5RGk0NFNLCw
ZSFZSKgx9Ef9ds125JFnqTmyr8WM8BjOXMA9hFUEo2yRl1R7CqMNfZMLII2m
1E+Rf0daCe/4HGPb4FduBrHUvlucGrO3WwEYpEvHEEEymgJdlk58ME2+Kd3X
bFfyaZojHA6x+6yzYyvrEIptuzzuAYQALHA8E6d6Z1ZOWpsVTA+kOruCJ/91
+k5I63muN30NVjVKpbbxkR6TBtT6nXh5H4Zr0NVGZlwWLxL8No//IlvQD3WW
9ZWh5ePkP+tSA+MFFb3OaKD+EvEToXvAKiocqNrryZ1/obbCfTVoguMjSmI5
oKWn/FFl9ouW+s8KRJio5mVehneHJukhTx2T5i+78K6bFMg1HwtnucpbvAJo
KlqLOctBG+eR9+WhGOeKogmq1JDsoYwRbZ00xDq69zQR3CDtzwByVCv8UEgH
xSpGvt16MXrZ0VFAbRxXNWMhAcispM40RRPbD7iXQn7NYBsLNHc6bf6UVskp
SYAUiDxsGDTSMt+mttgGw8h0poo+YQfn879youRGblM61GQAw0Gwf4Ovu9pJ
qTYfxFW3Uppk0a8EGKznb/wt7cCWXKEPgdebDQ4zwVmTAyp5ZBDwCUdho/il
s4A4yWqOphidp/EJMaqsAgPUhur+cyR107f0p8IFOsCCWGHp4eQ/SxtalacP
NLXKq9RMFLDNyRawfKcbP55dVvSoxB9zPmzVJB/GEGCyMDn5vM3r1KVUklaV
CQFHh1FRfdffnVGts8HupIkQCkPBvYLDU3T7Ub702AMNIFODop6T3rfNhoJt
O43aK2k96kzjPvShI49NySvN1tG9RvAivpzO3UnrBoEOizSGHX/7HqWgnqnu
VjqZa2k9/rSoBieq8Hftv5VXQyIX1u1qlXjTSeUh6y6fOypNNhmCbrO8tSib
4pcB2EsXTtHKIKN0TNzR4EHyneOCmjrRNVSP/V88eKOZxKXpRkYbbIDsf5xs
NxfH6K5FdrEzu7i7qx1UaGWu/ZUVRp0yenYTprNbAOXaiKEDzTFXLNCkAXzz
Q4T4RqKiaeXeBNElWM75iVyXtrbkhc6r02UPuewsd244Ig9+iy1y22EH5Mcc
4ztC0VRE+gVwRM5iPTdf6HgDG+tKhffMPvTMmxOh/uBIvxO56v6lEsUbDhQo
4O88OK1OrcJgXvBuQCvNP70bIhyMjXHqbX0vIeeXl9Y8nJcPkCKw56iKXpIs
diNheRgy2rHDosIIeP2kolrx4o5TKeAvuWmnbi36N1D0DGGlYw6sIJObT3yo
GHcpmiaYwxnYFhhBVekVNXrbb9KgA5CcYzbJQotNOMvN/umb+ryB7ztv/TCq
2Is9lOhynZJ6iCRgmXFvT38JPrxuL/bNjCuGeesD3Wkb15+SqwRhtmT7cFDO
JMviZ5PBaQ0Os6V1OtZmMigBBpoO2UOe8a8lLKLw8uhYx8J2m56sb1y7mm43
iVfP3961KsxBJdAWZg4DNspAYOP0qDbknXmf3DGsd9z4rbuMrDOzycxtEsGm
nl+x1JF34Z0qZhxNRFEkhwXryFc/N10sgfnFJfR4oW4H4fS9LtfbC4nNMj9g
S9VkM9e3V2o0H/x9GOpklCiu6HB0HsF8l71IXw9Jter/FUh1bk/dzKwyd0n7
vTMT+tIdB+UhvpHKw6j07gCuX5JcroVwiyoyuK/nuWwbIt6NzLm4qIFCuumr
sAWM3mFCjo09svLfiJxqnIQOyiVPNR2bW/HJAaqXYBiL4jkFG6c6UWSkYZtA
UcoJTNbNRlfz5sFa5LAmeKtjRwUU48QVo1q3PRQBjRN+QO6BwHfcD9SWqSPS
SIGTJdtzGu7HWtUp3tfxaUznsMeiSJZRoecubf2/8wY2FLaI+IzNbmtpcw+m
Mbg1BcZq0IsTBdRPgiSrm+PHWSLmw8czDez532zFezrkrnFfi5UvN32uUrRe
jHpVIy6vmoOWf4YaWLQMSocVYtYI9ppsTdKKuiPTOTSPKcJf4TG2yGWW1Nzj
R50H+oJML93PPzngCsLYWuoqjR7VU6BAbwlE0CkG3OWBmtEi8mfruWu87Dv3
KooUF3GsIiLUlqgga40B8iM7zaaisXpKBPQd20TJggziZc/My2GsJvyPcWC7
PMWgiFALkypLxVIrJ05IsYAvHlQSueJOoRXn4OVEzzxBj2QpO9hge9NI8Hdf
Kli65Fn46/sTZ0FHqlC4tGvIyOSWPc2cZ8+hutgV6aaGpe3x2iznbqnjgxEQ
CD6UvFw+mhtEq1LIhqALpygUUCvoeW4JM9zCc7JksgnO8mljRxjVM5LZYooL
gVhcMSkWOyAmsDGp2e89Xzgka286/xFmOXkLDz89IighGbU/dTgpFpIXgmzg
rjF6apBUXq2bF39oDQPlg/b1X47WTFzp2fmO+eKJ1zPtSkTSHv4Enk7hQfdN
3p9PaUWVgPiTx57nxLrEWqQff1B3BGpTtuqdPpHlOH9jY+mTzUzpahiwLrxi
8+cEXAEOnRXfzz6y4xG+ThgTrIUY+uNrmZfYs8CeldGpTgMfNxXVCbqLovVr
VGieBvCNMDXpQN8BJ9BOhPmIgNNQpXqvYkgfD2I+Fi+DBaJ4CvPJpV9nok9H
J0Lk2uh0cv+BXDL05aUcd5TzAzoaMC/SqWaNDR0W4tfn2RE3EHndRcnG/Ndi
Qq8KNCT5W0OD17JySHHeUfhYPtGh3+KwuxVvasgQphxjyz4SEVy+w/0U6wT9
+l6wjlGrdxT1bOKVLxMtC3YfsNSsFbXYN7BPXoxz1WmSgAmHsraeaWgTKBEX
FX3FOf5UYbypl9Vl8IqdQmihrDJ6zNrwFPmWsN6rZKPkiyxXJohp7kCHGhku
mRnGJsrqKKsbMNIgFEAji+o0oFoowE2w5ddwy2Fu/BwSXX9R49gw5pPart7s
KFTiXky1qbH1WHhCyN4XlriPoM4ya3+NIsLOfh/09k9PzzQqCN7rNUo1+P4k
dqjzZzS1zsCcBnnq+arw9hUYCwIPHdTKaOE1OYvqzRYTxdI0+/XSOnJnCVxy
oGL//UmettUCCAHE+/Lv0kprWXhaoKQCTlmenaxtVAcZoLYFy+DUbFdMrFZh
LZvO6myx+CXBFJXt4sllhtX0T2F8/8SsK9BsKHcjeItJ0+9y+hLZsN0CAKFn
PnjAKD7cViDmSfphl5hBZw8VTG8ga7ks6EIc6iEgoUbEdwhHZnyds17iB61z
acF/xxR8U6pp3Gq3CH1TeWrhe/Rxl8ds3He4aWSSGuWsyPbm3hY5sN57kr2y
VIxcqClWWqPMoZfpj/maAFqKQOqNfqBaZSU+ITK4wwavoOVbdpnBg97egPMz
h7/FyHdXsEuO39Re4lK0QA+BlCB4CnHGPPnWRSHp0kGj9FpP//OiwhEIcmlj
zm4zTO2ygI2/R8uV73cquK+Ea8pcjrQfbg73yQJcCETjp391YLGhPCMAY08t
tgmKLEkqudGsH3K76bDT6asQp2DCAETH6J2kPR26BL5RK3cAHOgbjrDZyheK
1zdfKmZHjksaqG30vmL+/KS9Bwo/PFJ9jxGn3ztN/kDtjQt9Rt8pX5XeXLgk
DvlQDMN7h5tGz5ik1WtKY25Ou2JSUijOg0aQ2LbYRfNGqGv6QKTk45/u6TXH
9EzFnNQsmNaltCj4gOnpNSnpXLJFcazKNoiMGypp3SmRWioG5KQ/qrU/WQjs
bor2YxgytOx81ZpN7QvjgcK1Bmiic+gPLdLMGu0vLH1Sqg3rGKTH0xezSYEy
kF1C9sY7P4DTQgnR7EOn3ZMPtT1GYW9CesLhcjvesSRuxSuKZ5jwaP0kPqv+
S7EfKQ24bhwubiRLsfQ7oa73eVLJVYlmNmxZcJsfPy19+OwsMaUd/k/GHmRj
uoO1Fzc1aMq0B4/YpE9GVj7SfTyn4MFpwuBsprFNZlqGj2NDBHCCXmY9Rxk+
Q22bCgiQhEp/UuMWwetpnHMZy/FYb02apTAQxIyC6A7Uh0nT7TQfHpHOnHz5
rG50jpX9mLroYxK2B3Zdi8SazdtbGbHhBaHhJYe2e+RyMXOooy+ns9l1KlgU
ch/+KuAnnfkqVcx5J+70rLVIS0XhF2dEfpvCo8hK43HwynUCPVBo83YdvLSi
o/IFKRhD9l7EPM+3/W18EQYH2WDx8K4mXi0d5rcc12nwPEdbsyqZwabTmDuZ
PnGnvbfq/uXOkcdmBvboZ5UJdsLHgg/o2gUGQJfmOXMFdBesGf/JnaFbm9WZ
WoOLetY72vttHrF+XTD3jQ5O3lHt53l4ac2YePo89dKeIlOOmqDSg4zUu5za
Symyjv+fUVMXsje8tyqT+rsAS78T/JFcwSHxysoihckL08vAfswXEFP9U1M7
+aEeC7oJ1AC5PEgfMmu61RYjseOA+UoOGpesc9CTK+Yo5WN1xldWC1H8m0An
O5lvuLTHf8XigfuY5+1CPewA3ph0gPwnCugsTIKgTVvJL+z0WW8Q08ff6O4n
VrKYfe8cCeFZeiiuyPD7P1e42aiINxtX6f81Azqf1H6NfjL0M7ARXTsRoOTm
wSSnr2T0vtd/tVLJEbffje3VNyNc40t+tw6hQ5uRLkB3shdgcNjVglYVWDbM
nYSp+hoI2VtXBQNQFDZxlGIbWCeU8/qe+IL3OucE+pEdsp0wGNxPLAyWAtku
LzBW9E8nxFUe88Qxfpcy4sc+4cEAt+y9EummMxW3gBlmANAD/6F8jdVDWYG6
zA2EgfyZ6BbnwbauEY1X+lTB0fl/MVdlFjp8Rvek08RGtkxCLYhJ0AGFg0iT
UM5chl9SusLEsDaYysTuFQMRUhqkKB7vUwde+0rXsgpLyA8K2NTZ7sQ3/vha
Q68xtUMbA4dLi29grI6ulAz5n/H3awhrkopYosa26BqTa7uE7/cc0qJVtr89
LS174aSVSsykb1tZajsOu+8ql+z+E1T2g2L0UQP3Q1R71D5VTG+PtMiA6hP6
qxrfQKQhgmL86d0KjPQI1hJmidQdCIlOT8MuRqeTwUmRoSNrjO649vdtb2Kl
xX+PLsIJrk/ftkMl6aPgH+j48hyRGQPX1pFHoBNHlV0Dw5ylUIKYddzrGgjB
BRDjgKP76eIDyp4aUMHjP9U3jqMekVYxJcMwVMmrILsgEcHNhX8CnyCNuHO0
YchCbdEAR1QN1+HfTbTCw6yjyiNLlB0IpGzaI9CdCdSJkBZEPjXDSyiXn8aI
C3Yoh5JjuJlF4hS2TUFUIEdwDOYegdU/CWiLalw7DchLOoAEL4fJ8hZW90tq
oG35PMjCtQnSITQOo29ITh2gE6dkoVXW6S9zauF9uLAt25K4P8gjkQ9eBR22
S+40blqJQwv8M5ddaZM0NGU58wOknhJee+dyvFc5x/T4aupuxks7OkqYk4C4
kbIjYsAvM++3w/oP8FYhd5eh41DB4qdt1iYzA5StxYsfuzCBF/5xs2a7CtJS
GHSSzIR5o+SeBdX/XtGKqE6Qu170Is6U1Oah2iwGLJPM7+1YIFCl9F+V12U+
o6sIWzyMQ2lGv3sxofRkTvahlMEZgvZ1ASQFgqVtKQykbs2gV+dUVTSxJxaZ
KQapPY2/aObNzcM/HHOdvJet0Xm5+PSnF86EedOAmqOZSa4mCmrc1pVNkl1Z
HqA2MKzwtm4WlCvwQWlTtkNvFESbIF1VtLO8pg1SFS6YDkNh6qC6Eal0BCb+
lJoNpV0Q8t4M4cDGO5V4Y8UWm9T8onRVF8wZl0Bv2vheWapLpNNkv2mh+frT
xMLCinmuxFdz9eAeUnqJ5GZoyD2lR9G66bc7slqI/vP6PLLwcYxRN9DTWRQe
rodRKfV2QxUX/Aaforr8tId5R78Cx2YuuV/n3QR3rCVXQHKbKfKpvHpcg/IJ
B33hpAJv8HpdxbLNwhxfDTf2kHGHqcBT+bwR/ewck1VpBJZnvvfutNj/XFWO
z3+k+c7u5xB/C2ZWpq28bhUfsYwhvS4lxXfqzF3u64lqv0BsUcEkVi/q2rIm
FE76mZJzWPD/q94WRa0Tgo9esLQ4LMZraWBR6MxyrrvoVh2uBA8ATYzLMrzZ
2eLz7Ng1Sw44D391MBNO3Z8BXibQFpDZRQN9EjIYCuHW1C1fnrZIcld26mYq
6OZ+640QUf+oDddks0O3w4ULDVnIi0FP1EQB6aWfQnnMUOwA1hAZECjPl1t0
8qq9rC/HeM7Bs3oWmdfKenvEN64O+KVgAjEUv8h/OrPZga3wh/4uH8ZrU7ra
wCLrcoj60anqQwML5HWqQNbyNSQbn0kylokFz+r9TBm1CrEZ5lchPSlaUv3h
kp3++fmlELu5hzKnDQCHgxFGBDBreY/vGwEgTkDj2J+TCtdCJVxBzXwKteYk
8OalT+VvONBMCQA1fxBomYh0MbeWp3L8spNwsneBHW5FHmuvEESeZVFlvsvf
otQzHlVJ5ABBKNucBlc7PJoh3XzNLfdMrOe3M9zsEYmHjRe2UEFpXotw2mWI
rEPweWCP2Iy8KjoNYTvtxHvKSSzgQWn+5QUx0WhVBoQ0ArA9fUBNadgAV1V4
+mjcuHQqJ/EPdd50lU1+4koMcRgYg3mLn5BwitifOeX6ltRkWPmb3j9Tz2X4
7Ry9pr4wiCmGlNHpQf6p3s0oOr+Gd2v7KQUhqA30Ynm7LN5hJKKRhYfSLRh0
vG4oKvpExmbYam66VZA7nt8RysAselqs6PsaZIhPJXophwggStWnv7T3Bf5A
izfj4mJQq0Jy2j0HDA4bj5T/dl7F52QYVa3g9IyIgGqU0yeUnxLvTc0ik+ws
thBSiDMntapyFDnbaq/W0qTAMjkn/3LlAhr4bPO9s6EzCZJW4AevRSSEyeG8
obRDKoT8hWeQ8uzC/Quz0pXBTHrICbBdww/JnyCr44YmeYkGyYhG9XvmaVmZ
K9ngc6BcyXvqydoIEQovgTn87Z/zt+e87OT8HqinNTBkw5F92K2sux4QM7AC
+t8f/9RG6rdBDpVbfUJ5JG3H/hcnRUEygtjwOBPKSoD19vjl+HhlSL/iGsJ7
bcv3GVfDvWfnR1pCWFnWet6CdfiXzV3wFYBTvAzt/f3xSkrxffVpIdmuqYkc
CLxGDYM+B4kZrdcoxzcsJG0qCAHAg0OoWAiPEJ20KQta8CikUogUqbl4zn62
4LXGI9dEYzhgzDFSLgcO4tJAAnURHpE4ISGmsLx/99dzjGd65HILgkxHJmTY
6Rxtk8qcT1bVx+8FeAt8NvyGwloRZnMxKdzxKyOJEI7t9/qgOUmwbdhGXTPG
UrZ4fipPKpcQ4sN5X3lJNCNexIHFoihrsHVCinO1y3AirdGP90Ty5e2Kz0N5
POZvyg6Qp/2nGPIDxSfQKEbGZxV14OVRxf4pWOmmN0xEpq/Q2Lwqk1VCSYH3
xqcItF4oMEArS8InDeERNxeHo3MohoQjFyG/bTDy6qmcGctQA21/GYpp7SXg
QE6/PCHl7SKD9F83cWKMHvPV+CviG73BXSvbP1+lPq+29BR6MkLPQC59uAVy
1Cgs6m5cyQraMXrPpW6rp23KzXrHktRi5dWV2Zg4Bh0ZkPIPjelfR6hS11zs
46ojt7q0kiZU0s7qy5IqyiTsDAnPE1QF3JE0eC4kzXXohOGhfJ1giXNmG8mm
GNXlWhj8Hz9alScmzkEBx25v/69rERrkYW3xJi8tgo1E+VBcwCunDmh0FPR8
SooGMeMbMcmUouzHM/MUI6S5j9x24bjryWuBXP5CQrW4g8WzzrZ18wx4ihji
jMHSQLV2JGd5rv8LJXb/qqiXB2ey8mLGQNhFxLFnRvN6EPPf9gMZijGxBAni
wK8+lr9uij7OvYDKcf5wvMvYc1W020F1HbBDwZcTsFqs3E6AoKqU30KLFqgp
/CZ1nsiTBsp2w3x0qxUqPu44fdG88IGTwBVtZtsjYiV2OSYJU2MrNqgY/cps
VT+Ih9WU8oBWQP1MN/MSspmZo60tRkKvNnX4Vz5WzgxsTA+kbSQIPo4kQR5r
VrkTSc/4unB0SSTrTLAoglFMhviW1nOEdCVyR5O5+6ZqV5H3MUeYO2S8Sp8J
ewST/y/aiFWKbX3LHXVnGlSqTsekGjw/GF1YWsQ8u4L7dRByDY+quhWnkGif
kt0uJ8VO/qqOOvkwFhaFa4WLD17LqrKhRdppAg3RhscmxUwMAKzFj2P0ZZI3
dSq15RK3aKvEx+hmCzCOgH4cxtpkmRDCdCDZY2cLhXyP51O6hW1TB9CZkpkQ
gGgxaj7KKkjzrvoE24qTtvwCfar7AHevUvBtjNFIvkE12m4RO2hDN2iPwd0Z
TAkBqY1prEgtFxwSH3TLRvbWhiyHVWTLhcNxVcuFlFmNzRE0EYyTqAfQWhg6
luGITLwxTmpYrEVvKmFxgxwAwxJqZcMNKam5HH/y8HR7qFcaQD2BAA2lzkny
/xSnuMQuQtb9xURS8be8ZnslzBF8if50AZhhy6F2tBfJJMG2hj6DDaGXPKER
ndgFv5ycgijxUMHRU/71/um/HW9PWOsoOGCtqHmBXb53jybT9ID1tHsv4pOs
smrG2bOpRI8lVJ5yhEkOqCzGjj+b4HZZm6PpBe7BSX2anTzoKudaLWGRInn7
Ll6vHWHo6kM61XwK/0aVObrtovVltVvudVnnI/iYCDpLqi8G7Q1OSR6akh41
64H2oZWBjsl4pGmAYLYcuvCdhYX1XYd68rduQPSs5UJONkk+m0sOwb/oCIev
maeSRMA6YL1RvSbVIDBRi7AFu9oUNiO3UOOymq7nZ+KsKVqbQia/rZJDZUpJ
Ge61+fOwJNkzLqhAcmrYdUcgA4MfhmyS62MUQdLdpDtSRntIZKvnQpiV9GFi
hfg/GWRaEUQVBBl1nnx4z9ZRY6GyUviuL74DT0ICcFXdEPWi+RJY5FeCsT3p
Ai1uYoMQRmfG26+7/o5rtFVyLE3L6Ai7U3RepDgH9LoxMwgkb5qbyZV8UaVu
9GXv8i9Y/yaql8dQnOUWH3V3fYsXRgZWaKkZpZVETvhsm3Qg76rcw/t8w0ch
BE8bMCtLiaFJfITX1oSE4gW9jR4pyZYxoIMyIzFMLJn1PnK8T6gzffpoZ8mq
2Qn+0BgLF9h9O0tvs+XSUxhLeR5yPtKux7MyPFyGtQXETnNIr6WN5UQrkOj9
bUj3IJEElpWSimVTAsDZwO3Rx/5fRt6tMGc4B5KB2bpTid9LvZPxY2d/Am6m
IO0toQsiS1NGj/eSv5GdwNccNbzYbWMtulbdHVEf+DItcSpYwNPf0Yle3hQR
hgs83vijw3myk+pSLCi+QL3WHfZrs/xb8miSen67Z3HHH+o97fgxn9Ul1/Vq
QtXHrlcOUeW+2qwWU0o9f+RY4qDDvJ7Xv5KgC4GmnoRJmKMdxhSglBA+X7kq
kUpy7nvpsYe5TPHrFhqiwxv5/zIimGXnZU5H6HzuXU2zqRc6pdQHWEtVIOAa
735A3sA0TUSTK+AiXspuygWNjSVkyDPq8rJWMKy4LjW9RlFGP3J7+wvc12MW
bfy54++SXx5Tg4tV9zOBQxyECj4PsP7QIwDha6uAlTqimfYx7j0jK50m9tiI
JenPlpG0idCfNW4R3uwla6wDAbPpVYa0oNrD8b35I2gQYNyZKS6XfRxL4OkN
E8LOKaCqFn1L8Dz6oPcq/4WCC8NJcCuQjQ85izV1COM8WIC0z6o+p/fW8xY4
hOAezBwLmOd8RGHOEnTB6uZYsENJ+7Jho/3QTTlbXo+/CLOGymIMLbYk0uWn
liqd2V0vSQ9uOPCD2JuD5gFHHwXmjvzRvsk8fw1uzFcz9S5S6qDgCkWWmVQ7
HpQwZlffYflUXCrZIUQkjpJiBUYvjEEbLAUJuASs9ip9k65BZ+a0RaHojjI5
0xjNqYkJ6QHxQx9+NVTvjTyZ7xesM9PgVzLm5dYkNjLqvzHAKwySsDZLH/A8
Puqnx3xY22zELzxRnOfk8sCFBTA/3RfJhZ2O/A1rpZbeca3/BB/M2OfMqery
NA+Kwjha52P1ty5SCLNo4pJSEXWNGclotLUL0Uva6a2AtDJNlJy+rtkEExZV
PHhWEbj8omPjIHi/zztepkw883xztuWBMWbPjaRVowP5ribxDRD53eFphZJr
+JNmxu2VUvK/DxIJpaGHMlW3BvEbkor8njEX78+Pw3hwqZNcGWrx/NkgTydr
nNTpXzzRxemMx7j+489djMC/WjSUJp5D1fV4i2RoXkByC9Q+lXZlj+BKESYd
d5DkAMDxwIC/sItfrddiuR/ZMpQ8CDyO8wOh5P8r/GLUjKQ+qZyQhXSBdeQ3
scWMgNiwSAXvpXN8FahDiJ8dsDcyaBXzhuyHCiFvduDNHV7hhKyF2XjKkwqr
0m8MJC65sCPBgckrfe7YjYZaYIMdi+FqcIg8aN7n4srW1KBWv+yh5UqhPPT5
wzMCsFqdOZ2ILZkpXOtLhRhk9YSdpf7Tn2iSQSLwiWPu/8uK8JfWbAV6CmHE
K1f9GVDHd88sMH3Z2BWMliTA76BwXUahcx8Yg9keOCraupge17Jfg6Q2/RdC
HA/ZBk1Yv038JvqIpfwx2nRoaTLt/YA5Tq+52efqXZRulJkkOtwe9ULW2HaM
mEt2zdGWd+FCkcXe/R4JPU2MFXgwtHx7F0tJfMJdJp0Kch3irf9Qa0Vyfc1n
Uyq2ZYhlTT488c4AfSvsJRUCueKPt1sZ12lveCdfzRXIUY+5dYxBRROSbM67
okS+WIeEZucXKNJg3leOcjZhrpCTtjCbmw/K1uXmWnHlf7pTy0oIDZZPLvA9
6wAQK4yPkSlHPoZQbJVBIOnA3/91L6d11Hg6W3Li2mXXyefYi2HV4hOt7dFS
04iSjBwuQxUkl9eAyFUQkxsNm8V2UMiPYbTd72W56BRPM0HU4VxoTq1FWcys
sQkpl4NhGMgrroBtzW0Mo4BYz0scUAuSEKbYNUBq5+AlkzpE1eLMTGt2AjrW
hOd8ATjylBnwLfhXX6Ayii6EuXufQOS/KgVFhuIeosdQ1BRftEHfO9qLEpMS
5SKcLlk+LytsipehMZxHcjcHf60zOYiWxb4V8D61LBAYwbJI8rbJpPL8zu5e
7K8YQU5NMo28xrA4urRDo7BWAs2vR107TQR86iLX5r5G71netZS+iJxoBaYt
+6RbunFBkIcX2nvNrK+uxbjP5E+k1L2bLOBJWZSm81HXfLOxJmgWGK38CqYU
E+NW7W6yF4tAnyYVD86sZthiufXHI2btnXXQBuaBpLYVEJE7l93efgPAfbnh
nKSx+LtRyjnWnzN+r9Oi27d66xtpUFudWYVV5Bj2GgDT9eZqJc9LKmcSGIzr
Bvm/8Tjy35lS2NvL5z+TpyaFj3DEWAxYqfhMhgQuGy1cnAoQoM93ztPYTmbw
TxLR4US6WWP/Jz1FiZ30FjWbf8Q/s8tKkJRRJTlH6auKEk5Bn2lPSoEmVUEa
zzQRMV32r6GVus9uNyJim7yrj3DuwZq8PHfzSzW99AMWYRTcHPeNHVCoQEwc
nFmRjEOSIf6xoGki7rE7Yl1S28zDcFno2y2gbZnevNzSs95m/CZMSQbD8KTq
fx29LqTXpdj9eXSLsbsS7qDMCvmM0a3ocyKf38Ivm57mZcA8vDaROCZMf2wq
cQCb4OFQDg1HTeoOyCU4m3RL4/dzWwZLrf/c4AzNlcxqdXicz8FlcoNQewXY
1MVr+Vm71ktdNFT9cKcCX1/5JppTlHmcUy57H0nrQHmvPJ4eHU+PajL3LY9f
+5u7KTK/g9zlt5WNOczw7ogkAIPukh04/NoXMG5D8jqblLI7IrDZjXQ+aR8Z
6N37frdmNX8OtSmGs+67ZL7XEDtzFNz175msyfltpKqG73H1TVarPfWt+g6J
JLJVdZf27iabz7hN/uAdw94Oy6Ub+BwKjVquY9RLkn6voM3HibFKM1M/Cti7
NR9iA1NYbJXuXfSbT86A2HYa9sFRaTUbUqtJUmTfxOqEXRc/XmqcqMvw7BMl
MJ3p1Svd8NZhgZ9RjWdx1G96XTnf4Fnw+MEloA8XkMCsJ3GR9GQbizMV4oSS
8kKNP49De/egqLIIiMtgL3sOXfEB7aO2o+m+JmtnePu7+lCu/H59oxKAcidH
1GTVgf3T1ITC5WSXAC/Lb7bI6vRiFPeRYnfMrSUzXSPNK408M2rhooIZP24T
0nY0htgE7KlfsPGYQHOUptMnW9vOjHmpnfrq4lhX1P5Mbk7/d4wA6Tbr8I/T
nEi1/ABjSnqrjgQbge8V0pbz2zqA+l+mag4gfp6wH8QZKBheCQ0cRxKB4T+g
al/8qoGtKJdN3okAulcliNJGL0YzKfNaTBrd2OQhOZLoUPeSMI+z0WJvoFXv
dbJO3hERncSiczzGl8g9wvOlRd8Fy1oAL2D83HbooU6Q7Bhqx3Oqke25hBFq
Oaaif9s9PmMAYbGJU+KgJM1xWSXT0d1ZGDZ5eXQ3ACB4v7Xu6kh1ZMVtr+gx
Tnx7/iof0zC6dPvNMcnzRB3Qtxa9pZdT9SmB+6DfMiCbhdIB1Sv80afsF6vf
SbGPHkPB89zAPs+O+1JSbbrThgeS8Ne54G7lnIJHab9gcRP/wOxPMpTw71HU
SUskD6s9WayZQPGluiQ9M1mnsysDB2+IJQyrXVtbaV0rw8hkZm1IBuzPiRd9
eW7L8QeFEiBZLB7wD8MXIBY+ILda3c6pqt1DJhdLd2GJxmo90b8rOXataWmO
/rTmx0jPLcQcciu5RJ/2MTwEYEbqZcOKIEu2+6wVGIKZkS99lTP+yRdOrHq+
ooNozMaFrbAkj/L4VNSZvdj4xLRRkk2QSyBQS99j15U1a2UJpYwv09ksFw4y
FZb69GWL1SC8dajqTMgyXnoa2HuTno8qKp/jjo/OTdihth4tBWRquYvud/G7
8uIrSQNYaMjQEao0Jqjy+Hcxxogrq0TWl3+UUQpa+1fdKZ0+a5KRBJuNccEQ
++SWYNEMYaA1fFJxHKAcxktsOOwFf/tHLx1KbbAWZ/mWPbowAROc92GdL45S
g0k8CNK6dJbDRG9iRyg/bkRPFaS40ldEoh2otxx1RqZN252JG92CUmdQHRD/
E9cyQC0h5t5wskL4azcGiX6+6OrDtmi5/QSnUH6wzDlNlgiagjRNfTrKhkpl
s+sgWI4nGBrev1iXJpEm8NWi5g9mBHrPScEDYrpQg2esHoX8nr6V3WvkssFu
PYc1pDrtMMdn3DtnJLwm6sR17nlFYZEYf8cBZ7Y4c884TEjj1uHaYuBfQ9TV
NNnbL7vCnXXia50EZbyTSS3hfqW3eKz9wLq+zH5wZSX99FrpI7gsUFfaLg4F
sZ5QnOzbDm1cO8N6bOCUrusWz2i07K0DsJBgm32bFAHjO4dmuFtjI4zHme4g
T6qabaP2b2i/UQdJuabPcTglK+dmYsOab5tfqw8bMa0IaxfPOhFaYjn1P93s
YGBwggQQTt7jd88wZbMhiJJIcTb0ccU7mSv79iw1WzM5WPUU2GL1z5wzQnhR
f6PrS4JqKcTBDAcYehocfJWuOCkhInxk0fBwwkuZClQnPKkmY//T/Uv5hVKa
NiNw2SnPde5K/rcWzTUDtuSef2h1acdc5JM3iTa/U8cEgVrE45Bx+Qu4+Z7p
AxxXgKk2FctEQjfds2t241q35si9f83ruGAanHMKA8W9kBd1cyE3N6TgNZad
m51uJSht2YWJVJMfLBSdK1B7v82LdeTb7+IG/R70WwNyTvBIYTSw/8xrN476
fZXeAnRBP4khXM6iwwIFepiHuZEBFlftQaZGpMGT8E81zUojHCkm3EF9Ov2O
tm1HPMHx3n94QZQqO+QFsFRIAfTIERLcXCSWO1WqdmBjT+v7Na3vaz9jfOe2
pij3NVlGMPao7Va2s54PGNEP9TUaAChYuYSFQF3LYAB+1V9jVpzqzZGl+J69
XJDiulBjemsxUWv6VUBusaOK4VsZbDaCLUEVxO3KEOL1g2F047sT97ppNfQM
PwgsyOgDRXC4x9vqfao0YxCvfy/pF9s3vnTwPhzlVh43JfNegzXCUZdT3ORc
eBs+ACRkpPf8adFKR+L+4ViMaPnpF2YOqrsbZTQWdAVodoWEPMCnbzEjYX+S
cevlu2t03o3nHDGjhgena59RIJ9zPFI5FpuL3M3q22YDSNABs/wEVFzYQDcm
gWH7761CZM9/69ndCyCsMB3UicNiw9/mgBRxHdgXgu6X/LvHAltWQkiDtkmi
2NeSIfet4/cTYNr6Rej072/ACZJmL2qlLBFdcW7Zq3xJMbqDYZOqh71idoAE
TfpWhyohO5eMCg+9T/Jd/cCDv4MJoCfgnp3Tue19KIz4UUaRu+y80a7chwHx
Bgbkpc9xiyG15JotoA7gzpH90kyarsBZfT3w99dfuwxyw5tGprkhHMuPWtud
FSO7Unq919IedXqVEIB/Y/Pp7Et8n73IMnYfpu9vCYV7jNXTeenpme965dwj
CSlbGLwgRWzTSbwf6ShYxOEjQ+lhnBXHsTJCNSXaWLCxdt/XdXLbiqyHy5zH
oO2CZAkbCwK1SoFhUh9E2G6BJWKKCoc3vGWB/8wDvFxhUMaGuOk6A8qANsm9
4roxWn/9BN/m3BSqTZrBT64tF/9DdXwGvO9hw9Thab+4M9Ud4LXNsOikRbpC
VwT40HlUtCuqqb0Vyy/ZG2pXyaJ1edmwkXAB0Xi5z5b9d272erhixOVWrPZo
XSvVaHO3ZimIMe79fEiuIyzvkRg57KKe3US6vgmglXlKJt3Gj0CAjW4Kwn3w
MWKxME2pwiR26DGhEZQmJ0G6UXRY7izp7IVIwfwjWWF16Dn2+Qgp5QPqx/3W
YSAYhEFH/eChOMLSNpEHBYunLY5gvAcWqTZgrg3+k3hwpnocQX/W1W/gDrQU
8+psPH2So6xod0UsDJPhldcubdXjGCtyBhTfNr6WgRkAt3pYFT1Chv1yor3f
p9PTS7qN/2NHowQqOJKaJmxGwFroShdKO7Gk9UQAG+HHqwurEojAd+P5QNqy
pooLan3bUuzzqAMdowV3L3XBQVB5AT3DO0hDR6N2UyvL5J430d4tp+3mzolK
KKWBHkBTj/5QU0jyzterA5X2DZCAhoiAFAskdpY63duIEARUMNbwHkMq001d
lKVz6qI+3YzJIn0KbD7IcT0MDxklH0hznpKAgpiQyeXb5kaMuLKn0t7WSNYe
azJLDLS3AJCkOVCf6x1sTDn7kYGUEVmHYoJDnxkNzjcblaEysZA+fFO9r+Tn
BCE8zRTJZPz2ku4V9LVjYUwecOhkM3zGB/7vCdjAd7PP84C9My86VddR5mZE
mo4g+5tSR2YsFXVJaiw+w0sZwNfEeh1b0WaQ/hDp6+g4XKTSfNYbXmoVEVyu
pA7mjdAaaMzIDryKXRt9pG/DPYa0C6bVVaSmfKVosrSkU2jawlRjpCIR99Ib
tkshTDd/XRydhHgGp0mj7BkxbNhnGxlGRQOd6Ehb6pvbBT3C+ycJJcwuTQbb
6ybgkiCmAKcFn0yqOmA9I+RJga0YYDEaQiiJwBtvPb3ueOmOY/gDT8bD8NuV
0D7758rwyBAmJEHMc7V8a7NyhFhIQyMhFSxk/faGkXXxIWCBtGgrcI2TRkvB
3mcSxDGm7B826XvlFOp9JRAq2983uOQDa2gRmW9E38Qt4l7UV26A+CmXUNBH
G0tvvr8kLeXeMYcbaFXljr63hl0tW2XtIJOqcuslCIRKVtUJwTjco4ON4Lyh
zDFjLsXMuKKq21dBCiLuLfaYAHDSFqwsKey3x2y1EJ8ybF7XWDPihu2OJR/S
FmPGP/OnBaPXn3UsZcJg7uiX/UlyXvgVznyTeSYk3sOEunPSaO1MHGrB+C9C
V4Ve8C5WJZYLSDcl/CmfJjpKScEoF1Q4KEZ+/RJxuUPvEGPJkbxv/i1pJANk
4MlntXPjew+xmXQFpIBRXm5B7qpduACwpYgnsZ0kk1BOZKE3BzNUvDAZR018
rMG8VGQ8KutRtSza1+f+vFRs73VRNtS8DF0Oh/nBrfp3z/DJv80MxI65MwHW
VPnFz+cT/mhK6q+Hpkpm1d1GGvfgOtkHRzOFD4iet4gWanjKn4HW0SzHWQPk
2Jxg7vICHWEtSOAACpvUhThsdpoYqMpPwqArznmv4DPg1C9CXxEEthgQFcsg
1xNkAqs96AFLsaQOQCGYW9B9xypVFAZ+KaIHXQ4QgZ5Q2ie0faErOub4dES2
h+jvAEFfoknoKvlqBFrAdo+qXwz5bdU5mQvkwqUAIpbdf/NldHdDpHqBF6HY
momeZx745ZY7tpcaVvnsy9y+IYrwGJLu0A5Ex9gS3z2NC2YXz2ucPDT7ceEh
dJJe9hJacx5yFY+EEfeEBSAdm0HRowAPNCNe4e3dByjSMW2aLsznpBq/bJSl
vyzcP+UfUggKUO/6dFXIGDFWyt3tYjHGh0KcNgvgQ4oRIj6MwpRakq4n+EFJ
3azbyfzPoGknH3OEYZNqWl6tKANZ9XP8gN2KLrQFVh3XewmuQ4B1orqJs4nK
2zBxIy5eaNS60xNGOtXNDXXBg844q1vqCeoSOeFzxFix4dtubk5zoKFMBT3e
7bXz+a0iPmbUA+cmBiFrL3bHJPTi/AYVld3o0l90AE5je1mZX4F34hyi6HkS
2++/6QRvgJeDWXEx5nADDB16dpki4GypZUsPdGFVt+vH/2HVxeb/IEmor4c/
E4ERpadx+3UvhIuYao7VeVLLwuwy1s8LmBywUyhCjoJySPXeGBLGb7HWBUDn
p1izKM5jl7GrY524ekNyHvWq9YYGNTCJCx1cQNnQscJXQJ34QxeZ9IGqHkuS
b6WhvqlLgBeiixMfr1SjKpO9UqFfIGQELtEG7YVA4FFTHFUKDCTcT11rUwo2
wP9bY2nIknFjMjoxPuaTi7k1HTQp0g0tfuQeaVbeGjRxL9Ke+2mSc28VFIp4
ptuUasvHphQIH4vSGuJCeHuJjzWCYkScIPeV3+eiM8JCcWNxav44ArDIYemO
KGkUqA0HWyohYFMtYbRadkUReX23Q9Ej18C9O2W9qY/P9IES9j5akjPT7aA7
27cjG77JZkLuDX8ocC/3ECSN2pRBWiDGAYxns1/HQigfo8srn2xRSuhgHw+c
B9RdNapUoWxJkixspBGYR8exUlPOP9dUY5HD69pOxUAma+gGVdCCF8TyRoeb
3PY8YQKX8efMdv71JABtmw70mZRPpKgCREC6uTcYbM90j8pWXr4HiRUIhnZB
uvERdL6AIKawDEvqeTDeVi8/7f8sOg6Ic30KSKn9B/Cps1lDpGXi4WkkxFri
FsE4u4uqBDl5CXD0LeEf34ljUXT1AeTkR9HaOt6nT/Ck2wLgKblu9blfHYYM
qOVQuoRVD5hsql/CUVvvebz7Qm9xXd+doPW72oYMLLLZp/rW0b4VhyrXq1bi
yNgPzQJMyI+3yPlH9S7yTQrVvCR3PRXzW4pb0I0dkxsk+ta8iTUJ0LgGzikT
nYm72CN97b8VDC0hbZ5QJiJB5nu+nvlhxpqbzj0MU2llu9CUC7wM3iEVMxHX
PNtPdcq5ah2I/x+Vv3rhf+Six7wMvfHgA28rKx28B9jZ4BPHs5JwWOttDAIa
V3CTZpuZaXoDywWKvmEyB1dqg7bGRhb/uD7GrudL5RB2O5MToR614TWxfYDc
Wkyuhrxve6gElEpTkvBeAxgoWaC7TcQW58IHwUt86Jc7KEGivP78ini0NE3v
3VS/yT0/hnOcaMQp+7DF+iHuvv6bZaad9hcGJQVQKsaSTFViTv/PAApwJ6km
l5mhRhkP1r5Pvby3vYA2cPzcuHJqTic3ALY2Nokf3t3Wm9wH7dgqHKx7uIh2
o2vfh48fkTXNni8dYsWyyorrICL0CNM42q7AlMpPwdXUG5/YhaLorN8d9Bp0
SWipdIoCg1Z3qrK7i2MuuWvYQdOT+lrjHVwACm/qhDqrpG5SkAVzQMrjTxch
KbhziQYHTEAiz7jGMoaW1XXzYeRVqzLrHFAndW7oMRTWdelqpTwfPzmQzBJO
Ea0CKYRyopD2aXQxirehiQ9WPCFnbsOYaPNdkEadY2LTgSSgmzt+lE18F50X
E5z4SWbSiL+6pBQxqpBzpKV6H9kVcay1KkQHBbIfTGlWFQw4PT1NC7qvyG4i
TJPxszJhD3f8CtfPL6G39ZDQ4jabuWaN/V6Xm4vpNpiYmVYcC4Hyv8ldNywT
wYWNiTS6MGXdZD0g8cFxGHOnyb0tlsjAGCJpBA9PbyUY2bJ7UhzWLknProN3
8246yqxnoBjaCUAhyEAPgL5YHj9dn3JJ96dG51MFHUfSJqVt0mI22jYEhJDY
5JkQGVQcmVagHt+M/rnYCPi0m5iA80/fOnIP3jikvNwW4yb11wPJMhaIYOfj
Zc3v5F8TSvN+wqKslHKnvShcXy/NaWXjKAwXSZUjSV51yrffruBh4ynYXIQ4
jucaYYZi0NcUJKXVKFohSLxQ5OrEcjctW6Iz4MCh0FCJjXOujAm00mynDbxk
fj6NvOK5g0DILcQWv6cREAvPW7p/SUn0aor1Jsy+KaMuMwcFNyrtlgTwDcAz
zANcsq5TBjcZQ7+q2O8zHwOyix3f+OdwLIKMthfwuINcy0GOUaNQVVZVuuO6
HVvK9kZCY8Bv3EbS9eiXRT+yOHMIioowTig6JCsFSMKWl0vzqJNWco3G4Xee
R10IWoBIUmcy8nl7aMSHQO4VEwBJUrR0UJeZWGQ6U3iBfoCzHuu7D1+CE6WS
zT2CZIZjuKiPmh2eWCUAxDyLXqmnr1yriPmItpd58bvm7Xp4K0ojkY6hboBs
wmX2Bg06LuOoP/TATd9JHYPmhCjK3x0JVT25VhYx8b4OeKLEF0Y57eMlfR03
LPfUvyKK8M8d2Dy1f76XyXoUDoIbpshi7YnC7nrOUm3PP7nkbD1r4bpwk2M/
Mur1fSjq0Jctidr+XfEP49aUh85DUgxN+vJY3CjJqaIyfzDEWaHDfHI1Vbzo
kQOT3M1p6ul0ZioyAUCRfBDCayMy6D/qtfcfOGIRl4RPe0Dm1nk0hWzuU9QB
qrYus9I68Mp1q4PlkWa5UBqXPy/KmkkQSxH2pyFP7tN3GCwA355be3wXme9j
GaCFD7Ojprsj3iqHjbkMaOV6V7LHHbEqtEAPavkNk5otcZeDSJgQ/kf2Yd53
FAZbZxLNDSERHK7IaCfYiaITvwGbWE6t1qfQQiZh6fJ9gK19i3r/78aOrTXi
33wrG00k8QaexNQ26KES4yL35QsiFJvoTBbR7bg8FNDsl1vTkhkxZK4zSQaz
ByHAd+lFoWQMS/jZLNShPCiqfv3lp+as9XP1YiiDiNqVxLRmY4YDioLSIrZj
CGv4xaganZ95yatu5P17xIxi8/mBDOE8ZvanMTtcX3xTFbbW5IBtrY5Z/ts2
ssbHSzmZ4X9gK65Ivoq+4RPYMN1t0V+PKBtVQpKPz1xdhs4k+TO7tou7cKw0
w5tBN7DIOiSLMpy+KwKsX6sDJiXAOfQmdVyrj2wKn3J6kUYfnYB6OobUeqE0
eAkHc3vuhYbt3VBpanCSxu4XXAbUXzyWCEX5N9IbZ5UIuwYSACKJOvSAkzd4
4eKNbcIsyyFQWn/CmW4nP4XXDg0ezgtUA3eV8C6Vy/860Z8X6l3xb4DBc2O3
k3MAGPOuiBBQm61TfFW7YT6qKfaOModE3JV+wFRxosR0tJpGFQQH0zMyYrWr
9jyyNuK5SI+wiY4SHDXtkyxeis1Bqn1RAaqv5q8dMReQBcMGD0y7Ae/T4LVk
g5YsJJ5pKU+Qz372CD3yBif9AY+amGikT+d6C3ZFX72GvqhALn7AiexO/nEB
2QM7dLoJaeCBn2WNECDI4SGO4Pt3nzZwVPS1TjIayH3or83K7JOBHbeFAqUt
FqARn5IHCBDCuTcMLQivQcjC5mWb7e7NIQJy8xfitfwEof0t8NGxQOUnecwt
FTLVZB4A07VC6bSValrnz0VSbmyfpxgRFL+6i891+n31Yo5ZznMswuRBuMEE
8/RTi07sSxFYwX7JocOq2NeoDDOhzr/8dXgKg6LjIn48Mua2cmddWU6oRBe8
heCH/0MPakog75Z3jmpMFYIVosIqUIBw43rMUtA2+SXpGDPVDw1foTebam+6
lNIUmi3tWYIfRD6bc5K+6AD0+H9qnSPit27R5VB+P+eT+Jgb8AltYJCvXzGY
eunZOweEIFZqgHnkAsWxDBm03ABrNhVtqjb4oXwLWNMnB3fQT/v8VezNs3fO
gy+rC/sfh9H7WteVT5mo7g3rb1/cF+w8uaMgd48UoFqkZs7kB2OJBX2AvXUY
0elmmos9jBiy2KUjgMfMfKJHJa8f0aFOFxiS/yW1pzna2/ZMtxImjh6JNGuC
k/k0Ov/jpYghGbD1aMtEYJOX67ZS95aHGbgEjaqo7NKRdzz5JhLo02Xa+lKF
G55MnSgV8rbyUuON8ELpQ7zo/DKk/1yluOCmHtBkEVbIHZQhjOA4FmIsmpQ5
oIJ0VM1CXptW+jbWiPvhSvcy4jrccxGPm93AdDA+LixHhodImk6+4YZyIgXM
gObbAscLPMDF7OV2G5U/j3Haqb1DUh79vJ2kh1UXoOc1w7JtqMGsrqu3xSq/
DcvI31QEs9RceHsJJAUsvYdN86Uoe12uvc9KimjxehxFY4V2U1FnNA6fhnRe
FgANFCKxUjZuJr/GdMnxjz0/rEIe6mxM5B9jx0mT/Xfa8Sk4lo32nbC1kDeB
+Y/SQImkctixgeO0NqJKDAsN5U8hc9JAx0CTpGkeun8pt5q2OW4G33eCyTgH
++4NF9Vvw1gxmgORA/fueJzltGkHqYSvQunmfTkuRCLQgwBBwBM+mGTqLW4O
AsQD11AKvz1DmVpoKWCEkgQrc00cTti8VvDz4YE6dEwyvDZdGrxOCqQxpyGW
43t90XVE3TCMZoAkf+Q0gP3WJkIpCsjXARJyiSUa2cL0p9d1+KRMUG4ZUWmf
bAhnDePUv6NL/ZrYdw3F3315cd4AukTzhK/h8DmgEiSLHp+lQcTklQfUmkjB
WIoW/mjmnqGh0zRMmE4n4KkrPRZRYajOoCEldgs9ykPT9r2e59eviY/cCr9i
7wZw6V0FtjQ/IbSeOvgWxkCUxEButyxbkXgT255pY1m7B2qspeRKYmZ7MASW
y3lQFq99vsr3Hb6cr6jh2PdUEZDnAGz2FI+PcL7XNNdB6BmBAKhoYBK2Yv7p
YOnbPukh4yAMFjLjRzvpw5QOtcsXAUsfomEKFtBokfI7Lc2s5N1LFd2cKJiZ
ATthj83AEpWRWAe2WQNhqSU+qhezM2J9oga364PwSAr8FIH7B7ytNTAlbYK9
TeuDcV/n5mVLVQW2YYFq9Rb/uA+kaaft6dfrZUF4O6ebHLF6b3JycXmFCMHD
/Qeses4q2qfkpSjC3tzZ3nRsUCfBa0OQmokLn/zeEFXXiz4UM7G4b77HhLMQ
JTjBgIQM3kqv5RmRgxFF7jgr0YZDUYTlfe7YQWhF663aMRMY6mfMIQGKQBfv
saR1hfvwNoxzc1r7EoW268We+vi2WUF0W7QmDZnxSCOe3qLHza92xdRx+sLQ
9DzTWtfv0wouYwOlxH1YjWEdDdiVMYN3EvRi5cf5wUipedS93B4+Vfc6S9Qh
tEKwb+5fWf6tnOow+Qcz4MXEZwn3cV9UH2mpEeGbPyJG/KUNykWAoCD3xBrp
6wraJ0xsqxbTCQs2C7jEC8T2Fnz9UlpGEHhilpLuB8pJz5gxLnI9MY0FVfNC
oJxngXTAaMRwMx3e3zgUNY9Aiai0FQHcpS3h4pRQ8HV8SXN7fJRXS6ggz57B
l0p5viuV+o6zYoYKG4tWUke6E9Jg5y8SszP+xJQS1C0k2K+CYnldOoZ+zoTk
Qyl6MxdeKbkshsnT7tsgZwPOq60yuJ/1pbn2DqT/rQx64Ij43NtZlD865p85
qtSz94LekwU6R2TNOdpn7f6vNTuUAlFTd2ufxRi6trYCwkOOe/TvjhaJmo2V
/FYSLxwJMMHRqkPN02gNTDGoNL0gFq//op0HHBo9XhAzVmttc4EcrcPiSRHk
7cYsV45G/SbpSyyzu84GM4Bmt3Ncx9AuUFwVdPCuWjwwqqVwz1JtzD3C+GeT
TyIMriwc9zAAKFaSPpZMQZr0b6ePOwkskh1p4Rpb5nxn3LCuK3nThbXdQsMe
lFs/i2lUEL7EAtyQle/5z2Hw8spQAmkQAVy2Sn8P8u00BStwoEgM5AT87naW
KIxA4jh30zasH/44nIT2BhqV4zZWbVyYbxX/+xGgoBdMayIktJAe599sxdro
8YSEygcXmVy786cChHhfnAmyIRr5gh4x6YApCtvUW2qXWHYYzwRAMXO3JEqO
O744IF9AYzleg1peSDPC4cLG6L18uH2x9XtwVgPO7vWKa1MxjxKXJ0jr2mmJ
kxrDVwYM/b1uGBgj+RXW7ITgFWVkpDhWu5HRBbq4cOcTPBOOc0gWmz5UaDjD
C+DUG2rqzx5h535fAg3Ucm2HHJ+ZsDITBWM2f0WInAfaFyfhA2IKuiOynKsS
DklIzluVFsxF/D9hkch7FHoxccAvPIEocZ+VFLBF9UAkcwHgDe+z6RHKTnS2
asgWQuWYoqtPHeNInE5ZuTg08XdH0ReaVls58nJyvrKLE8OYSPhvCCnF6m98
lS/r96iI5dpYeIo7rh9x32l/CgFGPT+JnxUbeiBgmDdFpFfNnM7Ef5DX1giP
3SGduFP/wYAPdHQXEJdiICrjvGGPf4mqcS9j+JRaYxyTtD+/VhTSx496r+Bt
wRQVNzYT6NElO7P5wpC0JGSxyJT0XneT4T1yhWcDsltrhfqKbl9kDVZjHVv5
q5v4d3YLt+JDz6liWhSlPCcSbOnDGS9MELN5qPrr2c6/Rov7kM8nSQ7hxfpk
XPkWhIzav3w9BfXqphBKf64LGrfNIKyM7WPjQNeC+AFQgrs3XEo6vvhLJZPE
WnXn1QkMsDa1a3DJdIg2zdWfNlFlF+ZIPEIMN/8ugDP78+PBTyizGwYsxQKP
ft95AL/ww4/clcZ3kTK54bnmhOrMnNWUGcr1avdBUJRR6lj8xmLVlzg5Goyk
ccwaaydndcSTvDzbT2/EeM+rrTabkfyWPnFMcAmp/xRuAJR83xPQjzA6ss4E
HeLdzZ9oPjH4frJfxPwQmJDC3DEIfUS892ganWPag+IPU0fb8yKh66zUtMsQ
Wy2qi6utprUbUbo25VLeYVfWsQDG5O7IceSQHV3OgZZVRMIHtZS/09EYkhHe
uEIi4B2b5yU2jS/t/2/MMmkAQFCbXCFPZ+evPKwaAwpUjyG1V/jkpQT6PpA5
J1rE43zhhglFllC3HH7GGu5GRvOBaa/Lqu6OZB0mBxwgvtg5Or9WHr168Pvp
doDJuCUVAFY0C5pg52j9mvv2SfOzmqocKP54Oy7dVOBHCpm5ixVWBQ0evkFD
ZMuTCTlLzBHzCKsrM5VQSRwjYlxdVrI6s9HfMJI+IpYPQ4udbARYagWsbqwR
nvY5Ss3zDTktkuUw+XxUkNW0PCgOiZ4InnUcNemUw1FMLrYRzB2++V7Kp/73
azsA1i3JVmR7Cy4LsqafRLy1uN3u5BANagbO2BQfhpi0Pe0NiBF7aHujsngD
E9JQjniTPY4OPgGNK/BjKyjeikNAkY80m1m3++I3npgWtCYzdO6LtLbSJMsq
Whw5VyX5ZP3/H+X58UuILC1k4T9ukgPci7albhQcwgh54t4guN6HTEyt9as5
4eBFGZgUEQ+6i0o6zKuZ55PZyD4jCpGQ9M/fpKVyqUosgpqFDhdQfqBbbqlW
qxBvzJGzgjXQnBmXokE4ATBOq64qiAvc3YlCx3da6GwiGHOB79WMTTikFEh6
A77nTZyn0YRzLcjBR+xnbClBKQf1gvXmIOYwRhtSNYiGIKmK605Z+Vg+8tOJ
l3ChI4B6avi6LO9LDQydJfmg4DmRjzBFOVsRyMvyMa69GyYyuq+lMxqQfZpq
pbOGUrMPfnkhUGWwHSme+dIMWqnNvexwfT3fMLDjlGYNhNmTxeGKoGIVpy3r
7NkZE4QISA/ez4q1R7Yj0DpVpR4S9jjIgAynwnSI2P+CUrW8Lh6qZuTEqST8
0yG3mO3OZBc/v8BJ/cJc3mEG10lBTQHm2jItSj1JxvRz+BgeqlvoNsJADgrf
kckjdUqR9QZvruhCBkwUMdaCmzCFA2tXRy5nZgs6mYfQwX3i2QYJ59lS0AI3
pJapndUSiZKAkpe1Rnvb/UesgtuuD63mSvvOg9OZL4rJc+3uSx3c/RMSZJJI
JcWeyGkjyPSg5ALAIdiT7Gp/XJNaZnfe7oCgbOtsUa7l2b5okwm+dttIPk+L
/s8D/OjCNkqOhCc6iRHZ567fo6YoYLdovVjiXEyMBcHqDsjnVHpRDd8KbJET
dpGvHtIHbAwH95o2hzxRagzsZmhbtDS3fYP9ZOtUdcYxhLtG+WaUzpQZI/g4
F1s0GVkpbPHIuac3H9LrtIUT1UrIIoP+IQirL5CcUIv/HPIY4Be+8exDQ+bz
WiZUsiNJ4Uj7SoJEJFYEZ5uKoYLH8kAvRNFdoPpCds68gVB1NAia+vSrTtM1
kXoL4pDr3cLLoJYL9KcHM1HLVF9DsQ+lbSWdsopkF1FPyxvE/Uw9MajehJ71
1u+W11MSX4c3Ij+Qaqk6az+L4ZyJDl/Hxdz4laVbz3N8EJZdPLpcP2xpcwdY
tCxXJxlbAGlYtzoIJcs+HFIjXPIgsuXuYJEzzSC0ul/WlqFzkIYcJsE9REld
xamHa0fbCR0qGmEGzsKJmZl+hiDNukp/V2SEA9MYtAY7CN86aMkHwLipWvUq
A0UB1KdbnyJZ7PfJZGMS+J12JaRdU0RXdOAyS79p8rxIVanPTB9jfnpe3DXs
P8GYkno4CvBGFy/ES/Si13V/so/ErXNwB1Wbzx5+6rcwFsoTU880EDoZoAPY
1DHa4V9j/cWPdAMs9RQTvCa8HYVpbZISzMMwRzrV+zPpiGkZlbuV6+mK3zpA
9STPC+BPSouQP2+TVbjt4OkeBYK0tAWsSaqGo9esC+L5S/Y77GZiQiZy5IWB
gDZHWK/7kQyj9tnerzIKYYmtIA8yzaODCEhiEyNhkdzW9IAyHMV3JTucaqiz
S/s2EfhJEYx/1A0bOijvX7CDkjo8oVIE19MUp1p9hcgA8qss/niNQbwLj7HP
EMLB3pOu6D3JAlMZz2knE49dxYkNYuqS9da5RCKE2xxGgpfn4w3+1WzCB3ZS
Qm5JEOqZkB2WqfL6vxJMs5M35lFoSNqTRuh6Y2AxSo/jVfp4WnmiKJO2FQkO
9upsHB0Tbe6wYqzK8AgEE6Eh7YwE108plDtSkai9FPFyK2YmWCWPJmkMREth
3YP+FSmTHZ48hmMHk9Qp+Pxors4RMOUWzzTFHBv5kafqDukaEXMjq+TBVsfm
8cRjEgND/BIGDNO0ZCKh2vup/2bkduyFxIkNWNRxUgOVeX99axfjw9xxnxtf
z/eBqFRbiVYTfqyhiNYCvCll1RHQ6E58114ybWZMTQMFc84Zbb22eNVMj91m
yb9J2sxv4uBuss6rxkjPkc3ZR08jhECGj2yMpc+v4Y4p6jSzXP+yL3l+R7W6
y+1h614NAt++RehRXatQdAg+MzYcRVfuXpIY8cuStEz+H4/El/Fx2ewBLATF
6sRiUjMIdHESLP6hMfZvK7gvNMJmWS1gUuy+4wI+WASJMVy5jl61ql6uaoRk
ZQGfjsreATxC1fsSIaSmjGEm0CLICqrHKEUUYdMNvCT9uVlr21muE92v1nAL
Ky3ucVt6IOCK/qw/gHpDhsD6BKnsYbCdsg6T3QlRZgrRJSHEP8PFy2hLc4Ja
7lvNQIEn8zQR7TF80YQm0/nGLpitBJ71bzU0cWOgpPUDb2wAMFu9bJp47xBL
CxLtZ40NshcMR8aPvbcj+e/IfSOS8xSiEix0QtPAII5bLp3J+rKBmZJlzwnu
QHMyL/7NHJz5iok5kZvv8f8FwT5mPPefm6OfqjaO/Ij131x/GSMnfpW14Q6O
gsW4ENyNv6vvc0k/ADshybZ3Yy+yIozToMcM3s8S1OwEEdfQ3gn3KreYoJ5t
IWB6SO8V9TcnlUaQxDHu8lsVm6cVxmeUPjiehsZD1zM1zSCRObtJNK1BFeKF
N7qpIKytSk4MG1ZdpMYpGYkyuej12MsDoRhUDqU8THvCAXJJH11HXVi1XC0h
WwyM41O6R4BKFAAThgQZ1LV+NL7upIGiXtfH5Rpi8mcX1hdSd8QnKw/iHJUS
yp8+EDevDEsChAfee2ji2fMDFQr+VhK2pVVe82G0V9IxM/e/4k/UFhYwVNq8
9KoqRj93qfMBAq0xTHcptwC7S02btz2ewrsj4LQmG8b6DIHwxjaRoH4q6LFv
+OUWzb35CMcgLjj/pAEKPgPn1+cLOSfjAkeK4bhyrttotg3g6YDADxamP5vI
djm11wtR32ZFcjrHCsfU7xUTeJvOWVaVVWIaiVYOKyaRXpA5m868P8vDc8GJ
k8p0g3+iBOzHXVN2x1tvZS3j0D7uxjqf0yfj7pY5Gun1uVe7NOny/55o6xf8
byIg1Hb9D+CroEJAnhpJkiiLUEbyWH6j37taWqJZjxltzNmEBDPHl1SeQ89Z
tpKwCcSwA95Fhg3vIZaur4Z3JgKxMRyqhQYGVaNxXliiyM4B7vk0krByRR8R
lNL64dED9yAlwODbzWN5EIE9resEYX0dfYB0IMwDX5Amfqj3g3PNfZmzBbjo
yrETgqwS1jh4ARGD81vZ+Qy9NLSwZ4UOa3+UUvozHUQ+KTBoH4bXztd6wopm
zpeVrWClP3SWjTbNu5wIKFl1VXN9C8Q5JnGuh07iIORlOn/pjHR8h3/Fc1Y9
2LSQ1KxRF/vtZ/we3QlD4rjWK6CfIHvnKN6qiViW3PFjXIiu5rfNAcoqGeTl
kfDSeWvRZswBmATFBjbNwKsfL1y5XdNsP4zjR7jhEDf3Io0/RXu5ORwBIg2E
S0S1B7IIiCDL1ro1o96+FmVbagUM7H0a2x1Wrz1KxDbQzTD6rBIWp30Qh2mK
io2yGvQPcc14jtJZdIc3HFAD4/v/wAjPTYoGekfBIrUkPjoD0V4ReoTo6rPU
x2X7sd0nOLUtGLRjpLsfmXUbGn8213NUQmW7mg53ddFxpOI5TEr1+wYsl8pM
EYSNsnF7D/IIf3e+ChmpqrtNsXLxL4ofGwqFs4MQ8K3FTE3D8VxO8nUYRyOX
F5ZmZmlQ9rc1mvOZpYfUDc7PTLi2IxvvW4YY2BGne2Kiwxb1Bhp7zQwg5xhv
rGzx4YTVn0u5XoF7H46K4HRjZPuCvPvOr1YSfFpEl15Y3nSTzNaKHK3ui/2V
0ev6n3RM8gWUimG75S2tGYYRn6w7U6rRCXW/nHwXX1Q3GNmv7R4DcHLslKab
1Zx3sHdyRLaaM0GMgHiIK2zO75lL0Kckctv/aDEh0wPJnqPv1NLOCYFS3NIl
GbljTmkS1EAM2Lm54da3FWlJ9ZzhAGky/T29ckiUL7hZsbe9zyxn0Pl40f7O
6hfHhAYRh2o6GajWmxPELdUwPU8nCAHYkOoRV3tlk0lp4hfUrqSsmaqVd7ee
Ou3Rjapd44FPPWgV3yqHEaGXjjOZiJSJvgYhKyQ4QzAaXwZI1/oJt3MfLLKt
H14brMnQ+A1sGfFSriCvgDPo0bVYiM28qlghQFGrsgSYW4zDB2RCWamPKr92
+vwAAyfmkFN9N9NvNqtm7cIVn3nfArYm4yQQeH5ZwP5Dwltjyt11A+Wnrzzy
IP7nW4j8Ax+cOV8cfj8pbSz9kuVSxgG9x1F5fvwdlz9kIE6DK6276i4XY1cj
ujTmSNNzwn7amPpw5lmlmow7hirKx85OGOy0jyOnvKMF8TJmNhMmPn09s/IZ
tLAuUQXzszZAFiygKyzLJHejVaJMUV33kFx7OkkOVCg037c9LTSauTLk4dMl
r9VtkVXmIm4he7sapynSTuxVxGF/IUjJrmTDW3cPGm4nHjUu2c7JdKTKXcDl
zfxeDG6ywQHFjTVXPd/nHLxQ93OBo4kfQyFHe3ZMRdFgVEbpopGR3n8k41L2
250qacywNGjH6YbFrzI2RBFx9hD4Zdvhpx+2ZYqAmfeZA8u+0RT4ye5PcmE6
GlWpcVDo6LT0GZWF6KVerxdn9fTL41hrVbVHVk3SkBfkLiFVwAJUUdqb/5ma
50GJJgsZN0I5PHdylnjIYMdPd6G6iD56Gw+EIzkkqznS7xh1vRxEy6z/QGoY
fwLXumhq6ZR6Oex52jTXhnszX9vn+ef154NijfEalOdrPHvUbnqdueMCF2QD
nNgYCCFBs99Hgn7wI1RQTKTtqQTBewkflpj+NLAvTI8+V2e84FIqfcqOOrqF
fSFIQ5lxtpzCHOW+MAtDsmM8Sb0wZgAHRVPareV0DxhZHXlzrZCDglebFsMN
QUNUKSHuS9sC0VwFsB1DjSSdK9jVIiGKCYkJaAfi8O07wkyObe+cNSlV7AkN
XuSJvRAYObu3uddKH6odllmzPeAtJi/miP4Lmbp/ZtHWzArlzWiVuIOBnqfX
1983GfWfvWKEJp0nqY1VfcqURz0g9BcgOhv9rPF4oeSAOmbC/dLJije2kBoH
iHYZtaV7rztb3lII4PQyN9clCR6xVA4SKkt6z+zdjzW/rQr1TU85cBy1udB9
aq/3UKndJP481Zt5olsKnmS29Pl80yRjeWIB3qnFjHOOcLdhE3Syhdc6aFzt
0Ri9iMvaYLfWFn6+vi1gw4U8XBW0ykcNM3u6UD4zwe8V6b4rTtnwFO8yo1gw
oUro7qCzUUUwrKqQpchV+Go9CGqOcbYhC2Zf2OYylIlgZ0UI31mMSHoiMCKC
4/tGlnqWuSXY7TgsS+cPIPTCVEXFrT+o1XholK/QWezrT6H4zEehbaOQzcC5
wGRRjfAbuoo6OqHbqwMOzL/G0y8YC+xSkpZ439ACexSUWqrSI+ojHMvlcAv6
mGZBl/maXhU/v0EwIyM+y9hqufEcYp5MBCjOpgarY450JQRYFhcwWp63b6nq
Tz+p4PdYtWpFYtmckirlbZFLfOVuWK5SjbhEIU46ZT7urHnrKG/L8Vu33IQI
qT0amEt/RHq0POpS6b1k/jz4/a6LZr6KdfZ7jOYtiQag7ccCHNN3UViEVsMF
WKonYZfUizZRqsliN36Rr6VO1shp/g0pcaKiG7O8UrAqXjdIgku3D+WMtUTG
qaiEd+xXMaKP40utpQ5lsWU2wBggk4d4AX2VE4IhDYJs7kVkgm0f8QNZFXBJ
hoAenjIRWYR87mlOaWWTuDjzXuaQMCFGsqz4tWTrZlJvf63CHmeXnJdCW/Ff
QiiELFlY2xuUs5AURI64T+vTkQ51Pvn7rjxxtWkdJEidoLW3O3VhQRsK+VLP
8Hirgilj0nmbTMw3IEsVUR88xsHKiEj7Hf+b312LAz4juh/rz3wV8Jer9WIc
CsGs/oACrE2oegLY5kJqdx/5n8ievxacgVBvd1LHMucuNy62z0kDt1sDpzmS
LusoiyBhnfkvqkN6j/d8SLLnaImn1+WPYgv39a7mKngurc8SEstptcBhcxrt
2bzSF6Pco0UxXxO75cPSL+saLDppIOj+XhExXD5u/Bjz4TDoWy+7d7c5wtnK
9t4TTjDSOFDDyJvBq51RByYdBoViGh4bzX7TI0OhbL332MjtIp+Rd9Tz2vs0
5kuSAk0PrgAoWQnWvp7lbcpui9X8AfT5+FNs5x9ZQb87TZ/OlexMZG3ZENI6
3nyEilnIjILcfVw0qscmr+o7ZIhg9Ntjalb80ApzXtB8qRSt0PAyD++9iYAC
1WLBxB7ScHIGMbOh3wUIV/70ifYDbwPm4uSXtyMNCLUL/ZPtCRurRZHVVcSD
gX0WJfIDpQY6cIEGajASJp937GfzJWlF8d+oDf/sA5T9oRP5hZvadnF51O4L
V7RweqJ3588LA4b8sBFAKKIPJWpJjnIlSP1Kh9Gn4mlSIKO6PZnhYvURWAh/
294uzjSs+Sv/x3h/xZkuq9iWjODmLDsVC5JV5muHqrg3XNlmVgEJt5yQtOyL
pniJ+MwwmqfOe1FFtzojkP9Q/X18n5RI3gENGvtJBMtBgEm4SZm6WmG3m+Q3
iCfeJxAFLQfrIr0wo9gVN1/oWpGELQq3dAVh38wEYS8+NBXvbWITk7kdIG1i
268r3/XgO6RLigprIjLeO0e4+GGBbaN8ibeHe80JGpPj9DTlR7KRoPR1zh6e
YS1w5yi8m7o0+uSH11r/BECATMlfcTEtq7XeR5rXR8GISWt7qcbZfZaP7dY6
YN9x9GnJIIkPKqXF8HsaLpbWi6hZBBVIp11Rg/rpsMKbjsqPAF5+5wMBdCd4
SG916bjhK2KS8s4q3se/Dyn5VWJAHFgqQxxo+hb38iitZ8vHFsqpdXiCULE+
T4marlu3zNs3ay4NELvJqrqxF35LWGuSjy4JfYOPaPl1KHGCHTXwUm4sAPej
bX5JRXjYNd1I4g5j+rQH649owUruTyumRABK7bDyXrVqCj/7QmLncJbitN45
MeFmebKlnrBF1JhxqrgmQ1smg33ypn08ZgsfYdx8r19oNgIw3qJ6daaSVvG5
o+qiB1s5nsf1gkhA5iuc8BQwxg72eoPipETW8gKhz+rYICKlKp5UJU0oVrCi
uglcI3qGzbF43Z1pG+Wrmb3YtADT2uD8j0C1fttRUPKdFwE/ZnfhJQzJCLuG
lD0ZNSxSypNZwSMqVwfEGkQngWO7PHb0Gtpu09EYjBYDQpdBzPsnn+9AXxbf
kSwdHW6S0DtdySmifDgRJ37tM71Yz7J7RZcTmFqctcaCf6HC3t1UdvOgG9ni
lSCNCeppH4zhf6HN/uIYRFCqH2b5j+oUpb9p56/HFV2WV63naZ0+J1YMrvd9
OoAlPs1jOwn1d6EPeCniRtRMylEqDgXdF3N62lW78MnBlocprS5GZ+OGHDFM
k6aq18lk92hTUM+mDs/Qt4lxgDXHvulBRvJWSrSyE9ZIOgviFm0nZwpyYQOm
QAw7zFztCitFA37ppf59TUWA6e1Ya6TLDYJw1sVMSmJMKwK3TfkB/WkL6efD
9Tikb5u1ExeOC/lJEchrufvaWKGZgBnZnS/634K3b5d7mfZASPefpoz2Hns4
h5Uhc5zxn/kRksLcakowbj5NYrCZWsp8JhWPhWVzzyp0tHNcrwnEx/GZAxbo
4v1j8EpcD6p4lW/3aacV8YEtZgK3DUv1JVmCg8+PXfRBTiqqYJMeTInvedly
9PIRYAH2Bx76imEOwHt9IRtxI1tGVu9S1TLvSblvcuhRwWiZtEz2EriXu07Q
zGmV+6yQ68+ZhSBLrHHRmkQBH5E3d+URi6nwcbT8v26NTpZw5JTa7sHdthe8
RyT2ZIVb99G54HR9WJyoHRbUJ1Bo4/SUe32TBpgxMgGxllVGX2QpkR8UUT7a
25pj4Z/5sX/2ZC+cIf3qGGazVwpscmneDYtcWQaXykWuLoUZ2LtpnnJJT7ir
kocMYrF4QekR7cvVAN1HBUBf+Y5/X6oVvODYo6J3dHDdDerXPk4Y+RFh3lPw
5Yas1gGa1ShqWnTE1M8MwyLzuz5TXPva8GetfJ9M/D/Jt1ZYehr0WRvXpKKb
Yhj9y9pA5f+aGwHE/wXB3E0b2vUgZ9FKuVwq6NMaDjvqbnFvqNgjrL6UY2xa
mneOCHvdZkTPK7LKun5iDzD5cRo6eAlGQ4+SmgWbFwYuvQHjPC35Hi8keaBT
YXLrrRFdrfgknYaKURvqrwysQZVdzHNGcCk0LoCrTALsa/KwTaqBNfoHohTP
jw0itFhq8+zXaOEffmW31WIx3GegXPAnCq0Pe72W4sqa/cPjN5c8K7yRmxCL
/J/Hy9mekZrl+hPY8SUWpRRfsCCDg9oTRx+Y/srHVG8NCGDnAdgLfNLKT9tY
nZFumVtcoRpHludH1aKjc/tFPKdlCnlstoKtFkTx9dc1MPoAL+4f0n2yQReD
zw4uu+/IyXX1CF4mTykpr+mw119j6KGHRjHB9szqmrc0JLmI9LXzd7YWctZP
ZALxRffDz6m6GGD52UFYBNxJ4BA2qfUEC+1iAHiInXdamtQchZNaZxy3ecZr
nY5EPeH953XdtQFAsLvS1C4W8EC+dfZFDXVsJaMqqZ94OHyx73H5ihtPmYRx
Hn5IYn78pWLA8+V4ZL2w+vYUorWk0gA3TVa0KRHIq/E4/FSkgO7gb2eyR1PF
KyiZrhjEbu3mJw2fscIW0JiRaXjXTPHzTzvit1d8iOPbwZsSL/Ylnk88BvE4
XvPRC+d3VNjiwvvyl3sdu2aavf3JnhRkxUcsOHzwDYOLz6RMGnzMsQ8mufsu
wsSr5XIEVkR0RubB+Va4QIojmRRQ47EniKKnaFSP02alHsMrHMxILpe7U6AN
Gh6kjARxq6Pc0jtShzXSzvZud9jeSuC58ylEEMM5l83d+lOClwY++Q8DYmY7
O5rrYcqr34mDH+JKnxqGryaZfl+GKVumocopx832BK8/xYHOCvDin1BfIiZl
PUo92hUnbKTBe8SBuBA3Q22foROpDXlNwV7TKRry52FqE3Nx7FBFM4Qr053W
ee3pYAD0TRWEr0ILvzsp1fNjCZmafejE6oD5VXbDkfd6DOvBUFDp3cmF6MI7
4UjFJ1LKph/ZagRdbyQ8oLrHBAxBiyHuotqW3EzYczmDXDG5p94nRqPkJ7jX
aYACfCZLg75OJMoOH6AAtAu7iomJcG1oBv/eGyojhkGhf0BRMg5nwvoJgoun
pnmbzA9xVfQFwMK8SFviFWflQx369zX/8t8rA5cXrWC/L4xVrJls6Rn2Wgb/
HFhK51M1f6WQjiNv5dHlQvl9CUfzi8km3smsa697NVOTwfe3UqHL14mUlKUG
puYif8PEt/TkuJ5bDs1ziwCnvIKn9eCUD1vBek45w+LBXy7F281BkXz2jHjE
TbmrSRxtLUqJN6jIrzIOUazYHfuSDE4aHbFBBeEwNWYpsW4+keH0yCB+tylW
zWNKnpHUIEnlyD/UdkBOA6BHHaE3iSHvutCHpqmbwC/iQGIoC0+zRTtuLLPZ
q3u+wsWDtn+VYuEbZCxBFlExag9XhBZyl6qHT27DzgRs60RyHQszJquX0TQi
US2ZcKNSWbkmdlkUIo5h1jst3DbsJuSKBnCx4GabtGG2OzSUy5GPZ1v77j9H
URmg/clYnAiTJ3xO/2P2n2JfBPpuMy3H+bw9j+w9BVBIB15nPyoWT3fVXD/k
tUzjPt+qzvgCISNWdgU0E+I2EuU0inmr78QF3aTA48bS+KS4mj4+l+HqpJxc
fyn5nPy7KB8RC/ZtTFK0QMLiRfBAQOJojpTNkk+tOHSxtPUTnbwB60+hbdUu
crAf+1WJRr/LzlZHyvEggs7SMDbvp1EFFLdi8YYlYABaIfU4phe742EXXgs6
Tm+w0GxDDW21ok6vSIDIYdQsu2ToKkO/323NEchWOL8dOZZ8XzG0bFelr4qo
T+xHKqZzIZWi0W5k6+hF6lEiAiABADgRQfZmQgkmkOGRF07aneTJLFY4+NSh
igF0+i2iUyAQrxk5VGR/QiVTPJ4yCM6sueKDYZDbnCIuSVnzJvMy6K0FzOxY
db55GQXp4LdgRruMVO7XNvZlLXH0BC1aB2Ckb1OrmGGr8EPNO+90Ne5eq6fN
92Bf7Elpe7utZFzF3qSi2GoqRq5AUN54FYjcArIHCKOH9qQvgQJpI0KeMNMF
Qtfvura7L45hJdfShONkIZF8mEc1mIpP60twTRrUfYykC6R3W26H5eDH7wu/
/qPDifUI2MV/XloTwPaRZLRwzWAMehwpauyRgZboLnjgE5ap8fWROd5yOeKs
KKXG2TYSA/ZdtL5hv7RHxDO97b/w3Rwxc+C/u/KIJAl8BFMltFZRKLE6UL+Z
p8r1WvRB4tZWIRn9AINgyop+O5vpCV6yG4vrOF6KtDremlXD7WMOASJbjQdq
+dGc04BNHOPruxvStHJdAKR+MhrETv1sptwr+O7EPAN7yLan1FVGn7pziRUw
nGb9+yQeNe3rc7G8gpwmhbc5b2lMId7i1fuXCzcnyUmXyS85krJG+/w4vGJU
N8kJgJsrJUpsErChiutsOd2Rf1Mr0bpGt/7kY7NVAvEz5Sr6iOvlTl8AzeRz
7ImVrC5IFZxq3c4zigRu1GuoVjfp3wZErGX3a07P9kLzif3RBqSVQYXsKtQM
VOv7SoWwAgGuTT287Yg2QZkke6OBvFZbsNLrxQTckHGOQnogezQyHgtcdKri
T++HJS79XX/2kRyU79QU+m4UG3C7FNUxrZbHzvUd3wkHG6BEvqw7h+gnPpUg
5qofmnDcJ2QKtHEVLcBrYNUe9Edxl3HcpNVRdYuPoXTZuPCK8Ilb5LJu+Az4
uLQB632T7ht3JJOf2Rusj6zFVpFdfvSNzPTcJqRDRPbOVCk6l/tDorCK6mBE
D/nt5b0yibyWYlUcyjZ3QucyrWhebO4Rsv8FlxZw2UXym3QhLpSP2v7lEv0M
Jp/O+t1h9b6Z3z1V2CLWlzFZAT2kpYJcUUNEDtGssik/nVlIeQ5pYD/oGUlf
yt9hmxc4Ky8TPhRBy03YlJ15WcTYHzgfuRza3wFV+7TKXxIBGG7fYEf/wBDa
+RRsEA/G9/3+DHR/WMSpWBNyc9eAH9GRVhRUJ2EPhcWAmKnKlpXOLBOux97h
L04hgDSwPU9vCYAtDT2aOQWE2LLqO5lMKpxHbvdtSZHMEuqzLRHaTcnhnfe4
FRvKWQpRn0N5TRYlhH4GvFkfz3McCF3vWu5lNK3chx8aqWot/dfp9gS2rS1t
gdrz+x6Bkf93CAHmaFp7CShrwqCgGiZ59lwAANaGx1PxFFqekhe2UV+wIV7n
l0W9thvgWz8yb/7O/FumoGi7L51TUCyEk7zwkzzcV+2pMv9BLv0jCQ9Z/76z
QC1o2se/lrgNMmzPa9Pi4Bcymoipa8SxBbrdwGxe+QGiBrgQ1Iqpeje8K7sn
iwGJzZ1nsVOs4juhwB+YVBPj4jAhQccs4iJ/heEpnLlHuQNlCDoBMibaRKZA
8hYRy+d2Ix7Xn3IyOIeYbEBGQcglqH2Heg/Qs0abFNSjZyrh0XyAdh4IrWOg
oT6vvEHp+5BRPrwuF31L+tH0RMHtmFmPOX5KwluZkkj9t9uoSDUkE2cnu1MM
Jf7+uXrVj1p2V4dYCA2VLUAgpy8vmbSQgjXoeNkZBWprS2KOQc2/hvzZB4NM
LlnYJFUw7LPPgAw4zuramqUbzht23Bu4mhZStGA+v9S1DqCKKsPoPqWi6Wi/
X9uoCzbUAuy3yzcwtxm9YvddtfxJTHwb7TsU8IIXCN3gQFGwTCiZ0zpw80LT
ioc8So9B9Oc4Li1kuNof08sNGnIMciguif6DlDfwVHEgy8tX8pY9WqEQS+Jx
WThHs2Ah+QkHcY1s3Mm+4OlXK6MIKYTVRZTQMw1KwfDzA7Yh7OzOMUH7TE75
8Ao8Zj7WNd6wpOi/XN73aG38ajP4DZA1qAs8KYQEdqV2U/1XOJ8bGew2e/2T
k3C4MXTs4hGivn6Bcj6EYsEvLSk1ewySnOoqM7PXeKws2t4cuvYHu0JxHKfZ
hUw9rTcWgPEkE2ethyPYRmO0S+hlNov0OhiZ+MiLCIVCEby/PAcVhNY0PXhR
LXp6JGmQ/YP4KhvuywiFmiia6Yzm/0gLbyqGPBhjpuqjYNONSF3o0sRYAcLE
KDcT1/6qF5F5ly1mYc+gXgNceCbwmlsgM2pFEPkX27SEYZotUBB6RxvcdJtC
LKFwnZMuegQzMS8yUqYot/BUxFDlpL9Rn+LQsr6+eOYlgzEG8BTXgimdaysi
4y6otOKGlVfeGyBId1BgYf8kJUEiH+4GzVUD5OrFRL6FfftPrzFZEwewYZGs
aQwp5TxzszZRJPnEseDe4xovF8f4Mlv2R1PPbIpoT2Gy7gMaguwVQlEKdfNZ
UN9tnflTfeDCJz4qJrMky+oPg4LGYqHqZDoEWpybOeNAJ+O50iTabk9eeixx
CNHJXVDZDqG3tAiKLHCXtvHmwcxanJSE2sBZfU32aqNwXm/LwL/f59ByqK7R
3yudWWooqoW9QDv96OJ46IdGp84TqDN6NkOdtZ5Dnjg8GT689Z9KVC2aC75a
8jfBeS1bre9g9TgZjyYd0cA33Ijr/plf896ncosOCK3oyUrGwNyFl23VFRXe
dWqAqbacTovASXJR6XrPnQ8GeyM8NHlzrNk/L58Csb3xEN+C2xshEm3WIeBP
/2IX4Ev+kddJwzLWuiqb23jZDVL/lm/syWUKmu76eRBxziYczgUVBwEh8tON
aPPmAXTNp4WE+KGYfYH+Xuue6y22Xdyj9pg9j7k1AQiT8+6OxGeCkDSMN8EA
ItbyFmoJKdb5o6Twj1ckUW8/o3UA+urefbH5F7HpSTZdCV3Og6E3k6tvm7PD
oFEzyi5YukXoigdB7NjwtWLgyguGz5soHP7oHviYvHyinhXKU4+SCB3MFnJ5
SZFgkK8kP+12NnXTvUJkNNCfPCiMQFWHRUPkQdsGklA6CEbwmP3AIA/KS7kL
TQGyYQQJhCGm88lQBwklKqQjRogHFgxgYfyoGpA2oUac66ZO31f8UAHoGyqz
OxYACj9Uy86qUgeYZBPZj9lqYh/zPwPtRaujewXokz4ycH0p4oK/yOoV7CIP
7RwEQ072GDwmON48coqxIdgaAGO00tGPSGL7VHYO97e9S8m43bVbnJOvVQIC
QBFlwL6NJtugBF8ktnv+HmFd3kbrkT7yjW1+roEW9dC+/VKtwC9j0lFOpBMa
iW02XMjKyXGGuwE7nphAsOslIFNxOY4KESRzGnRhwTzbxhhsYRCyvp3g1YET
Gb4qDISpmvgbLXkce/FZHwn0id7k2oaE+CJcC+RacdHdjsDVbR6GWwmUwi6Y
pVa3RuddWZndqZ4yxh/SaUnQOxnTNnHFgy/u4vXmvNAWfP2ysEtmSYAed/Al
WOHTg4fL7+qE6ANmiqSW1OLctnWskrTXrDQ78jvewzd6a5gpWhEx46/nv0jb
rfEetBn5YovmPGKvk5Yk2L16GceTcYCv5J7ps4za+v6isTNq/mSSwY+LLoTG
e/RBqVQT1HmEoVnIpH764VOkQ4aIHi/oa1RRCratl/nrOJG/OhLrvMU2fgs3
oApk5OpMcguH6QwTL2j5OjPAPUNA1a5HZBfOsijJOY2hErfvDFMFZQSGFyZs
H4332OnJCfng/whZyxst1wiFzidfBOh6j0ktDVFz1958IW84fi0Ez7K74LQL
HpY3Kur+B9GOmk5pBnRXcH+rUwGKe/NCbHiscsvkCJJ1ruSs9jW2virB3Ynx
MKP9Hd3yIne4kQBUQg4bFYKpZEdr7vZYhB0He1xsXLBpIVNA9sQ9uV0aKn7I
QAFTbK/lbRoWz3NgLdDXsQw6c1eZbphheLZW67UUXIt0gR0Vjdzrt30iCaaJ
tCpYbi2cWhdnV7ntNitZCTDXxFapm8zBsatu9fZqlNBwMiGBM6XHyfb7x4gF
FAMaN+O7RJgHJgvdv9PkwBhWN9Bvx/blg3Ri2QTl5jCbEqBNwGsrUoUl+9DU
I2t6ZdSlbE6H+lol5NNlC4D4fA66YpUcMSFbjc/5SZGtZNcecVtOxRlArNPB
6zQ+J+C8MPMfz8GdOutUY4wbHyIwPcvbwkvijphcs7ufNGOnyyv2hTxhLo35
LBw4QrTGFfaZvXFFPfbXaFCrfPNfP8OA+SNJ6wb2Sy8hCQck67zTjcTI4TeD
iX9nLKnOBeA0O/knFevOyiWB3pKEZwSAEmdoZ9Pk3UdclQ6CvZCRSii2sYKa
RBm1l/EO5mBYpM3Z4D+4RxYT83kcISstKFQ/+fQWG6jMht1bHUDcv4lqwfw5
Sq1NRaN3zsGYwRO9m2M284fsHTW87KiJbLbVyl8h5BUrOhhQ3OlHSSMomzRr
i0Y+vZTbyVF2iwRnk5Y9G0R9cWW990N/4UHt8htaVI7YGZjGJ3NqQ3T1c0iA
NsPN/vx1V/Wu5zJ1+Z/ZtYv5Hni4Cxj96azH5NxAZWqQBGEdsbkNRRb9IOzn
piDcpnZ1pnfhTSeN1na6dZkQMvlWx2hNoXTiyeib1aie3uXgt+LsdfhUu8fm
NvelCTTCZoiGS61I6KBhtWcnJ62kyMxVhT7wfu5BlTP6c4gbVMsVIkMyJ6RR
4xbb+mRoXJRQE0UtXWCIEYBJQ35tCJDXXveoogNAjW0Y9gCc3aBb679v/TkF
sEhed4Oa0CQJ6b6/MtLM41DFibv3WBZmN9I6BT0+jSDUyZpHn78BuBf6WdQM
OBsPUritGbINjp8KEGYp9QwkMAWNmKExi5DR2nhT+ko3I1U/H2QxBKNU7WVC
bP0W+5yDu37Ipb2orqgt1tEC07EGLQwKe8FolvuLF6+W/MQzn5umV7Pzn06d
j/cj+bCXnDhFhK31E1FgzHip8n0AAwde8Qno0znsFphrLdaiFuFkFelMKPId
cNHMiJnJTA9S4V0Lm6iie1ZNv4g6KU+OiP1ukm9McZ3ZmW4ZRJ/pikIsjpdm
gCRmHhvpTiZOSsy7UEaPaOdBfa2YTLKP6kKoTOBLgoAHPm2vhhTErVdQfxep
MRmxkdImHIibBnfsvSpFu36rV+FQioPPB2L0tq2A6pErDMimmy52ma2l4Vqm
c6wjwtrz9Bcy+5glcqw42iF551sznFhRxOQK6rHEfwit+iAplovzwT2bdhUu
BtJXHU7Ca6Zxs3FG0L6lFEwwy+c0s8MOb7ob2ZNTHQOeuOrLmeQBEDBBU9DA
duQUi9ncOeT8iLlE12nm6gd/LdNJ5/tMRMKmvkChO5zeRmPEmCL7DgXw4ub/
VQbSrF7Ur83Aqa4PP3X7/Tmumpk9wsD7BRLWkyFZ7AF5XSSWoZGTf5Hw5H6W
8KKWO/hksJ4Dh837Fbg06w06X46iUWz7cVXfbrQQxbMby3iW7xN+vGocB8oE
NdFwK0d/qmoibPOfd2/5eyLBH4p9xH2jpH6FT1y0rRy4h1pxgczV3zsv5Fai
K0sRSDekeLqegmQVIsGyRPf5pghrJyzbIWaAJUxuCudumz3xjvvgdRGrCqdK
XGOF1vnhMUIPXWI4M/dK1yqh6EabuPHkZNnbMZ94PZmzTv8uH07ganHmNu6r
G5bp1NqbHIEcMYEi0HxJiRU9X6olNJ87iDICHfdKDb6BO25zjUJ318fdKL+8
YOmK/snXJllE/Nv8hA3RWfp7haqC/vQIopB92iwAqxZoLArkTjj/LgAWctOX
paJhHBv/N22W+bDa0/VaqsK1bG7VapIVAfftEongkZ4IEsVN3TXr2piU3V7C
0xzQ8xSfIjg4qsCHLt83xL0sktgi8U2RBL5gHycvq3C5UzQnz6KJvrAMW+Ye
kbQAh9eq7lcFDSdUF86ztv3qRAqOB5KHx+K6+AoWy0+xzBILU9dXynin3IMc
NJjq4ou/VmYDigGXSuhN7/+5DWQ7jWbDg0IzUzMorRYIoRE5k/JBtf8LqYSF
pCb/6Rx1fNDH/mmyAAMcOSmMZPqjN2VzcS+9qFfPwasL1hGrjOHKwUSyWcfQ
sV9hTEMBp79+ycokETuEOD8T9v0tCkkON8Q5k1wPbpdLeyckFjYvVU8LgdsM
p2fq3BcThWaMaKjN6Nmb0sAArpMnQA80i4LJnMKVTRlEXV+9SCJ0Z1gCLP9m
hLTKVwaVvUVHrkgrGKYtSkn+0/R1sjZhTV4M6yCTKMdmj5Q2XVsqcNnVlDeT
yLN0aOvmDBODKqhbXcIG2VbGhMT7JRqBd98rxCYv1x4rV4paozjRNDFB7zSQ
usp5Ebh6qXMx2XI+x/rb1GdgGQi5CLGpLzstE/WHZ2rnDIEuncJGdltzZYpa
nusF4UO9mpXqGymgaso4v/r13S8lGXcF5FYd0AFbUdRVKilG0SJ8w+frXS0e
MbEB0JIQc0cMsGlJDW8YidXmiO2ulq+qKigCT7mgZ5LonTlBzZDuegsvF/O+
alIu/sTVrlcs/9r70oRzoCelGjKAzyh5Z5LHSRNzj5Hvx0BBQRkkc9UF1HrN
iTxu1Vn/Rg1qV1V1yGBS2cf6A/TDeXYwwyItOmsfK4eI1DRievPnikZjJzKU
rOcGyn7K4ZjaFlx+Mc6NX8gPoff0ReDTc0vNYF89u/jSXfjLB3+qIIHCBVKc
eD0UwMlXgAlyoS9O56G5TGzE3+G9VHLXlmNLeWSuPtedUL1BbD0bNdnlCMXO
kZQ7LFMgAemJCP/FBpG8lZKxVHLklwdGf55A7MfsnlB7dwhSCjEDiJSB0avL
yi0QwLUWhmcSZ1Sfw8RKuJi+C3OpKSF1uvh4qTIOOHuxFd6YT+guoE6st0z5
YrNbivN+oIeKNegmBaPm4YTAPZ0swepRNPVi9/4nFr5xNcgGpf2Ki6WUULuO
y9C1hqLNZq0csfg+avEL7KU/jGk5VhKwhwX3h0vXumGcY4iyrKAcZgcy8VWO
k1As3ud8Jth8v3CiB6SOc3z8uzMWXoL9tsd9UysN2duwwGW1tOA1bEx9idy+
wvAnuxbOGZ3nqFRuM+Or1l0QkMRwQvNG2FtVJ19MA5qpHW/9JS1g9t3Rx3Qz
bx/XFy/x14DriqcT7FdQAnOfYSWD7ToaBjAS4RfaZC9HDX4QRcOQrw2GNkDq
lh6bS5G7qAM9TTu3Y2DW2Y9EYtEfKrnMSO9hW0GsAr7FS1jic5zXSQ7iF+D9
kxfIgYFBRlEIGAQwr4B/w4f6jhjG5f6d4U6FvMX1hKaCoWcYQliPDJuBxgGa
VHCEP5hsKk/1oerX2XDuCLsZiwFW4bZmekwPR7QSI7KVNvAHCCbDoISNiDU/
iOaGQ9jHmMzJNcMm7BfCsDH2uMnSdRjkeCbj+0TCBuOY8BBOdInfdfZUe3V/
ubpeIeDvZ7uiow6ufhqaeGU6IHjLQGH2uS9KwBoZpo1tEZcfIgK5PwFYfLkl
RcH8SrwWq3FFg9ngxKa6V+3LnvgCiDTGsL3p4gnV7HGf2EvadTf7vLzvM+Ur
LFvVRvDdx9UkDG6VMQBp9JzaYp7H1r0xSDQX0GiGXLNBSg/RK/UeGrqdKMrp
ZObM/iLXmIJ/bqlhm3w106jZMpsCUKOdwMMZpQeS52dj0obFXcT9gtw5d59W
PWw9F3zKPjFNpXzYhku90lNognCKadGtaQF+GW9VIdFZRajhYaPBGiCd89a3
YWNrPYDvOaj2Ew2AFQeGv1Kh0dYsjElBwTdM7hY56NhLxxCnoXvazcCzcAKT
/DYlaXAWw8j9+ytttEtD3aUyvXZ9U9ZKAiRciaZ0/N18TaZSSvyIWz4cNns9
icBJlaz/e9elr2KZIcL8nZsajaTM6fpLBY5fTJ/dF/e+1UHpvmucGDuzVwMg
58NAot+604GVFCC3OCw2HtSx3OS3VrkhyPe/Z4b/P/c1dBx2DMpyjnFtLPyf
mtiMfZbA+sNDsA8VyL+h52RRiaguykroor+jgC7ynrPiiT6TtLzB+MCekF1Y
0TAztNsOpY3zaP72ZEdP1SqlLF/VLY4yWU/BofqzYbO6T1BeS33nJh0nlT3o
rvXgyPNEnzZaypbYyS/ASSSwe0rYPZe5kJhHbxHD7BEjnW6eeo/6US3qu+dI
ds+0gKfbP78wYJY0fCKlL3RzaRUyzrs1Dxz4WLjlkJSEmFpiJrAKeuA7m6zk
UZTwq460NXck9rCodH9vmeS3EGleyUVWiICgKY0nF7MnbSAJ7gHBCnTKW9Y/
uwsTNeth3lS3SQhF66BhjiUtZtOiWYlNmHEnq8q8BAG3exdTfEG1J8w5iPB6
IJA0W6whhbolTa92lZtDpnR1kI5UVMbLQRTc7jixUxHC0rYx9CkyKu8aBHSZ
WVZOqkaMHS579fa291VAhgjVkCT1oKLUWivP8cZ4P3zDNPdESppfue2MQu52
g1tIZ2hoXpXQHsYiJVV51olWolVTdU6xXv+zT/T/zevMGfVD3vxl1QhDLnb7
aMxu02A7ctACyZCwA4zNwESwY5h6cTtVuUuc3RZa9n7lva98OkrivWA6mal4
ZWo6Rd/07ZsybiQ9MSVW5ZK6BIE3Z3QUDDLzqwV1AKb7uyir/PBBm1cCFRNG
UK6pwUiPNeUFrXq2mrMeysfHa4/NwlbOFLWHItnqTAPNtNZKldXf3w7pfcMo
Ymh6tOXyxKsBW9pkmQH/Z8PHFyfsePeXFtp08BF+kVNDw8KbCrJV7xbDrbp6
toJF52TMpp2Vg5lMObVcCsYuqs8N/jDRAj2EftXt34xTWpbs0YmVFrUKvoF8
2oSdSLCPKs9tcLWZtkO78Jdufqjf2Ts0kHiCm/maSbPr80mz+Ne2RWm99zkh
8ryqQyARZ8a4yTgxPEEj18E+c0YAVdce2OzVlHprxFj9c6st9m5Ox3VdLt9Z
m8pc7iwYbiTKi2AalDuX7HmhtvIfHm9TQC0nEXwohrP5dZ3wTZEg167CDlLs
i0ERdn+M/J9VJvty5kZa2sYC78H2benO02BX9bM1w6teWkL/EDkSHFITof8p
ku65kmddqh080tvuysI782hl7xMvKkF9XVmCueNwkmD3J7RiMmSMJFxT4xx2
Q00EXX+kVcs+9iW9XgYObl6TogaNAS8Fm2V/6QD1v3a0qNAoFyaXzLH0gv70
6hEZkCipM95F9aW6aVSRbr+ebsKHo1VZKUL8HzXu6IveMlVVJwu0xSi6ynRU
aejB072q3bJUc6pX0EHsEqbXMFmFHLHkqidocs/l6hK1+Fsch3ALmCfjMQF3
r+IfaYDm+bzAiLsxZmWSzOjxNXEOUcwXnvOzWp0CYtvzK/wOP7+7Y5ChnnFS
tuqFXwkCYpRtTpF1gcKutcLPpuMWFHefIYDkEgDqOpBFUAvRd+mFq/3MwIr4
1qZw7z7JpjXFTdQDa+mRg0qioE7KZOmRn6NEvPpHs9RFgNx/eGlNg2KV9x+l
mSUL2GjXDLCdQU7cfZ/ub3g59+cjI0NklwAorA/cM1iGqfAVJ3NHklrI2nTD
XFy7oq3ZJhmlo22W7WYWRWGXkdrqpdTCNn7PD/8BmmI0iUJq5Whk6le9o+mk
IMtkcGWrrFC32TivdqZndaOOpp+SLrm1lU5PjJQpSaJbkhdIh8Wx40C747nd
Td/w9SWaVEuF6J1lno1WM3gsnkptTGOEmhjJNGSzZhuphb2krvqu2TDnlBbn
FAIKXLeaZJnWLZUoEVZEvzNQ8N4EJjLaDBMRDj3Ssb8GQEPOWxhExEPVFYOT
UlRrgPfL8J0Db8sW6MkR6+i4Za1E8BdzSffJX6kgtV6uXdvQHkQYM1f7KDTb
h88tam4CVP7Ne5cElTiONOvIxbPqfoaNZBcgGPJMyZur9dJeriU5IFIDzP1N
lVotJ2e1eK1phKmZH/x6YKXEjm/bkj/papqWS8AFsRmEMFsDmbPmDjrowFUx
Dp4S3On7SpdBBhIom7vZQBriUyCUWjoDVFy+EYH4AWDUjB6+Q26p+DT3BL/5
fe75DEi4I5cr6wDG4PigC926GxYdwj+EH6vSIsHePf674FSmIhjVkbIjg5FR
abz/8OE8gqV2PTbPRW8vYroe0yBjTN5xlRlYDmqLLM6kiUjMRfAQ2kZCrObm
NuUM1xujg/yCMRzChUfC+wThfGg4RBHDVY9pVLovyBNUK8P9b/6LjZ7S6Yrg
xkAKl03jz33h1D3dYXVlGJDGoOa8tNOeAVkPjcfbmHfkPzQbjn6jkby8JtTC
i4B8268vym4gx3txasDKZ8hySLa5v+xRn/cydYzg+82MZxsT4w5uGGtJQqsP
KlnT4xeRztNoYc5hy7taHuLYNRUbp+TlSQTnT9jZWcR8NA4aOzCgDxVPLPPg
JVJrI37J+8aRvIQL6ZQKuVN3jRLExOz5C/FDalpL2RAc6zkkb9fogq7J022m
G50PIn8XsNx4khuvyn9ANSRrgDi1csE13e4ysnro+87wD8bBaQ7faj6kw3eJ
XTbJEuTGBeZj8AlXnOdpGbc7PuMJm+py0mQlFE53guXbqAZgBdgfCe25tHgE
ltQM5t3OWlHFc4+48k/asQUuIceVnwA8zISMEwzTjXgGHaK3tdkSOKcBVA2t
gp3RKO9m7FzFDRQidEzGTJ++MgBmeiMcQkcOzTb9NOmaefEdRuUhOCaGFaeV
4/2ARQiJ1wg3On0eek16gqsEP+7aezV/8M54ApIgww14s0DhMB3/39Apo1Zl
bvrVDdQQboz1o1AcebFUxHv08I7hpMtSHJacuSvDU5DpCY5UspzIy/l6jH+C
o0MYTaIdl5AKYSRSeoKpOwfraqbXd9IWpdcPfJgB40TkJdt+hdYpJtach6e0
KHqKZ3C9tnzmtgl+2Osry7HIrVxWrquXPc8RP5qY6cd2mHKGcEkfBhF3DWGL
71IeFc2KzUGBJze3foU4WkD7nEhpkb8BgeXj6S5x9GML+9ja2pPexzVPtnbK
qTEyCZfhVz5hwRXCw9XTZupTqTVvMHWMcvIlLq9fG1JrURPbBzXAWqYk8ugG
S80ydn+gcX4k4hIqz2xdGfmrHKvlmnR6DDee8EC4slDM0P6Bei5xbZKcuCtc
4yuJIR5xyg3buEyCYAJU7Un/AawtyO+GZFhvvezO9PG0UNHLQEe/aMJnPj8m
Agr5sBxF6pt6frqHoK2I54TmjH24Df96UogzW6rYxbQiG+lS8cVPvhznliTf
MVrTqRHIW1yVtAd26PU6HFpk1+cA6oOuIbpsrIp9p8maL0G8CjBkjXIvg96g
ghosiZ70N0tGaPsSUI37LE47697grc54Wwrsdjbbu753WiImZmLHJq7YKOuK
aHxMFzyb4Y7UFxgArKFE1TPOyoe2X8n5cq6MP2ASvqkFdr8lRk8Okm6cqixl
tpStWBWm6NJrwPl1C2BfJoTpFviEyDvHlOxLCcnOWWHGemWTDLpAqnlGPM66
daDCx+h6c77r7E1zzKwyRBYJw4FW0Rc3KUtMuDYx1DvgI9DUSg5xku2Spi/p
pFIYJ4eAgXNkN8GJtUOWLRx//1rTooCaxfUMZPTzq6DGI0hkduAgzHMLvJYs
zaFgmKruxYU6Ee82k46yyVPPf4BYewnrX7aXyHuO3RQN+JLxnsuBA4JJ4yrE
mP9ZECIIEJ0hLEP8hjgwgAuPvKPrNrHbo1aBJC30yR77A3c07wVbn0SaiIaf
XYlVHcF3id2Shx589uxVETLLL0dPXQMU2HI3M4z0QGR3ewWDa+nLSFH9s5En
C5d6KW0lMJ3dQ7UWwZRs9dpqgJatkU1oNMkvSAL5pRWqe9BaBJ1HquildKcN
OqxevkZlW6Uj5rfbcSh5xVr8OlGrOIF/0SXdbk0cUr1l8a2IjCXiSaWwNnzL
1WnirPGU7LH0JEBj955WJAms6ivdlHv/VsKESsnltz46cKMPoDXoYU8APMnl
hNoGfP1HY8X7qkRYjO4A4rpVHt6kRSh7Pqjmak4oWt3MqSWrZ2FB6XZ+pfXl
L6UeYj8ljXnoBjCWaUJZl5AebK9HQd+Rc8tUlavhH1wijKwQ3XE9mwr7Q9jL
QsJnTZNRAe19V6Cu4Y4FrYrGFV7hEhWVDh4lg8Yjm6J4Np9EE/NQVvo8cKm2
o0SwOw3y1tAH5tfpNzU9iuP/w1JWN+W1dwKO5jqBIcPgb3U66bjmNYW0iCs8
bYOaVlsgGmaxPkheK+TeWjHTgrf/fuBiBgmTyQHq0wFQCGB+4UEXlaKgEAn3
dkTBUi/50qGr7WsNJ93v3KVoST2jvZwozkKzCG5i0pqhJLmxIw70aV6T6OjS
uwPBKx6iuG5HfDv2YCAURPLDpB56pIpv1duJ+ZszIHJB+mqbvaTWL90fmPWy
WoduyM1UjIDX1nK1eBOx4jZjCekj1xwao7uEnfcCmO+qkf/fWl8lUyPe9nef
HLH7BYVl96rAfmBsNP659QBSON8QYJlHxn7GoOyjBFrTxxQG4t/Oon25E3Xz
ehO+sz4nnTYx8+GijPZYfekX26EiMv1ILNPh9GdtVTpR/bDHVpEQtlFFEZgv
JChFuU7lsDTy8swpnTTIrDBUDQoVZBFuIdiYB2sd6tvYqT0/BTwhJVHwpwOs
zDM20a24pVJ1t8I0Dk33ayzW3rujGLEeV8/3SGT4SsvYoMbu89XhrYf8EU+C
Zu42mq/tjbJ1oJ4I5GigYQWmOzuMtHwBUa2DrIaGJtHZN6kiaMRN7NTM4zli
CPcoGuy4qE862IQn1Icc5j9eWe74Bo050YmP5fL+vaWTr0N0Jkr4LBkpqPt3
0l2KLkrLb6S1zc6EKhHgSbKpj5fpoCXdS1A9mDydOIKMQrVBI3DZpCRedCUK
r3Muk5yeJ5EOlJbsXugSV3T7INoLLS/YvN6dxDGRFQwiuHH+UR+aZaRu+4v3
EY3LcfDTMBjGhFc6zj3cVSfvlxXWwcwb5oD2vWN6KIORU4UU5thuS6vjYNuY
UGDShik8UU4izyH5Y6el3iD2FoNA2N+7wYB0W/vNzJO6pFixB7P6h656d7eE
SPFZgQAJ2NUSB7VGvkCyY1QMMrfY4yu304rk9OyZBt8cE6K1WJsNkA5tOOVb
rYr+Elo+Rhax4ehAVK2xPOFVPScwA0R+/ZLEJPfdFxTLjMZ679mrGX3wHeBf
OgG0DtWYXK5+1T3JeSQSbji9iwIcMsmmGVXmxgYcUeyxyOnLDyIfq/CsN1yi
7U3/Ar6LNIuC7Yi9JmGa057oNMxG74oHVt1ml0kW38i8MkSlsp8Gjk7qyL2S
bPoI2/Z3AMEJOVudhmQgTRrx1IbQ6OI3qCaVsHsCj1VgIaIibeQjNVaXdbwo
klRKpemHgEnUDwz/WeiB80smUpPChrLF4qmrl2906zOon7L8VEvnisce5vAV
ZPf5FZ6g91re18C3PXF4sytS9qT32IhS/P22cSF49kt/7e0LYTGjapaeAoPJ
Iv5U8cc6ZxKQTaflPvbjOLtCbkcoayrpGxTzGgVplM8oVuwo3HY7bIhilsmC
+5erwnlW45UirQN0bsYXupC/XarCRgzsXRiocw8Kd53y/ZKPApCzvxanhMmj
g5W42T20wuANab/StqPdSlPHNWBhoOF+606R4iB+KnJewO7MA7FTe7CjAdYY
/E1DplWuYEHk/lCr2aawt3iyaCKBcAz1D4ONDLQS2iUR4jTjpn4/lsYZxkx/
CqxWdRQXEjdKJiqTzaOfZyrXSjsLHLgbE3lOxh8vEj9W8lPMqWWyg8zwxEOR
VB5GddYrcSRrV/8kWtVO+re+52ZB95QHKwymBEuQZM4+XY9LVk7vkCZEfnIL
BETNRZ2lJw9V2sf87PDmt43puoZDlxnirrNkySDTJt8Ao/fJeHe855wg719J
DCg2PfL2NyboLGDb/3ABbwvVtSztRsTb/QnRkdHXauDIp2KDy38cXHq6Rc3s
h4jB2J4qqXYjQYUl7TaUeXBOK4BR25Un4xfdcNGLzoHj/cFz1QoTwmmaK5p9
xKtEwwySSh3J+Loh3d2eXLTrppblvPHMus5cAungwWblQs/x1DDyONoOEBF7
WgRvw2XWYWfhqR4f4XRJBPQdF0MxuYpu3+enIKkcoLQLOW/ReOZHcyI2nWlS
A+WWXGDFyAsVe7WuTPtw0bh6o/DrZ1VXLKbBCR6DioNd4jHC1ASs3Y2pHHDC
JbWWAul0WOn+hxTRpVXfsm4I7WVH15Ff6N22RQ25TBH/CmsS7fJs9qnSf1Vp
QNFcYCHP5Lwogxm4BwpEQ9OAqJAwWVFn1QuqWKY65h0PMog7UeO1jCegcOjp
0iyWvQuom8+j64de4yQ3VL58oppz4cp68zq22tWNnp2jAVLvhUcxpIMSiDt1
bJIUJ3Eq6nxFv3Ucfam9n+LLH0Z7vimSRjo9KVAVDW1jfXYd3OTScZTDOf/V
tU+mfz7w2cx7wKyl3OKXTGp9ZpYw1YqliJqYU7JKZSKd/tiliMOLLbyVJKJG
VcmD1Ftsbnu3sfnx1/49UCeBExEPmNf/EhIgJn9qo527STjmMgE2TjBMlxgL
7lqcfcCkwYK8DeMDWJ3rPOnGv6SfrqS/LC3Sb9lBZTgeQy1rVDokT8g+mM35
kFxM5BYWg5GFyVSBqi9xIX4UsHrn4y8h+ZdRmZM14bs59uc4AnfH5QjNqyY5
Zz38rqIaAvX+62rVHp7H0fy5efW5Yn/wyYHCUy6LkoNg6J7tCqF77+0l1ixT
shdDMblB+vt8HEnU9fu814GFDYax+Fde9wL6YzwiLNEvA1R8w7Pjcz9cPf/9
94ozHiMl8dSLpi5PyMKPzI99m9Qw6Fc9xn0RZe6/ofK5982SnqwO3XOhxcFs
L5CvgAwSSsEZq7BtcmKXGb2GoMqWDR33ypP3s2QWZcAEv2i9wPbW1sGZKIsu
Pd0M0uO5kvoS1SzS/4gxPwQkizWJWk97R75srH7OoEWe6uaXf2645t4bqCqD
2ueP5vwg+p47x58OgHDbJ0JlNDIe3gcCVGyekGDuV2eSg/bt8ChYfav4eEmA
XKa5DT0bhrZJRAhMCWQPQrxCXfVGIZeR7goNOyO1rRZtO4dmBzJmt03hkbYG
oApEF0tpirDteZLhqnA9joOeVBoJ2h9ULPsM42KDLo++vunIsys2TDFSLJlM
wjQAb3FRQgdcJd4MQC3Tqd988uxDOw5ALwXqzn2GDP34Mtv26L/erq25qO2B
Whx9ZvHbvu3qjnnQmnVo0cnrAqLNSSp82+sXyISHZFV7D7hntPR7L+wyu+9e
seDuvuLES4ZQb1E6NJ8+TzNaI5IZeXCaVNE10P1q4t6JkBc6j/mF9etex/VL
abUWOXZAYArmm2DjMNkbOaudo0wt9sKdHTc6F9uWlgSSjSg15wsSazKk2YSE
Pe1uf+FXV6RuBshgwaMlXB4yWurpf8rF3/bCpjlMzc3LYVt8epImrG1N0GJl
MxFuuhjp3O10yDa/rhmfqSXOJ4y2kZd4HqvHEOdSyp3trGcn2feZGvqlAj/H
kVX3IeU5GaX818d2OhWTNX1qDsCI2dMNF/c7E+SNZqCEUX4jB0eggRl6s/jt
BbBmJksvcUOoAlo5cfHL6py7+w1xsvDQyA8qsmN8tuVOJerLJmdMSdvgG7gh
l2RWT7j4YQtn82MhpUX5heuwd2eWlzhdDdGU5YlXe76NPacCcbg/l987+lC3
XU9CCiogucnWLg3KAUwhoAw1HDyZLb2aw+X8MQbORIkYFZQQ7B9wIdzgu0SV
Wi1G/4P0wafbTKg7Psype3XVbWR2KrtGnjokGjgEobyXGbvoBIeVIRcc5JgX
fK6qRLvM0yHoVRum/ARdCQaRDfcL0HFCZZjARWP95UJYk0bnNUSgwJAPWiyH
ARcYs3+GHLNhxc83CKNtpYQZUzOJbiYwqkcZFwguUWVwwgmw1Urm9mnpNoqU
bdF4gOKWFQiOiIPAxY3REFW+qGUBdpg9JD7FxE8o3R19gnskVm7WnpsShLMb
02Is3y5KRfpZ+R7VS2shJY5QWNBY6/9kdn9s99hokeDkKYWD9pjUWU4L9Oew
gKvn/K18xf6UprOp+pPU38XQu5kXtOaYzkOTnVI5Pm5DUApNviS4x1K0ERzG
J4eT4QSuGZRBQ6Uj2Z2cW5IrFyMKj8iCwEDRUjyJ0PshE/32XIb36EWEo0kh
7Aip4k4L2lI/Izy/8ZiHuBzuYkr2U65TwwmyvhIfrgQqZTop88ar2/hEzy20
knmBlupP7m7b/p20Xf9tKuy0Ig0Uoao1rasUTBNZZpo9wAL+NUa+rC6N/bWq
CVy5ZL2GDwqY5L4Vz+yo10ayZt6b7UgtqwD6he+Dkl7cjCTLrqerzxzvmVi0
LIQLLdV+8yqNxwTM2rK1VKZXD1aLSdGxiHKGeK2zJb7MbmCTGMtY7sxHqrRk
I9Im3H9IFo1dvMnC/5M94dYrqIm2rmdbyybtD5qoqi6SdPffrMdfYKTmAl/g
5oR/FLWueO5YQvnsOagQU+h657NyYg7ZJGy/vNjGT2/jfMphS28k0Z+Ii8Qf
fof4UXx4WRnyoerYxp4S+rKMd08p5DhfCIx9pUVS9ZGB8gd63WmAN/IXm+Ia
P2r9viqYepwEHnHwv8DktuyFkLZlUU10gvnOMu9+qsuMNZvW4V52HMa25Qga
GQGF1MYUzaJ9//arUsRRdEQxBElf9mqzokajmn17TAhxT1dFEPOhSyw5Hdm0
tf/uUkclS8EdM2NyGkOWEbJUts+AIPw7muLUocbicf0yDddR28ZQGz+eiDf4
huSPFezx61TyW14zL+m3fn3BWItsnu2V+c4vSyr2rMNwa4rjL+xd1BrkVhXp
YYDhmHotJfLosbRc/eLME7HdIi5e5btvq491A+egrPNg2cPWTEQlFjg4cJ3c
R7+UApgNlg1NcPNEASUm1XP6Yh06DK7ynRz9a9Gtr5O/nRqjiL7Xi4v+cVQM
Z/TOC0L41uDgpZZeyBAAPr6LyqRt34Oi/xd7vptDx82aDgZfcaym79JY8E0n
0/DD+LDJY0hJv0NE0aF5mLwXzhvfAphF4IEAaq/SS2AVoHNyEXc/UEOBZnZC
FnEeV+WBWQObjUIAm3vrEDB2PGPnfSEQSGkn+emFuhGnofq1uedv9NgWnX/+
rhu9tin6eo27rVHsLkGz+NkIB8SD2Uqda8fSMrjDZ08jMlVH/6teufYUuemp
I0ppQy9IQz/8ELvP2hAGGVIRgV6k1FzbStb8gjavoQ/sfRsZyCA8OaJtDmUM
vVnpkaI1IuOwj0aRCSwH0H46NS4BvtgAOmNu5FjsUoUHWk9PpySe2DzRw5F2
J9C7GZfkepHLJNzsBLI3fnbYlR4tjf08Ar03j7tBKlzHcWqPPk022sE6CG8E
yxmxSK5719JbOv2m+3EznDtdo7UwuKMoKeEHZB6zecgCaLRw7r+ji8Ltkjz4
vCJAbslJ8B+DwIpF0cfYF2dx0ZNCyuDyqjvbWJnNJlboGo5ZjtKz0sCJ6hpa
6QmfUZpoBYxI0J1KyZ+dm4A5QCSmlpPDfmNr6pqu4oak3O4f9R8I2Ii0agVv
OviMCDd/bnpLT8pao4ChV64e74bb9KiftVTPcua7Owrzz46ksi2telHVJZS+
nG/q4VgrMfm1jxtMFCv90twp3sXV6OJhRAvkJ204uTuKBpOAHigiqa0EL5ZM
44RlktRm6/j1/sbnlGg7bzg916cUeJkHKeQajg9oUP+ovYiwY4AJLFEyPpQz
FfCc0uZf+yMc1jJm4yjxL7jd2UdoQov/H5O+WSkIIBKE91+xY+ycnh8uFuJ7
ZVHfcXlHsgRdillbz7rPMIP3ukLpAwgo5olNBSq08VJ5/U40bsclAQ08rN/F
dmbHHh9jPq3SUgPpueMpEzlIsouebT7LNmFksEv1Qs6N+zBcYEg/wiQEWQLf
tD+OiFsI2k5S5oezsVMQ44a+D1Zi2AWec2S2M5QDTKJqDnvEPTMd4U/b50bp
l4cYcwVscLWUM9nwJdhQjWyj5+XgWpVB0e+a7+eHTXi2qhssvEKDTlYXQrvw
cp65f2aNP2NGMUJxQFP/mUhijOBOzYazzwZo2zBZPezesXpaqJIU18nKrffu
o3+wsU4lbrQEYgylN6Iz4r4ZUXncRViFuMA89ac9Rrer39PQv2XdllPZ5kNA
tOL9+HBJgUO1E9sKWAe49aEHRyBQxLbbq9u5LWLtpDYiFRxm5FS554UQ6dhG
GEeNDE5vCRoHk8i/DarW/Lq6eJMv0zeGmOR0xqDOENVhN/mbX2FWEmW6g2by
ytp5/IR0POXdYCeLDnwjMPlff6DzDVd5xrxbliN6UCQ4ZJAMURTioD6dZ4Ub
VxPY51y0tA27PEpLAmZLBkFEo1yYJ5X1Q+zJItHNhoJwi5UPodZI1e+T/7zy
iQUOsorf6R6QzyQtNpMIduzFH7kV2swX381ohIjoFk21/uCiTR15Cdka51Fn
tyG+pz0VwdwylP8FVoxC5/7zmqDujnOdfMvZvZMVTA8klC4OoQ19VPR2BPyb
oIkEjlsndzjAcphPwSGQBRCNk/DcCi8y0BkILVYf1KTrwu0oVD3gu/v/BFmp
QoneXefRIWkvUzRtakXh1KktOGTGi3MhX6W5gXyuAmZprzntqsYQu4uKOD54
YGH8C2eII5zSme5HqQeK1eULMd6QpsQJ9DzC83FLpfvts4X0oxSz1vPy1tzx
DuJCoxd0hAJuIzdOi4Z4gCh8J+nZ3cgCz9jXRFtrmWfxle9a8iQehsaGQU/3
zsC0AG++9RKtCL3lCpCsB67nqiikKwDP/OdKwajSmNE/n9cW7ZLXPEmZ31qj
7rQ8tgpOWJoHI53kz2pRnxfL1/1JQMj590SENsCRd9EWmvxr6U10C0fCwYSL
XFsGkdXW01/+vc8oKF2aDAZVVsHn79mTlb1wKdL8RiyosTg9grDRfqgkKxy7
H0hX2GWIY8l/FSXiwDBzy/ZJp+KwJr47IwUZAUWiIJfmuUPJVujcHa2HDQ2Z
kkE+mLSPz/RopzB1zwmpOHJZq1OmR7831WZCX1aBsOMv5LrtjhIJZROuUQxo
Yp5ODNSiJ/G+2BunkEcLe0eVNPhJQsUhKdoHJDp+nY4iZppxE6V+HEuaqaeu
4J2IKQ4wStXF/ZcuNoVZnm1gpGJ24Oh7mAUHTxyxdja8kdTxUnSdh5Jj7h9e
IQM0U98kmTttypjzj1m4/GfDRB2naCIQ/H1t3QgfKyCjH7hIjo0By1Z2Rx9v
wtszPD6EFZfzNZuY7/+yr+XwqOG+Lj0mYqm+qI472tNrWZ7IjV8t1a3kVsJU
btC4K/fBEqJyJd9lkgYOFmgnnJhMgqRbpW+UFsUmCLqTXgYJu3bEHMVrNnnC
zgK1uoZ1DNbu+A/3VewNvcJGbxvV9pbf147qu60drJlfPQOzQz/vAbBXY/Rf
d2T9W6YgS4Vj30z1CzFXRdbjQrpIineY/pGD5qWwcp/gcVHTb5RkcbPrWXJ9
MX5q5rxxGD19Kp1tQtah+3jT3xrBrzt40fSQqzruY/IT1Ktqhg/aU0VUzWmD
a3sUOIDXr6NFSMuwQIRrDhWueirdRB6Lupb4ND+0C5PEv0tzuCqQP/KV5Wsc
ToEfQHWOmNiejGHCB4aB3I3CPWtirXYxQOZ/tIIgXstpkDmucqjLea9q1cN+
GUJo9RHUfQVsUfdl2j8gav32THK3xR6W2LRg/ngVdrb4qlJlCAwaWOUSmzqp
y0n5u6xev4a3htIXn1jDstbaDByUT0p5JMPd6g9dH52XZqQJznKPcaXxP5qA
q7sKdCWMBahO7Ax3JtKKTFpO+ZYWDVJflPIAqeyRTnL1bmbxmOTZ6YEg/+Bs
jnQXFl04wkEaMYOfsf+bhxW8CQMXY/mmaOb6DooNFQqtL989CWE931BVUefA
5MTSQKy1eHpVs5tBCHhUAByl88nVVjkB49us3bI5BXbq0St1EwJdxgZ7TR1h
/tSxLQL8kSTeVXUgs5NDZQcfdux7t2MLjMLUcEOzW6KFac0f1SaAt/e1SNpg
rzhWIRdamfTrP2NE21P2n2YWZkPlb/te+9ts77yhbFEl5m3NdR1SYzjrqIab
lIOIrbYXqphviW7i1K58bhJ2LigVU16I8M67WAfV29m4VKtF/pvNkWpLss7X
69XTOd0DmbqTln4ktlwkusKEJN5Ynrd4uTyux+aOJTfSzlpzMCNqll5nF3+V
2jAmOXqW9WdYnx0xcvACljEr9fepB/pzyKrLOawHLLp0kRj34p+Qe8F7eJDt
9QtXbvbwszigJssidfS5Qf6S6ww6gRfnDOcjVX3rx+LRYRLuvzA45jVs+iXs
zrGsMvqkhyWVF5zYws5fpPPr0lCVmyw2tc8ktamGM/Ij9CI5Vdizl6l65p9p
iu8RgCW5INDcIZVzkWe1o7OUUrj2qSTGegC5gPVBH/fkylu0eSwiP5klU4ez
2Pn34OctjlFLqWKRDbDOVybQDCZ4LRe7x6U8kMABkmIgJugSEuDGW55B4TL9
PZiMhkEJn7ZdgX+f04xh57ckeQAsqUTDYb+whra3YdHM/1RXHiJvZ5WfL4ZY
AqTvyWIG7Em7Kj0umoLI/i4+AM9EcRRRrd3gPip4iqcDrgJavCKKolB2QweB
mByesQV8O9HIF2lpgGeRXlS/RrB6XD3jdC2al0yE6MM5WZsLmzI/PDCpRE7y
qyEx9847/x05R4VkPMhOn+4K9OcLJirE5O5oaA6Ng/B6LsSP2ZGtV1hsirzA
VEukdAIaTksVHivLEWvL0VXpZEDQr9ABaLYFPtVxBIn98OMaHUPoLfdQEpHN
mr4VxzFmSHGu6Rp2BCspd+/Wj9DghMJ6PqnexuHGQ5GsmevWKRBcG7LoPml5
kCw8mfYBt6cx+ZrYpG7UyYMLmk8asgd1vRshtxkOJK/HHl2AzBeNYL9iOIH9
3eJVO11YkUoqjXyCrXwsUbiWEdpH/+aaIQl1hdS0SACcUq+B1gqhiGOLKFhN
Ykyfjxj0OqdU4hJiOSQoLESzUFKiqpir1KVXA3QiKqwH9Hb62hs1q3gS7iAP
cvICLcynSV7SwTYeZGj6rH76wtMUZVDOi4i14nKvK6VHxvngn3cvjQRB0ueU
rsGQAM96GUz6K4jYY8ieMN13yk+UzlCYVEMuysZ43vSwHl39ed+FtdxL0QB5
9XjiNgYlZ39b0Do78nGguT+D+jxmh4p87KCDNRH6Q3y4/KFbYV9Keb3SGzDI
y39wVNfDDZEmu6a3A1O3Cxwy8MB3wosObv1rDY7M1sriNugsuEN+0bdOaN5h
25LLAKfPBOlh0RuebAcUw83hTAliakBQGxSqnJJk+Ea8Zu4wRVz0Ff1n/Ah8
9v9vA40DG/Eb8P/UAVpwLYl+ZRxel9+RULC56lkEWFsvLV19tF3On0WM4SVz
Q1vNHllxtiLC0YIi3teKJCVnyFhnjuArf5O9X9nTyH/Ugw6DO+dTa5VRZWvd
BQRo9Ukpxh0uOtSeRZrc0lCx7Uu7NezjhqndRRPxJwuZPYTpnV49vzM7Iwhl
lKWnt5/+eEJWI+Iep2PeLzKC8ak6uME8K6Mgf/JeppKFLe6ZjzRi84iLm068
LtcOF5s+WTJHzffXy+ZDy7PQoegh1xLlY+gvevtCrvfxUzQzYRqx20jtTqYH
GbbxXtbsFr8Nyg4F6isoznKbS+T/Wmz4pIzaku40EJMGuurqOjDkoZqUhFrv
+aJiao3Cvhx7cfHc75ralkzGNjYGJn4Ac4lU+6CgroVMq7hUKu/SSKH7wxJw
das1/X7RvDT9uZoTNwqApBvUdZCfWNz/NkWYodQczcjoSwfkikXZa7yQddYP
qRP6hT04OukQxPP4Fhsx32Zn/uLi45vf7CeNw5etmELYh5kV3hdLkSJOMKZj
LTcKWC25UJCodN9eypR2zWchlOBbngATxU5RwMOz+b2mcjpUgZs4IHsJ4tCJ
Nhl5QRJ/zW/7fJjy4q1EcfIKR07GEiDv66dqgAPUd0U+51uu3nrtGW7nmC2X
iKeK2m0gyajRaNOo0PJqgvl+0nk5Wp5gIlbsjyIkb5JTADlXFqY4wfQ2ucy7
tTehQTk9OZFMke7xI4CIeDpXQlZERYUItkhxvBoncwhAuCsxA1wtx5awCSy0
gMrp1fjeIWAKuojB68ruCIBQzlDImRVVORZx4qMl0GpqCs/iQXh19wvTBGyB
u8phIB6yLyq5EiTJwnkWNL+1F+3xLnRXKU+aE6s9f1GCyLgUMI3KIoZhMBHc
VqpCkFQjbd/1B4pPTqgqkTP7h30fXGZLtJGC+Sj/wm/w3HILyYTTx/n+MYOO
LjNNvLwhZsfTUQ/XKM7RiBV7HMMD9z5ZWg2X7mG93UbN9m0TbxRuFvMWF6F7
pfz7S62Po0CFXaAw2sIhWAOwoNUheqYaZjcZpJx3en7X6VYIEDUAM9e5ul24
afGQ3m5SGMTkoI5A2RKgSPOqe5JzV6BrE/ixHigSDARTLQ8f420xLrqpAxVR
kIHRFpksaBIpXu8KerQ344B50ezKRoBuHLHBLUVqap8CVKumoDRGBgfZV2hs
RhRqTpF3OlNNkkM7XsqtKPgAz2Tf1PThNaNyEG2e231vjTglUuHuputS8TKR
e1NrNDNbKrY5MVx6m/A5Um9+HF2/Cq45ahHtJX9QtmZT2XqRUk9NuuBLsBi6
AL5gb3uXR0Z7mxQMZ5XBUmZBpgV+x2feiZTY/KPah26CAerGpGVy7kj3DLwP
h/+Sknv+z4+ouDT0ze/fL8LvRSJ9oanO1S+vTUbo3+15TDRy3XCjw5nPSIsx
rd1boa3CsQcg5hSYV3oykN53NH04E+yXF51+yE+IyYHtm6gk7qjU2Ju4DDoz
oxROyWBKkkovatlKlrsQ7nud/1V4F6rXb7L5WHKo2zblvyS8j40Agv3lQCXY
An0myV1s3QMoz7MELGzqKLx1G7vAkbLc8d6eBqLRp1TqyBWseP9TapUFH/FP
uULZTDtZc2OA7yeX0Q7q5Tuxh9AE57tTB53Mo0s3j7Pwk6jley0RrHuqEJlP
ztZ4lHQg0ViTtio+qNSR887FMDrpSfPzkwTFFS3B4KnUEc0JoU2TYupF3Vbg
C9LxoNoQIz3b1Wel4n9y7EllNVH8cNqW0dloXDu+lkkw38mLN/ygQ+UPGdKh
FdPSkYm9k2g4rFMwU7jbeIJ9CoBSu7YPtADnD0ui9JcE1AJ2teisxJxOiTHQ
tUWxaVsCGbkSvpzYTqzRRsfu8C2gvg6uZUn0lEfLKsAS+8hNxWVyR2NY2CE+
xCLoG/Hw4VQHxIFU5OyG5oPJd+e2S/jNC4noFN5sLfr/SnBoPJ/6Aexe05cT
keX9Qg+7tAEN1TqXX3PBjcq8S8jfNuPENgyVw+0qL56y/XpS2yPR62wkrHF4
xdzRtIL21mryJu60+9HF2z95ZfaUWuE+8NBlgbSiHu42z9DYeZKqKbdhbkCg
MkL7I6ac+pLaQ9KmeDETe9Rmj90+/wBbNZ5J4ne0ubW2TL4s68QpHelAtv87
zW3NFXMNcDdia9tYfI4wZCei5v0KFgSnlRC3eOdF86yOymhHN4eElg6noaOf
PAAdpi37K+QOCWx9WMqr4PW9/yVvb0iBgrQU+rMNfMGfWYvIW3CrRmGLkf7u
0VbcEOl9f1XO7wHW7JBTwgCXZf+R3WJWfW5M5DEF5Cyye0J9YDU4AZPss2P4
KyGCTaWtGfm+18+9Q2io6YQIIsIy875g52ANdqSbP1BLJtuFG99jRnq++dcq
IQFoT6pc/XscNGnwvK8fj5EWwjbrWs4p3/WYYV7yX8gFAuYmJPSKn1qN5TyB
/bdY8Fd7+eyqq8jjGah1MuLomJ1LCZWXVsOG4miO7msiTOvFizVv4Bhj22jm
6aHrFZNll9CJ3pNCoS3xuqkyuWg+kAa4P6La/3QmuE1F4DYhjlhi+VE7cTHl
zTZq7WcUP+TwDaa9fooGay5sGKQg95GVYdM5GvrAkF9XBci8Uq6K8yoltDLc
1/zYPDQruLu9hNEbOwm/GAYAy2Eg9zVvDmu8+QiPZojZpfV5vo2vB/twbyNS
qYt3z/v49exufYJqnlZJLP92b0SU0sUKYaXYDWwdwriyFv5DZphSWOUiWn/s
0UJosw8KJAXI8mImjTo5cKJXWlOaIEcJGvOzt15KycrFdVpyfQ7vRczr92N2
DqBxanRQ5p4+6t01NhoU6cMFfeAAxe8e+m/nF6Lp5ZMGlOEjgjr2cy0q8d2Y
Ye7tOj6DrMTXTwdlAlORpDjMWyOwIDm75U3txL6YAdT4iQJbL1bySFJTzW03
lJODveofFIRt4cBLGsXVxgPJG+XblkaWnDcwazV9+rcAukGXbeldc5cQRmT4
lUhKeFhgY5jV3gsl1Y5ew4zR51lJoWNVwdp6BXlpfMUb6EZACvQ5PzzSsrEQ
3UnbN9HuCDVUZzEhfNRfd9E6CCDUmwY/MAraDtq4ukgt/0hNGrcWLbh0KlPy
5VXaVOxW8lo0obG7I6NlaWfZdwvODmKQVWrABc5iCsB6kh9F2ObVTuPpUUoX
GI8ns2I2PixGpeYqnQ/vC8VBt8Mbsa4IOMkt1ZXPJba/Ws3SB+l6Rire64He
ASLKcbd4bFMkgofjaWaabEoEglX9V2ASPr15pt+jNsfdVFuZpueL80w9DOd8
m+YM4/xSAgtTQTz3j9pLCgSSnAAU+gCQW1if1JoOJZwyXgF1Ip7DrctXqw7r
yIATJk86R1V+n7Q9JJBI74otkNmh+Tj1Xc1yQCi3QYJzmgkMTCDH8/P7wGP3
7dNe3HxClaYaN8YscKmTNNCFwPicsKhxjmaTalcjDKT5KK1HOc3+D/bq1KIw
voeE72J/CvyoP+FQY37mCSd9ERr+B5CesdWE2YmKCzC1PlgzToNsF/RVBBIF
7kFIHhCbOYSVBencrbU1NrfJVebBpj4qQfHc2l3osPqvUDmJmADUBvZ39eKw
/ml4hG4qzkzBDlQG+z9jomP0R/hyeFKNU/d3wScUYF6LbUbwabR9+ZXuYBBJ
CHF1UDRIIQNF33fULUxn9TUsifwC7rvdP8x6T5cLHhnr73zG1BXvp/5Ay6ba
Kofew4EXkD4jo7Q1AhnnsVGE+y6us+fqieR4D/IOClq16EZX7qA2bE+5dZnO
3RYCwpTWOc/+rR9lcWcbd2KbVjQDbgCr/eO8ZlW7/o4TbYQyE84P2zvrYfh3
sUjCmSOiLf3h5yQUupUxYFelSvaQbdFRcfxSckcYErOHVvQYmz8zvvlVBotx
cVtkm1KLnxE2jqpLoV5J2HTL9kpXLWgNIhdobuc1muZvCAi59ZQRPUEli9Pp
nT57sLezTaljDx1YpmJrZDvc38jHMcj/8PBAsiBwSsBRK+5pKJGubD8T29+S
fLhsfLcmRVG58cgvTPg64afSm4RNPlCqjIcWSwED2kaG0iwj3aF9dxj58AA9
AWTHraKMkFB17pJLTtoH6zCI2sbKwZAvxfklIZmUWxAzWd9tvWiv8ZCfIijA
1hkQN4YOF+2/a78m9NXUqBf4/EMjbD5EFVt2F7Qu1BGq+vDVr1vu2FFIlIrD
ZL/046ZXwg0R2VekUmk77O7E9I+kYV0emqWJNOjhFmu5cMU9AXPqnP1n3n94
vEFxxWoAZW7KMGDVGbfheS69DvWU/0FFUx/WZfltZ0r+oacGKYk6JtFI10ar
r6UEmvvhkiKjh6qNWYSg3pjTwFcc5LVhg728W2xbSxFT7af+N13HkMWrRFkO
h/NfRroUiGT70ifUocURSHgAsHTxPtiQMAkj2emcGc9QeYQi74wkq63zCxUw
kayRti4D21IzdzaHC4q2BtfAWhXF416MJArLmbyIaT8n2csaxK+vuB7+VSIt
nhTLDAxxuWCpYSPoBfdHSFyh6Ly4VCE//sMQDyaSFotZEO5bJUmePjdeP9k0
jn3+aLoISWNFUwuVtca4wFiM655yCjHTFSsZp1djQmeKI3pnCfgTS4vjGNZu
YFJ96HpY5o/Qs6vmcEzWiwGUctScfyGUkHKMqLRyv+fEGE+ZU/0P4y3kPRmZ
tBQWRumV4y5dZ5Lmd+rKg/pPLLfw0NLiWAILBNEbul+VLvbTgGeDSPfxIJMc
3mx3AfdaS4Uvf9yybUW05CBVUxcVgOn92k1URtsgX4ISZXS4lZ1cD1vLXemH
bj6fN8gLkHk5GAAkMZK5CbHJfiEGq6glIlE+v8MV4oF9hg+htLwxCKNyha4E
WAZy1B3kYDEe8apcnINrUtnUPC1px9Of8uRfcCKGae9MIk6FDb83EWlW8n/C
ktlgnBBZ5IW7fehSh9WQsTHn+c5UKSNTCrZSmpkBdEKsQdBn3yDES3oIN8pf
AJyxNEd/kcaveJAYTPz9hxcGTecv+SUrFU5ykrtTlsc6lJsqj5jAibUapCXq
QfDbHN1BEouy1CY36EUtpzzPVfKyh2I4cEHIwIKbX4DC5W+MWye/A1tukTYG
nV6/ENyaiEy2rhDlhQIE8iSICqkIllWz+ZggktglbdkV7pGyHPrKzdREFNq0
Qq4AUdRkX6S70CWa8UVmhIkB+mgl8g59tEzzQ8KLzF1zD27bOJvfYdghMdSz
VsYZA6MyWSUiq8/T3tky8dql2rLhXdzayS3Ic5thZB02IlBFYLNHxd8iGlF+
NliyJxHMWst2k9TwMB2fDrKiOfW/p4e/DbIQDF3eU6PnuD/H3sr+RtjoAFCG
uVstWOTf0u6+zMqSxM1a2VLGgGbsY0UTBcYIrHsOqyiPcJrz9blAs/VyrN7h
stR3+R+GcVqWEEgUZ6yzlBKJvoahLf5o4i4d9/5lEFi2uOssQm2nthem6JMp
QWLiL3O6H/vzMSUk6ChQ5IyfFt1LNU9hQxLpsGjVqnFxh08NJoF21dSgxY1n
n/Cv3F8suYqNpTPRDKkTMNErSZav9XLs+Er/iCQd2IJzHtjnOOcSpmLytag5
i6Ja59BGjkUEe3lvvzND7Z/OgfffJxFag+sBiyedQNZxbqY9CGDcBGMapT0l
9Oqk69+jP79wMSEklnWqX2KYXPkNDz5UeRjHtN+at9cgtUFsT6ysw4R0DiYt
t616TU9M9U7E2rKw9Fd5fvXvjr/1hM1S2ak21w9jSM0ohAXv81sbVAXo+Y0u
fAFX1qfwJXIYvQkxdHgjE4qdH/zkpZfBC9ZEKwYWKcAxXpEzyVX3M8jjc0mH
NBPZM4Mai3iRc4R/nL3+xArHEVFvCKAdDScTvoBBwGuJP8DMZPC9BZriwuhX
7BOMeKkAf5vG7xOW605/pORX+jr3C4smsYAkKR7FRHg5Y3frTScmL4zFHhOU
Gto7KEooBoLQVdJqxMfFjXnqbAmizQ2uhvjyOkazNjhKIe64JGAAvrXOAxco
N8b4EP7cWb5qe6o7MjzVQwP1SnUYlL8+Nz1/Emrr1C2+IFSbkriOLsqhFUuj
0qIBz1Q+K0eYINuTCkFsV9aLnOX+WcBSwmOc1/whw7Be5RshXg/VkSKPvfST
yp267K9kYqlzhs/udtsTOyWv7DVdyIC3562DIBMi9RpPWLQteQwveBDkj/e6
P0sxdmk2GwbmeazponnyBO2Y9Jl0aNPbvuQAxYe9K0c2gxP4zUdIWJ42pDkE
i22q3MugIIYxmn33Cdr6UAnzhYCC401DZYN5gEiMG13alvgyFVY2tXMZ5Lx3
JXEQx64+ORqoplsPkCVaVdkt2rwJCAH8GwLJN4QUDL3ozsuuqtZLB2sxeI0a
B+vw3puS1xYTojkPQWxlElKe+VaF+ZRTFqYeUpiQsK3MOrcGpflYRleVK25/
JHu9cCvzmp4yTgKmlIMNgPuux1laIfTpfAwHOUCjIVghnpZimqamV05N6mEk
W6XFoOu48HqetlZeF/FN7vDVaAW7BgwRyAbpfCrviEdaJxmggvsCKviSAR9I
rvhFoNbyFqPujgV1gRZhlbE1UfpPz/rsWsC5yj+Kj1WgzKYiYciiimV0e/Ej
KGcbZ78E17GnxV9N2sxhFHqh/S2M4ai3fW6v5XoZKi+CwYYgaqE7MTM+rpWy
vcvV/Yg5juwNxsBTRkAExYSa0FLeyq2uA5Fy19UMCdxGZx6pjEeYWCAhUeIq
DsK5NsXusB5c3lPqeLyi/UhKcRDJUNwFMFgSNc6JNjvTE080DHaH03mWOPto
54aPBUd5VJT46GU3S8KgV2IRLR0EVrhzvGqfcTRb97hE5xnQHI+csIzsw5Vo
XJr5oMtHAj3JhcxWNKDX3RBpwaPjDyOkUvQVrAFq9Bsrlh87CHxd//hn96YS
EMxgTyzFZA79tyZgp2VPCDv536O1m/lydeCEQkK0Ft5O3p/WxOAIgCfJBibW
MK8UBOz2cU5eTBZVjcNA5OKRiBhOx7zpX7+LKY0PvuzhMmEl0jAy/3J+tTxY
X5UjAWfhoU0jo1rbPyz2M/QYWPTOVjGhMzpoIHWLjvp8LNvNgw5PdnJL0unb
V7HF3zjH8K1r3l8rqtaWLfj3yN9pYzH91bz43C3kV8KlYtRvXKWbHmsxmSMJ
+M+8S2QaB5v/l0bW9vpoHaRNJcMjN6ATrn6yueVCmjYkIUbHJwVzeScY4pIj
/pFw/U4QXWuOmMqw2FxlCBY9rCgVd1c/8nZtzYsR0m3lF5l+I0PmgOk7uhZy
MpiFOK/umrfpD3CckWcczONfbK+QMUJTDsiep0Uom5UU15oIxnO2LhcJixr9
nAfI+3I5XTpqF3dYR4X1T/XSDFSrPRLNf65PRt1N/oGB5rnql2gjw4uwacME
KhpL3jFZkvaR23ZJTZTZi1nnHtae/giD5IG6tmj6LVUqvjsonrZxCP82sEMG
m0puNYrAc8thzMwCe7QTnXslT9bGVSOwe0D57b1QPfZ4yWoHu7qx0n6tkI3s
29YsPUpuwWazqqQ/bhkWYji/OR44gdO2woxU66Q+42GamGR2vmsnhlwZ7csC
Rlc2GeoqMaAJb6NpqZfy7jTri0WodKejHGtGHup7wQ3WBSCBUYO7Px9rn84s
Dm4lPAksVSagUNvB+u1M+9PcBuk/0PQAa+FEWrRP7xjYmBQn//NmfYotbdwO
aWDVbkBU6FCkpUHjH/iblF5mBJ5PduZzCrse3iBp7x96sQ3vQhb2vjoBOdpU
2Xxy5QsFpJGQu91cRhys2YvPJwUIJY0WwG1v7jWhDnkUFwIglyX5aMHR1FHF
S/tIRqZtF0YRGaePnA0RPz9TNoeEq60QpoNH5exeTpikv+y8xLF0yfFna6n+
v+ADYy6gLW8xe5YNIPWB3TGlgA9xzOwLGvbBoFedI5BnVdwqh206Vwb+4PcJ
9RcwnjswnivVgp6q3x5/03R6ZRTdlKwHB3e21A2IcYIEbqKnj7WlGwON+xms
SY9TQEUm5k1eVf5B1jUkJDWYXJciGrzaAuoFkc1Nfu1KRr2/kRuOtEIqrcbQ
r8Zy8K8EUMleFcsJfJwfKf6hUst9jLXnRMdSWjkIImNRFUBczwISX0L5iRRB
qapFMQoyaHYs4V/kGp5FEbwmL21pliy9iaNJR4VuNLxPf1+cH6OLYBcLII25
RjFnJhuaUxHaP360rgcl1yeVQksWgZn9p0FP/Z10y9PNxVmlSnR26ECNnWaL
+tJuwPcY3g03Zk+usSIxWEHmTbY6SP+jU58lLifiP4wp0fNMqBrfMiaDs2uj
AkDcIjxmV0c0rUEsSdsU3JSn7hSvZ00dfeClmS2uWXR9cYBdP8iqGPxcy8PA
hWIGf319lX9jZ75oeiLCxTvGnOT8YwOvE3vlKVhPLvGvHjfs6onGsEIf64e8
siaoSUmiYQPvsrLWUuCswoGzPi86IHN+QV6UJNNk6nOnRAnjbM4JZ2gqwiuE
b8q3iTEdOcOiOSLzzxIAyCTR6ZetI4h/LAfkEIo2dirRy5jbSNaDzopd6KRs
ehaxiTKu8Ysh1C2sJL3ic2/MtJTD18dF2Sq6DmYizzGhnLxfCTleQujqQlAl
oF2kR05tggBIrQ93SpNxOhTfS85Via1j68KsV0Ga4ZHhzeE+IGGGhEIDZ1hN
Ou/PZ/yS+frax3N6IEz9ZADD3kEUF6DkB2Z6OlDbVD9kG3JOl/UN54QlgBmK
cft4ZOTbm/rKwAF8YFAxxRGgR+rE04mnnVyTHbw160TBKsjrw953eyfHMFKD
GWfQ/0WO4K8Im0RRsWmX0r3ucpCaBz4yDdyqhVRBZfO0bMxraCpF/pAFG6xu
2iRRkUhPVQY6fIP6ALp2Vcz0W8yh1YE1kZJpjTr5lIPPTmhPskR5K4X9h730
8vLv7P0HPIT8M8eB2wDy6x8WbCoR9UCc+7V3UFWfNzbcPcBmgdJpeEsIeH28
I1GC0MdEQK5aL/stZ4DcJAY+lUYJxCkdtyCeUniHapcxNUPySK9sTtqFboc9
I3IJevu13Ey75Q4IYPRY6BSiSiCjmKyARm7jDm1WI53K83zJxsm4lRXPrK2V
oxz8ys40OeZylKguLQMKgjqptAzAkfwhUufMaFTMihda0UfUTAhXsmc8NqVM
tIjTJQmIf16o7B/D+xqXH+kygmt878l0L1cPvcHR0YPOmBkDL+uOlnbQmGC+
dZXsO9S1zE7H7u5B2Ij8XqtzkRUj+uCS1FEU3DvMHcP2Yu8q6a2ZWIXZWSQq
P2KDVIvzvxi62Ef3Ov5lFYortQPiP787hp9J48fvTqaqf+lmB8EwrvRuI8Nz
P10OCSmsGYDQGkON4mNt4xI9IJJt0Pnh+4IxZD1wlK9p0NqIjr9ipAO9xpYP
Cx5fkDUoBIykMwb9IgbV0j4HolqduzUuYYAw2pVbpEEbdZZ6xR7RMRJAyV2+
2Gca3JUlHykyKXanhKhqzCk9AfYcbxmP3V6uL1PgIdcEXEyp6FzHoTFuGn6D
1TfN6lBzUYyFS/KOTMvP9424mf33cHMMsy7HXJHk1NJHSHZHGXCkHRyvyywM
Hygwy0Vy/t8dqQCxXo0R4hAyBJZ9F/UxOhWpNCJH7QKaBp4C0j9KCrBwnuan
WHHzFar1RkWP+3ArjolRGclwmHvy/JRM0F6+HRhTZgomFMJ03SomUk3BiXD9
XPQn456sZ2BICONWTGuRLpdd2jBo773OVgXnhV9StfgFcGy4sguvjPrHlWeU
vg8jUREMDOBbFTW1AQ63yDV/YsHC5xNECoAiD3+3PxvQf7Ps2UBcZC9VKvJq
YVqVU8MMsXdppycBIA1W3P7X+ZkGyo+Pja7SylM8Ymu89f09HSKZnqeg2KAY
3+nXfTg5ku3SHEJNTNv0wOYmOIlcfgpSDIjZInb21cF4qS1HZImRlRc84LnZ
nIeGZgoXbOnNqFDsDbNBqE8ByFOVIMdMchw+VHZls3t8Ml2RQ1AMDXyGBFV2
rUoR0oF8NhQiJ80SeZWVW7J7HGi4Cpx7bQiybd0qskPz/y5qBsg9CP3gsR4V
RJiJi9/QBeZt/aW2VPNnFAKYJuNpD7weAQFOKH4NledLLX3PvitGdsh2si+S
ARMFzsWduyghJSbo7deubkyv1WF7LgR3ZTeoZWOsyrOmpZUZE1/SqzIYDK6y
NqGvkKwIzT5CgweGKuYpL3dNpDwOD9ITtDQKtNe3YDcWFpjgMPUJEcbc+BVV
+NBtMlO8PlsSEJ491jtXCDgWDNwtfa6+hteoxcKY+yzXUnm+kgKRnJOaC71l
RWmhhQjkxSiktPx/qs+K/QrrTCw5SiX1aR6jI7WbrvpjSP1bZ2ch5cAo7h6h
JddqxkpksfWZgUO6HV8bXVyYKXpX8VUHbZGKvu7E+Eofuilnw1a0+B0/YCdo
DEwqD2COInnLBhQqwYCgWlE6ZzTAb9hNAGspgS8DqYS0d0buus6BNHEeXGKs
Axbkfh/W0w0vU9B824npuo+oTX7pCk069keaibhCy7Tyhw2ItpprbwzYstvw
zQ3y40Ze1dtzxF/eJSZnnPeCY8guVkM028vOsAcxneF5fqetZuTGHyGJ5zhy
zCcOzsNTO9p//rY65thewOzpZP+6T/Qiq3xY4o8PWjOvZNaqlNValDn6cZJY
oTIQKqHnPpSFeC9PW/Wp/9yUyEuHqjz+pePpbOifVYvE8mNrZpwdI+q5QC5F
msffAEZyh1wLmHyKG6RsrKb/vDznjnT/QvBRTTjaIDB9O+AOHt46u9qpsCob
F2KsEBuL6+P3C/WfxjylwyfaA2/X8ZzXIuZWhTl1PvM/NWRmiToZjG1pEouz
6mLZIdMftb80IpR2PBnNpRpdIuQS/e+BInrHkFmioH1K0b2FZ10izAy130sR
LZ5ZwhekzfUT6S0TDULDXeSlyH8wVEMiu/Z0CkM3CjdneqIhokqgClw7PEeZ
tedl0Ekvzsq3dUlRPt2e4cn1zMhtUI0MZmkBqPH4xkl9UAbO1uh97YKgpFFC
FGE8+YWLGjGcpGP7vLDybEtjd6xtSHpCD4S6o5YxRF9Eb9MbWIt5Y0p5P6UC
3BFbUk/fRkJKxradHpDdK4/GxQ2WEsdPwSeNHhJA1HGhZJxpMWgnv/ffj3Jx
UmzFj3nnTyQtX9SIfMzyuaGh0T+jDTiDhRFk5qNalDsAXaqSi4hA+32RFLWs
p/JKsw4+1WigroyS7x1/4XdMUJl/Z1ruROct2puMD6T1CpM137hrpH5jX+Nv
YJ11p6ZVbcTD4vgLkFkfDj4Qyl3CCBbPVoJTuUWY67hHz8D15AMAlF/jTWyk
8IdQHH4YVPOFqcPalrhJOmUwF4DvR7eHd493F3EBVLYAwyEPWfTI2ivZzyTQ
TgVmGkzyX9I2Vk2fipboBT+NBd8TpfF6k+Z6Y0njWtgknb7uET7gl7IL9u4q
Y35G9VX88MA8q7/ReuzS+0+Y8PY9rjXhgut3bmDEdol6rkr5GxKTkcKNVKyz
tgsz7613kVFJwyUKZdbxhTlrWC2XjDTJ3RjINbQduh01cJ7Cl9R0AQxUX026
4SxPehYRgniS+lWyIey5zYUXJNExc12NtERiPhf0YQSaoDsIE6HVBY1AhCJu
z9dcSiQbZqiwLIe0aFygae32m3k9oxARcylLkXVl//6mZhYHjczQmvShL4vZ
S/y2Eac/82wyvBVNBftk8S6vTPp7QmIt86BgVxXg2jd6Fj1DWre+VosoNppP
QRSamsYWjKF7yxTLdJD/KmjVuF05bat5GuOKnNT36XNhPMpuM4/myjv6NUSW
ejYCNaQRc/wV48GBjv4c3KplcptwPLOfK03fmLb+q/r4fcDWW1scGAEaUE3g
qz73g4MQ6rMPLILMa1q77fMVo4bziAM8nCcQ4V9BwufGw+ovaUR7oq1UGjHg
rU+f7pouE0EBGb+7u5ZxWm5COM4bgzS1f+AyOBLqXwoMyqeMbdFbsiDGEgHG
c2GWpjlUhjIWxGsOUVHRILZRxgZMAMByy6f7kuYhb2qjXhsm7tWIzLDMFfm2
XDvQJPGRNXpjt/fijCf6JZETj7qXfhKxyo75mTNxA18ZrCI0v2xkmYsS1xe/
qR9YiN/wRkk71zWp47MBQwXjI2tSZhxb1L+N4jPUuzcD7lRKWcOXkymsntJl
jNFxECODWmcKcHBIWowqWPSmDhzaHklJNMmZxlsEju0rB9f19G1rCEWZTOGo
UBHDeeYjZ7uIe4/gAjDU81YcTW2ZqcYoZiPdz4kCEBr0u2/p8HS7mM+SOu7f
Tjfk0ihe8bYGIHakZ3Ev7KimSpHvnhKQ3NNauWleId1yKu1jXSdziSWjkBRO
vII3/qG7p8hwZCMAWYJ2jOwRqsSsAIeMfGshCGv9TyGT87etZTgpEbfp2x4W
971Euh6zFWwpdIWC25wTAqZgWhfw16Q4EiInM5lZEq4VCm7NJOLp1HWJAS45
989ldDiwl1ZUBOWMN82GPQ38i09uCIzUAm7f6Sit2JtyltORgc2hJUZWxqMK
9AuV7TwIxMFaMt/rqlXC+j0Oo3lftVO0tAuYkrdub9KdWHmxLpVW8+P1OjkM
RrO/0F05NwTY9dwQ/FoXGBVBwrgAk8NIegzDwgbd89nfiHBVsPyxxByjlx6e
fhPGIlh6oTkyWCP0KfMuDIarOnEALzGUx4skf87vpBr/AVXjyBIc6bWmdr5D
KfF0bmMxh3Z7r57tnqNyAeKHg2r7Xbi64fcnza+OQI9JCBP7WnjuMwMqiUgq
lpV1Cn75p/RFw/R3tQ7eB6k3cyl1vcQqLZIFK4sfiWUOfmUz9VKN7T0vmA1/
4KUcHFk6c2zoIFZ0zHGOWEWWu0HnAtkK9f+zlvypx1T6vd+K061/c2cN52QT
a5L4OZj43zggdxyjtVTxww78v7euXkSxF0QE8Y6PTU5F4k7J+6b4Yd1glx2Q
AOmRRaHRb/4Wk2xWwmHSlTQyoeCUEE/cAEehqw85aNlwfj5mCzbstpKldXaH
COblKz0R6Ka0SkriU+nZcuK890S6nB6fI5/npFv979ngzGyQjsNwjNOHS3gF
6kNMcloxry5t/mOix6BRv9JSd5r7NZmNmH989lfcq7joNaV9bGHFs8mX8peB
EoJTwVBOtL/UVMdA3eRksEe1w2gYUUCQcCY3h1CYmzzlaNj7Kk309d3DKW2r
Nee6c65XQcKTcfCEUrkbpBC68fGNjnAM9VprCeWtTbABXtepfJoq2nmlHHYg
D09+my6BY2ILgIWtqc7iN+1affejSS4CHpMZYOZGAMEOAfcbFVw8bqy83MSD
ugLUTrLv/muG3auxLsTfHe1GafvUAUMjHq1sGzato/ib3Dl89FA0IYqef6Aa
O5hm8aj92fRZAIku4OJga8AzSoH4kdHDNpCBJp+zi421Sz9oKf1WrsJ+I0K1
S4ua/BDL8Q8crG+sCfXPGlTDXSzgpKyiiqJ5CbIXx27BGfs95T2SFupAu/c8
9i0SEfKx4NIDMpA46i/LPekPBeGTpBm3E81uaPbc6Yx7XEZw82MXwGQaX6Ll
YaYwL50pxy0HStX9meGK6Q/oAwXVQY0dZD4ARU6tSfQSs3tGp7VFQSDKDEfN
vP16b2j5Se+IaKFY/43EbqfCDViT+6H77FTUQZLLjSSZUDO3iF0ztXWokgma
d2haoIrE+SJnB2Jyk7YR2XYk9ag9P2Oh/p48X8Z45BdIQagl1TmCJPnKnGTf
Y1VN1yyWOeJLgcTYVILPCRQ3OLmDI4mQItVu0XV2j591LAbWlxn4AyLTBtzG
EE73YwUicbs5cCbkPEPKAJTbXSifNqhpORvOuIc6DkxXGz1XwO8izrgklQVa
eenwpEwpP27PcYpjSrGBHDUO+B+Zu93/4r159TwNIqCzbIeAyLgvS3gn9E5x
Hc5SYP0SIXdSuhKUS4nuzDHLAVCUBn1HSOqOOzW6SZ+QcU16cZDZssgXofnp
XhmEpJQklp8zQ1AzJex6s9U2gPaxx1V3qGm27CTS4QG66bEUNM45bONFLJfX
xYQO4kekPdjXJ2K8Z0cGuLurSSmirnUnhLXZv37j6ab/uZGElXF/reoprJ+d
AX+pk4OHPIyZnAYBbrQso2wPXbMjU5gwkpSU4VsIKZfs63+Gdpu7IqBGkRLH
RsQRD6QUcWQc0R+3ptc9LAslJhDC1pEBJcBMQX4ojotPebMNi67D+TDE6YBn
A/f7BA57N/WhB/uip1LiUXB7g8ucZ9zB9OTrzSAodU9Lex8codYQqw3lpZ9B
uqFrdyv/bqyVSB2+ASp+xg8OqlcPLxazxhYoYNL9I1RI6+TLlaD1+LkX9fjL
kkRTr04WUJKgb4SgiH6GCecxDSQ8+zuoI/yEl9/tmx3G0jnEzihKoHtwxusq
F7VaDJYKkPPUKh91ZzyDSxO4X4lVxdYjJPCaaWu/nmecO0YxjLl4q28STD2v
410tTlFL4RNYBDmpcMEJA6gTrceitE8ml5iZcurtcoWI9rX2d6I6Jvy5228U
D6fRTqHzfp+0gBfYwXP9Itzv0QLgH++15CbdZHip32QuoXekkJOB0Jo20CP2
jksyNPEzxX2Zo6eY47FzE4EZ4XSpuLkxqX/vV/2/USCwcXcfh0RvoHiuFCi8
brQlkenQPRC3HvpkQmY5tKIwyvMd5aOQNWx74XpGykop2aWfNUN8pqNMy8dt
FFn3AediarPvf9ieYPkU/+i4dKhIo7QeKpAY6/W6Z4Kgt2DYIlx8epERCmdg
jayD2PxRq6e4ihjMezIBgItOQ7q5gddLSph4W0UxU3bqzC8jfzvVLFRYSFWa
a3f5QLavIVg7nxxjzE3Eto9dRko6pIgUYwQnjpuO35ksZAFKAtgVCSsKaAYc
G1C27uBpYW2uX9p3l0/VeO9UjtCeIuM7ip6VIZuN6aAozcMWKfNg9GwbANmU
mskQHFYNPw5yiscLwJmkaCeIdD096eNls2wecmVinCe1g9HkOWOYZoApezI+
8XWHr6SgJIDO7TWyrLy984zfFSppPhJK2ODDh+V52UpovCq7SsL9I0EVPKT2
npFyYOi6A3rHFA+j/vWbFC1QSlpc6Dnir7NAAJhpB7UxcumWIIuFW7EG9BwL
/pI8f+lb2XvF2LMhYjCDvX0HEtFN18CtzRTTMhRbs12GP5V00zoxw+qPudvg
HXoqaFvGaVRJc27tDJK7IW5T04JikdneI245LnqJ5IP5ARMkHwwStz6fIQmu
8KnlE5knW5Zm3kyGx152+N+REgZDiv2O00/Log89YhGT4Ru+XZ/PMpd/JbFH
1gRpizueDkOKxKhp6b5q4JfVPBq/1uop20aWcMORbEfog0b/g4KOIhWwEXuw
I+ARBkcHagkdsyERySJw/oqwY2EM630ysR3A/vl+7sbFvHgjyWA/Ncv+iJvi
RM4BhlQH8qwRL1IwDItXTHCoSDPeTBU2oITh/KiXM2oAqj3iIwrZ+RPyR+sj
drVq/e4rahP8S1jF4fpA+IxKTjFRp5v2/HA9EwDE/ST8fN2vQ87gci20LAVe
TzbHMXavxRoXAhKdAMj75vVtjk5qhzhNUCol3MhKswfuXs6BENzckcWB2eYN
1vssBONjba5FedRsfBTmxRZ7p2DrE65CyWyn4g7fuGdjrl9F/uu7GPdE/pHE
yP5YFLMRSIibR9KOx+dB1SABba8FFxsLmj0mmJJAThakdxbAl815KDdxnbRk
zNvLcDPL3enVURKY96iQpXqV6S8P+rKk6dhXUQ9qNxh+exQox9ce253/BVUb
oZTTcm7oGyBPFDciiTm/k49kmuL8gRNlsZzmHp9xAzLFPi6RBeUOfjww5D5v
1dS/wDDSSk3deMsub2TmTRzLjnipb95JtpK/FKpj+f1cpBKeXQxwCKLB1yu5
/d3m2DQZlhwRcjigQSRZV3EPlFqu8PTdydY/vqHDRRzpunTykFWdm6BM0aC/
alD9rpbNHjH0qjPD3pdeQ+prX0FevpVYKlOpEe/sNdwTJk18tLzncq7V+hgn
ISu+i2Hd3swcVFmDTC/9fP1aomTEUuSKb/Sdm6jG6iVnrLOZOU0K1A07ByIz
qkpK2rBLeV9sPQx6sTrWWdrldSIC6dQpSauqvPyJaX8+VDn425K83qVl/qd2
hgg9+peGgT0aOFgb6/QzpPE46Oc9PiiqBdNZ4c8ENgKmqonmoJ2GsGz4HSDu
7XRbQbh08eYf3c261fDcnUT80HJ+jcgmiqQrZorbnccjittSjFHpZhDDGYc1
mZ7NtVoz5Bl3ea4DR4tyh9m79I16lk2Ll/i/qbQoGAx5tRoiirIft51cpBYy
hbPvYiiV+rUmplUO6n8WUbAr1DOCFHL0DoSCpLuq/iQphL+U9hmrXg5W4IZ6
1kZmsufb1qWq8I9+xPq6w87eEPEUM43Fe3WC05erYXpBK8CgRU2j5GG8uRk2
DwE6MxoGbTobaOrAm7RDbMUClqtq2IskBRuBDUIB90+pCSnPP4WKmOPQ5/Sr
stpAFGr7A76vtSAvR29y4qIeKohTTfcR0f68RVbZ1Zgb0f5NR7qeJ0ouLp48
fkSxtMBnZnyrKZWPUzqBC7bYrFNbCEOBFsaVnPe7HFlOmx4ONxMu019nqzmy
T7x2a5GjECltjlxYhIntI2VsiHDYtCgsObcGlkcxE+NMIGQ1Tclav4Wharru
aQrfp4MrEvTZYJogzlu3wcgRUacuRN4d4klOJpelOvnIoKBd0+Uha7aKrnNN
34lxJqLIv0q9Fvzx5N8/kfu3IyJ0Hm3BC1M0zyDxL203zGKtZtK+volfFc40
5606x/kEg+aibo6qq61c4C+GmYrWKMP3E4lk7d6Of8x0EV2VgB7Be/ohF8yF
G+6T9s9L15JjFHnNeF1mPtgUlgbXuJC4zXaGDTuqmPSFjgxAvzF5l42xeDbd
KiWiL/M5996bpivKsrmB3m5wo0mDIF8Nr6QqbN1lkkl7q8vr42MxLAcs7BVM
zROX5pd56xUN8n6VoKVUaXolEWV6Sqpd4DTMqHSVrLmoN5zJCd5gKW59y8/L
1YpZNC/FBMF/dGHimFWTnVD9q6o0FxaurqFE+rQu+6Akq4DZHPHBRzE8foj9
YYEI4XijdP2uUnWctbNnh50wB7JJ1GMG4aMyMKRjoBE3kORrEL9BSmrNMEEP
LA7+yPW7gsy6H8SyoY8rGDUcZsy3ZpCiOp2Uojvb5liqRU+6L8rY0VrV+FI2
msKB/6Hx9XhimkXpd90dy0v9W54csgl79m27rM9W8ZJpOtutXbvESRHgcV3M
iwMV2C62Rh4tMeYqfzyYZvWpmlfKaVLIPyHmEFW40eIi2YinRpfb3YUE618M
MVvCoLg7gNkjODlYWNveqTxMhMfqZlDWEiKBMS23n7dK7C0m1rFY5DfkPK7K
SEE/J2KgfPiPVatkdja8fSuTEzbmfSpnV2aBgPQ6yrw6/e+wZuLzh2S5qzrt
jIMitimZ5mV/VW8cv/WMz1ym2Rled+C6rXf7yNEUhMxWivIIXTXO+j5GDLh/
5LnWMEZrFbGAkXWVEmim5FnnVQuvIzTuO0yUE5MB6QGcu/LHBmuX9fabNG8x
PuKX0AnfaEJGxfONHN9DoaAF+xOv9/afbnGTVMCfBJM7xUubtV79tcXYP3eD
HEkY3zL844GV2uJIMuwUDdFOsPTb7dA8Z9+5Q/9XAie+2zrLA6/B9sb/X7vP
cQAZenZViGoOJwM0oTziUk0GfXDlRpSi0kbRgAVTbWOnWQ2XdQTDEX4kv0K0
2bOFk5FxcR9BFMecfqnez+rKd/seXYw/bBR6/YWiq+RzvJFQzTEeuZkCPRwc
GzO4JXQqdG/CXA4wkwkexizNuQGc+W6AlnU4LtbcCmU4vhautLLkhsbZRoxR
y8K8esJyf+eLo5TtKRRo1IJliXhYLMm6NYn7sBMZP1XFZr0WdfFIWT4sCajp
F0gEqXIQTOpebGOeoO8ID9TzDTTVp3jTkUZ5PJU/lq0ri17M0TfK3liZYYYm
SkvLcNM1Bh7Hq68ueB48mv0k1faAzW06Tg2dHaMZmiCtMHIJQkUF62PNoV0W
6OsScKsWBM2rjBgt8N3Z462/ldFTrSVOi7Zg/21FnHeyDIGB1cjcFiDEVXR9
sYUp3ZScOXUxeRVUCajJ9RoT4hdvYhrY/JO7k64qVoyi/TVWkHlUybo8u9V5
4MOa1yJY/5fUwzKigoroY1Q4HcLLjsgfvEUkq4nlC9p7vHvHOzV5VuJwvmXK
1cULsgqMqVC+fdBQDXRva+k/c+8egFyBsPHCfnQ985P85p1b5MTgwt/l69va
5ik4QaabQlWUBoESoqpS3QVx0jDBxf/wvVOpMaszK4xksN6tVWO4D3xy4tUG
RKjMHE9NdTou7JuqUi7CRcM7c5KXiosqm3luBfmCjACZ8IpAyAtrkZeSD1fB
UCga8I27HVHK7IDfz/29fk86FnswFU2SrpAm7cykmmKe58UiqQfSXQ1Viher
e7TjJy9ycd1OLHmSKK0z99wvJ6VBISsSFHvy1lvFap4+ywtn9EV1NXb6+iJe
QeZ82A7QvjEg6edBUVPbF+5wGKG7crGRYP+sziBlfelM7tkViXzVeRfq1+1F
t9AfBAtjBQDtf3OXhTUEnI53X3WETnlI9TEqOKpPO2s/zs1ueLLOh8Fahi4C
hEf1Kvl3+76WgVPd/8rmVgsxEdtJgBRofHiXYKTANWCrvcxkyfSCNUhntvUD
4xkCyhQBzDOj/if/fTKSpeM+Bf5c6B8A0QIGebWMfJ/Gsx462U8MDQFsxPUs
w/KxIqPr3zGYYq0bq5UNVgz+CK7XFiPKcabPTpGH1PGdbhlpDtcrYTNCtLvC
LsLKyj/Mp3TIKiPukTjtzEwTTNBQ9nHMjJvUF1IqlLD1S6OGwKk6oZsuTaSc
PdbHFWZ/u+/qtKKY8QCdMuYCj5XZ2DRRikHo/RbZ70Fq62lAweaNXcowOZXS
Z2NGE84/M4u6fBJgTosolRXtEwKo4+UWu7OiKHSwvMua7IxYysCBzUlVAejj
5oU8zYatN8dY1/kSTwCZL5MPbGsxToewBB3qiHj82rTGqtKVQOTlqUcWyV5X
3ltFf7jel3qtHVt5IWwllgPnIRNC+7Pxrl+d3mPLuCltYL0+uScj6TWNEPoS
QpS6/9YogF6Fdqs3Dce5QKNKp6+ATw1zVNUI1UT/g6LCHRAxJ6z8qiPZUJmL
k+i1iTCfojTHk+yhOj0yd15paAlkbIoKNdn2HbyVMXW/FAsR2Ee/6VCSLkeH
CEhIzihBBB3pY3TtzpYeWANgpwH+jz3vvGNBLSKwp9ajgeU1Jrc2uSEcU2cd
GQhONhxWVNu+rCNRRva1OR+JELA0A6f2i40MoWaprBdt1nXqsOlJDBveDFnD
TbKKbO5/bkL6l0FimywbizT7l8KQEO1wIs5oslB5GjW757/13xfhwyXg40Vq
ngom89n/7NoZUyza8dPxO2w/kVfIq7Kor7KCwZtbUpWvxEiRLMxfO0zdTrfY
Fe6eI70G4OajUVwkX6nIP8s12JmbPQ4xyS8YK0BfP8VZvOoqBQbYCUKKIXxr
YeeixxMNUSaGCTErtRfxLioNNHk+YZahcSoLpiZAda5iEUNYJy+/2wQzxH65
tHbFgwUCnyzMm23nPFLdUj5oAGOTQcVjmCjNYBYopH4/vaTQQ1AlFeBIJT4t
dBcjz4AUMNBt0xaIC8roN9CEE5bRBq/qcp6KcJSJM393ooIPSJ7uGzQIf89P
llgRMNFvyfv8EgEbhVFzVQY1wAafNWeFW3KYLLEb5j0v/bvT64zbrTNzDex/
/wUfIO/XNGER5AIsQ/mq/mbk8ZDe5ep/bjeD5Jyf9xr8bwpayB46vlLe16yK
oOPjs2xCj4Qt/rTxCGwCHtT0CTqVSnj9Q5MGEiq3zeUqetLHJImzgt46wXl+
lhUg/7cp299RfPpm2j2E8Ti2AJVcuzdUDROsJF0ud0EEuO+FeUQL9mL3ClUt
UenY7l4c1aIGmFZS1ZqC1/bMX90hrgVXlKLB0rnsA1IONHVMBxOC3+Ov8IFu
LH2eUC/6hQLcreT9pQU9W+88HUPk6fW3HKMD5lFdSFZZ921AZlPpsxer1jFl
ceYBmRCi+RqSRzfVvbr5vTrNDlSEKOK0QgbOy8myR2exx25iGQXuj39tgjqY
JRLcnzkxugYWBbNKV/MjtJTSH/lf+z5psRrpxoxV96u9B5cpHG6unLHADBzS
fOUViBZA/632dPGmKqe6UIwMbzaRFKywVqgWEs/jY9YTpcdJbFNngR1YI3RN
vBaKLu4ylepkPxiVqrl5kdKHvRgniruIoRJC7dcdlW/00p6fedSRM/zcPGnK
/opubiAGKfDRkGemWBPXZ4PQeEVXYsJG/CdTSYIv3L7UzhzS8ko6oxTL6LQk
kunDBx4BgI+CwMmTemJaPlpOJUt1A6IMNMgMtBizNGTDOYWfGrblHF92PQ35
dV2ViNv8Nch3djx9oSp5BQvFi0zKo1gZif7iqZlntPQVAc4aCUVhydP9dm1g
zXUp11gMHmJiVmTzxxYVLcfXNVqhlTpUfUV4vGaS6oHCbaC7mr1FV+wA9d4b
5yEGpBO+O+37jnN5oukmQygR+c4GBgmDhXj4s+ZZdYX6Ki0xFidUgtWtpa+9
4DsGMJj04J+9HDKNbOciuCqq0vIfgeYkhVNjVebuX1hD/muPgSAeNzGbf+1J
KJa1nMBmxEFRexVd0pHA+x2kK0RYlw1C47FUvbzmZ8CztLGPHMiG+LjWr1Lw
DRxqbXAIHcVEDfccO+02m0uBetCYGu6Kaqbbofq0iOoGBSFMl2CXGVltY7xG
niPReIAzEZH7wB025K+R4qoOHXi+BCWsmIPgEZd+Yz9Vdt3o4V498hWN9ugc
Y0sE12cB4hZSybQO8YLE7p0xLcVUiFtLcXBnPtEggn2So/iAm3gvcgRgRGV8
ZWz5GjzFzPPgpECssRYo6J3ekn+ZLZHp5Qw7C9n7804m+Tl2arToBiVdVg1c
cFIr+DwXqRKBD5g8KKo7FekwcZzAlUSg852dE4TewWneGol9ppMIoLaIHY2V
pscovRVq3mr5r8B5FMu0qNXveGRAj6JQ0GPLtLHS9IJu+5u5eAV1O+Q9vj2u
Rs42emCniiTEfBKcHNu6Zj1TFUOAj2rvgxuwsB6/UoG3CZoyULFBMnfxBxaS
an3HbhJn9CYUjN8p03etESx1b8TZtFEaWvWnxRo37rgz9jx6wJB0yBEmcVFJ
neGLRB2HIvE1s0C8l9yN8pJGkBmHF90S2TAruXhQFBOm3uTFxHnlE2jrWAE4
hBe65lEnMGw962SRft8e2JdhunToz+GC7/x6ImzjL6EHKXSdyf5uZW5L1YZo
fkgmygtxj7yDPAF+pV05sSdI6pX9PUE0eAkM3c4gQREs/BY1AVGZA9dsbtXI
lMuCNCcJzLMauZmXzuUUdp7ivGQqlZOJLtNoCXM7tN/lXQlOz+VynalnubzT
BU0xRB00lQzoXY//3DhFNAvdWpFjSRfQQqZpChTftl+PJqsfvag4+helCE0+
M3f0zAhByzWt5OY1lkRbXjtHBOqd6mL0AiPf1w8F8kfLFOiF+uE4deNSM3zm
0hdv9+g3tdOWPybN9d6Xf+gLhGBx4ghAJG4hXyLBkYwV+5U/EGQ42ZzJUEOn
BMzx4cz7WmE9CLbwYkzmUmtuF35Ls5048MhNCozwK2TTOsu5aZ/UtKNSz8Hw
/NEci0aCXL7rxcHpk9KKxc/QYyGuOLuDTGbF4NJaDr+ppG1fuGlBaLYTys2y
ESWOaPgODBJ/CKMVw4zQcenr+O5F9zRekYkPKqXPOc16LzqPkJ/lhvrEm4SF
5FczXN9oFFh64zLPGA7tYe73JBbBdA7XlCXGqH/w0vRrFYhCraheNGRuxv0l
G7HpFZrzkg0TL9v2xGk2C56xDWjS0LV+fOdtcryfB57DZVbVsllPQeSN/LMD
8tL7QXfavo07pMwyH/d3ZmMW1jHZ6PUhP7PkC6SyAwJaSyG4JhJS8iqIqa/k
enK43/xP3mj8vyiLmODVU/8Z8ipCuEhkbnLJgqsiZGS4y1nI5b7JRCdwtF5K
1KmflWqm5RjsjZcVqvllm6pLVA02Nx2VutIXxDLeWQOXPBDtY7FEv79ewxci
AIVi7i25WrxLvStAfKxEQpVC9KKKCvbRHo9RZKxPdirpEoqnSgTuqN72mu+W
BYBdDMWW+65XZzj9ZD9izFDLWqlIGlFmEulGhkfT62Pnh/XMoYGqV1CFlXpy
ggJoWCz3hKkKHceq6aEMoXAYryRJ/DyIhHtc7GPxlh4KOxzO8rroKngc3h6j
okPbpn3vUpDHnzmaZwS03ZYUFHX9lnpFfYbufw3ryztbdQrLiB6oM6qNx4QJ
T1F+HUFaA/U13tD6tMp3oYTHE+QhhN9x1sqdi1OuWdKVHIcpULzHUAP3mW5j
nh21NZ0klQEhTouWWso+L3OUdE2GJO4HYKGXyfkXvzO0cdnc/K4IJVEiv3TH
45YeaQO1Oz12D4fu0mj81G5XzGUJyNnlkZngSI1FBN8/EO3TJ62J2rgq0wAO
gPkKh0nU/lWhlI2Uy5MxeXmT4Z+xNzbVLjASpcl3yW5lpql+cSypWWO0iRFb
GwaK2PoEjYhuZUA07qkPrdpxqeVQec/XCEwfiPD2rj+0uYEx3LYLU44kZVfv
cRrxDVriCy90Az2/knf+C+rErGJHtUGlIUC7FlaunALWz/v61+ZcLyj7+YHZ
DfOGBUbL/LY+fRJZPXel6ZrrT7b5b03pzVSckFPEaLA9+JAkG3QOH0Mnq9d1
GtyhWqI3MgupSh1ynKi9R/PsW2SPN6z0JJfmsRqW2BpnvTmWvG13+Xn7UVai
TGIa0e/qTOHXU71d6oOUv2Aw+hJT6SkOhXLHlW73JC44pjTblczfMse7K57U
533z89Kf+52VHSkE/+fAvmPrc/yF4utJBos0JPiEEbgFv4XHmnxK/igQY6Hk
zB1CReopwIe0bp8BhZ3XuQRywUIzOHpyR9/0+JUNJ9/JzA+r4ivq64XBwQxs
ENBK4//FO9Hh08VMp9US56hAV+IsZgVl8Dk9wJ7x2OCUm13PSSZnSbG088TG
jEeZW7JOrqJUN/DHo7pRE/NXT8nfQb6Nlsx0GSvXYyYZZjxgxhJbSm8tiIx4
+HxqIOWBqQtRAgH3TV+U2ZXl/mZF0WirRK7jGRhrCQwouVnK/8zO0DQfApdm
ZHB9Qj111rOMdUBUh3duqCBbzJwHAgJ5LJt4mkrQdtCs3tWL278/iQUlTJnu
DQIEFKnGXNTldO0N9HJ4x3+owQf1/rfVFP5mJDuyZknbLHStNOvsVb1hEe/3
HSVyhHHws91v+o/XkoLhwf1gvv1/aYqJrNsVWtQh2usdbB0IdldZCr3l0udf
BeUv4++fm2Tu9wbksFKTM8jKU7zQHOcuGfgbNkiBU22lH5FU6jvwKW13ZVXU
ZDb9TEdyx28G5Exm/YKLvXeSD98Dhgjs/nklNDf4JSeWLdoxulKPHs32UfrE
EK6+0s1+2+SYVG7EtCsERu93IvRszEeyuKIeRvqIHZPzAIp6m5JIMW1RRvoS
UVjqONuSQ7fEwA6R0bV2TQftEPs0iusoShsnK074lx4iciNllWSh3ezSaoH8
ekrBlW5nbgBg9UUtfb1+gUFWm3mdZnp0WLSPtnm3XXIg403d6aeKWe8PXV2B
CmBTILzw3CeYi/ZZ3Pte0MpM8aw25CGImMv8COTVQUZLnhwwqnMdxXChdALA
PLL151PhvE67rX+CdCdB5F9v7fo7nxeXZ5HnD95Cu76qewAbezAbKk3ZPwJU
qFbMzXmKAcZ23Sm/5N2nZ43nHWe0xWiYtZYgcOjnBXQRe/VsNBhu0myrtWRT
zLTGxXryyIi3DpTd21nJ3XIjeSvLO8Js4MO6uwTCnixjl3Pz50KtXU4BFMw2
QfWWMjL5uWDCGrJA13hIX0J+xlmmP2Rwv3HjOD1MfBMlp1pWBg9K0d85FQYe
UgJpBVGIss+QHvKxb1wJb9763F49CKexNDsPN8LIy5Ww6qhlR3MWR1K/ni0+
ZSyULvqVPPNKnUtV5sJvPi6bmm9cBKasFdQ7UolBoOY0MhtPY3Tp9C4TAbFc
/zWneToCfUdnHqZY+k9hoV0P8gMBFoGde596PI228ZtD7Kjm/V47oAS2dGQO
c+H2UFUTDBdq0RXRm3rldNK3Sud9yZ8f7JtLdd5QGDQbf3vCZR9zJUdxxPwc
xk/RB3JOrfUPmxgOZjW01E4s0l+VeL/B4F3kRaia69t8Kdsur2cjCRGu/mf9
EwQ6uwYFBeEVQmEuFplSU5HvxYObGPU50L3RR/Km8sGXtnOVHmS099v73b6H
wMqcgvTkq2UmhaCaQq7qVdS771WViHeoosUS4jscEUmJgZH0FyrxvXQFQ0E9
Mb/Up2vQkjN1CU52e+C8h64D/UJUHxT6r9EnpW1CXGcmONeYYTRwQT1oKXIb
Ol9FkmI5+mXo03/7iXBVQSlEN7yXMRyaX4AaX2SVVMFpzob+8ufdgLSbZ6th
so3LTofytRA9JY7T+Y7uKeGl6lEQ95KZIIj1lZW2EpHWD3VL57imk5HAO0ZM
ikAHgCfNdRFbhuHyPKfNuqwesckkCVE9t8/cd0QGsz2b5VqVt20Br7EGUq8y
7pXBcow3EPLIpzNBLxsQyuWV+Kpvox+Aa7ERH7Xr4lIZUk9jkEauQt/Gqq09
li85F9BvW7oPnsqc7QC1R0njL0wS5A8pso8Pel5uFn9+0r8/9N9PVNpXaW/C
RxufbsgVLGhp+jFLbySg3Ah/GT3K4UYcEMahF1IGzlmlRU48fbdhZ+YQBch1
zz/x6gg2JQy3Pn8oNHJLXrZs+ZjJ5B0ZBm/tg3ZtdWpEYycJ/t3l/pBVxEum
vRFbhhnuDzZ5ltEvUADKjmDbAKSYBez4mjsouQo0HgG75K7/Ihs/CMD7gBpR
j3n+qWObNSe/lZ05L51oTe3r3CT4pN9ewP7mihNFxAsXQmwinyAZvhuwH8RS
5CTBYvsgUFOMpGnrpN3v/xN/db2BGUpvBXX6wFI3fkf7qn+/xfoq4hjnSbcY
4PCWwg9YUc1MrtSab6FIwrdfQ+PUEodvU3wc8laF1vyrJdmHw5giJMV/4zlJ
VHxjdFaTSVOiaDJYAPg0DNrzxluMMGtjYN+Jz/MAbbZl6ROcbbsF64xflS22
UN20UdMK/HptP7JqgG9E80zdeTtp+nLNe/4zYWPGen/pRNE6Jfzuk0fQZsFB
b69QDLYp27DO1oXAphRskCzlIT7dOXms508EFyDICLio85T3aLGsmcK7oNc8
+poxvksKIbV0PHBnH4H1l572EwugCnkuVRLbRnROxFGGVzot4Z7bgXfX1QFp
/P6/vrevdQvf8Oteox4gleDZTUX6I3qiBnpQD4sI+wlV2AH9due08XDB6r1J
YN2fRN3JR3opK2aFTTno1WfFtUodojaI2YK4GjqdEpNpNWPuNt44V154keBq
RdZ41091tgHlqYGPR/rEnz56fvzJlwhBsI8Fqlc+kRM8mLNJ5MhnKajTSrUK
/Y/gvbPgjogTiMHQnAeE9bH/VspDETxpwszWr9Xbu+xuGm5agnglsjlsY/sM
LIXUxXpX0QtkNBZTQayDuqwjsMEna0uFIrGoLqAzM7xmT5E6DsUhGsyFAZhs
Bopk1tekvviJK4QmsqnBzIJ9IsSkawSD9X/H8uZQXxK1uUt9pP+PuXdnybyC
gFllZPWQMM5npdxEavM5osLAnBh7SMY/D/vO8q7zIGT05ZCPBNTn4G1id9er
M9W9f9Xm0vXVB1EbQr+M60mxSxzR2ArbFm1nI3RrD0qr6N6bsLd5zneyjcLU
ffGQYOIbDDnu5hrzt6G1l1c8DrmNyX7yJZnmkXn9v0fD/1CEMQbApNbqIKPO
h/XFfm0n83KQzel/25htRK3nbcvQm+mm8aNM4txmwmrtSlcZcdsGz/feE+Cb
Mwa0SDaob06C7y7IVBJcReVlIk8hmmhi9oMv6sO6sro71VAuEgXudPTixGR/
o77haMCWEtMO5t3xrTi/WCyN0hTKuyM1DSwyhPpr6MXTwRC2mbvRKR8i+Htx
41yNF1F3PTXE9EmPAzcgCzS52LwE7+pfC1f3Le6Hgj2zDci9QIjPanexTIlk
BdWzBp6dESyGWDSE/fKkGo4+fGqu3d3QdYIQrCYL19e2kyBLpBDCO9kDE0cf
m+maupW9ZCGb2LqpUbEZL4jxu+TP37ucXh9oX63pdaPpCRjG8yT5/FcWWxU0
ZOR9DFdYe0uC7g1siinhOIfS/ccXu3FP+BqeUqbOP+utFPcSmYJgZr8lKyRl
jsvTBcDSi1LudsreGrWcz6fQkuZXlpNUcZJ9uk3Bny6uf/J3zv2zAuK+DwP7
7mo0oZKCp8TIj7axRaRWLOUf464NU4+WWzym5EEv988crTkE+7w3J3GNSOuu
I1vByl4KQkvAtf22tFI3UenikWIj3VT82zDW0PemslMWUQAby/YtbYNtvDnk
ttrFW3UPpWJsSG+iw7yhLqLf3Flg1RNgDjyj1IYLMEXbWNqhPjjg6Uva4Csw
l7dYJ/hVQCm1l6xDLQBhUbsPpr3YMnUa4CfO7OsqTfZl0TYpVlLmq04Vhzb0
kAPGRU9L904n/ENbQ1ADTt1lVG2diMjhGUDyatKst5igdYfR6wu+plWGFh+J
9uG1nL0yQihLwZWvVWzrB2jNKO8YRgAZIqudvsnyhayVVhqwzK5zfI2eNgc5
PdbxnUnHn6B3Yw4Td0DY9Yiqv0086QHjlwTaxrLzZE3c4hp6+E5RmTemMZe7
X2rrVwyu/CZgVtwY2OEnMhH3Txy7FCoFEnXzV8p2oEcwXDautQKzvqrbVGdc
ZuSQkEkuCwOcppETTEpaovBb4nfX/parMWJJDC2Uj9gdCDcO4ww6J1W9Curo
6YU70TZemu1gtbuVn5mcD7g3A7l/E1L6H2Yl0VEmtaUo3pk5S4aP0H4h2uti
089C7HyJ3oOrKvP3LztfIAJmViJa1Sjgm1yN0MkSFO4PbqxSJ9RmDRCIXbsO
FYx8l+kUeGXTKNpDoedmUKQcVh7+9JHj9f70/Q3SVcLKcBOqkCiHfOzT0IWl
kyzYsBx2ShuP9zvVwBqCXnK+21W/bGgP5gnmw1WQ9zFRXQThV++M9tp2WaIa
1yPxJKkrCbhBglJvSX86NzX0D/Yx6KSjzO9lcSfuqZgNYyv6qzsFpBuEWrbm
Bt9VexBkQgupR3Ol3DrxXdz7iYmO5Xmn+rvDgmSgaustlUzPE5T8ASFnLApl
hpWuAZ5WicwrWMp5g7dBbDz9Ur0BVEVVpyEkuanO08TIBPCmXHjQXYuExp1o
zZF3zRnmrgmZwUXNlApk8LDO4qrRGgAV9dCprYZ5kNh7Q8it1m+o+dj6B2H+
/V9HKy5zWcjPxyPbZHRt26cQjr2WcYhF9cpbjktpVN57g9WlLJxojCxUZY8L
qhvUqDdf+WYuk4uWHMc+Zt4ul6IG7rKaj4BnAYYBuLxD1h8TIZnyM3mSefal
Ug/UhmlpOQdgEOZaIrkgd99hYD60mFDE5lMf2oFCSt7SqNuQ5yi+EMYewCKO
bXeVo3OBlJVuwpA1t6pDViqs6d5jKN6flSiyCYAmeKiN9hMhyiU/q27bx5Wn
9gGL/KS5eU+9XV8ala5KpKdQ1oZi+OwFR3wX8RaoJBkY6+XBfzoVQS76mtU6
uu8oc0e38geSv/oaf+0pzh1dNv2Cvj5ZKGv+EWQWVVUcorrCNMic02ai5E6o
Gly1IrUtW3hk38IryMnfsITl5aUyMwzXkWB4VDroTdRN0UeAvqe8x8yrehwa
sgaphHTrRjpr8mRrTuW2uiq0sMDLsfCMBXYbopSjkt/yR5c+9P0Eha+kqpT7
eERkWhW/rQ6bDqgbf0bG+RIms8MXLDYKibPmQ9RFDjviYs5m7+l53W58GigH
HkN5uTV0i65IpOb1RbBi/mv38il4EY2amlrrMaNEMAL89/tgloBPsEFUaBNZ
/8sUU3lJM+RMiZ34tQuUEH8LhlwIOVI60Hsok2UiS905jniMT1++eY9zqlmV
NqnDedZ6kKCT2TqOSuuen1WXS307VRRTLKbI29VKAQlF3GGB+7sCnxtugmDd
wN5pWRi7h5czQytlkfLQhJgrMQwCDRYeVK8ND04NfXnHJ1cqtQ57MfRY1LQd
MQl3fnIWhPxsVNcYh+wOg9j2vwl5WJbJ/wGGEBzFGw/9mo3J61JeArv4JHIp
QftKwtU5+9d2Wi5i7cF4rB8g6hVsYz1zlUkTznfOshMegg04wOQkDOtNJ1II
qRVDRyXX9FMcHi0OWPU8kQOS4yDCFYsEiIz54qq7vn1+TzNSlXDFceDY+Say
1KdUCCd6/J3KKiDhjV9Pk/YYkZNM7qVoFcOa+DpUOrvxIVooKW/ZRG9lX/xO
D5xtlBNun+1wTUeDSOXOw6QRDTsS2Z8BQhMN5+MuMkc0FLPCxEsNPgsmJvYo
OR7eRtkwkLMb63uPMe5fyZ/gKl9Zm+g6Va772PPClykzBzWcPGnEgKkcEhv2
yCbr25qZ6biY47HGZYfAqZPBaVZKoA5NqCptI75YrU3PzH5LSP+r9Qy3o4jJ
g9jp+UWp1lQc6bFFRb9wpdiUIxGAQJw4Cc3PBzH2GA+/LMpu7avQQTXiCnYD
dpzwJZcyKvGb+ZQzrRsxfiHlLNXcjyQaXekXizdlp0v9yDt1c5UI9tLivSqM
6vwEp8EbFaC6ZwustRvzB72yQmtjk6R57REk4h6eFPsbeKEHephgWfCA7r13
HmZLbnyUSU7ic7NexV3JO+6CLqOVlV8iph2SsnJY4tQIMDQU45tfQmsktqnc
8URf1S72nwiR7AvcKbt+GtvPjYR9ykNaYtazHfp5d4JBJij96O2KiHrrNrje
nmB6znrpGbjCAHscuip1jS5HjueEkAclyUjYAS+XqCQGPJevsz3qEn7lujiO
RH3WrfFnlXubAeBCRRe0Obv/scyuIWW665kiJshszTzYpPs77qPZZMzGLnVy
eW5j6ZoqAN1s5taPsE04uvZS87GGB1ESqWgzbn3U5GMVQ8eopM+MUEkKZKbC
v9Dus2m3OfyEoCa3v4WdUeETbNya6C2U5T1T2AOM05McGuFq5JiWpvtXRfRX
/m8kKyg2PtuZ5SOBtHGlq4W5xFmCnL/JUHMG1KvXJcryrFt0vgxAElNldr64
1L1da4LMlZids8Tkzl6yD1x1XkumtgxVUMX8EHHEAKVemoOR5YJx9iHVyC9g
wca33Ds3GqjKRCJ+hWkjlY2nzWYUe8qVsIYOO5wMzUz5WXqJq8qMvToefqyS
lOuthny8GN/46vV+9uZ1JICKq0nyeitzg8gKTAmQUA84iww7AFv6MRRRD4eY
w7r5isr68tpD+dKNYjihp6WR+I/tVxIldtfRM3dME4zmHyKSMgqLDgm0WdAY
1k8rutL0FA+FEcC/fbmPWB85sE9fbRfDvULFGAuUZKmz0yAi/+kmiTcPnlrf
vPaj2GuphaSvKyiLentseMQgmLypxou++LzhGwbT9O/ianWqVr4ThNKG95IX
hyfcA6JcI5CLnNe/QbIuEl+OnhkmJfpsVWKzfmLK2UWVAdH6HQFxT+qYzXix
RoL931knk+v/KfIVJ99h/mhro+ds2ofXjn/X+vPxt6aCrMCZuzccwAVTQ2WM
dBIvu8FaROMM8tgKYK5T3muuVc3ypXRmaT4gqt9OENg+ebAfh1xL+dL9rJO4
PipZwBnF8zhmpnrz1uZtCiDAAvyozBJzEnFULPz/n9lFhH4OpAlfC3d/fl1z
QvTKSi/DnIsf6ZjyZYjaZe9pKiLxwAP0Kl84T34dpqcoWmWFH8hUpmD2RvSp
uUyCmegooDxYqCV8ZdRrvYySdtZ/V5poxX+xMu1CWA9x3uuP8ezeCUD55m+I
eHW/TBN3abAC84EjZC9JOhWyL4Kj1bfOvq05Ruzj1xcHJon4FhNlJ2qpVu2T
ljhdNZkhqfobl9ClFQTjqGh2p/aJJ+tjx9YDTmPsWxS201AtENServmTpOSC
ZssTtYc03YBlboy7BEt0dat41xxx5lznCK1k+W6u8HZofeybujtE6qGKFgwt
6Lw8CanWXOxhq1ZFWduKNYilqYNF2WW78lqDB/zpU6wk8RofJWxbYxmyDipa
pSzG88iSMNQcgUdxgWNC8QBO5cExjW+JQZSG5uCXXfMD6K50E5Tkjzstd+DT
9eOvEuV/N5EKAIXxxvVYPkUdXtazpYnZIe4Cz+8mPLOYGfql6zZahmWlr3U7
TLtBERcKPYH+3Y9AZtMAfoqtkVdeDVXbCZ25bG4J+pubNlouM2UlsH2Ojsia
Pn+51/jYwYNMiLFse2ePFHoqmohnYkDFrUWh/49m6lAFZND2TK8rGJG5LYZR
UeuOTw6dQV3eSeNJAZ7HBtKxN6CcNobFBmpckKPllG277FAiNbMDdVmQHeEP
V6SFHI1le5uum122MkFMq3QanKzrcLDrOiq2njEBnuQVc3bOTuoRIL3vTCCq
NXdbgiD9Szx7pEGs4ouPf5Dsg5V1lnDgyzBMDW5fQwnDlbdkXLS/0VeLOr5p
wD+S+ugwfXn0peQB6KIme9J0v1nHN5bg639t9X3gwq5jYvv02ysc6M7/dyoT
0eqa3Xkm6s/u5uRG1WPNoFsCCh72/Sj+AqvtYsXCBVSFTnx9ys/HTaaNEGXR
wiMkwmrNNKEQ/gfuJKfd+IlkNYdflWMjH0RRZ5Q63zfULj7i2j+OmWPtEiPv
69aya+oz5/cIf8rtsDbY7CLoTOtOkIv8+sY4SGCjU5XniafG0oO8X3kocZn9
V0IcL3PedOIH2+zP8HGhnTs5HYZP3mBMn3RZRHyZnfb9CHDlrjbbQsys3//d
A44rQ2g72+f6Ft9/hJki72Rior2NwsvQMG057NWSJooC8wUuuqMiLzfiGElt
NJv9XwkGauPF9EtqFUMMK5CgHt1CKGMImi58xRdqYaUMr18xVBGMkHtxCp8U
9jh8Zw7EIz26kQSN6M6cG/NPIR1FEwhYMmGj8tnXiK/1MqGB9v4gH87LsOk3
kAq5G+ot8D8dcH+YbGkAx8fW7+0rDDYpiuCXp5u6y+e8sI9nQfglKpGygk+B
8sELw8Yxsy40R2OuF38GETT9fBQvA4Zw2dXwiWutINw45QwwK3kgATX2QQrU
2CWMzhUqve/2z27vyQwCB+Zpewd65qL+GNUzH+3pSRuYX7a5y570AvKVKHJZ
6mzsJ22ZOmKvT4dRPrwhVjPvkq5AdtyIziEMqfTt8mnmOYP+0L7HO3EU6rrZ
rK7b7c77bxaCp5AckVMuBQUf1p4GfD3XOv3KtQi/+fuBGhUaJcWN01Vd4KH5
kGFhN1CAC98iPr6E+/csU4EEIonEi11+5+rMk1YgnHKefinUV+8H0mjAd4rl
URqsyKZgf82UAAazX+qV8op0ZnBLuepGbtkDqS1p74CgFVs7KwPuh5HoK1Ym
FzbAnSeFit6YLjxzVExEW8wNByXrhtjoSmQQlcrpByQIMnux9LxAJTfbLDag
VeH3IWhGd8k1FKh1DF94ltfzV5/4HgF2rP81uktJBKes5iCJMBgRZNdQjgyI
fmo08INWu1NciWsrULnYIUqnLniD+S4+3NiE3fg89umnexscZUOc4BucFfjS
+Z87s/Yy2Bin5jl/5Bn79RKILuFDEY/VMyoniXqYn0lDacEfkiIabPML0j8A
0Nkp8e3OUi8mpoOJQgGFErdvMgY37rCgO+f2ZZ5WOFlc2g8MR75YTMop5Kjj
hOU669sq709ouMnQp8Yf3vO0wbDEiFPKXWoStGjUmZjTem5HbqcaCBVvqNtl
a3nQqP+FxLxRzLgPskdNubSBLVk4sDobCLzbDj4T18GDhWPjmRhxKfpurxrA
77Ni1d2AoVAAh+Psok10EBpy1u6YssjGXmsoYhKaS5Dq9qZa5jtFJitjNpuC
Alf4PFsA/0C/x3IdxoerhxwQwte9WBDfyvIskgWd/J1Woip85jC+VsbjTPHY
inawCozfoes4ll6zFSuzQc/flEE5igxdV0lnqfEUu8FaZ4OEszNszViMrCg5
DVNvJNQT+8487pRCdQeBHJIAD1vHAPI5hIbZf6yd9L2TKdKlY4y0qH63krrO
E2u2mNfl4XCU2dCpB056gixHENnML8JqR57fstlenj0IOYvjR+2f3Qmuj451
P+wpMZaC8yM5YWQ59Eqvml1ET6uK8Ez7qfC6fSYSAHx7EBlP3r9cEzueo7fl
69KbRLp44WSR4bXcLAWqGQ7DJ53xj06i2nkjO2mOdwSML6uQ3lUTFY2mRvna
ozBHWWmRowj2Azg+mnnCZ6OfQVW/zIpwUnLm0OuWDZpfMyZ+vNv8tDt3X1nU
wS9G51mpi67lvEJzUQM30cYstO48/6H8UPsIyjxYBlJHVfJyfHipawk0H/zJ
deeLBPqIE3R0HpOndW3kkEkG84dwBHEvAcRPX7e1iyOfO6i/EdOC/6RpAJMW
a0Ekfznvv99Z0cWJS2qtia9BOkKN/1MuXpX1XpzqrYl68G9XBz/rS84Ir11z
G775RgfuU+MU3L+5FYN2OVk5G67ulZl4wY/BwEAAcSAOaFpRySsdUSOXXVfd
qVWr0oDy7UgFErQlARtzOfG5weqoIM/vJUbXEXEBHZ6se1PwdsAgMtdpEEeA
8NbJXXp/PiWC8pFQhiaPjWPmQBRHJm3U08MzE/QT56CwAqUHJSBoCjjOR+FZ
zcaVUDakJez70zonXi/eLbYdKtudVbYc9J36fPa2qGdAIAOtpGwHywAknnY2
UmOorYWmsPU02wKcY/IPtku/0+DN9QnCh7MmhYl9QfH5C0CbtQuy9rEjSpo/
Yxis2z7yE7Y3WOR5lKqWRE3UK7GcOoibpijdRM5fv47qLc3wjYHytOC4gFqL
bXp2HOZ3V1VH8+Uf5XB2McPvouM4RPgCEHM+8qvr3hbyOVs4UXRuD1E9z+4B
rJb97N4hEJXMUE/46NgRm156SmhOcImZtUc4xOGSfRA6qD3GWI+J4IpcyHxS
/P/TSb6OkpH7AaWE/TpNe4jHbFqlQ+HC2nfsqhvjK+yFeJI2SUCLMb6QM75h
geRXG43uZ91QF9DtIvTUfrae977CsXUs1kOeyYn/nmvPqcRj/E9bJzyPFY2S
bTK+TCHz3NwQnGdow9DFkCnRdEvlWcbUk4DbCOeI2m6S+TqPaQ0eeQQlBCEk
9J7Wc8qyOLWJs++pEfGhVX26Db2QkEpqZFuuCRtsYTKKqTWmIsNU+Ci7DyYw
BA5OXzBYbfGLt9C1Rp/aLQKtMgLhKhiXbh/Wfl1RzqK6Ecp1JEsmRiyF2A1Q
B1I27cEHV1huVVIp2qHtBOW33sRGQRoq6PT3GaCsAgFr5jC02tDJo8pHY8P0
6dRG/XdXdfhqfvEIA+KLwOIWwCwcMBF1ccXEGLlfCW7EGe65HNYyZw4hJq43
qBJbqr4bDrNNuvzCfY6fddedmECjZ/lTPPScG96VNvACGm1muYdvRrYMVdF6
IkzrgoOoxvUFsb7RgoH+zZH40EE6cCEbXTGHqAu/atsuHHLd9HkOtfryxHY6
zK2QyT0sG1xBpS2apVXdr1XJokqjVL5ZEiFS8gjkEFaZEjeEr+EWMQyWFac1
H+RCp6lcqs+t4iU24caioijdfAtd1M11VavC1T4VIlR+xsqqkldAtIr6VqXX
VcUv1J1WM2x1F+yV6RpIZ84ULVh0IQ9m/EfYhOKK20yB+kbgIYoqrwk6a0v/
Ub8rZ2LD4l9OCUlf0+U+bk91G9BpISu0w01sgiNQksYWGV+6K/s0XrF2YOxA
D9jFzVD1ytdXKwoGf/Pn/vd7Whe54JJYUQcx9wNP2ZC1qybFS055W30Hr5Wz
m0bIn2/pCOnFfv5gMbubT/gy7NGSxdGTUBhrlmjZ82vFPESKNVeSd/wkdCD8
PKyAZNhWWMKC4e4NRYDVwu1OQqlOht05cy27Xq7ihgG1e092u+SgMghOa98e
kk9K9+LKGlz1hqfNmrQRqlVTd8cc/UwquR88xIYA3bysGstnOghiKUmTLT19
ZHoWCnaJugIARAVbEVuVoJ+HpsQYmnEbc22yYvDxWgVHuXfM5UNB7rIZ1gB4
4gHuRCHwr8N0xMKg0Gx0bi24sQ0QXJLUrNc5KOM64nH/g2xncal5oKK0in4n
f2FfLV38flkWoqbpXnHN/htHFTheqvMUATIvnwKMRF91Ld4+7jd2eWUxR9/B
3H2inXT7rqPEoW9Ykys4bBDa07x0sLxTUFUgySEyNO4ity6M4vRhX+6Yu5Kj
pVapiv6kjGf1+9s5MmU4Wp3njb7MzqYSkBmwuxMeSqKMUlsHLFiqlEfZMS4W
LmZxkkggOoAERXbSiWqH1cP9PkCeKkVKixR1HO/NqRWI3IEoJkf7514nSscV
JCALDSl1SVKfnrWyb6Olh1ooaxzlo868mjYacLtyjiN5BWea15ZXkb6cAL2t
XABQq3qZYu3NYq7uY+ymIcmNOB36CpSLxndTgLzILy7efsKphxKmgd/opIG5
HD5S87W9rt68ivtMwm93zXl0JJB29YBHju89XFmITIaoZQeE76keo2Ph95y/
TbCOlmIpYqsOywUlEb28rR/cSvE+j2W6yrDjTSzrNRJ+KIFYGTDc7oTCDxGP
6Xb9R9dMTEqIV8I8wJHLokgin79l+fW7TdCF7svXqVmOEXNOrRu+Ps6m4X+r
9j9I5KzEfbhJgNUq+HjS+VhBiKjl4X40/xH0tYaec72N8X62Eqqrmssg9az6
5cX2zrKJAJDWW/rkerapd1kKPB2PcNG5nU8W1oujX5HWp48cuO2bDQ08b5yn
7dAHV7YhKThzon9zBC5a15s023Y0y5bG3/b+1TNhWImu/F9ZyP1+ml2o/nxT
Dq/juvlaQdIdV5KowUk4FTxhkJUW4Lzp6W2GIfhdxE1DI3f+9OQnwwUezEa1
iqfBGJiz3yLtUDrguzBV6TWKrL1NHijtfHfajeKlROxlDVkqisN1biKY4GEt
U370YQFEWUJvEBLT1Hb8B3JlU5SGcxOc80jVGC/KQwZLAmom2JLYJfSgjrGf
vH9eFEOCbq7kF/LdKEkDTuHFOAkjN76pjnZ6KdyUR3w1Uv9zHP6ZPC5/anTy
LV72rroVl7rIxZXpP1s1yQtE0jjM34D58NzIDWzV+530cV0VJtLv8+4WZ+pS
YL+FC9c1QgvBKRPQ34wOjlJxUIM+8UDg4MCwBBYoRTZBUBWZRNF8Y+W3/VQ2
J8cYoYdSMPcMWcqtuKEup/orgAoUGD0L5shSyFFdHuKZJ4enIlq3IPEe2Xtt
3bg5UM/zSujkyUX3oMtCl4FaeOr0e9OOT2rL2/4gfuKTNeJROqJXgUK50JVF
KaZoBvSdRlwXIdojfYp+Q8uJHyC2VqXF04htLty7hs6yOCsiSW2+W40BZjAm
G94JsJMIfK+Pi0P+NOvPRNcm8JFhoWAF9yP2C1H/xU/xZUNsrohK5uEIITNW
Sig/EcNP7Yw30yI3uNL/dE2En5Tk8J3p9060YNZhuTt7egI72qAquOhaHttO
lc6l/i02H36XYGkdBNL7xyLeacZLJyeI1hXI9WCF2ggOBKpChw+p8Bqu9pNw
WLyuli6zviz+qYmavp+cYU/cZlWpCS5QOyG/6bKpjsVSJ95cz7BU/0R2dxUB
veeE5b0kkYUalHmCbbtwZzhBNwgsmtxM4gWj4sFIUcDemIp8f8B43VjF7lHk
/mDioBQc0N5dqjMkmi98khG6Qnt6ttsvgU6bRoSvT8OHyN/CM65MaOIyNoxU
g2YXNRca7L8YtqbP7jUJyVVfMYdAtmVrSyLlDQ3ayMf4AW/LK/hFbE20a+PT
YdBAmSBOZW1WWjvXtv0UgMoUap/cPRyS65+O6cJ2Mo3gqqiOGIKLs5pKRF/v
EqcaLkJ8A/E9dmkBpMcrsl/PhZoOCkoFRMW1kqbkNaY1LuNTaIjkwgfAOFlR
YBCI3aADx+qfrCFT/YjNAxOMVn95zSWnuFlGJXcT6hDlxK1K+TBsX6lBVjU0
pOZ8Ydt5yEQpH1YtGmxqvHdwshlgcNg7MgiS9kDowxqHu71+rtjgPrygyXb+
AXfwujI8L9Fe6txBzSWFyXlQv6ea2MHyaRjuxufPQFa3T45afGJHtw36ff8X
VhzA5VrjRBGjjdCkwAvjuqD5BjBSOcK6S32dhE1mJ0Y2ep+7GRZnIJbRPea+
oBa+b52HOElLmGq23xesX1qwBJPuojvBeDuX0KNlHoepa2TTcYFUPfmevE4C
d6Hmb5NdCvjltoOhFHwIIRLPyqVCvBWeaQyAwUv9YENKxWJoF2KaG6z02Jx3
vFAmTY1KYWpe2n9JweLZieMFqVmaYpHq5ox0Mj0ez1hfznFZAxYXU9Z+UYYL
zq8urf/fNl/km8Dhe/kCH3ymnIPa5FgU/fBgnTLaFWtvpIGkQzx58Bbc+18b
fvgPMH8IH3OUhhbuNGOA4vCfOOIIhDzJINHHFZOnuUdmx6AkIIFSv+QRGBm+
eQsWNNq3yRaLQmVBcxA3TTTVB6EnydZ444EXQNjihILDN3dSmlJiAgLEZjIN
L7gtoo7U9NkpwGj2U2vdu/eaG+lkdsSIQfLaMFgK8OhcI/cgXj8Q92wn/u2c
Y1j4uPEHTjizx/hCNEk7Ck/TeF6ibm+20q0KN3adXoqlF3oBerFFHzp75mE/
bFoLWdvJV0vaJek0PPcbmaKhkGCnzofvJ2fxWPb38M2xTtOqQnofO2gZP3rD
1ZOi+vDfe1mgEPHi5RaY+GxoUcgIpoZEKQGlN6mlUoduNn/HEZVpna0Y4EGy
hU9XIjeJUvH0P0e4y5OeCvT0LD7X7Sa3fJPwsBvPrkCG9rEI4w+esSqRUIkg
mAmhI4GLxom85/WbAxLYyoAqB1Fs6qQKJI/tUTXuqhE9egDfVCaLdk7t7KzN
NAehC+l/Q98sImZJPmpacfjrTRBG8omsuwZ3YnMbly+u3s2tusnDFAYIwaD8
WwlXI+hAYrfTnLU5B09seqYTuqF8wOXklt/9ApzpVOg2vvWSlfffg2yPZS94
iGS8isK2ajrIdhTu4VQx5OzYXKjky8oyAfNYuSxryQiE6/BVVVd6MI3YoSLK
dZFTg6GEjsQIludDTL7OAzGV0a2sLIdhRb4Z8elbiRQhvUD3AvyoktfrNzYY
XVXmEWBrBjbfOyDVIUeHTXVswe8EUrX7b1kxk65LKCfRT1ZVtyZRvQvto34S
81ZqYcZeugC/iREuqbr0x8C1F09DLOmiyH7IRyC7T2sHOV+TunYcVstdHQ5/
2B+Nn3zi6wUXspJ5Ul3aU93OOJ7xpthxRA2BgIYdZ5PpBWtURlE66YdI0Lnv
K0qWQKSYUObaP8rOgRrsbrH/U2y7ZNGO2lNuo0JIggmD6X0wPX9TWAwDKYWW
yVtosQ8ML5sLtxbbXeu7m8X+ZEUxAd1h2HIqB+gs7a4pL8cnsJrquBkDkcdi
Z8vKGq6ezJmd13mDhfESP8XzvwZ+J0zg9Lg7cz+pyqsWs3nBt1HwZPVRE8up
y1UC/qPtgfUV6ztssug5oMIB1GcvGro2oFU5pPorda1Gxh87bht16ERUvUqo
3fRu0hdKfgLOpT14YRRNIiMTlt8CSoZnBS2zRCNsHlvPFPVD3WINfKEholnH
gxVgZFjXHhuWLW3ybrDVr9DD8XnUEsFuZfsgBwsQ9VrX2jlzkWILHZFLkHnc
jqmtMFtskiWk0lIzOmRr+B8UCB8qMx+2GzzJzIpV44F1E7SIsxOEn34nU9mE
1a8kO8tVInRe0AU/EyMBhOkSn67pEbWbNb7W7O4hWANph8XrTc5fhCQUY1Gi
oDVBIb3FhtSpHcWKW94Z9MK87m1hR2qQL6aPYvoOeEC+wef2RjONxtaYS8zT
PYB96wss9ZnTjuvQzWfNDQYMRonT4KpaxeE+VYpHwzZXRDeEzSo0Ov28rDac
J445lxQpENbbG0wAdV5q0VJcslITn8hUW6z/UDEDzXId+KS/qzmqBg/l+WeD
TELOo09QK4DAB3/w8fHz8HfAhNyQx6674LBRLdDXVP6/GvSa6jZTDa0ymOqA
A/QcwDQd7X7Dg8d3sUz/o0edsp7CuzITZrDe4cAO0X7yFQeNa6poaegkBh81
XDTmZYUI3X1yLQn/Zkd8QChxS58CJ1RweUDpzjaJRS8o1hrfNByDJ2orLzNE
5kWKRYIyAutrkRRC50GsD/AyitUyRgWOl3B0Mb0OjGP71qeK0tPnaUfTd+y8
sC9mSGbdyXDqW+iMMd1ltT7o2s9xPfGcl/S2ObqnvICtWj8x+pJ5NTidJjyp
u1syoNxmbYEQy31XaQReUaY6s9k1mjHew53d8YE+BYD94E7qPLV1fbKxaY+T
36AYkYMTZ3uXX+G3c95F2eGmFy8vY1WS8uWc+l0qDRt8nY1vROVUL1LEUm3u
o/xpRPbBxt8DwQgTDsOTihYuztaQjktiOg6OleKKHm1CtcKM3u+t5QK3tyG+
kTFAN5w2Rq22sW6ECgWk4p33mCFUcaVaZLD4JNrVi9KBD8CGL8e4ZDWX+G/p
pWfrTHmrwGT4pZQcrJJ95ipV95TCSRYjBpCo10lbWFMO4a8MEsgf7EEczNto
nDGBhh6Z8LQUPRZXLVbkOnreEtU+gZ/n+j7g6hqg/hwdglFC1J0j1R8qeLpa
2k7DHUSPi221GsuqBrnkoA0LEx+70TzpHcBLYqRhUBQezV89j+coQczufJ5q
nkegAvHtDBUZUydKkPN3F01IkIK+9IQO/XyH2GEPYfDoMtdQSo2tFpCXvZR4
sGmuCory2yONmW6sRnqPwmV2prI7E/3Ly542LhWgRknbBmj/IBIQ5KU7L+bx
vu2pO7l6Qc9Bqs9veK9luqHUH9TLYP+Nm2x6AT08y6Y5sEatmzwdom8gjlWJ
esTullw291r1c9BwmMJdPC0RQ99SpuxYq/y9lKR8OcBSn5RkGWtGarRO8uBm
sFHoP20FXXMM6JvYPT8dtny9LLdc8Tc0dpuemPpxegKeUy88w4Lngcq6x9xc
Dlx1tCot/yKY92XxfBtFxaUoNIS6S+3A58i9wuPgO89zgh2qWGRRNlT3G69L
qPKJL4/gVTH2xHtwQSFe999/8mv0ERoEdbomHfiVqs51q4l/k9awpnAr3Emb
uEYpcTgwwgvsxQfsBBeniHUYKWr1Y1I8+HrKyY6jMtTvrwHd8MPyRtxcT7Cz
GVGRME7qjRdaHjsugaDSo2zcHfIo4gIfNKovmqM2bfgZX4GintDGuziqRsdw
lqfnObX+PO/qARv4LMBzZhp5CcUuhNxlEUMJ+0mvIvxUtvYNEcUCCG7QkYMF
sCJqjaSQk8pIjqhaarMfktCJIWgFohVOXgt7ec2BFI9NziAZDh6/K5FlFu0B
FIiMoxo3UDholPrvsYjlUYodyWg2NPUJAC6MQG+Wsm3GSUG9ZuQJ4VD5tzm/
WkyRrsZUo5qHiFx/6hSyv6jvlFNp7DDiv7uepfE2TPsV6CBLB13ys2CAR/gK
1AMEiZ9peQlNcfDUiMf8Q9GsNup5D99wmaHsT1fnpmRyicbryf/c1nR0wN4K
0UxgWQoOOc85DlIschloolqPlGxU3i7xKyHcQ1ZvR70CAwDCnBP7uhOulhHw
lBOqU+U1n1LEz8NSNLyJTQ5+qtTvnce8TkXkq3UgKlleXoSI2s6IJk55JKJg
UtkQOCpq5aKXhqXhK7X76KUnxaaKuk1n2P99bsehhjaKjzBvCZlaefs6QifI
gB0LOQnrTrv6nZ15w+juidpk5ob/o69ATvIM46gOWHHxyH7oUgLJtoaVjCdJ
vx2PH1cbjo2PTy8jPLtiZ5jkITc+BfstI7UhnpIfn2YUnISOOK/Jw1YXtdCk
EFCGbOGTJITqi2356YD2tJ3aW21CDx5oSMJC9OSXYETWhgGkLgFLg+UW2yKo
yMIqABHm8LfvS9ogalpiCPWBNE/Ejrm5ME/iIMs+6mEzAlvAkXp38NOZof1O
otSM6C55eBcVus8PmdK+7zbWsxy4oxK9/mTTlju4gzH325nI77TeZ8XB1OQY
Jps7yyESwc6xESm0XLskHYQrHZFxF9wL+nedfEndRtugrdR/KixNfAGPjLzL
rDr9o7dACDIHzaA9lHy1rIh6NEPO9nVWP5Izl135XxWGN9JaDfuSCeTFPONm
oXETNrTFhuMa6mWu/PParBuTEvQ07SOwvCOCQlfKZkJDMaiX4SquA6MT1PJE
lD9tRSk3HXkkKmAfMg15dHEViQQqO9DW8NItxFLN2uTC4RUf/nT783UUJLsV
Tv6tDPa/qw5ajG5P9+JdJ5mcPkBnJNTuh9sNWE/uEmY6YFLHA3GPJ/jJAWOH
gx7CPeLBjHpdq1xkK7FGWH/y9z1OgvrBJqUXazWfLLQoWr+Wpqkk2Sw/xDfN
32lGLdJxoLlgJsW7XEYe91SS2xjSGnTE218I2EEGi2VN+coogH9xnB+jH7/G
uNHU4hPrYJ9yhK0H9HwsBWP2jwybaN8bB8bWXMUiwC5WZTtg4kreaoVqOg1x
dkGR0IyxUhCuQEQYlFYYzwrS56JDBzes1Ykmlm8Ps2mBp05QFhavtZoXgrcF
jQtA2R+5otGUk/wT/2xL76DiL9nbhQ3J9v5oLeLrNN95NdnlWPwLK/RUcQb5
bR3sUt2IFbaT9/KHEKfvJdXYO2Ai5nwHAX5YY5bXFA9yGgdGn8c7uSBdEL1U
DNd5ynty18UOUbobNqJlu9DkE/4w6oXBQkc31/Jk+P74d6q9/ByiCxj24x9n
hJ4XIxlXcQ1AqlNAtcqVchLEn5OdavMx+ntpdwV3wLXy+lJk2nbympecze9p
XjcjR2VcC5H9a+6kmAevzDgy5gnMx/dweAkLiVZe5V/OOygiS+XvY+9p1aQc
pgvgXIGJWCOc+fYZ18HVadsli7NMAD7etnrnfLvbvF0E50GxB8P9waENVWtE
cpAV3O28TBflL3WcOr6SHCbR92/ga3zCzx7wr+gJFmIP64ISr3Wg+zd+F+ao
J7KpCjVcg+PmFTG2Orfn64aBkkHLnoVLnUPw2q6FocqykbbZHEeDq/KS0MNp
N4t3rRs8RXAWkSn2wRg0IhhWcfuCvEpxDsrphlmMEq9jxIAXVVDFdoT2/VH/
oONlyszyjx0pRaOdRQsD/Ir5q8d52v9+tuSdAQVBdkcK8sqjuwTc27M92WRH
b0IkkgIZ0/VLxQW5FV7h2P5khEkOONkQ3DCxDLIWCFNz+hcJnKa9o+wCvqwZ
V/+wR1PpTlf9ImkWx4BLmp4DeTcrGAtv4Bfkk/tu+K8IvWCB1YlFOf2wBpqA
xI43WvSfbXWgwVtLQQoazIHguL0LxzSbr8GREEwRy23r5cbm+fHUKzx9cy+1
v+RIQx49NWkwELlEiLWNQ4UU9VdjcEFmbTVBqM4O+4s3mA2LiY1YCDsjD/tb
bkw2nmEuWChTYQcBl4IDN/B8lU1+FyIhWVWeCy57V+b/3w/53+55riQyoEWh
t1iPI6qRKdCHzp239J7D+CxPcWPDUk7Apj01MIrJr5MRLrGKBebHLlLg3wMd
hY8491tk9jfM+huGjo5FYJ6O1sYIboHxPasAkxi9eJTmlqXs0oQfb+Dob+7u
9Zzu4u2ScaHpLnqHNcWVbl4I9TeaFLhLIHQxrsIN5PupjbER7fLA91TFxsDs
5UOQM3tABsqtKB+hEVgEH4ge65/vZwrG5K+fIYU9n+Kw+y3X+HQjWXeaHYG+
lrspz5HU7KlRgYs/CAz1/miY6G89v7jXBVAwdMKw1xckTDFBAYycK9MQv0hn
0lwdHV9qJuGZtIFY5DvppvTehfu1LeSJlxMVUCS0B9PR5ldYTp+k9u2qTYpH
ogXGSxh1tLt7ojkcHAMa8h18nGSR9hVXGTZ7Q5na+ZpLkbZNeLnBz5CN39tB
GcCKFLBVPU52En6IFApSYSV7o4RBg/nNklXi9RF7DNIPXxIddleqOaHo5q6u
vR5MmORWTH1lWfgdGe8ttkGtWGbFfHkR8lm1kIIC/HJydFRlLmAnnwgAoJ/3
iF4BokZFwPWWugQMB2QSlSy6wQR0tz4PQ3QKA1nT14LaMTXzkqTEhnWe7MfP
cDT/SsPUp4R+PPoBziODGNdFbVbD40qUX+lV1reJ+1X5rPZ4SU4stW4ldPWz
gY9qgOnwLH3WKK5W0CbxLaAs2XTpahTlW1Mp+coqhU4lSGAuM4Nkvyah6Q7K
DIBGFB8orV7ZV9CyfT95D+1brZ8hNIHRJkHCClCgwnpJL5XIy59UJEQFxe3N
VSSEwbDyLkF0DzO7hIOEbG5bSbtD1o7eyzgLtQaiajRkJGZTkiE5CGAMTHl9
FjeSax5RSSI2mnBjqUNQP2gzgducvySA+RtJxy3puJjzh/y6KQ4Z+/FfUlng
e84x3Vnn5ep3XxMBOHmiuLZcBSRp1MOowk+2jSkOqL7woB3yY2R7rU7kSLqS
kwC/9GOwy3sfoQvG/sQQOgcrd2gbhAAemJxTYn8SoYFY5tDpL42XW1r+0/dt
n+zQh7yFYWxvDBL2rcKOEnxtcFytg/u0F4Fyc34g6fg9aW8l8bGeuQiOFwyz
YLRUuv5F7FvUpcUQbpkjwYRqUKkHQxVRggP+UFw4zhFOu9dfbc1JZQLl0ORv
7TUq4TmeK4YxCgw4bqhk89pI7zMaujdlFsr3hSgReZ7Bj7fwX0jhle7YGLcE
OQGsmvwpQnfUEsWAMRIRI1n+DU4bdYIKCIS3qdCM+0B5uRnEAtzRB/eAQkKk
z79CdysDVeiTvMpYCNsJVl/p3nP4HbXoY/1dmxxF4bM3SeS87pWtD5EIZCKu
xVjSq8Jc4GZR09iCeskEDN5laVHCOT52JqdJNSlh1icUg9HwLEugDNbOjs5k
Gg/2T8s1vCVlrCRJZ42eCH1mVWzoYxq563XPM7d+Neg/Ojc8RAB/eo3HlQ7l
xiuJTyQPxntszK6WCnYgIivSPahMa6KHekTM6ILbJMfyL02YnVsezt0pW0/Y
C1JfTkHT/QCvbpIAOlfQr8rX6lyYydt/llKno4AolCAfUTHq8jEIjFybkRyo
4nwKlVWYneBtRufgw9TZ9jF99ntFGVmcdoLghs3tx62qikhvTen+ZK/iDYKD
OYMDGrLv+RNowrv2fEnY9wZnG9E9NjXCCmjZFKuJlcHdEbwFfLvpuy4S/Vn2
gaG1aIrIXmIitRDJHygY/hZYncmhDaukDYzYDgmX9HtMkwtIROvvARRX0eFf
8kwdVkfUWM1GZQ12TE4aPZ7kgsUqzWhkZirwNJy1QrNG7dw2niO5XHB4VE57
7L3ovDiR+PsOPb/bYRnGKyziDoIjpkQu9lmzs+JmeSrMQ0UDkHX54gTDNdvl
1qGNB/7v9lHY40OSXH63IQRZ44FV72+asQ2HuDs5U1B2cttBaj10X8BOwCvx
APDpdHVoqe27PbMiw9+/Gaad5DQUB/nRHqbR2UorcUk7kQheaJlx5MH/h2+/
A7HZncEz6uwyHTnZI9mBM8d6hNZhdZv1lVJkJ6Ga9zQR1Xa3VU9st6tPwHMx
XABwcfdBGNR8qbZbGy61U9RpsCZmw2P6FD51bsQV3dY4Y2o7tLkAIYhCEvuW
G0Nx4iz2xHy31jeYBtB6VVly0wZFdTffUKgSI+qlGjeNF3FuAB++BF//pSI8
Ygcjiqih1VK6WDepQQCgyM9jH6jdRtlCIMomBDPfi1pY3rzYug/HtpK0Tdbl
6Ri7MDlcQrQnLBSUVWP+I1nL7Ms6Px/odeUedGiUtzKzpGWql7CT1pJTb2AV
s0T4J7xIcKXiI2A1JIEdHKXEqW21dskJnpdkzLFZlqKbVmGqyjo5RuH9QRqC
Ay//OrUfyw4pIiNT7h7V5/TfaQfEThcprhq+ckTycnQsGqHQFYvBpf9DxqJx
wLgaHiFdhRbttcKXnxRgQ/mHqsSXU5YYbyWp7WQkdSPgjLmRVpEd/s1Pysy9
081jofSfPtTSnFhH2yVan5MOUt47tn7mvTqz2ym9vYOPB0v+0dU/R3hQD1ga
oeee/9lrrNT/FFiMR2FTjwjLbUiCfRe48FEN9Qb0fnJvMdCGCIxFJBpWAJx+
MVbTu4xckNbH/edo5h54HkVaj9Cr1cEJHzteAZmEXZZXebIapiTi51IfI714
J3XtkPUwawihdyZCQPs1URAL7e0QPs0NuH4BYd5hpcHzoBDv9Nzg9Ja4drQe
HzaAZbMid1CWpHm4jqB3OeUG00iPjuFa9MX2Wv87YorW3uuNfCmDeSTIETKV
KUnXvs5eTrHWrXtnemIFneVBs9xPrGc6zVq7vu37VE+dZ+f0xctsBvb91HOv
5l+5GLgyG5yals+b0ziq31m7N5vVOjHr13PcPajZ0gLj4m/1LF39DkBX3i/Z
AWkKwRbcCJgGFjJAX5/ZrRANPtuJStvSmlfNKpZfafuON6vKb5oL4h0nh9KK
VvC8ZnoRt62lLwzkdTvLnGLpsbrMMbvQTn4iiLfsCLruccyLWsVtZHaWbD7u
hQY0oRbFgJxY7mYF2wy+6m0Sl1y71FbjGS1aMnOs6mcynzYMEnLcBZQQIRkc
/YrhvJhR6xxHtDhuK0QIyPjdTjfva2bDi23lAYnshqJ3ehRl0O3/6xhqVQok
RyWNgpQWRKggBExEePa9Un56db6bTQv3np/cUnMp2Qcemain0ohMHS/XSkR4
Otp9ceehs9ZQxWwSzmlYm3Z0WGbvEdonGj/OIuvSPDPgOneYeJD8oVlA1rTI
CRxdi9Rvvqb+tR/mpedNGkc+pAtmGeh6wYUeqS4AS1fg8Qlwz2TZ471oe+2A
ri+ZCdua9wtZwafJDt/iHLL0SAuLiGn13yKfTGHwNdceGaceTckalVvscbJr
LH3U/PTlaoo9EqMguu6CY85htzsGJ4THC1w9JNDvhGYWFnj7xx0SO8JpA8GQ
lnJ/ZYJxD5VfpzfHg6BSUHyOnimFKMf1DAnGF5gP0GcCs5jecAkD9Gl3fHZq
9Dvruz4MP82HTaZCkntZknd41Y8/43ZM/vz4NLbYQD3T6XS3u27tJm9zgeYw
HvbYwNmZmG9CKBAIBVi6Op7z6VbgT/gQhwSveHDad+DC5SyPy33MMbCstAfO
rTrIDaDhI9H+Wwo9jn9H8RTdwuFF1dbatzfjc+gxwCz+qfJxFcVP4SG+le/t
rPnjMgLs/qqUzPgixIlc/lKt17q/oy4zm5g4Yxe0zwlnzqHocbr6IoWor8ga
cQ6WI3ehJZdA8EKd0an8X01uKRRj8/Q4IYTEZCui7FW4bRhuqgpyeCA1zIYZ
2eidpqTY7DblV1b9u5OhsZMm/Fxjcwuh81n9IY41RJzZmgzVKhnK64w3EGAm
6KshAZwWdtcKGeYilFMtU5nvGYEUMJo6w8cRgMCqi78/Yx6LEaLda5WlijP+
6dcwdVffGz04oDjUn5JMMudL6wQS6nf7L4yICc3yh9lhsgfNVWQGodg69m7r
YyWQ66Az85a+Sqztf5lxbWzYY+pc/K0iP3ADvMvBaiOvT9BZH8/Lz26VTHeo
EgOktrtQMvhI5vsCGDAAhO2Bv5hlF6zfBNrjlIi3n66XTmmomXgSALBV77QE
pGD/YoZnhxP6bx3OR6+3TCRvm4zp1BepbRcCRhMgFMTR/HnTRCEIZ7NcymeF
0YtXrv2grzLLeKeSqr0k3+IYdorcP54MA3xysXBC6o8opBbyOMEao+Zt0LUm
JSXF8KObes5h9LC3Xq8GXVht2Ec7tay9r4VlTGODVoeeb5U/VQQVadKGqUMp
Jv/uE0swiPeNB+UU7CMUOSgC0OU1K/ND+13b/eiPs1FQBQtc1KgaWVxeNzR1
2Exeqs7Y1LwzF3RQ50+6G+HXUFvY9HRSt5sQaXpd9MIv8UgiUJFOn6irSGny
KIdarfFh64BBJNorYNScEoSv2jMzo158LOeH11duEmS7TZ8XK5LmEpchVCAI
e4uDt9EDFcj3g05f72ECttIQLBkmmcB/wRtF7NxgtYX78/0L8UggqmGpOeo4
cXZWiLWVWREt3NESQPOt9x8OPWciwmVTT8yxZmjpIFGOCBEkqetwAfHpXHzl
ZI5ElbdZ9omqkSnYSV4YOBMOpXcWUqVm/GpHQzGcNvuhrAMvTbSLWfMYwD3w
ZiS6lH6qtSXZMj4DQcE/25v0Avr5gg+8Za7tm5LXCQcqlz5/QjD1m5e/hK2h
v1HqkdkIvW9ho8YH4kH6Qeqdyf3Y3BAdPEGHioy6arFbZRtktmQLrnj/hjKU
Wi9dfE7+HVzWpRxeXWsr/U39bMzJlodEbgCyVJcSzZEOFWxuLB1wHJaSzPkJ
MvSe+fXs4hEAUILEZB1X9HSwuTuSJWaJ9fHsGvkrwb8JJOivaYUnUWWIFhba
SRhz8m0yNIbHJo8ctBb2SZR0Z1ewVVO7aMW8BBhG+OWxsKrr7o6dcDXipOfe
t7wbY/CDav4EvhcYryD5lTOpE691eBhjINUD19gCmotTx25UrZdNR2L3oYJ2
jzXRJc7HhOmfAeGQaJACcjNnBce7BVn5QsGGrke41YaFwKPkvne7SG5HuCKa
TVwnu1OYojfvZyApBERFElHfpkqFQuGrfphiURw1tvA6v1PGgBxpFzPo2bw0
Dl63U+aQwwK2s42AxB7G8DJrtMTSgWdaQ7sQpVHDHqCH6ATcgMvZhIXz96n2
pHBl2h1UhswZGPY8E7rVjLX/igdkA68YWKSlCQdN0ZRkGBUSQD6Is7K4PkzR
dA8wOGuOItoMJzefi/cqR1bpeDCFIEb01OGLiW5Ur5hGmnGbGm4s/RslPRog
KybJoU83LDil0MM1p1jBiNkGS0Ov1ZX0fh+IxYvMdGs0Ov0UKv3h2uUTOolN
6aUbwUFNZQ4nwj4v5YIpOzzACjwfq9dBr3+kjun0ajD7rlzopYvxUO5c650E
SM2m5bSzRfZPn+6N9F/fMf/+6xQ8kLE7hUX04dNahago/S+eIerDXTHSMYjS
vrwmGinI0mqjklTfZKx7N9oAxWhkIE6WTkpa2e+jCPM5QZH+SWm0JMvqoo54
FrupuPizw0vCmBn5rdX5GZTdFdRsDZS2POiZRN485srtYDPtGbLsLlIWVdcH
FEkpgFkWEF8ETiLV+gaiSgxzteNG2VRM9dJpwdkGzGncRBEkv7NfhXYqAkhe
B4pIUcopSAtYnKkT8z32UBAu+tEKun0byBieCEx/SCkdR98/X90Ie8l89quO
MVGUYq6K4jNYalxfyKsAipI2jhYBZFZj/zSVQK7ccy56yuzRU91UcFNAKSgs
US/MdejwTboHcPGD+8hrC+NuAy/S9gduNeZNqbah/teo+YKT/q2oFi1hUi0k
81BRYMtVxMhNVjo0zLQhkeEycgkTfoGjX2uMhVQHnk2NQPoeWnsEQxDmkBDF
W4X7kvsrmMQa+6gVDqmdhdwRmKEtkwiJYjTsk5SM4u9HXQuS6GgDDm6/ZRYJ
co5R+LGVnkS2QTSWpfg8t+xxY+I8YshBwpQXcQh6kGbLQr+E7YzYbsK18cLo
/L0nB8rV4Wezja3qb+KQYkBMRX21upDI50BgC40oaKUtTLYCfoRTWU+RDTlC
nrIvPm798BisPSsAOn98IERHEfX6dTzPXxqaP2XbykCuRlTxTIetz3NKDxdW
vRe9ZWAUJcP1DVlijeDsENmro+eEOG7hUvlr+I4Yi60kBVneKkCqMPqTEsIa
hen+pfztujs3PaR1oGIkU28tmwpcOgUNRmxaTXlX+O0/p/j3ihxCGnhZkFBc
hEh+crauFDG08b3YA172YLaV3dkIikDgZxnabHVWqEA2Een0mQqeblxpF5hB
b8lycGRvgyBnQ8Gfgzse+3EnCvKY9gn4mAOrPqP43EeIR1m6ylSVZ26454+n
Ts1WLngBRvnd38nb5AFfKO8x0Mp9ZPOIfWbYUKEurMBBbVIywM+P92aGeJ9o
mnguG7gehdzdk/iGz/ycqtTmNiieR/2ickmwhIRJ55kYq5Kwxqhtz2oNEcOb
muz1NbyARpziJuV2Cib0zUHrhAhkuJZUjzAV9B9SkdxoHgLrbNQl6qYUifMY
/MzAk/PGjX+4vKYD2f1njQWpN9hRIpq6mUPn/aYesapvAK5lvOUxDTVBFiSx
9+xVCg3cQDdFv5uySw2KrD3neaDI0hzrVCJ51ueFfqrVT291zUMFU0SuHU9o
cTze8Nft3+D69OYVv1iE3AWPmN88lf0psqKFU8jo2d9pZxjME0C6R198+b3n
C6xqkq5YbdFfC8sL5sXImbvrvPh6799Kkta372VFXMN21UItk9Kr65Md2syL
rQvcbjrTyUkdYVhgWflG3S1KFsQXiorAZzDKEkwvGrMUskygb/l1WdVxdNdW
RFI76UI6SFWaj4/4SpQBN6lKni2wJpz9sxBf3VBc3rycmFUP/6g0Ww+EW1x9
WkinB/TwB7lPGf7KQO46bQ0GDqFkMQz+VKPOEH+WirG6l6rV3NmFz7P4jiNw
zXLp1XJtz3TnM/9gSne68dsQDevds2jE3oKpMGUKC84DFu8dWsqSCdPbUrUy
QfuZTL31QCnaVDmmrJZ4XMRX/2Y6P1p8uT3kkYsgnr1s7y1wM27kkkQsc83X
HzVB7tg6L3LtZM/pmrSTrDLqDu7Lq8V6uuuZabiylvqH0pHalPHAbS1/XMTq
VQkbsAQTcT6qx2904Vna5ijSqbONb68Bjj7fi+6OctSTKUynyDMj/gYSdM5i
achGn2QEYD7aie3S1hujXiBoefD/U861a5zkDFSKGXl8PsSujJQkMOJ9yfxs
TQS7q/S1O4lY0aWY/912yld+b/1SmOw7r1x6LtESR7/SWEaE/I/N/VTxHLup
tAcQkxlFqTU6d1a/TAmMC3l48ijFFZlyPUpCtjFGEOJYkRn8z5V8UGCfdxNu
9dJEG8myx6X5AX/bniy/dGOlePrN+6OIxFnFIxcIc+9jkYJSePH/Q1PVPH/o
10e16w8COV0HohKMSd7ertNWZI8XyouZESZEhIuQYOptyavB30F7xZHM+vV5
mI4AcCxXgwNthyGFsL/qpE0axaWze4t97druDhUt2GjXevYdVIXc1xNA3N61
OhrhOCk/qG8hUgMCb0O0bsnpkH/b88lkHBumG82Pklhi3ZTLCJ0vWFHd2pvJ
koGNJ0L30X2fyT8oNzVoQTQdX57Gact+Y3PNsCwmLpoo5welPHEiXyIoFnZ6
Ja7RLXieQZtj4Lfq9dD6PB05tPRlHcPINMF67g2+4C3tXNeHaIa5XPbdZhyj
xrrO3mxoieP+DS+F7NaqpH5xFdpkaHzpsZ3VGwLnTS5ujDyymNlnkmzSk4yx
YI886iy2q61Mh34svDvamJx3LL+x8A3ELhsARcitFQEGcbnc0oBey8bvL4Td
pWeOqAsvuk1OBEQyxyI3IjLnoC0aj8FoH5mBDD+NY5b8ItRIxA/ncP9hciVx
SvKJRhf9yNiU0Me2I+y4QZ8xd6+3abGAtlaFJA3WcqXG/Hjzgyln/GXVkouh
x7UK+Tt1MfCrWNJNEcqV2xEOuYPLWR8DyEwNBNnJm9dys/JTy6Q0FjDcBGOR
gIlmL4Vx6dM4MW53wOAZfDRce5zq9ToabPmj7/WjbffnVuCAi/Qe9GlxnEgh
3qzC6I44+YYPZ+P/urEbnnu8r+9KRkq6M1ASkhY+Mc9tqH6U5WJ9DKAgUzb5
jTqXYURidDNujZDYHe3P7bWuO7Wnro1srcU0wlhS3sdnipcsrsNEAWLXRyLr
C4UbKiGzWeJ0oouepLa+DNMRu3K4A5aPWwglpyDPeElLE2pXbWWseKu9p7ei
JuGZinhpT7nzUv43mkj9OPPU0xBe4VzsdOgeKol8TgqEnZabldTpBZnZaivC
zlF4I2f4BvoYAgDVV8tj/qoFdl7JEA3eYb7R7BT2y5mXGYgH2lXyrnmw/MW1
0+1cmQ8zaF0NV/WhZId8YjvigIQnHPvuOVTLfsou490X1lh1du8fK1SN+9fs
47Q+kMNZ3TQAzDQI8hswnh2r1DDDeLFQOjqRgqcLSYA3Wm9I9qvgKZmMyKtt
KSAf1uUH6c2f7Ev+bpIOOpAThcvljtZKka/olpBB1981/XgtUkkadp5wMmYJ
48fN8xxBLUSZxBBlFuWuE2ss7mYLPc5xBmcbyr83qe5NxB/EHNeJg0tPgbQo
NlwHz4IsgZ+xRzcZbH88izq5uV4Y3L2XWjJqbDMwr1lo+O2X2SjG1XELdK0g
9mgKlP9qgSD0mDw+TILAdBv6R7Oo7TV9TG2AecLJlkR1AXpd5nIzEYh9RQCy
+8oFH3HlY6T3HtBey93Yj50RfgKsoMUsQ4WTd2lKCWZ2pX/oNdsMP0O/VMfi
3XTX2GQunM0/OQY1xKAGUxXec6I5Lrc+NPxhzugLVzMWyKSjS8HiswMgNCon
VRPlNE0Z6A4Ms50GSQstSwRqCSFr+Eu5cQhf9ENMwbjpsEcBR8wo2qPdyrtm
dRGU4LTp1HMSR9iAvRKXkkBz8Y40WHwlDI4rkHVIhHN0qDDd48KaMkNJKZ9v
pERdHYhP0LJv3mJSQmihzv+IwJDS5Ds65Ufx9zJjreSLU3SQjT/+oE8AYHiN
YkkZVDT7kaUOh/wzH6GNAvnIb0/YjnDB6FqQGT8g9epO6LBzWPIqSxPxz80z
MlsX2fD+D6FJMheuzs6gEEx01DdmXcT0GmeYpA7x+c/fQHMUCLJnNCGYqxHZ
u6LuuCCs0LvwEtrxCrzubBLk5nZWvscTx+E3jFIrC28326oCfbuqLIkSG/f2
k4JmHNdC5hC1VTojObohJ983/eXThmmOQ9/zwEzNSEZArDf5LSf9f0NRVjyG
1zZe6eieSOmTI7Z4/UMHDDOuCwT6Rl0/DtaLTHFiOi5EfVP8LOVVWAqH5F6v
NkLs5LL72HzAui+k9D3kaDMnuehysqb8IigF5FGxKnhYe4cKQWDgRMOdx8kP
XlAYIYfC0wy24bdZa42zk4HAYVTkhVYIeKJf40ayiKsqJCA7XUwx1OiqJ1Zc
LzIt7ekmtx7GF9TZxL+WZfZ1PoonMld2hPMBdLOTxuUKG76O0FoxEFXKPnxq
2IqrTyd9P5ScT0s8GEqZ9sWq2edP3R1iUtwm623Nm4N/AWPNDXeDmfFK/YcR
9JXwwO7NWlJj/SGPfH34IJME3nWx3q6pTmlL2s26oW1ArDFyfOuMqpWO6jr1
2jL/XyrIOhC0DUK3XE3/0KvGIDAyIP7TjpmMrfpEYHDuE2nVg6Kn0e0re65x
eTmbqtq0tH04wKFsyWiU71stoUotVe+XYWfX0Vdl2XwwnxOui1G3Ok9/6lbi
dL9KKkfGROBQ/4XTYht6Tro2dqV/t06MuiUBSyUWnAjyS1kL5zKckHpF3ZZP
buPj6TEv13cvGXJyhEfbM9HaZeukrnUgj3W4DEnbfSPpO9XNHGFe28V4qE6C
/L551GEwjBhG0FdwkxiK+raQmSOn/bdm/x1CNt1JQYTtf0QyXuWputnH7pym
4LTVUjd+woDFfwxMmO/Vv2c8VM7ylffiNQWzvxo1ZNTXy2Ii9amSWjIUfMev
SfCf0UI9lGeKosp5yMiFklxIO9j2yvmlQA6R4gpDeDJONmNsqqO8f+ID+V6K
T7nY3JIm0iQVG1rV65er59M0xjZwtzNVMmym6qRb8Zxi7E2Dnl9mjGkugpbn
WVAbeF4kuwBTQX5QIDs5hZSGs3TDab/2xLrkO2NynnpJuuL26jtE/GppMEFy
VnXbIiJIFORYoJPi98Bxg+Lnplff/x9/n5B0NzEUEiQUZacfYMyz6Ad4AA6b
DFls8rrQWaCUmuHDlRqWyd1ACi1DYq7yMbloswkoN3bTgl0oD599HQg8uyNP
eFRIQVdme8yQDEFhvWIh4LOc8hsWOaMVsAo1cWhGyknEdERJfewET6F7c5QT
DZTEjxKAByyRC/B85uOpv9fmCdcLOtqxWykwAhAMDmoGI0nUBu+bY3Pr087q
wUXXxuD675RhR9n7K6MGkRuPoL/jJY2OAhl3/NnolwBvRHQP29Z98aGs2O74
zjG26/Q6MzP8qpWP6A4Id5pJHODIh7OdllGNhtykQUsoWzIwoHAb4cQVnvN0
ACIhb72T8eRfsOrIqaEPa3fYIXw5uZQHWLD3LVIg613MMXqG7988iUJp5p2B
qStrlW2Cbel6Qh3AwsSg7mKuWu2a4V6rSf4S8w0r04PU9dXpCMeLckhGpn1x
Sm+rvoaQ7zdlCpiMTfuh+69dkDdUvh7h/R9to4UzyXROhq01Nd8oHKsRC7Em
3jfaS0jXvH7Te8tgHmEKUYnsqooA4Emdz1baPhRJe/A/lBx7p+OY2R6Bczus
4mQXa48TnjNgYmHq5bSihXZ6LJvTLdXUbbVaAoWvS5D15gKUCQO1EBjyMM3X
jBEjs2lC7JAVupODocKFHUpjWbcz4FSqg6M6S+Na/xg8RMRRH0TzqrdSFjjS
5BWnFsYKWtYUDUfofnNcPVonvQwBUVLZ7FJC5FcTFqvCIAEc0aocW7w/zuU+
dqsUvRN1mWTe0hS3/3GyyZyGOpptR6UTkgA1as4Wg/u6vZ+eO3CaBXJCdGdK
4ob/+REGxTtq+Esei013WB5PHr8Vb0MAP721Yae7mbIuNmSFDCBxG7Z/Bo7U
1lNldkEK+5DMYxvHe1BUVzVOlw3WAk670cAuQkcasG3HCFwDezGa5N8S6PjF
INzSAk+HXa2xHgDop+4Snfn1B5MxoX6AkAYcvfZVAVO8uMHpx6XuKKjqehWP
YMOa1ClQYVF7jJwxvk9KEnU4BeTycAnu86OTRLKrNDYRVEn+g6d68hpyuSfo
U4ZfreRiuLrx+lsbfuD/QMmsv7lm10IXE81bU/e15ceGD25ZEPHF9BjKdPun
kfmqlHoIiMNiwnVpjwD8fDzmqqZ+y4eNdzvpXda96EpCivJ9jrNHYhMSxGBw
E2C4Y9VvLDshWybBaNNmwIErOwo1OIhw7BsvOEPsjle+96SDvG694TYnCXY5
ZQC2Z+juyDE8KY7tfhtBNeGNYakofdlQmeTQZaz/mRFl2QDHI8/+Xld/zxHl
BgEQTMoC05V0kekDduZvgn52mO+C/LPKy4VamjQ86yrW38tWkJfh5L6fMF/H
Th42NNC/9WqQRWhYxXlqFU/fkjX/sQUdsdOOtFk4FjZWuFBJ208JAmn44dTF
Pk5YmCR7oXtiUWSoFjHfPmevRo/Rp5NQnIsrhBoXoh4VhEt9A9KnUDSbSYQd
IRMRgqQ9G7y+A231BUgJC5PF4HzGPBHoE7RCKkn7cXilFPcCPMby+BQ/0b0O
9NGiADw4tLpTYnwXDe2pPX2330cNS2uEtc3NTuoIJvFWwH06Kg+zEwurEicH
2/GCocz8Sv5DStYoto5jmj1l3DrWGQu/v15VMFv5B1falTDP227VEPZeNlIl
FWFIYtXKJ9ve0+hrkn813hXAPaWZXwBk1A2EwhEcAhu7Nzobd85Ws/pELo1Q
NYpEMdYY7AXQbiVhdDZtv6rEBugLJTQefRc16Jtf2GDfA+ZnUSO5AQeqTwlq
yJf9ExEmDVQN47mNIC+NiZaPTNRgG03VyrSmqqXQHqMJHhf1VQiuLr9YQp0V
oJsUgVEQDUXPFfEH1wrTQgLJ90nj94/pSeuuht1jjg8Ryn53ojvvfbIC3ykO
f4jwbtRKOqzp2iIeYM6A18K+WTuqZ+4kRiVdiZmSU8D7bSPF/wMMGCEzWDda
mjpa1jQY+XSJ7AQx8UsKUrO4aliQes13pBoJP3fu7b60+tdmU0eqAWccvo7S
JJ4Yfh+wSOenYieZ4cP0L8uZb+I7tGHaTenwhmXa3bLVNj4z40GJuEJGIj8a
NkaMAS+X27bwc/c4r4sdcUPWjTk6c8mMA87klAaCxSvUuTu+YjJqUiT8ED5Y
DNmjI/iOUCo8tsa+mhLA0nQy45wqm3n7d0h4O7X3B0AyVQA1CBZnmFPJ2RmZ
b4NoYmqRxQQ9nsw2G6PqQ+utKhLaxleBlntkFFWNVNyoban7bXp64K0x3Rom
5r9VjBaZHTP86VHCDRiu+GEL4KQiPSf00U8B18enz43MGnaXrQEgAO4VpBjX
+RUHIfv7q8BeEaHRbCOfPtaDPxBD9c+JgbgpXBNnKzENjWstDbED944UK4xc
75EVexSCja9Wlh0AufsFY2tGS9UTR6zPcjHyP/p5gHr2DFAQVJF+Bnx2ya6L
4WaZN/CnYihTZvo5AO+bEOfIL8VBvCDp5U/7UA3aMMkPkMQ6dWI4Bdo8peRl
4BGAoXikl08FOnws6ou+GWHJA0nmyWa4SCWmlXIHVukrn0xFdZ5uxwuQKtJr
BGxg0WFeLUGQz+mtcmA/5WWuDw2X1ptSCGRUW+azi8aeNfzISk4qeuFriBoZ
Jo5sK5qqq9xXIBmHLJTwiC3kLgW+ULmsHJw0b5IvXEdM77tpBA0GppvuqkIp
OXCD7oxQE7yxeMAbJ21Be1l/l4jw0d+NOR53K7A/ajJph3qPhCpQzpVETKHM
Ojy4ZdfMKwPBhSoV15QLEBvxUQ7OBvM4BPziELpFriWCTmK/YxPQ4c9kNtwz
FXjQL5pRmqjHyYm/ikebpNV9jdvRPUlu8LIm7Qa2fyGbc1QfD6KFPNLaYizo
WVlvdumgAYU7tBGOl1+f+kIG1QbqqVDitFSsSc9hCjVwzRPI1pkpyzOfoYfG
dyfLU7yrOjn0GUjOTnKnfaXaXDfVYBs3/vwnG9gucRD7F1ONWP8d1Sic1ZB7
uB9wz19qO03PjIwx6Y5L7WQECrxDDzDPLoZ+64VJBcgFqB1jLBzuGiFnpPER
N2JRo0v5KQRPFI0v7y8UyR1gOWdoo2uyLp2kuF4fuaYeaoFy8Yf+usN7sydy
WKDK1owsIIg4RkEhX+dIdWhcfRvS3CK/8cfBDI24aYlwO63UOKfvNEpN+Bro
bbc7RmAYcMbDxtY/eGaLxrvshbMPed+x1wVO3secmGpICoapq/RnLimEQAAa
Amp5Z1djNpB5QJiFcFln1ioj0z4JVto6hHz2qiX/y8yBaLmzyDEOtde3IaM1
ZgajLghvWTzn6cbErU0HAvMwo+MAtvd1uu1LTnTi//S/dy/SeqY8WDlNDuSm
hT1x2LQ/4CIhcyQKJ9E9ZMSKoiqqK1n7L/gaHB82g+GAZME3tUrkJoZ3rlrx
M4YlDmU6EQtmtaIOUM9FD9SYKUSGSI4pAwo4lBsRiLztRDTcsa8cPKz5+z5/
JKF/ttPv6twsKBJP7yadnp2L8MW7fg1LtGXP6pN6LjG6cZX6yLSFi+GkjiHk
dQqWMTe3lQGw5W5cqgv7zdNBVTkFF1J8mM45gzzielZhXDCLDNe++Bt9/aEC
52m1aucQ+HFPcL2B5ekZeAnqM2mQUpjIJn0rvO2BlmB3aCPHTzufz9CdFUSx
LjSQd1BtF74I5ShDUh5NgKiuzI79n5UgKD7+nECfQ4Ej6rbhzHjgIFXidFed
az41OPSzu0zHJWptvDWye/PgIUJbuJrRQzXZrg9Ahl1Mgk5ToFBRCKismUq0
YX5Am2VPmtmvpLLgnAGN5jwnCSNNKV8SEoHyHKZMpyDNeB8JQfu157fTa6vx
MHTe03eG2pmAQ3hxZRjESEFm4fl56wodLphO8Ia+cFH2Qv+tCLFrtHMhcXQa
4Y/E3iYQxNPSvzJE0d+YIG0wDkcoKcMGrMbT/oZCnVjt90JteQ+gv3YviXx5
0Z8b054KrV0h58gOPGfGWgl1OyLHUKywy8uBze3WoHgczx4zv3NPwXSGK8jq
27shnqffYQbLAKFiPjforSv980ZajhR+fihw2946TNdwPNQJYFFiMLLN1x7f
QSZFkAGyw87bPReO5kE/DZUEIhX3vNtf75DphXY6nNZPRKHahrrhtXc/1SGY
0QQNnRYR+GiKOlUC7Ft7/a0LDeDcMvWdNdU1qlKl2exG77AHYOZXWW31u8lf
tHpTiaof1S/YSgSySU08m7X6iFgbcmVKu3dLDKYgd5kNE5vRutYEsN4wV5W9
S8vw/KieonEFs25RLOTxtSl0xh5TgJRVSQPdEvse0fCbpeUvurY5wupjQPcl
6qP6Q/QHsSddWdzDjcCQHQmge76Tgw03KYC4aL+xM8eK+0prebt1dxjCc/Qq
l0xwaOioCkWcvCN67aAKvEPXJtYIjsgSbZnobj71MWhJcQDLyz7LhgstMdUS
1uYQyxPBsQF+m5OeZ9r8+92y9tLaueKQOhx7p6wDEnIBMdMM3W/tP6qXwQhe
fvu2MDd+ef84qVtd9UMXSm2q6p0lfPMPrIF7yGBsLq1LTwGyu6kt5APMKQzU
p6dKahCB95oruk2KFMMWQ8IsFBHDG00WHltXgnQnSkPUarnKbfwZiUh9f6JG
dOc3CiYaA8ssWnQ6CD6wRXuM63SfjWmYJXIJMFIs5c6yroVDHvvRqX3m5x+f
COGMxClNqOfaQiXBzFfdi3cQhukXeJe6rdwQrjJXqSXgnScQVHx4pYdlTBMD
pxBY5r4ncvPvP1aTrpkEBXrLYllmXorF86t583MZgll6JgWkba20QLoKLSkI
MKGrzRdrWAYzL0WfiEceh85f6UQVvpoQx1D0je27WS318Iqp+fXNcZOzTn1T
s3EGwHggy69o+y9IJmMhPuHsWTnP55zvs3uWJb+3rOdBovauctawp7SfimSS
NovtanyyFQO0zZxvAvc9r5TFczlJ/2zO7Kkdn2JiFooJnE6EraxZdXGPy9cl
jrczUl++yHQfyFP1zStYwAkpsRAXuQAlAD+0MRK9d4Ub1Qdm/FNn3R4tLrom
gtfhRhFdty/rQusa9OhEcaA0onAX/B3mxxiwCxwdXbKa5OlTqmxwNN/PdiSs
3kvijxU+xm+twQ5IuKfojqNxnaImbfc6VYO9xNIy9W60ztPukdrkGx2gzv1v
rxTMXcC3eIuNaTQall4Vw/FXudb/XKs+/B165zfw4zixO+D3rrPXfZKO8nW7
LBrlE7PGiuhy3SewKQEhyNv8pabupd84XbJX5UdNx7R3OxHs6Lb7uRLVk3U4
H2tV7Ws+v1Ccqgjl/ey3ztX9aFzaSLjc5PbDBw72dG65a2eWNNxOnoqTMAfA
8i2XHr3XivFZcZ8rh8jn6ZEj5Py8V0UlrH7zKGQZrSTeMNmfdOT6dtS0q18J
KLCiwP9ukgbAq4ZWubsDzn58BXxOZIzG0dcu2kn8W0ftJY0ZymquN84SNofj
djcr6OZpHoSxGFEkqqADbueDZJzDMZvMa6iC2CJ9oOGnTSzNjoNakz+ViojN
q7Btsmm2WSgoN7AiIq33SOeVLbs2HRIPU3zvP0GNyKOGvOxNsXSLJYv+pmee
S3YAMPTxYWssnObXA1CbJsre4ge6TxAJ53OLP5Go2KEf4q8f9dMVduDVFot3
ioHV09wzK+KBGWbmxALcHTTPEBK8+y417BkZqwKGpDbkR4Lj6U9kPXwqJGg/
2RE2UrH0rzYLWknBQJGadl0ly0lHHdFYVo9bNd+4ukaIcO+pdftBCsbVBc1q
/y0C2IgVbdThqEiVl9s9o4GMgA3DkAv1ogjhnj55vAThyh00wcwdFbOlmO6U
jJoO0/5+X4YclmpUY2dDgJwxuE639+F7NzUF7INpvAo8iM9hK/r7G+/BLuBL
MxAqKpUyLEw40AY0PcjHfjBQcwlvEU6QtUHHmRGcXRxSNczrd8weycNy0WXh
WaNDyjpvOb/jRdqi5mIcSPGuyG8CIC9vJZmxzmujQGr93VtvD4mJprhVQfEk
yXhQ8Y+2K5eSvP9M1UHOdME59CLlDopYvrZ2kQCsPmUKWkLAj3dHxaLqm1pL
ZMA3/d+ef5Xr+62gPE+0OaiIEEdudyWvL6I070BL+LXaioQVnVdZBEWfZJN7
4T3P7rNgSchQ8uOZy+MZP9l1brIrynlgfoMKFBWUmeFC/af9hkd3liWvgp3d
8MDv6PSsxg6OeC13XsxZS1Z+/x4/z7XfamBGi1Ee+pE7xXogNksCBBGH+txv
+pKBjozenexz+xADc2qdE5HTdmX4mfQCaOqU5PwMpwHSmGMu/vzu+LMKipMx
W6xWWzhXzKFPtUDFVb1DeoZSIS45JjgtPX4aJtfZaLOq7WIfigOYLIMWIxVO
fHZDB7NVFesRY8PvQsay6yUN5Gluvm49NsiDO5N4SV5VNjLdO+DTb62Yc0HR
fexO92jIrl53Kb7jQfGqTyP5yexQpLN04Evr3Qu861Hq273LEMeXlqUu8gPi
HoSg46zPepxPR/vfVdNG3JsVkeJayhMTktF1xl72DTAS/pqZWZiZ+7LPZXBj
QtN7ytdEmPpCoo/WGZBDmsnmoRTItqiXxNycEyGFc3PqJdJxH3G1QF5wPefC
oUpg5PDl78lbxzjhr8TiJ7SrQ2oqr5Z12Q8luN0D15P8LgCHIPHwTlKbz397
p6YZ2tCoXzZWz3Js+c+Krt0ZCEb4bARmUWn7GL6zz6mZylDF1Po7xGemeoIy
pfmct+BZDG95o86mQcvKSN/gwuaKrX1y8ONri6WfEwEnbWSa86+M20MAJbzT
EWGQvLOHbtM8xuR2sHieS9msmQsLDHsHB+GKMV4M57kFDOddPC9jR5VlfEu2
nlO09tG9aKIrBePckFe2lyIYIIDPHeMErv8VJt0RsOlMHpc/lHRMdpakALjR
SG/Q9ab+KZg+p33wbN4piwaSWlszXW2vPIM0PVywCcWRUtIvrepswfCR9+4M
OqtSkN0vmd1HAs/Em+pxcFFNVQvS6dInZAXIQqIoUPz+S7tLRUCBlxmxaS8+
L4uHxkvjhjaa/VSTQvtR8UKzKtKh8bIXObkpUflr0Y2e7+H/mJTjM+DEQMI4
l9EvxRJTWuINQ7nb0AaM1hn8uEEmkhLWewjE/ix2dyz5w7NyRTkTZPnbGRzE
+hamqJyooQOwZBzj/TiuRim6jFtB8vHSYyIZVwzvMrDtZBd8tK8mNJzcofU8
9fghOqatxQr0TGV9QhtGwE+5ys8H6WyHfhKkjYUktqRMIlvfE8xoKBirYz2l
+3wAphkF5EFqHrNOKSQ6VLr/UW/uO5Iuj4IR7bIbVKw4YVACFkdL7XxmoAvv
6qc05WOtp4iBaJ4rK75L+0tE69M4+ZnMy20i/CjoiqdafA/ydaWJ52/pkYuw
78uXnRXzHMZTOnK43HA551GX/DjOGTOp4LTVhb5m5S65s1SV4/bgwHpyx2mM
xxbeV4t8idfTCqS0hNqdU5vi1BmTHt+FpplH3eoG2QMuZcCOBMr7GkSfNXxy
F5PENvj/wJJ699eRPf2n7iI4AfZXdFlUoJ9IY3NS9+5vVgLiZ0pZzRdgqFw8
N/WxsenqzEGiSHqNkUXK2l1QDkreKjq5jEfGVhWOjNPNRNTu1avdcabroCRP
HowjuJ4KGZTr6/zsU3JNAlS/1BHDiRUCUIHxi59XE6hRlXofdbh5Futa03aH
S5SPVj/q3laSEyIl4ZlWE7sFPkMpriMfD6VEXX1uhNWYL5JKBVt4UD5y/uqe
zi4hMFyxZHk2mNvO8Vj8LtOQUppe48vvGWfYcebP5DZWWelTYtx6lC923Hh/
QmXOz4MclrS4XqEwtDvAqbvFAmqgAEQdUjIR/og/Jbr5epFUa1a7XG+2BMLr
wO/mPzpA7ZyCW3m+2vt3aJwJiIT5p4JK0L/pj+a/L143bRUJnPGY90DsCTwp
ACiMEi5Nqq5PjjKd0DhChrt2yYvWPyjvuOz08Vhq/sKTPtxP1nhlibHCQRkF
MFWoITx5zhGl7cPI6asgvCIq8urz4KWthzYBOcmj6UQ/eqagL80CcOfdocUW
D/JWAQAcTRgFm8OHLgAZCO3eHEWGk5E2oPIia/hVKili7DLBMFdODBqwLttN
uRFLkcmFjLE+ptnlqAKtpICAHcQ6KIB+eY1KaXoGXNyMGTMtG7Pi1cVwdDk7
tpAuyHeyKzC2k1+qI9YWSULGFJEdux0NONJcjaegIw6qqQEv/NSP8kEZR0bG
93UygCLdy1cQl5ehl4zjRWiuGwcY/IYg7sO7vYEB8KC4HxatoUYYkhu5XIlP
YliLwnVB8Nrw57SqXQ1dWE7LckmsrTLieX6GyB3GChOj4QGmIRY2x0Xp5qz1
mycDEJrMabvpcEC2o/KRTSQ9XbJqOGcOxyy6loN2bIT7BWiMrcmztMuB6TUA
ynmoS57859xZSVa+ldvHPHpy+28QeSOObv0GJzCFstAveAYThRAHjZsxO5lR
Z6Je7qKU2qxwgg8Gn6FhNVKkYZpnOFHA2g9XPQlOizpiJ/iH3bkAgECpcnIb
Bab1RVNwi73zhTBw2KToqrf0Gms1w2hqFN+lKqOSByIc6xsaPQkH/Ep0g5mg
HAhtz9qZpRcPz0SkIMjkDKNhRPyRxKJUOzEk+tqd4s7KJb8iAoMtVFLQ601D
cKOdKmIe7+WkyZGQVpOtR1lvnNGGNPyn6WWuQhBGkbakJwIwBYDRrBctIBr7
3dTE440FeW3ZrNgU5heQnbVIfMKavYzF+I3nPmg5ippGZ4TYEDGkTuxN7sR/
uY8dB2q/uV8A3u7FJvDMrYUt5LRGB/yuUeysgYFZ/dDEBbsRB3IgF8/jItSw
VjhsDcgTRTSo0U17Qwpn21bziGPXCbvnsdxZ6fy/KYRZCJorZjAAulN6OW+3
8xRyY17d625gNJ2erfneAKSQPJcQFO1gVHSma+w4zxVmanO5mXDpYP1RkEhX
gD0Aw5QeoHrUUyLJkKZ/jOYXBLo6SBObbbzmxCYV1wH/GiLIA+uHHDUC0E5R
Nk088FlptOKGWZBF66HziY/H4ZXiYcbhGhLFfqVvf3h+RiNq5yr47PkhoOLM
uAr7GFQwbtOomahEsXFQQ1eG1817GRwjR0AB7Jt4slAPtYRA+SKmOky8Is0h
T94Hsc3Lm1Cnp1rOjXP/2S2LKZI8kmHxksTTMp/FJtSo1qo/L92pfnwYmPvX
8C0gsMSR88wNBYqAGV2xNSdjSLdSbAoCDs+5VW+yvw1rol9EdnNU23VZUwGX
3rpKtUU0M8C/Hj7bTxF00Kp02+XjKrVZjzxNBmcsQhBVGMEsQUu+p5uUIlj7
ojkM3NAY7HdmYSCDUL7+/wzkni10f5G2YsuxzCxNya513qO2LCNkD7rshH1N
73ZPtxW9MLYYx45qPUkFa5KfjcxbcjNi2lveKje7vbMIByILbKtcN19KEgm2
xLWlAtx5zOWBXohsPKPPFmmHMC04/CQsrWSoO+RXllrbbvCEd23NfJJcRmbU
crTxr7/iLOBFJweYJ71SkWT+MCLsIksSOuq/1/UtHtRBozBoBZ6QBlYeDK8H
Ajh4HkTRcmTqVHwvCyTWBqKdD+j8O0615zVF5v7fxYiI9yRyvQOCo1m3oAgJ
fotJNZmcKmYInDOb40YxCdp/T4MNvU47UCjB24jQRTfXzx4VpoI7d9ybAKnx
H2GVfAEYTZdu2BuvRy7aiQUxszXIoBnY3Xv4n711jeDOO5aUVAqPsjeHBPp5
y2YZB6LnYwXEeT0nKQBUJLlCe0up5NM63sQ1BNQU70qb2KXkuyrQap5g8FQY
vsivLwVoP7Ldrq/VbNDdgEothSX2+nEZ5+4FiztGGdo+lWxK/WwN5/9NAT/k
r/DTbPwteDGS2LDjLpubqZC4BuVHs2oHT9jYBjCeuo7uj14Rqkerw76kasj1
PoTEIAq9cXkk9w4YDsTwdhryY3VJrJorjMjATRRI2VTkV89QLKkoGT2N/Vdh
5aXdBq1+1mXjpW004XibU+t9/ERo/CqJ7tuAw2BXZOmPOmw+ftT7Gu9bBqQL
ms4nVBzMt2LUKje93MoHK1kjALUMELGSSa+6K9/BalJ5KQdH0lTxx1h9zRwD
4EVTS8wmmiGol6QBKOe6qWaIoGgb/XClV7zcDwfXDLm/qWozfjNosD3hia45
5wK1pO1ZfZl8LRMVEB3bGihFsmR028pHKbeAKB1tRwyEbykXpbmgoyTa+AR3
A1LrDcwyE4lF+6LMys4UNNNdFVjk3Yt9uFdnsJkwOrNp8A9PUYU362mF+pyX
amnPm3tyjtZ6OzlSnFf0YhsASuwBHkr63mS5+0l6HfHwKBj0kcLGPlcCIPvh
6w5yxbKWqqEXwYLfIMz4bJOBoOZkmJ+9+g7/TaDzVDh78yhByt7ZzOS1f/Lq
yWCzvSk9W/pemkwYQT16kkwdc2k0SBFCElxySuM+G9dapn+KZgttYI9q++/P
wNxguS8EbAqRvS9ndR0bCcPwoUiwzas+78+a/Gz1QOWCQvmxJknWNbXUTN4p
bv8QpExbFLsFW8DgEdJYN05/eGiySqYmz0wwM+5+um3WLvhh2bsT6aFiBuzm
LWXIZdRnJWtiVW+4pRhmSm/kShQE+vu3jXFpk1YrLqB4/2jxMhqx852Ja9tq
Kx/dWO9zEoNnU54Q2NLHeKUsALzbzLMxOXroGnSY/9KQOqsdN1qtWTvjRnXd
jY0HkwiPndJuQNRwirEzM4f+oMZx5CP1hUayvJqAANEsoZ4ZkD6DDzzwBE8k
0+w//hr50RiTQe+bYHBfWEyhovgBH6jG8C2CHmsOsMT9r9wH078YvpxVPDBb
3aJ2UBHLATJihTZt0DacR3VO47OVjwq+k9fmmtXSOBI5VN2fxlBGRmUk/ks2
TzEzLBonjDgiSq3BLJ+trIrMHPIGtZiUzyogCqIvKDc3j8Ou1YuxHk2oQlTZ
l6lPF8OKNgbkYjttUmeX8gKaiq7jJr+sMkGcGiXmYwKVsbiajjBSZRkCLbNm
anmUpVDF3Xw2Jz2z54gq/Il+KM53boTpiONBgp5tozvizCadY9leAokE3DmC
DpD4eWxnci7cLewJuYyAHDzs/4x35MXt+Uw8UdrQqxCG8nga1NgW6jDdv16L
GKJwxadeZ/PKaUAc+pbkmBw8Mk70CGWWIIBRZxIjm6gdu6A762OhIdsoFI1W
MCoDm5RmCUYMlp+rRJDwHRS51574gM8/srIKHUau1pcRn3poTu2UjEknaied
AE30bR1+I1SWJ3QnhwGUHf+Gc0xcZFmjyWBhMZdxgTn1iv077OJUeubWL4Lx
I3+eqXQVr4U89F7BLlheJ7VUZxMTha14cLsMAihywVpRZdWXaxIrfieLe95A
9/5ET2w7Yio0El7FVEierukYeqCovxzJi2oICtYRZyDKSLrNtraBe1Ma+Urr
A7KqdyPkFtWdwhoASwkwB5nhk6EH+PQrykhR5xiq6TuZ5QiNR82SjgPln9YP
aT4PL8MMSNgUfWl5CiefYDwYV2EcTZQ/gkW6ohOcjLqgcTs+pBW6Nrs0l2JY
I34m3dw08KuAjv8SIsrwQszM5WJG0Hf8trmBZd8mKeRiqNV13oKiiU0+KXNG
g0oUxjqyd89h+LJosIQdHggK76da3yd6e7AZCNpOnnxbf9+NtytKg23SWE5u
95tK1vL67FocQ4QND02kEdkDJKat+DGTMC88f2XgXhGZpelsb1HwvlQdRF7l
jWIj0mRJFYt18L7fONK5a4U7D/fkYPunGF9ZxJkb7mvxxuKkUMoMAjBVfNeA
Kl3rIRkd9TJ6F9LEP5ZxYtrvNznN80LEoUUS24500ot7/xFxzK5MSa87w1p5
RT3S/ov5FjfYelZqDayqv/MQBBdfAas1J0UFm+3UgFOqYaMpm2ngfuLaqst1
cec6qlSYpx4fSIfGtlMVV1dHwzXkfsInPn8rRJAkqVcnsDttCmz0Pk6bDzPP
GTj0kUuj0xrhth6mnzccqJeQ3QiY/GWnaJDLxD0JL5390jHqD65tBL027PqI
JFUHH1EE/uI4HrqQecs/HW0SFPrS+8k7r2mQpZEEzwcSAQHiV0Mz/JCS84Ld
hyEXgglYS4yONJNNxbCYbBv01Awwen4XelkB7FU4vYbsvefpq90Qm+nXcr0K
CVXk9s9lUlrv/F1aIQ9DvTP7F9B3IdQQk8kNq89vZ7H7ci2IbPRirJFn3Y8B
NbjbXFrWW8IXXNFcOljDtNnFUD8nzbWyOSKGymf/9wCnkPb3NS5MR+IlHNIB
FezSb2r1TSYfIIS267x4B4ge80iv/7q31njsDDRoxzAyAmSTQFksDQ8qQYeG
A6cgZ3phpogEuK77c5wAVb3/PDck8zi98Z6oZmRDlNKN6qVMwsh81MNMULkl
2Pi2v9aUVweY0jeuA8GWMazZDOytWBJKr+8RLd2c0hFMsOYLVel9/5iGGaNV
n3hg+MrAk4MqHyQZs7HPxRPaOAONKI+d9E4ALGY11zIAvC7BDQjCBEvjHqj8
LAS2dZaqsuSvWK2tZbziqkWbx1fiEt3Jt1C0MRNuKPwvZ4cY/EkEMYA8sGot
96ggBw2UrKc8dpezCAqboPsLcYAgVfnF/VIGbp3vpAOXl4czR3hBmv2qktj1
zKz9vaVyZWE+Vxbj0bFfyGthcorBU5IRI9mHFrxPRrZcDUSpITr6iR19/og8
3djvrZPSKSVRDp6FRaZbWKBUv8PqerHcJG3hymttpD7Tqfy7TrjutAASyRRM
Wh3hc0cTi83Kw6jAD9vuK+V8K4jBepHaNe91aU2Odr1RGm/+VIeMt7cnj3uM
fErzwILfa7GKH1K2syAq+F2qBKOUatnqAMchhW5fyKE3JiWCbarptggSpGSo
LoPuLZST+K5uySLvxPKnqQ5PmIi00hdetmVWxB9+tL9lzgjoGCyXRlvObgu9
ihH+A+VAVWboHRYHkyOsAS7ak/bcspvrRm7u7u1JzR4ez+Y1HTOMJ2laCcTZ
NLjBJzhV9snHUOdzyICo4jOhBS8WdmmHZKcobdXTUi8aL05mVcyH7Y0mbcAX
acCcmQCJklvw91K5C/VQZAUDXL/NTBlmYGn7FrMtXB27KL9XhtwUqTfCTaDP
50w8L43TWU3LI7OR9Nilb9cgJ5YAfC1Oz40o3N1Arn1rJ5XH99YpH9/Mg05B
2660a183opTbjnUff2xOAIJytoSOxlih1C9WyDGqqG9heGo7KDVPlYMaX56j
K5NnyC1TfgY5EI9u6j0WN1ZIKaD0GJownC5lWLE0nDRAQXw/uTUXUifNMECk
qjBgU3MlBa3vC3eVOP4p36aO7oTB08Pool22tF4M9aRGukJwq0xqHYPV54qY
H3wpI0nNKjagBILPJsu0s+JM9apvCXINJ4x13LBx/hjUaPKYbJU+26tj30zV
vri5e6lv8aAEmmwMIyJT5UrDniwSmJjgPCU08E3I7jdnGuEN46mTL5eTNrb5
eYVVFcTwfbDpf98LmZu4ECAHcwJJIpcH+jjhppkzmfgh8U4EPAYQM5G/QmwU
nDwW3fFpFhihNEhlPTK7iWYSYjIcq3mCvOHHna7BCwVM7h+Yg8VZ3RB4rLZ2
fdnpoqeaX9lUFaQOwkuMxKAwc9999p/bCgFdG9pZ9u3eDUI2babd7+qEy5JX
4OWC2M+iK33uq79K0w7f7fI8ADx0wj89gAaxOuEfbYL+/mdT2GfM3JMb03NL
NRSLv0IiA9Px6p3frDbf5Oy5GwOThKZqtZ5a8jekXEIHoWZ8urbmWXNH5Ch8
DIOJySsttKyok9YxxZLe2vgL5FT3v5jCkUCYY1jAhZ10slolvcNdbMgSOm5T
A1kkEyrvh77GPVeZE+3Qi4do4v6PsZdcXa6VbJ7v+hEK9ja32d+Ej1xMa8Fh
BHBvuFK56ete4zczfNF9GyNaRET4OVs0xRrc5d4LMMio5w/HD3obNX6QOErM
AeYmLLEj/xIgjpaWVbUdFqNNB90WfEc6mFYphSKjL7JdGtTiljfbKc/iJBuz
1D03OiOO8FFZ6QiCbNmMXrdqciafSac+i5IhvpsHZix9BBNE8pXUBklB0k4K
LYwXAjRWrTSFmUHz8F0XJtAbxF26Jnn2XpAlJh1VM6ZZs/cT0XXeEQKFnOGE
2mYhas4Rqi7xdJaEosmEOQm7XANL4V3Z8vw4TcTFREqM0z/XHVSWpsy798Wn
MU7++XC0BTv2QgFhn5tjWyKgxyBZfXlenodaaZTCXGHZhE4YFCcN2jiC5MTB
tstoNMuIu/MXz2wvu9uGZnSaCcjUFsSuykB1Guckr/0Th1pLLasvXByF94YN
DeDfaU6rd7DmI2uLJtsPqJiqcG9KEtIdnCSDkkcVRfdi6lsdsMkaavk91Bvb
fxYPWCO6wNbttFgHC5zr+aqFXHhufnmeUCBFYGCBsxuKXk5C4JqMPkp6MG4Z
JZsSUmPUBo1moAOWWNsYqeL8QcYOYh5/YfHd6tlq8ePuIH0kPSDSd3wFgZcd
5uGUtTWlTaN+YRctM6iUnP6/d6QpvbvVj5Fb4mJd69DRKM5Y7NMlKm/E1/yf
F6/oBRHCGBkm29z6dhG6+2+t1k92MqvNXB0laWY6Pxzh6eoCDHFQva42Bt4r
tz5KncRZfe2N8+U6KQ++DOr2LUVaatC3dtUH1jLkossF4es/INWdUsRbvlsz
lgm7aX6/MKrCcyP+WfNAsJkabtghjhll3mEburf/QDB6BmmiHR/GfT7hufbP
pE8B6jo5z0ABgAHoFWLpyaJZG3FOtmFskFqsriXesX1qyc8aIwJh51OA/Axe
CF39rZKIOHC1gxUqAuNPKlP4I8YYAdDZSh9spbihQKYWv5IS7RhygG5W3Q2f
ZTumsMRw/23o52s2aLqT1KgC5Y7qUhvmTBciW4kES9snvmgMaJkywgg1UQFr
6+GQUy7uUvOrc9iSePSucZ2ZEdPCfaVeH0t4+DY91L3JQXm+a9KokMZbq//r
I/Zs8Ih5r4ND099NmmARh3JvtBnbMgoJac793MTh/adshdOl+zvZYArmje2o
qrfZzKSUgLd0uB0+4Z9g8Q96H/YTca8dJNztx0nNZjDRkKZh3LLCQLemOtAP
sv/1WwD8fafIw05XF6weRQkyfjQ2ZathHLoWw/hxonhC0AX2m81dlleUEQNw
5GoTkTANE9iKgD0iRmO8KsZ6O04WzDc5dn493iHFxBXzjFSJhrphoRuJTyb3
n72fgX9aIWg4BXGzRKhLQP2Ju7pZmBKTTg9FtAtvDt9aEBZzKCPgQk8frkY8
jB/1ZDjbfodBC4e1zDFoGGl53+8eIrKSOftkVHZwmS0JXswJ31su/yzN0ZwU
OcxdwWDUWLry+9XdeyZLAQ3aIWEKKOjqOyfQUP+cpI1x8Uy0ck87yUUIJVTi
NZQNn6pRJxAsjYKe2MaelpyMhMwIHDnFLpRPYVG/GevenCvRgnuqPTSELDAl
s/O95NmcsUMJdpgh4/jLBfBh6faKiZukwV4RRnSb0RNzSi/T87psFLxiimwC
TbYzlpgZRihcu+D6gE6fvPSNGEmEe/dGGI0FWZb7ChcanV63f88MsjEAuxHk
YAxqCloOz4gVnLk77X6U0PC+nMj5S5NssEe8FohW1wg3cXldjGs+ejpptDR+
tE+E4g5Y1O0vXgqOhsMmohfrlSYn6ozyRfrhvoVhwkUQJf/A991DmNtr9l3z
jlymrTEg/sOYxJGTwIUDvm6KSwyEgmwR5tEXJ/AaDYIQlCvNt2h5vymTsoU2
0OkeYJwvtgronjNB4msRu372RiI1s2K7Ai4kuyLeASBIu1oIbgGLBDy5avQZ
TuEBMgNMLLhLkNSlxUSmohzbib1PgqDLWSuSWJr+lTpAwHhwmNRoEKcZWisG
6FRxFp2zdw9G98lrdE0wm8nBUxO5jTVp+RyPmYAZ5Mj6bIsX5akbjmtDEtYN
ff8HAQ2I+B+LBYVF7Ehz5c9pzsekXtz0xIMCmhIhlr4o6UnkGCfxYbN3wAhK
PDL0Hu+/xGqd2CXsSeoU7gaeFoMO4nAWig7KFJVvPlHZa4r6T6xAMnw96agS
QrgCQaho0YoMabDnXWe8StoSy2gsj6fszFe2fftGm9Osz2GhRz4XAfKRJMba
CfsQGUmn4k9DAkunwOWbQcNNhftvZeYnlh3J19yQ84TgJzc4u8Y/ALUwrBXL
O81c2yQ7dBHxQkayLJGHQVC/wUc8CfMqkjl39H5GLUGuHuiuxxq4C2nGmBdX
xQA7ig1Ci/uJhqweOu+YxubXBiNIcsRCx6KJ8U+u4QcffHYFZYgyTWXQEx1s
9pljLwC2jaPePF5UgAH2h+qlE9TmrU8L8PEpBkf3e41wPHE3n/d1Kv3mytCz
yl/8tkPQb2amIv5DnafeyFwIvoAPqk68EyEoX5EqVH3Kb9yhnJQIrq5vMyZg
uh4VPy+qy5mrBlngXL2f8dkTg+ZEWLGM4v8aQCL77esn7v7hoLvjxlxUz0yn
4/WI0/1gxqZovWVGIxK9OH7xARNw44YvmH9NsubQ819EXlFJucDrbEhIupxM
zfA0dwzKgbEAqS+8Q7yVx8Vv0nGn5U/nbH5Mh1EXGw+GpKRyIAgle3A/kndk
3Pq8l4ttURjZxFY+IpxM9ZMc5L+ce+KTE7Rjx8W+yJ2jS/jbKmp+tJgX/Sqh
tw5CorqHZB8/+gHYN3CwVYDVptWYU6h6A6nPZ8royR8PLO8tHcmZzM15A1ex
HbNt7XDcsuPUMRHzOQj/xURuL7aKhvw/e/Y4Vznb/xJUiSmIfTyGL/lAYm+g
ds1A/5iAAQkI1n48Q5Sm3dotQL+SdwnZacfF7IZePW2BXkRWotXZMSr7ffcv
Z5afi0T1Bf6MCWdu9IIV+UrhBWeyixBjdSaoLWHdOjaIp//ubsifn4vMgfRO
l/BlXPCr0nAuSCe0uCkqVP67rER16xzIVj1zYcPzcuk20aw7C19fYxyCDOD1
PGtFdhvSgr4L2JvLmjsWYXt0EsLhJnal7SdEJ8C2E06c4yMXIMKAgFWjAaNB
Y382RKgKwxVUL0Jl+mBHhwhaDXDwyNQ5b6DFj2WERY0IjW5vfP3MT4zLyMWC
ENHAixEPOmLMkuQE0f+4XcFTlaLHI//wIDCW4ALP+3eMVo0OleIoIRK/oXZk
QVdTz8Lj/ORTdFcI89pkMNeckcFnOOmQGUEmVNEDcU06Bl4jSQfo4Y2ckXEE
vCB6TsfGSEgNCxN5Lqz4E33Oow29ZlJ06FaHjQ/Luyuv3cgw5HTI98kPip1O
I1ecdu3JVhM6GNvAnelg8x1dDDKt376Y3UvV6zh1RBzyEVKQ8NrNhtGw9siW
iWzQYbmEQlv14ic5PBf+PHb7pHSoEhecjPIPv6pTYh/NpTUBFVvkrZYk2l5O
fFyPmw9b/RdU4eKF7Th7AVJM0uvoRuqcYgwPja/sZ9gpUQmNVNfDmoKzEesJ
1dLLeBUC7d/XsLbFSUUbGCMRmlvjQZZtH4p1vGqQFhyMfz4hL+FvwOhPZTiq
gDCORrywJsfhIUh2taNQOTcRx21GwCwXCT/3OBV/0GLuOy4f3QIKgSJx4Jya
rvnAdARHFNWOhpri65JHcX2txdNhMvaG0EDNRaOQXrLSTda326NIgxQ85YeA
6zXGQmk9oUyK+VDawxIH4EnJWx04X+2nNb+aFI8rbH9BDyMOWNgASHfoKHRE
75WUOV3fBPbdMS5gY5RC+EbpjlufEGVWiwFawZJP85ax2M5aHCyGWgoKt2zb
7A4so513bl0YlGVshRvshNKD3eGsb8vJ74LzHc0PcdotIgJQ5/epSsBDNfSf
aAAf9WY739fudWH7igQrAFRKY+A5YnPxwrzaleNe6/fv33w1I02v/aJ60wnY
1Bot2hypRk6rH7lV+VVXJdsfKVpgPGBDyTYxxbcZELSa27a7O5YMvLWxmkwU
if4mcMl8LNmJH4YT/FwAyx4jtKsV6Hvr1hclkDnjuEhoph4wvWSyp84uRqy2
t/M3vbIiPxWINA+bacBP/MKLn0S+9lMLUTrihJK3OnZ4MkSBL/UfiNt5/wKy
PBrT8q+RNekWYEcSNJ6kZ+pY/bCekO2YS6c4ifNPIKvTshFybioo2LOHcFab
pVGMNKF+sF7kCUL+WgB6F4Rqw5cBJUy4ugDsBKMffAAhOjOhm+5vzYpbm2EJ
0R3aeBgpHco3yp9lnY7zLlrPuJwtXrq3yhTH7RF6odQbY6jEsF8GyYNAZyP9
nvbyjPirpO+tOWN6sry/IqOqhJmq6leYnfuq0xpfPEeWfYmbGMabEH98JsDp
yamHzwvDXY3gSAbvRFzEYjYUNgc3DhnbYNmkCgPuRWpMeJ0o1220PT4Sg60b
qG6fXOmDVnWdhegEdViNkaRWkmoEt/YXBy72wIWKxhCkagxpj2H9kQh2XOqk
215KceEL28cP7kFuCipVY02ZCPkOXbhrmz+xdT72KuFaZDuV9gL5vZqWcNo/
0zngyDws/pm077mZpS9VrUffmnq0YpHcKa9qlZYiGZQwMqP1HpXFoZSSGkoJ
Ut7Y10155tbN/HFs6tKCVdh3uh5c6FlnfgRfbd0S+QgSeGTUddl3yLsNNuVj
HCJWj1c1+MzAVxaAACeVcsBLEyy6oOQfDA2cAfdev0r2eCpIakPlSKxNxIHH
jeZBmoOrtpRmcK755nhxUMucGx0Sd+erm70BR9RcWBif276PEE+IDMVnxlf9
FpXyqqC6EY9FCkEOAU0+GewLUi+ApDuAMInp1UamlOc7WaDq4+uL3SEebhz0
JxUK1+Y255l1wIsjb1aPnYd5x48Q4bg68JHvgOiNpGiseBtRAQqXXzpZqEMR
1g2SHvaZjiBfFLBfXnUhVTzZmYTZZbB8Iij8hwct0k4YhTgR9d8BCOg59oLR
qSPz69B+NdMlyr+Z7gA/zxsw4GxFjnmLyVlwLj+bhZbkZ281Cmt0kCq/rywx
Xqm9ogboxe0mGUazRX5QWvCkhAGG/GVxmzDGor6z5q0jE/smTFZsilpcZ5o1
D7ZIysG+hi9dvUNXVbwuDT4+Ncgdl0BaYiS7/1Ye7tBFUHleaot78YjsukhG
RuDImxQAk0bff0Qbp8dQMX7/SxkiewIRl0CAqlNiPD2QvIR1NG9EtX2mDHiQ
VwgszKpfiNZYnMsBKhVoZutelY4VE1mOd1F72xI4TsSmnOANhZ3tRYOPqA4d
6usjqpTNKvtFvJvBkn1/G9PPZ+MiFJxB0W/tW65vPwEIf7nsLUlHx1hztbQb
cBed3C8miH+S48VpC6Arz/pis4qFd7+nasYFG26m2Au+o6jTtqPm7tBpO5VU
df6m7K1rIxyIclYD6ICGSFP8+ph8hMAcnBD6JR3HV6tKamGxjmOxN4CC8N3n
usARCjdKjeMf8hO+cw9mOT5waKzL1vgUwJ2BpFmdpKs33E2ZaBphJUJDIHxg
KMvFLvqNf5UzQATmTJhRBqcvGBaGQ4XdId0Z2n9iDxUJI5lG2+dCryavXTEG
dvvg51uD+hWh2O1N0QdZYfXqr96Fwxipqe99PwbNI9PZ4WxqhHN5V7i9gGLA
mUxFa1VjBpbPO5EsDkZ0Cu/PlHP+gIeCsDC73qj8hsl9H8OhLMYtkKkYDPQJ
/MNjgMKyWKVgM20O0nWJRElovimMz4skuSIYZGMYWMLH2C5pUeSBudYneoaR
GkHgF+eTcAxBWPB/cYshWCZbcFqQWM/ivg3t2KgcIWAMh3Vry9kxGICkl48F
/IoiuFMXSimxB89kqoqwFCd+V2ZrRr7DKzmN0sI+TXZQ6fAGzjow/1jWTNtE
l6cXGQJRhqB6TIAoxjBcKHspTJNAmcTNgVoOKgPz/pOKtas9Geh2ntrWU6AG
LdINOrBPyGqNirrALEVJdqluKASJ1iMo8x/XEIFx6poya3JmUcdyPMufoOZ2
GIKp/B+66f6PViXC2ZmJBE6SuDxUaVzPlhe4oZgfwVYDJap2MJtOMm7k0jpi
/TXymrqkjgeG9Bjn88LOcIenCkiBWqxIhfNUR9XpzkRaKdJULxrcar7VO5EN
YtGEoPg6Lid3RIRbGm9+37WApexQw7XNWRHCtL2IbM2E6OquoZj9wY5e11dc
MKKkW0k5v4R88PPSDfVVTJjq9T/tGO5rklWtCs6hSwlqRPAKBszOcRUuIMS8
Fojfz6/hJdywCb4Or60U3cK9hNGp2BJ1RH0p5a2u7xqu7U0lAoAS4re65jIw
0qdN/F5ugmXvSesebXFNyMSGn9AgLfUqHJKRsqdUV4yqcun0wBGz8LRg7GCG
+hWluTfVEbYnWxsozCYuA2jnYQC/kt7mCTZwjBrwv12xX+itY78OH1P1Abhf
SNqkIRrjB3YIt7qk1nQXGXmj1slGBROBmM/CV7gYXZY/z1oEBitZrXCiXXc9
AsJ5rGEbp6RwkT0T0IT5oyJ6uBMWnvw6CLW16kmJWsdxVBQICyaSQs2Byhyi
zfiPKCcz1i3klq0kU/UfHB6ULCvg4kan/+UisvNdM47bw4WT+GS4nXbdipHG
EKmf0Vo5RLXxAh1pBDlJipt+yitskSjyjyVrysSqQZzvA4FwWFHs/0p8PGhu
qitiNwVqfhpAQ8+gIB1vRjBlVeKpzO/sE+GcxGFgsaiOuKTritazHMjZ6Opa
WVa03WR7wIV/P8SaBB8b3/KyO+nxGVC1QqsQPskraZIUtztPWI4UGxr8fTyK
s9hsPDFZtZNNBqUt3mrJxf59RYEhKEILCnGIveI/1Yj4nchjCiQr8Lo38jMX
/W7zqaB5+rfl0sEAcW2MK8vF/dmwloSk5fCuyXeGiXOzMcXFdYEExPZ+/5IH
QK0jSDYzjtbd8KikXI0nkm9ct1vMTdzEZLAy/9Oi7FNJTtDMPcANhGzjV7ql
jU702/+LoNESHXBD41TdtdnSorqOtaguYq/xa98lBSA3DdIG2k5TjignvQhj
G9LIBm22EFnBbVNEd+/8eNWSm9bUbNGDzjN7Xb0yHxGH39IpnJsFfCOb6q8L
J9tmrSjVkZx/Qrl9xsle/DG35fo8eyTw2NS2YNfejyFcbQqeXuU8y6xiw6BM
/tYig1GKCQ+KwfsEEUJDcCgivlP6LF/MoDAiCohXEAQb8AP5DOGV6JgkZp17
MY5evqKU81Gh+vl5FATn4Oqg83rPqtcjh6W0e6E/8NLpL8xdc2eBvP7pY08s
27PvOy8DTkKX+7U/gcby0PuR4UJwc5it2AGJPc5c+492BRpqCl2K9jPm7loU
PQf7pMmL2xAlkxS4eKkStM5lkw491hVSepOEvAeAC6fpxZ0A+cYwJ1lGqn//
V4D/4eDprXBukINWJSPUZkmq+eqPMDjmiHf883wm6kiVqs+oRpKJCGyCTPe7
Dk7EVunXukTZVS22Ro0g8iO2K+QMEoaN+nMP88Ys/5W5xv4pbK62b0j16y0E
kFC3naQ2VfMEWX9i8vKXKRPIhEYp6V64lRdAyg5SZFtt+r9CRbb8xphAe4At
JfJKb24jiZb0iMoh2Ehs3NAqvgJjhQYwJDX6boBvgvgAa5S2lH0u7DFobv2L
kGKIwV/eEAce+zemD+4NTGv6bNiKASzYQBlNbOeiiyMP4tuSH9iD23ryeB4A
0dhIrpgt4gYqUaadz7zJNj1P4/bhH4DSyhQVEd1VE9f37MooNjnwbATEMSvC
NdhplUhcjM398DzU3yVKob9ZSbv2J+dpubP+jl5mJMuUf3OzI/tpP9b0Y0cv
V80OiFQ5if7uGo9llVh7s89eNEj3KjbK7HBLYMhaHZ69Jv04aFSb0AbRKZT1
Z8wpljJdeZCOKrZT/uAhcRIGgsvpD2rMGIFEbvae4dGCEWXBEfrLEQp4pJUP
6YNl8hD3O04jQGgSAS+X4TLSVl4IpKRx5rJCzd9YPk/4uqyMOs7KYXvujEXe
/k7OBn3kc31rsGArHZ7HjxOPpSnk+mHu6ppGEd+rqJB7+xohgLhpCvtd8fMv
F/zFySHhzIiqfXqY7My8fV+rIH1Ge4o4z1Ok+LB8Zqztc5fIHgUupX7JcYyB
8bAlOiI7a3c6ZLwyeH29lO8Dcdx/0a+XOBuDZyoAuZhcznIH2sAGyGgm1EYN
e3tL0p3dpLmqXqjnxCR6HkKctIZi/t6FAtE5/NBlMs06TtKcAVPPtOTi5I8b
YzaPBS/HW+Gt7XTQV2lnnoct+su01Alrc/0apBlM5khgM+X+szehgZllxQ6y
j1j7ev4GTkt/S9aiYa7jQ3q4OCTJWcWw/pVi6IXjjjS84gl/Lr78Z/Pkjdj+
fjwbohp/jKplXNHwJyjaVVF2SxIn9zu2ZFdOu9bao/RSCCCXxn4p1hp+f3nL
VlX0xhaBBg9zA6kMUbmB8HVs8EcgEizgFUhJW1as/jOSffdfu/9O0A7IpxyU
GFC6aB3cUEMhqE/y01TYlHtdy2d71XjFTXNgtCs3EhnL6gySPiSPTdF+nVU5
WCPY+WOnkxxi0Wn3E3XBvmmGPpYBtjXluSFr8AvW+VubFWPI2NNa0D0edB+H
vlVHd3gduV2CEP4CwW+5aKnoJMTA/J3ikMcogs/NFSUpzd44nUxsisSRhT0y
cUvSjEFbysczTmcC7SRLCvfnqc0q3e+CvFDC4S+xEvELyDHMZV0YaGpVaxXx
7vXwyYII4zzM8fysDQKtr38PP1rjuyNtuq2CO8rJcodt9DlI/T/kGDaG3jmf
Yjp51MPOp9G/R1Zy4Kl7QGBtz/15DZGcFA3wi4nHtuTqSJed+ILo4j9GgDam
uJswj3md7mkiy+GIgRObAVayaqcLVebtTofVDPt2QRKF4c/t0fWqx7y6mEKE
jDkHYnp2DcbB910dZoWHL6C/AqoNMLi4TY6oS+a6XvZFyG/nGrX/7PwvcQzc
vU+HnXorwPPf7Ki6n7c+CKVBQ3EArMapq4roq/pVbtJ21oil/k3K3zZluugH
8okumb+LtbdhyHmM0PhtvOmGdvN6teUMdoqyb80xGfei49JXqn8RRrqf6xax
RMZOj+ysJwf2BOmktkafMhJ69N0ZkpUX3TjuHtI2yFw4iCvT+HxjiWQgzOsX
7+qRM7nWAqYyGaSL/Eb9WvRZBDomiEeDaVWYSMgGKav6fiX9uFO5pYPqphJX
2b83FI9KRX9fjUrovkHN1gtkmJnfJiJd8Bx4+OmE/dPxUKLs0l8o1/4UpMFV
A0NCsl0F7g+v3DzbIEjFNEQMs73PDSd79ZJGdy9C7f1X9VqOj3ff7qUsD2P8
wsXYcD7XGqQIpJZ1mw391Kqbw3H30MK01fOqvgx50MPaWIfYk5fRNVE36qZW
WYLCp07qIc4C9HCw1YOs9dLROtnzG6/QybsRU/Km60UkqVrkOwPiM2WBKUkB
krHoJSRExBUT3dARCADtphY0GYTvuBbR+a53nm1DCqSIKNKPT1zgGha3yruv
1HBhtOTo0Z77M1lLf1sJBB1zDj66Dyiz7ZWlwEARc+oU4vJOP5EZvvUQRAEk
eTJIPneiFMueZ9mK07MF+pQqYMocsNYMMi33g/wZUhlLJSZsRLPA4JrkTnM4
k8qceJBe26uIAueLlTTTVEIqm2+OrsSR5LGCSbeaLTr1o1FqD+mnEvAo5VWn
D+yHjLKh1o6bH+qsOZYii9XIyt23znUClX6tUSXgRcrCNOFk4HvfOGQkvP3s
7YITYunYvt3q2Vix9xM6BpYilDP6O4jAg1ZZu0zT2tsIfY/KuApxY2VBhS7S
Ok/CE4TXjk5PuSXdGLpugdnQLX32oxuNIQiogAR88v85d53M3ojhS8cgQ8Ta
H61ATDqCEcCEIQWDmzp300/m/XmfxquAbfHecQLKtts+dE7hqTtlf+tUBzAT
yi6iYGMVzvg1bxtieEdhj6+EsMFLrsmo1SleWK09ZVF+sAt+l+UKz4idZPjG
zqVojUp/CA+Aw9eDwwIlKj4arl3SrXOKb4ri+tzQMBhvt+4EjwZDY72SQHu/
yweK2WFTyPwCMSLIyd+UhXeLoXIfmlX6KX9FZ3YFlKbr14AYFXFAosXPb08c
ESu1GmQQKhF/zDoV+QC/1drJSEAbKyynJ9QrxfdbG/nLNhw9xwZLgCLmYjfG
jFnVRO1AQQuA2rGvMQJPIHFdU3Czu8JOFAK5rYxSaNDA4oHMUn3pbcvEaC1D
uusFOADMGhX8XWCL4QXXywFc8beKdZ8RkV9qwgfnaSEFjTOeNAV+62exsNVM
+K+1de8qfnMgGBIdtNZlgG2oBcnW71D6YIbgcO8GM1CEOsaeOnbd7+Gx+TIZ
roA1msB+jGWiU0oNLbKVkuwE5E5e6+qKMv/s4qa0OIrVnPR7fL5ZRzTt6gRU
/4gauz40csXne/H3RYZVN0sFWxm2IUsmPoc0+OtS0CaAjHc1KcwW6X3QhzAk
Fh3Ezsi+yqwNnSJghWWoNrf5+4ngT/0zux/WuQl12BhyoVbQhLk2AWH8LR16
RSmSNJFt72qMuhd5zDefHEcyiYMydqGPktnERrwWaNMQwPiIAvHX6pcpyUEo
mSGlD+5Tj5Zaeh4uFvMJXWXqQHgMFHbGkS+2LNK11852Mkk5vTCSVhMjWEg1
d/4c3c7boZNBq5RKMZbAe5Q2vx+HFWZJd87Z1ROSdRTyPBvIQ/dmQxf4ekof
ZxYkl+SLequ0ulk6t5ak/kc/4g0PFI1JaGns/MiqBMu4pmhqWWDm7kpc+ez7
+ZjMlYSvhaYCHd7zkqIcpsgBRs3JEYjnxbVrZMMoDNWz1wTmJSNbswmKX7xY
N+I4nkr//duJ6bu6gcRJ31YLjvz4Lf6MxCM+lGs4VEb4uxDvy3O1mJdjj7u3
WlVhMYoySh9M7l+WluHjwtPqd7CN23ePqthur30TEIlE0DWFTicGw+2kZV9x
U7gV/eJM+WN38f77sJSxV5shsmP/5CQl04KAXuSqqfwCyonkfa1uLDFmmiKg
jBsCFmGhKA+GaTuDbCuUbn+ey5qaHo3Wf35LRRiMfXd1l//HubnW5SVlB01P
/nUq8KxwGmQRHc8DQsHXU8UzOJfXIb7nj21OcHAmd68ICYDTv7/Z5nfB2T7v
A2g9KzNwPRryYJKDGYV7t4UBT1Vlv/9bDIRO8kbF6cbMrqQ7AJIKIZoNsDW2
7NqUYyX3OyshvVHTY5fuO7x7FPmFX/iog6CEQn6fdQTVr45EPeASnhyd1QRQ
aZ+4GaYJcZBVeKpRoLuw3EBL0k0AAhmsGxO32bJEkHxlqZJg/CMGJf7D/JxZ
RdEpfyCVel0/f1T/xj7aGTFtYW9Brrhfsa/t4SK7Jnnb4vY8xvipbk13V838
RkVrnC4y97nEkCylopCudNqVCznPSMZCsArNEbFmohL82QoDMtyrdy9xafjC
1M2OtTzy+O3JkBLODf5WCbkQI3o9l4CM3lxhFjBlQR5jAy0TFQEcNXdRstG/
d12d7PUlkTQQETMhXwnohELEHScy9MEzc59wCZy4qdOhTG2/ztAZ9JmFQ6/y
ZUEplUaSKGQVogrXD3USFQDkuGB8KUJSyJzB1Fh67yoUb0t8/3bZwEEXVH4l
p4GiDVcb/2+SPEMfUywZlYgsWCG2pq++DSsQUh1t4qIXIb65B/K7vUVTR1m3
w3ujDY6YSQ23BF2Iit3NBUh/LQiTp5adqmisE0ygQlIQmUiF3RTC28nqX3wD
24iidR22O8oJ3oAQcLbRJxof/GZ0q483qEI0Vw2E/EungevihtgmLcVG/NiK
YcOmRSAlYJg7HcXWP86pqnjwteDVyijVRxFSzCPBfc8B0KGjvy7MoqVSbqMX
BrZq/GsUvkgFfISBKGIqCRzU7XXVqfYi5vSjo84e0a3PCwH86Azv9cTdNpU+
fLhvWNp9TOK7dEd2114JFP1UPbLgqMncw+qU9x2QlHRBSW1QLxlBmedG2bwx
6RzL5XGadwHUWDfYhtIy45kLNc6u1P0c7h8Bfzo8sEWwksbO2KumPhIRw3jb
u7iLRvAF0iItnDYNyoryzf2FSRcmwW3ox1RtAMsYTmKVa+Sb3Tt2z4JmKq7z
IuVpcINTc5AMbwCVaWtFl0LfRgc6dB5fN55UXa/knKd/Y74BLwtVYK76phPz
roTmJXWr/wXHTC1V1mzdS/xlmOddEPxLpQDWtLB48e75xC4ay0aVEjvCHmo8
d7ePV98zqFlB4MvRTh5wp8h42KAeXEMINwi3lANRRxTaDQfmfXPBH7Bffxsz
rYTrmRtLSfpU7AMPGK0uhVPFcrYVNWWn+r8TB6+uB0nvVRT9O/YoHXLNWXNW
BG18IiBqbaJp21+6zrOgAfv1qXn/1nun4vQPIz9odTvEigEcHrV3NXy93uWG
ihPSNMYaeWdrN7IhbP5+ZMyLMuB3hCl/C5Elp1EUPWJoCg/kwFPcBzHScyDn
blsBthfps1gpYVcv2u2rt7y/sCBbl84t9T3r3mZHTnTzdsDTm1HOUVQcrXZ+
EJLkU90o9w5+OWf7aDEVE6gX0XYGl91TWImZwaITnC5hcTZ9zbbY6HvCfM41
XH4yqrxTxKkTztvWnM+SDJZHpdm/zt33LOdWpy29fRGCpXU+XRL+LUw0+ZBq
TuKVK35AhQ43QWMLcC7RH8fBUoy+IlqfnMtbxfZh9UvHnVR5nTqeH8LtninS
HlA2/qFW1m/mRm9YO+ml1UG/p2NuwDt7hGv11X5ULdJETqsuG8CZS1cVSJiD
TbHi1LMOyVze+qQyfNpJDX+XzuOL8CYKWm1ZHFOSz/UAtS8P0ZTApucgGAGI
iKyf6umPWe8iS8Y0RdT3Kh+EmsaqzsC3m9E2nyVEe8nIurEC2KwUwAStsq70
MTrnOalpvCj4ripQEpA4s2YA+gq9Vlhza1sAHEc95cKTO1WuhjL7jifPd0nN
DApzaOUYC++AXVVik26jzSAL+pjQppjCUSlbBREEsEJe1p6enoL4TNWf9hA5
RgRMW9tTd+qS4+FswqVNZu9MJBbJhIZo56N3BwE15Ob4W/5oe4w2kbKC9ZC9
VIfAaFL74V4wG4/paII9duECIDP3t7sF76toy8ZCtGrvNCfuMs++t4gU8Wg/
ukQgjd4XK7oEfPpakHk1HHti/7f6jkHDa08VV8o5tAKjD+uKyz4qoPlfw6bA
mYKEmcWGlYDNF5rCJ28wtonZXAjFWA86k5BGEkvsaDGpvTLKObAH6FVB7X+3
ndNoWh9/QmXgbElSZ2QuknabZAavV6e56Pen/STGcn+YsNwNiTTLvlntyx3d
zjRv4Nb/B0X6rDZRqYo8UkHAy1kRMlf1CdXDk9JUZLoXCWffgI24u11v0+QQ
4n8IcR14bc/PrgPINw+oBcgJJUOE6kA+1Riqm/CMYrLnY0+RfCc/Tf6TLUQW
2P72AmD/fubfMl8kO7bGrnekOiAE0TJPHjUO49eNK9DVvN0HvD1Leandeyfz
KwIBoUKlaSh9IAlZ86+Trrqgeapg0RrWNjWjwRCxIVVmtY5IlaCb70366dRe
Jz7eVrdirIoonPHzD7A62fO2X7OXtRpzT8A/P6qA2aiL6QrmUmXEf5j5Chpw
Mz+eiR8nQBdIj0ZrHN7AO62AtpuLRAKQ5nK01U4yte3xavjwg5lccAXTavvR
N9N+WjK6RczoEMTrBu2df+6md5x1yWl3+W4rCBDZRb4DPiQffJJSvLdOaOyh
iZbC+KotVGEtg1rQhSn9936ufXbfJtJPNefgxUVKnNnembHIlGhnBSWfS68x
l3kEC7dnzkXC0rUF41CQigxXjNrLFWSc8BEDnUcLxRwRb4cnAz5NnP9sHssY
ymF7XMkpdIkWTTakcL1oa89iM+2SqQwiXHUjwpWuJZ9gX9MGzP47hAke93wd
j0ULqoShnvgtMlxMZXxtC9XwxtZ4JseaYMVunmBTItSyEO6/t/zQ+uarJBOc
+zqlDviGeMDO+AYlw8wMlh7+HB5kPx8OMpL6Pa6heIhcXfRNZeIuTOT3U8nn
BZ1lq9zCSb/Y+kMcht4WTNr1k4TLL+g10ahOKS8SfT/X5nHk9JCO19RwqaIk
Zm6qgrUe3gap6I8qwtaT9KjZduhJ0A/bslLjevS2sxhQkNHGxTl1pbWmP9nh
dydYFCN163wyzEbXgSquQOTaWX8ZtCzX9f4S96OmF9zdzrJqz+qohFi1LeFO
ZXcrxk+lEJ6VnHrEKmkQFEMOIpHpsWYffQEfd6zH2YOyPO2IGb/eSgFujQVH
B0WiD43VGOeVVSZlivW7lIzrd3U0WLvyp+uNYh7dNEydLoCR6jw2JN9ldBcz
HUDhZXbFTCUmdUOtcmCVyNZGlcHaJtKwgSO01LegVlLdRqTIqhgUYvEAWGFV
scnoiI4lvqrdrYtjcbTd6ziIXiLY/MVouQLZpZo9/XaVVIUJeywIPU4fJaZ7
4tWm37iDfQcqrDALkGeBXTYZ53X/HmmTeEr45BvmDhRiF582YecFFgWGro/D
8xy+H2FQwMF6JlRQbhW+b7ek+ILRCks8wy62pAk7/fnHxoM6xHVsznLFpquz
e0xfIf8tf2DePeaqM8CE/g+ga27u1yZVlHjS3DpkA00IKrZF3r/ZKqGHGkGZ
/1srLvVIYMsFEZJrqF4dhWoOeQc+gBBQjQYs1sZULjDPwMZ3azY6sOd/aStd
FBRmnobp1U+vEqglvBTF61cuAOTwSUKoxnCICrnJpU1Yd+hrq3f+fE8BfOc5
fP+ZO/wqPBfrB4MTA/Db8MGns8RFuxmp9/p5NQK82VJt4YP0o0QsDg4EZjJ0
hOHx9l1N3p++82lSUWQFgI6uoY8gUKTRZuKf2phpgkWUlQQ4/RtcoXNW2LrK
fPcdSPs8qoTRiinjUXYNuJ3BRAARYpR9J9mItjyV+e8CCDC8uNapMudPOEVc
C0bERRFIhCRgiskZferJuIFzXSU7b6A85n7+atVij09aIznQRJ55/bysKICJ
nyB3XpzC39I+NT2HgtJRLicE6uT7tN9a8mCpYETOoH2mbbmFTtjzhXAB09Z5
wQjeVSxUdYaV+OuZ9OxWBA6Y88SVBfyP9oPRhx739WmRoUuvcK+VLrpjJ7Xe
7DMuHz7Rdb8Y1zsN5AN6LIWyBQC2PXl060xLewjeGR91PDVkMO7XmJTrdcXv
EE+KPetbCfRWWYJF1AXjq3feMtiB3pI9M6ruRNNpeItvajAJkO54FPYexyLF
uChTRRadRLQoMsSzXI+M+CjtvHUIQ3TxdB0IWn2Xsgzu4kIW3q445WUOVl4Q
Gv75/sf6vattS+8ttOV5QCEMs8B5uzg3a3Dajpd7LzSvP8DRMHfR7FRWkUny
5KR9ewImlJIFc8EdokpOc/XYn+koihJTHkontPhjXzvos6gt2C+Jgm6eZHMy
Lleb3DDB40qZvdcJx3xDTQ7/9HEvyJG4IfaGpM18oOcuTTuPFwWfUK2tWseY
8ha++s9typF1f+NjTzL710yHiDE6rf4vfzXc1qUlWRzrJrJZqL0ra4Dl/jhr
UbchRgB4tkRkOl4k8mPmIzin+IzAxO06qdcBKwW8UhWglw1hypqQ1Uz2r9CK
BNSxNaDoXvCccmmKRB0HUzhEFls3OACnn9qBYoVk4MZGE+ugnSIdL6R8vUlN
eqZCPgYM/lpq71F2i2qQeREmM7tpbD4hR3IKpUTIVjLu4GW7kaQBYzFO5yBG
NUUlT4fGi3Bg8QxCJxNUYA1QSqOIOlWzIeptwLuZQBCISizDejGJx6XlLwwM
Mr9fPMTtFR70xa0sN1pFdNG9Dv0IKk51yqru1KczsdM189ikv/8TXi9R1ixc
3z0Lyqrmbgp3E5nnmBdIRbvSXI12wGNErkKOsHUkkZFwq5K3BOLEnhDsApj9
Q+EHQgss3kOPBjI6S6I8CTQJoo6ZuyszDzufd7Z7BIaeAisQ/5NzwcGfllIR
CxEDmPWA1SIqaJZigTDNAADxDRgNtkoDWj1g6DdN1bNEEujNjEjBEDUldw5q
Z0zNRv3dyPN1OIlqi6SN3KHdc5F6RDfu7G/pTi5CZ4cWOsMNTBZJREk9wBu/
cLacx+1fpIFogQO3X25ssIKcphi7/MwdkRiZO73y4u9baADCADhGRwjIJ+ei
gPk/5NhWAgbVJsMhZh2vMHV9R2MnjOl8f4+4t/TuRQLUqgbq+osj6PWit5fE
OAo9cCXKyMTRpkfiagnBFUbDgWjlnpgDxs8M6pFPbeMegObE6NkzZtN4xF4N
pmWsx86JePkFTZoyVfIpgFpfZ05ERJtLox3acbpycBpkxCTEpxEzXXKmSYn/
RGOalXowrZ1wXo5dURU8eK5kLejUrsfE87xrgGtl7gm504Orxw7DZJ3sZ4IV
5Tsok8Fuy22JfvzKCLK6uoWMVkb/SRBvYGgFN6guU7CCaNdRqQr1hqslNrR8
GXY5Uf9zg57nfJz8vhlCe6cMSgzmDuPV++O5A+w/rUHrT/WIdqfkG5wzcsLg
+AoRy6HQKFZC06wx8j8PfN4hlGJ+/LizHTr55REoQdBrb3fHWL0FJpxAb5Vw
tVeGZ8sZ9x7HfdCRah6t95A92FoJcPGaMVAFerLwo4wwAZ+QALuS4BtsKLa/
GqS+U36krtYm55s3rPsFyiCv3iEWmw1ynoUcOUgtE2N4b7qN4nF+VBXWcczl
Uk94yKElswhdBIyhbZ8G4hX0TdySQbgjdIQHrCXN3eFowOJp2GXu3ciBig9B
ZqhdLgmsR8EzWvpOx+4USSz40yadBcumETKVvlQLB270R0PR2mJW7eAnn+Pk
4E8F1Byalqz43kU0R5U/i0LfJYZXIUMk3jT5PsEFD+EbkygWnwd4xFvDmj7e
yXhFrXict0sD9ikOygQY/qj58SvJbg3pxasqIQjuhK7PWxSDiclSh+vnnJhQ
z2Asccy14biqnDtVwmaxchTeBKdwZraGFr3q+m0eb61xCc7FViJiE+uLwjmU
Qy8PkDmtavZ33K59u01fsPDKLZswtqvbqmNm48bPhD/HQI/0r9CVum4SY4Xl
GKAkT1ywzlPixaCeBTbbiZ2oETso7przqv5kwRSSK+93/LDr5CszA4FquvDi
F3vuax3q/xIgX8IfMCZVmJ5lSGc/TV0cKCspE4hKjH7gGo5Bc8tY6tel/Z5d
hp60220e78z2JfpR/G35ZsqBVoD5teLp4mrHnERF155KJ3wZOZIld3qOLxyk
+27u+AYwKMb0rxdeMUyQ7FBjFts4+3WK7mOh7YQOroyFvRhkfs4L2qP64Kw/
DkA2VFDCPHJ6wLeNm7RtBDK0iZyzheI6yXKWgXPzQls41zGkaDwaZ77hUm6Q
RtTnXxkSGwOJ453bPIyolemwnGTQQudVaAUuy8cEb98uwoT++QSP4EYdGCj3
Xd0YloI/guS4WhOgmI4UR7+pZl21XBChAM9E0nwyXtjV5X/IEl3HK1GypUGH
DLb0ITO0o1WHY1sbS07c2TjRP7iBQkqD/tUexXCeRAwcEy7wyuLMZglWRtu0
PZv1+X9/3+iZjOFGTIptor6guZ4PIKqiUsPtWpYFAwpqPHj/GUk27KOESjkb
UjGkQcS9XX8i0dFiY+m6rGhHNV0xVzrgpEl3e1Fv+2PZFfO/jtWMc9XytJb7
fOB5PSdyRsp/tWjvfhVLLvtRcPSx3BMo+C9zr7v7q2mVhZSI22iSz3gJ2OSS
R6MpgHeVL/WvqqQ8BLEabooiSkHiJ0YAOVdeyqfe0h1yhERTMbNHmiDfTe5q
ixArBr+yAQEDPt1dTMYw7201PeOIgAnmOTcfo2401LMRQ0PAAm93+3AZgvTr
Q6Ii5dPlETR0KasolWLO8d111P0nHmEnke/VT30p0oMFuJq99Aj9ZUkCJq5K
siVXG0DDlHC+WADG0f/5WQlhS+MVhUtSCPOXsaokN89Fbw+yXF1InSAkQj81
peJk+LAUNiGsNsVTD/t+ypTPdbC5MI/yQb2F2xj5lSCL9qWe9NeeFXg9cSAA
8SAbLwskO9ARE+IRabsmKaW7kvgbMlmosMSi3j/T249Vj6J0AeWWuB6IdB1x
pjOy2RaTKmCqh7Sa3ecPrUf+Rmf6GnEGwlc+7e/vHYOqki1vKA7W+uzNqxWO
5Oh3BMUoXZp+oBpOsDSRbepXwHOVL9BSaXEiAZWeAeuDj2evepMku8BonUky
hGgSi/+1v2+okSaRm0nDeMrOuVCWiVSgprPywctKWwJikCmUkx+DR+oSpaPa
wgUpJgH32ciFuTZptjc8VP32ltozyzbX6fEk5H+urLquYAtncmCF/VawMU2M
Q6YHDD+leR77fZe6Q5YnUZe27vhWOhDQb9iN00PGsWR72cfcca3ehu+ZMeZl
A3fykAoum1XW0O51Vv52+hSHhzemnYJSsVFINtI8QMGZBPMk+ZXL0aiPbqEJ
q86jEyl7yfAxDK4rPZ7gXbNhp32leRXzr4oL5s+hJFZBKuJGlAg/hLibHFOR
13LIN13vnC6E1hahHJK5cEmyz1rjOd+DPvuncCEZMBqJoctqE241LAmMojgy
XeqD6x2EKF6IIa2D1swmonT5GezoLYBqiY45byRYH9rFWDws1J/FGzYIRtEb
ZuaanFenLd2AJHUgDia+fFHRYEHgLrmILzChxkhYlrlT7YeaudcQ/UqjWliN
GKw1bOyuLTXhgcHwml2xKfo4fh7RUcJQyNjSOOoes0H1DehhCn1uMZG/IPQT
QlUHKtLNTLu8qO6qnINUHjUIJNnF+1HumGYB1wkx3U7a+6mRjpdZ2t2ssZoZ
EZ54VCEa1ywWY51IaPHogIY6KzvdyPdMWN2qwSnsXKPTiAjjuAdiDkD33gQu
mHfDGSl8XJTvXbhQsiLkeC6oj97pCDQ/J0bf5X2TdF0K3ZJPadHBTYih9aYW
NsRvlpW2U3XliJnAAGXbmF4damwdIIvSGXiQjBfvK7DTC9ICsNTl8H9fwtu4
jP/DrDVXKVKMZ263Dle9qioZdnZF1gittzZ8r/quG7edEb6j2uRfDomw8LBK
XGGKCHIQUBw3lkaDYZ6p9zLtVxxtpWOClNnJdp+wdq1x+/u3Xjqvt2jS8DHp
eFACCb6jycNRU4i2rs6mUCcofAhEYi0Ryqm3YyQpVeP5c92NKv+A3H1hhTlS
RQ+WgRsnHoSq1GpuVRaDKIUwmIWPZgDOrR5xbDPLYOI3qusiqBKGVJ9j+OHM
4lTvBSuWtzjRh5lw/u5m4fqL2qkul8jV2prhidM3qwAFrw2BJsN+mxuG99dy
kHgxmFBgICoacXHD50AYi4sou4YTJYMhzF90nYD/m7iQgDJqBqgRPPXC3vIP
CUdnRNnuhO4HA7dOnNxuc6U6Ktr9UfBlJJbMqHfWESRWWqjxFNSsInvDJJ0+
FRYOrWkENHy8FiuDLp2Sk85CHVpzSzH6AIWbvOTDzY5BhCxx+1r7uQvXvT3W
4+a1aqXR690t2DUrI0P/IEWCMefNPKb4RAGyb6NrjKs+NgeoVZaZhvF/t9YL
VZV+I8BDHM8mJZ9vVcECV6FJu+rQ6teLAXl6UT1SIUre7FKci6zWYCTML6id
P0hW/veOKaigU5fTOaYYXer1tww3/I+6WrXCH5zCrKmeZxidFO1z+AoFUZsg
0wNdkTN1Ykq+DD7CoLd18JTNMpv14XJNNu7s/A6Q7CtJDRwHkV2Gel9GUPYQ
58pRcq9KFhVyknXq/kpc8xZ0ONksQWm8zscOMmpUx8+FZ7d49aCdirZ53dU1
kxuSxqmyKsds9X6xHKr67ZtTNSByirU/u2Q/vsScV7w7QVzOVMSzqeryMWtu
IITH//NrYOav+bqLGDYh9EaUPnrfVCMkQSfBYAdrTbUXLOuQb+FfNXDZYZZi
ysD514Gbj9mOc8oZuTrxHrVMRZZ1lOcR+1JztTdgCMq6d/5SPhLkKqFVJb3u
wqmlO2Vmpl6/EkLPpGIs4I8TfJZM7UtICLKlJXoodFo4dr+rbzXAY6wVwH/S
g1fmlSoHGBOshV1OG54Vm0TcmdrAyzxkKU1k2JbqkkDSqXiI1p9+9IiFwQdZ
aJrB4qXIkpQZTEcswzr3Rwjky2MjkU93p01kfAUHQP5g2n1rKSLzOUmuVayh
tb23nSnL0CFSKUnZ045bsnRAYNZ9A7V1Je9n5n+9QLXqlxVChwjh4rk3b5GM
0Jjrb+s1d0RxTZyglB61obv9t2HoKTUOMM2j+iSLXeJlgm+/8NrzX7uQYHoh
9cSsV28M4p2qC/JCRyFJ+ngvP03i6x5kjNRtAHzJ/xcaV1rJ0YiavVd55txp
YI0zQecl2SjpXR+fZrwBWChsn6f0UsjfiwNzSfqYVdLJjZNnJXUBHtGctYUU
/+53sjJArBT/J11vOIzcCWlaxc6z1sll19e/2fmANInRlILdoRslvyB+n9u/
uZp8jk4JFKKzL3fazf6sICuMBhjiEJSYoIu8yBqCTKCskdznesOzDbQRIWX8
Zjlxz+Hrcw1gd1vVnAdAFil/O8o6V53MFs8jzgrUbxKi6FjGCOTZH5xGc6NI
MxEvxh7hX+y7ZJxb+97bokHrM/t9idZmpX8j7Zr7MWhg5ju6Hkn5DPATQgM0
Kk77SZHJWDM8GAa42NO24fsRZWNCMPkqAcODSWFM8sdiTHzQZtS2TqoSibkH
+dSQwBo1/nBt8i//LRR2+XKBPX1XSa6zr4rsayY96ZXdDT20KAUxXlN6P8y2
A9TKpDDz4ioP7uPN86eeRlif4QvIoTE7nRf+n+amPY6ALp6BfRQw19/PNO3X
QIFRDX+HXfajTCONiHeMAZcO06VEI4jfWXWt04MrewbxXgcHv1ctJv1YUVjs
tKIsT8tMuejMmhS0H7tLhMAg0P02hKDCXUFRhFQ1KBqE5isu6kOvRmtfHeKg
g9cSk7FPyn6bGUMp7wXt7IxOGkH+wOEOengmsRnhm0wf4ztRpg+hEbo+Cah7
9aNO8uJFYCyqA4xO8kb2LPtt3cuTWaUsHTb2TrgrHHmMRgVYLgUCe+jEixg6
SOFsgsozscJmHVn+SmzNCac+XG8TTr7yBKdMu0iR14pyz2hrBZ2VkIKxNJHg
VZjfA0CFI2POnG6RMjRpg3MCRZiJM0fb7f8vQ7Jvui8z3XmZZ0fJ0jvFpmHG
9bWlmki6HVghgrPQPZEoPrHgs9Y4+UaE0b7zsPS87Us0z0kkgaWac743MaNG
+PjWxxbTUB5+zI0QdZM9HNtyfFjNNYxbv1RrCbvJyDarhmAGe1cDQww1jLZY
Zcl+G+LWxHTxZnFQAjIKtRWp6oqIAfzyu+4q4mlE+zrPxrP1sZWR26k9tCWe
NhtBqENyLkVwFZ66u2xcFcM52QEaqRmyZzr0J85vehHC6vRYQGn6Me7oKBm7
PZp9Aulhziw37fQfA/z3vigKV65QzyKUaukhaY/9ejVRoVFnzkM/TI8Fszt+
/qKqZEWFP1NaksS1SUAv226GcnQ7l30A2F59SHD2vklq5bpqLVYeLtNaRfzn
hYxVFrDMbWVeBa5ao6ozMpXoQABitarj0eBjSL1lG0SnsOfvYnAI+Yt5vEj8
NF1qC/QPDFt/jdirgpAL+BbmN4x3/iv+8AMYjO0F2us5TJyche1YE6dXhq3U
KHsnXiuVcrO4Gta9BSS0ZDd1QmHX579zDDauluyLEibE7F9FjtnBKBKBJl4R
0S6g7+505p8Ga2Jcz4E3DlS0wDQ8Rq4iKQVlM3+NI3hiea83NVsM9cszQPk0
e8oGPmUmgsV9kIv+VcakM24uzW6T3TJGJ+G/oDXIuvVIgP0fHwIwQEznsmoY
8qKVbsqPTo/oJdMdqb8VzdeyNiFEZlR/yqiO4i5vBzAA1V2eAJV1vlmaA2pA
0Ay/RNyAPXrco5rhbHNscoz0//pmmccWDFHw2JAs23DWAa7mIhrQgY4o6bKU
sNup5oEztaHyHySrJDL/PbW8pxDkfwt4G9BlpC9YO1p2eQ6v8+Dnib1cjPif
Lj8L2gS1hCp5M5/T76JjazGeeovccptruNHCUu95G8leH1O3oNl5M1MI3RaI
iegNb4RtmjxeMjLCc6sxffL9V9fBdR1HEEfQ6lsWyHmUoZBhac77QqR9tbxr
F+qqoHin9lfW+FWncTTk1yAJ5WVTE5Y8ZhEcSnTFUdTH/IiYKKC0DG1Spsvy
V/a1aR9C/7SBBasu41ftW+1AfUC/AojsaTo+XsZaY3VMR1JTYprFQs2kNVXp
vewiGG2iQerTRSCmjtOWiGSbsocta50c7FAuL3ZQWCGMH/9+f2h3zDjAV66h
Du/fShVP+DMYSKE+SnOOzVTNHC0UbXYyGu3QiWFc16jGOKoD1imFoO2O2cob
svtSJSxQoNbS0x0iLSKhYjto+0R4GqRVSNKYZFQZzWgp17PntFVKaGILq6zh
JSAzF7L18jFX+lpcxt1Zv2iBXAmv7BC+8iasHoGCz6jKzBIkuDXN0fJ/sA/t
MQqYPpR9fWpOg8HbH/dnNnqrl/zjNWBJ2toJce0jOW13zxk5EE8IOGKZ1ccq
4RIGuoz21KA3npV78aMSgg6zrMe/zfyYjR5Uw7tgCUUOlgTp3Th0Ll+iXqYc
GIQQLWeYe10aA2cqSEy2lVIJKnlBep3uCvSYGgDoYcM6Bl2LMdyNKS4BRbWF
MGfiQt7tzTyimyBpAuSevxNd07Fsp6Jr6yliKoB0sLBGD+t2p2eeb2AyjCR4
lkp7uxBpuvAiQNZkaPEyxZhEmZ2e6W++Wl3ELsTaQyGjEW8oDCNvDDA6v01z
vfTUkWU5F9dRW/nHAHXl/Mzztp/EUJDHyCuQ3xXeqoH5uEFpU/G18uZTKeow
uzbp6o8MZ1NhQQDj+nWRDw6LvmHndgwJdkn8pKgLt02rpt3e8mYqbRsD4YFO
cxCWPDM98BRWGgEhNhemyq7KZcsewJEU2SrfzJlTsbtC6HmBpeMvxTbUwUmb
Mj8uRsJCKin7A+glSobiZApVxMEjPaWyuFl5RpupAHBxNq3iQ+91OAto3IpU
mxg3TYUzcQ/4FWggDgzwdi/seLycbmg6WfoTm1TKO9XGhgz1l2osNkjPjxRl
kaTfhQKtSpVKs3Qw2UjwaTdeukZdpQNFJHP4VoNg4/IwKgeY4KcG5OZQSdns
nZhQz5sxandUu6LM6n71ALjCPp+K/8vsRinfKxMHxdjjgi2igKAqfI88iSVO
tcvwdAG+Kuj0zFuvlG/LAjcSoujUvN3D4vfaBTRSKDgWr8nA6jqqBJOEYPk7
alKN7yr4AphdDF7wcfCDY2ugXmGmSRuEo/+r9jjSJdBSATWUBG9bIn29qGJ/
4mTiCtJKgFU+eDXYGxSgrimRh6BLaFuTOtUhCaxp+4FBxii0C04wov2gkx3b
ltcJn9sNNmQeIFTya9Pnpi/88JT+T0ggye+Ip1e/JRa51htdZwdjVFqVux8s
gqfdEzWncbfLKTDqacRr13zvdSamqmSqIclTJxkfzbzUJBhm71P8y4oQdYzk
gKMfkluK3iBZExrZno61v2GD5cuzDr84HAaFwMDlgocETQQgAtL/xsplImIK
yZlVb4t5oViWFUFll9ZvAFiDwYIjuMcSQyWRdd7ZKmBXqGyilwtUts2/Eh6k
M9gmhkXA5w2PMd1yYLEPN9mJ2CXOs6ArNduWOLJsrFD7q5IlPkJt02bOaWWb
PKdGlPT4h4eYxfZrCog+w+5UHVkmmjms40mGgvzzUjpSXd1J8+gyYcWBD5Z2
jPd1oaa7jDyhaY5eeMUiDbBGj6QaVSls6QnT7m3zn07fWpoUI62y+QwmMTtG
KQoXHsSf6tpIjBvzHaGn+pcaQ6TBa+qX7yoRt1kWIjYHXkCsyHskLpZkks1H
C1aYLCuLZc4W4q39NPg9UomZnZKL+6nRjxxYrrSu1C/xw5CcqkVAuj5QhcHt
HxH9mdzdIVuy4BjgyEvysu1mdDOi5cCr1997AUuX4cZo+WKtC+5PQxUEtZoI
P20oqVdHPkkMalWquvX9oSKni2YInuF8lbWlBlAmKpuc2XdbNmERw8E3HCF0
eqdYN2cpIQYhaVwCVrCDTxQfQ3OWjt03BA6rDbJkpEQhxN5EJGEWo5NPZU3v
8E8skCY2+46xivFAjf+UwIgNqx7rtlXMDmEe7FoLgGbt19SKWBuoaQVF4Pzt
XyJb/vbhrw48qASuSztdpfhGN1O9eSMH2Y4wUbo19jd0dtU/BFRSsHLt6kpH
8F3atl1pRzaU5oK+EEh6SCicZQ3R4uIgS09C1fysspQsm+V7QRL8kZ2YVeEs
w5quo4Y1o7QPabxeeUgtKkEGTREPpPR+mn3e+ymEzaDRq/yvePzRokgneEWM
QX+Y3Mj4jSEhUp5GX/wBwPFURcIsIO9Dkx29MlwfzBNUlT/UVOjTCEn8dZK+
54CueV1Px0+VfpZKGVL0bY24w/RmnKNOF+qfw7yhoRtPhBQvdSXLUNJalgbN
WJjOdWrA/FCxKTe2Ix3CMdQDUhczYEQUp5Cy8VsN1DQDGFsExfqiCqJl2aer
f/D1hFTTfBNC3z71TtZYuB+II36mo2XcuRBDbKqd9i86eSVzGn27NWm8Obj4
z0RSjlse8zCKT/XYIWU2YHdsRk3SvONoeNr52d4FdR1M+FpgvfdDzE2w5v7+
GbRVvBFdd7j4fJwkLn6hm+xVwqrM9iyw1XGIAS5gF29e5ukk/tQxZItIT79P
4NTYUFvbb+8u4tHzNGQ/E7GZiNU4bFmTn/dUnpLtFxvpt75vffS9PccV04yB
Fr8ziBstt/2IWlkR1c+sxxP4Li97xoYFIv+nGqdqi+Q5XTFv8MtBv+eye5lb
sOjeJaanT7iSTK9yVKqmDb0OkWX3MNp7DAuhJoDapDRk+umX/TPZzlLfGMY0
8FYgOMeK5yd5eFBcFd2joPwKIBpdKQVnS90x/T36eph+sWv0zlX5XtKCEaQo
mP8ydUM5M93X01/gmkC+aJvLp7xHgCf/KsGluOGN4UIOmDYotj0ou51BfrH4
xJCeiHQzgNczGTRmm8P4chktMtmX3Z454TDc0UDvtAqG0heG9V0KK5zukNqh
M6fRcguezzGAloA5xxSYGAEsPnPQV1A58rKXlNU2Szcnb40Zva5FzUIsVsIl
s4PwdLGfQ7QPm6NypXQs98EQHSHbII6agWVTXXMLUpUgkEWqbrLZp2p8xUTC
br3LmS8bKfUL7/VqtBzig0xjGriqqBW+CBkqyT51V+X4VvB8Xrt29u481QsK
VveRhYWXNkzjY47eL7X7ESb+Bw2Js/cTKzT7hUha+0pk/wS0SN/ntUAiJI60
zrZkJNhQIFjpNYud6lH6g4UbhKJAEX7z5UOOftBnV3B9uITn/UwrzVUyLS9p
IEwMG7KBvLC1jjv7NvgJjN++iR/bBqKIPzYXlBorB1H5r31ES1UI4078b8CF
WLNibc0sPLYVNrGEyFP9+SFz1Tg8aHuW8C3QXE/VApEWxlHl45ldu1qhwOrO
3I5Gw5f0X26yjsLyL5uutDHkz81qinnODAt/IBNsV4Qk9WXmFDbxO9SMvJEp
r8yVhI39Q/AMkEaWQKS4leEpECqhYU76lapfihnH4bIwjaOj2Y58l/4jmx+t
u37WJc4rpmzF9rM4NZ9voxOa+E5+F5Xy0WwWG4J21TZzdSm5o54uNBe2NFW1
PbWizWkPcvjH6IGyD9jN0KF18qYNFffz5w00NR2knLO9NOVmRMkn+pFBLckz
Jx5J+B+0x6yglAzXc7wHqMapTUGsDIwcv6ZmV8qAWotm7mfG5wFom3pCWTeh
2HvYghE8zJk6tbrgsblc/wgfDSM7p99JhbjpWhVPZpVKkBCgJa0LZXYge9Df
AWINk9F17F4H8A+rPu/EzOwLIvyNwGK/4zwxe/LatFzng9+NvPA6QsGxjrHn
n8rJhs1MFpdrsDT99jh5wVPfrG+sGkWGdYZiQQ4Y9wd+ZNO/n2QbTV7UjHBQ
Cbrk/8OlJjNmFdHmtiDMuqEpoPPSH6igI6AVA6i4XyLXkDboTy4liZOOPixx
g+bJxxu1Nl6ODfoE35Pd17BzwKiOPj50dGXhQVgbtCVpZEdZ4cTFXInhsYiJ
mUW8BbnXVzhtzbESNY2LT/EgXI54jkVXbfFU/duZ8Pw+knwMvFlV6hNoyRNc
3vSj+fXjWKYXQQJTjHo0oCxpomcCmsM96qZ+WBPCdHQDdAd62ZdAoUSqyiby
IoPrN6rVAjDhpvgKwpkicpM/T1Ab/bAc3zDFVUSeSzULckORIwfNBi+YB40T
6kAVtiKm0oCp0gA2ggJ049nDA8dK0fMObm0FK7Lz6WZCKuliZ2cq3Xtr0+48
FSkFlOwB96TfXNV1nKzJup4/KX8dsT2ysIwK05iDbHiuRtcPwqnQsJMuyxMP
6iATdQYmg7fNr6utMBOqIbv03yj+vXydm9FkBlpJWJ9+OHJ+KmTqkUTvldK8
pqQq5dk5bFw+wd9MJSHOEKjkcS8ywvNvxrDxJ0qusD9sBFq1sXQsLm1cDFlU
K0HxO5bWM2cJJBlQHe8mfaKPcYfoG+9TD2RPNq9fn5QPD+uryYN5F4A9h3Wa
KuP3cIzd1lad66lInyqA6sIdnxcn2ZVz0h8oWHOVKpu7wMv4ZGb3gjcPOAH6
0wqQ8j27tr/QkYngiPHT+c10xkNWsy/U4Ron595VFWtLzs12hL8p6y0QY0DU
G09UeNT7/nZc4W7epKX3QQKzRIlzCrpzZpJs3cjMHdQxncZpNBVqkGki+3sO
2OlC2pE1DlgvMbQ7iSjybyan7Xv/+tm5vAvbepZ0c6ke/2v+RiouwCHhQFOp
NK/+EiFZ96LGc/K4B/rhC+bnOqmG7nhZHcgKGxVD/yVAcv9q6AeNbzLNl/VD
ssLZn4PQ4Wqi6TF5qJJy3WZ+CMBTtBRNrcicaFppfrVdD++lOgHPwgOnhW3H
p2U8MUeLNdZRvHilS5Vxzu6mWNprrAoL5iDUz0vZEu2hoYD1ITe8ABhl8TL+
Oih57HkifmgcIC3ZKSXYCk9oWZQbaYuR4dtw+1JpIXx2PvIhlvb6YJi3+M9N
OmsNT3EeO8Rk4lq+siW+BmVMn5OzFdCVreoRASBI6qLmQ1R+OUDj1Rr7lCyH
C48UCNJh9WTTQeewQJZ/jSG5obG87RydofR8wUhkKUl/q+wDpysTiHGBsK8+
ZEf4cqTwp9Yp9edxmeHOzhayt4IEUHg6fCN68rkdg89rYnsqsNduBvssghYe
jSRwPI1k3QYH/TazkIgFVzGbObiixP12DaPcAV5W+/IjpfdNnFl3pobYJdHq
2TAlxdIR+Nqfoe7bpJWAvBkwqtHBcZixQcxEWMHvCAhOxUJCfX/NKofbRzsP
Ys2h6ki/WUiQ98rV1G/vvcec+18yKTA1yQwbfrtOXVg0hw+V3ETVf1zbk7Hv
WuRUTmA0DPAqLilVN5LRCYR8FBIwWGbcA7RAX6YvcKuPB/jK8lqV1ak6QZFA
V3MnD5qKAeuhyNUEXXuatfwBX7XPrIqps4YgqLqEJLqqMoRmxtKbrnk8vJ+F
E+gc6kJ3XN982E8KmQ29N1vmCitbNdfWLM/MM0Jf+FrRXeddFPKtxFlaxIMR
613/eQg1QanCInf+nyrI/ujTj9I9fY1vRZM/j1VUvr79qHj2EJDxowSya/UW
O3KCATHwBscCI68ptN7hZujPzCXwInHLvRWazyqBx1SSIinUvRpwh9njtqVM
VNLQ9vyPNEqRRVwYELhzC580hRYEGU41Cylr96RjZsmu1+e23bCMS9yzpnra
IXSQZMEs+kemqnsFRgx3zUnKPAQU8lC0YUr/1BIpcg5OnzoLFq3UJa3+maR4
0IiTDNpREVAbaPdJprxirYPXRFofu2SLG2OJVKQ3sqioEygfD1Qi2VFuAlb2
dlua1DDhyHPeGadie9Ybapb6PIRsDMxLCU/zaFgDODckVYgEIJmXWK2UHFJm
jTWCRI5mXHCY60OFoEwUqo7xLLzwJStTbIUPrhvTNekpeFVOEfOPPJrt/GRk
5rctk7CcVVjezHSK9kGQjfv15DPWqkHVd6s1C2rPUtVQ3ZfaK7tN8jVFwbDg
W86lpKZwxEj0VE6tNrJ1Epo+dE2DzwUVH6xjP8LaB6doCjb36+WKzfCTLh8s
HQA7FSnW9JUPQnZTEepZkOiRjRw/cSbT7D0Y7MRxBtnMotOvsqbzKBuzGFou
LsuMdUikyIvVIZkmM+oPN31UMUtb6o+I0u/pxqeTmSO11j6UxPEX7SMMlzPy
Aj8C0+ySie2vv7FR6lAif3iidpe48TCnvfZhlaze8zlqbOoDUHEg1V/NT37K
QwDcxwgYdSa1vTEYAuXgPhPMt4e1nzjzvE28KM13m/2BZyNfRFI95ccuAZhA
DeFOfo0zxDwabn/dvmednJs7brJmT7x+QSHsuqN5pB7mCR9QmRMUFeibuVJd
KvzzbocMupSWnq8ya9O2acsfdKJNXyIRrRSsAOi++3IiRpHY+GZ3f9kBjfn/
Y0i7aw/yUdYh4r4/Hv5sEc/iD4ETSECCJgJHh8zuyoB0k3MPAr+NG8CINbrE
G9jYF/Llxr6ONgkqcQKOmfgYHDkIC4nM3b9UZxSrHCzoOvyWvPhqDf/foo7K
5oTKFbydZuauwUe6qfDaAYpP/LBJ0EJCnGWCEC/p90iVViiBzth7LyGcyT4e
ScOAc1Ca5xGj+/413OINtP1Ed65YkMFo0GPq2euBJMAbn1e42gimV4RWvZPN
+YEIH8xpQHHRxDSDfiK/nm8RAN3L16mqChzfOrzq6KABG6ij6M/n7lZaieUg
fy4WgHXP1HrKDoGSe0Jj2GLRoTX4fo7uYRZ4VdKLPdSHA9QxgAnuyKPYR14s
InwYW2FnAZJKrXqt2buJqKRTBWIJczVqpfqqDqAxwPJ2QrGjtTkAw19Bcd5U
UhvoOHgDbfsTQOTEssF1VsVk63lYrH2oLigNYSYTFIXoI5R7vU+unLMtHUou
86WmrMd95Crb76jMypV32lveL05pwPpqHh1ipVP6/fKIVJ/oUdJZBr9RYbqJ
zfgKjxpcQvlC5gb1cF0mNxKNCyxK7VKsQEnA4drNQETRpzUvAlp7mEWeiAYn
d8GBXsJc3yu4SsNQJIT6rgolwwlZmGFXyxi4MJSGQqnTkpy6Ztk9nFZGlDp0
LFqmc95cbVTtVuXgLTB/cFDNDV1pmzJX6Bcq9Obkiox7pZrIQcfemAbFaUbp
aW7IpzCII2MRZOJFqcswJDACm+0lG2AtXFD1rkyhEO4m16pq1dsbB5jxBU34
E7jCs9DuWaNSuXiL9s7NuN55QlgJeQ4/UHB1xkVQJFr/F2njdMnGrrzhx4q8
ysttl8Wa1mmCjb+tFvXrn+bThdctFO77lvozSorYIfYdb92Y6U3Euf/NbUDA
qAoLbJEYuweJosNAhFnnvTHGL0lvK+B2sDdX4ab+/KLvF1KcDCon5ZEmMtSk
JRp6Oki+MsAwI1pzpWIoi6ToHsw9h28MOli63kTj7mizLjaaDdIbEXH6AOn8
UIEh76zbqT0ymv4BFgSbEpo2aP83CCk15u0Q2H1xraCDtAPOP0J8zwFn1nXI
Z1DwiGUZWiU+CRJOWwpuLwEiCS3icwqA7tALp/YBClzb3Z8JH7u+imy2aAYt
TqxEIz18fFF2ar135P1fUot2NaH+9GleXL0g0kf6iGLFpkkfGZuFElovTOcP
iJHoAxK+H3Xy80SKbFFrYJxdmWyODhnLkWJdrOz2rTbLNqUXGscf90Apnx99
GAheoSRiYnVfP4k2avSDUI+7IC4rocxmUkUjtn2ku+bzLJZmFZWOd65yoQS5
WqWmSjbmyicKZXAaULmpb3Y3qK0zQ9Vvcf4wreun3KeNYOvLGL+0fz7I3GbU
VAXTWa2sdODWpjDHHJubM6qUNHWt1E32FnwlmJ8pEc25tuqCNZvV1n9XGpPt
IMS26uecOho5rXxEFKHa2X+Ws54dlE4Uxu7t15Rlct32R3Evi24STLwHyjRF
dAFvBExn2rBsjml15peHaiXybzZy2jLDifH809GGSs2Kuikht1I+e9pB5u8a
v6LRVEDpzMIyseo5rW+3QyYItXjFdDN5+j/DuQOfkdOHhyMR5BRTFPOgqEiH
oXUJjq7gH4wANBwH1dM8wSg4IUP0dvoV40UMBt6t3QGB+n4sjsoqB8KfX3a0
LJzTOIrSRcAX6hQeLlHpM+Eq/rCG5yMz4A+SOwOyHbigdR5unXIhLgDjUdfb
Z0yr8fFH/N6ofEm2eFCq3THsX5m4N/Pmdrw39Ws9ew4zV50gAmJdJHJMTklp
/d2JlmT7O88OMT3qYIKNYeyg2cZ9TMycwrzPueLFZFw7j/5IRv2AQQsaJ9HC
DKlXSnJXthwOpxp7SWxGDecbbCDBwen7Myv2L4ztaur3z2eyqdW4k9PuvONq
/ABT/GRVB88iwTF0IEoYGmsYkgFkHPiBRaaoEDQngnLfrcwZTQ6bQHU0EBnY
7YzIbkxTH38m3fu47sItg0gmzgA+NEKNHzqcNWdPIBqijj8keBzrmMbmepuA
Fyj+VqaBlu3FEuuvUHD2SaeEM2EeGMQ06FYG2MiSP6CQLK2IzKGP4TgH5S+U
5yIZeEpYTLNNvn+NOb2vbrP9OCWOf0t2XSvcWCDAALF1BeIS/dfx58ZBWaNy
zDfRpKs53n5japvP8dn3TOXoHXT9+aB1XVmaUiAn//UAzbtMh5KwpKgYD0bV
HgyPJh5rqsIrFSaHdMh3t0dGmSh/bm6uDRKK1/Af4103r+633Oc+MlKzvSFs
mSULBcUb2Jj93lq1xBFhO8QmBBq41deD7uhbSwWwXzGnbOZ+NwyfIjF64kgv
oEFxAgZcX+K7QZieGfEX4ORNTPEz/gt+Wim6PNMPoJ/tGOEORx0g6JOHnHGb
9nU5tL+YSxj59PLfWsSn0fhBwYAoiM+Ue+5G+e4PdjidKzGk8QQQlg24i/PV
/7JiU538atoLbpQVPA5ujBr41GNMoMG+FJsxYHQeURBvzw5GI49iit7a8NJ1
g/UKgFkA6Ud2DuLzSPYiXMz5Ly0JcrWGlwjPEzrGbK1e+w7+fF31FNIUWN4Q
jYkVMUThawmHhLcXcRJ6UwEqO9Z6ArgLFof5IXHK/FMvCgkmwTHNqzo1nAEx
CtzgaeiNsZtIWKSvkf+bAz9I0tlq89y69oiEJQuG2H/rGJ79LnrgDnZ7DkY4
7Gceu/AF65mrfN7toqaC0YOZp5n4vCH4uWQ3It9XSFrbHkjk9m+RkSgrxjnC
wDFrApwqdO68FSXVhulfzd8VTmfPOyb3MNzAqolP322y1rc6RvjxDWHObr2i
tWQfQd9u7iyrYpC8ZJ2U5e1nDvsoa8OXZvve3rlpaddVNqXOpqVUg5xnEkTj
46WeuO6BVb3d6umfG/OCMf1Mdz2ytMmuvq3fuSb5XgtGUUGE4/kay/hyTvTw
qMC4blEv+NYFJSxH7kVnqusv00xX7OgyPVwsK75QAQa4TLCJxIqGu59mi84+
/0kzEr3IrksRlm6KIfSuJwyqRfDpDh0brxNe09elX+sVh/IykOG1XCh4gx98
OK/cmeAXj1YjvSyBEM02nXOR0+VLOy8a7P7guIjCA1PDs67X/J7dWjfm0/XZ
DcG7DRfa25w7Vyx0XqfGSdD5J2I4Dk0NZfHyOqXh9Q25uk+BuAS6W9dBN1Wo
B0DV7+IQokxanuodKS+NCzskG9VyiglEm0fwm6CluH7NNb4lMkLTp80XGImK
MRzVBuywJsVRYzljmCpY/Hwu7TM63oVn0UzUPHvFbZXC7Pl/Xo1XRheG4L/u
nOuXGsdv56UfBDQ0KPr3sIbysB5Mppb07tcfHbbRPY//JhFdM4JHjwF4hq+k
qAO/JJPlKavuTdTuc/NcWm7jkJXlfpAqzImMwr7nKY5jU8tyP5EIVqheFYXM
aHhftBzXeVN5QcALKCRgJozQb2EbA92uKDMeJA4ToisACH1AW4tbZbp2k55j
3ScATrrgnSX7HhQ6S2rfP0BiLIW5TCkmqOVut4MsRUao5ew2dFMNYgwc1IDT
OlcApeg1Jy4wmuBXwbCfsxsdG9ywI2T+/FjA/zjKASp3X2lZPnfWX/TSmewV
S73G5byyLppIuAqzr/i4Cb12z3sG4SEiT1fu9u/5LIxVJcBOXt+lbjaQafs9
LAIBSzpYpz71FS4kuOMdR29pmduuWIpOkADBRCKpI0r8zZmhpoDgVnoa4McN
gPmuwvc+vB4RVpwmsDRc8gwd5goebnMWg/4qy6RyJEoQh6ANQgTADbCIGbei
qzUWvTXXnscc9F3P9dQ3/PywH6ncqjaPuhv76rb5O/G8ZxdfpAKigVfe0vHF
ChtVSNCihqMoOqtBt1GUJ0TJhmN9a2+jX4KDoyk/z/5DbZ7DAH2DnOf8evkc
AnHZuaUDK86mH9jJBotmEz71F539q4/1+RiS4QxjKjoJVloQrlSxz1x1SDXL
BeSDYq6YSsIyMC6BxBb2tBU3KXYypsLqvaAHfiMGXsrhTtORyGcd/F4hsOyj
T+EVYaxS+tVeUc/AO4JHAKw4Zew5Sc9+oaAF4GPqia0wbVshPeviJKBc3aB8
EGVT97Vpi0tISBkaf4F3x33w5yYdWbj1hW7HRbUqyvjiQ+fuVs1eVCJuKhPc
rkzxUTCoaS2uHCg+8pxRaiCyT5v+n94mWd6e6KN44hP7khhKeRqugr05xV6D
vDnq8YnA2ceFiFJzXOHOrhnqPVTCtT7wOe2zPnZ6SRgkj/NX4aVLROQrF4m6
yx6sumy4onx17EVLB1V5F2y+FT2tkEOSs4UhqxIVMh5XdSAvTRZjLiMAKSMx
DIhAFinjcRS90VMojyW7hvugI9T9LfjayZo64yxpbN2/voNb4G9qE5O9j/vj
oeqLvp7uWz9Adf1XTfp6E7WQK0HQ1TSWTREsG7PfxV1vCI2QxrLULohyeyN3
QHqupPalXDJgWnlwhso83K9Aoqa6e4UiMAQuJRVSmWhzYxaiT/wkhyvop5Ql
7ibyQQaH4Aj4IvuXO69yKMX2oYEBQW7W1/MXYOOsDBCU5DYMzlZNWuhl9rjt
9lA3WxvF5l1Gny+5+kYtuAFwSclZCF7DwFOPhPReggKrzxFCTTtsew8T8knP
Qad05yYfmsQO3fHLvTe0Ntw0NhHvRncZGMfd6FZahcpakKDWAJoXsifjS+Z/
BJtk4oz0GfakVwZ4SFtl/yJkzRLvhCa7Q2er/ipWm8vD4Lgc1DoB+8aSMNmW
BayNB1q5khptPhR5D9xXnklYw3Z0QO8FrjtviuMf2HpXhGqhhzNV8LvkVlmT
gsIjoMJ//Ktgjy5GDnGoofydETJ4LA2mGRWeasdQpR6GX3vCrsLH1614khxw
TcER0GfJIEFInQ3I2OHiV607Mx9M/m1b1PBsmuXCjYcZzKurZQYUy4z8sYqm
4TGPzX/gR1Hc5ETR3vxvY0C3eeZOkz3dy5ctCKynuml/mYILSoNWDxP07r3h
UAlCb0I6jz9lNKtYpbSim9Gi8Lg6G70UtXDsumI1t8elEp65bdiFAgED2w/k
lF0whHbvU39F3iCDDNPE7YwM+HEf7WhWozPhp+ttBNsHIFk5ckU8/i/i0I6j
RtngAj8gS2ELSkPDulkcsFf/9f9tl0wRXmKC68oyIpcvqcfOQtq/LFumI7zu
V2M08Aix2W4CB0dd2hSuJ2scTNilwCmYVhuHkfiktrhQy7gEIdVYVbjM4q0H
FpRx/M6YXsD7gGzGcq7ZOCRVVylXMhnAFGPw97x4vRlNcRe3/unVjGrTmzLv
rcS2nFPYL/eQYl1HjejxJIzcxryzi/l+g23SuqF9nBg3kGDMmTqZXm2aG/ax
NgC9pGPhN3xqpcP0UaLDjlhxqIW6ntFALenVxU61G0IDuzE/h1GcamY+23wE
7nWixuyLTo/6NOJxGPkfK6VM5mxU5GIilv9FapLDWPByHh2dOAgKgK7R0yAH
JKGPphXCicPN80Lzp7AZ49rOUmdMOYfOIblYMQ5fj/xSfyJbwShOJcXdv6yf
42qjVRuueLgXbRpc/VfOqLLZp6ai9m19GeLUtyePkkcEVXeC2poMbmjYgTGU
Jek8Y22qnNu2FNYXGaVIv8oRAON5IdNeV93Sctpv0ypA+D9CrGCJqfd7eBDK
msH2/hhkSC9Oq9we+dv+GidSRYhKftXrkQ/dDOz5hWywzBRHqMIOGHnv+uek
FVt9vfOhBOP7tbf/LPDqIaKiTEPxn6OCPEL38TYjAPte7bO+P5ayRNbnIbnO
7sp/yvdnWaSmCk7AWFNO2kLaDV8ZwsytmDpTPx4029J9KLCEW/jJdCZ0/q1x
IhFVfCZBaLlvWqqk6bFet45QcF/nKqbxub6RJAv5wkzfTJvxrJCKfFAG08pi
nKy1NB/8pprQVWKFNWwFAK96Z7sQ47Ad9TRHO5wuGPQcwYpGW8L4FsI+QJB1
j+QxLcuBFz7J+ea/HenctBWQDq7TOiTWlYw2JhsbhyYFxZh06s8IFcNESqiu
n+gDfTqKhdG6BwtRiUpFkbCg3jTD2H7RXRegZf1RPOz8sBJ9FJkMOJw/YltL
DMHhYHo6wfosGiTgya/hoNCWC9SzdBE6j4BrQ0ZBdNvc5Z4fMpWXlUuBWDxY
Jy7d45VibwTvb3nl/+FYjFg+CgDSVjQPC+zas2znTxLMTv/3zoxNsNfzJc1f
tk2+Fj6Sg8mZ8cqTWRSiXi3hReOV9UqudfLAItdJ2ELIUPQMg1gnQzKyqbOB
LDFJpj+bAu68lIni25Cm/evzhdR23DxCa8S1htpxK07NpQQij7nd3OYJC3B7
JHstorTXDE8rPdwVp/XKdchodt2e0/DlRh6MstJu/yBdShxRW3ZOebooX/D0
fVQYLuDTYOiBPHKO++vcFzcLXcf6l8IMQmNSTt0v/F1IFBkuyuTJmr4l0fhr
87refBW8oKS0GKhM2Tc9ldyCD0ooAK6AMVcpQM5tuNKhZaje6wb3Hq4+RZvp
5Ekd3thm4Sk0GDWP/pQWpb2ZW1hhh3BGh+W5k4gCOgh2TTvF6uNHe3/sEbFj
b25M9Vtw0KTiTBnhAO3A0wXeWIM68y/wQcYIgQu0mht5oOSIFX8D8Jt4DhYj
UnOGV3vyNYLct1vHIfkMF4XqWPHs9sQ/4EX1XQ8dhWTBeERPwaDmQBuAbpAQ
nMYGAZ9EM5wJSMJkSgc6swuOMafcXcWrooVcd7ckUjOi45W46277055Hvkvj
qfHUnPymQaM2kfQQLkidPXWP5YIaY8abqAoD3Ww9dEpeqYLVaEM0T/cfYOv4
AmdGoSVurzQ5ICPjSh26jATAtclJrp8G+6a5lqiRuqC9a1v/AgqyRsHqqbUQ
29MnleF9TO/gzzeG7/rgS82LzJrFclUgrqIfm2WBKg/3sAH1frK3HPrf6v9A
sAW1uDBpfBjHHzCEW7+Yzi/JbsL4MWHsq7nKGBK8pVGQ/ZwIrRL2/AT2XLgt
cqY0IxwQrJLMvr7BkAwO61gxIdeHtjL0UqYx6BB5kydzhu3exF3YaWUug7/J
t9w6x1g1055XAFp3SOM+BXaAExeogHE5rioe9qVldZZhGotADB/jpcBBpFYP
HW06dBYXzeDIs4g8wD6RJZfzza8OHGaVIz6UHVKC/WOcMp5sI2fGyRnLYm2J
lnUK7GHxPzcWsnAjGkyio/r+Y9VgagqvVwMQznZEpkQCg6JTFSgBwtTJ+Kv5
5P+fkQl0TMWw39WQJz8xGO0l+3y2nJRMdCuVARG1/ssr4YVcrDRc7+NWfcU5
qiR7oLgrcDrx1LwG2iGJAYaoiu0Vw1PHx1VdHOJ+wWwPmVSMJ+O2xFVsceMO
CBuW9mf0R1nLsd2hXEn10YLuE402YHuA+GNDfl56P/Vi3vmbPZNxp4575bQn
zg8+8iftC6UZIVgqnmUEUIoXq1RaflVuZvni0zqh2tXvTYFdVbYYy7VdhPLo
+RulpWZiNCwn/Gs5ifpzVNaHGkyOV4AXiQ8vFz7ioQVO2w3+H1/TiNDw43OO
pi58TvH/3/W8GWW/XdQeMps7B5TrNI2GGlcQqH5NrJ4IN9pOPJRdOCyUeIAB
Nx6aItpalMCnVq1gk2TbuVrFjkYsNhi01hwllrPRfbANrqABgF3MkNUQ5E+R
s0ywir9Nl2fceNYCNICrGEGqtXlek6hItN2P5jH2XPcHd3DdzQBB8l76uphr
YO4jVGVrPdnOMz3Xtxz+IYe+02wwNv1OS2YhSmOfzpuAUef+tuiowwm37RgX
xSpffpLlxm0AMsircas7CwW/mJzkTowi+7CrnuxKv6TKngvrYlbUjSsLI1iN
iaY47mYoAn+BkTYe+znsU5XQZDniLkUg6mdUEY4/9lHuEeR9k/mUr83hkAJS
U/H1FePmpc/GyCXBDvxil9YGYmB+ILO7k+KJkY3vMldX6UpzXn7Icle093DN
EIrjyGqUNuYyFDLlOjbnDPpZGJKjSD2MS/XWMPCh3nnDeoncsQPpYmrHN5gc
3DwcCMsx0qEj4VCTSOM58jPJjDutRuINY9IVwquMm28ZRkLw72l61sn6iU6B
wiIIvyJBAUJcvpqhzyrlIsXpGw77G0KWi1k6C21CEEk5WAlAs8lUE4EjE5vU
t8bnB/4PAX2W0Q/IXV44zgcXbeErIlfGZjA9TvZn3DMslcm/R/YRSRlbVTOb
HHSXLcB/XrD3yltS+2Fbdi2eFxzVxX3keo+SC7KJU0OxQJ1JVC2zGNxbiwie
OeNINn/52b1crLeL+OBdWT6QxjTrdebXc/aj1MBqqTs6B3m+2kcBR7H9fuqy
682vT0fuT7SHr6D7C+SWLBNmrqxbZkbK0YQ+y1XskLKDwZSMuk66CTkH721Z
BXMVw4zvjWYL1jw9PaNK654TtsD6qc+biRiKFKgliwB//k+P7v/Utd29/k2n
U559OZxAD15lUIYQ5Oo4xpAwNokW3MKY2swSD52M24PN4HgWc6TJKPbcmzrU
FmYDa/ip/hrOWwphUzXi6Pou1L3+g+0XvB2X7PMnbB0RhIjyNpjKTcoXiB3L
Ijq+g3vXKEgB1dvssXfbY+TTNWr1nkiYKQXDm1fgaWu5PvPO8njbJiQ3Py/k
7bd+7TDvrwJ3OObwa7KxpXG2b0W5f86NkW8Z/7TioYM5nM6q1IBQplFqwU+n
DLFNH845bhPEyCGFCSHP6VFYY6VAObqa5T/C1eqW5HPWck+J4e4Gn+6ikT8E
B4nfdfwwUkTsKEemrCT2pVniV7cxeDMD7oDOePLkOmPwF1dEKRgmcdX+sfxR
pjMaF+NfOQ2/dRRPXEk9rlSJc3Eh7tVeQjYUMACmb6A+ZKV+n3iYrYkvd7Hn
J+1n2AcxL5DfLn3wrdmCUgpqZMeew5U6VfxcWYeGyn2t6/OUdbAtQqR4pWdo
s11rag0RQfMNNzeXtDKbn06PSgSl9XzXx8ZCiFQ/RgnYW1mOP/zxCVgCTitp
VMlF8jAdIQtp19I81PY349UTLCUKipDSMP50KtqV+Zf5WLywkHBFQqnS8+RG
mqDMM8TJAuNf1ZygA8V16hMG6+HUlWh7x0UQ/hw+9581FZ1qDas6sE2LZt7G
v8OOjlMwPtYIHotKj90DRRKOPoC6vVV6ec858ZlH2hvgAyreg3Wien+k5AA4
jJGT8QQIagUsSibFmxfG9Zt0ZAl7Rt5kgoQ1fzf5K871ua3iktgsH2N4WbqK
sTVXxaKb5zovEm0138mqNIvfgDTke1RAyh8LIjC/uIzUZLNizf6XqHrlDla6
+vLNPaIo1jN4vFssCeF8TNIQ6R0kKMxa4RBvgmVhBJbuV62jtk0cte5mjy6M
nPuBY7q90KHrYnCasnJKYHOVpnC3hwWRq5VOBBEiO9ATcTnDrymXhqE8kNvw
IWMayC2meILgXSHO7RLY6Db+C3E26ALhUVz6w2bgGUMyIfWyXnkjz6nRfp5+
HnK9K0pWMx8f9OvJKc9j4kwh8eojNSTxBI1aJIjFaf2VG2oH9vwrhkqH2xIM
30x8txeLe/k71VEPifggK+6GUUs08vzNTtBGE5/BD9MsAGcfaGqVcE/8yYXX
It0CTM3oFR1z7Aja97QRy2M+J/e573B8lq+okOMgpW4m4u5fV3YHoLgGgfJM
hYM9ksb7zESM2ExrdgD6lRQ5OEJ/dqVv1fqa4fCkDfDZ6lkJlePfnjRkPmsx
G1wPOnYNAcNJmSNpe290a75wgXf68fdyw2H2TNy239cZsOQWuW7K7LxcuMhR
eAErtYtNe6n+cwsvxvdQZ3tGDIR0YDuZMy/q+j20ARfySNpyU7/CpG5xFAfN
ZB56VpnmrxB+BSmTXZSvAWXTZqBagPBIbf3jLu9NFXexKxPrA0TXCD/Ut8B6
31tni69noGBMQoEw3AgbpfqNy6zeXTFnATA2G8NWnHQVGLq/MXx+4tPghp1x
jBHAtUMro5Xsapratc/PF8hsi7xrpNlrq20Wj3edlPwADN7dBUSNvhaf8oAi
hsptfW8q1nSVicBWbCpNWTUDu8cjpqwLXfwLQzB100Ai05iuamTEsUBoU4JT
VhRN30xsDpD8txqhScruGtem+PGmA7eGjUya2qDokAbr7FEXq59LFlXKaUZ/
u3Yo0brt3SYMufkHSeTFtX9tfm2cwOq1nRaPRTpcaC+rmbxpC75xtQodECDJ
zU21kWDZNP5JfqLnc3+jA9rxeNvrnaQPbOaX0e4p4CyUdOaJC6+RJDw1WmI+
Wb+vuqNOh3hL66oPTKH1Aa2q9LH4X4xXFFsgXpj8Eza8Q5GnUxxd9HuXtisw
u20DKvxu+3XrZRc2P6UoCI5Ww+aeqY4PjWAZOQvT9lv9e7hWLzBzM5gQufbv
dEkxx/OphmBmdWm5e8SA8AFFQdDV8lKoh6uBpp7lhQIH+gPNBnYtuZdzsEju
x/aA6l9eQ2mOQL/PR7kUIAxC7AjPdJAVMAZCrZmAxij6GXlRZSy+gQ/+dowu
TvtOb8OIJckizvOm843ZaO3CgaSDnpfKHuzpKP6TwhMYBS12tjcsowk1bUiM
vASk6ngYbsEBd1PD/6DQXbaziFo089TzVGVj+0crNphJXUZ+J6NGNC00dNDq
CtPO0vZgVM8EpSsQUB4vLOloaY5zK3IA/K+N/4bGcACzyn1sKC1DNHw7+jDh
ty8UoGWIbUo+Lr7H3E4Qj2TAdjklQNyl51Z4K4Vifb2Y2j+KEzwUuOtpar0Y
Aad0/BcPUSwKW6tiol1eri16FMhvqOm08BzkTTJwMSxFlAmmu0A1NlytInQC
rbCmF4NIAHyCgV49CHPtItt+FP5fG6T5/KNYIIBeDQ+6YS7vSBgHM+N6YGZv
Kk/tlB/YeLuWSllDCg4s2PKaDn5LpHl1iCp5kpKYHRYwSAgSlrbujBxhXmbW
VkAvXBEnoy59EWygZ88PN/EZpwGKJufZqUKbYz3I0WVMZrkbQd8QqBW9vEKo
DWlpWyOd4b4g3lBO3RnRTj3wP28MEaPFg1/fia7Vb+FNJM3DT53cJFw2+8If
w6zX4kqAp7IzDAw/U4jNLvtX4g1gHkFmZ2DVdxbHWQnSKkA3G1dpx4TC90+F
oVcLY2Ba0RXPAMUh57/AJersJ9YsQv4+hMZXhwl00Tj1hnmKp0y1ytHqKEzO
T2chf06RGmDBNlTYKlLM8xgaTQCHoy4m1Wgdze60gcyEJIYeB47TxFxf67XB
gAdIs2ElbBGqp52YO8/HqzMHf2wYNoyC8kl1lSRWGGZeifyQe3qry2/Xb+D5
h2zDudjKVJpNZw0Us7/9Z0iPf/kqoMuU+uuPGyc7C7e2AMv4MUWpa1H5XFBi
MrJmav3Q0pdfkHUQOmCz+R2CiyG5Z4/I/yFoLILaNXh0FY+OCJ9sczs4ab2S
CWPggQm3O8hoUSIrSCaDyKe8B5frn94ENrO8/jRQIGA+2p7EwiZGGdzOy2mS
gwMDHBFuh+n+nzJ9Lqsa4bgJvEYjj15cMVTAZKk0ibsiKXiwxtTpbocOl8w6
itg4Gi22WLoKz1iAMqQ8G2fmJkRq6bS11e6vW7dNo48Fbe4aQT3YxZSySj60
0kQfxeMyiwuI3HzDmENoFSJ+qF1m8h3WEVIVgwfeqRPbnEBl013pJp2CUpfd
LR6dcoJp1cBy6lD/Q0QwxDYu2kM7dvmEq44pBD8Obm4gGT/4D6XUUUXDL1Vr
95mTPLJhZA9m4xrvIAI1WSMF1STQ9t0ZKrErX8Y8t8iItqRobUHu7R1sNZnA
AzIcwYJ2XCWPaHaDrmWUTUS9whvXi+CNEn1qevMWL67FC+EP3CmVlvFy/udC
Cm4ZAVxehqcBl/fiNCxaYjJq68YdmQERuuqSnCmgmYnl+aZVNfOWTDPEeWOZ
PMGg9F8L5sXr6L4G4pB9zPMW18YoVHW6roR0YgJs+hi5ner5iqbAgvvnuFLT
6k409sHalGYTe6DEkCwEclRtzoTBqBioX+SmArwB+Puq9DbbgJ3neHZrqUi7
QVxaS7Biw5Nd1EiTY1BdI5PnAx7dJO12sx4E5QHApYimUjt4l3cvK9YugWoa
0pbweaVDsuua0d/uv2HVUZs5zhYykAi7nHjND0sYwTeHmiVzYraAANfl1GvD
vRjxWISCB22Q7iJLjzKYw3iAO4+uUWygBVuuG+arGTqfITN9B27QqUSBK0/L
J34htLtKfxBMYhmG6fAX/oE/SUUU/M4ybW7lt/x2X6QpToMcsE6ogiXteL+H
zsxZBlYVR9HKedkz1/gQsOR6jYtJERaE8Y0AT6wTuqyC6DXhmi6XoByIuWpt
J7Y4KLTLLCNWTiGbVlIG4p+rZ9hsZN6Q2hiDxxWzOpSMHim7/xexE8MVbfcJ
ZU8scdL8LoYd9xPGCIwUwcdmJgDLbNxMr2q+JsQUX5BBBETFRpc71M9s6f4R
n3BWLyZrHR8wdhsJzDvmESzBZRh4KUpJ119OCZbyN8MP1H+eV93Vm0+ZGDhm
632UofOUX5mmKdWoaITMXCy43ZFm34PComWsB9nlQkmeUEmfRNZlJUHl1fYN
VxoJCV7r2hGW9d4pvjZBfdwwbwNUSbEpQBxbnK74WAI/W5wVUZc1bU8MJCtF
PQAwkTmrpSHNWowFrEG6NnNJPAZVUhohnK8dAv8qZldKEiAMTkvh2Zmydamc
UnFWBz3qO4moxfOVJrt0wYJbhAmZK8M4qhRs5RQysdMxbhNTbjkILAU+6NAP
ZpPOfOsg0n/XDLXGkS37I76F7c/YG/WMmw+gLK+NTlQl+HVO5Ps/BuDL2U5b
2vg2RDcVdyQ/zxdmDutlvSykfXu7R+iP+f6Cz9BWnlBMF1PSeZWICM2hdkf/
RW1zXMNVhqEgJIWZTc21/+aAdJ48LHuniSOELF4insbbm5hrH+uiJ7E3Z+zm
UdQAyUcazQPFyB9I33wbl4UJmWiWHhCDf6gQRuKRXfLWBbSztWofxA09wGpr
G2nYmjqG3Mf1vjNj1ieJaxugK4A19AUo75qkMty5WYDYwex2HJIYE+oN06t+
BIgv6oQx5qbE4lwIvIcszjKiLXu9vxUBod/HfxVt/J8kZi9S3JUWlsmgIYUd
4+P9QBH1WRVuYZb9l4YJOiZcV37bC7ntoRG4nzj458Ai/WYypbUb4OXXHJjl
xIqkOyEAWq/MudYY2Xq0TBoeraUAeKQ8lUrs1KJK+1i5VYkCv09L6kRKDRXz
ZT2Hugt73tDDzWZ00aDnpbdBzdjZX4tbIuDXw/XwDdHj603vWrpdTRkTO8HB
tUrGBXKsiDI7nCIJyJyMdDiCT7B2gDETOlhSWAaaHCRPFUbByvCGSRZRPrS7
wjNhOJ4ADWEehKbXJ794ViQg+Ii+K3aWPy36q2VEloSl498LIjTVD9M5qVIG
Lv2DsMXGsMQUVxtjanP8zUW5ezWmP3d8JcGT97Sh2U9zCBYrL2zAmfyliX9O
8rjI7r2mEQJM7FMA1xqSEfG5RDHxU2ieeheO4mxXTpdz9U2JD4MEf2G8eBXe
uFu2D9Ii2ooLddj7kUTFzzNZe1zyM3impjKJEAXCxphi0jbWVamiYLQC6j7s
HInv+0EQj6ts3yVl+N9SX8dvfjbnl3kCBJdoKp10nu79K5cqVXKSuivajMTA
8rrRc5jo/3IbkgwWFLF838X5efM3yiVRnmaF550YeFh7rM7QP7HSlEUyKHol
rLoyWRWXgEwev5ogcmDs8m7BU5OQmQwTgnhRhCgKcy9VyvcQ6HxIs+s8aycC
a7gPscpRytuRiYcqKbsWxjtwMleRYLwfXWBkEpyvG/ZzXRmg7zh3xZ8ZFygV
q3u/5H3qEinw53Vn4nhLFXeOHm+zv/62ZIkv/u44GNr4e58NrfQjGILpfgy/
PKrpWLhM/Ol4hUymrX6eRq4KHBeRnaAxmsQXtaTuvfXhCGEM91NxiBfC6y+c
V2Th+8GC/C6lM6sj71HxilZXPFo1nsojKGZjxDw7u17/2qAkjlsbPbpMO0jR
EtjkA+jU/N7J9IzcMBZsUU7tQYtWZYWoOBWORWC9rQBcil9YosyDqwWlp3iY
SaDiP047JaXZe4QrOp+8DRfCutyiVI+QgiqKVUJIE8AW7FijtLYSxXlB9nkY
ck9iALaj/nyObVIcI7Bdeb0hM0FMh7xG6KCUW7cO5rweWY59+0/mywFZxKj7
i0QfJxaTISvDrLId5nAzEev53pRlpqWQNvDlckotgS6v5hUxsf7EA0+6diWd
c9RVWPEsnZ9idMcR8cxwqabx5VbV2nDGCekFU+hMTg19iivQUzbnluLAPqoM
WbKHKD/7xp5iphIYgP7+j/JC9qErd4pziikA+8KXx7LVt2cKAb3KhIFBJxGs
jBZt0+lol/N5GnV8pRdoVtDTG5awTObmxtAfpoCvfRuBE7KlqxzadfM97wC4
SWNFss0rgXyiT37OkeuYhOrPHW7Bh8kqPoMctaOZEYFH84Op1LpUToBsh3OM
8a5FEmnw1sUOZ0C5qEzmIyHEO3CK1cFitU49aR4IJgWhTo+52zsLRicIz3Js
Z4KuwSzs8REASGJ1asPB8MjJnwRr2cLPo/KfwzKCj75iTs0Rrsayhnon8vWF
h3k4T1QjcXInX9YnoGMXeBoWSfBy74wNjscyda8FxmMdNZzWA+tYBVc5BEV5
h8hsbw7hpxksgC3qCf2jv7++TORkCga7+zhJhbw4S6FLR3093F+wct10hqP6
B2m8JfPCe7vNnEb+lG8JF46+TwCsVc+m3TJ7m4kfcUVSy7DcRT+ewlTeuLUw
CKeaSMkrrE1C7vj/l0dtVl0IbOi5Xyt4h1NkO2VqOhfPhTDjvAT0vm0NRbuA
K6CQ3r0bvrOIXiY3FdJP9hnFwiPbNcD2ziV18SufECdF/lODCn1nAm5tJi7L
Qx3Msmw213cADtzXmW8SxBTzZkJ4fsPGTIBa/ejUAhCP4cCj1Ad01xHebeNX
PT8uiOlbHLQ8YAfAOpEEq3mNZZkdY2isvQBLd2u0RwYUItTuPub7AikPylBl
UlHfnepBA60icXyoS0OS3Q4solWi+IbjMdHYYvKf1F8BcIFyAz/BGidAZWDP
+XiTUxHz2hKpclwiielXjnOJtACxNq2WYE1rN0yhtxTvFjBQ4tt1tZfGKE2h
squhwv0V9SuMmAt1VZNKIfPPgOM+RxOrMN3ji+fzNeRY0i0cHwptY65SpPnr
RW8611gX12V881uwV9ie4DNytQgyFg0k38iAztc9LY4jh1tZryoT4GW/itD0
a/pYfKaUwz80McjRuPfda09MJ1NDxEn2Nsggjyim0ZAnMlrM5Pi56WMls9pM
0l7b8ilasE5n6vg5zh5FxMLIhT6ccYwLeEq2w4R2bTJtGiZcjfSq+Hzq0zHt
Qsryw5Cuqtkz9fhJyoKzCDmcQ+28NcluiJQZD14zuyhxAoGq6L0ifCsyuUWA
AW9y3zYt48NxcI5KdjH9xkQ82F6ayTDbDvsVQ4apy3kEDGuML6+DQ4trapkg
O72W+tAfqOg4iEr6XZxrQl+MgAAJgvjqSpv0yf1I0s15GFRAEsdg0EgKuplh
FF6qfC0p0hKwxURaiuwuED5dNef1aM+cbFmljKuHqJN0bJRcT1BUyXLybJG7
7ZTw5ahqSSoMtMjyyYDti+Z6fmeAoZMhBw+7h2mSoLXlcjoW0jTEfqyQr0yc
IbqT3zlRCfKQW2ELe8ntSI+HThEmPernEK3t5WQYZTTRn0lDe9jYdl+mvMj6
9PIMQDYX2H89NlGXUarnukHUWVux1rq5zf+4jWScRvWdJbPKxugFmgO7Vyha
lW2om/qfEJJmdwC6nyNeDwgSdW4BAt1NklcdVJP0zaTURU0hk1y+lIGjoNcp
CYyPv1c28vhidtsMQ0I5oZkm82PIbdMHTRR08hiM16IWT9Z4y6ZgnBHRqxyV
e4q6b6+9wiKN9TqzRrQqbPSrn/gPl0RbtIQM3vUW8zOjoPuIKHyPAXoMbmhw
LsNMNFxXumWXs/scB4AzJpDzEsa2cwd0nU4YNErVtyjNSxVJ1sOM6axEpSPG
PnPTpZoJcDv6KRQEn5BHvCvEBF7IIAoQY6jRw/zotOpOKkz7VWePVZm2fAR/
52nI0FR9q8/+Odj+iuIndaAInYzBHPpa217DyDoSk/EZ/v67be5FkSWj2yci
t9A51zYvzboX5kxI6I3SgY2WcUrQkdSR7MijzQCr+vhk3Bo5sO55ji31kCb5
yhvX0X11xvwABbYNMboCs7+D9ytWdCPwY7/ZloRZQfV5VjQC8O/aHWLUSkSu
bw10htiZLCAATqv+EJCcKJFr1tqMTvRrXvFiqbdc4oOqeZ4nwP+3ZnR6tIZ/
HzQLT1SIs4Xt5W09s6Bfj3H4ejk0j39Y4RFKhDXIgMtkc2+frmABxVSyQDE8
2YuGOvLFOq0LsTrhIxOi6q2z8PLNgnzve4YddDHn08qyRejoqHchpmzKrxxz
nE6rDooKxRO/zM0n/rDJS63bcbpe34ZR3PtZi43X4RdWC3/z1GVMt8cxaQ/r
c07jckirLrkEg2+8PWFDPeautU6/rRcAyF4XqGBx+DoIf5em9QXZmKLTSOSs
AkR6hlAPeajiUbTQdPDg7h9dJjD+yRApMR2HQKwPsvTvE7jAIlamG3j4ohZa
jRv3IBnsV8cN7HejWd7PodjnXC9I9cVFBogahCiS55ArLcqtiJIHynjjv7lD
T9xbUobOEP/Fyzm8gY9CjIZi9X7VycjLO6P6MedJc4YJVmqOrfxn9PZh7ztk
kdLGBgBw+nEEA9wH4ldfUddG5vcLxaN0rytGbG4BvGmLUYn/dKD42iK5JLOQ
CjmoH40NXCgs6Osv4Qn02EJvIbV2hPXuFl1XgUBP241vIEdhmgejo4dEPBoN
X3QAR6t+NZySTpe+CZ/zQyeAs5jC6V4CLNWP4BLEJZoFs+y/Szd08vtg0fpT
lnR3/LuWx6pi26ge3CwOKjBFxBAaWORFsQOVAMH23mkIw1sdDtkJe3ZpiI5L
4l9IMBip2YOjeH8HkNxPr+8qptJgQUTe8HWcono+ji7ScczQSxplHlk9vCms
JXtOBSqfGh05LwiMmyhKKBgrw8ZiEhHNJFXmNbtHTvjc+HY9NhK0jV0eM4hx
8zli57FtwKTxvethN43/37KNumuitYPpzBfGghp/clZSlInKyjwlDxbiB26V
wP3zt5Qim06uOyBHP+b2EkfI6SD8nH0Khd+V4KOkea2qwW7aMr+hepQ48rTN
3mcENT4fCzJZmL68PPxHf6dBQbznGVXI3O0bEwokBkvmokhjIVo8aED4kuvw
/wWXaMIhqkwWOteKWkNdd0fvSiGlJrOzHRQQn/7VDz8cVMOUCXftaTTXFeyZ
CYjfs89HezDT6FTUUvwjNG5jXTsDs/JGHOJyWUEhC4NI28xxArTQ5OfoUolx
HapnBxmRVOUibSP7MCXKvhqtHQ2iU5QHj7YuUQfxmJA9aOS6NFHNs++lTya+
Cgx6YoXOFS7CPyYV0L9N60PUfA2SdwZ5NAT2lf8VKFUdIOad0PM9mSGTeJz3
cC/Wmx7RGlwMSWNlWWTCTBlmmopFDFV1WKhaOuntC90sck+je4z3jPXu5bK5
xU6L9/Ho8J87RqM/FIB0WE6HEY/9L5xywmNPKXTamPYCukoBPPqakSkAZK7m
DgNI2K0fb33rlv5zkNC56XZS0YJk3aw63t+5aCyeTKJI1wIZz1IobaVaEvHM
LxsjDaMmCdnNuAZs+x8yotpdXV4sEGlfdnLVTr4wgnnbqEmQdLBSUlsoBI4u
h2+yHYxyDM/C6ZDUjBPuddWIQsosaxEBtOPPL01i/j16yl6BZ3Yu86J2OrWS
nXK48gopydM4XgDj/GmtZ4ekFL4Hso86PIDCdbr7o/3FgwuPRXDBNi38oWuW
1G3XquugGh0fBSbbmtNnJlGrGwlxx2zzWXvZI22yhL4NSkvFFPbOpqp1DgAv
bU+VsWkXv0RKP6E5zdtviDSwh9sz4tiTx6IAxiJ7Cnaq6WrUVNlDgaiCazwc
Tzdm5idzFxJPbT+2VrtFvyOgzrX3ZD6JUA3K05H2Gg9oTTBHFzDwe2SIowo/
fWmJX8dh8nfMm9EF2XCTfJbdGy2y7FpxI0C0A1qwyHnCb5H8BCIpZnKecbLj
Pe3ba7eTQAaNqip+E85+nr+RfrSVoRA2Bft64jh1L66edAQH8tayxKcqADUq
k8ZK9abU26DLrMmY0C5zDSjYpIR+pmwY26lHrMuQyo/y0FqmNqasgNIkCbzo
ZnMhet7n9VwalvUmUU4MLnedvefgWPzsHC33n//fMZent0UjGOFbnlGyuIBC
treIJLaIm0/LE4w84rTGWQvcLfkSPNPfhJW2qb1YvuHdirlQlN0l/uKaTG9l
Tolf5uOUV1oqwYNkNXrI0KMQ2Z4MZjNrTFQmHiaMAD+8Ow8kCrPu20VToSoC
Hvot9RFN4czasCcSB/yAbtTkU7NuPOZh4qQ3Cak40wuWmzj/B0LhtBlFrDUR
fMRY7gl3wU8d8svqxi3wPKqncDVfeRmcdi2NVLxHjybfsQcPMqt8ayHlj8Gd
0mjxJSVftrMuC2H2oeSG+KH2jddoJBHISEpFl/ZAv0FgMkYTaDMhWo1Rs8lp
piVDsFszGgSlO93ZHEGDfGbIddlP7+aUGUFSIN7N+pbnHK1zhajZxkNst4Ij
h1T+1u7XVzkAejE/JgcQPqLy+MVwooPJqef9oFtFCNQIWQ25vIDKofBz+vZL
1eTjkx5ebqqZIM2xqoifim7QYXxBtWkY2VKnslCU6Jp44qfmsfJdiAgCqi80
JiyEhsbGeC4u2l/IwynLPTi+xoaqLV0RFTzcVIJ01BXt6XvU4ZZY0dqSFGkt
Zwu3jnQPorx7FpFlnfvT6PVFgaJEm5RPw7gbD22dmD1Eb9bN7+/aAA0qtVL/
wVA/T7nOwD13rtwJFC/myDcIEGUuaksfj/uGpyFuDkVWxV4dF+m/OcqNU96E
tllBH9LQorIQu75BsmgeBVcHT/EZEby/LIcDM/UwS0Fz9SZWStL5QJfcyGUL
2BfUEHaeW7icq9zQjO6oKA/4iktH3HVr8kBcC+H2Tvb/Ejqi6ZFfA4GThRf9
xN8vdKWDc/yruHhMN+vlSQh5ViEMSBOYAk0FRff6wsC+6zH6iaoGh9EBO5Py
k4DVtQpc7iKY0HCUqxWDYFtRkA4XOx7lH6msqoQz2K/Z5xlMLjGQ/bwTnBWR
I8eJ0Q8qPntmhVFbkcz7gMf+t8FHgmh/xCOuBNlZ3l1HucGEO+l3km1LGotl
DYh1KOw906eB78V+01aoyGewIjpyFOsFu2XvhQJi1j9vXK7gYj9ogsn3WADq
LaYeNtu2untJKtQXszSorL9fA/u61MCq94mjsBT/o9lN+5qQZuyB/hWlwm2V
mylLYY0xxtqmhpqBzK1qW7ijuSbCkuj9vfcMbOy/NcN6biwCgr0/WoB9V2id
PB99jWem28mhB9EG+a1NxwMZGA2/dOPBVOAmRWu6qeBYNOcs0+CRb5Ev92E4
YwgK4bV7e7e3gcm754HgAd17tswB8W6fA7Srhs8J03kWGZtVSBqYwh4mmTfK
rwa15yjC1ou/Eie/SgIVbv6/6PbXu9Vdf13sOIGAVZuK5C0IMDL9cArKChfR
y53akF32y5HoEWKAWR3ArHKvEARNiaP0KNX5xb8C2hpDzp7roh6XKMB7RPMP
zjMz6wVO1LUfnK02q9712LMiB0tDc3jzfhCLYV2SoNjtrXIdEx2zecx9N4zY
Rpr937j4wdaIdjL8d47QxXTmOlotB+iJ2yaiH083BTEHAxcl34/mdvPXXk/4
xdFcN2v+IsFIuGJb0tig0HLgUxjHX7ptsj3FTGPPcDVBKJP7vHxMLBtQCAFC
2eTKauTtCoVYGbDvNnWPdecFw0dHu9AV9ZeiCebYn3gJHc08Yvl0Gv9zmJvv
G2fj2AcKaLYRaISOE2Mn1ztO1KAqKEzsiqaIN6RlxW9MDiPv1fiyqJXSluQV
CjuN6zcYagHYxw8TPPymd6Y7EpvleTdSasA9H0c3m1hLgwMutwU26FBC037Q
mZpsbirMvtJJB3LfN0celHVTQy+IKKUwStKCZYkTdn3zyeQWj1s8Wv/1pT0m
cjNeQf+Yim37sXQrb3mZtaMgCrGMg87zaipzn10z8NxjXBymA/nTgbxr7cmF
8EN8t/d+DjoZ4RnqVomZD/qN6KQANTidsV9rcJ1393q/OWLMdbfXP0ZYIEzx
DcV9ICsCbOQquVXdXqrP4O8x5BFmXRl1UZuynlH+WDOHYzMIaTVaJoMQPxMF
IigQMK9JdWKqX1AqniWKQc73tm8aN1EmmVGtijjBATfBgCUWrLPBOU8nYePm
RD20qD3+bffp1C1aLmFh6LpfqsoUo6QKd6m9T9i3lHDJPm0c/7JhT5P065yZ
bBS8OslfhtM6H4mgDdGRBYy7vgKgpXZ36OuOKCsHLhXk04nT8zpz73F+j1Tj
qLaq5dAim6Q2LaDGkG97cLQO1gTn3+u8wZsXCbp60h/mpVyeV9YZdpr6tkfL
vVGfjDmsfGebjKkrWBd6jyOtQ7+h1bTaBLerZICmZycFBIN5TPMcpEf1D9dZ
NAscFne4jB0xXEmms3NW06vQfC6DbBp/y7J4E8dHfxcZSsrQjGbbm9f4HQyQ
k3R4udyFRdmi+wgyB7pHv0dqhtNpaoJ0jziTFG5YpNBQbkSV47RiPgKdF9cf
xdux4yfTYwi0LcOeRPrWM8M/eg6LkCh6sTAZGV8cPCcl+GjzzmA92JL9BN1C
XKVv8K1KvMzHF+a0qTU0DHeqUOlO/VY0LAP2hvtj+OxJ/2sBfiXuCnkqwa3f
L5vv0K7Tm1vqPpiUhDUthoyhCZH2RLuNGlov3MxdwQplvvbkbLFKbVzMR1sw
uGelcFHMwyjM/5aRd/CjhFWSo8YGpHPho4zjsx9uQie0YOH7BPRCj5avLtnP
DfEwiimSuC4uLCHe3EvvYMkT4csueEVEdkncDEUrizSSyj+Bmlj2hetjjsqm
ZffMDjoVR7Sj2qcAuk0sJC7dJ9+u+1pLwYjL87SGXJfJAWaRolTo5lzHoS/M
D/CO954i7ZISYU0/98WEyeuAS+p3eA+aY0CKlgmi7WeHdAKC31EJ9i/8CwTc
bw/asV3NAg6k4CKHyx3uRf6sDROfjT9+56LEJTABtIoHon37NlV26iAUnbir
Re8cB7FRzh8cwb6FzFf83u21pXfWMvGSOSEg5m2BY4O2CBNCiy03/s/RZMwO
EMOlvW2fZPOT3YaZhoSmbpzIer6p1eLJJB5HP7sAhXYcCNr+wWc7mJ1sqo7N
gzC7GaJ3o1eJu41YIUjdEwZELNhKidnvEd4Y++xkVj1BR1FsJ14iFCFnJsDJ
I1bbLszfnMOOYZNwctTRHBEHI61oOx60WymgARMh8OT8NY+gTJVz5pIe1Rh3
Tnp9KlHQQ7iZtEqnR/bQCxxiluIP8l1va6nW5vU8+0hNWflhTi6FOQZVORPl
Kz1sot9RY8kVcvmln6sl01fZSPtGG9NrLuE7HBzqCbtcBJ/lmyPzj6FzumF8
3OI4pEvNC727CnDMNLTqpvrHDBrcyUcu5QHGYvEyD01AUmvSs33E5hYj8vVv
jX5PhkOzY/GJ2DnipWoafPbh2fWFhQWXTuvTvlM36QJ2zvZrTqLBH3MTWkpQ
+xEuW01Hbdhz+gxjRCropM9BlVM0VbiV6EM3cff61jMIEC670LZD6T2x4Epn
qak0C+tU4A40k7S4KTjAPTEbe3/oU4/cQRYCMj1nyo320whQm/woilAIPgH0
cwGPmR+RL0jhiD9GXUNB4+6Gq39pzp95+AaLbgIgNj9lzRyZjvUGcIm3KaZL
eYNzj8DjKNlXrzYjokF510NJZI6Y8jY/BBDFGo8pr/kJ+hEauGnOk+FDSUhK
flKo+qYeeQ7Vr8EAjx1Y3bTg7hsMB6zyz/Ymt7/ijxw8a9ZK6Jkgsydjiwn4
HVGATPKoLN35GjziWjBGrbBQ0F0GXnvx8GjxUGebKcIeASb/ZkWa+Qc2yjoj
a5h4XqcZQ7IrpaJdaEcmLAQFOKuZ/gULU3vnkMrqVb/8t+wWd4qZh8Ya4GSa
zieUlRAlhkiLW96BBDrTYdHHCgdCiyTfPZu4iJ2gxavD6QOvtMyb+viprImj
NcSgvdx4SCCZes/XMIpe1fzHB5HuIut/Zz72k/rKgrLBXqMAe56OzE8uhXDs
Lp/bc7hNrtmu8b0VOd9WdMLwHuwIvy3caNikWnvnpzX5oBEvlS8XjsJ9mUxy
wFtDFSNxplAhsg0oBmwEo2MdJwJfsqvLmHqgjSJKPPAK/DArmKHnpgeTbf61
a2pkoJFEb8HWh5ZAi2N4yaW/FP+phic0AQTGVB+f/Q54JrSd9RUdlyup8J3k
VF98IJv3tEU6yO1i80YgYWdC3G0DcNaw19jkxbgVNVSDHm6G7vcpPAZ1c6cd
NWzvlYUJj8w/KusRLhRFQn6ODRUIjmQZ0HdSwyFs6GZe9wCpC8dEBpMLDsR2
pICM06RLAgFWRj0onZm4BJYFovt+1dNFbotVHLwXKfLiqDd/amAtP8LFTYl7
SHo49RMIyK9dDkO+l8iD/cZcQfTosTCuL9CTKxj5cZglwblwSD/Lu5HIvDtc
slKEL57bRXXTWTERQhc2Pi2BwgAF1+/8KSkAwEk9H9zhD49iDCE2Vzc1Yn7D
eIr1uMQ187LGujHnxYTJbjyWJGYsaSTSl/sUKDgZBynYcM8itAMhoDDIg97F
5eOjJdfQgAnz9QnCh9LWTcRb1YHc/PcRGzUQFuYMg+2y5Waa/ZfvMFcLMcs0
Ahbh4AeOH9btT0/2EIo6G65cv5T77x53uJaVCNxzStCUVRZb/D9tX2ux7Agw
+szpVO5lzclhGc48/reT0HjCboor/1euht+30kSQFPM+FmBcKb2yqwSkRNDz
GwBLdKLdjDJuqjBGVzv4KXpzKhSZwJaqIzpBlCqdBH/bcS49D3Im8r6eChwf
0JU+agaEyiBv+ZkQ+6gV6hTTXamzviZG00LwhNNiRG464hZhgqQ6ZKiR/yqM
IFNArbsHFd/wglhQsa/ehGlhFoJPBBwYszp/kQzAaNUeRjDW+Tm7h+oi+uVb
JGw9QRyKGmY22IEKvBVw1KFzHMgm1HXrfoUvPdGfWED7MX2J7HAbJHgZV2VJ
7Tu7gI3AaO6eR+hJWygHssyMTJSx+1ZAhZ3u6YLcHTLC+RJtfZjmrhS2oSfN
XzCt0BOlZMi+noAiMJIPxVSWVcJkqLM9MBe4kIl2Phb0oqAcGVVuRFIXpcFG
KP3QPG3H/vKF/JreaNQe6UTc/0guvkIb7s8uF9nQQ93b07ZQyjuYVPsfPxN3
nqe6wDlXYPg0FtR87klFInejn/cph3+o1AiZgPGoH2fKmRYL3Ri+jD0aaceD
bKaMJug1eOZwCOvyiUxKOuS5b5hSKvkzyd434fXnP9wzoNUt7yYogV0Ae0WA
ex8EG3AzwOU1ukLYlRSL4+HaSF0c3+tNfyoK34lRuJUd+CwivbClfPNHNpHe
QbY9O7NJJ23UbnXEole9yMTO1wGUSfTpcyN0fjntWg1kXtY+VZIe0HBqeYR3
shPyYo+iVn/GRhnT/mPNxAQpqD4mtGPjxmMUEKRTSZcwdOSsuUeg8anddvhk
joRZeZKmQq7rTOQwJkvuD3c+542aupFwWOM56DVMsR4unqWiPemuoqDa54vJ
WI5FYyxtuNye81YVvfCcJOeKBXGd/cEWD8SAONOURNIBhIu2i+jBQhvD1izr
Zu7PA187jtEUgd4uzwKZH3Zij0+6uUjTWYdN5x4RaByNsiBGJsXzj9CT3oFI
Tp+Wxb1Xl4IGRnNzo4rb82Hr3t4HC+BOSyll//36cmQun+9LkcSIUkGBLsMP
TwBKakbFGugHbSK/kPG2Di69zg/r7XM2SJXXmM+rHb0w0AxaPxpiYrgfQ184
fRgGs1ELDTjJn/lIlDpAevtjtLlg834KggTR/NWTHNdqvWgIk2+2cliGt5Xy
ldXlU0SwRq0kUMRl7KNZrb2St2KhTDlusTLNAxc2q24BS5TVlfUgkz3MCgVW
mAsVK1l54hUtWQCRfTwJTIS11LkP+LJ4fZ1nANePLSXSFf7T45yHw22J9a9U
0Uu5npOY6GByQFP0kxzFQ5+2gvNHutHX8LbUuRs4p6miWg2WqnlfvExXsDD8
L200de3h4RUP7PBF6IdK1CdIudhZAUcLcIfl8oH1RPNS3r8LOq5YVrC4VO4i
WoF1Q5NHNjcGmWiv0cfrHaRdQ4IlZfnXm4p1mpxecbAaS4fa9YXYPtCWR944
u3hnwTAj4zzUcYMzKg3T4Og2JMyIthUBTHFMsQG/w5EPgwMYfmi6sZhsXW3m
PBALdlceUBI5HM3/+y4ydldYmJ/FLmkh5ylE1jp1aPh/x4okwyJ6wtLLdeod
qipxJoOvFXcLTxoKSo4YUCbaWOXPXHk5FpX/N4ug35vWazm4bt4KpfiXsppX
fU/Rsyq2BZj4FSWDiF3iLhW+/iJK7dSFKIZ5uL5axyXJIb+Is7BO/dl8Y+el
vHhCqZQsZHWTdZH1xMDHfhL3iWNXvjVzDDyPqa9CvP2F2YR+zsGsvS79mwGD
CJ97bhXRs0Dp9m2oGKhjYVP22tMIIafjjnUeOv+4HL+03xHWGcAGqIZ8EiWB
bEnbMApbJUore/0XUmV49tXp3F+XPyMW4Tl8OaM8vg4QUt2AMn4WPQEVJ9Fm
YqlQRrv+GRpZFLjCJ2shONAfGuFHRp5K7n/sPASBvpKQJn3npAwixI8lWXZG
igTtGXyTy5TZAyqeX32jzszcM8j98aS9/2VC5T/AfuG4cLioWG4z54g9amz/
KBBAgpUlEbOHg0YcINi3vJcEB3TretHtKF0w+wNYByu4BaBmUdatLumPHEmI
u+XSHlTSKnybKpdfKeDgzFbmT+udHOys/K6zJSAmYCQae5oKJNv1NuCkgmjB
R4CGwSLgbQ22f5yZAG2PEeuUvxMFmKV+vzLNNaCl0+nPDpbpaZn+fIVIELAr
SnXQvMsTcs04bmDkFImkTVBELGtObH9CjLjUqutwDRfclBLnWa+Lg245Qucc
KrCktu4jXEjX9h38teFRmQ6+ixJPwZgkbxlgCpNehomR4PEoBHfxt4EBXGPS
aQSBLfrgwtMb+J7aCNZ5B+FIvJWS3yqtWXexx2H0mXOin4qYXxQbrqqtWLwV
3WCuZwS22VTRHmDgYQ4fu9fTljGLChvMf5YOF1p6/1pnYD9vSN9UbsY75yhc
8/Ht2O/koiURLeaAs8zWjT72eIRmnVJUj7smWia20mon5wJaDxeOZO3YBb+0
m2+urcdJ/t6AeEl2HqPB2lW9qxZBf6LyhfLPl+MeBc8l2exijooSuxmQeozb
y3fsAoAV97/FWpjWWkqE9TjN0T8WJRHU41ocWelKLG8asRNHBQ3KBwTyMrjZ
+EjFPuh825qRsCCQlFmix7oFdLf1cSYarf6wnakGSINkxIcXtaUO4nUpB+lN
WPxDW/f4uxrV6dhTZJyA4tPmtn0ViZ/8Yq1aeI77rppPXxRpv/NzhOBJrqSj
5HnU+Ocz00j2yrxl/gx8wAXPLns00zpba1aicoFZLTf8Efq37oCjIKXRfcF9
8dXz1HjAl5gzxGQtEndkIMZNgaE+ONvcROHcQY05gGsVM3B1P/8CCOrM2zHi
n4IlppSJH+nzHnPgaZlSVpNYvi5rtT93rvUEk4jWdBGeWR+1hYthWsqPmjsr
gC+0mYUQJRCcrn/r33TtiVDWbBRb38p4Dqv7oR8g2NxWTbdaohqY1TX+0y9H
BDPlGNGWt4eMFNjfOAGapAf4w+yyyb+G9DpFTHPhMeGtF60g5aPuX5WjEjdV
WJN7zLsalBKVdq8LT+LU2C5bORWucTuijUt9OWlCN2EBUVTeftdhD7DyUGCW
uBw8lOqP1bnOTF6QRV6YqSD2ff3ashKLKr7LWVeyTi0pN+zW0uTvAfaZ0q31
mCC4JzpcX977NU0S9JbqLTE98pOXEKdV6BOdYhBsN/WCCp+gbvC4xdtum8D7
V9VhemrIFrDxODURXCMKuuPeHSklUPQGldIVH4TLtrAyCsNV8d+suCoQ/6RJ
d7UqtBnkYew83A6svKwzST3PPMKLd78HSHSHownAqJPjDIkV5kKeeqdQ6DzA
lJ30clyo0hiwUJZGGqbI/MS/MSuh6p7x526fZqhwVJ46LgRzyjEQR3u6MHTX
4zl7YwQjQrQM6hvHXI2P7w/kmkOmkWdSDLp3NfhY9mF5crdnaEnPw1wPqzo5
xZioRCTtCxukDpQed/3E2D0/wW3D4vPC3piIBoCaqFoqusjytcJdsrw1zfN3
Je9dr3gN61+pOZETggfV6YHTT+5ym6PEgUN6T/vHmy0e+tG7yddX3wuHwSMd
Aey7k/cCERh3xFj1nBnZ+k8q0XQxiIEw7IUFb7xAaWSAO7Wbkvv1XxUnIYnO
ivQK2HCffZZ80B0DOd7pnP/G93SLJ7FV5ewdKUrUp1atKJgDR+FLAnXwVPrm
FvETLAnbdFAZ4f/qLgCjw8Y8Hu3WVNw4LN4k73zGkfODUioJOahyIVqG/rub
9bZFlzIstUXcvn2CiTD917CIcOFHis8ld7Ad7hVIpvmfNqXWK8UQRnMbvAzx
GTPcTpvrnuiu9891tdbyByO4HAPfCjKudpvG7J+yvo5luyif2gZ830y2rcwQ
yDbGFRYtYciWx/R/rguWVDeO+kEA110scIlq5eRKdZf5X5/WUFLirrSACDp2
SWmOCe/bEKoQhDPRGZC/2xB5D3CzmrvOAL0V8Ey+UMicx0kYnO72Dwu6e3Kt
L4tx3t/JK8ycGQ/CVzC2ozVwCh67DbwtwbXA951KuJhjjj8fn727jC7sdWab
flQFnYHawJnjlaV4STdcS0qotAaNbOUS6Nsep8zlTprCaakQA7BUxdRIg6Mb
azCM4/O7a7jiNQlXBycZiWLVBhjrojsq8NjyOBVLc6y1kmAfqNIbui2//4jl
r4UZwdf/1piqKBY56ciN62/IZHFzjC0aH4Mhw1CTV71hTKU3UnCRmVyx5kLg
oj8hJQ6X8CZ4zveHNY1PSrczYFH+V7I47+FfwFxwieTXQQBlYkpJw2qAlseM
pcWq6bmwupmCKWwjWPN5xiSLUhpn2u3/L2gcEL1pIXkwUMeuAXcUxJ4eqHco
0IFRgVudyaykQXA6802w+mG7R4Mqfm7AvfWfxJPNYNnYp7OB57fltiqX4d3h
nZE0A8nHhGe/1KCoIAowp6SEeBSSBjFauD8S5/2B8k6Dsk6HcVD9jYVQQOsP
1HYdtBuUq1xsO1ew9b9wdlcQCnHjQXEARU59EZ9tTXKmDgn+S2KM6NGjjcU/
MTm82+FT0IvXL9bxiM0y0rVLenDnt+DqJhU/pfhjmMQztPSsPZqey5Fkd6YI
8tNOD/6I5SBgqX2+2WoowwWw3GJ/nUhJT6vAkA5M3F7jvJmUJ/Rz4o30mFc0
AeosRXMwa/RyZ3nz6sOjwFSRbMzRZeM55CXZnAk5aTz8iCQwbOATbpFh8Mvh
vlFRmcE/cAAcTcuJ2hgJzVIVqys2QbxoTYBDT057C7VVj7QTbC30eZm/vSlx
CBBkSQbpuxUGS19l5rxRTZqFhugvEDlNpg7qRsQPI+wCn120NLxsOb64qfMQ
2EWeAxpkASB3lKhVew7B8uM3XSYh8/Hq6z4OdTNF1z//k3cgiF02YZ37e2ef
1yQZXy2RnqZ92rKYLECFKbE7cJGNlxmOh+lgE/dwyHSLRX933qQRdBRhXgSO
31GRbUYMufZu6iEZ/uK49xeCeBWew3sTKzMMqPWw/g1KexYGYvHVTFFvvRDQ
7M/q8hyGNMZdCPF4t25cWistHc3GZLQmYS1sOaM7yC9/FjlTu4EwmFor0jhk
eyWdAtPxK0RDcIsEJm7Mw1POe5nK4dr2KVaH8g0+q+kAnHKoEQAgYFhWuoqT
nQt2ou1pcOSrU5laYioJghxnBMXMiG31BhxkKPFqyc9jj0/Csp6tcjglmqgg
6NJUBYEy8Fxu1SqetCdSsbC6VABi9SZLYxFNCcBnrHSZBfmG3P3Da1St2+WD
G04IFZZEZ1ezcYkSIHUeJQUyohLtyB8pnljMtPUPMmrEBxHRoYBhcD1gZf4U
192OMrbqSCZRVlMuUG01JW0+zUB1a+Nh6JpfcCy1vve62q//XuiYmUjscCnD
42xfgP58EbwFQJlhraRMlew4oXhoE+Derrb/dw4rhEsb9yM2OvGkWp5GxbnA
w9YlQ8S1zsn6amwpArJMycza3Z5voQLSPkb09V8cSSRi02gk7oUHlZev9nlY
MtSuiJfV/hTNs+msAbTAUcVZzljpJUzYwo6AqEiNbhNjMUe9QUBkMVS39znp
2u4dUJh9ETskTMJOq2lOJdJNhloJhhpiQdpMpLDHdWdM4Tald3CeJgbv2hGw
tgX7xGgVkD8zTNdkzm9c92ngAE4Wrwkj+ZThgF3yoFgQvE35461+tUXDxhmc
mDm71pBBtGlIY0xwaZw86BNR31urRY7x7+GF+uWIDmDSIDZ5rCjr2oj5banO
fETmISjqaFAW7JgvJ8GsRQZJzliBnIUDDZkB9BymIB73iKbNc2F5FDdW9ABm
k3VhTjbJDx7bWZBtRXRBD0ibxwoErbnpKbVvAfDlM0mQtOYz6n+96bU0KnY0
aSz56Gx2FrQYNowCiXdiVi9rZtmMo+r6ASiA9L+E4nXbUgU5wIiJLdRtAcAc
XBZXHk/g3m/wUih3zFkmyvqRHmmPVnW4Au2zhBZ97kjqrl5oWaenNiDGd5Gg
7JPcc+cdZ2HCpZ+qopZaTTtZxnMmou1VD0NbDAVh9+dfyWDGgiCH7epR3E2q
Jd0384x1yKXloej11y/xYxcH3wlweAHs33A9pyh9Jwg+658SKo7bIw5s7lvE
b9kwUwB0z+Ozjmc+/mkkrRIvUUmX8553xqDEnmvufqUKB4fBFuYVAvraiIrX
v29cocis85BVmYOuR0A3cPtihaQj0mkyPGSsAH3pLHcfY4lT4tQENemxRZ7W
5NgzOAHoYFxzUw92ZJNTsIX/Yq5fUoQpYwm12PbYxDYZvFDNQE3J9zG/AY2x
cQfWvr2Y652kPtChD6oobW27NYREG3HtMyRLY9umRRUA3OhfJTuHBGAkuKKT
gdwyz07aix9JrtuMVlO95ZUkdhyq/3yalrMH41YYW3+OCFm3drxJHtT/iDxW
Ip7lBb0KJhX4CY1S0zN7ySwj0pWDWPwYHFC06LOr8GfR+R+u5kzM53SBaQb9
PloVHPqL+b5hvN/6yQVvZl9nLyCoZWWHVzApumCYYaDwlNsbkKNyOoHJ+gQ5
4BKsa5sXgOiRL0EEKsHt/NK/T3yr951hyNgDDUByo8tUj5eoS5tX3aKPWjc2
JscVRMhdyAwGPBcOvdsUXFbNTqbzu2+BUUB3QWpzrCvLUgNuGQnj3RWI7of+
sB7oCQbhj7kQ81DGq+b2FnL3+692WQfXo9CC0L4giHXlYyu6sVC+AvOVEPui
VD2fJuGU3f8FWZduUsOpnqKMZ9KT3ngTH/e5HWMLOkkEkjxsFGUkpOr0uYCy
MdzKCo+CftUL0SOl/S1FJI9pe517oIw8UswIOXmu6ul01/pyMcxjmzQWKVyr
ZnHPvT+0/o3QEpSRYH8QlEaUAov8+FQslu8nt/mUWhRDse3m82zSc67knopE
r6mZVLcpmARWy/+qNVweLjhGrQg5AQJY2jfljMJTCHvvt3/eXHdbZ/GZqmx6
F6PTUIJLnxsOBA0Nl9HcT4FvYr0k7J17AcR70XjLsvAlArc6g975538VZJaZ
QzmOBTWZ0a6KXIziB3wXZp08VBTRqCejVms6OXQGlCFF4q8hkTbd/kEe7ZRB
cjIAbu0JJVqnbpAb2VHg5PY2TMcnll/RfW2jKObABvHmiy7U3+VZCrz9qQ66
PHArpsBSyrwGHD9rsapz8Rkme6heRCjJt33IlF60HPB0vUw8hDCLA2xRrQWv
kiGK0d7mw6vfPOUI7eV+np+tOOuYGZ2RfskInPhv7MaT7C3zneDj91xifus/
e/xfb24pef9KfLDNmrquaursue4709ly8E6Y2oA7V0m5rmGDNCVYehVuoeQe
9LJoMbu/hU7Kjsh1lc1dJPCyrIwdho38R/9S6foPrEupWLmBqYFKOXy/RDd3
EOaiuvc61ae+BKEfuCmBtnWRd1ejtFLpQF4CT3llQqm9d4da3JyJbuyWVL0f
4WniPVObXefDIoEbbgjf8Ym838DbWxU1RG932LpuM9g8H4SAhqPtifsXJQ3N
3spxbdoFpspbq55OmNUBBr/Axmugka8GyxYYgAUrI8N2vTTMBf4zhMd/MDGa
NxGBAWVgSc8v9+YJCMz/cKKla2Cd0HoYHHq1RNz4dqEvr6UF4qIgX13gOU76
sv6fcVfDQ5B5rjkM7qkrkBNXBoKlShcIyMkOR7U7aLJGFfnPRHM2HkHtGp1y
QeWbNZnsenm68mYJlA1lSEaPwJf48KuwNucQBug3hZWdWhZSZPWi/VVDGHsB
ghDwR40ekbm1d++FPLT27T/qVRpVWNpExVcLTDxwWOCoz6ITdmx3cEAAdbiR
aTL+arWeiR9l/MYbWEjnBDSwAM2+NKQtIg4gar64WXp9Jz8bijPTc+zsuyts
AGPNodRkyDeLMGAbLmI0tQKdvHhG+FB8FLCJnceazAc19U7hbYmiXmWjen+v
ip9+hnIVNvGujrajzAiWfywOfg/1GBy0Q4MJ5jifQwSRfVCZgtAa2jty1RZH
zwAAkeNC9uPw9riNSIb5Pqhhp5JAldrPcyBhdOBxXq/vVNWWuEYgkC29kp1z
h+4r8X0as/ghol+XtATYSSzWMwdQoah59hjjfVPeW8TrIYGQAZ7gRzzyUhmd
AVEhINkpcjgkGnliYOqedSuPAsQYCrPHcNQUrhVdyOhF796fEo/3fCR4M9D7
9C+SPbdSHE3e/9D221EkYlobr/KBcr0fG8GRF8nZlJj329+5Qxf38rkHSwbm
DWTL24IRk8JMssak6YrGSZ6sfCevMe0MmhpRxnyuvARenrSKGrOBdu4KG9U0
3DeEVIlwrgrh3HDaKHlXyBsLhWD0k4t8VkXxGZWtRj494Zj7qZ3bVPyk/YKo
GCc2BWwpNVdcA9glo8a41OQnekIhBQK34FkUuIFY0ojX16+sRQiCIUNcqQqR
jrp5J6Ta/qVyMB3mXzb1q8266gVbEPhh+jhtvpIz8vBsw9EayYnkY0nVvzit
98XcSvmscpBloWcbrYQUCjK5OCzCFwlSYdG4ZDa4neqMGBxm+/emFSIe+JCy
Mg2ZVEXPXNIFUOjju2ZWELgqwEQlN8/35RNFpez1KmDFTybDgDIRM1HGJVEY
L84/24ghnxIFv0BC+TIGeuiQ6UYrlLoKCRqaLUtRHk452/KXw3MhvcO/Q9ty
/LLTE3JJJaSjRckvcfr4WMJiHgEw7kJB78q5rc0vpYT5wFdo+0VMZbki9YiL
IHl/EPAKFjFL99kvKD8BSFgr3lKzZn8ePx/NBzI1Hf0eZw4o+B/4HYv+Tlsr
Fn6oSF40VKhy3ku5e+GWUcUWYJvdNXOmV5DQ1cuUzwX2pkEfsYG2q7A/oQdj
cLr0YnxDYsQHkf6zi86LiFhs986PgY5/7mZ6yvPDet5dnCVFL0mRhEv1X5fy
mc/AmOvrebYCgmFtp6N1bKVNMlc/seyjPO/v1shE5b7NFV2cjR+Xryai1egg
Ih/znZVOqwBWG1sMMixyjq5lVxi+6OGI3Qlbca5gSItdyunkVs+ZcSw58MtB
ctVADMBlxBK2zP0gaxXxxE3B9fhLiKFjTD+uaUlmakcUQFnVrU+CNZfcxgYK
lbzmVb2Y0F8713eZpzNxSN8rc1fgA4nDwpLr71RySpMIGAZOvn4SFJwhul4r
iwjutSpMKUZhCpDkW6oDxJXhQCMTjcZF4nFkyMc+zdoZ2YNfRoMEh/bWq618
utLal+ASNF5mjZoZSpoQDyrHaj0vLI70lAw5k4/M/RStGEibxdcjLasxKuth
IQXb+DZMPKA/3ezH595vawd3fMv2iJwU/PVe5wFiYCtmbsJysr0/V4hCOM+f
zxLC6rCRzjpjtdP5zr+z9CGVzVwEzoVGBSO97ccV8AOBDw0TOejPIcr/yynj
jiehEfQDUSAhES0/r7QYS6qkF5P7n46RtQ6daytiHJk4Ibrv62ueRmFymr0V
84ZIgUAwOpG/eDrF3HyEpg8fz7MdXcozNqelks60irZsNYHprrUhVxmpdvKk
+AIcgoDw/cJJxw9yeQV638CqRNOj7jtDbpvusuBmGG3eeXAzuBGXKOw3oLcx
WLu6oXP1SiJzmkc10oZh5q92sqTMiGlMvVgw6dclAFLqeS+RHAvYdWdGiWYk
Idu2+GfKBM20lOY6x8TAXIPCNoaMRGsHGIt8WGqtYouaGUFgBIIc9gS4t2bU
3iaPJabMfUV83kSusejYN75zTNtzCTKMq07N3lJ1T/fICmMKxrCEOqy0al94
SFkbvFIhpvgIKEp/yhNTwgNoZJQ2/5PMIaKTa+PbPRXExO8HGf9EY0GASd/o
44cMqbFM5JTpIvfOF8vXv0aM0VoA/agaqIhwC12IANJq8M9jS8ctcd5SvhmP
6F8YaThMqbeLHsaXI2IXREiUkSYzgb3vWtxK2wA9HZFbC29zsw02Wogx+wlB
ZxIhNCQGaq/6N4dBvw1CUTxrXDUL9N1MCteW++fhftJwPlanRz8+UOFPVHgo
xgPT+J0MdZT16G5idBpNb83DQt0UARNt2JOaYkscMBwTSG9KkmrLK7nq4WXb
Ul8fVSipXopidD3adPHVqo4xSx50aBGmZEzXFYeLLwVNwKtcV5FEMU0B9NBl
IgW+30A5WFvgwyDCNC8OZ7UDzEwmE1ZwsDpv4LLnzgZQ+WGJIdztgRHoesan
UT0pMWUUHL4huOGRp/ihUnvAq2hNc6R/DnIA4jDZcjew3pXfPK+sC6upcXUz
GJXEN7vtzRpDXGeam6gdKUUPhwHkcgLA2ZBhf6TNiSTD8x/DtYyPbc7qDKlh
XQ/yYb5IJA8zT6wrJL+CxcAsexN7SfGPTiGM+EWLCqh9PCS7rOVG5Bt2IWf6
g7cxBYTdvuuV824QvwCq1oH4pydf1tsGIFes0eaWkWyvnlhKBZpiZv5TMtgX
jSNzCBa5AwqcVAr7S3LX+8eGe1bWe3O6hH4XXdvJSvy+aZ7lX//pXwNG2MS+
wcPVuqX1lzxS3AzHGKaBvHJa3bC2G1XZBQe3BPmOj4XbhLYoTg1gg7duXC3Y
ocuEpjpgCnYHRUxaD4ql9sfWiiKtbyoz+xZI7YgjnqxNemp/ICKA1+HQoyhg
twnEc38pSnhrinErmYhVMvGxmS/nIz+Z0NRHHlgjCy+v719Ln9zSBm/mhf9k
U2C+/JTDImwM1NNgpZSgIG6IJpiH4zv2yKpGAS6pL2SVTyw9Mc63H73mvaGu
jnqO4iGoM8XXgxqwcYD8bG2CSauFudbwR0a6yIXkfBLIvYzdJqm01DFZ3N2m
+R5hLk7xvcrukLsFt/bHPtROUg1eYLBHxwkmmTNXhXN60nOSzj0gHNTkcz7c
J0ZtEYDc7RnRidzFjZBd+902TIovHjRsfPLL8dTxgGarLSSmfcKGqO0mIVui
yXakMGK0XWjGmlxYMzXZHaNXioHRqQ8Z8odhi6xY41VO+aV7ib/PVIuRfsC7
Asbi3qpYkT3P2NarbF1g+fLL6zJBLZub2NtRurVZ3dksgM+WumzTXdOINZcn
KZBzFKZZa4LrX9ln7cFva9M/FOBFZSCKvs65u9NMbKV1NyRG7ciyRa3ddprM
KUpbyqOgkJyXJvauml4rD5Hcw94Ig20Yis6kWAOevO63cvTK3ZLXACl05xFD
sn8zonJor6M8bDoIQ7HhLu+Gi1zVVbc43SkYVguw3XVYNB+cQKH48oVe6SPt
36Y+degOyiefbBr69TzdKtuOaPLTPWdxcuRKLPnPYZV5VBkuRADsESvb4sYh
nYZMaBoT+u2JCf7+a1RCipb/shZDOP/XRRtt6fpm5NVocrUUQEOFfT1FkBgc
h/NH126UA7nokZYamuLQEGWr1XbZkdNa/BLwYZhlEo42Xn5G5nhHiH5pHPgR
g/Kl5iciZg74a7NU8M7MzfJ2Qg/rgN6z9BI1g9S8MUr3Q8ULtnFjFZGlSvkl
1CIrU6MT+QThRLmqj0pfJnxpOZTzmlqQYWi8A33RWWCVnXwtpjbAdUShCX6a
PgvjbMXE3jn4Hba2dIrSSUrs199ut/Kmu+X9dH1sTfKzFbwNZPuesoOWFig0
Sc++AhVWL8xoBzlorqx/K0nFRw7QO9MYkSeCdCMUsQLu8GjXxCH+pdcPuekn
YtyBZ0kt8gHMD98I2Zc23bQv9m6RK781D6y6Baht02v8KshzcYOxZNH2PBF+
bFxeY+C7OvevD8/pBqI5ct3c5gK+vHHz6O28Ssl0kHiusLDAmbTStpKiIjyC
OvX7Pm/2x4wJU6a5I9hiS7rM/N/fz7vVnotnKf8+6lqZqSMXZpDBQ/noTSHI
ar5h0bxA7SMm0OUMHVfujXKtg3lEimitAiZFk5evU1SE1hzgGYCgVEOHgsno
gmwM+vtXZF8dc1d2sLsCZ5gmblga/8HFgnMEyN8cZAV/Qv1cITz6jbi/muWM
iWqH7TpK6R2b+5iVCH2rRCk7/wLvjcgYVTnrHDsYM1E+gO6m2iAbF1RPSyaU
lpFPqaOWZWav8gT4uL7H1oVbJjUdCoOEB3S081SsXB4c8qTUbNMxNOTH4Dqm
mhHDrfPLEkiLz4tzwSJ5L9HRprCx46vvxyYWuQ/FA6JLIoXZu9x5j1MzKf9Q
DcQIxFTumr6AKwIOEcWJYAq9yd+Eo/GNPhMRIuAsdaQ9ejwCyWnP4YBBbzEy
NUIIL5dLRp1rNV0aEBENmUDWilQXdzJcQpomgjJjfkNDrkiB59C+A8M/enhy
QhpKm86/M+HWe660kn6oGbaHpMzviPYefUqVZFVXpVe1y7bULzhvk/u6a9U8
DNGklj+ya4lvm+d3p4k3m+Exn0eYtWkG+wVddGUTO1OSWKbp7bsbE2+DUeAn
TxRlNXofnJ+Zm8yIr9WxpZjs4Ljx2I/SDEaJPmzknjpIh7TPwItBkFmdf7W5
6wXK66WktTjYTiXwJqo38IoLQPtA+5ZxcWXfRA+eHLKS0XjKwmYpzvjpP98U
Ia+sZ9HbYqiFnuF55Cx51uWlN2JoUswaKLPAnG5nMMwpQ8qy1cc782wFcslh
nBGaTadJl+9RBCuihH/rjwpGKYIvgf3m3T4mtbkeWiC/nwRPj3BH049/XoqC
irJJH0H+JHxUJt6WMaMUZ/bRoI63pv8AwAdz5km2adzDZTVbC5PGSUQ95QHj
jvdMNhdGYBC/m2Qv/TPBQbz8ZbvHriw2lQ2sIhitGWL8ZstNq7wU4egKpjAP
0Lkc8qdosPWnbkb8Szq/5K+fMfCcDzlYS6g2L92cfQkIpzjE7jfBbpP6kov/
ShxtApiMk/Yth8mC1TIYBoiMjYuXA5BLKDFOZh2W5E1KLtRU4tSJsF/GkPNg
qTGLPtoe+6LGVrtagC28+265o87uF5ACOl6vf3J6jDicYe2XQwQ6HPSOcQow
DWJUs9HO7PrTeBkcy7MiDg1+bhiAew6sY819bNLxAXWMNu0r39/AznnRiz/J
ReW5o1X6r0u07r+hNU1gVR9OGPnEH5AIDoAH8xm0stMjlRAT1iMwewrcyWzH
BrpUkDdVr1fZVpIPN5LMDBUjCvfpyXlKJd56l5j8+tayBSkt0+SXskgqPlSL
fd7kNWrQ1ArGomwpyUmSZccusgtvetL21YIo53Pmw/EPmVpMIUSJDuIoDgbg
Qqsvbv8BQ0rcpZC0lFYmz2OaAcWNAdXrGe0zPSu7VGKJrp9ZQkYqS7R6+KOT
rkJUk4UwTVEaVnR+3GQ+LJfVvajs3aJtbgHxarwcoIIg2qcYxn3AAdN0NpKd
7Knl33v03Xpak8NA2YYPZTmlVu+RFd5e0IoLd8Xn65u9T8nxUH+C57u4zg85
HrP3uFUM/DZdbU0xfQ57T/emPbzJB+mmiowofRkITT/t2qNLCpv1HV78hUfG
swVWZ3s8qXpaqtpy+7QG4R7BmBg8BTQhUs3Hy8lgn7rB5WcwHJsWiSeMx2p/
N5FvJBjShmMfr/OEV0hWxbW+5zjRP66L8cdugzCDtGiFGzKJaTXhCI39Lbl6
07wpdVpiKKCVi8JwGt054CgiWo46Uo00QdCdmPeYdBDE9jUVuVx3qrnCSwVe
IIRKFJmT0v/C4dXwDLQng6a3nPgaucfU1H6L8rMNHiKqzwU0tAcLfxK81ARd
p86xQiVg8whIDStJAIjxqoGcUoD7UlrkAW+WwyCWyttdIHu+F/PMOX65mwaQ
Yc6xtg4EMlnvd2xSpsIbCm0+qS5pMk4Arv80sNJMnqzp7w9xohz8XnWSaj/4
OZZ+6hhDXx6AvncdAy8KPTeyTBpil0U4lnBHqjmmxFnEpPptYEGbYNQKETAV
S4scPyDbqi2yT4q/RtChFQ8DNgq+7QahoWEoj02gxo0XnRj2XtdJAx1CsbkF
hUZmO4pwyMo/nKETTUMI6PFZq+dyjDuNjbkaJvV83c9QxxZrYlXOUWScviIu
sBniSJwb5yelK9r6vpB91Gp7Whf7SmjDXuGr8UgmSrkPjp+j58NvVk8bebTe
QDGzeT8dLnuxuZrN7K/HxzT6uBqSRY0dhxAqbElzzcLQlKzPSqG2CMBsafJc
vpB/uep4ALCcHiq6gG6iew443bHEIuCEVhD+vLQBSTRSjzu7Ab9XcwUIdeH/
+3ny65b+3Pr+IqmBDpj5kFA5KghFstmUQJapu/DGpoz/TpgJ3VzYhBHNLfN/
sBwQuLwmm301URBawMveDGMvkFhOfBm/c5sIWDv0ExJ/QZc/R7syf+X1SBrM
KUyeTqd8pIFzVUj0EMW8pIHvBnWTS9TlZZVkzAl4G7POYLiF0yshx2PzPrfM
XyG9/sReteAIPYz+j9Hn0R0UKFkUdI6tzpbbk44H4Njq9wA4VmTs0tnqefU3
AQhzzK+LSdULN4f0En+2RfGhHISZrlF8bO11kZ4BbBUU/c9PgV1Q6y1Iqm+z
aZ092ShlrIWpUHdIsaYabJJHlsCG8Ix9s3JBsLKFcWUIaAzWtstFNtzre7PJ
s8UJtAutcCm358FLW11bwZGoDSLFD8SRiwtPFA1iuN3GWY6VDBUTYt3GvDeI
55/4nwSk1sRU1/5DtJlv/tyhq5t0L+ElG0RReTJ5G54/gnqKUCWw8+NRzO25
WimwjSypSP3+LHI5FmuC9OvCyFGkECw6KiO/G1ghRmbBWT2hwi/1MwNWwlDC
GtiuMyBmR12Rjeax/hvh/4eUvxqhb9uI7Bsv0+YKiKPAXIAYP45QBO7i5U8v
CjHcQRweqgRTCKnSduwcctoNcUpKhU4+vz2esCDlWM8s+Eyw+2GTiJaUi9fb
ANoEnYls/rojr6ggZ2eEncGdahkWaXrONQmn2S0XNwFrtZvyg0kxhmHNlKXO
sx1UVfa+UCHvviJqklejq7z2Azz0Qoye8pv17nkinq/PW0akArsKhrpJrTLP
s0cHkJ2rBnH8Z9+dXKiGwfdU867htm/jVgSWM8t6j1+rUYmSMbUP+JbRkUbh
qsPS3PZGksOsxmw0xHLm49CUv54oazFI1SM9yWhgTYPE7BIoSDAzUB+403hn
oc78GqpsuPOPYL/WWZrajROheOyYinZGi5ECbjCKfDRu5MmshuJifUtXhR/e
fiSHnQ7DnY+kCfnNWnCaV589e2is55FypD+hfB2wopj2jQBJiNRlcJzp7xgq
/uWKTTW3q/CBta81K1UmqLw9E1u9CqOl6PZ4dAfVejvnrca5ltOtrfu3KIlD
D6mPT8IoER/T0d0ayqcU1wjTbVWofvlONRm9BymF1UJh4RVYc3Tk3qmQxJFL
5w3DH9y58X8pjFwaEu//B8ptWKxjQ0uwT19kDIHwcggscEeFo6NutCRrB25J
rs0FmQpkkdPVyWeQ2NYbk1Tj2k3xmmaHtv/S1XhkPvaCZFmxlwy972xCrWz4
dWZLwp4RmFrwVURY9GNBM08cysxWdR43JBZCGqhTUEyrWzsWimRC/b9jtYPu
GWyXRrZDebI9u8g3vmiMsHBmYH5FqG/LItDoWENfSXEjK2+SSCXxNAI8mqg6
TEniSX1PsBQ3dE7cmTIB26X3HXXJoYn5bGdN6k/uW4JcSzRNW/Bt55kfO+6m
EnVcxguywfThTY7kqFEvlIZSIq90rhMp9bXA3QP3Ev9K+cd2TSSRjGwqI+7r
CsqvPdelkVuf8qlMvDLPfWxZFHFckm71q4XTChg8HGKbMgy/3f5OcpXyn0JU
W8m3eFyQYSOClXpaDE6K+t6ZXsr5lE+UeRY/NAeJNjidaRI/QlMOWXreJ4+k
qbrcSgK45kbpPZLbDPbgMJdkyHEPhCdt1wW2p8MEkV7I8NfjeyZsdrMO4lT5
NDXUIDY+kLMluEWVR067CpuWlldWR1kdnKR2emBwNke9np0TT9r10S/wmjAh
iSBhNMVXGAtAHBK04OaA9/ZkW7CVKlRF6Irhh5lNNy9bqvQXkzaeA8EtCp98
jc6/yO/cPalbKM8zqwRrlG+vvtE6dQgnZuaNOkKXKPYbSOFJq25AbrC7VLs8
w1Elvis+1YgkIOev5vSBAJP8vNH8JOPZHfdsfLOAPwgVy61VfwI07Pg27keR
aV/7KBtGxc8shjlIC9+QsYzijYiSIbkkSnS/r+YMfkeqBW6QYsNLCUu+s+Wk
GAGceLeZDyd9N+1GfhcfST411FzxUPnuLd6QV+HUwcjtUOHTBs+BoawRXhFh
7ANANgrdQqwzhbhEXUtfQc7d0r2ombHc3jGVwuwniSF1CUgcmN3H7IZtMWvS
k53cxre2SzTnb6Y8nqkb43EId/He9cgZudTJDr/Bpw7or2ETLTgwcurdznc7
R8xF5x6pRlwDXXcEMiZhJaqFQ3XS9B/emVKJGkLr15H+vvkuGlzSY4o/i2qf
HMLCx9VII+byqzY8oQhY0pB2yUBj/G7jdoL23gcmRGzJosjo66LBuBKzv0fw
oKXrbihoIdS8pJodiX3IYoxXPr1U5OSBHG2ZLxJX/H8rV816TKlwsE8kdh8Z
Fb2abL9BQ4pHqpCuON31b8D1t67mQl+cA8+YiY7jYKLQSFIBFO09PZGJL8x6
SQDwcra6zUMaAuAErnH1kzN59O695I4huSRFo3rDONDMwuuhIyZl9mH79pJ1
Z4LQzRyXTREq5qxUcIlIV2gAP3WYJXtdsXk4RPyck8oPqdvyaDUby1MLwHNa
PzMTckHC2EM/mmjMCi+jXgyltzWqZd55/GeOpwz6/hKn+WZsmQJ8CJHIh8WQ
XrAjUD9i7NWtj3VkaiyznOcn0+PEsq8+W5/bJv85PBK4HpjLbmGhva7aKrdX
8nuho2auDJ/M0Pie+q5yc+aFNgGJWJ/XgXbntudfITHxoJ8iYFld2YJ5FkxF
jaRroMhu8z08BZGpdeAK3IYCwEQdadFpLggqXWhLyVRXSRKrJTyJ3vOpwQ4H
/Fvk1jmWXRMYqL8aBGxdcCP4m6lSg1VM/GNCOiuCpGABGjgS1yBz7Dgw7Eul
trkI3mKpyyqFtS1H3sczimpq1S2LiOyX33IVfZ5kwfIDl5gi1sOc89JSkfoV
CTgz10JAEUTUoWAMvPcCAw1al9c6isUGlz8sQYpl+d7ieOg6BM/UWTVl9FQs
ZpqHi+bp5sdweQx37cCer4Ca+RWpi8OemacfploMahGh9u8fK5k8DSYylb//
lafhhhuTv0weEUhOqrN5jkjIBkdJyCVQZVPiUVphXhvVLNMm4PpfltyR1RQX
Wsl8lC/Et++isnRIEmlmVbrLiWUtJhxBy6jSdVvfK7WP8K5+HNuf1zh5EnBw
JnHzaMSgRteyYBEIg5uRa89ZW51Ae8tcXmVHvb73OS6fGKyCIrSMmCyJBpSv
4a8hwMELSA35whZdv+oP6aHTBGuxyE1BucREifPiAmL1TbNq7iSVeNH8A6VC
QgAqAI/hG470SwSap4kS9NkivHhYvMPHjcVsEsjlz5hFItCvynFbU3KCfdZ7
K8loEwz3IUi0WuHJVO3os1d8Yk136OFhhn7Td5EYytu4TU/thCBVT51rsb/4
aZqzcYwBcuoJhWiRWuyI4a88DT3OOUxBtMkjzpXZNq2WVQZbWkvr9t01QGsJ
awRm0smfVXn23ZdgLXhVZAu0A4vcC0Q8G8q7IV1MF+qHtwt442cmhqtRT2KG
P1uJL59V+8dMQCeD+7EIGZsMD2J+24yUfphwMvEUdD7xfcbinClsqKoPgS93
4thZNWbblU9+sNdA9afPa3+9hQWJ2eQfHWufdmvz0ckL78BKQYh1WFUg0riB
ir4+dwWBEvZ9ZxGhsXCcyS7QcNGUGzTGGKEGqHGWoxEytcVF+GsvM2i9bjUR
NEMY1xH2Zid1WAaD3mtkN66Sla+RNTcJYJGrm4PP5MzzxtE/9yOhZ3c1OeHb
s5Ax/ZTBQ9LVCLQH7rYwZgo3MNp5/iS18W8rcK21aoFc3dNHQWjYj5y4Rhn4
edsYaLf+B+M0O1FUmd/NXR0w5yNVr4LMmRUSoEg5liqHzfZue7/NzY6Ezv4S
3LHlWsU3qO66uP6evpsnwz48UfY+FHIv/yd9m2AyXqsXMFnVS4MXp40b4bSe
tWlavUs3APWU9T5xEdnKE1+J5DdpQiLyTK8IvjYmC1sPcy1fGPU9J0GI4eay
sIkL9FrYjXZAL68fdF30eiWtqgkCV9mfm29BuWbAXU6U7CZRhy2yi6v00wvi
yBUvTgkNwsEMIFFZ1c6T7+9fb+w8/ODSOHzlRtEVXIeiHyc8LFbVEEI7kQVN
VgpMwX4lBur2miy3fvm/I0BdDGTZAcJQuGRVvBzul5cD5BZyjtybbK/w5tgq
lkqyuRJjnhzaV4WAmcvEs8zjqqlVFXFgpMDospm+x1HL53YCummQlScfE0Vl
yHFeclxJukHmyD1IEcLdJPBMWv6X4IVqLbPbMCZxTMZr6Z/b4UWKIDrn7bUa
k0f9M+MfRkmki6APheNsroGAp7W4IllInQfSkdVPVFFeqDdKbeWz4tAyfYHa
HFx70OOv5aK9T/JF3tvV436C6d6gDAQnhrBttSzeG0u7Ly8ti8KEIzkuyI4L
74geT5VMmYal6rJ919829zKLFmTnfUTAiLpcKfOCMOsqGSZmSezGXTFFwW1s
+sASs+qBibo0Q/JLNaM60nlcA0XREqAm0uJcX69gTS0wuRWVOj+iziQyEST4
XJctB0lUBkEW6mzeeXXUPCkZ0v0jcvEozWE59JFxoz4/+Kktz+FVfY61OTI4
EQ0f2g/LBFrwzKk5a+/pN9VP80DiO/26qH4XWcCASE4CqCoDgCuWNp/Iod5Q
qmKndvvYHoy//V8gQzOmWmAvYBY3//U4TXFODPypAUQcHjBb39hwjto0BGWf
/D7CGyMHmzq+t4eZDjRda7Z4FKD5Zu4YSKNWjmCTcSnItInp9H+CG8BccSQc
fy8weBF2dGUGnm2qMTMjmu52yxsh6XrZHOQeg8jYwgEMkK6/4yCQ/FSt9XQW
GjRUc+IMEfVy2wh3YP1E9rfFKiQUS9M0YTsszGFuGSCj78QBCVC0Nf8nfJc5
OoQ+ni5MCET6BiPuGAuQ3IWy5m9PFixRkz1uPzpmAj5lC3yyczEoawtJjJNj
GNP+nwq+sTlEkz1W+Q2q0WpGQROcFFWFAv9biU+ZLL3pSpA4sYBl1Nu76oPH
af9aJOVRz6yeDJwrCMqpczQ/WwMOWEmVhrKH2DvaTQki9tA+w+Gl0Qpwf2i2
MkhdkUjUC5mx0V6/knLb3fNiLcuvABA4+rmoPYbXT2fN9KrlMaK7NJsXh6Cu
tF8D0ULryvqZYV3z4OoPFBs+QVBz34XQu3zsjVudtrB5UDNQgQi2amr+5qNm
brx23ZDykE5E4/1w4j+HcdVh3B/9pau9SnVAnWZsuqljv2/jb+LCG3PkSiNH
EIDaCyE94s1g4S4mLPkdoU7jRwrLz9Bsa9lGAj1M4X+U3odZgUeqIWMXfGr+
8UzKVI6YCfgWWV6q6kFZiRykObiHcAl0FwTbTSPLv4gKJWowx0/uwWMsfjcI
5Exr809BHHJUMiLIKLsSBq7Rbym8E797BhHuQRK+OOFKqMla7pKk35B+CuHF
SmCyrhpPPvuidDJ23/YqfoWb9KuCmbXXUJiXRxM76P79cf83DRc4IWGxCkwh
6GSRye7a8/1fPQe+OxysjbRqlWUe5bbMMPUfW0sOApkRsUG3HIf4Fs2EI08Z
eZHMiKfEWvDqJRIec284xVjHspY8kw+5n8j2sHF01Irz9OfdTLLfNd88sCU9
oxqoRMqF5kYNvDPctZi7NFYolGGbZe3bMuMEKYsvcDpZcBL0iuwxJjRjIsKF
zV3jTPYFghjSxmjxcnvVHZaFBRsesHZqvXYneLVSSkUPko8ljz3qHDTwF4tC
jHwUKQ92aLInVjjkCvJBK9jNWBDjy52jt7r4PvhnqXMRu/zEJI/5xAUM6MVM
VHnCe6ZhDRYngM7HiROWTq3Hd8psvTyQpP2serozsAnkKX8/bFqyk4k4wDQC
9+bIp+UIN5mZTUVBPeQQCuw9+xLVTnpXahorfk4oUl6rPELqMe2KS3cjiDc7
Ut2B5qtQj359gINnxfBQeipX43/VUJzj5crCmrJGwwAnGIeZm6K32PHM5hbH
66tWivZ6wu/02EjFI8ANYjZ9TgLvVFy0hyKFVrE5d3LBGc/pblpahNUuogtQ
XloH8b/trGx+mJo9d0DoYtrgvFC/EFR8/ljWl2tKJXJEaSGpHqhKO7nhbCle
VIMp6r9HTlhiuNFZi9ct5BzQBHR+ijfNwgsT7h66ckQIw0TGahMXcnjupGvs
AUkpMIDR9JJv1oLPTOvvlZK4dQZpfELeUGSMDkEp34y7XgtBlCyZhawkq9eg
fE0nhHlYE3FBevowRhDuDSc4z2rb8ZesU3SFiwVN/48K7FvPtrEjpom3SQRe
qjfi5wBNBQ8axDFJbQEvzT0y7Pg01TUzLGobWWWFa+leGZErzrHMz7Z7vrHS
k72QKqsjos5HwHWhQ+6TG+o2niiQVDCCxpcDBuRgbicnUwdcpDmumL0YR9zs
YwsPHlytd8bTqtmIsJmSIYSxd9t4nFD3bhL4ly4kPt9khn/xB3klqAMGkX9w
b2UCQdmc+CCPMF+XGW2iF7cwUW9WfpwnyZQqD1ucu5sDM9EKRFQdYfHIwVda
4la50MURQCwJd/AsclIkJlpBPnFhyurIt1geex7Ty6FazPgMVmz2Y0jqxFjg
k6XXB2G2WFwBIpEOkOOceiGZ8PYuai59G/KKANm+rUX0EC9g3ZYowPlkgnVj
N7mfv948KcOaAyNJM1hTU5aIqok7WDp2SG3jEs1+SIkEmCRflshfG+R1+JAF
0KMBfbdt3nBblbAgMYHgpWwMUuQm0g3090PZM6QQnYMteF1fv+j8DUfLi/68
RGrVJrHMBFQY9Lkfl5eZFpVZSLPwJ7A+/L3Ogd5Rg1CwrFe09CYAqNOmu4fi
lIiv9DzyyMLrCvhc653YrrfGRhr9X2DvjWzdshVssMNCSUnqqUFEsa+ezMXX
Qwab9MKGs9WdyWn7TVkhk3znOECkLwEJ8zyX2UXG9UtpUcsD7h97gGnNKT+g
yKPRSOuNR+7Wjn2T7Dsh89P9KntJEc3gA0Zav8q2iO0RAKac2H3KqacAZIFV
lmRjp4Fx+N03CbYT0aRBSBM1+Hf3gAQPP9A4O6ptz7cMLp+aZ68MJL04bjmu
7VK2TCVoBc7oTWNLiIsEBl3d+XxLWzjkZFdhMH2YCbkeLOnT2KDi+CzvS1BX
p9GRZLe/Nw93LCsbJT9OKSgdveSCuSV73FX+pT6s5AqfnalRhIm+quNUPDaK
d7P3jYVR+l5IO59yMXmnAlWZ5qDpbX5/vvrPzHdavSenwEgaLFumuRAAgGEV
baKvCeWOCgKbgNyB6rWnmFxzM7Dj0bD5XWqKq92aoFAPMkJH2FsSgy6EvNxR
lateaP+n7ZhDKlKWBW8DbdrSjHujk8ZO7fwCUakPWN7+ecz+MpA9vy2zkESy
o67LrnpH5YzbelTBgZ6zHtV1pi+B7iJ7bu8KCAkL8exSqO3jcdPnZR9gH1+t
+F/t+dF8pFlf9HDv5SRhnbphGwpZ27StVfiFjXtzsgE/KkzFL3/OjgxRpVWV
DcCo8lmX/+E0Ea+zhwrKNpXVvga0IsVCpf9yXq3lLGTBVNcSHKZ26usUU4uY
vdvkxZC6B7BPm/nr6rO4GcOzZ/oTexGVLvt2WdtKKx6mvQH2rbk1uNY6tPwU
sWj4amuS5czGeeFrS8cUephlRO9ATrssxKV4my6oUsLpWdgk+Dp2owC6l3qN
onBPJ+qpT6JydPVsOVyMtGtwGe0dWYotMtlDlAzIUQbhOODZYQUQocYGVzDM
LXA9mRy1b1pMx4VK7g4NjwkIeKbquMbKYIklLcTPKmhRTSyYUe2KNgtl//O6
/+AH2NVno18CDPbDTa5hQxi9gkBgObyEXokVrALkaGHY8ml+VwFPnIqnUFdR
NkQQJn/GcRgHuPY65RB3zNHK2LSXMDfLjP9Zz1rDOiu6W0hF77GBxLBXtFb6
8PvG3r5de/V0nIry2DYmp97DmRPH7hcnK8WJgAKi9kU9MHPyplqIPVmt/9n0
cHO4/lrZ7WAAWhKS86rtQnDDNo7JorGrRYHn2DP0Q6A1jH3il1K+94+YClVR
uofZDglMCJyi9sWFIIoueoyaquCJrCaWpQhJcCCIiIR0unbLMhBLey63omYr
HdBwMm2+noJqcGAbqojoFyoMxiYktVI3XcQSEysDC8JYWfLc2Pt2aFkiEG3W
yP3koJRabRFXPFMzvjUfT4feq/2ZmJJLXsJ+T0PRNZVR7kT6hk6kpEBp2GqC
8eRjVtAYCW8beRXgudiOe83Rf3lj/CeM3ihC17klfXDo5GURLolhSQIbGb7A
63nJBmY1xPnBoCub69PFJNjMrVhehIk9eesorjgkIB+IWoltaZ0nO+RqrcIh
kcYpd7gqXpNr+VgiyVuhBWwyXzvnoO/xZgj4RF0qLJQRUvaqXLTSyU8NNn+h
QMJVnCqnN72BPSO7i6lwLlwriey2mjESKXM97tMcVLDiYDD6iDsq6PntDh2/
SpDZpl0rH69cYdeTyzO78TCeQBj2gdEJN5ojnC9i0Nd9napQ3GHQD0klYa3W
SeDWQsXXWxSKhyppMtzwSsRcMUWsB1+yHJGyD8pl5JNFFLi3Sqg312EaRX+L
E8nSAu00VZZl+qhpANwPK7V5bI7ZqgTjlzX7MstOkjFOjHomeLRCh/+M4llo
OmEthFmzC3F1dAK+7aovhA+YrN5KOGiIuuhIaA80Zg3QuAzzbzsjiPQoFdDn
xQ0IFOkfhrZD1lXqNn029IkUmPCFwhZRsNZ8F4xoaD/sw1b/S2tUafWixhZF
wwiYwg2fpGwJjGyDGZEWgFQGhF2Rl7y3Shr7zvT7ANCWJ8ikSr8xl4vzJSUf
3mF3K+lOH3p7iB0KmSI97jWvmO1RIlY9D8YKnpCmdAD6+LQReNUs4ZQ6w26m
4DCuYdUx6Cs57/k/dkIdEDXVJP5LANRHI3qVw8QUeL1EOIqC+MscObMTkH/S
bfrMPIY9olBCtiaGt3u2wIR093Grd41gSxoP9dpDn55pYpGtHfeeaqgeMhnM
d3GDjqqBOpFHtzFoj5/7hvGlHrS45AkGh67gjL9nT7POIKP17+ySgY08AkuW
SlRBzGszwY0b7Up7IDxVi3NxaWDUSiO2iYrGZTonYiZk4Y+RuqDAFbM01i1N
pfKMeHieeHfMJNRiIORN7jl1nsiSUer5NJc4kRrQcHl28mugbO0ULoXK4rb9
fr+/bqosVQUA1XKr1IEwibSzQCXW8hei7R3jN9JJuK67KuOpo1fUglDVl8u6
Arb136E1PuR7lDbLNlBjUaWbz82UL4m3HbMtATdEHDvckwSFeRKFtKTMvlpX
yYY1fosSDJkMAu4HtWyL6vbHsL1BdAzbuMDu31DBN8hn015G8ZGes9QBWAOH
VGm30BiBsdOFLiXhYko+ZOAhlbkL7VWdDFsIzR4sZ6pGAWk7w5G9vvT3G8tY
54Dg4JblTWo9f1VudyHIzqDo0KbjD8Os08Kk/5gP9mqBhDBuwaKfuia+8Ssb
CnMDAbuHSoRwTxOgUKy61+ZjPdJbLPrsjSxL3yWn+aZuwk+zfEPpma3VBsaH
FMRUjRthLT0esIbVrBIr+Cz+sLEmZcDkJIybo4XRmoGBLMmvwZAyqV/0YDtc
5wF7gI9inZ90IsKMyvpT8WFkiJFb+WYP48toQYR45yE7ozgOzVtWdaKZneKg
8y5jw4wN4BTutzSqS9ysNJjXcYnwttJTdXKXFJaT9Gb9P9uwBERytn1+ojYm
sYl8V1DddJVTn5odEviZM1/Lg35en54eka67XeB52ESfSaLKwkpI+WzFvwBs
08+w1Pavdralk7hr+uB6qTycZzrHjOf6uD/8gt6BJ5n6dppQWH2e8oOwIlHj
cjK355azqwT/LpglqNVGoAU4aH3pKvlBRfXpH+K+n7hXlaMXeS32cPfzA/ve
OF7QdFVYtNYpp+QIQm3kW91iJrCasvYjJ3GZgjG319ZVkVytrRKdU5atp+PC
2fiO2l+GxoonYb+j1XrmySZAmRbif2ziBOVSRczQilat0gwc0bf1pM8rGe04
5AaAWPG0G5JT0sRSsY+MagWpKg887WTHxbHxUa4xsmp4Jm483dQqYn65fGDj
x6gqERODxmSNucx4pMTdB0x0Fl2FJZsAYzLizzNUDIhC2HdQIUytVDIiXo2Y
/jAlibHOKkue97mzN3UeXoLM7uufFj3/f+OdTcJmZnYioY4G+T5sfFEFgwbJ
fXk5h7+6yqIgngjIxAG/IOJ4CmEf/HE19GyhSKCmmM7LxxQZJWTTgnS32Tzp
hiXrUfdp5QZXYyEk9mYEXL5C8FU2sIsyCm9kK7lKJAYxtLqQaRhBODKIWsTi
EmKbQekKlZC5bgc1xWFgKvmDuYg6+I7JixE+oZNxngACw013ZuJILI/LxBVo
+453drHDT1uvJPZYAaGFbtQgix9D84gmW/p6X1xr5tauZ8kkaustbGdLrpfp
UXCFg++japSxzoJ+LFPsE9P5R1cczYDpH07oUtqD02DoKFY2dSAavh5Q4Lki
8f2dRmZ66GOESK2YaQ2RqU+Rt8GHyYLUDel3MR1Rs0i1DvpVl68g3VeQTkDh
scYne2E0eua+7xYd4VPdNt+C3nFeVezn1e2jRMwvfXx/J7Tn9DqnVTJH5u8j
ViNljjr4++fBZkUuRcf5Gb2I4fXjrDB6PT69RFHkezgxIu8d0O92aT4nySo9
1wPwigkrZkcg9M/75o+N3CC29VdctpubiDNfY8JP/8CYWvJjLWr/b60lmIZh
w75R9ktFos+2lPBR7qJx2eaM1/A7B4axlh+KCkSK9be72JUx/jQV5y4Nvwx8
78H2hHjyOtEYNHM6cExaJDuHijBdx8abO4YTliyA7kk2M1vlQRLJaHMEpg1M
u1ALgJKKL5sI7QG57KtFgc2SZ2ViA8Treu8VTrbPkdJZ+l1t+9CS0+rtwNVY
47G/nqCtVqBaxZ3owU+Uv51Y/8iXpy3JyOHtuuZDeS4iN3OPv1M3LAfzC0kp
+AxLzXbiMTH2pfoQY3AY479PeMVr8rwqWp4i2gBPLHgY3ZmcVrfgXf6s2LhE
JqGpNEI3i3PV2/HPdwWq2RA7mDjF6DFivpj/GofRlW6rNLbx0AhGp8He1EmT
bIwaPWSIMzCxYJd/bxT5OYSABxUA+qhspHz++D3IJjurgPgG+3xOMVbShAKc
xetB7d+30p49WApRIJDGeYvRgW4LPQOpycVJzkqdTw0zpNsqE9h1sW98ugrI
OIBOxhEh84s+gJviF2zvyPAsnxk4kTe6x7P7FsEjYc0TlfEfUEwUDl8soYLt
VIGtZJRFxg8fGZaunc8VsqRo5a7igkROCAco2Wfihyv7rA6bax5Koprw9LrZ
kjJyOXNQxHM2aIAVRwfBi64P6lVvUyjglqNsIIPXecaSUl/jJusYGy16akDK
kus5AtUrslI0qlHOIam3Gz1Msl4Arg/ghmX44/HpcBNLtcSREOFIL60VUOwW
3DZiXnkyiAgZabYR1P9PfOEfwZEFWB+8AOgU56P0PQUgPdhr0S841KthKOB0
+JpbZH6rjoIaQS1z8mEM3+TNgfeXMqfw76MQ71SSXij4S8VBNuBbsVmNlYD9
F0YcAhBXWZzv+Ji4BbpDK+oZmJXtdM//EXCLXVPQ+28C8PWQwYjuMWTeGjLI
cyt29Jt1DgQ/4AVkri3fsTlp1/XFMCFF6KggLPlSEvXma+Ni1JnM+VZ8m7R6
mrr53DpZzC7vLcXxC1v62HfdZXwXfykqZmiyxflWPrxymTHZXj0AaPBIgEcZ
oAzy92ViNUepN7gAM3dctYMHhhMvjsBu6wHzPBLtQjLD+pBtJ2GdzEK+a04x
7EADDD+9rX+lgh38aH4e+ZQ5Zvmk7oBiTc+gY9lOLDPIfVZhKfzF4cKDaZF6
ckZuwRhFwBLnSbIcDJdtEOy8Dq6/05OLClBumx7Mv8vFaUe6aE5M1QfONEWW
BlLJpovPKE9N6btmtct0TAtlIutT2gvpNQ64yTwtYQZXkOyeAWfOCgz3Fcci
Dkv1TM4VzbMfT8SNFSgcoUdu5/fIwioLY6E0YujryfzEGMatUu6wd8ibgs2A
6lNrPSgukHPUy/k5Em1wDW28gEX4ycSUzBULO/RHQnNdp8u+Ahv6QljHVTDR
GKNhpCfB95wKh/uurIR1Q5sOqTyLyKDIDtWvxOb+x0Y/7Jz3dhD41bwzzApF
Z9tdgQsrNuVACrN7nyGj2uItvbyN4eFOXamwZXF94AUK71xbBzHLPVZv1hWb
dOGLL0A6OsFgLhGBqkyxI38Ibylp69fN3u4AqkhGy9NameRdVq9Vs3An4nCx
V9t9TSpOKZRpDmsZsReHpce9m+jUxkc0gY5bVoKncz2SDUqpL6HSyxPBgd+u
dLCO/5exmzRve7M7XB/kRff9KC2iVFGrzfRfD2dSwSnBtcGEzDaJVcXS1i7t
9oDJXJBvK3JNXCwopeflEBykPMT83GyikYZvJSNMPFmR47Lzk4xjBsXQy1L5
uZWwwcGAuJrdyNp6dlc4BWSn+KbbEm83dv7rJTSt9Q292sF10AF8ELgfwO9w
Y8pgZ5qPxFNghoFXipw63g1MEbj9BOCCpbUss2CRJE5uMUOgfmQvaymVSyxN
zDOvQNWdaknspCKJMVP95CsFkcW6glwgXLFgnlyrLX85S+TYZkWoKVqdVM9P
SONsFgRpIaH0STC7n1IkmGw+adgzy81gcswGttd7O2W3JcoxDjrqjozvvDfn
a6K4ulkQyk5ID/KH7OOSiLvIqaRa95m7fmIzTvHPr2NHymLtLDW4cR5dSzt+
LHsC1muXCMYqvalQJJh2bvGylwoEltBaLXZ1l5rKriyxSJDT2JqRQNME4+uU
uX+zRtuzUEJA8A8e+0ZpQ6H2Q5nFkwRXPP0pJ3SwvtAfDETbYbjN5eV/iyQq
QxdA0HTz7n7YwRPsCW932mPc9RVQcgxIacRcvzfrKWLzgnAHkje+avBxkHcZ
+aWAtUx2+z8O6OkzdzMfDtYcjQFovRaKCozQV9gU/VMO2Z1FFgm64LTloPkN
cBO12sY8dDhSdR/cRL5X8Ccvh0lSFjLPSNCPDE6f3bkNhX0lhCSa1rQcXLHp
1a73h0nFT2ALN/Lq3NmyiF4rniV83/+84W26naTYYtwPGJih+2kPn4MPtcrF
VzQEGslWlZJYL3uuoftoV5aSSdU47nG3iaWoguM40UP+9qCO3hl99/gD5blV
35prB8mQ8k9ccm8/iehVYKj+CnSQFZ/cOuliqT8c47N0RxnHq+UWdvpEC95c
VMbF8U942VunhKf+skthNToIZ3gMAe/1/5GdJN90rFuNIQJ8Spoxbtbpv9zB
Coh9UdMw2/DC9GkiyzYj1O1kAeAvMimN2kB8s1ZvvqJHICVEDyeyiRxKsU6h
0M3wSP6zZ4CocoWzbuNe3cP4OUYhjJu7sC/nyUaHeF4eK+WsuifqHHbKAItH
AC3/yOy2Sq9bXeZu0Vv3h8OldnDDhP47S4XwdkWa9C0R4q/hlP4stXa7USj0
H84HK0qGvDPiYAoXV7O4ws6DZW9GGkUbF6P8RUsRsZBwI9w6R2c1U1KicunP
q984vXLMEfGyZgSg+ZCuoFjl3v39gEC6AUHF0HIjDoLAeh1OnfX2trh5n4U7
wnudxuDP91ghlKj4GbqUNrO1B+BN1W2FjBXLItHiVtx9BZHwDqXgnhx1m67L
Z0lWELprpVqxqdxfa4+N1lESiW/ObA8ho93lwC3v2gHRcN+Dyp3Rjl0keUVa
xltuQdNUsTCrD7re0i962H5soQpE+R0KI0jCDO8Jr2FKjf+CoeW6PnKG5a69
U6DLbA+NwllSHWWpWs7ERhR54+TaAdhN465NVYIkCimWlQfa4qokjTAy57JP
elUxgUyjGX6387GwhaOJzxgRgcjiYV+vbviKmwbGy16+JiuSgPx5ZrwNi1x2
l/ZRFkj1YYOWfnBEtYr+0KdKQwhX+In4bN/rd9X+IlUQftysU7Ev8/j/Myv0
Gi9MI0iBEpUEALalfjAR9soO7sTlL0j9nrK71oQV7is9NGE4sp/x7ANKuWRE
DfTKOrla9rc80qKXZkCGB5D6b024tub+NGTiCgV83cvH4jspAnB9Lb30WDF7
5o6rjllqsgmDLp0te2C+2/U0nHtz7kxtcRk4GiOtL/QF/gD9bYwFhTjf2RYY
rs1lzgxILR3biyXJEdiZ9HxYg4EXYVJYlYGH4RLSLY0D6izpmzmpBqh3ASek
zOu+gzvFesds4oab2vmG0DCITHI+Nf0tZVGRFyrogwucEdJjiatUvKv9/w3U
4OLd9k4j59kVTzIF7PtEQ6iG9osUQYDGySEqZxCX2eshWBCdHVD+ZLJGa3WD
mV3aehhBeqvv8m3S4/hpMcv0RbDekWmWKoV5sYdmfjjoctgRJwU21ItV324X
ocC6tV2gNA5gFIqOPcMUslDP/SPytiCrX/S5GiDuJNjki3H6UprQycjd+PXz
eSEZVD52j1eeS8UJ9Df4VHN07iZ20gLLvO7fObxA0mvCi4ZjGNcZNdPBDa4b
4/8dSI2EpyTfbnW0c7BuINM2Zq4DFdfk9LejXFl4jtpUGz97Ow3sr9huDV3S
qBc4N7BqyJO5zDdHRuaKCODmrhE+HeWxneJo3ItpjGIK993wpi2CqwXsoIG9
FcXcV8r3s/pqk57WmMuDdnJmKSJexZhpvtipB6t5nVXVziM/YV+no0XrFsTA
IigbDXKnJ7Es6aD3dxd2aGg5wgJkaWltS5BPLL9yQPc4q4ZIwkgfhMEQl0Mg
SUTv3mvYccwCvbzvLepAk7DCB5ZVQnis4PQSKZYyILSzfGb5HqB8Oi+JOEUy
G/0jOwpk43/5qgkJUDqhsU5Tj9YZo9UcmzTWvxtcP0Xk5t9p16aVRuyGobc8
NyZvxKDZH4ckm+PVXCMLirKVOQkx33y2URAbXUo/H5iIz9cDPWpRThzjIBmu
zG26HUc6HdQ/gbYAjXGz7uHP6Ktoy1bCppJBv295qdsVfN5xW4BbpgTszxk3
KlxqUDaIYkg1PbkmUPleM86j2+Z+tTlzoUIhealcwsLK760fMxDMnIvePRg9
MCkkBROvK+YDn9K/IHpPvWa32SBWHZw1EdylTua+D6DJefo8nzkZUUAxe4pM
3jFBB097ABPR2+fSIlQY45rbIFsiHPHCxOJ7uVjEa23n4DSAQShKHjbdkuvL
KiAkOVzERJGVkeld9gELycFWn0liXQEF5x2ETJvxl9wzqQm6nHRx7Rm1mEQ1
viaSCnwU09ooXqx6uRyMgn8XMXFCcSQ1X11O6G+n0HfehZRCiy//wk5bk8xe
rasjLI8VCCq1dSUW29ttXSX6qYXaHkZ6QwLodBzbhmhhjQj5pPz2mJy+SmeC
Ph6Wh2sQ/8HozLRgI0gD/Xa0QQINnezMNLR4BlUK7+xTvYRYmhMp400Gb70j
jo7HtFA60JmDRysuCUTU3e4zwub5+cOixuwxf0I+axkewC+MaPQSTHFBe1n5
hJJtP0T0TpQm3hhVOAzMHBbTJFVjl4dbdFTG+1NsYphBnTdjwe8yHvNx6w+r
XfP7PqpRZM39L1SyuqvHJRzMCoEzs1HVX0hCCbvhk88KZJEY7wn8IrDPH7nA
YBvwCOtTMyPSXUW4QovsiGb1ENi3jS9d0cqInPg6wFGFUwo56cUZmXfgIL37
yuS9bQzs+pIekkkMWED+2BHE55mbhRTdtOOVLDNPItzWY1CNNs0vsLGOS0pj
DgHpfZWqIi7sbFqllne7XJ8qhYe2e3O+k7rdPKHVn1WaRqV8nQ8SM8waZ+Zs
WyUQFGvoBISI9UPEwm1oKgZtYQgdnl9Xw+YTBE5+/clTSBv8n54qAvqZErKt
62OCBRXbmIjF0ZfTftVJ83kTXBJiFM2CGJaj1y2MonAqmIVQkagTp1hrio5x
DAvW5jc19wMkW49tabamVivliGnLLrw7TFmUoG9wdF6hgWsCyYDCZ3400TCm
F5NIB8HGKmvjQ//+pIairlaXqEJb3aY5pj0/ITjkBLmL1qWfKvAEx96TCaqL
26D3hzlYw36s9AdmSVDD0S9+rR4dxnYCSg2emDUcN4IUwSRBKApHikbeclUd
J5ovzQE4UxpWZtEBDMNVkiGi9AolnZuFddbBCxfbo65Sv66pF2XteoSOQJO8
Gsu5HrGz9lW4gYtEEGRZP1NXRy5qaAweGgyhGLRaIhAzTS0TokhcYM8xuv/b
A86O9pe4i68Qgq1i+HZ09BRz4DOLwOMqzEQvn69qSv9W2JYmeEMBQ/V2hHxh
T5lnOoN4ENR34FYom2pueA09JPSftWlUZMAn6zxg5Rj4ItJWvwEtHqGRWFu+
bZPNonX/vFEKW/E6tGGSysrcEmc7Uu1zDHeVhV3JYNELKV4kkry+Xu7REVs3
WHg84i7BuGASwpAPmOLRtPkAa6UTvUZS6Vik3J0LVZgg2UaQtyGgJsqTHB9H
dMn9VGkw2I2lrc2DsbVIWYY+MPxChvpJ0B8jzEsIkpS21WD2psuwkl4IXMzS
7Vo+yGzO/b627O013JP+1NVrjma5MUy00SdA9ye9SRSCE5Ngnki4s9oL1QQZ
dOnvTuXuGpSgJaewIx3Gwqmvufbz92bSkpQpWCtKT2Iid3AyMl2YgBoy+HlN
9AClpCrAAvQa7vQmw4czFDcvN6/M7950CqGhJZKIsJsu+HCw/EXkA4KHtyp3
blhIWd9B17G9QgGVCPa6aIfdtJ0doyprKiFOyjECoOhvSuVgkB9rR+X44qas
eq52x67vefwxOdkN4UgvL6Zwg80YOOT0bMXjxqG2pwpDh9XA9AcU/67K+odV
NSVkpSZ45plVBFRR65b3yGBpg3QBAHrZimn9yUt9Y1qNWLUjjMdfaZs/8+ic
oXCW4HMjTlJ2zfUsYda+0tr6dqrhWEjcZ+EsnLp6QIvspVezoHb1Y1jxE9HI
4kzeLNu8aqq6NpCbHe2g50pbNXu2ivDFMyQircIlM/uHYuFHaPfwpLjCLx7m
Q0KGtQ4RmkLTHZwSVU/Wuzzid0WFhlQjC41+WpIbir8j0yybxPc0M6EW+D2I
0k4WGw5sf/qxpycO9ElYO0G3Gfcpnt30Lg74/Xj2DngN22TzGQ0aX1z3WXMq
AWH1ZKAxlIqnaAcMwxr5JC6WRDtSr8qX2XM0Y/baaWWJjMUQ/Wapvx47pz8d
RKxR/VfB4unw0BJLcvSErZHYFCcdmHfuOdKVFD+mUavLdaprSEvdr8EN1yLg
F8DxpDFmP04JehRUXuXzCYF8LojdtAVOsCikWJR+efShM8cE1ABd8eaKDMm2
wmnv0RxmguZHN9hfldvfVJrgTWjKxEikA97JqVJEGQGdqdnCDZSR5hL09Okg
QLEvzKLx9Dwk7etUoSkYavaLpg7kBCsS/+TgR/4VV604iqXoJut4Il4OduPy
UqAcuTPK2hxQZ/yfqZFujULfRjHMt4s9ik8krbTi19tigpW78iIEI/eR2Auc
qxcVBWbh13SGs6bP4Wi05Zgja0yvTWoL2bYKw/6eAcE93wYTR1ZrKHGYQ5Xp
GmQLu9eFhRym/Lwtb2vQ9LkQh0Udh8cvZRo1edgAmg+3rG8+g+PzvUdmhCHp
Wdad2OBOrPonj9KPdf62liDlm9Ys+RXMZd9OVb8OQIv9UayqR5jiOBRkPsGw
836gokEWE8jp+5Fi8b7Qm+R6AYPmkwUH21umjgzIlHommfsSDDbio0LkRuVf
1efRf6KTM1PjsSG+B6VaWKegB+wtx+uOt5ZU+YZvOsHLWkT/D6TdjdCtAGVh
TQc0oG8YUcu+FXNsT+F/elkhNblYNGwfGuNZRthNsNvsM16C5Pf1IAx+Bjnw
YY/djSXVRhQZx3pNUgqN21Rarcxk308iDhS0V4qFLk90OLh8QpUK34sacYxC
OUteqJg3h3Gyyjy1xlWOwBictzq9Chx9An8+O9WNNwSmEl/D43bo6o1l8k4e
pGX4P7C1NU7n6+WB9baV/PxOO5SYFc2tlBTJhLJ06suRWPL6KC9Bh3Vp9hUu
s3skJ/LWbcCdibkW9sQZ+ITd0cu6e/0rsWrO8eSQpFCFTEte+dalSnVKyou/
jGalBLwb/+c2jICP3P6SrcMGNUVZS12uihZGsl2eCnDs15U8wdXTCwoTL7ka
x6PY3PEQ7E468BDV8ds9ZsabxhmsTMAFnbftX0FDQroaXOmrRPXtj+DwjhI2
VTVXi3kod0bCYC1xZoWGl1uBLOAzVOWghC7DdMtjhMOtUNhXp2vz+tCcmUbn
2NWWuYW3kzJVslJ3bNPBYNRNDE5LJsykn9uPn7in++kEj0rM2pN6mmb4+Xn3
2umTpdpc2G2Dr+1eCFm/LcEDPDPpkTPj93wI1O1UC6VxOGgRTHG8Wy3jKa7M
l2I0BGb1Yl2+rXsrN5TwMo5QOBgU90fPVA5VYlHOvZdM0O9Fiwz4sfKqJUvm
2ZCbx8illhzIxcKmBesY74bhfoTV9CTZvvP5BxuWRVdeAqFxi/HGUJRTzMBy
DSZ3V2NWS5o9CFhG3t2SQIcfkYhnmLewhTPLwANDWk8e2uHQXAjdNf1P4eO4
czG475jzTaIDsrYW/jg7YMM9vcyq7leEV1uoTK1cir8D4CXkZGldBaRMReIK
ZGWxGoJcDXeTOl8jHdijlmsiLm6CLJ0e4Pu3Bw2Yle8hkbBlGCj0GdrI2Y8K
k3bNSvz7y6+7hLVlT+TufO0rSD4WEzVdT0nBV0BV6DeQBCet56wQKS4t6V8B
ZEaH7w2KmXJm1ZiplqmdyPG+D0SmxfpXPtZb3kwE7v/rrX2jPx/9xg/YxNWH
TC76t86pFQyWPKmiavPl7MGQBY3htDFzE4VX6WNSb2R+2LOCMeu1nqhBJZZk
S8qPrjWrxsv4J8zn00KfTyT4XvHeN5ZQYV86U+iD2xQtll1ZEdJ+YnEsevkj
JMwNzUXSr1raQDWvMpsvO44etgIj1saM7vK16mkgRI2fbF2eUK9WZo1mUf0a
SQpeGgKCjYPR4Q69MsIYIbaTn4WfpB4N6DhpZJf9KzH90I5k11G67osc5EjN
EX6XzS1OuSIKTErGcD/VFcRE1LwEy9hDycE5mksm5Hu9FX332s1Ta73zrbkA
/kjocBo8rke8jz6YUdbO9CF6rg24kEEFiw+jN9RYEMLeCgi091tbvLbh1abP
8qTLIDwlBTkuvF45GHiRVif6jHSZvzPU6kS8R8Bq0S3bN9iy9ZJDNYwnU6Mt
Hd1VYcYt7L+BaAsKMeSto/sEe7HvZSWe9qh27WhHsiB8e9kRZTOhnE9sCoLV
1RMqCh4UJO62UzrznMzrmu/mtvWUNB8bkTFYqSFGxMOzC4jm8RJTwz6Y1Hby
VE0rHVwR0quv0VL+T08PgPhcmD7a3YOYUXr1elCVX6YdzapEqLyFYiRIhDbO
9Tw4GYjF6f/Zp62YMCvSXo+uFQV2rHcXZaNSDatv0TZlGIyktInRr75LCPPe
tExM9Kq8DZEccKHp5U6ZL1nif4JPiAUYGfxB3NQbH+A5VUx7tDYNuVsNvRde
jX51OqJNn06Ql6NtCFmiWlAXv4S3T4sfknF7MKAEERsErPl1Uf3FE48g13xk
clew0YwxD4CoCcBD4idthpxIESac2zmVlfvQNpeDNoNn9ffNshVta+2r6hYz
USnyg1Mm9uOVYtI/Xl9uL5jR0yhgF85IpXFCfub8wVTbxwEmnzgXgxxWVwzV
w5iivwJ8UOlXpDi8fh/GMxIVkBhF93SVC2X+dvQ/h7Il/jyvUxcAnyis0xRy
hXxOTTWq4i95/6oDeYlk1zeD0GsZnMFa2Uog2szEkKV9xu3GDY/nq8FLQrE1
39++Py9LhEfNj//L2YpI/mnL7B/PobB9Zy6qnSQtqJVPMsmhIqiSiGjmt0eN
zcvyB3rpbJJPoOMuToK8nfipvfjDFj5uqsZKxBLnEOqD+L/AhnDQ9VTbsZr+
3TXc00enqZa8DpLmI0H6Ax66RPv/xjBCfy2bK08pmbuIsROwP6ZuSVzU6e7J
jF1Q7HfJGXmdeknhbC/ridzsjMj8BFM3u+3pUpOk3PsVn6D2f8XolCTck34M
4NPYufUNCFzjbEJI09gsqyB8Px1+NXJucL2qr2DVbze1NtimpgwG48VRE+WB
OJzUYhx4k/j46fs97taOdLlg3/Ef9QawZvrjCR+Mnapb7BPYOGFDBGuBrZaf
wXHrGI7MM3GXK7eVoTcZzdnuiu0O5pz6eW7GE6vwHwABvw5+5s1PbvIZ9qE4
0BWo5ZyfcWvI5I0zXx9hiElvXN4xR90oWd/6MQZfN/TQBWyyKNIp5S67G1x5
KmtHYgglUWEAu7u4Q98mI5kzcf4vlOhXNPmNlB4l7OPRzqPczxXFAwsGvHRW
D462NefnmLjoy+YZYvWDiskivwwI+geZqc7uyxKeEcUIbmyS8SzO774wfwcc
E2OkcR7TQZW4ZA8iLRYszdYNsXDOnjZQSrXb1mS+rT8MQMOkwxt9C2zLuA49
Pc0KghweX1CfQMFJG6cbi/nWYcay1jldw7pyV8h5izGrQvKS6zRsFRJ2TIZf
BQAlsnKUMy4oxvMPuMixiumgi6Rw6EmtX+Nz+b+NB98yh6+kA7XIHYXfPMoK
kTu/lgrEfyCieji4y5sPMffpfFyZBmEEaLPLRb6zneXg3+rb2gA9C62LeyOv
DVIwuvu46oTg1raWgFr+mUmex7AwUKB7fSts+xM6dmgomPDUgBFi2YjYCwOU
i75tqtMvcean6eKDzsxnSBIWt5eY/4xf2CcRaXUGta701MIj5fuIkExK4nCS
QUeIgIg1nxS8/RfqGxkV/Gi8Vxv68SXH3lDzKdCuWE/i7wA44BWgzkkLkm8j
DsYPZdHN8vPyL/N/2aJIH57bZGserDxmTspvdY+5gO9AMxOSCz1rGqj/7OQD
gvtvThFnUFKOJ4Wai5/8v+Jk0tKy6hC8wb7f8RZGLNNIvxYpWl98YD+1pAEh
yMY4yl6aIlCc1BEAjZ2saCox3lPNTxD5h2QWpU47Ha1DTrIzJPdHN5qBz053
SplMpCJOG91CcT6pGy+LIyj8qqa4R3N0oRifmbVFlMbUdoYC7CTZ6ldx4fKG
Je4X/k0OEhjMpCgrvJbsCO+UJkPb+AiFhN/V7dygWzTsuNJAy+q3JBFZiTx3
qRWDcIMLpWu9Ceje1s0ijlv7GX7xx0PMX9E16aUrbKeqB2vHtkajFbp/EDeZ
4wNdC+5xm0wt9VhgDwlt32NSsPtYSWjarN6MxuL1k7ByotFyPboxnCIjdhwI
xcMcLVUyQ7S5a1QQUqoutsYgpHKn6MPQZ2/wVvkSDc/aq9lsXQAAsciutoI9
AdULoKtLrgm3ZWevdc38mHDuhJZpD9asq65lVPSC5O9REuQmbmA/HKVkkTxK
ci/wx/lqi4Sq2uO+KikwnVFE3l8k+mIcVdwPzJXV7Nf0KD2m+h24oKI5G5C3
fAmHtI54oY6aINhZwcSYFXZ16kafkQSzOELivvTvuwqfIxHdo+iTmYDgsnQf
1/diXPov/KnMedkmhx4QecyXxOYUBp3owyEVz4n9vOR9c3e8I+plukiuNDlB
lUgR4Vc2s1r2q67Ef0somQSHT1iu0I1ggnEdyAhybhbHu5TJJP5trw7F6gzk
g5/i30sMZuM7e7gEA8tvgzqPjy1lILSPEA9Mu9keDk2dw2AELPHVdwJbYqPX
8wgpcLQtneNnqvRfdaF4+grynECMT8FSz5g9eS+1kvvPdq1KMP6fplCHFWPJ
BM20MVeA8JqsWFP1JfzvjCLa3KZ8y5N2ImquyNaZBmKfFQG1xaFDh4B0yVn+
aI+IJLNXm1GM7txL2Z9214N13iL7RvkHogw8/JZakR176cp5WFKieW0QynMJ
iABPuuyzIGv4J2GpigUZ6nk74ABYprBA9Ax9pm6ZOfcN9K/fjCaRkK1JPyCj
QI5Ul3TPcEs+wZ2GkUoRGuL42k4rfZxBH/kCkU8oaHeZTZRb9Zg0KnLpnKH2
gOM2aEYFhhV3TL32wQ8kPTj8T3NVYeGnMfXh4JkbdLIXmL36UqXEWezs6525
E3TC9wgYU18SXLrBHdhSiUu0NJNFHCOzDQQTnz+Z8mfj/yoXg7v2d+qK6sPV
IrLUTc5aUO2nrF7k2dH675c6dXjY/qvSYosfC7L6/YZy0mA+lcCx7UmHd2gB
Qjebpa+8O1Fy3ji0a3E1s0Kznp+a9oHQeMijZ+faldeEmORCpe2cpCm5S4yk
/ajQPJykVHEn5MZKoDLbrEpGckartRw8zCftCKtL4h8UFUOUVMUvXWvheCkl
0qiknUlf/mL76Ey8Gj5brzjTseEKyPrlHuSv5GJNYuCHoU0Z0iFoaj1tZgyN
o9yw3lZE84e1gHWNulHpfqrnJXQhIEAIjniOQfHkaH4kAoCifIz81MjNlz5Y
WuIPEIH2FzL+prvwikAARTkT3I4LI8nEw4f8DdI5wGvpQt4EPkiVC5qaFb3q
C7v4Mx2B67jUkyJeI0qpD1elnF7gI/ivG1Z+g7EuaN+YUjKlU9LU+chmItVs
bzwAB2QeeGTPTVyNDKc2vW+KV6nDW6GBn44JpE+ukfRjYNdVD/i/iG52fsw0
fTuoeeXmnkgc8Jjwhn8PcTzyniSAi6hmr2Ku6Ltrk6yCwK1eYlBXqus9YRhu
cqh/bQbjftWSf66S2ONuKU/C3aMdrpgLdixCz8NKglNhCnviMjNys9wz6ncK
xkLhu1j6M/5bC+/niL3ddUDq/XKP3F37xt1pNRGikjYECwaV28uUWDQ+IcEX
l0YP3w/FrbDdHpKA/q/3KWTybxi8J0dWFhsdaJbCD2NBthrlMsAhG+2rZtGe
yFm5PNDvlZo2l+QqhZZc7rl5i/U5c6yg4eRanc6izPs85Wt4EjZ2IELd9McC
QPs9oP0Ep5yuwJFi9AW+f8Z0WKHexOBZ2/4KcjhgXeh0BItZIRexgxLJC/MD
teuy+vITdT4rlbVFqAYj8RbghX8DqVxjg0wYIYxvUg33erGQuOAfAnKyHX6W
zuOlHJCYfbMDf4yVjAWYZaFrT5Kj5JkcUsNFHGa0bp8aWxS7nS5kAEIgohUH
NGhvUov0Vi3a9FCfN4b8YLZE7DSPCV2vxfcoa2t+mflmpXkFv8LliJ1eFfrd
l/c5duz+6izqiprb3EQtFLsQiQ7PWQJgXkxPjG2JniFN53v8D4CyVGKLz87G
r3AQ9WI+uOHZwNAd5W1GbUX4Hs+CGOk20gwVRQJvJ1rsNQH4iZa6iJoTCgoW
XOVav2CuI4jTmaMj7HVlKLXuOfAmF41nftKYl1bDdCOeoE5b74SC+MawCV7J
uDWtCa7KTapbGMJnqUjo1I9mj7S0cw1td39ptWyma+zuHSTwLI6WEjwOKzPN
k73c4cNQtr8FrNVBPvz0oiOE1m/lUb6BUPJPo4HvzlY9jc09WP5wMFTGB1aH
7rZ3Q0guga+1Sr0RiJyfUr/O3Zht6Lmu/S5fShPZo8OYyCh6++5lSAaxzxnY
6xFersjB8/5W87Q4w2dtIjhAZXZiOCvL3MgZyuoPKuRpnOpTeS+Hsu/Low1P
zTnRLC4RRSL0L6ZVl92cBA7NGwjM5mW9sF8gK8PFhoZ/TppKWzBfalEODVEj
Z5RkwSlNsqrMj+zG6sChnVmueqqiH5X3Y5mXYKkAgyXb/iL0lPXhJuJK63iK
Yre5vN/alW2TJ3pBqfQHCXrOl+erWGqgUgNgwHV+gOiSUti0KWFXpQjG+4o+
phAFIskxkDYvGTvMEeKeyBTScQQ257LvVzrYWgqjp542cR033Y0BPukaUEuC
VjV3EmyiZX2SUHFdPs9wNBLsX0x1dD0qHMP42+IR//L8g2MEZznUgFpQ0g7O
hcXnAFVEQ9aVcu030wsM1ueXFG8OkJlGEqTk9bzjdfbZrey2QvSb49X4t2Dd
FUadJ/nf0eiNgGoHakJj+1zFZ4OaSUiNpSIQnLEtNAyy0rixPD6fjzWPVcCB
6dCq8UqAYidoINnTO/tvXJJ7kJ2Ipgh7zwfDYVm/xFdkuiOc5YFFl2K+NwAY
lTL1XnZA9pqv1IYlRo3dBVrfA0u9Kb+i27x0bXc4kX2fhjTtJv+tOdKCgdgC
y67X9aEUHn1jsYuKJ4znMMrMb/8t/UI+5rcUyyX+EecI0/kMU97x6zUkFh0A
HFjZV/3edrhTF78jXV9jfVZvfpBvwMLTf2oIJVVj3CC1hl4S4kmoFv9j9BWr
3/9prJHNuDokEl2YPkrLbOrhDRDgPaqPHof9z0Bu6DhL7BFYhBiuCy2/Ngy+
GtqM7oCdA7pz5L3TdYIAI+o/pxjd8xEc0zvUxDyteEp9tBCjHdK+yFyWLETx
yiTgMeto9+eFv5m8348YTLhZ9SKShS0AMKausLMYmAOj3N41ybkAEdth8MX5
qZD9Zem8sr8/zo0tURyKH1DvvH6lexAqeiCM6nl7re5XoxVN4XrYMP8vR9gQ
TTo52KpOR5tkwt7a1OTB5vS5+HPcYC+iQVhYx335oTStG7l7UlYnjmgT/Opw
eyCD8yjsc4dYzqX29gbNHFTlyZEhKv///e899mrV9HaZV3ZFYLEwGRutj0x7
yhnkDDDLxLZpACdueFfQ2qx+qrOd1N3OSph9ZEydz6gnEeB7CV/pPjkTUwJj
AnByXhUyArrb0vl1gRdZE1eHpoCsB4nA84VvAn192Z80nEfyX1s+2HLoRST1
pNhdDJB/7POC3jM9sErUDo9UdvHL76zGKd7RVus4Og9xUcyG/D4aIc6Iec5j
f5leWoUYv5dFTPEq09TrSsBnSjpTaMvlyObpvZcK5RR/S+jF2IICNZhr/mPj
0cMgpvVsncmiPcqnLHEFzrOTc3dIMklH8JSeT6iOec/fOEzvgiy4IjuBeeDi
b1S0BVz5l4+UsWFTQNulKiKbGsTh2qBoO/VtY05j9jWwNgGMpuXnP+DXHma9
XoT3DZrlcz2MlXSfJoJpwaC/MMG+AWeFVvJ2RkJwXUdtdhA3fJqniManaXuP
sWTVcT9ZlU90CWBqnISVpN1VyauetGkwyUivKPHJmvmshYUstk+Uqd2GgW7Z
kHOJUesmS0jRSlovlHq1J0hNlW/7w6aGRiKHiIMBJVb+yBds1HYvvfntQNOd
Vb87u4Q7QTNsdF9dkDtd0HKuixdtjUQ9yNovrgaK7jEUiM3G97ahET92ve3D
sj2Jj0MXLRypj+BumkxELqeXxXZs3CiZ1x622X5+gH7/Q/GQUGqMg7s8aAHj
RadzzVKSAZSPzjvaD7aQZJ5XWwCh4PzOumhGMGkteumxztKO44ImlKcdBsiM
XtLdVjd1VNQG4tbPsWMGSBjAYmuoKkJ6yTuAvAxLAi8ZBbjburN0gzQKWB3e
L1VkZKmKY1lMM02fwPdBy/v+pzGnbvE1iVzIC93/3RuzU3FdsP/NEZC0cf3z
68ejZIbZlXQcAkA9aUrc38S34AJlAYP/ps+EJ+qdLvb47EfBdLwlTlTGSLYO
VHgrpFz1b5ep1mmQ5q5OW7oxPubOM/g8Z1K9B6xWuhAp+ES1VsWzwlNbywYZ
V8FALz/bH+k6hvWPG+sQagwp7x94AMF5tN+cUyVLuOJblq0o1kaYWqolleDi
/S04NhMqr8SVUgPUIe/yesCNeUE1hvuhwvH996qU0wYhb7Ni13CTk/3/u5WO
wK81Xb0JH6baq68g+Y/3wUKCkYJ155ufgQaI9IGCi6IpgSp2cuLuHlMVS1QQ
jQclMV/aWAikoAQRwnSZnRYdv29emzkU7eX8D3qSih9llQe2Qm1MlCjHKSim
UQbmLkIRQIPTe3VoGTddeFFR2/BpM0Uu8/xRNZQoaW9jDm67/TjBXt769dxT
ViP61qSTaAKaDWTltZebPDTw7Sk/CkYAXVlr154K+kWSTpeusQBw8HH+avv5
sOxC2yaUBEs5bf0evr03Vr+BxL6t3XN2OMaeu782OMUPAJ4NHZQuE4/7hLTx
5W7GkQwW2g8Ob4EoT9EfvNIwla0BucDUkbzmUpYtrgidXqrEo4vOYOquy8Vo
xk4VIN20v+tOJ/qeiMpbW7Qj79TcoLuqh9imv94Deo5u1D8OjHpc5Q1ZRil7
SF09ztKBJxVCNJdw/HopXb1uQdoW9pr7E8fBLbGDO6fzfibZEiVl5yU03kEN
P8iHU2iCKCfcaxU/mfsOjPOTXm/g/Wdn1COJXPuyq1UhSwqEjci7sr8r4xcU
80073Of5zaCziXM/SWKCpH7wa8RK/WARUzp2Sj9KzFfDHc+DwFkdzH+by3VR
mmBtmH1Cf1A+IySycqBEKuhfJBTbJbOrqN6ymxE5IFy8FuS3lE1Xi38bWR9v
yDgF8zY93TeA2Ib8VlG6Ka+2X4N6acubowJcMZ9fzJtVBI3AyhcGys4Nlooq
K6l4petLpFhPqULn27W70vDdF8RpMY4QYx7oXtRHxAoBlvu9z/XJr/eKw1tr
mt4W9WjgxfsxJ/SIG8OnoMf2WnhCHV9AIJAu8/jTlmAT66VUlxGrO9QmkYjH
6vSGzl9b8Kgc7ztd0XzOCkYiOe9aXcYJrzN6eZbhYCLVqek0sffmNoHr1l8G
bL6Ws6m8lzlY0p/CD01VJiugLFPOv8poJDqFm8ZmoapGqzxn6MHBxT60XsQu
PQ1j46TNxKRRwvPflzhAinCtU5p8BrR3ryr+ZkhQbbzf5LQUvvCOgplf0Kfy
9JnYgJcVC5EnzMjdOEzGjrodPPbovb6R/DicIBUKpwXumV0rXiRyXGkn7hIN
ZQwjYq2nU32JwzHWmV/vZBO/PcVxFYmAv36X1vXsjvhWaUChixzNQLvNORc7
mW06xpioT5wR2t1dddgBPVbuVvsdwA350CXbPhmIU6dpl7UyE+uzcwipn8W/
ekur5Po5t2pOgQMh1jwaVanQEu9yQ8lYu2/v76CFuW/YPba8RONGa10gkfzU
qdITkZGh9ZQRuDje6/ar7K1jAPqnVJFknHLkdAJj1KJtkXnyfxfzylAy4UW7
fyWIrSG89POtCjzhbJEeKbVa7kWBLiJNxxKw8g+t5eAAlGAudS9oN+qWlmWP
ubi4MLdJKIs14TMKtqPy7Eqfc1kWBEJZfcwjeMWGRe7jcHvp8VBY6nPxPGwe
LbN4LsxoZnO3U3jJbeT5+MnujytZiArAdKITOJ/EV96PawCpREiHJMeJ9M1g
lvW0e/DwmUEO3kbFkC94/3NPLaWc2V2uCHEBrUj8LunRnss8E7lAlflhK27j
h9WDAYFQqCrxaaYe8JA7/9mCJdiCvjv9Bnn4SO/wpTaeyxf1IQo6FPhLNgn8
Iz03rqL4rAzG62g4aC9AaQCvOmc4LkaYo671cnIXz4nT3Q6vSDgnYtYaxaEd
Fg9XhmJEEDvLTMeloTv3ldok3Lmidgvy7LgjO+gsH2MZd3ymBNHUxbDynQSS
fAXgTirSizBLtRyEauJA1OxdpnkkWI18f/5ANQBRQNMBOTVgkvmV7e7HWX49
sZ3l3qf2yb7ti2b1Ivtfx6KNktvqsfG8k83Ao46buEIccmh8/pFCqWMyTXpa
/1Zf33KwTfx19a0rRfXww9SAX/RGAiEatf3zB8oU6OWqcgqys1dZpRlBqaOq
tI2a4u8BAYOnu9x++6jcNOP8h6bISbleL5GpMPKDyMD2IsjpSQQmZI1/3cdH
xWMDj/88NHOYQCah0IJ9bdPOrSKmejPjOdvHiKRP3zXzpN4C+io3p2Kciob1
GwrtVGvZeCPJEHnUbsYDKHTwodXgiaI0ONrOAQAT3zVze5mx4S58VRT06riW
PiBbWIY9n/YQFgVcyq1ayqpZrKmm3zU/8RmPTFa9uWqY+AkQF9Du4cnpIH7Z
tqS85ycIP8oXrCraNWyr6Pc88EAt124S+jc06vbeuUf7s3FBe4bQIZNmIJkH
SvV5o6ZEz0ww5TOEHC7sGICS5OweBKyItwlpNJOcPo20KPblMYyijfPAORJQ
4W8fkuXkkegdNLzIglxrKo4hMoWOXc54Js9MDFLlIJuX93WJhfVwkK1tg2p4
wP1kAxph26Qp4VYD9Wjl/tPhh613Z3N6MWmOC4dT/DTkQo8Cge8OMDk/HAGv
aXEgT2c4rHCW0mPMybWMaOIIpAm7ApJDilmK/0VrPsBVajBED9jreZIU2t7e
8C7cPhl2d1E1X9Q6Pi3nYy7+08Q8WkTQagVGFVDPbZ0WkXSSXVOAONYCRmhS
BCpfZQ7gmJ78Jxmy28HsTN5+U7+YYFqqNZwHL0TYAw4ZussDGaBbLvkmaFDc
+bw6eXE5vp2C8iNHOObYo2ZeIN6QJ9is1jvM175ubSB/Zp2IvVMxBDoV7CPo
hbIB3R2srnFJnGRGDopsuziuleuAsDKEj/HJLV0J54dybm8KeLlSQpwdwDqV
xffKegQzWmWyrJDlxCWBj26CitvPZ9GMIW4ZNCenD8V0gBlOvFiB2ZcrYDu+
CFE3gPQ5VP83b6eMquusAatYycClb9YCt4b5ym5Ib8tyn/UKt/IrpwYMZf8r
avuArMld73MRzIT1wGM46Vxlp8xJ3CNX/pWq7s0uX2AdoZD4DZ+vV5s0MhOj
4jK+PdZHAQDuG3kAvWLvf+8Zr1LeIeHvc3s62QQAEwPJJ/6+6qQLktmrOxia
FBVQGp1e6rdFFlVNacgoQ4ryH+28b9CtI1YYX+mAM5ejF3ZCCYSL0QvIOnXo
a7b7MChQTIxEAiR+mvxgmoSF0EN+Z+05I0+uYnTuF2H39RCMZ7604u7N2cJy
h8muJ4h1WnTCkunYC1sw/FJXihopJVxRh6akJeQiPA6uWWpeRYFKVJzyj9Ro
CLAyfAJOWOFKdVDG72K7xAFowsuNjaw/JrRxHuohWS0NKTW5E5mLC6eZ70h+
zWHuc+OIV8cElIrnsPh4SnYI0LJgNORArEtBWBBDsklIgCGsKN2IQhF9+E+Y
IuU1XttlmheB/ltwFEiXvGvGUlNLmGfdwaTBEqkWH3dEimH2uR9EFGLn5w4W
KA3Un0G+YoOqurnwFmlSCRG6ZPD0+eAqCfPrujQmNpqleZ6eoSL78OKd5kwP
eLOIBqwLWFVHOkjjxY5zOK861hnszxZfd89M2XiBWRVUzPlm3B2y+uUmkFEZ
A+KHwe2yaS9xm0Vbc72vx4+gXbxAyox309qAnXIK5h40sYgMdFdpt4WlbG9g
4p88cNBSvOgy8LvKtG8icTvf23Gel6RZ31XEUtwWf+IcPiK9zLEau+rvsION
L2PWIhgY7aZOODPlPVcM3n+WM+eIU7z+uugXVHvXacUrtMiLiLF8/9FfnIyc
wvkXodJh86OVBNejwGPplA30ggfxRlgj5i1r7Yj9Mw6IIEHGtr5zDxlThHxn
PAy8ujrm6VmVvkv5+4Q5arPJnlaBvvpq+XE0mEri3QSM2mZDTmGrh69eNvS+
wNmaRnwRbY8bh0YkOHUIujLcGisCTSYwuSSnUwQ29WpgHdpCm32Fi24KL6xx
9qiEG/alnh7yBu2K7bR+suae0Pf0vry5kG3wIUC/oiA1Sr278seGAmTaP6NM
2XQiRhY+ak2Bh7JAI1rHzhh8T/MZfouZVxLedVdQiLtuyUyh4BTxZ0Imj1Z3
V5g8yg4vDesBb+cyk2v2B99jeP7EUAfDUYY1tBTp8xLAV3rBu9DQX4agkcpC
ick7XBtW3wmngJmLk6pdJfaWbke04F+hOeEREK0uyfPtaFT9QhuNcJc3yGV6
YP1EzIwlaRgRYvESETC1IPrEDE8mu6yVFQHnKllYZ76aTzT+rAt2pRDrikSk
RCtDegoOB4CBijAaUaRkbQGaV/oV/OXnKq2bP7mK6nX7/RGKGicgcyHaP+vn
ifvi3gAH+f28JUoZ7dBumaHnELDYv0rtsUw94dCOmVfXh33tgqsrGR1NDEJ/
FMC2+TDj5KJd8ornbHhpyL9sASLa9mW9o8PaMB4x2DLgpq513AbMOUf23tRD
zysOKXAAKXZf4e8P7cigL0+pP/73T/6DYvHUkLAwqTsSICKlMqgXZTMO3jyC
DGR4ZflmkPZlWbDEm+9vJPBlt2cVmtHhpnGqSn8k4HVx21gcNQXbx+81HLr8
UvZDVsGDV/wN6KZ1GaHRGLgzOmu9Gvn6/aeErS5ZbfdwZdzOaj3p7TZoh+Lm
rrWui5yUybeVpD0e44Z83sbfrmqvbu1rGTlO5nQSn461fmlPwDSWv7DcuWf4
UCZj/HTNVnRF2n/1eDuUgFqQxsJywJ8Zkb3obGxa6CyfUQtgS++oOM1/vs+p
PV0x0l0UIe20JxEO9F8uPdRg2JP8NWidgBmL5ylLBB9ZS/FwsDHc5C1E+RFm
3dtV2adEKDGFI+UAW5ZPetE+QXZyTH3n8v4kBCY/5umfqJLjmPquXYxv+Ird
gnHos0eBPuZTi5wZ1oDivJiGbT5Tmqgmqr+r2QHAs7gWZY8kvFO8MPJgHQco
u0tf3qhe3zNewQUW0MTdhvQg2lNdbEZPYlQuS5ZxDmgd1/sNw+1hpG6uaCcv
+GBpwHHIGARrlythQvv8qLmgA9tFwLZ5ow7kK/Y9BAIxZUtGzk44nJ5hgiIV
XrARnrVJA/dLQeK+5M5i3FBbhds8UMyINU5C4fRtRMig/hzOXg+xAacxw/Or
yuRmgsYyahaEVvsJi6Qq8eGQu3ZrfdoNSZGkf2Ze7SMJnIfU9SlFxHZo+WNV
Af84gEZlducRhCYRvaIW9/PuLiS+4W2id36q8cAvSAjYTulYqEFSYHAYLL5D
6KJQR7s5BMuzfhjBi6u97XTfK2d8PG199q2QhwPbnBxSk1BsDZhqJN3jg+hm
J2Zm4vgupsNuX1lGOa+SBc8Mlf4BlAMuUtlJ92D3lXZVeot8jRXHQncmBew+
76tVgaarKcCw9FxCkYxbNT0dIEW+qZw9JWikiOh3z0k43aDTiAGIJyFEc24Z
XD9a+nt27yzQFfXj17KQnkNCLkHKdguJnrn8JU5WXeB5qG4e5xL0IJu5liHW
amJay70wPkhIKE/0cw35V5O5nR8DR/wDOM9GP71B+//D3X5Bv64uyeGMCXIQ
gqKY4Eq2mYcMG45le++9I70E0kg7rmXDCoGS9eM0DiBGyXA5rvLIwezg3AAR
mIZRWmlEjM9vkYndwu4yXMqO5EhUo9KDgSGOWhkMZ+nW39voZCndM5LVf8xk
bkS9cpgk9Cg6rgUJTPj0DNFbtwv1LsHn75sEY/jlm6ChT+ybmIyNWFjIKEBJ
eQ82AYkCqExbtuOt9cBjh7V5mMWo2yLupDNxgNgCqXecGskRzBejujCxb/sf
JSStWHKfNVUtG6csTgkP6TNI2yS9O9VJXxNlGtWMBIvr74f8YsHzjivMUz9K
YLh+rtxiqE8ZpHWDJBoPRQDX8DPjY5hfxDY25nabIbc4/Yi/kjbPZ4HbrQP1
gv6++w/BMzO4BxER1xT9WWtb8FHtEuPT3R/nixxIX/fJQvMErp0eTZ0qvbBe
D3mQExa2zByjFhhSXl0WfdHh5i0nX9xHGQ46RwYJjiVrVeXyprW/q0VMc4jZ
Wn8hiNg4z0vTeIfjK2y96zUw6rJAUAULsUUXDg7ilGK4d08ATTSL02K0fDdi
HJrImS3IxzoEickMlzS6Xi+7dsmVWwaV+DWMku8tK52DugvuLk6Y/m6/fBt9
EBXLEQG+U5NwrcDzfxHgAaXOOww0B4jjvUeU12UA7VtACfJCKwTP5DrC4JjT
kQP0wKsYZyCSb+b/wp1ep+ar5JpLnNbTQjflq/j5/FemFWkQmw14PTU3fof+
lPr7ncKvV97oo7sQO7k+1so2r8nm9APsjRNkVaDdd+WtVYVbPNUlK3uDiIwe
1ZsVQu2vO2r+DZO0aQ28u6K1RKYHtGVanMD/ry2V/S1s7O86T7B36Y0xqof/
xyzdewTqdI+Cf3BjMou2aPV9Q50n8d1gdXGZxWP7/BZdcR+aXY/qnIVsjj9K
CW7QN699pPWw0KZMyadShrMy4Qx/VwOyU5j/CZgK3GZZ9+EjjMXjm7BGf6Cv
WVrbNK8lp/gIPblEBjbOkirOwrHA2lHCqG9/nQH9B9LtkgIWmOsZyp4muiHe
5A9yDnt+7Za/0S//kPrri5GsdndtEbe2dOau3IxERs/JBOpfvQfUkE42wgzt
vqGUiqtTbfetqkohMgywJKVkbltnsvUh/3b4XkZjtJzKb+KCqQOh3t5qiCu5
fdxVC4dE1ldl1x00YRUEvBokCdbwvjqNYCKwQ3M14lgOT4g1QLOWFo+GCoto
gK5cvBwDxbki69/pZvAq8CsaU/nNSs1xHurP0UmOGkIldyif+X7zbt8uppu1
UgG2ExTvyyGF5weKsqjJ/gj5JhaEEYwff48DwMnJs89DpN6+2ZsD13rjD50t
QeL37BiZnKvjLI/ySEUTYZwcmfzWmHvK8fPN3dDbEttR25C9mSnuq5kfFZg+
CUgrRowcDLzUpEt7YA8hh1+fTqEJN0sg5Na3e6bpJVIPNT1HgstLXwf0YSBb
5oOHE/Ry6WR5G/c6Jz+v/zMKoBaEfuZl6ugRymOxXl8OtQPPR5ixKQtCgMTp
7Tz2orKixeLt7L2SZEnIuxyliA2ojPVpTziHu7ZSoeux4MmsXlbdw1k7NmSQ
5JMun4XP+sTo0Fu0Z+PMpvb2oMrr33Z/oPYGv01mflkQny3ZMaLs0rgb4kWC
9/cQrIsu6c1eobeZkDuf950LhJYfZSMyB+Ok+63XwN09I9Xt5qIH2b8BJzbx
a6xyyiO62E4M1VwKjbXi1Cm7/yoKmTVzrEee8QYn3ExgfzURXaK2Ke7aVCw5
wHykl9S+huiVW/uRxakHxVhg0Wu6zBgoneRkwirhjTXiMRGqjdnrN0vXijrd
SmX6p6Xw/B0dmTvdL0pStUVTlTm3OAdd5NwBDLdQfB2dUz01+K9VURUTI9ZJ
mzfTjEmbcUTPIRLxFMKvXMIukWKUtNNmfMVxT8kRbDmsB4AHQBn9t9w176gJ
i5oGlq7DALKN3wnU/nj5eoHx3JVKCd62NkLx4fqE9NSMvVWCXzeH1lBvmJCT
HNb4VfCRGswYUT+DYCrfttUpY0x5bZKukDyju0+vKIw8iSZvnOAReg4Tdl/r
+OHYmvvop96ZId1zvO7fqHBgE1J1wpGXivQhduHpQhHgKOPoHUb7mUqddnXR
s+DOLMREk6DmBIpD3mqNn4sjTI3CSUWNhQ/nh8He0ZxJFguZIH3BlK6ctn6w
8jlJ8nJAd99n9dqvA05zeeL2DaHtBmGZxRc03f34y/+dcR+NIx54OzxiZMg+
4alpTBJCOKNWnQiTIeIozerVe//2qtomb6tucFIcrfom+l9P2OCpv33i90jU
ThrWrm1qyD/xMDiQmMyOeqWPiOKQz/0bqR1XgtlLD3jXG84ZVU09V3Vk83Yj
qR/wkIRcDpdfABAuxIH6D6AScFNAjRs4UYYX6rBz06TzX6TKP5LbN9jG3AVm
VJTPNJp9o+/TUioPk9VsnV1Hov0V3SPdHdNuVRR5/pQdfcb+cBHd0k+b64vH
nRZetmh2RuHy9HSE66T2sVxtemK8MJXz7SaLdm8BG1Qi3wYr9z42QZQWxUkO
ywwS1EKSx08RtbrsXpf1/DY4NMbQFe3FIxreMOP9bUZaCtyu3cU0rhYUD1mR
Jv4XQ3VYGmcUJ/xaF3EvXYo+aq/hd5iluvlwM9t9S3k3SsQY3yXPJKT8HbIX
y5CLRHV2JOVxjhbrS6hZcnHvY1gChTZ6aYtwj06PvdNFwOSfHO19O34kPON2
f4HdoXgQQ1By8ahb4rCs+JPOOz2ABD3rupuiHUFXw2Ld+xhbW5QS1ooIy+RJ
yLdIQfNFSpozhqDo0kFikOLJ4gJLCPtoWThlSLsqSZ1D8hGi2XnXnIXUJnbH
jJr1rdM26sMopWLJqYfiBrzGjnzw18WT79dpDYyH/3o21sGJ6pwjx+r1AIju
PvYLkafuUPeTwZF5L1nGKXGEq/mHbvgF6Iw19VwwbD2QxPVtz+7oDJwi4Tcd
2+Bygo/kTLz7pzkccUUP3Z8RZNalQjWmbHdW3IVOEZs1YzwVpvRCzsgnsDAp
+Bp+q/EDlrsbq9hcWnT3haXr/2thVVt5hZdUfTpyW7G0BimlA6u3Zmn55rnS
ZvqHzmmn1XVnFZ5ZcibWX0QZObvzrmZG+/VLVoifDX4jeyZlXYizaP8zsl+p
U14rbafM9hn8BPHOgLBb8y3qCEbvywm6wekPnQcgyb5aK/4Blhfu2qeSmFVH
hwC8Nr0Wkz/Ec8UAeHWInlTssEsyIZr6c0XAQLQU6QqrXbdMzUrQA/1P8DGd
McuApQLSAMxPaKJWGKlMXf+V2V7s6B3IvtYcqm4qK4rJ+147e9/s2bJdC1CB
BGqR4gx2HPMSgvjO6uLkRbIeK8utnDH5WEQ8DcEfMtKhz74XTzfsEQDG6A3P
hAjoaI8xxmFbtI13CXZooFUQWDQVODHefrsIwHz2sWOLrin6CWLw4d4aeP8T
MrT83fVQ0HkoiyPLVSbq35/j7cKyIgCpjC68dkIosCgcpD+6utkiJUDgcE/1
Z6RyuMjqw0+hsG3CoBm9lXmRsfMFLQhQ7AnbR++dTfvkX00r1d9zDI4S3dby
3QSoEnMnLhHFAQb5EyNO9fCnkECLp+vN/Uu/Rw6amHoy8pof9zRvTOltPpM9
pygCUSRMW2hzeTvQGibGxgIiS5Wd/ZkATQntQnJ45PtdR+7YkFpA/PxoDUAq
aqGj3RKMoWgTf0xr4ZcVgHfkFXsy7EWmkCVIlXFOZDHzUCckcFOVROpOFYhS
a919xgP/rNwTTfGHn5TEkpAJq6dvaQ+qzvNeK2nSK6BmH4JabnpimkHLNqLN
c3p2Av14OIurqj435F2NyrhN53hQpB1LZoN8T9RrJpUdq1UT/8qpJH5Moajo
IDaX1aTDHBgSP7TII10SKEQY07DtHYGirl7xW3v2CB05IPyVh+SfemYVz9ll
ViUw3VLmqmncAaPnBxRy2KmviZg0nr/RAcwJ287z+xwNj5rDb841FGksAAmt
nbQqrPpOVpYk/iSbjPjDwb7F9C36zYITRrb5aYzv6aCwc+2U64xVYWnOIzh8
FsLi3WuM9EFiX/Jq4G8koqR7n+bQq5NckarAGafUrAARrsnrO9/BKXlSjE24
3xvN3zah7r8tlaBGDjQi7L3wh75psSaS9zI4WzrZS2jygSpGH5aIw3/tYyMb
dC40gjresymRczIhOBWrBs+oFKb6MsgTilv2RU6BzpukO3aPlfukfb7/mnUh
Oxz+sVwQNbT+izBimSRDpGIomVyneLJ+VNi6YrSWrRa2uB2S1KymRl6Yb59+
QXeG32LIqMyWjtdEFUZuPXDPDKyXqRcEy9yaW6DGu/yBN+xcdwVvxLacmdLJ
arAfPv9anVf2N6XvhlZZlSp/XJeL2/4hDnPzyqb2/5vF6/uJj+Sq7WAXi/Ga
y8Z5bFmXDMQKhkgMzhCT1jO/TT1iPnk8QyOx7gplb0cHAU4N7k/b42ZKZ234
51dSFuAnec98L2pQAz/BN6g506WFGLjWcBTKhk/cNZvLm+tZ7QyRIOmMX7Vi
rxRD6gPIzh18iCwetQlQklPxlB/dpck/5L3CpLfTexjapIAEB4Eps3yDvHBH
KtxeA20RPXhXt9v53E/D4DrB36yBOUaViIwMxRXKhJkVyi1ApQsM/Uq4pDIR
r/U6X7gPwS5AuqZta6NBWx/R3AaUipVrxSXA8lpeipuiwWms5687WVhipe9j
n6bNZeztJiWyB/3QpkapUTR4CE5lUT1FeF2XYVJJOeXCsnVyab24UUotbtV5
XaarwVzElJGP/xMX8hJSPEW1RukKFNJwlbBxJ4sMd///R6Sf+1gF5bIjlGKm
JD7bCBfndsW7I18TGNuBlRNAZuZEpPxkp4L2N4SX2PtEOeHzXF5quMRIy784
V+YQJMzUb3vU2jCnP1so6Kmu3qvE6oQF9yebfhpa5LF5ZvIVzJnypeFk5jhe
uiWmG0ixTnZp3lut39c6kP7SGZSh7UmP0/tjtpic08PyFXuMEPB6kFb3QbrQ
YQCkt4I+FtUUJ8Vuy5gNxq+6ufU5t7Zs+w88eJEzsExMn/78iVIA6O++h6X7
vEEx6ZHxUVJnNE5odmTUwV5AXoybWtmxgum3TTWV59r3x4lpAuSIG2Pr3bZ5
A2mgkwZvM4tSFbC5VY8dLXZOhq61fZO46rzo1m00NiOAr5DNFqjqh1O21P+1
ED2ROZ5WwGPecmZJWVzX7cR0qnXaefdMfEweC80iV+7DL7HO1vyVIQ27twDm
FIE4ceoq3m6nadEO3pHE7OIn9ISRkxrflWEY96+S20VCtT769gUiCCscLbM4
0LPKILRegNfubNvLsEIwgZ6IfZykApNlhbXrmaMCbh+Fmx+oZ+4MLv7aGb1w
B3m4Tx/2Afx0FV/IhLTi4gPmjquGX4TkvkJnHR/2Bs4cnME0o7SM6DWoYPMk
80vw9x0QewtliCqbDE+P7TtkDSxfRPvLpw4uFMRdfh3faIz52eLod0YU3FUR
KBPz+0J2NZTZJ/BaYkOXO2KFkHudzaUe3BOtVlzc6Klkkp/yREp3wLE5ALkN
Mg6LuG4ieQkluvz+5JVFSoRGHXcuK5YkfIFFFMc00pci/hrgbeg/VfNq+4Kv
OgD1WXJPZnW511epzeQetJ/yAKhrQlfObuUYAZWsohb2XOVGRrTaQ+/ZuZSl
zSUyE6LRoAGH6K04TYc7zsK/XHtjDrQo4PKIX5gNzkunIOnNtAxmO5Z+0G9Q
tEBbDZek5GiWryDhKbgJMb4nsQ9660pKgi2HA7+LuDpAQ2S+uE5RPsL5zGiU
wb5hUuEyZ3tDE8flb+hVPdzdm+yJvoxS8WvuqppCj0KLrsyOEeed5fFPZMcs
qbY15gL2YShTWWoEIjW9mMMCFnRM/aCWR+393noZkLaoZS/fEk0lwBNzPnt7
YLWlPZ+6Ii7LCGLpZWk1e+pKoI9UunJa8oheeccHdhq+bj8G6QAuZG3Q+QsJ
QMoX+n1CUDTEmQov2i6ji/36lPuVgXmfIKBKQ+4qAyz/irkv+8Le0LLB5Xvy
PVgJkKtOkFK1ds4AFzRRjZ9CCCYCEgKbVsgr3rXcKuYtC9HuAHjZrUHfeFz4
0Dh8x93nUQmo9aqSvbXg470cXIPTIpHd/K4G3jzGU64BCeMWTNW1mTNIHI9N
HmKCSe0ktQw6xZV3R4y1YFaU3rHTSYr2PudYzamCHp9B5xPzw0pnoqSQQxNn
QVh7rNO8su7QRpZcO/adKy72EfQ6WlbDE6XdwJgeg/le/gUfXD4Ojb4fZ9Or
+fZH0U1yUgGtbhODVtrj3E+6L/O3QXvuPWLik04pnisVJ3ihHFHZhVo6tJW0
XzPOVOMGZk5ZVZZnNGlk8Tao9BiddYjkfUNoLOJS8p8ly3xorEJyCmKAR1dj
mZ4wND6FgZkaseWhYiEFTo9Z7uFgXjpJeOK/C2ChZbEqCHsk7celCnsi1zdx
WAEpfsVf148T8YZZJZZ65CUk5uzK58zKkMSEhNtu7BB6+r8OPlvhiChLboTc
Dfj2pAf8L3JR74VVD0enbDRZgQjwByBsRV8ozqZcbeZ7BddXOrV2D3pkuquq
mDuCruDXOAyYC9PvS61uC/BzB7w6DcphmEm843o7QzUZCtTmHWHl0w7xnPwV
z5IvTXk8nxZVzKIi+bot1JdlVZPsSOGcbkQvJIxWtxZH8j8DOiHggK3oSBHO
BbG3SbHHDe9Ye4ESsCBUnN8nQRV4D5WAyoOtYt9xkuZDM9Ib6DgeWnv6ZhEg
Bwa0mSpdfNDMwfLeuRxjCLkXVWVyAtpjbpVDKNUHYXMM/rWotlmbM86KnRHn
lu5jXM9Tup/3TChNCVipDfTb/U+91PYwPsG2b4DRcVO1MemULq6+bNa/XB47
tBu7Sqm2I6XlUsxf6JHc5zAzJz7OYWycjGtfYvAUoc2vqVdJ/qvXHRBKzgyO
wuEmN00A6scNkEnEwsOpVANQpbuURh2mES9+Av6sVXMwri8fZFuHmpEYobzD
XMZC3ZCFZVr24O3hyisAnzMWW8W7UHL6QyRTPGIf64vULx12RC/fqw9IRw3Y
BwdXQ+gUvg0Ozgecp+Zy8T+oDjTEbGBOqPiSJaGrQkIQtE5gvgjnHFjxP5hc
Nf/uxjwFYye6oEjRz3H1s69f16yo3eY+7dBppzLEpmPCLPBrKKkKW+ThzcCY
jmy7PPD492ByeSdAQTUkwnC0RYwlyeJ1bqT3VH5XxxVEmv1YufjVEW/Vr/wj
I0TfVjobp607z7ugGBI2EGv3c5GaRUippf0zg8NaQGjWiHFpfXNUhB9FFwnt
z0+buIMYiF/tJDKAmJ09eP0TZ9u9n9n6vtDTK87C1OaYxRf3AQdsi1hFN0i8
mz53aDB12mmvuiPwyOJU2YT+vLtMAFd3XV385mvbeu5jQyEvVjDQxGWMdMMe
HUrdym3hyWZXEW0+f3Up6daZEOyweInP3DUeUUl+JtCch4Bvqvh0WBfzgDQX
Q912ZvuOCFPRaYSzz6ARqb10Vcor5IM7OiPOV+x/Mcm6hk7Q8rNUrH+zUp3p
6zPhQTgJw4kF7oHeI9uD7ajafPMiy26w/NslfmRV+SmWVWcKoEgZKJywoEQE
BJW8YMOUDAHRYAZMfWl9uf2OgCqB6Sz05n6k1B3Zo0roIr0ubIEb7P4GSBnG
HVB+IxAnd4+czDbg33M6r5ApkHeM7b0+VA/g16HwEHhIGcOpjm7SNwc1T5aP
K9kz1XnYX1LN9DYHzzL/NodVbK80pC0n8BgShYDbCY4Q8QV9TiQr8DANosen
0OdcRXrpct0kISs1ymHkVXuvyWkMPzIURjGgP2zy882ESGgPaqmFNDfEvDR2
uFYbDgcjCK/X7NqyWVyqxx2QDGMk1MqyGdimCGnNr9LMJgd5H0DK+ZZEepLA
VnnJRykdN816IInhgZbaAwiH2l7pWTiqiPHAsWxdDRKvHhThxQY3QiXMOQX1
NzUpIN2nrRBbaUPiyRTp6uoU6uQ1GdlOO7V/HF9yCW9AWjxzHap6IG5t9KdY
HwgFcsr5MEefoGzK/kFmRiZlP4+jDyDOFgUpxjVP0p3RMmTcYEPIRE9hvzZR
+Bi5MMvjjJKQgDehA2Mdxt/q7DqD3LxbYLErKugg/q3U0ZPtBKt5faE/FZJE
wJ/vY35ddq9+tDa00lK3+dDOat9z9oQ9QV5EyFzb734g2F+5mfdTcoCxI+/6
4xj5QJPdZ6XM6KZjbVgHWeNDJAN+YF2cKAam9xinfopwSqGggn70GHraSrNw
fw3xfWrBamLZTLFIpoBovLGNPrfy6CJYQ/eYYaOuzLszlb9wIqbEZRRG13Pq
d4deULjVDdJZlSgzxc1Q2RExk/iiNmocmsAxUcasWy16aW3TLjXjuKCK517M
PwonNs8ELGc4/JNEfwgO2KZ00vZBzB3EqaEKFxf9OtOkYqIU/nqa2S86qe6d
CxxE74+By9R9Yx4wYleEkHbwq0vQhl7vt/950Ctfq5M0YuqXUCXrUUhW5lbi
6jtmHSDX1iKydFbvVD0EmW0vBxxFEul6ezas+5lxsxe/1XocN9Ahkx4LqR2l
p9qqrWKrtlq/b9fn5TBIY9CaIHWBJOYlyZbnXd0lt/crnQj9Yo4IEab/lTKh
yg3cF0KhlinWWfR/3syyoxfZwN5J0UBO4pyOo08164FbrtILXDhTx+yrrJKp
wy9CtOoXu2LQKYgPhZanIICjIfIubk/HVv91DWvUVwzXWyC0U1DlhljlMc+h
pRcjt6zSy6UjDJvE69c43n793ojygZAcFbpugty6lmYMJzrfm20/GWRYeCUo
ABy8fJeLrEPm398vVFKRotYDo5N8Jt8ZcySCp2vxpzFh15fZ9EvTGwjIr7TV
9BdFvRf2V5tZsJiskb2qCV+Yp2yk6KaAyOCcFzlxHJn7SCUJwmxAfuF6eB8w
KWJS15J9yrRbRiRPZiYyRSgNY2a+gCoCw0TSfPWWsTroaUQWCZCjAMkkJP9c
09oEm8QrKyTE+WwC1AHuSV8UwQkDjLjcpnkIWhPHwKJOeB/+EIilQhMVUNVw
zLk5rlHZJACT7BnZ6QbwiIkq86MCb74eatwxiRp2+IShJA64eLooBD4Pkge3
3evTEloskQJej//yULM8LVA3QSvEattdk3KCEF5lXMQhvHz/3B6MkX6rovce
FFkZlvMUzL1+Xt5DAWs07YQ+zlOmcMHSYKkcZ9DtyLRj2x53X9EGhjFQAcEB
/5csd8AvU0tbiAgGybaIJVoPZ32C3rK1XXaJFAJIY1nXljlC7qT0siBF+qLR
lzeUpHOOEzZbiCDuLZerQxajU7UIqPYDrx00pdmDGT2Vn7fQ5Nn0HzlQF+Ly
nuipAf3YBH7ms8aueRzo7dXrSZU9WEcQt7BkS1+nwqLZz4aa7myxwTQSiP0+
+4CJEVNn1v6ZpOH85c2GnU7m91QK4p0/gbumULeISpAoRYth2RDFRG5vnzyk
T8vPQJN4dULSk2s4YhG86+7G5qQNlgyHoVFUEd8ATpLqGjx5T18A3gFLpDeH
ASmUXBxrw49SKZTMS/tbpDXrQFpqjCXmp+iNr+RMBr+q9Oq9Wkcb6KoshEqW
sUriX4NGJg1oHTlJinB0kSXTSzmtVZcE2UPw838u3G0Q293nH1IGeYC3LT7u
UooGk2pPdQ8r37kcO8owW+OnphmDoDdElv//anDKs7Fn/Q3H+/3M9TO2Ss1f
nv/R8D+jGGxXB3yKA8zO4VTu2u92EJSXcUO7p+6s7D813VkZj59C6sMgJJSZ
IBG0NcBRnKb3xVPdSFR0tnrBGCeVYlI4sgnQ7qUdqvwmIfLxMAwFHZbQW9Pl
n/t5WSLqA6nqYuFmYGRae0z8unCDIiaSrDBcJ/DqsRhaIp19uvf4KXY78Yqx
cwTIzghmIKU4NzQcDSGF7u8hGNzyv7PA34Y5vpefqN2w6X+T3PozpibKDlwv
ftA4/IrHwfl8y556cmXw065TueDLiTzrDd1zhnBBNH6jVQ38mvERGNHTvp22
J2hxX3InEcweQzp3+0EIOgnHgk+EU1X8i9zxn8rHUyLESQBHsT2Dw8itDWrv
fJ2KPXupUDWYVZFACawq/kjno8g0/J/eVg9jGIDE7nqVN6Bjl/EZYkC/a3SM
UeaB5ofLS+IhsliVECbHo68E0xex3MX0tcm6hGe3V5UAexa3wQRnHX8N1IdK
DkpBbEAhV7RdecKqvgS5DPTtgEnxI2hN99mhIyOnYeQ9sGoUwbEflfU6In1G
XPm9AZZeeQ9BxreCkD0aomH6gLesfT+sQMitPL8wcN1wpP3t82b69DLCC/m/
dmABCXySJplHL//kBb/z3l+IVRz61byjPvf9j2DXe0RhzBiffWyAu6MqvXCb
tsHsZejmHqhldjNxxYBRh/jVcD9T8vAls6ZdtcYNqrVBwZX8mHDR7SmZfqKD
U6euyEzBDQVte65Tn/dVpgELBJ8825hDmnoixvsP72B47rS9JSojcqDSMYtG
7teMWUDVKgm0f2izYUaUdi1edXwTPlRlu5sTIS20EBLLlQfLsMO1qVeYgP56
gk5f0KIrHA1vT5aT3w0X07NFzdCoZaGywy3owhZA91V6Fmof+arxTb7S5G2Y
BLZ3X5vU6Vhws40ha75JC7oVyN7SeUuSuPqS19H2sSGDbcByEwN58uAy1nmw
BwwgElYBGTEmpXXgTjFJ+XTYODpy2KiFU6jiwkR/GqbIdOauI4R95B6v4XDT
ywshYuZD7VEjmkEwWeHfzSX2Ze7dlhNFiLKrSyuWr11r4NNv6RvKOYQOTI3C
xTA7LD62G/8jyfE/jlBfDS1rxV8+m3R2EfzdiknmQrg6k5UBAFNq1sxCwJmc
Ky5X8cAB4K/uBFfIzjceOCJReCYtedVQ1k3991it+FHN+iBz8HqyWQ3plUlz
z/K2F2xsWpts6+IN2MGOQbhwGI30XnWwNUDJSBSk/3q2x/h3scKUdwro7PZP
MwhOlSbkUIk7vZCqxaoayNwsmMARXXKYPm6BB8TDfwwoO8MVeN3ZEUmsrDys
dMJgGHZsRppEe+9EJ3c1zir+fZkGrOon1joCknb0J5dHaPYF4P7GQa5T5nVN
gsdWn2paRdF1iQhsTsMLWfKekykyhBkV2Oy+1ATEEIoRZ/67TjtkE4KUKHqf
8qKVAH1Eam4YQ5fsMQ04Vq+0+7ZSDN6iWiVBpNLdX07HHJwLAPJxKBb9wHUS
637vCBZFmhM11710LpqLBRidcBloAhHMApzO8KNTCo/Gpqng2Fg83/jzsR5j
z/iOlJTWqVb7UGuvccRxZ1Rp0F639/oBlW/468lvasYaItk4SNnXHXZkYQ00
e+8TFGp0EDqfA363/mz6g9kRAUMFOQDyK1AxdSKYY/UKqvKiqIQ4Ur13NZ6g
ly/ypc6OrWX4UPZvcJOA3Ulwq86++61ewQdw3K9xmDncZi2F26YIHrgqMH5A
zKfnFFF8bJmqffPwoel+LpxST51udfkZWLwGntlpc7U+OTF7xfJsqUeQ3oUN
ptE29IfUe9b2vodA4eVYv8qrJnkki2j1Y78RdTWuLD1SHKiHI8ZfiC9bZGOY
5rkRmNZ98LvmWwuVX3QvZNff4O4qWRMIA4JUhjogMsQ07w1q4wE6BBuMqeZp
uZk0wO/6Xma6XsORV0JHEmwQAhFYshwmW68uO/mQe/mmS/a8YfssRZf70Cin
drUEphjaJiDbu9TTcmEmWi/F+U+zKDHwFcS3XQzoPHEtf/87SYXV1PWjSZjI
n0IIrE0anlkhYpA5VN+awtlT0++0FP9oGopGBIEbp0XljQcFTpPyHGOofObH
qB4k4f4VcLOxhzFmEiOm+9eKTCi+S7s7plJ2AWjXZM9B6HHPsNS8fMSoRBj5
JC8xcOHaCUhyUZtCqjucJ00aWAPH1vmf6njzvDKs0OHQzMzvyJFIIeVn36Ik
o+3IbKywiwRx2UiiRXB0VzbZktMbAS7q+xUbQcf+CaX90hpd8FwnzvRI2W8j
+8BRfBciOixryqkwESY3a5e034ODGTkKROgvGm54T6KuApRpxe8XP5AXGKwR
I6jkbETCPKYCKg1kYDsKXuFJBxa0HVd6IGAm3nSZn8djkAU+xc5RVt+nk+Lq
CHLvLn/JbT7xyR1n9YE4xVu76j6zeH36rbQpJoO0WT5dVufFoUH+qaRNfMyD
HqUJBaBDJ8Z2dOkRjCWQrlUlgrMYGSKkhKr0fiFJXLeMCnGhOHt31f02pbui
SyAUBuJEEJoslYxyo7+0/apjE0YS7o7nAoflOawAG4TaaA+4MTv8wFre1wEg
EEwKvLr3y+2i46EqeA+Is9axuO8UWprcACTEOxm43ZHJDerbrn62Y/33kKl7
TavH0GEaFLZYdTB0PSizTbJwObTlOwalxSFD57DgdhcYGwqFZo2w/NLKrody
MJKdNkcBJzgvqVq3V745X4dj0DO8zySAz3Q0tK8MTckCF3jbo/MWFMPqoRod
ZiGv8fThCkvKznTz23GGLCKH/DiyLV+aRAX1wlEd4Cih2Gm3cV4o1nhWLg3A
nA7gNuXm8F1KVRpm17C97vLuq5r9EjR4o2tyr87ed+vQld3I4uY4UseNfNXm
6IoaZMNyTboA5LYl95D2BAAGJxZo09HdCQuHpzGuzgptnnDOMBbPnICPT29n
NjrVpZz35ycw+TdXavyNu0FQAD1yUvAv1/p9S1b7m71hdrxZw7YRMdsV/oGe
9Uz6QMvgOVbl2GpALyRFlFU5eAzuhasEPN69QrvecHcTvrb6H1xkBeQHXZby
3BCOj8ac18QhB+m//OBzAXkJj5TA+BvYm1VVDto7tCMV+4Y5qkTuo0IG6S9v
h4KltxofEgMGkYpsBekcDPe5ufQnmLDi/2nPXg4OCNYlaRCtVgc77SyN9apB
CqujCMZr5cjY0J4CGxOJs45Y5b6h+NizfqNxcyMLeLdDpa5YtB1KI+d8CcVp
eOremz54/qZliwdHakuEvF6WZQ4vkUW2tK2J841i2wA1G2vTMinwFonycHkE
ZkHnCxWmNhkA2hzmI7LogYTGR6oGEd9XaBxZbTqOqnpHV8udipaMUY6RxkeM
rKYHctH9ykD1D1OPKTU3vWGO3ZoCc0VYc9dStJD7LTyv4X4K+K4xyH1Yvx8r
1/5gfPurlV48JJukeSBBUvm7MGeMdNnMFRISZuZGcsljWjL1T+I3xfV7AsYU
Tr+3uk99cxRxDGP1vKbvoz53UowVpkgX/ieNxXmrqK5Ay3t3SiK3fP+qpemE
EkI6w+XLrgwxMMtKbeubOuXsdPTEakgTp7stow7BRJBCDQynFH9h24TWXKNi
y6qb0B5JI9xcip1WdMmibB02LbXQPVhMsiY8jDt36OasKtVw7LaweMVoEjZv
xjBRg7LXek0WztqSukcLxxA2vH27W6LjOU1E18/cdappPZoCxb8uBEeOiHKS
WDrtywWJYwEcuSk9EyYkpgR3j1SIx8kz/LYDUr8si6Qair7CUPEoT6sDQm+f
TC60Ctb7jTl2GaWwklKDDHHtFW4h1s7TOA9GP85GNScr6WArSPgd4CQX+yKR
N+L+Ly1JfKuJ4wMI6AS2kibjHi7+WlSlXqvYf06BKVRQmnnjyOUVjVO0NyE+
nZTnugDEk081hdYTxR6sVvX6Bgri9VeK6G98SxVdJpQ/CGXzLU0NneRz2XGf
aVpDV+9FxluSuDu+Z9vzWMvn+Mgz/OI6Lsro7nch2uzpn32rGNgewrpIepUx
nl++GlJvOXHZl2pO9vmH07j1T2DjxRB9OUrm21veSi4cnZi85rxHdC1hj188
uectmPdw+cBIrOBkGSjYq1hJLmu/BXsEFBS7qzBXSBydz2dMJaxGcUJFHgGR
QPtG/FYaRRs077r/32gIMtpnOoAAbkhffOUT62Xi17HY242J3as20OyKsgym
VWCUi8q8r1bf0mGHvWz96uXsZZzW1cydtv1CB5mCUaMhTqdM07wJUrOx/wH+
7qloGkR5PusUfWym5uA1juAbAZJbb4LcUssfzYLYLOMZ3mqhOOkaKRXj9I10
fBvm1v2AG9vB1tvQRFVuOSpLoOeTmLPO5FZ5V38/Rw8PecD21c+hGx3bEf34
zgt/+jFxUdkleRo+oaRWLiKE0IxagNxPXwx43emp59erkerdCeA0TEYrY/Qc
/CdzIlKoFNj3Sq2aiJjS/R9wrXLhpHm6BSiykPP3ouBZ0a6+pTeU5na963xQ
Lq6N/q9qu5ckhJke4Efkg2LSYCg7l6vt4GbMlVv/v65opyux8fBWp8dlTGMh
E7yUDGbzRXgbJQDfSERNJiLHFy90kct/N1mbo7o3AohDoppCkWmOzXK6s/2Y
IeQb+idomwkak2eVVlduoB7bBWZD3+GNmAXLsjFCPiUiJSn4cI6YFcHLlnWq
V6q7W/QgqwXY/pEFxGUjzZBBmXGe1iyBWHk09QGpUmkknZgC38aIi7gqNdTW
KjkvyBbWVNPDfht02hsmJrbhl6K1KkVdAHbNYbiUHRmd8mV8kiwcUhjKC4fv
EKg3rwzS1Mev3tDJcDFfcwtc9O5PQwFBgkCZ7LvOPzA2g5uh15/nNojJmWpg
e10bv2y9ca1VUXiy24FRs5hs98BKrQV1xd8bHR7p0BvN2ZVhqWhe0e96ig6h
zkSCbmlCHrEQ/IaITVBYq4SuCU0XwjsYCraosGMEX6Tc/0uBRMpwgrcQqlOO
2paBxgepUwca2DLC/xFr+SSkoWXhedEqpdie7kLK7BRbk2WlxUXq5YnRiAkD
+hYAI1AWHsDlgkeGzOMH0BwtZHOWNGRWoAXw4UF8cUiLWjdSdRKRTEEAGOou
6FqSeLsLNfgJzqHPMm5pSN+qJmRqzgNxIZnwGcA43z8a9mG5eVEMMkxqglM4
ybRzr/PseFa1/zUOX1Hxt5OuZlMfokSvLpSR8bVvMnH7O4LW3db1cppAntGL
wtBVXmofh3vqpdAbd03PEV4qL7nCLgHSJ2fKAfrYD+T/x2SezLhEphrFhxB1
Ww0UCllKuPPLlLZgwoCxJkY+TAmAdmPMFt0jkK8jd0cQ8tRtYSvAkAKDNfyr
ouPUgjbaYeWuqaqXSuzEnSK3NULSQlkP79uk+8+oKizv25lA0KJ+FBh8vaYC
YsQZ1uQcAqwz3IElPk7pMo2VNrto+NKm74qCJy9NR2AJtMwk6WVYpZ4qlxZF
GEEhQTNRpqVWtAegL9e1XY1qh+GGvsZ1pIVRSA8b8goZ3vuSh6vd/3A+N7Y4
/9nj+PFXjfWdIDxwvWcsrL2MXNCN+YoAXxMFGrBwlY++R1rkOShxHrH820tG
/kaCVKV9m6MsHOZsdJ0akTOoQXSRsA3LDCbQSm+mXfCYyp9FAmzYvyvFcHNT
GqC8EJzUORC50Lz0zQJ89oIQjmahnoPZrBb1FtY0swHi66sByDr2V7nW/SL0
8fliACU0bfMF0FrFo1RiGkdilSjd7Vmh4DQXDCNyCbfdOw/SQjjxmgJS+xze
i6ijzu9tsmqlAXTvbf3M9USMG9hS6Jb+owskwvBZtcnS7lWkVFe7xj3M2B32
SXbVTKVryjmiqmXp+m5aOVaBh+obfvjK2eumj5PDucM/dMpmvseDRWj5XgwW
b0futtsuVZxQWx1oZQqBdkHzKokX+n2gsXNFK45aqTnFh9s8z9P0i/UOkpFl
SLmRxTyVCWS7LRIjk4Y5JlhcT25TTl1TRXtuNDvIV3tRCXWGRhxBMXqok10F
i3deJYlw18DOWFSDpp+7yeA2w+Ya9SqaJ708Pa3qa0epvUVqOWzTHwddNGbg
F4alniWtBZ5JEkJBxvbGzLwTK0NdEehL5lBC/SDxGZgQjtZ2QlpQPRqcxxwG
w5Y1Jrs5Ny9vrW+TUMORp2aj7LqVv8Go+KgLCq27Vele16BVjDAIW+65h7b+
gXhG+C2AoAZ38mfGHxOY5TLUOv+jIvW5Q8F/OprWfwmDlK5G7msbcBO3wgFs
8ELcjN5WACUbONL+G3zpGR2p7/MoQoH1j/F259ZKmT7O4PasKPpNqhmJi4Vy
xvjp8FuNdd3G7ghSTiS91ZV1UQqibuqeB/gcdJALaSkEhjEYE9Js52F0rD2B
07D6ZTOLIlmpAgUqHFtQ44A17fd/pCwzxUCzjFWp/JYl13qwlbjWEmYy+Ie8
UnSml9UeXyWfwvp4vq3tuDikh9Qh1wWWZLfhL83DLRrJPUQJHMOvUCUgs3Kn
jaT334+pwoErvQGHYk9fB5abOI7INO6jCGQknbdCbahJRMfMz2lXHWUF1dad
SQPJLU0dvNPZpWRh/NxXeP52nW0lHeWdBiCM8akgbvvqaUXI1e0EcxTQ/4Kp
jhr1VnlqW0mwa4Vap/uD9IyLFuiwi77LT6TLSSO0m3lGPh/+ZAYsjaR3z33x
A3jALLoGLYogx1NxbhWfZxEsoYYwDKlg/NZAQ0/nEvl9FEAMc0HUu6JjYilU
Kj0oVtcIYlbj+niMXPKvJhj3/gdNIZNmp6aDq9zPYzPeEU/gMGRwGUr31Sea
5rWp6ya2jys8Sj9JFFkPanKbLylIAdtiaA5K+uGNTFDLXha86waG+ABCiqW1
qy76p1DeO+H+v4+1ZzwV0MO5lO43m4y0b+N1olrQ5M+rgxhT8fYWllJZV5gJ
7jNtX/InLSL7NfYshx8GrsGLeNxR1rVL3xz8Oc2O6/U56woGnzlURAguI9XL
xAZ8TR10vosKYBesEXMdYBLvFW7OXS5jamfy4LeCP/7XSk8kSiOkaG7NDlIo
EyQTAOFeX95oL7taScZWAnEmekQH/OMbNykgVRRNzRv0rbeybS2Nhxt9WdLe
UYHsKPjMSVeRNF5Mxnychn+GnfkDi40N9OC/SYSrPy+9luah9ZtMcUYaJMkO
4u7w0E2UourEQqtU1bMmtZ9jVWjsz2OuE/4eB7Z6NSpftIVpizS0v5F2+ugW
kMztK+0Hos/HG4EeRvdpsYN8e8voilqeQOwxj/mOxCbjcSGAr652SEe0ZFy3
hGMg1jMZb86fie3ZbmE+DNAe8aEX7E8+bn6eBBerI4+8FTDmedXyEFCYNOn6
eo92F6MM2E50SbDnmlrtf1QYPf+ahZHMR0TrJ+GLWfGA8bm3s3Z9abwaZb2m
bsYcIlOewRj2djc9yUikyJ37oCMe+OOzQv4ajlCURpBKTUqYTWI6TA64s5YG
qHnoSaufyfmSnbD2NRqKZNV123r0npPbGFXO+KZZLUyBmKvqVYW3AGSfMg3R
ak8hsyrVzC3951ODn0iXIT/svWZTz1vrV7Z4y5fL8DSXb7gztNTzXlYVj68S
KISCl4pcw5XgRz1rkMgFboX6g+OzRWp3uQzq9RHPUw77GuoxH81AG8W+wZuO
znYQPtrsVYfUIQyT8rOW8RLIBYBOSZGrlVNxh5fB982WGp22CghW4eFWxSZF
sVvB1a+qzU0wWI9hz3pA/dDcIyUKbY3xEkaKHB1x88ceHaBPu0PyH9XUp0Ia
1IOzA2oRjiQ8v2qufH1V0mGQcJigVn5+RPY4colLJRACA7lMM66r81oOEQ0L
1oLEjNPIbNIfrGjvJoQSirZgj3z6NcQNHfVZ/lmmE/75PirUMZJzWLgnOaAv
2bGt7JMQCw5i+BRGABitMwsZ0jseGH8//YYGqw79lIBut9C3PJsevIuvKEwY
bFxwXFD6Y9xek0pdOvo6iYEYX6ubx/IBehTrQZp3JC1luqzOxjo3MrjnzdUL
5G07EhNNJQd1k5Y5+GQEFXthnUU2QIBFnqL9WEkMTDkrkZLK8z18Mzx2l3h2
k3wr0E3MAH2iREUlhkwYSwnYNqDkGw7MtdAgbammlDoZBm62kS4lg46jNC+c
DNOjE+OF3bNL+OxF75Sv8OFPGqlJpbE3CVIGj/6S8eJfjKcbrE2FgJLyu4yR
vFF8kvHBb6gMtMdsuNLKPKCNAgdfGUPFVf6qcYjQZjgEKiHDoA9DXOzW19Or
/dVM5u+yFB1jRQesFwnOmfAsONa24yd+54o47mcmaU1scHlclq1I6MQcmW+S
eFBTnoFoB+C6KJxZe0xxghUmbLRb6gkr1oGx4b2eaKcpe700jWZ5hKvZsGby
vUsqvjNvA0F+jF3hhEsJJjtL9Db6ktSUmIv9D/Dy47QEGznUrG8hOnK/E7B2
e52JS7PR6C6cWlNm/DO/yilmsAasrLBYy81VnxbOQ7kC0M1RSMbsMPHioPzL
IB6ATtiFTkuUQXqRWIAZi6q8u2cA5a+p36I7+RU1HekMbl4fOfdl5gc4trSh
G6odyY3zhR62XustGiDGV7ZtFXhKIcCdoMbKc32iLznvfFlW/GNj6QaakJTj
ySMoCorRGtA28h8vD4G2cnt0an2bsZLcwK7bgEZKrgf4nZlpVLRk0OIN40zi
hEk1JEtvdGCmI2O6T3RH7pZCp/Vntl2R3K9m9pJF6Wrfx2TUApxIFA1EZ8g6
wlu9IFnTMGNefhguDboPWmd7KIuEPJMhQZ1Wy4kILzMhglvbq1Li6fm6LsdG
Y8wfM6G/YKUQ/CVApiPOuVpicFhhM7qpHa31stbF4AIRj+phKK+Lot3XSI2g
RiPuDzT6j+KcBLh3ldMiK0HgG0Efo/qqRb7tEkdp5F17wcXJxDmyHAE9rKvo
layqxum28Xeg2ILIrLcZ8LLvuoToFHwc6QIeNMfe7gc0U3vzOfVIt8CtUVkT
6WXX4ja/GfrL68agj66cDg5OLFkwet9nnYHx/RUed948c6kiiJMaSuUvs4v+
Rn+gzA7q2H1S2ig6SxEYnmGUOr5XNkLvU7iPVUq3gVgUp51kyQ0CnFW4sitn
SEc1oEtls0wmny6HVU1d96Oe7PZbrsOa1iPG4Xb/m57LzaO8s/t6LLsO5bp2
NtaxpmsFENN1VYpTQ+7Cbr85AoqhllGTVxJHZ7dYdiwGDXAj3U9l7KILH5vz
PdxCWimcYjhcy7JMZLrQdRI4w+KjA5EONREpaqbwxk2c9bdRxBxr2JS/h7Ab
75xs59WAFwwYTZM+zJV/gkBrvKtjVo+ZB+v80pQWtx/75B53Hi22XJBg2Xtu
2GRH3MTAP3xO7lBeHc5WJ4fdP2EBcgWUwGDVR5lcHkp4Ff/5OVFzdKhru3Xs
1FmKWDy93as2LA/8vp2aWtVRK6N7moZOQ/KEdkY4yDFeJMG6v4fp3vNh712K
Vy+3CxIPVgi546DL/3/AgPiCML9GXl8u77pkjViEm87Pk1LDbE73ofubudu7
T0xGCVozSxfEl6M6NsHjsL8iErX8igITDAj0drIVmBVb1n+vqE/ufTPv6FiM
fn1lR+S0gps7yQs8lHg73LCLcWb1aUg0GwBdL0coFHpA1AkN/u+UhcgwXX2l
JoZIJHmkUS8FNJ978cYRc//V4VdYWozE4RI3yIfxtEqjsGLs5I3wwFfk7ZI8
gs+Pf4GqULQNCAv+btexHXrdHR1c/cdjGyl2j/bG08cgxIPRnUhh7QvtWrrj
PIz0M3OuS3WpvpCkI1AjJOKuVOAVfiYArBDLNdEvG5Vo8rXx/yjqDCJosfAa
q9M3d3Azr0CrVwpdx3Z6K7Fv5zPkZho59IN1v9UsIqbCLIlxp4AI036ccrFK
y5zOBCcGYbxpTEnLpM7UZ/EnZRUhIBCj0xtUERzXyKRat18avTBRDUx1iNDJ
aFavr/YhKTr0efY/WERSgeQA86zZ5C0i1eV0Ht+RACQ4cJlP5Nx6x69Umajc
FltVk5JItMesLLCmnKDHeq+tjC9WZfCtV9Y4pEvJyvEPLRD8NBlnIGoTsav4
b6S+pFZqjeBgWoxSw1K1VPWKQd8jmPzwamIQEDT2CZPtZC+I9iHs+Zdco51W
ZONyDQE3qfu9xG7yb3dl/rrbgWGdSPZ9ohKvegVmy7XnCAcUGEQgFSIgmhUz
8P2I2QD+wlLKN8jdIXIBLhY4iiqtJdm7vdOPjwr5Hxk8lsuTWMjmNFLYkqWz
bqhw3qtX/aHXIjuz+REIg9Qzeai77juB4dPmwYVM5zJHPaOE978TAzkEv/QA
bnxCPmF9qoQUTnbvhRKoFG2KC49kNYQuBT2pTRqfartCE5vE+TnnYL9TOYIm
YKE1d8WQvv0pjc2cgvqNDM51Bm/26iRFzBiZoIj4vgPFhMLSTkoW10Fz/Z6v
B7nGuOjRbGEiHut4cak234PJxLQSIHINooFwTql50ZetQc6sCIJWssc3cJn5
yuvRS9Amg9ZdIK+jKQQnu00ZVPlBLBkRLiKO38Pp8DXlKbltumRCpvrcMfWA
Ir/PhshoEl0vpuaKY2fd6fnJWx8NqX+tUEtd8jURg0+UVVKa7IQsJialy379
jjIM9TG8fg9cyRLH5JqkQyna7nbvxHP3Ce2q5dPwl01gfebdAuO7XD7DjgGh
OJeHhJWVNwvkX7fXaRxCWnagAPDvvvyH9c7OrNTspWSXMces0VpHAD3mK5Iz
aNZ2gnksNof9IJ2AQDynYfcAMw7lgOEBRws8MeiojdSbz07+eTqA6gYetMKU
+XOsQ9efeABdJreYpPOOMO8iPqCEMd1CsvgQ15yhFxdg0Si8e9MiMfBrhFkm
4pHydTzL0U+AdWkpmfcagNnh247qVlhTU5LF+WZWDFkA7e7WhzIy/F6GFqho
pAqNDSJQby/scU0mF6vrtSmOn9p3E+xfDKcxwwq8Gx1gi4xPc9gGiglsgnte
a1/C1OzO2glBHmR8vliCIG4Ad2Lccbr8KQyGZPCa8v7kh9R0vaAkUNDBSJMj
Tb1ygB8xMUfFJDVgA+z152J43tkSgEGljAOXCR3aBigt3pnK5/uhixqcanA+
SwXCeg+s2YEBbTBAfqKqF/bAdF+av4nylo4ZwOVJj9YPX0+b5EAiBtaLW/37
LF5Mh6KCh2P3poT5mFL2a8d6wJWSFelqLc4eiW1jV6+vwtWqhlL9IeoQzeje
kwukyChfXjqnsbg9h5pbA6aKG3baQVX5atni7z4FluHMgidT0K16/RW9YSHd
MH0Hxha4cCtdl68la//I/kxjJwXggC6zecYp/eOGMpnFdtMci5/j9Ym4fygr
4TDDqrCgzHQZpXsVGSH1B69M/pyZzwD1BsNCqyd0c7b5xpnQqpOcAyGWsJ6R
VMiohFBTmI+fIyiGa6YD3KQtJKN5PrJJr72tWwEyPsUeL7XwabSB29CKp1A+
g5QS5dwxTFPem5droxMg9ubTVVVDTUwQf4ajqmv4YvxPZa4mPLPoBRG2sUPo
5PqcfTDOycUNteDERoYVLaZWR1eNTe6EZ60+EjKu5GSmd95msx2CaOz9Nd0F
lRmqAfLcpNBqLHPtPuEYrGTu4OL+UNXrWQ/9Bc2rWPq+52o82XvCP7sWEfQO
zQ178ZY3sDI2UYAhefi2xw+7USDm1sWoWZF2Jr4xYAeMyqOiaMiyXW+/mLIm
Enkrp8HL1qHQXkgN5iA2FdbWyDkj3dAjom+iA+V1rKOR7G0QvucT5DsFUiEb
Vt1Mou6wVU3N7I9DixJTTTJiTMvagGGznDnXPW6vPK07q+vQatkgnV5pqb1q
KFCN57PHR1v1YUhTjBJWe+HHYyugvIhwxWWIE2N7bbM/mzb0XLNtdZu0OBE0
kV0JgIlDlqccA5DSpO91aWf/mDnovji+h/mBFYdOK3XPSwvyALOu5rmjnBrs
Qh2BngGwj+FsqwCU7VH5llavJUgBA7o3XsRUHYHo4foBInD4GTfo06Ya66LH
aIt4G0S+WunuXO/7s/I9/PuJSOkSIfeILklsMAhzMNaSKXoIDWUDUsoWPge+
zpuyKuUsfR0eU8ICR79pYQMmnv844IIQgjBEPe1cmpYeiURzqQSdr4tP7nIA
meRWc9gnlWt+bcGspbb8/a5K2VDkWnDySe45bSemkvJe3TjpIgt0QEw3v7dx
6RhLi9omO4ZDay4cO8UXEctaHQMOWjqkmyNthitHjE6picqjl/xzdeTqp7Ug
m3lHVXfP4MuaxVASKXluqArj1hzLEBRU/k59F1H7Ltl0OS+Ohw5Hkm2pdg0i
Gb9XcSByj0bwQQdODKQ1x6OTWwdcE8NrZ9ERjOZ8AMGi9ipXGGZEUu3LDYac
I9v9tjf9otQ7V9xezCcnSlGPeJlL0p8+6qQNbOrKsuMBN7FkkhIblkdziJ+t
ByhiLKBDZIOF5W7w8odLMxFT6+wg06x0GpU1XoweOgl/59+rc7uBljhIkIwb
BKhmNHbsm/oqBQkOo2YFQWNFr5Cg89uoiZX7342cOSDqllZNstNnnk6Sznfg
Q9j4phh9/SeDXhWInw/d9R2pZNKvUGSGpwdEm3YRrtfBaM8PHvr3hnJ6KNhl
HSMqMbs+Sf7o/8QdNEW5E37nb8rNDHcvshQl2yk/+jS/NZA3WVUWZQfcfl9r
+9/GMn0tFKZmsS69YIHuejdbgNgTHOYtCgftyM8dCaPJbvvL6BmDoSa7enHd
9XCgjEgoiGob9jk2t8o7YXd6vmNrBpfyW35TAiTS9Xq4ctyply9DhnUsFreW
tkaw2iJd9I+r7aYb5zwu9IrmQP3HsRMlObnCbEZqxWPmrHBXIuVUGpkjY7zl
GUbRfbYx5gPtTTVgQafW7O3LPoIdDqh+C20lzRDwBejH31Bbt9/ks132eOuu
Sn3bndKt8L44XXgdWdoFbeUjHHAEnwqtm+lts7Aa33v/ULBX15LS4CrkCJb1
HZFtSmmAq9FJMVkK5gnUZH5ZnqIQT3Y9PKH0RhQWZXZ6sIItMjYiND6veuLO
IasYsQExQiLotKHYZ0lGBfdWUtYFQ/Lw01mujLzbwMWrRV26+LbGJAuON7Zd
4JwhdsA4LZnL0GwWoSLWLFZ7jmWCesg/MdcY6KFpkZgV/tSeDV7I0oKrr5dE
VtU1PEikZcwOMc9egDyeObxpmsX4z4MXlvqvh6kgm1wGGcIPHeQ/trPO9Jg5
NcFb89mG//uS4iZeS6A/o2rajEhLZIpbZ49X2e0kFJg1d1i+X9Kx7mO/wfmb
NWBP7EvQt7jyN7o8thUM7W+RFpr0Pa3675MOx5cW+UrrGFeKpmBvYPmmY1jg
9l8qh29APtE4GzopMSOzAr+zrts552SMLz7+ogdmJGUnt+uXhziS4mslAfOl
PY0dZHb76ZXHh743rtO8fcXdI1Z/eTtwRbeXD/X/JXimCLN00bNsXaDBnkwk
YpFeqImT7PlwS3ygVEXfr3WNr8uJuNJCMKJ5Q955SkWcQeIPWxUVXKI/zB8G
ZbZtWVGDlbNUo/25dlkaFb2zEK8cAEUBAd4kIdBCtTEtXjxdl+B+TRW1709D
8ge3bdir2GGq8+msAoSyJ7r9VVoVzhrXYJBwmosE0dn4qPZYxCCsSwaO4AI3
x6Mx9Q1UIGTcy8+PQp0SkstFwcktS1dZVbeBMIwGULBxbN4eQP1X3aZmSLXs
XWazdX7dMuluduELJkTd4dWJs6O+N+YLnro8n7205dnBuUSB7eFuJepOrWPQ
gK+A86m8MaOGDkYAhFqp0dJ9oLHqVV+mR57/nOWLWBKJjTPWdDZMahgcw6xR
NmG2TNaJ5HYeB7fVcVvq9CXtut46du+rSNJ/NuUSd+tR87iJ8ibTWMn5Npy7
5T5QZzbuJoUsnA8da3Y1C+jTSMFfc4EOu07ZfZvacQ3ATkltf/74Mvy33G/B
qmUMXEAIVpMnp4yptcUBqXYsdeUOGoPJUL2rfrUWmCNqpYjx2+vjmw0x/oux
07clKoQXcj/lE1jZxw+N94R1MNQOjyDwpIYYge9osCorCJyO4jaQOWt4KBD+
XGCtT6Xy5b+aOJYuxz6O33/eSxj1flWf4m5OnKYReaaHbVKteBWYlvHBb6Ox
2qBPPrGXQrH6n/XS2820FryhjcGA3on5zu0rck6ztb0mzeWzdEn3YSeXu928
v70a7h1MMRRZ5h0DewKVLKTTGOJOLc3bjZeJHIVk5nL5aPzWAxbnAGISKLWR
ged5wfuqbQM6dxLG3LvgeqwCrBM/nSzBqm4hUjJ7HCkibL0qa0pAO8wKUnMh
y6oR8pN1Y6toeKnYvbjT2XQYid+yRacJRZp0L6LDBIi3/PSsUC3P3Hce+GD+
BY0vZPxY3CxKG0UkEVhSba01qVdN18mA0oX3T9Yy57AcJBoi/HqDa50icvcm
TBvAIR7hF+psXbgeyCsiZuI9NVyKXoWobucsuMoLOHTjOO+0e6zYztZHvL2r
VNPbur3gUAdaQWr9YP2AhssV+KHyMpPfSKPthS8A/G8+rErDKhgdCaUu2DrM
dsAvBw7J1qPNXAvrS2/ndYmuz0353Vun5XKl00VZWVswJdlsqtMsABfe8BEP
UTk/5KR9cvzdOGOusDgpsnZg/1SjDzD+65Orb5nnj7Aa+goyT09U/JcuREh/
GpULKSSL8TLa/4/UbakGR9jI680GP9nVAwccIpmlwp2HEmPJqHI0dFxZ5afF
1xUeIJGLRS1PaaRo6jE30pGEL0eMJaYkAy4jPSywUcXLTVWCYhaSObgafpIO
J4zbDmDEaA8FZl1o9AgUnh0YyFxa/YxFLs3CuW3K08ctGktwa/0TM8lzmc0g
j8uDc88DZj3MjKLKNPXb/Ys6btGU/ZtxccllQeAvaa2XK6VF6Auu/k+ot0Zb
siGx9yTBdLQy+MrTEtCpYZbPtU+tomrZ7lc7q0L3dY3l2SJrsfEs1JUC8RFy
nGh0P057hgsq5tBXhzZ3TiwH0KQsv8ElAXpJ5MJ/bWTf42fTF6JYUO+7G2dC
pXCSda06Z89vWUUwvne/uIDXfg0Cl+h+giwJt0VhRLzXtNXNODHCAVnpU1Tg
vhuZYExViQib0Bu7oqO2Phi1I2l9Kf+upGjIS1XJ0DaKfvhUa5eejvCzsUeU
IDGo2guPCRMd44py1RU2eJb2irUnj/aEQB86zYFTjN5dWgW4BUqS2nKMYFqn
gplrgbVagJzteO9LOEX9MHbw6BKrswWC6b8XYXCyar3zJ68YuZdmt8whKtza
mzhVI5fTmVZnPkNyLpsLPoMQbciCuqZ/I0k4ORI51bDER206dHI5GG+6qQnR
AZ8ROFertEVXKp0YIbtOeBzb/bqq58wYvYOLIxY8a4+J3ZFay+rCUj7qki7a
FFnLG1CS2NJWe3PxDpnTFWpt0jM7HjCZP7lQ11Oy3ooM8PRSfPktjZyGZZX7
60WQ7atGB8lyAVzglFlkhxnp8bpWMuM86U7RkuY7aDCs5JOFcwmvLBYvXeG3
ZkNV27wJC2h3qFUMCaiqqKcqOCy8y+RrT08GsPGIbMVuOfa+OYJiM97p2a6c
QgrkZBEihdt/CHIjSsD761qnkMfoW7PcLUBVg/md+Z3C7tYuoMOih/pv3sip
mD1D44rXU/+9Vwwm4kiGvW7te++earMTDq6+YrNjR0mRQX7MucNTBcVWqNK7
OlYCCW1/1mz/tWN4rBcPlT8GXg/ii2BeYTA0HRy5jemJSfT039esSEoxXn4D
/5pUSeu/Kd7fVPlweVM6vYhgOMM1pru8fYM/1E0ZpiL9C5qRDdjXtOGV2uG8
4KpK1Aa3J109Vfb7AbiU4kTjEUlWFTZSLfYoC73OwGdTD/fibVCFKeBAFpxR
jqXND5TmdgKG9FmVvHSvh+r4o0PzEXcdgp5/bg7VrmNJAojpDDL9H5eRas24
4OrkY7Pg5D6uyAcqesFdHorHfUtbRlDhAXwKUKA9Nty5njtX4YgV4GJOKMyZ
t9eg72WdbIE1M9ZdZMSgtlkznhIau3USu+33Yde/qhyAbTYHsmEH2kZwJDO2
3nFNQQDjwogOgWOAqNP4PNbbn+8P4nTURXOVO85nIohQMRvZ3jkbQlQR9W4R
1YJfpyN7dUDvUC3fYNeSO38bN9W8gitxikoamldXJJQ2udm/iAENn3kpvQfs
ZaIsdQ8iJ6TfRTPvxIs+011++CPXk9yAarIhvYJbgfLXQ0B14nPdLwtG0OKF
79c/V17a01T1RK3gxRHVbMU/k4SUmsIleqtjKii3WOnSw/4BRIRvDOyj8pM0
WP0db4C3AdOYo6rjEKNE20pft+dsIIIgWA2tEU2WVSS2uEb5GpE6Ov2KfyYE
lF5J6HVywmJ8c6tUo63dAKfQPU8Eg/3y5AXr04rdx0c88Z+AEKmQsnER5eb8
4ek5ve3bwvjXEsv4nrtbF3SfvPawqqeb2p8a1sivLhkgDAiwSNQyYVBsIByg
J0OhYxZ0LHGBd7kILOfVqyIAPnChfZsFAP9rRHOtEe6uUHSLPOq0jpiRIonx
+a233TdmlYVAC92Nbq3WCVa7DNWbti3HKiGibJtZUoFn+byPhgWHyjugnbGC
OCCMvJMDg8t6j7Qm/NpVKrrrkPbQiVwIxRJAmQjQbXHS3B+4AM7cgpSNQGpU
lbnpEzoBA7CFMQPf+zPtA+pSDEoKwYnc8VgOC0uLQel5i7jn8+mxpD4Ht91l
Rab6cQlPYXzsxNLmXzqnunL7lU8EQBC0fqcYnFSjaMIYwSWbJcl+qcl8TPgC
9uXq2uofaDCZey1b6TkN2KjJfwE/EpLrODncQHFW7tqRVz5GbPkV/18s+QLI
mle6xDMM49zdzhTTkKbW5X3Lun2vfuqOwkyGPWPbaUfJoPppGpHYvHGFZu5Y
s4oK2OY8HsFAzsupQHYHnPrFXAKAnxPt4McSamUlY9ZDEWRdHzUobUB2tzrA
qxKUdYRIZANNAMK3hCuToaKQZKJknmQ+J7EodGKYmzstqAD3INKuqGQ6FN/J
HEENQRx+9SleBSN/FF/oYmtB9C8gDNm1vFi9aNbrb0Eu+jhyDTgEmiJcCHrz
A+LTc42O2DyuhzJCUeI6IDerepDS8V8dlwSpJhf3N+i6ZcYpsVg9KLeuPT4i
Ym6Q2pXKbXSQlrs9pZKBqOLcAiniVTfjc9z5ua2dT6ZA9RnvZ48xUEaTXuwn
ku1Ypi67d/ISl3ZJsimnVDAOkguhHewAFuGDKxD+fqP2mH4nLKlYWje5P40d
0KRm+f3bCXEdsNSnFc4z6VDA0z2iV7G22/iVqnDRCissjLS2WSKbhl9GjOQA
yBgLOFQhCqHyCpd0kyBuLmUdIRcnLOWBpbXw1ZiVNenbiVG5q05SdDuZr1wT
zyuE1cYDTRXb4GPrC2/tERrw/X1umMUArrBBQHpx2g3LWPPeM+SLEjzJ1uXc
5mW6M/b/8VtIoCAw4PUSCnQmNlZAXjlqzCpvGFGBsXV6vmVcUj8BXzKX1ErS
j1KTf1sqidvWPbjMAsg++4CoTf7hTUdt0hM9ELBddSzU00pjV26TewHLJxiT
zWFxD5EonECLTnIktVtaqCFr9/5x/tZ+VZgDewuc9s0roK7S8vkDGHVYkNbI
iXtDljZKiMMZb9P2UcdJlu/P+DpYmq4BB65PmSwFXasobmHDz2s6UNLxDkhe
xMfpCZABMAqqAWNO4ZuqbxZckoLb99z2uDbzmhpCFw3QWvjETAlSmvGeob9g
G8eehATrgkcSR+HSu5z99TCNz86jKtFVLZ/CDjiC2ZAfFwucKwpBNbX5uhCh
Km9GGz1fFWs7ytWqPmRE73v/FnVDaV8ka7NVtIHUIo/BPRDoSIUSkbH1jZYt
QQpYV5hTHki2bMBKnMIskzR6tZUmxa7NWhFAc5otl+/OkM17f3FDpsTTvi7L
QbQKt9jWsw+Qvz1QAOX+GKpLVeY0O45hOBE5D+jZI1sXtmX0oMDEN9ZHWGeC
ZAxCWTqEpzBayavX66A350tRFOh8RfpdwB+nsd146MAOaJggEJRk6+YZxyMX
LukHPSUdU8Z2AxDWnnCjcFFhj2AjAOCfGUDzgW1ki8GBl1fh4zsheWkrQqUx
aPHFzXYqThD0Wh+pQqHa4oQSinpM+hYHOdxFH7dcuzBvqxhqZLgqUll80jMh
KY/QW6RAjEW0CxkFBYdcLrIIIFCGlMI9Ty6L0ANg9EynvVz+0ZCCT5VaHrpz
gTkny26mJisN8vDqXj4htN/8qL8AtjZlm7Xx2HrXGbb8gbbjyZGGn4c0iYcz
pOGI8Efs15ArefHfhDqiMXb+FSq/xkIeSPj10fxds7aOC9C1+EnJftLkH5SI
DUOOZ/kL+18+CHnRFYx0ZJhzCWiPk6iyNlMJV3MbsKOSZpLEM54pD1Nhp66G
/2XPh4eCbBlmEAgkONTY9n+kN65+1qoj6tPvCAEsXbmZSySOZKWyEU7pYeoy
OC1mLnWD76uL3XipBkTd6V2QuMpH3WkH5dGECwSQsghNxYH+ZdRoWuWyINGU
aXSDeGyHE4rNf10OtTVE8kXWiDKpFx5NoWhmkYguMGZvcCcotzVFEqi/KsPm
e4IS1zMxH+ux/Ur4QAayPK5U2Pt1egX32MvUVeCJNEDTTwjmlAhOxc7WtDOX
nQIWPcXXkowm4UahXzuwHUMNgse0R4QniD5akcDf8baDM3BoxCdkDsLMMgE3
aXgGtxpqwFRd26MM09erpQ+Se2TM+nLMZUs7yJn6WUbSyBSTZ0xiSBuE22nI
drw08ozFnQFK/9J8pgLxfJQrVgp6ziJNQ/KN5z7vFUueYA2c+zdBlHp0cY06
U5XJp4eCdd7Wgv0R/2SZUe8r9IQs/fwXLsXv2jJBdO6rM4iqKgfFvI8ycRa3
25MF3ekfTFb4JNAvGz0a9GpNeEoYXN17GUUuQ7+w0JEVCfkIQaMVxrOQsLD9
2yYVg3GBMyYPW+Dz+HMibrZe94llGrHjbSavBJ/wGXjctale0UYhZYhLlNcN
NU1kpH8kuEr0T3utMsbl5osv97KiKoX3oOzgEwl2cnK7OlGIDztMDEqFvhn4
4oDZU86mmPeBmRxWLlnUFhTutoZBDQHFVuLtszpwYYy1qB9dLtQ0S+miHpre
4Er+b0byZmvT+d7iLI+DaxczALRqozemUmEFGEZcZ+vqSp71zpoT+0GPH0pU
cCy5AUzyNXHkPsboBkEZu0afouDvfnQk2JYr6/VNB/DYVL5xbvvBu3hduuJU
juNLNaboXiZhfGUW/t3/2G3JrZd+Gdunzxmx4j8OTbf+tRZboPLAdQ4FYOOV
T6o3GhOLC1Uw9FqN+w2YIEawqwoX3WV3/4D++3/KeJh+INNPkP8QNWrFbUI2
p2pzrFdUEAj5xE5c+u9U0mX3nxIgyPv1M64/0c9yPyhbo1uqWCZc4Go1T9wY
DCtkPan+x76LCL7O1I+cNbqPiHnsw0vzUZuCg3EHfmIF5NV53xCNSd7Dk11t
nZwTWWjGH0foI+T/G67WmcGHWqN1++oBq5hs+I++uZKYmeWRPctnpECnIDyC
LZPomXUy6XMSlqpPyzYBf/CIvvV/FpKMrTwECiLF82c7JNk14BlJSJozRNZZ
Sf2dH97Qc54OoZwHoVE1wows64Cjs8HVuJN6APza0nR7tO25mtlTsqtsCxgx
7VLvKA9EQ1H/c6KZL9qLDdwnSOjy5MLOTYVH6+WEATVFJ+OfkoM3QVcZAV+S
KfvvQ8Oo303eotIpqKDc4pgeIQaUrcTcJ/jdsjQhyw8UpumqeTxfOo0Q/zgn
VFVJv9VhUvbl4QYNrd8JmXDvvOh13e/+2Pd+I2C329ofA0s9yqFZHZ6uSS09
35ENTCcv1q8meAGG7tH7VWeDEoNFUaJ3M+hlSc3ta+wQnOzIhNbCWInPF9ta
WAbphK00RQTBNU/v8QssC6CBcRg0WVW5nr8T9MxGve2jGC5DzmNPFMMftFmV
orcp+P8KbKppqzGh4F3zZ/uldLi0F4JcepWOteLBeOic115US2CsVA3R+LEu
mwT0eWSkzcu5N4J0Cta9VzUe7xyZcfwrNVv8IHUM6F80DpYigcSYKymhwusd
hAyrr3x07Z0HEImNxs7KrXXEv2ZNqQQtunaRWsUUQ6pb7/5+KRtJX/vnQA8d
zWVAMdEQrt25Gwcow660wfkO+bDeVzDCeiySQgQ16diUji3N+dB7xACmDoik
+TYIwONUEtVD2eGxClBV7VJF/vKqbmkyBmMy92Lw9ikZSJtQANqVkgIbjelQ
zo5z+SISkIztSHdRJ98FJk7XBYwuHQ2Pas0sfmT6N7B4bqpRRbEVQR+J65n+
kdZwe7AUPDRW53IfHAJZAm6tvdlJ0EuaYq7Pa2Hfx6i5kc0zXszY1RFxiZHs
jlHAg5k92S0rMiSyNxAKc6okNMU45CXYreB+7UsEzTEU8iDGC41d7OdzDDN/
dnqh6dthc7VLO9ucAHYdbr/uURLEKC7NTo0jXNUEusGfYftp9cfnf7uA0dpC
xKobzs5pa3B9s3KVq0v9QZ3pUEg8Yyul/E/SLZ5f9OSYsBYzFPDcaZoKX2iN
kX+QuXVYx//ItuFckbxTVEsxd344mfqajQWgsdI5Wr2Di2TATBQT1I3TQMk8
S5U4c9Xc5hkztyrecPYJMA1YCNW6iXgesw8KVj17vYIvY6ByqlCqqWBaQz4Q
qNL/mt3sTnLjBmeHzYntN1MTDoJt9wohAmnLETx0caPgKWnwBaGz7lsjCV+y
u7Q95g4LQG/UZ44QrZqeDY6e9o4PhqHfuU065JVBtC4fyrNIIObkr91fcxyw
kyPBxWFLI+wHtuu63X+9uplJtuUmh0knK7ZGPYfgyVwiyztINfQnoi8CfsFO
RD5BoA6QS4Y6m4p6K7xi2kRpTR5quGBh0aaPKjnPv1anuNm4ogBW/P+Nouzz
y74IWvsZlNS3QnZrushoFugVyy4aVLLL/nWxiu9g8Sm13N1KmZLGshtFTWIh
9kKIDhxYwQ2lKMIr0BYBmToLm1DLOQakp4VYodo0h4m2K9WwNbiHOXYtM7RR
ed4EOOp1wPNq8v/h5kCG69E2Wvnc0hTsD8Vukgc+Yv0pg5iNY5PMImHII9C3
doxT+/fdAu7mhEaYcJ33YEwgbnafOwl8xo0mTp6KOhG6B5yGORpmBD1+TaJc
iSiEeHkDchNtSqOYMGXYjs+QM1UQfQ5VTBcJ44W41fbjRIaVum0G92HYyLY0
12wQB5QxFGsGnYTZLISpAb7itwJgRDUp+Y2vJV0k+GIhCEXNceWWhQjygmw2
BVctwHEIfBIAa1cbroiHpvHpXBHTBwPLapLk7LW+WzP9IzBhzShYYk2h12SF
4wybf/fgEdIGx4lefjrg0RZu3KwYl1fzlof9GEcKPErhudRqiCQC/LcTy81B
XQ5qK8+3S0Wq0lza3FqiE54Vn9Gp2X32R26kP4IVnDbsNkyK4ET36lpfSkmG
t/fNRg0JUcZKSIwI0Cqx3feeIVpdLFhcyVfSqf/Ci4nLJ8D1jxv4ID1AUZT7
YOLN0vOc7KjGDXYn+y1uGEVIJ0ZNCwXbwEwBsegZOPbZUZFsJdjpm1dNsVMB
TanV/ASbuT2DKXkfSR4lqFDW8CuSZkj3LouqHJr+aKtkgBwtHTAgZU/iYFjn
8IDa8MVm40pE2chE/a6NhpXXBBgh+rKpv2LxBf7jkHYoYA2eCq8+CyUuu/vX
ptRzVpO7YcgAUvzKI3SpKbmOnx96zqTWy8Pio1cTX7hEU+Fb4WPuxw1dWIoN
XTbga8V/QyMWga4GNarWN62PfrBJN+CP/vu+Cssadycw+uQ+SU5hY5J96lC8
szpzeXya7yTxwwPFXrR4yoaoybIXvhfqCu9ZdcT6xHmDak79eI3u2paJKimp
/o84cHfucPq0SMuZgfXNGvVFrR1e+/BZu6lSg4Efa5Oa33iNTHAKWWUsr4Sx
t9ppW9LMbx2tFyg89q54OLA49dCBZJT1LZeBR/1HvG6zUET6OAL7zcl4YGcU
pWhEbY4dBLDsXsdE13z47VuEPkuj2+D5U9FiCoji8z+by91FVItFlVaCgKWA
DVoCEAepmlh110CA+rqvPpCA+ABQcNCDJvP2wlX63pUbDl/+YUX2o/kHHXVm
+ZoFanF+gfHSC62PbF2KhLnPQ/kkPUh3mCf+zP4hMVhDN5JldfK83NFKdpHy
1HCwWzwf6Bewp3H2Tur6fdUmI9CSrJIOUt64Mx+riY/SZJAxWOPknGHsna+G
3w+vhtQPrBcwgd9SKwEH/y7/hpwp4AvoAZu35psVj9joT31mCNf5mRlwNMTM
vj6WUDUtxx5/FqxGB0bCWsl4kledq58Vd889rSCinK3wBTbpzw4u4uT8j8MT
kL5lAdksMqynJ+NhdTTwRmCi2aCDkP/NB6Zz9Qr/yd9FTYQmYcELmk3hMju1
rn31SDc3njRdg2BmQzTCYG63bfRriNkJ2CZgiIpXvTl/7vIM/84WHx7Du4o/
pwmyN/bzwcWSbp5GPEOX6OCVMa9FLbt3ih1gsPuCkoQyeOp7ASADirj4zlQ0
2BNACToSoVC793cVUTUqgV71pi0L90A73kZuId9sK8laB1bi+fFMPmlqyAsa
TyzFKM9+/Vul7Vmn92HBAJOFqEC1Egr7Mrdwl8/g0kQ9Yejh9N93wQzFTwaa
a8M6+vTyXW+D0QZh9YUoYWAF7tbW9y8mBPlBQCi1KfnKBZepWoshDnwDRcXF
SJ9RuwcPur8HTtIKeL8nJflh8+HVMLZaOeQMaf72nFUhBvb+0LKHW26h9SGS
v2P+VBaghbJzB7AXj2rziG/9cUZRBAiajZyR6oxF+cA93JHafgZewI7pgLDl
k6qyQSwi28VTVT1JfeMDtpP4n4Dtk8U62AbfzFVAE10i05u97gi0SvatPCEM
bRZTpJPqWCyqYuOl0ZOI25LVPGF0AjI2Y94rZntwMq6e103mVYn2/xifo3PH
sigiDvCIPmK/NuzH8QkL6fgkl6WQQs8XvxORq9Ko+T+GQh9qcXjzfdECHT/Q
yJUpVx48p5DiDaHgzcP8DBoLuTylh4AtHOGOPurMmfWuv6KRgUISiHOabtLs
1GpI9V6x3FEfbaWQjZLTgGHHlys0COsrIM8wA052clVva3EoLUEGL9XtqAe3
gCI4AFWhyDHWJYdlUynyWnyOtLieJFNP6/l9hskqmcloH5UtKjotENZErJOK
co7aedHe7Qxu0w5tAbZWddQcq/BIktgQX5WiOe4eq2lDYsnk1EcqvI6LP0PC
t1EHGE0GbdYcyqg2HnbbIsURNjjHS1YcAgU8oCe4b9DiKE+YeLsvYvZQ1dbR
p0AuKA64X215PCYF5GmsL7wLIxNkJ1mzXeepXIHFXjDP4JQ3QstLlmTKLFpz
HBRvjdrGmqsBRZcoiRWo6xV04wGKXWbvsDwMSLt7ZNc7gU/aCwd9bNKtwNRl
cKvDKdbH8E1hLJRKW4lUeBA8jw/1MK45k/ax2mYOqcrBDjuXbl8eOCZFbiKy
3OTk7teGA3Od6T8v5vIzRJKWDtBd1MJkvc4FmhGYZTYwn4br2YHltj0XnbIi
nePFy2XJF1JVWP3YHoimchaMge/m6sq8SD9Rdp1XlMcHxcVwalX1q1d5mM8H
Y3IMhgCUuv717c7iMdZJ4iYWZW4SYorF2QuNdcPnCndqjDjF741VxYgbibyG
jFJnNd9ibbK2TCOgN7wacmHw0R/Eb33mQ8/uD7UoVzGSFZGuX2W151hIVIOz
anMPG8vAeFukIODYYHS50h3SQvmx9mct4u5cdJ+ZYUMdTlQn5L+mTwF6YUYn
RVBptZ9185c2vzFs3c6Vc+Ibo0Td26MiUtRlpDh7CjqD0RI2HhihQAqZZFVX
XI8IE1POCiWpYxD4gqYLqKijDpIohOuCA2mUkSm7s2SI82NmOLmp84ghYf8z
YBGk+U9WLSrHkjVm8ak08tWvr8njBsnzX+dAWQLEWcF7vFJn5Mczppn37+mH
Re4gaIDYKlbOby2h6ujfBeWt6xJ5nC1SIHGCG7lXGXGAADYOwfpzqwVgYNxJ
CobB4D2T6/AKn73R+f11Aw+lRrNDcsMUjCHO03C56itobBcktw7yA9e3ZsOu
MJ17q5Y+McoWr3U4mYx4Kca97tkdhwq4ytajhW5GKkVdSlBjtbmmeVQWGQF+
0jUnjgUMkcX95eacEYH7NIBDKev451l+6t7hASj0BJBOftxt4SwOC4uhwGTJ
oVmrDDDLqe3m3xiKo6iVT2FTJ4+jCOmNLI7iJQpN2vCMvQzvj50scrLhIHo4
ZpffoM41TGvcBR45AZ/MprdRlCq/deSF68qWr7pjgl6PVW5bxWftEbWG6oxL
JZCcEtiEExycPJ43qqH1+JOB1ei1tSENdLcqxb1f/t46dzl5+L6DIdVh4dOQ
VS7zh5HpeeEyC+lPF9duiYi7XTUIPOxh5tXaJksZMt69N72TRq2PKyWFIYip
dtJIxIiusCPOjvZ+9FFPky8qwP00EKvNL9kZBSlxJ+ViJMVrVNYhgVrmSG3G
qCAEo3HIy8GDy+EkxVqqxGeuQ3DA+VK31lfeGx7Shp++7k38M726bNVNlHwY
gIyck/F8qAUM+IMyXZzgPPSSHX3ZHyYTOkgCuKHnsqcVPX+6X7778MJ+x2s+
qJogM9Yn0qj2AmWn8abaDSLjSBD/nLgCYET+j7J4lBrPJyn/sAtAmxtxo5ny
KydfAzC+ev7/aI35GUidUnZlL7KVJtWvl7zmAxGtARMPm/+mP41xeJ+ia2EK
zGXOVaco4DxR8+gCXkFT3u2exNzS1K592ekm6k2fy4l30oIW3uAQUrF3934i
u0ENqX3bLzQvC4GqfyYj9QF0+he4Lz3fbMhG9rcjVw+SktjcFmJOxnE0QygO
uJne/KgoeHOSZt+scLufsoYjNSzyU47PrcBkfVxQclCZ055w0K2zSjUAA1Hf
MktINr9aKhj1f4tptJ1DQUsqOuxH7uYnZgCfbs0Y9akpFXuCGpwziIxr6J0r
YNqWoNW1sAkVNpklWI2qeol2J2tR10uSqfH/dVGvq7m5COqIw599/1zjfG3E
CYCiBPxk195+CzkkhMlMD0H8XaB24m/vtkhOn3jhUBMi/fy3wmdWkDnTjNFU
HnoQbVScOrl2+tnA4BoYqmdLZ0YTcjgRSIGu0g2BHFPGE8sDtEvs6GBYsOAa
xXBNz0lXEz1/T6XJS85bTKighPmNacH+PPd+tLhg67Ntkm7jqkMnwXK50a+Z
sd8K6FXFQqh1vsmgI5mWcWlRLLsFEIkatNGfv87kTl2Lyn6GrFTqLpzaZZ1q
MnyMYj8YtT1yIqwKSnoEdzWVdcuNtEun+R+11dqvnpJ0QWfWDIQfPQNE7DoF
W94ibhE95XaYFqxTkmkDm1w9pl/WMVHAYhsqZ8oSCKAyvnqJ5YbUYCrUiZr4
3avn0SLagziYQw5tFw7oqpuKFAjsvkXOT+OTm+9S47uFwTu0Kjy7tWo9DPsg
KZ7nePEL3e53Q9Hmd0gKYxOXmBjH/0zEgd0/5DKYCD6NIwM1EG/mtSZenMNI
TQXZNGopPIQNbVLaQ868CqWpHCAagQc86x/pYeYhbOoS2msVsRThLi04XsBV
XitwqoXu7rzlKcGWw5L+R+Ot88vwYVJG11fsTo5X9RRSz1FjrgtxD8Zg26qy
glNP1J0/aIxttWdwx1OX+1JnwUssJtCFR6JBkmYuPMFtmtboQrm6PgNPPol5
sc9vIJMCTq8DAZBDOJbc/58ZTMl82q1ZcY2d5VjWz0uJ7nDyRxZzj2Jo8hhI
8ENBYkQhJfx5cDcfhxZkMujP3WmuPOejkJvZ3UpDm1AN6Lw9g5bR8bDLpzcc
aSwK76GnkNaq3AHmrLJssRLgXjC5NJuuwRvqUrImRgpHZbWjkAZ/HwMpbtTA
pHKIECBjoLxUt3hGP0rmLeTXgFMyRgu2NnNGV/BibJ2hr9caXqE9Uxxfp4ET
hUgMZ9n7zUObkPgQq4WoQpqdyjjDJ284gDv5X9bZqclMpiUb0QSK5r8T/Un/
M3aVv2DVRpQysX9ufKUCa2QR1/db0/3ZxcG08S1KiHVzv4NOF5p7lsNQuC08
JI9HK5XcFk67SWCyDJiuVT3GxeD/A4iQzMLxMwCqbAtQ6jqziG7ut/TTc61H
WmF9P37CAG2z4uG5rybibMV4iI4Z7bJrjgTOH1Tm+542WzYdk5+8sPvi3+zv
34n8Y63fZMg4sLlqUkMpgZo6udJBpUXNOmIX2XkvlzDjJFzqcY90Ma0qq08A
sh50B7O/jY7THUq0Yc3wNC6DiqnwqcmkPj2ArV2qXl54ukBdCpKodokKSESj
vRpvGd5L78bgzjBs0XEOQYY2hd/yHzwhcQXJVtXRQQ5J2ahdmaBpRPpZTkUn
Ae/mPwtQ9sxJ0vDQfUB1I3+9y+oaAEMh76VaPYXHlRlz5QNnhbbrhGez/9p0
0UWI1XHSrDFEO7h9qkP6Jgv5LuIYIakoRf+SB+M7TX70OCyr8TGYzdFOFaui
mUennt78SBTgBrcPM1gDesqUmmlrKMIqHH5ycNi0vpQaFu48aWNBYbyErRuq
FIZh/uylddFHsHUw39XJgeUY1sox7uKHE+qy+z5uTjMZFOUq9JAbTx7Bqu8b
hkfZFc/b9slpRQvLgV0vzDrzDgxiyK6TbieEn2jNm+yqZMDy9C2fKQG8ERZk
oRdwIa0Iw+vUkoBp1O9CUje4MzQUwkjLi/HpcsJfDowdfmrpgw2LaJaQIVzC
J/z/K3cnNO/Jl7q972ALFbhjjZyLIUMmfiNGZbi/U9FCKS/Ri9mtmJEtRAPU
0cXvExyfAE27AscP1UXlsWIQU5KpokByn0aNhlk4noK6CA9spbMsMOYQIb6K
umFNR2Q2bPs45yxWefa4l8LzVjlA1BadvPGNtpPag2KlPEhnDopewtYzAVEO
JXIsh6/rhClBn0yB+ZGV5e8US/5xGCZ/WaUo18detv8cllWsYTGp/XJRS6K1
FHaDPkr6kJbXe00V0/8tk258q1IGFT3mKJ0zy3SE/r8B3T1BrJHWkKQekKCe
gxKt9ZFV4K+yqA/UcD6N3CgNqeDBE2EVJaWAHpZfYsmVzecMVPVDWRNIBUqY
GDt3I0+1IUDWQu0mM6R3YCHU8ca2tZuNKiWFvrTVAt15CFoaIxYHD05IJQLz
z518yULd8KgURC5ur1v2cqs9TDIPpL3X5xUTAP6US265J1h7iZQffVIWJZod
WxB5Vii2+Xr6dwwWC05NesJuQzjC2ID1cyEmnebwCCDeOS51hFOdp8FBcirr
/CaBPAYC68DxwB/FU/2uYGb9PZg4IbHB2rtxYrWpuu88HHITAxMENqk+7uUv
YUivpXSWqHWuy48/GCtGrjLCppS6TSzWlTAtwF4ysFbX8pKPvlmGUU0bccuf
iwG5uVLgdMTYPYYfBQezxmBEp0K3G5jMYAEsShnLnmoftGuK7SwwS1o2Al6M
ohvfksxErAy+FLscoM+UnggXeFny2B4US+enKwh39T/lrIZZ+pyHvAQrpAMA
jGIPTiXF58ijmCtFNL5z95vH5vMlqSPgr0tNFi0QzcVkR4iY8KeGqx4p168R
9hx2LAhGqH/I6aNiO/548vqKAG3oI8qCzJM5GQVpKVuo/IAncMLZj1kWXyrm
Do4rko3YfeoKqxpj+Xvuw58LCCr5WzI2ghJb6+InoiHiHpBV1EQYJsbeXP/F
lzdGEqeA6Q+3Ynf60n69vnQ34W7YMctKhakQZUAak/Qc8SQyywv9n5NYETvq
z9FgLictIYyYot5Og7iaxWKqHkfSc1Dt0T72QrxJL7JDji6yoUTzzGQnNRQC
IfzOFPxYcgovyVdCiGofBjge1HRPiRNwNRLh6GOCTpVdIimMi7zPTunDCf1r
9p4w+OdP4+RUjKPm271ZcE/aHOHmD73y/9eQHbAyI+CgLYkcLZgIjwCc9WI4
fKb4IZ6EvbTaaEhS/XBZZj5JExLgyupsjU4C0W8CeSzvbNiNKbortS5uCJUT
SRj6OyzzcMtFbix2NvrQ8Y2B06h2aLzXsDJ4YIYRLweoaGbeEgYKQ7T+oGRg
eGzOYvVNMHGTdOzNIzgq5TbTsGFw9s5u2E6FXM/fwYqZcgogar+4gjtJISvD
9mV7bEOrJmsHRMQsYzUym+wGoewhrfos/SYf2cZx0xnimBoY0clP5fFIAVfn
jp2NJXDseD+zhSJou42lzvdbw2SgZxnz7qLasaAze19Kf20WzmVRZD0Baw2U
8bhf/iiJZzdPvdVfJ+dkEu78IZvjiEZx66n6ThaKz0YtqcuKpwQ6BxKHb6Ly
uLWpfziGInrtgrip/L/o7w1UmYpxXW2NeUHmdbF+GrWjDrhm41BwJyCYN+wW
y9oOZeX2bfK81Qu0yEBNl3AlfayaM++I/i4rNz3SwnROw9zkWiuffHL0sMIm
K3FU5+sRKfVC6qzbKT9lQviFR6DxWr1aHJt5Uu2d4gceKc3j4E0W733TrSqs
Ba0FH06Uynp4TbdrcPxvGmOtotWLjgiSEnAyRRIR5o1n19Ky3VkAaLqa1jb7
BSRWdVsjB/8bCK1WtTRE1vhQ21TW0RrmuN9mjj/F/NDL8DrL4GfJWyiV78wA
SzV9q+wtH7SKlFGIklCBvbhMLyoJpHtqIggFNaIYk2uM8NYbufdWB8kGV6Xb
5HJPkBSHmjVLOEXZSwzqhuC31S8XaUqacHz2zVnhhU1Xnuoa4WCx44m20hzC
NHNgoRKt8FxytciXiQr7/MUsnExezfOtsZKSBI9h9AVdcolK5/3oGMTwpJey
oNPsnA+lrovDZfZYp1hJOo+bAO8Qsi+t1i6ZRamfGD+eAr7C9FzvV9TtXllQ
8YJAQjMEGpQLeEvs+MMY5T5qqeBrcgKCfFBmlMsCSjPXDrhCVkizUuJaVbmw
+/BvV0tG+Y6X5RNxY5Besg8Lxfhj8EQ+wFF7lmBQXHeu87cPPcH/v7aATGqo
lPHSYFt/nOSJV4VP6e5ebXFgOyEtulcNgUR7IGgnqas+X/+4NdwL1rY/4P15
FYj8ZVd7YpJpH4DsnaYUR/Ns2R6rTx4bj+yqYG4SRe2Ug6kY3TiJg9B4iMUs
6r4CxUC/cqYHjptoCAFrtn1QSbAV8+EMh/Vqo5oti0tmTp/UcYqZ2WtKFAoa
trWrbm4HNYdW3PP3SG7XNirOTNCZvEW0UsbeG/WmFwRndEsmS2lrZX7sRmC4
7hDmpCy0lg/xSk5B7RS9cu6+HMAT45rw08ZERNkzgONp8lYHMUwBSXZqIh4l
7lx9mR4cvRpSfEKyF+OKHrv86xh0WA6kMvztwSTly7TSFh6ZuC2niA9TfDq9
UghEI3niIGhcn4kT6VxlDLG1Cnv+oNgRPiKmOvHKzXuC8ivbZ/FZFxbTTRwl
txfMHQk8XM+EV6ggyQCIK4UFTqQb/4DOMrvImpkrvDd0Ij1iADPurtL2UACk
h7dc7sPdkk2uDJDFJqH2ewH6Wgk80IlF5557e9juw4vWOGw1chFPqZdSQpz5
E6VfoHUpA1VQ2tc0utgfGae+enA+29DrKiP2dCP8Rsc+qrgRg4IWiuKv14Ya
q4VcHOI/2E1o7wItOIDqS911SR9Z5koYJ5uobHx5lSD97lFWLAh9Lem/J9NY
f3sGAgLTNiRcr26BEi4M7Pb8+AmaqG2RIO41ovdpAnSmhljZXUJdEgqHgPwF
NIYBaj74pznNzgCbYGg/tDluKeXHdTng1Xl2rYi7+INuYd+4noC6Ex6AxDn9
ItsbGVOdVO5Zy/0jV5Unoif2yv0rUrk8qt3D17P2lM2KvmSttt4aoBCF/0MW
bY2mE1qh6YDjPTnF5n+09zLTlsovIFzXfpXm6Hl/pjlHeEBL35TdqkNMv59c
M0G9/yWbL6KM8cBADhMLzzsVKIO+ZDyVIxoMTfxCyFg4SWUAgZ7P/Q6qtPbJ
8Uc+psU2iV5DHDrHjJu8YIwvYnr8/6n3suu9PLAYIjh+nnQEmzKRKWXDSLId
ktVDA0B8SsGwpBjbUf7wr37TN9W078TSLAHqj23nUTdNtDY23TlCLAX5K1mO
Wc7MJ9ZSNoTwqMLliIrnlNf2Cvz40Dkgbcc2YNBTsSq4G5/udz8BlK5i9kQE
YFnWhs0lh4bgnPkBMgd0cBABxSUNokCerD4TYTMGn5PEeGhTLOJAmHL2Fl+M
MAxGDnBxAIN6qgtqddeoc1wZffWunDDVGHj6CgIzTCoaqRs6P+ckXb4y4lVx
a+5KlcuC1u8tDNQY2Gdpx7GfpDhvoLpJd3kkZoq62U3LHUhMIlIcvTlHCvhI
8NW9ccDnaYqP8su7X4MxoPMm/NpFIQFeBuS0Y2EzUWj0xR72Vtnx8FVYl1BU
FHlXgDGcPPZDbqjc3WAYB0br+FvTTWinBqv7+QoMIkluTH97JsGv8w3U8n+r
Ma5KgVtbQWXy+YkqPDiFDw/kZgOB5HKEcWO2e2OxooJl3yXC5d1AwXUvpYD3
IWNp4crVk3pF1NoMsRXIZAr9rLAr7TlhicHb9wlm7wI0ZWu1HbWB/U3IORW5
NOQ/+SHOC0xQH9w2VjLN8I/P2FzVqImFYUUk+qweCFehE3yTxOYwwTfaEjkQ
8kcrMQvvE880aHkVvyAJaQr9S7kUdtem7p7IT4KM0htyVzyWmgc2GOBBOYUl
gcxuhjpeKst+NtPd7PUwgzu9cN3WU61HXVa9giFiCHZFAmfYX0oNYE/1j3af
rhF/PaTvvQFQ95+j6OTNmpBXBjMCuEIZEx+uJsXetKxGHIzfx91ayCaO3sy1
dgCC9A+UyMXZ+YGfh8hX6HAkKpK3JEywumYs8iGp2DILOdkasnRgeO7Mtiio
YkAdbXIkhHPmxOOTkwf8affu014xylpvgjsB4DK4UtA2egWKdK8hqbRhkOmy
JBPqIn25WmC1gx9Ys5egGoePZbCg00+pLHs6lznIoR69VmR9OSk4d7cjmlzt
2OQYKIr89ZvaL1wdNF4hRRWhYsblAqMgCjg3Uj6619CyRK6Vt+xFwD92Catz
mgbvZoyBL9/BmFEHWtb6fOEauQxTvJ7YZeoSz4PSRhRQ6WDQPHOAtVjRvpF+
IPkK/rXtslf1O+waMYY2Ffpire7dFg8G0DlKSCyCbKVwYEpEAJ550LcYCX1n
d8FfsYvNca+lEGwxYkZMCnFksLfMMATGo5j175dh66kHVsy1Ye3SwrqUZ0k6
hLnILBSZeAlIykBWBbgHacHWW6HmUF/6C9FxbjciMg/fWMNeZw+4aifj79zV
0TlhOOHKzyg04S0shFGkXxFv5H3epfc7amf34DvLe0BW3s3PlagDDvuL++9n
JbHbCiKT4UGQ1zByMsY4gXGMho2vhe1FibAfVJN5wRjnKWKaF1FXPrSIHJJP
TdmL1neoNAI3Z7+AdDp3mj8AbACqVJMQvULvNongBexdJXoVxs/s3RqmcCqe
hLNKFFjcFJgbnISiWgFwFHUvaFRKvIc2Ba+YgJuocWmHUC83J2wz7ieV5p1n
j5maq4j1bNAyztK7COtdOKJ26QrcgtKjUWeoF08M4/lLHT/z9MwWoOD/LAro
W5aqk4zpAs2Drw2tUxX6WnRoYEwceHzoXAfOYMHGeZ/an58RISqn+lpMy0ei
SiKkEUYNOU6Wg6wR0AMorJONY4ZxCVi8MJXRXDCesV5UMULK/niV3A+x8NZR
xndzuo1ALudWCv+OIdmIxPM07WnCQLv9ynJ2LGIEL8b71sb/w866bKYDTcvH
fMoZeqW2pUDwQoVG2tnrxhoqlcw/O1AshYGKtip/52E9KCky41eAmM1+V4KB
389T+ZnAcTSSH75JxmMhiWtksPmj51/1Q6iZXhnoEmntDbcgrBCprBnV5Ets
cIUdvzkX83y317OIcyVbtxHvZgRYTepM2GP13DlcNbb9T+z9j3ZJIDT7Ml5B
QuKa15ygHQjLc/jTaTQUhIaNBlJZ0dttdX+rcezLd+aUqalq5Eolik/qUpfY
Y47c02W56NbRCSujFwC7vMmPkO0ekzoDt/PC8yQaa7Q3txwiwIbHKyaN65NN
PNoZi86gUMb0CIz/wxkIYvVQmSvrnTz9C7Z887tN6rs07Lii/Mjlu6+Xq70l
qacmkKwU8lX3RoMLi9zisxCmYycdD81dHxptkpftJCoxEufPI79JEzYdWXnU
nHnS6a8RA7qgaEhPR0ZUyRwAOiu+ENwrWxh0SeKXUjkrjY5bzbaK8wO7YyAy
4CfiQhfNEUxwtVxMLKZfgZt/0j3JGRscoyRtCMTlVg8B5J/3XP2BfQNg7H7j
z529dHUm2XS1F8QKIdLt3S0rr0bOLCEefaSxN/R9wJw4eJcIzEZvt16DCVrU
D56zyyFi9ad6sVM9d90/J23Zlq1q5P0gwc/43D8q+YyeWH4Ga9xSL+5HnWlp
ViLs5miIICP0Bik0i4C3d8RQfog7spe0Rqo8eOpeUptGWdbR32tGwmysQHkv
CzxmDgCyk59+HRVqJScj1HoRPJTmN0nbKgZ3txb+510yPjxZoeEL2PnyV2K/
OLepL+lktZPDUxdtZJdIQ55HxycyZ26cAxZNpxA852HX7QpV0i2rFMNbZlGd
R7O0PXhbE2FpgkqccR2oncG4AtagG5kpsWi5pI9/MID6M/kb4WVZpn32YnI8
ogpSp4E7QYuilOHG24jVAvroLpmPe3Wd+dA1JLcVi3OHZ64EoMbc2GVju0qj
cZl9RhRke952Uba8S+vsgs0GBn2QysEMSLGsR9pYmRjVIfvJe8sajckYG3u4
J68bbNxWfiqTKwZCUIR2NM2z18DsA5hLDozCvBQj8tNwBVXTp/RjXVguyGnk
XS5UKFgMV9p04nLcQfb4Y0no7i8xSUUB143vf1agn0GHnDgb7YN+4gPJOxOR
GUn0NhN7y04Vp4Z/mmXwEBi2zSXyzL1uJZh47KAhdZ5ilAnwYlGe0pP3TM1t
30Xxh1H6Yha9KE9FvCTZgwWt9uoVA8IOpHhdaKTZTPtSv3WaX9EdEnB1QULV
jtrAANeZ6BtIfCjJpoQHakTGs05IQ333FZzoEhwKq1R+HQryTwYJM4+klIFE
8w4WNf/qF7X/mEYTPkq3iGlaS1HM9GQb6bYF73nq1ASZugSkiMbEZ7tgDOBI
KfaRQDfxQzToyxMRiBcmY/wrSSPjLUpTbx9oMoqz5D8vv35D/ZYFmJuYucm9
oXzGCBGxdoh5X+La89TJV+EgZn5PToUva2xlACgXEchBlVQirCUFT+lpjb4U
5rqHJjlp1oLI0V1c/HrbgHCz9f1E64bfVsGOyRsvlf5KAdamSy6r7mAtjk29
MT6h6a05EW9lhcJfQeYt08crep9h8ilhM2Frb0UPvAWxw0Kowh25ZakIagnA
XMVHDyx5MeFLs+1x9nxfvO56sQs2YdaITRqcynkJXUfJyW8No//MewJnluq2
zc3dLKRyVvINq0KY0ZBrND2R0vC1ssFXcYXp7WJdu8OgcRSgl0QQ0EFlASNa
3NGA2X4CE+KKk/fyV5kfHMLXOstXQlIPDPd0S5ITZRdW7ag+aMvOKO2preIa
BPAYAlIBfH7zWTIPnF6BFXZP/6ykz3+t5Xu6MHrjP7cQLq1degraOkKLY/NT
2WCqhtrKSfrioEam5C/5cSUA89nGmeDyN3CPkMzq49sdcsEZmrRC8Rbix+H2
ya48QE0I/ihM9iJL7RLqdBmvll0nnqRi0H+ApvqJ65OGWZC6gdswdGMif4Kq
An6BnAFDZLU0yLD3rBE0H+uLutTs55otcl/3iuH4LVbsHOSICvkZt+cdD2pA
BdMUXa21vDWdKTuEjuDG1ogtQBSgXSE/HvtSMfSDmKIxAQMv9Plk37RFct6+
OAU5UXotTAoXLxIWVg1Lnlb9Oa1GYx9omUfkxFB3oKigweW7NmL9Xki5g1KZ
157Yw94BjFm2DDMZBbr2IjxAKuIQ8OBoXdgqlbhkqoXBQS/5vhij1/kZw5ri
piGLzniXB8FpXrW2pL6tLe7p6mwWOA57gXhVn4aQpSSOBP7RbvoII51/cFos
4dh+9j6znLyUhUv+zSf6GNfLlAQZEe67YGSTNezgB2AxuEHWKCIkK2XogQbi
JI5fCQt2QsPgAsBa2xgVsj8yWGGQJYu78QqI07VInwymrL1+dF6pCjAKohL9
f9O2Qh1Cz0BjaXcrJ7u+lgEk9lEBnu2QCScHU9Mh2tPlCspxpdUoNeBT/f+K
Yewsb3tlYSB7szGdKByoBIkwAUidWedd7bsqz7sDKb4jtvxo4PfCEuqqzOtd
+Y/9rDG07Pviny6tzoKaktbYPoGteIAgjagXDv921utjY96/3gNupukoJ/VF
+VTJG7Gz1iYk2p9w1LAbXOzlSvnxtG1kvUhiu+j7AR6zmFa1CmyYd/zi+iK1
NT5/rRV14+N3ZHOPNFj13KC51PjpgNYKWFPnnVM4fodRy5jIbFtG0MXedvG3
o3U9zMveZGSadLZfBU7gyiok1ifLMQcDIlrFC5vNaW+wqTbKTwy1uZkAFyvV
gJW8uSpNO0EsMFLquJP6K1matZWZCDIh1p89BkM3aXS1pdib1pT1K4L6vQ28
iQB5aCgqsavtvyc18QUhU6tSmLRnjN1ledlUV2oEBkWpWn4DcSpkJ6q6c05V
chU1KwYtNmiw+hCfOsHm6SOL3bd075j7BT4LwiCn3JeLA9NkD4H2uwXZ3bxr
FdCJAkUfoubtBx+plH//1ISgM8GyrWraecLAmfrI/rFIBDdTUB5GMX0WGBpT
/W/n0fuxsCnz8xv7YD033GTWe2kViKpIyFiIJ65/jt22SmRF/1e4Y86/CauJ
IZ5DPA33zYZ8KrFuT0Eq8PdH1B+OhSDhJqtxa7FdDiXST5FG5EeDOUYqiIVC
TwPR0DkMou7Csw6ImifYaIvwka9HaZ+sHVD4sRLTPJi5zKs4sG2FL0osuzgZ
/Nz2Q3yBi/JpMsz6Pgvt183mDkGqN24uxSpS826L3giPVt0gQuzux0gJsuxP
Wtl7cwwadGL9EP+Py8D3oEYQ7X3tvK3N9berEgOCMsTxRVT6k5D2Lon+5Kp0
JqDebCuZTCcQ4EUWf7aJgztrbNntZ2lC+/MJTnxKMYuoF2ahjXMH9a7t2QcZ
wAIcL1/Q/An/7CBvp02J2w7MfQeIPiggsOvSoKvOTgnq6pqEwm4TMf2lrzZV
1i07wdC0Te5cntKeEqVJsNI25Dl+OL6TswV/8myl9BDzIQdiMLMyImRkFTim
XZhwredPJkzXPFeHzlnTG8vuqJyMqQm6nF4el9BLL3EpdKsOx5ps/ZsmQazy
rUIPqf513VSJAsPskc3lRn5Jr8s5nYtSMPv1QiBLu+xrUnjK5v9AZU82Sjrk
xVfr/T/e+fqYuzzN/6xwt1HGSrFnC0HxJPxB3zSzpC0Qmf0IhaJRdYppcr/F
Au2LMU9ozrEXVEZhntSidCIzMcFdsh+FAHDXSljfK7D62mDemW3UqmFIxwgn
Rhw5T51B9gRUWdsfhgkNQxxaA8nKwa6+TYq9nL0V+gx3iNMMXVK1tuHDUi1O
L6pgBc5OUGowUDQb2pLVFs++02j1ZZDrFuUUzt4U1HBDF2JOJhoaD16+S85P
Hl1k2Nkdp3+pV5nfEZr92dbYYcdHCimVCG6T6PHNZNYKqBENXxpYRXMWACwn
iZiu9T7ze9r1z/5Ji09RD0vsGBVj3eshnMAg0yNA6fQ1eb9jTlWYFkqElya7
GvLRvY/D6YDKF+nmux4t/48MTrdiEVTMLVL2jCC+y61mhzmnD22gQFJSq8Bb
X20RUFrDA9QPbLpjP7DN4+VkIgWposD23IzH+cRiZRTOIVfFcPK2+rZkDhUt
/RQ3qibU2rlKn2XMLkEZZ3j/7nZFHtoXLVPdXFRZ2RPEaapp2fs2S/cs3tRn
sH+0nJZ0va7lK85hJ80N5MKqlo3TGEvvu/gYZxZTGD0UX4gzpvFROnJ9ft9K
jilKUULewawAPQ4iK83/1wP0IY7YIALdwjV6shf1UIFwD2p8vo+mH1QfYZe/
CGVZNNH/1I5W8H4nUcQOilNW5xvoyQXdJkzuTPMoSlXYp7JbrS/DesPr8V0N
4u5VM44CBA4HjxTwBfjVUquf5l+FR6IK3HWsae7EoJr+YyIZcsSQZxH6jvuA
zptr+lHNN6zMK8x2ZYJ+vAFW0B5A9bbnFtxT9WtihQuAg4gOTZa22RWMm9+Q
34iwD6kjo47qMO319G+3taEZF+Ov0UyiWqOAXCWYLTZry+IWG5GtLdrtGTMe
MdEAKBP6KiEOOWnuxJmHkUqYOuMtV5Hn4IgKOz2rjsBz4BhH1PTj+zvzZbsC
6FpKbiDucA6CZm8ObrJp+ViP2/HbSwBFYLEwW8Hjoj7feZov8f9x0Yz+FBP0
1Rqb/SYbgaNXkRKLOXY9HiyJBYtA0Sdl/oCbEF9TxagGI3rvFr380IagG3Sf
O4x8uVhWx5m9oyex34mhCvTYFye/sI1tu5nCvLcQoMeNj/VUoilbCd0uGBpp
hAWSwT+1mRb9mMJR/6CAot/PphS87JJCedAWlps83k5pCB7anuZEGBW4w2be
EVA3l7t1Iph4Ao3dTJ8Gfihlv2bp9tFB8UP2jZLMdTYqEjYtMVmqtmJd6T28
DcNubSDGpW8uM6TIpLzZmdhNEKXz0rTMJv++4G1MiJJHZ837MDTyVRXPwX6V
15MOB40EgG/5mUrR7IjpziAOPf8Td9uONBntTnxvbIXRZEsyyTYF0JRJRKKa
FM6bvp1uH/SHmVntGxOBimGPVm+EgbP1rsKffAPouPS60MUDdlutN7zJY/TI
qgbaUBHYAThX1eZHRSC4n0v0qyvVZ7miaR8fH4wn7OvmYvrNdVuTdILcW5u0
PSXekfhbpYw6cEvYNwklva5P9xZx51X8KcGys4zlIj7thEbVYa5F9tssb/lb
hLju1by6n89aoY1SGjpQRcRYmHGpa5dNWeoDGbbLJn3dUV/2ndX8e6qlK2O3
2MX8ur3FeNy/8nJu8yYp7xwB5E06N/758xs0IF5YvSQ1aG4CTnPIt81UUw7S
LWBWrj9KPWl6iRn6HDDZ69oJ85aJFrvMtAJnYZDqRksYUpQQ8tSs3XO55Ync
x5NxVwXResSsnTfr00mMq+jdPiq2OKPALWVai0qJJQKEgUpbxnIHA4R54iAS
hLe0azysMxIFlR3NuDAdt+S7yuWkDoUPkp09hDH8oYXQi6rfxbvjR+fBpCTg
KTEMIpf2kLo3k8TtGbpodSX8eU92eYch1oKOF7WBLoF6Du/mlSqet7kUaKjh
DXMfjUqacx4CK63D735DE+e9///gS7jPtmfRaHSVxKLMHxE7eUYKedYHJ8oX
w3V5JiGRhLZZQH6KmGx/xBwOLtGUw+Jgx1xfSzs9E3puvcYZcU9y3HZ2mvpv
MxqZWXl4MMnEvMufsqCXivVGunKVBdMvIib6jZ8LGdpypa6EutkDbxJUOCXT
/02KduO6RQkdVyRJvfHMECCnfcxCJX1AwbCCqyeGgRlb7OtJhZ7taHu7vPT/
ilWFjSDPBwjAZsibMK3TKzst5X9CTpZ0MfuT1Z+6ge7T0GLZjhvtGDz3wYG9
kCiuHS0V3HRHqOPq/UeFQGnr6Z/10WEHfuUO954UwzozYDwt8J6yVEds4+/L
Uij+brf1qLhT6Vy9Opz5rp4PMFmXbayRw2GxFHziD9v/j1C9FT/viZHXZ9tt
42kkD2oyNqdujpkCGjtIKEbGuVSrdjxCJlYq/iAFplG5qU79LayhoYQ+jJ3B
dXV6RHnw5HeDE1dLUZ83R4tDUKlP9beDU5DGO7Awm2RThaS7a9RImQMhgWzg
Uh9y5ViD8hGsn9/w4kgNZfwvQPE5/N+tgPXF4FNIGg+T2QRtGeDYyaoRQEPO
YNa24az6Xy+rW8CDOEg+nTsWPdai9HpJVcfqx+Yfj/LP9OIr5Rle3UOMNgv+
Nhti/ddCLlrtm8GHA0UZpsTO4pIllb3d4qHzFmTVL4dOG1oUn+qCBFy2y8hr
9fKwnsDeev6a58+H+8l5FcY/CjXH/dryCgmKbqYM7SPFtP0TLbGppbFf4OIN
KPiYDJIUaMbKulbI5ERZynyycDJVRmOJW7PESt5JL87S6du0TpqhgElahCPr
bK3hiBP1u0ioqku2U7sh9gxHmdvNU+2Ov/XyU85zlChcsAWFZ8usoQhDhrkR
5KFw7lUS4OFh08mSaPZLRdeMpJ/F7d4VYom/i7Lc0+eWchcVrWBLbPH9ZO/X
38IbepMhRc4zQSH/UB2luc/0+JV1L6BcbRaQg1Sq4Ieq8C1MKX03nvk1OAIP
naIoy4TDhThPiswj2YMoxdLiGZGOqfSto4Iap/VqAs208dPXvHwJFVVjgZ8U
H9NJIzYR2RQky3mXi+bWHR+t985SM7Vvv8iyqSPR9w0UhuP2S2ZEgZQ3L0Bo
nLTR6ik/182gxJSxxcRgKH5KxJCj3uJAhfZR+YmSMKa8EKI4gDLXlIEiCpy7
2IZCwWJF5JAOBZ7OmY+jiLCOYvG+annPkirue1Ji8TPHeRmfr8GXgmNFqCBz
IhSq150zGw+6cbCkCHfui9P+ybdSe9Ei/kEsu3Uw+LevMR5X/huF4+8qanY8
woxGb5eQcRibWPr+7LXzEtzoo9Jp0/BsA5SEpt6h+b1t1uQpGBGiTLJbHYlb
SMMLen2QuYz9dWRC8tR7XLtBpnIQbyStoMPttKtSJt96A+D7AAseaaopioFq
I0qvmyP2eDK50RG4Is93tkCuQ+MLGwnzNsEk0jgqgep3aXgQ+8oMq0HRXOrB
svP2h6CjYUImWMsmZkHsvVViAZV0klhu4ib+HUlsz2nk2eO1/BY/55+N025u
55DNvfvzCKSO6/Q2X31+thePnkwcbSEA/vjcoxWu5QWmHnzO/hAyc6sLnCNK
rDqR92RGxGY7N7Du5ApKkubREysgaSEAsux5OVON0vZS4NOsN3tkkZwYHLhE
+zUqGLW9mth5SMLxGcSdnT+hGrCyXq9AljK/aRJxgMsIRJ4Iubg8ZfAtRzV0
QEiOo1bqtwyIYkDyZxaXCYaOy4KSXT51H2l1W+4FEU/smLbwFirBJV41izHM
GtFfIcUyHb+RqgydAeY1ir8RYK7ZamN96QtAbUqMeoWxzK6vuvA/RlsLtFSB
ioNzgVrdMlCpgSFTsMwoYLSGGS2Nfxb/h6EUruChVjNlx4kIS/0Yx0Zw49hr
/N37Rx/I+7hdvChKBK1WXwSYE814uILWsiLHdw2MqJgENF5NDY9IQerVdpX7
k7mRXoLkgLYeBb1H9glLJT9VbCnLtyC/PN8vyhOXXy+WLk7ZYAbd5W8bn9AB
q001mdQOWJLr/PCsXPEBlV+6/vQpxZS0e7pKE9z5QzFZLOMLeBPg0M4zPzZg
guCOuzCoo3IXLLvrJ+k7qy+Bx0OdfRI9xODbjYz7BNFTxAunj6SQN+jEeasn
5LAcQgxi4UKss6OKQoghi/WTlq9X3fdQ7bxZPbaErKjLT4XkTpiastromaHm
lMn0MtXHaStRBT0t06F2/eW6YSvfgU8Ejkm0W7qu/8LuLwUUCbcM+4MKnC03
9Wvvj9LWLBLi3JsCEyUwJDDpibEjdx2d/Koc/9KnwoVipCbaRIDmmYf+MQEe
Hrh7KaeQr7nHchsc1qrlDiWSMETC56JT9fuTHuN5d2OFq71BnOfG5WIscrbb
tLCFAmFBHsyqSCpC24lkj3yY6WNo6d/js5DZPxEsli3ij8Na6Qy8btKv10/F
qNZPGuindmo7J/+gcTYHqzrY97qvFrkBQDyump8vaTy2XnaLe4gasQkRDHif
Lw7gqbtjPwTdcLYk/LaGdflGO+Py7mWxLcILSEf3c3NZljchiqeJDxaM1Qq6
SXI+3qhE2kz+wZWV9N9FnRElsaeI858YcFMAXTgBBMsTAXp7B+geu6zTvRVp
pQT7ZYN7m3IUKIkHtmk1Zs73pvH8dtOdsC9f51MO/zms17d56A66LjpgxNhC
bnN3QO61ek5EoLe7yZXEsApo6QcG7H+9Qhq7CCK/T9zijAjNe9dEXrltO+1i
2y8+ezTFpVBW6yYtCsiEH5OWmjKvyO3FGCbno1oQNHZ2ZwR+dvLw6Qao3Zm3
vLutfYs35gyJZn03QQPAlwPr7JNO6XsRrlF5YUD+BKTiTziYDN6kTfwBxa9A
dCwsoBefu5h3F/SdQh9zcFrcf3Dm2rXTaopGl28h30aqkxw677H5ulUoFiwq
R3Ao7cFLgKbBmyqFfWFbPHInPhgY8kVcDqc/e5TBVCXyb1Y47HwelstS1Ymy
xlJZv+LCimotBsVwVuPtRWY2owyQiHJnvC8Z+jzPsoF3yroE6ELXt12IBiKu
eCAD0wt9ur39UXLNYJu7C5wzJZ4WGgjak3K663eiN8vgsuTG19Gyttt5xCTL
PtZEcZnxxKINEeDrbeueGCOutNRi8Ub02A4oFVT/t1MlanGdrpsCyQrDNZE3
iQVdsCVAws2HsDCq8HP3O7aUmJWPzujsNObaYqgUvCc4whONFiJX9S7oADwX
SP4k3jF5LD+G4dnrntieVLrSkiU453gqafeHl++uKZV2rbsl+F8eHmUv3ydp
DeO9ccJPbRWRSvlomRpaF3j/HuZdpoLGcQOtVuC06W4FfCORThseb85mRfIT
NU3pIzf3MV7TPRhl+D8LHOOluSeXBo69iiDTwgVL3nLTTHB4DaPkyZ3asz6G
zZX5n0txb5uBvGSX7s3qvZU14OSBTBSjSygZtTH2wTBF2HnKSOfAMQoZ+muh
IpgqdqJGO4Wb+7s5TrSVX5VOmInx1g3nYISl1UKEChycjAYjovNCa+4a5xS7
UnsT1HgLKv/KpQHowjGgbxBfNTPAFuNjfOQKKWH3tkhu+98GKJaPPx4SjJxm
M/lewDEP4V2gYYLynaa7aM4sQiyhVnu15T7Trg8OwFaz7JKSV/NjY61qNavw
5Zker+B+oBeqk7yJAYS0lPlnWlu1S3tId1cnyPEtGlVr9FS44ut3xqIMh122
gIxdjdlGZZ3TBs7MHHnu7gAIhnnVgMtvCB4GkuSra91QfMJ9TjtzM6CV+FVj
3UGfbsrNnbUaSOOVL4c8dD9ngG74q+r2Y1AfAkm9BxCzB4ZhdDCbj80hIk0m
FOazAIFOdGr1HM5zg+HVwYBi4Z1eT62mExe7xauLro8KP5ZW7aCbVtsxlRKp
UUYyTM1oHd/5e6pYzELAohrdG9OS0QOeNFMehC/UlxxjrFFxzaAv+ajgNOKf
i02hI8OJochzCHqiYpGlY2lysTGEeIBjVmCRpcEJ81XosGvzpc6JpL1bs16l
35X6oIzw7HNO7qoVXyGpwCY4BbFyv9vvEXKYSyhNaqT2GiBhG1B91jx/teUY
7lFznyQ7wE57reMHCNvNWSU4F1n2ZAfs5uqyDbl45oNOWuDe7mffDN+avA40
QglFAK5Uh2Kbc1eIACX2FsS+gpf8axJ047fzcvDcJEAXD8BT3L/Fu7CuTWOv
PraOHw0epvMHzKfGvOQhckHLXAR+KI0clf+0lBhDABUlBpnaFN6mPC39R6Qj
4uPUFw4BygLsV4hkhsfTM3r40dBNpec8PxVQc23osY0akVtU1eSEOx4sof6X
0YkepnpL7i/qsBvVlPApmJPcutioBNQL6jn+pfKf/A/n/4PPtkoybqYNsPkw
JoStztuCsCRsJkbWSmyPehWyaH7DIimV5vaX5Ys32P+IkgHFe4LIpSE8zbM3
cRdoKOqqTS18AeeXWM2nq/ZJ0S9tBGIfMN+3CVfFrXPPmuZa5yNWdkjS8t5z
Ygk8zG4+OQDc0fsWDBYLGBH8oh1M68tuTsfrGIH7FhPrinC+uRVvyrQ1aDym
ciaZiFV9OIiSGTWQajHMc5j6cb7RdUAyBqH2rsJIQcCTLVO8yLgQ4kIRMXkw
028sHJeDevS0E/+VQTGAuMCLfO5QX2BlBdS4qvTRJxmX4+JZCBzNO+D37SVo
8xueXf48AqGPGVeLewgFB2P47gSGywEINhHCeHySbRUOa4ZH5Ck6pYInqqWz
lo+HlrYx++64+3NK6TRUeNY/oEzUYFEHKnxXxIW3fJTDbfxa8nZcw5W7ned9
EOww+7fsr2JNHk4damQkfgPz2UmQVeFkyRUn6Dl0RLcc/CBqD5+ew4RXIV8w
tLBsdUe/SuBCZxl36ZMDljfdVlD86sjGds9N0Kxzc1CSXttXI7kEXwYFZBzr
g3eIT8LQQ14j4oW2L7pTXfO4Svpx8SHQ/e2ZVeYiob4uV2SJELCC2p+Jv9LO
e+Jv4gXUWfjwyqpApYujk0eWctlXfUiphIJrBfAl6Kk947TRvbHgvada4Pn6
oW1rN2hLC9q6CZ/eqrm+PVIr8TfRTm3pzul9wpEd3eeg5zns8bgQSgJ2uzc5
rphUWy70iEwNGIDVrWNuwvUuVWtMFFBEhuDusxCBtiS0y678ZOyP2qxV7YXQ
FdjChejK5A9UxcyxOOZnJwMiqa/MnHLI/jNoccMeASGIPOX7WSovhnoVIWzZ
etlefr08IH2FP1NUUGuAn3+UHhg9S4xHkzcVMwyacHABJv63svKKkc3FzfEp
LOUM/Npde+dMFxNtjTaaTDm9PPsY6aUe1ZPuhhyc8HM5VDf+ciOyf0Fzuywe
er9CxAeKx+iIqnPDV7jjiEDXMQrKM4+oCtNZ7ZE7qMEmMg5NCRifHqYoDwY5
1zB89GFjb/USXicevO4fxg7AZCvlgNFKpPebRdjA8zLhcslYyoZfN8X/IbLA
lecN4Y0zp3ZdBPw1Z0XfI1SmKhxHPEm/QxZY+2iUnoIYp9m+buTjLNOZCs15
yo5asfC0vDkaH3rtxIAssIP7R832ZY7H6dcanr7vAD+YxBvIwAKbxHRvFZoX
D5fuoCuAZg600fWoYCK70GdTxE2ZPg7kYLXUm3igVa8sAr6x0+O/csaQDt+t
2b6LZqDgnOMEi6PiVSvj8DfWNBZWq42+2hI8DrdrVFMFKgpJi+SnhmAgHIWN
azFFHemFf3DL26Af5KH9s9woAzLwheO+u63twXXSUh8Ist/yf3XjMKQtPMbQ
/8bgAwOf3F0uQLLyrOTaym3s1q0gDgYGzP8KpXnij+l8yOMBQpxhIdE5b2lh
AOORb9yr3BggywvjTTM0youRKp2yhRK6DECvEpE+yGlkSOa2PHZBqjnJLSJV
O/Qgr4ABEjxHFivqI7Qjl9tj2AgCta7U1v9lUShPXePgejzQdw0wsMFIdkNs
AQcvCmPSy3E3ahS2POVBar6tkXt2BuSGPuEvOn3gjMJvAIYPBG0vtniVTnzI
ogL1R3UR7+mp0pNOvr6D30hy6o0n88NyTTdohT2B4IWNiddgC1qM+Y5OPPYb
ZzQivQKrefb+CvzAsG0OxINdl0ZwYEwGIx/NTvVy3m/U+YlqK6+4+gkCWHyM
KGf7geWarh9qbJLFvlb2wypXOsohQLtTf+GpLR9KXhjylEy2DVbkP+ahstdm
xFlTevKWsffOLaIom7Oc8WGsCxr24PZtRdo7xeNylkSye4XkHTCdJ2HFjiS3
E4k6dAYO8JW2hBdbcUO+VkeYjfMJBUogkPYRpFrEc8VYUcci0zMaxO+LKWXH
a1srPMr+kgSk18hRYxxn/TVHDm85yC5CfTMYsOUS1KsybXcsEumO1+uXyGIo
F9mxZ6nUINlwie1RT3wtHiGfbZYIg8L2vL3hELmltjjwWYBIiQhxMsx8y4s4
tOD69MCOebU7uLS1SfQuovo43YtATEMsNqcKLdkYxlQAWqXv8KMFOZD5vW71
lhO78M9+3s8kcataFtTG8ZsA7da34Qu+Bbix2sxnKfamVVaUiYj1UhsbW+2B
l3/NnFTTlsSjs2vJJEL6rzYxkx/l8YCvn8wT0P0SSPqHxMmKA6IxDi55AODu
wYvJhnuo+HXjV0NQqijta7kTSlWKkVzaYGLAj4sXV/XFUSOHTtIl3mxGPwNa
Rg+Bn08ZMFMmH/TIYGj61maC9V4NsAqvr14xYSAOXALexDKFUIrvBT1stroj
5QzFRWrqPGMZOMUnz9bn7i6rYo7CbjGvMLt/ymUIIfx3af9Ge6FaP33M/ReA
5XRoW7NGQu2hU8BfoaAtr4W+ABDYDXiCJAGvbL0/b1iTS0O8e/YG0U0/sz/R
vhvVa9YNLenpI8W2Aq6XCrTQzo+2TV1SPuheSPBsIShILFGnsEOI2N09PlGb
LoFxeAZaLVNVIHm6opep5Zq/bwrHitg52woSwpBoopzyPKeWb086FFHA0yig
byXd2FFWUObJkz098ATiJ0mpIheKpqBhjTeBI+/peWZdXePus2to10caKP4r
C/Bppa1LLHqvIf1PrTBWMOcG9MsmlES/Oi7d+ABcADdrc7ZRyf2dTb72OwQx
sl9ATJTUr+mJnCo5GUY9zo4rFbgYDPEwnRBQUqIMGvfZV9o4ri9N5d7ExCpN
+K5Zhknt3O4AE2IEna2EMyrUB8/I24MHryaTYK1BnVL3G5f+fPDdyHLs6Tq1
2emsN6GvIPLJiRiw6O2to5AUb36DbmlxSGlVa1ep90Zziy+BQo3Ca3VSWNFd
pXoRiV8Xt9uLL74EtVLvzQvgPFT/UKOK/uAV3VaIPboiXsdUiBAIHI3L6lhQ
sHltwsKl4BcLCMZIORC0ZodMYNxTAgftRcZDnShxHdcWYg/twZj4NgD9gbzO
AB4XH7NMQAhIOw9pAv/nD2UlQ3sXPYxyviMm0rnLP13rQwhB7AdQDtF1vLoq
vvIibkTf2wEo6OBp/UNnIrYJuJUpdnHz+yptAxLTqYD66RpGQ6Gk//7vXw1G
z50JvGSTID8pwhrYmI2ZyGfRsl/oh7vpB64rkjVckdJt2kkZt8CyzZ/CES3o
slE15qh1f9bTkfG96dTpLIDV73X96vsxg+cpMtIQIqqzA9LesYmRgXFzLj4w
qJTfV/xe0z0jnuNBBKp4s/o+pDqdMt28dx/AbRBLTdDYtkS01KcJtah01sAX
hiWdm3gXyA9eR2byoujoX6hRI+uWB0iI1XsM0L2t/nrTAMXybs0mZHK/KeSO
p6iWqaQV84N5ZszJHe8hoB52Qokz+1fRHsuo1G7p35umcneOGBIQIKZCLSz9
8Qgw3VLE/nf9eQykUAZjVa34KVur2OnWmKqbGpDAoqFxgWia9xbML5DC/amT
2PRbz/xfp64Ve9rdB2KW06TGi97S3GekFSWLAFqtGr+XipzidW54N26rhba/
nqNM5Az6j2e7nIh0WvCS0crXv/3OuJl0UmL8UpKTsH8JkmwJInt5mwCKmvej
X3emNyC5aTwbztON2MkVKUMyR5aK1bkbRUJXyl7LwKe0B+RFIq8zzpxATV6k
pu3d8BOxuXanNwofPhSZoTI0XrC9IrYxDbdsLPMyUAr+URLtPeDLRVOq44qB
zgJWAgDo2V7Gi7D64/w+qKI69mBBsFK+jAnxWHz0Ei7WSD0LqeW5Ku8iumWL
xm4eWyXTa59N4jkESvVHz3vuvFA1IYi7tCTfavFoqYxnOEXXNoVQ/pe3+CGq
hcQp6qQ1Joa8i3y8q1WaRBnJfPRNMTWNeUQq/DVtY0zyxBhCv1+HQX5g1Iqc
esObLkIvsQtntVtSyJhzQSt96FYUfeqEjC1mOH/Qsej4voyandVQimeH1Suu
iRuvzHzsGvUOfbt+HuI6+Bfn9uiyuJQwlciYnxNRy/9fyA9FUDLY//jPtuSt
LvcPhySZX7oe1iQiRrnb+ereItE8vgBXBiEvrhvOigjgglbD+tMU9xbbxBE3
6Bjuh2+vLY89uD3tt5DRODUvOu7tz5xXoVOSe5RSmlBAdBzcx4Z3jK/hlbT5
8TaJDD6sZOMqRlQdTiGExTR15mFIzMYxdR8g7KwD4jkjFG0tCrunnLDYIE14
ttl7mJw5w3KYJy6b2D26ybdcJGB4pk+oUbE3IAOLB5/luhelUvQY+mK2DoRC
AQeCV1ny7BLI8/m5TiUmcv0czbPRafAlQguJ7OQQ8I4w2X8ONlhcap85wpKL
FjbzX1BZNhU18GibyzChMABBjiiIVK0WZkFkYjfhMhzXyDcxSFIE+W1COFpy
Fmla+TLa5y+vnp95lNHifNFeUB0edFwa76gSi8ddSi/pvB51i6h61xFKs8J6
lF6S6OKs1ZGjpHW7scIxdgDZnWFsNqanQx9W71yT9FmSjUOLnw6+xxzPUBdo
GJDZ8zpHYxDGsJkGKYtwjzDubSczeOfX8gulhOcW3ew345mgw/J3xEZFXjSs
Zl11UvoGHb0V+7B/aV46hdXLcW+D+cTmqDH98bLgpcrGYKfu2S8ZLZwgMf/+
BFMsWBhJbe1Pru/E6vW6fIGL9E4YtxFovd8xbiVt4eJnHb5tGOwucODfL2Tb
rAFjwTgGlTq22GIBg86b/1ODhdRSjvXxObhXzA7/4Pnoh38rSKXVtWQ8yzC6
2Klxtxe/gUH5gz7bqxxNdqloo9xFLAWzaz06frqmP7KgcZYdGmNRtz+Xmtr4
R8FGh3S2i2gx0/CakF5c/soT+wFhL/iKJcCOkYxbaRjxnP3Q4ra/0i/qjhhB
FvE7Ng7/e9Dq7K9NvYjOvEtAU9SGdanHvvlGsCZhznKP+aUnb30Hj7X3xwfH
Rog7xdojEwtBoVCl8nFQD0ZqhhJIHyYizb0tkTQjPISY2AsEL0FINtvNitOl
H2HMLRjMKrL+6i3Dlchngpr+pwj+PJ9RjE30gg3TDFiEDOhPdhmcn+v3IFLF
7PLVuUT3cBe1dfv3o6onbRZHOUq4Dr+cjjO1exkhGchlMYhGq07B0SDSAgy0
q4+2hcZNhTUyGrEJYXpA9QBAtg89oyl4mvNUykRiN8qlN7jL4jfW35Ar0pxJ
V3pC40jm7qo4zjUmOR30b7Kf/JCGQYB5eW1gEde2LFqfCMv4g/1WoCqxMauA
sWU+r6GKl6VX1zEV0+UFkGiuydX+9HX2r2FOoDifDjjJ9a8PE+Ljc1rtp+g8
WitiZJAV3ry2gjA7jgqvN9lq/7xLSUyhH4GKUtLh5oBoWKAfZT3S2rS6I8yd
MPzUPxC23zRL9V7wpis7cimxFOw7dZzIFOdH+HDvMnVDiS8v2Vhp2Vo9XSDU
OP/1op+gR4i/Zpa6fdGOBBep7z6ctJlaOqpHcjKxcZcIbmEU2MH1o4YKj0tI
c+Keo3VzfM+CFVzdF02AHJT9LV3lNoFkc59sYKBmlDFBCNl3UqL0fVutfxw5
rnSXZCFa4K/T5fKWdlyOXJNH0SOyzBgmutAGhBsuLnwIDlMEL/R2SqjaB9Pe
K9SCqJb2hYJi44fxmWQIxKHo1c5UngdI1uCAx8Iknq0lPuF6zsAn29eLlks+
FX6E3WrrOv6jQmLGoQRSwmn2y4gGgA2C7iaUKS9m6CPVUuRDdYlk49P9vmvX
nVsSA+cWS8W+ap9m+5++589XCW5+e7kt/tIfw9pqke7b8pPsIvrNVvPWnziI
dAjyyOx5FR3qHxue/PuWitMTQBdjwpm3+9N1NXdPScWNF6FBxGt/ZyybwMUm
ZXhnVLbAMhtJ/nBabP4mflOzup+2th1Mc8tYlNv7aHfMcnvdZa6T858gpR1L
jNMcPSFWI65v3pELNIGIKSkl5oG8J55ohslQdOnRpwc0TvAYNtOZICeciTJ0
1cr5+Y7H0jnIkjt5TvnxxKA7pAPIOcNSpJezGqgdEnh9vBAZhEmxr7QiykHL
IaRX1BbjJNnU0pfALT3iVXSsIEmoLWEY8id/MM2G6K6NWQm7Q1+8FPJosyiF
DOkzHTuERneim0vqD1/XPIPtiDMc4gEKjIxjyQsfxWRb8GiDeW+KY6lVtkTl
cXXAu9VjbzR2rvSVxbtY3F4kDWUj9mU2pq1IvJjxVLLi9tX6qTPKCfa+OIKY
ISFDAFzCX3KiHNfgDeOhoIqn0v9au0Ow2GH5xAiarYEt06RckSx0b20xZWf2
cDVoTWaI07tOnWYTMdZWZS7F8iN6setyMrqtXncAgTTcSHW95O4AO/pca4gx
2jANXd9XbUQjuEKDTgenisXgpuh5Gwg54HpLV/WMDCM6g/28WN1W8yWAPwcP
g5Vt/HyBFFFYfIcT5qoBoiffb9n6uSO7efDHlsnA1SdbjWxeohWorQqWja6r
MOW2sxSvdBAx+dkWijKQFvziVwNKsOJL1rPn+Pc51fYJq2o+MJp22qC/pbH6
iYwa9YprLdjcpDvK2ADngOYmC+pifKFlPYmRId9qdJua+1TsUvAZ+0HTaAll
5LFw6Sk8u8yuJy8GIjdaNIAZUMRO+InErq4WuvFV+Avn7vAwjLu77Tk05kIb
bJVDqZ6gdqHPhK4zfjz5c0Ii8PCo+jiQisBqmMaVxr9UhnGWck9Nju6AhDVN
xcJ7pqHR+aiOSwEVKFrD/WU5hIDVJX39KadeDwhDe+YJvptzFQo6kIjK7FwS
ZomypbR5LXUKA44pUxU/V6YxzNOMIp/SNPJMzUbtFoQUZ0ZCL3ZXb8PFFGYP
hEGZkSSqEzh7M+IUcWaP9d72gkPF3jHJxOduv5MYoe5wh6UwSEBRt+XpLUTU
fkcw7KBEIoDxSz2b27HvgV3fjMIxnvuSm53pNV8SDtIWvQdKeTy5Rr1/cxji
2OiGvpHB4J6wj8Eg0JVsOERH+j5hMKoNalalbZ/dr37V0xN+F2p2IoXQIpxt
OQqCwIGOKbF5L2cmLB0hkhLl7OZkoPw3YxRdT6d2Jj48DNDjT+1lRD1P8I0M
U+HB7br4RbmzRM8y2+Hj10am/C88FJQgvsRSahtoijA0pTpFG/Riia6BJf/2
TqmcCq2bCAdXuRwHRWcSKsqxPrUbp3DTbV2RZE2WrpkBOoqA0I6aErBaMpyB
rWYgSYDHYM03DJVXOfaLWLNK/P0cJrG13mekPZTkHvLLdvVaT/zjpOUOtj55
fQXKhQuOrOLN8zkjEy1Od0zKTTfpVfwuAox3H5QlBwV5vdjQaUUMOLksdOYp
Pew496ndzYpnFkxOFH4/qvIwzklG/ZDmcrN9tqFnVsPei+38Dla1F/+zghkg
K7mvpmoUSa9FssF65FwdD0PRgKusB0RwJBda+gHD+0gOcszOmBiq4uf4JBer
B6e8FaaDFo5lsdyZ7gIBbLla6TA2nRSP9PjlouRa2IYVIveeVtVBG4IlYHBT
7jk87/dixCDPlktDerguZpmQQ2bOCg6cpcavpquFIDMO5y4Q+WElgQfnGN4G
WV2qBdlZ9RZmD3jHxMJBXky7Fax+iwca0jr/H8f0RTo7VgTnHV+SIp3yV3Gi
vFisgJtcnsS63aKJ1aMZkySxH5HIc8a8VOVQt1IHWbRSmtWIrrHtgdewG0Vp
7+bTxRImRbA9r//bpeWXJ9sQZF6lJYX/y0K3X40tABtgp++kvS+is8RH5pWF
qruQ4jeBcSvgobxEh0G5dDROoHKDkDL61u1Nq/wjRBE4DV+Mbr8Ly1D2FWlE
07L3DcadQ5d9Z+HjgK+wDGgMovjJCw+sTGYHEkK5lGpfY9JgviE06+WPWMV9
2VEl9Qj8yWxmQE5BK7I7dtAb7y4Hm2GVWNDDsJUjYIGdSoSMFw31s9MLupPr
exW8zAdQDP0jxwAa6wnckHzi+3hErd+Lbesqi0OLWStwvyZVbuEFruSPNvGS
VCdeblNutgwNPFu+u295OS5ou/bx9cF/EzrKxw2BOdk9lIKVDF6i05FhSYIV
Y7IYjltcx99Cp4eGM9na8SeqkM05mEz1eNibFMkcWTEE5XO619QjzvyaeetR
hWJaf76rlJofR/JUKoPuNCyt9zykpRxsJN8vQTPFMvS+/+6jQ0cnoD48Wmaq
GaYU5v6fLTcNEdyLcA5hd2Lz1rEYUIMj0UGhyVT2zDO92GN/y/KrXN5eXCa/
zcalNEUuOEosShsE3JdkLheKfORgTjA3o8+k8rg0vjnPXYOMHbZvK/eCYQFh
QDxSJ1GXxYhH7ALIuEKNAuPy0rQ+CLQqWLL54tSOxvt1s1mDD3L+GZkKpFzc
0fzmhV4NShS/aelzyob61fdJSCCxGN+u1Scq2EZnxDaQV0POQnj9RSUCu7+D
UQlDNoWTKv+437x9sS7JrQBrEoPGRP0m+we4hcWQv3qf1cZsthc6PzkKC1bc
19pHLnUo7IaTKLSqJz4U+y4n+ZimXlvPN4wCKu39l0usvPpPhg34yxJdqgoa
T7CAUrBIJbG3n9uq3XwywXC9+XRz9lU9jsA8W4vNid3WIP0DymgT+yLvRnlt
4pnbQyOunbNOek9bJhdWGFg+umCY9MH36vc/ri8BwxjOqFcS1AJYtqs7gFEK
L315TJ3nR7CdiF4mJ313D+qXHctiTEbY+dUGR2YU5S1g9FuX9VVpqruh0XBl
Us5IaIV6M53pOQOf3TXTRzK6aTkOQkyrqctKBTQuKFfMtc7CZVCRnBh5iyvl
+89HELkVzAgPoiePEdRx9MKiD/q3rdP6fEqXHL1Kws16YSjIsMv79c+6MToj
B9p6gGqqJOStBZOq6phyr7Yoiobv/HRO4AL4f7abulAi7rjkCfwZ1oxUVNGi
d562p7vS8cZREdMGn9ork2fYV0yiaeSZ8/vx8UOtdgBOrKhWPpRO4eBZnejr
F7zSMVeiP7/pmyECpFkbGSLPdx33eGvIN1cFHsoKRSKWZ9GICBtg63Mgzvlm
AOQbGxTd2goBlbRcCsdev3VRdCBJ4vZ/chuyeii65EgsJtZCJ/MR6k9uHi2j
FXjSbRefor0d0tRiVyXowpwlmF5WUectvxoZkrimKGrnHW/5CUIfrhY8F2Iq
G1OVW7xl3YWzqL+egTE4HdmqZuDhemNOExzNGG/YgRxkKCX0dHqZX5TkDn/Z
Zmr7Nn40RMZWRR9tBQNJeX/YQ5lIkxNGoCgo6pPrcCI7AOtx1X0qXicNAGDH
FNYHPbjyVrXMNxKjr0BOTd1fRxVELzZgUEKC+0O6vTM4DS7p5k0w6lNTqncz
F8CskY3MQOYhfNMK5BAUdtd4UFz4dcIDhO3xIumw+Smv+U3quEi+ir4QspHc
3BAVeNCrFeD91KmUGImYLJ2Ks4mp4qe/loxkQwKQ1iO2EjVGuD6kUXV5So4y
/re0w5HE/9ePhb4hDPrWDwyd+BTZBHRWsA/aAY7cvS+5QsezO7BYtjBj0B1f
1wyFJSmBc3SLWsVy2gsy80iezk48lZBuH0tMoKIldfpDH3rOKAJtIjr69A03
AULXPyBRInPoBcyWC9zGSvSGalqmfgb//FXWIMaVZcA2uLGg2jdbjGN1ms8v
Xh8QEkGK8ut3SGhJbRujYcZjJ2aVjbXSQKTmC1L0xZs3n7YZeUE/JGtu85T+
aBTU9cONcXFY9kHX1bVjJgmzI6sr/rWmjK9jRhCJBKTWAJokUCa6J+03go3l
MCHh7lGbPRVEm5fT0vh9t4OL8p3MRigjY8maE06rtdEhV+/cndqbsGTKPM8l
2rBn825qtmRceheGLtfCIAGfKpPb/ZMn056qPnoSSR7cAVKgtLF9zmLjacok
wEFfz1M+QD6Kn2k21IZnd6aXkNJnOdeWH4miq1orl5tBWHZpq/J8tcaD2cjT
4X+92/NmQJa51jtwq3dAFQo1sj2qnt3zoP9nnT6mReWSq8+PLA/MFTk4EU4N
8yaR/FjGU/g3G+KyT/FVoYxcgbsOmxPEXyG4nyDHtzKfasc47VflW0Zgfh+d
+mpSgIdyGLvXfsjAj9xPUqFybMwsvyMWgriPADuFDmyNtFH6SPbgUAdhyf/j
ePSqptteBoWVgqfZEULYc9xLNDhoc279z/8APed8M5kbqh7W7tCfGgKWrtie
+V7w3WV8TFlEzqNKrug/TzoYWCL20dqtq8H5tuRUQ89hzqxRXmHh8mbwge4w
DfnBn8UzrDsnYdLsAid+YlmT8Y41/k6Z3xo6PlJDa2ngaN2Yqc2GvUhJPylD
DIPeqHY6xR8vN7p+tf4nruspNgtHCoXi1LHLQGrHZfWIUG34DEYpxxHJEJ7L
QkTDcwA2MvZHkVMQQOF4kEbrAEfSlEb0Kr2c4IrVh08yQiERxIXQY5zRmFsR
g+4la6/TzxDW1e6PN2S/Pfq/gt82fGhCoVV3x3DOGwi3ECXVC2CVJskjV9PR
GNMsyRHI5f1PYACdYbONYm5tL/P0/rVuCdV0e6emGe6D720VKW7zuME1prl7
Z0PRzvUs7Oqqq62NZE50Udd3gVftmby7rNZd5Q3K7s/sLNGvXVEn0ii+L0WP
2fXJmqmwuTQul+hUQy8Aa+Y6r1JYkDA9XQIgn9bkLs/C1YVa4gK/xBX9kPvx
oC2htD3rCpZ0jKVK31dSYfnSqvPc3uV0OfPZC6OC7TFzQDG2pBJb7+eEs6MY
pQigOmwc55Z3upUl8TXHK33lJ5PMHzHVDjUvP8i0vu96UN5a6Lh4VBrNZqnx
he5V4Wlq7ocXvkC5fDVcuc1ZLBTve4RrWnvunVBu79NfQZk/Y1EtI0fCAYMo
mKQgPDphaj1/JsfGeqFz22cHixjSf9ilSnv2O3GwkcnH0zMOlM/3mtuhWXg1
rQ9Jyc178f5tDBhA0e+WjTuAmY92mx/x9Ol5R07T8qk7BB9rUGf9cIn5ODdj
SsGbwB6Ql+7UMV0/qjxVKZYS/Dn3i1JcY+ua8LiQuJAXl3anNryeL70xPOaY
Wt7ETh1GR3XrVJD5snQhYDzNHUsdvZ/wbYWxDjLTVYQD9tsAtLjVC7K+2UYf
n3YVSg9Vf6nzkscsaasPowQ1UAYfjhaNepJFoz5iqw7bIZkQFYI/gPCIVOFy
Hd32JR9eAtB/TzLRpzdori3hvBwS9slKDfsAroGUgO40HzZ8uQFQAhrAi1Ez
j9l+5vNLw/ztZAp+Chr+QN8FxsTztGeaDmHGj+jSZfJHkwq5JdPNortrIzPw
6gSx/QSjvjV0U4GT4Ew/subOpRNzDJi7a6EzYf11GulaqUWJBgr0/G4iHafd
n94J3MdIrTphGzE/SjgyqjHNAgqvinN6SKzRy545CyfV4fTfuaUCTaGQXf/f
+bAh65I6trzvKQ/2F1qsTtXidoVo2mA4sxEF9aFEKtBqY51Yx6yp8CjyX6/l
g42yd2A8UCAMNFzA3l+uVdvHpp4rvohTb1JDYVAYW1S+GMODRJv6FSMyHFcm
UIzdqun04ez4QP6XG3WxxPT1THohawxst0iwe9dJaG3cEbRsJKz3d+jLlv0L
0C2tCeIFpGtDkmUcE9P16ZURmaULfWisha8B0I/ZZpPav2c/uIz4/ZaENn4J
w/F22M9CZhkZd/edLMzR6QdCnxVPjPf+WmHSyMO5J+3JFTv5lAl+Om4q40kY
NTzJ8M0Z42RovvX+zjqYRiG//TE9LiUV8XPAlNEmtAeCd9StB6P3GCOTvbFJ
iMQjXeaH0Ds0sSGxAWivTR/esw1exJJPA0cPq8v9FPP5pc93tMzW1sqrL15g
NZz2K2UDSS3ytg8VjyruH2wjXCBpN7ovErxo9K3ElWsc1VZDk0evKuOfDvtB
4JN+YouvttN2qJC5NH12AlSe2E56cDxsajtkoF+qfl9n3lRAxUl/hb1Y39sT
u3K1GSdL14iWfxIpez3GpEj7hnIG2E+Aq/50H1U3oJJw1tWsR0S00AI73Hl+
YFVWO4VX/bhV05i4zhO89GWNovRP7F/q7dYZuTvVDZ9qgp/qwy+vfJAPkYWZ
dT1vgoBPKtUAbE2NWDPYwgNLFFqJNoTnfRHHWcMDb7FhuZ6txOSRWloTx/n7
fqZLMp38JbM+YIHQiB1H5QwCWS72LHGRS5TL0AniTaZra97SSaAHOh6v4orx
UpoU5zK6C7ORkPZjm70K5CZ8j52Z9qyUqnbMlcMw95u3ADA9YwLzPlmVmxUd
dKPSZu1NDK1Bpn5OMAgGnLxzew6ntmkBKASZ0i1XDyWeB7S5QfAYN/z3avXp
N//FjmKzpNsjjPq5qLMKgPyr7m8c/Kn65ybIU42NAuoPtkt13mx+uQFnfWOK
KyP/2A4hvHALVXU8RU9mXp5z9zaTcNitpN3mEwRUnK0LoO/6mC+W8mv4sQJB
OoKFa+L6a0n3L61uA0o42zkzagtfo8J2L5qxEjkD7u7LX5BlA0wcob72VtER
pexrbI4sWH+fgUsHkmKcFliMVZCu63n8r+cuQI/FXlieoOebJpbHaE7d1NSi
5vkEIGBNtJPPKnTwpkROz5ptPQJszSM7sc0sfj32C7Zal2C5s0ub8/ZMGE3k
uqboPlVW7mfcoUWtAve8UpDxqGCfOTgakcHyRuWz7TmxapXjfmnO3w7KinNQ
vUwgpK4sQZe7VKkoNPhzZfq65YaQ6mj1ImtLMYAoGCdF7d51JVkU6O7hBSFQ
7q1IUsJEqYAq1/PZRzxwebxann1pZe4iur7/2KLAQnKWkBzPIABvwW8nN7zR
GZWC7AzdEZ38eSgttpGKWW2LWdg3+cwSBpqLD2Esj05k0Zes0L4ry5nLnaXE
yCoWE9XIMukTp00nkVFn9WQbLdXUIFYwqMflgAZGxw7XKaZpReO5TAlfhqSm
WkCOYfnPCQRY/olQ/tYQAV1O1Cc74TSVBPW7ezPnYMMkqAE4tSzkKbYgpzFW
DiXz1RNU6oOhnQhtS/pMCbUQIiRHQfNjBC8ghsNBExrMzK9qc4aJWMERbBij
ZfvnS23paX1fzq0EQc8n6+E7bEc2VzWptrYrMB/ERbH2PE7kPXS7dAIV+8A8
px8icTplMwnWw38ty1xOUNVdMxhojA4LiwoPlrjpS1TyaQuIlSP/fFHo5SEH
zu1vVI+eS3XG51Kohg3zK/dCQ/sIE4GohGpOj24GxD6sPhz9IntoCE1VXNBB
QhuqFDVBaKzYwZ1HvDrvTxnM+SsqTuXe4WIBnCI3vT7/fNzq0LJFO7dRkFBz
cGaSsRtUYESWlbmlPgwqC5gv8xAlyh5Umhxykoy/LGNY8Li5+PRavmrkvUt8
BXfBFhHvKGzFaNenc4cO5J7Zd7LCNsnuAZ9ffBJ5wKokVc8f8mfW7Ec3Md95
26oFiU8oHw+DbAOBGKLJIgtfUqqmds/UIMyGEAvJCUMVTbTBwJjyZkOp9bV7
ZOkHpameXdmpO+Rd/hlWc9M01biruEPxRDIsAiP8eZkD3nudo+ijtbSUhnQ7
mQuOTtOXdRFVQ4PzfVH4rDIPY4nTwfdV/qC7xppn6KmFN+5WJq6bOfHkd4R0
TAaIOEOeQoLlFuPZV0RCWqe6smk2N6eNf435HBZLoxgnvfS19aTSk0s8Afbg
PltsQctSM3W3JQIIan8e7n4OAM8tdIB/OiC2Y7FfS6eUO5AcKaO/lSB9pW50
BdVY1dxeGRmFmHuQUMq9gib+5nZuxK438viKwcTENPr1IHpBy73AgZsw+D7G
GMQBp9Zw+a0UkFUJv5y7OrA5PL5RkFK77amOxzIn67Fywq+XMVjeqGkZtZcr
6Xow3QxRvMn0kC2Enx3LKy8J43TrAos1ybT1kx/VrPJy+kauKbOSNhKKk/q7
BaMU3UUGsGkuNQMbrBnI1LuXVa5yjYIZDwkP9tR3GI7kcivL6e7aZV+VY07h
xEqkkj3hAg7lbuS6BpbrVd1bmzmT9OhJ36o9qvHnCdD6kkgASVQ35oo2/gW7
IQIx4z+5lLfoiBXZRll1FyKvOtq+eHJnn9OtLwQ6fu9gnR5DqzN3O7YKgJRH
EWLjoT0DHlgAXcrJU08AmH9flOBFt1JuMJxzt+OdmgZLvUZGxTyKFq1kaILa
uYQTZRMsaeD4xl2RenzxVA+skKuF6HcbWsRnPHK7bMWgRfstYNNJxVmB/VvR
2IytegZ66omBeEP3AM5NQgI0gE9Nr4XM3XRwq2ciqPbX+4wFAjACkYQE+FX3
rUrcWuaUEhn13gfdLFeedruGMlG4uz7wAWfBP8UL4/bu7qy5nDW/G/CYlwrG
2pC7p2gMagfE7Od2JMVTUGW78ImwBnHC0GJNbCp0FtwxzFbAEWgpjq2Qgy45
0GbW9w3hP1qEtpNTOa9uLK9G5cH9zP93Y4gtQb5/Kprb1FyulNtyR6tJJ6Xf
0mp34s/B6fDThGxm9gnSaIf+IbXxULx+eykMClL573zFWqkuppGk/F+p9eHQ
FqNdxvHnjZ5fhZMOVE3gttorfpXTz6m7YtYf2dhbOU/BTf/L//2tPemltNnh
EG2xHnoYz8rgvTInxLQ1s88e6zrhiJVMIPRvKjgDhEINn3kG1h1ZkQjlRKqN
eBtAmL1U6PiaSKu4PDPMO2zjvG4vorwGCuqsW7W0eltnuB3SpFAwnCQVJ8Qv
FySDoUR79Fl1SSdzNsYfMDy3p8FV9CX64v3Sy4zQnRi6Gx3R1W9Uj8WRwmoU
V1LHVgnKkvgpMoMV7ZvVl0MulKCT/47KXi+uewjsAAC5ifvXz5NX/6eUr/79
3yzz8sQnJSqQbj/hJEnTtLVW4vCLsNTbEB164horGc3u6uYTw40aU0UjPMul
efOB3/nVq9U4QAkFaHizssqzh1EZ4FKmhVREsfNIjbHA2fpZlqaqBKUirF8p
w8vVyduJL29YTSSA+unx/xvGAUajd3cuxtSOpRjPHVSbWofhT8YM5Mynzs0a
gJfs35WHAW4pMFY9harWrS/GqCbDWEtvNz0GiNWNNRcX8bCJtP/CH+VkyMsu
+5jXkmuAmuHNCvYL+TVXi9IxDeS7+j6QIzKvmcua/skqY+DOejnjPZemlxeg
rg0DAKsSkpd8Tt4j7vtGByw6DtvaFtqWzlkSDZg19oihxT+YHYM66OzqwdD2
VdAma2PkD7zDAN9uMLVZ0z/ekeQXY1JYXh9lPBQs9Pi0Qdq7Y/DMiFQfONxs
epteYg3RirTZj+5jsGBOtUGS18R5qArFZhOufSpb0V8VnPGinnA0kQ8IS5yk
dgB0uOwpTPaw++OwXM88s8IJ8jqntwQSBNVPog7wtthYFidQgBsB04AYuBwD
I7Q6g9J5Mt3nm6QXgnjmRWoe9wGWPJhIILNMWLIut3yigB9Zw6iX47sXrHfQ
vlQF1y4GSK03rh3bOzAg7DdzjlgB0aP3iihyOFrjYUx+LriZG3GY376onzV/
dXyml96z1BkV23ex8PMOGQSYhqQXF1wk3NI4I1nQx9efRct1xkXa8OYUV4Jz
YJYc2clRLOe6tj/vepEu2IFZoiXlndGJODw9fo71KhRwaPV7znNZdIU7Q2Ts
5MY3gaa+BfebtOoPriEyS+zZOinkJYApIDwEuyjpTEt4uRoh5LDn2IOg1nLU
LH+AImGNRE3SARMQPrdDTywueZLKMKRoiO/wNqqkJMRDz9JVf8TUjy+cLiMm
rw/ac9TmtgY+4aebBGLs9BIimuqF1mYZ2cunJY58Xd0646hj6wwy1DOS7NDA
tl56qH56m3Jjh5xNsva1C1xLelruzvLmHr3AR2ZN27p+0gciLnQ1JuZ7xbUP
3VJrn3cJzig5uADAf2fcBjgaABGuWxOIrNBPChVwpsMWPu2OSLh5Gf0D/pFW
eBQQZ20EdC/o2ZibZ5Lc3jx6geVESzKu/GwMNAACMFVdJh+fv9sTEGEX0jQI
8qlvP352bZnQ2u6V3UPmXJLG8fOWoCsZKOTKWd+oInejc2qpVeIjEmqhFXXz
80BEYKpoFGn7AOFDOCx0tLBzuBYY2d2gz93uMgm/Mp80pUMUAxduDWFIaSn2
GFtb0c8aCOlviEwkUcMCm68IfdbxdDoJYkuu6nenKnmN+l6UwhlI3S0PJn72
VsnpJCsng/L51yJ+YlSQi0uDQoNq/E77NM1BQwROi+NQ5HlCvN+bWwl3ZPQH
miJld61Vns0Rge7StRu0lz3RoLoObNPjRqIKvEoxuMSjjM30sfG+Rx6iDD1M
04EiJBxFjTPsDIEG4FDWXonR5nJ12thwEBT+MFPZqbZGiyLl6HgCjpvbIvv9
oiKrVDuA+71WvD98EYlI7p0VXDYUtGEpqlbv7MQo16q0YkLeEuxYkIV7NGwb
niUq5yer2uy1suJPAvDcF4NREOpfX+PiWJjjn2Gtjk6ureNMFSKpYvyC++sZ
wt2g1DgTtIq57BnZs4lI97qjSXHkZtBjfofs/6OkZdjI1xh2Rf8wXjqSuNxn
rVcBFlu4Dx1twTaIDRv4NaHo8ElYRMP/b8ShPb38DIaCG6AUuGBbzHfoi+dD
PsikWiXfwk2RdUZ5q3zasLOKtFI+1yVh36AEMdQxB86ewKYFx2POOw6RVUdS
Vyad9FRxPK+j7W8/8WARVVQRK1NqtXbjAWka9PE9ccRq6lPBq3JRMgaNhlqT
H1k38l9sJeYpvTDEvJtCBycFsUFv1E/tBtlL+fG+U8SKcQ3X2Z2D+MhFoEn1
OpbpaKUn8vvl7qsDjdWV5KAAFP0WRwj/RMzm9od/gssH+6YydFkpt7ejdotT
+9ni2OkvAn+20P/iuZkUldQor2T8DQbPBCv1I9NzoRbX5hUCzxohTOJ6EAxR
z0NZsPoOL7/1QWYYf48ZEIdtYBBvevK6RYnVeab3HLGKKSmCfvnArkPPysms
PoUk4Z+eoNumBRJRCpIBz3f6U5SOadELRnQu2B87XFHU1GWo+GSeKVLj+8vZ
EvWjbc6n2FnlvC7vbC9R3NdjZA2JYMe8LO5u5H939Z07Xub7X+tpgY54QwVd
Yy2nfTNXJvDb1xT+TGNbG7Zzkg7qurqm1lxgxy/I5hZmPr1FMXEhyyo4+Nqr
3nEuCXPb8X5Xcs8U9pejt2W6PemCxqmzsmTG1AH285FaUX6YDwYyLyWQO5xF
PeMpydNlV6yU1kKJzZvEBZWDYDcLOc91YFhJ0u6AyrJd65ncbrx74aoJxnC+
iHSc6x++r4elOAPEqUSRTK3POnqrXVq2gI1VPcAstO3SJjmyqakYyXHkgVcR
siH39AV54TbSVfbYW3HM1s9nO1MsGWeHin/Ph2t5V92ysOQ1o6Ug+1bYesYe
lYk2A4OvJ1XL20amfm5sa94npmrLClTmo1+NYh2NjnCyFtlbVJz4F8rvrJsB
viHF2B7R2fA/gM1WGz3i4dMPEnUC1/oCueJuXsJNxuKIsSpOpHIdEsPMVEuv
zN4ojo0vVcvLAD3Ix43AJzzwoxSf7283z2JIMFaCF4Z9p2+JPpEdeuO/lob3
Icnjx7g1oYi8RzHoTmADXhi47811zH3yq/35A5QO5mwh1laO8rtR6Otk3MEY
ucoqFECbyJGI0xjt6DhfC8iqIFMGcBA+Tst+QiPFTxLGsLVyAnj3fbMxEuBU
j/7+NsleDS1sriAZGNOqJtxFh5PVuiLkMfqnzRWniDC2LfnOuCrO9qEk2As4
2r4OVV9R5Vz04kfTfEjUFaef3pJXSNeGVWwN0QgfQ+3FnLaLW/W1zphd6oSz
/YHFE62LvXuBCleJ2FR2HxvDgxeGsMO5d97zqfpsjqK73WU6MU25l3UZRmP/
lVTJB5PHoqevB8v9QTZ03tbjFKHWGpYvYslsS2oPIHJk94r9vjUThGAaXNJo
j5lFSr/opILRMkUXFUTTVrVwzggXcbRIRW+006qfkmZ+LpWfq1ddoJhXuZvB
qiwbemgrtqi/dIrXg80vwZRa0YlWbgR5EAc+8MThg+GPaFNw1AaR5gY/dsy+
WfTmKpBZYPJCSbYL+ZN0fxM8B2/fkzv9sNxpwiks/hVXzj9ZBW1GfmDp+XX5
Jpg+t4tuU0ToXxwWkNcxnPt66d8ykFClhx4vRIh8uvX5d1JVH1WhciI7wzp4
tDD4gnPg61riyvO3vufK34sBcL/UR3LyIhgCSz3+qmbjCE+fc1uqOc2ZSZO8
141FEXUXnDgo7BtL50aIEfx35nNPiCAA1gCYNIesJpVwMulY9fX+341CdUx/
Ae530ob9miMMyKbKDZJzVAN+3XKv9MuXHEpIucdUSzK1TgS55JihKOr72s8I
ajzzsnXfLdZcR1mCfwU2AgfQjJda3ubV1WzJhKWzKbfXjK85//Z4/pBhJX7t
t6RhvQwaXOrPxBFFnAGB3E67LqETinvUHsLbGTggtk5fSGmieliqf+w07/xr
lLYnvW4MfPLvt2RAwx00cgaaZBgphtpoDsIk74r17uAEiH8TGQmTR1h3cBS1
w//RXilESq7fqAUCcaIECbCs0Hmsv79j8rjt0tCOnpsPkXnwO1HdrYt+dz1U
mC6Qwgc54YuXDDOm8tJwXuVZ0cgscyeztdRvRDRuc+ld8Eqzfpoy5ISnMDY7
3XI/dQBNsJEDYZEBBR9CoWTSFwkuKm/2cYX2IyBcWoNhBPD3spZ5Ge3TzqLF
q+T7JdFds0FPDi8nzb4gA2m0UShBfUSOfxsombo8ctgcXsGSPN4MlvlMKGuD
cOCG+I5Pd5VS65O3hMoVkcGIL0cxlhxgp1MatDp7kurwGmxV1sRmV8ejIyAi
L6G2uZhT8BOEIm8WRbk6PvwCNUnucRk+Ii02jFUpDIjqR+gxausiXwZ2WjEu
CKBRUBq0lqntdC5OD3Wsr4ErC9qLhbjAg2vOynnDJs5H2YAucKVysz08Nm65
EZOAb6UijATAAPZahjTgxMQp+7R+wpcKJG/qtXjUc9L2UvnrHwpDxPtjk9RE
Z2HJ5A+bCSnA2nTZ7LAxuwQoKc1crwC78Vg+oRwjdsFjF1vQtXO0KVsJYlAh
6Do4+yXlWRfoVwEZL6RLZidollSwF2TIpNPd6tnAoiNcitfszmEDAOSOmYnk
djeRdgxIWKtuSjQV4xPw8aPMj6fqXZo7CQiXcT1DLs+WQLcCNW27VEyAvDrj
IkJNNkQlXB/gIZ1Lmjxw0pdMTBX1esy+IjHLt4HclboiW/0cRXUj9SDs5YGk
njJL/XBkAISqTunaovcG980pWMxdGLH3ZA0j7TbvTWnPR0pU8p6FkJbTnufP
+YMPksz+rxrnxhlMXdmDCVAiYK9NYEqy9RIq/bErc7AtwWiSxctlHuEo6+A2
coNbanU7E6Wpfogzriss7KaZKrLqN9aKecnlqfe52I88qnxo54oIJvYBgoKb
rKMBbNAbj7LWnPwhUeYv76dOjRrvhpFVrF3q0ReukuxirPpqu5oanldVwLqX
CL8s0Lsfbc2a2xfNLlVzghHdBt0QNxOas0qUjwGLZUnSQLFF70/VOmp+l9ZV
djjz0Ixmsz6scC+U9cKEFSpavq0tV6HDuhQu7hBIIvfpdaXA+B+9zxSChMSO
pEvY4gBCudGK0rX72jgFsryx08B7erQMJerelVB16sJnPzg9VR0d7l2pcrTO
KE+GrUzZLcVzXtNdG2gg+sEqJ8ingUEJVSGZHiVqRJCciCbN/7/4ExNUl4GN
lmdlDhyOk4nj3eHYmblAu9iyj+UjCbr7nam0fbH/kPS+xY0nBsCjRmWUS/sZ
4hX0XuEDLIj+pEklIAg7sQvjgiQy9r/WL+XxFD8vzKnFd+OLCqoDlWIhpxp/
xH5VMrcHmW+nv3ljt8Rhzn3YduRRmMgsszUqLJl/ie3Ymls9C69FhEsLnCjp
GU8NeNVvt9eljpr11DOiUiBquoZiS8+NclGMM25sKu8IP9jgp5jFKZ30/sUL
K4w9G2dx0j0KvypOGGcTiZUKFOLQOfK0ZpQj601YHZKyiwWhz2uPhVLOJvjC
RaNTgx2uHR3shpNj6llV8/a6A9RvY7rQcLUritTghRSya651ix+DwLNLaPfj
D2b2jw5r2dj5ra9+t8DEHVkitdcZT3kuN221+lkWCDVemm/igG2IMU897/ON
KhSJeup/CfIaDvDjBskyqbTy/DUkdsnXSdbFM4XNVPvoUjDoVQjsM1pqMXPe
E7Fnlz7ZiOd6uC3YAlgVVwujXJoAvNXLFA23++op8wRnLGVGge5MEb5zPDH9
lxXY5q0zWwtU2+QbsQ6XDP8qTkfOK1nFIHxY0+y04LdLoy0zVQF9/v4aytPG
XV1GKM9fmUg/XpxHzj1/n1L17fgiWbneWEBjIOqDNljyZhoF86zC3IornCC6
TuiW8f5aDnNVTajCs/oF8N1UKlxhw/oQAvl0+sTRr4lVztNZlN3WO+kyqS3q
tS/0S1ri7rHe6jRjdPKtCRGBZyM0+HoEToJT6sQv+VcXazBgoPYEfdFNMPkI
2d7UxpU5f42V/xboiHF/mZIlKotd6BCmzE2T+G9c1OA/3zec3W63Grk1pldd
Sz2O/7sdMdCEHxvr3JpXq6k3mleAEh99ea6FM2cpC+8wIgb1bZYZUZ5R3AOl
Z452iB74y8CNXQu94qh9yiuGMNc6SiPpG3PvxxY30sM1v3A9rj6L8tv2NbNx
ug0nYq59l4aozU8+hbzGuyKWdhn/PFdePdXrtCO+t+uzayHGNuUaomSkUK0q
MytPqB2hF/pKFRkF2Vwr5/5+km+qcB4jnIAfP8J3FJlJC1T7oNeo7ESXOS+F
kfwTGQLFXnU5fw3smN3Gqkkrfd1Q+xVbZxim8tOuuRLV3AP7KgQI5lhMKhRw
WTJUyN/UdbJeFXeh+Lnk1usRUwV0aUyGTb1PstTnDbkLgG07fgTd/EhmfBnW
YMq8fQkfQaYx1QznE89x3dQtbYEGOmkrac7BoHAYicjmM70KDdYiV4jWRxl5
UR6OU7P3Fvax/1LkT4UyIP6HszVqagG+taSR3Pwmeu82XnDolVhhK6N9EJ6L
7P1ciqRhB3/AkajDuhV8DFkgKxudBL9l7H/OXb3eGGdVIwGHab825Idp6P8P
PjuvISbPbqUJlN50L0JyyORz2wqzSKUIl+YCVt9JEW8jAgbnL4iLGK9JsjPF
tiPusHifbXTZ4DyW8zT11+npFysLtZfgzVe3HBb2eggwxIe2tYM3I2PXP/Ju
ieu6rliQhVZVppRZXEj5YclUT4oZaBlezElOyJPw/oSce9nLw7Ihf4jPkenV
mRWWrcgfWreI5waftfx56jw+CY1KSbMgdkzZC0T3btVlBB56rzwP2c43MKQo
/v4eRyAeNEb4Qzp5D9pHNNSkPaIw13xpJxWhxjrdlpj87om/HA5w+8Dng1r9
DECRXXfgm5PanbFdHf8hUOjaEQGNo6Xp0rH4Mtijw+WnXRw/0s6/D6+1BAJ9
OMWSbPHJDuT+f7ekM1Ezwg7qh4SPgui4XwKqBGmfDOHEquKUsoQ6XDSbukJ8
xP5o96tAvjTXCzM6yMvmFBAA05tuSVHnUxHMOHIiCU2t9idQnATdTTfjnq4Z
uCBU8z0DmJHKkYleCCI3bT/0SVT7Jg6WsT39QlZ0prdZVNpqygOM5aZeNdJ3
Q7AM30MFG+Cs6oftU8vgZkp8fwvjMvDPZQPGmfKs818TlhQyZpxBYEKpmhGr
SqhOziBgXB1ajczVJicE+zA2SlYR4pgdedJQ2RAxh44u64aMlyW8oxHpdpvf
LMYsLT+1fQMJFNI70kylEk+d/ZrR2Zg7fKeNmgrU8MphB3Yqght1LKpxOLn/
DWhtd7CN7oE75sh6Gqgc5QK6fuS1rMEh7xiGr7ldGXsRf2WLaqWMDejCxj8r
Q2r09Pf2x1XMOH7XT3hckcPNyGNVieea5z0lNoVw1jzpITr7kh4HZYsgP1sf
dqhPL6c+u72FK+ArQr2dJhLsBqIdixzhO7QodKroC/1TGz4o6A3Z9Tq5bOtO
C2BvBPyh+UInKIpUlo09YAF5hdDYrxg0QONh+gmaV5X4pu6ZzZjzrKkFshht
oUv26HwPVaATbiMJRtanmxniOjcmpv4+1onyqdKu1cG6fAqwXKbnNI2Gbv8n
3h4vLN9bwtHDzSzVoGUP2Ap093Mwh4Lni0vWAAQMDa8yLAIKUQqZYzzZ2ICM
AZTAVknP6hLJQZkLT2dHkUa3A55WWWVTQfyaEeIS+bPq+j+7GFEVelHBoTVG
sVcq22b1MjJWSHp7+r5B6gHH1AVVw2LhkKoIizjwUH+oxpuXegOhmsmRxCe1
IKggwrHyhMNGHotCcpG4+r+witjhWOPgRtw46erbgQ3p1hllSXaxcvkXWehB
ZN35xHde9BqksQYVRcqth8VeJbpxYEde3qNxHS0rcnugUxkuasYnIyOug0YF
UoHWBX1Dx9U3Hy1Yy02VxPPqVeJbFe9SqqwPJVmcJa/L9UHet1yC1FnPXgq9
SIimbSOvWpYOnOnnTlD3E74MDvYrM/g+FT69bTHx9x4MqFQDEb481CMB3vVW
BoCvHL0aiSTJJs6aJruQhhakJzmhbI06tEyPTr5splC3chCPMV1Ni6ElQYIa
S7oo12YgvVf3odpo5Yi7zfM7rn8PUsYJHQcBuNIJlytEgQM2m5WELGM0+SM5
upKhT6wb0MxNlpZb/29yLcEG1ChX5PXlFlJRZRsjZoUzTNgoIPyFu0GcTdWC
78522Hdj/us1EWKACUeCabldNnDUWYN4YCq/W5FxTBzU3eH2zw4i6IFxfMpU
mczlnlknWvtv6J2pUyWsD5V9YMRSpOGIbjFho9baEiVEQHU072o3ZLjqe/rh
wEbOSLy/KMLoa/K4fUmhH4x42ZHIk1BHlYKkpXc2lxfXkA/VBRAfkjKH9iX5
opyWp9ac67eswkq8sne5019Q2NXgY5gM+z4vCg+oipbBg5bJ72bCgvbS1Ycc
jaAXsr3iD/vDfgnHwGMvo6g7svp6PSH6Qwu7f2sS04BzMNbqmU6OamtiO8IW
cz4yNhGzXh6++CUSvV8vCBVgRE+pri8D398Cv2tChTPFIqCDEj7Q9Vw4UBnN
hOvcOU666t0zzGzcuE3arz/fmgpd3qC1bVVtHW0Gq9qJo9w0zsP1qvNAksnR
uqx+fBTBAEr4PjLnE7aSon6wd1WMj3xoZYuCvKSdjmh4fg92S2m4bQUd79RF
9+IXf1WXv78oXmgPkm7g8qTL6WZ+cdiaYab9kWPLKWHDJDp6diDhwDuo/OkV
EawmLLYK9GwZQTmN0wxdOEb2zzEjVRISOc8falSjaZtbznXa/2b3ZflbxZHL
ZK/l/IV8Ffj82CKtaZCMj+D2OrvuNVQo3dAlpVii0wzShemzsdtZj7689E4Q
QI79I5qlmX77UkOezG91Yp39pkhR7EWj3covibDIdoDDclLtiGU2egVXiukZ
VQlzNpapPptLwIZAf8mUf18kunJhvu776YOQ9s83whRHA0dvCQXTLFyGTv6z
xAkF2MHSW9I6fNRv07ah+5pLRdslgQBOeA6H9UH2yS+fPXtLKX7W8LRqNgVF
ou4+ibW9FOW07CL/yoFpYuWgJ6pMIINnbtG3sdUmFoxeUGVqW0KCuVWIgsNq
nUSi8EbTuVXEsulrMvHqwEORB8Xlz5Kzx/9Fu4cxG4yHjgxQSnZZe904291a
S4NiqPm54eei3HRHweNWUWPBLX0EWLZuDmVgQ0NqKH93taqyHC5kyDi1BH8v
S1MhzZhOfmPhdOKkIXWesHZltFtla1OIPygDG14Qx0yKoKAar7DhPXjEUy2G
1Qx/MPNT+qew+ipU9eGVDPydA7hxOy3nlMbPIJg7NLFf75AyeFFqK9jq542w
fwF3Y6z+gprkyLjohFLTB0hJu6tf9nkdzhKX6vj7TXl4aFCF6t4BIWD7lgM6
mXumLI+arUGE3BbRh0n14k195MoLR0X14SLr4ds4UpZ0hEu3zdAAlu2u3gRF
clMJM0Si5OJsDQtImm88wp0y4oRLge+nl5SoBkv/MtAgWPdjZVd725mL1obI
m8qlZgaJKOqpySeM7WxhYXfQxv3NjLfEjyrwCKPRpDA6pyUEZTa+2YY2kdlr
Y+rt5bA/gjJLzKET5EuibdukNZ1/jitoSbeaqaH6CshF9LwIuwF1HRdi/ixe
iRZqab5s+gFaekvSqRy3lNirGd5Cmj/S5dNYvefieM8JHtlROY3rAEJQqJGB
75ycvO7dYWH87d8DnxLEwyEt2QEAu0qdYCB+o61jxc9/bJ+woptWtN88cT3e
g/tFBDWRA7EerupMMM8PthnhkaNSM8cEY2yvW6ef0oL6tBgqjHKdrIaij4ux
6d/CLwgfa0oRoFIFm0KKsekul0Ql57+jlG5W0EwTlKYjhaNXI3B6BrfsJA2t
s06dLuZ9LALgQ7YzAhnWNIaESZ00lgxXDNnqxbKYfaKHC/kCeAnQzmXM3Azc
F66uofVuK6ZmUq5yEAX/1RiZhCD327kdtvB19fyDBb89+TZ6GrW6KhggzUS/
bTRe1gpceQ5PiPfGcBzSF+iDqT2e6qnppoXo2WKZpJy4uTMG7DKJD98LqEVu
9cpHKBziq6ZUUDTh8mi0DWYXLeexNGaPwzY8kQFTiKJIknL2W5ZYzqoRU21U
DWwS2Tmxi1sHDsxEIqkYBUgObDBw35lJuf+gY23Gqvhlhd3Y38W4CFVz8PDt
GWWsTVXGZJ6iIBOah0P/HJpT5mk4Hmudte75MCSUwfhm8aXtyZACuown5jV8
XFG+GwN1xu/o2Zm5O7y9tqJbMjnnFFkHarKO/gyAi1DBWKS+PNa5xWsQmdQh
S+v4RnvZWeppY7Wm37BXdrW0/3ZYGeqJwvku/lJka+p6pjGi/RXIqTqO0fwJ
JeA2NFxxlRp37TogSWFZ73mWA0Oe1oY0lcJTkml64ZT/o8zUdnBg4jnRfWoa
75q8h/HgzAH4ZBjF8xAYIAADnFZt91tWIU5wF9Z+DC3010E/geL4H2hafZcW
YDx1f5Km4wttmC/npefQHQcob7+ozyMvqHdEX/mBXOMrZ2lvVUBit/4DLS+Y
8376sZEwiR3YbhA/8vd1K2R907ecBtf1+xQNEPRMQGQGlrfEE2E4BgNnMx8/
aqGIpIWEIiah8wzaYZbh7j0KJNxnAXYOd+wg94gyMM8YGhRH+x8oKw/0SwE/
2hC4EjkFjI5y0LByuDuysY2HsqD8zADvsYukB0Fqi6JoABZTTNMW3jb1IxIE
JraeEX/RPTFWtpSAJuQI9dOl0tDWRTksJqWyYYlvdyereUbz3CXSa9yL/47n
LwUGHN7PZxpHoouJ8gRtTGBfNRlfP1nE3sgcmZaSQ1sdVr4esJYhRWhJm6qV
3ekkHG5SUU7fpyglN0OjtFAAwSEnD7Mv4CSMmGFa8FY2I9aNm3dV7rVGqjLa
uzCCTzeSZcv5ZvGRRwJvHL3y5a3XZJOYCovJikWauotMVQJ0R2xXH1RIEmRw
5sDzwmOLpeadWCtXTUrXETV8EaXkO0b40DSKJ2w6axGsB4rQ+ULQN5okwgLt
GOgGazBT5RRqLlxDqsXsfwwq2dpvBlQy9YKYUoCGzr7chCwqbI0BxdypqDC+
j+IWmAwrjQ/L+aeeNe/ia8QfRFIUY3ZmICrOO7AEk0g3S2oOv4fpsOJkDEIH
CdyvXjSYP8UX02g4oayCqDDHlJQhLy8bvTsKf1DLmWS3UXsRd8SIxwF14m0f
rBwDJsDC91HSflBwzN6H26/LofViB+0zBcQ5mQcf4e2QOvtlndIYqkjgd7df
X32qkuWp5tzku2d6K8u5E7QtgQ7VmdIOoE5m3taOYVIHUirG5KCPUQXr3+1E
0C24p/Bd6vYVlZk4QzfsoQleGpTFiwdPW+MgWBnjvRdmyNi9lcKjbaQ7o3Tc
PHl8o+QzcCxQgpY3YrG3+kIU+CeR9iPfHePFOAMef2KpjFpX8SAlzVZNxk4K
tp4JDgiQHvhRmLUrnG0pw+EuPb1DxtV8RkfDiYaNKfoDhZchalUMOSU9RhN1
J5mf93pEplou34V46xwkPqBtrvvNDK83hlvalB9pjcc2y/Bpp4ZXky5/Vv8N
P3m1BzEdTfbnWZcigyZfXbxSFcjtJ0WrXNPoiuno5ROjdsiNuP4cCplODFur
2n0Ol/pt6X0qkOJg6MY+NAVFCVoe7Xh2vmbhAo5e/QC9WuTSBM/CYCCy3VFg
5e+KByg6AO1JhD/gZ1+M1h1dbFd8qaqEWRjlPTIm6r5NIXDzJRD7fQBp2N3k
Z/2P2xoWIevvpzZ3WP7we5XrgIKZUQyFoye5jBjWURNyaSPJvpu4mZvgAflI
Xe0UEcemzvs8JnxnAd1faLAam++XO8+fxvygOlTSC3JmFB2z+OFNQAHspdRM
cfS03MfLl2C6gupOT9sT1Ux5hQXtI11kKjs+QFy/nD+o6Y2RZY4K9wctbEBm
H+2WJYBFEAtGQLYPJr99uTmHrkriu8F03Y/wpC7ohuuqh9d99RC8PE6sJGKd
FYwdXw3L8jf5uMNG3BtxsqIC3OVvRadBL3B95TBGjYcowFr1Qf9AKeJT/Bs4
p3cmD8JZ69sUJt77DZbh7CKGq1r3/ioudpIrwaGPep/DNBMvMJopZxtdJ+Ok
JFZqSwpPOK5d8r605qLkSQxMFDrXbVX4SzxzP5n/eLvypJ+vTa983lsrcmZh
xCjsolAygPoHoLEe828j5vkeHcC5kLYTkLn6+lTt3An63wpH0B1JPEs52sQU
wrzI8Maf7LVuU2QlVu9MO0tsk+8crgQ4AYGMmxd+wT2FEMX6k35lpZv/ZGew
5NWzApXIVThCniwtXausTlr8JC3LExyu2tFYUU7s/flz5BZ4moKVC/zeDaGf
Q+XdjnIch31vt/dLOvEyOGPiXhI4/kxLRYxPUesN6WVMJECP7PROxFOCPBtX
d7i3LqaxQLPEpcYD1VsxTRB/NZ/KFANd6xbyu2Z5PWTMYuwcz+5sP+EJH6rT
HmeqZaGjZK2pdg6J7/q88IkuuLr4+O4K/nzOta2KUnGET3byuLDd8wrG9sT+
eQIWqMbDVMoR7mHOTyiuiPCCHjL+OWI4OxMbZpXsbCTKBMSut9ynGW3Z4fzN
TevQ0Z1DZPvPcagJDFZ+x6ERzFglLPqeY2TxHsk+IN57XCFpnUUYiTPxI/S8
jb18kR4HBu8K44wXOlpScDZ3ZST35PVUpNwvnu+hCamIWEheM+e2gx4ApL7x
bL+jFIKfR6PqSRIbZw050YzFUqiq8wePvP4FiyGpcZGJcFJ4gbnVgMaz/iuN
tB1WC5ItY9dqwyWF1ljmNBYGAdYkYHWXh9UPf6CEyy7y1Q37g+iANJrpzKKc
S5AvLvt24+PsgBVU88Fndi/LVyHpKWZnHwZUykBWdqhPPjLTCEH/4vkosy7u
0iC6NCEhfZmFhgiROilESAyi6gR3Yvk+i/r1bJozxgLOq+ybBGNOf9heJmJE
KJtQQLKEjTIYDJks9Z997S4RMFw0vk5/1bhO+KPWyFDG2gxIYzCFzvo4EV83
hMJZXwWOMJ0pLmnUi+v8FKtnisO7mPEHC8huqeHD4FDauYWKsTw0CxFzpivD
o7KSkhFFI3e0Ps0iAdg4lioElk3qkNuR6PwUfhEluSr+fqXXf4e2JIVCc2n8
27wUYhsWQfKoI5MwN7HnVKgqKSf+dNE+RQ/IlVeMf8e/ewLYKUhtaynHrtXu
r4S/MRNHO/8xoZj2zbVkcvPcPyD2qNq18zBNEd1AlM0/2fhxfNYJ4xA1w9gg
uI+LdzlRSpyoVldwCeNDR/54tDQgsQnE2yhIuxgYbThKVeGxJ1sdzdMYWsAd
O50s9TiVZHHAALaVCu00u1ftZrypR0Bzv4QzNO67/ctcFF6JUF9InfnLf+NO
HiTBrQ/u740b9oT7z44vra0alNNcAQ5PgXvgxnzBeYQGFhP+WYxBJKemX3GF
o1YSFF0ewrxL1G6U2yZCKFR5wv9nFBe7pJwOBHpg7zt/Wtpkuw2LCU9cAD2o
O/YOXyv0WEczcMHLXSNw94XfYOBsfuxyTkwKYKpqRv9U7WrEE8qePv3wpwPA
typVHp47WQe0eKemBVNlrz7/F/8PniCmhrzrkCG7e0ZptmcJsq60b8fzAz58
Xm7eTXScxqEdTxwoDRZFDj6imgjs5oppdQQpZwsh3QpdQrmkRtMwUjXppMZh
nLDgahb5OpfBOeIEIEB3RJEE+SblLDyUVx0/QMD6XqxaxaLvv00hwz4/tMKu
k557POutFJiNQHVQBCEkCSxOX+dr0uDmwlVzRAbqpArftI6nTlw+eDAX8jSh
+vIdh6M9ygOJMT7NHginZEbNGQe4lDUpg6uh+2KPLkP9kKc6ERBESyLwwL5j
cnu/h6/qrPdDxYbVmD57IF51OALraTQdRV7rOCVFMAukpvql3vmz0C+8HmBR
Ml4G2xlA8GhlR/KzC4ZqKwczg90/PYAnvU/NUgSqcmDAnbKn9qHIPhn645WW
l0m7n02ezV3ddKKchRqDTSqzFSD8X749OKC4hOcTU9iyLQaj/q+pkfFUw7o5
JMKALwNYPNQdQJ7ZNGEiGpGIfBVgWQ6w/81zPPTyh8AdKGVODexQww2sfvTj
xAqeCXdmVge186bdubKEM47/dSpudL1/X49fPrJB5fHjwNI8Hg5G3aiePaNd
ViNfJjp2XMzwnahKjI+JG1ra+Iuk8QjapgQvaxDlIScF1WAqQ0ALddpAWNPl
c7n1HwAsL3bCbVShpbN5P8ymqO6MSN5KwmPltApkVOOOh+kp2di5kQvi9ypk
63mQ/TGPinstdXoqh9wjo2PgzxZR+JY+lMdTHRMpENv1L60Ny6cswOOTjH6/
esIsIrP5gom8wPXyCODQTPX7XkOewQjsi+U70rZepkXckibyIM7Dd/SbCwEA
DUym4hHgc1zXSCXWdWvXYP7MZ0RdMwW96SBzDQ+UZkkRDrAPuCaq0g2hCx2w
guEJuc7r8LC/RyqWHvPJSfqSiTk0KfTl0PkJG9K/kf6gvQbL/Gerxr81kaJL
FON+lpUKrWZLICkSPqHHtrWDToT+qOGa6pidPlGoiR0VAFv9UiED9mNxJEVv
waG5jvUN/X7nhY7d5TrJqWDr1xd015RZFzFGGYXl5INPGXZOZu65+OaK8Ejb
d81KGx4UWpfjhmswHkhT1tbh0xcNUD/OYrHFPTnaK3rHent+TQTxhtRMZ7MB
sRjtlV/5MREa97SP6wJ3n+NZ5zw5gcf4g/tWylXdt7hghSgKf7Cf9qy5ZMc7
9TC7tM1H9dVYTqldWiOLze9a/Qom12Pk9TFGkP4wn8VsH9h7k00iXvMhD7Op
pV6Zlk06UaKS0SwNhfsrJUpXFLXCy1slDBo+v0XtNQo9rxU1QsXH0ep1ZEV8
w1qmQnu6sDlt/3vZVPrgegk0kOYOSPYSV/jAUqVlLmgwEat+QurIPFRwrucn
FKDPTwH5ZSvgKfLzRJQTqzIgWFd7eB7dpUym3mvy3qlKngHLvUmuffU6eeRp
b+3Zx/2cSJzio4NXwKoZaI1t+CgGfcYsXTVdLLgdTg1EQSnJ5zzHI7VX8rh1
gfXssrvQLCM+Zifa3GB1oL03Wvul3wf9D0AovKrZHl/n3I6m+pSb31MRHCsi
HymMt4KW1Kv2DvG61at3kPUvKgnOWin7kFlV8oV/Xl1JF/LnF72aRpT05rsr
dDzW0pcmOudO6saLN7Wwc/f5N1knvhYbAXuwe2AZCo0rSPcP6aU/P+WmP75N
36RSM4WraeclDFxFzyU7HAcjMRpOwS9BrBkwpCX6EnRgRYCT/r2iMXeJ+Xv1
EH9eDDhqFQpoKVs9wDi3TAgrM8UTcbA0OY3mMaRIJPBsd8m8WuucboU61qzL
1OtDYTMHIomP0aN2cQsck0MP8fzOw910yFkWWL3cBkDQOxoXzAjYYyHJPheg
xrcmi7dvYItAw7PmdJqWgftMCd7/vxMox+pGKhufCHDvDpIy6nTtgZekC++C
IywZKf/i991EcoAsV28JKT/XHNsCBk+EgcMmBo7c7zcR/g3M6bSC+ypUbqvx
c0syxqR7/KjKYUSYtz9Nd1nRKuIg+ESqCjwfDl+LEnd6fzfU3DW5y70C4tZx
0iwsACKQBRVmW9ozsCaXmuPEGeLhcXr/hlHlnfuvgZqu1shuMDfS1Q545n9P
oNAbqQeAG/251l7x26vJGwkqkKw+PNcKRKOMWoc/TCSLkOIadPAcjAx9RtfU
NTKToa84mpyHo/LPBMDp1TpJGQzuZZJ6JnFrIp63VnALh4/w1bD4w+h9T/WQ
Rp4UT30RS9w425UfjdRZjiFgAnDd2MH11YFZ28XBNDv7BevcEBELKOUJO+xz
PKMIirbYicGCZdNFQ0M4pmhtK2C839drF92KWB834fDrT9NTDm42i33ZSJkI
IMBRaRGgN9OnNWvHGNREOyso2aCTU3ojH/JYL08Jr1eCwfCxBq2cdwFw2lCm
PfJokM1pTjdFmj2ZplrXvrjd/QabaTAPbGhL2SjTFnW/xSkdAJUxewuynr/e
9CUktjMS9YfMXVykrZ+JqSDdN32YoRQBsSioJm2xn3GoNvI05z4hHao7zfR4
FiGGVxaIpZopvUmA6Iq8YjDIBb5Vci96kVgNHL/hLzGrWolIYBpITnlyRjUW
GZp3U7A8XJamZcaurs7AEACACey6ZESNi948jZI6a2Cg33aza4ZIHcbuJBb8
vua8nUw6ZURPuO5YbvsNwWPOKewSc8IwH1eAs+dsLxTCIr0qctpKrxqDY2CH
LormussZ/9rDH8ZN+tLh3QLfAzZzYH7pYJ/lE3TVokcOk6C0mwVQDrQkTEMP
9hqZFKRPFWgzQWmX39cfpE4QoGSRyw2v7QC3xpMDjWiGr6OeoUhBV4nk/2dE
PgZ136f4swswrugLfLjo/ZV85r5KqH1j/g7Ue8N7IlNXE6WSSf0DhLBI6d8q
ZRf1RW224ZqZOGuH+l+MSZZ1YPEonCX2+I3LbbHGYCDffUQNA2RNjjpui72K
rqDX+LcOybpcDFsNqeH16fjAY0V0n7m5pntoxhK7bBSaOSD6vCv2Vc/kg4PI
cGy7NSrVxOphg0RS7h8MquTLA8Sb4xhzelBFJzK4lqzfDWKFHus0h6DOjQJZ
Qd2XyUEXJYkB9/l9CQxKh4eynRG4HNO78nJf0N/juHjofdDWBMRrjf4c1WjY
QO/vYq+/sfRzuZCik4oRMsnoIFVJHfB2yvWg+YYfAjvOrS+G8mun+UrmvVHE
s1YAr/8kvOCW5c8TEkR0aCsv6qUf3IGD9zWMIWEhwY1Kwy1KZtlTxpvkO82M
t4adLyR1xM0EVKpO/B1nRrRRO4dIIueWyKcXtvCTRL+pKnWDLdKCVXxqhHM5
kiheN9QJyC6k2YH3mHUukK14TyU1TbGQaDiShpHU/tlrm+oFDrLP7ul6MNpY
yBlzn/cb8e87+NsDQm5PBbI4giK8V/sYSqEjsiibWSQBgUX5eEwd41nxuFbA
prXznP4vKcHjtA82mDA09ILNh1bXb0KbHxW7pNV7sSWQO4/ww6sQEX9UYJNM
gyg6mQOYz9bH8DrW9UQrfqJLaQDP+L3plcQ7xRGhnKAe7qjEuwZUK9b97awn
0/Eln4jsns6/VsOdNnumVtHzVUdfnSU0aaezfpQopJe23pIa27YqWv5y6V59
hBY04/f3IAwwaMWMNREjOQKJLKw5Po+akJUeUF0usCexJjbAjSx8eAGB0EtE
RC7zDwHiFqRDItT14ZcmQ0tkDNGf0TfIdU1oeDdWbK9SzG9KzU5HRPYA1GCS
h5jlRN9ymDIJBT/19EofjRqKM4jjhxY0M13hhw0DIBt+b+TBJPla+ltkAXPK
dTLyqcdpsQwuamo0A4SHpIayXqOzKHkljhKU8yU0HKpocsYqHn6jPBj+G0g1
3O18kb1OFjgyLNvzFKc5fsNiPMdMQ1piPTMfWTiPxuSbIMsD4qrNj5VIC89D
/ZUCEp7IAzyML2FBiB1PRHNES/FCigz6JFCLBfSRX+jDzToVS05obj/eTlu8
eNIDj46MVebA6oXQmv+JddyH9P/aT7B5DwC8FTmSzsKyQkiCUK7fa0WDGT6a
Wsoe2v9+Mth0JYf+zlLMwggS7URew4eJV99nWVWAdM75d89o5pBbABYT4ErH
5pAJAQnflDXGxc2MARHtIBRXyy+ZJLp19q7chncBD/VGifvN3ZWyoSyqvgdF
H1m5+iPeJda0suE2/kLmq9uZJiRkYYMaZ1usviznnvEcnqCJd3Sjmcw9rLGh
naHeQbhrBpfNvglyBhfp536rhCS90KoH42XeylviggS/DEtIwfC90w4dZFZE
EdetexwgDUW/vt+LGh4hUK3QfmbdCR6Wx9yUy4Ff3jj1iFZeo/y3+NOzqw4y
8jz7UEDbumhqMBKTaBvEhDPViT0R2+UvHQQS88FslkzefFp9Ng17YbIoxlbs
Up31eUXSZ7FTansX947yiNXakppk7fUK6GBzRug1iE83rGEQr3p9gBDIGLw2
6sqA1dweq4IbdfHEARS8cF1Bs+B2vhoj8sur+SjpkkaAir5Z88ZrD2lsqVy8
Rz9qLd4vfx8nSjaSLvhc4MIO5adnyiFwJ1w+7fGfYjU9xwyJuyxdh+Llpe/O
CbN89EZcOAnDssH0wwOiN1G2NmD+Gu7GnPTzTi9h+MkXNHwH1yazy91kLwNm
WBaq6Zt7iM2tL3ys9sS17zP8s1/I9bzfGbQy+jfnypVKnaEZ2OIy5KDSRLzR
1pZn7Irzm6VF+JBSwZXEyzJo0hQ8qB0injOzKVjQf2rauMN9rF3J5Gl2/Hu3
qLq74NHbpgl8KYPB16vqeVR5JpdZBG5O+z0nNiAr1ii/o2IC8uoD33i4XM2J
DFecl9y82m1yQPZ4tqXqmXyL/oGWF4DIu72koY0BSqhim7dk/hbAqfw1mPUl
HP2idJkLy6TL+0LyMcLdogiVjmW1kNmPZQPJ9MH87Ir6/xUuQshvW1A9H5bJ
cjkXu2vedRauctI6jOLs+a3Ly+EmugJfeaEYf2S00t9tXFhETj6Gd4Dfu2Xh
WIqRmmRU3vXWoY5T22/ENWurjDRQgutpfgornB/IRqsoMm0eyzJSt+X+AiJm
utrXcRwim61c5ry0jUI6RjTgztWrrPR8op32sCfK67DmgOZv0ng7f9W6C4lR
5b2zI5uEN1YRUwZjvoNxrkb+IdFfZyF8xmT1yKNnaK+jREo45pdyyHmTllak
DmPcczu/AxyUYxxZme5MeDx/GGmDjwPChSf3//NH2f53TzdL9XEe9OI9Gk3N
wTJViWPGNJ/SzaMxxeu9l5+1oGB9tdaIe78E3wM5kb6zztWjIPhR99oJiwpB
JZ3xzTwdmA07ZpKBYppeq4+4d4uWm0EAV18ZvlQl7EQp1Lb/Lsuu7gzBhEd4
geawv3VDi2bT0MKOusPwj/6W4+C7rrByjNRV2bJofqDle1EJtwtzdjQzz5UC
ajxoqoS5u9BAknGZJ8L7l0T+tVqRIeZckSPMBc3bUm9uwpV/Yp3r6Au49DPs
LHmn+vmyOIcwrhKqT3NiziSGQ4PQUGN6XOv8B1i8z3YM4U7RYvs5J/qiOWOc
ShxBsvXhagZaFXPP2CWBDQsimhxR/o0yQQTWSV+HWYcA0NwjyYn/6kN82hEB
DqZ2g9jKscSHyPcpj/63d7x2tJ9pp7KVqDgn0kEHFX0Svs2bIypjl3CiEPZ8
6t1orzwjYkJlwVdExjQas8zkWZ6ZX2lauNk2tXz1I+dL/dOBbj1/JsTGAbtG
rRJn3ndu2wuWTwJcdp322Cyl+VCuvdshJj7ep2F2PUrY2r6MCud+0anF1zNr
ttbycmJW7h+Kz84GskY6enHLpH+wWC/rZO8R655/MIyp1Q53uzcK/6YI/NX/
cmTLNKXRHlYaCeWXz5ixpoMuqEzJyZoWHsjL1pZqMJyWsC+cu0hjN7Bh4YKL
Iad8QnE3OQDc4Bs8B/rhLDgAfkqenJr9r7oBfle7WNeGViHsNM/pp8tXUNZS
WQn/SRog1i2nKQsKxlYunl802DzUqTz7cJWgEqGfEgBhiUPWO32rZq3dU1uw
nK5wD9pk2UUvwMVPrRxfjsaa5SRpnnbyXXYsghnEzM+/b5VpI+bZrCnHo95n
FAJ9xit4Al9SGx6UrzGHJNPv7cRgZYXTfizhSn9NFSGDGyPr/ujWJbPyw77k
Niabq3YlDF3bs+hHYkV8NvqqxQ6V88JZ+eTo3sblxXzUonpgx3MDR3BxVuWL
Q8IblnZP83bMT49szJ8MKX71YB7jKedVoi5MSKbLLCdLAYlInPx6o+zZ6ghv
y+qTw08DoPOStjeRBT6CDp0movnpTWWI7fK3ybGc3m+EdXcAqkPPE1Fyb+Hs
k6SqTZBWUfxQ/bKeadDt+jT4wLU6hW56Hb8FEH9Yb5gZ2kdl5Vh6K1QpKar7
9rCzjkAUBdO3pVdqKBchZZCW0SZTj/1bwPzprsM3TejG4cX7sWUDSiLF8hwy
w93rCwYyHvKc682gYUm7y/6ZWScmQiU1EmbFwVaGDR4JwQH6XNglSwx6KT/f
F7G9EC1JBOx8qoyRLPrDZKbFIPNyXh0G+D7dlmGC28ye/1Drl19xp8jfHWWI
Cf1jIBiJtzCK7KXYWZUvee/x+L2SoEbaW+Z5ByedO9GlVsyxjixzEsDUxK88
VYwbB+ZVgCpV5UNgHb+C5Hfq9CWm8ZNRCJVkEJbeaSfgOO/MLECtjMgch8C5
sTC5E08VQn++031peAFjeaABHI7kx0CxiTCQyIvG05r+bFv8rSWCp212cOLE
oWr8wRMQncaQh9mnc429s+x2NTVORaZGCXMtIqALTs6Q9mrtqfGaHF5lmFbg
rA4v+ADRv+Xdp9HBzHbvlaPE+qzzOBMtZjGfPx9kTgwnsmDto7OJQgpg2xaJ
umrydUDB1HpD2FPiN6gang/aXI/M6FUdc58dxH4G4PtbjFt98SQZk9CTQcfF
FH4F1emcPcJtc49TLoWq/DyvOfwXjw6tji3vwJ55Bm9AkWoKn4kOYvYxaiRs
E9mhT8/NveM7LlwNbRVmFCmLjmat0vqFpX8pC7fE3dAcBxHcruAaBv9dDCGs
uAN7wssV3GrDeTz91yEWFypA/+tpcxnYEplnzhIpTHxx+RlOquErnh3XFB0y
4CoPfyVlgqG5ab7ugDis6ym8Hhw9dz3my8Z1x4IiJ/CprBlk0KX0ciw4UO4k
WzMTod5wAcylz4Yz4EuP4JMZRZiJrsb/lNOU8TU4IbQXJ0zLV5o10npfZYGs
phB1azNR5zMOZ4GTQDBLG8MyOe7T4nODskoKxBc0U3f2Eb49LnxbVcs0SZib
t+ubYodqDgve70lSS6RqckpdjQCETgoe7wK5bSaQsgX8rUXD5WxWCzRX1XO5
mZgNw+bD+wz/nCsI5vthUfpXoiZfQs568TMkAk1nRM9nM+aOMN9QqZk4ia9d
jQpMoUxAI3kPfU1ILsnqx86AG3WD2bW0YEz3El4vw1dOj5kNXoyWuHNQ70Wb
E6rYq1a7GZ2W3V0qMtilfSAPVeh3crKjs8hSMHsi8MC6IFRKFSQAgxBHQXFA
zduuOFb0iT4lg9AzTxesjcA6KNeR4xyUKujooi37dGnZEiG1gZpOJo/iSNkb
8GhBvMNCETNVGcKacqYCNPbccuHCsfPV9VuNWk/NBtAK1clKc7QYkCSYbSZ6
r6RwpJ0z1Kmf7aPxxZWw5lygk90BYhOm45YFFyNxZxYddCavcUpbmFBXwInx
b7ESY9eymcFHWnJEo7/5tCwj6w1cus3ZNiHF007ts4IEbCaqRK/b5PDqykc2
dg89SbsCpm0774oo/KYiLVyWrXRAQ2c3k4rgq2o2ITTxdzNYruXsxWeGA9Xp
uANs1rqmi7uhfy/TSKk65X/Y1mJZbvuXLLaDJYRyUCxG9ONxrzNhS+kBX3c5
sxxgUSyGi3YOGb3YVUE3IH/Se8w33k+LQvXabHmBl3kLclfdzK37c73Vm4OO
uXOrv1xlEFRjwlJjXMocECS4Lyq/Zku2G2UFYaFx7ftiaFRVs1+CAUEF7+p1
R55a56bd5DqHI3OpAhMxaA7FyGzdVKHd8zHbzhA3S9YRdpZTrWeFBnxzad2I
QMbzcDiwLHa83yzfMAGvjvAquV27mVUsVvwE+WHbgPaYmDC1ieedLXEUVO5U
N7BsXKu8fT1Cx5cwWssLa37oQg/YbZQbNJrgknr03w+NxQ0JwPxZOtC3XsCu
oA0WTOx1R1Dm6eXe9F7RScdMx1xZCaZPGHczSWVL04DfOtyuwo/wSVkKlFX6
YtYBE2h5zZXOzIhVpVfT7FowcOT5KjuDcsgr0kZfNBLVdDNGn/e5fiBDZ63E
2VoYJLo3UDCoxMjExyW8wW91euVF1nIPQnXPnjVo73Hnh5FVa4hse9Yp/Lix
FEh3MB4roDGuwKTIwlx1+F1z/YwWGROKSHnZQ4XMDgCjRv7+gtJENROlyGCE
JeeKDJJQjPMi29bpYFxmNBLAHWaZZ83po9VjD444d9rq0KHJ38QjpktQ0U6n
hZI30YgErS5WhpS7uL2RUMaOdPKJJ+dCRe7bumK5CZQYjzLLJo3QRDnl6cEe
LRLICRMh4PLHTCirR1bTfCBEbazHHeM2MMin1rmYWqiBPs8vS4kuzZdX7jQ9
PcwvWtREz2S19ocxeSp+nCIOKb+ZxBWYDBk+fnuJMakz7H2ee8e1qtpXW4L/
uo5JsrffAAOiKoYkCk13Q/8Lah7g1ZTEvP+/4b15iCWCeuqo10WeluO7Izvp
TKbEzAgZSjgzeVCZcMG/4gZ59OIEor76dz7y4AkZKkIyS15mBSJx+siuQggZ
rTRUKuluzyM/NoGXgrRxtxtOXzYjLReLvOuhWOFayvGNYNJ+KdvV+j9r3Bt5
imaUlTBCF1+C2bdUME1pqyksKkgLLGYt9dx72QWI3CW0iAONm4wb9qsdpPmH
Hp09JCOtUJnvh7MqXMHaLNOndxzlD9Dphr9Qu8uQRtomytf5aRbiWdY9Chvc
OV1yLJYhmexHniq4ONsX1vE6gRmgNenmeNcsB6yD78VI6wz04SGOrJhUVRNT
cQbFL3Kz8K6lF/erhZp/3+v69Y4M5Wo+EWtq021UOqT/IGOWJLZWTKHKwGhk
MhPdSV5HMmMc5uiWAuA4lWaFk7d6A7CzUrpH9THFIKrgRHsuELpZu0/naGuE
GS1aitTfB01FK1a+Gs8mr+mOcNMvjxj0bFGryffYDrSkrqf5HfYQjSqNLD22
2BqL6OA+P0JhxVtssmiB/q8sl/xD7mQIoriO3I1JMTGwQDd33Lj1EHozyCtx
ZDDXyj3x7UAQ/rETizjg9kBdPvbHjz8yCszBA4WmrCRJehRQJn9iBoYVyReJ
pOFey656bEuG7NV7d/e+Jm3B5QUwJfSwJGMPYmjPsUKOfRWxNf8N7A+qmuMO
6/wUGimHRvUhs5KSLxcGN69lXf3SLvbRceUjyyIRZzE5x5XCat98z/s+7CPj
cDeXo0SkQ+HxjP2I9v2xCM/xOPEmJA29m2pPMIEjcd2KaC7I14TRSCxhEDgd
PberU9vExzZnMIpoEG4UiBX2+F01CpkLUHA2jJlv/53Gt+ILrh/mCD9TrG9Q
/7+8oJmxmbd7wUvyDxOiLDTnAmdQG4S4EKpgZx3f8OookRA5IKOj2VJJti9B
rlXhgMkuzhxlocWKm6qilfaoHtgxo+1B21n8P4cTnvnfbbtV7ee3vIB14aOA
4UsRHTiORG2csf7bpjYYLgyDsaqKCF4Dd+cxj+QXaMslNTKqoOkYBUpPb+0B
8Kj3PhYcDTOzdjxHaV1N0aA0CWQ4Lch1GD2BqP4LIYdMbBiLI/q0bKy4vi1v
93pXg6hMuShU4Ox8JiU400wZCcqm2E04vzf9sOr+sAf4wAeKGz5KzgH6EfA4
uKXSnn411XccwPOqaja4cfT4/h3FCPsrbqDP3DjWVnaD5F0FP5k4x72Hzpd0
j/idLaJc9Wg+vWDKx34ScnSycBcQzS+wmy0XoXxfzyO5G9831aSKe8nvaHyK
MtAQcKBJavN5VLckmZPOiPxih40C/Ddnba2+9yx/5DleTr5XTb4oHirnjVxs
43CdDAqBfGmkT/3kSeHzqTTBIe/jjwucoEOw3xAANkWFKWMBDSx3DEZxNPRF
XZW04N2dVQ48YnXt4lJyEIUFGItTRG0PdP8XPx0TDrrGN7XnTp8GjNBFXrn4
paapSkEHHVKStY5M1RDQ+XhzQHUWlIKOAihvStBkI41EYL1ASBrjItdzBHEA
ypK+XM9pALSN5PP0jCPSKKY5RfdBsedWjoNTideVL84q5UhUmD0zMO5ioHON
r0oUJ6XnbjSXKMnLKTCABzjSkd9iHVb3nvP1bGS+dhfSrj+h6Ev+aUtt8gV3
ULRTgtHuk2y3WU389LGUQgUazczBGU1uM2GbqS0P33l8nrrUH8fvE+k8eK3o
+xPfVnEwXgmehfLEumF3U3N2r/zukcdfid0lKSyX6udRixAPKaxEFruy0gju
6OdzPc0EwZtLY9Db7UFb9TcEWOMxKORtyBNLtKhBPlPRBIX8uH79rjf7e/2R
wmCBt/d4LbhiAbs9F8EXDN6MIHgM7FJpwKCCUj1yOXSWI63QlYvaK8nuOthC
AZ+8dTkKpaz5x5MDcjfLuOimdcBGptHcD+1PhQp5U1M1RBE9oIIhkaa/ftdX
ShJnk+7WX/Zem+SQB4Twg41RWOKgKTYSXDlHL4CA/prpVIzw9hcd3AgvBTC4
b+/5jiKAx6vXmwb4fM7TeiPvI0wo8QuTxrvnIeLK+9muhclzEf0rLxdQnAuy
jqUlIkX1IZeLikNaBMingsWwGSg4+1SJ45/C9lj43kIJWUiBcfk2CGb3g2m8
t3sT2emn32YO9FdOF8j/81EKBlJKBNCy5GJteKyvvptOHXaEZFUKEPiCcg8w
FPwE4G7Wmmqb1ITYnucsJkTkVOrVQkOnzjeoDiuDR/gIMizJEmTu+0Ll1Ysa
UTFELTuvulnDW17tyxgWVt9yncGf7C0rilNtxYC/dCUrGdIp4rWeNtVc62Xd
gPXsXr1w+qLMmmntQ+3zMa4BBfqFlWsufWuynZdLl8G7I+wskek9QCYSJb9/
R9r1UHXRN8Wiqfcp16tBfC98UO5Kq4DjYrmnnGLOlRyuS26q5Npr3dcQiaOr
S2WBh90Zm4WnlknES1FMYMFiobGTme0Jf8CpsOa7m8QMq21zxm+6b8vvV+GW
Spp6h7p59qoTpI4OA81cfzz8SeA/NDJ+C3SM5uNLPcpkV1PifcxhUFMO2dsX
wSj/Xpryp3795KT1CWtTM2zeq1ELfYNzQM2TFhYq4I4+3SsxEUZTzYorYQJy
Y6MX3JkHqUtWe5OG5Qk9vS7aGHaMLQ2zDGZDgV+mU1H2OaeQKUsKu+BR+gqv
eagJmtT0gzdk6WqrTYBJbIo5cOaTihxOjzr/Uuv5DiSL7TbOsj9YXKw+De3g
/IT9Ow16K4S5vjAaeOBZ5ZvBgpoVDnyTjXohz3onGwKz+8M8d5rBNR93lVWZ
z4/oAlGOAi7OKmmvD8LfWtaxChY7RuMv2/IRDuIMvlMuXDnBj1Qr6VmtZEOO
6l9MUoWK7O9RMb9cx5OcKaNyQeaccC/fdXPDIyh3wkcjf7lb3hKcOJqW8nKg
n4TMq9RLrL2A9a+XEC62V2mK0QWvIgSObOWFPhh3XVwQ1GrV1rJMVwB1yY/y
xb+qHl5RtIxIjRwdWCS+xDUhscNCIhaekmulqbFEBh3kfB7HFZ41QLUguE1o
fQAHc3giJLtLyIueuBVK19m+EHMcsRymjhaQxrjkw3+oPI3Dm2e11efC4X1Z
c6SzLMUxh4PLG2DzITuebAfjzoPpMmhVy0Mgh+rLP6KjjruqGFiEAO7TmPEP
nkCXrTpPCgq1i+19rzeL1ahDiKhtcIxsn/NacHVHShxCu4dO9kEVioXc1zDK
nQ0QtyItHNc6UO19OCeH8U1Yvlo/yigC0JiJ7V2TZdL6e50rXNYNoGG9fEZc
ss5OpWd1ZjR2VBfAaN46BYyF8ITRYTnBuGe5O3lxbn5d2OrywW0cEZcyTb5a
309k+yHw6niS+gVMbhXBUECboBvwHA3nMpvBVm+EWYUJB315A5eCdZMAjTcj
1YDvVm5+MwnHuI7d06V32SkO4B6jjLNVUjwoBu17ASFAT+lKeS1TPLtZUJ8Q
NlJ+Wdu8z4FS45XhH4Dda4PjVfPB6wI9Ir+HDGhhcXCpytL44Vc6hEM7sBel
X2IVsEEdLC39vgFbGkhZ+r7kDst5l+ow4xc9Q3vROcQsnYeuTISPdQZTSPzS
CM/ItpzrBz92WRZY1x4nJJ1tcgL3zBo/VMVNANaAeiSD6gvh1ED9D7+D2uGh
6XfyMUD8cCHpVUuCZWvnQrRMrKOaM7fIZOdf798cTj3l7HzaLGn5FZRdV81g
dFPmCWnTt4tJuAVcP0tbEkNOae3qg/6DKCuyCEpA/j5digJPav9qPrScdIwc
7AgEgnyW1Sbnm/tvU0ggXU3A82RVyGrH7FZdf6UzsMKjPNI1veK1u0tFbV8u
BKrDZrr1A2i9AtoFPDFvaYv5A19TidRzUbgwbcxgw0jyvswlv4dOUOCnsXyF
jVUH1nseWL0Xu/MGycUPNQrlWkpeMh6IAUnZ67dBPiHrJn983a5mTphxnRO/
F7mxlsbbrXAehei6Dz4sfCPXPL+VBujMhYowRx4snn6iqRH9xQbCLzZfg0By
gO0kQfyTeNTR3HWWqVs8wf1kaR7/pU8SR9OcfurPQqC9KfpNDoRwFO0aJo3x
EZsu0K3XoSNAXTln+YcA6RqfpxP5ACDPlsFM1anxsrFP52CfPavGcF8UVDQk
ObPRpYrIz4hbe9Im7ZisbzF28etALjSJ1rsxA/5TYlxTM1+eur2Etd62VP3d
rH0/LsPhAxHZxlVkGepoGdqQHceITAYJTYO9Nkhh+6tfWbhwsdzGmwa0yrzl
RrMS0zFYKHgKWim77k6YwxZv9QsZYE5FFFmL0pqbnninzmMyTX3dDjwwfLNP
9duI/1J2j+t6Uk46cZwj0cJNhRs6P474qCdJJTPOJs6Cvinl1RvtBuuNfJ1B
c6eHNj90HTddJJem0qni8b+kRFb0GOxZayvHNiKzxAJkjNuKrebXZ0OCgAkV
+t01ha2J/Zca952cDdKkJ/hlmMxUALMUP312RVBmpqFW120v2j/Sr/p2Gl8f
zUU7aOzsWkxgY8upv91YO8XZVlJiwZpy840C+e4l1WKcOX3+RrPRz96KltPB
5EWezsH99m3Z7Zjr2fhdp/JnKBHouO+DGfiH8I+PbnOz6Dit6Qds7alBFbFJ
s335TE+0QMQnMzyK+M9xSkwqAT0XjWJ3IKBFOyCEDTkh/yMk9rbfU7T5Omp9
JBWnMVtj8vKvc/XfBNFZxIqSQhnzWlcmUTW1bhNR3XhyBrPbGkcWTOlqOKpx
bLVtdrxmBGlqzbLQCZKMypjmibSRS8CQillNNmg7FpQhe3BoaZL3bPLSf9Wo
cZkdTELBCBGurewLb406OMRRdrU2ocivHNi0bcaMkf9FJg5WnkdofMfLU3Rh
6o2ldV80c4TIENxxwZH4ZKLf8Rn1sULI9wBeV3wKCKp6T9W43BBVYkJJB04r
bNLjAADe7XbrhSFcwNUsIVqqL8Y79KvDe32+rdUmxfgXt4fCu22JVI6pb1Iv
4CJhvKfXRsiQ/XEdOAiyEYw86PyAGPxTRteKEGirapcPX69Cv5T7wdqPHeLz
ucmKOav6ykddZonX5azrqz/StDXo4c+dNE3GPm2Giiulfs0kyB4bvH68/Uvk
jlEh9zwtxIPI4RVLIgcqfTUg1IMP87aHeRhHAPBR9QSYYxjmMh9CUruzLLlE
QHrf1tam1/KSTmhfU2rVl1hdwmANzyreljyI5Y4B4RZs3Yz1LpZm67alHOEl
mJglCnvuwC57nR97fvQcUTszra9oUTOCxSaZuVUkrQaKmESJkKAEG/bs4zXl
meIAk150BI3obZHNRz88kt9fNrAPa2z3JumoxuBVMtVAoEV6QGvOQ352hJXo
oRMEe7RdXoqP+blfvV/FGFvy1eS6pdNG2oGJ8R8JqgLxGqEsDkV/O9wwp/ba
4tNGK1dA3XCjf0zTlZTYZcFUjIWYP8YhAbi0WnA9lVvALSoyTduMNN0it6XR
VBMqYONivRgK+9YjVF6CFZAI7ND/XA2i6ucbbZYGMG74uJxFIrL+G3F24aWb
8EjKhAfP/58ckrrQzGY2l5NsY5iqNVACuXMi/cLhLF62Wgsruvx6wEatEneN
xOLWXKFis3f704IsntrjpJHZ8hVztgfwcB9NyLNDqt4YtqzKDmLqwo9Ac/pA
Zugauhcd7ERQIfwYmKVU4O9u873jM/M17oK4hjp+CbqUn+BBy/KUALVDDjI9
j/r1ceq10PF//iR/8cyWOjmu5ln74m0YCiqcDrSza4M4d5kgVM1735ANmucl
lKFggTyEfo2MIKeijyAw9JLnz1aP0mUHzhra678jjstOz8XRwKj3Hpb3kVfR
1UMEfoIqCsIgyG+pKVpEkQ83X16Hp6WHkmcm9vnEqE0msFqnYm5HdFrY3VEI
6pjZVBg7lk8TnCXNk5c5h2Vy6D6uqouIWHVCca6tNhwuqclMMDi7HTFY3EqE
2wyK7vIjflPJEBBdWSFpp7zrhhW1vUbjNg7fiojcQaMyVo1uTAObNAZ5Rsft
/4gBUvFt94/ZebEv2ZKzF0mDEu2icCiFA2f5TKqXZF74xqMVliEjfKgHXobX
23Gw5MbYUTNbn2DPdtJ/bcSVEaAX3Ge6Prcsn2WYghAH1NzYsEvqtEkCXBGk
lwS7UpA8jHmIwLQs+QEeARB1aiNtwTykcsqwGcYqBuadlGjsco8QDeAknNbj
ee3clOaPHmiKEkVGt2EHpw/tt5s7sso8sdlmq5FSG9JKI+PCkQRrUpnPSoEm
uDq9ICQLPly4cf6RSP1wdrgB7615ClYZsxCkbONjkMrFiazM2uKC2x5oPV6S
+MyzX/PF1fUvVp1hMnJoypT5MUSBszUh/wNPvRvlA3O6BBiFoDbI9wJI4a5I
gniHKvXXb3jF7hNEwDJiDMAeMFVwZLC9W3/qGNVTTRIWOlU8xviIZ3Li4G3t
eUM76YqxL2ioH5ZuJkXz+1FAEa/X70MjPoaThNm4aHfjf0vscJofeeQ3DqJA
kbVsn2RXUDX5zsLemQqQdAn28PCJz7rtUbxA8OzJVg/2HFDOblGrVTLW3RRm
fLSpcYvISCCfBYuk8G8Q/WSpKQ+BszrTnUc+2PpgfdgwImFDNGQKcURMT++M
lYpwgExbRjt6TA3KXF182IXh5HLcUolWPbaWotXrmjSP7C7eC3O0EQ/4UCfx
QRkfROuBUA68+Je58Ez994RMVwuBMZ5/TwLrKwFsIfhM9Au8ZhVhdtQqd5L9
PV94GhYfRYSHJk/5wKn+WVWAQsMVkEdkp7HBlRMfxpqYU6HOEg9lywnnkVxh
OQS0Wd9QASmMFiPsk/lLBNfknzVj9KQ0xiDUEES7ppdVocVOp9HZezFkVkaw
ZW3hEjq4og9ix0JjTvdrUZYyAICp35RgBxRCyCbndO3JvjxpC/+gYXBAnCc5
RdXhYuGN/alAGbvGP/5NTS9k3ZKsQedOyYjs5W8uNPxj4Gyx0rFoeFwK31//
Gn1I2K9LyKTGPkIU7ckdsoMXKG8DKBpqdSpCr2062jTbJAcvMKs9sE6vFYf3
ECcUvpORjsqAMUNyVI3H7Ny5wLKy2HgdXzupNbxhQZcM+LxhfnRWOyiIZs+k
hqMEgVuE3dpLz1coFnHPvpUi5BnkuFO0qdvYa4OmPI/vR1DaP0QDoxIDDWB8
eqMVi9CE/lEh/OZnXEV8uY4fTFe/pdmc48IaqsOg9WZvN2HmXdMZdYo8wjO5
2Xz2dFFAMGUh/cHFQty/ZDBpvN838qFySEejZB8drt1H6RvDs2DWctF3vTTR
66F+KkE8DOELn6cTG/66t9mU0nlqfgS0DSkwiOJOezellbzzil5uu6bC4hCT
CECZMRHdmFaoXSByFDwgYxPxsjKiVIlxw6JHP9YRUwuV6gGclaurOI27FkAi
kq535qhFalyfA/yT2mCY1ed1wd0MwJVvOMyaEOSI4uRt/IjulphWxnwKKu3c
A5tddpZZ0ELeuhButqBjbC3UlzBd6TLXe7fB5QIa/w2gQ8i0HBSpNrtYjGL7
at1wJde23OG+e7ahQyK61aptr8uIShyTkkB10fu5dHv4ccZgJG6gJZX/o1W/
XTqKhzYQru8GgG9fkGA8/J5+QRMPc67SH9nfUJ7OYaF/NQDn3zUm0826YaOI
2n+mi+WakTkXn9Je3oTFOz4DxjN2+7qqV9Wjnz8H6YK0KUipCqeWcyMBfrZi
PB26VxEgiqghKFWx5lNYQg1Cpu7a0pVGBP3w87n5AQlE3ec66B7EkhxCs3LJ
9H+4pTObaiLmDSh6wn1yXFSHFasTXG5rMLTBnF9f79IQsDwUH3+XEeU0Xsy3
gUK3sj3p4mO+QFIGP5namlrrNy7P7194sY6oNFvs0FmNex2aiaS2o5nELMaC
cWedTV+QHse7oGdF8VVuui8a+8qKFtij8fzERvMlPOBhZoSdpVBmb0x1lfbf
WeV1XP5XJdU58hRVUVkHz3eu8yzIVSEIhsP5/ezCPNTK0B7uQrahrlnIlSTw
X+gux8lZFeli9NO49yv5VlLYJ9/RBZjDLp2aU053ZzzlREmuyLM/2FLdwabh
F3PYzTDOMYXC/A0AcF9qSiFthGbDQMVFz2T6MDA7sKS3VoTHgWDLYxJPyULG
CaImOjsg365cnqWS8Ap6RNaGUBMnoZuUTXgZ7d9cAo7CO3W2vxLBMEp3IUQS
2pX2Ux/LieZNwSPTK+zQq2Coe+iIEkvyC22YXT4hXpnGXNTNg1X5YZrfd4Mo
fMwn1PWxrF8FauWDa5dXweiRMOlTp4P+8OHUi5tDwbG5Tb+j23Tcz46BkKwa
9RA8kZOFtmQ20Nas5cQ5igQJM9Q5KMbDDBDVl4pEdc3J8V9T3Wg4+gywrLRJ
Dt42vc5MqEo+ldWt6QpMlrZ5srrDiuDCETnSy+LsjmR4CsuVkWTNN1PErmga
/f3cSbBRI6HCg/zbnk/7ah19PNMnzKvwyi6YD2RNKFnKpilaSiqFIsfnhjf0
iB1aD7COPKWTBhV44TgbPlAoy/XiTDplfOEQFlpRLVsLP9F4J7JCrckDE4tt
Xk/b02+YMt4TqEKMxx7EqagWsfa5ziJCp/7vNBYlStVIAaRMohYIN/G7jCm3
E+NIYf8y66eIMXltcYcczl5eAAPKYTsRs2JWvdtAm3/p1qAHiiTW+MEeCdSD
R+rzwCXxlAOkdcEsWW/mTMX6VpyimPSEJf8zYxvBIWX+c3nDv64KvNgvOtMQ
abiTGK4H2OE7A5IjU+b2dNa5Lbo8OyY7iv4436Sr1u7jZgRlsWGk+u3T3QDz
4imxuwmlchZRf1azAJF5gxJcG/OsC3WgNYjqZr4OkxTnoc523mhP2Qu52//K
zXKJe/g+qxnR6ZKZ0J+F6MFkPA1QHR8/xYkfb6CZCD2QKsLzo1oNFFDtf87p
CGLS12NF7m3I0dy9bqIl7TP1PSK6xsYnNTaTAwbk3oNP6oGbQjaPazRdyzl1
OpQ7SeMGKs3cfRUb6s8+VNgPpIKLEH8iPNs4RPr5t+hNWkC6hTef6X3voCeX
feEBaBV4cVDgp5V2PkFBRYasQXE3vQQD6uaLJsZpvUBo/AW5479UQSl85LfJ
R9IhjepR9D/lPGyU9z/z/RcLsgrzvbNADRCKtLPnYa1Wkpvm+bkCJAMuNLB9
IHobee4EwhoQbD7D85vssVlxAa607nJiHmMUvecQGqbX4+goiz/oAfg5G45v
IOFg1Qsou7zXH1l+8PnwcGBLu+/Wx9LjO8onwAc5twStOqDQ/F+i653Yp2to
KBq1eg/9b1RpXf7XbHONbm8bL61dlaDBYd6P31+9RZ/a/RgiGukhtncAJpH9
QdxHTjIFXF0uYJoeFo9EMMdlOmo3cf52c4aNahfZJGmJ77xr/raTLYbOtNFS
ZueKOB4vtTgn1s1yfV6RwSCF1uteIoN9RQiyv+sLwH46H+jS7K0sA4ieVOfy
uMvLXEZ2b+5OSNXs6qt7IVVtnpu8eqos/A3mkMhRXdQpfyAtxis226Gfnr+A
uthyqDzuqNoFKqBlUuQca2dsxJOv8SX7H/l6RwOpxk6nuJNUxe378K67Yxi+
xkdDjR8umlsbAIETexQIIoNr5xD8KyrMq+yxpZjEaztt1EZf+W5CdjO1N7sz
ye7f+hNvONsWQGm/JKPTK+5uWMshA8H8JszIwQAleW+GIAdTbkka7qeo4ASM
Jpw2JxpxBboKWtmX4IooLHb9W6lK627whGFXf3i8sko/gR+60tl3xrTG1D08
H8wWBidFUpHNczp59u8BvlPDFAyOyYodq1131JoL7tDHekZazK4q6VFHBVEw
kabu5BJSreulMkX1v8p626gz3zZGUUy8IW1b8Su9YQIPgXIqtzEo2iqFwGdd
jWmTSgax+H1Yx70/z+k7q57K+Y1LYHLBTNN9vISEs05BUe0JWQ2Wkhl7tX2t
q3Wtq8ClMNU5fwB9oDoCpiHWQ/QvOvdoeCDzBkWmusXQ4HqWDNZIw6F9ld1F
53vdxEX5Db+EBsvYMMXLGrFVZ1XtAVPITho2qcXDABbnjXrXoNAF3Sq+I9x1
/EbO7N6GcgZc2I+9hzgUgax5nKF2RWkiPDjGJDA/coHjVjR0XX+ndZ+tjGHw
qVy78jB0MBMlgZTA6e+AAKKxviZIkhsqL0G7+kVduStQHorO3XhIBLKvbwBD
H4EUh5RWTLiuFWxiEV1KXegDyxIRuuxHcJNjZ3CYkxTKH7yWe9x2HgMxBQeg
xiknaGK0ZvWBwimbM7cDim8z2z29UhFJVC8kJHJazmEBwEsko2vrhQSJNS+H
NY8iMD3t8UiMvR7mdqaNnx4LlA7MFLgcDnWF6KbaUIccemSw+KxBDjq9TD6g
1XekuxhtEChV20uywFWtwooIT4YcZe+VDygDrkaB/E0fxusKqf2anOBPDZ57
U0SWhip+XwUmjuT1wrwevx2SlFkIPUVCIt5zZow3lYH0yYfQ0TMEg8iniww1
vWrpLgbb/r4xwQogiNZZE4a00nbOOg9OJ0Q7MfMpNolT9S/gcx8/G0FBycWL
HXlEaJIHvLcQ3YAeM+escdUS40/E31opGgI7kIGF+8ert0c3hh6cNT4mqfDh
UqCRSNs64JFIVD3b2KcqN+2ztBSeiW/cbGM1B3+bmxx6eBXe8/k5vhkbS+HD
m0feQhEm7dUlwOu7lo40CTXXtYxtg2IgvasikqKYVfGjaMVXmpvFIxZxD17w
xzQZ0NDwnNBP8AHCn6QWtitqCcsM7Ep2yNqEyaiFdiPjVrw6k/zwgG8XA9gW
gNRtnmk/LlOb7l92o+8wn3WHbOBJGphQjisuhfnj5fbbSa3ldUW/FmO2Xo+7
uhwbx96Db/hGc3y606O7aZqiDI6KaoSNyIcsoHcxDHiZXFG/3FhSZyI5cYBp
uzPhGWCGDHIxnmhyBj3x9Smh0nRPhwANM3kooFYYFQCwnQle+3Df7mIcMApd
rinjQog9w9I+E8pCAjwjXefZMVRTQTeVPyPRRsIfPoFK0ibh4wofnmo5W10s
WWMG3ITiOsbQeg8Zl8q+7JcfnwkI52g2e4XLfSzNV802eVmHLiRr/aK+wR/y
XR2u2Xy3XsmFXEGbkXmQWovqxGypQ3HKpw8E1PUhOrqyGoGCP5G/x+suWt3I
A4Iu/1Qhd5hcEKwEUiq5Sum9xmiKVf0xhDGOStLrAoS5L9sqYEP8ClcyOnNu
n7s2wQHVrE93iuzDO60H37Zju1hn7U6HvUyNBEAwlyfIOJ+W7WYXCu6E0iS7
2ctsqJz5Zd3L+qyuPQH2oxVbbDdG4WaTwiPfQyDwx9AQWKzIA5O4O4++9r8s
VNxOvhWJ58/zGp6HRjg2+1VHC7DhZoK+zky0dPdHldyJD4H74gvUgjGYFb6U
8xy10v5BhUOb9Lpy84plSrr8oyVLUY5c5AP2bu7JS12EMi4xK+99F1FbPSk7
1O9hmV81zRxJdwUIYgGkAOanuwVLCYG479/9m3NyfWFHnR06I9A/eU64vVc2
c3K6yz7NV4LY9y29Fsu2Lw7ix1pGLlC1HYKRHCiwBO8xPQzGKk3BEF2nPXpS
oZJw9mpVD0rfG5Iq3765DTzJizkfGB9TZ4W4NXI0ENap2Oomr04IVUJV4LZo
92XxK1FHPbxTblI+1DIh45PNML5b4+7dQTOPMBDZtFxJ4eQb0aLR7fylFC15
Aw5HoztWgr7dZi7yf/C9bFEBYeFwfSANFIbRzxYevZ9b6BfGdGjawlErYhbT
pykaK6qV7NajfUvdgMn+sVVEudoaPE1v0CAfeMhySQ5N4JRd+WTzB2T9mN/T
oPmanyUAYeJ1uJ+9jX840uNeLEufayvyxsSl/klAoUn/tFg8zn9UNktitQYL
fO6CkwWRmTOcXedFCVMbgQQFeEU3NQqqv4KMVNSltGqT6JWk6rVqEwGbmDlT
5VR3mXhOfBWrrXww0u8cEDwRfk2BUf1BRPdbQnf1Xiz9DsnDaUxO63GZuxC4
oIMSeJFhEcaafT8FFx0jvmswdYsStMQVmcxPzKkN081Cvbg8Jgz6wcd3YVoe
RgMESm+ORqcXdGsG978EQbYrh8JHX2F3vgUzMsHNMPy4a9blEGJpB5cVHUfP
N2UeX3kvEd9rSiQXZZYFyadSNvMaY/6YAaa+81hPN5/YKG5YOSn5SHQ63Gt1
Px7B9F66LHtIHq1q7fJrJCWcU0Af2E8UtYfL5oWppGhQmES0SQ0Ku1FywvVO
RK6uvUSS9xZVPrIVJoKCcNaOjnCMA91QD2m6SW/jVh2cNSnDDSHtJj7PcJu4
kwX+Vsa4d7v1wUdK3MeoetAHPv9bFp7WMstBfkLyIzpclesx+qa8feL+BD/Z
tTXSDxYz1FwYLWPsk7GKSVliCySHgQEctIkeA9McCfjjooYC1fHdtdZB6ZkQ
fLdvWuwY80JaLsKqdKAi9xarKcobx4eBTbP5OU/NFPIaKGGDLptAMQVD9nio
AdJTdmsxmTLyrW94ZbcOiCtTryGOV2o0iciWIhMIu4UK2iOQqMkvvGWdE3hc
Dm7gzK5p+pBEWTQx/cUhmHS1mMfBvSeeRGd0X4vNPhSoGxfuSzOOPeQxtld7
SvHJcvq9TfODBMADF26rZKbYwe8684t7yfUQ+ju1l3mZXrDHtg5stLNmi51L
arSwR8pfCGyOX4KrQUDF7ailIbN4wrf20FXiC3S2YpdxW5cp2VxGR+m8AoX/
8pULR7f253aJA2QpwegbKTIBMCONPu1bgHADbcBZ8Hs5gjbGgWT9JVE6q6kX
FjZazbsyZFSoelexxMwGXKEL5iBTDnDw0F8yUIxlpoL4v4/pKNY1uhL17RKP
vN99Lij8tZKXPaH+dh2O9RupJyma1RmWCC85UbKSYr4kiN0u3IlfmV+YEgSB
HifnOB6tIjIE3XamDBBwDwETyi6Pyj9h5XkNgi1CwFB5pZHQE5IrSjl3jeJK
ljW50N6V7g3SxBeUajiXZ3EWuglwS2Yx4uYDmRTuAfScTfzn2/CR6QEHy78m
JZT2J7fv99/mMt7qbp6bBy+rxeg8jHRiLmStGWLo0V7bs96DYu05yf+Cjxri
rvTx90qrXkxUNceN7zD7xN4qpIT/8MGLHvawxgvC6DDLWplOhhdpXthIXiip
2i4e8wrjcjHpgOAYqy3L4wc7jIP/XbCzF267ZfJIV/NnTpMWJC2ZUdiWfwCT
vsm1+qa92LyF5hNZ+xzpUn9VUU1YxgBpB8kjjhA7eOaoQB2Kd02NLtTnxD9C
hBZ971qckuSse8S+elcHOXYknet/3VV8NnT1uossp+eL+2MKboaxjtirp/dU
wlUda0WPfawOqHYSinH5NrFDGq8bGjVZsW9FhwnJ191qhj5zSmBGr+ybYEhD
aC6m9eJaqSReWeK7diFXAKwTSs4mqSt2doRmkD9JgIGJOQW/x49qQuWtKwOw
JdbuhUXA+lYE49z+zBSH/Lsi2mGmC61naqGcR2vx8Z6fsgzk839o/mTzYvj5
7SKWEt+u9HSLtwYj8jsH8GtZBVBaTRNp/87gC8ZuDqIwZJbL+9ToHDmvt92E
KSuhK59IGb9vE5COVUo6I03gzamBudymxLPrNEE3V6xUIYgDHR/5195NDdxu
KCRe3gAEt1+KnylqL+2wCubRagPqU0OcsG3F9ih7ZIET2/1xk5laYicG9JxR
D6ePxWZKSjkgZll5cM4+xecN2hxfmkKregBO0X+JoOnv9208oo5rWeYZvlDE
whIWe0xyjtJYcqeEsetHBmbl3vTTufg2zmDGllFg5ToHt3/DO6ct+CtSW/+x
jLd0c/dcz1AmkpRnyQJ6yF92P4XH1WY7tQcsbuHEeDmpPyjPp9psQGz9psCC
vTmiLXEpiND7VH26dhOSC1aRyc1TyRCjylzD+QCcUFpEsELeYOoWMRLZuNzb
zEFVHLEclfmHVOE9r044MnyHwrkRmvrUWD83mpdKSOR13VT5nCYggwRjgCTd
cwSgWeZogTooN/fkMLl4V3UBxd00yKw0cc7KlV+OjOoJh2nxmR1oB+9zkcKO
VCW0eamW2jE8rvjI9f4lKtZA/J7yffpPnm7rfmoR38b6dYgFkss40NSXf0dm
QmmErC9TVAEP6DJM3N6pELYmkCGkT/c9bReqSvCerLSZhOAT7i7hybWRb6fm
NUDsmvUPzN9CxgFGya72VS88UzAcVFV6VOF4AYKdANuP8AyGSGk9Pn8g+/78
M9MJnE7fCrE4/CaZOwHlaBoi1qU6+9yT0cLWG/Ki6JvJvAbARRi8h7GQksIq
WC3kdB+hx51cjWAunWlo+aiFh+JfhXPR301/KVxB32GWI9p4jELai10RLGqf
uATeVAVRSdL6wf2qs821zxPG6N5w7cTt1GB85ZmZ1mi8TopSaUhq2kY0IblC
IbuMmAv3Xt/DHuoz8FsivXp4q1wxPFdXCoCvfWvo7fQCKD+UgU4GzaMgb/Do
y1zy3JguMniB9C6+TDX47CUvyw3/byeVBohG+VpqXpw1jPLQbCqZGAmPtyAS
j15dUrcs3am+QsheqikJ5uVDqhbhcaUNCW0Ux7gcS8Tbb3Dg/x7CqJdEhAYN
U9dGi0CDknW8AO/m87ZJiVy2FpeUo0/6HXFn4pKlDVhvCAx9V0qBr0mfP27W
ZgWTYEBDwC4ghmnl3qeNPbPKtgzbLCbB83Ponb7ZwjzGSIqyJ08QEdB7KlCo
2nEu+lWjwmiW8ZHNMchTdc9Rgx56PIRYgo9C2+TY07rVYf0oeWxx5O4RhLCJ
XJbp9omhJ/E6476Nc5Vr2mGWUlSDEW4OxX7AG+J14t+ESQ6okkGLfNcEkhzb
IguOUtuLC76uzvTvZ481GOMqfqzMRFf7KapmQxhAXp0VES7zv9rrwASy086N
vXQ4pVaetvZC78WMKxMeOlJ1uoQIX3+z840bDTDLQQReTN3PZMSosAOcybIy
/UL7fn0WJNJhBfTYYlA7GiFgWJSNGoXNWfEsFumshKxhz68D09bTtKO+sNYU
IDl6OY5urOEQZvAHfoZWCl//ywaoQ1QV2ny27kgjl/3aXz+l/f/j5MMSfTef
sfD1YujfLa04PAoJhstC/HuocOqxUUNMGZcGk8H9t8VGfI84tj2AvSGyL3xJ
CGIOWmE82l+7+B1DFSj6vKSFE+19CGYNAd4AZUFup1c9fwyoO95oFCWQ5Sr5
a5nFn4kp36awN9hBYpV9mDK0LEqItlb9mEFNE3TvtRqmlwbCkrDMgMQjqcOM
1qbr23SOpLv2rxUo8m9S9EgB7emv19eYfWOOgb1bTPqU4NUkfLxngw9qqQoh
Di624SKKVuviR2nxXtf1LT+csYP3sZHr2cJiXkO6APrpWQDt40JX8tOGfkWi
a4xBXMnusdxDYFJoBNs7d+mdvd3uD8rDYAIdDxGlmA7230u9yonWtGzi+awQ
Uxwl+fLDORWGwTqHiuuInnigflu2E9b0rn4uYUiExFHGZePTEw3Ad5EXwelH
OC83idWU1VCNDZWFNv5WdmY6l1gAaWzPo2OsyMgOFM2XcX3BNjsdY0qVMvj9
WVxZdA2mbxth03l6aJ3EtgenEZ0VCwVL0FwJTUfyvxaLssMYdxiGTiy0/88K
Zw9PsIAmbCOKZiuVr2jSTO6JbAYtNG3NHU6LSQGOsd9153isRJj5lbjM8AoT
VGE0RIrHIs8ko2W+iE71/cRHN3xEG3Sw1Y2CScpwh7LbqpMivxFEqWBeqAOt
8pNNzhPdNZfzlVUw/MJ8w29VLn+FFF5Q64/ULahGr/8RiwsgxrC5vIwe5U48
zcY0/ofUypVysZMwnniM456Udid0lA4TYOsuYrnrLogjcz/pYq5rpVfU7wEz
k18rAsAJVh9nqeyCh+BZyaRi4pZsumvpI/41VvmYuo+0/7juqTNGTxjXPXfm
RK0yb+ZK9YyyiZ8qx7DuPWed55c9J57HljMd3WkfgP4K9k1KJ7RGiiqEb/Pw
VRuS+PtHYxrBA7D7Xxhp1uutzAxocEzRht4yvM+dVGG1rV4n+VjK68SmSI/K
HNLHKR/nyT7wbznGcA0V4LdE58DyUhjCsFC5qagrV4xKHf91h2ioZ4sCbW3k
a4w5BN96fox9u3AO8TFdqfCk0Pg2oultB3KV9/n0DmTI42FKCparFLsmFKKq
n46EKXzgMGKUT9EASYy43mK2teXr8JbTI6BS5P0xRnSnL6/SAmSeJ0K+/uHg
/YXzojp4hTjeB2yCwZpUxDM9SHxPBHoGkxIbosXPAncab1ybSB2AKB4Jh4Rm
YMNG34dBrPVb+HudvZGjdKsHKW5dJzz8yWFsHYplZQFjnTzVLkNOaemm7YD0
A1UzRT7HwzYJHrtPr7kQUFWDXjELUe/2KEXo/ZaoUPjYgJHPfraFTXAPh6CK
Ga6c8uHgkcRbHIyUmbPZAehQTYzQSDH9sszZqwnjY8ighYuPhAIUjACDWZW+
ztkximdt1JNFtj04kWEZzqx+ZxP4TWYO/8W4/RowtEGmQYCXOx5AjM32UKyi
jjGZy0FhPnNzzvWsTJAhGREYmy65soIAdlvaG1lbzxk2FNK6xFbGe7W1NifG
329EU++BN1Z/i2ADz3/jA9IlP0m9lDmY2ahhZ5JbYTV0jvvAfm/bZT4GWDum
WbRigjeT1dJ5TBnUpmPE3BuvNsHeuCYRbp8agvAdvlYGjPPZlBWgiU6Q/ecd
mXzUsC9tAtAdlOlykBgWIVqFO21I/FqsAuvW+ZlEv2PjBzsSG8ow/tTyk57r
2jVhSNPrqA9Wa6vy7HydLwucIVXNic2DNqGEpZHv/1ohWg/fLZShP/0imE9Y
ZIICFfYhdfGAEl01DpogG6ohk1B1lMoBWmlnW+UrtL5gqslxSMKZv+Ix7GVo
uWmnqVlb0qOzQqpRZSMH7byUGuZJaPxXLkNbk0runGLSeRVCzwD/6y8d1Vhy
XR9mkczrYS7gO9pCn6ME7gyeUUQitm+tKxKUfwHkEk46CeGvJZ53QzmY20rO
6AqhtxPwDV4uk8VhPKla0IqHtvxDaFFen8/thMrVaN3DsODJMSf7FqwLkgOT
b5c7vbqBY1Ne17NzfjXnYu74quqYe2GH0t7dkq42CFNrWCZj5ijQBHn0Q8fD
wFZc5k7jaLnLiFqdXNK2gStidfj0z/afsJ0ki9oGw4zv3zEnB4DnvpkMvfvq
KkNyhktVZPKP1K4Bobfq1VmI+JEJugXXR9n2xasSVKPBIg6BkVCwimJdE8Uh
lQvEcOMBUwcpEnfw+ABWYT4g/tM4wzw3mCXIzhq3I/blfW7kab7QwmnqVxB/
cX2uIeMiy9AExhJOe3GkPkgeN5CElNyi8z6ZcyhdcO+1Zvh/FlLFXu0XAW2C
j6qSCeMNbVFDkqn2FmiyCh64fM+NN9TqCuufMApZcCmOB2j4V6FsrhceY6X1
EWPZnbxXUPe0YNHGGLMsBaB/9T/+fmt+vQsms3hnd/NHW0a/vMDH2PAWJ6j+
0XTBY0vNq9yMACfwDvvhoVyXi33xGqtzrFg5QI0Lzv51W1P8MHO9BKpjb8x/
j2vWhtEHzyOfOn5qI2gbb9CB+AOXNK8r7j30brGTVuqdz41X/bosxXZ44/KV
UO3FTyjfxVWiGVNg5JHTFovyPT0u8hA/L14Pg2zY6QKn/xJuuK1l+VHV9C+l
xCajQI5Rhuhdc/Hy6h98ufwbORIWWKyOQql/+Gdem0k2BbzZ8VkueCRWtsa9
uyAIilnHtpl5j8q8zp/WnNSSBujKYb4vMNMQQ4m+MY/S4/lix5UBK9DQMjKE
WAt72oeAJSeOO8INNISYrGwPb8tVaTn5VQjLSANBp35NBARzwVdGuR+Z5/16
Xd5FGdIFk6P3HYvWtCfwad6SkC5u11BRpZpNRLxsDTGRJgcDqe8tyI7FJwY3
3/4vwn1xL/wzc5/M12KLVsXytGI5dz+nGH5mhMj9DxO0m8jKsB+rCkkohPbD
RQNNIqJb0q/yXez6iUzjbI8DHlkcN3H2avHUFQUdm2nYdh0vbACS2lIDwQ+b
HJ5RqDXHho7dzAqxUOFjjwqU2N/kX2Pb/9wvkDR9nxz6Ut54Br1CBJ9mFJj4
tpV52trerefTuWcJM8hpgIFMYbVmAH60nG+KvgZ3A9xBXt/MZPKgs8ZdSizV
sGkWUyvOPi7KgTBWT0/ioe1kFxAEfrqNDg3aY8uU1XYcafcNc50CtFDAY4e2
teeLg46gMbMqBoi4bzuObE5efy8L2+wy1RtvIgU0Y9XAwydt48X12XoOr2mw
cfOWTMrEe/HcQBPxlKctWM26LUBNZBdOHPLMeeVCrS5TnF/SRtdkYOKCUUks
iJ/I8mcwlIXVnnE7xtgo75pAAKGQCeGmEn/jYCze0RL/KDvZfnbUsRzSd5LL
oHYBnOMhLTCa3Op4Tzcxx9p2Dc22mQYa+G/O/ySBJlYdPqsLp+7/biD/P8H5
S5Hu9v/5qOrEjv+hLp+nMaaiuDvOGBppGFoL9hjpPP3D43imd1dL3YBBaQfG
mSmOnHMLfPkWGoDupYkxr6yTHVqOI4jU4xvccPoMaahNgek/dErQHAMh5D33
6u6zyMMWCGL2sC/lY/gSxQ3VZ5Kgi3uiedv4UDKkryX2HCKnyo73d9bW9xM0
xj2Hyfk6BK3AOBrcKPUONtLXVJsUspbFejiQUptsPmtAlgfXQJflVkrYLWYT
BU04fbeRSMeMdirfpXzyrhEhKxfpejll0PMOW7/1pFEeIFwhdOrc5Kp4hPLR
BzS1CbC7O+Kw8+WIhL3CrWfG2sh5e6NobJ+yhpfSzFx51eA0WDKlrRHUgIU6
PWCmSKsfzb9GXgnv2xQ3ocQqvCZk4QCnxXVa/lzrfVnXib1WGy8Y1LnO3S/8
MIHIgv2WfgfZNVmT+IyxuKue0NwuK9Dccpc9ubbdziBzDkn/L12XggqdwlIa
ALKS+jOd59bzFls41YTYKoe+2FeG+0OfZBHvCOGsMZ+ooyVcQiIJCXSC5+id
E2U6R5hOA1hoIuj9v7juDhTyyOEFVDb55SlcPX6HYx/dqId7qBrU+zops7kI
6BYCdMVNb9r4OM10KqWGNn1EgQ/bnglTM/3XWf5BIpA0b+1jlxLEn5OdvRzr
XBOqQDwniIS3AA8N94Wvhas1ifZl+kfXPE/OFWIplYFdc+zmd/aE1TA/vnGN
r3Fy3f33vmNs1mHGZNdCrTknDKEo7SpEdCEeOF4G+laYRAiHKH6vA7/Qs4+l
x660jzy62PG80q04iZskH8O8O/Ve5ED7LmmYNnEsZCRoQR5PDC6c48MC53eW
AXL5+DuUcWOilK7O/Ozz8QXp3PfW+yqBOaYV66Y7PFGJiiBoY/2kCnCxAWvC
V36R+iKd7yy0J7GoOwFf/fJTpqLalgj+jKMe5ttgM46iBaU6YNzFFfX0kcEn
LuaOJqJOUTdMWLUrIZUEzjb49u+qdcMd58KiPbPDqlUdCQIS67LR8s+h95aN
CRHKbsHGc2l6Z9hKl5j3CMuaBLODai70JwczGL7hFhKGUxzIPiD0dymfbcIV
n6RBnZs8SsYuSp5NRNhwA86h6tIvuBTYxbhh3GBfB0ybfxRww+sBhPjZgy8E
gK6RF9h1SQ2Bt1WsBYYYWgIvcKI05lOH6NtC12q6uGMf7XPzTggX/H+Fp/kN
5fIXrcVcr92+PbvKYbl9Az+a6c5tsXnyjlU33aRME9hx1Npg3gu5nqa+oqMF
eV67bPd35CoAvXaq1ZRRnkMagQFLPXCL0UTSmAlsxSIXiG24kVXYS90fUgqu
XAQnI90A5LwKFZaxKd+Zv05BKVeBx6pCsDqZCmlqlLqBCrg+W3EMii6qVJGp
R1LbFuLi08h3CIC0JGFBWUqPe2+uyHr6KFL2T7TW3s3zHrV1lViiFn+NvYfN
ALcpyJqPyQYnWpqo9rEIELZA29WNOkRCEOhst7NXG17DEy04yh3vyeRIDaS/
9H4obx6KLrVONe4e92K2NuJW9j+2pjG0ZqW2xtF9Zo9+EEi5uM3F813ig0B6
cl+8MhaV0twXv9Pyz0RR0A4t8rvPRMryYtgPVjJfGfxrKVI3wZySXxpp1Pzy
5GPQL8GSJixPd0iSIhn3jR1NZF7F01tYC0HR/0+fgyyEHPo8ptxGcNtvLcJx
IdedcGhDTBjiDrqbI7tzNs69cc5zULEkWqLXF60bLshBiueGAdbJ3ZlpskTO
z+awVVmbCefRN2sn4pSEmOorHaN83RhIZw72cBR1J3vibIDV2g5KS2t0JroA
vgXSY5LLAnK1HAaTqjcJu/d0dU6qbKUn15cCU6notJ9riVUCCUDtgRReKwfS
uziFtfsYyQGkxEOEThaag3J+ABvATDwO8J+21SgZAQCuCUXrZhNCT5mflsr6
pmXzdvwKZ70rmMSzR5e84dylK+d+vTtuYBk/ed5Ah6d1OWN/lOUJ71n2T9s1
7BWrFHHlUq87+fWMYJTN6i4aJEasZNwVbvbB90jnEiouqIC6Xiv6Vzjn8fVs
cZdq9BeYfYJg1TMMSCB2/LqugabS6BPYFBA4pQH+ELYk6bLeqb4xaGsoKoXh
Xi19D6Dkm0rV4BCJjMmo1DaKAyId1bDHhNrLmsxRlgm7Zpv2ZhC8V9X6LD0T
V4oE4OQjjF8EdFUKlnFn9XHDh1gesGdzjfOTwBM2l1ZMVGDkLOYYct5e3Qwn
itaitkSjplJodhlJW51sudnBKeGRlDaG2cGjtK+mQkcNQTtQIQEUc3jbtwXg
/+m9+ERd47Jp/nijAUJyWAc2ukLVUo6j44WkyE+2Jl9YtncJyhVehsrXm4+q
Zu8fIb4fMkhfAoM4PQjf/8/k1BoNC3mvPrGK4VJsP6PWH6276sdW8FbWKsr0
XSxb1/GtZsQDoGxgEk4Zt/e2w4FV6O/E+h1nTP0Uf43J61AsHkeBWAtyMK8Z
popSw77FSRNe+nMacp0m6fNAQUWfdwD/Htnk1NzjBn9cm7kjbOGr3TgirXy+
s+Ut+QmFRhNLKYX976GTFAoRjjhmFOokWXysRo3F6QRwZuw6YGz7AM8p5AQf
7uCBrmLNqEiTwDZ50+aiZugDwgISBLSbGy2OsP7gY2EB5UPDYSyJB5EgkAdH
kw0Z2hOUvAy0M82nEPlJidvRc10kI+OBRmTI6wUN9zqsmDB72R/WTDZsW8Pp
BDcZIRIZRyZ+B1Bzcz8ysgUUE5Whnk+cC0JU+OX4Oj+hpRRwiyQscUcKSmv6
Y1mdTd5hI6ub7zjTG+umCPFtmnRf+4E/aa+ste8frKS9NmG1w3EtU0Cvb1F1
UVlc2+Q2WppGNr5dQiBvkY+s3Kmh/k5VQRz5QG3xlStyhZ3XS7vUKN0pZJjS
fHes7BWAXLjHDQwgoocGWJhyWjRfpk90z2I41XrFkuoZcbdJ70qPy48P5khv
KA4tEl/4y05MjLJYVdi0YJRt1nG57LEz/8IsJs32/IYIT5mg8fT1kkMtkKFN
u4GyMHTcZ2Jns5PXeGifEmM0S9YkPcb8VE+dklg/+2vsQxJjkQlSm0aMSu0w
jM7vE7VRGYdaCH53Scdq4EPfUcl/1NWbGxbdnctuGvvet91+3gEFqfGkwLsW
xjCLw3NlUqw3zavIdC+bVHZrzXgasD8tUP5IdN4MoLni1n/Yw+9Lj5skrNr4
8AWf334NUwJxyZaFrhaJ0bSYsR+Y6qqIMXDrRBcUgwqW2N5ULCGvxQvLzWC+
nITWIMQKWfKTacK69BUWRBHlwu1D6uprbDzzA1nQX3ptSva4r72/rKCBhuRQ
O2JfxHoF2pzZuzm9Ua8MzT+q1Mdvt00sOjgxgb8+kQzfPPU+D4Vq5EYTvpql
xQqtQmLVzRBa9M1M3zeYiNkpvPUFzDfIJxT5ePAusnOSfWUxWAoHbTnHmZLz
j/ROIPNgqBpqu31uYEtYiqG0Zgps1VqRWXRxNqQwa++D/trlWrvG6c8syxfg
vwiup4qPIT/hkvxM5BlKGc0shj1XRFIugnXhJOUplDmztAOldmJIHdutQVkA
F3ex0xnf+lwtsViTxg58DTBseGao6p8IPV/XZT9LmikL3MtAandoUeqFFdy9
Wdag6ko2xDu9XfBqPYcO7sH1xoNM3ZU4CynaNIzl3g8+uyoWASxin93MmIeG
2DB+H8uUgYqtYuyDB9kmwAH3Om0ZnZO/BEQRgBqXz5shXHWfcXvq2ptoz4am
rSUBXfXapTeOpCSSTNM7qJsXSdHeIreDFYWHDyKWb3K14+Ieechth9no8G4R
Tr4JoPWNFvCY9QYEpkRRHJkraNRofyN1c6mekhFIKVjcc3Kwut4JSzwkCIka
9lCnrtMt8wyFQrfrA9pkStbhB9EK+j8TBwdq6006TooHQwdE9P188hast/t6
gfOa5ZlrTpwoL8q7CfVVtYpUV+3EyvNpuD9HNZtk51a/nCDTl15ns5lz6zk/
4XhLuKhrcQA8X9ggM/aDn5/YCcLSFt2hdGeLJso8CCfhtNqo82wNldhoMBfe
EqsAj/Z49X5fEmIquwZr2K1Q6xY7gpOURixAafq0UCAHixdLebIlYA2hO4eY
vj+N8T5A6Bg4Wr/XDcMKJ3B/qriz+eujIjiwTpUCJfrJ5hKJVT/OZOByM2CK
FmLiowI46FNreH6WHka1mAZr+hXmyx71YB5d3q2GzaRK2ijxOWV1eXoSsK16
QRDaHIUWkC8xDPzislAjAgQw5vBoanRnocF/tqInop8snfUFokzC/GUvGmRe
o1FqIrA0BMJmtadk1H4V8hjSEDIfvns3o63deuvGmLRbIMLNK/pOjX8/7Vcf
vVCRpb7IsKCb+H9UNh9k4XUqM2oFXL6iNAIxWvs3MSeRg3TqI/qH8+oFm+qz
xWTjTCym5JZR5S/JYbwKuLln4FkyCN5FTgw0f24n7lwOzyUF1+RAxVkRVAbt
SFUDr/bGWND88THSlMQ2Y9ZzsJjr7SDB9P4QOl1ucmyd6e1HNvb8X8rAbIKB
I2fGDwzH6zLJ5A+/rIwyR/Wovr0S7On1ST7cjYMGkWOMx9BZ0pRrtJHibl8t
JwfGqUXUjh0zphHEalLOdZmYFb3bKeQkYHMOsL6M9bkBTgycJfCepbmx3/Nn
f+h4GE/3C/ts/3EZPC+DziY3nDGAinoB/QEmTwk9wfLREAuQSqMB9Cu8KJha
h/J9lmz15RTbPLRqROnVP3vwB3aB7b8qe9tIy/FRzhAZ9Fm2JfXqECY34bXU
Pn1CipTNZjXImKr7R0nGiQeAiGmdB4xDHpTK5MUxgH1TL9OHPgwlFJRKPfNy
JyndTFXVqKw6i/EOwxnSNCq9FMJynxdZI6BvqK2pNinpxhwjJQtBSkAH2yWW
9nawtlFDFc/1jt+06PoZBOCicDXsqLRQ/UuG8/YGMvkYt3nOFYBtHTmI8Xv3
Myy4cBYoEVp4+F1CprijZTPzJI8f7XawxtnaRjgmcSAL+Fp5YqKtWKbSwFTw
7ZxCKCW6ui/APR7+MBdQIV0KjnvpOCtV6SooSCvxVIUAbUYMQVLYyiSh2YRt
4pnyCi49lr5llhqMoS+6idaHo/I0G20IilS0mPfNEv3j2tL2iMeUfBy+JF+d
Eet8JVnnO6WFcJMDzr5BwFOWITFzHEsQqRq5SHDGPP6glOidjiro7qJZB7p5
hy6KsWpoHIE1C9AeCx3x/5aSQ9sPdL+LKPxt/vBRj4axTa8gtVvVFFWjAY3h
zZi0MQ/pqTSRXCOXeUvqsuR7b46v6XaHTc/qTl+inD6rJU5jkiuLr1K1piLe
9scvoH/WRA8FCVtMvO2PCkdKndWFj+RCROyW/qkBVfVmSlWCkVHp6y9qUiKQ
ztWC2op5IJCvhuGDblZuKoFFrtTm2ev0E3yozOTFOi01dWAAnR/NkPHnMlxn
5LC+cpUaoIYWnry4Ov21d0l/VszbY3TH9Pfd1lBdkYwAMG94HzzXL5Aa68wd
n3mK57S2DPlWPZ68Ir2UE6ejyYtPq2SRXn+SdDeOR25dxv6979psdJGH5C9P
mM1t0dIkVFR/LTPBmhehXSKX98r0I/vZtUsEsifpRxn6cJVijud5GTneJvi3
e1C3b8r4Y9nBDYDXQXMMJbsFtQgVKEm8SbGCaznIgZOgFna4GmM1Pc/v4UJo
rvry0Y+Haq0MFILBFhuQgo8vkW3WhpPkL49TCAl6RCtmXNV+tTC12IlvIHIN
tAwqYwEW1MQkttc308ap0jOOJ1+v5BfR5QALzD2QX1jGldOjRs/pLalIgaQ9
4wEQWYmQOYQjgi9I5531cMXN8QwDbGGJGDYxvKBDyDSAht0xZ4XQqxWf1UTe
yb2SPBSPunbhFuKfpG29wQy84IOzXwAoO8S8/Vbq6f+Xiefhu8OkWEr++d7X
SevQsj9yw+jsST27ae39u9IaEHQQgdgMGUGU8ZYGy15YuhBVRLJbrETQtw+t
pJHBicGO7X4TBBK9yXWQTeTfPlcUDUDmuqyfM7qOt+F4daEsXt2xC561eYEP
9HKdiNas/pCeVFwk0gmiU1guLCQIzVeFyRblloFgey2bbp4Xq8M0FvurDvi4
SfmyOUbao47/nQZAD+wrI35j3LJmC6me2Kj4j2viRfUJweMjE3Z0o8cPwTzO
kQkKO7hIlZrcb01V0i/3R0m8vH+AxOp84JESqk/K5Zx/X1E3QIcNei5RvUPI
K+4UpEPx3NJnpvXOna0cSAmO4sxnjBn3eQvl84sTc/WW/ANXYuvtviY9WS94
q9iHM/Cp2IoYJ0SnJqI+UoI38R0E3A5769xe1jPpzpua344hbN7kf1n3lR4p
st/y0xsgbk5eNUP5+Vt8UCKxRpQFLCRP7zBFsg7p1o9Hqd3KooVFGbADJx4a
rYatWzb5nvaU0kutZ9BhK2RgHqS/Og7tPuvrMgRK6LqNyEZS++xYnJIDBVbZ
vTNXNg7NUGgs0c1HqmrU7DssIYrMrAf5cpq4styuxa2V8ba9BHC5kR5OGzIl
jQ3xKra9p/b+5MSO0nPJTjdU5r2YlM1we54vcprqA2OhOhtl2iLxieLbOL73
MiTYWJxaMjhYCrjVTqkqZa/DVMqGWzPoqLB7he0VbWzXfwk6RwegS2mYVrnQ
A2wnhw0MqMPD0unzOqpVScNu1SUMM8cnXqevPwZzQv84pYhUFvdYBQx41tKw
Ez0DKoefetzc7TmDf8m8wLPLxsyD1Mul81PMm0Dvt2yYuLB1/3Vu5niNDq5O
n/EgYH8AaOLTASwpM/3fPeH0bMRUeE2Tb5WCCVmuSwW7wDT02VxObdT1+/dB
PHMn20YxsqycHl+IvoJkh1VrI3P59lGTu66qd3QyhlcwdOrRdKrlmNJqF0pj
29WuScooTIpAD8yYhAVcthoapnLrOjH+Gt1Tn8fOa7kCL4cJDxAuqiKZlzOO
DfGl0607HNsSSCfuCGbeEFPMVTpNj+d8LHuZT7HJPmd4s4zpwG43Zg9g8n9Q
rtJ3rtbywy1/YEs9AERKtqMjzhTz3+4esBb8DcjHa5aXzv6AILUsDKDo2mCT
7yPMbYJmLNHfTDeMXonU5UmlnA58qq4RTqwr/LT1RfAxAQ0mkczhGe8HR1c/
L8RkIL2SK88JBP2tKyGoqhvWLRgieHVoTzrbM7voNR3zeg0km/Rvc7Qmnb3K
tXlL8kpl3i/VZAAZBIOqjjZnzcOONxDN0vAk6O6nAn7oY8sFnJp2uelieyjh
UFXOcwJxNNeoKYE+YHlS3KdhJZ4no1xcN4ht2bIvexJsTwFSGZ9Ddk1IRnv2
Q2Nd1t9UI+6xIFo9Q4nw3ZwCsMMDfGCBBZI0zNFcX9/E4FEEeP20hLE0/kHm
ixx2GoDaa1ReLCYTkguhtqniD+wtvwcJrfavki0XGoVa7NeI+cqwWteNWuBg
/ucOC7BMu+Q+u0g++mVGI9waXFWwJHzoyawetAqfC2vYMH0PnS4l82W+hsQ+
w9nWYUgpJnnl7KliS3NBMFUOeBAZ5bbsxfZOoh5/B8y1fZvk546OJqBGQf+u
T6GURUfmpw+iQRslbn9ACSXP1arHyv3azo/MlR364TYVy6fS61oVHV/wf2rD
v43Yui8OeUd0FL+3DmkdURQvCZDGCHx7V4AiPmFjBYv8T1c0lNwkhvX70y+h
y26+PooGMHl0yJiAgoyXcIf0eoxncnNbfeg/jYwtsfm9ug8Hrk5AUwIwDqp8
3YPqxby88SsA5Le5UaEiA6K1qQb4tl1aOTKqUjeHrpkpwZn7UOYfQWr0YhGv
l4djWzRLibpS1ONm8mn5axlJeqxoUrdmC2a5z7kgE3+nMNBvaaVFaEhkigVt
teZz4HrBVnG8kfi5H6EjKXDsuS9EWfrvjO74v5qRFtxrcNSkbAJOS3jWGkap
NsFJmW2+l1GC/e2BNiMEMwoD6MeYGs9saSVhEO7/wYPHFHwRFzjtO4udfiyo
xA/P1kZEOPCCzmDlUc6nwn3+wml8T8SNdFrKzDBv7YAw1T++ZLtQm21Sajb0
weXiSmXhk38zUlFUPjiinmwIiau4KrcOeuuCyajeOW978yy+x15NLn5yI7DA
ZNYU0ZZJJ08uoY88eITS7YbwFz43V+8pIAaCxIXQKwLVS0tsSAlblPvwkyhs
PzZoHnJft6Ru9r/8PtqEoxW6+JwpqYIzhf8ddz+Ru95oSfVDrn2K7Ek2Qtt0
cz63r1OLT+5AnTSIsEDTKUUzRRXgiBsYS4CCGClVvjsxt+de4T96CR4kq9kc
6sJ7tIfbQ9sloYMpf7yhjQcReloiCRiSfrSmrSdMDASPPgPec8WFZhALOpus
8nXtHtttr/LtElbC9Gu5BC53jWm9LXU8T8GfdsFHxoYTp/nCV89F47emc3xK
XivQ+6YdVmBkxg3zFihvgsVM/WpxdlEqSdqkagup0ElinuOjlMpENeLIi9qx
t15IDkWxFi5/nxI4dMRV4TzEynwC7/HUxRcAeCAUNAJvj1OdG8B69nmxcnrv
7i+iqYA/m/jc+VKIx203N9PG4dFghpZneDRDukZuidHcBAVd7JoDktA7AqGU
rxZRyrJH9jJvpuS3DhBtR+kQcUq2ELVj7NYx3v1pd1qxg7L8RNDaM2hxBGfl
FY0TqQSjFi0Xy+rEY7yvjqmobp6iNn/drLGUFYshu2dS1wdkUpuejrpL4ZYp
Tx0gD+UmayNuv5ZTfcn9GnVcMZKdW51kEbrqXO8xE+SPXE4FD7270aKv5V+z
wHZG+USRwb8zc0xR003YOGcfS2SEZSZEB5V2i8PC/gjRWZYou3Vb6eRBsoqp
pIM7abJC/wR8CyTSaQvmoZVb5fXoYSpmDTk67B0a07TmI2uroFYHotFIijvF
K5INGIfY1wXpA+OLeLq0FENauK/6/QpxuGeshSZ6U8MSWuLZOJiTM5hT2XDV
6SSuTwGcZ4fZjCzPOEhz4GSRE8GWbkBImX5gxmqxyXda7f6xQ6SS+YN/7VAx
TrBugJkCHUzGT4+UveDQ2fslmnqiIlRYiE01zHm5maoDdMF2OxKNcoTaw5Cx
Tvxka7tTOBJuiJT50xgCi2w3RzstB/UugEuTqiEU1Vha77tN2+lIcz/a3GX4
3FIJsg3suRtF7KOHNxcmOYn4/xyvHm4I/tweAU0q3icpDnX5xdPrSKjFcOdy
6Zw2Gx4WEnAO7a8DKnWWWmbPxpkFm774qyQuHqXIeu9prC4cYDubJcxSJ6U6
wWriHkMCUMaR1EyAg+QqMxXII9WQPVLOopQWWg6yZVPHQ4JQHOvTazdI1pgS
BJxEVCp0Jkv7b0FWbnU6PMdeqO1QqjsDJi/dXphP5MeAIWp+5ZaIuxG5GRfx
gKABADoYd2GoxKxKYuqfJmfo80N2SS20oWoFU/6Bx1hRu3UImNlk09sLOwhe
W0gPu5TkmfbvYJHwuBTGlsFkYK1SWU8LRd3WRiFk0Zcw+Ffn/Oc/3jdkq85L
1J7rbfSWtr2pDchbrPj20zDRGNcEkBLojx1iVgQ1VJaU2GEqgmh/DgxyQar6
uF1AcOhJb8pSSt94x0Px6BeaqvbTpW7i2x4y5D/3F0FRxpz4IIFnRpHTOsng
58BjDJTCwbB9YxiElQ3wAm8SEIdUXVWgaSIj8xa71NUTNTd39Bz1YDtAjaYe
+acxd/k/ify/hc47GOO8DSVctfh+IxbW4gzy3TDmtWN7T42N0ec6CWnZqHeo
eC2u4CKbdc87i11AL6L1EutSOMvBLXRJIoqix+HW+j0TTaBZ7F26leB9zL5m
Cr/1jG09MaCW/n4ZfLerSBKqABYjxBxZSEWqNmwkGJtFtAb33Bx1xqUfQjMs
9v81tAJ1HFM2rosSVOd1+f/HC8Xm4digGJ+rgxr+VFahwuvdBGyQujhqbHMW
P5vjeIycUF6OyqIBrQRnbp2roHoOxtKZ/dLmT9yS+ac62MaUH76zGQZ37Yzm
9AG4905O0dypZ4zG7uVq4sbICrHDfZovgsWJuwW+E8LGPdrvO+844Tub1xp8
uknamck1ATeMYwtam4snTPRKbexavnSyLcbVjZns+ivlX720yjGULc3tQkcu
D6o7+z1cyFo910FpOYc9ko7z/qj22BU8uMLlYSuY5ZQkkvaa8dpDVvcUb99P
m41R4rSSqwiGS6KdReyUdaLpBTeCJPGDlt6bLZZkRWdj9f4NIkVbbgc8PwPh
QBGqPIKHq5+MWo5O+/R7iiR3iniH/DknRHQ1/1BIhFy8ThzFKdQ4ofr1zIfX
Ke/bsgOFWPmdEmLPNxlm3AG/uVDvcBvQE5CI3lYfDbOgBh6uolq8qGcmfaHF
9aPLl3LCmB2IiB23tvIEvjcKyJKi8MzHRCEhNgPqPuGhRxJ45ieJN5UmY70e
x0LbuLiQdGBnWCT7CO+0Q9gt8+hsOginax15KTARlfe/ss1P+Uw5fkqVNe12
f3XHI/gz/XyWD/6M292+bFy2YHMurbyw4ZNoNRxJT9jAzdXDwrlG5E5PzSym
ZyKDQwvdXUeEG4Z79mh41z+ZchEblImqVW3oXYE9atbEDjsaQGza0+qOSvca
Q5RK91rGG0cH1j8crUEF/Eur74MYl61hmCcRc8jJPaOOVthfa5GsrjnXcXHj
dXqXGj4cbGaR8H8qN9a4g+WaTNjzWltnXfP/ZOLIBIs4sL9/IR1Q1hp85y2F
h85JQb0V2HvV+uNTbTECwPn7rC29gTK4FyfcPPrA3NmHkqFE/2Ue791dL/iD
Zuu1Gk27erRZ9lCKTA6Po5A04qPXHhTrrJ/VoO1RPbnE4CoLzgsDLIebRoan
bN0UTA03E+dB5aY1hmJAHAxf07+aTvmVjYt/bUOgpHLAv6u5Y+fr5/TlV9p4
/Q8K8IlW9Agh/XviUZjdjmHVZMJl9lTbNQMVY9UYasSXmEiPzbCkaIkhfJXr
0MGlGYyFnJ3yS7bjDSDaRQhHitUCGdprPZAoTqE7NNocr5LtnYumtEWwaJ/E
BsQRBPgxbeH/r6D9ba9TvA3VabLmnKT1MPcsQYB8wQ5H4A19EwxjRFHv6/AT
ats4AYRnm1vW0ZwnTELYei3cXedDEiC9Pyzi57B/xnyDri+9EsH3qVK+kbPA
cMDstK7XkA2eNPwY/L93jBMYlEI8qj8yG6pzF6H/Udr+gWzfGaSe6tTd/aL4
ouKzG5LDqDrwpaFz5xWjFUOKFgbDpf7069x5J4XvycPUK9ZzgRJVYUmmhA8j
oXRIQnwGc/f/Hozfp++MwL9ZVAr2xGH7r20UmWZM8osarbnfBg5fCsBPjMvO
9U9GhQ5U5FBeQvF7hGNxZSc8o5IeWxeY+JlMY9bhV16ENX+ZncUgTwIHrHic
CBPzwkCdgz7vZKz+2r9WwknieaIW7iwBxWhr7p+U1thVptbY2GXiGOUWKVVL
KwPRMOa9uVfFB9rHTRNJjKBarNH/I5qOispKWZVPrm4iUlx1FlHsuY4m7dq+
rbnB70AS1ImlrtVYHHS7+hQ1F04FiOFLS+GAvAmEY7/Ar6ALRUJ43McHWzOB
DmUKs90w85JCJBSHryhyof1WAKIVEbWlQzFdL7Rtokav5mF4raaKDub6c9TG
RHSVsuGDhKSwJSlXeZMcOP9qFr7shwqMkohdRNfzqIhbop7LvFqY5Aef/Ix/
++gwZr7v/3RmEq12MWg685FmqiigT/hsZIp8dbWoUOhUqBES9rOzHY+0emSH
4YaRxZJWu8Nv83UbPN67yND/XzBksvyM2GzaGtQARRdch1ChMUUyUPDcW6tH
IlNv++f025Php9x0zk7DnH7igxR5RDQ2YEes6L5un7VCCevtXMpXVzmO+52+
N37BUpSxo8d3BbZUTtw1LOk/DFyYyt4VTLovPRyCPvZlCGJx3JKU2BiGSYsl
pOPW0ZC8jw7AGWcSXNfv5H1+PAhqvZbr6rQ08GZ4QJ54JuSATF07vxhCi+Sf
dmP2N5pOHxWVpJGrNH7fzgFKlq9RzJr867p7JOmsz1SeskzWKrGDdcuRkM75
QGkToPfPrqvnsVu9Gum9K+k4KDvPuGZ6ixB72jLyn4O6QHTbIt2sq/Dn4ppE
f8KzOx4Hckj4FlV/ssOylswot4EYMuNT+G6xCPo+nknIRwrrwRzM4jdBc3AZ
dSNIHQ0EzOdoQUtmHn2Cvvna6IhwBKG1kbcUdjh8K1YtqFCdFOOTj8phAy7B
lwC8w0Z/FTz8eW/gJNKeF1+VegnyVj5M6YUSJN2yS0sGAG6yKBoSPe5vuutR
TDYI+BxjX6oK3k/C3ANF1xn8f+PNaRMbHm8TNauTfLKT76xV+j3Gbfr83Uhx
bl79W9K840yneNrC7NfOBCjrSJocdYbWBW+ARSv57NTUVvzbimE4r1Ic6aKl
J2OkFRLbV4y/sFnJbHoQC+Zk1AMmDsYx37IJeDQvvBEgE6V6iqLZ558tiVOf
OqXcLCksrdGGuqRqPWyMGSyluMx8f+g8a22ZfBJD5FhPJmLbunpD7P74cCIj
y/wgnVrsQt7akbGHIi0h/ArKjmQRJpx5mwtqPVG+eVA4s5APSNcPNUub2Opw
I04X3GWgD8KHWQMNKmZoc/Pt4OckcoQL2z2LqeBNOT7HFKbkyLe/LiMHXjVU
CwIOND0rTX8eSZIg8SmCC/XG84q2NyfL6yg7eY640cFHI9w2Y7EZp8zoofKA
IuaXVq5hDz1N57E5bXG+Rl5gGOS1b0nrrlEKoLjsMWiMbrcCfam0Qy7/fFdF
jSQiAepCK3hpAKS1Cf/g/N81/WnImkrvKeThFqssHXFgMNaEGxp63QPA5W4r
OXcG3Sr28YlaYmCN7qnXlnxQE7Ex72Xe3pz22/cvTlz2Wd7Ns3hRTAsj5ACL
A4AUXw2ImhccOuZJYCyuPvh/Yhq9svx39r6QiT5Bx9kf9SbKOk3c65GyoikF
6FRGiUCAKjaU/AQ9RBjyet72Q5Yql434rSkAMrud7gmiabHcz7476tnbWFrQ
h5hAbLBN/yKnA4u4/OQpLik29AoRTlwjbVcbAQxNUZ5G8BYakUAE/O8ugmXW
6kEPfY1iBYbSKKBUKdDieb0ICUOMkkk+N59gPnEsJ2V4fetb3+UEZ2QK1KY2
5Xnyz6ATNWpOqaK7EW9ojBcwh/98plEmhhyEs9wJ/WEHEQaMnSoJpuwyB0fw
MmgGofL1dE8XQC+esOdEIXOOAMT37rjXIJJQXqkrr5OOAt08ubCdoiLyaBTL
u7o1pyW147NnPJu1eXn1S/k9cKtUzj6/TIsbIXAVooQ8aQokOL9Gio4zUVB+
gJcXSR46ueVJK/AZyiI95KOpKjiypAtnzlAt2GBi7r9ovN25ifIXVyAiDW2z
dT825ZGPJsAcqHnZj3vXWEF0vSStQ0IU2reQv7v7lzzM61ZdIcU88nUCGHBQ
36lm+qReHPa8IFlBLL6alRH/QZEf8AnxDn9WcxB0MDV/MwHHZX6BGfsImAyI
5gp3bjWKlAKW0ld9+Oy7D9K8VqTDv8bu7BRfkKWbkwXEzdj1511wEz2LcO4C
OHAo5pkAg+jLaATBJxjBMOMzxONmi9G/ZWOkj7+8ASdZK/n1luU7LOFpzmip
XvGm7WpRug1g+ULoxDCiYzhIrWxbNaQ/AKc2UcUTBiVDJeQw1D+YimzTgL4L
v1mPzehJeT+ilmQf8KkWJ9//h7YSQ4aKzgLod/ItIuv2p3cCCkvQ0YgCUCSF
22bPInoYCZ+4BW5lLEfeyH8d0dJZOA6GmAXFxPgOP6s70eq9XQ9XUmnV+6bs
RwoE5aSYIkMBgwkPzlKhwc+sErUwzSd+NauYdv/Nj7IOAV4Zz2ljNn7Udzr7
7eCfs1d3LW0GN5uJFzqy/ZLg1rEHz0JlP5SWsFFoCBH+TQYuu00bWniBF0JY
dP69Bo0ZGijZA84+4VTDAQRtfHVouxGYM2U93MPAaz8LXStA4q7JIi+4DoHY
fw8/iQbd0LSU4Rz5TdfT0rVcWxcectiot9QvYNw6PpfIf9EFZquvrUWkPrbZ
Hdz6kEf8YCDQsDfoaq7+SPgLXSbMdbKfHZB3pObsPa8gG55Z0MBih7eh8lN8
zlE6qIXJcfL6bKKPq38CR/Nu1877xKtvTlAy2PJCUvjJeqWkdb8AjSX+2IN/
y5cSxoUcfKdZ7+BIh3eHPwkePZr0qrvDzExljtOqd3bS8Ls4GAwYCKPr6Ghw
BoQu039h+BYa94TpSXf/7bITKpA3zZd6+3Vk/qrhNSujFPG3zyCJn6fgXV5W
8l3ztdiANWU/yF1/cE11PmxhXTQZPgKz6BjbrT9TIc0LdaR9huqaeIaryKOy
bGDpHZYV4eToVeTBk993NpE03DZ3DVu4/Ickwl90QKkgP2sNzDgOOQRZk704
PbGSBjN71tKzboU1KePlildA64j/cnpKjiLcZErbnRoQ+0wdrJUmrgDRj/iF
uXZN1KD8KvgFb1YsOC5PN3EGoOAhZF9iP9R9A/dwM9Wxu7J7u7ejGtY2R8lY
9u4s2nkXjeZiXhNbi+OrlSkmN11KyUdKtZxvoQjP2nsRjmGkpcMoqFnr572W
D78DTPuVSCASynDmdRHvMiM8Qln4ZGpOPuRjFbmwd9p95BHpJx5RLGHEzbxz
hpeY7+TZD3vsbaZbQaxS5HnRozYF/F+GYTstiYRCumlGXz9jS5DBmD1fwn0e
NUvyRrK/t99knaa9IrnUDOMpUw8JtseNUDqJbebAWMySbZF+0xq18WmzF/Fr
tUh//rM0t7OS8MNxoefo3PXGNVhbYkIAOhfBZwWiXDtO7BEPypLv48wGDynR
eXJN9ZQxKzM3xJVqhWA0cJ4SQYDppG2surUUogQGZBQdWlQ+vkK78BSiTbS2
jranzJl71VetYOWLvBbmFimaI4hZsj7f+h4DfvdWUDsPDyMulxiFx19KTXDV
pH9nLvvqBL6sw6r70OPrPrcMI71chdScNOvoUEfx6x47ExXCtCckuKy3sSuY
6EdXMAZ988wzdhm8hQ6Zu9s64KomRw1cjvLlzoKqRsZ3dZlR67Zpk7FNyIRH
QOBnm3zvfAFNMNM2IjvwqqU5tAFaoS95J6EdnRCOxVSQRBZWsL2OD2Fu2/Ey
OpGbWYg91QWgON0waD7Gh+pc5za1yajB5j5JT5PDdDLm4Gx+1WfRohSAgR73
LjYKqTQwcg4qsPPDbw48j81IxXfVb2LkR45RQWbFAXvjaOfzfmMNFQuJ30LU
2NUd/mGqGm13Uq+HP5nmA96vyBJFjhWHCqvrI0V5Koc5YQHbcSYyz9SAX3yI
oNH2K7FCq2DPDJ44crZ+L0MRMMFMndtYHCSV+bHqNAmCYzlkpTr0/HwiiQvR
XJhGeNH6Cet4L09t8oXqjBl3npRtUHk+2HJiXtpvpJ6fpAhQWj6QSpvXWYg9
cWyjOnEg2KmJlONBdUQT0rPjZqTukMR6GXa9I934uWmucVfukmMg0Gg+cdUL
7jCK5AA7lhbPldAQNvqaUMG8OM6WW5HXkH8yELqFAyFtTBk6of4/roOHjMQq
0D4/nIMyAZAg+SDtI+UnwIEZpXSS08BC5WtzHJqBUMqSyIiUQhXuuAm/Xp8e
84vgMt5lexUCb+BQrXrmKfioa4+AY0x3lTaSU98jx5aKqkOFGsdB7/JJj0Ud
F5a8qYvsE9adgB5B8SBMNofKW/JSbQ9ldVj5fM073weX7HAeq4UZD/XTg1pQ
cOOv3ZkigjYLI5aT6Zwk5APtA4jeLPOLwSVtg2BliLoKFcc2T5afSbqZvjN4
Y1u/r8964ELzgM36Y5FdUmxgONKyyZy3LlCpIoQRK9VD0KHu1Gll85BP+Vw7
BZUazE47AwmYTYY22u9tfMPqL4wlm6S7ArabkrpmA/zPoJxtCNNbFC1X6fs1
BIRmbwXxj6q1cKyd9N9t7t+0AyFGX4UkBGT/DYq0MossRJ42dhfSsyJGtqUV
6PAthWEqLg4+uaaCgUbSWh67zwYo+qcHpruFUzno0qTFp4+Lhg7N1QpHMXDY
hfJW/iB+0CH9URtm9Z29gmVQqkYD9NScKJ4uJpIOEJ4v6383mDnBvxLYCxji
5yL8i5WaTD7c9Xy/RoffEqFT0jfZH8oH0XfoyMYCCNBhrtuAgWW8nKhvlJO0
UWzz4fSLazzovb0CdW8z8S0kys8CeyBzy1pTbGtbH/I4I1JqYAzbWMtTa4cs
athJ/UDXQ5XYDElUnKgd7lSoyENtSJ5CI+1oW3THhRH38NlX4McIBz26V80k
UDvmjIm53dNG0ljj+cK0lOECeWxKVi6Dr36CR9cqDId83rdWjXF9OLIoa3Zr
C+qdNYGqFNq9kHEH6NndwOI0WLdSZqBt/ppI1AekEuM7EaghylzI7lP5RoCB
n7luXn+bgZmlQjVFMV7g13d1QrWCDSSXArL7ZzqKYY5AnPSOGbsjLqseKnK5
nIiSa7xUTwp7e0G0DXQZIMGK4cDnIfs+mGnPBDIV5OasBjyNOijCkY1lmMFk
5b3OkqvFqTAEOKFhTEY5XluwjlJWFbwtuv8cSz9eOfzZarKBaIbomSPvxRWW
8dQVSjQbSCAA1dmYEvpyFeddLm8YKfvNq001H8OEcWeNMkL1ytoK9Xp0RCEn
eLLM/GMBrkuWMmuT2oG7cHv/qT/p9IsxF8xMdTDAqrW3wdji0ZKsQc+nZZqF
8cvYigx9TZkjihsbJFrw6q0sDwbz2y3qoQJiqudgkkchtf3hYJng8ZJ8+83h
5KsQo6jc0HDfvRBUCevBLiOujiuT5XItpYWwG2Gs+mFHShcZLHJV6mTdpKTG
FURfn9kcH5qiRx4GtkQyPcvymkmEFzs1tggWs27OrB22mhxiQcx3unMHITs/
kt2bhPmt9fo1/+4kIM4l+hBfDqinMFcBcxVVZbjnhW76FtKlNai3RCPFGq1O
RzHppK0gWS6b2qkRqiGxOAxeGhLkZ6tfJiUTFaIyonIWXM3ND9dDsUVCckyZ
SmefOPHPpPnqcTAMSHgNvogUJfpgVXqxNyS3iBM3hlA0Li//6oHSi+f0l/JX
UnZVcAmQQACHvl2hsLhyoIByn5fgLelMbznMhGOxavMl/hl81lQh1gA4tY0T
Cy931msczSgn/x/hfG9p8OxAR293BWt+w8y+RnsJiyidqxZ8PMm2YYppDZVo
zrxwretsVVokVK9csZ1qFoLGuaia2Hbohncs6Lb8g8BhU3WPmBqZEl8PGi4S
SqCgLna9mqJP87l2bb6c4XBjqtm/Pn5WYi7nrq5OPUKXJ04EdeaiwCNc+PFT
EN8BiK4JuqCb6oRdG0TAlQn1iYAc1N/VeDQvWdvjVUtf0tqdv0zr1auSSAKg
GHO1iYkELUp3Ztb33CV9QQ4RCHC+ph16DxJEPfn19Hb0cHIqiKwbNrc4FRaa
7OzTYdUOu/TvI39Tyc7OuOxd7xpmwaI/0woAgAZOnHfolFXeSxlJ1iMEhNkt
jBLq2P76qlVdshH9ltLMH87DrotPK2iN/y/qzU2Kyk9zCxZnqbpqxqUHq/4j
N00hh/XWT7S3FI0BPJTTKoZUb60yd3O7bw8Y/ROidx52yZPSCJQ1UQmHpeG9
CdcspuirZsuhx6fQyBuwRWXbZA/b8ifrTozgt9jXM+R1pAFbKq7tx8D7savp
yDLSYPZADP9Rr5D7ZilglMfNhILrGY16m0oF9N1ZNZxNCGuF9HOo6cJvO5jf
m5ctvuc+NQ1H8dcEIAiOkD5xwwASWZ5/IIjrILgOc7xWdL3clvbdW7dHr0xD
ffGS3WJkMCOclhUQNYVyl99mw4kd0PGJ+Z+fEfvSdZVI9S6ODlw3BYS7+abG
M0RuVWaEH357hwL2kVMeebnFkWQ1xd0PxtKwHy4S1hZs9AbEhU/MNOijRlWQ
mKyERW70DTdA2uVBAA87KfVCgLk9AIyE6eUcu82XM3fBmFMVdENi90Pf/rUH
nNowrGGVYg7VNUq+gGQxSQilv+RqokqAbKvNtTivK66JxMVFDMfT8RwVjcBU
97n9Pw+DIWbytrHvpsGz4AnqEJTcwxvxLXzDKvvTAIaShtgkHnP4y5p503aR
8c8Xf8VuZq/pZC1jDNzDlqGS23oNcGenrVOh1sCm8+56ier22DO3v0y0a8Eh
OWa8gpgBZQWN6MzSUgpnAr5VlZK0EtIq7zC8w1tMn9aNjg0jjyuBjqJtjVSB
JROjqRZc72Bmh51M/wsxkt+fetu5HcEssPjuqhKxq9x1ZpsTvbe4uWDYyA1T
2i2IfPIzHOcNL37UBrX/4fssm/VaqJfVoRkbNnGMXIX/9PdZKtCjY1Fm9eNK
L0+XGYJLDdO/vryFB89QcrJ/9guW6aXs1OUDV9AWalsG3IHOxZe1qGyjO+SQ
m3b3W4OnfzfJdtQjpYh+wR3sHGkYAIDlq6ViKxOAbChlz4yTX4XRiU40t0Mv
mTWEtXW0VEWe002oMezUAt1IErsycF6tWb3AsoAEnb5iUT0nzw+2IKC6g/FJ
+PrV4HHpm5IRJxL24r260HMyFCFUDPp4M3mYifK3TrmdKzafb45fXzL4DCwT
906mb+YVaJjU6ZF3zirhC0ZP/KTbHIodLbfqImm+/sccbJksl5ejD0ZBnVqr
4ayIDyUEBkfQ/yEc0I7+t79fDFM7nJ+DygruwGnPnzwRZnij0hOClyi+zeYw
kWaCCa/gq+I18+4FSs+tgstu3NRq1ZkbHeC7e+nxt81wh8lIn2LBDGIQCIR+
lVHiGw5syNnCjCuJdeWs+l5rPtjSARgaiYIJaXLKd8sJx5Z0Ov7+zzqjO7sK
fVHhnEg4j6E3Q5n+GOmrkvQp6aj0nqKnLegZZzNThSYxBBSvNRkRTKr/tuNE
7FvDGjfrHgQfIdcKP5p9V2GFZhm+DLEiL6bvBVvOqIsoF+hNt2Ba9coDs6a7
EmfxCcbAC6nUDv2Z2C9/tGL/gLNdRiZG0HVvlEh1QltOQHbEVJV8pqROqh4X
xZBR7O6PUEsvEKuSjKU5LEzMySKwWnPdgDqOruk6BTBG9Gop5ULX/3n0Z4sS
8ueG8Q6Jg7oCkMyxHa5NLkAjpEcrCfnME5iw91Xd4xYoMp3MtB2D7g0CpRjw
AD1RlMpkg+OxbIT8QaPprTbtkTjvjlKcyQ15rl3z3pwDOWEpavdkGJ6Nv1iU
ka1U8xghPR9ItN7zg6wyLE6tNFvPBQ1AzHGrGy0IGiq3Lgs40m9wFpWmbiYz
vLVldszfGrOsHjKuTcTQWHWa5GViYGBeFhTiQCwzjWw7+0S1J+gFkQDGCzsC
k4JQ30CUuRwoZrqSBo5KZbO7PTVGfPFMPudAcmLvZo4zC9utqOChg+Ayd7jn
a03af9fAy5p0VmsAxqKKiLDHiYxBYY6hkTTc5q6+zyZw1OdVujXvxgb/bbEn
lQegxKPXqr5hfNtcVQUDrRab+DA8op1q4teVVAvx1RhGLm1PvmUx3VFbADzP
bjIX2b2IAQrD6CE/LVm0ZdSrk1e+98Yu/HAqS4NsYp0bq9srmpqpVLRX+V9w
mEqNLDqnvTwXCss52N+AjE3X108nD3k70Syf+cLGbBjw60yzdoq52TVabcxb
vFN7Xa4RJuPUAWBo7IumZOcyUkwWC/ruGI98D/ENjF4Q2Xcr9tNR4NgP6Kk2
I1Rk20O97Sr+FNskSLv0itd2BtihQBEcKWYs0sTVStST2choJqFldOSH5q0g
rBJYwJWet8WVLLTZZ1rHdRROYI/7d8MFlGGN/V20lbpGWiW6Qh0lszJ+l4LH
eeLi1dU95zV3TEWqRclEvsrGPKFddt8ZIi72nybeKdZXRkUBILPNr2zv9NVW
R4q9vP4KwxSZM919cRTS8Q6e4qJ+Em7IgA/rL9PeK3LAXi21WJ0QdtzN/5DJ
xPbitrIikRPau4fJdpUbxvmiS+CHiG/v37F6KJVt5Snkt75mUY3wnl16lSCe
9zWgOaWKZQvxjJzdxZXIRcjF8ah3wy/2uhsv1bPhBSABr0HRcE6uML+BXT3+
47YeWa3YourOaqudy0L/TEOp4ZgNOy2enf9KZFQMNpMouNLkLjZw3yfWl1ad
foSwI3iR78u9ojbb7VoZAFFznHjMi6S4ZsjVUeLy586n4Qa8m2q6dykSOztW
iyJ2lVdtAe0hET9OAY8m839qFReXH+MUlXuhf9EpgH9AybP8qe6SeWhcbX2w
i74OhGrMPDb8aWDPDBUHWBlBY3kLYbSZLUDR7ePMQgchqoIVf3S6b0jL8/Cj
c8Lwah40yIFP4b1fbtkMm9vIMPaBbrQ3CcOYD7cc+nbkjoPaqNvIx7LVmK9l
rF9REfB/BDD7Q+0WlDUwwe83DI29To6VSMfATCK7Sj6ENcxR8aYrpdDEJgOG
RV5L8Vxv2RsJGUmAL197IPDF9wnTHhEmgDVcCWgEVmuprn6wEr3NPjVN2J9U
2QXoxbu0mabWXxDkIlrX4MUgqOkVpH8KOJOGkfHgkYQj4cZky5JnOhvhC5+J
n4jGz2FTUcU/990Elyj2KrSPNfCd2ffNaWj8p2bRQgksLUN2enZZnVO6GJ0X
N+1rSGksuXUR3bywbLbq1JW7otACYnZsdhmqWQeMNFt4Fn7mEjAgX04458rE
zsfaFZySLWflgYsPnGL2ZlfxBN4kKCMGNzebEzYuC2rTp2YoNYiANhYDd4yE
9eAK38PtRoFhXDiHnzBlS+PmT0S972IUrw3XHa9/IU9IS656J0oXNGKAZYWj
wyOc8ObA55kwX8+b62svM8nd9oCpcbucB7/JO7TNvoF6+Sxeh8ujxM0dJkrc
f/KeOFILGcrtdqDafFRGlzdiLnycphrFwfb0TJ0v3wAfb6E08nKq+Np7UEei
W53eKlPXpuDVeJX2zDVMpOxTE6z14ztNJvHIairV9RuwD5+oR+bh8dgs55Iz
TU450qgCOZuPt5XSaEMv+few5x9sInaWjrz3XqVXqUZeISBF9jh2yBpEN1yN
dYGu2+z/23J4Gl9UDMhkHDNtj+Q0lYg+DweeoMOcg8z1w6dtLSfwkPaJrG27
QmIZszgm/zJNp74QGRwLqsPk+Bac4T/7QV/OMMo+ZabSwA4NuR440BOkGekB
Vtqsu22Wl39YYF+ttpqxcuavXFoyQKt9aRGXZOAXBNaH19E20dPNljQChvt5
D2MB+xV2nsUeDpci0Tyhki78G6qD30ADEhGuH7d9f5oiyOQCZoc3wnItW8y7
fjgMr84gHA35YVhDUrtdrlqD8niqgU7oEORctMv2jnHWZTnMXyFJgRnQhnOx
moydvJloWhNccY5y59Cn0h2HJ7RkFYwCGksdZGsHuDXSSE4k4OuvTh7GbNHJ
VF7EML3u8z1a2/JiU0CTWMB5fdQS/KiIkrsnZxnu3f8LZEHQ8KlLU9cYXJex
2i4m3KNEEA+6lF8lCGMlMIrIclbGWEKLoVVuFhyhOamta/xeGEM9ZGUxJTBR
K+Hj0jV3/Sm25ZkMQsf1kuRQWqkN3F2oOAUkO/Bx3woEy4Q0keNbu46KWlJh
ruDn7DP1JtVPfAwwkBjcyIIfx624xtX337TbtixzFhYQxxb2wkaxao8ifVZz
StjTease1lu4ZT82+SZbJ0h+aHrYb9oTwR2oDMAcMleH5ffRnm1OmzDbJOsK
+q2HONWBBTcuw0x2OmxUTkVHXMy61j+EP8Z2Ffhu8rH5yqtkGLGEUJlhKvLi
BWtH7ct7wxt6G3utgVa62sBydSiTSS9wzHLcGDBV5olAv+0rA7XF9qKfUF+s
BvAQ0AKiZjI1QzXpWIzc1v0ll9vxSXs+IEkEAA+vBrAFR1AeBeMegt02O9+1
luqQ2Z9LOac62uOWpiXZLB0TVNCPFcRgnEZ4XCpAY/nAbHVTl1bbV4UViwxZ
tbelbiIgPrmDD2QEZCcwy3rGUF2mDPImZRKvLi98gM3oQnNskeauZhWuAtmM
eyIb13TnONEPgnjEiaTLJfZhWV5/Zc+HFmpAq7IIW08TgM6Xfyb9C9IdMPpG
v2DsBA75OQj4s4rLD3yCIT6sNvGVSPUiBZ49UM9RLagGp1PG2HJd+00GXQHl
X8/SfctbQmRJ3eOfWexCT9h1WK+nVHaLocLqbFBI+1XFzrOJ9gSBmm/IpJmB
/HPyIwRqVDlcVe/pK1PR/oe0aQ42azsz3N7sMNvpf+ZeW0qPWsi1okZ2k+5m
LCVdFOkB2r3ucxfHl7OFZtYvTGAmW6vImk+OLo10AvE1Hfbz0YgeY9gyrn+R
kxou/VkIZL6K+Z7NwpEaXeKAnHUfqOIMFu3BF2DAjm31qpPNNN6U1NbatlUV
LN01oIG2btNYtz5PNfmrC8bTDnoRsJzqLa3MIc/wkrvzsYFnfJ3xV/h6/wiK
riwnou0N9TbjqP+3CERy7WCNdCL3LB57tmdDykgb8M3QDGEXz8xnraNJZkra
M48j4ezc03vgNUdqOfGSC/he5rapiWuzjmfEfjWons2sqeKUEWI32R2nmv8x
iUVK/FuaGX9+tfjR/fAaAR8uboGUeIQYHlGXcftHmGaye4TGKarrL18hZBoZ
apn9U+1ZnsWV3mboUyiBF4IxY7m4gWMACewYElNB9/KipwzVAUK7jAP5z0aZ
6ungbsCkX8h/o/hjT1lLPQCixw8yLXaHW+Xgu/LqOEtuVkKiGKhVLTfB8/wJ
ci8Z1D0kRkMVVNS1E8NU0h3JIH4BfX6XypPeUYHBV2Hx6v1NDeEsDZyLbOWt
JSemDhDe0hqwpwSoH7FcIcMEwyKi58CHIKeUHfc+I5w5AxrY88SyePNQh6L8
GPeslBUMacADGQbMUh34ewiq2SZpad4JD6qeiNNKDqq9VGsX9HtKCwc/93Qk
MtYJZMIEuXM5fRYBJ0CFdT7lbC4QxK7bYnn2HvF1CJW5K4UqWksUR/oSBM3j
Cz9mnQl1gI9DcjdirR5l+3Prq6fG7aVXst7590JXeaKvOhgxJ+ARDbgI+1Aw
lgs8HzJYH+quJKaB6vU3oiTBASk13POKBQOhkqCBtnTk/jLz8h+bypVJCN+s
ExlAcj7bucHrDd5VxQpxvzL2u8V1Jp4+ohTv+1PavqrEqheEotrdvqIzMdhf
iR9FOKIbRPBS1/W7SNF17QcV6eRtGNlviHLuv2wO8ddrjNu60E9XCUZj+sJx
IRPkj7qz3VyYXqCJpnN4PnmvT8A5vbA4O10yIKdJr5pAg94b1ezTRQKWw0Rt
7hGpNXaUtC2MNHt7NZZpGN5CM4WlYeB5Byxpooppf9nmb9Gz4S3hNzdoKI5V
d2M2uhvqYyeoLV54DLOEEWYLpMb4jKJMQAl+c5WxcsuJd8Wa2DnhanFTSAQE
eYUP48+zikT6pLEkEJfIVCquR+2WB9Js8q4XgExlQ09s9E5qMGRtLF061VL5
VU59nxHepnsTW2BbaA/+vVTt/3nH+rG3b0Y71GoTyu/vDpr2ThipvLTzQlyg
fUYF8zepwAY/KRigZcmmtvwAaK5VfGh0UzWTgNauVWn5CVkXiMaHlVHtagKp
uWnJ6hOEhDCjcS8W0IesURneRpF5WmzfOXZF3CH3TPLchBXWH8v1jv28cv/k
bgUulbx4ITSuS8Uu5o6YiNQXdQ+CC4sYH060o5B3+H+IyACpLCVWSI9/X3o7
zDcirzaCFqQZrbB+R3iPdIdSrchut/nWN31h57RQOCmdJ9jDYWEAtXujKDUZ
7+9Ys83FoAKfoQnj2iO9OrfbX9eRJL+4dBgtr6OTNi6iNZ1Tr5Xhr/tGo+s0
Tjske5kmdQLNKpPhYGYwEjfU0a03xnsw3Ipaq5fbAxmECnJuiuhfs+ZE66yM
8Qkx7a0STt+gKP6YdTGTb3SSYwHUdE2sBZYHRU1FE7fn83CJoxLq3d6KuaY1
Qwll7bjX3UKdq6fvaduSWx/7DUxCB5e/c7a5tAAuV1eeA+8zIYms3pxAh8FZ
TKY9kXObDKkeNTLUUPU8TpyfH6j9SoyH/NW7DZA24rCm2bQHCUSO3DLhVMFo
4hTSWz6IHR+/UtHieHCsRdhj+z3rQCR2fqJt+UW3lYNqEQo96+6ya+zzj8NH
2MH1xak5jXRAKEy7A1JIyIv1+DxZ/G7ouzlPnrsf3SAcieaZ3AZlC4+wnDOZ
7mMQLzAMdPVWavxYxiQSGolp8kOyb4kIq0YhpJ6rQ0lR0zGcvFM3Kho+g0+z
3K2TjPef9yHQ+ey04VwL9K4QUhomTPfBoWZPhS/EzC7xz32HOXwVr4VNnIDY
WEZcjI7Nd9Ex+/2V646l8LIuI97wtKpp6KUS9FVxiq1jNOrhvFmAKYdvIpkG
Aw6U1YReIPDA8hqW/Zv3IT8EZONoNkm/KWLfMXoJzxYrLHQGjwffRdRxpimf
nZoX1scnb1C76Z6Ww15i6RFF4zhCBLYAifc1lfN1y7WrpM6+0Eev6JYBaNWe
0R8rJg12yZM9S1rFI9HFSIaRc3t8x1J4vSyoFbhND2b+s/QceHfXGEidk/cj
WBYVPR+b6DKYbwEPAtAVJQcPsv8HU5OJGvRlNlT8jxjhD/xw2Uu9uZMKYtqA
HD1L6aSTEj4R1rtPvGvcPzdujDSIhJ7rps17KxWYA8b7L1x5EXaVpjJtkqiU
iamKZe9Os9Zfej5O9KB2RMUkL9J0YBVBBYlP0sSQOrlcbAfppgwF5i6dPxIc
XDeis/LE7USDYcvE0Hk9oe4Qdxo4d+qdA6b0+gp14ESA7q29ftOAFYyWM/cH
l0Q3DhujrajGQEip8lrhbHKgZOBGrlf1WaPRaUog8+7/qMr56uwQjrUtLMMr
AY97ZJ4cFew5ioFOa9kY7xEiOkwWla/N4oSk05Yo2Ktrksrc2TnOiMauXlkP
xIoALvScfevDbLDkRya0Wd0iqNzq1W5EmXi7EEI+1zO6wiNpgG2YEWkCv5hd
39boIEjw8N11g3mHsABNpso5j1auQKsUENQ2242w57yoHK9BOaqz5X7yok0r
0oT4MvVISAdkmkWa4pilUyj5K3OIwNe1TVytZkvsn6BkrFFFBtcpHqZ4TBkT
yHPJ9h4BIzpvf3jG6rlLFdW0NwsaboP75HRUsL4y7XnEOu5rExtMF4RNATiG
5CB3hzal54UaI28LWeWIsQUgcqmz845tSL/jQT/OA7Y2anzjWX0Tyo0BqJ0m
BlHo76L6fjkDoz7TFAXL9kCaQK3zROqdWX/RsgBpvRYSmEjHYqcKUjC0dTxX
P4OSC47X1RnYRN6fk1TZfUmkMvfjxIjn98lLEg7GJu0eYHYle7gA+0zz4rNV
pH8tLEFUpf5Vp6gpo39m6ddNQfGyN0RzcSwOciwj9/eef69MKF8DlGB9Ftbw
w1nDLYvYfyfN/FGzROFyjQokHKg2awaT6xVcmeI6paUfjEedX3NL8szP1ecr
fiTgjHP0KLDNt+dBFmtNtA8Sxk5VJskwkCVmjtxO8Ur+PHkyYtaa4YpyzCed
0TbuxBxExCmjKmU7O1L9LifStvNG871qsTmal8VLuhsPgqf0d4J8jtGRHgkz
53kk/9kC2XjRqy/YG0C/zwJTLykRmv/Galf6V64VeCOhy1nqyLYbvCXdsZ1H
YxgPcuxQItF/NhitIPa1g+Qyxn+awqbM4LKYaNrU8UE/Ic5NCUpollSaGaK8
eLf9LP5360UT2tZKOIabkbTgp8ggejM4tlQ7s5/CDIbPY0GqW82cTEKAxIvs
fbHBx76ZSS7M/j84E4udQ1lSFFnvNO7zP/wu8FlszOniKjmR6u4/DaJhOUOb
1wCWcyT4iNKIBS+JS0xC5TEi0e1LDz8xVBC2xPtqUv0iOOzrZmSKK96EwY73
MVo+SjLWGWZTDOaqr8eyn9qX5+CBEPGaLSw5JQ/3FPuiYX6Hj7ujbIsawBBd
KbsktsIPKDpIKfZ958YRSu7tglbVW57Dgo56w9HK16qnn2lHpo+vnCQrOMxc
45Ej8lmcCczdfmCxOqK++PG3TSNxGtcUYwGHhcqAJgD/ZvNS/qFYz7b2CyGJ
+K3OKHq2nzLEX9WYKwMZa6cXAlPNaampq7uYV+afproVU9ZWlEqHAezziiUQ
RrAdRrEuTTR8tRGuCvjPgo1E4FhFG/R19sCT0SGY+AtfuP3Q17piFuy0Lg2q
CHU60SnQQDVrM+ERFww9HH6h7Y10S/zViOI0hITeo6OwX+hZwS33UGNpIEvd
p2sw75tpiidHEkEqclBont6FTEAPO7e8cUWNdDtnR7zLv5BnMjUzVvUAiSHq
Rx0dDM6nj0g7T4MzyN2h0yySxsVrlPHWBZhi7SWe3X12x0rpIVqbaYITjRQP
0grL2XjuTGbabwY25xBXV1jTZiDTIU8oUmsw8wIVxyCGY0C5HuRtlsJKW6zX
yION05abrMR7copKa1DXrpZQUWd4yfuC/w0XZL5jZSEAh4tceXNpuy9YaxGk
Wi6NlrSTh2EewORCfPHwfvNZsjiF1siChs7ZLPgDuiwWLS8KzApVbDa8qXZh
RE8RJ0U8T2XTus1aD+BOzl694X0j70/jUSZ+AkIrRHTYP2z5aPGlyYZLp9uX
truPsw09fjJxf6GWz0TStnRV4PN6n2xtWVflyOBhFYt+8Y+uuQxQd3LBWgkG
Kbv2gCs4S6dsCmyOaMvo2g8fwFJbTSegh0ytncbZ4zZdj4cKnLfNcWUcsiC3
7aWo8SOom2VIvrFlF3z2C9NMX+IYkE4oi0bNH/4vFwIAtej5gZRGoC8lFq6k
WlMkDcLbG3EnvMpAAekzbXTrhBwyM5Jg1NggccO6Mya1CUr++hxTBSkM85k3
FapJ4HVrxpvDoNNMHrTTJU4HyH3id5N9AWOoOtCNeHG8rrcKXpU8oX8f+mC5
YejTtFDA5X5WZ9T72wlrsgrLZ93IG6qiFb/seOeBVaFKitpUbDCvGwiCllej
5zu27M9ZYeWE7XrncEZqdjbVGefzMVskl9Dek4lQnwgQeFDW6+72WKaCZYeN
m51TM1tlqtUIc8dEtYZ0qDOoQV4ab65wqcBkpyJB8sZZ3apk5dvnGmvK/Vjn
u1vzZpRpYPBp8hu+Ry6QcDhFdTHRZMuVpsexSclxtG8qlBbyoeiL8v0q9sJ1
o7txvpWoHxA7Fe5jcHIuqYwCc13rHbL/M+xZoYvwvB3kEgA4flDnKocjW2tD
D6XJzGyHiELSxIBi8UOS5/rngfAdF2C7PwLQtDk5JL2suwyqkWYU7xCkysR0
7cSCwIozZ6yzSFjZMQ+X6e7IqCQM7c5nEPApedbk6Y9bWWNqiERvo2LP77LQ
r8G5cUPPZRLg/1GtRU/IUQ4vvXCzTEHfr7HBf/QfGAbpwp6BJaFuIOw9PYiu
ZUzn3mQ/aSg2ne7W5EaiAgzOaVHBwJ/mSXI/yf8NfCHhKzf/j92U13lwiIAq
dszqfBNTUNMnaDOCcgXbQEI4hH/7iQUhOv38MpYcXHnQ2GqRRgC3rVZzsbb7
22U18FZkoGpHQgOv8L/Gxy9oNFx+P0QlMXptBh0IoPK4F7R1x6AHIlqyZtiQ
mApcH/SyhyJlQynNEYKiwyg1XqqE9bJNLpzCvu9nLTMS7gqKajkXC5WEqUS6
vdTSJc5QbRi45A4WjrKgg2M3LsO7MLvbwBpMK312LHVDMsAnclunomVHSLck
g0TXe605d0BwWSLn+ioLjn2hlL5MQY9G+igbfg02f5ydVvQBeFiMIE82LpX1
68UxTODxinZhHnGzPx5ib0N5MpmohJewj9fL1aj0XhHO3TPvRK7UXul/GeTv
Fcu4e5LRnscPisZRLm3Vy4HPvcGb5C8iMkv2skewWbySHagM1aRNuFkSptXx
swuRquLlIXDhQJg60BLWB+M2lBcUFNAHx0s8JCCY4D6Sx2UpHo1Ls9Vf2Egw
SlPmxLmkj+uWFODQ0dPT2h1bw6Ff4UxdZ+lxi01LN4nPfX+6X0f9cmHQubJp
EMnt9qpHTbEqVwyvAcJu4L7eSP4sHaoHBa7/IZbHvc9RJ8EooYjCZ/Cs1HL/
8t46q5IV1E2/SC6RsCp+dXDHZVnPmu+6zgkJSbrXgHyQ+IV23kFj2W2oJx2r
b8e+c77Uw1qJoWm2DNuad+dzk1Zktq82ZtIAlqiB/oysAU3SOx1PgpaNmt0M
1iFUvezftTcRF4FW8Ub2N5bZGH0nImkvOwtt3X4YFAetk83wRSQI1/sOfyJh
p078FPeRn2z83Ew8xGwTVumXV3jjzcHoLM+bvzcWHxXMSiHjD5+ictp3pt2m
rYozTkyIEn+KFqthGOE2iybgHK4RYKYkKrjc2PjKhjxNfxgIX9I7EkHF1txu
VR/b4w5uR9pHXCioBh2LjQGwV5SYa1r2GPoA43I7FuOtOGZ+HznVc4H4qA+i
ZmXL1Aby4/MH98TMHS2OCsvjaqkoM96TdNKMQUOtsT1h1Gc2y+NHQZkxFojN
+aLyd8CqX9FEYrLjgU2gfnAVer0AkFOGhuVsuo6/Q1WTGrmxkx9oOpc45i8+
MQ5pyUN1dSrW6ppbZZ2WobTs7UOglOnieODavYqs5TmB2igL9njD+kg+nAgQ
/HsYn0R23chXrbtMfgaUGypZxFTn0Ku2uqVToDrefKq66ydcDpKv+KDaaQXD
lyziH2u6UsKgrcLOr7SXz1lDFYAiNIPfufLFAycn8h6K5PHlIO/qYSYFLWI1
zx6HfRxZqiDKjM++Ii94LFxOg89lr3bD76I9tID0BX+khtI2KDJkn7R11yth
oSEJezAQ0O3ke4Cj2K1Lj/KtZm0oL92JNsknMu/CD268eQHw03UxECf7Rkwe
zd02EfsWyRlNQYSMq7Mn/3S60JJO6VPkyj9i+BX78nMCVWhluoddGwo8Oi1p
7AlJYWIGhndRMvk66kYj0KLcLA0GZwy5KPDOV2d1FsBs9Od3BsPsFw03bJn+
ZdE7kb2bS71U6jIfPj9oScJUcJHDrowI3qJiYjtxgsPSJLnglbLlesDogivi
/B35FCKFf1eExKBrz70HRbMg7MKETaDwlPUOvs7/tQCb6SMdtK0TBbbAJ0+W
J0Z0rylLx8VNQpCmCHplrTpHdvQ/6tZzkLC7ZvQnw++/W2FKtIUBPNLDBza2
79KDRyI7r0bTyyRQxiCmRRFp/1q/sxGfLjIN+I5A+GusQhEMrHltNXJMF2pP
d5wq/ydysg1k+shuO4CdvMHvBmg+23lUROvn4oDG9m9W2JcHFpTTVPEhFMiI
b/p6k0XhJYgFTRVg7RZ5swWbzGhmTmfBB1hq/P9OdRVvaM/WIaXH9bRSlh3O
QmyCM8JYeweI88lv5VNIwWubXVf9TCSZxcNP23uWHaAtRJjbJnlEx4koeIjK
Y2q6sw/BMkYlUZHcMndqawBKOXJ9tien7OvXpwHcOCSu9VeMS4DtEaSfecw3
hOiQ2MrSQbXzHAlb3I7nqH77nq262TnSi6WBVdooC1FWy6ddHucHMRMPSqRs
MIHkFsAOXZm8hMFGcCn5yo6dSw063VRywv0wbikgUcQ4Zb81VtpGItJXHwAy
BQN34uMA8ZQUGCYCHiLiFOpyokij08WNY6SQ4A9TmRwEk+JTk92hUAOKtO4U
IGrPZK9sXxSgrY6iZxqcYMjg+A7lx32Boba68CzQy4Rh630lzQtpo3ioXUPI
psMoj3B+VHB7FS0i8Of2HFmHn/3IEX0J4OCFJRK13IlEX5InGYdX6dPPqw3Z
zHkcSAjzSXiqNJi+QcxfaOLo/yjtx0HB0ypCldtCslSxwzcQqlpPbEysMFcS
cPV2bvktBVgeS+8vdI6dklUCZgu1KbbV9ccOLefPqFlRev0enaPRhL5T4naa
Dqa9SGHdmap+xN7aU1KMHfl4RrAH4+9iv3ylYdlwMdwD1BdACatXK9EKlq71
y8/vGk7YVNLZNLNkxI+iJrBaDzyqbGgNXYQc13NH4ie67SnoWJmldEid0O7n
z3jmfxmCmfQth8oGSB6bHFQJeYcJj4cJ40nuLBbAuRCOcAH27koILyl44N9Q
Z8EY5zJGc5LZzzDoqr+voLbI+xYwZ53mbOHl+sqsxF+FVaBAoiXVjX4Nb1dn
T5j2zs29bfL9jjx4NcQoUAA1reqxg8DHnreFApJccGOMPAyjDFXTpo58KLD8
dBM6V3slYeFHp5omj1GqlTMBTovnzl2MPfPNuGjSoV5NgrLEVv7i3wWtVlmA
y5DWDY9sUfp1oRwN/TvBq1LmaTTpbSjGw03NRaK4mu+ab8UkcLShQQ/FXULu
jvtMmP3eiVFb6u/IPWgIA8Hp0/PoPkLSn3apzGPwManaG+6MLoAWKP6t3i/F
rYC+yTIC7Ak2409U6AlueFjkzb06fe0n0Jcyr22aHOVZWFMPJq/MV32DMfw4
dHwuG+pdkMdzcAQI86sgzBsphoBKESWUsfHkzE0lDJAAjiXOqAhK/TpyFer8
4kMZz42WLDLfm/EpuGqLmLCyi/X6agrlku/WfFqDnswg5hiSKp/v2d9fB6NJ
MyInct89ZhnZ5q/s6bNkJnbmQWdztGbIqsjaLwD7L0lPuzPs3+8Ly7rdYBxz
rNDlAfkT83b5PgsbQpUnfBsrpVZ1Bae+sOQKY+M307rup6qvf4S+SV2sKYuU
9afIMtAb2W1cTE1WB66YO/jcVHWKhZOxGF4TB+/B8IvzvA0tjL7raqCR/YNC
j16Vak07u4/g38Y9vgPPD/ICstRyok2YcH2oU4MFHK/NkQwtTgPX/3P6XzOb
DOlAoqboX6ztHMy9tQttVFesUl0jAI5dogxQO7fR+H98lY/1t6C1qbd/UsIa
v+l+HCo5n6z+ERxsYObwy97zi8UP0Sf29VPN2Q8Fx8egArFGmAoqCYKy5Ila
ri+871mg/iGLFByZm7LOkeeDBeNDtix+Wnjz6tGIephQaRvqRoSy7V+9aA6u
Fle832CG+0yXAPJaMbivIKtfynZgAcPZ7v6SK9W0RsaqNuJLBE9C+eIEwjX+
qgNsaatnTIMRJm6qIwwOD/bnid0R4anq49SIcGLGnbsklesA8X5dmh0E1NOA
PGmdBzdb8b2ZaGwhHauM5mDeB06aiKdA4lyRonJT46nppntn2Zps1hsLCnWm
OUqx0a95uN0TE+NsvglKLbRsmMrBtCKauZvtcNLsbQgjrb4DcA4v3AzGdCXi
HSKQhXlRsYvVo+0YTrf3leDU0wEtnZeQVfQ5+0OmPezD7jPGSZCoQHPq95z4
dxLfdcTR8y/0nNYsuDb5/+SUkuNT+/ssFKURLX0FxfGszfpOeKYB7MMTvq1n
0K1NxVJM7Bb8FQZQWjhSYURR5pc5O6GOEkCCnP0l5m5ZaKOnSjJIr6+Vz5Z3
YIzKloSN1TWHAGGfzW8NFLO/ysObau1kM1t1eG1YAtZNaBRB3tc9kC7o/BG2
/jnxJc+qfwYR1SapTKmlQwoFWzR5zmZShTyR3cdlwXKCsV2iWP7oDt9BFTz4
HbhY1X2jTfXXgtnqOVQYxJ6JB2O916vj7leJ8ZQtwboO14ZxlYY3rbUXN9gj
6vcHFG7/JexDtSMyUiUygN2mjp01cekANgJE72ig3jTX+aZQhSYnTlDrVQqq
S61FYgXZaDlY5XOkiduZ9AJSItDpi7ajvM+SJRhbVJPG0WKOZF3tF8ZgOeZu
TmjvYfIJyr2YOIf3nN7mUron7ISspV+qfVq2vTf7Ocp9h/uUnsg0I/a6jjwW
ZZSgy0uMFEhYZt9YwrdOf0P3X6FVbPbyRFaAnOi98wBrRmbDMzjTnU7Fg9fl
DHWMHvJG5GuPQan3JACwW4RePK7GUJbTit8RAqsQyw00Uep8aowKjAaHOpQN
fmiJH89CV5Nh5OrlA2vJrCV/ZfjSm4zynLzQCoD7x3diNh5cNEGmLVzLN6DO
Fz+G9V0aKdrOL82t2Ei7IhCuu8tCLYzF1RMND3T39E+4s8G7BRhXTo8d/MMb
tTycCO0AJ2kWTcho2dJgPCuFZcMlvAv32Zn5+Qf7aM2A+dzXMSUIAyrh6HrJ
J2t98E7jtgHbLT+JVDx47+MqMecLv9VYbR99plddYinXzyOQnFnXvprI/uAx
SNPQt/4R0q6WKRHdYU12G4AM5d1zstOJFPQemJcdB8gRn11Z+FAY6E/JTWUj
jIyVkEDgkcZ7nGWdHQWrrRiRro9+1vOvGYiMlW0VItpk2XLG5i5qQBo84ZpF
OGd2SuvMk+OdcutHrpBX2ugSycjwB7Q4QBudQkMEmuNAe/1pUWwPs9maOpHI
TuvYCzarNnV0qxTPbWyg0L2CBN/7qrwSgWlJhKKnCltGpaO7X2Oo7jhshMsM
ZMwqdKPY7bedxjxWhGGdJpr7bNhAG0vaAD9uwyyWRLpm8pIGv0KQQrUloiSf
2GaSjV/Kdhj1CX9Ii/205aGEuWJ7glCMTGEjZU6kdaHmk/gpffgh+5pIFElc
NcjbBPEfR584ylZNtU7JJP/n8acv94VDYKbjgeopXYM8T6GYaWj2Dl9K/qJq
8Tp99D7onjKUWqWdYpTBsJXEh36nAfXrQ/60D9SUVgkeeEsBtDDmwpOg+mjG
poEaJCRbR1ZYA0ftt2fQ81S17T7FBgtzAq5WxR025rbDNLEaIfhuT2IHedYb
PJwNhMQ43tvZ7u5ILtjH4NUeybPrGEBNBxc3jMlYsw/UiACq/v6X6cJLaz5P
07Zcfyj6by3WcE+I95xtPHT+OV9cqGGJJkwqNKRqg7py5MUHY7LnrSOpxJ0e
64ZlBQEtlBR4bUpDfm0IeNtSh+wKxhKk5k06AHQgTJUdk8pklIDHNjQMloOh
TSsdoO5iS1zmng9w6myePUO5ttGoVfmYdzTW8ia6A3znk6Ru2n5X2b1gHF+K
TezM8CvqEUvYwULT0OOHs2v4J3fXXXF+xFp1sQ8XRi9SSBbNBTk2ncexkEHC
iMPpI/wJZvIqw1bN7skFYMdDc54vzF7iSoI3HHDMUJ8stCD92CCJJ9aUHtpp
CkkjP12Nh0YF4MIfMjnMGW7ws2dNmaDw5ulcpghKzDL1RtTpmYVLtQlsJE0b
QU+tUG9GlVQuiMvwiGuuAmv41N/V3kW4JiuVpaT0phVkpE2sXgJpRUD9TW/Q
EWgH8AcsrrLrFPEbso4rtnnGFiK4ydoyuRq0vEbxGhglKH0Bnqw2XHDGNBZj
RyVMNhv2KUNr7YrV9pVUlbNZyT9ekpgO5jpB4pblFvn4aNOALh8mwE4yQNHo
iwVWXMBqtpAqcQa35dXzEszIXysEH01QlMF3d5QZERBDcr5Hdbi2UdoC+aWR
sCDn9Nd+ApD3S5wVXrboZK+Z2WRtoV5D3G8SaV0R0/ggUXHOdiZxfkfH5oB8
twXwfTAQRccY8bTuxKgyPkJuZmuacaIa8e5iMRf5TJ8UDv6wNcNK1anQvMzh
YDuGkM5ojYN98loDdSiUBKoFRXke3k+NpWSKWZuunxEa6qaRdmej/neW/Zw9
RWH+LLLCElwF7uy8KJj0dZS2buIy6tQPNyFAoQzY1zmya6w/SfNUhzWCipJ6
9y+qnFAPLVRq5TgUMtCEV7uh0cA9OHqvzgcz5VMdMNTvFTH5dKRGnqv0bhcZ
io5iOgzq1NAerXlqenXwMd8dAeUQrXwWAf3am1Or4WMc0KzwlnC64J47sEa3
viRuUMCchqK0COtd4IgCmidBOSfm2xi73v6qH8SbqMg1Gi6CgxZIZChoPKyM
4kqpqvdu2emHXSk/AMPuIUywau2h446Bi65WNQ1ihvclQpJW7QUn8Vbwq524
dH+F5bNdUv74mxj4i0WZYlFf+flgWyfWzPRZ71zFAVPLbhWs2zB5JgXeK4q5
Ge7s8gP/3Rr6Bx/zSLh9XjdxdhiaOxxMUYgnq/XkLXOdaWYihM7OuIhRhQdv
/6f1g3k6WKYv1nR/Jgjo4PASeJK/ZxVerYBht+coCkNSWXckmvzE+0J15Krx
ZLyW535/FJDCWVoAlOd4Q3xgfF8CCQbYol0lYUKri5o9QLfS2YswFxrAlA+S
XcYL6qkUwUYigGpnAN4LdawVGsFLf2KFSqu5IVN/L8ke1PdQXnIfoah2EGDz
3XqjLOZddeutJ7IhcRXj0TDq6XCodwgaVqc79qZEHPhf2ugh/qo4MkFi+Q+D
bxQCNZvMnntJR7YWlmDQJDq2r/ai8gc5mm5TCv/Y6LGNOa8pd9PVzNVED/IQ
rCkNC/tsxDI7jT4A/FxDCcPKv4kytRegGVA1J3skMlc+AlqHnGIB0SF1DadZ
8F2QUBo8+2Ro0eo0+9sMvcQQgRMTefDaVrX3XFpLAvewsfpcjsVdCovSCNNn
T2wycpgi+nUGIjGpWY1umFqMsTKJIQWbXIzdILUAvO/l/XbnhckCoO70gQso
/JmiRqJHqvh2tczVNYVKVPvmCU040dh3XiauhTMtiUDV+DPqtN/2duAMBgUt
1pu+tvUpEDPZyxPi2VNp9jpREokCIrbFzn2kU63k99UBbfyCidBTNAX1hqEN
1ZurJv7DMzfTBZHXcqKnP9xyYhPUH4nrdA4r9nW/tI92n8FmXqf+hUDFqTfU
b6BP1dP7VQr+ib0heNaSC1og7Deh1LNEYWYAdV8FW8m53rwDnyx3nGFavBJm
+66khJkYfUrBuT13ylpWSWYMxP9qGqjlAVQGgP/GZHDKUjhuSghySz7Dibxf
TOoKjit8/7Gv8rUeSR8hu4scRGtPLynXTG6RQoMn5IRfsCRSVJmXH2v13Ldk
dd9lJ0DEKiG0a/6EfkFy2u4ZJ4MA9S6/Z4/A+0DqJfm29l4GcpdiDvBLFYKm
3AgzbYuNoHMmBcSpm/Qwxpcxh/DmLC4W1/ZgrUyMGdOfnKJf1mKY2U1GbJiB
Q5SzKBUNwV5cgNRo1LLVjBtlHHhUzCjOtlxgX+3gBVvfAcPQlIhvzqbzuq2N
ATPXTtYQaY+AbO9acYbd79FfFAGT3uHRDIw6NFl7fX7wGrCbTlqV18KyOUd5
3Av8WDKxAIuvQG3ZPb81ln260pzWoUtFBhTXjXrIhUWsNg16XJaR3rml6OPH
uJZWISopZ9XSX3wPBXnwDdK0SmLXC4n1z8/P13nz/dgmqk6I+BJ3BYc8z5vz
Pl7ycQPT+rLtc87C0KwtQtWXwsxYSe8R6NaFFpzWlBC9IqLjVvhgsHf/IgDZ
091hBC2ObW2peFLGowo36R8a1Y9rwjUw+scFKseWxpgdXD7i/ZrsNRJkPQyH
liHBZmLMtQgLt91sOnzKIQFGJe55Uf0kCXAFSafjPFaFLBLroecvy3bVlYI4
qPN6B1r5YjW0OrI5z1MP2tc8APuuD6T/UXQVC7uJbLgxgO5Pp5RjHCt4UN3s
xzd7DaDVW6jspdCBCDUQuofldgxQTeZks7F5CLOmFPPiFi6JKb2IRTfxnWps
rxofkK8nuDPkkqEeOFbH/v93Wr+zEbYkjR6rUkFQx7bNNj5DCoDmI3EE5oUC
vAnHFUWCC3ehLU4sqUwGtoeqAIijJ9R7C3aK3EXAGdyfrxF51v5AHUMpXttK
8ByFmyRnTF6A8IcfTf+1PkKa5tJ9Cy+4i3KkyxXhWYko/F8WgpehjofSm8j0
TPFV/Ikz3Dqq40ZJnNml9UKphNNR5RhY+EN4ba7aJMGPuV7JWRvLCFqRxGLQ
4oaIjfdFF3UBEeqHOti6X+8YZN4iwnrz5Ek36Nivez6G5YtXNFeN83dvYTF3
i0hkR1JvrXm9MHMCByAoJK6bfOUD56YNcKYzPr8K0BKSssMdl3HwKCZviJM4
FnP4su8foVFSHEBpgFUAdplXaGI8Elq3UVYtWSs+E6SL+XMx0kd/5XSJHYHF
Tx/bnpVN1PpsuqisTLncS132QJdUTCK5B+1y2wWh19bhhgn1t4Y9M6uKSxN8
1aBE+b4Vxg02Cf/JjxLsV1oI8R0yxP1SVIR6BqUYKCO0l7nE7dZJvJ6oocN5
Zv/OpnAZ2gbH0rfnPYKUDO7srAx4zW7zV0KS1BoNrBeUFmMwOVlpRzGlzeTw
zXSTZok0uDFyPhXRJCQ08B+GmPtzZqTr9T8/cEKnF3H9HaP2nyxihl6je476
HYnQapP9OD8QIrePOL7fqN1Btyb+wUPUmSB1t4ZpYwcRbVj69KOaYssnWWdz
TqFBKkMN/WKCy/2MPwneFQzBsC/8kzum1O2Zb2tWnwBoWX1kbnVetuOE2zQd
vv/wyGBH34DFx8Co4B52z2p1Bz10uC46vwoj/Qxqm3/HgIvgXLQkqZJkObIV
ERul8HDqSNB0aRsgLUwHYCXCA8D+YttObtNo62LFj5n7mGwqyr1hpOV3ZmF5
owrLiD0rQC70lOXcMKS4R+WbKtdjuCThrrJYY/zsJQcpqgGgP5H7GdEK0pxp
LeznnntHJ+AFsuB9ETJ5/QTnrVLkQ7BC8FKdf9RglvnsyOWZdHrRR2EV+Cp/
7OeBdUQutCNin6uV9I6oIePW2eNjWGrO+09aqyLH5x51DjwmlgSbnYSqrkbl
cSQ5J5Avd3aWVuB9cmxcOJ12LGFHfFiWBaSCUZBItwjQGTcQgGwn/aoxAYXd
N6CEOZsf7W/0xisUtC10SgwmvEtwVFLidT10Y3Fy2JhIzIMXv13Kh1p6zEnm
Isfkvb1yQA0JQJ6UFPABz0xl1wxd8rBq9aeDmaUdYr7OUVkkOLmxwAsL70V5
p648k41A6dkl92CQNQq7iJPsB6hsgzi27AQIPQ9VItzUy4DE+Hq/3h2PXoOo
7aKRI4GeCceERL93vB0M218iLAd/JlgfSBfRnR+nLkk0Jc7LtRwvyRiKPQPv
cMi0BMsHC7ptz9BvCJC93fjU/HqnApjve6fHPfg4HbNyLJGiX5oLo3XSDZqF
BIhVCBI7H7PA+1F2oQ2pWDcYdLMgHtwiefGNB3y3qvvcaoIARNK4M/6g02LF
HdB9OWjJpKYyh2iEKnjxOH6pHvVk5JtrpLGUAoOTF43fi4XUzvqJHgVOx2J2
4rt8Fl5xc/bpzd0iRwrI20aBXloxjTNNruPFhRTzPDd6LZb2BbuFhRY+z+qV
LCleqSgtCM5lOWm5PWFW46A3LH3NzdSGDIB2jBeNTUMb+hg3aW+yibU4XTFm
QOukyZ/XVgBHSV0h09qObyV5HSDXnwh8BCI42KSB0gvhkHwBDVuUy3F8Bd5O
WP4vZVEvTMY+R3OCF9zR/mTnzVJNImqVRduX4FsftUqWI6nN9zX2T9/3cQJp
IOV/JuG7t2WRpQCGRr4Rc/qiXLqbxcg0khbhYiOnMZpFvTrrt5GgG5dSHNR/
y/+afVeTGk7ggB5KSv5mw05nmXMKY1j5kRf10Pu3a/TP+OK/h14Vw+HTShQ3
4dlsjFY5gdwH9FuaqPVfAn/7JMPlbVLn8Z5rNjTAFkARO5jYikhsLCl8/phN
2wjbWm8ZqqWnFZ1XtfM7R+nxPHQLh/n9/l3cUFs8M5inHJi/t1vz0ZwVXw53
nn8N4Qd3sKV9LrdDGZEEMDzFsX3S4N672Pg6mMbwck8YoWemEGmfT3rFhmj/
TJaPMV2njgdUjmMwoW2cZgFQq35uSR8GrDiCAKtGsBtJCeT63hPgeihF+mJs
8megT0ayynygz5s2hKE9QOyu5EjPJkflG1dpAqKKEnL2oA1oLucWC0xkWFb3
h/RfuU0GTORPjS6iUcwjVxLW/YHD7U0uh5h1QE6iPT2evEt0rCHZgdMXlwCU
bIqZ+vn7rq2dKpf6kClEo88AJxy6ASTQYa3ntXjuzoIub8ZfaUDhlD/LMhp8
088wE/tn6PO78zm1xHHan+t3bkAezbZJUtghRCLmgfYPusFiOyQg5QM7KpQh
QCkm1fm/VVTZWywNSTPmm7WNFcrcM24n7lG1q3S9R/eUGZVtyKcxTtrKKVJw
cQWXuJKJqA1OOEmpG0vd1xmfRnR/KQOIFNBDro61oF2ZguNGn8WFQEZYuqRM
3RHlgenMDfuh278PMgkQEnWf6l4IXij+XF2ac+zUrQ9FGIsdqYPHxX3Im4Ny
nXMk67BBJWjVXG1CDKpeLDN98ijgIo8lEsk2lEjxJQx4W8M9lAUOksn9Y0pF
6E+o0GGU/NBhCcKWgjfDNgUufBQTMqX1sishvu+h8M4WEsDjIjTTa4DSPKpV
1T24WeUSuu6yK1g4gjNNAtuWi1/PFhlVCG4d9m6cNDF/rIm9tr9cmeYC3cti
vxBzDqjL+jDDBGO9GdmngPKaQGPgtVrb0UNn9Jyz7QyX3rMbnY6q9X3PfyB0
LLcpU20N0Dfv7/IjuUWQSAdB0h0OfJ0US3i9RQ+L0o/ZnoPbjkRhn3Qhzhwx
VsiPPw2hQsBUr4u3FopscH6l4+tlTSiuRVlTjRRXE7XPDUapaCGAic2IcwLh
e5Ker0H0PgjjuRVkgsoNziEMO6MHd2SQBvbAd30mXLS+oByzg/7I4vsSRY2m
qGLQoluLQtrybGtGaMRTyr/A3ZV0GXVA+Td7KtzDVWRlwYaNWcbeOay5mAgT
lQZiqdI1ZaqNMJlRASOKarvon+Laqq4OblAkr8rMbcAKNM/ehb6IT+ss7S3A
iHZ6upUeofGfHcQUbhhORGqMnhOwD5iVrxb/6z0/+75VydBxn/Vx5O7HoqvV
o3F2Ko0BF3xBpM49/Mxoej0yldXDde8pUNV35Rtd1m00R3GJ3UgV5OeUKlMY
5mdC/UyvG/7Xu3KIq1o22vp6G196yAlP7NO2X0XLBbrTyaoHsbN0lTEjqaC3
lgiaBA93FlLrX+AAYyrYKD6GuiAjcws42d7mZtMfz4q8SawxptbKGG70Qn5+
2Vx9NOjyStOISYNIXRoa/+LzI+3vLAj1p+nBkE//+7KAFn2YlvnVJdXAqiBp
A/9BqvCnNHAJ45/Pcb8v1Y6VPSmzqrg3Cvlhkk38fSJDHtrJ1a/xBlj16PYf
v9L8X91e1DcWs9l6NwduB5CJ4pRt7ow/C6v3Av8l/Ah36sCJkExoFvxGLqES
PwBXHNl+SHB7rF4KhFkBc0ZxtkEaXfokLYNrU4n/99LLJXq/s4iMrTu3at76
voYvCiwP2q3UxutGlvuy5rga6SHfgY56IJnx3RBfXqHXqnIi8bOCR0Ev8sll
kbIQoUOmNqcC4Bi/CmMCF3Jlkj2sRctQ+Hji5x/hldLF7RyiKdi/+sdVRiIS
oHtsTimqt7kgD71Ur0/Xq9y+tl4UoND9RyOhKPFJwF9s2EILftzw35EQp4pn
mgFJi1p7O26Zp8o5uASBhsReCMyDQoF6FmQYfeq+gih8Joki+DmdDOWn1Imx
VdFJXGXpeqihyL/0y3vGrKd1uGmXqSpWp2IhB75cba4pP/pVec7VfGtLq6vy
31HORZL/Xpo9Y0bDgv/nDfvhEB6hskzEhWwmoQIhYmLI9Qr/EprRK6RY4slk
AC6fA8thCMIEtMF656W88BA3FQ+T6DMiP4VeA7OsN0IzSDCh3w9LBmsCHqhM
aINOKrtZFx7yadiB277oa3/KaCaSlwg+sMciEe633QoeA2DmR5ReIZ09RXGP
hsFIEOBnU+X8MFeYwxuZA1yTPyr0ikVE6hxlxs4i09EGGlkb0aPrsU2y7IdX
5/w161/Ynr5URfVlgbFAw03xL/aO41fSL25tNoPGEWnyQbP7gGe6ANXze6OU
LyNpfGCVSNUfAwdLyqIwk7r7N6BoOPqLMSBHwvI+6GgPrESEw98yGkcP6ViE
pkjMGHO6YNRhmQanNccpCOy5VRS9dt1VSqYKP0cLczQ8yC/6P3vgrbe0MI+f
RmLpA+8SWrysJQe0QJDKA5QRn5lQPVU4pmxzeAztaG9SIOPJJbD9/wZyAhTW
3LURVneKLfnyjdjnnGhZics0eeHUOhH4IxCdszgQU+WqFwVkqO1cSCWeGsIg
rIK2tRnaSsGt1FAdXNlAA5mS/0uPotNqTDscB/h1gIPad9gEq1K7zdHzVhZF
trk6LbzDmD+mSiQtj7BYvCTPqDoApvNUu2jS4FkXoS7Xpmwrgq7pGOR17JDN
VvoNCvtAffIVRODq+45s11wmpP84w8kmfXvp8L49K90CNAfyV9HnBhVuVxIb
vpbezuV5TqMC/3hs0jJcvGpIF5KsRI+GYcVZdaOKjxZUhX3GYKSJrA4pkQTM
yKpbO3mMVZgWvRqExksm2jk2CJx6jSZjnnGGEunqHWUpBldWnKxhYvsFE2Dr
PIwPdqs9EvQZb6nqz7H4P8I7Xzytvc9iHY+kc3adVcuSdMUFc6rr491hlgIp
OU7q3IU9cSvEqpytqQtqsOCHzd356oNdbcGxVTdtrc2nndk6Hyo50KAPe01T
efY/Q0WKAmYwhGo+VLJTCW8dOjJJKmiC9YmEdOrXyPBWbfswb4yd8UXWxhSm
W9Mznr67D4kwpkbzy7JjQtzID0fKUojti8+GftWmxwbRfDgzgEUzTQnTE48T
XJlYfX2Nm7kOUyaTG1Wu33BTuS1ycGGdtq8m/rIb7bcE1expxJRRDuTqzzOJ
qrv9TRZvMeoSVi0dXNyHN9j50o6/Axrg6zqEsZdlilfWrByLjvmod8MH/kIa
J2FB6eF+eDZhk9Ije3HvoaOBMka8ABDini9wPxxMEyMSBzYPgZ5dbIXjw/ez
9L6Ue2BSx80zznA2xce9j3ttARyM3Q4zZQGYuQXq8uUpyIw3glfAutkOpnBv
WhYswowKjthLCvmcV49HLZla6SvztazzcFPxihSqNsFcy7EFx5Ir47RZwUlA
qTv5/YEh6wc2RSmIthwa4x2fwVNjdccrL4qZT57RwU+KtLAum8QPNec5snsJ
eyUbxNbUr1cazYAZJaf/5gVRxPFNQIemuz5x+ow6cSpxMUcJvmxGAVeLRtTg
/5uQYKt6e3iELCQk+7TaNyXpg7fhn6tX7z7/UxFm6kAzwi8acdVeftrKUsoP
a3CASj8HBIF1iusnP8Y9znfvf1usQXVyhkJWcu8EPkxZDBNNyKtdBZjCfIBV
5UFaa8NCjhq/pwQFDuVPRLQ+Vf2n6Gxm5qN2buQQQ7XKx3armqlE+WK1UcFB
kiEEnz6OcbzzfX2Cp6G55/LomKOul55HCY+k54gtpKbe1eNlss54iBDQr/Vb
TJ2D5dvw1J/RxT0flTR12h3ZYyDuWK5cpd2LvSyXDkr0oaOlExZqFbkRuQ+/
sYFvEM/dUq3SUAGR2lhtIEdfmrAvs11DeaniJ9MUs7oH/4yizUUh1CcywBqz
6TFga4HnHi5694jekndsrN9XSlSJDLhNnUnN9coakpeJGdGL+MJocXPJhv8U
5sM0gPCd73DKIjKQMAbaRJRxMPcFnlfEViYkpSC1oNmkVVSRUQNgU3iSakzk
4LjDTeJnzd8dt2mINQxbyXctIlzIlmBejRqHhw4R2amDyU06UfFmM5uUonoD
vbXUzzX8eKWBTdg54yeXdLPfScH4M+G8enzyhAYroW+uD6FiufQxYyHenFg0
pUbxV4/MsVBf3Z03RlMtI6einsTkHlGdsT3RYDnR9kdx7GAO0xaJJ530K8h5
W9/PSWehS/DYHLvvyH1figT4UaGOPmwHE2J/p7dlsS95oAxMnACNmJVIYMkZ
7dy25qLVuTKzWk5z4qCiZgq8hmJgToyZPtbLPI2iHKAvKcdkds9DUoyRR0ug
A6VtSMRIhk4QJYNuKSBKT934UsdxHtUNEOeJmeK0B/GnSAdo7nePC1Vtjd2l
tuZ9DN43IK2eYc3m09ViWEF7fy4wPo4ptPyduUQFKCvxJlfZ1FO89txtXAaK
sIdbOvGnKIyx90vDNW+Nrw3sXDiDSBZSZCm4tXkVnzxoMBju3uGypdsNSW7a
tKnvucsoE50Kr/09RTRYoeJ1z2KMbSmh3Je++HJjicW2oHB2POMY82MDYN9O
IUGvr2z19nyxn1Ve8hWqv3HVAVnI2uLDdzetvIAl4nBwqzJnt82yDGOSML3d
EGfv510EWvntdml2v7xoxhYNG9b/Mts3nap3xWQgQxTDmnMppDdDLoC9Ihuq
rTOw+pbEWr6y7g3ZqIv9QiE0S1G0UVJPnXyHF5Kv/e8uEbkL8AxMGAIN2+bt
v7ieNI8iut2J9PD3yeYllh8CjlbI6FPuwxAzXXKe/QugUojgapdnCEyzio6u
k5YJCvlPrj5zCLoRUOWV2NHbGyYEUQ3ObBUeQVdB3zgCdl8K4DZPxvUVrpis
uYhIQRy5VwF9qj78oEEOTvl/FyPMm/2X138U4NHk8i5Pu5ShdUXqWej8kNtm
RRvf7gocLygHQ6RQg73zDube7yuwnUCu2S3tJ7oeeONnExeUrdKJWgrLAmKs
/h/gnokoAQwXvahNscQkmIJvRDVtIA56Y8S1Ng1GFi3vW/n8ql9ta3ib2Z+x
MKeC3P8eNQ2LhIyeM54QAXcNxf2OVUuK9qxzQy734qyeciERWeFI1Z5yvnNE
bUBShIfZRD84jpD/BC8jJVZk3GM0nq35eJdFDPE+WxhSxgMD4NdCaijGAGX0
8Dzn8Wn8WlfFiT2UneUFEjazay1Iv6G5wZYr8XJvUEmOGw+unYzJRS1Fxa6R
MUB8K3gwkrBhInzbyptdL9F2z2hDHTrYjjqOhYJVeLn6VnNDDjOL1/MEI4uU
tqhRlxUknDKYGkxLhkR50E7P/Fhkc0B+nsPZ8bv4W/IO5wTfLdPFOf8t1lXt
1dTFtYlwW4Sz8JJKj+govRPalRz9iao7lDHQoDnHub0GEhw52uC4RJ2ajkVo
2LjBxXQUt+aJIuL7GUuRE7Cm73RfhTY+sYXXj83fC2GzPX9njIcMi6Yp4n9y
nT896SOzBVqkT4SvebxoVReMlBQ8dHAWa81RebdQRRsMkhWVu/Caa//T1+gS
o733L7t6d6kPdXDs9moXeEG4kRI795ez/9RqjFKpUU45VMpQy2/z0GHaFZy3
0EkOIGUKpctC6zCxCdugicXWT5BAhGi8hRepydjha7jIAICFLM8TLTbbzilk
Utaihq5DoD8Wpgbc6M2md0kkvDZhJHNa1/JwmF3WW+8sw5AEzHCNLMbPtlXy
KgZxUH2gnplKUedLNzIV5TE072egJJv3lPWG4No9Oa9tEhlw9k4U5U6tZ61l
8kq9ORPYlOSHtoqouuq0RMdU+68foUP+7xWnleZOr1I+J3Kti7AUhjJ+sn6u
QJoJC8A0ZA2wgswyzsxjj4ojG1L0w7X961EBs8Knhq1ApeYMydijXkr9GLyC
umtOWVVsUgvOh7XJPTvTzgbCoGUzIRMm0HR+sRfi6CGLlkBJruANx5r8hWsq
Sg3NOTSuPV/LlApzMWWI6BNRdgDaLpd09dOt4HeYS8lcK+SyRL8cuhiDsjgT
UrA/JvJMAAAYLvYH+OaG1q6n/BRr4PY/JISUKBkSwvorakgxLkF16epmt/aI
lI4DRZ5PxoEZfvFK9tNxl2jp12VF6YVcXOYr0XLIiMo5cwIPbYE4WvJ36t4l
JDEVcZYEZglWx37gzxWzgUll0U8K8bnZYkcJhVSLLBlAUYnXQGmfwujIgNPY
pFFzRl54hI5nznAwymVAXoLacTi8rJHY7dXpxcasfIoN50BKh42FQVueVpHt
wabWYpRy83xpcVSjgblarpImBd6GhnnVGAlMAhWvADiU1F5kF+1G+8ic3AY6
Pc8yvh+kJWAvtnNfOUBPK7nNv+kGM7YoFX6Le/lC+kXSQGv6l+tcF9S9O9wN
wgqzwM1WNPL5UlyXifFFAeLzVf7iQstchrvsemjjR4E1gBes1XUilJGzHlqA
bmzhVVdo2jrXBN3TFBIaM1zBj762CAah8uTUECC4zsRICUO5JAS+0UZyYdhH
XDjQbu1T5s0G36gOFlsAi8Bs//aO3zp9iyoCTH+DZmC76GuriQ88tONpGedH
tZwxLxmC2WhDneKNj6vWN6B57C3h1COcP0x1mLY+2A7zQfKNU+ZM4LR8wB3o
aqcNGB9/WoUvflWGayVSKk6hcUc/6/ZAU/B0WZdflhKMdbhibvymyBiI4/Qh
KVaVhmbYaJLE8ank1UPptW5D/v13UTQnWtI7kNyowqfdSEu0AB8LtUSJlGX3
vojC4Rk2UGUAOvIj5wqFHEaL5OT+fQX+D1/MLgvDWVP3tAPRBQawRe59bhIf
KIRV2xK8BzYF2es0N3Pc72wnNfzkKaFSMy3z/XUgYIxoNS2A0JMrxQAVdAqp
Hhw+C3K1E5lwkkQwXc28QrcRJDdPl/2n1j9ZqZIrmQLkybTZ4IqfNw+7dGdW
IaDBQK3TmdOvNJ4u/9wh0z/zW7f3DWCiQURz2Tyk7KzUsC1c8j20szXJkDAC
wCChVw6Uw5Bei4EURqVK3WBxGMswUhleN//pIgY+0YPQTNqzHBU8qjI5lcAD
7rETZn8L0zqMzzzYGyspmfNcWgeWbOnRVa4nP88iHMZG4MprlL0J5A9MccKZ
+3O9NJA5m0kvU+jRPom6QCEFI/lsg9Zc868P+UKa6F0eETw2JQBzXCUzSiKP
Uqd9cjbGt2Iiqmu/6B2v0oQRg60h6bMTrZOCjtxeGbPFnWzG2oGoJhgosU9t
ZxNYv7KL3HVe36LmSlBxj2Rjfj8kkbLKFS1Fu6vfRtZ4kCbvY8z5CS7p8flx
MGfEEL+DR3rAlmApOOSmZnPd7b7VRuJUX8bY/tI5tk19GUidqfQWGTidsyCH
l6XnBorEKRj/kQU1bIowgcqvgkzLYywqgSniLOuCbEimkc9wTotx7peaVzyJ
KWlB2UqHEToqt8KBLgHQ6ttkb662pXcKu5EqJJqXDP/Tat80A3kkXEIvlUY6
0Cuv52wCJs/6IegDmn2RRCqqSZhG3NGIaaDm/reTIO+IwmX9MOpcENFNzWwm
prRVMLRNuar5b1esaqMkYJ+tmX9JlmbXmA4JxbkIz99ydcapW6T87uM54BAB
PxhJ8pP46Mvj6sHhwE4hr/rdVSVrpP3PD6BDLnSeyIIfYVp+1gkix8/tlseu
/SnzLv0JKy3rzLQTliZrDIDvwJ+kBy8PvoA70ygwAFsUqTgtQEAlxDKt+87/
cZtd6bz3lIfiNoZ9rulZGvjqSIBwlCZBYrS7m7+fEH7eBEdXFp89wc5YtECy
ZjCE7aiSj/DHWAUpI+YA5JFMuKMlTraKzLCGlUevf8R4SsuCyOosJ5GJCb7T
YiP7H3f5y/Si4bBJB/qspK5ibu4jsorjFpUsY0EIY2AaaVkRBmZfxEJksDiw
DAsiNjarPXui97d8WZtpR9t2Evhyxu7NJzQvob7W0o78UTQBpnGhpR0MBI/d
IwjjVKWykDjkWjo9RqkJXhVp1YE03zJgSLPOY2wxipPkNV7YdlazAw//3en8
j4/DKe4L5/06jd2EsjnNWqCrfMRH3Fp2+X8lF2OJ/S4KBj2kOZ6EuMfwSlYb
Eke+ij2g4uMe78eJvEjHUDeOe+72KQm0RCgjXBAfWbnEV97LO78jhTi/1QWz
CRvBoxmQuoO8dcwWdN7e00B57p3NBnXu80JIpukNj8Lv0+xAHJ2O8KxzjJ1r
Y7UVVPgzM1d87KyGWHGvVmSAfaaog6xI5/cTXbKRbQKTJ/+qDglbj+5ihZos
y3MDUP1pNQnCApMuMaSSYcTplw6uA1EiwSVy6snqUU4iTorURVdrPyQ1HjuA
VkB+S4KneqPhR1KhGgMIZvcp8+lNwizD+ElvzNV8SmTBZtIPFr37K8JotAv4
NqX2xM830DJZDbbWCDh9BQ008cpugSIl9cTIbXqIiSQq4U3ZwcLAGIiDz38S
lW4qiYcI7YDEpuM2A+9/BTNhrDT/xzJPg+8sTBAJt8uE04GWuPo8J3y+YfFF
g5A7pTfmf/1Cka1Jf+RJ3vlZwAw6qqTl2q7LopCCz10n/72TsONZ6m/kRdzS
W3OJAV+his23lSYEi0se5eXVOIu8xZzGym2d0ltCiISPLA5jx61CkjZETs0e
CkgIIAoYsQ3uAe2nWBqjdpPJbvrMgGUefqfgXlJlnPziIyJakdShbiExPrgI
6oH5jc2WAyjofb9kkw+BgGtw3hSD87pDql5QxBXNuiUK3syZw8V0L780GRjS
V9Jw7dPETC+ZC9jo05DILT2DPiC8Itj4VldQkJwO60nVojPX1gurBLki5x/4
vE3qJVifx9F4xCz9+EjYNjgjU6YpfhknTFic0CAIrxiSWfgP5pXtE9c+o5Qv
4A9vzzh6m2vc5bGmMOtgdYdxUqHKnIiTkBQQnV4PXAGq5NmRL9zyefzt6XT/
2oa7gszHmoF5Z2nck/hV0XR7fUijjLhuymDH38FOdHQblrAuJaacceMKPYGd
/Z7aPTUssa+ei75JSxsiibp/GfJV5zLtuCVhS5WyvCC3NGB04WlO2Sob04LQ
KsNz1C/WLNhXenBCqI7fIZohPcbitQH7KF5yoATSX2BBq86o3RREa2HWfUde
LObdoZdVq6POcCeV33qk+Fm4lQ0rDXhnEn226eRbXRSOXyiJvbnbdbVOB2CC
N9iOiDMtgSk1pz04PI0cIN4fS8Y81Va54wAsfSj//qRtfF1XJ6LeTX8mRYnU
2UnBsPFwyOV8k8jYCBaU8spnmPUHIfyvkfPUGESlmOntjneLmjqvvAOe98Tx
6MFYmIG20qRB3zj30OMLab9PT+ZbiWMaLDNRnBed+vbZDshrdBfPkOqXvF3+
OYPCxeHEKBL/+YWFoUmtfM1qpQO1Y7xbettnqAQkJsX8sSb4d+SI5xI1PnBT
z7WZxfzn0BoHBH6+bLbjT17P0DY4RBABEIzKvLs8huNgzmPkDyiHAfpvpB0Y
Ju8qlGSS57nDPJzpg1YvW5fORrwL/IST1RrdUJn76yvRDlUxDwZX9I8hj5CV
lAQZr5oTyOpdXmvCJ8+SnxeFI3xUfVg2tqXpKuS3WVQedy3mztBqmp3DSaoV
GGXwq4aACgMcmLNIP2+nk9PmN0XIWi8Um2bwuUBmBPvhwBDMA3/K4+cFZl25
6Y0BtVjPXZ4uRynC9bde0DMHccELhcSWPAs5HcqOc0yyG65UIGPQWdzY4Qz6
Qxgc5FfeVmpZQoxiW07N+qb0iBcEKw7huGI/4h6R0sTMcw0sr9fm3Gr6tfuR
MgLCrfWAI0DjRXgUqhuNHnu3dGfyZ5RIAzCn90zVdwPm0xX2XOm4Jmor10K+
dSG+MSfNdFzK0KCV8ITYI7+syDtIDNpv7ufHLUcil99b0esXqsFSSfZZzOhM
/ZYNNlS7FoKIyZlC1UM+GYoHdJNfgzEO5GSDnn+AC4c9fSY6FezyZrTYOpWn
cNQm0cobUZyOvjwGQ/9qv0VY7skmcqeTaSOtzn6A9XlSXeQyUSmVUOdBieLJ
+iNGjOXQNzWjBSaUzwPTRn03dWTGoMdZ4M7T9XWmrDLlu8C3iyDOHmxaLHhz
s4bchZDsqGq3UPRf5ZS50nl590+WCClmM9KiwpcZsjNedSB1r4AJC5a5JvQ0
+XO4mKR8d3hw+S/0CrK8IcU2zUgVVfn2zU92/Gyu1kRTXbSH2+SVCw5vfmN1
NfmtkpMvbZq2yUcw2OI6hod8teaMAKULCJ7ryQPBxNskEpRQ2dESbG3aQPDB
bBWOX0LwvY0DeGfLAKtRYud9dJRTqait5Ba8HwXYzXJjB/ZtINiYLgCLGLv5
dKqiFRObWYk7QW4DLRAXYbNdsAiy0EapW9lElM98K+g749McZMKSRkOmmoRc
zOdVzn1Qaj7Y6c9wmTf0JaaSFE/QBXU5m4ifInx7ecl8KwWFnD7i9l4SphS0
WyG7Wl5C9iC74Iz4T6Ae+KrEtkVmcoUPFOMQHNSOBS8kveTPp3oYMdCD0KCk
YZbbYsZNHgOVybw8qx7sWYoAF/Blw2JGGbfqZPtBO9/lQmRFdNxple9DdnUC
pkaoRVHmOjkZK9tEwqlAeocaRjK0NbB1UEi3vbSIhkmwH3eE5ZVOg+x6orf3
CrB2ggEJHDTw9to9n0G93MiJUEu1ByX6zvO8tUCNE6n466XyqwE9JMEdrNUY
Te9PxcMQc6R9vdyfmGXZBGU3bBUE/K2VSYeuaVEXHdzwEwXEP3sY3Vi384bG
kQxyJkkhp4fQcLAssyXKu3FwifGpyiYE8D7qVxpPGIjsG3AsJLLTSC+KYPx3
RxawhsabijZPcx3hIWbx9ZdYd/kgoGiE7w+OJjDQwVtw5cp2Xg47+m6dN21K
RyqF80p0c8hn8JOXEnJ30io8sMQwA8GKDpQsyLwGYyButYuAYON2O+PABdP8
uF2JF+i8etPqwZK25nM5Tif1jj/w81tqNVVKgDNWq6BvAtBVVcH0y/fpJHjD
H683HMxqH28WMpreCCNp/6y5PemUF6DRZ226QSqFWRufCRPkQ0mZRw0bXQ8O
Fhurtko0w49m7x9X+4JkwSrj+Bp+tPsQjkY/bvp4V0/Xs7476rFVD+Q5RKlh
ttkG8Uttty7sC2OZSB0L8qYZr74j8KRi8VrnxMQYXHTkc/UvlUnf1Z4SZ+nF
bhNBqRoyS9oSsZxqjGERxydw6B4IIHxGK5jDASrU/FrZ3dA0QH5UOfOBGmqp
dSTqhDJ+sMMC87rO+kKioTMmD8ABisZIhqPIgGrbtXrB5tYcAlPYCZ4H5exR
p0xUTdqSOVOniJVmoQE+R97eeFTzENXPvLVh42CExSy5MilzjcwBdedu89r1
cARvoZfQErorQPBrf1WH6rHPwYasBxDo1HFi0SQ7LzlspQ4xyUH4DL+NPbuo
GbSMdHaGcgv7g3P5d5NInb5lXRKGS78kCc9+goURhWODo483icEtG/aXYF2v
LXdb/Oa9zzIrRL8Cp08doJ6jH7TOzjUYlNU8VWsVbXPiqKUtleynMEL+RwPi
6C2ho/j2sYUx06MmggRkle543AJfriVtKbv7nyvPVvWCeMNC01taFzsc4IuB
KqqHpKx2kpDacOdnEFXm8aYB0DoJEirIBxBl54oNs0NZTMmjFfyTtZWxxtxA
oG6UShXR/NW7jT/QTUxwdL7OMGJlp5aqWDq4orfSp5deLsxOxdqPr99bHhUa
XbDwBc54WiUW52xzvE8VExIE9MVLIFa8NS523YD34BjdU4A6y9c5TOhwVUlH
sHTKFpwjyevlqwM5SB3ioETlgS0XTaBWZVEtcGNK5u+YNAW1zdmjFtRqog2n
tC4O7yMi7NUyVMU9gOu9D18GRCLDPvtR136LP4GSL3boDYk/58xI9/I9/HbT
gtvBH+2jVh1u1fEeyE+SYVSbUdi0WPgEXd1hMUlqd0WWnRSjJmDLVEs0+p3j
qthK52mhCoI+QDyQ5Zle+wO/gW0YOuIN3GMk4zeKaH6a6sGrp1agNzeZYGtU
2e7xhFfCNv4Q8VVGJRY1OkfJU3mx+8ZYIylilh7PdgbRk0eDuc0X1B01yrI4
2erTTWcdNlY4uZJN5MMzHjRlRIo0T60X6auWrLHG9n7RD3tRmYAm4jwFg7S4
OldLdbZ2Y/mqcatDEyQKaUV9yzki8M8aNqfwqRAYi4th1aaJQmaEpRSfBk5i
aTT/O6EfRRoCIo+76dtzih3y3AX87S2GC1e9vw6UnnL1UWMME4kKcmswdWdf
gIUKD45YwJpGtM0TqWCqkji9x5yvBjaNPkOvOC73/H5QwjTUbjhJmzk4T1o8
yw/6sTT5nIYciIsjtNGHbGX2v6UBr9YS77dmE7eNAI46jui3/GNolkeYLTYz
yhG7dPtkcssfSV5P4baFZqJn5bmli39zJ3OwL9Ec5DAqA9fe4lr5eS7lJCD0
EJeKgI2d7G0jzgKkiBVHhvZyRVnSHzMsPXuUMMF4cohhqKrEsfownkh14Zae
x+U6phDa98+Fj6iWLDD+ZmAzQrNna05+cOjYRfjgDS5OhkxRWzV1zlvF7bDd
JNxO/Q2iwYw9YWJpHgRxRLrSX9KAkcZcQCW8JECNYpf1xGn39b5VFoGbtPf5
FheFAwPwB7J7ibcopVvQvztaozc+9MEliwild/3nIPnnHFqT1ZyJzWgyGoDY
OIpCecTlonydd5C5MJPJoL28TL3LJ1ipcySlA/bNFiDGvj/MR9+OhINlJW6c
+Ps/QKOeOGwB/di6CxMURflMC5aFZRFdoposSvI/n2X7a5rla7bkOYPo11Xj
yniaexiNSjDBdYjaOOX51jrWudURaDH2qfKb94+Sy9YdoL4DgvVaaFbFleGW
PVhaTZ2vdL+N1qMAp0KFWy/zdy7Cp2wClIm+BjZS2NK7uh8U09cQWkxWAN4I
bomcNkKlWLtbsdKm4h6Q93TWRQy6cQX+f9t6JmQTYsD1uZv5IVHKb0SBHWTm
nTiNtVJuaj2+LmfMPyRpX5D609O0RbSS1h1WyKLOIichScNTzUu7ctgzRSBC
hA+AOrTI+7w3vQICXfC6s+WpaHlgihGZDKRSyx+z/f3/Lo35tQria9EGztvW
PuKUsRfsCw0lxQp5ulKunD6Ia0+FhHR1v8H/6ForS/sATr/v0Pwpt4boBUgi
5pVOA/DF32i2oITleXrOuXXM7PoLQAytLXHQEpDSGx6nqq2ZcPBCagRcFxyn
OAAtZkl25Ky4s928GRhePDftyRS8+4dFrxXJ7PcpyqQ3El+N09EgXCc5RGRH
Sxe2mgb7C3JgKoVT3eB88IRZv+m6q6vf1N1eEVqxt9zRPZBDwTCjZuYXS0sG
OaJOrxHzh62zFt1obzxwNpn/lvGahDKaRGA6IwBOu0vPrW1x8NcN5OLZwW4T
wR71FMlvAHgyyzwUn9JXq6sipYYLEPXHUTd7UJ0y20R03pJ8Jxaln/8wp1z2
gyDkFuU1kXrbrd0wBW2hnstrCnaeuiEbGNU0Zh/1mnHfTSULVl0SKcDbp8Dz
hMxK7CmdVDKHbGnJ9Ab97caXOwSEyuewbRTA117dh8UboabwLHldVuZf7xW/
630cp6EHF1exzCwDn4Zq1swJQnqvRoQGKElemPHEssBYa/iutl2gm3PyahcI
wSsEUCn+zuoZXAaLAajrIsvseqbLUfF5dBKUUM0xp6rOVrBITVXlS8PcCQBz
uzJIFgstsjmfu+C4sMsbwxfq3mdJTE10T0XrghwcT5EQjXpca12DOas1EUOs
JvPi8elnYWtQE4wV7uNHLhSm8UD/GqmvBwfPdYkRS/5DY6z9/vGvT6BtnS4l
iOZO9aTGvGPnjRJp7xiu8TTtsMoMAhtiuAi8/hGEQOOnB8PGQmI+iv9CyBhW
OcyLWw2rq5tHiKOsNKvMgA3Vj/EID+9FK2PxZ9qI0MeUcVjtNDsPFIKivli/
fuyvpJz31YDa+CU9fmyRjYqIB5DOfamSZmZ5SBm3xolgioAmq0vDVjtIHcc7
n5b/8aLkTbr43ug9lvrPW0z/xp7Ddgsq4s7oa3eV4FtLMqPRNPEEC3vt0bO1
T/EwHRTU96PBvFyyy9HWR2EVuBb1Jj4cRC1I5oV8aSsx+snhOs6SUqXVQTC7
AhCrwL7IUn4e4/7IZqO9AcDXRi4G1FP+LbkCX+pQLuyADKwcnQ+TicYm/nSA
nADQIxkw+WasWV7c6kyBf5LhNVD7WlnkO81KGkum5I2WcG25rMMCgl6/OUF3
Cs63HM8Hawta3p6haecPzMCI37uJtq/zR8niGqFx86WjBf6r1ah/lwiGmBlB
L3TF7zCGMJvyc/ZZXIMZJ/UdlDA6VdWkXPvwXdZm07Akpk80HxVsBrs5elFQ
1Pg2DQkxGZNUVPV0wtZxVhVW+rQfklD1/xnm5BV9tdAjsvEUoITgfq4DjlXP
HiF9OoxjIkxZeA9R3xl5OUDpfqcDT1+586cl6ZV17nVJPA1lhlVVXyt6PfmL
HBwM/YMP1EtmslDE+1jLa9hyHdm8nnui9BuLqix1vvTRbua0ONZA4j71fvTb
8oplPlX3OpmQpDvADvvaS/chjhoAU3FciEzi12A1ni7frzZeDcjOiEu1Igpd
Ny4H2sYd96AMsKedOZmdol7ANFGnVsHIVQD8IZ2kQu1wsD1Nr3/1P2oIM7+o
69hheWY3fXWHiqKXQdH21kBz5nU1hSRMpC6DieGPtIe474CpbSs3KETUWk68
GXF9ZvaQq2XDIA4hOmvmgNQQn9HMU4JxyjJ//ze+ejT4cEKeLGoXCUxbQEA/
bliVPamH2qOhBPK4bjV1tBrNfxDb1Y4B1ovT6Zx+obhv8EAfApmRQA5MZlPk
LdG3j3FnhbG7dfGIxhgiuLsy05bkeZbvPx/RwPYu/zL6O+SnEqQmu+yg6edg
7arl9qoH4Lohgt+J0O4JH+GK7tjM2DF2Br3iECkT3KCRX2trKnIiBGT+9Lr8
zpeoRBASS/hthazVZiHZ0X9jEhhgQh7r3MLAKA3fzvbkFTY9GxDecwLAhWF/
/y9eWtXRbx9vWoP2S+3m8BjgyQIDLMBiB3w+bwxuJGUBeswxKbhwMImXAeRC
+L6KhBur7k3Wn4ZiApAA/YySDUKLNkAuNn9JtNTRLrXgSn8OGAiKHVnnq3GS
r/125hs2ft3AnJnUeyCH3V8j1byGr5jANDyZRf0VgssQPlaa6pgNV2d+HwWG
dEzu0uAKnydnzfsMvnqVkWi6NcH6IX5lfKU1dbDPELtXw7x32wDLViTW45fV
U4SDUYsj7mDmqEaDkdIygVcpfdon3poWqrZClF/CrZDO5eUHZ5U7OrP4ZDD4
O9sxlT7rtjIk/WaqrlGJbCToL7oV1cjJX48XJiCaYA3Z15Yq+fuLFqJz1nmP
bDimS+Gal3IyIaWldt9KNOjsQLaJIu9xCUK9EFdxS4Xng7488YJZ0axfWyLA
dGVotzd8woK1hDk4H4xM9RXEBQOy6IWN8VsRRzMZVwBwfSOQOZOiG+FDyEje
5E491APScYIijiyll9P/fhN9Io7pHpH+VzImvtlqbQz7wKOqJuWZ4HGvhhGb
cICCJ4an4mPdt/gGZBuayBugtHvS3T1E0pZwEot4LK6YPhAj283QySxBbh2c
gTduM9FWEdRjlDYWImbijaPA1NcUYlXPPS9iH81Dv+MdEHMSHiaPMP4g3OGJ
OD7I8oUqwnUXtOLRcJRd9jpLQcKcvriNm0QerrQ3zeJgKUFl3rSCmnNz/ZDj
EoRB9KMpSqaWLBjYSPC4c+0AwESBEfKYEuKIUSS8gDJUjN8KPjtKnxZo+dMo
LtBzmjvJp9cI1CnMnyq24+MmwPhBEVsiwSP86UN5yaLKWklVFlSgo/CDMOKv
wOb9P0+9TZNQRyl4YUJEx3PTMP5ZomK45lJ/mazAykzIrBKLhEEDSFsdyjBT
cvUTXAocFeiSmbU9nm83qb6rEbrVq/HeAb+YAXJV2dJTYFieKj3Uid36DJEz
+OYqNO85AZK81HyEi2OcJek/3d9oLj5Is5zYAQo2rguiPZ8X3bXqpSXMrpRA
gckUlAMHX9AULzUyuzc0jqiXrlgdasxELtuynfUSGUaoD0znlVbTR9hfEfUS
6TCR4rgMwBoF1X5+gcQjx3kA4UWfmYlLQ/PxCvo0yno8CT89uedH8pZWGj21
XHgfgpstc3mgzf5hm+aoEml8CJ8118UiBA6peeChof6CGd1OC4Z19S3pCcMA
WiujUJ0F4KqhJ0x1wA7F3f6EHe9bQYJQD7YW/+TNS2mZmOwPFfZO/jsQK8Td
GibMNdAtYGmys2v7CHPER9FM7LD70NMkGI5ZpQpeFkfgaoKS3g/tu+dkV/Hu
T/0ADrSl/E4TTKCNtAHGosflrg1bKxrgkkJqf55yM0xyQK6bzZbp9wucbNJt
4lREh/gJCe08yu0jOj2BsOwIA5V9xNnmdw5Ybj9UrScee+bZLfyswMUIxkA5
TMlBi2vnQeaFy+LLXGDkeoUG76xX9zaPC4RQp+4VL10rnR3WXztZbBX1aChF
lEAkcEwxl/TosghcLR77jvAB84LVOetv4UrbdjrNyJZ9hMeJkFKQj4ye0DTq
/gpoBBoNBGOCbTPcedbIJ5cr9HQjyDKO4uOJw3HtHIStEB7sZD8/ER1D66kk
Jvb7N/+jAkqOtYtwQd06xBKWqWnMh/l+iKSXDVEPxyduyTjq3xA7XTUe7YM9
l63UDCdQhEmSrP+mvQcO53WuE71L51DFkkjtPPoOsoBn+ZAS5XFh21WsnJVP
gDtaNAhWmhcqgPVMJoLETlWQKfmPDDGEL5QU1qt4ilrRp9lmWJA4lsHaRQH0
QCdRXogucpPD//LtDT+bAGqnpNvU5xpTd5AJfr4TNNL+KlK7lLGxHFBLm35n
G/kTOGZrQ2HbBn1Ykp2vndZzwAKcviPEIYobLdc4kZ0L+9UErw1rRKZNJ4pV
FlDUGQF56eFkkKX9Y504BMNx0B26Xz0RcxfOOkZOhKgLppyViZDKZq/9orzK
4XjKcngkzMNnBNeH9Dws48eryOAPzCCA8uNuy3gd1foIlmVB/pw+pV+1cjOc
Amer7FLx7OpsUIoNQQty6gfhSUS2VVLF93L9ocEnGQSVqV3bbfdZlp/pYa8y
MH9I6AXO95rMYZUJMI0LTfypoD1kEaQcD3GkKuJrqKvPbgxUsOVIseinpj+j
lNXJgwmsLcATmYrR4e9jhbXFgV3hayQyri1MD39JA89vI76h30YdOIW3MQWH
52EsL3mQhSyUxH0vtuj9e/+BnqGuihcQ28vpfOlsvTYtJF7B7qKnwuGqixue
ruzeruRMJNzBJh4dS7Be4zKwCrlCtsl3abwOKoOEgfDhkoXRQVIwk+U91IK3
j3Me/TyfngYoE9VvCdw+omexJ4/yX0d9E9ZVnprkQn31XQKr0cuOlrGvnC1c
+T1+MvAKZ2gUMcSwbceP2xZtrX96wb2DQduGD3MjfINqoolDIUoRiX/CQT4l
mbUuwgxg+Er3QOKWOasoaDTmXnqnuvjs15/oM/NJUXTDk0HhB2nVSSuKs3JA
gdVUNPQ5sF2PJvvOTTciH7pHwoBK4dNnxTX6Hr8vjO73QanSOQ3o99WIer45
Q8yOc7Z813Yp4ni/fqY2tYfeWQpDdndwnt4RZPIlBapeR+HfMZVw+DCK5rD5
c8Zv/92KWxpu6xFz/WG79V2zBA/uQpRyM6Hhxd603oTfHOi50+3JvuCduxri
XivFUEWC3eUg9fvEEceOvFADLGWKgrkDDnx/rN1/YR281k5b4qsYZL3iiq4Q
B3zh/InG2FTbkA2Cg0O0ggh16ypx+muokJ0TnljQoblcVdEj7iK/hbcXsEl4
xQt2qeM2CpIjZEY0NQz49KpV07FeNxviEcz9qIUZmZjQNDffIzsCep0A5O3q
bfRBHhTsQRQeclfgWF7DRbhe/FSNybTpi669hyQ0g+d8ZfT6z+DKJXb5/5tz
ftkCDgsss8UgYbXfd/ut/iSnoyIFW3AM52BzFzKmarlHvG6/7yisWhuyHL43
XXNOtV4SgZ0H1vbFDmlrD8YPKSUYBZ8wGRLMh6o532kf9tmE/npnHKWvSPYQ
Nwr05Pf8lxCShsnnEU8+zFubBb/J7HE68gCZ3Xx55gQSwRTu4Nqg+tU33d09
jME7DbKrtx5RGviRYqPb9XJwZyYQ67xv0sMrc/ny2ynX5v8XolXYG2gy8ZAG
HKkFGF5tX7NN92S9q5wBJ02Lweh6TAWCfoOk6ReJdSlC+dkFcmqnkLgNH6Te
+t1jha23RDZH82x+3dr+Ly3N9INJrlf/pUGtL5MJRF53TeNBqjeXcrAxGSF+
zFDtufrcqSQqE3lkcBtmF0HcuWug0+CF8Plh/z7/yZ4DqqpjxuyCKn6wfZUU
rggJO5mZT0goS9qwgHQcpnrkxJhxG8xofdssrLK7V1nwuU8dY17fWNfuV3KP
/DPO2s44ZOo8VFB/lz2hNOQy+O5rnemrdbT/v/JlEX7mqXTjATb91waZj6dS
roZwLvFkchTW3/v+x85hv6fzIgzAUcscwtAp4g1pwminFhWFtWgQFZjmX7nE
yMU0/OF2uYGnQlbm/6i5DgxR4fyATfnj/Ur3iDXxNwzDr98GFtD0Be9fhgWV
L8V6gpgs+ERhhWZJSdApBKK+iIHyD5S+kinMrX2nk3aFIeZwSOBsiX0GnfqA
apIkUbZi26DiaV+4iEIP36OaysrssDWegKbHZXFBN+0g9R9jzU/ZTmb90hJr
EYzxEgxcn6zllcNFQ8i9lcTYbevG5WaFjMIyBtD9YxpUgax+rcDzMyA2GT2l
yhmMTSdLzd9if2AIurmCLPM3e34HIRW4xEgKzwsXQQzxy3ZOcCrDt7Byyl13
Vz4uupGczo0HerNW7IFttHO1bL/pptu3WyitdQwbrz9hW5rqHFlzw5U3D/wd
N/3KeaV2EPrqlYtiQe1rtAynETYlr79OZkLAvBpXXtHTKsgMM+GdQUE1sE+w
2Q5zklodApuqKANn5992Gq/nSUD59eNjOp3ZnQigckYZR0afKAjqjGB0W0jE
mi+2foRJJjySrR3T7RUzSqonyl2iDikagKLCsgLeNW2dawlUinTQCyhC0q3Q
KjSKiiZkfc27KfOOQFdg3bsBdHLGIzm2mXsIJ5q+O2B5Vf6qS7xt32RfnCH2
A7DBEjZJgCOSL4K2Z/oNMTETVq66OqlRB9gQntaO/arDuZjTrPURVzQulfsj
fyGlq2R+2k0Pjaui6jTjt+xBUh3/+wOaCfh2ivLoLEFQkNqh3ZRLHw/BFjBN
+w4/KsAryxLuH+1/ONvpk6q8iQFzoXvrwUW91FJtQL1LxAT4vSw8JgtXo8af
cfXqiMDLpVJXaOvf/iESgNXdTDLA6dziuKkpgTVSNx2hR7O7kyi+DIQwWSTh
JHRNZmKAwqo8X2v+0YBU1zQ+Bnnzi+ytmmBDhZF4VUqWpoKq2z4REbRnlDtT
FmU7IxOTPcLXML+eI12jO2kLpxCLpo1K4z431N5G2io6KE6PQ84+TRJ+86yR
OmrBSjLQT7MfrefXbB670H0pCqTpSQChduGZU1qR0sHPI2m5AR00uPfOjYm7
05+WsK0UDsvsIBhE5/j08yIxnK54j85JeurXHHz3c5ODlkVlnZM7nNFFEhfS
xneLgjzcswF8JH6HMWz2taZZWHxPUWAa4RZ/G6N9Qyo26a3i2CsIhfgfzcwE
8ekcQG5WZ4gZO7QqVN0ty+98NxvXEXG/SWUYkT2TbAh8MviTJDvT/oE0iZoT
YY9NDjnwtlQ0YllNDcul/MQHVPXCMXMsz3kyCjG66+dTIrAtLOZtDTMgL4Av
wu3A5pJ7j3AxMTz92rU3sXwSZU/PJVKvs9lyLlaPmIzZmUptp81UP42G7ErK
4iFJeWHX/BEDPaBeVJecRWX5qSVOEFR39B058SgZOiXLxc56s7qGkgAxliI4
HDLrsBGxHG4GsJ43ctjiiT67XEiwvArwyEUjQM8Na8Sev08qEu4rpifalTXL
BARjovuVySURyLSCV1WAh5zHy72tTDiDMoFe4MmwcuNo6LCu3HH8vaesR5Ep
oBCVj4Y2Ca5d7GkiPDbKhypLoN9kFqIzsLUDribFMhxShdYjRuhb425YDAqh
H/YtxgzMBcyx6D79jFiGbdmqGAjwdhPPa/eZm77xHbruoZBlNXci2/K1bdzK
XFAZuBSA1jpUjyTD64nbvyqP2PuIl3e+Prr1wTxfN406RvzFg0eI2EK9iCxw
TwJ9RzLOwH+OYH5MCImL6AHgLW0LM2Cgjy3zJGAmquHCzgC5FmHSUgCWUm6N
mCAyWMLPQYPH8tQ3Y1KBunWagNQVIx1RjE6CPTkN+7sV2X51okpTOKkUYh0X
uYIeD0Ap9wpDM2Ig8PF9jwrd0ePgnKP2B1VlXygJy2hs21NzxhGhjZlqZrA9
aevIhUOhDeg/zR5jGyHPiqP2TOtWjlJ3BdpRGyKIm0luQzCskfmv14emBAki
czf98Bun2z68wbZGadP/6fB8SiwRjoXT1vaF1NejoqVLr/hM7fT0spgr6b0i
oFsH7saWcMqw8wwphwOuE4NIjrGsMdprCZKqRKqw7F9x/mNB7uDQClZzzgSg
pCfcIyyT5g/wxZKwzGjTgBr0SX1T6H36BoFLaCihX1CTGt7UyadPD/g3shmN
TkxbO/Nb3uRIpgPc9IDnMjB+xr7ZYmdzM452GanlJOgMebZa6QmdHnj9tRuY
HCYbhE6/AYDLYE/mREovwju0qnI8FW16F4Sb24aHlbKtNJMupVL+oTh87uVF
NAJBLekkCm2plCzRaUv8iC4csoFthOdTISZDCTpVABD7oOlPnijAt7T5PkZm
J+UdfC1mArjn8q72e5UX1yG5V/7R8Q4xken1qyOV2J9mMM2uGHx3709hxsNJ
iXdU9DeDslhrZOE3t0HaDjMTfglJoa2RzKo7BDd9VPgBOnCqV87LdDCFBRp9
N/kST+IVEIOtRrw5Rt+r5aJRtooupgE2sH6hU0s8GnglqggPFCLnRzge8sge
sqoPm8YolapuzImUCcJgyXmarBai1PD+RSTBf12zY5ceTF43kkfkRmEwo2qs
kUnG65hwAouclyQ1cESldG8eFi4NcVOAClGgNt1P4gCU8531Ht0FPjayr2oS
8QpaBqf6pTU8DR866TT/Ut8Qb76hWPYs1QeJFmPW0+cGXsmMdTkcMF0qw/jB
7u/eWaClfVwwsKKitCBQxeJnUfDMTRMipC5eNRDGl4pBvB5DR1ZeqtuLUb/x
Ucs+sm22lSvA6pPx7Wt18NvxQNgnKrPWCrDcQYMdVbqTQSXWPsKvHymebm7Y
n7X8NuUElBztXdNXA0Dm0MeHZLR6JkQe54nHv/IGTqy0rvPSCj5l4FN8S/wX
eLSAIsS8XDgAmBrXFYPn1ssvPo+2jC2x426Trl+7aBkKnOK38l862DvuNl6l
qdSgDj7NUk8kthJAFICoBJvBdSLKlfqm0eRjfds3GwijCyBow/ebtFUDB+iQ
t2jY+qe/iwu20BSb4Snj/L5k8xI9gXnFWPbBy/oQ2ZBnuVpQS+LgeWuk9QLo
oDmAJ+RbTqowfqdmsYjjlB59Ko+kWTp5D1XZvD1SWATWWbvSYwGxBbBTvQZn
KWO4+uNI+xRm+7Rkayhekgqz5cYKGxzHuC96MKnqvQOVv9FENAzc7MNnwufI
EwayiKgYWOq1wvRo8aBQEY5ZdIZbLAvQJ/jcZMxzrKsusM2PHtDkcAIEMOeL
7kUfzSMD5wQflfqjfNa6wBkDBAIWM3k+QcyXGVmZNCssEmTtL+PUBD6dpHiG
tBFiyySVRxDbpOesa+HllsHGSlbKSZdn7aA1R/+NaIDv9AWhfzvhhS/BxOZY
7q5uxLzbZMrgT39GF4hsAsuXTTK/6d52U8QpWf5U2y+B2n2XJ9oJDh5mdVkN
rx1IaR0VWXKYF2Y48Tp9DP10uMmP/DPnUge8C5n4yHDOtdTHM5JA17cpHCI8
ZLMwJbkC678ZPKlA4o2oH8gSk9Ej/Vj/PpUG0w8uZh8uI5ah9+2JUNi0Q/rP
10gEtsO3FRbnU84593ewcPJaE9XrAIFypsKC/guMb3vZP40sxwFRUO8sN515
ql3LMx5uu2VpQsLKDV9M/XsYhM+BGfFTIVUnkJ+NkyDige5NIyZO3o6t69nv
osKIHmslmTGuZhxl+V0vJJQT37HYHkCXA5i3B0eUBcnvDhiJ31m/U+yPIYhT
fKoWZmLhP+MjXvCdiP3H6sSPy945JTZ891lVVCBw3wELfIlQF4ivfJDkiDb1
Y6WNwswNEt0EUopexxdWn1ic4B1WG6JBqinpAEuuV0dElQ7ZV0Y+tt2vGYlc
Dg559DlI3imfCh1MqeBNfJYEVQxS3LUJIB9bkUNztW+Ajiy0rqLNrRTS5ddZ
sJgItJjt8jJgYPtcn+N26IBS6TnbiD/4mBqx7oz0fHjyy4j9mgL6u+7QeNVN
lLqmjFDIF9KA+d4GwraIU0fT1uFqYRQzucDXLM62kLhmcqTmzbD/zlVsqabA
CeRzyW+zTVDuVCoAv/w0sNfd6oEFumTa7n4YldxOm8pVjHeND8/nk/PVKzWw
75GLVDeX9MTLULQqPr49aEw1aGPg7/sT5kop77/uxc7yDdTTlB/GaQ4hrsJt
xZriOcuTW2aG3OZWgG2gCIcOCjckhMmTBKcW6uanhCP0+LnN6b4NGDp6Vlnd
ieVxVDh2qjeq4tqvZQZpiXKaVsBcLbQhkoAkuD6jz8sc9QGMwQiewuFJ5Jzs
0px3CsbkOIUIp9jpFBuPEkr6TXWlZa332kN1tySddp2QYf2l9F57idb4OW0w
blL7r3/FoR2q1nNxgshxbT/FiBnJrezkI756aEJ86cP05WQfPwNlmtpuSNfo
hjVHAkAx9p++9dzpE960A3GsMo8ojFF/rYbbEnvA7HwxeOfFh7TKpsfJoyCy
p6aObClNNVHJupWdAbJ5+2vD7Iio1AU2ysRve2UUtZic2WVpq43Jn1apmuwF
/Cgx7xd+AsDOdaIQN375eI559CqJJenn5ioA736JHXHAGXzovOFtDN3krDmE
if77RW4HPQSWvDk1QH8gHt5n4HfEYSkwoif4pJq5OgY2VaF1O8o3LFd6GPYU
2GZVaWLsL7lNrw2jrwtm7buJulQxN/Op0GbQxKjuYJE8Sy8JrUr+GtWztNVj
yuiMrPm/jnHoYK8W/y/x0WdlNGy6b8xn8ZGExyaNPpJtwclTFQBmjWR3luJt
dPuJ6DEsAzbe9raueu7cqWq4PKpYekw8JQki71QxKhLj79KjchMrJF5OPcn1
/hHEZ7cVYJxNJbI3lD4dMIZ/Cnl+fLACnvy39ssdTrttvG7Rtik1Nc7cvD2q
b/HgCFTVwl+tPir5nAud/WOcCEYtsCZ4kUiUtHCJ+oZi6Y8Jgvjx8tDzin18
dYulE6HK674VvQLZNVE/Wl0Vvdpl2Br852mn/GXe9yMc82hoaqXzDZWWFUfe
Z3xTlsLHSdoN9tOPh+ajYb7LMfHLj9vlb9oGcoLxSQ36NLwkbhtimRL2mao8
1f5ivc/iIGW4xW2ww2EFVvk+86uShDJhJXWdJ1gUwn3vKRXW1gJgvUGIqeJX
fhJDisMkb7Sr9tWRgpW1SLvNBBK2i7SBPjOvRdYwwilnGiy0yWARKW54rM32
tC2ggESzUAjLvod2iearSI3XonPiO9aGjAGih3ke2Uox0mvorAY50F8yCLlT
NvIlUDvzv+bYc98aXl0icdsBpBShX3oJ3jn8dcuyDCHtQOYOW5TKrFgGSwuH
ywwlre95ALvznK70pXtYWkp4QLmefLpgKKOj2UMkLFVDmzbVU/FgEk86ERFT
pcBz29zYZoPV3XQRXMesYQX5JYizoQC8+DZvlE8BLNMHLtfGDXH1lqFqiFhv
CwrIz2YHrQ87FXl2DCvuw/WxtN485PrrT7LPwmTx1yQf/tn4xKuezz3adsJF
gJ48gkwylDktae1mHHEtFNCSMFLmqCHTpPsue41gW6x0eYktdVCq7CrHzr34
khDz5nSSMFwBJozOhJQNums1SWKWH4pSOF+xn6DdIRS3fyx02oThiZ2fR02N
HZJ9xVxUKiTZRyLKwT5i4P8wFjhSQQOO/koIxmEgUjoAyp0etR6pTjg4DiCR
tsU3R2oAYnPZ+VI2ayOg9wiz//vrdtVC6VgdnbKWlGSM10yl7rLWuWta1tRe
NKh5la8Oi4AKu59bmxBbZTPqtMYEExHls1TItk7R3PJA4zIJ57kdN7k9reXQ
tjJ76EeE88gCNbf8QRbva7tx5xSNrOTUWy+3EphJS0HvlTYJOggCg421CfA+
4rbBK5tGuvPLFNKuYJxbIMQU4lrV+080ec+ravk3lQKZbCS9EAaF/hLKxvIX
xsVnH85F3ftrlEWZvtbSrQDRL4SC1xZeX52J5iF7t3XqdcoPo62pMiSrgB4C
DUzD6uh5SUgHnq2fe+gPbIQ7srdveR+9Hh68Z1mxZUA/uXJySIB/OB5dXw/S
4H9SYHgaM3LMQsSOEZgwRdztiFDwKG5IHhJGorNjJ59/8Vm4XDZTTmvmqXjm
O63fuuSlfgJbvjYJlDN7W/FnmQ3XNWOVyE7xQr31BbPyJKsCM2lcac9oCODA
jlKJeVHCuvHnQmo2LzVB8shypl4UVqQSsYG4oTdkHVjPpxHdAfeg8t3mo/I9
G91/LxujRIA6znw1AAoNMmZ0v3sPK0aMO0GqnOuZFCZiQukXvnHAtKEDzB0z
k9rucIROhdUyt0npTUiyQyGic4hjnxgf5YEAxnYNFoGu7icDJOricCKNgg4O
UtT8e22c7ockGXDVjDjT2BzgFFN6OxSdZv/SSAF1/aUdiiLLT/AT1tAjjqcT
Jy+jgQNDHt3Mj18VtZY9GJZLHlKo5hG2wmNuYCVdcQxvl1nDI3sItTGMwATL
+m1SPFXYvvNMHkCvQmTO+D2WJufoDsjbP0Trr0+QZoNYcjl+W7PvF/sOpeOl
/jiVRIOgzagXwVQnaRoLpOoYn23UHqdJgwd3sZGMt7KeoIWGp4PAtbdH9lC3
d9saLzZDQ3oTbE19NISLOieRFC1YUA7Eg8jFq5Wj/NeCDxKaRu8usJ1K3Rwu
AoMwGxoq6PngYPXBZsM/M/jXqShDb/TG9LSOCPiNtjHfW46UCKnYWVlvf0OD
MOJGZ2E1UHjYwUDJAfntiKjdzVqsJOVzo5fMgYa27TLMfm9rMw/klDs0egux
7DTNbRjLTXt3S8fTQlvEgvzqX4B7fVGOZhQxVjsEJyci7VqqDvuTTA5xQKjn
T0NdinRPY+bFyKlF5GCgyopIT7z4WBZcVWtaKt5JZCd0Qqrb2l7ycQWR/+Ju
MVQ0aDl7Kkr9udXfoOHBkoUGGThNA3hXmTqTvB3ocXlWlruNrp4rxa7KAii+
m47DwDVpExMnnR3pEV6vOGSwZKPA53qYqNjtpNF+AyfAwnZY/1L5ksVFEDlB
vre9Ij6GxsGn1iqtMbJr3aTkUlw+CLZCcIXuyZ/PF1lhxKBv0Levph2ZiqXX
gHdbU0orXS7hnEMBzsS6mpKuQIf5KUuo2vRdn4+Q/lvfPJ2IErMJKU2QJJXM
RczUO8Wt3VZ88Uugdlm1WpKWZN2JRoWf4GqZbfdkOxKIaNvjO6mAKLfvxvVv
BOE00Q3MaDwh8RSdU3jTgn1zkGxQx7F5HkPMNE3M/WMbrXN7dbtB17ndqLBq
TL5CLNNEY36W9Z8XAkVim0r5kZtqaxmRHADRA68PUAEiWKiH8oUNlbGKyqJ0
tJE/zEtLZs3rbEI6JYc8+IT2JUaHUWhjst++nqDWpS7xAaNy0WQn+hp27ig/
HBeOU+KVWn/ezgQA77gUASz68TPDS992EexEusx/M4NgRDXrQRi8EUsrW+03
2Ci97cJAVosQ3yPBpyV4HVVYMDWwj0MjZqgMHeGa0Sdcgw7bXFrCpqtm+x/e
QlAPHDrwmHLh8TinqV4DXMQ/Ab2DQ3ZXpTVSWJt2tVh01kCAMmNRkkSwrTEq
X3bQ8z7qQ/dDG367BAl7NN3JJZQI7/AqdBPGmqm+YAuLtnEgV1VBTtZ3O6gW
CLKhkSaMCqnEEPKNjMg5W+c4Kt2MXXPqtGLFWIMdOUbClfrHeaSOMa7P+xbf
BMv+H857+/b6rU5vlvDSlTSUKAlZ4BnhrzU3PS/BLm4f49xYwu2i47kD0KdG
fGuK9rlUSWMlDXeQnV4AUvHiqPI9//h7PrZJqA03vGKIOWFQ7RWdTBKHiutq
r1gWUqzWJ77N6KuN9OoTTQyAAaI/DrF3VlMxxH8PY2Fj75Q8j+CyL7IIIkqd
b+/Mg7+FmRKnC7zPFUKAB2jFh8sdzHrhmzeDMzpocNkajOnsYsDxpxooBtAF
Ia5oEtS7EZTc+as91pXNxoZbX0kC6EphJ7YiNlGTQLW+3JTdPpgo/06e5zsz
PkpHxFmnj1Wffd1cYaaPxAajweTIkIsnRUKaH+gL9gl/HWFvdaPYRozD6CPS
6Sk9c5qLCKPWEalJ+Sy+LvwqX7TgpNHMBHTHk+byK2J3mOeGAn/R32k5Nryg
tfnnTNkCG0p2O0PaWwL3sv5NopnbRjHRqenJZKoj6mPWR7RnBUpd94tIejax
moqjm4DHmcb+T2Fj8igdmEP08rzG7pvSr70YHyd/RfNPJIVAx7xYMpybw8f8
dzu+vwy6H6C3uihwv0geAsFwfi97GZJNDI6w+75RQPksW3hHpGCTSDFFpNf+
qwuM1ACJc6oKsUswiCjN7hc4HdXAH3o8m7ARRPlCjwJxtDs8KXiViQU34Bpi
+PK+w1RJYerhiHUDIsDRQTabnvh2aUW4ALQlkxItDOSIoI9PeLnhKCZFG2yF
QW53kviyKY702Bhtume92hDAHJl+z/gAlVroBdqpxQ1zOdqk7vBRJmLwG+o5
77yDmC81c+pL38sMGwzgTDge+pRTUQTzDznP+CHWpHPyrtuUSebBfdLnV8uH
Dd9tphVAh5ytwlzbbHeMmhzEphx7ZbKCbadcyZKVzgGyNrJ9zj0rEyafe7X+
8zOGSBwgUPwVOVpw1iBsQ2O/qKyYpheemJEHg/CDoHA0XkUGCTqoCdiClLxV
4RPdgtAEoKpfRXcjuKq7Vd9iTsDsycjiG8LuU7bX8XjMzb8EynICI0tKy8oT
Zlq58+Bcpg9TjQdxFP6FN8w9oqNNZ/jEO/UQveqhcrWhqrOQxUkyePen69bO
vnxDnLMH32rksi8Rm7UlRCjafumZU3mMDy6Akx6Vul2V0SWyZosNZkJegEsg
C4YD7f2cm7yIvyJWuhAo/0laKF24yAEhXxL40afJNEveItbzeqJHSbpk1ESI
UFY/M5LU7LJKLrn8gbU7KL1VKrXeOa/AXAJ8qvrBq7QtvLeHPEtKMzBl2pBi
cEF8ovlqlsZgNI7++7VAZj+dBKN0M8Ua4gJpfVjjJmu6M+iPSWuBt3Hm07Nd
Sxwava8f6rkKjHjuVl9t56oeZ/31GfDq7dpMQqmdVNIbnQXMg5I+ZCQxOgl5
Q0SijjRh1Yu8khafash5aBXzysU/gw6dyLEZRUsCYmPsQhmkBT577lre/THN
CBkwC2CEkVvzCBMZPWxJH2Lh0nLcGIKyV7XFIB7pXTvvlwYzXQcvThLsoSX0
F4292g4sn3d3F75y8sTmiHAassWXixfUzgL/TQAEIOJb55rsRnCWOC5udmBY
jMztjBerJ1+DAXUcWUq4Nb1Bzg0AqnjdTntD7OoF97MP6hnTb6vBf7N6cNM8
lwj5NAwlLa+kckI7wuVlmibcU4GGKnjafyrNRVEupNTPJZx9nlvNqb3F4Syw
WwIA8e4YGNO2PF2PF1hLAjQ3xyWsM3GbxQDuNn4Knhqjy9ZLkQArhvaqKaOK
QMOnTOvCnKhcSbxvnpvZL6Z1QuVAtLa+gzfvhjNOJMU8rl31ea16w7vYxtqs
b87qZnSgHNNRmZ8/Pkjt9xVFB+cM/sYSZ90MyqYsW7hzCd99i8mFpmV/QhPq
4fbc64vSf+im8b7gBnNYTpKHerRhISIFKFF70MS6FeKUpGxUjTVhicolCJNY
Aq/ePyOdFUdIBfhEVjuc1rIiTMA3owHRZE/kbfUrEcD5HOBMaglwef1+A4zs
RTyHQTQNBGvdglK2olFMvJTlv28ADNylZ+dY2j3PrNIOCOHwcWwJx+zSvx5y
42pHGikOLGh0tgWSqjQCF1LfWZDMLmhKHFPH+rdr+LNRCZy4RlN7nXhoBUhw
gaQjYnH8L3up4HnwzJIHfAcJOAK5VfESiYn+dohx9EvJCD2vYv1dKo69Eg6l
J0iLgW/kYoW4aexZ17oQxTGSrP28idn1IhN4uD4f5D2aIwWklSMLJZCpVGMc
wjfzU+2G3/fiqM8oyCPxrkGZ5nYkk4QPZRCzUL1SCx6XA6fxWiSAn17L2ZB5
2yr/E0KjiLiPzVRUUDhMMF7kFOW7puSv6o2U/k8HYB8uGA09IBRDX/va1GSL
ecKQ0sHxzUU8puId+nRePAU67/W2JsW6Z6kBkEwLUPAxg7Qg6E+B6Luc1/jZ
01jiWwnBExhiB/N0ZWijqCIxBMEXcfUG4dqYItmhR2wIfAjzxuY28S5Tc6QS
ANU0h6wT0dpzPwaGu2TrMgfNOwSdECJxmyc8LQONRCFD2PFYMS1d6oHbXYLW
rwgYps18tzh8Tux7hIjea22UA6Dax0L/BDtUETmieRrumjaAIt4+WfJLQaN9
riNBvdeOKZwAp7r1kSJBQqEepQYHU4I2Lzn5EdYruOTsSXfFh47fQyVmz2Zg
Khb9zpFyf7YkZ1VARYDdIetlMfoQSfBt+FuW80gX6WbbGgyPxDE4XeYsYMbb
dS9ZOQujk8M8FGLNaC93P0X0t2svQVZVOcoxPjm4cOpnxGj+EW6t23XFfIx+
7jcFE/4WQAgv8nX5t82q2/ieyllpXS5zUBlKO/DvLPirBM5Z06ggnukAvWVL
KlHCQtB24XgclG9ZFERKO0hfvqcxc+wXA310bY30yZ2Ug4kwiBhqePH0jFx6
etHQHHL38n9IUdZLUPUe44KoOdqts1Qa2QmEPdCF8pmjQ5J/ULOcc9bhqNBP
+ZUyKNkmV8zvtYlyEhNA4YMKcI++tcucRad8FQnixTb466u2XPc6+BwtguTD
3ftHPudAMqo379uGHJpS5DBlDbjn++80WZwtHYROofXGmGuTtcktwiG5DTHg
cZO+IFxdcOQxS5Ut7Y46ZQdSX0ukOTAIc5PBuhInb+D+dWTf9JCGpK2Is6rY
Qat174JDN7GTyGXxDnS11oaOvIrCYhRFhUDPEsBc/P3hA04M0QT4UABaHssd
HdMaIFGp3D+MNu2zc7Eze1aznFPMf5Oxxr+lQLrR5U3f+0O2vFWedelprvbV
qohL+MuWpm6C6caFJe3IvjXQYUKs2tNiST+Kka82tCfXxqBbgauWtp9l/Lpc
BofqHOdIPlZUVCI64zF2RgM8w9vH5aenH42IEt9AdD+uetWb5LNrquk3sFR9
rgjTkz8EVRGsSB2azXN/2lqAwgNdGRslMFj3UFfXDDSLEVuZmz5c0aVZDNhX
TKZ5MhJjVRnt49hLiWKcuAfXhgu3Ec+5oTFpqVEQOuVNQA9r3flm8JqUbY5f
DNfSxNFFXvar40gwCL5bATEF+sPhBIGqHYZmmOXpXiAjlzd0K0NSRo3zjeYi
uVGZ9QDHXrKUkFPaHltsZl9dLntxAolX46nOwt4QmRVGFbyNySdlyWNLXBli
w+A2KKdOYS86ozLw2N1fU2lXzu8+v4AzkMKW3ocFTCFIIhkkUd+fiKRRSaAg
7wuHSbMPZcOSZ4cRriKTGeSBIQygpF8r4jx2DOmWvjWzhQW+oVQgArpCO2C7
kDZNhQDfP5FpizGUMExqwdhgCZh8Ew7osBJnYqTIP7tHHoeSXYeJAsPR6ZkD
rQaHRCu0w9Aek9ccavUEFoCfsnf147K1kf9ZxiRTg/C1lQ6E9kqQr2uLTExQ
NzZ/o4oHXMv3NBRcdSG7NgJ//97aslQEY+YGeZbYj74Tw9DuGeSDOTgV4B4l
U6yEQBoQEEiO+4DrCa9Ju7N/xpOYuoeTE/YbsL+b+oToC8lD8QMSPEEuI0ME
i5rgAPhdcgBcnLpoF7xcCdVL+xfiuP6Qyiu2nXlojY4xBcppmAZJVZCUtvar
CwJ8FFqUTMFFIHO+OlKc1kNvoSZL8fYA6/G495oKmvCbHJLHWcNnigaB32PN
4boB8hoC0AWbJJJcSWz1R62XA1NCLRnvlWmyYgA2Mlb/rSVVXGI5KmLSI1g8
GvrjtyK5fhkyxd53903vIsMUR4CNOUXoiH9HCp7rmOMbqzJXp2iP5lcnm0/h
mEYDJqRGGWET31emBVxc/1NXwar/O9/0PIEbRgSmgNv4qPCGf3fQ23JBhlqW
+Qpe577dd7P4yO5TT/7givyAlHiEDca6e+GtQTWp71gmOH1cg+QJOzlWQcVe
luKnBEM5Rnk2jRPs3nvhEK6xnKnE+yBuSH3Cmv3OroCZ4qGhIP3tYhfBH7Qw
H8wZ7hyC/H8zbpk185N/VqcrPt/Z6/bZBbYwO3EgUdx1Mbbfjhtxbb3v9uEL
tAIMcdUziqfF0/7klVeEdLd+A8lO4QO1FjJAM6vB5AfejEIdvO7ARcLYkvgf
Gu8TSxVHgsiOdNnjYck6qz7Srcv8UsfZEVDB+wDlGDCKEnNU2PZWPn/tiajm
KSJUPnDCn8vWrgFq0a/MNLtl1b9n4Uld6BXprkodqe3Sz/KPPiVDLJYPcojA
Cm5T8nHNmi/bNRIJafT6qn4m1cmQ9RLA3qJo80x+vyxA+ccTeGLrFFwaqHvB
tG8vMFGGuBtoYGi9W4j9DON/uIFCHoQjC6gU4PRehfpAmRh4EGWl/MgYZh+G
91Ss2c1gK4UIUSzi/mVJnzpZ8YzZkamSZLHpcUHH/EZhmoE7v9wGTyyy9ClX
BBsA7HQBonlAFPDx/MuzB68ph54AF6/VifxObJ3Pn+MV/mAOqLq29y5zGa88
EY+n0awwmDvK2fntnG0juHmkHcWV9beZPivonoqDhirCYwQsixVB4Nh9ZQ7l
OEXveozZhsV6YJq6muAn2antzCHdIG7ZjTbbexg9ef25udk/xC0RGztrX3zR
aFm54Mqs9t+5Mbt7kYLEydwz0wV6xAxuiohd7/1eXUqYZlX9T7STqz2ND3Zt
G3OYLdlRnnlRX41b4JYClxIvvTYQSefdbrtN/Etc2HG7c/8UziVzNOwbdoDb
/ajoMLlYtUY2vrPONTeZrRJ4pReBj7/WUEyI3UWk9IqmKI1+qo7fxbc3X2UY
3xVDfGXBJBKlThfSKQ3lcSycoWZwhsj65cvr93kfAa/CIYPt2fbarqJNo349
qDAy5BGwRN7SVV6ARYuJ6bQja65MNMYPMcXCcIr14Oeu23gE9/CgS/Q6y9Cb
RHSjXWUWhT1ciQP29Mo5IletJkqKqaTWQFHBRjD5zo1Xa58I63FZ6TWfyvsd
I0VOPCX4wND6//lWpuTCon6Z0mZD9agwh6VyuqKXKUWoV+Y9aPNQmwi5tx1i
nEKvf5wUkumpFT2+kN22rzk0m0QhpleNCHkhz6NxhrhFG7AJi5wDU63mudVY
FANF0rRV4ZghL4hpQpmiDUDSjhSa0fU5ZDqV1WN02IazfVm0mVm1RTKB5T/8
KvXulIk72uhJf/VCXAlEsmmfgDHfTU30XheyVesZ0ciylKClnM0fxC8aosdk
iMyCpd5gyRprAjYLwIBK3LxpDbV7YLxtWNdTqEHPoDVklTTEnD5e0njbSDaR
mVGunFZWDJTHpf1QYLfU2cLx4VZZTiucZZfkVfUh40fkMP+OGPyTpFs198Ds
qYqPJsIOloinuW36i4oVPJwH2udV4KnukQCpa2E9uasdJxllUD1MFUQr27H8
XeX0jKeFqKz1M8grJqoT4mkFDS0Of9dfGEXn0l77z1SLH4bt9hkSIB45NBBb
Qn1R9aXwcAaGyqGE1gc0Ss1Mp/SC1pftOLs43mskpmzqBBo68HpoXsZwmsK2
SU0bLDN7PJ2rIze0z/P7FHRYjXPsMW1V+kt6IgL+Lkv8wK64K0MVAXnlljS4
32N0cdLPrv4fRKMT+/fb/7y0eYwl9FgKWP8urqcstJiBI/iDBXsYs1KQ9LnN
AmuhA1n0WKus8pkEXGR0ejshe2W0qkmzFqDN7uThfcx4QGQju1oiaXCPm721
t4rKt76jsAVge/c0NOFROYQd0t3lktwQpzfDj/4fnPpXLqK56cKAVs40PlHV
Ab3gza5UPS7A2G1M65uxp0ADj9yWk7qB2xTvgtvxeW6434Nb0GyVxvT/SD/8
eYrJ0uPm9Nttd7Kk9RKBOOZkxT1a0Nm9bTZfGMPiZz1OH/hzqfkB8dPtuY4k
wA0nxLtmmsfrOxnrDFDvc9ry/N949ZxFRLl35GEoUKRWNfcefuqRpR3abfwS
5aJIpEBUKVwMb1/Dq71bvnQb6JPGVz4ye/zrYGFpSPCEyF3YLfsP+lK5ivCP
1Vl4G7DlmYCAACCcrsx2WPtUZmABfp6GhCy2meNekEI+j4oIPQaoQT4ugrse
kWRO40AZOQVPYAHN0CJYAwlWeEhv2IcUQ+oyXYGZXSqo8jW6F+lzDeM4q+cD
lwuFVM8TJFHm7BiZ8yHJA6wz3vLNXfZvwweNZMMtTcU2+cfpW9sdLtOUk24T
+p1iUTFGLlgoImYEQeXRAsogzMUhV6eVsGyexgVEHyfnIFsWy9JfUgjjUA9E
f6Bvs5TBfIyKBnL+bxIfStT5M7I9eK68sVGGha0dPtp6g7JH4GhZUKTREsgE
7NnqXPZ2xllGQVZgrJy+RE6Z1mL0rWaOc2/Lq5hpEmBmL6CtLM6SqVo7LTMG
CZ8gnLW7vI1CNTR6HHwpDFpJLS69HNQJvgSDnoorcJreKB8E89tPT6fio6gZ
aFNUpsuhDUU/8WaLNNtmYB5W/jF4XOk4B1IqxpWJE/t68YEj142MHigoRd+Y
5VigWW1MAkFTL+ZwvsV3+2KxnjrHsA/yOwIt1qrQQpTxbOwDT4eSpyllrdbY
iPK1NVzAh8NrsA4iAIHHVFOa+VBo7VgCGLuwbynyOuOjQzjQ5dRB4BznsK5W
6+YDFLj2D7zbouyQHRAwVazG7wi1XqmYORWu3FrH2ZWDkyieeTMPTH+6Ohqa
Ggj6rlsRhfIV6x6/oC2u+kWiDnW9wR28XUmdfm5dnUbzOgCuCMpOn7xZgPJc
I3M3UlTi2SHbbJO3VfQZG04ZfC5YwdcOZSFT8CJbPA5AaIT4sSXdCxWhGoO6
H6g1V4L12pxbipZLRbv8Bo7B/urQG3sR1o8XGzozwG3vT9WlmW4941CIw4Yn
D+b9vzt/g2cIxc2UsXcxZVVas0+3mxhjJbVxzL/IDCaIuAMfFjFSRNGyu/7i
DedipzQkJjPoDeJWyHg6EUT4i+4s2iJPlE/koVQDj9gGm7oxG1rPygc1ruSM
n1zTotMSAEi/8CL3dHM/20cSRyOYKlPPuj+9UsxxjBXrr0XtWBsk0/EX4nr5
BKfVJ1VE5PoIsejiCln42IFQGkhF7U3isXBTv9zeS1DwlHSv7j3btqoQ9aCn
rveBuCjI/ouw9EV3rKwSyxUGuT6YDJ7kceaoeCQE95ZU02AGJVshKjg2jZxp
mQnd7DvXOLFWUZmxzbd8fyrBPQ08172cfOS2PoKWVQqkIUY2pXnOidizoOtJ
8AuyB/VN7bkxctFgIVMu74HZw6PyRsFb+E/zoKsTqqAJzIhl3DZyqLOccIvT
IJbO5B5ZgC0jyXwl8WXJkLNmwUnm99PJ36+TvP8pwzP6wmwiV/eWWS/VkE/P
Rxin6o5jakPtjKY0AKFxrtZMFkgarYGvNgL6twYt8THPbRfzPCgQuQK1JtQj
ekWyHvlLF52TuyBk6hSvQHJQb+UEVPCo32ldcnxCJUD5zwj2fZP8/6cj7A9/
pdk/YEwvQtIfU0McbdL0PVrDwm9o9RMrIH5bxw/ZT1czSGHWA5JY7pOG5Sz+
qgxz6Usg5dgwr9OVnesD5CFZQmXIb+6ZQIHVnsrEz4OGWHa8igHFjN3Jsrqt
1+2Vw8yrno6ghIS3JALaAmcZH8ad6JusWm/nw1lr5gveEKR4FtIYbg3rwRYM
mcQd+EZQg0ujfKpDvmWxp32dfpVvyf/XDlhkh0ev4Octafaab5AOKHGxi5lf
w5mf/bUd5CLsU7AUST4tKMxwZl2/xwx1Af+HLuyoxCduJDVyvrogymP88SUJ
UW6yPD6yotwRoDVLxuoVTMtF2tD2s7ErDDUGSwrn6zvjtid74QUvQMp0UlV5
nCN7ATO0y/YX6Ug12Dz490eyDMkI05DtwMuIr/1FQnBFVHtjgHNm42MmRqIv
qiRyeL+VPsqRll9Okp3WU9jCte2ZEdT1rz/Ilo835CsQzrDRtJFncgDJYBdA
0bk1PANeFUHIK/tMWfu71lTw+yHYXxR57H1+jd+5DT4M2i8al8D5+iNcYPbh
6uwHf3h32ObATFtfpBl2Nxyk1Hr9yZ8OYu26zOqubeYou00OnozPSrNJQw5m
+S8nd3LHklxaEiR1sP+pi9YvsMtSTxQetRUoJF/vRH4oQranLJoSQpu/67DW
fSoQdeAAf30coLOZ5Vf855h18qw39sYmOOAW77Vb8YthqPxbpkGYnrFWWdWr
Cy7iUbzqYO/HfEFBPkBPLigfcgC2Tp6Pvxk0ihYBG0oyC37BAThnU1yPXbMZ
I57a7dhdz6ze07g+GXvVaJZck85mEhA526IYxJpHrnvN2lbKNdWQDtfYwFWB
y2qqN/xpHpjgCVNhxWlTLXCCwvc39fxithDXGGtKYjB8jZ0t5it3Hlft4aCT
PPkSnhocltlxd7bAQf+HMfEpySwwU4UijNcvCQeqQTMF1MdW9xIqbL76XZbd
UxyG+6i+t4zTvQJMvEoBCpgXsog0+3HBiNW1TvT/L2m3914hGBwYsv51Ckyx
61WFNocVxRGrX1S5ixki4qz8cNDUblRJ1EO8+JisdArSad04gqHDOTt5khgH
sFs0vW1H58aXZlQJGP9kPTpI6F+ZHGK2oHuuWOL7ZL/0aTbxG5LmAPg/+gih
M8+twiLU2krtgXOX4AM7UWRaZfbt74VUpUNN9l53WJemLxEDOJ93yy/gnF85
Str9DHqZSJS2l4GIMFupNDYBBl8umuV3PuIxyeELcBLITJMpMhxYgR0otERR
fwhMXRt6u7XY0k0z4Yd2wY8C677+YUqbgRyAKmK8f53xfDlIzAO4V/bzHoqe
yjGfTNeNPo7vCOSUzkgircMs24ceLoVjGt3sTDgty+jwTZjeN2NprqNk9aV6
XeUfBAObrhgTwE5+UkImbPFDQL+uHmnhh3e/Z9kawoph1FicuOdIvnANkmje
HLmpFvjv07cHS+ELmOtc6BxGZomLY8IjDNNgGTtHunUgkBs06bbMPonExwU+
CFrwaa5csOduoGP0tW89KmBuhLg2w2bX9y1c+vUXU0xLoa84tWjEy7sfxdt9
Ij6zs609Aow+Ki4xyL6Zcn+n+PgTPQkW9cpb+DaSXSrK30nt84he5gNCXuVR
ed3gpT35GoWTJlq/dD/2OWIJmnJBimrrL9932qlJdsHGC2wx63DxMtj5FtNW
U1jjajMRueq1SkbwL8abHMfQQOksSNzb8Mxk+qPemXXG7tlxCns313kw0djc
UlxxVrnxuJInKKwCZ32jHk1sEPEKd5+Zwt7l6ET3sP7nWNCIRBRjiBaBtgxc
ZJFdpCysHXEBWw5nYYNPVxpvOqtcUHYhFa1/edqYUzIGzBSZrarOJgncIYMf
ebztZC3Su6ZwfIb2/yBHvbpaSMuKvMjPmrmU5nzaL9aAhCImEOM1Go0ndhpf
O97f7jZHQFRHcjTII1v0jdO5+Adj73xyE1hlJT8HP6mtvPHw2Q69N6OK22o7
dKXXkqspb0rj/JF3+fPifarK03Xk46QIO5Uq8N7vNmJXHdU02kPJAgo+iax+
MUesV6a3zSFvaJkXvvBTeic9cnGHc6ro44HolDtqkgg4nQIhtcOKlZZthFxf
r4tLYcOOM+dPrIt3i6Q9coMHiPwt6lcWBv1qZUyZAZsp9zHoiuyYehhDxDRD
I7CR0M9oTnArNL1VRXJeFJ52pFqPwwDbeCOniD638SnMy/zvucXVnqVmza/X
WgvBxFvKWXLO7egT0M0/WTkpfFgwvAEXef00qZMeOmjQdYGO2Y6ynYrciEZk
5k4CXjNG84yw7YRQPZVThMHA6d30f6Gt9png8RuxOEsvG0CZyie3i0toddPM
uOEmLJScTzZvE6vYJ9ikxwX6M+jrJ7nz3k7PGIu5m1vriKb09UZYs3cS//oA
7vWCayPFdv4A5dfQPvD32198k3EwvISujrWvVkY0370AYgGVZ1/gpYnev1Ae
QO4XgzA9dYe3GrhvP5GLwcR5DO19Ty6t/RcdUHmwIXU5MV1G+57Jzp7pmQik
5cqQKqXeK3HTQDlJhzuqxUiXeIVqaOaGezvs+F86UjhNfTR4qf+RbbZsdFnv
P4/b5UIqIVgwFVCMVFqCTkwY5+G26KQFvMqHUvQaMqpJEsKbsziK0GjhZrUH
TAHJve3Gi704iSmx0MCwe4fZ/lxV87a0w82rbNpck2OTlJk5zP6cLRi0RIPN
IB5aPCN0tEiG1csQOs8oc8AaWaHumx/FHuPPTD5hSRLbHrFAEoeDkvx15aSM
/0Gf2QDlBJP0U6FJomq0DlUn5BWUnyYL5Lx9F86qdDJNu5ct7996sSj1W+HS
5Ii4wwUoyq1+BFkIVcAPIcg7kWEV9VbLjBiEPTt5mB2eA62IwDZZVVAOkBng
IcN0B0zmZIethnaCjuhwd2JJhC8FcWAPy6LtiQicYbEP3VTPx6w2J1jN3/KG
YyWUhiOIahdYhlQs1bpGh8N1Q9NCLVXExF3E3z4F8sR6AN2w2R6DQJkpFIvo
Jam7ZOoDDBd98J4SxgcEoj+GsSJNHypfhT8kX/bmPcUQNiRwMEb+f2zuQvdR
vPYYggLG1r2XR21MLsWTOyoNbkB0yLLlay/HzQtiHR7R/Mk/ebOumwOy8vTX
9HLT0VApG+41h6g3zDuY7b8ERWCPIGLpsDAYxPZtVuuz6pV9kQfRpwU64g8g
Qb57tjq2TOb/v5S5VF5GwnTrzZ1n7jPRIpVf0PiE2DYb1lzqlIfmqQ81cb8c
JN+3zUWMPuPYa7gnfzDCcy3+QF01kkI+310awtJXpZPBanak9PKM5pdjKh9z
6HlvEk7OLq+FAYa25KbmuxnznvwieQ8XASBxnzQbuWQ/iqEKpz2BqArNFi/X
NXLjzqvmdWIFaKCDH6cHlxhcILvxd3qrvlWVQlAj2FxkWZijI/6u/UTiqWjo
WKLEbxbOEzJGIZA70xxE9AoXMbrYqc4BxHHzGg7NV8IHnAJfiy6r7ELV9LV8
OGgUMdAY3/Ob2YMnFSr4Cb2OcRx11WSyDUIMo12Hi/2V3put5YoN92/swoqU
L549fFuRpKfHMVlLDyNz+WMmDUeoYDVc2Kk0/wVujCDaXa5RjkdzAG6HhRnR
d/rZUrnl18j0TQcHbR8AXVLzf5ZFxJ1oM5dmD30E9OlmKfKOp58lYRUBo/HB
uJBNKUuDc/iYWTPaeI2vq3/IldLR6+Q4e+19qanGh+C9//TNpE7JvW4trS8c
Yavyy4bDHFs3OzYnMix4WITnK4ldnGD1kE0bqP9IagDncQiEFzihs5g/gdtZ
fXgQS1zk7LQbbCYdEgyj34nI+y8UVKIs+2otsivD159qYwh5wzW41Dg+mQg2
6b44BC8+QC7ZRdiAwQbi8ok0XbnG2xHGfsSN0dfFRaFkZC8en4TxZiNCQyhF
nEbpi2rnjRMsogBplNP8p7ftrQN3zWKevb5AqF9GwVe7/eeAJk1psfNfuQOK
8jhPpMGiyFHUN5lZ2n0bcM+/VfFeHsQfg0ypfWE2VKnBXU9n4lrhRGR/L308
B6i4f0BS2jflzxHomngshxM8L0fZQ66u4w017txJ/M20CXcFyKTGDDCN+ZyU
SdDDugW85okL+A8DJmxpVoa+9WFjvmdv8CvnV0yTGPrNGQ3vQCX+ZRxsO0zx
JIRDZou5oDJ1ixbP6uOcskhfbno8jzpuCZJnriV6JFK4we5l+sVXm6PqI8Rj
gQVa7j9WLlMCTs/xYtbLETDEXXTf3GkHZJty/c3I7XhXHCMeGTwXiTmuQPde
hKJjPCdLaTSbfI9kW5KYSS3xwZa28yDpIdb1esAV7i4WRU+XTJ3wY1YlakBq
qD79tWFsmiG75Y2KWVNUgXHlXGyVbaDrOlA4AabEj7QsE3nNmeNKOCqfPrqG
ZuaYYniihaH/uy4VZNDwj57ecWE5Hx7lD5o/Fh89T8smcqJKyQSvQntJ8nMp
WvkMs6UsrBIypGscnRC+nlE6XNMNCfVZni9PQoEdnV7aXBsdZ+gdq3nVTcve
90hAMNpjVh8QZ+X3ubOykXGmWJpjAE+599LHhTuN5eIgDdAdUBLYXyn1VP+O
lVcFLLpmW4Sr+mEGzPxkyogDyNRBTavJAHCzYlzjeTaryc5jol2lnGlhsOeH
cRAAzkLobR+1FY7j6eTQvbQtbQN7NFWEtO7m0+mXMbaARYiUV7JGiQ8HAsoP
7NQFI3Z8ibTKgMkTdNmNXGCD91KVM2qus0ICUM/F97EmEWe+oJXL4GkSSscc
W/OR1oiG3InbiU1VZFc5gmSu5IvyqxM0N5b+Y1vxK3TIkVhOPqryjeT4rxol
5jGHcbdeOqLrKw3HHs8SiIf7f1zG17cTu33QflrbhbhpvY2BH+nbO6qcobWN
j9I8x6j2trWKeOj+r58cwVTd/5h0Wo0Y6A9mG2vrzbnzaQeSXm2QnCXWYAYX
wpGvLNc2rYgGf44eM/y4TiJ4P0F0FJwxGMzuaNpRLC19xBdB++6t7Z02HHgc
K08h6VXVaUgkJZW2xiPmaCs2m4LR5JdBFI9s8Qcr0/PvQfzG/X9JapQY8dU2
CuG+LZS9FEWYfGOd8msfv6Bx4ApAuRZQL/JzLOCHtWV4zi+WPpzP27ibxTlI
iY3W8wqDCazpCiRyOtVq8OdeN26/f5UAsAD5csHrOz66ZQyP7/FqIUpJ1kOh
atTaqj0BtCfwGpAd/CWbsdpeQeNn6HexWS4e8NV/hFMQ5wsDvt9jyizUaP/i
r81AjxUH85yYS4kMf/sXd3+0IAhaRMmc8Mu1Eugv5sRr+0sOokeZBvFQNDS3
yxfdXpE+Dt9uTsUPrvz0PRSUqLoPyzG0PxaT8c/+MwsGnpNNXSdYefvlcC2J
Kw7kSbifsQ9NqcqkgAgEzEY95dBY++UVo3tQ42VpPKGQAblwF5Y6OPCNXYfV
NdQxMOqUt0jsBZ/Sx2bE2suX8RvAMXnnIoX1YhDVqGrsTSK5erWuwBL1skyu
XLFm1XJd9Juhl3HNnQ1ZGrl7Xbxw+4XC/Fe1ukPrYT0StF9s1K4bvjXY6+LE
bRnvJsUJPKEo8d+J5XYUe16Ao/VUUxmJDI9QImsQi7olLJeOnvvv/kNJDdEg
QqeyFbL0UZudUwfTnA4JgwV3Bh5HtpmbpHkBAqEQ4BAfJlnAUqaloq957Z7y
h134dp+1J8z0gmPKAa3n1Icst7d7Vv3Xk40r5W+wmz5tK1oqso4LVOipn5eI
Rn3951HbfR5kJZR7KFT//Lsox2kYEYwQCX8T4NgPxmylkT9RGwGiVQgBXodx
KeeR/YcepzK7fxEsxySKkMmVzY7pHxxLiKd7FbRsZHr1mFidY+nZnPIKNgUT
1RWVk24QkfS+j1BermKDlzIMywRvQ4LUuiMs6rudR3k18gGdUQbkM7hmeGAn
6IYFEBvbjYvSzIsZaNaXDq7+RYfJnRPjQDPJMGtV7KKLdqwrSLFO2SPrNDsn
BSAWJOyDwcLCpV0OK5sAlMIkjOZE+a45QqjSDbhIYDpJYou5mBkyI1yi1SV5
qxpDfGHbwvHQGn8Qd7Ej6e+q0mAkfzTxSdqguwiV/i8z57RBPz5je8zIlH9H
qR0n4HiPW8S4p94APBPhx1mjSQUUqjDGnOIQBOjjRspiYWqtbi8Mjv451bRE
h32wkNMq1g5ci3dWPK63YVUPO/JXK0jP+PAW0CxInWtt1X1ULkekb7kykS9L
Qh761rIhJDfa1mmsOg+12ZxVed1PGc7kltLjbjAjWcMpxUJHSixaw0vbDBj1
v9sWkx5svQPJP0r6qbezLcTpbiyZzykk45E9Jh80AvBwjMnI/QObCKxJ6emj
b4grrYQSu0cRz/6XraTD9ctVlKtV4lvDF79MK8pjtRQ9cA9psFGZ0dYkxl4C
ScAbQrf1v5eXPhlroteQh0vdeBlIxZrsH0MK7NBdOxM77N7HZesLINXUbA7K
seMIHXB3k46E257+qp77FSOjYD60sB/6mVwN2Plq3flygGPJ1UQpJN6nAkYL
WwJ3g0bLeGwW4STwiU2jVQ9OYCO3Sk5MMQ6wS8OeG2EKeVQ7TcdVXsFakTon
3boAh8hdALjlVB00s0a0uYD/Zt7ETp48JSuPVBvlydpn91F0qvGEfVYPOZ/g
6J+rwCBf1aZ4FcczUMQPBzc5wZUbcb1lgl6z0GWNFryQOpWNYDCxvyyTFj8i
uxRtAFoiIW2PdMhklIWUIZJuZDCQQ30xp0x+rus4gqHrmlSKxY48XSSBF1qV
YpGEsMsb7AMuAqzFVdXgjPjO2qGtXLLaghYI6OvMXTloBmoEhYRCAv5iOfs5
7chjZ4vgaGCo5gep1QkvumBAMW0UPpimPDSZPokcAVv+I2/MsoFiC5/aH+e3
9tOHQRGbNiMd+bxuAI9uAdhK9NHMBSaZ23G2/eXQtg+WKkNxURpRhEKlHIFt
WKt0W5KrgUOtIMfm1weWg6yWsy9rsxnuxaDNINWxtWvVitW2YGpi8AXCDVFh
tmym0LXmCnXAOaDiDsNWwX+bMx2ftEr/iElhkLg08iqscOMwO5/UkJUtg48k
STTEecrM0YM6fsvzs1EvvUFnMJkUD15WJFgJNnjKHJuab1k/0s6WAFUeBV94
DHr8PnFf7e+D9D/llkNcDB8ZDhDo6TnKoo3CEMftgFqUTbOhlzZ15w087amE
t5jlrVAcqdyZmvn9/BRk5bDGvGTbGnf0twx4V991bi4DC2/cXfjbh5EwuE21
js8RsrQH2002tWJsy+Rsakt8y4Ytxose6hwUOLSBYAvsZytpS6sK2fehAeS6
XoJls4pZFOx1RIkBKJ1uEo8ZwN7lpUiXGQAO3+hgjj7FoY8RWeaa+5pDbnVS
1yEh4PAhiTt683VpiQ4Tg16mSASLoNxbeLjAo5HHvjGkz/0McAVn16Z1nXEr
McWfRQqBZJxZe49neyIsdhkEaI21gCU6kP2URTjGdF/cGA84M/aRQzMPqkRq
2BVu8T3USr9iQ7P0p8GfPuxAdTfqRBQVquPY5qbcxUCAfcaGmbmCp3oS4Ply
c3cpw/S/a1nXbmNuUgqpSy/1Lyuqu689M4bxaEFE7vLKeZegR6aVvCbmEigB
Wc8TGkTWUq6HUhklp0ZLWJ6rHqaJveVDyRA8PbC5oQAHyRw1OrxZL2opUUUT
YlhWhBj8mPIlhzcEfhWGqZaAun7Mv6t7z0cOl2j+flMGFJVzLB86Snf8blQM
aN6/KbjsyootO7jj+rWy2YMi3Dtx07uVgE+qd/h34st+t+1liHCmPsFeXkLX
HQ4obUteReFyw61WEsHtCuJ7G27qALFrFvWRgkDCDuDqUtRAZlZIHZ+bvOvM
MwtPq2uqEg5oZaAclANRV67Zs0d71twmKockK+r5ojjEvFvAy7b64E+IQQwP
5AFYc2jiI09K1mp2fTBsXoQ8cf9Z+qOx37EinoUElGTNty0fIfbxcxzzfLQH
v9EcrED88NRCaPdcHfEr8zp0GoTypIt6sqQ4myYB68vlYRgJufOXklmHAckC
Sw581hk2bjmUyHH6V5DgoA/w9mxNmA9u0GR+O6pKuOsNYwqwIl4Q0o62J5pp
ph7dZqso6Ni/E0nryZgX3IWN++ee+PEeHSSgCcNKmXnroXXLvlj+op6FmBJn
DRS4tMSSE7kEGpDRNx5jr4Z/QeANMgxYaNrJr4lABvZmxvEC1KmoZWg5RTQK
CgxuFJxqy25xJDl/RuTAElk/pYBHlsktT+PeQYa2c/JNWtJvVJCbZ0ZH3NNP
OK8wuzQtV0V5A9LkYB/CHntCMfPS6KQFPhdYV+5Uef7fXQjoqbc3DNY2CX1D
WhvaIBRP+Ka/hGNKjtnOaXyrb9FbMm94OdfYSwPPJ387BrQzEejMKA5CL/BC
h/O6wRS5GlVdhXqTgD2uDJFhpaZw30p1fiolJEDOqmqZgImvxnLL3mvkpzhO
KyGvGZLdbgIbuQrhedShONxYlZfLLs2m/f8lGvdaITyek+Ov1IDHHWKH99Kb
MNpys/SDsgXCFYSjvkFPtUdRUhCaqgkgmd/M5n0ypgq9StmEgy+kIroXU5jk
qI9jAyFzCqPaSa4aRVDHr7DnezZT20Yej1g1fOtB86PPpGgyPldycSXRB4mZ
8h+wAnu/ZPLa4YktXXWb0wa/x4oD3hGuCApAgVainTGxUtH+zBvDDFpwBemH
uIZKaNUUncdhJRBMvazF/2Dhq4aXNWnLpE69uxE+5pmyiany3xnzM56lV6J4
w62kku22u+61rDP5ZEM2qodX3Ri+QoSuAXLQeCDYP2Dcw1XPv06wLlyok6MA
l/zwAd7pQRkdG4QHPDB0jFKtsE46uYHAJAu2hsZcdvo6oPdyR0YL9y030LFy
eER+bwS+xYFzDDxN2xGMuSUyO51yy0uTYXe2oi5MUWlJME7y111ZRwko2Jl6
5WtZUJlQohhJ89o+2RF+q0ojvTMLLoYOZ6N5luvjLTZdlsfR/L6HAqBGHXIh
LInh8KlNXvz/RWGA2SlEEtOkFyb7/JkGaap7w6sXTwgF/2uoqbtP1xHzT1Lr
C3tKTolzFrEY7pyzi3YWLYaSz298e5DYFWf6PV2nDEUipauw9Q3yV4BsxaVV
FjS3tVDEYts4SeyMvtwNo1qM2+rC7QeK6MgwoN6Duo/ZW6EQw++bHdNrWcCA
W2pl4dF3OFCMilTCPxmvNPSxZFQuxPE+HEXaZJe6QIX+NHnT/SfBu9O3gVGq
7VOnCS59Wknx5R/4uARr92hgNNjH208JpdIq16ufNsxkuJiHimZz7eswzOrH
VH1s9ZgE+yMZ4c1FESMrHhWCxfeAxoi9oG2RTK6XreMdAdYw1eap00gNKuO5
6pIpRDeU4P7CIDm8JvvObroajy8cZj3WEY4gbRssNBkX2Eg0O9awD188UB/L
h5VwiBKmhnyS45AxS5tfz5rrE6WSsUR5gu+/slXc6L10G6WjMURFQkp4ykkm
rMN5qr2f4PNEbb+civziJ2zbZAZDZXSL73w/EvIdwV7601nPG9VnoJJDVOxj
oEIYkeNN66j+Gm5IBotEbwiA59b3sZB46qpzWoyGx7V3/HxGsJxoXFEH4Cn7
CQVIfkgh7H5CJODvv6hENhn3HXItwd+E1fC0aeLrPUpr/570zHNaUq0Rv/u/
s9g8FtDuzVafGwsd1yROwvHZjAi5jLgr7LtG2c5QRlJdUMnZlFBgLYD48VMZ
H6gPBwAvLRIYmj+ojKCn27+z4imSbVMmA09CrWGV6w+aVvyiS8IIwnm1J8dT
3r5TgZoF2d/9Jro1BIl69cDtC9pCyUVfpZUxlvgdDRfJpDsSIRRILObloQsg
Uv2u4XOqC+C7VmczcwtI/sxUjuCVzEn9vm3n3htGT3p0EFJkjCxcZG+7sTGo
aaUxbmLkM7pWz1gIT1B3pU0140OqXS9G/R48TF5oy+FyN/3bTHpRABQtdbbg
0jrL+uLMRQE5n6wsrNxjHIRl83Tr7eJ0Zv2862Kd5mPZ6bNlDtgjhVyd9xSM
Jy/BVsV3TTytTZyfzdQvN4SAL1LeeR3S86MR6n1J2pvwxipgakK8l9NZLbMO
9bCHwEw98npWlpmjDkbwo/eYXDluoTIHPl9Myqufs8hzoapXj73GWMJ/79/X
UuqsBsQdr6GRZTfMf3Jj/nq0q1kPWbv2v1m+zHfxrfKbEoalzF69HZ7jfU46
sa/rrjwJPyMXPUVEkVFjbjVDUY3zu4W0fyA2/6mBPMRP8haZ7Y1ILM6wsnX+
OHmsZJaIvc1hYvaZ9Dl5ttvPSPRyCTIVvu57iQune3EPsNH3nzJg+95VdA7I
I2tdW5e2p67YmP12WMHXqXxFoGHBaPjHQ9ABEAUDn1qNnQBIRrXziJrRlFAh
spht1h12jbnHKfhaawnYlcZfgDGiYOPYzh07NpOkYyVWzpNxhlq0SthuvsWN
hX224O9pYnAXqaLk4Eq9BOY97UnPD4n/c+pGALORcGjc2OMTGkSy8+me6WJp
dSN9PxHHZnuz3RkkETp8CdR0yXGJAYW1Bf0OsgbdF8pXRFRJEu04K3ZSyy4W
owq7EMIY9Ij0m5moU3Q0QJpKR6rNpciRrEjl5qW+qjQAL3nwLQfxTexG+N1f
Uq2J3eV9hIApjZx8dhvXAjUHL9Xi3k8GWKgKfmLFxr5ZcHgHnafCRKOAQT19
VwRkuxONdwf2tmobZ17OYM/ToYc8dYYl2p+jYea1K4TY8Qn3XVFwOhF9TLSB
n/NDTyaKpVcas0W8IOLDWjONbofYk0GHAiFdCGQSrHI6+c6XtmNqCGivhyB8
boYkWjGRAD/rSoPDuTRkpso2d8RmoXqluLiRy2Wzv7yTc4GOMRqVkNR3E9qZ
60errHPeaV0F/twTnv5DiF3tBXqlHM6CkKHXntiA46js/IwJpw0uk5wzqhER
V7Zs2lguUe5C8B/GUcD2T8PJ37HgPMgN8HEuL0aPOyKcEhZdJv7KYbO4ENI/
LP7lNNb42wimG8rKNPVJ9I0l+elKXB2yi+7dSQ2HL4vbirNIZSlNW0u3FBNb
MJh74w9006/p2q5RizP+jWE3x5V7UMQTCj6imVssTCrntcxAQPxuoyYNoB4j
MtY1c171S3XaG+tkbAx3acVkFGTOj6wuFCyRj0ZvAsRCHlmq34bUe/g3lbzX
yuHq8nxMtZWM4rJaDmd+yz4KNkfceSMpHsjl2bef0ZS/38O74GLVftio1QwF
VHGKECungwm2UrrliD+yu7B7NnY8SIEsp/G1+cWe2mGSPCgfhou8bOC/RlxN
f9f/CxlOqozQs9Mra7buRnz7jX8aeJxgFUh4JDpJfl2p+Z+Y1RPIThn4/n10
yG9KOpfE3A/jUIXYmAu4qaPyEH7rkroDGHgOP1niF+74VwLQZZ66BsIcb4L7
TR0AL3UskhIgpkxC51nafyKcYonPsxQkvEGc0WiKua3eTNnKleHyCGYd7p5k
HVqtd+ZYIo9r6YPkbuhFxJKurwzejNcg794ddwbirJMIaEHljQ/doJe7kGoV
E/t6aMsEmPoqaa8TaL94ZC5w+pqlWadyrXKellGBma1MJ3QQn7NL2UiMNUZy
fWDvijOa2b4fNaEzp14E82pI9rgiLDm0O4gkC1D0aYttDIpR+kQo4BT56uby
EdaTpyq2fSvtv7LUfe3+MNcf5VRdPDs/Y1/mBfJeulwHNeic4Uh8Lkgqj7GA
5k7TDi8Gqpxpb+/Z0NkJ8Jd0rZGWpzuC8odc4kZI1h3cgaBHq1Q6MLUJEzHM
KmJK6VreXoCYm+S041DJguB957YtBSIjs8zrY92ziNGHVAob6icXQnV23jBG
WrPqKp6B10uVKvs+0jg6dhKVlJrhD03IaqtJR/Wggtds7U5sti4jt6n6sEq8
OB+MPiVK8HQGgXjstOMmVZKKFDYhl2At4/o2LphGxPRNU3jgo0DQpEyVE15a
sTWaFMIHBLh73EwWEh6StYc5Rc2a7RWHfpvTK84aEESVW3lGsrrTLLRkPgFi
GUcLOQIifwj0prKTxrXwTgBbwnXTaeV3l0O4MgBiNPEY5hHJvem2w7PY2laM
urVINpiGj7GPkXNq9WBislcTc6+TR4oBiom+cL0+Trr1sHAuTF0NiI1zSUKZ
+lSAWryPIxms3AkG84kqZUyqUmvn6QxeyjhYkXAjq37ur8bi6klsW0GX340n
E5x9zSahsWMvTk+smhx4DyGlwhjFvL9Y6zva2UOH7SUbmS+J8a5Les068MVr
0FDpwolLrEsIUCdFB1G8HygGdXrrFB/hSuVxeBMtHJ+zfAUiMj4HSCY+3vRr
8thIrqs7ePGuO4m+EguP4E4+PTpb4s4yRro4VMfb1Gb1iEsIfqt9DPPjb9Ry
tW+1Ckapgi+J5sNVT1XcMY7keqK/oL0bBcSGCBSFvrMMgjGnEI32OSu2VxyM
SM8rAsZw8rid4yJHChdQFNJ0ddlP0FV4X2lb1kFkPSPTdHSiWAx5T5NG6MuW
Vn4L1pfY62QHqTxpNs8U8fkSjB9qy+FlCSEIkxzfe2rN71dx2HO3LrTdKBz7
UjZNBZGkdKKRcE4GSMB0rKMyKe24MHJ2xP1XeN0OI6WB/vzHNyHjEudCOMXt
O1UGhtgTTgxPofVBtwY+cWlCugfhLtUhm9gh2xO9Bdeqy9dX7eHtVc8NwjZC
N2zewdqfyX2IwL2wCA0xWdENJL2HG6U8mYZek6pckqkZCRmdF1QgBsRn0irJ
JIT8+g2aXYKLa3n4XSVwBBog4ElyN6Di/XmkrNrvlqpq1wPH++UV2OdZdicd
5klm3VTbv1FgcocfBfYO/9vO4o6cld7VfW6CJ9+5YkhHXpO+ZQoG3dfBdDh+
dTaQqL2nUD+NrUxwzgY1z0KZsbbM/X1tf34OPa6CPsdaH9jggdJbLSAMywBM
ckCfz1MJrFedQY6vJi/YwkZ+TB33Nq/mH7F0p17oIhas8olHX3DNQsb6BC1G
/SH8IYzyXgDzDZvtWMNdz4pbRiVyLRWf6XWCdqXLjA8xdf+vnXkABUFSiINf
k0g3w0BcpR8Bg3KFKkTmM43nm1d2ShQw4rAENLddhigP+3fOwcnKkjWoPQV/
RchJqWzz+7+zzIEGOcXOJe9welptceqMwImJkKHe1yBZ8J4VGCxMjB3RDLTV
KH/kUt4b4jUnnl3hLHUr4qb2VZz9E5BI549EySfUGeKTmrVfjRoayJG6e8oV
iQY4I+kmHWa7qLu8FsL04Jm6FJ/79IGd1B6/wb/D8XYONrNOql6Jqab7OUtQ
N90erdDBhC0nz2xR+TfapVVQHITzhXqXMbNNXhkAaf7m3rwuJoragkIFSeND
gSJEAjauP539Snx1q/Cn2F2kmLsxQ7JmEE1R+qkooCvt150K8qZuHhbK+0iO
gI4nZUYISds92DjDx0LKTzVaCUeCuVWZorfhdR/97CFgKtGLkVs4Z1vCB2OJ
nYrjrFhNDOZ5XRbzqYL6LkUHteanNokna6HJULZugkDzbCWtwwG45bI5dO58
7YPsu2fMbm9DzszOTmIvk7d4uUGB/D6FiAu6UrsWYxZO/+N6ExAWdTpeotRl
K/fn5u1aJ7Jd8HcsBajelJSRvRyzg7qik9xMmRuLT6iZFf2++BOtXejCoSzw
BMVggUxhD/F2qWz6YlhXkBrqqS/xOG9OXdWFbfyoBF8RrZcVSl2UiJeh23Tc
cJrfii14Xy8CBcAm4/N5iyIIoASf0W95/3CocN8zll5p83fSGza48nYpvcYH
mU5UBuYLNZcvzPI2fNoWJNuyyrCDAWgY8tb31j9KATYtezRi/QdC+CG4EJJ7
QLtClv9CQmEELe0vGfRtMz55/GQ6gnq6W2MFIJT5Tr2bGI8yiuVL01WcZkTz
P/NVm93VHs+Hl5lgeKEBPVpWz1vyb9CwHFSVu9XjlqKZyxdaWN/sH1f7fM/6
y8CDXKBAcKuK/4gy6YFtcPH22DZXB6jOAnkuGG0GrAvLu659GEtEAYE5xkXn
UeWCV59qRSa2K3uyr+Pbykw3Mn4PmhLKfWLS3QCYMVuD2W8X1E4LmkC55f3o
VEcRvhclEL4nJ/5YtVprofMiQUaJ+38bGH2//WjZVKVGNSOkyG7mGdg3MImj
CGwgXvU2wYAPXJShBtQQt0kMfl7Kr+t94Sr2sF5qUWDHgrQmwwP/X27M0ZYk
FjlzgY1d1dXIqf9WdSj439qy7aTAFiwIYSwmPQT2/xb548BWRHLnHLO8832v
EOb1V0/JQhc3b1E93zN87kYosscMrNE3fJLrfXo1i8Agjs9zEzhL8tvgrF9M
gemFEu/K7xNU5yH8FIxDl96rggJjMPDzpFHHXyZeAMgpgTkqb5IOMYSN/odv
aqaWXNDDNlY1f/QLYqrNFjJY7tGnOjqeQuMKlS8VvNzc85INOhImwqgdh4ZF
I54K0iYLflJrel6q5CnF5b5hObr54xn4yvo60m/n36Xe0VBwCmBrQLCnS9O9
IEQK5QYxtpAgdj3QV/hIenQhk1CDnxkJ435QD/APMUCEKqExUeY3m8LnO6b9
prhgHdZKyHZiKNzCRTti6vMQS1FF7BBAA5JcBoQNHrllQsRKk0ZwWU0D5i1a
PzT+nKNZ7fH1U7HFPLnED+d63sR17fyoz70QaOGBzfd02f7REAUvdlhfWO7y
P4P0h8Mvj0YX2P46xYrtogZP4UlkIjV4L7A5wuun4y46oCv4OYomNtNcLCxV
J6++Oy9wSDZPEVTpwbhLkCtAofmD+xfutF5Svzj3hrFo9sskUYPSP9VWxR64
/HyJqx+9oyQbxayHw3x7DGidH6mt++mNN+QkYBmRRutB8V2vdwwbwNSCKDEx
Vaf+TCDn8pjupxb6msvLoBK3PwMz76Sp0fu9D0Tp5SKKqSmNrtVerPOLWVzp
FGqMJx5x93oXjZ81yj5ew15PgDAzbjvulFmjDdF25V1j9gU9mehV0nHUCR3z
/24KLSXBsp06NlZbvrPuEDRjol6Yll5FozDbgGkWnSF5i8iboseSj4EZEdv2
vuNezNKxogu+XcbiG1odSsabjcAy6ggjE80yJmMBplqDHG5UYTKKmH6vVTIS
nlr6tGHUlfItgnkm27Ze6cG7qbb55ZLDs0QZ56N+QM3HFOC2LFQykG2kSWnj
J4QfvqlS2wMGEhkh91bgFId/NjLs6CXhjOVkC4xIoUGCcyrjPuMcJTkC4/jK
vgu0Ow/dTuxh+xOoneU2/N/p0NsKXhcB9D+ixcZkW0il/kggC23Qw15EPXQh
aDY3np4dvbDhYJUWeAx1+VgfbkAEL2uzthUEkQLQfAhw5sx/wc3llwFkN17d
z3rYV++GJAQYj5DDVPmwKsEPr03Hc+4HBJ20gIfdxjj+GtSABv8Xb4lHsZRM
lo2WTO/Zynh0uRCqlRSF7VM//keWQcZxTVb2p6wGvqDmP/7rWrs8fov1rv7R
f0liO7vL3WNGDyquEXluZYd0EiSbS4JEuQIu1wcms8a3wA/gxtIHZaSyzfhX
MacOo5123iK1h8uJzymxiqft8+aSmZf4omj202774HQteA/jsd4yDREDvGuT
o6Tky+fjC45Otu7omRnOxAeS5uH3C5Bjyy8Y2DIEhTah+HFlAySLJwFuX7tY
FldZ58sKamqU6kwNGc+W92qYmbNIFHfThjbJ7Bbo4vOp3Y8jrvIRCgSPRaT7
lQ/u+Z3CnzaDfR6bU5jJ7IY5mwj4zYgslUcaDCnLZNo9dM6/wnxPMcc+h7JK
oBtlP+bUlXfd5jZ5fTXcSLqXVgqV/dxJhRWFGXeMji6cLoB887mqn+DQp4GR
7MRSkVWxPazckWdxN0ffLM/u402g8HFLJuTmtNAAFc7TtXfP3xWv6uk6fQCw
KpjoX2oVxqLI4ED81YErQOhgFqo1j39fELV9Id4fbHJNg1mguvqogbF8mCIM
JF62Lk4GWAqbJdWSP2Om5AWUthLF4VVvg4dWXo/krQzcbbgMlsirwdxO4sYE
xaKZuZtj0mWsLqJSaVTQQ6GT1FNwqJk+DJ6WG/QdbO7rV+Z1RnYlWCPO9a4f
ibNwuC/X+Lri0KIHKolmBwmEJlUx7VUnEOMnUAuePJLAxcoKmSCNNcjDGonR
H1x4N1mV/zXuHuBzuVO2Y7YPFEsg+WFvbuGx/1+q+gtgLw0PFh5ty35NQzyb
Kyv2uuTokvIv17Ku9YWgfviHyS4vj2qRiCEJZH1rh55v/ctAnteuZOqMfhw/
yw1Piiu7gpV+O31n7ucc/y1DR65PFjgDzadVDEkFqhBsBqfd89MK6hWxq6uY
pM6y27Q+3bAVhD6BUrT0W1otkYpLVtcOBXkvUdZKCQYve/fs/OWDrxVl58yi
RFNLBsJYsbugy6zbL0tB3JcOtqTHr9KBMmjJ3vubOSw0K9SBAtmF7mPWKoz9
FrYFG9dnMa/gLrC4zSnUhZESslDirPELszwYGs0bJx388gdt/hLdHyBj+hFk
IbYfSOGdPV9SQRMgwGZSllZIJuotQfCa0lWN0aRn/4mVerwK+UVgCsRznKRj
2gAgCVCzTmy50gEiurYxOApQynszjO/VqN3IptLo0IMiWVZkzJBbeVBSdBSq
F9dnptKAJosCyNFDTn7QZmjadgtYKT17Zd9MiEHU3daiuLO4vCL54MIP1TAV
uIYVygrl7p3ZIC0iQyvK6ZVWFWS6CgWUyVG0MP15YAc3UOT/gIpyUsHfbOPz
MmGAx4PE0nEirGqsreJiEwbdQDNXA4yArTw6ROSbonApblvlLDYrNfO8b8dv
njjpB4g6xu9KxBQhp4kUkMrFTKIGH4w2zT14PDTYXBt8KR6Zn3+eR7KctjDk
BIcfnygUPR9Nw/IKDVea6L/+5bjSvQUReEca8Gaac3RFUaa/rjm1oxRtrUhp
lKlAJ+A5XFXNacjOATGqvkCuacMJ3ixs9CwKeFjoHGgYZ+SaHdS1Kccu3O9p
SbX3RZIuuY1Ma/A8R24zNRW08iSC3IQZAbTQT5Rx29Znt3+2A0j/aAXJKQd9
H4oov+xwVrtt6L7RKm289jBWnIlQqOoziweAfdXxpr7vP0wW0Mb/ym+n8iNT
WcAUcVSRtewddznONQtCWUcO21kEpkGCDc+/4jzrMZcAzyw6anvZKuveXeIS
94VTRWjzbTp5sgTo/NOz6IAHycKmJs4K7/pSKzMbA0YIPNtEciJGaP5erHyt
Jz0GAp0baYeMqQEgYxHfuVZ8ZYP0/HinnWRybYHEuHBZDsneFGTjo5yQnqlR
CyA4/yDrmsdPC4I9j8iG9RTGb9sezYp1975yex2gZoaoajTqnJuNLrWY5ylB
ZaJeySHRCk8isNOYrWCn34Rf5TB+eMv5dazXQMWWhVgSKA466lRC0bt72cLJ
2vnQQgjmFvlTidq6uVkSttC3cWj4a4Vlsj70qEZH1NA6gMzQvdH9vpILUQXr
1gw3M8WkZIaOH5mO6rmtAKtgXFM7K0Mw8j9bL4gu7g8rdB/d7OEg0IfRI9oA
bEFY8nIQLoMqdCcNHcju9/d1e8NoC0l6oXAQtorrNnSOfd/kUwwdMJcQ3PX9
z8kYszjVHPxKWSTpLrJkgL2Kj2TKF9LisjyfJErG14xElZyKzSCZAqBbvJyv
X9pcHWoVKf6gYvTXJNqSvIME8jR/msNRy6kbkoNs97qAQGP8E2R16a/v6huO
WFGOM86xE7tGHzo3xxuXhM3V2cbXEw2y6/4FbzPQGqzOnb935oz1uddwKf+H
kBhb5dzllejqBfNUBCmKDnzmPNJk0ik0pPgpPJX9IQJb2wvwxE8EOUW5FVcd
MVktY8IsD1htEDLdeWGZf2yaVDGLkl5KtKro3FqX5nHEhTprhNCO8lG2uinB
Aaan6ZcEKiodYdRhuvwqBjYmeXccy7ENRzLa1dHLMTh3hjO0noNPEMStX2IZ
J/D/T/IKRjrNdPoeFxtr7KzrkQkTEkm5k/HtHdZpi1y7a+bu/rXLgzqDgCN5
6aMLRQzIpczeCtrukneGlr/ZLqwyd1sSl9TjdZOHbwgoJbriCD9rxUGg20NO
Rwc8p8z8syEV1vpJQm9yp9NF09LC0+P2dOCYTYy7qKJL1pYVs3cdnMZWJooE
3GGDkOtdvsY4OPN4ND24MQDLbB2ez3jIYoHVbiae8knx8FSid9fLycNScvYn
H3WfiwIXDJ+vzvOS4uhKuvxzVoNEf+nvI1L76fARlO+Qd2vrfINzKEKPf90N
ej3ZxMkxWt8D1G8w+gxinwPS2u1o3j0mUNHwrKnILjDVAnR3mABvsQfNKPC6
rL1Oys9GA0CXShTdY4RxMG8r2WXOfzRjBePYA98b2rBT35pmUQSQysuKGoG7
n89gQeHJlnAhw3PwHCtxSl6sGyNTweL8VDwnjjiht66sm+jnOZK4ICwHrEfw
I9zvC8M59wUhp2BOzFlCbheJ/K5PST8SrycG0LzNYH3nsi8baDEoMXvA6Lyk
p1iBZU/u1NB+WhyTP+YyxMdvOw0MFuxmyhlvZURHlGNMaJ4naIAZu5aFLNuA
Tuej63ltOusbYWjQLuKQw7pLRfIqkAStBYNNI9j9zgV04j0e/fLHTXp4ft7K
Y9LBfcV2yNS2h25PCCSNx7r0UpVi7S08WovlmjCV4Ko1ZZ4mNb+4sStPwYTA
BQoVEgWW6D+WMi9zcMFhU2G8f1s8+UQSgjiEuA0vfwGnfjmk6dF4zMTusrqQ
5y/tsjsyrOnY3wcLSqmbvNK71MC32metfzcAIFP0m2M/7bK3zAqEmfktMf3N
vu4a9SD904rhiEiS3WqmiYfuymIhq0TqBdU38qVugWDOXdYS0EHS53NEzNHc
wZ+mDaaIZgTTp6RKZn1KttdBKiXPBFpxHHXkBBS2oJvPvbrKlYd0XbvHTSGx
NXzCipQ5OMSE13VWn1ohNYCmLTUUh2wsfgmQSDofGQqBQZTkxD/+/3Yvhg9C
W6+9ds9ww7PwJNuOGgnqrhN6PxAR4CFNNEmhTMYArPJ6UecTttpsaYfUMqW8
REdAZ41mrY9wlrPLTBbwVGBI7C/o551Pso4wsDCSlD+FiPhkZn3xI3MCYTpd
s0bIt/xFoE9sH3dVUrexsz2KL+XkbwJmpVeLHemUp/V2C/f8X85FwD2Y7gSh
d2pnblW2/ohRfqMtFWLo3lFZHf90lG34el7cgcoKmaFwSg1QQhqlblcuoVTA
erKSjr2y5oy8JvkcC3U/Krb/lAJUvUSoy0R+wJvQtVT+pKZ6fnfq+9kiBsfw
wNpWM/CxT8lEH1155R0j3Ni4C5Cyed6EnV6Yzx6y2l5bOIHzXPJMMgi8JjCK
5dn4G7W/F+zf2nPPnfEIIh1GnfVrMDoQNHNkSR9XnII5N+Wa8p1BDYom49hN
umaMFbqSYfLtOhNz8LbZTLs5cxQmBnvuLljh2jcz1wiDKPfBDiMQhIoZSC4v
m4p1O8NQEx/Obhu9wbu4lLcGNNMUR4lLUnA6M6VlRNKJshrw94/msOtV+uyh
n9oweN1V2KXZuFP6N0Nn0E/zDpTbroSxcNBlFHX+CdtLsuB747adhJkmCsnF
HuIy73gjecl4LK/B1rzzOAz2THKwIMynUMakt0r7X46vIFlWiSWLfoDOJ9YK
61CZ81VF2q3l9uav2g0md6vHZUEmx4FKCNPcoDzpm0R8xjYvU36WdGRoXDYW
TIjSeI9ZS7klN+nkKUE2vAjoScmFVJnc56/hRkaRQ1UqfDDnVN+CUBTbL5Dp
vzcDaliiF02fTn4aPEd9MRbZKwMGbKC9Zv/Tgj5HyTx3H2Q1JCDNdt+XpSuT
S1lUsK4Mg86W18HQ9k9jV+fVC/0RmpE1X/YLul4knObafhCimMka2DBffYjr
ll1SbSDmr766+FC12iTv1DdjOi5gRqFM9K2UYU2iXRrabr2MvvGeJssfPCbE
OMZdVtehdO9CrMeu2n92i9CEIjkn4Gzg1xLdNNggG+opoPK9pQyG22ZUDi8n
pQTwHjffMVCgwtGslxxmpRGgqApY8tqTbiQdCe9k5zfxmqO2HzmsrtdkCgkR
acjN/WjwapgvSt67RaXNpgvvTs+Cdo59xKyNqy+A9w7NV3tAQomR/CbJsuNR
eFxWt/3HPd+D4zmp89WmizJQPNsRs9R9KWsQD0EHwacTC9zBvtDM4fv7mQGE
IkB1QSc8oTU8EoPvpM5t5UWnRdixBJnH1iJgw8nFwmAuFv5AxkdaZNWvmQva
hhXBWUMMbUCViUvofjKMvSirn5WcqHpZDNhKs+EIcXXVt3g5Ky31kdYpW6Rx
ML+3p03yAIwUZOgZV7vp4kAtZOwDJHa9W8NxQDxmxKKiMDVzc1UBX5iCf+mG
yTf45INLo1wf7hpfjb90vyrO0X0DT/qmOSDtL1AeAzg+eXz834nMKM2ZaHju
dMTagp4Qp6R7ZcSykJ9a9RiMnUuAWoCr+EoDAxVY+HjOWFeq2llMsvLXDQtK
z82fiXhOxJIFuMgGLu/ywC6cHR80JJaBlqwEiHZQeiBPfB8pVzaDNxZxkU7V
L/5ZEclAFuLBRx43QmKFFtIAKcnlJEWwNR6eiG6Jxjzpa1Gwo2NgKrPRIxNn
91uBFgwon8iCCfBtQ/49R6ZEORfwVABDWMembGVG/6yq8MJ/IN+WCOWmYGUI
WaRktDAFxdzDcNH8/pYnPMbbSMRzQo7wIDKyyaa9Vlq5I/vQS49R/1IAqxDi
/9Ed7BB0nazu7A76xveb53wnVW0f/tit3s7NRToBlDyArRIk4DicyVhZeSEO
mlQ6N0y+RLmD3yJ/Y+pY0URsBRXHY5T7nnDdJRHfa3xqhoxLYP4V3JoRjCQV
cEAuO0SKFn7JGOekU7W0exrg1ddy+GAWVs2ajiIc19UWSeCMovzRKZ3hwOkr
zObsugKKIhY0q1zpYl4BpGC+6QZWB0saqRdjzzyGA9Px0PKU904W8LojM/HR
qZkpNUlQIEbmc/3efs+ysIgXZuecAAWco+OVwwHiG+ReW2xovXuM7Sc7r4NP
gcFkyYUOPI3p5C69Z5vUMxZA8pshDMRmQRCGKPdmjFchQw1vHf52elb2uupp
DFq+3LrZQml7590Yx1iRnBSRGq5niapsHULxaiB7rFWGow791IZEfAwbBU2Y
Ef7AWO5/SHO6IS3AbTRXxWkfN04fNSyuazbqM0Tw56lR4W8yAHzWP7ZL5QL6
xUWz3acQvuvGEklE+wB1f3q/rgVCBi+p8EDKaLAzcegJe/7/wHKNVfN/LYy2
aNJZvhde0+C8osHf4bDF/gQrAiyhOM6n5vmcKHv42+qjlWYGRdwyylgzk0mU
DA8rzF8ZspyPkK9eorArMNcRs07cLd4nC2UtLlg6YI4Qh9XP7uUQRZkedZ8z
pCitQa+5z7O0FfLcAuOtWRWa+kkM/avzTWBa5iElflX7fblklYzD9yNOZJw6
+Iiq8db5+H1JjX+qzFlonsCQi2nEJ8fNtzV7XvRCbVlx2ljGC0c8sEs6nQY2
RjyqMsrVB0GG4+L8g7lvS2V/WfNqDideSBfumWemrfrcX7xPSO0TqajhCf7H
5LW10NVJK9mgutxrOE0EMvrlef+7HystG6pE1eLYG2UtK/MicLcBStcP1j0R
H0EAXB8Zo9GbJeTDXWM6W/LZ/6ohuhPd3vq6KDeYG0tGlGChaSTndIRvpL6x
1UUITrfssqa+10sQokYUDzlH4OT5bc1vks49Iw0vyVescj/J9cPDXbuRfY6y
g+KCSZk5oDz3XmmccIqcBOe4a9b+a74kKxDqbtbO52Q8x+qFMXB3yzXXWCMa
oueQ3ZwyTUBSkr/8PlHRYSzMTKXO1MA1wGSXYkwx8rb6ghDyE9Wd2QIesOGj
+Bx0gXnDlJCIXfVY+2kIjo/JRwn0cgzzg27RbZr2hBWzMYErCWBrpCJ8uXFh
R89V2YDAgpx+17kK5yGRT4rSWDaVrCeze6Nx2CdntfU72vPZeKpIg+aZBeq2
+6G3LidMW1BkWLQxBS7QGPMDYB8PSGpxwcGhAN86KlharKhEyXpDndkeg6KH
GiFURlQ31ChGc25JjqZWGOac9ZosJPkdkbc0ElgxjYXMnyh42YWB+dIBXC/h
OMJYRuK2TFQdcTWK4gJLmxNFKd8Jpe1MCKrNFd1s4peGe9dZ4nT32cIUqaPB
M+2lXVBwkwSzB6hnKTnSaBqJiTRu9SLwOw4H4RM6WbrFfJKi2VyVSROEhQOV
YHfC+20PTjCSdWcHoa3lW1FHDiEyj1L/4E2iP+U7mkC+VNu7brtpUDdLjD5a
fIkDcs8M+lAT1M454a+aXucfI9jVvCJXw/+ZROK/Gk7/6P+F5RaZjsEXsj5r
f9a1BxHmScXqoe/hH8M+ZBPRrvnN7JEEQgLfGCAIeljCHBSIg7pNuVm34PzY
xZB6YfbP546XdZwuqVa3xPDaSX8V7zsLTiTufgc6D2yGscVO3heuEMOBIOed
hqD4KDUEV2nZivfsp8g0AaTZSdbCc3uX1Xi9nCvLIOWSIbZkjrt+E3VCZsaR
jqQER8wL3MUdu/56s31DbDMFWjqamwXqOYKIzTOxavBynvtPwt8njExECCMN
avyk15L9kEN5Rakdc1zmuv5IKhJS+Xz2t0aQPBqMca2cbg5Pm9tJMePnOiR0
GxLihXFiZUhRvYTG0ioXypKEL3eE3KVgtvGoZIMa6NkVjlbdzp+4rtG9qMjg
4lO4/aNwLtSxgLJRYdUY8PDOT5tS09TBvdY6luCylPBxXe+6G3KE7H/ddxhK
FegvVcjS7uN9/wHXhlVq1KPxVZoKsriS/3O370rvH/LHIjqSejyekPwpVQ5/
DWeyNa3wwdCmH6Fo3Prw0xxdAM6i3ukobu/37VIcR5JAwOs8oIxsVW+SIWvI
6GSXTEo7AP7sw2V909pBG5YqIKYQcybl/Us6bfasGdHCkfvZjM3cIeFpiUsa
zkJiJ4qBFXafXBNMuzaOAkg5iAqBD51PbFMhuoY8qNWil226VD8HOgv2frYy
xUOs4hEoQrShK7PH74zEycZTagBRKouFFFXi+fN/4ylK1dQm17s0JFfPeTNZ
b2HDM6fEUOczlRckwK2xIzJBL9/lmh+m0sOpkt2C2aWAQ2cGjzxjc6gMbenT
9aP2H1L6AT2/Xf+H5n4WTo2gBus8HUoeIuDftFQLDk9vaSuySJ6uuwV1pukV
OGCLvG9Zb4oNCy2D7Hgamo3a4SGAXNfEnc63023fJoLI7ti4nAr4KL+ktrAh
Gv8CSSCQS/WyRjDsEpMRSbPa1/LI6pC85/ELmegAXtXyl3RDpwVDrKWdE9SV
PkbsZwFcemPFx3XdQuDavt/lG/ThJDx+azlWXHNBTPqXaQwCg+kMjPK0gJ/d
e9NG6WUkyyye11rLhc9HauxZCTN//rjUX8aumkMgaB8NzkZZvxGz6H6m2ur6
9oM4yOVaXPtIrIHG9FWuuIysMLzXR40gNDu7x88vDiIOTGC7rP7PashGvqnf
7qV7a1k+xWxT7oe5KBOXSC7ioNohEsn1e2kWO89aYN704N8lgLYY2MIxduWW
E3iRqk8pE/cI6TcZPsrEMHtk6emPnZv2oRyMoc8m2jY2i9OcmjzZkRffB9IE
r+N/7g+SIBDcPWLFhtKPv1bP0kkH+FqUR2lxjkjnB0S08WxB4rPuDlEpvCyA
b7AgReQWuze5VusnPo3L7Qw01uc19RhgXQ0meTrhsAliN5dpNPFPoB/jbkKm
xLji1brwrc9x4R573m7/C+Eiw9xCbmbOhC5iqEc+GScZli3nRN47XFKqplDt
pjw0TamQT9svsXDgbbZlx++Kpd6fd1rC8maMAL11JJs7yGyqSARdoqTgCgme
f12oVdSYKn8RCqCcBdQVU8VslBg+DNwpxic3vM9dfGqkdFuGE9EVLahEAlzP
b8zgSwa+fH2FJRBW8jnn9UT6lsLZ+6c2P9314np2KHArdIjEsD2ugWdiScqW
vOgpNZDxD6jApUapw25KoEDxD8Swe5JMzIY2rBsM2BkYD+OUO/1sEFPKFSV+
F1r7xltWYnf+l9A76FPkdII2ig+6qwPJxCytEcORaTxwOmDnnqNxbSobZKvH
3Q6PcYwZ8xRaPySefWF4ZayGtfYcpCfaGu6T6Gpdyghl6Bz9kX73W7Bc9byn
79a/zJsqdgeQhI7v6MYqC/lvDwm9CJ2oYJQ3TjKSggWAntB6pHCz3h9Lpy8O
zhqXacPlZik9ICie0vbVi+CewTx7kbMoGUuX7qTZ+U5Gcu745ujKDsDXDAW7
S+d0wT3/SSXDRvr9KGNVRnLtJG52odqxDCg6pw5kyvhridX1DYtn+ZMOMo3I
3LsYj8+hoYn1UXKFP4qe7TYbJSV8XB5YHfxYDDDPwRCE2lrpRFEGjJEt+l17
IXcNUDQnOXGQZN2mG36XwfA3sZx5niRT3rMyXn/MKS+GnuyKif+HAVvtVs7a
KvrqmkfMsWZ30nOBbDTI9qNCirT4R9FApOZOu0tTXR08vCso7le57Z9fcMyT
PcEfraxFtmjJYwB6Elo9WCrl38wd0+o6b7TeboV9TVm1uY3UZO3kzUPef5Gx
meD8drNoq0bD7Bp7vWinzqxJPq6Dh0oxi2IaGKpLy4HtXXYaeXvaIyhyjskB
J/d5UroWKRRPFDiGIUmDX3yrFvzbR7LyqV7CJIe7mwQrgUj5j1uSGrOtvBRS
kUk3/XPCIElWboeqsG2pYi0Db2k/ZdJXYYQNe8QC5Jx1eIj3Sa5w5R9cj8DO
u3bIPna+SoO6xgTrKr+zCGs+JPmtuKSZvRQwf0UmkgXdeTf9denfK1hlJfYS
xwxarpjf7DrM9bWUeV89lP/bpxsFUWV08O9pevyt7yF98UIlvoozWo7rLyVE
a9GjrGZyz7m8PxeIa/pKELsFIo1q6Fi3mOe4yfaJQlnGrDOOeiViVt71zxSd
oGBGy9sDV+Wml+PYgd6AgB3A8GVLtLOf6Y1aYb9ho2DfvISz+YP5giXjl104
2Yf8HB9+W+T7ngAO0TdqUb3cBM2DcaAsxQFx3C/CQJi/V8+FUELeDfSkG+Rj
8DrAkkVSN72WMkZb8dwXgSm3AaCZxqK1C0te3BVuU+BwIfwqBkT+9rEaompS
h1IfADTuJY3maiAEltj+bM/ottqOILJsa46cs5mc3Q6H5Vfifav1QbZqS4aA
CLW6uODjwp1oTv2sY082wGqThudfaJE/G2fgvotlCdZqJPQRG5dcyqT3As4L
tNIzJiJQpyKj/dr+mBxSb0PiNsp76r80w5GMC3z3mo++4g/KCUHXGAfLis5O
22DbP4nSDQusimPpk4pA6nZQfQ6HNtEvOfkQv9uXeWKnKBqG1y59eI5tD3VH
wPfxBFy26MoYaNBlr34/8JeDb/G4YBWvDzelLj+j9uPEjNOV2SFdKTY3xdAu
hHboHgrkQr2tpM7DdQZ8na4gyjHQ1lGP8gFIxK+6klp2z//RpxJlZ6BqG4JO
FVS9WU0JtMwq86jxjLQV8+qeuR0Z9Ds2ywrxHErIjeH7jwDxZwFhvEmEqnd6
0vQLRFqB1GisD/LEqJ+o9qqfqs2PVxYkXDDc+vcCT6rDbxOCHKZjr+gZ00ch
QhMrvoTeWSDBjX49f3h/tt2kqG17RCuSI5dLZKX+q2PKL8JzTrdf4r5f+vFy
BMJBUAN3nS52VfRPLi1DKEo/5iafbHoGLfY3rEYKug6Xp5JWbhuptP8vKQIl
AcWx9FcdyqtdsU+GEjaj+KUwyElaJhgCjV9OVVLgDHJ2hDvqcomj2ESnpBv0
IGbScIAp9BJgrWnpuzveF8HhVtibkYhIUAim+/YKD9eQwZFev6uvtjpCRz2J
zEwpDIyp2czmoEj6XQ1EJTj47lMgLUFEYo+5/79UNHkSBB7UNb7/8RW5zsre
Ae7DUGnwoEWdo1gAk98/PBU92pc0XB9KTtXZO2n0STd7WEdP/bD4fFc+xPxP
ikceFpgUExD4rqzysS4L2RxfpxUWhbVtoPMW9WP7UKyC0o2LqvapGKwKHru5
fYMN3xpUO6P7EtvukFkTk9WKPmLflkaoOuxhjA90o9ZE3vMh8VjeRJeZgG+6
Gbt6ulgrX8Yqx0Zk70h/h3OFBlVc4XpvYP8G8RRdNacojrEtPABombYks34R
CmwsEll2TjjcBj4nTzQk7/rx5gqBv7SasWaCx7MSVHLkLJac+2qdkCPzKTzJ
/nkOUAP95n6CcG+HTw2JufVpcvybESKlH5IcVdxvMgqoQwB40enFtoEujKgT
qO9rO7nwly127fnpi8CFO9DKmxxngkVgOPp7n30qJTp3BX+Qr4n4WMwJWpSL
wgEJPtFFpWlyLuQfxClzf1p50aowMjRvgUuwJ/Ziiq8InQY5mIOZNum016Nt
+7fKoFeeLhHlbvSTctlSeV4cigpReKzbts4AIFXqsNC1fn099Ocvo5aPqCyh
w6mvi3wULBYQruTFRCGw0nJslh97UXylj5R7KeVUHBpAL+qJzNfVcnTeAXIG
cuHQNLau/qt0MGN9f8i5g2ugNGhfKRJ5nv2EHE4KpPv7hNXZHTW8+NFR6l22
RoCjqHW3gip1k6hDAjBK6eQmeGazEvtP97QRiyPBCPhk5Xwj9ti9MnFig2ya
ykwbX8wxKOAgB5WVtkmjkT3NMsxxEgniQtLSwbhGEK9finGulMS4TxOnoAdb
nSFVPe9T+HW7ugYBzx/aXACGYl94rvQY/1tEv2wfcxczVCM+j7wNymxO5Z3X
bv7ajU2gF0bbHxj+imtneUafVgko9SNCw9LGVYzFP6BIoDI+7MFbaOriXnOo
Qxph6Gq1W3dIU5yi9WGxHzfCzbcaj4Fe3ilSr34f8tLthHYlr+RxlABKnyqv
tdgJQRQZbUEv/Y5JM+LspXerR0ZX54HqPE8TbPbzAyd3ES4gMvwcAHOAjFyC
d/9tLpSMJ8qLBaMQG6s/d4YDNj1GcPuVsa5PJvQ4MVBwd8oU4h0FEsZZ0UFS
H2AtPWksFq32VaBIFMLVP+rQ6iHFUhMFJCtod37TEVy+FGjCplEPyapNxzAH
VwOEpmkNVzHaReP2ul7iy66D6mXJzY5LmHPfvIyXL0MbDU1EA/jWps57160R
G3t6B0/+6nYVs9qTn2yc/NDIHfqjNY93l5rVp1O9oMejnLpTOtNvpNxG5JbC
9YK33SNT/jZTgCV9Hh6DSvRffT4mafbZPuZB8b1X9fXyOqLUsp2MgtBLVbRg
YC/kBGnfhXn7Q+dxJKxJoWDNtEQwOz3XXL0SZihDpRrv81Rtk6+uzBQceklA
kOeWnzUWXLbFny3yKOEOoQDVooJXgCXU3hc9ISB4s3I6fRGR3MSGm4ArIXuR
iXWQn0+PwXGkTpETNlERvib/VGLtYAIvEk3DRXWGVelCzK3zYg4sjarDKABa
ff/5JriStK+6PYjDi/PdQ9LS0b+2PvSCk9aTjJ77ZDu2oEkN90qL8/6AHqP8
MHIZK1JNizFsvqD7OPiTbPmWSx8gfP9p/D4QTzgd6jQ6VWrS2+7PzpqwlOVu
v4zhuuqE3zvlB2YPcbqf0DIMAVsduNxzGE9/H30ebCmUxqc5Q2vimuumqXXp
sBVCy97WjdiTcXuOdj9FhkjXxT8V6+4V4BWbFuVQbR45UuHwqUlm3vy0C/1a
K/XfMDeSDT7/MCeJv2HSGwWfQNYcCIoSgKwvSzfGkjXRlg1XeHYzmz20h8J+
NyP1ud4aq/QE7VwVbeUaAXsKymJFh0c4l84y3+24r7jUneDP4YSJaYUZFaWo
rrE7T3T0y4XffK7B+w/dDlRBIo7XhEcpAWqK4LuK0PuMXdjFDNbnIYhdRPSW
NL1+ttIScZfkozNypVL0gU2wt/q2TER5zyUFWiMfN2MnaSvHwjmKHmArS5Qt
TDgasIxKlFQhspoKAYMCKnILzqpF3cLplX+gQhEnw9EhWDNBVNPGZ3GAPG8W
aEG3T7Z+h5IuW4hNcQKBZj4abw6ksba8wa0WcOS6blW2jOlAitsZ780HoR2Y
52bdTERA1lmPFs5SVJpV8IPVfPSh9wY4CP0NPjUwCc789BTgPfCInn3ufrzX
jutEMfHNVbuXLkdeF/vyBnyt+GbqdhqQzvm/mPLKa9sU/UQE6gP8luh3DIJj
G8NYT0X83YcUHsyfQb9jZpnJ80hybHfTBIjMEmIG83br3ZaW5meSx3j7PkR7
reIvOaq/kS2ItKA4xZ/UyrMyRX6pH5ilbUfsDPwwcglsWbZgjUpwzAL0NoGt
C2TGAHRJOk9nYkVwRnx8FdNQ9riLYyq2PE/rr+axdq/LDVTk+nH7Y0ZBWpy9
dTzn4ucYlaLqkhVr82PSerMTTjcnsEa8UzUC70V4wck3PzYpc0S/N9MHU+GW
U8stcR/W8w4yL1zMY/BB0bXB3tKnI//7NMDyUHTO5KKDl3TjLGWGoDNTbV/T
m26nBQ63PwZCXyTXRSCF5YczTuuLc9RbuwkEDgB/Y/TdIUk+ZdXfumEdHQJ7
Kuy+i3pU8esCZDpVoU6n12xBFwjoGC6kWxfgo8TvtzW9HW/vf6IVGAhl/PJD
bL5v8CrNaogbSJihRydBu1qcmkFqvjQnm9sdfbKDz2b/cPm+FfZT7cs8n7CD
53ejVAwShg+VS5UMEGSSHcgKn/3cMiank094rI65+VTTk4WotvvUcizyYWTf
WpJy0r0bRb9WmxVgRJhQ0Okuuoza1HJU9zSwY08F+MCQBjtm5/3juBaGZwER
SAGSxcB7o6uIxZeNwTt8MeCuHTK83HbtCn09cMAnJ2Jh8GkRYVbpaDMOy0Se
AHMrRLAZu7LuKK8N/rXl5ZjzoCCXt4pXllzuDXx0O0P81o34ZLCP7qZrAzjG
WV09OwKqt9fbNzRbktHwYI7sDszJW9Kb4h4/ax9M0r4aPeyeovxBaqjN395T
HDIb3E8qTHK40AQlKNsKfDAoF+HHPpIfFxzTzLmBYXupYIaoXO+nU2yIGgiI
0iCvss15j+R6vWaXEDOLKuYNmiguU3evKvKN8+x0Rfmd5vx2xPPn7gNo6VK3
sNyCYI8JdoDty5S8841I0VRaEDKgMgKPjnFdZVgswyMJ7A9pLfBRn2/6y6Jw
7yJsj6kfTUjFCgbwoi9/0VAm/eWc+KwUdiOlz9uPWBTPo7uTq49sRmJxAGk3
A6hB1sVcfdY/XO/OEBiqneLOc3FSz0mQFiofM543/VnC61q3v7IC8PMP0MBJ
P4gigS+EY9621Ueir5FhUOayuov+Rj7LNOdXffpzeQSNsVJfmhJJn2eyDyxW
uqJ01O5kiUx9xng0ChKiNyePFzB4Cym11fvkrh4BXfzpMwoufHrTkK24bejn
AAiBIuUevXx9cyazQMKDRDDGnrQzFAjrLEL4qUMeqAIhAPj2nB0sbq0J8Mu9
gu/tl3EImX5mCH9OFSMGCSeFNsARARsuxuBhmvvskjmbmbGANPLeoQkLwCUy
ng+KIrHAcP7ZPLsRg/8h2ZLLTe6lmZ39f4jATCe5/Ox7oFyI8SZnjKxxa0lS
RCFQlvAK+hpRra+JnPtauRioDeAMtgtkH4CwCMnoRjfQXMbiIdEPh9GIjpqy
Grn3ysGqauehHLhL0DYVDDtYQxvCKvaroDyMniXtkO1PjYiQR178tQy2XbAq
Wt8OzLGgUX/av1rzGqrvHfO9vIxqI9ViQ1DD1K++orGjzlvkGYC4jr0XmpfH
NtG9Up/eJN3jXH1EZSjXaMMEK0KirbFV2Mxpw2Sra7OOaeRBi1W3xPpwTYg2
MvSzCocqGxC3ShiDqZpV32hSwRHPXjqR9l9gKV/0OCcBdj2FjGZFT2GMh+gF
6IFIEtoYqyeTQ52jaeNb2YODKRI3EGzgPns53HMxCJI0t/Fw80UEJCKbEAxV
VD4yjPpEzg4IvkhW2WQekaQyE6xjq2SwBNbWA4DmD9xYaxqZ48hfByqTo/v4
EobjJYJtUBKPJ2732hjRnOPyxwDvGqHuKr1Syt1yhvVoRHP+BmSE1MffbVvg
G3TV46g++v1pf1SiWD6Kpm1Mej+WAvMrhpK8SjjTy9gmXNW9aNRGxVa30E0Y
0fR9Crh7GMvruTRackuYEI6XFg+ydtfJONIaapgml5IP5tV4nWy8Qg+eyMgd
LJZ6oBq3qNBeO0V4W1S6fi9oFSLDVmrWwOJVfDPU0CpDS/sbG23qh9xichV/
E75BiJ/I+2FYkEvXUXfzXgG9w8OGlKWXBVXD0z+kTOmIhpCw3aItuNsINIaP
ZNNkw8gWzspZCwc+ocEwXKasPLIyWJabW/dh9P1hANPVbNDI6TfVAeRuz+Mv
26r9cFNzwxYLIESeVTn2LIp8vloTyjr2pQp94EnX7bIjp65DK5YJypsisXe3
zGa5CsNXDvAMGRIr9ZTO+CCtMZeYqLsUBZvc/bNDUktUwVnmo4l9wIRFV2/e
99bV2KCrVjeFVa4zFncCE+zH96wYDWHTP5ei9mQpNdfGKZXYGF+CYUsJHWT9
yglnx0wBTH9nnMho3FYVN2QsfeaJDNEQkTz3qBLTu8/jTS+vQrEdmXYwzTOQ
pD4N5v31+nbqtYbLeKjawV1FT5EoE2CvBn9n1OgHoF9uOww1+W1MnuQkIEke
nbBHPeK6fIxW3SEwUJPz/Wi7N9l+XCmgoOS6wl+wQs3GkPqw4KmWIFqlu/Lo
wadxPhk8SUg7j5xQsz6HSnF7XiZQepkh9S8EQ0pX/+rdVeT1Eq3fPu6LfD6M
GdnbjfMUQU5hvTWlh70mMlZtHOyX9WqsywMqNkn6HCa7/kWWzUk3eAejEFOL
TfiLWxmefkf32T3aXU95Dx6PriMBtQ+RAY/ab/fuJUUQ50MI4FK98FIx38oj
UhCD3Mb+sARFY68dTU4b9yVATT8+rd7DaHrDJzwZwAFE0xQ7BfrMLS6gxROB
ZjpGkcf9tbR1whpI6hngiAwnlg2VR0qdLeHqfEIaKe99mbfcow+gCw3v9FqS
Yiqf6mm7J6ceGadFoYxCf+8BhaD8gY7OogowsJae7Pxc9yRDAtCIZfsP82zs
w3lYdNA+KEpZEbj3k8RwGlgJ85igXZUawEwiqSE8oI/nV7IpAxatosDNmdAl
wTp7a61ezK+4+1LNxhKX3i5gbKiow7/6c8aJ4vnR/0c37IT+0+vudN9l11/w
XpgpXq5wEHFwwRjpSGOrof6f+GQ3n749rop39OQoZGPfcZKEndU6Mvk2vz8L
b1ZQe/TqNJV252S3SfEe8WXkNf2F96RXVtgYWvdRjLamKynN4sEISkMXTlVJ
xMEdB/0EjQio6kitE4lcYzbuPFv0eMLIUJz1HEUt7ek2DdTIVhkin85b227D
esibOoDYQoc6vqwCbdpBPhWz0xFgbaZ6OiWkt76m+T/b3FLQSj5nnV99tJ08
WsNma1x+lFq4hObLYvNanZ9+5eQv63sYAE7ji1aw04/J/tQTy3p6PFcXHXwe
4Z84x7JLT3KLkqojSotEXdytKR3d70UIF5di+n+WiiklZriHbxTeMI+WLJMX
/tB12B7flLujYLvs66AS9nHzZuWSDgaJfd2pkyeafCQydqEizdVQYZWVcUOZ
wssBnyeJC5dMKz7dkvPqulfyNFUZc9tAb7CghyYqGN3zUiAt6NeltqR5m0JF
zoD5Wm7YJk3JYGKNZjRDrzpMt3mVrWxGduC3BUFDl4YGj5DiOgiHf57ggamh
e9mRD+g3FBaUPHGwb1Ezc7Dr2PJF4R2ZXxoYcPC87V64YPkpQ2xAfvjiQlOD
5kTy8zLzYLbKmJX+rIlFC6HE57F80SN2XWUu3BNWAbJnUC9WHNUZTUIzloP6
sw1h/+E6Yumyhd3mt5/2LlOWlmTZQnfxR1vAhFD7KnK1xz27GNi3TweYMDDu
quhghuuZgogD0ksR15XcWePz39NIugsuQa1PnOqK/EJRvWtL6G5KFDTU0U8U
gO2dQDo4MiojMmTGtaUoQ2K+AX/me5v+rRXUfHsBBJKlkyxTYNihO+Uw2KUY
TjKxluMfXxjEO3hDnWYRSuXK7WqJal8qPo0SpfDX4wJm1gbgi4g5BK2UTjaU
GcTiYyf/mvtzGymta9upCA3FaeNqDC2BcvxDOpRp5+wGdQlxeSXVUm/WHb8H
EcCg5Wkc6KP+f0VCazAosIihB6330Qph9C+0J8hEaMfeHW1pTFPbLljwvHmY
1Y4fKBkxaXQFggE1DnV9tKgfou+0tn8in0yvph02r8yAExk6oMcwCICXtutA
1kIGGwTK9hKJ9Fd9rY1X/PeTHg+jKfQJlX195P2Knbdw3/NspcYsMRZLP1/F
WpdltkxrkjHggz8P7MlGTfgDAsupVwQlReXRMeaIZXJfD5iBFS7hFl+CdtIa
yPqa0Ms9HXt/xAvIdSzzVKBwD5dHd/7dIImZcrkRMpgjhhIa9SgEwCo1J/8s
1dio9zM1IXKjNRfQwoYs35QpcAHWSG1s4VbKeK6i4hb9/6QY7eLr8q9lmyAa
FJZ6/QbfmDZSNSya7vf469CNMoFDN1X3SP5F7mPTEpKPFAYfQ+A7wBQ3yKDI
NxfFpTXJUfUdbTgbuNpw5qmS14TcqzebD6aOmKkZ90lhlJ220AqRJx9o1rUM
zSwQ+zU8PTlyTPP620S1b2g26dewacblTUP/A+p9ok4Z0hq5t1saqNp/74hy
VjL5yLCbJy4Hl/BXNhVHp3j69AMnx9OUNMTeanEyjadR27O7lodw62ANDhSF
7FOAqLCW/Ya6xVd0frIhghZ51bKtC/3HCkaJ50NkLoSIjpts26Ehbm5g4k1/
n7H9d+Af5+lq8l/ZaCJPU4Y256exX5qFNvjHjrH0I0k/5AJzXyDEuqCbVHix
NyHebzElHNsMfg7Ay68Ao1+nWryvw4nnh0dKMivkc1tuBcekBxxCWoizKPNF
l+vIBriUuGLuL1ef93PjtTif4sZqBw8jkl6dioDrZYYyGUicFbZrHnoA01pc
4yC5fHPm2W2KNqVXgKypiAv5aOn8714yy88AoTPBlNZJWmcPkVJpegsR54bp
A1yUrstD3sovH/F6ppHHPWYdQ9ip1Um1m1sSsGp62Gs9N7RJCmimmkI91Taa
cwgV5SbMEDJfyO7IPbaLgj0XUwOE050erqW+OYdLC6CBEOS09CwlJWgABdrr
qnP8ECWgeJ83Drimoe98pqqXbCfyd1KqLBucnccRdiRgMZVCVLQMxbZrRmSb
GzDUgM/5fb3wmwzvQQHOp2jS5SfDjf4yaKH7dzrqaTe/LyXqdJaMbKpGrUpy
/4uWmqnHVNb93k1CTli7HqqgNdW7crRNk69hbppmz9cw1ejtGHAANsTdPgIn
dpp2RNWnr0X6azqaSkPlOKlguipvfri5co+notyABcBcSYL3PpKWviqt4I9b
kdpn7ET2mZ0IoA5VeuJ0CzwvNnvhi0Tsl0xiVHR3Fm6X0+csj/0YiSmk5Ya9
avUrZ9O/qq5ZasUdviOfjUI1Dya0usXSRbYcxx6yUe+szyIfSc+dj14+iQBC
9+12l+MPq0GzBFwUZtrFGcATi3rNCofrMecP9dpxtM474Y9Op2J9d4SKSScA
bygXjJlO8J7NOBokGJh3yiohGIPfI6o8IivfmCGP5jJa1AiMCwuCFLSyuK4u
E+qtw0HrGN1DKZaZhVGfSTG8YtLAH0eNmZ6UJdR63iijZ0FBnBUAni9gxJqi
5I/scE30o8ks5jxzmFfCL3qtSZH8MF10nXqs8LiCZp5P8JiMQTHTgTmlhaLx
N1qTQtbu18j/cIMwkvH0Uc7Lh1DhIa1qUTLCUHbB5kR63jMK7gct4Nhr6IEd
Q2FRacvH940HIaSjCnuttHBF6mr8LOZT+CNF7e3/gWoKDzmhraGXlEtK+NpL
Bn3YggrODzcesqZGgmzg/ZDpj0nDS2EbpXhN4fRSOMPmbmNICknUBmShF4sJ
Fi1DioDc0JwKyoHoV5WEItWchvHzw04sJMkZTb1ugKHl2Y0cymrdeRURzGSS
KokrCGK/EenI5Eznle63DYkTFCEDq+1U4xmOYNUbtEJ9moABSKvvG0VcKeQE
X6nqwsqz2zOEoiNuYTAJ01nv1z1qf+dz+L7fADlD450n5ROn2ncSglPU581/
Pv9cWdZVdLf+5pg/YnYE3szuV5259cZMYOpgO+Ja9iR3pua4PXrcZxJWMNa2
1vcx8uUoNYqrkEPef6WufZDtKpfmm8B4XR5ZGkxWJ72FH6DZGsig5ZDO/LvE
1nxxOgJsThMqwMAoUktpD1KkMWwwCkN533PVMsfl2g3Qwv5z1cSSGZVEmgJG
jztsH8YBoPrlTsqWH+AbNL42uLaLr+w3o4KnZeGO6PGxI5/k8Xi9Q3UU7qL7
SBitkhEd8H9/iZazqOul7gak+Ot238gAStpRs38/N52YcEgfkZUHFAo4yeIy
Iyor2D7qZlHTKbYqVQogM9uZD3faKnRogEGky+ajpkTEcf0CkhBY+anUwJss
u5uaTMuGJ0CxgnJ0kIQ1WZsHRnOlDsRZEn3J4UeIswF4P6MNp0lACW9MJzps
nTw8P3crWQscxyGu/M7lLzxEifkH2/HVzg+MjWQpvRezRh0wqf6OZNOkbSwX
/snOWN9mym6JrJug2v5ZRP7XjGRDy4udDy7ygJZs3VfyOdHXsh3wQp9ba3Ks
GqzrPu34pKWRFWH+poAsVbslofmmDsNofvoXaiEJYot/PhtJtine6pLhJFaq
Wl2uX4fdsLnWKGDtKfNHgdR8rTTy2A5Zuo2ueEXpKjfW1r+YkBUyMAJg2Bfd
zmWdN24RlE1cHZ1mm0/sj4vR8uJoZ6MP0RNCRdGyEaEP1xf4lqBm2sDvLjQf
y5qNn01MrGMsE5SHa3P1U5z7xe/SC0cWK4+hOrpu1VWjgFlwwbufA9ujj+d4
bhHtYwuFentSp5f+GpcuByrZKjIXXAbRUwpSig/gf7uGdmEPMf+S1ckcmJaL
d7XRbQWcwT21fFD2ZATvOHAEgdR2cXcNvTNblbDR4AcErL5jnL9MquL9w6KH
H6zSuAeDMBtquVXCawx7x7F2yPYiIkE5EIKz5TdtM3iqcDyqNU4ZTiWw8Ymy
uMvduRQW8UiMPCdPis7ZtLFz0SwXH7xhVSbC5blOgg7GpAEZy3mfIpZVyPq/
SrctU3d7v+nS18OymabxtNaFq6/rw7iaANas8nkNCfQM7iATOzP0K46jfDx7
SCnTZvyO78a76Xj+F6qqNZ14Spwz+bszeJEn9H00VXM92EvZ++q/n0FdufN9
4wy7PP7wqIHhap+9qko7Zu2JPN4obQNx83dwocWz21k94U2hdbUU1BuzSFTn
V7lRxU5QqG5A3ourP6QQY7uBgQzmi2jhr8B11HygMd7aNcUFJFsBl89Fd9of
LCtgeMcaBXOnDB5LeSF+Wjx0eC33ZTj7WzmEhks/zA0IIXvxEh36OjCYT/2u
MJsTyLsL0rTIzK5QRla97S0m0SZTyyTNeag2gz3hArXlMQibVCTlNWPkO1/m
Zo6/EsZ9j78CAofTMT5P4sts//cQuvyK/kIRSxWAJa0y5iWc0tTA2+4xyYJ5
oj5QT2Vutr1MipicG8LaHlVBVl2gdnF/oMa+IRbtmOoMZTHZDAKBoraTgMxL
kJ9afvUJvlnjObCQZ48o/4Fro+lcLs94hAezN/TMOSVXdovjQ8pJakHxJLmN
DTvFv3z343oLrHynN5eVHXlbqL4rg7wvualcQPGBMxGo6H5icD/pBNt8e2v+
ezY1FS0ZcjAo00cUFM0Vn6t0DjiY81w1TABkFs/JatHDvctgY4VqTobymEBq
w0+F3MqGmhsMWptceZryaLtdZn+fp7bMpNtSUhhMQNlGPtnhbtaWEmrn+mal
T2EBv0i6u5RRRA8eaN8jJEkbte4+tquRhe5dUgeBfdKelj42HhGfl4yHFFCW
eG9Rbr4XSNIX4pBPzC+rizoRsUnXv9lFRGFC/KL4RaGWciDLGLnIBCtkiSD7
2o42KHGKu+OH1nmMiwr/73AEX6xmo6PZdjSKq64V9DCdeQyh68qQnSE+gcYq
udZasj1N/QnLEPVph8xeMKGwiqWrNOJNL6hev0bSJEZ2W0KkN4vyMloM3IwD
far3Q4t5SsC8lPQO2zhKhgEy79DvBZZLs/fgViImDxokXKN0EiA9wgTjpq6H
zeUOH6qTnsbmk3aGhtm7G3/V/wkLP1VaVjMCPEnkOiy1ajY0x/kg7sOUWCmJ
iqhot8vsadRRdZNqFkOJTTUjIbb/6lXrmIN36b9EiOEPxkEy0L5n/Hei59VG
6LjyibO/0uWFmVfxfen+CyuBEBD5bFYVR61EuyZe0l9uQ1CyWPSMSCGCF4KW
3oHcMJWHN5cHVOfKPq5lYw+/MYECq9Aepoet1XUa3UlLEIHjhUOuZqtwgc8o
gn3DuMWZWHXHlc+Sd+UkIpd12SHe3mBT4JegWV9vG8589+GsQTQiRdRUG4gp
T4IcdroJKZ8TWXQ/UHu0/DQkCghdQlFM5Mc8gi8qVHWdBMjorNACEf7nYhcr
bo/okfEQxyCFK9k5tv7I0F59zjjSYzMJ6AfhGl0Tb5cPf1pTgBZPrBkOGiJd
MGYwo46Y1HVX5b/UQa4NqL1RYbfdJoSgv2coynp/5HHjxg4w3PV0bc8vJSKy
JF7z8q74TA8ToznJR016r/PG6V46oYodgMm2twPp2PAtblHBaT7sGoexSE20
UvPwpanXQvaGWkjUSYxYdXn5CW+KsRrjx5nwPtwwuxBRGKLWBjqYYYMc4pHf
P5zQpBh3UJFiuk/OZzhPD0I65zAHrKr7okbYHyiqRiQcruM6xHYpu3ygzq2q
nwu1FvD0DnDXZyDKTCR5vCUXdEelnCWFXcN3uaVP1WidOI+ycrt87XmT1RJH
66LLksrN+qXijzgOx2eB7ahbePzjpLnKfIpuTr5jbV4LLcfQ1xK/HLJlbvuA
LfHj9XXv6KZcCD756CZ1x880+7efydrde580b16x9aUnJN5ggNX5T3hJdEW+
zzpHJFDBqA8vkPbWRBHkmEpuoGNN2tf5jJOtFPk1xidEpr4UTb0L2ohCsiDI
CGQGax/oUDL8GUBA5Dttpz0IzyDLhWkkTpxnb4gmuXqzbA+iw3wwgfKVnca3
AVHcN5owlhv7uej6dv7tNC30XscecaTFMpgp0qBtSfhdnP+/jYRssVPlb8p4
1IWbtjVe0E9I33HKtJvMENuh0XH+214G49HTUXBxFVajZYC9yn/3gLXi/rgO
PgJ9FrIHNTqA9Z5ituiJBo6ZpNF11kQlpHeLW6PalM46LxaIAlwOZMhQEuIN
j3em9hyQ7nmI8mvOg0hYFgElOuQydaMzv4ZAcdMo1/tfUuJfaUjqk3su2xt5
xGakOCwucyKD/zfqv620ffqPtBMx5T6QoEay3nI2hSO947BTs3tMh/SZ+61I
98RrofJxVC9b5lEik3f9NTf7TE2vV6GiZEi4VbAfHQ0X4YrSyq4JXpVN70xb
4QfoffQ3jbfSFH1pnMrH5sbyJ32piVVwTb9lndzIYRswtZkswsg9a4oEXDmU
/9a/BYYgqhlSbAvXXFq6Ev0Xb6Rcth2pLjY7O5zHxusTDh4Vz9OPpsPsfGf/
rY1REUU2G6Y00Vl8sDasRXw/890KyVaTyUePnD++6qvqQQAo/OGTLAYjQKpR
6xdEycLlGsxhq24AsxWfTyeBNsTvwRprMIwMJoRTd6sSO4F7kptcvGD9H0QE
2zuNPtgJQI3TfHZX5XORvHFdJ6NoWfm8yS5EpJUFkkg/vE2AwZaCLw7leGZP
hetExNSS50XPtv5qKjTjUSp8VCCm/4/y3gvk4F4OAVwh77ShCw1a0212Kyor
aeDZnIMndK2Wt3LhgHXxDLlpoY+moVqao8LZDixPwyRwhfJYH5knqbjLJj16
J0Khj2nzpOXcaSSkWra45uNhYwAs+RFCIuzLvbJ4fk3rcVqE0jAoC80zN7Rd
LukEprKTOGXSeUpP60HEUkGzIZXEdjKaCloNhwMygoFLFQ4OCzJ3B1UuEaY2
ELWjSb/GkK9Zn1n4N+nvCpAi/PD0gLndviuQj/08LL/xT1zciV576LEBpmwA
2l9TkRQXvome2o8HzFA2Xc0pX++M4XoDs2cQLyWESn9ztKEJpUhzVH7b9oXN
jBBILHs9f8sR4OdZ6lqVzjFmxd4be+6a7Q5jCVPixgDCEDQ48p44H2YK+mzt
VXdbdy1KPZMH4RYP+YxdQVy8PPMWSwfcpL9qjK9m4A9ieHx9KAcgi3Sz9Ze+
i/v3Evnnd44b/Jh6WH5zV9SM0js5GR2RNgfJgN5mQEpcWBFeMz8a53+IJpcD
1bK2xwJyZIrA0A1r1yX//bHw7DoUiD+49eH7JWcvLmLUkW2IZhtzeMGdEexk
vjqc8j0Tz8lsM6U58lhNckMjNhnsR6C2DzYb9usBkSjElq0TtFXzUw+ry3Ri
gN0fjsyfLhPYfmipRmtVNOMk2gLvcd9EMViIR091O7HNMWhollM4Z9BkgsCO
pcppSm2CUPw7XcqJgsreTMOAd1l0WvAmyCs+sUD4JECq2s8w2Vqv/1wp7DO+
u/+4eXtGouI9vpY4nGYFyboUDcj2BTsGewHo/fO9XrZVrCbi0YBPCVAg6Ja+
2H3i5GO0ZvzoshLg2/p6RlUnoXAvNTU6C/TTgD44E1zQMUYdWZcqWeyvBNfD
LY0AFLeKNZ6iIIfHO0rwklPoZKCBrrpg4SwserdgRpmxDRK22Vv8H0v1WOOZ
pdNhi7PUqV0PQkpwlTDiRX1g//BDVf4+frFqyimttozOSrTyTQuAYG5lO3c5
bu3gNDptBbcyJTV1aVuATPojPIK+j7fr3FpvUYjMnQ8UFS7c9jTQ3mjb2NkU
kB9ddWOV/jS3FNDQ9jhL5WrNxD5hfrKNEQ1ixjgsGrJ/8+IkUo9dRbKzMqp9
3n47uPfEe9eNLYf5lSNEN8TWIH1uo3/ZnYuJWJseAOjF1+OT9V13FEVFTdqm
yTq/1267V9K2eDndpZr6aZLI3c+IqRMHxHRlJhXbAX3Ib1Ug3H0HaNv9KkuG
U0ws+hQkfFwappzG8cSdF+xp2WNFPwmoiy4G6rotkjRRvixwJrMWH4Dj4WkH
xGPpBd/zf7cShHwDFgrbUFoEWgT8vYjr/Mk/Z5/iWYUEeVKC7wQDm6lUFuEI
a33vfZglC8/dAIo2aoOIG1gqsVr3PMjkmJiQelq+5CHTkgZL9h3L3ggtugCw
Id/1T4RZPGnjJzrsAxS+uyy2iCUJ18+v5OrDVJ6iZILs7HkSdCPNdmYyKpkp
UUCP4lShDu10nlDYlMOHdcg8kcvLBWGMX3V8dx5N+jpr9Xz6dg3H6F5eR/a4
fnSN5XXCNkaXjbAwlp4/feDnoSkYGKbboH/qI0mZ3kbYmKH4G0GlOHVOY3jg
5B5nTjA+qQTfJ1k7OCV2ygvw5RK2CMuMNU1UTHDjj7933U5V7xTjb2ISX0Ea
v9rYe+PeqSTcfA+unTBaWyEGsCtBeU8Sor+tQlQROk71lKy5N7R+opNWFYPA
XioDRJdhjtZr38ApdRrYxwuhMi0Gjl7BdBHMc/3LcMcy8diIniECjpbhf+N5
Ij9tumlyQjseOcN7JRhxFp3X9ou25Lap7vNOFE/ZPQgXl4u7eFXPkJkDW/+9
0Hlof7aFRLS0lS8j2NhBk8iMCdoW0sQS15nqNb7wMuVKkCf4/2jU9WLS/INB
YX8JEnA4H+l84Cz6SwPt2umYwdki7yjpdxQfoicTFKjBPGY76eb2tqU8ubPV
sJQop3A/fLNvkDyuE77GqEoaIeXxMlqkgAUU3NOzoHp9G1VX8Bd/fRjeJcgO
W8VhAHfv0Qv8t/f5WfAWMdiYM+RlcaZnyzpE4z3neZKW5f+tROyacZ17MsAO
HlrL4OY6RRdNdKiY5P2FELdWLrVylS9mLTW7kc2wLiONhivX/DiJQp3wA8fx
2ZGfKgw9lZ1fhmZ4DyGTY9XTNFaNAQMnKJXxofwo9NTCnLZBVo+JGSaujTJC
q8Nqp4LSS+dESFokTqC4qTOTM2cCFGRrKgGWRFc9TjmTEwn1pYK/fNqzSg8t
oUMoHdGzikElxihwUy8L2mKAmBluntTF75AoxVUhJm+Xsq0qwzRndf+++qSV
r0CVglAEtLYU8a2cqBSN8Af0+bxoFYO1w/ohYdcmY2Cgi2OVmBdVNw3rAzYL
5KZycRjQVdXsUjRr/qn8JWf31iJmdEbi+awGtY8Aq7NGlSHkjiquor2ciHTu
dz8f+JO0HkQAQpJJjwuRD/iTeY4aWzJdRygEEkdqbK42DU2uLBNB4mExHrdn
b8nnTN1HrPZ+DtWyedKO+nc/tCvcsKaa0LzADF4Iqs046RIwgR1CEUQDTRd5
9xMfA2ycwbOuIGCmGouWrDxfCbHfxCL5V6MZEB3SYRURRGJTXB9tsZW7hRP2
Gm2Db/ycbX9EoCT738a5ZFwN2YmfgDDSOv1OQnZNgZps113cNQvxCxpDLi9b
JCFx7Os6WvHESMpFl8Rwase+bg0K8zeMadgFMaRkOm5LBnbzIHWJZeyCbJ9I
niuxcDeFc8hdTLrrMnBaEN8+Xd+dXUtem4ke8TBVbgyUX7/xRrWYd91KkQVl
3fZIM/1r70XzBcWsVbHvNzQZk7ZKELXHjW7mJDclcQeMlOlI3BbfcPiybHMa
Y3tkMu2t5xqROFP0ool8y7nYnbIsOsg+sT1VFeHB4IDcKpr+tJnftMuWJ8h/
NqJvtv6lTAiKwGdCGtgMKfDbz92ln+cD0VuU57p/i90V81jYua9DfBcHgfWx
KBQBTqkNXcD11eNuQtTUzyKgO4JaVAkR95eOQUmBHCfHSxjMfFDdcKVpmFFz
+8pnjExSxqg4kmBX7ZJdxZjOzbVsorpCVR/4tXfZrkXFylwb1KrQQluotXBb
HzD2zaYASuCgYJ/GQ6K5ZEMXhymEP+KqDenGpWPOPN8Vp7bdITITDHPYqqNO
XKZU8Qs7oxiOVutAcNMKkKqghq5rRy+zQ64h8QPjCqPp0tdg29ir/R2hhusS
Vg0kRhEtnk09+WbFdIUctPe2cInZhDFxEqXvMefb6zkmUm7SHzMIpOP7pjow
7JTzTDKVRdA859TH9mjX0AOUxs0UDfGuyUBTDCdrgN6wsugogC7Gdmei0ZqB
lYFjAojKaVtNxUDu7+FJYyF6GkVjTLD9B8nF87jF3yEXCdIHQiDQZm7K+0zi
fJkATsz9tz7vfPoJdScQfBKI41KGiyHnxmFYkE4JJ6pmNFgUwrljf/bhX9A3
HWzRRi/RwC1AgeTW0nVwpR4AlNWxEslpGPuXnSZV1sup9uHZ0ltqb2i1huXl
FLGxzhHxbC2gUjoO5oyGzPLz4XqvdenL0/WovBWFBxyDl4VjVnz2UREoeLa6
0UeaGLxpCC2ADlgWb8chc7QTljTUgaWl5R3si2A3BIHGXVWAp19XDx6n2YPr
FJ0kjx7qHVYPHpEAmOGyZ3ZY5uHM1Sjn3ufRwR3ziWvnqhkmnjudC9n5ho2M
66YiW/v3EHj1BtkUA5PSD+YJFq5yarJrlIDYcuyFoLZxwRcW858jfJTld+Hy
jC0OLO4zEXQ1gLoal5uWVM0rbbYRXNnqJUZR3iaT6OFNtKOMWpQK1uKcCpkd
gPWUnTvAPvzPY84xGN7jddWmagpESrsA4IwmQNUUO2Msup/m2XoP0ng0GCr4
parnl8caerhHL6g2brBOZYft2dW8kneL240FxjhnNZw8GtBrwFD9r6Ej6TM7
wtlWr+vmGfI6JQ1p3wo+EO8391C+U74KDNH2oSU4JWo6SenyggqSJZim0G9i
/jeaOEWdgDmUN45RhP1MkRyGfo3Laz/9X0MH3/y8Svks0cUCG9L031VquQJv
YuCYEKGLNOw5f7BWxscLfiA/0bqhzVLCYTLAfbH+f4Ar4zg/sF506yLJTQ/C
8RsuLZptrnCkjbcFqnpriUzs9wJzOP9lIyIjgSljEQK3DK5S6v+X9MG8EBae
EOwMlcmWoUCSoi6S8/V0LV1RVrxDXtX73rgsbK/aDs+d8duV0W9oVBSjkXss
f+liNkKrzgXIBOih6yq6+H/dqaUFN3DSszd8n82dePcAgatLV9eDxZgTDKFT
s4ezhLfi1HgLuX+W+BhNA2ZldKF+Lu9OR2hrH6NwHq+7Dkc5u6ookqpDcOWQ
P6scpnOCFgWoqSRcxQJE9MNxnKhT1gF8rcilvT1/TOQwac/syARJIT0k9/Qt
vI8DKrKX47pKCE6vxQSDVtaOg4QYshtj3UJOxnqfr9N7Xekxs37lvUhPo7zm
54htzP4d0P537lwChfvwTicQNB4XkBZXDuHyshcM5VcboivzpzjAgkmg7m4d
CyTqE0TEn/O0idmdb9U/JKNm5kEigZDCHJ3soKqRiOsgAM/YGe3P8d4kY8iV
QNqfwWLnaJMGbNF36B9x88By/OZ7jNHFJfcm6XSSlOqokbfU9cbHDwN1/0gu
F80GH8NpUFK4hJBzglL3e2XBWbCPQtVEWR55Xv+18sJRjyoa+nZ3Q40cw9WN
5pRgNvfEQFrYWJSnfd1iKzi15OyqTR15nVoFfZPnvGad7mLHXPNmDlPZgAnv
o5yZX45oc/zD4wmv7McJ1igVVNW2eIa1OmKS/9v1wvgiZLgk3JCnApAu+wH9
0BsSBp67b1V7k054ilrHe+t2J8LcI4Mwz3yln2KuYOGYvdnyXk1QpAPkEcbe
BIihLRAxnsxJBQ79C8RJM3NQSU2hUClzWp0c0cFC848kP+myAwMtDd/L947g
JUdwsnZvuODScytzdgucegsizU8bl28evlbmcJO7OPrHr2xhKOE+4nQ1D2U8
X+GdawOBYq3otzISnuXG4otQAF4S+phnoE6Yljsi35QQhLnsJMaNHJGra+PC
bEkgYJ5olPRKoagCnLU+sRYSsx6zhBZ2ZsGvf8g/HH/yOrHjYKcLGLix0ZJH
UsqP8G9MIGsOPjChWLx3YggmG8ALFucELSTYEOEAtLAlcecMMf5Jj4qMiGdQ
7job0Nc4AKtN/cofD3SrPp7Qir+c1Al4aO46mq5ine2osLhSk3H/dyNrTSwH
PdjgxS/BlM2uhi65VVReUn7BMMGKtBbGXwH2Q7WF+hnKyj3vApXGdeBl2auO
03XEGZlHnaMwvw5C4YMJgNUzYqwDxshG/r/S0ZhJ8v+lo9rfAQAtum/MwW66
T58PAzLhby7FumuE6sgCoIG8s75svVSjwYu2lZGONjRcesdrNLuZ9XqWrd5J
rAR2MjAGlCDspvb9X8Z0PPxDQGft29EbZC2SMdD+5Ai+chUGATpxvj/PwRYr
9+baHvcGxaBrCiWxRYGbaui6COTV6c8d+vlbgaI576fE0Y4rpc/zA/sUwmqJ
SfFpLpyscWtkypzExP2uQrMPBZykKL16B/CDBGQed97B8+h7eJqhPlOsnHdH
6EXJWrQHrFJv+LFDUg6+8rPePpswDI9U9V4StfZCeDXChRJqWTNamY4hR2+D
tqGL0CXuAHczWaxPYKFTLY2QGb+0Zlvx4f42pUV1rNLDMvy9nvCKrhIMJYqw
bWhQZYx6R9jeAc8Qve9LaYQpyOp8dYH4RHYQhLUBB+UEM3Yu8l++6cOLj7+X
Z97uoN3H5ObQIjMHMiay+3Ug1pLIpkca8JIzwRoH0J0rSdrN+KNFcqA4S3iV
N5JqYE9E8vHcECHybRRP9qkFAgGngkU0PW+xdgEUCKhSSdymZErx4klrwC0s
tvDjxaujAZmVYlXh30JzlWGH+EjE5AYY3OvycWegYYrrIbOYoLryqMWZSDnx
SQ0RL4jiUOE+POWCSOtdi+MlrpnMrwMPiLmwKzpBFNp53VHHePOkkbJa5UpF
sOdTYNarXLMUpe5cdCZ972maisidvjTw63AbKf6ZswM42MjifadzgDVdlVgi
IO9qdmX3ur64rlqSSAQipD2eQviZsu1MG53J9pWddi/oLcQ5y0YmFLGCOpBj
d5PkEIrjHsooogWnF2VHzbXiMhxZFfdbiPxepGfjJ//3KEvQR8qpuaw/GdDq
xBXpHEPJkrhRrlP9yQbYJvs+lLFadpB7TSTq7If+RTPR1TDTL67TwumBflkm
S9PLwFBQna8gVmwg5sTl7QjCxg4FMm8DeKIg4l1qUHRnlQWv6cgBriLEVAjP
8dgUy5vFu1/gQS+75crUMmrqFl0Yv+odURjvZRcsGvIk+L7olNOX2ANK5JI0
zbij45LiFNWljWuhF67u0fU+W3n1bCRlBGHsEcniSy+yhHMc4MUij0oILWzW
qvGPuP4wDQS8yJF3IgY0LGjr+a0ChNBi/cV+oPIIV2MmiVEVDKdlmonWArvS
fXN6h+fK9zCASfAm3ji7nFctl62BBv61Xy2CsjK6uy+qs46xD/R5Gs3Tql3L
gMbxoYKXuyw+cD3u/RkxbHovfb0Fvmp9FBFW+K3mdllPwJQ0aoL0voUdmcLf
1CtBeQOAeC9x5SQdAf7gRmWIQ9/QyDFxLRNDt95f/Y4BfWL9PHHxvqgikict
LmBc+U8ADq+eUOtSS+Cwr65eJNeHqAyB4aswQPwGnSOumZLmR54cD3JFdInx
eqB0kApqaanrpvBTYgpTZQPKLvULGjSKykI4H4tnwrREJRWTBNBdXCTSlaFO
Q4FDsKTUQKOnt20ml1sm2TQqNXoGFKfm2q7gKbLul/pr9xX+U7eKK2jCDgHR
Kj212nqdKfE23T7MFrk23XA93x8fHh3GlSjvaxBmpxpoSFyaIYrQMS0hYMlF
R2PmEc2ubDHYyJ6tjBmk8og4oOTHjYqdifN87xQs3T5UsGBI/sGVOGh60rHE
sPo1RVD9WDj1Z40ne6YYTHwSaUBJLX2C/bKUnKORnXi9R1fnxEsIyxu3QE8X
tGk7cxwAK+Dut47FzGuKb3TuUebRijY9xtoRHVDcytaKinNZtbyIrStycHHC
BL0kKCO1uF6bDKI+KVduj7ETQEdp4usKBEtv1oUofES7HKjJ//EyoR9gPTBD
mK8KOpzr8QFjoqIWOYOTZNn+u27YhGiVuuLvxbLJFf3bN/iJ2rLcMlInpILo
GfXHmWAaryX6X0BaQ4fLM1qaNl+AIyn0GawDY8CqX6B7JJiwAmLvMc+QvFql
RBSEAXsJiJqLRFt/df5MncG60eVzMq4smJi2+m5+oFkf7K3UydtdIcoPXtif
O8VPrGU1gvMZRDzIyvoUpNypPlbpiGKVWPqP5aA2mTW+JzZjJi/QaenTl5rl
z9hI/A78dnzUW1KIIZD+2XT8Kn0ajtx9tJsuxy+5Rb7mDgdM7RJynW9gdoEO
0mcQ+b6WdJ7ssRbPudZpoECHicFItwvFly8qboWDYTDRhJyFuNB7+t4wxHq9
KRvY+R10cXlf/Y9BJhP6PRvMB9tzzOBmxDCrxnCzxpWA+iGCLy+UxctafpRO
0ZtUBNb6HYULKYP9e3Xo3ElrompJjKemzLe0IdDfczaqxa7ckYneYRanFGRw
GBRYBtUowSYfU8ZPzRTqGZ91zGRIG37RkWElwEFvaMpe9eIChmXiCtmLgGZq
SxuzE0M0s5D+YH6yV3ApWyZqdXXbh++pxXLoFOElKfvR3HOg+t0Xs4iWBw8O
trYHOhDNldz7GAE/NiC9aLuC5ThS6NdTpAfjcMKpIz8kNyIimgvTqjDQyRWk
gc1yjEVY4XszLvOV3pVzPJ+jE+DQZKIUWZSRFV+Lyx08H84zfnlkj2LixQjJ
fUcYEkzTnZtGe+ffOun5VD7Oo8VnOmbKHQaE+mF1lo0bjL7EMi1U9jxxY0ox
o3xw2/dint9DA5jLcIWwFcsDPEozKBGBgZcbJEqIgLUanlvdsNq9o5smLqKN
QsUV8O7MZKNeK2c1EdDEESAQ0WmIJjvjGZqyqs3wW3wALD5TT9wdXInAIa2Z
mOPjeirn4PRUiBf8EvjurqJhITBttz0moQWrs87TQd0MT16ItAIBeN/eDQZQ
4MP6wIwcnju561Nd/zQQr5fwC6jwv0FjE1flP7u7p7HVNKMD/q5T0IiA9mqo
6dhOvNuu5ONf097rDbnlNcmkiuk1v2o7yX0tB9yzX1OXf/E+iw6rRJ1gPsm3
a+YxbHn2SArZKvLAWHwghPYgF16m2BuePstfwA0cHAYjmmXVTNLw3jzthtXG
5WCIlTvAZZqW337Pykh9jIrS5u3LBQ7VJjAVjjgV8vJPzTu4H2TK/HaAxd5e
IHdBwwnWWQQ1cIBXx4Um2CmZiRPdqHHoOAlcUi27Yo5SdR8smNiJqqmK0lCR
LwUCqor4zCxNA49hTiTLXoM9h0nlWQO/44bUxB/Y0ly4QJZLWqdk9YG1eAMV
zwr+reb+TFYsmZgrwEKGKHTNmbLlxArgxyfOFtBk5mK9AmNvBXVd+Rc5v+BY
j1emZFr4LG4AwNEBZK70mvprZY956+x+Fsy0cpXQ1bw5SPPpmUaybtCMHVgJ
jVKjXrbN+ZzvFCplE8oeugKoEySZpPid5HEhP4Fa4v3a6pncRHhIqRM3sGa2
C7pjAiZ6kG/MFsgXwqRAdjAQBFAe5hz+eNj5NoDX19uX5WQIFVCYoePtClAi
m+32Nexb/lNPw/1OrEwlaWADEo79Q9KfkySCEOJwc9mmssVvZlMg83TQLyKg
TMbuTpxq0ynwoAGIvIWFLE78wEFcoCE+eV4NjuVqbu3UVuZyt/mF5KEgcrd8
Oi3VCx0n6h5DXbIOAI/8ULj1QoxaZ+wKBZVc1xkVhwlfg2JFnEUVI0aw+vzy
dWKiJF6R871HODnVTRauII/HYaFSl4cpd03CL/gI9kJHK5Zk73ftLeo1Eexj
3Gx1Q4oIncpRzl/aZCoCCqIUjPi8o2dYUNOR5kARwXUsZKkR9bSwven4PYZD
QdkxUAMTKqj2n2L6A12e89IiYyaxtdE1JPJEyQ8DIHN4/V1/B97uhNywb6FJ
VVtOyOewbim73wjYJdtYLRIHc4B3xr5kaoFl05gHE3JZE59LW7EmaUA34MSQ
XsDRwcedoi+5nU/XNVyL/bvP4vtLONqGnTegSGRiBB5PmbCZ7id95fi/4cNA
piLvs/aIJep1rIfwzIyNQIXW/150VNxCvRYFsLe0O8GZbFZnXATBe/lPalWp
YnAqgfUq4Qizu+Imorm2ODZhk51w7V+++Wi4cteiZ5CxCJQpnYtSPPxPsLke
Mk/DEuDsY40Gqk7n0zr85QtF6Tm/l9cED1pSkhsjaOBj99Z0z/sWwVGFCqKR
5DDDBUvaLq4VOvKiNe+IUC2IoK83CClvTA4qFU11/B+s+pmTCGk7bWCEhKyW
Z7XVkIZpLLC3ZxGm/myXAxT6ioHw1k6IjI32huJROQsU7ow5WC0gv/gKHbNr
kAGG8qdmALbkdGiCfqBgUUDsJAvZIG9ffh5a584LTkmq9OkkUyVVKIKpNWbo
3GuzAZToH2sXT82CtIAWnR9YMoG3p+BoD9+PtyCl39eR64sNU7EEyi1Q3vde
f2EyOcnSUOkd6SXl9Fw8s+19YXJPcTQ8dyUNGx15D7SRVLQDOidr/b9IkE72
y+gLM85WN6yU1od8Xch58fqjLAr2VN30+nWQ9gIgubkwGpEWMjbMPT+ACTIZ
SOU0QLVGup6hdjwopiaqXzDERTsgz8HmFrydcD9InIeylwp7CWpyJXMxn4lh
8XW2D64RMJFwqvg9q+t93qtruY4JkQVMFjkroIHQDeWqBC3hg/s2P9H/6Fc3
8Bcx1rF+NQgKSDE41fyFl7LUTXGBydGCex8YcbDydJLcT2KJkcmpsWrxhXNa
v4rSWy1n1ircjJd9lDpd4pzcuwzJBSBcjjrbT2TKIUI6/JF8UrzhKHI9xCb5
I2FcCc94sqm3RgixRxSBTA7y7tW1ocBT7aMvK7fkTdAroThbrSTCtExDVSM9
nYXGvaLP0gRvsnSXINsFop7TXs0jyRvU7PvfcCcp6KAmttB9zi3PamZyP2KG
F/Ok/KABnvUPzAW/B+477Ng/nuUdYvtTP2UuFPJ2VSRbU878+O1zlgbuRaAX
iIFV1zRL0ZtjjuehsAmKKchp1G+wlqnnSOsv70ltT3fZNGPS8yw0JBAQi4S8
2ZQiVijfNPg0J3lgu+/dHFFIkqnxkqVIdJY4JgM2pX4zI1uXV2TRZ6jkcLET
mHPCS70hLvtkdZvc4p/cLUfcuZDLB9TwDHPA4RLc9/necOV9iernNvqVJScX
tOERa9iny0w4u1sbPc2D4cJwDcigGGOyZ19VS+a/DvIIVlG4+AvzmzdJiYlx
lUI0snY5FlsV8vmQ3db/q3dhjPe8NGsAjlK9jGZqqjFIaCPzEQO+G17m9NvK
9Y0tD/MZCMI6Vydgjn7ipx0OXiosE/RX3YJ121ZfEgsVOgh461zfYjRDhSQb
jlFN1YlBidcGD/y8Y4fS9KpakoX+z9Ypnf6wR0cpL9n4zDeRrIrEXmsIzR8q
ttTN5AdoygiTWP2s+qDpn1f9lZi1R314Q328i0MgYQBQVVob1g9JMbz6/5tQ
tqJLD7C2PR6CT4EWCyrGAF63Cyf7+y3QN7f/m0YFcg5Z/yzXYoVxOC8DWNs9
ZOr3SrhBtGOijWFoEZUuP58gUWzMH/5DuEq+6e7kQI2X8j2VMuE5tWaE3pMy
k0+V0Ya2qPHqdapR8vtIGBcjIlbUBDtNAJ7zuhxM3COskaX8N21DobhKcjFr
SYHPh7xlVE/6vhsIBdxu5+cojVLztqIl014ntDUMlNxrKjQCjHwf+8GKEcrj
itb9Ylj541W2kaR/9+BizLrEI2AMD+QhSeDlCtURfraNO/Lz+K3gTtPUSZu7
Z8qENtURkth4AujZDn6XTJKTOoeTGXWoekTVTB7vIZdP35G9ReLoLCOAJa/A
PJqGqBR1s3ud9XBbkVUYVDzIAl+1BgNq3NjBGoSu7C5y+9fYrNRq5Ju1a1aG
IYbY4DYHzraec9OImYXV5MxbDWFZ9gaR6krcw7N8tPqphqII+DJ4WNL7a0rr
/PLAW15AWeeUezhHp49IFMEW11p7kwmEdKPJvtOpX+aC+Kx8TB5qJyI0gW2k
Y8FoG5xvJtplU+woiFDZxnCLGUk/dIhA/lQR89+cp38HZA5i1Gkho8ctMZSm
EEIwn33Ju442FUBjcAadtQ7u0keuVd/qslA4na8h9FLvjhVDu+VB4PtQgx9P
Qk1JD/6DWfkHePQyu9YuvubL1gBiecL/MdwqG5hR2zlqWYQg+QbVRa4s6NQx
6YkLUWHjq5GNTeuVD6WyGZobV2Ke1CSt97RyPNEnww8g0BTIq0FaOIySFbuQ
eqAStta8F8oDD9PVV8+oxwyBP59d39Sm0UaCo8H4TYOYyY0Ix1HJTTvDneOU
JSF66VQDFCvs3Jbd8nNLR3c3Yn79uYgsbMmpSFbTlizWPRB3vQf+2tFfsYQC
5nA861hSCla2a1I1ckA8FCREUiuLvL96e7Tdk7yJIMIIkhsUe72GoMpNam0J
Xa3QHAjmLwT0EUQuTCcxDLlLNP/Lxq4yS389H1nKR/u4D2dypagHAy3JTqk2
TAnrNF5jtOUO2KpjmUv/eT7HEE0Mh2KPEAzAOV1vdoIRFKlix4zBkLDaWjBK
HQzeZEnA6/OtIyZ4hq5mzsY7boTzF6loUr+q+utVTepn5TiUEUmF8l1mXSKU
LVOyKpcWnKGK/5Y3DOek258FgWmWX0PAZx7j+fq2f6dx/qc5SFnWXpm+DNv1
J5tBTikGQkq2UYNrPdGYYJE5gw+JIPpUJUR9RRG2M2yZMuvFQhnlZc8vXyTb
lHF2a994F4AJcRiU0YvwnzDAMLq9pR13BkVNxXhJmcMUyt39GFUscdmzLouc
SSvpSEVf6dZ6lbR4qnLXVjeHXAISBwySrQO/kZkdOm0zdk0NswvvsdCltslt
6TH7s4AspZKuUZn1j0AjiYMVYxzkiOsG07yrzQys7p0J30S8Y09ZBDJum63k
VWhn2eQAKxdqLsWLrcKUAAxP/KUIsh5YlI4Oh1l8f8DivZi4nnbzV80UkW5o
cClL96HMqTXRGEXlX1NUx4bkLj8HU7h28xcwy2KDUw0id76fvfHcpEghU9Nj
5Q4KRfx+aWRGsa5eKlpNJZ7TA3jvCpc5mzIaR07PGFqg7yvBGzLBM5lEVRIq
jj8G8wXy2PiB22GnjBhkqxzUP6rSpWd4qX4eeKzgNKDq4hjXkUpbLx9MqMKG
KDRqQcYtDj/xfIFeiWWSltsAEh7ql7D07piLElgf8nIjJlMxpn0XyVfWoX3+
fTyj+Nq50xX6d8PtgTHXmd/3ULpMpYLP2MQJROluf3bNTSutjWLKn+kWAfs6
y38MGL8npmmHVztVo2l3MvFggOcsjcUq82MxF87QFTbKIx/f//0bC57qz/+K
NS11ddoUxMzaAwhZO1hn4k/sXlQEz+FPxSoMAt8zpTfJCeNqihN7Crkmx0BX
+cAHa7/LVC1eROUbmGs28lUc12s1Sg7nUTaqCnCkzcp8eY6sg0WFloltiGVC
xDiVChUOPLXBtFSDbXBp9D2A3sxiVt2xzJ+aikceIHSNy9Uocee4BVt4/iIE
LPK+PGRE8VIAZR9z81YRwEZACu/30fHIxqPhpC6OfqiWslDUw43mhNhcFsMp
2vepT9gPpEWr5rZPv0l6zzbFpKIN9ANQw8K2dQlULUj4Dz/tJZmGdXnTYS2a
L5rrmuj52G6VESTw71H76rjWcYFk/Qh9Ce5gE7ILsMmVbrdN1zH/gK8a3HN7
f4tYtWyOXK5PqLTYFNu1P80CnWpbq9S0nyH3fL1X5juwgo7VIlg/V0GbtdNr
DntZxXwHS8ZS74HjPZH9kF95H7mcxAhX8olQpUCTku7+5ZxpMb7rqTfmqxWF
psMBDLuvTGU3LnTRB6H3O49SpvLshZKWtEK1HDVJ1wAgizyo9IAPBS34jEp9
Yf4PGpKC4KW7fDx68wTkaUudpd8U3s1ePKxD/BAO8Y33xOJI6HuIMTIjhb2Z
U37F8GLeGmEgTvaMIqR7CuBZPvHr6ClEYhYY7VWmg3IWBwRtdoVV1kHfU/UY
eKNe1H5YZRgJoajZ1IEaWAEYR/227z5YXFjoon+toMvIzrxOHad2ogcjvEOy
QhHb5Pl2vVj7l5xrzosR/bsxBWqczjierKMyttMZ5Pgo0UfUvOEpy7ktITrH
8tRJxJut6R/YDwLoq61DuhAEquOW661tCamQiq8SKsTfNPzdoAbWw24o4KRr
fq9w0pmq3PKv9CR7iarYELEno1LcNMi/OfWiv1cSgPHuIWlaQMAh81UmGFn0
FJ5a91FBhY4ve0YIQAflpNTekmRlHpI8VUq2AF1D6YNZ+ZKXltZq7VYXeaTe
ogUROvMPyaYUBhrduV2LkDzxcTQdmgF0AsiKBK6RbW0fbQzeDBxe3EDOcmXr
3ECts9wUq4EUI+zW9JVAlTWO5DYmrp8X5Wk6PPQXmId8Bqe7GLkQahjI/paO
uwFrI4xhnkxUrWoKJPZ9q0Z4z5sEIM+Ep7Ev2V7KDJlBjWVCJ5yzqEdSDEzf
YLjIa3KdNZ9DG7+bWhsOcn/He7ij4wTNVMw2jPyyi1va1vclCFvE6tOiGn+J
0AUzbEMh02aC0Vj029co/YBTSD6h/EGbothutLQ8k6ohSwvQtDmQblWg8hRq
t+OsFhSUReqyrs80jWgrRM0BYM1sY781fPJeX3OQiaIc6VL4x0n8JLzMxC4q
elyYE+QBvdmANNsVskYaflSnfkbLi0TUDIDQQB/D/Xk3hM8Rqi+4qvxg/YfE
7E5KLESRqNXtDUr4ovfgg7WZmepdGQkpjPGeCpweoilqaXA3MmPSMX0QfAcy
h0uA6QIvXsducUloIci01wTgYL4V4ObC9lSBXE4Bd7UMtwf2aJopPksulewi
8A90CNXcvzCBmja0jWs932U3VcFOBxXK3SUgl0JY0jDoK/U6uSLOb25RMVas
jAXDJhUCjoE/iTOjFulE/FpkYI7f7JvAzSu06C0t3+my8diB0rBaDhYui4uc
zPK9E73CsQQcw0QZ8C6dYjhzcoEw3VUoLlgxk+w1iUjTYwg1N8K86ECYMAwS
cDpaC4BV0y/qGcYJv4y5c0ylZLDbNsdZKAGz3V0rTaOOMCmc2n29gxOti7Ud
4OUcfp1QeYZ/7cqBySeaq7TCrG3dg5IbF9yNwuvFcZJc/i57jZKnE9KK94p/
jxrev5t57bgZ/3LNAnyhp8ufbRG2UQPQhiGW5JBGOwvASit5T/jzg0fKAWx4
Jc2L8r3Q4bDs1O9BeZEsjon57bETUGgZNnyEwIVYp3TdBVdiq9JqQUrHQt3h
WDSuje2nkGxXHglHB9aGKKbXndH60LRmLnu9TKamzuO1R0Jf7JicpJozV4Vt
ujPAb3eJZcgbiEudXVq2gTvomKqXjGqowhhfJIiFSauiI0t0kcOGfF1++JlB
A0QIZCly5eDTV1xB9V/6XAG0ear72z+KJQx2HCMbyw11lbfd2JzNZz5aouBh
cQphPHRgKYbKIIcRI++IYU0mWh6XlRNjPEnPQz4VVS2kb1twnjP71beG1OIw
Dpv7rbRXHffDah82q38Hl4/YSK8kC2TpNcGfmmDHF/DYqCX44khJgHyHkK2B
jRnR4jBf0rP9bEvpuutLvdEXmLwA4NolW8gs14JKWGG9wuxNrJGKAYuqZdcJ
xqu5hSndHy98M4x6ZQS+Cm5AeHwO2OjtVp42NmXHHsgsc6BYrMhcJYcDKXqP
abqYE1g4DCABnFbaf/dQ81pYSLKMqalkKnPcD83iIOl6rM4pu0lSt6Mo3ofy
F9z8pF7yGWxsmk+7ooPSMOlK7fo/d82hPXEdNNoGL9pI6Ek6DNgs2AEHAZyB
CdYEC3FMEM1/nKwHbFas2M9z0ybvW69BEb7tlKq43GA11CM+TZzef4VzWz/6
YjHqMOHDHt18Nlt1DMzb7AjRrVFVvBahtkcDAP45nd6cJdHSMYA+XyNElIl0
YJEbITjns5BEgxJtMqqa+zQ8PsfYBEq4SRoQ4FnhXYf9KIJ0PRIEaSmSs3L1
X46+vB+dGELrmCSg1n81dzo2kFhv6MhhRr5WnzoiTNP+SjA12u0ncnB9L4bg
XTBTNIULE8x+SWRxl4Y0N+nH6ymgP+0LBIBNiot/BZpoI+eTdcT97dIPIFFf
lNQOT3uDCSaVY5UjkUzNHFol642sClknS6iJOKFHMICVTBEviqxetPOltc3t
LUwkVDvEXA5kUvff5kLiozR6e1jpGaERv2cjT+LYfsO7V3rjH2SWyhaFfTGT
hM2O1RTQSoGQIeRjB3xBm7P4NqMdyGA6S22yRXPL4UCZPa8jCYcJ9lMnLi6y
h1ZSTYJTymkOu9rQz6kws5ZynlS44WUUP8r/7y0ETuvIPRtmrvZjprbOiQDA
z746aeykmvNx9ZZ657rSWlLlIgln+HVnJAIioX2Wg+2DREw7HEzBD4Jb//mT
AXDNM5/W5K4Vt/CeJC3WBo8LQXKD6ifr/TU1Rc508A/R5vMMHgjPM1NKm3rP
Y2h35Wsx8X4m/23idKNwmWu44BIqLyyZQ/gYWoEK5Zr8XQyXDiv8MG2o5IXV
Tasfr2h5WicQkiViRPICtEsRGMbrUobccAYPOewbDa6DapFjF0Vz+N8MGvks
lmuUi4AuTgVaQ4ecLGVa5YQ5YVh37XXxTiaQuHqAyvNlBpIpy2H6aDX8Xq/M
9t/xbujSVpuge8aHtEM4J/uNwRjpQ+b9eSudsovuHg9x88E+6XUY8DHxK7h/
U8VMIR7GXcNTBaTDlAWFSJY3IITfSHrenBc5ZNgzJ9YQM9AOvPjTxXDf6UWs
M1fNadvzTAQTNT4SSHP+arbbqTtCVBYCZueE/Mdl4nFvIOT78TozLJPQD/RI
y6eplw/LL1M4M+9dHTyLcNuC+ixyRyjWzNy/4LSRz75jGiegCb/TyUOxKL4C
97ZALV0GXqe0YG8Y4XXNCY6oSJMlQr+oKt5gneMQ9X7yanVy0Cfj7vcmkaO0
q+AFKz4WmXQ/BnIJtbjDwJBiMyfNtcP6FYnRQCCCAGwAqqdkBbUBVRNyLot8
s6Ka5eTwavqPSNlLesXAB/If9Dx6oxvPCKefpIDFhJpPd/RKVb+AiFUUVaCI
3Czg1jWZpDq0Z1EQKB6izNhDpJvVgIeoKsrI/1g3yQa2N/dulW8wMDFF9IFZ
fiWyH8y7J/a7Ogn0bD0PZva/zAj26JfuzZJU/NQYpbwl91Elipr2N0y6oGrw
RWo0luMn3SIhJFqTVbVZo8D1WzL6oevpkrKQOwVmxO1ek0fZoPqU+DWSL1Du
o2/0qjKhbm4ci9w+SBseHsZ4UPbdroxad2P7dTZdQxpFpAp8C3Ib9NBzs+MW
kJEHdqfXq8k4Mj6vPTnrFH4Wcnz3Gh1T2kJSKeeX+BTmla4UwfM1t/RhBzII
qhuaOKTSdd6aAZPxmuzlsQSNOIjOVVVlaAhdLh4ljWRqFMYPyF1NtP9J+mcC
f8e/ulRQymU/7wV6ioNwvnGSjGgyu4B2MJM9lJopKEGyoaK3b/UksdCQ0p79
x3kIl0qfpYxfGTYqFVCf4zT8Unm0otNU4PRN/JXkuSnh0X//mlji/esBgwsU
24tHEBnrpLHP3gWxbANCySL280JARhEkHaeB7ZBCssSk8i9dY4mVfkK6IE7X
N7FkhAAVxtDqaLItQdhHUDnpW2F53NHezU5nuAzR3lZrjYhl2um3kYaWTcNy
g5i+iuHevdpYG87FVUM58yo6LH9f1hMnqneZNwjrixjRQrwqJeeTcbD9jZ5H
Rru2MHNFRAeXfpbLBrE6765443wA1ksK27R/c3nil6zySmM+8WZtjlCqimpw
WvWernGmgNkSe8jwISUGVQm8wwIwWZWRE47gWiwNtx1KQvTABF5TZoIfbC/t
KaqcK4wuFEBH7HOscTY9MCV8wznvF3C25j/f/5YbVrGYJk1efM/mPO9lHDEg
D1v5ZKQU9AZzHAw9M+FPTsELngN9vT6SfotLT9yfYFFnpJDY5c88MXb/9LeQ
e78+VH9mxe/DYawlUWAMAVSayALH8YAlHLboFbo21bPInKecijZvGOM94sBI
Nj+pqr+whGRKxgshdHkd0tatByPQD6vocnUpMA2f4L8bqWvc1AU4/86ob7Hs
SVp+Ue+gxq4cRK3b6xS2stRMONT+ckDuZPkSlyzoRNa3B9mDz/dbOhLn4Sj9
HdrRuJNIFrSuUrEx2OupLydlTTJ+tU/d9YRz1bRM9q4h9qLhVgOtCGFlV05F
96YYkDXwIYZjHKIlUxRi3OY4/dyV75/D08cMY69H8RSIWdrPIrsIWhBiFxdZ
goya/g1w23R4Oy9H7sIaDbwRGqfcyinsQMNAEvTJ2Ke+ZscmFLY3a28g4ogm
hO7UeUdLBdcj9EN4d3956UbGGcKMt65dZFVSrvEv2p427KTV7Fm3JT0BQNLv
H9uOMb05HpqkMZrD1V19kZDOhSU6oILbFv40JrzgLo8YAPw0sMJCkqiDQzw4
Pp6AIwO1U/R97LEQe7eEMX++XiDDymRwHwYCiG4e2zxwhSkbBJKtyKiaMESx
skA0MkhJz7iG7P+JAR4WIY0jh40dFCrzupsCdurMRIMuuAnHBoCysv6AXh9F
KsfeYR1YMP6jAHRgZDViUTscnEGQxyOBkpbuhGbO3jG6Sl/za6iJlLk33lps
FDMyWazgU/V3WIK8n5bbURwaEvxT6FIn7G8oe8DrGa5JnmDkgqUWMamq19TV
q9Ll+NzmHZuvPCx2Dh01NV04CKtB9nZl+kH6343O33DSHxeUBFgKjeaX+YNP
aewMzXVpzSnosK6y1SpD/SyMEI4I870lLgeWuDcRh+SZYnj2s1W10PUKanw5
ZKg/rAPZIJmSySGFgpSk7YYIXi0Cp/rSAWYulIAU6wrBZTx83dQGcJJo7QjU
m2yL0bs7QdznF6taCHgMCOVoDUZaMZ6lwhHwHe9oXngabNyF6RGYmreCIns1
DduxtONi+Yo2c/83Mb84o/v63n5kiSphvTdKP9/qTvIsERBYh4Ca9UIZMLkZ
ErdOU2YYPAwl47WtMAYFoO/ijBc2/XApYC2OfhEGfu0fG2XoYSgH3UIAk8Ec
1eWZIf00YEyriol1M/HhAsu5prtX/7WTdnGY/XppwKxIMeXwCLUfW1lvOEi6
1gonsMWscfYilDBPDy/3iQVnCATof3QdRLZqP3JNGe6WBGQC7vyxKWNQB6gc
fXX8tpFbZ5E3qiN8Ls6rrv/qF9D5NHWa2Pr2PqtiRIbwt9T9MduvzGfwdzQ2
ja9v6+7bf+YU9qrtkbZK61+eo19N1cll4cguQ2C+A9San1xbCI0qffGsW1gv
lz89PdERkTAuabUT+B5JfwsWoV+TcHB3eo5LrmqsaiwKF1RGzb4XrbvKBYnW
w/i1F+BW1dzoJxoePfrHVRVyadB8ZyHDQ36kd0E9+4jRoi4okzP9aYn10xF+
IXxv8TnBqjLU8b/nR/OKNX3qq0flGKMoBNPw9wyqfnNZ1MY8ivH8CBzMZJ5P
fV8c120MMTG380X9pz6G2qat8GYp8Bg0oL3IEhXgm6/LBEoXs0ZP6CG2vPvG
5d5S2oqoEUFgg3u0sYnu8+h5wEEa3LbQrlcuvdS77T/1A0zn98lWwe45l1d3
O78Y4IDWLxnYNM26AwTtrliX05FFtIJ/SvqxNOWCkQYH68KLLo31mgka9Qwc
TSxfcRMAqA3Oof/jIFIpPoKQ8ObicOHOvsj90uNpD+IILTtqpCEWSwik8Tdo
bSgtz5H88kfiWsxVw/fPxYJuKqiHMWh8mXcvbqKVisAepyGGTrY393Mhqhjg
+FLtQMdVyrJXwQrMzZfdtjJKXa026rxCemaZUOELBD8CildVjKKkZHJZu2GA
JhmQCo29kFnjYzNP37JLwiQU65/CFs0e5FD/VYSf4vmwE3iver18DEEMqGEx
xzuxxOhxb7Kw1EwWDHZ4OXpl36YKWH9CwgeDHjlU3pCu69cqM0GVmc6nh3hv
lc5KDmEkhijrfmFCEkClZ6vYD6PhsAvuLUa5JzsMdXmMd1AieKdD5opvLH3L
gUzqhuSy9NHIrz1IIDf4GwXw/bvNSOco4jVdOoa+ZP+mmRjfjnKo1B80WZRV
wt6x82/Yti3ZC6CcsiordbpfaV9jii+pjB8SY5hVtP80DcfnThHA6tvZHHVM
zuRSHChXMPpEP4n6hQyqrxwYe0H3OE3GuWgR7aPnEKv44I48pSvpwCwnNj2V
lKTjvzhnwIJZvklTGPFpIyR3eNpREn8F+eAi86y+7alBpumE6OMuClVwPrzJ
gwvBv/DYO57oUHBvBlzT7h5mOaHDWm9H750xnXABi7kaOIrLEvX9SzbjX+MS
iAAwyWBQZYFxFHoPhLOR2S/6JiL14GwT534719REJFNfhFJokdd/uusLViiG
vGnyAb/Mn6kBNLb9GJjoSmVAFPjlPuhw3mCW5kLw1B8JLb38jzU20lo9QJkF
+K1qFnFCE8tuKj4Fkc4WjKyHFmxCIFRxpqXdzcbfcgbRak2ArEv1818zdh0L
YHaCJEjr7BiP+43kEMduXvFITRIJ8SsP/vilBwg/2Fy8e07J1TfAECXtoaNp
q0bvvlpsTee3GmDm0u3aJn1ST79paG/SxzGgAmgrQ3QnZ9wFRQtVQfwrn4pg
LagLFYFXWAPm44gdgXbJEfo+CVVkbGCUFX3uaYQRDl61qFaf8rO9jWYm2paf
RAGWPcLJn7lO4PCXOHZJMn7abXDoGE7VMNc7eRbZ+XIW0wpgjXRv8pdhMWJs
hTvst/q5mLlydyHIkwqxkEBH2GQUPIsf4nEgKkh0kJLpI0Sw72UaP3UhtP9f
oeToJocur/9G8bpQEnRwAOxDqH7FegvEwwxo8T13PNI1sbmc7iAEkcyBFHUi
jHoRkVEaRcYPjQpGAzrPqEn7CeTerxomIRD+TiAksEAH3PWeiJ7jxHWDzTQ8
0SmskHmaQi7bZqm7kq6vSPo8DFU3WRIvIICT86+2nwozSmFkF1bY2oEdmpM8
Cx8Bq46yy510qV7zzZAmeqxW1tqoIRXQCoHw4i6e2crKFcnP/Kq83TQbT2be
Y6q9mIamfmGfzhHUjpcDbsJ5Yhv9kbEBb+9Wvf6bmraqK8+L3CGMw3P3Gkow
rP4lNSw2GWKjFjgFssyah/b1SoCpOxDfBqPFQucKywNJYOHGXfh7UMxYiZHH
0hnh3hsigWAD1JvhkZRM+WTC5qkLEXArgOCIPnLixnhsneZE7hNAh/XNsDem
GLZC8Pfibc2xpSEb4lplyPFLCeYu/f1LND2h29XI89hM9y1yxuldYJvMRkr5
cH5HTIap1Ewisg4RIhpK6rDs4nYPRfUEiehNHKnHeBFa3r3GnixtzU6N/geb
/CQGc8tnSYjnFJXZhuDOBsuV6zTd9OOYpFjuHO4LUJ0PAJ28gX5mFKq1bqNe
pe0odP+47R/RJ4j74RJAEWz+x/1dGrRJnZyf25+IIxdPr2sX7XWQsVgKWdZ5
xt1X7hHBbkIjJjVa9/TaucxieGf6HrMwYHSnJZYD507gkgWPN9FHDXWzxemo
7zS7cBV4JOa1iwYgEtJ5xctXmLSDNaGb/c4rlBmaCmLytdhAzgxrl79w58Zt
L4dZ1i7FwqxeyfmIrkwqWJ0lXmKpPLKVO2k2yMcfBuVi/2rA3BbUTzRWvxof
ypOOY2t0Yj6jVLQ6UNHMz/up7d+eM39LEO1dpCcw0el815cODUK2b1lIrgZG
eo+C8KVh/mGKBzYWQYj4VCuCBqEZI5SgT7XvuxH0miQ1UvKdZRkqADEbTWsa
lQmnkQFFYxc2h6Qot3OPMpdDr7OXAC4E9cJArVsnlE6ui2jhHFrw8nx2iCAw
fTzhrJ4NkCEQOWT8zjVNzMtjMY+ZMOt9+bd/OkHm62fr+m/fidBvlMgHy7uv
AoS6qNfOOExokLwPdL7ByPANKSCVtrDUwvipEvpP61ho7/MJz1u/Nfnw+Kdo
6b8y0jSxfjDild6n4NNkQjwLcXTFJIkAE92GqV7BrhuMp5BH5qrgml7OIURI
Jx1runJ4KoGk5pjNN65mIgKLyxxDyrofKhdZpwcPpqZjKU7yDEfECS1aSkUR
pidvnfo5bh8evv6r4UAIdhPT3FCw5ALWiFjeNm4pZqYISqhj+MOun3o1o+mp
5/kOqn9njZpx2g3fxr4ejm9uU/FB3WDe6f3ZZwFjx0twA/00wjEmZ7L6OEE2
dryAelpXtWutWeHkDlg+jTj/a08W/I6cI2EBxYZEO20tx5XOwwzPQP74jn/n
6et8yp0jer3PaNQv22hUzp17ZC3Sy/f9fQz6kOcSfD4t7rDrwwbdt/Pa5ysv
PO71okMdqda4dSZrjDD6f9xXiVN1gzRfpvZ1oKZTqDQcXip7oI8S+/iFDFHL
gvVoO2tNV0jxJeTb8ZucxzbQf1YeI/O5Lp/6eoGSqTQhVUq8wN/CQf3fHF9d
A/KLXRueq+ljYgYKLZecZP5MvJYtwsg3iiVT+PBuCUAYaS2aikBbDcverpHQ
sP0v7amqtuR3KmPO6npAfU1AY7NMOkQCIsFcwZs8PDtKwywNUrl7DwXvczfy
a+dZPB8+qmdwquiJTH4wEd31TGhYQOSxUkMglK/Y/z8FdO1LzEgjQ4fjXzY9
Wdfw1tby6zar8DtjKh8WFg9/yMWkrolDwxMykgnKaXUMn0Wd00CZKvsGV+2e
yOE9Ulk88vr9q3HYRiZsFgQ8U/jFH/0olibbWK92Vx7O2mREB+etT+RpZOb8
qR3ZQDqmqV0XNmaaYPqJHIfkwx1fz1GPnKuPhuMwX8MZahMATYYcE7nKbbWm
fnVMW9x+FOtM/sWfEaHY6xM8NZLE4x4tQB8gplYDM/MF9kIXeYV5H/HhdRLo
a7XgLl/Z7bQr0scwjTsSXH0hsl+MHkFBk+PXWvdcUEUJAOf9H45f879rwyI+
3gLOpvli9XPrz/tGXS+XdnRZwIZIwLgAf+QN8TR6rsi8kFA86Oa8phOvJF7B
v2wKaS7BHWlX3ceyZN25o3g5VcUMs0GTqSEtKO3UJHxx7ALKMdrDOh9sZ45r
D62tZ14yH3xMXSWGQXbtX+qVe2dP9oTyL/q7hMPmPIPWnrZjLWVUY7DxupLp
Fh/9vNBEfvAeCOXPnT44z1DnCel3qgTgY9oDp8yEVW9ztsTj4KrIsRROcEm+
VqOYe873Gw7T5o01YtfkBsYCwjo+NiUNCTSjGourPquYQ3/pmRWPmRXrhC3N
wBrIYnMYSmx1VxwJc9AtEQSl/woMFZBDFa/c5j3eJsankPt2qZjyurKRnZvT
41hdii8c3EDZkKszd8JFJyZhvqyiX+6SLgsqP4HYu2v0n1EqvUIAJR06pQNa
iqxUPY8ICCuCb2Uj5V88m/sltr/wp8Lan5D9/zQnhIk5oFqEjoKLy/tLeojz
1zBiGNGa7JD7DLggDnGa0T8aMhJ2we7QaZd1nYUouVOQOIW8c3U6HzPGX1G1
2mBGnVdkfR1lNrus+o/8wqZ/NL9tFMvqXG0XOVgV+zyBajiNs2Vcp+odkDiU
4GH/RkZOSiYG5R1R9j3zJ0FtUYxe4NrMUoCZsxOkD8H2utycqNWSg+OuREC9
NJxyE4J8OKfaqbtiMncaQZfQLSiuwTAsGiWEMzA1dqE3STEBU2QBgqSJUwmV
g+jx6nBsN42lHPdEa960kH692vfV1CjAYd/ckMaAaUaQjFm9+w1JJ2M+H6Zs
frQnar+S7jBXF/Fo4zoaW++KnKfoBrgqa98MvTXXxSnrwJRP5yMjy2LfZkvf
HnNWZptDfowkpgxdHlnDl9DcfJv4c4Rcgk//Ggh7sYlkIyMyag6tWHjRiKV2
+4W65h5gU+K7fhOK83gckdP7Qwi/cr06KItkfDJooO6Og+/ZPWMIEQLsQmTG
9efUpqSKAWF9jSmxRW0/ME6Et6UfvKKouBwqoxAHZA9uOgaEB9naPp+1DYa2
QcnuQQMATFqdFTFD5ALXFAHRVFokRRqfGpHYMURaZv8AiMxkr55+EESYpQg2
nxSM/kHYM+DiMBCVAkSI5xKdvxIVB3SM0sRS09tVVcDQnFP1rDoVXDRCE2RH
HAcGXrfcQoVeQ3K2+bPKxQ3BasCxuRfs0cFp6XiMQvYHsBJnCFaRiS7/KkHk
BxsaTpmbjaKJKDYVIykZZcqSPsYgpEntF4ZfxCFYNegUyWjAmwEDkJycuRIN
FmwNzFMSTF2XtebKXTueIW2EeNWk5PWKVFqkHEJToRIgd+wN0Dhxo+FitdtE
DKnnSC4yD4TF49j1WMBTYh3QLxRdiByqVKWN4KJIEnHIp9r32x+66MtrbqwY
h7+4VZAORlcY/Fprlb6kjpYREcbk4E+BVbDdjFHZNZuH8QdJMkV6IhmqzrgC
tfF9D0/zxmj1rc0u8VUgyB+SIJwe49QFi4VoXia8btDc3X2jjKxL2XtZwSyo
59iLWcjs0KRzC0UZRtTo9OVwVCYzYx8VU75FCjt3gMZ2xibkLIo5by5I4bK3
rYAYyO8T+v867jdX1ixy8ewVedqRq8Jy77zJ6LY4DkeaU1kM3B78NJI50qAB
BHkY/H28ShbueuZq1fbaDnjhpOivurFrFCL+VMnYWnmKTzLpOWuGRGA/XuPo
57rl6hSUyQdj4OV3OnygLZ1m5ljTdhTMCAStekT1ZAQIJAvqCpA0115+6lPQ
WXNPim9qfU/4OT+oTQS8yHfb4Q43SFQX0m2vhnB1mGo4tiAJKXe1Voinjc5i
e9QDFnzUeRwhmK3Wc3EaCO8drC8u4eTSkS4LWmwNRNkpo5Vsf+crclSNuEHn
MXN0jbrpd0jIJtPq88F5Cn/7TgA9GunHhzHkv8Uw0CbmB22jPY8+rHIQhJFN
Gr/bNecj2u/vYImTHshsBq+vTiwA+2TYnNC831pz4n8aOcfnb8OGfP9F50bM
9EUfmug92QRGqGUUbueOIlLAt2rR5eFywCm65Qp9ZKZGAu34PUGToRs7wusK
rauf9z4Pqxv5BzgAv/aUZenKKwYyQQGj3A+hEEOHlrArkfENOo5taf83W0Yl
aUcSIW2eIJvKd2DD3KdOVAxr3jj61LxMDwUnUY/wCyQoTvoqcrRNTOWqDHdJ
FywHWawgRJJ6N8tQ5VDm0otEORbz2EmAYJd1A7N7SAbRazHpVHWFFQQU5WZK
9LHtsL+34HwRTJdvR9eM14SzfafRwKJOVhMziAYWaUZ6NBdW5SPwWvoJMTrU
hRm/xZJp7046xBDAOvY6Bc4OWU/8S12tQlH4LVGuQnJYj8XQ1u0aipeE4VRD
0z9Poz8SWoUpEjF5LALhcgK3MzI/RhGZP/5vWAfQ2mbgBqch+fzHpBNkHj3K
sF4oQjBaT/jCNz3Om6/hUtcouc7XPFN8agDlP8FQU6HwD1suzgzeB7Y/11Zm
+KjKNkLkQHZuqlyoBZQjcftYq+q9i8dl69D3BjBwooifJleke1tDA17hclJh
OtfxJDCGa/SoSD2f24xjdJ6UfVE2RMzlc6Y2KG4iIssu6Suzm4uvJMLdDDr5
1PVxyb/O/hBE6KmMYCWJAjtlXpZKKaXfOhHC6Q8//ndk4+O+XoOvIswBQEYz
vorzPfsR1xTbsgelfIjNjYnLK08gWXsp8Y4IS9n0BYrKDUGhgvmKCWSbt7nB
i3s5zuiF5kazBys9w0t8mEKOKusBKL8Qg6lf+m15lEY4ktgdUsMePSqBto/0
OEkjbHtEWuLPAOepFvejz0fTvWYmW2pz6pUWTF/VIVo9ht4z9jjZVGjUrnDB
XFs4zoTGhoyhwjynhSdc5nikroBWX0Y/PPPiqtdispJZvNDl4UbE0pIYV8kW
UyvrLKn8ZglHA2CrFeNVOstC2hdMMsR3Hl7XLuJYNtkcWk+YQ5hY9Q8f6sKR
uUG1K7ugRjQOnugg0ds1xGU0j48tqjnqM2DE20gzfMKEeZn3U5M7Yf5fcNm1
rtqjabLWRk/8SDQnL99gG3dCyoxQZyS4Bm6UrugTweut3kAp6rK53J1BKFR9
+m7FmuwcBTCPx3G9FX0LVkU4/Vu2+WPRCSkogIkrl2AmNs3EABghTuYim194
sH1+g6A95aqlpCCoYx75lcY/1I994Zjp/r7JqN22wNJ4g9NfSldfiCCwXpU+
RbWd3X7loH80cnBvT6NYjOeAbVSQReaNhb+7mYYfb2RbNJr76u3UQM+/QRmz
syIfha/XEFBVeZIrkG8Vtr1xE/D4j4BI2HS0KYAxLR/Da97AMy8jl9iVvJCJ
CD/N7Gf0EtbB8SosyStn7rong6klljfdo0qjt6UOKLMbIuVRnzXRJhUxoy9S
GdrqqQNpQtMHcp7gu0SVHZrByHcAQiiGErQCCppoY4wUyxg0o01bCkp5hKfg
zbpBC2Mcz0QxABJJpt7/DimtiHsUoZPCZF/pqevE27bYM1azrUuWqcUNySbC
dbxdjv0zqze0ytBtrargpYNX3UocwbICjYMRtr0DxYObbZLQcAcDrlPy9qxb
ATXUQSdC/cNLZikecpv4fwC/KUTbNttmS/T9vFEb+WCxjrT2AwQ7Turfx5A1
9nHmDJZWajQhvHSLV13LA9qP8l2CgIbjkuXKmp4hPiYMHSl081EVyQlbeF/J
5nbHC6nj8pBjM1u1cvRcbcO08wGAE8dg56TGQk11nv4B/pBZ3yQ2Qn8OVDRV
s0JignwdOXwdIdJq8sTgWuEbjtNSPUXW08pgK3sU27/1LJMEEj/OtNQk4TfA
nKH+4dY7C8qCFYYzTVbDVwQarnApNYSv7Tbfa5pFoDceQWUoUzoglS0tP5N9
wTQK58mC/a9Cs1abJFetoWAuewYyJUiOTlL0ZWHkvk8+E6XO60D8ODLE2Buv
a3mj7a512qAeRW66RVND60sMVQD8+F/ycdE6IOnPmUO9YQ4WqOTXCnYoRBZp
AwX1jE3RLxsby6Q8cbvWNYRBf7A7HS/5TXsCuDTeVhZzuyQOBdeTtjObWZk4
etLMuGE9feQptfSJSUoouB9zZkOofAa2LxHB58twDJbjvgOh6SnydkAdt4UY
2y/KmZCGlf3i9FUysYgBw9HZXnZEQ12cbt27OpCZFjD9XMi7Iik4SaM3knp9
YEQIqPgSNGtzn6CNXDKyRuctfbOAfALuA1TnCnFAeakjAac1KlbmvuHX8WMa
ppMvL3xckczq3fDaC2wuQplbE6jfJICO+3AX+FW1mgrz5MhFjCWbBFDfa/m0
8llrW86TR9V0R9VHVuX07YDO1sS0Cin4ioN2KwsIgO4SGen3fKopvqpPLjqk
Lapw732HqJ17vnOCY4f6FQkBy4kzA2YsTCTK/4WIQygCxQf9NKRq9yXx58WX
068FXyYnZuibCSbIYBAvRjQGiotPHpNpklgMKuSqpZH9mrxHCm5/plmb22K0
kiSibQsw3F0klH/6Bjkx5fqK8SwUf1UHl9yMLXgZbjG47ewQsX/fo2krLMa5
eXnfTO7C8L4Z3bjd0X56f1Dn7YadsusaCj6VrwAnkC4g7GB6nWZYRpV9GrWO
1eZ829IQBGc6kreZBqXHq1NS2+b4Sz9crHdImy9/x+eDv5S7WhtLdfoKLjaq
cQEpYPyhIIOtJ7XeP8i/lyToKvJ6ynUqEQOPoiesoPQ5r6kU6Mlt9iWuVVwT
Hxr6azClT8rq6EKEBX1y34x3stWfLfO5k3ObdRZDOcxOQmgRzDdpkruoC7bG
z1wtjIY4ccMBpJM7FrwtYNVq4JhgcR4wKJJS2u18q+Vtya0v2lgz07gpETTE
uR6Q+OCiHZOO5yGB4wYDQOimdseKbPRgA0UfL8liZIm31BouWYk55GvEB4b6
v4s2K8nXG6fnAC0336EATEs97TSIQC1JjfCwFIgab60JP72U5Kz+AKupdfq9
CbbDHCTt6dhSsm0KOtZASqXmX4XbLRinHMt9D3FHy5uKuQ1HD9Ab6M4HDfoz
MZdE+/FeEtsiI1qC365kNkLVFuyHq1YTlDDYUj+O40BjCxSomIbAWp8dtiaZ
HgJ8am6IaBDWO/C1IHtbHulLfAFyrwv8LblYgbEoe872RucyAVqhMHPkAGom
4807Gz3esuFxepW3rxrXiCfMhe83LiQKxV5nl2krDuJwXeKaYXKWrk0sLrKe
8/NjVgpsimcSYe4hPHuN91XtWqUUk6Y43n/RzfbwnkIKuAAiUheN0AHb89j8
OtEcq6rWkXJwf/CmG9zZofukw4xUuAvzyZe8aDD2Bs2obYMtzwKGwsanspak
jA00u9bpEM1FDt08nuIffwQxN5mhFwTaR27eJEuicG7AQQUXvhz2fBNuiGVO
nYHuxE3ZMV6rK9nIpqp0HxZ4VPB/U+7e1cj+wztEpWji1BZ/WvnOssRogFGI
OLoZKtrk5hpj8GCgBfopgBJYoQj2lRqCEBewmYrBi6VAYfeuaYm/Robi2JUC
zihdaTPWaeoffaUAW29h4RYpbYH8AJvNFZjcw7c6SgjZ36qBOq1ESgmai0NU
EukST+ZvqBQ9jU4ZJfji28kaA7Q+GTYvd1DC3DV/N4OCWgGkJ39rhz+dioQA
OXcGnOUGajz8qc3QHzWYV8kvtO+ytXakgzss/0EUkpjN4zxRRskwpGsiSm/y
Zj9cB85OkRUrAzASoVybanPs6Yo7Hf5I+etTx3v4nkSHi/Ana0Pi7bg4PH4Q
0mPD1dCcXiBbxLyItLcu3Cxl4iW+36fSftxtn5c7HSF9o+TFaDH0qn0sv5w2
+SskQjlO8fVhP1X9+B97TP1UA4yVjFz6REpaEjJerYyOpN/TrH1LfCy3+rQQ
k4F0c59I6N0vaB0s23KQlDcP1qWyKiDqYdqY0/kfate6c+aFs/Yh4pCJJIIP
PrYJnA7qM2mMU4uWXSF3x2Uyu5t6rwE/+lvLmZHI+UVgaQRVEHEi54Fabm8U
kTd86WDordOxme9grTuUCxGgp/TyQMnn00OhvolwH+ODf7PT/2mcnnbi87Mq
EWAWilIiX4STXlYpYtuU59g+2y7UXdNYIpyXrL2LCzZESptsisW3xrPlTwex
gy/KZNuFz4M7AgP/mlBiL9hSZ3KP5RwiRq583uKpocwKwDSvYLLKCIlb9/aa
HnfKAtARA/gvaez1PdFbX99axfD+9nQRXqAo9sxICfVMfYLXEzPGSzlra98p
KQ7zAqEFJmH3nm1+7lFwzSm6KUNMN39p7wPdfjXoF0tszeKIU1XWnyr4on5R
zslO2mQOv7ijYF9v+bfPyv15h/Hq3pvoELrXB6dfD2wam1cgJDsp0cXayc6q
M2VTyd8lSelt1KiuHBHYi2n3yovN7yqK9jRPalFGQAlIaLvy8fpLaGKTKBkA
C547gNrsoQ+ri5d5PAwYnr2dNXoWaewdZxSUkhj9JppmCKZnkXKFzlAEVUN/
KODHv+MI471dzL3ikGs7pXwe2Md7rtM02TP4s/x5dVQAtsiLfL13P8K8lQjK
Wkjp60WS0pYg8HmikdxFK2gdV41uMG29/mOkO8fhQjun0I2+fM0N2LgfKvUa
olcyFfJXJc3Tyf1rrD8iBKOIvpy5b/LjfjL+pTD7hcoXdDKKyT53upbMMZ95
TGslaqijLUWZzKKkKfid9h4iEWKlXmKHuxJ0bVJzLJRDfUTb5W5GkmXyfM3L
5u5gigTTwQk0iJzi6GNVGcSvIn0No5ixMHcIQH8G6cplJoB77T81m0vkzxyG
9mtl4J+WO+C2q4hHflyD7v9Po1rbPQFrGKGd9h6TxFJT7C5RlJjOqwkZYw4P
oD651bJBtqzIRJU7adlXAA2ujW3XZFZ9HkVOlVnS9Wc/Tyb4+cZcQhlInDe/
OHF/gjquRHaIvhxh2D3oZ6xTMNPhK/787lUA2kb2Xmwa+utxmtEV4z/yucFP
Ix1JR1L9nZs5bl4AifdfdS9YShi/+lEnXqr8pBJgleDpqQeFxI7/EDU9IXKj
lS9MS8hvd1vCp82QrwHSUuqIDgHVCcFGRx1QKWuy3qO+zjj4vcGXereYxP10
7w6d7ayRnUBKkcC1JoOiVV9jcxZdMOP9ZKz/i8A5FFEIU4/CUnJj+JpWxX2w
zXdE5rN9WGQqFmiUmvIe71s/+Gf1VL6jrYZj2ZDDDV3twPAIg2aFIaRUDPXw
ef0pCnd+/oq3uzj4kHhwAt7uNYiZDA45wfGPEla8p1bVyvYbcN7acjf9C0EP
1rsPtjaJAieCfzlbAEGc2tQOPswABZmTtiVAzmIxSHTqRPTXJQDjn0NeBUoH
Y3nIK14npdorKiTOLtgl+TLJIT/qnifE5tUP4vHF5kjsyZBhN79HVJlnCZZP
Qpog5BahFluiUE/lc0TBAooZMxoVfLW7wHb3XKkbAgC4KDqIw125C0oqvUlW
0sCFGyD2O2h14WSDowrw9ycoaTIO8HfJ0+OSwLh/m+Jrg/+UR6fNs7sK/WOj
NK4atp6M0YqVNdaA2T0VfnqllDUG+92VtgZyLjUYuleQP5kiI9CQuHGAxtqE
V9axcdqkZuumBov1HM1i3bo4adOrRseUIN02YktY7B5dWnqncgLh5vWPfFWV
8u1diKTT7V+l60HI2o5/mmv6SC5KFQSJNu6UnuoVl+9yULxRFKbOz+1K1ZsM
ft0UE6Av1HO8flnZ2cpV3qUNYurPRPbD0BsqGaCyxCTxiQke2o4tgB3U4SEX
23mmsWjzyhpAYJi3SB2o2780o2VraBd2/Z5y2nLfk5ChACN9+VGzILx1WZ27
7o9lqNRQaJTpBXE67A5/cTVRilUBHaJM4oX4+PeKSR9vOhnUvVqX/hz0Jq5s
QWMDpW6sGPTBhRSVgO2onKIOXzOaL8clUvMmOTZosbyLmuznGsXzW9FKveAc
HAh741X2soMntilCYa3mpNXGev+q7OxLJrsDXNxd1hqiVT01GX8zKYBgYWrK
POj8m0uLa2BBSjW5JzA0J8VqJZkTg6/yuNubyl5gVeZlzkwdrzzeE91l0qNi
oMIgU+VJIe7nZdDwVpS0OOBmKCjb+nrifv2lFOhbbViimt/NgkDHCWtmoq+q
0WdiLlEU+zJdQIsot5OdUpfGTq7ppGIACa/EIJMec9STvcUD9k+ck+BNehGZ
fKJdNJymIWFfTSulb6+RBndJDN3pSpIhILGIArxVJa9VGgG1xlmB6cKiSeTf
mh0xgh+ay68jWzKPoWX/E52AUiuaeFgHGMjAF9uuRWOO0I79EI9VWsRFpthI
dEQQibrwilPIYBxJb0XxV23RcbmHsv96gjFT6OeOBGN7ED+s0mBsoTxCQfAc
+se75yaKzWOpVX8PG78Or4FaFyWuvo6o5Mdgpzy1cvWQdSpRYOTi6WUKTENW
AlTR52hUtg7YMOBeTC8/QOC+3tPZhaEhvey8qXsLjF5QLkqQ+wHo1axF0YN2
tNmZaJpLxqQboWiNu6aMWRzpYl2E+J8yoMnBeXjkdtyqedI1hMUJ7b6QHsL9
5ULVtMfibo1jexy3fZR0/zzNCvCwzrt1W5Szxz6YrxFyc5jqzIu5LKP6D1Dg
CiNbqUSuuy1JxiR4xkpWNX7A8+gsBljO3UTA68HDgVQcA4+UOGUVc8P9YowZ
8s6WMjQv9Q2tZl0fRPI4QqZb82Ft4qbWFOmOaQxHC6G9JPr8yIvhAxBxhuIQ
SwRyPZDb9UFi55Ww4qv/flWImMIX8dd1MJVd5o35JhVFgY3qm4cSOh/8LnwB
CnbWVxIWvlTY9JZI+xdi0KQ6Mg7ZY18jGL7zFSS9EA2CTFW3Eh2qFNCkPa8a
UbntCnonGFNX2q2QhxFQ5k7IQmkED83VC3WXb8KCCm91I5lUzGhvoxZ8asWe
oAa6sS+AwPIdsNvT/7SNmZ64blgQ/5QPfEIvaKG1Y89sJci7C/CTgyArR6KF
kNXlt9zIlac84FEyI25R6qyxW6lDGrdjeDawlgpbsWmhAEVTo3n7f5bdlx7c
m6kkZDh/N1IcgZcvd5LxkVVSZI3kX9wiF2bWVtcsyFTll2SCCUEjhX7nlpvD
f7H9nuUDnYEmJSkLCaN1pZgIoh7f4aT02ctCeCqM2YpE37NyGP7MAu4uLWcL
dGw+277AU6LtnLTM2O5vEtbX1K/BL7Xt9rX23hk1lENXdSsjCQFyGai3vfgq
KYoS/3ZcbDfQy6nxKSKwt7VJLqD4/DxNGgLKv0Jf0L04Vd05oSSWqA1jnLxK
u0+6hRXzw7052cwez1brXdTPvLRqDtJbPJhThhHg+4RqK9B33GtjGADStdX4
kF1yO7Dl73iNxwuOcFygys6PApzW7KemaRYasmaMRJp1B0+X7xUSe4zEHNIS
+g2bR4mO0ddGFA6PhZPQ3GSoTepeZnneQGGSXHtQBEMplTneBdOrp6c2mxXs
kRjpvrtrvGDlhVH5JCSR+MRj02kQ2BRwTpEJ4FUAf8wtq5cEPs9A+V+qnacL
5rhg7ryupDPLGdr0QWLwkNbSunn/yzWTKsuj/Kzj5UehJhC7wCXM9cHe4LQD
yPaO3UPCCGapyCiB4YyGpMmUjm77yWILhn3wdOTzih97xK56wgsOffd3ZPwU
kZE+RIdclE0vYBFrby1HMl16PVnzb6AwAH3RpI8IrvqDpQIF1ohg2yulvDmv
c7btm/v1CZj3T+K2TNKYY2gAfZuEEhPMMYsft6zc0johVTJxyzfl3BbsgPBQ
tkt4gEqP+kDtZ6FSnnFXL3UF8q1Qy0mwybTtO0VCqAtr9Rn0h+C6ZYKm0Hb1
Rs5objxuGTTwow4cF/Q4hw2PFk4V6w3VU6CGHotYWFooSa34aJvbZhwFiXNA
WLCETwEsOdfrtLwma+s6BXPGjPDCoypsemi+36vJwFB+0ZdsCBKxw7fWGogL
vfyg2MSkJQJnNEeXrb9phubNR8TrT81jIsgc+Tia2E/xmMmZnlQYm8mpGvFm
q2guroZJNWfgtGwQskq66Al8oUp3inLzFFMeXc3kwUflfoWwCArDsr01CVo8
xaBT+dK8pgvrFzuBJIZp/5w360znpp+JZvS2MxGawhN3/RAYeTF7zZgvSFTt
Y8xqD+rRwLRVh/cA9AbIbrb9hhPAXXVqNM2NAM8gvGkA2UPK0dhVeouJGZmY
2rwtu+g3l4B78Ln5mZGCV+TG5utjPaHZB9g4d7a3mgcMOxcaw9IcujoxvpUf
yol3mYCb7z7WgV0hfuj0hWFaNm/H6X9Olpx02PZlZwaWkaAt+n8PqkgItlL3
7Oawzw4pCaFa6l9zZSgK3pXCSE70f1MMtoPr/8Caj+B+CqmWaLRwgPOCoUa7
xOy1/Eh3OWWRhEky8haOd9POJszkXE605RG4qylNnYqYtsqLKT1P0EdMPI/g
Lh34bFq9dqasbP4SA9alrPpqpJIRI9qQJn8EIruOIrO3cHPAAXOpW0SqZVEt
ptif3qyEcbQPZBCc9uvTimbwDqoUrUCJE0KDkKAGEXiFPbru7QpLjJIgAWlA
DeOUBYc8C53Cxkb97PQ9lvGvzDarlkqhbJ7XdbUskNNuxRtJw4KQYF4ajQSv
8b0pcZ3bS+5SSNxRLqgih9nAVJqYwsJRY/UxdeiwZpS+DfT8OCQLQJS5fkxN
48ycXGUYh4uMYtYqmCEHE6Krb2sBJT5B3HBhdoHv0dRmHu7ftljDFqb0qZav
v2O05xK6iP5/TUMdoL+d9KwBUtIJEg3zaVI089W/EDKeEkKJjszPRY3Q1pr8
Z1NUVw4nn4UNtIAxKDre3H5ecAVRS7+a6oQ+PLWFRYMLLCXq6z31wAQ4Ag0Z
dee5Qhq+weMGVEFLhkYEvWz1rpEqFwu7vFHP1q7++ZDCMQiEv9mLsIm3g62s
GGUmRl/FQRDntVquc0JJ0Juoe6ErLZvkbVqdrtcrAfpOTFkNxNxd9QQ7gagu
O0/Mtujv4WtbbsVaF9JqUDnsyqkK242WXdU/Lki2Sog0qW5aP7bVYZjfkbGw
UYmzB8CUXYGmR0EJ06Le92y3FV954Ut759gJOUcRh6RZ9r7MYdSz9qF7sUBq
QYkk8gLOtR5dB7+rsIN4EWR5AlFrVTcUEisvncYzw83W2oIAinpmG8Hd7I8Q
XmFHA3mSHTc/dC3QCs60prZ3Di505tJbLeV6/CVz8DpsiZAa+lxS5sAcLcVI
OsCKCpMHwux0ZNPsvKMjcn8oTazdGbTp928dX8n3YnyzZre6tHee7hH/3eEs
hKpLXDs3Ve7o54FGsTa6GvSTBQwyi2H8wNuRi/spYm4hXgDYA7NwsZcWZ78r
LS89bbzQI35NXfzHmd8EZfCnjUl1QQgYged1YRu9UZidz/+8hJq+DiSM3TxN
9t6p2ivBSr1qE+0H1Jgy2yFwzVJCpwZcrMFQPLu6lKs0IKPMhA3/zLeB3fAD
Trn9XSvoETBXYwJ70Y+N87dIu06exuiuYJ3LdZeIKY4nMycnsJx2A6SC+l/E
04hvf8EpHdReIbANro+iwcMBku0Gn6U+KK1BTUrBOb3cwiWqtRGY4lqyKFr+
FoYkIbRFdFXCOUIySRtcv9FLjBSYQo4lFdqmgDPHwe74GBxulZvpgJwcWsH0
6S0pY5IL7350VSzwcDPB07hTZQHwgBiw9xwHSVfFHyLjyVqDOe5ldj83PrY/
Ig9R8aPz7M2mL69ru3p6r6NBcQe9qATGi5VP0BuLUEV+oex58A7QOkdjcf3t
thHOtovaMWzjwNxFZ+ZMGEh3IQ7xeq9YzmtWgQR5jyT/xd45kLr20v0+ZJSM
bKnkkTWq2sBNyWPjrNWfu0P4Vvxp35/FqDdLKX3YyCQvZcRwj39tao6mAghC
feG0NCzwnbpy3JJECci6VBxpEd//ws2/WbUF1kTdAh5psD5LBI4I/gaFyisv
XNNHBfL+EVDFp7lL+OMB8xaELD7wXSic9dTOIPgEbaE0FDqJ1cxAbSe/iOi5
ONoq+zftT/hqxCNnnpE+SVBOBtkcgNVIEZLyxVEgFGDl/AFsXvnzRaA6PLyx
zBk8SE62ORbMmBA9KDIOPmJ97JWp1s4rAnSJOD3J1DtW1KgtITJFvbR3ZO/w
wSLwmHLWzhpii1UzK8jS5+Zbl7K3nF1yiDT4k7A8e+XYpIlGyxnRh/Z9jfvy
8MARunLPM98GhoVywhrTJYtA7AhaHBwH5cE93LJhmakf9sa3JhbId/5305XD
3K8cFWYRBtuxZLCvHwVucq5dvvWFl1at8GarfNv8OS4Fgw7EmeDV3v4SEEc1
yJoze0/NqJywvhz3VS8SV+qHbdfIKQ+2sRz22rXhJr5OBe9+epE0wBtutnwj
hSw6lClqZy1as72tzf01CRqVrZ9NSzPiYfeRz81V4sfjZcKGt0Cw901P2QiL
ZWqZaOxvQHca22Co1Qh1IcZxan3dNTKrNI+QKcBAdeh+aQnndJa8rMwmB9t8
mY2m93b7sbFKFPbpKqMnHEXRKCjyWUd/yk3VBJKx2ja9qSFU1Z1VJfQQOA9u
oFMOAWrEU3kySoDwsQzUukpVvtdqrSRElybS9kV5p7O4TnYlJaXBgORraud/
AHVPC9KSGbe2EiEWfXusoso64pZEdFBzh6WKfCon4fDvsXHXFVMfdff0tdDN
d0WZiI1F3VdLzLk4EkusBkzpMaWFP3C4Ea7vmDPglPLopDGRYL+BC8/UobAy
w/rRnoBmyzsruUEWSAg73zBP3wN1ZFIDyBFeKOozmL2nt18z2LERQSBexmx2
5w/BxGmm+g80/iTsUKqk6e/aEUqO+2FGEXtTfIH9UfJr7mcDTDHWZDFooSOb
e5ZG/0y9O9C15/blEA7ja2R+NzFLvts1asItUdtX4mIcdAXbKpEokXDZo5v/
8WkUQ1TJOW/TMIu0YVnAEYXVJx6o/UaQhsRAbGHPO579tDvEKCvhtWvWP10D
YoV1O1LXT+nxbXg5HtYFNVwyB01XwPq6nOhNBA7ZTDjIVdmUEjMskGfLXmf4
Ye5oAQAjiMtkRKOVyiM8fGCOBr07OxduvHfZJUYApa568x2J5RC2l8aVaN/c
cw+8eQHrI9o/IJWElL5DANMPSKImccqEyhHe0JhtcEccobGviDL2D3pQfNUP
VHKRce3qKE7dm4HZwG20HRl6hf3cHlULJxskIW7dgduFM55gN37zqcn/7Inc
DBa4pcrvSdbNfc4vneSl484PiRKs76O6+iKK5r8GM5lcL4DnoSNKZeQSIgNT
bNbE7JlhYmJAvgL2Jd4q4lkbZsv2QnBPqgGaog9DSkuPHu2BoSMMKKyHOGjn
ooXj/dOWN6ISoB3b7A7ovv6xx+Sd0JCsBIDh15c+G6B/YxXL1UmmTowJBEgX
txOfToyGOmp+vPjB1bpPKbZC1A9dBIJOKd6eQaxxS7u6udfugQQFHq2lEjQj
Dc8isicPjYp0ngA8tTjNKgP/9yUDtMW2GL0oXG9/jrBNg9vaRrLgqc4uRNi0
D2tLVWcpMevOO7bZRhuH6P0A8EGp4on7PUjfvu5HChiAnIGsIjbfixivis9j
IxZhHxLpE6LFla46B58zYfG9Qba5mUqvUpvzfXu9JzLwquSYIkkCLhwawMB/
IRVJOHs6HaQguPY4BKd+xH+TEMbxXYmgnziRO9JtzxUp+qWxVnUbhoB//EHh
31rVJJdakcd72JTGYcOeBIyKx8C5TCxoeNYfhFZM+DtJVR+ZudZdAkH6RKF1
VL/ymy+EzGDURV47bzlYMEWXi4pGG+Y0+jirzsw51RXyakp0ftq8KmMg4aWa
TYq3s9FJDslTXD2uCUTn2TTPOU1GcA0xpx2uNNTwaolIhbxjSZ5BvMVsah8o
o6EvhMVDADaPVxPCkkNYf4RaEIl/rNDGKhNbSEkf/yPlF2je9Hxo0R3LC4Dn
Dw1mAVw6tjEaSIuaB09nCOG5CmnyxkndZ/HcH2gBaUNzRJrE6xRZmDIbkb6e
60Fvr6mMGFDtZgdqrA+LEkmhO1YdGqa3SsIm9IbYFafZ++Q4sGjlBIfaoMtU
Gp7LCKvw5xNTVL1t1Gj1k0LvdCcOInsbKbyLa4day/ae9u+2uKPwtnN8W5NY
kqiix8bQWJQ9OmaFmb6z8tzpfDo4qh6qeh+rWSwqzC3Fr/pRnyDnLG/FNaQc
NphJPjHk5Hun3K1+TqbjfX+lFJIKDCosxknlWjPbV1D47olhVQz/2Cq1JFSO
fohQI7TdsWzULPnNEYKaZ7T14TTB8J5RqYN3vBSZv5sc8CbK4FtM/aw2d0l6
guUdmTVXa9qroJSZSlPq5zleM+P5lCOqQ0rYZy9pZJsWCWrOkjzRU2I+RzVE
AQMYhplIjlPNEEd2MVhTs8lWgaXKfKNnSAsnrAaSZd9yRc9P0A6vk57WN9xK
0F6mn0NkY8hTIwZM4/AQMpBD7p1D1pUe+0XHwnzDBEQ9vq3mJI/QEwQtCVbp
JyTUar8Q2ZoxE9cvOpCVO0WpvJ4huPKgmClIWjKdPihKlJq8jEwIeD38pfrR
vbZm6Wu4x16PE2W+vl3MAPln2u+/8d6qOfBPuVl7umLoX2KIGRlWZL+1Z/Ct
PhrTpbONmUZA66HfvNEE2utyB32qa96t7Lb0WoNui6I9h+d56fPig8mJUdbb
+MMXpp1lTcvn7Se+Jzxah3WMHGQnHwBncr7qQS5+bExgE1nNiu6tBynbwg7c
3n3cqzo/sRvdHVdIYg/rNmSD/AkDsEno+mQE0jIVeqpsZLXkrFCuK8HH7P91
0EVaNC0oDmwSconSXNqawAQeQ7ly1YiA0ngaxhCvGX48FjNMV96zN7zp23HL
dlIfKiEsywtL63GiDz0IjxqIV9H/6CfXTygNCvfXRA4q/vpeFTID/svos/OY
o8PMFYnGnmkU9ngKcQ6hTYcDU2S3XIhs4mwSfujTdO3uEaE0qYFqarxHOmk5
IaN95MYBaFphv9uBPapmWXPJoMv47EHja4azi7sjTyjjJ7Ine+n5ickG5k84
TZiqvyPModXTHvpHuojYqXyNHWWVKVTexBO/mJK4Ct6FCeqAxRgqrVq8Fp2Y
JcwKwzNPG8M8OxI2Oxn2S38GEizS1xR1pP7tDg7/6NUD62/Fs8w0J/5kZCPR
7hwrBIMJIhak6cb+AIjnzYTUCU/kEzQb02U8jN4OqH3ZZE5RxkDlLroakuPJ
aEYQ0R6EViOsgxDAVOpUfim/PtCXK+TzPPsbcsRtZk57zves6+gAfEWn5pcT
dLdfYeGurft0bfmsBLuhcSGh1QWg502ccCfl9SO/PfhI2iw03onAL2Mtx39G
XHWPVgLd5kxM+yFNDLAoDuf7eYUvCSZGPU5YtVHlEiAgQEf+gt4BJtu5XZKI
RHVtqTl5bZDB1rNCjaN/hpb4uE3iKisPVGC1guqJDGI3Ya4DRNvGXMfAzzoL
cfX8dyEEef0unz4/US/GbdSdebPtaYKK6/wlAlAItwXOgxVLWkq4cgNADSXz
GK3PHQnDQ2NOFCrWWYwtuCtu4GUrBXNIxR26gUTopoQ8t5l1eZqD9PV9L6a8
XlpZNuezOuQ9aNzdxrxan6LHBRvpNkUK25T5LiP+YE8ggiSHq0U5Y7S9Y8Pi
EbW8nKYMtYpSa6bBlLU51XDYRuCMfthpl6lBBI5NhgPulKk88k6cIJOTIY+e
yCwvmZgVY8dh8eMKtBc6zzjcc+r4VuycGvp0mizvL/TYy0Ds6RsIM71LHxuc
ZiA5DuBojKjMVipgZbOMtyKTXN1+WXACRiE/0JvTyvMv89Ptcn/4KP20Wc0p
e8FiS0wG4D1em1dIhLoZmSN746xrxiRG4pXctZ+o2gQP7SLzGoRdl2JJPIzV
P9yKqQUo6fgIs6AvO2dR+twxszmUulxwOBJIQW9lhitOxrN9UpN5skfv7vqW
VOglFXco1JyYOLwRTw6JXYtyLUpTN6CJT0ocyfkOMGxn8LfIHYXztl7PRNIH
OYWwRUsyZy9senHBYvedDdsyjt0c4MaZg6Q+8XoBTtTJHzgxoCmu0o0oJrxT
LijePPlxatrIHbYZwmfkKsHIDtojm/K0Cr+GCSDZguZapJRbWP278hjR/4Uc
sQnjGw50wrjLOOfvBIWtRs7v9HdzYjEdplVrBFdGnmmAHqqTEHCyAcuPp25d
tCJnxjEOH5148JSYQaC38kVI8azyI7DUHs+Z5Q0N/nhWcNd5EU68/GxSGOAz
IQYfp37texgXh8SDQHBdYWt3OzwIx03wpP606BJoAZavTK1qUCd4twT5hf/0
deoZe210U+I3eGFGpH534PsHMMtUIqiVcZF4WmgD9Bgg3Gx0CARKCIN28PyC
Udh3IGWd/H7pn0Dmpo5F7m85iD2Iq6blXZDnUgFfWfGxZPuqS7Q3MBtORUbV
CNAy/xpc2f9rc9y8WW61PX9ApDi6mgnZkQqKZvxY8djC6lsp13xNmWja7Lgo
2e5twl+02QkcTNoTDPGqZx0s7nmXHATSSG9D3W0JYqUIOPhCSsrPIafLhjIX
31iLy7XdvLn9oVqdgD0atXfBV/ZtQrKtjmO18VSj4SCGpdmyJMVr6vvNkmTl
WqNxqH37GV+XSVc0zwJvaM0kKSF3LXreOzU4EHu5QwaOxWRlvt+PYFHRZuOe
VQ5vzztd3mXALk/PuNdpzA/+V2y0QwdbGo5uQNOlqnPqJ9rmhK0orHxuhnyZ
kaaifpVW+0cumzH7DRYRqnRDBcQ0DwtCZs610OtXonCI6KgQO2wVbcCOL6T3
Jqh8PYgyzKRc1nr5EKupd5rrA74XuYQwE7ESuQGQCGBb3Y4PRLin78JatbwE
H9bPlwVmyW8qa4gdw6UBAtuVhj2L7NTeXcRJo9GZDXgw1hXPEeFOzN72JlB6
Uq2xt4Cat3X/5DMvODrzcHQslWCcdR85nqgjGZlxWJiw1CLAI+3pqvvyS3T5
kHEUsT8Cwr0s0YxZ/krapBnRQgLrxi3yZQNpXeJVi3rXHo6qYXcjAZdfCbyW
uh8+y/09dMxbJtagVAmKfebEDOzt5LcTnlbDGHDtHCtwmX5elwo9qGQzgM4U
23+chdzlq8VcwLCuFjeELJoxJhZFdobxFas3mt2KeYeAl7/y5U/4eEA7kn3d
DIqCuVO1yYYrPnV1XYDm8y1os3YWZY2nzfx6XZysItYaoqbmOAh1CgXMDBY1
wO7cmnlFhNlmKcsPPe4tjjvsCykUqpyfGFxIwQ9SK1hU4IbkQQC0mJHKJaOO
pxW5oPOP5Qn1MrbCw6d+X1AJvs4c18mhP3xvYigS+yv6MJGTxMbyPEFapX3j
/3U4DDND4KF7+Df+tGoVYDN1YLVpNcihm6tO1ubj/FcnCziF8mTAUVx2At3e
mwu0zs2DwBCelM3X/hK7W/3hsYj2p4FzQcdqAWdZGZujVhX12Y223M82+7wp
yjEP55sq5X+IW9IHXdNu7gwzyHxmfptq837kX4n8EOW8VpEMv414W/Sz/vzW
evPQc7eu9Iw7STfYMOL0tEIPb6sGCL/g5pb9jy6m4MFqL1NvpanZD08zF409
6MNG2xGHvd82yWm2ZiTybwmcZ6nPQU/I0o+fGxGq+dd7iavmU3N+BWuE4tVq
XshpWCAgype2Qm95/LuPX0KrMDihngqyIZuQHXZlW/jqQm/Hgk/9hg3lqDYg
oi39rYMWu/liIoiThcqxYu1GXAsyEpD+7svO1jFU+9gzQ0K0Q+qunIJ3dQEz
3FtobBrAjt2Duc28hyj2FKUzknJTaqYvx1t0yNoHfvKIn3IpwgT8IsgAi23c
/x7wkAx/mJtIA5e+viQ4qZdLQnjBWJPS+Bp5EWta/IxixCcK99igdHpghW3T
jASV9SNomQZJGzeqXT0+yFNmsJbKe0C0HEYgWPb9qXScylfm9GYPQPkcmbcd
PUS440HLiUUZZApi2i5ydfGiNPF3/5edNfA7RnQ02Ohfn++HW5AfXYsa/cUa
YFfHVdg2p/K/t5ThC5z8kjBAyvGTn3CCNG0uS1MIOL+D6SA8Apdj1NBwa3rW
gWlnG3ZPLs5tW3XmrvKZ/trY+8SmfS2GNZj+fVLbDrG9Qlvm874TsA94YjCt
MaxvUilDGXdG3hPWueGdtl1R07i5i7xRyE8Csx9UeHeJEe4hu+LiVSu+vpOl
Cc/KtyYS9OISEL/9vqnXrbyPFAq0x48aHkr8HHlO0IxGIl5lRrsJXkuthZU+
3eGC3Xnjt7potBFjV30kr56sQH7mQ2qFbyCdBhENyq3xgrftrlXG41OkCrQo
LWDd2/Q4mBbiSC63kiXqBkqRskxQ9iYXm7OKdGcKvuvZdvRlSMDhxWWqMh+e
Ryip7suCE4AHOFWtY6+4YzeL94+E9XYmjzAQhCL2zNuIxUS+6AV5CoehPiby
Rs5XQcfYv7h6aqox+l/Eoxbb47bd7c7XlLPGiZMaTDo5/kszx/3ZhvQ0Oxu6
bX4BqlUVWDSGTMxYoZcsB+LAJV+qB6+qDLDTaws3fA3W4dP5/Yzzivp16CH/
HDDgNct8sQjzVzGRyIGyW9YXcwjdDg68LklgQ6ngq+W8b1GqXEhZUKz2iRW6
A205gtgNV82Q9lRKo0VXO/VBPGjGnwqdimV0VzKU3SlGt4VKoXkEGsFEQV+3
p74mE8tM208h5qzOh5NESvteGB4nd7Pgx7LqB9HN/rJ9JEywKsZ9JUJx3pMO
vRMn7cpdfZSevNOvLZILCSfc/w3ZwGJ0n9WO7BOcSdBY4PZf4SZfapXfsLyo
/jFhwCHEZ5KzbpVtJqGCAmfNps9a1TShvoDIn3AHFPwwVZ+/dJZwvlzmBKJN
ztmb0HY9LsYEZHz303bngvXTbdR5fih72LO+/WHlCymw7ww6zW+NyYjA6Pjm
pYyUZQSNhH0bJtsDQ3isT2VeLXcE3TZH2pRjr8yuFRj9ZiuOhp2ehkJPDjEZ
TrzzZT+AEI8sFnSd7Qrje2bzAbblcSKOctTDUIZBOVGcPn2U16zO3vCREUqG
p1r1wqp53EWN4TsKwZHj4Ut4Y7KL9/VcCStfBLIevqfntsRshTfoBXX1PTEV
zJlhekz392ZBxnpGddWaeojv1kZPhPAVU57MzWbokjp7D61bNiSyhcAtg4hf
dDadcTHElttb7MQSgVF4UqtuZ9PC2keHrmCEssyLfzScbPTgf14X+q5lCUzs
/q3yFT+eZ5NX5hKUbOP9VqeY2IB8nunfEMj+IpcAJBBsj67FsrCSHExt6OtK
ml7836lUIX2R2CisQGiSwrk0L9co5eMYo3t1+GfabLPB9WF8hIG3kjLfqYDB
0oCnAjoWAL6XbEhXyIYByYpVuzn72pfzcz5RaVKcXskMuW1chpWJ2VyiuqUQ
X47cL3/Hc6lp0l6zOqYGPIpy3ymMXDRnb/QsLBvBkpxd3PmuxxeiY2XqIvdN
U8c6fGgoJ5lYY4BmXuxx3vSl6GDRn4toIymdNlnHOJxb7/xxXSpIW4HZkYXM
dq57V3cHQ1DFIE+hqrjd6ScSJ5/jqD6xUdeJFr1wZq3WOnBHxKg54JM2fEC2
O4iX0B8sdUq6jih0CAOasPcw3ZyHvOK6p2TYK7VjQ9+vZbTbRIA1rnsYl1uP
FyXj+MCeeTySnLhR5bqZjZ3HKrNQtVKzqdg5VGwbXznTLNiXwHxEa92FLs0m
ZD9bTkEiRgnMsb9zhrTQUAe8Sle/9AtkSMNJ2bkl1RjGhxxxvCoBmMVIaemU
/MmCwmrL3MHDXkdvEwpW/9LnHAutALZRvHrY0NEc+kbCYAhhVBwzlbFHWB0H
+AqGPX0su0eEXMZEDupJRdKgOGUYUHfVG5n0klaDreAUphR26MXNEW85gk9x
9LG9d+bhwsmjDRrIg3CGP2JI6mgHlWDdHUa59BsGoh+u+SashOkt4j4HxHSt
PJKk3mkSrPLbKBYREb1BGSdSRMdXhtOkvghCzkYPTL1iMFdXcZJcWaaGBL86
pB4w+xBSF7Wd0zZHQszRdkmKpisAORS7xHIq3Bd15/+8pT7ANde6ekF9cCAQ
gyZHq1Fg8452JGHQytLUGoNC5SbujULOa0n2L3lV/zbdYyYkbF62XOTq5TsD
57l/3rWFU6AkMM1CQlRdMW8nun86dgzktlUDOB0KdeQVNZqQkRYtBxZvmuNc
bTttZ4gQazixgUTNtRPOn4flUbBXUE2Alas6/dg8m9w5h72q8KZe1Jjq8s5B
p9RIH1kyBMcisJ3zTjc3nXRiq/Ne6MEMtP9MYum3+zlyAJ9W4GTiKTYxkCUL
8rnmXs9/lpODfLc5qpZkRCsitdyBS/ezVEJLlNaqg73HLLwaZQn9sBOdQaj5
erebAgFC8JE7mExhZd6hE2UVjaUa79ggF0TnwgOGefmGHarwOPh8lS9NjzgD
bfsXwe1oiHbZH8a7/NqQ4U96m1zqcKi18SSVXPrJJSFQ8EM47UYpEo0IZgdq
VP4jX3inNQS8KLnyjnShdjNuilmrn9jxZxqkVVe3ek0WTg5OgMTrGHjDkR22
2GOO/GTJ0pWvGZFG00vVXCpQyatTWTzDf3Y+A9lpxmpiXEIvvaN/sxCHEFWq
ikrOg9dOrI+5ybKPwvvxduvNduN0dI0pkZ+F3HQNx70WJYiCcfhM/xgewICh
31AqHuAR9DAGbB0B+220HZD03TBLJf3CyNoha1xA0P1y8LdrsXcJ6yoBB7Lk
MiTIcZKqmJMJ3W0PNL+fky/q71O0vXjGVtT2kNjMuNL8ZE9D7Ew0Lo7RTAio
URr4dbqDRk/dXzSLvHRHYIZ73vSAgjljgppVdMFxvq6eAXgnu5FkDWsBoXRX
XzcAI28dmx2oM+0hT7q2KZpcyvbTVu1ZiFQ7bD4u+vOH10SiEc22HLxM7Xm4
QAklfiMzedrcCwtTQJkVEA4o3dsQF90Q9TbpHvO0fRhmxSi3k7cJf0gNGHSn
2u5nKz0HLVEmW07FE3rM9acP8sVCI/Jl6In7JsEbnMhsMtixcekyPNj23kAH
oRZWMSMy4Ij9zRXOFO8gxEkNqHW7tAtylyAeuuymtlwhmjvQAvP2ZFO+QKJN
cc3eszPjO3AIZvCPPsAO68JeEbBbtOAJ2VSYohThkH9nel4JOWQUE1QscZWl
JtiBuRT8mmmTqpLf1DjM9ZWjBfEGWeLtKyEzjg8gUFxNqD2GpiS4x0uGGtF/
/SX4gI6GdWwZdPtFALWNhvJU4TRrH1CqhKi/mKM7HDYsDaeDKHmexoRphSGi
HSwNHmoj0/hbxmU3qIez/L+BDffyQKfJW88mWTbU/XhGSpnwqlORPax/7CFB
zM/rZnpuABU4jiQIFDjrzbc2BOODJP7GMiajoyRGjtfh9x3WLOdhcqNJUVnP
91JTgCGmgxASkRHSkAE2OB8u2CedonMMnJlSsQof4VhxpEUB7ZN4wfbm9QXq
XLfzm6tdfAxJDHAUctF2ZcVC8xdQnJhiiG/Da/Ly46AZf3ZSL5dI8I9CI1Kc
P9binWOLkbIsf17mq2wB7WjcgyBw8N0EyfjEdTLFscoHcYpbf121qSUeHgbT
m1qoI7dKlraqVUktqpVkKoqw3igYPS1R4VPisAmWECNuIAx4PKJes86IQXLm
J5B0AZ9Min0dDbpKkMQvwyj6RPsw99S1nDFWC9c4DLxyHmTzjRgMsLChVrmg
dGu9HbWdRf0OlGOqix4jndz9MYPv/yaaOzAlWvFwT0qeZzYBcxMibQ8MhNpt
5MYJGzWbstIZFBbGiN0vxjgMv2L+LBFArXmG/ni13l5lwhGkvO+IpY/Tyaku
DRshb1ytr1COFbY6Fm7FyUnKj+2+/uPl3XoFEuNitPegslcfRbHVH9+8cRpm
+RNjf66OKwdRvXPEPmE4QgwIu39B2kzzLXYqFCBQa0G+JypNzKBSofz7fTZz
fTWkituMCWDRz5KuTEe5JO9DWPeZp5TGWhU8r+Zwgza3gW5xqMDdzQNbaaqK
KW1NpsfkqJt9z+r2LqzZjB80ZbDOfxmidOHPVZNEr4fxLIn0eAZQxGwk0h1u
wzyu6ZlGRnjMmaBMIHcn5uUANCy9ZO4JH6qFX0cx5O8qB58ZFYnjWWUdhwq/
T1XE8I2j2PH8jYbxy/894DyLlKvNAFq1XoBJdu7wVPeXBjU4Qy6ecvt2ZeQm
z69JPqLBYxBS3R3sF5QbZWU1oWxdDBMrcsM+FCrewKHus2jsDKaxDJK6OcFh
UNaRCWADwvHpbub145SAzVq4YOuds9T8DBSP5O51O/aUHeFeaRII3gYVmj3c
1SYx1CJa7kab0wx8KdFkuxtv7ZLF6JnLGtUF/xm7W+dGpFmG+S9RbQQ9IvGH
tajQ1GITAyPdrafoYdx8SzMwcQ2zeiNTgI7Trs4IXjWQgPN39zyF9T39J4pZ
Pz5uofeYNMuqD8UV5s7ClIYTvyhXsOwWWwJoaw1hoJQpMfTEVzrghWj7fzSx
8VhwFiBkdf53WukNVs/1TZ/CT94fYuX5nTlUWFRkpK8IT59fKrFC239z4Mos
4e28T5Zo/yYwg2EJHlN9y+/bPtQKFxvJdpnilnMja2DL3XLXwH0VDOrH7F8l
Agsq9DeFJo/89MMmxXMHMRPfUm+xsecYyMjpQa6O9aO9zstM/NKPdR+/kT0x
2Hzhpn3XQzRSQ+rfLJpNIM1XQ29eJ2BMz7qpYPmpm+jFIYqs7T4ByjyOO4mv
YIcMG+C0YQvfcVTLeDihHOlIOg+jYAa0XavrE7z4CmD5TaRMeFMmjNidp8S6
OxrUUQnwawpBWd3t1VP5+eP5aKBpW2l512Mz/ipx4VbjX8ZqtubLfFyiElap
0GE3K+H6FDt0iqdcOmUGGvoD157LQ9CSmkFs2KYTt+9TAAmI44O82od1pTpl
molSTqF2KXxRxul6SEYduKZADXa1THbeXbh1Mi+BFjMTGcGmp0yLNoKf5Rza
eroZY4JnRDVYDpKZgXGbai3q1EM13TnvFoJvcalxGWjcLUzhEFv/wFaIh9Ku
Oj9sfjhxUlXTGLnn2yAvq56d5Qbz8MjVun1wKemM6DAyYQJBPQglVSIpm+d+
v7dTbtRDbOGgVDpI3ScRyvDVNvm6H04ZR326OmBfKTyT4A4b7/YE46WEIe8j
3BCumKqHnAhwBFTtBgvXcJQHjZctzVFgETL+9R4BE4kBllXCazjd0ciFVypF
yN+3V6A9jAC9ctaDxsDx5NvIAS5QEViVwI1r1GCLAJNg1OXHCM/Md7yHrQOA
Q+Xt71AtzV1KhLaXLCL8GnsWlgMJFXQLmm6EEvrQjGChrmo0ykCxyuOABvvy
t1kNijXRspwrYKtuTnXjkqhGORXowxo0U0y2mfxttuZl6Mz8ohzRZhq6U/Xv
2eGLVltMPUbHV4rnnwHDzo14MDvFWwUlfepZ4L0M8AH5Ek+im3SJCdfxEJWo
6yydkQuDOiNQV/TbDrh1UoKlLZJ1udlizJSuzFblTvNK60Yz3hAV9mKkAJ09
3XWrCOpysIB7fQL72AHb4i5mUIAgO3rG5/6+y1BNAx0MjF8z6t8n1Wnedj4H
gKasR41BPLyKE5+St9EQccQaCe0JMtpB2K+YpqiIE3yul93YLz8A6bTnQPQa
H/BNVhIW4zIRG4kCmCq/9pnnHR1Uejl8FjGsOqmqqKH1Qe01RpB0tvxx67YE
wMkT0ym+9jcAHFVaq9CxshRlWrjjyi48odAr072DpzkDyQ8hSeOZH2q4DFh+
193wgDGBdqUpcp2hmV2PEnL0qqPlzVv+qFf0EswP2kMpZ4KVenHC0XrDF0p+
0oKgBuD/9gYFXfYAFpgT/xON8HZhDcmf7voImQnereUvjSyiKkMmM9NsUYNE
HqRxMGSwEzSVycY8dYrnAZk2oN5g0uqqDHN+zle8zZlndoqMzN6rK2w0d2ag
zUp/pb976Ujl4OVvXHyZZzlnfZEgxoV3l2ooDr27w0BP3X+w4xuoQHlMTYOd
10SF/NTy3+ScxIUP8eAetO3zA3lON9zZTusI5KFNvfz6o7in/JZuTR3RlPrs
8Yy2LtfDu5VKmBNvB2zYOuaYUDdlypjFG+EH/OxAHBQXejzDtqB1rSPNpouJ
mow5BIcfIqQZ++eKfPrvczL0gg4XhY2Wj/e1oOnVcwsWmu6xI341GojRrHJO
op4f5ZCwG8IMTB1zZsYVI7C0HmIeA+nXzHkdYlvwXtAs7LUxcPGv25Fft1aD
jRZqViM8Cu0sgR8LBhb6k6VVyo4BT1P3JJFbTGFE7NpFXF48ETXv6YA7Ae6l
2oFt5aqLHcFnkNrusfutFOASchaePmFuNpgGGrphAZvWyyA1iygEdmW72CVA
6+KTX70mfr7nSfn7WO+PBX7Umjj4XIy49N2wBGVcesDk2ax0ZjPNSD02fD3L
jD024PZqGEbnz71tCJ73lyPz2gHbnaaNo85xtPytqOX7f2sp95pqnBQ9tey1
zfYmMOPBSCRUFoOYNHACu/dF0JEH1HRhXr521rj+LbhquTH9h/8ItS5rJnVN
QVK3p9dGzPWkBoNSfmerKnVN2DSBcB5IUAWtuLTc4R36BXKGrESJA0ut8FrN
GtwpTiSsXGce10Ix3DnQMjC2RHoPpe9Z7npPU8ul4IuOLvo+AdhXOQ6lC5pf
5GJN4KgSYNyBIX9TLlsgr5sYDgKM82mjM/B1mUe7eX4tq0bPONzUn+p5yd3k
D4h1NbqUkgsf/GHvlKEQfEu7N5tDNdkp8CyxDjgnjMt2PaGIj6RbK8u/amMq
2QpkhZ6Wm2rv3xOCQIJ5gzyPP7HQBn8iBsL0HMWnAGyAACpzEVtY1e8jkUxD
+aNKzwHSYz5TIq4qzGFp8o9a6ba1ItcfsTwflMAX1T/JBc2fFW3mRn5M0ZjX
pX29kbxxa93EpSSqjYybQ+Tl+HNv5CPiX0nCLEiGDZ376LX5J2U8kNAdeDEB
/n3jKnIy0J0zhnfE1V4aUbys8hLAJRtkzOOnT0Z0c1Zx/FfB7SRSP2YPyWQI
PgPcd1rZVaMsBWmGi1nCdmDmMDWGDpeNjv5uFR46VEceabwGdZm9gTFE4fJA
9IBr00+XkeBtx2wgIom/sU/EFqB6J3Nsc6VhQL2fNYR5QQ6pdaHX6Y16vGab
Djkic5bu4Rcl2WXK+22NMwVezY8TlkSjdOXjGdh/4XApF35lEKly08tnyeHK
8eTHwySEfL5AZfx5S3kS0bgRy1oqkKwW/L83GNlI8VJjd/WhiPGtjGUpihZg
f/3xpi4IF21FkXjmED7TQqwWIVuO2bdITggZ8Y3d5X/uvfo59/3yJEo3L63q
5ztD9fmnnS62hQd1KDHKkx3QVakl5GMKsjfUTCY3BUnH6/HyiBEaiwQLxctl
uoXWKkptq/XQsCrZRRchQhk3jSTiyaPHUBlOiADh2hQMlyrGfr8mLgCRtdh7
zMs2j8YkVnzuOAmjsrHuuTqih1K1ZfqEY3fb2tx1m127E4g2Dh8gl1mpB6gS
FnrUxGWIMSy3IEH1jURN+HQelMJDHUBZDNhY7QPhLEFUrw3uMd+5qEEOWu8o
nWqn95ajxKe79sGYjfLr2YS73GfGSjpFtsqu1x7dr3WGjHpinicMOi4njFG/
2zgxpiAXhTaxppa361P2S5XNbLHyTLLmxrnuZp7pkgy+g3edvKHbStQGpnsR
P+jv7voCKQpXwtGLoJUnjkNvXgGx7pvUG8IPUm1NncWLuJHGeYSCrl5NbR6T
0xK4ufHomaGYJ1cVE0pgo7r33eLgbV7BQcKVEnKpQfebphyz3cjNRPiUCqsp
t6zawnFYwi2NjMwdKO12GUta3sjBq84mBwheX12/8ftH9LkjDv3FBEBJIRrB
Bi8N2yOWmVK60hj0vtxwKaZN1xSvxaGX3TbctsgInSQzo1dNXoPzMEY176SY
AVnCMdAgYBAHhmqT9pE6cPjRNKUe6UmliDqYPoDKIz/xiCj/zRQzPxJBpW0/
T4jwYHacDFlnwMkprynJUmq4cgXAttmT8BUM4nPO6Qc2n0CSo7EwWWHYTEnC
7OTo+HM1bYWeVMYRaq/Bfwkj3Ok6eJZ4Q4IXSuCyl7aHtayaPw23yQGQ7Bmb
SM938cGEBllqJ14WljDViROoFtNuMg3NTcyU/sKCrYpGi+7PW1/Ps0bIt0y3
8QpzGC9XbDDiofkQvhVAgIZAzXUOMTpkqq/5ICWCuh34gyza8WzJq7CMkOzX
NQWUpsM7NQGlCFgTgeRe0AmzEJ7VandiGKGfao6z5+kP2Qn5ryPqDPzvSkIp
RG76thOJSmyj37tixzUgVkLI80X6Ulfvgh2X+biVbNmla54yzlniGtMVJ+pr
2ZXoR1+pMnskmGzGT50FS96+LRw6U3IXSnsu3nHFQbS05xJZqPwMfpPN3ial
4y7gPQmC3c7dknTfIOUrRoJncED7RcvtE2FWgB4UZ0ywWpyKVyDK/cmQBSjR
XXya+aWGir7jGyZJhNHiB4VNgU2pEiinQpJAnDzIvm8mEhGSFn5TLBu0yp/8
3XL4lljct21HODVuNRcDd3MrJ2RYWIsQmbF/LpBSTBTSCqUEiAEDtFa59XlZ
ERhJcbvW0FzBrLUNaxJoG38d8tJITfZBkEqai42RoMJx2agXniH55qvxpIb1
EjQhAzHo50joOn5LEp91gWQb4U3AQ9v7EVWGjeiFFOUJHSXDVOFWxhzPwdlU
rN80w9RiWJ87HdvKcsbVcpunelX1hAv12CgHd8k9oV4C5JBG2NG5YCCErHtK
V25roycppUISGkLFGAV6nPo3Q/g7DNDJEwW72VOcJfC7uToEjsqPtB3AAwv4
bpMKllrGLTYAPXvuT7As3pKxpSfa66PQKSrt/wqf8gcPn17vbLi3uJpfNjuE
4ZPrEe1tOJtyGETOh9mvf99wvgVkVlyPEoypeXw70GBQK3/QrTw3MBNcxwpl
h7MsNmOXffcLtLOfber4RdbSdl1TUm1hjKG2u8usqN7iWOuXkJYXcWYy2Ioe
f5WewB2FJvIaDoVbyilRpRR79cJ1l+W3dR0lizyjOMPhM5ViwYb9Hb3MYXIF
IqHjnpCiezeJM36alXEOgd6d9WAakwAMKqBD2kLw00Ctz7F6xVCe+Ez97/Xo
xXSc5QXAnetUPfL1SjEb+8gq9wiUQJb/kc5FAS8DPt2jte7naXj85Aauamqu
/GHcpONRpwRfALDVwefWbqiVDoxPHU4dpMlUUyGtxvydUobQ2r6o9FomMmNX
oIBDlwFmDqWV1w/4616FeWG+YeRjQS/H/IUbCFu0T50YRLwTuscNfmUhaUOA
XzQTN6jf7k5wV2pKAP0YslqiyqFzMZQBrU/oVMkyBnk+0t2B99PT2tIYjbZS
Uzcow6qlJy2OxCmCUBrzdmoBNitX3gpua7Mh1Zs5m4cIX+tyLw4MrOyz6e2x
+tFgIbj/BdHGfL8EJ9jZeYHeCMZNh01+CEZMHG6gUSHoEht2tv2sja4PQDuL
qDUMAHqYnKsTP5lE9AWhiunkgCzu9rw3sF7gU+zfOLVwai/p3/DiW/cPB6z9
Rjs6R7q86DraixQ+J01bYMvdXh5glqhCpGhR4v3cMsEYXE22ObaXlRdrBmCp
D5v9lkwqjdVz2392ghN/YIJQ16HENxL4t7OvMAqaamHJ8GGFxy1F/wYiCNBE
YZHy1fZSSyKzIPBkdIfneJAo0IF0hFKANAJEoTcp4cEG0t7r5ZLwwFJxKICn
GINX48o47NQiE+yqFRp26g7tnondKrVB76FLUbWYnU+bdh+pVzViAh7rtLTW
FaR/2VMbITbTDeIBejPYOputqAr9d9ABm+zbyaxqPqm0BOSUFDhhDmlmQHwZ
AhbmaD7XlYpTieFzxpl+v5mRkkekecPS4xCvmyFXxDimeQDTYr3yb1OLo/2+
PtDiAsNrqqTa1HA0b4EyaW+yo15F8miF0nMpJkCeVx0QOag4AH4skR5NVQmx
2bShJviZ7Uj87PiCVn4BGXxvh2dAofwu5+Y58V+b9Nro2oSn45m3HkO6uNER
8AHVjW3xl/nV/knpyAJ/su/RhkUQQoUb/F95lpf+X2zUKt9GV4WmjhzVoI/r
XWv4H/Ct99zVhQZDYUuGQNOhVX24xGAKKan/TRmt3/2rm8Xb90/8Amr21GYH
YhinhhitJGiYpBlNzy0Jf8nGfRym6xBjO754bLW712/6ZFVgmKwVA5MNIl2x
CQxPQudrrR2alT4vc8R3Kj0tQYZsXSDQwMczucmecqLYYfWaWILGRMJrngkR
B1sn19nrT94xjGNRF8YSWgO8PgZYDzkO6CfP2BhmFF1AbTqjLjqx3esBVSnb
v2sCHg+++H6nRnnlaWDIJKhwtGULhtEkyAhJf22pCtKgt154H4pukhF6RIqI
EPHd/rmqWQjA+RIO/3GncAvKKnq4t+sT9bcFaXvBpbS42Q4VF07/mK3bAKo7
++82QSvuiMyBB65FWb7iNXrs7+W0lv9/kWw6uB3oVFFbQ7YLLEAfxppIJxKw
3j6ykwwRNznDfYHhGvOsRjgXczj/49DjdSUwolwdE3Ot4ykEYA+bl6zopa7X
Dmqff9YmJf4agA1/cWhwTxa2doILk2ow9pgFn8HarEs93/z/iH0MJ8h/eigj
4W7PZbIg9E5scFx1n2JYBGApdnEOvi9G5L9RjoqpoSfV6qXSTaZ1iFfQWjS8
AFHsXygNluZUxDI4LM2uLUsS53ZCvP6Rl7nXW7tqKBEiiYTXkOgBJeYhuDIY
992vzG6HUJ8LbqYc63/Hnj5KtG2o/KTzXRlh8QphEdDlBvWs9nCYF15EEyu7
ChF5wt3oEzL2FJDEHkC+tCD9VctmyzpL+DnXeYWP52lSJZpjVrkN02zJ9IJ/
sNLlM4bhPFVjZY+pHD+8eyKE9O9DBp2/Ra/mEMbOhrovsAaJmgwz5ApL9MrM
G9RF570SdoEMvT557hxLVoJ0MaVSf7R7kVPGM4/qC7s9PHVJRdxr8iJ/s4jN
piM2DMdGROZ6GvhOLBU0RY2jUuClloKmihYz1EIYKwNFXSfIVEOhvcIeBAOp
uttu8dAOcYk0qWbQvm6ddkMBg8lpHzDQ4zOq400kU7sFLccHy3Rq4VBbFA99
fQOBIJxMxKsfTZ+rFeouIO8cUMNS5oYXXrqCEWXTemrRP6c51306kh8svc7d
+pVkte7GndxZwZZvveU/AlpiEPZbQAt7B30zdftkkK0uT6VAXY/8669nNy/o
OHUSqoZgdhXR2630Z15onV/2c7dkwF31sJdw/y02wrIV0h+wKB5KtiVFIYTp
qQKcOflXKpCVcDkkIy+esQ6JRf9j7IGO4GY73mDvfQh579JqmhhQX2FXze90
aJOJqO8Lo9rrgGxzlbqP2pWo95Fu9saLkt3QxCuApJs0wZjkkbgMrNH7AuGG
zyAHWSAD8pSiH2lbIuwrNbbYSLgv4GFb4ugqM3sELTtG6XtmbCdIlgFDIO6e
ZVrCs5E10eqWtT9UPmk7D6o1L7SGlw4G+8WN1+uK/qSNNSqPAvBhcasUp4Bd
sBUj+SIKGPpq6g3NN5pi40+56fHnFzvCrOd65H+P8wnWTt0pPGvaSgP3RUx3
Tr0BC0c0t/G9ju+oHGukG2UGJXtIO2ViaBH+K5+CleMykx5f5Au8iHxJB2va
HYHKWSz4UrH1LbYNmOX6RBAHVew8H7tS5YqqZ4u8ZqbK624oQytyutupOTMq
YjzNi9+YVIOLyRJ5SsUMVEeECuhCRX8WBUsqhdTPvYiOk292WS2f8RLZJ1TB
iGapHA0AynvLlXlpcbp4lX1iNcMbkH469fo9zPQz2jbO7K4NMxA/9xJvRMRj
VHrY02q7V3L5dRzyTKvlwcjhIjeiZJ/R19OwiX/aCQVGZpAfb/IaAwyX9Sde
if8FliAeUB5Hb0HpW7VLJ8wJdhEEfDhaFtShR6qKhBdXGDFVdE3eHdh/O7V4
hVJMHgyxhyoUIJd2q+gbN5f/EbL56KosCcXo+xcJqNj4Q5Uc+x7/Sf+GDoVy
bn6yHKuAReM7eZ1IMe3iegEvLrKL1jd8F2dp06H03zpqz5gRsIXfaL6rRC0z
uOK3hUFY4EcRqXU04HCnSpaIXuWT+MA+m2NDxoSRGTZWJJ5IKwnQMezMF89Y
8wKU/yUqwkSeK4BrxulkSsUs731MGm4ln2Lf9gmSssGcUoVJl6Ms33o+t3k3
O0V5rdJ3RVXoeUvX6avo0UjxDhjFqB57GiDykzMhwA7hnuL1ClIYyR9uPLgu
dCHWKzd/uymNFmsVO8D7TfV468w6tYr9JrHk4Fh1EAFg2sIJBXzgPNQA6x4V
YTSC5bJhOMhVmaXIPjQOswvko4SjLu1C5+XnvKIQ73+9w436KnrC+qnj4212
6m57zvV+4ZIxcSTYfWIrtnYuBtnr8Sle5wELBcWxzMiUdMkNkpZ5EXRnem5Y
Kj6qcw1uhip25n3K0MyHxAVF5O39K34RcEwOKklJrBbbP3+GxDcg269n1dAx
a6+QwnAI8YdKUZDuNQpaHL/Q6QaZK5+Rb6mnO2aJ8tABJw0Q8y7gTKi99M+o
fcWtu/7AD4BIisL1F+jETSJrR4cjypTVqM/vYqu2hRwQ1G2WNqBWvH9Wpc7I
nFNkx48hFN1e37eP6C9QqNjHMOP/icJ38amE36edtsPTRHG8abOZwlVYWitz
2e2rgI8OvbGZD3h+uyUkGfWHbtCRtoQ2/3koXxQelUvym54E7S4jzkqfYw0s
Nx1kTH/lZufKnb/gcH4fxs0TFJ07MxSMTNf7DPtstS78SNnxWsHNMaJ9mi/u
tSytYD6lIE92/u/1xu8c6V7qX0f9ypnZPRcXadgwXoX2GaFfY77PipIJh0l+
OATIS/LBqGzjqs8W4fSxm8g1I5/4uYVWZIzeZpkuPcasf/T3HoiqT+N498Xz
ewoCoZxWjD/SA9nlWXME/ZctUFVyfSH7et6/2yIm4o8ElLdpZRkTpAMsX6kc
vQQ1UHoehNd0UkEfeSK8w/1tvl3XSvcpaAvO/8RbE/rYoYNeis8gbmZMy2ei
J4pJxB9Bv7HYRSNNs8r/dMwBGQ1Ydd81V3SJ3KKcgf01ADRHB4UAW5tH1TEx
uMrLjunP0SrCFqutp+qibxjjLFWF+gxiHzEmhR9hMCiNvwkJHTR6QdnjbWjx
DMvGD5yQAxV30uKb8xlOvaqw+O2WzzOvlsj0Qi+5pMUzeBoRzEtepwr1mBGA
wN2+09Ug5ijBhOKEllMatWlpDZknSq7RcNwmeSm2wJkE2j8HVRFtGhYJwQWD
n3gw8c+j2FtcY2ev2ke49Eu727E4VhqIyjsHrtjdSeB6D/rNJdZLNPR7UA6A
h5Psm+1qiy3fy88F6mFFuSPImCWGFLFve4jC2E6HFgKB/Z+NI7Lzbr3QqVWg
dW4rpn1vYNBn8E1+J+8KHvXWSDuUu08Shr5By3M10Rss6rxqH9/UWTixDB/N
9XZ0p+MPF2p15UxTI69/xJbWzW2GzJGu1tBwKu1aKRd/evbu7P0Sy92jhQWA
Zu4YU3M7puwqabkHWXYIY1ZRIQbag7wl+oOVe674guY6VYihWkcLHV3Kj8j+
RKBCvmTCJI+t5GVnGANj+kViNGLvyU72WccInMW6ILS4zxsa+79EVA7E8A9I
Q2H08ZuKMgxT1+wZLN6dGmRHDelYPSAQ1NRrYGI87N0h841i48vMWLNtllno
M7dwWD5af9EG7pBb6zD3nuseaI2Rp7ydq/sWadKsCxrwLKAM3IZcYyBNSdbJ
Mn9hlTpC36E5va/wWQoLv6mK2WgU/wjb49vJY9XbdOvHKd5QTL1faok5tCrc
0j0TogfhB2DbBXqSZYhbYmySCtjga3jXmrIcSRowXQ2cCioBvBTV44cYSlTe
yC+/2kAtO9Bh2NinbOZrOzrZUrzR5ueii0+HgWv/6kRrUy62lTJtvgDMPhl3
EbgBb2tS3DcWSsmw6xdzb8FAfb/Pu5CJAQLX/SeFKryuJ7Zck6WAdP3aJxxq
cr7uuj085LjIw6jYCTFjOJ6A8m1EyLdyWiOYdz9IdqfUu1/jv8PSxJ4V0wyr
oSo+Ya5o5L+zAUdxSe4uLdnLjT1zuJGP7+EJ2YP4SeOakoHW7k90+dC0qo54
9Y3YPh+3laTqM3qmwIfnrh7u4j4r46M+2qtTdb7Lqw/wX9ebAOFx0d/k5Esg
sLdp1AaINJK1jULXm9g1Q35H/YCkz5Eo1T4/TEvon6rYBxh9kFGFmU62KhMz
tvU323WeypC9s01oeKmPNDCux+nDALQauWmzZ1pG/xOZdfb2iyBnVCgPooXR
im/D7DEheCCTfcC+lKYrCBBiTUdS+5brF1Z4v5ZxoSGS7qXun8+JcSCRCZFa
GQtWUBoXojCMs2D0PnNFl6rvBDMn5ulSXGOKlYq0mqdiHWTz0Bf74DEEugKb
hSF1ww7b5luqvI6kQY6s7EofNlLmfX1xXCRxrUDWHQbGp6mRvbtCugQ9f62W
O56ykdSybO2Ewxugojv9GQEn3xFs1Lvb8+7sW028oLQZ66NcnL6We7iwPrxu
UhKGoVUsNHhaI7seopPpKmth4Do2vlI3mT7LYLK/ZC/ulxSPd3k6ydWSTMwy
9Y33fyEbe0mS+1m+usT5jNyVDDQJV4jqtIqyzQrMxVrSW2O8L1DxyUq2mfu6
jaGJ0xmBxhkwc/H9nmjlaK2cDNgRkv7oHvy6WtxFJUUVSO+nkC4CrGbRPVLx
eMje98iHhpNo8TCGu7Ors5+H+VgL7kwe/QavaCyX8Bpg/ipDUmla/ZlrZBVh
1h4ZtfpvDfQuohz5O7RNsgPJFktihZ3RX/0URqTWAL8K9jOecg4x+niK685y
DMMBGPcIlqyNsyZaCefimU1UJaq8vT/xHl1NT6my1slB71cXPcJdeDVNSoT2
AX0JBCJiK9pvzuoxGK7cVosNv5SA1P8kHc0ZKYkVteDFD7df7mxKHoQ3dlYl
klh1iUQBZ7bbmH66hlDXIHLa2fsT7lxczZoxZBco4DYGk9mq8Z1rkYZ5KfLu
X+9Uw38MFs1rgqp6BsF3kU90vBxMicnVRzLs9gdmf9pvqdGHSHbMPCAQ6xho
pWw2XuM41YLuBxjlss99YQ88/PcPEgPlYTZT5C0TyCosOVzEqKw/UbpIq1N7
v6Vi1RIAci23PHR5yO+PmVTrYQMOdPsUUdgFcKRqEVAW5yxmWOkDcrFXeA8e
H/YZwYtMlCXsvwhrGhbfQadz6uylZoZbK4VV8dUuN7klj0ELOj/SrR+9eeaY
+MD11H66EPpmhir8gReCIxygDvvfts5PjbE5X4qaFg9b5TdfWeBrGfpfYQ5n
f6T12cGvSpsk2efE3ofE3rwj7wUVagNktsGxEmwGKY7b+ylS8yp70348wr1u
H5Fb3n+ZZVZsGgMBtVGdSZyVBy8BjxEcgIdHb5k+TQULIu6BlelpkHn4SYYO
vBTwTxeeTFI8en5tdmEbQKxSIDrNkwxgesxnOBJH/f8eOklB1PmF4cO66lVN
keMzk+z+OUChcc8OJmLVuLI5/l0+iuTgckZDgay4dtqh0lUjc17auxdB+Hc3
nhIitOX914v2pTphZn+lvlCkYvOATk3xv0bUz3glXFAq+WdIuQPWVATfAhvz
Gkrqb6i4pqUQSkI4dgp31NtDj3QHTFlU1PBdZ/6kAlvKP6YmiIuGufDEe7je
vmzR5u1Yt8PjhVqERuEdpc68qEhdRhL9PD91v0wDG5E+sRRGgeeemSBiJVFh
VCiQDXWa5Y1TLb+98eQV7WLaXFqxCNk4DzJhNkjHEhFcfeVxAAEsLdnXTxXV
OvzpaSi61yOBoY7raT1Vk/lIa7kawAAPu+AzeN7TPmsrH10VjhCNCTIMan+F
9Woi/ldIoTDatszLfYp0oea2G45Ijs04qUaDQd8BwNn48fiZaskZZJlWjErC
oSKX8oiqhTyMIL4NfvrgBONCm8IlJwVl6+xvlnDNjlvay/Xx4PB8o/DnNcdP
IvyL1jCkAQy78tEW2hPQymKtNSIF0rYlAwgnwaVXeUx5m0xBDiDgko9ZDBEW
4UrKZGqPNzokug6YrUNXe4PjUg8/zv0m+hRNwTdGAdzYWyuDafS0ROJav9/H
oWqn4TKYOySITnqxQeGZ56pwKZ7fIeLE3ecFJKFQg4nb8ZJSrfpJwZFBZhL8
Uck3tonVIbXKZnWjl+6iJiXaVvaXGiOUloOlQn57kvsJE04f0Hg+JIBMCwlh
YMF/+9JpiTdUHRwlmmi954TJERZ+BUJggr/wSQ2PhLHv8ho/2ei000VshBMN
NmtK7vaTVfF8Ku8Ytn2a8nbA73pPAC0l7S9dtYvuXf/KXmtrJWZJuGp0cmd4
MKF7D4SDdmK/o4CzAaY+ud+tCgFAOWBkdzUuUpMRpEeAdJWQSwxhHRqo4Fk0
5zF1CWTqcSnf8QW0ZnHqeQ15aZAgwhjRaBQgrMyDsIIqKRE3njWFPMyRE+6f
hqZd/zOr6sEu8m7cvfld3NuPAY6IGQY7tWPqlHTACm2lxGCnsxlwredhjKT1
x/IqSLgzjZ5kcDEy9slfQYpM5QnD0jTCcptsAjyW+RHFnE90awccnDSgHywZ
3mT9myOqrWJVo1FrlbuepG3LXwpmwXRffEh6BZFCXiyyVSkhwDlxTIkz8TKY
s5LBsJGVSgbms5MXE+Fw9zKUbxxe1V5GZX6LDMPf9Dw0Ezy0Y7U1DzT37HzG
dXjiE17RUmd21rReYsUYxkUPMx/rcC2Wljuj3h7Rg7hgyZZdYib0QVtaW728
TM0sPMAu5RIXXo0GGLZUTlzo1I2cl5Z5rtNUsfOq8vMt1/JZMQFTa7aPdFLa
L/jPRr045/VNyq3hKSZq0ieopVRn1u+PCuwdMjmFbKLQxUyaZhk+qp7yMlJu
khyaen/4CZ6yL4vkj7v0/6ANE4Bb0cz2gV25Q21z8BtXGVAgnkJkNAcmQn5I
szWOzNXbd5V/oEN6l3NXyuWg65u09kYWjuKoj71TGMPlw8t0CogmygtnNyoO
4h/K5HfNDUj76t8rcF3AEWmohcMFbfeYqlXGp/IsT7DGLTuBm5y7MfanEOnt
A0cNuSfftr3i7SizqbbJn30VhtUXUxkON1sokVQdJAnEArZkKcW/Ja3eY+j4
vHxkWhpvmYOgglZHfqMqf5r/wpih3AQc5lKIm+YE3TtgBQev6f0kmxMrI8Ci
1Dj1PvJb9yA0fPvJv/RXDEo84rM6D/AkwwBSuVkwjm8RoqJjIYIX2BQWNRRh
hy6GqU31cEuNk7M+zpLs/CqWpP+jvi1m3EdkGKJlZ9rHsSmklb0fns89VCJ0
L5cmW7sI9bRbEhOw9BJtFsNU/fmiQ+O47sXn9naM/+YJVxQcqdBiXYfsarNk
mdgQv9p6DFxa1xIe4NutDZvZWBaVaUhGZOP1fqIn10wgNXs8MWHLkjVVnxX4
lR7ewjtvl0wB8bU8toCbQHeYIInLzQeioWWo2VlOtbWrssuZBZZICC1uesws
aE25Mje6xd/nDa1vEf14hlHt0V7uAnO4n4twOn0x557+ky4uPOZqiGHGBJVV
yaaEKbUKPFUVQKonCC0PcSc6iDkIi5ZwhZcOg1LqkoaiRM3P15M8I6ig0Q6r
ho/1VeBOFVOa4VGEoxf/tptCtLuxQiND3tnz80en6hf37iGtbt3QYRja8tR7
Tu3Q57Fl3EgzM9zqub3khIA5UG+wsNj1EsLepneqCfJWA88NUt29lJLkFoJl
QYWZ4v+dzZuqHb+Fm3LKwuMczuHY3XKANh01pmv9RMHzUICl5IP18T9ei41x
bMyFxaFZ8U48uGYC/EGpWVIGSt4OCpqjZ2N/JgP6jDE8pj/N47ZogwBiHvkc
BenwifZvfaXcK2d/GetRPL8SjhHdEQOAsEVWWnj3ypKeHdcz/pKTk/7obsyT
PlDgJpVB4al52z2Gaq74j/nVESLMuwqVp95wFjZL+F2hfnIBW4EYKeLFqZFs
bkiNCR1PBgQ6BmRxD70JpgnmSmO+QQfpj+mr69L3MLADrjuHkwX2nGWjT/1q
t3uG6WlL8Jubb2QwvndnJJ2hBjbjT5kAeC3JczugcQ7AyPVAOohjzaPB6WQD
LQivqx2tDh1yEXdOmv5hFwCGsNdl/OBP5m5MYXBR6OWJQF6Gg7WOcuwVicpq
L5cePZIMUDYVhpBnwZ9oRjvqUfvMXqH6UGLVJsO/dsq7lH1w6P/7pE6o471s
+HUDeiqpfJo5LFZmH1Ox5dBoxLp/Oie3MH1oE0EfUlDLFzeP4CT7o8C6ROaE
0XbKxM0au4SMQGnTlrwFq/RpebMgEhAOPpVsIN79y6ZjqZmjbNgqN1ysq10t
+MuCcsbPkwKwR17gCew6ZLVwdBRAtMYftqqGiuA4lASc+gnNU+wz4WBEQSbt
IQxNQhrFJU3nYQAREhKaQqaRjY/Nisrz9RXJwggln9sokJs3Ts/YeWizlVk9
GEXGVzmB2jd8dk9ExC7bTgiw8HzKXCw4V1EOV+N9s42E+pvhuBjUJkHYbTvf
VlkqclLJzMJPh8pCV0f00jNVvVeiGuahEmtZCItOBD0BhR/r7YrJr/SRNWHM
COQ8BsBGlI5PxmNw+GikR+8xpyA3ytzlzRBMKHWoKA5kCt/MO2QsV72y2AzL
pdpVNTV2bs03u1F78iA1oh1TCWhJZpb9CEGipkIIygd5gnNFTrT5VKuCgKpE
iEZJUbaDODJ5Ej+R0+03DyixGyuXkQS3mGvA4tPSqzCYrVXwPHW8Cn5LbXyV
uLbp9TFaGcxS8UEBPfzWkkN8a+sc0CVqPRziQaBH9SK66l1zGhhBXocKguFj
74tbm1kfGwM4f0Co5rXv0I3qso2Ook6tKWGJk2INkNtJT23kQHGjo3jrFzcz
J9pGlinxs34WhkTKWqdVc2LFoINBsXAqiZaItFqo0UgdZ9AoYWaMLYgU2rnG
sCqMCQukZYZflwSahgpLaw+YrkrLk0MhUC3SWAp7ttX1tTLun/XXc9OYy96D
fTJqoYCztUjl4nfinJIcVLJnh+Hz8Nd+X4fRDAOyN95DjPDuOE8FWtBwz9KG
wBNbr8u7tYKMUHXrXtEBMwX2yt2yxs57XRVOBjVvpA0k1fkpyJkMcQTmDTxB
yd5HsCtBmZrG9wgHXU7ZhUvyKgRR8b90fJbnpPVsbyndr7LrUh69XrYRpLqH
hPdXla7PiuDlNJJf/HePEKA7GbrUXP7NDyc3LplRHYlq8/GhjF7P8porlhss
uS/pW/SbMPvCyDZUpKyX+9km6MCzGjQKta1lcPuAK6MBLBzSx/jq60ebW9rJ
l0tYL45bJ+PZCfAt8HOXijnIg/8n4NC7CGD0K6hVeHSTgQglSZG/VY6q/33s
mhm4quKT1EQIZG8Uo9UNAepnGKhbnDqK8DJ0OrL3+mnlx9PRT3MPAgqLoPRM
SRZF1vQzLYBKzUftRI27SoKSqZA9qPa1zUKosHMiOpxk/qSi+IiaxXKLHYA5
2Zdt0zT6VjkBNnBYCrcFrFaeUD1/UXxTqPAXt1Tdwch1r0tx2xMqDARG0gu2
ZGwmOW2Zk0iDV7vM3WeeaYEFGAnG0gkVp8vp2N8N3sNHXnRTKVoQG2Hng3et
ucyknPsexyz+RBUjm+KX0zfgHS3T7R6YX8d5lh8p+lkt1UkPhGLcdJ21JEZg
KkHLtlasmE2qETChEqmxnqAXqfur3ch+V/zDPn+1KY7WYW2FS1EHPMC5VYRM
UMir9/yesQ5zXdSEDnxAiH9FlpP8ckK5OF3UAxGm63MCoafWDGkq3P9mD8d/
97YjU6xjUrBomF1wT3FKlWl6SCiB5veFqJ1bL0Hvm4Am0rM3W7ti4bROtm1R
T2i+ZEvjof7pS0PM/YcXVNWHMR256fWH/w2RMxB8bFTS/FwjNQ4GbP0DRnJo
WwAACOc2RYivDMS9aXcKruKchJjpyiHUtqXquJGIG5eQrBL71VP2+V5I3KU9
TS4m0cGqswEpF3wTpG0TEg4jT30PoXvs9dA+1UTLrgarqoe31cA5DVlR0T2u
r2p4t3uHXKJqlj2B15zGZOCMZ/B8Y9JPCFchenNfq/9NgdrI6TTrKLxrBcyL
kwKwivJ/Q9lG6YxXU6Qdlvt4FKkR7AfpB2PwXvoVAfiZS7Qjkg6O5z2tLNZG
hvVZYsvUp1YiejadPPNgcFjj2jNdwAxPSUsZHBr3Egi4e0HtmY7v/f1ervHf
IU3OPbAkIZ7q5gDP84rzYNulUnZM7VpiQEcsPagFyGFhuQowDLBEIPVgMRwe
GcVWKlw2PnKuvdzItKKguz/SSbfKWwazZu64EEALE8yb9n6Erszt6kJzNFAJ
8y0+jp8yuUAMY31ff7N8u6Xn4Ik6f4cIPZfua1shdJZUGalvP6tf+0rigLvU
MidUOU9KA5q32Uy7S7oZBdzGlKJW1Bzda0cEKBmktnh200Pfb17mLGntnv6Y
yuRuNzHtWrhNdQVeJSNCTNECgDmB+U/ZBjS4p1KyyLg49JGne28N9MR8wV8B
BCV0kbKEBYUyiF0pdITtv0LBj4lM+k9Dv3XINmLf+eF6bqHh1qftRpJxJSwy
9JTjU/5rKbgiLptm86TdxaUAiH2bTcWuZGckR5kiJTuxd5gH23SkmBLvGBic
59m/fAw0crjgXCTBL6kyGYff/6cFMveEIcwxpmdu4xSl9lGyZ9bdKuvjycCF
K6bWN7pfiKgmnPd9ObXnXio/eCeyqC6c2en97C/HY7mmrqqgCTimp3O4bZYA
eQu0v1EmLgOG0XlKighwskeAxlWIhL2RfrysfyL9srZmQyWh6G7rt95omhbc
MPoZiKAO6LmgxVwTOCsE4VcTYovixDKt3XD0FEpBlSESVD3dP4IJvTbEqe/5
sIso3ETTcujMijRh8lyEhQHuEl4g14DQz43CO+VERL7JBp6xsoyFEdmdbhhl
O6yUM8wEjCB44rkInzNSz2F+D7RmN+B8uadshuuitZeJR7bUtPZ4TKG+m9rt
Frj+ZUBcV8Bz0uiuT2HcezpC6wKPRAEOZtv0A4W6JcnV8MaTClvTYd+2RlKa
rx5fWhq3JRHEpn6/VWOKtCBRnSoOujqtnqU4SqWhCXfIgFk6YWGm++EczKXb
AN0NexraLmqXIGCPcRkuQ9goYEdcPhq4tZ/292qJSmrmMJaBFL/dYkhBlNz4
l2tPDdeBfXlUfYqlHq0R36CuREHduIawEjjEx6poZD32JSgrlnDYv9PzJ8wt
zCndRq1V8NF2zkzlDyZ3FftrZgLffT7WF5j0HsmMzZhJAxwOiY0f0fPPgooE
e4uX0f2HaRHRhml5wylDJuKka4NPnLm15eLRUHg0Sn28WXt0u2hkPmic28pN
CEtC8q3Rk6WWiPksvzpkyd2QvO80PB3RzFNOrN9ZdW2xmPM6iaeSS7xp8mYo
2407zh9vtKcWZI/Xl+6jtF5QmcVd5P8ovAtCEeB/a75FdmjnIOciQMDhEi0r
UTQQ0XZ49ucWFpCJXlHWJs+h2vR7AbqDlRN3vVWX43nW9ZInGIPpjCzID+i7
wCYVR82l3GEEAbcru/cWK9aMyTkNkFCXfywMeIn5kJjEKc8psNz4ltzwyQ+B
d2bycwdApeCk7t3PWrT6smi0P/qJ3ktQHmz7yA6z0JQ8W3Q0OJWl0BJ0Rh0V
TbcVFA9xKgTo9ATyRN55vLt8bDuZPQ0xkvvbu6SBWziWnyBQUniQ2Gw927xJ
HGumGRLk7U6BmNLq6FGlzmCY/SXKmdYf1mc4YPifjhd7k+Nx/MVKxkYlkaZc
caPouXmMDC3vDH6QpklKyJJFkZb0sBcYNlxXpRtZu3hK9YRzb35njapwpSom
Dg54uPsQA1xNUK6gzVDILCuFViqIs/2HKDskSEmyeOXR7DAGuIL90x5si2XF
IkSFVvvqddwuxNA1FYPenyz09MWPvRnHU+iupb6RImVm/iMB4KvwZXF5XweB
pXWfqi28cW6A5kenDyFasxENcFBge8gSvU9UsPTjynpbYymLdQwaWGykSP5T
nGxBpEDxUoFrQnOqpmuX61W9btH1RwF4DhzpsFcbBMcLZUrDMtNquScM+pDs
T1p2ijxRiVsLPfwV/AqrqBgdnBf1ICNcuwQNn+z8pbPa131daEoBSKdw7PyA
mryw8mFFkfPUEBZDVTtug/kxKPB2pE8KbMTD6NGpt57WxO+1ED/vTg4CAqZO
ld6JxTEDRqPYeDGL/oWZsQ9M7PsSoqpFSkGsRXG9tNZLqr82NmvVfmbauX+p
eSYxJl9TNsWTqW8vbGDW0u09g7vteT8JNtjIgBsNekrcNCNv/eAjXZvgbOO6
yfFmKLe8Lve7ohCQU6GtRhW4NpCZPkxgFwupaRAozNwvleDJQeJ+r8fNbJgw
/YQnAPh8+2nTNrZWLapB/K2E/IG2KpcJasINbUe8UxBKjO0EzBp4xuKqOpWC
xEOt6bx5j3lMc4cOUApZR65WtuV1JmM9e9QQn9SdApb7fv6lJfSjC3t8j/tH
YiJgd+5jg8yn14dyWlR+/KkaC/TlH1IFCfSWQZMxHDwDhmJm4feiu77u8Rdk
5UOr4ZIniTQTMFKAL/++cFGN506uzM29AMVFvhlNqUdg0q9I4ExGj8wX4dqP
kJgnvO1Ug6LmRcvnAgIoRJMZ1iy/M5zW93hklGMM8F6mMGp2gTlxQrbPiNZr
SFdggkTQ4V5HfyrWoO8jLNcRezWt/tpkEw+327w7iNP4tAVhYUDqOVtBArQd
n6HamhVeyQOTuxTGCfRTaMvos++iirRZynDUL+wT5kPfkfH2Pr6pzxKWW+Uj
pk/y5V0TEkP+gQ2sAoz7cdv6gWjQeJuHWsDNphzXCXA2vw9kKQSZs/I/M2he
+db+eZb8kgqv9T5ZrUpiEUyXWzzgTr9iwj8rznZgjcPwSx3Yx7rFbZM2q2XS
yigMCx9iWbr9DJk75bMW3/ph2C+xpaDXoR1aql+Jy7hC78UqJtA5hD+SeRG/
i8yRiPGsWLpS3oIPIcswOebxkMLnFPfhajIYiijcZGbpD9zl0Dsj71CQg/oX
d5J7EOuouuDILELe1w8zZwQrKCCoMMSLqtyR740KSr4G51frnwN24U9IqU4e
2uWtm9utb31ULdA3DogStK3ZrchGv0O+faFNQx+vQNwsKF0S/kVjt8Fc7eVd
xc8HA67dKpatfu8ilMt70eeXO8owu6pVjbUUyV8PzDv0YtSHmCdntqITiSfV
eOVcXKfWxLg92tmORKemno/XnExZBASnDxUn+UnX0ilpKbvuXbJ+xd99EERu
VvXjj7IwWsNgZI0Y+tRJvBuZoI11HIgpmimjNVfNFcn2iBPv+bgMg5sKsDH/
/mXnyFavZTdi+oXvXJStyz8ugvB3PqJg6ogaWqVehvfxvuunVdTcFvfhvSj5
LlCBmH9SqcetLlEIyliSqiN8OvI8W42cx8QcGMzTqHseXI0tv9ONlS5/V3ee
JGFzZO0gf/VZfC9hKOMYGUE6lx8Yb9fIw1ubsYYDgAD6pCCgDNYj/Yl3KqJT
dxl01re83jbbQ5ZjMisJNzwE8pTaOzUbFkTfqFdiFJ+XMPtg+rnSsS1Gxd0w
CI0aiw88XObP6NdTrsiLlZWKO2BwclWdTlA/HY97YEnMkNpcmbtZKSigpUZX
P6zPYufbeUXRa4O6J8MzkVavDrOyQnaJw7tTZwBD6H0dHOpGy87UWtFOr51W
E9W60A7Y4Oz821J15SVwzZOSIyp0OONGtGdPFH82yxAfrJTDulsCs/psVISS
UmWEu0DhJb20jS6kaM+nf7ckyvYxSCAEm/BTdsCnL1TI0KcH25AIa/6nRnX0
+whqGY3KloZpVlE5fR12V452vgy+j1J3Xns8QV2pevQMQMrNNKbxi5QGBqGK
ZJpIqG2lzBV4j8y0fNdekpAtnNiy2x6oMzg32ZCuKpzNb0GimFpRmkTLnUXF
chUR6DcQza/czjJaqsAlwhN5VHAdaQn1O394gSVuCijMBYieS6NXR+UuhSLK
6gcP+4m4km/lSkDa0YQHpOfLH19T7RGAtzxhGmo/+PtPtSpW0+jAmTP+6KM1
PaLp5Hk8g0iFjpHHS/SiN9q7l7Y96JXrQ97OT8PZ+up9estJL60vKlqI4BFa
cD/pvLJX2/NLDzQP0gVZQsgbxtb+fR3D6JfAF7MUcD3bPfE/cv0WRJOIx3SA
WWNKIvrG2hiIkKdjzcUoRNIihb+H5mzozjqnPABVLjraIPDrkXyjVxOBKNXE
88dPD8DoP6RT8EyQ72/Mv3LCc/p9DQfiof6Qu4AiIG4tSixChPDDtlVqeohN
bWEFvhXyqj2MUw2Ns8Fo6x//NN7YALE2jm9n5AM3KA9Ac/z4hzulVvAhC18f
9GpVkzmyLrpxXd508UWQySS3gz4q9G0AozUP4ocfjVI7TJJLh0TWnXvMGOMZ
BjxBEU/UC6SlmuxorRT0onc+4XNsJfvI9OyUzk8C3lxQOd3rc3v07CAZwKLs
SJUiWck7e1LqaSHjfYTq01EQ9JVxVPJQaKyw99IV2iQzQSinL6PLXmXAJuJh
0kefVoBE/kQJumy1zAvPjEb3hQRPG+I5/rn4oY3EJqn9xx9OwAjASS/Zvp2+
NPzyxqoBiLycDtreMh8B+bG6ZQu8zyrjwdGDLkgYxdGgoti7viv0dVijvbAQ
EebimXypud0whnAIMXdJwl5GUZewBKVA7nUvSU1pfYK/0mYAc+MnKIlIn0Np
yk+tjLZ+qYjAk3X0FGcWOLlQSSSCeLnPLpzS92+I1BeADFp7eW+BqCHkZRJk
1Kihles1xGqN7Kwltf6BsZeVrL69bKNq59mSj0cO39kL00GTDPtvtB+PtMm2
OGITK+nn4s3ABkvKe4R/kRi8enRxg+hI8Vd3tn+a7H3mjcDfYk8s/neuMiDW
MKaenQIsKuNeT2nN5NntG8nUXEWnHZ0iyGJqPdwG9CVjTtqWR2n6ui0hyNW6
fVKBsHL7HHLYxzOGZLd4A1hvoht3/qErPdvcYyXQUVOlVdUElxcCVs4Gap6p
Z4TpDf22GDgi/9F+fYtVyxiL78xnui1txBMECrr7SJpEG7DlNGdlUXv2DAOu
qRWlEkkBD0dbTTKIZipZ5R80rhLyKw0N0xOy1yWyyKThI/GAD9JFAnTLZsPg
Yc+uNK+TRs1ay7flSL0mMI1SnCUT929h8QnTS3+E3i2RjA6X5NZy9l14mzNu
4OVRsI/OC6EZoaUozQUDBGrwNLZlBE5WtxTCmNQ+giK12rvgAe4R6WEYmo5Q
AMpfqbxn5/AnwgIcuzGCxuj4/USL3NIHJX8HmjqeX51AB32JQ09yfx+NIVTx
1KRLnTp9atrbGAvTAY2SgwoW/3awCwJV+zOOt+mIhi40Vk4k8M+nz7tybUuB
kww5/moFZS49qxZ4/pru2LxAJkg23eoAOQagLSX4ujvdxkHVw2R+FiXyMU77
2Q4egGDyztPpeFM13dfB1T4ijpEW3e1J2ECvYbXnZNtCaLMaqHtAVM3cX8QL
0U54YMUx5MpNJt8KFqd+78sq9T2macWyY7VDAZZmQu8CoQrBiIRP/SK2plgH
ycYrKkxg4df3WUWIAA2aJlBXokIQRTivyNCwhB5Vf8CoPHoOd4dzvfOsdp/M
UFA70i/EjjUnOoZzNva3aMcuFeNmw6FaEUPgPVKYMypNN1DbHBvSUQwXat2D
CePGEiKknqpVAvZVGKnpSQq9IFSpXIuNQxfUHQzLcr6il/r8SButxn4WrRDu
+ntze3+I2umYc9/mwhDH76WAuEgACdvzLqnXdUP3SIdNHqQBzzNrllMTXnm+
iEaXhjh3eZj57T5SXtyAOCFJ7mKsyUTLrf8XlTbvh4ojKhYLx7HxLphjRY1E
gohrkvBVA24bKg5mj98AfAHuY6yLliPKSPnquYoBB3aS57GCH2dtjJ585rSN
JjCVg27R/+ac7cAr4lJz6KjPxsncKS3UEXf6sIHUGTTLyaBdxnU1lbQOhbb0
Hl7MEENCxBULlcmk3Z2buHDbcwqaYomf3I3B4MZwh4yb4uTDYGsEt+Y40yFT
BNfXtamVdAMloD5TGakE+GWWqFsuuGALqPTKKbVfya9qC73jYLons8f9FxEP
Xlo2lo9O/oLr1PGyaTT6PT8pBOMD1wVlgfNcY1dXNoPcfi8eL55sKaqcW3hZ
BKnqS6ud/UPJWVbz4tafT1xcPyzzhHPgj91y3ryV2HUT7U8XO8yskiQPFiyH
2x603e4nKYoP9xL1UUoWznH0mWcYazIvwPNZUVRs7xr/1nfi/GdiwKaHeWY8
VpB4OGWQ0puctFVzDuH3nqgGeIF/KA5lqczjrT8fDRyiVZ4PZpoyIIvtbvJQ
CieHryOwAdo2lybnoKIeIeCxOjxcFdDPqIEgX+DUNr8Qz6+kk5NlEDN+7duB
xZxYHd2fwWAWWYTIqdnBMXFpttIApb1eJEEkBX5/UcRBzWjukGNw8qVShJTd
Zn+E38GE98fWjylixDuxFvKzXawXVWLlvTVIF1jEqTsocmri5rSq9oesABg7
Hq/HIHtHZHkHZHL76rnlS9vunBhgat6klWj1wK4GLx6Sky7bc0Q/9rkgIEu2
1NyuLUxRS4f3801OLQ6PrxlZonzfXi+LvjsojMpEksZfEDh031AEzXAr1EJ1
UzDVNKd0Icqqe0yOGIZd+iKDwKPninQZQj0ZOuPpCS0omb53hPO4UKC7gIO5
df7fGXuVfisMox2tOOrLjimr6nhfmvhlb4M6J7hvng3UVvK+UQPiCDpnj2jZ
3LYVhjtDCBLMRX2saZDQEjk6h/dWrv5mJ1M6YCmyBVJNsfwL03k0H9fPpsGL
KffP8fGwrtt4WrO0FlRt5D2AdTYtehVM/d65jXTpLVVQP72NODivKt35nIkA
qFZOZh9KeuKlJf03lML02/4wKDUHAq63Y6TaWN3nqdtIgg+cHquuY6o6Xav7
LEn8kM4S4ShGxj9RxvcYxAWm7TGentlIU1JhheJ2G409NqqhUWIGL7qKnGWA
B9nHtatJNrec2s2XCEEW/AGKXe871ufHs4aeL6Sgnl+pmp1iEx8IiieNg3dP
VTfyQCU7qxOOsZlW0xYOiwAxkVTYeTkWvar2tQNmx8qifXsLy7EY8Zu6avFk
16jOlKPNsTMs0CF96yb11aBeYLDbE9N7ofgAwPzzPR6q2JiHTJ5FRuGNEW+5
iVDTanLVbvAsONC99QkgCKk0lBLH5B2rWIBn4a8JKFXDhFBiQhHypOAw/1w8
552CkXVi64NxHc69vgMNuDiasxrkxAVMCJySfIKkDJJ6e8+BI5yqNbDVKKO9
ppbRhKVhN0V/OdQaS4fGfcKhnH3GJ92SrN0p8gF1tDoY+wdFvXJ42lq5DZ7g
83wIetHnM5dfrGfZBrOiUAWj+A6OLDujc2JfP/xsduE309ruDpW0c/T+eQb2
PxNDSiSAVezzX8s9JqphunWq8RGqkFHLSC0aHe3OVf6RbjdBWmDWsIcbWGeW
YoEvXLtBkBPoX72uU4/NLkhujAbN9QdFrnZ3HPkMVfWO2XqmWV7HpvvrOp6C
ljUNSF9hHwmYMBayDyFFEdrOdbtxwzLpllY/JZezk879vfSRVidiHovJPpUl
giAzycLsFlAUzPYS/MDliOHcRTQ8No/2cof4QlGhEt3nIj6w/J/gXaacift9
92qtngATaw1C00ZHgFyVQEzFOJMy3c7VIbUayoq8z2eFAgQX/GBnPSbWOTQ3
Mgd5uxgbraqKifbcswVQ0AHQo5GHW5swLtGHrAHpn9di9P0QZIia9dIlBNHn
qxmDLGJ4kTjlentHPzgSMtSB1ybe32l2ut4eq7RoNqmtw1abookZfFx5LRK9
kEc40K6T+FoVdGxGqJNxca6z9FLumnpQhKDNlCzyWY6bjvqCbjZzLUxaMCpK
n6ILPYMKmVSHnTeiuhShU7LgvQ038JwhLnUTOxEnksVWgOFbfqBtu+RoCjc/
YiGli0YPBn1ncTihUmIcGO+vjsbysLHrYl8kCENbuLaVXfWGtA83aPn9pwTp
+/HhCqzJXl2GISdK8KtA1Bwxu98X0JM188lxt/2bBtuAIbE+IvVjK/baFgj6
s9cL06HZyPyt530Smt1ijTh/wFiSsJftUy0eLOXJUCg5PqjD31cUVMRLwMeb
gSdmV0wrAZECKXxT73e7ct8IJ1c/P6X2hShhp4ca+nJgda0dNwazFf1EJUA6
RHZrcuMfloIWw/58J+ULdBV4BLsODoLxyPvPwuimK3ZMEurm2/5m6bxwpiT5
NN6/cIw8tos8qsRoTD7AxWZ4V9ueUQ1wfBYNSI0Mt+z9FR1LC4Dn4a/wAhq/
OIOAakNwzXwF0Ysb7m8r8FInIp8CEV88IrUjLnja9vCq3EhGg+N9oyTVWzUM
n3oy4vAHsPz0yiHlu0LqluZFYUEdHNdXOKRHGOrx96X7h5fnpKEIfUtYbYYN
plFocQy82zgypW9sYiIjyOVuMUbIsQLEQuZMwyLMrkq3AJghVZt6vlAk0tDY
tHwO2dhcyuOyir7aBWvXbbvUlX5X2gVZ0KqpXM6LNweU9Z6RY0Qiq169Y7K0
IYHhhlkjTRleh7/H7H0ji71bFXIaLX2NR40KwLOpyx6W06UAnTmaAu/ddcoG
rgQ1pc1i9HNUarPlp1PoZUzEWQzbBnwqV7m+XW+EmyvmAZicsmMYcGccRuy8
2dE+afk9nV0aWg3KrcXDfh5ixkbUeIlN/GupGbSSi0Tjo2aW3WgueJvKs5Oo
OmfFa4ezeCw0Yo2wKasVT4B+bfAsZZwaxxrEOQh2kCcftc/iFLL+YmCIT55y
uzVIQOR+/VcvJm+yplU+GqO0IiCI1HP8Rb6s1/Qkd0V1iey8Q74dVmDIuxBV
CMavLZ3s/IQ1w3TXBuz1nrBvOVcoYlYQUBFN85/R/KKEH8AspSncBF/tlBUA
VTGRodz+qWaJRnCd6+Wz8BPMfOEcVqjspYuYAJc40VcfafyaZztMrZ1scwb7
JGWioOZx5JJQPLGPVeUm7aPgZwjixqfwzJxaGQ9qa+KJuF7kqD//rEOyd9lj
tWGZcaNnWI9ivyMWThO9zFUvUwMIDMuHkqJfgHcvpMIuKR7eJ01DIE2x0eLb
kOiXFEUsY4tf3kTxRpjNqtVGaBxK0wWzhvmdrmk8JgcG35AJ3MZApD5TzJ4D
rxObVXhh6OKuK3P3dxvzaVVPLYN5qSBUU/5nC2ES9XG3fQPrD2i5z2dIO7mh
x3ynib73bjS8gDhjAZzdTSX2puB6/HcCsF9+BkV/WVfb5LfHpitTwP/w0WjP
mKrOI3GYjKpG+dRTzzfnHTnZVEHDDLYjmUuefVs4Z8EBStL3mWFd8bd+keDG
61BNNRpk2OZV/G0s6SUDf008wCSECcJgN+SjCiBSKbDZni+EBdEs4hFsBT05
U028gvyMZ7H9Lzaeyu+ZvQXLf7CvEfLsa+N8RMlLfJ+CF6x/Q5EOEjcnsvUH
VS/7I6Fb6iLETfs9JXS2FGiNSyivDbJK88TYgevej/jhHhC/QlzNGggM26wc
WGR0VlvMOt5A7cYPxAf2Yx9IweqXtWMuUlnAcubGJVjoYhQCTD/jfvSrdcW6
DjcA9ljEqQTX3DIPB9tzuCqLlbqSJCa2M24TOrZHnejD2Jb8b2BKeY4kXvYt
pHhzxxk9O+buSpsENYAqVNCaXvZWA8IyXXmHj6rs2zQIm6oN97irLhNDiSl3
xdQzldUGtPAHbZrTcrD2gnQ9OM+E+RkeDMS+gb+oCLDZRAWIJiYLozZo8pQs
Hshpctl3zK4PEazM1JN6CIdFjme67VNWzZZLrOBCD0FISPdOrb/FDivchXqP
AFl69cd3/5/UmHDCidTF5e+W1N4hAGRpaODR7F5JfdqQVU+CJFNlvHt1CETQ
N4u7o1RRIhkxDVE710of0X16Lkm2fpNcIqzI+yFWw8b1dRQ5XNwbr7NFI5Uo
hBbgKn9XG0X5D2Yv46yS3DbLVEwJPAXQMY7kwNfo59PI6CMSHh0UsLHlfjn/
GSsMYLIMo+yQPl3uER/FJ9KWa44UlJRQhuwe14YgypaGQve6E9dUgbmsAjJ+
NIWhYshXBITSoeWBP9u+aqHq5rNxsX+1IvHUeNy+ZuOUIbZ9hM1vjQgdC/VX
a9Idn/+yVLfIU1vRvSYgdJUTgm87/2SD5vD7TIvbxGCs75ZSGQ/9QoQCB8/q
HJiwUBhUuGH34nHOVZOUwsHOgJ4tZDDoA7IRescBgpkpVjufgH4F8UaNKb/L
D19QvPTpJOp3sP9ujq1/gKDab/FiyoxFj/OkM+T5oZRmlvZlmVG1LsCM2q2O
2gIgPlOv4vbUFJpUwL6dJOdSphIrj/wCzU6TV/6RwD4ampOUIkGubZzHh9bn
52qpaBLVsgKlZEIYh82B77E6NAZGggRkOVO1gez5ywhRWWMNt/B6VJcvQtff
e/X5lxfcw0G1ijMkRbRggkfhlA56DrOR6Nyi2fe2nKLFUt4tikrALszMfTkW
s/6mY2bt7VV/sD3/pbjjZ+Do5B/6aNcASA5+S0WchE3eDsY6nOJqUcda23IT
BTyAz+rl/tBnsY/TaBzQvWbF4MBvTiMlPRMss2ob6caiGoSeKADHw5SEvYGI
nYmsnRd73Y42xn7Gj6LjnfbsAQcbsMEvTNjSzGg71RZBAaay75yoZ5/0FzUc
r+MF7/OZL/s+dLKlEl0J19kKhj9W5gYVwAhpdc/k2lBz27Q5u7Kb6nJbEiUy
0I8elxpmnvVmQ9nLv1sJEiMcFieYgyOEA3MIbJglZvYfV08vzithkCG+avr4
t9yUbMft9dBNrKSKtRvMmHs0+ms7iphP2FV0bWetE8tDmjNWzS6QpIi87laq
Ceos1qH2F5PZQJU8GxEyommwQws5y6p3CK/dp+yoCtsJjA0IAT6WBN6085Bt
DRg1KJw+kBxzAL8yLEjodnC4OZQyru42AbsT0Bm+DFU+ZeMy0zQIzFXzS0zH
/krCbnLZY4nRr7K9n1rXaEkPv7TTNiDMQK5H30USQfWZwGBrznTU28zag7FS
qXRDPUyMhnFH9DHXCRrzlCvEyzkcIES4YRK6XsTn2EOfzPkgUa8Kd0HuMVEU
wCsCIGGYvrRDyRiEOsCqv7sJLPviieXRVIhPgo6IGUfPw5BsvZpKcJ5IzTqw
0yTLtpV/jAdNSjuhanA0f0latpgHbxProtbCzJqeu0ngCVtO1nz14xbNNNkt
Vij35MK406o0fzmHRDd8XqCFm/C/FuhKFPT2Fsli3ar61uIh5q2nPXCGqP9Q
n1Mk6FdbA/N0kgoQEFi0aonxEA0cf3TeqMdZ87zpbcclQ1j8E1pxYiKODOfl
Ldx2pkrm8ptnKCRtFaOn9/mxZTZAr47D/diikfZiSDqDd7F3/LbHsCwSPr5A
uA5R9e0XH/fYqeEjsoI8T+3cB7vc4+/RdKjyiXnrjxemvIoc80kF5bN8DXLJ
YFoA/j+D03GJX5sS4TUMSjsytRFg7zO+fSlxwbpXT4Pqo6koZZecwjII1fOP
y8tWcwEOTRvBsvUsnzKJqkMxAp6oxcI9HuRcv3RYShDt2OQARUCPemG41FBR
Skvl+6/eNTM/TWGcjBwY9nYZhs0/+2/t08qOLbIpVhV/pq6m6aJxrSjMqqRL
Nj3z+oxiq40V/rAVvbTYH1BcabDaihnIvGhUQA6ixtoY0U4fajoGwnBFsnAc
IzyMRLzafOhbSjIlvFBDQ+LDHbQsUye607pJxKKvs8d07A3QjdttQqkFi3gV
cmeaN3pSjhTXTkb5iEZhlY2gUXmx7wVAkUYN+ttnzK8bcaPLB4Pca9zu6wXN
/NMxgRtxj2vIKzi4wFFq0D+l3jhGPdkXPYSKCkDiCTa92CvtRha2lCOUqBMF
F48JLQZU1uXM/XcB3AN4TrUkAZP1b+lTsss+k3PKrmEPaAshVAlYuGyrfhgZ
9j2C//V4mzqAT5XtKcd0BGkLZTFf1EiCiPBD4SsiIEpUgJiJJYiGh2NqnW4G
J1KNpDFrQGbQ9B9EzfroSmyS1ymfvtty8UWEQ1WeoYOH6Gu8puyG3hxQbOu4
6q9E0dqVlw1a/WZHiKR2vg4tRm2NZzGAvkdQEEWNeR5ItYe51QhXvp60QsSS
rouiZQV+hY/pw/MzxwKLRLfeJwrAv4PVOt9EbLFxCcVoq5iYNodxeus2muiA
l1OVMuncOQ+p0UIIYglBJO544Q5UoKCV5VKomquR8P/vYa7jKGDOKUouUmYc
LCAIARMiLVq0/8lJY+CXi4PibGz47inythwGseQq7xGz+zZz/q1+yFUlyrFE
G3OfOosJ23PQX06R3dPw3MIsRP0Y0VHH8F6SrMl269F766o2G/nJmwbG7f+t
WcqmHVLmnxdNNK6LfMEMR5MEKhhXRNHdALl06v95H2swtRZ8pxINOCd3qmNe
b0YpzXbbQzZu4WrDh23bKOvoOVbvyu9GsFtgyts/+pp0xza1Wbk+rSOzoiyx
L17gYmRK4/mK9XNqn1c70WC8BnY6qmpmu8GxN1b4XaVASC+1z3Fct+9CplcN
3aeFpnrBUjUorDPcp6DSsprQCGz0O2of55orl40Dp8fStZEHo35r9EHESZiW
OScc0fw+UcN9M7kc49KumauwTciUizFS0xLaXkAN3VAEnqEFStqQ4P40g1TN
F+ztVfdTHHuCzblxY4vdRHr5dp/mqKeXlfAQdvcnc4I6Ac445egqwu1tKPLr
iY601U6iSE+oai+MgYIhUOwfO+dqybAWY+sFFxvPUDbRNOElNoTfpoyWi7y4
XBkKxXh4P9HXW5++87SBQVBURk5QyR8jrXeJP2UU7yOvQhc+1m7mhdXPQTPV
xBvM7V+xxAkFY/4L6GZOuWdSnj8ayFSUnUZpWp/0WQZ0+ueKd2MY7J+uVkAU
gO4I5ZaKm2vULZ0YzwSrs51cAh5LVwUNxpWl9pMOlWYkAUfEczV9EyTiH22w
Z+KO74LJ83fvjwJdNBIS3erj3Gt6Vk2HHIijRhq7IMvfXGQp/BMBYxG7NPeU
t1kuizbmfGyV/Zo6ql4tAnF/mwcq8VD6eWvmMplpOOrj4VO6h/MbR9rpwPad
FMtOIHt/wKu/97a0E0UkcAeGYvdPt9nAU4v8mOv1DWdmEdDFe0b8PTyrNP7t
ORbhfkC4HrMjzdWvpf/b3L3whB73IMwznPrdqB8yw6EqSeaklvEhWX/st8mN
Tx50MDW6rXSmJ50ZeEcu16LR17eJobBqgzt0ZPUmjgKRX24bdOm54Rn8F/rP
P/qNH/UDtCCA/FdIqqxZtrPBAwhTlnUJ0kqHEJCiOSKArmEHozpNRmzlT3P0
77XQxbZWuX6HywCoAIpKb5eEf6yivTNcPso05DBjjKKjG6u1aCtBee/9E5eQ
w4bj8PTEzq12XlydPLxCHGtDbbQSNjZ+2IrHjgGDOx/x5QP9ptKzjsi1Gq9x
lfpvPdAQ+IHHpDRStjfJtx8tesobjfyYemQXydwnsIOv1XJwvn/NytgFdsQJ
iDDluuXAyMC39XPIVjqdhw1CtdvbIABjD0pg/JD7lVGGyu/TWgTq3nWcWA9v
V1tx4qd7dEq83Xg2w1zU5J0teZguBU/GBbl1dBYzNwhRrzQcUM747m1/akll
wwaCbtJJsUFsR0hDbA1baryQjZG2J24yxQmtcfP95Wo7TF7AoJZ7EEYmLOnC
5c+KsxpVc+BoJHnpoUWeazqWzLIwoemsxLH/VCm9+0V7qehDCjvir6O661r9
nwD+ugaK3t7BxXR3hbAxTS/LAphT5S8WnD8LM5it0UG/6TmLAFynALch8n+o
ZFApQNIgNwKPe/DPrv1+TaNcfHIRlR3pnI+57jfq8EuQw53nV1JnUq4WeiPB
VmwXY4Lv/cGP0XlQLsr5ehGOuapKY2xvG/smNiygK6ndSeJw/wxvN32dOTjn
e2of0GUwpUftGrR29qujE+lCTl+vQSNtRQoA8/4KDGAcPdHjEgvFORI6AM1a
mmC+7xGeQHYGI27Y7JGeS6IvfxtPa6HbcAcWvO0Nn1tPxidD3nJX/SEnkm2U
9spDaVAws5v2d4s+YNPRlMwJT5E/v301mS6iCDqMTUl6TQc48oC/PsCTwkhX
BmBe6lmS4Av6DBubckbaARWbPqTkILYBqj4TKMh4R275Gk/Kna8GszeQpyzN
r+gHSjP8ezE4kxdEohJNphqhBfPjIeshfIv3bTAWpkc+Ck9jWZ5u6RDAeLjm
7HDDQtfvr/e+8u47vW4K5rWm/iHZGwaE0ZUmYd3VDIt9gBjfoHIVPsXlUT9+
n9j9+oy4uBuWkwMhXr5y36Ury/Bpb2ieWBI+t+xGgq1zRXYZXBqsCpsKaWv2
zlfJNCYiy0OpO9QQSx3TQGrwnE/NjyGYlOV+anLCLBzy2QwgToDPw9fXss+0
zAgm0gUKtjeL5UW/mmIuFrNLVAria3uHFY8V3DkVDzDXvsOF9c21TnX13KFh
GfJvd0C1Z9mYuFQ+a33sS0d2E6FCti8NKGI69WADKuxZRcrtEMNO6ow56XVW
XscQlfZxEEn6HWvPIdLLIvYdesP6VlP5U+gsfWa7ZkJZnXUoy1ziK7JiD0rR
ZujFCVAehah1BbHf47VAT7b4V2T/ec0ErfuTdVPoqUp5e8iLVul4pc4wTyna
Geu+ots0PiR2m3rgXbY8vZzY8UHHFaB7/1BKD2dsnRmJq6s4qb6hjIWRifYk
7eGYNyoSXu7P8g/sAsilisKT1aNk761C30SfRPVzWQCnkzwWGQqZd6t1vfH7
z85rD9MBi7Yk+H7x2/YTe0hK2g6pVpUC4tGt5pprKBZJB7GAHzlQQSuSVSid
uSCtPR1ZWiGfEN3HcduUAhDLVCLSkYkbpdy7Z5Z+Qmimi2w7ALSBNR3kJ98w
pNkRumBxbT0mzSQW4W9GYc/HnR1F3aPVCDCXPpXDNvTBcL4xuWSjDi3LALXe
IB7VlebOmts3au9lPoGfzhAP06GvS7nTRlqXEriHoT8eBr3EybXthasJPEdG
lCaTFKcXVk+fQo/auOmbnsxwxoeKEkZIJUnuZB7Qth2fxu2Rbiv5UDGUYQAU
8iLIvQiDeliRsnfpJOQ4dNYC40UnXwRKPGqQzWSs5s/fl52STmj1ncAFxrLI
NcWYVZ8w0dZp+CEECk3BINCkQvW1RMKGRWJTheDfjBsZaxHX3ytsV/0NnreN
m/lMFJZqnOmHOdbteG8GSEBGclAb4uIzPBmhUTsp070k7v6swAAPo9qChaiN
VNtt7+mL0FvyiKP8ojzgnZNHRABNbqvvfuQ2fuWVRGAzznkNKqm/OCFC+vVw
pBfzW9Iibcpo3x8OC+dN+woPwlWk7h/z8kXFHy9qx2TVs+9A/q+OzLecXgxS
MfcFnacU8oCQufFDHQQmGgk6hGiBr0aUmhDIL78T/F1u0woCpZfVQZloxy8r
syp/yU2DCxeVhWdig7tXm8L7QqtuisiOz3FoECQ8fVb87ob7ksqvUxCcdoCV
Qdhsy0U5N9QTkrz1bJd+bmrDeK12c3AhrB2XKbg8wp/ey/tBH9w6SAM6P4Fx
xeAMUdOQc+yJ4cfrLOq6GLcd7gJQnbYSR52TJcxt+XRiK/HX4upmm/16FCDW
LBjJwzbb+mdi8O4Oj65vv3zT7FrKwGCN1vvRd55Km8KqlkXJ74/49dqtkL1K
m8UYHG1eHhb6gqpINqY85zQUhoYjB0glw7OnGLAZxt4+quZsuU1TuJqASiNy
XGXXa4MMeN2hswZhYn3oA3gd/3O9Ym/B0oytF/NA17N7RKtnUqiCv2vmVGdB
7JVIheLS/TwoDFhYxJfJUaf5mGV/G36T6XfTc03Nvbo436HOnmlJEewXfFru
BiKsmMT2S22TRfNQL4EE8VgSib1FYu2zBZOTuGrgXQ3l5usMWJWcs5ZTtZR0
tZkkSSWdO/39AzZlbeE1lsalwtP7cDFW2T/LzIQZOAqzsEdyYYRgA9mkAw2O
Bzmz2idIp0uBnGC4+6Z0EZpx+FPzZ7rU0gdk592RYS88u2GYWgYFQlEzMr8/
T2KRgLypxu64cuHkmQxzo04xs4lR+oWQSe3dS7gQWXtat3bAiWp+j4bra9T8
BXFgIOQOO39OPHeMsWl171oOIV1AAiOwoMI65alIbtWhmFc7MMUpNS0fgR1q
xTONNIJXP+xbZectgIAPkAsQa5+V+pVEMw/yfkBHle7ZOInmrA4Z6Hs9HIwy
hsMJ1BcvmBt2pjlHyDgyR8gvBxKYK1+tEQGdPaFKLWIym9jGo54cCzGe0Ps0
8wVKCFRjkQi6Oyxi3Q3S6s37sc2wOVfWudRvfywsKBCiLHuVhCpMdxh28fje
EpZrxd4Or4Z+OqlDS2dDwzSWFp1Auyjkc7DYIqLgZyjT0XbK41WzjBZH0FdW
2uLGQ8cDF7rNeS9C1j3mf5vVnGIDaQZQYE+DN37VLNrfG2r+W3kYJxwKp6I+
LaCbJ2qcwQtKIfQaO+GE3VOzrOFU6W8A+b35zbJs9w3c9NBsAJuFT7Okk+2f
voWOhZDFsklpGG6PzHoOWz5X7LL0oF+yM9Qwtllsws9RN7Srb2p22Nf9qKvE
WKnCiYVTIOqGMzPr2/nM01EM+c9G26xio+mYOVXO+IrWS71WvqddgbsyauDP
t0bjaVJFj2IDF5hlK4iGYS0qG9SqZTd2X1VckTZyvkgek7jsJMsQYhzAKEJ9
dZ9pFnKaoHkTGkgxjCzK5OIGR0jy7t2RUKROp+3rX21c+TZ9wfxEXseg+GjS
sP5NWQxC98RprWjpdtEZYdfii1JYq45AEdNT4FJ5sLS+3B1HsQBOeiCNrudg
jSEHtaXVoDv7v5QVX6OV/akUBC7WkucEr8wnR+w9+TvYyF5UehfnvAruTGo4
NEaFSG0lRGgMOOyqPw82NXWhBcswZpixz7N/lPax6dNmXiZ2ic/CkuXyoST1
hL2qf2PE4cFwNtoLKNcXZ7BjI6DoJMTZx1TC6B5vQ78tmrCf8xGrs2sPL1Qh
NP35hE+lBvssrDTDr+uIiakywleR98PAHfICspUB8hQfyiQVZDuoOZTebcYj
zEBX8WoMsetok7tOsUvGRKfaWsAsV6we6m1yzxkgpu8zkBHE2J+iFYk+c0qe
mozovLZWt1FMF8KLm7yrR4p8115Hd1zf8IcdKKDeQOr3C/MSw2dvtKKRY9wy
m4zAaDykLaqlyeztPmS+Kq0QvTNHjR7QCrZNB8HcVcImNUrNG2Pdz1JtoxRS
z9kqEnXDi1pUvvG3wSbaMA8wkw3A5R/re/V+xoWIj6aIO8YawshaYsmheynp
HW6TN2krs5/Z40+xuj6qcF7cCyUn2GZJSCYnXAZci7QueHavlMiWTZjcOhc7
ewE2qOWGEAd8deM5ynE8XbgGDp1MQAdZEHrB75+0AzgJv2Chl6X0P3vxusNo
MqycO7V7hdlCn5eergnfy4hp5SUx9Rve8dEIGuSiYvuXcNZ5/tPDL87tS85I
4+zvd11s3uwQ3gZmm7+WMXvoe6CkVzTTqxtR0qp87orMviuM382LUc2vvZ20
5jaxnPwCr/H41hjpT1ncYqGPoclifaspswr6rEIs7vrbVliK6tohDg2cy5mW
LBUunzqDxDR+tEq4iX0S+Ft7IJdEGpd1Kzr2wcSR1UuAwakeCgm77OgQSWx0
dqZWX3J1ieEzNbVeUj113y7zsw1LSEgDeviBDcNpCf+Qa3DXluo3J7EpmlCS
ytT0xwwg/Yif5P2byaBaKoWw+LnRO+Mq/UIqtma1YuWnJYfRC8lExV9juGn+
TjUwTbu4ax10ETP96TkajOwuxvXH8m+pdL17NvC5YAXSD2KxiyVoHWOfTGgP
AD+Ylf16DQmLKza0qz73VMvVFGfmBMSNEIeBwQTnuoEjxmP7gXZ/xIOIiyxM
JmyA5t0MHvsUBLPio4hx1eUmkimVRlY+Pah8FA46wvFqQiVjgilzUbVSS2q5
Me+O6/qrb/+xZgOLLevjdYO+KIF97iHIP8uy7tlc9gVoEeol8Xttn/8MxcY8
I0VrTYJVmafpzb/4Tl1RI2bxCbO6JonSMCp329OSUj8M4TN1R43ZxU6iyHpK
N1TG3MRoeZvRxuHGBXQ7xx/17wzmhgi62TIMsXPIpM+k4CD4crCHzXj413Pw
3D1crmWZQNdKHfO3vi27hOdFmy2FEjAhnkDCPcDbGySoUAnmYOl6TQbE2mKy
keZY6sw87jHr0enU5ng2yd4ACiWLR6blcP1uG/41s1hrYNzvmeK5QfoJ+Y3I
++qU0dr1af4tVJlUtdUfzXYb57EXQGxUoCgcO9RlGSpmE1hePBsbScQLjLJS
3IQ+GY7HUziOF9KdafWu/XFYATJFw8ELAuiPJygZw+lXr1M8UKS8WO+QTIqS
wme6SIbkRpuk0+clXrCgCn3zALHKKl46yarpjynW0WsS6a85s1KWeowaGdJV
wX1unJIze8ri70G1B3IPLQj6zglbkuzdR1KHrnAzNQ7ExWDEif0D0eELaeuu
/Um7tgDV3CTkhoF7YdB15M/I1yJAwoAmRWRiS8gkiJkNmyrPEVAFh2OoDZlr
ETM4aCJ0I6U7BvO2jkjw1j+w8eQfpxhOSrezUN9NDtcGYCLSqoYfxtthkLro
91d5kFnm+/o5Pi/lXat3ngZrKDKJMQwYh046QgtzfIihYl28gTvGZ3LAJbNS
uYl+DwAMU8n+axqFAH1CcBmsUxa7ZrGYP0NvxS2whSOgLWs5Y+FPTo5q0iPh
wrMuy1LIhGAYimUtXEL7Uk08NkaDf5HftlEjShyIHe24ciiuSf5rQV2JiUFc
MI1ydQxAu+/Hsjikrs14dBywqsTcZyn9Dgw8rE2cglXRFJXzXyLmw3a46AFT
0ck3kzbOflgAdx8G7H1LhZIWiSvXIeCta65AeDMPomYaxmh4wbtxKPgh+vhH
3BPYk0E9inNvGH9wsBLaj62WJ08xW+tXtQuip/cQKgCcrUBLyFUs1/iLISTz
nht2XOfGTSvBoO5LFHstr0W0tpYkfysEoUx9wJ5zGVy3El1snYi3lwo38nLD
GRrbY13BcZbAv1oEi4A5bNzk5ae4yQvK39E09IoAd75RUcXpSNbpV/iE4b86
kQRYA10gb7ByukUFiU52qxgjG0GkQlgo6PW4xibaMZuUZqClzntKrLPEu6sP
wBs0fg3kzgTHaM8wfXfe9WkYRo7LZ4VsWgsKkD4Q+FzOAWVWQCBdDH2lIcZp
7PvAVosinlUzhf6SrEi+oCh2BSzlVK+bSKp2BD8fSnzhT7nOcY+o7r0c8HOQ
81nYsb8BAniiUyqoWuUJca1pOW3tPkWgLNELWtdFnbQ2JkeOTLKz1IacLUBb
QcwCpxPgXRKV2GyRsnuvMyaf6LjgP40I2knkSxEQiNp62HEYeXX2ygT+Irbf
zIJcRfMnFKvXa28OANxymTc1IQCkTFo6kckHxy5WhvR/tocw5qcKuwvnxj1W
Aq7AhXY0AkiGbTjTYeB8NSE9WEQRL47RT32Ju+8bznOJKjes32uCue5rW7D7
7RXGyJaca/gcaVnjaEQ0WgOuEeojIpj91VN4fRYHC86BngGKedfq25OLvXKc
DFYh2b7ocSX7q4EFaF67BpeIOxYo06ajjUgm4Ne6WSDo1QlsofDYjXbSb1Df
MyIC6Own8X4mo/1IreZkFriWpUrweV4AzcjBW3+HSEjTDlN/VAMB1KZLR+pr
w74+72pbbdtoq1OGy9aTUIaiCv8wxGgZLb7zHJvco1SGopazVlGwyVR5xFax
Bl6mrASIoQIMLG+WpQkObYlmqQeZl5s3vfDg71SCiOrQBgjrzmLYTHqJMSR5
WloT4d3mbKnQ2cOVr8VTrnS9UyVkzOwCRCAVjL5u8gw2VBVoJJo/LQuWxWt6
fh20wg0SCVmZLUd0XSh2ikvQND9djYt87b80r2vR9QyUQJNW6MlZ3PbrJHmL
NOBfKiznGDkzNxs1V5ixf9tME4LIsHLuAns8QJRi5pfPvT72qh451o8LvOM4
bdQE0baC+MKOAR032orppOI0bhdyQ2hSBLtwGHvnT88RJvkuow/NzwkPsAkb
c0w6U06Hk/Ue0NW7r2K9pbrmLE3XS591dQ2+M8XBPN/TT/mFphGLn4XVJxxn
R1AmGQwk/ot8dzXnFTNmywYYnn4Z2B38rhU/2TTCo0KbkO9OxHdOEEGlq0Gv
2AIJZCrk4e6G+FZmXjyRjclvXsEdGrJ/XFl+cghJkcg3Yeosd2rlOjcL/Uga
OWSiBu80SoWz12AU4ETX1pcQShDwZLcznzk380EyYFi3sXZ9zlAjZ0fkthqH
W9Fburfir47ebwBNhE6Z4XwoW8CLsiR5S1zAz7PIALKXI31KbXSiCyoAFeLC
ommjOIyA9foRwctCGr6yeiuh71nUKvW/QF98cyrV2bgBoU5plNwXvRN/l6HG
vzzH3BjYkuNIe3p+yykaJVL6CwufSHdnmd724H5YVESIwY/FM3qB4WAzwoYM
d8+Z5RRBaMjLcjBM7KAs17BD4xiCl7uOi/ZTag26duCRkkjSZcHgSaLknrYu
V8/n2kvNH0iiqm1YyngSQVhL/6Aue1bPLvC6TJjWZdv6CS7uTlUW49+YMO3S
dHONBFqJt7lx4qa9AJ0D13RXWaLwcb68m6ihEsNaYD+C8O0heSFxfb7Ul5Ls
9CtfjRp2r8/uKrzBFTBpxiEO67Wa/vDU6i993D/4LXZghhzTKsVftHOlAwbC
C8JQY8z7U2uzM3tGiI4caA2cXWR+0kpdxHeZoX8/DZLgHD+FXsWrISt/w2m+
RrEiG5RRGP53q0vVVrRYVeDuqjm2tnQFw3Ti6KQ9ObQNtjwO0A9fvrcioGue
Z9dvOFCh70ATJg6XVkHPaA7Yl1Lki2QLA3HldShcPuf3hzRcNOct3aiGx22O
NFy3VKqmqUaOr5HhOTV791AZfAcaYqFC2aHRqK730117U3zu+//kle3esuxi
jaBYNX8876ZrI54zTi0aVU5UhIBXlYgdjx5qr1VLpQOqbzhv2m6tmZ9TIKTn
5MAAf2A/ytRhQNUnwlTZps+A19rXweNUaNxfrasHCW0hlW6TIy4qh0qDoy3T
FUuRZMy4qblPh6d/z1h/w+4sHr3XyQTOVWPUtkEfvePbcYaGYancw6wEKhPb
P+d1OoqnRHAkF86vHA7earIDo/khwm8LFLDYItFAqOs5BnpqMDPe6gaY5MtH
dYDhtlSAXsW6J/jFOw+H7H6GLjJjQEbwIXTZ30bu3SLYif0BKrBEJkI9y7pG
67eZljf4S80LTmhSEc9eyZ+txoorVNsWM5O4qjeE4gx9Jge0XC8q9y3afwhU
b28qd7nhK3d4Dcdj32nZbbZV5SB8cYOO1pEyvOkLAD3DjqCprPGHdMtzO9l3
1s4c6roiIecTTYTvAokqj58xvYE8bmW24iD3abLEWLZAib4CWElK+y8k9FWN
6/w6Z/TlyIVskW6mY73Shv1C4L7HkuNMsh2jPYlnaIscjEItHM7SXBz/p+lo
MJS47UP0vPqc3Qjb1/e76QbdUmfvTih034GC1RCQ00i6I6QP5MuYdgtYdcii
GPSVGUPpDsKHYlOE1ggyrm5EfovhmIAn1IxYMNZw0r9RmiVT6mRG3UZ40ahe
UxRVTECvAZD0Iu9Xcv8q9LSjPGzlgO7FOhWPfgPpFHi28+3AED/JR4kGZCJL
2c8HY3XLgosJO/7UnGQ9MPifW/bRB149SFmzfJ/zusmH1rKopouyBi2dbnRc
C/z1BYhO1APwAe5D6ZITi8g3c8KjJlUi+1t2tfiTSfVFjk2N93Pp7w1KnMt+
w07B05ibnsejfKLbsYFCkyal3fqgaOSSYmrLtzHqnXK43gp0OjTPg++fkGL6
zQLfDoC3zpMY+TI75tvNTbPcb4C7FzHtdbok2oh2pUF6faMvnbNSyzbPmhD4
TxhlVK8tfXhxc+spkHSZJ4BkDYSVyFk+vOvAFNNxRbtr5aBAAR9pOUFJauox
qJIjETg75iw2x+5d9ggiTjMSDR00hp5C1NJryTmK2Pw6ojqfW+jaSluEZfVB
N2vwJZgtfPsRXUIIbZvgQSJjSlPwFP0fnK6OiQ4KJnteVZGHLI1ZQdzdPzLE
HjOFtbubH6lZZdJGKMvHgt9w98y/DYRh9JTbPHji4NcLZKh6p2fiT7XxyJRG
bqQDE6Zlv30NRaTg6CgStLBNInV9u9vbxGNPbMc9xpzvNiTIaMhI4Zn8jzR1
nohxJO0cg4Ixy4icgu6LCWLLpPpWzv4r8c9VwPl3gIDd92CBM6pyVsl5D4aX
MOAIPMpY2LVwNjR6x05BG71yHTN8Em8lyNN2Iajjf0i5OLpgeO1HVcBpZiAq
qRJRVuBrd4hNuwfJ/L9yTcV0wb/+Wwhergcj36nDJX0l2UCyFH3/qc6QDLDb
RGgCW8CzOdlUvsKlIh1BG3NJiMy+EZeqhxhzFnZ9ZGcY4q3uHZsWvbT8XHxh
0l2PIdjIKRA9t9zkeg9wiXBkQopMBUm5sSb9/QwZpGSqXWR9eyRLnRrYL/G6
uTpGLFix25VI+5mWZiwvbyyOoLdmeMz2mZELL2p3o+5Ce3K96TwHvEoVRH+B
44Me+Rh1mXJuQKjSOTyeIbqEW2kFA5Gc+AI2nNUfVsQ7vq0eN2L4EsKFtiL8
iQKPKzreqwLHU11fx4Pr3dHIN6KfsFW5wZCVwaZHumOFNJN8BFLRB6A1diVy
kAnUghFjy5noZgTSb7GL+1GXXfKHhiDgH403UiVzeZrjwsPiJCamijKPpYpS
ZvCFnwo5EpeXW5Hy4PS0MKFZnpgBNWTUiCYCiMmS/FGh6egA0+ANcG1Y58ry
z3b0OQK8MF8JGHSLJsUJTgebjU7DZ06BEh+2OOQuLuHEV6hqeciRSCN3wUcZ
g1kV6R4u1A93p9goWpO3aNM6IYb8bicXcbGNZdMTq5u0kx49cjnyeEzhQ7MJ
nEkjFQ/HP+I4IHL2sXmhsn3s7sQUgIdLhT487O4bLbx4tjixlGyDHmM/Ajqn
7DziTmwt7Zehng9p3VAVC6XZkhC/fJw/335QIwq952Gz0VkPPeOrY6xf2pZa
h+AJiHuERnUUoaZupx/sqzI5AF9G8ems7AxlwHPyWmIABSSQfdt0RsJyufE8
LRdqWAAdMJwfBHzXF1RSvTJzhK3a3nYl33Nppg53k8lGZssgSouMlY/shiyh
gxndBI9uZq6ZVg5x3Rglu7cnWq84WLs2tn4h6rtE7ok8wehSKeO+8ErwnJID
mz1euU0RwRVSTMEK99PMbLrgWxN5cQ+ETQ0jM2c+09QYTiKHIxHLy1dtc7jD
HbkGZPTTqFgLPu5hjHKBoIKb0K0enQR4FQY2sbdG5Mx0eMC5hjav/bOgfQ/y
T6N/uTCCatSYVCdyqalfQonrgp6/pj5r8HcyX2DtMsHqKjjaGdOsX3/ZNhvU
Bk+rDWEwCj7L6/ZTxJtJvhqjTUmHufJGZG7WB+RFUKeztIc9+SH1qL3hteSo
tknUuFcWhDIezlAfFGo/EbrMejPnPgtIR658VSa9

`pragma protect end_protected
