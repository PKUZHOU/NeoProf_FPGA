// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
SitLNhh2NNpSkhZshWVuaagoeQGl1HOugLwlXWNfAY6xNJivhuaoApYVE8HSv2ax
z9a9BgyfQtYZf5yRBvBQR6F3Fwtw7/gUbjEzilyvSxevHO9UOaNAnSpt0HZn7S+g
InnnoiWS1iFuFHCdl9pHp2szKTdyPzAICw1rmNwq/5aSk9P/kIOXeg==
//pragma protect end_key_block
//pragma protect digest_block
8xbJ0oQJKzsF+Nx55wOnS/sBzeM=
//pragma protect end_digest_block
//pragma protect data_block
glxzIYSunAxREcVOZ1AUKzq/L57lj2L0Ihff56gczNQ2DrxBwGYB2I5vtzYnOnGk
eSn36KRSxtpxa0K5LI527VEwj7/O6Q3EV/RDBg0QZJ00g7yZf8xR9Jr6aSMoisBC
baPsgfct+au3wg5mwR1DN3x7MmGRZ/qUR0qStFr/g/RkSkkfF3uJnNGQ5E7s20GU
07XDwnIHGSNtMWnsMt+TlxBn8v6RRhseXdjTijN7FR08IW0diHzFFaDoPkFrLCH5
66CNZ3ADVYV1Z4UYtYOCBQE/AZR/qQ5gNydVpahzvdMyU3/dEa/1DXetKkLbRuiL
LR0/z/Ynuw8NB3lX5hJyBFvQ0ydMsy8tJ6rc80cxAw8tadsjAerpP7oqVL2Veoyg
N6mSVs+HSyRHGyqAgM9eBfb69fStuDr9V88rXTDGHfH98UQwvU5rg0tvnoAsqX+q
s8MKAB7VuHGxPvYXMiBwsL+4wLNaCgmrRVgC285fD5ei9GP3KSymGWNJbXmt8NKO
jtD5Cx6+hjzzgbBM5qekC6fXPATT5997FJJQJSHxG4pK3olQQGs9nCWBlxNLdpkW
uPTHLfj+1rnxOvcjzI6akbaOkwiMu/scg3X0fER6bV7O08eUfj4AEvTpJBykfTvq
9Gk030hnWXsQGbBMZiJIOdk5U37L0Wn9p5UKUmsBPy8flWUIKC/cSJNKN2LvE2RA
2gXueoOWk2KYe1BnjOaCLkLVrY9BmHXBjfyufGGSSRyETFY4wzSBKLO9pEjQsCRG
CS2gW79OQRdtGepp8wOw6eGjdzlz2WfDFzRtRF9/U63mLWPJOFpzlNIddXHQH17V
OqC0/M1u9jg80shuionA/Bpgj72mWiB+m3YWJObgN1iZcgI2keh2DV4T8AqW1cv3
878r58INBBmQoH+unePo9hGtUsKyOitHwktBgAJ7rWDlLfv1ELVS42SzAcjePk4Z
8u5jDf3Jh/A8qkUt7lVw1C5NQhDXLD/33s9nAdRl06S9+f3jPnND+hRTr2ejbCoX
hi6JbRO2gDFQfoY+GS7DIbFWeeZHft21s6RulzYczxzatZiN8ZC75T0Usn7QE0BA
BEfZ5pKm09/r8Gt/qMfc/1rTCGZRcNgVmzYYa34vN3EciiGXM1YLgkWGaQ7Zv6WC
jScm55VUP+TMKEp2E1C0ffe8ig3fSLlDPLEnpAp4qO0rowfatButPwP+Z4TC8Lpy
CHTXL5/cpBLDXZcpXEVKW06N5HEJ7uH9HSDoKn3VY/1xdLurg7rfy7OUaY6CFhYh
u+8+pgDoVWcVPlc3WHq7zuPimXV/n/UESqfnez3QVv+PiPPFcG7wOUlJe2GsNsTi
xyRwqMbox8f5nzTyNA2PG2B0Eh7JYsgABJkAzq7P6s71UENW4CJns88KFQP8IVSc
bdYU5nQ82f2jzkbWveIQJ8E5oV28AcCdi5XlJmdCzkkxJNPApisWsxr8pp0etRB4
9AxGFL6i0K8JUJcwRPi5FykXVCZCJKsBFhAXhGiRSsKIWP44JK+CmeVBNhHBAyRd
e5PjUqIHzKmJmjAZQm8KwTfsZPrgPBRXFBJ5ZdJu/nmco2dVu1g5kEtbloz1/uku
joRG526x5/asIQzVKXycH2FA8XYP4ZfZ+dc0uoYIf9GrXiwxG+X8cnxWPZ0XIP8+
5SUfSoTU4cUb87pUiKPl8GjKd09fc6abOIEPioaBbbwG3B38t2PpD2ZsPUAD3bTD
eKEtJlexOIfXgm79ppV7qo40efXR9ePb5uTLQlt00hMi5i8zQCkoC26Z1C5OqZkE
ZjSM/oi0GBzbhHfWJGZMPoH+hbY+/TPXVdtfcVKIOMNC9lPFe2crqaOjdKizCMPZ
al/LNrdZT+DoETiB5K7O7ufJ7QkKIkKaCGc2B2A0LFYHa+bkFlCtVmOcIPuxQ6Bi
Q42JgfYTw0lAg1bM1LCw2I50ii6vU9xMXUMHn2ZJIPmwWVMcit1yGhK3p67jp6IY
AGGjP8rr7aneUaqBM+oNrFRMsXOfY6Wji8DvkLZU/CQIAZjULcGDGbFU6XZ8paXB
44y4UeupUqNKwplt2EufifYSsfW3oFUCpD+56inUN0j9VweXDBw457yYGywRRzSq
4KgwzZbbL9keVNv5sgBD70oq1erDLUwAKbCxZEWaoewMQAD8sf/NIm7qMcv5+SpS
Y10N7rEQAIcxUMhk79TzalbH+ZVUgRPUwgWXPFk+eBgiEgTL7lCQsU0PycAJ/59c
VQ/RjoZsFyfyjnDtM1xxqTXg5u5OPsIjr2jojR9tHwW4xMcib8gzbhNzwJjvVucx
bnIjaPrkC5zsY4rEYK9GZyFHDFblPK5Pcvj94PrkLKrsTPkmocuhORRes48NjkFS
6Qn8v/77lsifjcSdh+Tw5qaEpLiAmxDh5Ye5Vv9IROWEGvnoOwD70cE04qFj39AO
Ae5dUgtvRE5w11wGBCV98X6FQIf7PFJepzchmpHze0OW+ndMefUnbMzSf9/4bV0c
LXrfATO22ESxtQFW+jFyinHKlszXVxkXWbzk0JjnH2LWbhEHAhXeW4e2lh0lwUrH
Ms6n13+tCThrm33RSU0mEJuq31tbfdDX1wJ3Y45usYirzAVt4Iq8uncTzoCjoiPW
M2H0/PloV++HjNieo/tpDwDuba/R4Zdand5Rar3mTtb/xq+iNbhwC5mw1MUTu4Oi
3y2NHghQbpWDp4rtAiSTfDJwY2uPiC9N6f8V1J6Ctxnwggk2OgXJEE4X1eRJmx9+
2yd2cs0eIqzMethodfgt/e9j+3vkJUlah1xZrSbg/sNJQXWBj6C0/qkm+C2mGXgD
Eyc+Gu48w5PeAw95eHQKUdP+RsaMWniQdp40aeQHzYahw5HVORc1kOs+NnM+lfqU
GRmY0T/FHYBeAujanwMNvBJUQ4Bk3kBwPDRe+N8skN1qshbcM5yap16UkxwB4WKO
tR9KXuISp7GOeGTDGi9AuEppcUWnUql97L5Z20E4FVfOh4Oj554JKqSFhHyx00/E
oM5+vzSmEbXql3O6k8RKPevg9ZKr16cFwmskDu0uf49imVCQ1EghnHXcGhHnQn/N
PvIFrcsx14v8ZR8pmIrXTfPvVZrnB0f8zrpM2NQFmzIWCxIJNzYk7OvCcg1qyvwe
u+sQpN1jdbWol3RbgFHTRzsukUj9U5EHofBbn9CEutAyvzjWZ/cX1eHuJqZoeXVt
gi+qkIzhY/wMwBs3Fgs2SKyFZJlZXURD2BuhCYAA1c03Dah2GUNtLyI7FxfyRxy2
OcYWtrfN8EE/yhodyDUII2jwuDqil8PSlJKOyjReVnnbPtom3BCq9r0JaSfGjNAb
W8XgXtxi9T+p4jhDEqBlpj8mgcnI/5Ol5Jg2/nYK8j7wTeywZB7zToLvfNqg/Btp
tmujgPSRQy23t+zfG9HX3MU+qyzhZyM85QQeTWkYUvJf5jHqkbz3s8n5DYbHjzTU
fn/CjLHEQD99EJ6jETxgR3A9m1zFRrYr1xgEg65BKO+xbAaqaRhaqTppdnMgOvhF
E06EvR28hn2XENmI6x0THlKzlt4YdK32oI9uGcp542YPvVvIx2u7YYs6t6aJRaIW
rou1VC9qEDfx4u6KLwkhQ7/vOj/Qv2IHkN/SUJ9UY81w8deBpI3l0muPY04pBoXu
Ip6OlEiKc+VJnsTy6n7XJ3MDLGAnG3UMrrqsyZcfN8en2Giffmv47EHz87G5RAON
6FWwZuOeS2Us9UcTWLbAEs6t3mfrfVpYlksahiCxTyAj32tyj/Ki5E7iC1/8k1zy
6wA80tdoD3mLlB0NuTas7ZS0z7FRIQusvUWxNeKrjfTIEcTMPHVSdKARqpOY06qk
psM/is9iRcmArM410Hdx+jukUErV16LEoIbzACRRzcMt8KtzUE5nzydob44akyPU
3LX1kSgeh/+U16T6hdTg+1w+UN3117QSadzdXNhxwTSSaiUTk89spGl99UJRXskz
cLVj0y5EfH3SoxseXhGimd9Kg2jT1LT7dseVVzNpMoT4Rt1RIa601iVp5SWeUbpP
RgTM5V0+OLZjqhOwGMIhrENfcIIKVcczfETujtD2eNvOukedyEPt0DwCl6WZKXO7
xUg829soWl/RBu/lcozgeLujhMbdtD6MiPuL8VZMnA7Oqh+aEP9t96+iBFCGvKKm
g0iiR5xKees/B9wXaYanISVd0n1OuaSs0SS7e8RDQIWownbZNofOMOQno7dN1SL2
m8GYTh3LP1D/Oq9JCCvvoMLsCU8jxBuOd4Jzao2oldgFOTHM0TgqkdYOZqAQ5yN9
wSKHXSYOJM8tGyQ5sJE5nMVxDyR3c7FdC8QEHH6IGf1nIuPZhXeV3TSGDeXPlfEp
m0ZQwq/X8pj3SDjT1GewhvApn5FxSDJw9/PHW1IcF4jn1vbOutf+XX6YnNKfDF7Z
6FK84vj03whUSGVaDiUYpYwS5RjS6nd/RgQ+eDTC6XzrExoBwMAopPn9oCQIaz9m
X1gl0QN0tEq8Du7166JeFjZS7TlwN7P3W7tgT4B1izft3z6/r3JNL9NWlAuOiw1E
kJfSNaK9TV2bmrMiC7ln6BNDRBkcgu5LxRXqCc2o7/5e7O66EsMdmY2j67iFcWlu
0ArcNEO4ibGhtG40Rv3q+4j59Y0DMdNWB47u7AgBbbXUd6dq6T1aI+ahVMbaUy3G
3KWTRypPBo+fGJZJammhO74EJgXPT0NpTUYCV3G53wSGnUfNy03BihaWOa2u2IZH
7lVhXXmMid19UyjKnyUCKJVhDFSgz1ieO37lDvOsImfKU+HPtMoGXkHoYnwSInwm
iHwhzO1a91rZLg4wserx+R+uAnFy4m9dhOA3jaO/UFGMTmaMVP2zajpX++NuWUyM
eyUjri7mOgnSgqqFYsecP4Z4RZc7kkK/VaklyekRFYPoT1d8cAIP6HBpJG5uynMj
XqtIIJmI5gJbxE6nvkk1+OIjDwiWuRHiZl7yszoXMFUX3+Hajn0cEugO/yos0+4q
3H4EbvS/2N/+KS80bR9ydJblEQpQwHmjc3Xl3wvZFFGDtNB56vCDONqPBxhOPSKa
xne9zqmaBk6DFdXMEFRZHhiBtTeTcrcdtBp1OvI1CMK8fJ8ExbK1PDh2pcbjhb/D
ztid11S9Nk361Y1oUrQYe+a3+mBMlJqCWr0n1ueigBOT3/CX4GG8WVZYvqPYo5MJ
duR8KSb2a9zF44IbAcj/+5bYJVGQZskf32HojQUxIaaaUH1ip5gK6xzbHmIa16nG
9AHVuneFJvRpA5ZGlK1Wx1Qv5zSAeykf7THZmfRVTbo/s04TZXKurY8EQyGgSLIu
p9TWR1WmbaM2TBozSDltB2rVvHrp2xM+kmQlTvGT6dbLpssgkEwr3P3ja9KBA9qQ
Y2veMTgM9JmuYHWgbtd/7kNB+xMkpa9zSsZACHLyIHdWRwB5huoKTEvmtsUA4C91
3/GpuALOnqHp8oA8yeEKdAMNCP9InNRI3Ru1zICemK9F0NCsLdTSj600y4HMkyBh
7FcirxSPU1v0m6L6XK0azY+gDw94br7Bjsprhv/3K8X0zDFzyFUQf5bdewg512g5
PDxzYHBvzhJv05vhsTcO3OvVajltI8UWPEfJjDT8DPQ7xTOcASr1kE+oJr7L5A8+
yz/CKPFOiPGoCmEw/mRnUe+QGU1s14vufynj03VdA3+iIWF1msw0f4XoJZRkZPvR
GTF1tTkd6FASGk0PIF1la9UUj46Urf2goAPK3OILiIVXA9UNZWWJgdmiDa5Zoo5m
fc0CFzPUEPrUqcqJHYsjFDjcWK7LIjPJcoPW9OFjLJpKz1FSaVx3O84tPQcDTAlR
d/6OmPVdnLqyvuDruu1rmo4pj4f02ziDYhl+64LodtzXE2u8xcA4rcCsFjU+soOQ
sVfMMSBnEOOyhgJgYoULi8yOL9WK5NMhEVSn8tKqj1SdV9qpXssQwVJYGmpUXUQl
JdegX2J/NbUHmiMQaALWXo4T3GUSjLrimGAN1heCmJQdnQwKzrJgKequu/a3R281
KJ5FnDXpXr/HSRWVyRpkzYw755IyTKGS637uRWcQVhKw6YIgYNN5zOxeLHq2aP5h
JXIbpLO7sT7PEHv3RjND/Jjl+rQm1tVuiPFJeW3KDq6EyerSbGnP2Ghe3nXvAcMp
e1b4jrFFsZQkpyp5q6tMbqm0om4TrRcLsE4mmlOAZW/Uu+AGwxcfT8EgjxyMYjUH
0UdD34lfcozfcqY2fbF5HRy9Vya3ppIzbkploFYg/0NYLkog4dNn88o9dPmpQPKL
Dv2TqScByeiVMsrk65RHD0gN0E0Eu8Ekvwn+ZMIXVXSEcYtr7gIcbuW6dCKjVZKf
CyhS9JCW1RzTXr++S3/0One77PyGwnlUsmfOs2xpr7c6xauzNNrxowqWX/6rL74q
rj7fL+Anwj8k1t3KMh+BzvsIk139dJ/knTgdKnR6C7j3qzKX4qqGpQGG2UlMUBv9
SsO88AlzgShOQGrebSabbfatnNs1SAebdFKONSZO1vaQeTMaU6xIflVLiswdKswz
N5ACthzyFefkq9q/aQbNTkAHWcpaJuUNnsPuqMSDunA4sJAK0oy0PncFrH9U51xl
Qg4xJ4wlD5mJP6KTdtikSHVQXsYmmnTncL1fOg6M4h9tPyKKcbl3//ALOkC0Ozye
u+jadhByMphx7gINk/8xvn3XHbuuwX2LX88+yJcgXZki4yIKJSYaVlLdqSJ8QgXW
FP4NRqPmmkvt9wYBWkPNIT/W3ZtiJFeUVVwXPHXvcr+cvoaeZdXsLT007GeOf9AT
CSP8dvSXjuHibZfQtXM+kpGHhxFts4E77k1yJd+go/dvmZSg8oYEiQdcv/KEzG0l
0Qajck4J0Emrl8CibDviRy6+GRbg4T8iruvFnupj+ZA99e1PwysLONXiuldYS4jv
sKWU4q7s6UJK1wncg1vs3FhtBJLgX2UDhRjHq02Pr5N3fRjqymuAItxsLraQVYN6
uy4eHh1nvN8F4pms0qSbZDoyy4oroC0AFGxaD/ZM3o0E5NWI3tfk2psxE5CHO5PD
j9z81zgKysnRaAj2m2Kgk4z6yVkzB/NkK5UFDckCUBNESGDKzVk+JDsnWYlrQznb
qhAYBR1mmEba6V5eWYW3B48FDoznZz9+1Dzn/jAp7ePe51vVKaypgtpGr1tIhu8c
htgZj/Mvbo8np5i8g4yi3zZlhf1pBXp03Ri6RnBSfc8lbce1nguT40RT00TKealU
lVee3zYValO9i0GDrrcnLF0w9RSKQxGE5v2LSqLhaQyhFMzBSyV8YN8KqTJAOSjt
CQGSFYfT4vBaflT9Os65VfrICD0OzHNOGYZviLHLP4U2y6IEYPK3sye9yIO0kXLX
izetW9Y+EF0kWy93KtRdrgm4MmSrmlCXJqZuV6e7q1gBf9E+RiCX/NTuju6S/EGd
FBiv1r65JHmfdFpHKYby6nTxLpMa30wpZ1tMbY/2sWMdgAOK7/3HuVxqmhnlqn2Z
EMXK5Kzj26c3zo4nLLTDVhqP4xrtiI7CF7of/3VQSQrV+2smUUAyupdNHSg5TruV
y0WSxNLBUQEop0i7BHza+POPG0AP0FKvZQsyaLammUMHEykeQJtwlN9t/7yI8R0O
pOYuLXDlJdmswsVS6M/HPRFEZmnHMYf80qUmu9SalmKuGpYVkg7zf1m/PNlwsZy/
/vigZDekLSURgJBNCFVp6GDaMsUQWGiajx8jzcPGEoiXeKamFD06VFwdPLz+uQ54
KFal+FKtH7bpgrShHicUfgcLMyAyrZONsC/b6S1SwIIba5uvcS3g+OGnApMdfaCa
mUQTtubQc1SZ6jTb21Xm+VlRaIlqCo6PzNXZyqq8F7LPUiQ68vTjZ8GKLX7wwrIo
FtoF8KzJ9tEqcf2+SE7Z9gR8xb5F4MJzrbHkQMSnW8ty6yFC/u+1KlxClI4ta+ZL
ByFxY6XlfB7LaLUef9E9CCAvsHHc5368ToH+TaG6OOrrDl5luLf4caxYg+7JeuTU
urvpTyC0CYgFsna0BrDXjY0SkE8Sd5JnQt7Zbbc3LF6DrK0tnoTovjufQD5MhCV0
NOi5T0C1sD07ufOeShAJJL1Ag7WTILbRjQmY8YFmMyB+eQTnOjXGqNniqlFKaLh0
FCsSgNmhtkaQBjBe6o70MKtWyFUFrC69SuDx9Xqi+WtPCvrKZxYy0Xh+qkBnncbw
ggjG5JHIZW/eII7a+VKVMIWNIyps2sn9kllrEU/Uxj5KoSB67NgyaQTqfJXF8c+l
CMysDA3TfwlnhAPtD+wo6lLBqtH/+M0cStsMLtGGIHmglycJWr585C47mvVMrX04
T/uAipg+1tllUU/rGDeyJ3J9W4tm659Jn3PxD8JVx4yfjnu1uR1+6zMhuyVudVXy
nINS53WWrHhTfwqUEX+hc0ipLc7RhsbXAUzSSCYbUfYkttQn903Di4BE7vyVG/OB
pv/rACFHB2I06BOh6OP0f6h3bUq+yM/lgHVcn5PO6D7EqFRAr/iiKdw5DLcbAeFp
32k7HKsWUo2wpsEYdkHTxPqe0dS+LDHGfZcNV3upWxHG9Fdtbm+/ulVNxzaR0QIc
vMquCI1n5TGjFxAO6GHHqHdhvBv+YUahNmKEiB1wvRtA3saiksEj3c00KgYpTcw+
Kuubcsg6F8qe0NuN0q81O5UGpBF5DZA8PKmAW9wfhuh7bsmKiG1PICHnCekJIY68
KSEGPSvkn4m4HaLqyU5u6zOG1exT+0MRXLMzLz5Wg2Sdoq4by0viZAF1fn5R+W1a
iOnakFmYUDW30AaIJe2PBtFeOGQ3KzPDFE9EKj3lijjCElJzgwONRmZRbK5RC4xR
3s1pCHWN4moAQGgXjgQ/k2kkM3Xbom7rPmtxDUrrdhMmZLuLVQMxhzHPzwexWoVp
fy8uoOEpTyVYTSB1CxXz3aYW9JlmswmpeVtzMLmOLfX5rU3Bgovyk7vPKEVPuPTN
AAKPdUCscAbUKHEA9faFGqRURGlK2XSMeB7p7B/CVaNudo1hQRDQv/HfcCz5cn2F
JCHJc7LuUDwP3CI3efdb6pLX4p2W5MhuntG/xQhL3zLdky+rnU8xV8HjE+A+OZMQ
Tnf2dKPZehyF55kVd+bFei8euNgVQeaQsVGhFJBFe0uLO6RdqJMBQeGCiyX5QkMn
bNcV75I1sWSW6lczXO1zq8Q2k9yOFFw7Hz4sIvABn+vA7FMeRoFoPDcI+gAsDVQb
F8nWxXABfmnLeC9+HMgHg+JExtTJ0JmyUXmOt9po7WsYC7vHGfuJiUAQ/rLWBPp+
hX8d+gnNcs93Kp7/gqxMeQBOyV6gCglnODWm+7xCzhgRVjBAndmQf+XBL7M4sh13
q3LUDBF7Tf2igPUvB3VJ9jINsprH64ooRR6cMuV7oilAk5HHvVBr3VEoF+KliwUF
lfsCtSXG9SyxpQbnVYSlviJma3DCX83bt6APj30k/kAwPsR2o9ZMeLSwWyS8TY0U
JL9BrceD6V1Dwag8lKBuldJnORkvZPDI69/ovqUZQXapC8bTPy3ulgNVROsBJFE4
KlwnMExlrlLxtmYkktV0NQ73KEByzAIvSx22qiCAHeJZWprNAZdmgl1ffgRtmJrJ
qRDpssrx4u1auUfZgmNCLiZOrNLVEumGK+UVNz4QNJ4hUZXPhW3h4uHyobnIVEc4
lQvH4QWflqLx4dBIeuAOK2qJXzFxpyGPjVIqYYd2PP3uIOTBJLFBylSq4MKZ/Uc2
Fj9/8YPcsWvUvrhouq6rUutmRbyL4Nbx9QQsukQI0u/jtPCAJ5YiiGH0WTAF9xri
+5YaoDwbqXJTHQZzhLI0SA7oScIJzNxR/+FwjTJZIMpVQBjD8zQjgPzwaNVKm0kO
U8Y0HPfI0QT9BQII2vME9qZUjqrXO7OWo6iM77tpeTKncWKsk6gS/mprElFJbDP9
rsXUXXyGY7DEKPpnsmin08zk4Dkk6ZGdVT90xsKUoX5GqpYU6Jlx11U5qLOO1HK+
3WYqopofkZp2j8gvRhU2dh9wHZN+RxRn7w2Ge87JELhHy5hw6ZudKeK2ZXhmSsPi
SxxEPi90XFMf0AnkgaehS6MycTMcSM220UZlDRx97hVH0jcjGkRhk9mFGIibEPay
iU1Q00KLLAhIntfWbVBakUseS/vPUpeccNGZ/viE2VDsPv3fp335734Y/voI5IHE
uhNRpz0REZWP4YX5Wr1/F3PbwaFKrcpMFJuVwVsoabk78cQaImCCFayI9nVwXHPg
6vm8C06UfiqquK0zAO20Rn+RmQrXxuOC3ya87PmvXlL9krPuNLQ0Hy/9WvI6TViD
/4lUz4afa0HAMNSY7/t0qSDKPuAwysNJ/NiUJKYFDQb9iEHU8zagLDpZa7SbOfEn
o3oYbB0yE0yw8UiniIHyXq583f/wy/q5EuTMPLEzAE/M8M/YcTP5vC6mPxP7sXVA
Zhi9dwU0JcyaDML7eezFJ/w1nAM9MiKdT22H8k9tETD5jApcg16ChRrPaDHCkhlw
esyqMIzvO2zpJswFH1p0fbDEUvnI7QiZ3CxlHYEuSaPDpXk5aJRHXD8r9YHyDlRN
GVY9SJxTmXb5pgu0dnN6gpBO2YOvra/pnQXX5NkWFRT/DmD+GuYibZuBHLPnBZxd
r9kLt2o6opKtPFNXpPrz1cJuzDfhj8ptyYWx1tNVyO6KP4mf+atcjgpk7ocSatfp
8gLexq+A9xvvLug6F9vwrOcDgXZZa7Bl7Fo9XxZZHSZhW5nMCWSsvP2cusSAj0tr
qLpqwlUtTADwTEWI4+Inv1oh9+IjdjhfKBAhtLwtq1Xx8ZnHeOheFEPwN7nE2IRP
bEXGptn/bDIZsxtrBfgIi+Ap65WN9HHGEQKkuKO7ScIOFbZyEMCaZgFKrHA+M/0i
4tClmSeZ/3a+g2sjmFkvzSV8LabKwRUQP+rP7Kz61AjLMkIx2CBtaYsmYVOtysa/
m81j/S4vfi/AfU0gwP75b8o1PRSG55YTyvkOU62A2YxTziFL6j2TWX2MEVOHCMiD
15itIdYfOYk1WpZgvGVk3KzWXTEX6NIdaeSDqgaCr6d72853evyggp12hgPDXfh1
bGBeIUnBDIbtgFa6/uIPOenNwnO9Xzwxx44Fr80OQD2hwQ2yHS3wLUTwnOBwFxDe
Z3OP3zxL+TSrWlVezMn9FqOJcHTecv27uEkemT0/4YW01ehpCk3K0TE7XekaSP/b
JvTrSGpDg9JKH5dJ/Q5ARSgqNoIXZ3hXYTB1Ewnlld/FeGcrotzmR1gaGdjk5lUA
yBA1hwsKOpQiwpY8D8VrwZ6ejAMkfAHNEXonQLDqzbgJEr/Ti0ouTTO1PESB6qMC
mCsUmjH1/H0uEDzZdDN/AQ8tBNquDpOFYPDdN8NGta6fkBdkbg3JNt1G6jMhADAl
Mr/zkH8XB3RvyY7fn0Y/UvAZp7CXAoRwo+/tk0Ult9pSkqlFJuPIGCnXItvIVLXu
TJ8D4dae3gDh4l0OfkEptVaAOn45gIInFmRmFye5o7lOE3kGHzFwwz4SMYz3UBkH
yP2597F1MnWcdaGAXxs3tw3bGoe9vORa1Ds0Ruf8d6mJi/tPxkRJU3ghyRv0dAm5
ShmUwYWBuyHk4BXO3eRlOS6rTPFP++HU2dBoZ/WyGCJfABwuzRx3mIXqEk3/m36v

//pragma protect end_data_block
//pragma protect digest_block
ynnU6ERFbCnn763r+atFKPGtJCs=
//pragma protect end_digest_block
//pragma protect end_protected
