// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
1+NEYc11YNNVRwC/8riDGerWb2vogazjhp8TTF5SFtDJr4ItK7EAXWBoOy1X
t3/uzlfFFY5yteqt2Y1/km/XR7VIkv8IjIrbOJbTfVUCdERlkhxgKwjQ6Fvq
n0XnENkqUMEjLAorz6+94/tUz+K5sLXShQ3nIOhZenLr8u9DGDcVDW9hlw4y
KxIw/oaD/DW8bVzsy/+PnrG4vAVQ0tjJy74xgzovwknEh8k+NsQCta61tfb+
IwNU5Fsf2QPp3S/EqpBcnkHiERQCxKLGPoIZ+kWHAAFUXtQ+CwhacrVtzA2D
zv1fUrFQSvFvfPF/0Vncv7/YmWT+Na7qwZBL9QqFzA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
DvdvLYbTjv3h9ZCw26XDVhaBrmHYj9z/P4FcBpY0HmISUPDMVJUaV7Hn67Vz
iJttL2KtfFwzgVzsrPZARLxqW2qam/Op1ddqnayozshow2kEklqHAS9F8T6H
6UgjGUudNLBXcJMW5llGpMfiUumr0nVhucicpUhlZMDTNhsOhPMaXRBo7ZlI
luBFUm2V3DtTY1qR2J40m1Ujvk0WPM/IygxAa5z39ol0HN0ObKG/mskdET+7
VhowFqcgHcjD7rKef8Sx4Bhqx9nDZe7JtiW+/Ki+2tPpnAWbeTkOocA3UR/M
TRVVGdcfwqb+OIhG2zabGLef1nj8lNf7W45wIqD0Xw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
B6OwGpKfTpUqDZcNmQRg8+mqNvbSzRAQrearvnklWYHyVHDO5ImokFOvtIEl
avoxjir8Sawn+IVlHw9R7QAIl+o5gawhQflS4osWeFJG4b2MT+LIKc24Sgsj
tNkxkofAvP2AqRAU2WPMkHp88PTUfo0L9YfLmcdi3EH8/EcBIUc/bjS0bg9T
zCGHZzqOBfkDidTIKmD/i0AGd5LIIqla5R2EdavTcu1Rm92+Fsl5RlEn10uH
hOFB5If3zFjJx5TsR0GhU9TySOH1spqbLD1LniO5YInVLjz4oed3Qz2bQ1DR
aYGDsxBcJsA6OKldtsz91GecrN3xoxrDCP1U9v6JNg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
kykh04YgxgP+0vfyaAZi0zqqOoLOBiEKEerIjs89UnuyKn+WSEaNkCNPMu1m
a5OxHaYDTQ43Wi/CsDYirqdBX1Em/ZlJGUdKx7mcEF0Ej8rZ8ZjYu/KNfn86
6bhX57OLQiw5IPikS8igif0GPXrgtuanvBfSxyo7PlCXn9urncU=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
M8C9sjBUnX+KbVTKp+SPyUXnVQhvw+8ofsGr9Us+1yVTLXpHTPulNE0ZV/Ot
5kHya3ycTDt5fCFj6uNQ4AHthJiZNPGWn+zpKFJX++vydMRVOpKn6Q8n5ELh
JJSS1ejV1a99zN7cn046Bk2Mjkb65lghGdWdMohGX0on4IkQbuQDZEWGPY3R
39eP2PNiwJKbjHqEvKFVRMinRjad6PDW3TMBlIxWGfOMt28rnDOU5A8Pqff9
lMvmkpp7BfJjzH79nMxnbvq4yFRXKAOtdIatYUnxJafbGwJmygqSvx2jaXN8
JICzO5tAC06nW4KskSXk8zG4sPOwVK8AKslv3QBxZOWCvqB7bSNC9PjcWa6A
VFMYbiXL3Z4GmeOjPIJBqsmmtD0Qy6g09+n+50445pbu4VoYAiRcrfzfkII8
fmrS6lMIFiyOBDCRrHXzsMFHI1H4G5sqvlFMdVN1zkJqCg1cWp+Zi1k00ZHN
LMTdQMex+nkcxlXx/6Oy0jUCKNjz+bwR


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
HR0UsOs4jBpfSUoMVDR3FGL+D3aBfVkj8u3YUkhSE2Nmtz3eXk/B2/vOvMdK
birwyLlCalrgV9daZfrvUhZ6VbNbFLaUr8R9DkPFIv/2BBDNM0BSrrMRl8L5
As287WK9ZJaaImibtqgWte8ODHVazXmSlR28+bKcJ0yDWYhnjKc=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
cwGT3CDNGPXh3Usiaq9UsJczVjmL6SeCxF0nEKCUaWB4XLoPSRgJ9UZF34cS
eJun6EM1FlNxIiEV5y13UX5AQEgJjzcvumRWSgz1nsD3CHKgcqz+DFeR3yhB
WlbuOrdcTrsnAlVb9JSfH7Q9jghZ+vyTHP+snpHMwpBeV2jai+c=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 65472)
`pragma protect data_block
ZbarRnuCzPjSfzhOXIajeBC+ocAWKmkDbofy2CA4W+EFmQg15y+bKz1PQHN+
YLOICFhgw1l1QED+IbtO4co0uk1qgaiifvoOLAyHAPURM/UQWR57jXZnXRAE
arXHjdPNL/D4pldXiWrVtTrVi0SXPNcQTEiTpxUAJzmn0OuPj1wpNakyaTfs
EmjRp+qBzKyyPODkrOfINvd+a2lhmJ+2Oxsfjory9xjF7TVEe073Dg4egpCD
EyHazvxiTUrb4/DDUowIkTuugDiFwqfvs/Akd9h0PCJFzKNjRcLgHYABbbzK
H9uS/pn/QmyruI444mw6eheI26midKKwl7iSXM72Yry10rmuQk3jca1CDEUB
Xj94QYtnfcyKpWnvLhqgzYEDm8Ppqys5f1ox98j677cY9fLM9urwGRzbccjg
RKVc4oIT1UGLqx0bSWIzBxc1wIKDTqoUNlbcDG4NnHuH3L6IjZoHIC3ohIdk
14gNiv9vlz1FE2v8YGF9HYlGzAv5WgT13r4qaDj4HHXpYOpdBLgIp365iSfN
wQxYLVUKL5jEDSU3BEF37w/Z+dBiLpI5CzdBNAipjNoQyOEEc44qSwSYPUdf
Xu/ZVfUGrGYSS1ULN51XX/7muYlEv7ysQdsrtRCm4RdJyEh2BYUkx6040sSg
XY4SrsFFMUtAhvyQv1lyaZu+v4lxlDdDIV+dJeSlgR6GFva2IuC8LVsVQEsG
WN7tSLFGO+BjqL9N/MvFRPOD8edo6sAkUIA5wAApIQzNXvbYa6L+3nqWx45z
foz7QVIfnHKUriLTBdJ9HUiTO2+APQywA/zVErxtoB03WH57gT1ReW2C95Am
3E4VVCZQH1pChFOh8D5nyMjSyjU63PX39qQd/Eb9qTNuVUe7N2HTp+sSqBXy
/BrsZG7/F/JrmOXaHL63/6t9qKmVMeQkRF+C52R58p/tUAbsFWaP7iwy2zqe
gAEWzWSxAvQypwu6hVwg9Oq7TwJR+KaYWA/cMwRbY1U4N4TdUs4niV8xDnTQ
26c2SzCSrlo6KNuJ3tdOpBS75/bSEt13JZ56HU7hw5tu1gkChgDRjtd2dnWG
h5q2wUOZ25+F0cI7WGlhL0K6dhg4uO5lDd82NdfJG0LvFW6nQUBgotV5zyPJ
YmEYIbTZp5sOLf6tIT9bwCf2ciDRkNNQItspwxKHJKabam4Dmd3mn4ZaPNo6
sfsEzDbx1FXLdbzrvkr9TP3dQcUPSuI1gd6ocJFy9Hk/cS3fVRP9HSMpx6LO
DMOjLuey7s6nD0bT/X4rcVNlAGb6Iu7XrWzF+KyYSOT54XKtOJuOBDY52eBN
na8ZJPiLHxqe5wNfip3dqKFmqbBMUY/67LjWv00jFuOhzTQ+vCE6N0bTi5E7
52JNXCqYUJQBZjd/RyecMytoDUZgcDwlAxJRkGMyiG23dg2c+NAY9CWAh8b+
JG+kWlghAUIN7a4Jnj9STuSOW8sAMyjz/IOv4FbF+zWM4d8Xs9i+ua1cd2aL
Cs/lzuUo7amPGIVUQ5+rOB8vdzvKb/wsKk+yx+c23xyr9Lj45fDl26SFn5hE
Uad0NSt0sqwHXUlJ91ER8+g86wZwr8LK/bsJxwSxLLBNYBqRra5ZXMXc/MuM
NclYXkpXaLEtkZs3yFIFkqQlHBVBO/cgNHgeRkq7FYiR8+p7BD2c8s3r+TMx
r4bXFOf9O8jZbqHt/KDh39JRXe4ezqavF/96ZCVxA3udsxcbEEaqoaJseyeq
bfIkpw9MHqwlX/WXBuQNZB2XSIYH1YHdmoBygp64pQA2KAZpsyVRZjtCC9nx
T/yJB3haV0/mxziB2UqV8J1LJTKd/twK3ke1BxusPvLSic0XCO6vgaRbIfp8
3Y0oN2JwSC7QgK2uAkhVJCC3VybxIhvDc9K8x2I7jgAdpGVZNTDtiTgpetrx
6G1k115Ke8tFig2Y1NGSi8Ry/1/B/hPtWiiQTqvEPwzb9Gfv8XU+Pg0Unms2
Zu+CNcSAxm2C+TdnhzDHn5lJMMQJc1nRqDXyJgdXD0uyhbtn0m52Qo496+Qm
4zjKKReJS9+tWEEsWQcS0rFFCw+OBio2uKe0y591knu1dF0zIvEsyU+s3qpT
Q/gDyHsb704w5MRbCFVlzAYfU6VbaDBGKKes9gFS+0r9gZvpR61B0w7F8NXv
KAlx6peOm7cm1XVK58+eYP0inPNGIV98HxYH267h8gw0Bn2Qud52yvQ29DCw
56x4h/cOzPwyzYfS1rPWIuTZWMQxUvNmb5KkZYSZG+hX2FxA8Yl8AJ6HkPYP
ASus7f0kFSxmbhd78RkPi7xC68B5A2HvibLrUDBr0zKHWbADQXN9oh6vkNUF
OgnU1CyKn5EdZFdAb6CxL8rUDyuE4p+wQrAcTSdncWeQQQeDRKIYgqgstmu4
jKf0uSqKH/IJ1vxBoZsSrQiU0AJrD6llnJkpLHlzTWu77lvChmLu8F1nVx2U
DhOlW+mm/1TKzZmF8nJrf71DnJSr6T68pri3ztck6X0BZrqSF9PqRVDMy9tw
aiLiClD5bw10ILNkEXm3tR83oE5ZnzvVnFKVkZXP+YZ+d6ek5RKXjaWzktsc
KWkCQPNQ8fVfImtgR0Fv9n7IC1ooeEjM90BzREnSuDih6ChQrflhErsyqN6O
gxBwSnm0UCwl2CEwPk0/Nu7qi5PqUpjp0IC5OLTNfad4jllL6sZdpaErScXA
3Az+zPuIF2FmD6c2oJq3dkrGeE9OVmbyveNDIdVa51j1fMpTaWrJlajKqMsX
QpW7tjVwjhuF/p/96am4AgcOlyAt/bVWPWg20A4sp4t4c1+zjs/TzCXzl1zT
0s2MKEtz162s0kOmg/p2epcpJ/VSPV+VVj7Gay7Da3p3/PIv7jFTcfxuFHDy
8A8NdDBISp3xPQIXq2QY0N8nTyQ+tNiTemyxmT5AhooqrNUdOftxykUakb+X
kU8ai96aPsvEx1riH8eXXYVOG0ac9uFra3ZFN5fWHgp/uUxpUINl2vJvKkVp
5zC1wWSlxROZjkQER+AEKTySXUv2svJOoUFED+aQXCGWb+5jNSan/wzXpcw7
DAJpoIQe+4sec3AAvZETCz/k+XBDai1+41bqTt36VPhtbiS4hYm1xbY70308
fDFDeDddNO/TsFXvaDXBZ2rJN/awOFWiRYpWpxdt/w6vWef9g7b4LveFFeYC
MRSfqpvwV6P60FgvJKZpMinUNMYZNfUUm/3SFeyQlsxQ39sApUCSAtCHYoGj
2U3iU+89AhxkO9f32GgkbuaHNla0lvKcPAOsbmN1qHv3ss0pxtzD03i+1Yfq
WVMnejD7EMMURp/cn3ns5bnDNw0TiELPiCx7lRPtvMBin4Jv7EopdYQ5bsom
lZnzBVJnpEQEloN6wjKi8AqGfFesjO+5ZuK3jQLe91CI86U4PHfpYahzbPVp
zthZbavMK1FRJ2I39QrDvWQ4vbZt10utsxG5rS6zHeHNrqLpswmYZq7jVL+H
d511Qjf6VpNLTev3w+owbQcOlqYDmZp8GY+EILyWa04r0HVmwFSNjpUZWDYC
58vY8fYWCXqRRTbMezdxa8DenqJ1iU1+FPmlLnZx//dMSNllQV0oimy1TDI3
yXQmZkcPccq4iI+mi1PT4RNNHdDuzXJis+S+I9Dr/L0pwe33IiHb+/rENOkK
dARU2DyImwSTidj1GVx2KwrVSiAHiS+HRUy5Oe78Z0yDlz7uc+IQNKDpCah3
yriFFgQ6V+Vhpclbt3KhonNVpYu1SBbLSL8y8ZYqhq/M1xsdRIKhI1axp2nl
zWFKcTbzZ1DO2rDY8TwHYIghuBj1x9WJ9THvQL7T4CUUcgZp+lrUjQ0mtUUn
6zSvpU127nxVTDwX33/idFANBS8d5uGo0JQOjwVkJD90UgokNQU+w5+pgHGo
FndhwTHtErEK3UA21dvWZA5YySAar1T/jO1nCKPL9Yr41gJeVPj/EM9EQi+s
LjmcaYXJ46N0DfmQ1LMXu51zR59+QG6O0gyenR8ZP8Tz2FUvN6F/HDfr0mDX
92BPYVfQp65wfLG887+RH9chqiHNXdxFr9tLUy0NShnSlyQsMGorFXkDXa9d
f9WxZDOZz8bH/v22kz5fyW1sBOiHgrKBXi1qF31/jTFAeL+peumpekWGaWFE
/JbPULIPJvFksOQ78DGU1Xw+d50DMX8m0fgSxigUUi9Bs5njxAM8YG6QW+pJ
z/UczSbzkhofG1djasm+4X1AXF6LDvQ9gggrsKCrWgFM3JHaG4DFjsrtpxwK
tf991X3/J2WY1ChrBuOGzEB8VBv+4ioxp9UI34m0D1XPxiRaMl9Tak5YO8F3
Tzy1iCjWZRf/Jz9twFMlZPpqsS7QnG8AUsCCt994ISgnIVza1CfMhsAhlvHe
eXnt2Btc3soy7AiqUi279jiDoHvjG3/U8nGWE9zQ9d73XJwi6Y6W3GpF9mBa
IAOEcqYg9qYe+D9C2br9p8hUu5D1Xs037Xq3/CzUCk3SBbS7kqkb1g4CSQ8y
Qni0DS6/CV2cC+wdJMi5am/gQYz+vjKRxp5jRMgUXGPvWx0DUtJe7FTCMtrz
WVD+Vqi2wHXVllQwyuClKo88bgCHnlWoKongmv62y8Qb9Vj7uK9ViEVyvyQt
VHG5aJeivZlgA2wrHInwn2TUyONB7Xlu9BVoXGgexTPI8nLkkWruzsMSHoMx
g5MWd8Am+i1/adysU6Bz2fWt+6mK1pgrWPLohyLvbrN4ew4yJE4tyYDd9oOG
L0Wg6qhkKvNMCn1xY1Vj0b1nrG9eE7duQHIAEtyN2q+I4Tu/4oMs2CMamMdj
PBWKQpedpUJ2P/9JpB6I1Ycz3n0hotzTnQMJCF/rDCcYv7zfFLvhZ7occZcb
xETMVb0lFNbx9u6CWoCRoVduEFHjQM1kwaA/OKdCLFP7QlbBwoX0V4ZESoPN
UefVFG9eYzGi0XwV7tyZabgGcxGS6qKOOKsVk2w5ypYk4RgS562+XM1yaNwL
Z/YEEEzRVnJRUshcppbU265zWxfZzs6MtJHJh+AlvCJhBbdWNkxbbRhO45tc
gjdglLwXx9mhJRV+o9uZtAbShYYqZ/FjJPHBOjuMjiC6u6rusve58R6JT3GO
awJnssPJYzLUJGgESWvi2bLcN3D1Xp0/6Nr6ztfCwLOPVizgY3vfryQoRpYr
8sSs0w274UgaD1phPhI7u1QbC0+QlPfJiir5XMed1CmOyRsKlP3ddmkkaR6S
6cg0NLXQKm+IhtsTda8MPHaJ2BpB2DDtmqHdmcU1ZIMaTShx6c0dWA2IG4c+
laQUdhCi7H3jwhi1dZQPkJ/WNpW3Q7GhpR/t217DftD0gLKSnFWRFA3ctn07
FNLTrL+qjP5uO5/gEe1tR20KGjhoIVl0p2I3lQ/Wqw6J3oNeFjFOxpenCl4T
cNVhA0PMzV1GrmetT3IIdS4BHzp5bZfROzTiD8w2hJjqiBeQXbtiEBNdMiqJ
bOByFQ0Uphqmc5o5mxOwQJKQfI6O4G1Tac/bbDCTRSgUYOgEgQ3PIzU+f0wK
2waGkVXJhhpzS+nVV95Henu79lvMfPUzVpHH2NngvPPBpMZoTA/bwpUjzrfL
wYryhrethUkA670oI+FwMY6lP/kif4/pTslUXl55alSD84TwmONzt5kLHUFT
5Sk4prRMX0Czxq1BRe75AUO3o6NkFKchRtHyGkBvwQy5ETFkBYqVeVBgb7vB
x3K1RRIbA/lePKIlqZPvIQqJjm/aHLtLe+Zw7kIuZVb3/uxEHKYVnMO1FxQL
iExBSCdZgm9+NuUJQSHdypFkj9531L3LaAdhuAZn4j27P93qYNR4xE78srq/
VUxHYdtoRI1e/38ld8jVBx2CtTXX8lt3J8NH46jWc/2NxeiUUVgWLIgrvlRE
NgEQcY6+wWQ3R5vYkJa0jTcNTe2xkx8gPxuaJ8SJe8gCuZ5e+gRtQwj0YvkT
SIVf8G4jxzTPz9DDkgaeJyImxf2EaPHJT4T6K0Glxnpu3wj/hAXQy8hiOr4Y
uThN17VRt/Z7Epw7sK35srCl/l1nvf11YKFbDu3gYLI0DY7jm5Y+8SD1kV1Z
Hf2HEg7b3DgU1hByQ3LQY9/32IMpM5iMUCDqXdI8V/i2KktkvJZqS4YBYW3s
+F3niVM5UBBaFed2jV66TVVRoGAEFrDQ5Y+i6s0CVHIjXxbq0sjeN2O/vvUE
DdaHpNmEbHApnzZxCorB3AMkBYpR8S3wcIlEmOe5bVmqZDfore1HvG+n/bsJ
9Ir60QW99VBp3+ZN2PAi1Ic3ILUOqmTtT++r5ujF0w/+iUhDWQtwXG85spfq
ceKCg/jnIaN+RLWi9DcYs/83p5QMu3CMhOJ1QiWDRSFfmXgFY62P9nEaqSIT
PBw+4FMBTJ9cM50jfJlB7mq+qKb1ZsbKiLPQJ982G9mn2LzrRKZWjrw0vqlZ
/eKZN4xWdME4eQDb2uCIXoNL+DfeghXCey+sjvHOsPAJdMhtDvr9XA8fxjay
3+BgWRF04q3K5lPqpj9e0KFmgdwmPg4VVDRl/esn/YVWUTag9ke7BvfGEu66
w82/MaGdJ246HrzdHqBYHG6s3Se8g2d0Z3snTrm/joodw513NTJpT62Xqlsq
WyLYYSSJle4t5lQRwNEO/XnR7oJVsd6gT3uiubh9M3lTFZYcJ3CQQE8F0PIj
FP/CLmDoam8Ufepwpc4AWKIo5ZxhwjcmUQcc9zIUraEXKzAu9p5If8AhMZN7
Z0y23etu7NsD81WPup7LEtpVk5ZSRgiRBuXxCnz4p9QFfccBgAVqPcMtis3A
oIq3U8WyTAmVAEecwJ6ZYApqI/SWYXtVcTxJkGW4A5jVlBoRoQtqYq6LffHQ
0I8x3+KlE/xmx5LndprVXNsqkDye/lljxHrFai0E6P26SUt1bMFN9aZLvNU6
ed7gjL4LMFR8EzI2ZXrdfIBrl89gfgX1AkY3bYGNfrWVP5oCKTWgL6WNWi/6
z/xSccrndWH0CM1+xCqKlUy6YlALimcxnRsyW9XnZHP/v97mQOwzpWRdehs0
oWiFkqeSFNSHJG0o3uKk2zH121o96JB6qEQfZEGTrc+FitgMrLyQWJVjlyFI
5+ihxIscPyk6gY9XjMf8yXiz9NS0/FsSBPe5dcGq5AU9WMIo6yvF1bUPMLUA
RnHL+RCsTBwgtKz8tPsaEnHMpuYjkFKhH2SBKPkuhnWiUUDHixgk3AeHrzaA
C+mkgPOOG04aPi38fMPS1K05wb3MaY2vLLyg68Zvl9avSM15PqAzSe+4rPu4
Kmpx8+xuz4++y4ti8wh0+mikSbp7PVUbDbH4qc4KlpOryAnqgvUByNQQCVc3
BjaoAbngQV9IwBRPKWWHrHOxzee0spgml1xRVZv0DM7BUNUZ7hKFNau4U6Xu
hcB/nnd9ZB+rr81rk1WO2NlF+6Vt+Hkk9U/HDwnLzWKWyixU/+EL87Zn/JIh
Ek4RylOrEK1p0ODotnSk/tQ9sUqmj0ynVe+NB1A8ipGTDo4RPnHa7zwHOrgQ
JkF4mVeY/ew4dLwX0AOXy32GKptbrACilJtkaZtZDZDtGshn1kBMv4gfD/dD
m+KiecFtiUiivaQVi1GCkRn+Vuo6N/714PRf8h/CeFirY6CeDIwuLlgHUgbW
DGzplNJN/xftUmVPWxwqAcN6kzbP6U8JTMCC+dGP0IS0vFRtbKa2NcgCm9VE
Ao9FPt9aJd+6gJBfOp9GvwE0agdw7VdqVmf6jppfxScgNK1XO2y2/vC+mje1
56N2ZZXgLFnD3hhldEeNXwTYXJ52bxom6rJSyw03UODnidPbQ8QxNTqDaywO
ZYY4ZVRUsZIuFjoqKJAsip63qgd3bDQvmlu9Y+G7aD+HUyQ14BKyuwvgx2ou
HBuc+cEHF+yYZ+hLlU+zbtU650KcsHi+GHqR64cbVq1U0rjfdYXxP1wjnVlY
6ZxH4fQ+FQq9C7n4xG9CJaykPOKCQN7n0ietjrUCKGMbMD8Kh8BG5llngToX
5c+v5rp5iNmsVr1z+pr5XnaCTyeXtYQX03pp6cs9kZ5MgsaKJi1FjzmHg2UI
Uv+rs2M7L/OeSGOTIAH9zSZbdtM7aPpMDkydFzh7jMx4rrApumV0SS9egg6N
S/T/acdk8KZZC7mCSnFQp1XX0LWT3ed5KvNRCmlEmeJ61Cgz5PgXvoEjMRra
PjteSTpH9J3+3stieAeNEsA+ARAx5kLd98/tWlNRhDKxBdmfjNwUMFVsh6ZV
sOgmx1lMVwevdUL8g+8OxPT7hTspt25Tz38WvIpx99G7stbso/MdoIpCLjNY
JWgP6/fNDnctJLwXw5UF7IWckB3rqD4zUBDW7xpaaWqHxmipjtY0EIttwAeF
Dj73F6c3KSq78FjZywedGGlW+WKKVQDsptSYA7oKc8t/3DHimizfn3pBgfJ4
DtbQZe6Me8Ioz41ptrYDbk17cnrJB1bwzYnUtKh1ztGG7eTgSKESx7vDYwyM
GRQyKIc1cKfv2qOrwjnLjhWJ5zITC6RSKkrpLGVLrP3F/qyMRHRgHIRx19IL
iSNwPVj1I+w96KRxj0uGcQvljwV5KfHECsjjRy8jkN+sBBZ2lVqjY3vEPfz4
Wg3WUaJ82oavv3wVDkNyrESvT4W2Lgc7uJfai2km6X5htwICuTCNSjd1dWPj
NlNPnf14fsYr8IPVdNawvqpygDv9l4nLJBF3auIWeLwQ5q2wQx2uorAWZVnz
8ASdV6r4XiwuheNZv5+GtVbzZJW5g+FvaDaOqxYwgkiByIq3yArA2qDrqKT3
LS7VicXs49AmX6gIb60o2DvXhxC+V2wQqyO666AmhP2ZkPUqB4ZBRcnPm1tg
CsxoG6wRGgk7yw9+qm87nW6B+tLVN48RsQoUZTE5TaxdZW8RzDgPS0BeoLbx
okO7nm3P5xNewzuuithJUrXAADTVBhU8VUXfmUG5JhT9ON+oTzprZbvh5rKY
hvuxQJbBBBTNRd+6QX37U2PVzfl08ggP//vKwCDz6hOqnhtTnTI0x4DhLEVi
bSf8bRpSgYX/hOB7QGCsQwsplwYqeDnZ8RLTpc6zteXpYXnaLUpTg0cTC8B/
1QudIpt4+Z5aj6or8TI3ixWxhlfWDQPvcU57HU80d4t7MnnkXJ2OoPvEGzOx
vwGW/UOYp4xr2fwHWL+cJ7kMgU6179nRMDZc78hpapBZMjB8vLx3B7W7QePJ
aFr7ZZNH2AguqGeglYxVzihN/QGDBjhJnbEGehtXNIN1SbiMDj+clJb1St11
vW4Wrx9ucKkjLk2Sxbf5z1KTERb5HFQMw4jCIrACpODq9jUu8Ja54Xb9uJlJ
GSZpxcMXa3K7eWPyjhX4Brv4sDW2mV8u/KIB/h17MmOjoD0TqjUVoDo/d/oq
6FfO9cmoxPK+gB4UdF1xRDeQLbc8Wx6+zQlw3BzZg9SeVnyhry9EznIYYGmQ
kF3d3g8Jya7gxL6Kmpcdji6pUhCzgRxgEY4SXICl2LtuE3x9FdfenKYRQQ6m
tnRIJqr9IeORcnsREn2l90yKJJYJlGqqKerS/9VRnAIlA6J4h5BCfhT2Q7mY
v1W/FRpYI9eeTnRh3pMbdGcK7/y72r2omR4ksP/1faEMljWm4+SuDaeIIvYf
cVbwxPvbLHgq9/INEWyobVomVs+4Uc5egTeCp3SuPpLvrcR++nzKYk0gOYBc
Xfwwu8S1Lurgp/aPgytF8behODdFVZqL+ert+QeoCWKCoeKPvYtp9WwufUcz
ACpGzXqzIS/wOZeLjlLgmkwZUecBNnXU68N9ZORw5mslSADQ4I/++IwYJ6Zg
PyJMbUn3wBd3EGSnJu6rBU+JCYrrsLqArtC7GbHML9NHfxRfPvLUpjY+9f9h
/LbiKy2cbPMT2TvvNGzAJgrRLdR4Vzl1/nBqumJRTunIdqRH7LdXKDc9mZh5
B+Gvop6Oa8PhOVYjkWepfbMQseRi2lYNE7I+dc+G9/KzGu1WpndBPGlXnPwW
gd2cwtRMJiqbG3lSaYLqH9+75ekcXgtVDZRvdJZefNWV7vY+wG3krAgtYldd
/xmLdbJjCIxXn4tdGTeuIbCXKsPlzpwS9Ho2ibkJLlPa0hQlGTJUm770WgJQ
ICNcegnt7G4LtDl11U3GCES8rR4BFOmDz1C8FZ1CnQgwGXdl6K27Me8nrjmF
L2wvlba5HO7Xl9QBqp9JyUHzaL7pbw/HnHb0qzP1mL7E9BsSokfMpPj9UgVd
2JHud4nYtvS7B1Lf3UPcguaeP6LxK356wnr/z/6KWLXlMYQIwcI+HgT32drT
zQEugjQHV2GGzTKBj+UPlVJo+NB8+w2Fa/sGxZ8l2TSQ0Fz+lyCR5NgL+4oo
rVDSvAxi5bWXCGsAaC/z611QbjOnEszFJS5Tq48Tr7+bH9cRNRklI4jDJ8NO
0UFbnOby853HsHx0V7gtJlzItaLwOlV160IOwfay1Mu2vqj+ySP8a7zfNYep
9CY02Aj3GNfhd3+6Oi4+oSJA7ULRLZoeF4rY4RRGxB5E3gPyoTp1WjsL4n9m
ceA2U1JF1fcFC/U3GPPyfNWL8gAcMZWfjB4+xG1sv9GfcqGh87n3yZL4qL+s
WtGnm68js/G6JoliYlm76lXelzrUlY8rlZKJvpZ4m9eDElV3/BfgPHLbsjbi
fpJhVx9bzqAA5Gs315LWR8f6A+tWviAFbDfJW+5PwvL8DwB8vMJpyEfiKww9
U3xX9MChHJP/Cm9IUP1lAldeyzUBNBtzx9V46W8NgqGiiG0hdHWVNrxVDkVG
QQnscgREBHf6FgPNVFJ+1rMUE2Z3wXgSU07VF/MpWur6SeSR5kxGVJjbJ8G2
GjjHqFLYfEwixw94JN8ta0oTqT98+TKAC1N6Ll6oc4X6n6z4E3p/x+M1hDxT
Q+mQSRL0dj0mdJyAlX0PonTTsxV9kLWoKRP2qhVIB+D3m5rZTacSnfh+n1OF
8AdZUt0YbnY96N/lZ2eSHf+F2OpicG12AmE/M3UxDpbnTIm8wKqveqRk1SVF
HQYWFB3b2xVVRiTqnYpU6Ss5xOU3PNvxHFjD95+Ngg7vREByAkjI3k2YbdpG
u1JXImCXAOOmf6Vb/aXQNO7ieSMdjyA9mRQ+8ssMGE1CtlG5pH37nc5e5uXI
XkggudgGPiyKstazbuMBakFrBOfggYj+K4A5pEwKE/eiBjnyp/MXhrhV46K9
v9uYIN3NJNclBeNMd3Mza9TmU9bjFIqngnuc8/VJmsTVSS+SeNfLPSttSS5R
FXS7gD5PpemEJ9hG6qNqk8DXzNGW/X6y/z5nSTYx6AYTWpBCfL0KXZaKXNDN
gV99Q/desNrqcAJ4SLI6QlCW5FSdlAKcv1Its+kdOGV6efZv9MH7K87YTwTi
jyMCA4u4cx5H0nvFxpy6rr7araWmZvVnKagYEbSIjNBC1LKq9BdYFe+1+MP4
eQICNyL0fq5oCklYW1iF25hOpmv/jgO+NJSy3hwrxQOIzND9k1ms/7813m8r
Yi+vjkPKxMIgr02cjhsS4BMUdrjx3lhnCkQQw61yUUzFssK1jCKyf++3EEsb
UyLlUTTD9kjFu1tJIv4X5hPA2cgBxmhKBfGwymnf6aGBANn7sbLMSH8BOmz2
H02xHoC51TdRMQNSMGxHmPio0mNvWCwdY88/9LVZqOtX/l47VfME9kZDG4h7
Z71V2YgQqZsDJfhc84tbBMBcmRG1Zp3Urz3lD2bOj7tATbPrMsl4iaBMjSE9
ri6HSzfAN0kF/2aNtIBkow+kbJwpiudIjlfNXnLiXV1m1BPmM/GcHtM6IFtn
ysix/eS9EgIl4rXpIb6lZbvNdTyq1mLzFDq8XZJv3EL5AC50mqA+Vovi0ykO
vsOsWRTpABl1tF/X35BumJVQVprmup305Pdxmn0YwfV5sM8CnbCAJBp4LOW7
LpTpFK91/bmAngHBHndt0JRA4D7jws+ulpFRi1v1TKk2YJUn867ULPv4MxZj
RKoiGZatpMEvSd2uqyKDVcysohQr9fGuV2x8ZcDegl7O8cv+v14cYM5v/l2f
a4ulhhCJ6R03eWSddTj5WLmvzXAelImEGlQPQXi2EXbf3YXrWmHL0niKo691
NXRyBBSwTVyH0yu1wbcUTzeHnwCRFmJnndt1zqqWUIzaDG8hEpWjuaExNq67
PaOu+GOMikKEPZBHdIUcIGPFo/i5B5OZ5sumKrLJku1sbAnB/KEkCo5/b0ne
pqbpQswgzmOaMpihs9VPFh80KkQ2I9Z2cg8gbfFoc4M+7HuVjHIxe7SpLePw
bl79q2lLU5cH5I0xTxLqop5XVo6jZ43ZaCVjrmXbWk/E3NAWnDF7ncBfwxVt
+AzZHSvAMhJCguwDIeG1Y1H7X920WAD4nh5KIWD4u/T/1X/PqzfA3ctsbc+p
Hevbx98VtSx/7BMjeo4o5n3K0+Roh+SMrTxY/98dKhBDTViINDM5WAoTy4mk
HGDO6uM2g3BbaOhoCoR5l7c8DKOfrSyh9atsuKuAMRQa8BWVkcRb1wAU3/GC
flcjEsa9T5vq9A8mKeoVzFHG8K0gEzxAwQzi9bOd9HmCeent30z5Oo2B/xDy
PCN0r3VsdZUyi3fY8CwpAu1jTR6rMAG1KEYcJWC9lrvscOCJiciFoNlWi/PG
GRIMyy6tPt1r8DPooQzU1p6rC09sORZWo6JwVnFwp7ZXZa26uXc/VaUoBpc4
fgg2mPTYvVj94sF8oQkJrx3zVIZ2Rl5TyTTrak1Q/Sanmbo09GVZaA9MtB0P
jiIE6xd8qHIBfgIYzeoGenrDXma5WgIi866ch+RVcNTC6gnR3zs6o2LDVIsv
uCQs/t2R+LG1wme01SIK33NkHJZLtqkOyvjt9257ce0q3ZfUPctQshY7Tw3s
bK6RMNtQnPi/hvIa4plGIg0hsi5I1GmKS7WlMEyBf6GhGOsvNfMyZpW0CwvF
R907OHUpQYuXh/15G99+bLqz5D7TLA5Qw/PJcgQLRfX50zISpFex/kcAo9U5
nxIgWUCwae2iwbpcbeaex7Aa31vNnWQ2hYT533wWQEW1glGyymZwkEb8uCvX
wPEwVve+X+l/u/qRM6l09dhV3wSPbF3o0wrtFRvcbT4Up30M2qb3BEIFANjE
GLXC8aCS5TNbdZgbvCU+KQYzc4iAYVrLTZUHl8Pp517gTm1j35f84zHQOmfi
Qwb035iE+btLE0iQtkVCcyXWSLAbLc/kZxWZCEHo0YGIEt1DdKlAvXcjp3gq
itsJBLqahwt/1htSEf1UOmKuikWQUKKlOSwUIKxThULwpjUU3K4JgqwT7yHc
cp2qX5Lrwpx/E1zvPVa4TKlaMlylSbUofRxep0/8Xb62yOum8Dlyvvl20XWy
R+iwEMxlo5lczJPa43/g8G+ibSYi+6NfsYG4ZzDXQuydQr7eDaYckClmhQ9r
Tu9DQ7SflRVZLpg+tfrsCuXgfCls/COpVbdgierWc+J65w0ry0CGPncA/N6v
bmnD06e1ib+d+GsGx2iH65mT+Wqh9EymT4ahMa/Xt1LFv8SmfCIMw5wiTZDE
OGVvu29PYeNXdpgnm9wEOxIbQj6+1wk8x03taMYCbRunFYzlitadwARxK6Ja
z04+tCODyUuFarQVGUXcepzkDX7kNKE50uMhmCjg0DGym33W7fo+/wk+9qMX
ewonN8AQv9ECPd1gEjZshN6yuQAqruWUFq9UAEvj7ilAd8Ia7CYtYvwL6mkc
W6lnapFvdlgGNeLkzdJ+YDgYOIsuY6C/llDlbi8a3NLxFrNdNuN7pjjGXEiS
HKcJrEXwZzKlYIBJOXCiQzXYzgdpk1obPr36fu6ZxPkRZR2cUoB7Q1biK1+M
5f9rUU1q8VbRutICAV88r5OBjGxoMGkxEAnxsBVaQl+pkCn3MnjR3Iu+Vj3W
JJqM98IifjKqCJkrjR6sPJwnHq5a9eru7HCG30EQh3NW1qwGyNWuIFFXOoRN
eU9tUl+W6aHVjup2SWgCoA8LebFP9Pc39RBYiCvtrB4Hpz0nJzZ51y4O5h5w
phh2LEk3yR4dcR4QOMox9LhthnkojoUJgDHBm1gcv/CLqLRczhW0Gh2ENDpo
nM6CsexWzkxX8cDNf93obCl1fUcKspyDPLhtoWBcguYxOKZYcRi4AmPIT0Y/
HlL9S8JySJCwgTNyuCBW4AnGDXndcfD6aCHPG4zH7Ou9Ua+SRcsZnAe0Laan
uN9gTkEdzVxfgMl3vrWHCGWz2hm9Vi9nfh0KKIUjCUGP5vysEHWAFUXvaIHA
CzrUsUCZ2vSkt4CzmspduA42n+/KLDnHvmSeamoe24x21azNlESu/ZRGM/MR
RtDzp30+wV2ocvwylUA2nh4uEl0iw3KmR6ugw6nD/FkFr6G/LXW91dsqTeCM
2+f0qoLK9DmU4RoXFDRLTOTNrekXMAuG6FC6uTyqwUefhC2E+NYqj1W+iP0p
gXXXVUgLO2TFCtn1F2DgFBNPnLKow+llIe6I/WPOAX5I5jksEvhavd2C2+rn
9qB6Kx2NZAr77bDf/ItM9BO52JJ4qpc/eX0zBZnxcKIPxkNkzXTTmaoTqnTf
SLfo/KwV24ddHNG4FaJblLl4kXk9x8f1sbs62I4wo/J3l7giQ8fesib921hH
CXgCf43K34aBvgYzu2cx91megnsdD/8NfPUy41R3qGn0S9hmwG1OLk0bwvaE
QSapIqC/L7wQnikZdMa5K9hS9xdoVEQ77HaQc5iNySy4LAMQv1iqGuzqRxC7
ZU1EXM2uQ/bIEovfTQNja+DDNfrtByZ9Iq3hgRvNCdFjNO5Fby8UNWI5cGA9
jqWP5Kv2Lu4POgeDUKfNd8mUz12QE617tzcwrtrwJQ2o4SI3eCbuq2syIpKd
UMAxvRrpWV8+qldgf4cwlb/lJHZMOeyec6vcdyFJJkMB82eOQ3oIcO3HSl+x
NcChZt3ZJgLomgN70Wls0GBqe/JBYQAxUJ7Cbv3sQriiadtnW/e8OamvtTKZ
Dvi5vHeQfO2XoHLQix8O7MPrvi7beUMMuL3hTrDftU83Privqu2I14HKKlHh
o9hOZdWPzL3nOOHS+9gk2+mr1YB/6qEfokmCqtkOa1j3WU8RowjabkNWjxdq
Pl4AbwuBvSnkCHnoasGlZq2y4wdAZq9e+mno3xwWHK3SMPNVyUr3d5act2vM
+tv9Fs2luMGfAlN2js3Ez9D8oEN6gu6SP8O24llKD4qCANxeNH4n3ORMBsFv
bB5t4jkOdUUI76XdLk5lE7jVaAqVVa4zMndK+qrgpgLMOnUgrt6HGgqe4IYQ
teqhSHUnIWnhTv8vk+uAl1MfFOUBAQrlzeYA0rpL3tinm/GaPMsh31t3KCEh
ak6ldkWk/cbf9YurdCbFg+STlO3/SiL+0li5qPDp7w1tBkWoSqo0Zhy8X8xc
t2zBeX5my0Iajw1zYH6pjYav7O7V5uLuLA6am+arnb8B6VVhSgYwYLTKL2an
b5HG5fuyyy4hBQovdtvGPdJUHKcQKgMVS8OI7yB3dwHevAOCJnARUeQ8ffdC
YZDMlUy6VuuZAdsoy7jtuHo9sK3jf20B3UGVtt5ebVAfBFIXKywC46wuT9MG
grbjtkdiSfeBYIY/xE0KfPiZc1nzL152e9F7kRQA1RP7hFRJePjJBjvcJwLp
bGBkz8efxB6bD7TFsjPfvoxGZZDw+pkoCnmij3Hv9epLE/u3/SHIQLE0V7M8
Cv260EfeH8M08X/DQH/gEnC1a89ov6f+th+gR6OavgfdT2MnSBcwgMJLXfbf
cN/1sgi9LxxvW2f9dCmFhLizQ4cCOmM9nLf6ZvMmYBQFIhdzO2TWcBOXf5yN
eslHNLQEwObjVrcKN+XPHTD7OFfbSY2i+Hd8ezHLXcZpGGPGPw01jtuf2bgy
GcpVKwpJIQiq4hQzz+HhP9CulopfaJ8xDdFf7oOQmVMfQb5NQmG5+OgDWoxM
lA6yRvpke45ggXwUo++5GvNsEcoXGCe0rW572+GhFNUxvntJllBvjFO0+U2j
uZE07W1Lg+GFKKCM7CmfdeWwXQ/nLByP4au1/xYOXeY+OgamD4ZbZRilNzWk
dfoysmmd8iSO33I/rbrlbL2mBuMYaSyLTNdYtx5EmVPgWCH1MS7Szil5V1PT
yNHozBIldCtqSTLxgXfLe99LLcjuWEdYirqufakixHh8k3HUi+dWTminIRlo
CfqSd8qr4Ozz8p1IoUwoHA9zZBmugXcpA8fcIhvouRwjYYB54bY1rIVU3bJn
6cGSSlN+pwEHAubGnDziWqj68YHAm6BwTbQVAQkc2+h2iaLdIynhYausGMGb
kyMzmrEAhNizTL3R+joxQxrDYxTxgVZCkq1mx07zYFRQergtHgpBq0VfLqOU
vWZ/52xgYMxFoLmimNljocuRQBE0iTyXfZhffMSnZTco5S2nLrtakpAi+FKW
29Rf4VqBGZSmFTjLuRtCwlle+/LQOqfvfyImiI/mslYOczJRSnBDXliL7ccx
0GQuZ767h4HKEJ+04GL+lvW22QQTTT/+94PzV85ULmZWvoPPm+qzQLoXHYgJ
Ujjc256oZXFY+hRIiTHvNsRCuHNV24ITJucQ1CaAMUaLQZE2xDNuV3BYIA+O
iZOTtwZGNdUXL2Rl7XX88aM2ptnixc7YswqWIGyh4pmhr2WRF21Tn/ASPeWv
JO9rEr3XWt3Ym5Phu4JkWjTz+mSBsMvPsOxq0/zooS/kgpa+kipSMSjX9u/Y
9eyu8EjoWbN886vVv3GELJRRqMqLWHlSrvoTBRKiBiuOkNJ/CJKE3cexp4MN
eQncNJAhJiuFH1gZjhEdE91uLGFXyASL0GhygQP+IttbcbOOgurYp586fuMJ
ct9wYzdPYc8I7ZduKz957idyy/LXcyWC6YAo+J/dTS8vwm2EJqLra8i8VHwa
I3RVflOW9jBAFPFFGR8DzD4NIrov6v2HR06cebSXtw8QLEr2KBsYDJOZqgfr
w1pCn3QaIwGgPfKU7u6whIkVR+WXmnL3eSnA31eSeZKQuf2bmMAHTeq/ASnl
EmLFedhN8igBsOx5tya9NocKAgAkrybEc2eTaGpuDiWFUupCc1eITVQZcOLd
edBziRzKopiyGe8TV6cSB4NyFk1ctlvWiPF47r29OApJH8kO/0JzeQIWfmBb
boyJQqMKq+ZxtoFeGzgXaWqY8UflgD7PvN4TaZGOkcVbTwH9TlkAhzqzMtxc
pm0k9axH2PwcR8uPafUNk3+kYgeyyqkTcHoTB6H14eBbWh0GoftdA/qEViwY
aqyckvO+h8U5JUYU0ZZZPgtybHuaZAOO1FGzvd+i4NHgSVe8jUgl90exdwiw
2KWtuT9b6kn2rCXVEJSLzonmt/FcnB1am9sOHxjNKW9FsF/3WPu84ZHM5f+8
6kNVJc/e6VXaeQKBCW706JVywYwI0Ga3vAx/fUUlhrYIkjfPczXKy/NbkxnM
iE9+t4R65W3D42tiDMldg6aYXMHn4vBx7ryGgpzcMHbDas3ZZE3Q4Vzc+uIL
WyCyIxaBgZRYY1Y3vTYEpImGaQcKRnOEqECXbFBdZXpgdhZvfSLAF4rVcNIS
R4hKK09nXsJvHAFMl0luUE9f6LjUQstOetZC7yGRW9UTTBDgYKhuzDEWh28y
YISBarSHmcv8dy2p7FF4wYpPD/KiPAeeiX66Efyy60gRFD/aMu7/PwLkQlYs
5vuCKJEdbdHEG7fU/4CvERAG5t8fsrFN2t7zWaHWk5G+8qgHAeudFXs34A6H
tggfcdpqywKIE1avx4uGkIc9k+40uU42EML3BBDRwmhMXnvdyW0Jo06FiGP1
+40AwpUnmxzo/4SAkkc7GqH0gKMf02nrT37g1NRN88htDjblkKFfR5DpcIdt
cFQiOEYw/M0DKdTCg9uTlXcl3FLXjv4WocSvXyA6ml2zMz7O6OAZAgmul1CP
i4vguSFUiTN6YaaEUkwsGWZpWH1kgT1T6VvRDedwOflqfmwuZ8n4wuktBqAx
GVyt6xHOhS5/7WIYXMrTdssPAm5ZE3p206SwWq1MO8e3+JqQfT6O+RfTstz/
f3JVflzpxvhJrN1hY5mdqgjsyzb9kjBNThrdKmwfqvAIVTNQ24WbIqs8rNlF
lylUeT23SrJpT07rYJtO8OEbs8Q8fB+k9wJM/rNf9PeQne4tfwOVc+4B441k
N6WrYxtwOx4OjM5au8spBw4Gb4S7hYmiSxEkC0gHoNCKcwTRRdbPF/JLCm2t
O5c13Y/euLheHWZobTQDMurrLZJB//ZCB/3T9T3rgAvCICN8NEhCfOg+X2HK
7ZdHAVbmTAeeeuNyDdrl6ZNOvKfEXcyGCP+FPg9Oh6HLplGYuPa/YQw41J7u
29mDm2BQ/vZHVSHym5vLtdefYZigUsJ+KEfAVcGrRVBs96xxlYlvB3h+KuBf
roa6OuyVLZqCxtFSIXp5XppED6NF4Gil32YN34nwJ7rAOJWHuxiK6VBG7WI/
CPaaZwQz4/Weoqeeyk71BD9BZDr70GAgLPGChqDJMvJeHfliKTx4Q/XL6PtB
jETgIcMy1+B6K0awxc6CrCzBAKyvVwP/9PyqeLHGUXqpUQafQvOIOW0JEu4D
PNNySvZuDVrsH8A+aX/5EJ9nebnbUZxRcM5SiAImo3kjnCMpr9qa854uof0V
5bmQ+qbARK/VFrxaEem0pDTx9NkFQKhY4ZnPqmdy0/iEDLnUyoIzy6LDT2JP
En7yjQRwsL4Dc7vBpigTv/CFhwd5j+2UIXQVE6xWNB15Ykn5zJMxhaYVk/81
egnB47MWfcJ07OlVBIbIW8LtOAgF+3c4h8fPEdJn/4y5Xk5sz8snq+yKY95o
MFtRYrWDg5WjV8XJC0+sUNPQgLhu/H0RPAsLtWd6j3Q2h+Mo5NYrc0r/4vrC
NwL9tVGJh2sMnT6GmNn0ZDtH9sUPF1c8jfO8zi4xbXIFC+KJFclZmtCLw2G8
O4fz8e2x0kqMbrXzY11IlNusx1QN1Q8IYf/xewNbYKgOCcUTwr5WtO+uhkWr
tUxLWw06Sw3rNbxxS8EvJILLEPO3QZmYnVQ38UQBYC1uV+OGihh58zQ2dHdb
piN4qkHvoQpuXhNAV1VsYo4zG3n2z0gebELUURfyZaOsRu8e01j85RnYDiNP
1r7jdHXBJ6eqLamnja9qcoo7rhaGckM+f389BtyIanUWckpcgIxfwIDutxz6
oqpcKIkRXGhiE+6wtGXpMDatOSKYuciImi2KX+18ReJS7memV7ei2TYHt4sC
8GIiW9GYX1tlZ5x9bcPbhW74MpgZQZUQBXbwk7u/pvdPAOMEa9t/amxuVTC2
DGijcHKHQG/xRjl437j7O6QLQYntPf0aBvJ+LOVkmC8itGp7+b923Tsfu5Ju
lnnDni/z6XXAWSb8DBWLaVWOWm0axGwzva5kZmD51H4ruvQ6YMZecodqopno
m0mC5oDUg7PyeJA7//rmvTLG6y0+IwKnEpmjgamkPOPw3Lt/B2yMG6LuGRWx
ijvp9imCNCCDAaEGmTKVX7fo00XYnuarWvi37tViR4sqPehzIB6U45jgKFQq
XEX+Jn1CgGUcYlE4VXdTjFvnyAsEkW7rM0fJpkFXtZXED8cewJwMsHtG073l
/IQ2QMnImr625VNygte1uIUBoUwUbSJi07/i4JMo0eccdWYJ0SRjQt94MIsv
guiyqay4J2X+msWHfsnodSSzr2nygoOn+W4c77j78UtGBAoXXMQTOB1xLAcQ
9PHpZD5AumZIrif9xuAUWTkPrVrpXNJDdK4xYZzmS0QYVUocl3OYRvIs/bJv
2jZYIoe203soi/NER6X+IB9Mn7yoTAMZYdycyu3psthv3bY+Fwb1E3dvLCUY
J9dApsTnWjlKQ5/XzFT/1o9MlSA6bWwnAZFxLj46pM/oHfzyA3WADO7mJy/1
PIGGht6SH3iU2ZBCRO0NQ+rrKYhSeYoIrdb9wbrvVwniEehGXsyVVe446y+m
5KiaOPsKiH+rtJc6K5R5vhvoS5NPVOk8w9MP4J5nxxTLsywPZsMGLpAOHx4U
+dGpah8GeqcP7C8ZHbj0PlgS+Ha/ErMlFdBXTZm+VRju7fWr20FAAzIWd5xO
qYZRDSGolubL47xpVGISu4r7gb210tOIGy7xuQMICNNXVogyClrWf+4GuOwk
Mm46iXOwnv1ENTi1eLkbG2BCjeR2JZJtNNk2/sB5EDvuxBa8s5H0ySjLn9Rq
xfNid5SrK8YniEKQqghUMdR9lufZLWmrFtLNwl/7qX4/BhCIB1gJGq9OBUas
xnO5DlS1emUWKBuK/0KCGj6w4OAO5a0MTMl5+sX8pO+11Rqep4IoJ5d3FsnG
utvrt7Obw//4zDWiuUP0TWJsVCFBb3Xaqyan/4tGMPUtpWFgF0QhSzdeCn9Q
uSmlZ1r+9dcZ36qgc+Iko+BWfbNARGgoTVaqINnlpRV7YlIAud7y5FHaQCeD
4pLScpkOp1ZPQc3g0BMdJB0zlxJUBllNwI2b2e4Bag4+2mnz+l+Pby5RNWOH
UBWoTBO4PNF1a3PImB0UMwRnFJLw+jJfPuleM5nRc9SvQPfRL+hw/FDBoFN7
pTGOmWTGrmXdmBZF5DzXsGlWTwbZTPzxWB3l/Aqv3Albt5iamAIH3H5vu5N2
RxZpRn1nJM5lyP85EVV6YWKh+PyMjLc4nLgalYdHH/gHxotIDH9Zy4QdSx/e
Gy0nHlKP6MFBXEPiSQ/PYxMPBlxQhdHFgfaCzlPAv0nXwWmPpCgC7GKGiux1
bQ/FM3px9HGPEpsTRI/X3vN60n9PRO3DTtqamb0DZlj2YbrxMbE8UizfK9yP
GvOleDIF7kg02E4vXE0UZVLH1IuKI2hRlaxQ6ET6PDQct0eNN/RUjPXzKGx4
iQGcxeW1GM+iN3uNaEZwiMmu7f4rJ8qoQb7aJXwjcPl3+UU82bvXfMVAUN8h
RMtxnZ5pMlrRu0lAkXMHEiRLkWGx8kt6gB1Dtj6gNtXwgJLJ7abXtkery//b
9vDaUBYOVSLoECu8pOs4jBE23lSXHQCG8UY9PNOuKuFF7bR2368g6+DtLbTF
aA4gr0iJfDNoTeZldFqWcGGhXZEL7hegYMXZhsYjjf4onGd6ioUrskg4BA5m
+bJJHWhXwXdscQXrny7EB+JlRSW+2nq4Ld/QpEaLQXtvkliTFOweh4FHkkov
o+mjeRGlJgQtDI0nwC3ew6gNtmWpvCOSMU0Nza/yPQRBcrUVuE3D55GzQjOS
ZQI+t8K4r//cJ9YgyB0NeNfpxRQNIBWDLtgKCojOWm+ioZw8m4TuiXICKTCr
VdNo0nH4yBNppcKbkmEmNm9f6p6VSNTdWoDRD6GtEDWMVvXVivFr9dW2Qea1
MSgm0K7AI0zkI6u45pba/ygIukMKwdpDoNCr/604xW/0srLQ5hFL+n3kRtK6
JsD6LDyMQjs/bLK1s1I9qMxjHGOBlMCR5k6INRy5SxBOiap3lobr/1ygX666
QcNClH+mk8lKIK7zGFyfHty/KwJvbFJ0dabu4cayHmV0hZEclQj8iTgAW8p1
89XK3gxZwVxcJYQiUDr4w+aGECAHnFPJQyBOron7dQ/Qq+4m8kvT+qpCdo9U
bzkmWPtSZoH+/OfOg4bsFj2MQF7eEPdIwQOm52g3WAxcGj/r9WtcyIJWBwu4
izTKxILRu4+EMybzRbiDs/splo/WPbBWOYbgcWYJD8O3IRwEyjLgTz0n2hKs
F9qA0NUus7timoN1Ouu8LQ0DnGvDBR6UOERcrroHUvy3A5vtNO/5NSfSho1G
Byat8ZaTcaXM0b4Lf2H8MNZtIV67hy6zwxqIwQ5TTkrBHV+O0m4W0wYWsUAt
KZwYEjRk2CQAWA3gEQOrJ9BCl20OyPaohc+yK+84Xzy6KryMtt8ebpqmVkYY
F5WUmGjQ3mm3BgdaPsNLA9bMVJ4i2AQ04U8Eg4RrJox0xZcRwbjLpgURfxBG
aMGrv2f3pOrzAzeSWmx7MYHr8x8OlMEQwKYBjcliG67GNVmp5qjHLTgMDXjl
wTdi078wUcbk8Tzl8zAGPKC1kvl+Bs/fNslhha3dWbYjfwYNNlXjZOO3AsIU
fxgEw/Av4Ym/uXMtCNDEs2xTpjeE2heTZxTT5X5wfhTVQmk/+4Va/WeT0Xdy
LI5hzoheAvaTuYQcDNvKShnB8HZD26WXfDqPpjgXECJTGWLl5aXKbI2XUyah
AyE9qQ0PI2NfMGrfr473fDs1KZ4VxKznPOfZc/SEI7/+TqpmH0aGcFOAbbvY
fVhaWSVLqG9oqo1z2/OO3gwXdKFs8jD9Drnj0u7UcJxycDMTaXllxJcPbCZc
anElLzhmSSHMH87LLgPc2FSV8h2/QNyMRjb4AuKr7bWh/3Rlh0caqMhsoy2+
IWJUnm9pFntY4tCqhjTaBE+t4QVY9oq6sjWs/hghaXQN1hkd5bzsGoGDZ0/7
os/WIvIBeeKxRAG4gzjwZ5zehJ0Rf+wxEsnB0SC5NE1MA3NyXULryQnruOma
rdIUIgZ7iIaGDpsHBro9q+Yaay23jJV0Fi3tXNyhYjk5rycTs6psL8IMELMg
RdAd2hqZN3Y0nF8ETkvH4RhfzKNd913Qr+0kQj1TwMdNpd38C5z6fYRcmUgI
3/Vi8Xm6k+8eHX38XNUo3/NbbjJs/u+xCVpZwM8YgLL/T6KQCyzKaHNs8Fs7
bvJXNQZN1PenX0D+WeY1UdaJdk43GS54dBhlIYYC7v/Yx1hlsNJWlKTg2kZL
aoAYNYKEh3ReJng1uFJx4uG01+yEhV9T+H7i4sq9h2UIF1YRTwPkPPR3ziZZ
HRFITVi7JPB0ImxTEadLagpIOR1PhervqwOMN6dPcWwxDvAvdNPGiQKSfleF
B24MbAjf6kbyTzyVCAlQNLjG8jz+p9Nof56YeC9hG5rBfF93vxcR1dHsqFbI
NlHKPOrv2jsjuFWBDArmwcHmOKNmxoF/53vaINo2TDc4h9aTW6jEVKtqgk1R
85lxztRgslNnfcwQQkw8VaVermdvIeyVQzYUj30sf+J05nksJ3zgrwsLMQpw
RTPiic8rjvzNnT4lmw7J5HLeVbaP2W6Vru1C+9mSOR5Ko6k0hAc57BMrI7/U
UAGg5BXgD7UXMCOHpjnpMiSzBJOgCRrMc7uNmGvVKs8xHDjwuW0+eumg5+Vp
Pc9izW3mXiTzaDnu2DL/Or/TRUypzIQaZa8vVsadbg/5TspzFh+/DMW52J97
uHpQ5jLNe3gWTwYhA2CVxWOQXV+OTLprdI5gvTMzUF8hIO5gTlGEfIdGWc/B
mmKyHkAxor6Xmysp01yj3IOz26qlCsEA4lRjbYMsR3RRC0+ZqxVIPav66TMt
/Wzxh2mT8vlj+9w80YOPzCqh63He0Q6NxIqbxxKg519kRQFC924lzs3+VPBL
P0Lyp7M2cuUHVMwTwvIftOuVDmfZlHf22Sz8odleIKaZjlHlXbb67six3WrF
7XtWW9WKdw1oGmuVz21MkAedmXzthtVPUwKn6ITtSeY9eR3ISQGVzvw6ys+k
RhG1idPRpd/mg5+jKUWVSVVVUGwt6MIARDJSnYde/Z1p69xDr/ruS4IoXEwX
E6uD9pssT54drgokh96ikxq1JBIxkxhsS70Hipy5Kdlsd9SeBB+RTxw1tFGP
xeh/lG75r2BNAneV8VJAhn5H1SN6r4R5YXwb4/oFmo6Zh3vBPsDleI0WGhNO
Z7HaqLFX89XuUk+b8DW6Q9JZ/SwtugBCJxNEIINOwhHHqzf/x6LvgUwBwYgo
yv7n8uCbDZO4uIsOss61emWsF0uNELrkR2nwQD+LINK3f1m96ICOxBsFQ6fd
EYjH6Xg8OwrCDLt+3SaG/Ece+1mSy4+K+VXXdE02PP7YQiOUnu4V3GfTxb8S
yzQDHG7XPzG9w0W1MeXjiRFaGU3eZ1N11liiNPyaYPZZiGMlu8hcWdSFYAnE
fcULS1o+nSlc+6igw+KcVdYAP5EYsO1dKqFXracbsmhkB+1ULlQFUitnQ60i
H2cRnPZmsuwSiMDw1lPyG80W22WXjGGGlvvI4kHRAeR4bD6FBr9ITyYV4Fbq
qcxVGCbY2i6gcJToOCCYhQ/elOE+uWbWdDtLAhiChau5vcbJMVPuqITb6St8
wGyvDJR+yXUam2eVxrERs9jj0l8Ya2J6rBUDTvFIgmfmqoaCOnEOwhHy7Bb4
LtH3HksEqR/zdrXVTxGHgSNhUWoXYGTBU71A4wjVK04MFfmHBKD6Sno2TbGY
wlnQZrFyecFYaMBEUy1m/kNjAjQGCvqBZuYX1+Tnp5i9gixUmEsAZ/tQsutI
my58lC2uCVkHQ4BXRNJAKEsNiOkU9dBvY2SDrHfh30hvLAPOk/9EaN5YUCaV
ZcwIh5YUqdCaJ2PwN2A2a5BBU+PtmzVaeEW06+UO0mRkmAHqyPJ5PDxvj5lU
C7F135UmPzHH8FdjWA4tkFqZGjeykuQu5YmpAfEG3G1lSqmR9SIuYQhv2QPn
6uuQFYeIKA1psbq46Atv0503Fcel+He2RFrMfvmC8jqyaYkhKh5crmiSBgxw
J7aFFStm+A6R4HM9erT/VufEXQLIpG6o8HfB6pdsqJTj6O2J/dkP3QCEWlcT
/MZOH0yDAFwLsbUmg2hKSdjFz5kgtzFa4IeNmcwU67ZtdptMnlmYgFm245K1
GrZIWvDX40FYRB5e8hCVMI5GRZkKTYNdqTez8g0I1c2wth+96Lz6vGL72moh
c7iHw+O5sd4wtU5NqxgRJ0Km4DiYPSKwkC0ySrNaup+Xa4Th4fg5VKTcC7SJ
f1EpDkmrlLi8C6QGjvDqMQGwND/yErM0fxIuHcxzeLe2wxHngdsUBDj3FMO6
8Yme5flb5dF1Xfg76cPCpSQ99L3359fVi6B2J/Vkyw0suxZXt1nEjSY1NTA7
/VN5Jn5H6y72DHMpdlHnBFxvzH8Dn8OEdZB1BnGxXm+Cd3syanFijNJQOwan
pWiMiqnBD1AhaBId/Z0L3aZd3ydpLWqXO/wFo4A3dcg5VTK7r6Dkene2br6y
oIPtZxijHjtSyWpes8BXtAHTXb5E6f2JVhbmumwouP6UIQTy7yFjpeuw02c8
yaYVzMET6aDoeyjCUb1bGXkysnNq5LBV8NLy+C4cVP2s+pTYB/e4m/AXb7lW
AdggIRwt2HWS1Evk/NjtFuBW+9U+JLjDd7Tik5xvt/5+cL+SSnR6sXHib6Zd
9303JHFZUgMPSaLzOuW4iSlncqRA1ZJK8AHm+pb1lcu9L0KmEq8gBbfjTEzb
LKUPIectldbV4MaiPc7XpoBVofjNT+CYS/XMYuO0tpTbtbMOqZe9KgE0Ib5S
DVxRkotBn1ms3Pw1AhKenEZZ9YkQAvNIqDg47Ep1e/Vo0XoaesS5Gb2jkTC1
2rJsDNI3tc0yYc3xKT+NwT04CPa0/2F3xo2x/PfPnUXwlylnkZRrg4DHTppw
LddgvjU0T+X1/Aka7AAMXRKfqfExuZogm/dH3X7SZXq8DgRgD21cP6ZamAK8
TG+OtnAszJtbdNUBrzEJxdKJHxt6XML4vzx5Q6Rg8KZHZZXEjBnpIBjJzJIR
recSRY2pZbVBxnMaSba9rTqUR3gIOs7nrlGTZZEYu1fW+w960yEtgjGI1F4D
iXR1KgDD3Wpv84Q8E//4XL2PQ9Rsm95gOEyGVszb6sP37bckRe7jBHC4s2XZ
+7zUvYLfRBy6oCTYcNK9UyHxSgbTdo4rMeErkxeGCgx7n9eiDco+/moYHnlB
9aSZZolK9Jg+7aWcwBxfAEJfgzcbuihF1dgYs6LxjqFgjghBnYGUtaPeVXDO
qk5LGj4z16UQfwnYff9YdUmPKpV27VIoRaAX7kBGk0znJvuDU7rdR0sT8wWR
2NgM6gctmviCEpyorF46wjUdVbt0g3lGPQTJauRr8Bv9UQqRzSQWjWhOuxUI
GTaW1Cqm3iyP5KDH5f2oSy6SPmZiZoEb9TjukmdFAQ4JcxnczclvozBSkedX
3BbFW7nxEINlFuNs0lJ7oIOV3BEKCAXUz2ILI+gm3fE8tUZntUm2Lkr/Dx32
oJfDJu3BS/L40y51ZwgFCB/Pg/K4o440o+QyXOTLX0GxC+hr+NyyX/RLe2RD
egoHlEBqozvxmiTWHpbxjJCePNgM/8W8thr3Bqdr92L46oAKXoThwDC9GkHL
K69fG6X2m+rRMM+H14uUiCLuFmwdplOVS+HJHQOjCGy7UyGg5lQHJVP8MNuS
fBR2AXqnzoekFA7jN+zyWlrkoHt0tXveib5Cew7i8dLSl0ito+PTxwlmOG9x
BZb+d4S9ai++cNE7QtJERdsUPQdw5EHZPpJJ2ln78KzNUTJzFdkFSAvYqXfC
eHzPqs8R2xcGaHAf7jeu+ovVcvfNV1bLa1tOWxHAVI5pcsdb4sxvg1e7Nh7H
Xv0BQhfhwPJwWxP/MhzqaWvH2ECUVc43eG5go8xLEfZutHimXXL+5vnwpyZr
YqBc/t8nPezI1cO766SFFzSq9pmLK+nRFG+pSpNl9FY2BLab+MzvCy8H9K2o
g6x057as9wUslore5uULNChcD7nkNvER++Z+JmidRJGdPYHzQBazu5i4D0UU
QOVceDvZ5EfsSe8hSWUY6DigTiDYcArIEJy1htdmud7fJnYiik68wVQPTIlY
toVC8zCEqOFp89BIzXJUKHDnP47VnU9H5Z77K2w3zAx3Nhn90ts9cAcVK0vQ
4ePaL/D3kK8Nnfw+SFNupR5Lg1nD24AmsETYgTY2mhkVbvGxpPk6owlIrB4C
ojD7LFTHdnEcHR74go941LhN1P9u37hatN+uiOQsyioPcjY9CmJxxt0cXI4m
AilOvv6CKm68RpuyRRr9lnsc+T/BfbFu02kuipKi2Ijztq9e0PHuE4QnRnD+
JV8nd/CcB7cAmLziZ32kc2+KrqLC3q1K4SiShrsxlKd26HY+/6z0AaQF3CQ+
WADujvJj+m9bHvKPnKzzhUAFVqeZngUOgXhbGxKO8R9BTe9UK4wjXARsaFSY
LEexNAY3Z9n9XaTVOO9cyGtJNwKfoQ6kqaEUqNs6KDVEk5XO4VnmtXuoBVW+
QFKIW0KjilIXuFu3K0WuDn7wYqMQXWZWKB7+V7w/KKbJUZ2NU5Tv7FAfSD7e
jHJdTCaNk+Sk5T3sJCW1+ocqjsK8xDiNJG0PS+N9BmE1YHuitwAiwUL49BxR
yZhvJlip0Z1y8chCyA46D31SWMfVuEm08s65G1sd1qceE5K8fTh+3c2a5Mwe
97Mo+7+uEP9nU7Eu2XiLoO0N+oj+pr6PVgAhO7fvDSttWfe7ppdDeWRoFO58
M/+2Ao8Vdk8YaU6K1jPqec7BV+eT5oBOFGmPe8rouZuj6muZK5CbfCBhOkBZ
KZcX2VCvQ51++rxxuvPEQ7y9lxB8RGG8Mgt6y+3DfbTq1lAqf887aAafO+Wu
BUOE+QBvx/siXl+zvGRnqkjyjQCmf4+gTy73ZONfSv6Ch40UD2SIsJhpkEIL
0Zd7h/BC9lhj+XglGxtqFNe9tE6WdR8UK+BNdFs+cIuFdoBwOpeOtBpBBDih
Y9OS65G7VEowkAsKwawYYCjKTg78KdXYUH4l30igY/GbvM12z5ejDgHFeOmp
1+LNHWR3bvFBVSER72XUh21YFdye5St0IvaHs9MZ4I8ruw0wgxmOeptwM6xt
PeAODiozXHVk/+XBtbrqCF5Vb+nkfyosbpjAHzHQLSUlduvru9E/B3ZnCn0C
s83P498Wg6bvjwDzORnhx/T9dvi2xZBU7xzmSielZLEw1jJtrpzsVoawYjDe
IJ+W5bsIgG241mlIDnNx/MrhzA3GCdWdbuopQccCieeiOpnwJWx0INOxGDqY
AIrz5MxVcDt3EyxHOcnhKgkETSGP/LZKVUEmcSLRdmZb/58Hwmk9UbtS/rfE
u4m6fJ0P1aw/aEYHPj1wmVT9az61Bl5rBdeR8JQGg6OMZp5Ys1FUxlDh8ibw
PwkIaZ6s8/IxWY5PlTkHmjD9mRnwErF5ZBXxpsp+j6KH6n+c8rX1Ot/A5x1K
z3LHFxHBQQRhIdvnusUti9q35fCaWuFUC1WlcYq6XQ38S8WyrrtB6MUTWqMx
vK31ogEJAdQ4DzLAcOgbdfiSKYW3+GynnqPbeJ4nMOpjDLMZ3S9B6YpcgZ7k
3wT9xNsVajwDRdNzSGmJsWzY3SfiwtHAccAKP5oRdi6B5WtNhfPuEY+06ygU
JTbC+PeG7vLa+ANrbeTitUfLLL7GaUi4l0saGkK4meF18xb7Sq9Mz11osjz1
PppZyhrHH4ujjsGN48k8VqhFThJeBNX8NO8SZx7bsDK3qG4eSFB9UUH+/JvI
cbPOjEScpFyoLIdt/IojcplnnqYm9MExBwFsaalhbc65WMfD9pmUhMmd66aI
DqfkYUhVKWUQYoCCIeZVYHFFPBBivio/gLB/ZPqkEYFy+J6wiE54xu8590GE
iNQPYQAx+20Nux/gpsl4ENKXcFo06+Gq1zI6iTp0YhxYlOV0xgcyfdykkhXW
faNDKWLIYxnQFVnp+d8k7TPXWXokXeqgT1b81bhCRf113rqIejdqTpe6VVjS
EXfdbs9ISeLlWx6gKQnsS8b4nAy4qmgCVu5nWA3ZAHOfIt1yc6CCHwcuwugq
n766gLgPwAH8ME+ulHU3UIDa+EaY71yrJyF63EYdJOprRjgA0DBQxwYVEitX
SUCnWzknbw/WEQGwJZJzO9islN6kOzvalkNy646U8tiQzZ2epu+EpOA5Tjpa
eZsaS6IN0vwwe9/hX7N/8ua7wOfqJUbK8yTP3QDBmEZH/iaarwKkRwmFp5+b
jDz66oiDpBVtSTugejFqblvRl5Sqky56swrKo6TMS2QA/u7jN/AZnlvU8fot
AcqlELyNjWTtn/PDSz8XhG7rpJUUGuNAztLCge6CRGzQeRd+zjHDLIBhZL9L
GiGJllqEO9fqjSgn8+uGPZzqTVa4aKlZXPOtMmfO/O4ze337LdvHjWeGOrzJ
t4Xre+5UYcxVzlG2bphwLYie6yhov3OqmSDYDGnxxoh8C5K5y0UAWd0I+B0S
oiGSb+dJm80DyOMVUn5VQweSZkv8FeUlL3a9e+3lR7cwLVMkoMkVvWP9ZChX
3PIQQBCytOMixcNAaMzix/iDeu9k28ev2Xtp2PTsPEhcgszTW1yLRywfpij8
HtYt9WTFNSml8u0nLueRg/2DoRzdOIGNr6TtpIFp9W5ujCjiFYsdkGcbaTIc
A4a27lmbLu9U3NYfSEC/NPAku9fs3UrGltcAyJy5rh3oFkXZPi05jDbalzvV
PENUxHMjTmeh64QRj7sxL54KI6ktvlgK7YgXOfyGovKTZfAeYvcUSyvtdwwE
V2ZIq73FgSA1iKX5iOjldgL9phsCNCud24zS9ydpBcCcMX3+d16IKeGayhjW
H3BJafDowO8O8eS1Q6cUWWDRiyZdP8PxsuRIk2Qmo0Fyo+SJp+NNrlt2xs6/
EJ+O107OizybKvmN55RkERsS4MESXMEGTKMDqToiK1RkTRew+MKtRf7yE51C
Kn3LK21PS0G/XieRHoShe1uypG9bqqGXw8dUcKvPV1cPj4+L+1nS6K9cKqgz
gu69V3vOELNOAjuni8ed73D1fXV0ZzKrZF9ofGv0NRdvcHdqf6NdSvpxae1L
MHF98Vztf2NJospiWn6hDXymP7Ux9nhGSMIqOEKI/THHxWM7o/jHD+YudGg2
bSgSMxqKbepavrvcVwQnwC1drba7Et0WrnDZzJSRCoC5iPrL5ipHu7/Z7jDU
ytwWUoVJ9F5R5I5ydFyh1AnVp//f3E/1dT/vbpCLEb3XznK3fvK51Mi4D0ra
4O6mSpQ7EErPeOf4fFK1AeKwWW+1Ji4gvo2Gz3iptCwjFwwW4CnKt77MNYOX
cqlwQ6Gl5DdLJ/mzkKdoLnRKmAia0EMzNVI1PFxlAMAOJalv8R0SjSSvgz1d
FSuv70p5VTEZDOVS8rHhc2HL36/l+z8xNJVrJ5ou43nHUuaM2YvKirz5vCdL
Hc1G9oywizau/CtiRmcYSXLeb4kflOnozJJBur4DOytARjThnJua9xmHmZDp
gyMOQa7FSoODtxjcPGXtmq9FtrQCp5Zw5hWHCu2LKYlPfLUBbREVGgW6QOWE
bI5GvpP4CCJkeoxfxUOoGEaIHa/muX3EzGbBRi1Fw5qUcu4BtBeu50lvMx8h
chgdqltt40aVA0rbPP/T5Qimyf1NofjlVfEUBZ0uydD+QTmAWlEE//2k/FAe
96GVMnt2dP8JaX3XCg8uTWAARgW+LSHmyo5DPGztitgFMsBqXRJvHcSnd+7j
YJRi5ZVfD4d5qnk789kvQZKgcOGKu43Nm5GOvRLeENoQaQcxkbNRUSRh4EUA
n+M3Lc2ve5aUegWsG43COVado+qt0wDJfgEpjzKwsxuKHTEG0yM5lCzuyzEf
a46pWtjq1doiEzJsIlpvwBfRmWI3krMgYvqsGq1fYkre5kf660oNwY+dlrTs
6incQ4X2oNhbANoQB0KrZB6P20ZFx6pbbjBE8Ff810k9OlGrdqOD+097KfUM
sX/6YZpNQbALG6brG2FpZ8Eakg7+n3Q/zy1OaeOYz6PBdJeJmiGolPUad2Sy
sptxBqLYMrbU4vuWDRujqHJqQ0E4AsWVFM9dUNw6sse78hqFiM91u27QURyH
RMRL+te9Zdqm2RqSvJ0wV76TyhtfTziy9yaCSGku1bCYKVY6yWmzYg4lfjZP
ZM0Y+/1RPyQIzWgSOWP4nXziFIt3RcR7H0igTLG1aAOfgQzookAN/5QbuWRk
TFUd63P/dXXV+I6HikOfJBUl3ZzemruCFcdUvJjtk2JAWR9QvO5nR9fRUDFj
TWCRgT5/3/M68SJX8ZMJMr3s8xJzMomhyTpLM6K4rz2bfISRkeV1vBj0inFx
v4ffiUQCo/wbrXS/EMvXWUu+VT1smBldL6n+plXRd40JP2UnhSshNFjz3Q+i
JDbx5UfF6sQ1TlMBxJ/+KpHtn78G+FB8YxTReSD4f494L0isajmfakcoGw8h
0hsVB7v1kTdArxml1EzDHtx+UtQKmGHZzkQLTQ69g+/wL/AjZrbLiHPklXWH
FxosFf4hLgrqvDtoLr1hC/sS4UGsZuGO/PBHIRvc59XSz1iHx8vDQJpG1eNL
hb6H3dz9UKCyfRJXCFAsdvBwJJuToIDhpYO+62hy6i6k+1jzjYVrW5WRN4qk
gbpfSSSqptGm2XloDseTwvQYgPxDdcsXDEcb9x10pxl/jcg+Vabw8O1Lc79Z
/oSX1Hbxq7WrNRj1G/n2/+2N3Mye6U46V6w6WJe8/mowpSJPWsFsCpZbt7iV
p+MQkgmfiItuo1CvsqN3PTegRvIrafSzyEwxOu+JQpxT0tDVvcixvkHaQ8c9
OO+XJpi1JKiLvaoX+q0qBxQzRcbzPZtBttPcJnZEHs+iYJGmMMyzYVAe3dmF
G7qbkAjmKNW5ibUN+qnnTuc5OYRkUC5viVlns3t7b7vw3qprS02ksGhLGZH8
axyIDlFVqXXlmae1YKbIJ6haFD6nelJvweHJ9MKRRdxL7QZleUsSWyImQObW
edIXZvjnnSVNn37LUp/jRAV+HvinmyewWHDv9Pdt+eTXbcjhbiNuRWg7Gsdf
sm0ImAF3TcT3qBfH/iG2E96C6vHWvbDc+v1Q64I27LX6ZcMxWVJjlJvuGF4L
r7Fa7bVZPJ1jW9f4fhEFY3/X7JHXJJQ0wFwfHOGy9Yiw3WQkMbM3klAOTOYw
334n6CcLkoF6oBb7DdWu2ewjzEcYCUEonb9BG0/kT31Z80G4IR3EDxcoWsot
jU69ysq+uRQB0KF4Tcuhn/xcprBIwLO2V9P7u+X2uoP/hONctRVeoAqHb3eg
xVEaJ528EKFXTCzauCgD2iZ54o5u2HOCIVwRkbfvokhX33VDxOyebDogilVK
bfEMtdpkGN9d6iHJdpbmMk3r8gwly7hvhUuKAmNTs0JITqClNUTbSYbpa+jN
yqicRRmOMQeUhM4wKXKX8Q8c+eXIoMLCrmmv2bAvtrolCHQS47FP49sGXR6L
We8ZNIoPgA0uMpaMg/ok72FFS2o+hf7u4pmrtlch05ZFsvSLzYcNWcIiNjeH
wcOsec8cgdkZa0Lj/HSm0+Zsr/OThVvMym6zSpasvuBV5sLUmdH0NDVKpyDQ
lP+HwOiOq2TozMu/Gv2Wk9OP3+Y1ieeqpq/mCqVhf0aBPqLaRQ/vJaQVozJf
sVdeyLjHEwR4Wsx/uoZeQIhVDYKKhKXNw2M3pcY1WKtV21BHKxDAmZiRrqjI
ZW7k0epXMHPERV0PiLY2/+TAIlI+tB4fD+opawRAxvHgKrT7lvXrLM9kXZGX
eM6PnQ97Y2+RRVk9nmTBCLIzfLQWi8cBOujrSrqo53kv4lTyozer27c96hwp
gtHIrEyLc72uv/wVctN7E87pVofKYGUs4bjLyLdiktEJ+h5kRg0TyHHn6sE3
O1vS/2MCKUujim4UZtYH9wg7/d4GhCkKa2rDyT9BnOQ11pZYil+kf1e6C6rY
qljuL2eo8zX0IACxGjUWmHW8S6ikZmwBvICKoNf5pa5EoEf0iEwRH+ERL3YA
C+V7Suj9WdVh9/O2v7M1psNuyFZ17PC1KX2vtUY4eIa8rk5t+QOhRLCpyYmW
yrZfYkdjiWk8BBRYDYVNpFBaMOwoyIu64XvdMZfFTgJx6H+UzosU5ACa/9cd
1sS7l3FSt+6/11f1S/Q4hTCsOBy12Ba2rOeon1PAn+kEd5horiGsnWK3ohhy
jTlB0QlJny0V+WLFebCvjupriqd/ZzbAbPl4NNYDRqwqAE8juCHRXabgvN2z
vPOBGaIhRZBjv13PRJR6oKAQuVPTVJvP9xLkX3Qmwdz+PvsbrQ8TjV/1ptd0
h4/Y/0dliIl4OHb92bpQoIfmKTVQtD4CNmMAGKnMVa0emwCDlJ3qt89CHmfV
f8OHVQnX3ZpuhpsMVHvT5Bf1bNaV71ye2NmFOdunoA/yRETNyQwXeI2RYfT6
0EmvDddZHSx5yL+mPA0Jgekyk6XK69YoC2BGfaLnZqxTmL0CaMXMv7sq5WUE
4Rof1p975XYbVXYYNRFrX+cvyMQIpJnjvxAkoYzOnHiahdgzKDsj3RMttjDL
wz7imCHw589tSA9NGQg3e+x0CtfHq0SKGemC+XYP5Q8sIsn+EqTjwXPwJN+T
wLx0AbjweE+Mo8lQvDHLkGYJozILGX+5UUmhGoxYfUcI73oPcnGws7NIotnq
i9GyH/jdkbqrw119HAikI9wLLliMzuoRi9vzzDYiLCM2DYhYtMGGabS5jSS6
vfAI6yKQ8U+8ulL+LtuALcuUkE3VxNvjI9KcLcuR/jK8dbiXGfdrq1+xdFc1
vNpOOYAHAYXkAk1Sa0fU2tdRS9bSKsvW0EKYgul1nR71X+SF5KpB6z9rHfII
YmbkL1A0vl61sD8MvbuN78LSuhy8P318axOCAGhJxcGhx+kh8ylvPn8Bd9M8
C2a0UDrGLKmrVLd/Ov9IDGl2ChCOuAdlpLH6f0NnatZV3eLim2zXNBAt4Gt1
omqupYb4yH95wNSkk/g1xBqcB1ruiQfJvYsZAckCsQBUNBNh2mY68p9YXh8m
mwQZ7Mea5P64kLFgb80ip6JFy3EFWHCXKQmyc5NBAhso3DA2cjxUcrU9U6XT
JaBfzsLOgMcm1FeLvW+bPTYpmf0CSRG67Q9L2B1ggL9Frg0U8uFv+0g8eCxn
fsTbXGg3VWHJvmme/eX27+kuRXZ4wws3b451nhRSKf5wCvBw4BjiTjlUh+jH
WXIHrkaoPMjAMHzLhu7D1k2CJyk72sAkv6U6HXxCbOS4b8SlkV7O3wJ7eZqz
lNfQhMVlnYA4uZmY3tYuWqAP9r2xLYxEUJlyogphmcYijQuEYDU9FQbINwUg
uZF7g1hlhTVM4AfkIgoIQhtBim2EN4GjYV3weKMYPHlUjvmBd2gkxrScT243
cJYUC5xUXp9SR4nj7SOzladgeHqpZ10zfkAIiN6EaPPFEd9ozf2w3bwTj5v0
dTvw9xyKSqM1aVGsqt5gQ6nERP1nvv7GEHEcOEo05Nw2GT52iU5Zwte1eRDv
sIXZtqgQDBSFpTytS/cClYd0LE1wW9Y10E6erT5VFHVkeTNX/J2fgjzMv4mM
6icVmh/09wDAt+gfKCEX/l4FuHM3nhYxWVb/d67kgFf77dynlD14N0FBn+jX
rKB5f0TcqEm5VLtE9CXM1QsMQx10uFOfsBtQz5gBH9+cFPpqIhqzo6UBpPxP
2d1bQv//h29fjdxc1QglG69Zy+i/niuPYXpEh/gTl0OiMQNFyFOU31rCl6Xn
d7pq6N69gPH2b8yCn6XDQD06pcceAdRjmYkKHnRcUwV35eogU0Kx890SXP1z
K/16KJ0VGMN4dzD1RBAd+MvGIL5fdLK4UG1xdS8vdoIfiVwAANpdFispwD79
JHKyg9wRbMEUTAQNgemfCirL1OwyFWKRdTLQ2x7Oc3xr5A/oyiQ5b6vQDLxl
c5ogJCj8hxvvEE9X79x/Hw2BEwNn253Fe9KDJUkhGH+cykrvD3uSALlN11mX
3GA+4KJJO968K/gEsF9u1iy9/s9l5u7YZoCTVdc0awo49MIAqAgneJkjFFA6
MWj6woSKgYNkslFNJLesBrzQlLh6yxuvR4Eow1aZ9MpmlPgPIN17Cmd/Y61l
NICXp0fiPmZ7vIRCyKjKxUCEIlp4yL/OcIROEkU9LwaFRX2B3C2KgUQE6ID5
msJ2QfRdITTmZ04Ulvi79++mUgTiG1g/6jMcpQp3z9REa0kcyF0O8MC35kYm
gWYU3CoZb4/N+vAMCDDPfssqCuVzwwOTSAMFhBBNC7IYbk8mpiG1ZZxLoAGB
Z1ItOh7CjBKnNL9nQD/SiOM6h8+Av98KjjPa8t0isQYOMh76RZrxobOgoruS
oTifeAXVPFH4Iug+6kukS1U+qZDKgYyEwoHck7reR1nxJUYOqO8jQO56NqKb
ScG3yBoHfusSgl3XsDdbG8myE6j2oVG49Yg8iRxXHOCcBuQDi44GfSwxIICJ
zMp+rByIz6NAw7E3RYq6d3GJlqaxWzuWnK1KKWO2mDHki8Aw6u9QEYD9iQFk
QIXpO540YXy5zF+qAVKsyWf4WwZsqYgP3ySgAjtzAJ+M49QBU3v2f51gfEMl
ShnKNjp0aUHIhgPuM0L/KnBRZw2tULOKE8CfdYmQligZhF+rg1tbmf30tH+h
Ac/vinShHf2CAa0dV+LrS2xOkcZdmIl7XApU5TRLc7fvsMYZ+IKQDIlTsiV9
zIRwMuGnDckUhCnUuY1KRdODhIDKvB3HNKWY/3geBjPUFiWwh/KuIRfTAgvq
XtvEPoOjnDNueUbBPsRfVQplWzhMGx2igviXZFjYASIQeswsl2Pxx1zWwEbg
cH7c51feQQutOcFI9olsqVlBNR5OXxRdgzBwFWxW4PKVLRR2NPEMvFiMARJu
bExEcGYOyOf2wEmrGV2lo4zyhsgnjl42DqzFkWbU5L1rF948M17QsQtjAVN9
LiijChx8gu+yNW9v2HYzPv9iNuBemMEd/atMPycIP9MQNs6v/1jfV/QCKO0h
Ge1oFfHVq9UXiZslwclTpNjac1VOnQrIdqCxl4OOUIdxkx2fm5pvIj0qHnn6
RpW6VAzq6YCCyYxyiC5qfARScfEPMB009a1rpFHAaHsVyAdDl/s0WGFcrIzs
bJb3L/0SAJRb/rd7TAcT0gRa+YzQKfWbKVYGBLKt1ibOQKUMUo34jRmsS5hh
I7rSwWRL5HF67QP6WyWfBLX2FRs+rUbGvpidCywbXxB3Ll1mwmFGcUTJxASZ
fRQGB1/ihRMkVZcv39OVOygSrfaOe7JAOUwaqxARI+ZDJmJQDxTcdrfEe918
HbufQxbSh1aQ8OZoUlfxAKFxuJr/40N8ad7Fw4vijxd2OS5eaCbZ3ZTIByDl
RXf4Mn1wFjZq9DX2il6TLlmJ8ZcYjBM4XqjVwc8dta726jw3wRK8KsWNzt/O
Qp3a2OV7h2eR9NPgDVC8WDUPvB0fmpeQRiKoVKlFmUINKvhiU6q7c3UC3F0D
PKF1pihE7e9WRNGQN4RT2DUXFsLvcQNj1gPBpZA+h8utQlj1T7sRZIgytF2P
9RcNcImO/X82WFnT6sYTvvJzN/MEsw6UM1g9v5jQcI2YglhCpQVA7VijR4Nm
qOFNBEbPyRsw2FNCFeHhS6EhiY8SwBVwJcHur5XJ8ymvNa0TBI/czqyX9FMf
7ghuLOSYdd9BH8pm+EQ6bn2nd7YG59CRpqXgaKKEVmWB1wcYre0hxVBSbcpO
VyN8+IYYqKpAg7EhpytnxCuvJAWT6yEAuYE1SecubojuhPKFLNguavZ6+cWF
hS7kI173fG3JQjQOb5VmX2b8t8KYZWF/my8XRSsUmuJlzYNMvA9mIHUYfQTg
qxZ1hogbjf4+fhQwcT2uqacwfvtKhuOwzXyV/Ghx6RWwhdrf6wXEUhnQzbmU
DsXEisckXKraIh8wjPG6qQB7bBr9ldFlzIQ9XQHLF5MLtvjVuJExmkwLTYIJ
rHw6169KtDsd9AaNIK1LxdXijqQyE94eDnZPzwtIacOzas9VY5czjoWGbork
oYEZ5SXHfRN/JNYM4t39mWuoKsa0dKSCmCmHHxEsgFZ+8bbh5tGebarP2HDm
xZScBxYaUUPtuZM0SNtfFDCvKObv1671Ikgvn7LXVbtnBYxtZ/dcQ1Ed3Q6C
yOykHGtOq1esSJJ+kCUom4OgAVJn5Es79kq0oYgVLHp81NwQzNAFrpo021ei
Xz3/IUqlklR6Clh6iuInOiG3RiwK2nZWb0sM97CxB+Sv9mAZ6E71nA0l66W5
AzkLlk0GVhw/jLJyjzgVf7irO0X4khcoMNXAimc5CiO0MUJ0Bmc2iWqGspMA
E0Jik2XsoDtjEjW4fvtHg9fnrnerFxX7fyVpfINTFjTuL54BUgvXJp/0ywUr
MEYXiUKHfFNRti2YFDtwq91TVJlChh5HmSvnNfI42uXm06ttE1vg4a2prZbI
jEl3B8bFfsI6gpsqDqytvPiZCPN3XVtvZYErXJQdYFR/8M14tw1JqLE27kPs
0XnYUlFBfOLkYNt7YnVGXIMZcd5TBqDCfTqgo/aOUFOGJQP2LSiAtBP8nZKm
IuiFDvxzGyGoZVw4XmFNk58BATGpFq0/ITqWIeA4rHy7M4hT0ttf9VOv7pMa
uuHN8+rRqt9a9EIMpLHkbEETZmBQQM1WMeXLiWmWxmhI+ALaf73T3CnRujdL
F3vJnQM8TyndPc1elZWdq7jgGTa7Z674M1SaMd9guw6q1ej/Okg8fwGIU8EA
/+PhH7s3AoDsoxdBBpdJmaH84lnQmmAy1VKSYpE5mC3U2THmBUiYAcN3k0YK
l0hfF0GNw5xRxdC4R1eRfyXxVylte6/32t6vg4OxjIQtyyOc6qXV4Z9iDH1K
PgJUFGeiBNzCg+pvSm4BN9FTGIx/xyMHMQVDWn4liKxG3XqTuJDiLPInRXD3
A4J+sq4ev787I/BfTjm5xB3hIAJg/wNS8R0g9lFkuXU/esVDU7J93Fcqcc+f
bRwPeVYrkY0eSZggs5TGBDsurWQFyXVih42M5UfxRIZEEQ36zHdlcd4/qDyI
vBdKNJBdjHaFs/c95Al9IbjylEM3vEg10U/iQFk0Hpv0k3d9zd0NySVE2e2w
nVqem/xX5Nr6iKEil2P61bFcmTJ7wvh958sGhXBRiHU+6rGoM2vT9bfe6gVv
mtKhGpL7V12XlWw/Zy6iB5uPo0hUvsCKRUmsP0GoAy6LgxnWI8+EBzRf02lE
DQ9/exEl37mDTnwKueFnP71ukkW9Ggd5jqQ9s1UOZJnclMyRLCepNRf94ReC
t7+7IJD8eWuuC8xzHwwl+0m+JiJVhYFY2NzYuX+9R+BeMNq557KsQA/7Ener
irc8ygs+6KKln0D2w9DFuSizzR1R+Bw8AwfUF9fuC6hJGxuLd3z7r886Iw/f
CGrRsLwPa3R4Hko824bQtHRG3JpmC0wTlKYBFZahC3KSJ6NthrlLqjsF7EI3
g+2W2wlqHLU82IxT1jezNpWQ7YZ6mkym9GFFuT2GGob7PmVmSbZQ4DzNu0+5
r8BJm94KuJuTj/i/OVtQPc8xwREkoVLgS0QrN1zHyExV0//GGce89zCBnNN9
n0OmpGBde9X1xq5dVgd15w5sRSH9uL5+NGQr1buG0UTovvDDBZB9RrArydSv
v/NPBOkxTxSDE0aC96yKmrbSZF2WyBeRloOZwrx/8uIWC+RqjyihBb6DJPpp
M67H3wCMwNIaIjLgoCNasqUENSb+uPD/g6SkgjesarilovZD7ib1fMF5tKWg
STe7ebgvdP2az5gFp1Ls8FBuB2Fz7FFSQECkrmUiOyXZz9hm9PPE6iOsZUfo
Vsyd5Cm/1fgmzGpyoaZ+cOA5R0esAw6nkuqpIcZFGTbFGTBzY5eMycBd+xc2
wDmxelClb56dx224wWiD+yrdOBwbrRbZn8unucnwWLbI2ymzbDb/6jyhG6BQ
RsKwOrrxCiuwFt3hxHs7PPsZZhvPD3bk/nDECNXKrm/+woGw8qdq4WzAXUo7
0IhxOqNVNzTbcr0A47KfU1BYJds9gP68iKvUcKZzmgwQZgta9UXFsTjsRLPw
ooC5s+XlyPCXhbzowvBMkCZ1owk5lpyPYazIBay5eotxS05GJjqfHVkmn/+4
nbjMx9Wnd42g2Ggejib02KVb7Cgcy8wsvdXMUlm2VA6TZ5lRlLTfu2L/UKFY
CELxeLXleC8zU4nP0wmKa6pyfxORGygnJOKPNHNxLnD9GMmx/G1D2GiElJLf
oqGPtkQZku5LNClex9fwZEQ2DB6kimgmIj1CcDWkYTSt5HYIgdDFVYDF7znd
XppgOSFzpfDL+3EvrU/Jhdq7A64CcOmngY7x56eoLn5HIUJmOuTVDjl/bRTk
aDMkVp80Rnx/u4Xu1Yij7jNyNnMG6oLLOGjxGpEAfwAdHimCiMWVZU7nO539
yl40Nd6KqQvaZoERdUJpKu96JLuw12JicKhq9ISZ3gt9mwmXsHt3tSoecVNx
9I5ergA5pftQSFLJhbMEAEldL6qTXwuOdGiCBp00sa5w+Y8QCxbW9rUvMMNY
K6RU0J6Vkfiob24/WLnlO2hqStRilCLZEWeCLnmeE+z6VpLp2Lhptz8Fsp4D
uyohPNhNrY0iraU8BVyHkzsUHdMJpyuFb9lf7W56rMm0+/1+oXKYZyCZmQYz
y5tcyj63Fr7iQTkuOCcxHJKA18u5Pq0sutzv9jMhxdFVHlid6v+ohp3JDqym
3kBRxK/ZgN2kPeINl8cUZcqf3NcvZ4yVdJgWFhf5QX47pcKFJdxfulFTt1Ev
3PqEZa2lIkAQzmKOlSN3ubUOJ2yHnUcCCLGRoKItv1826X4qYQ8HO1tLLzgL
gSkdaKmFI/ibyH2lqkEVJjqnmfaqp62Ywr7VJGEHvDyTx7tqlgx9Cw/LVhwh
e1zrI5WTQT8QGjmzGoWDqSuQVfen8+XEl/Jk8CtwEIpKQPC3MV4aFK/gAAdH
3KMlkJNmsUHNeEDh1RDZBJ3rHmyFz70ov1hDCHy2ZA9DGI8kLWmnYLNyQMsZ
nJlHwcEnNBNJ2uuf2/OzJCOtV8z3GzjkF44wVnCXzysJ1bmQBDrdsp3pUBvt
Sfx1s/u1s1RQlnB2FPzScMbDa+6MRKEbpbksYVZ+EJzAWzUeVTOJEuspPu1Y
9CKB+lvW2ZLghcHXzDLYqpJD1lhHZOE88dtPqvUuhOl6+zzDRwXr664VFb89
kPH4JZ6HOCrjoRNiyBjm4pxRrvJoQ4LtRn+ts6v8fiFa8nP3hDRfHdbUjpgE
6pefp8LyTFqSuhzrsyrW99PMN0ooG1h6NNm8pD9q6Fnk0gE2rcEGxyOj1jtA
DFGKVed47ko27WUiOUNN3E81o687mZ2jClaeI3n2Y7ihMM27DMo3nXHHU0VI
xqilL/1EKNS+hEVprw+u8l2gc01oUCdKL7PDsUz8In0STLjEZMBQORcObh5F
PvbnDLgT3KAgFHWrGBbbDMlXQ7+EsKgLj8cejibj75OVGqeKGuWGv7gOIvgb
CD/MxjTkWpjydpJHr1kEhNb8+s94FWWbUT0WmSuvvuscLIPdm355euFBwRy4
qeWk56cfMrOxEw7q0d+xHTZu1Nn6kYiWu5JxpcunGPwe2zgLVdIzC2t9BAGc
1znjU4dJqJ03g2U1N4yrThS24wtJwFcKFdobKDGFM+zY3gBZNjM4WVWemH3i
qAEM/Ldgd6NxC3WoGaV8iUYUm0+4b92WTfhrMMXrRa4POoif+LJNIVD9tnhQ
uNw1mYXeWt7c51qE/nexNYZUxo3aNbPVFjB8NGD9mcTJipONaiVme8G63RRL
NMBsF69ScBuej5vASwkQVt/scNOpeh+eDR/B3lNJ/iagHiRRxibG2qjMUivx
wuUG99UpvP5NzaCc/prnWw+5JkCF9HtK57vQyaP4M9lhvE+hkgz9TCAs6LOc
J6+Hc7Qfys0irMkHICU+8Xu9iwsDYPVcOykWlFpTeONL3tZ5/DjgrYDrCyG8
5bZ5C96bBHFEXMDCzxcwlIlOe3Ma7WWczJAJxkEikSsZdfosbtqCqpRrGDu4
KkABnHRB+ROgIcccpo3HPCl5lY3v/7Q/SZvJekL057OMIO9COMnBh/SFmHJm
ET2dV/XRxUjgIOxMRd+Et/gXt8BKnoJosfq2DmRwCxalOKWDH6tqR61HqUxY
48h28We//GlHejZvjzpu5zf5o7u6ZcZ1VxbrQbv1pRpuSI/FEqmKqCPNz8dW
Ll3PUfZBwk4zIt11881iknLjXc4e/fr9szBy3MVbsWwm/5hxGCQpQKCuJ1e3
e6zYbd5PFKLy9YN2kF1THwsLa6w+rebkECj1JuVYtAlw6HmrA++PLXSIA1Mg
HuiSrs2WRmyL9xkRVRt3obg+OuWxhJS5OtOdd1LlZRiWmHHXQCEBnla2h2AP
S5V5h5s2Oqb3K7KUeo9DdztAo9GOMHN52zqqKSFg/bhneWKnDws73vVaV5H6
J5Il4zOhFNqQcB7thG6uFfHoF11UI4Yr1MKiRQY4CubY77xNTuAyYiiS40bV
s8Oj9qIO9f+M9KnumVc3mFODjNVnj59abJf2ZqLI15Xm2tnOuugxAT6TmUbS
hcezfeW2EpDsQvoY/g66/2+iuQVaGtOAmUYlAE2lLf3Y+kh9/8OHK7fCAS96
89oYoGicH9+GseEMuvMuH20OMdZgMjKX1bSRXC014Cgi/QCqELLJs8AYCJXi
LtTv6YTG7CM50X0ulXhbCUq8uOWLB3TzbYHt20uRUjJxPck/K67tJGaV+y9Q
YVL8CYbsEo9ruXscf/xRZUGNFIajLI+X/VkzLw4+e5HCJKII7UTsGDOt70kX
ffhayIYEKVJEgjVKkmKkBiv0iYnkV6+21YhJR/XXIWMJMgbe0e4Fv5M+2gzA
B3/FWvl6DXV0f2ZlEBxq8oSHDaiE4ziYYyyNq3yhtTApeLyw3eSA+bzXyil1
cMZEHEJwwJjuohT8N7HCy+go70KQ6IPEKiU4APExNgdPSZjH9R8odeLfB2tP
3Tq/VPqyxyUszdW4F4FoOsBf5q2vJKtrnLDpSJgl+MmurQCpNyklkVswQppM
/HezbHa1bSXyx64N6Oe8tYKI7LElDXAM4J8D60AEbjloefwioQ+WUR/sWHl5
kz7fAds/BUhX7mi/+lEhRO6UdU095GbTuvTY/8VzPWzhMFQ4Q4pTW+Lkb9j4
IVKH8EiM5CwH2Xd4BsSo+XWoTvMDE+ll9+cQ/Jy7bZI4PPZ3hy5E/dlg82xV
QiAaBBt/F1V/hOYNZq+UtvZF1jBDHrxpcj6jvfQt+XJKbcchMRGc7a5bTgjM
Z7JkqtArLSN5Bq/VbXnjNBCIgWLHyutinQnBoW9N4t5Y6lUi2mvRN3idAlzT
kbGniTdVr2h1+xowiZdkUHna+GHDHcZkgCB28WXwpe8C06eDAyWoyq5N/p0s
pT+7Lgfd4gux7uXTej+D7hJnf1ojnsFY4B4t0gQj9kPCp/RrNywGlRBzx3rS
nvZruBjqmO5eIrOOivcb82vCzMIatytpHgYCYzgfkG/kWFp2xLRXG+8FGosh
aeHnfA2W8DKzslQ1epZhvctD5FguF2PloXGsQb+5BJiGDMMRGRHhLIfBL4C0
lgvs6k4qCn3lygXI1BmuzKHyBOiCHUIbD9j6NnOxl5V1qslG3c1Wg3As5I5G
1fX6SyJf4SP5VhFeW3LV7cd5wXz3MaRHDBjVYm1w+i2O+5jGEDMjFyjOV/tA
43yHIz0tpRShC3ko6C7og8k0JB4JsdCZ9F5t1PwgY2SjR6CiRU8vlIb/3YAh
cuH32ZwoBamWegqNPlXgZETyxLm1w/EV6TZlKQk1VEQYqsTVyRPSD1ZrQKRH
RymG/NBYZvik5l5aPcK8PzJIFU8MyESGDRn6wgmTzPGadp4fHz3/HIxaGhI4
WZxfra0MpgBsT8xHJZIhdKKPXAahL2Pz5LpG4IfQbCvOXTNeWbynavpcbVKm
o6g1FgnTXSH7nHpa1JrVoRQ9L6N+08pwnav9ByPhjXuvezxRvPDTLYG8gbhe
XaxWKVMOkv8h0Nn/lI2DfBMAL0DJTTooOkBn3cvj7YqEqP51bH3PQ0ky/29v
N78NosuIbhO4Ssqc5wV0UYvl5wxFANJRFZCqT6nkPXsqALIHoiFK1JiQMV0Y
i1eWdaKgonQpjx9iWItzy0aPVirtY7PoULbZEv6v3up+CC81a5JzpMoo4Wa4
9FmyXW5bdLTa5IKuvFaefn9sxSok85OKfU4sMWdiNg7v6FhYeXmShSQWeuGV
mTyr8TF1HW0Q7iA/kWoui5jpZGc2uq+I+Z009wKqoOWvPJWJ/25O+I/1yXRx
3waHBW2WNmPjaTsDYAxqIZkrxl7gwArb8vyxoyNFJLnPqnAnVLoucEx5dWzp
YlOBjwUX2mCS+fNe1V91hePQuY5AAb7DC92z0hmG0VRHF4bEDnXziCDk5BmF
8OCzOIGWSBofEfxZSSwINcYLwzrVIxshW+AGWyZicOMhXownHzoNvBrPKPZ1
eWihq2j6u0IEXmuBCVTzs4NzPmOfvZSjrMqmMdXTfO11d72YRBLbVFu+7VRj
JHxQ0x6vGr3aP7/CXUarSic96F4oiUmgPz8Zv0pnq9Gh/KSXHWqeug5yeanY
9SqyfU0VWmrIBlATRPXAYpJCfpBNBB5FSU7uC0pxlP0fI5auCJqza53AmMDx
a/PiLV1WMQc3rX/XUsCLN5vm4jDJU0IRDfj+ylnf9iSmY2ez6fOIBNPsAx45
1ukRo8/4HgDZfZVAcPAyF/umj2gjm54k0lIUsKFESKNy9Kz2nCFrX1wJdAlr
bXGwWkzPYSBi7gWuonyRUThnft2QGMyj8ojAIbvpdpfgj4/3YJZqSgIBBHRR
BSLZHV+5I8L/8K9xBgEqRVWs+MsnTGv1ES4wuzFNTSNVRFsgUYHF9lsZAJlC
h8dI2Z4dHIMQxTjJ0DgolbACUTxm0SGYeRZnagPcO0Ar448qhdzdPT19SKiL
6dbvk4X33biB8cbpuY+uK0oG0YkM1SNfyYFPIkw9auudbQD4p08AXtqCZYO2
W966fo0SGghRNgLXuuoB8VcNwAMm73XoM4mtuLEzdH9WS0kg9cc8j73I8lEj
cYSu2TyrGjDfyWUXprwj7g8UVobCBJh+LzzE48clwasvOZTojx4YHdBPw5tW
9BRVes60ZfBZAPKWWW+K10j3t7VzVBVEF5JG7qwFqkepXRNUgIFTltlak0qw
Z8EBCf1yIQTS9pVST4hO/WUHubLosM+1nQUeBGoqw0gXtuQPP7kQGlFjm1eU
9tWn9Xdhc6qggZ+5mwC0rDpI0wXKE87p7N7AdB1x3WuXGFglpfdrVV85Fi4A
mYsk6BEf0TtPr6HE1otdcJ8z+ipVAofKQ7NH7STyBAe74qjWPsMYJiOCb7OO
dxoVKHhCjvslHEvsGI83Llwu1iNa0YRfPv+WAWA2M+ECQDf2mN13c5AkLOJv
a1v4vCl73jGIFX0M9H2q7bsZ6YBXKn0G2rAK+z3bJ1dDhz88fS3JMuSKDgZq
J5metUt2e7Xa2LmRrirnMMVzNWKcSzj5QJ7OG278OsPBnLybbMAHgmsQD3eG
1ojq1KJpoGqM95Zml7tRoYNz8dVwgUidAySY3Bu3CsfKJspkzGIIlTmxZVj3
1Ah+0Mfrf2lU4jc+IfwzOpuKu2ulfmKTIJ5MTgMmTtfZZ7rUyr4GclikMEAp
wdg1JoGCLRsKd08X4TfrXpclysQ/yruFhRGArrxT973jKVfDsBGpd5wWqmhO
hk74WgEpg1PXrS1uPTlTYObErYjVyHcHMQlZHXxRA3kNsdbOlTTlgDLOJ9Dl
2ns+/IU/hEOiY7aJ9RVyUFBmi4S+oauljVfRPnHKwX7IvhakVgJ1DPyBWp6X
yJ3JAgyAmouHqNBWNJ/fxjaTm57Lp423cWOuz0bIlJ/RAJZdgeeu7Q1fnVcu
u/asBU6eFyKVoTKeZyVgKlU2RLVozQ8zGX1LNZiR8gb1/xMUXsjoEpKz+hpp
MRRcDACOh/dvWL/KRsT9rVT4G5c2iXt7/AchjfwKGkctwlTh8dYez03rUoYT
UUnALWjAc2kvvFdj5dPPyFfHecd8BXP/6NHmlnrWCs6c+Ma+0YEokLFqHFOM
0+r37Ttaepj+JDNrwiA9fepqBDHU9RFXGZ64LGmwXQ3i+yiTgw3QOcq4TRt0
CZjGQTjDLoSmauWWbsI3/7E1QbxRRoS2hHBOkeL8jMgjXvJ8quN5COcBONyF
efq6cDHE08MY+t0MM+0IBSrQzIrXLLo627XNRG1xmdXRVEqvQk3WwglE2+RW
9qtUEDPew/ZsLwavOe73TBG9QPwYbvEwCwpJEvHmFSZgblJYtUMB9hFJXljx
UQY9xA1YrK69qeYVERbAeWohYOwJwHSI0zlRhKrVRNGHptwj/nZOqEIU28Q/
UijULbZdRmHrrfRpOKSbg8f7wd4SQ6Bwa8ym833GBAze8y6Kl57zEQZWXurR
9aHVVx1cOK4sq1Lin+FFx27mAlyCL60IebvNANbYT7c5dmrj4vxl4i2Xx24X
VYWd2ywDuZJr5brxp1jqln27LSmoyKmmKIszbSpBjFpH69xD8uIRy/t4mUNN
SL4lW772XNOoN1N+mjnGL2W1uplg7rUhVVygfPNINgrXnSKmlVcN+nlkAWpb
esbqtaRRhqRcimV+nTG6gW0kjP40eOAyVvzxVodPXCYb/JtPbuuqMdyD4F4h
8GPRKhsXchicJRffATZ7pQ4GKMrvBi8nUBgKFgTloBDLoZ3JH1wCze4ZvJff
VfdX3+0PkFKnayyQNHrhW5nJt79076cKfgmqhFLQfPE2ACmtTE1ChfDLSPSg
zTjGPI5OAVOZkhzQbQo30cVcmWeRRMCpBVcwadMRV/I90bu9oclsGtHSwlTe
2M6QP2hWhD3JUl4QSUz90TwZbcw6GwugZqSXXl2vrsVS05znT6VXdDddhyHf
rElBEPGy63D0ezMrYayiPOuubx4nLlSrhdnSSvOUoFWB+w5YqYDUuIMGaCyt
WQfLoKGzFw/S9g/x3xLkRHeLG7JxH9HXQpTGgcHZvca9W6u+yjc76uZB1Qmj
FEjS1YubqcufnFjMjJhuJFQKxPCr0VMhooHfsR9QEDWBBg5XTxK9Mo4XUKXp
GxxsWs73eUz+VB45cuKnLFL/Bsua5My1eMJ+DbtCGfFTsB35Wc6yblMwsPBJ
0z1FUH1fnNWJS6aK1T3GftL/qA5EP/0CcJzPWE7Dxy8S8ZNmbmLkcmpqOU8K
RqA7V72ZSrsea7b9PFNUnYoWBJZ32OJMT+inXk1rkskOPsx/GVTi0Hk/ihba
FDDJtRlgMK63GhxLOA8N4DZBQ5x49q+cdNpLarfBx9BoEJNcgYXDJeLkAoCu
i9Us5kxCFpNWdAxNgM94XsGVUGI5FtgwsT5XU5pQf2+pgFjpLZivwzjJoSqc
rJcbg5kEOSdMaFrwLHXKURJ7yAvVJDWPaGg4B4+T/pKudoh6KrEHUReqzzQK
Fux2wLm7TwnO7/Mu2qDFcqCzVZey6C1bW+oZ05jrcMP09eXaRVZZiaxEUxJb
NFEVFxXw04SmDXjZ0BfkcNev92hiqvdULfgr9EOsY9z9aoLQ6/5pjtOXVA1C
5SXiBJhjNiircMkhgnYsuDD0LkrzLhBAyZ3DIArBmmDGkZbqi3MUabR5umZo
LMlFn6lU7gAJi2FzYNBw0adEhMxYwAIno4b6AwYsYUOqxauXyQ+igFrW/R/P
8vL5oWyMel22wibz20fOZ2GuINNW/TWFpvI1lEZlJp9x4XAiBj19Ba28ZUk+
nPk3XUNsR6d3bM3GDpQt28NForNcwb3oBc/aF2DZETylt9GyZO3KU9XEoY8k
6l7443Z89iXGBIMEsmrrAkV4CFAF25y9Pe2UV0/VUMbKM+t33r36mDl5FRmP
CU8LFkZVrSx/q8C30jNKZSErxyoBjyPuO07+XL55xWz1aORr8NlmRHI9ng5r
tUmqwqRTZffFwmeTQgdpGyFU+pSH1fqizYiu0ZJPJNGVQb79J4vD8lA2mdVG
PkN04GWq74AhyUouT2NUThAX9H0P80u7wLkqiKwdOGh0YjxaQPVKEO+spBSA
C6p/bxsSCnQV7ns7tGN/vherrNGOaGF7Yy7qI/kYUQtmR9qnJV5/WAsaYOP3
6sEprOGiKvy8tUAdRRVJze0YISOQFLbbRcTogH3Vv/Vti5L1BNG8JK0po2MO
zTon2ItTNugNFNPXxSFG03O8m5KmRGRWBPV8JAs55Q6wvLUIfJi2sAEVG8uU
WhAscEVQrhNtZBIlYnrVNrykV+37Vbkw4rh+fmsI95FhK8IfafiNCEp/ZjXE
FZ/6CNi95kyerTgdUcI1QxsBS8wDXhzEfRRLIuc88R7HbNOlvzsHXAscdze5
Frqq8c/HQvQUyUkH6mVHXhEcbcEvBfD4roIEeVol/1A/todTH8Cjm/P5Yukw
aAIX7QJL/LKXHSo3PxnbWgcpakJVY7jiU8P3ovEiQU3GguUo1FIeg25ErzHI
d7wVwZIbjfx7ZlgouawEuZscn/jiy4ky/yHFSlgPqO0RfQ1CxGfKvr8rkYnF
T+D9DVhCuCAzeE0M0tWeK8Q2kh1J14P32nHYEBpp+O4FMuFXjYuNHC5CncbQ
4IljyV8eStifZpBjmM9eLUlc9nGJ7zZVa9YuODHNX6IMWH1qO7U5quv4dL8x
MxZYXkJqpHbtRVmwtRJgjm3s1xw7ETNpwKrRB9WhgHaxXv/xJTlTFesIqmR1
bKWinmL3M3oLHeEn1JzAjMpPS6qVgDyMT/wuznD+3HZDdixCUiRtvlkV+7Ir
YZvQDxB21N8iW5ueTWHSEb0uekmO9gCnzIOnukzyhWtbyDdXVb90u9AyuwZy
hMNqHJBe0xqpJfOeWaHimgwAfIgErja0MmziUU8J+u0aQLAxDZIFSjj/3wzR
bIdlA//F14ofPuPzqJ2aemqyFXij9V0e58Prn58KLV1DeI/Jouq4nkSg8d7X
UnLmIf5tV8oXvpgJq5N8kLi4i4YyMcSRLHMCZVau792TPJXMkvivuzRdeO69
5R4KOCCD1YM17tJCdXIBnzUCrwQ3nuzOBm4mpKzUsF69pVVGEbAvS35Y5JiC
IgXV8nKsfb2sa/oV7Ha+dTwFsA5SaySLwLwlD8R1t1SOCkOGVqSaz18jCUfc
LrX3mBjZAiDAfhHb49ZhdVgZbXsyaQdI6lWEAviOsrC6AaEWZRb65DsbS8/y
Ay8YK+19I7V3bap5vfWBBZUfBzuGeXWlJCw091b97ZpY6k8gsNRlCj1WjTLQ
PJ7VmcZXHQQSASlWiuLHx1oBQ2N0O5YYYSyHAae+ZZ4sPc9Fc7u06PU0lnNI
bj35twbjvgNJOeVDL3i7K307V6maNWGukoZqllXeAjvyXTyFMn4nbDgOH5LE
/4O2oTrurNjdo22ptoBWByQvSwEorHFxj+C2n3E71gstGcEUoRTKM/DZrcbN
9OTnMgDIKP01STLBV88HV8YnNt2nhH4SyHVIRFcmbJWAd3i8iim2AfagR0le
fUae7Po3ligZX5F9FOVXrdUzSgnFL5sx8aUtpfe1ltWO5tOudej8sfkiDv6+
kuq+hZqlbR4FIMrxo3WTc/3fR8nASakAhiZg3aFOwxBc/zYmJJsYavqK9bZ6
D5IrKDnC2jYY29UtZXdoVBbEehq0Ra9d/bjbKzQ2sV8DFXsYDGn1mURRDGRk
x0KUNriAGkTLt+J4Bmr6nJnTZwniMuoBxgmCGMoZSXlbCduv+uSZMPH8hFRi
2pr2N4NUwBwexIPvaiSXEo9WLAZf7yUDDNZ8SBuAwJMXcq4Y9AZg1mpgTrUH
ImKMs6zGuq34aQltFX+Ixq50tITlKq/eeQ+N7/SYtIDJ0x3D8TT6KRTFi6Id
UD5lCemypV6vnfdTSeU4q/WXK6M10cxogUB2BtkWIlWAAHe576B4WfYrw18y
3flT/Po7vrNlRfZD0WR2frApXF69jUYW1BDjndFH/wfa1P/eqo2FaZXp4IEh
QmAxcb5d6raLQHpcF9NAnrfQDhLAtNZVUwGvMLk1p4Y0hAhq9PP1I9niU8wR
ILr3ybwL22Gxvpark5Tef9DFlpITTdT5invRM89tZY2UCbcxf/YPA6d2tgFZ
mBR/+T/hRHalFLX9bnXm0dsd3XsLZNZRu3tCDZPNNauY2691HwHZf4iFlzIY
t1iAGx+JSWP0cAEsA/8KA3pQ/mUNTQrbcRVZyIdgtiK/+Rymdt7gihCQVWEt
rMd7JOHZNjCLxe94S8s5sSZvdwcy69wxRDC5+FLiQRitvJsTDorrof0l5Fuk
5p2tbZ01HGAu+Sv/b6RNEPyHyZVR5GnxId6efRlfGrydW93UwSYNXmjNLloo
gzSd5lV9BKKmtLAGG6dsshMiPFQfVCTJskGUiDrRRpXywozYgdCRyV+9zaPe
E5/76YuRpasQvTfYWYdwI0Ehve76U9BUNtXMvnvMHCWhK+4dzpArAe9FePN5
gkV93udoo/GyxKsiI3W+Ede00DEQ0BnnsnvXlN1/nan5t/wOaKq4F0nxydc2
NDBS8yVUKsLHiJo4bjhAf0Xjzwf/Y0C2DPJKKFfO6zwpnCy6lvGLDeN3F7SF
al7kPOToVNRg+OklU8rzZZa2vDO7leYj3FBQISq1xTD2o1+XZG8ffnYkA90X
dzHAtub9AQz1dMDgWcxVNkwYfLVL6XqG0gNkB9iKGA81JVm/UT+SvHFrE+2G
AWwlHcyM8zI+QzJr1K9ZG/UzR7qF6RlSF5AB5tbDcrV4IZPwY3JZZMTMHcAz
XWVyw4GuxiQkQviB8oKod4026QmtAePierEQXOHtnLe9JLNZHtvrFM3rHAUa
l5OKXgfPGrOuGexo4t1sNYaebKgquMcPwIiagu66IMhkY4JBKbqKm+yyXVJ7
KLjtTCIaWcvFcXC2HMiDgLqbk4pFNfGpVdndEzTYsmnQ5sF55jsY94sJL1Uo
vOsFe42NdRDauBB8Xvx1rq8I6GhDc+3YyPru80WkEiFcfM2Mw+VCehLzew2p
KggnYDXj4Rj6JDNNjWaOIPy1cib091QZJsu0YgHTYvKiUtvAulf78xQnqtqS
N2bubfn+1Ujcx2iHChaZt8L/KHP/vh/DOLo3DSQRcaoW6aISSn9GyMPrZE/2
g2rWrPFeRX0Vu4+/gUfGla8nOHqr6Wfk0tN7xvrk2SATt9LNfw/VuTW9DV+J
p1rwgh++7a8M8Ew2h+GYdD3IMnbq7RSQNDZ7yd43EpxwGVM3RqTmFgnKdYnQ
9oaE+DuMLyGoIAudohsfATmho9iL8fWWMOWrggkdoMduC2UNyLyww5P6Dfpd
D9hoQtsMqxLU040mlNXpVOw0CLoZyqNYh/ZLVHjXJ7azCe11Q7juJkLgriYy
WrtezxipeD1l0fmDbuqbX15xg+J0erukbj8DXcP0QguHHgrdnG7/cKbdPKVa
u1Ain4cTCzFaxXlyy450qLZG75IcyNn5ZaogqNX/OK0lgYWnGmBli09TSZa7
RswyaHSEA0AP6HTepIYqhUZefCBHJWvk/FRVoUKIMXX0tS1ib/L5g9fAUCXV
C7wdZAeXNRApljeAUDC/ISC9x+O96PAJ6ZJxHhZMERBI+rdD4678u4V8l+No
YAHJda1w97v4o3/dj4tYx+FD9E5gQ9P8jxOuzlm/IJ9Fb9+m86fFtDmt+UuM
tpvmTs55/3lhmUrfsr0clfCgl2aaKFXqrxwUGbA5/rOnRX7m1POu32Cg/PDz
1PM48XE1TMWqlXRBhmoTK91UyNlP7HBW27CrQAPNSmOuE4igr56iFgc+HdzS
WTk+PJ5fPuh70p7BmZIZaxZF7R6tw+nkHwG7SsnXZOatO3mKkfNCSkY7chv7
EKBFfi3/SQ0nb8cK4ehJ7VHXeEHlemKX0nOrr6XwviJUaDVtv+7Ae8lgmb9X
Rjs27y+L8oJ7OE+6dAP1UTv12uPqoxskRajQH1BYixiYwtX78RKF0e/acXuM
nFhWpdtUnAjB6Ojh/hYcQyqnEgRbcnUM6qqIQF++2Oq7x+tHxqVSMs8/xA9d
eXm/5PbJg+iJ7T7U/UlyvVxA9IqUYGuw9KNroeUWycs6/Sz0BSqFaBPJASXU
p+2KGoqNF4rIa3Pv2ZRSG5aIt21fQ/U/lsGiwygyuDXRpCZ5pVwpPf9g7qoJ
iCGDBFCCeEjLCATz6mXvvAhPSJjS/4qIgC+so4EOnPfcyU/t+zjX30Q9/h00
jP6j7rvBQpk3UCslFxMDvse9OZWkDgsGR58+GbtonBm7eEilOqRSTMMONTcw
aoxvv7Y5Ce6Fip/wSUPhgaLKgOCEAEYHTnbCfaOZKW3DiPyguGDCiKoNdAtQ
nVCWqq4L+hLQ0IHsvTmfnr16yxdp0vBiEugij3uq55inFaTFPyoPmSNaMjm+
OYlYh3VctdkH5bQH1k+jeoQoahd2n3Ebpl4lwOLHzQN/fTWshx1+C5+39+II
h/GzjfA22YxqebIGkZiwX5exLOdeZk2eJGyon4OAQ81IZ9Ft0x0eCDvEm0gv
gZXqpnMsPHgTnaOY8UHc6fcBcE5Odi/QL62Sma4d+CU21CV6IU3TUz9fBlZM
MvTX856Aoc2fAjEVWGZRmm8//zjriEfHbG7HDOwvXa8kYoJBFQzlt02g7p5I
JB4ucOZlUGput2Km1MuRipcfOj5ga84qGV4KYwDcnQYo2yaoN829rInQdPPA
3C+x3QfuYtk4UTPJU2coXQyU0d7LAPPij1LAOYXm6YxiBB2sEM753xOTIlXK
VKZdlicjoynuyvj/CqT5gTOI4Xs4WszlsI7KT8kL5N9aUSiQERBkk9rIpXXt
BZ3uoJZQ34YyHCrwE9ZOY8elYCNMZd1ODtz8IayseesriKtoXoBOWdAb0Fie
rF/z+c2vMukS3LalJySM/0biBs8OEs91Q8Ev4Cz0pUfItCIoooCyPWYwyIG+
3sHc2j3RSK4CmgCpMoDJHNttUE8sM3oGssjutli1OwWY09p9RkDIwS0DRUHt
ec5y7et94hLazMyhpurTzsSVfinE8+GJoMFSIwvEIB9+FfZ2v2ST3bF+GPkq
3SyCcAKJe+qIfaFSBK6yTQkG38QTDRxT3PIclN/QvTs57qUTqpidj6eah6Tk
Z2zUpSvDwmQJaX/QCwNy0OlDl/swlb/uWKbuwVHfrOx6Fw4SSXapbrJdhIiu
oGjT5GX2ZMHa099esGY0lJoWUQz0/nQBh+HoWfHX49bDq4tj1ucmG7DjR8gg
sEH42knQUHl6ikvik+fMEuzR21redDpR53T3K/Q1stQqJu/bJ4pDf2+yII4u
zNOE2vQPURb7JOIuGA29duqqbleCLdjRQ9Bt8fgUp/CXZfm+CTHEkrhDnDz7
6VdNqopxpU1iR2OVspU+nejLjaQZ3hxA0X0UsZy4fQ3KyQzi3BhClA/ErM1H
NdyyuPy62h53X57espNHfsgZGfRn1ksgRCYgPXCQzhopjr0oxxJXLGxkTBct
FOs6TM/LWlDqxzKXIdgWlTmi1hs/seBjNzw11ZqYFOsVgFA07vHF7okttKZG
C+EkWM06aVZ6eqmqYSaCEgDhMV+NiKAy90i6US1ZXMvNpUWujjU/wHY9wrNz
GCBniqdX+BbHJOQMivZESFrzwdC885pnYh/DMggqv1r6oUMMWnoEYw4WO17I
4Q2qUuVS11reIAuOce7AlTV4e0jSnRVHIXDo01+1GjIWlNbn6P7MZh7o5/PE
6gaxjSp40pONKYN4j/FOb7aivpCwOHSFSLvIzwkkb7qpzTAUzAhlmHWzLwRl
xnywCrNgSOZTZ6z2JFRXGsYX3K+wB+9EOgXFrTSKFAzTF6KM52DZdk6Ciate
qehp0Zqhes6xZz1esJR3ODG7EYODAFvEgOiJSh3kiRmref2xEYAQwKjeJAM3
NgIsRuIATUzrEd9jnyhofSv6Mh98HakKGIF9P5loshrlpH76tngwTUACh0Jw
6Aag0iiVC6L2MFUCjJNi1rFzd/VfMKc1s/0uMHtzfBdoqwAWlw956LEBS6Zx
QN+x9Qj7uGimLMKq7TAMRSRafdgNcml+DDN2CMMGsp6xdRMdhjoL55Wx28nb
CaQOThb+FOHbdD8lo5gkKFKpNgvG162d14WjBR3uzVwCT23HPALdlDGy4DHF
NoZ9fYpU+Xwu/sWjjJj+WJViQ60udf9EX4Bp20NONJOprLaGZHVC25go7428
U2yCuk+0reCSZtva80RhtGQFrQdmE08mYhgh7qxs3+lm2zzLRNEEO+nkpqPA
JgIrrRZENnmEvD2807F8F78bUxp+BiS2A0NDBfUeUu/1IVgd6K8Sua1XciNq
BCW7e+eSPJ0bEBOUARWnaYYfVol97Qbsg+CkwBtXGigq+gwSaOejeb25Gm2n
jiTBUxN+3VA91LUTVb0s/DOuJ4SElQfBT5d2lDdsPXIf7T1e8gOxtzwXnu/6
jgMnRRUIEAPHtdzFO6h7OKw5laoOxFchsbkPjpVnriBEEnJyK92iaaDXM5yc
9czqjdGMpQv2BIODp3rc3pMM5ayOh5sB2zUN+ZneO+pGxNwX1oIUKTuHG7TT
BQkanany2MT8hJ2S/TcJ7NtkaexIeckLLFo2Sj2evBFmvf5yIHGR7brfKkuZ
3MABPU2ovlMI1nWCTi3atrynW6n8A8/DeMyP/WBGiMaN6R+c2Hil6arNMoo4
a9V2GXSRxyuuuv5TSVMWhQtl7ZkxwhxwXTcNVHB8iAvQKTeD8Q0cLW/cU+hJ
2/jrHPVG5NrUKn9BW1wN+kKXYwu+PM06EItav5+7ubj3WAcC8XXi9CU3U70b
qlC4cAlELgwQfkAYhqA5po1kECUKLnmxv7mzVBxCzutQDowfQVWfi1JVC09S
QTNLn3a84E4iTfpLto4N/8OkUX4GqLrsRwpWbqj3i/phXf9l/Diz0A6SPPO4
IPcx0USTdDjKGqVTLB9TIVtwVB7ubB76fdFlLZoSZqZcAxiDRTKxlYcJ9TjQ
iFp3KwHHW5IKe5aIeiIObzcla2KUQytaJ+L2T4MCV/7fVCFcGOM5+k5l64aY
lVhXJd6rqZRvLV2OeLZTo9wlHRfn7cpfYiEmc0U1Pz2d100w54YFdLkAROY8
jN8w/nEqW2AGhcjuyNfR9okpO9N4nabc/8PGkkPWqLKmQsvG2Psba5UEBT09
lf6N95IgNLwVzJ5K9ekDIPxVVY6TFe2u3/3e1VgZLbkTt7ShEt1P8Lk/ZNsL
zY+0sjELjMbEwuu3z8tg4HkLQvsW1d2mEZTgm42PAGZBd9H31CfyFmsVDag6
gW8JS6HOuh+HYRJj78jkkqx7YeHe86LjLXXswARWu+9c/lwN5L3WHHrTJbRw
rsQTSARUdm1fN545FEPjpVd0YFynZ9zcKqGmR9viCpr5bybjRKDNOUPEK48Y
0enlZYCllr/gmPyuJm4MVwL+3lOqIDp5+H0r6SB5NxPxnZ0vLlrNHbKV9YSQ
DtnBUw4CDNhyCIvuKdyH1kcRKOwefhUb30bsnuO8maWYe+UUhhOseNLVGwRK
kIQhfcmOp0qnzqo3pDrFVxKFvri0zUBL/sSyu6WKCsTEKStWEQpF+AUAoU0I
IZzPaHBh6aGLayi9CLNrPjSXqWi7DkzeoZ9VYf/FB1kWG+eV5O6U9Hl0m/Ea
9AYtvJIwUFNhn8vmOrTgtcStOZysGp9TpVkHf7rtiXCvQm728NJcJ7Xlxysj
ZYyo9pIPohO1RXOEUPhvHzFihFAuq0wtnXos1lMi8yRsDDVmqaeTW59rv2BL
0Db2CC18gKb4P03K3+4140Ix2+C8F9Fm5JeNFW8I9ZdVoNAE51CoiZo+R17E
kqKYnGHdqxlRkmagl4+8F+hU5bGj7oUxI/HANRuZ2ibpTnEEebBb4XnFN+3w
PUPy0nsEjHaW41H2pbl9O6W847x0fSDB6XpX/2pPHQ+EY6EeQIOPs/NTqAyy
BqkjL+o1+4grDztwDudGVWf4eRL58Rw83z/K+u+86alz0xEBN4kyDDOy5NBK
Smj7HcGPNwwnIiJp4ybXsao84mBK476S+Zw1SDzLmNyNzdlMie0IgXHJ8m1O
Xbs2EVPYLxEnv7+xfDcmeoe9FB6G36XUYTaSJ4Je+DNhzeeqriyuzetPPlot
fjH1WxidgJIG9AVSfjrytA7S8ZrDub75QhuTfrTqIB6hhGMRCJn8FMUGwgDa
qJ5U5eHNeCrdkIJTmEBR5D8DQXv8U4zC4s8Fd9Rtty9EbX4W0znRPxZPwlix
CcQ6q8kAvPKP2NYiiTeXuqDe5QlSalX7YG71t8Wz9ntGTT0qQDSjGcCuk317
hK3ZiU11uS6E1qz4J5dx7iSxisUMydhxeMW2ELa+1FHqTwf+oEPXm6BDc0dP
hf93hUpXWinSv96B2IX2Rb7MZZDhRRE0Z2vFU3bQ3w6ZlB6ZKq6jlHrPlmET
u7SRrWpljxbDJoeurrrKjlNplje3x5mSkymDv6a9JhxVgSklqHxnP69nHlxa
P0Lev6RsxaJ/PgimeXU3Qjf0HlvC4v/T/zJ9U1s8mV5UKvDeTnZfliCQdUtt
nW+FuFK9UZrHqzYdGSeIt/c0sAPV/mxdD7D/2YpX4bP0NBqK+LcasJiWZ8cY
1VtJSJ6LrA8kGuGL/9qkdpKBtPcNjy9Q4eiVky04Kj395+kv9w1XF0Jb/6l3
kmA8Td4Wn9OlmmFwuM9Xv3wD5Ja/GxjdSGxVnRexGyxPFGPjnqv4q3R+ebdU
8b2oDBd9bU+k6iEIfzFtS8jYAKM5qk8LW+cqQXVQoKyZ12gL7UuIoPAteZaR
chiWCvToSO+teFVXKZ03uA5IO0+4Kdh2RTDrcknDlICze0rhqbwH++dKoCX5
6/SUXdpzKxvALkjXaYIgbvfSW9OFhRAnsABJ0gb14GZmxrQ7BzKh7UVyXAic
FYAqL3acdKNzV7IUB42jMYHMvO51+Am0ab3iS8dDeWBnUp8fnrH7ohksy9Lz
p0sKFJdxduS6wMTObc3jea6bP8enJGq4++hbvxZBCxcvI0/t3va3kIceCgmP
kPOa7YzeLvQZDtLrzO0d5qb5CuraIHNoBHVJCwpuHMBYGBP5Kta5Ol7soFe1
kIiYcmbK4U159DxLlehdQtmre9Ddm7YIyOSoRqMfiPTFAIp6gH8I5ArtrrNR
RE5YiZBwnBDM820o7LK+/JDF38wJgN2M0ngpov8u1JmpskGTAIuSmAnglHOL
qvvk31+1fGSwgB7FkHHdFit3654+cTjYPYCalfM7b8fmgUiD1PC3bRMaA12t
NVySf/yE//ioUlh+h2xOhFU9HKLP7KmyAu5D7dqiXXcg1p6Tz6UP1N2VteWx
sR29JPjGOfsoYp4rQlT/axrSpEZlskd7+WSS8mm+IXPGwp911HyLngVuoBVS
m+sE6ePLrm1y71RQ/S3yji0kfERWnWH90XVkG+bQ6uDZRza4vP63H+zIi2c2
1dxVbU4C3IQsmMBtvGWEDdi9l9+w9d/S8UM9GYIiMcc8vZe0e7d+4OsfA2yj
6wXG/u/emcvYc8ywtIF69XD2zyg048hPqwpEYLbyLk193a3/qv8NDIHHlEvY
SKk3rFVueAe0PiNVHJMcYJWGdyClim7MTGZVPHNBqice1GTSgHmfJSCYUxWZ
QjN9/GiAfE8aBYPH+/47zYSLkFKgjawRj2Z67R8Lk2ig7TgvCvasPXvvV5q8
7KRk77el+hPcLlLv3p90Z7QBq5Oz2azo9yozTwu78nchntAxPfuMi70/8dGO
IV+1UPurmkOuJVrYno/NL+izia5oibDXGOSXcMreUS4QAl1U61HFKETnINeT
dqBUNp8PuORsGCTc8DgJqX6zlHbNCa3Pof2JhF245Y1RSCwytxCBR5IoF3h1
uGYAWIL710MjPqEfUHTv/URlzQQL/dC2kN6Uj72gJzJv3RpvGZiqrEY2qHS/
W5NUVSQOtlTuntTLbgIzAy+6+MEB82d3Z4mm5DC+swP4XYp3rqqAMyFo/LcY
wtpTEinKzKO3XbJOXGY0+F8BanKfmZcXS27hHQmQcykwdA58cM8fFa0LHQrT
55clysYOTERY9658hJZTvpAjeSm2Fx9aoy90ZujF54TNsD/Pwj08mdjAjFWo
J9iTTQcpeQJD/7GzobDkEWPD0KFwHR2cOQH65mplKULUq49gHlzhSHP+RGyA
coRhv7WP1qgfhwaRV1+R9kN5opO7USWreY8/lLXgzz6i5PP0xU7kY593kyOA
h5b1pSwgbvmm5BAU2zCc/vh3THV7Jh2yPJ/yQkoNtCqCXgJHmL2CgZDbr6+D
qUyt42VYQeKwkYhiz6ozjtql0UKTwuGpkzsSKBFOdmB56BCOZeemZH7mTpa5
s51aQxP/cjRRRkwZmuWBi1bGUBEsCQHJOqEzhj/ucHkJq/iUDZJtSO5Qe4T0
XNCLrevnuU1mBCmzENxU2rS+f3RcdEIs2t2gZVS/mddR0nSKkn9LFGnuaPNC
sNt1FPZrRwLTyqRwnRF0AodsvYvlMD3HZhFuwSqigOVOCQoq4/37AGNyDKu6
sBeYs5GGJBXlfDqEsiNMVTcffm80zcPzbChJQQuvip+8T2+d+83a7LnYDbcs
DZDVDLBse2y1daY9EgG98PFkXhsA5Klc31v33xg76PPw3723MSrZlQMJAsFh
ef0XqZ0wEeImKmAv8lvdoXFeMIh0B5gyrbESLqo06cFwBgXWMZW1de9lakFC
YUoPlzdqssTCqSvhzhSv33NXyeIcfZiSxl3oZ6RpQKXFEubjOcCs8AMRMt+8
J0vpig4L+AotCb8xqGmwN79GKxUISmfQ1aegOJ5V2WNN5tXoRNwjBdLt6COG
ZLp4ezZw0d1RNrY/p437crd+lUYX1yqrb20nn72igT7o66zEHvICVocaL8qH
Ur3UDZrjlfgxWyRUSQ952sIepX7qhZ89b654L8sumV/2yi+HuLzjwcPlUsTG
4PkLybpR+GgSm+FFUVUBXz+ktVa/zM+dDsVqqwwTKx6yepv+LufVbDoamHfi
GdJTHCpp5SyQohi09c67gNmtSm3e7CPCoBNz4Ruf5rDpSs4YPkUSfneeyob9
MBCavtdW1Dgqf+UBfTocBQ9B4HuNLb6Z63qbGvSwtmNeYo0Ac0Mg8HG3THp0
CuMWSkTFqcyPFHWZ69a6Ow7zf0nmBgzcuheMPJ9aAccn1tUNzwOk6WNM2nEy
hkVXU4SLXuHmEPq+FEtUbYhac4t7ixrWQZG+PvbvtezwqMFH222G7wd7JZ62
ovq1iPhR9FJDa4Z7BTdc3pElIOwoDYMPhe+KuFlolzW9B/R8BMdfASOZ13g5
bqNuaYEmgonpD58AxPC2v++jVIN3eCocRzOJPaf4bmS6WdD0CF6fvwjeqBL+
iYT72mo/VAug+wwsd+ZYD+I76oWt6uk8MGZPEcZyZdydTfkY62Bh4zbHLrMB
UVDZUMrKwCENAuNL5p9R7jl0JZGuJo67Kv/ySOas/HZBdk9JsgJI2r6X9VNw
nZbPGznsGTVCqyIykXKTFwfMQkddxYYFuk6zdMv/EAcP/zQ6wWD1EU9eEOPF
EDMGZm7vdcVsSabpkTwbHFliQ6Qlz1o8hwCHsYi75/PECOUFt3poAq3lA2/6
Ud/Jt1VgInLAbnuMRsUCeFiEh0KxMq+0Hi5jjM/wq+cQi7oBns8TCzv5p9mG
kxPnQnnUcHyvv3bGZMcA4hNkoszhkMCAmGqn5xZrTUK1o2oDSNv7wduuuRmC
8CqbYdIwyLHMYh79C40BRVTaX8mnC6uFEslsH4SPRsvF+uo9R/VMmBc/4vFb
HWiMTxhmiOC6Vfcjgb2RVzD2AExd5iZ7/k1gpqb7ZJfsUKYt+6qki1/Or+Ic
nN7vuDotpWl7NeZyLGVUhBqpZOfhUL5xyyR1MdyBA342b/kIXs9VDF0QOr1I
ergCcXCzKIbfNN+LQ5ZUMcDfCV/6aYjEGx3zH0kEp0YUibjpWbudayTGcX6e
4x4Ekx3hWg1Qi7CWCa9q0CTayeZiXQ0upBUPFzIJZcKVuwcfisQNL6H0v89y
+PWAQPnms0Z9/5jRUkUHByHgWJyYnegbzOP6n9apOTXCR8C57Mo/kBljFNUT
siu5awaeEgnbpOF2YDKzVvf7bME/INIRaNfGaDJL/daxRVY6lnfyaplg97YN
s33s2APZzt6uWUfVrO4ixaziA4ypSrER9vtmRJWO/6TkY11Nvb9EfufMN6pS
zG3v0Mr/KJcfbtYCJpjybVYLigsReAxtriQsu60hg3VCT7oCiTBY1NNAMkHg
JNbtDV27wMctwzfvwHDnRAqcuXM4tZIfxlAmp00SCIYD2B9z/TymsI0Y+a01
Yf52j2RryPSbxcC4XKDylnbz6Ygi3lwKh49OX2AaQ9KriBICfgG1lwy5r/bB
d0bfqRtyOERcTG5scv7iWjs14mhU3WYXIHaG58drZCEtvIqBwTkyMTHB+Cct
DWjeA1DbRkZfFswzNWzl9+owjAig0yDj0EorzBKd7nWRuuP2Pgj05LzbZO3+
o2gWxCg4zsNBA1JYyF76Q3IqQmuiTr7BJDCN83+zb4xFhsCsd0DuUB9ESPFs
QoedeuISh5BNDobcHxIjTipMybSV2dzKqgN7MbUNz0RETXHYmBrjkiAL6iIb
znQj2Aa1xRRyO4GuBaQ9HfcfUNLf3Bh5uL0pd8i1405+mGntXChIV4GzHkdN
u4BO3OUDqEYvAzSACQZqtFOKlDyTjAFEbMUrnM/T4qJb9OYzUxWpRI4BSmIg
zPnqiVe0dL6cNvJu5aV+XVMl2L2VNZbhJQ0VAKv7LZkFC3aw42VItkcBTfca
umy1jPXy+s5LbjS08D/HYwG70cVTLHdgfQ4g+ER6o9l6gRpX2hBMz0xr4vJ/
xQb2PTOA7qEkRmOn3RycIP/VZ5UdXt31M9MP3+ngny/0blxVGHFlU+C3eheH
JBzofrmOPNYNBGgNHtXFi85Q+0BtcuJpMYAXF0kFwPXJ7HfSykQM8qYXH2Cl
M1GaqCScS8lasavJ2Jj+4Zr+yR2KfgmC5WwokLosNsSeVHGB0SxGlCdKyqcF
I/ygL20Rd9efQYMIrsRJBQKZ8hUGdg/drmg8u6KwAUgNhbF2lPrUb4sltxSk
NpEYsuz1yUUPc/w56Vh9iMv5t46yV+jWyz7iZN97UX357l/RzEqqUcUK/hi7
Wg1DATky5TfBLWQ39Y1te+kPvj7AKCQhm6EPpd6PMt9HnIHxRolN0gUNMoXK
vz1BOtp0Os+Th4OxeLVXrClF6jladV9X+Pasa1UzSzhgVZia4of5wJrzIXYI
qfZG4d3DiKx5ofOeSoxLOlfWc+9SPP7V9d67ZXVkx/fLdTIODAftHzcIHsle
d89/sVAm+jIyg1uX2BmhQlWTEqsiIiIDSduj2xWJY5O0GUFORLXQ3DLHicQ+
bXGdRnQ2jwk002vY1lIEbQf4K8hnhoU2O/AWSwRK4adjFvYkifzJdtZ8TWSs
Irh/9rY5mjrthb4TmhuLv+5+kHK9j06+ERmc7uNYr9VWvz02stLpKdCVj61X
ILszEBWRks0U9Z/5eQ9el3ZoAapRyC9eSY0X5mlvG4TiMurdOw3OlyJfE1eI
zsWRKxIeSO9IiFDiuBgC/Tkdksai0rJycM1cSS11703rksZJOdek7OtCAStS
y/sSaz/UoE1nFb8sxr/JoGnMtGLSgwON8FJyK2ZjDp0QqPwh8Ai5mbDfuc+z
iD3/ETOU2enDmKZGOd/7X0AoDGsigIKwt9xaztzDUa4IV6LUKGyfZbjfUbnm
dsuDFSZJrNl63lUFscdOPq31Jn4fgL7E0swObHX+xAibMUKY/lM4w3Ta7YUx
mGnJnf+imJVOkjKF6ITQxyCQQ3bPp8r4zUiZnvtOFMEdlwlf7RX9lhQYSLd+
XkLmbd3pohDUooVDuRCrcNE5dMIuaFYuUfwBMQRNefZEgoilO3cz8/7SwuXx
fauFm+4NqZdRYvuTvzMF/2EDHcX2QMecjoAP0M2VRgF/HdJP4rk9CmTPLPCf
ZD2D9F2QJX42rmpiG/FePZf0uzSPHhQ23ruz5cqGz7Rjsd/V12q7mGIWGyAK
vnATyCqjsobI4P+3IEzD/92Jkgfu3ACOmedntvALfYgDM36RcmIaE75D9CM9
uI3qzm9Y2VBak+JJVMNc4cQ2QLJ3fPfu2ksSNzb+4FiS0BmKfK7sHk5oj1RL
8y6SxFNN2/E29vj/uCWAMTm0yY5+RxEsC9OwyEOj5Y1B6svo1iI4ZfSdar/W
e/P7qBt6zkWmHKYAG4HaSFBr6LGF1GslcJfIsQqPV5Y681oLC1nsUASHSUgS
qquAzg4VrKDC10p20AJ2mDp7+yVBManfp6WVf+XgcSWpa3mSzXVjHRNcY4ea
9rbmHEJnI7BgK8TXfSzdH7mH0uIlQyiqliK+Xar5FnH6Z+6kkInSZVnfbRP8
SqTSvf0D0PWyW3U3H+gIhXvw/ta6n1UEnKQaXfSOeTewRtN4QoYu4d26POoy
3N8fbQaAWgB1AqRjJ1gH6gA3sMdBXBWjTn86QtAp/iRo7Ce8dr2p87odfVMJ
tbcFn/9++271THQdLKqCLj72uZhH92x42n46R1B3FDgtjAR5Cyqa/0jtD1VB
F2JbUthhf9mqt/eyX7VXgeNSiGNyf6nr30erZSppYXJJIlNTFeAXFiFwM5wH
xTS9HH2SvUbmRmLIEy0FRZovpl4vYWxOD1cVH7bL1aad8NoQq+RajiIrF6tL
iQK7IAXqxt/dlvRRwKVJzZNMorSbjLl9XIN2djncMJCT0aZfw409+5J0DzvC
kkwY30gp4CMxNGlYS72LKHHLeoHCxEKzMrS8Gi3ML6VoeHaNeI7ct2sa4d4h
qglwvkT8emxfOzbOavr+0OCdGtKc5KcTJIA5Cd18wN3oM0oQ8PPc2jejUwKi
GYZ03R4GT6Fg9lHOh0/sXd0fnuKGY/nxx4bnfwGb8oYt/dwLEao9P/F2+wQt
qOAkT5lEj3OpocwBZPMKWpG25LJjvgoHclGH/aB0ovZ4sMlCAPjI6DRLLq4y
FNzi1W6hI671VMNC0Yf5pO9pNOKUIsHKdMeZhHloraC5vSNDsgvMONMCk2VR
YI0k1zvWAThzxffoSAQ2OmSaiE9cVPHf9C1/vVyRpu04F9MM5PTKlYoXTH+N
JUiveekj4vz5q55hAnzyMBCG5/wcUN+MOqAxouWJWYpQiRFE8dXRuDV+PiUu
B3vqFLPmwPvex+IrLDyKwkAAOloY186HIVwKjXsg4C8AVBWpZosDBKKklGcN
gwhJQvcocV6oYHUaJxxig6jZr5YwMC52zPXsiFP/w3zjVTnHVDpjjST2nCQ2
wgh/76/o2oW/7FVl1OFcFLFXcHAcxKlcuuN3nlFJUzRCYcCs2RFtgeWSuF31
L5J/lpvhJCBhUtYVvRks0mj1cLHsMD51phLArdHJOkf07gY5k0ViArsGeYzE
xyV30T4huvUXMXs4+FVcy90+GXz92LuxkYIDAEdpn+ZEJwpuL7dwS4do9Zl6
h4zZdCmctJlQ/FXW3CZaZBYRJpdsHlJ16qzRBLoMckmlEN6sRuNsgz9orXTl
21sxkqGXV8gls+syxVuUBxbcLkdVUco8UBRVbcsAwDSIpiemiPxTXk/rAH3o
xeTZdPmor5IFB0D8rqYkmer/UwP7PZwgbmF+RMPGhYyZ5fCZ1GDqENG5y7GR
JA2Kvjb1UA75g/OqibpSaIKTXtHnzHHtESxDJKUeRNI+ZgO1ieXpt0N0kJg+
FplbfyWbvF8SqRugJ0QuJXse0yPCNyQZMKj1PY8R0XXoGnnu+YMprAroOLr0
7QnXQucRx1i9QQ22nxGFwFUjhFcc/EoJxfQeFNbJZqyn5xj/H1E86fPO9XBI
KzgEGjpp/N6vmT5fnuxoX7t8HNzp2gOko0tRIBpF5xXE4jAa3jNrbDpu40Oh
79Os35PKjTU+j8VvYzdFtr0RxZjJK02sjYAfGVT8tg6euSSunem3qg0Cawz8
Ua9MYFdnGSKCUxantzApBjrjiIV3AiAnR+lqyHsppX6jkSOaSSBULP1jXrcq
d9NCCrtkbfyjSG8puzjtxLE33LKHnqhxjHu5nWjmwsmkzyuuf6mfsKy008mW
FV2FYH6pNAmNzHGe5eaCB/6yMRJNdzrQdmm3vOeB8Ppdr2Dbbtb4d6F4ElDK
SBj0AdmCQ19M85X7bC0JeGSzIjHB0dtImw2kmc8KNAmAkb/AWOLtj+Bdxcvi
oB1R4B1hHVVIg9dX53K3AfcMubAFl4x40sUboLYoNGtIsNirYs70fvFeiUcJ
dD0bV4h38AgIBVWIjsSKuAPW0xvT3XslPbtmbDlPmUcn1xEhjF4bVD/3SRsn
1onvUjHHiw7q5vxnvv9kuWUvvF/8vDZ7L+VA7dX8rkV6rP81miUXbEuol38I
39SJER9OBOg0Y0e+hxwo2ZvbjU9rprTSXqwvyf92OT+keXZUWDyz53PUZJui
T+nvaz2EGQclZT8yayirJhuAWeA57IYpBQ3T13gsOmIkxBYZVJeLwEXjYuWW
o5p/3PwLOJrwuwgMds/xPcK1MvPW/RjAic82JYwRyrnnvTQNRGWKNMeYSITc
Lg8hNqypn+msJHz4pLpY51z3BSb21AsuyOD7saXRHjt9l1XNyuWw2zecubDJ
DOB7fN6M5JfEttyW6Mtvhl71qhdDzINT0fZZAZuGAYKxgnmX7YWeB9ndnZON
bH8MX0bl1EYGvZ0pyEFwmkKY4yknXulC+ifk6a+j5AfH7UT4ZV63TQTDGy8L
PCte2XF7HwC43SLdhs37EJ/Hs+UE89Eo2CQIrUPWDLnIsvswv0AOpfZ6rptT
3iA4Fh926nX9n7yWjiW0bzNZUkwL/F6qpfPnXFDG6ZLCaIxSR7CqNr3hwglU
AflPdMmDJ/uPHxDHxO9Es3XT9wFqsVq6LFXiVI6QYapuSsTGY+Fr7pD5uJEu
uLK5TBLbYUn7yAfdH67jhAQ5H+r/WmBtBDUnWvNKNHe0dn+hNQ1EPssQ3CAF
j4y8p0CKJOcTdY8OLdC4GIzrOFHNEUClQbEmzrNhg+0ug3SO1q4nkG8WS1cE
AYooykp/ZxLPH6T3mB5gzuRv4vnXhGrxRskzRF9en3HflZik+bgx+bTzWXF1
oN/6apfcyKr/Zl9I5qaRPZuqhLY+6zcDilTHOetXoyT97VuzuULcrXVD22wc
WQi7ZFmoAvZakqQA5J7lCzkQN7s4pwL4UY06CxLG+h/Xt4/GxwrmpOjzll5r
OLbQHaRhaxffTJ1iOQnX9VCuUMSfPi3uUEJbqlx0BAZ+mFPaNXlN4ECwlNqT
EIcNqvjFnxW+gJ/dTLi0oUBdHNdGfbe6I91d0SIS8kDXF6yvgKzotOQgzr9g
vHXChJRcdR+sGA2KlnTguwYj5p/XqmOBtX8ltonGeiSpT0ASBExP0VWe+in0
p/iiUypU2h0JiOxKeoBGsVxu/4rIBxnt2zw+WEy4CsmhLvHwi1DuOzap4tx1
pgY15LMilQxzOTkTr09CwZTrY7BDuJsQDSlbZpHhaIxumqxN22J+RIlozW6A
7DZRPzCqp+ffLKtECOyhwzWUS6CHlQXTxYZcUtXsA7K5NRcs6LBkCRVgPHq4
hPsxiTsCfQSfQacBSQWMu4zwvaBjrmkkDAhWm/w1zpiCPoSG07tXpUqEsH8S
PXdjyQFGm1nEMpEgSxAqCskSKy3QKGWNTMGF5L3igwekMBibDk8WgopqlA1y
6UCcizlAkPOF0f8JUPrtDWohFdHjjLSpjkrSErUeKUe/GVuylXje9v/u6EAh
n6K2yC5Ob0+oV7GzUGEZmbGznD93Om3uAmGjl76nfyXqn83ELCnSPztQd+Cm
D/aTdU791hudP5IpN9NdQxIGRKleSf4jwQwFJAfmUacjDMJTTiUicr2kpeIJ
Fh/nKbLNyElAvkEWbhHoL01cX+Q4L1jq1EWM7Wpr0zHZf8Xr5PK2ND/k5TPi
VdfwnUrkeXdadCFKN9p8BxAm/HWgTTNQ7l+vMK2ZJt064lWuYypfL3dSUAv2
EWIYc9xi7bTyxNp9Zg7y+J+lnx7Xu+UauFK4yuB1u2iSLSzfThWlfjz7QQmm
UsqixGT7NJ1R2qOGL52k2Kj/CxAUpheVdc9UVe2+cbK19DqaRJa5/J1ARqFj
GE133uxTB4Jl1Wm0gibr9/WyaD6GkQFqvGlRNof6bAI86LjwJePFrvWAuzSM
rVQMRK6zykgTHd0FQDxAlDP8NP/+Hx7Cue3L4lA8tWHANpZXMhauIwTrBNsh
Gaunj4NT0u3hJLUU0HVZeKsU3MeFic/ppxYZsNKosf7/FPloqzc6AomPMwDi
TR6fNG++cRzMoPLe9JL+7476eTGeyGYpq8dWqnoVdkC1hR4hax4v4lHldQlh
vl9ANvgBApxf7VuD1Ll4QfImuCy0w7aImfC0dmw8KRWWxoW2Yr+H6cl8dwDZ
j+twwm9BXl3WcUKPtsOpA48C++Zok1oRkXWSgT43EsHOrFg4JrjmoFYNING/
1um6FKkxWRprTcwnNFDCBIpSYlxd6TYN0MNo9QpMpMIKTCFMl6z4LVyfIWXs
qHG/3g/KaUKLIhryYlKEGlX5vWyDtQWzHQxeB27rpa98B1ofKGEKX+yfBpmW
s4qwkawBlFbjCKbCODGm3LvOlJaVr8xnfA7v75qx0yz0/nMyCFt6oULH1eMh
/ND3hzwt7rl29AWkdK1KqTMIBVxpJtGnnga2KjXvhAbHwJPzxwN7DflfPq87
f+RB7Zyu84KILN+YioE8/k8CHBmdewQVABzd+glsIf3y7lZ0mZ8ZJ7+ExulG
lysH6DUEWzWU6tBcxdr1MHGQftoLqlC7EQ5TuOBgdN1eN3UrorP5P4cFOzaX
NszHBqcYiIP2RVafHznq8D4j7bjpPd38wfPOE1XyIpLlJwz23C2t/M+MyGwo
MbMCstLPEflqviAT6Xxb6qWO3oV2W31E2JDfKugg3DwOBzAkcTVYd5JlRF7u
e88RQCTV4wqHifaEXptFDsPfX1apZ6wNorPqcv8c1WpV9Tn0E45AanffxLZx
fWyvUGe0c/Ubgj9Ee5juWBSjC+9HdrU9HWHbU+om8mQJWJ0rGzGl3LMtyV7v
AbjU6eFZ+vvYHq7OoNsZUfbEnZo0ZXZyNZeu6baeDCc9nXDHzN2t0XYv38Cw
2Rw4DvEPxMn85ZyPtPYOgxg6JGby+qKzzdoJhBuYXK8SRF7R8IYHYmlIx1hZ
G70MegTpLu/VmxOTorOYDXWcoAv6cTkUsd7mFm5e9NH8O3JKZL/RlpSWnngj
o0yRjz+XDJkcxlWq0ouquckqLWsqUXjorAAu/f1oWWZwyMTibAvqTo8mESqq
SSWqUghV5VcGardiQjcEJywkayp7aqa9BiWTGeMVzp5VhbLqelJwuaNKDkzE
r+lG1akm8Tw6kfhfo4vKDrzlOmxrwlZMXwB+TJtq/Dbo70pphbNHOSxNaQKZ
0XrMhGv2uC8cy4WQ5sauiCEK96x65cYzZ+DQE1MdFpHoOTbmd6vmZtx7F0+t
pcOHsbCJWIcNKGW/8+6QOIvsPWA2ILc4xKwRT6qMqLdKZRRLZsVwjEnqYrW2
U6nGlWacBmGPnS6ltGmAgX1fdWCsaESppZGzO/lWsLe4aMo1ggbpg85FrPKe
l/946Mx8FtJXZEe6K3RPI+7T872L1IdozZELMgPtD7sD57BBRroCgYw/9opE
jQtxYD/oaVzg/UYpqaHVJvIHt83J/CV7wzsqnc7PFYEd9LQp/228MT8odOeI
YXhynlYb9lie2/M6zFdJIqal21WwWcDDbw0msGWmhRfVevdcOE+/WWDhPN8J
zKcpSHI3gdsTUHgQMOCFO7vZi5a4hO+thhWtXkcmmpFhswfpSJnenT4IjrI2
CEWSSKnnz4s8xt+mT7/S8/k9woCbsQG2m8l9e1bYon01yAV05zYflOolXLlx
HSDeCSJkSWpmQipVmuLi1X9QlMDG4Tv4s+ySamZ6RmvDv4R/ueDlzGCSrl59
s28BzzerpYGhMQmgclHaOFgOQcAQsu8J5Rz4eqkZCo13Zi0/FdRULjDGJ3ec
hYvs7ERW5T261k/dZ3pEOeKf0Q+usodp30pBQlxFsG1ORD+4vCbgiFaup8jY
kYAG9+KQHtT81o5sRBWtUDKOfpyAKQwDLODJTKBUwV9wAjpkWcMMKLeCWn/u
b2dAr2VlBPxTQB0yBnF649vGdAV4X/3fN8SqPI4jHccVzREHEgEwU8R6EheB
avP88vdn39wRbGnh10YBQHRIJwHQb25IS4tgNUQcR7pd+gnGc1aSgQe89JRk
En2WhHeO4SXMaj/srguQA3rC8uZk+0KCnLN6K7+VRIgVt/nSVtaF/zzgPp6N
hQkuXVq9fYpgFeFFCQrS6kw9Mx5cA5tDxBa3YVzsMaFcbNBqPSB0keUiqsfa
JmsG9qqlldi1UdgjFtNiDA0QxYjptgpnC+rIab9Cz49OltfrwSKrbJvxXR1g
kkk17K1m4tYqdYr3ACAOXXZL/xWWMJekMQVN5zEzUTBeJghwCoH1pWKyZ7kd
iWciZzxOmpDv9kTB9tG4rhGEIYOQeMKwGKSgE0uIve7jWxiviej+1IueegWO
qok0ijjyKBPIwuVp0MCP9cgv2eBiOC3vaOr+YadOtClRTixjikA0OcTwtJq1
7nzLmtGOqEeOWEm0MAkqBc3tN3wH25WaHGr7xk2mJUW/ZA2Q4sidRO/ioGhb
lAcREBycIkTOznzx7LXh8bam0AP6AvaJuplUYne3pNhcSHBxFjaDsJs9KBsZ
HDL5hyBIOVLRCWd4FUZHfuQ3SC6KP6sc6biz8Yn188GGWYKLL9+3WEGw9UOz
o7/JlEhsiaaEOrjEqjQy7KhVijc0f3OQyRu1UHv+uEF+nldn7adc+bMFz7Wf
UCiLz5xMMn/fIhzurxMl1EutXUbb3tjkOcMVr+0+HB/VPCNVEyGg+rnp6cnN
rmRrP1bJr7bIYooxzn97/c7YM6pQjK1DZ43EYVMxReFyBGj1yeL39biXGyfQ
B2zO3J68ufEfXqrjU86pzVjF/VbsMUmPTp9NHoO6hx4z5NkMK0IoUWIErirs
aMKE1OnyKXGTL9bJoQiX4G/Qbm+5dClgRvhzX/WFIAy9xcGUMO3XWYFOOpM7
dYy2sl/5hKlapUpngNBHXfxKODQRcUPs91fdgZDkZEpuL4hOW/9PndP/Mtwg
kAkxcZbA1ahJLwrjnoWnh08Ro4trBb2hcCOL1oWjeiS9b5dPUrHCycyKmp+u
FsnHYLRzIXPg71RSGlZLbyCp/ud0rSwM+MLLLj6W34mH58Q0QDrD3WA2Tplj
RcDgBGxNjQRLvBhqfamRe3bYogJlMlee3i2nNd/XS+K5pLyb6ip6rvIPKPNY
noUHlv7uvu3CVYWql+dQ14rDlrXnx1kcMwZvNBOzESSIHD6NWTKU4sUv4ZL6
Bx3yUTHY12BODrTarHjC7L1BpMme1Qo0B4VsvWxhCiG5wNMWW4JZpZyVKHkE
xz3Azt6ZZNZ7JZukdiHnYJqpxL9NhqBnbxJOJ382yePSa0mCvGdL41NU/w/3
ZrMmNHgxFty9PjftTaUyZ7Z/W5h7ZGBzSz8UkJi/bi5ROlxApJEjMzvfuLYZ
OR396EKXFusE228VAaAT+eIKoio+4kxIPcp1vU2GgDUWUIj30I2JQtmex3/1
wMgryK9NU8uqI9goKZcvKdDsKxtObBI9LUI5q8UUaryRAt2HcO4Sarco09Om
8TgV7jRegQqEMcssnJYH4bBamkCqYBBwJh9MJws6AAaY0v01oMQKzN3LsmDB
91tfCVm81Ea5hYo70NhH/rnhcrrrxF/7rinPrjRIUmNKUu0HWnuTfWeIr54P
JkJukPXkVQRS9e8Nl7B0Ls9CBbupl/B9V/bsIGEHl9HNXulA/E+A5InNLFzD
MxEAXetzdLyfqDrpI72lZeCqGSv49R90VIhTpSNsvg/g30rpFkoLikxoXmNl
kf0KxZXElqVliRuxseQBmAl4CLzmAEyxGThzSxZM0snWe/LoEy1P38+gOf1d
NLOBFAZjf5oA4Jpzvr2uWSa4cS6mBHSSYnoojPDt3PbOcPRdl+PE+Ve7J2lr
go53L0FQSrsjCINEA+giOwjIi6oPDWBOGxRi8jslfb39DrdDt2jvTkLwmfYW
SY7460EfOHRfcjrF1e8i7qoQJAP/Vw/HKCs42PWpnx/8YUrB//H8I6tW/amp
w7q1pIc949vBV9JOgcDblPtSJHnCjAx7RC5hHcQ3UBxRopy3BmCXkJMpiOzP
L5Mep8bbdA1OfpR76pFYHQ58HXStfOie+UxpVWhWQaownAl6yNQ4yLm7TtHS
cfwXTCaWSokQzSyZOOXzWm6urv13OezNkMirOOLBZo9TIhSE6d9zjT2Wd1Vy
PcEf8bYnFaiDnKHkD8eB0mG53i7YuCCN38WXLpTx2fJxG02JGA/lfxoC9Ixh
FXXHd8y4z/luSD4EFuEYQK9xkz1wSg3oe1AWgfNmYWnrxB6pnmumi6zEJdu2
omkH5iM6/Yt6X9/gDOmCfFp+uZ3VEhvwEWnrKmclmNii4bm+Rqs0PDYXR4p7
wHEimrpQPFIKOOEzbtp59bxEArW1tf6/X1xqoK8lD/uaP45vUEaMLQxCg9PG
OQLDg84CO0X7z2FNyCRPPTkqU+QEcnKjiJKrodFMhe2GWfvPB6vBKhfvaOKY
wscdyGuzKUntdeC+H1FdOa9IiioAS85NOm4Sj7EeHV++tmWHvSVE04GXS5Aj
3caH7Hn3A3LfQ2zlyg7LZ/PONIAx5iFUcsbpd4trM3GtZlWnk2fjlCZYruSq
WO/WLVH0t9Y5LTfzy0tNan5W+ABPowlXqCbEhBod5n7221K86+yMf/CqZwuN
LWSm+9NGAkuMgjRosnmlabaN1IfiE50uxRajo/xfQSpz+4OL9V6Ug2uMQ8P6
vPKtcja8klAI+Wn3JIglsLT2hLYPU/sJJQInwCK3d+gPEnN2WKpsrZftg06t
Y1NHIYvKGa0enHYVeaa7aZarGdmOA7oczTb9oG3LwiJck5l5M9TynHPS+teD
GfdPf50NZXCSXXtr22xmCnrNSqAmpt/BO7DvjlamEMtOaK5qC/qxNx6q2MQt
ZV9r4/XsPCMquADMRmcGwM3cAUyq+L0XbyKnc4HT+tVxr4atTrNOuCTXedvs
b5EgBXGwYCQyBlT/RKusAHLIKHNXIqsVyReMsJaTNhbRxp0AbRlcU6TwIG3k
z0EUQyVOowCZmJGYN3V5KM5GdeLgb4t7OTInPyIQ+sYO4oJOra7jn63EU6w5
oQU33xs0eG6kcDdCHsLUTjxbMnkkR/qEYBYTMa4ogGOFSTIOZ+L+4goldjtD
m7xFyAbNXLcxDd9yj7zoueaUHSQscd8Q5y0C6J3MSl8dU7DjzuTmBOB2B0Sd
vzhIFqIQg7sDqt6+HTQdehoavuXn9g/AzW4mV+IJpgiSQPIDbq3Z1X5lai0v
dnl02xFlDyOYR5FYa9s89GJ0WD2ul5xCOtO7GLCx3AO/n539IFqfKiUfY7yw
oJDX3lTSamVFDoUYpu7dftYtu6JM685NI1aZr+GVv2thKFKtnFaEAnW81IG/
fES7DE60lEgLGssrrVxmsxvQrunImUQOunWXe/hKhsHLFqr2mcnv4AynzNWc
dRFcNl4sybRUImCqwcnJAvmRnALInDI2e59QF3ZakaYFqZhi2QS/sM2Ux6xY
OwAuTofmRXR0Pv0jPwFpfFqqhaWTAuOu0QKUmEMEPWNGS3i7IWAppfwz/lbv
JCjtUTWAekSnWMUaY3EiWowL7wd+lSdFrEu0Iz9nf96UJ5ATYe/eDSlG2enj
5XUw6ZZ3oEX/XrpkcTuDhpFtf+3qTm9ls8Ha4xgcwEqlzsberpXvFM9yjaWa
6dtblg6XN90HV5nRxFsPJFA9iZq+6SO2n1Erxd7sRqlSOJ6F9QFLWxNuUBDw
59BlKee3LLFOPYI89IiGBT0eh8UHXxA8/+MYsEX2KI5GB929yE0AGv/NirR2
+Dz67kPP5ALHNU+S5bibnobhKsW1zNbb/yO2GMfMFv10CESKb8FiSdK4RsCS
JSWDEwZqI7PJsW4X68/dNNuRDG1w1zTJ437Rc0pg/7p5J+nteYIUNNY+v2B3
dwbrofRrd2SoLgeWMxlTYZJRjaWmkvWy+uWaU5zl7I6AGhzrXOV0KIUkxdft
r8Pg//tct1xnOeyyu0J98qt+bl2DSZgWLoLlfBNlkIoPsusZf+C62oDc1x76
URLGVfHAIKrOBJ5WgqOt+ycUZ/0WGcGc3FK/agcoRSqsZGJhVKeQ8L1oYYi7
aAy0yUOfDdElBOlWZmVVzsTaOqX9+fVpF16Bmej0utv9IE6rbyEJGC8TdBFT
rkYHEyzXLd0oUjHwTmDbj5QDG9NR1tddTX3eWRMDmrODDQCppQOxGNocFjb7
NVdk26kKxYfXXKnIbunwVqpDTu/elmDtfHxVBOgHFUIfzT9RAD7PV/bc7qEb
DgFaOvWyKWN0nSp0IsRKpfmdC3Wut2qCBzrC4qMgPYEulyipo2/FDP+lHabK
KAnOjzBdx2SQ3JVplAz7mUEB7Qmg83PAZ/ADOQ9vJLvJGiez0+CsPXqSkAaJ
g/lYNJZOcYAWpkhPXx20rTKNei4GE92wiwNX46kw6BYhxwSadZ9vfK6InPEg
M9diyHeuMZSl84QMOCPvicdmOpJ67He+pyqXCCx7xdORkXAvbhModIWwJlGh
qUnVmdnnWvAHbSx8jDkGai16babxdE1Rdb29wzBfg81OWtXOJCnY+85otEUB
pxZ4ZpmMjfTZ3Ug1sD19bNB3WtKiyBHb22eZUNgMvgwbwKLf9dbu2igqYTrs
hASMUBe5A5KbRvVc2GjcPghgwITVkxWY/7N0SB25BEutsyYiwY20yKW8xZef
cAEd+3Jle5tepk4C+1L4q9aLDg9Rwcoat/xpC8IdNGv4FbGC/Ld7g3/cH5sD
hGYrpcJ+FVe4Nj5rWqvfLmKDHI9hY+fPgctUvcPHvL7OBYoV8D0YTlJp9GPC
seajphvJ0/yoaI/nr/I6yQKO0YWh4Oso2e0uL831NTdPCSvt5eyG+3c7GYJF
8Wks4FP0yeKi84QwbRrJBe1MXS2JnsZevFNaIDrnyuNlV+HOfP2tjLQmJ+eo
JRdw8URKnQOxy+xdKIrp+WOqFEEhJj0eudwhmRFDWuxl2TQb0RN7Tfa48C2A
mxsh/giQYi7qK+egVocigAEffyRIXtjyOLe203z124gWwhAMq7X/hdUZMVPY
KJ52LBWCqv4+IgIEgRv4As/ABUXb4I0NA9ijA3A1Di1wugCyCAaTkMHi197Y
oQh3vbIUrQTp6h6kpn3W5McUj/cQp2U/hCT8CsP6sasxiPY0tMK6pcCIyJCg
BbXArJkkUthGZHFy5vPi/sUBp7Pf5FP2yfUDtRFYVFNJHLsvO7cWPRQUmjzs
NdwVwl/j2sLaDHzyQFJBPdYOVmFmAg8NK31NoYmGlZr8Sr3RPDAVZm2SxN2Z
9sorZhmiflJsOFp/H9VebXCTwq+YsgB7gIPkSetRSqg6D439XXJWwo4xenmT
M9yzX1OpeZ0jFzcVE89qTrjBPQMHOAY8OnPfiZzf4trFsa06IwmCK/EtS/c1
Dxw6bPPRbCx8CkzJ6T0VA/3nO4hUYuNVTmgVhxGA/JQx3sOnI7oIwy9VCjWQ
6+SvDA+KGA0kCKLw7D+53TQEAue5X6o+LAUAuk1ZnoW8ZlMe1OZ7/FaGXRsB
pujBXbygv0w1KHKQbVL4XSHFoVhG9YMuVwWbjBRjSDXLEUSdGpqB78jvZ9gV
3PjtAK+7qBM7dub4GZvLkVt9Fuq322ZKTR0mb+xSAjUogQ9vV12IKonp/Z/V
/DCunrCgLPBr2DTD9DpNH4VuBLndFrGMSXcIjBpAH3MvdJiK5PE40x3yXyvR
+tGYFp8G6d77qDGO3UK97pVBE/B1qv/exInYeDOYIXS1WaHiPe1kHoE6fevV
qodC3ojcOazYGn3d9o7VxE7s+oVL6rAUQKCTuOOb0C0l4U7rac4VhMsFMBJy
/u8ZgjZl88k6bjNHbEhpdX2+ETVcWKk2J4CmPI8tavicsvk9HQmGYCHdioxc
qQGjCAOcGLEKp7J/2hj8RDCm/zO22t/wntV8t6rt5wYzbRq0kJ/jZakoM7mo
s0nMOVVA6rcQNHSOiP9mgchtJHxHkRYYTYb9E86wRdm/+M8Ql8wY1a0mvgy3
qJow1bfamhsQIaNxZXkNl2LsEbuZRdJbVRg/J3c2u3IhUmKL55N8XJctzmrP
d3eDld7m9YB4mE7bU8/iuzR4lLklLKZ5w/LPLxd05Sh2QR20iyL+JshVXFxV
J66oRSkPSP4yT35ER8vhPN0OTFGHNJIGrNj6dc0+HU7YGJ22HTA+HI535nuG
it6UL7Ig2/U6d9AW9FHZcjkK5JgXCMKUT/O7D9bTVBDfTFPOmtF4tl1iPoKe
sySCCC8LmiBz+42D0x+b2JLHsLUHTjmmbq9jqZRFXfqXxs7BY/M1rgOs5JkQ
i1xGPQIVme6uHBFJk9k88o5RffO0cUSx5sgoSbSMXKJBWF2VctCAmgQPkXOt
+EojShfhgXplFJoFRJ2pm5tJtJr4ZS2Y/B0qZdm64rrH5+scELY15/5tav0+
sjEh1ROSIT7frG6iCasBcwcbMwR5r9GAkUXmKAHu5hJnnJG3FPJJ1clZ02Yu
JK4vZPIiLxg2G3MJigUKoZKPJ5yAPIyLJToaOUgmE/QzBlsEepswqDfb2Fc1
dS5yZ3TBE4PWKHqbQkzVvP2cHv8pQoKwgruqozU1xQ3XOXmjiaTY7e+OcxIu
iTyyxywg2jSwVpkNDG9BNRhhQQ7BN4T7PeQHw2ey9kFh7eaGz5DIdnV+Gb+y
GMS0xAUj4yLbwzpwplEqJWe/9fVmiKQFM6B6dZkwKhBLpBxV0OgO2kODG+Rg
R8dfp6fome36Aknhm/tPyHumR2KNWspxjotPVfmG//4kXoa61R/VZkT46S4F
qH1iGVL4hHKHzRqySxB2HyZmKAwcWJ+sXZqYUY3sSdJL992MFabw8jUrG46T
VYzrHcRX+srI8sn6V7Rvpd2c1Y8LDa27B8HLDYb4YVq/paRlpE3XTXLi2KdZ
Xet532mqaB6/pKBCzA2XEFW5FmNMZrr5iuB/MJvZOwT0VwNYsy2/xllxw0eD
TUf9JKJpZVFd5DTMtzCexKiDZI3z0u3fgkxcnn9fVoEVKpkJwYAGb5rg1Oh/
r1uhPpqDdS5UQGkWGDa2KCC26hoBsqHXBLf9U9QqJVy5FPZN6qrV2zhHqomH
BQARYr5nQb4TCORpxoD2DIVbJmxWk4hv4EFBESDSLSjzuiBXMAkDW8wZNop9
tjeAscKwpPzP9sjbtEJ2qUDGPS3NL9DINZrzj/FIFwfOl7Og6T1ZG3L5l9ZX
SP1MpokAmLZZ34coFFEuk1QlgNfvt8kQXPZTQq0W7UZqDFbNPgp/bglKuQE2
GlwGHz2UUiG7q0X7WM7xMgI7ND93GWFIahMyAbtTs985yn1sF+q8rSydqk9g
7iOv2mp70B2LMMCLHsQpZcIYeHGpq0U1aOQKCO3KCfXgAIl4mlqSdU1vxVZS
Y2o4zbza+RL/DZE3/QIKN93pl9TYM8yu3j6xSeP3Vuncsmsuza0fBSpKnxs7
K0FuOJvLXcj2K/TtFTLTglZ5pIKKp3k2Ad5igdmdqTnU1meQ18dNQMnXfDXv
8BNZnMH3Zf7PN/AI+7nIRAKWBpcBq1wn9XkDYZ2RBpkHA5afJ4UpkbRN7Oyp
i7+m/IyrtFHsChbsxyWEYcp4qJa6/dPlKDDYt9KhE/EtpUTU55NQZ4dW+i7B
i/Un3MapTq+gok+b72HXpr3l9zgmCES5XmcD+OTxp2hlXXc5u+VqetDCMFbU
pTpTSiRBR32FcYwKhpyMOBXtmORqdRGYUsx+Sl+pzxsHZvMx3xnI5RmIBcgw
+ejVLZQUWrb4NXOIDWrZXSbgUnvKidHioz6ZauLid6FDYCWnjeIcTp3uqKij
UJYUf3xlKCiZdOV4akLpoAd3Xre93NtfDAHsLp8dMK2Utob2jW/QKkcVEaEA
aA2P4wGh/kgs3cw/4d0IQt4ha2Mzn3bkYo1XsYvTU4n+aUJkDbnYiIt5H8lf
LEfKtBVpMbQv18lGU/N1T0/8JxMw0mPD7KpWEZc+qaSKzKn7sztaKIc5RMHW
je61LOkEMHl6AjJMBG7aMwDjVR/y4G6yOlf2RzHqeXobB6D+gw2TtU/axyls
YmajJ8x86M8p5olbnWEPTAZocmLX7OQEm72PpeQeoy/P/MyicPHx+sZzg1vF
1JV9R6r1nISv1KaGDsfWWrJLqIiA4QCz4pTx58gc7dkaXxkrQ76cWottfzYt
VIlz+Ou03YiqSfODONOyajrZDKI6APCWANT1bkKooc1Xzc9vXeTVBwVuVDED
rnhe1Mf4oxHzBMF2pHjjCvBrQs4Vu5y2CanEbkUm4tmtwNBFUQMo8jEHxdN+
KNQAkINNGJO6xGhAufBgHdD1MLdwEZ074kJTd7XSgoA0i8pbMsZ02C2Dx6NL
g2op4DKpjnQrJTT4HyacZZphsVuZzXorFGvWAbiJ9GGuhtAKuW4NC6hlJKnk
6DhFXTp9pT3KJ881+JRPJS+UuIvbeKcwEny+Y4lV5syoWddTMLfPpWcGfZHA
ULxHK/LTovvU3Apu6pgy0fTv0rIITKdYBL/qytEu8lSFLFzjHg6WScfJMIAb
Ir8sW+UQaW0N4UiKbCvoN7iDtiIqq7C82rjE1BuNS1JgVDJFp4N0qhstrV5S
RtVZ6oDpyuOO42BDCzY+klIXGrTdzPKyZJedMjyp5atkhdeq0cldM0tpTpZV
7G5BiQH8rdTZrCf2uwNmbESo2yjw+ZpVhxC4DUPC8VHcXgY0l34alUphdil4
MD6rDkPaTLp2AjnLD/FxjwC38EFGL73auQ+kAZJn2AAKFU4KFs1Ti9qtZ7Mn
ZNmJq+1cvp+04tDiVxRqmKkRnzNXqCmFFbf9Xgl004ChXfO7rx/MftHyM+Wl
kd/XL+eBSOfYZ2vOEcpEk+HnpXFuec5hJrtmhT8Vb/1lsGaz7EsDFWNEQpio
2Hat0Rb8i2Tr6JRfoWz+cGoUNLaPbvK/CSI2fc7sh19Clv/NVzjea0dSHKPV
vb6XFJ4LbJ1I8n6Oek3wHwMG3xWg+9/LbUXSWVYKBOlG1CH1Yi3mfarJxsSK
Vv4+7TM4PLio0BBtiDdJlUzFuk24pPIgQKEZpoBysPhOmUbZlBiGLsN8fZal
6v0iOJH3bUneKkLP22IIBQnASRfKvkudeZYQITbFIKbs7Mq0NOYre02RGtsB
m7aFrNCdsWPoXeHFZ6mVNpPBLA3GhGC9s9YgYh/BDjinswP2OpC9KuRwcOcg
jsRaHKUNrlHBNB9n7aIroAO2I3mebsFNrlm1uq4k/xsZi9mF/GYHpG+in1A2
W8Sorh9o1dngw5GRBOPhTEiv/lc9xI4it0wlwi2qzJl9h8qW9TqMTZJBQ/NP
h4J4GhL/Cu18ku6ZtZ1xmyDSY5yh7wRegkE6oXpfHqObWlm7mOD+GmnoS8xX
5vwX1yC7kWau/UDOyCUf5e8YGyfWG3IDD+jKDWc+Nw1jqbZ/92AnO/bokQA9
/O2wfAvFzfbfTNz6OkjvYslWvIaCAfUIeNjNnu1tNAz92Aiy79fmK/IY1gNX
I/a/jYcWIm0qHjoOmtu37BvfTi0rMUoKUaoMYefY8o7n2UAFTvEMWfn16Q3m
ZEaOwbCVEXnTaNN2+YEOmM+Z4Gji/ZtSzyrseovtl7SXRW7iZt3hVvzU0Iz4
8NZKyA88B9adt9Bu65eUCrk/2mUxgI48sctCBwhxZ5eEtDCqBbGjo/+hmJ2/
q8+FzPHyrxSFF6Zp4xsYWX95eliU2DEyYC/5ycuUHvTV5Gc0V8MVFudNIsw1
27fNRfyjUrSNkZ0weFhp8uKy/+xoAb/9afp2jBdoPXZRFaAtc83ekRwJZh+c
SA3uss+3KUzb52o+1+XTSgFc5rmveHOX3MKql0O1goishVL/Tkr/BrEYtFHF
IAGQA8vmbxz2CKlLaA49KoIobCNUJonAOzkDbFQhridMgp78n2Yjtdbt8JtW
bqYUTxU4JatYLo7XjuIJIv4x8Eck6hzxvmdRT+QX4aaTWLJIP6DRshTgI3yN
DObM7qkvxfA4LQ4TlVnUALz7CXd7aIWoQXV/sPam70RWhs8dX4ZUewJN0Fos
EnZzSc4dWr/wkBoPjQ3Tk2SEhl1jGHhV0dMX+u81JUv6jze0oLgqjfnTKwkz
LCFL2oKJowRRXd3lJC6YQzJVstU21V9dhWrxUVxkQFS8tLmBwxku7fP6y9nw
QhH4cghw9wtHypn5cekeOt3JVhe0HLZeWghASFEjlNXZfFZf+m03oRJNQ/Ia
bNjs/h6mhTLPWOdaUdbZjuUyUIZDD7O0Ibz5HkqQH4ZrU3qEY49/RkjrUo6S
kEJdKjmkij3IRzwWFAJysHFLYCm2AhhxatbdAqwlR1kouXTUqsQc3nfBP3IE
ms4wJdpC4RGHJdqkcueM5NqayCqSlewCqZ2wM2VJSepdg5ZiIXYRk80i88tP
3I+1cCFEgmERpXdM8LFgy/lgH+56UhD7ONotqA/CZPpYo4sBCavudgvqXCJh
Y2wMCUwoR6bIvg8JzIiYnaf8rEsilUnWwZsVFrNmDBxxiGjpRk5mHJ1V6GQd
7J6KKksFBaC7iAxkBlABeigIltLRCNjfpSM9sn1f8DGkgXOkVr4Wcg4KXwbM
lSyfq6Nrns1VW5agJnncUyBrv+ybOlXs27ymeFGunxJTxVK+qgx10pSxpw5x
QL5BJ8/dRW37njWxPXS/DFecmM01uXxhgUnUsQ07WDf/OBlIgwJwS1t3+l/x
+AMxy/9Dn89JTPpNRsNw/w1n0qraeOd5l+1P1riXGqsck+DN8x8xcDiiWLeb
9tIAF1VMIuv/UjOt6UmwWNNh9NO26ymKqCAuhzYgneB4i42xubE8vTM/Krfy
AM3wgGVrnJtM7SAtMbemt7Dmvh8oq4ZAKaDbGT9/IJ1sLTT5ofV+j6Ha2Zl0
RNyFy6OqtZhtdfQZlIlIrB7k4ivSyQWy41WPdlS46xKI+/Lfs0n9Rvkt+laH
AnaaNZ5XVRkXxwkz60Ncd3dFFSV1+NXEwvHDzpSEonVpU7fV19YvFp3L/tXR
v35nWVnXPOTGiSA4wECGwSt3wo1FVPpXB4SjvG9KQOeGgSVYXehV99FKW60t
fnWvi5bciXu5AwwhSCyV/XCkktLkTInVnpCZ7MxH8q0T6Jvl75MnIxrzM4Nu
h1tKQIhQW81COT/VY6xu+cla4vFZlYq39AF9FMUu6nWASBNEP8aPCtuHUeeJ
B25VobQucV4CrCfDK03mjldE3v9Fs0EtHbEHgXp7YN1+4NXlM6RkFHowtWCc
4W9+jaHCs9TZuVOtRsDG7HOqlaCJyJp8x2PURlF/KtwIP0KDJjolHlFwAAQ1
GAY81JBEnDqm7dQ38Gigmk8AwDxTAEqd5Zmr9jWSfe3zvoZmLldh16hJ4g6x
R6UlkkQ7wdZx2f1Iadgt04EjVv206u0LJC5eVwLrW2408POpFsxxlpPzxm0n
Vs7hTaM+KzGblAcm1ix5guphBAbbUe1oqoGKvD9i0g61j7w0VkeaQp9Pk0vA
upNPd7SFF4kaNsM4/U1HFM6YuyQS0U9nV14OzINDhwPxAPQFL3Aq0d2Te8r7
GVvFAcLYUE/SRpZzXskiexAS3ZiAqjMC3NZHS/Z/NwIjgDs9jWRD1hkEKhMo
ESoVfqeweaLhz+TgC5EGCXuxKfXicM+2DJs7bVo0tF7jl3TeBsCZYWjqlIlM
q2PnkXsDtO/D3lsG40pn7i8H0cWsh/cQOkBTPBna6Pv32CQaM9yd+b94BSf1
WfwLhC0jSZ6lR5orVjxTe9q0LZGhZhNrmYlmpTM/JnRG9rkEIo5IWomh856H
Z4X36K9G0iaPTBS0hGSquKLyEh/AMExCI9TPa0b2VnKM1iNc8Z7GKJQMf3Sp
qU3tmdI1pNBATDAOvEq1uSMcCAQ5kA4ed+YqF1DXpLwEm+m+TJlYxXJZbFYa
YVIscOUB2Wzq1K0k98d6xaVhj4anoT/rnx088DMLIby8NMI/vuq2AdQqJGo0
CmCFcsgma2PQSdGQq6FiLXwib1Dk+3WL11t+cTSU4KhY1oeGgkXAn2N/I0cU
JTcDG93R+GVTIIvkSOB7BMXHpQ+kRBrownfeeBZqycDa4Zqgs8KMYX2gnujD
xccfOftWB36s5vNDTZQ5Y4UIVPyAeoBF/8H0LQ0qL8ljIEoqHGbtAeGvSFcT
jnhMIhz6aFdSJjImibjTpgu0vqUA8htjBZJS+02ZGa5SlNFr4vJSAfrpfpoD
1YCszHLrKO9b63RZcKxBMGabNtDRtSI8D4MMc5crOnH6HdJQJG+hInTEmYhK
VtGrpPeVYfiJ6GikeuIP7DPl7P3aO/ktaf9ZedAROYnDyUVRUqKC1BKHaHhO
r40Nrsyx66O29nvmGHBDeVnbpD0GYEHzM8EVfQeGp5IyU9K/PQT8zeMCjFg6
jbaq2iqCl+pPb4xispRnTgLAIulR9ftos9N5e+UTCyWiLcKkIiQ4GeFs2Fig
Das7CL3Zt80Goo2DfXMvOOgnR5gK9QeOT3gtHIbBlgHUgxminkChYXzLFSNl
861saygskUwkbGEHPY1iai5PG0nyE1kZLJms1c+kkQTkrVYJJPwgxdnLNAOs
A4wrVVCQB/i35G6SBkgm9esGHFsMO8EwqlWMWmxZCf726Nr82H2krPECCtn0
Z41VsvkB2k5g2/gAHII7ORpsA69gMqB1tqEZwJ+h8btKFXOjJ9d71yBOBi7r
G7jiS+5boTef5n7LQwyN6vz0Z9SDWiVE8dQcnO2+wAdg6NuBoDowCEG95zuk
c3VwNZhDsejq2pD4F+t3ZUtROHtz5mxN1jy90KOt9162apVQdHCsS8Qoo0SV
ykDi/a/A1lL0ltNEGHJJGpMVDPY5/MkJ3GljP91rfh5ea1FtsLfwDJR/Q96f
oPFwCzfTa9K/T2F6bTBsntQIAT9GCRCaIOIpMEnITzf1cBy3RjnTGgyMLO08
U/aH0wq6J5syB9i+aQyT2qZGvFYeFA/+XQAxTRoQuMmhfbILyiSMgqeplydD
MiCS54hjnnA/LeluP5NgvRKv+C85mPSuEVjTDr7f38b+4+Gy49cqMPlyaf9+
wAJdKQoB8i6WvqobDdefZ0sSBltCQ+5HNd24TpTE3yJoW+bjizWBoUebV1vd
gYOdLL5xNiDW0HrJ1O6axIRaSDFKJIYN6xeyqoIq8WZiRG8C4l3UHLdYQnN7
o+yLE/dSmEOUQopkhl5QkC2JHbbWgRAhYDHz76ZMBxfNAe5zz34sEIwtUWoi
xZ0S67MxzNR7J1DSSkRFdiXv3xS+OyHnWpn4Qkx8W3zbbFVQ+53kvFuxk+lI
3MvAfr/oXs3bUMDHFydNGNQV6UnSHtdm9sP/xBYYHsRHxAdraJvGkM+zpVJB
b03TFBFGkamic9cvwLn1QzXVKT3fi4sMBF2IJiJdLg1ixr6e0U/WqUT4codw
rTiizx638NnQbgDdy6Aw4xQ69k9NIIqd3BQinWBeKHtfUzDP5m5WwurZGfIo
2QRTCI0Esc8Mo+HWFpf0pd2laRigHd44SHvZwn/K6Z01VXaJUJ9KXdJLRGAY
Y1Qk5Zx+hmtmUpf+UxJmrGTdtEsv+BtKhlNs1S13jVKoqM/E/ZeEHqN6bLR5
H5AYAlZdBGBw6k2KB7gzoZpGT8mBwilZWyt3E4rxmYO/m5aqgRwxlz+Kdx9M
R8c9J+IhNw3EFICwIT5CB0KyosEYuFp8LajtCeq7oY05iar/+wjaA5yPH8Ko
njmV0ETDSrs8xaVygVGviM1mz+YbeOLslwLDxqoHsjp3z3bFtgPMgR68OSIy
W2fVIP1n+X2swv1/ow3MeK336QK+TAlOJ7ZXleR7CrIuZgdfdKxj9bMHitJM
XTKc/VM0XFFfQrMgoqfLZbZKGQb5rvrqRTkhQCVW7S0yNLKwTi8x7Rb1FfJK
4TaKDzUHnz0Q5NZg53MkTB5+cgZaxsoMgoxp114fV4yC17SmkpZJk23gMXBj
yNMt2P44q94Myjy/qMg3shLnqnXZvy9Knj4ADR+hl6giLvhHyG6spYs/z1Aa
JYcS4s73gXpT+zlaYhJscQImgt92SAavB00k2JrZah16N7e/HkCz2o08ly6j
IujNfxyiPROzuDn+ayaonUchBsRATnvoSaYDrVVQxrK+YXw9RGTOd5jwhkbc
CjEzBB00W52/iCWTFI8U3JpoKPU0NQwL7JSZAZJxcHxpRG6zELhaio7Y4dA/
OJROCme4/SxJMjCDMvrSoSrOK9Jz0r8d+2iVGfCrmrqreWd1L57Qd6UPkg0G
J7Y/f9LbMcRo+rkjgpVIImm2UYMXCwNVzqctu89m5htjJP8a9yJzFKLidaPi
HEwzzaLpK6ywqXpI+56zlCGuwFWCiIDchGwbRQpokB9tuWl0p+VcwQrM+NJf
ESKt8YYQWoFRyQyh1jaE88bqflUb8tHdUFMRha2WK+uDGa4GsyTLL1b2S1EV
wd5KhqtfXHeLz5eMuQkl77W5WM9whxKZL0t2kxrk2S0gC5gZfPHZpkeGtqhf
te2FO0PinzTAWGlo9jgy1uJM0ekU5Ky5sh2EjG9K2Sna7+iNZbWryx77il8A
h71aZD8awSHSVpMyvjZPNsRJmA7lqDyBMZL1cpQRBBdZUx5vpaMZy8Rq0P5G
NLBn0jK+K8WL9tO1eM9BCwRiiFCYZ9MNFwetuyGGC4hzyQF5EhFQllFhrLL6
RALyDziiUhWmXZCYcCrpT6VkuZP+LveS0hj3UmeiuB7lre+PMoz66M3tSKiE
IvjiEzfN3P1s8I0luBU/Ov/YP/ki7xjjkR/KarJOmGsKFrZCJZzAyo//TVle
Df5dWW5LXhPqIuKbNmLaV9bjkIHGk76Uyvzl+w1RWHmuReTxHbwQLs+Tg3rz
Q1o3QZF2okpllthHa8i+NeFbQrj1n19YsJmrU9EP9LyMrozLfSWJ4RQlV2G8
iQKSM5YWj8MHN0TyYlc91UVSrZnBqUVcB+1tCLEb27dMKHM1SX+NwUwzil1g
cPQG7bwkwFVZOWvh7LywoAC+V1G9VEgIlavWxtpa6SusgxDW81vqGuCaZayR
h0557nKdFgnrLNKi7zRGMc3grPwLk/ZVIjlgi1qt+BoCg6bUC++lkgca8uEY
n67OwfO2G4q0BEyex35IHhd2selScI0oT4/DwIoq8mEnTDKymdRCkrwblawi
DQGvuc+2qr7aBt4/1YAbneE5kLFKBdr1PMsDZNig0ypWQB3OV/HjsV+Ut4HR
zsZslqLkYg5MNGTWxdbx9511McwAQ/jSxvjqjI03SMIV7NNIPLimzkSS7CZd
RCT+orgT9QR44mPLw+e3VUjttrrces/7bsYB7cqI05WbolfUzwptrd973Cov
XkNLrhwPeUGoJZTbfIwTbCGJIzw4YdupctWUUX+ccE9bYHjwswKzHgwKDN/1
dbqUypGAX4J1qclpXmZSCH24gVj2WylvUXXh1txuG9dQ0rjIJMZpN3DkruOP
AskwvTPGTWUDzAFlT3KtY3UnwUmOx0PvvtB5Ae3HMcxE4fqju5Zpc7WEXwYT
0D4pk6su9/VSgIpAsJQJtSRl5WR25IcZk+NxNJX4k0f6DlaTeZ6ARC3ygJH1
iP5sd08KdGJE/gTVf7JvFJAvSK10cakS5TA0ZmJun/tQ/t3B4+tVCLPxJ622
4R/nZS22uiZj1IgafJdVEidFTmwtRLQY6jpESYmDXiLd6n79DiyABKA3V0N2
IrP32JMIT6GglaN48umc4+mb7qFMJx5i/NtLz4gMa0c6Dlyx2z3q/xY1C1rq
9jRAwcJHfwSJpbwqgzry7aeIg3TgvUmXVFgse+DHfBoCemBu/bKwac/h2nHe
A++DPsIkeNUyQevOAx4ImSkJCYg+SEtFwUhJjUmTL3rjt2oU+O+mg5aHejLL
sNusw0dBHIjzMHg8a4hcrjk5Ydrf+zEWCHfplGNXYbaNMoYnx4odXoVhv9KV
2zW47+TqvLg/Yb42R6aRr2ENztdkRmaxn/JqgrAjj4LAZfowLEjzi20nCee0
i+9WwrlBmcJhmSHdfRlG2h25f2IQCn9XNMaG5kDxTPjm3DNp9m7jDQOEq+0t
/2lYbf8bS+5oqYsm/QipoAUbQoW8Job0QawX2yW47wI95kDbxtkKNG+rxbRi
sTWDEsfanHOiV4DIenhFTfEmQX9iNrNLBykT7rXjqTCLc21wtSISUp10YUxN
mCz6nSkTJB9FjOyE8PPos9PyCOEGMpyWz5SFqMpeb5jd4UGYGwjBbGL8Ymii
Y2AGnheA9tfE+YfepfVIAjVwgYgIK4G5iHstxN7gXwcULOtykxTozD0XQwL0
EvenOtBARLXL9HFGhyaETMkJ1sq+MPf0cDYSe6jTeVUIdQksFig7JUx4ZzMq
12iqY2pItrtqHZXNIWMFxJOamvUONkrJSf9wK9vItZE+SvKsIidEFrnfHbR7
fJ1Q07nGFvnl5R8hnXnjquYEOjJSQ1xK0Kq2BTBnpgqJJXT6jsj8tZ8mCXa1
dtPkgurw8dn4m5ayRd1spycAd/HtAX019BDuuIxbelJOgfXt1tS1kavVZyU3
uVOQPWzEdkZmtLWI4oXG7SyfWE+nsmnaCD5chvC1/PENQsnmAPkGNT6O3z6y
KsFPnwZxzr8A/hj/kYVApxOuti4SY9LGBkfHqd8sMsznlx332B5QoC9x9dR2
6rtIwj0FjD9cUR7H6u+OxnCaaVhM92nQbY6ntoR00hgBv+sCSQfcOvRGWryU
zbURLQh2R8C4lPeDjEUQDEptvkWNKYse/XY1rfry9ksqfDFXHHBtkjCGpBbk
AS4rBZTuIo9u+QxnZi0O4t9SEmiAZAXEaRvcKhXY2+fjuy9OSv/yJa6pn9r2
Nz1l3M1qcn1+VvM8J8+htuLD07cxO8s3wYS4DfkT8DsRhy6mnUiquUgX5+uZ
S9LIO3QnEwh9sHvGKgdFUvTHoc/JP+SZUEPL5hFqrZfPzpLESm2BhxufTz5+
qI6shq0TmSwWD5PtLiQnmCgwNZvVUohVN+YWTLv3Goc8Hc5tH2DLml9bJGpM
g0Bk9ob1aNiUHxL+TtESY2vbcx1pzs5YFrnO2XRLS1yZ+YrHgoVC9HSvTfYn
kIRf2XhBNO+9PeF3tjws28eUGEuvNHbTqaTGmxIfV1UZ9CEgeG4UA1aUPxkH
0LhdSa75hBIDk99eYWADXMNObkZIbKRTU9gw4XH+Gk+Nv+cRVvVJsOgNDmBD
Bt1E2zYm638pR0nJ3NKvgq92MU5mljNqCHUUjmdXEDFJY90tlUlW2tFv3jZt
YJ/UB+6SjHCBZCd67cP85hzQctllsdp7iXVDJ3UL/2Ai1HPQ/VVO25iWg9sv
SWV3V+M6aGYzRsWDKzHpH4yS1x8cN+529nScc46QHo5T7rNOIBprrsCeLZ1S
VOVmO/S/z3s2vFJ9UHXZZ9x4X2xIuJOEJ/HD7joiPoHMC0Nl7iDa2rZ6aIgY
b6dXvlhLobewyfr9Nda4OELu0i91qYdVVh7sVbkoBRPyeGX7zVuhlNWC28Uy
8jjglmYuZFwv09QuFv1D2INZFqN8xSJbyMX5jguQ7TT73ap4RbLsxei+e+yx
oRGwRrCInNXTuvEOUoRYA0oBJ9EaVlvzVZoeb+d7luSfmjyNq4j+re3od7KY
2pspUu/xte+LUp+dWqF6IFYQX/tXy/Y6FC7iXStRaMv1aLTO1hwIuqg4GWfl
p0UjFJY5GB6puENws97sTqAYz8DijW/+QeEsCskwr66zRc7Oy5JtM61TV7PP
MiSPSOqw6/pnvlc+FgVMWGDTAx5oonYSvbtgpbZUaGsYH59x+2BcMd+vWWSN
MiC8lYNHLQyGPY9SJlRzK5yI6qS57bLZD8ZZAxOTZ9jQYvrdSp6p+JX3yy31
kyFk+vJCQ4ndLhGPQSnMkwrv5S+UjmOu4DPVq51Zrr0RQBr2xQ1kGr+EM7mM
emFtw2IzlNdSBvLNeyXfvv9IS+SRPn6IrYI+40XunJECV3efJjHzXo/9PRwo
o/ayv+eAZzsTioE+rGJz60GKKyKj+Ox463QPsG5scrkTFd4JezIBPOHlUX+9
H0rHerMwB9r89NU6bCtU/5AY+edfHjlSu8QWHWvtUId1r2a2HRwgiLpoR0WX
cNpNXeAP1WpI3CvtGC4aRfvD1yrPsNlfKnR7IYhhd4BA+ngWTNKDMWHPUMzs
uiv7c2BB7luw5FDBYVvVZesHxdCI+U3xriTAZ12/pWKrZBOwk/obbp9bLt7/
Aaj3X5690TpUuWqTCaifN1SGsVFXM1pUvWJEFpG24YWLJNr+jOHH2epuNm6k
HkQQ7sBY7/TgD0/+dv3hGTodSBkti8BuG36DYC9pHs638icO7fUBFL/0c7M9
7e29zYXmyBzsJYrqX7vWjHvGuFOfmNNz0x/24hACMpcF8e/pATkyONv9mBcK
jeqjdvlIpDpqLWsvoTqqNyRnlmgA32bVI4ua8wE4zMXj8BfA3bfeMpdNFr2N
qNr8Yk5jsm4dUh/MEN2IlK2QUpSHlUHMQ+WwXWqxhfCEEPx32eZOAL21LUdg
55sNpBqpIY3axx1xKn/oPsvfv3tMTw8hK6Osg2JFuTLbQljOX5oHbMkwjK8x
wwsoGC/NUyAUxLxYBjUJOoG1iKbyrHKkytRLpm2LV9D8PIO26rzJsQj/FTjP
xmZCzvPjKhZS/f2sPiB8wj8L2Jz8m/MpL4ooxwMMQlHpjixe8XStrBfKxdGu
cwaNCl8DSNVS6Y1PlGAl5K5Mp1PsY2RG10N73MtI3BdFSLyup9snfgKusXot
g9TdNlsBpQATIRRbP8Z6wjTBuWizeclinm39/t4O8q0GNvPwAhVUpTornt2y
To1BTWAgmegkmV7BrzFqkAuhQ/TncXv79BHb16eWn4oeyrGl+hyA/Z1En06D
WfDsbPeaW0U1UrlltXTnvbotdfuTl0jnwHx11libk36AM/AH15NKFMbWN2qe
lmkC9PBHNeAY1Qmja0wVyfU5yxlSZAd3dBJDVMU1DqP+J7DCZSKOcH/LT2Qg
9uKlqNrkDEZKHz3dYmqKiD3PpwRieHbZtkq/vR3ouL4rcopYwHm8Fk76Etd9
QQLQab/kxneuOIs4McS2i64DVkiZa+D2K6TGYQMIyzl9kcSBOsyNguPxe9dt
M9uh0qHBHfluXtXeVXAh4ZiISjulm/tvin7jPHGww9yg8rMzjEHYpD9rLiwl
aoosIDY7CNoWyf0GUkvl4Oh53eQrzblgWET8egj/Y9Vqe9Ak3LCJTCBTW4YX
iFm11Fuj1c7Tp5ZgDj9tfN063vDXMi9tUGiv/20j0WxjnZwdGJEDg9kuW7BL
0Yw3VV4nJ0JsXsuDIvFeS89LiEuDxOwUmKYHpFvJraRF7tjYXkfqii5LT9bA
Xite5i9+I9tsQjukAmtsM9FSC+mEV7m7D41M/R7So/bxJ9SUpxE9QHpJm/cy
p7gdWDYCqOrF+46ZrhPtLWSrYLdMNREQOsa6ZcQd5J8e5hCGvy7CRsflense
aeX8sRir2+HI+C3oA/r8ESVR6ihGf0c4oLdAM7ol+uZ2zR3sKun+XLjNwJem
EceLQg40bNNoph7d0/vlds0lYjzQYJCHzdiw4CgmPY93ab+VwgdhMfDKBk3a
ULbsqC2Jm7RYUEga5UV0+pgzppo6p/vOXkLJn15MqkmzMdClIQkDHJn/ttgq
ZxQH5+LfyZoJ7lrLhiqXR2bPYGnpNavLPH40vUDRiB9VwRbtriapiXpAcntP
c5QRcWSYH0RUIIS6ghvI6UxFw+u5DiEbyd1WL61rDnQ3z6VqhD9nwrc3ZCCO
rUDrqiYPlJ0G6J4CzFnFCu2Qa4u+hkJSb8/yZROPrP0l42UPEQI5IdMvWWuS
sRn0Tj+Q2lGXqe5oQims6E5fOvESbIvJKml67iRrwwST9/PMGlMRsR8UXOj0
FtoV+rzapPNwN1su884TfZamlignVIOW3lMnx3OCT7jITvEsDEQGW84XPiRO
4DdksJcdwA19yxLv6/TOCAioIVW+wl34vGqNVcgiQQgOXmT//A7OscGVulNF
dUHaiUdMs6Fpw9dlvqVUPHK9/R+ZvNGiAOjblPAreQeoa25/uGA0DGdsTYqA
KrmlY4djOLpz+7kOEAEbTMmcz3dsE3sihUdDXdCaj6QGBpgQzEgRBXCWjsWU
Li1y7QVPGquQN2X5W3PkUAEo632/Cno/wRT3NWvLtcHGvQlz5eHObfelQdP7
rLh18L4CYmfEoF0N1zZBT8Nb/tpJJu543M1Yr8RH6Tqee2OoZH9O1SPXtG6T
dMfycbfLlzjnIABWtujBHxB3VRfcIGVZWVvlZhJ0oLgQ0y7NqQjuPVE0qleH
oYNuA1Ib5GHgWts2nRgz2NY6kEM6qcdBfc3w+UMogRS5jQVXk1rx7oNhibao
LCZHIcfLBqy0ViuKuzMePiQfTuFlGqYSlzk9aEhSdfIgUngGU0IJC3qs94fI
3ZTr/3WA2uuPlenkaFSP0F4VpoIg7yZnp5PPA6guYseZtgnxF0/e0juTcbz9
yPDZvgC0H5pDZ/7dE+H95l5VqoHkRtunZe8mPN3APpk/gYl3g3E5tJD0

`pragma protect end_protected
