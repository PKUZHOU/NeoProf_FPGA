module intel_reset_release (
		output wire  ninit_done  // ninit_done.ninit_done
	);
endmodule

