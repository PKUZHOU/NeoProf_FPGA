// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
vZgZkJkCb41EL3KEliH7uKkyZFME2577NRd0XY+cFpfurN+X4sguO3rUT8so
KrVtSXpsWZe7lgQQMNUc2WdXP4+Sxs5/KTpvVm2m0JoxUzLOXv60emhsmoKB
gc/zP9XGWjUZx2nkcYL53pQmlYkqGjGTNdgCZx2ST4uPXP7Bz9XC+r4OiOGq
6GFs9e7qU9QeTK6m17oep4jShppNWEoFe7wVpK5HR5AUjCrnAfiucxeJUirc
LIg4XWI9lbmlYrCwGkXT5fs1FvDA/cNVZ3n2Y5mUXwT77TN0zZZJ7LufVYVc
vcs7+momhK20GIPZynqVsWmvUoQJnbO9SaTruJ5+xg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
dcF1iyEeGkNBDYUwb5VfI5IcnfpsWVx+N9oOQ6atWuKNsj/3LR8izuNdO+d8
tHXEzSnEz0+80LwcZNVOkez1PilN/Ng2agSMuR4JiugB6P12D2TbhIqMNOY5
xeHpwFrRIDjAFb4ZpErnJymTvSDrGgdTQkJBrdxhAlonVVqc9aFWgtKOMvnE
0N7xPEmxvoN3S0+gwGG2kbzKhaiwvDGu8awSyEDA82yxL2a+F2Sxj5XUEuuy
thMR5WPWwBdoEr29Bfxv1IoQSndgZ27DJoPCVZtESJvUvrWxlHOkC8ORru1C
jcg61sj9Wnq0lpmcmWVzLveBwQemRZClbqB5ib8A/Q==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
eZEfxHr9I8q26Qv3IJ55RfzkI/0ibWbIwmq5tt8AG1KC51SonfSEbQyR0XTA
O+5CRvieGLrJlZ8TS80bHquN6ziyRt6l18W9o/d+57cW/xR8zWmrjJxheDL0
8rWbnGQL3yP/cWC6H0JB04xrHNn7BC5zSgCUD0OBvfaO9FEalhZlXyQpoGJY
oobmHBIal9dYuSZf9X04BTLybPSWQZWE/oAvBMVoUucOTRveqOe3uJ1cKyFB
t7vd2AVvL3BtUONek3RbRjYLpWS5Aofd9xHNZPNmS3ufmqv+ci9yRbCM17pQ
jlD3nSqUkyeKv7/aCFLwAI3hX6WdSgiLke6tUMK/Iw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
X6AD4njOcYv21FvK3LYSrOe0WhHTWcB8L0X+mMflfrM2ggXcX7jxKnF27lZt
CdR7m079UBVEUJaTE2d6kxNSfA5tPBGnZiGBNNNh9ZSfmqqj7O3xFwycWCum
c3Pg7gSPKBZxz75kidlb6bs9Jlwki8D7ktC4bQ6dzu2p9oYrSQI=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
MNWT0CnOuR/mxoXCAtElFFK2eH1R7RRz6GGiZjrBwf7r/WqZozMhFb9FO+6x
5h6JqMhEkeRLYVORCPzoKoKZypxgZI78/nzq0MOLh5h/qUpKPNkQTf+OOKkt
C3XyxddxSOjEoXCkf6MFB1BlEzEcYDZ7mnbI6Thv6vFmGx3ZoiZ36Li5QuC4
KTqZaZAwcXEc9gcWeH7WXa8LEgZYY+aDOFsxVysH+q/QBkzQg7OcDYIzlvwn
i04x2ztdAFJTxGnQjKO0NO05pyHOvgvzH7Dq4mVWr33Vv3zcslsMy/Z36AC7
/ay56w4AlWwgFwqAzwyD74K4FF7UhYDjNzGxU9yTK+J4hdZLNdu7r/hJOZHa
ASipjc92oU9/v4Z5kIycQ8vA9D+/wa1n98QEAS5StEMYklU97bem1IHHh9ZL
CiYYx6orYXGiVYYaehhfMOwCWGUdKpcko/9GHx8/tKqbGh5Ubeh+B091q+nu
dpyRjbGVTueQk661zb85xhF7nRYLB1hj


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
eGrgPh2GtWJhFOlpeMsqesfOV5m2QnC3CyObL6sb3+vzQWaS+TkH1NIEh0rA
wNnld/kTL05OJjGs/k3CrxlWyQR1RBpNFMPLhInd3f3jc0CM6hHt68ylEfq+
4WItdEwZPPDrLsoPZv/JvRBLngW/SGTvqKVXhw5/mcYc31kdKpg=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
E9uErTEXUwdIUVci1KjKGmNzA+OuesoLc3jrOGZgBhX5Fz9Cwuv1YCSwuoQz
2ReQwsSTHFXjRsM6CCvomfOL4RYG7+knMFwjXPV6/cTNcTQd/nonESPMC6yP
OQGzvCvu5QzUQh7jDL3Mgko6AZwlNdPVEZgoP4a0Y+01Mv9EqhU=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 84400)
`pragma protect data_block
roblFlGxvvP6Kt9DF00peO6dKJPLoROayE1oMApiKv13d1cdLk1N6LssLUBs
YbkiB8I9FL2YfxD0zw8Et3/9jMSMSCWflNRo9uvT83O/40d/7BIX1yUxwJcj
AE0o6d56J8I0JkLIIbvzs7/JDOGFucrsrFJ2g4nLfKeFgW/1228dFHAfn8Z8
787LmQQq/K+uIt6ZzrJUUA8plzlle2uQBuEuXa4eLj/zsXaQNweQNKD5cu2P
AsiCDVlojaGAb/1Ot43+ygX9yCAXnlOOKjO6UtqUoqsuQSrp6+DVG94qZV0L
/zJV1kpWxAgeV1mrSa99x0PaxPoEAFIClz27lo6DrhpJP/Sa/SoTJNsrW76l
oQ55ffYU6vLCLrim0eFAvX57Ci4KAigs44EfYPdHpQ8h2KYVsOqoIn3oZus0
puoHBXlZtZdWCtC+G0d5WJnel+yrTEPKf58307Xw0F/sIdlKgIXnWcMZCe5g
lZWSbME1QtWKKWMKVRZlzzH0o53JzD9OBGA32RLme/WoFokwe0P4VT0CsPvW
Ij+ImyUH2634KqPZCraAKhtPylpua8VXAoOXiZUT42YRCrreXp0Cu1dBsIyU
z+4MRx4HvsSt+suhzkhGs6cwunb91Qnbw25zJFyz0w5h3psmY/RQWzyRhKdg
jUE0C2B9cI3EekT7n3vC3lOQCJeAOC5YRXQqAHuZICAPv0WsMYorrcDX3hXT
ZX7NkiXSyce78ffti3Ann0lUFMPuZMqkaac3v671ri1SmTK5fxCVRFZxwa4q
8wNzuJMmUoxg17qwbUCv2BWNlzSyao40gI2iEugLlCE88QyoSaCIILu9JZUq
P5IGEG9RBiMZXya+WPJnaIpze+dqndSwNg6NDAApDocUpj1+Ylvmx0T7wDs0
vFlc7B3lfgSpCqqoEUkdu0+AXeEN6QcM7vPHoosI+4Qt83gu54jpb7BPP9cA
lfOUqcXeXmKlH8VZhlJL3gUKfWFC9cLdserU3qKf1OHXx4rsylJgx5rOuZ88
Tp7X9yH8a1vZw8dM7hveEaXv/rkYs5uUk+m8HMcWbqpV012AJcZl4wtHl6tr
BjNNuu5yNvG0Q1/+43t9MAElqGFoO2seXx0M34pZn4bfrtMHjDXadtUkkDi1
EGK63jsCljmyrxFl7dlJ8IuZgrVYGh6xSXMBm7K4mqkFn1fTKy2779R+U0aY
7c9G76pAc5ZkqoerSsekXHfxWnQcOrTqNMb6L+Ab56/Le1bkFWOBiJRAdTbu
1cCW+ZgXhFltH/ezwI5EvS31vXe0YeY5T+sbomTfJiC8MUIGZlQHWraH3qAT
bHBzyfHEGiqJnxIgxHRA3YvtNS9pJcqecv+rxL5ORRBo3et9ZZnG3gS0+klE
s7JPFEziw+7AxMBcp3wQhe4jofFFUqAwTn0bIJItW4gtV7FoeNhTXMv2jr5/
ffiVwK0Y5e0+IKDfjYOGhknZHt3Oxtp7n/GGZPHn9itjiquFh8EOciSyAbyn
sUzVN04DuMsX46rOnLZ31cfBgQ8Uwif6MtLln9fsAhPw7gqOciLaHvZ5RLF+
VIw6y8XncLruNXd7rtackj3k2DOfTWJj3YGXFs/TS63FkrRmpOYE82FgKvty
OeNkuzmKvMmNOtNacNletqa9ZPZK74rdc3YdE78Gl/OnbZbs7KZyEpzPluiW
57vDpBEsbfelo19QgvSB/+RVsW/XytrdTWRVTrPI8Ij6IOrQmXA3D7vPKZ2e
EV3J9jJ9lu54fVEQoDHCR+cyyk1QW40qZAAAblXKhXoE25tLKJNuw6Uz3hDo
th0x6F8BHD1nzdEursNcOHr1ltAYoeL0FJtCJdU/LzJoaKhcNzNif90b228I
uzPsVI/e85yQlXBnjX6drpkBBo5+5waew8AzeaNW+OYZX822otZzyxCViapA
3TGaH0+LNTQ+kmudFRFyMvmA+lOPg1o5J9Ye6ViS26rEilCY3lsUQtsMMHZh
CcBL46+G6mF71As/tqlOJkLoNOxU+65X3ODuWLZMY3hGRaHghxTGAzhPOEBd
yG5NvR6g/+44lN541lmmegefyx9hUrlyDUBSIGGsXp2VSbi650Tez4ASaIN5
zk1O2daNRTX8jh7gxt6ME5IUkFaMF14xXQn+dMy/Z9rMBAAZ4S1XDLpAxKoM
FW48msDaPmuHXFDbLO78qE8DsVnCFgCLUVWj1l7XLa6BP3IuNPRGFW7G6BL5
glyFPQFagegOPAi2j8A/Y3EhndSsnFINnBlvDhrICPP4rU35aP9r51YCUSrT
kcmtbgr62VjIiLW709Ef8Zznpt8Ha55eSPMJ7XqE9Xim1w8g7V2O99n9KaQm
wM7M6ZWVO6cwi+QNbAm6m8OVSEOn1p3ZnMWoTeqJ8qy4LhCo5ZJ8DRYvgbEb
xJVNTYsD9MrG7EbHiwI3DHBapPmU5Wp7TN+Q9YlpHza0qJDrnmUoCONX++vF
Uj8Jm0fWjp9b/jNO2rciPmz4luwO0ia+HK9ARJyyhoO9Jc4iugneru3JsBS9
ItyuURLx6BUtDneJ5EIuwIKTJQKpGItEKCBGbwNqkSpABoYVehT0NHr7BQrQ
yeVbe3vFe5Gho1qHQBbYy8aALXQOap1x2HvEBrhK3L3bpOo7hsBB60jQ5iir
rtB2t5TOVeB+OqrBBx2QrIwiMbWaZURdiIGZZUMoiOrnTdyorkS8urmrQXc3
i3puFaWFHdon155NzwQiTm1MolNnec9K4JRYP5Yk3CarPijGxXsMkKV/JJjJ
B8m+Xu+B6cVRSDwBiKfcIl6oZsW15UYpSbq5q5Obn2ijGdQQbKkALg0XwKkF
CWz7Af/PHAQPFioqClUdP2tm9wC04+EpUrqNr/4Ond+rlfW8xYrV5y2xpWsF
x11YCjKAU/s11EUhhloT3IpeNZR2JkirbrMMjJdN26RVBEtAEvS2G1nByyyS
LxB/fPb9QmvlKX/JY6I8LmlrpvmPxW/ZUSlJzEHfWykC5I1Lv9axOctmTz/g
ErWBiTujVyk0Puvo27NwxNsKyL68ulIPF4+nu7WP148QooM5ip9MYh8scPmJ
vv9TUZIfbYjfaogdbaC0ob8J9SSYX1WElKipIhEliOT+mG/LnTvi3ExFMhfW
N0F5j5sC7IwTB7edI3O2XixSI4nodGDXCPH64IhxIwOQwCCN+3kCuAC0t2wI
dgtnDiGseGpUM1LssA3bM9LL1AmW5PotkZG2hmhRe8jLdDVzqKws5cnYD9aM
UhWBNWzWGUGwGLOGY7RT+8d+2Gsfl2nkCZhnLTXnJRi6fi4MDE8aGJCovMLd
r7TDpyCZbN/luZ5JeW8xNkJ1/NllBoJeZ82ulr1f+1SlOzLsw1zBTzuxCN/R
sD0BzXOYcgTAjeTg+EVYd2mRsy9A89HTkxgvNWMRORUjZu7RR1oCgepBa1dH
27q0DRpochsPiTA1R2jlqoPaGcx5M8Ms9r2bH9NL3UF1bK1Thfzzh8kIF4Pv
M0DF6PLI51JgX3XbffHYfGUs5454sEJc6D39MoAYhX3XE2F5r4auqjTd3ZT2
Tu14sp5Qb+MiPW2cawfxP72xvq30/ilmkSNHWRUSCM/2Sa3+3GbUiYN6IKnw
4JL2lPojvUpN91eRnVtLZz3jebfpPOP2/r1jtwEvcW2ZMl7tVcfLxkgufb8I
0BwMAMm/tetHAwGiQo/AFisFhwEv2iCliqRbWuNdktm+ZkzcsINIGZ6rfc7t
8zKS0N++C0bmGdkZnze38qv0kcY3EZpDC1JiMUIN6kjNzc2D1gEPgIjAFULa
ybw1EWQTHCUEySWb1UKUfOV6HlyXg/7fKNTVStXfLF/uvYEyNqkl/mX4GiMw
Q/iCq4w+Ikb/1pAc1VGWuS1kGS27AqjdOo9WimVjvyQ95b/rmY/SRTRKlqKw
uNsWXN674M0cVCvezfbATNRDMh6D+zwDARftY1yNqLy28DG/9SpcDLZ9C1Xf
Q+EtmWrGMlSbZ01SZfXMb6Hog3JtVy/z+zopGezPjrC2nsAx/7q2Qu7zQXAp
oih1spSupl8wmE4iHyt2nOJ5IXNqy1SCJuwiFXTuXbkgaEaDk029VfOqe+Gg
HclbkqQ+cp9L4GepOSgV3ROLUzwRtkrDMMi3jwTmEbzeDCcsPI47N/28riMX
jxG2fXBSsqsVd5/f+EjvJuj4AdZAtzMkCZHOR6M7esCz2dpyuZRYyLeMAn4D
TX9sTqV5x6s3gVuxsg+vPSLjfuUN1VOuEVTUXLYzWzMx8jfkuTHj9cYmlWs8
BYTdOnCQwsh7kg39pE01IhhjfRexjlkj8ZoRviSelIHX9vyf0fFPJMazInV9
A0st7u9X4evPErRQgvkfY6bcSu6zdcJIol9Fvzc9yGlQ0Ni6uxkpuDb1o6K7
KUq0IQA4WFidp19BBpBiBhMX/EkwlwpEZGEEukvklWpwnJPKheZELKMpvNJ4
xSuwjcXpMbVaxyn54Y/mL0/DFmxtCsKLzB7DeOIW2JwaIVv6Ir17cWjQifZZ
JvLCYROrw3D3kbI6injgPkJHWUdVPVKjkAV2AR06VvRY9XE/Z+0LXWFYNTvg
zQbPvetr9n7oRYXClrSAv0Kde5OxFy3L5L1qUHrUrllNs6od24lxQ/47b2RU
U4BCYLDphgfX4D7CEyHjMUvBMoRT4YmjTqfKwjghjPR08+EN/3AkhfKfz762
VzYPIXZ9wPRgN2ur8gF7Jpj7w+EH8kHDM7r5jcXXinV0O+DppVCg8lwdOw64
vtJ5ib6nfNG6LkshrMGNdRVXPpoXRqtQTtT9uz2ICf6J7VkbiyBbywSPTgb1
9qKfBrdUwhBn3csls72+4vn5bKkcKWE9c8+SwLUoFyrRykCKT/vStqoSuREp
JcFVcHzHRlXGF0rq9y7LZpz0QZL3vS4tNioylbTw7bpsCRNMU8LMgCL3WCyZ
tmbDD7j7M3tDoRxoFcNIyic78pPQXJvqPp5twLrEfw1lPDDy6+iwSuEA9yGP
sGq1NUgHgDFUDHCYAcccWv+1RbF0uQgifKnicAjq44+30mUcBxcIhG6zybPC
E+uQnmb8mnFMaNgZvm8DCY38l7dTIX7e575eNKTzZwkLomgUpc5PNC9lLc1e
ZTIHLgU1MW3DZQFp/iiKy5lEs/WD/2352NcX6kNV/oBbTfXRxl0ipSNnJc9V
Oqz3qRLiuo8/vPK047uvqjWl+6Ml29lJWmy7qSONRo2QuN4artS+amWuSXd2
S55kQ926/ZZHvezoFUzb0a3BksdN9Twr7mkKCHykdrizx5GPOppkG41A0KKQ
u5qIdk912bxUpSNnQdlyltx10SMpTAIAAk2ss+asaTmo921SvFRO+lLk7SBB
4G8SEduO47KWiNdxqoJrEjmdqED4Su7bQKfLrdopuU8Tg6VZ7IHTYTM3UMJe
iwyfqAkUsSzK1PXPcMAX06/BPDKJHUymtTXr7q5CQGekHoEEKO34/K1cINZW
uWx6NcdDTE9EDkvS6Eh7ecvYb++sghGcCL5f356R6NojcRuyfW02HDoDvdUC
+q+AELXp0KAG+rQ1d3E+CaWWi3OpwaHSiFaeJYb9wjQvMZL6agLfGxjowXpf
GQElF2q81yN+cuC/VK9qqg8/OXKt/r4sYWIL0VMg3sOv+ypfvL5KvEYdFscC
ZW4jeSSGlhi/xY3jF9DEmaYSwY2V2k+nXm5q/5+yoUuLRE9qCws4VrowfFZf
JW2/wYwBlXKN0Q8bd9hoARB00A5BB8BapdssDs8YbjL4kxG88bPXycZkzmxu
i8tRRi4G90UKyi3juukvmCuaTvtdZC0AErY2qOzQQLOZzr9X7NaL96gbKEYj
umci7AfBJyqZXEwrp0njRRZIfu4Yd5Dww6RI2AwmcDo92pqY0QxnDjKTNUko
sHb7r/OyEKbupPmc1TcO4UfhxwjFCpGYk319WtGzNCsEILRjfG96VV3JGAsP
ptjQgd9kf6rzQtMtRTIkzmFuKxNdV/lR21i96wT/SJmAEJWAOoSMhOnQVo21
Yrjp5BRBMiMI0osBIktoX338B1oyCoYY4KxM/I/l3HI54fYtU5CtrFL9L2K3
iRSBe40jRBAkT3juGxotlZEfvpu0cPisMmBBR2NzMQEoSZmh2OKDZXLP7rCj
89lneAt6HN9D3pKE6DGtJC/NSleR5CUca+ufMY6EdCVTBh+pX962jCUm6f/g
fJnCFsOp2wlap6ROiXFab5kbguiBHMvwz60G8/PE+jgk0hNRJleRbjf1hwSr
ag1/KzeCXrKiwa6ibaQdR6+0L5+bj8hW+USavfkNbEhfl2fbpKE3Ke0IwKx9
AJSpuSVuns0n6d7Vc3RRU5+Fe6c7Z0qn9tir782KaGjk2oOSkRpw/pneeEdK
6a3/vvzZCs+NkUFWQszZzUkDnIdF5Q7NezT3PI+yfOfqc9AnXktU+64aoMRj
K/8CfRfJ8zoWcxRwNEpJ5ahuG7Yl9acTkyzCjO1YKUNk1MRSHF9oVb5qSuu4
7Wtgqphqi9HrBeP0FYRZyF+ucPNh/Nc/cSwdQdnAdwXTtO2clm4r3XOuPD5j
5WaLPmXm5yyPXSbbwAYXuEEef28XR/FJ7BqK2+NMMlslQ0/AIzAWIyyeyL16
AEzNdjf1Ggpg/Wn+sRLraql0D8UKT6xOEtHL89qNxADs1ImXPoyCVXIuX5AZ
Js236LXIhBYSuydkysjMk+aRaaixWDDtZXEDDVOhWCGHPoIE3BvGjpkDpoeh
pL9hHWakFxJhUF0bV+YvQki5IuT3j0Gy7MF1i2kTbvvTT9qTEB5lLv8Fk8uC
BeMRmGXZi6ZMF33pNK46p4z40uHng5tAI1J3Stf5RLTRWih11AfE8g6Gn1rr
d0WwWk4TDYkznPd+4w/guZhATLSiDsxrNNeVNkffkY5iMKgql13M1ujI4Owz
IWeBf977WMP3D4Q3XVO4D8ZEOFpC62i27jdItbMaXZY00jxozFr+EAKw5YWw
VWYZZ2j28PiLDFkcLjXiACtEOu+iTwqW39cDZEK5cpuwy0soTzcUuiZ2W7H/
u//lX3NoJdfoeZx8sGyUa4OLepeH6HkC3r5UpMHsC9dkHzyz4WoQ4j/fFH6r
8WtSvnv1I+DxN+oJU0gjm6WgxUrY8s+usOAuJQQuRPN32WFJ7doxZVmsn+1m
alAEcBhkN46xSHADeHdd1xHuWzDBQRNgJ2CLj1XCxuBhIlQfVm+uE0o8am0r
N6d/IBGHNUK/yZnUEsjEVWZxs1XhyeRmkXl0Gqf6KSc5XeLBR/Di5k2PyMSc
nEQ07/zzJM1pXCoMucoxzCffFFAIdQFXM9RquC12lV73ILigg7U9nqOYwBkh
GjxHqDtAD2YQM3Av9IymAcW7LwTVl7O9/tHTuo5Jq2uN5s+B6TtuTO6SImI5
f6G+8kYKzgFRpnruGJGgEuLxrUcjGr+EX1cvHjFr34iW+uc+TrfEFKFbFnvm
hoNR91HTvT0mHQlnc+0SYAsZjeLG6/Bmu1DeuIXVY6yiZc/FwYCVokWV181J
jwJ9TtRKac7xIoynXl006edZglDHrGr891T9+2CKktanqmy11MjUO4095h0P
VYQNbgwmwNqLm290lsUMEqY4hRQvUFwPyEqx7ZRD/369f6MRRMqk+8fMDe24
NH1yFyvgzJKFBBrnhXDUSGIXEgRg6JGL6o5XTEtsr1PCyGbPYZeFCcSa3/UC
7vQgGcA5wp4oO3AFAhAyEd0l+bb9tgnJMiX6T3cIloIIde3ACWVllnsvNnPG
TJkq68KTC2E8+eXi4D1YdpGK4Oz6xJzIeStrcQvtXLL1UQPZHQRNizvnZVOY
b8sgGCn5mvr6I9nGSgHoXtN97Zd3VDJ5e5Dbd0S/UkIw6PSHYTv+QLQyrEYt
IIinaE6l80Sv5ICg9/vqibYumtSFKRr6sIYUfSstrEFvufLZHZxrLDowly0a
/D3cuow+kDl2C1XvnzPrzxtY5sGKPSE/Ee4ue8xEESOnBI796Fr672C4UDMq
6V8AAmSJMlKhXoIRy9eHcB+XUEbmAc0duadioBMvRHDMH7qc/Yfsv14+4jJX
GlZNeJvhwS7GH4sgbC21Pd5+EASvQ6lesjeiSE9eBK3coJHse9UNEUFZw2R5
yQ16XoRm0yKya9NyrGkU4GjAUqc8Ql3WUD/D/BlP3mRVp1SJJrkVRYLEM4Vs
FV/5Y/pN6GlWD7ayVhKVOyEiz9G+BBqIzvfY+4GnpxeJoxifI8dBpAuNAGDc
/lEQSyppbP7yyk2cmNDjBxsES2ZaZ+Pu6Cd9IeYpUM3mKcmuLqyU2CVIwqZi
YY7xQOiP6WkGNsSirzfsIsqh5Jz7G1MZGtyVx4IF+aSWazi+NSy9vdeAcaJT
gPgbhwBW1C6PSgBbygq4J5HfKzobQpCSIK0clIUgjdY5mKQkYruaq2LP9OTU
ZgFso0Sz5JqQ6xFERqFT1SfglFSRaJMAlBcjjTrhwogvsq4+eul5tvNZfwrK
3MMTIUI3ugJCXyATlZ6/9cskPd0afcrGGHEFTkAnTIynvP0gFrNxCv0VK5sS
2SDZoVJUj2SvZlaUyziDG0UFgGJbc3Daim2yay2NhyqzSRUVwzJ1FZgidu8D
bX3j+a6ohXvVCrLZGmMuyM2KIjeuIRqXXOsmNIA5SNoS23xCnqtpZKZhgIIr
E2mieeqPavuUhNPT5SX744Ds+/LypdMdw/a5OkIU/xLjaTW5lgqd4mnC1zYy
aYdKA2JY6cQL6jN8nb0356xy9sXJ2+kVsKM9G0PfgkCjJW3CyDUYSz+RcmVC
Ay5KrC6or/h7SdFtVcPHQGpAS0yNcjiqncdPn5B03y8kTUYnaxuADP7k9WRX
5TGW+Q/4c713BNeDvG65HmNzCDDCe6TIRaA6AbsiUPH+4n27ldZLyE0kgyMG
4x3R/t9ao55Jqpa9kZbO4JRdgzlDLl9RF2xBvCRq31jlYyykt+qZga2DCyBP
c68DyfaMo8iJqsWFfEeJqXRAGf8qCjY5YGhk98KhQLkX4YjdbSOonriyjxjH
aQ7C0p2mWzfvMArCbit0KoUqQb0Y9hYVZGU7FcJPi/gSiZ4I65jqIjV3ZNio
mfJkBWTKHS9CuH2cn+7Jxhd5b/ZCFoMYcKMqzhW7Lsa/ajTOSbMlfeMpdBaJ
Ya3mm+qnWbDLfqT+Z+/cen34j7xizfFuGpeEBY3INaYjQ4A82TjUYYHsPkDN
QVrKEdCGtA34qkZLSQMTNytGXvjPlFJbTFtUT6k/m5h07R382ZNhySzr4A0+
qRcAiUcW45uFuV4caRyjBWNrRDsE6Xitn6wnU6HzIwpMRzQy+1u8YGrc6ZRB
CbfZdnQkrhEZefp+KLHmr1jRJueXsO2yfNwGSm+OyPukhotDMEQqUZUavDpT
DJe37JeWvJJyE9HXf5rtpAD/MSOf3/OqVXwaus1PYzgurk+CWnOxdFPa54fW
SqJwPHvm2Z5JcCoFWodjaZ2bkZAwlqiQwlpHOr79TBMWeCsr9meRe9JxGkpk
0KFP4a37gSueF1bBr4xc90a1B6PgRGqJKhGGz+L6SJkbETnfk/b0ls/vu4j7
puTHboP2WWU8mhk5xPr9ag8316iDkrB8/I88nwa3QWqHs979tfF/3WuJbcz3
HjwAvU2VDaI7POs1ur6IgO/pea4wBWgS6mLfMGmEgxmUOhn0UeD/VxZ88lH7
fcMF4dagYJhYUvj+h3F7+r4oeyqrUa0BgrQf9AfPwkXCZ1HdGD2TgBXb+1AG
xI0b4IezJ/eocs34VwimIsFfZ7nrCrqyAeJFhzi3G9h3trwgNgk30Ii8pVoZ
jouU3Jp9FH26ckI21+ko8jpES9v+gsCaclSUk/AKnAjwKIPypNWZhri7Cy4/
FM0A+uSH5ImyddZpjBmyixl7C9hnxn29vccUkecs8mf05QELCdbJBJCi//JT
PVR8j7XbjKMoLsGqmqDtCHwJT//9SDHgive4UL+sJRZNH4PVZGN0rdGz+/vt
ZEO9SS2HhdGnPTYtXGbEAECb47YPaZ7qN6jt225bfU8fDYXAOHzP7pzfd22P
UKOR56y49fFee4ljzIPwC6nYtTsrdRTWiDNwJu+ac0ok+0huQ/bniU5ZuhdS
UooJSXHywhAo1O0H7v1ynu++qi7b498WtUunoBMfTaHcWsdCaYwUqyQJ27Cf
aWWfviWfTX4KWI7tQ5dx3bZ+gkVIhvE6y2O8MQwImyio4hVBzIW4QYb/jcka
GmiuTYjFe6PwYSq+vbqrdivfJY37Q81oL4Erq8GCc7lfK/14wulZByzXGizm
qzCrftHOPxSirGcst9eYVzq/0Jzgw9twI/UIrpYM4g8CSsw3M0LUr8TqRh97
YvSVA/84Cp+pxCAzFd+dZrdhV1rCe+qgbdfcqRXAVCX5DKN95TT4anOD9FJe
hcz3f95kp2nkumBMRJ8ozgcCAXs7U8z6305ML1YEjlXOHvUoooEdB3ucGPNi
A6r6y31jjmiKveAY/Em3wqC4Okoe5mhUpdnsEmY703AQ+SbNDiT9pPcGy+MV
GoUlEQlBTSH2yF/fpCURpsxUKSAQscSM4MpcPTqV6XLTe041VaB1cWUpVX6w
CPNVbqynK/7aTRP1IOCxjZCWpj46+E10NdlfhVmXlFLgD8tVIlLcVFahP4uE
uS7473PO5WYGNEI26uvqWuoDK1IJwwACFNZ4ONjpf8QPVa3RYd8kNKoQ1lS4
OLCUNbAGqzBnehQfqLLgEFV3SRsuZwxwb9xtDo1WzfA8nTk5PH20mWtp4ciO
7gvYFpPwo7d5sQH9Wztjdff8lKRp0340qRRt5oXUDKkUPdX7G4zOBd1kHN+t
oE9ZO2RsTtn+8qwIj8RrHuKL+n2c2teBJ05cxSZUdmuvjYJgwqICgJ53sZr3
BE83W9xSeK/1//l6ItaWzB/kalhEHDIcVtzSle25vNYNK7PIAk4kqa2PliTs
0Oo9Io84oTljGMmb/2c+PplbMTAN0DsGKXe5+M9cRjMlyrEfmixXfVYlt9W5
NbcYGjNilYsS8b2AfFYmoJFdpMBbduJnFK8hfoFjUVpiE0L2EUpu9JR9ERHg
5rDXoW0dFt5+MpzZV28iSm56ezYLkpVSMWtL2zdCuBWU1Va0DGQ2p15rCOur
avt2hBFZxTaDdKHwC2hNK6WwEacxlpfOaIfP8m6qxK8Hp1XOxDrA34bO58dc
syCLwJl8uNJVtUNXJ5Pw0qAaruFyVYVdiMBC6+sEOfMUpeWAKQJaODTB1BbE
Xu7NoVWkkiRev3HAFCFp+sR+qbXl6bG83YAiGl8OkaBqutHFUp7yO1PUyuBC
uVzCBe8OwkrWE1Y86fZbUIo/O6wb+nVhaN10KhPowkoe2s+HOOv9vZz/xzoZ
Yag+xKxV85/RMbA8nT5tx0Td2/5/U0r1zGKFbVi/EhoaKW0AUhJ10X2eRXyw
+XysUFFghDM/s3tDtORVaaA4wknGeHODsSjXi40PPFYvnU4th2pYmQyVY53z
CYIWqsyVIsY1uFbVwABENEnLUFfjuHzQa63ZLRIorxAZ2UaDqDr5pZC5iIt9
FKz1bFXwdAa6h45eoS4XDti6ux6+Ysi5B1xnnodrkXQBpJhFR2b7wYNiflEn
TC5xTZKFCqUwXVd1xdKuYOFIfUFhqdltYG4faoLsOEInj/9gYyBUGb/oSbVP
KbZoGnyyA0i/a59s2OaAqrUAfpikCm+Uvv/Y0OUtyK+raEPhRz/Ol7WYk5gK
uiYLDoDTanc4Nq6AM83LD0pkAotaNR1XKkLYJXf83TeySfRrHPV1W8I+3oXA
9OLdlRSukq/y+RrInDuL+Yhe9ynfMCEuqUQe7uyb6phN7WidDBtZMaCCBQpI
twbv+Wt+EAHmmlQj1uINZbz5sAsfjOWr2bcHWS97qTAmhd81mbl7Z7bXtGB3
IsJ8FIv1MxEuuZK7dZFxiE+ELTPoFjWieWIdurD897Ah2oIAHwYg082DRZmY
d9mUzxGt2TSL6+lgQ/Y6qe1dxMbNql/09niXw9XKdVz4yzaCC/18iKGIz0Iu
wlJ852SI9igFQbO5oCzHcnbzKf2bPAorYLxRiTtGEo4/zmEOurTzxWBBoyc6
vy1h5mAeHMSzuEcGW+MqtzkGPTOs3f2swcpUdqQYdXv6wqVzL6Wak1l1fP2X
RaNhXfhISwcnLV8hQ3Tj+g7tVGQuY3joOoWIXtACjmOKq2+OV1r7u+YLpDES
uCza879azJYI+hGY/OP3Qfs6UhirAawr9wh5M1nY+tcggn52kbnDNiOjNbHP
xkLL+2YQlohJp8n79lFRH7lJAbVXyEISHqUdr+afSY4BA6Qsb+99XO9rK3a5
Izm//weftkFNnGqAGm1LM+xrdFA0OgaDTs5emx2K/+qhCG4cHzdB0VA3VcJ3
V57BDvty0qV9d3NlN5/7yhHdk9m6N1hpVbgurrKr2Bqoi/7zsSL2tyznVU7I
CH6cFpLV6n9k44P1euhJQg+U9AATYln/0Iy7+13EtgEVYpjAmkAfXvudzLSE
OudSIX9rgPwKLEW3o7mW8Xq/ZwbzaB46Lu/IqdKWMXK1WMtXgnX8FSV/J1I0
6qrnDZohqG+5FMTSLEFJYJWiYDs95H/wxiLKJFwyLnAsxl5QIGUpQ6V1AKVc
no40MMenSMBsBBv5Z96dtk5tmLon4m5pxUbFEbJBa4Pjg8rZ92RPRuWljeMP
3L8Hq1dmdN5LuPIWNSWthY4F/lPCpzE9bjdWYaDX5E6zbNOJH9XcaL4kO2Qh
OvC+pxJyVFN2RkUmVRsQJrsrqzOe3ko1xtgeEjsAqG1ROUOaZM6AIqnaycRy
fdfiy+1luSSX0gMC1kbxAs6I3W9Lc/HKK4ILYc4ntzRWCecVRV8AOydbzmwz
XZMk1Xl4prYsNcK38u20TvT9eb4ARkxn8agfkRaI9XMDsXC8FyUM5pY3fTbS
EVU1gfQGB468aF8I1OxAKHJnDFgOJZsLtm2ni1XilLHJeBnqg/UdwXP3yi0H
u+BNuWwPYfKsH7HvOxPL0KI0Ua3Gfhe5Pe6h2GYYGGA1cs71AVoLgFvIfsSj
Udk+OFfp2iT4tR97tT0F2AjdoPYj+UWMFaKu5CJkjOgZxPa1aa4xMM/4j6lA
KHM5CbiGcHASX5gnTbPCfPfJfL8o7y8a8n1gH2yWGk2dsorJ6v19Jx1PMfBN
xNb8rICARscB1g7VjAdjs9OH2DgcuBGlUY9MEY7PSQHBgd+vGPHIQq9yR5GP
+f7Q8P3gNVQb2tB5nXjTlsbUIla694UEvNYGnGTxS0U8dMYB+Y7NMaiH0DtI
31S1gimLNkCNZl62qHyyW0Hpr9ndSNdtFSDWRL7Luw/DG23aGomsoe/sVFy1
+OQGvcUxb6+0nHpS8UuULPzbfdXfJRahmjwH+4CkOlMztptsFgR5Kzcrvo81
q1ar0gBFvbGKU0ZcXyfGu0OClSsUOrAMRc3Wkb8HaFUCmiBdRHe7P/KZ/DTE
fnBfNRpGLp8glXlirHHFvoSiBzlL7qdxTBP+k6aTUBpgIOtHGGaGi04UHBha
iJGTY8BUi23vdlnG5cdH9ndq5R3mJZTbMr2Ny3hZTCcWITfQhPeLmsBMnTQr
CnX5bhhz/evYLzxxxUYJ+0NzkFUAwvlJh0ju33bAO0R1+GyWSkyxhLdz1e7I
xJPc3J/352qxrCBPYjTJzikA2DR9J9Mox+uPaFDNCBmQMrP0XS1kqiNycW3b
kGQd67GrBjcfLfKuUECFhBIPxam8AK0toRtNRTPArapbQx+jTDfy9l7fE9dg
f06kB6uL2OzdCoIZ244alUXavkIfXoCPXqbI/WMYP71+KRL45SSg+rxc65Dh
ygep76ejyomnBFdIJ2qzJ/lekpcoPejBqp9hPbHnvJTWZsmCuHOTaJnvSXxa
viP5zY40NLn77r0qm1KXQNyAZsewedcuHDl1aJgrvCBPT7jeWLB4r3HYtCoP
Ua2qXGxnHRksW4UEGynHuyxmClpbnC2ztxyEB9A2CNcSeiUedW5Xk4/hZNHt
9jwAZ+3g3Ucw/UZdneYFn0LS3izif8LzRlWs7rKyqPOvtyt6Zqs3EphbDZZI
uB35gpCwaerNdXXvoonz1iFJH/3lDk03Jkb0XOz/5sqpLP+yxQH+TTbbclvH
0hejULfjAEPq4F0qpSlVhqcbAEE2Ma0coY78Sf2qkexqb8tidURjtQ3Q4THR
mmQe7uMOLfd42/WqGxaYEHxb69CWp5wvecAQh8/1jfkfy9mDvzFjt1/28eAr
/4UfACqEq8f5xwQxFqTm0NvO24zCQGCBIKxGqYz6Thi1QB+eiQnPtVv4NUjj
HU7iV7eQBuTmhy7eqN6+BoqBz+LmTFIW1JhxqvwNO0BNcrPmbU0UsiDYvdiM
msS7diNba9uLtW1LmXVztAi1nY3cQzlbgd9XGf2mVWZAR5tdA0HB1RWHH4kg
0J5XLI6+VW+0QN/SRitciLM8VmyeiznppNxBIL+BOa+gjix3NOzKSL6ohkQ2
OE+mHbmQcgQ7YLpyo6yd99bDiBBHxN4M75LsrJUItnFUZJN3p39yJmTw7zVH
1htNup55rlzYi9yXTtYfpQm3CncqmVwiZQRff7fg2e0Chf14YWH7gAKtWA2m
opFKw264Tp7QUOp5q+XzNBG998qGP8q3WOVVV+c4iJz1N7CsXtZkJm6Omcr5
jyra0Ovy5QG3ds8SpnPch0IebwHLDto1gfy2kZmR7xgEeHJXjdsWDuQ78E9N
TwtcD5VJYZl35NyvvyuE3c3CrYlB2ka+eDuQgAzRIjhekKZM7SMszYCqVA0h
pQgiFFzm94r81lH3tvdEiFFXkQ0SGw/AxMZOtLoDtxMONBfYZjoqtHCXs4oL
zLDWSb+eAicK+H3k+1WV6SfC0kl82pcUfO8zk+oPgGapnQ+ghy8vgptlxspr
rQq9OILfShOnjZT/fNAM9BQj+Ozy2adUnCWynFZ7zyS9FQ64lH64icQ0niG9
x4ZFu0VLaC/eSgZbCHgySNGiyM1oKJGCat2/ZDj0VMweDSHlfDwsNRqd1CVm
XC2lzINYafrHqlCTtJ3YAGbIhepK0vGVuadIfSUnKXfE2lUMJ7wgai9X7QYD
371sBs/CUr7zeVMiFMJwP80YdJff+fNVpjscr/sPA3z9sHuK0h/JllhYjkRC
2G6M/06iw9jeVoM50hbBWqp5QV0XvxG10m0C9hrl5DBQ7gP/OQH2gyT2uN7W
pzZFmSKBNoLJbReJlbwCUjsaAqMxLdg6DUkwo+4hUCY3DqpFVWg2a/dQkax0
cLnfqtM19O4q7jMkWekbLmJQ3DdPNlNda9sj5CWG7eGkObiKo0oQP/2fO1cU
/2Hx1GnnJNks1Z/1hQLU3AxpZln42y0X6J4UdFFC1o4jvt3vpkWHYZmjEdMt
9O9GTMMCUzvYepG8mkigwTZ+vWsxYS2WWMCjQeJy3DMAcQyCWcQVQcLUrPAH
DCt7c7ifI61Be+DhjWXnZevLDsV6QhcoHcxGwz+H8N9MaxRFMaxVF85EtH7j
R+TquOwaFCN5IMsvp5cfLfsdkNbF/Gtvrbf2xeMR/Xz/3hJwjx7IzVmPJE8R
CTRHtxyySMENuYseGzd/IlY8HbnPls0k4PcRs8SX/xKklzjO78sVliGAuU8N
tSyN1lzAAfPkAr06/gLKBZf1F2v6do8WlXE2InNYA7Cnj7iFOTaNJyPy1t2J
/POOQF3KhohoLoI+1OKNeXM/5rHKBgyXI1IgfhNFyJxphFIN6UWopZ4xz6Yk
BfCLJxPL699FjDgvKv3cxrgr49j4Af/780Ku+9CVQJ2OZI2jfhUwrOi3zzv7
hJ9tZ/7H6NLKQSL6DME9rMsKPTuZ9UbkLpBGCKk51t0LAUFqf4peSkkRMo13
bZdMfmvKOwDz1xCTuqK7BNtEygbb0RysNuO/bm6qbD013HBC604krG6Kg8yd
efdXL2yU7GHZF55Hj+1nMntss5pn3XJKB7Bq0t1x/+gMeuwOtVqNLiCNm+T7
QyCVOF4K7dRntWezb93fH9qdlBA+wv2pm0yYSTelyIZe721qPKRvMbBzwsvN
ptigGncxrwiB75y+kP+p5PPhkmjjXHT1Fxwg3yHv1PdpHXtg5MVvZL1XvZYB
xP5zC8oWQ0i6yF30+OH8aWEjIlxB9wgoEbtK43EIBjtJb9IbZUFfM/SJZq0F
ju36vgoGvi2EiKvcOYtpvlzS5yVT7VGudWL7kIWGxO0hFhWe8QW2OlIS9nF9
HbIDd7yYHjI6zSwe/MC6PGk0lcRK8XOa88tkAYX+TZA4n3OA4V1LssgwCkdw
8LOVtB+wo8d+1C2Zvkj5Q4Qw10og9tcyQ8rvSZoYJl8BNPDcdW0ZEsTHa6Fk
e+W7JM0x6uAV04pvUr7KVre7ftrQW9hZiroWh2aqOLIZUfbpY9WTA07GPX9P
dVmmH5K2XpVwljgW4g6QV8BbfaRt72Sk5NwKDE4TjYYeTScxGpltEtam7BBG
bd/JHJYz706Im/a2DFJptEryvc7HSSXGbJ9mCqcwh8sgv+j710EgQZz8449J
3hO4/lHTLO2DG7yOc3Y9OksfB9Mz4/jMpTMOjyycBEAY4EzGKCUeQn+10SCQ
q1iN2J9jQBvjGtXqhkF46ZJrAOqhCWk4BpBZNbowsKKTv5koLHFglL9oRH3A
hENF6NedAguGCRti7t/9+6LfevA7oDw9Mzcbxo728zEqUWHgI46Ihjo+SY69
Fb9Mlaedma4otcYl+r74/Jvla2xqn7bix7KOKOpOxAPCNFXuxQllKqimARPE
VupypfPtJFGRyzX2oFINw3EEkUa7XEow2bQ5kBuD3Mk2Ee7SGmda2GHXOdje
Y7NuvPmIAXOOJC3aOq64YDU5FNv1fL5aBGLhDlDsIhpjpaVskG2leJvH02mz
XJkV457PoyJSzsoRK+aXh/2A79SA37/crY3vca5sU5s+d/L2Ju69R1K2FlxK
QrFqbu+81TGGGAQpYvGfyXTlaE3XbR35RlQv2SRs9AbHPam4PhVkmGmQcgtI
gYIpqIOOJDf4FSBQoE2hl7ggYk+mur+XfKgcrsS0Ps4vaxYzaVZKtPTTYlln
8Rx3e+WP3qCSpobODFBFMhAVqJ5WQSPrcYtmYS2JOrPEoPvSzpX6AYzGmhO4
v1ijpz5asUzuSCszLpxCpFiJpHYWTABc5YALu1lL29Z3gzfprFX4uKxulmjp
dLxtlDo7VNfVVmM0oL9k3/kSB8u4X6Hb8tMm967b8rlBHj4B3mxWjD1TcLyk
woTya0P5lYIT/OLJuwe4B6Ptx5sBVvChbwdzfqE3MMWGuBuXNkxMfB7SIsNj
rIkJ5udNm79rQInHRsT30GeY5XYPqw8cCxG9vEpE1PkXKdHxbH6TKDrVSOJk
8xT2Cskt7+x5UUn3G/yFz4tKsGAFX+VEBOys+Os4nwxIVu0kP69MaZ86rWRf
7FQPKFAd/Z3eKtlTBtRnO5M0C3fjpFLVQf99W3bPw9ZRUR4LOH4fFaV5s/Cn
leLJ8E2nuKcA/690mrkwOXcFJ7c0mjQ0vwLvov2PxFYSQ72oN27Hg8sHfr4G
+8B5wnNp6PwkaGnsxnGhtMO7/qJtqa83hWbaQK5McCLkE6WzzTqa1l3SDvLJ
8EZe9KcR6o1JYvNmnMuSz6nSGiQlFXvG9Czdt9+27lZIis2bSHnUHC7XsJxK
ajrXAKBS/Uqcsles7bzjL+dYTYHNSCuVeLqwzJSPKAm3te8O0DhtXgeQtoca
ZWGmLYtrchm7l+w8AWyeaAeGNSnrXIFM38naffd+F9BYqfAYpxWe49RCg0K8
iuHF0TLvFSoQN8pgY/S5EWmMF45leLxZTYYlkTDwdCqr66xtykuu9nsw9arh
jM2BBg1AdbVDKBGVd9gLohtUrCThoOtM4H4xwjzu7y7WBsSq7EFkV3z4J+Wt
5zoo3hGC9PEe/9Bgl0tKygXF3AHZJhsApCXqqHNb+Zt9RsO2hNAjYmA7EDcK
fcFbIJ5KoxmTsX3NUorPBOYEjZAr7O75bkdhc8COCi8asOVBD6XAAVAiBYBM
tafIRwtKlbj8/inXG9Ld5swgxwIgYgTb4UtKZSo/PjmtE7yW9MtE++AmVGUs
bvvVCBr44suQfFq8Z94vf3y30V6gGVQuyCPfPgYHFevcoIzXPr5U7adMpDR+
UnLZ1b467C9x/IqwjhptBoWRZh2CCScp7d4/QFTfsS52IwjhVVftEI+DC7HS
3FUKZK1RUtAai14mCz3Acm7GkyPId19WDhKV/eWtgMUpmK+xiMFrfP9pg55o
xTBvSZCA47OHgyQSPPrJtftuZXeHLXw//igQhBjfGU/BKNZ0NRenM2AOKsKQ
31w9gHejrhw8fkAv+3+v3lJSaMzNh0ZFvjsrIqrBK6IH29QFp0sRO5nPlxW7
9m+QQhKfg5lkC7/+67QQ0/QIGyWSjPgploVZr3kcHTLK5+gcN88AWrJ3pJ7/
xle+NgW4nf/DjbmLiXp4bhk994xBb4kxBuulEOPPQ4zrG148/8lKs0uRdrmc
gBoplX/Ub6skVO94icoG0D4SMZl31uiMWVf2F7+YE5G9bofpsPTq1ylC0Zkc
ImvzS6AfNt9tLT4Jew84a7FKsYgwr0CRgaLqduawBA0UcHx8dOWMws4qYTvE
jVM5+2crK9phfNXDoOAk6f0Joy+uOaWz3/uDhPl/mGQ3PjjSOQ9BotnCRn3m
tlZAtptZu9mZ9luMQrdmF23rLIs2fJygtduYOYnPOY6Kyhzlryo8LPqe71Um
qpcCAdwBjLa3zcGXW/e9DwrOpF/xF0CfrI9MhzGWPoh1Bdd5Kjqg4ushaYpU
bdN49v4H/pd2/vFXLA8UaQqEvl/ixTdRaJipPEyOWtVaoxGpNRmW8WgRk5z1
vyz7gLZ8m/Ge8/byeji+5+GQsil1msac4kw8lqMe+YDfIgvRIsoLpfOS8U49
i43ttmv7tKI2WLI8oHU/xx2kUEpeaNlXbwguk4CjrSAqgaQGT8PNxtTohYmq
+EgNxToS2jtZKsQ7uDjop17UvP1XIALYA81rrsmuvEN2EYF1uqy0TXX2e8iS
5p3O+YUWiZyP9dxuU12lwA8oCFwwSSGan28FofrVLDgkdxSsgfpH9NtxZFaf
TkpW5aaOvrGOHICTA/T7UcKldk6gFDJ1a6+hvoA5xziBNB6U10Ctsmf7u38o
fvDB8C5IEjWUwVoIMRWpr0xMITPrUrvXGc9QHHKGCmiYDEfhFlmst5nBBCII
SdV2CHnaNaIMdgm4H6kS0TvJJvXdPjIGFoEkP2XwGaxrhDR1RujRn5QlM1g+
ISnAcAU/iZaZlOpMf/hachCa4bb82tT2d8Kqibm8qJOT9NdFAxYf8b9vfrwU
IUuoVKUOgHnO3j7Nc724RyvUXBLIpSjcxSkdUzLjblQ6BjVr5gDtBEou+RJN
RL758dXzziQN3zNMN/bUqZf5WbI6mviUQBQ5ywLR4mMBE8lRfzsrGgmvOZjW
yjE+nNq+JuX581rMPuv8nADklqsljACHDBfZU7Kxt+vSnGj/sWirk9+96tbx
IvWK1C/fppuY9wVgRRKuE9rdCUfepwQt5Sf/y/ynbxEF4x72tFBKweIiqE/p
KiNgENMqW/AbWp6ryrxY51j1F2fFacFbIsgQrUqomQRm7FmSxlWThEDf7361
RT2ZPrwrQ2HKHzal3jA2iplNlt3GDfQIZHhzWfRxrks7PfYaYyEZiDDZ4edz
JvIKntCmzLLrxxRwfJIWbas8ShxbK2z5ZtzJ/aBUEv9Rzs3FvZNCd3gtH7po
kAW/qjvObmFVG4tMwYhTchzVJmIldUfYwFAEitZGOcHrgw9DxNN8HI1M4taB
nVBFBt7FwJd4oxjrD30l+4B7guvm0x83GdirIgufHEFOYuOvGKD6tylH/bST
JMeT3c5cJUp7ZpTUnY3xu7L9QmKEdui3WYq+Z/uF5zHLa3M6kEm0eQWCMhLA
eT+4qz6q2FeuYpS/YwkaUBvqv8pacIEbgy2GP2Fs63oS97zpSQS7OMQ+NZEI
iaWWWTowxuCZiYu5/22iB9ZaHb6QvRJ02h0UC03OL98RVQmODYO5AS8/8vy1
1P2fzQll2hTsMpezFvF0NXxUabKHs3KWiTZqBZ7sCFEi3lVHzUiTZmlVDxba
/UQx+oNWeKQavoIlBOhcseXpWoPvGK42GYKMs1JHOXK+j9HugUtdg1q2rH4f
6VVbhCwDTBn4qazA3j/u3Z13rP9+bAmZ91rloSNG5+0/7asp0CBK/RXCmJtd
0IWE/7N4W48OyY2JSN/jyE5is6OXilhdCD9VdSAcVezOPkzhbFVFUAhoxo+j
pMvuqOHH7mXLTFwuWzFHQCWv9sQlqZH7ZiPLLsTrGyaq9ZkRdDXkRX/pT5OG
DF4HeuIl3qm1DBmNIqZMHVTj/Ke5Z3qyJPj0rncbjbdOo9HYRmoz7DCrEX+u
k0xrQXrV6xuxcfsQ0ZvFCzqeX5CGfmDW1M/ECgkXHxjE1XeyqCws/di1RrRi
ISkz7xRIa+MeDyAzNwLrvBjz+O0JzrcNOW4A27UDlhhhoc457B8Otx0NgrWb
c7zMiK4zuPDypix7Nti6Hw8QuicTr/X93hx/R8j36V3jrmtDxh2UVRa1L2Tq
g9y2DSXb9J+dkFuBnykhpfI75K0NLXL6HVKuMBW3xqJJTr8BpPpmE9ctXoiE
hG/V2Hy3VfWInogMNkyt34+tvoM4l2wEhQKebE2/cwmWpOmOgtW8B8CpoahR
RRvoULWwBy9ynvziR9Z+MkwY9FeZbAKpPn+jrbqvmap8r/fK96tgH7bzqn+U
iPMLSt5HvM3Pqz55RD2hUFzGrgEQ/QfQ/82Wt/AGsbvVXwBwUaPh9zMoHWVe
eaF/r9/mMLWp2z1nB7cu4IzwuFOXaMKxz5raBYCPfOGvm7kGoBy/xJ3lc1Fq
YeVhwD2I8qPIPNtJNWavSZ6LF6g9Y89o2Ucu7AOfQ6i5IK4X5UoMwNnqo+DR
VJhUM33QGjfst4D91R0DJDtE5/ok4oH85bWZvi6hzuVmE/tQKeS167865hWu
obhqq+JXqWlePaKFF0ZfZos8yy93dTG8OvOluj7GxCOI4Hrl0GhPEFROMP8X
EJRH7BUIPiktRdqLJT7aqJTr4tv/ILjkLIDvzpXI4HWRIxPG+nWp0hb65JTQ
ohJAmabjQKn7s536PXpoPGzj0C4uydcdPfKeCgNz91hiuLf0jlO05E3ByRax
pKjqZXE6/PHHQOSqkxKPrJvP5U1fvRZD9sam9GN/A2U82xbcNmQPbf6Lf+Vm
JkOI6cO8MndWYF+VWkORtofIssdo7rKyn/RCendS9FJUDbdSKBakJ3R5LFUO
yOGV7ez2KS0vJWL1sou8LghXZ07YjXk8RxteV+7ODg6mTlOys+4PemAOocg+
8Qzjvr+hHvAivOEwjLW7FuWccSbKAK3hePhSGx4dnHc++dOSqTzZOSTsJ9X8
LfnYXq9abcPHpmZo6oMYVDUxdclBRW+Y6tvDRKAy3zT1eKcARmLgD7VQc3QU
9bjm6+y15ml+VUXZUTwH2CT1+QU4NtjsygaEZjU56B55lqyNwYh4ELJer4P+
WeRh+xNyRu3MKKNKdWprlTGOBrmcEIH6ftIH6C0VSJ1VCtacAlY/Ck0mB2ti
2ESjvttUK1soaZ6oTsq+FY+oY84cxffOh925D/QlI16/lZmORP8NePIMoYM/
VwryVMljIkC5aiEXXSoCVkOr30C80iZlWZqeJM1Z9kq+UlmpaX8r1gKJEBBh
4Px9kaQe1Ju0s2pB2TjM2Tbdn/o8+RZh7ZIRh5fvT4pxXtSuf7hbB0gVa+Yd
UbpKQkIMxTf5Lapyk38hAjgqdT5QesBoPsMudJGPyjSK2bbdopcVhjV4doEy
hT2p6RMHeA4UGjncfM3sntC8lqaRV9YfT+k8y6UVRvw7U+1TkEvCk+6cMPw3
jZ3NgcKXtR1SnlPY4tPWyT3dMr13a1eT9r8ckuX3RWyTQPhEsVbdjO1heeB9
KqoDjgDndr+Py+2uhuVoXyRQEk3nEyL5NLgG1dzr0D5q0tlk+AR7KN6e1lXt
Wqh+v1Qvg0fDYK/0XFx1D8M0uxPoxNI0heuNc8gFADu8EEf8NnyNw/5xjBVn
e6vAF2xjOIoI8sfPLR3NYq46//AAPq5zh+ENUd2QcPN/h581gxjthk5g19kq
MLGiwTJxVC7XRX96ebi1cWcMqzi1GbUYpt2FopjaOiYfiLgpC+UgSBAHc/v2
lDa1V6AOkKE/Rk5DEX0SlKBTXCuxk+dZTQpKZoyWlnD1fIEAAKJUYUQ6NNH/
hiVpaVyh5D5ESYFov0trzA1ygwVy/WHPCie75LMM0qsCMs06ZPtPngRQE6Qc
RSPbKmLrRyqcHttvCZ8Kw7utY7yiYO9Pw1i+Bd1+yTAzXrg4TEP/HXmBGFi1
2/dGxQGP+K+QV5xflQvw727lSXAhiBqa9+4ha7jplRcGz58rPCJNvpsojS/U
a4fzylXDXbA4YgvwDAz8rpgXxInCgWv0jvHQB8wpkfqSNROTr9YyJ8quNG1r
6muycWiKZv6Sdkyzsr9647L5g2r6YbOT9JN4mkUBylhicWHhAJqwL6LuKiB1
fyMm2EAdr0d/zKl4mRUHCnj9ifGGmp2o+2q49Cg1Smq/1xOXbQuxlbwEod+Q
q6IIRnB2hs0Kp7eJsy/qUtS2CQw8vpsBSx2egexcLG4F0oG4LXQ6q+8FRbGF
dLZGoGmUI0RPbql02sSv6canQpTiUIjwrKlJAhX/4kItHoqN0+JsunTiIK1M
HvLubNAxcP+1c6Xil9RL7WnVycBBCQNq8yyB3vz94Db3cJyHEqOpyvf89pe6
01FO0NtV9PbxsvvtA/g0WrvLfCpsYTGl71SI3sEj2512SyUZdaez4lYiDkA0
oTTe/8sBoPFmP5juOvPIuzK5V4cEgwXAVre2V3nzb1SsgNNVM1KyZBsqOmnH
wzOhlb1dYy4qAwdDPUD/LCrppHoYZ7xNGzUyCuPHOqYalMOhItF/s9MxKrVE
+VPj7xPdu5nWssIykval8ochenLzb/CMmO0L9/WeTd3nkrUxQuSr6LeQKKIk
Q84B8QPOaYHh02tox0DWnuWFHSKfnVyG2/dhwEnzjfPBm/kWYtTh4OvgM0I5
0+A93+wB8q25V/OrawGmXOPBScqPV4izREygrZK4Fp17nlMh9GIl4A6Yuisb
wsLRnFtHZ2NiodtIFIKLPRaYur1vFHZgWZhsyNVQQJnnInK7UECUdKHH2UFF
Slj+MNC3NkIa6P/CjxlFR3mEz353yXPOSKM3R4nsu6VCDAPg/NXURH7670Iq
jQI/UA0+5haXPxd1UVImlvrGMPqQbuXilJhHtVjyWAwJuBwVUYAQGJcFJp82
OWAZn/TjLswVvnHFBWvXig/CuMYat69REhE+msmNUY6Fu+XmBWCxrTQ01Yrn
hECqM3VNWp7/EqZfC7yCTllJ7CixevOO650OdKnJBroOz/P5LFq+x/NtFJ56
6ekQaxJE0lFtddZRkp6Ie0jR2D0/ZCQyPeWD+1KtU6gRAFhW/8tCQxHrP9H2
JtFgbWMJvKvG4P43DSs5aMxk/0ZiyC7ITBKbGbfNRkKrJapxEYcwh99lQ4gn
AJuX1umQeYqM1dtiAqkCpXTycQqhb+19LE51cMwuLOFBlseE5hmXiCFMWZV0
zioqkGKk5hErPhubDjwyqBIK4insMbkA8gTmsqYvKRJVJ91Zr1CDAI5GRJsx
vwuEWGnFfnNPa6ygguAhNCae70tgujO70A5cEmFfCQKvJwQIcMkA7vx0sobS
b61FLTwNhfnU1n3KZ1PfMhMQYQtho7MpqLtngYZq2ojkonV529ODPHZlLqt4
pu/0QJw4O4yCzCgyECdrG004R6bXcIVGPjv1YxLLpONt6KNdkKoYbXM2On0A
L67vY0RgEkEi8h17o7GYqSIjNhOZBZNyeGjjZ+UG0EYHE9Qtaa/+wfuf4kl7
zSos13Djw0e2JywiDkddItS0J/PThyi5j0Q/tW9MQXgPvzFQvJqKdyW+pXir
SyBfgjJT11Qgu3+FA58s5e7tTMkK1lsghCXIIPCRKld0d1wbHUR37LxGgGY0
tiGdzJx64A7uxo7ZreEzzi3ATmuLuB5z0EF4JewvTM9InotHfwUjKwlTVfhH
/Uvx0N1yIuWm6gHlvscRJbK2dyaT17ZVlAoW51HQ0WU5QtKMy8/tdtYDoCID
AjYMy0tqbV8mcm8mtAFvykLQL4ror52Xj5wcLY+TQrBSwfXmqoTtYloOCTJm
czwTJWpi3cbrz6vjaJVKvmMEI+7HMGfAT+N+n71esHiKOPUX4XwEmV+HKd7M
khk9iywMteZH6RdnVRz3y5RI+Jl9C9IStiaSUjYDvroDyma+cTNpKQLQnYD2
x8UACTTiOwHVnlVsrfyXfCQKqfyXosX1clT8kCHkqs034uT3w5c+Utq1wHw2
/cbIPb+OwfxvLj1VHwp/YQ7Fgcls8s6BB1j+Vf4q69S5oFZh8BrSiXgp1Aj/
e/hTolyqY04VJ69cK37g5gN/I6BdMg8O0IBKjaSCIhZsQq/OXnvmy3XbsDyM
aoZTyHeMhQT/Hdq/U+WjoPSgX/gcdnw5zVksVUYEAS6ZvgxO8uFzQe+/+4hG
hzaqnPyrOSl9uREeL7h8+8edOvyzXjcIzIk9F1o2wpEVV7SnyIEZuKRSBm9H
EddwSmLrT2TUlp3mNtbiGvzus//eV09/Ve8hkhWZ51jvSSO5cqnsGU2qDaG5
eaMDq9MzvptsbmAqULChuzVuXlALpr2gmh4P7eOpyCIppk9vHAd7nXqbRex5
qbZxVG9EmvPMj/BhaDMmw41VnBIu+qqURm4qDTEkX4dyOYrXZBfgYs7VhBLW
ldG839q3/yl1H9dpifPG3D3JSWFTS7ma3Of3HLmcsLv36/4C3ITfaxkRbg4e
X5tIq2ubaznvg9dIKUnFRHWEUgZIduVsct68Sk5biASrptathmlYQ/HNhl60
N2okUk8N8kK3xsvobB3Qcjj7+nTih0Kpa1+f2g/uarF6g9psZrtW4VlXEer/
s8p7Aeilaodk1I2DTFlOkgAoTlKIbmYogJz2CbzpM05LDQIqXnuHhKIANLtP
SrgyvNEn05BjKIQAWwN4+P5dvqvi/YEYc9noQM5cUs4hpt43D20UKcv9/BE9
YElFT3LXt8C7Nyu/07vpe6jkLJiA9dFiHAGR8f6p4E0P/PdVrJEPySaYxsuG
sXN7ui/TOC2mybsj0INUaA+yypPpuOu8GasM5UnvjTcSUK0zkXvsPbOhNhdu
Vx1QzaYfmjxpBHn5fqnDFuT8VCOhKL4jn+6O+UGTrmMJ1R9W6fj+9VIiJEhQ
hGtWndZ+tff/9SiSCYYmCHy571rf8TCMZ8SN6eT2L+liMd39LGMvRl+KR72V
XnFgFl6ZPH5YNz8w/8QtxEDuMOOCBnvm5QLU8o6V+DfzxbjlkD2LA6S0QHGC
EPg0SnkuwvUioqnd3TigW73QDffhH+NK7GFzsxMZi9FX2p9hA5mAZ2iYYSyd
D10oae4RfHwpROf7Kf9uJ+3aCPRwi8AdqGMXd/jUoC3m2u2NYiKaIQtd8010
3LrFAjeidM0dIOMK5DYjtIYxVvxnbqz2CmLWnc7sN3hhbxdcIf6Hhu9dacNx
AuPssg5Awf/SU5mFFikIzScjEjM2GD0ECVE6ZkgZanIXzfHVKscHvn97FnGq
KF1KgYd+/KJiBGWrdsm7h77hkkr+DLv43O++ISab9iVq/yFIW8esVwwarbvN
gksdrrjmoHlKM4gslJTY7rOkMlLOcfhj8MA0TIUEuxT3g/J6oBLSTgfRXrO5
9gh2xT5krt+GGM+Y2LMiI5llOsB3p2d9Unfd3HH2GplkkAPLTWkBNyO9WYCI
dfA+drkdSyTMLfTpU9gncx3IwoQoIZNmhsfBSJRNGsoPt0xK/QhBuU6soDRl
1qnpZ54xaby3IXGgFUfZyD+alNdGfWSUhsfB7AyWCl4/qNDCDk9tPHhWU++K
Y1niQ2Ui3z2DpMSBIIaA7c9oB91gy/1hya8BQIQS9Z23t31V4/XPycxhulnn
jEDrDZ6dljiefhyWd/9E/hLEMXoYZpHIvSDgrDOZC/IcI3uwymAmllm5Gzqx
7vrkEns6FTaZt2OFuKgWL3rQy0wYP+4X/8mENdNiPu9HelzEHgag5tav9R5r
cq+fQDjTxG81+rht6ZOmPfatoG/8TmCLFhQYsBpXKCKgNjzsQSfKl8BVJShQ
3bJjxS9TDXpAv+PpwtI7cyAr5drGSRO+Wb+U1g6iE2delokWJ/X4AeesE30C
a71u6m90rJNMiuDPuZQKifpgBEkuvWke3GDspAjI/NrOkFEZ3VnbL4LCOhKp
wLITjK19Cf3hbsrWuib7h6vkIcnoXZrsYecVEYxSGFtFR+pwfaRpuRmdnDAn
ppW9oMfvgQHZ2n9CuGmT65QT9vp8AmxS71j6+Z0jYEQ8FJSXrJ8VfWxXn6Sg
9Cc6EGzs0DrQcNiGvvGXQZukGJhVOu39PeKpVBm/gGwGeTc/wK9jFfbjzHgl
56MefPdVoiJFRHfPdOIgZKwCTG3SQNGgOzUkHg1iZuN2WoEDpbImVpfUCu+J
fk4UDkYRDxtoGP96mdS4+80UPTMG9jLz9sLrHEc2rb+WqPj2NBE/15QL2jv9
BD/wT5HUudA9wCM/WvD7txD4S2hbCuIflddgCZS+t65b84RfxVV+5/e7X5UD
8/WaZ+E30S1SerAamSvtyEtog3ydAMPBPCDIl5ELMPDcgXj1ZaO28Oy9XDNL
cclRjKgZjYLrLqhNNpLZfGKJ1ac/e9/iA+bUZezDWst4PwLp3kNBHKRNnfdV
5MfAHxHFjv2MZGB7OuI0n1CVHYxXPmPFKe9rE0vfqwVAyCKcsL+tQvdZz4Rd
KYokTrn2QLo6066nNwpVJRCuETR1V+0IvG1SCzTUO7Tom2rLE4mnAM2ld81i
uVhU+RFD65zeEU4+e2nUMph3MiUJedX5gvyqVYU7VPv73QmmenuoaD6Mn+qQ
+db7tLTY1KWvCKHAiHL+myiW9CTZV49WvJLIVS+trAUARY6xOK94P3nySUjb
Ic4EpVslKmYftOQtCcBkFMPv8Rs6bTi82rJe4PZZuMAAWMdt1BP1KKNFFYxl
E8Vmc6jl8SIduiBz7GjS4lhQwRoviuCDMCRGJ2pcq6jwkqen3T5IBFlAeAlV
3zbIE1LdPKhEjEh2jI3FYC3Ti5FobzIRZCe/xBUC1nK80oNxONl2BZFMyYSC
kFhkf4JDFO7LO7Mc8GFCfuzCSxXxXxCWav7mPEyST+RuGizNvfdHwyFxTMZB
0nO0BqnpoOMgMxx4TZqgE/XDAYxD/sEpVLL4+tUC8nPrdRjsDSUvVPaOqwHU
lbZ4Vx3AB9d8TdazbKqhQTDUQwHhDeKBRM1gt6fTPZPavEUpb1Qs6JFMtYmC
9PaueSiCUgQdTdVh5D+WCvQaLLELVnie19pLoH+HS67eb8IlcyLuAc15N1TH
Kei4lPFt/i3sARViMWCkEi9VGV4UBOnJu9zqodqncwMz/Nsm4A2sOaw6RVW2
4Bn8YHRofYIWbmFwxQBdPCYuA4xxrYtuq5SmrnHh98VHYIIidfncpvV6sRs+
j3V0zLKjcMdm4/4ZMxwFll939jnhaWj7+9xpFcVUK8aDd8sn4r9C+226j4Wa
pxMZnSmij9WDbekO2IkE9SKrRmETWg8DwrOChW7JHaGt+NCLHsG8OtFNwYcy
HBn0G/9OT+YFEghgf/C8MmcQzKaS5zKkCBBAW5YBoBE797PXDkfoBOsClUKa
piEWpWChqneZygC4zcFv/YPmr/u+7M+OY45tiXaClIwUnho4AoHxEO9YWl/n
GnxP+GKKQvAUo2IMoef1J82vfmevNLHj5zU8yrA0P9sVF0lHIapeqEdPrUo4
oWdeumjKdreBRBv0Ose2CSrUjFhIOd1gb8lohHc+HaV3f4U7LC0xZZMKtLZB
ZUhIpgpenobdR51aENNv2PREGaOUsd6vXAjW28IdiMfAMGWsRCpCPzVidvUR
4rLe7xI6UCk9MYuvgQYNHK4qA8KKcl0MkiJ+OsVWJJchnMn8hjwh2/MOiAXR
cTMkAXQ/Kqf2lXNCU/nI0nzs2BG2fFfufciocJirNP3XQKLBc/IuijcwS9WG
Nx97wFNYZtaR/soJSIHY/tBbBIRSfrNB2dJy8l2Q6y0dYAmqW8qhqnKmJlpe
qw/uk1EszYROdk1EqC45eqJo7/cLdtrpd/oB87lmpT+Y/EUclwABiwtJ7P+P
10vntTLvOv+607qQNxH57s9X+p2nXPvsMrz00VyWDp8GqOP0VLInj/APthn2
9ah8bBbrGT8CxsT+29GOMalpdoamnU5k3yRbkwGqnc3ek+u6pDlQWt09tZhk
zi0ly0ASvNa+vJj+rZWLJNiZEh2cIyy2h1BrDgG7gsUcCv5TNxvZnSGfz/tz
orPWsRrsFj9CkzZgTXRctnizeJKfoWdjNY8zjhSPjiv/jWjBGGRosCR2hPh3
c9oauwupTOdb5bA6HMi7Xry8f7MkgYcx4ikQwXgI7WakWUpCNnKMxqIVRtm2
ap5O2Fvsxbc26GXvsjiAAkEl5mJ+gBDaNunyivaoI1KGG3I5Py60WccHSJYP
UtUhsLqNLecKZObs0LIpJOsk14aSHNV8xGw9kLKNqzCpwqGIsOXJQzA7cK3n
+4NdsslvyHQlG9UeX8gilo35C2kXtH6gXdbVL9Q7HXHp+G0pNOQ+Fy6FAzrt
fdOcPhaISmBHdNJy8oeN20GysaNZ/EC9UHPOV8UEn1AoWOJL4ZEsy2dMkSGS
ZndbDskBQCWnFkKqc4M6VQ0T0kqoJFHfyyCaRIbexLs0scv/j4t1IaXnmrva
Cg1yiBhkDagedd8h5wv+8lsuE5JVlIQVsdFQwNERk7kKh4Iw+ZvJIzBRHrZX
SSOQwzObXtWkfKk7sxRn5OAa47yZB2G34XgpuNI+zA8U8TLKT9HMevMVkUq8
Zm4fkHVBW9NYP2voXo3DP4lgo2iqJS8189bzDbIWOgLyMYran/FYjjfTZRQN
0QPVp3nwRvS1XDE7Nq0/rwwOaAKP/lCrnNoElE8EfKRwAMnrSRO9Nl32zqc4
4LDrtCLi1Ml65trZ5w0ym+OVHdvz0Q8cS/2Wl0yfppniyEYxkk1jf68+zN1y
3oRjp2xR6VuSzN+kI8OsTTjjnzuldrOKrqEMPijqKb7qSbS57qrkw8THNR2I
uQaI3p07vre3lzVH1zFZrnf5X7pjq/ZA69xlkhIs4xrtwjwYM79VebjnfQWO
sF04ylKp79B3XP2/P1Z4ifO1KtddKpA38nfvS7Fkq2MTdUIg+5eKKVLuyo9Q
K5lf5fJeF4eQG+o3nfrP3Esg19ZuXFIv+P7B2l2z11JVp+B6Dgr6ycAqmT61
MBBoA8ExVdTkE9LjXzMdByt+J4Byt+48uwQoR0doZru7gk0OM2e62iOglrnU
NZXEdHCDSzrwJH/4328+bMs/lTg2eAOcRj58yt/k/kdFGKe+x9oKNw9Jj/QX
6Jep9ol3D8l9dnJzF7VZzh3j1EUUAY/Dgz2Il4Zt9fK5RXbuqBpn33Kuj1ac
Cbn0te6KiFeiBudmOtFg88XPmvmRBd105ABwIZ3nngTsUNohgL4WrUnwTBv9
awgJhbAGp7WOSuWV6+KpIZxexC1Z5/m1FHhJcudKKeMiMm2N+qf3U0Uuax/D
6bZPbYYkDztW3pKBn3ctsQtnuunseFtFG9kuU5ABpTuXdBEPKq4Xq93YDTF5
DGPK1hI09tmEpWN/340tTk1h5MwBYDr3F4YE0sDJglgmduHo8vb/+luKt9bp
lRdOtMsinGSn255J0qxrmN6BeTMLrUupgUvqMmZT4zNaO02iGxeEk5uQ6ebG
dVO6dIijJy/iRtPRBrEgUnQYpmaAd2kFIK+PogZyhI+RHZoaJsPEyX926Nez
zni1AKB4cMjmUJAUA5nrQX62FwCetL/YLJ28sxGocRIK7ALKga4YrZ4bYjr7
YDwlkIROkrbZdBomdRnZ38hlpdfvgYLzdNVLEjBasrW+PWAZuPE7/2rT+M1u
sJ0yEiC/HXFE6GVL+n8f2IZfC0vjex6QakHnkQnaYXRmlA3kAhzcZeiQJI0l
PB950Nhch9bZFtvfrHQPa51XkwiQGGcfHKl/L9xHX5SzP2KqsbLk5YH8u/o5
7eB9iW7BiE09KnY4H+RJqTfZuLQNSSk2OGgebWxHqnYAzeUJXUXO8ZthR/JO
gtH4OE46qrjt0nfz/vVN5ltARLA+oCun6MBltyFLyXx88mZTfvOawhlfYnjI
dc3JoB1knuEQVQJTN2qVMrR7/udzMjlJoVkGg5D24LYMFMvNs/71ODzpAimF
cnWTDHCUSZeEnM7MGXjYiGR1yOSxDdlUqEegcHZ0wwJeo5xFBcemdfCVJ94m
d2XN8tAVoRj356QIujn7xt8AdkyirHAeI7RIZV9SBTVM5iHyPqqQcU9apxsb
nFwyPeGKMXg+o+zGFkTAl97I/H75D4e/tPjchIG3cYb8ydEPTgK9v7ZfYR5n
dVLIIb9rhS3SwpJL5gC8FOF5johuZI9xFjf5XYh/Wn25nIhK+IkQXw7QZhHI
6xL4BhdIIukdP1LAsVq1D8iC9vq/Eozds6k1xyGXmUJWmrUrvJrKGAq8wxvB
XnJIIcdSNSxhgIb/Enmm+S0tLywlRO9bHx0QpaxIi9IJKwMpDCTtXGtfxAr6
U8waeLDCZ9Kgq94nVUSCYYinHCYb0VWMepGAlbu8yZDTyBl40f6OC3izqixd
nFGZN0zLGuqWEo6b5UFJQYDS0TbYkQgKw5jFoWM2LPMVVbN1IebOpj+udO3L
YyG0vZaWkb6CSMp7Zo32ZzD2cmcTdpMu0sysPgSR+0n0xIWkBPm3SGi06cg9
hYRrpM2hkZV+D3Zn5+RlY4wGyebId3X/Aeo2CO9Hx/EAj6dSqV7+FvKcpc9d
07lCJnovIY4UqcmPiKFBfZfkmD+zdQv6M+6RL+L9rmZQI/FeE/E6tJ9JHwgW
fmGOFNGZkIYJ4hZpLwe9Sywbq2OZNH7uGKtelfX6RZnjP5STExe4KAFlMVRY
tMuOw/Fnva6bVByQO/1YpXdUNHjyzwCVEgdNiHCY+6Tc0I4Tp6cfZDPyZcMN
bZz4IMCFuA1YRrRv4AygDY6Sb0UAwC9DzwiFh/jXV6mnrEIT+FCScgUnu52p
YghYcoRI3v+mFjyjpN1Qvbx2yoDfg1zI+RbBEFsDYaKIP3MUTSYYGMspG2ll
dKFXnGO2U+g5Lbu1Q7CfXORjenD9XBZ849w6EoHhAAhq6UQgAZkzcods8rmb
LzMndCW0MWdsc0RtxyZEyaTegCKaPMOXtJvX0jhVFXM7A0xNlRNUksyGi5WD
AKD0ej9vdLVUyBKHioH4cnjK9CjXd3gGEWTtBuwrPJumqdIKe+UCPrq9MaAQ
SCHcKi9xGmQKkbkKJk/OV2NtcOFz9er6YsjYnDv02RLYyJrPewnMtL1AikYR
CyueGBjcgWtV4VLb5he0v5IJQWbQ9PRFUQKi69ew0MZDad88PcTPbvITlEfM
x6Qf+2Rz+YOMrbYqcfOYc7FOce6FfZMYJ4cduUsmI+ryeyEy6HkCI0J5J7tr
qIUM/OrATZPE5naWKLPBjCDVAZa2MRwBLzIawGzpcPz1+uWxWskCdZtQOtVT
hxrl7TGh4CqEGNpmgQCK1usR5Il6al/SUb7sd263gQUyQ7uZyqyAyM6z9Yjb
AUVFcyC4nqnHw4JHFpd/xIJNJtj3SH2rKZ7faE0jLZgsiZ9lzzYk6QyrS3AI
spbmHA3C8lIrYXXeVxPTf8mxB+1TqSLw9EvOJYx5Tn+kcOm/zg/BJJfrA5A0
+NfSeQ7/QppKYDPLYy7O7jlLY0QwkTp578V7fC/an3qwomsI2DLl5ch8F3ZE
1gMtjA0Pn2FqkWKzNb6vbO3Sep0HRcoFVEsnIfyodV0Bj9Rlm0vLrC8lQ+5V
spBeeYMp+3VXdUeqvCkUb8JsatpUdWknadUDj8DlyMIXj/j8TumyIrfVUbev
XBbTLbpnScEthJSCzRyR+gHIizIBvbbKAxMepxOgwBMJ3I0X5gwXaj/7TaG/
mqWNp/2dzXQrDAMcVM8KVABdfsyI1PZgdpEXZTDrkkD0K/Up3+p7mFSpw3OJ
O9zNjDAt8H/vnnDwrAoz0GVjXaDuPNSLTG8421ac6XnIOmF0qYRzx7zLUeXx
58OR0qwf/fsth5Ys7ZogomkUn4p/gP9Ds99jbdWV48rYxvdLuQGWk6JwOGDv
TecR3+obEiIUVzV6sC1PCoCSUYbOFlqDA6YkMKiP0Ur0thx03pJpHdfkw6om
su0jLy95n8aFI95dPRE434AGQDLZG933YNezoLY5vogC1mSkxKfyRfmJmKcu
3IoZFBjJgxksndllENIGvFT2ySjsxXcxpKMi/ikB5Vor0pawfOh/Yh4FgaE7
Ca/nedvlCUAMehM70A/XsaQL1NSr/vkr32/RsfqRQ6Mhcm6lGsJy/0P7adWB
klHkeRS+0YiG2/8EBmtIOIzWRiXqRkO71SaIRuPSfo5AhQZ+VyJomkwdl1yg
hFT7Ddg4zyJJumWRGKTrnC1Cz+oQ6mWe1zQvZscJvmEXl5lo/2tvWIPtsMan
7IS9vIyfauNdPNRuOL2tonTfkedW+wxel5cRvck/VOOQnnow8s3S4tIl4nxT
OVdIAK4nOLCN0ftjpACyneSpmqusDdkRgO4zLbEEa6zML7CeB0L8rRN4InXi
naq27hctB08Dk90rmqCluYtewxzuLIuGSiS7OBkk3u1VUaWIhzQnUSZroE4/
tS2xaaFMQCmD1pts1Gq5b0JD1MhX1k0aKckRTIdHGDR9u2f8dC1jdZqdA1IY
Xx7aabsfm2WRYWhf+RcutH/xCCWzY4dG6IYOfXbLJUGEjmovYxZtewzLyjFf
sSQiXdNkTKHzCuLpNNcbFfWaKgA/9rbq4LTqj1ZfxWxUco+ppLBkqh8OuEkn
Zf/sphFIAxGP6O8lugmtsUb9gNJHvEUGBTnP7ArtRNdYl5JPaBWSQ5m2ae3B
ZSJQ27BNPDZfHNpS65I4DDxE/VcTCI2+teyord0a7ZJS4uKzebQl3v+7IA6N
jJptxeXNoCVTNaTT6K6ppXcL4jInLwmUg0sb6igYXBGMZ0nUMNR9EFXE+K1v
aOhqtZH7PiqIOaka7c7uR+h29XoM5dSo6i+NGLT4hT81X+oCuiz/arDBmR33
bHhQiWBohd1t2rMTSpdfVEUyWJhkjnnnadzqevdw6NtgpkOqTYQbZdtVbHiq
S54S25GIokr/jglZs6tSjcoIVE1rHRCfxtbR+k6iLyrZaS8D4jTngPPSGLb+
6B/mWKoJ4jTni6yElQdQx3j+SpLKg2b4mgpeY2KQvGt2aPjYYHlihcDVAzSq
CzffH4suEBpgPaneJ54Wuz1cVrzqVe8hlTOMD5bjXcNErV3xeRVhTX5HxyV6
ZwGN6qryup5lVCfBQpFh5e2zxRfeLaeArBpyB4u+iKnXbUAnsKwA0qLlWEzy
wQpL5aH1AWDeMxDj0rhz7pNC5iif+70uHrEplMTbdF7RrOfRg6j/Pq04vX+t
BHdc3jIGmd1r63zA7qtwfbe7s/Y3d5B4loXhSKDnS/8s0l/DWu7a4y3opjJN
MzLDPNB5AXygvIo6mXrqqo73pK/niR9swEU7iMVmco2ArgpKCw/zuxfIpFd9
bol3i+2Susqt3sHVqx5+2htdOQXVTUM/0don4iiGoTsWE8EE2KBrkhpXUAxJ
g4smQ3MFrQdAzxM5FQdmCmYZvGWKX7FYwWDUl6CzwgTBBPaznLS8/5TlKlM9
pRSz05LFzFog32ojBC+KpPpgtiUJ+RSLbMI6s1wviXzIGtVNAsFdYJanPEV7
I3wldMODc7nrbnzQS1mQ4JRoWi0Uhv7wrAkeELOEWaTygBk6Ki5CQysI8np0
sIGFTYSE1MeLoxc/6TuxR6MgbWVayyaD6GflDueZypTW7U6ZEHSVHF4XReBc
GtzpLedRS6KJKW6sHX+esLeV9JM5d5pFErGiIeUq8uAuGoH82zRk55a/aD19
cs2UTxLX7LhaOfkwR5xWU4RuwFj57xoZ9imLr+rESc86vV/DdTBEekd0Zwul
8pnlYkt/TAFU0K2mTI79SzNZ4rL1G8nlvreDiMmOm3+n3/E/rZsxQSGbsk06
8ntxHRV9HPl7jgYE//4llYfD/Y55d5Y3l34v50uG4yMFh/J2lMhRwtw0fe4s
HZX2+WdV9zMJRdcVhpCeisfMitkKyTDBMzEJBMbtp1Th/TT3zDsrAfssmFIw
36dbjKclx8CpT63XW483YlQc2URUrse25z4DRhnQA6Z5ldJg90CbnEYIhALE
Vbv8MCr3ACX7U80wEhMhwSs7PTAmrRZkRcLwaJLditRT76bxVMpCtn+nkiG4
JOIZsagoUrAoz7F79ahb5A6QSo5aKjp7f+9cNIFZmjkvUoluzAIZddodonvH
tEqG7tGvJHylRL2t4szCth0RSas/blWNNF+A3cpHW0/U2t6adl4htF5Mpguv
yRCKNSElbbdtGJCvEJ4Gm7mdhlhODvUsebDPpwTt7Pho/dNcPuO5nac6mERQ
akYpv2jS2NfaOj8JKs++o0pgkIjSD6Z/9irDOor0wZsEaLtYtFtybpNIDREZ
XnLU3H2Jas5VubeF6iQ/SVO0Cs++x17d3hkjHSM55C0fyjOz744UZJiik8Gn
pw/QMdHJ84SGrLbBYdXUyrB813I3sKELi3wcqevWs+m4lOm/UyTEjHwe9XUA
3j1flEVZfG4pa9MPibaID1vNV2/pKWyX+XgVCYuwW53nXgU2I+upR7Hgl6cB
FCd21EEAQwrKERPxEe9UbTn/4l7Ot/DyyKbTuf2RIa2R0zk5/LlgX2hzRt1B
mH2CY69Y1qq8cRUd5dQ5RGMAIxtQLiTWeu54I8pam8sNC+kH6GhMby/WVwej
h2Cbh2g+gMLqerooTe/V9b4cgxx7ypWACu5WHF2+mp24W1DhPgPgsSu0RoAy
xQ90EprhIstmdjMGGxJT32qr+KHCfrSv1M8crSHqmIvBYf7KlF/Kkh24863B
L0AxWSZz0GCI71pVmGSdAIG6RQT7YorewwJHsonVMeISYS3cUfamtYIOBDJ9
qUeFOmmrJvKbkfHtlcnHSpjqKayxz24MGsv4wOYhV4GOfY3ejs03ViituPOM
lGrQJlvseSri3yu2pCSpyHXe/pbAWIFD8l9TkoBjXqmkD9M6T+uySoGRJe74
zctaMCWZCSIQsFqIeiLo74eAJ3uHFEKEbKEo2ak0BhbL2mNPF2E+I8mFKwx4
+eROfxWFFe/a/X18xx/EbyFC2ZagW4p3rz2jzzpWEqhpwb9iZpfbZp6UL6bE
4qop/FR2uGgRG8fIQ3FFxiLahHu04/ZdGuo5JxTKz0bnsG2bZ6GOAnOER7Mg
N91itJHIWNMLCKLzzFXr4PzvzqbFly6/QBsja0dvwsf4y9FR5BcVT4qmXhlQ
/XdqCkHM27s2NDjMZBmvGAxiYDrzapcQsSKEbEEQinKlrpy7Jo6pJmaHeSay
ULmHf6KZsCTYofXqgUaXjn9yen/XR3el59tRAsYbcFROUrQHSKqt+WTc6sLz
MvtaL806nXFXRwuUr1BJpo6B9QGxzX1C3Eejk/l3/DUyDYoc29NYr1GP+eLh
rvP+zJojVJwHXQz9ZkQSfN184HPUZgZw/sP2htvCnyZtQ7h7IWLobqAjpacM
6B8lw55CPeO/+A5ilQJWmP7hjat6BWaDSNNqU0YgPjacu/wOXxHzTeBGFtnu
eBQqoF50+zgVOiNLVvTPlBW81s8hF9kaF+25xjZeEVh2b7J81Jf3CR4MpHs2
ONjCMGhUeWfyRXxwIrafDKTRetHfXAHnbNFWLWwfGx+TIxXfU9YqMC5dQ16Q
zOpIbzFPGc3U1G5GTdCSISYd6/Ek+lYX44vxEBTP+GC6C2MPfMOCgJ73fas7
1xqihodMi7InUgTN4j4UhLtwxshycVQ0eChd4RNrEaBaaGkibhQxzZ27Epto
blUNNKlD7pXsHTwZfellNL9ZvawTVJaV6PQXnzi/RR1bhxWsZhabt8AIRm6b
x9uEOlQUyQ22UDqLDsD9gAtCcjn2XBwhaqSh/z6vDlFCirjLKHRIxdtjyD6V
0OW2CP146OB6U6TyCZX1IFKTRsIZGymoODmfst6D2WQxeSnnIvbk7Z77D6cn
ZapEWZCOzH1/sKz8jCv7OP6Okh30HZXFOIKr6JJFlnW+eGC+7OnLz+d90lpf
y1oZ3+uVSYS3WYjcE3GhMoNgbaUGr0ENh2lztab4fNvVutnBb1UYecYZGKhZ
VY+TTnA9NpSKiSo3NuuNjLu95t0B/x7T4x10O1f2zzAZRDFrQR6CBj3n1M3Z
3HSGSmGceJgLSZzm4/xsyEgNGgQcy9dcoW58TcqUeOSMv2px6+pJYhBiXek1
lKH1UH5GXRR6sY7rPQA/Jwq2ZXUooJMc2/TQE5k0RKl3I1HxzXoXbrK34RPK
wmhPBP7+P812AmRClgXQ1bVy0wI63Ib1Z45n3cgnSiWAp+eYIWFC35VqSaYG
MEdaRixOSTI+crMGC/1jFG3n22kGiHyRY7yS61DFpFvVZqhicLqh0MJaHu1e
qBCvdr4U4iwvDLijPO2vpRJhPoPZiWV+T4CnFxq0Qr8TZ8zyCi8WqBbexu8Y
GVJlMylFgZV6FXYy5bJgm0hSArGpp71CX1rjIcDVuoPr1sAaNSTV8LCLlZ1D
CeQDAUi2h31PzctjwY6Z+dlRQczTiF9Fsyi70GrFMz0RRSswypgc0A5uWqbm
5ejXmfYarhapD0JVqNckaDINh2F+zqLR5Nv2VsDRBsgfu3TFDxN0rbrKs0+y
7F9xMatCmENFWHWm2hqsqNMPXsiRWqEmtpzLM62Et/MKpKpLtsfzGcTqrAug
Tr6jIje/dr9Eg0M8pqbyqd2JhhIHkwgCcztKXe2n9dV5jXAfQ3jzX2CXAF2C
OoHnQYMJdxPDJiT7ycn+EqT59EVQdkX1556bePXtLUXet4xlMy127k9KwSsD
qS3hoHO1CTXMxqhgqalImtmvus0adXamvf0nEWcYmqSgEfnerC8YyQr3z+0T
v24WU+UBV1X0QrQrWyY+Ymrmi+HKeGTR5XSsLi/EvuW5Sdp2R6ViVnxpjb20
QeT0IcMAjn7W2kqDP8tACCkqkg40WnmJW6c5pKh19hJ7QAu7VlMgRugIMdIQ
28tfTQE6BwrZV36AsIOuEq6T3oP5RvznlXMIruhKp2zH5zzvwuDuYAlkNV+1
zUJ7DCoHV4ay/obgVCfYjeD0MP/C2P2kHsSfRowllOZV82A/gvP/ronVY16T
IT8jHiVSidl0dsQcZc3XaETmVgUBHVIbK1v9ubggzV0BpWdrg/FV5cu/8Uco
1f7drGQUy+UOdAQ3NPcziOWSrGhNmb7kNABANmU6qnXyCui/ab+fPBcgbKn5
R7yljIqEjTW1Czly6KQeVG15WbRbRFfiCcxzW2Wa6V+R9kNapoW2O3AQUpZY
yb9qLJM/2SbIl89JNOMXmLwAsJDITknKmAfabV+bCsaAv5RPblqM6bwoHCXp
oZ4axAUimcmqFzQoImGheA2yWTjIP93dPD90o0ndnwXAYm03e889DjQx/Q3G
jiBDJ59oJlUFW0iwaTWekpTEj/57E+NdUV3msrANqWGx6SNDJ+PEK7Jw1Ne5
hNwJPEN6P0QiIylgwBbyPn9kl9BE6QMAwV9Bj2TTkWtPMKTdx/z+N9Gf4/U3
AHVUDemtNF1RxQZNu4OugerpOBkx7bfmdNkW6sdULUYm2fnR04InaX9zLPhp
DBtNRw8GQE3kOvMZRkLTaJi7x/o127UOzPFntCQ3/C+LM0WYBS+bBsWFppWp
bmAcI4/9FpgvcxSZ/ocQf3ctHsIaXVSrs1j1FVxovr9HSNFioRVDGoleoSdU
ozo0UcKT1N3ZoFE0FrA/X7zn7NuB4PUrPfb+oyO6Nbf2ki70KBuheiZb9B7G
N7fAslXVuLj9uTCK8ycM9i6OQQiPnp7oYJxeIA9ygtbWVuw9UM8HeXig8Hoh
VS/3/zQfYt1kNwNs7kPaJu5qTIGTMh2UpjANWVdefx9z1Wu78Jh+n66hsWp9
l/vkNT+PSRF8fLrdXuKJsUsIW6jpjQu68QeR5rgzRZoszCXGS+iYVjAsNnYn
sxJrAnusJgeEmQardVFuAtqKXS88+y28Rp7WtYJAqsOpseXGks8uOLqtnLO0
RGvpVIrHrkikK3w8j5NTDs9RaGKulVoNvVWgOoR73UZl/NYUan/C1yjCAc3P
tCtVCWBnrZPXa7/mxq0juw8CKUBR0db+l5tJ9CbRsWt7De+qxj6VDYUgRTgQ
NfZ88z8bzkCK7ogAV2jN37g4hz2dQ8JZX0UmdG0CRv6X34A2ANcT4wpNNBEk
svYzNAMfa1yWpQ3YUdm4X+bQXlOdrQ/VzJHcWEl+BsMMRTXNrIuAzNHPOZqb
M2gisQavnAucPGjtF26qkDYhReTQsGmweiPe671d9wtaRBcmYN4wGapDZ8RX
edwJORj6TYHahhLEPdGwVEuTKbTIWRQyuSMmsDzc5Pgt8BAqMv4RlFGBPEVF
lX0L8HSFo6DmHMas5SeuSra/lYGVUpLIhsiMM7BAr8GbDNKYnLfUSgbzt+Vn
X8Lm5JHEnpdi4aGX/kDFGUE0kU4DWyKWlvIoKlsZ7kB9FaXeXzWXbexwy1ve
7/EO2rOhiPOgU9GDARUwWKaAqmHoLfbe6ihpwH0FlyEX/8hWY828hS/rkUGL
4XSUE0Rdf7RK8YvMW9ddEi8C+nlN74VKJUbOgzi1sm+J8MDncX5hMw5itQPq
wmtg9N0blDfjCwuTr/Z3qWSF37x5YO7nfum7j34FiVRQCI0YqcDCQfV+gevo
V6YNAU4TuA+kN1ziiI0u8DmxgSfs+Km/sjnC45yjvjIGkbq/zAHoHFgGFko+
d+8/nLe18rb3MQ72+ppBNFxs4/0zLDxsIxWQmV6P/xU9o3ysAdqaypcY/54F
FE/RPj7j8jKfq6kAI2pD+ogkAl1rl65guRqjFIeQ2+e/j8I+ESSJ3XEeuVbV
US3KBMiT4Pfwwy0NOHageuH28OfmkiridXo45LElwGWf/XHsyfgL+C5VgZlm
U5HsFzXWfcp1NCQZ3zgQ+LMMBxAs3TycN1PhBI9PTmJIsyBJTlKWC8fxzvfk
ukQrZTK49fbG5g7gEbH0DsbhOhR8wWbvD6KRI72oktEf2oO6qGXCsXDV9ndK
JGLEXdE7vBQyGZIiWZNWPrJbPMhIl5an0exrpNrCuQejF2UQ/iySBzRaYrYx
N/KzHfOKX8885ChGcGgBeOaBNwssQwdAtrkzytY1/eV5MFO3HPPHXYgcaG9t
4+LiShDkEz/B4xjGRyxTggd0aRHuMzbLLdbwPHAjtIkZidIKecPYnXMnO51O
W7LSmy64SbGnSWnaVKGCIZrOnSr8nG4UGzvt2tq6HuS+JbatY+0Zq1jUnUGw
eEwrxzvlw9mkX/WUaF1/jwVMCIUNz2mEdZlib06JVz76QOd9wex4k3uj5dtx
gXD/nwQWKOY5zPI6KITSuEd20KxY5CNs8dAlJyUW4o++WUHpYj0pTuU07Pzx
5VntwrE0eSev5n9s+3XSNkQR1xWKaK8LEy9gKOGBBeZDCN+cAv2rDeYgpe0M
Vx+JORMi4OEVv3GH61KllO1NYhWvpr3rj/4XrvXeZzShjCumS23hwhgVL/2N
DfcRrgoqSV6UBphIH+ICLDq8GgMaZDIG8pUWljVqIVuVfSwbjCHOqndmI+t8
s7JtcXnkeobP+JGyc4H0f8OA+87/swkGRkhPvVEnfdIIp7w89KZukMorESLZ
WTt6rlmTp+udW0wfGr1EAFNLqTI/hpSDxcx3aPiteyqp67/6XEEu/UssnhF7
V8eSXzTEp33YtPMT6R9uHVaJv7LmzhL2VUH2dcNoUuMIWk4F9UFgLVnT3wd7
j2xUJzpavbRM+bBXbta0GASboVqnMRI17ygXW+9F9GhmSblhD9wt9nBH+SrD
IJW00Mn1fBsm0WP7b/8015wBalhWGngEhROXi1Db8jWXDPSNMSk3q+CUkSCr
nN8ulJ6gDY3hPW9i06ODmP2J1sh+/zvJKvFTGDz2rgLC3aj7QYmqJFiotEff
k+eN1j2mGlkkOuGCieBTa6/6SfHd5WiV1x1qxus2UQqd3xZZno7Z40WeKsAM
DV2Kyo64cJsuunagrKmwkPkvMJFW4qM2JKECZAeYZ9Vy0JyRowy5q1QyncmX
a8WdDCfPVM0GOcUbTOP5xBVCfJNTmb1IWcjkJBghtFwuHxF5EEUl5knz+jwx
vV2FJ8qZpLnRQjsXJC6FxT87jD4/V/jwg4BcSt/ZwQzng2jcad+y73elFV83
6R68zexj2IMot1ugb0sjCjdj05t6VRG1aZCSsEtpBwCb9I5uaLEEUo+ktUx5
Y2OyOVAIqU9YmubxnKcC9/TIehKK94lFffiSfaunJy3CszOSk/zpaoyTspJW
/ZYTiBWcx72wYDXBJZyWVx6jWBbDGg5SUgm84yuJ+BvQcbxXRuNOrQBBY6XZ
T+laJxskigCg+XN8KJuPQAMYC2EJYPMRAveOMKiJL9zHEOXjjjsxmL6bmVM9
00OUugWOvUzgOY+lQXq3jxKmhiuAGCn1DOdG09gilkYHwL4oDCdeOA66JOhK
AjLD4dbBl7qJh55kW/+H16A2RMa0nuUqDhQJq+Spd6CDmqG0O7fx2KrBWr9O
JUq8VrvaE81oFZ4lb9SV3lZ+TzJoDShN9OLpR+8fyAQ/e+C5lTBr3SoLqE1I
w9X7n8Lj7IvvS43q2RhBvmKdUJ3bHH7i3a4SH/2roqNjZfWV+r/qc/tCV1Wh
l6sxkr23a4Gn2LZ83ZstoiQkXs8+5I/aMTbILWlDtWKCblC5kkGGC4fsyO9D
LIFm3KGsSqR58fX91cmgiY+MOz3hNc+jbT84USkR3mdK/z7Ib2N+4ypu8eTX
7iSpcqL2aeqblBkcRbcKK44qLjy2UZlqW/v3Gr+pLD6bfFeAc+q1hvQB1AKP
DnvfsyefAakQnN0+kDC8eoA+58FMjgikUMbPtYTB4E10bRtSHvaQ80+kiIzh
fFgYvJOK0qvj+07YNnQpgsuRpN2bxp+muxuSGuAF/+oAUX8s9f6D0V3GkaOo
lGvWGK3ElY3LZvLVqCGJc3ApX8ZfR3agad3uNguD8oY6dAdmN/pO5i8G1AsL
NikqHbLjTkMTYx+Bk4yIcmPwqw5Ckn28dAcbN5T5+wTVWWBwjRSkJZO8pmr+
GmO16PffTpHrOXNVTDmlSXSyAid+L67w+MZhiMiQGJHV3KA5y98/n1DpjriZ
z6JMIHt6D2MaqHh/L07J2j5fQQF+k6n67oKHKnrCIIuuEyZ6i7oILTTfXTNs
OXQ4tA6N+sGPLlZhPUTE92rHa+oWIAxjxjbLlGQRi0+vSAOnwd1QqKRxREir
2XQpdATxNriapAvXiKcA2z82kaRPRGTcITeVrIT5Kot8hJcff+G+V1hkDt1K
nGbfOwCoBnw5vB3YPgXFiYOaFze8m6cHdMmJ92GyA+ecgxqLPH7jbPqrA8SV
tZBK8m0bO+8aCkiQ8K3IBrHk4ol7G2k3NzDzkOOstCaymajDrUItFLpNwoI4
TRIC28exejccUzfR/e5KSB/+Maawjw8tuj1ELQxPBvyRoHIAzfBe7sQlt2QR
h4frolmtxhbAcv7tFbTJ8g++EegJZXCKlQnJ1OQZbqdm2E3Ov2ldgOuZhBv0
APRA5htDigXmaoalEM84O0oHt5bWhmWWFyhfBxlzdXL9aw9is/2wZWmpznzS
eVzKwG424S9gBmx6kOXruha2Nu1J5BvqXbMY4tXvEvP7mxnF5fpVvpPWY+l/
f/52lqMXH0edfYmW1BHrkd3R05isXJUmExovNpujlFfojT5ZBCsKdAjK76LD
J09ABRnXQ8jKQC8vx/0l8KkV31+uxatNc53ZXqsAfungzRCchHbMQyR7FS7u
ihqWZ7OzJpbNpoEEkS002DOdoyb8+4p5O+ybCrro5qjlld+6R+uOvdNqSJI6
M4/kk4o+WQpaSYTjaeGHHXZyHExDGK2uuag5cxEU8uY0D4HO5MAwrOqfuQOq
ihzH33GLX1LPXcO0CU86PCZO76rx6KXjb3E5cdbkZLpKDSctNyQNPmgVeOQP
xrG1xY8Xierq15yefeR//4sqjxeZeXTk2z8Vz2MfT8/hhjIyUz4ig/KjCxU8
AkgWlEuWEawai5tL7LttmubfPizHmsO2x7Wy5htVsIDqdXV99OzELnk6ycVq
SmY7MxmX2uMojDInh1nCA7q0RYSM2COsYF/lYVqB30aJH8jE2OPeTafHByOk
Ow4mrx8vXUar4Y2hITZbDaIC92AdvkHObeOagUxd9DrF4Vt+y3/jvpDPRQsg
fImS9/0fcY999ywTG2Po+qHJbW6p+jw7b1ASy+NKZpxul2DQUN4jCt8HMDjV
PI3R3KumrdJHgnIxFn2rASlYNcn/tLIzMxBtVEwI+sZgEjyuMxpOdDZu2a0b
QeBv0E5Gfo66TPukExjaJ9BptoL6H3V2XxLndyJKia5StGaIsvgjJg1wRfv8
ZjlOTyH0mvE8KZKuYB5TikaoJ/nl81xbJY54wgOnrVkx0yeOHSTZJ1vQATH0
S8eTi0L4xEhzeVXOSq0ngyNoSXgLyQGUd8EI4iS1lv5yLoZyCMaLvjceN4+q
eZeoHMmp9Y+FA0MOZv+G7UYRGzVbN8P/PSo/qj223mec3nWNyD14O7YBo48i
BPPrgM4WBhFw1HCFQqnwMjpFv4Y8OVKe3aoBkbidJaOcWu8KsxhP5weBViV9
zFz29Ddp21pdxkw2F289klxgwShC8Rp0bVejKQZU0iS54yVLF2lJGY9PHKOu
MrtAxsHuHzXU7+JXx2007DGbi6V2YB9h+SAZCPFSlhUgaiSovTe+QZ5p0dVx
T7AnXjjc+Ybr2utUPnODCysZdL5CzOPkNvEnnI7HVPPq/Qpws48qWLjZXAr5
EjPGZEEHFrmNNtxwgmStHa2xR0uBFR5tEiVYwqX/Rr8SQALm9aPGAQnKI9l8
jyQmebtlgFXj9QUza9d0nmsCTTqMyKoxdMYAxZ1l5gRODQt9j23RuP2QVAHX
d4a9fNu+e6NxOs/gue1IRoLHZVG/Wh0ajrli3CQ07ee3V9hyvZCz7DEz8CSe
xGQIDIr1npVHUoe2FG0GXyu1ztZuEEd9g8tBfXtaQ09mXuJGyWA1W7U5Jjd0
2im2bHFKzh6O6apVqQpDCmJKvaDbgJPsvv6aJURsDXPWglzxGoCpHiy1ic42
XLPLGPwen4sA7ShdwPcrej2XNRD7fpugIaQK2dOXmFzlLxbHAnbS/XdWF24Y
9qTzpt/Fd2P1A7tuJVytjqKsfnbrKfeSI5Z1BAha/s9sGZkySvQBVo4vOKmM
F9km0RC4jqGq2LN4OrCMZp9Dm4wvCoX0ypd+WeX9VCzPG0f6uF+FFkNzCa90
sn5TJ3MXXDBl/kdWAl7Oh9KFdxqRx00Nk8BX5GsR+Qmps8TozoCinzgBdWdo
iWAqyJwBZuwaschSI4Ln3M/aoT28Aaq+D0poeu6tckBEY3I9Mjl7OGLVj/FA
bOxl0br4nQae86j5LXkZZjmmCezCi7kNSUCp09MAYO5/VQskKFBgPoMOoHYw
XSkNDEPyykRv2eENdiIKh86B1CqciB4COCjcc0+fwZQl5nNAz9a2CCr+cZ71
UCJECdDijXx0slTWdTrumZIeQXOZzpSaMj6WoeEPuZJqSIAcBprYffT3N8qC
LoDp9DTy69wcWfpLw7DeVMp8Qyf/gXuHWZxtqlRkz3+UW7KZF/Duk42OjxtT
9FU7blGDOUBzbO2Fh3nRCvcWqRb7N01AU2iQHI4pfz6qweXveUsTON4S+Mqw
6mgiBXxMab+fBtyNY89yXQHE56Aj9ZdfiFICoAL3XmeYOpHpoOHSAOGCMvZM
ns38RrZJXVum2V2CQFipquG1jVkAFVSzW2pgkGdyVHLLk+FmqDBAs6qb3Qfx
+7KBytjbvi0R83wmFqG4pq5XDUsz7GnbXY/b2Omygg1DkIZUIr0XvTkBUI1T
v6rd8WN6GKEu8dL2+P+SkePZBElVB1QmDGTK2gyFPaNF9AXWEAzppK3vJZ2m
5oNNwfcXV2jztTs8i3FuyewZUkKF0ncnDJawKoIvFEAfh0rdLf/M4Rk2d0L/
vWAlkoX3x3cAByvPsD3ChI7eW1PeAQwFde8xGa60iMw9xsxJfLEMLtl7AJFp
D40f3hXg73pAq9SybrdH89UtBWBkqQTHtpKLc3S8i5CEqTxHuZbn2FrQTQB6
FJ4F2DZ7TcjWrmjSk1EenqFvNicHBOWhSbLggJATaXS5pavaNuKtzI+6qzJ+
PJd+99+LbSPqzAFAb/9lEibLTAC22fT1nMNjmDVIg7vX3WOKa8z1vsgL+NBo
6cQsUfcLsQajubRWssNGgpCR1KYTc13W70m/Kh2ltsF4l6FS4jDFUdxN1WSe
gMz4iLf3w9/yzMrH8tv6+jjH8ngGnV+DVbqwEXKuXYNmFAs6B5uLtBoeOMvE
vZgxeJJdWad3L5kuSeAZqVjUqRTqIfd3h14ASKuB/4E+uG1gHhDubdkXDwMJ
acS9GQbX2rCHHJNS+0i2Jhk4vpVoq/9HSp7Q8yhWTg+2JQglFqivwE5vENUP
FUJ0wYt/jRMwBFwh7bcNbCFFIVjriIga3fLz6OwJK0Un9Wz18aERn9k3j4ga
ozyj/i68mmzdbBu0/LHrhAgH31Noz+vSdPSMQZ5I5F7lHy/hq69o/lrtbbaO
dOkHAZYxn+BAg7xF4pHnyNJ+7E77lGkFa1rVSJKYu6DdqLIKq/XOtoe2ZezH
GnNiw41sNEi5PJmAwDz68dVz1PKrXXERZwcxGhlrMOOaODOP16DPmYYN9pJS
hUDG66ioFEV8kgKJTWPI8Pr+Hpso8xhsuc7Nvx5iaLRrdlTfAHDsfriaI95J
F5wKmtbm1ITZYtS1945iU4P80AcY7R8VfEHw21wTyrqj5RVjniw/vcB+Gzzu
tkcsAsjOK/JT7co7UY6TI4nNvKbNEAqn9lB4+fsB+MH2uUl5efPg4JcuxpA8
yOnbjZJ7Nl82/8Jl3ffPDIeSpqUlnVNKP1iMvRLf5NTSROx5BvbCiRBJplh+
mN6d/HdTcilbOb86Bh7nuVTZ6v2oYyCgt3eYeOI8M/obUbiLwMAQDfxSMNc8
L9VvybDfuuwC8NT5jaLuc005FCrizmII5Ul9gY63WUA+LQ9n+3nwJENZZwGL
9Md9TywfU6hcv6k90T5/31VTM71ozwDcgAfl4h2MSAnh6mNEQT8coodIfMUA
9efkfikP7i5KIxSO3ZeZ9focQheqlpFxere4F4OaApDJa7XPjdRfOj54dHuv
JrJD8i62eMGdADTk8XCeHDbDUPiOWxvvf2hVEmKfC67HuzqLoNYWWhdl3P8n
baDAP9/NuegazTA5iVhEA7ehaQbJhRvUUf7uDla6502YslCdZaxY2k97z200
MIevfQR0pR1X/nb/5D0F0avY2rNuyU9AmiLpyZroDY6smD6S+h5ihmUdLIyB
7/yZwyqwmls1eZC547XRBojV+DCrRRIuEQrYKRCjyqk7b66ROqsNqV7TQMAJ
Kn74WBoNrdHKNqvcPIsjiJ+ZO16gy8ssYmBF1iQExvYMDr14oW5PGZ1cuA60
nP+uf2+YKfLwMySmU6zKZv7oQ9FcP+6e4wtgK5U8SJZWD86dwkLKjNX3hyCh
rdH9y+rlo2UnX8h7a0oNL66QUiEvjrnyjHp33bLreHnq2/Jtvj946o5KWPkg
HkXBJwwePa5RXl3yhdsw5c1Slr+U+YlKhM/FRKnFr+z5JnDqiaPPiKBmeBA3
0M5ylvVDl4mSx94k+F6XA1STAPkJDEHPxBO+eSzlmgdXDIqrBEdCT+rYdG4j
9GMNxC5ml9Z0GKocjrd6LIdy+XUQflO6mK3KbeqpuZgFBFvp/XZZVBfa3EhH
/WFOiWrJynNr/+uB7IdMqsJzf4XnHIF25rZsQD6SavqGwaCHS6Z+OZj5x83o
7EU7kR7opUyNBsfqdbPUlpAxxJBhg6jHXyakTMmyLeUSMSDw3TRMV1gdt+SL
Hl7Xv1fxhrPNrYUhvGTslJQv+B5Z0wOAXSqIs40Xe6YYiltmBL1drSbtjrR3
8ilDivFTyeJ+UyMoTiJT6CezKDGImCOjuakqtO1B9uNrc4eg2BrVimME7UPT
KytyOJT/ReEtHReGb/zLUVgRYxeNTeTMpW7cTXqh4e38QR56XZGANil0tYdw
FBfDSCk8iOT5VHBKv9x7r7dfxdPPfp/iCYWb0bW2cegnJKIecg0cvQIGmaJ/
BPFPz/73KETfvxvbV4jdtgSGjlghDMfBnIVNyZzp09ojQBNktqwl8A45KKBj
7mv1y6sI5K2wHR8Ob4+1ZuEcu5Gwlx1fuJiiuqjfyyK4QbSokx/V5JUIGqK2
JblmL16m06nA9HcJTJA/O7p8HgffuM6Zh0QtcpVGxWK3E+7In1JTljA0rV0v
np5MchoMRpO2kJF6itI6S4Q0NcLohX7a3t1Da5ZLfGoZBqop4h8T9Vc2pCoo
OHkB8k2wyl2f0wyZZDX2dV48ZyL+k/qCp82I3OaUMaY5nMD2U56CMpRyK4j1
SbaEIlwwvhKCRHw5zjMDva4hwVY3I+aP5t/EpOsqj3fFjzwPTA1ciAVreLHs
figAbnMBGHd73rqMg6RLK+YhjlhxiVhEMN7DyOUT5tGJe5Rc+qNARPbH6q0C
v1XnHvytAwhixbAxXPsH9ksrd6koTi5S6mlX00bgoTalANyaYz7g/J34h0UZ
mV8K6EL9k+DU5LHxchwZlQlmsS/8BOCKQ23u981KltfNetiepvIhMrzpzOpS
vZypQNvI029y7BOXPD4/3uXzikCF/1rlGsqQh/IdmH0rNnE+yFljwZ09/ln0
YgMiNM6qhPsWhAVSGoikD1JMLdt7TRwrJlkeunfT2dklYi0mWoIexK9xSyS/
ff3zYURo5nQeaBJBh+FNgToomdZ4BIeloblJegbVX9xkMSb2Yr+DMjpkSmn6
D0g3LH3PBPMUmjwkPq4KBUXbYMs1PcPX6vJNZuWvLP8/Fe2AnG+xO2wnZRsn
UhreF1AoL7YB6N3E41phMYsEIq9AYGcppA5/+tQrcJF7kM1tpGidu+f7Fz3r
vRmUEiYooRmekGP1qHUR43KQ9m7gzzfoKxfs9dhRYLWb6f4SC1YYJlhzGTHi
UCGP9d1Mxmzk4n0NmFSl6moZlyW1HIrr/zZ6Cs6Y6gHeMwXfcwATkFE55ZAl
WW7JFjHzgiCbBoh7ETVQMuK5GHAzGUMjRWbyDiM8c1Kokzwr3kknTLbGL7m4
sjXw+kmfSQcUBzEgd91pAe1UvqqhITWuTiitJ3ig+gyalubyoMhjxNCycoJi
CekThvtl2NJcG8avIC2j3ssdaCNQSAwkRLbBY7NxX5o93GROtJX8UIkeCEd2
ATbAL6T0MEdOb+s/IXiD7zvkTU5krFFKFjbLjZ4ckHRaGiVe5AQoZEbz/+ox
STd+4RC7BkSIcsdz5RA9ZCQ1t3p5fy0DIaX4cDHaFt4XliC7CEPlUB28hOQl
wvqV8+7cexJSbRDeyZRYKbpC7U9Umnih/FNHtH8Y+raGzrN/X26mKU2I18NF
vnBMPzSQ/BB6ZXj15cpyWYnW/gZYuvITWDbp5ZDqRoYdec2vRCHvUHe9EUwg
WITk16/iXEOTMbls5VtWLLkWi1xw6cr7HoN9kWSanxnLhlhhyq3Kjg4yBsHt
nURRbg4VEy5FYfwEBMJsm0h01WUaO9unWtqGPJqVgUn9h+GokxwzFn0fqdmB
87HrBdvodi7Kn1UGuk0Iub2TNI4SNxHOmqTHWEjr07O0g203xbjixLL5b1+S
URZXM95bIbAOsh737Cq/tI/+kEXuebBD85YJW4aSOl0dpWjEpQBjb55XocZq
K4tWxGtpDVlul/xvcX8R37rkbVJ7/+srTcfaRYhODA+aIYQybJROBcpY2aSE
WqQoWso0biRvQa/4HAvn4u52lRBWt5Bxvy8jaJkuUCxkRQhnhLVv1XobsA2k
CrMvPq9BEyaoyyh1+Hp06ebIuM69rLfaJplVXsS4Agig0G3POEVNR0Ela1bq
mQosFboSeKPOoSV21bpCw5JMwCjZAuVhtTfdbKP3kDyOZxDiovJfwRvgY/Tg
c7qTshLAQ8A5Q+xlxHCmmd9NGsPrCZc7WgGGckcmu+lrKD39gb7KE9Qhwc55
fwRffeRT7bdLGMeqOUc1JBGIpF3mwKpg7ZZYlDtBef2K8pJIq+VUHEQP4qek
hY8GqpYDNuEFkGfv+ZfRPeJgUgAlsto2oPNQAhAwUMGVRUi5Bi7ue9h2c6la
DuJDpCuI92tOx6cSs6n+1g+Uvwh/hTlu4tuMwOhG+mtra7ybXXsvX+Npgsab
/b4DwlOsoq+Hen4/7Lien2ApfJ6czRSA78KeTs7E/cASz14BGMxVUyz+Cud1
VNuxA4McjesByDBebJlEn+VwNFXKnwI7krLRWsBd+6QW9xpFSm9kTy9+0YdU
Kkc9h0xLy3ifKyOwHFTNxAT4ucVeCsJkhiMSvwCv8vgYnTAlERGHGRmVVDc+
ZNTrm7RISl/d35g4Jw5YzTxhhyEAOjmXhGoqgJn3OVPC6SlRsXDqxrE7TKbk
ndshtEgBqA+M9RhtL+sp/1g3vvl9npM4Ms3RkdMfs7iYJa8tA9UpbvgSxXRa
RSkMGQdgxribtz5qEdqTNMg2LCdYVFh6EmE0C6k9JAMWxOfigarGY7sHXj38
szefd5gIn7rCoF5OWTNLS/al3fNMwZFFHMTWIKNjtxtuCLqZ3wiqIhUyQpeQ
xfUU7EUH54Ts6Zbhh+AMl1iPPO79outPMBEgfdjYcEfiGb6I42djQCJ2xtpE
0shrt92ZiP6tIZzjaq+lF4vPGT5pBve6y0tuT9dt69sU3nSfLhqm1CkX2sin
f4CGQ/WcWNZ2fLJY5QbK1a1p5JbTE69KRqJMt7/uLyZKjeKiVH+/309cwLGu
IAKpCSxl9xhkyOgBQZAt0xeAF3Xt/7eE9zmf2XGSNs5HCSGjpSTSh2HCOlJB
Tm69Y3W1gtW1EpVRWBjY0foq6ZEdlIJcPR7sVz4lZK931TotIHoxuFan7Vvy
3yZ4/nsVAiDPQqeoi5KP0KV8XGGeQScvV7x6pqXOe30YvVIX7JLD0rhHH9dH
b/1Qt641PiFmNjJ2J2mXX2QwbeEpTyUqMvK3vDagCFBQoU9gpQ82cy++7ciA
RJG7CV/1+Kn3rdIf1m+ytJLlC7LJ5cv1uKS+oAR3V4tATpA1ZUpql252AoEi
Pe8nBtNFl27/ZEEw10z78vt4VHt2A1bfgXyow09wG5NFajfF3q8D2xuCjYdx
fzSDmXYa1lZzbEFF1aeydxRpil1jcoTCrI/0Zm2tCs0EGgZtrxF925cuKJTC
TVbhKHHm1N4mYE9zCu+efJ/N1LTRz+Qa/h/TNwqvy67apKYUJi/VERSf1cR+
SrUg5+UG/yyDZPc0qM7ymF1ghJYFH4K39cOwDS+Y66G5pOZNRae5Uo66gi1G
LYt9bSYmwTIsANFxEibh+3Ycy6ez8w3N/8vNomY5XsB9YLGZG99SlyCo4tHo
fakqJRxshquAppldEje5VOmn8jwj/M50eSTgHhQAM3Dct5ddQmghYtbc0ema
5e+quY6CL0Qux84Rh5oE1KyQSHY8BsIUQZIOCXs+khxPvqk3FutvcMu8k0w2
9pkbXtmCZVA7kbEKuHPQzOjnivwwu9040QhbzbLc2tNdHAd0kajEaIo37xaZ
Wx1h2llximNWYyhrGMs6l5vBjVU+Dnav/AVicUNAqdqYHwP+YVrrmhsA//CX
Iygz+1sV2XDOL/ub88r+0m/W5z/GhyEkyuYis69K/O7vrfD2SglMosCdExTM
2SNN+cPMkWD3eLvVKYXamSMZq+Nvs+QJ0Pn33tTwjqnwEj7LwKiCwWTDN9gx
pxAkRT3t06BQrBNNNFtRw05iOfFbVktwX62/uLFdhWKQ+t1d0xVWBjcRHhW9
VcH1krhBxIYook+JdI8PGwxKhfJlEWdK+QMUc5bPQIuoHjDMP/fyX9i/mtXE
os9dzT2BZPLkqRCRfr+ZTRKY4q2zhCd9uJZqbKVpRhtTf9WwUoc9buxItu1w
svayNe2XHvLYaiJ0QwgnLcGxAWUsBu6PeRpdk3TOioHMlkPurFpof7qZ+KxI
IsxDZq5dMUb1vZHbvp1KxKRvcad2dJO4L4k4QbQfWfNBEG8WEPp7tMdXbaOg
CNpV8NEc66WQ5UclONGDhdGu/AygJBDrUKaazphBHAaxfwerkikDu/avoDlg
fPZ6C5NnEApmwDTaE+m5phf3nVA2WH7R+DugXNVorKP7qN/XNGvfmHnX3FJN
6qP/oGHbH8QCLYh2HM55zHgRnzlqp7i6NI7HoZVkrEZrB/UEckKgYoq06v6a
dDGsHLVawMCaoFFuK9ZOHSfLw1T80NN/kKITb3aznhUIGlckqUSs7Aa8JbV9
UHWKe0yqTHb6af2HhgWNwNTg7Ru1VVmnWf8F2cgj6UB2T0FmrI5AzsP/wPFp
+h+mDJY8Ng2NTOO3wiHdj+srjdfs7yHFOap0sZ8eAxsaTJU1cme+Fmm4Th6S
C/Rwij8LQoKVbiqXwtWfbuYU3ULL0D3iW+vKbWrV5NY6qQbkSKNJbX8UgHQS
i80MV6y7C87EF63DHNwzckczzbXq0DDDxWlQsUcbfp0BkuplnFhNJLTlmojy
iNbYDhtdqedBvlXL911EIKYgZK2RYzxQDey6gECyoxOTpgquP7slwiBKgd48
A2G2DeLzogBwgTRAhQD2WIaziz/oQH/U+o7g1uolBF5Yj/4cl86jpVQpXD8j
52Dd8d62JcZvtH0pHOS80aGFJ3nOd435F1WhgVg1DjFoljc1D1oOHKGLN2oM
/tETDEL5Bew/D8PawHm2mZCVMesybn2FhtOqjjOwNWogodqs0xa1c58ecbtY
MVWlov1W2Z6Rvf9Znts61NQ4giQVGBIkwqssS5Mh6/Yz4JfrlHSl526zkRH4
MxgYwJDdwptwxi86KAtd5L3/qZYY7OpS1xab0bi0mtbH4vKic7KFgOzP6jQs
gCQltmyc5uMNvhjxICHxgjFLc+e1tz64omekJ3q1Eq4SPwzgKQommDR6UlB3
7K4x2Q1oL9jbWhqq18w7JknQi5k2Z7uFmUBmb18eWnQBKyOs3XOeyMzHOMTV
TsX0a9R919bUFE9fbU395TtEKrELCpWQJFH81IJp8kAS7Yx8A2ZuCgIq3eP5
uguEcF5Z44GlHKusbZoJKt5u5r34cqUte6m1xoJoESXG+wP6A47TbI5SwmdA
h2iSo0mf0GYfBNB2DJdMo7bVLZ9cKADUNVs3rXU+P7nsLzd80PzzdDc6kDL7
8U1ydpovikdt9ei0voTtHq4rRin4eKxup4p2cX9caG/jaXzYkl58OvE9rdgQ
6M3hcpWfEF9Y4MdGcNADG+P1bMjWyigs5TYu5G1wSY9xs1+UMHg5boXNURhF
q5YIFYBH56VzZOFStNM6/1fgSFGWMwapXtfwrj0W3Z2TUZ+y4biZm1L1rLgK
dq7MFL8o75nMdDohRA34qeKQNFCF8qt3jWGcTZe/XNhE9RyyYprLLnLxruc+
qTkb/DR3O44MXPT6YwvWsenYiyeqpdU67duLfUBgSoWnV3fIBsgwryJceA1i
5U7Q1h2Xp1EW7ktgWKfuY667aBGeKk18UNd0i3vkVOfmOKr7EEdUkiMG1Dhi
7gwKNOgcjPSYVdA2Fv434Qam32KHyOgYYALoTYOLlXCMFV5ka5csEEhLUJyP
3BfryuTFYONFfXIezt1UX5b4kkDhQvNIHnv1Z7X1EH1mVs0G8E/YDmJnXJ7A
3sgItXYkhcoCRzuR8TvEoR2ESHM+iRuqsOLEPYDF+jcuycK7Q2HKDwuIQjg8
XmFuwS50XTTJASw9Gskx13FnyU8+tEkHnRpWN09ZGzC84vNmTQpLZzwvDtko
re1ztOahoWFxjwizCq9xch2pBtyinTe+ZlAxEnItNSyiKbi8H9yebORi/RyW
JaQWuL8CM2vSKOH4IWCVx6VwT1PwCca7jZf23/kC0IxKNym+WCmHiVtnyHhx
PZcVEaArlP3uBGNHGQGsu2P7fb447g2fL1NUQ+peSAqJWZsm10Q9O8LC+ykX
7UWlKxnR59wYSyoLih7oGp3WdMx0t+KkNo2Jyhc89RUswY3hKBTsMcHd+jdy
YHybbyzYLfQWr3KMSt692M+0tf2rm4HXj2/vl6ORYbc+ouPFnR8QFkYPlmyW
s5pt99tAXINCd08dmd7wSs9Zd6mlp5BNt/2RlR69BGoMxTHQXCnOqvYtVf60
W5g0JnN+DS4pfaq+VcEkmg16nlh10uaJ3o6HhbOmNOkFjQ57BxE5+3K3WM3F
iu8opVK1+JDft5Td58CdRexyc8Jw0uM3Hg6wx8ynbtLV6UXszjhon/upTD7l
8DilthGVlKGg/u9jnwuUQJ+ehxs0ANslo0yrOKLSAo8a7OZu68+VYy9/4KmJ
1VcpIS7K6f9sYw/MsaPEgs5RWPJuEAPa5/xEQXKTOuXZpFTgtS+9usc9iRDV
yk9XGK3zbt67po+QFqvJeYziAKi+Q3yLDoDEfwoCNUWMAZBgVZgoGj/oevez
wpUQfHLxJ0z5a2Zqf6U0zIIQzbtiVzk4QjNSnPLflj5X4cXgHJbApoy7f4Gr
2q88ieFVWCFogPjOlhdJBTaeRfPbn5qYq7hTQUmpIjEIGSBFxIhtlaDCWZjt
OITZ8JJdCwTcfIPYi+VanTpRmU7sfdjlnyWucDNwXppLoyS3tbzKfmBaOS1q
MP+EDv9o416TzKsIKT/GvXxcRN5OtAEU0v4AQGF1RbVYMMTAWECUsVyGEpgO
RHwu6L+fL5gFE4Ierj8kOqs6lyfhE8dtU2Lh8NH0VJr38vrp8HjdB9koiicT
bESuCte+EjVrtTa9o6AV+lzZbqHA2a9G33xxvow5o2wieM7H1QKExeBRiDbj
gRXVnpaudYrABh289nLaagznvUpCyKFfaS9y4BJ4+NKJbI22FiIEYE9GxS3P
x7L3lvTHiGhulNjmfzMdtLIEUjzK9tXwhA8Eov6P/CA7h/3sOErX1F0K/Fu3
vlcizaKOUduba8vdbBBue4LilRyf/C2vuWMhao20xjwJKhWQpr35rAKchaxG
3gGF7llAXbLTF6KqHxOx0cWcgRdVFfQH3y0W8Y1rIsnHX+DAbAeYmfnByuh0
M2E1JOBMUdkVdOSMwe/2AqhUbqpNRfIGInJRZeD4yymX7C3dbtQdEPTDp/K8
ePI5VTsaeJdCzZQ0VwHQM8JBm2TXtrJFH5d3WUufn9TWQxQAQas+7/t+P6Nh
HS67iX2bJx4q7zRmfBAUwQ5G2mO//51HWkEbQoWhwJNHG/G64XGiRv5Wq/8Q
eaSesVXl5cCadeBBNf4+rKVNF/XJOU/269RVb39Bulu58inuJEcaeoxgJSvB
PJNamSagGhMWMBLE1wg6zdh3hY2wq1axr2tQxbXpJB/Lq9HD87ehgqtxqoVD
f75pzWXgdfeNHpPJvbilpvhz9X2rVAsdSnDsjubnRjPRQFhzmnQwHvHTr5WP
pb2ebl8pY8lW9ymu/acCN5aoMLWQDEYEmuWg/G/GNAKL4CWjZ+2RQ7khUsoE
/FFw0B050NEP+49Sd6cL2/g2h1u6TCyfxr91r94I7CD2o/AujyiuloOVT+Tk
rgvptNtmVKmadLLzq45FMw8oLSxTaaF52+ccR5sESAf0b6q3Pc+23WsrLk2b
PkMo1HeB7uNy2UZK/nPFD2K2S379TYskw7owcrHTwhOSyMmdAZ6wJAGk5t4M
1chxKPrdzFlclH3lXOzU2PQXW2/rZqiDkrkzJ9hSGCEnql1f4JahHR/KP69P
FVfqwdzTh/ZehflkWFSVnQm3LzP1/Pn3EL2syi7RhFq7TxFRYpt4OXGl9oSI
L6j+JiUg+TZNoHak4NL5hyMPL9pR1MHH4qlZJ1JBVRUqUMy9tF4K18Mo8Fr4
Mz0Z8ywdB6NA1patkgXND4Yz1NehDujREPZrU8rWhdDzXghvR8YHYxFh4kQl
9YSZa6l5WMXAowIaMSkvQgMfE85qmUTUbHTu+W9nKh+b7l1o2pXaLisxUHOZ
ncUBb/LT8l4mEDYhwqtO/7hzC11V5M15UsAUMJCZMkOtlG0ibpYFQh/roOA8
sDL9gXiNgQ1birqHVznBv/n61VsfkFNYIwPjnGtzM64ElaSqFwLnlyXtq7XM
bjwDDGfl8gLht4oj5mQRMreMiNkAoKerpXgNWn5S04Cz7Se4H4xzlGsaLAiD
OruYeDX0qY338gfN8xsSMGwG/HvosCVMEEsk7ZTAlC8BLB2gkSGiSXrhUDIm
FYu/Zu3Jjm8gfUW5mhXsf1Y28fz8+ozrb5/2NtBZVyQB/mTrrClVQNxce0hA
rLxrWRItJBmvqG+j+TZG/fPTHxXioUmq59u2+0eMPgJ7Kbn+4bxmvCUic2dm
7nv9RQ60WDzzS5TnazRzQENBYc1thgh0YwiSmoNJeOuD350jqbT5SIsRAqYP
eKRRcYxbxriQSJQh30XEdNVSso2xHwEjOS9AxpYWTtlzfSjvTbCfCEBbG/jr
ouey090VFioDXPktKx7WHbGiotnzjl2NU9ryQ5prQARjZWtgSrJdd6EG+nnV
1znoacHRDaJAewfh5KcIgMZQ6MNm11b7g4/9cqAZCQRIKyaj+mgqFl1gbeVs
MdAzI1r73Q5lD6/iOT2CRpk0+DKt1g29PAhHyGjNY1ManE3Y4OeOrC3bbkAK
Ot4UnNlsSfbKfOHvPsiAGrHoJQ5rwEbnAdy0b6GLAEtauppTRjporxASnXhe
wh/gn+RIZoWfaY0tpWqwG6d1yc/3QYl8uepcMyQDmSeA5fqJq4ieQvex1TmT
XOo4/vfgIp/0dcw6A+PNX8DjKoq72Gm97mcVv8ijf/LUbuLIBYNL2qgUxp/O
hs0/YsagJ3t9nqG7Qt5xdXZrl913o3oaXlGbxiUM6xeyKQUx+VWfIvqr572p
22p3idgYB/GqDTPR6peOAYhFD1drekl9bv1VMFWcacHeV+0DYoHM3qXfl3kC
zFj/hBOcyAWCJ0DnSrVPf/OfGbVJQjZ+hx7W3FZFq434Aq1yyV6SE/82Lode
GpT+pg1aoUXWOJxzAessUiTwfW/Gahea+rG7/OkQYCt8VDWM7SN/+vkrN3Zw
5Aeh0aswIyGfmgMj0kZeZkU+GyfqRQ7ytflqbwjeHTCV7J8Znh10exaXC7vv
HAvWHqUZbOxMJheAml0tseAXl0h3HydA1wGio431xTposUoii5qhYNOFEbNn
P1uNat8Wf4R3TwRsB6t+hXOJaAMPE3fp4nbNLgjOB/Fmi3iYdgRGRyx/R/Sz
v3/P6dffvXQtM9fbDWLv8rFPDxk4AVLCUmpoPhFtE1QblJl1moDJZZRQsPyZ
7SEidF5GvdUL8V+OxcLCUv57AH6/MqgLngPDLpQXzGQSRcnzfdclSv/d+uXA
OGatA3dgrzaZxe9QMqpnZnMhrsSUrjinJcdNhdMCHp4r7lKUJPCSw3gdyA0e
RB+UP5vnuuHrmjImxcSSq94wG+q9BUiLQQrGnY/sndJaTMLE2xPR/81DY5FZ
nCmU34HnOAmJHGmdY06JMcG7ManSvvYUtS6WKB7BO0rHp7SeXRVr5+mzw6d5
gwZBw1oZ6FTqVHAD3ziiXWrgggZXPbO2BA3Mx55bxLFFuEfgCowXC5r673xd
MxEjpXwKRSDfJzNBhybEBLPStnoo/0a8BVzNna/lkbUirUD/cOhC7KMF0Kf+
lO5CEX9TEuP22uATef8/i1TCldY3YoeF5zWpQb/dfYpeDnBE+p5AKvbcIc9W
prNAr63IpQZ2m8vK3yr9dsvt5UEgeCyImlI8KkZ9DX3gFxqGvnkGSJkzCgkJ
ZQbau8w0Cbpt+BOP8eindW/s0lHfIuB5NmEQqg+gtyTzYthgrP3DJv2glV2e
WE6JfrqTWFh3Sf8WRabnNbfm2Uy80sANb8ErkThPEI+JKdEl8o/jXg7a8oWa
PyfD0k4Erz9OlPKEOsuzRXYk8JVf2XKpj6GtTDL3GTx92HfIRfG2MNw3Wcae
X5J2TQLqhODtjzmfsWnQhlI0QXOuNKKSiDQhuSX5rmlrcnziVDO2ZtXjGoUw
P7oAtrxYoaL12BzEefUqm+vy97Mv7MgTVIJ6ukmbezYSUU4miF8+b7Ur7J9I
qjJs0HqYsJLLsMJAjDvKrayJM+MXarvGFAlCE7/dLvIBo7NabTKF3+mMeGy5
ux43Z1gUvvNVuNUimuSVYSjfVWM2lrERlq80ux0PObOJTxBd8FHYWltUD7Rs
hFc4nAKc+kP/DLT7yKwrzoqNRjdb+vGSqQMwWNfJwBTW5WMFlgpEEOlsPXtX
aHBRztYYeXPm/4IlLSquPF3Eamkh3snXcw6lBiBNjqxG5cN6e9vjlLwUudEr
3f4ikN8L1zP0Tvst6E2l/idWdFtoB7pKOfYMEiMOXk5WCEoRJ6MhXGdclRnR
QT8VXDtYluf2Gy5NTNZwvo9l9YsxLUiYTRjyxuxfB5g6r7mNs4N/keG6t6Dc
b85Iv7hkzOsuyrImzfnYHAi3wYypi6B5WnEYztLxAK4omtVEgQ9Ot5GZwQyz
U1aG9k9KMktZ7n2QKn09Zu7j7ZbTVU75ZXa5qUc+YUrdA1OpfMUusRXYQ32r
5b3wgctX2YDiAWt08IpaCm6tSyklfMej+BCelpDbThK9P3R8VDnWVSunS0B3
ZXJzAfkryYOxLA4c8P/QMtj2e70uj0ZKgm2fg0z1k2IwXPF4k96i068QJM0e
zTFMvPfH2ESRCQJkEMeFjg6wpM5fxi/BcsHuZP/9+haAEG+q7Ry23XbEZ2FG
KD9ay3x8sq+ZZqbYa7p365WoERXHcG2QfRzSYiON9FslZ0tK/rNRyCvr+l05
XxwsY8W+tLgxastHsKd4rjZr9bk7OnuMtwzyUMBRvG8t7ri3Azbw+w0brCwR
5tB1txX2rRoZgxrzKvrFlkHrXyIXIWfkppeBBbXeW/AGkIEGaXud5TB/o2+H
1CHGWwk7ooW6fFzUrAMhLhXVAiJOGjaHbbVAche8DOb1eZ7neScy2L5j7GP6
pbl29pmsEX4reSnTNulFUCJco+4SAIuuWIgMS12lRtMdyQqleaMRVrVGRGJH
uya1pcQb+W2oqAJ1HR8U2LV2mLp/WR4eA595Y1rTklh1J/lzFF2t7a8Tud8+
iTQNhvrjcorHFZVuawN9UHX58MgONiJz31V6W61AwezSDSHkPFqRV5dSjqLL
JSNhJ8153wZImp/Y1YhESSr6M+KzvB0wdYxnxcrzqh8trBE8XY88rmpr90DI
tEdW4lf0PMiikzxQr/AYPq0WV9CNQMhDXjbrP5/rcpeUJIr25lifwuhBJsAV
apQVkmG2283cDKAXT0cRo2aUKGDssFy3CFqVB2wH2QITI6vSQIG20R7oUOnH
mJOKf0EpyIVOD+PaYBNktqzV6mFe5fW25+zo4azhJQDb1o8BGOSsswsoY7S1
Z8MsvdDOxbCgGNOMFmAI3lhT9i4VkTcvlAxcqjp9LJZ4IXIMWFTSBBESa6Ns
Bj0ivyEla4oj9wUtuIYf1uRsFwZ+BG8ETaSnlW51j2b0v7uID2sGxCC1/CQA
iaaGgn2XwrJrbU5dPlcK62s2PclCh6gTLuRvb87htHLD7fjIVRJcvfGw5B6e
cy0rHb1Xam7zgBrGJBM8+a3Fih19rt5AImTMR+v4MkM+W71iKrjtrWKpuqnr
jQm238Yn2ACUxWvCwEUnKQ7H4/0deAax+x9FQ6yFv8859SKlIviplju6fGjo
1iLFJ1QdhyCO1wSMaSsJWr3mm4Gr+1Np/TyXjflH/f/fiFu9V+cVz6vfq3BM
fYED+bvtKgpBdzcCnWjSBRbq4RyEMyDXjNcqVlkk5qSBar1EB7foSIIwCNfd
tIXOHQHu9MsfcWKKAHjGUNBnTbPJNi7UKvp3XmZfi+TtzR2c90LDdtjbL3h1
CML1KeOJmU22iUmC+1d4QvdNr43BzG7tJXC5cON3kIOReOGst4YIogv+SfNe
fLi6UR1s03gzVOYbnw2K/tzqkSCNl65NAPWpHcf5eURIy4n/bnXu1tKMCiT3
6x2G1o5UxZ4BghkVnL3XPuPScTeIYMmN8haw1roJtmfBnuTvJ3EkVsF9w9la
Ir2gU/rlu9qOtEa6hiMm3okazHxunqyIw2lnWNGvqXKFUuxdTyS5Joj/ahtD
zzR7Z9UANTDGwDJojMxto/xB0U0mTI1HeuvnM8JuqF1s17U6bRbiQ8W003aL
vM3P3L4bCWWY1zhH7wyJSppQ0/lTbXY5rOMsJktNM058ahR5dakV2Fv/xltY
xCKC6J8osYidB2mWQh8IPotHTgBAfkXd+xIpDYlLvVZrN71iaVLJGEg0psgY
5GvVRKCfgqsF2f5bstHQnNyUx4ZRhUcCHn7Vi+xrEXlWQ8jU7Bczq5ZmL9Zb
FkuF4YdMclPSyh1q9obx8O54GpImpqaj9py9CfvJWUD+NnRjATqAUMkyMw5F
xWM85OTDgVkq40u4gvnUU1rqQwTnEND8HhVnpGW0pKsSfMTmOhkgsxj5S1fC
P+6z6opRzwCAQIXsVirQtzpuNI+OTk5MZT3gl1R6BkltSGXAIp+vDS9RDY4/
xDj2J4uYNo5juGYPDDydHFjH2hYqeoW7G6VoksvezuYU+dIC3fd1G4Dt7HMc
TYZfYmxyTOuwrzjggeLrsplCUV+Uf2j92CXFp/1NhuEKuKgjonxnidx21Wwb
ZHaGohN8jKdyfptchWMNH28Y4Lc31AAkOkcpefEnAJiiLuVyzbVy443r/C2f
j4b3TEqt7/JkO2COtuqqz5eRCRiVbKKZ+roRwUXUpU12C5pLDtK6PLMDRRZf
PtbKFQwXSaua1w2eC2mRNx1Tr3n351IcKi/FtRBTKir/uM+uAzhDpScGJqfr
/i7NcCw/vPmrUjaZBdJ9KNIrhrdvfmpo5Adh6r4cc4yEVesdr3IzF0LpTsQ4
8R77pxzOZxAae/ZKOdUyWVghn4CnSRtlGlI+Qjl2Bf3iWmtCZYPS+gZ0Xx4a
dzSNsSzDN0ZXHFWyNzlULqi9H+kD00RzAlwxyOpk9lDKrgfNpvXZYZvvZjF1
UAQfT1EntOuoluSd/bGvfuoy6a52DVBzZMTKFm9GPIyAs2w5cCFNXgB7Wy7Q
fTuBAmg4+T/10zG6IOgjIYyCc/7ZD74ZaFugQO8NUmGezXDqg5Fl+d8ahAzf
0Nynrm09anqDgYaYeEGrFy428g6opyttkN0NWPuMDcqnpESt+xazg5/ifigc
u+E709JGOThCEQ+XgacsOHeuUdrE2qVvX/pQiT3/JYbNI6VmqA+uQ1WJEAcj
BL6IAJhr6AtgbUmfN3o9f28a9ezJjDfO8B4QJJNGtOun2syVyxf9etXtRN/N
2hE8TY44LTY4FZU79ufxdsH81H9OERttTROcECo/rdwYAR/VHssf45D8rq/q
+lM3xCyhx4ulg1FONA8/0lz3OxDOnOi7Bv3v59oR/RSoOYfih69KGmgyyt/h
BTZR+Ov7o3WK3bFA5B0ecIyDqB5K0Pz1KLSUdK0+R4uR1gJACNJRDZQhqDpu
GfubUzVJZM3TyBrK4c9m4bRrRml18qEGHsYimGmRGUIRsdiYBh15Q2wpRtU3
NiRMVjuchWAGqeUmHnrkQxADxdszpoDkgTeq22HiCufs8n/KDViB8DJfnfH0
9Dj/bdTwsRf89OSPPAhhBC73cWpZdxOLkj+ttfsQ9EHQ0aq+OAjetMvGLBWO
V8ps8WD/E5nSIwRNylC9/aR90SHhqJHmPtYARGUK8dkrrW1b8K7HTZi0SJmX
wdfHoZK2KcQ7RHr7aFr7m241AI2SS7IK14Wb+ydC9x3+RMcanIilj4nO3gbA
WslqWyV5QqAgeE8G2EOOJza9fjUVWtJh/J2DPGBQr5gKArcV1Zg/XmXWCuUy
Dow6sFjvC6STIQdxMDe9I48EefQDmELM0BEUhdXFyngeUTnwR/bvIWVTZ9lK
ho6+U3jlSQzVgMrCuo0R37nXnNr/tH1WqLc91eq0dBq99Whp8UzFLUQ6Ca5S
o22vs3TI13VlTO1DQtvWa1V8g+ce/EL/43nmyxVuB+jGvnYD1pbz9eLxemlP
wD31emYdsMyXbNA9QqsreCGtJQdq6UK3r89couUwPnDjr8OAv9APaU2BOi7T
nrlinq0lMOnPLPpdWH8DD+FI3QDqUQ88KKYtx26bGFZqB145YrvEsTWRZ5Vf
tb3GqFwlcMiPSMHRUhPYcCBjfmaj3RODepVqqFpM63iP/wEoZjQIkFuJPyV9
ittPF17EJDBwD55XUmyZdXYoOEFuHgZTDhcIN4VaqQNHBZZY9pGBvbKZIaoP
6w26xF9KJT6TE2Aioy8iU37UmiwOorRTMaOnyAT3OF8hfQwJBg3D5HBrUYc6
FVSb48tamtQhnRHxOa60/lNX1Bz86YiVbHZ0GrOqnaExtMgvh32Kn0c1YRMm
kIlqcW7eUh7oxb5F0zZotcQMAlFgocntlNWLZ6mS3IbcYgLlu56JOtXfF0IX
FWnnisg3HWcGI4yYg1qsCByA8NA7b6AhzlL9dJjT3eIuPyfddx63Jwy7wdJy
zO8rILi5cy7uP9nQzlbVctDh/G5h0rd+Ua8HjY09JvYKRKP6SnqHj9pv2v5i
lHXB6U8hzVTWRi7yakyYSB40P8MmEm83n7eu6v7N+WLt/EjuE3gMifX/Vtju
NC6cJo/NgAbrZKP1uMxv6ii6hZcZPv9jBKCg4qSeSab8jq4e36KVUjmO/Qv/
hs+LCPC9PNVT8tRlpBLkIv6UjnXDKJbVn2+k8QGBCBoQSJg3UBss3KgubuBx
BCNUNAZ9vpnMIP+9MDCZIr+SaRr1LGqiLUfzWPf6WVvyFUKD9zERlSD07t55
afZZ5aClE+0HUFmR1B+qK41mnc6yGXEmvHtAOA378UdMIbi4ycnRzDYuUBKH
ACZwba4ERyOnq802j1NWyD/I+H3spE3b7WlNZDGF3FyqwdLx/0b4EtXb1XxN
9CS0T+gIk5boQshfjt1PSYRtoBVQ9GQ19NwFHB1jnj/sECvZv6cCH9osChZ0
7xpdFzj8mpk32xSEIiPUXkrKgNmfcvjGh8FMpdbSrGS5/UQqW8BYlVLaQLPH
AdeO82RcnChChyp/l/7T5BHpcgALf3eeeYmXMuyVcwnftxbE+TVcOJ2o1R8r
yG0Q+s01uPKxr2lMtT5Mi3QRmPV0Ayb9J5COSe6XyA35rxcDYOIIxhoPDWRn
Waln8KDthRzo5rUZs1iA0R4KrENtc12TA+88u+0I83CyEIzA21jC7t7fOKIl
wF4S/mc205ip+3ooKBhMgHgfRSGm+ZA6d2EHtosJr8UNcKeuJT7Wqo4o5/Nd
i0jhjsM8M2kfJEPNg1ab2e+H1Qhh5SZPK5yMsFtL0EQMBfBgUwgP5BSWhvS8
bAa5H8ZUhLAx4ugRrIio1jUxAdFXnVufDulghSK4DZ+HoFniIhUUwyVJj2SI
bn8fLF2q0KwIiDnRkN8kgP+crh3YoStE0Ec3DUlBYjpCVpB0M5eARuoEw7wk
d63MGcYdiNWv5s84dlud9f/njPz6kWwwdTDP3o/+9Um3+CLR3/BHO4FIiGO/
xX2hn1CxH8OTaXujRV/t6dlENOY2tHxZO0/1NsntZ8/9MHuROlqg5fn5AsTG
2HC6zcym5zD+PwGanggC5MXhly/CNbhC9WFT8kxQ0qhW1PTPtIjLxT8YMR4q
7+DpkS3CDCi958Kmvsq5Nu/E5e8/i/eExpMIJyGaoYMI7FfQrXa3Vk5SuW5r
N1sadVEVQ74hZ6JGSBL6ZrU9EG9UKGYqjfqWe37Z4AjnNsUc2GAzZjh/Kx/B
jnQSkafrxrYMM21Wfox2Wt+GCzfliwNOmdZ6oUk0uTK81BQhbI9TrtsryAo4
NKVUAFC3Ri/1vAwhMQRVa0V7sYCNHS1hE/y8sZy3JsOkiv5Wjq4L1wd4zuD4
aWyq15CMUbUCM5yPBwrW+oi2uAOAjTOKhcRFYXQknIUk/yUVttpJSKQ+SPwF
cGbLbXCQuJZ23gKTz/SZLRdtTlef1plYeVeK93UtG5LTkzEgDuTobkiMR7IN
8BwHt6obXq2GWQ+5YfDpMTLhgWQlLsFZs9K6d8NC/yohXBcnyspZMru+ucmq
Qtmeb/u5pbCNjGq4Ns0rltjTJP67uZbAHt8OgwArSwi7dVmFB8Aif/C68STQ
i6DReTSTIaTJk2fw81nnG5Ln0NKToCO5cupBPLoyd/Z2zznZqnXTnDnEx9wa
R26cjnplvQ4cCxjbx7FiiiEWQ97bBKJzYZED6VXLqjwOacF/GL6y3U8Chf0+
9/rxM+4Ozw1EPxz0e3gvKupJ5/1LONW1qlTa8ZJbNDLwbmVFOv/ErjV5uebg
SGjkf/I+g1nFY830LbdiHDPL2zwCxYhjua/uWjcjqSyobu9bgyECgxaFrbjI
QtCl/oTanOXhJZeQuS8+y22/rfxdLJUSfR0ket9X052TyMzfSq34iLj1rzv8
NPgqhIg0xhkSn28S/tpOh3XY+zfq2dSZHtYibscxa2gquHWseulBeaPmJbu7
UFvRpyVgX+VhZxa4Un6Tifekuq8rp4HY4oGhZHhLwivRaev3PDVp8AFckw0p
jANsKNZLKG4V9JCLzYLHx3pRRA05yT1I8wAeOZT/FfEEnAtgdKZeFZKCFz96
G3brNwX+gxIYCyyE1YHM8Cf7ygSoZyoNoH0F5f//VlARK8VMsZSdrurxzRmh
chP5VuVMKsrxVeiqMSiHBxsWKLnaWieubc8MepYQcL4JYI8XPxg/v7KW1qE+
02zaXB8Bl8AIYNT7rlJAL5dop3h3xqeDqh+L/wloC/tcMkthhtFhZiYJxKqs
58ggraWJFXVhOYFi4JeByv5EZQjC+1WibQnmHMI7R/Bp+pWcG3Z+csTqkuMm
SpjGIA34iAUPO93YxC733H6FtiWhVyiQO1MbjV3PYtWVYm93z353GJgB3HRC
R1Zr5tM/plW1JaCk+c3hoJMuv5fBwVJOQz2le8HHwH2h7DUB4z2fENRvwS+L
hFJapvtEqu1a0M9eDjXJCdC2fDVCBrj15UKDk19d2Ee7b7WMgTq6lI/1QBN4
/aX1v5YF7lO9PCSHJN2ClbvIW/8OIZTkbuXk5cI0Uzpqe5BV9MfkNoUiUdFM
TMmMplfJcEaapUmilLBknlaeUGA0GBMD9NyDS9Ppg8bQi5WBclOQ3KHrxpRf
wLEvRMIqQ/QrXx7eYj+rLJskranETjUo85y7IxK3VNEHaVS5ObNsDw7Y6pu9
GcdFY8Y/v++LXfeU8r0G0FyQN2hd/eC5275/6uJGfVv7xsikdjhEcw+T5WMb
KC15owj2bQTIyrB095sjArGX0x5GLYAT6xuJ/IfliYtCprg4jp6lf22RjZHv
y1vdfjSssgheF8WgXgn5IVTrT1qjRjayJQPEwgp5i9jXvdaB4H+O0RPbBZxP
kKnLn5oRAVRBqryItisWyT3D90QgfKnxyXV+JGrqkhxtGTKX2sYWUOoTo4D0
KJicEbECnQEwwR95RzT70BpE3zQYCZfW2fLFI9gagrRxBRCUuGAXegOm9yQZ
G+HLmwLvanlpoYJsMWFS25FpmDtqxz8fgm1zlbYccuNqRIYyI0Z8eBP5avnY
mQY5N8v+KxdMwJunx5GnxBsbSyfYO22eV9yrD+dD+F4ZLYiW6VZ02wYY/rMV
w/6EQaf5aJsUjOcSFmeQ0elCH6ZvNprtGqa1UYj4GViaDxxjqW3qXhp/s1/x
EtTYH4P+YIX2S5ganadT5tPOfFqXQ90UxS7C7aJ52X7sXXaAc34sUu2e3emx
DJKeYT3qmBJR09bpYzu8RHSrupWQpmJKKYuisKssuOyX/6GHyciVcYUCKcGT
hUUyje/Y/0fgoHZ6db6/Tc136RjX1eRQdheNzC8eyQLNuFlGsNxu7sCSMnlx
I3o8snFc/jJN9sMmOytKDZgU2cV9VKK96GAg+a2hhFOPVCZFVQM7cLKhXgMA
OPCs0BquJhCZLLSTWf6xBLPUt+QXTHIEUQcHI8AjilMTqSFKRksaVMOBkjXU
WRAhW6jfUY16uNJBsEU2jPw/6+5o5lmxy1PrW5HXotrBpzyMsWZqquPX7N0o
n1zFQt8tMo8M3R0+X4OXkTtFnBBUSJdz+3CtDe84USfixv8ZNzdLMS/JuHlD
Xa/rXkyRk8DCnEg8Mw60degie/kC/zoAaz48hegpMGLEapmbA/PXQqHI6ddO
MU9AMhQNYh9ragfM4she4D6S8pvvh6LLOl+h2iwcwfWiUU03h5H9MH0rfAto
HzEd7HZMETBhV+v+S+5wqpKiPQvp/3IhvRzMujmCVLiLjPdKELBtFyPCZDJY
scrsd5wznuPFzp26LTkMyu3OOXMSiAjk/gOYU7vSiXIYXtlkNuCB072GBK6x
8Xs/bTpbYwThSQ8Wu6TaPQ1i/GvYuDzEIN/M25SC/P8RTHSwoZNu0oaxiq6K
dSvFHC+MrvfYk1JQAMBVaF6tOp3RdvK+d3VUxrJKiYuDSDHPhuj6ggANny+g
EySA6SBX5em7k69j4cC+zz3duuKDfDu7D0Z9t7egYvb5JuZR61ROi1/dHq7g
5gZq5N2Zf4mLUrUJhlNOLFhoRsfJmDL8ETuPegkxpXZQd1hcCf4IGVPx0iVw
wdFXt/kx2VHg6aI8eXtG0Ddnv7q0Z0fYWw64V8E9TmbxPcz7e2cNkjqt3Vpc
+pEOAT6IRGRmMS+/R7lspVkLFzA1LC5AD9WkOfv4Jaof9cXkSxgh/o8G1Cql
U7t2xLbHtNOSD8yv4b0+nWnFZFvWL3i3uVgjKpFWyOyA/RnjMiEQx0KaRJ5D
rwQXjBCjTTiMBdd4Wr65cbEQzJBozwzSWh5+ep2zL/LHcEhJYng3mclzpsrD
I6FVtqu+hpUlWNCn3cnTxrAk7j7TbqdFupKLtIjO4g412VQiC6gUJ2b//TaR
aC0aW7riI+prhdkEIAkRdlphySTheYESjTAuh30IN+Ehf8keAhCbqu8CzHOR
q0ezFSdm3x7ghK2/nU3qrToHhta1PadarEAqFvY2JTwKt5w+gZKF4dyQBdWf
gdz5VeSPh/jnxBzdHnHPD5lXCZd6M8V+uT6WXK84TXIHl9DMLWcEiYrlRw1P
D8zIUNcf8/eRljwkiZOsSRDr+8xzSYADWZ2Wl21yKJPO93CS83B8qrfexvOU
mmDNuJ3Xt46pE2lvPjC4nmV1m6jGQuQ4cRjipGQPeBwhXDBGXHLM8aBeKCNt
o4aJ+/vGfNTPgplkT+YMNGAtJO2FJiwV4F04kyOiLRHvLilJPgOBabO4+VOJ
rrifNCC1lLXwZIgYQSUzwgBw5tdtSydS/ZkxzHQWOLpQXpuCfy0remuEv0Tw
0Vpg9hrBU/r1FJFBMz11bMnrlFdg5SdyZ9gqtVGgxYCWynx7pfo/GZUMbJwF
h79H0VBq9GO3hSULBM5CNm7Prs6vPDMezp8sQGhHH+ZYMAvCMZhP5B0dpb0G
AGhwC50vhFYC5EXRFdIgKZ03NDg7l2Zne1Z6BF8CJWtqJVjy5Hg+yBeaVlv+
26YPvp65qFdpXgOsi/VYd7FWNtcLe9V0fxjb86JFjGNBDW33g4iV1TYBQ4g5
SZHY7u2hy+ZXaRdFcmS6H0Vif5M2/Dp/Kaegg82SoFmC+77ToXmIvJQJ+qnc
EVjtfjOj3Ps38t4aRLA53NyXxJmUffZdi67UHPJBTAiggojEgFX9+YrEB8RT
UJboYOKRTEimngZ2aFHgbNEf3D24MuUmw7PFDfaol+ZsWE0svWOuHIcfXW9l
XlwVnoHv5Ix4w4eR8ggfnsS5CTtGFC9+awGk8/0tIkBgFJ7O6YzEsbcTpD/d
yGjhbaD3g/UtxtB0Yv5Hb1k1xjEXPLCkh95VeR+OWImh25XIqNkOl2F0aDRq
1RJfuqu9J7wPui6BOzw514Q/g3vcAxxSDWBw4pILAWNSQZQKbpnds0x86a1A
K+Zr2DQnjGeYa4t/vYEyN1I2ZFweuj7d1dqCh4AlcS9FD48ggedsYgGv/oaC
v1qjNQf+wjsEtxdv3iWMpM5zEZl3BggCWO4dXu4Qi4+PYcgUm8EM8sRco9H8
ow9dzckcl9YafeYne1BTN590Ry7uLyoilk4wdyvteaaAgMyfWtI8tudmhmj6
VPgSmZjgOJQh9oKETYLuEXUvaEGALvykA8I/67INHY1qlu3oXSkjpyr2fW+P
iDyAVzHiREhNsQLK3ZBP+4d3SrU8Ils3gJGn02aUbSM6IrglWE1xajQhaH20
88iuCQstwNaiZ0RzJ/sGXiLOE2C9vH7ZxGdt8NZNCn2Tfd87y83GlVMe2KjJ
AheQy/OFdJcwEZiJwCUXphtOQN27rbW90q0oWtgjfIo+YQwCaODqFXSXaVpT
RFI5oCyymvZSkI/yP51XIgUsrGS5QRkjB4vqb/E27Wo4b1WM2F2NjYwxW3Bz
ONWyvnauBYE/1aMa1fg8j6j3Qh48zpK4gJp/Agu2Oa2HKozRr4HluTI+ffLT
pdJUhl1FaftHfAIGDSfrQi9Zkr/s+DWvA1Jw25wONlAeP3ZD6tIkegUdAVhL
jKjJIAaOL1CT191cADd0Tz1Dy5cbvEnNBxrXaoGGp+OuHo3iAKzDCZDbU4/d
TCojTz0OTtjI8wwCJ7EXmucm7N7/Jml3k2ds7p95vU7HslV0ic4yJa2RBAHA
O8Zo8SqqlvdrCufJkkDYgmxkvXDnFp01gqlkRFfHcnYs2KuftK7Jb4Ys9/m5
+r91/zxfFwbOTpxomornce2o4NJ71nOwtHy4RnrGPquxLqVU324YgMr8mT5L
zudKi2cKf8aCKsWO0w9jGTXBY0wSyUUKs9N4fhnmBlFuDz99B0AMrF7Vj2co
I4sN+kB+N6kb+bB8WMowGmbDVrCdDY2aV3aDQWXuicDyZ9LmZbg3pBCzj3pi
gwYDlEcOyY5jrNAcuVTAKN7BpCMPRSiMW/heYzHG9EChz7nQqAUk5uCvV+q4
tzzBhBTtzjD+vawr5JbEk8GNM/6VTZvQQvGvLdOJO1FjMHf/XWoytAIvdcwz
bykNeEMZThNaRr10wAXhb1kkixAYcg6Yy+cXwwrIfSsvQcMUesWcID08Pcrk
vKlUXfG3ZcaUhBhkDEuCGGrmMqZegIgwOM+Hzjl3Yuw7QxYBUJuSiwYkCAGt
DyTAwAsgZsGYWAN/S6jO8PN029G4PHXLTJeW2Dy8yYfApyqQw5XM9fB3VQWt
vB59fHRnHm7IKk9nhnYA/0eCx5S65gwqnQCR/pnpOnqwiClXoGzVyWmcGbx1
Q3OR9FlEqhzLP83z32oO+lkz8Fw7Qrx8HMKnCUvV6iu1PENABrnRahCJr29H
FwZ0N3zQkI0VAVADYBj+OvsXoMYUQp+MHh7vG3f4mwC5J6kRxLpQvbU32QQE
JGZM4gLyaq6M+KAaoLowJwCpHsfDgTHAweTFqMqrfyWXVXX0LVK5T9qM+yd2
V41hM+VGZzjY9Vu6sJoCHommwY9t/4lbF7XVfGg3IYbuC7lxNvoKjXDB/S2O
uQMCrGB2qWzV108aCNKh7gXqz1A8gB/5Jupo/RGNEybWzSQcJVU9qkQVQ4vP
nOmWaXmZlr1y69UgWk6jajRUPELNLupVJ/NGEUOVlaMfXzWdCSk1HvLPFMpQ
KPdLg8A/C7obN8pocVB4kMTd84n9M2X1LUWabJDVBELuny40+I7QxoYQ3D1v
D+oY2Xoekh6aY4DpZsWchjgIE2lIb4lspF40Z9KC9nYQzlev1VuIZMfLSgez
wF7MFI6h0vIMGsQs897rEIH4zrrOe0vA7QZ3QBYXWE9GDsGrS9RqIaLPt7hT
6sG6a7CB2/kWMj2x6JyZ48LWz+lCRQr+dFED1JgcF+THG7kfp8GdyaJ3jS/n
uY4CYt6CmWywxW9vg9uKRnlc7FYMNN//QTHP6qRKz0m7YO9lnS5wLmAk83+h
Aza6UIvBMMFoihCpHg4++JhgYTnBfygbAMTDg3hZDON4f54BvzNmzYhDmMe7
7AcL4uU0I4qqSe2DuJ8Y+mvzs92avHXFGlgt0ytVBkCu3ojXHB4hMYexDUJ/
x29080MsLQwjA9KoCzSikSb//TYywdh7HKIBywqNcoPTaMwNWRGN+rc99RRd
1EotODaTCdn1TI1DNqtzx0uEVMKkATHDGSVFSVmwj0JHciJDgaw0DB5GlDzW
zRRhdcbwdsqmaz7ELs33nLP7NFl1wD9xWwRZ1Sdb+jBXbGUR6YFwF7RxYdAA
NbtpvltUutn9lX8DNG9BptpXiPS++wA/ARj7g4XBTIg+JjGCUYQcETrT5eWF
p7S/7P0u2wfuIB4RuTEgIVWTSSsEJCfkEjb88J0FLgotedeJycnjafezVDsN
8MUbtdywbNB2GgTNfqVRkD6wdhBVaTceQT3jqH2E3L/gowSvNM1XDCvollup
4IQ5NMqqQrsmAo0Xib4QmeFv0FIva4Cfl1LV+D6xqefDWqLiDLTVjKXd1rw4
xjNriOD/faaQnrVQPLtn1yNWOJc4mrZeRhyD2GxjSG/9sNkVbQ4NW0PBaLAq
VC3gYwL6NKuZHxEqcgJc6R+UaFR7BJ9GHPNhVg0/pevV38/sCcgsX2+I6fdt
0Uq3+j9yxCLuKj126owXP+tAoLiCYlfpZBGNHaDhSgaw5Bm+wYJYXIrQ73/0
SSWRbqr05pT0jYKMY+szgz+vcMjN/PAcD7pXLfMBHsQqsuAKFWSeOssUb8W2
rRNsGVbwal+mueseACo/+vTnEHg1vwaN1Na1xv+yVtmZMJRnKU69RcTuqpE/
Jd7SXaZiWPedREb+YzHhSBwE/Yz9pB/+ie/23UyQqFBTmISok7cZ9ZJeMU26
+UTCZEtuVkRmwdxfXIdOWAq0LgW9NQ8KJsR/FtRDaopelMAuZrdEQ1IJ3a5V
4aS8H2Vi+YxbDPybdjrgrYXhc/9Y8Mki6BU9mbUedEz9h3OV6RCiy2QF2iJW
DfeNyC98dNWp9sYHeYWnhNdERCwPxuKdbPobSagg8Pl416BXYrKzhQ9DOCxQ
GJrKbMQMLo2Pl8T46QFDC1xa3iY0eXVSW4unjhdmpH1GJmi+3OWjKY5aLiee
Nr8h7CBzosPCQ8EUfJ61uvCz5RgfCIbP38BVhJ3TKmXv6Y60nwSefLCSElPB
ZQcg8B2f9IrbbRoJgoXIJ0AI8xzK9PMyJAApviMo99XXhcuSIEQ0dnJxFydC
6owj7Ole9nWgvVhW5N/qjCO9XzniNznizO88DsHwtqy3mE5RWTh6sV0zceDE
0kVJYKIQ20V3tmKdEntoqQvkbNFL7nr8W9whC/soNo13mPTYOs01v701PZ6k
Qxe/zWW8RLPLn1k2JrPjyiCT7wbVS3/KR5Tgm7lAivzVr0FgX9cIRSlmpLLa
PhE38mLObHMDA0/zl4qSyHq5ORFeGynagyYeMiYRvgAlOq1grTZM+sLIxSSK
Nt3sOc9Fy+TKP8iLW3G45lAP41uAHyp0oJRBzB8dJdFQ1QhxynslqZJQHUqK
Qp1ZpTaokF5hlvT3CuXVwAFedhWc55lp3QqMIsamJBrm8dDJNpK0kp93HQmV
yYZGutohVaMeL4J4WuH8swP82epSg48mB6Bct80PIEFmYO3rXwRrzGjKW3Ym
7yCua3ESHOg82bi4Fqt7OI2c5+v2E1g89PlYJcuaYXGYaGBsjNFGbiCaF0D7
fZ3168VRsLLv+3VKJdPZUoQ4337zc1wAn3qdvSTJ/bG2FhLMNVwxSVo8ChMl
sCkDuzJzAXBTfS6MsxC6/ULwaTI5AuK2uLqL6Ec+PLkJ+8G0nWtoYSCWR8Qg
vsvb846PLQz27WynukcLsWxlYSYwXavn+c/OyRhFVIQwE6qFZzJnXsxfFQT6
rKe7ND/1GYv1NSk8gzcePeSdeG7qnQqN8++T978jMC+32iYGL9Kh6qDDc6hk
bqkbRloPWGk2G7KtXvfPFUYVnhLK6o+hoV66JLXos3C5S5fjvNoCEALfhQRd
qoORX7VmtAnW+4ENDOQ/TMfJmYPZ0uI9zL4cosGclZlkVoWyb4AuB9Op32+G
1uifurhx/wsZKZ+H4xL9mr8up5Ni3ukrfUYJ70faJ0oCZOOsr8S90wfX9NjJ
8zywpMWd45+CwRpfvGgQeNe6bkug5kQ0On0+JqvSVrazyTJNBBG8oUAEo95v
jnas3+q7EcuiopMRuWWRpL7i44k8TavlYWNmdFlOpAoZOfyjmDdwERRMfZ2q
8OU0fduquORMYwauvWvxpSK2d3XZ3E9bFJH+UjOrda9qHtUZFA7ELG/v4xOW
BmxUf+umd48YLlNqlUmyFyGGrPgCG0T8Vuz0zRntt+nJYqMMZ1FOgPUKSkqq
hPIajUadjGulz3hmte/JRyHz84ywQgy+SKTWC+h94im31P6bSovYVYsDCXLe
lsJMkyzW+Vw1rU2UsUAx5wm8giSUoGv9rKa2FvKCLybbSq30IgAAEAtqnk+u
nO4yl15+MXsJLlFAzKDPZe86BdqzTCUhHP+hmohMv4eVSzO43i8HieX27hRe
mcVBVLjYC5XKbfjeNIOFD6QPFAq+CgUqD90wYhD8DDejhloeECfqLztM2xBG
ANmV8DRogxSTV+nUb9m3YmH8ehbAJH+crf26KQMqV8H00Yaobw/M5MNDakuz
7p0yMrmAU1bbQNYok/QZGVvdH4f2dlFyAAO6qKMNfGNQw2t7WGD9AjoVI6mH
GPN8HDR1SsYszapfQtJGETec/uqNhUCVsBdAbn2XYuDOdUfPEvPWRHohEqPB
CGjvC7TbVi2FdVUS2DB1qzYiWEYMD+3gUToMeN6ebWX/z9xt2pI+FAuofGjW
p5fiyL2RdygjQukt/dAxFev4V6fWKt0xxs1z2hDMbwZFcZ1ZEiRABONeug2L
pmh9FlRBb12DTcfFCsW5wSuCE/L4DupqFB/dYdNg7gKUHBhnsVRIhbfznNBo
RUeM0PlY+7vdinju1n2kH4QRwHq0TNuesDHYLFC7J7EvjcpqVSJvcJ8sD+7s
/YT+njIyipqJXjQ7kkGw1gz5HUumEkKIMgbYVwQaqoGzG0Jo9/bUcI7bjwMB
6A5EfhOni/dMwn+dl4ieu8+etCOVSnUkClIkA5JHDojXdmuql1L1MwN5P8i5
nFeQth82iDnm4kD7kdjjQjL+0r4VNDXXspwNOQjBDv8LnbQX7T37CGL4GAHL
x1SOLAHGiW9OWYm2cA3kn85Jr5Ke0M5nVp/wdHuQx68YzMt7dZ+QwpOBXv/t
XUmjdIVcqjfN32S8AD/BBX0KjbRHLFSZ9t0NJjg0C/St2hpLA3O0ldsTSVoB
+qldmovvO912sw/NtwE286UJus9C/pJStiVa873uc8h2JDtBhQpsJN6rZL4n
0nM/fofloI+m4zrsE84/XMCrDfadt4T1a5GnnNsFbs7tgErHFa2yFI4DtBot
cQnqGmEd+NKXI6edtNS6KmdFOSI0B4hjabt/+J9CFKAbX4OG9F0pMm7Q1u4A
bRlJ8xQHA9mAXOKQ2OJfgWYwRYkkVxm+Y4grUlFHWHhG5G3eNNGk/5S0WpNc
Iwq0joy2DNJMbubMwqoum37fyayKTNCLDqZZieF9uBMTuPkBcUN+wNiq9jPZ
SNu/Z4hbZFr2yKU+OvvPE7ccYv0QuADLwXqTgVjAEajil6C60JFK0j1yqZP6
BOnLH6IajPsu8gG4A+0V0mWq12WhYwDUYH93dwdENIMOCZqfz/gmugIwT5+A
VIQTLo4/al+Q2byr9MtNvfrIqpYiisSpYskJ3CB5mCGexSyq3oH+0YVn5DgS
adChJPr8ZNKlvcth07AX3ghS+AFGSqhaNBWaZa4kmSLiAtZd5izh+BCRfuZu
L4qB9jdKXYPbShJ3ZCXaT7aIeA65p7YAXEfXGiZ3EAII4JGOpDR3a1htJ0xy
K3vpmPmoZXjJhVx5bsQcpwTFLDGM8jz4Su8ThMgfW3UgIf2hgSvrUYEfPdsT
CuQHtK9L2cyGJYfmonCN+vAEpY+CXefA6FX3bxi8i459qQBe/Z/AVqgUwVg2
pVkUcnMJgktcwIdbrkfTFdp1cqQ8rNsMQVHzfcG5Nw6gICDTPC+UZkOP6eIX
bByNw2w2MBC3Bu35Ydqin6PWyUOMntSLJONC9teOQVz5WRXjC7kMupdltrkT
81t+PoKk2XrfD0kvKgsmXsPk2b1J8CC9XKHAOVXmPp8YbpuB+/zocis50R7D
iItO1fsADHGXqQbKAQ1aL5217ED+Lk6qlSJWkqcYI1d2TerqVCrf++7DDsSj
kLrB6QSHq2olk1ecEOllGxTLp7CXozLfB7+HZvlSze0Naj3l4c3w/BSCWlE7
C1gPLwdsS3t33Ko3/H+raeqRe3pMxwArzIGJ6I8Ztiz/rRrTun6FQd5+2K7Y
3gyqLao/6EvKiAxImPjUS7TzAZBmFBXqR4MN0QV3tF/ojNvP1e9KamHC/QXF
MyDAlNHPiVUnEKemBYGTL0vsJ5OJmrFxxw7wxUG1xa5KIlGaxCDDVjFDw3rb
naweG82DO3iIHcgZ0FcJLbxU4z/iZp7ZISu2bb17zkxiYF3BaXAovgFQXFYu
NPIfRvcbynJp2w7UN8pQk4I77Xg/ECNbdlNRLPUSw71E5NKRp6q7dsCPKDPx
PH7TCQV1JIAZWwxp5j5F0/Uh4V3iOHeZQSa4yV9Th6fi48wtLfRuBL6AHXST
QDmGkPTN8ZQfSaE02chDjKnzrwRo367yNJG28P+c9aF3eCMAznSC8Hsdf801
7jWoZz+gNcHkAgJjf+8Iwctt4ItR8k9WXQmWBeYLC6pXlwTu+pDjeFC+MXEd
qjC54hEbuHnISjfK85iL/unMnd/JuUBp4xfnqE2kYX+qrjWYlvObRxqyHKmY
G9C9ND3snfL4tZTCz/FgdOM2rNJ943R5LjTAQKPH6VClU5xx8f1WehYGddmY
WYt7cTIMwmnopMQsrluLqEPssk4mDlAbA2CMli+pkoPWvJxNqHtfX2lcp4kP
jjDyF15pph4i7W8jUPO4espQYtEK0FK/szrb+yMUGGc4gV7qgHrJIWive3qD
vJo3R8rJmZjjdmpwaACsNRK5NcRo5C0211i0TipOrcQHyy1AcwenTEle16jV
DhDigeL7Ohva8pbGl/SHoAreuB2qKGcwWAqFLDta7CRPDLFYyx42AbvIFAWx
l1Wd23ZExS410209Sbru/4LZj+g85eOsSBCBqfaJxHSRNNHBzw8Mpno3JZmj
+kelmIqGFrjXB0iVXvbm6GHA5SCIppSF+4uP+L6j4ihfHUu1PVWiRmGByFQc
nReyGV8B7WLkAF5ByfgR+ciL5eXCKDf9qFNdyMQksp8YkN0etqm6iXTW1Zhk
Uwv514M2s/61xvOpjl8MF4CFSuF/zK0e+3BkXd/hhNlKmkGISEEiKHvFEzp1
3c6MPWMLPZ+zs7G6H/pndFD/Rbs8rZiUuBVc6ag+LpHg91PlWllo2TO6y3jv
DdQj1KXPOyr+f2FbMgSIa/01ijwZf9AI/uE6OEO5sygQUuI////ujfd7SD+6
JqLTxwLtdleSFNxBFxtJzGxvFdh/87VWu2o/GNSDvQx1MPOJRXtfxGzUvR34
iioHICRxUc23MngzSQtIDEZdGug8N2xx68Fgj9LYM4+mk9AXF53CBFytDvcF
DK/0FUFY4ODnzk/g/stTVG1sVFxkQ+US4jQ2gvPqqKs1BS6Bjtr+u+NIEBC+
uBrS3lk/3sW9WGD5D8uLqVXufl33WdZjBx5sK/iF/o+wSwZB1J67VFnQhHEV
zwde6WjluhyiOIjKlbRcxOL89r1r1tWfs8Axh83xZcHvLqCf/FgotGsfp6B6
m2J8y9J0MphpUqc2NDAzLhEPrwBH+lIGmSuALwxGPIBSM5H5n+3xHmwbz9CE
Vcypr3dr3iIv1woZ0sQNPBhBCfV4dZx6iQbFyITe8AD7j6nVRjYqqDBriICN
uvNefOkCTTj1F9mD/73XpGc3um2bamjCwiO5c3w82OK+qLECrAQL7r7D8HMT
JAxRIavi/zfi3IoeMA+TFkeD4MqATkHe3Bf+mSlqAzvLeKZcWaXAasfU74rW
GxcB7PRFX3yQ5AesKIcdjpttbedrWk/6HsMb5RAABkWfQaM13fCkNhHfjOE3
JwtWPgRk8Lfn0X0sleJtXNub/zgS7JfC65jptwajNTs40Cuipyho7KCwz25p
Rze8BQRLK6ehX93qvIm279TD+jSL4nqQ0Rqh2qoe5Mketh/DsVbPf2yLRdfg
WIufC+I6VPlSMx+U4WPnYY4bnInX7mLuxhVCROKwyGefgiTm+RggdDx3FwFR
EgqehEMEJmUSDnWU2TD65hEAbs5g2OOG6vmUDfJTGIWQ1u4NobT/+PeEgGvq
8Pf8M+0id9YxRGte9+7VyB6+K6iusdZfiJFCpQOuSygvoiFcGoOzr/l54v1g
QbO5aXCtBjgBrdUVTefv3TtlHTlVw6FPLkbFQCQdK3pYzu50JP8TLC1iELvz
l7kOeSLinpjIPWEJ4v6h0dGDeOXqkS79lQMnJFZUDM8+suZLC/8bNd65xn5M
V4Vg5CnHc1u0ngUjdUifkWcmf9sxF4FxmU+59rqhNUNjHob0n2S5TA9t7pbS
jMr9SmUqPefvycodHhApZ2nchTWnlSEHDfncnKx5x4GwSie7gSIefsnqxjXH
vbja5eUn3tLnnTAolJ3MY34GxH2JOGL49fh/1V7lGQti1qyx35Y5AtviMHA0
AlmZJoK90HbHKx383GiOd8+X1OKCj5kcWyY5FkmBltRt4yqTVlRfhKTS2cJh
XqY8CeGJFvJRmBni6Yeaj4U6bjvTtzlR83f8REbY4C+/RHAs9hP8/GjSmBb3
E2SiEVN8u2NQzTb9jiqdZCPVvppn7fXUwlJylZEZ96/fgBdfwtBU7fedv7Wp
cfdNCDm54E8SEDfZDD1JVIYU+e2JQHJWL5nweG37g4ZGFJiH7o+VIlZT/aLW
gDmW6rpz1U9sYHM1PaOI6XpBYFFZboXtrq1fNV/Vvnf2uS4SYjKzcSuWC2TL
4Rr+Wgosfhc68E6uAtycNnV9M3J+YnXfK1HQBxKeNO69kpHR4CaEcw6kUfog
V+Iso5Ev/NxufxcnC/kp5Dm1flqNxyN+AJbQM4zP2AGZZeQ8h1uXQLTgyfJV
4/+miPP4cOlfAgk/vuk7OHLUf5FsvIisxG7ivmeXXalED7ps2QYalK9jiVya
MpNjY9WRLtMelU7ufmI1ywJZDPQd9jMwWZMJpxvPUeKTbnCc88RtBciA0qAs
nXkw/KkP7Wv9mK68AyWT+/Lb3OP8qdE1+QxUaKm7xa6abfZDLzj+mLBMMjZn
RkLLBspO7+YRQQMB2cXfWpHrI1aM2qE2LMoxQJO+A3kL/9rAXZa/p5NuGdpV
zap8iR4LIGVClcCwcDE/gliqMgBB1+nab0fkvQzlMwwNcbvqMQo1oS9ivt8D
zJJNg2rptVjHmEGYNU6aHJB3rnKGhsJm3JKlF7qAKbSLBeJUrQAer1/F+kUN
LKflNq2GynzBJWR0NNAUdN0KINGuuFUI5LtA4/wvHpqR15haeGUwjHDPF+Rc
Tlqn8AnlW4pmR5eLt7KAPNwsjgY51mSsN+m4Ftgk6jpVKJsBqkTaCjX0gf2+
7aMw3E3doMIF8SiICQ36mQht5Coqw2r0EAPSL7hCD7eVBXXed1DlbmAznVVC
jcjvb9BKptH0uRZYDAsqkozaTsDTfG/2dDpionC7KT+TY3y9kU3Co/7HjBJo
Z+6zCkyWxASzbh1T+2dca+PzOj+ILG1HjPKSRuH85FO76yeUo6kovUM3r9b6
4DHsC9CKxFx1G8dHqg9eCMtx+w8JFBx5BLJ7MLnnCKsEnGxxiCKN5xQ/ChU9
NqhB57UfxJuDTJhaVqaZr9gjGo/yNkBJCA1IVcNwvhxpEBRwVnbLnyha8Zzu
scgCLElgVI77kpXeG16kTo+5ACqoMR0gtWC0Focd8vne8dKEzRyKRP9IibuE
ceOGwzZgzYfDiWU25/zp1tmvpI9NegKDJFk490oM92JP/uDdOn0T6my3n239
Ue1V12eLPf/HHEcFSEthb/AK5iA4jAJjfv4TRfBDkg+3tUdiLmHGQ9N3lttq
8Fmo8WKLzPCyuxaYitq9s6bUgz3/zTUwdegLYa07li85tJdAoVfY3H3mIWjq
Hkr6Z++1Nc/LzIcDiQ2delRukOSvzmPnKx6mT2dCSvROBAo2rMvyBLYcgVwz
V6St+lqMoVO7zaz0Uf2haL8Fh8aoGyOnFakGKPRhKxDECPamLjWLVmxG0AAg
Tlu4hfhq+htBoHFWAyL7drm9Fk0ryXIyucwDSJmdClB9l53G2TykGorUxouk
HDOLwigjFwCbB8MZU5ZMYQhVUsZ3fcGk5DHXB0W5l8YYU3NDzlxobgpw0x2V
v2Ygz3WD54lZA+qNt/S2Z15efjoQlof2s264uDluTx9XGMsQOSJ3XIxL6Usg
DUrgkmzsARiKYKrUcIHM8hKb2dPXr+WE2sDBWjF+ldmMMsvEIOFzsBk+bhGe
HOq7lLqIAjTs0yt+vNii3q49cBkJ8fBF/ZDOJWLuGRLNhnyuwDy8SX0PqAQm
1bnSjy3/HgIbjEkxWcFClIbTYwmH3IRPbWQ0SzTnAXj7VZl8zwqBVi3cfOxE
bfhjNPC5YO/CItvxh4OPV8t6IPaqMCPq9GMl+HRnntHJ3cQiDXDJZavFvOMs
l04czG7/hxiH9+yH0VdSk1bMLBw6YwHdkdS05gohihts4dYk3KvlDeLol8Co
tTKlPvJbDeX4PPk4i76nTl7pNL+zUN9nGnRelwuSf0G9aGbla+rMdNj4y/mi
Z2u00nZRFVztIx1TXrRW737uRItbeN6TO8igVcVtAozZ/Y0FfIgcQOq39/Ld
dcC448cNvQuMMn+zRpViYj5vlPUaQSfAplsTQbJLK5SPtLKZJrf3QOy12k80
GasDAAlYkBrPoxpyMEv2tEWJLiU8bO9iRUNwvewxT3jQi3gDc3hkt8pqTbIY
xbsmSk02fEfRW1HUXDrHM+O+vRkJP3dugOM3yCWFoA1/no1sVMiHoKFfi7pC
ZlvXEkXsVYaRrCY2Nn0NCXSeYYShxPz1aQzhfcbk0T0zjoFeO289MmP8RtcD
Ixo8rdelrUShde8wEtN8u+KQFi1nsdXZrovvfbxRJIEhHSPdmj5PMSPDWA99
VMqiNDNELy3UvxeRBsxh2nkoTtMp5foN3sMw0DItHjluYMG952PHkJnUmejG
SGZQsjahlvlV7UOF6YEXwn1Pi8yoxe669uT6yGJ2xaL7OGVERs13eyF8qwQf
EMWmZ5KMDvGC+9qVo6+kEC0t5PPRYcUGwgCJs+jApQjerBJxb/lQetmXsPbA
A4373PiLhkTlptYD2WmqlWROoHGrYW0uF6RTn8cQOPvAo4mCQznm7cH95fvK
AnFuQ9u0ZckVvS8NwZ2arsGjWtb+she9IiWL150jI1ifdaOwu/brUV5ISFZM
yaAL4rAYm/8sQFQFWzwRsYWDjJehhEAz0M2fjBD8mJCNm/HbqwrdbtnZNzR/
v8CjYN8GquzqJ5K/aSqKPV3ORUWrBCY0Qo8GJMN1CLpf+E5hWelRMctyK8TM
kXY/iQiZ1oQNa9dJLd7jmV1x9zq/Gwv+f1FkXC8+zdFledfMslZEKTngEGal
3OI9cqA1YFHq0P8FtHlidvXUazeAeLlaV8uIUvQbgPw0w6rk8LBFN/jj23Bv
RQP+rf8mXPpWs5M2GYt/PV4LV5W8o8Xo8Ivk6170K5pQXV3lPl0s2li1Dq7I
B56VKK0SwyT9Tm2doL72Yvl2sL8/bE/2xefT0ih5IvIzxxeJ1m3t5HfZVllH
PYdJqcdRpW0UHxaiRO2SJUZuEcx+X+WBsxsfvsM9kOm3RBN72RaOOyIYUQGx
zOFJKxqjC1TkGSQLVgpx9TFqElgsLCBO7HAboJAdrmHSNglvxcqtTuJMeRPt
OMh+SFf3XuuXtRLBFFpt6DMcQBDRaKiyXPemOkEw6OYwCKB5lMefv8C4Xzw5
fU+AFE1zQWvpZyIApVjMm+yRB5ZiyTxTx3qyJXCAC9AJmFhWE0ManDHN5e1m
p1Wv/ddf4jUl+AVOeBT6u4JSCSSkTV+k8W2N3fO3VBF5F+C3A9yLLQBhBuoZ
zFif1O+mHYqEtRAcBjV5FhBFI0bfBcImdaqR8CbUxt0rP0QtscIJUmi8+bmp
Hni6oDfr/prJShCeEakQfibTqcCcIKznM4f4eW/27NSFA/3geUje7njizwnx
IG4KTtlhlsTLH2XKCKLJmECB792pbMxZXnMIBIooeExE1WbxxTPw5SQyMUy8
dPd4M9A35yS+D6zjuBZ+hlE+DueTjRzQgTOUmJchUhIyVPa93KQiZ84MrlLt
XouUlYVrJ+4llDmGeJk5j2SlwNBsiBcCF2psXpCOeQlfR6nhvYC6hRpallY7
cdwUvyBuRWal90/4AvUuQx7ycDFhGE2mnYMRJEkmEn2GZRgDxJer9vMNe1m+
3eCyhHW4bdVSRaW8akveF5vj+fKddOLg7ZOGNwodTKrL6S0M0YPCJR+DZ3Fp
8VpVKIfd+U3vG0aRFN3TNrQFVOamS4YTZ/PYk/5q+DZb+BxBA8PhNRW4yk7J
xt1E0FrPG/r3Kkg/zpfiOz3/2KLhlUHEBf2e46TZ7Ccfm08llg9RsVzLf/zY
u/qaRIeEywpQrWyFqmZlNUMVwMzIzZM+8bUv6FQmDg51E+JD7mFUf44eDAo3
u0Jtf2Fe9xLcV9tcuohTFyCVWUWFIZPv9XzYu91Qecc4DYhV0rp28DbZ7Ium
kP8P7IbDwZTz+0U239M7XkvM764hUSxoM/BjtK1r7MRsdFrFzRDPzlV4F1p/
phAHGO8+MDaHmPcXuidgOdm1x483oFBUSYcfXUgc5RuU1YnCBIQITLoWg1wU
VsAh4U7YBvaur2KD4NDd+u8LvaXvenP+J1ampR+rXRnzN5/6dNhrkKfRTpOM
9xUPJQc7ab9x8n8EDMKKPE4bdSlqlQLeM/9HRZbh2IIzrA1wpKG43JjYJ2AW
mBAOGcucV82KoXqw266iI1f2GDgAPTJ4TS9KcZpU+0Ja4lDIba4N1N0gHmUj
g9cd8mINF6WeTXNlKnxGxUzG4W5F2yJq/2ECJl7HCAANfjqFXhgVD8qzzzqT
LLFopppnWm314oH8NFiI+dnPvPrANSC/Ab6boEongVCkw8UkLm/ZTNB2SqFB
OXXL0+LNzX0aRBrBDQTQNwAFjRYbO8kJcqRVc9eovhmWwqJAm6BOCX12waa/
zENL+oVLyv/2is3MwYFc6HuTDEoMepXeqceK85EzJgi1pARvY2vNAXGM1nvU
FOQ4aXAZUL3DqKVaYywlnC9LtcfrRHUCUcKoEfqjl77hSk5EWSdufeAQYv0l
eXIFLq2YQ0/7VGWKpyeRmWxaT+4OYzvHj+O79M83L3vyZodDk0k4eVe8m2ct
uNw0RLIskmPgwLB3qux75fvb3c9zE7IusGtJG96BzfM0LbrAkYS/71uVXie0
2OZp1xae7vGv+G1QbxcPKa262jbAGCtYQlxaYUrfqoKSDSoAcqTJUqPbd3k6
zan11JzLWOiqWBKQbFyMT51qdjudVc91VlFwuQk8dTJopNhy9pWDheENBHpS
Lsbu99LNnSFG2VdnOOjc/hzTD1HZohEVCXY0suoBrKZU8Rc/f1h6TYF8qE6y
i4JZTorkXholvYmtA8kljPckriON4DWaoNp3l3Yjy88y8SRex39at3NhI6dG
b97sdRPXcYJZhkSBMp75DAFFaRUrDv5w8Paef0DlsfycEVb7Ft6yGHLp2qVE
Aik+GHXcxuJWZCNuUwLwbrvXRzq/qEOudtgWw7fDYpvzIXe4B/kAIoznqtEs
5l/UmozE5B3jqgjrtmzu7mU89xOaNgLuRJ7uQSaCvSgmN8RT2bEEAYvKTm0p
REYcasfncrji/vzg/rwYS/d43vJUPxdggS5JQLueZb3erA7xkXFUQoxYjNCp
9BbGCOQY791k4oRzL/1vlz3WtLQ3eE8WcrPkWzoPNLsUXNPDuV0kkFrl0Tbc
w1BAu4EipDgKQciZacftjXRsArs8Jw5RPeAu7yODftUa1i1ndjrI70RHAyWG
VZ+dY6paWcMm5sHxq+m8wnEGoZkj+YhpR/w6m6uTDyYrFfJxFQso7BIwnzwP
b3+spnjm0+lr6JnkPVH5JluVkGGRJ3InCbtXvDp6lxLrYcVsKvamGL2VZKxF
wB8ZBIgBaLiR51qjosefvNpr2MNICIfg/WInIxO++k8PPO+tcGsJttSYUWDy
Ouu0NL+hFF1+VRY3QN/pzunFjKryxABn71XG58gyoref/E2gIgbkUCGOB9Pn
hc+v4XSoz2zo1IcRPYNWq5Q3+WDaNHxemtC/p2+3X6kjo7yGYym+iHr7g24v
FSnBjYlCAC94v/1n0XReGO4eJ5Kb3bBs8aN2cd4CvuQBTJYp2QXzxUiEepiF
UZlB+texEOMnsk8lyoFkiloqHUomRmc5aAW+Myqy81O3YM66tJeJLRQK9LXN
sTHfsGZW8AcHHph67HkZGuHNylBpRBG7wDAyFrjozp0gIy85ArrAZC2bmsgC
c/tyiliwVWkXvF03G4wS/gQ7r4voyuHEkTTKTRdqpN1uP7/FkOJJlERZiXdY
0lWQA0GMSe9ToYyNz7QJP6MQli86e0vbJPh5nL8RrYNqDnxL0au3hTh62ITq
oNAzTDyVSEEwnjlOAzUVzuu/0TKNe+ehnWu4OTKBP8PrKTNQZNam86O5Rzzv
CY+2x2uGOwJ4rT5G8ux1Vnvi90gEe3zivoy00ev6oAHFHyaq52aQvDYVBM1s
xKodMLPZxYnRPRJ2xT9pRAPOiaRlpTNij9FcGJFCb/bAe0Tik/O5r7qtT2yY
BTtDT6S+iFzzrWz3dfBDRDi06A1Qzd1OQLwQh15K9MjN6O1i13lngP8oocHF
qcBWOlo6BCYF+34ldwOHY2srks23EEApmajkVjpQ3+qX2j5jBh+RvOiq+PDm
j5QpKJ0FCCMi22SdxWZ8+aJ+a2hsbw3J1x9FcC546UHhnvVsfKfEXi5y4oCY
cJYXE+7Oz+whWLZv/0DVIXb4Gnt0EgmUKGo9Hen8ADBYQnzbeXV5iatlAGIP
+VzRihxLK6YjrSUzxTYxkgW59BsNiELmV8i4EIciDY09Cxthv7lEb7R8Ysez
rVrPBUZKjTV0wenmQnO5Um5OAgA5BsZfblaW3AKz4QmtWIhNVFYVcgvggNNl
PeCVgaq5XxenTbn1A6p2Q8bxaXjXq5gFuQxzFwIMP3PBMQd43A2TEEySgFhV
LKSkekxVfG3gukKnHtegKqgCoAq1oibLjNgksfzdco0A0xtfvHd59dcnUWQP
tuIzZ7M+oES4u7CEF22qA7e0p4fzdWwLcCBvAlTgf/uyXSnLxoCaF+g8ancB
RWabVCAhhwD8cAILOYI2XBoyUzUmSwp892iabq9t4zVxHar1SvjPuXxCSBQs
kTsGNDub+Tx6jkKEUUx8OxF0UBwh9TpLY5eIQbBym7NitUnDyV+oo62oE5Mo
DPPiIsveG6Oxo5UXWlRwTEqzN875SqbKUz9FMjGlpaNrtB9Pzb1+Chg2sjOa
daq8ls1Z4MZGbw25Hnx06Y0XtsPvRi/geETgE3MigdgJF1xr2POCp7qVGdxj
nK72GezqeeK3QMYoXMo9xxgW+/HZ1j+thqP0zuX6L5ae/WcZroJsr4nMTpqy
CcQJMWsNyTRhnPJVdABZtXHZG5o5AiaatmdZAttNZm5ckxGbTqKqQuFyrJn2
uJjAmt6UVrhXT1IhCFLAqpNugRZt1/TRss20v3MNnm7wn2px0SnBJn+5JJ4D
pFRWk+D5z21IcMXerYxFm/33Q1w4FXZ2RPNGMzX8NjbsK7y1xDpapGMd7jAa
UoAXX3EKYYw7dQGtFBtjcUubrh3sC16YfLpeTQbZWdgrNakD1vihiqBDfrj2
GZOWj1a1EnfzV9N9VseWSX4xhz6UEwMGN3TbEuOlnMz/zoNuL+DYYGAZ7j0V
b8QWOUvWwPjTN1BH9I2IK+WGv1OdyeD6ha4g1ON1KLjwa783RD1kR0phFV4s
QL5YkPju6BqKKmZT59KJox62erZa1E+GANqNATYQvz2A1flrOyLmGwQpEZ9R
2ePs4b8hMMFv5wjaZWJVdTyn9wP2knEmqaa4iYvqEoctAkhoIVXAq4XPyfbu
YCOB973Moj2v3LHXy+dHO9JDzVTchbamYObeEwvsP8YRmGokK15bada1I2BH
17fGS57KAdUBU7h8IOksNOsY4i9agBQFIkT6VM50j7yu27T+5V4jO2/yOIiJ
VmeGCtQ94OPHfQU+Na5anuGe1fhny6uMuCn0AvLul00EQiYUsG9d/nXqypgJ
iD+xphdcpFnIafaTY6h+RtumPurcMExyNsay9V4d9zL/K8ICeobX5r8ZP+3G
JQHyRaLtVFqWK6AVJSpTMeXSfG+dGmbXSwMv2j9YT9OQ+5pfoZ2sVhWLRu95
jYIXo5wwrzjko4ByJKVVhaisAUfxWtUTwWO/GXgK2GZy3ixMHRPzgqhVY1dI
1EnamqYJl5KR1ujDzhL6ZTBGFVa4gQwBAo/7OF90pDlSgj51QrTv04+vXdHG
oVmVKvAgA4QssRiLMMPDWUFgcJtZAvaIXF6+jyB7PlCgP12cJktOMqAouaQQ
dq0sf8a1l0b42UlCYV/uGaiUkHcwg71P819DFEbZiHn+v8THdKTCkQOLuojp
17JtR/rGcix+w162akJtRNczpFZcPh6KCiUPv+98Tbig2xZ59pUxhyyW6FmE
NWh8xjd7HomSrxShPG/CCbQsa+mEvbXsuE/OmarnvNd7NEn61KBUMKM6nvC7
gJGixom9BfRwDXjNSqVhcZyxSu+27KbbYBxFR1o1QEb6g2oH1gjAM4tutk+R
a+yI++w6z3ObzGmbYgNZYTLQ/b+lfIgOlIVqjOyavcSS4ms75AJA/wOKhDtm
AOZI/lKuNvEBrpHigXSj4DH2ChBqlN36tJHni1bCtPkW/JfodaFJWBtZJZXa
0qHsZfAa+pFbuqRbtdm0Y225WCBymniySCpiPWuR81/1Fhbt1JiTCeNDhXEu
FX9WqrUd1E8W1dFRC/1aRKH2VwPP/iroirZS7flXDTxBpKNyFLfD21fdw1Bd
xJY1EohcNxRei3j6WbCglM2fUc7VCE981Tt9CIXKS4jNcoxYuWoCqmHXkyK6
YluYQluQnGn9W6iwlE6fEMqfd1WLKIt0/I1ph8e7eI0C+5Az94Y5GyqXEjlN
M0naM0YWkBErBuP+yqABhpsLz5WjLwsgj+RZxEDaulClDyTGyAIl9/Kd0NHH
B+GaTAynFj/VeLeXBBM3G70QjviZbFamLahXsSp4cy+pJyvawPgahhcHw6Qa
ke4+ELTKcTyzoN+PY88dnWKJ56eiB6uqCVGWislHngxixPymmzTts+jpDz5s
j0eVXxfhlbN1UCNLrkJTa7T5kg4SuEUgmhivS3PEU4xMpeB0jJezHXptZ+3b
GzgIHiGdaJtUV+pPTGX96kHB9PAPDKvLSFsu/CT7IeucE2o5qh/PfI0CXiqc
Mc0JFsZzn2UwDO5iSNCkpU6nr8j5aqN6ZwYCpbbWNRgyZcIwwanTJEZnK9e4
W/fD3giildLB9deJNWyQ+fu5Cyj4nOMoOMbqHEBrPXINg13lkWZolYC3JSi6
DhEF4XM9OebWBbz9V4No6K2ad9dUy711BgHFQ8dQerbWJ3e3K5Vwia45dNzH
dBlQr/g+A3LyHXEYMXQ6DMNaOtqEyytAHrQDd4MxVRJhTPe6Il9Fgrs5Ur3Q
uMDNwSMTy5lzLol7uxERQFMXvIdNn5bqXHglSS4yvzOwqpwYERIindDMFBFq
+Y7yM6SnWeGpJKY6uoTlEVoYk4MLBXSCDPrxXsAwNnBgoe7OzdV4gejyAbYi
RFwGCU3kJDWF6UsprOnm4uOBfG31t+ia2mSUSBiJUzKjp9fpTTXPzc/AUEOc
F70P8ab+CphfmxvZyPb/IjwS/bCXzHhnzqayEf9aUWpM0d/DpzsJuzQ5H2LW
Pt1urgzg4aixVZRNVnOC9wC0Aw9goFaf8whvn+BlgQfrLacyF6fR7PRr7q5V
S5qUtMbffU+cL6hfFwUGWIADSajodQc+GqYu7O8awen+Z8FQhxLJYDCXFByq
aqgEORNZsIvdKrpcC2aWN7Il0MsWV6+4A1xND6v77P/nu3rbuZzyqZ2MH4Jx
TeMjBKyxVsq/6N6yv49Tez+9xUvl3gCdKrUWmMqx4fB1JFl6P+VHboYT/TEu
kbAS2MiDKzB9FLPsi7M1RCDYsDhEp1/vxgFG44AD0E+B861mxQytgcu+pqoI
aYKzVMOEj6/6HssCx+5VDKE/LAwO/wuON/5aasKdggfe4v5FPrQuu39dWjXO
4Sq/SJUtQDNa1ZMSr2tfiJhXKSQ12k/1j/WSPmc738iqPMmmkLGUgfDfPIWC
oplhKveC62+A/kofjy0Je5BLNykSC46k1DlN4rvKVLT3Q2YgJCb5l2n7hhIW
BYKkpbOBNB7w1/VJu2pHtxjm65urYs6+6GUVj8BuP7kiv1h7DpBwnQp8ARBs
fFTzgE8RnbtqsWZGW/FlmNWIJcPdFNdGEaUAYmMqclKbY2P5opjJ/y/KSTgg
BbRIN0eaehfE8VwogPjm3k9ga1DURaRO3Q12yQdbjwj0rzfiGxBc0BzN1tRs
WFncmkxZaBzpr7V6UCbg3g/qVUJLnMpkwde0bSmcI22tbgy6rEJwgdKGKUc4
97121UR45Tlic6fVXwAGCIdkjnmd9OB6FcGD3KN6+xs081sU1umIr2Iw7z3Q
0voz6EzbFIOifzXqK4/RmfdajJCXzhrrr2uJIzZZgvXCncc1WOJO7gP+PcMS
TIe6Kgb/ii7UUuq57q/mVZi8AaG7mTDomlUcmvP2EDjXeJFbyxs5pOE4Zkzd
6NX6MnTuZRgntTryP8Vd1/YNmjrsAKHkc3n3Nwwr5O7PjyrgJX1GF06Kkp3F
gdZXamrcj0egVbStkdnRrY35Jq0Rwrli+TnRfhtKp5I5EMAFVvhUD1HlAiGd
ANmoFDpxqJtNaqCpGy9DZKEGiZpoKYeTVqtW/01CmCsl3FDlUBEyNUtogs+w
2eO+KQ4v1GDNtzaa52c39XvAUrtYUM/UD46EEWPn6wjhvH9VsyjaCQzi7cdj
Pl2THuvo9h9HdzeSSRPXsk8554Qa9+aSjFKB+mYIsoErl09lLFeDjTQ8OE3/
3BD38Yx7FsAvG1HDqr+S4QFMosa8MDEVxeG3SAiC1UYWDAZC0KI8e8RNOXN8
kLbKd0k7dEEmiQhWnGhvUHHN8Zz7TBILpxATqH43+i8AvnHXeZqzrtqna5ct
ShRY90hjmDxu6oHIjwHhISCQeIzked2rxoS9Bk+M2bqAx47ApIVw0K6Qz20e
tJ8YJ3DbsA2bxAGHWpRBfTgi5Cv/aGfvYJAmlGPax5sQQ7N/tb1bDdbYDiuy
OBc6HeV0rP1a8SpcceHZdAWQIz2WXstCrZxqDbN6yFW9YbvCQF0U7KTPKcDv
fpvP3mt6MUUv+rdPMc84PiKZl7Qr9ziDpzR5uoO4r2+RanxqgAGDxcN4BUj8
P4vwEYfLA/nCz1yJcR3sBa0SFoYUbxv2rhI3uUKpAT+5ldgYGGoXhfeLhIHj
TkGb2sGDWaIZ4k+QZ9diNzFNzQka9IWkidZaDZCCVEvZWXWIom11Y3cj0mQt
F7CtDnwCFx4XgkTdSAshwNt2nBg1oiR6nSSaqFY93+Yeuh4jQutYTTHu7fbX
4pA5io9bKcG4aF7cD2wCVQQFIu5C6ECxBt2rqyAXlZ8sECIH/oPuR9iVPgEc
nqZdTaNnBGHrB6YKYbXGLyhqktQnwuNMvoFuwpkqwRUIgXEnUfVZaqGfqnUA
EBWTN7UJGoTb4EAHOL7aOgD/TmMP4Au9PAROLh09neLf5cEMFOjMF19sQFcQ
vbtZY+2GgEGc3g7v/N+OEXzSiX1vH9nl3376Tt1EUI8+NFA5y3PFnDWRw9Xb
TUkIiruc1DPrZXyexYi0nFpaFa42LYdPrp+/qRf3t0zNqGxD2RmXYb7cj7MD
xYgGkULotYPAbLNC4z3n0ksD0crrznbERBnoMUDVnUihblv315kDCZvkycvK
T85KFXAuoz5RnoEBN5UNrQjjL+JX84Xl1jjBzkp9s9sti1cW+qrC7A2eWcer
y9lGTf/awBehTUOfF45Ba4UB9HcBuQeFWLuYXS/QcjVYOHHjscOP91VAHRCy
Oko1ZxNZA3JkXSmPYnkVmEEBVYIgQ7jSw5ZkdWCdsEZnMwQHow2jzwA5mOcT
8btkWmDiRVWZS6NOEV7cvd6TrrgQa0908TGKk18X/4hWK8dUhOW6kW5T7Qtd
7v1LPq7JhgbDOQd3K9JEtYHWNZR1LqmXrEkd6hrOXZ4W7zsfdvhSLF3iU73j
U6TvXG3tS8L2N+pPMfXYYB88REzR7z2OTOR/a17HOehUw00O0rZbKpcU6wyR
uUjt6uVt8QSQal2yHgqFQCsn+mZCTCWFnR0TXqTyihSAuTvEN+8JpYcHs+ya
IxOxCb0C3mfaf2kZgm27QGBZalba7/ZE5IbHtbBpOS29qUQgECsSbZWUDpMQ
WbKF2y1IDh/BHMwOwO7YDZO77GVLIeW3wfY01jGeJqErBdzsNjTbM2Ww8O39
T0TY59epaB7fj9XcOEanQkKmxhySm0ApqpFJ+4Xm4Q3FYMtVRfuYpMJbQSCk
nTptzLT7Dnz2cmhYoeZiCaF01im3+VlKagwCp4P14gdge5axGdiaMLwnCFUZ
7tMWLkYLSMy2PbFOKa48aa7Wff3JETRC/gQantRhMaIKv/y9toil8KwGdXPr
xanyOSAY8iBnX1SBCxVDYsLUMQcrLgmLtaDMBBleNwYxS9btaDbLhCHN76lF
bJDaVdDJ18t6AwpUu67FCBMcRpuCFcqtynoyoO04b0pFq6UZxUM1AB4gOhLv
kXurfPvDiS2oiHrQ+mO6Nfg5tRc4sU+Bu1RTBfgbzzRKVli2hv/NLoW7O29G
i1LZmghGSPf7VoyZhulZaEQADhELRDze/a/tZwNNushrvsvrwYQw46T1C51V
1zCX/HOCU4OqzLI+xsIbANRqPsvgJjL3cCIEwc1h4109JhoHprXgTm4wmimu
iZGG8iEcBLBQk749rhCquE/y6o7FyNOpI026tf4Afu8+DxKDyCfLvDdTz1h9
GipbiqqwKR+wMEuw+T476+oUifv+GbxIe2BpuA/mTVUZWwe20IUqUMkVuOg7
+FsV4PEx6FgAq4B5NFddFGTHh7nJAS0jWZbPlR0Nc9OGgLn36FAgX/Uaz+1t
5iK0XwppH3wWbNJYlV3cL73Lahn5vmJeoiul21mxcgppcpFUZLd+68N6s5Pm
1KXRsQXPdhHGp4oqsZsOaGok+zS80tDsBlI1wakjLxlN0rrlmkFVSGxf/HUI
XPq6EQ73g5K52JKjtbIgceno0tJnVhkDTtY+QW85XBGpaRmZ9a2tl+aaLodW
moEbkvGc4u7HTwdHib/SQ5TZKIvaiACcDU0pzQwrDzVX6KF9MZUuctFd92jT
mxOQIEYSGSlZmSKk75s+zauUQKBHEhBpIG8avnYJkAu71T1aAlCyb5KSxngx
fluX7+0hdP46IWWa2JloJ8G5Who4Ai/+dNoJeYTEP/tGaFMGZj8HSqD0/jxv
Dh4mRE0cIDKy+QHI3Ig6N1dZErX4nWypn/KqeUX5C9qqKFOIkU7znEXyS4oH
0DCUdDPGLTabk7Ydc0qU5rv9eRGJExkY3tnFLkBqYDM7ku/eup1hQPIqObBd
I1Wl8h6ov46Dxvh4gNKEqhfJYKIj2gR6bFARkbvTtbU/yYq7iQr/HfcX4WL+
OAkaaPFidKflA+JKnqgIBrHlH6jN1LzPUF87Ebnk5XrwrN2JPRjFIBquNt2S
vbKc3KtknN/ezk9JNNbTKjgaHK6JwZTecv0hrhjVjzIFl6MwU8Z2tfnm3Ayi
BRrhx/dnPaLzpzAx65hgVhJ2HRE8QaHhJkLkHth/m8GbNzBOIaRMWQABr1J9
Y3ILU7vJBCIJUS/bbE6eJr6pStXdc/jIq0NpmQYCC1Dk9e48tpaLRLYKvX+P
NLVcUCdu/6xJvRoRtSD9nSohnGyZD7McmCXk49NAjVhTjwekb3DW8OAGI/nI
5LvKua3fMPhS9CFej665ZfUNsokV92Tl5w2iQlufwumxqqPT+MOCOChRaVGh
D9r5+pQCeS6Q/flaAkzcKuNJg7Mm369rumFUyEbNu4FMK5/KGnMDlGx8Wa6p
oi85fyrvUOOVmCCCzD4G3fTNtHQE3a+d7ZUHPzPyTXBERS8jOvxjrGJ/b+qu
kE1NWZKUxQ7/+bSHjmUZdTrlw/OvstBjoft9zJuLm8rnH8PsRpWEHDOfpR4+
HyXyZu8xa8fSCt/S9QmvORyvc3n79xy1KqwduJpJw46JcvcQeDe3zwnKZtLI
+aI9vw/1hKJT7ANIOUBU85VDYP7jpUzr40YpJrHuR/Iz381MVxtXZjxcWUuK
McNlMyLLtlns+Sss6o1GqPr4KDe4rWS8mBi69vVJ2hgF2mFpNLlGZPW4qdM4
RMK4UofE7BX3wUfBVngOlVKjoFnCFQeS49E29Tky9x6JyAZuE4ukcYzOY+kk
Kqql6UjFMOZTx6iB/DuZmOGoRxaEVjZskIW4VfsIlgdPDocJY9wlG2AxO5fV
rUuE0pocW4LybBILrCGGMtBqw2zdhMaaUN8Qx/fcpZ71XPmw5gb+nu7UzGqu
LUqVdWeQ1pYmkfPl75/g9YjC8yWPiYCLkNMYaAid3Pf1AGBVnkyqZCliR0vE
cxJ/51vQHL4dZpBgW6Qnu+bTvVwkiHZ0GzVOmKWLHlywXYgZVzgOlUMEDgtW
mVa4jfu+oVr34XUcw+409Km2QxDRz7Oee5THwZzdRguWPV0LWPRDSZto2Yzh
C3yErUrbMdf69zZJLu7KrCv3G+d5qD0n0XPf/Y4iF1fBJsNALRjvkVLWlc5/
DLJEkdVuPchckcCk5Wpmd1V96UqR9hNqtA4CEcDas8qqXEjroVuEMC08VUdY
P7SC0MWqToSrCJs1ywW2v7WveR5fQZjSNyAe2vWp+jhlLdvz2ZG09pf4a1dd
fEUr/ohUByDuWtYUt7xz6jXAyVFqZYvmciGjclqs+g3v/tBg+i4q2c9CyH/q
3WGyzkMk1QMU4NBuNumaNOc2uBr4VOQNaTSuDFvcQpubqVwcH++1NPHcngCB
6EaaFMGIKyD2ozgTMq5s76DDogNeJCH1dtILX8BwB4eyPrO9NvsiFiwjnXuC
+CCCt8TuMxewrBOPoWDCFPV942dWtCbz9IqPg/h0S3BnQhqrJ6BK+7asChfu
mKKMzs60qEoDF3d2zl/3Wg7edmZ6YIfJFCn4MgJhOMwTvHVUtSRwvoOG80Zz
gEkN/QgOAYFLgjJK6xntgBJzxzSmPFoEFNYu5pn9DKXz2zwB8q0FWy9Ws3rj
0P8FGZpQvWQ67DoVRzUoYZQbFEG6fDXgoKEmFQvVv15kl8iHX24QtEbFezbk
fkWNB6HX9eRrEZ+CIPHv2Pz0CpRNBfoFSobJvMN2GEkW/IFSkjB/TC0YF82l
J5AqWHrvSfmrCg6RFrJ855Nff4q+mDvLG27jfhxLBh5trWkLtEiKM49Ui/z/
Hk2x1oMaTa582L5su3cCV3iw+p5X7arCnhf0CaPAZpqCWTncxP6hBI1U4r1O
7pejlN5eFulP7MWTSPUy466k9Rs0bmLbZb8JytZOYzu7lgkQ3FAKN7t7Hu9k
cltWUDfppTiDHDNGc/qh4g1S9rpcu7UOE4UKfdfH0vu9nfMXZ7nbF1nA0nte
UCzfnE6CkIHh2C4KNz550fTsNLaooKHUibGt1cTbakOITlAta+/NvFxnXP3s
npXwXAaU8/6MoqxbIiCLtw91Gf8TnXiThU3Yc7FSIkqBqyik0BKZ5tVugXUV
+QenltR8aCxYeDn6/2rAWIm0yPmMTdsCoeLzjooxgTrudN2o1eZXZGiofaCV
unJDNvTQJqOIsN7/MARtirvyH8q85QxiijSGWDYBmAj0HwOhLSedWm/UgvGM
tm+jm6j+X+bpMeP6F/RyPE9uIoSi+7hXXDlCgDHc4yqlbrngC6clCUI7nyQt
sAIT0kF4tyQypq2Peqchr1f1p4DfQsRXxViXnSDcGhlPbkCpQsTZhr9KC0jL
bZtHppONvOyX+hZPxAWbGR9ls8fn0/YIrrV474yzV2EQs7edPafnH2T3oU8f
9zVQy9RTPrTcsXW9bKQWLL+A3GphN8fRF5xawEcJvJopguAYalx9nXMUl6By
twCMb+k8b+MCHyun46sD+Xid8E6ilKi0mIOe07aephJlnsjRg5/NL2/8q5mM
lJd8Yr+/7dZt68mbyRX9RU9gZNxCYyswNVSoqqloQ09xZNfZFun12JJOlsV6
d7qPwJxZy1lBoo5cnctmPlEAG9tAi6UFgUoxtX38oormO0X89vLt7b4tICZY
2Dd53C0c6BtQkms8Dd1nY9pKBi/RlNSzc9vGud88fTmxYUEYK1CGqAMjU9NH
w+0rPOWQBZhzmotBiu6vSHK1VvVTuinWrv7OisniY1E7qvyv1/UofvlNq1w5
/v7aTCE1s83ugQr28I4PFaFv4UQVc6bDGKiKO7mAy86ZbD5KxUaN5Jd3OJ5v
Uu2fR4yoh8P9Id6FR414xBlFHb3N32dEVR9ZRUGyms+3z2HbcD7m6IO/gTIJ
1WO/nIssPr+xMeI0ykjNKxdoT4wa19H/CTWU7lewpuD7aCT5ufGwXkB2WZUU
OoQcba52hjsaojI8j6ifglz/C4hlPLuuAuLgbl5XfLMNDgvw4HqYRH0vZ/+Q
qZJp/4fv7FciCt1ijhfJZbvCWnpaI+VzW+d6Zmm9voXSwGPapgtQZDGTQUm1
jc+ujdlb+ZFzHRDMytYcj9f7SaLzDyInFyMhAzlPMbW1agx1OFdBiTg4eSLs
sevzqOzsmP9VOEWD3XiK/EWQ0I//YyeVseWGPVx1YvBnJXbrJJMg8SaBnHPt
3sSOMjknj92J1kbNV+6pDq5ohRj3/bWncJg7BGDgICNoH8ZlIHRU4JqXuphc
mXGL7kQQYT31QYSrdMAM8VlpmV8vXtcCLZBuZnN5NiOfYo/FxBEvFIYAEXkA
AnWg8EFlHfK/xjF8EFSKNqBokR3yztYHLWHOCfVLtCchcTVb1JvDybzI9Biq
03tWR/zVHyFAl0Unb4diKiO21tcnUdacCpcd2I+eYuzLIf+LEXpcevCvKO9r
KVX5FcYQZZ25u2ew7A38hW0MGgbY+R2EHTxJ6dNwW7kLjYvBv04xktzjtcxZ
rqC5qwifWbNg7GhyTBXVM3CrqmRpbl/xRxWEDGibpM1Com/qFOfgorBYpoqx
FG1rgSjv9PigbHq0RJ/tFLN5BBkNKOX1tA66Ks4XoUS9gOWB5DC/VTyMiWIG
EwRw2mNNJ3CaE30NEQZF5xCwytKTtgY6NzRjWIiitHwY8nWBqf3InoRd1xU7
Aof6gqgAWyB5VIkJljnyomt4J73oXmv9U8Zm8KCdm6CZoUcQRfE53Pg9VctE
DKxiDJ6TQ9hhxuMzL2w2DHy55VPa5dQH3Jq1uta/c6J9qcihz7i6eP7bqE6b
SuvwiSF2PTlU6yUZ+NCFYiqD+sOxlT+DOQ0IbjLMCjdvw3E2ES/VCGnvAF/N
WTGXQz3e8SMVXiXV2K5xGiJu/U9wT1nbjLTOGrLVCpfvVINcZoehBK/uYBtc
rwYXkl0tABaXgTc329qW7UL7fSYQmcqLsG6aoRLBG+/8cgOoMoMtm9xYVIWH
/fm/cxUP/cZGAcvBeX/n1HBxyaDgop6i71dc3fjLNWlL32F9fpmU9QgJM2ce
Nf2NHqWMCyZ+tW+5E+19h4By1GdM+Axu1JaMwV/xryCzD6ylvMbS/UjYugSB
fRM8TFtGUnPADp/HMGzZmLUBJi26bq17ofUei4Riuk4fnp2605mwtxEjIPuo
L7Yfu4emYInkkFFW1AQQnE99FiRsfaY7SRsSdLFPUVu2zfAgYonmkAsOhz6g
kG8f5a7xuRCqmtKCSBmh6DKbXQP3kETZZ/lhKJDc9q1owy5KQGWsG3KGlKd+
cP8qg4psxTUzLHIHsi6fJ5I1g6GigDNcAwPNU+2a8rs3yfI7zRjFM2DbbqJV
w9iHYRssfSBDBFp9oW6p7F47G6zX10LME/SYiZ/H0/0cWDOOWk31ZqnSrm1v
I2ZqPuaxiJycWzYKlFwykUQiQ5O1RdfnBXt37PHtQMzfhdr/wFNzkLdnB8MM
i9+iZ1njQkIqk/x2R4CBNQjpP7TXHIjExpErm/BEavHs9ZGI2Wyrnmp0bWzy
14U/LbHouTeGeOaU46Wv5Z/sF4UnNgvm+cyPPviVW2J2YrC2vfVHlgvjpqyd
FeRqWyuzphREGG+IZ4nD3Y3gxmZSXDbgD0UJ2QF1bNbyF+65jQVZnRg3l4jy
lyOa4x9qbnsMYVl9c1V++Gaid0+bY3BhR6s9aEwKaasZZbwmEI2DhMg1z2xi
PgcUirzZjY6P8nvj3CmvZL3kjZ1ploQNj1birvMuPx0yyjSzpgDbb3LM//PA
TUpDXwqV50p+T6yUkx72EJGl63Ytt+2aUCXr08OpOSGT0A7mUSEn49PWM8u1
uUXEJaKQxLEIMqdlJS0/VHmPLhK9NJq5bJf48tCAvxxgzvsnFUbkG4KTggpO
/yZV8a25KNHMBr6uzA4OprwQfNJxt3VTIaBoYrJ7mJoqUjtHlRrC7bL50FaE
oWERgdwO4v4OFsKsy0nhRYjr1eQzHVljM0k7ImzZvOUUxtm0m5t3ZkWwz6wx
j9PXxF0RoylRXNiyhEf4sypSbNE/eAJANdQ9goqKIpYDS7Aa64b/iaRhp6Rp
9kMfAMZxoqWyGOTbq9CukeM6Oe9o2wOKaPdZzXNHUhdmOm4xInPSLzJo9SQS
d4Cfrs3iqBqtrJaR51FtvEYsAxU1fjpOEzRpyOOawoPNk4cRSJjOAaOFj0Ai
JB9DQ8p7O7OcO5JiiHKIYmUvhqivhPdhFWfyZ4/bPp3cZhcr4LpUAYJxExTu
0my5I8kixG3jjilaHVTK71nW/kD00vZ+I1IyWMWmOqE46zBIvszGlcIqPDap
ZR3tDYA/ZklQ3r3L02P+8QxxRHmub28pOQpTaL87MoYJXN5AA3Vge/yxhUiu
XSZqoq1mQOS1QlAlMHa0EVRuzN+a7S1EpYX2V5YzzRMLVXd2GHzoTupg6KBJ
AWMddbwM3GcoPwg3WTilx7WToLdgPZjqI/q81grsRX2z+RBlz6CqgtykL8WJ
4UJKQ734hdq+0Jy77g22qVyBjIwXrd0weATTQzZRMsMndm1ioLX2tHpumueI
kZpK2YgDpohwj4F6NZfhxuuLZl49j5aBZVROrT1VaVs1xpsPqe8dqT3wqCnj
DJ8AZpT0LLLVJKHynaWaG6PzyZ8sIrb+S+4xkcC1dX57SNozU7Gyym2Ez+S9
CJde8SHFaoAr82wSQnVUMK/cjoiz/9TCH7Q0I4ttuslQxUGTiWFmmnPRUxLL
RSFDl0pcpvoObdzMxQQ+U0QQwQLUijpLHeNxRr6JvhecnUY7i8uW+7M4EgeP
oDn1awNLDcDwRHrfW5Qb5P6eyc+1gIPhYUfMF6Fc77344nQfhGhxaRktEQZp
5LBTj6P4q6pu+zXEViYQWt5cQ3W30BsUJ9KPWX6edNBT03jk6uDm5s7FfGcI
uJ/1c4S5N65dYwoLxpTw1DZYSW9ufFMxhpri7TsksIOl8wN6ie/wEorZBWia
YlLmh8fWkPFpzO8lf3ToliuaAebfOLtkszTYPD+mnk9hUHxpN9+wnC45cu3N
uel6J6kHWLQzPYJKkFcjmPuk2oqujXx64izKRQQm5azu+st984hsmDL4/+Gm
f8Nyoqt8VZMVYFQqtDrAahHEc+Ve3IfeuTCgoGHKOu30TCdtvH1IWf0b8FtH
TAgn7Y/Oi6EdmyyyTP7xSDlSijMAm3fnDYpSSFERXCip+HWAmWYswBwVgwY2
rQuf3nQ07Awff4un7jm2K6uhFgSt4Bm2suhjXbYHb88g+9QATVgGg4yW7xdP
Kg+QAvP/f7kRcB9JvYsD3G6Yf6zLbQs2h31GiZy+r4IWaIkFC7arU1lAiiys
YbQ/JOUJUMVW9TKiH9AyiaJCKDPfELxmUKNsogPawqYDRYuEghBpOzNenYjo
pmoKRiUp0x9otzK4SoFsO9NfDdsYPIJZwoYPYqlr+5C0L7UbJ+LKJ49ARD3j
ysnbjvGJIhodlOygqXEUU4LVtbrRFGMSresqkVF4gDPDFhKEMpf6yiCOL+Zq
3NIY5XomyqfWzu6ycsb20nu6d0RBI/pE/GN2Nq8qM0lLHDcUv8/SyVdLL0mQ
29Mo0eqLHg2Mq4gKP7ld2VaR2yNbwtuoPxiOuADhHHxHGNzz9qiMXAOMBuvr
Vz08s0KUvyBH0JrW2b9KtaDDPqwkIzJYXFOLWfX4opvLWuDPli8MsZfmrGBx
yono+ynUEXhAsQkkWfKoHzlt5bkdGTIaGSToYHMOgIUVWTp1GWqsPlHMDyxK
nz71CkfwkZ9tAdj9i+y+lPCgVgDgp9VBN8LnUO6UlJx/Wz/kC799X76cckG+
E4YwAqs56zvI8K/7bi0UBGn1GByOZJfgZtmcMsUtfiO0dFHpITOEyJA8auUM
IqXS4lqoURwSxTQmH0Oy0+MEVue9LnLYtvvr9xoio+2hwwxGVAAUkFnPQptz
gjBmfcRUJDXe6oIcFytimLjExvBiEreBFqoPiVtI2KoVY72zZbUKq52K1UWT
1l4pCstzDf0t5eSbJKQXRCKzUVUf3K2/fxySFCo6ZXENfwafYeL890OOcaov
uz7BioINRWmAa5GODbElSl4S4C4lNKpn45pLulQ1aea/TjkmaTY2ucPRjTdV
5ZLIMLdmTeDb1Vpo8pE/BaHLt4IpUdDzX7NGCEgSStTm/2n2+0sQ9MOXArv8
4VjeLXX6so5UDqo9UW1SnIY+PTH8NvPWaFajRvV0Q4qWkjoNiZf4qx6HcvbF
MQQTCshU4kKAObtqbk3UuLTlm1lPpHykL+zRa/uN/gR05DLgeVbvIfABkEdX
zciyoTIIAeflUTP2+ltnwkFPulUMYR9SRD6m0VN+bwkZVJTgNqcNv6Diuabh
GmfM9wOU9+FFpQDgHMXezF4p0kXwGP0I2jsj+ye23eWumscfiCrNvyHH3F3J
z0aW6Pc9wPw3XtmzeFx4ZC9F+ACQzSu2SiZ7+o4aVb8Pfa9ebUkvbRmrTMib
Pi62ggYHHKHt7ClmOeXRQtDpu4T9nucZ4X9AbNK2zlL/7txIgfgA3E7czGRa
r7aZUmj2B++UY3XrRjRZernaKeGfTc7h5jWhNRWBb6lsxZMs+c/GsLqIACp2
W4rbJ/EuU/ElnIXH7JqNnhB0sVTSRmp5sFtWHwruGfG24Jet92VjEyGmFqhz
sCCFXi5weqcwI7tGNhe1b5bLhQRgqKqmCqNA8VbRkYyKsKlirHmzdmT6hTBf
gotjk5TzoxKRuR4CP4Y+S1g9XvCZw+BJXgUE6FCX86TrWbLZQwRz6maFhZvy
XwT3EGHXBTbowFwbJRpQn0u3phhfZxjZQcQLxccJfxaQVDt/gtPC6DMvN5Au
ELSKXTvcKh9W0cHJH2fVuQz3Q2UHVlQTkfvWoAlgK2rDOX1ipEtqFJaBhS03
4UjA9tpVpI94qtvdwV9afN4WFqewMMhMDhj6z7IqKR2K0IY/IkFNAzW0w1pp
k49TDtuwGwqX0u8Gbly2a7PAmxqvhwdvNfKumYRkBi5ZN1AKheQwRuaS2mq4
pMq4k1ftWm1nmLknGpTvYxIciuUcUqyCCf2rNjj5Bcnt+5OLRP7WRk8zynyv
IcaDc1MZMwseJ9QNbLVDOOs27+nU2JSTBojuVyhAEBbxYPBBvNZL8cWU/v7J
UzpKUc6JVRBHS5movde1vZsarwUV7cTT6u9kFc3blcqWpqQJBjNKJh0EBK94
hHIkOOhSCbtPev6Da4vULpnRPC4uQKAywnBh+g3msiYDWAEHgrHeAg2/6NSn
/PK+VbKkZ3jcdHDV9i2lx1szaij+iqwRRa2zrfB3LuKyEeIj8e6Mp4M0Z7w9
RgROHnswdafoYijFvqMmAKqBP2BIfNoXL182TmdlKbvfPviiFrJNlc3BE2xt
c2HcljuG5+bNAByEsQZ3XXyMPxjIUDRUUjw/RsCmkhuP8W4mQjz344jkfiGb
zvHWNjwTQ4JR2+Kny4ReERhfRn9QZTnNdGvOgDmcdEGpWarh2AeueXiezR7N
+0+T9zhG0+EShpWW3hc/9og5RdGxS4zmhZpIQj5xPKhPlE0u8qbHfOL7weNP
MYaUGfL60wDqVkgAZDMP6N3NzXciUD29XR38mZWnOI3QIALXpE7HehFiM6P4
afqBl1PpwE0fiyM/qOohkvBt94ct758l6FXYU36cFbSzHcugq/zxCBGQHsrH
juTfNcv2FL7mb00gGspYfAEh2Hi13hda9dsmXzJX6wLmyKgQK8W7UiBhhE1o
MG5t9W8R9OCs4pKBuP4rFU4T7UvR114vLJm2QfW2PMAzeI4VEiyKFkcw40WR
7H/cn5ORhYRzbYisW682wJWEXXJwI4q06LhkAVfTgH/7U1PJ06CJ+a9snVPt
G06y5b2MLoyVSAEQGVcOJ5xe+aRtqzl6Df4xx7fVTmLigcXpXq31wW3Ju7y6
LTfCRcmA73oNIxnDIu3+mTej94saXhvr6SLkeyKSwVKOpDPauMEl/V0MePkp
Glbz8ccVBwwjYF3xMPtNjMg0F9mUVh/H6gwR8cPzBGUM5G6fy/PntsTn3xBR
+GlgeS7GIOSnU9aywiPgGQIs9y7Mc8kOOZkyiVAvqrdZvq56UsGcPfZDOj/t
6p8T1bisoVRelQYTJ8eQX8ylljOtKc2L75LR2GOiUHJmBAg8WKF1j9ezpISk
rilhld0ICJ7puNLG1VLfkcdhB71vRr5owvmp4fJU3Q7aDZz9tfHJOBWhH/kG
44LQvDubS0y/UKNJM104pBptm7N7l9r8FmkwRo9YqF+WDU+TkkNyZvdu/8qd
XJ6Q8u54qINa8o/33CeXCdBiXnTQn5BXxdBLzayvX8Cni+4o2G4cJh30digR
ANJaP72IIEIW/+TFq9Xv/3WGNNFeNMv+PTpe/rsMHU89110tnlh3eFqIuUnX
fr5N/7GQ04ZrhFkHKW2Qppulf+Kg/XoUiFhWzhy61MkI8p+gcHhavMKXNGcE
0Kx5/U+i1DqnrrCR3XEGHsgtfWrUvIjwkV3DH3fQ3WcH+maR9sMdGiKl1Ifd
PlDHgD9NIEmHWQHE6+xsMpXKN44kPVSjnnHCcvPkwLaVMWWyMw1modTDGtb6
dePwO62qZZ33Ibm7C8bVdxZk6yQxou53S5Qoy6IGYch6K0CO/I6Hc7xj9L7W
0HfysKnq7rpH4RwRPEvmTPmEV3iLC/W3sHDE80wI8kCjUu/zs7wQin8KkLvl
VLddY3SAjn529+NXbLGjH8n+gmt2mZWN0KtMYafEjnIMmIH5qXgXfwP6ImZi
gbmyy0o/w586hwxIG4CATOyHvOfDp2EvCGChUvKLPQjd4COmtEyoo14h3yiV
HtRMMX7qhq6uP6p+rk93yVptekA9r5jITyaBMzJsWjzuAiwpVDIAz/5MAs27
h5PiyBzmj+ZhecEj2zu+xvnojqversp34WW0+yleETG6WiiIk7UQ2x7M68vL
Lov2/J5mfC3MgRQSv/VwDm7Os7hRGPaxc3BFYYRVpZYbIm/JEsfFR430q3kt
yWD6yhT6oO661VwoakxRx16tEKoFEUGIs5F439xQbSFIs0MB1WVYQQGOUb0+
JCYCjUzP8S4X20dQnKu/LsDLrqrg6P1QKHmRiZtC1iet5o2n6j7pUcu/HX33
DX901tM0TopZpsGR+axi53wBQFgTM+QqMGlLx2pC9MDEaWuDrhLoIhCnPEk+
ET2f7nVVkyXmpr+1Zq7Zi0RiC97pgP72mKSQozJO0x8EyQ1yHLCWf3CPyMHy
Ea0RpvK48PFeStP/ieKhaHLfvGWimR2Pdb7aBfFZElOyeqSWTurMR44upass
jrfRRm44H8Vw7Qsazul1+X9GDtP0Y7PEWwOxTpJ73DiBGCo1WHR1rFaoaG52
IETuK1wdKjL7d4NgdUL+n0Er+5R/+3mPqJhjlukeA8DSOlVaTD7Rli6X3UVd
tH37DbMM4qfCjR34ReIdeZMRvt1npgdRJVwpTkO9xcSqqoEPUsIKjfVHIaJ2
p1KibEKM1n9PiDPawLPzYBhQaj0qfSO6BCYm/fScCe1FuHWncHbJsz900Hxq
5//nIbXSrinhaT7rKTZawMylpOdv3L20e6Rl/jX9hg19nKpH3MmxAOlhtj8I
IcElHNTfW2ss+1boel0qHx/fiL08MRHSZKSVrXyV1dl1CivVeCopVWEKyBNQ
w/RrS1HVH3KslNY+DbSxlDLXxgqOljbFme4wlIqDRaRTBnjZMj7GJmzYCHjw
CG0rZCvny+Jpe9aq/krmzp1j0CBq3qEt1S+WxXjC6Fzx+CeTiFK4U/kIi+o5
C2ND/WYSuSwPp0COn7hXAe0Z0ZEMZ1weq1j9diohXim89tnGTXP3fwzlZLQt
yrYRRwKtT8V7tjhL3bkAMreQxga6dZdzddaQSIrZOcBmrVX4GhEN1vZNEtus
nVVwD3wKAgwZ2D1Sm05KMwXzKC3R66bgdAnIcJv/F0Z9wS9EZtLr82Sp1C6N
kfw6v1gEvVQzLEn7vOOBIYEggZbrngxfTJ37ABU5XgzCn0tL6Hjt3Kkkidot
jIGpCNt9TGugadv17hiNF0U12fXT46Yi0Ux3c+46Tu4U8Vi5ThDXx9zoLoJo
6QF9exMqYlKBoecTNE35XZw2ndT8tcJjNg1pn62myepAPqkZWYj6QbE6EhEV
ZrpRRK2Uc1t3uyblsgF7PWhJegWtqq6fu2bbMeBAJzQGf4yYtNxQhi40AABt
VHcDxPU5Nsr6x/ckp1VxyRFGE3ZeiUjbLnNo/KAVN9Y0+qvSMmtK5D6KVvyH
CqNWJCy6IQw8jWQ7a3auXmT+Lx4mkluNcbsTQ8lxN/FeClgJYteMFZj5O/Lo
4PXqwqQzUQuxZnOIhK6iBXrTnQtYuEq7OpzAHuoccz78gryfmOQzRpbqRKK+
eytmSB99j6/OQQYh8xmMl7uBwBAhFMSnP6VZ3sddWVC3Vc0q04Bl512k0Snw
mMzZVnDXYorgcy/JbqQdacs7OjxoODB+dGhV0JpQyYYMUwzHWjPlrsfoAl36
7mmuYclu3lVmTHn7MZVmrf7+HAso1TIr/in2Y64zALxoRE8t1m1WHvSQCkGA
kuWYleOnPs6Ufdswr40UaxeOUIulXh3Rb7YzA3TyIIFYut1V1D8AN7mzMSqb
pzCqnDaxp0BKl8xRri79dxERdZe6t03KFTJMfvzzTgr4dKeGu6dquJY7yE3k
vfdl8S/0uu/AR/00D1v6daEqcvlCECqS909lAbdHM/OF7VML/i7kgpkYsWrw
ib5bcDSN4/5aX5ET8i7rnGzkANm2LyWj0Ycrwhooo3F4xXacJbusLvE1E1Db
avNTHAVJNnx5uWHX7nMhf++X2InjK0W3A+aPqAzPzeOKIrnwgE8xdRVfi45h
hMjRhCyo4yOEdnD5f359+i24sn5ZxTAnjv1xkYfSPKa1pmUC3Dw9j92/YFYc
hYA7Ou9f9e0HWy8PrvvnN2t7WAADnX9CtrjN4EkqZVMgeAkX+T7srRbNkT8v
iNn9z3QRHMlfwhpXKCtG3VDHeAhYgsRH+XQHMmiwNNkMBi78DA/a98CuHQ4e
kfyWodWBr8QTKYWarcu7KZNYzKjYlBvUl/qEeuw+rziF09JKgPsATLqWk8Lq
YjFnDTOh4zIMvpcn/zRkZFy/NpZYcBFwmGc+TQH2GCJ2p0J56vEiFBLh+s5D
gagBG11FQdMipd7Z7mc+6/7QaYKuW8+z2Is7CC3JyT0cldfIgsjv2erEymb9
Q3ugGTaLazfUjoSOe5I9qJFQf8t5EdG3Nq7TZCbUMKiZZUSX0SAdVaheZxn6
ieBEIcDveE8qY1zdbVkZI6skADzD+vAHCbei3uXn/ArhnJsQeSNORj4Cwbu6
ZPBgUN1EKLRZ3Y3gcT6hGvB/3zNXa0sGkIX3UIKCPKHYL8wrWLVvjCtgOIh9
IUiklIrO7YPg/6LemhoMA+CI+tX1bMjShJ57RjrvV2nmxPQ7U0NZeopqdqfu
1v8CGxEBZt//dbQeHMVGqF+G2M6Hy27+5Ot2voS4/C6HWJ6gnC0xpN3GlgZG
hAfcbfCyz+MsnqJH4mKCrz8QecT4XfAxlIUPED+vzxuzk9B7oFz3GD+BiSEP
KZkXETqqOfFeZUi0FE52eSHYPGwZ0IYzwvzASt+2mMrajvijE6dNDYt2m+fH
In8CSYRMCEULpKD1ocl8rDx31iXGEdePfpe1reYh4seaDwyOKD9RMEhmmbnW
9RvoIxs8/RBuml9vI6oK3L0MzjaBfj27CRCrmEx5Zteei5fDnbKFOBxZRjeU
RuLI0CNHgA8+mcdIfaSUtUWms/D/6xCXaQufQG/mvP/jEz4I8fQxxVlXSsV2
JLL9b6XU1KC7YLSVB9p9A5XUtytbSS6RBizYWmOzMlCkStsekdNfZmUY1CYn
+d8hRzbP9Vls3VM1/lOdmTEREMseTAoOU+I3UpdhYUpG5wXQnwo7lag8OEBs
Kulg+q75JLEsW1GgKx9fsElpjV5Y5IAITuDjBHaAlD1TRgj8OfeDr21hRMT9
aY/8r86l8KBkdW7+gotS1H21QfvmTZDAd7zvh/2YytnwSJ9Y9KpCyjJDGAbH
im+raYpn0R8I/RF8khcNqrtsGwHKGs52vc8ambNGIu5UeuxftipkMjzh/bsj
Sx3uKiM9qoVoEMPtTpj+70oASRVoCiuAzQTXkzNwEwBg7EUqsZSnBPp4nNFP
L1Gmqgq0mTmvpHf+Cv2DGuicQusWVrgBpRlPpUuiWGVhjJfhR2SNUUJ4QWfJ
TCj9uyocNRy4HVWLuFLqpCVkU09D7Fnfq8maHKg+8DbXDtZOVDsmvJmOvK1Z
Swloj7RZWbthaAW/GfVKShBbDY5rpVWbv4xaOpoNto+aoNNd4tQUcxBhr4D0
PyV/E5e+jyza/jBS9WBtpE10N6zPdqStPmbcW2HPwaJEW9zWQI5Hhf7J3QZo
+QSUbRfccm7yv0wcUWJYE+VJqSdN3L9A8ILxfNjhwbQcSNkMrxJfCYk8WvGO
aXgP2hbPkUu7o4LWJ/ULTfbsfKlyk9c2TK52k1xivFdt91RBtTwbKaF8b6LN
yfgzxYrrDE7AqvJFIjvtt5rw/z2sL3jFrQNo22EoTOe61rdjqEeKbrUyMY0C
ioE1WEa3UbqpzWP9ON7uncHwkgNBHdl5LYFc4gPdO9OulylMc4AHFzqp15Iu
RyxDC4znle8utmX9W8RYo/JKLg21wEAu3deQSpv1sOkdPdwlH3RKxMPOpjjw
dhLfkDaWo7x1J/F92/uVMJlhApf7D6r34K3zi0IdfZIvHqf1D73XTYZ9TZxk
OeKE0YIA+Hk/4hCyO+7nHQctriU6VHZiYNYW0mO9DkQEx/o/AhyJVcVdAGKh
HCKHr8aJ6JkmmWJ1f7dMSXOXFMcUKg6Vfck0u4P3xmhP3lfhSS3/hLrgHj9X
ssz5AvNkNMFMZAP9ZQKLRe02h1rFfd/wNGdhLo5Wg/lTGGJEgZ2jWVsjTrBQ
avTJURz1uNMNSiru6DsJ1L1Ia21S87euN6TpQYBwgDQSiItWjn0UzNLkfz0Q
lJaBb5r0a39dplBUvBTGcKXUFvt5CYbC0d+v8EJ1lQcowUaHL1/KIpaOs/4f
8MZHSPfkfJRY40s2awygBM5CCkNvuAGCtwUs4vKBTYoGxIjH87xkvjnkD+qw
dhM8hsbkpc91FESFH8EDhlas8JhTz1JkQwfuO6Yrtc5cQam4wl15AbM0rgW6
fXJ/QdI4j5j16oUFGX0USR31xqxnHXeWLc7Hkmql7n9dXnWK71BDir0LIxcI
UoCHHyoJkmFAs4f32PzI0/vCBZHA2aqu6YcEwxntuAEK2txfklEABdqoxKSM
UrPkzp7KDCTnh7L6loT95NGCTux/ap27oYSm4gzZmLPNWbjvsF4EE0UxvZei
Ic0cvCazSTkYF6W9Jl2n77UyxCvvvbdIcNd0SoVFTuhbBIwxQYnNPmyJW24a
Qof/Orv90ewKvVJ8oAX4OJiSpc5XvgO+TVgKLxcJ6DDbhVZ+zFlsuXBW0lTt
CRrJn08wGA34qPEz2kfhFHNQmyNWx5nnJQc8lsR0u9+zqZqeHAsYWEXtsm26
brFE5U2dVyQrY+oL8D7NN1xYX/AFjKAtymwPuF6CTzfZyET22f2d17qmE7GD
nYfSe7mAlqnGj0DHR0V0t1yx39wN50/gOW9adaM7mQROxgQ9/XPfdXmAoO3r
09YLcTS0nfR0duKRUXxo8cfli522JU+30iHcNdK6VkQup4j9seJ1n9ubE6K+
xOBYw23IHpBrbJ7pVRrfPR+PPXGRFsSw2gzck5NDt91Ci3gZjzat1SWp/Buk
lRX2blLrVIJNp+02F96MiDESCLwtdI3GjPc2lzLi642KjE29GPzv0K9+EKrz
9PckGfWT3WLdQwP6ycMed87jIMkr7ac6XWmu0Oy1iI1vti3R3hKDjxrx6Mwi
gCkcfiYNPmcbrttCFvuwGzgxdEo2Areyd66m75zZ2HzPtlL/UX2DL4KQdjzb
gDBYj+nt0mDoXWLlCaK2yrbHoffOyWHzQmaMM3vWrFX5CGFJw+cxecQHUZrR
ZLZ9X7D6gxHfSDc40+RCaFK9x7QUE92gvcsMipxHPnQucZKo9UxMY/w+WepS
QRuu+sdV9J8rPHOaH34XkYnnJsF5+OLEoQLBgmKzDTKv0QHk2TfewfywYruQ
NkvzSoaQOWdBjMy+Y1Hm4Df6uoDJT498cH+MROQQYpXeMK11c+4dnbKolX6Y
+teoH3jLKHpyiJ3F80Yswh4gD3U2/wSJl5cimXEX1QIx6auveqOtn3J4M/Jc
tSfdjxwherLZHD3XfKinU14/FRlMtg5wGzXMl/YxSU5ufCRWn+XVkI4THuZq
hwoVYTSSOqO5HMxardd/d4n1hg0BBSD/frihB3HJlkj9z2V+/2FDuOrHrmD4
iWUHPfjnJ1QUwNp4sQUKXEfeZ5SM2mtNmLQ/ZTzvOrsZpKKwvpKYRx/0twZ7
N15ja6q3P7DFRtJmK+EpL0KYfILJ8tnGV0JXn2h5Jd535hdzNqO4RO3t/2Pu
sKcf7aTLeiJddulQU2+G3UANGNPvY0nQgmrpro4EnaisvloKq5zsklzS9jFG
Wspwkp5ug2K8dfCfSDpEDHjrQji1vh7IN5j0ei38JAeM/Fcvo5A/fc74eyA+
Ed3/Mu1yTP1xG9DPdPpCLoKe3NfJjSuv04ZDNe3f84pB+r1b4cUrPagMHmxW
A2yvXtAcELtfGxK8fTfRIbOanbUh/A0DOm60YfC8ggZaLqpf1mFfKoj2CSgw
LSRK8OOvUw6lHNAec0O5a64ZGA1GEwNs3xtxZOuGBtp2oA37pMlARjT8XQWJ
ukszkwGjx6lyR2dafbs+bXblcfzSBw30c5WpHa43ss7HZ5ceJ6BuDhAlbxQ4
eUoLJR3sMaBjonKG8ruezsJNN5MAzRqs+BfRr2JpndHpODO6fJHglyXyUlFX
piuuc++LhnuiXuKckK1ADSwAN3c+6WQeE9acYFWrGTXZtvKq/kjKhtZ04wyo
WVyO4IKi7FbK+tp7mIZzr0dW+Vw/6NujB7VoR1aNrN/4Ax+6nePjiGbHD78l
+VCMpVyf+lQPlKJvqT0QLkDjo4Qv6oI3l9o0AJxDvbSKz3iLijjmw11kGRhs
fDFs65iODg5vlo3LSLtNmZDJOxyu18FDTqjAcqu5dCKh18aL5UmypqDPHZVo
7SkmavZ77aKCw1EbKsytA0Cu6IsdRk6EtzxQqXyPyw8obKgc23Ipj2G7zh4j
jcLUrbjvSzG6wGf/f4slYrLnlR1l/7UnOikk0Tbj+7hRmD/6X0M6/BmiTxNR
VA8b1Jr/8qqFA6qbccrSFSykcCVJQnTyJVrJhK3TJ267gNGjIH0ABP/Yjq4i
3ZtY20kSgUluYe5qO4VwrQoQLvQBV4GZOwhQ8B38csOW/0YALHNJw5pVQDHg
Ydd15IKH9TsvDzx9iMr19nNWYommWabzY1qjkm3v+8jEto35666gKBlKHRtA
DRCiIlA1b7E6kKm40j4y/TJnLvCT0gsp3/Kx8gzK7yFv+L1ruaFVWRTswbwr
udpmlolIOCh3RgpdzIrBRt8fd4fHna0xm+lDaCutRXJet3j79iSavu86+yo/
QTjcvuPSeQ7gJ6yzjc2cDZ3Xzy23NfujonRMCBn3RLNCX9B0mA1KsrUqHG7l
9demsJfNk94V3QTvuQfJ5qbkobWzycjCsR6mpvTLcD9vLkm5/MFbQCY9+QXH
QGW5b862UGsCOCMznQexD/LnfvSvdNzKb81BP4tN1y0S4Gl8haAd/dHn4Nx2
RBs7hZxBP3CJD+TV02KKdUfr2dXwistC1OnLb415HycwtYtC2pBQwgF217GL
NLdi1rANgdwxmH8bsb1preI8trjEu/Ri897V+QtrxIi4obVN/XFoUTtRctT1
2n4720DyVq6r30XSRfK6y8V0YHicL8RM4PzlyAcFId+VmRJy5KG7qkSedh67
uWGfd/LeoSp085Vvo3Wfh/BKiz9dJfEI8pQygKUyDwn7XdXZnIpZaGGXN66d
ED2c9BSX8F8UVQh24Ve2aa1VU5ql2gDWkZcrJ009INdGqL4QNKbZkhECiBhv
Q5rjqA3jM19APMEg4CBc82JRRbF3WKaA2FxTuMXR7dnBh4Vk/4g3ZDq5ErbY
yiYNOflV3BVmth6qmDzLHuuzc2cEBCj7fy+fMhw9H4TrH9J5FUby1hgUuwxV
Y9wHhRP/6ieiFUvmYiQo4zs8Ytu7E0BkXkl+fMAypbLkRKGqqs0T4X87i8dC
Hbh8TiauxFfA2nk/YlnJf6m9QrcqQG++tLdM6wEBWJD97IJhHTMSPZZ0Ajt7
QBbcbLor+0twl5OZVHRbItYoDIZUNOK7XDQx3U60DFPwYI6eCoLLTF6PEVNS
crPfCX8wP1990CZh3655cRciC8CpNil/tvewLofk3BUoNCsUqMy9cq+brf1S
qvyz0jcuFxu16ohWHeJ0Buv2Ewqu4knID8NT3ewsBRt/5s0mjOrdKNbUpyFf
0RKLlJUfFdfr721gTlTXHEU4GJwLgT85V1mr2bQoktzsuMduK7AzegbH2mmX
7qvGTHhxASojOOWNE80W/iuql6MPeoGl4cWRG8Q/YZ9R5fRLSFNV6A3xo8/D
oMVNVCiMeW5DtBUEvDBifj72TallrmHEvAVXLpZLtjo9unpSED0OIkOFZL/G
w6ooPN88Y3tHB6aq8CTrlDqrehMSqC6QKMa14Wrv4Thlx4sAEhmEQMzn96AP
TQ6dR6dhg4aHeJYpIh2xzgkFZIF7v8XLu041u43IeEhik0qWCVWLdpzeRxWD
MxlKXFSaGN1aPoWgMmRVbAnemPDxTwqicdmyNwXkDjt2hUViUga2sGy6BXtQ
+PxRsdTg6hJ1/GFyY3TjVfqchYpbkkffuvQkUcIZ7BbLsji0C2+UVMWjQYYZ
nJRuQqg2Pyfz7FrqJkrIwgRLbEtAHzzOy4eGPhZ1eb5PplTOcY1qOxzQGIOT
FkqYE0EVFb0jadNtwwzxxn8mFZAyvwbIzez0GAX72nNcZxuZBWcT2dKkdXRj
hdR6YMMcWz8oYNZiiyPZjgQzVa5NEfCpmoqtPjDk5PA1nELXyUuxie/xvi42
v8WoKLTbYOTqvEw9PFZOh4ALFAnMcjeXB/8NWYTo4AQnOO96TvJCeDC/JQSB
GCdI1Oib98aL+afHRtfCI1abvcuX6SV0IoRKYNOjjBbtMrBK+8e+5UVJ1RT9
AYGxUaL8vShEFS2t5V/eT155AtZDMIoYe3BP8l+AmuScYozUl5+j1XDnfk3p
aeZU3hnLMd9qYMaU15hEXPPUoMv6AKaAlgqapCuh2+UoG8A1CgKruhd16cqZ
DU9zlqCLw+OSzfcrhje4enlPk3bNglVMa9sOcEV15zoaf7dtSRfSkoVau0Q2
Ulz/dMzYNfCkt53Nso8ohpN/Bg/oLSHinItSOMOqCViEq+PpwAYJiJYwffEH
1UjPqsfEq/woGZQLWCC2kg82WITCoeI/W7VoGKnlQaOYW81g0Crk84xMuWZ+
fyebsmIsHpf0FO/GQeaNwx9NRNKNBMUcnmk5Niw2Qe+342WSy2ZszQqcz+F6
i+mG8Np67FWKf4kE8ggH7CznfXPGKknhHd+7jErjd30IIT/vd6I19hnhjXHX
lgaFnLt8mhAP/vwAR9N6KHP5CSmXnKG28jP7yKTsc7ktTC7u/V6wvu87DtU8
XCsUGV33917bJ0MFA5C3tyfjhVW4jyZ1TlOOUVT6dxsjBk5l+kpE0NCJpHBn
506ws/o9h939tgMjSwjNfbfQuyTND4HvIzB9WVZBpPk5tBVip4nwF4rZd5Er
jVMCNhl+zKWkafZNyNyTeGS00F/zf/4GfyxGvcoEobgtMbniymOe9D9rLjvQ
7ElisiY0pj+YpFkDJhOxDr+M6+X7RlLY6dB7mTG7fc1ukZyWavTA4z5Jhoi3
YtDGRznzQZgyHvyanNNwhpVSYKg4Dwa9rllDe3/WKQt9Ql82ed8XPVnaesr+
xzYcDtpE/dPzMvgx1CfKLTk6KeWshbanSJ8j00QhW+gsW1sM/MbEBEsiRidm
XeBwRm8lpH9T02dmulySb+8lw9j/KC6heyXqJKNdQz/FD1otaaRsceHY1AtB
zD777czU1Ti7Wl31USq224Pbhp0NEBaEf9t7jPxL2PIA2bYovoe90pbQ8vs4
QuF8Kl/KFJ/dHv/tMEucK342yAbN5dzAmgHNQFxjJ0ABCcZ4V0N5Fmtd5NKR
6s2iv3Vn0QtjcgdOghXzJXDvz5UFhLnLQIIaUryl3ShstmQJGo0h1/F1j2M5
px8A2QtoQk6vXDrG3hcnwOYdna+wIv23HlPQXDF4JCHh9IjtLkvgLDDHYwpu
D0+XGban28cCYZJSeVJJ1kbmPcZ8jjB4r50w2EUHg40dWsuc6nmaUpc/Wm8p
5yDQoST6Uu+MuR/b2dchUGI0A5rbVm3QWuLr1qtpvigVWb/D05B6TuR8Z7kO
8bEB+fhGXADvH63eWfbzqleZflLH+b34wpanamuXh8iy9HaMvW6Hiiuj16XQ
sC3eEr6yZ+GTciYe1HZgI3otb0/fr64w8IXwIJJ6pkvbuE/lyNOo2UAVX/Tq
H7sKsTJpiB77qwWT/qdaPL9BnrXCiPfCWFmm+q9Z3wXFh6oex5zWmunvTfe1
gyYESLYVOw1iccoEjYUl4pCq4Fqw8JSy3ZnU1Jbr3utFkuJZzOzS5PGKYKCw
GfsLmqxRFHTLPfJDaoRJSY9bIZ2UR719vlD4zeq7GoAX/13xnw4MTLsiOFJ1
XbvOqC2D96I+Phpk+DHVYQb53cqSR9h05q6egvooSCXWZL1ypm1rsDWUFWxD
K0YUz201UKwgm4q6aDYfCof8mquosM8jDwUEpuPVmtj44lO5xTkdgt5R9kai
ah80+pu4sMZp7reeXzANyuzYY/XgMQcgkp3nkBmHICqLf4up8gbH2p7KUV89
+aheu2J8Uxvyl0TnGvukH9rhNJzDHUEtFR2hYDm65avJNbH19IXEkqJ9irgl
GbUDTUygIGdJ97e+J0F9NMcys7WNWpYSra9aXQjlvgd90cUxr7X7tOS14s+a
A13/DMpWY7+cDIbUn9MEiTzmvsI9kGZVKY+Xo+1WgaItXivAoN51xvxhnba8
pa+r1KTSp2xSPh1wax7qwBBJ0cg/nTTEgp3WFEL8MYlt8UJS4FCWR3n9ivyq
YZ6Ds9MB8AqTL+d2sQgce8v9NRVI4BZPnHgpKGYRZUG+KlvO1iWQqUlMyBsy
s6SC0apnksOcVuVUTR+f6fK4aSEMPWiD0i6wN1l9vC3kXBgIAls3IEKTpWjp
FSPL8M/6bbS7C8a0gnjpEsij/tWhacmkLdpX4f9BZ4T7p88vqnMSwmddXr7e
CkEOrmGMBd+bzaj3JlYqruiqDeOc/KS+tMJ7eD387eeqOo2Rf3hJBzSLdzRw
W4VgS+M5hYFvuLgSYd2Nxgbk14KqQAKi+kQHnmQgYOmXAejHaPKg+NYDbVcK
Ux2FmqtKFUn9j6G6r6WsdfXpga2lGfkRUBOV6zwXeQDbrzCUTHjjPgRc7KR8
oBvOmfWfD2iTpCZw4SVFedBKlWZvRGepxjo2qxmXKyYmpTbbDPN/XjenJMpw
cYEdQHqZ0rrav2/pPfwvf9ZQ3o9mD7jlHkPxFh+lszESkomKSRlo45WOacdn
wLU5JUG7S9WOz59xRiqOIAIwwFZPs1L8AXuBnW4xfZkkmnqzEAMtrMdudEyf
F2ml5+r6618ESbWfvwCGFRpFPGDP3zkfAJW9y+fMuVupZxehnR4L98nOsP0S
nTkbmV/fVGJ0l7deN6ZDUH9PNsreFcvCLPMnazBEjMTExrMSjN8+MAjUSPJy
bdOqr8nZQpBctDUAKTYaLo7VYQDmu+3kiKigOpeFPF5cCzPNOLu8AS63Vezp
iBoHeXuAJHt6R+2L2BHST4eb1rqAUKzE8koY1CVhgBGfr831Tm+y+h1McGpt
uFhH+Dz61YsjKg+mEWVIsPPXdWMioAV0bE55Xp3CziVrVAgEy0Trj8YOjYcL
9uSYjq78iRUlBK+7lcgiPBs7Mm70j4VTEoh+Ytrt18BmFHJIjvhWuAydzyFS
Y8Nx4u0FKJeVqzvv9O/bbni4a4/bLgLI7KhRZJ/wZP0hk38cKYuyh/cg3xxc
tzs5nKxkH3gbx8rnqrx6UDq+v2Pekp1yvy4NOrh7cruOqysgc9AvVWVDSkL8
jAerBc31nm0jUgZchjmBC0ib9YjjDA9O9yufABi1EC9lMDP+kTOujL8dFCsT
GpjQzFX6HIa026WUbS4nHz9uKGnhIpXRIgSUXdQPAGUZHtmgYkPoUGPEjNT+
UxCbkXpdBXPrTebdKqiM6VgPlckR70joSEFq2DY5lgPevYW9Pg4vIOYd8oAs
MO76nGoVyzWHSUZJVCGBAFp1dzoj2dTQGEPTceMo0e9rf9YCXfYJi1UyQY+1
LzcrWmJZmdv4YSVkfv9JLhasFBGVb+amLY/mii/zWfyXShKq78S6pwb4YaV+
raGmQzb9SF17MSX57oG4tLzlFdY4oT3dv5J+koTYwzTfwBLP8X8rfBn9l/NX
Oye8X9iQb4jUtqkysiFuqrbVC2rovZX046tm5q5Ff/hxzlxfEyz6p8J5H+Pw
y7UKw1rqD3nfQTllh3gfh2S1HVvfePM6RSmi6vLooSvvBgyBHp7szR+7bblA
Lx+F+9K1raXvx0Ih+oJvBrWdi4RyRFdkllOINBTXEN9XObde+hdHOX7T5D3q
ZbBqE0d1iMyUEOXmC2uCtZ88l1aOijb4kpKEEFj9zeZ/NKTltiSfj56qSK5L
iTCIxcFdkC4Ki/QIaI2ZDcuIF36P4ndEc+Q8fwao4KFrdfe3IypLcF4Gti9n
7L0x9l65us5YcpskN7iSl7p8eroFHAr9u64HqTiVvs9duxW/AAspRdJmparI
WbYrLhKwGf4GCjtGlKKvhnAG5NqVUqFIYaVNp1vgejLBUKPV6vtIJEphn5L4
pc3GfWEJOwJ8jQHHe2ftR9nHgE5A+mWzp20koqswZN/QgQO4JLBmZY3lKdLi
e/a9eiO7STJ9+uIAaI5EBvmQs36U372wZi6j8+2EZm+hS7CWutoz73e+vjpf
s7kvXNTrFoaiQkHl6V5BjLo6JxH6QCfN5srats/20fccHnIZsvDM18fwqlyi
Gh5DFzxZDGlyDY/eS0TMe7+W6EPv4wpknjCpf2O8FH4wDV0tXutnkA6N3AEa
3ewdpvDbrnNgw1oFRFx4HeYcm8Jj8D2zPUfc7NCKKj6N3Q0XGPoRdpqAgE8x
0ZFBaUXe059N/G0eWtqmuSRUw2/3sQJivV9FilOZ/wlKujvvK3PpwCDSxh2w
vwAne3WNNoaPuyLYrOhGmjvHrSCCsggh2xK9sYfbIahoaTP3++sgAd3l4udr
JXXJictoJCDjWI6fRnsx/FO+7zkPjVPtREaTdlbl8fGlvwhAihXzBmVHfXo+
bY34ScXFwLSPs1GVIPVpRQx7jSYxCYOSQvTj2+JsowlcDiwHInoYZf/2H1OQ
bP9bpjIKZVnRqJ41IRm/QbZY5QCdt8jRWhnwtB2KFOKx7//hdDYyARNOessy
91HMWLZfkfRgLv/gMNv9uGNMdah/dXJctWffZp4qBP/Lic3dJ/8YgRbRxrDM
ZYU/GaY2sRA2LMO/bopw5oBkGQwrsIfp2OTr9DbZBXFjqS+YOvZ317HZr1/r
WznJjXzXIhHZp+HVZ3yq2brQykNWseLivGby4TFNWCPPDSwXugyioNBwXwcL
kFBONqmz513v4pIC6d8EIXV6ZiFH8RuANVLdK/Y26893LZFPgvdm3ivcvS3k
D65dFVQ8EbeuOUAs7NwP0Np9Ew4YUvgD7k/3XAAqR9Ou/VFPOxm4zZDhKwye
MFzPx+zZqBpcEJ2QXwG9Pm5ChqviD4ejSsI3KhT6IVJVJuPta7HXI5zRbOBk
GGFJCNXBQ+AKrN0oggCIIK2YdVngLJP0rfqbnwWH9LmXYowNZBVlbGmi7FiZ
gyEvuXSkpdqz6OvkPSafqQBaT14vXCR0tV78SmqAmIT/DUIxkvNL/V/RZuHH
qLddHe9GFQLXcm8SMNBQN7i5aJM8D8QXNWbhJdDfQw7uDsR96UqjnJx8fxrG
Weh0ObsTGwRBNAo9DdtJz/BrWdhe/sv0DJn9QbbnLtRlTXvDerYWnygoiyeE
ja31u8UPz1c/bGCxR743Vwn1wdVKPy+WsOZMHOkoWRClfSMVB+R6L/sOlVE0
okWCe4LfGhXPbB9llaxZIyIcbcvgLSbD2sDcmH455wM9ON+GsPaOZ+2ozvW5
cv4Yuzms5GWb8oLnc8KMnxtCG8+gIbkmrOOkkET5jTUBzBAZqvgxTNiLGarG
wj2bGrdOQmnP8TpYMdG++JLlthnByADqgmUkRRdNQsS2Rjf0YWYMUVamTJr5
od88iqAdugSqkTsz3DExrmd4vhKWfePWRyMPZF6lVytIwZyMxZDx7u9sV5oz
Uno4m1IEc+7x65R1+HRr4ZGgBhkeuwr39z69vptuJICy8np7B7B6Vgx8vEXR
9ZYgO2LFyRt9dgd6zet8xEQD48mhuEggCUuTxO/1Q5rguvOqiF3ptK7JSamH
XvF7lJXTGsnyQ5TG+VafbEY/7veVnhlCtrinW/e1SSw90NsHnkLL5Q4NU1w4
/JwEHY1AC9osB3M9NacRC/5lyQHYokaqnBCG41joSvWZpiczFLkTCDcqCFKC
Q/L+rWVxV/0KwMqFFDKIPN97a/ff79C0kZJLoQQjAbgrQkiuO6FGR/FkLDn6
a0ojIoRgrEwnMXl+RImPsnNBcTKX5yL8QMbVIvdQCXZp1k4vPou4Ab/1ciWP
heR81wSD5xWGtJUXLPpfInkM3OmUI0PTDOyWq1MZVxxziMvFEiNWM2qWu0XY
O99flxGeYVPaxxBZbRMu2B/ybSfLnmwmlc2aRsfq0lc4P4tzi9x3EBwI04wc
WictzqPC9Ihg3hKGxKvDqfVvHG9YjeTXjuhFSTEbhFTVGxkN3x673cTdiKWf
qn5dNa2nhNm2c6gJkKCVHYVDnTuISbZffNmwxO3KT+si+RKyRwsFOept4F+I
tGcjX5uMCvz0FZJWj15qagTwxXhsLZaS7zmlW3WCvUISJjfg5JuLFCBvuTOO
IgPUM5RaOPkJkmDdTa8tZ501H7TGsNAe+tBqv5FYlwZkjNfLU3HXQeLGKUAV
TvT4CgCo44FOyf7AqusznJJIgPJd+pQu+IoZCz/Yxzikx7HjfL0RGwy/eVBd
qAQj76FCoxdx1rcftWfJh/jOl8pJykT8zWmbxJW6IzkKlfHUdbO5f7dKth5k
0mjBQ1Df9f1+CwiGKxZTtCt+8T0cGeKFjQ==

`pragma protect end_protected
