`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
TW1YcqU87coXgHGEr0sr7cErPqwjemFY5pR9Y1WUaZyQcMVDS6hweXU8pW9TaAFQ
+VCbpNi0f+fBJ5jmyz+XRiXJbSAugF1K0GP4IkTeFtaZAc42BVtffoOWg50mSz9E
y3aW2g4C1QB5yY4sE3H0RMFKzyEctc51AIhGaQF+IGI=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 10928), data_block
LsktV85SFu80yAkkolIgroOZYZ1OEnOv+6dGlujjuWxbLG7VPfXUZD39KNC/pgXk
WZo/Egir2ZDqwC8bu9g+zeJlVKn/U4157fvdXYA/+hN8tcJnJUgdAb9LjU2eQb5c
dQ+n2u1Ern6GD5TAPGqBPlz9yIh9PAIYVeSiaGfaBqBCanMRyXTsT8jX8ffLAF5g
VjcEi8xgpnoh2ME4yGqDh4TZYVDkYfTQVgyBJFcrDZAmNzTHBfVah9pewQ5598Wq
q3vjbPPh4kZlAMWe7QC90KdC3hVjEweUPXybBtbu6QScbLclP9yZfUOWMBKgFOM3
/So7773YbZnPhW2tFH/du+VhvaKmJ+T1zUjboEv6ufnVuV79jEKvZiw08VIz7QsM
OIDxcLmyvfyEFJxulGshslGz4hQdG9lsOw3gtlIWgZn7GhaJGI4EJU1eUzu42bH1
aexQjuQf3YCpyFokN94f6g85bObqV1g4wzsy3s8sKEn69mR8F/LXgTGoXsqFQLvO
Wavrg67yeAT56fLjgCkzaahkUofp/c8w4wmJfbZYXAXvVHQcggsznSvN5Adjjj8G
W6BSKGj0+1tUoyvmucR8Om17YkoqUpHR+kmTudbOefzGuzv5/H45alfBdUjTgvIi
HtCsHFU0Xe07Ye6y5pGdL/mJjCG5n1Bdewxo9sbmK2B9j501YbSoT4QbpRQknUCf
eptei8SZkfwFeNh7u0gywxX9LPmydQMJ5nRBwgCHGzZ5cdTGvWc+ULuY/spg9HV+
fTYL35CrIhCwdzOmN2RMzlw1Xrt+J8B0cU+I7PnNWChNr+aG1it4Xk3ZzZ5RUaeW
SdvzC6GGoktBAVULqJNVL6wWtYL3Zqc/bOMAqjMFvyWiU44FPEKouYNy4uFIxZ24
Wbsj5ZXELcAOxTi7i/2iuEyEI6jzqkZm8yYnfgTB4j9VERaj5Gh/qcN3u1f2fZtb
ljQXAp64w3QarUiGXHfU3BzvPfP5n9O5kHuBnDb1APdXw9IpiupWTMHTNh5FNhOD
s0AlhWemnFHtNHVadpEal6J4YtVfKzaI7BteGYCJgN23GFlcAJ7GAPAnhHE2Tc2d
o76LFNQM7Zv9uuvm/0zgBsmEFyGrda0Z14CPBwpV5v4wWV+G+4yEUEP8WpqRHmiI
JMVpxjkxVfmGgCcy2szKO5ob0VsbmzbF6CVusur2jc5c0Krt3VAZ1TcZ43vmHokV
UWqbYsGzHQfNRC/rU6FsdZVLwjEjuXb3LyDiXFb8+wb9Lk9hB0sXyZPXXILQu0Hu
GXjupEQw+/28xwWcgNPxnjC3V97Z9BUpOcSVKTDzp7GRhY08m0Ee8M/K4GsSPi3o
yupze+UvRqdAl4/x5VZlpWf4wUmpt/KXtU9Hp5WBkD/OornW4/Zn4elD5PajWFws
e9d6mIaFHS/U7FKz96nDC+w9xBZ+8G1R804IZMQhgkkgxf/uBZ3IHH1ysth64VM7
Hsh1dkGI3nSjo0o+Xy0z2gVVGPfoROTkgDa+YB3ZN96hKkac+zeaI1sL2S9iAuXf
+sLvFgmgzO1HHaYl2F2dzGY6IjTBkoni/U3baL9NgkMErrvFx2C6FJvcGyHtD2BQ
PqOr5qyLQSy67VIFnMaepwnQi3IXu+uNRjJ3AWeB+z/fqBwUVot1jVmTrvyEJ28J
DrtT1uxHSdktLOOm6zteYTm7xaNeAdAFcLcT25A1Udnq0fWaAn9nR+Sc7hTKmwAw
4Fz3IeN+gcq+M5hjbq+Xt+hbc0N5AhhPqDuOFcF4tsES31QIDVAPr+F94g2xXY3z
dLdEGOibT4T74COZe0yIjV2+95kVEpeCXKyJDuTJp/ctXBAivWk8OxBRdgEQk7nr
bL1SzQtWX3pPFp5NerGIkrhlvlryYDYX9+LJl8RvXpO4VVN0IwlCzMZMICJ/bNTY
+cRLyZiamic6s9DmJhgX/rIdXE55avki4cdsK/GPi/rZM5Rh0O/TJ+R8Aa+aLbst
iZPD065pKVl3N5+noDEQ45D/EnYaOeHQM/jqPvTRYfG78NNDQ0zjX+nQfnqyPf/a
EOIHcSdmrTAXUCN3yQkNflOeSQEfxfz0WbIWIJZ7RsKViljKO7/Ecj1JfFamfMse
QRIE49yiv9HLy0VthK5U8qjnwwcQibXPWRoOFllb5FrtabKmOwvRL0E40D8iwDLD
cdvr48Hux7A+zS4KBjAvKcUtEjlkQNc4dL9iWIN9LSTWITvqTTJLf2RqPvXo0MtW
TB5uM/VGeXodSGKZq/VRDdtx4zdOd3yBP7RFWhMq23pGSQ0C40nuilJdizQ/V8Gq
f3n3BJBRAQBXboewxvZhSRAkcsjTRVBuHvkQiNW57o1+ZgD0KomyCWZaWl3nhVBN
0xf7L/wKWSAAyKlmdi7TG8qsIhLbN3MlWTtzgvr0si7JLIu6hdDxkhAu5b6HOzND
kGSAHILM39/lBm43SCF9Y4pGooWYR6yEfqdS9cTcWxegDFdZz71OL4TBDn6XLGq1
XSBe88fOn+shv0ZdZIp0RqAjFx0zW5hjKpTaHdaSRcuzFQih5sbii0FbRCFtdaIx
2AK05cDkJ6a7/5zfvJjieOQunRCAvn5ZvCXxmohHy+oAk+MJNUe5n9mjJg/h4X5Q
Z8GQEyS8DH86Z+AoRDmMQEt+rv4iiODYf2qzNBM4kr9QPCX/UJ1dxUah2Hxkj4LE
8VtjCpOqX0TgxzBw/RfQQW41n7U4UBk2mWgEJEmlulFAAttsi8ZcJFv0brKmj7oh
2I6KaX6iPwulYie+z4YHnwYHHee/Eqx6MgVNlsKEmEL8v+MMVINU8YIpqmJsoB1T
t/q3YOdFQocszunTlvav/vI56TAiXX1jvQ16BcmrbsRiOE0YkwT6KGn1HS6KbTFs
fWuE6DJG1H6YR5XTK02vnVIRO4ZMR1vIgH7KR/1DtEqXlMR6mb85xIgEOQhaHOwJ
nwKrVrRn8T5U+BbVyTBygqugR85BR4kPNHv16bXO0Qe8zYk7wCzJtzxjv3qQ9H0C
MLUmDloTk7mJqGIdG7ykKpbSYIQ+CxpO7i4g/rpxpxPdpm7z05tukN9dFd/FXxFx
ovlB1bmlfWO7JKwWsamqBK8Kq4NgELw9Fq9zBAXNWGbctH4W5z0OxHRmgLSRAyQM
1N/yJdCBqd9H2auTcee3ItTV6Kegnd14XY1wS4ztPxW2AspbWhhJl1R5uZLOMibU
7p511Th8bCSGn7ywRcr9JZCFYYZKDUdM2tSH0/JrE1Bq8uuwDmI9pQj44qtqytGi
4AsBt10iU5J8+NzxEfa5LYO8ncAYvVaVq8fTFq8yJ0et05be5eRi0dAbJZMMkDcg
KL5AhTufbHH3R5GwhcLNBECZWTn2WfoHkh4U92VKQ3gSQRVPY5DBB0nPXUMb/2lZ
CYwVnSKJsn+l34peBMLVuZrzeLabpdZ6OQWdJhmNpRIIeXu7fjNZPjq3sAmPuDcV
UWY0SK5rEVh0WNCXw5bLUvxa1BaJlv9YVKtwug1qgTGIODb4J/oX/PJ7u3g6L5cK
B90QBfyuGioWhwYvSZsxhBDxegw081qofzqv9AZTQ6qNHxaOH6/elU3IXfOAomBL
mo6+GUQkiub9DFedBpoODmWCtXw0d4lwSvXqSgUcxZBkfHY4ZKBfXd20qvEymlVS
vV4Hq3EKIG2UNkoHgHshZoy3A4SC0FiikfufMvFnY95t0lJdAdB/e3DP5CXFbVsp
OEJmkDb8N9ELJshxEBJVNtY9nJDXu7jPCXCVExW/nN6tOdYo5+CEEIIduYD5ZIPX
Ou/edCdWiWrkjJtrg36lUO9qBVdJwuEECCzWNqNWkErIN43cVywT0g18WER/DLYj
1s/cHDLUQLitL7/2A01ehFeR/VR66tg/F68WSwY5IXpqQUiUOqL8rAnajJP0mqqm
c2wqLUKvxuiw2rQBJFlBJFA2QeEdw2AWWC8vPNr4plKxtc8qsIJu71AQ1gwK7JWH
aPveX7fRDORcA/gqrR7IFkiuCus5N5MDJ2QRHx2ywuB26fsrDX50GwvdMxxbXP4w
ugynwx3Moa/KsbKkuLEA7zy4mrMoQS69bMSwxR3gE7mbO9LCPR/ldaRE7uY4e6Ys
4qYcf+P6mrCV2FlInxRzrfUvdwclYE1H/U+maBy0pZT8MIYmLy8PeuPz1MaP8xhC
Hlhwckel9K+PACGRYNP9LcC0p7HXkqX9MGqOvriiqWLHOfxyrPRrLGaazQee+0B4
uKHAPhMMtH4P+AqiCN0vGKGKw8SsL301QK/qmA+kSvMFulBgOn4VxU1FxaV18NJI
pflklWXZ2QtEUSOWvjf+by9cF9P9TCn2QMwxsEZXrrQ6+5F9b1CP5o1wmSzxMYnx
OXlhNUzEhVCRz5kSDeoWdTT958m8Ig91YNPDuPHMkRPKkZiD9r08msCB48J2Sj2S
32sbelFmN5bP98cKMhbG9N+R2v7qBFbayVG1ptIK41w+n9WNt2PdWs+Bm0l4/y0E
kpjcMK5nYt8fuvAvEl95qZRyyCL3sTMoRutEbCtSJuZoti/EkPWSGzrgFyCn1DzV
XCBB1vJr/G66HOulk2xRbcD2ndWhwZhHkHXZS4nLtkuIfPaIEzYHdWACxMuCxdJ5
2bSit2kDJpzCFyw1T6wEptFyu+q8gaca6OBITH9upbRbbhbaBGLNSLnmuALBDGGr
7Tex7ZV0PavrcHvl2WGzjr1baxYIHkP2j9QKcVARFG5uUQuSlrCM8TJ4UIkcj9a6
eGOol6b0KVbiGd6GB0JNaQFkeAgageryG/ladIqnDaG30LvzqjVsU58Kdc6khKER
/Xknh1VGgDYR+Es82AG8VU/a2BwtlbHfGfcq+oCQVeh5z+kCcytbd9T9Lkz+MKNC
mAqoTJ8+IShTX9iea1/OZ8Ieh1U8/0LKslMb6gIFrAh+ihUfLXBeEl+6zjldTy+I
4buf7N6UANi8zg9acKbotocj7RyY+PyWUClMGPTZVy878X8iC7VbSvgVRGHa2ayT
UvuFGBfQYh2PNpuhEcmlbdWjGw6U17rnZgaMe93Y3HnE2n+ySJvC5oHtnn9ypP+s
b0RrBvhuPwBwLAxyZAAZS3/yDh4lVTOhyRAl71rccMxoHy/kq4KkC9YjqDCCXa9W
oMxGTfjZ1ChE4LzK3AUcrJ7n8f8B1vHQi1zDTx6mJ3aCnliS3hjFA4HtwbsB6W54
pEBbswRaIbGFtG9Tnk+OSkUfCOBNq+9etDSHgEEYJeRCdbtboRXb/ADQFtUh71v2
zOGePzSNJI7a9dBGZL2yyBTHCyj4SlW+o7BZBOxpKbI75UjwMpOpPIRKmGDmhEVy
5sTFgdsUQhRWJdksK/HJDOwVzINPqkwZCjXJCJDMbxKJFx0NGrQqP0k8TfGFizYM
rwXy49uBFmk719L3MNA5JomyPst9BmE2hiKy7RCu+/cTU3LfEohmEw1DNi117Ddt
wLbEb/+GyV5aPHvrgBXlvBdhfHWRbvplgFj+YvvPTXqanR4eBtD4Iqo3YkgB1lEE
qFEb9TuAaB6sjaR2qS0byp0JxW9mKmqzO2oG7n1VFGxHOShf3eNpz9u8tVaGpAYr
vWIRe4X3WIPFIQCWocYGuU3zyvWlPkRsHE2eBpgmG0cTbrn2ZfVWkTcTAVaSJfz0
8fd4epHCZYLeHiadc8syqYlFv3A8rN/fJrFCFFbxUZr1JHPP/AaGdZ7T1+p6HIQR
XD+iw5df/CLq1PsmV/gh9fcsync0d+18I3IzFd3AiZ/WhPEOUyb6BYZe5G0vaKSz
46Pkw0cLtWQ/3v3LN55OMepFhgNfM+OkUlxmGfOVzcXdY66O8WBiXSYlrgkAk3d6
7WLvvY3mDTLDvMd3b3547qfGJNQEdBViPlMnkLdUiofUul7tOfQh2u1i/EzrgxWc
zOqD7uEniRopa22AW5UuDmb7oEmyi9qk0RaxPtCY/Xv4ilIVLtsJWJ8bEmRHUo1f
rdCM8SbGqITkFqiTZeZqR2H4nsoSx7O7s3x9UVT2nUx0DTd9Shd5WboQZZWwcVoT
50BXVZ8bP0ut7N6Ag/xMmhO/ePWyDzVeb0/R/Mj7/aU0dBO4e3V3uzD+8mmjBaLv
YgC4pC7D8tjSG0pEP2ZkxnDIi7LNs+znBbGpIQQOKe0rnK2TlvjaFWGLRDz/CCmi
P3+Nr/yiVNunqQxYR5nY6dbm2Pio2xJITb+jm7Elgwlt3z35H7tmUS4eVCEIg0Fx
+hoBvH3w9zn7gHYqYG+ICZBt+G7hkGT0Fn692ymNGjzpfrK3KbeD1RHQ8l2EJ90O
gkj/eQO2X2nkv7sLFOgX52MCoKrd9WhDX0uVN0n9hTDHKR5oVHZW9IUH04waQEKH
HQOps/8uKnmRX77FCOrc54XULgUk/24mjF+ib6untj317BIt9hg4aeTp1dTOiqHf
17BWqF2Z0T4SqgBQD/pbOdIRCqGgAoJ8NlSzcM1zndCS8XnIaFIXmf5xuboVA3Tn
QbXr5+3KOsSP2akiH5MnJZLx2uNm8oltlfbuXzYVQee5+a6foKllIpbEYGjJEBNg
2pybH/ptDh0Ky4hP6t64hM/BvRbsk0juFBzZkBXYvFXXfD/inMqJvYoF1jQz2bUL
Q68Edr7FIOEfE7R+YpakAdVpvNXdh0Ga+clZDprrwY6OmaU6AkpQ5nufIazORAen
J0kAOqWqsZXSd6SfLOS7S1hRoKeL4xq9211o+HAYTHaqyLuUKC2MhwyzuNqDvvWc
ssd6iOoyoSU4uMMIIMHgBJhZ7BYQYW1rxyV2DiyHbp8bxtb5j+SIwEcOIzs5A9DJ
oQrJrj/qWeLqVGFD4hoqSXwuTReybPQt9ATn8qoSuF0YIq8CE8kkv4d4El2cnhpz
Nj3eAfICB4OPkKhZpyskNUz+Ul32KWrjuimMMuw8E8JQndhf1Is4Hg2fivsDD5/2
PsjuIiBCxoXmN1Z4OyVSEurR+7IUOVAK4PdaoKeozyhS1a9UMILOafXKiCK7an8b
h0xhBaUateO/h2ozdLAEGg1ZjXxD0cC8iutSNkBJgyy4n+eiIiHgu81hJXU6/YX5
LVKwt37IL/SLHs4uSs6esPjfVJ3sJ7DbnLQ/JbJK1LTVuLx1+z2D0h/CvvYrvNtt
+jATmU+UwFiTzlG/fU8jT83KurXvVGkiMudCSBfmSkeEwjRenPcJlietl9p3yxbs
D/SRsQw/DXLO/Ai6eBGSNbQGyvn7VJ7A1I9BI6gVsnMUVH+I9GCPvax/qTp9ZfVp
+2nj9CiNVP5du/MLFlzwTEKcjj4sc1l2PueylkozSzfO8O/MU8pXupEM/6tY8K3i
GohCULo6Y7Q/WRuwiMoQYdZZ4RuqX8kP4rSxQFsTgxerrOsre8XEttCNUE0iBMg9
MOaYinDt+iigwZ0brnDtMpuO+0K2pAVk7MZcC5vnHL5f+fRZUV2Ud07TqupDqMav
TpMkrhozTOpI+ggJ0ZodUPPSSjsSm9P8I5NkMPe2DBfQCmDgQ0bHXP96uaZjf9Gn
Wfi6vQoTeY+rODUKgQ+BL77KiInFWCzB7P385Qh5AVrY7Mp6XRPij9Jg+mEpPykK
dOFSCn3H7+GN3oaUgi+s1M7POE3IS39ZD/xo9/C6+T1W5QX6wdQdu5bqIf/NblL4
9VYzyPDII98lZWc7ivYVsmi4YK2v9D5Q7yqJo5FoMAja0XJOdTixN2BM04QqqTof
EI2OaB9Xa5Tq7XkvZ7eLyE/3tKLclbcomt1PnIWtYCNrJOhBHdT2l2rD4f9H2BLy
KGFv5MhqhlEdv3XilCs0YGMCePrQRopbbGqs7XDD6fG2UMz37De+4PGtwU63Oya9
3XEe/vus3JHcLlKv8DYLJAAukBD1Y7SwMFfuLpyjM3mlRHvgeHpN6OFgpnoFBP3n
D5dqJ8ywB2EY6RWmmaK3A7w2DyNmSkuEP+FzHH2Lf6kCYrz177Mox4MnVNpp8ceE
z2wrTJWwVlxvJyJgrElJGi0iucZ5Zb+CQ7FqDI6jv07Y51wdMPVDaqmdWAtpa954
BfdunV8G6PVY/4Y74LcUIuG0XXYqqlrUuHero4bP90hsQ6PlxRoq0e0IqB61RtkX
7KKqVoyNYGfU7Rt6qcPeJ6UTQwfSZudI6TbSzzL3DdQPz74AfzbCRTcMMiDkluCN
cq+20OwkTY+8MgrdsWqZE9osofmJBjtnKeQqjuW1pXrYSro9+nO/e5hta4fu6xt7
lOvf+4z2v/fvZK96zwDMkkxxY5dLIuJkep26Q4Py8JtFRXk/S3282AZLHSxlNKOT
Y+4f68XjTQq6Heex0RsSfSGmBNt7O1qhJjZEaif4p/8euLx0Zv0dwGZbdyfhVC1Q
w8vCVh0t77EKQs5FWaD5r1Hb5igIlfrAsod89vN05AbOGxiU++zAU5rEowAa1/19
72ldwbHbAU3U3CjVzhplphQq7PcYFFgJ73h2VzZtR2tzVLGBgJ9LutbBNsu7PsPN
V97T4PSVcx0LOVVg/cLxBNLqmLcNn/tOd2tOwjOOezfTTTCU4vaZN9Re39AnbOqF
JPISvpf7UBnxdiTZ7ploOIPnD22CS+eQVnSNIr4hOlpyh7g0RZCwhlHfW45JZKuz
F+dn9FmgNnTSDCcpWWMxm3+4u/LP3NrOOOPl9j/Io/CLntFgXCbXehZUaO3tylq1
uP8mmBSC/vEzUUjM5nQAHs1FlyY5M5498EsRXR4DaU4Q0B6ryIDRKs09wvxD6Gkd
6hdBDypAex+70L7Ho50I4fvHEOrKd2tQa6g8gcRbdRn2omfdem2TAAibYaWAjFmO
lzR8E1i/xnh75IrNka3Si9w038xqVoPAVIjd9ah7wfG1YoHye9vmbD/e+mtDMN0x
cWXLllSnRyjYuMldBBTkjI7oEU8KnImYYPEqLUpa7bpFHDXenFIT3VXWTMOhl+8k
9kQPdWe+UjDuAjd3GeFfB3LVsBB4QQc3q0DbRS1U8NFzflSRxuEqj8M9pFGF+wuJ
BM9fncvubpoTkYNVjrrpB5oi3Jl2t9UUss49RcpWLtTuZZ6uEdd+3PfXQemsN3Ib
WuPgQf/qAXXP0MobEtRumiwHaAt6wnldzrkD725aXYYlPdpRCDFgD32FfuirlhgO
w8w8fVL92JTGufuA7Q+7kyoqtkGXSpyzV1Xec1xkibfY6wEcuUkkcbJ0VE2NyWYk
MJF841DsAU7j7VhXVBYqQimG3Fw3XasqRA/Y2zx9uDztbujCEj6tAbZV74+EdYG1
EB4laFjz60l3yLAvF5p4CF3p53pptY8WP7+7BUU62mqlLnPlv2U7kHF9Zg1XiZu3
p6pJrML1FeAWhJilJZNnES2/jeKo4je/xC6o5nBhdumTEOi0xXUC0UcFv3XK8K9u
rDIVwG5lR4/bDp0TuRKdAB5be7+fTp2xwIGoFW+sSEemUBf9e4AAAX+mkGYhNu7P
w6q1fzNzm20R6F9GDrK0Ralf8SUzJdyvzEKU3Ot7tKO7dm8fziJ3dyrixGTe+gbP
aqN5sWK7JcN8tCSftP3zhnz2Ryg8Cg71EY5k+r9gvWp8cvc9jH6fQDGH/zBTFVi4
WkyUiSPRfB9nFMlNNy9I9d/RsHVoxC2hdw1QwEd/hB0r+COhuu2ythZpnxlmQBNW
w0BgdV9Znvz6GU2Jj/0kpV5eDGdI80n1XWNkJ2550wVVdINxfsS2FWZMxag/kIsC
FqbwmPxALRkM8H8GyEGoc5t1GaPh4NXDeWiIDw3/kRgQG0T5iNBP+smE7F05u6Y+
F+6tuAM7Sj5tI5F1rIwUSSVYhge4UJOZyTYdh9vZlld+GIdvsLTWJ4qWSDNHHKyb
cJHCl93R8vA9yB2/yOEYGIl+FUctTpecTQBBXwN7ET0PcIEARK5Qg61yBvbPf7dK
5AAS/aTK9YfzOM9KJ4hwHJUdCjHv33WCcTr9WP/vpAf7LWYKhrwOKRKsb6lPnThR
XLwprtVjGysTCadn8CZ119Dgy6z3uyiDtXZFmbN2NVb7xroEshlfXrZivAhTD2Dz
FoVlyIajw+O2hnuOHukZ+oXTR8XdjYzSSgT5Ne2wHdODX6aP7iC1L3M/CM7gcxxt
anE8SF/nvThRLjIXM8hw6QUdGJA0NJo5bG/V6vLhFGUCxHy1W+EiDh1R+uaSIFBA
L/SxrIxTZHRH+bn5ys2obZWgSYUXNF1ZtgYqvMEiJkVnPJAYyjEA0hpkaGi50QpR
CniAQxtxvxvx39sjzopXRajd4oeYrgc5rKAqnAzgl0awyzIP+oF0Pfkxu008bKK2
DinNb+DDUTIZjr09cTZmiV54Mt9qlDYxZURdQZnCKo0l6w+dpEUtmbbcAH+K+w9F
WWfRLJq2H05zYWWkNwrxIx3scEzKvKL6DcC2giYQfBikDL1sJTO8TCEIDlpQG+EB
8+wAu15ks8HzOYzb2zJKa225KSP01IUmdywPqwklpeJ7ge5pUpSevhlwYOspaWBE
ovhwj1XBSvgtfJA/UoKqNtJ+elA7DkqWcWgLVQgQw5DuNEdC9U70+QaP6hK+RFUD
WiESrtbpdTQh20i7NF0uTyVKGy3VukTztERJ/dAnUFuepRM4drOV3cHoJu7ErqiA
lWEEgsAjG99H8HMIvpgFxPfCABAxiAs5Soz7yit/8sz2G84HRzgdhVl/p0s6cYba
vEBcJwPtEeDUXJUH52tt9D7+E7H4l7JxE/QJQ3kuPbTHUeC6BBBUES2SE5P1Fckk
rIstqsknWgp7+7LsGLr8J8o4m5jAx+zv4PG8bmXo8bp6K2aZ2S7DEB6pOJ5jEj3l
wBaauQWput0laWOqMBqUDHRBAyRtvTdX2skPSNLX5e9xQ+SOSkyv7Q2isAPd+l3T
Pu+nq/YAAJo5GB5F6owuE3Ma4lLokRChmxa2PgZPIr+6KVNUk+3ryVe+9AMe/El3
nLBO5TEm7H3IDu51760M/F7xPz5bA3w/Bc65MRassZHFAUzZVSq6gQOx2FyZy4zE
pIzSDiNXKVzyNcRqKz/ABmjFbOKo3AQIleZWQVJnOBaopl9FW4lg46GyWIM770FR
udhevdev+8vHUFItDrKhZZI47kyrcbw+zDfKQ0F+s0OTUKrsT+FvfNuosW7jB+nP
YLtjtPzQCKO99ECRufcRMY75w0c8gvKiMW3c45cAZMkhGiBcKxpn9GBknlnrOiMF
+FWUeEXKXwTvrybA6JMEt7q/pqPGbThLRh2xv5/GmgwLXuGke7pzJ87XV4N3l/Um
OOZCiyuPwk0Ui1N3O39zk8yXeejU+aIOwz6FYfDRyLMqhq6Eeq7SFg/yHbJ2vvWL
Ez/HXrQzCz+JdB+gU/BBr5EOWq+9jeWdOfSpBc/xYcfJtyP+g1Oted7Y8yZEVs4B
e6typCV2iZp9h2xQf/wBdfBlgkd+gynG/bP4AWrQL/D0Nm748+GeEid0rb2WcsY0
uttnkg9bZV98QM6IF7pJkfjZ1zOz5rqhV3n8tchk/skzpnxN7ggijHmf1Mu5cQ3e
6JL/B/8SEOqEd7+JKhgri1cx1LrD8Qp69KjLWeLCbPU68V4BqkdkAQX0n3DmXcan
62ZnNsoihK2DGg7t0nBjhX+vRe51N2+dhhYOaxGgWfoiyNs4D/sd9qaV2s4s/dEW
eeqHrD/xMIvErgm+BvwkEZv8KWsYKNedEC5EEinxMUmh3TeT36i989cpuhB15+kS
RhfFia8T4yIAdvXN+9poa+BocO3gT1AgkaVFJfDi99d6vCSXsy0sGCIyMp4QnB4p
4Hm7cbs1pYvTEpdAZNVNMdEU6Buu1yV19RSjPemUjm2/glKH7Ec7o+qJtaDGtNgM
LJ2OIwLdBQWLQqS9I7tLdw1Mw5SOtpCoaynujf1iQxS+0OJukuhcmyl3rIS8hdKd
cEmIVxMz26XKyP5/WxTP3WBCZrZbXlzvAx+HdH+njy7xfsHAi7sUk2IZLFevNpAY
3VKiMvoe1VLmyaQciAcagj7HE6XODgzDj1QC0Ue7C6aAFWCa1kzbDj22fi30oV9D
GdHvqonXFmaZxRBQyxkU9RhfVJw4nillpMMYCgQ526Th2CJ3r3HETcWCV7fwRzQo
E4b5iOv4t6IL0iYyLTmUiFB7sTn9keSXRgel12QJgvq0/rfGxfFPjTtjCphmdOpo
N4yxSUrb7febXvKt7Uf506cT9t7o+QooDgCiUUi2XICO6LmrDHlrp4nwZ8oz8oTo
2dow4DYjGFwyqxKvs8CkIHEG7jdCJMCsYsBa+LVysNEcb81fAhgJEKZFbSl8yJtw
j0sY2zQOP/15Tz79He3WpLWyZipPQy4o8OIlAQeTmQEyftSaaB7dZqKb3J4WwKb7
uWUiy2SiMUtBZ46KFu6O2e027qtwI/QHywYAftXSbqNbl1P6ks9qdSCnxUrvQ1ig
BNUDdgWmGUb7owYeLarkNi3MjeoFbBHRipWOSKrNIQwvaS1z2OuGaYorL1U0i0gf
TDfbMWsKVij1+a/t356dG41wG12HftGC/QIgiIABMrm4pYb+lPSonFuf0IrtiSYa
5TlRY4vxTRLDfHAL5JDdbRo/MUbdDovV5Yzevn8Xua9IKIx07bMU5Whw5r8JNRuq
Qg7Q41Lw4oA3hW55epFfXJZYtyAaNklVulW0cDBTmB2GTIdRcEz6ETlgRqGJR/SY
RUEU1i1Mi71G8Ir4Rhsp67mRWruE26MRgCeDSTpOnl6aShZvo4sQp8c820r9IZTK
poa58XdIz/K1IIb7YUECJsmvAFwRSe/e3xdPYq9mytj66/Ogh3ii/GyGdt2oTLFm
y6m+BPVRbc5+V1EceinWgoK9Nw8DQ971XQ8127wnpkUtT7Jkk6nkE0DGE5H0NvJc
Aiud3X+ltvmdq5RZjbXFQT9jaQzhtkYWtIFsVLdhC/7GakuJL1FoaMwtEbuk4BXZ
tNrGuGM6JEn4EzYJpj0s2CQPQO2Hl1hkSSKcFxHbVOdSBkLm4bzFmoAm+RhvVHPC
hYi0dqujO+AlUeOzssiErgP8qaaGMqEaiEsKmC35JWf87CMsbPQlGTekajed3EK1
JObME6ckz6EbkvBtGWPwIls+/mCoRwCC0nOF1dRy1xJHyVKgAERof9Mdc6y2mLOw
7CW9/97JoNq7UaY9Dl2gEpeZywu5HIXyyw3GST9ZT6cjt6rr/m4t/3ogBX/EYG/z
GRjazsiO4Y8OGUxJA8qpmEXBCohUQGLnucD+1ZF7OjnyBvUolhOSLIf4zCipHjbX
AyfDqR3aiSHD3f34G3kyJ50o76q4beomNoKH7H9xFR7MtD1VeB8U+hmIAyQQGgoQ
Df6ksPJrhqpcRTeiRM0LCTi2Qd+oTEMeO1414O8u3o+kny5WWOf60rYEtk3R/0TB
zJyYCZU6uE/xG9/MrRQucPKB5rwqLv5dlN1zDqHbSJywv3X2IijcxdyB94RaVIyS
bpHOh0NY6HtxC4da2zG6k4FOYuIf/dOAKxMozncz6g+0mvqnTckNXcCIgi22BHLE
Q5dJO4YvaLk7l4JqS5PQrONEb/2FV2jinrJGHwa0VqnE5o1DpBEZW5HHcaNcPn5j
1tdcwiNKhwTW2poQmE9fAjQEulqFFC/2ppJsKqlwjmJpOjyllaEdEOAeAz0EENLY
VGwcdgaBe9HBUQDmxjGzqMfj86N3Ah2JL1YftT0OMIUOnZOEsJ5TEjyGsLg92DRN
Y3HBXckMyWh1mgNVKbgTK/yppnJxZK6GYRJ00nAmOupt5N/ZJbvRT54QFnuayTJu
ZgwjedKCt+wSgqXT92ffxXlbkUQ+tEMs5J/kOUPVzkPXIlLxogSMFvuKDrBZa1YQ
v1lWQDH8SOg+eZDSRamFHOgzU/PEyfanVngl4TxykZQyl/sYXEb2uOwiibBWjkBZ
zAXjuhH4sV0LJYZ4Vs+1+c6KmPAvo4OeH2gH7d8rHmjq61Lj3qVLMY05fl6GuBez
rNOz6DNzu4vPXfq+8Oh0xD/T1V6ozN8Yue5smFMT3Yb0ZCVr3ptcvuDvlqmt7H8G
05eYzovyoqOn/+Qh1VtnqC5woBN0G6Ql0ryp4qanOzXdP2JO7oD9TZ5i7TUGUxFg
GqPRNhDv0DyUFimArKswaQgcWkl9MZIWLL/WBCydAkH08TJECMPSbNGzXrusaumX
o48XqxmiqXww6bfyWIM1oacnhujtG6+Mtd84Fr/FtpKf7RPwdu6mTAPl0zMtOE/H
fupmu/IgqIc75jSQr73L4heG8V3MS1UJd8x/YL3mN7MeYZBumrKZsAJYZhqbc4CP
yaXTPCBowG7g+kB5NH+axnNmhO3oJTK9wfjS5sdAh8qIyebUuRIGCgSZGTbB1DLh
ytRB9rBBIO8VdRSSLSvzPW7lbAkE/bGKcx/CSJKk+Ub6kYfZtdvQrgszMnzeDKH+
V1xB3v7zeAFQMRGFbF062MkfCbU+0plZRNi9iVQITK7FGM42RjsJxYkQSixQSJp3
frZoklwGPI6JWR7ujye59Y6b6bIpaDtZLqLW1AojLaqxNImvV4cKcjxCzXzDFvlV
EB4cSmNbgDdASYXYU8/AH486UWC2KsumH5UsvycGD4Av/lRqm966CiXXFJhFH5FJ
cdJ8uhjp7BrShQfxMP51QuIlVbNEoA8TQzgljGHIe28=
`pragma protect end_protected
