`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
EsK6g/Nxp3/JGXwVyX/tqv/MZPbkISSOrkw+sQBu4BQz3dKdGlBdr0E35xEdVO/8
OIqZbOQv/otCBJB5yFWTfTV9+kP8RA7HKwNLMMcqTSUUlloSpHtnijDUNM6bYHMK
vS8w9dMRkdW57pu0HPqRohnDuFvZ2q9cmHGlN64quIc=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 4688), data_block
rHWEvjX3W1O5Ts9FessNhalTl16tK4XVx08HChN1ricg3KP2KDgC9W+Ga5TYWT13
N0mGO7QkxVrK+DmA5Rkk9TxWJ/BnEY+uzflAjqoWewudBILhXVj+b7f0UNoiLyaQ
9hHuJpOM+npPF9Iby8kmBGwwjfAFvPEECEQvBaYjtiPkdUAhZUiYKzqT1oo+Mosh
ZvJ031GTpKiQ5QSckHEy8HSlDYHz1T5AfhH70AO/lVQWLJxR4fMwPeFZbuT/wx4s
C0+WgEapcribIf5p4VWheye1d+Hv1JZ5DllNmL8Fa0tOF16WbnKDNHZ7/ipTzSqs
YvK31yCCRe1g88wG2fTMiGLvlm11eBZRrC2HtshjsTeiMx1dfdcVhl3ss9eqzer0
U1AvTQ9w/3M9Kg1SekeGzJGqz1DHQDdCR7nE9yrt5dVIWKvoIwGU93QAUTPlL30Z
EJxTKjk1/l2FH+zeL1/XOKZgKYbPr/oN+knohbPndmuFUYgOzsDZopCKfYiJnR9s
NH7iGSGb1UPXWKZRIM1XhHg6k6EVqQU7YQuTom4wU3hHPqw1mRDxkSZ8k9ntRFKc
Jvn1l+wOzi9fMlv94xTPMymkI+2RzF2Lj4E4G7cF44YICbogUqkykRsf5Cagzkhk
GZ66J2ywQ+3Aj1Lo+bUGEWn9MmRDgOLrAsJuGhV2Y4ilvtparuIclXhCgPPZi4TV
DcygTk46iJ3IEJdRPFhAWSjbsOhgsmADjrEYAEHeZEqcGDiKLfY4NtPzRRYuL9iY
UAdM+70M42gSWz2R8VZrXlHaZPpCRSGOMWGmKMj+nZPWO7mL/BwN9Zq3YLi/z1XK
qInH32LOyWoYs3nVwaIoG0AG6xMMhkPQPCJKlqjshmlBnlJjqiFcuCezuQ72+6A/
W95oHNPllIHInLp2LfTwHQOZsBzpeYIJX4coVX3NABVKYotdXNhPpg/NVa9m076j
EWMPLjQk6s+u1DenMAjeNMmj/a5H77zHPqQ5gT5E9aKjBHBMJ7+Lr5uKffqzmbZk
rWCmaEOKN/2uu+1IcfDG0yceY7slJ8V/mqWLzGy+Efn48vOvxDmlvIV8xnvrjlcQ
F3wV5s5QmgPQ/ahiI2ZLliYw6HUUcEuWCqDalEsGZJMVTLFdAeyJ+ayeyTa2l+U9
l/VHSoUW2xBVvRk32n7rhdJZeswyUoH6dE6w/P8LsDn00AV3dW2E1KAhku+FKQpO
iiXtXW6MNU77llv3DoDnz04BXoTjFOhyypURCARSUzbI+Qdt7pX9Os3SgH0+f5X0
E9UzwzSf3/91tBvw0/gybfVFHn8hLXqgCK/7hmrcDJskqXC8uXXCZtmxOBnjrH8k
1dP5ZPfhoNXRcwG62a6fU1GZsCeCWPrE276wxwEw2Uk81cFwgGkSjMj0jgDguc+R
+JDb0e/+XOshnDGmRJCrcf2FA6mPqeWAkf1leHcpzveZ/RznsdQrB0tHVLEc9yhv
1QD/AkjCrVzUiEczxUUgDDQjKIRM4YV2DV6hide2Bf6wSQsns2wAJgMKsgA4HW1X
xg8DZIwDUHFTy9Z5kafB72Hwg5tUr3hgrmJicvK0HnwVImiVHRo81iZFnNj/HI0k
da/yERWx2G80CXJtgYKN8XGbfg2e5FV42YvYDV08ef/i9u8VFf4RrxvSfiGP/hLU
C24g5glSjZb7dUpoYaAriNui7SvcACtevGJPO2Zif0TfCnL7Hkp8ntp34sKG8e7D
HA+fxU+w3lbgT64dwTZnr3bEar6XBVyBoaMOSOsi2gQc3NHpIkL5ZJFaeI+Rux+4
gxivI4ktp+bQzO45NGjRAKQY9gWWJ91gqYBd2ammCA/tWj75wUmITXiLvWk//uTE
ZkiUwXhu+QnjFFK8CTkaEZq6lGoQFyEqQ0Y4gyaLjKjGelpxazcO8Ow6IxxGpgcX
1Poq+2PKZTHPPH0Qeps1P8pegFW9CWvulbH+BTbP4zgsxMftoloN4FgWA6UoIC59
6ta7LvX5POpInY6tIb297aSqI0sayxwEeMyl0FhZwHtLgeyaloQNXqZp2ZWOShru
pgWlKBw7OWWmW2jpKIaJphnrGIStKAbMVfj4S9Fe8/LOgbjPyZNTVPKFSGFP6zoB
+/meeZMW0mUJCv7mkKOt5XmkeQuLkk0oBo0pLQD7vx2f1+vPxGFgVOLjEtPfLp7Q
/m3JzYsIAMjqY+uO1yvRnNJY0K2K/QJX3KmbuMyTjFURvARfMVkBNJqSgyLFO/OU
2f5QOmF4AHDdwsmb8NMjsYyW+94Iv867ya2gOdFNtxzoiZ45TlsQluGOdR6IaomY
4MYg41Ft1bTAWloTXzvySTq3zYeZGjGZrcA/hOW6D0pJ4Ew2c6kNYvz1fuHofD/B
sIOtVRGjyb3AEhcH+924AQKKvKO0jAskTDkI4sOLMxryV3EAMUZt/JFLnvHgYDi5
xcz6dpZlQYXLJ/pVHrLa/utZKn0if+F/RkJgM5CE0m8+bVRoPI33+F7c2iHdadre
xfnDKZ0phrAlfJi+IX2c6OBXRqHEpIBOSNlXmLej6tPs5ovwuvp5/0ydJmCKU+P+
vgB9Ie6fbYPOXrY1gG/g7eeO1xgDOJ6/f2LBPxM8f/2z1197M3Nd4u1WZlk4oCq8
Top5yW0abtzmwmZi54lzVXipmP2KeYBlXOH1ALiQ2hxEyVUeSkJYLxkq8aIck0id
gIMe3fS3CU4NZF6xA6g7QCBX6Hvuf9Z8fhpnJVvveik/Tw4L6JPAlfvxY7e8wBQU
0k11mlQ+2D0SpgjQOz+drvyXG3s0bArVRZKc2LrYxIVusyzkFCUwoN8UMPKrmCxM
blR6/FjTnt0gczpR9LANE5bwWIv8Q4Dcg/PO0iLtOoO3ZQiFDFJf+hd7poBopYGm
6Wm+oAwWD6OCB2PEhnGxIgYCQWKk8PL+il87KLPajEuV+2izTDRM8Zthyommi0BF
R7tJ4vJbxYLy1JeKJ58VrSV6X4uTdKhJ+L7ZfwWMHAI3CEjAeGhRjmoYTog/bLuu
gs4QaRCnDBwglug7rEAi9raDzdPoBVZ9fwoIf0j+1d5t4uA8FWXQwGViHe79EbWu
Y4PUEBUFm2vdsojTTNwjw7AIOWZZBixsxnNl/k0YklJkrv1Y7Yn2ci/LBGCeDwa2
/kao8I8nVAuOYM4o5CiD7PTYqfkI8HymQJaFF+6YMlrOGV8C0PCECGSPIxZTe1/u
XNXOd7CIfZLCUf0DEFQSamuvgpO018APrHCFDOc2nfvPeBrYHhgyS/5wuuBQ+UjZ
46pvmFUxIS7PPpQU6ozLW9VqrVXIKjNWvW93Gvb+fMmlbdBxPOQtmg8xKLTZpYE7
wkOywribOpG/+OrhByq1sY8wbuIsColZPYSE+SHfnC+T2v57/i7Sm+pep1YP5xht
cdikGxBqv0MFVFGuYcFY2uKCszxQiNhNqPPf7hzf/2ykwfLnrwzZ2a92oNkgTvjk
DVa1Ms1zYWw/NOZU/K2ddEkwRE/te6Gwh93QqWIQ5FlII15vDAIDjIh++TgWf1ol
4D6cgFssiux6guLNql/pBsB6JySAutOn1/WqA+j4NDKhGkLajvw6rSG56smWngqD
q5KdiftGQXE9ndBEndQWdpE7np77vdNJizSc9dhCMtDgMJxfG3bR5UfTwmCXKq86
gfBBLYtLFu7T/jqPanCYw9AXHEUZ8NPyUiPmzyaDmhiVDfJ4OZjePZMXOyI+vKmy
0SqTY1SzH3ZLFSV1FNUPPlpKeGiBz/EKFUsV23+Vk+NxtOnRUnqmAfCCQ8t34pj7
I5dv/3ijvKgg3QyauQJ2ga0fChQmvn5CYdaKyxXVxZltHPNB6iCfxJgip685TxvK
GAzHUYLyT5YbyjAoBdLqCm305o/I056MalND+TgmklXxE3vbDPF7y2ptWRI1eRi+
+hQ7/sR4Yu+IWspvu3TOw8syuP3rOiiA/z9ftfEHn+SNyirC6z4etdg3hCXV9jj8
Sb8A8m4VXB5GE7e17RIUTgo4c6mzjLfc2TdC0uS3f/sy3Kx4S8/ZIpftHwgEGb7D
dzWDFuRFo8JVQkTyhKuVQVA27Nb6tXgyMx6knLxy1snfzQTMjJ8XQPp20BYDZvUF
ujy/bVJo5Sd7OGwN5VZiwzWaJpCaRObsZewH6ZjN0y/ic8PaF3ZjD6hFtNgGtk0G
I3tZhSdfMNQV2Q10pq4buo53xwzXlJ2DXebdoGgFTa8TC4LxPPVRUl+3n5wzprrx
ydWA1bEvvWAEmzUSc3bbLKesjaqLMeadUZDPOP3P02p/oDxDArwpqv2JzjS8OARK
cXPKe1hnR8JucXZP58Tdocrlqoyg3v25MXF+i3k5N6v4QTCSf2PY0SqXuFTihpjd
LFRducK0F2ou8/vufza/EZFmLemWbEe644w8OEHImQRk+y5f+FwaZtQSKE+x4c8N
VxoiYJJ8BHwtbOAAhnHXe9n9D5nRFO3X/24aJH5I9E6g5v0/i0pAwNcylEb2MWfy
IYMoX0VetD99lhdxxzjxBhfIDkX7CfhqzxMDDkX3FlvXT2HBpkrj8GuWtdKkpDGW
/KXiTMuqOwwhGk8WgcfSvBnR5xRPVrLWWgDtX0tcniUSyhOtHYL7DipgsddutCiY
WFj7rxC9jOgNq+NHjaUW+mEUzT8Qrx0Iu1YC3nZ+7P6n9NkDgLXEaW7GJ6rpMk6P
xnLhv1e4FJ247X/KLMpHiFnjuFoa3bc6eAOeyosvYBk3I5u1/2MDbkyPrftRSJZB
igS3QksRTTOOapfLhZVDCGEaCVOh46v5drEPQ31ZWXjS6kEjb4Cvrdlo9JQ0DiOw
+mxLPestEduDjTp9/ZV1J4YvR/b4CB1PLP6VDsO+yxO18CGchhj5iDeUtjULIher
f/ImbnHApJMjw7fWkUQ8FzzZnAau20t24gKNGs+7HuihPulWixrsMNu+HELGBcQt
HkU4GGG/EdtlyR1Nv/OTFQshad+W5j8KaNTZQ9otbl/m4ZRqPHyBDKk7ROcHwBzE
dhd+QHf6BLgIbPGpx8XXXdXlyz3QSFpaIcYw8g0KKu/Rw/80XZAQfqKi85nvtWdX
3byMo3dof/iUf4nuk988jVdvolJOeAqtt1RwTpa/ix3rRY9lm8jRhFiFZ0cDleOE
uCJqF+9F4c9IasjR7K7Q2m1wmFfctuiu/C3wNwg0DjUQtrvE2RYvnEkDLFZo1wD+
7n0kL4+i4NhH6z3TkE2QZ/GBum8axmPRBWq6L7o6F3H0763RNHozTWKOxffSDFtO
MJA3NC735EobUTKRIMpm9Rq0qLzh9ozCjTz5pO6FO+YBg238AsTa3CUuOML09PrW
m5Ej39fTWr1puSBSyfdsPV2cjymYfrweyPE2mNXDwCWjvMR+yGhaAwgvGWtqmxpx
2HPvI/4vU59LjJTjLP6EuftNGK/mDzC11ArgcjlhGoSpGjkCy64D2c2YYPaImnUY
0bHMqHrsgQrtMliGl1ryxTz9YbrZwe3zK2KWZSIVun+iYZ1x2lSMq56Proa7tNYm
4ASResgKli1mgaUORbSAyZQ9HxxH7GX1RCIaj/cMjtFx2gxpAskZ+6M5GFSFi79u
24qSFppCp0e86BEsxpmsAK862Tn6ReFGaPGZkPlPnBp4NijZu4cWFoZ2ZwFwp9wj
RgQ6c5CwpXyli/HK6eEDoYijSmtN/PdQL5j+g39qCZAStvFU9BpNtUth9Pcjm/+4
4VucfuazM4i3DpPVhO2LUpQLQvrZ/vsL4BzDpKbT3QaPxlQvMHfD3Nkad4zMU/yU
42EoiEmfNHkKs/eIeSBXGtVMVwAQNqUQ7oR0o9t02sdN1ZdJVKLuBjhG1IADIA/+
ptueqWrXqGgxSxeH5VSaKqLpvEMM9aILPkobRSHx9fIucuK4mal0lHsn2x/uf+/b
X2maNwPU77ndKxfqKvCFApVQ2YSaU8Fc5dc69Sz43vQfpIAsCQ4NeqMhRCrK/2ei
IZpJcE/78Hq30nLmgXWks28x1DKZe11g4chd5C93rWskLyfM1PpPFFSAYZhseQs/
E8SxMQO2csnz6gV/hsun+cjDiTTAOph9qYbubRCJADQ68l8IszMfR4FJ9uLXXney
BUJ9KJK+3gGS4BGHuhZ5ceflcJ4Pqg9hyNVh2vyYMxdMrqT6TgjXTTEOKJ5nhEV7
2P7KJ7c6hChTWJNO5jcYKJD9cm8mHHFjtcKF3wH81jUgZBxpCIG+wP5n6PPmJNOO
idq3/385whWvrNTkHWpu5xoIdlnfP75UEpR+zYRzmeU=
`pragma protect end_protected
