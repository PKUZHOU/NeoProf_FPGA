// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
jHc27de7c3Rw5tvFVKCnEXQNA/91G7h33XWIPxCZ52QNQIkNH7gaUx6wg5y2
wF9kAV6NbWme5KC06IIs5/oF8yK81qtaLZQOYic+R4CjWaXXb2x5/8VcccHM
bSITCJBFxpHe9BxN6nPqw8bR6QwbZQCVDCc0IPQrcf4B58rF2qQF9DdDbLn2
yprvUoJ3mteR1z1xXjh37dMpp70yag+sTMc6L86pxlkVJBIeFHJu2Ldwye1u
lggFDtQSSiyr0de7FRmSxl0YBEiSl/mmrANjr/HC28d+UrD5SganOvQlM2pq
V3lE0oC5mp9VNXN7ilCOvMGwbdnjQRx/K2rDOKitMQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
inBJsyZW9IeLW1b6/c35ELNEqxIX4NUIYDNePiE1n95I3O0wrjxLU4vglLhl
FP9jAlW0daCbWBO+wDa0/TuAiA63wepUj5pcO+wQsyvpA+2vbUd/5X53EoMO
gWqCZ2JX/7/T6Y7ziPyNaNhXrqISiNc3nA++9g9n3RVrX3X/u6bf20jexwld
EWnXtTUkFhnIRs4k+saFpYkQ0m/ZA+/RAJVjttW2u++j9lx+95zpB7llPXW4
i2CvJtIc1VCcrtIPb34TabJkuq29LXlJLvEHtHU1lKMyC4tB9plZwU/Vj8N+
ZixrfGYb9/x8anTbgLJPgKFqOEnFAoda1oJPIDrfdQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
BbR+XyXcIxL7vgWG/AoeBZidRA3dh3xu2F1/s/ZUfPOXtPnNkJSjXKtT4VbD
upgVZUkl0SY02OoWjOjNPM3s82IQXaMxlAgngzsmYetkwTEl/1MMpZTJDf56
evxYiBKRtaT8abWZ4CZVvGJHPUAwASpYJMNY7AIcKjdI6ZZ2tE3rIrrlZAo6
0At2oT51JD/YJfrKguQN1CJX5yPjuWleMRYAQO4nPtKG0uxEECWYNI1lqrO+
P0SnV3pXPabT4NSREyEJn3rxzUHDeragx2spG//dLSx10slyBjkdylTEbn8K
Jsk5i9jv6JPAZ3Y/3IA9yIwcb/ZIiPzWDy+gIKyN0Q==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FuFTKkRfXdnp9N8q0YXymeeQl72mvnvw22qWq5J+FZpeaqJk5rWZI4yQJbti
QsTuD8bDWx24hv4GPdtOpJt9PbgdQL1/xY1eJDTBO1H7e64KkYnR6GeAfeDA
RLqy7QD+fCk/OcFgdbf7qaGX2D+esfwU2x91rgj3u1eNR0ka0ks=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
R+VInBPR24WN7EU41D4GgRhf1BUCeZJ8MStB3W2yQL92r4ltx6z0qkNzgK3f
8vZ9D+DpBfUNJknkK9HYBzJ9zCxLB8S0YGMqL7/7nbJNjUqW3Udv0G6RBM/H
b5jcPXDCXxz8c6utgdDWGFhfLcumTeQyhSbEDbz+1icgVfs1ZEGwL9dctauY
Wx/RFOEcw+ZFxyC8caPLDQLn1+YOa0YnOMjyiYa7uAxYDjo17Jyav34cn7I5
6CHBSZIsxmnuiKZGm8LgfYPS9yMED81dYxaMjQe/tml5f8SkQrBYndsRK3bN
LLh7N/NE5vF8NeGGVNlECWSMpgP0jJmP26ed52bb0Cv+Ib8Gx3IFoXpbyw9v
9uly1I8COsP4rrp99dMVr7Ld3njcFF9p+IQ7Kwb0lT1j0ilrwalGavgG4AeX
d/0kVPqWTiO/iv4//tVLGCGd0BdECJE5cb2QG2Y/5bXl91G+J9xV0Vi2VPfS
+loBgTpMCZTdbTv+lmlHV+Y+bIAfNAAD


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
hlTbzxwSAdfneJte5A3G7wOMtEXdEiJqwT5T+UfsmcE6D9LQ1PbLGuqbTRGH
eyYTv8emrVkh7weRPSI5yyWACxcEFjjMUxP90JXcrWYWqKAxpPWlgzxca/fT
8VNTxWUV+s0EMhR569qSbtEV+9TxN06ToLj/kdqT3nXPfN7EIe8=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
rMuMZVnULnkweaiz6E+ilR7OAaAwilxUysM9Ax3rlz9QfRoaZtgzy+5iqvdj
kg6UFSnEFVVBzvj2W6sgJTv4be6vSSpuRlutFX6FYn61/86cWGKpXyJ3RQV1
hL2gwReAVeq+p6JFe3RQ8gSYUlA0rjZym8WYmigKFuOqkwkGcyA=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8976)
`pragma protect data_block
tTkvP35aLIZdLHbxAHQ4rTuDgVKsfTYqGR4PDTUtLrGc37fb5AzhBMYLcOhf
hRHAd+vW4LIganwXIjRSJnFOHZkLbSF6efAPoQLDMqubS9Nnipr3wVrVEVVJ
UHmhHk+xdutSotgnJIr779H2aQUoHowOHF4T3eZ5HCXi7tJXXuK4RB/vtM36
39yDDABh5htTUXR0mqSdfRRfb/DIBv2cyoG/k6f9oWJcFkqniEG7F9aZOv6W
vs4hpVSxi5SRyiLCz+gKGuZP7Gzusn3JWZA/Do938kOTu5V+5hEw36z16S6K
NOIlQf1EnO2YAb6y85vfLprN8/N2Iqb+305kpBVFuqJgTo/N5uvTmDN4YgfG
jqQiPFWvhEGmikRN9YgL3R1D8EeircAzNyAIfLAVci4b4vHuHAKp9X3QX9Aj
4U+zCSs/jNNPkWNhKcMijywGvqOPCSqdkt8bzKVHuC6LNUOTJD5g2nwOGXbc
0fLs982sdkv/jIzQB7G49ruz31sj0E33MgmX0XvOwz+FFlGcdIC9FpE6EIlP
dhgdpDhPie3V3z+92UCTk6SPGyFzlNqHbsv0pQZo0UNKZN+uvfEjbxywPONd
WPUl1rlYeKrFOCUF+hLsAovoKQ7+Um9J0VCFL/YsqYpcCykl9u+7lndmMtgV
Jnv7Ir8Syr3YSlhfUBFmpzcfWf+hLNcOhfzbDSYGy/KvceYULUNrPR4pNNsd
phzHG7uECUdFPMrZuU8bAIfTvWkmvjJ9/aagdvbPP8IH4bj7dUB6U3+A+Ebu
bv+eUJng0HAUSAtHFzgq0048kxhBwIN4BF+TbPWpzh0JT8IP+C1iEmHlV25M
1s64+ijDqLlQJhtWyW+MNiHxNVWdB4JiJx3f+CBLZMvXyQXhO0IB7ZLgXlli
TF45OqotLkM2Wa1zYvhsMfMv3s4oU+wSfN0L9DDPlY7pSR8ZEQD0MpbT+vK2
Ih3doW4/ZAQRueq55KsG1Q0vyQrQfM+0xkvpQvq3Ze/LpMC2Xg9hjOyzJmis
/WvmPrr0jRPeg4Zp8v0k+dsPm2PhC6NqG52QLJu0Y74LEDrui54bJwnIAjVO
8CD9dDxvc1AmC0KwPHBF6nT33+6jYFFjbHRP3E66Wqp4DsZ7NlFKV1yhEJM4
OTvhOASC4ujV2MLke3hSaL0KpCb7WEVTV6S2EinMRIcSRG7tRF9PG2YkavLS
T/sd0MSAHq0jDTRGr8UhJ7Ie2z8X4ZXzjQoDdsWh7oui3rJAxFE/EsjsAg76
jiEKxDNgkdQxWOdT7iL8cGPMWAgnAEat+WPeqGtHUQPCW5LVhB2qhDN/sjy+
16AL7GMXpHmNvwgetr9xRag0D4GhrLf81MPxiC0x7GsVqDM98a3uQecG+5vV
BrVHLRo9UVRNjbP+UKt+sKJDpPHVicLPbBBq//ofRRuhNm9JkdOe2hnliS5g
ZSF+F+4+3+X9Th+ZaX//bVemfq+SgXgnUap89Pr/kIEjPtvUXxGFk0WZk0S9
bWFyY4vNfkAT7tihzyr63m6i1RHv0vKMKMxb2dbvvA1Tnmhu0bhlFqEa9Vm2
Wzcnz75gqQ+lo02beRDSQdnEbMyt83ZPPYyOkHM3N6s/4e4v8tFUZcnkz1Lb
Ptk4snYeHzh7dgmwlJHOaFx4jxRPdhRUNzh7J1bQChspWtB1Cx1Zb+Whqnmn
H/QHIKoTaTPRHXU/tyL2O+7VPOM01xZu4CHRy0eF8wfRKq5Edpq0Ng7CUyJH
5uBh0Lo+ou9K+t0CixUKFSbHFqLq7+PEUPXuHy3z2L24vPu9zUWITtp8HiGz
Zgs8dVjv7IWHHcMrbRVeoXT8xN3WTkO05oJfw8urn1Ouer163M1F5IGaMwP4
SYqh9c+XySzKaw9+C6Iz/i+oukacaz0gt9RcNUF2ht/cb63k1alktIf79pCx
1W3TO8IiUc4/FX2J1sPTQVtW02iCYd6WOmVx0pluq93TqRJgwJadDg1o3nTM
+Hs3XgSAA52D3JlJOAGmXX35Hc8gfoHiobFLtat5N7n19JXw1tT2+S/pmxE/
ntc0E0z6fyIxeLm+1qtufro36GFLzibeUNshGHYIME1si36/+T/zNsGmjy5D
SAe2d1PbfmpiNCw0/+aaPW/2RhD+1LBFOqRTnYh5SoiT4BLhAlqrxCSsMXTA
Bu/wJh3c9v5imJXecWcVwqL8WO+P1Dc0OFP0ki8IjFZ9rrxuO+nSX21qGqmN
i6rrSgcaVwP+iz8oWdy8W7GBt3dGK2UI/WS0gsP45eny7v7C8MPlBvLi7kYy
oPJUv29oXPb7JTbKskAr6PyDGVDj/2McR1F1ztPzcB3KYi9MPHuELVei6NPv
fHNdCGNS5G78/fJJC3/Qd6pIQ7YR94WOzbnwQDkANlM0gTV5ce8HLiNCNfAs
8dznlosHtY4qaXc9IL3r268cF6zMl60mBR9sOx6fawRr2PyF/f9EbJ/EyRl2
owJ+KkMzCe28FLM+Xk7HznpKpRt4bh8dX8KNaFryeDXtt90iM1StTRJja4MO
t3C5SBKB+kC3ktuvJLkRci39UOFu1QMelKkvk6d072c3cf+muf3dU58kEGDQ
5cKd+pxV8IwRMv7x9BNB1r7RCtdMh3XMghjxJCLSeUyBWxQ2dcq8rQxm2VuI
ULcC71b36HGTAfcUYNQB/xyjd2uaJrQhmYICceOovXTJhFFvsqmuIbp/ozy3
xhsT99FOVjlVllqfJMBzTGplDdiGQ6H2VmS/JD2sE0sX5cJQ4YwRjxKA+TBh
zWOJvTmdI6X44cfQOwT2G1dyQ6CQWPXIr4jykCUrz+1gAVoDluX5ti/0awp+
zfhI+HkqxuqEA3SVxxT8Nh8EDnlmY6aUFp8wgzjnw1cQgKWMOVLgE3vaF0qf
BC676VGdm/aYMkhkS8oZw+5Zre73hMKYZE8W6t/0itngTSJIatIYX2lDV1Xc
ECp9Zns+DtG0QF+zqyOgMAnKCDyrQE6PjVZafmqlwLweA7s0f+FmfvE4zeZp
cxtmy9p1DZFjwpwPvoO/9abTOE9FU42bGROBLGn5N6gGFbtduQGKPHPKSnf7
0c+yyG12XlD6Sr9/GHTQb91eZnMyYOZYCjENiAAgr+jE5bsCbr9uYqxROEyZ
4j2H+vyYP/WfcqMp04e/RP+gz5QtyEYEHozdOUChn58QRlzC91IyADwq3gvA
jRjyQY10GiHWTWjv5EARQFb1JCNAJdqA/XMw2dTpwUwK6vJoUysPHpL4x9/m
YLtVZ4nCvA+fLppX1nMWmGAdXrMwdyjsKBnzZ2M7KPn8KR0T81Uh09/Z5tGQ
6cv39EPlQkBqppS04kUGoIUG/8xwxSJTBC8oI8q1ipvqM7KEZ0qnuyvdVzbs
EFysA5BurM0IXJSLs9mqR0orA+zmJtt19ufN5NbkesuLRHcVJ/3sic/b14Nh
XfVJns7RQxYA00AXEn8HvI6y7wnKP7BReMbdM589gpLdMwwE/Rs9Jqhk9sR7
jTmJMi1IrbBgxVccT3gZ+n2/NL0zWffwrqzDEgXdLAPH6fKjhVIxsvW1ngcj
O5YiYsMdLmtWYUCZ112XiWW3WqKBW6z5STEax9NbhLo76fFze5st5cP/u3HO
YzBZp4hJWw4hbXzJbdthyI6jkJwiYjBwJiziERjs9toP2KIdkrrbPePXk5HG
ZO7E9dIl4wk2d3UI30ztxuISY14iFf44JEnoUBX0mJsVGRNzcwe9ixSMNka0
IwKFoyG0/EVqsJz5ZEdS5HBp6Clp0X4HlQsJ0UVQ/BraYgFTkiMSHxKOG4pM
UD9/t6FZYXXD1m8vHxV5tpR2WFSLsduFpczr1FCyAdi8yAtaJyNxpO0fjqJJ
eclt1TGEtRK/7FuAv1p6cQaR+cyebeLxzw5LWDMxDejqMwdfawbWwDhR/Psx
SvYHw03zRnulJwLUbjK0gggQyTwt0vG5N5hOpb4/DAh0g0Xx9di0VvxO6o1g
1UFmGX4uKnTImpTNDohrLqOkW4R6duAiYL4ZpvkwpCAtLNtWg/7p9J7pPyEJ
deBazdE6/HmAVZHSLaKdDbtl4I1q2LjMDMTm9zCzrSY3OuUqfxeO1KClYCH+
asvoVCu3QDHmuxu/pTSn3T626NJ+Xeszd76j4XE1xBfx8KKTJbLXBbA3PtGP
QVAD2LT2h+I6CXwdZYa9DzE8XYT0cNypc/98rQFngD6tAAO5uLykkA49C35T
k3NRpWTd2S9qkizxBy8gVOh4q4fD9y6lu2BhWNri6cB/VCDIDqsMUXgsDWXZ
BUz7vuuofavHOaX9G6NOMNheC1T6u57cNZhuAnNv0X1wYegDr87seFWTGbNl
ImOkwgsO4a1V5GqTsUjXwOs1Qc9nRlYXlVz3W3s3EJUomOo6gaRrO/vmpiqc
GsjHqrFkY9d+bApCI5qFsvBpytmkTG+Bx9xc1YFG9XiTqj7KCv6iWUwu2fTk
JmqgW+zeALWK2SJOBw8PhOXi4QVsr26vhBOXkQMfHLZUAQuAe8lYb8Ca6h10
I8GVUWHyrkFBiZ6L4uoQsD5UZhHZpsouPh7TsmhjNIVeA7FWMF8iHK0U0AIK
hHwKvhYinaSs8BanfaKUCsLSsvSKuptlmIP0wGS4OTx0xTNuldo9AB/9To2N
s5d++M5FFkvVb1SqxDnOZ+ZedmnOti+i58T6uzMUAw/mAdptznmCmL7NJ9JH
HlNX6LfmcDVl+uYa9uQhmT7X3NYgpL5ysKuH9M4ZEn1vsFqag6jdIUOM5wkS
C1fz9xPo0KhOVrV0qlvbQZ2je/s5cM5EoYRajnchBA21q21D00EYjwNG5Z/3
1tHpJTMWHBQy+8Uiy0iDKe/GbkcVMSHZ1ovSHuk4BD1e4booYGtlG5fwnE9c
qzg+K2WtRZgtmbjTpVcDSxMpzQnD3q6yh0+myf/i/cKgKLdg/dRHQT5cGAFB
/KNAylsQO7mNfpY6Ubgj7K2J4CCNGxjgdEdO4Hp+9XZunGthqYkZ4+YSAuWO
c3rcww0CDV5z6CfDucBPqp4XZP4eimTgBXrk5ZsiDejoarF8QnLuf0Oq4x7q
SSY4SfaHqyrlCxx4yDh0hEd5AfBvPHTxk8JkoCIjQ1e1CLdyeyfUEz9r05xU
jZTnpAYF3SF00WRZ2pUGHfE7M9tx09WD9CJ7Eq+qdRnd//aiHkr356qMRWKF
Wj2KkJ8sLb5hQ+LgIcDbROTu0j/zNlUYec+N5Rz/0KfrYNibrAF8UIszAAos
6vVRikXUiaDo3orzyE+TVck+ng8RAmiclZLpHOXpB0krkO4HCTbEMPveQfG6
JVhED11y+XkAhsyhBns5eMtcg6hicJh2KSzSNu2pykDwe6upp5/XG262G+oY
rEtIj4UN5ZNgSop7T7r8eMsUm85WRrxCar8VoE3+xt7mpTSdQOinRZkjKiRU
ev65is4FxXhOT78TA7RNGAvMgrT6dopTS4OYy/uvY3wCvQ/IAlUeg4ytQiO1
I3wsVhaAD8BCXQiWbk3osdwmr4WIcdZDsEJ0UgLmU1mn9u7w/5NHJp3oOC7/
QaTthG7eUXYQi01rSWzVSb9pXsFEAmNEYp9ouaHjUEk/9zs2AW/f51eU5gf2
BNQyBj03Hl8GP1cXenZcMA0AQhuE+c38h3mPE31WLUvieUZhnYM9x5x2f5wS
/CbWbayBjYEyRebelZzDteOJYClhHjoj8YxtfYlB5hBfe32pFSgbHf9O3yMj
05uo9ndvWlAhAlxukzc7vffk0hjTwiR1hgjgAYAryNf8Wi3iMVHeSKFAeY8h
ffXuQh5R7Ji8NWMJ47JyrCLxoDdhJmwkVELOG3Lk3ebgxW2T9dzkiLXs8ob8
aFdiOvjoDLalLjLuXEohAaz5oxnnWmxwROcXfnYWuMJS0cFyDPa8RyxOhljW
hGIzEA9GgFzJt2f8of+oGEBvrfKY6509zAVbTc162uk/qphb2mty+oTWMq/L
MLJ9yyT/N6dLF+QnCQF9vuJX+b2os32+eAL14NEDXhb50E++lVZHyTPDq/uv
1hYDEFDnIVMZl34bTn0lXqCk8amBC+rCmIR9N398Kbll6KsIubpyDcc6uECw
5cCX0WdPMqIMgw6C3JfsooT19TjwdslvWAJ94zD8Zc6BIJB2uGjMDUAgfqK7
CnRYMmbCHw6m74PMsrIk7GyNoMFIWb/mZJGTdMJu3Gx7/6DRqlfQ5MtzCF//
ZeUXJTguv1X9KBEnkYkvGktrCM65ze+n5yy1N0YCiCajshmfqBb8csAyBZ4f
mE7n9bpzplkDjOPFDSb49PDMggqUi1AZ/sfiIFHGGv54GJ42753AHVIf34g+
qUCSrLOm8pwaxHOZ2CyoBBepAQ6qyqkXoCgoN9LtjiLFI07nsgo0n4/eOSUS
sHFsBlo//nYU3jLMogvOZjJJV3XybewRxda3B6bR3iELsd+24NkMR7FqEmBl
FlTLB8VN+Wo8jem6MvUgNX3cdiuh877UX4FGAYt22MNf3KBvo2xG5NCzmgv0
gz/9hJ1oVtceMAr3j0WOpN0qCSzGHuCGvtWuKva3ApXuDO92SI6RIcPkdwbF
rQB/lGvtKyOShi86Shr+FJ9Y3ivnjLOVyvVHX4N9qshjYXtcJqHKvHvmJ3Kh
Qw0VJmeS9MO6GmLMvDcw/DgABej8TomUAnwnsn8HX5W7pmicpnUPItXvEKt4
5e3aV5ZI+XrRzAAxQaYnC4mfRbfdpLRcN0+tVHw4luQka0fJCFWiinEeGWwE
k+Uip2URJxpWKGuKcW7WZg2mBYPXVQnU1mDLu2FmnvYNj9rVL4BP1RvpQ87O
JlGj1D0OiwSBinYfMr4ptat+JmA5wz1apZrEyP+YOG29QlIuoARQRLA+P7f+
CSB7zI5pTI+G70R91lWx7A3rPkftsCGDoRB0s5Ys2h6p4QnocIzZsfX60Fol
WG3DrbB/7gjV2sisq4uj8671yzVnsghFW+Mn4j5Sy/UEQFGmkBdIzF3x93eQ
AfL9/XIUDvoVDpEbOTi1sFlksHZcqhdF7Dnx2hASwPD4akCxOG7x8Xi4SO7m
75rVbGxEdvwocIi9X1CXwSuTUpdFPoeE0N3i1JYoReJf86w+mnfGhAnaJiiE
F28sFOJm6/3cQUvj8kBTXnEf2xfHBkd0o4gYraoll5/xmIPD5g4aP3IatGIy
zAc7h78WXy3y4ig9sGB/t9hAOKIZAIX91pzjDYYx8rf0ulVVVLXi2Y4PIn33
sU/lvhTafW3VGmzctp0iJxpN7cEDamAGVweWyS85bi4vuzfrlnze+QsvEzji
hJ4Y5BHbTyIt7JFcIR4AuOBc3af7TfifGK7ReuyhN/OxCaMQ86KBq7+5XYnl
Qsjrar+PZRvyySbvcRFwYupeS8d/sFvc8eS6C+Ki1h6XOR7vldymWB8lx+cv
2B+3cywph01jy9NUEBLEzUf/ORwY4kOf3YbxNwj6aTfLI3lL4lkG/CxxYXGU
t1FujUW72BzOUnvtb8IXgG84kwMmbWbwV+680aG+IAD1hKhMet5ffIULpJHf
tSKHU4dgWkAiccqq26dG1pLfc6HQiOEbDeWfa6CEM39gZ/N0pf4BYwB6SL9a
rSMfNn9xk/t7S/Bjm17QydUkbTROrLkMvWksxwWaq5UY3dLUSQfsA3XKm+wf
A3QQ8WwsjAfe+/rL++pChN3z3VJhxZetw7aIeJk9GcAjAGvpukSJunaHYqHp
/ibm3wvfQ8yfa88ZVNWBMq+tMss1BAjHJKQTrmqlRJtY6o1MdusgpbP6SMmP
WWbed+CASsLXlu/SBNMfFufvELdX7yiEfkuGXKORVWxbdL/+ishdsV/r4qkU
FMALnkMWv4GNCSoXy6UEvUQLFvmDpFzKLzRE5GMr458FFpsTqy+FDIFZHyN+
M4si1ZOOx9uNOok1yKieb7YbSdoI0b3/MBHPx6LRMrgXfvpWK14qrahgaox0
aUCNAzmzSojpg8R4xC9cKWP7fb8t27nqEZ2nlDP0c1qqPmQbHBMCrCSMyOa4
iSjC/EM2+7dvFgU7i0p8odxMeH6JOUsZPfgvEjYN9yU+GPBkCBgn3qphRW7W
CbwdlZOaGyQIH6zLYZNdhrhbils/xaZ0lX3y5BetGkrdC0u7veBULL7NA1Hx
CBHZ8c0CGhXl+4nJeAA94ww2oE/k1eGqETOlCjL7zL1XyJJtrh6y2m95kOeu
zEAE7T+DkxYhY2YHVD76P88KeA3EQqLJ4uujAr6p0iJmaHiyklVAATQa49CN
0CEt3/F0HUadeG1SHRuToFWPH2QyG9EBDJKb4t2lXA0+qqSIETivbi3uFFDy
MxspLJzqEOTYS2Voccs6FUhFfnCK6TAuBnpz3m1u4CsqO+8vmBw4h7INCvad
viTlTBbzXpbnD0qPRDrMHQ5uhw+sC5NOx+mw6WcBjvcZkDSZ6pTnAr8I48uf
+XPGQffberGvCy1q5aM1MMYOGGC74WayVgtI9i4Rip8XgB1pQXake3RzYZJX
0vRHu9AfX25s4tzDPyFYyuPezqAPEKoLxdpbeqi4NF1sNYet0Xs94QmrfOmi
IgTONHjADD2aziaLfmiJdoiFTxHwHeODotoTPnBGVwZZmYkmXqFafUeqKuor
1cP4DRtGF5JBlIZU2xTCo4FI3ySNLYFKbGpeQGqnuHESDn8ZYm4hgqFCsvE1
eX70OrA1E8NoksfPpZGam09ZDBxERUTOCL0XjO3Z9IcQv6FFqJ3Z8HmVVEDx
DnrsrgIfqPDeJHHgbqyEReWSSQwIo5Z3AEYhbKF19EfdbSurbTbimowg6BBB
kU5QU2O9Vq74bBzdBr+/Ad+dcdh412BVEQ/dJb1YHfL4cjkwnNvzeX+OMGpY
8An2oCIupJlaFfqAyif91NQgJqY++erV+crF6fNSCBx3yJUlaoA/m0P3jWiQ
RJRuNNm9QX9oyUaQmhwsAmkc+fpcGkHouHR/MYNYOnTzBVQCEeMY4flhgVQZ
cCT3AvHmPEc/h5XBR2h4mjgOls4meyre+/8Cz0cvY75sQv5zI2xsoGeiO4XO
Z5gzQ+DzmuN4mshzg8j08FbIjfTUzqc1pKT3CtHXF2Kar60WjlWNVEVw1IqO
N6j2llQi1YJwyg197on0MTPW5JzsfZ2Y2f7bvefluZawpaFSHRziio9aMaxL
ihorT300yX0aXE9lCBLXp/VF0FRU8m5u9QTr1NpQvO50yHIzrb9qOD7eRFIJ
eX9KVQiPOTwxUhrQFthNsu1x8jmWmIu9Cw5CJ4c6bny32Y72BLA3mL/SMGKY
mDL1BtvCGxDDZQkZWoJ4llPzQNrYgXoxy3jt5fU7uC4ojQCscID37Xs/uVgc
IfoGzwNsOIrfzZzSjQhvqcvq4qqX+YAemcw6OzKJjtF5W466i8DKd+NnzMe8
qsSYrttGVdeTFMTdTPcD5qAWiawRx0oDz+O+i1mD681YuLITzEMq2k60TXXP
zzrSY9f12qJIUr6OisKuvV2VqDWhJ6ySJcy0TdaIu7LXg7ww140pPSsj+fd5
6Jz2uhCaytg2LyG3bFkBbhraa1SFdHOr3Zsj8Bx8RNieTIC7BFd5pnH16ldQ
+7e+uAMhDGY9aaNzhfpJ8HrIQML6yZ90UflJytrq/HoLHfhyz2nDeCH3Jvt7
shx6G8wsH4Y87G30gtZCqWtxs1yQtDZvYVE2MpGwGzJcAmX2oJ8/rkIVDpXa
T3lOYafucbYqZf5UyzHH5gV8wUZVvSGf1GvCTcPgivsr7+j1CK/++8YfRbT7
V91ZEXsBBYjK0Mn2/A8sazpe54ln6YW2YBbYGhp2T/cdlqKvPFnTEZVP3mH+
7/LB9Cy5HU5WnRWx5Y0aRz/QJ/Zi977iDNsL/HWaw2wRBoKULQby/2IOsu9N
WORxB8Q5FVIuvOOhYHq53mOcm+3KlXdzTMDkmIQ5EOqWPzYBUnkTrK80jtHd
PJvP8SPtUWIU+wbhXnw/1F6G/2RZgYCAjG8UNd8iAMwlWXPXrDgohIJ6ALRG
w1C0Cw5Ze8uwK0RGZUxsvsGmDlo1UzsLd2VH54qHXy8KVwWF2d/J4kbBWjfy
RDSUDZ2QooBvS/unKy+Ab9rcy5uCinE1Eazgq3lXkCzP715yCTdL+Uy11cks
+WENtsWJmEnFe+2F75cXL1NVK7HrfK5uV7RJuMO7mDMdTQK/oyLQeGVzo74X
HqJb2Ar4drvVAugE3ze3dW7GVh0ASPeRRbx2ZPp+dB3/WZWC9+ZNYtuiR3la
C0PK8z80754DXf59VBakT+nCb/R2aX4zvcwEsPAdtv1ov0+pVivihtzcvRjI
AAlpUA+m2uhKHxG7A/lBXANesjsCPA2DIhvI/RJihIe6vjbtn0QQc/dIV0zm
nwa0gc7i8bv2LxQBTiLT4baIXQd8pQBU/QlvvyAP/7YAGyGcIt7nyqwtt1Tn
qGER1PePppkfsw5LoqtiVKI237quWHG2SozaJqcW8q6eBr0KfL1IdhXTpiRB
ekk2eXd02S7EonDJg7/kTS4OCN1r9PJQleYUDSKBQgN0AKRuXsKzdePC7cr6
Fo4n5p+YmqVbKLEbmuL6oHLOFr6M55TWAArxtyrilOQC4WehgkrTwOu33Qou
Tn1SFcj49m9M+SfWqGNloYvwl3PeHuKvKFeummCUmPOhNwtg+MZ8Ml2P2J6f
w03eyUEbDdDPv/Sh2JzeuGumU5yy0NGcih4HNHsgiC3wMmHUH5jFgLxJGXoo
11M45e5HXVAd9fFhuOLQxVZeDBPiLV72uQfSlu0oReDmicv0lx8ilja0bdqe
XNBTZp0whbcpBS+qMa2o2Xk55vN0UgExg74Z+7knbSws30RvfKkj4ru4VcWq
o3MsiH4fYPqkC/5nLdj738DqMikCBDMg33wWFJljj1zfRIgC14P+TPEKASgo
T9yOgsVHQuCIO5ZX4jXqdMoyENk+gxfTzbwfZ4IMTWFmUT0cbNinETKr7QHS
Vh9rd2/Z8SjGDMuhdfbK9mlQev4+nllivjkQZZlVu6WntL1NX6lUVrpGSdF2
0RmgKRztHxt6KWfN2XTVauzw1o9zlnV/Ge4GPO2VchStDfuIn637OZhnG1Su
u6H1nTNQL8udbcNcfYsv9Rh2H+dBmhU+SjhEiRhQMcpATmrwaDf+dcAu/h19
tRS1R7LSRo9+6rHgUbDYP2UrsrxR1ujFpnVmKYf9+j0Gkv4gJ6oIe+C+PBu9
S9POU9X6WAiJw8VMtXRHpaaY3ER5BwCBEE2TIP8dilK0vWuPJe092A+jJ+0X
i1p+n5b6AmSnwGwvF1KDZ8bHT3Y28gSImqy7YYwhI1KPrxWajxmuEDW6l/lV
9Hat7scMxiHjkCp1BA2hyTSs/lqmRjgvedQuhqRiiU/0qRSEln7g9pan0LKP
1xvpwVf1gbhab8AbHsHoBToHskr0oq0KF+AUeekftGPON5oWk5RmubjUR+4c
K74d4tfKjUDw8KI9Dqd2kpKY2Bs2od+urLmZg3M4A8IpHXKmxJsHT9FwML0A
2U07yv//Oov7MPv0ZK5/Bi1KTCnwWbUTjqw9ekS1Vs5MP4Lyli0cFrNO/lwT
6ZLl6hD4nXlH7anhkqoxMrcHww1tNbi2vePnBjk/cMbcUbYIHbdodNN4VtnJ
vkXtp53fnQReGitPT4X4JeCMHxBerFHzho2GJvL6/PIkHoxGqLhZ63bcn1y7
ttlVjnjjo85DWz2kpWgfT9ruJ7mPUPJJmXarZ9gbvfwYbcB/pyFFv6kwboLB
TO78z4jvXSOempro+rAD3BajuaSy7C2+zcN6y+qsZ4JmvohsxzUrPYWE/rTn
2LeanmMoM3HqtiV+8OnKuVwsuM6iSNXNM01sddUeexmi6MqPz2c+Vbaw+QhF
ofw8Z1FD82m35y+6o5EL78bleo841/88RdGlecS+eBaYjRN09gcMbQnTxhkX
5BuBaRbwKoP+L2qwdvZOTVK/oJe/U7DpPeIcYV4nNKDT1Kwcz/Zk3ShrG9tw
7tjbINq8WCJXXc7ZBdutvOzoGt97

`pragma protect end_protected
