// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
hnxrEX2BG8auRmrioY6NDH5BTAN8C1W7Pp5BmHI+G3NJ/EngkPIfjauFgkWz0sqN
ekALyxxvuUdpU3PywG7O2r/Ruhu/nBAztldUXSLxsg3lKY+6gj7xbb/23BDSWzf+
CcTqcS7I2g8zJF0FP9ueZB19v+UPfrjjZ9XMoAerVow=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 6896 )
`pragma protect data_block
G3wSVHCTWZXvVUq5xIok6ioVprt+kvIMLayhc+FECOhFCr8f6OetHiCHmP/r4a5q
fBH/4C48LtR72PRaO6A8YHemazfdzOtk77gB2dPZMoeXumiZAzD6QYfLxWJeD2z8
C/WEBS8a+xLbNlLAtSri8PDKXsi0xRtee/2eaD3OUp5og/W3bS64ir/Dp65BnGOO
Q4jzOkrT4MXooy1M4ZiYGMqgQ83nI720scHExxcSpP9Yzpr7oxG5I7YHVR6FpphB
bety/49ypXEHtKL0NgLtLmXR64F6bdGvgi2CVKKjsyqHjfqjEZiMOkzkf0qvlq3W
953h9mK65SvE9ESq5lGnZrU2vl4z00p4U7rXqVxkCF2S8JjGEvTMoTOlg0SOUbpD
5eDG9ppX7lfu7leSmYmIWdx5267jGNPvMYk/BK73ZUpVEJONgcyXOMzqEFLfJ+H4
tGx+0cVd05j6kE2oWYaEwRl6NMH1detMFdiRcVE8ZQ43t2F1j3Sq5FxGpEJCm9fI
1u+Qzuvrts0fXbBop4ETGMeq/t7kRtVn1B5IJCSPipDQ+WdxKJc1k1Dimm7zFDbv
uBObFhZ4sMpyuDhelym2/l1t2px2CBCtI+srmiVuN4+bKkrakATuzAije/Prqfvo
MAKk6S+8ybKg8QEKk60mgz1effk9soqMQxINihVouoDkkxIgz2nZpN6nPb1NOSZ3
7U9PFpyRxvkPStopJGCBskon+Twnu1lrINZxx8onwYgs5QJrZukx6rd0l0lc40vv
CY+/A3+M6RsfzhpD/dzSdRAwfkPw5IwEYk8lUwe5c5u0v9ib4AmaRBBtp/pfWUoQ
QVY1iEpnrdUwgV8rV5Keli2hDqtDWRsH/ZTRFLD7gm/Wmmy9CD5CuQzeF4eBylKu
QTps613eQyRg3nQEwmemZwASR+Sf7KDarhHGx6EemUC+pWDc61T2XLJmLXNPhKc3
GZnHFyYlmHkCCqnxGVyNk5Cr9DrBFJBgkCDoqs7NxoWww4mfbqRfL6FphyPwbXgl
ZaGGHV8suL1ydLjzbX+xNkWEaVrMKxHwxBK742yHPeBR4SzkQBLqdKUVkGpSuuxV
CVjMQkaKClozcyJkc5l1VuJUo4Bimbza2hyyoTncfb6ITx3TkHP7gX2CQOwnM5iL
AJYeKc9g3vayxs0NaZKBxTfMx9yn1qhhXFnvmoXDT5lDytq8lOONQ2vE6YXiFPzG
FGJY5cuNNi3aX0MlaqLsbPqRadlDBUGLMlVd1vNMMvK26han0ZKD+tWQu0zt7ITz
5AfxlQ83vu0VWWHACGLn95UMGXL9U5sAIZvXCbvr6RoCZBDHub+Pwzgrt5OIubT/
gWNkVy0f/tdjgoPW619b6BnZTJqeUTQUEXoqKyB8mokaLF/IgDiTdSKdgux2LmpU
l6KSc1OxmNCew2tu12xwjHyVfxzQFBBKSGhIdanrh/urP91xkZrHB9XENTH93nSB
RoEV9eKKe7EWPwYjOihrDQJVFKl1lFpvubznitPdS918YAYwoFmstHJ9WSsGViwD
Baa4oPnhGshJVpW/2DNI0UTJz9YQblDFvJYJ9sWNcm83UQoDUR3FRZCxMTVJEXHg
YGwyOcLTilyPp6H22+bkUHAy8fCvwbfDUEF+gyeU5X2I8NXZ5RU/7XuNWZfD4mZx
oMMLcpOQNRVwVozc8enWvfTH9beIez/iIX/r0gk20YlggNN4vVZNZXBHI85MYGNQ
SuSDw/8tkgt6sEaSBqV3lW0U/hQBEiEXNt7KAdj3JOge8sPAvILuHmxRG1LtoQs4
Pdb2q6hdF4sjbAc4dLBOvCTdYSCuUVG2vw3otO9DjGk2M5VIzgfHvQ2ObG8xCfUL
/9eGHANL5wt2on2PiDOk+H9Xa2/SK7wIz8kLPpKamo81cVDJD6qbw4EIVwXYFLS0
uwk6ANdegeG/5FV9e5WsAytro7K91yyIWK2WGwQIMJzPOI6kJSJH71fP2pWLhyaE
GFH+NG1sogyYhqvrC7XAjCFbbLO64JwN5IQEtSfYv41Fz6G+wpcjno86riDJG4E1
5c+pOTwIDsX6TGR5/El2wcldNWx5o9yBrK6Y4si52WnyapY8xPr3HkR9tvgn9VTU
VzlSNogR0cCJvMWIUPl9DXUOAxAMw61Le4jw0C22yx4UU9ADgBU4xDn/tJRi6w4x
DOaM4MfqGB/aV3AKoNdvKdpzqTnP46Xzo8zEZNeCtUn2Ro+lDdsMJCyXocRjZjAh
OBF/q5jERg4xQljvXGNIOI/crLREddhmg5GDlKCZh5380ZRsqYBEO0JUmtni/sQr
Aw2F+vbPyddWKOoYppmsfKoQQy/V+m8kyQjFiO5zJttpIxp8wIzHHtHtW+sXxASJ
+FsifUk+lAXvNiqhQ3daHYxZGMy0hETUyP3/z+fTxci7OKHVq6VuvHvo0c+XKbBs
TaBepLim8CSRS+XH9DhGtmzh9krJ2rs9R200uO6mv/Zt9ll943cc8KBUCveD8nlL
j/hsibFYVTQyxJz2nkNd1QVk122WFw1NpCmNbPgyDjLo2v7QnW+/eoX92S6Ey1wO
dNyTR5G+yQjeyiW38R0Skw90rIpo2+v+ePPCoQWD/VxFfVYqt5BZkLpJbFROVceH
HEdaPeqWK87J2Fp+k85CWPQFhM0NKjPFbe11IViYDhZmjp8BzAxShtR6GfhYdrld
//uG5G7dYDfF0ZERBRGMCbogT/27QG9m5tgCoFlrQikQuQ1nYQwChBsnnukFCjiD
AgJPO544UzRzBYgzJ48gj9dIhqf3bZ/dC8DdYdSYOox6D6vMQVqMDXyD54agY7vn
HY90HSNzmbm9xLpPEn97Zvk+dNt4GNJcapjCLdcbbbPcZVcSNGtkhfTD4tmp6V3s
quTcVTjNCca0XiTX43wnoRoT/+h+aMsB/Wx9SfMeE7euTDrqW0hI2Vy3AwEdd7Cw
jp53N6Med6JfF+4k/gyFJdMly3WVKW6IrHJCSHuRgIYk5zFrRU/2yD+3hpgnMUi9
5VlGrWy3kb5RRd3d+hawnaXpSOvACHlkNFz4Ux3ayuEgEswXb2hCXYYxz/Gtf2pT
lWsJtM6SgXgcdIQbG3FEKtQfwQqWdqW7PbxtZWsE9NjSLJ6xY0b2U4cf82JUQR4B
ljP3QwWO99FvMvplPuHa/ExOGQdSin84e/ZvOA5W7nL2PvSsCvFaRqjy7jzqwcWR
qk/gONhUUv2a0VrHOfYJ/uSqLZxqkkTvdJozq5SKKpqgx8Z3NhV4qejUgKer+X+7
KxzZr0LoogrhM4JrTiYmMLUgEKe9o39xmJ286wLMvq2VBEsZQ/BQKBjSkYu05VWt
/Z7NrYd3T7aZzuMMaV6NKlN6whXwmP/c+xc5gAoAmf1Lm/NvAYEI+WhYSAk+zZJk
NCNEBf0eLE01wdskdd2ujK2Qn12DgWEqpIPadwsVZ2V8YTh+QBVnoyNSeqoJH9Fl
PEEcGwG+cI+Bt1fRWyCKXDSOqCgV45OF7DB8ZLGFlmS46S75oE4eIs1hRlCu6FX0
mBAQEjyUyXLEqOfQhrXa3upqbQ1IdEYHWt9DoZn9y9Kemnuaqq7mdaxgPV5zHUjv
PLze0deOksnlEXyTEyoeF3ghYue+eAmaagZB4/8ehbyCDAxxelZ/NXzuDBSThUpv
zgvHxpkM3E5jNJvAq/80yHtpP0ntqTV2yX27yEq82gm8lECIq23dS6Puc6TpA0yu
qkjmMmISV7IjDf/mW2IYLzT0cpV1SwPGhaW97yglWAHlepm1kLOarnHJ3sDhGKbZ
j8HlpTwkU0UDENkbYI7TZd6glC6lT5jqhsAv4bXMLdWKdGtBEnuUtbpiY8r0XrsR
dITMWVAqaxGpoc3PxkNve8BeOexxL/ucz7i4dtie+7Fa7XqkKuUeHdtMMM6gFTmj
iDC24wOSCTBBPQQsrKSKbUsMz8Poa+UWe0jrcwddmikIUrnjkNYLH/Rzbdy+OFXr
qR6s5CvJQr02tN5EwIg6RzsM+h6tmqvbdxEuSJp6ZvCrpBj9N0a0dVwFXOlG3hkm
oUFvk9b48eVZniJagLSrDmwGfPUEYInsoc8Gu1CcLcc3ZL0isZAMRCbnazxD6rd9
TQHPgZL6ubLU8fKpeiJJA8QNgD+Thk2zVlNucW8pffns0X4b7X0d+YYxQjgVNg1L
8NJEHWMADSXAB2Del6pE28wm7+0xWXeLcGXwaGn8BH40QOwjkmnx0SmL0KdUxej4
7Utz6ul3zcDZshAYtnGX+dVgM+CFbTSVBEDtrhDMLcgKixmowOIC/+eMbjvjhamN
3ZZaD9n1qJBJnkv4zZkrXnv3hVIm83KQZ3o/EsYDwQSer4vuZKpa2vaZTjx4Dbdn
i3zZya34+T6VBqMa3MScvvuv0/nsGH/OGPk3TAJVAU0MHbzNk0UN+SRNfVdTItve
Ka37c89sy+IV+4kb320QpAOVBGDAdyg8NaKoDLhqD6AtbzFEMRWXgB1/WXlLpT98
Vi7bQrUyPG80IO3bUYrOD49GX3FMgCOUMgfk03hMawWYPaxhLFUk2/mRtVgVUt8j
FiQPx5+aBKW+5VO7wQvi6QUpTxTgzOIekUs244pZsogAHdHxgFRY2vCQMETIoL79
TiE48VKEjyr40Jerdsh4qZF0aiaBqNsoVLe2v4qV2xzxi/4DHEPVCpf1dgdrT9Wy
BIpFA3gEyI70mG7eyiOQlBLxoF1ryZTG9eD+MO8FDgkJJ8IeQkX5f1iRBFd5Rml/
QD8f932QNvkvvo1UPK5iF+8NCS+Frp0V04+MWUtCZ87oMmwKCyJv3Ycy0L74RXS+
chNJGZdMKqFK0zbSm7HVDnAbuI3JM9EgSTNImU+XZJ5PeZYjJrFISNzhC04/rZgm
73vKerAdVEeRyhf6pHlKpSUSuS6rJs9OltrJQLTtjHG2hKQHhe3hOzzA6PxSMpCv
+KMw7zETzDKfUAyzzTpzJVe4rgooBp2oPjwmQsb3SN+C00/yvJDEHYcNrrlRAPYT
+PTDNtNmcGF7fTSAWaQqmE6D5d7LURoJrgFhRj8S2sJb/I4IK7eUV0w+Wz3iult2
Ey7+sMLZz0uuFciTaxx+6n6CMETiwrvXpPZy0efps3Jedii0avOkmkIWNlZSUc4N
3e9bNufp0FxzxNin9JihyKv3+PVAKkVTv8b2E0su5hZCgGrOGEQgney8hLf2HXSo
9qf6+iu7LRHop7vvCG66QufFSOYFGkZGo+S+9eL9imxjQHsoMjR+XbpGx4exK5B9
MknIayJQb5v1yaWgGy5x/Cg91aQ/TYhfZJsklqB/WQR5lMSSVgwOA2I2QNnN8vRX
/LyHowaF51SIGhC57A0ZdSF1e6zk/1D3iW54zVhJlmCwCJILKFxw4tFWTIDucYJj
rBd728ctsTdMZ6Z6Sz8b1ZxQhyLGIkCxvSc4SG9WY11witzt/jr47lBaquBQMrrQ
xMxA41e+zuzAp86yKSGpWbhY3xKF+vWfn464Keb2DeDbH6oHNQo997QhFWL6D1TM
L3aZ+hEJ6zdu6RqlHT7fJ6nSg7BPGGRVETqOw/TrU7C0xxFTAvYI5pfXneXmnfrI
LcLLr+yuHk2aOX4L570Lm+n3hpRQRBHhANykMxRBncSOCQlgpkWH496m4zHVvWkr
VwmVNj6XsjUS3/1feQmFn1ETnASQ6yO7s1LPf41q46BCJ7DpKbDezywEYSn3jkZk
+FH6VlxJJKImWODMrb9Q8Oe+dBFQCIu4arh4Pu/Z8ENbbjkx4gN8VXiFgirup4if
vvy+2JuhQZuUNyTDhMr1lND6OlFSkfp85B/t6AHzQU/hwtPVxVcPuw00760/Ahf/
TlWkxoJ1n3v/UCYFULyTnvsS/Kn6qKTmRDo6xTEf+3Q55Tae8axCK+RaCgdX+Uqm
0oIheQVsq2Qc6Z/V3P56JvW81vM6Az0i7UnRSqwaKn+7ZLVj8fUmunbYB9/uT4Ak
e2RQRzpl4vBv06EQT5QT1vXZ6o4u8fc4h5mxExwM5U/d0WV4lkkIz5KkQ73OyGeA
QK/iHLlqoxbgKR7ZtX7aP6kU0OnBeCVIc20pXf9CjC/t4H3RhwMoOCe2BvXUqc3/
PLxI4Iz+helMHKhWCfyhVTQD32Sn5lPDiizq0IU/88IezIlrl75mryAviFciCqHl
HH3rn8di+1lqoh8wX1CHHtarvXwQZlZyX6xznllZ5yTTosMJxhaQAfPbyZcyiEOf
hFTg50/Ze0u1++RjlwpaUUVM+Hj4Re95Paz36iHAqKT+hbW0jEn4I4H4T47WqLTc
73USafX2sfP28U8+2JKZWozp5ug9XBNrCvFgB6MO5bD4cnJL2+7OVZblCuCc+Nio
uam/7Mb+HvOPs3PN6F/t7I+/miZkqmVYDCF3aEi0usHKPWHJ5JLi04eTVtgtWH9u
Sud5SVt2IkCyuG7DZexlDFmvRxqyyFXEU6R3QWKoz9A7Q7aGuKNXTIm3+UIRHW8e
9dqJF+NRyZyoS/KIR7R7MiV57D0UVWjhWitPgTAE0lSvvznJCHJ4/wuDJccxg6+u
NqK4AN0ccdbgcBfh/3MZAEfMB5cYqYpKyrJ2nXPf8SdA9hDTzUFm5DcNLiSiZxVE
5levyKH3mtF1wNV4PNGzgCLHPTgv+JxO/omQOrG0yi0jkpDq7ADHx7KeOCfdukTz
VEEgBzmwNXu+PYkz8HYUS+eV80F5zB+Rjm7l3Lp2ApBqHDi9GOCQ7lRqkBeVNSk9
NZJ0ZIO7b9lItpTR4ov8kKYD0KD7GRQ715OxXnI9o9AIw9BZYByxKsnHg9kOMoYP
mi3k1VNyOvkNeiojJF478NSb43viqOh5uvltx4tx/lg5gzGnS2cPjagiRMRuUl14
zhM8uGZj9hdOuEJJOHqqXo/NG/hbEmf8ID6yu1BKErN/aBD8kCbNOTzvuDzJN59u
nH5kDZ5czkROipeNxvtD1qWkMHx9LJvBURuWNlTjSXjzOmopagCGLfohJDHFq/ep
0SXuEG3U/gz5YwsGrX790uubTHYpus2fIa3RTAmKslJjWc4zqb26RUtVeVG5aC9P
X4NzZvVPilA8fox7qkpplaDEE7tX/ZIFT4AWZ3W0LKk1nX/iYb5CHrm930TXTgj7
dWqzgwg2FOGGIkOTJQPqlYFP3N62+D0pRvRNWiY5gD2NCOKvMe9AfDBkrnWnbSkX
yaxgiNnssk6Yg85xgYdGHu7VYh2daquZoUcTOOMOWI1PVk/Dy+1/OchDL2qrrGXL
/1cx80+HjIfY1SKfAdSr8CTcG63C15RbaRKXWGQeQ8ywV0MV7IYdyN9Ml9hIB0i4
/RVneShS+CBJdDX9prjrmkZtw8Q+PRgsOF5xPl6BcFgmzV06Su6Q6H5r4GTjcGn2
Cnt8K+H3hzzWsqxvQE+1Pknzfa2wLSFFQtxz+HNbZjk/LKbWWv5eVSweS+JP+aG1
UAaJ1oBwtQ1ESp4WdyZO1MF2ZY3uLHgq/LaddWwE3TCUJDc0rmjuhCAgJE721Iaz
VRDapAVrUDHGmTm17ptntIkGQb46McFlIAzogbmetcIW06O6S2pL1kqLiC2hyFD8
hJB1c46+TVnfbFatsSP26KW62Am1oS5lz//JMgnDZ87dINxhwLJwgSiJ9bLmISjb
LJz8Q4vPzgSaeNcrUdOcPaXH8ODRYQXZS0QtiCmuGEqe63XeuqxGlc67WcigSGg5
h9QvVHuNY3FqB8hdN6WwFVIkSpL9FwnY2zIaDsKHxM3+baGLkSlgsz79EkUFZ6DL
p1fEnfJkXMmifYvlDmN8hfFIknIVK51+kYPspMZuy5zQDXsSIw/reS/Y8ZRuj7OV
NJTTRiEFzmgUL7rgFkR8irEUiZVUeRy7zI6yLd/5I3xkc7c7tMXbhQuXtUri0NVT
47UyhlE3Ar2yUFJMPvV0xTuNHUhUU523UFl6oJL3/9hnMe1h8eXTDjdkp8+RprmL
o5TP9fFymjuNSS2vHNaOiZ55FPFcVPfh7IvRu/X3T3xMI49LPehDFijMPT9+BUe1
4zhoLbJxM6JqTwK2zFngpKVsQoBcPekZFvvBRUYZCgukmMhRkY1lY8mi2WCfq2sQ
8AyhxxyWD9WO2l7s3biL2a/YCHbq4kzb8sBjeUoDFQyOXC2dr3IHwT/AtIIrjK1J
2hZRr+XoJePuKo0kGmRx5VF31dd6kae4ABEVdXr8bE2byH7AWYZ0owMLfpD9CLhm
0RRIKrhO2H34kllmQxA2IcAO0GktBXXGukOBWMAJfnO5ifDB9Q+mqJIBEB0rWsVj
ucrSDgBReCCksfNWUk6OpbpfQkTIwiOFvWLmtd0V1J9yvuoZu+ShRJamvTPqkF3g
wQtd6WR017+bgKRenceSzL7JMNZW7z3zhfMIYoGR6GMv/M+RDGmPwhpotNAzxWsA
+OkXCbt5kDeE0A2vhGeT0423jdtAa0LYx1opjcuJtWefuj0hMmawjREMkfearb54
+o8TEbvesKlJJLsAdeLL3Nv0WSny6oF5Jb7qyRzHD7bxvsOzxxkb7e5Er25ccboz
hLKslE9KWsihN5jLf7kCV3Cu9KRbbezyeGmfP3lY8K9A/tKTXuqk8DZAVr70SHz0
N2DuS8YPzyjaO+9nH0bXdKKEYf2rrfPnJfhOzw8vtti6JWlogG0hjJnx/6VhVxFV
iRJirU2CodVkiYmdUc6jXpWKgxb2nXnsnCtKtCe5TmuyUIj16gJ7rEL/WXycfr+G
kWXqfFZIJILrP3u0feS6RdhQhWCqJilmx6mx+dfy3Xk/SxJIlQvvSOE8CcDk3ffl
7xtuJToK4jAlaLkNQRpuj1GaFUH9I56w2AsDBvDnYJRYhXqW7MToHgFAg8jZ9MKd
mXe+DgfPgPqb5oRjxKxtNvf8SxenTszboRRx+arKKnYnrRKGGUN3aT6StvQ6oOkb
k4JAVJoI+nNjCMim4vRKvbheGUST1ch304Mp/H85j0c9kEzrdPeVsYVuDK707lOH
MrrM7FbhZxeFEJNmwfqG1N3APjiTJK8Aul78WiR88lTVdbNzt4vkIjZsJYmZgFox
s4o72+QyyyJDGz6i2krP0+CEVN9/Ggv3mtgyI3Az/9UDpuO3xRHs6+/PBqfuyMuW
+ERrYj8To8HkX1l3kAuTYYxA1CtooeeQc9rJsfvb4fB29B2xZkopqMqGJPn2FDPm
0bywOZVXJddQTbLwMy2qwr5pFObMX6Ev8enUCQfJ174=

`pragma protect end_protected
