// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
R/Xx7TD5hcuiY/1hP+86XMapDf1vDmta1O4y10mNvrKH8ZgYOboqRsApI8CnAhBmqlM5omc0LjTW
4UTma1x19+AQkPRXX+Z0c9N4Wy3zAOIofwW77eEmNKDAuC+ahQoVMClTXv1VlCG2IEXmhEES47mX
jr/1xLyG+DCV6Fu7t4TfUuP0VCCWJcoFzjHqwSPX6K+SDkOyq9/oe1FicmgA2o2U+xy7rQqRZqkf
GdVq4W3pvqExOPrmG1khGUflv/lNrrEWVZyUvFPkeWoEdNVk8C4yG56qAYJN+ReCh7BcC2J70kgG
MvK5FwYTb4Cc3sIQ4FKAaj964QBft9q7e2ZZ4w==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 25728)
CNeChA8VKGmS8fm8RTCaAy1P9fvLw3HUbs/kEWxsl3mORh1dNtB3wKAF8Lp3xP6yKeleYYTSed1f
lgTpPohyhbYDsL29fOOrDQb5vEMTEuxOMy6Il2MdX+yGWMbtBWtd5hnOVHKzsJTUwj6TutTaGc9K
oLFYeH2d3+v1p3HooF6sjPH/v0J+9TbRjWGzzwROU/WGErKyW+KYpl/AY5iTpcHYnMTmFxznyjRA
D7z/tqAT5YRrAZc1SUBGMf79giHgQBqeHq5eBO3eAAimyWiLVm/WuOZK8hlJg1AeHOt9hIPxI/DE
mtYVQvCWREW3qfqLwR6+jofBMEEDG4WnkRrZEzI3bMd6FR1N0QfU/rNXAx3X3TE7Y8OMd57JH+xy
nQ++G4nU5QchbUR2//jLagQ+yvE7Y/ihCZ8RzUxYmqbu/VGINz9mPjUjOnjOuq2dbxiuakZRAbbd
Mu2O0cfbvA55ytjVqziK33zWwuboMwIFT2D0ya488RGIIy0PiqZ3qGhK4RwFdTbgAfD6ZuAimdoU
sIIQWzpLrrkVINxsoGleqQZuHXKusdpjRxqFBJilc/ZhL+/o/mDiFfZGl9uzoux3yLi7dHCwsyx4
lI55EUCsTMcCRdRZn4fGKK0mIoq61HeRWkIfxdcH9ybFJsw6XMENwqVTjf64If84Q8kYcFiefr8S
2LZxlXgMeXYjDm2bnl/n5Gye/ivvUAs34P8qWUo7hXZTfOZemiqRbL31A4HbNbeNI4KUQZirU1tO
0oegjbfe7SxDHW+AyfXitA+KRCV1T2iBFmelAwd5VVk3hBYapwm8b4WYOjueUntKWdH0Dam297fx
Nst84G6OLKusTue2g4I3wX42aiFALYKvP4lHFh68iyELjKm16RNyB4zsMuy2RyS2BbX8FMjRToYz
YyfyGF4Xlebq6gsUT/cEPR5XBfAEuS50+DBbDlmboYY33XRnQdY7te6im1quXuVXodDvPPCpby/H
5gid2RST0HitA4Uy3GK2iTz2KIL4b1MBgAR838j8Rno1dHDhlVduO8MarXZZNeB+D45profywRiO
9F50wU+bxFni6S2PzZQGGkvwnix6LZ6/eZiKGSnKGHb8pyUyo7llHgm6lUNSOhW6Hbrc8nBM0aZr
Va4cxnS8JqUNgMwC4i/I5fwNqDoBlmgWTUqDAwupHTMcDWbLNY+1B9sjD1ajCyphqTM992IC/kYz
MWq6fcGZpz3/Xx3B6rem8EcmpRvbSW7sQ6xv4M3moy4zbQBNbFP2wTR86TZo1g6hQ1qJq+pZCbKE
+tfRp8T3w+Pff1ENgCmX9b6knm9l49HT8wk5mCbPLppM9si5k2zv0fTn+6x3SnQnUQK7u46EQ6dh
zieEPveSjtuyGDaH4ZvogU3/4MoAfnHXJEIJw7La4SecEs1BGJCJiMpuXVYz0VfjSmZDRgSlTm48
wTEpZwKNUcz67OTbhx4P3kDuo9jznL8q8dDbUTmpmPj1SZEaKNCpyjrCAl7TuuvAsgq4xk+kwNZC
U7H8wRghCuFvc2G1XB4wFd/iOCB6CCbAvocXKuD58T0+MfgaxgvI2Krje9tkFLpCdoxgnMs1Ufpw
y/oDVgdNHFoqXlhbsEuDi1dOi5M4pA36DsY/rX6cYu1lSnAGbtTqDw5fHH3hGuuiD6DGf5BVbw4o
6AEKLniIHG8jB+b5s6QHHg12asUr9aJS1VRuqnumFI/NmzytraPfxVTZ7H0uGRCKTwMyNcIkYupn
gx2+hCUtBCafIvlxhoQ3kx0jNHJIqEoAqOFwnXtBsTmsOfLgjGMOlqu1JfDr/VS57bOw4kYMC4uE
stDD4CJ5xR3D308Ymyoj419/+KvInUsc7oolrVqLhyEMeA+UPrCNu9Ni2SqrC0E/xpJwS++PXV76
C4wJ3MbarGKqSFiQ+COF6iN3+rcz4zUhSNn0A2RJLz/f0vGKTPuGTql1JAJ/up0SRxpqMSudeEYf
GU/iiBHkJuGpdOXu5vE12UX89AjQDymcvUeQaM0NByw6pl9BGhCwaDr7FJHo/mQ3UUkS7xceEKnA
4UgPQTqoh/E6z6BB1jO5WveJ/aJr2k9Gw+d9l9ZoNAauHEmMJIsX3HKo8MuMky6G8kKMcxmXUBNW
gMPIOPn65Acs28s3mpBQ6SIyQ1P4OaHnP86t4LjyEn7IWVTRnAfAxK/wvagYN0vKjtuXAX0Qwjc6
svp7rX1e6diahxAPq2CG/GAd5S2Syxtk7QaYDQ+8Hk5gzXNA4K+BV60MkeoY4bLkSVDY0+HRDeh5
3X3fOop0Xoqf6Bcd7eKK7msA+gBCOTbDAK6Ru20Dpu9Qtm/sasF/R30xVm3GAeu7QL1nZAfL8F0V
YlAu2XIIWYR2t1AQFyg/2eeRxWlGgFSshcRl0qPT4hR9pOjR/x0VKNYG+JYll/RiC9NWtu94x1/k
KuvKAIYpDlLOeuJOtecDQni5zddg4kcMe9sBvb1lzqh2tT8teNWeHUHqadolm+6nOCooKNrkwMdZ
vFvCYWFv+ZWJ/9XcuyDDWspPytNBgfwlbRNsQdUUuLCuVdfmWy2wAg9l3AK1ryY1h+CWyrZKjik2
cBGaPWekisuzmu08ApIneGC+Dm36szJKJ5msjbcZpd88yq5DemkzjP7g2TrRZvTqdNhllkfUWH7A
6mvfp5Z3dhousEybvldoZQrv7YeOjAnrIBY4/0YOqtP3r32g3WcTmZpyWOfg4oLkPyFnLU4Me4AQ
RkvcA2xzc9Pws7A7jcHfu721qhOJkGRpqle2dQoKoKSc9uR1oxNOJhaLNk0GaneyQAQ5Auhy+Xu+
uAnayM3VuIDmVJ4s8C7z6mjohKHoqRAVtMORhJ2Ht/4iT7u/7UecGK0PWqk1rkJQhOiLwdj1Pmny
6nPOzTY4Ruax4d6dALNV9wlP9FjTuNnGLCvqmrMzTH5LNddT2z3T41kvbPSArQj+iZGNSstbUbC9
6aGXCHT59y/Q+E3AzUGac3PTpixSoPVsUBlXT11GTIflKUUgBwWjP71NBugYhFKG+I7lW/PjmMB9
+vjAh16zyb65h6zgGwJsQZo8jKtwpXZHI1VcPh/oORJXUd5LzAKfS3+zyCB/C7/ovId4lEn0ZmaW
YrApBF4BTW4GE5SxdDAIL2yF+5KVAa4UFdmsGBewQ9P6UPZQ3bROyp2sdofYS4V21vWbp1EcLYuJ
4Fxh51/j7V5HDCIce6d2cNnTNH5AylkpVSpowiOch3fez71oyXsinJxyNH8OjG80dJ8UQMwYdnvA
NH48MXbfVMbF5H5Iov4y9G/X+Br6coa6CN+L9g1yVwagQ4INSO889UbUGwf6bGhvZdMMGRnRjCaA
hsUl3qbcbYQLCCDYW4yKWnyD4/yW+0z3h9S0TtM5FvpJCK3PUFSJ+E2LA1BWR4wfL32mGMXojkLC
dKCYn/Yl7b0FFeDLihMDQauz7AC9FWQBCR0l0/mXmUDrjQQBdIlKvFvY8OR5nYG4Wme0qEslIzAY
F7iC/D78TgWnpKQIlD/xL5goNvoWM0h3CrNF7boAqMNz4QiKpqaGz6G+Bj2scMIY5VXhJZMZ6fyd
8TDL+VmN6pamtXWle0HHdLa2YVx5Fh036hQkfZRaECSLYNR9TXUuqphkgR+uOIa2ub8PvnpV3HuH
ynm/ViYntvden4How7jJTr1QwmoIljPsejxA0s1ODuCoDc9WWm8dv8pRijYP1fuIvzaNwFlhES1r
PQhQTzVpWU69mcu9QV4RtyHEnbRJNztubsjoBfqALJeKsHylFwxtnLiXm5fzmKkto87uSLpqrcno
N1ctudLwsZmEpQlakKFmxzWgxFQZTB/od19ed+Y5WJ9ep1tUgwb4pViyhheoa7LpmMqgXZgc5FAH
Ena5VZFnC0vDyB07qtJ9by3C4BBXgP+74FQoRM38QplVLOcPrfHSI72woPWlwYeIPGem4FFRB/++
6PRszdix1NLu9ymYx22FidQW53fYBl28Y0GsoANQHDO4V6FsPUPzUCtDtyyFAV2Uqkd25xEP0oCE
Ex/R98mgCKbsSNZBdtaFQBrBK8SR5mxPvypOJ9b9eFD1FFERRK2gdH5AaR8kHE2HRQeEotQhMtaH
A3QcS/WzhRQnF3WzlkWLxIP9HDzPunv2HlQEMBJUWlkRgrcgQKOe8OMrQyDAukl9ZzCqU/Qkawht
J/ZNpPNlw35PWbz62tP7gtE1BpR/Z9OD+bV42HdzFNMP2QqB+H6kD67DcBFsy/NOn7sabJYhY4nj
mXtUwnEc2RkCVTsJEm93PYjChiaLeiO+FRRT/U4P0M6ih8MBMk/FfyRS6l4M0a5j/lVwFM9JtQHY
bsK6BU2zYqA0eQVokodD/vyiVjTzJkUSylsHi+e+3lEfLcXGYLcT/19m393o95TPpTp7SATjFBYt
OvheV/LxREjQoJyzjRuwnqXvK9Od53tLucgRp17TjF6Wis2lngfo+78ICMc6VVNCOYxDcrZIlM9v
/2aC8qJ0KjLhweT8zfx5aQDEKQYPLws2dXmgAIz1+4cS9eSJJaMXV+2t7qi0X2uBE9i7WKNxshpd
QeWFMVNYOfscoZKOa9HEcipNe2s3sAMIOS47rJyZCvYnPE0uFe8L/d9iXQxmPpKS1qxbkOlht70D
C5+3SxzExycVHKJiNKl+ESnnjIjI4X2iTRhn0wjvUt97pzWnYTBqn6SiOsNeyvFbVebRkFvsmJD5
y4TwUYEsBparAPqJbQQWVtDir/tCpVdFkQMrLZ90YSOonuhGVKFTrSJoSAhandq4BzAYZtIyMI9t
OcTQd/DSrj1kCufU5CIBkUQyvGj9hyTxOQfJwtohmZ90Plsj5AnKZQJiC29JrsGWZgmek5XzEu9M
8KMwIG1WU2106kTrRuvkhoBB2NgUN6E6kWnPuU0Sc7NaARG/y6bczUt2bAqXs/WhXbISF4+D+VdI
l441hJUJfJbsB5s5/8YSJTMORQB8Vzc2Shlbjavid8EuJDgYlcYcBE0f+ApBIG6/0g+x6RVt1rSB
yj4yd8+kMneSrTPpI+CauT6L2KUYn4cIBUBFlEC5JLieHA1RyxmpnXybXtQm/qqf+hcyokO8dTNC
TgatebczqxYC6n+MQjBLGJIiD+yhQQ/HB/642dbMTPXTyhEntPoDUVU6YbHO+yYHMyn23E14y3Ro
eSpu7M4Gc7A5b0/qG4Ieivj+MLxjUwELZxG+NQeRML9kuj/A3fXbcaeXpPbv5saLxxuk/asKho6F
rbpOxC1Zksygf6kgeL5G93hCLrk92GbbOp9NStncP1++AebFjcCiP/Jj3vU2xE+TKseZD9wwzNXL
AQX+q99tofCZ5JDzhhfEnEo3VDSV7tTmMVIFm0BwFhRF40FdCNtfgFgc1Q/xldWMP9wj8Wr7Vz72
J3zHOIq/PShenPuJQqgcZrOsd4+0KM2dP2MXj+QthMDxLccO/Puxo+4DCJVAnGWSZHQxLWkW1FGb
9IDrNPIEzD1sFLC3/NQbEUTAvVm9GkLWfpBCY8Ykg0ahenJX3oodWnu47kzhFZtOgnKMHGGz/mXp
NXijdVvg+jTVd3WjAQcb5KEcreTrgjrjqWZ8ZeP8yGqStuhZrsQi+4gVXoXlWh3qvs2FGA0bN6W7
gBXw5VqzAmIgFGS4agP8ggS74O5Eo+JUEzkjs7w7WyGjPElEiSS2jto4YXLkT9VZ2+7+D0Wom0fG
304bRFeQU4EZ2imx5tqUvc+gmLXPPpZcOU1pKJyIdG9b5wdxhDAOAmzWseVO1w7SsKyUbIZUO8fX
s33s5ZTx0vIuhFvYkp50eUtJFQ0SLTqQMbun/7JxaXyupENMfOU+iWrTKJMfIouX5yLXxkGfsuJI
QablgxJ9IiggKJyGKsRFr/FK+l0fuOjbtjsZnv1Zypzd4+31NNIemxzd3HiKPYs/kAdQl94gZSXJ
HH1XOTOV//DTN3pgwLlwIgyYTDcPuWEXNg6m5MpbJCCN5+TQMXsdA4uJyxRgeAU9XtJyG79XmW/w
+TPnxgmpPXppoNe9Z4607x3iTYGeDYfKX1OoqLRbc4AGqAhfGPJZkJP53xzo+4H+MXq0jnxz5yrX
gQLljvn+nPGi/fefwvx0CBETyvXTeKra6p/fJ4js1X9cUhNb7Cyc+Hn7zCPW7SORwQWOoe5D/lAX
HFXyvLg6CRePNgSph5k7NaE6faIXuJ2MNBO4Igo4ae1f9dM3cyhwScpchrrE211Ln+HJ8oSqBiyl
pZiE2TxBK6UnLhHixDjIMwfzgpl+dpdOHVj3r3rMU/8mJ2jzZytybG5GNM7OlTJlyo3t0DGnC9uT
EWdKzawqXJNz83xDQh8N9iSfGb+UK9e3SCWucrV6LQ3C2Zwn1egWS+IdwXuVhix3xgyhfvLSUpB5
tz0JklQjBc+r63tvYbVzC3bnLnGU6kXcmiS8iLVIdeTj15PQqWpmrhUCVERP6PCxeu+YzAzLaOKy
SrJxrh/UpOJWj892lEXrRczN0kqiENgeYnXfVdsB8Oddc9SqvhpnBb44KbW5hEKx/NxnmSA5EaMj
uPrUpZdRgziqWUU4VYUDsk5uHBsXuGmudqftECc8pCBWdaz24onj19/u+LFUMHP3zn2uvNSiZtA9
PnRj5beQr1dmorkrg+xKklnL0Xg0GM1howlM4BZpeQlD2Ulqj9zeNYdxPyE5UuA56Ng3lvaeNvyV
Yr1Tp/gnv2w458O6gxqXaaQkNezPGQKo8nOq+wu895HwDBtMr6eLdxHc7OYaVRhyu878Y+t5MRRG
gjbkQM4fS6sJ9aNcGs7ZeeIcDVNtXu/LLjn2CiYcLn/JNw2Tt0jlb6qRJjuIN11rQqcCTdUWqVR/
bx2p8wndiOywcGTTDnbUQ5QETknvzqNZ1K4B4zx1J0NLTbuqSdo/tsDeIoV9u0chTFBAm19uGt5a
GSh37YxKs9540PDUPgL4/fXiAtyUQOxo1x1uFl/S/LMCMUJ4w+Mfz6pyXVi02ZHl5Md+Qb+6zRgt
VffB54Rl0CgVDIXdkgNDtPooDzbqDVlsHAEShAl8zhe9tM9AoYg8Wr9wCQ4Dnxt58N129nTDqoem
ABhPmJGzkmctE4lAOr3cEk1zR4WvoGS4yvl3gN5KPanARnGKYgZ98JHJCmbUP+GoRAI1Be5SDqKC
pOqAyDuNjY+ka3FvAV88dOUfvzkjmDtbgBd6AwMza6LjgxEsUiYrorniTMiA4WJUXMgmW5X6mPxJ
Fo0WJbCbqw2Ngm7WoUoMcC3Z4V9iz+bW3qS1Btqkg4r4CwLEV/KRhxUj1/yIpBvH0Fal+CR2y6iO
8YEk8/wP/VIuogOQKollxwxtejbQx+5ZM94YNO4+AWnGdYYx3lphM21uh0abJ38dNeKo3Mk0iBPh
96/cr15Ducv91E5FVtnWU4z/jPUbKCDTQRZiSdrYwcSHQRD7XOdCoVilv08WK8Rh3uLYn5kwaWRR
wQbAJ4WISJRM8Y5AFnMfD8XL34B9iYga2oQyDdO1DEkolQH0DA/xFiH7Hlck9VM9dBDCUeZLNO8k
KtcL4kp4iZ8SAzB+Qr13YYYK70sCMt9j4LFuMYaipn+wQPydg/NGZjTweT4ZOf8LXtJx21xa5xKS
Jqp6PtK8i+fU42/Y684nRASqLpwZ3vSued7C+DPv5VfJbfRCMRE24jcj6pee1duN8dNPDumeasGt
uwY9hOcs+U2O46GBE+PYcbYLeD+Kuy9FJcqbzkeYToCFwlFofZjTcuPODrJu4aW9zZC75ijDpG29
NP9RHViBxbdyNRA9lLtyrNDMM8xy806fKi9BxyXipCPsVBR6+ldLXPGAcuM+If/9uOPgLGVScy+d
XbDyF3KOkcakvmXiwJkfz/URv9xIRTZcEfTKC9ySe57ZX9kL3SQp92iyCNaleHGDlEgg7fsqItRi
1mHazSKcdQF+gea6C42C7i4us0fYsxPcHGOrxDXZjUcG5VOZBfUSZdmbsRvlMCSmv12JkvUOyL7F
tYrvVMTU058v6DeS7/DrpvJC8Vd+QFT4LMs1wf6WTUUQlJzOI9QVIrUAPn+mNggvG8XSRYVF6TCB
3xk/98/LUM83MgibkJKXryZDANcsIsbNwIuRh4U5l4mqQFSHGzWRpGEQwUQz/VSnBEZ4g9mj0ksi
UleQQhsGKnkU1iK1stZiT/WZaU7ADX9BP1qTKodfTlVD6t9yS/9sS2PkiXeO1nEDfLyYYLitgGU7
nPXGbN3ako7a+U/aKB6uelZpEDWufVGRhic+5aADrja6I3mpf17pUWszlvPvmoqTta9VzXlF3Zyc
azuqGYe/j9Ax2pfDTP1qla/lwqxGKbDQvbhliM10nMvsGyEckgpSS7IC5pSE3aEc8eN0q/3oiT2X
n4nEsizPod+sgptYbsuL0GQvIYymz7k2N0RsAWJD5hQPl6ATqlY2QOjKHnZJBCFow9OLy5Wum07v
1+iU4ihtm7nI8bqP0Hiup2eSJ14a/JeTM+nh/gbetQKMOuJ72ryr+kHpw8UdFcCfV/aGWU2VGz8Z
EsihOIuU/OFGtGomy/Sc1/kqfVKMOp2IwFuUl3CNH+IfNj3VIJTg4c5SH2u3V/gPjRiZKbxI4z4y
lygGsYulNePuU8N5qP84VFrIwyle6n+/+Vu01ZzZLgaCdp74wfV6NI0dVMFTVPpO/FJxDLSQSBsK
trgnKBro1YAc/4o3YonMFguR6sU6Yx9hqN9P/K6pWKUSb2Qnv2RL+UD5+cLErG6I5Eq9qeLZOZWv
B/rcqQK70PhqATvHHCheWJBVY1U7uQ0vdBaweZ/tGmreYJPH2S4gPzu1R7aMMRGomsfM1peHdlY6
WW+FUGEwgY1qH7/X/8xsJTzypPrGVBKd1CzmIt4AP/UXchndcIAxIy9Xmo1GTXmi6H6tQA4vTCN8
C1lCihdrj4CYGiWF9j/MA8XVMxKPwb3RDFPeG7F/TtEkYvlm4zC5s4GQHMws7/2m4DA69ah3YLlK
utvIQXQR+oZ2o+prqfXpNSgrd2QzF14+S/X8MorUlGoNHP5AGLpiyD6TD7/uaPt17XeX2BX6mZyR
fmacgHp1x7et8DRHMiCkP8guACgEckARs8IWSEI/RLNt025UpJVUxdyiTZJXU2bc7CSiUwPUacce
6vrtLUcwTkQFESRw45kuVtGLBQ/Y5i9afybXBkwMEa/VmKujVSoEVWBQ5LiPAeKx465ZOwpVpjqz
4Yw745LuMDEJv24sM9u20lKgVSAt6iOrdfZm9YvWx/mFVMwCxZ7xs9Op15qAgVvtlPNRIWmq4cPQ
XMlRD+GT3i5E4SOTxG1F7lyyINgUitM22UsUOJtrByFXH8eh4Tg5FDqnGuj4hrCkDwj1jYuXWnys
fzjD2P3MGmVk4E5E5AlKYDVkQKEYT3l2kSv/QOP4uY4T5gGbaycenmvgeKFDRz5+E+mTatS/BrQY
f+uGKwoWJc29N+JScl6d5Iqdnhth9hWbqvVQSuZSxL2U1vw9PpUB+Mrjzsq59ksk4aZ5twz4Ya25
CEJJRpDLY8i3jwP0CtOORkjFxp9DiLuHZLklSV69Bp7D9xERm2zpARPqKsHyHy5Ypq8vq/SwKt5x
ZYOaa4MEtretHxlvhTZ3FxJa179veoVlu2bpXN+i9VKGTiOOiBMq2EuBqnps5vGMDTTwbL8Y1XMU
QuIlKUXBtXECszWtLIK2u1E63Rkim3c0mzYHLYWaSl7d/YZK8nCmi9BNBAKml9JEgxUeLgvdQ2RS
Gj0gDqFL8tN2x+290tdhGVlKzEPK5dlIIKP5JC4TokXHzPCSHoTJyw8PU74dM5V0C1kTZEjm1Zaj
Xabw4GPRh09naCUro6ELU3JqPdP70V/olW2+h61nJfgJdPoqWef8mnOXPOfvOlxyauEzzaYFOgtT
AekFXULLNYnnDX7Z/qU4qA9UuSXFGY60oqnVIhL7mKSX0I65PP1WIREkAoOFYwg4J95iRFZlHlfm
bsCBJ1smplmIzNUSrr+o/M1ZV9eOj5SyLnI0ZwNq7gr42AKurzyEdQXlMFHQ/Eso/TPoJrP5odGL
7mioUUKaUN45S7MH8Q9OgVZLn+UWlJJZVTdyiJ13by6qkVjwh6Hgnd2GYAByxCjj8GOm1xI47ZsH
gnqNpo9IEPavb15VlPox/bC40/YbNHGN0Rc8AmJG8Yt1Mz2sR3VmPi2UzNGg3mziKEsmvj7bPzJD
a7pGWXxF9TYJ7kl0lmg61fhIckItVJY3gaGXOqu6a+56iklwSGWRIr4itbKgZTYgWrjLn3kYjTnc
+IaJ/EkUZh/yXAJauWd3let9JVtqhIdndlvh/9c4EX/661Oi0WBeQI6nvPZoepbidWYdqkur1kko
uInaewC41PRzBkfStgCSwXHsdEiJAaXxJgBIRyMDqR0zGOL11BUK9RyTVWJ5UjLkg11b78/xl2gE
QtEkLDFwQyC5++r9u7OJ0xE4wPuR8OLTwiv3dik81NSBJIvKwM782tLCWD4kG2SnBX8uiV51+Tpp
oig3wspsfYiUThh3Hv2jl26eVTaEqcr3+FqXRGmrW/7clA3YQAkcQXTlHosM50tHN/QrPC3ao+r0
WpaXnvh7IceCjx212gNQEj5VZRyhZs1URVJSsKQTtUCe11N8sQcFNPWqkc7RxGqkXrlGOveivZ+3
Oa2Q50jx2tD+gyaeQBLtVc3UHujHUi5fq+QY4NfcUDII9vdrO9cfI4C/nFTkMCypCPKwW0wBZku1
YqX/LlYufwRgrPX0QmAUHYP4mF5sgn0xkhsTC6wQ5z/sk6SeVBeYiEXjg4uHtGGZ09J/zG824UXS
gRwXWs/8oTg/b3pP/ySJatSXHY23UQxUZvhyLcCE9EO1KqLw2N7rtEIENKZCBG/+NabhGK+0mV7h
8OqPVajGrFBpAadjlLVVXAHa++8HAwebWVWG4u9tEf6LgBCWK2J9EOASKv0er+mQzbo5szTlRnTp
Fgr7fkEH3UGTwYe+S2Egzyczp6rPb36C5m1VWxhIBZVUkYu3Z3Mf5pLTD0cZZhl+UEckX8tBnB15
BO46e6EYIa1XjWD/iyOjjSnhgbUh/gGxLzmKdFw4Vm9psshE02YR+wV26thvffmOUGe0AhHxQKRJ
MpYdzwhafM2TYZI5s+jGE24Li9PakKwP5vrNhHBhAKDweRpis6rrusH0tmXlW/+UgER4Nheuw/ad
lzWVKqTyRj9qKEWn9jM6xc85ULUC1FgtvhEeaOg+h4QE3Gecogy0/uJU+HSlW506DxPP+1tePJvf
bm5lYK/YXejSJ3m/AybhrDgSk2GcyFyvfv4mI8wBEAYlcMHU5f2h318FdHoglMLJ1WC1hKEv2sf8
NWc/TyGLD3VQIZcWGSKfiVbnuzURuBojCSumSOY1dZoF5tfW85YvicduArao0x7kDLseTge9uhBU
+kw9FRA4Qj67UIYjWuxBhvZduIm4FE5F4QNSGf2vdPNfgj6mbcrLcHfBkzcfXa9LCSoyGE8eQAi7
0PHyF6Vm4m68+0mXa/QjSSOxhG/LBCq1zrxc+L1d3gsDOByHzdEZ9ZzGrx3YOkCYe695wLLn/bJW
5E41Jjipnb/RAZ4AOwNKRBwkWLGjSmvONQmqngGQjHv7g8pPZ3Mscg/c564FACvMi0jaJlIc7/8i
w+YizeQfdN7st3hmj3G36QgrCVQ3Waqj+w5MqKAHUIGXa0VDj+/rtz/LYbqzu7kdSGJs4+2xeG8i
Su+GTAVCVtEFh7XzwdMhpN1OttCJ6wbBPAMLLbCmF8OXBPVZP1qAFGz0ogXat/INQi7vhG0QvVQN
7Ai5/vTWzqU4MhLLKtdofCpBin/6S8wdZRlBdDO2KrPQ418Q8klbsLzXTxJWXSYt51mvzIznBV0Q
Fi9gYiXh6oA6kCQZGmsySbYNHIp31W3WWZQuazWNvtpAicUKZVyZ+6EnQRtnpQN4EUz0Bo4j6tLE
JklmAHVGi+2U3EZhKJPT6iTGubHzMtMSciLKVZ4NyFqEsLqb+mb/YBNr2XEoFd5EGrzHlLav1ZJE
vSxJBmUGG8f967c1AezdrvqTLszZHe2tWYbL39+T9f8BrcpSAGLy9EwGMq2uxK6ZEGEOpjpDSkcs
xM3HT7GhXl3R++vbnzfxTi0nvDcNCiTnfYGio+9hkLoUKRfnig4LpdFP5qMmmnnOSPgtwwcXSszT
DnaTx1uv0CGqDGNQkkynuWYSPP1bQs+dnRXuop70YWJPSEGGoDOm7BlnH77rUDTd1Qceatt/h7E2
9HmlEDVb5wUgjYkC8VC24+zbszqB+QraLHSXdsOu/bs0LsPT3caynoucRylS85vCp9FxvfXjphjJ
ug0UzWNGWKhVglyrDILuQoyAsdYVLZXZVJvRC2pOqHgKtVr7uXPw+UmglHZpCyHoGaLoPQQNVaoF
0vPNi0bdV7519mK/f1duPNt8O3Aw6f064GRw3FN4vVE1kMfOd62qym6Xxplpx4Sz62S8qPSlPqW9
91Nzj5Fvj1R+zGKYid5FvjYIgAFRkpLIZQIYAn7ypy6+3pncvB8zuzZ1xq/IWYMNJeq+Du5QG4JP
1ydFnhr0quvH2R0NjAhpkS8vN5/k9cBod8KOtVHJY2Rv+WzjetyVaka+AnazqRgGlqv3P/JZwIno
LY58p42hJKXM0/o400PpcXWsff4/XH18HberF+5b0oLmHQZ5a5923KPqXT6dKl9chnTRO2nKE4Pa
xLZzoKaFPr3fx120VXsD6yMZmsD1wrp1iBl5N7TZ1jqalJVFbWDzpodfI2dGGSJCWoKXrL2tF4iV
8jhuA6MFSq1rZC7HdBZC5CoPYmGf23kXjMPo2HfsQV0H5d9ubefgoxecv85fBt6tGlItHeev5G/M
0NCEi0IQ8zv9EwJg40sU5AK7KfT3QjjSuonDkUcwxcWZtYQszHel1EEgEu4Irb1HttrymqEr/8iI
lMjNFVK91zKEWBVZv62HjQidFFUQYlDxZFQ4Nr2jUg8Oei3SAeq6W2yKOOJlNLwd4fXDl8Plrc++
1Xd6nV+pJ0RhxaVLSYMZeZ/ybUK3VYgpjQzg52V/5dbDcmRXq+4KLCPTpDRi5mHKFiIGEEgd88j0
XblW8EPK9fmG7WyieHyq8iFSD+R7wVbiQ4s5g5SQTIxXfo7nva/iUa4IVmgJzLRX7XA3a/RbkXcF
pNo8n1dCXczXeHRh6L7Hn0L0YI9MG8rSOlVPWbzSSkFKtFDY8TzhdRboChZKYJZ/SKJDGVzsgmMU
yQkmKxKGVUBNAP/PWTYOPghRldQVSpBC4pB9Lpht1Nx/Eh/ckFCiN4oTUlTwGQYGwVna/5b+daaw
oGv1aHFAbN2tMrMmCdRfz5E4nzRPQIGfcBXsT7pEywpAYG3PxPzbQKvLgC+cBlsP5r/GsLHdpGFp
9P5j7ND42vBSajvm7J9bJAt6Z5OA0YjYvqg4JEeAg+IEkwDLIznv9KFOhuLSYuqROQ9S4XUM//C0
zyxuOnVP29Lp4AdLKHLfSCu9O2XJfW5FibyWVxjKv5QNzhPqoiUPhjB0OJ5AUV6Tg2d7R9C6wDPI
7BvAJi92lJ1DUdMnTHj/WGNBKkzZK2aSmqWvmo3Ms5p0tG1DpsK4DPAg3fyBoxW0pjJdnBn+svw1
1wSCKen26T8RjGd/l84dsnQV3AAa1U8Ehe+lev5puysiP4hpg+TUNrwG+VEjRMCa+8UjWlvgDT+I
Sr3DOFp23fzaAzcFg0zPneT46YdvKG8TosSdprKXH2oKmv92Ikz9v7iS/C85qihK0WjevUB0pqsm
BTkX/VgH3486PTzG4P2fsY/J/X0Nhs4W/hAYGBUPMVnWY6Cx95PjEaoShulJXfFg3UyZb0pPe+nt
Pt5jpSz5ps89OQ2DKqXtEf4aaKvDq27lcMnB162ysNkzqAUpfSFW9mlimHc/4fd0ShsjoqebSLQF
C3Z0Zv3RA9r535E2Oj6ssLNP3c/WXmCR1t499hEv4X3ZVianMyS/uFuXXdLy5XQYg2Yi2FL9kKXz
25ARDFmaRoajMG454YNsqVQmOS+OIOGj4FStM2bVrsRFXZdhTrCq7PtoV0RKdbO0UKrov63CaObO
KwIniWK7aToR9CC6qpuUQlNfpsF9YuWsV1HCTrXYpDh3x+4NPeiVSKcNgZ887rbJU9B085jdvNYr
NORmmv/m74vJ/QZ787cIaGnaEFaRThZCS+f1rpR+RQkaK2kv7RTHCwPmRNptziIhwdJ0VJIrNRrW
NieI5ZTCYuOqfZ/NzzuNZNbM+ice5ln0LXoIwi5WwG8gyZ1EO6vu8Z2whTJQ/snyO/Nyo4J/06CP
G10huXLiqARca0e5gEdDQp+mUI233MNU3LE3gpKTr5u3SfStfMqm+qWdTRJCCfhR+3dsw3nbhefH
7hDHHv9d+y4qJQpEZq1ehPbk09Z5+tDUT5525zifVdolIvaXYMQMnMnS/VLg6VLyjuucukpxA9vB
/0iuR45JUQgLrC4Z+hRyeiSAcKgShLQ6VzW9TubNFBEgfg/LrmJmel/keUsypaB2iYpVLe2veYX6
v4M5UQlxbTvXNH1vy4yyFH/h8vPDoc+OsO1LbiNVKYbQTIK0Jyl1O7YKFnylhvNvNC+X0STsTaNm
AekRTLzWerUl1xhWYfrc/8GB1ZBOdNwaX2efpIczEARJcLG+zxOiROsW7IuAZbrITvWMWELQzNYy
w3rPuEsjfF1hDKw/SyZU86+qLeC5fd5Ne8RqzRJGr93WYRdSPvOZc2cGFd6xFntQiZBSlj8BSskb
SH2/S03McVwEahQNQ+Zr+DZBoeJ0d53VRpDXo/DWIBuT46yyoTVCqyVG9IwPKAYvHKfPg05Nmh3i
QRfAgLzCfYFM9I7bHrnkIyOA601mc1UKGx5OequSJqffvLo36Wqk37qMRoh6Rfa961a3wuPh+KKd
hV2xysvVimI8X3t8YgRqOOK/codlpaq+0Z7Rapw1mM2FIOJfN6nn6C/TlKKxYNjBXpdpPeP28a92
YxcwoIIco0Z7P9kUp6j635aBiFoDZVi7gZCJKdSxVy1iE49zYHV7RzTUKxT07IcQ6Ygd0lJ2F5V6
SB2R/jPJA+WJXy0PDxgI8YjTN+4uuBL7J6qfZYgwKnCB7RL2fhx7fa3qaJHICQ//a6VGu793DrXD
yOTNZA08PiEjBiHXTfyoc69Gn4DvVvJ6jPSDHz2PNOknHPZtJHOdqaEkit54Q1O2OGOASr0IWXU9
Zk2DT3g9sdm+kKY/UakJIZHHPKSFBzBHyCiq9bMdM3VLXpnsAYqT/xrNeNMI9emudiGrCP8m9l/4
D5M7GmJrgB/vtdzE4SmHuI7em4Qe7h/gSNOiaU3lpkmy0Fk4g3emVfGEUr60vD1Gcg5RcosiW1y4
C9wJnKKatVR1neqUmGD0tt6cy8fKoJglbB9v9pb8PsJlSGpITJzl9uAS3JJ/y6FXp9Lt+fJgmAjA
ZGHBlh6i9SZiqOuVOh5rWwo7YRlpF5bUUxXBvEMx5Ic9iUtg0PoE18KmDPQ+KUjB6aTp/oJKiA6X
e0991E+6MOknyERqecyHN8P273UMCqlC99suat+9P4jdJQbijHqkv34bMEuvROubnMwavATdxuW7
nadSycH8JiyoNNLFtvOUjiM3FI6GDJi40BaW64WXpAfbq7LAIvoxbH3hPIKx/bJZ+PabD3Hn+tMb
hlr1BiPfptvy2JaqYItCpCv1kylepfH1VeLvbBiTuHoatR7Gy+TsahXnMrOEKzCn51qXd9wWuc80
1T7JZL5RpGL3XWTPfrbGjjCh89ixXnUC6bTinhyX2cB2U6P11wsdhL5eu/3X5Dk4LOqGvuOTNtqr
kElfmQ9r80g/um1L7LGrpXsRBwuXywD51eB3LwisQoYWS5yKe79qimsfE+UloMMTrFvWjWP6rM61
ezEemculkPrYB3DCzfJ8HvzGoKk0FHg4al/McYII3pREBvaEKNsTEGAfaHNHYJzAc7JXDxUTDD6A
8J/YJP7gBXB5fuYxZgPXEAtNzjfGdUtI93qkse5zACFpwy5YnvkdO9HjeSBdy81zhuruiDb8efHw
8m1RODz/tdDvOvChEflimLSNwLkYh7yArgKT0NGPEPy9lo5rSIA8h5FOr3oEQMH3vXBILVVTuwfj
kIBqExHKN7rdGd7llfwnPYp7U1JL7qAGQA9uD6d2NO2jNlViWBQvTPoxQesVnTPqkd3kE2YHh7OQ
VSnjwvDjDBQn6LKeOLgfzEWyAXmOU1/zTRrCLhR6K4AebNcbjbGNplaodmpEjzOA78R+XMLK2I/x
s2Tlcf94G4p2I7Q/ENNvovemcuTrdBMoPRcjoRO5yQxz3n9VVGecRqo5j+//zh9n7CSeKwIoY8Ql
ID3i9Q/nf2CvfEkZb0QfwEmOpk0wAnOyz2B5Wi+azGl1F7RebbqGLs+rMjWXMmOJRfUqUgAfr5v2
sh0rYWtXti7OasZxpbK4tRGnR3neowM4PaJNKycjTH8I2/7tzxaj3mun8uQReeS2NQ0+q6f9p1YR
Q2g+2DQVP09cWXTkPszT1xqqugzxsUDrDXxEBLvZcDsIuk3RTTV8WB4S6xQjungpOCQp+nYIAtVO
RUD8jUgTQFFKCT2FnMkC5z6IhyRn0knTcyPOq0lH+UFReYO2/dwBYMAW8wsMyUbc/qWitKYzjgqr
WEkGRSBfk7j+VYZvS4QSC8b1JgQV/6sJx/mvORxRxue+nDYSEsud0gohpN/WsKoUj7HC2w/4gsTL
zsD+0DFSbRADnqyKi+4dlRYdAeCkFyhM9faX1UaU7WkXWlHya+FgsT4iqs5enEuM9hJXOuLbHHrX
UfCyFzGlRY/3hG1pL3qPLgS8uPAAnzV0e6GUOMVVJiDya9ruzWITDwrbIJ3AMrxAhtETlM7DUwvA
qbr+4xFX7Y3X4fdKunZKMualgoOJiknzn5+3OEIuFYHpR3aUO5SWAlr6TYxSnxCvIPh0fxSMVHhT
HjDISBlwDNxBSOnWLrrT/PYWCGK59rkAnbhDQYJ9pbocMci9/2jaM/dMm5Y2y4bbLkZQJxqN3mBB
2GGuRwe/Q6KgJvtsn59olDXic7z1DRwYX3CuNLz519s+OI4FJae1Hy2C+SNY+/kBJc7MX3BoKJ64
WUWqvWu+bUMsdiHkBRGwYZcJH9HELM0sz6uXgrlBQt/Ds76z+bMXOcBwAuZOHs1NfraO4bJqyujJ
cicEC5cHYSEVtytvNJBP/+fWiRLiMVREYhy1vYcHxBekRSfy7pD/y8zheKyIYRuZ7BsgfG+/eeVj
D5pOlROPr4pfD30NpTzVSwGqXNu2XrR2y/7XzBcRpXyXWqbca69hwiGfMqrBdlsbS7IT7SkuLqya
NRhmtXG5hMVRco0INAbYsm/kg1vJQLyDW7py5qED4vXWRkXn2zgU/dGnCTTUOxB0ar01LBjeATyC
SIhkrQgywOF8TE9OOJSGcxaA05OnJxUJ/xHbOkO7HLhhgzYO06bmi/aFRZOhbyzRTcAs5YMiiYFP
6riAnaOgVsN3Nl8y2iQmMrnyRWkZ2MHBcig4EJKmxmhwDmC/kakHrkceVpJoJQCLBU0+ABiisCbP
7i/vreIdxqgw1VB90KAdEU8JfU2ZFaPAGZK4CS0c90m5wyB6ohMtcFOQhUS1b8ufQoQ0rw6bt0hc
yO/4rWDdEo1UHZGHbn0s0aFTBqxcyqBG471c9VMoEd+c8IIt1+BJPqN8CsqZthRo8i2iKtkq+SWf
n7YyjO5pObL2HLpEsQbufZc+o6vkZO6bPgcdAVV/Zlishh9Moe4hngDkVfIQ0dBxT9yKbiBbeZmR
lBMlOthhnHlHPfjFod+vd56XcemhdprXFnJdLHqNLZLq85gEUpzJvMvt4HT/FIYaxbeg5S2Hi0OZ
zWRjJE1khKUQvjTLfcg1KRWi/OG7QBTYVyVUvZRcGmllXYrsvwrimltLgQeAfp/e/eLq5U4mTz7t
4Z6CfRYCmP1u+nni1WBzQfhxR/AmiQQ1rTYkx89IdHwpN9gItAkvdzI3qCA6cKxcxfIuxcjpnwfG
65dHcH4JSGYYQpF2ABHkYP7HL50/ZBq6b8cC6BfsL96VMhNrJ5fjeaSytrx3UT02flmOua8qLFwX
7AjpuJZevlhZ53cNxiW/dJCGhKa3wnwugZ3O7BXljDN1uUpvlAa1CLX0JXWkDDxYJr7OvF3UQ7mX
B2CQ+ft2nNavYoX/hMQaDLjDSz5iy6BdfSijJncnOM7u1UiLOA+KznnYIk0rqRy1akKvQbGYvwGn
uxWwonHM0AdcDMiUyPciyalPItEJpV+fFJeTcaxqVehumTzlpBmscqPRIKMRWLCOvWtiCezcmaZW
oHJtNLe5Xxpw8//eTshCZjykSLRNo2U9OsGYMW5xXt1a1tZ7120n9Wn932WfTucioH5k7eeP0Gx5
0LEVWH2AQ728aw+cr43Du7N1GVemqLDlJhig9fHhJ//HFkfEjC+jwTtGBJIrFHP/uq5X4XH5MTel
XA3BUcA1ZUWI9udVevt2ytjEiD6unrhrM0kBu7uMGPg27Dq8cB6O+NK33S7teso73+dtNmd8OO5l
sGJE7pJe0kdxsDQcNoaS+diSf+mXf0TJEQd5JUvgrY0fxp/4wlTMJmnUAS8pqfiy3piw2/Z/Ck+0
iZDxANbapvfIX5jC7QXt9ScIlEEKUUGXRKCpcwPQJnFfl07Fx/SOiFOuuYSFc1ddM2aNcC9GKpHk
A3jHeoA0mx6rilqky4xpVIeRjwod/MNVZ8gz6eHj7WmmyLKPz537Nl+PD/+ilsQQP8gyOfA9Fvao
7JHgz8vR5DuqrEhZMhvsnH24vzGLEgukp5UQYxLzfNm3AltvI9zdxiyOOeEveR8wkcOL2G7nh9jZ
2nsJIQ86iUcjzqgvnsR+kf8OaBwyozYu1FkIRfhP1b7BccjbDmRgzCM9uLjTLyiWo7GL7sLF2T7M
UDxtG0mMIT1hjDKt73hypUhXhU2v/ev0BNDVZqFwqLRZl4U4UlDH0hksr+NM1kdiUoyfzljnvGX3
rvsBF6gYTDkHLJ5+7pi78FjJ4JQEsAYDr81J5l/EQTIARtHTj2thTbDKFYtjqKX294QuLFH8PDsD
TYfRuRzuDsmsX4tnucn3mb1nLs8KUAbW/Lf9+3Q+qqVv8e1xRW3mkUjOb3+PzBiz3/Gs0augEFI/
w24X7UDwtuKaWQzZQeVNWiwPjsvwKBv49rd7RTWjZT0FCXsU3XJ7Cmxom1+iLp4eDyt5g/CPmG9/
bnykKuTdLehPVzwbH1DUguXsQLbcZKIJKdJpy43FfRF5FCRUXhweWCm7ehaCL5FwX4EW4hKgxXE7
cquLjT3bXC3/fRTm72mNDsqsMyh5k6MivuVxdkhcOusZnOKI/uUmyRvLgOMZYL80GmtpuEEQCfKU
Dql5DlDe73W+U+FNb0vxKMnbeZ+kr3OK3hVMCKufkv6SrUzWIxgdMhkBBCoI/2cJfpaX0Vf+X9/6
vDJzblFcdLNmDshLnBdMDZ/6vMO1icvAp5rxfEt002ef9G/KAwN0e1YgeWMnUw3ZEnF6aeMN1caE
dXmUqrd6qTXeh+pLOO8CjWsEC28z9tswX5bWkBrCIr5aYOPNgtwQzFo/DaB409zdfTLoxTq/M0+J
UKuuE9saA9V3tH765c4JLch1QQZCY77WLSRubMiHhKG9MO56XpJ+T8/nX533DItzQdjOCRL5wmud
yK94NjWkLCUxCA7hAqlPTTG1ty8DOz3mL8oy7Wxnq2zNnq72ewHRWEKLpiQLvqw5l2yWGeCM/6Hs
AcKy9mTZlIqnoiE3LUFx7GOB3MJjhR9iZn8cNdJqHsLF0skl4bB7+uGoTmepP7VyVaVRFAHiwxeT
ZFbsNkxxmbkB9jDdcEDVuAw+OTFG5dHnq8zX7w3rckvYstqbbmF2qmmChGmISZLnLg/XDAOxU4LY
s41jvo+/+vZLBmOrCkJU7AElKQkNxn9HnnPHUO5scHDCTtcnLVpjS+QWQHec02ZdKTjRK2clCyqN
X1CxpPa9s7dFkMmk2ZmfQLpdWBOJ5otkM4a+VbsvfQfIsnWA2o0B1BdyrTIPcbdYqsJq7MrmpbWl
wPmMmleP6jvG6wwzJk8oBn80j5svU93Jp9XwiBkQLrKFmRiJkzP9lYST8QBz8InXXJMIkne3/FbB
7mUWVWweHk1QBO9hUiONVvBD3w9GELQ5oSd92Tw5bZAaPjJ7oy7MEop2IptCsKvnW95ndlwwQFyK
rmJY88GNLaRVd2hbH25Eey48UrCoNWkFId3fkFKA8jFStcRQJ3a40Pr+KRwkAEe3UYBBkXqBF62L
9lslCbYUBBPs2B9gdE8IprAU9ouIJnPuhJFEdgNtDWrqWxT5WoL0WeeeMAGMoJPbacb7dAOHB3od
cdQsagz3BWIzsNeEr/5z7ak8HDoBFWZdUKG2BOIVEKdn+/enyuc0e4g3HLa3oFa8g0M6ZStS77MI
bIEywgXtY4sYWPmazg5IUFyRPSyJhQqITVJZInDB8rgPlfJUhT1fo6F7oyyxETfakPpYoc3gXxHX
97tVCJG2wqWrqrMbyizBk0Tf14k37sb3wDGqDKObWCRWhIfDSx5J0WHrPpBZE32QNw3VEBQlwQK9
4L3+BD7OFM4SnkT7tACbEgF2q0SPlbEIt2Tr15UbWAOfrqEP0wyZXX1nR8UCKZ3Olm/lE6YUT2zV
ueJG6LH1lMAp+vVnKn6JdwkhYY33N7FuCu9IpZb/g/N2+A+e8Kb7Y56HeDefd5nbNYc+JYaTRsqB
7og7Hy1Xv0x4lIPqtXNyBninpObD6j6J7Vp5l49SmWpAN8qDd0u+fLyxqOfO3z+MoQiSMtKZNzYK
pWs+tScOewXHQPES0me/KuXyJ3sCFrwSyHGG0/WS9XHHhQu6suBMhbOtRUyVxB/l/53/oUwcvYvb
IE4FhQ4TKqUjIkaAtart6qDrxTRLot4bBayVO/0zmhCs9/85Tgix/zWIzx+2wrYN5y+azvGj1xry
OG7PylljjjMfXcOugDiJQwSXi8v+WcI2FU2keHriqLuRdE1itnHyXL4sYw07VZ4G4VXz1ntDYQlH
12cehh+EmU/JgMisZHGxXi9ViejzBJOTTuw1kiybsu03OiFjk1/IWbyUJYY38MXCiOHcVsYE4d+y
/xnlZWSAg1pyRgff4pbIS2u8YEQbBoy0SyWa0uMIQGa7Kvv8B98hA5DEDGw/5FDhiSoF31aFcDM7
tzhBb57y04bo/Z94CE3Hj3L+g1hSlTRaSgNGYaR2Mr/JSgVvRRc3Yi/igS6oYCoUjhSGhRFOWY0u
pWaOtBLi3c8WGR1Jrcp1WpNlV6Ipux7mt0bhSpxUFsImXi8LH/DvrjxNN6VnVNxoCxZ0lBD3Vxja
7S5/oE7aPf6P0C+AACxX7HSHekmysDb0X38/LyaZDxWMHAj8WFhfl6c/9Prki1R/S8C6emHNASkz
EvXaSp5bEKUdXyxRwXyKAIcABRkG297gmGefdIUhaKGxt2TujnUFaQv/KYRpcxH7439JnfTweoGo
KSXEikxLPWy5aFdUiosUGXP5VZ6dKyBGk0kO8waUOKcOGySk+XApq3QBnSticTEz7zjQKviayt/y
Rt5Mwr6GtBkqcYtOKb18fB99bo3x24FjoO7FmdBDJ1G/E6y6/5ypEUvkZfSbmz4BU3HPwLiPkha+
7wfRLZhWum25BekOYon/LYrcBSjSM73Ejbr2uwsbynmujZPwJ31g48ELX5YapkYcfbMbzjIbskHq
F9/pUYQtNGdkO4ENiUfkREu8w99IlxOA9tIabC/FsGUV74dhuoc8qsGeB2K4O+8kZ0JoDitY6MFU
hJbYiKd6d9LgR1fOiR3m172AXp4reUbtEqv70KlGOo8WBShW2RgPRvBXfjyO1XR3GhcO53HaKZAK
ahdsdLTYAFFB/MWCYibpHEaa/04fZMIuJm0+1r+TMpJF8kOPGUKYVnFYjWXoZltAc+26b7af3AUT
WaxBP/wMxqbaksBCmDafYwiQO7FLVJMU+z8YgPjHGefGoyHAN1lD5iP6hy/Kun594tgxZ1oaHeaX
ey2cQ7Iovq4bRKGNWcUG84kjAAdo6DQ7COxpfuU5yjvlHrBDm2FSntREGU2mQr/tG2I40hp0artb
HKIpHypyc8ag1M3ksOaV3N0zijYAHaqXCQB1/tR9l8soUirF2twMNQFZnc60eGClHZ7KRIGECK8P
ezuUMJ7t6SrTlJIG5+gF88INZoJAI8vRoACy3bNe/pMVi1asxntmzOGIDVONBIkbXb7DSAfHI384
V9OCptKpsrM6Zn+AAnvR19V653A7Y9x0qcFklIz2cYjV+FhBhsqg8m/mSk2k8dUoIWHRVx0mO2DW
15vXOqIrVjIsenq3iGsBofLUXO7D7oohAsHjBewIR1KboYFilnz1mgR7bnIRtZN2nf+zRI3AQ03k
Zhl4W6BH5RGWtA1eWJ+iC0rAFUS2Dp96IKNIfpxs6qupgJileBfsJ4/YM3RtEoUlv6xDkIf1dMCw
CT6eVqMOnCFwU+QxyN7ze7LmJrKOHaWOJFBKTahyXmwteFEVngwppVpVxtp3sIKI0XyHdo1bNJDC
FQ/MbdZGGi/HjASu/A5TiaIQT/ngSg94bYU13XarT1FjDvqfAEpfn4BETktczBFWX3xJy3NRcXiD
sUr/zOdC+eWSxk7O5wF4tkRr4HdY+9anPBJgilKOSz9YXAzHPn0xE4PTb6A87W2EsbBzIs93gwAi
PMBVtvijpJepKzjoL4+n1BGgNNw0qlxZfDLfYuUdhz/IxjXqvU0FiYMPTqw4s8O8AzwfnE4e9C6g
izXEUMP56xERBldtYfnM3OxGnvMRGWdRupcZPihN68cM1p/pPg9CRTKhQ7GUAq2idaxZTdZ3yQ18
iJ7pQuntDiVFzJBK2uVNgivIlOf+fOH0XToSfz4tAVqUzgbHWHuNM+4GEO7k96VF7fMiY7myNviW
y0SCCUZEX5GnjN8WID2xAVrG8mFYkfH3jEpJzHTPPmEP6k28F2sZc75DZjLKZBN9KpSvC7J7p5nv
y3DYDvvjA8Yfqlkyuo7hBw6IQe0nH2AwEH4fB2p8qsXZspCOgw14maDk0JV4eESVF5y2ajNPmDsq
QcBuTwWV8SUUBt9jNm8pid+ShDheVNgp0oirZy0AhmaJJ+pBEGMOvYSYf2NWAw7BSLogZ/vzqUQL
Z5DKXPm9zBfW4/nCJBKASNo+Allivrosj3H+PfzjCukUcZ7GxI3vyD+Oxqt6gzkenJujdfd0Wlum
+MLk6ZkMM6HtQTu9E/k5/iJ44uxs5EMD9D4kYV/SipICqf0O/59jgcLPKzTaqbE2MUIx4r0EOLww
ZbVTsJSlIxyRL//bDxL0Hc2m+HjdRbXsEN/ypQ54b53zDXT5mfcm0qt6qQ9xDi7cYv/hEwAy+ITx
a5H9JffbZa6fHntfMWFidhj71+4R4P6V9LqHLoeB4HySNpP99azt+lBKdwVFibywDcEqR5IcAshx
wJa+LikJoWhLM9x6uQVt93TpWBmqbTXF/Dlul0n3rwDxMlOJLf+eo/NJH5HY/6n3DL95QzNswyNM
T2jjZiYeKoE2X8ndJElVWmM/XnEg3EkHQGbmssBhjqZepFMWvWqBXyvAPveW0JDyKy4QKRAk+ma1
BEnm8siLNR+IdbqlE/8XgSpd76A9TMowrglXTD2TgoYdY2NGBvIX97KWNLvqkvoYUbJHX+t59sGk
sjE9mRFoaTu1/58XzREM1zw/5E1QYsCyZOmPpqQrv4WAMVdYpbVrrWRJnyQXvarVh1bEHV/1DDI1
ToKA6K8oLh/I1Ri9+JMAbFauG+hx0QOhFvKUYyD1Pl7DBJKQY+kMwxaEOdkC1wDxIMPB/2MuOrPG
a5E5bigZclgBXKyGa1YczPUYsuJQZQ46EOMUY3peqR/R8IZp1N3psawq2B6fPLYB577IkOOafo7w
6DApWEiVDzJBNQBfi6QlGgtaUk84bRbPwZdfcSnN00yaFnpxEt1mW79c+Fb+i5FfeE7yXYiKlqhX
ZpNst3Q1SMv2rHS75lA0wM33l1pkW86t61n4BWklbau8No89U0NEx9Hb/PT9GVANSo9d/cCSJyYW
Z7FsTDoGB+p8V+KG3SAlp81YZNfFfemW+Y6FE49trPREReFkceBXdacopLvus3nJlZZA9kqKiw0V
Z7ysAWs08JvLzXIg3ZdYXXIzw9stwhOB4coLlaLmr15eS5CbgIO8I1QpefxtOxmPFp1XjtA6+OtY
Il5inJgqXPbWz6HA+siEmfQKSHLBsNMoezI8L8RQ/rkUHFMrBzMWk6PB8M/gyXyJn84f/3qUl9jY
HWtvBPFcNEDR8Y0upraP3MvRvkFb5LthD0pRVD2vZ/rTY/SuNlHFCKYhLYE3GdXbdrcn7nrt/ubj
6ewClq++6+7hfI6RPcB9spJrB0MQKrbpfUEFZ3vIwTSdrh6pCnwdx4X26CFtky1Y3LU3DztQJgKA
OK1TkzbpmmFv0TuM4G5WXtFborFnxz6LIgyUQtmuyMOxrmfiynb4z9mY09upTB1Ez661fLGI+YAo
QBL7xwRuGAeBKbxzZ1SLtcNIskCvNQlJhK2XL6XDLGoFDaZxA5nSklGGb5geM75L6X4Z7Qkt/J4+
khK2oE6wo0eGD4Y09Wcc2CewiIlS2A8Uv2dq4RibrNDyualGnv+qIkuJONOWZ3f0oqrXPdjRJ+iV
bOeBGwK1ido2HUoLjFEGWQvfAXPDcsQLaNh0j3uzSaj+dio0BZpEI/k0MeXSpxwpqBWypOVNZ3ig
SpmT0paxycPNah0bMIHZ7Kj8QJenZpbcj3fHyp6qwqvGWrSnzg90A53FU/DQ+6YmqAGlroXS1Uxm
273OVll9X0YthxGq34HPmmCLR7guC8j2vmlL9yk0v6iiMCxPSvmilD0yVTQOvnyqcHVM4MeN8ATx
npuPEL7pluQEmjduq1MX1A/+N5yGFfcYY/hDT/eWWnM7dJWTkKTahmMXC3hSlAlxG+SRcieKymFo
1OeHRl4vKqfqAPYOXX5CHv7og7eGi4FyUL63FAdt458c9ty9PwkQ7aAVlWehpWQwbsryf4cAHcQh
kKucvhfHJZHkHCijr/WncB4tzcfpSJT1O+01dNnLbvO1YGorUrCSQk5GWfeMQSRDztEBkF/20zKL
H4SEP6lcagkLtKygxg1G5Bch6y289Vbwz6WVrIeUJsllp9uSwqIZSDxuqrs2ubOcKAe9/dubYtOE
Jp8b/HHFZAVnmqTa261LG6iRVhH5b0sUnpdxKIVSuqiK/IFhp/RWrMX3Zm97ZZNTJyFfPdyTdSEx
0CzKsJ9ShMngL6o5ooZwWBDbjVeB4SRtrLwsetIEviaUAoO4tNohnjtLVNtFGvup5QoG5Nhhdw5q
s5SJjnBYBNv1AJCr5AA6+v7Mf1kCkVUs7dLkv67wB3PFbtv240raVmD6jv7W3a91i7RBiFSzkAN+
/i4UNXdEwAym1ZWGD89+ykp1kJOeWjDxiiMYKCdJDvtx8K6xBKR1rCSiUmZ6W9M8cUUEl0LRPv9P
yuVmvi3D59oNoS4xaL7Fr+DFCyihtjQUHaBlRz29d4W8b3RyzJV1AdJZANV6NMDgSD9n5HLLJ87E
heA8dvkve3S08aloKg/+12ExUDo8LsPensSOSIptwS1RTHk4mWcNqfljhBRUhbNWd3hHM/9AjhWW
uzW8CCQHthXivVGdZvJrHMZLOC6iNnEurc6uvoF2jTmCMw4jeg/Wo/Th76oKwuclz6e6hLry/fE8
hPCWcx1FZIh49Mv0GQZmu6CJuEnMPGePE1aF3fjzRoNVIc3UWOT4igPz8mxAZfLt2fKaJ62+3ZFo
+BTGSV5cKzX/MV1dxnqeh7G1oSyv5/0b48RCkwtWhzFpfpS1mJGvrm7qvMAOz3Aw6oT2GORS+Xpj
0TLTsiXpfSivpD/JwfbYi5PT+Iq1MSbSMDSW2SdVmYvdag9mrT82H/hzcwgfYNkjiuRFROe8i1oE
iEnJYSCY89DsAjrhBRn1uHBBEnOlaaclir1ZFu5aqKS3TqOyFabm88omJLNi4z+XG6hfycofQ0hY
f346Wne4YWYX4Ak1u7CybzgvDSfL/DDR0zQYr1hVJJYam1LWzhho+7b2H5Rl/ABQZW32GgLRKrwT
Oo/0S40C4QxS4eWSwdx6AQax9uVF4Mf8FIlfQv5KNZbBc4uDPO9Rz0UkM6PBdLopJQxWT0IgrkR/
NaI0rpJmku0+Q02nVJswK3BrgGGbSi4eCRUNsz8TU2By6wy+w6rNWnlcSBYc18b6aGgwgV4fU8NO
2QQpovadA5Vl/aZPDlag6VhDOaT6iWPs7IScnmpNya426V/si/92xRcH5E+ddfWCg0ID/OEvpJon
8M3IG88nnnbLsBMh2uCCi4yXyGpib8TIzoTWmhhhj/Wg1BqR5DbNOV+/qNUlNKdrhhPRadfWqGGU
2UcKfKTq1DLaLy8bJPLosjFPhB6lWQPl9UOHjp6gQ4S9W/vtRWpCjcjJYL1JnIf9HnjvnKHH42sa
EFIU9W7FVeO7x5LZTaLjCw+rpI6lM6AqZAbZSQsK6pc86XILSzTtyya0UFy1gE+TM6q13L2O8vM/
Sx0ssAw3boGoI2JFoBCOCEawPyNnfGPJny8CLnMy+Ovli6nvNTiCDnIyPM/D0wryWCQOcVBFxQqZ
msq6ZzTF8eHZYEkEStvzT1H1/Jd8i0kyjxl6596za3nRoV154XiFBwaRASlT1NHelhLScApm7+wI
KrWzDcF/SmVa8BpqW1OdEqKH5X5RreLkFD7P4U07owKOGN81aBYnl2W4bB3Snn48dxauxi0aFTpH
2t1kez7HTII0S6S5tuGSTtg/rK8wvtjmEnFt4S+QlKPXCjJ2xfHe3ZIK/WsmVAPNk3futWnNvVHe
MwDoc/vg/pfz3mK7X9EVh0p5CQdBdIkBjwSGCD9z/Y7AeNEu1Kx3facWKk+tmHROn5Q9XR7poUoh
+wzcISTBEAL/h1HClcO3br161OjiWRyLIOia44ufJSS5LPPnHRk2ULGqYOC8Vfxk9XrBa3F1cP/u
lwqmdcXHtwY1djY1VnBuXrX8/a7T+Te2mPA5sovgJlsl9oIlvoXAjRQdO5rx+YEjlE2Fkxr1HeIk
A5Wn/RJ0i1/q8qojgd4PIgh00N5LgmD75zTfeJC481MtOJru7MW3BHRyBHdaHv+/eFTV6/BxBtAT
TpsCcAAmxG449NP+jg9pdm0xTrJ2FLE0T2REHGYK7MmXQEpKbV0mxs1y64wnCRfZV6PIdJnXdCss
Sd43tAVlhbMqUpmb8dCY+BFilzKYBD3/0KBfVruckDa7YUn8x8tFsNxoIIORo9Co4xf99TCdA8nV
+MAuS51qt3J/VOMdDI85ZLMwKHjjL0XE8i9mrqmuTGKkV9GIYaioXNBCWADeGhI4PAQv2zSOq/0t
vNP4idAN7hCTAxjuNrtVjdYLqDMva8Ql2GtZ3Acb1i/Y7wRpyWTf4KoYPvdnP2Isjc0GRsGm+7Do
v8bdhDobetxMRyAPD/oozkK5ijt2YFLfQoRz060H6/MPI1oR2GTmC3Mj70EMz+sex3WPZKEz7xlb
Q/NAX18anwShupnTIwlP/maiJRVcTIVVoXt9Iefb7d8Dm2jS3QD3NeMgvGJ/HWSOwqX92K6Pg7M0
NmArmx7WnchPfDBXGNrlGSHnn+Rq7gpIKMWKhVyyT9gP2WEmH8twSG8+M/s3+4cxty6ELUGcpm/Q
nCJ1DpmcpebWfj8qBi4LXQWPhRtSTruTw3cQNaYogAgvgQ7j8VYKzG7L4tf5CQf+ZcHbQ9nBdBVR
+ecOVMPtnqLeHEgaUKQ9vRAtn1gupdXV1qNbSF2VFIrSnJZ9EorxQoA4hsGgYn65CPjjfEi++JCI
xBKGZyQn+Zxjg5b5sGCCB6++XDEJhSNC4J1uJrvQsSxibQKbnOvXq4tXIokHReyc8QqARDoPlz7C
jSltai6FwGrVLL9PwhlDFFkhzcG12NKHUm38nppDBtZJYaulNiNDHT9V/ArDhI9vlOUXBPsaXOM/
uNXa2i0dfey+H8wnR/Y1923ey9QriWKg9QE3GN5xbG9baN/upR5IeppMwGh6DcVZl0bgaltt8TGf
AzU2jCBd552b5WBp2msbN39ScWvGXtDU9Knnd/iFoAT/1yyb63ca7Eck1YhNeX5ao3XDE/iStzZ8
VYnMTgfFa4Z/pBcVSuurjrrFe1w7pwHrCZPqQ+1JaLcWT+LXx9vlHlR1rzYXRt1dCGKXkcbATOme
lrhk/RfwHrqo2ZylAkW+4gMCTNdKhMrlf/Hdp4e5rbqJvgNh0bdmsBTKcOHUPwZdpmV7k3B9DqcF
tDaP5BfXxTFYoXNQr3YT+yFmYhh2fzDjqWK6mLi14fiGviqPB6g5TyS0+SAC20sstl+IEK4q6nMZ
2H9qRMkPsxTXKBaIl7R2RwA1rp9ojipx1fzLBB5hl2Eoz7sjo6sgVza2C5azWkNELN+jLw7HmF2X
nkbIMjXnbEBugB1fvqVEEqQTPRBra+pSjS3BVsD0NIwWFiMy7p2fK8iPLRTReHAYfLAwVmgF6Vnq
2w8r2x8E2jQExe5lzJA6oS+qF7V7CQaYnt4wr4syEVCsuBZQ9Y8yuNc0rqc9m7M1f2sb0hvhqH3/
azO4U2GL+OP8OVzqqIalD66YStxkMxze0I9hywQ5suyJGY340gRd3o1WCqtUp3vEoXY4dMNi6vv6
pVE567W8MR8vEU9gRoy9UjgRfmaS/ualW9ULy6NnDiCBQ8MG39u0cxJ2yUjNRcr/vyRqb2/mukRa
OtstwCTVXdP2KJ6kmzIntQj1rwCkR4JhzuxewaYKpjk38AR1sbbbuVEaHFW5IYbOcTo/5/bYqtRz
4IfPITBMhDiDcMKymlSvR7LJvYKmaOncZoxs+rAFL9ZUo/1+XXJ2BiK24psYj8cTNzunVjQy/3pM
0mbSHeUM0JVOEdDqIBZ0BTYtbVUapxF1+sUJMllYn3JeZn2MPUVyTm4ie4CXizXle43/py7UUeEx
FmldoKab3ON+7M/u75VmgP5o9eR8DXucIMDU6CD+7YzMCRx2j61SQO6hCrdftsURcmOIsEjHqWci
CSV7XzNOJqsedk9u7MJBgeUKmeckKHSpgXKLPUuoDyl6d80pi2mHCoCe190Zlfi9xe9BNdV6XHyY
m3RSsdbWrG/N9VvNyKeVvDhM8bKjEXl2+KhtUAwJutU2ihPoBKAhdmYf6kdowpaiCmiLe1zIlYtQ
tkfWNcSQoAG8Qx+Kwdywx/+7ToQdBkEc5jmMK3DhCtEkAxkMYjwkH9ql4BIptUkdjDztblyRScOw
4XvOqlBO/LRm+W5nfjt1OuoKPqURhrkyu7cFOAiIujPZcutPgrVaLNepBcvreJ39gHOYbw8P4Nrz
/jYmobDMs+07lHowNK6SjwZI+uWBGt5ysH3aiq0rO80B6g910ZqbVxImehcd6SIN1R8JG2T6XNiK
nBdjLWws0zpUDfjRItpK+m1dQbSPRyr7s8qHMs/zi9kMEiDtxQ15K2rSM20tGvCOTuqf81a2k6lR
uxMYlOa7aekgn4++ru88Jus45Ky3sU2lLJwBasIE0UaZ8xdzVXhnTj6WVal0Io7TzpFVA3zh/SOh
H6ZE8k5OKqT9ACtLD9BwFnhsIYcunkD01ysh54Na+ByJob5rPJMxkyODKfpdhme7lgqyJks41zN3
NLn+wJFfMzGMYmWORC68/RcHy8RVHIicq7pR0i/iejyemPnXKMmHzqUjokRYRxtjo/XoiaZtWU43
1K0zeo86YFpzG/yu/7waPp8F82nJmZ5MIHFB15h6yxzHAj1+AOcr9x+pzm2KcRv22Ri2NWFC2Prl
VJxwFWfQjQDGJIf6GZnrw1oFBY6hWmi0E8QB2bkQBQ8fAz42UPG7vdgiEWrdugCJkEdk08en362y
8UddjFi29i1IwGMFAxh5qcDTUigyCBLahPPaYKSYuCmVj2ArKGEgU45J40kgLMEgw9Dzx8Qpajgc
zCRD9Loi8CVNhsLDLTxIyTGkRowsmzMCljS/fnB7vfj2OzXq+44FMMroJpAHeTJ7CCo69ygykp/I
9Zh7mFCFUllbH4SLgnVbjRlmJvnt3qEiphpZ+AQsJu74NV2BWE+ujK8l9VhtuzzB7UGytwQvJ/5h
CroqOtYB6L9iAaCx+6crYOZgavrLk/KOZLVLRQd+F5a7gDvdbNZPlXo/Joy6UuDru90nE1eT1BnJ
6GXr3DkTQyptb/G6D3Ol6m5zpEk74Cct6ZqjUALyjTHT2XewaKFpo6Td92AIQ6xp2vBam5J0PBdg
0HcxA+xgVOZxbwQTgCaeGPWgePKJDDC+/GiinDp+7aewpqVHLP6RVi4CoNbWmDeu0gIcI63l73N9
Wiy4nQjNKR+EgaMev178sAlqvIdE9d8eqTBwU3jQlL8KlBO6u1poTRSJM1xswgq6N8LDiGCeqPF8
WQUlN3DFTMlzQ1MwhujumCTlMp+SRhf62SFxWJnqCGJpQzYVgHAaDlyGB6ft3adzKRrlnsUsEuks
5dSXyYWsa6Fh2ASjbaA+80y74rhH+8tDTKtybnHyKBIVFwNMRmjfJ5j4mNkuIjaDUlG8jftQW3gL
trBTRc1RNiJtItwYKb3yizAM4qOlD5+ihgnmzLfLnrRQ2ZXpdUyw4Ln+Yn7GguWO8Av8cBiJo/sm
xkxiZUzNt/gO3ThUngoJSevZ2Kgbwx0tHI/foqWDNQsgZE/uHF5gYG1pClfqHWzw09rz5xDi3L3b
q3sFyUtzPl4HhEq5ANLX+wFKK6J6we4XUhOa9uZz3bWeTSnQBDMookI1ZR21Ri2eilqaHnQXAEYp
on4n7QDBx0cx70ygseefuJUgwbw7gehCQyTiwueG+aBi6t5wQR3bWSvXq9IWHt8kcuroQjYpZFP/
mIvtzLwfn5Icdb0unuiud8AhyCLAIvmnISf1FT8poiKaXMHlLvPw918lLZv7m7vTbmOYd/o+fvkR
3Y3XoVsMZ6KWSkhgDPBWT7HhzasuMtQ6NNZTrM9a5MlmbJkvVO8GUiWRIr8+70msLNFt15u8tner
oCtFgxSBJ16W2NKxtqeGnC0DICxoN9ZSkert+xb0uv89Lu1AMxxvrqHae12QN8m08wJoAgedMvjY
Kf5AkhJWZu7X5wCxYRRh2GOQqmwI/yXucH/I2vqV/l61VP+sHENMjxbYlgatpcqV9/1Op8J7Kyuj
D4BkZZGmhTpRecQ7lypoYndtRqBd4RlDDjJmeU8gAFDPIenjQZqfzdwGno9ykpN6MXarHzH3+Puv
DtvFvEWcNoJApZmIfpd+W/5rDmhPCXT4oWrRpmGDUhqsI79H8ioTK6JaP773e2x0Ofj1rEluyLq+
rjTYtY/qNMeyf4tqLpNlZgA7E6KJ6OOki3p+gStNF2yYzM+j/W4av/zezD+N7whcpvQIBYQac8IW
GBKDzGR3zcxKWXUxrGEPEcjV9U1k4TtoQw67c7uL2ww3GuHMWCoVKrjs9/Ow0FtBos2rMMrSUt8w
qamzkGdBXzQJA7F8HZssH9bic5MCxF1UFIBEFBGdGn9BKe5ucWqnC/bjatztOq73HfDJk2sAN2YD
nA2i4QNIuzemnhyY+xH0GUlfW3nnq2RzoZxsLIO6I8ffA9D5oow7ucIxi21yqxhpK7VEZvQyA1xy
rYHMzqqdeZR44xQnRqAt64AXj8K82ykbrrJpH9xl84LXLxBWz3lp7HdtG5X/7YM5qsZ83oKhttnm
J1HfAqhOp9wDkbPQkLBp7yLULPCXAa/DLEYTlaNPgs/zxpeSbh+Z7LEaBEbbOOdvxUAS55MRj5CK
YnsXtbKsW4DdLnZoKnmJ+39ZrywevgzZz3xlquTTNsHV/R+ayeNkfIrDYcT+LpAYMaNLQ6iQtc/P
GXIRdZzOtL3EidGYn3sJBQRAJXyBRRU/MJPQ4b1ODbE5W7eHaQKChXb3dh1nKN31ZVUBX57W/bFI
SzJXJCFwaiJb0DeJ6D8rh7b4gTFAULbE1Yrua9yUjSw1QHykBtzOjUSWSvgBmObM2U05wlAMMGKJ
4pB5b4Jf7bNeS/O2X0pTm5VjRSZ74TB8uzkZPw4u6RbAq/QDvvHBT0nXqXC468Qxz3S8AfH/hski
nsqnkl/n87SgKUIM9VnR9lAfCMyDxLOnNb1w39NrrWtGtzs7FkFjImgQzV6+v4SguBRVuubLfAOc
N9bx4xvFgvpJ8sFTQHIxs1qKctB4kdu44Nh0OB48gqwmu1dFG5/3uU6ItC9ugOzarPVJI+cuk6c3
Rakk3ThN7k44qeErvCV85x+UuRG3WEdTlacZKbUsqILGvNOGYr88YSz4Fw+qZZwSMFCJ6xtnNUpL
SkRaR6rwfHX3dQrsDcBLiLahywwvXYXGsEX4c6j/hD3iEREV/j2ZLv9ttFNNPT8s4LUn2942Yb20
1eyFbXYngacH/q/VBE9qWF+t4OfIg3MkHpe8nH6+MHsjZ4I8oQok2IF7lvZl0qLoVTJT+FJKOhvH
8rfXRBc3PSjonJ0/MC/6VlMeTZJjUPi8aglb4YsI1SCwZE4wRP4jclXJHcIWGoY/cK5KtaV5huU5
5PeO3KhvXqXm7Gd05uzhMwrlvtnmud49gs5Q4ZIkjj0r7IX0AOD6ZdR9QH+g+JXC78mj5/x7yX7b
lHhiBDGRMdRvsNREcEkO0KtBh7mp5PsUcCQrKarwqNCNKtux2/JD7DSnWQMsW3+8OzrKQt5PK5gK
kYGHOzcHMCHl5b6Utr2HQTO/vDKcTMVp9riEBA5MMIH75kHCVULga+frTnmBzJeBwJpNFuH2VVOF
YKc8Qsd86XViJRmyVFyU5Y8bVxAL5BLdn5/4b2FsrCMhPXXUiWh/61FHAhqmCJwxFBEALzdFbRSf
bwCiGVyt/lAD6fUTG8GBv9/3cr3lR5gOAz5IJZd3z+s44bdOslionhiXGRiH2JJ6EKkLxr0c2SnM
fkGnTiEixDkjUeqzpp0QE1sEFyYCc83N8eJcx5unVJ51DOdFbmEeA/IOCk/yN+JFHLfxLs7m3CcL
2ofVLx5qJT/3zov2RzTQAU+lH/AnySTgL7HUYvMuPHvyzUrdqYfVQfChGMrpKGQgPCEkDxN7qFH2
jdyC32eQPmOQAc0oVqs1vYLDu5cq8DL38lWSpk3TKfs0OiXxRC46oPZjU3dPjZ1WLUsWv150MZ6B
FUr3I+ouZWRnJSIAnoMhTTKMlKnlK5XFh4cmnN9QfR1NiANrQNfN7/yasw3ygjEVuGZUOFXrrSVR
SVsKDvczMdoSpHJ2fd2HdTu3MDKxQw5XaClCmVxgkmHSvVl1Uqdxlubo3LOxG0FEGA7xBUpmsfZ/
YG1mT99O7efOHHyvQas/Ho3r3Y3RbjUeshc2lL2DEG/HxeL+gv9JKD/UdDZEZ/WSvlP6h9wHJsdi
9YX4uKKHeLld3nYDhHoDRhXJwGNPb8GE8rYIYrR2eltOwRNBqUxmkQHmXApKb+ZZNk30KhA1U23W
XE+/echGgVU7RbbE0j5q4fYEHuW31rzN6gwY4e3S8AyxQBW6VDxBwb8iBV/KTyT2oPD6Jn2LTaSR
xJaKXFPPFDOWSl/smq5RSseTTqscdYcC/jhv44/1CUdNcKPjeAkS01k2xmETha+HJ4eRFH6JX1vN
a6XGqr/izUzprtTZOoLVLYGUNSOffmDbAjOhu0eVjRcp60LLSZIAeuQghKG6Ff4KTBLEtqLrHYOx
LaGvyE29OxKnc/VFWCE825GhWtpLBl+U4gEkLic+Hc45ZYiJ8Ovps1qw97QrdCvFTs8+5mhME0pO
83laE3/+vgrizr+GtrcwX2EoLg3hlmEXnAD1GMojdPoSEmYK9FmAtMPWQjhDGAn+oeVc6sk6afAI
BJazAwclC7BI0w3Wlznofz0EWQl387BoPdnhjaxkd5MZMNagoibjwMlrvc2zhc4DI44izPmhi8Pv
VFtzWfqIyleKm+Rd2svRYFGrxKJKbVJJN1fstb/cFI9NHXHDvOtV/k2eu7HSVSpucMVc10ZoQ3Or
k+0qrjW9tMe7sYUVtplLuRxD8zNcffFo5+fhe2YeiX/rHsfySYo5CqauPP3mIxFcmZVYKxuz3NNC
G3lzTDoC/bsNN2pd2GJKjBXJ70041iRQ7qH2dswGGliD+0IhdTXKN/vTeqbXaHru7ZGFH9tuE6nm
th/itqjtByd3DKaNvhNy3EGFcM27Nz4JfPX+NSA6XOgAsV7TN/uReg6cmBkQMzufUlljAg5ucDZL
WBH+FWYfQUXKQDcxDUGTgG6gccyQ
`pragma protect end_protected
