// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
MlcKMJ2FSS99yt4+hdIW+CLQK3W/ekYTS1Z29tXDc5su38au0x4Hx1EMlTe8
kqz0j/cMqb6ooZ0c7ILLfbk65W8PIUDeUpA4+0zeJa2huLArOywA1Ugqr1yW
opCj5yRKLlgOXSmTMX8kVuDq3e6Juy5OGyrNw3kKSPsLzgTRsMnjnx6FGQBA
0mSYiXAZObQwhAru75I4tMbPn++6hRJ/mHsh12hDrE+5UxvBw4MnEAdlG0PV
dXyGEEvH50iH3e7T81iGH6sUlNXqILk2OkyCW8SjhBsM6olPCKLvu0FsDr8E
wZCMX9EBuHipZGABUxwnM7uuB8hUNn0KxKjn3AXrtA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
iXC7qJSeaZqa1YpXAdEFmlJsvjRFbzprcxvd9pTSstStfIjUaVQeVWgIqe63
Iet7S2avlt9h44oeiEFZOcFFq9cjL9eBl1M3o+6XpNQk3umQyaV0IrUI5iRi
aAwpx+ZtWFySzkVAeB0OXqJ2Ye9WY3EkDgwqCIqFyjuwx/EGnZ9/bAtTBtQF
R/sPoZwD53rIxbTwXOR95TWdFFwo1NVIinUune8NyIOD6A6D94zjFAsV3b/8
vhCL6b1Ye1gesZ6IfNeWISBNs/79PewykHI2gcTfg1g6XcoJIZDpwS86SdxB
GHQr5iWV3CapWkYCrPOeTHpoX464thO5OZI8+TGTHQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bj6jIrh7KZbIecVNKAshxOA31R3Xc+to6zWQPUGdzZlzcMeEPk7+eT5O2EHe
GExEdR8m0Mgjsm4HYcSfE1OJd+pwlZ3poBSKGVP+360VomPgDVrWdTmmspTm
dw/PHwPi4df4GWh5I0teX27gGTm8Pam1PGdPyAHB3IUtagISWw0EcN5izNQA
uaMcp5UVpb3pQ0UBgO7qXty5OLe3W3WMs3/ird748U7FsEFdPEryPgNcPR58
i+vkLcO6oNKPXE+wDNbgzFsLQ1YbQBX9uKOCz+P02m3IddTMmGp2pKUGV6BJ
6zbg8lTXV938QwEIE0mq0p+Ddq44fFDJnhol9RVOUw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
A31xdvIwtRbImDT1fKOuk4rBujDk+TjMY0Ci6dFVAJwOde3Z8tOzwEM+lHrm
ByMg8DqCLTA5Mc3Or1Q6J3pSBYxW5DYKuEfllHygxEM4uYCu9AZJNwIGpXg5
3BuDrNfDnYLWsqMANqlN8kr1isq0rmdSMSQ0L03iquxaTs8uk20=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
gXY6e+2OyjgWN/LclPyBHDMfBjMDQDQKE3vthXIG4NdPd5QRc6rYYaEICuhP
gSoF76kl4kEf711SHNDi6dm61Qe6hP6LuFROyOBIgqElioH9gRWk5EnOpGC2
dt2KtUwOJDtcW0d1xMqFXtTz8GNM4GU9uU27c0lIoyxeJV9AGyINIiIdRlUW
lO5/77+TNWvHGCImGtvzs38VP5MRWhPEPjEibFtROKFB8+EmKxlw5frcIeTp
UagBj6MZB84bYFN+mUOeK5Li/rgigqXigy0c+mFx97+bwv5mNk8rwj/KyL6g
hFsDb9w+woUw6Z+0vBTd4isnx5CP34ump6gYHZwDmLDQZyemXCWa3v+d0Fij
qsJjIOWvfbswf/D5+umAQkiCq9iFrxyNA4hjImg/5WttHDQkSZPpuoWAi36C
xP0RuJnVya+kpbyJLEb/2sCVOe+pGHJrwlDaba6HbMG+zzkvjFLXpCsX4+v2
Myj3lJ9YIpVN5qs3p20JHUqGhaFRgxWX


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
TMh3mfXfYfJ3dXazT88zXy4xvEjiMTpv/nrkzqbIiM0b6fP8l/bshbYG+shl
CweujT0Q9W8wbnj2kv1rmxazY0oexgRO3x32ZzzBt/j4Bk903OIkz2Fm3emL
B/U9zDbB/Ot9X2pZuCNOn7iYm+nMxofZUL+NtybBdiJwRkfS41o=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
G66vCuVjz/1K5E+Z4X2cuktJW/U9spDFQ+stBEvyaE07Zc9lCKmStcJFNa+U
o3R04CTZ4grc8i+wyfP5dQeZBN6I2AZPNnKa2QW58dthE9P5uV3ZAoMxKCkS
fl59vaj9qsXoP1NVzEMypmUjYl7t7zvfi1iLDPbGts1sXlGg84g=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 2320)
`pragma protect data_block
1p+pmXNZrSS2Sj4kBOUE9Zi1+hQYIwfSBqj/Rk+9zT3UgCA2WDq2+jGqj1h+
tz43WKy52xxFCScP9lofv7iLONMsFUsGnTjK9aVPG+Mc79Y0AI4BhONB3e1q
koc6S4lnhD/vw9SgxFZWlIDqo0pY2vC8/a4kDBX3YxGNuEHy8y60nzRv/9G8
mcLXmD+c6caYWIajdLtuRgZKPbRNbn6ticPeqjm9vNuT2BO6wGjCEKyVwic/
nb8yTDqdlMk9v6DulcKwDZZL51DDcaCY+a0WuKdgbSAQgghZRyNw8M9A4Ovf
pEgcPecrc6dkFDRt7cLeglU5EZnpmurO2Bws5K3fM9rdTYZX9j917a+cxhRl
G93tM2qzTqN28dNsuhLlQ8b7hJjhMfyVMfEKZNLDE3ROetVcjKEyHiNY9MOd
FGlLIuo0WiuqnLlOZLXRDboc9vRHGotZy5ApD7VqJA3Odeqw0C1e48G+Sw4E
U4PytL4QqxrFNil/kT7jvg04qopK8WkRaTjk8OgqbFFw/VPs30gLuX4ZW3C7
6tMFWsO3P1NJODNsb7ND4ixBCdUttoaLRWB6MWUxfrQbNDND2D/stTNdbheK
9BOSBX4s/YyHY0WapN3LWhZfsThurTRKfttBng6r6yGiY9u7GChnG6D2fGyP
VQnv66rK4xjVl6L49/NZ0BIWR7Xm0rx1eAv9S5ymv0y5WyU7YgLM9k3A7Jhb
FhUZ5rHzfMKTBVcLm0Iyqb4cqmqFrsw3Yj1x2Z0zrMtgkuGxCgaOP5NGvbcm
vhfR36gMS6JVEz9IEUvKFA7WWDuXnD8BVLvAg4djhxbdWIkXY8Dlqf2CB+t+
0oFaZGTtN2ror+DHnaF5xnSkmZqsT4PI5ki3ySEY0yMEoCeBzhdirN9SI8/H
X2vONCALKT9we9U0Oe1fSmzP+fhqY2EpZRmGtFgozrzmf2nbzp1vaT9vgYON
wfxEXJHBvIpS0wfTbtUuApy0I+1TRp0khNqqHW+bzuEEfMxhrthitQKYSKsd
XNVlMKfljTCbOHJg64tpJse6GXwIXvbZmUTYIwBLOGbxvgCuOqM7fXC40+01
04TM0q9vmsTox3ItwfgmV1NOQPRNq/mmyeMaICbELXN3BtNXGJDG6Z2lrkL4
F0d1XF/jAnAiYP2TBjA8vnAdywGHm9ju01MPZfLSHLJPw7QAALFIv3HalS+f
RF9jscxIQSGx8ngVdZKp7ERpRb4hJxENku6AX8l31xJn2J2ulccZHFfFlLo4
Qi7+tRkV2BvXkFg96Z+z2SeaEcx4yEdV+YsG8Z+wfWkoxj5kc8/GFxEZnDdm
bcs3XUCP62DTHD1E2W4rZ+DUzskx1HqXZB2IfjYSorovnyImArT4ioYpMzkZ
rm14bx5fM+cnfCKTMg8I0lqXqkrWjp1FM0yQ/iSY4JI1pfEgS452D9FDr72C
llGm9/S2dYDxi9IyiOvJPQzKZbj43Okw/JwRD/NE3DJCuWkUmkTU2TsdlwFc
GFJ/JFL0+SxD3ifGrR1Kghp6zxJziQvKiGz84X8l3S32Wy1VWdlJrstSUaRl
UGYeV4VLAgi4l5Z4r7fi1qqy7PPOwGVcrwczvlIQSs/UbFxL+TenTLty6rhH
LVz/CpXO910+79kGFPMyzmdSaPH6huVjDdJGzT26g4VNVa5C4Cpgp7u0ROtp
VWAsbdI9cUFRsHtMhmuCFFLZa8oMZaOitbzyviZHHshBgu1w3fdWeojoXWE9
HmhjD/4H+vEf3QslcOyaZQMV5YJETZPxM210xDyFoI9cCfz80uQeXR9JOGJj
FlBQKBofakKffIJtFxk+7xn3gOJiK79CZvsAfqKyvxk/l5mbfwGOkvS3RTfv
jVVEcrs7IkpsVXwFWpoDNGK1qpfceGCYY5odEA/PcZCFvXL/hfJbPIHZIQI9
WUlaofd83JiVjipNtavj3xKx/0cx5vNTMXnT48qPH5ZZzPtJdMzbgYWMtHer
WuqJDqKWW5DvR8pVkM6SahmPMgbCEi1vWd7r+I1fzSndoPeZTgpHT+POvp1C
va4htnDYzX9lq4toDDh6MhavhqYduB4B2Nl3UFHk/ZFl/hikmytVKFu4zV+L
6f7kzplMrNffRSbwsg8PmVZJFzBopwjN8NCwD41jRDivKv3F/ykhrKlVebma
0P2XRyHswDAYhdq1XoSxTyuM5Rb2CQZaG/ssXDlYI1GzEUCipU4u2TDUBvbQ
ESNewXy/uZqglGI7Eyxdo4MfLICJR7WRQoZUqpeAnuPplwhfLhZVjAmZ8jdb
K50HIEIXxvuBShMPr0IpXf+mM6RCqzh2IGUS+nr4dwltSw5GpX47PHS6F3AA
voK8bmKfkPC//p8XgrTB8kN23bESxglJIh4N59w5O3zzReZEAeU7Rfz3KSYn
tVl51cMZUvInP6AV9OBjpqE8OxpNJoAAW/e3X2qSlJYVM7WkH0I2l7CFmJF1
Ndte6TiPvRptACBTW4a7esABzoFohCh07NGqD7a/tf0JBz0xwJxPCdnPY3nC
+gERVUhoxdtatM+qW5yuInDQqrP6mTD9jLmXCfP7Q76nmY11r6I9FxcUAKCf
ExPSIQx2BQ8Ew7pbFxOtfZ/+T/UztgWaQDXwr7H9tcedrIaqHhgUF1CSm02G
dLKOouvln4j53iFsSf1hR70nK2Zo08MrCTKu8YgKpQChrpA/eJ+NnCsTiwzs
o8WdwWekWnObAiz18JugpDWHcq5ltoJQLt9kXcrivmx3RfOGVSo1SCe7qTxh
ZznwkHyB+koVR4xGK9XRcRZ2P6p1rXkD85IcNGTGlZGz5wXUmTR6hhLimN7g
zalAZ1brDzq0/XJgwDW5vVILLE6Mies0/p5gDgTHn9PQRiBooSFLxnymAoCl
7bhIaa1MzbehtWrKY/X12jPLGSEWnf5iCTM5hRSDTfRMARkDw7Gc78uUG7Hj
xe9gRMJIyzTY+xBF4s4YFtk4H8UbzQ2ND7kP1n0uYYLndZXgw9Mu69/wyL8K
1uMCkZJt4yaB3Ygcv+gdN3cGW67CYemuHS/sGcFWBbG/wbcOGkPneFY7GYBw
W2JUQvusYZYEUGUqCs6hq4/rIblY8sINhA==

`pragma protect end_protected
