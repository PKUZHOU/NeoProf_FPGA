// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
un0yb4A9iy0Xj99UEuTin/kGhfNMRpggmqS3sJqPZ653Kb3lcdoq7i2wT30vvcYZ
GscFo5i3018Kwp6MByfSVvfg/h0CzXdm8GM4UjJsWtE/2jqv23I3Ib3dB3WfgIFX
bqXb3fLBJgC0RGcTKLFlQO54c+Ir99rxNAKr4zGBiYs=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 46352 )
`pragma protect data_block
Nc6kx3dgSRy4JquttD9JPkzOVnMRa5FajCiLjHQmO9PTjoIg6kenkuPZivxzawR8
X+smNxwKiA+jXre1Vj0zVkIs6hZhN83dpbimK+HIgjNPXNigvsGMIZS3iGSqain1
WI9601WpTle+qA3EFyd+Uws3wXm9rcjSUaTtlQWziJ34dvcTq9ktjQMkLMoznQjD
B+Xv8Wc4ve4KS+rl/yAkXIdi79v9R3x86IEM/0g2O3Pmy56CrG3D4PeIiUbCenXy
fS32Uejfe7zSO9ZrtFGpt0gtljhgNrMelI2mdN/cQoUudqUa1On32hHMk4qOJoWN
2AIzLdZex6sTrS01rDzqnspa88VA6nNo8xdoc+7Us7pMwu/jEt69QCpMIYU2zOv9
64mfKIX9QTnGUnnRUJRoKfIkU6RBTwk9nQTZPmwVIfBe/uQK847Ja+ExVKDevaxI
9MXwMvA49MW06fHYrhVFF4BZvfpLq6BJX1N46Hb7NjCxG72X/eMvl588j9sl6sm8
FiXNuCT6Rppu4Bi/x1deKzVUf3G1L/ZMo3QhR1nrMHkeDADov1vM8jF84vlotd4M
fWGD22icJ95WpwRwSJn6XO/H0agM0knfuQRwGpcDiJdazfnXSoALMxpGQuxfTNeQ
Y0Wz8P5qePq6np2LnIFGyvimFHQjIK9BIS+xduhbCMqv2JWWEv/FSNobY3eQq3Wx
xyvjq/jFEm3G6TAGkPGzUCTQBDhgcvyJKg6aubPOxvLA7P0MaLbn/xxB1Sm0w1/K
fxuXB0LYOpZs8eSDcnlvLdMU3SBkfvci7h50CGpxv5uG/N1ra0VcraYdpTJApIZf
wDyTV5N5X4A7jMyFbW8UCxrqvMhuO8VV+wsC8pib/AubBrqvnBxZZRn9nxpoINK0
gCjj6C8t4SksU1slPfQpqtzkER9uhWU5pOFoVdNyl9rK+KNBaUKFy76qpm+HEYMk
qr8kNQd2hSkMjenSKXcWPG/zPlR4VozQnDyZT/U3ZHe/XolVEAV3ERPER4k/WfBy
haM+GPe5boHkcutfjMwWDOpcamj7Y8af0C3SXIe/kj/ScZ+kz6DhTH9F/AXe+RgG
Ak1TStbTgGOsHri7qV8xJ31E/9NpJGAKZewkekiWUqhw4n8n0DJ87Q7KSHfHpbR4
MGhMSWs0mW5B55KA0c8voaig79Jm1Wn3vvcDcO7GjDTzsVAt2SOZ0Tr8sSex+jSR
sT8ARzc6PvS1k5XEvb7nD8SJDWdQcjiahYyC2phJGQ5AVhT/LKxE5BzxSFuklyHH
BH1ELp1orMHVfSC0TohYlffxEbrBKU/k5L9P1aLQgatorl8Fyqn8Rd36vxEsw0v9
3C/s7HkcTSa4zjf20F4TNo/x7feeeWA7YA6R0CWyHTwPWZcSvPEbRnMa0tCzq1N/
rK2W42dJuqgBlfcJ8rRqVYAvHHoV+dUxmntwrhXSnNY3jgcNZPfzi0f+7TtT5g5h
mUa4K7xeqgHbiH6SkPu9lTY5cWaESklEgP/0gh9oVehR9HxudYs94j2pib2aGyty
WA2VTqFHiBcfNTVq93Or9OcKb6BJkNN/fwOHaYobG4bWeZmv3hg/MhNpyJWR3Xb8
Sh38KSsGHe9EmJqWtz1kHFPBc1SFwkPCeMkNocEW9lBiQfO+BYrwsljqfHW14AxF
Ft5RWp1pV/qxRirDw8s6TcjFp62ut8Fq6HvdWM5sT3zDaPe5CVP8iAdMYnW1yjRf
0Sxu6JWvdTfScBKRKIAd3rWO1tsD5yzhokvmULH0qPtTSfev2MtXQTYG02zWkoGh
HJXqK6u9fbnZNFrFwOCoLXgD/EJ114zHHESfCEn4VhtTcmloVqdOEHOe00ubr9d5
YVCcJYUQcYn85maPwNHebU97f1am0gIwD0dlByC7Ad1hLIqUmi3apR3+Mv2/iRKI
+QRG/IFyAV1fk2NnqfU1F2/J1rBinMvm6ikdKPpA65kpmDFksrIraxeBSbw0bEWG
zd07lqpkGxSPxeryQ7p6dvat+jpL0X+V/DSXd4XW7xu4Qp5D9FunJlbUzR6HirqI
98GMWvRqyxsC7Mm4d3jaOlg8W8pbHpfzPn8fQx04RQrLOK+VWdkOmujfGDAcBqyH
FZIpoetn2221XQPAQlnAXu0U3kPdSswALhBWf167FUKSeY5q95vwm9WCdrVH4xia
PmHP+g4XvU2lEXh5kH4RaoPV2ChPvWSEFMKNDyZDf8t+N3A6jziceAwO8z0ZLsmI
3cw26Gi8c85r63NgA0dIARjay0dcjULnmcSciYmlk0CIfAHDXy8gWwzCg9nCw6nh
4aQ5D5/0hdeiOSWEvx6E5Ale4MCZCEQ4uMu3AZIlGDV7A7y83KvclXY4Oy5zH+bX
rNz8eX2eL9JOBWXUcXORHhdzD2ycB6C+vzF1pVOFh8CRw8pBp85hcAoXcFGjLbPk
hVnq2HzFHsgB1MDnkJWrnjqYcHd8PQEZ3usn6AuXLpeGTu4Ou15ozKdUmXhYNh9e
AdakL+824D4HCNqyfVICArNqluiV+EPSHubmc7XJHiT1+ylU/JrwJu0gzZV6UYl9
DWMe7pRHfdmtUFRIpv01VgKsPXUy1iNV+f+fu0UEUbm4VvqL7rbkMbmxKa7GrGZ5
sQp/5ChIzTeK9m0m0NfyREwAsNrqyPEqfqOuFnzxbPjx5LelXFn0duXrWkIpsVRO
dZtIRWGgmKSwPiS234kWIvEfr/tNNsCG+SJbDabsO+XnhdRyIvSl6PdqQLSZz4yd
37N+WqTQnlerEVD57UM9/V3m6MrzcWeL6lHEM+Q8W+V5xtFyndUeOHlwCsDBUHBc
9mRTBIcZBsqDfulLADWmpqaaON8yNicUzNT7AQKwqwIyIi5m+4Wa5gaSCJoOOGWI
G6jca+eXR2kY2jV1VU2lOl08Zto1hb9vdKGt8gMlWHTzIdlTR0XYr0ftoNItuX5J
mk/jtdtcBBFb7gsY81YJRU48iFRNVmCLK8bvOATaQ9D92v6Ea+FV9VSCg3vVfSWl
eM7et8jPs6JYuyDEfjHOyKBtf7UOUojtq/9QSyAQWwaZgnUaBBNdRh7thns9t3lB
fB7MGRXoCzLyDgMWjy0xLot8kEp7kc4L2EwbJQbg2GghkpJBha0MKdqFBbIiJJdY
4QpcR62erq1KhRUDohUPL07AEpw1MehM4B3LT48QJOrBlY8eBKubY763UjoUBlcK
eQYMcXu/vFZFeSyWRvM/TrrWd9PiUpOoe13MDGGthlmGz2dyh6/32RqQfufCQYbL
Zn7YUivPyxTiedIIdAMfBRecjDgq1yh9bWEIXwpTUNsjAMIWATKBnDGUkttc3193
iSjik5c71VoYkg/x4zqYj6PgzWYCsljjCnzM2OT3H+pxUTvi0Y6ruEjBsRtZaPd4
Y8E6eeBhIt7ziYkMnEW2MVwA4FQ8uNJCzx5JQjn+e9SOw8l4jJ68gw/PMSm2IMJp
hPS+Xg+fly4NpqZq2RSOubTHmlxZ55NbDJXRuSECXzOIvAjuE209xcPFoq6BGR6H
yZa9Q/huw2Htf8u/7cTgSRKl1qUHHpCoU3D02mYJDq5nFn8osXl1kIghc48tubn/
CLUtdgZzCHhW6GSVlsuHuEj6Guq4MnPlBu6I0LXuxU7wTq/nzdSMnuG9k+OPXazO
HkqDFW5vy32rVQS1PFys9o5KhncWdziHHqJ0SALAQKtCfzMLigGrwhN+8BLa3t5S
wvw3JCsa2A7ETgFdDdB04xJD8d4593cgaO1btj7c+eABGomx5U6TskGUMV1SYFus
Fhu741DOvW93iG+QpOLRhisv/gtdD1vIMyD4Vso93cTWSSbGaGE7Nht9ZWNpCbUu
AfPQvO6FNKzxpJ4KbOz6LcE2uYkc2p4oIv6qbqpeCrp6K1aPkJWPfqoPka2vo17F
j5YJsyHLW3kdqf+CQAkg0gbxHyrG//z7Pcl/MwfJRiWaqkPyGH7LnLOKhh+ObK/s
xQGFwV1VIYB3eQSNHSSRgcOCFXw4DUh699GeyUUCUf6/islSggH7qqhySobKCuly
L0e02wgQT4Q7BgqzdBqiL2mAlW7QKqwoHCb0usERDxSCqZ17qurzanK8cX9R7XK5
3CEBZ9KLuz2GodgyA0oYTghYDeC5PnjRVg26c51KFOlNSRKXGTTBohGcOVhpEwx0
whdbhxiKButOafser8oQnFfRxm3JckR1F1U2+lQ6Ui6N/Rp6IbgrFOYCFzS5Z5Os
z5rxl3YvPxVwFmZmPYKkTQDP6WqQwqLb1I+NSk878vy1l36KJClisfBd+w2N6s4a
QVgjt4VLBaQeGtz8NGkp10PqybBnPqNadGO30pzlSzUf3gbWCXThP4vgGTCAtIYG
OZ4njYHnLp/2AMeiuIS6JX0ja9SFGEUUf27y8c6uF+Kx0sPCCqhdpjGshaN+wiTK
eGcprwcZnkkTC7Yk4Bv9RB5wrYotP0TvR6yLwbdjSto0EaKfcTUJWX6HcFm3ArUA
k48RM6aZ9xSIczEjUWJLpABg16QVCGOJ0MCplcc4ZhIHW8+AOX3sLY3DGQUwBIb+
yRNRCQwBjE0qMNW1ihHQg1LVV/3qNdmDIfRCMIocgoLHczwYdIZcPl/vELg9c463
uyYJNNN/f9KgSRLP3l6/OjhkGG561KB7CSJawHYpO/X+QO8sFLEf8fhCdgrONjL4
jN2BglmBhoGqL13cvA0XTqcrF8f3DYg8ld6I0h7RvOhJAyTeRCEfyLdm3UZQNk4F
W4ZTEM7/eTVKPJtf3eapIYQV699JwdCSKEKW7X8K9lLzbO1fVXC4hav4gT6PozoU
MFlvv7n+1DmPI4QSh1gcOSbqbXbc/xhTHB1vCusu4k8xypj2DMK1n/t05XKwHwuT
SQ9Ollth4cH/ncswWMahx4+XdNYfNsNgP/kuXBb7vGEMJwMW7Zs4j3dA4Szf0uwd
xviNcRyjRD+ZOs9zIZu9ZL+Gbypm1DNpSGYBPzZCYDvj1IjAZ2Md1P+ke5WecLP0
V1/Xsz1RFFiIKmJYD75oTFqa1Mo4s9Fof0A37vSnYUl4DGrL8tOasFfhCF6i4HPc
4U6VtUim+uJZi5hTcJw/ykaVQJovBOKAx4kfpERhDtYhmfI8/EfOOWr22IzTC0O2
+SX3jkRQBIxvlw8EgNkTXm0XqwM60CtMs01SFSzrCBM+y36HIijnGaAu4l7Ev12S
DnShK7d8yT4OeJzMRE9OT5vGFDPVJ7XTOMVA0ucl2gDlqrl4R098baoA4rGUovnE
311er6lg2hmMJfdtl0WN3ts7GljOnawGBFTATbMVp1E+50GiLgTinPvcLmN5ph0k
HiDkSE7dAwHsmReFBjBsRHQIPQ1bCxPUM/MszOR2q6Tvucl4SxNMNKG6QfT6byfu
iZcaK5KJxPceURmLdWluSCCkC00e+RAf5yVBNVznweV/+nL7dVovSUywO8Nb38ul
nimhOWVh4dHdq63h7ForDuvQ8m9nkSyyQj2sF8JKX5pWNQdfTvqSF1azJ4R2eC7n
WDYoPjXTflUwP6dcdUcVSUwlgOPfL/3OxdbOdLCxJvK6mSbrZXrdaQ9WYn0xag7+
WxOySsj8Yg9KKSora9iDRAYsOAs+fRyzUcBOKKMmT72fRJj9snAoqbvd+GgQ6x84
N9HWYnejYE6fe+Oonimwonrf/6o40kvCLNVV7cGUgxBQWKvBbyvrUaxl4NQV1i+4
Xx1cz68lLdf9Wf/UwG5f9XN2S8Y6h4DTTjFIafNOI3NK2Lrr3Er7QyOTkII+HIDt
KUHN/YZBCxwBpGC5rBEjMn0TCmM5rpzJ5ShcoObF0OfeaqMNSA2xltNzZcgOuS+z
d58TJxJ79b3GxzDvPl26tEc+zmi6nDh7I5lQqmE+DRjHwEspKeQ0TvLTsV4beN58
yLHrCPgeOg8Wugnk0IQIGmlqWnSLRc14xb9donYf/El/00Zd+ka36rLcOWO3KBhB
ix1wMuYCfs1TKNdvVtfWAZrdGcobyhRK1YGJA7Xg58PvhFkTuOoglbydDFUNKXci
FyKoS8oSFJgF9B9SD0SFW3R286vSRt+fOzM9UnB5lsS0UF/3YDjxs0QneZCHdd3k
jCOJT+mB1Nj+gcDDcwMEs0MBsoR8h8tK3gldZhaCAW/d5lpxyR0Cs5LE7RfD4n/E
5SFAHqP1Ev863GFgcohgKWpva1E3K550REvwMDqEw9yG75QHiX9xJh4fuUCmGLVH
l/mTpxfVtjQ3vg13ggYcGYO3LOBdYEjf8r+Q3vcRZW7qDqkqSie9k1fTkp7FhrDf
boxWdjVTWjWO8dA+vy3ctjtN9TpcGwphG6+FrvKx1P8hj0zm7KmxmgtQx9Uaw5u8
OmO1tq5W3piKtg9EV7r/7HIekGzf7uNcS/byFrgZcvkVZCENhlOaBctPqB4Oi9SR
W4ry/HUawbsq6Gq2mrUtSL3PQ3/sfPx/mtUKNTPJkC+nT/22yr5Rzd9Xx07tPoTo
qv85CCXVSBVQ5qkTTJ6WizNvp3bAva5fPZm8eqLCi/x717ZCguu7vaMBCw9P5YP2
jmurM5w13EI7pElbnWXJQQSSjsjX5hJhBZI1XoNWaLuGdTlNCHOipPez9Z2hStgW
4eNeO3q7vWUJBzEj8j0fjCS9Pdf1mCTJPMsQ+hesmr3d/zaERsk+riPc4ZlbM8qr
/aWTo62oL1z10WAD6WURHUmuLfyCheOSDfoGS6bvdtzTFlkgrNp3g/L18aZ6mOkQ
EB+hBfGgsY8zMATk/5o0IYKrCfYVA/5WCBUpkLKcBt/16Fv3VixTj/q0xB03YsGI
ff4RVAqtmEhQn8g+qmLUPOk4Fys6ix/0jeMbo3xjrjVi9HnDApyBdsqNKaW+cBoe
0eVldfQ0YwrHTO8nk0v9cHKjoxp219tzvr7RLl+WKV5yUgII9xNH5daosg+3B5sC
xlBSedB0vK3C8AkCDM8y6wJ9ilfT4iaAd6YLGIfFLW3XYpQau8pJ2MbYMS2cGTDz
IZ47vDOR23TSBaz+ncdF74GqzaTidaGh/Zatp5oGVbXL9DGok9dtnHgxx2MF2FQv
PZNv6uztzxDnRylEE0CEIBckzcHgoHleNxFT7z1iiReUfs+5tHM06cx9zrE8o9E0
Rx+3aN5LxpA2o0ekdmI0P7Wyu5YE/lfmLJHToWNy+Mw4cHkX+w3mOFgHFKL8LWGs
Iy3/r0d4OejZ8N48LdP0fE8jQP70oz4elw7C12zGcKU8Kauvdq32VIaWkCgFrksd
ML8vy0key6md7thFhKlJYo2oVaIIJF0mQKHNS4RE6v1XG/xfeS3xC76vLFcE725y
d0m6sUfdMHsMqRwG3TwMzEah1QUbUv+smrgo7iWDLMsQUB1QZakDsInYkXXJvhzD
/ShNmcAn6Af19QHyPj/Z7BjALXt2X4GYOLI3TvDJ7HmfkYyqE5WHoYKrz8tuQWgz
v/Qkvjc0cO3YXbrV2M73Il8FXHY0n984upkZhsuaCDltg9DOXqBoceFZ8P4XGhQq
f0smi1pYmfrpQx/F2aE1IyOzxO2uznUN2Adhu8CyoFIbItLfVY3r4ftBFQzm/Rqc
+TcVcLgDFLN/U44Sk8Oxp4ZvYdaOKBPtqWToIAI/rCBJopAaQCLnXiWQ+Vp+n/xe
FQTyetzSnVo2PujcGjgjgzQH8FlE0XEhF2G6t75FFP2QVd9R8Yjprj1NKq8ZjsPs
KVItdV6ig1Yy9UrNiMVGHFy7w3EgWvlMQHav+Psvljdc+VsIAovPXjaxIQ1L0vCp
mjOfXW4E1OVjiji48RLC95XxA7/4jMOHMqgo2u2vbQJS6z4GwrVITxhfJr36w49Z
fdG+jKXEWMujPgFArUKbf7Ik6+ywzOLSOhlThFQRi0lSJnsTV/n/eGimjkmEf537
aCQOGz6R8P8H+vRSdJtISG64mECOzvjBNBRZLQ7RThkmZ3TXigj09qZALsFsCVmq
KufTJvRF5sqBzUDpG81KgjNiNrx0PWBeS5XdyjAcRh+0qcZkt9UYMSX18f2G8KET
EhGL0D8BZtlz9lBxM09GAbmClto82/lrJU0Ui9uW/TfnqGiMfXgXKvPBsFSMKca0
np/2VY6dSVrFqYtrbf/TwYXdbYwW/lg/qhd+wd7zeIhjWAaEDOuBze88Zseha9Fb
+eXut6n20aKKN2r384FBx5ESgstJW441N/3dCQg1GStF/7g0+1E1xzHvMlZk0HCb
Bg43z/HXo7rX37E74aJ3FRrluGXckbtX2GNjcFCjvtwruvIMEKyPD9hA9nW8b/jU
usHv38QRDtd/68lgBXlXE+p9dCFJO7jqKVP3xEyr4sL9a4upIs10RcuMH3uCwqb5
3ltvxYjtS/+B7dm7bDsjVTLYy1C5F6kj4BTEDAhLfQKSNt/OoLq/I37MWVCEbPXz
0hgwhB7k04MqIYiUvxcxlFvgjJSzDUdaZKPa5wFX0t/2gT7JhhhCkuSvDVNeSm2N
RRDysyq6lZQRiLq76qKkFVqu8xOxDVHNds8vaflO8gnWuKKbBgyy55mTRnOCBq15
5uB3tFf/JeFR+BRvnZxXmUuDBShTRTWk/F5O2mO12kL0TZ75ZaBCBO14aqtjCNwD
CXDZMwWcETNh/WVAHWyJQZ3miZ9S1WmWOBrug0okqAEIJ+nMTx8TlKIK9y1N16h8
E3FtM+dLWC1+DIa4SB9AiPMAClkFEp16ZZhi4YddP505Kh0oHtHnB4yRu4DnRQcA
/ycQ5gSc2LjpOg6nMqDQPXCPPQOIbJqG5ucRIbXxJl4Upl0ereFhQUklQwGIQ90p
CF2xcL+HOWYi1kRp9XHup0QYFvK9oHolaBOVBSEY3faDRCTp0p3MzXJb9P/AWklC
Z0yZC/pel2L3qbW8UPtatxBL7HUNZvkIHKnO7eYfqt7m6Oc6p1hmDYa++g2FnBwV
iee1F9kC8xgKGZOmID2vBH8eAvKD4uTX6kKVIx37aLVyW5f2HZBJYTbSNszKcQ1S
6HNuYHMgOjTPnnuGk0yVIurmLY0CvDcROpdKVgQ/2McbD7IF9YbEUfAaWB5CIKWJ
CWl2LQyfCZ6aEo43xZuUveBpZqDz722C/cEVC5TDaXbs6XmSrxfVEw8XMxapmKd/
8O++8WNBJy8hfL8tSqYSDjnqfP/v3lZowBpwrKzobL6TIFnAv66G96SFAoIexpm4
H3h4oR+Qhv4OoVQdeohwJOeiniSkfEztzTKX+FfAoHsfXwSNEwYWjruH1LaSWQR9
4QzLvpL+I1afV8QhsT3aNOANySplQeV6FcZFJjzIvpbx8/Yl2QsTG209LK5uxBrO
BesTRAmkW5A5PiggVlVjTNZegqlNr3sWeCr2t2x8wKOFzVMoko3IaNmTSnSbzHKB
aq9stWVimGrzALnsMzENzeMzGtFtRCOjPOoKF3ekoiC8GOpuzQe/Ur77bFlgCB0P
xVUbwY11sF+7JZD3Z++hyFGnXKIKz+0pdF1YXIS54v1UDNe8DJUz2D6v/pM/wdkr
nAeJPvgN5nSMZPzZdZXYh4SenpMpPhMySjhQXzwGKDoPpu0kP1k3bZClKKotGRDa
hoC/9JJHksFVK2m+djWglTCaNISDNaItGqgVUQhcM+N8ymCH9aogofwpDgFxGdMV
oepFRkWfgoikOcoxZlwC4K0nrrDBfjALcg3bujc5GF/r1t26mIT7SSrOZgNuzyJ3
WngjOEimI5e1kvYWaH3oO6NQ9EuJ/q1hpkjs46Lg3XOw3cha0CxMXlCf7xncsLB+
WGtyXmsiHBUdwdqfqfEWsxN4uORbuMVsp6aYlCXOVCBvWBcXFkQj0RKfTlAaXgdd
4dt17KhmSw+cif7fOINsi1dQzyKugpeDQ9K2svO+0PRIw0opEAvTCSPuoR2GESUm
wD+uhG0aSqbxQFCjYqBnLQNy7cBz7lg1/myif8cbHBSkCdZ60kx6CKaOMEjq+ppT
xjgSAMW42HYzTNwaKduGyzwpW/1g77GGF1UrxJPqnetC03/NgmOWBIclUouEIK1L
+KZTCndJZi/7vkwcbMVh15OW1CzDWy/uSyS5usQaEu/Vkj7VanWasn31NIRoRhwR
ahXKk0nKPSS3C3W52M6uI/jSOI0sv3bQ+rvMePrOeDQkQ11W6TsMfSTxq7+cR62e
FmSa1ie8WnCjfp47RIxhgWhf+PBi72Za4S4TwoeKEDYbdxRbQi7nHFoo752gg2Oc
rokt8J5EVHMTJ3u2pZEYZzADgpdHZFjYXQNzC5LsHs/A+8/r+NMahDYDYcZ1w7wW
I2SsPYAIrZs2DwwoHA+pyPuqbcnv0MBZ8WdJ3Gz0yVi1aeazP9Oopp+wVzFwfg/n
G6Rfg8RAteDbJBJy1HE6lzOMk5ivJjMGWOkW3iAiQV2UPfvCMWID8x3BJpn2GH9C
O1hkV0LAMzLpBDj6Qcxl/U8HpgS40kHBNzWy+C+4/rrXxZoQQMMGXPaE7MNzJRyp
tRZq/alpf+1UWGPYvVIAAXBMct8p0/sfR3mOC35oWuXOTAW1dxJHohtGCIxu3A7P
AvO7sW5J5P3NyE/tfYoia1FBzqNLgyC6fLyhFtQ2BoDWGn+b/KluE8on9q+/i7S0
sAgUD5X4VRovzrmLRiOyo/19C4JXvSmv5LIOt1KNcj6wcYWzwuEjn5gwHJbXwOKg
ArPhzuITCT+oXf7Q58K3wxjgGPWRPL0y34C9i9n0ABV5ezkGYruPocJC3WsM2TJy
Q00Hh/I+QdSpYcH5UePOTPcJ3CsM97PqntTdMUhV6u/zrHwba/kyF8mK9ICboXQH
cLxdSIuJ7CNebY8YUz8iQ8LeaGf9ywC5YWampgTrRdDbBGf2UeocD07Z88YIvZfF
1gYdn90DAYTXqQOeVGCSNt04zUuJZdAoMP2vZGHeFEHB6638tswctHy4Pz1t1+40
oOeCSppvYRVkNgRf2EHfEZ+5QSxpa3LA9cDPleWXg1ML2DNsgx3nUKy2zLkMVCVX
R7LgQL8pm4qMB//DToQSNMp6sywhbXBVW5bzAP7W+Ks5zEvdaYMpvpk4jZB1v08I
SkP6Q87GLKmSvqurrcEKtynNxZKHRsXPhm3ugEIFE82TcAGCya6HZhAs21P8J/Fw
oSQ9V6a1gD+ncWTxnrm20JRN9h9bKr5JPWhMuuWCWQYxP4B+nzdpqvqWlh1fcBMy
Pr/UfA598Bp6p2X61pIId39MvCBUgbcagyqYt2KSJYxWOWVDSbM0r1RerIuT0UH6
DxFLHY/DJRYfIIkmxzkj6hbBEM7Eb9Bru/mnN7Unw33CfiXvXN0ilqpgBxuWcWG5
wemyxU/LXT0LcmWdNk0GLCcSCAs52V2Wp+kvGKH2aUsT5RpyQnQi4ioKg+JNrDNa
X6BLfoQl3E7TRpVg26T422FMXDEAo5JAkkbG9s020oszABW/ytaP3Zp/466kYVlJ
eUKCh0BCNl0YVTD4PSJGd/P/FPlLThL8Q0FlIjIaBClqAfro1VDvBZ68G606Wo1Z
Jd0E+LTflEQr/eFaUT7wMj3n2sjg0JcMvAh15QMCgHjOPgQiY2cW+9XHG4fNR85K
9BZB8u5EAlK2wn9TTK3yuyOFNsjsB5Bk0wVlLjVmZ18tQiTkndLnUtrLF1eu6BiD
6jMaBV+y0bjR3TW/w+GT+phOmpLnlDaMijLGI026FITXsqJczT0XVK5z3cBPfLoG
kRgBDKfKCWfUcQWyGwIOwYjd2mi+fKDmkoiEbhH/ngwp/S9FgjD1ep7ojluEH2tn
f3oz1K7GNYLfiKTS3L410JJVTHfu0lPRHXh7uOdQMSIxFtOgOpF2QDvGvfWQpapR
17qyToFU0RvUu/aTnIEixL/j3UHy8y7lY5zUGJXVgh8eV75GUAmT48w85w3hXT97
IZHcRGruqPtquv4DqXkdIUWFPo7IJ8uZxmWkdjoI7U8gJRMbz2nUNM4mMBwaraWd
yWXmsHQBCxBFXzv7FoaO2Y8adE0NuWnmaYcRQuept5rj+NGCv9hkjCfBhDSN2dyr
Ikpuh6GD0FurBGGLDNzkoj54R+6oxC3LE6YZ84J0lH8MXMFi+GtjE+Y41dq4lXrc
SDL3tcNmIYX48pFGPI7nfPJsVyt+5y+Q2DA88T3tQcKamaVyCdR2DPLrKTtMKZtJ
FTon/23atYuev6Qbm/FCHR/0Qcv+cPMcCB7nGUPSUreHeO9RS/nPiFHZidm9i+Au
4FAJaKMR3E9OZ7VpSd6EBjBakxq3KruO2Exz7TLScOASALudAZpV7O7b3P3Xf+rA
A/sk6FHTgpHg8gaVb72pJ+iLEIk3dP3hhHkkcLennRVtAgwJpOvJ02Bl9L2hDmEm
XgYYY3hxSoFaUEmeafOe1Bk3zPjMuHRWohobz8ZPsTIxf5bWFsK10qs5U/RP3sWs
1JJxthakpjAopUrkygzJJaY4RRJhiWa2RWeSmwzPWjpzDBUCCoe9YhrP8WmjAD8A
YWqlgqLDJoe7ZL5P4+9kXVNVzE0Sl0U2nAKWNd6wMJOFIDo5g8N//ztKGTaRiBBU
A6lUwjzpbyN5pbeLch2QhC8I0v9Gr4v07S5rTHrK7Kd5XjI2fzifIpHtinZWevnl
U8ck3UWvB3efdWFOQSxpqobTjYJFXYKE7rJczKnMQx/RwkJ482TWb961gRweBMSQ
6DLomRwDDU4BsIGWZ/RXGO7rThnjqflgKVEwYf4K3X0OkE0ygCOckiVRay1x/ZQD
kDIq6Tjd8qn4dOnbh+TO7rPbxcsTWbY8AVGGcqY/7dCced3vczA9AfGLR38TeaFd
aSITb8wIob8sVUerKbD1h6a3lc/3L9JUGzZVaW/uwLGYM3wdS+YQ9ExLzjuMfzeX
rfftp4JtoC76ptxAA/aZU31EDi1UHO0tEqd2lzOGON9fqNS3W/ooSQ2CcQlnVCmr
tZCXKyRizmgL9SG0hzbe7cLfrkJ/2zz3hhzd8gtGUiIYf+3Tbb79+bJDQzv7Qngx
eLhW2ChwX62SPP8WIoZYYbNakj1Uwxj87U1iGiVi0j/f7N0HUAUgJ5C0uL4TEtCK
3WO9fBqQtBpW9AWUUjKScj703J5db9DC9tZC/5iatDxPhiO5+fqNxtXw8/Rprxej
TS1voM2+w/XsAwAGxX5EBEtZpaWdiftJ+qv701/B6Pbe6wwQzNBmd6U2gxOuPOXr
/GYKIIE62MbQplNt8r0D+AAi3fciK6jY/Q2otr6iY7j8eSsfW/EZzPe0F9bifpQh
qstA5ZB2T8/AeOkarp595kuBxWeZ0N9m0ZZRtVu+3jTdIxlxdP6BGPYTDxeSbPiF
v9gv/NSBjbu4vhw7lLg3eMtSwOyHgPjm0Ilq84tM5DuCS+AZappu6UD83VE3UaZF
fltEC5GD4ZYuf9wF5whDK9O+9xXPCyvrao93SxOftvK7lX17vPE5r3vnjJv5mpxj
4rucqvXwrz39SZtkaYIhWf/Qm4RtF6OSUvM9DnaX954JMS/GuZCVPAnsqddTS6wt
vOWJ0SCdDLF0NSjqPU301/8tbjwfIMr4Bs2UwPMmxiOfEpuDgJL8x79P77jX6nHF
TgfwQRFafRlk/5jwoeGhBlGbvqJGwQx+wZiErQJs6gN/0lRoW7xHj5xUShSbWYrl
zTGmVKaatt3FrtXl6dRYZ9lxuzG31S7Ao70BWCG1Sg0E5aaJcRQ8zOAQQShBKLYH
MMdnft+lwNmpB6hvNtFEsV3XgtQ4yRaxL5ul+jvgoG0bxluPHY/WCvknF01HZ6Sb
tfumQInFo093a7fspnMMmF88v9glNEl+/wOzJFCM/roocSSqjN6CLIoOCej9Z8Gg
NN5DXmyfdBzFhD5qozprfF1yMVhVyzo1AcMguYPwAIEEJY8CJuech3ibfPRq6X8J
7aknLN0MCe2U8SOPZM0JsNrEfBiwY4fHjWXmF2Qg/RwSHDV9711H6RN7OxpbXQyo
sKEVwdcMcThYvCSwfKkiACFriTg5RKHMsh/VIEwxRT8+2PqV7e/VatPfEkd+yQIp
skamoSaG7X9ZYvzsY01Kzew0yrFwPn75QFoKQpeDLAeog1WSFD+FJg7xp7wcWMQd
dSS13KPmRGNt8WlDeJcs1BZlxnBnWTd+kWbIsaWXiQzWZzOl1JwVY4Ex8Eep35zs
SpGBu+Hy5iZdbNEZQrUf2mFfwCyC8FSXZAnRZ14jQfODs1vZKNGtGi3hptWKiT9Y
Mq6AGZ4Jv/vLvur5tXu++yoPBKMfptSsvYPBpM4zr/Vo/oThbwT3jpyO3xZPeYp3
vTqqCXDYch6HvV29lT9gAAV4LvSow0Ja07HdXrn/kO9aEN0ytP3aP9/DkeT0waCp
ijOV1HUJTFEFJcNB0T11tNeDVz2+Qt5Q1sg6RC/RL9x35YQKZ0NFBeIM76QXKJfG
A+2GTIfnZ/IfGXPB+RLPPHi3cmy8tKRgf5Sq+ax0IYjCWBSqSDLfam+83+nH4bsL
wRhAhRMIrgYmKJf2smb1ep+eT1W1oJj/aLG+uoY+hNwiKMjAiCtRYY2TiYxrdmY+
wU7bhxKgTV78u5PIXsOgRTSF4hTiaDYpIqBFsBjUPug4kv0DPaaRQ9pauPYbyuKS
zAgxnPva11Wuk0YUgdhIIRpOZuRX+uY1mL7Ilg2KGumPMDUubH+XKfZRpBPtLp1u
Bf0gGQFjAj8/YuySmTrltV1Va/LPmArJF8YXjRlM86P8zaeWi1RlMQivQUbBB3RR
gLzAdImRyslIG3mPd5BGh2sWuAZFMxV8QodFcPzuS9dVoYBtyn6r93E+KZPSVtRl
DrCbWPrhWWpJHGZoKCNZGox6gzBgQXv7bhb63H9ILqCyE5RTcWAYS19xm52W5fTp
kxN4/LFzeR8dUA6ovnHb4+MKZtNUcvwYti2I1IgDNi2/6UWit2RiCU/U1P8DImo7
73QjhohgRQREopvGFODLJx3b9nts2Zi6b97ffgGmLB66UC8jB/u6cS2sKh+qTg7i
dCpSegM03kGgbxT0LZJ8ALkOCm9O3b4itB7uFD7A3bXE/zZPy5cktd+TgvIx1KAc
eobD7Apt0E3Jthsb8rk+ercY48VM1wkX7Z6das2uG1dngvSRZCC/ViqBFdDt+XX+
z3GSUS18b4PtBtvE1IxYxKVO/Up+psCrOCepGd9z+ttNJA4dGrcM/OMAU0hE1ni+
XTP7D5G4jBDBFThd5LHmLvPiUSLmPFmIABapsMiV48KuT/kGMZVNRjx3YyoaTUur
I9bFz314/6YuArW9JuMskOFoMnQ1CkmjxKdop8JMRmvjPREBOkyP5U0ZawnfZuUo
g2RR0y1FP1xsGkhLjKs0rqQd7vhsK42wIQdS8rj+ofIURPG1GAXwmH8AUQ2FlSTu
Vbj7iQpJJ/tYRuG3cH1wCNPEno3M58bSIRzrq6GCGYKyrWiXgSexyfQjBSjXC05x
/xYLWWqBpaB67fOq3l36nu7pyrcmocXxO8OiNjY7UpeqSBpbOF1QMuD4W9SciBIK
yBqBh1/bCf1k0MiYKrRv8SZKW/vQw5q/1BiiJ9FQysDVvN2Dx0XA+DZ7emSTmUeH
d1HWgXC58amy+eNQfN5lDtglaiWVzjXBxK5yHnLq6p80I6xd3q9X8FBmbt2fE7WG
bywnYRPstVwAvI++uSuHLWNyzgqc67EQUPhqP74QgvS0ys3ZhAve9azi3DlsTqjC
8ERUpWBfy+R/Po0obDlpavru3NzmiejHGXo/4+F/tPXDKBPGc2tiPoS2G/zxES9a
Myn5HSDGpub0eBHr7cY+YkVneoexEzEzukw9af0gAZMtc0zetE9rYzBnJBHEojNU
AOTYDTK+V5dpk+gBH5fGbW9bHwIpgAorvCoBhWH474EcViu1KWJc7xK8oJLPohzc
mCNfoyLmP+WscJvsCqOZPsCUsH3Dl62COZpqujw+GfzdaYjE9HQLPASg47pI0Ctf
RoWX0vBGFz2y/8ZnPnIX0yFmG82s6kevExhyEPMiOTD0YrywZaGN69n7oIAsRLrx
HMmhCBshLYyT0Va+8KwfVo3NdwAZKM1aq/OhLNLPhoMHt9QDByb5kdA9is0ezFHB
sNnL/X6SfHj2+LwwLTnoE/A9ZPhLaGoJ2vS9jsRZbl9LtalVx6j9atjf5XLSiBSb
/u3APJlScUlxxJwDXQkJZBUuKUjQ/518xgFxj4BrZ1z2WkWY6Ht0Xy3yhx11GKcw
jGLGJlRyGU2szap7iM52gbwFtO5fUoGva3qdNSX1TCU+pZKncg1bop58j7NooDns
pTKPOlD1g2oH6RN5BoVKStVQNKKi07MGfwCQeyGVVydohA0RKVUJIxnyu0iBMnDy
T0c7IAOyl8ugYWeuRv67Qittyg18piQU1UegXDheTNvug6KrRhEhpnWWHO5viLj6
SgryFoFtzqQa3xIJQFl6+ad7r7aUoueGR2eUVxObRxX9T87kBWgrDEpFLF52gARk
wp0bB9zU1g1qbFfK/o4AChzgs3nclZXXINdi9KZ54fgtmPnZuMgQ0iitmmf+3ycw
uZ7g02w34EnTEtvsy97hzsRgr81kt5kvSNHNQ2i/biavZ2ZaTL61QWeCgXiOHebP
67UlNalzDJZ1iSJL2Q0Xuq7Aae1ZZsnRa/xEs8Ht/eF8b5vdcethQhRq94/3LgZ2
0zD/TO/mZ5w1lK112uH2qwguLc9ubemvjfMxWoOXZySfokuuv4OHtaJxXRPVPBfV
F330fsn/ysTT1pNm/nDdNctVRgYF4FaAg1Iqo3kTV94WO2V9Ux3rY8MgaMGzPwgM
FM5aL2B+xxpTqb4kpA45NaVVKXzbt/txqVzcwhQMZvIRiNK+2ygn9puqcLdURRBp
xIvQWqBxcEScVWVv5quqAlRBxhTGtyt8OqpQb7ymL5K9Eh7pZe+KVRi63JIiXCsE
1lIMhdJaY/eUf57XPhrbIuA1nlv+vsetanXnlvy5lVUzpC2LkuwiD+PNInjY5f4T
n/N/S+on/5cptz4y4Frwb9LTYulvGPOY/0DgxfbzblAkjM3cK8FkIRr69I8OPNo+
2EfbznK5BU113J7Tm466vFCp1iEx/n42d67CYV1LU2jjkBJGUz44Xk5mLrbTPEnh
9PF2wPi3tuSLtoTnEYM4mseAdQJc5IRck+AWKvd0lGcbMx52RRYv6Wq0CmrTssgX
NCqS8aaEGj8HKCvQFVElHWp74sv0vnGeB46lqq1Nuc1gJ6EOj6Fj7lw/jxelxHG4
Obm6i0T8IvhY+7eP+KzZJQOzH69NiHiFzb5QyiY2yGr9RLy9bNkA1YjTm4ffIwkz
cjQRHhKM+yDNdbzbJLAtmwPARPlzSs3UYXrWrCG7Hy4aR/dZVpmipERNEgdiFohf
OhgMMQ0awrHc60CWgOTcm8gKKcjSlmecr5COlvBPa4r7zpMwHivRmNnmDjcf1w8/
hKmX4cQDnQdXXVRcOidRKZcnM4OCmX3LtEDJwCsD9cCquR4MYc1nPbx4aBscCPbO
xa64hRvHrQseeIG30bXeRcotvsYNDE/Dpr48jZ/ZW4isNkRg+SutiQkXI0vQQcYN
LPqpqp7CxNb2E+PF5HPkbkuM5Gw7+fiZA2lM6FWfdWdwl3KX41DDxel8b4Vxx+74
sepLbCgUdZQCUALWJEA73fWWlEM8L2POpfseYGWzo7lJhv36ane0HbQuxKb0doUv
XsarPq+O1URJ4jG8uRqgQqPDx1iVgsq/qfC9aKQkaC9jL/aLh6TiRmiJODxyJ2Rs
P0lmAyOybutHBjR7b684JUJG+Rv8SJjJpNrRo4KcIUmpxQxPl2iGytnwqKkK+IeR
vxIENOU4igecYT2DtYHyAsNKN5ELGWni/D9nJwlArw5Emqy89lfCtTJ44YseZaym
NAClkQ0oYfAaU2t4sx4RGYr/Hh+zjYghXFD52kxL8LB7jWyUoTOBpcBi0/9SU2Ie
6lt0ICl6u9OP88xVXPOBMcFXobUGWTunCfMr3oDdUzph1vUirrkSdi4RBMrMBuhj
8zG4j5lYqrgXea4JTYI8F8Xr2pcFbsR1bfthUQfNcweo0JHNLZ/L97fyCPG6i4xj
S9f2fgrb0sk/viY6pNSbNXqotczU3xwzF0EjDuW4jv8407aDB3GEWboosJt77BTU
eV7UfJtEiD4hVI0LPMqb9R/cJm4CKkBjypT/c/AuUCJ6Mxdb5stkArkeEd2BzfVo
GNNMCC+PsOQBNjNHOliV6FweynH75uP9Ug61hATWe5weCBVoiedKKAd4JmsXtIyz
DMdXEOcAQf4asXHFPHzgagm/JehwvlXFfx8M05uO58PEZMFHfNkGM6KcbXHFN+/m
KEkhdrcCZZMj7SyCKTMPM+5fjdVVAfJ004zQDcjGaZZGxn2pG2y7R458ZU//KT2L
p0kGrem31B7fCQNwhXIU/ifdH2MXjGeQBUknh1gkcNDy4m4EaWP9MMfW+UgenNKO
us3NC18fFiKi/CI3fg2+bbdjcFa4hAq9Ha8RlJVSSN7v/S++A4sz39qeYBBazdB3
ZXdafALhcUHbEdxq9CA2SXDtkZJmfQ08/yL3FtwmmGj8myIWGUsWo2Q8Zz4I3l0h
FjU8hT6biHyzXd9257GsHPf+BXoyub8KGewDcps4R6MpB/luCqueea02kegheIo0
szrDMFEwLmX9ch6Cm8MOC+Q7dTbxGqjApUz5qOhCwIdBj7oxwuY02gXh1cvg8WD3
8oM6AgkOQo+C/+23rP3/Jwo1jj3j7u7CpSesEycoYgtPS7OAJTbgWFLRBwwtm7ds
4AKl6MN/39l0SmmBc1AN2TcsJc1xAACis3VK1lWjFAzvnDH+0yIrOdItyqmM5F1x
eChyMPhBiAg3hcPRVLNiassn0yNqCZ5BB/PIs9WQGGpBqDgKC8TPvHJR55gA2lpf
9sgSeOg6EBl4X1tsYPu0rdf91nGolFJknSmynHFfpbVvhT7YfDsR1s0OruwFAU0l
T+XhdujaFuG2dxmDp8mhG2DLm1jO3DFaq10qnqZc8TqqFuYtGzxUaEAZDHyXt9oE
pC1YU8IE421MKF+YJQ0P6fS1A7SYfdqAgjqZdt1hdBaQjcbjtRRnU//vkDt5Jm+l
Pnhzk2PyvsPlS51mhVETSKqsIDnbeVbUXu/faWsWwuWHFO5vyzD8p7m7RMClK2J5
nFwxm5uMFBFW7rYi75NWn9ehRVj7drVXox7b07W4krFnhY4epr2vm1bv9tAcSoK6
XKB617to49OnFkS1pg3Ruo9s4Kd7lxtnLDW1GoLtjMJQvE2rfZfoz6VqW6BQhvgb
5f4LCtvOZvKSnuAGWqYzs5hXBXd8FbGlnKsuNvZBk9sGIYG5MQsOKoFGx1ot64eK
XfMND4KVuM9nijCCm81MOqNUtA5hcs+tKgDCKSP7ac7Mdxj04ZoSj9VBUwxELAI4
cXFaWGQkyaKrR32ua0QjQq6PrDW31jI2Zp7kTSN4rg60VJuFXud82sSt6oO4jFqa
IOvsLvry/05GWTLJILl2Z3CFaFwjfsK0FPpNJSyf3WyoWlwfPEnylRlwMb5E3CEG
VSI4pBH5eXX2neet3xwZf3vx7vSuVSu0YC30IG4KtBW0e3+AqbbOYvBefR04GqWj
rpVJdAC6mg2jlTX0YY3/71huEIYVJoqIH3FFs3UCMzC8XSNOypq7SFpZ9bEKTmys
gA154nlPn08v5jruhBmnlQn1M5XKw63ySKp3mTZlM8hxjDH5Zg1CdmsUkgoZgunS
7mUNJS7+2WHzyJSUh7zWf184M2EH7hpUsh+zdfXn9YaYRlcpycmgRPInVtM4rPna
GIlxgFK/uAn+WXArLmq/RFfKamFKmDXKo3C9csJtaNW0HV7DZtplciusekbuSsJ6
WQS+iHwhV9WZQCS+c5zZ9WUZQUyfIww7y2+xe3MJ9SwXmHHPk6rCuFQiZKgoD1bA
YB2R03C+Jy9giaYvjqiuUfXqQ/YUFVBBc8MhL7VEGG/OynvWfVbjaxPAf3DFj5je
0W4Y42bbMyqgfN1ZWRCnDK3tVIkVyqGXvnAuvr5L9Y4BrnrRMkyb7C5fhx1njxKw
BN3Bbz8apZP42oiD6xVKXwnbV0E1GNLSB10aSy8CtcKjOXfkuhyIPboas6a5V/9+
Bh3/3sb8DnKUvFP13JqTk02baRjhRWtu/82sSBXVOBZEqLxdPNXqrMLfQawaIksL
hjZXpxwYPslTilrZi+dGsG7srHr3JNiVOl1YUIbSgfZ3gdkV0I9J+W3U2VIKvAe+
DTWpAoGQif5CIv3JW3wdy2dzhqyGB2FB7RQfy87OmRCWObgJkbLwKVUHQLZh+DrM
ZPdv1zA1zyl7H9s1l/hQv55x8LhKbSoSCtIcTSmrPqD3fDTjNOSiLrkjJnKjoF62
TU8LdvaeaDsDuH+IQ4AVSFc5GffnYsqm9a4ljeIq57b8YXVzenIP2OQQNNhRdaGV
/CtXAgNQWFTyvaAjMI/3+zXp8d4wO2wjxOfObvSABgLB4QTnjJNAxpxFw3pdvNUH
TDYouAIO59D28xF44ZdjwYFuGzq0Rfu3VKoNaZADaTOe/ePYahqovjcwMNOnTmpJ
tP2+YNgc+J//wvPsJxc+tR1DqoES1LQTLNZMBMJD1l3knPmXtEqyxX8lm4Gm7YCR
741xzTqtIvvE3K+HMUMFtu8K8WKPp2kc3weZyPi5GaNlLbFC3tOEWOO9XMY7HNDT
b1oqa28YrFK6Rin8m5Zt15OUgAYXiLP612F1QqDvKenb6mnYMNYRhop64DNSrLB2
YE+uI+FZZrMSeEJLSc7qDHD8bgOCiEsrpyj8qCwMgFjVHhvSWUfIwPp2Kk6mxmC8
h2MH5rZWFF8kZmDopR4KhdvlngCaMKOB1nOoXvoitO4/T3f+UEPQAlbNAEClFSA0
NzwN5MC7e4le4fUmFveCt19CRLVJB0o3uo9FC2BPF8RhkKlBpZVdTOn5rlmA9SZR
dweUEEOYyxUNZCenaBdIRh9wm4j841KA4q1BfNKobvjpRzg18Jk4xNknj3RE4rfu
6tw4KaryQcoyj5NABGCuxFUamqA1Zm/Yli7RSX33N8IlzsuM097gODOFkyW7Jg5R
3jd9jbCzkctpOY6k0AhX2GgiERl5goyc+3xHTqdOdkts55CTt+CW14KZ5JU3Uute
lwbxfWKh6XUz1tqzaO7pl7qpkNKcTGa5d7aibsrVx3oPG7cQZa58gMnViLqkXIBn
6wvy6g1lTf64VeFzj7LX9IZsdFo+2LbSW5p5GQ7GhxOCi5dsKOK/ddNUcN0Q58mn
2h0M5IJYtHTs3eQLBN92Sv8ymQyK1uGbZ5/rxdsb1GtdM+8fQhTT3Odr6lUy2ZkJ
JP8T2oszQDfk43Ft68X0gjO605Rcn144kRMact6DqTA+XBdAY+6p3Ym1Zfs+DcQ1
zB9TlDo6WbqMvsq0E6dvetJ6tu48M3WyLGF1uf5CDGJWNwUAERRrgaOHEiut8sv+
27OOi2OZGaGAHAIPe6c3LfESyvDMRiDPgxtOZO0no5NPvsoPEBhaQitI+MRGpR1D
OEYQnyXQ9zyoh4AXmt8x+VOEgNcmUQLZDRTmuyHq9LCgpRqT6aRnoA9MmsamGuD/
ElEmqMRHD8gfOe/v1XH4UpdHIXP62w7uySOr3NLxX5/hX82ViMJeYB51RXB7/ded
j251usxlantA7y5CvLSAybYDRJJtfZFE0GIRsocqhqyZx2J7bJsUM/tdekpjyryC
pzsT0306KK4ao9738aSqndBrIIwEu98QmeaiVBAlQY9aDGUVHvAAjfjnElCYm8aE
0wAt+PUPumnbcfsG5Cf8DsEV9umMoVuOvbB7H6ptTzBfBImX8zsFvDEZHM6t5gRE
PSsRplPRV0rB135Bsc27HdgQT336pi2FpbbnnrON2yZLPjD9KnrU/ihGes3D8zYN
ZpDgAT/wZWvuka4lO7Nd8i78l4wEcj/CbTufFbH60Ya3WTkSByDGTU2EpA56PXVo
F2ZuC5SyczRM38kcC+RJwvroGenxmdoed6mqb9C3jRtVN1Tjvx9Sg4Y8lLvYgvlT
fDFd7pYVQJIjQM+bQCpHFkm7Mr/rE9Tm2AGtPu9G6XsOjjGtYK1r3dyBDfTx6D5E
MRCr8D/TFoerxh6J2K3M0zuuXiWl2AY2D6b0rzpXsbC5i33z5jc1xtO1nVzQQzSS
jaWnX7CDAaywS5h2SfiFD4KiYDQ47/J0geyC0mohfnANDsd6+stVE0uclzY+ardp
y+WX2wc5CEuTMNzmigdHBGJJaspI+ihpZV3RJwUpQELl+yNve4bye5ujxJ5tAXOx
gnXlpl7pDVuUooji5OFjqHXaoB6sxKfKeUkd9myIMp9Rtc1DLSJu6vX6m1IwBBWR
KXF1ppOUoHVQRYz2DlM+hu/VtPip0EpSMeklaYG84tv0gn5ZAtIOnxE352o1uxBM
JLHj4+YcGpYT4bDD6IEV7zk/WoyjW5NWJ69Rpy2cgPKcH5w44YzxYv+eIZlTqsLZ
UheQ6OcUTlPEVOqMvPYnRhDyU/SbDGuKPv7RctyNqrcmNzo7sVAKY32x05EAgYAe
cUV6GS3yl1Yr7m5g0vGM4fZ4L4gCVR0DLzJn3upZjuSALRHFtfjY30iDVb54jfW4
CYbrHtS2bPZy9HMaIekTJwSL9dBydKDuCSJm1tDho1aMZPRADP6AVBnaixDrHj31
qtI1DIR5cyvQe7D2aujI0MT/5ZQ0pm6lyMjrR4MV4GBeVuwlFjeKL6NwtyZtmR77
2afsHE++a+YMWarU2z3Vk7n6KWvL+nq2I2qUVbw1JEkE+eLiKDEJ5644Xj/vBoUI
z/0HUGz/ox5srRIHr54ESLxXjswB7nLAUC2k0+HX9R5I8OnGx3kxq2py2akKtVXo
JU8q9WhxQ5/+u7cd63bpjuT9DgB6SuTw9qi64GAmOB7kTqdoYSEA8od3KV4pL00w
KTO3bIXaBnDRU3zh9ErLPBFF21ZWTof58ngccOZOj87nLaUwRVmNh5T9CT9Le7jy
KOL+V6x+pv8c+bEmdi6kgFbLiB3h3guw2W+fh209DCxSa8oqa5wVbNRzsqhXywZQ
KAHhmIRiquWIzR5EJHtIFkveD1+AdGasTbGywfW8NiYHF6/uJSd4Zh3DvDiZHS4f
LfNNgjGIUDn6X4UeV5TfejerIHXlMeNCIkJKm9kbDxkYcCoMWOpyHcsIXWz62fov
HBOvTRw6+xUdNsEbu3MJHwi+DXZjcJjSHw0rqIO28j8nV4RoC1FVMx4cfT3pqWYF
o/PjzQUsSZHcZVmfNgNO45mm9FfJneoIDFmy2De+bYxxqPYWNMQq4RYjb+Adqvdz
DsoG8IRuZcGK/gJN3eIaWCueidK81hXt6BYRgDCUf0g6vcyYvB207Uts6b9QYjgP
UOU76eoDvr2FPzw0qnFHXDjfF7Y/QaF5EDNV9G+0b+8FqNlDJi6yGg0kGt2gi1ii
+Yk+Ur+SeArThb4iSEazlwDYNce3FLoQUt8FiwagNchSvnannsFIpIQ/mrY5Si9k
Anrx+HUPBVmZJUtgbaYqPg+ELMwHqJbh38knG7MrnUdimuoNLHA/j1x9dRrPRGoq
nl65Pz+2frUA7Pxo+oF5O/DQojc+Z96zV09vVyY4fxQyIPuZ5HHSRJJYDXAazmW5
lpQXHsEp2SaIEe7QVtTDGLrvqIwe5ex3vaZ9cvvE47WrWEjfgLqHDrH+ba0HSRfr
AniST6+lJNMEw+xX6PCB9yXrcUwkEy4t0jqh3PyaLEu+gR8ipXSqwaCXEllJpatY
cZ0OmGRRzp0rctBzC9fpGh6otHduHhW8lCmX8/VaIozNF2GyVT2XbuLx8CF/sUeW
QYgqtnrGFfThK7PR/kzMFtrbNTzZcPuv5hOj/yIbe9vXzoJYGIr/r2wWzmkkpcFg
8kaAJu268hnkO49myTj5b223bFVKsA+CEYUigaadJuRzSYzWkC6/zfdUpMkTQ1m7
S38lCPc2rcXUI+dGksD5mzYxV1x0YabHybg5wNDEIQ2O+WDvRseuPhgYT0tmlzHy
0W9BMsfmvaqTu4EiP1WErWzxx+4uutZIif5qPY+4Xb4aP4qsAL+d4IcKwQftSfvf
J5sR/zgGttfDq1upmN0sTiGUyqPbhGD8UXUtKjbDPIIwkN6+ghkapjLs4+1qv8DZ
dkpEk2J9QG00Jpo8Kis9vsaPDfcBdiyGnit582KvDxSNRfOFDj5ZKa4RxHaBiCtj
UG6tM3T83jEq/RwKcATQrYZ065RftTvCYv3J1uzM/X029azTyaOOkNu8h9UI0Vtb
BzCOubJhLzImuv/7hlmUxSIOKkMyCUyXXLPKgl2M4sBkmZwoTP7tkiwsZhrwbI00
44d8mr6+WPKyHgUe2eLUD2gYecrTXGNOy/+TvgHVbUdj1s3LEvSYH1jdaC9xUv+d
L4WzDkqVYi2PftzvKhtNco8s44URACTSFQnjX4J1xBxsy5wTOuFt1MJMa9fd8h8A
PMwYFex4bzEwedVC+IJIjnO2RCUXpmlro1G48PJqmBKBHxGm252mg1jE7HuH3OXX
dUMA6cx1o2bKTmoFZIYNJklRSW+nm3IGzK6M+VmIwdDnRCULDWC5sCbl+l1sWsMh
KMgwambysVyehiJPB6RMbjdqNSKFWP80eXlvZwiUjLRlB+F5xTEUFw75lomR3ImL
8b6olOdTdBxBbXuneKcLCX1LjOtkC2ZGiIJwGd1+oBQGothei8Mi21lF7vcJsXTt
hTfTxJXhjKo5GX/DLoLklJ+5jpAn7KWSeoNDtfbjPyZxmj1sjtRukbdwW+YP7siW
kkUN+bde+l5LLqtD6/wjphOsBBkkhz2qwfyEjLsDe34/Pm7BD498PKTuJVXZM12K
/g3X3hIshgcatRZhCR74k3FIDKoiuGvnWqnGwNVNgKEp1OQHCQmn22Us1CqM+Bh1
LHb9NAPnwUXNyTiwUJjQmFiVBClQM/PvTW4iaC2joTQdyFz0iC53t2QiDLbHyln4
yM1khC2ZBu1hCPzKfAUhCktYJKIfe86VyMur5FJpE/NWDPtvG239acDSW4CK1SUo
/McWFemd0XOHjWgLvfqrQXxRQe/t4rM8WMtvtO/INHZ4n81QYowk1KW9risI/DsY
y92XzCvaGS0n6GwaBgfc6VaNxy4e3jWkMQ2VqWK8fTCevjVf8j4iLOxKRdYGfqm2
BW2UOKQJfngjKIFdHZiDRvHoFQSrt5nKOcgw3ZiHAFV4sJnj2hjxuctVkuYFOlD6
fztwK/mDsmT2yt3lfFRYMC70tGqt16CIXY4qt1J92ivl3G4wUGCQYaJTjnpI57AW
I0ZEMjhP0Rgxo8GiTRiM68XD1m54gPHmvNt/H0jq//MdBI+owEPnmr/NVqzde5Mr
Ybyx7lKbRjDY022dIqCreYlqajct758WJ+CE14u84ta47WgQoM8fKj52VtCCBiWj
IiUd4lMkuQ5faT/EvSc1lRzS4y+DhlHxJKVQiJdAMveqJzIIo0TlNWP4JC0NX1zf
rwhU05iWVeZJ7zb9kwQMz/d/GAR7kWjYtVQmCUwOfBK5SFBQN9shtfnmoQy2A2t/
wkzB5kFhlJfQgpNKTrTdKwvhwcRkfHGy9jYxvU/IYX0iYiEv3ekUvivkfczZv6vk
VdYZlJGVQGO7gEehE4lN1B0vtIRQ/D+6EDUaZrq4aEEv/QIKdeJKKQ1WyxoKXRkJ
NKebec4qREenAB+5+r1d/gKjkIFcc+vTL7adSEq6MCfimwkjdo+o+kNDH0uwOuvX
eeF6tj1H0AvVTOvCc5lpKLZi3UnhAJ5KVij6kMWaGBGilQQ2LleuE7EgRqeEF5Aa
ofJp/04oryTYyd5l+4DpXi0fKIVDD2dHrhIP3vEWEUF9idWFTZVl7zsDKlTftyYl
bJ8PZPcYgbbODX5CSnYDo/fFYfHAgYJHa8BCFVupVi16HbmXM3ai7rOZQ+BxLWUQ
HX1yBPH0Pd5uyhHMH+wQEWjf8lpHnQaekZ0bjLN6NRFi6WsG3vKcE96nItEsPGoU
zAE7l7DFCH0RuJPfw1NlatcQnrHQ5mFiovjfHhrSCVHGBjptN5+MK/GBeJm076xm
tYzOhT6G5Z6VPgCFw49hGYHxP86w0lurbFkTWQ8e0w1KWDpPYmfwXAoehVzZYtAb
awhH5g6R86a0WKfPdG2LDz8K9ENsdye61jL7DrJ46BWgXCEMFoXZFQ7H1boJ3WPr
qQjReUoQEwD50N7k5Lwikcmtvfgl4u/M+eXVNZc2/Ib7gkXqophae/OtwTu2AisR
x3V8XlODBH0X8IlFxD4EiP2QDKy0BNE9cj5r1rAuKZA2TdSlrEAJ6f5h3spw41zA
9BnCkWxhLBeJ0FbRNfTrSw9ubwqbSpiRjeXWjqUpl8YWeJuL6PAwD6LHsdOCBsEs
kzIRpjxxv8AthNDzDBEvHS+BhQayVzdLmPnBUa1k0LZzBrKjwFuWUl8wd6qwaYp/
fb4tMNxPrDTF62R/ZgM2yp9ztWxz26sMOn3z2Ld6SXRpU7445tW5/rYDkf07osGy
mvtj/atxh9M+ISBJXmIjl+7zE+zRp3lBUkVmEDcYV3G39F2CE19fxRdTGaziKOct
rGeuckqOmiwje+myBcw4I1EvqtgqCOszQoz+o/VZN3Dl9zg+wzH1xh/Wdb03Nu28
z4PTSfdwtyKiI5VEXFHB4fvcfR/dN2I2N40gxWggBSqolSzTsxaZz5X6iBpF/U0I
sVpyILrk6QfmTmYWU01KpUBQBrRZiyQ0jj402dayPjR2oSBD+tZNs85h5aTer0nI
+kpT+B7RJb6Vri/yTj/nBJZn158z5bzhC9jYVnBS4n1k2e+JF8FRWVvTsDrdEGTV
/iGI3VcuBYsLpq0mH/Gn5jZPxtDMdmhvcRozuR2RIHSuauZb1OhM6W+3UMK4rijJ
hh/8lLcsPA19E0Fy8pMrr7oP0HI48C8s+YfEI969mOFs8mtCsbczCy32teiWbPJO
mk2iJLW+WlUxn43r5Ou7sw5lbfShqnIvDyjUiirXeDUfit3aj9OYKDi++s/U+2Ef
FbO7khszOSJH8lFZIRFUwgg+QngGyytiid+Owe2NjK6r8cHjTnoamqigNH4ftfQp
bqogQ4RUcWxIsadxhWsqluj9/rh7m/pUjbxE9yajnIEle3tIRku0o58W+w2s0rKx
qx9Yr1uY4obQuHaQ2XQyQ1TzjUfv53Kw5JwleJVmwW6ZWyJcnpfniSNlzHKDcLs+
R8p6r13c09a2oD75YcpibW/xY4iq7nalxlkQn3bHiYFMcKVIAED9nXFnsrmPAz2c
Agg2AKQZQ/+6KQvXJRdelEzPkwEMfdd6PUYKjylVo0JfYaKAW8sejNvStKMblIfF
+e8FHh9sDveZqN1W2tqatSSWnkTm/hTxVkS/dwNxTyrSOek3Qt8wPD5WpmxLwL9U
46uMc4xJkL53WcX6U0a4rVI5Js6oLuZdmhBUbpJ8YUewi1dppI+avPNJoWItsAH2
mGY7vW35YEftXUj2gdq2Hhhg1Zg1wcjlnBQZFFXYjcFrHQhKszWaGqqVNGfLUhiB
ZvAde1h8GCq2hl2akGCVEE7JsQvxFdZFRcfy0KD/zk4a1rd+AJBvntaDQtLO1ZZ8
is2IhbAy3k8416lbAFwloxcfjlmuR4t4wVHj/XSHwGDBJziIn6ATMcT8Sr8r+fQE
HkDtpea7CIuRXEQnXZmF0X0HUI/FKjmBCbDsnMr+F0vK9fXTqzO9YygEoKLFCs3E
H8DSR6hISstRtgvN9qA0KWIqB8ZhWRplQ5bqmD/a+A39CN4Cf9qZfhH/520VNlzB
E8s6d7Ox5DP7IuHxG11AvQi/aD6qJZFhmwMJkchWPB5nJQ5d3tKlazP+79bZ4lfp
JWMWCAeEI55GXf5a3Zh/Bc+8c9cNs7/Mo+PX7Usudev5vDyz4wWQuMxNmEui19zJ
1PrxxtzeSgg8n7qmVVs71zoLOc5G6bsZdFR8MRLT4ttlUzQhE06X9G6cqScSmoKL
9vP3LU47JtP62URo+C6qeIYIZjMWLJw2OySJhCGjJY4kiQpCz7j9yRbMWvVXG3Uh
ziKa9HDA0osdE5LQX7mY3zK0qn9rKZlX3WZ5vh4sW6EtvdoKw7rfr5QgOPYlQJXp
6ldV0Zbh2bGjkWB/xp235BC/AJOCn+U2R4svcgE6RYvi0rrHbeWqrur7uZ+2T3nz
t8js2AWxZ/4n8c0McBfYcg+tQCAE4jX1WpaFSeBn5x5EH0eIraur5xMnqaVoJpJA
1n/kDRMq6VTXa180Mttjn3X4hq+5h3dt8TofXcNIIfRo6INWOnIA1p7Frxuwe/FW
3HyosbcGZjchYnrAG4pTBIbkxR3CEJy5Cv+DqwchcWxX74buEhgVvKPTou255UlH
ZLS9mhL9/05ATPawg0Q/KPuZ0bKz7l4Mkl8K6pBQH9L3gEeXkzueb3v8BQspkyon
bhifGdlOZHLZEI744xjV4lU3XR/r/j25cisQOIHziTmIIPoz3xNesU72wpoKf0Jr
0qcJ2uaaByczzRzc7sC/m05heyP9zAI3YG/62zERhuS3ybXWith0crxNyWy4q19r
F/BjFzJCOivNApkRv1JrXlQkyk9eLGLSJ65V3NyW0xf4/XXGCOnTGo3BLl3QCplM
yeTRA8LUdiCCphxAbThCt6QlVWCpCw8nwcmFfYr5jc56rjSbYL2bjMQjJrrTYyoS
nFLJqPfoHUe424bnT1OAYRvPVAJwjy5cx7Z1G5O8t2RT/eRQ2djTT5i/uGYJP89h
8A7nGi8DuufR4ZS4KJId1PZHX6gsywug8a3VdWobFXRUINHEHW1uTYYKcgyhxYcg
j26Cr75nebdGPmRYCJnanZnLEjBBpA37Lj9+qhlGV6g3ZpKZa7GgebELnY53DWqP
eiEoV3RWG3a/OZuX6C2wLnJCLzKJV8tSEO2e7YtfUaOvfAuO9afLUd/QNbh9D9yh
n8bpQCsiDbcWISsRC/qwfk39tv/F9eIwTjiStfVVhWuNDjBVYXIsYGKWQYRrlWfT
BvU03bDXVZ3kTUSZaqtEt5fYHw+V4qq/+9fsQMXnUTtnQ0231TfMWOwpoNiCS2pV
qWcAhgvoXhCdgNx3obPGeRc3qTV9mMDJQyVp8mrgDYJpq5Qg/Y4DZUYmcgBZ0zJq
tvaPtWUIYqPqhdLitn2i35uwbsG+rXY3tA5EaiWYIgWD6FpIb7ey9zrZYRPcs2V2
FXp3J7I8Esae0XveMLLOrsHGz0IGaiiIIKDBpdPRyIzp5KaaSBzQviipdffqqbmV
nCxA15LcNT2o3T0NiR08knky+WCaqInY/GNCJyLdc0Mbobxf1PMAY2Ofm3pSJQOB
o59Rxi5G1lr4yYYtgk+2VG1IwUYlzEXHyh4jkaQ5Ah4hUC22pAiasOlETMTOjXgK
arGmYh/O/w6wy7OclHCQIcEkrmSOanlsE7v+94q3EEIfTCP5Z/GmyNltNDOCq+qh
M8YDc75ii1ukZ4DAdd/M+IQqZZ0AiuINpgLb7o7vxZ2vO4rIDUZS8W4nHgEhK833
it0dArKlkxTxJBSKhmB+WQljJ+UkjqXiXPXMx20axMFDaPbt/tO94zzWsekOMU5X
hIzxamg5TodTqn5nMMJ/XaOkXVvprwOPZyZ6xNfuERVgqqueKdcK1JIo8SkTaUlY
Hv8GsnKibk28h7DPwy1FbEFUFFwhQWChhJT5hsDL2kXRXF17Bz1lEt8Ezyf6OybB
/YQvZeVm5MGZgbYGhed4oYzsqfniLvAnJNvSCIs3ipQXhrYEki5QoL5475I3JbIm
p6WuHMJrtc4VuxIa5VrrAZ0MzG7KBHm5iklW3fqGcYFxVXSH7n/wfFwI/aHLXw3D
OrmZ2B+iM4Kn2c57QHF4hNeafyyHngQ7tRQT9kSBOEzSxe1bYvmXGTQTm/RCWGDa
EiJTQ+mSf+Sbbk/0bEr9BYd2FQa9p4MXqTfeBcdFPlq5+vuMB7Qvw304Y59swlVX
6ZwFW/KHaNLkOS/PEldXlNskovoCQFYFDMkp1PoL06HPJ2HFncXUCBDEBLxGd4rU
vLDwssErs4AbXgtzpZ+XzWS63pYNtT/9y7DeAyng8Ul7cStj3JXTxHvL1pVoAMk6
zMvi/cOUJiqK0wGaRdeLzSuPzivzPpReqkR6ttCr0cDQkdLjfU25rT5vjATiS9uc
jqrANPxouolmzy+Usk2V/8j2E0fJ8wFLI0TY+kjXCSDPEa4d1S9TbTuihLyfGdpK
sah99AIWk37nnL/c1QAS6Rah18+qtTlqIacMjyBuWo3VZHHdYYHD0z5ZNBq4y1ej
zbR1LDD1tqAj0eZ/2BOLSSUwOe05Bn/yQqFHvXsffMOIodDz/dX5K3QHkDrhsn/T
QATJyZcbicsvRdhFSjfJYH+fh2gcjO8H1/ieuqL5is2haxe5gLX12XQpEj3KpOgl
vV5k7dgZ2wsSHmtvWHrbcpEot6KyD0YuyI2Hcj0Q1h/oK++uIt/Tq8leofRVOo2i
zTClCu8SPfgfutvllDBo8ExIOSwXfJKtP4FnqGSi7T+7leqUhF8S4y/0gt8Thssn
fll68JA80sctkm+snZ/JLAum1oYWVvDMZo9t/XvNk+3qEw6eO12+sYUjTsWABBvf
/yh+RY/UCvsX3vrnnzoF6+DLJnZ1P3TgI/gTRitRbTDwzYYV49fQpx4BwzuWICs5
UsdtFaW4zIIymJAhhY3qpmjnS/Gy4zxM296YCMMEYVRxNxHc5hqT0mDsum9E9jyR
N7JHJfHVY92mkJVZiPPyLDxyCbnVya/N2+7ZEFin+fM+cb1GJzJctgtrDMPtbvFX
sMFrCk9l5HpYhMmQl9ylfYYgey1sGNE0WB0ZF3LqasA2tYZdSy0KqF1sw3dXUGh7
ofont8uY+PY2XUrFvGZ6crIFKgBWEeLYgc0m4m6skRwL1WshfMqMKWEbfnWXvMUX
HqTN/QCOIJYFhq+6VShmffTAdbIlMUsJdhHhx0Iw3kVIfsY0SQAkXOuZaFG4B+9q
5mMro+sQqPpH31hOMRlIAm1obkYL/G7fqR3JXCacUUbQEBYQGVessHuVEclWJQ3l
fZPVWsqE9LFHjHUWLwHLKNrQV6zO7gLa1CKMOQt3Bp0LWW0UZpm3dTo0sCrxWnlH
UzYq2/w7TunIeFUMQWp6LuSni5EZiCmSCLX7cbxoAhkvfl3JM9m+kcrpXOJ0F8pf
oNSnzNehfAgbsLiarAu0NchvKaCH6i1hK6qUGSUJt2cK32zLeIUni3HuXOtdK2FK
Xyfj8hphuspF9E/TRcrWXyGXpvu+dJuEAIFBbdivY/XxBDs+EA1ishiNYtNDxIUn
8kjA9WW0UlznYkhZcwNiAHLnpAgK7PPdayrzBcpNyTXtAIRvsA/YA1gfmyspjuTW
6k856grX9VDLAzyOJ+jQoH8PQKWSZ/ggghIPNnV0Gci3Fd8LF6fxB9wDbwL3Kq/5
vI3H5m8TCLswj812W41mlAcg3y5d9hb1pKTUKolq1KmlzXJi8UPhgc6vahDSRUtq
qTuGbmxkA/r02Y1JSfhPmhhQj+6bJNjdYqHoDfXfWIL/xv97P+FjHS4+zKrpXf4w
d1CxWuMoXrViDria6fythRtWcSU7L51oYKKFkAoi2NTOO8phd7xnoU6NorWfT23L
mj4+QaUZQA3btrxqxXw77a0QSWm6aFH5D6qH7UIMndhCnxE1UPgUNTr8xNbPkmT2
eobrGTg06ChwOj5f55bx4aLSXq87U0PoaehhGhL9mhQJRSjCZusj1yjIYlr9V09F
kXfgxUoK/WdXI4K5w/6PqbKAeilB/9m+K1RIW4vE8ctWqRNjcC0CgoWnSqQublZP
GxEnKEM+A6pKIx0+jyaYRseBuuIQ5E55ef1KLwow8VpFGOyi8K2Pjz764pnTxfCu
DJh/kxSCdxXJN8Iq9Ku7sla1OSBUKr9NOjiLuVTCbbbLAX/Pa9XY19H+SfxgtJdO
AYFCZUBsrINCcgRm29PVrjU1IYbdqcC617BdrY4G2c4MB4WJKUVjUxx428txOvTk
QKKBR2Prf3mLBOSIOzDPRQHP/Nx3KTLpm/jpR0QKAkCsNdezySO2WP+W+EmDBzbC
Z+XZVZ3bSyHDY7+o74pEVyytxEQu+2o8h0A3RqKQBMTr6X0TWkzNLRwvYZ4CCZWN
mCKUkM0ZvZIGBZcALhS/K+h4sgaMOz1e8yEg93BEB53rLH134t1Kj2Ixtmxl91PN
ybNJku9ByQMj21/dp76mX2l9nJx9x+QSE7GtG9VaupwPfjbWFPVKQZbXXCQvNgKO
zkFtqag28B7gUxhTHAsDy1okUeu44dHtsRxOPbIgYoVs9JpM5XUsqbm9CVceatsm
02FjXcskERCRXSwkZKQCr8YLg93cmNenIjgXfDpzQxTJbtcN2GQS1HaUg14hsTQb
O/dDZgYkwmFgp8uhEHpThKWkM6yMvNMdvZi4L4LRVND0y39UIgnLjeQXFfzcelaA
GofuzJ13C9aNkzSdEGL3X5ADc56atMg77LoF7crKm8f+AoLNOZn8VDv4x45YqU1N
Z/jp2bHOIP8thKBh9iliWmPVLS0hHDozVUmHc2fxhGKQgBXjhFctY7z+lOQfGwNe
0R0TIKc1dYIPL0ONhGjYFThWz8CfxXPoTDtZ4DqjAZ4mLZfDjNQuZzyEWhrv5hzu
ZJyxcZLLA5Zi5qZ/3LGleCY51IieIsusuJi5U6HzwPJIoohvM5TMIvKBrnJDjCuR
r6C9AC2gS5RTqONFFhL+C87s1B88azecBaQfJvVb6FvrBfP082RymZcoQwEicWqK
n/GyMsEmLWEvHL0xQjS8BUElwYjPl7xDzjNhWKGzlei+wKefJMLnqbqX76QMl0wU
Yzb3b8tAI71hoQDOjr8nxxgQ+twpCWYwC/tjVYubXgPTDr62IXcv9tAwCcK9jzag
+TdLdZVct3E+FNn8rd/ksYVHAQxKuROSbe1/AhqI1+gYNBnVg5G3L3yq7K8IxO35
LRDAAnM5XJ56xivryLD9TiaDwUxiTEI1OrzVsEls8AmrctysQBwYu/tf/IVdNpwr
QUcEllYPhjYnrMHWikdL5jcg1PiYEMYtqdGn4PSI0ii54hWuAL8CHYoW6N/9X7Zc
Mqpa7+UVJyjgHLPnTGnFVY1YL6u2X2gBwkVugk/jhWcq+fdaK1vQJil0S06rV2j8
6bFSZfH7F/SERXgWOaW1tXfytd3q7FoK4LEbpUIJOKIGaEnZjq9ywAgn7Gi/M4tZ
cgts8KqCZELA2AMi1+vm9asT6yei31yLvJDZ45wplubuo5OQEofNyLCwyrqw6Ky6
0N7fBAHzJKSfpUU8/wqX7tAyflAsv8ceNyJN9xxMZBBphuO7Gh0TumdJEccUAn8f
1R0C5a5JlJpd8ZwjMngXdchNLoT5cYu1j0n9w5Uq7oHlg8diNI7cq2DJC/t7pO2U
iDIGyLR1axrDUfDldvfShxcLJV1CG6HnJB9vcbllCEw2wZI+G9qEduRbXJtqGATB
Kp1XGGRlzhYm5kyCF0zSW8B1JN3/ph5lqE53swgNta4rKdmsyKZ1E4Pa+O9Lh1vN
gXq2mkeeA7t4yCdc9pGwgJ0u2wF8Cs26IJtP+KQ3r1/H64w9LTjLWJissmeShKxk
L5Rf8jVLiqyw1g7Ol9T+81jJd2+roUWkrsPTo+3USui8o9Qca66/0mVLwBhIDDHt
ZpPEFJecri0jCaCu0gbZKggHX+QbzF7u2DQR8g1bJEbyuA4hx8/03roJ45tVdA9w
i/jwU0ppW0s3E2R9LLJS2rg2KLVHcxMEBSrZnShqmnngR2dkJwSVg3VLMmtuKI7+
mNJc57UO0cgxuTStue3c/NcOUcJbe/dGri8Of7vcjPMyDLQHEbSrfXiVeSqOwJIn
q7NkXpkmPj09U6kA24Yv/gCRQ2noMztcFkmq83wnq4M1Nn60HFPDvTvOvp1C5kfG
8wVwQ8dpb32AmyD/wKqRmq1Yfg+n7TCnwm2KSyWuvSMbc3XvnYGXFHwzBp8r2tvV
yWa8VgHpoQu29102eiVtQbH5steugJlWqPkR+R0AenI0py5lQgvVDxzR9kfnoiIH
8lqGaVovOBFubWa7pDa6ZV9myqgm+fqr4RZNBgQOkPYPgsoxThFRyafev5nJw/6B
HArAdC083Bgo0oBEvo5X91Idx3EUtLHlwtdwYQL9xU0l7RRoaiLzPeHqSIQdFF0M
G6AssWfZzxZYsG2/0TvW2HJwJc0j1vIaJqTxFyQfg/1WmEeVTa3f/jLrOYR43k+b
QoOYyGU1KOB8bih53pO+wv/3Qq2sNaXb2I8DEfUQIhUF+Dncq8FzLpV1mtcGwzhx
aL7Jo+LtfkbcDk1yN9yjr7AwE2rUM9gjQ4yMvjjiU9y31M8XGDM0HVAt6leX2xiK
xhdg3rpMoSxSRTCJBCli1zzz4klJ9XMecPHcZB/RdVRjBHVpM+EOV/uOtztI2cka
S0UPlw+DfeSCA8+L/xva0g6vlFZlUpbIU4S4MlFTC07GSdm5kE/YHrvh0kr0W5jf
LmKDkCGl6hZ/AJeKjfBHCkLQ1PQqmqLORHTeMXV7Ztb75N4baPT/ILe4+3YVMeF2
99/Ca3c3z8dGRsUxMogCuIscrUjmAHcObm7bmPZpfTr0sxC+C3Uqe0v4kdItzxL5
LbysBeu6V3c+xmEUaJgWPFz+r6fLyLISRYD0QB3tzh+mbVB3y+KQQvj31/d6k/X+
hPW2K1DCGM3FC9kwzq4+IAiGZSFND9IhdeW9CIpgir/ybX+S5MHHP6F4GgPv4b8s
2ZIV63HSTfA71PncSF1+wQOphLU5WtrW7ZMXIJvvXuecbP9AmxwcxNh3GJtuKSQG
j8IK7ESo0lQL+x+GMaJeNjjpm339K/YwNlQwXjZaFKtTFCbYj7WezZuGg1p4YIEt
dmh1nWbz+gt7OiMu9lr2GKd45Kk4RPwg5cSu020G0sBXz4j2w9CECuJOLyzu5KX3
Wzz/rmv0ZJk1vl8HV7HQGhekxDg2LmJEr3eZJocpBrry72ox8xz8XbJs9gBda+9M
XCcaHRPK1YHvbRCSAK8e/5gLpJutSMsZj0J6BoQw8y+O2EAB0xMqLGjj0F3DvpZs
hp7ti68QlW4uBQOeJiPJxFuVvO82XfW0DHRLIfxI3/j4sylBlI+ZzirT5u+QKlwg
MJ6lVXr26AOhYZyB26kbMRTrP7X7R+65tO4DzW1EvFe+5PvOkX4vC1n2tj7si3Oj
Si5Ivfa7iFx/ghJG0EqH/DWC6ONtJJmzTRhXFboBBdBX+z7Y+/OOVTLbOGlpFY0v
tpRA35zA7HA5rp0N/yu/8hn12IxCl36j3Zv0GsvesIh4QVLDw60V4O2pUtt9kIzL
SjXfaFom1kR6gR2XEYK1KxrLMqjkpE6qVLjpbQwqemow7MsgSjLZgiE/MnWtLFqL
+7wL6LjXjNmV2pQUg4cD0AfsSauw4XPKLmdLTxWEFRKMRTesWxrAJCYDHgKX4yb3
4FIln+K3jRRDmXiw0EhNJ+57spCX//3S2t1gjA7kjYlhAXs/hFr9txbL5G33WZWJ
WRK2bKaWsX3wuAmmS0aESXcN3IhpABZAIwS1uhk9uN5Ek0b9Ei2vc43vXF54BsLl
8TXY9PjILD3Oc/JWk7bcghr9QepxvjJAA9YnOo15PUxlR19VcMqVhLLLQpPuuO/D
8AjZIQrsRl9fgS+jC8kQsSI0vf2NC83hKrOVfZelFkk5rJRsyZKQGspxNU6UKUYM
3owoRt0yLN6jZEOHIkDSc5e4fRWyttt4NHGiT8henajWkwnEXoGrqQe9hRWfghPR
tEUAYza2pQvM9NxFsIGpv/Le6iUsO7NgYR7rBxqALQdl6Xx8pWvR62LFhCp8/uI/
UHDC1E819083mregh3LfV8USbO6TXC16AD0P9g8+hrEUG0Cpi2jIhkznJXq4dcGz
hfsOYZTjU97NMgJqTZ8aFdUj1RTVM7P3ib4XqlTJhk1lPzJgMmnpTqi1YZ5fW3CL
URB6Qpsp+4zEkU5SZcAyDh8nY2d1mtn/0ZzmbHpF8VKO6Kh7i9DhwmKHXqXgMdBv
bN7nL2h4b2noj0tRkXQUBkPgg74+Et5HtkVOUVvvuv7Muv7EHf5eNgKTvJtKWdbr
HDsUeOufhWfkxgYSdRi5ZOZ4eTlp/32Qbv5WqJd5ndVp2Et/nZZPobWCR9vBvW3F
+/CW2E+MssQgZI8rvkIVZnVxUtpGoGJfzgfES0B5Uf+nDNZDJaoekPTH8pkJ1+nO
LLv1gpt2763D+N49htSmGNMKTCINMNV21rY1H2vPNQ8vvkfww0BPQdRlC6ofcY1A
JPRAkrukEpv6QJ63yp+6uLvnr4A29Zlurpx6sUuzAxfOlAtudEwckSixB1+VKc2D
U1PS7a54jICIvSTr7cGJH0OUR3vKlZ1rOgOruWHKsof2gtlxiTfW5reW5du+gKd0
KC/d4NtLDdIe8XAjleXHnBJ352SLR7k0THKjIubPkrfS/Ieufd1F2wEWIYVQC4xE
IZy5dvQF8SHwuPK+asvE7AqvlWsJCsIQu1uaPZEAlqynHYs+U261wf/y1YWRLJ2P
YHpNi5IslCGaAWok3XezAtj/PYdKz+CA/Tdgb3c40aBSx27U1lfHSSaPRu83BwZo
92zZd+oBWIEZ5xfoFtAN5KAojEgZV5M+eTy3ft0qsVsvoTyn/WoeOhIfOIJ4Sd+/
GxvUxDCUyw/mZ5WtsMOzRa/avdY/KRoVSlWnU3KH0YR4+3RGUmgxQI9fksb/7oYt
PFdn0gw8a9nuhzGrKdV1IcRYA9pvsjcmfJT+TDCreZV2ZofJ7ZSAvfVF3+DscxlH
eXnmEPGmeCEvZClpqK/uDdqimw8fk6n8eW74lgfGAlGtDAS6N1XzYziXHeNJGb7K
koRFTiCSCDzK0LTML3JQHo8EgIYUiWd58u+zyZ3bazj8RQcHuDm6DWR8gBrTvKJb
mMDvLaUHuXAyWb/LJUg3MTKx0yJ+BKn+PdCg03lzOdEqiq2SmTK3+AvreI65VYm+
Jl+iPyd8ThV9xeoYI0ww+UoDn7GLgfVhg9VL22vA53zkx5VWOtvWRXKuQ22km29j
eVcXfRWLgf1N8wNvT6IWuQh0gIl6LLmZ4WVWFUdRyHJARCT6ojzDHz+e+SPhhOyz
KP0IIyNwUnBfo2StcI1rsepX/MbnETGiGUStgSkw6JGdbY5Frzgmdb/t1GiPMK3k
xYHYyk25f4UYHfAbomHYlQ/0/NZj30VQTTN6bpgdVqrbRTa37UxtbphOOSmoeQlN
1oTRSWzDm3jrK78bc8CmAP7kKIBno1QKGcN1hn7mNSaEKaDxw27JEk0/aiHG2NP5
KTqXH1v35gKpb6cciTPpqUYs2ZWcV5vspixe9hGhcHoseQmBCtY71aZaVz1rEhfP
wzy3ytieNWG+o0xbcRZ1UOfLT4LeYWQ9s+9XFRGjHIAFcOROq1+7VJKCA3LxuqN2
eieon3/ZvPfZhesDeqFjVnJlzlzzGOMKudGzT91Jf8fNslp1yalRAvQXkwtSlL70
IT96IN32zVnCM7mkgi/I82db1M/Jo/EGCFodJhdamxaTV5hRfJ0+NCjDqN78wkGX
VJ0WZGafsDVigARItmfMQSzsVSv15Cai3OAhpoJ8FcS40LpvdifdJ2OlIyABfdFK
NXOyO1FGH8i/n4xFEMc5bDa74stTCQqfdAdMBwJxLZfqqb2N8upJ22RS+Opd+dMY
QXE/igulM3d91xKsKBXT3+1nSdnr1liioBu2DZ7o2Q4Ave6jxRcaQbnkM6WpjJBH
Q6QPxXTiM2n+vyiKlHeR46jutoLWwjdRLmqKChnWdx4KY3m6VNE/nd2uT5afzDQi
kDj849U5jWSikpEBKZQJ947of7McRTMvOE6VV3X5g1qBAXyrx1rVBuT+WuH7RsJU
a81ge8uQCHVZZL9X9S3SMmP7ynT6terhxvOXrGhaO0bvA64GcNchORONzPe9mLOU
NpysPuG9G6gLTDLVi8DFaBFlmwZO25c1Ktt1d9zNsyW/UImicG0XUYtXN6JkKcVR
gATvaAQLE2XiEVJHL3pKjY88Ev0YhgC2CrNG29JxThtWpzIpOMi4oO98cL3hHdPa
1z8ai+tbW2PM0tDGXJ9kYK64cSBSAUmYpQm9qtQg6sJPi7RjJ/GBIgnQw1WxSg2G
O9gIhpJl6BAHWQM6R1lx7hkzWPVdjIuFyUITprra77CE/S5VgK0bmx21evHkEIVX
RFNmWiBAX6hudNLt0j5CXmkb+lAzAeXHe7RH+XeoKxxi6iKE2s/oSgEQv8oePjKH
eq5JIA9WSkVZcztoj4JXFXxVsw2CQgTicsXmOsUuYyfu5EBrFbIJR1V0zizaQlas
srser4V0S4LlcOPbi3zr/pXv2fWqmPX8lyMtPj5SutM3Bo3psVZKGOp81lqZod1R
BFoEF3/IHUFSeWbPWC16iPL5unS17kBGawWtcgKletrKbhCVBHKT+CsyeSLe25YY
5MMd+uEXBpvxz42qFfoHWf4qyeJ5OGoDUQe9xQucJWnZIlYzBn8CG5EshD6UZoFf
Xhv0Fp1bxBZHrQkUWb/Zszb5SNQGLTLZHQYpuUaxovJ9pijySFwGLFzwHioKgb+Z
LrC1SnlEuZaGkMN0KoHOM1+wGpyuGgPdXiBjbTX3S0ycHKVOs7cVLIn5LoK/Hfgc
1mDknZnv56mCXF/iDXFRws0fSl1zkC1xvI4lo9B6SSX1Ivg2vzUfmOtyKJyre0Xe
WrRfaA1ZFOIgMFsjnQHYMRdz7uvrvDT+uNMKKu+HqHZjt/YYQ4xI4N6RVaXrl2KG
hl2DNSOmRIrrgDvOH6JHal0F/FOPhO1udHn05liLODRCOPRK06DMIGvAbNvMJHEb
7CeiEyw34vOuTAfj9fX7dz6BM9luxZih3W/fCkcJbRgRlcET2Py6DDNqK99hbqIR
+BVYEMAgyvcRh/wdaJ8sHJU/gbmBhqutBRIKPvh+7H7TJd9TWlofpLcLWlMhvt3y
PVyBEtUVLdLQM5VRGUdGyiEcnv1ct6gnfzaMfMzT5uVwWh2EJL5zfvRgysVRAElV
3QR6OC4WWWyfMoh9msqToUm2gtZglM+a4IcWPl3mceVpDUtYg1N9ctMl44uJbPBs
W7TloWE1L+G/b7rBxHdCPc41YWLyYoXObcXGGUkKLFbs4qQEhF5gDhySTfz82c8i
zOV1s0q1TM3rCRNNYufScIO90AJiLz0O87t7ldIjbKGJz0UjNXnan+gm7rf/hsBV
ErKdn78XC/DSFwSXicaQX9krH/zkMpPtxO3Ep/GDjaoh91Qpj9mV1r8MsgaLqXKV
efviy2+1EZoDFGLXV0SZ8l2i1khxewTJ2HnH6QYbQJWJ2cg+j0xhqllLXuu23gj8
veEw7z6xa8bKrgXqI9ueiyoqNI9NS67ufFJltpPDwTy3XTZ9PORDdkf4rm2r1tDE
wNJEcFFDsyczlEsMuRctPan4zdrj2Fbc6itMlGCgrF0xXAwnydFdeOEx4pm/Ww0D
sv+1xK4duMCN/Lb+UpfX5hxwoE5vQa5ranCPvYaTzFpDz+2IvxIR1EpImPvqhH7J
TZF7bd201DMWpw+CJlIA6FxkgOnrFHQ1CxE8YelAMHTwVxreewmgz31MZS0trJVa
9KUOlUC4Tt5/z5fFx4IRNAwYWxd5JrUodc5eFFgGSJC/5/wVPSYnOQLIogdPEguo
Yyb3FHv34W7lH98YWN2Q1A0S996lg8CyFKZd3Ta9zM+Ycx2/Si9+xS7hHKf7PuO+
JiWLU7iI08iphh7/VBjK38s+jbeQaL2U4WaiBJ+il7m4HcNBc892cVdOpXIahraT
t+RN9tgBECCQ1I0KIQOp1ffZoCzFa3delGfsszmB0eQ95GGshIgdVxl341BS3A2m
IvWwCZW7qtMWr71FpRQLEfVnPnOWyU4EBloo3Bjdtd/cmYDSjcOV+EHbGS6E9Uqs
mv6Frp/CqfHYc1HCBAOLIwZsVEAgVuoqufSje7iRv6U+09HVB92Aa/PfG58PsSgO
hK/3tg1S8YH4ee+LjMLAkyGG4GocZ8mWLkxB1riNRBl4+LKFxjraqjRO9Osbm/We
q652CzweZsyOTIAiyro5+cXopv7rVNGj93El6paINsmSIzCY2wNmfe91FA27Ygpa
RdMd4yQ56/8yPH3clCTJxc9djnDur7gpAPKtH1wiwjAOL5xCG++m87AsalOHYE+A
A/Z9Q6P/KvvYh1uip3By8tA7qxlJcNfcbPhNAZxGGS+Ucp2nNnkJqk0y2EUGnRvL
v9IO5noldgrF0/vw4agWP+j8nTRZg4gB7cws6VopUxy/W9PACFtOWu/4a1VwX7mz
j+Z/fx+sLilvpiZzwYGvozx86ZCN5tBS52v262UievHvDE73b/yrFdNgHkyd1gyF
d55wbDXjiuMVlOT7OmqPOpG3JxCwAyGvleBUH8XkzJFRGtvgRVAxNw39N62pXonr
MpeJ1t4WCJjcGg5Ffum1jS6M6hflk1eG+FQ+Gr+50IFRirlkLMApX5PQRqpnKUwc
eIbIW9oXR2HkGiXG+yUJEYQGQxpanP14AZwXmrpSkJdCDfVQWHcVcTsOYMdvC4lF
Ia0ANkaMe571me1VbdNQA3j/ev7YjmRp3xQwGlgQ45n4ifIAqpJOZA+OOqtMQ6bJ
BLKwquShe+hw4/vqociozFCPKyH1XFW9Z8gj/oqsYJcdV6ONdH6h1RoMhpfCnE47
jh0IRz/8nZjC04gHWCq4AA+HLGCvq6zc+xI8l7HE5OFchdg8Z3guCQr03diEiPor
vCVqL/10fjirSsIC2PKguhMSL++//fd0W1r4eBiX+/gG491nV0Spg9xNNJp1bU5e
AJGRikHLCvzvWOxFJaibcjDnchrUiVmRoQCjFD+r3eU3SGwPO0BeYLKGW73Eo6VT
Z6tP7WVWs5DyDpLscvZ3/eviFMNK2/sZF1ex9c7oNKtbzLq9iiDddXBJ917umnew
7j/YeS3iM1mvoesoukBUjSxaZ+rAHUTkUeIxaLb/1U+5OtIiqvMLClb5gQyofcdg
GxTvB5vObz7CfYm7V5SN7zpHmQTFiWD0iqDYmVGum+a5J7INPe53KTLCX64pmQLm
uma46l3gPedpyeXEr3tGdHJj0W83zJpziWNQVqK7Bbd0Vird+cS7bj4ORX5RU/og
jdnNnLiwlT7jZj5Rvr3MdyLkBtYODGqR20d6UzeRKttVFGmy3HO5GQJtwQdOjKuH
H2W6yiL8Dl1I8a7d01rittVj4Lgbbtf9iWAu8j6KP7vWJxUiMvNSfJ2ou2v22AOT
2WKIgC9lJFtwHbg5GejkGF41eNcgQfxXjw21goZ5iNv2l1eIZC7F869gwnFcUNM8
m1vIWSlqP1V957cYwbkIhESVGz+DWlL/GIucJ425BmPjGRZZACKN/KjdnQPUeylb
1UPMPCqR9eLTwZAUoqwO386xwtal9t7LiC7vnZvlIGDJY5TDcVvOMpL7pDQaS/HI
PgZ0vksRDy7guiCiMyQW0eNRODTyFvUa7LHcu7QZt58Sbxss13F7NLYN795WFIpx
HG5WoXRzd6VnEAxBWsndlr85DsXp/jAHUGyYAYx1N7Whdf23Nb9JV0rwsNPxJyoi
9/LYJj6sSpwkbtiOFS6Y3NyYDRttzkAEai/xR9iwpstM2yha+Z80ct1Bcbsx6+Nx
xdjf7SwzL41W193EYQxIgGMzr8aUhCgnSxHgSC4tU8OEdZKNsRAewExnHP9G4Cwt
CR7tgmhTflp0G3EVzJaXKJF43FEHN6cI1/BQYcPf70b9B0YBhHNJpWrJ7UhRY/ha
PgE/r5RltLXsitrdfgF3Lg5WuGO1ETkBo+Cw44f0S4O9KYwlgJzgFQFXwXf4uDKV
xmLmjU/63QPy/lNG9Z7zJUgrnOQ6a9cafPXBZWSSPq/XAQ1i87QpLwA5hHFvxbmp
PixvvGaukniQpubflu3Q6vDiklyQPby/OWITfJBu4AvklXftoGj799lgPOCryA1e
erASvAqxrxJ6+v/6W9BILQ9j0liDk7eBOgWg5Dlu9U7zCd5Onqb9I1nG5yLwD3BW
NSt64ujhuisFYl6+7qegQTO/gT9W88adwlEjg3wXIuSyNK4P5bAE6ji+PBNo8NtT
hnAiIUGNWp5c82oP63gc13GPAkATa0HmBovWuQ7uAJbNeOnuI3U8ZvdJLp9g5Phv
+B2MpG1FrEYS6nJtsdl1DPoxFdAyEzb1M4ONID6OhJfqxDYnQrrEFmCSV8o0DJkp
TJOEA4GuHIBtj+lQVwKQhA/6PfHWIownfAj5TXRR44aoo9kmB0oJiSJLtkkvOED5
l3LYnQ4QkTlN/PK2QmxHmbsXU2dvv4zSdvKbXbvK1zLe4pl1okFDg8PO0e0r09QI
ZtbBc2DMt7ySyWjvQQTaEp+0utHnS3bsypCs3uFfh3crveyGyHraikBiYzntUpQj
a+gNGOU8aXVasMfFjnQnYjxA9RyEWAf5vlX8KPTpPrAoJog9NkeiMLIfI3YWJjTo
xfHPeYFSYSe0zPNFOnXWLUwrEWasP33zAmBpVLRmnw2glNKuIYaQ16V1THxOTNMe
zB1hlc3pqpx1Uz0IYD7v9lIVu1hmxf9Fk1z2JjdoPxxME4wRxx96nzd9U7fM+kRH
ttYud4R9931TDJgxeK2NGzM/ox65u/OqlyJK8jNSitxdPT7TIe327A7ofAj43H8V
Ty/pR7nflfoiRJ96jazKi5IlkPrVg8LT0r64er4Fyn4Q8FZJvR516Q2SwSFBh9/U
SIQkqRVNZ397OaMp3Gbq1S7kziUtfL8WUv4jWoteLPHfFNw4J3V4S6b5qQLG63hG
ETv+REMwJXPIB2OGF9a0ixvDR6wzm9RKHY3LllruMxOFSl+myqjY/ivAWyVJr8oN
TdR3qR0J9nfhoqB/wvnUeHom5r9rxBIhPfnI69deO/iGbBzth6gXOY/ceUVG1Qrg
L0ORkuZz/0nanY5//a+dy/rqyaiDlQJ8K3I1UP5t3Ms+hbnoQDzn2hKclX4ctChK
4one2evKx2lvqQKvuyRVGMMR2WzANlww40zyx8/buP/iDnvpo/uLl77L7PlJfmfg
72NnSND7/WWNejb0n0vddFUaP5kKU2nUHyv1teA3TzzHcuNpSlu5ZQ5hmrl49kDx
BSQbh8vFkwyY7jr/ADse0NUQLwdgNRMB5sOQdkG3TI97muzeG2wJ41u/9DVcXbYk
DLCRc5i2W0gSyzAscva4AyqhQ5czq8Vp6tq61XRIGYHPvTNzyb/ugTgjavkb9+ZK
3r06lWTv1tm7RQy0LjrGgXTAcgi/avHzs/XrosVOGAB0UPYT4SG7sgwi7lHJw2Uj
BEZGWhhvwDsSkNOyt3Slyn9NsiX6pRnx4zb75u2XS4vkLaKY//GuP6p8fQSiIuZH
4hz+mIwIJnBU9j9z1DwwDRWdrn30dhhU2JB31YRmQjskGDo+MbY5+bJ0Z9+VNCTK
CJLVtF8RCSki0cPFd1fQG5U144rxDBRTeL+JG9qVGRkTZIU7tj7H3NLEdmw0Npa6
6FbuaQZx/UbO57aPuzOczfPfrKxePluFgOxWvnts87UV15ZDc4tR3YUWqt4+wtfg
Q1NEQIMQcyRPbabLoX7eOPflRTQS2zK8JcXLrNJ/mDOKMdFpjnChoBNzohxwNwXo
CpFKRRHJnnAYxw+8Gj1i3ohATlYdAnsvQLFJUqb4xlDURCNx8EEC+knaynzqxFld
9XHhxI9wtTf+TpW3caEHBfk6Zht4cQzEwzSKWW52Gq3BvrrdC1MfOnrMjf/HIyCs
vHReuNT5CXeWND4vGeFhA9hALdcVgBWJM1gHOisZxUk5kv0iJf/FPB5W0EwRaO+4
pF+QU+/VXeSFMfzQehQKSMh09rBj4BYXAJsOng3dkURXGdnRwN7SLeF3RuyUvzTH
1VUV3oBEPgdDpMHV16dZBJN5+tmioE69KxovhxS/5L4fto9D36J+rKkcdZ3EYc2r
s8+gOeH3r1VyRbkOryTiuHbx9dgDnl73OV8DgG0rFDI29LXIVAuJHoJ80nHj2e6B
1qfoXRFJX9g0EV7+moWyRW6lFzckKTKdxAlK9mw/rMnXp9uFownAqJ+FZj+pvEA2
s0Bt0vo0uJDIpHmJBVtT+oDrZ8CxSM9dTwRWZ+KgULFLCcbXUXitn6nzka6rymnS
PbYt/hqmuPZAbRR+1URTYGfL4kFy3eMdg+hJper6IoYG5KwV0QkhvItt1GWMt8Nd
W6K5dT9O87QXp3/zwQNyCp1RDUQukBh3FlIMh1H6puqEg0kfEsoRag14GOHsqvBd
r7ITrRAlpTJYBi0e+hecghZu4q/aFguiPLA+qJSfAuk9ZNS0mbWL5C1yiF0JXYKv
iZcQ2VoOiZZhZ3suBxc9PaKZRr/m6vYcXltOu5qTW6/HeRA+1/Y//T1kjBvflOVT
KYBiPtCXGkObLbn2VaoGI9+Ov96gEVXzHIELz8U1wz6iizDAdD0n8mbvdH1XMdy5
GmYPK1Wx05BW4CCN4EOxU+wRY9hiJxo9PxhAVuBeN8XU38YXGo3JsF751LMjVCEi
Q1RMWfI4yLSErKW12hFvSexN5Yx6GvXJvsWZcwt6t3ZhYDTum1fFzADo5fTdCfFC
OPqdkxgy5t8WbN+JhoKTTB0qSsysLtkQWDFvt5L649Toc5AFrn+J1YIBsywlImYR
R6lT4BHR8m16bEpOkBqgmThlZV+RY7W5TOnf+TLkMQdg/VCwFwz0OB+ZkzW/01HP
P8VOHv4r/QLq8/QNNnt1UqpWfCi8TJlmMyGdgFQD6KKEWqP2JAZFWRoehycDCwVp
/hMAV17jDSKGAz9XnVSE6BjlF0PBMuI/U0GXVt5Qu6kdePNzvrYh2hECStBZExOO
ttx+kxQ0b7xWJdT+GU7BUZshW982LaQkgBOAD4BvJZC6pVsO829QeNnA+US//GNG
0OMQQXcVX83MNcON9xXBpJ5Mp69rA00+1fbFmDy8HOpQ8hfNBq1KGlrfoz/nuLqw
/5kQ3V23vjTmzRfykX/h09bNJeLrvwST1BTxGpR77CU1R3cUkXF1e7nbUvOTGnWf
/J/ScHeXAvWKKOlHF8QLjujfGxW/yHYXNEZeN8LSuEu7JXPPopAmRRprBwe0wSvi
1NB02JNG8ATI1uExDFr0nEW24tQKMKPxphfLjZ9Z66D2qJCbIeO6qnIrUFIXPKMH
0n8hn1bX5odHm1787MHJkZYV/Oe7cv8AhrvqoiDAZRlRQzXGN0qwbewBlVPCUph3
2DddF1hOJMDMdSiAm0RqksnW1kv91J/R7VfPFN69031J1JKNc60wxXo0ZgG5QThL
qp9ii2oW3rPx9oioKGJusSrlCBrKLw/CoHMszdoKqYEFqT9eLz+xFsyrQg3cI01J
tVh6DuzyniR6znu+4ZmyUplnPqfTdQ76TWN/10aLpucytjhl95YKSGVjOabKHCVv
31M9RVictObLT6i3yViB358/4vhVcoNKyFppPjvIt4zNdKIkcGZMX2A3JJmjmVo0
SLNOn6fNk/h9qT7qhxnxM9N6NlAzc/EhshAzukxBCjFtj4EwnA2QsPDiEEz7xOS8
9FwzN1dOJq21kmqw2Pw8v0xatKLzS7FVwmOZyz/FWIqbiB2ZU4Yd4EbHtSUcFOjq
TYSrnF9TVAIPokJfib7xNt3uiCjmlgWnKOocq3VKDjGiBdDYir3A0ANwdH0+44bg
WDRUhc6RIqcstzNDqH1zpVfZrGbkfE8hoVODVzhnJrrs41sjcPFITNWXO2c7Z0rv
qkPXsecnjjUKMcISV8KQ4oMqIFNNBz0834uM2jnKCa9GvNNFWJYciIHSi/qb36kj
HmzbreXXEfWu6vbjpprGb2jUL6w3yI+zPPEsC7l+hk6QR2gPNgLu+rK5vNvWsJAX
b82PXYDDEqAbWdK+9XmyrmNOtMpPa1KeUTB6b21wT7z4K4YSroHNmTi83zk70/qO
BkH0lsHBOGbBwyIrTOnOdaM9KQo/KKXJY1q5NSdou+k0t610cFzrB5l20Z26hPOY
4PnwNwa2ERKLq0le52Zv2IXLYgnYLowZ3sWd9Vmc6P9j8UrHjHQHZaXBsszYtSDX
UJDGR3yQauuFiAGzMt1XyiwbMKuuFhlOL6DUpgTSpaOp6W+FQCFccQ7ezzhHAc1R
reR3xFWW9sRsW720urbhtFAM2+VIpaFzgdGU3tTT46+IjIcc0lu2TYeiCMlPWZ8a
LtCKbxF1aILVKnp9PIb6TT0zJo1bkTfKmRhfS0/2nOj+vBwU/K/gP2hubQprhQ19
YcKIwx6wuPhOCRz123x92D9oGauUnxsCepkqWxe0USQpQzFsSXjFRQvpF36x/4cq
e6LAXofUM7xsc68+lqNlpCVwR6o355XdgVSNRwcZ9yx5qYk8Q/GpU2e5GlLojpIe
JxNlPvGlwfI6gkm50rUXG9DcR6YPX+rO77DrFAp/e6XnX2MLoqNITN20borhl3dO
qvIe39H725PKfsVVx2EjdgFq4g+a33tfwQpvUjaacIL0Upb9t7ZTINQMZwtlhdxw
zYgWmAa5kdnWz0xpjt3QXZVINY0/Q2eKMDi5yCTr6287NxSsVNkHl7aZF9844Q/y
n8SejkJ4WGbdGNkXg4HhVf72CIrBWG+C6wNvh7WHP2SfZ3mv9vjkp8mJIuSzxgLP
jeBu3NoGAGEiei8mWo1NtLg11TogdJLY9u3WhE1x4x2uzZLlKVhuEvlHTqvOD3h1
JHCaoOtsaCNeGMEWXqQk4RRQrx3CsxA6kSSgm5x39I9VVqs5cC9nBt+ucl2tEfgg
M6kajf44Xz/7zMd92C8YuvR9gTUDTPrERDbWVUj/j4g947DuRT+AhbbbiTwGSWup
QQ36E16Q+ws/2oCZHHy0hgIKHjHiwcpGxro2yF6cO3BR1E1oggwPsLDcdIWbqfE8
3Tblv0Cf83NGD5mEOm/5lAf4AbyM/5Df7DbEnC+7gE7p1vhnzyr/GW8N/6lDRNne
iRtwTjw6ssOsRXhSoiMqM561Y7UHg1Xqu6Zawj7E1WyNVMwGUhy0wiQajZ1vQdQq
wE95a7M/cpkCXpBa8rZCbGPAgbA8+MW2VA1FLUntUDsKqY3Haur5nHvnWAqU5d8A
OBXxGpyr4eRfBXdhHUzMgnROg7NHCYwEcgm2/lp5D2mtkSz80heOIk59yzP8QhYM
A4s/CckaRkzLytfDoES66IesWvkunO2wIPlVnkg5Z5n7l6ne8C/81lIMfiZAWAkf
/LCtdoKjltW7lLAFX06CA6BXAlq9hqDsvjHuW60F3vzcca2V0byJEY3Ydl/nfdWk
XVkIukkXR5sULQBmTeIwQ5DbI7JcP5UgS3NNU+av7dcOZLV3WWzH3ZWdVHRlaW5V
oC5FLGnqYBldJF2W3bqRGKyKZkrLAURZP2g0P4MG+8RPNDLXb1vk47wO8GAbhI4h
93yc9zb5W+Oi0F3smpRERkPWGTnjKPfZDvEOcFF31Yl70nMFJLuoGp/3INaE+y89
eNpgr3QIEI5hb8G6Jh/PYlEMFvsJrScqK4rr/WoS0IeYDC72N7ndVKDwjCaKyK5y
PVFtLrkrPqv2rO5IefwnRdhnVQVhXiQvXrR8V6zYJA1GKDUMW2wjpVyfO5EnSOOX
T99D0XzzoLXG8NUkB3L4uRHG9e9bA7LT5tLcTr1UGvwWUqEOpIZbRHyAc130q2cv
2kA2W+a3T8YbT2vHZ32/Vgez4DkHgjGgln1Wt/zfJrNUjRnbCpcBttSG3Uk7FhOL
VuMQ4R5sIp4TZ03/rv9wMtODOcgsJyANCrXkRUCcMCPM6ICngVcLqFx/6w5MmL8o
5DWEsdQKiIbNgkX7RotbwZ7gDD+h0Q0EqHWg8XyfaETTXd26iOgI72ZjVfP6EvWq
ipUMoEXvCS2JESC5cmxZVLbm7bUcSAnQZavQ9zE8JD2h1wtpTeb5nrhrMeFJ1aGe
/xoTbAUCj5BRro0ibojQyXnlL1D+xmVwlrlvVnTp23Z5IO03Uw7fdQUon5I3r5wM
3fnaFpFibPVGLxCee8fR5TYudLWrUgif6VceHDSm1Ih6Q/dle1TAVHd0z7MoRUMp
Cxl8zPBDtExHRVERinKveRvO09AfhmCjSe1nP+Q4Fguo+apt8YEsY62AphKK5yq2
WepNSMhQ9l2B+ewNxQ8AXzGQVL2u00JsmRCKNTf/SAHzvUfvZi9tbVA1lXfXXagt
jNrjcrRVSFqT7r5L0AFcfjv+aUl0T+MHaIKIC8AGB4pCzi0yKvPUMrCRkURz1RwO
XVxW5S/yPlPxOIgv7s4kI5ovVIhgGoQ4qGr/5fJMBzn6OHDsvOWYXdkW7+FyFc6Y
hinDzmPJNmQyZbvhPMefo9eTvIUI/7i3Sn+I1pTSDDMwu6n4DVJPd288yFaVWdD9
BPYRi8Y9S3EEEiO9lBxUNZziugi5HAaK2Fu53cF3QCE+VSXDAy6J5MdfodOBBH02
MFNPWUiQHtz6nwiQOv6zWNKRv+r2EAR7hsmWK+6BBNKyMI/jJIYSmdRwEMXM/en0
4DlOqKL2OBdyvkwFQJme54ad30O/ubb4RRZBndV6hoPiQ5/+NBtqQyrBvpe3E1eX
R+6Kzcfl5NUMG+1zs4fomAb6qpjWg75Xl6cwCVazfZ6CG7fo5GxDOMbS4Lzt9Kvr
Lxiz2NCymowEOHjMpFTxx/nRuPYBt9YqlrAFnVJgce/iNh6dMdTlMfyLUrYlLz4k
TmZxjtYuRlJFFytWOVKPQgOejLxwgJwidC9CxhRmH04NRANtQihdT0yTUVEcQgGp
Gz0ZMsk9WtymL8e3pMjcPO108gJL6pfkfCZAZRA5mYQi7LviOYSyS/5T6KeLT2NC
jCACw/nkTqOEN4GXf8ADIxUNZqvcj0M/aZ+WVW3hs+Obr7bpimdX856Rjt95OeRt
HToB2cV8a3XF0VdOKTlazcwIzeWpYMa996ckP5Dj9eY0SeDYYqQTrdsSraPYByIp
ENWUUm+NCMt0T+DO73Ya7fugKhugwxNKpOuoqwUeU0LL/UKKBq3G+Zl37pGpOa5a
Nw4kKvIo+6JjlYjUIsP2g8m5dRtdeNj1IKJrDF/8mVbVpgTC0mhihbprEgxrxPXJ
tjUq0mJK9ErxkEYSxLYyM5jfmTa9nApSPtD4BJDbvbOIY4LNRY4BwDF+6oQpo89S
F2wGj21VdEUD4gm04R3V6UMt/k3K+ALNCIlK/Ekst6MgUj5Qnn990oXpv+OHLEQU
XaM7qTPDGQHQdxlLBszO9B7VQicaHzC7bWx+SThWThBtzFYrbwRhhZgLpeTULsMR
dROazBpVHkvRk9uHul5KufLn04c38fT/Nfae20TJSiuMZicoTNvUcq0OsyjzCEVx
BPHBot/Pmh+lZFObJKemOVHbT0Y4iJxEoiU+5n2laJvLMFCgMGaOvNCujl6mydfK
wIgcrhjK+JEi78D6YSFAwnafVi78vmBVB8HbLnMVXbb3P70VT4F+C40iSqUcRF9X
xLBQort8l9hstxEdFm+2h0BtCz9nhVCtE1tO2z8JFQ2Ghx+CfuXver+13+u/5Q0X
p9HG9gq2P8zpdnvNDWy93jzC+De/Zhy06Q+IEWyYoQ/ZPdj7pQOyYMs88obQp1bq
HExtt+S8npQaNDIF97FVUwMqkRRMairKJ3FKb7kTyt7qT89SN9Mgx45nrxIyjM2u
Jy1QXMmIIBRioSa0wXlEsTerCTNVJgjlJ47ZoEt6B04W4ESNqEVf2TB9otvDNiOo
FET2DR3v5LShxcDJwdKZPLZyQ84kpA4X4B43xmcCcFyrXCcahKqnJhMug2bR92pe
5orh1EHlyl7qNMuKitimJsjTti1nMeFsTZ3uY7uQXAsDQuxofW/R9SBL7B0KhJ7Z
ZJh/9Fl2poZVQJf3QjWJKG2Xf+t8yZFSHTSJsysiJl2AMpqerqbkJtmGejqxbwSC
0kiLtB49XHLG38hGItLZIVfY99hCtveMJuB47QTdoiOXHW1D4ARIS/8kKn2TLpUQ
YW61inHzH1gl1lCf5YS1dL9i5V3egfbP4pmykxPwEV9QktYtcrRqTD7VwckheJXG
cGTwPDfUtUoATybXALYJaUR8YWUZO0L1zgAw804Z5JNOXmcK1GGlBpepm1vDBa2a
2bBUSq1/N+WP92Gcm2ffoSWaDqETRHcbHtOQ47i9qmnjmo4AZL4E4SEkpSIrnGs1
BvyczGYCLEdSZgmcl6/QE7fOmORoc4rEiooc3Jl+zUro9FoUiG59vO/xWCBFZVkS
v/2K3/yv0ZL5/RBxswnPmEtd/XXsipLuAEPZ/RqcKiQxpzM5JOiurwg5rb0lev9h
5ERIXja13m0N+gqfgz7p1jw/D0CHbZ8dDfqW99Mx/KBnUtJyZSRDgBN/eQ0Dxhx+
BWOXCwpLikGg63ev5JaQPhF5t0e0jdc7V9OPiNwG81vBolUqwfYFrOUTVwUf5cKu
1KyGzD48ePPqIebwHJXUo0laMAxrdCP3GZOUNa4ORKX7h4F5VrbVuRwkKtkEJ1F9
U9yeEvvRWHSaDm64M9SrGm8s6t9wWzMIux3ZkF8BzhkjSjv8fCzyZj/vRbgLM1zS
C4XC0cGiP8vYn3iJmxvyf82JiE9fnrjAfNNbaUCZjJtQdHHT6jVofU7vL0lWm3jB
R1JEiVZsYqXrN3Ho7o/0Dmqvr5/DoJBFR+otVxg0dw7kqKHUSds+j1sCtzy+pnNx
35fQfzTWjpQcw3Kz2P9Is0qQAWVkoqJ/xo1ZOQYFOFv9eRG1JWlbheLzR2XZGVad
M8rPfEeH8on2ia7QF5naQ/45GkUd4MWUAj8iEYGnP+b3ksihc3CbzlBRQ0j7rjp4
ziOi0wW3JTyhbJzFac7vpK1X7YMj3Bt+8KxlocuyQFSoEOOGQwoF6yQum0qICOgD
MTv5pOmAvuZnMjrM+6PFB5r/lt/Q3PcY7/V2jWmRU3pekI23EPRGXygL5p5NDNP6
F0UnU+1pOXUBVEbF/9aSJ4kDHS6f2c4JzNA36o6W059JS67f6xPLHTTZ9fZOSTh5
l3s+48DlH9Bh3HTaDlwGEmbBzMOt9uL6PFNMcyY3QgnYjCym4KSvEqYjxMjcZr4z
WS78HvtFPp75W+0I8vLoCyojfRIb2xhIhgMP0fsWqWW1sNLXIfSR4rwsXB2YovH4
4pZ6Wkk0eC7JDi7pbYNCQSwnSCsrjpcSEwBXenKnak6k9Ip0Tsu1aPLr+T6R5B0g
deKq3KRykE5X5DUGgQngGgq1SifM527BoOdVquMIe18OGCQemylEQIM7Ig93chHt
fiPgy2SPTD1QeOVpH1cGDn0w+/TEZthxs08iwbeejEMNB4ltgbwAj/zCqgDgb2nA
QNvWcrD+su8zkISomYqiFgeSMnEbSa7n+k0Xcpa/ZKNpz6PAHWxo+M4drzEc9fFV
bNpo4Omj8GkRgwKEBvMlPsrRiVNPiyEPEZ5kqhm0F2oot06aOTMZe/FoXRPb/LqS
KGIBrF91dZpPZFURL0wtYsNiiRHAF3IhYZtR8Znr1uphtm89z3E1iA0Upvi3KXe4
qc70WPmDPQ3fKIP/yKzFC45jhqACTa8iCQb54eidKxwUe0wmkXyP+jQ2eZLiv2/d
gUKvAyiLWamHzp46EZddP7O/0N6AaeIeBY1jTnnnqA7fOyNZruJxCAJzUNgA6SHE
3RUGKCcrv3mdmAgvnpr9Buvw2tQvAXqugZjSeI7bIlBdqvsfkg8UwPtOwJB3QQS2
YspUccPfQ2h8PfhX+6GA1y48W7eeXV9rpCsM/ZBMlf8XemFwbj+Q1FDO2hcHuJL3
5K+PQeUz0uraSWYKxMdpceHi3qK3oopIdYKD2l8gqK0EB6O1RNURS/UD/j1ZjDBY
+Vw7nQapIvUBqI/rxBzFYd/Iz8G3Lh6RN1uCyxL3pk1+L6k35pRBDSwLcfkMt/DO
uBTfruxKjpGQrybG4SQI/BRJdJDOP2u4YTZNxOCorFxwaM/oN4GuBawwZ8D69EDA
FpPN+EjAxcoDldr1N/ade8dKEcQsVXdR2Fm55LYiXp670xzCtYv27OQpMXNiDFlw
kWznAmDgyXM8hIQS+1O20rgfRPG5ZS47n7jmlGfI0pXfQEKR+LSiYJs2adfEOGWC
0XvHpNzOBC6iNzJRZOyjtje9jYvZV1eIYTiVAqwcBqwWkxqQgx9CT01RkgCeem8E
9kGP5EwHV/TGCQcJgFyKKVc1PM3AcN2zmLwyVR8vhyopJT3+C0vMHB8zfMgbdmeW
Y6VTJm9yxwXi5InqIU5QnAxESp/HXjXjrzbs6qpi9tT6cvw6NHZwMHxZe4ZcD3oB
g/NaR1wxi2CyE3hmhAEpihEZlcGh5JdXYCPaQ/cwpf2Knd77VZWVfPf/uaQhpjce
x/qCXIw0pRKSTi6X+JSGZf3ehGqvDwy7NzuAEZUXquSpf3TsExL5UcJdqhGTjroZ
pkHFh8BQJ54E5IhdtUy3RaljpLX9sRYu6aDBijqi6/XvGjLUsF7LR1L0GwAJQam8
1kPJ31+JK3HxqqTU6AhHc1BYCK6GHZcZuhO/xXbhIiX6bIYon/Y6O6IXKgt/p54I
Ug5Ob2Tg1lym3jch1q4x1AtvaXpd7nwbFLDh6HRROS8TnJAsnXorAFgm8YpQLc5u
8mBPjC/HMobMb75ZshRNHPoE7i8N9jzeXPNcWzKuzIYVlRwlcd+K+vfN5jww8cNs
023EMxqj4t+Pu4ZFhBOiJ9VezNbJ5z59M5mdnJk4dUYt166hULJHjhzyPPOvgidD
x2w65dVbqGsuDbWKuqZuIrlzzZuPqQALJgn1oV4xdWJV/3t24+xfoyKY79z1MYcL
etHlPpAw8uZ3PNZog7stO55nUKSUlpdWMY7pCaGQufxd1JLbeKUkg6g1LpSVZ+8L
LB2Wej6MtNwuaQd6y3ByR4Cke6QOoa2X62R72wdrXdx09Lm8+WmZJhNmQTlYDx9p
csbUwQ0hMPmO79dQPY20oA5t/8KcMI/cpS5tEvOL/22wX4JtWwnhg+pK/myQ4oLY
oo64PjCTt1ccev+vjah3EwlRF78pAGXSDjWyNKovueEf0NR9GQg2jEd0m+3pI86w
Jxuqjc7oSSwLBRnJ6x22WV0QHjLsYzT27KkglRtyGDTTZ2JN83xPxFf3InKCXDbN
HJ+jzWXuRu5q51xrIVRF3l1Idua+erMluHhweskic7cLXACAhpD+qEiSbYpB1j85
Bats41oSTkaXKTgnzLjM1F4bHOTL8ViQLH1r00OZpQRaEpAJ5gn8UZCyMXcntquN
LbVNF7Xf0RaSfYBOt/JLb+LMToeIDmr7CZ6h4M/wluKTw8k7OcWSB5ZT2xIv9hq1
y7NjwI8lUoWtDdW1DVZKVqezB7Zzu5s1qWG7IqLdUIFQDncMj7J43HgFBHCopuWh
mxBuDVmxAugAnHA4hNDxCJkc+uSxaRvHjj34VlxvNrLoiPb4DBvrC7U4CtRBXjNn
XwlzfbTPyZaJF0+6OtbktGWx7+xjeUfEArwrw8CdEvb07Qy6BAfZGu+PJybfY/aj
gjTlGGmgGL1j3i/25hyY0uEybz7RvLbt9/82uXWUOujxi2F7Y0Q3lfD0ySoUloKk
H78WfdFZYiCorH1CvydoemoTw8e9vVNb/QQ1czyHKfqizSgIgAD5C9KZ3AlU70EY
N0d34rxDdULzCLNthJ1KKNhV3lptZrxjhIWDCEGaOaXAradk2HNhCf3qkPdnRoT8
JehI8dNcB9NfYqvN95RZ81Y7rgf4xFciZT9BJJZ+HL4+jH5c2V6m0QMAYI/W4t8T
uLnyBlGOi7GHJ3mnYvl5FsIXrvKKoWm0pGkwqzsVvW5jEIYJwhySeymlq8SkqUBn
BMJuc2ISwI/V3RJV4nS9xr3lp5wDVtZZmXsaEeWKqcGMzgDlzAXDakMzqPeSdKWW
WXZ4GPTgUceWXXlzUC5z7zEJFCDKjtqoyCSlAJyZBy7BSGbR2EXYMbXihLDtqZK0
0PNjpz71lZneQvCfwAH/6LOqU8de9u++AB8Dzy5gZxHtRJRtyS6HcIgpGBKWkaFn
GgtudiGZ9lM9k04zKKmGH7EpoAHaKABGbkLL/Y84RhByJ+kessu0aPIkrN5kQZUV
lZrMozaTNi/JuuRZxknAl00JtTeQ7FYZgWSLUZpgWpF9uwCy0tKph+Ad4nmsPQgR
mm4Ac3YQcpmWoPTPb/XalnTE6AJudTACo5va+ZQ7q8XnLwHfOleoYfV9HtpFb+Ex
ps0IXC3S1CvCKk8w0Zg5WLrXk6yd98z5/nkgg3OFxOQqfy/+gxfmiohYmsk/hWHh
qMpf+i4veYfiUOp+Sm2ZAwtbURnv45Fw0pwEMA3O0yzKPXqlJHnA83U7TIlkLYuV
yZ5TYyVGAASIRJPZmbfVsELYW4gEzXLAKXX5GL2lG8OYHkEFVa3lSUWVFQHnSp2+
F9CY1RUA9NDQzu9efZQPdGFWP6wMMzG3zEMhGFRkiMLUxDZlDndi1SmgITKC6Q03
o6M35h4QpC30R8zyFzhyB3TnYQ99/1ABMhIIYLEdNg6nfwX0vR38nlz9tEFgHXbj
/saRG73cTPNg+O98mFGP+prJ7JvjSAUQ2dJ75Ps8UljhuYQD7iSY/NDlHVBHREVs
YxsXP+oNZmrzDg+83By1dxvKAEF+NL/pSgiF1ncbswIWIA9n4mCw48AnFgtzlQ9Y
svIXVXUrUahKNcLKAy/EnXHxzHBY1Atn2X3uKZd+/TOZuHv6iVSG1T0Vy1YEeibf
24Np+8BNUcbIjScyUeEH0+DZpBrYSXTHFncOEfQ9gRDrBOvq/hq/j6yTdYO5YaJr
/PB0w/gUSQmry6iAupA5waKMrQd07yiDzjtcN1RymUDinrwFs8NCjx2UVROoI5Ym
Ud5MyOvzMNG2KUJ3oVHDXfkFQ6Cb0xg08XoqGCpOaERecFbUMEFh0DQMZVctGlN3
NWROop3PI6XjxpIEoSw89KAnaSlBYwADDIHie8kZG9EPb/bRfLRaw05RZkGBBetZ
zLxVl6y59+tGa3dR/iY5zn8fKMCQJoufnG7wfu2iKNEvKrnIMwbvwpz+LsMoYnio
4FFeF/LM6gbORo6dVm+gwd0UjiZNLlfPYm3/KNTGNHogKaMvacLJgYvEgefWh8qf
3HM6ijEDtt7MskomgTIgB5LXrZTAOSAqYttn0JglTD3azCRUfR3JQOj6w8WBymf4
fCFRoDnxjm3MVnM+q3VVN3VRh/Fa9JGCXUcma6QtrZ+RCyWFVkLPL0wrXS4mSyIt
yjvJhvuldp9ZJNEh4MX4mHAE1w4XN+d05sTMsFzZq4rOJ+gFEhc0dCyjCMqdcngY
LeRkiZPdrz6irXbh4XTQIk0p5p01aPThhCi9vAv41qlpFzVUxA7PIxYy4MZAPvI7
07z0j0WOYyXMM1WE9Vx0fiIk1r/t6eH9zMsFQ0rGi0S3ehnKryW2/dfo91IHI4NS
LvNnNiZ2oMPpMYYxrDSC0uCXjsXbgI46CNIoXa6Ov1s6NYHFZgQbVAhsgl2m1QbX
DoUCv5p/eMQQzlDoVGnJrP1v12glA8kUm25E9c7oQYtBVIzo+VMR62PToAveRfBZ
G3KdLSuMa72Q0lQSLXqUNkGdeLdin3Whb2s+wkIYcKkzaI/X8diMUJpiJcYmODol
YvixsBd6LrAekfLO3q44F5STymlqYG4BQiYT3/OjU7UukRFCdQXpNVOgIrD8SVhc
phRHlBO3QHRNzZL7bI/v7XcqMJ8GbTfR5xsJPpyitoPkzB9zRQL3JEADJgXEutlh
KVNPCiR46PgD+Ix0Bye1l5UJRdOFevHhpbR+M70bH7AXibcWo4quc/XJExjqWQEh
3vwLjr2pJKCwK84e060HcfYMC05p0TslybaI/izJYj64zwyVi87dNix9wZ5yrg3M
6DawKef+/p5Te0RgDeAF0bzW4QNrhLuqLY67FbmBfCGgtd36+wpvmKuauUSKw2mW
CFTXwliFt0FfkyyGPE0x3tJ7fLxyJwbBjpRIZZM07rQRA8b6LkwpKhd8vc3mgXCV
ztB54z40S2V3AWuP/AnrQdf2uZoTbLv3KHIDhsxidTfMlpsvhTuva2yOMTpmXj4S
4LG+Q392VcryJPougB5O6WWdo1SGK+7j8W6BDh+52RUKXpGurhVhSPmVUV7z8ssR
s/TKVXoynM40IkhWQzphOWRHpmzBB0KofuORDXX0UtFFwM5U3AuWPbKu5yyxY82K
ZzycAvSSJ0HAQOwIoHWRci16lA6YFkx5DPaXp/JiJcQfJDvziqRsHkCsLylxkrGc
SkusBnhsipJwfVZbi2vYCUQnTqt9XxgzEi/ynLwW7fdJ6eOPnQqvimPYY6RJ7G6s
lKAHwlFRfpD2KJ5CbKOGJH+6zvv3qQabBFYu2JmjcbCIcMEJh2xHHrhWz+8OlaGe
MGHrLdpBKBtulWwqiplwetT0PEd4L7Nx2ufpWocHgC8/r+F3agTeuLxotNiNIu0f
p2TJLU+opl3EP7sQW3K8ryi2omYMetajulftSyAfKscTW1ohqXCU3EEZJTWekM7O
riUj5AM023jZBOS27UPI/oQaC2jLr1J41U6dHEJzfgOhnNR92dOov5APb2wwm/h/
c3UtnBNd76StVzhxaYJEHQ9pKCmuFoIYeaAmwd4v+ptwxvJpjYd6jX6hCqvq431F
tjxnBCuGePVziNvP/QcfNtkkSsjd+jflo81c1kmyPQC6o0AQdQdc0UWzOdkhwhHC
3CjKET0DFjw1zK/256a19Zjp5kidhKpzlPwIPpNJhapqhJo5eja2qlHQWCFe8n8K
QMJ95qJjyVZ+SeDkQVS/aGc2LVTIkuGGoDnAXWTGm/G2y+Srsg+Frz/Io891HqmT
yYnp6r1f0bm3TMzJetO6a2fDKfZ2T0S/dysrKueHpYQePTJgjfLjPWUUriuYKipu
984H8BTDBIOmyQ/tQE/cmYWOf6/KbR6EOogUgoLKkRXloXdTLBxitzs+ahXb/FCE
FDlG/FeYjhXiTNOjdk28Kt4wmX/xWGd+qSoUA9N4HKuLNNvJQCeK6ueg5MLjs9gq
Kpk9t+7M6gMYemWt0lBgqe6wp/iLF2guwXioZnQuq0z+OOVie/DCdY3nbEQn1jGM
olsgYuJJHa6ua0lHf/BTkyjeDa9XQeIRe4eLXTU7jPhPpE3g+jxT8m49i96bqOpg
eUSFEbo76SC48NgpxG/bAKFaxOS12KL1+t49gitfxxlWB+74bmOKthtCwlvMoKwe
5CulhsMxs+TynWiK6PfIaUmfu9OmhPN+766r+TBQ1OM9n2C47If+BS5BfcbSu5+s
PPcXudlHc2+Fs/0LKZMBJP9ydYfdfem8RuscWqgUwWKq5zX0lATpKN9lqBml+sPv
XUSG51rWWrcodTfd+DBt2IpXf3v4fKD9rKetLuzAw/Bs6xsNo07Zk1AcZ/af77nc
Z8imAugXjx2ZXHYd6IMVF/bka+6wsQb9qEHyv9c/l4mUqnJLpCXcgtVjBhr3Tr3O
Tlkfm6j6sP0LRVhg6aSKBR+axGTCwsw8dSLQSR1Dbo8gqYoVZ+3Oxo/vTL7FmlSy
hZtVuvapec2mMpRa7JVqgXlXFrM6sYRbSkIT/DJckHCo6DNVyHuSSxpVdinuy4pd
TEyRk5QsJhO/xEbcGhB0yRc05tBQ4SI+SKHDm4gmJRO6rcM/4w3GZAIfxqLc94Ja
HtxvNGkLvCyEF5dFkvE7PsV8tRV+CNGAnKGZdj2AaNKG+c8W0HvVx4jVqkekuMV1
IftedFiS3prKqMNC1+CY2SuzRkGd/YSxxYLctNII/6hsWvsFfW59uLeImHeZs9ya
I1Al2/PdWbkFcUK/fvCVI9VAGlQWo96QMtgjRuyPPqz/BZMgj44hVvAzgb8Avb7E
MVmf2bRPX7uNfzH+btf+MaMyR4xSIw08LOVID2fqGRqx05XmlFrHV/pZUSpUPjvc
T1FHS7U5c5kLV4uFaZQRHoTwqqUOUYk3DVl9MHXoifk6neknFULgSqqJTJn9219F
iIXRj8YYXYtV9hZGB0lVTDc0LH/va5xqklcv1XI/HbsDQ/pboYZYJf0CrfoSrAdI
6wz1gVsrb6CnuONq3+JlYykd6nVMlt0bf3zzX83L0vMSKo/WQczIwgbBzYPWUk3k
S4F9PabKTX2Q2ti3y4vYsK9qOGJow1TPiof3eDRAFNl3StBWt/n66KIcin+9tcpL
MjaNrRxQq5X7ntQoKKRhPGdyiNCAeViN5SD/phK2TxuVV8h1gMPz/5MaIoK4Nb3e
2/8ptmH8H8ycFlzabcKQX/f3S/QfbAqecTGUmnqhoyqbVBf7uVzf95McTLasLQkF
66XIRp0MdQGuV2R/iIzEVMIdBzQ6DGCkYvgNGaCkFsm+eN205+TpqeaR3K/ZjeaP
QlyKQttz5EOt5pJSuD4g7PX2lS6g1tYpSajWtgEBTKlowzqrWorSEz5RN6xPb93R
bss5/KarTTxeTzLEpXhskX50lV/apxQdRqAISXiNYZlsQOHwmsbP4Nm1GC4KQIoH
oee8eF//4/VAzB0KfmqmX9mNDaMezebwtPl7TZVmZmAxcMe9KD9LcE3phdNlh+RN
cceZWKJw1COGma9zj38dlIPoIB4Nl2jhkQcjgrI7df4z5qWLKBSi+gkL0UmtkRy2
2hBFXKDZhGlDD2zGxHYta2pquTI5W0h0erMxuxy+P1ejy5a26FJfZrGYNR68cgJx
6uunY2O/ougqcp2FnThjGed7BSmU4Y2jBYsbrj8JmX3/TTOTNOmdWdsp8kkcP7rW
2U7vJqZeSPz9yI/j7PIbdFdGUrXVVwWXySsV+Xetr325CrNM5rRsRYKty3MerzQi
45JVtoNwES9VcTHp9jNi1CoiHy96RvwlEypZVDueswdzpj+2iqs0Au5CZWgkrWlG
BsIeRFhqa4hy6ohGxDZwMJWSL3Qh19/DI9sJM+isbfy/QrYs1LqS+RzgnI02W1no
X2byMr7WhDYAKtH4mDaCR5AxeD5tZArI33r9V4o8dYQp+hVjWEu8Yjzi7UVFDoMj
L2JcrKKa8WMHm92VWTFZ14MOR3c/a9bdrOFACoeiHc3FH3J30nZKThGYIwdbp9Cf
ZyCy62MuxND6Lwj1OaeS2Me2P/pL37+4uoGJI1jErz1AknG54MJtR2Ky2wFvJ76Y
joc4utLjYzchUI02e2K6Hjgt7Ev90oE1dd1BFN/OlfSC7X0J+XeKJo7IeNlfSJlQ
EYcaSSEVJY2w1wajRPqFPYlQWXLRbJpRI9fkg4y1iQkgQFjfMt5T1mIjk0zxF3wF
tLvwsJ2mLyVqH0l1QMEC+2/vpL3MfzYGJTZt8NPGq/qDZ16npd/9s9F/+VlfruKz
Pq0aHzgcDCb830j1YiRdZmWjq/C24zcMnNSn+MwTLK0bkKsvR3mn2unJ/UCLwicK
a9CFN437Qc0OOUy3pJ8wJYtcwKOdvoKKcwPrRxpK+ha0ComI9pTq887EOb2Wsw6N
XGZkfUdL4AExYErA7qXqSbtuV/d0YN0r9u0RDdlVqZRnbymn5SJCWtLfs6Zx+lrW
85HAVgh0KSmWM4ne9IwUcTdYUssU3ei/mx9/xrGDC/Yj4scOm5xOm2MqzgMSkOpU
uvZo3kZNA+EhSiCjDOKS54XQ2TTyvtRT/cqGQd13cd99yvVXslJcbEATx2BpIEYH
nPpJAtbwmYFwXy9gvPbzCOheSAIcjSYChFSttZvzepIAsJ5nxCnu9iGEOQBIZZFT
TMoHjhVD99arOPbY7KK7k0+8MKqYrljQSWMjdPA+QqqCianamy17vR07nzY3IgZp
3wGjkE8kNOwStSSOre3hI33Jyfwzy0lG018sgZzaOJIKmjzaPq33slLkDIvrLcTl
LAn9C/kCNdDmzK2InvPyKqfYZlvIEeRwZBP4db+p3gatsF0afnE+ZFUapXSk0HzE
G4PSrD30B+wn55epkNMjYiox+vXKhQOaZcmiM04Nw3SToWZntAiiA6ggNU5NMsK7
73J+vdjLvCC7nwGwA/VTYBI56D0D+TKSXHZhpF8+AmF4aW74QkCt/a9PNMRTG9pv
okK/Ko6y0UMQyTt4EWTl+gGS4zCr5/ctwBTnyqvKGbVnwXrJ3P82ynbJ5f5m2lzl
e3OhalRFTfQQtrPRZcIEHwP9tGPJQ0SXCi3FBNEhIdpNtwxfCZsgVdI6/kWY67lh
jsFqPWgxDqAzGaeOywmlYVFwcH5aH7F+H5C/W3vAyZSBAdX4QZLC61YJUp6gwD0K
Dj9aLnRxiFhQoxxIsVQGNOZtdbqgECxelq8h9zcIS+ihecyL959dtpBCB4MqXZeE
V5snhf8sXYcKlkziFzj87BPM/nt+rbHrSQpG7uKdZdN37OHgxBBrElETmC2iZflV
VSMgu+p2uVB6opO1rDHX1nIW4pnS4HP6T6SR7aShWmGbSdM/wE9N13upjyfmDJ/7
7Q0eyuY95ZqC2qcDUt0FmrHAupKJjAJeL+QzlgWIx2ZQ5xLROOkx66UavWa3YUAi
2OThFEcOkjGUH9/0GxqxuY+VqtKzUO4fcOsolEKz9HHp0UCeoImrSSQsTf33PEuw
7Os6ITcjnnHIpa35J2YoC9pww3QJnkIWjvIfMxQz9PAeRil4jta9YjxgBU4nWJat
eWSKosD9Of1dgqslt8TLYVm9KyvATq5YUX7UGn62M1IQ7HLPi472Hviz8EyaFB25
z6kagXrZGgDkQxwnrJEC2qklIJtc8yrAM/CIJKQ5lYmXVlitVGncxfB2y5YGQk8J
jsYIw0rg/Rev63DKYtY6adBPBg2UjwLmCYgJWt7zadqD8g9z2PIT8ESqUqmjRz33
2JyVCSiZi9dFSE/2kp09yvnQ45xz995WEYNB5lAzpmnLTZhz7fD9EyNLIuDmbfMM
jPkyTig5QSzHA6ZNoFPuadFq+CgLrTE8ZWmgBRDqfmgKre97hIaZ9rcgOsFd/wN3
S5o+eR5pRkXExlbSlQEbi8dYfLrxOn/HUuFzVbviPL4RHsyxsfNFP7GgEC/iwpY8
ZNDpRBXV1fsHW23PJbX3Hnfg8gyHFgnLlUaWJBc8Pwb2qYlUYavyTLUPSHxy795G
FRsxQ6xZTMc9tlL1NqKlWJ9FImEwZ+Vm5X1Mf/5lBEZcP0kKNHf2SxMOuPootQdR
5du/RwArRGJnWNcnNkVHyNodtVShLDAym9I5s01Acoz/Co3oaqKcUL7plRiK4W/K
HNfMXugU2FIlfKD0xnMoQ9Ybrjy3afnzuEiuIbqfxaNLXq16M7TG8Iq/WOsFi0Hr
batOclnJETow964ELG4O82n/r2y4tWayKZWkDDb3wX2q0sRkmRwCw0Z252NSxa4o
2RtAJ2chYdJhJ5m8NUADTCPf2Yf255n628r7QfuIE8dm2J7lPrvk3f3VgWsA11V2
1e44P9v94rH3sQ4HWy0JI7H1GJ+E8SMfOFzQDJUNEcS8E/2wS68yYxXShOSRuhXP
cGE2tEpou/xIWhKypT2BQ3kJZ7fejcvwXWHX5wwZVlDXklnusjiCbaL5QltweXuE
lJMWEdY7LDqmCWaIxa0vBLD1Oke4E29Z90Amg2aasmD9dGagwpcUYuFJa4h3rQnx
O/MhpOFm+nHdAfmvTiuT8br7IpQgsPh6PnweCfztMU1VXcUp15VP8fjii73AN6ex
w3WDprTULZ4X6dP4itCPWVEXV2iB0qkh+JbX3qhmX5QfDkHnoKkgj51CsAnjFXx+
pqewlklGWme+VLuxctbdrP206/oIUQ3Dx6o6U4+bdrMZBtuvmSGED4QDH+Ak8KhG
OEm9nUFLEKV0y7v2U9IP/SHc/vzWjPwUJP8APVrldFinslIH8Ep8t55uTpJbwiJh
CXYcDMQO/RCmBDH3LJ6DG+7Fc6JEyDB6PQMUGfeM9rU=

`pragma protect end_protected
