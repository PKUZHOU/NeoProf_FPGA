`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
fFKA+SQJCxrszxASjDp46DHqIvVYH/VpwnSX+jJCwF89hkj/b/K7ec83iGXpigLI
qaLQPp41iBtniOsRRTNDlvYz6FIv1ivFye+kmtWvhKFZP6H/uh7rZfS0D+ENPl9K
lSM9SbZhmyCSaid9+Hkq67AJpS4XbKxqEVp5O+DYQn0=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 81536), data_block
SmyqOofctGojV4PEKkTI+qhF+J01QYe/lY/g1S1fMuj+JCUr1hYJZEhylCByYxwf
uJLw3T8vDFv3oSx09AP88BaOthz9BdXjpBCfufzD5/TRtVQ2WWpI6IkYlK9xJqGv
ZS9WogLuGo/05ooGtCl31VaD+WvN5Jpa64Klx+m9asX8qm9IqJS/4ZT3j9Z0oyYP
MpmXw0IDB020MI6I/5n/Sgj5y5L9jxHbmewGUxTKwxwkVwg/zSeqw3o0SZeKdtb7
2m4MoOO6Y9NeuyEAszB22ZRPwscZU1yBb+p6rD59tBkt0Q7odl/LL5tjhCPfNk8e
MceL3Nmou1o03SRctrGXEo2RkVSPrAMFIsUGWjzbbGn7/TpTPgzotQ2mdUHqNw2H
zNF3qD7NSFaB9Rouwssm/sy1tSYxn7HR31PS7nT/duaPPbHUT4HyFBdslQ7fu4yS
aXzwhwbAGmdJwtFRvWUBTEzLHVYzgv4TfiERF4dPmHps0t4b6xzHe7nJqkKeBHGQ
8M6ZCJ6SU9iKcnV/2lWNR6hN1dZqsmcWgSBEd5GtwWpwOlNnUlM9wxetQqqBLFP5
M7V10Brs+3YaUjboFxHVe65VTInbOPXO3rg3dFqg39V//MoiK3rUfANhBPjJXBuR
GuxPdDk1O3cqYjiolQ0vS1YQOxvDs0J1N7luejpAxSH1xZichjxlHrFP4K2ajkf6
ifeG37VAzb6KYeHrH2yUrb8X0bbMOjVDihVFK5lQpfjgfMWg/X6VfPSz6s4owuN/
6aF0Ht0bPYgTR9rBggDpLV09oE+wjUxgORoa5HU3Gus8bo3oNmQupwsO6lOO0ZWr
eiSrHXtZHFrNxr9kGK2lzpyRJnlkW+1/Yx0QdadUJ6hQJp8DnNkoViO6L5poWSIE
JKg1rOgJmE3jC4eIsML75AH2TBOqKtm3umDe5M0TkXkXYVVLoQM3q31efdJW0ek0
cseGc3w86xbEJTykgQqwYgc1SMYff7eDTGNlWyTCIj/xo+P+qQqnPDgJ1WDbwzmh
Jv1gkat/fYr8qki/NhzQvMdqhzrZzr7leFTfAtVD2eR0Xqv7s/BHki1gRcJPsuX7
UGMl4Q8V5lX3MmyAp3UaZwHQv/pb15p5ds3ZaZ5/y3x/9KhThD3ZjTxual1fh/+f
LBvta+EgiR/t6wd0hJlQUWIn8OI6669OL+0NEybCFun3BM3+mIDHPRLniN3i8E2f
SZR0JKDteap+8onp5RFDDuWjXfIAgkc5V3rYkQ4UCKqB/9vHVEtwFk65C+mGNUbr
Rffsh4L7+4BH8uijiVmPgRbqAIVxYAZbVgeJKpp5AeuE4sYGuY9VY/WSMLzCrSbr
eWhpUGCklhjP4ovPRoKoPf5F05SvpLR91BbbVTXMivPhsTNhUaLpA/uDRJW6YqLp
RlSWDJxPEyqT5oiQIuuj//csmbfHCGtiFhTulL2adV2bIZBzVH9sU3TBs6QrPOA8
BI24cQKait6PnDnx4iDJ9AIYSBMsm0B1hxceD0fnpl4lSD0KFPbsGTo0V/cg++WE
vx5cpL/RH0tjm+9B2GM9k87dlqGTawiKxE5rDXV9t/DEH/noahHJM3aYMcrvJ+Fa
exkXE4h49zXRCIe5p+qN8BHxNRumyOvRNM8rQVgo6DTONNsQZCk+clgD1zUzd1Rv
+IUMWE/IbwmVwGf8RYxx0TiGPUFX14q6yFs4VjxAtXNo06d8owcSFHCiWNpYuq8e
lqmWs4bqcYRuc/wYRof7IKOFBJB1OcNrsfKyW4t2pVXWebLORh88ut/3Px07INsd
wIfthNrXw9le+6hNF3hMy/SO9I2pyD5QyRJkk+gydn8cyZ3UzCjWrj6FqRcTSuq5
SaIRtyUh5NpsICmdYzpm7orJEImaYzUTMwyDtYbBmU9Nes4VVrRdyBi/XLrDnIS5
/GB2khJ0h7F6toQ6Ot8qlDHfTBCrSj7GHBdoB9v+rBCx210j8DQVHZSB+Oaojios
MoHk5HMrIZfCOWGjgPa8b5pGVyGGvQg9T620V7yTBDhtQMtqTvJ9aiN5kD3MGChf
RtzpuFqCGtKbEK1kfFSTo60IKR5Ls42s4ItYgpHtwG46dyCC7jrp9eLqAviGaaCT
pxFXaMhseJDdQ3p7yAZS2wjPZJunRlkhQ7D7w3/KeTTRuG6w7AIaHPYTNAbKNaV2
YTOSkGV96B+u4OHhpqD7f9eKKR2wqx+t1vin+XC7YEG367XWHQsjxZMQXMB5ZIBO
vs79ofCGpH9EBWLXDDp/I0g6ZteEU7NXMwkk1BQ9zPPwwEqN5PajUn2Z81ACdOwr
sG878MOyf0GvSbF7HP0PERSllEmSnUi6fN/d3TFnZ+TxEGegGkVDIDgagdefc+gi
rbJH8zelJKMqXqJWnzj0mokIlF6AeAmCbFcnZEf8KfujD+Ufccw+JMxYS7gzFZIU
bDYO37oNFGlEW7A/SP2pCzgbyMhVv4gnu2MuSNtwLuKH8FMh8rwSO/8hu0DlFN8U
lCfcdBjuO057Bp7bS3n7KEqJhkUfqrJxB0rN5y1qnAPphxZrdpRHUXXGr2XTq6tU
r4Y8WNyg/RddBWm7B75dompM2NRePBtvcKlgOD86lRfTowTJkWjaAg85JbvP4irf
n2ZsBryTibTYcFCQm3L0LdFsyIU/gyR7oZy7jm6sgL1uPTrkxWA7CtaIAZ1kEeVj
pY/ZigTP6V0lYLHQMJR901lixphPfaDsuJydxHWuREfrxHjeTZlTRmoDqKnpZASs
03uaNd3n4goibJYnsznKSUTgMWgaI5mHLTdtOqQ5LThbhTEBk9Akc/Q/zEQNaIpO
VOJ8UEkC8r8iotfUJYz7r/qACvosGA+ZlkDeiQyxz2/TYZ1YY8UMeMDWk4FFcfDD
X0755UjP52Al5vRsDOdoWebpdsDbtrBpJlwiBsN/MH3ZJfgFdKfUUJwjDLxySxgb
7FHqcRHtXbCjTwD8ju2YQ+Q7MVj296JdeiE3L+0g7ujvhGdQEZi9eUoz/2Rl5iUI
F7w3oU6biZrPBdyZAvBre5jQt0/nFieZ/71yV+fMLi/uqEfWZ+ACEOc0ojC9xz67
7sbnF1GVyBUMNQ/CrgaZkVyxF2DCHVFAOdMEamnngKaLkaUmczUVPCWfx0x2IQ5r
A0WUuipkpw4SNYc0dHUXvHuji1Q+cLTM8vxH+GzsFoD9qGejcx4BxmEvY9ZJgN54
+nK19hp8syDeeRHmOH1EI07AJn+lrHeGwXid0FCqb91e/+cfX11yVnhzMnqr8/xl
/pOH5fRG5LdwwFiiTxkHDCFe59T9HRJRD2krmjM9mKUiaIzBZA1tdOV7FUpybIjD
bTsk/YEphZOY+XpMoOkglbLMLv1v0JNPfT5Ar3SLNk4GvPzhSJFniDp6ruzKKtSa
wekrE60B3Bi7JqjSHz2I8JM03m8/ZZ9+tnhN5+ekE6egxW1fK426RwZdlibaZU3x
2+cDdc02Khl5MX7GbMQYOYvbsCSli4XnJoqPBZYwL0H6InkCVmh7RES5zNUF/KTa
knzLUB31HLCKlK8kiB0DTt4+odLFKMvKlHYvLB9N6Fkuj7W9ljwLrtjuK7ev+HlI
kSxkTCsByaJqZc7tVKKrRBRa6q8sDPHbKqhswcf3PdTQ0p6Fitp/iphPJ5yLsGBQ
XrtzlzESTw0w8t8hSlvtYPWfwlEDFz0ytWnPv113s3KWYbTyOqqMfXWvmuCFWdqX
KcRdkZ/Rsp1TTEgxRDEU79Uq1RslEoQYQ50qCt0yjntMekR+UtpA0invgY9F7HLg
qae1kpmAZ/C5j3dL7QNvqY97fOfeygNvqJT//XRb4upAHxWaTPdIqwpqklaWl7Zr
vE39ucqhmex45YX1sgfztmFLV7VSfhQnV+779ZyDv47x28F/5WT7/mFfkvmYuFhY
Orx1kjbEb4TGjWemBduatRqKk2C36fzgUuVDcXeYTMJQ4FGdHgtj9ZjCdcyOGolR
iCsYrzj4cT5STINFTTYxjsk2CYbZ+D9BUkGVePucUaQP7hTCGmllA1yJFHAED8so
wjcfBTlPZl5LtVEfU+267CfSLFQL6XFU6+Rk/1cRjPsALtaEBNLZbe2Xwii7mCyH
6WJTeLtDn587ebDgMc9LvEpMSo3yd8E/fL885Da/k+vihP7m7Ukkco/63Pzh/sW7
i9kEfBHuX9BM12RafB3sNTeVv7oT8O/QH457JdMzVdiBjNsnChFwNSAQIo8q76Zf
jLmsPkzsR40ui8HDiEH0HzK4tqmeUltqgJDtphT04eDqRnJDKRI9V0/dNrWoAiAg
ksIm0PWPxWbLnNcaDiPDAYd16Zekq5RND6sV/PSqgsgFUTJHNfe5xdjvBNO7Kyx9
sNuDaxUyMhpZA3DZjSkSMHR2AvhqmGkjUaSgzSpAZWr+rx1znBGXIcqr7S5YbchI
P6bTsnchIJFVBeKOKEVad+CKu0+R1AOictrq/OaB38ZlivKILizjJn5pfngAhQMp
EwsV+l3WMl71CKmwgF/1088GgbAHgAzMDF6SE+bC5TOxm2WDi4J8DM8DduEHRz5y
vZpX7YARPejFHYX936DsglyJDYZPi/FEtrOoWqY5c2lFOnOKmPenaASzmZ47sJ98
VpBP59pb7pmNFNp1uQpbBfkFENIUkzQ+zIioEDEMCjZmgqwjvSA4j1EgbRtRHr9u
7gEAybGmWh43fIcHoMdlkgLoG6xsXakbLo6OQr1eHItmAnRQyKyEc8L+RBvQ28dI
m/rQHamXUAGKH8CUK8h0G7nu+Yd21+fRR9wK6SFIRgISZm/AYdUJ4hU7Xp7V+dHR
eOezNoJPbrjByccL6Peiof5ZyebdcqD7Skzz6JfN7Hkq4aKxSwxMPHW3ZlmlCqOL
ARgSPeUsRv/4j7Aeigpii6HCnxY+dr0vBezR5Am6vuyOifMzLPmGOYTIxTqtgkWT
FnBA7FooE/Ce+UATE0NpiRDRoje3uP+yjgDRY4zN78d+7anUkM0Z45LVtdiuuH9l
S2uu7w5jtBWDPDg8O2h/MlMk1qf6rftFy01oDEWgUn4R885E04K4infW7sOJLlsY
1Y24RkPK6UiaDJ/MvBfGYfjPDKj0WKFy+K0+mf8CdwWI2Cks7DqCTrvwhznbU+nE
07HkBEMwCr3tKPI+3H+ZVIhMWGDJ6EJuMgXIN1snET8y0psURtqjD7GGnG7zAvhE
CQfb4dE8Fs/+LNCSAp/kEpUAonYpjFOvZoc9mxilHt3i6Aj8CNXmDislZHz2jr6f
+vDoAO5WXm5HbhkuIIBS5oq62u1Us5p3QPLyGisaHdapuIhy5/+R8lJaciPl4Ygz
wbtCIqqJW6cnz26mtTSHeLxBxEN7LK4Ml1Z+sjo3vpJ4bzI8cbLDnJHfATpHPwrh
D8mtlfoVKapWcayZFBYkbnsiP8yp5rBKI2qsFolsej/qQ5rX31rPCFRgWiYIIKp6
leMdzJxABPxMfsSI7SjPFHJFD+13DdlhmSU7L9V8DUV8rBEURA/qdyrwXf0tOpoi
5myVW9fs72lukcYpKwwtq7lAK1cI9hyHJkUYrgYDVcmncwVwi+4d2JgqbYtu6W42
w4CNKccsZwrVpDBcY71uEbjlESdLCGoghkui26tOi08o1+2xb6SPs+grsE7bL/Lk
Fjz3gjRvgxEKHSq7WbW6SYVQbJbuXwkkzC7h8JQ+CkLmWdl2EIzbpUKrLj9YyXWa
c4TEbVALhQkARjdTGRv0XLC6JD/d4A4sX0E1aMDICQdlWG7Ybv2TgiJdI9EDe/BT
kVQyuwjAWwIRoU5JTjUy+cSq1UCZq8ClpeSPMi68r8RslRrcE/WxBsTO46sxfDNg
p/Ke7uP8omoPS9fsY2NQZBgrgAqjZm3YPHLNus9MhiRWjIh9xqDxI4ZBIV6QQx3/
yM0y26toYbX4G99pkCUfB/JRH8W152JkL4/gH4+T+Z63JRKM1v58fBQA70DcGdFI
10dLPf7x/I81BVlrczypkOmiffz1J/iBPNock0Z8dalg4lt3BOVtkAFfSbH63dLK
OrmMghhznm5/LPJnSXJqVOtGdUVUcqPuKcwC6NyLs7VjiYaqhPpjzq8RUZ/Kt6kU
LLFTP+L9gZQwP1ub8GK0gzDse+4weky+sedKlg2lk2tS4ZTIc3XEQAaoLnbo9zFZ
92CeNgpbpJe8jQSoKGgCupuiPpouLtVrw0VP7w0MkSrOcAcPx/B7u08iLF3EoAnb
4nVViKHQwArAlrEc7ftVsqLNrs+c84lXZoSxwewhZgFffPOukPMd0eq1F4Lg0j5j
pDbIB5iYnom1cq+8Y09BBIMABnnS8Ns/vUaLz1rPwEV0EJAV1fNF5yCYJNhKtTfj
EeA2XTkgKv7q3euS8TJvoNKHCyBEo9o86GW4Ae1pG8m/1zqnF7DgRofBizpiT76r
ViV17vj1JDQ0nB7YBM61Qdo4SMmXFJ/b4pDuZ8Yk5w+BC1Com2wSszvJYuDZJzgb
qwM5Ea2uVP9LqOWB3slMzEASCmCeUaNWnoeTM6mY9etuDfn3EITtoViPp4dNzgVv
Jrquqxglogh5erIs/FOAzXSsc5uhZ60bfnAvJKoTdNNIWFfxXlc2SuUh9gYpjDql
9uX9pmru2iCi+Olv7jCNbWiTClpGkbsi/1L4XGjskcLVbHWEJ2GO4rx8y6cX3hZO
eXSKx1degIu+A9dHWyQzwoTf5UBS0NPa/IDyIv4cr0ctBT/eifsMPoFYBpWgMLwx
erFDn0tqqkxtF0AJ6HqVGoGVp6JihU3HjcrVVX9+LyinNDhyU+ZReBHKhKXqJ9U8
D28g6PhKOI0jGcM5xD9CgnHw9AY26TEL7rsOQjJFA/6Op75MgiRf4Rtg/01Ll4L7
x22FEkJD5H6nOyhQjS/Ig1LWlimJ1qaTx3xKuQL7N0dbcZWlFy7KdKYFTB1Yni5N
CmRXzAH4dd7i6XLnNGXODlt4MljWZM1wfczPRcybLyr5+CY92yk2cwnr52bHTQ/v
I0+LdIg0sCC5gixdeSvSS0PLph7Cbz+MnNcG3aLFHeH9mY6Ghm9a2q3PlbbRjRmU
ysqXEkBGav0y8UUszn03KtKaI/LlQcX9TvY6KKefZK323SGKLTPd+aFGiMi+3PEP
eYwI5sDmA+Jat681+mihadgC60V2Yh4rYFp+V9NBHJFqDM/ELe3CHQ3jXfnRVNs+
E0Ra0cFU0UifM4STuC2Qgwk3N2XlIKqqN19LDf+WKbr16fUEX89Phof0J02QXd9+
jwhX4/ZbirD9UMbme4WFoLYJkB5R/k4Y6s30hlXWrphY+crjEAR3Lx61UbzgwxVr
v0l4xdys5aCMWQ/UhQvK3+nmvNoLHMhLC/OXPun0Vej4gPLP9MXuaAQR6ENONCAT
yM4TqeUT6BwP6+jPB8+2pWIwvHoJLHeVVcE6lJG7br1RdmTPMY3+Lpg8IxPCOVRB
NkHjeQZQA8BWh8Op2KXIiztBczKHScLQNYj7Sz6r31zTK6QlJcbwlpJSj4D8ZRF0
34/96SWyPfI+bY6wB+QE6SCOusuqbfA+GezMhaAVZTPKZTuRjRiT05IfFpOJesFX
urJg0IhykVpHlGz1SgGFGefAMQ+nKzmxliPmBujBffY4vRDQ8VMhM614hhEzVofM
gJybg462nPSRpUw+gnr8/eYCpj9NX5PdviYNXMs+X2GOv873BGgQ9CC1ENXxLuME
y2F4Qz7qSUSMnwo7oji+Yll1cUiLqilIEd/Qevvsb9PnBARX2GbNmvjiPsYMPW1I
/X3Ymqg75HWNbaYSS4h3Gl7YkqPGbZsK9YLtU8FnZzshPO9b/aPmLqH0PX76gwNs
rShAfT3/b50LKWWjDQU+SXJscqRpVc3vlE9lQeJps7AEMWelsnZ8f+jnAILLEMjr
85QV6UmLusZppJjtQEPKRCQX0k4EMCUK1uU8dRZgJdP7dBmJ0A0w0PcEWmipOPdv
/Tlun4EZ6FZd8Uug8AXSWLqgiPw5DIGE4WTLBe7KCOJGKKMBwM2qgGw1IgfamLO5
CoK91xO63zP5b4vBUp9NvUte6TfA4MD7FOGG8UX/SUXyKp6HZ6zrtwoZ/veJsrT6
FOTMTpjnx/bBiiB+WxRbo0Hj8f/omi6a5BieCwpncrsK9h/Ul0NTjbWMQqnHP3XN
tisYIT3mEqDHV5V4k0SRrG98RXDJDsCSwtRuzjrbW5fgSlkulkzApXjZeEJ+dD7i
UQJzZ+t6tjkOM3voRdyD2wCAv5YYe/YMb9W+HnSeOpkUrds+KER4m2/+5c3HYBBr
lV4GZ3Oo12G5ej87n7SCnCBzY8LKf4/qhVQHxHTIxEG2scVyMCZNSPNOsRsq8a7V
fw5voaw5C1dP6vLwc1jBfpwQ7srxJ77+4aBOUp6H+43t1ucT6vcF3eJxAjy47ubs
fE9R8lzhOERLI07XJEWX6f15j8/q+jxRLHlH0baBSo0btR24GjWGZxVIfK4q4DoB
4RzAIexmNCNh5soN25Da4sHhVdbGeGw8rsuomFSy7sp4l5mmx50aATxkquQkddT0
P8rL7/4/Bk5i26s+Oe8WbPqLFT+U/KgCCsBaL4AeS+rU7kyjkZ89gSRIHVV4jxtX
54/NZ90wfmBUrvKxvqwl122XZTvHDd+uQ3EjlGbdzyK4MYcwiVDwefzyXk2yR5uX
MwnUySVf2w3GMZMKuXFQPwKtRTQqxqeBksi7OO/OTP0CMa4jk+daokczQNBtbQpo
PDeZyAvduEvwRDDCY+X/QtmKR91IXusQSoMKkyAJb5e17zdeoMeFKe7VNaPTzxVQ
rsDO1iahO9Qqbke21hHf2pKFfrOIm/nlrbpD0ZYHaPqsguJUjVWf2hDPNNIwBL91
cjSqXynt+4SLXfriXBwikzr9IeTVzzrYj+IZ0tbMrr3GoWpd8ySD5/GAht9bhok4
J8UnXoXAtYw3uNxsyZbaZMQY2bO8krooERGsX/1GZNAgp9LL1zSU8a1beDTStea3
j9uFkNE25xJc2G5HS5wqOKwq/bMC2YVGXnRvfTrpKvUswsz+Q50fVvck+ONLgFRY
N7kvu+djArSoaBBixEDTHWaQ/bKJUtC1Mx+aP6AlAzxqIj9OndeDm9cXYhrYBNJ4
6kwrrVARZbYIfelY6IP/GBrurcu/rvWAsmXaFeciPf141sakOJJQv5kuO9BbQkyN
opU5HxJeEc0EsxG/YafDbYuU+nBFSjBJQo+burGoJbPnKTmYeINADd5Khx0aud10
YRPEyc1b/PQbxg0xgZcdg998aHZOx7nPFKbrDb/eU78pEnu19H/5jXJYw1nSgaAb
zdS5ooJUxrH2ye4+MvutCB1rPwc0ebAYyYlYRJ+ObABNSGZV8xjOyvXw6u5Py8/v
GF/6aUl2otxVvl1s3/TBjfZ//va9Rn7eLdvVEIyM7FXmM2Bx7MHfGmrs5oNua6Ni
caP8kjKcJVefrPsFNmlLVSaJBSH9a3CY/LOEUy1x07+YCMuoHVS0i3oIGjNP8GU9
8BvpXyjwCgU1v7KKwio19DbhsX6uoq8sRpywMsrCLd0qcsrVFH+g3X99s/53TU0s
Y8LKuS9Ghu9NJuTKjphSA1x3C/CLZY8oAjkfyPYVVk9gsiv0Up7u3kGI3ilp10l2
QybgIXMoorTKNSENMesyiPWg4Kg8OgVuXlf+9zoZZlt1Ow046QTYJ3CMKCZSIPs4
WHoxNBTvsHHbnw9OUZEjBrvDv9zV3WaWHbVLbfeFfSeMKmym+3bFPpMgKrWVdd/S
QYyuutNyljDdzFHTpTPg5tcKVRCtSf8e+ygKksyTckevFvq+hDgVe5STbHdOfoTe
bPlE9V72MkYB/k7gSMtyBbyrBZ89tlybv20OP639+34coKD/z0D7JvA91b5Nt/LW
GT59bqW1p3t/Q+bZ4PMrn6ouCu3KAvDaJRWEs8ERO6XwbyGSWtUfIncSOixjVX59
fKBbMiXmrcib36FAIS1brd7yBAlN9N5D20JvnaL1b1kDafS3PiFjmMcvqa2RF5JH
5te0kGwEiXWRGamyUGqjUJaFqFseqflw/czXrPq4WsSa97Ruemc8d7c9xxCaArg/
R6SDBV4iJP0YR8g0bilDZP5DUFdfuI4fewqOSGmh2N4tHCab62Kd0H1E+qkuppfq
t9b5eR4jhRA26JCFLf9nF+aQMOAa9kHE/kp8UvDM4+Nr+WoHmHu+z/kufYDvIzBr
p+NH9FSQ7Xs0xEnlPEP97QBZwDRGRgc7MI2XZZD0CmvLssoGxar6wZsrjYTExgeq
fOm+POyZHt2WTDhPTwYacGZU7be3ArtelYOizHyIY8GcUeeMdqQmMYCACNpnPVip
25RQzjxSRiBHdwDp2UipLcq/fNeMCju8uXGLAdjOsQpdOeURr8+TMpVw+yJEA7/X
WuF2GrOZxr8xwluW+4wRVLV5Pb0xFMcjF4ce/YE6RUMaQUt54AKJYrFEGFG8iw+2
m0krNrZfv2Q/Yc6X4o+Z8H7RTIC5wSm/a/kPTTvjdv8oyvk1YeLMB471JSX5L3qK
phwCSWQ287MVSGkXv9g3D3ShAburouhdOVYhVL5/wcdmZvkLRO2sVsh9/F2ugUL7
7o42bqm9MaoiXBLGkFIFNHiDReWtb3ZfHXswOR8L5qVQQ4uHhqqtY+x4L9VAhvwt
n6gy6KOYpeDxMokGA9V0s3272BVRHwnzM1Q3jUxp6tI8/nTxxaJH9/F/rhhSRp7n
kic9v6xvd8XyTfkbLVjEZ1L1JhOXoz3Ve0J7ycUbRCyELvpKOg5IIRD99fMf0X8L
OIsRr5tYP7fCEj/C/slRENJllZtoeFoL8GKgjmTG16NnIqcU859+z/n4xoJZmTke
hYKRLQRofeAyxxvmI8hef43Tu7rRDSr4jFgs0HYGuLYVos5JwmR2hSH+czy0B4/F
ny2XEOGKnAKlZ3+/xtqPIs29KEP8PxxC6OfPpHKIC48a9a3VvB+0L8UT36Mpkuu9
sFlLd6bU080pephxnCeTJ7ZLC9pr/Jsrh5taxVu2hEkQCS7DWBn7sXCXbKPkdtBC
89/TgZeeV1DZ/HuA6AUPYGPpJPcu/g9jKA/SrISpnQGbBUw/80gZ0qqy5xel+Pqy
bCCtdyXZSkLNxHmpkYdR6wKzPGh9LR3bt7TfJnp6mxcTgMmXm1SFmnYouh+gwIA4
dBO/67tRmcCOsxvW0n6YUcyB+mSnjUyox9MWDDVKtOlGoPfvliOsU7c5WYCYAa5g
i6iFPFzAM37tdojnjYvUlRQ3QlZNvq/UV0p5Vjb34wFOC6OjJBoV0KrBryPCxB40
12aCUIWA1tpsOy6/XqmByJ7rnqTyRVnGRjghVc+Gyo0nD8C2VUn7YfcxK/OFUKvO
wL92QJ22/My7Y6WM3XRklJnu+bHc0nFNCC3Yn3HKw0s8NSnOV2Wg26uMcmsNuXWO
B9trGPPKFb8hftTA1ELH6JzjXa9zjfqPCh/9qztsaoyJpiylIOpELhqySYPTGhPX
5OMYpfEnxS4s7Y33+g2iwXXKVKJXAGbTPuIOEWhOVxvyqRYTu8UkPS8mA3Zamy+1
VybO+QSyGqT5xVjMVFE5gC6QXgQlIEguVuUG2N7hUc9hZTUwoaIN+IJ9Z9PpmRsL
HsKJbCiYCmdWjLpp9yz6EJEz56CPiDuJw7/VYxQpK367NBOAe8kfivVsspgc3QDE
hj0pC/vI4LJCzp6tNY9mrb0h2iHG/Q5zYz4GfwgjaWuKMAQNa1piJsEdMXuljx6F
8HUiWU3qcL698iev6IZl9OCXl9okBLvdcsSQDPBZSn9fnzdYHp/ihjE0gRScqnn+
gZcfiKsnY0o+ok7nmsZgZjkcmIMmFJn4RylxzUOXngaqezjEPQLNdlf+zP7rGF+h
NxISri74C/pgrKPaMYZHBxOdeNpKoo/9NXJ9FI6bqXAu9E7ycnDJPP+x1tlM/Ajl
QtqQdRtLD23/vFofcNsDJu9ZiyNgKGTOe7i1QfuTFiT5Ogv0w0SkiTLJCHESpT55
4PrJaNvAG9iACLqqV+WeeWa6gQaNDO/thIotSR+wCJHAZst3r4kSl4DIwYDWRvvW
kZyysGp8HkOuRcspR0R/lbIIfWzivl9yEk1G7Jj5m4AUgE7Qk0sAR/bkRGb69WIt
m/W++Cb3AeLubw3EcjGpZZ4PViYtFO5kNnSKlc7pYgFATgIoGCQCGlS/O4fRfrAD
R3k7EtkCFrmFuKcWVDQgDB6E9IclKLwluAJLBczubAV8MFMsLOKYLk6nPHOdnul+
HbsrRWDnMrynC3uPMvFpVnF9pX2Ake7risfvS9cPBzhQSJA7FZ8dFs9Rtp6SCzXS
gCDHcXEi6sIh8h6Ksu2G46r0m9EXbbpdVxPbOnesf8b7gTn67RU+nqiB9EFOnCX9
fe+3zhXX7YBnbbOAvDTfJHma6CXBjMmSuoGorYE7sN9NqhUnneHveekoKAVEaW1v
K3Js9xH0VS3k0kJ++HE/M8NSyJDnjbkNVhGOznT02UV5b2QD4KRMR7A/tjyN7OfP
F2CvbPwRIzmMd2f8K0XI6r1PiIvxqEWMndSL1h/Apvm6vRQG5oPsO0YhOkNn3B6U
ym5nbNMZGanlt2ohGleG5C+ykgfGGcwK3BiWI5pTVfAqJRvKk9cx97ljzZ941z5y
FKuUKNR4ZSVlBeFCighO6YSreyJuZxuvsoy5ig/CH/iN1lJ4IPToKnq0cFECHShb
gfLILFiVZ7xegnX9b93S4ArrdYPjUtOoNcDawpUmfxjcQvDueJ1UnKbOBdm18JIF
ZydhiZTMvvH3QyjyUHtzWSm+BHryumC3JToROE49m0LnUgu2bJn+WOZJ5Lcw0RDj
wckfhYLjjU6MsQxbHZRiJpwK/0CeJ3pncWi1oilctpcWl3zhCFOHvMmDpPna/8kG
+ZP9z0gsmYhVGuPiYTT2T/ms2r1lbVgFqZbkKB3VKRxWu4P8Gj9QrZykqyD76Ukh
mrxWI/JlZUYEGN4Zkvy901x3DBX3bi7r6Fb1iH1T3P3x1oB1Ud85VrkTm0iZvZ3F
1ioINvcfB0mA3znf5jd15gTfide7wsClCGJJrFjwXbgzKcAZkiTrQPs1ioLrSqVh
XcdX4RI/QTzpdhsxAJ/9VXJej9hK4DuzuuAUtGS2phNZP0uXewb58xOqRVqvyaj3
/cS1v82CDR0P1DgcoKEN24qIjvHG58Pc4IuRRgI5Wvm+Tk++rU5oz84DQCXnYDKC
LdqMBN3iC9lpOZXFMCAShwiSN+U4XGNvNBX8T9iu8IC7S8zH19IMG7Ean/l1EnBT
3NMKEvZEIvMc5LtQJaqXABSxRWpUgAmRX9dRCJLjdKj5d19mgr81OD11ydcqFkZk
YwT9n06vJ/9QYj2rJe22PFS9AO3gUyXFe1dW06ik/MhMQC+2lydRNL/f8SNMeYpK
lNi+W6VBTO3wGwsUL202WrIxX58csWdTRy4q0M9Q9HZNKAh1rfVFyhfb3Hp2fGAd
5hVZPOsyE4EbesO9cq4RrwnXL44tCAFa77JrXVfhxGyvD2Mh8wmAzwTUeqB0jWd1
KoKDj8pOtUulZPTQdl1LK0lLMNAg2K1U0T8eVqESxF7aZ/hNGMNxVjsDTN4KXJfy
VzEjL4qFgo2S4TWanG7D8NKLzfTISetNdI7gc8N3fyAPeMo/9W3HBxzh1aiP3QYR
wGcG9kK9aiJkPUfWDmtBum2qTJuMYeyt/3UkFrWXEYPjDOlzhb/pm5ZM4Cp1HHTt
/DEtqPXL8gkDbcwf21Wi4tMvLIAsPqtjNnR8KtuNyyKZUnowbbb22yDr02GOWJdP
bwuRbLwOg8mzUp9lDRvkLfr4+uZLF/Sv3bBpPrrnf/HMpVpu11/Uwu5VpVNipK0j
Eg4crWTHlWJVBUBP2vYxDO+jBtCG5tvIO8tmTeHBPvK1boRedh++4zaPH1DE7TEw
QeGptQm/MpHdQ/BuF0YRvUHl2xsHNnhTj3HFHC7qy8q/QKcgToojQp9Vk8p72SAw
FcsvfGbqBZcBM5pXF9QpCzxI+8q713ie9FNfQkWqgXZ1JDNFDykQ1GA3I9T1frfA
SgrIQbR8D25hhoHUs8S0udiBhlGgETl7UtlAnaMeR9tPe4eUthoV9W+WIOJjMsUj
aDr4RHJJvg/mP9y2Ae3ntwBgOJK8cIQ6HFkVTCSgqIhtH8y/Mv2PsOZ60FWuE5TH
/rqYgiTVRV/VLyz8a+SHb9/Fatf4l8OYX+OoY+fTs675grS76G1CtzNBA/Jj5jzo
j/jusMp5+9NTnDF5oynR07vc3xzu54dRSHMUz8ZWdhcqjizHooAeMMQEnRU/KAm9
5KnVZCgteMnJOgXsmNWewYNaY8hkQBjFLqgZuQnfCNnAIjZMLz8oH4Mu1Z7djv5W
wdjZjQPIi0BR5oBIphxdBFX8b4Sk/Ei2h4rnQ/2PjA0aBgIACA8kz2k7k/TL4vuk
cdrQ5fxa3hM3BoLa5FolRc2Lgettk9nCYv0Me1CDhdMHb7ZH4citXLzUi+FRQ5IH
iJ9NWmhtF4iyRncrq5mDztIqevxadACiTbi6Ul4acIeGzYJx+5eWdq2WIOMFECp5
qsXzhU2UypwRhc6YACYoYuNq7W1H7s0sOYPtOU/p6G8+A+RVVkWaPoM5d5u0BoeY
Mo81BMS5D0/8yEmTqyvY5i4NnqHnNeDcEausDp0faIj0DMEd7E/BGeu+uLF8RwcP
mmG2SdGaiXJjWUwc4Uc+MB1WsLi4IkF0RkUy1MSD0PagqpFDfq+sUwTsFt3IdJsY
ebtjVYPbCV6F2mNgY9IyER124cZUCoU6aFO/YfpPs/bi7krE7Hg9St/g6s0sA7jW
Z5X74X0K6p3JPXyCn6o52RLvUoYokaNwuy0OpUWlvfuB5FVrJpJCteDWqzcHw1uC
wiuodmYPblXUUdv4mHMRR/hkW4CeP7QVUNE8brBZNGBt++QtTSOYUB1WHv0NU63r
DPTGzlYp33pR5KUH9evpzPvMrNDZ6IJGaTPuSbE7kMORtgrpgqiYydSNStQW5EEm
Gm0o5LVkErpOsP6cPQ3bS46Iq51WYKH7BeGcsX3oWG7LhPnDK0n3XXuU7JNPqNTn
oTjBwtjlM+5QbDMHMMkAmSwbxeoSZMj/vE3eZy1ZiHlebY/ycjQ2ZX3nSefu884f
C0ynXsGCxiAZIaTUcr6QF8s1NPu4+cJ0gbip82whqWcLjqw4Oc53eMdhFIwBLEDo
NpBmyGwtZx1Viqecq1u205k2i0+5aQUU+pvjEWTEs6p91CHMvDwIKBioJAcuRbpR
ST1e17Rg0b39aNgdXwgIN9Z30pDo0fjdnCCQx1mv/O9P798YfeKGbWK6Q+R6pHUU
JVTOexurPb6+W8RW3vRZI+H7j0NYI7Mx6V+sevYtumKK2G/jakdgX+ZiFXjgHQTS
ITAYkbSUzZqugpSvTZyXA7CUpQ43JVyrgkWHfC3LMoDEjLrlNA2gyZ7o5wP+3xXx
PcjY1/6jQHrKC2FWuOlBjhNH6XKaFru3hNW5f4VL2MUqjB6Zwo+hkhVOCiIW7Gb/
V38iFjb/2zCp4aPJvZFuA6dfwHJnSmvy9Y/h4Xg5LTZ8BZ0CfXfvQO8CGWiMBWTh
hvs9PkgD7Ja4tFdhsAdBjLSa/36vg0oHw1havLhjokaajBB1Xn6nzcXbTjekKb+f
VUnFHxskXELo0upZn3Wu52MngYUFSzJFKMMfwOHDmMDypt47PWvX+v77wR6H5RsO
E+zdpSdx3d7LyOHeq119opIO4/V2i6mGqYH90lmM7UuI9VARsV4PffyG6bL99Y2k
pbulRMzWKkHMFtwE9PhWkhEsyVFIS1+GRW7XrdK8UtIBXDemweoKeDe99q2caeCr
GwlUhEQqH8BEXaqKg7+oP7rR4jPqfevgXxEKFAjzyXgg5me0tY9vJSBqrMdiVB4A
hPbmNhkShKSVMn64nYPA1bMDSJb4XP/7vNwqnRMdhpbNSejx/AP+30tqvg3cWNGP
CcMIbvNGExL8T3Ocm9ANBer4gP98Q0eYwprIFSvhZ/ahjy2dXp38V7Ata6IFpY68
BNFBPwVdNctJ+C5eHC+G5BAvMP9hq7ZF/LhC44rqpHuJ/eNnHg3b7syoPDzNa80d
TG3ovI2NHyEPXXbgwNxahMwHD/uhrX0S0o4e+ZT6gNWQxFK57uj3qbIIJvCHNwaq
ng0Qe1WAKA/jNjjjW4u0BlRLQtlCuFwjzyFdCq7rs2jvfgq4K7b+qG6B30k7Vid8
W2RVwBL24eabNhkeO3PpO6Z6G4QylaRyQ0wHTdlEthCAF+mKXJQWhDxvdhN5Xer/
5O6tBkvwobzmlv46OUU/Prqi+5Obixyob2kBZHnyLju2i+vZf4jAk4cYHRChqW+c
jQREvkCiXKKqfiJ2okiwAmDmXoN3XP1nKha0kuU4j/NTbXFbuReECdSieb5e7UBy
KBsArHWVI80zEgYxaYvjwvwBhGr0RE7bx0IvADEyUTfyD3wk8U0EvN067NpPM3HQ
zt/MYbDTSv+LlOa7vmuSb2a19LCaM0aNl9a7C4XKMIZlHsWvKet1+RjtYRSQKRAo
GKx/CVWJVUe00gaufzJRRO8o1Ucgr48H2GLlAFoP22669jN5QelDZrAwob3mtS/K
fTVCzYPuZ5J8mjZ1Fh8k66fzu/UCQBtJyrroIO+ONO4bbsih4Ca9GrLmk7qwWY5s
yOhXIMV8RrxmWPxO3DPvAjMz3EMPwpXy0kcIuk2UinhO9fGheigcL9UUPwfLxUFP
o2JWBV5zYmDpxIbBP7zR7LGZClYVadRKqNQJ+MbkRoJfCvkknGqgKUIaiikRJYRj
OgTpL3ivKtWEZw2zJ8NHdDqt262fhljr3DVmWHS0V6wPYTwn8INack/0Q4InbMYf
WjBGHaQYaZP4TgaAW1xti9Bf7c/q34khb85eKkQC+/LMyCmr7XAOiGMRuMJySl0j
qt/DrkzgZDThWKwhJcsVvzhorH/ll8jrQLr16rtKK1XazZ1JxhRR7u5B+qD5qOhj
eXpGcTbSqovIsV/Iz/VkXT0jQiCIolWSAMIDwuUxEGzDs0gLd2w/whkqjzelnysg
K3EEu9sQEhteKFMYw0g/XzozEe+XG72kVAQqdv/YO2C0NeXs93e/DGvwXnScPdyX
4rZCFklPG1v9rHmAbVXwWlCtSFm+FbpO/GIIYFmaHep3ajFf7pQ3Ywq2743UkmP8
SA0nGajRiTvtdDsxTcqHZd+O8K3ZyhzbiccDBO/gg5NjtmoEBeJGtVkcV5XF+xy+
erjFH9QCJEt6KV96CurlZafB2g7xT/rATo+S1Z5TpLQ4i8AQH4nJeiPIz1T1nzGn
zYe3fBg2e84d/8uQQjRSQ/W+rHJyFvyLmIbmw1K2qApp4Re4q7lwER5P6DM3GsT3
MuikdT+Z6+uDLa3TZZKIFgLC/PLCKMW0PpKfQQnWgcvQJu+BrT2oPAm6W+NK6EPm
JiFUKN2+0SSzL5j4bhaNQWxcA4kR7F51J+uAJ4TZRYAGg+A28GHk1oAt0N5m+l/r
yMl1zi6RjqvLPaCd+6Je7xfGckVNqhTyzCQSLi4cDTQrPQZFZYIFWa8H1XSWt82f
cAmVXTSAZ/SW0mzCuiBWF5iOEIoUy8wqJ2O01XqGxyAs39hkgtBdZq63FLvItFQi
EtG9GK4OWTazIKEnhmsQjTBhe6YBw0eAy94d6ZA6mp/etdeRcgkWrELnB9114phy
8cR/Dxbi81yOrDkbyrQaDdVSjIdoHA3i88vRs4vDQOe3N+8Dg3/Hvm6aSnevh48K
9yv5/dI1VjBsH527nDkc4m6qag/BCccFQCmtCXH66f3qBL9luXYAFoKQPWL8Bp2m
Q+GCGWK5bIuh3cZtBTSEZPKF4c8hx4eduYUMdbKsv/nkrDzyUA7MdDcpDXA8efx0
819PoxibI3GYtVt7SrXZKPuxa0aSv7Lw0LNJuEFhQbMGrTSirm3kzTYoRvzLGsgR
K//HhXdnEjGGlh6A/rYa6N/m0JcFiG9tcFQsGW1hjSb0QdYsxGUzPOr0SkdWCdgG
GJMKltJuck6E+Igs42hSh2u4tIr2TvolR4W3wZ0UBkWe0Dsgr1fxSL0L+IHxWrVu
SKwanS52upj8IvU9MGFtNLkgwtSAmqmcfuLhmBJi798jDCQVtWrWEvEDAuugInsu
FfjG/ccGGZi2qy0qcRVXnZ6qGJ7chfRZR0bEMwlcaslw3pE6ARFru/srKr1PmnBL
tI9QuvQwq2AfPXFIaSmdTHdc4od/6vZ7fU0ClKsMgVbVb6tWAwxNmAB5N49KS+gb
LITCVzhxoODjrRwbwH0PTCBaCoxnmLRihG5vtN6cfpbmdwQNbbbuaFbKKkp3eeNf
5ZHFL4y6m5HUd0z3Jv4udYVKsKEBYAhkHb/PvtmI+YbpXjqWUJH7u6u7GaFAagvZ
tMSLsnAdr9D4LXHsvgy3GZMmzLzMVez1wwrGwBTwyQSNXwUchyPX4DN2u+szeFnr
+I4V1Hr8ZXB/EAklzq3ibR5c6X3hE1xQPXLF5XEuOJXW0/a4Hw0u41Txs3jB+aTj
bBzGsmr/1fviJ6FnQwiyqqJDhjAXcigrnQliJFipUdrsfkkyqCiCA/7SKp9ay4n3
IsQWIza7upfsqDc9ewzUTeC5JSNTdpSYhFQjllyM1U7cKEN0ZZn2KSqkePt7lf3+
3peVnJeSicTKSCgKgI5YahK1MyrM0ZQoAbfuWZPvTEo3ijVcFBDJoJah29Fa5pdv
rewYbzBwWdBCgrSj2+TNg2DOiVpowwTbnz+YXhXPk6ELB8VrwNPhBjCmCADxZ9q0
RNJ3iHE6QJCmGd/RFYsJ/6qN5HSqoODVrfUXtzDffNh4TgZfKhfoBKzNSv2u2IUY
RmKBb0gb+K721Sb8PCWeJMsWyHd78Il1oEGuV0Y8q8WALPMStzIoQyP3Gh+qHz/H
1EMElaiDC4lKEQ0zIo8PZFmNorKoujT7i53chBqM4GnGxS2a9kX+KbskPQby7D5K
CElRuN37zY7h7BfT3WVKXZuJBhmK6sgXJzQJOAhBC4MiVeqV3k6418JJK0lEKk1L
7uxK81zQUe5VspVwQdDM7RrW5dz4IJTQ2SlC7UKxuL5Ysd8Rs4W/jesqsrDRmnrA
Q9MrMaamG7z+dkVY8w8r21IK/Y6yyv8pYYpKuz1helSTAM4zEsqbcpcQQjyTRAET
kR0czOUUiR5fC3dVxR5vyo8LGB656YF22J6eHdzGlHID65kcD01qlXNZps7KOnbH
yPS6o19Nny1TFRSlbUzxmoQojTBGzWwfOnLL9Q0RZatGmyIeExHtTMMd96LCcBun
DmiTnvWEpw8IFwO63flv1ivLoJTmLuJeKr9qPAX4upoIEYjcKHxgGnpxvTYhS+uY
XYK5/L06VMSRn5aL6YOHQmRsncRNcJ7zXmX0B9YDk8mGlpTjJDOnLztPgkrcqvnq
7dHHknV6N2tIbO8lnlASoWcLNjB+S/+AzvIqPB3V/J1HMbu2ZuVEU6gTBf1t3Ww3
r6YqOr+MST4pNVGddNnspfL+WaxuOyIRzJb6TY8qXL6uGK14FFGKihDdQn3fcjgj
auyWvbcSBuakZ30b528UfSuCFVG0J3kWzgsAEfLyjtZJ/zVPjYcsXJZszzy3Ok9A
Sz9qKZZLfR/qqn431MdB78Xe4MY6gquLA7Grcs/ZAaMrtNimIXRVNvsM93P9yUC7
W4taoZABvOj/sDg3ssu99xgL8BjDmr0nXtvsNYxSpnkPKhT6kCw/sokSykaWM6Ux
h39owY+e9FK7TzaOTUFHewSorEWogzhouQ804hPSoM2Uzoa1ldvOlslKZZNpc2N+
yK7qZ72f/8hv+6ge1mEChiIKYTETT5u/N2jN+1dV+fsvBaqZQTqX+3emZV+c91jk
a+rJIHW6ycLGF+YBdgJT2+HNH8WjSQumZZO+d1us20hd7iohx+96z+b9thzJUc0D
6Zd6N09VT2gGzEDwjQaFoW4diqJu2oHffxw6N1j6RHigoHReqi7PPFYTEtiE5pM2
O0Jsd8qiL4r4/oLm36nJOvbkaoppRvkJgFYs+epdt+28Pk0JMfRmexsZCIXCVO/8
Nd9EnU1ywUCNOF9w/mHQ4fQrYRKcTvKuA8FTaz5id6mcKlQCX5dLFpWnv6QXyB8S
r7BemSx0EpDsrx5LehCIyjGj4/+nuGrtoRD4FsEP+pU+0ce1LJ/f4992OFsAV2zl
AJrKR8/MbJ0lhMWyDCY2vv05ZUinKyMCIRlxbbYo2OBnvK6tmHhcQKuHZ7kLZF93
d/FmVdFg5kzU8ibWI9x5ZFrcD1Je7XRO4E/u7heOk8zTK3aQGeA+HRelOVhVY6kn
cuGmoABZcrAEfqfT4Ykrc59/aLjkUnG0kx7UNmJGYLLW/a/k5jnpyMZAeOc9rcG7
4+gdjyKx1JxK6z1gTNfuz1yd3uZV8fsG11z0pH4RU7as+7+DeJW60Jb3S5hwkAJe
R7ul5Bo6U9E+Hgbmu7nHh6fb+gL8gRpqk36r6Lrm6k+RTb0zn+eLPiepuOJJmGGd
fQKsjoN6SOUYIwu2UJIx2I0jBJR61Qr7EopqeCTUkqHwEFiecWnwdpt6L0N3ufqb
qp2uzu07Z44Iw6bln//ILcjNpVi+a27IQCMoW0yvDkP1P9coP48ON4fQ35JxJ+gZ
Y8sjXYBIH2qXlPxrE4LnyAaJJj8J4xM9Tdhe5lTfbABf4kLB5Qdp+C4brhYyo+8O
0zgc2uknUUDHN9P3f4SZocSHUCQdTddIA/NLNPc1PY5wHHj5+D71pHWeiCGzxuu3
d2NW9e5uEeh802GW0jiC8D8fZ/HXNvv6N4lDOofOrmPS/ASxxFjsHF/Kd3zezUqp
/5cLn7orzkJIVrzjkRdKBIo9YhxOUsuQCCqIXBlbt8V1+f/TexbDhJ7eQaviDE/E
ZcMWuP4rx6eN01VjYHZVR4hjbeMOoTwtIzus/+GLP0bHjR7zokCO5H31CsfM14mQ
mka6rXTisFfW5VkTyKib/lRFwxfgBnH+VU2IvDiA1/H68eK9EJ7EW+Gd7Lp+KyX/
tJ1R/VVsG/FtQRfjSKKH+LtPF+PQeb7x8ZEHY0JFpBYrnRk6WR9fKgxER+x/vUPu
bG8HzTepSKlt9JKFve+jvYLdS43Gg8b0/kzR45Nmf9lTTJIkDiOTIaWEfxLa2QKh
5PtOSypbeCO5+tXEP7t/Ikx+4L8kisWC76RCyHtfue/lflxxSPWdUcFvA+2JEILt
L+b68DNm/li1k/nR28+ejwpyjEyDcfBIq5xEmG1mBDPmVIV3X4DITJzWDfNPRPSr
09x+cYvmmAx1Rkg7OSxRoWHspf+XAB8qPWYSHNNLQaKTdJIYP0o+Pd2nLioJkb4N
8tL55Hio7PP52URLdLfwhctHlob1Cfzz/bURO6T2lwfWmRZpRjX13fjPKLGxwl71
Qigb8r3xrkp6VaCtq+LsgnO+w054aeNXDL9/62dXSfxBimpX6qNS3U8r/ZDmzoZz
cLWedB1BO0Ltwb8dyh683pVc16M0zuTHA61AZWfkQpcYkGkQwPnE7uLyuHF+3N6A
cfoTloGLZy6MLiveRyN+9eIOYrh0NL4wrP5TGwuZ8xbYUQ3II1clbVVUPIxunlXU
MZqzP3dQfzCO2G03HkWgN0fJGnPOYDtylecGg27bwiqAZXpAlnZlubSdW8qYGYZH
dncI/IBCSXUKRTbwWDFeaP9wB6fn7MaJjTy0FJkK3Ie3ObCzxG8FDKLtsE4AigpE
GzLBXUZrLO1s/7FEor6E+wRUqL0cPN7LyYZZoLY5Sk4z3cr2fZhFV1QF2DIogkzu
v/Xa+PLq5MrTed1HYKC3f/hMPB0vOtdNdwZTIz80AfdTdycdx5o3CNIN7xWC99Yc
F1o5d8TEeA4rfmkSFcftVKWvrMee/6f00SxIEgXURoT7/+gLAH4QNhOK4xUAze1C
Dpgk2HtkoEl5w0/+Q7Zc6D7kGkinxcWSgc6/XGIFYrBmb6ACubksW5Vuuu1OEJhO
VkYdl1eoCKl9hFYGqRIZ3UrrMl9E+k5VwYC5/lhS+FANrD0zBVQViL8FXN7mtoV0
902Tgr0Hj3ZGj+o+ilOTcMr9HXrXMkVxN+Q6DhBV6vCRZtq4H1vQAEEQ18YF6CFe
Uy1gt4w8wtRyrB1QnptVOXv4kgMUpCthCIZbsYvZWH386q4zndE1YIdCNWbitcfu
yGhsIEtR/F2/WuoKxVuwuH7zymPYT0LCJM1ELxFtCi3kGTQ34OBQd7uClJzBw/pg
FKD9CsdgdMV2om1WcMIFECPW8QKEew9V9m7Oh/WEiUT/nZbvoCQ3PgR+nszbEvSN
twrud0h6f0Gp98STG0ed4eIsKc5XMIcr5JLlvmtPTDnmCOL5h8Coe661bLuXOwzV
w/REnvdYE8eOXcZN0FyTnmEusR6sGFVy7pcTFk2hXUSxhQKTv91RQ3hVacrGwDTp
63gAIIA74ToxuU/4jQz0NVZO+jpJFAofLMsJlE1cizdeZzIE2ipKH+yo1bdiiNIh
hhukW0uzKc9MANMpIHV68xkgmLZBhBoUQkBr4j9YJBfHIGVaj0/Tg1alVmvBDXHD
EhMmikAJtwJ9g2s6t1uEXfrdhJAhIca22ITPrffVuOkIuUb3VxXnWuEdw/ig9oK1
uhMznubQYJ7KD1YMLXcP57tYUWxMoq1eAKvN/9wVZV78vyzhTVkcq3X1oChHHl2I
jDoPbZWjrk+OUL4HuNlOfl6A1/Thp8mwc4aPmO/2hucE+ybyBLZXVtdaNZpEBgcX
A3M3UuGaymyxHyO5mEhan9Rj55z+UFpEA1WEyZJ99SxudvscBObasHbHjv8GwWZw
Fd7qfYCWh+ODMtSz+l6zyuJf0B/987nxyhfPMNeP0tc3y/Gm2hJaqwj0Sft/+h8B
zAVLVa3MUL/JLvi2752NuUR3/cjmGczTRjDcPVdZTQcR+gVP/iR52bPxTxcYRHa5
44h+qRdSa2ekGUTgyCxrS2ioAZHdIbc7zcpsP/GV6fieOiKa806onOu39oOjfZ2X
GkALukqxISbbr1qfhKv+CdI1+APJcvsBdvRC3qEWZ/DveVq8W2nyEAFTkhrH5XMm
h1CJ34BpDvzQNz0l5WM27iK2c83zP9p1ImaHCUJwNOOUQqW4PrfSFbF1iE1oiuEr
Pcs636aNEKqjo6zOIqbztZdYghx7RjycVY6Lucj+teRUrq6iqCIUf4e9Q6el8CCF
YQGF6WFRWUeykuJ2KeLUoGXDbBpnx1K3RbAlvBroJySqJaGBrkaYhuB33bLBSv+W
SRR9CD50kDwEXsH1pNp4MO27xnWVfVJMCRY9LVEEB2TVpOD+7DzI24E3syRTsmUb
OqpgA6YvFnKf2O238iMLAmRIlzls+FaUF9keqaiJNz5JB9RsTRKy4f++yqRdLaK2
fzzxxsPeK/6rvKCf3xmAWUDcRzchWUwJTqix6Gb8EthaTHWvuJr+n/IBNrY2W8tN
j7QogBbYUZvOJK0XnEaVkptA/fQVlcg3Ux3rcEYNrH7R1Pi0HpDwZJ4WzjKGFp3Z
5PTgd4pthfL7Pcg0EL1jGyJTLxIJzhotV9qhxoLoeHUW1vwB1YqEjvtrRZx6hoFF
Dt41pm4mAEPQg/EEnFoX15oeQLEItiWhpRB9iAaBegn9zCVgisl1tBqLkXUOJev4
g15hx7AAHKNDjiwtgglZE02BXKW67BJ6ZvTlqo9/rRubaV7DhrqX7Z99OXoO8WgU
W4C+OM9eqgff8ZbA2/UWg+ai72wDw5yauirSl3cjZC4tYbDy9jE6HYdbONMzZkzz
ji9iQjgylnPw0IOo65Yhd67CHcEZGOr08IQKD3cCzrztI3Y28aS79c1KVF0v7zvV
vzMYpb4aXvvmC1nvEgjJWJiY1QDnksD+qnIrmMN9PGQOEvyAIQDr8u0AMp0D4da1
oZ4eqQQ+CiotUjTXtiqjRxDaVyxlYF8xiVb1VwYHfd3720mngyUFLtoHqHcOlZ9D
gUnavPaG4wN+0ULidXoBqf9i7hUw/9OgZaTMXQSzk9W7c1FX3PHOWbat0Opbps7O
ZiBgygg6kvIykFfxMyrE8gcjuO2iaF1RPvdwZ5fyYcH76DCtT9LXN7sy+a15U/ca
79hMatd+uWeIP1J7nxuJLJcvwrT1C3OjxMZz8SzI8lns40xXFrvnp3BC5TLNM2v3
UejqJEIhFBGCyiSkLFbYYzcq768nYs554/ajI4N2h5tyGabpg2HUYgylCTWYK4ZG
b8o6RCbVSXgZzE7noTlC1m6q9p18JYdjQwP+EGXJmsWUm4lnkv+l8GanZPjwNVhV
CyVc8J9GyCzkil8D6e8eZHPgJUUXMvqGYcYOj2OzoAgKnXkEvj8X1UR9QLr9+CRL
dWbteJd6ORZY1t4AoTMtBWFY2M76ezdJ63bDvJgfHAdbpeuBVShsKNTKlukYC46a
ruyKNLKTwdrbiXwqQkkuiQKMkb1S7dm4EICgNBVugA7RaciOyXFB5H+v1EKtk2tW
026Lsk95KEwu2SvWKTH/rpYq9ZW+bdriwllTQs4lBPnf4PcUuhicF7LQjI1yjxCi
EEl3IFuVGyy3RGrLFDu+Q7wmex5CSksB2RKwSP4Wg68/XOke0AkrUPzEGFZ/fSt4
IsrcV8R+2v+j2fOrL43pLi/FDdgRaVppLGYGEYtfX+lnjTE4mg2kopL4wjRteNgf
o5aQtUtFn8Ia3Z0GfKN+2/UdZSC7I+/kNb5glwM1xlLnWktN5dp5RXc+KvtHDLsx
TolEivpIS29UnnTfv0fez9J0zAMGkPEj2bMoDT3KQyIeHj0Gf3xXXo8LwIku3uLS
tPzkzAhqYQJ4TTMMK0ao5Q3e6WiqfZMtpM9pWqifchakU1Mgia1fbh5wGbhmZ1p7
5RJv8CK7gAWdE955/V9mSv16JBBiBGIrmDLBSB0FMDB9llx73+fMcIwLhXLbQpUg
DZL88ETmmHlvfXzyoq4V9R1YijhDkhunI0p+WLzEm51TBgluZ6lI/j+6z1gmTIeM
dvBMRHRb8oZPyQkPUd0HW00GfEAm9D485M5ZpTCkHRLJvLzmwMG+gMFM3CmKbc72
K3cAHfrZCriwSBUp5r4Fh3cMFm4aLgMZc2MnSG5iHgBUF64oYhi4WO2hBiX3jyq0
cQ8Q5GtMtbl3JUcEo+c6EU12h1IkD+xeI6+5cNBxH2VQrYUTPf75kIsnfYYdwUfh
RFc/X5qXD8ow3nJJa0fwXOCzTyHaPGOSZAU51BAeHpd3G4QvxEZYdnORJnXRqjiO
1FGGpfLuPjdsiIIomyUWVhH6LmGySFTwL78pQ8YVSjvGExP3zzHEVB6lGQeOPn2b
9W+Dnneb1rHXcD/taooEH8DUKyGKgVN+DtKaPLLnpdQA96lvC4dgTcos/CC28bnr
jXuFbiCePoEthdwlioN/L4HqW9O4bUs+6jC1kaP+WO87wiLkCbFvKqI7jXtpKNcv
L21iyBtC8AIbOitESclygqE0sMg55YdWugNiOJFVcVWS+esZvylZrJhNYOrMMnj6
Xt2hDr2aFcofgq62OadPCKrboA3yE2tHxgQYepYFG4TjJyIj3uL7hEuybUvkPJT3
SpiR9ztCd0r1t+zuHnUjbC3xmY9fs2WFYe7oZ4Pk3S/pZr/dzxlkJNq/1wutHIYd
u9mLRTaX1zo4ihNft/l7rFnaILz8X7Y21HL2Vt5f1mZx5nusGsFGNnrXZoF9+zMG
ZOBPIjOchzv08qRrMHEYHBeC+Sxlo9tNI8dB3JK2HOKFjSoJyJRqxYHFRm9KaU7s
/ZBRNg8erejmfW6lri8C8+1fO8MiSMRPnZh5OjijY871bbQdYdFPwY5fRIE/nUi/
53H8dB9nwI4F+oFiQ6nPoonK8bhl0iav2cbzVgjBfz6HunZi/dW9vx+mRu1CvclO
QXK5JUB/9qs0ymjHO12hUyQrzPm04RqsBAcfNIvr4lvEXinKDsW4YMUZ9bIDD4aX
vgLf/hK3UPo5EGwyoYEa6omGB0L+rR3RcHdGW1N/DVEtpeMCjgjDrCsPhukUyv8g
+xIr3O9NsquPn6aAjN+n6B3X4eG+6PTFeqM8ww0rsfbSyPwN6OMYQwciEanMDkzW
2Qvy51bgOpPorureH6aUa7z7LkaoxMaHn75/UFRGraDV+CsH2V29At1ojctTuiFv
GQ9/NDOA132eJ15wBAP7DfGVojmlg/AMkPgJoQYjPzrN0fy20UPK/E5hR6Kq0WU+
tc3jgAVnqhc+IUMaiaf1P9ducbp9EMpWpY4V8Ovho48HOmzUpBFlAMZ5M3Dxv17R
8IXM+iQeshipQhNmkv94TN6nbAukFBsMOpXWXCsHIv/cKRbjpt1H7Iw9dWKzMXWg
ly+09NIvudEN8vibxaQ8RhYOO/xY6CvhUdpyHOZppqqFNwI/tnZBMoSFzXv6F/o/
ODXhJJUSSxVGCf1tK5g+Kj2YfXRO855q8yoR/Or6i+t8tDG8i9t6hGtwLj+LKRob
7elwSP1stn25yfjnHHSl+h4btpgqWb/+BL6MgwmuzjbfxrATdTNdDWtkdyibBKJ0
clXfkVzevQMZPl6/YKZch97kV715FaQFydh4cO5UZj2uKhvuyJDTRNBVhkVZjSos
0LLqe3z3YOsWohHmh8XIDYaP1m9BqGCIBhY8btQ4VGFgiNIS/siDNAsyY9kakRI8
cKAJVbZDXz36enWydcdgLNDaP8Yk5mJp6c8dn7agSeJogJYdUg9g4lnWMUyENwf/
T7FGredPLZrMalOuGtqeQvmQPrjIDl+QN2UJ3K56UqvqkxqpyyqgKHvkcnrKFvFh
c8V8T4ZfhuRvg9C34+1LSpBnJ7PEDZcf8r08HHfKHkhWD2cnu7s62ZLrwWojOLYM
uLAO1EhRrdhxa1O3XNJO1KL8X5XemESNg0sJSgykzotnqAjXWw3C5e8SPoUEbC9J
8ky+1H+D/3Zx9dhrSXG7IbxkSqw2E93ua4eqpSttuBG+QSb5FE2RChsRqqRkNgYw
R0LP3CKM8+zHOkoo2cEiWogS7BmoU4jSWwszPhoLeBIgfZOHh8FbGs01GBS69J+u
n7K8u1kotBBZbpdGfgw7IkyFVtmnF3Rcxwb3arAJV4I/gbcuWsayEvOvIwtgAxfY
I6/vRFwR2UvkZR8/PZrL87VIC9anAP2z86wRvO4QpIFUVXe7kArd3ukP9GeYKfUB
+FdbRzWq67FjLpTcgFzQTt23uT1POiX2Gx8ggPWmOhdUxG0S8/NDn7IJCqnZscwt
2qjQsIMgkK1F01sc1fohr6dWA2kSht/DXdfGnxThOlCqeYPAGvL1fSb/AF079Y/k
Y5D+Yh2iSDzHslOcnsUIlu+qbVFUxriPphHPElsdIAqt6E6UtXJNBJlBHcO7ibyp
JrlLjD0/R1210wEPEZN8NGlX7HW45x2e3fa7Rzy/oRk5DnTHMnmfZNo/7aoaXHbl
pfLRpJrTzCpKr2/MK/10akhojstpzKJG8tSLxxuGO/jWxImbch0fMkUYRXocEQkF
QKZcTc60F/AamklZZUtMiE5FokOdh5l2lXs1DTlM3iocp1HgGdMX9LGEUz9PtY02
xrDvd9hd1HqWt5URdawo4Ch/auy3bCTQDIGMvHO/684ORcZsfMmZpLFzyuPi0daA
P/8Ad633+ZhtBtgRg1+4JT29oAeA8WPdj5wFSIKolM42F2IK6vD6eS6fWokjwoVv
b3giwpmGYQBfowWiKx05o4poBzIyxwlRWb+g80YbIeLGD/81IgAeoE7JrJ5QxQg3
h0hcMLEy3IsyrldMYrmuih4DTUrLn8+FasG5VtV1dncWEDbIVrdwHsF7C/kjG5m+
WRWICjzo3Pha8b1UHcBnwhFKX32w8QGs2az/FJlcNMMIY72a3OaJIn/PBqP+7mDq
lVKUy9ElOCMvQYSgUxzqD2iBRXETwoa+Oo5F0bXjz0RCXeeljAHAq6iHRQ4Muyzq
h+NFkGpbpWTIwDzSjjsFQXeKhW7W5cNFFeoZ17v0NQvTaBr9FTT1Z8PjMX4Nr7Pw
eZZ58wx1PWodFSlSk9bztMifMcFG0FswYWX05Q7wHaitvffq05PgjKerUwzyOGNl
M6JRIHxIHUc9QBjAg3wM2uT9dsso45In4hRCzrTU3Y6QQv1FIxrrJ0DbdlgTl3DN
CCAXo5Fwl82ZBUQML4Ad0LA7YiH8ONfEbyig2ILujuUiKFlk92LTZsCleH7eWmNv
15vTP4cHIHWYCfpLE4MNFK2JVWszmM+GBsKF0SmmFxn0LhW0JaQw7T/uPldeldii
iw9BYvTOcK+EeaT26b2y6fjIMG87nXRY4IulaCEJrs9xcB3POm0AJ3hgW7bC9Y6U
lHsEf/VFwXPfPm4TakRAn2qXF/TrjPctnShH2P7HkO9HwOnUsXvG4cpGoCi37E9f
0i7w80sN72QNBJz+4uX6No2cVurozgbO0t4tUNgbemaeZPuVc6rOPz/tU1VcYEul
BEqVlTqNXJX/tRDNazHxBd8tIFOKTm5WFJt7MbQ4NNsh2R3K7UzyF3S4C6uDcg4x
vSvn8xaWM5WvnE9AVYqLpZ0C1SKKlV+sSlNVBKSsWh8QViaBP9Hej4AwsRNTX2IT
aSbsyXveafcmVOklQE6XtaaykZApAx3vfqcg2YyaUUu/zyT6gTPZVogi8a/Zui8I
v+fZ+ScIrj16TarDNxATkJSDz30BLlw6qyp7kZFqoT3Ecf1N5RQwF0igA3FLwPDr
28Sr4q1plCD76ETIduL2x7ziE7zra69OSqUo8LHeFdHzmX9xtEkRPvRlTQtzaitI
ySYr7wknX1orUXX7z33LkSRgn2pooGz/+MSZwuuIUwpZogDEaM3+zMcPz5zwSFyr
jaz3yleevMNcnREp1Bdxj+IlhPBZDqo9pE9y0/lORn2c1HyqyloHXkcKmL468kIT
1FuPsyACPwSL54koJpibiQANkFdzHaUaMHnC0LOsab4l1mPA1f5XEbOBvnMGcBAf
AzQtDg7Up62iBn4dfyJxpJ/ohEzSDkgT0w4T4drLw9dG1V8lQvLyvpiXdsbYTDam
kYxwKGm4mXXI0rVBxvyovp5/He0WLq4Taew9UEugWWm9dJSKZF0S3W1twyEPMltk
j3S/OZ88GjdOkm/BHCQNJ9n1ZbEblK31etLM5+as9qWS72z+opK6dDDi0Lqml2dW
Axdf+RdkmMREELuOPjRF6CxVzCI1pCsR7LWE2hNoBt8+mHGJa/aVGWU0YHPuYZz3
yciY7FlP24WlLzWt78HqqOIA9VVWGaEkqDgAhWaeDZtlin61CVuKC0BH3ovaVwib
ZdwEyZD+yRm9zJVh2rLIueOKLqEQrKNAx9XY3gjAD/aschzxUrQ6Q0QKKcu/irhn
f69L+C+oEff8CKrCtaZAD9y1XixQ4O1191dgy57EkQdd9tKR2Z5RR7zfUmFTi5Xi
GtJ61dpcpDrn8eeA3kO6A2dypw6gFT0bxSsGsWY2QP9b/c8oMmYLPznEFmxSlW9c
5+sgjsiDbroA/A33ODWVhT5O9XtOYKOP3Zy3EmbBYD72MZdvVwIPefv/xv7EGB51
IdFXh2fapn/ralMycn5JwTS0Z836b/YbZW13EI84WXnaawUV4LT9MUbToRHudwvt
vX297T9HD+ivlqLFKWOgizb3BvSOKOkbtr0tElE7Aily4geijMchCOjzjT4MbQZC
aLsX8LZ739IecLkBXxVBiPp4KZsBvDaQDCXUEVALQ5oJrJotL7431DP4CKVcb64k
AZu2++/3TK6HmsKbpFouSJDMG+rADZDBxgqHL6Gd+E4SJz23xeWtnVOL/5VOpEGF
QTMoqIE70LSJoazCvFx5G9A40yR6c9E/3GtuDuJzjY14qvxEjELx9M9spm1+S/Nx
GHKBi9Y+HX7RBWGYnP+1R5Xmb7DuzJ8S5NEo5nd0xxjElF7XGiG1ubyp/ufDIhsg
DmN58lB5G9Kds6NrTmlf0JBDg9fkN1gvnt4zxahGdXVKmkyXiR+m9W7PhtIgJKkt
xpHB/M9PUU4D8omWft2AFjAxExDq6QeYpYRK5Y100I6kkXe7Na+se+VRALNL0+c4
d7Z4DChREc8j0UEjcuuswf+Q29t2rAQ527jmOyRWUyxl1c9xcx77KVWEi0U2vgT6
67+3zC7WMG1hmi/bfknmV1OuRXfGZpvN6n+nkzg7EFOdIdKKidUSMP14lgXvOOGb
OMkaMfCm7m3ehzsPxK9w67cNthf8n9Bv88gldhrpO0EbLCqYsqjH6+uRjjguVdGV
fPCFLMw1vnl7KonG65v5TFXOSa29JHhVkYuvAFJ2+CTvzoEL/x/AtRrxIgB0lZUI
wsZRZanqQYAv8uI+de8yloN4NLE/j3HFngcJ/UQJi0TrktpON2Zb3gNcYX17izox
GZMs/NywQVT81gTuF2SxpeTdrapusprnDBXAPaIYIHi3uwdnRZqo3fOzkTQk/hKD
YTV/BjVNCEOIH0J2nuYj/iFOa53wH0uYAWNFe/i0WcCbBSfWKFLxU5FHxqD/iiEX
vP3wHufkBXR6OFDMWOUGkGuYdyHazJlJYcFJXbULc2zGADO9x49VR2/WqgE8Md8S
iwdz8Z8cE6KRZ+iReV1NFTm/PX6FZvBhrhQGIdN+4u8G6HBoT21lzVWRHfXPF54J
lSIZSKW7QMXFjKRkw2WrQ4rpG4Hb5LU+UF88RlwwoRXX3ZJ+tUqfTJz2/87IKZQB
ADlhbuGEeLBX/K7A+KLVTcFWJZxeaXfBlz54pzt8vDtnOk/o/bCBSWxhJOaIeqA8
5ie2owQIZN14TFVSUz58JPokdhFGUhsF++in7VKf3WEV1S8VNUBvOa7ZnL1yLVx3
Vf5h+6IHSWDUNcAWQj7LH3ikTAJwl8iYn06Q9BiXMe3NQKjO6kbeVIJUSGoYh2PC
GiAFOaBc1N/KQOGmH228KG69K12MU1ikNUYXDpsjfjKdtMmqSj07D4O2XMnkdG3n
6eTXON4jSbnk7AIPIxdH2p1/Si0dNwSHqKaRlLyB4/UW56zHdLE0jq+ps7/lkyjc
3fee0WLEvIi2D06AkoRKVTr1x0JptyCuK9OQ9ngXux4qKq8qH5+XqpF+dSf6quGM
t0aKuR43FS5yQVod0tXDYIFCGI6XQq7NOYRgPVyxpB7Zix0JmrEM2KwMR0YhYFF3
ulpyMa2jckhMjfSjcJWQ1JPs7cxbLaKDDspowEqXKRQ741PDqjQU4Sm2BEmpZ+Vn
/as2WEhALIahNxb7shNU3nSl0nxEUZtKA1JNbVLsNGiLggV2nKfB0JseuBjsHRWp
lrzzQtHYyAHjEyDlr8FQqCEkR/94uQWlVjy99Cdqg4j6YuDwKAa3V8EK6oqtADq/
8JQbAGBpMWEj1J1Egl6UWbWY0WusIal5ixoL+i4++0AjBREt2wTvSQ3dJNaNAezs
vMwqZMQrg5/Jg46twcftJ5RUgAOY0XxUZBiBUPJr0P9gb7bN9vJlRcCM6gYVo5HJ
O6zBI/nbgiO+jd5yulThfz8AzjRDZA3tlV3x50vYrAYcksCGEW/g/lR2t0MXxowq
v9w2yorMiK3GzVVm3G0YcI4MfRtEutZlhof2fQe8xj7+04u+qLMx4zvu9JnJwmN/
OfxIHR4/J9H8YD1sF+7dmugs8vol9o9hry/ScSbGw0ZlgmHV6WR5EHJS01LpwMk8
AVRsmwKtzIxx4PTQjtLP9TnYm14hZHYL9UrkalTw/Oufpk2LL0FeEdW3JzSrwgI9
XkguBRh3fP7W1BoegXU+IOug3miL+dTt+fHJtJknKyH0LZpId6PJO1DKZ356Ujrt
D5MMXVz5qTcAss0vWLO6I7h8TWFEq5YzVvG+tRSAMOZOqUyaktcYoRw7tSHUTpij
R2mtyxMveY8v7eVzJpF+/ZCaddeH2n37f4nceXhLwCZDiB7n/+bAXlENlec/zzas
RjtVYWCpfHRBc/o/lKcbnKe1WmDuzeWaa1cVYIgYQBiY4r+LpE6eg7qhsdjwgwaU
dKR4GN6uHSw074JUZKrGt/9HFt+4b4NikmEAUODXgsAaXWS5zPhCo2+wlXHSn12e
ca+CFCpUe5M+n1fk9WP599EIi6NfX0eV4wn3Q9PsSOoLYssQDfgKAI/rB7dUusx+
MJCb8+jtW74NYci5UxiRYiUY0Vh8/MAS2Aur01Ry9t5bpRgohB1W5ReSevyMVUFL
NnV0aAjAS71HgulCTc0jpApefrhunAxFmIl0m+8r08VdiC5SFQ4socXOWbjlHC86
5RBMrkcF9ar4ncr8z5maOsT/42NqadE60H+CDETeKG0BujBRKWnNgDPGP0BrawL/
6Fh769wh0fSflxRRhusUd47CEEPFFB08EH8rJSVM0OKF46CHFZ2GotyNckPA+4gN
WP438pNXH8v++PtmmQXnfLgI6aFgjV9rJmyw4spuOtoKnMCApzYqrW1LN5ibU2QN
7K8RWyJS5EP/15YkufWZrZB1yQuF6UWhvuFFsnpc3xyaGrbCrYZz2fgIvdZ9/rvq
sqtHeqx9iVwLEWbf8ijfIRsYqkFGKve4OIAz2/0JKVp14VlEC5GQ9ejUfKNK6Yrz
+tEv79iqc41qNLE3Sy2ULcb9cJ3VNes86EEoXzIRT3DnXmN/X+NBShBW34U65rqT
C4bG2OBT1LIY7ka1U4GBEkMXB0Byc24UgIJhNmzxm32176+fP1kvdawnRV0Axgie
NOwMN8LqWKfW+CvhG9bEthWebupU9VQ7XOX79hLg/dIDCJ7qNd0R0P3XW9bzLNPN
xJ8gPILsTF1RYi9LqnSw2OBLarAtAl6olO77bnMgCRpgNcgQ7408uc1/2E/+wNx4
X1w4wHJxMdaCBfZb3xdfjtaMwPwQitrt6X2PN9+Yy6BB/TRx8q2ag0eq8hDYQpVh
h108IzfGfsrGBgjL/c3S183g5OlBOjf6B0ZDHhgNTLCAbIgpHADz9OgTcM+PCAwK
YZ8JGxk6NLnMsrjpvrRnt61VSkKxjjzajsPYZNj9h5RLs9xYFh2qJjrayxFKJvuF
q5eNfRVB1AvENEleJojb8wDOBwhNKvtVlAL51z/gemZKTP1+yMWRUUZK21eR9fz5
97tuQETta+zDeoKz+UkGVaut20Dwf7sTv3YFvqwmExqw1nXt/7TS55NXONcmpSPO
Gxtl+MYacPWqDji+1VTKIT43V4r2qHYhlE848i6C/NrX+fORTcHidx5guNMA0Lr9
4cB0COlZwKAi6QokqEkeZdn09YDaTZgcb0h7ujJKHQ/RtENFoeZHkgmrNTIJ024l
ES4CheQUd6ma10Ms95H98aIrRrbeKQasNRzMzooXNbJEyXhMdjg85yB7cr2+AYyW
T3oHc6+tclr2rhSVFGFc7oSWcb9WX5HqZlYDi7zuakjn8tVrvHSSwNvkDJ4DMC4R
Iy6G/oa65DQUha4Qbxiz/kK4Rh0rgyAM0xcwz41IWdVVwoaMG6Cvp9DMg1FfDmKs
wVjJqhmUL+bd5nyhVZhqCq9Qsnk+bpimLKKaQae8d+78Vr0E4xHoD9b8UWzDZ+Ol
ZK71sBuG4/fGT7l/ASrQErCKE6AQJHwch1smSh2kEGGDVcgRiNmSPIVIxFmdo7A0
w/AAb73+eVr5LlHI8CnyalsafEyDdssfvLTmETGZG6BvrHHLhBmGpBqY5JOoEgmY
RxjfzkraD8UmA+bH/Pb/Ge/kwQ1Xo2Qt2K13RM3KSQ7sjM4iqPQbayWII9QursZb
b4IlqI42kPh8UCs6eo7aXs2ifgWRlEn6lWlZaluS4+W0GtcJtDJ9sj0SDUlmf892
cTO0fzc+TB1tUurPHj7uqiBNypm10oWCN35d2TyLStP3fby4f204iQt28n+oo2Fc
/gfpIfjXuEc48yGztTKZ33OrSOxIkvDaW++GjcSYLYnrUEtDX2smUDgZqppgF4iJ
HOB59svBJG6kywTBn/GRdBC3U5bUpJxptdJ7VpDsW+Anv9fxDAYfC/VPSHhrtkvA
K+BnYVShj5FZ0vuh9UIQFuCwiK2KYzTejERGUqR9fFufdEPeSMrWFIxJ/3Zopwb6
wj/mgsVIC4b/lUXSkq2GX7aU51i4CwJE3ZormNisTZP4YLybvCRScUktmgn7aNN4
rJurtbaV4J90DiEfvaPfHuGR14BZY3O9HOraTzOtLb+dgGNbmC1y4+AXsygnRWIY
iSGogJCes+JXH1i3hoBi+V4iC0srpTSVoO9hqNVeft96c1q2wbrqZPQ1tRCyv60g
/lIGe1hWjXdJUJx3X/kABQ0HPlV0F38qEqQr89Z10Lx/RnEuPcWing5oBpSsUIPZ
25C1nezdq8stMzJZAN254iEfp9AZ9Is1v5z+OOk61G1w4AhKJUoRvZ+GDKJkfkiC
IXEKehXYXuyL/Eg+utpsABBG11pzAbkMdbFpCiB4H90Rd+zIxck5TQXfiKd4zhUy
GaQ7rSwLblpLWt3NCmhbeu0YlskRksST1eLjymCLbYmuIIt8WbOTURfTQs1+GYJz
c/dc/+R7P0p51ylkKMmBXuJWzSWBY3nHj5ced9CxM7mz5+xkWzcOvLgiuEDD1gnN
DLtsfSgBCU263eEMdlLTLHxo1tL2J+k3mydoLVk+G6N/xAsyOijVjKO9paG3LRsP
qbClbvmptjQnmVhAf04L2Eikv6FTaVKcWWevDQoOLgdEiMfF6O32FWY8G/lYt28W
br9Q6pzpI+VBRNwg+khkXJgM6ketptpegiwZDNxd8EmSsIKUAkWYxSlB/prZt6C+
DCSsw+fpEUl3XQl7E1+/tX56Dh4rzzy6vEBXBHiNKqst8F2jRTo/k0DNsjLlj7m5
e+Ya403VjJg7+rnfRtW5bHsKQwZDwBILOoz28bF6i2I/q6+AlG70/a0mNBeEdFzv
BJLpARRJ6W2gVz4khLb2zZ+Bk2xdSmeX5gA5qFtdPypo0gavs69dBXCcO1b77oXR
YZHiiy+p57D7NTqjTgmscmb40xFjjF5wqj2RyDFhaJcUSym3omwcjF166OhT689H
sZ3MBG6dzG39Yf3EBpodBBLO5jR8/B2uqt6fKwktmqSiRlFgWO++sjFUZoGst+4p
hmUpAONROmyA+uxvyKhaVqLGtljlvmN1GUa9PorBoS7lbhuDT+d5eHThPxT9fFHp
8bYz4yqhsecXhoLN6cKoy0jZTILbGbu6s1MQxmHodXO3BXbl8Yu+8ACVEC+dQ5tx
9RpdVr1r5FTWi9+cpOCUuMCsU1Ydx77lPy5Cl7tdEBh4XdX3NaSMnVLT+FnJuHin
IhJA97BZmbUXzRNIHhsAJLOExJrtVE6cUhmwSa9mVoQv9tD6FFyEpp2MBXcRkjK0
4AibTaC9rjlVOTlEtTjCXoNEJUedkxO3a6ss/H/c/DeUSssR56ErSS8lI9L6/Ygh
ekZ8aeWt62Fyv+xBggNyV64EP2lys+SOkl8EWnPOMU0EfXBoBXnM8/IfuhNr7usV
y9w99U93qTUNFKUh0rAK7n8gQuBAWq8mpDRmvtTaq8o5MKRTO0YGAPSOid8URoyz
GKlnaZKCUUDz6blLbVMF2TPA91lfntQfS7c7QHbZWaOjCXuldCkxL8ZR0u52hJCk
MDHzSakpUl/TugH0nlX8Xyfp1eyxfqQ9dNV8T7dFita83Aon1BiSZDN60LtDp8kM
HlMdUI6H9FP0vTCRsdZPbcWI5h0ouCyOOVJaMczYp8qyi29UFdCeYYlRVWwe7A0j
WYXnbPoKOGZ5IDg5bs9QfKy03mTLJyqGZzfizPPf45HbaYgL/1ig8GqqfXuGgZfI
mYZLT8W3v+LoHfBKfRksCZGlwbFHVaqAhZRdaAtdSt0jniu89kAOfXRgyQs4fxA4
24NzMcPqjXFqOOVbWuxwpQd512LxksanlMjx3KmQmw75fYV3Q+oH/1iOPXz6WpY2
KHJ2HpkjdZCHabu3eujs4l7H8impGXSIHCyM+1LROWGa6ZcFkOt5VUGqzyMQfbic
HYYr2C/jD6mKrHf5IHupciy0AYu6/C7yddFMomHIMJl7kFmjyxFEKKyTkWK2l/Tb
/qoliut9ZDu7+uUICd9cD73kDpcCbMpX4nacODqeHHeKkcGlYMeMLkPjrNipeQNz
YNrIKnWjYzX/EFRSLmW19LgU+oacSVjbtbyyoVlsK6ni+TNn2i2uBDOw91HnSTOD
h0FxwvUIADmNnIcI3oQp87HzQnc8od1NlQixHGnRwmeaPQFkVi+l8Vn3rt6hmn0p
pHPQrn9PCuHjcm2kv3tT2iEr0aNFpQD311PKtmd+WoNDpFPlZz4YK8N/SaBkRKwC
Bnsu+RU4RRsWS618OVHMkI5mrh8RcLlDHCOTOwi87PFyWvJygN3g9XUfkcZOrLj1
ltfUs5R8BdzO+qF+pndeAJcvxKIfepRpxbnXQYanPcQugELjndxHtwLBzT5SJ3cx
RGnKO8iTJ0WfR8MpDViVa/vP9YDiVbXrRr0N4O7LttWiVnjhv4WSS6LBqUnz1B4s
Ngs2NhWLg0oPRxHIqWLrknKj0kpFRHsFSnAqYBPAvVu/gIRgZMrlADD0I0oBU0hg
hu5hZKPI5I+r9ig32IMVXKez0hWcaXSTeEA36pXqMyVGvZDB5oi5Tqvuk2Lm+0F7
mAUJaI3GCCRrkOr7k/172zWQRUdRO0qFaPNxS1w3eEBh735CbfQQb/Dr7nX3aMVF
0YG3viIyBitbW7rEOYGuQewxZEVVnJxeUOmFE+Vp4MMlpPTk8G66V4RHekf3LL1P
skx+yk1NFsuD5yQDv6zYOfFkiydBwt8mxeGdXkSXyMZIrjN8FXtj6S3W6mn5WQAQ
E9KmDmfZtVj8cu1X0PnOqAtIonlEyvhzld+4o2bi1yPb5QNn12wv/b7M8JxsmeI3
V6elOHWVUYwSp13wMUcdf5dtnylTa03Uy2ewqAId1TQGon32x71yd8SpgWVEoPCP
HdjdAcuLraXbRgfvyYEFRo2Uqenu9WEtYSsSVau7GJ2Nzpkum8iD+hBXoyUuSiHn
9LxOMRcOf9chMuVdmSkQR7WJyCLcmlj9NWCCmToyyQIf7q24mZ3t7hCyEwl4B7JL
UxmrBE//BYs7A40tLT+/sfD7yYedhdyrpyqB0EWNmeigIbHqe2B7gDgDRUEoXTqQ
QoykCvKyh88gPsX2tciRvq+AXq5WFieBPO0aCcbZyOa2EGrGwKLjVoj5ynycsurw
ZhKNgGOIhWMTejHi8/0oydCrBqlDLFO6ugfx7RKwRKV8XIMFAqVz9c3DlbXpc44x
6GDcaepobIv+BjbhYIwLK72T+CJJZTzqkmhd7jtt/MxcK7zFyl7eFAOCYK3shnx/
4hPknCr5RV5+P8JEwq4KuOD9TN1S6aHIKohseRAbKd4GBf7tlCufajmIVwWBX4nz
pGW+NUjfA3kGy0nh1i5rN2p+HiGETmsudl3Ah+pWbVfqBspkr4yYePmcwKktPUHa
MdRxOEOkJKqjW8SI/xafm0HmJoEhXkeRKfuLHA3fqqU++cwML7+NDenV7rjVOph7
aO8PIvQ+a5Hzi4ssEuZWQp0mx+bs2W7bQTbOQNFAi/zz7E914kc7U3GZaw/iDW04
ndsmxNnig4ifpCeqSEOHWO13oErs2nfioUf3nNmTjfREomnjD9+z3mIXreL+zB0Z
sxJZ2HVowmNqpguqr8A/LpnY7T5G3f/l6hfnM4LVBqhhV5tCgIzzFaWlqN/+0ebZ
yPTHAX/ncs2y5+R9qe9gFo3nqWSFrHFgFEmxIVVKoMQSN6T8/C5S5rs7YRgGfLgk
OCI/XLpb0CRcxnFUVLUSmPxvgZippJ7VaBfNvh8Vbb8ETtMn2qOgJmS3NPauthOh
eJHfuxvwEbh3jss/lRmYP9vA0zrgkN1JlpzVDIXwcHgOfby5Kka0pk5GwJqsf0g8
CSxKhvN9/poLU2zVaGMKiqsX8EDa+nfre6h1xqGt07lgRrQeZowBidLCTJzA3GGE
+XVTibWIJWOG7dFp98WFxD42JKcdMBPokW7yDcja289M/W8yELXmTG70BunCHM7S
f5bPXhrBNFVoKjz5zUAcp4L6rO+12S2Rsxcf7MNs33Dm1ma4Npx0gb5t+gA0gzIn
jMobgz9CBVh/yr/1Z4ZCsHh2m/Zs1F474Ac2gt6bYMD9OyxTuvfTYhSjDCsFN0Eg
MgH/C/3MDW4oicR55410ri6LzxcxGzh0Ig7J3HZEK1MHah8rWZnWdKKia7LbTwSC
uHdN+ltrKeRD2pS7Jj1XE60WOY3FN6MOvs7Ef+YXT0d2ssoTlO26plUTht0o6oMn
Y+URDydIZanZd0ml+lJn6XuirYR3ImtFC2/soLreVuYy4tuaqIBUJCawhG+1A51O
Rpb5g88DMtpoBcN9wCpSMbA8mxqqLU85fNYmvwzW3eaHOHBvkbjF0ZvX6+rfwMMb
7i3bQbsoEnIjveaK4UP8CWXVqIigaQyJ0HOHX/BY76K4ZLwtPxcSSWFD6rQgcX5/
f/4Q1NsnxhHjoY9/ahLtJKmjyDC2RmZywq/p6qwdt5/PiT0FouY6wyJ6tpM2fSTC
rGuAd2Sg4Jr3NRyLmct23vfRGS/UKX3+tRBZ2RG/2o16ziIEq1Rvc3KpzpUAQ5M/
2cQGekRFjmBvXSWfrIdZ3EVanpdhTwEgZ/AsrnfNIs+1nJojZP0lMj/fjDLKghia
AQxVuddHvTVKbnRgP+jiQvmGcjR9jhUAQKNSut8c/2gP86iXl1qY7S1pGbA91G05
eyPle4pSdBEep0wj86P45V4Ho4/32nIsFyRS1TaobSQp84U8MTS6LvI8783c44bk
pKUmQeNPqFyckOiB/nic/FwYwaGk7EIF5uoB9M56lXexJ9fqyxZ7bFcbCmkln6pK
zIGNeqP4qoH0GKZFt4eZHkMxrM7nho7+XvaWc9RT4fDvM0dY1DnBkhI/rokWyM4j
srN3H+q1QpHNP/7UgmRA/Q7/L033scNIrjcLDuJz+B97G/GmBBlUqy6OQXAT2FsC
zjx6gyCHCxFtHmoNqUcvRjLzmIOhHNAerKt4rfs4XhO4ar7x8Or0r5VSBHfsk0Hj
IngLo97Qf+cFiFtHgRGOykWYWNPSqY4QjRCR72DYkEAio7JRJAlITFhu/U5kD363
JTlPnl6EsMZ9aI8UwQz4QtnpKivb/mfYvrOqCKJFbR+euR9pJsWxRsq7dBEFwktI
N/3s1J8gP4FTWtXX/SZLeU3dE9cRhavzVNjrMu3Y6S50xmXnzlyhfIwe0dPzhodd
5uRwWiZ2/8No2XvXjJ86/EBdUesuZeioVIeq0NTmBqAbggzgy0yRodPJggLNRBOe
hj68i9JJexJCwTvs7HhWgCVAcCEUy3fDRU07ujq1+YaZB1URWN/zL21+bj8NMK0A
9OwQFj/z2vzGQhJy9Nxsdb7A8CcaBVsIJBbVFf7+2Yn5xKXsu9LQkgjnCMfuMagC
HjZxgl8jvLtErBgCnhSMNV83qK8l90icl9Dv3ZNwc2mFF8dzS0ZIHUc4sBAdDnpY
CUd6MOVbvhEnwKv5ixZcyM77qw4vIZ1uagrKl7CduNhTIBVy9XCQ4F5bZQdsThuA
Yd6lc6wKdvfczfclPqd8yCGaktDtHo34iikWIINctIts3sSbcsOnvhr5IcEEzOqP
gIWJVl3pdc1GtTv7+jtC6K0HcUP0L9/GhR0TGbo1MnJKB8CFpi373VcXt5qp0yD7
LfOfi5We+n7LE9aGVEUFr62vQcQ1thsBW2ZAn/ESkPLifT045r4uv67+d0Iw6a08
7Nx+VcjVuwTLc8HCmvgMTIg+HGoI2kjutPYxjpyBXU9LhPJf507xjBaZnunlfPbs
cQwrH7GLu9i7a2VxLZr1OWcuNz5lbsp4arNmiMCbMS0vB4EuW9mmPqJHuy5bE5Y6
YaXGMHiL0XKLAQOX3yLaFLGhbeMRW6w++znjM+QB28E3zEMY5bkVEiMSVfhxfpsk
axIonKqCg2JJ3GpAjyioJ/FnwKpWSmWZqyswiqicgFFOuxekK3dm/AIg69eZqGdP
YgB6VAnmR22cTweUzT+aMD5quXEDSNRj263ZZNZxhimw/ZCZlaIL7xIUGQyaMN+P
XraOuwvuXyz5QJ4csLAHFBmiR2ID0AdourjH0su+dssXCjFH5leViC2X76+qUqcK
GKQSt29McOLITqBuXK1z0QdmA05Noj2ouD+VcBBe1sLv1hQKmMarskNhhhZU4YYO
SEzSQXiYj/sPPt563PtKnR3xbUPLJZr4DvF1spxeOnlQfRrq7U2dGmk6KH3jOATn
YNmPm9h4BkPG4LsyHOfVQ+E6mLUCMONrGK2NCv54QBlVcKfFIIs8qaYs7j9fZGG2
nqm8plz9syw6xUwf0NaF0BD05NR977YpxuxQYvLQBe41tHIsKnBRTWiliCDK5PIH
kxgsbAV2c6j5HbArDoxtbopSl/B38fWaQZ5afTTU6BHldPSeK78KAGiR3H3L8YBd
Ms40V8/G4oNeXulNSHJYit0t1wE80XbxR0XKP3AoBQNwtRBs4u3qZn5XYqondbns
Q4ECi/RzDBO/6XPUjd9GPeJkMXT/2nPBJrhJUKaKyq8Mn2vtuDZ7ow5OLc6EPulG
o+6MyjaHWK/UmxtsQDSPJD70DNQEW7Mi/SlFTBdrfGYaMWRVnCn/JYP47+QZJlnv
7eBg8B71XESVHQ/7oSKtElORnJoaoFQkKwPQM4Tabr5lwLzobHSyzd95cfvomH1D
JEOCdxe+Auay4MB8cV2bAdmjzXZxZ6lQMGQh8Q8m3MA9l9tlirpNdDeLbfMkP43G
FSRsj4Fyspr2GtTswzICSLtVjrdJOBF1Egr0L0U8ucmbtKEmLCDtfBIl79biV/+p
SMPaSHnQ8kb8aTVphJdN5u9+nyBH34q8C3+4LEx46JfmKPzLWYMw3mDfPLhE3c0P
5Ca+b+TtKrM7N30ZT1k2/5AFT5qTCUPYHwSKpOnsoV9iYh+xIsZVt10URq9s+V3b
armP8ViUCwjQqH4PqjnIlmUxxbIEARjf7IacXm4UzEHyOjyYhNNykhCd8aUeOPRQ
kPWnGV0KSRZzG0DVLuKmCakURJy1qyAa0B1XOZJsXNs+3qcpId/yCw0ECuF13uk+
dxQ31uvIU59IoX7cq2Gfsx5iifO53FhaKwlpDZ1zlzxPhQs7WAlIJ3kOnxszHe1a
aCZPZgVui9VqqSQSHvB+7gFB7stSel4JzSlmfo3weHPmWYRlWooTLE3agfexiVLx
2mS60FkLnRaQfQ3hEXFcdpePhsm3LufoWgxU8ATqgceHXGz0qKVzEQO5zw3AEdpf
pT5LY+lNOm1+TGSFX2Ei8sfWIEaZfrY+BMSk6coFSC2D3ZbDRua0+bb2lUIHeGYQ
jgEJpxDvk6I2jVPnhxCMXwzJSAhEAKHQd1OHSMiMdULpvI1CxBk+Vd8c4Pj8/g/f
qa1DzO4UNBRGFolqvgmE8TKn5mBIwPR+S5BJPTEIZxgixw6afjzMjpS4RtqacMkt
26qmfmXswKIaI45uVNHa7sWFh/42ahTQr3BgQqukKJZVjx7ACdfOTO/iOnespTvd
BcC+t+v6OKvJohlwrNwOaFVViY0DJ24YRlyxdHAVmKs2I8Gvy2xqET7YKTIqXPbj
ccaQyfDnr+DBrGWTQ/lxBjDuJ3Jc/jzdcG4+YlLvA8zSANRurs9l7J9iIYCrq+3C
UN+YvPFORP8Jxz8Vg5UJ3fhP+JxwRUNPNNweqaqBJnLsItslcPP/vPrvV29hhLHe
fvBJTstkj+GNNy6PyRqy5JX6SSa6OZzNpHX8yD89YLpNfLE8Ibk4wZtTt7DJdEhm
HWqb38Bts4BwNQGeZrdXjoEMEE5DjqlAickkQ8vZN0faNGkeeM/lK11dJ8Iqw2Yt
c8Jl97SzgpdPE8IxurLxstYCzMY2T6sT5AwoHSUthBwmVDyYkM3vvupLcFvo8k6K
fQcYKhnByw75PGk71QZ21UmLiQ4efG6PnmiVzwMibYjKbXVf3IO6ivvauZABYGR1
39oO2ZwFhSEfM4CHLUQMXPq33X61CBAUiUuGKsAF6lMt9Aaku2kmjRhvM/r/WdV9
s4ZMySP7j1csa+tOzFzwcDhzyP5LQmWfvR2iI85x/Vla9BI27nBl7KfOt+mbFQT1
VpXsFCEt5DKUWhnbzu8CqJ3tWypjVMi3zqeTovmHz5lSMYTYOSWc5VBOWCvO9N9+
FlvZ+HK4TJj++b3lnsg1l+jWVMar7MagyDJABOysywUDW8CfRprl1JEDD7/aTtkS
Aj+//sRgd1cVDXp/Lk6bLVkATO2l50+7Zzi7Rbv0/09JfajNARKaCASUx347elwl
XZzd/sGBZZOaS/tub2YuIua+aSs46Cx36el0l7EX3u1bvMmUB07cDtH9oYO2OSVG
JEmBDpjYPUvIA46kKptp8ZqQor5NSfJ7OB/XkWOBQemVs0EbFBpBi2BJG0d33ghq
nP5bDlIljtUM4LWvzHE9MaStXnFLge+puf9URKVog+qb/DdyWNw+UzLLJ0g48hQE
DEWxZ+f1Z/1O9h/JJrxT8JFbJ1vzHNMqkscMQn449ch/9wFQ08a2mJG2pYQOL0AW
2PGkfWlY8623eJ5QSgPCLhCtUcMd0hP30jYp76JkVCoVB21qM43O5WICyVr9O/K/
Y45MsmaQYsYAwRbCx0CwE7h4AQGF8s4ew7sL9yeedu6uusfDUWuzDCYnntlkn7N2
R1Z8IGy853ltnP5x4m5P3FYfkeUg+vE9U6RkOuQWVEdSRTvfuA7kctNtT+oFO2n6
hdeAqkQtKLxwiaVBPkHHZBJlc5SSpZmUaeDaQDIA44vupvn8fCtmS5vw2Pou5zaA
Tw2R4cPZNfzr5gYxJRiBjs9v/PL/3hftWTV9LsRAX3Ne8HMh6dV/xHiaK11ZUaHE
/Biwu3a0bsptAyOqrAvmkGsRXMZHMNBwXib7hBWiMC4uxVBLSAzJE+DuhEIHIa2H
XxpWdEbqVe8OlE+LP6xp77RkKrbTd01qIh2jDR/QVubrHy3lW1PLp8THY0+XS1Av
66ns6Frr/G3wOXvBTZhvTPKyDhULyj/oWAxQxUX7oj1xqDMhkASAVf4CIJ4pG6xb
pDtI+6RhBB/hBu9QWCv0wg7ZD9RgAENP7Wf8g3DG6XUMVOW8Mjt/S+LKjFCDN834
RRuhSzOfkBmEjLx9zb+1Z4Q+akJdaHq4ChFh8pc7HztFVKSwQ1h/M3vVowfoyjBs
vwnuQrj5je8Fk0wWnjxu8t00i48a6GWOgyDEXbe7DLSwQxUYwtjWxmR2DLsrRV0M
5u+vQOd+WONlrF+sqeowYKyaTLlnbaUTcMhSntYX0si+QVB0G8aDwuVW8PNaruhz
g71rVov7Im8iDCgIMyf6OYkaPi8z8aPVUd1vDfnlvQr6GIQ85XAQ7Tx5YqykXvKp
oaSl7Fi+t5+l+DkoAH+eBvH6vM1gd6UMAcd+XEtI1WfmJqfprUoLw8/IpEePAd0x
P6gDY2aGCu7DyIIvh749sPK0bXg9V/p+HCd185+F0579QRHIV5Gh+8h3KVflsDlU
SEtLT75GmFlIpHRUIcu3WsTDCMaYoGmDYsKnrhDObt3Zmg6YmuBqplFOTF1l99Yp
HI0fnrQHEO1a0o4frtUH6S57AfhF0WCJwWBbuKDEklq8V2tgnqsW3V+jq936OUF9
ADlXeb31z7gon0gQOeXh/h0VKSvT7lR7ASqRzKG2P5KB8xxmYM9bZiN8ZB7qV2Km
E3aIltjfOxp9ekvWzMJF2BJJ7VrnLvuQEo936dnNIM714WRVRBcHU3CAygvrHxcG
LaU2OglXX44S0zD9j9qLdNtDcuAW2SdFZuQjVAEhyt1yNKEVC6cPdlKc858JjUnR
Sz7i/9BFOzMRas54yjsX1Ic3MThdME41bduS9iRc5Sw95a2gAx8d3bZ/abjis00Z
okS8LyfOAwL1jmHLFi2X1RgVJptRQPnJLjwFpZDQtkunmgJ19XYTE8ugu6UilCXY
QzrS5Vltt5p/AKLWA06M6UbmdahyVXeOATGyjrlUqGPWar8ZzVDwpH5tEsZwUH8x
vGMWsa3Vvdu9X2TyZRgoz9J8piMaP8t7LH102Cbt0cayVMXlgWEo9JhkMXu3x8ki
8wmwaj5oUUlabDrHp2BHUpmU9vPv6Dc87QijUHOozOdzRMvLakgT7KzXU/MgW8Ug
RO3gs5AiIVGmOJevbfACJDedRrEZLzC6RwP7g5wkMAAKEL5nSFNyq4xtm7NsuMGE
OlLnzK0DZY7Ocdk1igtWE6aNP1pD41mq20a7RZggzo3ykGi0x5HF7bNHAIGgzlKP
9PfUQ0/Ygs2HkfOguSyTe26ZTMN26hah3Q3LHXDWwRJmF7997Cl/mtLheE5VTElS
xeKzmTky0k1y+pMkafZjGCa2kyqHMwLK7mXWkA26/liplQvaRnBv2D1S6mUrc97X
gMZ/A5vWgi0EVfE7/aOBXMJrz6pLiUEmMZWcY153RrylIJQ85h7EhLS1hkXCUUfM
dnFb+vgnbv9l9axCsmwwF1WWzQW3C69QDJMsKQRzXSryyEFXJk6Sp7FLgAb16zfQ
RAbPrdd6pfLsaGD6y+TuN7zHoOutn8llBiSv1L4cs1N7MlUrB+hJUR8r0vdszFC0
f6vTQEwHEso8aGtNQtIyLE/cEoCUm2YB3wj74LhtoTkf7FRagBMmFvSoq7KPmwPh
8jBkrVPbwp4BiUAK2mppyrR0eEA6y/xcYiQRz53vvTB5t7LJJ9HtNnBso9Yv8icR
2SbrD4ICBe/PCf+D9iis5lGqQ5/urT0GhhD3ljCYdP7c5jBojWrTPZcvzDnfuN8b
0WzzSpfWSF44lPFDRK+5pK8KIM6zesOT9O1SzHS1lUEbnD9jfW2yAQjm89HmJkQ7
YPkEMW7IpF9ph8942mPEpdV62x3p2GbqZsENjOkx1MLKjWcU57vZz59Z7SMgFxUZ
FWgJwKXSQ3wMKjtz15oaaPsWcgWoRXyTH9DM1duhil32De0MdQ2QBZibxpBoWLW3
odWDmvsE6PEkX8Z7FtU7QojS3jfJEUK/PctRvyFFIpzL/MAAVctJxcBtx1KcmfGQ
Q+U5FE8+6Zm50mX+rizYx0UjZXmI18Cyz0R62gabw0/t2h0IaSjlchn8NaHJpyQv
Az3pUsgHgH8STcLpi/ZPLzPAA5zloNomV/D2gkclMMmUQV/tqRFVMmE0c9aohVGK
I3qWJ2TRaz4AMMdSZbVxVBo4ht0cMw49Gg7347GdTaFf8Zrd1qmOMG0XGQIxxYDH
Ne2opx3HWmxuxbLsm6MmNZs1dk7kIrFMJ4uOuvIxvq9+LbGyyNez6OUN/bXKac1v
Zc+RdBPrWWUQm+v5iEeEEGp8f4BqHAnnstefi1hI+dbzcmVLY8qCloPSur2Mkis0
rUsoK1xvt4zR/uq2q3HOgbe885sblUv9otaj2gXl/iE3KEQHCLwNFbMMVDePxXTN
WFnPy1Pq7KKpVVOmxrjkEuOLQq+OlnoefMELdsEgcnuSCzsbFWXIu0AO/XDvkRHh
uDFvLlk/DQkuAyM1meGcFW5KUO5VquTqW5sB29MqRJGU1U8oRMJyOH4s+G1tPc5z
4QwgtYbsFkKg/5Iy3scgHqG9ObksExuSP11eF9dFWovC3YAWh+uaez/9XWENq4Mo
H81ifUz/c0imlj70kT4NXIx2eaPYG5WQKdPIMXA+bycLd5xYq46ASiZAwbthDC4y
8DsL1Liq0VXQaHZHV+B6D/MFFWy/kK43WE03BATxnOvmASBjgPD91CfIi9aKYhlG
Wp+4fQNCmoyXqVy3QNYs5zwlONh+G2tr3PEg6tWze6n4F+HyTSvAgWvFfFdCZUkJ
ofOKqnzjMCi/GgZ2rs0ZoCPUD9GbuVXEwjlpyFwwzRqI/Ku7gWJfCaJGoxCs0PLr
4gzelGABgnpmc+Y59wbM9bISxIV7wHWom4SemrUx+N/30+O/o8RHL8sNeNAjWy+q
j/XB6vUAmRojFjPP9RNfHkEUCswooeMosOQdqduwuqYpc5ifO6NZT2pdmTTNcW3l
gIBevrG0p9awePY4xjKjiNUKhZCjg5BhX5Rshr8u6eDtCa4L6egUsKGogPbYzP2P
8PJbPLERp+kbKSOP0ImyddBMoh1KnE3y22vVVobxlIgYLTgxyrRAySsLzlEpxDFu
y40y8Kqi4y085lz5etDHLIrYcAroL9BSfQCdSpQJzZtcTiNy2RQfT3xdn+OIzc5q
ddmO3ER9TVnMYqllblpAxW2v4Qmswcq8345/wVtWPsQ2rj6PfWKhAdnaxxTtJrU2
tNeCzlXqMtCZIuppJo24VyRTBhBGaLOEkCWFmcOYxfmZsOYZhSAHZOV4kxCMsj8j
NS+hTzarXBvLy0LXyv+DYfOhUceYe/04UYQuJileGYp5rMlgAJjAtJ5Yh7dBxnuX
8KapWn69xkrke1mfrf7/cRZkyVFL3OOoq/fStFZDMLuxAAN8RpepzOX0JLNs72Hg
btk5NPlI4/tYGf55e3uXt4MuAjkxN8TX9wPEOAsjv4Fnp1lZAFixJKiISG40LuY4
qtcPDycNmJ7ZqvfWRyx8ZLEfj6pOGaheyTBZobR6R2hWXHRnoHi4Ea3C0rcMS9yI
h8shdKETK/WFp/tTcJGeQVHrp6tsszY8j7vTAsM42jF2D+p56m1707j2pBilO0d4
i1RNAxgwXcpJ9GO3GpTBepQ6kHWPFWt0nq0QFI3xImLV8N6LvWVlH0kNr6iODsOq
kI78sv7KIDcyZgGAZ+nOOTYAXHtADNTgePx7hA77U+2n1p7kbsUtH8QheUrFnDaz
LIPg3Y7pNIk6KWp/EyKsRDVFlsRKn8GWAhvrDdtiWwL5Wft4dDT25RJHO0Xff4rX
h/4P73p4xT8BZjIaQ/2T37UKQf747csSfaqPqnPvNxqAypuuY7ytM2k9kzCM5vdd
WkqfRJkKo3pP5w5axtiF1dfOWIMq4RRtzvqD++M9U2fWc1IHn3P5mWtNN9UaKZLF
QJWBlKErFfSQBgg2AuleHnvEfK6Ur5lLPbIgsSXG6VZeMzu8DjyEeFD5dvXUsBz3
/AeBmDoWzQTnvUCOEJfQn3LJMex3mLbzoDhCqcsCWCBdZib1dZNpuMXGcqgYW4Qg
alYxBddv7haIS8+PUlXpIW7tarW0tzzeSgjeaRmtaLaaS6seFR6irgSSKzqIfYQ2
1zzzrngXzZjKqwkDnVu3HM6ZY9nWILiUfVwHiWGKvNhiijX5YT/fBG7NYVzl3dzx
BStX6EPwsAZzGYKFfKoZvztGmzFUjO8jKb63KAdTOKQNDngt/HumqlKiaO9Mtar5
SHQZY/CQUbD78h1mPZ+VpmaYjmZZEovoDU4J87ZSqhnr6XsXrqIIAMACxxlObe0m
wwyyrn4BDC7nmNUXdjO3ecOWor8ZWzp6dCs8zw1+hvjqS3udirZNQleWeHTzKGzA
C7nZBE5mhD4vBOxhtgNZy1/fl2m3M5NHlCWQcSf66iI/7Af5kiAEzbGfKxb4D6jl
JVnSghZFIH9tFyL1RG284Hp0OqfDdjd0eioFdhkjGAAeCbyqFFanA1KFRgFBsmvu
VJmB4IfTfiGX3se9mYa8nq9zZpJIvw+VeCuBq/cZdmHXFo62Xxk5Kovytp6PTj65
x/C9BWuLa/8Bftjh3njzyKX7vbTMnMJKKWwqh0B/nUCiw9SDrbEU2gF6vWqoiMq2
KdjfwFkB0B8fn8V/udc7MDoYyVkaDIIFuX96kqhI9EAce8PMf+X9fm3j9997cz+7
CG0f0yd82TcH/+AKmT3GNcW7DbfSrnD8ICRjd3yWjRSwb8CDJRVjriVIb7TlM2P1
MC/ZcUUUJcU1EdjxIKph+Fn7FATb2C4sjkUEohNes8zv/eFTAOrTZq3wuAx2Wy7r
oWw523EBuuWlQ2/uTeWIgbxFWv5hzFp62VpXB/ppKunHW0+UOZdCEYEr1ElLsDxY
3uKb4vzh22RzcTDG+rhpM1trMBqCoCKVptGS1lxZtwWSr90jcUNohYyMzvneMLpz
UmRqbd67YVnDZQWLUk4WU1zvdnVbuBsvVuY8+26ZagP/q5kQRgoKfwaCNO43n+gK
HkLdxdOapvR2hcatwrL1vF5HyXhZdbMTF/wXIAZ4CcBqsX+IFE7Z0IjZhYyOkanc
mZLf3sd0uat0emjoqBMMz2yBZDfyFpUFwES6rl3CNXcA5R2yJ8fFvPnvpUOyuEVy
YGrmd+NW0SM/tkXSSuRvk/LQt3AlPqCMBeTf4Vv88SPAfp/NsoXjv5PIspd2rmOc
Z7fW30/bZnrPeburn+5e3dMBUnlFHsipYhRogaMOys9L7LMiLZwO1s40o9GWaEG0
H6h2XPIPFR23uvytaFsvpbT/3cd16SqjW7s3VGKR/ZVWCdXYc8/UxvEsx2aqo7QI
0XeRA1L16+cZ5FPWteIDE5DtP7ss0WqxsQ3GTBPfkrBsKcBUbCv4HL4B8fTs7UJh
vI3A0Q9kgnkRYhmjH/9TcIBIKARFzD5byGoaPXa2spfnxAWbcnMUpf3dqzLDzmrt
rYsYw4LFlGR6dtwClttFjzp1wGS9/lJmtJxRN9B0dXD/7ZMfABlYF03bV0Iz5cia
ewvTBtW98lKte+Go7UWpmL0eChQCZUyqKAS8yZFo6f+7bde0VZNOu/5vGYqDh39a
HdKFrODj+wA2I4+qXuMbrR2gbheLOOQPDim5EEByiEzhU5hRScO3DCcs5fI4q9MP
qBe0rciR/G6Mxx00FCqOzG/jiZsp/ubC1LNyJ8D7lxC81jMLJL64aoHMcv/w+cvX
IimBBnsU810E86AsMAW6VGd1XO0iA3fxf9c/paeVCqDuyO71lqUT9C/vqhyS/OOz
N4gHE1sS1VR+x/rr5b5XMTfHsb8+5TiOmd+C2bFZBFR5tu5i/hxB0oJSvgc5LcHQ
Tf9TnvXVspCTqhb3K7rX3NDYQ5yvxGHNMkDBFRF6976EjhXwsM2TzsVgzN0xh2C5
9v985vrX6r7NwEewRBIc0aepPgvgOVpDBsQCpo4/o9ruAVX24/fq+FMOsJfAVf/i
r8deATf6XtLIh50lLjX+CAYsJUoR2Sg5VfYxv57TReO63EBY+pTu71ESzzvMPY/9
R+f4ipK3Sr0xie/6KcizaS3oqs0+6hfO9bUmYKYRjEVxo9VcSyM/ECPofCGg4Nov
cgPFryOG04lnOMPu6k260ACopxXh8T1EBn3sL/lvbKu3kW4/Hgl/8TOk+pWViFiV
ZNIMR5RuhGI1odxdkq+bDhVOm0FKGLxCqf8afNOPgaZhwjMN8BbpmRt13s1n2eJ5
AWXn4Y/nlCjYMu/tydTRkdTqa6IIUCeS/rY77wS82sUM6v1JKv39u5s0s1cIGuve
R88NOJA04bXsPLk6txQITdhyPB+SOMY+reYujnS0Tq4fjMOtY5XuzdlYDsheBsoo
djo+Jw7zFMuLp8H4cmdv9GWmq0kCg3+M/GhXeG349RdCOOATzb1gqkTWcx5Nn8KN
u126vZuTXeunmRddkXigqe9ZjKrUQtPISCXdDLKcfQvMTt+dOnu2zdXNsa0Mulu0
uaxg9aWwu/y5n/3fg07H14P8tI/PTYSVDLzllp1kvyeZns2fqH8uRMnsSol4jFTb
qj6677d7l4CKQolYfch54hZgMMAKki5wt1qzymsB+TC0mo1jKGD6e0mZkUfH+3qs
gjXS9JVHhy3pTjamUMZ9Mo6KuD8qXh2ToapEVyhvpZLWBsA1Nilo2L8xAYny/JZa
ppDabjxdCgOatWgfSTfYr2t7iDGAuyZU5gLMuUN2z2b2mF3+niY9PRZ/7ewTDOpP
2eNGnH9QG2RPUFYgD8NJ46Z3ZTWQkGL8PS5wsP6Q7S+l7+cMKbzODGY+pmJ/Rv36
nYWGfE/4b3+V4dF+icnva063geTtaexJfwGCrrAO9A4QCvsILZ8+Ok7WH8iaAu3Z
iv8P4T1fIBeAAawuVBQo7zQWU19fUUDgicDctIUJRWta7Gcx9gbp80FQT9zSug8S
T7eOTE8V5WWMSeI1KIzzhkVlyTvV3k+hAozUyzPluS42UpmatxIQFzThyCDYP2lq
B49CpLeiHt0DRMdLbmBm6ZU0TFy3qIu3otDyPjQYnI2eEQ0HTlcYwNW9X0H/EWQ7
HqMdez2uqsdQtHSGFyF74qPqJehOusDjdk04x5+Zbel4fsEALzXxyMaqLkKObfdA
PEq/MZbwM+jKvLCrjkSFtgywEn7795oWhdH+lEluQrn3Z4T2T7vUe6QI3BLVkquq
m3Q2aGEEyu5peADENy7RtJTF3KfGOh9h+dOASsAj5c961DNfyIsOvpv3wUDjw0w0
XEHWJt5avwWgEAouXsoxrHEYZ7xAlb7rLeRfsAT592Szeuz19n1umHOKwNDjhBvy
aZsJ1JqeFSG0mjmKPOh6mF1HLSpACf4QE5qDM96uS4206/UODLvliCjybEb+g3ou
tCo4k1cXXsfWQzQMF6W9vSt/4scZQngePYiVWKbCQ4LIL6BNBvyPpS1oVpVyGiFV
CKiy1jS0SV7oy5ZA19KQarFEaq4ywxe6bvrWsvRP0eOWxkF+kXjXeEkCqEIhGRvQ
4teJb5OiYe5/JkDc9GAPWwQWEtIvgILfbFFv8NS4W68+821aEgmo3SW9DqdjwiN+
1kBt2kDzxt0R61Y9EkCzkGg7FU6LmrYYndPRATI4+NkN9Us1fwFax0bJrq7ZiAKw
PFMg2bu5lV+mDWmlX0FESKNzlj4DKRVlm/j2Sbvz4RvBsnbdMhJXlfOnnrdX6is2
aCPfmsXQsvTUZWlD/G95+IVZSsxbPAnKGXM/6uv0qDcY8Nc897JZNaZWp1Uw+a+d
xO43oDaC7mmVPwj8TN+vlDJDT+XEuBL5HBC3J1YZEPMQUXL0NOwVOIQF97A48e0z
RGWLcodVxzLD2H8LJkSSkaHq05iWZtGBdasj3MMt2SSsDAu3zCXpoWG9raVsdcOK
7cSnNToPJtEGua0hLV4yEusWr2+usGX/iHhPa2xHdYxQ12p49tSmjF/x3GwCV/LH
UqTp/eN/k9+KXUpaiTXfPTzdPUSPqJrBfECr2oRt7UZr+pM4aOiiEat6LG77l+G6
49+UYbipfsQFWY2ywFVtzfPCbDc1WP3lEPHeVNJcavgqjUjvm70hk0lkGA6ZPCxs
llweoUSNIiLotw/8mlMpWw/HFMUy8iCS7OT++RiLoSeNOpEPTnrAfkD/G8AES3OJ
QUyJ713J0F5ocUIbz+YlMn28faaWWLevQfZ4tF3k2dM2oDiwpJWR4dN7zT/paSnH
SZdes2PLfd8QZaubpQmZJZ0HCCd0nqkTjY9TXJoOxLVRDaA0pS0OwAlQPdY/CNIg
q045+EJTXv06jip0WVvSIeQPvrKrVy6R7qiKgvKIx/vG7Ztv7Nj05VlF8IdMVivN
w9yyOTWy93y6c4xq1eCVztP83Q7W4xxdz1l6+p+ow+otW4mlDkJIfLzdElisLPLK
vbRvusoGBFY6GTElDVZOX6fMPYw6Az5sZ7tI/8HF/lAE3sQsEnMeEz5FHo7n2u2f
aa/Raf671fIB5GHm8Bj5vyIhJ9FjMfDVHYO21v0sMcwdjgqIu21gTyYpVAxbdDhl
3HDTOMRM8iNy1ZL6Xwr4u/sd5+M/LQ0vO1CJATJUaxQcvhCwWKEr1EeUSf4j1Hdt
X21nC1AAQuZ1mjlwd7SCpCXDWiNBKXSX+5GkCWgABmtrj74Br+lKJBjNNnnIixjl
+d8Ry/dwqMs0FwJgJyDsVMhr51DYR0FQrJxAXWdSBwbfyP/axupBF6gb2VzV2/0A
ivPLlf5z5uM23dssyYs6bECOTXaUhX0gwyFk/DkMLTy1VwjDULkYyi5rCmQ+EvhC
Q43c5amPm+0Fe6ttNZsUVZC9iyje1PubMJeVL8KxP9O/7wKSxRdkxfVUfYUdihwi
Vu0kT51fW8kFlthh3rnCEZ0cyRdZUR2DUhPqwh6mttLO6S8+QzNT9EmNV6bxDTm0
YFufdxKyIVtDEvRiCXC2Cdo/wJ3pL1rUvcpQHGZHe533WVcZCR818v3T1SAMUMr+
G8KRnZ5vWG/ZUGP3c9mDwTMgZuUZNtHi/U5f/YxMoelpv1ZKGWVmFUVFH6QcbKAh
N5xL1e81wo1Z0dvqY0uSuiLUJFFqoUwqr3DamI17T1pZYhSe+9EePkHcEpzqvZkY
bKy5+UsOQiusCiUvEN2m1jUNyoGIU0syae9I2GogSMIkD+DwMQsyBe+ytiPQmeza
mU+s3hHif/cNtZU/2NS9WLZ3iIglpGdFaOBGHx6hxu6KSvqF41lexLVuOdNtEEMM
3vxVN6AdBbbT3SEs/V9wMGpdgW225Kc/k3bl3aD86ydLzuovCKG/r4CnDaGdD8Bg
CKr5eSua3uAh6aizPTz4cwEeVFwV5fI8AqH9eQho0LW8gxV+sdaRmqjjemnYV4/K
ekZtashCbfYmdEOGD8IXS5lRgeiBm67x4U+HE3QezQzqwGQ3jWSogiJyWH14ly9E
wqGmv9mprYOOrnMgVF4QWyi6Nt6a4sL/zOhr2CLoTPvpdvKj1WPT9Pniqe00wrSj
aaZmr2Amzo/o3fQH2OdAaD75KucOM7h9LCjZG3/Xys1XrCY2IIS0ZIT2uF+itEAD
PuEZtt8/pYTlIVi7/aHYOwjDH1FpxavmcBvOU0nZa2m6L+4Z34HxA3SnbTnTwMMx
e3oaiwKtv9OAYOqhtp/7fYZr6usevX/1TwDjIUnS15C3XhHN1biSkx0s41i9lIbL
pluE6RuHIZ7LtKHf8MiQ7+i7rxQRo5nINC+MPp2tTpdZ2bAkG/AmMf8dCUeRHSQf
pqkMGFmyBXy3Q0G82syLXpJLwVahKafWFyp/sJzBQ232r9Bk5++8TXhnLAVVorlD
rOluKZ9PuGWTY1KAprsc/f6LyHWIofYQ5Jk0yQfbxh+F1wsGQyjICxdUHTXVaK9g
J1Pkk1sEdPEDozQD+/iRVqxJgr3xUzcYPgvI/rXbrSvT+8jEgV1cl4Tl01dmXItf
EJsPhJNP0l8NJia71QiKlj7QmZOmVSqRQG/sO+nY3iIwXRgpJHoCm1cRmmuLuA12
h9P56m8c1yU8ZEEc7J7fYsQH83kqbrh3flDK4h6z/KkORVsJQy+WYK6nUJpm+Q2J
TeTNiPN8gWzaYD722nd1lrbTl5isDg40uNsROo+H0/PafHFcqo3hTYgGHql1XdJS
TEEbnlxL4BsZB0PTDLZXabuizLP/earoouKd19lpVyfCFOmpnT03afXtOLJmmdS3
8BM9Ty8PeDblWSsXHae7W1hFNrv7WT7uMTkrBvwirBB3BUzBpwHhzHA9M6cAENIH
R8N5DXYr/Y3nX7iZzwazcl1/T3Ixy6yeVLPU8BNSb+sjHTRg8XtkwD4nPJpE7kKc
xSWuBv576rJy05cB7l2Bmv9EzGk6wBwKJFedJetJC+uJ4HT6EjKb8vCbsUNyKdXt
JfrcPF/t0CqUWFxpxA4HoRMyS2E9AM53Ojyv6QdELEXP85s8r3ImS7x7LLFBwJV4
yj9nHHoeLCp0RO/ZEDDguJ6WUA1AYQe9il2UEPH5+fyg0q5qph1tvF4Z1v04XPjT
+Wg/fpswwl53gA+UsLVvKdDiVHUR0bnc63iA7oUa4RMvyHO72utfNGOg+mabDG1V
1nUoxk3EApb2I8yX1t1bELgj/kJBYu+jjnifm4L/5RuDjWjqYbTz5W9q8bgEHWY7
EjCw9sykbQvT4ExoVlqXhwEicRJWPXpG0hWyd6BsrnXRuZwK9xKOr0N1mPVPBgo2
JTmi7R5v5X8te9u1vyL0QbY9jQU/DL1tJf40MYGnuh0NrOFON/w5lFZUIsnkldjF
MjpGIwpDXK2xgl8TLu6bP+97nsOfbVSyVHfClDeIKPnIudZYugVVvNtutuWQsms3
Ov4Ykyj2/SDh1jZZ5AdBus3m1ZhVPKALxsclkT1BxugW8OUnttQwuVG4epJABt97
wyAJdZqaOuihEQ3dXkCqKeNBASHKu69TlXMA+3tgfzBGkeF9Z04aPQZUABLgcPNl
rLRyUob7R8r38JD4QyoByWmBb2BchiliXzUheDY0RTKdCUwll4DYEyxh6tZ7MxUM
l5/8sgWFEs2IIcQwJUenZPfsjTeveONDE+6PKNE8X03bOPPv0rqpL6qOaRyj51Er
UiB80mSRtntdwTzWT0Yri147+oX203gBXOhOeAGGtnU7JPHt+lldF9dnZBE7Ubwg
phbfy+sBo33p5xKJegJu8eg6CeA8I9oawrSNPUc160DkNxl4rhi90+s0PlnxQ08d
5G6vL3mrUwwBezmydz5Afb/GgrnR3TSM0j4EqurVuCzR20dYtCN6BCpVfXZETol1
SxCE8dYrU3QWSxglZ+SuudZ4HviCQe3UyvXLfnYAWUocnfIwTmBRIhHkOAO6HKa/
rf+SPuJKr6rhFjzgQtC7FFC3QT4sdUiGSGIOzaJC0/rhk76ml6rPTF9A1PMInogQ
1A1UT0+VFt0SH2n/NcVVDcOiJ8MCmoa8DrklTdPUC/5yEFcQvpus+uhFg7cp24Br
oqNu5wymbxlf+gTHOJ86ZfPWHnWf6OCtKlEuSYNIqrPFErPQhCYd83c5nDYQ1vGV
p/XJ8QIsoH1uQGs359LS3IFFhAHqIssRc8Rrl4YWMHwmdMJBaznvInYKGWTWxNAH
jKDdJ8cyMHyPVOF5sSO8yp5L2VjodKoXCkjCGVInqq0YdH8/HJzITUCbvd8drnQN
OepVHHi0n9YUzPcigg9MsWu17lPTH/ri6qtnsZsKZZG5Ku7nnp5v9UMvfo4pMgVl
UY/U1IYASjDOKuwsEAXYYUuuRrW7mVumD/sp2OU2Nb4hT1CMg5m7aX94EZosELmn
Fvg4r00Z8/f7f1BGIQ3XATLLZnzKBEzn59a+kb2cuole6dnn+xblOnxpvkijqGc4
5SKPLHmAbvU5Z+97shwq535u33KyNqppdhBSN0MAJBK+9VE/lNg21L8PSuiqUpH0
F3K1QJhC9F1OKgMemRDEj8uZnga0M73VcZesyPcVseyn5/Q3572y8H1SsAnPJOzY
r901C0IjGp1F1BBXr+QkYHx/zADgmR2DBilWTL/5baA4iaZgx+q6ccwD+XdF0Ytw
ocEJHXx5V1+0ZK0gFWwo+6YTnIOolrrs8xlQzpx+W0vEq9CGYbA2GJ9ydChc0JwH
rtqSbaQWSseiulvLFKZHGyJrpeRZTugXII18iQq9EutCWjx9h1wNjcJ/1pL62DQS
GRgYV6lqi985kf5CJQcy/XCElSK6Nsr+40y2Qjfou0z6CbFU+YxnkQD0OEJ1gKFu
CZPEmGsWDO1TMAuococZp/bFuXDU1peMgFZYuiAgsTF8jJAt8HwqTgWtKQJUSim1
jyIKdbJOaLto4wuANcV0yPO6igtE7iYAgXVl9KT1hRMyGLBpvODr0N1wPD3TSJ1b
xwS1mC9GFkXhaBuc7wF8KXSDvwr2A9mmAQZtWxLFMsknP5wnYJMu4xL8IysntLcU
PwYnekNgmUoUune23go9MA9EEf0ZW4whAmFhDWlTQe0KKsPig7n/nmhLaR0BNJZY
XKvMkmLea/klFztdRsNazdU7KCuuc99J48RLJTS6sCYW1AgB5d+f61GfrIns5ZE+
AjT2bTQScy/c/59vYDILntz3VAmvTcIS1RyIYih7/dfAmmYGf+X7Nkx/WMTqVVJw
TRRKrrLc30/+Sh3piGHUYU6VrANCuNiqpbrCSheZ444bY/nEbdMMPCy8PPsHk+a4
NizHEhUZJcymGKpx01BRGGrccE6YMzQq2JF38Jgt9FYqrsuMGixddqnrvw7WzUET
PqITuFAUKLBrQt1N9BWIH1Aiko8IrLArxe9bZ0THUEwBC3nhMWEd0O1tXn0ZT9F+
v83xecI1uZX4gFFS4AUPkZik/qTGFLFPHGL8/8/rPZRsh4k/zaRWdLhq9nNFdjoz
Xj+ZxyVK7k4I9q3kUjUZWfN+e8vtL6s2VVjOIJFZ0aKQQH2ZXTL9NpUCTYOtbFSy
Hlnkx0Me4VMP+g+ZApDefx6nbja37fbm9BNKNHgjXI2xg8NKUQbrX6UtEpK4zzIE
2ujfl3SrE4ZODLf/6gzQZHG3GzCaEgxnTTXgqQBZCroud2gTR/pnH1P04eJX/s/P
/nqDg9cbM6PQBwoSF/tJAnXSco+ekyEO6CBvaqbFx4iYGaaj076gAXKYsgmPvZbX
CjqYZnhZUW62YfvROTozJIXndL1X8BQm82PEjlTgF69+lvVRQO3Dn0qMu5REPF7c
8sRrgLjUfmXfHCh2EJuXVjMZQKu5dIg5CfmPo0Mned4v1CBsB/+YbjwF0VkwfPUN
SIaNaL6oigMhQOKJOaDuVbo0Ueib7Ds+uq7gHvYFzoQhcnPn8ClF3wVy4VTyu7a2
Fnzcw4/2csWsD1sJOFxZI2PEZCrzzBxnFgLSEa1YnTV3FDcJ4QAgNiO+bq3HtlB9
T7Lam2CzLq0r17C1tu/Oc+i47n/PzeGHb9aIzVAsDh+G4Ec2MWPYCB/jt0jCqzx6
B5ThVy4B9/wB3URmSjLl91xdt9OUl17bYtGzqaS86d3ZqDj+IuYt98ML7BUGppT1
FoFTQktsSFcSOX3mwajjsRPyecPbOvjuIOXRlJU4MEEK84/U/aYeZb2ErsoLyxI8
xdSGvYslZNvgafgHfsm04YghbTcjrqwA09mhzW89Fd4ADMCiDNeLKLH8VVN4udE5
0KaiGC4CnW8AbfU4HC5p1A4UhfjjcLJEOHmUYQje4c2rEKPw4BlJg1Mq2MXGurpi
qUB2ud73Fuu53t/u4PwRdmoNJbzgFrbKSrdYvY1ylW6i6P8KVrr6/jMOsX7W/IDx
G2HYe0Qhz8lvtGaBygelKn+SODRceztA3xQ7eHV4khxVBAb3+OO04VpH4LbPUS4k
f+ORJp6nsixcG78OV2xCLM56MTKbAYYF0zkFvqsi1nsgaQrr7mirl7u0KLmI/1ae
1PTYyiv/B6EtkC9ZLHMmwWD+382SbwxGQEQ88NSK28ZZp6x9ggexS5/THK3wscZq
OKXf4alCVdP/YZ3lBexqzLWg4vb16ntzIBxFsog/JSG9jUYyPg3csmmz4AwePzVY
RxNsgkeO0RwQ5oAjtSCqISt9TUSW9gEowFhfAahV4Ijf7TeZMoeTy9EZ/bJsVPu/
ThhqcaLmn1Hbv7KNo0j/24QjkUwQNfkzMBvDd2k2XblKOJ8GcL3WlFad12uG4DJb
ZFDSv4z91T9EN+zDFgZzqI82p0BU8k1dUYk30X3h0Tat+T7oWYMrPZ9jy25LJN06
jL4tdv7qD75Wy+XmnUhW8DLzjLfsgG2ySyNZE0AKV8t4OUGHO9+ayBinIMHfjaVv
tVhEIFf37uHraMWlHefEKFDMjiwZWWeJGgE+ltek2IAIDlnLmDuYwGpS18eiDOyW
U8haUdDY86kMolhm7/R1R58+9qIst4uD50SS8sFc/Hw463GSbzH0sM1x5z17y6Ay
BYvqXq0jRHHoD504PDzPcebyM1OHHRqQA3gTXLQVzfXPcYMWBVJSh4G5Y1ri7MXE
B65oLUsK2DTveoRv1RJ+K2onZEMdiAFncwcSW6DR+OfzJ4bhw3h/ImKlOG4nqbem
4UDOoRV8kfZMwQZVkatEOR10IDwQ3GbrrY/jR2EyCdcTOvhD2YnuRA0ngPhAhFp+
VIRUZlLVoyWv6U9l5HBWhRQlxcY0NJQtAJUS0k4lHI7XXGHYBOuygy7Uh/XCsaOR
M/y1IKO2QHjcvE5Fm/FcqpCkA7+Unf/CuQVimbgbmPLB3PW2z3jg4FBeJgWiLQfi
/0n6gGqp96g3ZLpJb9SAuCcvYu48fq/b2S2E60MSZS6TdzYmscMVXVTaYfHBYY4I
sGVRuLZiBA1l2Atk4zjhJblg2g2ZcseRFgK4TBn8naHWfnhiqCOSlcTeEufq3LGD
TvJDgxkXuXGqf/LJuoytuMxKna32WSgvQPXWiP3MrZBgsWhv6izAmagqWpHNpMBT
VSmvgfmXZ/sPZemlPdS19lQrCGyBebzj+BxU2A7JgPIc+MYt+X3YyBVkQamLWGdr
ShgIFgdMRPD+dIlChq+90Lg24FywFtcdnOb7kEbM6a9xBv9evJaOhNmyNKBm4Oft
vllDdZiuBhWRIkf4BqGSOjPCOUxT/aTGMn73ksBVHXUSdq66Dn/YSL26oGK3jRcv
pa5VepgRy6LDXqpwoOVWRxfAg8/yKn3dffPNXA0Al77G5DAX9o95txR/hqMUTRJw
18hdMjZvAWhfjqINnvxzhdD06BsNRR++42gDOrdHxxf9m1ujznX/Dk9twJZPuHSJ
3/Udx/DtrPQivhF0f2ME5KewIGqGnD9BWf1au7gQ40Jkc0Su7clXdi0oBAdEr0wB
WvVySDrTT7+NKwxbbVh1rHxrIUbWwDCh5qCNXIOVW7WYtauGaJh5+ECVptt1VoPY
XxOt1Ggc6vuVC/iOf/hvAZIDzaV/ubJria/XM6KJ+XgZbTiv4HuYRgmdioGtMk/F
JbCV3jNvRxLP7jTX3PhUnlS0O15qQSpuIsxMpySf14/lbyVO9sFJZkG9H62+qZ0Y
AvTMdxipVKiYuia1NgX6n9L5eMBrE1lqFoPXv4V3xJpjMBOhfe35piV6dWw8Qg7w
1rfw0Ay8F7RCp1laPmETTT80CKJ63TquIxoP0MeG0Z5HjB3O3hysiSMjHH9mkd/Y
p03/GS5w5C9oWHy19LwC6N2esMJjKdmSReM86uUMHvcAxljVj8gOlVFetIxV+tUV
Z3US/Ztx2UTkKs38tfZVj6nUy/H3B8owW6wfoe3S9HxpKg92ro8VM8guaMdHaKxf
c6pRcTIC/J9bMXwX1L+pwPKi/US3WAJqE2pv+kOHo+BaAYpLhHBIBLNBkPOAw+Wi
U757KthmvRd+KqBXYkwCXF9UNwMwtkcomNyLD54kEemcaWg+VQdajgR/SY82Iki1
wyaWdbxvlGrucwRxRPrCZZcOu1liU6fpKa799NezPaMPpVJWFmUD3GkVaVAOeSOB
76vmOTq5rKiJr+E0tNsyz+KvhUJUKew1AoqptU6diR6fXaKMG++WPr5wLM34mNiq
gMlgpFgj0VmX89F5bDaI5Dko65MxTte378Jxbd1w17UhC+V5wYuo82kHs8RSsftq
O5s9VsE/gE3+8N4kzcZzrKOIwx8xNQwZr500kaWjDfFSRndqnbEscDyTHANSjSbu
h3qDP0T0x5NZMfD5k9J1/TZNgvA3MOAc+t+7bV6rXOUb15hF0pAhGsRDVaDCvopa
0Hssmf/hlPXr/7MRcfJvRfpIIGYSX7zVGw1TfYH4Jg1HNO67qeZGOyCSFiPp2P+L
9KyHrhtsQ9bzYpf2svhr8OVw74MwZUJ/C8rw1oO+KxsM8iSJ2IcrNBeNfx4lsl8D
NM447W6bbVCiSOpEoCKR5f0xiJOiCc/o6Br3CGMdjZfsv4k04MXa72fOo9qn2Sk3
tAzrPxqHmFwxUyqMZv1Yf6/6ZvrpJ9TOWbCdTxav1OxFEX2tJ7FnbvskD7lF4lF8
tF4tCzoBXQMA+GZaDgoSIffZPgBThnfuDl61TWZO+18mOMdUiVaaknoZblbgI/oR
/Fn6PaPlUCF7yOwylHfKgSyIqTgfmB0Ad2HOHWGI5i1YuqUFF2T8pyfbdu6anRvs
T9lA9bh+PdwxrzTXcdbqNBxug3Einv2UDWbCMrn9D99YgY1cVn32kxrQ8WScpvVY
swR9EETJAeCI3BsWAV6JpyhUZxMEJ22Pdagduz1VkKoZ/8ESIslC284ncR2QbAKR
tU8yL4q9uafMCdGfO9gBm42ld9UcVYLnb1a95sBYyDgZiJ6MMl/u4C1GvnXKdk6e
yp5vKb92LfYXpzXJlpFELysppj4vDkCOO9zdyeWVV3J8JKMzRnsNwjCNJ9MgRv7B
e6f8jxXhg0cUOCDvX/BSAwLx36U5uPgM/PrCg87fVMee89P1Zj17srM22gFZ9wMa
w/+Q8TlPPQCTfeUWmgBQ2ncsYCvF3bzxi9QKsb9TgdBgKVIhUs5+xz8+1GeHh/9j
2mDN8nT+iwKI2r2LE1ZLH3z0lH3aRq33JtmERsTB1ZYOQcxfmu8OeOKpbBZ5tXw9
oinD2RZOCaGbrgzABbF201X6U0nTXpeIEO5rr/gN7tYKFYE9vQ0MirdsbJg8JBdR
STKo6CT0s4S3a1Pc8t4wjgkifBYw+nfaXmSGSB7RsT/pKNEBoVQEWrrAb0uX8FUt
DuaepOafzp+Elv2MlmELIJU3JsGSJWSBKj56WDJB9TWYMvU0GW8Xld0h3x7pYNtq
A1bjs1U9tmGRkbDcDmVgpy0915mzntv5RChqnAn5f3Tg/fcd36HCJ1RiRwIPUwf+
XyXYUDCkAtLlEDyBuCMDTt86ba7YKub5aiM3+PN6R0Gxc0Vm4BjsvNN3iTatqh6a
Nl65eeKXUkOl5la5INdUfhsa+reslH+bjWf6FKC/JZf3h7DWSOLG0ScHmsmQ6USL
VGRBaNrQ6kPj+9ETkALGk/GLGKvy7J8KSJHIprdUB3uC2i5iipiKZ7B/1A0YvH0u
et35yXcT+B1l03toZJeFRAubX+i9KMcXAqrQgGCCQfNUUTLuAAuKCYw7+bIze3Qa
Wj4Ic7SqmihCwQKcKmwmEQsvApm7FB/2ALBuvf1wHF3xxtaKydW2jvafJPORGX8W
291Bg2YaKZQ1U2VeGoaNpeLh19yHB0YRbD+ePs93+UL05LE/EhmuBk4GZ6u1LkSY
+cYELn3V5A0kyaoZRThnqs2lVoaQQd86TeBcA+t17skgUjZva6EDi8pgUA4/tQfs
tK5r/yLwSWiQc8dtIMpzTiAjMJI527DhMA+yeyO1YgBOxiYWhApkK+3rHQst8z0E
fAB56GfKH9/a5UdkJED0KxWA8+zVKReIIb1gVp6tideq8g2mH0s18GYoZgm8VcGQ
yvNTEMjVsG5boGIXqKrssA67T3L7DhFbdY/ASfoXqiXE6OeRouBVrTCJZWqJ+nd+
AZGMvd4/0tOO15jwrV0Y4/mnZRW/2ka62wyA3QNODw6DJRadkVdnh1KSKEupjLGk
J+ACkIltmup3V8aDgjwmBIGjovO71v85BeYi+pth/CdT/Npu/nKtLdTeB5SUIC/S
XBu89OWg7GczcVNpj5hdbybDak2KT1kmOIYcEJ61awZt6Wk+H7P28LLUqdknLXip
LclGfPu34/PLNEdIroHeM4FNz0ThRjWIQ4fyZMqwPmc+qQUhgHFL4l9IICzw1jgb
CSmIN+FXJYPhGs0TILEYgFJypFzplV/cuaq65Wp3v3MCVMvg3seWNFQ6/NnXyuyj
qZj+rZudfzYwIIpD/hfzRnxwsry1OvPuUF8ZqmkqsVjmgYzUvPj8Vryf3ZkkKBZy
MfwW8XnEo0uvpN/3gk96zJYRqJLfxslR6jgaGSdKzVZWLoP0IVDbQ7XgUbXIg5ta
oEc5LpWd75fZVP0z+LGj/9BxKATdQ5oFEBTDjNQ/OUedWAi3lvuAAEc+HciVDpLa
0QboMoPRHMQgMZm9+km+TMWMtaaTcPLSIACliQ0mGFT0yjQ7/ZqLyc74ovrpF3+H
JnIiKKFDaUrQQz5PD+AmXMxa2VuQ0nau2of5V4b8jCGqiiSM0F6ZbaTuFlbA5sH3
ZVz68yEe9ZvYNTI8Mi5uXJ0N7A6i23GPFvu1Kx/8jKpyWqgkqJkhYOgzrz17/l1I
/qLmPtKt9sxJjjsEOhzwaKOIMu2PklUAjlrIs/kLCI/vsnRUDlQQmAlgjL3XXR48
Qkj0y0EoVfRfUql0N8Tyvmz61FwsvXndOBfW5E7CiUmy+MwOeHFd52VMwT1muCiP
qdcLUI+JEDaUxWK8/N/q32QGvyW67PqlYM64iWiDJT8YMnn28NQ9BRCcFy58ci2i
uSAqkbxux59L5UiMkBa4lEY+/pLVLpxYIvKKuTsatQkvNby6r9T2Hr+5Vu1PJRxA
BkAeVEU8pFE29rIeJfhRMAn8jsnAVliAzReI9owOWlmLMeFr7eh87WX2ewcNhc8l
N6HhQc4dQsIbgljWb4TIQVyQLHsg4htdA7aQjye4SEoe+SVcN47++rKA1CH+q2er
ATNY4QZyS8TTRuwJ2tVHn/4qkS83fXHX1Av3ls0cywx1TQoKXcMR2JQoUBwQfKmh
UzvhFA/M1rQKvo1qQdSkbTOeagrTzibeFhOuJ075t4cYjhV5Bvhfv3DW3YtNuZ5Z
u9b4NhzRJ21a3DdH632wrDKCp9deovqMFx6zgbVML+NToiV939cZh2KvBFRAO2az
S6bd5pnxFmsrnQgN4+pHUx462p6ERlPmw8CatCaMJTJgsr40CNERmdjZWGMiEZgh
mY1w6MN1ckBqaoIfNK62OzfkJWhyHUgy1ZglPOxxinSPCa62hhI7GIiy6uv/TqE0
znmp1oPA9WX/q+4uJRDiEDZayVfH7aVY9Zg24QiOATntHQJC1ig78uAOG3u9otZ2
R60XXLSxodQjVlVAt5WvT8PTVLnNuiJLiSqL87OlnmDNtKyZqXRpHpK+/6mca1Vj
U/ZZWy6pvOXHxd4vIadMfLSXQ2Q0Cj+Df4579cJs/d2SX7RglpJYbFe4kkH5tHjp
F7Xagpp8ibaUXawwDo6aSsVdVvMtBc25Tt24AB6+5tgWkaeTzWbVDNgdmwFdHDSh
nZBI1pG7Uvs2Bsdez13Zw30p2cw6XDhRB2Zm0kosbRwWc/Ko2wdqmvrCmO6P9Odw
qaGBMBjIHVrnx54t1KKkXQlBgn0G+XzB4SuwxnlNHFAn+/SswndL/LAvfF99vhgG
gYE0UOfQWVt98W1eU5s9dUTpNRYgzRoeOaJpXNLPlFKxY/wvFJAED1D3JAoB0Sbi
BWmesnBrcY9e4ls0mzQkLPts48PfO0V4shgE2wU3wZEaHvExr2H222HrhruYMNTX
J9I3x00w4k0iFvQ4EfI3cKzdCikfsFgtmzwwOLRRaXNc1TcSWoHPy28MYrJcbD2z
JV8KRn1xWkpunFdvpjN22ETGVATmBZrlYUdtCXwHxU5rs5OUQc7zuX3v0Y8cEiXd
xHXCRaqa+DXKHOVZ17TsuggHTu+Q2zk1vZHcOGFaJIdC7mvW6FAiVw/9nEjpgnJ4
n5OaHE5qEQSm5r9202aZfJzUZ4Mn3Wswo3GV3UWHjgjy5gkxB7TJMSEyKlobVmyu
ErmcnFXjkCaT9cd6oAKDQJdIIrAmxBhyOZtljvgoGvW5zPhiBlTwodfsusfcU1qG
6ljeno9B1QPDRfvja+nWMyz6AVKGi2hJpHrc73/BVnVFSyos4Es7pO0D99baFd5d
ZrDKWgQKZWh7P7czWnlwgGtWwVEVyUdBMrr8uQiH5lVabiBIl7aFfysj6iTkLvvp
OMhRxJ+RqGxBmb1XDtOBEpsOYiE+V2K5ptHzrvIXTkQtw4tMBmxRKtHDsScyInLX
r0XvioaVoaMux3NCfaVRz3nBdb8mhkTfDKaXJBFYrMhCg1yPayZZm+J+Piad9Usk
i4MXF8xU37sSHUObLfTRgueIlhEwf6lDemQyGw7YrHEOlMvi5ZaFyqhK2k8VHgBL
7VfmemVpB0xbWmE8mw7f9KIq8fIi+cufYOr++i/NdHrp0+Z198Lx7ZuTv5TzDZJL
zU3Rqq2fiRSmGL1VsHbrH/25AKKGy2uH8tt9bd1RNM2y9Ikl8ihmLfnZ3BLtEpZi
SCoZ7612Qfv42zv6j+t2e+JH6CkWn+tL++R6AOQewM6kdv2UUvxWHXc5NLZZehjL
PdPIhyLoHicki1E/GBwMMwGzztj6GI+8a5BuoshSmUVchEo4M4UmImuhljR4Rfzu
NQu1w+nvTZHqby8P/pSRCB+0SzXzmbaraQNevSwDW4o5QE6pFfZ09hZ//ypzuQU4
DiPdzxy6g2FKasr00MgKguRmyGBUYzXHoiFoHJjHXlSYJS2dRpSgeBha+G8sM3BE
m+YJQsrbMfEnRDbaqoLXjq0Jqbz9P+GipP02qNIEE0wal5CrmgYQ+lmgA7K6GuIo
QCsEqtGNA3fYgaqfy5jAc4zlmqU1ES3IDUNxFuKV+Xr5YKU7+C5Ss2Lwd1/jx/Vk
qwMwNukXBBjlgyuCTuj9HzlbqXo6fGKovcZqjE9Rt5fhlOaYdUl3DPGLrXSVw0cU
Z7QswEBDG1x61NVC3EL4SMzOO+zOc6GA27yY1CtkBI+dxc6zWorg/r1KxHTLuDj5
zmZKnwI2oiw1RxwAP8any8nJlkc8pH+AxUNE0GKD8j9S6zOUmbVqMPE5ngpC5YcP
ST46fbZQU8cnL1NWsz7YYazVJqO2aYPMN/gOEc3/iSJYwV3KvHIBnJE1t8RPOhOt
n2J8ed1g3J2S0vR4Amq4asU28oSWLEl2PLLYhO2To7u5uPKDNhi8nabMwZtmHcyS
MVz5tVsoh9Zq8vQMVZWIiupj8qSvkiVhkMC0wC8bnww4ckB/nz5Ff1cnv/wUyOuK
XjEBQaWT6jAW7Qrbc0qi2edyyUTSmviKArbEyJFG0V8iOpY5GcPuiYsUzGQXHRQs
wc9PotU8XxvdVDY2TgiHqbozU262j5TOlhzE9qSACVeBI+FR/jbgHLu1pP37nVum
vwKyBWHVXzfrTxtd9tSLRROHgVcHsk9HJs13KpAu/LT/L5Hu2z/g3t6FtApzX77x
V7KxGhAF3nKtf0fwrKbotDsmd9DP1ySNGFdVOHgb0Lw/8WwJByH+mBM6k8w5FRuh
zEgfX7E2jcLDV3mfPnrzugV40yG0konqwn+gsjkXWLSmZM5lttACAwx0g1q9nrTE
6RUYcQyKVerkCR+FFcADIr8LPhDXHLsyW0qeH4dnJIJ8j+hVC3FG4ffTJWa8A31V
R4ALx2qmlo7ez1deOsbhQcAQ/KxCN4hGMFVm9VDbBxIaWrK1UvElUWY8bas5SiQv
eoGZcGE02f34/o6bgROwlFAbSS8EDF7bD3sezNQiOV2w/HUBkzbjxJ7xag27O4bY
h8nhZc5CKtOYYP9xCI+Y0det7KlYAbwPt26jndiJ7LcXMfr7GbFDPCs9XxZpNrQ2
M8uvOC+VZhrbF0zgEnpjnP4jYXBOFGx5CUgQfPteK82BsF9SKhnxW0isC87fMSU7
DS13Ah+SpY49W8sMUbaj7jl+CfmaBa/keKy85nPZgkLcwUWOOBGLO6RBnwF9xCpf
W1DCmAjLSjN14ACpC7bejHFu8dxDc/UNUM6wbvgfYh2bcuVBSQRG7ljw1ifyLD0B
4tiSXRdgSMK01GhddgkuWWaSXDpvqtT5uMppkZZ/LMEI3iWGvFlRAiK4ceGVI31f
DzJHX8QvLg8nCaT0um7X4ISWl/UCcYp88GslgvB7tj3Iec53FFhC3DBYSRt+Zo0T
VPSkqXm0bikeCNLwoAaHyEZYt1Id+9AnosAsGQywF2r79LujsoQwdRAxWmdvL4lA
yFc8ughg90eieQ7qNeF/O6dRZqGYiQ0TqMwlBXyJsTfCIrIyYA0G1lFmn+7CHk+W
R+wgWZkA+Hy8gf2BSzKcs6tUYkWxalGMGhAq3hzcjNydx5t6WWrrIOQBKHuCd6xt
5DLK2AaO+57JB9RZy2Az1qPY0+e4x4cHJKun38gjaBXx+Jqtolu+NIGAquXWQFbs
Wem9VTmatfaWtexGj1795rIWki3EJhcI2HPmIo48ZnEFrDOuoExk4hfAL69Az5Hd
UUQhaDVyslcI0OFOq7jTj3WcC85ECracEHfWG0IH5pyhmuCY6+HZF9RgA5v4Z4R7
8trtSIdi15tGI746Ndk1oTDtMtuPq9oupFKuZPNPInE5/gf1ypXbSQZdDNQbO2kg
VFiA82fbfx1JW3TbsUv2k+C1lR/X0NpGsqce32X08ouQTLBT9jFs7GEMdYvmQ67A
ThSqrfDQhiKeaMKhXooa1qGn4xbeD8TePvWtawRwSjVQTTPDnL99He6fcLVKY5gQ
LwAHuRehsjo77Xt5J6J9eODTuL0oP4ab0I5/brqSJH/CfLsprxYrbFIYxciQv2iU
qV32xd5vtOwWLDXbGbZ6qW1FQoGFHtxA6aB+/eAUJ07ZCKsDLpqdZ3gr1yL31H2R
GiQXBgFMBK/hWVVpUhYgbwYa0wcn+FizIjHCJiEW3EaLEwGZrW0QNpu9Q/VJ6JYQ
4XphrKkvIvNvwMMeJ3ZTbeWdv0a4RHFGzeztoEPMgUPtSr6L+3gbbsVVxQG38G4I
nGWJamqJRtnqYopsk89yPldUsh/FcY12XyTIbbxPJVGKoroKCed39alV6LJTRQl+
kwqA9ijVnSKJSSgC/HePlBcnjxIPoSeYkl955HW6y3CTo2aEjlyevyRBUZxHFXlj
31yw6SyUGPOuqnJ+hSISIMLQA/fIfSQqMZCizkoKJMBOQjaQZlNYQZj7j3jHjJeN
ibYnfD4aV37p8CPcQE5NJb7eNjeYonK+8YwmlFzddhGqjUG93qtC4bVvGvKxC7Wv
3oG9aOxDUmUxrOUXih49vTm8PwVxffZbL4E3GBpuGdFm2lK2eV0mGQCaz6AvVLph
9+5IMTD6Zk8/KNzcl0zk7sxFhkZ25SxzurW/f2Dj3Bk/s0+TkXfYCucNoBtxhnJz
O1yFZhFNUeiqAK5UXiMwQAoiN1UCJemZLhXvcZKpKjzoSt6aQaqvDwsOpAkEMF58
65m/MJ3gF/hEa6j9Q9s4SSldxZ1lUZSuRpfB92aGeIgA0qtSp66BMfj6UkjiWpfp
vXtIhiiozIcQdxuNBFjvpPDR7MEMY6uMC5ecwZCVikg+lxGoZncucAcApSMFrz02
rPaTaBb4p5AL9TfjM/HA74vtlBBFepASZeqJYEARzfxOcbspbwChpy1LwQfI9Cs/
pC9gJ1IBtiB8yXWOKDTEAJ5anro57VgB1QtJKJ0us4fruOvb6N/IxUbdSk5dIw2+
Y03GgoBObEk1gUBLIleg5K0SE0lHxPcJhQpCjwFPG6in4oX79sflkZHCC8e3tvEM
Jd9H+pyN6WAgavWMjlobjOfwQWvP6+yQ4uCnzFYhNbf96qRudPytvd/3SpMyKKWb
N9g5eyGOtGKNQwj+f57nZPEtUJeq+6lriVrbLQq/x3TICCwqwQV+q+oblOflJX4i
CkVk6kfn7QqNwZErf9Cwsig+0g22WrP2i3R9jctZoCpM7EsYaLGRx7QrMlhE8RUA
dvcG8hFnDwi4i1QkpzNEkuz9fUhVCnT/gCN5gjgaZ7N2J/Nb4zEwfTyB2vpSsykz
CNoulskpKq160Lu56cYbCqfPjg+CiGRm0NsZh4cymqjPYXsMu6+vD4XVAcl2RN4N
i+H4lB8e9tStwsRZZifyOMMnkgnyF+sS4n9lBzKukck+qEZopQ6UAsjGlvXqjp96
qWRlf9cYnrnMzYdHwTx3an2kjWR3r1CQewlBFjH1Ms42lID3CLHPlw1w6XJIJX9p
1IXEXJ7jNoOa1h0UkAvemezodoazMP4vFmjDREinAuKnYm3k1v74qWows5nifID5
MU30w6pgj2G/nsu6MPTZQAX6V6Mmri97CcEmkVy98N2YOY0J5dtmpb+0r2aK4zHj
1D/oFnIk8+OQ5iT2RZSZcw1TOPr6nSEVYisezjHt46v/1Nig4mIffDkFmv0xrlsh
QKUM1cn7RHaNVcuUY+kfToqb/8Pq5pvN8tFbcgu67ovA1RZbtDGAN4GG/6bMof5v
gTs0Qqs+AqDR4hZu8fldjCHjDdGd/bZaogNDr9W789xa4KWN0yx16SyNe5cq4MOs
8m1o3UzPgfVQfsWFcts5W3GQKvVxrpcMxtMMayK5NL1lNxHiWcPFrKexokPtgyNo
qaAajLxTOUN/YIutAI9ZhLquYVxqS4mEPV+OCO1Zhg6uMVS8HFcCouB9SC/qpRHq
1q5M4IEaA1j6GOxCYST1nHkFBO6lhQxy4EeVafPNa/i2Nimu8UPtde4ML0Q7fic8
VZtvuwZEb0YL2gKNjj+o94gy0ql9GZq+1Zz46h1CIn1yGvDFc2CffJwQyZ3Ab4SB
1iwfiLUx1PNVOuzjlNwoau0RWCF/s7n5tuYiqnVPVczrr/FXx3jCWFjAeCFZ2S8V
1P5bP30PoB2+HLamSizsCqyXvUDkz7n7/FkmeonLf2vE7kOaysBihyAk4wSpi1dO
ltomj0O5p2AmV3X0g/SbRtyJZ0ZeBGif1aeJWYhWQwbWI44oiNazHYQ2EdAuKLDl
k4f379Gl6jJhABmqhoZ6b4xdAqox2OxYSshzXY2hm7EgYzSt6EKOzAsxPNfO0sTG
+iHH9cNZebl3qFKnNF/TJxoHSUJ+ECZZHT+UEOS/Hfpw+yYDfCPPqUl83QGSz2lq
YLDApXde3TrZAYhkqJJY01S6+F9rHGw9/6Iq6wRuMxuHPLAo1GEaZy3UTHXPFqkJ
Im44KLs9P2gsGH7vGEx7MAWm4V6bDX46PY4vNX3NnQ8mgZ6X02R2CflF5iDQcHtf
XG5/grf2O4t9xpV/aE1g678lZHu1CJqjX0imaKI7W0RDuoXbNU5F3imGdm42V8YF
e6R7X0JAD6g2/Z3Y95IK2CQHIK4lNJWNigHdKYyUPQmXCxqPkgAq4/0lq9JBdE2n
Hn/GAgLA4Fbszn+D2Z4ioXxvjZaq+1B3mlMXbEUZiofZEacDQK3JkmlWEbxj+oti
pAUdCObABDml0qq/uvfNS2vFhtKr9c996+1DrYEpIVyQfxkofz8GJtrqEcn7Xh2o
x8Q9lLXwA++5CUAIbFD4cptKNSM87HhtF3wpAt5sOa0wP+K0Q8EvWfztQa97Gw9x
3nVvyHGv24BXJdvKNYuYf43JKX2WikieRAtOGpLRcK3YWw+ZEFcAbZg8YYtR080L
5XLrQBED2GM9qMdLdweLaIsH0BxEM/pjGEgE6pL69YBDicDam8Ytj8aHWnnFlQkX
NdFdPUASvVJtdp9ewAuoouibe1NkuQ5wOeeWyFHfcPF6YrzodUZLUJoYw2oKRotf
YZue3dMMnOBOjpbJDPH/ymummrjyBjaGZi5Jd9HvPtJGKuEze0iO62nsqaDEWvkn
jMHijDXHIzo8FBn7FNA97hPwffBJ3dt9YniBP4uXe1oZutj2SuTVpXpDPKYs0gJg
rZ0zt8X8wsA6Ip+kOs92JVGjR7JfC5cKxxR6OYXcS4I4DebJ3SJK+VF7jV8f7/9f
ErMdVXJeQ1c6xIm0516bJyTXqEZ4jzmbN0JDQ/+c7BIJfMm62Qgfsf4bJ9DYrgMe
Jh4vWxCAoIHsMZejt6g/QXDh8sFeAnCcnGHMPB7W1vPMM00WCrhfaKtV7ulCLJtH
IZi7ec2IFdiXWhTEJl80VAcR3hT+vqEJyqq4PadQaykqvObUzk0nrm6afqMH2IT7
Uz83IBtnI5efVqunC1wC3t4FhQ500yRSaC4VzXVza1DTb2XhwCtUZRRzL60b2G/H
ikmUq7L4m1y6m7h909zfB9nfjt9gatWuK5A/+D6DuKA9ZO18SOknur+07otTG4AS
BQFvaGKMu2j9xpYtZRpQ5Hgow1uvO5ocGPuQEluUwEapeYELl4ZKg0G52r0pUTuv
3X4V7ejCgWM74a36m0rYTO3BpAs3DDJZ+F1zXhMZOKmQ5/w44NKkIwikGRG5M90U
KLnIyvRVyNKyyx0GDtszS0pyhU0np3+NP3iAsgzdQBe1efkFunTnKimFeDfxNbNZ
fKAhvDjBW4/po42eYKQSKR7Sr75eIZoPvPq7NDBo3j4h4yuZ75efOs4I87wp8XLE
yRkDVCxGsqvFCD0+/qFWCwKWzX8g5Z5uNmFTUH3rrhn5PTx3Pp7kUuhgcFfCCVHk
mwWmESlp+tsRBQYpPXj+lrFhU1x4YLoj5o24Ey7XnWdGQaENWtlgsl/2eWThu9oH
6v7jL+qQr6rI+UsNzqotXpinFfX9puWvA48MIjNk4RNmPZBp13XqNe/0W2yN3HTk
Oz06nNJTSiGJ2Zioq1lPglv22P8WEvKVE8pzxNxa96PubpOzzBCd7vsaMWuD+WOn
+a8KlyWgqqydd4P97Qyt25AlY33Lrx5ValmahEtJM1RXej+ymHxr9xnFoHEh8pnZ
AugiYuN7dMZEmRZNMSfQoTBgXSu0f3dZJD+ioWMsDs5N0QXdAekZfNV/Jgdt+05s
uVR/lG/XKYCLinQstid5R8UhHcbhc8gf+XryWqM+V9aIg4IcgDy9Ra2esawiGfrN
WU1dAdeRlQ0ObgOA+501FAJGxCxNlFnbVl7usS/hMIFtSk+ngXw3KQfO24bDxdk7
TekXJ78FJqeODr8JOMBLX3aHPICuCtDUbYbvN4pqHIi8cMIS2kvDDpfx6Lvgd9H0
+f3feH2wKLPwqziZipgu6H+UYCL7DgAz+u2Y+jrp0lPDpsFG1rqGjfZlwrP3uvjC
T/OSa1/nzwnxAdFtgPqKkWWgsH6KAPYvNx8Sge+5EzOxrZf+HikDyz2GHOD+ViW1
A6ygyhr4ZO3EMLaVd/o+urWtt+0QVB3Jlqmyw0yaHk0V2Hs+KLwCXzRzmXai+vNB
c0QNHX2+9MsREgvFfM/JKpN+CpSogVYrnQUFXEPyCnwUUrHhs0Jb3m6/vpCFUyPD
kPKxAF/Qy4jIYj6mHXl0dl+jFnOIZuJCzACmo5MP0puruYB8z6q/eCfRQEtB5TXX
FIEkdDfg1HS1ku3jAOyfYp0ZNZGEbVSs8ZhKcbd/GiNqCUg/N6BJ9viZD6hNQRJ0
WtYaYRiwX4F1KG+zhrAZSPDfStqYWXvOeVNRTjuccfP9DerTpJGSZhLMZa86cj34
nVw2bdhtORDxeiL4yXY40vn4UV9wpGCzQi4+UA6YkOlfZ4RyoIvqo5mMQEms2oOK
lHBMeSgSd7wNBLjfZecVeC4d/daruwYGVZ1WC5nNYXUguf3rm6SCuE/5ryP1de8J
RgWwiKV6nxcnDazPkooJPJp4DLW0fg1k1s5j2InpN6GvJ+bknqjylo4S5eRbHqNZ
Sd/ofNFHPJxko/HNRacWbBPFiqfGQAvry5ey7pzkCZVABhQJwpXvmCeXoB2F0IYw
iX66ugKWh2CmQw4VFnTC/dqtANMkgAil2+cTL+UcHVQ4+tEKllKX0C5oRrYjhWk2
lsm2dQZYkiMf/GeP/RVNNibN5cDWUFBEfmyIlZSx3zpB6GPlx7PKToI8cSAPewK/
g1SMqC/pz4x77emk7MAdwRfMJ5B4KYDVUZU/AWtHmtx0zcCi5qkJ4/OHFw5YFihv
6SDZYBVcykHx3plqT4P1AP1QzfORNwbXmjtHVkREs6BcaBW6h/JfpyJy0L9wfZL7
HrNlE3S1f5gMDf4jwszldkVsm49APGYP/b0aLdTV3BL9W8IOJ1RdTlZlf3iHv51E
BaP2Xpw4jGyeYee89UH2UyVRiPWtj68jFLhkseOxHyrIrBzBCLgwHtRLy9cCtsHa
RZVqAvbXIauLaZBgg7dAEki4QegjWxWV6Ztb9wvNBRsTE9p8NUbsh/ba2RxLPfag
bbWeKZEPXETdMu1ZbGKU5pr/fht/norv9XzMrlZQCPe9LqxFyHf03bfRq0RTkf1n
W+1l+FEuG/6tsfj7Voq7PbA24lGFoiUQCImEp4JwShDusS2Ptbdai204W8FdqH6H
pID320L7A4/mTQ0PvpRRr3Sr1yodAbc3gQRx66D/TOIfOCvuRIDRfLpRQ579eoJk
VSFwjeZtd2ZZmFwVIb2WXwDYG0lQ01lPtoDTN9Qs8xSTKlVCARp1XodXCo2Pgjlf
kyeePfY63nz7+QV0hmJO8cjdme986hzeVvDCcLupLnsu66JGoLPx/9+5DCDYP+B6
QQDXI4t6/KwMyqroxOYCX+ACC1v9ej/p3VrYSh+DIf6Uc92/XRBXjjP01Z8CzuBb
g4qMmuMgPdUFyCZLPzKOh7+4EWbOF7SogvDnLmNlBXeQoCh/9P6q0jqeWn25w/35
L7XJUxeOv4IYvTaqmdOQ179tXBpR7My8FCwTvWsbF2C5LDgKEaXQdrtN8F7aovUF
P3EWSp6tcAIQjDb46uU70XMqIkaFN1y5nkIOeB0ttVBlzKXv6ctPCiwISu+qac37
2spm/0vEQ44qXaxHb5kcO25y9KxH+BDvWGZGv7lRbK1BmLyDmMKuU19jGYgoD3A5
1YjF8nyH03zSBgqEtnAeSdKYTcqYY7h9+ozFmuqCjMpn2Gz58b1Za5D0/fiD6ixN
6UM6DeMqDDY7FEFrOXOkqDQmii3BY+5TelVDyAWigARjoUQmHL39T9kOaT/+jUzk
KdW+Bnh4UlpXxejtFr/acbRgB+cqB6Yc1jDTNgzeOBKDf+bIOQtbYb0PuXMCiqRs
EH2RYpbtimd1/fZK4cH0h+YTWmt5FFFANSYfmfoOTgFXBOaVCcYsrkPScwcA7wwf
ZU3/3NjxSgAqlo9kR5KHVcLH/9zcYfKzPDg2t1Vpa0xq8z55nbkS+LqkMaBFIejK
uPGt+uTD+z1f1jNJT1u5sb28VInUwPIcfgs2JgxaUaT7JWdgz1Y9NEPxm2hdp5Ky
soDQxItauh2FkW12PW4JD1MLe3GbraAB/x1hvhekmBdsW/eZnkS9HTaXCAdeDgDw
0IAl/HMQV968RlBftpHNO2uhxYAoIl7R5bzKHzD9opuZqx8annAvlYh0cxS7wjlJ
EhMOb477hO62rB6Y+D47C/92Upo8S6lWNUW+iPLvvQUh7rTX57WLn7GjTWC+nrp/
LQ/NVX24aSDpJacDKTcyPXCEXCluGURviRWZgnVbMQbf/OH4aqpGYBfrRMa00au3
tj8H/nMzWYlZnuY7g7CZb+N/TNh1MAEtq7pjMap6jVtyjHPrsq8KYjBMjOBnICf4
n2wDNyg14q01iT3u/DTCOFHtNE63qrtrFW+sfEOLXCnxXp5uGkSNlwRfhq+8Jmlz
S4Qhrl8rcX5j/BOjVieq+u19BWOhXpo364YS/ZJwZeYJB0wMvxXMZZInvvDyPbyf
OPwpoDYcUoOL819k+KbIW3ZkmfWsRdM1nfBg9iSMIEGDZ7iqLuD3luFnZGALEcXm
BP7p4hSLaC4ZUZ3sF2CAxrsQ5Ly2n4F5NvLgmoe6Uu/1Nms1+Z4uCWttVewHaEKt
taGR//Y3fPP58QcCR/LrYn5mjuPTH7crTPVHqKDiXxbia5qRzGnft9f6iL9Oidd1
0mLUMmY/Q0Bh/bHI4vD/JRJ677f2XETaWPzr1qZJJWSPmlHov1wcx6yudSvOhtMb
0bY12yxp9TpUwJbv7S38/BcV+LN7xkfDmOKD0C8QvAn9X1kJjR9xoF/EEm16M9NA
Io5WqgjbcoyOzK2dfNJLBUvx62BK7NjBazYXZzrSKrV+kQfa/kp/B1aAry/ztCn3
H0d2uN07SsPIBDBJ1VeqPO+KZ5H4SS/l6Jwop3EqjdfD5u9InF8ipyWWMbNVf+t8
dL3XFScXFTRJnE9aaxHxn0XYw3zNYeYfb5a0kFGlFCCR1Fje0yEQnd8y8YSAcc0C
JIohpfafcqor8gItjtnf6gQXtn/IT5pIi9PsX1bERVFpa/pmKp/5PVUl6oqIbsOR
JXvfw13XXFrz9/5TjC22Twc04BVKzxtRoPY+e0bejHq/ig/K9Y1wRvsIh1VR2x3V
lV6bEr4uncuzLOBTb5G2JkRuTVUt6zi5UlJ2QdsSX7JvKXhDK2Lq7vnNXWnEHxX0
tkzXmzJ8ivroZsN7g3J51QuDj2Glvi9G+1lfS/H0Gx1icI8EHrXSNkTP97aIiJ+i
DUSaltab4r5FM0amzq2ErAZBuHJ8olK8PL2kysWP84FvV2Z4HQT1D1jbg3uwIWAk
XkrY5iSw0zoOxAxR8PR3gvM3BSHMsSRJ/hDNd5Le5xwxTgwRHuaG9UFk8U5sXB2X
PbFwThodB74mYu/g9dZZw+5qye78QxXzNn256E0BnZ9ALZMDHzzLOlrBxd4iaxs3
Vcdr3Iq9THr9KyGlbpwW82LF/PuX7jgz9FAA09krWoHAa1KOW9uRUe1+doPtya5Z
0c2C+CC/5UcTk1SMP3P5ydkcM4qdmVvEQbuB/KToY0IJBeB6Zxdt3esnSMDfswNi
qZ1gmDq9no4Lsa1Wc6WfLiMTRic7U4hYM9numQJVG38QfOV0lpVnN2vU5lBM6gJe
rWzwXYPt2a/D0ovrcs2kYxfCKOGxWrPI3U80wCGDMtqQr7abpEeuExNpGpOn/p/v
tV6bX9IUFNoP7zJ5LW+hZPVkXsrJB/Qqhvt7KPtr7DLB4F9AamqEq5SgvOviLPrZ
ES8PWq+2/v5SC3dIMqKxZ7YEh/bX0ngOQzvicy71lOqdzlHC0bS6mb7kkuVaYoU0
WedFfrSG83/ts72XxZ3miAnPY6MBS1/5J9b0wfnKyXRlV7GAZdYDzdJHW3qWMapJ
BnmLR/nZSe8MaeDt9/fyWvr9ViVIDhxK8ufyijtFlUkELpRCyoFZCbc1AH3d30Hd
L4Zen89J6AyG0THX/ccyHS/yBGXARl1zMKea2xm0spcIBez4xLrC6lSdGt8UXVDG
FQJBl/rVLpGRtLO5dAp4EJPY/UbiG6vUEqf2c6mXoj3QxWvlep3dgB4mxvd3PRsq
0gbj09921x/uN92QgenVjLdjxu72fapnRJwP9HqGwH9s4ByrtbSZ1Q56YJKwDJKn
ZlU7wL3WdqzOxZhXtabsWHTo6JigIbBkDcZkOzxmsaf4YyC1cKV6yVUk/SZPGkEc
oxDjn3VUSb4mSbNcLJKtqbo7g0VUtXAKGkVHx9lOZVsDX04zyE+74l5yyXHzPd6I
f670dOeFVwDT+Ti6DiMwP+K5NoofTrsrltwYSa/CHx5Ut4XyvlK9nLqRVChzxEEg
Ard7nbedhDbCAeq3HN/FplaELraUxeJvyNrOe84mN7fSX5DYOxPsxvEjgbcH+/on
yO4Pj1/xodaOx45a1RDgMrl2MBl5sLUyDJaSVOwD5GDO72RXsdJdwcKSJ+ek/Uf7
hemvTHRnPijfwhcj0ayiGysIA6hGLGluJjpV1ZHaeKk/C9tNGwlmFjMwOSMLOn1x
2cnnr4GRkEf2OWwoaFlgbo0bCt44xjIHR8og55T+5k8In+5fYys2x+eslKs4+GMX
jSKt0sC6zjQI95PaIf6V+OYlJgjhnDFeQnXRpA/mhVYcS93kS7X3jqXkATZAeYLg
I2a7LTkHPKaQqXOiaWLe0iTOGoPVophCoPOKSUpvcDdaQ9TMdizkbdWnfoZNobNS
UFmESOwoUPyQuJXB8RZm8GXkjwzFE0W8Q0wOL+vclwN7FAsHc/t7yfhMF5xH1CWn
JTrrAbIbQYdWB8apEENbA4ppIEVTr06iRAkUs/crCC0xxQHFxauA3LIDMhPmZNuU
m1j/FtgYdC34d9OUXNC+ukE0eB2zIgQrHAzD4idfB0BK/MPCUuUI8SEmeXVSN21v
xEfX+GUWBe5dpfTuezeKIHGDxw/gLuCDjYfBJnAAvenFCvorJlLovDHCi6qA87mY
MugsBSPw8okecx5JqPCIWvttHK2JwGALSAm3Av5ubdQXnmJ9aD68+OlUVvz8MyCj
PlqTIZtsKXCIGt+sPID42+d1RteWGAlD4vRXt0/xmQSuIGIB1qu2HobmkSW7fHXL
FiJh5qGSEfSE/gkW+gxMp4zNVpnujw+Jh+onlT3QnJutAgCIo+8MKxAdGKUaWXbC
F7Kv34+czJgUudZYkG6WkMNI2rOiy5XK+PTlhOEuDKbYefu9xjMh7rX+26eSEy7/
VyrRqPCPFXhAPTBgVe/x0dgIw4yi/qCbi9z5mSUMzKcksVs8m3aHh6PPKI0TMukF
WQ0Hcv9tM0D91Zucv0bQH1MIoCSRdUtak9Vt6An14C45TVVIeBcm+pJtSC8Fc9jy
XKSdrt1gYSoPbG0wPIJQYvtvq2FyI9lU/kX6ogK9GO13dv/kr4jjd2cSM4KT6113
YXqet43xtBCojsYszT8xsgFDETK4f1X53HAYfTJJaqRBb0au23PpVF+k5bTeh5xH
DySCfqH2biaCp17wVTTols1LGc9iNFTpmZhP4zOUZ/YdF4QYLdlMqPBwat4ewWjz
GtIkUUGghtJv77UZ2WM1RsszIJVwkEjO+/g3OZ91u+gSP3UojPmEJIrD5y3y9d3e
AzXhFtq5OeTJhsHROZpc/LSvojBVg7opd2OqOslx4+1oA44285PwVS/3y2oARFql
gRC92+vuNaGpioVW+3StptKjjU9xqnGnfAS9ERD2D8hz8DyAt8YEYHWKPvQCpA2J
30fB8vr7L7o4tHn4JSzKMCaQExNUIxKe+Bh6tJQByvt3XcAVihW/3ndHYfrPuZ/q
eAr5r2ju9kMC+wUHRgwu8K8Z4xp2OnUL4dTJzBfyoBgYdMFy/FZ+plNKv69WbetA
W6s6rf1zgFCnu+nJZ+bmseUsi/1DsDMmr/InXmNyzj2ZokDAzzv/rUctiWQadikI
+6WUitDl4AzkOcMcspPppdt04C558cN3U4UyI9YPuEl3+KP5XCEOZkxHUX3sqAec
diAjan0NEjpMa2lGUJOvKSpvhFnjrB1e7jbqvzb9yq726ri0ozV0c32tM6vPNE1M
adlUSLTF0KRP6mV+/0prGAbnIxBr4WmTJ+fRXzTJ+gku3hQKg73fZzsE/Jb54Z9E
6Yx9ry8p2Y7z6bvnhzq+R9RB6d7zNtgOldr13Pur1Kzqt/YSfBjqtBZjoI2pa2e2
/Uxf8WPzp9YX0kk5JCjsORLb/05nHfsEOXF0weef/Ifqyq51ghPsHQUWxsIfxup8
Doe8qO0i6c2kODXANK9ZL8Mfc/oaJxGQIz1hdll7NCgnNCGXBjufrTkBsqq9R3H8
Pru05ZAXbrwxYJOuwn+aW6L/uaq+4E0rvobWCoddWA/jMtpv7wQB/V++I6hZxOUN
V1HA2ylRvaktUccgbGRtW1O63cMmgBx8giSu6ofFpX3QqYe1riJ0LN4QgA12aHz0
88JjH3EMuULMUBScuzwAMgns/lUk+gBPjtgDZpAuPLsp8KZwugbWg7TF57E7tok3
aNAgXnHl6EBr4ZpRZ4A4tPurqtScPsRAhD3qIrp3wxQ00nXirxr0dCp57G9TYZPb
iXPRPCNg1u2sk8wplGMhIYxfNPf8sGuDh+r7vYtt2oTv8Atq+gwn02YHin8i2fEI
Ots0vF7uYkOHO2XgSO/zjFw/J1C9ZVYEhM9fntmzI61bib/K/lEeVNX7FK++kyaw
SvtRrgMhENGrYH/lJDqLlCWa0xzGomXODWjcGGrCov6cwYDbiPjB/ltyzfO+3mgD
lZHi9SIYH/45U5ZJf5mUCLw2IOzPYQJuq49iJxe5esND3a89ELk02/n18OziaM9+
GnkYhrX68DqdaL5Hn+gCIzguLakE3L4ASWOMUhNegOMe6SKsieoPRTsRlsdzR7g1
4JfO9y3X4Dq1B1F9SsIYGBqklJ6YsNI8jdUF7PhNt8sY3mh+bZvVNug7tA6dtfCY
7j8RvKZbD31fa1dCpf+KMxreD6F2B/IltVNgy1H6qyx29sXTFOZNF92uxkH2WBAR
sm2YJBYyYm3HbVspy1ynK6tHwNnuY4uRa02UTE6Fl/FibV1NIFWhMumjUumMITQX
j9PB/Ygo52eiMePjsqKMdmL4+RrtEbiYJjyhQUb0K1PjuBzUbDBBXLFOPB3cFTwZ
iVIEXCbx+XyTXnAINW4pVVgMcD7/fgkBHiROgYd6TuzqUeLc/ezKIL2zl9iPPjue
cvitnKol+CYkmBEcryS7uQm2W4ldb5HzSGgPhB326eY6UibBf9AriSTsD8Yldm4W
foDEnBfiOa84pLOEelKmuXMuGBZant2w/2oqBykNkUoEM5bg+Dm4wwvZCucK6P4S
U9WpXN3dh5ZBqq9ljt+sgkDOg3y9JbLdvPIPDZn4sJzAKIu0LVWcr0ZQkoQ0dceF
+I6wQcAyKdJ+zTR0XnK9LgWuvnvgj4ii213wk5ERp2SfoAerIrnz+O7XPrwu/7gL
MGldYFuDfZsnFOGFpqpvd6RCxXddwHqPvgXyk1GuMWV454b+9mDVFhesvuR9aOxz
Bq3QTVRfU6zGI5c+4HTCcfhGheDUHwBHbSDK9hhzU40Hf6O0DfKG1HF65CCbbcHs
DKfYdbEBjUQghcUThLMsGlTpCU9MlWNMcRe3OakfM0UMqaSpVOkxfnZbuFZ/jvEK
b4/df+HZ3e5HFt/j9tvrn4Q6FVDqjdptb1xZObRy3UqR7bSz4oF6KhIeFg0uWYWw
yQ7Vb7ReyJi3PTnN25sRxR7n1dB8q5E+qIlUA48v5MIjEhNf3D3lDP7ZsnKm/aDx
Gm9dSFZIJrygrq72VNV8u4IrGIK8Fv2BAwRI8mieb5TBT/buFVd6nMxmqo36gwlj
dAFMAGqzc84nB7YzZXa1xAuRo6Ig98bxvVROZkf2EmEnDS+3wftDDHMJYaw3jgUJ
5Q+5CPGpC0brP4zPxNS+Nbi8GBnOQyZFSm8Jd/1GiOlJ/Y2hpFx76doZJ2d4sZmj
zLR6YjRGdA2ATzSKbJySxJ+CJYlF/zfuiTrdHpptlmWSmAacEeP7DIfn43+mX7cm
MD/8jgNdgtUPQvSdnaiitk8ddXk/2hr9+THVpYboPYFDMhrMO+2ydg8rdK7WDmIB
UnNp7l/WtMIJHaT4djX4TcDszpFkkvoaGm/TAzABekIRqbuQF4re2bbbYgCB5VOC
Tfgpx8B0Ue1CfcfsREG/qIUAB8G93WNzSHXpElSRCHqyK0w/DRVEFx9UbP4WFsJ2
3cV+acqowSa+uMlG5Tvyp5+LA9jpE6L+mOWlzxLp3nF4dtP5V5QCiORi/RBJv/kl
Fzj/fTcVzwhq9fRSfGE+Yk/ywcyEPermtvZqSYRQl4QR8hYr36QtcdStRLyJKOgW
r8CxiWda26o3VSPIYWgeC5PQyXGsR6zwPhmYDzNK1Epmv7rl1EdVGBZrc4Lbkw5f
gN75Fa1Yp81Ky6q1VJbHj1Zy0Rq7NBnLB9aQYLKMQ4Osu9ZWDnM4Zq+c9+JLPQ7c
R/if1rfk4iJTCWd8o9V/fNBHHCrT5NPL+fWtcLd7J/bb36t+5bi4W+GN6OzHmV39
X/Ieei+XV0BO8VnnLfuS7hUNUnpDq11qTdyvAO2tfarDMCJL60q5JEFApyFBTueP
FccgRNu+OGNjV60QR5r+eQp8uZ5TySiHZoJPwKMPN9dhMvE5/5r5SVHuwXyG6Ye0
eFrVDdkJuetRRJrm/hrpAyOrQDGT7FWRwVXRLyRo/FOTvM82j4Pex4fkrK9OwfjD
5lHABBjp1w7QgxmNhHAYBqZDAMFV204DzC1VgD7v6IcpbF2M9QphyXOhEV7bvXfU
AlFlO8tSheEhOJzuH86phjxmsqZ4LuNluC07Z+0/D6HO98RqMN5Um0LyO5YB/+CU
WQphlA3EkEbQ/JAh2QqGOLR9dgwJBLlt3Lpu4hMOYMuwZVOjh9Mbf5YYz5zbhcKR
EafNDM4Ptdwfhmh+ILzxpq7rMAet2XQxXSY810Dk6XUDdrJ68tOwY3vVaAAZp+q6
EzA/G+AMgxdczS8ZfP/aaszqiTJ2VvW8PDI5MkoEjoCj0acVMFgKkSsZ2+T0EhPE
zUhLwEZ5CXhhPh9f+SwsHOWyKyJ97StQeLo6i/p8WEKdEToCGGJDCypOWNisAPCH
Gk+iX8IWDweWm8Zc9r8y7H9o3mBO4KZwZM9V5nwXh4n2dR+thFCKSiPQNRRhBmZx
ekfTdJaBfJts2og2XO7vrFhaF0VavKqo69XoQZFPjqy2FtIyYAlmqvKoV28lvVUm
BXnVxgtLuv/yHNUmRVn23DYDANvwlUJ+cNOkdWYPORE4ThIQ3F+VX+eeGsWyYPX8
mWNq7nHazAoDCHVyUkxBNHuty4w4myz7DzZMB0cykWpYpu6KL3KO0XnC3jTpIFBm
dXkBAuQVQm4P+/tNkOFGSk6XkeUfykmaXB2FJ6kYY2WEax30vW5pj78TZzhmc/ff
ky/sWftrsAzd7dv73FooXjsaA84aKfN5p6F4or5oDmyuvY8zU2eOaoto+Mw6a4w8
VV2hWUWm8OuD0W6NDn0bv9S87UP0sr4J2g2DC3YGcUeb83AYPySmEbT+B2+W0h/h
HsV4pn2L3DE3ok57/q+KtV7XRwQdZXKKzpJGV1jtOmr9Lt2AF2Tca8lD77BSJDr4
geLVPBPyDhzWg6lzPm22wEiPqFwbHklupMdYc8hQP9fk38aP4px9y5Uo+YjoCYaq
Y24+we/YadLlL7lSyox19agWmsg75N3fx4NLNRl74GBx6pea1pDvRxZaNQ499cyr
RbFzG5O/ZXIHSr1PDh49jOlvto4+MVAoMYaJvtKikI9Oz3shH7q2eQtgMP0vLQSY
+Qsh9BbKHsAFIWcQJXQ9Q+iQLsXFCT8GWJb6w1iPmf1+LahfBxtrP+SHnODcP/9a
Yg5Nl8jOPTksKV0/14pF4P1N1K+0+BZCiNah++nVQu2gPo91/uiXlIzzC0H8byPK
Yt7NZp20ajDvU+ki65lHgDi7d5Ga9g3PxQN9F1BlcK/TkKW3b1s7BGZqWNR5rcFq
l/jYQxXiLRMgwxf+MGMTZkFgX+p+FWS+3n7KOL7NnajCLo3+hM6KLLmjFS6oeYeL
8UdqjSj14LAk4QhmJGck8HyjmUhxeStBmSSN27GL9li3krcZWoVjErx1ypBQotnO
M02Q3Mo3/9pgJkACNj1Nt8e7iONO8spd/WWwcrPhLYvV2MBYMH8QSbRjPLEm0Ymk
T+B2XpnG62SFIKawAFeMlhRqY6/1SSP9HOfFnUoBhsgW9NWkmZCoHs9FApPNvInR
oNAqsoE0o85ZYxAjUOu20lbPCtaJ6WWQHoJxawqq1M8toKJgQMjQMRJXSi7Der9e
rTnyz4945Fcc4Q9wYPMPCYgKdbddXzanHPu9DPYpB83mysuVdHMv6dTsKtZ2iwvf
VAWuc78FSyGxtEawIJthkshPbZyk/5s+q4oP/b6e529p5cpPLPoBqn+bz++OEXSb
Lf8f/gtlvMs3+UYSddIZPJ6N/Mc+KOOA7biEGLgH4BtWsWKrNiWLcQ3VApW/+/cE
d4COcgqTaFeQPxyVRifzt8fMhggOXJGVHlBikSdkEWsAmmMhjp0v8nFOHg4GIG7X
xlFk373UTCNoyCYot1S9sJdyKnUEToerCQ0Ci/MrthQSzqrP9hE1i5Jh5hvfDhCA
+bE+75bgZ9fyeLx5v257rlYjv9kdAi/6F1fJv7tMWlwvmBQYNcHqx10+qEV0ziI6
oCD7Hsw1PzL9WItz3sib+hl61BTndY6CryZv1Xz3ayzQEDLE8Z/zvv1XZh5v0M5N
pUJrBdwjweLapaTi0TN4qY19tNAgNZowkOW+31Vcs8gHl5N1j2ckGHkYDynQ9xXZ
OApntNK3UdxrzIXfFd1pKIxlunOoD4mMOjUuR6crsyEwmgwCMTBzSoWozTkgBdbX
9V2h2wr4WizEoQx1AqHbovNbvRz7rPWvQVbCcZLkVc8IN+usdf6zSwxLhmsqiely
gq/YZcA7yUvvNqfNN+osFUUbfFx8Dqny5WiNupqvItDmIEZ3aCguHoyWifQIpiv7
FXq5AFS2V/Jsgd8hO4ckPiiF76uC+cfKu6wsI+qciHW9IBWDMxR1d0IbWibF6psU
8SnH3jhlbF9h7eA5YsUv+Ln8KaFCkl0wszRiN5ZS84FPZRUdKTISfz1ubPfP/i4L
pRk6V9iphQ8JJ03lolsbCBBQER0zT7vnkf3EdI86vUV5hMgiAL4R868s5n/KzfUB
iWzmVOuUHqqlQtef0oJeUkrx39OaNe0KndLPVMqLbg8zD3PB4xEv28JJdrQMeDES
ZfD+cVTxSmmEhKDu+tWBzyfkwcw4MLNhmKlW9HuaTQWQjCgiJSTxX+izsPY1t49h
JRpLstnl0R/xEw40SZKH9LMD6JiR4hYlyLgpVUE790dUVi5lgTVZ798UPZ7fTNf/
c0QISk10RBa7j1HNuub/KjgjPDLpVhirYXeKVO9aMtNoeEno4oQCDg5kS1HF0VAN
EEtoZIU+4h5ok1k4JQJRUoIqX6TgpuVu4lbuScu0brw+Pwe2u8tRO+N+yWPXWmrb
NjVViF4xyD8vjw/UPBPnd1j9wh4FqZbBynyMNLa2zvdjjAbYiFfTWdCAsbCmslV+
GwlQeiuvSAtnd5cYsMzgle6gbG4R78tZBKyp9cq7s6FglcL/qoP98qZP1Tn7ZpC9
iF8O7yeZ+ELq4HL0vUZfpZ4ilLDvQdTWMoKpNEX2o9CfdUL37dJN8eAPudn2svZl
55p5jdK3e/C8YAEkaOXCEniKqVRpdESg+1bBvXeP9TFrBWAfVYE7kzgFEzRcHdx3
UHxPbnidzSAOKnufSBnEL5YXwDyOGG+rSjfExY/tH/TP7NAQCwXtHQIGL5polORG
rmVFJNiZLv2OvhKeqitD3OJjqy2i3iXHYcVDndXE+NRmplFC0fF2vzwa1R9jE+8L
+mjW/bxNOL5xDVD2innxjWsPSzhc8Bqz5QiypSFaO760zLc8Rp5rV00gX/PL3q9V
bAK9BuhTIrn1vKD1RD3ZOATD/L+ScH+JpPncpJ+C3kAYJrq5iWuvzi3wEmTKQXt8
v8z2bxoGIoPSkfKgDATRXBP0fpUGyuDZfaq84ZBXHmnw3zQ2Tm4hjbqyCbWuatpu
varP0MOmC1+Bkg8hcYdYHSgl/yQa0lU+DP+BHRU7aFFUIXUxIsGuymhjoxde1bVB
04NxGpCj0CM8S1yurruaqz+epWLUl6QAv/Kg/I3d81ItZT0T9sJmZRY2uZUR/WDH
BcJne54UtsC9bvEbSItCVEublb8uDoFp5oqJcD/a+RKCWjBP2kxQOP0+j9B/UrXQ
ScCosq8RGH1+20kfIQGwahxaEwbaI7FDQwOaYzE7HSQoQEDDliedLsaexyiDCnq5
HAwzkE0M14JCvkFg2UuxxOZb+lEpGZmdJy1lzA8wll129jbpCmcTZGtBbNRiGul5
raNjC8V7gGRg1FGOGr0SByfUSD+FeLyQ63akZ+S4uHm+rDHzNZECTU7tnRSR17i8
fA3UsCHW1EAWurG4l4P7DP2QIxeLLlAfoL7557fRuhxe63D3wQZyz0NQ8hwvD8Lb
KoZmn61lAQY1Hwyy81QRY4O1Oto8fe/sQsnsc9Q43pMJuisDQkBcmCIh1uwKpp8c
a+83ae3mZq4SXjFCqinyJycPK8kPeciIRRF2O/gLAxyHqTRzgFTM/Fv4WuBmlDbV
kr/zH6lk/iKzrHV95bcwXKU1XzukzMdlLEXEd7qLAK+a8leZQU0QpJ3gqid8NLN/
ia/MiuM68DBy/+RwwbceGzuborbAfefXJbCq7dH2B6fu/mJoxd0pKWUovBO40B2K
b4fv3mkazBGfjjNgbZTVO0JkzToMJ7xG65BIYNELj+aLhZ/HC906IkdoxP3u4fQv
gKcms3aC/0aWZb+YG6KnUW7PPBdhnR3GVuvEuszSwCMyhI5Kh3UhyHBuhc5ercdr
HIT1oh2CiehBhOrUCJB3JcMXdlPqRVx6XzNu+m0kQ0ri8o6UNEZYozGxBfe55Zq5
wsC5mjh5tapznWO/3AKbOuqWo3YS5AP64ZfxaHOOoTF4kBNwf4fS6I3a9RHKDVy1
McJpGmoMSBhCEd5Nrf3i8MnmqoZfgOJmNgi2OxcGerAqJ4fJwpMjfCzQMq8U8dC7
Z4Bkl+YP79RFTR8SwzeoxdLxWoPacga6I0k4OXCBCIRBSkLo3R2MvAuTsqY8o+Tt
e83E4tH5OpVJgmwtYN5PPDZbQGFQ7h3TfVksa7I0OlnXLrG8gmLbl+O5x0LWXZ/I
HkrolSc42iO73MdrZfexkYbDIuGepj9arE1HKEGzbVbx+02c4//vWQFiD+qJ6Tvq
91pcoqFgxCQuD3HrE2IozBUJcp0Icyh8TOgEk5AtaQ4beNUsC3srwyMr0gwJZPNE
HWbrBVxKxtkU32+V0z/z5E3mmB8WOnSCSn/t+Kv+/7Xkll+Wma7HACySlZ2AdNqN
PJ72McZlGGAHdFN2FTUydu/1h76JWHyDUD8xw0/46QpraWymiCJrYahWUZFPaSil
h1RwUCdmEK498mkXWSe/NIAwyduItTE2rhh21WKlI0GhWx7lCen110bXJYB4IXjZ
4T8rfx8d6w5hLrUzqLyEpAuUemUMVKKI1u+8sm1TOrkdEzWTsaBGkUcvfCkEeiu6
XCJLcuGZ1IX6uiy9h3hqtgtsLW6XQGGR20nVIE//2IQvqzNdnxlUhsqHPI5Y8a7f
ouqnTiKLM9ZKfgBZt56S9BEeSKAAZ5MSVbFTnRd9Ab7c0pAZc6D1o2SY9uEXvzNz
qbPauMDYzkN24WJ/qR5qZTehmzF3G15XFXpwPvvO2tCyKGV9sYfHezBtSiXO8eeU
f+iToPh33sc9lhuZJZBapu6RlyxmRzJVKn1Ad1NP8BCP6yfE4KcPPxQBCIc+udci
ym57VgGNyn4ttdLFym75A8Gn4I4RN9y+nQyw0E5MFvr6RterbwxG52byvH+FMOHE
ILLwopbowmGJIATNIJ3CO8Gmr/rpvOuBVNQRXD1OYOpzlSvpA0+3fPmwdu37qCng
a8mMs4LoYah0tLHHMbIH0aeL9YozRDGZb2aNfh3Qjf740sikZvz9RJuVZP2+IjUR
eFMnk76+Y/HvSgvhJ1YFC4oxge4eGThYTU5Cw7CDzN6qU8nim8L3h6s6O+TkWByD
mJyVBud7SkWy2i3HEreW3gS2Myd4Ju9T08vFNrnjfkS2uM6bAEmOvfly8PO2sJ4N
+EdGf/xlR3/e15AYVAEaMZPyE3ZF7qin8581lB8jNSxyKW3gDBmZ+9+16oW7GXQ9
ywQoAJYhcDOFjDNmKyJAeHlOZLEnTjaOmvvfPowrI0+r6KNbwRW9PWM0AhB7BqKQ
OmzGG/QoGfKhpOfS4uqn7Y0FiO5kFXiD8HLgcInJPzEAilD2RBlwr0wTWs1y2lgW
7fwc+NhQpZXmtzS03Oy8vth516xlT1KWhPIoDB6dZ2TNymk2MXGxFy9dKI3bIYI3
AAtzCu7t2XjnfFCzuUREEmoje3aVVsvm6D4zYhhftdpGBW90DCM0pfD4EE+kmNZ8
M5WjkQCKRphSQvjPg9C7IG7MTprY2QXbTCJZaLyYoVpHUrzwrdFS/NXzxff5sGz/
nMQeH8mnzUAadq4ctSQ6YGyM7cefkEnm8ykYCU7vFB7rhJr5YKUvaOuVXEKVO5uK
vLhl/vVyOKvSVyWdfVqlbGCAqogNOWrHPyYQWZU1pZYnaVjWledbS9EJROyHDxlV
Z67Wv/dte20Tec6A8ToIMizKlSMjPKq2MRUHrJ0eQNc9nFxPWYbb2xpl4qyYF//K
GipUOWwlctrM/yr7ZaZaPWM1rwyM+gqpNbtndLd9vIxb82qtUcE7llm2HVw03s+X
16aG+2NGAYmfXsyvpjpLHhsPlzVgaXkO/f7srbPD6RMvj7+RSueQ0sVYOhEgEY1J
GfoEyha8F7n3P7VPSXpwlN571YUCsjZ0nWcHVqKeTYX6E3uufRPWuPuuUnn8P9qf
CPf0VaRE/+niYPdqVRS2hlHVCl3FXvXfo0RmS00t92/Ab6jzfybCunCtQCjwlK+x
ysA8W0UIgRRa+HenY6e+yyB5CJ99RH2jlHcJIIjmD18YTff+YalYHCEQa9ux1Gty
XEnX6zYRMqcsiJfT5BZoH5X/KhccusS9y5cgtL4oTIEi2dKW2ZQuk442GsOP9r4V
0UGAk44Pb4uukNjxP+XZXp64tpO9gE+qn6eOEkqJk2FIS9V6Zw6QoEOwXrV8Q1Am
T+JLEv+RYE9tpZ2v/bFc/zmnIx1HwRrvxcSf7o4j27g0troeXM74XNMpQZe1uN31
4X0zt9hWNcUA7diFqCwGTXZudunOpSxVFG2VDUXpGqQB33iuJIG40GLhdKYLZAob
tmcXwbBytG643z01RObj62MFhiGJx0qKZanIUI7lxgr6Aq18ExJ64UuXwvKn3R00
NU7W/ODSqF34FEL1Otk25opsnnDzZ19w+zUvn1O2NssiZQou1BweBh814KVNsSV4
0X541yJMe0fwlxzNFdkuYGzFB4rRLQkWbCGSaxLMVuZLZ0e7uBzipnSVL59qPIi9
84rdEkgNPoc6/Q5xkpQJyzzzEX+svj1MsSdmsxvvUoHuS7/I7XnVastpqTeNi+8H
NjDSbFmH4N+uqP966CxOVbcSMRTWLTooV1Dkr/SN0graw+HjpAJGeA8uRgIM1my2
P7ux0N24FCn2qOjV51QYQkhqv5IdIomELgHThpyCibtZ8MgDf6ICy04Km8e/A0tu
BuLUIuKQqJtDOS48WPwqFrxn1Dbo76emvHCGPUHjo767+b4rEe7bM5/aQBwKlnLD
ynRLlkXKubaNeaIGiq5aK4LY0FN9O0aDm2Qm2f/szTNKm/QR+h7pCoOi2U2CpyDC
ouS1MPUbUHSA3RQAU8bWmysgM8y4T/rP2vLCmHdOrdDM/f9O/jt8IojEXToTlDyx
YRmTdJTcZfSvssCre9evREVVLNb1FI0bEJaL4Qj7riF4PwGNxAUARRd0d8IjgvO2
cEHsZKmI57nNkGn9UVsdP5B0doyfr5nliGuSRo09p3JOUnGYIyEfsXMJ9WWurFYM
7chrYiz9IAx6+VNkyoqAptiMa8X6YRdXmJkuHYMa2kqSbfi3i1WQ/DyKMSAOJRwh
A6kIm9KAk6dmlgZrr92dC9BKvKLjfbkDon2qRQkcQFE4biMKCAg1zTC7L8i9MiOX
/j7JBPZJfzHXuvxNwqh7EbzpWr72vrnO4Yy/Wq/3mcVd0ZfE9dX9aopfla1igt4M
NEdywucUWnUt5FAbivOeZfVO1qdYO1acnh0fTJE+VK/iICx6h5xaU/dcFbO3gw/B
l+uz7YklWzssxlPx8WmKvm6e2xUrESH4pg6zYdg/StGHaASNtCv6qLr+rv0WGrMC
zEhbnPITsHZ6bkToN514YYeA6yIViw5LG0H2t4fZTpi8TEd/Th37466y5uGv1dd7
ckVOpNroP0yEHzLKB/djFBMI95U3KrKgP40SX+WANam/eAOqzvV9uRI+gfIDm284
ndwHWxiJfFiK34qIYCalJPMopIxq+BUEj5sGErMH/co1TglKHZXagYfyH2zV+7Fn
ubtHFY/4bHu+dCOMppq/Fr18uCCw4gXe1jStu4jm9GFRPcjGjvnDeRChksk3rOZ6
G2VxCupF+sQ7ZZte00h/oiyjJNa8mZsiiHEUUYzhMyLFq1g1vlZRREWK5JKStOa4
ShNlQIOZcLUuoC1JG3uji1Krm/MhdqqKAHHmpAmtykJHMPCoHNadIjlckd3LCUzc
OXGg7T6hZtn+unS4wSRIH7aICh+RwbmESAuajcuQ1DxxnB1LLMSQLWcr8HozDb9E
dUfOJBm9IEOH/KGaYW7KUcoNmCn3cIDYbFMO8K5o4gT+6u2oKD3KDxwwlXcS4XB6
4X1HvWgQJQKj9K8dg+hd9X9lIJq/eH9WRyHQrgzqNMHBzy9Jp13TWkIqal773vxu
COazY+/y9EP2/wg6LSLWissxvdKvR6pYVvOeVyLm1dJuqFAqxGyNktfZzQKSyETw
vVZgIFNujRXcv6ZMIHrbXYTesdP90wu58OK06ubJBE+IiB0zpO+geE6emT6IJYzy
HqPosBsrhXmwwm/lWicVUZA4upK5lSi2iG6u8JwoKS6o1XRGsCW5NuMSq0GPnPbx
aL0KAJve4N8ME3JLvq8I8nDo6PYl9MSiRCned5h9jSpKu5Pixk1VvpPOwHo2sAO2
3QZDAaef5wfpRafWMb7QHm2Wcz4ZA0awthEVMGINQdis5ki43j1JK5JSHMLiuQJk
h3HsIu3+O/j80tcZFMnQeOKrovKP0LZQbheXK+dPIGetWQnDxfPXrtyJrfgwjIw2
db2xZhYzMpAKS+k9pKWOGIWWpszLtjDSfzUSrrEYrxiQmj0P0dgIH7D4Sjv27eB6
RMQyYTZcVramc093FVSRtGmRxOpXTU/A97bLLcZHAXqVYu3Gj+9qEr9CdLKFQxws
OGK4iY36HdY9G1hqYzCrwyaERN/FWnZ2/xMwwUx7skALoXkkCjFQBwLv8A5P2eva
wjUxuoqbn7UEHzzR3T6rs647YBtxUxJLc7e2k8yBlQGk9W0kgnxSE8yV0tTNhiVQ
Wo7CyOVc+kw13bCz3w6Yw1WfKIAV5uRl3wQJ2yMk0IqC0BJJVUeYVZOpR6ctVJHX
7Lb4V5Sn/faGULjAlc2yf1RW/wsLP4PG9gjswMIb1sjpbnWBWlrWpLb/HIsg5Lfw
5IVELvsFCuDdD9u1q2DQ5hNZb2yGybG7gc1YzU8vwuItumbAPffQxi88Yvtvb3nc
dZYw6LUI3sXIX35j+6Hn8c8NtTihO11o/0erjYPM2txIJBvvUdbOK3tgmUb0A8gX
njt7vMBSSXmIv9z0JODGKslyrsvvOZl58aY5zSp3sIaGw0CM+e/EC1rkFDcVBEge
3Bo1sGccdGcDWLsfilccjS3jg3tEcUfRP2/a0eb8Xqxb+Yg87hyLJsfDLmhm5tOG
6G4QHYHmP+0VcbEefl4Lji1Oo0hr50DkR1CkbweleKSDnw1rjlSCCdIOVoFOhk7O
1IqvaUbnd3/sitBVd41t9JxCfH1NtqcRgMXlsbsbw1m1GScYrXi+1oA9g3eeWGlU
1zxgKAGyT8ROD8nllhJR1n3ytp4sUowsgLiyrZEGrUyTBDamCFnk20pp40KMcxbW
fWDDt6ud3JT3nOgHeUmUOeDWCSoCLBa4646+9njh6yeYiOmEhj9H1z9TRV+C51g2
0qO+/ji8IN0RShYlrclJyUQP14FA7JvR6UrOcxRMOOXgekq1ey0Fac+C5jg3SRq4
ofLG140P0xjaLhqNySIZ2rWYfebjqgDmBuxQe5ZVNg25EzWN2Q+wqR3jQalb6LDc
zRTlTIY2nlVCh+1AkDF/fwpVWx4LJiZDIZuqL1VEX/3AfEyowHSFiy4G1c6AtlWV
BxcWoplTA8p4xJDFuFuulXoU6yaWb3EZZ4P0ARhAuH8j2xyJyVc3/GT8VztibFob
LxQLIHdMe4OgFdpoA70MJoqCPLtdNsi/lJpro8TJMJWif8R/wmiOw+8vSOEaf3ug
q7/2rRNvcjCrkhrQ0jwa3BJCgCz4xWkSflPC1C7c/D1JzUr/8H3aTRrY52OqPRM5
y/vRwJzyRC5W7W9paMhKFqLifVceHmUpMGVLRV+0BZa5q3j4AE6srlMJnmTF4lXI
xdKPRSLJk8ho8MWvXDP8rlKDPPqcOXS/y3wf9sYWFJFBKuFhlZMXifonExBCcqpC
sGKABUtuB9uP2oIIcrirmsT76YmW9vM2QJjX62jeevWroc16wkJu7L4YggfmAq29
gsGl49Em7gfSiGM1HA57I9Xy/T8BU43rHS7oBk6eUcxaaHZ26M70BI2BEQ8VYkh7
jSUnxI3CctQY4aP0Ctc0XFtTIB3VJMUuF9nyWOKeh/d2moDe3CxTC+9b9j/Jp5o0
9TEkm74F6vtTQpgPw2Q4z4KSEilNp46AAo4M+eGwvz3ATgeRsw23RRUYyg4uzNzW
JkbXDd4V1fL0q8By3aPW55rHiObTgja/fxkjHriETUqf2chQ4Xa+stx+ktuhbT2r
5g28xjtmv83JlF3rBhBE4x6x3r3LGfArB4jEKLjPQwh20S3MnbeH2/el9GMBBy3v
lc+H0bkkOEtgUFOolLV5TpFNGs37K50JundXAQZnq2SrHMIVQotd3eSDGxb7f+ew
cbF9MCZFqoOhW6s33Y0m3h0O0okdzhuT8HqlQszJ/U6qZCsRHo2h+qa2Ir4ly/BW
KcZCiVXRAmsk5ZjSC9ZI4c3rzYRZnVNcafcag1vO4KXw2T595D+v9LJ4qf6ImFJ+
prIv/yj+1GKuMRe1PtdjKef5+Su5e6zlX/tEtmkz0P89YYt4Lko18wHvgk/068Q7
WILtv/N/BfAH0DcYI2TOGIOPcBZL2MC82SJIYFLvHMbSeqh2CgpweuQiICz1oOpZ
rf/I+XdiucxQ3SIKO43SJmO5HuZNhGNDwuMSCrWka1aOD97Ypwe5dPZMhDA/JoKR
4fIkkfr4tGCKHkbcetG1FkswT3VLa36iDHE2z38xfqF7Tc52yscrNiJ5aXm0HIyF
32gFya6q1r4/XFXXXtclFbS3sQOJ3rPegbyFreFugJrwPhKZmf6MRU240xOICFs6
vXCsp4n1IJ2c9weBNJddRGkghUyxxVlJZHEDGm4cku16OfZRfycS0m/wvVVVuRWW
16Q6M+7nEMgmO7WbmKD36fPlpP3L2koWRqfWhko8RrUYolodBushhxjmZucnEtWG
sXfMY2qrlAdMzKJnwfPj+PDnCy3tZqw4QJDdPlFqJqKMIYA73znNDIYOph8M5H1/
Q0RUsHxtLrWo45Tp+nRb8PjINngl+f5l5febHnuQQnztWj8QIGfF9/Qq0FZG3X0e
Q5OqDkzLH4DfkBbIzgiEObou56bHjYSLTqyGOhrq/i3aj7yZOb2woYhJ5/KNJf/v
jbgVgbMuvH6UOweyVoY/RKHFHeFiEEpm4WgIm1z6xtO+zBaqDgBHJ4eBEi5vrhsN
kNDgIA5dq1Tf/Z9HSqw2ul4kbhB3cuZ0SbvaRh5yBJn5MCn9ER2YkEzjzUmU+fGf
+pbMsmgFu9sD+xqe91OJh8/tHYh9KWELTk02/zP+w0PY8yE/FyKVLdFWyIYWh9KC
LG2ZkiqoC0hub9HavOut/xWGu42BUbVDBuJR+NmWFSWNzBAR4orBJ4vqikeUPPC9
XTyovQEvd/XSiG2p1IpSQl3nQFvKTKIqGO6NtXAaTf+hrZpYrCa/SXVxpQ8TiRD8
mSnJPPBicckCb8SOnZQneofevlmUWOGGplJU+QI7QgLUnpRDKTxkXfib+otnfHeE
XL+ic0ZTA0CYHlvxx5SGCmBlB5OEaXujJ0Q55cBvh0pBG/ELf7i7C2it19/y5ubL
3/SvHU4jPLRx/cjPq+/ipmv9PsV0ypQ13oeXUbHrc+O50sA4RH55gRYCs8NRmbYR
z5+GrQ9r9phUJ07ArTK0PQSeFdHUSiKvnyjwwB0YWoMycXYCkD4Ho466H8QLl+UC
Mr+zDnD3Y8E7OkbAUiMegpz76/MoC79Q3p8AcnNM+tOFkFs6nxuB7h/LcJzwi7f8
1SSV5IkmBz8vUCUc7jG5rHP3Sz0g22K9iqHaj8PKVndYzHNUbYps4t5wzc6XhaeW
iIZSyn1cLk8cFqcKwXVI3Kj8EBy5MONlp0MEjWkP5qudnEt9Ipith3FHXSkrh8Ck
BioAEfrsogRR4wsHwHw2w0tD6vACMRJBMR7rqdXDpem4xAo5Q2KDcULI2Cv/g8QP
4L1ZRXs4USUOvzIYiDwTvsb6dtFltc0kwzkldDbsMsFNnriupM15eTAxbjyD6fCS
q/1tRICD61+wsp2K7UBF+uR08kOZ9DcRhYHAb9RcRijz7ZOwjfhH4Ph3W0aIa2Ai
e2veCkrRHc20/LDsB2mct9GB/tzX84waNKWkdspVqIGjPtU7La4dBxJtx6/BApHa
JTd9LhVwnTNtD2DPJkBD0qvMA4li6iTuZm2PHbQLJWZ9zwI/XWZEWT4sMQaRnwQK
8Aq8s7/zEPPtYsJHv5n+G0RkPxd/17P/VawPzd2eLer6IH4JcpGiwUKpR1f/xIU2
iE7QzjRz33gSVIJBDDbzKTA5xC/cPNs0tRkTavqXnavFp+Xf5p2mt4yg9o9Hnj0Q
IWUwKoKadKtO33+5ZH76O64zMswwTTmPLcWELfGvTqfvaPXCBTHOLM4Pn5OUCXLR
8+sQMUnhOv4KixhZ0hfqL6EWU7YwXs0Py8chTA641qseS0MJtqfUrFXMqCSmEYk3
fQ5yV/ZVEMMqNw/mw95TOvfb16TEnhS9pwQc2XlSoTR6D9GMKxwD+LwLbtDefhmk
AyRLP5w5osF6oHPKqGOHledkb8G+elYRPkJF4b89Jv8hayXonTqY54q7s6jkBoKW
BPNOYdt3cO0rxsH00Qs6g5AsyQ/XSZKntyDX550DLCQFMCcH3+gP0nw9FBHikwYu
787HON3Kr503id8qnkw+Uu5MFBcvTM7BlffxON0O71E3fN8oAcUZbr8w4Ft8hdeI
4+AphNNDVt1rLVNp8JPDGqeSkO5KSoNtpCehJycWIR1ifEh5o2jUPOZSbktqB63z
8brVALzeURX62bucbuJzafNI1GjCnvVmVel58RUx33xgfNSCkkbJnROkqEGiMT4/
eG2kcBetf9M0DKkSkWOwbDfQCqRchYb/xgPRmJ2tQiewzw/XdQbnNHAx5tfIOJ6n
iXig9d2RVQidC34CQB+qipubk7SRRWTflmgHEtvprE6/YriIL0Uc5d61F2GQQsJA
3xveSunS/LmBQ4RGJPLqu4LEPr75ojUxWYaltt0Ok5x41ax5pO8uyp+ggviGQuF7
S3VkBBS8xSMQy40amf6Ypb6TWZ7QNUWjTN/QMl6QRued41Vi7clxYlzuZvCdDzcN
p82KZM+lUvMsyj3kKkh7M8tBHnWYruRXepuNhx9ChBQIo5nkh6wBtTwe9o5JJ1Zv
zPeRCCA7e4Q89QHCFaNVX3+vN4sGcdEIKT5zxIECCRX69hgoqAQ8C8NE65ukRf2+
soQkx2ue7CvAAk9wTZots8SnRd9LdB/MJtuiBNbxGNCMHHtVn5tapd9pbKDXqEI6
Ewp/EOtEl5w3cuKDiotwzOFkwbnVSRKxYwvE+E00mnwT1vdfzjI44NWjrlwIq5KV
8IVr35cPVCgCeCgQFqNi4EJHmRf1APE8YYoYzDiWhgICfXCXIT0/0/C+zQSSdyxq
x4nqzYERtxYn97HFNl+AwwpAXh2oVQ0y0uGPEYJG/wOHKSMrQoWHPcB3TpoBTo3w
fNn1b9Kb3UFT222kS8xGPtwIZI7PXY+cuuSOjAsmMVsUNmgeFJB+yDtG1cCjD+iM
pcRi0IYjrdb7TLGIE9snVqIsaKJ9/j+ggkkae2FeuD9Pay3i0bIC3AQyPGaexlG6
eIVcCLpN+s1evp5v1VOfp5mUxtA85Y8oyHFK9TsAaGUfTCeBN+BlbjVSmUB9LtnF
OOEYHcjvUITs3gc2CPb/1xQ+zQL+p8paUAC3sg6DCazmzp0yKVmAn33YbA9KXg4u
lugZqraFDrxFiafHIs/gmbbnlK4/H0FyxOx+wHO059GsYlKBZPFrCZc8e7+a/fFy
5vIyuFSw9Mp+xUyUyn+kF6tIyir+dZvm8LezkwsEpSY3KqUPrv1tiT9uyLDr9ryI
fg5S20z3ub1AQDEEPemZPLTRDRxAp+df0tn0ESWcB6uGSYgK0rMa1/ydHuWJz9Dr
SVRAoHktybQ4MI7y4dSBOr36kDqBzdYCgVF6ejAHYdgT8mkQPUFc3/rkWrYLMIXs
QIAvHet58OYRtOlmEmKL4c0I35Kl1eva8aM25SQBtEcx/vxw7pVKouCMX0uzoonP
5x3PkGygepjl6gsU7H/ifxa0Pvd/KceZ5jVKUE1RmwG7fUR5eNQnJTcJXc5Jnd8d
GoXnki9oIivBY7tbqDZA2qzyiAsOWnoQpWivVhEAO1rJl9VU69KZt04KlkC9AoPO
7AszXbnYadHw5SwLxfMmznQDUcc9+6IFKEvMMQBH+jmhm9aLRv5gcwKJM4lXqjrH
7xiwQ8psklJgKqhWDilS10Z2uTqCj+9DvaCeja3mrREyJqPj1x5U40LmGBUugV0S
xOXebtU6bzu/GbaMXGGhe0oEOltEv73ZKqiarpyk4uWcwrWkkkX29BlDnICk/jkg
hFIlw/rBUfFDVnhtyWn7qy5qV33UUss7hkFgqyPboVA+Hem8auchHuPyaw/CFMU6
yDrqTJxBMWHEfcaVhtCCKOjVrZGAOr/K+JXyPzSmvHwcA0lqypAZyIJsjgYyAezj
wjbEDhb9Lj8sqXG9p7h/DKdUHfpbdbLiXGTiEJc6l408lIdSZeIFHNdM4rqTlk1g
ipLIlqNvl9RtO+U4Mkbx2woFbrWB2Izqjb1Op84FO7lvXx1GHj5LSfN61kfOrH+W
OJ2QXUz9ZpbJesvOkH+rywcGf+9on8mOBIbj36H2qVMMMl7uFhkX3QsIVulvj4gR
NkKATgyp0MCvk9zBwmH7A+MP7W/MaD9YKfSF61jw56kCnZaPfkoRkvam4pCAYme0
9rFjgfaYfnucKnV5QTDTLtSQw2wLCJ4jk/vs3zc8A6ue94seBZEVasZmlhiAof5d
SJsXck7XBUrZ1btqilWkKY+AepE9Bz0BWyQgpcQQieR2TZO6iQPEiDRx9bvB4GW9
2hG7JOpbpIauTLRZq2p4jFmslsd7R9KmmFTcESVflnvzdlUu0+/dKxDacynIGEGt
LUPp5NM5ZQtB8KPRg+HS9fFvhxD+K0baxWKx+5hgwwiNiSv7IXwAbLmIsbZEyLG2
yRwmu9SC0RCvszWUDsI21SnvQJElglc62Mt8EbXX3MziNgu/AOIEX17HEnISh/zQ
UcYoWPO9cGkHYtc9zy/xfzecihwlLRGLZL2c4WX14e8/u+OnIJlo+8owloqRg5N2
LoVV17uh3QisgIqjv0aC0is9r/Qi8NzomPtGLv9+yGS0K/8orHM4CeAljZdx0LKK
TU89GOE8PR25j+12/IawELhXG9E8pZ5tsSOCorbQxdEjPpG7aPxVuj/uEsOgHl6y
QHu1SBD0+HQiR/ICt7nDqZaBZ0ZOStOLpWAKQFBY6xHbnZTmCnbjmLYJoc5sB7zm
KbprvPm1waQVSMy+x0UlFcmwJBteVRB+ySCi2+ReMqBTPa8cxudzugO81qKg0Uvp
G4Myo4x86uNUPCJwaw44Ez0PPD49lRDDrhuxhGcdRRqJFQY5+xHXsdKG8Wd0RWp0
mun4iPuxwuM+1WSfCGW/rzXLv23pTLTHBQiah2rIUAsl1f9CLcidthL6zTZHeDPX
ZhQ/TF3GC/GY6AcEr0OKuEQEOXjx8Y0wai6zAq/GnLpHsPGqPpAL0I4Y4cAa9RAn
vP97jdXjJFJxkm75H5SqRpuCmkcwFQQxk3y2lOdvfmsIqZbOdf79geWmf8ZpcUJF
gZLx/EDJjLQd0wWDvD6KQjjSV7vIRmyHcaAzMVZkWSi1rBF0ce3xbkDSp17/KuYW
bHZQhHBzEk7PtGg7TZVfNcrJsMU7Dpl4kvU64hL7V+uZ9x6w8z0H36xsMNltIFfC
BWOTvMTYtZ0+L+KRltciDQo/ms/NNbM0y3hGTPyZyOJamQQF+ijZEXQMzMIiywXl
1deYI7N3DXxq00wLTim8z6O31EpZTDsFVzlVf+qSzHEGZwEe4eKHRp3jjMEHXCoL
JKK9kMjF5nTQz2uw5HyHdv7J2NW4JKnyY3AQnwcFSYBL2etSz8Cz2gjkebqUli2B
kLQ1top9GnfmSf8fRIkcrXV++Tt8G5JakUreNniuFYv+5DRg8qvIL5zCJUKurMWV
PTiIG6rGj42p94oG0bpc2baOl0c5Gzr5I2p3GHbXLv1C0h5XKqPlUmBZCim8ffnh
Il8tnhIWsncUwX5mdEYe0q2JG4FF4PIjMfTF1MrHpEczxpe/GJYuwe/3oZeacLoB
Pfde4XLlmzTmh42W/TcddYCYNOvDL5isXvpx29QV9YvH7OxEqarCvX+P0kwqJR3w
gG7L4ulhmOXgKeYZDE3jOzUzYX5UNTn5y7HF55w9T2pvQ4EahoIPhSRM8x1un5r3
/pOlR/iQbcYOLxUUYOafyDkbbl5wqLishHOyv2L6RCsGzYdBKnSWGjaMe019slDb
/uAy6QKbGPqNd1EiuTkGrB22R4z0NIXEvlcBgWnqkYUKT4PLtdVJUvgLPjnvjZb3
ejMIx3rMusSPyg4zgzxbBUlZ7B6TLDNydxTohUgIMQn7T3sEXJ5DjCnKfTE479el
CY+VAKlNFOP8mkGCkVIwd9zUFfUspa2u646gJWmNjKz8srh4YTJDkWsS+jGz2Ft1
TJ9nO+G3d4CUlEgQXmHgONjRVLff6ajFPqoxgt93vznnU6AWpt+cDQU+dws9jA7z
w/zUy3D8tbl8OAP2qBp9VjL7fLif3juoyRtM3ASCo/8MuKN4VbiYo4h7ZmRUbtuW
VOdyWdQLBsCbX7UZbpX5FlWX/GLFOXVOZt0yfXSrPmnnDsIq6uP6mo6AA+iBPSDf
LN+JEUajqUeVHdCtGrO691xpCROu/DF2PQwVKb0hij6fPFfjDSMXDgQkFxesjBU9
37jVwZjGlNTeq5xRfvPyqrrEm7+VAw1rs6CG0oxG4XRhWPSFZmOaoW7coYzfVpMk
Nx8fCboiNF2EtClSo1uYWAIdroYfw5QDHqJnorMpOeo6+TZ/EGMnFgJB1joQpiA7
n0/n5oFM845LgOa3efhBDMydXNCfqyJQwSD+4Mw6iRfcwjad/OUb77cimmoIKVr3
is0UXcIUi8FiqiOP+45JcTywrXUKoxRAyXPCvh7oi+Rmupzxx1Tqt6H8zQyl+Yic
bm97wcDrSV4/p04StBe1Gvmr4B34T7acKBykRSel1hdTIDaDpSSRYiGM/oZj8pga
A/VfV5rKRqkybSNfmP9ZyoAoYiMrmMxdDS1/nqda9+/jiwH6qI1ZOtB9ODVk5qgW
PlcXy/kXb0wf1O62mX+c0/of68C4J1tHJaSRhn3/FvmpIrlR/v7xkU75D52kK6ZX
mmXqQSJPke404CqnSrpRpQ/bhrFcb+Ac76dL+qpG4W9+N2JOU4rDLzhMrCwNTfNA
WDMqc0GV5enOf4omwU6NJsQIwPwVuvfpAioVXTT/jwxOz46zHbmU1ln6XYFYzQm8
g2rODaFrr5R5WVCemRpYZGDf77PEBEHtQRnvDE5PxKhNi2Vse8YRdksDYTCHG9+J
0zuvqYqlPeyJaQDq/EG9tYiaV51cfmRjFeE1obodHmme1AzBynrOjzXEtmqL4FBW
0eN1D6CXCpiDlSKXqRLoDShllYPkUskyohZoxv/0Fs2j/h0fmyiBr8vgM4UT8YEv
46JdvJPX2HnAWwQIxrj23IH+Yjzfs3pughcS7+W6Emx5ANTea4iKApdxYIDtg0P1
SX/nfdZySWCYp7pgT6M5bAa0/ZU6IOBz1cX9Jp7nKBFUgtdTkSY79Qjg1/N/A1sB
bbiMnKHvPVIRlfUc+pqlcEK0ywF6y9ONe5NQMK3adXfaeA1zEZxHu3+fOQf609XD
cgGi3aYY/FAq8fuN8E+E4g91+fzYabTIWKjegygIALcML4Jt+PK3lyqfgaamlc7H
iQ4+OrwHXsluyXCaN6zzWVdYSoYnr/G+fBnsbOS9Vr3rXohJ/O9wZCcRxd2SrfMw
U05w7m7naq38bIQr8getfS0AkrJXVJCp69DUuLLt+9heOPrr+nJXTU9AlkG77xFc
6dl1AUEa/JHY3hfDAEnh8IPSw/yEMH0xduR214OlCemyVtyEu7NpgbUxSJ1kmTSh
J7AWah0cTz4UEFxYufupgowQzYv7Y0bCumeM7mmjeQADxObcQc/aThjWfdew0oSB
UyPiDQSggtoj8unXRfQEPnAF0BRJ9XFPGETs9bcyT3zXePyqTJ5xYrVOfCMXpCvA
qGEHTt3WjnzNWLj7oVQpZW09nCN2WxOT4dMn0DlUZQbDt9FZz0nWHP74Vf5/StZV
+jLjrz8LPvFJiQBV5aim1btXMZjXyrxkg9cjo+46jdxpHnczTENKMG1Fk5PBMfvT
TdJsXlyZ11Cm0T6rMTkg4oZbQO3PlQQIQjb8p5VO90LMbcSHLZZhWInDrOpu4aw/
AvotXCRuaUB4e3HM4OU09HLMYzbRmXblLjbKSoaJZRCaH8NlxXRt1u+PgmHfbXY3
xJyV01djqijpAhcmyTov1cWvUx3nk4HkbPwBPZPZNFjh6JNZNb6jEO9lkAPtaqAO
xlCY38O+pEqScoC40fxfzG6h/ds04oGsSVp5reeEVg5Lha1nk0dEVBQVzAuFiS5X
nrGkU1suE/ku48xg93339RMuzQZ+9z1RQa82BdFsTp82qO0fyspK7zVDDUfoEVf2
5ngpHmmRJU1nMIsq0REOKgpO5eDPkTqPLe++XXK9QDhNt1T8TaObGtWHbrazxKOy
FpqYb80bC/EymkUblsPMIkZyoElM11z8q6mU4WFv+6j4iHjwjLNX07VmokGzaCnu
tCBtQEVm2jIcY+q66Bc4CM/og0Eym90grQk4bH0WoQJp5klr7J0E9jzyUrE/1UXu
M0ZEMUiMIRKKVUR0PO21S/viE6nvcqcWCcmXkZFNWQM2aL8EjuXCafg1tpGJL9iA
nTR2N8gAoOFmTFGIDRmxUjvJukyptJkov9myiALwUfyqeqXNH8fsw72LVPkl/uNs
5brs/v3Y7Z8FtqPPmsrlDAkhkMWSNFwg9wv0gH5tzWagE2LZwfCnUwgcSP4zV/Hv
JSY96DlJ7in1xFQ6WBzGqOXrHmn/1j4MYOKmEOqL0gSAlf/9u4TkQ/lZAf3aUaY4
q8w0Mj+fnVasgFvaisiLS7rrCt/NS2GFIUNAi4cdX36vBUxONQIfl/YUWgb0dBrt
xJo6nf37ToXdSbgRp+mNneokBIDQvUnghZIowhPJTdu+F/Og0MKyF31vBhoQSYZz
eWyTlHzxWObANDAKZn9BNbZxubSNcKpos/ZgHDPWqqpjR96nBjxrscsrm6D+Q6aL
CAPPQT179MKtnFUW9o6qMydVebtVblzQ+4mCLBa7fgkILn0Hmaf2W9BzK6Nqwa2L
2mbXrX61mdZlytsTvdQlnTtuHqpH5f9InVn7PKgW7BXERJwHSpYyROhMp1YQ2q1J
VSn0y/7Ss1Zwk6r7biq8+M9JnS3/Zues7QADj2OwhKC5wmnTw3bbyNahB+Rlxc8G
zUydojGEELN3DxVQ4qkFffFCItDRzh3L7N2ca1znCSIZFssW0riCLKaBav0Ghb+y
kTH6jN6WIFAZ7IX1bqjRtIioI8pYdalRf1+J6eKRtYRUnfTYf5peQqlvLUaJcUWE
8k08WqFCwIqzIMLJlq00JzyYv5hWCQRXdAcJrBJFtyt1tesCirWWjRGz9QdA6Fs1
EGWiYUgw79ZdTbAGUxEfu8ytEhFKePbbORi3IeVIfOma6gUs3RlS13vLjPEJ6cQU
7uc28fuwCiVIpLqtIv04piGIIAq4PhNgZcCblEyInL9nekPMa+epnS5eEbLjinln
TYQBk7GNU+HNnrZ1+rjv7cgRCsfYF4vYae3B6JycOPcQ21sTK2JeusjCEdCq5gKJ
esdWyQFvd32Vw9UnHCaAtmfZz6lroPbmHrjRneQ2n1MGIoqZZgbJ0jxZuDjAgDYY
clOqy9flfonBLXZiWxDJtoCewLoqwJXM2YPTlQTsWHRPM++lA6kT/7Ao3tfDkFCC
iWT2c82E9kezv2V+WVNj7EZFmlMcZGRxDVRzgpgtla3e1rfQWKqM0HqovfWB+byF
hp0d+sH75au1mZYT+DALN5lkTPvgMxkoUZinxXcES5t2aBuL/kyG05qaG5Ge+bmp
MCy+YfkrYGhzKwQKTNGPiRSOKLP2dZgjI3zDtOyvpCqWOqd5nkyAu4hS865pmBUU
/uq9dkudviNhAjJCBvcvX2qb7GFeG3kI3xWOYhTLjrNwZSHwczUp3zJdacHZwghE
6bPsjF0RzFxxki7sQOBbrsl84WtAe34R5M7K7tPMJHGxK6Yd83T+SiQCgKeBp7vW
Q46J+EcLTzL8inftd43nRZQQ8zcmWa3eWFfpaC5anB1X6vn/aEB7/fwcftXDpDVm
0vld88KxkvmzPe1X9iUPsHaioOrh/YP7Kfm7cjuWRA3jdVcog1GNDYMhFPZLZ761
OlNu9ysRG3cU4rd9wJq05a60AFvOT02CAsd8j4CiDy2T03mZDSdsO73S27sfSiot
BS1YT2hRlGWODssV2gpLTOahcR3JENN0+jWoeAb2C+UVCDCIiZDvMRsAz2iCfy8k
wZ2uVXJGn32XdXqiLYerNrMLP7LX9VFa0zUuPYJRsgD8db8PycXfZr7LchIJDFjs
wLB7izP9riwG9EeowgRQbxW3mtwNxG6k92z2e73CEyHsSyxnlkdWFuBm1gWt77YR
7g96FwLn/DEV9/70jYfcuA5BBl3tqL2YzHXxRYCvQSOV9KdZgBLoA4xlJgucsdDk
GTX58hVRg3nq8iFHnkhJzR9smpI3ga+eAq5GZU5sMD6j5tAgtANKvA2g/5RkT4Xa
E1M3bosElbD6qVxzHQMssVjRqtHjGg9/uBB6+q1MNquPRhD8Zp2RfcTiuIDAzXvP
uei7C1HQnbFhH282o0cO1oRI9Fk3pcltcKs86v/7UHuPCx70UhV9z1hVR7u4zXuK
vTrkG2C1wDPgGr6NMRqucxPtAP8w15VvGcsi8F8+4DWMUxBn8uK34hDdOudKYVQt
qQNBfm8XiJqK7Vay2kiEJ5gnJc5YzxRi0Dohwjfso+YVfP01XLvs/MG7bJo90xkv
NT4pXBDIoCIZkLN1Drl3pyxntz1rHducNZPsEfo2D/5Z4aAsU6SjjT1iJvBSP6kS
7wcB/+XPn4IHl/YeQFuxQZ5pomf4YAdVFNctspW0QZ3UwBnSxWpW8ehZY/up3PNY
l2k0NLlTfJv+o2FTURu771jFZOzKPppTmGh0qoRVh2/Uu+MS1jrKHksUNY/eUo9O
cK3UOQ+D69NXeNezYP3ocCYDe74T0rL1wee6pYYnJVyN5pCzPEwnHeluErepUZld
+cP0qDKoE9EDmAsfr8YiKLiLu4IT/+sPgAdcJgIn28d+JjBDRV0tx7oBqiXU5hrA
8MfZNqWg/YIePC50g0l6Bn4HXrHQ+QjKj9WCb+D2krwgjVWT4jKqAouRgrf/f1a3
TsYAZvJNgM3XXTpQwKVKVc7BufeV1nJuACZBIkTbrkCQua191eZXLmjr1IG1mN+z
xaqDCZMFQXQWZi4D29/GwT73lHH6C8TYfoshCpFMKqmxBmX31UNy/wa7blAPL713
6MC1pEj+nQ16lS/GbDl8vPczxCPATdxxG5mbYA2HxQRWnZZ60ZiTmPAf0zr7773y
YM3U2A37FMDFuiEqGEA3uN3v4zcSoW8y471kv/I2dxVDFg+JWRT1bC16OlhFurEy
3kxxQVwy/nrZY3ILbu+vRkHpZl9wnqErRZ8nFGptxpQOdMbBrlMsPQr0zq4I1UkT
n/um7hJ2sebpZ5I72RTlQyrXgA3TKc4UkFa9+t16EZah3wPvu602xChZv8FEflYA
yj6IaPutWMYluGC37sm2eqXb9KyV1TCWmHs31rsiunDx7NKBU1Lh/yNmRr7DzeVH
3QdHt1jSfqQZSMq+8HbaA8RMlcyXNxuKlHkUQU/dkXlGdBoDvn1QJ9PEnHRTy6zF
rGq48T4epFqA+BjP2lCbh6zozrevwDo5XljYZfWFaLU9aE6xk8hm3SMdK/Dgvm/o
Gn7lATTZW6NIwyawRva70f/u8yuxJrlKw+Ib7kycxiJX91dpZ0mIznS7CZbtY95Y
FNDA0xIoOOhd72QlS+XbEu+BLU+i1RMClPr3il7fjo8Eq6bNxK+CK/zK/2LeF5+E
7o9pdpioYtYCWzDqWl1XxS+bQGzLzZvjZVUXeCbii0qORX8XHFVEOiJpfIRgoxXI
7gtFpNXmLYIzfO1Ai0ehyjlwpOTOONHvBz6ePMbegyFOhncFzH2tcbdP7HOKv+jC
DCnH2+M4T3ac+aVVsx/+LXrHu5pnrtc3lt1Y/4uCN/Du6g+Q5YCSpGv8Qdr8sPOE
1CgmqFRg7dqkrvb6JKso5/u3Ov70vkGNmwCj0yMdqFao8qH/bc2k75Yc/5DE6bWv
JqoiQcS50GrXs3z67xyrXtF6dW7SpFQNr5al9Iew38uEtJ8Vkkp278+LnoQao7HT
YjDRe+bpqYafWvVo3TbC4Iet6el7kD+3FCfrX3346tw6p7F5rW2ndn0lszET/Oe7
9dYPArN2kJP1Qo6dCaGJIuB6FoOxt2oASAXRDc/jBpuJzoumK/pQ1u++nnt0oNbJ
bv0QuX/dIJlPZuvfmEHqntAUOJQ1h+tN10QxgXUVTy0u9ovfvbKV8rhSrXkEnR9W
9r3uFS71qDOL/7tTdh9kl8Rjr3g/FACBI6Efl34+KzThT5d9m/pAKZB1bJ5YLBfG
KFVuNVzT54/0lpRMyu8BdsCoPCdopKJXd4lnrupZ7iqT1USKmK97YUAFrSy5QGSO
bODLPWHgsVGmoN3uqcsO2cPTol2FeSy/R5Ix3a4TbOw3nzYmuZdYGqB4aJLxocKZ
FU/NvheAnmR6uP7/vggs9/5e683R6cGYzDlG0gGRI67QR8xRpyXTSm0ExlWN53Db
aM2XLzvOn+uHSJPcj/ZJRBZIi6tU7Hxq+tlek58xDpMGa96Bv85jJgKvCdMeG7i6
Mg/ozhvJ915/0pn6wBRjFV57KBOAVyhPODQX4VjGfTIzRIqmIarEk/VgmNjOBCP3
ElXs+4VOBjGDPrSbJWzFWCDGv+1gc0iVgrvFGUGc/cjp2iVPPq47pB4ey9dmGDnm
NQnsEJvb/G3lp4wuwaErRuoWA/mlDw1UHW8wIwmbkzN/T1CJWfxp/9Iufxk36FsQ
EBRpXYmSAHwlzRQzhoWZHKa/XSIEaFIReS7NxRyyzj4iRv2jlf0YjLTqvVhNO+/u
Zri5oN3GCq9eS4z7w/srIwKCoM53oRZ5qTYJON1UqhI2K/kzhMPVk0AwlECPweS1
GIEKJNFo5Yn8klf01PqXJz8twITLkNrzxO4eCKqriWdVeEscv5WZXesdj3WVrgby
du7PBXKu1E8BaIKb4/9l0iUeOutbywzlIV39H7tgt8yBgjLz2QsZg9xke0JEyLXD
owAZE/uwVKVluBMmyFd/xDE4x+FEV+3ixLDUCk9YU50njBZixReDAsDxItVKi81L
mGzz81mDfrlh2Bao8qdZrGJzuWw7CmN3Tmj8Ls+Sl3+q6+s4FjZO5Eq+TIydUgBZ
qPtnJx1MmC/sS+B0zkH03qMZqJGOQ/XYyA2l8wpWxtlTzrqkNhTg28o0Jbg4GJK5
FXseD8C+jc+dKGouhcTKAIiTUUuWvzzOkkW8TohLYIxfCiJIk4oYTU+bmlVfpXx7
V5k9D0nH9Z4wYObQvFqFc4xWFUiqp1TTPwePtSnMkNVua7VqBjC4WCrClFr05QgF
mfE/6mQLvsvhVMly+JoIacbJSbYroBOwA3yd7KevpqE8/1f3rEWS9slbscBlM1S+
ffbfHQH6qKGNC+MjWWXQT8O0TWhH/PNtMqEQYhLWUtlSYkpR80jqwJytDR3uAAEy
q3B3vIgNPtscgdzdUc8DLr2N60G2YxA/1JcdM2q9XCWacgh2doMAitvlRlaSsWsY
HQETK+BGhq9sAZG5ZSjsnGdnHJ9v2960sPORYXYVW+iqUgmJliS3/IlZJospOyQg
IJ6xwPfCStadXBFyVQTnNpjG9Sq6sEZnPvgpzZtiF2m/naHIJN1FFdRFeosfOD2E
enzijs0S68SOrX7ZPop2TJU4eR5XLSkaBCJInkYGir5uBRrGGuz1qKgZ7y0WaIwl
6RuUT9NgV9KGU4bhs2y1tc7LZjsA04HixyWs6b5yA+oK/yIJxHeZwGBonWsV4rrT
s1G/FQG2ja+bf9qB6uLVBBUlVF94i6+nyAlSG2sW5hgVdr4/HfhDyTxVkfCTvrxP
8dCngX8kgcRp8Ud8+WIZ3i8rQbGmnK2Gbi53mjatqttfYHSDNpLiqLby1LbUk0TW
n6DDIscTuP/ExZJU4i0Gg65UVPIcjXY7IZVNx8mohbWtgN7KX5vqoF87UHIHoh/E
bq5n0dg+LJJIdvj9r/Abv0T5V7CqhEO8/myku7o6FcGn6y3s0QD8EQNnOQoORVyf
j38t5drQTE1rw7ri2K/wf4mJ0M/0EoiM8rOU7q64PjGT78u1Guz7x4jxoosN47Zj
qOBq4E4FY6MfENOMNQMu9q4aGer6XF35SJaXxngQL36Sa/SAFciviHvNYGjBF8E8
F9L4jXMztjOk8eJUD/xcodZ8JC4+gKzqTGUu52hq+BHzsZ9MBWplIqdoBnvR96+4
Ls1dAlb7jMzsT9vGgYL7OiwOdy8TUYhKw+JgtQRuXxv0b83VGFmrffzH4XW5Qke+
L6FYyHUC7a+sNDBIySfYSvcN4wMVtdNiFCMz9k/BkwYYEUO7DlOfSeOVGxyAZVTl
WioUtWuEUm4eOqosCr1a/uCk+IqH44TlA6a3dIlzZQAZIJ4Qb1BuwLx9fN1q3p5k
5AZ2CC+TWI9Q4ScSbKHl3/1t0i5317QKagNdykzw9wzmNy607t3oKk3YTv5lciao
WhYRSDkCyIQ0OpGqN+5dieEZELQTfu7MKsrQrH0xfDfbeFGZ3QvcFgVRIgKi1kEn
6BQQcCYXKrisxgtkHY37yyG0QdJsHeKdQ6PatPPoinaCrsWACAuP6DHGMnmq5TNc
mbzG8PWxzDrVUNVTae0AHL0cAd0CCDVp1vn8Sn0Yg48lAkTGhHF/aHS0LpFSxZwI
t5x3pn2ogDhKbEkaFu/kQbW8fmYfxq3u9SIg5n1ve1APHYjpe0QoXnbF61sLormH
LKG4avqdJermVxGsSRJotAceMklX0ZHPZ8yxg5SaWEMnTduy59z3983PcXMNYNO0
zmRLG9AQUXcLlwL2ae+kQvpZOj/i80gafx4IQEHysc1NWDXcZkLsRgkqg9euSyf+
ZqSlgdAiNu1YIAPEOZ057ISP0zUa6PLiwsUv9e/gyLL6V4CV5ezH7hURcpLoRASn
7djDAkUJM5LeWCWAGyuNh3NcNdeZLGXWN+DLK0lE8NyyKV5JGF+UMfLnEO6kW8OJ
WiYlD6nd3IgtV2zX2Y74rjednet44fUTGrae7Zg4d6TlFTQIgSef2sxqJvkQHK9S
cwDZKeMLhRXFILdyt/MOWyiqeJw0HUbkd+o2lglo/yJ4yA04hGrnoZmdbeVOh2hP
xH8A0W7QR1ZJGJENNjzCrWTU6ZIkafklig9pnI6hy4WcGS/AbBTQGHnP8mfpKbe/
WXCRP9Oa4flciZdK0uGiRyve5Kc64zdr9JpDixi8W5AaIr0Xth0wdBy1qFNVYMmu
ByBXdsBMomo27VRDSBxJP8YrKRO9X0rN8Mg6r6AdV6A6n15JoObZlQ21JURJDzC2
5LgU5OW9uQdNAfACOin73MMmWWggt4lrFOm+5ffhG4tVYxfkRuFNbaKr+hFDiA7g
U9WlyNPT79nWZFaF5u8yCI0CIZChjxV/lr0XUzeu9Wb3v+9DxOZZp8ZnpAIXFlHB
ENVa6XrSvcTEAafzAq/shXswd0nT3QyHGsXQ5L9J8hU++LibkMzN6jCUzBOQ6jcZ
YZZyP3TtO3nx4DGl5WpSlyNS3yvCHC8Ss+qHIVWvH5Ff1fKP7cX8ZEe1KKJ/Seem
cKr3zQfQgmoLDN853QSn4S6VeEPzybMumbr/00Vx6DaECsxSZn7IRqTbwafXmX5l
srjGmn/7ldaqAGz6IrMgH5j3TqrNFCOE2nSGPdwDXm/Xb5KduYHCZcfsqjsQPS4x
wPaiSVmumUxmSzJcUfkPQchzCbOQOy5pBC5/xcDvWLhj7GnQV8aB58X3W2ujPO73
ByuY0cM1DT/8hVvkvCUcBcgdri2og0/lpFE98BU/45rnpE2YFlCi69qlyqv629Lu
0Oe9yEQdemaTcKMNFQ/AuSgmr1WomjHJZsoABoze2TvXXdBAblFRhcUbSeyFnT2s
sMEN316zPEeFO0JXKT7kVe0kFW8N/dTZdpYiV+Z2Vtn7UgwelihLWk1Qj6AnGtJD
I7/Qi1T812J6ztNTijflpvgt9YdJKhrfTNsNCaYTwzfnFOn/3BEb6zUrdoVKs2uw
YD58dRTTCsDjsOh5PEkQpfTWOMAY4MumJWu+WlpPvfXdOrN+cjs9r3oei1A+r7VF
ossQ8+j7XvuPozB1YflD6NVqz7TNp9lwNRZYe1UoaNLpmhb+Sp2KJFc3hcISFfPr
rxdhqrrPbz9v8+3oFOlZ+TVud98WeDK+g7DhVhFD/KvVF6YQDaJkfe+R9eaxAHST
tD6cCQG9QETIjnDrJUuEDLV4AmJep7r3oOKQrHl/kBlGPkF27D7U9omXPsZp58yO
2o6basQzba5kr3+RBUgVnyI+IEGUSm0hFbOvQWc8Rc9kbPDoXPm0WjUpbZS/Nqee
2tgd8BeLLrwceRc1RQoJlXaaDUFzm1t+aKdoc+1RWshxz3YctZk3PrCYcbhkjQ/V
unnugn1NxtxqpPPrPncUBWmjJsoJSAk0auObAUAlSCEr+JAfl+qS4I0UDxTcSS+m
ySEziWk1/9pqiLM2ewNcDGvmSKNkTW8D8EaHqtW3SadEhfA8aj3wZuxFbyR8qcWg
ZDURw3luoFfVR7gnMnLm7TB+RvzXPrLXoiquCi3Ic4kvYJTRCYFh/uoYYapfVZRq
st36VQCh4gb48QesFhJ2K0cniriw7F8+E4d1/3uEJJrUYnMaU/4r934EE7oeVACM
O4gVdh4Shh8ZuZZ3p5YlpLIbFvvlj33tNYXzAGBRuIBvNwQvH/I06+bSYwgfjOde
qKg6gHShicCO1KwleGJfNivJGkehZC63ZGGSgYbc+0I4s7N/Tt9+MF14acmTMoGq
D9LFFiZ67//EwasileHbcrMDlJUzqZudQUPzMBjCMF56vYiKD+WRiaKbGOOcZArB
GrUBZ/Q+EMgEUmWo/G0XBk4/pWI/LVSZOrvelBPsys661X4wNiCxWB17JssNttqQ
B6pu188/fkkvR3iNMElMFYXCPCybAO0NRr9X76tRYGqThW0YyBKCZT4vThGTWznl
/cMzqgY/37sZuVDaVBFBW7fZ3ZnoTEa9OOqIzs11ZTlncc/BmqFmYmDA9QR8BNkv
/5h+o5lEbmBXVZwxWnO0qZbMbBy+3WuHgXA8YOpPSYVpL5wT88In4j4VWqgij0DA
2CkNdP0q4doNPsg/b4bNbwme2GA83gEn1A4xhhKFiV6uXNLOIEOyOUYncm9P2J3g
KxGVJ1++C5De/TA5OrQC8iB70490NRcITkzp+qQW7XhN7hwZ0uKzeI9bSlajKR1C
QM7VF+H3j137wNju80tbK0rLqrZbNe2CsniiRKRLjWRI2uNLsn7GmlwPnkbNyWFv
T5A9d3O3KCGY/WvsuZjxFhqL4Bj7F2YW0sK1dAZgQHGSBt+5lJNN+/D+6xMDwtVp
q6WaOSxOtsGWLMlTADB4oiWPFiKjoobUVA4vheyWZp2/Qpdq316P4amd/ZAVfJb0
RfCxahOfext8AIuTeGuIuWVFtgvYcbiCDWH7sg1z17bVCVNxEVOcs134eV9LW0pc
pN15iBumph9TEwv6Oz/oLeeJG/mRVMYCi6TaphCSorTDfEtkQHVNlalg1idzGIiz
ruZhK9cYBKoWUqS21vJC2nr4bmigXG4csZOVLpQzc1vpqYHyJJXRkJeXFFk7lAgf
3EogY8bFOoI8FMFC35WMy8kyMIaU0JA6nJ9wtX3zyvXvuv73QgxROnzYylvO/WF0
o6b62YrCf61vbpTwR3OyDPgy/wY20t9Pul3BCH4PYlp+6OUN/H2ZFAJLRXYV1saS
Ol8lCBBjnJ3gVJtt87ubcqGs27mCRXPy3ehCzA+axi1fubWj+ACHbINGVpxcN2rf
QtPVN0n7e43eEdBysYcg5u7l74ils+3koXYPCLY2emugBQX0p1CRvdV9Je2P71us
4Wjp+UVl5b/Ye+puOzYNbuiH5YiDmF0kvUGp3u8vED/I+MpA1+w7K0K+HbMJhyJn
/Gx6FnncO6OaKr4MYiGm2d80Kuv6tUsGO4nuz2n3vmCBggsHUgc/FAQkLXXN6JFf
4wmS82jetRHyTlBrqOap6I7zOZ/Ng5zEO32YOb6dkxlr1TvyLQmuTwhdQ9K0X+Rj
sA1XTwQ6io/AwHrehwlDj/G5JhXw3Cd3xGeOHa8uyQV7BN5kWdizi5S/kk6DQm7P
cta+58NUiJzS4FaxxqiDQOznLyuLeAYGN8HKoln8Geik+2pta1/RGdP9u7bGQj/b
CV6sH39YHEzMv6H1A1nYAd6aFf3xPWQRw/+32V+1VQv+zG9iWrsLU8hmIa1iWWYx
XLiFBVaLM0yvnkQA0YNuRt8HCd2JI552UxCwUiGL2jfOVgNlDqdtVbbGB0TPMYQB
pumQrasczI7CvPt3g+zixaLRp07f4BjyV13ZQvNsxw7LXRK8fk8PNfSnNnynvXmG
IRocdBjAJAk7VZjrFAG+sUr3x2LqCd/PKFn8ZVfOC93x+zOPJbn3Gm+LZrhyJJr+
mKvl9ezwwupVCM7MKh4+XnmjtYl+qRFM7iMuDbBdTv/qtLL12KvxtvdBws92e6xl
AbXaxRRzj0NvoKcK9avrEW8cLg9EjgTuo0AYoSYzuo6MkQzUPNIhCN0hinM2yze5
SQf9ydYj6CvBC0bx54G+iKi5pdyBRW8Yd+9SKNhpLLaO3/YbbvOuYoHkF6/mmKWC
2lGfwygXVylBBRg1IICmcKR6CxKoVbZ/DKczN7Z1Hz22axXuNipuxZ/qx20TNGEM
CsCxOt9Q8umQF/syt2OeA9dL9M5zcIkZG9ZfSZ0nReqfmrj043gcbtevk4qHEQfl
uQtBP0NxxCARJBMEsyiaIuiynGvMXHIZ0BSl0tzAB/UaaF65x2dqPCy2NYW4AXat
I3A7x7AMGIyNFpvFdsmUG36JI0FXklK44PADkAlVk76zNZe0I9fhiFaUWkf9TBzR
CYfzrmv210pHb4jwNpRp6zzsPDgHFEStR4z6rJeJpb/+5uKD860fTtCcqUd9qDzv
NF3dKfynNh09Mow1fEe/QAFrEZPN/Ud61Dwl+EnLXpxpa4kGmIUZBPgMV7J6JuFG
Izm3q1QUUgjiFe6ZeiZgT+NbufMWeqWl/q8Mt3KKWJE=
`pragma protect end_protected
