// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
n18/snMIdJ8fdK/A4p4ixniFljRg6bo8btyX+Byzlqn+rGpqGRPpxRvvWTr2
2ze80yYtXI6vdSQTI9d798wmLm6GlTS7fCuPS2bJA0CYuhu2ztQ7BMKbhiqU
0l+0TgfPI9nWNm5knlup1tKrLMPDebXibbssXU8r7BHVxTYozoE/o6psXZGZ
W9W5OY4ovHkCNMXb/weHAgWJ+JjDQUxcLwb4i+wVMbtNqkbrjFWzWZ9cZA89
Bx7wC18tY6qPiaVjXBDnjURWpnHBViagRurHgVXir0mHmpyAWBORw8FppbZa
keAG06Ze30geANgRAfpGgW13uRbeQPO34h4PoqAZrQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Mv7rlG68rN/hLJCoFDyE+BhoJQfmp5rKxduVpKo7Eq/n1gOhfHFu+d2pf90j
P6XIQkVJrEXL+MhR4z2cu9Jzjs2vJwRR7E3+jHHHTp96H5DFrx7C1GA09SZX
TZYygoauGoCSLrW0aJsSBOrgs3FyOwaVaRQ5PX/g5N1OM6aBMUBwqGSA1Tv4
cgyY1rebfpiVOF6ch/Gvfb9Viuns97v2tsTvOm6SiIEp08UgphVLVnNIQ0z3
m2dzq+C9srgXZXNv6PkS3itU5tmq31mNgIOpdD3+2DHk2i5dol/Scbv8lB+g
ByqkNb7Lta5BJmIQNA6bXnYPnp7kJOTYkgZn1ci2vA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
d9ppX+XPPSKRMhPN7effqPpNc0kDMKm5phKEf6Q6vh6cPt9rdblklhrPPIpY
fSNRGnNX55a/UhktvvQwnsvB768a5Xr7iUUI89c6VFh/AQXIbMHE8rgd+wzQ
l6jeds8hO5jL63miGNl1jZ2AO4fNWKHn482xFQhMgpLa2HbEf78GFKn1+Yf2
tCngpuwXuNyXKV0icNRDb65UvTgajJGt5S0ncf2xfhw03baMFhIJexf5nPJF
L9DmIcoY75MAOaTS/zl+x7Qi7old4/1YFtF7rjB29iHHfJvD3iX5wFR/PDYG
Tlaf8Iwn0/fblB2sRcat5+EhWeasJ9+UiIEbkkU6Gg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ksgWoAFKj+5LQWElqqdnLE3Bp3sZQ3KUAzjRcIrALIKimkuKEOA/RVI/61wb
d925nDF4lKEis9fMZXt72nlfJVtKf3xgxhMDZKFi3VYriy6dA5wO8PrCfqpt
V606RvpLfYzfYgfBNnrjEZgSe6t1us9hX3bFeoRBXmFXDMcymhk=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
ktjxSBpfoIku5C3H49tanCNfrbAcfAaSoheU9joukp3N0R8UCeLKHLFO9R3n
UeyZ7GZKiLxHFD4XzaGvFKS0+FUw1KR2sJuYrIqjJ+UgDHjdM5dp3l2sG7Oh
ks5kzGEUFP+3/enDtKy2Qwbqdl9c31eHgq5/iQaXmN+fguvKQfwxgoYKtWF5
mGySlEHpkkJUxWe3Oii/GjZX9n/Q7V+/IqZOmrnCqTKJnPOIuD318Do4YS/u
/JSh75cnpEHPb4d4d5SD6/7V3za07iUp7PLMj9KO8QiYMqjv1rCvqPkZq3vU
NmtK33sJEgyWy9I38wTo8bcR5/cmG08zH6an2Fo4YUmpdMcfW07OuJ5OOhwG
1JDsIVPfoKmLMPeg+nSydAMts5oWpsW0Mx4zLsqRoj/KakdwlVr9fhWvgPA9
np84mNBCL1icnEsYVhqPVlvlOVwh3Iv2VBVSCkTRM2yp8S+Nrd8LUOE6pBIV
XH/f6F+CWQ7pw4htJkCg+W2JzoOZnUDt


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
TJHYsRNxeZlBNSrFmYlsLtQZUG6QXfdniDWgpNsPkehY7kpSHcQE6bf/CPK2
NwbcJrATtfQsR5FSpM4JxKmqgBzsq9hCTYsaBuu2YqiwuIUZEQQXHsC76Nx3
P0wLdVTmTzmL3YGnrj8OdSYOnXvzBXvl526jipYS/jF3z8Q0d1g=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Fow4FwB8Feg1uqZdcwUVnQNCAZjLejbdMRex+w9RW0UP9Rt/QOZLNGB3t7dU
q9yAN9DJ8NOOKnsYcbhwAePbgT7J1cLmbDSdS5fzcsUVBBeqsWs5+6POuauS
dddf3iJUgxs9buZN1ybhUmNkXDD2NB2AaU0P3lekppttA+LkxeQ=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 113664)
`pragma protect data_block
3JMkQN7uXgF5aICwDbF2V9UwMMUF4mHixA7P9Zgei5RRT2vZ/ZZPs6CUGSIl
WicvGsBEfprJmYyIZkQqsmu6bcUwlHjBVIUvfSVOucd6QDBYjHaCF/nMAH5l
EyyckFBKawgIpMA71QnkT+yGxTf625YsR0fbjXE6GC8oV3ESOkPwo/53EqhJ
1yOMrU3pLbWbBIe4ffzMlEbe6ytQVEBrpQpE96KbPAniHmVntQTFgXpKS51+
YEtylAap+ousTyLX2ZcVO2rFE42fbyVR6a2F6SKi0taQ8fLUrCNsW4qw9gVs
fNnQIoALm5G2RMfbxQdPpZO/14fsqwCHwkAvBqtO/7K+el8BFY7E9ZZzI4iF
2ce11LfRK0+VSxUz2xn2+ZK3UrZHRTO/NEHR50xrH0mfA5KGZGTcrH+Xzh1G
zEorlJ3duqmwh5Wp5jvHDxjDuHJZsCrUeh8YeZ9JWUdEjpZO1KeAyl7XIx/Q
Rf9WYDGfZ7J1h8l8vR5+3ZRW2IG0StWNW9QRAO39+Dy1t+AUWfRxWbqhXTO3
/detwhRxjx9kuOEbe09QIZIOGOKCNARHNHnphaWu3JyYAsVUatmOAQeBcJlv
wV4bHNu90VI9b61JFcADgbQyPZNymMIXAImGZ8xKkEdoLuDbZGFoZYVjMSEP
X3xQIdFq9W2n4IdrerfmAZ8AKNHoB0PyeOM3h4zPBVNOsubhwK7t8yg9Wu1K
lr1KwhU5ZYqQcV+ZNP9tOt8/wxoyiFVk8eR8gdZ0o6NJpMf6Mwts/UwApi/z
xQx5zAuFI8GhaZPMmQH5hQfoqOy7q00sg5+p8JYqxpfrZ6k4XDn1Q7UzWgI8
ExoaAM93HkNeim3Sj351OxBTHYM0cTgEnMlt2iW8Nvmda+6XBWCPS3XLfJkO
FgAvrOZmUU4Wr5QSduGIilStx0DADw3B6DDwAf1g91FmWLdDZgEKM4As64Md
ktCQozCkkHZ2reo6hHve6KnhudoIslebydxIUMtelktZSMhhGR1kYii1ZKl4
5oh5dn9erBV846mEY6K6P3SwZlO1RGJYkdXtH6B8Mjg44ntkAccHosL9y++s
TlpU3cnFM3Lx+7JAOIlaTWGq1HawFd/642q8JakHAodC4wzyFUVEUujEZEB2
pWMdjb6aeQnqdy8Gtjo1F36NQsTVTtAEIOJ7smX9B5O4jA6V1MST+BwotGVy
x91sIw62KNx5lzw75cmA+r5uXjwj70HIIxzqwizyhcFdBYU7RTLnsDxvLNTY
QrVGMMRg/BEFhlnBFjpV8Zs13U+MBa9YBJjk1bMTpWU5fcz3p1Nk/054WvAG
qPkue9QtRCxCiaY1UkY1z8hVwA+cl6BRM2zmxy4YpwrGElv+R2ctevTUCLF3
4YNlqEr/Vj62NIu/5zzE7e1En1pBqpGKZWoc88W42O4MeFJFPHl7i+l5YlH1
hJouHH1wKv5yTcqqrzab46sVJ/ivJh7aWZOMxiurYkkGuMhsHYNo3uAXaV2z
1t4DHExca4vDbGxVB6dub0g/7flxkF4PhB4ijanOmzYxVWWVPN6KnNQ03ogE
try2futnTqm0N3DpdgTLnrP7vumqBmeIsEZaYOBREm9xfzUanphyqbGJFaI4
URl4OPh+3t+utiZxom+GBT+EfG1Eib73j4oIGOmSd5Wa21ym+VcxiSBHkJUc
aTJZAOOQO6UIYV/dAP1x2w1PstPoBN4MkFYKZV9yi1sgK7nMfMHnk8KCc1/C
/WyU3hmFQrbRLedl+8V/G7HB3nlUziGLAUgz4UF9lSUIyLAjOzJiPdJnzhWp
wGWbBfVwcXvjDI/KyAdDJZUXNduwQTXsj3ZgdiE/BKjzj7bYpp8hu6P5c6mY
eFH7+JDJSQQqQUeKgEpsQmhjAadIIPNoJgdpJLHWgSCJDdEgXTcqeZB/Gqms
8jZMEShgKgVPqPwtAYh9tA0lhL9zUxRBrSzWe0qfUT6cpyrKf90Tei6fc8hb
6rEQADBqDzm6Ekt+wUBKAeNEFL03Ebdyga+sZZbaE6pzzQrA1QTJylIfV/uj
B8ze9TpTlXkAANgduHpI0AFRRFXGt6TNunufYr7+lgdGYd5opYEHMFHJ1GKO
wZEzrGyTqiBvKtNEub3Z+VA6RQBobLyAK7hvHpbI1EJaP6ayC8mzRFFdxYQi
uNwx+j1IF+GS6qgvS+rraODQD46QiimN65GJF0pq7lfF+kBYCnl+IE0piqvJ
jm9hlpiP6g5Och0KQ6jgkCpC6bI0Z7v7yzmtVumNd3TbjM2k3Dyp2cGSBPqM
+8tkmwJ12HWn4qTCKhcqVIvdfNrXhGPoxD+i3yuwLM3gj+UcwthmW53Alxfx
rY5iz5/LWaKAQw5C1YCyG7NlEjH0+wL6gLx2p1u663c56eoZB+0TF5nYLxpb
E3hsc5aXgNnByhIes7BueP1stgoVgVHc1nipffkZjWCrZod8wQ3NORhi/bLe
K4en5DB1sh0arjnT6RGYhTWkji4NyKOlRfaKSnfvfr8cKbFD75Uzo4eR09rb
56wCjIuOViTlYUMSIkD5bRVVByHMI5dy0Cc1Mg51rAKGN2Ig7izT+dG1SVWH
7AATD1AX/f7q1ADUIwqKvDGR0SJlk5lDOMbS/TdQUTGnqKyinrtvNFhsXsw7
uLw2649yqky68F3DRfVNMaNdREWjfp+Jju/psiLnOHctKKaGy7HfSTWQwS86
ufZJIdXhUpCoLgsovHPdyPOI0hVF0zdubA7w/YkYd3xXneXDsnYOolaG4tUL
Gj1mYTT+b+OAMplXObtJa0LYCkgDSsKSsvH3FOb4nWYYg9MMq/wEZ/tOuPIc
lU8b1iKq1vwnkeHKxfEcI6i1TumAWWUguCbKpBatXcvxI1g83gmQlfrGwv7I
/3CIz5yh9hMJki33oeohyNm9x19gqbtQBni9Idl/eEWkg9MKHLlx1+ELW3cq
5uFdKMyaszq/grPOJ+gAfuy3VbgftYBMP9WLrvfqss6DKi5JqeF+qFh1cpBR
bZ8wANPoSoKv/aiae0UuzvAbxxopc1JRY4MYGWDVZVpjqPIWOHoHvQH2II3+
CDthZpcf16Zgm1jBd3gEzdYKTal3Qeuo24G0Ypp8omHHbBJjtfEsrG/glmfe
v8d0j7NNkXgaD7K/5Gm7WsK09xFaYjs7L4B0P84Jvle2ZU4xTGTVnjbUdj+c
On7lIQtVVvepI199dgErCdsPhE7tx2ciOQ9Hx55RXhWfrur0DWDWuekTraJU
FcQRwCxLoe+WZBj3y6NCPxQVAB3Eu4mN74RXbMyD7dfbYYM4QR0u6qa6IlyF
yBMY5nPoPeB1I39FcczN1N1Ol5AxaifHOu3TvCzfDp553JMSlZj4z0SNxu3H
Q6uwY9z8i96DKBATRF06goHKqiwUDcsFaqmfD0s5FF0x2LTY77TbUSCkSvZV
26UXsWklFC8lOequNjvBhoU1YePwBDJCNgqshKvnYKV7zaBsRrWPZy7DiJ2p
jeE6Fx3ZwM8wQ2yzPwA0DzaEpKuTGIksWqYIp9UQmTAqvk/yhEHWkKgf9jgZ
gsP4cBzRmat66AGBoJLWx3zc8oZ1YngmD0Zn/2QjUM4UlbDXFxN/Hxoo7JzB
u4WTBWo4ox3GlxuYwMTIGEhZH6cmLOXDPD88iybbofKirHnxaRZ8ZIzZQRAh
FkSK61nzz2QzoIl/38vVOLCb/pj4nrGRpnyVXE0s9UW2J82aGze8rVOwC3+s
F+hwDsxqKlstPoWwHyaW4cJ1N0lwoeMHqJs751JGWDoBlxP3b7RjfdbNz+B/
emUTLwTmZGBL9vdhKQnMOwS1nSmTUXCmc6eNVOnIj7aDiCQYf9HmYGpi+OFd
C0BKnaU+9d33Oi2HayDf884X0BarMvGQY5n9wfpYH8FHqH3zjv8YUOs+u0si
Pi947weXamJdLQOtMf/TRbnIJZhTx6MRhN2k8Wjvw0xIP+gvPGRUSkK4LlOD
G+UGhtTlde5InQ8ssGHzerM+t2FFtbXkSXc8WXu/zuOgQQFrGzu5yU2P6sao
UALBvVug21z9wH92xiN6UUobKAZT9d+vejlMwMusdGcY4hBnWNJenf9yKHTF
bAwLDl18qHkJe+oIywH11z4fkb0XkogenMWEQ4xW0j+c2p9qqjPqXNEEmpOO
l4TRsCO7ruWphIaHmcKZOCQHCIqbnyzJ0qK/+wfatA3UKXx+9i/55DCxFdg2
aAW9yCB5uMqkBvEWslkj2Z2GdjzluE4HmVFsmx2Bt0R6T6xmA7YaMpxojfHx
4QAVXN/PDALG+noVvMXeGJXXorsfWmDr8n6pDlgdpL6XvyXpVoKvfyPxS+GE
AaZ+WxDPTXJ+L1B3ddDWrbvZpVKNX4Xj+FuC6GmtoJu7BFtdpAbVDVrc3K/B
N4PpEDrVdNoKumKujwZLAZf8HAp890XZrltI8qqPYqN4Vjy/PBDOmOekQN/T
uyAsKWIKfxot91GDOrbA6L8M7i307xER2yIXRA/8Dis5i0D0RWtEBLS3mBrg
4MoZIga/J3Pfdx4+IIua0mOaMD9522UcQgSBsgkYm6l7kxE4148TGZQg+J8A
6z6+X129DKe923yrU8jdsHTiKKp0au5gvXyDJiIWD/ok/KMF3Jizyamq03os
mVsK4AepP3sbcw7FEJg8OKLbydSFMpDhW6012q+fGm9+vo8RKP0Oiwlbzk+G
+9zbh/qlPtUPx0LMZvV4CJrg9ZQr58++dHwQiOxW73HoqQ/o+CWOjdwqwv64
R3roHr59X9Y2d0Me+8z7Yvh2dG7Mv/3tChPtKATvg/3n6xqKSquT+m/xr58P
IDvfLjQHx2iIInIaG3aqR5msSqBNwCBZcQgh4p7ELffiHFBd3NMepM9CEu0D
x+4BwfFqg8moHn5uO//ocoxLIcaPaedyxNAx26z88iUq4rV4QAkZiomPS9LF
v2BhL91mL/9rGYI3jf8f7ZAG4UIZ/ryu6gV9SHjs5uqHz9J/oVxxgSYiWKLi
SpNPirfnvPDgn2Yy//0GX/1dNncmBTKUWJaklG157eJL/aQ4Y1ZmkT3P6liO
XY3OmmJxzn/r3njgWHddidIIN9o2W2TvgTA/YrMaTHm+/JReXntWzvHwk8wd
jEo0RVkbjzIntXK8E6apF73NLpSVwgO37bEttVvvPj0hJQH2mO0w/HwfWRmp
UiO/nTbPX5qvsXvfD9+JlrvTUYAH5MRe4AP6o0bIsEBNhUQiRNuD+Ds+HOZZ
fygz1eJ9qgNHvRLD3DN90NVXrb16cQfAeqqMpZH92gOLY7D3VUuA99otoS9U
GcSQ/G4XHeVN04PhPenxccMzLZCSiC9ouX4wcfjqRCFo9X3EZoUP/cofeZVE
kfoLmxf53z0WfLfybKeOtC9TMsc9xHRkcWrRCyPb9k6XokAcfYKTIaxKuryd
f1kcPTw0NkNKz2QgUa3JoMfRSxBDU5ZA0QNXLLyGC+4pWSxrzJ64VVRc/AJ2
H75QfGZq4JZ5ihaPws4/lLFkVvY+YHabG0uhtK7dWpYrUcqlhRvrZvngyQFZ
tnm++nl13AUpUSwmKFiJrK8najZP4S8sJerMTfuq3GjIEV1UpOZQYvfPM9LR
5CZEXTeh90HEJ6EFmFVCG1+NVwhZbEEdmixG14y4+iny/EyFpBAQbgwBeH+K
B0B8m59JzAVx/53z20ByrKU9t1RQ/NX8QP45jBWmZAhRO8pgqYkpljhqt1xP
a0uBVOtDgfxHorGyAA5hrzXez2p0ugO4CQsbhBPKjqvfyuPxTq4257V8R2ot
0e7C/NN2N59iWQZ2Hln7ZwXeQzTT4/7QY3pVK2Cmscz/As3HX/FtY2ACmzs3
X0hMCp2DwQuW/vxKJH+QMoK8ZpO7ZLWnrYVmhjUPgZEXpuFdR/uVDtB0NOK4
qjlcoexTmq5Kr5IAGxOEasxmn2ZqdvzTGbDAIe5ryTyBRKm9/mNRTNpdUNMH
WakZHlcWXkO3ixvH4CPaZ1tFptvx1GEJMDB3oNz3SrozecKE2TCEKJcs1VI+
1vag720PmiKF0f1XdPS19nRunxKhMX5vO55j5Fiko57r8qf092ZJoUnIXdWD
Nf4T7TlN3mAeA6JbhgxIx8E7UUqKuP8Fot1tplV2bqwdwzZJ+zNHV85TkBmy
uoNmpfKWLYWhTzz/AnowQdDIiTU9/p2YQHpJAfqWoM45SkDwgkHrQRGycKpd
neZhSQFx4cNxjOaK2LZQK9FI/btU29+GLVguVpRVW70d8xh8m/TFiYgdPohb
dYLOmxu+X6VJ3iWTpq4L9yCih6tHGc6MA0QHaTZqdCPlCRrmR5gbSSUX0kqf
7q5KX80vq6OEJAuYNvPX9dvWyuGiIVIqNCX5K+KyVRGUAuLc8HluKNlLH9Lj
VEmWRxcwlO0aUnoOWDSXofc65CRFWcW/LVymZRg+PdF9Fds+KaVuEDJ4Q31K
VOIRmgzAvXTXlZILafLeVFow7z7RJBul1BAcQTQEloacOF2QhcDlNB0OJqMh
3rpFY6PGHHzUhYRftb/0i5m8cgnoPJtXZmDS1iCIbskHZDtGewFkNQ+Qeq3p
q4pxX3qoyB1i0n6njizrChmsmNW+k/0kLTHBXfTi0QSBhwmy0yrBKbIxAa10
/OVr9y7lKn63rD8NBOEyQWpstIFuiBYIXnLuJyAFqiOG5cNFF1D68waxDRJ8
85sP5SxiZje/cLSHc63zEc4DwDXsMY9Ivm1viZ9jyqvR+25EBYmDYLU2+zC8
tbi7AhyACdrBx2eqpE0D/GbX60v7B74g1S1eT6LU0QWM+1ok4/wr3yhPt5Hd
ik73PqsGsCejxOU/fUbCxN5DESih4N+SxG8j4z4wQpmR3I0D0hV8u2cW299O
WSPuYEQnUNIHToWTMzjIDOH6g/pvoTlOfAli1Y/NLcQKKQC6hEzcZnNQ9VH1
BCncLnDUntqYmr/gisI34S+kdr5//aBrCqgbAiOWRZmQgTm0f8ho/zeJ1m3X
vLwm0NZV3utePdIKaiYUEBZaXUEB2IoOoDruiHg3m2W56aJRcjQ6XomXawkP
n/XAY+NdBjjJMCwcxwLSpw2BmmBReoIm5RHIs6y2m17nX8BoV7uAqjOQFFHw
NZuqbKf4PW2azoVnWeL2rVsp4O3E2/JmICP1G5FrbeQsMg7QB/XvpBwZ1pci
WIg/uOWcxE8P/Dnk0a4dGJOiMCfU5nfpG8uWXmmX2rQNaQw8iMLZbFN1eoaD
fnR279zrEX9mJ9HKZ/5PPcGZyLmkRUN0AAVo1sxgz82roEOPMU8ZO45JF1wg
sSQXM/mUzcbTV99Fn9VNdWtcvu/0IWPi68cAbA94zIZ8ryEIJxlYubx9PNrS
fM3TqfcQyKJ+w0zdrjpFFuYxeoaaYHjRSbm7aX0a6ac7YsUGYiKBuqVhPcAq
hl9ftu7/tqMUzNCDS8dFcZmDJ5dLECppka7hjj0S8DVmfEFPuR4DSQ1u3041
YM3DE9YhbuIvBLlIk3fAvbCjxP4owjMn1quZe/vclepak8gBdSApRQExnlVt
MU2AHmhmBQyZRCkfMV6lzBiwvsxlvawZv6xqkzdqpqi+gmP9FGkylooKJkEz
xdQy403I9Bm++CNUTQTxxsTGWd1RqkJYI1fdASu/Bl8wYOUvo9Ivw4tmsmcP
aHvhgrDxQG3QlrDv5HFo5IHjFIjwA69bsfUOTYqHo8JftFkXl3E1eEaCEzwE
J3V4nsIfhkEp80iqWh7j6G4UxhRObn/fr/JWFWIxq9FeMK6Cnh2s24Y2G/72
5z485DYYF1LVoYw09bwpNfoOHFZ+QJNk+p7Teozv/1sT1rYwfGN1WAQIl91U
rJHMGqYX5rdJ7/IBQ5tbtnqUycInHzZy9uDUO5g/cnDYUaqxCuJBmQFYzIyZ
Tt7ucveyQ9g2LNf9NTBz1aHW17dJsQBdPMZbORpCQq0gGW2D6MN2X/YN4cH7
8YZiJX/OFnGwSmghnNMT2+ofHMf1wQTDhlp+Thn8ViH2fqLBozgDNbaR/QU9
Dc1OoiNUznvp5hmzVZ0D26Q5OL6/lY4XFKJUw+/s5a0FDqsXqk+qyICppwFn
UzT7LV167dLgpKauPC52j4y/0yZNapQHZwVyCaBQw0v3EUBUVw7xDcOnE/Dj
RfwVeyRb3JBZIW9dbV72tHtD2Ltq6rOR6xWoUgoV0bB5HGCTF1oa/uCUJmXt
edEl4h470Tht2+V+buP34p5HzBiFd+7Q7H4T2M+16/AoueQCQ2PdwzZDaU3E
TtmWwcf+T5ekuOxZrxSeP39Mp0SBMlEVWADaini5ZxjP8uoblQwMn9jdGF0R
hzgqcHYp7bUGY5saUyHDrNvMNhWM8dtzUQdXOhM92OKKubzaUWXGJw30euZN
tfx48RyND08MEIU+OUxXxC/cW1yQ1Fjor0dn2BxcQ4vF+2Y2qS0fqE2X338l
XnuFtJZdcpyxvdlIKDNmihaSw0s6O8CAMU8wTb8NEL7UGoKlV3w6KDWQCpzT
ByMswTBgwOt5W32aw3RVYK3IvxmJPxo5v+IVgOvm26oH+Jg+BlsF1vW8xArl
fFSwMnKgtj+fn20Isbzr2Ki4hPLA4TGsN7It8PW2LhUrLmlOKwA9i8diGCVj
+YiycKmd8wEdf0xdNB6EuAsENm2/WH/RkA5JjlbsouL9YkCXaQfVA1qBadj7
Vez/cFNFGM/RYDBjEq1H0RJ8JdbRqZkoHtV4z3RAFccfx3/Hczr7/72giR1N
LYBMEmccemGlidrxfr3pKXHQEL70TXjquDTXeTSuocI2tMC/KXy45H7p7bYB
4ykCR37/61NcgTlzJJDrwGU5i++tOCs9qvkORDS3QRbzxfpjMNS/3sIMjmNQ
WYgW253cquXr4X4agVzwVm2tziQ0BdHK44GoISL9iJGvkfPmgA6IRnh7g6gx
nBH6hug2vTtAUBjFw1qikrtHYiCiXs7tIt9t63K5M+wq9yOqANWRtV/lGznQ
a/CTGZgQLtq8gttVS0zBAe663FsDD01XXNqUOWHBDtP4vsNn50vJeyUpiMpC
jt/aSwxnfjXdfsu8wKpa6ft5tT1XZjtxBECFv+kQaEpifvKXMCQudEljWLEz
4JwMRtUHrtsw9kHrriMjIa+v0beXUfAc3Zslge6o0JHDabU+/O2xtB/tn/X/
GaRTIHm76qeBcJ1uAyQ6Rfg78Pn35aiLYcDWeyWFtPkaiJDL5kLqqKQMQtEo
Lq6ztBfrs3Wdqv3u3FBLVcYJYxIyk2pa8PRJjgLphL2E7b7W8RCnAlq6Y5f0
2K2Z4Fkd3/BV+etnYagwF7bRw5yfi2xnfeTRgO4a/GOXhT4ky+Dbs1x/wqFC
GcwDUJvzG3xYfXPkV0wb/CHIjaqUEjbPno8ygXASwYiFXDQ8dWuKpkAxRGkg
XTRujmN2pE55UbAKB3ZJcqI/g8GVsn5KlV2WxneBNjatTtrttxqyr9i5TrMp
VcTeUhIkdEQg0BmHWnE146y0aX13WrPoWKzMbkHBJ2+JW8bJv7f0vQtVRbIr
NtHXWL3YGFZ6WF413oqoSPuIYr6Exyg/vK8GWHwhJrR2IGT6sL7wVmumPKkO
vxJsdPouh3P222rsY/ZT/eWsraAOt1jokKx4UXNrXpQAfMdyNiJ7qaIC5P1d
C/bNMX4f2dTD+NBceEWmvvnbScXkhshQuQGGtiSUHDkZdcDtn486m1GNJUrr
INLZlQK+Xr/48F0BMIGIbFPyGrd/VHjNf/DjHTk1v+N8pVF7c5u/WKHeiIA2
xtB3QMZyLILvmALyR8QjqqveMh+lckJO4N0ROAzjF37VnCSYwGKsiOTPFiDc
ps46JucjKR9Thjm1OV/bQP86HQ05jozY6yEL/yyh+ucKElng7vtrrwERkqFp
ZUtS+q7MEbwBhTkyk4IgJuG48Mt7XKVKwfmUaotQH9xYRtDtlSsTjP/eETfH
0t+5faUPp0w7njqD6U6KYxrtyq7Obo1gsmiJzHg4E2azy57ohGnhJZyexEa7
RiKN832mpXJhkw5wI9auSjQOHU7tfM/IaHOWjuiNkuTd0kYL0jGbc3/zkQae
cYibYtHPsogfvEHJ6d5qyywe2eJaKD0EF4DqMSti8RcXbeViNk2zc1DwxY1Y
oBsui62U1s/OfDkSl8gihya2DIf7X+evcIVUiujbbrePbLXdXB1toYlktO6Q
h4oa875ZJIKFV0+wM2reILlonem3W020r9ylx2VX88E57kmt0jhxSoBtjoX+
mq20LyUxEOyip0w5/R11FhIe6908wBNQyEvbuUmknKH2FB5PyVrlrhz2WTSu
BYvQCx8ZBNv7w6ZttktrEj8iZvt+rLAq4XewzvHM3iMYvTikgkcf7VNoFlYl
kKZdirfvvECZxzzmQRCOWBINV8egCuX+jG3/pwcjO9cShj82/GVfpqciFP7P
OrNUchGJkikWmh5dTuMOJpUfIR4RtS3CJFpVcYkao4rs8K7cgHf7O8OXI6Ex
/1GQDonPSdtFYkccx+lO/hUMe1VozJsr54iyWFSp0choeiLCPXwk0vs0ykuo
3msVeHkQLsjqtLCt0RuD2zLmnTN0G/h7XBH4R7x7LMNi5TFAh0kRVNp/SJrJ
IHsHjrMJ5JbTtLaafeGhTbGhG2qc6Is3bN1REyY7Nfa45sKi9Z7M0tjgkT9s
BInuXoWZEDaZsMQFUqiIenvjhqwu8A8I65ZQzFr3gNL6a4Ez23AWw2+omSjD
yYIH69NgKO8jCWJqQ9MKaNlAbju6cyMEbCPSo4ePW78gcPGPiU/vLs048Gn/
TlHX7pJ9Q2mw+9fEVakxoJk1qGAfvlNPi7hTVYak6HkF9kIW/MnFf5Qnh94Z
89Jzp+t3nSxgK5GlGCA5JVRDMAr3879M8m/FjC5jjYpWAOcR7d9edQ8rXd9m
G/ne0lvCNRm7yJSOE0wUncAtynVnhcr9eZIgpRajgo86UKvxOFiX20ge/vGN
7fMieMej62yQruVSmOUurG4mdpkWU5qqq/Z+YjtwmdV6adsb+i1hmy+/QYAS
tjr+tDYoBMrwDGBGfL9eZMlPmQkyY+xb6Z8rLXSvkqKGHgED07JLrgS6G6LU
zDWeRYddAsbAy7Zlne3M583cJvEiWLvQ/owz6INXusr2pA2PDA01Xba3Fbxd
OCCXlLk7bgUyrWChg6mcjJXFgwu+QnQQuQeuwP83O6ubcAy6J/Jvr7hP3Dn9
zeAqyzmyDI2fY6Mbu7oenkg3lEoOCqyHBMw/Tgxl/zuXNSYfk1UzKRASHSlC
NwWmXr8kmX6lliZ1d7z1ELuEVqWMnBP/r7cjC6eGwcXMt32+5amTsWW1M3EK
hDYL5PK37Bgr2pYnupmv4S7T4R5NgiaBAkwFCcadoNgKAG2foNcd6RpLTNWb
QgVRvfBW1ioxlRQ2jbLZnX2Ac2GxCBjY/Ax6XWaccKDRsN9T4zPE12lCqWZl
WvN09l6IP7hwfVpg7Bw0yQDoQhbR0KfjaDNEOp7tckDt7ed+ATgOl7TbP0lN
Xsrdle2WkzL/B19CexT0sSSBpSQe26/OzsqDgzm8E+CuqPfXlk2PzZepOhjF
H0j+Gh0yMkXYWHdwh/hj0BPVLEtr1gjTo2JyR4p8zTjwtKiYsKnaMZ2Mpb6N
au7IgTtcfkLy73KGOpLzhdYTn782/q0Jx9eiGgGayraRCan/4UxJgUsW5hfM
v+oeMDSp2DoFa8Z10JHm9XFv2vcU+7OoR3Z/kSIQezSlg8bQxDkrT3H1xJUe
qMV63lIPKViGbY2cjkj88LHfN8Lg09mg3VJlXE5wBUWh9gtCa+LQeVpNE9K/
RaLwFS2jPuMIGGB8z66KMEMSpB2U8IfRVlS74huPclptJZbYma8y/V/RaGVl
Id8tNG5MCKx/Bz01lEt3+5wNX+HT9odTb5b+faBp5L77T43LMKTNj2FE8MAR
gHTMnMSiXzh9Z0GmAHNaw9iw8+BG9VqbQLUusdbFMZa4rF50xJiDmHnGusVg
vzumsrI7cQQNqutE2m/XwD4h+7/RRD4yLIbnS/EKoJLD4iqnEDsEib9LFW3k
zS0QauVBRg1tNYW4yY3j4VS4N6RUUXH0B3bikGdNcHNv9rfXOUrtwuf7B540
96OD+QduMbE3iFrQoqDucX7oCHRFeU8/Dj8vec1X29H2NqiE6rItDOesQOdr
TWXYiaWb6/S5JD1zWBncsHoIyu9BvZ1PE0GbRASyGx8wavVS9c2/lyV0fda3
2nQms3XeumFAAOpPmWUD1Yly2PvJFulLOfkXdSepnLBE/YAHrRYa5Azvp+1g
h55wzjvHV6w9wY03yWT54Yvs4txpHwHISbC1ujQqkPrgNEo0N9DpnY+5Ougo
QBP7CPM8SkjUaUy7xqfuNPDlZF3oMJANYai3fsQcJUOolqbodxiG3q+yEqgd
NmFk3Pw7jS+h0h9bejDXncKjp4MQVwg1V4vXIKeu41Cn3PqMp4MZcshBrqPH
ipZI1j1cnpZU4Y1UfiJeZZpmDMG5UW+hT+b1TSQpT5YYCnKYQuOZUpvsCH7a
M8SwDMjDuASbZiRD2sKF+3am3Lecb9T31RRgMjQtSTHyG78oKI7RDIX5iPD1
FX00yijfo9JKY4xVh27qul3lIytKrPXcWenWXcGx2H8tNzf7ba27iAEY7cDY
upKyagjJ8kJrYazCNK65ZjtYQIj+eLemhtATI1QutxHShPq0bUR4Z2xMAD1R
m0M1ubBiPWu9P6REQOT1OrzwOSwjW2sJdYSzz5iu1tlSGxm2D1oZOK5pXXBP
R029dqHUqrzBX/cGcRnKIjXaOIPPKqTOkYuYEXJVBeY5MSyM1IMIZ/4URzsM
Y4bIrmCrMobegVeZ/fiPnQuvShrMMkctbdAhN7kq0aMJKNjqO+NTAGFwSSMB
9WAybt/s0VgOH7QkkP/kYmvXLC5amnOwiTB/qAz3Oym874tc0vNfhIGkX5qW
avWaOrSZMa5oB3gIIeBz1ur1A2Ccgz6r1NRAMTdtFMldCRHDA5ICdotbXJ51
IAZak6P2EjpzzVekgMLJep0Ebsho3Fj7ZwqhIIHRG97xRbVoAyKi7OePRrWV
NsvdgbnSMtZg9jp3V/EmHkxdJAL5JZDpZrgX6GrBE78HTdPrONvKgRpIByAW
xaseJHRcJ9yDobynYBXEuUKDWR+zpW9nT3O7qEKoyDhkcKI7VKV+4r3sL5aZ
jdubrheekeDoCRi68O7fKTiBqZq7DiGqSDhPV3ClRiDC80U3TSQqr49z/Fv8
eAivT67LWNaU6LS0DbVQm2z6vb1qKYrxQhB5ZGlJxS/NcIBUZMA4DyC2oxQw
PZ3zJQ5JgMQK16rjVE4jSxD4elH0Iq4T9l9cXetMohMKEKgKuukXNdLrnVNP
0sftCjIY3gJAxWF8/3zFkXUFEe4c8/rsYda5UX7upAq7C4zP1/yYA/iEaONE
n/jCqM8IvlQV9z/Z8NFbwyHwrOh2vnBZIl9WSdnZMixp+n2S9mxRtC5MLcGQ
K0exjUMyuV680IrWSu4MnPg1cCUNUO29FsFvTrR0xT7xIbhKi3t8aQlq5zv6
2oJLKVT5A276nWZWPwLug0+YhBFuiqwphSzqTncWTZYq5qIn0Y1Owd9cqnop
YI6ByIxX0VdvfPnkfF74HamjKVsah+fX3ZXrFvOgdyCJ5kPH1Xvr5iJwXxA5
tRu9bRQ1zEZDZWtI/oXOJXQEZBagx63eRWtGbhUHoAIEZfyHUHNjjGLBw7xr
EpcszyCGTPXqtqyUWrxQ/dhFxdv5qKW5LfuJnpuo6qhzTQF9d3xo/snMv77N
QjJf6kKwgdrzVTWrrxZRQePt/ka+EkbSfe3j9afOYMnSh5iDL/bU6PsZgIDX
mli+5cgHmnCvc7CxIGkDt3gPrJhES5EFUF2rTS191jFI4Nv5Eyn65tQi8cTD
T5H0FQJGpd2YFnnlM3Ks+f0y3Eoikn7tEWqb7o+NZWvtFWjelusJIglMB+hy
SRuUqZJ0cNQI9DXbmaikpARl6G/x91ZjuQRdCaiUM8cKN5hdS0OgSaIIhX6H
WDBv/wvb98D4Kmffs8e3el9NqT378QqM8u1lcdBR2qAGGikcCOWMbKHFMZL5
pEX9ICv/XGb+mW7ZE1q9zMP+bCyLGON+6TYVZjlReEZN0iuImEgN27ciVelW
navlBrk0mUcq6f/H3fCog9zjp1pNSk8T9X+1R6THqiSJB7CP1/eihI5LHCXo
OltXqh6ShtS65f5aS9zIEpQ7B+4UrjwYVPSQE9CjHzlBWGA2B/EpNn4LoC2c
eJyL8ywNnsR1FwYdugf7rq6Zkh2/KcNuPpGNeGjOkVddAhvlnHV/6R6dQRjw
gblIS69HPqZZRN+Ig1KJx2mz2lMwLhO9NJcAhPaQohyLGFEMZ6i/gKy5MSSy
zbx8CVIPNgWLn0ed4KKVta/IuEt4Y4vIPiXkCvSka4HIUNRUTozRoAMfJ31M
UTEbasCNfQHkBQzMubpr36mY1bVG3RptidpZC5I2Xz+Y+W2zvwvQc6thdK9I
c1u5Eus/2rIuc5cHQ+clzlC1zEPrLaxLvhvPIAEAb473vCv497QgfinORUDA
DuxBozGrFKbBcmk/tIo8/bagLJ9vUBiQpdZoGCFSkh+hKib237kez0svCYkV
KA5XgWqusiDl0E2muFOzhjEWhNshcibEoJ4xLVgZ1CJDxeDat3H9O8L48+St
vqUXbjI0IsB7E0KSRSb+cOfXV89KyNeRMQaMEW7UKTNdTxpKqjrFAYT6p3rB
fDGfqxfRboTj4kdQd0eWzuMsRq3HavQtm0Un61OxzJUu6G/zjacxGmLyBT5O
HG11bgJnIm5HcRtryO7UDEoUtc0nkaF5rtNwDSI4xRjI/guFj4YJWx1QxwBJ
uE2V9gbhWHoIM7YhmD7oWG2NjsP30rcagzfcv7jKaF6kcd6Aal7BpF1oJdBZ
f845JS7GwusMfTFYLOuAIrml2knyEZDZeHyQxPZy0gusNWFO19bBZ8JobZ4n
IG0eM3RsD0iyF6ULyB26OVv6+qBv8tyIqZzTSjDTARzHuoh+/+riKPvbxW/u
eoeLI2ZY4dGqDR+jb+TXZBMR5cZQkyv0f4dr8SQ6zI3NPTneiuqxCdcY1dDq
+ejIfTfiRkx/8Q4ynsyvx09M57zZ+FBZqQrOPH5x3Zr6WffV6/qHD9P7eeyQ
HzTsPMmmGzTc4zCtrM97jkJGBqVSTt5l7hpbJMkH3zhTb2v+IfQEWZNBIp9S
QZuON+At0JxCEFdLkZnGMnUf8OAY99FC4gl1KNOhIbfG99ouBvt4S7h41VOA
4O+I0YFNGNFHk2i7SapwXJDgalCLqJyvUVXkfxlhH74Suid4M54vTUHil+Sa
FM9tDPQnyEi0WmadHqS0QEmoEleJPZxBVOqiWY15+q5hDS5r4oEgmy5aTkW0
DbduFtAUb2i1IHswsioRSO6oOJmlJl42HX/+ZNdzwVWC4p2FqEhJ7oMMl7Yb
qYG9zDOP7HdEoz3trVWJm5WrgsKdaYnvG5EKzB4xpNfhQ3/ZrUAire1FACYb
DOBYeBoGqBMeq72rk+F1M/RKMqYjppy3LoCeQG2x7WMDycmJSrEyfAnd+TPY
AHrnkahhrcaZtLfVWskAPqebnXi3XzJ5gRxtisqs8cT7pN+1PH82Xh8bG7e+
r5m8zoy4u/nZIebDTrAMzZppH/Pmyo5WBnK2dF9kHRmWhADQyHtYetF7IE+d
5xSO71eNxHOBYlPYnD0JA8wpDdaByz9j99R6MzUf5oG2Sj1wusxAXD9zOcc3
lynEIGT5M6HI+k/2OLm1fiORlLGXojmqLnrYRUB8/8QDqURMRfFdFjzwv17L
AYBoE/1QGcq5RvDo3BG34AkR+79PnEBHwmh8qsH1mfeiA8RebL1lfQ2PbShV
Bm5o/gbYRQ8WVA3fRUPCyLjz6R8STrbhc5cEh0rXIorL+o/dALLNM+Xt9tI0
4otaUMqbMrJWNsHJe8tZEGL+zEPqN4VFy4zG1aNBFeVjGkA2F3mR4wjOwUt2
J9o64/tIR4NT+vy5qWcYpo1AI8y1bzl8KxzseehyJ3Wx+hy2flicUOZA39b5
MK6oIJfvs1vsrFiZc5pr8OfsqH0U81TQA/448zUdEUA0vXdq2IkgA33twE4W
XE/hjSw6vndn1YKJr929/wEmKnkyyq1OnE86Powaw1G/PUv/qI7I/iBR8epn
ChqKSQ0fmSUGWzK6a3gTn6F4Jebu0PK/yafUyNZ3M0Y2/wQ+MigrXR1Fb/TE
k9u0R1Yop6Z6lvA2JOFPXUDE2EwM9kG5QK6Pz/f8tMUr3kQvS8AVD+0zEI4X
qeLjwKdu7/KXFr9BCzkh1hofmRMpMk+wKpweEXzJ7j15ZsMEydjRbMZ0qbth
373pC8IvWnF8YrkurmC97IgO0pthx7p0FKUnzCkyUnkBQz71r/JK15bgEN6U
LL9213YlarkCFxJO4pmqXz1RZnLc9qFQqVNW4gGuxip9dy4VqVOMoJI+tpOH
OZUolxW+R97RuxPAQuxcpSbdM29t1PV23rrKvdI2ntumtJP/yFp+N7vWgGlk
vUydt89NfeH2f4byQLpROy1CA7pwhlA58djYVq0cVf4yu6SggJnin01SfRw9
ihv1EKa5o5xGjo2OfcA+s1kahBN+KQeK4S9zCiy3shWL19PqJ+JH2db6OTii
qpPEf1wAG2aiK98jrol9W8oCvm4fjJ6ebZhXrz6E7xjfQR8VN10MB/7moqEa
3Lttd5oljBuuVq9tyiYNqVzwixpMPkJqc7IdzyslWEUdIKfIlJpVuKoT1iCm
MaZQS4DRUYuWYUwz8DO1L9vEmKk+FAZjhCKIoZjuUyAPss6ONj9T9ixdExvJ
is50JE/Xwe11POEdc6pBE8vBE0TuQh/RTAXMT0pVdo91/ASOQaWui6RzMk27
cl0OkSfkyIUkzTuAxMCOcXVIH5yqQ6yIUfdXBG7vtVaCHdjcSj+Y0jPRh5UV
OCo8H53adsCZY11MMwhKkRa0tiRqF+fVZUiUhSVKTtN9whVLTg3JQjdrkp03
snyQG2F4DseEfhal3L7gJIY1JAFiuTPclA6RyQShqhaNMLTORi7suSOCf6Id
pAAVEcytfVngJv/C0zdo4owQfwznfY1hsAJtJNDHDEyXuIet3a2ARWj9Iw/I
qmm7EHbtsvZEnfUO7Hk+11jHG1EQkxyPE/OrXRoCfJcOqrZ8XJyadE/QWyIf
ZL6LMFweyAkjF3NW4hKwGmRG8Ct+EvQK8ZYoFRMhps/2oz9UWu0G906hXXU4
iBDtFHtaPVoiPGfGKbgtkbtGC9DTw9tiZwSIPTS0kNERCplN7+ia7pyIF27A
vl3LZyK072I6MEQAh4N4rudwsrlDih4I2lQutUf3/HYiVyWj5hAxt7IM7I9S
8DsnvUjXct/Ig/rkudifLb4dJvDHKs4xuuSro5UomctCTDfWNQ26un00N66q
QMq4rRwFE86IYpWX81HPw9nCaEL/K/xpzyr1XCZIp6zTf3HJv57M6IVES3RY
YQ/YrRMBT3TtMmckrV3l8cOWlZghrNXIr+9sCqgLMH3ecIxKOuT4obJEk7+p
aNP0RKmI/hU7XL0ap5SBch/U7bKO2MSYMfByehkzz3Nj8yrc/T55ngoOYaoi
A4fscyp9OVdAeYlVE4wnYfOciABCtX5x5YllIRfmivwvpbIxDr/7S0/PWnQG
02AfVQkOm58qXZxp2ruDdrMQ+t0FtyHJp2RxpP0dlD3nOUtzRsVMkjnJ+aVN
szKNswKpfkP6mmEkuqVb9z/JMJswoetdHHLGr0/vUycgJL0gGmuUQS4tX9jc
GTWDGEPewyAwRtKs090t69uBCQI419RIi7VZXqdjcxq7EUntmTZi4h06xURm
hxRaiIjW92iOqeYwsa+sBE6YyJjn0UsF+bFqkIi4RgDeKx1hB4K8GO7mf6ca
e/Xo8Mj4KpIcNFXYjfbbRw+C2pZHxF/ZEz5WO8BZ1qVAks3r8paxbfZw/QzM
VtxUFGIzv9pHUMHwnimm9hDHGy0wkuvBVwKEv7be3wgzSd9sAxn24mdp9e4z
KbVKUnww0sWZEqBRJwiW0H3KlhRA1NPHGDsXKhM9YJoBwNse58kAaO9T/oF9
UWBq0HwozzqkTzYsvUreEs9+OpzXOMkcLEZUFLDva02g/871+yTIubEY2UcA
aYaqpxMqCwM4BY+uaTCVTWURreOHIyw0z8WJ49l7OMm8lMjw0LCb7k6N5/vW
AkR90ge1FplDR5S8gIlOs0jh8tYmi3UH/mrNWblvtIMWbva2MzWDFkHGAjkr
8Mc2gJxlUlfRFUjgTEOux7AZ4EpCIArEbefEWJPUO2R8XPm6Yw45uL2u4XCx
5jTtBddjyPdMk5XidilpSbSXpVEGUyjIY2VZDO4bbWNlgXuZJkzm4GDxFVYo
jDHQYgG4jC6ok9rtieZm6HCph2VKTBUMD1QuVwMsCP7YKWfA+Y23Meu45Bnv
4YeUBbRbgzfNdiYojVxwruTX+V2xCkhOaPfMv5+AEGqI8vGIzmI6BXmgRSCF
x0Tn6XZZiq+EBpigoRg64hi7YGuh8nPpevd4TojOyw30pITQqgBduMUSRC80
LrvqAidhEKdQnydTVesIxMvtCmt0nf7jL383mRXVFsilRvZCpnWVgPisSSi9
q5UIVjJfUOj2HOJWPHsWNdaBcQVkD41gGgWL6DYCmqcVZC9VAgElXJfLUeDE
gD2boexCDQ/vM+AsyGB5Smr8X8NMqezxdku6QL5EBZiRoCpiv0DCQU3dgWi3
d4HkA1f9mqqQ4nUsxT8KOyh2yjsxwDZQX5zYvd95WEU0ryk11Fd7zVxHzed6
iY1CnqkqMG9WjdZsosKstVy2GL5Z5IQBwsigy95QA00clLpMx26gpD8cvv3G
yHG5xLd1CctymEZXUlCd6Oo1O2+8FWTQTbXawkXtqJ9WmCvgy6DBME6Xjswd
GM4XZy5IEUpU3VX0V+n82/eSDlxDrTx7ewJ6SDbv6n6hGaBBTP/J7dtz+G23
8aliRlw8cgPU9byFpLXIeLrI1eUs8cNRYGgHGlyK7q2H/wExCsLJ91f5vpjQ
VqJ5stbajWyhCfNz8u8Pt4MQ3c+PXDF5gOi0Sqohj2mSD5UeoIRSJziOtEJm
f4YWASosk90MY0Uv3XKZVDefdrI4czjL0WKKnEKwlR840tvZm2fYd2zmzT6R
Is2IvzkVuLd3rBRCFH2WWyoJUMjzjA7orHPlX1aUsE/zA0jVv1mQ6qeDAZGn
9WYDcJRDpt0SggXjp5OVtzAJh30A9ExQV65FDvQfiaVq5MbMWkkJhjsVdl7w
g/z8pavxZE+wbb6bPhDSS2592zfRCZm3c3OKzk0UcQ1fyhkEiJExiBtHZaZC
XVjEUDarpprOlEhbg/7oVNSBX5L33NmxeUL2357k8mCJ/TUgPHxtu18vy7IL
qlkmkpA+iNEzkL+4aN+g05vWhQYMxfByw6R/WvK+qcXrr17CYTIOQTciALje
4SuebULlWRTxr3J037Nosjm/SkbJQ4QB9hQQ/+g725xjeI8csJmDlm/Cx4Qh
bA0a6fV+JmGrgI7WzY3iizDuVxze4eyRlRlXbFOFN+t5PSR7/LKNcUqWmNxC
HZRRVwq9S2jfnDeJWlgqMs+v5Nxj6zNlyso03QAkMBnblqkKVCQ/a7lRHzsh
8fgqey+U1qgo/FD4UPgT5U6Z/ZWdaNac9eR9l++LXQFwFOt6tI3GgIkJ4j/o
fF0iIA949gGVzI8SDpvOOct9Io7wIYBtfHT9+foKZmqGnHCBDrb6nitm2dRx
k/7POiyOp6q4dS7TJNVqrtwi87RpiiJphgi28jTHaKEuimjQfWpalAmiCFXM
NxS2GvZHs3HWAe/HoxXD36wQtc95O2nWr5Qsy+Pps2XI8CqWDIOXygVkac/G
gskXtXzWgMa1wJ2lTYv3dnUOwDJ7POpTjOdHwdKFgaio/oRTgncmAP9tcxrJ
3Ao8kt7J/PCSAXfl2bms2tDPTiuiF/XZ3lMxUHVFr6apvYrDf1I2POKRdqET
BvBCh43sUov1gW95z8eplO7NrIOchL338hOG6SMd5Jyja9TXDIBXMjGAIKvM
pDa40qdd8LSiMJN/BmQtzIBe+2MYksN1+vu70pEAFB6UqHMrYmEUwYr/D5KV
CZK7+2Z1TZtH74BsjD5vrbzDzpO8icmFk+P9jfiE8cvBg87DZX8+sStud77M
WRRUjatE2M7wmZLP3l08LQ3e4d7vWCAwIzxlJthIdIXvak2UvI5hd8qucb2X
NELpXirep1KrjB2ThnBkskSZvpauPMknMq5YhinZI1F6Qw/NkaKqrxpeDxFi
gN8A/Hiy9xhpUXOQhODz0O/UMjo9CmGqEfwK84KGai0I+V/aFp6FmsVKg5WN
i/aILepyIzzfH4BigVny+4jZ4CInC/q/XpOPwGNFVP+C7xXgOaZNlXCMElWi
u6hk+RQNujfbkBHDvqpuvyb0+3iKToMAlObz7RlAM+lFmaeyBuPZhmyjd8Ny
HBrpT49oaAUL0e8qYcfXVo4rIMx3s5MjFA1Wf5Yzf4XWi1Ya5scRnVRKeAW+
vBkivoEYYNqZ7zFvovojV1yBW5gxAqxm+IW07OF008xwMhH4ATYill1O96+u
E+JnQJD6GVquqL4yBiACQXNlvdWhPfiD0WJs8ly+Gp8O+Fa8Y5DmUBxlbE4V
KqMOcLRGTLlurjdZV+UVac0wi62HCt/WmvTjbu31zsIoP2/eS1D6vfjeY9Gd
pIvq0QRxIGKUzqMZ1p0qrtoNoGzK4+zcgRD+ucC4Sq2d1IPpxBlWnCfAkyal
G4gXBqPZFxsX6k4kKh0kIxJvSEzAcwxxdEtHG8oIOkkkVqWWIUzBZWi/olDS
i0QjVCDBnPCJwsp4Z5su8Nto7gdgP0ZMYiroDYnvAFlLK4yIA/ml/l1YUSfz
hY/+h6yk8xRfs18GH4i4kruVcxkvgtk/TYJnNMvMCPZKd3ftNx9Z4opbVmHv
SIIqIdFu1yYz/2XovtZenKyGmh38N0J7Irrhplv9q0Su/obYl+F7lkOkgGp7
YMgy377RgTp3w02q5PeaANcdGcez6cmMuRUTYikZ3Xjg90eeleTYMr8gxQQ9
jnfFLftvlTSGuh0WuqAHcokDbLfnwATtzIBYFbHa6Q/UkkIL4c0uIkMVDwMP
gJ4EdUQbj2cP6Vlxm8d9+2fxw0c8cWe+N4FAF4EjzWb7hByP0aGFrEdpMwK6
gzO6uc/8EQpzrTzIag3Qscd7ogkRyVUDqXMnRH1piYhbtYY5S3RDMRu7Y01F
zCR2ZwUpLi3Td6XRxxG6SyPb0V7VtKyJLjNVaBswP6PRSbVA2jLguE7/fyBy
DDne7ZmOKnEYzpi0IG3JqA9owFWe2JsEmNn9iC+VrwAQq3OiDif+3djC3XYS
jSijuKn8Pbx2EtiWHV9IzwAPL+O7EVe1WhrFZG6S4v23MuhNel/IZufGlDat
RajjcgR+RwTllYc65r3X3Fzgew1RYj6mOl0bzSdHn/iMwS4eVIcnDne4zvc9
QDKR9Mahn5SnpGH6G9bIrw4JL8tZY0bljuTooP4IJbXrCTIM2/dDDFUzH8Gn
AyrUSfDQXxvPGgdt6OhpEJkTc/Szwx/f2rTBnkAaxR8as1R5iYzUH8FWECIu
qiIubf2Zcqi0ur7/48Hg/gOLRh8rgEOSm9ONn1MT4g+AO30cSf2Z+zciQX7J
lfMoO3Xvzm/X+/ObfUL0z4/QVak8eVnYwtbbRzdqh8JgCqd9YMCQEtF9mm+D
RkDTSjv65mYFH7JaYirCvSyw9KEwApS5iu9aclRnWbuVzXxmF2SgkBnHl1E3
nwgCNNq5RWjCb6DqoTYQj36W6wmEDGtUAGIKqdY9yinH1asVDo4yIraR9QaP
KnA32kAxK3nPENSY9fy02bN5ZqYg+RgBwpp2UnpFrxWVBXkT0aI3Zo5KqWBT
PI8rQfA6xraXBmT7s16O5GLRUBv1MtzJwFjORCECNLnfl63auCibyjtujb4z
xkOEqbTcFtYyxctBPchv4P6GOOi2euQPWbGmAQC7cf+xSu4r5JZDuFXGNlJw
NUGkt4crzlVpZbsf0yRUo42x0h26m03Yl0JXAxKm8XT6Xy3jf/JE/cV8tEQD
Ovoy/o8AfbeuECYaw15xzdLHKhFdy5faaoHBFayrvxHuihCwAiZh1Jze++GV
KU/MGmRFiavMLNgPUwoH9DPtN43S7HGiO5/Y6mdQ0vCU3J7JAw21qIrALFzW
8kCnErAr/UaUeXnDTEkK3l+AGzF3YCTdeuNDfY1vpzqH3jUZ/K71PHTP2Lqt
pbSpDIGMEguzbJ9HhgzySdxSF/6lovwkynjpz+UQC+FAvFEU+IPH4forxzFO
pGGhMEvWN3aPXvLZfNwJb1hsLpM2Fo+SkHStEQ0LRWPbSl6Y1sc3FyejuaSD
Ky4iZyV7+qRKfaQK4WK22uFCygk0Cwzvb2WV5aVO480xZH3Yg/fnmCx6mFtG
lJnXDmtRaNMmPelfyvcjR+ZNEqsih2h1hFUhz3IkNUW0IZmJ/WQCIJ+xF5Nc
wsqavWrQNqBi3Z6sR8/z6Fydu+La4Tdb90R4YKH/zQRgFoKm/zlIlPY2eQ+A
9rsuHML0mBgKuSEbMW44zTYUytqBimeWdeKl3j+0//ap/Ugz1TSWLRH4Mnm5
YGWTTRoK8d+kqh+uNMt6L1o4WiJFg7Zav4yjAVNmr0H/D59qZiTDnziM9pt/
a5fz41OQxnRV2A8+OBZkbAU/M5jPSs9MJ27ic/vtcLcwC44TmYt9VaI7IXs7
p91csPx5KSYja1e5o8KQ7KPpuekur+QsKT2SbabAFNEbhOMPdTfenvKRVq+G
bG09OqEJZU9IY6uidAW/o8OXiBwRrqXstHI692eGQb0pmQ02dotArNY4y3iD
c513ggijbRGSDX4Y7I+slVnb7qMyunN1YyLKSmqFtvHj3tyGDxhiOEMucVuy
Q/sMIV49Nk80q1Bj7RYAU3KtVInVDmKM88W3UFK2OKk0jLbyZyzYohgH1HvL
QElG3wkejieWOYvjcTVD2fGom1DuPgOhQj13BVUtcobDBKSXgXTATxcoFEWB
93CuR8Swh5YeJdTzFA4aqaHQAkXeXOmUDgKKekMIhBqGRm2aOn/Dd/6Hvj+a
6Qs0h1V5m/rGMVOnXCGUD65DVvFV2pRo2Cl7Y5Wq6hUMLZ0876rSLjfQeBfd
tW6FxjVXpRdL+Q/P9pki1rEgeo3NUXhix/ofv+ErENA/hFMUKuzkaHCuubh+
S5HSauLbHERv+32qRxdEkyEeZR1CKNrOh7fpjKUDKYPVYmsZWGVloni8OBxQ
wvTNu6Jgzdakz1JFYskv4zTyhu67brN/seA9yIo4QyAJzLene/S1Pkeq9dJ3
dUMrruRsWowzziE9O+IpXXH112NxmNPgll20HlrR/GK9gaOWZO6CZqOi9LSq
gA1zB1/qJ4AExqtzp+/u0sOCm3gscVE2i/Wyn/NH2aE/8GxN2P7GvaSgt2j+
2M2nQYOUcZbKM6xLBaI/Uwt2ate9hkhCMcqCkupCIqLgl7jJJWuBrRRLMCkE
o2TybzGm0TIipeKGmNgObfHAr1TwiDSaxdci8UHlOleKxS6P8U1XFcCK+kB7
jgn7+iKikvSmZu8aUk8t4P/d0k93z7BOtdvHXZScK1DORpIrzsfqqLlTCCkN
czUZfxe+6rPE48kdDp25+l8Zcm/CRxhw6HMsAXVW6QvGrSg6vpki12uaKfcL
oduq95NzoyhyGLUlBMVvAv9rhKiXyoHsPeJZ+QVSBR8qukx8JhEWHupOTAsl
0WbJbsc3m14qjB1eXyYyCEhYoc5+43Pv0bSeMdivOcZ7HguxJG3Ho8rrKkBt
AKH4LPfF/8OekG+pXshIAp4ad0Eebp+isVwao1JCT4Foh49HcvpWyrw2b1rD
eVvqy6TYpaBBlL7LXvHUB0QZwa0ciNe2yylnt/jPGB9YLvF9rYeiFquo1LQZ
cn2q2HH4rIAEmsrXWcXkbq/uYC4Uqw12PGi1SexIbQ7L9g/OckVIQjXhiHOj
HEq/rnrV0Fl+B5H5lqrxHD4a1C/FB/vvpcmMVY4l80JmfhPSrB0EpieIXL34
OLhPNbc1FrWKC+MsJRexoqEE53VYuNkfZzKlg5zbSNx34ahoW2f/g8eg3Mhe
8dPrt78qiaj/YRh3g2OthUFKS4bO1UvASnL3bH2VrogC5WLnLnTZaGwJd3ha
FZulbbTHYxAWWDtuORuxiYDiX6wQpGeOrT6jZuD52i/vWj4sNWUHJ/+WKL1W
MLm31/WNzaGM2NLNtbXngwQ18h6F68KBhvLBT8Oja8OOyGTyQVxYe7K2WUhn
T2ZmoTI2j+ToLstl+9oprocamGoaRlCfzYwPpL+JQXel0K5p81RlrA2N331R
150MspGamTQpC67PXMKuJNC8/79zWVs1S+LzLDCPw2oVIxRxhaKtsK12vl4x
OFO/YjgkaAe/z75IAr2+wcMNnDv8UhWJ7Ll47V/2wmZDofgg8oj7lWH2dOTy
TNa8z5lXwbpAmp25731ylWTNuY9n9i9eMI1MAjD/OnFElLE2Fc4V5Z8oID63
K4O+VCEmuAA4VTyagdfunpjnxxvNHCmFTV74vf/tuYxtT21sY4NEi47LeVYj
iBHP6Q+ikxt7Vt3n22Eccdli1ZJQ1Z+4IiuppoGSvLdEMFdykELN6yyxvDTW
LcKw+GC+PH0BdCBz8OwfnSvdsagutQBj2XoqBfIbA18YsQPu7uSZLxhjhp/8
pAl6C1lmnbgxrREKaEFkla1B9HLvDl1y1LNGd0W33nG/tgaG5w0FFyncdpae
dWnuAA2FSMTz8Cjp4sH9e6Xtl/mj55mYUbwH8cIDX6cDxnOLM0Du9Ag0VSlc
pSjAuf8HT2xPOhQa47W1YUeCueKoeCIYqUnlkVD9y8+7lZ65Lzo361YIYIMj
uMTnMfw/HfWlFnzelgZNDygxH0IaGH7woYbOR0Ya78/4PdxG0PeBYiq33QNe
erCUZr30fqJ/Ucl2+Psl+tpJRifjZzubl7szJeWIyg3ZqEanCFzSySgJqROJ
KE2yXH41IMF4XNfN5HRF9kXsjsZlRPht94GYppFA7K+opnJQA/RYOEMTVT1Q
nvkF0EpbZ0lQOECnKrX4KtnIiJP8QeSDBQ2zZPtypk2uH1SwZ4Ae1caXvi2g
KuQZextxIIJbH6ScdDqGGUFpcHF17zQh4obpIVJGhZWCZWOSh7nKq809PpkY
IeZZyhiTPA1723ouO20pZUqztS1qq0mNH4a50dGNNKb8aHOepeGvxu/plYqI
qpeXhUpFJ15iaiSA7SYg0u/4txNEh3QoEmjdpj+RUvC7eUfZNbL56Yb3EZY0
6dQX2eZt+msfoIsq1xYe4ApOkqCilOQeU+svQ8/5GS+D1jpf4fI7qivaxfRI
9LLytBwkOGbxbbpxBrwBu8G11aWP0+K6pLdXzTYpmMC/duxbb3L8YnSa3bOJ
lAN95OJ3GVbSrL7zsqSus616GFcBZ8f3Bn8dH5GUZZTyCXD1jBgPt2SKEDNx
32+/KEi1a752baisCdD5oCFSWPBSpBtLO5mE4hBRLnTPufCDHc3Xi8F9Q0Mj
hmTk5jgTzYMCZe3s9wSTae0sBRNj+Im4oK5YGBntt1hbPI+Tmi0ok0pmK8Z/
NyFFz5Gtai++fw+vOTk3IxGiUazjcoQYmKAblZZuT4J5KTqHy6EE8evqVjMy
buj8QflPQR0AohoI7kZUCv29OB8hy9jN871V78RoZlqxNfWZWZghcTT2U5Qj
XnqayTJHczGJqN0sB4dphracugxJYLQ+ufUWJM2WWdup6TkHQwaQCGE3gEHA
FApBet7hHBIbVxkAZPD045Z0clGhuzDyv7yS/CcH1cGkmoLqfUcfjzpIU3ZA
NztjwX1EtvvUPxXOIYPX3stivclD5oJrm43da8XkxFZBKNod0L+1IfVDVH4/
herDT+Y8EGl6B4+wUJJPxQV764QoXSo0W/tHhRPUIzd6ICgtTcQF7G3dxx6F
XRf/1vKF/Aavdh4s9KrXU4xDlNW4cX5N7Im6fLldpoFeraMljaeGeuNo4tk2
bTS5PyxZwK/8Vs/dRG2Mia7CFaiNadcbgx8mO49ONcAXUVb/YTOLOHWVXnvJ
syz0kTuCte9y4zV23ctE0elZ2v+5PuzAQ7UwYDm4+3YJSTtKY0eBFEXP1cx3
iiOX7/gv+0T9b9+tKnYHGr9yzwf8af36SHy+G0JjMnbqHyugEglPiqekn5zW
Or4Q36tyxhR3X5gy9am6OU8b8ai4YPkQ3WTD7UE7WIQPhbv8mu8Am/uUL9FK
bWJLmQTMDTiUwDVk1Zv/j0EgRGD3Cv86KNZ7IqkxU3h/yuNk6fJoUwtSNVaR
JSDy62ILU9/gWZVyEK3MOfmLyirM51vPfLit2OFuiMl3Qrzx9YC6uhJbHkdC
JmVDqa1s6rbn80v9cMYAw92RcibIvNO7XmlFPDH7Kp23IYuxaCvEsKLQseSv
7aVsN+B3Ub3fJ6FjwYqEqM1XnkIiYW/SRZlIE55JTlK/6BtnIQya2MvysCj8
DRumx6TT2SwZmfbrNFPHjv6l5nzT+wxjwz0chviGIndpNiUwAvs2CYjuF7D6
Kemn/e3AINryquR553QXesclDMQCQ96tK1XRXjTN0JSvBW268a8ePhc/h28y
Fw9NRFtNTLzNHNy8o6ynFI493rEJ8IWKL+2NopQlrM90ltMRQYhkRsGUd5nf
weGp87C+qE8X7GVQGBVjBbgANXbURGd8qyu9IHxSbI01/E0TjPjiaamkfp4M
39zmvC8+V2gs/dskYGabHOsmPcc/I+1YQ53TnD9if5181uyoyplMJHBKA+0t
XWJ57wTrClzE9mkRdkuTAF2u8tcJ2grSI1DwuGrXheMclDBdqLgnEpx8SLI1
0uuJMmp5fkTUjGoWaqzmFxZkbmmpH5+AOEN1ZKRmlHdA35xF0clYbNZu+N5+
t+m2oKy8jRkacD2TYNsD5at3o96rqx3YDwHWP3zz9zybSBjBJ9jjwBquz0YS
oykKsCuQbi/AoWogJkg6RBQ9U4nVx/aYywsJDFeS0VorDgP1UgDTHUKnwEOw
gsmQXsA3/hlWY390nN9F7OwOcyOM/oONp3eaPjstXREkZMc2aiCwvCt3BAUT
01raCoCUMwiYAk4F4DUkwwkUjnLwi8iG6GWt0m6Bdc3rSTx1E+cvkWWw8+X7
Q/XgiGb6d7wHs3CdFVIja6InVQwsKg+rNpFEmxInN8SSl5zI/FLrHoMV5Y3m
PtAXQ0LZosbC4SdwZ9Ab+1rivKQsxNtB79QMFAi0aU1K4pgjAOjMLPb9mqRO
7tvGSjgjTeRvU5ymWp7L1AXzyU8B4EHg+PcHVl30nx48TJfgStJ2TUZbJ1cp
ut3AmAN1d09RsrHttbzsLmEulxu9lJDkGdrwNnvZtAF0U8aunXbzruP4Qb6a
WuEoKBDBfMu7nfT0no3kFCNaRAf4m+buRa0rduKT6VRrewmT9rVvCSjCBArE
uTGvmHqLPs7k/GOKEUpe9skroH9c227fqHEU/heTPxvBK0MdTLXEsxdlZmUN
+zaR/sa4sVs1HFnSEO5cdjDUXyTU4+Rln9JmCUw4HS73BgUtfDymyoG7uuji
IiUdZ6azhnCUF7UQHRXdl7Daq8gt2OimPcA4XQUTQp/o56NcXfswniXa82VR
r6pppojFDth04pzmETeP5tH1UhenVnUt/4oRcnTRQxudAjaP9pJQB5soJt29
Ps5Xw/40Namadn3nYi8vnEvFZc4KECVgVZya+mHyjA4zpclt8JLXl8p8Zis4
9zatL9LBoz35VOOLSpHDfiHsnDt/NeW2DdOHIjBR27roFW+6SuDhFT7qxtLr
vzUdvy1yH1iE41BYt9sd8jvU1lUuaoEW1JO5EpHSdDTR9NZ4c5kSUrtn7r8s
xoA5JcVchPqtgib6O0osZ3sCK1NUt0BWFD9E89LHL1THq4RVc4Dnu3RpA2fj
JuEPkZoScB9SAWmfzhpauVPY/bnxSLSumS8v36mp0I7Kli9c/bik6IV8SKsn
e30ENx2rcz55B9C+ZBmOOu+RmsD1jIjXBlbtrZr8Q9LX5Wt0kgV3NWgDgXoT
38cVerfdGQo0YfwVKKA/ODwL4li+t266NC6TXkP5ZQm0Fgdmo2eAsla2G9cz
JKJtPjQtiNaRTYn0kKEDIsbU0TnRtpFcZWzs99g3LhPL9mAbXpS81Vw7lP98
TuEdGsRVRWH1hVZCtMw7znZRUfy9Op5hbl05mQZQ/JdzB6cbvEZHvMq99yh2
Kbl63nyrORlsh0niUxwVCpTn0FOi+PYTDvx8M0TVMX5NzbiBNhvl+HrrnIEW
LlvZtTfqfnAQ4xH4Ww1d8eKJ6Kh56zbgJAKbJbj7737jzooiz7eAAXivg01K
i9ayNAVwuagOPPpU3MjaUe9eDvtk1SY69pm7oMZF2SIGe1y4T9tauaVsWwWi
FcIjXBxRWNhkHbvrQI9OCiD/KCecX3xcJQNMS/JfQWfpGfMMcGhTCdezyzPX
CHSVc5XFxCzQK1mpTM7ExsshnjCptyECaWcCa1i/iTcqaDq/tdYe4EMlJclk
uUfp+tLbhz/R6jq969MMOfLBqfFIsS5F2c3Z5OoB7tnL/GuQHaZw+XEy2pt9
jnUQoLcSfsFfmwGhJB98xnpTsLaFaNAk+MWEr13pm5WzjGaFS6+JdcdeqGjz
1BPBW0QVy9J3DzxJ7x4uMiB4isSWduXG/sSetvN6EVjLtl/QK9o6+r6kvkDg
QBKBtIE/ptr0ilMRh8gnbsmqO8FgtXvYyZg5ZETcYsm6ELZFayVBaBCnY8Wg
Hvpfe2rs0eS1vcSr4AHXUSlADvzOKKoFRgU/y9y3rCdRD9Hy+sNmx3GeU2nC
ggcYZTtOyufwNpL32tdooKsbz1x7OV44NQ2QW90sMcra9jFqFImfSyFDmEJZ
DWyBJR5zqaXh9nejWn/0lWs/NzYtac9AvmQnrazAhd4vFEIA96Kv8UhczWhc
etF8FqZ6vAiZAgFV5opbVQW3hDCTunnw6eQQEebMTYmgT97Ga+tlY6yQ9sQg
iJFUYeLh9HQ/2aDQdzXXFdtzC3nAWwInDbWWPc+UM362e5Yi8ctTK8ZUDWNY
fBRlA06UEttTfP9oeFev6ffKtnRqK+xtJOeRLnnKh9r6NL0vNNJwE3YGtfKG
nhGITgyDi9YvKnOeIvK7m1xErl/nM64sfzTZ3c8BAJDBovQPvJH1PPAN2gvZ
DMdoXAdh0ySHzG4dz8RXwlZdXa5SxUXwDAUt68pHbPub0qr3jCjfa/8vZk0F
F/BL+Y8I2rMsByhgEr9pRXlc+xwdHaBeFJ4+p/rrMAqbNqVnErhnu5XPL2p8
82b8h+yjakycq7jJajj6oY3L7sC4wDtZyXp4wAXgHyACjzWVUdDhgHt19BjJ
I8FpdBfwot60SaIjb4aZ2qObe3QjEJOcYRRvY4Ha8O+KQ2l9PACySUmTxtC/
9ADZb/KLEiETh5220gy/V7Y3E9gR/ruXPzeRjQICVYdaoYBWs14nOtoSKPyl
OXlGgdlzd+oBECupKsEcHQdt5XAXZM7orR3sa4q4tKV2TZhFruuNVcn+WuOd
/Gx4uW8nVMgM8uaSCMk1YBqKQfiByuwPKzBjB0N8Xv6sCtEAjjuxmI9tcUTp
Dwk35ENYzvOV97mb+IGGoSOyBHPTs3ochJoTk6wMOfNt0DCpyflPhXNaB8u4
p7Ncx6ux5DrlsiAINRRSI7PbNbDk7UKZ127OYV6UCR8jXHIEk+o/IariLob3
9uSX9F2H0ww1D2YWmOCTBUNhTSHUJPiWQ57IWqdC28snrjV+6janh17fhru0
j01eiIM6Ip5OTAoxAXd/Ohu+mSYvKGUNv2wX0Q9EDJkyIj+dyOr8qJMVPFr5
o1kxcRpvAziOmE1e8LYhwtyDEoiLM4zsZF7aQV+F8LnpXCLtbgUqz8EGR1Rw
ekh97t3FGMifrkg05DfWtBVsG4WpYPnqWLJ5f29oPWbSybWA2c8izDKhYg4E
jE+1NmpHpBaKb9ERXyOrIg/Cc8XQwa7h9y+8Rbv0hSWET8A6xnp0gbdL2gRm
W50C5C6T8owQZdHHfagfouBzD+A8Bu8QS01DKaw2Y+47euRcPac/n6P0B+m5
yf975RF1WRvy+3ZbU/ArASXmwBF6nQHQmZguzDKZDy/B8unX/++gXwx4aCYj
MSYQNK0LzV6JHu9oZFNQifwPfrANjxgmN60zPtN66iPEWfZ7+9I99Aj7nCVh
4+3jY0e6Ia0OudxtFXD5mgDRRUOHytzuu/EuPDuu79gtEQU+FMfQ69YAAiDX
RXBcPo3TopFSrcgfOe74524EaCne/bt8bIbWTb5+lu09sx00vECjfV/Vcjj1
7NDGob63umE98LJm6i2wYw9WYU2G/IOBYBUicJIdoPvvvC9yjSEHEafbpQ7+
veNnXsIVgyuYSx2H8+sTBHGG7y4GAb25JFz9FXXM+4kMdkt02LNrcpwuosVV
DYFnwXCXZ9wTdOMYrjpo5JwIk8UDuV3Knrn6wwIbaBgiXjf381LU0yx35gsT
khvosEYsnKdM/5iocQ1j3JVhfq4cHUN0wE0qX2/UDcRre9UO/yfQuLUmAIHY
eUVqn4461lC87o0OAWrRbVL1qfMnW66cWIzacmj5Qxgj1M3BdBi2IQwMI9+m
nE5TdDucJ8XfUgIDQ59uk7yYeWvCcs7goqEzVu+7SqtYNxF77lYQW5dQ/Cca
WgXj0Y972v1Q6Bj0/qOFWjcggg3Sk6vC0rwSClPbBTTGldlQk49UGjQmxgoN
+VJOEWfVwNkpSPsZcUOVxiZ+UZ5wyD8ihOcUTUBt453Nl4rCbxnNJkMCl6Il
/x1Mv73VCS6He5YdvSSaSeE0C/8kkBtUOtSAg1ExH07lhsn0QmsmvekT3Qg0
X/jPtFANrz1F2nmEL77k4PqWnx438ReNvWpuKeMw073kOAmpo28tpuHAhRq1
zTQmdvpqHw81I1AiR48mLPer/JBmKUxJC7mZiKZc1EFRf18CTLtjLQOSVdoL
sJx44wqk/YAbPecDjRU0yP5xKpcKgOLPquRzVTnr2GCstwso0R28af/92x4M
ZgZHrh1/2w9fePocNWhhYwRHuRnGmBVWtLt2MjJZCPAtsKPPLRyOGLOXxSFX
w83nCnbu/QGDwdP2vZnH5TSOHKQK50NH1sNZDCpACIma0MuaxggOTxy+EaS9
IB5/yIirJ2x9+vkIMu30fdyjTc5BRwklIW/iAlMyPFPREXNO5+DRNNZSMGWj
eR4rCw+5QZnswqUIlPAKQdwjc59ExDXlRnT161k3lHvCfAwLKkHVeqrNZ6Wx
nXSc7PXhnq9ooXHTCW33mFmFO4IppE0chAD9EUCPy7bVt1vX6J9Bsr8c0+6r
ZumZPYCh2O5FdITLXZ0cvbdf88K/DdXwrSMp0wcz6ydDzBHrgL1JKFqzwfgH
KK0yKcdocf4JsDjyiQ+p7g27qaW739laQotl/Wf9qj7s0CNzsra+/SDZ8GoL
t+57CyCzDLUfxHCn71a130N9G3quGc/zRDqmOLBd6Dv4TRctoaBpKnPomKL7
pQ0iCuNFvUJV9S4LeybMR2/atVvOVzMyDgdBGIFCbOS3CUZxratagXC9Cavq
5dnsqkTupdUjp+CKKJNiC6kEZ1E3MdY0mN5WA2JSFxaDIV7bNrthkMHxxC0O
LDCBX+FW84jJzDkQH24DfAOa5y2JvtjWIfP0be5MSSq07HrePRyyexvLFyW1
abnQMF2K3N0kOhZpKRJrzyx6WB6TAkTic23ZDCyc6l+nWKB302w54HbX6YNi
t2k4nIdBO73FLWbMvu6SrItRYlI+oBUe/VjaMJDD3ioII88GthMJ3j4c9DfX
fZFJZWWSk2v4MaF29Cc1vkHVXMlvxO16Q9kgMnNsfMr50jo2JUoBcmoq6n+C
64xPWTyTEUAYBKuRecQy5Oy5R6HCcdVIyL8/WdotKlSiVLQDKmrorwX2GaGi
nvVDIirc/Uv+ovmGfsQtiGQiRBzvj/GiBwxT2CvlC5MJzW8Ho5iXKee7J9jD
i2vJuoNK854bzqGp8p3/zD/24OSZ1SpZw4wM7f4u4XniQRsj8CqRa6yeFlAN
aNJQNCNEFCx0woCH2SOnIPOg4bE/cewBW+i9aWx1W0iKLtyFU7V+BL5b5EI+
O0F3KB/Pg6JRotJOnHwtPdRn0cjffP5CevgIg7GHPNqwYZslyl/IDTfnukMH
0IuuFSas2T+VVyFft5g1FHl/56JAnGmAqXh5tT5QEu0bP9PYoE+lu1oCJ9iE
EuiKLutw6WnyL8fMoRiju0IsNsUDE0tZBTCvBRjQAfKeBQnIMyuiagiEEKUS
lhADn1ouAyD/OpBf/IWNwrBJ0tIM9YzWK9DmEVqZKZQNXNQiyqT9vqe9q9RB
GdiC57uZ/yWK6elmmjxUDSLXUmHWtbKdG9R/AwqG+ggaCTn0NMiTQTFF3jgI
0te1VvXG2SbKRZOSmhfeAX5t+MdGS2I+8NMeFwaJp+GzYWtNwqiVpaa36DYN
br1MU6/8BzZVWCR8EjCyqQNL37A/udSPdMP8ZBFxorZ1BbwC3/Ln+3eVapB7
ytrNc8gE12nOSPBn+/tYIzhPv3m8RvkZ9mLwMX30FpZhXxm3w39kwWeFnBs0
T4FYpLE8zhGCJnSBb5ofqDeIK1VOIqec0WqkAeh9ISAOpM30qZMJgYMSSJge
nntOGrzdbAPfQ214kRznt4ZqUA6XL5C7Pa2LAIgX8k0VPs/muN39reKFrSen
YJJ4gu1X1gTGhIvQsTc59LbishzeIhRO0EZQnHsYZE/RH3moDwRq2SfiItgt
szB6jSP6zgrGLoiHGSXUxstKIdqYqUbmfd7VGW5qtuJYRbyKO8tFkpJr70gC
hnXCbL1uGluTxNcvxXCzPpzQhHBlHzKHZPrPbBo2RhkwsTEemviZeAt72dF2
WTxgkvk3yxi2Na3F/ZNUNfQNrsm2mGIZKcBvCIyovHPc4n2MoLz6KGFYkRaX
3ww+3qWNiC/Zg+IAqtVbOqguAF6Lha1lRuN1VNfji8Fc1OgtspolaTXRirdZ
cM1ImBgIuM1sbY8egV/6iaM8x3BNYISMxD9Xeuibq4P9u+w5rPiY1Fe1dIiK
cAvlXz/Unu1UUqHjA/v8RkSZYJM+MX2GgO6ISVcfLUBSJZzkhmjAYejEueQA
M1KgU0yNaJivNfUdLfllNauQkfXl2S5NwnmENSP3+99ucsWegtBG6NkXW41m
3TeNq70vWrbSldsdl2NVix3v4IXrCGlzZybT4wglJh5Vr1u3KJwaDyHM2INh
GmfuNhXJu+c3+3Cs7Wea3RlrSYF40OE48OsmmVvTSZ8liCMNRYnnmxw/qpti
tFWwywPJBrw9bUMj+Ro45BjxcIFvHFG0DEwsS8/WUPEXyFsDpf0IlcOWbMQF
z2hB+qbXJiheD3vxYb1t45AbKp4BZjGRseVtT90jBs3TSkCCUIi00onvRjud
D5IrA8HfZ7BAbrssuCCW3avkzZAoiZzowLfspghe0mnpN7LkUG0arbkZJpG+
UXO82MwdwwHxpp13TXL1AZwtOfcseblZRVv2XnUCFjYmBS7NiS5KHRx+X0NS
UaOcOto/T9YDE/eHao7xs46HbaktigNiXlLQAlsdnbQ2Z6TYFMTRQsxNdJjB
YsgecaDS3h5dHjdANk5gKCY8cngI5Qx4jHIxpG1Ez5ohEZlRnh0xjsKVlQMg
5hQMb7idQXKfXRoe/DfzmpbJiIpOM9ZNIzynr9GxY4pQrY8lGaRDwbLfRDx2
dN8uap7ACM2aXH4x54w+1fsyZKuFAX65+ZdaKqWVj266TmdkIAjQMhL+e/x0
xL6Kl2oOXRDGQjGj2ZHsnpc+czz5QwZm/c4Diezl5JiLA1WWJYJeh6A8j2Xj
kMvTBcbcg8S+jqFXEZKYE/fA+rpmQFOk3BloH6xokp2I6shQlYz8aR0SX5mI
1bZ6iEkMKxq6+isvUPmF9k4ccqj9BoVVaXa1i4Y8xR9B9+nCWaYyDAAB6DQW
zvIIIEiwkAjEAUIVFbgxvEa5GvGpcuoFymwwPMGxcBbA3z7HkqNNHKweip+2
LqD7+RkXD4Sh3UpR34GaR4mWhOlIS5LITOplBpGa3m1X7m6ljnLuhfpvSlDB
1A4RbUtDQQQENZ2uJ6AAK/ixTfLJbvQqRPj6ybGwFwi8C1wjgFLd76DbGkOm
HtaFEzh93/7CtRNSee2FYmbiSyDWN3OhkaoJ3rRtBZuOfMvO9/z3pZNks7ko
atQ40aQ+j2upHr3/zw3laGEFuZbkNOh/43M2DHjlQcgNXMYxZBGpk+8pEp/g
StAg8Lr2xks1+NAuxBwsWIEszhcIEUzycXbOyaaPsf0vquKJo7pNxqJrqhWa
2q/BkQ8mbh5bV3+Phu1Dl+BN+wNiK1swsKhD/KU/vrnunDpya7PUjccLzHDp
et2MCDYcknCHBto2nzg465G/CK8a7ayNxtkLIUXemM8tFnzDlprrtN8HzGrj
gy1W7wKgHoBcEBBwjnWF0QxSpssSxWHQ9BACykLCjKDN8kxosrYtheL1LSIL
RTMLomAZqIKZWmytKc9QqB++MGUklTwgmO/+1DLFTCwQXvBkvQIyaQlyRCvR
aZn8ttWCs36rtehylxTPO+ctyIGgIx3oBU3m0k4cnAU0cKWELRxJTFMaD677
84gvFUhRTGctUg/Dyozd2wjx6AwdGxdlY+ahWergaOKH3ELbGyecgT5BDOGt
NV8hNFg5PLeiCaIzC2XdyU6FHk8Oq1T6ZD+Ss3uSNERaUDVFtfBeFauIUaLb
8++p7Tz2TrAb4W1SO75KP/fPSGcMVA7Sa5VUC/DJUzfJkGMEX0omchyXp+8t
cO5+G7rSB5rdA2BVN+wWCQbvE/bMLmv/OHfedD8WHBsPp8XxsfFfXMJvoV75
qGJPnUdEzUdbCtMT+PugzEIav2n0J+y0hbfLSWLUgBOPMTKOm5PVz3o/f6cP
n47EHH8MobL6z4GfEpidNy6MjdOKnEdVQ0KrqW5MN1qkdsDT9kWndrgyeFK5
9BVN4+BQppX6j8glkM67ObJQ0FVEBQsl4h4lIQNcCCbp5UENe1qDmPFv4Dy5
TJaZxEeDVotgSxvd/0nE94EKcqrWi3wsl0ysaOPUiwuVTcq4dkECRYywLUp2
TEt4MQpQVuCaAtib5m0y9vmYpL0KEGx9Uh9ytkiq7iTmha8J5lm4DYT6wXXn
uwtluza9rDX/N9vudWlt+zzgp/cELOju8bAqq+UP7HYXW66QblHsjmrood2V
Fom3Q/N4HiVhRT1hmS84BwM+aPXJpEiTd2m449MQVp3C3l7Q2M3bDMiZtk0B
KBRXpSpXmtNvo+F2bUqQ/5Q5kSIPYiAjrBQTi/8lPKM+qoGLPUu45yKmWrRM
a25apd9eCGYxe1y8FqC5HdJZHplQSCGWQfew3Oy9z8Zeifbf6rTCRwZIO5H8
Iyx+siP4yy5NJd4qq6PpB2/ye99txMtY+kofs3FQL82ol8xwpeIAFtfCb4IZ
Kx2qlIhe3vNQpOtP6vUq0TS1kv+FFuw2a5kJo6QECfVfwkRXAQjfyc0EDA+P
crS4I6TpB/KvHUnZMVi5xtLCuDbG1u8S6DTZo4lt51YOECDLQTAZOToK/Qvt
LwBqaQkslsM4v1Mzv+q1jCp9IvdjM/UIOO/ZrG0fPWhplJ71vL9MhDCSgFIZ
MEoHU6Rp0Y8oeREbGXQQdvUyxjAMZ4XOVhueIC8g6q6P6J/9pzy6DuvcoSU/
9vERlllWPTjqINQ+lGGjw5J6zKBkRaGomw+G6umeLY0sY/jI1TLpY9R+BKrN
qz1BpCaw5ZEVrOYEkkg/IdRgh/bxVxgYOBft2qLBMkYUc8DClXQE+eLx586A
xC487OEZVSq1nc/WVoaPqVW4RfaPc48HR1jZudpzfOnLi2zzzoOFvWgU1WpO
e+moOoY1orp29rPIP183NTbG0OulcNdnyPCs30jC3I0YFm+j3r6i1x68bUdg
NpNEnwy4feREnhfKY+RLQSpqy8s15BTmsFnoOB+t2MQaV18GPiGbVX4gmsqq
g2XoWvfWXqpiZ6t7rTrk5zLrtY4Bsn4G40d2Tlu6yir1QDs5IJOdLQ2lGba+
VhQ01PBMCHQUDKFCKPC9zd3ROQxIxfHoBPWk6qWckja5KVblmSRTJHxEIyRP
zj8BxCiEEZEW0fC/pR+BVaIXGLxWTv0lvYdiH1TVzusA8HMxdWUx9IYRAdBq
HF+IoZfIK4zKjKjR6aRYuesrxN1tAvhO3o78tfczU/8svyKKr3FuegzYtpjV
tU2hKaYQ8xnrMAtsw4GXp6pWJswf0T+xBfGQNxKtl/6Z0BUDXvlYRUHkB4Qf
asVRIA7NIY5bEb74Oecg77s8EFGcEWLxvj1mwZhhYG0XJnHhA3XPlkgLGAfz
mNsjOm/P2PqM0W2OjZwcYwZOuicdC2KWWlNrMDp2FO/4g4vZQQSjQVyrrjrs
u8bdB2mMfyCXUyV+WhtoVOa1AfuGK7kxF2gztAFLma2E2/QWtkRnjbi26DGJ
rGpotD9UWQcJHLm9E7fxVXBQrCiwQ5+LnuY2tRanFTgOHWuMLD9OJXMsLHP2
hVRO/rBooedUx8QDR9E5FU2lBGQPExBcfnMpxc7hYxCHcKgMvIRKpsqIeUXW
X/5sZlCxDtemdPUeB+ZoERpcDu152JitwbDUPq+4EHnSAGeoJcuGbk8G29q0
8iUPXRQFkuL/4H9Lk7HoOOaRnqGmb40UvYpjDWh5HQ1BPmu2r83SA+CDKjH7
DgjUQn0OeBdKGA1hhKN476VsPIqCo7OJcePXoi17twHq6VGWfHIqA1pHypOp
g1uMRNN31ze8WcVcrmlhATy8vboSwltEmaQqR5kL+3/byvkkCxrY0AFiqtOD
o57pr33GOHilTorGdsHjQsusTzeqQ6OI3NwCgqjw2/Y5gNkbW3fh5zj/QAFn
yR2NWymez6pjE+I0wCNfls7N63hhYB6dcic+EDfn1YTZg6D4RxC7DA3+N33Y
q177+HDM787XyY/7TycfKK3iVJbY9u7wISCKO83vnSU/aXURwt2SfH66R2HF
p1z47BRulq5Tznbg6PGNtx/qCvt2KaF06SULxm5OkDJgDXO4JqIIBZNd+LTB
eg4wCKV35mtdvmrDr5TfIecuiePIzHlD4CiQPMMhEsZ+2sBnXQb4PIVv0EF+
RWytRb3eBKxwWcJcNr7KwmIr4enST9mFk32MksZX/Q98UFlSGkhGEKay2psm
kXz8wear6hSgE9RL4jZzleAJt16d96JoM1bFlbcV7yTOmBWHTflJDQknFrBq
uEWQwv2ApWD6R8bklVHoUUIDZaz0RDppyyIdCUqK+27vWn/q91y+Ay4F5KvT
rrSIqTGkGHfxD7X+La5CNnEbkQq6RyUDvsHrru5SnS75XnKYy0/rvd20LcLq
a341sXCrJuWuUIl9aIqxx/6Xkzq1JmPN2oydNGM3o5kxjnZCrF3MaDnuE5Mw
OGUmH+uHF/uQvjeTaDoLExRytu/S/bVcAAi8MWp67ecjtvp5WBleLHWlbh1o
B52tfqELgT5Yv4z4OUwjPh1k+1aext2O4ylGyeARPmoXvO75T34kUTI/r47o
hMuscmHLmv5ShVPgApwUazte4HuDLMjnkqjoBqWtSBJMOOYova1nLMc4cTLw
dUYjgnro+Bv/aCY+0VlI/fimJy26U0RMvP/hwGPbYw4rpBW7PTUBnK8sJMJQ
WFsPAJZM2vQgDvUksrRYa7R3AVtD67gTRgWDQPrrZQT/xNfrvUJcUl0LOiLe
AajYdrX9xxD7oAuRADAEZcTjkB+5XIbxiLO0lMTfeKtNwHNzPpiHf6I4ZRZl
IefTJvTJpJLT3s4sU82ocRvzV5/mW/jN0TvB086KW3YUBx9wEj2RjPg/iCMw
uLVCzPKgiSBZmBlfR/JWjFOP+LTyPMwSZqrLo01xsJzJ01xRC+tbspFATMhq
x7oZJLVLPLbPfpkP4tVU3KgSilLCUsDorxxca7ArfzaIepTjGH69hWiWYShk
M85YORxgQYShRR6d8x0wxM4KQN7Odv8Zx+M6il/KlSUVHYtKSBbWsNuM2tyz
jZTAZJmJ1eLzwyXEOZb0TdCrY/mKO0yQXyu04tYE/JzfSOYFmNCf7G+mCD9k
1nhMOkzib1EsepIbswfh27Ha9PgDRiIV2AUUflRHwLUvvUKEmhkI85qe3onB
uk/Tx1abKiOlzJJCzX/AuhECmhRK7RXNBztIoVLdBzUfwRBgTTtB1PSLzkOn
WfQ+fwWOmbPOUCIBL0IqewLeKukA4+IkeCxcLQCVlblskgcZ8hoD+88Cqcaa
ognvAEHXndIq6swGRw/WbNeYv33vdSW7etmrYPQTSuKh+kcM4Q4/nOu76eS+
f7+7gW3pS7FHjmOHP6HpdeuWYBEHJsCphRb+XjHDiEygwvQFu+RgpFa97DcE
TMo/sur9AXXYOStIyaN2b0XIsWpm0mEQYdMvdUjoepfmovIbpc9i/r8aITSx
t0OtXcBZVYKZYf/WqG48tnVYlvbpozu/LaLgxWLln/lmQrA15avhNYS5dtoh
u71AgKh2wNiSmaXZbE7eNspwJPdSz9NB9HLjRjC3efgiCUXXn5s01RAyCyap
Jo2xKZ+C5lOICfNZcaFrdB7C+xgqUcngGBB214cfG8GGLP5vQSTOv0pEWRHl
i/2hXCGfuQoRcavMvW/IL8/9xvGzolOniyKATIfgQ0VLrIDrpSkHwLf3i/9A
Fuz8ZhqDv6QcXMfgG5QNXizDMAzb+aqKWIERcjQWfIHWCXelb3ppdg4okQ8S
g9xbAQuJFe51CR+lTj2c8NTi/HC3ej9X9J71btsY9V9dZSJQn9Gk0HszAsMb
wTI8k9+3ykKUJkthJ8ajoQTZCdZPQ+rSNxOHfWo45+VHyjZ15vvRrCB7xg0q
IXXxM8ZKMkWUU5KgrOnOV8RfBT45IUoK35QAKfV7k3n9gudKI6BeW8L3O5IB
96iucDET3mBNNjO0bb9xAdvBKntR08syK/h94+3W4nwH/tWPENSCSlEs/8Bv
/8N5HLcV9dkGDgcnrUzlc0VWjYf1NMkbmxZ8hPT/9JW5/zjC/3J3TBhDPC6/
uW1KSbsig/cP0bt0yjIEwZXRenL5IM6roCKg4RpVupSGwqRlM4T4OL+ZUp1x
kXigTZG9SmmUc07GjfWSglrYrXW3XK2OscZqcCN07rcmXIptipbBDYG53cQ8
SkQd1xl9lM8tQPz/g3CK8VSIVuPj5UdEdrEUTbJNwJsE1Tw7Sf47qfVCdagx
qg1TFwNbIu8D5J/p+XWcNh7qQ9EqvlegeXVZMN+Rg4epVFeOa7kJzpUelTSX
scMpatW9qGLqrc1MiQS7Nf/7uJXiJrgy9jL6Ks5NyKtY2RTuIdnyBD810OBL
7EuRCLZ+2atr8f6YXUbTyFQfdK4xwLPOnYPPcKhaZ/n08tlVKtnFgr//T/Go
f5ZzOg3ID9E4glapSfm30GnnDE29/ArkTQ6m2GWw+oOCX41DEexeP+uFlftU
FTm1kZ4hustHlDRaiRVl3dTyo6URqGvzvn/TotqgEIhBjvFNQUQclUedZqTy
Bh3nBB+uRdd+2YSdKMFk2j2bLpGF13XLbhcFXz4lka+jInVJVPB/fgrOd8TO
H2ZWhg5tFeVwO2Cn1vwfLLiGihhSlRmMLlEouGXV5o9rtZRcvtJzFC2BuImS
esoTYSBUuxStz58vQh7hDjiaYheNyzqbkPjDttSchcf2R5426L1EI6b0ztPD
PrfIU7DxcN07OwlzZGJHGl8pNB/Lj4L2XohwiSwmvs9qHwLEchsBu1i3VOmg
o4Y8jzjgDuFR9uvElicJVaOl35oqdAB3luaXcL8xnJMZ1CmFKp8U6DR3al2J
qAEWR2qVVDgx5ZABKwTxEWfd3A2fHFIYz+cpNf1ARqHBQj9o6qx91aR5r+T/
Vwq2UNlx984i1ew5juCOAjFomeVqOYzGCwrnnegeU5ZLSFdf7XApbF7WbjKO
CTAVNsFBo2OM5P6abFfckbuFxjZbs3gWpXKYOGub5g0dMcviChM/B42i5f3D
MXtyoqRHJZO5GHSVKOUUsaU6gSfKwZSbf8pBbBRgilVb1kLN5/AbBwPn7/Gd
kVwmE+sWpeDmGmg0CDWJeDyBqC2Mn2jPC0LO4mWTtE0YFI2LU4rM5DsirpIN
tTNeQqkVSECNCnrjTPN+5tGAKMr5ehk3rMKIxZOtFDVD0sePUbn35jEVVkvE
TxO3Agjij8v0Aegtu36ozdSTskVXlODAc56We8vmFZMMu1W0iXCUso5Crmwl
/BYY/k7/yqHTEZbS6Wf5/HWh17VLiPdzp0ndkFpVHGW/zbGk4BXLFDNe+57m
zJQ2lwFpRCW5O4m4suv4IEUYRcHgduniNDTkUvIjloeZbGWTdyWdYQI+KPTq
eYvWlzr+K2Hjpjbp4/oZ/RvnajgZ2KLqo7nWvIQn780XeeEUrsYh/iyQgOjO
miZsFYjD+Z/zgaNkchr8JzO7FfoAl+kfdNUy67A1Xj/FWXrDAFW0GyzZVhav
YBjdPF0GAjNIV43JhUIeELxWas0an5IoCs1Gcfpl5JfWQjZq0Tg9JafzvcTg
3XZkfLuIYO8Wqatk0YraU7hsTfTTiIqNg8b2jAxiqlMey/aLMIEYBFIWYNUi
YwSXSMPX/gx/GtV+y1rqZ2P6C3/+O4KArx7uHKyi5c0Ll6Ze6nQOoVfPuwdA
kFXGfhDTOKn7v1QwsYMJMFD8vWXiGHB79I7ya/0fpCECXxl9MBAt0OHPPXAU
PJ8T3jtVDMelkYbbfCYkALzFAfNaWNbtHCnTrbid7a3bYDxQlderiOhA7QbY
kUXMF4OcYk4R8icjXcTuDq05IMB0heNqVG/8dDf9EuB9bGPhACPdGayVnTQL
vDrD7bEvviM7TP69TJW+GnFQjFUzz2B1fAsCH2kh368x87zmdbKkKh40qM19
fdXXybegg6jdku4aU1L0SXoleZTMxET9zNcwdVa/BmGIM+dNCtk2ylOzdZb1
AMj7lGkqSvG33DOHwkgKDQkT4ycOr+nrvZpXfL6H4usLssiLmRARKw+bMC7f
9H8Aq/AordF/+MjkjBTNYBoMf2p2vitCUo9vC2Hr5lg0VYO/vxwvlIYcWFux
ac8WveNwgK+O2B50h1D87LeHLNFny5rg6pSEtF3K+NWRLUeI6bJOPAmJB83C
Y5apUVCH0Qmo1BNKvkQOA4nCmVxgruBKdgfJ+opJKRYNEyeOb0OloNH+rbYE
QIyVU257CNT1tlBWHYvqjboRa1dSo3XnUPKBHl2L6GMtKEtvfJxGtogsP1yw
7LxJYK7GRW2giYGHvAS88QHJ+spCtqOGhCE/ALOBzrslnYlaQe9SJhy4Us9X
O0IOVrQRGNsd2BPGPNtauZOTR/342aII7twT32MSAWc2KEOWc2ItkPUb5YFa
Gus3oDo7x+NSJakt2B8y7GRj8ebmq/NAF/EQ3a2YyT9EglepzT+c0cCZEVis
HB/kQf60ypXO3iiTiYcuCXT38N5BNFKDCw8xGH5p0DRkSK+yiw0LP3nFXGIL
FpZ93fiEmhoEjgBEI7gR7pXQDcbVcDtlQjQBAN6fkuN3mZRdK2smTTzbjlDt
c04XW/1XuidFIcF/1cqxKOWQolod/C7l7i60T52Xi/158XdlsW7QxJ4VsixT
Sth9LKxC9qu9e22qZgQv54EBUE/C3+0zl41rjjHfM4FWXFHyZBwZJMuJQ/zX
1pvdC44g0x8ZAhaf/Ey4du6cdYaAn3cdefu99J+gO7JceXFDIFjCtrk0JQp+
XjfyN6RdvUDj0iF7HFOqIOrnACEgoai1aFNG1czs7xsX59pzABA4Uwt4MtmX
6z8rr84ADTIW0NuJq71Q5ha2bdTPOhYHXPXXJTb9J1fPnL6gNC4MJ/U46Nwn
GTcQ3k0m5o+oZzO3hyXwsKlkZxbzJHXXbr/RoAUBghNSYoZKZAez2XIyZYFh
5CfOHpv+2MwWNyPyZvSIEYYr7qQfc1zboZIw72Ellq0qXVG7LDZ+YH/wTTex
EYFbtRuetBGnwtpiZgks+bK2txxNc8X3UV47dm71H2P8yzYvUTllKShqOCvc
U+f1d2DOMex/kZPA1EFFg7yH/CsFfqc9OjldY5vrgwHSLV0fTPuMLLzZapdP
UT6SOU9cBD+04JUvJCYBIqtG3w5n7AMxmUTQrUOldSeqmL+DUMs999TXFZXe
QcMvOs8Fs9tS961pNLfUpxi0w1WjAMdM2o0BIUA92fDaWaQuCsOJhGOk9WBy
1AFTTgGh+3ZywqI8KHZU8lMNcGGcy0ADZa9yFyweqEon/8ZT9Rj0ySR/SaRN
Pyxha6c7Ido2r/4sNjZZMa14bf5dNGtg6FhsG4gTri0hg7qxcuo7LtqnOLx2
qbs7ZQmuRR9l7xaSj85KxMghzRfsrpoI7lsmwMwQd+RivfRXke3QJyNtQrJw
5668T7kUzu1Zd+d0NUJ4jlw8BlEsJPHnMQ480E/alo0d7zu99HYUcSjKJz2f
BakY+jVppUwjeOluId4Ob9vcNvYAHVgsZCy30jEpORcQJ8iDow+qKR5imZHg
GV/A3jJ1yvzukZO4O9GwSp52yzB3fgcEeplocIgKaVTpeAgTYdq9rvEOdcrQ
boY5hs7x2y2xaFp+5kCInlcklG2MRVbZYpmqhBfBgmRc2c1TUnA21H412rc/
9QhBW1XRnvG3aW1r2cPvtBY63q07ZweEw6qEhI+f1FK+l99VzYqIH53WAqlX
GSn/L0QeHGKnH96fB5TZFI/oZwi7zwj30J/2hFZVlrgTeOSE33H0novxfP+f
fPRkVcJXR+KsbWBVfuVxke4TsulubeVqJR4tnNRZw3zXpoMpmpCOo3S/asbE
xrb28Hx9pfvqp60pL2uQILxP0nNa27EImvGnVvkIPavZdQwe4Wmrjq21gnds
5c3aYD8cWNslkCyqE4sYgkrLlHyZkwYk1HQrhPwH+/I+jDOSfBhSrY3nrKwE
3MzzLoSKmkx+cKT6O+NoRFK0koZ3Z+WrvKwnDjnnpkn7N2J3SDwcmVOy3Oa4
FoNMm32OExlogegTRhRWRY8bgpa99S6clogBdyNZbGnDl8NoFycMxhvryJBs
WrinzUj6ycfHxUTAUYuTPadY18SvbcWeAu5sveojmyOkbjgg/TUeGAh28eP/
J5Cvc0n2DxbVag1iFdCmnO5UHRskLzuAzjs4Ip0eoYr1drY0O8swOUDiYrbi
qp2swwUJOOs0tL8R0r19/4ObzkpClZQsE6eTiqEHi51x+PONvnSK44AOXvpw
Fw0nuPzBrqEK8kxFK7pf/IacO7lZCzG8065yxGzRxRmBQGIkOv5FJQDxpAoR
aTovWZAmg2IZbqsqGCA2GY6GwAZeXqmKp3ts8+Io0P/fA469rQlDZK3MnyS4
YCEXusbs86FaNGaRwcGGuLbPJPvOXPPsqVyo9N1OoBR+OlFKbevLj2QMHpVO
+WkghjqXKB3GLuZH0jXHiT41d2ShuPag3Cm7+tkoQOqNVaKdvPoZQyaljUd+
0+eAXDiJH1ZM3y+WykfSs4rULQtIV48Iqz1r3luZqKcyPxBTFiyOvi8YePLu
+PfTTFqC8lMkTveoq5gzLwt8K7DzEoeRuTA9Nd70WH5q0lzaybgyQh8EvM/w
MznrbaplbXv3+rvdo0b1mEGnSbhof2ni0bi5UlYbsKfdAlvAaNvdYa9FHDNJ
2Tn521ymbnwrc2SuyQGg1O3ba1gJOwrz+wVcsYKZzTtpOe4FjruJz1UKdVmH
4bjdaQhy4g7aMkfIGlr1ZKdh2M5esZ/ybUUuAG4Hm4TlaXVXTQ9DYmbHFMM/
U3GyFFcEUqEZwNVs8FaOW37VSVsMFMSs7NlIGyKlvV/BBiVimBeivOHR+zsy
2XB6QMhbhVU6YQajKokAMJh5ihq/5HXcVdoBTofdw/lGIsFlG77aP3+3x/F9
EDvzwuq8z1e64PVjW9YwR5hR67WlYXzg/77Epl/S6bQCOX+yBLqmc4P8sfSY
jqA4XW/Fn0Y9YH23L4BdVSDZEuGPboVJFImJ2oJg3Gus4SM+FDp883vX4fPB
mpilqwrbPsRgkeeDEb7egWZWD83lzaQGT6m3k0TmuHNbXuJbfmkeTixedSYz
5+GHBOOQMcgn438bQUpaRFweIKovcC0m+F3D4+VHe5cS5yJp2ri5AKn2n5pG
xahC0E/4loWHKtUxoeNeyh788aio+bG9gFx+DFJoMWlPwdewsPirNbXMgIxu
SmoeEpHQs6fi7JyqIlMz9Tc1Yu5FeyfUeFIMrtznj2AD2xFPMC+2PUqfdD9L
L0Yu5DEwMEF+lUWYUzVB/WR74Iw6PfKxw++N9PaFA4GhHqXcKCb4bTxAdlSR
pmq9SSlyGHLrURH83g6QORE0ejbe+k34jF8e92jw7Q0gpVQUe4O9XnBvbhcA
ZgxXg8oYFzsmZCWTCkaGs7Khyj4VibcHj4jh0D9JF5qLyHXVepb2omL+h424
53zt0fHrhDeURCp274bcp/y4V3jLstpk1cOTNPbj2FG72cVVxdBGQT+qinSw
t/1JWZUXH+BWxzRBWD6nVBmXYWfXTLQM00Eqs9ZPO1kzS5l03MNGd+A8B2fm
/qJttZrwW/AIEDDpDleAX0vo0h2ayzNtB9ff9+wt1EdF9VsYddtBrJ5oaK8v
VGLE7tPaPnof/tuW3BTIuGhav+Vyy6X1glXA2p1y6T/cEIDVA02UjyAu6Zye
Pvcee3zjV3PLZl8TrzsMXXZwJRwIcN4jq2GTA2tai+U18IKuGDENAQ/9bO1w
RYPI6JRThdGhP9pkWOp/V5McswV/F9PT1QsC3z0/YmnOeSz5xIliP16+1NbP
bJEeSqs/78+GKegYUJm3xeaYufCFyFftNutg+J2nBJxn8gfn2uS4yhXWEY71
6LI44fQmukij6/kHb36P3OgteuA6+tfyLJD8blrQy16+lk2RBd54atUjfq6d
BA85166eZVEW3L9SVgDzdfLC9cc0YD68/YfBHH/TEAEMfBGOQQ+H5ZCIDpLP
BTkv+vrku085jgpk7RXvjE4/lFu9woAnaJzrXPvRdjWkA2eBccBCV1PC19DC
Vq6jWYm0l4Lz9lpfYYtZg/DOGoBSDnAjIozamhVJ4oXPWtrCchCu+MC2VlJM
JaNwBjs3Gsyw9O7nmS7crFl5PjUehfGi5GRsUJ/YpOaPHQha7s/VbTVRrhA5
fbyrleuPPq5vgeVXvLlJ4ESSsp53mNkYrh6YvUcAyG0PGlhVUra3PwKjwfe1
IF5BNSGnl8KNo7AlsfNN29/Mjk36CyDFAH/k3Q0md3++iGNcZr9jgQKfzRGA
1qUzX+ZjSLGzyxxkC0O35fVfKek7hUBBDkgYTLWqd27llK43jEnheFKQ+vuc
N4LknPzQLzx51qHItMRLy7/NB5lczkxcTWnMQtZzJMRj/CXLgsPZAfpiJlbR
yCG9jKt2xiEkkg0GSe3hFbxx2Wsu+egP92ULPjpPpDf1AeunQZt/ypuc41j6
Es19HUuYFG9OnLUVFV5cu+00LNV2ArQ85WN1kAWjcmhr64+gHYrDVFx5auIF
5DYm81C1eV+32+7s1TMKX/QVSes/5aW3hgNNcqXYsESZOB7/o4NdhhgSvpK+
sVkVyJusBiKr9Ov17WSZWbXnjKY/WsK1sBgbYm9y7T3wOPWQuozPzShluNDX
R2hw5j0gSy2yijJh1hoYeTeKB8usAV2cKg45xm5Z2Ue1ixotXZU7G3A4kZ88
1KqhtzvhuI6ytenffoH0LtoFBPqtcpH/s7oK0fx9lV0RGQO/6HaE379WqDNr
VVT+auJSP3CgebW9WNImXI+WBLJkoOgfB3zNPm+GLfq1uOI9j1Q+JXdDeHNI
mp/d0nPJdVpXu0EDuzVXRKATBzHG7l4kvhLJ5UQR0qLZYVeFeoNlT0/HbHcu
YcebyezYx6DH34qt7uf9Sf2+h9rMULhvBfhpC5MiVU1yblH1wjyHHS4G0egn
fILT/+0atYIL7xXSVWHPmo+zk7MDh+FjyYmPwE4hdTxs1tsTqAAt8QVcoKtD
77s1xxNKffceIu2ST0+ZZPnbelG+nPeMPJ1QGKKY4Ex9TI/XUL1QZXwoaul3
S/0aMEdjNDdv15zoxwHmfoFFe6CPcDeGxJv+VwahMX5Pgmco3z10VL4hErWU
jQGMAGJEEaKDNSLg7PS7xG2m/rsqmIWiS6rJd0Wd+BwHcES/EUR30qyKX9GU
Sgo+YbCdEhhL5KbTp36WwtODZQ2CR01dsqPDHocIzdA0tmKFrIk7QweSZZvl
+GQeR+v9BZayCqU1uCCQ2DfnrY1T9pW8I6Tw53GFQx2+t2K66DTSb0qNEPUA
89p5UjeNPf535FIUm3G4F1TEyKky8HrSkmxUuTEJeF1XkZxroz+xP5Pk1S6t
FDT7BVhZrmKY/JZZ0ks8K75ixHFDOd2zoAg8kAImEPDRywSSQJTgYr8eXH0+
C9K8ULJXbQgK4uPtIK2lhb4jFyePS53FErVcyHeE8fMlfzF6XBp/PrqDt72n
2ufpGQSBM43P2bmCbwewJ+q6ra6f4e8TNqEi0owLsz0nAQ29rBHf2Um8OkE3
TyHnCswQLAZfiMSCBV63CXyOcXy2zVCTZ7ndqHmw10wiQZE0dPepySYdVuTg
IB+uFEhAqlOM8GCpvEo2R7KN8wCJE5KLf5++dahDXMRGFCjszEx33awk/vJa
EC0/LBl75epYZtk4mina+GBNGUjpNQw2tdnr/FfGM/WnvqdnI1veOJulUPAX
9GHDNA/3fhR6zaTTSAB5rst/SJnmE0fXZnOKHgNbgVtSwqOpylCqE7gWIEFO
ubc98QWr80J1yCwhoE+qxuBgb4wH38s3WFcTN87w/TJ5zhd9+1i61+nW//ZR
V94HTcXDiJjzKPrhzI2LXyJpZ/niFKw48JlfwEQoPLlqIoeqysrPux3mFjoi
x46EG0LnDuWRno1oqNvBbeHwL9v5PhAqkXfuOl8XTW7PfXKFfLpNFnCo1/Wd
qB5EtuWn5WfrirGX6SIcZlFoW7Kp0JOMvvYH7YGKAoqfyWikOQfiq37caxaE
okKBW+hbsYNK4TNrfFS2F2MgxM7z3TjuM9uV92yBpUL/LeKpNnx2VZyeds2e
bPXg9sOSQi4/8uhdEU0bIwB781JmVQotM2yp5U08cipmzUB/iUoUERcJ6FH2
dgKA+g5Hv9iwm64ERN1TsLVQv7uJ+I6Heg7BLoF2rR7M3ymjTqtO/BW5KQYJ
LPJUnKQNQyoXw8Ec5FDxUruYEcHR3lJft57IgcId89/nAB2bkmQQxB72/Gt7
oibVQi7dq06ro+7Ca1CjHk7pstUk0XMcDbUrRl+Pme/NIAvj0Fsdka3lzSQQ
n0qvCc61bsTh4DSAYhfNy+jVwR+QujlJ45JbULj+C4k+sAkbhn1hWOlNLNdz
vfSoBhC4MIw0WahchIW64dQSwRLn2+FhNbk+PL/Dw3Nlske4zrajksOyiqdj
awVmekf3uTlcOBRwRm+DTWEyLj1R1XbfHxliV4jw1EH89hY1eD1/mis/6R3W
7oSjNNWnRvLIk6ZLXnfZuSrZKFd0cf+k7oaor2sd7y9e34sTdxhNvo+0pog8
UR+Vs+QwoJEa/zRQQIsehtu1xNSUaJOW+w0I42QDVKLT5ychaTx1ACYt4+OZ
QUUl+9ERE3TtieOeYeF3l1uWyum8Y2qOuPYS8zzi7m4XRqHGPl1KGLxTN8wA
IdySXWxsvNsz6eEbBvwSyrRKnqq69fdEN9dM9ppVuQ+1KxUT4phiZexqZrs1
0FLt8gyZso6t0ThBaLdTwZRToj+qekG7vVwbRY0RK00RbZ6hGjYrxmtgkUrB
Pa1zqDDX26/Ph/8526r0ecWh2PF9nU1shlI05AwmiwSiFGPDa0Q9LWQqSDF0
n2jxJCZATqyqxAgAHOVahPzbQ3P8y2NFv2wHttXefmWJ+jGW7chDaPtcGx75
W5SUi/9i6J9bbDl5KM/JK+Xk+2GAcR/NRkf588wU4949wV/0FPLU+oXIFiPq
OR9Or9oekw0It/5gTVWKyzGRz+L58VztDixLTnJEcecxqU6ok/OBeL5ghUW7
ENJlZJUhJXOF+i0rCl3+U6Dsft4DquM4z4m/2FZL0Jd2jRKTyh+x2MufaRdN
YIj2rkd0vzN0jN7CH/69XRedgU7/hyUebSkYwYTZ1zHCVbqSXVuKT/rro/Xs
2t+FsogUtV2lrzNE98QjoNeieY57aWSFv+GAm2YtjT8fX41FDDFRq9NbbX8p
QmSP1K5YVPFcOZqGksTRgObNnqUNTt1csWBEHB7b1xJhepjvG8PvYlBQi7YW
NxODdBkhio+EwKKQuPnPOha5i852i/O3a9vE8vdPOKepDN9cPnhy200eNjG5
wv1iRv0F4sQgp15KlXCSYsuHXsKfRjiE/UQ0lkw9OxcFLckSx4AnsBFaeYxD
2f4QcLjmCVQoWxnC5QshQtNfKzW+v1tKwZPM5xMOsPJhG6gqosooFahSQ2IK
YZLQZObteh2FhJ2mVkOisbTe6rLZ41IKfXVpMHzvG6lBxLA5/0o9PLOKFeiY
7xO34G2Fb59qGV01QP2NUYF9FvvwhH+YHy6sDTGQExum3HDuPvcAwhHxAcMi
rayx3Llc/nJ0pD2Gzw9SSQoFne53D4hbd1NIiXH9TFY5JWNYaNBEhrOaFiqS
E8EwCxkRWIC2ULpHm8WoUxB5tR1tUSA5yuHCat8L2IM1kH+ucuDzzJkuhh59
DCXeSEPKKa83TURXNxW/tVGFSQi8GYiz7PN3W72jf8MWA7h4hZVhHvub3hoV
crpJQdd6cflmVZH7Vn/o+XJnhccvGtOofEjSZjgMrNcNk7Gq5yUxlKn6HBqo
RByL1Wn+ojIc+Y9eH1/bTFHh1GegL3i5tXXHu5ueFKWMhepTEwfiJUTk/cQG
UjmWMPIi5OFCjtkdAvmgQID0qkAiz1WZfXJioom4rBHbtrylWYnD1o/ki0h7
B8J63+M3lJELG6wwsSmMrgF5hy60RwpID8eqOWdGpCaOl4Rh9W9u+GzjqRP0
/1OkTK9FnTCAyyFOFk+odpC1OTiOiOmCAnhIoJuEU20vodsbesKOfr4c0+/7
aaQ039b968PZqOb0FFtRJI7rq7d8H5jvyi017C9R6/g7sNkZjhmeu7dFkJz1
OZVcCXPkAZGsx6zozt7SaX0GgoXkm43t23zLYcFYYwQ48nnZ0cvChZOqbusP
nyz9AinETmq3AK39G5RpSQIUiXxS3CPrhNSvTY9q5ghYwRS0uVZCQJOphdcE
0fEszNiyw8aX+ByYJ1zYQsmS7L0bG7WNlzoLTXKzgrqARaS4kWmfRHdpXEiG
kOXF0vs5u4InL/woxUkcz20vaFLuFEzpTW9IXknmrXQ5FpX4k6Uufz4yYcDv
n4B6Wb2XPsRXlIUhkcQtIjNl/hNCK9gUYkjv3KH+OTJkBjXs8K4F3mVs969t
RGaXMJuKlOwDItWaE8AelOQcuT0eyFjvwqGv3aDSYfd0kTtFn4//5ksz0NP1
18u/kLM2dB/UHd1qGqqgylv5hXlVEs39dFZrqDcFu8J35LHdIHKTRXMK8vVU
YWta9sO2/BCc860p+Qo5pKIoAhBMjLTQs3J5E8bmNmhSrlQ7ymTUtw9IvPrP
ZVaQ5CVwzGT/c+k7DlHJqL2ekIpx8XeDXgGS4iXPmAkUCX5W089ZaiO4iXDR
71Lpn+8rochkdoA3zBVFFHlOIOup18wJDcTDdU75zGDrRW3b0mTCyTjN7sOf
QvQTNOI5LWyZY4PsX60r879y9iJbLK5D1lxLEwpfrpkDFzMmQf9rwOAQ9Pcf
eaff3iBsy2FLIYZSPSFXkcciIflpGY5kwL3aImp3eHxDlAsYP4NwBcJuc34t
SPw2o1QRQTLzI8aQ2L/GZMYRG0fmZH5tLNjw6wswCoz83wQJfqf8W0PETAVf
EaBOFF/BfmY2ur8Kf2y/jDHdb+h3nsHSPUwsqeT65SJpOJ3QBDsycjxcD0a8
unPEudZmNintelwwxexyxHsgiOe724yGrlIn2nnfZsQoaHA9amLRSRoCdMxJ
/S6Pw82inQkY4P2zDyZ6HW/d4DPDWzv1syYdZZeqPVXtQpHuHvRvoXVclCmZ
KOjULUXP2xGxhW4zqXpoyOBmyMilHg9w9A2daZxVjsP+/Fo8fTriS1WI8ip6
C24pOwl7frSZCBdXnBpUbBDU3faWpw7S1DQ7o7x6QDClr8ZBE1h4wBW9OaG3
jPJTBExB5xhX5nPKTTMu/dUMPNYhx7tkXhr4pkMRC3XycopVoAIzY6PTZQ+l
ZYLEA8vXeOU7NKPjMp0KcYjBwcoGBqdYwNxmn5S/pvylMiDwrRf7+CYnAcwg
5L02K6FWiIqpo72EE81KpOaDi/lmKn53IoPsAeaZH4hfVXlNx0p9z4RLMCPj
xzsG6xnYf5Gtn4g0JvIPVsx7JJ7RRFsP7pouj73iYuvNvtthriQRsr6FAwEw
rS39XaJuc8BezfQux6uwwZQUM5A+ipViibo1VGVbQuNeVqzKtKRvylIqgAcM
4h7k9ZBdVDi9TqM9SukDWn9bKOF6U+msXCaJGhED2IxMaWVY295lJIHRjzLV
xDafgwaVttirTjgV1Chxdkj/FOX/TA3PgtgpXPZd5ZafGw2pKw0zzJcgprOe
g0WDX+WiAth/Jhx6OEZpVyPPcBp/sASQHtdr2ANIDHm06TluIUZmHL/dDw4f
wlE8RHZUx84WCfdGXQVP0Nzii14U91Sspfio5Oo1EqjaEqZSDTU+kf4IVFNS
oeWtT2/CkuUU6xIT2Gacr6QTlac82aRsZZ5b2TM5sQfOEX/a9Gh/y4Cad/HN
mzgG1PUMVVNIcgwc7KRgxah89ypIiqW6w8pqT3z+P5T+WG1vyG23eceYHoBp
stCiZbLRNBHOGwQoXtXLvka89n2yN1XiYw/4VABkWC/EnMKAF1rY+J9GlPku
yHXgTihR57tdgxBFRkbbAE/MlDb8PfFI/Teuf2pgfNTlAvAVwC6HwicHgt66
0g2bZkrONdaian8LrQnE1OUE0DX0QSqnGw3spAeYcgX0MRinoVQX2r+U29ED
1IG26NAHKy9LLC8LvuPAB4aC4Y27CaEj4icdWqK2mNDRksAfVCJhrDCSkd/M
NFQHqnj7qAwCUcBW9sIs0iKqv724BJHZU9bw+cFOmGzuZboHglEbL9RjAJQX
/6QqWD0hyQOcZYynBv4WGAfvoZYmNlCZQhs1Fx2qwiS7teojq9+RuVFcsUsH
xdAIag0VQDVVh1RMj1tGWKCh1K4H/x69WA6abl6RBZrGpKi+TMBewuMwiSd6
vU3Vsiy2XfWCwa4iys/TjIz6EPCH5fbJR/NERDFdUCKsv/btCjxLxEmLEvUi
k1pIQjjvZtbokwvY4MTBgTuzw6ZMF+4FQ9q8FCZa3jPL6GsZ2VjdGFQdaIXX
hxIwnf+iYPaTzz+Gm112e3W/hAdnNbIDk5afSWgcBEyN0a/s2N7L+PMgK/gc
nDIMwKvE2uRQ3vD822LNJejljZtPg3rd0c85QX7HNptQl6zZiuGwsXIEAFJN
0nXDPKerjCYry+Xq65lvv6P3Xxot9GkRWS9c57uCZd/Fr1ZDOnRuxXs95wM7
R7r6IjZnHHyElh1Jfa3uqRr8eHEaLbGXniIl6MpaR8Sn6rvQg+RoOmCFHXSM
qP2045lO6N13tF4I3mgy/dGseIGo3sJE87FH2pQlcXAhFJSQw7f4mPV4jlh2
yx9xeEXoDyHbAFUIEgbWQljt8YoMfj5G0j2WQRcNph8ANs3jVYEb1md4jLt6
NQbBlNbHw/5IYabCW4ggEHD7RC2cMUkcyAN0yTn87qfpWuNMARC403j6y+YB
tzpHWV51hfbEunSEPFJS0fK5mG/xQN4qhNOcr+9Eb3OyV4M3pQMqvxMP0ICU
bqZs+sB/IuS8uvfYdBXh9BsiSU6/CYm7OF93tDjrWrkPTRCgu2nXDpFcw1vH
8J59S7CXZ6S+bAlF+nE+7ODC9HGe2Fk4NQpmKVyjGUZ3lKFdyKRqbl4aSdKK
98xmMabT25PuRiK/OjwegxnITzdIXrCwVOPjYkXNMMCGL1eD9xAZtDe8qbTN
JoUYq9cen0zIlo7O6exvBsdEH2YIv4evi3nKWian7EUd7StHYQBkoXB7kOwZ
dfH2NV8NDtNucTs+CULvZfP7XgW81d6ELHWeEDckuKiK8eWP4EYNSGv5s8zH
WcTAQV5/4cYTWKVJblaCTC4Y8qQFWru/XaktJKMnZHWEI0/6oQGnBYf4b9G4
vo8UNSuhyIbZ25swjhvCVaX/pGuSxo1IoCXptbsieQbZlEilFsq0H+hqi/EZ
1XoasTB42B60P+CTQH8kCfJuWqEEOSKXVUmOCtfRRJu6EbAIllCErKCMn30e
TmJ1rCG12ury1FpSSymlKjjjmTQNwgPHROTDHvkLMInEnIxTJTrPgZ0EbHVf
HhQpJ62fPuAjvHlY94/c+Gb6YkIvwRpNMVsoh0Nhu5qR/HvUmaQUg5hoS0rj
bPWCeONGmDj6F+NY4J8Akfo3W/HQ01bWWuMpa4hbHqgSHRWy5McSt98Vgxss
9wzhGRCTKTwuvr7rY9DrpAGh6sNL3QPWP63N+EclpPKkq8upQv2tMAwct3My
A69GE++aZpgzoCinHt0MbuowReaQkddLcYs+L2ysJzAWr1sMPtXqkDusLJ0k
9hU7SuynN6GRMQYxkeJ2dT5g30R5E5QhsI9iYnm7xhpNnvAT8t9Fe71xQR1/
G8GSpmy5esyxtzWzu5ROZjbuQyiAHTAyiRmGrQl8ikLxxBOutHkPlAFM4Qty
G5dGCmSK0DoBu9aXrtpkdLVbtOKRCvZBJZ4acJzkuKIEywkP6qhxPJ4RqNQm
3DRhnTgeDVnLc6ki2sF1ZPItGU92/1phwYiQeKNaKQSgsnbaIzT6tmGQfJN5
M4Pp8jJRFzV/vEWmqZSl5+rjG1n5eMtXyWuoslxpd6otU67Crr4AKsDT1ZRs
D0vn8fOyNqLnufrEC2A76bva/COW7xCcD73gIBk2upzHm/+PMN7Vk9sBIX9z
K2Wu3+xQbKgXmkGG/7S1lPwYQrZ5sZ1zAgjRpV1seWY/Nz7L+yYIWOxDQnso
DXpb2g7wfzTuhlhd/btr17kizqhuzTcEAT/xWbpfWD4woiHFa54D/EyIFxqx
aX/Rba7TDt6V55Rg0ibVADlvLmaodLN9ybijvWAdMdeB6WDEtAfuPQajVBLV
PgQgqbTLaNjEup96ZLfAGFy95CB73DJO16lXCc+sn20juXjR8HUcvZNydhR2
Pu682rz5mpEh72/ac2WwM0AAeD0+Lq85XIYPtRro9p1CFvXxlqjDDOD4nsCw
4sHiO9mHpaOLVXBhvwtXO5ZqUSFY8x3Xh7YeErRvNwuiyKcFYssHs2ZsUudn
6Ir/1TyfuYSx0jDvoq3AP6h7W4yO1itYqwuIW4qiby5oYpTxYllmuNxaMupg
LNNmQs7BKJZiffx0IlJ0R3sWQiI2XdlfzrcytCxfSwEWPh2OvbmLnbe6ygHo
3YSMPAzlabel6badoDtbp3rHnhK/yRJl9GsgZZnBoMWGYF9n9740N+xpxwgI
0mGfE2btFNIw8h+FOcx5BqGXLJ2STc3rJZn+2VwK0h/zDHStr+LYjkG1qLFT
fbLY/PwUio8MFsHlHjhOzslBOKxGH7rce+c6lzCM+yeWfFqgVQEwDELCACk+
RusZZjxs1k/00bkORzXBzXEHTQJhLD2pJMsTNgWytj6ecuJQZD5xkXZGQp8F
WW6teiPk4KShahpLrrC+pbKtQDtikmAyuIx1QUFmcVVx5GTqZ2lKpoRc9a6Y
7nY+TvsNnclED5PJz/7Agtp5T/nAAjE/q1INzsAobSTdY3nDwDuQNHTmJofU
eqeYir79GNJaLVCupAJ0M8e9T3CzR5zFUj5adtpEGKy9DtJjXX0ykBSu1Khr
vER0xDgCV/A7Jk83VxKPsPMeZp8hTmuJBMdGdQsyyYNkpZb6CjuxbgCmXUjX
eukQo2zziN0gluIRx98tCqYAj+JgYX+ep4nvpa1++iUCVnAiuFtZvU3KkRsx
wIyMGguBbC9tW76jaqNnK+6hJ2diWnrpnUqfsUCl4xRNs8Of+3xVrcmUO4X7
ximjZgfFP+Il2DhW6v9qNf+vEQlZ1wGYISfqMleSaD2dhEXBqAU88PwzGT60
9no7Lx98pkZnM6Xi1VkTMIuyNH/j52494ZhW+NUHkw7WnbA+Yd2EDqQjFGoc
7RdLJ0vgcemqvUNH7lUmjSpwJCUEFN1uI04gYDExhF8IatG7wUOQbe+VoTXQ
zUmHzm0dmh+rdPkfuQut0piu61f4pRQFjj2qG9hk0sNBHbJ21Fla0IienkHa
LY6XQtyDjjQCJi7SYMsBdV95RxdyPlUQFm3Go2w5o6C9pPCJ6FG3xHP0hU3y
s07JZ/m5AImVyNKyCWpLnkdsLDQB4TqumfSCx0Pq9T9X2tklUm0/Se4JQmPv
z7J6bVsjIskvq4QiMzhecrMLxwCshMONREtNQ8m8w2/2My4QtO/t9ztdu1Vb
J1LF9LMqBSxol6+4Fi3syTliO7OmO0z3jfbN6rRohe74spwb6PkC3O7vKeKZ
cLHdY6Ht44zBsrNX1mXEBnv8bJEQtExS4gPr7S4U/WEaZE5R9FZn17nVRa68
L/E6TkQRjd3p9l3FkVjdMhynUhG1cS7aGs6GQndzkktCOsucug5yp7IccXlW
1yI5IVpcv+Dhx/JsxO4WfpF9yiJNc+IYjumPt8lK11Tie5QXcOwze44dtfk9
dEznxAZadzSjp4MtxfJEltYyuLDUbkXsz3Nn0cBcuquPpYbzjjjOcSbegXbg
pwgu17RHNu03OH8mDeaUVmLvXrmtqw+4IreP1IemfUUiE5oue9XiST0y0pVj
YTID6I5cLtjm8NsjXGY3eEH6KceLAs+896UJMm6eYHMdjUmheApvfvU6WEMc
Kh5VtNecUl8uN5BOQHfgVF157R9FjvDP0dl/K5xGYrKcW0JDMWYa6aAA51Fo
8CIqreKCNXsg165Ni9hUjV8RRidd9Y1sx1HSFW1yS6/vOGhWXFw7ADDixTIO
8x4YpYO8dLjeYAZDbz0EzswwjYjXXq5RznKNpT1LVuthXtoFIMua7NybNMfG
1P6yCXA/6gBpwsSiiuumf3SypCyGxlz6SbZqVMTouJhH+lNqE9NUjcKohVw0
WJ0Y6T6/AK4+lSrobocLRwOPUZO7r1hoOY8rZVDiGYLDceCUD8qSS2K7slco
rcpn/3iyszb4wVqjvVNiYOasugfffZMKBTMg/UxTXrZg18+TIMq7Ayb2sRYD
o1D8CBGCMcIoaVJWLj+9ep4sxM54kag8Xsv5B+I/W5Kdq6b6stJMUKUmnVlv
zIt5beOTTfruNjR4eWa9f/KTJsFZsHK4nfeTLki29wMk6iP5aOy/4NAYkTZL
/YSAZzQYctYORAHnXSIc+SQvTamX+Se5QA0SovVxV3JkPk006FCMzUQXxuUr
EaEu/Xua+k9C+Cwd8MELAta2VqYQQWqdKdwBqq3ITRBQ7IcXseBZnwQX+JTQ
PCW7KaxYptCO9wqfKZXEzBrRAAnadowcmY+rzItP9crJNtnAwYGggKYptJxa
EOLh7qmZr9wF6tBjwiuwMIcd+7DZ9CTgGcdeYuFyjUxwGUQgmRR1SLVMYDjR
+r2PK949Fp0HkpHSTq7bqgZ9aCPMj7jt4YPd3/N0lZO/Rwy2xmc3rHMpJNcS
emwNibwDVntX2+lhKDt+X0qxHqU+WjgeSta+MrGkr+/JJUY/FUQTdOUfgfta
1Hu5wHO8bavAts0DEKMK9FP9ZLwZJwuwSCAMaxlDn8EqU5jSULGCZMnDbmGn
U5dYju/IJJOlx/JEDC4JzXMO5h0KT7ZJ5SR67Dzzf22Sh2Eva+azqzzgDjyy
LhXVrE7ZTnu0ZQxTQ2xMl4WN4ks7n78a7dK+t1tR2imXX4me29dp6o2EdAdw
2sHbe6camVvFSPvXuExaed8ZrdMLRSxmpPo0igHItiivBZrU4sLVdtIY0NIJ
UoOsPWfQipXcZmXv3YWb3KAcGHbvW6BHMxhHgLczu3YoS8gF4Qf69/7vMRqO
fsHqIH6cEDZM+go/FJlhLggy6M9LAVFmVCRP2RyaibptwGmHx/v7WHsoHc0/
ugDuSC2dPF2QvWsjfoNlCMWfgjiV8W4kr+b2um3EniB/dgdWdgn6Uk5lMHyK
Q3WMkqo9Ui06Dq9dQJ3KxAEYiImrt0rwPbkCoZORUGpWL7Urt9f13TkLA0nd
XCqmMVtknfevPjnxQAz1NGHVcjxfJdV027kNoMaILVW64PUfpRqLZ6XZATlc
/Y30YEI/XrvuxNU/Up69emKxtBnnkURXvhxRD9ySI2l9j6Q50gXbc6uH/DQ3
pFgdHrNEIAiOPKRNFAwqtRGAM6OlCE3BHoUEGnsUwdZVFqsEyBdSroWfKxLN
UcK8TAFWSQJnpkkwN9DSVx7g1BdyM5TBQ/UlWuXQvlglYY41PsjsqCGowXLW
pgXIrNrfMUVlFIKSmCOmC5NCJmBy8nmRNNNNOhC9OXIAtVY+OFhxg+66uM+/
JVS4IAfP2B2vFCm8sbigjtyStaC7slB2bvO9hD+nCS2ihyq6kpPUHxcaucHi
YtJp+Q4GApNv8OCSZ77pXGMRZc6hDS+H4E8zOp0zrRXRvHel15evRHD1bs1D
5Drpn8Wm//ITjmdxi9o13QoxkwhoJp5dP+GNpp6AGqtopYd37xNqJfCoZtR7
X6g7p8yXrx6wbfp9/1DLK7VIMxMH35svWBURgKyyDQsraStlKUskU9ai96BU
7C6tQ2/9HmWxhLxzmYDXp5Rm668t8Dq6vShxu558vE2XPN9vE1CGemK+aOlm
DIKueygw13mwIPapBpVeMcOpDp2uS3qONZFMNGTxUoSj61aeXNEUEm+lXWaD
WStr0BESqWIjPoE7T93ibwyFeVy8HkoNIpq6o56X3MaQCbW8UIDPc/ITqGO6
v+vpVqQHOv800mWh3RHGpZHk4JPJ7TwAEdynOlXISmPjNWbcuedcFJFr0EjT
Qb0Tw3bJ3rpNSgjrHzMbnRJoari/O3/eMEqubxee98aIEAArYWfoL0H3r62l
2y2vdckpOZC2cqX3xi/H3Yw5jbAWnSdeFWeNMRr7wBSSQh60FtfFb5CU3rkf
FW2a4B8I6W1dwy5pMMIThvMO30SKXomH3LRGreQWkKEf58FDNygHNXY6/Zjd
7sWuNaXHRTnZ9fxyDh0ShMA3pDASiS7UuGySjGkOf6tIsr2rcsEw5KUQ3hXx
U4j3qln89voi1BBEJGUrrW5Wp1iTx9PaLFM5645qBwvz5OE71xVR3A7r5OgL
6d5/jjnRBFE3N2iD9WTXzJ4FNQWTo3L5zPM9BUMWk+AF15ZNW0t6wH7EBsGl
nvU5Xz9HtD3F60sG6I87uQbKrGW/T+qKjyeW87IUFXchd4pd4oJCMThChEus
2R2Ew2c6KrnuqkB1qdPD/jI9nhrdVNZx60Mw+I2p89Au9v0gyqlQUYZWqShV
BClZXoRds8TMQr4znVFbPa44gr8M5qIz1wzBWqT0VOjnjAQADT4vaAe1BsOb
H1G+Bucwz+L+p2iN/+M97+0Ry6MNcAsKashw9XixX721F+FErOnm+30mcTSg
FlpaXQBGAcB/hhv1E+/6UVQxFrbHWWp40230SVqoWTmQeBgkCImNFmT/lAZw
sJw1TNbPSC5EIdC4kUAMt43oE06Pph/HbLpjaF71X5st5ThOwe8u9DFT9lit
Bj8pj1JC7Ed8bOC1NEsVPvq67jcoZMDdLsMfojh/Qi6/b6sKbrd/tT9x7ueh
w24vWSHBR8eQ+dNJpCujl+yraaQOpxe9vai3tPX20Rv471GIA737pcCsyCDW
7jY5eKhA8Rxuz2BIBuXPxC0BqEw/qnN5pUAbnkdpLgMZzxBMRVfXRMWmq9sA
38ITlJD5+FpRa77WSBlUmKJ1y4VxMsBMNeidsxstfGz5GnOmzGxWLVPkxsc6
IpZZR4FI4bjusJGRj6jjjBq3JB8vOevRvlwd84S0AgUTnwbe9tpw8xDIkRpE
2UijeZdHVUzGFp3IjpwatTdlmwru3Akmww0KdF+bYhvTEeVMpz9TFo0phWBD
UNKE6nPdq1i49xu5SBdvwlueJpZxujYaO39v86nF8hGrh3iNP2YXCisWhoaa
xWer/M3s1jODWkIhFMmZjT1NFVAI/f3BHdfv+B8Wgmy7kCN/1fbK8D5ZoP/Y
/4QlTJ7SyVOQzM5J/VdoczUMQCxYd4si0362Zc8UM5cS9w28oYzPN00nS/Rb
Wbohzkn8ar6f2sNwW9KA1WF+EDZeGn0ETCT1vrTmo1fqc6/BPzoKjdo8s8Gc
xMhvG5xc1h8Uepe7S3yWR1enPOuniDkBRivlH8zON4VhDUb3p89VxPgR4ETo
XCD/x32JpqGO1cISbZr8JQWl8L9Ez3Kpc1OymlJri+5nYo2iCGz+uIX2z3IS
gOY9D72htNoJrTQnZEipZ2DDFnocbKDXJbtbixpqNCC3LCeeJZiH1kP3lbkp
IKHWy/FbPtrYsyKO92qRZG4NCj+9K7FD1AtQG/xMXCaw5Rtyt1RiRVXKn5PG
wzgoznQ55wFlZolcj/3yi/N+439sJjwxq8RVcmq5XDp2rAbqlZhQ9HQbg7O0
i++pp4ulKI0DSfBWP1TVhOJ0ntaLCsTNawYyNqFULhgsAZCAqSJ0qUEP0HDp
L4/5HsC+1YKBq41UJu1vWJqqDsyjZh6XhXaOO5SCsRRWIrGMGuz/wQcq3hQx
DywfW7Fid+5Qo/YhJ6uSMya9Pv1CsUQFA/ii+mfITfH/bCvh1LQTo67NYAP8
Be4lPr2ZKA+vgwspACXhZfQv5zH9DZTjAf+YxxFMWDS6Fh7Gv64tOAjt/XSk
juxI3hmrcsZs5k0a8lX9SjPATIukZC+0DXoGjBQ7vGezPXhoWShY7QXEgduj
6UHkTR3n+9XzHlGRhruE2RckR6P11GZn/u5F2H0cmFZymS4AVVEGdrUGmRbt
1Hu+fjpylOmBvBzFNMhRRZ2dgu+K5tNW8BNN06W5hozlqzOZtmzhV0lXSA2a
nsrUf1e9dhOskm/eypxpRX+10EvpDphYVNtquJoNbaCdqeIZbWuV++3x48Qx
lvU2WLpg+1tSMBTqvP96h3XNcXlo+1DPJbIax7LJ5puzGq1kPqKjfV2NvwAk
Rvk2DxT04eF4s2JkKLDB8wjMYfW36YBT/5fDcoyPCwMfHPZDJay7R+7FkFBC
LtaBVClrXjRFoOJ8krQx88DMgHS1pKeFseYm3H9sdAZMUJTamJsFdQViQfLd
K3xMF1AwDSmTEaCuoSMGc3QS2SH8CRbQrkDUnUAa9tzpDOKRI3XPq0e//nOk
BV7nC6PPOUBvef9yGnLUCGC+jUdkMKmsLS3MnF3SP/J6gxCyfbVluTW9wGIt
7fRHGwv+Dqh13ySKsVRfzmVgM2ZqplWHQ5OjPsDPuDJCW2DFeET+CRNZAINX
CMEKn3E6AjccgzU+8ZtwM45OBT2cns15MYa7jr09SalXY4gzjfzvfSzTyy4v
trra7k1tiMxokW3A3lpxieV2OejjcpPkNGAuWTL64h8JX/FFhm7fBoZSXzij
40frWaFdhIT0zsOICjT2aHEio/0sIIFLf8k0/xE6xR4LRfkfB+NKRGxzJYKG
iRPfHKABb3qS1VrBJQQRsd9/XHxGhf6UfmDbcp0rFBK5BWk4n4w36MQGVu+0
LYT71+8vnzBX3sViKqy3ThxVLC7O798xJkrhUrEMj91jzgRbwy6QEtXveP6V
ZZP8FpGUdhD+OrQwN682b0wflAvPbFAoGhY8d8IFR5FLmXTPzko3rvKB+Fyf
1ts/64nfWvQB2LqEd/tUnUgVSBaZdM2KBYcgMuaMt5RaZwIa5AatZG1NUDzk
IpHzmo47feEPz24q1Wqj2IPcKzKy2rEp1VM0X0D4Kbptif7wNBKogo3n8ue9
08EQMxNWbvLPcqUCSmy0oVjbAE5WiP4wDV4q2a7j4SgIraivBUGsnakIcTQ7
P+Nn4v03h8DzvbvhLXDOE1bNh7HbDTw5ZfutaiLyrqbe/uvfPIcYQ6qumuPM
SosMNsPr8IO3Z4I2i0NvHW8l1Mj4suwvO6DlbH778cdZC2v6uqyKbcE3ybXM
7HLcUrTUMKViwcQZ3HICA5PXE1KjJCeNWtKoql9bPicjXSgNawXIukvhHqrt
0ZvARmy3+YAIzXuApDjg6+mhep9tz859bePrpsAgEE58cbQq1bdxNk6ev+Oz
HWFn3Iz4aVymgnKD6imbvB18oHL1qLrVmiPFVfF7ColG56WFIHNdp/MmWFnC
XsFyH6eMT66t6tTNNSlYEdhwkYau4vNl6cQCc/FIyDg5LVJI6OJthLxMfcaZ
0zWGTIhrIoI+ylxET9F4LDgnlGl7e5bPTtnkD3YRnrG1PYSZiWIoabz7ADhp
/snynhEJ7KE+W4Xh3dpqVl6EargbFtIRWzGe+i/7gSyeXCicCkM1sqZGcpZy
4lkfZFVKAQQIdlvAMLOJ5CyAilKunE14mZOxtUo8EyFiTLdmNsHbWVrr1dVD
Jm9Tjn1vMPClRa7ixmDJX747lEkqYEuE1GIY5UWST86Y5ifj+T/aIPHKr4Ci
NAeIKHKUjgQFhjvC62cU0Xgmb3oqXJcXtyYIdUp7ja5q5eyhkIpLdI3UePFh
bdUz85WMAgm6rjtMGZKkhbcx0m44GzIpBJ8bcbzchNQhzwfCVIqV6V1BqAZ/
TwJ37nhwij+LF5YqEU3ezM6G/P2dPsU43Qks/8Yq0r0HgwawwqSC8+1er9+0
aBEIjcBSDitWFWZVzKN/Fod9mNebhfZ6yfOPSWKRfX+36NCqy7uaeybVxSPU
In9DnI+aZOWwXQB1XhVcfuBR3LYW4BQxERQK2e0Q1+E0CI/rgc79YYNp7iAG
I6Pm3KX+ek4nqNEys6PLtcsKZF+6+dLRYsMCaCOXQsu7VIyxrsITc6njaPhp
FI0Qvykcl9bcybsWY8AKrRMwkSwqzQu73o0SIxIF5TLc7gaV/eNbbH4lsHEu
s2aL3iDHV8p2fg8wXjzZu0ICJJC6RydHuWzoXyb8q9YDSegjaQSvLSyj5+g7
1IPTr6FdETfGv0DAHDXcEuCvU4c+S5S4C23qrAkBPWUSoNwMHyFwGehtxw2x
+GiFSh5a+3FZKP5N6DfImLVTDxLd8MN4EPokbSAhPqBBBJ4wad5MupVLht7H
lHcGsDNX5wSx/Z+5d2LphCrmOeGRqaKhoS2K/Yj/y7+GznUVQVxOJMEIwUsy
nQb4ct2h4ITUbgiObyrv/1ce7UgIvj5vpiseRebtRoUHrWx6yE+UsOx7gVRz
nbQpPeuh8NDf3AICUOZfEs26Mu+ZG4Hoj2w7tfROdEbp7JCxuIzqwlxKBxJn
fq0po02K0S1qXoSrf4xQxK0oaP1jP7hB8zp78F0D4G5Jlb/g2q/PeUplgSPU
8DsSJrrLwC4+s+njliD44R5yYUv09FDq7q3dEEZGjyDklsQbDxhfuj3tAP6c
s7pMvzpj5UYeVfkmqM7ajl8oTlYZMLK8BBcZIICrMjs6xksdCx7c0Xyyywrs
vPo/4A67uEP5au/14Ee5IY2191Xyne+FpLGxo1sdT/BAlV5PyPWqLvALGQq5
yol7QgV54tIIci+7uHezB3E4hrGtV/3cG84BT/XqIO3rcnHlDKoNOsv63pw+
5vm9RaNwopzf/rMBujUiiFNprRbkKG/U2LJp6FXpxuVlKpKqbkRtanqERyKU
yxc0eG9UoMpPchzg72PGJRVCAU79fj8WolEFumoRjZNKJeyn5XmQ5PIQOyav
CwaNOtnm98KehYdlKWKjJGt0dkpvSNI/cbEp2NKqgq+7eMzlM+xxabq6b415
m8Ajre82XBQQtQhrtG/3u2HG/Hc4aDXlwS+Crmb6Bqw9pOd8wnJfHYEbr06b
G0fHyPahwQ19jAbWdVGZMZNyn5mTTaleuzE7Y0mmZRoYq7nEOzW307SCwRge
tUXY+RmHyMqfMTtnlkKW7eLwHJTZFQ2Pvcr2cZX4QJNQRb+AhNIgIzowTw9v
CY0UDNV8rUV6dJqveknOUWJ/Eg1Gd/q9ozX5UVPufXZ94FjumbUGDN6XBVBC
UTOe9Xuc9gmYk8ymSYPmMKSfNSdzLWFokwoZGZwG/ayKQB36Q15TMgnITaB5
CVOAmVf/ujbcszzGqLQVAHhH2/15tNvAv5XsFzoTPUwv3KkATmv+Sc1vQRQC
KkHUXEhQxhbDVCA1BIbiN1MF7xXzlmPLrdepCq1lZ9C2qGwSomdCkbZs2rxk
WgEYZi84hX+QCTIbAJYwhkrUaqrueLcr+v824FnlloSDHUjHE+poHoFgKyIH
twOLYhc1U0D1hSGlbLEO6V4gn1oXNnKzxKwmVziGZrVKwopwNzTA5YzJDXT6
7vXYTmjs0JaBIsfNCRjEyjuvGWGGH8+1jb3hS9N7j9WSCe8U+s74T8PVXZAH
M2a4lDOgzZmt+d0djcJ3iwTQVh1NHIl6+Mab0tKyJ8g69pLZ8OzV796cUXoy
/807+BQ7aWy3cuhqL5sebLmFvFRVa8tzUqDBpofP90xC5VElEap8jbgRtUcx
qKUohhwwFf56K0BvGsadXjtDA8tc6y+b0/QugtVxTaLTAHM6vTEzohpN4rIf
xECSyWxxcAaGshtHYOG1ieqh97hiOGTCptMGROx1tBODCfdZg0RvoXByasAe
XbVNypG7G1xQawO7h26Y0UtRywhASmIecSz8XFSkMANyKMEDP7QkYg6ogv/G
qjSIo8wqVIhwGohq6VR3mHSv1TU8LCMk6IEKw7PuQpo13fH75VThBv7yyZG6
0wzLqctvoqeJ6JH+jQVlQaU1oGYw4oBXV7QcC2yQYMHQYo6ExPn/OBswQ+zQ
wGE0Re+y7vOAOBmEVJW41g9rsivoVxeR9eNahdybo/PgylO0uZRzoiipDxvH
ZxJ6PnLhfWAQ6OBv8XFmSLpMSv5qsWVu2OfhPr+JAY07YjCwA39Pl2IY4ojZ
2MZNBele2E55tYeE4kEM6uRvms4AoSvub2NBhaq0CNhMVdktNoe40qXhQNae
rCz5npPrG3ye7draYysIPlRyI7mgJ84d7N0V9HrgSlQ/6qYcGSOplTS3Gkrv
SlE9oGK0LA2KFkYNr83q0edSJiOd7shEiFdKk9bn9/A0gIrbdJi8o8e5og5h
+LuTL3e+7+ThRkBGXxtNMutcOnS/ftZmeDpfnVyRc617euAzErh63IZWShGf
Lto2aUobSkkYu4mFcEm27iJZTIhmGCm9VGBkc1JdnXyXDzujqpQewQQAg2mr
XU62BHYV8ZvCYCz9he2rrg3wqza75RBKz70Y71zJfA+diC8zneZjowe0MUoT
7hHgNLzLjKluzuX9C9ZdgJqA21Hd2n6wMqalF1pUDQWKnel9PZ6c65TV22WF
4SqbJlVhsIG+UTGQ/m9e7P92JCq8uZYGpE5nJRAMmBVVthdCJaS1+8l0Y50B
dhRJZD7rJnOqbDFmXpU2twmt6gH8FSnpUg0mibhIfGZ6STz6YyzczleI8CbB
r2gFlOLyNXMBNMj+FuJLLLfdvNnMhqBTiPd1te/6X2YpVpHEC/zjbUXpqI7a
daggR62PBdudmibBdOAHkiXgS/E249Lv0ETdhRlUOYgHGxRbFLtZM0bicAyS
tY3XlSaWCbsd46Kuy7//1ZFwZBTEiMF5V/NM3ORpEx/mQMVuwdjrRtnibXuk
UyIQMB1NeSDMXSWc93/nVFBBhp4p7NrQ5z03NxOR7VJ+ZSCZttjJEHQiD6zT
P8IJRb1jjJGC0zlR/So9VnJ7eebWJVoWavX7DJnyKJBTasyJqdQppQNAeZ+L
dBvLhKdJrzjMb+bGY8SfF/flVs6B19I8DjvxJxsnI5c5hjDxuhF9HZerqev1
L0AWZGEPWCBhTT80XanNDz5WgOlFxa7V+NPndwFPC9DTxc1wu9Bp5dsPnF+t
71mAMUiAHpKOVbRWxLB7Bnp2WvA/IY/24zZH13BzI0ytIeGwDaGM6U7dU1WN
3S5jqVsbkD5wJMaF94L2YHtSanX3s038BDbZwuzl9AccdnfKzAjB2hVFg4bv
DTGAfLU0riAwnO5/sxHeQHHj0goUI8KgV5j2gtvDBiS0oK0P+Gtu+HgyYrmh
M/Db5aAKv6dwybCO727319RKiL7W2WjIGhg1Ert6aqGML7SyEKUNQrzcAkKS
INBaElXkGv5+eLcVpjk/5cCcFVjHrrppGk1TGufuW01D5nUDabMlJywTZLpn
Z8wbBlWUqTCsFqd7R8eKXxqbwKOfu4b6VqDMKV1se8ZHWGAu0FJ2ghymH7UB
srdA6mKa4WiixJAb4FlO9xpkfVITc54H7R62AqyEuXiVdR6d12PqG+6KQKOk
MfF2Qceid57+C/AAUxMF1+F5vE4I7bkjEUnboG8n1mqQNbZ5iOniNiqA7vJD
ilTCbnlwndkHv2JSDaKuYgE7euYVVQUdrJNmTcUvxd1j64iswarnXjVyky/z
guwbL6EdpKzNmlpAB9kS+Y3HVTGSWg/yp2IC7qYwiudQnrwtk0B6VYenmFrR
Q/7noo53FYsR+rgiB7M2JkKyhCr1s8bnyc3MOn42FLQNWoOnBYb7laOg5A9D
AVE56uL5EJtdzpaYT7YJsclXe5/uh5Ery+uL6nDr2gvJkshyWDJeNq9K6kIV
PNKsFl88XisGC438VlPrI0LWasYHwIMtMaI49ndwkwFSQ+ZdN6GBqLFWByP3
pubxAMt9YAOaxl169joDfWcEy+qjgAVvf4UXXobHEcfrQPTlJ83VpGVOBmpD
yKSPgL/YEOv+lOnVGiLHdCPib3ULBL8LSEG6yple4egeAEeJqYMzsVr30vmy
PKY+vcYgjt/QbrApWblPen0QARWhO/lGJLaPCEoOVLYL7TwTx4UTrJ0NUMyJ
U5amjPq7R+qH8VsDV3jHt2ynJ2YyawRDSimyP/JBE1sgMAOHfF/mFgrxp3Av
dDhX5ZjNYvGCAVX8okJJs58NcWOSCDIPSvWlKXDoFQgoUja1KFezdpYihDRS
CX+Ez+MCeUOSuj8EYCszCdVsmJI9G/NSYbAYR1PYsKZuzxY3+2wNeU+WSmV4
bBX2OntnZVn+0wSpQYnmM4gpuFY4oQqNvTG4hDFlIrRy/SEL4DHTvtL8braj
JWFi7uUizVUNwcO3yiq5nIHNHelSJuIeUhuSIz7ty6KUYRSiv+r+fwzNCV3B
Fkjy1Ehb6j/QJJqQ/a8oqF+Qbpv1qFc55M3fHMDR8ORBxYMITDBYhtJi8DHA
TVuLLUCTf6clhmqRTGrQGav4v550yV2czgYrNmMI17jIE1met2ryMItjOTvf
O8xU3xt0dh23p2Ie3lA90nIh1HBU2BsNeLHpVmDZH6mrM2T+WXzAKr7hiy1J
BB1+CsJXa0yqgGSLQ6g67X5WwYPHKj+YAvg0g7+PRQF+mjUkSAZOUX/f8VP7
b5KjsbB5T5uQBKipxLbKXH5m7ns046nimJbpT1FC9lHjXZTInqFwAvcUbAmo
WvYsla4tvCFo8p7F6ybX34ET3iBqHtsWM0p/IODbWv5zc19b4g9XuEMXYHTZ
pXMEcR16oOpYzcY/RxS6rTw7otPvzCmozHEa7QRi02xkDDj3X83yJRbMoTI5
uHm/6n4ilUksPKZ/Ps3DwbPGFgIeBqDSPLvUsJtx8nl3vyNAGfc887sOlx+4
jn4CWREv4VOld9mft+aVzFP5bEwmw8yVx1yQEjozsa9XyY1eQXgs3A+X/WKt
Y2wyFMmkRSQ7MxSC7TEusAcHjoCIhYzPPBRw/LSPPnfmDyTI2Y92dGJo62u2
9DVfcax3ny8QJnv1/htY6+VYBJWFxTOe6/G3W47sCZX7TsN/1SuY3SiaIQRn
rthZRC5mEzcMjaLS9xTxBDuu9l1F3vK2s3YAopLRkjiAL4+6/xDqjBFAT/1d
1Fkb9bIl+Meg76Kv32aI05kt6CVxyjUbiCNCddSeY4dz9+8QtvCWODf/mVL2
7DN5KrhN8P1eZxs2bGQtl88cuXrc070nxflX8LgAhT2mfHvx2RdsYcoPtIoT
sQKJRDOQLpIPAcS77HoJJIm4QrvwK0J91WFpEXLdzCxwOUwvnMUEJmF08Bqc
SUAhB8Kk9hhNhK2O2OTnggIaUNKQOaPcwWJhwd+6acCrO6bbFtbH3lBK0h3E
8Dnlfp4PtXKnnmHbzJfexv48tNPuetG2Ro+0oYzhwnzpr+lawDRICFZa7DoD
CDhS/iVnLp6IyVpRED+33vtgVlJXKmsABgvBtXHa/4ZxXaXWkXg9OPFsEOaj
ufg0ebzw/fWRyBUJwTbvu+g3u/xuDzw7eLB6gubHVsRCcWUJbWA8X+MUDpVm
fUit0magpS1l1znOaPP1ZUkUkUckff7TL83mSJR+9xXaANVSHEY8/XnhQsMo
bA8snE2xUxQrETxNYpJQkQ3Ald9Ix+qeOspsTdW1nYlfGMafMQnPF2TBOUv7
3URSYzmWoP+qiu1oNqaHAoeJ/VzP1Enab4IPcv6xlRLaIr2Nj39lSi1rf2KD
f7IPecEelyGj/E0z4qEGe62j+jxo8aZPMzRgBQPufXln38qqDfDsLw6xoCSA
exWZCF7TeXrFAe5AJ2fJ7Q3MzJbSIKP08MpzDVeql1FH3jsewpglPyWqwB21
ud0RqcP+0reEwPRpi2hPiKkTucVAYvkfwoUab0n5CU7UoPsjQHAJX+FfZySq
NO5TLhUorgDKibAgantGc8tPFp7sWUsvTtpEXv8ebaj/x1SkeMHkOoCoe+d3
aiADDXL+BfcwuSzsTCShhFHf+TyAXsQThuHvXA1MXiEXZjxogjWX4EXETF0L
/kykDFnP8hITCFALdQIXYWOcJ/EEhFZwZ7UMqcopnOQeyjEmPc4ac7/K3lWJ
okaftA0Nswyv2ylGxZ7DPwrxmta88iEx5p/rUjnGSpFZU0LqB/gO8EjVPsDL
q0FBi2/K3SVdCaNsQuZeJL+Orx8QVo9JJHcdH2slajfLQWkt2O9pBtZzR+0S
agNXlsHG3HskawiYr56A5VNG/9vWCcHZIA/agltdF7/Rc7/LyPpJmhypGFMx
NsvxUPTn6rGrZsBwNe+74tPFjTsm0PdKUkwuLGy+xJu0sFlWOveoW3F/RcCV
TimZQohJObYkcp6hYPDssLBN7hSX6RyLlU53iAlHaR7cdhW1R2ICNgsMm8jU
G7WAFQ/opT6ncinzi7xhihzwBPtv232IFmpoX/MI4UbLlp5TFEl6oJYPBIgM
08P0HqUxQb1oLvlN13+ftojsvqKNUFRLsOIzG7AgXapM1O8COByuQDlPJCe5
Izx3hxh0g56SZzhwNETVhdyeOAtLm0zn4Mcv+NQgMR7d6S9K2f6B9Yilq59P
RbN5TjRDv9YE8/B7/eaFKUHI+h/HgsY1Zk6PppKwNvP9ZgW6fW7ewbYiHEjs
shzMsT8WhWHWqeqQf8ZCMRsvGZfWj4iHIOr7MCZ/LDiqgSu7DS3uBs2hyt8p
cxOhhPHz6X4jKWzAtvoPKOrDbMIZmj2l18x+UEsd5rJ2OR801h9RoOTjcW+k
GIiGYnB4jZOjoXviqa8YJf5NGeWIyltLVq292FnmpaAgtanpeb1alQem/hPZ
x6zeH0FknD4xTD3OvRQGG7RZFhzKnivwkF5xlDTzwqzZ/5+VHEztIh8TGUdt
SIyn4ezOj6Vs0c5tuTsxt6mW2clB0/gI0sCOMnb1BbTtgcIV8MSvKORKRUd6
FPTay7N8kOaoVLorx1i8SMT3a1MaxwwBmTrqb6eykvd/Ad9FhtS6MTDYaYSC
HJ75LA+r2Du8pdtJ9GyLNIHX0Hy6tu3pDaCW/GBXfFf285UklK4WcvQowfK8
rxCJX81ULGzhEq6WIimtIMcke8e6vMOzeTGf0fdEgk8WEowuKqmeSNuc1yW8
6/DS2ep5DqjLRdQnmiRxxBbuf6b56LYbv8+IuCUVtB1Sf/NIp13bTEz5rl+X
KMhhFwg+SipzQx6lgeNTbpalsS4p87gmBS9LFWLt50TYfw3n79VexFtRM38u
4YZgD3JZr4+fhxsaZT86UwBHbkUf85pIj/lsJNCLwsWmcQeDdFX3QNZ0IzNK
jQpO8vzy/sEwWvZyu2TuXvVF0J2mGPn8h/tXzeQGoQA7kpCYSm6YJOVmn0Uh
9ol6jewDKZHDiwlFslzp/+gJl+sy84lBTZwvjUBTGVdg9A0EnX5sqFtMKRyq
Ekr52C4AFKHCsA0bMPNDiVIY/OZDBwWRaYBa7DZ/vLZFWdQbjeiOO7teVOxG
HDdPGGFIWLp4N3DrVpMfa++GIRVlwuG90GSbWimuX0xHvFmREDPk99rl72Ok
2R7GbdLFgdjsApWn+8+XiAaeh6HtiQ24bF65kAGtO23q7vy3mcQSFIwciJ+f
oR/kXpKZywI2jNyLfXgQdSucK/F+R28PVDvNjDef1MgB/zZRrhxE2dt2XzeZ
ryEaQ/nuJ/JCPbEO+xUx1y5qB3xstoA9V2z9JZngYlTW7dsbcpTbQ4RfVMTR
b8eN6ysA1KkAHSR1u6wsqUhBRUzd6UpJgPO76l+wXQ4+0ymSgFCK/8BXjB9v
wc2/6s942yduYbtaNcCpNw6CytJgRK60ToWJlDXTenryx4LS7onrXzkx2l0F
qPtK8Mb1OOfJSyia8pQIgPO0I48NkAzwrBTTXZB0lu0R9eS4u85YU8o57yfK
+zHxhdmAXzUwbVvNPa8kxHV4rGCKeYTjWdN22oHrFkOijXVxMVL2ZsAgWAJK
hTiomM7Ja0tDdKTH532wnGaJ+MZsf0DBt/Tpk2WOyVahzUoMOOoCDfdaQFp7
9XBzRWKOmU3SEL5n5XFRL5TVVDkpJr3LL2dUEfgspkTlWhINXLMDO0rG8Ps2
IpmR/8zOOY8Gnff+YuDMHMC5LADmVuANR2WSY77mGjEmLZ1RxZWPw7XJICyr
E6Vp//+rFMVxQzzja3M1WLnAt2g84UgqjaZdQoOFN+5/v/FHkTtuCjBmSpKm
+NM5yTjGV4xbPqalH/vRP4Lh1sVeAQOPErPMZ3LwMdjDmhy4IDl+zHYhPXec
7GUklENkQmDStJ3Nsygjna7mikiXy166UdJl6jYVR8SNpRav1TvklaW1xY/g
hRR+Oh6OXA3/tLnDRWnGMHrKN8ICf/K0QxMXU5ZRNejgPePT3r+2Ayk6UyCM
cmKpWesiOOKpzTLG371xoRPlWQ8xs5sd7JkCVV+8wP2JG5jrHifDTinNhF99
RdDB/817ZLrkQ7259UpHPDD3lm8iZw7tsYScvxnP6NOkSfRR21ceqPCEl57D
PI1RdQzoZN71exO/zL3Lve5GxQJbjpkZ6cBNk6HZgu1B9eHnS4cO0GIMN9fp
0m595D0aaM/v24Rc2Rs4dm1FwgfxoiLccxEqW160/9CS0TGJx72PtgaT6HjN
pv9whxXlxfl6iXt4hsfi1ARsKIfgj31o+JptJTX5AsKS0RiT8gH/fdJQ8lFf
RT8JMx5cPXfPC30AMZAOpiw93K8og1GyYsvUI8O4vntwyaIeZpJ1GpHZWaNU
M5eCVgBmhiFqUDDWVYSI1TT3fgyWiev94kSsBsw95TR2gcicHc0dSsZck528
Trd3jAPg0lZbmPhy6/QsRkIcFIjn+K9nugdoPFhHy8JyBVftFYMdFVdc+i/v
kc8v8fFPdzpestJG0gOa2HiT9fmEpWtue4k7p63T44cg+lcZLEak52VQ4J/Y
+99KYERJF+tQuJuyuVIb6kU3os/m9MoHZkgJzvhkdjJX+sJPGzpwEeB4j1gy
PB0bPY7NthSln9Xd7BHoG7Gal2LM7VDQtaL6LxzzXZtQhSpjIY0uge+GhILY
OnjsPYjmaTmtXmlFBj1lGlv/Qz47awby6tO/8bkzaGT3URtlrwdYKq5t6kQJ
mUqYmQLhEWQFabiYF17Vl2OJLkKxFR9zJY0i8jryoA05o+qBv8nW9FvphDmx
sphfZM8xs3R1lBlzNoNJcZw3yvsFNjXRzIbavWHeIApIQ3fI8QTY9zsnqJIt
5dAxTSi2h2I4FLGVjd4JKdXiF4ACJ3yJ9H5J4ikOIL0siR9ytZRr9zQdk14W
kt8c06Iy5szDyytG+AGsLpFEvMoItYqzXFqj0o4jjlw9SKpfySDDLCG2gdes
y9aFn0Z0TT1LN74HCS3wNJ64xm6IbKUcF7b2t0JAJlZTVvg799L6lExupGcL
Hyu0Nr+VNTIhYBZ5LDrrmmjunnQ0hEuI2iImeuRKTCKts6Xb+jCbqFCQH6D9
OMmTFvZQyphMuCrEPFBFoPTae8w2Izg6gLMILmhzer//5P/aIJHIAaGWvlQD
unDy6lXfdhXz1OQc+1SBD/oBB3p3yVMWRJWCBM55VetaaijISulavjwZl06I
4rPqyUDvKuDspY1xN2iZdZxkwC9K1oJaN2XXTdHANUjIPFAId0bpmllr3D9x
aeAlNn/Tf+WFxdHYVh+CtBNJ+dV6/nI64KLcNLz116fKb9mfvlbq6fGz3OBq
i1Yx4ylMRZ6Rd3ToXG1wavSkLYa3vM+xoadBB3w9AkE/0+0rsBr3n2wtRFce
zP/8IzaFnv2kEozZp/iiAT+ODJFwgAOdHR9WiqRS2RpMqHDAWAYCb4mu6HzG
nqyV4hgS76mDJIyCeRe/345c03uDjR1yfKS1BVhdZ3ptIj1a79XlqBUmjaQi
cooOfYrFNabAHIV99kMW9PNbgYdNGjmXE1VkR4rHnYVTsixIquUjjjZTWA51
YAqSYguDlj0HdlAkrgked2Cgx0C2AftLFP7dBEG5P0VD2PRByKfD8SOCu4ty
zeZxMUht+8Anr1uD4/WqexOMBgsSrXULjWqPgQ9WsilszvTP5mmEZgW+Df8a
8ul45JHkH5gxDKAMXG88UwBV+RNqiDxL1pGS2ibZSqggXaugKLPBPXdAsx5t
jAGcaLLD6oIrdnyhecqi+/obld9izGnNhQBfITGUyZZDS6TmKJ/8Nq2pb8rc
SDXuBsXueyivEhROx2B7vKlVtOlEpDDCxTWqQeuYGUBFZNqrtDdhCCW7mZx/
M7JOp+i/dKRn/VmNBXVgkRMCtDpPvDM6VTePt6Irvi2luI11U0fQNPFVHLyR
ZhIrYtscienb6RXh2wpgmI7RHq42N/HtTG0MeGlFSHQQDdTmuOvFZJNYfylo
R2DlNW3qHVjCexETPkFWuhapHl/wAvXpsw/8YHxz2aE/53r5y14UVUZb0CfU
K77WDmz/BRISeKSeLTahbpjMs8s94/clVFoFCtyPBsIqNmPH12m/auon6Llu
WHNBPR9j0VSrfw+NP/7jWkFUi5LKXj3gdXW4uxdEv1bzW2TSBt3Lvd7AeCwr
6p5EYVX3GQPjM5vnwwbAAeI1cM1+3mlC+QOHYSJUNCUHNojQRWEk1S0HslJ3
C2iyP1rjzrg8QWOCOHBXlsXZt6SAOd7T9WBbdcSLZUYySIFP4DBKQyIpjFpT
Fc0ZOJmOmHm/EdgixOVznfWyIG8m3EN97rHkcnh1ikfgwbSGPcH6EEwkU9IV
0Tyil4JjsOKI937N7XbUaUCBLVmCiEHr+/Z/7y1CM5nD3uivzPWc8XiyPAGE
ZYBLqG/LnZ50zlc4s91S84vxSxSkQaVMwEcmMw9EjnD6CbYDMZaQOcP4+sd1
m0d2OOKXJ9PCXOO2Q9bwdTAzS4BoJzUKeNqvumobyLGrTDNZKLnTxGyb0hlm
0OWp9IfslxcKKhj/H6BTrfAC6dzHgUV0+4fJtpMm9C+rBiuYrf6rJc+WYW41
qa1CW6oRWBk7FgzVq9WpE4YPSZ8dGe7be898fH/ZDDC5uEgfxxf2NUvFtl/W
DoDGJTDesUakwuj63DNlEvYkGpgCR0zCWnLPp62lomiW4tirRxmba7PC24MQ
BG0L2dHUgrnml5yY2l9/ANXymt2Ngbdt0n1JIybKr+lW7OyvhYBI/ph+2/J4
W6ERrBQJw9O1qYAshYK5afimNk7yixjiI2Zvy3fsETYU9oBfylIurd6icSMx
zc9LPCGru7VC4yTrBDSsLdqQGrc1TUkiQT1pI/D8hZgK3SZOufG3uvyoBlha
Boh5IDi6DaRDo6KYtn2aS/vtH7K2B9mySgXRSWz7OVJqESpX7yCQyrK3yRVA
lvvGIeDKKxbb94RjhwKPFiWVXr1uxfvFbpF8TMOyd3XS2EqP1DkdoP4z5RNS
1vvfpl4tJ2zSjDH/1aWRDOO1p/OcGJS9fKgay7ChRriRZGIMEYv3szwV2nPe
QvGmNzsvAADY8ZI3KTzgz1nJYnIrda0tOx1PYeL8kQVKyL7C7QSdKDVMhX1a
xUGY8kpIflsCqxUEIgf39AJSg5pK0SlnIDbvUQZn7iaNcP2X8/ozzMAC1EZn
+bMtrS40ziOnY2ABTCRDlvvVY8OFE60M4TcDj0dC5zddbq9xlnjYoYujMU5h
6QD7rCNfV6Asw12srw/TReazPXR2BdVJ56smMG1bapQPEH6t2MmpTb9rpTgp
itq0k1z4V1acmPyAtg9Dv6bwiqhnI+4hn9Kmg/mSBigDNEQ0CswWmrVpsjtU
r0ek55Bt5u6Y6h8Sk7HyYIwXGRW/nMG8Rirl2qDpaD5lLKwVQ3UdCZfSiW5f
q2nVWpRmej/23/5/XDc6tHFBh8tCfpX0TcHg/sHEMMkcCnW8E442zCvzkTcS
R2ub3LRMEQFNmdXKYSMIcw+eUt7bn+5i68niSWdpnSXBHiDP8dMYZDRRKcil
etv8OXbOfEB9H+7Q647/reDgMUZJv9xkTETI2/rR+2lWB6xLsY5WZUiI4lnA
WfE82QTsTK2L7/A78+YpWAX+YUL6rshc4188fwDVDB5NPyFZTByM35DaN06Z
6yT9P136UL1hNwfnBuYpzt3XFm8P3w4wJvsFaxJsIGq2EGRMJt5LqkQ1sUKg
Ioj/z3Bdbwfn50HkcfFG6MVcyaDP/TwqJPFCMJtmUCJGaOFV4zST2yg/+PeZ
4W0ysrHi2X7uwLwG+7Gsj1+sIuymPYWNnDnbtEYJGlQCPcZ3G3YpNXf8zmic
pLllr3wiiPFmbUTgculpvU5hwqhJabQmzmEXo21gxTWBYh3triSkm9+xHPtA
dN6hU9m5v33zRVh/JlcSvf0XPIADzz47kuEvz13fFtWHe3Y+LVZFlpHog6lz
z6P2PzRfea6iLR6d5CJOgt1ffUyczWg1bpzXI7XZGQ5I9sg2yebOVkFbfnvm
YoKRwFLq/VXTeTmKJySqj3QjyGqXSsHbq8/DwUSJOOltGMKjcMLcXa6k5PXS
ejelXxHOZYJjvTiR5HHQacaONU0DL/sUS+0YEg51btBaMpFkgvxICculLeqA
aFDFqHPU93vBpTOm/TGgyj39ussMHxayFs2wBubGaebANBlohZrWx8RBzfVZ
UJQ4edO5VTzRTw2DX+YtPG0c+YABzVr0sIHVC3KwxMXZnlaH2DP9os+Y7FF1
FYDvDPLUR35e9AbESjf/Ocd8qjLCQcNP8o2z3o8tJbhgLF64B8MJ4Le1RMaa
Pdq5ZOxjz9uKDzu48wfs7pjPN5zbpO8pU57jSBRXtz++UtzkkufYGBeqcqTZ
HTAXmISlnE+L4cZ9hKgJDN310plO3ublAKLGHmleXVuQxi2+AAULRCobERgK
7PL0oGQETxKY3OYYHL5Sh1ESMXfZeVFsRvnHcsbkhsl5rUNiZEkKyIWyqeIw
6ZeBjsksLxjcvTFjOJecFUg/jNuYgV1R2Q6HMQX3/Hwby/46Pv7zWyVCHxmN
Oe5FZT2yPbXe8aApLP1k0DBewZ9idh+Zn1+BCi/YVHcUwqf631NDPdNeDO9X
fQueJK1uuugF5Sndob7hNqKBlVmLcguNB/HZ4bslEVO+XkjVGEJuuXUBPonK
E+tGAyqV1OfIO0UIMqA5Wlg2E1mE3lHLnx4nn9SREJDtEAKM9sLb1OAC+WxE
uGg/Y3/52X2s8IWnmnFvARuGO6oIPY7BgAUI0zA2RlL7jfX6cQB9ssbi29UJ
MJ73O7HIxH2oIS1NTN8Z642I6QX8QW9DgifUtJkRckXm/y4ritRpp0OBKZW7
T61zVOyOC4J4ffusG0P6CEJaKV72jH1TPziaIBvRjqx0cD3zGraSy3WizuLf
s0mYDZL7ASJtf1yR0ZqoU1MxVinOOci6crM8talNfp9hze8Yub4nq/+dBfu4
D91pyX2DHh+haGjBpxl9+adAxNJain9cZkh8z+BeLu0KpfoIeEwFo60nWbsr
oIyRhTpdO/3mHyHBA9N401xEAkhPLjsdqSsYbpwLxtgJ+P1bULKqMQPwCrd3
wTpcRH01APs6Pwfg5nAiVG/5L4cyHIXp6zT99Wd/8i3DkRkNyneb4kKcVR30
GUm/3MDobK9/H48HZUV4jY6Nya5iG7tABansAUB0zHFH1ziJn3b/xX5QDLJE
7N8t2Pnrg3mRdVhdK5p7hpaFXRRFwDWaF6pUJNQtIMEms0InQvHsDTg8j5pp
7tg72R1tyasQVzvOvrMw/AwSn4wkd2XgVm79kRu/R6kclmY3FT3svHLyGMA7
duMfNkeV4bSIgvagTYd3V0qA69gP777RddOQtV7FazlLaInp66ip3pZz2jvb
IxNWAiJ00Cdqqj63ey2Ehjavxbb9F5k8yILpBcdi57pUXU2O4UsFcpHCFFp8
qrY90tnPeuv43YCyJyH44VLVKFtruZOqPnX/Rrkwhv3ABpzS0y3cf77bDX7h
CNC9kwgA5Lpr0VQ5NlTOr8494/RoEqr0wIVD/3SFyJaxA9ujzSrbvQjiCGZy
P0YyiuqoWKXZ0X4ZVgA2+thxEM/3FFv/MTsQzvwk/RDSHAgOcC+OzCepgfZ7
pfUEUbtRrkvWiN+CCWBXyBT2OPbvw2NY03KwfJUUbo/vhk0mrdxtNlPkJQcO
mncXLuPsijt9SXm1ZXgLZaJFTOrVEJk88NBbECtMRoe6+IgrU5Ab6nJ9/6rZ
oIQhqlD/fALybjjRNDUVHq+H+YNStWw1KyV2ZB38Md65j41qAS7k8O1PJNvj
9WMUwg9A72dgO//1c7AzK+djS6dNtt1LlmKBe8VDB/2RHfzzqEvAxHow3wd3
OmfOLFtZxVZgOInsDPcqG7Afc3Y+5+XFVb2OiFoTq/Sk56l6uw/OpROoTRZk
+bPupU5ESjk1VkHWrTivJxPsffw7x2TsrqJiVP8XZ+PNJHjB4B4L431tpEKX
BDY9lahvtOmMtAioQsK/i6KRJ/5qgg2w1qi69nTye4kD2QMSZsNVWWdFmU9C
4YvsQvpSGZpOrsnMKCRZ1l1y7PdzaHkcg49yQHtOgobrZA0YW2xMenQ3JaXe
ySEskSS0Y/HHmc7mKEDvIER4+UY6J602Eqn6omPVPOSw6PYgvaIIqSBOl7S2
4V5aXew9jJek5ai1JFfy8i8wyUz7R0i01/58cfjYHV164SRziXYNBRQBqCoj
rAY6lti3uinKJHsYnworX88ujhXePfRQI78S3KXAbJttooKbLMlFDasxsc2h
8u8LSUuqBjEGDBRGi4ugKQaj4J9vWurXEHQBt0yx9HIJeBkQAATuh176PVoL
JuiJGyC4b/23qznoD7J4nMrOMPTpDbhs9fHd7iKFr1I7nQULxONSxer04m/m
bvh0fe3Ut+Bv2qyUO73V2dw2gCJibIdqoNNnExQuu61GpHPpXID+DNvoKk7S
OE9DVsqZCcWZY85nZnMHlLXDdg3shMhoSRhTPQ29nwVDGqxj4CGfw4d9gknA
57ORPW2TMHvlWF67TegjD55BrJNfmTYm5XrkbpTnaDJeOX4rWkvYISuPqlVz
cdYlc49nkYXeHcQ1LThTNsdhhNY7lyMJw9D2bOXmPTW3KBmqxRelKWJpymmK
8NmZVPNIPwvU+H8d1fu7mCNpTqBifm7Jmsz8CY9UqKXGqHcBlNCUSkLAh9LQ
x4LV4LpKeeJsLVB9UKDbrMqZs3eHaww1McCZ7dX4ac4illsDsJxJfTNiVi7T
uC/hbc/kmaC6qJWhBOSwgRMyNDLMDuXLPl/CzL73KIAeUxOx8SXr8Sn0i/Dw
ioNs4agkFneTDSqOpmHnq4p+A2MpqYl82VJOufgw6w+0UM4UCruphYZAcR+1
zKE/B++VbdOGRpFXZXIhZDX+56y40JwI+JUJarcVjloHgSIHuYSuMSz0/Zs/
rm6dhSuWczhxyxZ9JdzZ/iJ6xoV+4R3+678i/b7HUdZE4N/RPEfyqVjm6X2p
h03VA+5jAQ0/XwyIkHDCJ5uMZFgnHlyaHSN4NJv/lMfif3dsSRoW0Tu8YtXa
BLyXE6AMuu368KMfLrBvhdAMsnl2wnZSlIFA7qgEu/fdPP3/VzKQF/QMPOQ7
QYERy4jN/aGE6Ob1c0qNlHnQG2j27j4LzjBdYXnLVXW2cSlaz9owZVjzvyQv
1gbIDOfdkp36UD5feK3x1h0IHRRJ0gNf8ZIL7UwcXfVcO/+niHb2kV2Awx+p
aXtLZhEza8+pXW8+lmll9XMQy+4kySmv8xYI8GxOYYtuBG4R4UVq28Lhelaq
ayZoy/kNFNXuXqp4kmFV6w8Frbzr/wkzHcsgYTL9ERjMSijAUAtE6OclSupL
7RgJSXqlTPx5Bf1TJOn4qUyr/k0jLpNwn1RqviXmVBwkm50gszQHSCXWziXK
a5fp15aRJ/9+b1KcpH3654MKvQhaK2ipPh3W00h3UVvyJgsUQR4s6MVRLkZp
nNqsNvPp4oH10tuDWQsnIywEchqr/oL07F34qGyUWbsBjE8qo5a4EnnmlM2r
L4z53kbnLb9eawARjVaF2ZMo3+szP4lFcVgoWAkrF4PCVkeotGri1HdVnVae
amhSAjlrFT6AqVzhQUz/WkeL506JNH8qZqRd0EHPE2/snCFkEzzZKfpsvWj1
RiBrGSp2wQFJKOYMrNZdGYYucWQSMOwcUhfyA1ol1ndw4+epMAvKR5RQet4r
am3HBzJACFi0zYXmLw+j8/XacK85ZbARfmQT632XsYXAB2RwJJv09sNDXQaG
5JebCqdAPa7P5XkCrTv30XFB+mVZ3ZU2PbvTYAhssDTye2KUb2c0RhKVBwyh
pHp43OXSFK8+Ps47phyv5zlbE7pjk9CTdF3uo2MZsTZrneKa4PnYtFSym2vz
RGniN+o2oMYM5hTMtuSAzi2QYg4BvJFd067sLnsSdmoVM3/8/rEelJjIcbrl
WPYYLz8pnDVJqdQ6ueJZImyHdZgte4BWCZFJIjl/p7lPS/KvAxHVmqCPcymD
xbk2SBcCeclhUXC97ArxcU5moHu+hx4dSWo+oAtIEAfRaClZQGysESBbxfDZ
lKq47PdGSRBZxUbwsB6daKqnyJQRf7SYHL13LtruBK7AFqoq5BAQy49y6ayc
KBuj90MY7wAujeW7jNxSvYuySret4fhsyR6j3i/s1y0syK3VWgsti5Tb0rBv
G6mucACftYHT/yaJEsLgmfaEd5Js/5UGlxTL4ou6tboWg2JPgyewODz221tE
Nr/dNAv3aWiVseGvHJQ8kx4Lihzo+cqBU90V95kg54+ycfbuhvYYEtwmLvv4
TUwApUuFWHLOfg4j8oZwTCVZJblBf8fQH4ILu/MFxMUeOgyTyXnV1hI8nEQc
MJAQ8sc0dVBFAaRBJuM6Kum2mUY5+LuIfyD+bBnF2IZcrdR4B3G7Iz1dadJI
lcZZGGbU0vt2cd+ijZaJGk7wYoWpXt8midat0zID8Nx07TAePc4ujmqXXNf+
ISbEpEj5idTLTunIt8HEM+WPW1yl25n0gtkjpSnAnvNU7PRtnqxfyR7LeXy3
Rqi4bzaZaNs9TceXBwEvP5T2g63F0z8G1i0OomdGrSzAZrhFAZ+kP1NCCeuO
9YH5XkUmq0lG+rGUmTPkQ7BD+J4CeiGjx3+EBvMiwX9hNQIq0MbXsI/4iJU0
WkHMNqXtrRjlM9X52N56Xr1eURAPIOlvoANf5Givy0PHofLVQjQWGDW7ZAZf
8XkypWMVecXBGEcUBpgDMJfzRhqNLQIt6i1SoqkGrjJ16gJcKM/RTCTHYOpj
F7qmeoLxgju+R6/ie1FEIPIKX1DF8BKx6Zomj0lrArqApW1rohLW3ItEmKkB
nYLZBEZzL9J01uMyEJMvBatsPXGahVCimkZnqbsbARhXQ4ebaUEX5LGGCbkq
8haHBOZmlqqRdtFIXHf3mKEtl9liWBI24bc7/uzBSMBrU45prBQ+spBM8Aoj
W9tMLBZGfd0ffBhBPYA7Cv3ErScKRtFkv9JfR/Le0gmhG9KfxfsHYuFilzI5
6BSIWr5iVBqjyj3QKlh8iuLGO1v3CutvEPj+BWFlvIsK4m0pEWjVzPJuLrrh
GtIHCiRLrtMEkS32BghDq6QJWyyomoLLtfZNsOgPH+oKcGyoiiyGJjJ8+id2
jMlljronZNpm1yaPs2Su8hY8YxRi7iypiblgYZEjIuKYDVHqxXEHWy2xCgnr
iK7p+m0c+FMawnHDfmC6Or+4Tw/e5tfo293SbifhJYD51MHYWQ6fKT/YUo1I
IlCUnnpdMxZceuXRyKFXua7ijsEaUgjwhHbTAVLUKcLV0XtsNBWGhfNKy++C
OJxNrMblb6cwNsnT29LzH65KKzc/36FA+iujMMG3NfejEAo121e86PvyuXPb
UUgU+BbHdnp4QUQvJFZPvwNsx8+mfs84wvHj7x5txADusGI/nXwl/zcWS3jr
leTKonw3NvzdQ8Fbj+MuKJqo6EzN/5Ar95luR3JcdtWmXuwjBpOMG6kgmLkG
JphWRMLpv4OGiP9CYoPYIw8SJUG5K49b3yMCz5S9FCENhalU9SdOc3EMFy39
RzU98jX3B2dDUJoYbBe+NDrPyXwpqhe87D9czHUbl38KhZkxx1pLw/hIYjRg
hXvvMIdnJMgiMVFt2JEJxUAqWqLOaz+75g+3B5cp6VYSmfrbcJdotPaDMamT
R2ViRd6aD5TCIIP1TFJhkDFzL8UA81x+gHQSK1lIjKE8oRe3XxS4DBlmXBpV
I3HxosXdW5I1erkIRfzmPk8QUY1qs3MRKzJfIiB05g40oBSiOh4FhfPc5P1J
kYsMn/eZzP03wzhBRq87lHQ2eLAptJVfKJStdVNsDOsZ45ex9/ZGQk+7+TMo
W5bAHTymKME5GQeNevmIu5ViAyRk47KCN6bM0NNum3B2kCXqtLV6sjeEcPaR
qRTMBa/fmNNrDJg8Q/BrsGptfUglU+2nuLnIePwcEg9XPdycXavVnhKkpI/f
VzbAD65wxSFqCZtw+AOiFw0LyiyrjUbS5nluyYoIpkaf92FjOhZvnsLwUo5+
3t8uloep69fMncfADkzYCWfNRHTtjtyeMEPOCr2B5YkWVPFWR3IKjORqdEeL
rHXhbh26/3e3C9Df/AI4lnwVzcTEHwrrVGS4lX22YJEHMDPueGpyrDSydLpV
8EHOl0hK8Z5gKjueqz5GbhoCdTK7jaqfC3fgDohmqCjq0jqii6gGJwMHEevn
wJxP9zXQhFI5jhIJrVmZe/3sc6o9DPhFb0yxqmQIkz/7XWlUov1fd5z+RVFV
Wy8Ym1v7/uLBa1OHnR/KXa1ptJ1/4Y/Qud1M2v7s5Qyx5N9ksQJWrfOniB4P
jaXBFE9JkDcrtlSV0/G+p69V1UVHFMZFyrrpSJPT+o6rxAdEgM7Q3ONoE9TX
nbFy+TSJ6PesqZ1ZPS4FWiAAzXY/y4V1l2UFpWgMFrRg5yt9+II+BYuJYlf2
O3yCQEI9NZCUttUebkD5iO97LPmsmfK5t6fdKoccTot+XwBdQp2K+1PL6A/x
KGoFvCMP0FlUS6BAB120qK/gpZim0i8aQcysgKr8hNYWMvnpBJcWlNGuGJSd
pVGwbQkhJpf072fdhxRQWco0GsZBuwk7d9Zuriajk+maN8HpbnaPCZu8EyX6
Ss0JtnLC+H2BjKFy1JvwvYN7xU3Wvf/aZkYEpOQDksKEj00Pi5QczQz7TMks
0icAMfW4R73Uns3Qa0M7fOzEWDE5AYnCPKoxnXnLPwXiSWh8MnXZs5m33tnZ
Te0HUtSeci8jvnm2U8cX3pyisfZkKyjLYWqThSeI+j20WPwiCFhAuSFFGetU
uNyb5IdRSW+RWJZMLvVDS1A+Cc9iF0iUO+DBHDkfU+o+wkki/RWg4MMWCinA
Mx+aJtlvz+myBDf3sovkLESW0xD/o+34vTNjmu+41+bPoarOstCR8w0LGKd7
sjZlTbj7rt91rbjq5/dM/6SZv2SkVksm9pOPBAzJb4gWWm8OebBRa7oo6uPO
bT4mme1eVV/ilmXPoKl3UQMc6f1jmBq2e75vGlO82fnNeWiuDhipkfcQglwO
qc8ku09jo86omM3jQNlaW1b03EIbLxYie8gG2bmlMEImqL1Wo4p7k1iTwXnD
ROy4prwkOrdDefkgHxATtXPMSIs4z2QXFi/4fZt1SBSXS26Z1YhZb5GjdHnU
LHSlh1ugKL3E09fLGYRknDSCEYmrvvAS/iVg1G1S202gZCtpTIX9MDtP7nLf
/qFFCtWdQe/orRf0TKkCOE8vFTxnrmGh9tc1+3NifaKrsTFd4aMexsNM1j7q
Xm3o7LKOxz6YgULSln9nm2z2MIJC5NbzYGXnHFJff24f6ZSoxPGOggwWVvJJ
WBNyObpA9PszE+C9zUxuX+78U6WEbwM1SE65sSCyDm8PhLKZLu2udAm9FFBD
60iXOGCnrzml2SIMus+zp8PvyTzxEJk1OeHODBxp89HhazYg0+dsbdggD+sK
oSUC0B+oOQSM7Q1TsKbG9Blb70kh2QblMBOYsNfDQo+Et38mnUS8GK4i5zMa
Rf1pTpP3FUwj3nU6aRODt2tEP9Oo1TYgjpurd1QHWEsbp14QLcC6HxgeFRoX
5NOE2vaAw2MPWz3Np50iceW1zle7GwYZqrK9j73Cs8oYM4x0I8Y6Oxf+bh2A
tNJxpw5trsmHem4QYKfVf9ph+98tRbQDcaWTzBeGVK0DzH12wkvxIqlhiz2u
nmpyJaNsN2lwCEL7oRllJdEIkvbYKtSSUAD2GG6dZTsKEnsOpBMJcImTvvlT
yt00YBWmr4OUfdKL5VeBqojuAYLsUyHllmphtAxfHm6do43HdIE2BTXEfh/9
DRiltiC+IaZX7wo3Eg0mJa/8QvTrIhgVtJp+rEY53bQVYaBO5G0tbCRqwR7a
M1d6YJl53DgfVg8b294GxoY7M63c47dVeLcrd3k5i7EzTgfZDjMzyHmGMFTO
WYDX69C6evY/5+fxhKP2hNsWYu82m0Sc11XHOoL2MBDaEAtaaFjd2piHduBh
Zpp7vkXonQLkkS4OJ8nIXtu6tNMwjB0CiLHKGYCoFndua2vjsBHqLPmDc2nG
hNWqR4us4ntYpoz/Bx/dX7BLw6oIZO39LWVx4XrL86+MxmyY+3+BAm23OGHL
eBisNPDhG5PtyJDGbg2pOt/d7qX6UmducQJ1wREZiit1VECJQXBTw+BlxSg4
ZAVVZCtHu7/xAY5vVpA62H4Mh77hPjlmGkd6nRmpZUkbl16xjh9Js20MNIa6
XY23VfsNsqFaHNkGbnqcLqGVHjsuWSamfqoC3Lg/AeMdsHDw1oIR+kR+IONp
Xz0UEnbrqbpJClfN291WnaIPX78SE8A/OQldlkeCd0nIDWQNn9Dhf2ZqsJSf
rnTVdPZX3ws90Vmht+hrMNVpfdErpBO8OHblw/wToT+u0vbCxfVbVCwX4MDe
PuKVpMtLSolOQqCRGAoB0SB8FZR/3YpCmdfOjB3W+8qD01wnKWPEo7CXRblL
klMscGgI7NIYcI8GXASMob21QCeFBTTZt+JgS8zWkdz8gQEz9hnQFrpNah1C
DHYLE6V4u1/fEicrOOf4h5k5YbYZ/u+1lG1qTt0+CLU5SEEQys40TYsKRZiq
VpdYXrxc57SFKXI7Nf8XhWw8HPOvN8AHSvah+6d0u19iKUI0rWrnl7WysiIj
gbYiqtwO9R/WXYFFnFW2oNly7diicJ1sBDyrGmLmNH9ainHDma6b4FnGyD2P
6NNnXdbp5ZnCZbrhbSQruUrq5EL0N0x0WkOjNgndXhYfvMWTzKI364ePOWig
JnMwPD7+4C6PjIXCDpGBTYT7b32GmsIaTTp+Jz95V+9ukHb8SgqKleSA0xgk
U1MBTKl0+Y8DN5axENZVlJJFdRt/iiaOgNtHIcdKZVn5glmnk9eMZdfErz3I
LoYmSiHoloK1Jo5ntY0/Clpec/+1DdrNC/MriidtaNnuIyrz42WvIA+u9FXR
QFrIGfBchYq8LvuQOQFqGSlaDO/03qW7d+MZk0aglah4Hl1qVKGfaibIhebC
RKcO/Okgb38y9o2ElZIYU23RZUIzFpk6uFvKbq5gmyHIEpTNkIbiNKd7sdn3
iB1UT4y3j5xyjo8EJsNkt0A18i1qBnzXm0wTIy3ty2przkNorjkRwxIc0SWq
SNujFVRmRRg0Hyqsh6JFBy79nIfYqEKZj75H75wMTxhXlTnulouUDy9oP16f
n6sjbNShrUIeTP1LEJhLhS77vRG/5qoq4ZKY8Dh6Ps+O7r2GXNtM9JNWA4lW
BmH3CdSCf/piTSX6rvqntpNaLaU1fb+ubN34F1HGZsyNoluAZ4PshotQz0Bf
2CDcavi9fGHDS/q5NXgfn0/749NzlMY98k32lOsw5Z8h2lBAqwqpX75iXQ3M
gZ34anT+/bp4niWkS9A14akesKK5k8pj2ZEMy+FZWXbDmMDzdVTNqCobjfgP
H79j+Hr8/cHU+/BeMSyURC4VJt36dhWexd2tU0hdg+OWG++NmRmAxH1cUKAI
2eL/Y928DCLddpwVJgqZeMjGsfw7rrPoIAXi+7op0fBdv0Wjei57LYxSTkhA
3zHoxRIyK4uI3CTGCPcSBxhzIUhIlKKRDEiyvV8maKVDTkVQKInAd1m/LVJt
auQFCPqR2L4I04+YkOD9bkO1ovFr8vxCP9Mu/CIsSVXZmLc4X/AubEJMumvg
X2V8BGojjrfYWKHXrnQdHQ3Gl+BzRR3Q6A4U/Ff6/wfZQ/Gs+kC+rWGyMowk
w8NcZBjFw5zWDoT+sDlFx8clGJMDCmmIt/UoBGMAwbD6pvQD/XspHy4Yr7Tp
yxf2JxmnupPrEpe0S8fWRfDDRC2IERrHkLadtCr2y8LgXcxvlNXoW0PCZ2SZ
9I/6snytVy1wknmV00BSx24wIp+C0+twiLGjC1XE+NJCGc5keDX+/6LLrGqj
7keUo5GBt1bUZedWVaeCoJ3AzaSu6Bg5IV7eYdGUM1cfBcMTQrLPkoo9klBH
Mpc2wmdNmaBGetQb7k4cMSlBw2OTWPyU+n0ghC922Uv7emj+YbT2P0X97HR/
nulv1/bj/ma35XdIcJXtIFMIvN6i4ZNTSVqVOSiewXsk8i7G46pXLAL8HILV
RrNKN14FcLPhWyigl98glDkMfixWj1YckThs/ewOQ/ab/ulm6PZGuPup+K7j
rtfXhK182NjIDrVfZGb8/cgtGJkArGfEATHLrVfSStYQshkmtH2b4pIUNDvQ
vFEu935X0y66OUXB0nkv5XffeHYip8xuqwPh1WVbMPp4OPn1HpYHLR0E8/Rb
BD0qptUIY6dpeG2Gxnz7cKSoKosHw6Y3EyfKKfm9PDVErvexMdZNWjwaX+5p
LYNA2p810f824g591szMrl9wmB4bzH4FCXhCCqmxrogDhXG+p+uicoLf9E5v
7EQQINH5Tt6SqXLwc6gylQqyJhnPCceUewB7vh11CTE95r50hzxuMVU2FL4H
jXTGx/JBQIzixkyPtqQPUaz3RmUmOivT7ya6ZuOQGm5OerTemYOrjc5cr2Re
Qf8xdJyv4dighRI+mtikXUUwH48rVRAkr5VfUfamWFa7UZQ9/yg+4gut5dcW
CT+FWTMOyCNv8zti/pq86/H8jRjtTr0SvjkDPIVh0XRyB7tFj9xGHKZ7ir8v
BY6SMkL+z2BM+blp4LwWsvS26cEqL8O+DidwKwy/BHYUoHcnMPOO1jZ7SwkX
GUFZzoQ49TLIIoH2RNZeO1GLKiywM1ANRLn7gveTsR14dyu4ORxEjYiO4pkR
R/DTvdlSn3W7Os5R9ODADEyT+enfJtCV/blmrb0JHfhKK4GdGvBshdIjqo9g
AV7Dwz8BBPEzm4v2oiwZt1Yz6HyXMyCyfyEiXME7nEZFxIcBjE2izs7cUnAE
HwyRQ9oVyVzkXLlDiukUEW+4mfshjzvYNPwqRq5p6mqdLcjgFLnlzMzrnwGr
2h5L0DF+hNoKDhdfeM+043ITOuRVZa8QXj/WGymY+KVhyauZsDehOd4PlDSV
XZiu/xgMfxFKveXG/GV+t8aF2GA4/VjMrPN07D8iFSQx4YTkWZYv/xtNn5NC
D4pigUkwdlqoAcV6lcpmQeTz+e7zX4TAP2YwYdYZjyAe+AL2IhA3c0/WtjWH
jG1eWggH0PNInXFr7DpVD9e8FWfknMAMBM5cDTPX5se7+YxW7ZBS/45nKSmI
gJAK6eDrSJB0iHelYKTEtLyVGhfrvLYAIi2Qzj9EbC0ofl+5KZD7kVPQ/3P3
T4qLzV8Wf8QwHrT17tE36GvEEve/6zZamubucSAeycwkt8oytkpB8qqfXpz2
b9As/r0LoMx1od/5Ys10I9AbDcE0gfOs8oPd9q0ank+7djvbfjmLWCmI6k+h
DVdPbXUWoe7KSZvtIHbKdC1FGv5+b7NIcWogy5ZaOnnhXLPLOUr88AXVN9ie
Lfx8aK5YFBRZpaU4XXs4oDaFEEoN23BE+juAYyGqaIba+d4xShmdQCsXzbbO
SpnhAtLmBqfqyOfukEhStSm8sDwBgHf8da/LtUgJ6WUmzEeG+ijmLh3mvnC5
XCWwMbCwmn3656KoTQz1ei90N4tK0aNbWtaNWew4Z5Vt261SHUDXBRePSrfj
OqeUHqM2N26Dwyh3QNVfT9GSMl4iInqlCLq/AlRaRIJOCCvmwask38YGt+41
1ngl4kQbG0PuD+PzgX8wnBWvxoU7C+hkE6YIYRLIWIDLvR7Qwpsvw8FMCehp
YNXKy3Jzi5MkrUVWgZO3OCcRfz1ujUOkQpAY5Y7zNoAYr+h71YCVfaiGrfMD
1K+iHcik3dkFhbZh8QOf7jF4zULCxTN7BXLIsFlj27mYraVtP9WsTru3IfVd
hMddAlmr0mjXuvk1Tk6kYhOxbGplk6sMJfK/AUSjvQC1Mg7IoPb2BoLmF2TF
RMRJMl843FapTbzw0O5OmLJuKG+t2SrxKUEhSRrXarj9MrAYHUfrbACpwhcz
LlhFqoasYyXKSkDvsztfjXigGbOp2idrpMvLMSC69tjT7OYgSasJuGu35IhC
BBVi9Ri0hRsxZmN5/mHmWJvPYeA/9z8nqCsbF1PsTnFt2ZiH5OS7F5t32TfK
JqkymtkQmyfCs2u97SugVYzQQhzbgcJht8R3mS6aLsiaas/X3lPlj6yZ/anI
F3Y+oaBcMinkP1PjBE5cDSN14QDsHr/nDmU+pGmDx7G3LNmtJ7lNyeAyCQR4
QnOizf/1e9BVjeRKxjgMpGFBwgzlGIaA+u6j9OkgSOzbvKYgtgcYt4HB17AA
q11WNUU+yXw3/F++8wiuOJ51OT4FUGwvu4zkjFCZrp6SrfW55SxduuzlqnMA
08m3elDM18uEuY+9I8SbLQcDy7L+CpMxldLOVqa4ELLEYaOCBpm2MZCY1pgO
eXA0K+zLx5rVIvG4rKwevinliNrxCGEHSYfCPtNQgdCBD+Lo2DeK9xME7rdB
Es4b8aifcHFWJ0XK6IPnQzvkqu35+4W91uerTkRBNhiFTuADvagEvI3JpGCZ
HkgK6uYAMoFHXGneMHtLhTScruFJNHi/VTPrznfXDf8/sRW6QTgrb0dlnenx
7/74PhZU1vRrwNB2p19PwhF3mmQNlP9CaRYDPkjUD7zeke/Ywp2/yCY0REzv
4EkScGnKE8sjkzgK4Jd895cDA7+W0thP4tPHJ9s8xrJ0FvlNTGEfPKi8InL0
3q4e0fw+vXbEFh5cSCbEVq7E32WFOKvsrKCqmLjfI1EolGGFQF8dG/5CW3tz
pbHvwxhLPEphU8a25ykimSeJExQmF1cnJRtXTeo7/tOGR12uylKmdBzi34mj
wQOundlPTO+v9m8vV/tgiS+ccwraRjzQcyhGg84CG8bUYzXQeV0x0widduov
o1l+KtqO3GZuST6ChP0fd8wSrICYAy8AoOJIUgOY8tsfVV0ZQFY1GRX+b24y
bB4bXRywogH8kJXRUwpogmdGajYA8s5vLKtwrFcO/tcYtcSHHKENO+BgAIeF
KqXcyIOF27TNngSNagbDRcmR1Fkc9eyNv1B4fP1VJ8KQ74+1Ig1hRFDCJifP
iR4DRqSPWmhmTaycaIn2fZS9o8ma72lmD+E8eKGLQVIiWK+lD3lvGmiY6Kij
dCHqa2vctqv6YdsAghF9F/phDH+0CX7DisPOBAfGIYMvd0kR3Ka5DN752Soz
zo3lAVP0A4mABJzOWz4mSu5eb7WdNcm940xIQdmdlkjOmNfc98YSVsuAUYYL
bJKTAbmGPp96qfMwhersubxFqu/FJF4bNmmqOaraJyE7tQFztItpr5QiAIRn
gDJSijrHdrYJaRCyPT02aYcaJd5HLwZqK4THFO193oDT7Pm2JKitlhIGa9Uc
xEWqhz9t2Wd87zOtZszAt2RKXvIoEIe+satDbiDUqs4G+Hmx7SSj0IaxILUj
SmHU42d3O6pmgDiTuuXHczqm8AxWkuA9TGcecgkxrW5KsBs3R7hXtCkl5fVQ
O4VIKFMqCkWa1CgKBZj+E++2lOg4+AmaZUnmbjZ1Pg+8v8N5TDIrPSMwf4N3
p6+O1WGnOIaN36jAjHuGNwltJLaWop2aQR+ld2Bl4kC6Vc1QyubOauUN7COQ
7lHqR10zpAqfGUpazlUFr1dKiJam0bzPnQY9npYSlnp1/MPm0ZekCNgWQZm5
u/QSP4AAIhDCQu+waT71bQ3KtesaeBsK9ryY0uxc8X9oOp4qzSEiMZcuzIeF
1SSnkR+RVcyHMx+9QBPu5BuFoFKsj5+LX47XieQWYZduLm0IqdQmLcmyiVb6
L2xQP/7LzWXEVwjweUFChx39UfjW29qNawADr1Ykk//SzUDlI4m3C6n9yBaA
7lknLFJGnegr3Wp0LY0oEqit1Ktdhu2iekZRVmm55P54SuSe9POxlqjN0eVK
gAvYwtlFA0p47lQoW0eYMCv+sO9PBIcuBGdwsdjPfZZRHlbFQLVWNFSfMdkg
tQjuiRdBkruReHLUVYflOu/vi90hF/SSqX3mv1TtKX7CA4+WW1LSdJ+WOaxq
E9WxT+6SmxR0mCZ3B1l+PewGL3FdkNfVmg8mk9Bnnh1+8XvkpPr6HfAAtKOq
1yTbCzPRhf1AJv0Iq1nz8rcBw4OTVbLJkvbN8cdvM7dSX6/dQ4PNLQWS0iz3
MkgC1u8BfPExPPsXupuntEPGTm86xnj0R0My83kCmfP5azU8/s1/2/tZkKYS
f6UhtIWkdMC21wptj11wOxbV0q4NdUMsylSdHXLZcoAy0i2EnepFcGNxZJ9V
gWJNb/z7SHhE5Gi+B07GPIpdKGBBkt9umPQn0E43kaxhB34cJA7OReS2W0cv
D46IKyFlrovmHnwrCE6/1MRvLeChnRENyseDWe79LoguqqaKXIyI82GRDi+q
xCe3eDC7r5K4MOX+PfIX7LfWfepubaqE+6WxnUIBgl8PG/fqJVUtiQRnt2Uv
Cljs4zDPHKHAQCnoJVefJ1gWHIdgXFI+aXaGDocic2nob+U/ZudSTPhzZG0i
m736JZv02XGZ0HsWvTFCFRFFKNkklwEh5pOCSUGVFOH/1p+eMdjpHlHjz3dl
Zt/Lg4h+X8E0zwzFWhc2Nnr/Yund3R5WBmVT5E60SU01zsj1GxML+79nzy0r
iiHxUg2wkZMf60CGRYyExnCnwfodW9WGh48x9QvPy9qHzvwUKjPec7ods/9P
6rszYRxjvRT78v+D4bmkrGVJmJPctO2xNu+zeN9Y7Ea31g5EX5PWqO8gKsNB
uSyl5HQbEHp+t2QHAYK6J/YdarYn8FNkIpg4nMpqrBV/mIOB9ixraiChFN2P
7/bcxmy61zytU25udcVuXK7hyK56Gu/Cj1B25ji/nDSSwuXgS/Kq1l99uI2K
elMRCXmADQyGSY882mPMrplPxv70uXUYEnc4DeubZh+UC+f/VLBRIyzjOhPS
Om9EBI+FKCBDgdDGZj04YqldRhCexmf4wC5TeR92v4At7sOEwNqoe97u+yoY
oAdAj0B+JRq9PO3813w9PBixwmVaI7B/OykXYTcVMXsM3GqNDlFA1VfuUWeS
0LaTvaZknUjQURa5UY61gSO5I91oz3sGW+BAscSCx6WdEfuM2MNEsjvkBSTu
/liNQPug21g0Wx7OFC1QJjlyaoT1PQ6faEyx6untHrHxSL7KFIoYOmrWGYZa
6IyG8cLBpCwgZbSydzuMqDInfzBgvv98Tr/7nm9gJCtfk/QamBRNdlY3qH3K
0o/vrN+fh8LLW3djEO4l9ul/BOWgNV/ERB1bBMKWiONgVgodhWxAfmCd9H2z
ITfJJ1bSAQIMho9OgcJh7AFYG3hBVqSIrESvIIxw5tZhlt9tuGz6uF8pCUeu
UGgpKwiE5EmVlUb51ux3dwR06qQzrfAznw46fl6K2iciAcOe3Es9Ey0qNlj2
p0srC6jJbRzJb8irhfhSie+RhrWifJ7lQ28LO6SRx20p9xxgIcUEuLS0Lq8s
ANKrauNmNDiWuoycGCksZVOVBojTxSYBrEwD/EvnmqJWfS9tm63PALMzXwbS
0cBmyKhGKtGWty+yU3I2Dhhl1nNit3pd2n0KcRitzRXjKVTT4FcQ1Wzpag/Z
e8MukzEb88m/IEXMEnGTD5UG9NF0rmjInDsjpvjskcHGZEqBZtT9sm5QCIwO
TZ18qnwvHfbLBfWJFnXgz6TJLZtkZidJUjUJk6xJYH9UueZbS+9JfZrVFVy7
Ipyw24l3LyPcpHSxwyyAzDQJU7TO63epSlCgfESVJJIwfVZ4SYruND063FKF
ZZTjIckaOfMyszB2Emm22wFYFdzY133i1MGgY1Msbpd3VijE3GSXWm8/g0qa
h0ei4UfW8DX3yRDlzjqbjIplvzHXvu9+UlIRNrH3Wm/bll5FBiPsPH2gOUbl
qykslZq5/b6tGAwtPBHmUHATltzsBmbmPQYTEbKnhf6igFAz8SvOzB8qaBaD
AQPSPf5frykL3iTr3jGwY9rJeZtNM9b7Syue7mo37fKJ9eyqFk76/EoF+uIt
Soza8IAtuGATIrSp8PXxRuAdF8mE4L5y8FXX/tYipBHGWJCBFtJ0y1ZdbBfB
pYh8K81qpwpqLsPk898WC6JfZiqaxCdcmJEXhx8VgHLgJhSW4f91fcDQ0kfT
8p8Ndr81RvqWRj2635UQSFvDeF/d+I6N0KImcbIQEzvF3sE6iwmXvWhOqsZd
XbGfqA/GmLS0Z+4BBiSb9IZRbsmsMpkFLOQwAiVKZNKrIYBtM871M5w4Zbp0
DmJdoGacekpLcsW+LRddw0bZw+yQZ7g0rfhREyUpVK5931Vx1HX0VPvnOO8A
5mxmmrFBwaCOPRtkMTR3hMBXXPyOe3H0c1SPh7cpqbbEpggbkTpvbQVJBQTk
y/EA6yK8HXRmokmuxscp5ccMXV2EgeQHsVEIe8J5CPaLE9Gyks7f6KeW0GnJ
0vC562wrreTCA5LFCMzhseXy5ViQm1QeakbBFKdlnIYAfqWnTkJmzQRE3iz6
2CMTKfgjAiTUapm81ULDMVKyOXEVxoXjW+fpKVrN0PZ4fgcHRCa2XEyzqSQT
A/v4cPV6VIvHwFGPjcR2tpM/Mx4VFFWnMUmyeUu+Xv3WpdpZi5Ufs4WPzdMV
Ka7KD+MunrQJ23DKnbqKmCwMOrMHmjI6f62VzTS5zSOmX6Hh2j3wCGG5mOnn
3xfGIIR/AfTsmN7VQzjlTVbRMgV8CJ/9QwRHZMF/fHpgU2R3jEf9IbdmnZkQ
4vPkqSWThqM7+dvFX33e2E/q8lX8FdMvuHDM6jG6K3U6LHGYKu2dDmOVhpBp
tTOJLS5hqedgLiC5dDT05Pr7IFGlw6L1PvQHN/y2PM+fxDxyRNxDzez+fCU8
B5/s4/w5MHRRPlulmjj7leV2XyFymwnfVnyXS7swK9aSSOA9hqKyJeoPcqcY
LyqWE5me0f/g5rNiXtdEdbai5lt4ECXkTBlLVuMSTAwfS9m6WntE9r6Bu4rF
cxOwbKZ65KuoQ+uTTGPXEPpiJi8alaBfE/ro+GzlMms6tdp1/r14LWsUBvhH
+7m9Iypqe+CBZTK5iFr6yEhiLqQqeWK7WqIYkF88I72vLAQYFph26dJfKi2N
lFCZ6Pm1gsTh72+njCO+pbAfFDXd4Ur1ZF12opOev1FwF6zkCaEnHhIm8vE1
xk1lI+2LFut1Gk/aVg796O3vGd2yiCevovAHYm0PUzcrXZ4I3F9fqN9DjhtA
GnayKsPz5PhRrKtpHc8gEXtsx1YNaZZiss7J63QNEjvhEss+psWVqwJCx9/i
wdglqwW8Z4tU3vmUSiozWZpmvvKm4icyhYRVR3GHT8gjay56OXZxW810p4Jr
3MVbRFD7+MBVuSzQIywmCC2BE2ADlOMbvXt2mGyDOOh5G88DHXAHv3TlmhXd
oIVFxpwyv+TIa3BUkyXQt1C5Mbm+qxMteA96ZEkINRnYWSmhtA1OZyTqiAZM
YMcL5V0Io90Ink1KAgeATDGWsKxg3Oe2LQGBALZeleM9JYfGHFuibZWymS5u
DbA7dxOscrFUdErHnPC957HRD6gmnrKzrdnlfkY2sWKmeNf6Z3sBXL3lMevH
mwtNZy7HLNBpEpaYkE3Uh+dnKmcF83641+1qJfGdF88wgVIM4ZMGKFOs0a+H
dKpfE6wdqWdaf9cUs26ruaVIkgcdlkxO3s4AOvV6h+iyHXKBlSMOKG4a8q+E
s/QuW0WDn1DYxRTkvhZruENkbWu/ZOkxOaHR78MDx/7ZjREh+/dvRA4ObGaY
lgYTJfvqo5FiCAWcsVFoV7N2cx115jLrS9fG/yuIhACqGhMfbrXLELQESgoI
xALzno1opcTOfYfJar9LLQ+rEk5Trgo5yK9UeCuubl1XR810ZhoVZ4CpI3io
r7AF+Gri624e0Pa/OkQbPFprKhQwMTz3R77VpvrUR6DCKHuCfRK6EeV/uCPG
Iu7ndVFxA19axP/07kYgHvuVIY2/n3W3wd95mB8T8GfMCYyvXW5R4lvOfUJ3
RSxg+OK/zgb895CifAR/eUdP3t17LaVQcg8cGYDGnDEWfdLcfzZ4h/Kqy20I
ig2je2OHgfT5G7nggak9kCzXhEmo4A/jG79V8x3SiTes6ls3xVUMx//NyqdI
v11ePo3/D5hzpaCYDWMyVeR+SWDUMT49db8Aq5aYOAxfGsUvUcNme7ux5XD0
saWTo82m2uO2GQbHt2rJvcNuV/RgQ7Q8hyrjh9v083AdQs4O5E7nYOn1ouUO
x0BFzpse7WEM832KCeXiNNhobbEFHwUtQz5yg5Ilq3p+GcYTjKy8/dWA/bS+
ktMTW7+um/YP+GJp0A4lsslGNZRSZLdRJc4w8MNo2w1Nip1MsqMWptwv3Omf
q12VkeHzWSLA2aNCr6rjPVuwvcy+c7Hc6xNosvErOIYMn2npm0GdEOTRM4pl
JNBGFSUBJIYbilyusFgFIO7uvgp+HpHSBCRtW0pICyKEG4QFDbs6KGtlyVJZ
ViUDUyayoRbjWKo5yE+FcLINo24ecBGcSDEYVXnMsArb0Sm4L3wZzfsb2qfl
uBhlFZJyWwZmz6PhOiDRJmNccIbvfJH1uxwN/7zBPp1+B8kjjlY7dJiKfxCC
ILFwAs0sEedZ6dZgzehwn+hpHSWEPh85oshc1JF/1WwjI4aM13YaMENcCT0t
ounklqDAUkJtcGayyne5aRBpGHH17zspDkgg7K2rSfBTqUNIWoLGC1TorvXg
+FsxDOC2KN+PBqgZvZuPMHUKadTkxf3mFOy+yFpY6rQVsRkHbeS5/lFh1XdO
mVSfkLedO4bga7EwlTvma1cb2rslHvnNcY8RpnCAXyyjPiMUhz6/I8B8oJt0
7m+rR+oTQjMCr2MF6L7FGNbiYA4b7LVeYBTkQC5hMsrv6DW1EZDJC7wcnCJ2
B6s7y9S4RBHNkRXofHlgmtx2fFZlv/omNyP9tUyIk3c632dULbv8i8jSj+gG
Lxi2DoiBgG5AIHbE4p4k2aSCWeW+WBYa5pveoMe1e8Rb1p6FoVYZyCd2cgjN
/DoDQ9hQENB1I/wgOwTNdaOOoZfpP+Ou9zLa12Lpg0k1HlaPlrIiG6kGZoH/
FNVQwEReyzf1wQk3NwAcNbVt4bSy9j8HVJFYDhnHcTy2RfAEchMqc8GudF7n
7G8QdW48GVsnfKYQ7zodWFHKPjozoZF9CuS7904qXWccYkgEs+WAIf49Ts+i
m8AUV/VNU6mHdMDABSwyBlpeHF8sUJrjvA6V7cvweYVq0vpJzEz3C4QZVrYf
V8jevEbxYULQDTh5N8ntXF4riyOTgr2UcJ9y2gxIRCAGFYxU5xGbyWA1uNSn
l5BDS8/gXy2LxFPuTR66ayveZjcgzAUok8coisp40NBM73fzpoXdMMi0TXg1
K4oQ1N/4gUSuAQLe7uIhxUfL7CK1jOWsILRVO18vnqI4gXfwQfnDDId5eUuE
TSUGvdIMdgssmSSuZWVrVNHuUg5068A/sEuC6iqh1kdH914Us9dT87gUiOtJ
JdNv/gB28bBn8Wnubi8rJIqM7QlbXVvXlJA1SD2rJonDkOr/Nmw04frd8g5M
cScYrs+Jqr3pwPUOmM1PoRg1Lq+WuDWDPZWc9KOYoTECP3zvf9jzmGGy+PU6
7PFZ4yjyTnHGFKzlAj6A4/vmgefw4RvYEeLWy2TpBqGx1svAGwClh45rAJ0/
43I731T+UccImPo8QnZu3iSDByI/7OnzMZKgweS+TJcxtYEhSrXfMC5CLVqG
mLG2S5/kkbG8fAZ51lba7RrrOAy7RhyMX3U3byrze8LKqToCQTH5eG17gZzT
D/7Tw/qg27J7v11D/tNmGWvRVo6xePTsmwdB3VzoiDYuPKmYlmrLNXH8/CMO
9mQUS4pf3OHR7SvRFSnyBsdpXi2778815h3+NDpmCq+Sxz1+oCR7TOB2f31Z
mdXlsSXlx+opRaZzutgeIbw2fC/VoDYajwE20OGvQ83aV2KCftb6fnC1zdRw
m3VNoy8IG2CapTlX+yBhDvxQKeG1rnEgHtkfmrSkcptKszz0gzIRGqckOXai
LeSWLYuRXYizATrS/uVGPmEubz8b0AfhpAlOgwTmmLG+lV5atPvyA6mKKsBg
KwT672JYcgX1m9FB1VO/H3rcxC23uF2lmOwb7I1zdz5V/AszMyTFRRLRa9aC
zuji2DjtVM0d6Z1SHVG2OT54BK/qCeulRIPbS81WKg7ZnwXV2Q8dTkcbiC6T
zQk7bkLzSh0AdJ9XETm2w0k7aJrIpxuSID7SF6k1Hlw3h+bnVfCFMZdAVDPb
YwDhZoKGl5axDrxuLsG/EOXX7V34rKn9+6t9jyQ7RAuW1xrmDuE3+3pU4sh2
X3resoSx5bZZQNzRHcEhVA+NJvGurhBeux0u4Sb0RrKw7F8FSZiD/IrM1NbG
g1vsIrO+qN6dyLghVZTjTyXQa3ZSJuHRqB1LHn8455dys36G+k37Ir9SdxM9
k/xX408JXjjveypMPA12+eBG1LD62V48RBBv9hLQYX/Jzb2Ts4/YTc15OeAj
QN5bT3m5EwmtqLIXPvlEJVjzzUlYX/EuVfXP0q6MiCZkkIbSDtxRDOdpfTdz
A1VepSkT9Ry8EIXEbCpjq9F7ENzkBfhPhF5eJQOHWR2HBurHj639E+H8hIcH
1eMgXGclffbcNzNvOqIrcyiCRlO/O0epxoNBCnGIy0kkkSRMmXfrHXNkvMMN
yqenwJvkP0lbs97I82uUTwglY1EIL2VTQM144QuvdnwopFikPrWIiOcvHGnT
4vjo1vGfKGQuLEU/Xsm7e3Lc4zdeBQerFhMa3nDEsRkFUVZkcZTuSwo0P33w
q+5jahA7bwUrBRaiydk1r/57CNd/2VoKVl02mwzGEujOoJE7M6uRGtiOaOpu
D4XKUKnsfrONSOAyxNvV4cGXeWeFQuRJ0NVVekXvZwwI36y9+JPsVzfIW2V+
Pbgt53euRb1xIfYEIjcVQECm3AjJTQsah0vIqjpdjzWOZYL8FhRac3Pt4nIG
qaeZtQ2JCR5Qd4vXA9xATpeBow7jh1F59RUwVoryQy/OnU9Sku9f5zZp/l2p
mHEToZ9Pnio6vPRlSg1HN0wZPojA5dj/ctOCU2Iay6Jpg/9zAbVhDaFODHBs
VAynNq/8ADOrGiRODIoLSd4mOsYdTHYM3SnNXpM5jPrXAZZ8ayGPgmNa8S6J
uPm4UhK4yWtYWvrke3YE86pkQLMVlIghgMXq5nOoQtKNNocx91KYS2pjshGf
zf5CFLNUJb34onX+OMiRkFggbGNnQtFTkdPquB3iulx/AmwMnRwT4v+kgxLA
4A6Sc2eYmye1H8JKIuCno/BTfmI54z7c681X8HfOXyFZ+wi/gKXSemV7oPVW
8wpc0Dm9NaLFw2KFFpiigBWqxxAZCjVNnv/iq3PeAWfczr/39/UAKgvX98yg
bfiLQmraqwj0UA/pK8s01+ZDxUHh82ENyF3a5SXMCAmrQNFxbEXyc3JenWM/
CragB4N06/NY3YhuSnT9xvLySOQCPTJmJjsYHMeOuEmHnxOVV+uPUwFUL2LT
E8Gj2cxGCC2xPONOS3rQLTBV3f7YGlozvZaH+Y+xt1M6h8SzFU7cnwKhqUcx
p25DTnZZ6cT6OfSuQ3bKDzJsVW79oedhW4wEhHoZxpDLGvI4ANKthFwEAJo2
IfhGntjsP8RGWoVB3kjvisyuhyXJLZiNcZ+hFcokny97n3bXzKor5XOye276
69ovpQ1J1ogMtWapQ3P0lxqpRtETGObCdqQ7/TKEBdPFQ0MeF8LlXIL2fuHA
CnguwIrWhS/b6siN7J6LTHJdug5VGXAwCm0sfcOgn0Tey/VllUry3JlIeIyX
cwQ43XuUlgKALayey+iOeSLofVFvlmO/CpNC9Yw/OnX7NRobidR+Tj2BCh4K
cppOcbUr9xiQKDyM+LsBAj+veOMFkzwSg5KglHxHWkJDQZnS0GlikxHZKBTU
Bn5KUC9SuMUTrar0pG7x1GvzK8ckmbLRwGS3OKHX58bnccsky0Nbo6IRDklg
DqaLbd5H6xiwpmf5Ua60z+GGekMP1NAIXbxBezVVdVeEnl9rkLCoWZPIMxUZ
H4APOPrzUoaWzBT+MCHXiZg9P27o2M6QKVdJU3AtQsIGlZxISZi4Bm9wRJIz
EO/Tkoyb7em2WYgiToS3ECVBNIpsCX9IYYiN4qp+Ck3o999gf+eB5eQUqqOc
8aF3t/qgHIgkt6OlNywvo68oMgoc5WqxvAUmtGclKFnYNSN7pPJJ/dv0aUda
O2bpYieGLH0SzPeg2rEBel4UKQ85TNl6z3FynPmh+Gz9Fz8K1xyFZ7WG6BxD
87TbdJR6Mo5qA7v4Hlo0i0vTyD5NaQVb3Yjy8aRgsnFW3sOpnKdNdkJm1VdE
KwrR3nuKoN94wXaf5AEF1RF63MQF3hGlIXTt3mLXxIwF35IPWKbRca2DV5i8
FpvznyLaOXSyREf2aZSfH5fCaE9CyV+V2WRcDtK66hYYapb2v3zslGIDZrUV
IX9k/kCikdcnCBML/45iW2AmrqXYGrrukgSnFAC4X/K+UGc9FAjKm3owrFd2
5nQ76ESoPQ1tMoU2UH8T1mq8u6OpwjMmO4AnoyowpbzEK4cEA386urDclTGj
qCwhZkOPlxYL7Z8Lhuq0CBuGomjeWHMlvZvC2mOpGxVAxvzJiYpSskoO5bcZ
LKzlB3zapODBRuUjt/srm+Uc2U6BfWg5kLD2i+Q0Oo2bO/CIFXCo5RiZDSLC
Lg9RoAGdqkC38EsBB6/Qy/IL5rx21C2ySZaMrJiFVLg4xgdzkXBoUiBxT7Nr
+MtDHJ0BKqAnK7/4jLe7kpJy0L0lt1U6Tl3Lv//leY8iBmXotxqbukj9DDwv
tv22FffCnNBXbyuVCVPtJHNYW4zW1uwlwRW094LIqwN9nEVJt3gZgU5P3lwi
mzPHKRkbX6n/LZqBMnoNwhxLzAthScI5MnCw70nTtb6NSf2+qAqzmQ1sD5Lk
KaJlm7Nz5ovE82k/SHuX1nzRY3uYXYvsmU3B4aq/9CMQohOwd8j2+C29D8jf
hIzHmHyw2n26fZ+j/HhKcINf2Yyxhduoo+whaeFT89N8+5MWUUklom3GBEB8
SJOiN+Frh8OId+FsXqPJX/JYwhLjH4zRKJZ8rRJUazcvoo3TsNKSdNCQegT+
QIFX5KwGkxbjC5lfSuXD7bpOJITOTwbn4p4AsL4GR6vpu19zhN+wcfViMLjT
EFy9GRLOxqDnlAUVqAYYUebkASTkZJLWw/ElApmUKUpIRmnTBd5Vili5pnCh
GoQUACeHy7Sde5vcNqqU/FXZH01lUdIzbI/PwCVP3MlqznT92+KDyb9UuHfA
XuizLW5NEhv+3XeZVx0p3RAIm/I15HCRqSP5dfP+AfZWZhDZhrliHPkuT/jC
RwHwAxypo8WHnZA5w/xdn2rmggTF65rDNA8tBz4Ar+9mJRwv2eckzcPMyLLo
ehPQm5nIQTvgp3qUCcSl2CNNLsQs8Fs5/QXUU8zV/4fTdV+LRQO//wRMMPR5
Qtl4fOrhegZzyb3xJkxwWHA+XWNgRataLstMu6qwDIDTjVhn3bz9dYKNxuLd
GP+iqmHafMmpJRrQmIy/uJ7aGm9Musj/LBXytJNIu8oBaIiTxd2O2aIRePTN
VkeKMtVJJ9g8SCR7+TBOZ739d22TfFvUljVw9jC0hjxM1UwIf/kQ+5uxTsJE
Yj0qXhYIyJ1/lXxkjkymUmZVkn+R0ZhlBveqtBlVoMF+NZb/ahRZ+Pl0C8p2
U0myKTChsgvy36WUr0hWYFsrjif6no1IbeLhD9vnJiTasjUQ4kfa/YCdE85e
QBtrcavAnTQKsJi83X87l3VrC52A5x34nqg+Hv3Uc09m27CqqM5ac9+0W1gy
Nk+osRZHf/nB9JNUbM/Md6Itb9JjmtDo+AnuDioOwlQkd0u0kFnunb60YZ18
TzVv6ZxZaCj5pDQGwFVantoWI07LSdyk2lWa+HnpcC10lU1KpVgySRSHR5bi
ybCKUUflskSMIVsAzdCWsGwN269dCnFNP2yuYhjDrpUInhS8PgC+Ck1r85b9
Y14vXIeaNdLPeDRaSHwJkTHbMUV+sreY50vo93T1jZawhmxoWaIEeqAfElbu
L6Wbpa1ea7Hfw6ahgCp18amHkPRR64IxpYVIKi96RtAi3uskQT0gBSSP1PFw
iVJQDK33XR97lGWHuv+pwRwtHoSc+pu9+gc4L9XYPK7zm1NaVlr4RbwIHGSc
0kWfJ7ow/nBrRuCOsSPA027s6of6ME1fI9CzaWFNa56ApAAISgFvXXUlV7RN
Hy5c5xT4dpNK7PMUnWpjm557CKQTYKbj20SWZi/kx8LdjqEG85Yrsqj3ZHGC
IfdZETu/Y3Yojr3rEMxSk0oOhXvDaSWP77Xrl0yfJQ8luarW1ZeDEbemNExY
sntId4cH+uWQpjkO7q7zwSsbObCzvWzQdMg9AZrsTOMb7/u4uGUrpyxsb0IP
tbufQfY+0GPW/+lhVOJUOh/aLltgoukBiiOPo61uzo0I94OvLdV9bTxNiC9I
A+s18NOWkZ9DM5vUZv2zEyAICIcfq06U1DmvEI2rBJf+aW/OPqvl+4Tr9m/m
+iwyXoD6EBpetCOiIOQCJqLNBbXWKOs4/FRU5aYFuW4LHVUHKeG/1zc3ATNC
WaRysZOOj8dVKvjNVo+PKU0DxB8sApV8Kh0ea76RJm7jKnJo6j26Qbye1sEZ
AMQgCp7SH75ODs5nlgnIpf+tUNFw/fVJrEiugA/SVfWEZQO7bUcQTu3zrkth
fHX1fC1daSGG/mGDzgU+usb/iFpIUESa5HjoiU+Pp40trpeRZAr9ToITy87H
48J61bf3EHwuTfX2FXB/h6tYYyHiPQb6NisKFu4SjnVo1X65GoMK44HFAri6
cOL3+06MRw1C4M/FiD28Ix7lAFI9xwITjyQqWccECOAfAb5CTRoUNIcbQ2EE
Y2BO925iqKL1A9vnHKvYPD76e8s8d2WIGCxvTZSi6mr4IKav09kElhov+J1b
Mp0pyzOUjkR6e1ijaSeooFiuui/Sp0OagKnn5wqJ2UMr8/XGSzKtAFLCfSPZ
7INwKiU+/Lxym0Mgh79u9PelkuJRLAMSdPg0OOHB2Sj+kIYCGWFSIcPZDJQp
fGgpfWx3DReG1CeH1eja42ny9nYoIOqvZefBEycCrw0xgxsoVp4ZV6YMeGMg
VReA4XYdj2K2jwfHJoxFsi+EWtdvPGSazClCUr+hblGxPsylKfwOnrcBGK2s
GuXNjXrWA6pwgGwwqcTlBMfRA80icKSRYtaebOrP5tGjdLGgXrHpuR/9v5GC
dSxu0q+nNTvCoVfF++GB25ByXYdlAhvzvWBuw+HQyyqVyhslgpktcM8QdNXl
7KlrZa/qSn93QPsDWwl9VG116Qtk+1ljBHo6BxnRJyk1RdczGCOOjXtCzeXL
W4hfTEV4n0BSC9PBMf5+e84s5B6rqyVg/QqHTS1gs7CqdJbl7hfu1LgUOJLX
Q8nFEFOoOoL25BfnQzkV8l4xHTy6Gi8bbq3JxkShUyVK7CydvTC2CqPhCPlm
Yi7OND4JvZDKZAdKTX+vwAKTrfKRXRpfHXW9Z/3NBr9JzbeONZ5kxSS7eBzg
DzLZ6BWf5dZJTP/KDwPQjJjOx8NLZ9mem0N3iOpmVQZMTtpdYgQPEZeUYKob
+mgkRa9yPbgspacQtIghyqI+rJI56h/Z5K+hNbkjfHKZClbsiFNT05oWReKG
jVDn1mGp0oqoMwxIzScdjLOGaCo90kTRJwHJ7lKP0TMAhWfqUy3odL4KEVgn
KGZBpOg/sWxhvyvIsOa6kligjFRTRGGxd3LX3RNc3dEmnfLbIZtIfRsrHGvz
bnUIWot/6/Jl9HC2S3cwxtdiY/yLrsZVXlNLiovLgZuVlfbXdzErX9yZ+WBU
aJVM82FdENMCjspAZ497ouQkKIhp3ZqmndTuHY9o7eByJzJEA1bNJNk0I0Kh
9XhWVJhHw/OOkjzVUXkt0837eGz0vdy2pTK/WkTQ/vaF7jMNGRGNfgQBH/ZE
U5DFofra2D8GM4Mf6ErAQhWkt/hEGTWUWgSpWN7GhT9iISIoWlTtO+bWwKgH
XQyRcaHuWNAhhnuY9hSkA7hzOSHqvOy+4o9J0hVRc7tHxUHXpqWfMMd4F3Wl
SQpbnZY6CX7f7N3XP3zPRSglBS2BcZeqcaAR36A5GyejvBS0RDtgJ0yy6D+l
LvJbWs1YuuTG0pEBGZqXtkD0q2FNbRA6nCaQMcTCj0pEFx9ZGPAMlaWZheTK
O9tFMvRNNapD7X3YeZQ7R3sdDs4AdMvWrB2L8iQscYbAwak66ahQMdtQGNHk
Twdo+zePPSDX381yYrp+VggdYS2cy+cynKnkGE3KetcwiOVELSyaGSt42fYW
nkYa2f8Wh3XB5Pkgmr5iLxmpdE5np75Se2jknUuqm5RFQRq/nw2WxbTgUrAX
FamS58BIfvgkQWj/FSwUbLKHHi9C5jIafYSOOW4c+LTI/gBEz7BTHHh01hDn
t7C/tRt3V7pEj9xgBooaAfr2VhjzLNzbJLpcZWMLoXES7jIjQW1xcyUONthD
cV3d+vmCiVoVhhuyqnMJsCcdKPvCKB53W86QG+e6wx2ajoYJxyBobCM0LFhK
p82taGMNH6nEgLpayFsDp/CB65a1giBH2gMDzDJiUGh7M4NhEYbPWOk/K6rN
Cd02at77P0m7h9MSD3ZHMax7tWmUO5eSfk/d4E+4CUUi++t3MdgkY77yCWzP
0rnfd0xH82VltEgj1Ak2FWlYYnstauLZZ1tYE8gJLJAOKrlgDOPezY69tCPJ
PfPfrwCdKy5rbEfiZdLgqT/Gp05g8DAukYOGec5hauwsqyYCgNtB2FPkaqQa
E1J41KTVFo79jMCg43yGSYT3pHlDojbu95gWkr8X7Y9N1pb0bgFG8cBjHue/
dq5EuA1cWU/L/Sx7eW6VnUy+Yys2/u83eIvDi77ruvBWKGm0jUflzOxyg7Rx
J+MHHbWcD9dtqxyNCPsQeozaGNK1eanXdmqAeeV9MJob8v4sv/uqYmSNRT+a
JN0MpBY3s+Kv7ZSHLBzFoKuM3o1Dob9svrTp2YgtJMJdZYRPt0No/Q5dZMX6
8KV9ehUf8PCNDL4GK4yXt5jx9JmawDb5Xm7scH4o1Ao7ay3yMFjnSSVmkNL7
9549XrqYqlJq2W51nhxRuEXRoaCSChHPeqqajYMbvovFcGI6oqrWlAecvfMj
WXP47HItLatINJt1MaFbixIw0i0YTVR+xLjDmGTw14cNEuekzzW7pV4wbRBn
C05AnW7RUkUk9FxLer1wTzuVld7qork8fQC5UUTzOU+4AvKPmU7awX0NByqV
hwmVTPf7BYQTtuJSxx1aZqURAh/2VhhI1qHuteYkN5eI+8/vV1ZyDtmcvHj/
QZGcSvRCMRC757/Vb2djNhLbfst3yJo8e6G4MYQ9mix0ZS11voQ1Cnm+UIQZ
ZxWrpPCOqovUhWygnHG5adckeHSFFk5tPoLzV1f2ns0Ps4bSdhAL6USGOG/U
mjbg3w3bwW1+8sSR9D+r3FjlwXsVpmfCCv485xF3QEZ02MtcMXYAnV3xuLiO
F2Zg7UB7oem44zMB3OKRo52bvV42TV+Ph9XPA8NCG7WIlK7D+aT8ep5+oMzR
oYL8qvSPWOyRJHlNn/QoHaNgiq3xocCoeuJuw0X04Fbn4M5LNSM7UYDemVnG
JAYGPOLhu5hgbVgthbZKzoONUS1HaeHBEGvAs14poa7LtByttIxzdC45mh7+
+PHjrpzXOqVKWTZRi2YTxXQKbjJmgqhuJSTwZItAbh5gRIZiVBEKjW4DC0td
xS4RANPytQ1gEsLmkYopiyh8wQpF7bGR0gPkblrHy8lW0PyB/Hhpk4oLyW6/
9owUEIL9rGteQjo7/KJnCcXldJEUAlsyngx7DYneAnD9Nv5QCVbL9J4znS+C
JjS2zGgWHo8/fqIsQQ9tM42QxQNpckmiQo2B5chj0y9Bg8ibG8sapLxkqUUu
2SAqNmguCQdgmqdnt2U20i7DdII/OwRlNE2Zp2ISTK8jqEO4m7TzWXrtrjJt
QW8Cjm57SMuq5Oq1bqgIVbStqgTED6Xn+FQo0CQlNX2TGhwnH1Qeqr1YjQA/
9AY29g1fxjCVAReyF5rA4JE1uKGFbxkPCdzS5jgN+oKs2Syxv9e6TeN9/oSq
j65HZmTE8MRUAENmr2uHUEUbi1NQnQ317jQIV763AmimufoyUyBWtNCgnZzU
LXlXnP/KoOno6shHVkyifADjZGbBP9nZ20zgZVoVo/TsVW7NaPF/Wj0fcw27
twJRVOj5FtZCLFdOoRpuYPrXZ9G6DHdpdPPlk/tu3sGqoWO5gCabl9Dm3i94
FYY4lHHuYfgvxHIXNaWmY8ozn3tBeLNkHFR9aWtHy5pigyhjUmy0CH/oYRGq
5TN4HSMb4sZLUcHIaHrySBohIkweC7jlqhfjJBkrwDyijM29eJwHjiLrL4SX
IPFhWfFnSfKGDt4uJBUtrrl3eSHbPzsRU/yOTMZeO66WqzB09fK4tmW01E3R
5cFxw0SAkF9zDvVqdu7iCiPL4CYlnX2ZCUqjHYn1l9KqjPaFTqx7kIHEs2Id
pCtHdVYXG68rmPDHmCnSf3+6KZYuBCeptm38PZs2oAzwe6Xtl0HGeppJs4me
y0TuTlYB5W6cpweee2MNekk+NeHzsTKon63EGgv5TUrSzwaw7VA60ps57B8t
wH95Gh1S2HMCAHR4CurPsP4S0RBr69d9/UArVI+R6R9CGpiUfnWT6bwYG8pb
CkYRlSE81E2ILHlFeZN5gvf8xHu3acx8ID8inzoM2T3/m7UU47YLBlNBP24k
xZtUYGmPLvU93PzfUIes7UpK3GACDKVzce3H2VykYxNverQmyNub5bSXTFB/
ZuwEEf1LYRNjHT3ogu6EmFAeFZiTr+rKwpujNVbSroPMb5CwxuhVl/UKgln8
31CRkfOhRRWug3+R3av2M3KnVyeVAYjuBHclw3kTGOeJyh9/fR58YoO3g8PV
jtGWb0lOuFoQkShoX+nVBYLcTizDjclZY2O+fUyjXMbNbLOTeiSaZKFft6KL
4gmUqDBT28YW9xrSqKvWPeYKPOelMTdkOgz+4eQSsZcgkAqdMD8S3KpI1hM0
+rDY12/en7djzi/oIiXrwS/wHYRNMxd/HRe32ltTmtAGSAx6pIf16hAYXywX
HEi54iMZ26qEN6pW8aC5guQ14HK88o63ZM4tns02g9yfoCNSuqq/pgOEdeEB
k/OuA2yMWTSPWNBM6izsx4NKbHZzLuMjlWwTeLMqgObjkzJrM0EGrkHkoeGq
qWf0x+/ZWfoWELEF+pOpAvGYl+oVtG0yX0X3nPNOMRJwHwbxpDgPvunOD762
aWsfj5u7hhpn5qTli/fKGvqxQqmFcSrKWrZpr0vkBWLl/8Uunv1SdDxoXGsv
Z0oeCIiAtM4f7VkCkRATQe8Ko0vz7IUHy6Gp5JcmdkF1m6MMV2skZ9wjxRJu
dNj7ICldhCjrND/OvYplBmcTdRIfjYvtD8KMXoCMpDUJyp1fJKqbaeXfJ1S3
LfQ1BRuRS0rgK0nmYXdMMH7/6YaiSTRRTlNC3UYt8NDDlmLAlkktLfWDBrmk
wAZ7tmMcLtQkMZIWoC2cyq0Qa+TQOSbQ6ThA+ARols9uCwlktdl2A+7xjkqF
OhubCu0zbpy3M+KdwcIoWSiigUH3hBTjfdkMD4MzlKT+vwasRYSeJ2xkPpY1
LS9bul9Wv15vvbeZ2I1e/olO8kPuVsELeIXuTr4Zxh++37zmXRcMFwwN4Nw9
vg0MkNRx6XYC8DMwXo3yl+pUOQ4F1kpjp8qN7N4x9ukqkDLpiLzQ3pCXweD0
1ECVZuHH9cl5Z7ppmDSodwxE7gmAV1zw7VCJXgTi2c0n4v3Pyt9GIm7fpS79
LNvj6Eeq32yx2124Su9JVUIjaeyV0CUTcYa41/FdVovyZ8srJ8n9+fsday43
B0uX9do3vZ5uJnwa+YVzVt+OyLDAezcEPdzMQmNDnrhvnFMc6R4I2wC/NXY1
YX8vIdrh+3TO3+BXDNXln+eIiSu25/pAeBXjANKcXs6Rt2KPoUK3Ca4NlSBd
oxdLRlQu8k1TlUBobSfVKyXXSqiiX+xztHt0hDhFk1oDeKlt0Q5XXKd4DfMk
vpQsagGh+GGpewy4KOFk1IoWGpn2kJvATbeRX0WV2cO0LmDzPe9l85Sx2u7A
QTcM1y5oDsrB/kZNlWu6FQpQmzpm57kXZwacM1Ls144/AYfeew7tQZhSyN8g
PqCu9UmmGyyb7zJ9MMeyyUWF+bw7gm2q7VAT22E2BKG0vP8Mt6ClSMSWUDMH
AW+prByCLUheZcqTulYO2F7M9NVK/iie/9Mo3NSysm8baHsyETmsPb6dPgYK
05ncMAT7ozWZAJf9pKKCMRF5aWeC7C9nG6yFcecXqGv6udhKhOoKjJDvDGF9
GdrpCI/QrZMbOsX0869O18l0/0DKDEfrjcAo8XMNrIYBGHZdeWa7Ks1YHGKF
PSkvFuWniaOHSt4u3QaOHFnRy7Q0EC23doISfnokVOPQ6fMtCjzq/5I7f2QM
RhWgqj5MOtA/CL2HFhhLI4984vTMqMZa5WyP7QRou5kih/UAiG2K1Ptwj8Ek
mrtziArVQV9Nxd2jXSI8JzSF5dEJQJh0/kE6rGa8AG9aVfT17FCILnA3fInA
IG48qddTlJb7lpUZ2zc//evgnDVII5kvB9TOW8haBSE6hkRc+BHKpqy2YAtM
+5yqdktpmTU+X8Jqve0VaAZDsqfHKWapw4Cf5uTIOrSKZ3hcxl9mTno2lyke
7F1e2AicutROFHttFplIoeBs+5FfGRKiuYdUOJDsHx5IUvXlpTSb01xVlPo4
3h3qMzSdoGhb16nCoohVvDREU/Xbqn9DQVmB0lfA2oAo42JFpaDCdw2rlUge
bhxuXECTcnHpxZyKTfkLsDHANe5kOrQdLRCDdObCSV5JCMtvHAsI/qds2O7n
QU8VGxy4ljJYRcUMFWa6n7o0njhBHISzv/JDf6HBsQiufJOxinEXWyGNLZ8n
cRIp+YmtVVjDoJfJkS03lZF64wK2IFyLmEYaGSpx3C7vrLbE8XjihPU4YuEt
KJGecC17rAiiDTr6YN6WGUuKY01LBT7dqjfPwjOcuylwPhpB2h18mF8r7Ige
pokq9CZhe8STkDbJhhW/cp5ddtWut4V4SQISir9ojB+E6T8hC2aaxuqsC+4n
MbbfpQ1cYP/81B2MPk20HXdANDUSDDgUBpZZEJqGhvenU778hL7rSwLLwxm6
x2a3hQGu/vKZ0AM/h9i+BFlI3Y4GkSpVtSRgBUXC0hy/YVPVS7fUMYJCtIcy
HLxF1r9A5mmP6SuJORnl1vP/gxlORX5n0YnEXsvUPFOQ40jmtc644ewqLL3z
CoJFhAZ4KOaVHM6a0XmJxfiE1TXRLkhWrfPF3aPJbc3hbNj0OWlX5u4gdjSp
VyEqry4biCkGZBnsNnLi6AxakOe3ZSTNH/75mt3FZuWWo91v7NzijfPJA0yH
QU0fcs1jxRHdfd5F8yoVfufth1ihDnvAeuT5AV0+cODPTthxiG3TGLCaJyFs
84QP1rxT3CY4lFS2vwWVh+nw9rtON8HdFDNMyN2bCFLgZPLOjZSNMYfdRD6P
7E9oWTFhbgrfeWID4wsY19g4dhGC4aJylJikNRB92AYFn6ttKWcPimziAO+U
fdbXY3avUiR+dskco89rGRNE8tnCigJoAx3UxSD13qfkyiw+emWF2vJZwxN9
GetWPGRrdAfECWEu5jwyGmIe39cj3u91EcRfAV5owncf14B7VDa1g4HaYELt
oCSaMjiAhgP0VLi8sKBfWduXdm1ZPh7GpMPUO6aAV3M+f5Dxfre9ZDOkUp34
xNLhdpGxFHOwFKFC2hMbT7MQCpytoNHEwMTCeApUAd2TcgsYRKXL/+5z9iQJ
6T3+e8nrclo86Jwk3IzzD/y9inlFciCtEXsdqWONZx6aCitu5MAJWc4ZCdHv
oLDAp7Qq8MH/5kxAf7x5AKHcTacdF7l1q/cikf1lcB9MwXV9+ncvw87JTU2n
vzKeyAsacq+9MMLDBhWo8GC50t/KDM+yCvAtYXnYp/NOB0llldrjZYi8gwJj
6e333vbK9sUSHsv9RXyqOuUrhN56gaKNAV9WSFBSebRZNSw2Hc9TEuwCOmE8
/GId6LeOghjUZP+l4Y4tomb3TTBw4jyHmcDrklFpogb/H+ArbvVFOfPd4Q5q
jXYEPE5s9B2EIeZiU0dj9DAd3+GLfGtpjqcUWYHhPldgMi4L7RrNTpQ0c/O8
IYdUe2U33hVGGQ0zh2r33eeUhVRZhAH7XszXzURyAE4zTjrp74I3YQ6fUy53
8B/1fPhBKdNTxfSee36Bf7DnSMHhAyx7APPZs074UrtZpT6sszrpCZJJY5WE
1UTFa3Jr36A+jOQKyj3fIE2wwcCe2SbCcdYj/sk9fAgb5p8T1SHiZ8DeQXH2
blfgyI9FiBvga8ZI4lU1laZHJ6w6FzafOKGwJXWYPB432f7bb48q7X8vzJjj
KoVuy0g8N50tpMUf3xe1afJxkw74Pwc9daBkKrsnF3KZTqTvx6z1f3hL9dIf
owpik48otxghq9XaeZqDhyP0TUshZZP2izIICgiUlSCm2dQIkqJ12eQVsj8w
4aJwTBtn0eayZVhZZnRSwLm8mNhzHpGFVnkdXM/9heU05lu7Ch31sApTZ+oZ
0szYEHWF4aOF9niTBa3N8qqsu+uVsKU9DmA6uRLdw4mvXkttK+04DNZPd/36
B81i4Kwb14XYycQA+x+YSUwZLdp+jbAH1TbkV/PCFLlhDuKaNanErMp44/wG
ilV+6vGTPeYEAKsWRxyT6C8E+uGtMfhktCTt4yOxKPkiX0wlhQGbK/9DcKry
UgzK9+MvLppD6zV5qlR0BAO+1ffZMECzbc6SGoj00oJAbq5KiRrBvq9h7Ygk
zBrQk7seCFmzW9tL9RDXlbXiCEpadkWHX79o6cX0sIMymobEHGodrritwQqK
9DDtrPzRF45aNwSTm+2BbUrObtLlzYUAxjNksdhKflYurB2Ut4zL07ffWNZY
mtyEJM3GVVCTIJUTbkzBdG7I75EpQ8thyC/cQchPm2eMI/ubH5TKPDuo2dK8
9b0aD0S6KZN4MvQIFJ4MaS526GpIsdTLZ1kg59G/285a7SO5+r3hsjQqxIaZ
9K4BcpNr6ZFkyO7xl4GKuqXQdnYR7m94aJ+VUPK3RibsHfKIArNxRY/G7KDB
V0yLWmoApz4mGtTQPOQWW734FuG3mLHGboAIKt8RwYjHwMt2zYuPbdHIgnp6
r2EYUAxVQ80WbLKyWl95L+ITR9I7GE9pqd1Y28H9QE1nq19CE2fO+b2nAVw8
Lu/v5vuy0EqkFIQWQrgmPyWoM09SKmOCItJ3LO7Ed8JL7yL7oaD5VPEamL7j
yT2qiKKVf/20nKzLV/1RkySlAP10Q+42Xukt5DxCj3VTGuSiTOWKl4v19ZGv
hX/i0/7ftyTyIbodrIhwxT6/MkuixFWw8xLVhGwLvnBsoe1QWEek9m6usF2y
HU0M8USL5hx/JitbSltL5wRABs5lojTess3vzUVX7C7ti4AWUVOf94ymWVft
USrcTqydgMaLLRe1SkKyWPs76tt6Qum0T681dUxqvBJ5lbL/0XGSlSBwCRP4
gWpzBvE4TGYbLzIJiKL/4uR8BwOOcfswaZXKtkYZpg6MlKLujRIfUTBPe63I
MSRu8bKChxZ85iJPuLu3yPlmriVJtN8U2seFd0LNf321AUax7tX9fwlfNXX3
fceJ7LAiWyYnSleiGXRe0v0R9NVQ/7O2clF4Fhy1xcls687UTlDBe/HLgbVJ
3RrvjVcXeZ7kV+wPI4+bUdYlYMZXNEVlN189NjGALHVJz3tqGxycnDoNPydF
GP/YH4TWwXrB8OghymSvGrnDgdPpKeewYx8o5guTXNYFdxiHX1qASffS345s
5R6s9/L7UAkvsK6/YnnccokHT/XJZHQ/Q/YnZ3B/gZguNqcbPtNhdDeqaSXd
a//NnXTGJuSm5GT5Emuw67DqqvoBTmJIeJn8DnYT3IjDHnvGs2yVwWNQBT/3
Xq6PQMsTCiaIlEXdVhBJWiqfz8rZsQzf9vuHWDSa+RIUmAVvEVRFy16GweQ0
D92qQFOjIOl3P3qhVjn7CKsrrqz5b04S6n16Xpr5WN1vAK4XvaOoEAV2RBZX
aaR121w+ZM/EYvLz5qZFEj8DrwjffCixS53Mg/u0qQxsLyLfz98pMbhPFVoR
U82poreOhRnSwA6pBW412k8Hwl7VeyuKG+Xxm0DoK3WFHZR0lWpxKdaJ80WO
ePDdQCgMd+m67VB1JX6tqRGc01YCnFR0vPc4fD5l8j71l2dhhd7IQ3FlvcNQ
JVhtBSL3e1ZsXVDxf0p9WyryXKp08TbfBgCRgJdo258sDlgTAkJEr+mm3Pca
h/qnBmDhXQPMqIkylKnRLBAIdVpUSb0KTtCR4whfJrBHGL91XLxZ8aEHUUai
Rxu4xEhDoqaZgdES/04DtYLHoTV/C+3XKtp+Ga5V38haNXWTwPc1aaU75jTb
Qzgzpgj/gxAlpm1IfmMAzs0QBF1JFNezy7phrgNU7tOE0e+MpxiFtA3wFK6W
emwJLeG4SWFjQb0upIu1IgVdwrh30CirX8CTij+MUKw/vvLpCp8+JiyfrEFv
t+DNqL7xstLOwD9XFY6aIxH2lmFmC4C1s5u0n7nzyw+0eUFlb5rzMiPhtCa5
bg/joLZ4rFsIeij/2tMojP3sFwtIWkRMwhpWKLq8Z2ypeOmRTr93OyPRVDtr
dNwMs2E3bvr6h4aJQyY/HwzLBHWwerRNNU0+i7MEPG35TqkpWvg1MLagBvJf
d+VMtDkhUwVX2myM5fWMal68DG+VIXYKS++lT7xM3s7y9I/ccdftWUtqeuLI
PvcWft5f4IiussFK5XtsuVHCHAwhsiMdXpMQKGAsYpErYRbTGnHFY3KWHwvp
IIeAWKtd+BVyY7mzGUtJiVUg2VTSulR1Arc4yAd++PkmvJjq05IQc6sEWrbH
2ZMrqvvKTQjNS9XbW+8jYomOjDvEcZfKxwbEywn9Oq7YDQpGCkU43Jgk5Tk/
BLLiwfmXdgD/84W14PU7vsWHdietqd4NhF/uhLbDIP+rYnf7LQ7YM18k1Hvv
rXaPVhjortslrYBa0VpnPz3JnIAqoHAaAEzLqR+Dtc+D0fbS7wA+C8+Wv0iK
65aDT8V91yXJ+WIGDELdLs+gALtVqMKwcAfkMw5E65nPfX18EZr40Kb1uPxr
P5ePP9NSfhQmQ/11i3G36Px3rOg/eMK2jGAYlICz08PYncIFGPgxgfOFH7y/
4v+1bsuk+kdakvokcVH0/4xzOilrWfG5T1V918WtY9dFeYQqztnq7ce8iBYQ
Ge15WM4vRZBn/1oFmif2U+HoP7SWgqCzqG2xj4PPP2q9a7ZAQFpR638DGEEa
U7d796rWG8IaVYN6P3x/pZAs5X2Wn7WQOwyIa58LRQ+KJ5za4DIkPH5CNjt4
aY++m6yPtt+Pj8yCIDljf7CX2gCVBxNy+xgGKp5Ey4iJ4+OPTVc0BRHDPYtk
LcT/vIacmPUFlYXX+T5lem91Q9i7JYdn38pw+xm5lp3VZihygAUJwmke0d2X
N+qi+/LysxjalJly4crIbMRAsTXMK2LdNXlgXL7ycHX/3DeEkJtOsQ35Z01P
kx/EaolXONRCtBDnSUi+EWlq3Ip1j/A6Kw1c3yySEG4kb8NyRK7mjCuk8yl1
9NPMH6I6bwmACCriO00HxyjyJ6kplyK93NJtkfhDoHpKPch1ON5YuQmQdtgw
Wa/QTIdTWQS0vmwPD0DFIzF5ewd7d/bjO5AeBk+szLjazCetbpE+hZfz8KSH
hgOViQ+GJ/vAXY3nRnZgRFbBzqGQG+Dom1l+eArVaSOZrOKvEady3YBCphdz
gKcaXPjpBIBCsBiBZbyODQ4p8ZhCp76dVBkBzDgAc40WHG+bxCte8r1GxWIT
8M96idXptf9DwmAfp5sEQmJASih2ezezOcvnG2C4p1rAbMelJbUYBwJg+TCx
OMXllloZC8Sy2AY0IfqpHlf1D1Ug/Kvb/rESll649UZ7lXx6Fc3H7vVId/q7
JDZxBzeIeImSPta9HLjYLW1x9l+Z8rfF9qmXDWOqSXvV09zC0YIlAd8wGa7z
k+Tq9SpXdjp5Z5cdaclAYrDKaPXu5p6ivlarZZ3q5B8mSFnbQDxgJ82vMhPj
jm6qsWGINLdD6OS+iD8KEOpdwLPXjEFduPlvhf2PTyzf/6uPErhTzMqfH4vj
D+35rGtkKP5q/x+t45zJeBwuPkgxrG94l/l+JUBcFkYvSrSJiiMo4tgnQT/8
nMZvDX0lUM8Ntpy6qD1UfmhRacK1r6Nd+n065e7kFlHY1NiSb+TW/tw1NaUu
A0/uz24YpGDCSTMvNF0FeImbU5ZIQXe0DFOgsUNkeO6rKCBj0aZ8teIPJ70e
vmbZjjjgq7EXPv9bxXUWiYunahdJLOi0q+UCTjrywIEcgrx7s6E1Fj6y12bQ
j96mkSwqNC4AYFqjXlAdtPGfhFKiFCV10pRZjQDUTTTZxiNRmHhu92PkbA0R
MTdKYQKauF+jdZ5Zf00nFGfKNXSi+Rquatgj3LwkzlBrd8CQTBBtrvtv5c5I
963iRDa7J0tlB2ut8NFB1WhIkjO2AP2wozqeyWC3KseqjY+Zhz/YudOAFAt/
iCQzs4QbIL27E+oOb741H5XY9PNxweW4U2CkO8Fzk5iuBRL13iEJAmyDUthF
IeRXOK7wQbL4+ja6FaHHsOc2gaevkwj6azyhKb0uLm8/FM3cAKoNmYjIjSU6
uNXiLNBFekkdPGCPOn1Lz3Sh4wO4TmkCCzfZmHDJX7rrukDQDi2D2a5lQSyr
H9BLtCnwcddQpW3G95XUL7Mk+XsIagODwX8OrPwXzjU4DMRb9dS8B3J8T5pg
6BtNiHzZtnnytgt005wPwGUxtIUV/G4fjrkPiKHygsBwwws7paMfrryItfZq
3rODwFHg+SuZtBdE8X5HzfvG6FtCC38V1ZeHW+AoGaKd4HJgQpi55itzYEWY
vpimkDzVelzXiOIo9DdTagnmlZ1QCFRFjTBC8oDBDH+WMQ00L75sHSTznVos
oeOf3UB/XrIJOiKPOrkCRLCP5kXWCxcuSwz2yJ8453dMXNiLizZfoTmQApyL
aZ9M9CixLVH0zXiRBMZSFvac4e/Rff8f23FINSSep3NLp40gRD1ODvHTBnKy
8/EZsnFUbGhWhLNa6/rXqAFCtGWJ6//rERkYeJ1qFrDB8yM+KBAqRb/2rpso
/Nz3i8/04+WfNS+qq6kgKHb9FLFuGUKSFlDiLpMQieHUwJt7CA874guEK7yF
uZyIPyje87KJBUJMrnURI7ihQMsiOt4zZ8JU1JCxHeKYvQPMdAv9QxC2+BFu
vnE5eGjRp37Ynbf2XuGcb1Wc3T+Qa0mLItQTt5Pr20yoDiXm5mMhs8Sff6PB
A4Ev6bk1F6hC0Ikikj81ykm9M48eJz7DB82yAuChWjyklsV3bxIvMLiJyQrn
ViLfydEsjANdViY3h1oN5UXVcgqPNu6PpNZLhp43x2/G8TC49ULlpkIZKwqg
Qdrnaw2rA+GxI1QMiBz/Lc0HVZwKBrqkdVfQLKwxyjKoubiZ5V66XQlUQYg7
PVQrKLwz/RWGPHTNUwUPuNNYmBFz+pSQk350Q/Zqjj5IPqwkpLuBuUr7XRTq
up02rwdOYdJN33Ph+dfLh4cEbUgpT8UgOdWkryIlIrWYuZzC+7HzNosGahlk
gMbFCVv/xcHS2RYEvGMaA9c1JyldIXBrDlnzlMEp5DtlAZ1Jej8tgYDJxTbG
KaW5c+JaO8lnHBBHsNzc8q0YOo375n6arzTNOl+0mp9YgCGk1Vd1nLCKu+Oi
CZmMTMcP6J7mUzsDsMHp6jT3xKPNfQWRAZ+VjM1Csrrig2YWenHtyA6ft387
MXrfTOdHWkAMg89qr80Lzxgs1cCbHIGOEjXejgQntwGIZSVzOVaOjBbz1z39
K3Snp8bTHbwIaZyHLOmrNNQiJ2doliMe87I4Btj/BnZ5wGCzyyIx2/e0r5Ra
L5cYm/8s68YSJ5fQsmnyYzwGRx3b8BKdzjLQemYYbmayzQCnODTd8s8jpGHb
mbAPgrvTr8vO/mXNIklDfkZqC4hIHSZL5hsb5tMGehPv7KLFOzabz2I2tl1D
C/u+qwU+PZy5aNpSFB1ETJz1YLGikJoDNko+8w1Uq3xVJ2gAA3DsaTnqzjFX
Nw9msu74dFXJsleDiJKtfUVGnYodLvj7PLqebKTZENV3bSs8rbkz3oRxiKUW
xSijaBRlacmujJVzVabqvNTsr87L77yA874LUypyh8rqS6mGIEn1f09purye
O8LIJIJ7LiP9Wy6k6gSvZRPlfb+Kvb5oCqdEx5gy4D3aWuk8FWcpobSS1qSy
4ixK30rfxCC5ZWMf8kot49hrT81HSSl6nqR8Sf8CzNplS4HzID6+6xe430ww
AZAq08OaAs6eCb3AqiDoQVYNpMJYa/Q6HpOxR/KQvj43NfKdheSjQijx+6Ay
fNr0cOy4xc1gxSAUADI+CEALmuZgDleM4KY2ni7AmByoMjQob9zdCRdi5rzP
gKhRG5wTvycovKsJFTIJoohcB8vXIBd0zOtZNcB4z7vVd+xVuNiW3hRJ9hKb
3gOfIYNy+SQmBboursohYeBBbilWoantyjzpVPMxZ9XfCEGgVpcwfi6/AyIZ
NWTGBADRSba8k6E4DA1L8HinyEi9GcOEGSqN1Sg02G7o04idOU+Kypfx60RA
O16hnHVMhskBNx4SHdjqwU6MTGtPi6+46reAFYCV3vCyGy+6TpO0J4EIEQ1R
iFbtMFP52nXV4u0O/M3pw/zUFxA0sZQjjCmlsltySIiGXB0fFUdHoCtcTDIa
gspm+OeFX79ds5vBR7eOojCr0UHtwmb46HcwUf6DqgVfe6a0cPMB8Ywahq5a
6psCYHwzU3OXo7H2h8+Q2gepgKtfI91JQbq46uMdqqcFAs60EJNu/v+fhv2a
g8QFJbDjCSxnsPYzKauG8xEaT/qjsq/VXo9vfJxSBOwJwp3bnvqKHDZsLJQV
cGFcw/bK2Q+v9y+c72JYCweOQlQveO1w11oPxf8VTf+K/LyFeZM/fiRG6eIn
aCZNlEsjxhfRaXsHC93heA7ATqE0kX/pNCh6K/CxpQTry/0fAIUv2hcuQytp
304ODzx0ABGAv81QHI3M9pn2gT6p1O4gUv9FtMuzeQsbvbEtk6RAfqXRndlm
E78S9iILRA7DEye7fgHr03W3ZjTlgunbNhJKZIF4/bZqVg5aibcuDuexbBlE
DK+qFkXPaL1FqLVqadZrxyM9jWtrFBP72s4p4OD1bUAqJlCeEg3Q8hlyDcUP
w/HcJx8TqvGIMmEMrnGGK772bGSopBt/LDnYyxu5fV2WxJzFdt/j7pTNBECS
eZ/iy4/U6LZVaapQYI/OKJwzCpZF23Kcj5RHySqlZ29ZeDgo0zYc4jyft3La
HBGaLSUuF5lBvbtIRIaipSmOQqQyl+KIruLj7+EbGE8t9rOiVHYDHbCMeWUG
pOPd/BEC/xvl4eugzfGIaCVXXr6iIVXCTfkN8l2Fg20r1hvuFNHeYR2Z2u1l
D7Sli/k9o9p/NSD09a2GebisUHsplnatdq9VrwgG5fyEtr0YwgnPAN2MUK4L
ju0Ov3dRJo/v6nwLdc7resfukp/X7GTcTXNnHzDrmrgAavjwXt+kNQ2dZdyx
5LF/Ie80Wg4VJRvwqgUAP72Y7YQ81229wwJxm/JqwRM3eX921LHDewoGJCzN
aWBW56SocCAzgixfuKXUuNS+pzyFWvlOd/zRFgP5G6Lw9elaCZ9H7VKFRP0L
fJCY5XQzeMzu/Q6AbDN9OKOeww5gDHY/T9gSY/HXRwIZ0wBpNy+iy+eATVi7
8EauqyHB6XuQo3vSZdKwTA+9c7t9NPKI6VdYGO2+xTvQu5nZ7Qj7lKMFpeYB
tH9JIeg3JQ3RRG/UrjMwjuwljrsqYIO+9V+1J43qTA52XlKLHlFlMg633pld
BOZ4nkssoFz2BevtlDDd7aX9gx/b0oRqxJsjXKeZ15VGpxBxTDA9+TgljFC+
LSvdtSNhSmV06pxI3e+lxPTkD0HTjI1GT04OSE+UE5gyRaeQeAFdOSh5Pgvb
gy/si7TCyRjLx7h1R3AlKd6uGvr31bKMtphSJkxDTs8/0kJvawLYGX3Wwdq3
I1yWxkGihRWdi0CkqkqGSgdBsFio0yu+H3G5tXGW0eC4cvAQ+yBMDchkxNw7
XRPtVJD9a4B1FxDh95UfCDIHeKf/36t854km3NtuRRIXG4F14B8tdodMjovL
FVw4uK2tHHrv0TgvWo5CWm0qcuwBWTZSeoWty7+vL8oAi4LXY5+lmuiCjrz1
V0v0SKaMDYE0eNThJsKM4BZnP1+feNRkGF47DwBKpF0q9G2bmjreCnI3rcBX
IQ92mwNyijgkkY29UHwlkWJ6ixVxVgYfe7Cn8bkPBYErWENRL3zrN7IegD+t
QqZ0r6KP2XoRLQxds0sydCybYp368sZINXkYmwYYrUuA2RFgfMoPvPKE+cjb
deU2pzq0QtaeaQJmReviRNYjF5zOKuV2X7+k+/c/5FZJUTYqQSsFx4prBSyo
NcXHaM7e47GIKkwk1t9f70Slc5M523meavKAG8COjkT48dJpCgDVD9WQ+OFo
YzthMhsY1UbOnJ9ZTCgVxLXcrSJeBZFImqiZJsATmjLZkWvZy9DGHCfiSccF
OBN3RTSRre0k4UE4GbnTOsAxG2swl47GZnDQSNwffDHod7KMLdVgWYa3QMl1
p5qtmiUEpxqNe2TAJq75qdl5MHwFtvegysc4IF1G8XISwMD20IWw5JGQSoqU
JI6FlDqx29/m9so9oZcoYCGxd8NTGgnNYnerKa+rMWioW3G3hecr6fV3MaLn
m3txsqFcUPs9XuZ3ehwqCp119Li5tx9DIfTCXEb4sM2ygDFswDeHB13X9LT8
91CIdMUoU+5hNN1i+0gVrYHfwdzRmIzXZeEIAKNiHKskWWxQzi6W+HGZ0SaX
e2bVVMAYurFbQJVW7viEcJea6DP914ISJ7id+e8HFsJWH4tpW2g0VAbFvrGu
dGY1GC1B8PJE8QvAG+4k7oXdkJ9Fs+Xu+2dQbEBI3zDRIbwbK/WFt+oLbVX/
E/HYxpMgT7eKLCad00wPD1lwxWOozTq2qsl1pb0hfp63LCUeA5ssbLz89NGK
kDWg/QrKHn5BnLWEc78HHtW9V6S60j9GVxpUcz5M1EIOm6og6OaDlOj82o/X
RtbWg2uOJpcbYTpHpaZFRjBZpgDn70pV96GeNnxMmq7f3Av25U5f8RmoLaJW
E654W6vXuWmMCpPcdganpKg8aSUFFq52Tp9HxFtRPxYAQaJe1yBNZvHlYOwI
WR2jQnvcFq7BuwYtdjSEHq+ah1CW6aIQVtB/nBAbtHnSkPusDC7F5d/bMtPO
axRp9QYTosZVqnYHtHco8S+RaQBPVy0S2MOXVp+EN5zXL8lcvVCfNdyas+lr
d2DdnPt8PKUBhA0SKicNStbVwhCJ7Ikgy2q0CdNpLf2n/DGDPW9DZWTosJnJ
rRK40dMxlaWCaOLNi/OliPbwXtya8ueL3J4FicI5HhX6Nl7N5OzI2O+2/i22
iMa/YK5CaSzOTEMyYYSOtVMn8QAW6pGM6+noJ3n237Vz3KG5RisOYgHLecVr
MmihNprW0Gun5rv3yAFG1wyqNmRsdRo0Et5Ra/d7st7SyoUg7r8XaF9J50iK
LQBF64oQVn+Bdh/aKSAMDRPyFyydeF+FlyJZsO+XsdLP0evFr+W5IImVPOCh
Ohesm8EhA5HNX2U7yMzr+M+IQrOnO1QhLli1qLwMN/CV65qJOMWvMKcDNmWf
FxP/Mde1l+MzUNk7lAs+DUHJqhWt8U+uTUk3rJCuFyXZq3J7gNze+zs0Q5Bp
PG8XUO/2zqUHC3MsetM19yc2ac5VzP/aCRHDkpLt4jPTwXWMiSbGkC7PE5Tf
qDV6em8jBPuBvghSwhSmyg7/PoMvzA0WgwzIgkTUfKYTAwOsEQIxsr0UIfD9
cuoAyxcCIzO4H7nPJFeWbbz82LffOaV6vkTJbynkHeWBz6ZfTzIqgpQXdkCp
LvVdomwx/M8rOs1ZCYKehN5u9BdESAf5YZPwbdOa42p4j4PxcwnVTMz3J4wo
0w1ZxtJmShARbIhpkd5hvkxPXqG95ZBYPwAwnYjWdDqsVufg8B4xkea2ELUi
6o2+gSNMSz6XEg0FMpNLkwYmB+UY+VGyVtf90tcdXAzBr6JEahYCZ0IuYTiF
ZsBxPyjiACiB6kxPLjP1na2TIuxFbnwgPjQo1eS2j8zW5WusclcPoHzJGrxo
JpPM9pChgL/WiF0odvpaK3FUkHCpWKyrkP8HklviL32w9Rf5bnfqgyxWEqst
U2OhC6/2X9OkxExKQTw3VjfRgCyek1ZEvg8rhIn0FQ2aOON8MB4SoDdYgomo
FmQOMMgEODynpRC1cE6ZIaL9tQR9uPhuDnN8IzvMQOfO8TW5lz4n1tQv2bh5
pgwpy072lPuV6Wkl1AlvZFxX3i1cw1DhJhjvb7A6igfENUtXYF3VOCd8LKuN
g6QOw/In7f5a1atkQ1i7crPOLdWGRB+wyddaZ2mMbmmsdjjML1E/ZReB64as
zHW3GXEPoUQRlKnSOAoLuoRAO2/JXWe+rLE/gf+CGz3rU8LhFJYBhMLij3zI
Z9rOhNZwCj/F8GKQqDGKJummby2lHUZTOIDe70WNTq1/zNHEu57B07h2N+I7
JbD7UhGWOrtq5k+brIsLyPCcKZFcrwhXP2wVxEv2ajUySous+hR5F6UKe8Am
8oUYvKf5nRjjEoCb9Gyzv5mW5FzlqELdMnxPm63TBiC82CDcZQNXcCGXAemL
EOUjdlB8Hlk/HMuZYoejWA9Rz5kKQU8CBQrDZ6fPFpsCihmzfsFTCY36+VXQ
XHobo6kRiQES4Er5lSwpIcHs4uQItktV7C8tHd6H0IEuW0ZnVRmnzCZKsAKr
JPI0EHglOEEqebgCkUPKs6EaFdZ2Fn+fWfPZw7dtUrfi0C2cNLutpr0mxZRy
RZNomYAgr5DIH1wZzCTa1QDMZsaX87Bg4Jzc3eOqUbcRF66Adslz2pp1y2js
cCDnNQsHPerZnLjMvB77T8ULzyTukJE/Hc8xO+f9/LCdFwDxH9KM1FgVy3w6
HN4D/KJ7sZAeDYVV4LqP4fM3vZmot6U+2iLXHolxyYtyHL5ebpXf3NyLx6K2
J3G9h66z182u+od75pWZQgYH7kkAXrgydyhc7DKqYhrB5x354rkiBDjHuy78
ApS3sCTGczu4+mPgt0aOAjoKd+Ppaa0E7IxrEUWTYCgh1MhUo1a3ij86FbLj
Dm1BtNB9VsY1wAmlMVml8G+Loh/OzX7LUACToKhyA3dBT7FOvHMncSjzOmQU
/BexJg9tG7uW7zKmUVGA/QDsawoJG57+mYL8xBPHOoz/ivqHIC7UWkx4nmLS
Q3HkSRfAOiqtxXlFduGVSadnJi31J3yTBoj/GNO2Sd+R1ybpGpyNZQ8HqoAK
DYzuXwL7CcMHcMHNAs051sgW4YN5TJIbcdLilxtB9YJpLXJ4v3jfTihwemPM
mxr/6/tiShLbqZx+AMlNLQdwKcaGp6EwPg5Biy6mGWC5d2M4Y54KwIZ+IZjn
YCHpGXSLHbTEMKrFJ9YpVy/6fOLacApepLFAuDw8Y/2FI30av2pNuH42gAxU
TXaieedn6bX/nzY2BAu2lioPF1eoZIY4JoAMDzx4TRbck5gYW8GR4Yv1sH2H
V3zPdnv5hM3G09kf7KJ0v8NtwzF7EgljyIwpFl+nkVEAXuWMuihfbpro3EMO
744ci4jxMoGdyFz5fcyvicykE2ZBEhboRQhSNDd/e4D7PMsndnvJgBKevY13
cJpylQHcN7VxVenCi5PHWMx3dX7r1B5pVK3swcG9h1JhbqlmEU75pO1bdYeH
Tso79fvj4Bd+AQhbEJwzJw3Yvl0tNV1HEbfMlnTSZJnT327DlNAnkbbzbUC6
n1bP6Dg908HUFf/kZCwV+m8A/8AQhDxRzyv7hhZ37OWFR8+H+/tY+pqkePrs
z0tMeqL91NwmBUNiTz+NcZO3kOFBL/v2aF/aVeDKKWxU8Ng4l4D7Hb8Ugiai
TxWApBhmFpW4Jz18Y/tZ8n6S0aDKYRXgO6+UN0ZGY33nQDfsn4EkD5EQNt3n
egsEt1X+TFFgSBoRWxzkIjSMPRVNWqOGKmMrSyN0Yaf8a+h87V/3FgfunIBs
sCv4nmUdzZiJlOc7vGiP82hiavltn5wN/ciiIxuQxmOE0ZrOV+15jdN60Sii
7MGqj587eftjTEZmvBc1Bn4NrCfNkcp/iQYw6HCL6Pt9gfJ4QY/XQkZ3Se5b
nSDrarFvO8VV3z0T+clM7qSz9BkViokatMHVyKdc3+Xzg+9g39B83BDAGlSN
6Ih1OveYMY2/N5FmJpDM1oB9hOZ+cH9rzPob6w9CeSjf3xR//oMRozdOKJik
hVKSadVLSkwdHdRepzJScT+fwIXGnWBpz+EZKfih89q9NShxFoHo1Xo82xj/
IXbQc+2Y+R+HUySDRLsmT/Cf5NcdZ4I2bMxESMO2KaV8cz7/4SXwvqI8GFHe
m/waGsWQTF3A6jLEuB7DXh0yw15WJpyQSaPUZlew2zXQhfHbDJDmdGRTZ4+T
gKn6eIbFM+lKWAwYVEAdaa8kq29oQfl11BubeJYl3h6N3PtFg24EeIfUg+r7
APMMpOLsM2udCAphAnX0L+2htrSBWqvgM3SXjtcGJ76Dg9m743WccK+UOd7E
iMsLZhhWKus9m9FtXSccf22iUwx88ptdR6uyjcCNf3VXLO/7o0uusqLW6Ucu
NzWv8+Abf85nsWHh61MU9b34174JIU8p2nJBXiV1DR2aTKUYuIOlc3p2tqBq
yFuhAF4dFStt+HQTU4G7UqXzj30AZ0q3nGsYMMT1L19i0qhF6458GFoc0KLQ
N9Q80q5C8KCuw4mDrq+dPa0EspZCH0TjR6AlTuSJvcW28fWYKXMF2Zqjqduz
UaDpYJsbDfkvlQ+qIxYmar1FoxAXsKiAWaR/TsWO4qAUsWdn2GF/AcSRKyuh
oeb3f/4M3io2yCRxuvZAE03F7SQFkbYj/RhGewiVCTL1BtOIxtzj0DOz1sOJ
JCU1IpBcizYUliwyBBxo0KriLuHJ7/9syi4PFqjBCYgNxWzJc3h6j0pQZqlo
g7vdCdL7wnUpfOrNkjkmBkSC60VhIMbYOQgY2Jboq9L/DZa0WhhTTNMG3aUI
p8I6rsTSUlTkTK/DyPRKSkp/hAbnJRR1um0T5tibRAg3cx9TEsU5+xV2NR+7
0WuYY+ZOH88bw7BVSCLwnuDL9bOWME/qauadHHtJ6ujFKZw+0ptc3PBjEOyK
yQTRoa3su4rEqd0YFcZ7Ih0+8FvGGrsJy5DNnmJOzJt+0eUhS3+Qgb8fzr6i
U6/8vQMi5vW+4kufjVoJ66RgHk1dZMbVAJhAriUI1XtLkegNypc6Oi9GxqTu
VYv9CRrrVtDaDCw3Jj7MTFv2dmfXzXVmy7pgH5lNLIG+Hjm3Z9OtdZnIgwMw
oPGzleiy5bswESuDwpUqLjDX4n8b010E9jcWGs8voEMhXb3t4pz0Pow15UO1
qgr810izVVsHMwnJ38QVykxP0cHtMnnLymVivoy5f1EFngcE4Sl1+YRz4/qD
MnYXpLp/XMZTEIjwM72qUy/xv0nGbvf4Uau6cvFBZ9cXahwaIW1aCV8BaD2F
pW22oyryVlBArZ2EtAhh6aHSBQQBWpqWIYIab2ekq5n8ru9F+x9g0627e848
mkZ2fMrPDk6OrU2Kx27nselg9qa189I7DaWAxSJE0V7wBdNReSVmf2gH0oLm
1dmTspG8y6TEH69/q+25q+xZGtl7ZDV+Cwr5RJI5ft5+n8507c4S72aJ2cI9
LOsVs+Q8ItK2m4J5FZzlU+mqRTc5YMTBFJjo54tmn6P2TQLTLJUhwrngxsSw
tweZ58iUkvd517+Io5JfWWtE0ll/EjwsPyp8/zVPyfPg8+TxwihOomIOU+5W
Ue5RWnqnKvHpaFQaoMrlPCDnkZ+Jw/t2cV5AqirYtFYCN+5J02kjDI7g7ivC
Y6MlmlpTQt+ebBmrCQj241etnuxsrzwo+8hnG87BfHKEnN3n2rgxL1IeNCpj
lvF/H1UcxgylJhqTckdLiZc9eWhxHT015vcAALq4d7zeBncSJRTFtYcUH0l1
j0+T9d1KuTBIxUsZRzwrbmOMsgjTbj6KiN76i9luS9rdRfioJfjwH9LqZKUf
8iDmV5SrSN1NoIVI7h36GbqNcuPa0606sS+Q4+jv6GBz4up7yn3kRu3PaEFN
a+Rys0ezhHDmZ+B6k3hNkh/wCKI8Am/LvZSoCNY4PW+DaozFYAOB7YDkVkU1
BhTTbnDjH28dx7geUNTloKEt4Y9g8iz81+X9qHWHtgqmXhZdMkhuM6/gAabP
WqfYLMAgNcVWfDdt3MtYMOEIRWZH4V0ydotMgPxxDCGu5B2Huu/NhlqaBaox
+lF7EhEHROl2Pe/0v154f2IhQF4JH/HnBLNmEy010uLfEAXrPJReG2IDFGbf
PFeuBww701JGcI9Mz+DmxhdPBCi/QVEOpedBNbPmJ8qZ0muM+xwgt0lXFYCm
RkXNqTwWk41RDdqG8N4KUZxXLwwwVuwD8tKcOC7btoDTzyI/QzB92zwYn35n
z+9SDWVpCngffJPUIG0RGcMvQGxlF3aG6bKgt8jcpUot3OKyaQ+VkVWD0j+T
T/QcwETp/QXGfFTOhSWy5H5qlhqfO/4cpanXYY6eZ7o0ThPMSilbE/9Apu/y
ASS2GaXPRHvrLz6OOXc7+6JwcHiO6XGfO/Lfc0qAq9Tut9GHM7SMmoeus8Pz
I88xIny2+ImFoOmqWtKTHobJRRYSuE5ZQMbCmCnTRvZdH7NFGz+RD8aS0iH5
Oz4LtESJgeMmvBY+BcJzGv9Pqmc3asMrOFPXYZvCJtpARSto/zpXNBdrtVG2
e1W6rq+tKEJ9CSwi01Lp3eAeGELYqCBTjVUerXJTEuLNkop5tsGbuGiamK2w
ZWz9hVSXSxxDSGq8Vs62WnXwKkXa1ivglg8kcs7tfJMyHrJBhAaHoGSlKHYP
bsGGV9QxFg5u+e3T/VIIFnNjbUlioHJyH31SD4JWRg3uD5Go4vXQG6nBck4k
iDZlAo0znHgwEAkX5Mtsva6h+F/Po077FvAF0A/zh4HadoYeL5U3uwEstvRm
vosuO+16lwOFyJpC9rg3KNlgGIN/yZBhq2jwRfEn4b4Ds+1mX+xqOHmTiBJg
GADzG/u1F4XjnFNhp1M4uV5t/6lIKwzr2QxxDQKHXUPdyb4U2WIOvQEPv35o
1lwrq2+wSKD6t5k6+eyTyxDfWJYgGtY+DjQb7Na5LRxMfg+cY1BQeFJdNTHl
L82JzOcMjO19F7Uogr5Vqw2sNGb4gG8FHTAXsVBX+KLuBSx02Epwol/Knnoj
zDCjkahVIw3k2H4fdyAfbnx8rxNh7c5hQXkHmZCOCKBSRFSkf54jQ7L/TWbn
ZzQ+3xe9z91/mhhbalf0WIFPqtwRpFHLQxb0c3EXRFCUByUz+F7NSLCy6NC0
r7eC+vulj+RUoVZLHSFTM/H7U81PdOESkpI1QH8Eb+7NZTCfXNGrb+F1U5zx
TY723mrYVpZyT5FEYowhkOknwmQpw+5EaSToolaXotxczzGW940i9fT+rlNf
aVXuucO3iT6W+Tddep6n4jKnJnmKXCEqssUWw1PdIT2SE3OJbHiiX2aHqsWq
zcZS6oqT9ILxhcXd/j8vWk2CLwL/IL9uJKFInkd2+LERerq/m36kaFBdzZUa
utZZnWy4i5lgc4iVxsz8CPGZy+6EL2Kei9+1mWPXUiRcIR6RQ37h961dNXi3
rSGwZZTO1asnB6mmf/0hU+HavCylQGNFptMFqzJZvy/RSJHddkauEiHEQyR5
P5DjUWkTvDo6lUF4Xi+BCTpOLKSScvl0OXLFLZipMGJHGsUUEvicP/pj8NtL
+xnMBYWxkkTAFR92wlomAzVHQoe+DCsA03YTmt/nDtEb/N8OOqm+BrYq+lp9
rvOiwtqaN+ZyF7qaYlT3yPkKJHuvGzhpuLURq94ezjImCOUPPUpz14aAKPIN
JPG9lo2LelxdLCbPeQWBeyVvVPwtZK9qv4jqfSvi+ooxEoXTVuyTsYBkS8BI
1v3czxSFgnIWHDlJvBBBT4LuIuGPdljH8SA5p4JQpr3s6jLl5/IJAh75Ulfr
tlmu6GDymX6iQBCGReZ3lINOyg7iLfigdv3AoPB/evnr0jdTnDkSCniHbmmy
373BiyXWjFrJ/OyedPAPpfJEtp+7/LI1Z1z5jS8FR5Xxh+zh/bvXFmUey6u/
5P+TNSZwkqAVpbFOuGfUTHLWrL4bbisIRNvnNIQhaIuBYGhGvYbfdlrg1pkN
JpE6qJgfe/oMwDZNs+wRRmUv5b92RR3k0b1b9NWbnVec7o2BhoWEbzw7wC3A
hp3rodzbQ950KAq6GTaMIjVDz40o4Hg2aulzqh0CbZsHQlmKV8wXkNBp8P/c
1ve2/7w2nyB0YIo/Ekmn/PvNOebiOG7ADmDkZ3PWznxTN994CWWdKyu4fdRT
EyhR10rot3QCF8majU8/pYm+W03gClVL48tv8cpsZLmGxV5vxyH0Pekmy1WC
KB7B+i5YmmSizgm6HnMUnS6+6CKzhQnONFCLIzQWf58zDVVMBPokVfrvBWr0
d/A3sC+H1JyJCShqYIhZATIOlBlqZzvfiqn55NjSB9GeTk3co/qW9lDMMmn7
3pqxiDTdRr1iAtLmWwI/E7WCWRwwji6ybth64Zsv7TmSXLW/lQf+LUcdg5f0
3u50nq2nkryvXWq5PQnAsf4919PpsuyKEDvfpCrrCjNT7j6qcprK6/ITIGRt
MB6z4CNx0Z/CBx4LdwTh2N7ipQ/qPllfSpvKBFwouPjzf7Qar0fQ+gUwRs0J
SWzmuwGzqbrLYNgoOzcnVeZLHAfjSy/iVlZk57ECoF5NXKb+XMcnX5mhaW70
v+XW6H+3FdKIAHtsI15XsdvwzxZXkMq2cdO+2uKRQwaWGoGHO2oDtusWy4Yd
/0U/vTimE0SV+UvVbwLntDgbK0/5JVNkwhdA0zEh2owDyCvLXNa14DCGVn2Q
8yhFNPA7zGZ4rpQauYomhaPXXMKyWqYIFaz6YzG8uVXwIxvunjvV2vtYFS6W
sj2ENZbyKvRao5yasNF+JeM1zMIWs1g9qnteiIUtlzZ9ZQXui6j0HBVZ5d2O
E4GnEoJY+bp8fTT3OFJLiCMSX8TAj+rWoqkrMWzAOd4TjurVKfh2e90qx+HT
+o/F7sAwVUKq7UbixEgWkMRAX1DL983jb35qWoptUzSZXZJmcgYEIFZyfGnL
IfqA+73p41os+2orpXHOUGEU/57jn8qc2FZSOtm9GvVcPXq6sMOAaAsMx0OF
7kZLAbyPsxNuoS6q8zMhjkYECyubmHUTVAc1H4iYN/PnLo8tS9+v/enw7EWc
BJnQO3+lPz8raHeaheX93QC6MC03FhFoh7dJnuslIAcA1OCZYDcBK3cnUQgK
p1I3oWBTl7t4rBUU/kaFeVdHoH48poT2u2/y1n6wXVMfdSrLuBXLpHlqzQEY
r1OoD9E8c6eee4AGZ/MdYZRYcWlLCpJLug77SF4mUoO2I2WvlaIcjWJpZ5J1
wuYiir2YSVhXUElXH2r66a3hhGt4cZuIeB1v8W6AhYzTzVTpRJO5IXiRXORm
UbY8i558gK5ObX8MeljwS6ArhXcNPDKn1GxLiTTNl+EPccCSPd63uqiOtWbi
uPUxCMZgsTss3FVfncjXu35RKMiYrjnTf40Ky+xvJKRhE06j5/v47vovhkl4
M6AUk7OmjrNV88KiLBA/bzrqbRS4CEzqFnQJmcS9tdb6ohbnfRIZGnD5HexO
J63WarinmmUQUTm27LgclPcbwE2/YWblANrwCDBoQLlFrSyGzcDhc4d+gCjW
nbl2maN/PBJFUfWkZJFpvzZ+kmTIbyOU8tQBsFU43gYpEzrLkKCeeHOqs4c3
jolRAEbpsZHCnE5tXh9NaUIgMtzu+FOoptVbIM8WrorILxy3/piIiR0e5LGv
0I4KDgVdIXAiZ4ceEDeZp+gf/kjtkKM/ED0Dts3+irfe7a7NY+MLUW68f5IQ
bOdT2J6x5cuds5bnNYo2kEUHCRlSn28XGFYlIJkPdahSqDdGpQc1wupw1tcA
YpBwUUmTH65bGH0kG3Bij0f3ehIQu1dXa2X4zT60SdvyfJRZ1+CCH/o9ZGRP
gtwg8DwQ3D5yBwmtJV1WJcq5qOmvtXQNhsTFFqH7VjQQa2Tx81dULMLcBlo/
OuuDVItyy5XDNLr/4kSnntvReWCpLheA1w6+gf1M7rzAQg6/KW9FjzM3UPPW
Bw9y6vI59nOdI/sbvHvaXDDKw2EYHP8hCf6P0NODCB/84DWExbf9/W+s+3Tg
KiO9zcz5l0p87cekUhI8+3m5NlVk9al19sIRPVrGzDsybcMcdIlWmQoIaauJ
+rl/mDMdhq6iNN612D75O1uMuxPidM5SuZ/gljNHg5ZyqTz83FsWPWPAgEvZ
+IiihAl3XCgyJ4VIjje0dhwjv5hnhxtI74PU1wPiqyKzOfgT3JthqTCpVnqS
O/eff/DCqYxl2UouIDYicnp/5TK+tR04zqzrM5mjHrhEtf0FCOhK7XIe+bMm
ZGpL5lD9uRZ+c5remv+9iMZcBRk0RupvJRN1LZYJrH8J+Bc1DNqoLtVbhzQE
+GvfTwK5t5hPVRQKgaIkubpS2+t2XFyCsbaLaSrfZk7OHlHfVAEAoWlhs6Mt
LXTMDMNRg5NiGI8ANTvpF5icdzzcG8L/FP5MPoGd5A3AR+K+PjFwjSJHNBYl
w/uR+NZKLT1fOdek8UwfPgWvl7b+3GXTW7ng4uV3l+m4KrQxfanXBOYGylLM
LJFntC2CxcmD8dxJaKAZmmzJrthvZ8ezY/9I9Rt/NDyjEXi1VSPYNIX5dR5p
4oP8TYaCgesburcpUhqPhjKyifj4UxbF74uqYiGuIA2c3z4ioT/m8LNXfRJT
e7wRUo0giNl6L//MTFSrLvyOzxSmHdjf3IzWDmRSsHzV2tX5p291MR2PBryM
IcTEfLxqNIsF7wIICgSLgQhSv2+tsF3J5BRE+QFU3wRyZw1L3E8apgHgwFC8
1UGM8wykRI2kDAxV69DVM0vTnbXYxZoa5hbzAP4QRARs3/qoS/44lCs8AR3o
A6vyPQ5M4h2sMp+Uj45uWVVYpezct3VFXAmmI2KGiJaLGaSI0jTTYyEOh03b
rGfvNne5X2wwGvS3GSYYXpa+rlS4C9/sk/fYSLaHJCHRcyw0rCF8rC2poZKM
d+j4rm63eSTdHi6kjTGCNPhMrDVu3NulwOWfkIemFM4220V/xlKeDPWPhSgs
dGPzxOliN1BhDzQTCj09KKBcYNnzGnIPXzfdSxcvhewhVKrKxiB7oZ/yIBXf
tu7EvUPf8jkDjTnQiCkvO+KXDTsMeL4O2CHq8AGpO8bPQCbrUe6uKMr3QJ56
MQNT/z47FWJvnN2EMTdvGIstCfx5syXZ/O7i2POHJr4M1b2e0vB8iPWBKnw/
JcIyzmE/X4KmqvFb+GIdNnW4SPkVO6peoQKXsBBwkrP5M/PjWjMHWqn6FqQW
77rp4A0cudzwnr72Q4oroeKh/D5/gsiWTDTfd/4+4+ELo7kLLepHcclapo5h
ZrPmDMU3hNADdq1TEIu9q1260popjoMu8CMLjdRptFIVxXbSWrZV6d/vkiMC
t4vhnfpE5AVcJhhoBah1GiP1p+SAZkIFf5U4xbahd+5juXDBN0Io9VnzuqwY
1zexACHr4AdrhEajNDntesXNjMa9ankt6iFi3v1uLoRnNaNgmNyWziV8MHWo
pXbzWoKGTEhwvQjWtV2fWHfND2nTbOqKj0X1B5WGkwBrbl9AhokBzcQSi9ul
jPHHYx01DnHpgvqnW7w7LZ11UO8swsJcKJU27kPFFMSfIpkEFV9infeunTed
c2gmTLm5dpZrR7510a2JmOtrQeffUHJJo5VeupbQi1s8yL3pZHp/0qPp79ad
GSIz4T9Qb1wQDHAJkezMvbRyUzsu14rMzrWlDuvINSYc0zD/scrGD46Ggg7t
cIn8Yk4NJs+AlqBvrypEIg9qNjk5azemDueoGVHOxksGAogZ+xAg9Ab8bO1M
VqpjomvNYlrUrt06WrO5lyck9MH+bJ9ZToinmgOTjuDCLyx8255aVIHmhpg8
pGXP8PsZdnIBrURHt1yy+y66z5W2RnkOKuND98xMkwkxW3FfEIccVI2OSzpA
VxdYhJaEcPfm6x2W6ezRGxtRj2adCCoo9DWFV+2Bk55Ttte7MJRB8PmEpA9f
1yXIlOeF/JmLmR7sN3x/kgJDWAiFG1zSokK8WCTdptNr4mn/on4ZnwJpx46B
ivXxklRzEMTL4vKLGBlC+opIPxkIhBXttDY2NVlaHjTIffu3toSlClFcg0Bq
JyxceqTpFBsg6Q2BqcE8T8HVcFC+dDEBoUHfih0dmSCLvJ8QVIYSNIjlpkIL
vNcmdZ7GJUesrSR0Hd6G6RXbtwqRRNZ/AVC6jWcIIvc2ma8hlXB0C90QBhL3
CVNSxRtr3sSXo26TBHfO9XJcIduP1t5NPAg0Ndlpo2HKYH29vxaPgrw/DIFT
ci6ukYgWP8bsSGXhikY6Oz6cgIfHGDjL0AOiWNrW1l0D0xCwk4T+m9xZnCRt
26d//eZhLL0TJ2MQIpMUm55qQks+2DCe+FX7b2ZTTy7CBrp0sVplrv7XiyhJ
cA4Ho+mtGn9hgzqF5BSFp9/29JgGhKZ3cJ8cmpsAlZz43TaA26VPH+JiKac2
+dBidZp7NFtAPOEtrlrvsDBo2xnybZJG9YO/VoWdaMFUWRPVTdcVgcT4hT14
t1nlgCIiMLSiiU1euBtOAFLqG0OGEJTX+rzPMA5J6BzdBD3uSjAR38QsFCKS
lMtxgiElktg0NqbE81FXdOxb/LnyHBYQWDcrkfkA4EmeTpu7Z/j4xeU+dMNe
n4b28vWRyYputFCOT/yT7JLsjwrj8aHloCGjRLMhG4kKO2EioLQKhSjQTkF1
SXRIGJSqAlc5WxcZAobLEYnnsZqpA5jZNnq3Nl96xB5B5TiaSFJ0fnomJmqo
d0Q2/uwx4s8BzXTnXBQaBpFpFLEjbll0dj4/A7PId69dUXgCiEzWJaT9OUaM
Ej7glhxDUGMfTbd9OQDe/lN5zaK1H8j+FpIKPptQC+YxA406aUbiHHrwsj0+
ZK8t7sqdyvOZzh39NGcJW3qN3BN9CUMHrf9VGq5i0bk+vA2GrrbKsS/r7ccz
j+1O49QL7kYVXIFJrz8MVVhjz/EdN4gjFQV9LdHyPJHDzf11MB6Sl+GBe/4a
4aJ/qU8TyYyaLfROXSULHPadA/Vc7fp0DXYnU6j2iWkEbiqSy/HP4YVAiQpA
OZZWFnRfIWSV2CSs0DhwWI0zpa5Q1QO0BnYZF1nQOURahtexmHgq11Ob5Ubi
EnsRQC6gNkONvbkd0KhHjeY+0TEFOD0DDd0YlJUj1GeNrdcT7G/4QXdRHIqB
UirFZwKAdpRNIDPkeyS5vHX6jRVdJZis4cSnkelPg6x4oSMPGQTQKkas6LpU
NyFQVxUB8/VOrMOtTd0GFjF8AMY2P5zzyOqJY0cRWgImDIy9hPv5MB9pCB13
Jzky+QVbigkxxe7jLM1Ew29fXCMqtiBm/9ZoJKZKB0nN/CuHtfGEKi3oSen1
KO6xf2/+Pj8Z1tRyAAuFLGJoOSiylSLyuAAsPVIoqMw1YPn77xywDhaOrWuQ
M9TiwkOLL7x5AD6ay5Joc2Sb7BkZTjfpg7k0oT3NUpi749hAYSHdPYsyfGN8
envn+UVwoBPXVdeGASPfkpBzi8ngj79VHXRF4Ho8XE29ckxXfOifDSSk9L55
nV8QXQf7BT9dTHtbXbvgRgWl7o0AHx4gMx8+2RMbAxBSVaG7PQqwlGojzIrj
D+X9m+mRaAd7c5FV58afUZbVC+Qein3VFsjShm+DGuwar3jXjNpLBvW8JJu/
6w8GO4u0Vxsbb4Rf6x1n8UH4eHpwuaTLYmsNDbLoAPk7kCNe7A9b1+CmK8Zp
9Lagp+bX4Dug+5cSNtsRsZHlccSoHhYlTpkRnWiIGMsY3oBwxF/ezzYf5Z5S
54Ia10xabaqGIPX0p0PbcP9TwhJ+RbC0g0IUR+H6gSUh3n9OGg+CKNx3l7FI
j5Ut0xeUqEJpx/EAPV1yewbgx7w+Jc6/Nxgw0+nC1PP8+fBMHokGPOYnZDye
nqnSMPDvxQeGcBNyp8gQvwGQ4omNUjuY9teA0/XKdu/XJmkmQnBWcl9KRCn1
n+EfsHSUeKk16ijUsFC2gEqoIyP3lBN1BLhOPoY+QjSnszf02B21UTBnbqmw
x4EjNrXY/2aXlhHRS8YbbvlZZ47ntaAOyf5x9Ij5ONc95ACAxJkVBj1aYbs8
APzstX0+H/Ckrlf45bWu1WAdIjj1B5xw1rIMIJyFDARxCYUBv9F/EPpowiC2
weXrqgeKarRkzZcZ4Gzaw8iTpgMHj3xYcPg3FgOPvYagSFbhL8R3AgdWQ6M+
f5vVDdu1wHQ4TJCbXk0YpSHseqR3aXyhDhYoLZAWJ767jNZY7sT/JlsGMhzZ
bD+FKOI+va8IKlsed7c75q4R2EH9lwnuayFJJZKE3xp2R0srRa5iI6uW4Rte
FF4EOr+Pzb0alkt7y99fm5PlaXmYWVDsPXWxniwO1Pnc4viQ9Csc1bPvklE1
CAWmsCw7OvBbJtau9Juo+sn+CIy3627qRcgencEBji/n8JEkbqbsgLXSwMh/
nCZMIj/TdCCpyqh+NPQtF3HgsX25JnJQl4zwVh+xP4LCncSGea4ef0QzQsTf
0wAsvK9DvaKsaPTce3bnP8dk8axjcD7Q+8x7nixMcFy68w9hspmoxY45FCxQ
PB4UBp/uLPg15ZRCt0Ub3+5FN+TuIKRuxw0e5hecfKJJe7BDr2uJ+CCQfF5f
LmM88jnuLCK3CrxbsbXBmcCe1ZVULA3a7hOkNDgF6vnWyMuQB0FDuhCdzBZG
Y0X5HOCCa8swiDRYV8YTu8VY0cDLXiOXFqf07NHiwtqeYFALeRX58oJ1aRcy
0u4rhVkD2xXJIZ6ohF0rd0bX4VVVJDE+lvPCkR9TIJFlxGFIbxFquxVmgRYG
G/H1vL48QtEbwFeMGmwC9ji0Q4/azWdU0oWEgHVqKVOv2v4ESnO2aTNZCYpe
waXsnttY4nvcGyh6awopDAcrA2nty0FRJb83qwun9vfvvltT8D5XPPHu2STV
EJbmYuDA//l9sl4uo3fAFywZOYyQkeSgdPn/68K5NvCYhJEqHyrCE5BfwXiP
4ktuMrAvln5bgxTXhEAvUMA20UvZ8LIMHFDEpQGH5WfLc5jo/gexRUYJby0o
T9/tKI6R/Ux+9j0ES3wYXq+DhkUF99Ma/vS9tnKWamMNIzJtFIPsWQFHNpuO
qkHLV4Cdb39T6EntRE9fnMkVLOENsp+7BF9A3xdM/Qgccimo1Ey8Oh2D7ngb
AnuiuDsizOFy30nFiFhh/DU9Vi01QfoxYVwEUxWIolvB69PyoBJfyoL1XGx3
7AIgAJo/ORIaKYUhiqxOhbOdxeUBWy79db7TKHTC/so5As1MPndioWHOvBw3
ZPJOrmESmQ9yE5tM31yjFN8uR9Xfv/6Jyx2JsKy8uotwLjEXr34gXFBm68B6
FlcVOYt9iTNir4zG7CoU81Oo/9XMuqMgCZYQeUVrBLXvevbVdL8OHWk9rluV
UYRowN8L1eME2NFc5lrZeEN/0ysOy8RkOfvqBr+sS+G5miaWnAr7ICtkM1uF
syiZlUsfj5Yco1FsZ4iA8Fva4HpYSGRURgQzGcT9umPvdPJy1Af6mwEUifAM
zHDClgda+yFIJJdISHfOq/ILxFo37HEe3sginL6qQiPuvV/ueDQe1Jzcwyox
XxwCnWJ5YvYUH2w+TXSU7uwv2aPJbDQwyQpY64ktDCGlnA5veF0WAh9En8S+
zPpiSdMmIL196259fLLNX9gUiQHpHZ8zFvE354JZuI8R/A+mwIZzAZoPzf/P
LWRdGJea7DhHtiZM9ozvw5v1CQoVTaEO+LuT2dZeVfalkBAthgXR4TBtyMJ/
wi2NxCvWtWAaG/Kq3b37+7n8T35aWnGyqdouMdAqK/matUKkMSYDTkhkjbD5
I3FKQNYuHFobCgraCFrpBM0axtNAy0AtqCl2wlxIVoXthZ/9pwq/HKWaoThN
GTYIp3c2/jH6ZMutOEWZkJjNnG72iZGilr40JnpC/m31O6xAxwXlIOBY/EVB
62jLS2Dvu+Ne7oeeD2CidjxDv6M4FUI/5Fboltw/7oHRUIikCC79MlpBy9nt
6X+nuYUEtdUbxkxbrYF88/ztEDe/LD5W+CkN7M73WNsbr97RieX4S+k7OUdv
w0JBB52pJIBjkCGcfCAg3X7LXAMs8urBGujLcwOF8ah2yuRe6UmBB+8SLc+3
crTssUVxgx9dr/t0b9OctVwP3hEVsd84qK2gBI0Mk/6flvsTuXBuy8VtSOBV
rLOvcP1MxjyrEBPilsjwN79nOR/IyZngOGOkIPefRTJXgktFl80peRBNXzC4
c5URWc17dcvv8IAGIVGt5JaPcRpCcNV5KOnBGO00TmcABAEjp9qlT0qricOl
KgpRqCA4unkb8JU4Tbp3Uol+ELDW4RUq8nP5zB3uW7Sr7ewkErN7K5k5rdLF
DnAfTpnKaXQpymFRdaGDe2XuTxwc+ydNZWfDsx00QqhRjoAebHNpMX4i+c1D
ED+VUXMUVsgI3fW18z3uNQ3ePXPBJYV6w0HJ8k0k4I5w0m4ZJqM2aCfdgWBT
FXzr9F/gPxhiivfZn1gTGbWMWKBpY7dNOQVb2I9md7rSoCaNQly8AnD2uk6I
lv2ZERcjYGybhYPz2Qm6nGzrZzrxflm5WnLVOXi0nTuwWTWgGIbW9drEOuCS
VzgUUIyXC8RtlrWx5CL00RG9fr4sho5xvHKBk4tJvskZNCe2nNY0cnFb652u
qePGqAjZD0T7ENsvbViXnJk3wI8ZHHzI+aG1h6gdcx5tEWX/KGRlOFzrHQh4
Zc0VWIK02YAlMtwr98w2FO2CUNu5F4whEpN2jQczy/N/3ChXwm/7SZb3DAzO
HLRAlPVYxlTp7aO0OBv5Isr/gUKUkzZ3yo9tOAFkJoiPrCS0QLlT3ryShwZS
neKWQtgypusw0di6B8ITA2dZKj4Kvda77LoGR4Abutby6R0Jge1AdkOuVtVK
rnDuoYhGzUI7YjJNpV0U5Dm34V8Aq9BTTaFK6R1F6HEuQWYXaT8LUzp0wWZZ
OQHObG46KB7epgDt7vGF8eK88DooHifELpuD3Kl37FxDS9eWf63NvDNQc59G
i/Yhkon6e4fakhawUcOfmGfr1hhC/0d3eyPTANGGQ/ettOu/dgG3h6+t9W9D
YkSC4nLPdBRFr0HvCxEkBr+rCz5zpUxraK4hzPDKIjV7QOpdR/ye5Niv+HkZ
j2YYe2jyiT/4bLZbldG6gpfbFsmVAihtgz92BMK9reCElA0AlLrTqncIMV63
X22bbfyTX+2pDv4RCv8H7DxkKGfWcAJ1HPPZnGWI2s9+xltiTjT+xIQY89vS
8Xt/NXKWofrYCLqIWObPmyWgngCy/IW2DeYFc8S6nIZ6E+T1QXS+G5+F+sP7
W9/oE7UDACLoV3wVLWBp8GYGDRTEfQ2f3FA0sE9HU9xsbfs3CYIIHiGzRXR1
mpwGqnF2NB0keMAIcG692Rfq2ByXSJM1IJeGQXBKvPXR3N4OQefZPsx/lgv5
FdlyH7OJ0MiNlr0e6QuGXyC5L7hDMm4GqdEwQ9gGiF/Obgzzeh8dnb3tjJGs
axgCxSMQX5vBCkMq8fkqrMSaYDEtNESze4ioTIEb+k9QOCYRohZnYCphmL2J
vITn8P/WPUSV/BSt7XdykdWQANLIyk3UTw+kf9RHeyOSThFWbRCp1vJo61da
bO2CzvNc9lZ9wuDNUDa58Pa5am+MSMYGr59IMykpu/FHdc3gZYza/dTCmrl5
aw9h0fc5404dUU4aVIENho/nM11y7RZ/HHQXvHZrfrQco0DUksb+ikN+fmhX
ZmfWsHEcyjUVHVuHwyoiKOH6OwhNA6JOx1/wEtpH5b0RswQTv4mnCbQMi+XN
ARxx6U7EOSbNCh6hb4HLwTvW2Daxm/5TkjhjwTf7ybDL+PlKw4jsJSjDDkIY
76DvHbx2p+iu4slp36QdBSidc7kXVdQ7WEd3lqh5VPwv/QDiIv812Ih7Hq1H
govn/7oInQO39JsIlJpabIkcWeuRgiYJzYLMsuD1uiv64YNGNaj75i/BfDtH
s98IGzZfh5H8hu7h0OOOEBEPONwb/Zj/Limm/zy65KE537mFtntdrycW010B
tiTxxQz+KvlkoVpXuM3ZZhzKL6hT5zGwD8hi5zuInFNZ2tIp3Yx46/jZ4i6O
o1n3S9JJNmlXsJevGtjlEsYHs0aqrK0j6XEwxJ7INl1CEPczJ2Z5+R0M54nL
VyLNFRvxbH1JaKQlelL6mX9JpppAanvg+NP6JiOY6BmfUrCX9M/fwoXU5JEx
GpCZhw4/ir6T+238s/5aCmMcVfuHsDakZiCQL2hGYO6aMOV4gCx5DilKnOuh
0rSo7hXLtof6G/C9ULfnu1Ka6ICbawA7xxFaZ7zWinuMfsOuY1yQdRHQA30w
DzfsKAvI2WouqUVPTccxravCTxOssaQrjdSvMc31ipn0Kj1hyefuiKkPAwyB
4q4SgWWH5a6TP1F5kKfZLRSdDJ9rzpwEV3UP7iNccR0xLPMLLgqgU8RXx6/b
5tavi8mEYmYf1+IxOmECC1W8BRKeVNcLpPeuPzbbyQEH12WnNSktVJtDCVvM
z3hpd9ox0aR2MLcAw1hE/ThFVGDE7JRoxpAZUwPzjkLOX1MA3V7lwSw7QKxj
zKzgpySCeclGPLeEqWmel4SoHKgufplLD0J5JZ83UgowN3YoCuUviYgCJQJB
n4iqSPVMPN7pnha4a4wPvCBbjriCYSWv+A2iRybkIRoO21Gl2vR/Qz/p5tCB
r3HRkVB8sb6KWe/arGSEj6HIUHLBdIsClLoGZmc16w+mSH+AlNf+ztTSUsgt
AEHY2kyACkoeC5b9Negybw4xutv2WxLBYRoRFP+A4z3qudSR4vahqPfkABMV
3NYDIy5wy9z4UfcNMZiBAuIasbcx2BT8ylhpaq7SOWnNBiLkLM+x8nq13s21
0aMsP7Ub4Coq2OPhAO7/2klQUOz35FvGR8jN0lU55bMt/tyRdUMGoDKOAI+S
N/tyKy0M3JbZsuRXATDM8yoW6l4RiFjz5sHU5WHUJ9jqhe37ilQlCPJHvNBW
sGcXrLOPhv8jQbZ9VsXWlWNlch97qEkQ8efGW0YAdWDIGihUsHx1m8+1JgKr
ctoik/WCSfDIxVEMTHenXyfoUu7KS7ZkAscu7JqySDhRuMqtzoZ61wlMdCWT
Ai2c4oqaM1yMj4RgBovifYl4dfP0pkaq+nuBh1WUx3VbWNPAt0nh9EDjB5lo
wzHah2Y1H8MB39iMKTMTdIZjmoFZFbQZjzGycra0jxnkbiTl6MvSML3C3MWQ
uFROAqfrcXO70Qu+hmk7VORvMVO+jhxJOYXzs1vwO27syc/WbCRqEr7p+ooP
ywqaMs0vEAVUxlM+BPCpaiCCa/ZoNIjsXXsMcI8VjRUTiTNb+Pdo2CRQimfL
SfzMo42VQ75vRrj80/qt7S+Lydf+pJB3omEsZmV2Y+3q2zrLHGCFZX6pxt3N
+FOxIkLviB+9BkDLc3apC01BJbakbeC8cE5HFIrseySg1Ru/OXkfgG0zGhyD
1AEMpSBLokXwtSWdbtRosGAPZTYicxGaOwHNwezypva0Mvp5xMOFba5S3Z0H
nf5CmGlOajW2ToQY+7jogEanyYb+b/Hw4Xbo6s8Uml3ilfNtyCFn0h9pPX2r
4KMu3D9Z8PDhsRH7JqF5kB8ta31lczHmIa14B3RjGBOumpCUfLdhCRvUyyA/
ZUcZ99mRsItX2LjZ8Cqr6ftlUcFuVWTCC/U/B+WpjYrngsOQVxO5T9QSBPjC
37e6WuwEotWeEcns8ODoqqPfHXOQFt9kjms3TZlrw4+jOzziniGWcxQHoylC
OHxmPWl2vzmKkZQaxpOMIOoFEXeZr+Ze0yOCsTfZmrQ4chbYJqRBfRB5YQ/9
AH8c5r6w23fHo48x0d8F3EF1ivMkxkDR88uVWSocOwDwWv9RNfMekxkLyKxo
TZAF7tHl0D+4pcUBv2b+poJc0HNEpqNYyXbUKukHOnzFAPbVg6Ss1rKhn7oR
YfAmkMcWdkdK708Ly1OJWzxUCWzCBnvL3SyoAj3WGAjrXuXLDyqZJEKxJThl
BW0g31BEiVdUx7TExyelnrc97qAKVpWPgvI5CRftfggUGqRGpfc2wth0sz5x
+4VuDiH9GrpuBXe+gV1+N9Su5aIffDMY9XzV0MN/4GURkTrpX4royywVXpP5
d8wD74RvWb5IFYWdxorCMXfMcwMzMB6xLiEYKg2iCI/ktELg2ObcsLdE6Lg3
QDd1lkB/CnS145MW4HREOIXZid9d01oTddCF+ye8KycJPcSn92gPPiK7nBdd
zMsfJAbCMTLC5bG4Fqjc+copaH17GBGAM9ru1Lmp5Nrco3uD3hbpHmbwSN8m
ZEQpbZqbrAUPbaAIRuIDd96CgIQpu4My5Pptn9T2XP235KPURzX8phF1fdfA
3fLhfFDNaNVoY4q1t2a1dVaQHnPFdyFtu2NLvbLtRyP4OXJJn1y1R8q3xtva
i0pJCPk3HnHubVFhJg6bNidQA/aJNZtZTCYzcAQ+VAUaP/CzVC6WjRq08BWY
89mHpvaWKrvaWDPm8fp0flerrvsxmjHkhEBywRs/NXlY5lgPxBBaG7Drgq4o
VcBtin2Mvpmp+8UVK4pXflObxpUeZS+PMbea6PVug7Snt1pn1Pni79bKFZWt
EyEz4i95Ge7eEE/u8SbYnspO09cAZKAXlGQvcr7/uE74yXunfaQNWCpyXzof
6xDbTEhouavTnKR0dkCZv4LMXmSDorgEFDnL0xzRldfShC/t9Y6oWKetUc2a
VwrUnG4vw0tgZQbMxYN2v1dVASXdzydY8vi1NXkw1FvZXl4/rg0KWUz7c0Jt
v+XhD1qXxl9HxTUb4lcrIYFjtNkzCYIu8lFXzhLq+4bhPMlAqh7lHVE7LXJy
dDgAfJdSsoy9fgkavTc43EpclsWjCvga365/FHs8k/6nl1we80lCKGENFVQ3
F6K6Wnk1zqcyB4kdRRsdrB9QC/AD+fgAHqmobjt1mdfGVZ7f/zJARVdED83A
PGBg+rdCers67g64EV4z24hmMT59CfP776L9g1mfM1wNBiUnhlM7PLTYivhs
BL9FklTWQwkc//OxGjfULEnpNzoYvVg8GYBU20L+tnzgVGYydcLYwVAu69cx
RQb3nouifeTT4FInbJkevO3OzewvRj4KFSxseTkYWkdMbfua/ISwZE3716oO
nA7Q74dUWXwJsQS1UXk3xlyD3MJxPbv/TF0VAb9aAf3nIz23wEoV7FDaj/IP
XsqMpLflyKWkmZIJGhXyc8fZwlTDF9Cf0XqKwQ74Xi2BKpgG1dr0sDmzrT97
/aveubn6rwkw12ydeC1dw980Ybg+rltQ5YdBR9vaMGSmFicUvOe9v7ufW0sb
Pr5tXSLdAtj9gaaZ+0SxP+gjxhD/0J69JJH9YlXsuw7WByuRGJM8bcmdHgiK
glPI5n42PRf1dMbjeh8xXA8/Dz0D0vEbv7XPXxnLubBH6IJ7h/GZx0I7xyOV
z6/NRFjcyvrJm0Sw1WBuqZYdkosNslixkKcycHRIl0jqK2TeeaOaqyB8WvFS
zNlwepY/WidT3MQ3YsmVIqLbkeG8pE3XQ2SI/Tza9Vt55gcW/jK/y0vsXUZt
0cAKp1NMP+FZcKrOOHZyLB+GUFoej1eck57fYdKsfuOGYhNmIZW4zDiJlQeg
dDrwa9tXMSvmpz5KRUohDr7epcpHaAuRbKew9JBzLLbS4/VrWaxFdJn01C22
wC5Ny5vx7TJI8OcsSHPlx6tHN2zKl1prrfsTwocIsggTxey08xJP8rgKXI5x
8GnDVGxVDo0gjDqzuhX36PoObX3j2iYY9ORzl3QY2C0scV4xcLmyo1lKzNSL
P0ldT0UrpNuR4i8bQ1Rl9J9nmP+KkCvZAnLbDNeOeTb4BeMrfaK4xvY09Wrp
IifymDun7iJiU2dYTURLyglA6RQq1+/DOvD+5cJNA9WPC+P3FSyOTvU3Gyhj
FKMle9ZdMxZFExRGz/8/E0vKV3moN+0HyNXeSAtxK/PXlUtZVo779NW0S/Kw
iDme2Sbmr5BmlINyjqpcdUD44QzCxbqF1oWw3xzqM8xYIS68+yfwGJsN465e
KN/BhVhNYa1LOuvFDuyXBrgj5CHm6ndXLYkcgaTlV7AfG3K6i5WpINyL1OW2
AYJxW6IkceWyRL1XVjj+rKYOIgO63QlDOEEu5IZbjpM+inhhfRRBrm13vKFv
Wnl61tDDo3EaPqvj/WpEyQp1iwEX2U8N/oFLuAKupzCinjNogse8ls+AxLsV
EZW9kuc27G+dhRS4O1qcnQnoTbZxHhsdO+J0OS0ckZzAx20d+DnxIwLblCgK
qtrSwTZCnNlJKTN3id06hiQIwtwFau/DBpEYxPzzwA3pVuE/ibTG6udEnT82
ReJigcyeo+CQaxPqJZOf7XnjUIesFs3lh8ffz1NkgsDfPKUlrZAVPbaRYvg5
9fZg+GXZ8IJ3TwHv1vOk7c+fl3n4PPMw7jFmiql3C8LlF/BWofnhKP7pIooo
1YIckVzRMqJyuUf5LEL19cLLJvsSK6wf5GuQqqc5JwRpmhgrXe9mWs26+nKC
mrbILebnC65tiMQv7TeDCqdpUOzelO7jrjtIbf3tEmcxFA6qzwi9di1NH/Rt
ZrjVd1xf5f7N80sPOdFZtt9KsM+q9Xx/pKTYunz5wif7HnKMBgwOCcZ4eiqy
8yXS5OYBgkGDH1dNJqpfcyybKH2lezjVru6sezbzlM3Af8z7x9lGSKGL6FnP
ZIqQyGSFSEHXUCpnUV52KYH2qa33USnia7jfSVkijyiQGthjPFdW+TT6Kgpn
lpI8DbUmBGpq9a+wByXUd1tgEJ5vk4IJfzTgZYnp3Z8q2OVdvzm0QlHDgitR
/kFL5qzNRJt9hLCHOKMV5TDf9q8sDTyWyoPZoG86ek8XWhyvEZN9MmobHlx1
52rBTN1gR6LsTrSm16MQKkE6UaSKN+Y+QdOXvekWV3pKFXCkvQQf4EzKAPha
9l+S9NRMo6ZrBv5ESKFJp2fWcC2W4nsM7dvKkce7D18yP1GmE5rYY4nEGOEV
hu+jLdXS9VL4ijjUnNR65smBruxusB2/wj6gPhmETpxxQMW2+h4s2AjJXi0z
5wpvQ9/FDgZRqDLOYBK496nWcZtyHFuo4EgZx/E1dtfFiNbJEGMuRQ3mOn1w
XeHeUU8gi/0YouV6oq2NVSYwEawqzn/6LUlLVhP2+Z74lL98iwipTzRj6QWA
hAMMQNMVijcPcaw9K408pkIQEtqvBJX3yy0ua3LKsk0YbThBJRYbdu/4nJ0R
OcoOAqjYRlYbcgsrJri2gQFiCV63oEwZhc78gHt16cr3inccpTyi6UORTgcN
nR+R05yziDQrN5AzCZM2Mv/BB0wWk9/337mBXKK+RpV6GdyIuDQb1N/D6QcI
XqJIZ8dEpG+zOpN6hZOCGDkEYR+cjWnYv7oNRIbV5catztvAwtBKH/V0I8MT
PjPdFlbLODQIVE01J31yYykQMmHjYQOHEQMici3W7n6cPd0RmahYMWYboJfo
y97qrd0iDtE3weVcL6Ut+HHy/DdCKzbiFb5ANhme8P+7y13l0u9B7agMh+HD
zyY3glCVzCyK9xRzDookHsSGiFMw6gPDe7Lir8qLpQ7A1Uu2w6EwwdKXm2do
G9Mx2Ldh3JxMb+DYJrqK4aLKxahVv86FRYZbLfGwfbHmP9P/Md9BcNiT7KTk
/ifihYkzbHxnP/FBNKNLnHmOFgs/enJLCh9EydBx7L13jyXY5QZGSMVjNa/2
+bwY7oRAQeB0CoWhyuz8Z/rAqR0MwkQOWyWcvBWfmiXfNY/lho74r1b95JMU
XKqEMU1k0Gk6erT2BzPjBQPfPvO94nTHUTMJukIAahqWJYUWBOZFyp7Ds1ju
WI4eXSIS6frsDkq55EvUvgC8HYbktYhAX4tWgGmbHQuo1aOKmhMdrYqpKGJn
Eq4Bosk5EnpRYFvr5NbTAqYjnteraLoljXRp7e6CsUbW/lK+zGLWgoSCknFN
y1qGRZ12inbyCcz7yItBeqY4Z/fUtrgMpSCkHwSP/rDzcGdumlyZ6wjDCIxd
IAwIiCsTsuIo6Lxt68QI3+wAC2HrXkff4iO5jdojzJlW3FPMx9tFIT/c3N65
3eZPoh83xv/cZ9czCM3knXN3UVBCdfMHc61FHXGvzdP9tgtUC0qU1yCvs5tr
SCtQpEQ+PXu5hn3a+FxFpBAu9X7DQjlsI8UHr+F97JqmSwOvhUteiiuuh7iU
1tM60J0EOCMVio5HVKd1u6wNyV6U8f7/VOXrAKd25wrUHjPPy6sjTO+xITkR
jtD5Nl0r5wOzcjAw3Qz/9tEWQIw8AYfUF/VDtAsLsCep/IntuNCG7lhGt4Tk
CGA6Q/xCk89IvV/G1CKtNwfXDlRvzxOgS3oOoL1LlzVtCJvbJkYv4fLO94Z7
KIXuio27nFq4azZ/+KpOJFgCU3ipKfPZ2ljyGjdeQlsUMNxlfGbsj6eTHQdW
ts1Gw4EagSOf0aFM97/3rf0gbvsBpUZy4OSk17SoirDpADOOGLtm1EDg72xS
xrsubX2WRoX4qwSGzUNvtZDuK8XVmqx/TILw62TeYbMI/+k9NxDXyC1u4fvb
+P7S14q7e9WsSuLVLsBLTT8oJ7vPj5coxRt7qAhyXDs6qLYZrZB1KnKckny2
oV3p5tXO6Hv8HMoZgh9ZtCFeG+w2CAnK8qp5uPdD0b9Iccwrb8OWxInE53tK
F5hszfigRX7Lc6tnZ0LK8V+sKWrxI3nDuOa9HqDn2VxA+DTa6u7J6u4ZAabp
gkO/2DVwKISFysz70J/YOnBW/q/bf4EZTUshua0OpEtCaXEnfhzLAqQ/hdp1
u5ffK91aMbCp6x627sTl151JpFOrEOPscyGRXmyd2f3o6eppJu/SGySG18O+
JyRg2bdPJFGyHZFM/0/6WwWh2UNtUVt4+r4cTV3C8RvaIp57DqKSp+y6bdMw
LBOvl0LSOSLOzxY2j/TXiFMXtcW+Ow9nuri3kq7M72vmeijR7o6qBoWryM7J
RklLPBGq2QzMFV6lMXWmFFZBT6QiD6HNMGZd75CroCCIC6YazaIKs5f9c+aF
R+VnudMtXxkJ49NR5H0ynxW7Fx0pegpfiO7WjcNUXMZs2D4QjXE4QiRol7B1
e6iMdtdrtG22wCZys2xH2LwTSSaZpHIovpaQtYSXt34rfPyF8lc1wsP/PidS
kqwzFM6e5JDjRn39puyDGIaF2/p0JNLBIlbguJgMmWUwp6mPKDxBA3/VlC89
sH8xEZNS0WY/6qeW6Nst/ful0XMlCZnFYoZlJ1i85mpWg2ySOhSkcJqtM5yL
CJzZi35FpW+EyXNbQN+s2t9wG0qSitFut00+dYwWwESO5lCC1IIYH+QAhDYO
SLsA//fVtV1KKoS68t2efRmF9vmC6PKklKLGSjdkv0ri5jIfiXnDvfbL9n9h
+K2c9eLIvguSAFMxViFRsTdDH14eI9AgmEivFtjxqVTt7hxFOZvwvm9Uw/7n
92ny8ZKE7qGUoPm46Ys4YN/v9SIBoyFSsNrlb63ReOYpDf2Y9iF2PDbmqWu8
DzjUAJA+yPnItr76YfuNZNy4LWEKxU7trQGJbxibiWGktTjSTse/i9YvECl3
vTVGgSVp0fpevJGHBaQUNF4WXEMrGSjcLhuI016iZmWbAGdD6vH4EKWew3qY
DlEiub9f24g+z09w37siuMaLFtPo11ms56GyMVqVqZUOOEJsXlfacKAku9Ed
dju6AoRZTz1hVeRTsrsXSfAVdEOiJT6Xi8ghzYRyYWTBOvESy5mgZR8FeHPn
SM2FmCqS9WgkLdUs+QRIi4FXaNkIIk+UBcvFKDZBNrCVrM9OWP7SSyWJq9lI
VR1KT8WlbLgF8ExYb6syFH2pC+9k2wdPAW51T+/TyNISZEnnMJNDUI0I67Qm
rUNChKtDDWiM0EZ/Ax+NBWcwQtzaBn59kFe1S+hecbI0OKhPU5ZHSZN/JCBv
HBoCkk/SZc3JTrOTyXMwtRpoddr/RSev3gK2+j56F5iJfaySnR27QUFH9UlX
WMglYAoZFbjxi88PIsG5FLdW55eOegin5bSFdQ3m80fALB33QftflSzMHAG4
H/35em8TtQISex1KJpkqoiuDmP8rc/NPnyOzuXi6a8UnBi7pLtsmNEpBc3Jo
ki6zDc45kGnDHvFYIZVZCvWzY2mDhmFPZMNmHrCc1o4a4l4f7upPHHcRFMDR
U91oGuQJzrbDBQOQ/59OQosbymsHcYNKaIH5nQfRGnEGSWS9z4l7zIVm3mzJ
5u2ZZkkVg/D1Xjix6W3QQB5FYPAyFmAJHNnRuXc+T/n7kE9K/Ml/djNk5eMG
8fFwvnMVCEm82E9UdxO9ywMKaac180KrbUvGw7NF66eOwNzlAIh47P9UgF0s
hnZH49hvytfu/Z+3Tc/MKrSoXBtGEnDAefDk6T/ZYc12C1EE/4cDypukEni+
T+v+9SXcqRcJg1/ty3cvxLAVKuZeUt64//JpWkzSUF06evoAz7763e8mRItH
fbiO0GsG+MOXJYd38Ad017dJF4OemnnfeGtwc51a2n37crl0gUpLzc+LeH98
alr5HmzEz1gHWmmDxioOK3OYdei58AqNTx6PLZ1Gluc7KOm/pFBJC1dZIuhJ
+L1ahRSvtFJjK/CuwMhB3PWov2Ju4KIf4Du7gE1Vom4Pai0klSQlPYHz3+Zs
DBffAyhQOXuoPqRpKkVm5KdSdzBU+gpglkDhqCeKjM2fbOqWXpbdlAE3rL7c
KE5zVV78qAcMBqvdAcrsYKWmIdLSoFxQTw/fJ7lUwJfH1TZ+yrUjAKUNgdxa
D2joxyLU0xiiRcdqMe4lA5IwLPX7Xc83M7GV/Bf36rpdjHB3Qd5JhghXtVGT
VmhWBX9VXF2qVspDjmH2ktebg8VEkc8iLJxXftHB2aRN+i6+dR/whTz/YXZD
XWS71pmVwGpiS242+npIWPx7GEe+VWue7alT3+Rcg4bXXpJT3ljUqQI3w+UE
7bG/8Z0zjXcpIft9tBYk66gztSo2FfH8kkj5yzjKrYwJ7UBKE7rn++lUFSIP
X/jVwwB4GT3bKLzU1qZlXEqWhJ9yaQbwzUbs9Pw5ZnP4MHqTKcVUYMytOL4M
k/P0HEChEb6sZ5dp5JD3dpH9KOcx5PY7qkWrd9t+36zwkug7iRuUdGhmCnUc
ozjwcQAeDROpE3YUJUHeUDYa0KfHBGTXDAhVAQl6fO+EoNhk6X8U04QraDIY
7eC7VzT2yFKU1VrDIuOY7otKu+tiyZBgadQAyldIEyxvmdxnpa2Y8WKps+Oq
AYCog8It097QQ6QoSeVtHTrAOTiyStB/kas4+6r1ALUkrbDbf9QzqlsB5yk9
JDy3/FRGaClZqVLC5K+YqJVKs5yYQJftOMFRLolQV6UGi+oR4wwAxKgRWVqz
obqVkrslOYSm/sGRVP837A7uMre6tWpB2XYs1n7lvc5gLRDyWKGNSahedsU4
bE6nWV4qcc1+5HCLgm+Nd3Q0+F9XLIW3hVqIlP37kFpwkvaca0SWNFryKSEH
Nudtgqa8rWQdjAXmOCljzfOhizKE4epzFxtU4qOqPqh6mhEYyWdSQlhYQq3U
wvOcaxbRcnDZT9ENkC4TuqqIOnv03goqOtAt2hc1cyS7ilkt7xxlQEzMhYlt
RpDw/Z6lMTngNAT/YZF9SbAcoKSfET5tYC2sxKcdlDfb7VIFiFcdZJo9Ts6C
5ru0HqSFISgld4QO7y8RVTfwyhjEwVblEWzDOIQ9B1F0Y2dfvm6+r3+rQ8g1
U2ljATZYQNJoUcLnzWEIb/TU24F04apO4++FfT/dbymFi0ClLP0JCEGk4wi4
NJDArO+yR9f2wikw9dhLCFOQizhISUDQyQEmGnnSLbTUJjx+eSIWllSXbs7E
AokE/NCm5z9bq361ADFCktg1NIiZJXnv+5oqVYOeRm/6lLcs5+11a5dg0cyi
jY0jbp6dQweA5GXZ4R+Rxno9XCEpcMpjUT25kmkVPiU/kUrX0KDPNCFo9ivn
J934Vuu1RmSyp3+eNkCdch53IZZurQ++DUtNwyuxzQfhDcgKWFHflKybPpTK
CiL6sgrlBAI+5+4eMRfirkefc55IwZB4aEbRyjCdrzZuFDeJ9nKee1H6i4H1
JCLxNwDAzs7Tgsd8/Yf3y+HsAYYQJI2TwgT3ua88yovwt+78VT05Ta96wu9h
A+kTF9ZoEWrffBOqPfg1dre9gQcGX/gnEJdngbFKQ7CspJyHIUbXq8mUkbEP
p+PEBq/S7x0L2p5mfcz3fzkLCnTFuRKPRrobUN8YPbqFhiBM2nQ+ORa1ZhOs
JbAEtIv8lXD9zX6qtVcO6S6CNjy5SrN7MbbQVHNIwOWtuAe3ndmZoB5eWipe
VUTI0H7zj0y7SY6EIvAi00Nrvgl0zHuedMZBSv8VrrhPFtWNfeW8w8pfoxCk
cirdZ6b09ChFpWKUPIsO+vvvwbUQ8Fd3gtmkOTAbpltynyFYHIwxzfsmluDF
hQ93M4q+5/mhHscTNDyIKDmscDuusstkN9hsryy7Obu1NrIQrAkNkHw9xca9
GEQvBNZbAyeN8UyIdl6MATOKEIu4BMRgMk65m1lUxi4R3aM8SkONwRVtLOZs
M5A9j0f3o64+sCsF/VLwZvmcYYzvHDZ4j+tijY958vcSfTbE/YIoWXZeM/in
7whvjqeJnTeDYGcXsQK5bQOSVpMBrL7k8lKpnZNavqig6Tz6mjGMfdPAOodL
f4HMQYKKFrsmC8jA368wORjvBylsgZCHrpP+khto67mB0ld5xqMgTydZzYgV
WGvOvJW7D+7KRQXVgJz5hK1lLznaWoK7zsYNUKGakIV0a12txe/aldrX0WbD
VasBgf1RKtHDGmtfLtBEFPjtOH67lgIWnglw+SBKnIUuHvVQXUROEX3gXd2N
+gkTXvwzJsggjU4/PCRhCwCZH+711YkLOH6bDyaEGyuLju5QerzSAThx5Jxw
xeYPCJ5W2G42btkhGvNfAyI5o6vr1pHRJq8p/4ESiss0MTn/fH/1eTgifzxF
aTfcf9QWkZnrSv+CIsZ2aelwblgFRYljYHfNyQ57kEnVbzmfF+04R3m89Joh
T6wG/TPSnqElXqw5HPUcrtRZMimStWMp66XAQt7f89Ki7/YXY5fx2yzvbsUX
G9vJoKklI60u0goDwSVlFcQTlKGeMwTXjbFsD8GSnSuAW5yVBFJi9DA/8XjQ
4cafjlMPZ3DKf7JetrLofU271LNyG0UTH5ymOfQgbcHI+WU4mGeVnh6peA4S
ff7XKDUw9RQJVGckFYULXGo+3ujo8ZLq6xDzDnctmPLc1C5MEafYMdcvRgmR
BwPK7N6E26JMKV7GAa+ukJulh5xsL/Y1OT7Ti7XH9ke0QnUnw9yJYXURrXFi
x4X8TDYfJApq3/NZrzZSmBYHQMLD1feJyRpEsk+wJNCSsY4UHuphEe7Fh96f
O2OzZL5+NbR8ecs3lZ8AWhI3HA2d1/XH7UXMEEso91kAFk8PWiT1ZIV12KFw
/qiJku8ojRneLmM0fLYo+ec6fm/c7d1BI5aDxlp2x6wQNUCo934tC/YIA9kf
F+L+9tp4mqd0rOhpx2N3MULx5dCu6UqPKfU/jUUSUHstH1al4WRHNiHoVOnC
kxHdQ5Gf+f8hLsXTU9q7+aVMN5CIrmMeOXaFtHRGB7BzjT0nv4KDn3YFeQgn
QiQhI2vasUBFb5b002PMYaLF81kk4Rs0LUc0EhEkaXp0XEs/FfDV0riY/cFz
OxmB2DZqPZ+evkxjKIGkalmoO74RYACrMSxHi+iAF5xXlon82cNA7iWeJr8F
1VaQW+qrOZWhxbVd/ZSAb+uDZyrkc358m3LLCtoDb8Ktb9ZRk1L1kmzZG3fg
OFmLY9N7RlfBFxSeW0WlZ+qpnKQZZ3gry4Uam5d3xg/Z0mJ6BqNGpVe4WyYc
XNZSiPbQ6Qlkd4M3u3xDwcXrT4zSvJi9bq9nujIEsM5Z8ee0HDxEcNdLJUSh
3Bjr+9uDehx5VLNG/GRmfrbvYziM02ub5ANo2oVVMMdPeNLiymroj6NuYcOh
mmxL69+WanKBaXRPnz/JckyN3o+rsCBNusHCl8v2TVOd22aoeUCGnrAbyqaq
hYPJZ7F83FzEhE1MFdHVQsdWEo82UzxvmEFXZUbv7fhqpR/Gh6wxCeL0TteS
82fRdrkEuNIW+qiV1LU2bIAgGTxq+TJwe9aVZd7RBkTNXnmVJGGpjNlYVs6b
5wUBmtipUUn9bOFULWYHalGXpSDo4rxGGwNRlrCzmoZVYIevfzRqbPJFMZ5T
569B5egfMr+/i+Wazt/fKL46bVYaSHnsofC7Ag1Oqj54FH23vDpRTeu2IiGu
kU93dUZzpcXrawNgKDjQrMknQc/7sZxa5ZTQhTVx17vmZiu8XMY30UDyFQyY
EaSx21tqGWY02mA8J9PcBb/aMmu6+OmJDeZGefDQpzd3xCoNc/lVN9vVJNGs
ryZ5NMsrhhIOlXNNkg77DHnL524+Eu7E8NW+laK3q/ZiYcDl/FYnWqeaM4+K
XhMrK6BridTJIt+Exq8/Izur4YJFgJxIt7hLH+32x3quJ8LvxwJTcLnl+zvF
fwXVIzRQPPwyFzTZbqicOP7WV0256f11K6wIylKpA6kS7hP2vzTNJrOyqTAZ
YFDUzzxf25WYlfjUVXG/iPqbiX29Y0/xG5X3n/kCfDOujf3Q0r9+X8P7ki33
MNBGwryyOtywfJKQBn2vkT5w8g1bo6r/o6DVT+x2JG9nluD7s2aevQTZa2YR
LqfMvtNyWQM22Bl6SenwpXmbWAn97xv9RK0iFAPYPR4QR8UD9/F28bFnClN9
jgZKZBoxIaobV9WcQNIAhxnG7FmZzQlw936p808/emstrKXL/8kAZgyt1W6G
vwnwCT8yU3Lck/6bmW2jnzyTJziQngTbt11ugTi4HXXzxr4M0SkkZBQkC417
yjWuS1xX5m247cPsJ7J6XRhIvpdZ2Hom+DQ8d8x4OMW3I9ashwnWPTxbGmWk
wrXWJIOietMoycnWhvdJm59TBhxtqobyFzuMlBbGS7njXb+BFDSA8bJ1EnSE
iDtHOWJuEATkBKFapR0kBOirCdVi5utGW8JXm7c/3yiPuJ/mw46DfYbtY1bj
ctxSFEaeUxXtKMYQyVLStfGVtsDm0y9tRbUytKU/KoQhc7T9aHATtUtoqa8b
4iyCLOY74gQhBjfusQppuK9d03L1YdMZuMKxnnMI3u/pv55XdEX7AKYWqW5h
QXHNST1rmST4boW2TQbbEDR15zhnoAgRtV8AGiDnjPJya3QtNZFyqDpr5u+4
4YWEKpwn5uXqpGe6sHKYiZTTopvHOBOu85ueU1kVtKkoekYDrCBwZ7igSsyM
UoGY/b5DvlGi0q2r7XSJfQ3YWFg2rm/zDT6r/fmJ+lwDmSwZKk0NZPvp3lTI
NOvf/zQEBYqAPsyTHwactZMAuRUoPLnTxGaiyUMb6grh4BpTYpSxXziOGZIw
i5wgSlY54qP5LADETMoJynnY0TkqMpEf3gpUKOeqvErUC2EQFR7wcD9giFD6
HSDT1nPfFZ9V1j0F18iA+4xm4os6Qx5zvARt++UWTgb4yVcBy1F8rOXc+DIR
rw3r3vLzCcQi8zc0AmJn7qDhYh/7cDW453EfLWOtCd2gudcQ3tkTSyt/w3R4
TFjSc5Y+vRI0m0MQh8w0BNc+OJMkJySH4YJpVvJnUYnUCDMpsoeSvuD9nl2K
TugF6pOLXu5XzyEGXiFn7ropr37ecE++FA3bTrH5mQ76kkFS6oMlYWiPbA8u
DlvffkTZgEYyQdXBu2LE9WbSlbZhYSgpGdAWZ0jZIPB6KDJtrjDXZL9rIwgp
xlCCOWvPlVUnBDKFP9d/pk1/3ZhywWL9L1HlEhi3+QBWzEFVxEV7WqpSy/WX
THDkfbQStdNB1JycC4BSSaQaRnQ+tVivfDmqjDvwjUtI9JTZCUH3XKe1DlUw
vvSdkPsvuJsONRBg1sr6G/aOOBjqcGpPEG+yknSm9HhCNa3pQwTBiEKYhoEG
/NbGZi2B0dILYAHf9iXFj5fmcVsWJtS5FTE+b+cYLzKMmFQELAkd21FmVR+o
YX6tnZ3qlkQVX6rFDXmnyAo9hLqTU7HT90bSU0X7Tk/AT6gsvMZkjlhLmie/
87zJ7NqBAe2qE7dAeDfeMgHelcdMRpNWC39pyqoczZkkCPygYD5boD6GLEkg
sT3ziFfejG6S8sMZOuZy+uNE5X52tMAutQ6lpxuFyl4ItxXhW4bVx0DZECQ8
JhrANAOT3eATf56Bs4BU6Seh9MaBuRlJ9Wnq5g3CobkNDPZNx1JlVC2Ln+nK
KyFAu8UPm/5GZAW8+P9tKQFQVHvAfG3/6/oLOSmZhU7VwDLxqxDL9WxFmk03
RY2VC0fDV2729EiL+PVokpvXp83lH9EaKgN6Zut6LI/VOClw2bxayx/s2PdA
FEjSa1SGv8OzWHTbpFVWUYc6zyCk+IJbEeWoBck2XTYzYwz0+NtkADrO5gTF
RidkC+LatWBbKwmpnU3Srj3ALpa876MtrHtwi5nYtk+AQB48EtWL0mPkCim+
6azZpZJadVw/DbngmpqaEhpmZgT70kQ8xMBBhBo3Uip24i23o0DFVmu2/LYv
lu8EKOUmDDwGoArvvg2t0utTf/WSUNQb4a1O0+teOe+4xFvz6qSgdU2bSmHa
OGRGPDFWPac2Mo5aiLlzP2fv+i9nrGSAU1rxQ8Q8oJPHgZcuzEWlSY8x6apW
jeC054I7YnAHJNhbPW5MPwMcGa6mnWoUN/Z8jBltY87w/KHyFSphj/HtdV3A
XYsKJsWeFn4h14+QZYgrhivhOY4V42haVuN2vcMqA61VS3rdWWiovLrBf8vo
O3S6tbuoPJDtIbQXsfw1NwbBbIxnLNkepF4L6eyYMfCVhuUy7KfhvL/bx43n
vSt3rqTKCyUdEYH1UjK5Qd8DOgLtOQVf36fMdXYGuYUbuv2RV58PNjQY2unf
QKpM74c4YXtJtT8yLyWm2/uva+AB2aRErRaAFcEbOnlYHBXExcBJUNV8vPdg
yxwh7L6695e3BF6m2mpsNR5terbo2LNuNbw8KOSc1Cv7rOf2w14UF2zK2aR4
sdgVCbaI8V2OV6GmwdUmQ7whKeyIUJ8YQsRsCYJUXAWd47m9XPgnYosNXpO3
nj/VA/ik4/GStYJ8JJO4/4yAGobCVHuhrYy7VAiEyfHmkPLsmgHEwJt8O4cA
FaL3xxhUUDiAYHSdg12w7UUmpUHOJQJpeknnlu4hPuP9q0yg+Q4kLRNjhDnG
8XOChKcKapULW8scjMQwcQst3jnHzLJ1ud9I8TaDKg99bnDjLhCVzpWJfPS0
qlwI3saEHcP96LuMZcWJ1PRrPZscH5a+KXIZLXuWzcSoPFL//nQ9IU9I2ceZ
MElsaJ0f5JBZUS3mEQDLe978vUn5MZyI3FUr5+4nytHO/UhVr41K0sPKJYGn
EUQO1fcAdLznJ0omyC6W8BydDDROR6PjMPVgvCGK8jHTCfCbYzWlrVfzo4A+
sWF01thkVrbByQioGcMsRtNZtNn29k+08vVjUWLOWxWLqxXVGvedji2Yqqha
3BxJpex/evMDXAYUjgyyT52zvQ2VUlTw+aYKvhKX9PEtDsXpEGyRtKHydMu+
Dz7Jw48vJODxxmIqKL4uAwW6WrkjYqzzOvU2d5rw8DAI1WtyQm68Z5KvZScQ
U6LkArAQVR9HufLRgH/Q8M9lwg4KjjP+Rga5vlej2PRRIfM0FYYK0KKvmPWS
OvNxp/+9MpUgTlB6lm/AdpuB99coQJkYddWP3sokQ1kjOqFA2S00s3zxkBBr
0XfXhFhAJhgPPcl6PgVuCgrVQfBNgcBpN5KP3mFSmW/jTyOuVFlJCqb65Ik0
ZxZc7eMMj8zbbFWGiKFJSXtfoKtZqP6vNrAH0J/mwoip+JgC7szDzoMZwjHU
4UMMHjYoSju2zvXDcA3a6MuELp160CBd8R4/q8hnRv3UCIivI3Pg02Ff/pYe
bmdZmEUV0DCVmOKJyzMpfMr8miJhTg/G7gf1GOc+ihP0lmPItB17h3RkSaIB
y3RS1M77P3h+Bp0sxwwjAcvi7ZkMQVjVfNRi9kho2GFDbGK9rthoQflZBJRo
YQtabG8ZUzQlUjWexVAHRM7uSqseVOUH5F/pFi9GgojuqD2RwUVX2CC/8yzP
MqCwSbh35tFTTgy2vJngQZYn1qAZXWIiQibzJO9in6Ons3mxlEOtL2t4clJr
r9+Of/yBIQsQKpwvLdwPDIUqZr3S+EyF/9lmuxeU5ZSZ5PUzclGKYfeI+sLR
wX5EO6RPviRvLiTVg7cOkCZ+Iz4Of/IMc18VCvVhVcCT6PWBhIxE4LO3l9bw
CFg3ovl7FFZArQgYhG0l9tl5EFf3dn1uczmikx9dxRNagY3uHCElNVk3L40n
/+LBuRqqn2VU1mBC7qS7MfzkT3Hv2xMXUK6YUPtDLpYHa55tyldS7DT+a5G0
4gfCrkOb+MlNmByAGrKErqvmrDrlBjtfB8N7EzpEP3IQY1l3+9f07JhbhCZc
TJgA4DxUzmdizHg4vRTn2pvSzPQUDEm11ipdIZ1rtuUUX+dr9lfoAG9lBfvP
IwzUDAL+8w6Bg8CaABEk7nb7NsrGdgBCFDMs9PBAFF8Xb1dIMtwDhooeJx+s
Gz2pIUhHhd2qsTWb1UKrc6zzji7uaNOZNc5bBrii3ddGb09ZbkAt9fyqaJ3p
gfTmEBsDF0tVgBGrGZVEQuIy4/uOhpTa2RuLQ47QmcUYGfG8o/dzce4qznx0
1zpFD94vQXLzEm/Mw3xtMUegd9EC7iLtSuw2/vvS7Pri9LvPgO5sZoFaRP2D
bJfIZapxFejy9hDzO5g7t+5PpKJRovVKP5kNpPmWbX1WXx5b863vtt0TkH2/
4ez1sIOqw0D0DK4vv0jYgVplrLVcZdAk3b+J5DZgKtBvM5qET6G3tf50o9Di
X2yMzJhaUB0NVlkqEKhBnKiXaCwTGk5/t/RtPKFYqLK4DKZfIrOTwRu8Ah+n
ZkmUeA8DuxkadBqzd86B5wEOgdYEJ18IUAzfPbGNyRBLLPwUU7BjNcECLiTH
Z2LmsaeGdZFpeC/nkaxXzR5YrMvbfcMoOhlKqq7VW94M3/palA/E/GFIgCAd
QwqgCqcWOqjKPYW80BozjBc2xWtZQAK3J/KaV7oMg9u5pLo5Q51dfpTUIK79
T/LJt2UmW1drecF1A7PUeLF9B6qfcBB0Hs5CSQZdDIb4yGBZy3cb2y3o95y5
MEUhGFLIrtH0Up0F5wqclsKVy3Hizp3VxYlLVU/2xJd4Fx0mZrDZXen9r+RO
GfTJnG23Dcb8QSdHzihIMVog8TQtls67RYQeX1TcR9GPYmMo3VOUPvAXsOs6
/QFevZfygFol2ho0VYPKvHGCYNpW0DVO9xiOwSgK+itboGwYcI5ISNiawJ/P
jzE72ezC4vAPhBWdtV7j4L+u9L+mWsUkOgs+2x/Tcltk7Ue4SSvrbJ+1jTLR
RthLvg5szfwy/mjZgPX5HoS5jc5MDF1zKtOXFS4q3gpA3keLvXoejb0+myXf
sEfagvVvI9lOySpsEgoVnu5up+XO4UQMMkUHcOxTLB4pMFpAzo8sheh4R2sY
YUQe/+VB5ET9oHVUk4ouYcOJpgOSSc9+7kEODy3jBFqayzN2AEC2GT2gNTjo
fBEfZ8nRDQx3trx2QH90+uY48qLmi8l0B//1KVehZC3wSNz2w9re60i4WFMN
mZIqf1HJIECcsoBnoyCyHQ1GH5UOMB5jUrKi4ce0yCaQSgh9x8yvVxZ0VcNa
RCPXC2zBvHKdRQZx89XQurYB5ND/4+mjAmkV4IMmPvDVVcMpZWfKd6zMzOI3
r/oJ0aSiwyrWasgLmfxahPS2q3Wv10e7ctx1HPzem0caAtnkWEwK6qlapdUy
4NdmrnWR5xaUv5GrlFLGDeMdrcqxZ1QPfX/M5uSbLWq1YNFYk6juq8NM+Eei
IlrKShRwg3fmhD0yp2QPajA34Oix4k4lNnENYSNHMIgSO//aVY8mowukoRKN
CweGP8bvjPwUTCIMidlJVC7ibmP76FlbW7PAf8cGC6Kx648Z2dQlvPRg5ZmQ
y5m1ZEFAQRdLc44ZPYaqLLRzg8BpNkhY+IOWEsguIkAsXLW1PKigUstHRh4D
OrK+81+R5jbH3CVbnUfLk8CPwoO7G1eYq2KxZ+JRvpQo00mgwhS6UIVRvZcg
DujAD3czWI17L51hmVdKmVMX3OA+4zDKBFMafFNfrXOiFTUwleuAVQiA23U3
o2aengAnI4Gu62w3EMlGur5ibokMOGDf0sIY6/DkvZCamDD1SM76qdlrRsdw
nJceYNSTnAWXQYqJo+JtTZ2CNrH9lsjw+XW/CjvCi2sFHnLh7FNrgEU0xoh6
NXDWB4P5HtZRtfbwrWkUU09LVwIBgZdFIhj6ieTzlFfkD1F6OeGZqvCsMn8n
Aa6PzWpG0F6fCt/iydIFKZDwlxajSlzVLz1tKcAvuKAZ6V8/2U1USZWyJ3Mq
bzLKFo1DndwrQLb9ZSp9kT4Wvkky+p6qmGqet/ZsS/lVmCzEOAuZp06Hmv5J
5G4b72Lb74XIbv6fentEXvmsaZ7BjXWPqmcaTAlJCl7ruht6UwtDsRWvdwTz
EsoXFY9OznH/vS+5CAva/jVoDXHH7K1ZAtwRTTY47rswp1uIjXfmkg6Wwfr8
FU9pXclk3k5OVvMw8LofDpAhHoH9QM5JtMSrfkVKS2zpBD72N/YNmYYUSd/c
zGtfryjvwJt9LS3FNC9vLkWelryxcOhbRd0VDHh8HwH8m9RGs6CQs4uPVpAD
POmnImbhtRUe1EuLwbq0h+2wxgSZM7QPJvgqv2ydH0Isep9emNPNnytXCO3t
jtxlKzu/xsk6vAIgUo5A4Fp48p0iaHmOMv3mM+8BEwu2aba3XVymu6fdxcyO
mfGzWgWRNQB4YgHyO4ntSM+8sxyT8Y9MdTlwZDpHxAcckeLODtN8mAve/ILj
BjFY7rokN7zpI8Mp228fQhDRyHJK3ao+F++vg53mMqlQ2qGhv0HDqlIzDwmz
IB+fEuF1+faRJxHn2iBW2OK1TQ+YUuss4hzINITb5yO+M+GiJQbuem+o2/3e
pGvVUMaX11Ak7W/bQxAq1xD+vmWgD6G6A+smSfJDDvK9Qz7jS/38VBy6JtJW
2xV4upx5FEsH1OnS+gG7dgkA2KotsWVjuCuNE3JGL7/kGnfq9VESZ16JVVLx
CKihZ5TGTWSiRFbTqBuzzylk1unStKiuzdsPsUK7QKZA6eFNJlwY4FX9sbCL
aCsLYl8mKLNEXUJisYo4SN9OlPKevC6m7sU7nWn/B1vTEzvc5uhQoiQo09xH
ivh3PLPtyTOjEK/2lG7BBZZ9Gea8emOEAI1/QxRcortFtHCMLroZtI35WTqe
DaRLqr2OtOo8nDHK4ZULOQ/4NvDcRqrEXt3odkgI7HuDbFTgQZQqAdgMgHeQ
zvdkn2RW46dX0VjD9RncEHMZuGP0bZ1SfgK4jpFfhACMa70XnK7DOFoLGL0R
r/n/pJLT9YK11T3sX9gf6RCKdu2CfbYvmrgKmvbFvtRtbAJu40rxpAZrBGz8
QrJJGCfFNlGlP+MmoOXkbdBLZKvrlvxheVm/yI+lBoFOp5bsYv8S

`pragma protect end_protected
