`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
qxwrmuxaABpD0BumOEg5bIFd8rmfflCzHzjJ8AKp8UL3z4Wr7Evk0ZbH89PchksV
v+ECLSgJDLPFLY3eSvLg5kaeF7z3jCNzIwuzrhld1alY/jYbB/pIpfAz9riGtoLA
f3l8rTOAxsu4wpoy7kic2zBplmzUEIrRW1vj8EopH80=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 10640), data_block
UC6cgVmBGUZ7YRe7ebClL6QIrFQGe3oA0dmXb120CfPRpVNAFn9mCtVNMF5JaXMK
Q4CRaUYStxQl/rsAPKgX7x2qNByfpqDO98J2R1HUhzYyOBTJa498xbuQIU6sUGLq
jMdvQR3fLkz1zRaGV7d0s0x9RCAJdv5hfGyYsR1NfV7GS8ZfbelnHpPbXnqCvHaU
PlEOavaZSMpXNtkFdxLrq4v+V5WD7Iqb7e7ptjItanFIooLf2ExlJHXoxBecsov3
IkJ6zjOhIUT5fhjdkziA/8rIja4WU25qK67Ll3jHcA0mNmHoQ2ZLru9o9geskM6c
uk1lnDQEh8gWHK3p3yPxusmrNcoSZObDIA21hhp8iAOv1AOPZpGFPCoBwAa/JIa7
MdPC2KB0tV+VEOL+PN3V/hTxLMaRgdJz7hmzlQk5PJZ7TyJ5kivKlSDEViT87Kqm
jIP/6mAvylEejXsF/I1XboQHri9W98yOTsNQwMA+W7xVRFlQJwz886VPiELZ3Ydc
k+S/ij4Z8WXFMBoiga1Z4R3ZLIW9bUqfbzOuXGmwXcbkoKVdgF3pLwafBhm6JUli
WVYn2zXcJfAR0Pvsx6wtj0Cud7Rw+RvhNAjya6+IUadq1b9tHCeX6RQOQlnLl/ZH
fCIDIl5EyUatFh3YyeusZ9vjK4fhgcK18SjWSg0oro+lbercv+mJIZP2lW2n5Pqq
84/E7SHML3aFLa6FnZprEG9EOEUzOPwmK3Rr9DWhIGhoUaKAwfBTrwQsSnDSd5KH
mvuqcS4KxPxeuvx3TcRHiJhtqBRfxi/OVZJX1YMrjBMqr1GoazYNIcnyxbwX9kyB
qwJqGY5exQ682xJen+q6qsCQ/aqsZH5RQ+ygTf01wehrNYaiVBN2oGzdpm3CjEev
SRtqImT+T2gFfA8FGE6jRMp1drak2kXdZaSnKeibh4ZBH5xkc+A+LyYe54/ZupEh
g2hvA3D0AC2Ff6efYaafHVR1O1depnjXpUFVy7p5IXloq+Dsm3Exn8/6cplrRqrk
3XwWErJ1pWrGECezKLjxCfnY7ESTRx5L78cnpe/M5opiq2WxSd0z1M+2hj0wAYvN
3rxdJ2zLdEQ9VyrcCWxbz3KYolLmpmSlja2Mvk6RZvLQ2PcbJZjfDl8B2czSLT0R
kfY27hRsfO0Zcv/EqLfEWVINyeaHSrb+3YFEIGlmcPHoM5SxwjL9Oi/y+dcEpdzu
pNmebICda3EakRT+UVDFCOYwCqaC46tSW6POv/QvHkXGeZf0RD/F94zT/MMScIOP
dfOmGeRnuwhEXCgJO7Z2k5txjewBQD0yrmjIlPRzpJ5MpkT42LLR7lNpvycWW713
5dbu5eRb03wigGEkcDVGoTV9oq4s4CbvYvV6w3pGhZhaWQldWPq5iqlGLYktu5jA
RVX3LzJ9wIsCwn/gjj0Z1zG6LdZ02I03i/RW/iGJdkP15Q7BAZ54qbtQeG8o8uyd
eADSKOn4M91N3fVM434BNrci5kf0pQ97BceP3bEYAq8f4pwMaYxbhbGeZJy2mjnz
Ljz+DLc+w/EhoUxrj6V5Lho1PTLjRXAM7OTje6N/dio/73xmPdj1h6E8B+bwrfoI
oRu9sJPYoZePR3lKqMssobHXHJc1uHOGg8nf0NX3zR2qBDQl7L5XSvtVmplciGAN
MDK+tnOkfoepHbUTjlW4afDFJjnRgCjtgAoJc3c1ga2FoUQGy1T9Gau2uPLxWFaf
wglRA0KdUX88nEuCASsUSQoXBBMWfXjsSocoqZEEgaPj76Kgk2EwtAUkaQFXrI/+
4rVPpbO9gE3WxLDry9tKqliWyKtLDf3kQ5xpv212HCoRx6AsyTnTXugxaPduO2aU
+0JYQRuSfMGI+NVEeK1ALN+VyHFILTIK8DtQsvSs5IjjhYvElhcBJSXhTkTMX12E
W+Qs6v2OnyWTYyaxFOlDhTIxnUCA46a4ConvkkFFMosf/aSk/3i0G3IdwOj5T+Jk
Zd6LhXMLXu+ipkw9oAMq9btHSPB/JB9raPKljRsr/QMAYXHtxLmQrj2ycXi/Ilgg
YUKLT9DH1SwU9dt9u/85hqBwLm3dV16Zd4MrfG2O1QtdNfkfRmWgtqGowrYYlmFK
FJNiTCESC0ObdSvWnAXlXZnV40CATFM3w3bNLE9MFvx1vAqMx/bRVjNxk9ZocrNu
vatIRpaxZzKBHuyLTrBI4dcqyiBwvJm4fTU6V8DnRVMO6+r6xKX/675Xj1MInXAz
NacaQp1BYgPjpVQg+e4iu2nS5Ly7pheV9gt1o3yyambgC8Zf+xDk5nSgYPgAefnX
NJL8pBNeFF4ji4+TCcipn4+5/OcNTRiN09V4BcvQ+1tWd+7Cg7zeALp3zg2HJD7N
YHsPoLOEQaIrD2ljoOPP/HyxiZ3r4+LQITVZmDwwkzPC8UbBVfLFAq1ZKnnrZGgU
zgj7e5j+LINcrTD6x/qURBvfoMaW6OKUJvoD7wg0Hr/LavH4318wezsSX+04GaUD
JyKaBCjkeICz52eb/3JPvDc4Mh1lT8ZeA5tkSMS27XkIOgRhpmglLa5p4Hl7cY8O
f5zC6fDuEJJ/ydLo18Ed4cxsI1NmMVPDwmp7dbOI8NxLYYDg6ca9F9Fqan6YGpsB
lq38pKyJQGu+ziYmbnsk4qbOsuvtQuscsZxBKI3ZTv/sdOGPNUx4LH6gphSiwTov
ZGE1ktM6ioeD5iP3jrUVX/WO5X5hygHORPoBNoZu66qjwf+poqqazH/zPJkx5H3D
jf7BljvSiJryhIHJswgTy1yisM7ALX5ZdN8RMaDRaaPg9mjv4R7qtGjrpcW1FXIY
ln/ajEIu2qWJuoO6n7PkWAOaDFxJKrmuJjL+5rS7LHLNiKj7iTQlBnByvocX8td8
n5eD7tqG8J3GkBODa/bSxX12aHqrJkckvhbFQF6YIM67VhxLlYuPyr5JR44T0Uej
S3/UnQbUaqZV89KkEnSomsoICrt/wQnOK7+vJDtqgI7ln23mBz0PeFNILNuCBUPQ
aoTkP7wWJHOEy4zydKoivLrrWrIRwWcbg9vtBnE8qx2FWwpMQnsV0hZRHk3Pu7Ys
5PYep8EehVJbJE9Y434vIOgOG8ZMdxBCcflbZNqMyWRfLiQx5BE4LakVeIONs3s7
A19IaL88eVqV9mYFOX073AfG7Sl8jA7khmbojTxb9EQO8Wk9KHa5t5gBbCHqYRuh
aGDonNoazC8+rZ5ETQX566aXWZpHcFUJuZj/33S6oKsqFss3gctsStlej7XYHmU0
i/9VZAqwXwrX5V4SlkvF5pmAtvGSksMPBraCztYbFZeBAK+qwrgXgCI6yUiDvCfp
RmsKsdVW2WL3Gr1tuC243nB13UXygqhXTFS53PQbPr6k/0kOkVlPfGd+8gr9OvjH
q4ArvMZ0DU289WXrIwr31qhCW3gSAM9GNIedkGozSZwnll+jmmTM7sTKHTLCvBnV
4H4viBfW/T3oy/vTyKs7kscX/5XVyuFqESIt3KnPA+YUX+si8Qv7lgV7wjHk0YOT
k0T/vra9uHvSo85FJUdj5UGwEJK/u0KAfLUGSNbXia/n7Wx8GJu050jKtjicjLwW
EmJsLjtdoDpay0oWzlDVucUxvLCk2a/NHgbt7VYvo1KkUys3J4XAwvucRmcDju2r
Ch7LQTEgR7xn3xaB29Rb36WuSXuPw+sNMaf5Z/0maOwN0lisVPjCaCLHK9ATphT6
SlhC+0iLRCAnwZtGi7RfqhVGGsqXUYritqKLRM1PmQ/nu1xrZ15BTT0IZG/Q+8U7
e3xiRvVm8p6fFmIeUMFC6RAtV5tilQZ1o6VUGaknZYpb9zheGtdpOdU9PVIRecpW
KHcVpeQcEwnTsDstwi7VZHL4HzOWfeI8vrWHux1ewLgYNZCesQKh0wEffFq1Csst
NMicI0HFJi3tr6bwFjXVW5zy4IpD91gDqHrXMaF8mgPMKcIUNhUhrFAPErgcACC6
2NzfUbw0yifrkUm9Qg5ygLZft85GZ0Pz2D2k8wW7A4cILop4lxqDbP5+tLdqbQfm
LLXbxPYC+OK99jKq65X+F5pMkIi7M7pRmEdUcv4xi1H6MWjmPp7JyYsJh8rzJBIj
RO8bDrhvEJfdrrRgmHS4PkgfN6TwQh47XWOHOMhk2x3wvG3GzmI81pQ6A/1TiSDv
jgcAzFG7Lo3T1nbXrXyzHlQOtFIK2X34VDE2nvNudlUqe3oHBrfaPOsNl5BmOukv
oJTkPiOoWaWCORP4U2zbXhNmq0ctAAwfH8wtoniHoqkQx3M1Ox/7wkFD9Fho207s
Yj5aZNRrz9/o+uIwpLQ6HiaZT0eW+wW7N5AtTrSqLZdUkSeJPNFs9Ay4XOhi9Gck
8XzPa9SpOWi2dU/zJYtFqwKeASRXvbswGrvv6JEU6qZqnsNQjjungrVraekbwlvN
sqnIcMRTkLmewTQm+l6K5fuCtdU6m3IgtwF+jlsTFXNnFF7//vakZTsz2HfSCMpi
CP7ks5XTYKSYbEqEKW1IK8BOX1YNQkJjkTQRsLIwjAKkJ60SBxlyisH6HX9B1zzg
Ayd2yPtSbzQ6xwZFD9fmcgbPX58vUddbeP3qh6w/bIGDF9NfmfUGEPqs9XOaJX2Y
yqtjW52ImIYWwxe1BmnL/X+F9hz/tRVcRmBdoqfnX3NKQnTohBYS2ep83TGE93Vl
nh06BUxg4pujUnsosAqZ1LcNZZTQpi8F4l888p+hZBIAPCI19zJQwyJ57IHhGwRM
jwSUZlGxdSJxsEwWfy/nw/5a6vKqIZVFX3wujhKfjjFoeZCB6+DtfIC01QO3joSx
jlpuIqlavznj9EMgGxKjSmkTjH9DS3pkBHBm7NQRP+NOePE1aHtOFOtNct9jdBOZ
SvLCLjaYix8EDqGtB/+UaSOMboQw4AanF62dnnMwiq+p+btS1dTUZixMVjJGTpix
fAnOWLJwhV/1ex2uYuqmb+ir0MZwvGVyDLkdGeyIx9Ktx9Te5mjLZ7jlCITIwXjw
WzSOTxn6Hjft3o/QTu8usYg/zKq+VweqF6YofAV2w6wjjY8bRGvgnyNppMI8ewhr
zQLezIu57C1aIKfSiPQp/pUHG1FjYVaI9U3mVGdQzHgdIQXwRmuATkzJAI3tJXqc
pi4eN04lSdgqWM98W3E7ToN9hbwmHkm7hcmkx2Lp20sPb9uyLBWc7IiHOby0vicQ
fYAvThbE+mpiTGPJq0bL7ZZjlMrmQyjrM9tfgGrUO9KXD2pdkTqcT23VP9LmyiHx
1i/q4aBoPUITSQ/5hzNznXNpV9SIh1yjdFYbi1CVRlO0RfJx24SapuAjoQuyO9DQ
dmBqSeh2FEow+ml/ZIHBEVUsooyptxMZv2gGEniDxnf4HSERxFY6NUKgAlu9rbsH
1V3G10h8YTrTnhNUTK1CYfcqmK+83oXLXBCCci5yHqLyiWr9LdqjoGCrlQw5e2I0
n9+jEGaXOMqmEtIyGII09o8z1bnYQdttxMvtjI3b5mUCImrl5vcbyWtPmEhgruww
hUZ7L1Hj87dpd3mTnugIic4f98lpL2cqzBlc7J8wL9MYNM1LP6EMeIB1Ow5vN/ro
9SnVmDmsXh7QRbhIRa4af0RM8XKv+5GEzxTf9brrq0mk0gNK9L6MiKqW0Msy+r3u
vlLXAsS8Uq9wdc5fEg6TQs9LioMbzAibNvZP3x1lskWZYOqj8yMGtEB4lMZaIMIA
8iaZC47imliCJTySy72qRNI288r6HZxsaoQoSp+WGZUHJDDvUNHS/QD5PsXa09l3
+BUOYM9G8OgiA592cttlpyMEkCIJLNOnf1Ls94UlsSHYRgHZbVr1/W/7LKsVVa7F
ed1RlDuO4KgeN4s/cMIlVH/NjSElFfZkU/0lIYdVkv/c10o0IMj+TFxty3otIzo7
ce3p1B9dVJIp5/qii8gEUNVwTx67fezGoWDf7P0ieCcDt/sdkl0upIraNqz0x5mJ
1/deHLnYMiQ5GlKKdJKN18rJNk6ZiMMehLRx8g0t8tTEcDz+sfaSmUFxKOFDpVc2
jgZ6pATE/zFBnqVvfgQTrGyQQFUr4hA49U414MIlawVLmcr/DmdOr9EszQUvx5Mh
jkCB7Mft1L+c3j3EIjXMVzutRalKOJfRFLZivKdgZvu722XIFLZPWfT2vhmgdnot
bnS0eEdg9vaYgQrlEr7bec7kiB/o5KveKb9LLp1KQrifDTX0On/gMTPBilOuRh6d
ZQiUTQ1KokQ4yhJm/SsiDtbl8IwgQxRVKPojOP/50FmGj5U4LfHfFcXGxvLC8ZuY
cNYdk78HedOUxrm6FRUAybngyrlmu6OOm60iPxggNM5xw5rkI2nWhn59WUtR279q
Prd7Oeyy/qb3xLtcNqfBTZuu8yp8zkaQDyuBp0x4Di28ETkabHXdhLS+joT6y0Ha
Nq3eghqQQU8FoWFgEiRIQ6j1qgF6B12IWDtGcBL9FY81Ep6Uk3+0Jb/DYlFxfKHn
swG1754h5q6DKBmzUoLo3OVxu6fZOvwY57l1OXn6rcbDL66zHnpmjDACjWvmuGvi
II14Nc1lwzmWPHnx/k3xwKmCVjhxfRMMuXFVqcnF5REIItk8i0nGWYkT+/eqm4cj
GEOCCFsQnsI4NpvsD4j/kOekJp90O4X7m0VN9jRdfF/aSrlRFOwlupM0TP6bvLrf
JeqS2lX37eLLW4vvyQlrwnZ1321oA/Ksgdn/Otn0dLcSAmQ/mqqogrIpih0aV2Fs
Zi1ksi6ST3mkX1BeGI7QtpO02WOkLDVX+rJAiUdVlAVJdWn1bCAZa3YxvaSzCqbC
gl/Yy9fyTeYEpkklhcIhp1ZCaK3oc+mr55sVSlVpKjhQQ1gJVOM99z3/65qtiUmM
959/ysj8ATDWSiDwsffYsEXISWTYHl3bEj5k1ObIN0Gj57oIKNl0tpJs36k/OM6u
utqf4JUIJX9d4yYJf8J1ggFi2gCuJMNK5kAXA8nPEIqRac9g+NFOkkuVUInaL2I0
Q5eeWAdDslixNrAmpt0e5xpJ3Cb+bLMJCfhKzjrzAIjmeLuPCx0I6MIP0w1CTcwv
jugsx+CgWICKoXTGwsj+snaow0ybdBQLSl7JKu4TzOQmMwot8eESCP3BGWxbR05L
Jwck80hHCsN5lQZHzCUPh9J+UYizL/qQdVNngnpjqQaAofDsdOJrk7axKZuIvV0I
wvpBiMlqoftefJO0J0K8zR/aojRegd0mRSFHDaR85BS6gx8nSSQACyQumhFwQEOA
ElDQY3mQlc3fgX2GgjYp8lTpMfhQuiUPrWkOpJcvoNuUDMhYiQQEe95f4EK0PnV+
TVH+RMLmkVIntsn0T3sQptMfzuy5fj8xNvwO26uPFucFnnN9YDQu8/rnNZXTXyfv
fCEpMtJC29ycmuBIbF6SEzuLqyzKSEjCSQoLfebUv6pFQMIWzqb6OkzQ3uZbVYz0
gkJpN+ZkptrfNLe/mDDiYcoTErybZyH6k3c3iG5lfKVcsKGbRtqYKEfy/WmxNw9S
5TxbAAkXPND6WXN5uAGrYTNCs7lpfttaCpPKYUMDuN3M6yXRqMcg39jzjfm+uqaX
6uZSmvHYTKSsLNi6Jw+XztOsGMA2YQ66CD0QQlpI4Br0NH4LKlo1YPQihBvBXOx0
7r0U4QRn450usrurN9s/F7ZhFeJf9SRrI/3SiX2QHS3FMbO4EVU+MDs6lU5T38Ow
SQf7o/U6YQ4lFhYEVB03R0tOMvAIxzFpO0UThRPCRCZ+d/X3hLvXkXi3kyX2dbEf
ZNhDpWwjhZUuxBk+TZOOHtI56Lg10BNrqA6nIMri84ZB12wueBOvAqiCETzyd6TZ
HJoWk7KPVwgPo9c5UXKsVMi+c3sqyvT8sn2oeDAA06KP5YKmvH2sq/XpN1vmhROK
icEbipc/RaSt1YJ0ByYZPJGNEiWgKDNNcVO+F0z9YPlE0kcOuQp8NFxuamb4IQ0J
/L4ZWd7j5/Aur3TpncrqzK0axneC9iN/1TiwabeSpY73RdMXcUre3ztlBsSExwFF
s+ZEqGUezfKv7ySzyCdLDef6fUfGMUtZ03uK1mmHBHMFEikf43yzk7hB6iVw3WVp
6PfaxmLVldXkCXaLieLrzgunjooJxUuC3JJSu+oegni7eXYj3YcQEp/NIrT5iU+T
4lTTR4ThYbfnSXwl2dBHiP3bzms6UKLqGoKZe2yKxFSvoVn1f9Nzdb79BoQb/cWK
UOBteG5YPLVpw7s5mPRWxNp43jJEaxB+gqDmBiRkc7K67PG0TRkaLjTIQc0vkXd5
NnbIcz7WB/+7J+L/g9QsoB1ah5gj2+fDbSN4sWLjM9W6ahNTtGgE8ylzW1dms+Se
UmDnJbfL2itZPJfq0Y+8m/oJQAE4qn3qPCCgf4olorUSzlheHLOBBZhSKWwVQbt7
5ToWVrF0Nwc2NxjuLrqZC7eWE5JcFfb2d4DazYdeUp+nI4Zc1jn7Zj4hlhZEvtI/
tiK5zR/uDrv057okblj6OwNeDJhaOWZKTrJ9YNCrdt0ohAv5PzYKPrapH/kx9CBD
T1qXQEbS8z4SrChMRSOkaV81QRP560GWj+YWcdIwuxfVgTk38xEFqeKvSgol4Uaf
QhTYH2GyRjqp+QOtbnZrngKC5BpXzLOECogA0fp9RzSQf4zAiiMCF9haVI+Ie4D0
E1u2RIrelP85WcJu1l7a8bIygQ2w3t5SzoIxg6vESLexqWec2ZZ+n6yQfC1yDZTh
ZjPmeJYSAh2ypIcH5xKbnt6jJi1FsysZnj6zPTfSerjDYdNUgTQC/64rt7kCOSWY
Ombv5JQXVlnQ/abAAgyMrba7bJJSX2rhJBtQpf+PryIirnhlUao6rK9ps1lQtBCC
y+Q7YBEmwPMnD2Wj0SeCcGddxcMlYFBxwNnbnu6l015M4ni2+2KvcBzZFwT7kI70
jdERuU8LuTQ39si4/wlLGvoIRsX+5+DOKU103Ny7PCBW8Zu3keZWxyijHCez9NMR
qmxoAS4kyHUYJo/UdeeaUGJtQo4U6ssHXKHU1B2D09HLK6FGXXM2cLmD+NCeXa1V
VyM/iC2E26k16C2xk4NUc3XvHjkHnklI8NEznDWCjx+GtwfK7ng+gnExFvqYx3s3
Y+ALVnEMAvIpot7WRm24XLwqF/2RlyeCD++WWl5/PTHYh31pXDY6hRQlDM6+5S4U
xdQsn9RcqOQXZZxS5x7ODjQOOhA80mQLCvJZFjrG6jlQLH4ku0KjfSpdnQ1pFoJi
8b8qbddq5e9MjjUStmVBtOM8MLZnICDZK8N5FUgQRImhHzZijKUxPHuGIkYVY/Le
n6/U/fwWA+JDxqgKJP5CfSuFBLUwZwSK4Eq8tz3m3IcYQhh2X1bDfEbGdn1p1s8b
fzHxADuzPMa4/UuvotvPcaNcsjSsQyDfRRT4+fK/uibzGRzeIaEbMzWHQ5CTInY3
sbwIgYNVb+/2V/SW7hOZOu6MVkOL6KAYC5hABoL9sLuEEAnT0rxXtoart1RaPa4E
PFREw4hHqYBoqsSaCHYo16NwsU8Au68qCCb9rhzLAuIZCA+6Zj4SxpJk0mg0fQSA
7FXxf9Xdzrvl20D+VFm+/YltDJWJgKxwq6go5UseL3gJ1rJXlTcuMLwYH/UeXeBV
EwzrmjGDdIzVSLQTVSiRo6Np77NQpAHORMTBLfJNm1Cfm56WB+AZjuPKNs389GMZ
7Jv4mBJ/rt+qqxvSUvqvZOUSRNoxdeGK7KLzEY0ppoSsaeje1qTpcj8HWbA26bD2
yw1VnA7R1TPsXcbi6p/7jKTVxKCwqmR0EqBLBXUxkwR7BavIM/JED3ot5DGBZakJ
g9c/OK+3sIrZ9AxeXocRaWTkQpMTss+YzJAS7ZG7ZBieZuX3cLBhLyKOzxmheALa
xj5CUO3q4ZlQIZ31J/C5cNR9pgJSZlQt3qpY++partwk3np7l3cySMVjyEw4DqZc
gNbRsY2jOh99kd4a7SEfEq3R9U//brWLueZQBviK17gGilsIcWXjUCk0onWnJ0fv
5zpOplEzJFm1vf3sQXRIJkm5jzggZIxei0hEx71YmvUE8u3N2cnBL0uEnYdimBX7
hN/RQAoe1RGvfl4MdkTkFYtnET/P7FHNJv6WoSgb8QIYBC64t0ky0vmO5cW40uBd
uXp3ribc5MvL+/qa3xLWvUWOOxZqFI4Ygnf94AJ4jJpKf9s64wsv5C8ROZA1OVNm
3SWUJv15KXZ+IwcrU79TrwJXhdxU+2jMEAcuPH7ZFy3GafNwpMzbb50OzCGMBPCA
hpQcaksIhFP3f8Mtwd6B827x2qdF+MHXRlXfdbmk++A2B6xcf7U97ItHdlcpf+lr
+cA/jxemIu0/paHyJjJw3Lya7zWSOOtMeotoK5wqlCmo2Vmosgo95zlyec5L4u67
7m066efeQO/q60M6ItW5f9HWU0N/8c7FFKKeDqx3xcH1FgeVbrxP4AdUdjybCO2f
ZBLUDpJI/7g7E4hLHb69HEf1U/lCy3BKJ3Nhv5c71GaLvzMsl5FRl93DdPYkWW0E
x6Rs3OiCn9rYS8nkmCqxiOG6d3sV+YPX8Q5h57vlVjZKmZ8xr8e6xEbTmRPpV0HL
8ChzBdFngmoq4UlXQfa0RJ84f0FN++ZPdcwnhYFIm+7FyGD9YGg6DMWM1HfjWyuZ
5VZez8DzxenfIhY6rC49Ro7Qwg3tbVW4gEsedbAHG9vG152+oXd6xtO3u3zn2gXP
Zk0pMtJTaqVupYOKE4aRAxJ89u6sx90iVETJcb5+/0HotC0p5Y7iVXp8VQiX86zh
D2TQcaL6I7w+zEbbt5WoqFAwnC2VBRIA/ZDYogahSlh5KUnnfLDH24P00mpJ+yIN
m7bXM3qHzSVaqa0ODyGlSKJN8txXit56dKn9RY99hgxu/d4JmMSansBBMWZnNXto
gN3wbcyvZZqCn27k1+84YImj6u8EL10bWzrG50WaVzIivv1Rve3kTEi+aTVoeEu8
zpHDU/a0RdK78Tbz9vLrR1kL7B7p/Rbiu4enp7qMXBx+PiiU2icg/sNDmt/gQxWw
Q5ZSH8K1i+enJeeUzGrOILkzjzC6AGQ5tD99tJngQOoUQINTv/0UwSZZIpHbRnYj
Skil0YDLZC00FLpksfFgmo7JKHHJqSoQfU8oJ4lyyFMZAPanol4zn+29NPzzp+SP
uq4w9VNgUA/IASvS9Q/G6EI78UqFWrWqNeC6RV4J1JZT6Ycod09Rn+uLEcy6xsTD
8kmP6y+aCnwgnmIdG6cz+Q3e6p+2mKLF5/9MyjySL0mOibj+EloxxM8omPTmoT3n
lXv7b5rwXNfvrTbiDr5xKfhIfD7eeYmLHHDq6VNOjhsVOIZG5NGD/soI8Jx+yQ7J
OwBySTsnispAkI8smQiMQxTwhHt9iUTuzQFTeTFC77eHEHc9aApJNYYfujKfEUWY
KwBH7u7/pWRLhYgig/5lzT4LmjccX9cADEOZhwD0btQEmJBo3SqFNK9SOVGpXRAY
y8iI7v7k2DPc0qqnCh9r2/DQBVgIlrc/GUKtO90c/H7QpiTQHPgVFmOJ+Tw/JtU+
1S7bNEfN/XVzwqN9y9m2/jTBk5KR02HXTUnhA5CSpvcz5k6mnsPiBfsYhKJYEFsJ
y6p+8VUcUs5IZTA5Tm1JbC2PVyMlHpmzeVzfOpXydvF0NcYlQkZdFrDfk9rQuCwx
babu8F0Kh4qEVSUalfYf3uAco3RaGy0Ah6DNsdBu87xKySQP/sgJXgyT2b7xZD8R
cTinnzOsrM9xss+ww5VHzL3kmKp9wQazqomVHfv4e6UhQ/vZH0wdKYZUObo7baE8
UXzHOpE3aYKeqt0aHTGIeobO6kyPzW6SQukl5afxb1GToZRxc91hV8h52OmJP+Hk
jBW/kjxoUwEs2h4FDu7iVmR0iXqypMIYOEiAi+dWtoTK3H5e9HSAWNVf112HP0e3
e2Y0MuHSLk18g+P8ZVsE5jdi9CWrfKFi8mP7y3bOKZJR/Am3a1GR7yYXbySQmkrW
K0bK0lkvPSvQfToK29bT1ZYgSVljYzeQn9ezACvWKJGuoXdx27RcoOfzpDWxtEZo
fvRiZkyCl8mS81DddWGhVDLKvlm5be21M5LzctO5Hza31o11NLBu+6d883P8N2Yk
MNVi/jDzgCYhuXv9/U4Y07Eat67kuDMQnjJhusCnFTmvjuLSNw7+655Sur3x6M9k
22FbmcNaHXjEfbem4SsMUP60Lywa1sHdwoegVlPmd1zunrYBt15HcuR6HfqNhdDh
MjKybU2EinwDAxx6bx5pnvr6EpicgDJRV7zMopJh699T2oup5qwNtfZEZvn2IbE1
4p/7u+vaZxI9ui3CUjVLxmqpvjjXbK59NgVkm+AuI9DNyvZUpz17bGF3JvVdffma
wQI+1F1ySFi+4vUpaVY8YN5gCn/7E46QjJWhO2zKR6wHqd5HewVe1qDsNG9H+iqJ
o4HjU2B2b2m096QDZ/IbqMKbLAkP3kY49kK9CaKNe6uCJLc+f0hA1U01Lr20qhoW
CK71wInwU3IFzlmtSfqX7nbpOrNgBbuuuZO6MKg+dp322k0ciREK5cB26ipN+FN0
T/TqJdrdLC9Q9e9adGuadBLEccRKtK00Ia/B5tqdCLlp3rHLgcANBJdiaQ513Yq1
fyTi08gSOOvX4OsdUj9fPd7cO1MDyfmmUjgziB0z5Mh+WYYe1ovCMRkdFsbrVUkg
nKqXdcfbXjdD9mgNhTCnUtdLRgm/PEqeyeCxfGHEcddRR8cWKEBUIWnq+Azhv/w3
LP3KA68DOTFqGw3AAZdaDdXzYTo/NWI0nh+6C9Vzw7tayBoTJr4Dh7hNqwlH72iF
q8kWU8gbmp3TfJ6w6Puhssnbgbfn60jJIQTA0VuPMUKBGjcZr4scCkWTOZGhcXje
9VFyIld1u9523zpUNUGCbzn/nPzGwBdrsnj+lJyF+8LlW4gAN2LAwR/4kaQKWpDs
RGugYk8wTagvOrx3+Ym1GTcNW+ZjcKrdPmnxOXwYmGifmGOy24akw7gJvJVQlTpA
2NcwG8iqQ28cFzjqcgEJQrGhSKuDfI/OES8edfS9eq9T53P7ByQwx1EZ6Wa2mhb8
s9NLah0G3j7E42Sg1Pr/4BZ3aXbA84NLyBrgPqyrzR8Bi8CmOiDnIm3NYa7+xy76
X+BkBv3fR8U2MSNNa3CYOAcYOUrcJQ89P2lpYSCiaLPcNTYYAHJtJKNmiNWt3mks
xysnRV2MhCsvXDBbn+07vmVh9PAdhzyc5bCr5bKTzaW8j6jQYn0x+ABAEtc5uMrU
aHqrQbsCDRoebXAyTXfIX3VSB5ahFifTYFEflnKgteM2UoE7Kqs/d/YA6pf6LPwH
1Tn5gFTt+XvqwFALFqBXWwRurKD0PQu1EvqHADoyuVRDStYLLCUGZ1/bBaJdvfL8
Taow8wMhaiJ041pAh8SdyL+tJUBrWNPfwbVqLGqpwGMkbMaC2uASR+937PBpSug5
Ni7CleOfZezs3D2rh2d07TNS+g6MWk6cu8UoNoJGnbdmadoMl7AWq8pKUaLncahC
5M4rUXsGnEB5qCswFXLA2VCvhG/+pB2tffxXbPPjjmuEnRc51d0xS6oBfqZcW4cJ
9l9Taz55qL/qH3PLfZSPR8F7KkD8KR19HDqruZx3C+ON+aVMZ2mb6HBnDqBIv73D
Oo9APIpVloCaCPQ0dchUyMF4gD4MqwholoBxpSiecI7t8Q97RGk4GOD6rgL+BSha
AC5faYonc/8evEiXMCOaNTD83qbW7lZpFrnQKjIi6ZYDF9P5wwwSCPH6f30+w4jd
hg91Ce6eRjUPG0U/ikJ8P9ufyLu/UzxbXwOdYPQOmHwiAEYbyUoqD2hFrq5LZGwQ
sd3EXhUtwO7xkhAXkPED9bYpFTAUhM25IJndY4sNO/hEEPuT6sy8Y4Pgx8Ikf2JU
b8u8k9lVlB5q7ayUEhH3rmhj+lx07kFJ7q7FE3llkt3IL8zqfoldq0jSKVoQqCZk
U9SeJgnpDI2s+WW2lgokIVaPhPmW+X00gCRFGGa9wk0TpGd19PfaqC5HabSuetAi
CQew6Kp94jrHC1hlOr6ELDUo3z+4yp3UnupQqf59O1aiWqI7N8EiO3Ek+rqrj1ki
9665dpUI1of9T3ZAyl81Ezm0mWgFko736DSJ+e6bFGIouQDO8bAfvY7t6WKovo1A
KhpbMa313M3Vdrcdn6dQDCrvKKfB46s3mvuzMzcExwo=
`pragma protect end_protected
