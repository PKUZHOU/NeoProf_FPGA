// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
NrDkKYu/EvAd+SY64Hv4HAL5AKvBbdGNV+VHcJpDqe+lw7ORG3AdiRsuG23I3QVJTBCg1779YRiy
q+Hp+p/VGQ0PxdoRjQ+NFkhJNLax63Hjci2qrtXxFE7ONLlMxodMEzPrCHFPZGLgVo8iWsZoudj3
GCdGk7z0ucZJRSOqQ7DwjMI35VsjKdYgTKN4GkOG00RE5Ij99pT+P25QH3ijOYlvDo6U4cDgYOOG
zpsECwxUh7k6OvqGzRubroxe1pUYQvwH0m0d69RcHX2bZmVg76kmW0DR72Ya9jwGqg6gL8JXe8C7
Dsb7dHZI8G69I9KrSOpvffp65p/epWZp5/Y/8A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 50208)
oIHuFdSfgyslk7aEI3BL1iQ6pNaBv2KHgto1KiYIv/b8xCppMk9/9euaOsKnkH5X4yhT0SWsM8k6
v5odTLXJzvYxcoibS2v3e65tu2iP5Emsi8sRDWLeseEbNCtFVz7TXNprTWuww3MlV8jm9M4Dak3M
BeCOWpHUZX8kSOhDHH2rGf3C99UEpZYDg5AqihpLVyBp0hQ4lVw9qV9z+/a/SxM++nbXnc8/55Im
qAdu/1fhgm0j7loE3gitXQFxUcgWGZOt6NqQ2s69JUBz4DSpepm5zZLG9u+TVmO2/2RFoBRKoDGU
ZwP8HUuTucc4W9crIJHMrJDn9QFRdIPDBIdXH+na5EFAGKXLL4N+RiWVGxE0hwkiq0Gz4sUSn4bb
CQwkOnPUPnIKSMOdLpbqK4CJR8e3hT0YFbixLVmrub/UNWNR4g7mZYDlGmYG6yFI9qcmNgsTMNut
8yeSiyXnvQnDoOTBeHWOuJBqxe9vLG0u9W6LhiRxxpGY3PHi1oHs0rGxQIX7yXSwsqvslcCkcxmK
kHo/plcTrRoMyAkXL2YXXcXf9v63tRPmQ/7DYverMNYSgEybPC3jADy0s8gSJJ3gEeucu1aLlXsO
l0S/Azu28gwTNCTIMNUpoXdX5BMwzXihs65qEk/kRCFfEIlgULxkzL+lKQ4SM6VJbaOeWfIiP6Nc
2Jk0C2sgtM9HpwLMj8aEJx3RcqZh34rQGHu+IazLhWZ26gpQroSxrjFAfJH2Stqqn3xa0kodQdgY
/WFXmxNYYWEb47f/b2Mji/kI89jODmzOoUQHtEaNa+hexooIOVR8ZtHT+hP/4l9Oi+6RJP72h4j1
CeirGCRWN9+VAUa2425/GEHYGWnCQRAG3XP6ucZAKjmySJjigkxBvhZsR8JFpAr+Ykju8dmd6w3d
KaLYF7YcKTU9duO+J62VIaAGtd4HXfPCLVYbiW7BVJv5AGXj7455TLfohoo8ihM78BBW72hpvNXn
1DWAO0UfAcoP8YXLBfpITg9cdYS/3/mRKyF0S6dZEAr3iAYcJhWOZNddQqfAbw+4lZUPp2zqrQ0Y
LpuTMhHe7YCD/hfAok6hgjBIHz5sR57OZ9Dhnbi/7nnE4yPRzPufHsrLw74tyCzbjJ4JhnMpjKfT
oMbl+eTR2ovXJDYnkPHD2jvDz2Tj0/xwFVzwPl1UvChhxt2hah0w/U73JIRJ3afPPh/jR10DQ0XE
BtdyWS8m5Pz/igHnXItitRezX+MBHOTIhiYZQDiY6U0xOQvdxN+53u4tk+aWPiIbkPVfHiprxsnt
EVFKSeKMpTIrBt+T9gFgiVUbFKAhuuEUgnosxLJF9xn56YpL2E6dsfsgiEGWknaAxMOVxh8owjf/
dSIYvZMzk8RgYy0qnh8uBrxf7Iav68AG+6ZHlyJmZCM13qx7pgOE9IK1dgWUQg+qVMeXRepZ9u8G
3xxiMOaNx5QmeV+pR+M8oiWTUwkF5eVmCqBOMifmhxlRSlLi5qtUt/FsNb4ztLO0nv29/13BFUVE
S0WYa09NcU7k8F1uufc1PKBlupE3OUcIRZRdQKMY2t21dDoIgNjL+DfxKbktRcEuX/EbM9w3o+99
qesUJgd7KqlWbDhLpr4A1I33XGjnPl96diiQCNs52E2ZzePU3TgxnKR0TntKv3jcNYMXcrU0aaMp
tiEEtUKapjDdauSmkKdSRpN6zJykyAMvcL7hEJny60jzBiXWfGVk0vhwBgjgYzrsOI4TA7LLOsWD
NPcwl9nSN1qjsMWmz3NkppkFqv4C4NuI3rdvvT2MkvxKSDVwGU0nE5sX+BFreZQELsdyyD2wtRdd
xAzLmpTzMOlJEVPjLymn+OBKd97mSMekzDwOTXKzULmri5qrjepAA/WQBe5E67i/T8NKQZHXwzm1
4+MxcEc1QSjipt5/x2VOrt82pz17ncJ6cL2ZWnqX5y6vonNtmfUbzFZWxkdkOpI/0tdHdoXxXSCb
jnmVRbLkEokOMahmOngY/s2gKh9JsKhqQludidqCjWBZOgIsSO79Xw5XtluqXtR1DEUplrhHzu9K
fTV+fkZrBootv1xCf7CkRfCMcqgEXQNNmS/6AvkaW5R2gl2ZrduENKfmTBInmdaaYTTd6PATM31Y
Y8WnVX9T+qnKgQvnxsoyOhlqB2wasdJw7x8s7xPkO3outZvj7JUpMyazGWZGZpTEo3iBaLRmTmzU
gsYorn7UD5uULASHn18GljAY/IqQuMZg82nVHf3sA/oYBx+P8ZZSpCyzG61wKHIqHbK+TmxaJz11
mJXAphk9LVOeTphpjO9f69reSNUSEERJZ4yenh2ptxtBStGiwB5j4GxNyyOyfALS2VbQ6Bj3gblX
WsoVCACu49nf29ZvmioRfKq1RF38RKlmNfUQFR5nM16ZEU/PReGlEt/LGl4le9hSAVOax2G5Imri
MNDjoKNtoTO4z0gUe4uhTYhk8gZ+B+Gi6dz7Mt82rjN+IxSICLBJKgSIoT5JQTjKpkgh5U3TO3Jv
YHOeGA3YkA6C47vigzttJqCoHF8giWttukDWquaUzjXY4gOsYdNjaTp1OszXxOXKGmG7FeNM2YnX
gJz82DJmRME2hVtMc93K4LOaNxF+eUYfyCZRyKKYGt+q6DXzmKd9k/yzV2x9+kt7Yv27b3Usudh7
zdi9Hbe5OXiU1NgBgdwO+UtYQMLn08jny5sGAoaZX1UOTzUYS2RjenEUtcNnC7AWng5xlVNz/q9J
CRFbUDoQvv623LGd3ngfUYP7eayTDJ790rpIeBPQ6wZSB1tU/qGR0gPJcJpKgKXVowaFRR5LKJtQ
+Xj8NmDPhaprM78pWgG5DUA5+ingBVD4rsQ24502XsylkaAJUORzETLMPV/lhScIxpUnAMt1rcBw
GYzhPTZlkRQaNEGYy1SkG/d0yla+vy7ahTTiq3y+uYPGSJccPkbKd3vVVMuE8Kp4HN0i0Ru4+wbZ
ZptZ4hIjo6pCkEKPYsm0dNfZjQVe9NW1RflSN2J5pI1kI8TG+O4OcdoXKRJdcB5fbGc9vhqIAyw6
p5rqOLA6lLROp4+Ze8PwI64dcu6V4fN6PlQEW7Rhu2mq/PhdrdtEsPeKNZyNzWqGpwuyBFtvxpQj
eMpPVOWkpMMDaP07EbhY5QU3C2RDXs12D9mVhjg8JfSEL+BkFEL7hfamQARH2LrWfqTV/4qDlvNP
QY4petctwXvRjaUkemVwsZlIhdBUACrWGnZsMMnYFXPLbdtaE3CuSVSlfTxjTjb7p1LN7x6KjyDV
YNM46goWV4JKcecQ7+6kUXDeKrW7LWCO4X6cMHHYFZw6vFtvVfjEPa5usJdICtmdWIUcZdckcRMz
5+Uaiv7TSQkEYs3A0jmDx1Sh0R+b3A4dlGWWrwuBKtODVmIVFsTDQqd5175TMKNAFp8bbfyr2DTt
UZB/1cZU/q8AnU+nH0XBqzef+gzIjAfTBWXJ2xGJqrqis1d737+EqNekpBpq7Fa5ZhQ9lcjgj8kP
trHC8uy3cdh2Vc0c9cjmparEeTGcmB6+K2cgawa+zqpBwkAHHzEyKLd6C03pzuCr9mJDEygHXIt0
i+kSRqN6mj+MHBrwrOl4Hn6cBqdHzORQnR5zxwCPjuuuFWkBcfOwIoO90zK4IOptGzRUN1WbxgiZ
Cw9Jx9WtISXr8LSTjMbaVT8eck5jIhDkp2iXplXunNLFpWvWbnnV2IPq3O0yMSEgCSUdmNotEzXh
gRwP0YbFQOV3GJTR1X9DUym3GLuqtl0s8xbLncoo7aHsy9lsOcnrqAtLDdOLm5GlvrvYPJufnGTa
6+PDg4PTa1ZOl7oCCYcHsWKedZogzWkgF+VpTbPzpbKCZAZrQTuz4WiAceWEVRWu6mEn9Xkzg8hl
Kf6O8qFJpzB1qOn36MxE5xFwS/gMuqS8o50hKAvzd0RfaYRVAG2kW+lHZHvAJiDSVMphljhRCjYb
EM20LB5xxYrlRYTQmRWolM7IEeHypANkm8gO3i33HyjrI1WgOacy6WkyoZw1HOYOo+3Oy2hxstFi
5sB/qqMDpUT2R2WDf33a0ZTpmAUapoH89NsR8/J+FtFg5lGaLP/H2/v7sEpQPKxv7BAxJkmG+Vgs
3wcqmEnp3hUZyk/Luyb+btRSOVKau5mBabKhY5uvVe/9NjqlM9WzsIwriiU3eOFiLnEv6u6pVI3B
ad9h4c1uO3CMO7COIBXcvCvaDAboMwy9IxxK6oOFijx96o80TXchohkp6h0ypA/pVIUzZTVWMKcg
1xPp9wXbjFuv4ZKlH605kSMo1x6tXJLST+b6EX1knQduoNCnMyAU5HSTA+EsgI+Dv/XCRgrAtTyF
KYly1tcnym3CwuaCooy7uLMWcg+RQUifdxO0Z+PWkwDVFW1MwVH4pyaPqrPIMxfkRxjp5EU+lG4X
1jUb2JLkDH/5MVdF8/ijqHGCi/wpfKKC3kTwny017PuQpIx/vX2QF7RQW4oILofGD4VVcWF38myj
qvEQEBcayxbl9ijqpS7038CAzv+6uZQAQq3ntmMwytyiIEYeKj4vxOL4eLq5uV8wTnZMc+CyhgSP
140A1UkBMjhQhJmqbEij5BoQVhRyRQCH4K8parlm5fiLPfjb90Zt/h8uBNQeAoVqWgbb7SLP3ACA
5GR13FL8OjeSAaQ4zSslBqDfqn13koSv7qOv+cvml7tiwWOYC6jOiEWXd4zBsoJfQ12He9c2y4+V
SRNoQ3XLgIjYbLXHCPklSN3nUoSivkGgXyHfmbR3UzGfknUyKcNWGT6kF9mL+hp7BQTybaahKMnw
DI73eG4z+lC/TY/uzYo8A5tjc38sdFq8M4vnZkfH6VIpdpR9eX5cD5Wl9A075KYfRb88xcFW9l/9
E+kckXlmOtp9rxot9jmKE76LhyqqRo1hAR6CQ94baN8UObWUa3AyKWclzDlRj7DR43b5fEfoZ904
3pDeuDnD8zs6k+l3T6SHh4ptF9NbjqG33/ArtvSKUx9BdVs34ymKfd5ZUbFz85CjwiFyRdXzYSuU
JXFGbigj12hbKR84/993Ils4ovhq/kjYKc4P2XXFaKA1ahv8pQZy73kLJnzsjM571eVnVj0I4ncz
WWrcIZq0M0ntVhj9ncYnYdQtSx6QrP/6hKonuPpfeG636R8OH/XvfVecqMXITduczvX3HgYA0axE
fRyyxeMnaxnTAqZulVciVmWtPl2i+LoOnnsFjo+4VeIbkU6pPuF9Hqe3xBZW483dHZBTNKU6jxeM
m8EeZuGVULVY/FlmPq8Ohx846WrLKDfm8MoELtBV3cP54c8X2xeXGqJgg2eilk87DpXpMVc5K7eh
CfuJmU37ruhQdWExzFrS9xBs8KV80mtKwgL2Y2rRC0fe4N5GVUJI0ViN2G0f4yEn+hJV9BBoXScT
1jwq2/4hQv55n95vJXgsJHB3PmPRiPnN+QfureC3S3PdT4CHAQ2w3A+QJTzFMUETAv/Eo9OnZSgr
XM/NpAcGG2PqT9Fx6DlfFcH/4F3mY8m5s6gAwRstutcJRRsyfWF861hNvZNN7xEwOnlKVT7keerJ
Ab7PrUsRPMyrcQfhb/0CKlcHL6z8YSw2uMP7IVSYLfQ2+RDM8IAoR9UTR1+lD0xwX8RQndD1aOOf
jpA7GNxCpTknYb6MeQWokAbw0b4jDGsRrpnckiAk/85soIJCoUB7kCLwt2xpifGcQILtNe4+zvgc
2d6LSvh8kNtk0jNqajRRaSY3edVkacO8RsCsWEd+sfG3LJtVQg2z/7ih6kSvmJ5A1QwIAe2W/ftF
kJWkeScq6IC3P5P62Yr/VDCuS4nyi43AcfFmvOcDlOi1QegFfdy1sbRwSqWOuyi6YBtU5RsfrKmD
95WArO2N/GwGqGktGTM4B9BAV1NOi1yTTbiOi3o47fcPXB60eWLJIa6z4bgN+IFarwmRueY7vKZh
bP4X+behHdSglLObf/AN1BBgJj2V6E65YOVh4b2aJ1LXsouYsCBuoBD2Lv14zcXsLfYrBX2X+QPc
UeU7L581CN4jFhuOLVeM14HUBORTBakL2Dj3gicam15RYAqNADvfpGPn6rKDwoeYZNvsdwmGZvBK
ALgP9y8QIGLW/8o9NJj8oO9rHL2VP9fOlIKMxg5rSXsglmOWgPWAO/yqSNXDcS5G+MZrpDbYUEI0
EoeuZtD/RjV2lF7RghN6LJiHJ5B7KueaNekDNy6bZ9miWSiLD+86niHeW84lCZgKhH6zl8G/pMIg
4ZueEq+gge6y8/aTWcxWJ0YYoKc2UC/FIpQeTvXg1OCi1WZ9CxpFWB1tsQHCrbSOITiAa/8JA3zI
FJihHlHlTh/fZSrQtWLRxmUfsaoWVDdEBugUP449e87cw6AShe9y7jhNnZduAit60ayr0Xbujzb+
Ekzka5QHhzk3FHHmGU881/6MobmUF/3p3XboaYDTl6GkFISA1nBo0olRJkwBrM1abcHRce/h49tF
UcNQAD8UiVsSCHVuQvGONqb9qZPjWT6gyG2c1b5TyyAcsXFrVWlU9hVNqHT0DCNYGEMyQBMUhmy5
Wl934A0nRrwz8jRcD7kEjIXpsv5rZjt/5dLzeyXshE5lJusQilih/RSN19L9ODihlSn5bcRwYHPN
VxslhOdLfjeHHF9ui/IPgItk7sSo2U5vVn3m1WeaPOpo3bgQqqaWFrapPYUYJtzzATWLGIeK53zd
i5s9sOxzFISqsLslsR+ehRYyTa/RNtAB48LIsBrQJnJgN/tRTBYIK+hGnK0N/gMhs948eutNkluP
54EasOiZRWJP4JdXYlkwO8l38MN9Y8juUNqNMitEGQ911bwdOAF1Q1DKffpNjgzm47kOFCrgXUMl
Hdt+uYT/D6PhDg6JT59dVwYtfYYxQQ0vEwcTuLDeiwzyzpZjirmAjmBKYdY4nf6jXA6KheSlt7tu
wyv9nDlqMP3nwxZQluLA2se1acu5qPiJTNoTlCpygHUOe0y06HQ3SDLD23zNNaQi9K7DHQugvV8J
shojNoowDPQR5Ff2J6+lWYemxR6ayWLKTVBeVaT5M/FYTX1hUAOT4LoQCIQQBgf1j28l1w1SyULW
h+ImNSCV9BwUQiRVcIp9ihGFzj5S7jlcqXhUtDk2wFyqShXw90DJSI8d7VDrEPI+lj6M/CNfLIq4
O1Y5dcEf0FGC3RHJGVvNCCczx20c9k+o99qFuSgfGQrggYCbnELQ8nFp5XqYAaV5Vkxexiyh2eLr
s4QNYwSKnfWW6bt06wPrbRj3o0UjUQTGTQ2ZXvMnjr76UCQRm2R+8CuFfMA+4zUmIB2VnQqHOAVv
S3ciY/HMCjNRaqMXvoJIKRhntEVit2N9Hw4hB5pIzYY0WgCL7nvwVWV9EZfjr2TmPeKW/cwiB6Wu
SDvN+SihyYXxGKVJ22/iuVI1TGi/fk3En/Zi5Ngu4oTbUviqxJmYhvobcS+eR9M7dYqy0MbIMIGB
bGtZe8K0OEkA4EHBsVVGO3B2l03aJ1V68SHRWWkWoLqc+C+8eWqwDF3xImlhIG8znybX5vLTXP2G
bhQMV6CxEkAVbxmg3iovlWV1LbwupNkIv6nNhmISwoCNG0gZsWVzOfMpa9ZWThxoH0GpEbai8dNB
T7+oj14wgo/JEuv/z8w9auP5PsZEPqraaMnJPM3ALMFJbcoDGhI0IOVbVEXdTlKimoflT7p2Ti6L
H9Uqc1c08qpO255mNOAxOuFY2YWSv7qtadJBVUhc/kghD1LIbXIxoMUFX8MAZzw3yHXCFN4y7QI2
I/CK6uojRgYEb7Z91JQJ3HcnktkvWo1GCQGWD+TvzTD8lpsr96yi3bi7M1Ss2iSwdjHu/QozCIgg
saWKmz99EquGQYQ6rhDnTTQ7SaO3Cf/N3qtlQgum+aj4MgYQdzmN9n1DqrM+iJn68d8eCD+hsknF
+AhV4dfOtwieJfO6Rmjkl+hv0mnMG73QACCCZo6rSwBkdByWXIjKP8ZL1XqtGeNaPuyeBWuVkU0S
0u3NDrIqcqGzx2UO8gns7zGlkX1Irki52UkXZMTP3BJGiBMkIQEIQNtY8DHvt8SjDMOMcowlHwSj
d4PwHz64fyYtuPhiZot4rx5u+KpVMIONQe7zs9czzXX6N8mUl4TG+y8ZbXRTK1UWoU3sRlaqh+Sx
i8aCESQG3i25h+9maWWwU/7OhuxSmf2XPbUhZTFSy6ZrTpQECwHmnqizlPlE3U3DSsRRjMzk7USw
xYn0/YN7EwvhUbEDRlZjBUi3UGsv1kXTeQ5lRnI4dB1umgEMjrLGj/exk0AZTjPjWhvl2M9ffOxY
oTuJktSVq8zQj5dyQuJ5GnV4xwztg+3J1yZeucK5rheLai5ZuGFAzLhdcoq9cXouNwzewNs6wBcM
2Web6UZ51sEBEyINHTdYiFAKcpc+2Lbcz1uVpputwLf4J0Uz6leMX6HUnr1sazW0fPZHTe+SprDE
ddyDEnL/17jtDQVTnlLUE88BEQBAGk+kIUK+F1y7rb6ONMslhb5ni26RZoSJw9e/h1pzwamiDTzl
HsqfiHib0TKQ2p1bkoNTH5ARw5MZ78O9gwT2WF8Z6TSni/asksFfxPWi+5hVPJox9bdySDaJKNIu
Z1P1vb203R6D3JU1N3aRcnQrbHISLV5uWMsXa4eoWFfbCf+fE9q9sVKWvRuRv6oRWxf3Xux5iFu5
A7N5OEfPGPMsF9ejx5jCUIgtpQfmyJx8SWBmTbxONQO7vb98RfUYHrT38I+LrErvzUu7FvdK7tRs
Hqx/70t9U1Dr2Wo9hphli/Ca09JhMSQbntKaYE01o5MPC3PnCZxPaQZJqSx/mw41KJ1z7fL+/EA8
+cBvXzUbm1w7vxBSxi5jXIYOeylUAW0BDidKAsUDsdeQGmzzMRdCByCENdrsC07WZIlmi3mYs8YR
AmEP4XROAEIC/naNwHH4oD9E2PW+XZmtCdhjyEWKcRHaAUf8prRD5MbR9qBeIgNxrjBPSrdOlTQM
w1nZ6KyON/pkIqwxiKw270JBz7njFfve4OQhlu7t6oTS3ssCOaMyCUpaLCt9nLl5d+B13b3YY7r1
YWOWaVnr8VNwdRh95IOco6K3HC3n4DcxWCPOOpqMUuOOAITANrS/iCDQ+gUApfcuFKCcrL03dE+x
T5yRKrgzojsNy4EoLGvzAgH4Q9NvlM9TM54gWvasCWYg33Iw0SjxtRVK11vxQSKeqp1VCG4W6Amb
mUijcErpZJLCHE0b5iXIxfsmqRpWP0Kwy2xG8riP3fcpO7j98p6y3P+97jPaoNqZM3BfnyZlUrbH
vGQ6PL7U0b5QO0oV/mewsPS2GFf/8a+941fpf/q+x6PmEB2faZktBr8zwjoEKTkKmu+YDGuhCQbA
/ajiaU6aIKB9DqgtyZ7q8dtn2CQnGz9XpicpxhbrLy6h/BE7K39QGjU9/PttBmPqpXcIiBn/3Yd/
27gZBEcQDW517zUSYUAWS7f/3R1mIYxxlvn2qTsGc237wQethzs4b2FIbnLY2fpyslgQVIsFo6H6
LHc4iSy3IS+4pu3b7l4WGWCC1wKOY7XA2eJdDvfCFfdkijcQ0AW9HTPfPdQxdYdQqd+0XWTPiMpk
A0wVvyxfVi469tzYWKzukpPZW7HoXeEjjo964Z3pRcRfdDPgXVga4wXcBcomk/1Rb68fkKMCZyZR
ebLABXOjWGZ3DqFPimOVdZlF0DYNKZ/l2WndJnLWwYeAj0CBmVMpPvMWpZJGNUL+SoHP/cEjYsO/
Mmfw4MSQ6FAhY80fEXva9S7J3pcsZMlqOLmhWRD3b7OPmHn8No8aRRr27HaDLqotCiu3Cyzt7Trq
93SUOQzD3AhNppVIQdFIyT8Y3vahtTdTXeFSppZUi1J/PRHBt3Av84hgYhM12jT2d7ggWsGv4c32
lXvBMMy+Am7lCtEi39kBvkDuISJ4L9XasZnc5kl1mAG7DKLtnj0vLU22R8xUi9/oXouCjR8/JD5+
Pw9hJWM6yeAlFhTMXG95IaNJX2EcvLE2hV9UKWYzYNHBTvCgUoe2puc4eO1W/5e73S1Kzr6YQysM
Z7r8XZMaymFt2cDRbibi54k02H7PhRkV8bTfRzyBM62/KBq2Zlnm22/LZo5bIMrJrtbOnI2KhFuk
ITiy9mVBLVzblgkQMrslPxRH80UZICIql9QgNtHjAoK88U37KYx4jFXwcehpX/nqzY9gPP6+emdK
QX1u/w+el1ab0QHgBJldusoIoT9N7v5AmNNxhoHscHs+j/WZB9lRCRzhMZzXcpgYwCPvXHoDqv6R
h9a8qrlhfac03yO+OkG4ufQdyuQ+EtrjeMkAhukq4B4HIlX2XtDXVQgLOcWk/G/pTyVi4hxCa1zA
HNrciDjbCpRR/33Velbnqt4m2SqkbwgOBACSMv8Vwg1xCEaSJQ7KGjKl5EZuwdxb0lKsOfhpMvhS
H31cJNGNvCKLf3U61yiKNM/SOXzNhSpdKI2V3tJYP05LkN0IfI0ktN3nTuV3EgwRkwBiLVJlx9wg
DNmB2y4Ol4aCdjqa1GSBtIwY8b2Ao2uIkQ9n9YLmNTsISgb4ZkWXC2JG61m1ZHV88iv8Ddsf61/L
gJ5JWbbylbWKSmHjyAL1+aAYfDxzc9eipN57f9BiftlSZEGWEdWjqu93ISiEz8ABZ2ihuchl6wPY
SgAaMlZi7aThRDaxbsjU+Y+fC7CuR9Lq8+R9zehp+ChVZMv4psIMrS5oho7YdPmUodXjtPwXqky+
Zldg18BBsn3UGkoGnUCTrrlQDhNbGyaP1GUbZDe67HB/h4YSpATkU4l/J29OhNmFFbxvuABAxhor
aTXqHu+qR5915uqd3PUdFv6D4d8mgwNe5Y6bZBbxB/3SmR/GlRMR7YXVF4lsZxTSg1gW+KyiDkKe
jOBVFhRDkhGhHsh6Q5GSLnSyXzM/AGUHnvXmc1eietZ1SuYEgELMfJ3osQn0o0RJkwlg94l0zJKV
s/tK7+DXcV1CJ8ttdSZXQYpmnmmShqqNl3bnwGAvco1jR19M+npUCHxF3GReFMW2YkmGsLUvCQKO
CUoJ3mOQap82KztSmZ2WrmImY+fk7Dnc6s4ISqYz8jFn9Gqjj0by9UGP9hrIyguIe5BHrEf5YcwH
8xPx5P1ZuWitcfaLQzj8tL8iOey7odF+au5LaiCAQu0o2Tl8koRD4snayhxmoJ4N19XANwMI/6DH
aiINahsukjwI9wEbSAYvdyb0ZbZDeLCoGEqCYGNDgxVvoffnM0IgZlt8ay63kKq+LgLrpinW9AfW
gkSUj3tV40Tyu76xkg0CSJkewKHLRgawc5ZeTIvDoGwgKdJvZQn2q30nOcsSwTGLd1gAvm6oRdkd
gL+WMaCP+MBh3zLiF8UycQyQSm8GdydeOxkOKKe6AeBCAayl3ulkCBbEkBPJ4oxI7Y/PyIA1d7jl
l4JnOaUOqLOmSNTyZ4kQOjmqeIK6otwCsL063njAd0g1KzzpunLpblHkBgeT0g78ECU6L2LeHVlZ
ff3ZQMMqKh+jlkeDymaBxhNTpT+A/7sWPYRDhoVs9xauuzf8LnJpOn+WK4t1fuVt8D9BNd5S8Z5X
tKXezpTTUZFPcpo5DLdWMgY0PrI5vH9HwUklrvv1fVuMwPgK1pDmt+DvZ95ZBitYtXnIefql6VYw
KEU8WPjnAkU3n3kST8dcR+adoCLAv/NoZJrUexbJCMzdU9aC47tgacMGpBAf6qDPt/iCoQ1lto9d
wZML1CTXMF13IaRxwyG5HVwJeLqMjJGkgfaeIqdTx3hFG+xLu7XH4WfvwTWRsEsxDKjLl62I+8QB
lFR5kcw7JW+jrng2ph20pQ7V7RltYhE199Sp5wyonf2lOwdDGQlb1UQp4crJQP8VXWt6n6yLBTD1
oZ4xaZOpkh9gB0pXcf0TXfkTSu86DEXeZS25s4LCHVFa6ySbr9qoIL7qc5c3N31dnJft4Asxpai8
C4BnXHU1fuLRhVvp6Nk5pPPvUzAwjkaHAx1sEgTnYtuh9mA7Umixprv50ILnD712ZqnpAU0kFclZ
X79oWP7RpAXAPyQbJQz9oKN+TFEIvstS+Xs4LTLU0R5cmik9xtTCbgf/ZWomkFznVVFd9U89wSQ+
LYzCt++6Gi8sMqXLdZmqQqvKIH5ZroIyFiATCIIhb62u/an/yl57cxyFmy2Jy7pWftYwYe6Afdj9
DVmrlklvFG1mzpJ3uP4Yyt4PimD3gfxkUPE+HQHRk4bQMEVBYD43ryTEihh+6OHzwGyf3jbv5Q4f
OpY8Tnaoh9mSYpBKGu7809VTeHZzAn2xDeC6NUHeJHfbUS2bds45oCTOo+nxOF6nVO4oIz732Zb1
nwg1DtERhGiky9wcplswo920eYdQnsuQUYyb32rfFF5vzERUXQhUgCTPfhh9ywyX0SY843Hn8mTY
uKjDTb0xOmOBivFYdxxcm2VQLw1P/Brh1GYaIjJqvy+9zWZos58YyxT2hWZejzaKJ6w/BAITuoI3
vjrRPwvMNTAoGRcWtFX+8Srj1vCg8ewtR+5PAnpUb89yup8J1+00Uzz0Y+B3r6TqWJqlFZwc5QBU
+IABLPhAhQm+UiJ3vL6JifTgUNPhTawKOP3xAzMhBQdjqZjtSiYMANRP9IHKS6dRArUwa1O2RV/y
SlhBFQiNLWnzBU90YhaoXe6vaj4Q1ctqD8nHsSgsJjjiupjZH2IlEnKx1i1h+F71w7xjDRA66dAj
R+KZEtjtUJD+pFkbiKlNNxRHEjOGBAED2xx23H4m5j9lkY2ERDDhprTrrbhPDFKvviBuP6PzMlsY
5GLBWsiv4H1c1bPwGMklo0nUECWApD5qDC3JUqvpR1dVr6DqJZBxKiLT+vtSLPSNeug57UU/orcp
MSNQFavt0sMfNpwX36ocirUYn3mKLSTIqCL4AAkAtbp0WakYbQBZeIyLrRoSUzqnzY3WhSUTxCHr
7zRi2OsKfvhlsB75DVTxLFmAB7zUqfl3NU+b0HEcQfJ1WoWM2hhXCqp0Mv1beLW0NXZmyVvZnDTW
RCk7aCSnwrNqioxPouu7vzcQJIFaJsBsnnMV0tZRqrs0M6YMz8g7mb5b4gfXSlnD2nGgyIpnnUQI
F7wgygTSUP4mXl7YRYwjB37JZSImNrNKRSe8qcEEuynx+749wPj+h1pv5YpbAgO7wKcd0s6XobhJ
tvYFgX/01oSGa+hq/pT86/FYM3kHtEXUl5K8ssDrJHomI1UUWuS3yhhQW1yD4Rhk8OtILjeXCLzQ
PxUKtaF9ui0TkAsqwee8w7zP1BGTkae5b/jVRlS/pZ/KgO6lfOxyYLOOMlQqwGmuM8HBY8+41fbQ
F5aOFWhXWbAa4JJVH8OqAHWZOLXaghmI8eHr6WOLwhKgcnaQMvXswemrdnOYx3HJUmzyR+9PFX18
Y1YhDudbUKoFn0Zv3n2e2OJVqNZjGgQWkZ3JvHtbkL0Bbn9xMnyixXvXiOFIY+7RSt5cp3DyI8Nl
az4LnBfT9IR7YHNCz4ubMGk7VYjVVA/WIqbuOimEHfQijIwyYZF3SKwscy+WjmA9hAFGO2trk3Nl
mmB4YI9l/BHkw/o7nQCVbA4t/fEbToIpGn7pkPuI2KXoNsRMOhEuZLcK/eh2Vhj1HmuYd7W9W+UK
JxxRlvqIhsPLdBFbu2gptd4jpmXN4eSQOzbI0dSttdG5/85hkl+yP+20UzD+vP8ZBoF4fw8Gi9ll
McCgNTJEcxIWh/gYzn2Bch6JcSthzLRKbzWJ9vNaBRtuRUPEofkfh4pYsE38sJDE2oFOm0gg10tW
F+7KQBw/y85aRBdOc5EvTYWt0hVPFwiszpWC3wFTWjvDb5OksygbNm/8OLylN892JX7x5HlOO9Ux
8bflBJJMdV/1qu7/5zOQS2IrTDxNQXQhH5N4qjblhWoJ3Ko7qsZXEqeGHt9HXH6la4sfogZHl4kK
lTJXiu5LLl2sirPXg01/h9O/cJQF4FI9W05x77p8Qyih8/eD+p5ttezpSNaGdAQXJ9MFSCVyV3Bs
nxZSU2fOqjebQ+YMKCuixLVIdzNllsDxcRJgmZeZkhEDAt+0lNqSLQ/Qwd2fX8mI7/jLBLBhHS0z
21NBdeN4RM+2TXjl+yPdWoefXaHBzJ+qykIVtiFmFkq+hGW/pviBnCsFwGr8VOxAejv9WOzCBSfc
ob2PRYqTyPTOo+pGABZMyKcjjexWSZWG94bXmb6HQG3WgTMYLVPQwL5J6i4NTO9jlKQfJhMluoZQ
es9N0m4QrJzIXkxpnvm7iPndL2v2agY83lMzfZpWsqc0knBzEEs7+xpEFU0OcPfmtSorLxdeBqPs
Ieb6SMuF8g4giYUR6K2gve4XcGFpcoHFMzD4XADZqFKObkR5PzhnSsd48+QN9X+2ee66xdKA1+ja
XqMmNsJlaCac2MeOPjWjKae39OMNEmq/ihc2cw3NXI60aZ6rktpQVeqPSFHiEDr+DOBihGSQfCfM
iR8c8Ko3ASPQpGNjg6vazbKcvYSUii7StvwQO7pkGLlSF91dTHMEui1tqPhK4kja/DiMVyx5rMRE
fzN+1K0RYp+hxqs28diapwwPdlkfvK0vRCImdEtnvZRBo1ynIlENxrZ0SowjykM4/rJoMxHJG3p6
80OL4yQj3Lp6thtRIMzlnPgOToNOdRmP2kwB6vOvblrVuiJIJm4oUH6A3w3SNfx4oR1D+viZpQ/s
1IvchpvlK5wHSm8gSaet3LKcEkF7nZAaHU2NpMvSfLzWfg1wcBwF+HvKtiG0ja/RQU91C29vJ8Y9
LOctrb8UETwq9jneX3hwuBEuN9Ur+nWecj3CGF7OnIbBjYFswMqTkGoHDkm3J5ASzJQ972ayu0gG
TcQb8DB8r4y6olV1urC2qKds4GBqNANrSMl5MR7X8Y4lbcKT/49AeYxaeJiuioz6S3bkOCm9G4ia
+EcpnWeQRhuzuqjV7vEgUCAC9PtekhTsvG8YnH7fQBNA5C4z0w3HmPW+W3RiXeO4troO8N2goi4Q
vWpMWNzoOk47LTqXoTBJD2nLOlazlkWE3wI56bhP/9u3QrUKF4jXl25riZeehv0Qwxy4Luig8/71
mzsBE0r8fbL9aWey1p9HXQwve95VQAa5WACTHgZJSquFB7eyh+Cy2lItpK5qKNKO1pR+94es3NCx
ZuO7TA0rlfNpt08MxiY/X8vlFBEkkvbkFlitaSkBb2n0XtL8RWYAftvnuT6AdIEwdDOGFDR6UUSR
RYl60ilXZ4C9CEnGFssa6gMV7uQPuKKakiu2LbH2hsKJ5NfUKkQdNV9QHhn1N6PP5Cu6NhsNhxPb
jFSr8c49QFyxOYAPMMUZ1nD3xKLVAnbAC92KienjvBINuYXebYKBsps7xMZRRLPcvMbqxmLdZxw6
wo3ufu9VjRUEjRdWdkAXZdWBKrDzjrg8EtpxBM5wXiWFht8MSusQZhtXjpDYqS4Q+DzJ7KueEPPd
jNXM9bQTkeeUCsBjJsN9OFoEPOzG2I2TORHJdEqBHuEwDzgZ3pQ1kUbKQhRJ/3ejhn6W7nm0F6BE
GcfNWo7TMXNnUlIqCPMXpr5WzuLdI2hQOC8GMUruXmdLT3iReKLZ96hjwbAxGoKIIOAlhMwGgTs5
thpMLyuyxa1XxknVl9MI6gwMTRnBlsTE2edi6fOCFodpiqHiruiq0f58Qt3hIk86YCnbeWoCtBlq
qXdvReSC8K28ywQwrenwpQCQanjT0CnCIM8j0aNTHW5E1QVjHWzgpgPk+Z2ez+4CeFZNAFc2Xhzj
OqP21notsg2A9tvx+x3ySZB6Q0HssWRSlKtdfeLJ55N5YbgyZutlBbL7r589WPc5tjtzIuLUeav8
wSbM+jQNXgtimc2BqC7qL7CN19omCZHe2dHTRe8dCivOOhE6vjgFNM0G6NVKJ0+pGt/Tr4afewt+
o8Up2hGv1SglVyB7kYmOm2+gr8qXaaji6JdbBIs5dD4r1sHth+AFsuJdbHuGkaqLuGWKL55KEsp8
NQ3Dhv4ty8mwgmlO7AMMLOv8Yn0JT7s3chvnIMqCQbrSyZS0KtUGHpDx5QVDpkFZP32kYkGEEt5O
6Y9f4fH/ZFznDsO1wW2mqpQXSvpAiY1aqrJhmYnVeF+XrME+bF5SY+AVW+b+FhUY+acCPRqk/EJb
LBuH7Ppc4j4IoMzLldArfliw8gP97SvuR6D985L9AK7pcAMul2+5qVzTFEmG6SEiiSaw6v+XvX5g
iBCeIY+sH1zsnNJB7NA0pPzwwg4YNthii4oV9RfvB7vQlTPZ/YFOQmw4U4wbqft8L/28qOMSp6KV
n4ZjYGKyofl/mJF/WBx+1fDZDgQdR2FWvDrBBg6ytLwWEtfygC8Yf5ZXh2hSttoZIUmUvNdRbcDi
MQ+LZIzo9zoV28jtFjgPR9vfvux15XQv+8nmXpNCbN8D/n+tAooGKoHtL00tboUNktkJqz2uiuK4
0Aj9+/S+okA5Yd1gwuyGmdl+bjNExwZSHxx+6Ra9nAwN6o4iwdOQEefdXglLjPPVsOpAmP+bXLwa
S9qn2fWng/YQEWrQ/05eJQXpTxypdHAqC4BfnSXykgrMGSVUi317NPpbdQkpointais96QRQZwjM
Jpi6ND7mRWslnu6sENCdX+9k/cF8DFeBtbA6cTsgldCp4eASt0nBmuSMDbkbBnlNyf9M7eX/PA6b
Ejg5VbkHkBFj64Qri23XcgKyElFBmHUHXfdDkw8gelv3N8VZH1/AoAo2bCxHLWzCrsTk0AE1/+98
3Ev3sLbJ935LdsjD19PE+hlUHPf+/B5gCIfqJlaowDyGxuc7pSPQ17ZiosyrrNCOj6pfdL3XBimQ
NK+Lm3SFRTgnNMTDl1vRV9/olec6yZ/mgKm3ns3FOY3rVJx09imZUr4c+kSwo2ZuI3kWa7GlDWgt
+t0CRvw9/8/UoS33i/eX3w8+8ra6ZdJAFuAhx2dCGVYEI6ZlG/kl7tlmhJbA7O6c5DwIkV4kttFq
0AmWDCTbo7YNt5qxMzH8Sx58tkv2hc+vzw0bVIHnbKZ5AQNiu1W4ZHZTVNt6Gnnn+WT6jGpXcJwT
wVL41/gSRN84wsyFzg2/dR+G4bENkx3FIV1wPNxCM4rwoFLuKi5U3HQ28MMn3Fc1I/XQvq1XxphU
eIMHb6HKZGbhax3vT8O1eTu0Act2dynEWDFnF+vM5wK/aLWXsh0BGxr/13pdt5QNRjE0MzxQude7
e0CtMlw9DoRRRIOA2aqBN/St1Zb58+e/aDbP9pzvk7dvnIBajZPYvMWTsdvQAJg9VaUsyMI0FcOJ
r8rLoMcxFhNb76KD/DdZnl/WFiO5K4qmGdJmFLuimp/m945VkpeOXb/WQcXsTEaZm/S9wU9yV2+O
g4QCX2QA49vVmB4wDm1pBtf/4dEwluMifgWe7RHfhJa7J0fbEJmuUcQ6ZK3ZjDG2eiffr6YveXVB
crik6ZzAshlAxrVDWtA5bDBdNEkpJN94vmadO5HJSSynjKJ//qCFBLWgT1d1LudK00LOfgS+vOgr
1brBpv7OfW3LEebJJDqyC4Qq8/0S2tbGMKsdRb1mlyqQ0yGT/wlqBVJB+RpMmhDl89NtMmHrBaRy
xU3CVS5Xqr3C3r9PSglLFvNSNM89l4IlF1yapuk0/PUQiIXfAkm3LlIYgh13HI4/uPVpgysXGlxZ
KGn6BYaUlGDPaF/XEqkl5S/EoEl9vyPCAG45iSOibH+xogg9GtPm+FG7lXdkLcfoneOGLPuQC7iX
X1x++jaxalgeByJQN+ZSuRqTb2sMhkAQiMcLOopx6SaNwIfF0uUub43CkeT9ACSkLQQKk8fhog/A
rx2OeivhpvWWUqUnV//BeSCXZPsVUagnGIGYKAEsSHyuSuvn5iFiQG00ahc1pBCF0jJbds5bAPfV
ANnuVCHtChU/j3hVF3DODhQAbOAfl+46J1rE7lGJRlwBeBJCqhV3y0GeL0BJob+xJ3Te5eyeZ1zj
mwbU+aoRqNXfYWGh1yA6e367LhR+xAxPauLoJbFLrIROyQFMxlFeDdNNhNhqgyP1POVA2bcu6OGy
fblfHVXW/m3ERWJki/zM0+yaGaw2C1ArTHgWAQnWTRIkJGhjAYWR98+4+1yd9D4Jpz3HQ1Ic1bKV
XLSGuHLcZxKWHl/nst/VtjuuSDUyN5cD7hpytVOaYvjkGXL1vAt1mj8c90IPMzzUmzr+WpUw3Edx
0UIA6+ezExL63jssO++YGFlwFe5KZX5F0L3MFsWKT5uObcr+sdpjUt8J4awRValBHnuxN0HCJ8Oa
LC7ofY9fr291Wo0CNRkJ2tH3mwikAzU/hqX5NegqBZ3q8gJBFKkTVFwATPGtoRhGE6gXmErL8Ubz
2OzQSZxozgOEXXt3RWHoici2oJv2YThuiJq7rmNgpzkmqikAemsi3iYjklvxVRqQXHDyX0XXqdJR
RKN3oVB/2jlZ5x4F1AJjMitoP9Cj4oXoUlMWWFkVSqz3XLjyEh0bY9kZAS8ynbu3YZ/ykg0iISYS
FJ9cUtSWp3Jg+QjGqmoIq0hNx2QSJIfiEJKhUBrLkBKkN1NowWNDKwKQtwAdL/1yxAsQssZ9ek6e
3tE8bErJ0Dp11sl0taizPekcIqQYWlG+W64Jld8/iGQd/QrBd0ChntSBJazNxhofCfwSRWhvjfC9
kQ2iqu/MtNRYN3e5wafYv6D4VsnOp3oGCA/9Zu2Fxr2VPRs0DZd72kyu18qi4n+1MWewEP0kVCkr
1k2aXh5qJzKdVdG/sooJawuwoBQ6aPUXV5eea2CrVPHpZNUJ/FpS1MWXqk4xVyTmaUAM1gv40T5n
vGFidwJYfF//j+ASHKj4VxVvs55xBbMe4F8VSLBy1G1ig57BC4+OxXJA+Qux/D/cfTzvWuz0eQ0k
WHbHvqeiQC5a2FEnIja43iFC03vXyVEqnkCbdByDukkcseLf/+r9cmlodBvV+PMB/mvAnE1YHaT0
4GzwYwEidj/1ubO4u3+mFK8WvX+gjrK8J+VXyeRe5Oiij1WZG3VfD53UKOjnUIvcpN21Vx0tiDpQ
WLIxLugfxFK1X4Jq4vaXLcrKZ+KyVlaW79Q+G1hwwGFpdqbbZQtCeWKk614Xy0FmoVUjypawMCg/
UKXuD4BKxr+t8uSXdkrNzWw1kXLUxGRrCahRbLd2CIpAnd/DSUi2FEeYsjL437k0Xg9AB+OCiqpa
RII7sqt3scM9mgNDFNQs4Z7DN/dNIAErSmAt/Wd94Va8trUj8aTa2HcvCNXLI3kyZIDy/xof+Lto
n0VDxeL7KTUL4Y2GpsEiCRCfn5LBahOQ3WjaIXFB7eL+Lic9TIJmzaRiLgAO8VCERindlLL4rI1j
eOiSK3hr3UmAwMGLJ01/Y6TKb8Dk+HuKxQpNoFvF6aS8KFm/7aDySTJwhCz0UUKj7eP4NEt0alOf
QxQlhp24ycwRvd6pvsb6NKJ13J4FJYNRhU9yvfgKJj/vTMmqH0/U9MOujAEYcY/ZYW9o7Cd6jElY
V56km6ClwtmgLn5M43L3//Rx4s3ke4AV7who33AUV1WJ8Zb/AAOHHFkn7hUh+m4aUodbM1YRE9rF
rPepZy9DC5O1WJPjfnSOzO5cDB6tp6QbFEnIxQmfNuUBCaw1S5xgOeF9iLTOg3Zv0PxTmr+ZnW5B
3SJC1fNbCyGsrbRNSDjhzqomrwNBf0tOW/dUuHLzW12SlSTjaJjsFe2u7+DVRpe5z8Uz/1XF2c1l
lFpmqRrlScGm7cx/ejS9M8gPQo49+YSW7psgbr5KS4A1ZfTcMi+QyTPXGh22pp+iVaW6ZbrOT42Q
mAlF2J5Tpg/XiFyJmX10fug87/gwpRbp7+4/2s0ZQsSTyQ19b044b3MU77q3Le7MYL3gKuFiew8l
Wln3RgSjSC8+b+T5+Mp3R4iFXqAos9iJMxC4bmauVmy62A8Ug5ZoVYbGztwKaHQEMyCxPNgLLRBA
ceZTaZ7fos1R7IOaCFzIl7vkUjP9ankGEhpnAkkQeMGfiSyVQYQRSA+TkTTvTrly95eSR7H8jKnH
qS18Sf0EgKcrFODLNiWPF4sfQdHiBT3H+GsSeZo8pfQyXZwIkDAGQ3ZfkChLF10v8ZHEq65H4VQv
N47rwBDP5lNW8l+WgMFw6CBYQ/5Kxw8LQaq6izDF81KWCAveTpm/LUji3KZhCrCx12rROTrlx8q3
hCOIK3bYvOF8/0XEdNOo8B+iegS0ihAdcRBG1Ts5qoanG4SEgrKTnrY6pOLtqFa/YDpWgtGLFHX9
47UoIvIYiBBjFQ4j8eehfhX8ZxFJmlM3m56uObCPuFSCQMDyYfbHbPjcimVspMl+CuyMVnZ1YH4t
fW2Qy+w/3sewDOQwpxSq8ropblNxp48xwKa4HvfPXtufS/i4lxxFo6ZhQr49O8gAsGL4dyihSP5a
Uqk++qRC+b8ZPMpvbMOX/lHDEzSSuHgpRy9uze21BBTl6DTJLSV37gIl0x0TmeNHaHvilkzlgZLk
iWnCvElQ4rPlQDNTC59m+31+fviTDLl/zSwcEFCPU57/JgpL4UrMCwQJEmuuIhxKTGPYorOaJE/x
B4bPC0nFBO5YsFsjuiBaQe/0mVndXrg8bD7N7gD+4Hp2Qu06s2A2zvn+W2Pp0Ul9sOEA5D4gV1KH
nH6RtlyLICqQnm2bKlNT4vIDbR/9CZL/Y3E1vevnh5So981tu4kIo6sILwFxGKmUCynQ8ZtMfHqv
7x8h0JbPbxe1PZfYA0lpUhBba1mWlm3kO1wgK7uR5QuMYHgpSgz3NmpwCkK1B80FmF/R6aYhUARp
OADP4V216IyzbhlM293XQG0ZbYhbdg1lkrJop6BuVCp8MsbsdFUqLDDYdUVnf/9P6mK/xQbN54mX
naIzN4uq0y8risO/CEMV2hNRq74rxTvcYJvF2H9b1/UIghQeBUNl5xtn2xzQN2p0Emai9ROJRnnG
15jfivdPlWtIyy2WW/enlww00V+iomtJK4xBuJAD/S8O0toFmM5W84WHLhpvxTRfpeZFjbcSLccM
SHBgoNG3akOFWW79FRHfB8ph8cw44nXTDIqkJatExMSrTPj6fBhhE6X6l4SgNPbXeaKoz/57Yy84
dfV15fN8osW17BUt3G6er+8R0G6hJ5G+i3Tx/qFBtMTRNuvu3V1xLjjg96D0gYFXB8efZMiLuxIe
UiIYj56tGzsPh6btKhyfnlUtKfPXMD5ZvEJf0oRHc5LieDpAm9npfn47tiwaS7Z0tFi//ygGlEtR
PbpXfQaUsr4FWEV/i3hd0NfuUi99umIgkXhJjuNRJAKgtENDs69LK7cc98LNEwOEO3sFyqKAvIV7
NoxUUEp4XTzE7CvH9hBzAEHxQvreVWI6YWzMXBMJPzLY0gjD5481ZOJFqBeRfihCsfqt96sco1te
XZ9H1ZbXfdZ+HptRCVHGbED3K2cGaiBQR2eg9xwIfoqxhPRS/FL+3JI8PJfOCWciQEIWcv+djyS5
aQJsVYxc0gXPf7t/FJK+Km4dJ3pNQeANp9saG8/jDk5DLsKa/TaICMOOUDL5s/WwF7wWATITELr4
+2Fdkful2vYtexx37ZWYp4DfxP+A9pwtpofREZYHWWFgNYpLwGysIfZ0mgIyg4te804jkjs9vaOH
5yVtGTXVRpqrbot4MeEaIms+YL/WA597D6UCwVkY12ltEW71cm98K6BNg+ndoWWVdT2ezeyKiJFn
jefQFTuaRYLv+BXnFYCNzrX5BNXZzXoFALhRR4y/tX18pXL7JcwUzBm9yQzm0zD3N0Ww9x3gQfhR
jbg+PMgvIxh2L7mN3BjKyvQ38tUmWlV/A1U4naGMnf7XYdptM13i7dkw4yHRjXZeVbdH9cB6W5rP
IKHdi6qMQAhljZvrGqyFKnwk3zTZWe/OBx9b12VpgeY+12A7LVrFFf5RFKiUgPzZ9KyM7PFib4+K
eZYP5wqX0kYP5W3b8CyXMO0Qm9AMRa3JnjLRSQeryKRWZKKEpqHqUPGM5dt4g5KM1KsOPqKiGeEM
JiIzdYtclojsskhKU/kpihFTpPE6QoKvinyAr/uapK7ncKFhkAkvtSj4kbzeMjy4Dc29vuiOgCIp
e/T3gpzSJHpf3bdQZMdVK9RTVlYAt01YVdy9KDf/ZvUwr4if5jWdO90guvZqbRPc3yKs/VgpoNSr
ZIe4tLwrUM3k9fukT2ubDIQcer2cL7oWPnWGQOf00Z1olgo6PnuKJcsPmHULh1IQy1GhAsb/3gBa
7oTdhLNUnbP3Sz5J9LX95Q1jc+o+cEjTVU/d4+G7+OmScOSq47Vq9lw0vROT4i7rjJmbNXSvtqTj
6iPLecrTa3jlZytlPRrMRTLpGyN+oJevrborbKZkO8Pwz7eyX40800ePE0gZWVLO9ZZaAqPMRKwu
SE50HRQEYt/7Rhk1U8uvgL5fTWOTdCkR8AIcgMCrAwVNO5ucEsyWCL576By04w+xqvK00dU7+vBw
AhoOfvFkNix65/P0gvf+jyjRZPv+MVkzr9OyatFdGXSRAvOEoux/UCJE0oljcwh/lbOmxI7Az4Ps
A7X9MEwpmnskHm7liHtiYJOBLFLwrOoBSYu5r+WQLSC8nhirSdrN6huTPRC5yvvz9J6/z51Eu+W3
ShC2B4l+uJM6jTnvyhT9CBfUUsube9f9fyK6OdQxxkTX+2TY3qeTIRIPBQlAAhUtIINBDQUbuwCj
KX+OGwesxIaDK8I962hsDnEJWki8Y9DizhhATTdXSwcIF/TRbSYP/Mto8JBIBAcnJ90hGqPywCxA
hQ+Pm3pxeLch1bscJrbKVjcSHu/ZZcwDUWlzzroY4RiHkgNZYMPvGoE8mCAFF+nHG6Cf8LaIoX4e
YT9MCZFfXUa092asML59C1P+skETaL2pYFyxSUBqnps+UpYzYC90Zc4QI2c3eKpNKOT5hspGUlqd
KovcjHf9s+LYGxbfDSSwhi1KGBUz6UIABH9ADE1+AtVQksiJF12D2KuKan7r4+mOizOgd3G+y/dF
m+ELmmVxuqU9dLiIQ8z1Z/NgLMmH/ee2DgvYElk4IUMbiiAgaK76uWhTl81J9bHu5a4tFpNH6qi5
F2hqNXnoSWrCSBcUav5erqLauGADIyfTx0rsdY1jtRiBjwwsGLTuL+6b8VHqlgpT4aRhl1kpGNVV
ZD/YFlU70a22Zp6hPxUKv4EZEgAPg1FfK1dcQe2xhzPe7bk9b7ud/kkaa3VmqPqC+MaaQ257nkbd
ukAuRfUzQx5yG1IYX7E7N5BbfYIFMBmM+uBhcpeXTkHOd2j14iOcTVX5yNm4xlbhhpVNhr0hA30o
VpIFItAs5gZa5yxTQfKTjR5etdmbaPy5i3b5tsOVFVQ+IQRmOctZ12dsL+TzBTi9QzbTWgQIXTvI
K427jNcMqh2+pWg9eNsPubEV2TZUiRuxNwWV8F1zA1dU9HYwrouYBi2dfuUPyMYYF2aIYF91hxAs
9FIG2CDURvlpDQeX7wjWWBpdEXycAec7uBONKRkws6jDdsBUtMpsT63fWJ6R6QvB3GOCtUgQOshW
Xn9jOQQYpKPCWzP/7Rim7HHDEV6iqXbiR+dgCLSFyYiRrolTa5ka+p6YpCARuWE+SW8x2rfsqC3K
7jYMTSGIhF7un/Knkij2ZfVOG4DLOa1ECEPxQI2TwDllz+0fVOCsT1qTs1ipqJVR1BtADOmJpSHc
QkcWgBY7i/BroL/2FBZDAH1JjLolj5T8Ima9JA6iOt7Sgzs4W6OjpX8Rg43jva2QMNtZebRumVQU
WjBRgNTh8tL2ldsFX/ONrEfpk5j07uTBmhyfGuxIMphotioqvyTG9C73TfMngzM6FrTmOFxZt7Bh
J2gTPG6gnW+ldgVmZqAJrwk1zbdxjJKUjA/L/mUsMe/ROAAQzaC0BqYc0dLM5ABrypCavegj3cXS
NPae75aehUDRO2wnNHD22Ll9tl6s01kT8Y3ZOYJX0BhdrmniOU9EMOd25cPftkqvPdYWjexKsji+
i7tVMtSNM/Dx0L3DucO8il99WbiSFW+wyVIdKR9Hhpgpb1HQAEYiG5JZAG0lxwRzBzwLSmmd9nK3
z3/ZBBWW2IW4oAcJrFjkvZdv7XVjXH/FCmtq3gVzCEdexBssF7Bv8qBF4qI2xxP+KH21A0mdOu6A
+KMAm6MemWvmuFYAI2NMHHreeMCzXXrvLnh7H/yV29aEcokI/DdXouBVPFotCTEnutuAfMCxIZsm
hrlU7bXL9Q5qBZh+e9Vx8cBRbKd49dBM5LK2fzNfVNZw77DECL0OEZvNlwpvgIWi41ZocCazeCSP
C3CZc/ddSEQ8q6n0lDXX3uJP5leeOnchMzUpH/To5cVa3zWiDVRTQFkbRJ3wpu+zWBcpvsTUahSh
M+6AxXXfqCMt13susE+4i96dWIwibJqp+hTFn//GvktcM3RPRj9VIuA0KV9X8upftY+808ZqmqN7
wFTVQKtnS98IUqlydZOOhppY0HglQhIfZFvKRKZ/LsRcj4O92DT7ZiWDK9NFB9695PaM0lzTOvNO
U8CkvQNR6FKFxKcZNRBH8QmRESPhk2k4/u14CPbxMy1h3Tb/7HUk0DyAPeFUkpQudXPcwqHHpwvw
2AYj1BQVCISId5CxVfNliGJJldgjX102UTp4fzQst3oNZi6Jb1dafamB9NwJ5gewUQVLeA2qaiQG
vdjVqBNeHwcIY3nQjuffFFvqXCdIZ//3RLnJ1EsAek6ZDdVtWy2ZMtdYZk07NlHQUF2iOuDxNqcQ
aWvn5FPEMivKvPW6IrpGVmp9HCkToHHE1d/vpkZ0nWOTQAEX/8QMYkGAQkwkcFBsQLSPkOSWj/0w
Bdvbox2yNBnRU9TDTvEQD8OJLPOuXncmLE5MHyXPCq/YdChOASfI8QfsE39s7ulC9dsiIPclOQR8
q66q/8csQz8oDxE3GyP68Eo00qaX+lpsk6JdxFh2BwChhQmNqThGnOcYnT6Jf5n7iO62Y2IFD89H
OEGr35N+grsDOnYspNRsOX0A1HlqKRrmH+Otw4sJ+NsK3MxCutCkonRO+59k9MszE82UvemGYJSV
A6S7+Ei7MwFIuVHDhGNvxviIQJwQDTv0CEUffoDmmdtkG9lY8JTk4yF4PS21mXo03uFukEYz4II8
qnJi2giVQokiO9uE+KxXADPo6XSDbfkoZEWJdKgVmC7rquEJMNR/qSo2jA1IHB26WImp1CpUR9FJ
VleqfjFD/FtnTEYrYVJWmmTow8qO+YxWET4adgsjQ1k/CLrrnzaT70+hIywTOP1knW6MSiD7Ei/E
aDzZh+JsEq5SpNUaJtbSqx+PbkiHoK9jgaqoxfTOelI7vFOGfcREvy5ERpwY4swJN2gfg3GL5by2
ZUOmLL60e8W63x7JvXJeB/xRCOTVPw2dPLZRvOg7rsRcxbBrkOe9U5SEHk/1s9xgjPcwsEfEMdGX
PvRbc377qoK5JRn/aNaqzu5Ksj6Dd/MuEGisFH/AzvXQWISIB1d4RXizjLngBnAgrSSwVrdC1c1s
VTXUU2ira4V5YicqNvYRVdyjV4dqjjsgAJbk530otU+qxKGrX5cJ7r0hF15VAti71IyVIYHeCUm0
uHx3Ut3OyOIqtsd2/SFz92/qIRwEPk+MZmbm55lsfegXs1orHCeeNPvK+oCL9tR3MlK4fGDQ/w2x
+VF1Q/CNfQ3ZnUT7GsR730frJ4HG5+8hUH1iygWUNXT2WdqVaV0zbjNRuqq6awpAKAwuk9zaumBe
9y8KbCCH2IKa/rfgNWoy83ka6w1Xb/QLOBTiK+YH8u26B0ydiWGPOcTTXE3Yi9V5Vf2QIEd5ELSm
vklJ+Iq1743pYPOxYpFd/MsdnygZREj4QF4w3p+UX1pAFPklZHmxKwdZZOwHiMXM2bvovcIdEMs0
vk+wu/Yk1paSPIMaBvid8+0gOW5qw7c+COmI3r4VIn7g8IypEgt5qJnRk1xpVmUP10yWDb3jKyfA
sPa+9Al8A38GqIny3IFPm/woK8iI2MsDfBAFzZy/S48qs9q1XwvEPNFLei3Zb63uuTYz9yurHBMf
YA86u7POgOQmw1T941CQoQ9e2BRqi4zCP8HoRUiXRSO1IBTXWNYLokcXU8Gsk+3o54opHe58dNus
fUo96DpLgrO1rRxLlFOs1A0KcPchiV4Rq5X0L8oEUevuZREWnIH1+TdYjpByZ5mZFzF2+TG4lSnH
HbYYX8C3yItln2vsvy5crVCGMjqs1uLlv8vEa1mgUaMm43wJq84Ous+PLdu8s1fVubiaqYKpAeUF
u13EtDyyOyRuEq8XDzxQ4PKBBGZM9ovnxHU228H4Ydqg/YVsnmwHnNkWwPey+m52zla0ygMtdRlH
aX1a8PPQQHy5nua75HAXzkzKpOTKr2hSeMVHLzLb3q3b7ywyAZjP4vmk0ZWzfxeiCsjTnNyXQ/A3
SxStvlQwtn95+eLSgOnIzgV9xbdSAZQ+CvS5LrifZkTFarHzmQ0OZHccLcgVvFA0Q4qamEb6vsXI
4zdMDIDLmTCS7Cn7wvJpQXFvwGI+RtTwVpqUZQihe/QqWCgT5Tu7tvEkdXAJbcbEuB7YaGbZAhpp
8Xx9UyfFNVMu5pMxoJLex8dczMLSb0n8VRwrj+u8yH4mmQJkjQAxG9Me3WcZQJvqupzaTzvsGZlT
b78105jyjsUnBkkSxfaNFUQ5jfy3oE4YY7gmifNrypiCYwpZCGrcEndO7dR2Z89TGsktZ70svQnZ
kWxX7YEowjPo6itE26g7abcBDrnynV/gEJ/v013KIeaknawfK/qahvJZEeuQFJoBlIae0Enltxm3
hbkfhOQ2hVnxFiNhk5smod4wz/9L7/TwkuGOwPMxI1criQGZQenjHf4RgjpfD7yRC/pPrTIHF4XX
6kzobrCLQH9QH34w90bB8O/YIVkaLq91u7ayqeqvOd2JlK8JmmqPHDU/CEBX5HDeRazu2AowBiM0
Y+TY5Wp14/PbUF7pDY3WrXctLOuyC7PV+Pw5nowSgjYgC8WPBsFBGp4wv1+a2S/DPSp/+icwnwNJ
ZguOEYBIeRZJEFjQkmHZl9uhzHT9ApNthi7JRwEROM5x3iLbH5No3PZmIafcP1SvMzCL5Po1yU50
OonhvwVzZpYya4iOTkPVFxv5RqDOs0U07IhCjIbHlEYv/EFIWeHZtvdBL6rpKHQKvTgVNerWPGax
HOA1BxkhxPoeDypQ+uP7c4M3Wnk0cJ+evkA5Oh538csiaX9qVORIZP2tXhW0T05mZBMIRIXC+3sT
kq61F/S9Zx3vBIRzxZkmOl6efdPG5CG8+8QD0LlyEbYdi+ImgyEkaqdeyFSrqFLDViFxN2Y8TNst
Pbz6W5flwaaLrh90X/FYuyqlfK2U6if3E7LzP6sPLAvkYdtCNwRECXXWugjd2lG/PGHOy447ruYU
dKWYzfl5le2UOk5hZUpNyvUkkKgp3e+vY2k14GHHb5M/BhHT7RLvBg3qPp1cGiHSRsASdUZeg9UR
AjxIYTPdT9P+Q75/yzhz6AT6rHiv7s05DmNcIFg2HCBCA42NoDEA0Y3tl/zQLgVsqGKkxC6aqZ8k
oBA4l5rsgGFlnclU16ITd47TibGbwJdO1wz4HKE83j4XWzodTTJsSfOZT2Q+6TCM1sissrhOGZWj
fe1WCC02PQUyb3xJiaHGQdRRvPY8bu5WL/Zho2WlMdapB13RIlgJx76yGe6NqRHOKuugL4P6cd1L
P9K0xNzIDBS/U28h+5LOt/qKxZP/Q6eGfvziJwYdDyiB8LM2U9PmKSOnOjW9PVbyIKT87fdkOgU5
devmbwJGCDkKimzJELqGhYZ8C+thf7MYBVaWQW74IJRmQBp2eBbCbRDgpA9UaHk5KaMiSC9yiRJy
HxTTypgNU14D7nKHtNLxvB+w1Fc6vfX1TTIq/rN/3GHRKDhHg/n31LQufAohTl8KQ8M6WE+QgxUw
VSw1JosT1jMng8NXbecZQmWoeyyydOvj3qBfpNKhh1w/9x4oi7uPX7OW3tXg0AKRZ2weSkk762cc
H7gRX0LVafb7kR+laHZdUhvFLuen4rFmH49JOWz86z1o0UfJwgeLn3n0TILC2+tNJPeV/PY+OR5m
4JT73Oj4SPH6ZWdRIk0Bp87fTWGexikOIEdympJbyEvF+K/Ij7HjRYN1REKc2M50Po/WDV28u3RF
B04xxFtHLtqohI2Cc0nBZnrU6QJ9xby2Dk1jegkhhQPjzXFG17c/12N8pTTWCDSospO0H4NDzJo7
+Cb0Fb8H8HWIiaqn3CaosTKIGdKrKDYt6rBYQQWbpxDuivA7G6pjQYXuvp/R7ZNpLXeP+YUvM+Ih
+9RZPP1EkgOSPugFZGGLOiXuatqY5rYw0nhlCAQTMHDM4uoOKG3qIaKlZk0JqJox5xJ5emc4oXqS
L19hXuobRK0csYWV8PS3+Q+J4nbAmWDgHemafAZYQDbYjauGIBYYLcf2Y25mSZr6p0t2yvNnW8us
HYJ/vNQZj5f2arTkGR/rRbF/pixZdVdVf3s14HCE+CR+GVPgr/hCceLZ7AG1D4xGAS71hjf4kWJK
Tt02yH7sUeAfNLDeeQJE+KK56dT3InP/uHuPLBV+3gc5/OFyb1GKteCIOcJ8tAjvQPE97SLqaOCF
dzNDIpswGJVopJOXFT9D3YiNt3KlFS1Xz7nLQWvvrV8AvxfTB97dJzzgW9jOO3xtEO5uI7sgjKOf
kHC2Jrv0J2Gd8HdHJcTGaOhuOs3z75j9SOtzdJhJK60QtOggcdaLgByYZRFCdBI4YPBUppXaNOJi
Em/V+WZ1DiHQFfAPLNJa3rbS3/EUyeKG5h7Xw+PEcQkxyEv0U5Eq+2nZJRJKBlB0AyN4j7u+aLYK
T3xTe2sxax/R8vHWKVbBDXcjcc25Qsz1xa1B4+gTQhyo1Y52gnLw4aO2ctxxW3VEyYohG+uT6MHP
kQXVugzOPW0wmd8zlsNrmZGa/stiU535Xo0I9Hx7FJUvEggDVKgYiA8GrC0TOM8Vk4a/Blp7Nljv
6Tg/oxrMLlqXtGb8d7Bf0gVB4reg1w113qP6toyyl+X5yv5mkfQxCFK6xvLoo2DBnJm9nirfuiGL
grxNzN3pbKBhHbh9kiegkwKExTzZwPVk6tx43/yLX31GIlJ0jEMGmcWCCCsBiCD+XUVoXoW/HKk0
6wHldd+i6m5rZHS1q4CIA0ya2oXRLUBO9GEejlHwXkiGWFMPcFAka7XcuQcW6IcAwcbF3FV7lbBl
YuVLqpTn87XlyRKX2PNqD6OR3a1attBSPjHLW3J0ykR/gxHk57vkAkDjgfgXtMnarz+X8bKRwZyN
9YqAZlGkrZMFoVYSv21NFWrD2rp0Vw3kZ0lHC1xmEA2BR0tky9rurdjGyyUYdJHRUZPrH18wq9F+
Gg5vjmF0NfG/rdlhX4VwTkLarec3FAGKBH2pxdBd/revx4sm1Q9oLleicudbcNWFROtVq0bVPE5X
OLoWI6Nho2jlktCdiLLDrS6HHw4NR2GQkpF1gcVUs1uoV1+hwaGaObZmGpld5iX0GHL9x0DU+ABu
T20RuohJ3m1674FImjsiiRdj7C16GbRTlNp1LUW1rGp/4cp4uvoOL6JQn0A6oYNNVntHEbk6ZWF7
/YI7JmpN9w3L1CHhsT5DC5fOy7axrMibdoX8ndP93x4jUBS5BcaFZJRgRmBaJKJiS7VssIsLYxms
S6FePDEFUgsO041y+rhL+1TDqrdN65O+Jgjp8FDiWBzJNvuCXwyrQlaZQRQkKscXVOWTFPDqaqek
zrbkXbUjvRkSR5KZDC2Ps8S076UAdaIYVQxmiKPQKKFrj76sG6ubFMxxQsXGTLWIEau25O7A5OYs
TSMk+LKn5P3tHA35mMNDUHymcyxQbJo4k0gDO/jE0CTlZ6Z8/8n907fEvzMiW7AUP1ndnqcdWy+H
DbyPn5Ufg/ycDITLfAdgcssfX0hdx0PoGKvYqqhR42zN5yi69YcSG5Xvfzr4FjMf66jJQDppMeQS
7EBhqYlwvYfHKBEn9JIi+Z68gpAVf4oQR+DFiEfSQQF/hMjy2+Gb1t3gixoqqUeDKy2eSid/xnD8
ej7z5k/sYHQ+TXN769x0odS9BzOJFHOGT8+dqJ03mWb2/1Yl++RbYN49++6kRPf01GBd+onsm2Ru
K09OTeLFBbWdnn3LiKCHEa9q2BImUvw8dPlrO1ncvIRsxdGgcvSExeUpcT36ACi9LeSKB/cvSNqN
mMUpHzY2A5rYql0QiW43tXA60GJ6KbpT+woiG6skkJYrAz9WmMOCPG0HhezYZbOCYY393KHUQKUp
o0TH5puF2LmGIhD9sfBDrarMxktbiegbp+M4qGt+hzi6NlosHMoxNL5yWvBYvqEycMDlTWXZ7fOK
B3wG8ZFA8T818R/fbqmeGZ3DSc81VKdfekuTvubuniljiXgwABJAIMQX9Eore5RkI6P9Hv7+DT9T
SEtT2/yXAsRWiSBbAU63MCXtK83Ncsy4MkPNJddAAKLwteUgZtfWFkeehSDPI77n8nJtxY6LsHuA
2Df2/nfpbrQ41a8rnpjXj9mY2RYKVwOErqLsEs6irF4OEEnPmAMHpTk7Gei5QZnnP20SP4S9k+j6
KPO75z7D2zM93wZWXLqdcExlcr/QrhDXke0avokrSRmDtA6aQSn7qWcMfqofA3TKkCUQyQCymtSi
/gYTczjf0KyfLUyJaTHRHP/1+KUXlrDUvSG1zt7UyX1hUmEcrrTmggQnFS4CJX6mnWVDIfKu0c+W
TjVzTcB7LGXif2yjP6d9Rh6RjZBf+sDzKbyyMzMCh2rHQy28Er5EVNm1/+vujuOdunaAmLZOZ2zq
VFZqA70GOlfxX9cuAY+olDotAdfno7a0cgQUtsiEdA4wu5u7tGF5k/YxaoQJisbmvoLTZv3pF8JA
hW0ElNAhC6hE+2nGt8BgCIG9hg/m3IFpeA1Q5JmilSItuertOOD/y0ZdHuf9mDBNRZVwXKOEVQx4
vOhzV8N6ov/aXc8us0lZjsFyb2BnwCjy30VMKeSDsGKn5e+yrlXvA0E82AIqnuKNOuPXviaohiUq
uudql5U8uP5m1fIvMpC4iOkqxRwsamkEtLr1KgEeUJsLwXwY6sf0BgUNM+Uu8oainLVUA1lPHwMd
CUcYlZaKzff+1RUhqGvyhE1565l9kj5cfZJHC+k4tHDDevxy5/Wy1Qk4yqXSkhaeixu05aAQayEU
cavfmDqkvH1Zhu4WISA99fp9n+oX5k/wPLlYIkvRg5iGHo4gOQ4UEu0EMck/xFqerlevQwkvuLp5
0zdfCpyxHzmsIB+hGtQkmr1VQo1NHHybX+JZooexYX22SR8YR2fKYmBQ6FvlfScFH2F9umbIkMuL
q96O2qAHvE/JaceS1+55euqRJobIL5+FQOjWqevyxjJy0nZQcqnqDkvXqypNzwMbAk9yoSIbNvIh
8IGljH5/OXGdMOjghMCvNEfbGSBRrkmSq+NaoCHV9MtigK2NzAmQ9ECkIO8hgqx/eSUQTY+VuMvf
Iz2f/7KVPb0nNqWEFltuCnyko1K3q0m6B/eUE4KQmZu4trTrYmn5w5wsCEvG6DWNzvz0QNYK56S4
6tspiJgAcRQLLwqmtvC3r/uP7QUREkOrVVDiJtn3JlOSC2TBW8gPY/E6oifkNJJTGFhFKdzqA2/N
bVgqGh7W0/q8Ln+QarEp2RzpfdSemHcdISORly8sY8EuFCG7YbGOkB6Ify/udAwra0+Xr5aUAOUB
p5K+rAFjyQOYObMEiGtmhcSyvOY7RxczCtnY5E4MDP+s47QVR3BdHwDOAwDf7c20ggyCHujaUZt+
wi4rKtrwmml7fLkYBpTv4CeeMm5Wei+tkc5Cb7tRobPEESiMz4q7mE6M/Rr4em9uh40DKMOU/Qaj
elIYtCKIqLvfhaCSnPlxogSQBUs8VvBVP0sRD8BDxMZXpi96f3uUuM1Uz9k4qT6kH5pYotFNYXED
EvGddIco2Lxy2bZd9LryufgRXdXPg4uGBy5/Bo7t4RK9sAoxPKVoTUWTXUi8BdHgBGnmMdYBc4du
uL53vl5LqWYNdr2w9OZ0pfS8XQhEoGpzjPVtKtYy2ER+BllLuGhfAzSGvJXKCdmRb+LLc5vWa/9p
6tEOUl/B8TPqUMaNasWcr4xjWJNn8fGV5oMCOATrjMQ+FReYkkoRvJlbcpX/V/AlB+hX3U2IrZzj
X9w4pEDvzT9ojA0hYoVaoalpT3dYDtXenzldCkByViXhdRxxKNi18PKx6jfa+xVG2sOCyCTDu02W
7mTeIJ7bA0GzdwAWk6ec+ex0oB7gVnOCBd7QScyhChWlruaGPK8hWQTHg33R5u0WBajw1QQocurC
8TPKc8zd/+iXY1sOcSOz0WWcju4nClumNCQqoM4D6yUJYBKXAFH+eS4XsM6fWTjGdw2APowbNguW
fWsrkSXt+ocfSCG/uFayW2mK/RtiGf4x2OWe66gTy9ZwdaCwZ3YDWZz8A5SJaJ4gEKjuJyU0hxX6
uIvQPeqsuqHHVJslx9+2BWNUwwhW9wS55O2WuyNJgZkXvesQsgsDeWMNFLns6rxloID4T7AruLgX
2S5JQPHAEj1V/fmTSxWfKbefWgrTPZpyOrTRe61Sob25rBYvmWL0BwngldJNJWAMm6EK1zv2gi0h
p766WKLhuCXBOrHh+o5+yCdzECFhEUmMzlqGV1MAZ46PCBMjs0fFFbcJkFzyUAgb6lV3dGBN3NmQ
AJoarTvJ6Zj24xNAX8Qrk01At7+N6iDqoAl+K34hjF9j0lEsyAFwV296z0fIytwPGFu9raCS08Fo
D9uJ0jUxVJWBLNSHKow5lU1MT60HK8aRvH1xZ6LkTCSIRtd8eunvo9eiT55GEbC8ZbLb9lqIQafJ
ETjiYNzxHP6m60TMGNbUVnfE7y2FDGmmhE6gsE/31qIMznIFdPwtpxtgDdjko9B8950weyqktCZw
J9IypV+BoDTj+57VZHso6kZMEpLOPq6sabWPm9ChCWIDE5MFCLvxqTcPx8Ptwmem5e9anap14wpR
so+wf0lOctSqyBN99kJX+U6iiN79bGYDo20J1x85FO7ljlQv90J2L21qCFnKjc0vOICRGPOHgmTw
qAxUEltMZ/CQ4VC0bEs2GLSnOtT2J/fot6n5wRtErG+2WWzihSLCgCvkj/Nk4q+2pmptKmSzzXX4
npNiNF/gi31MmIolif56T6cO+7KY2kLGWroJkCG7RNSL7O43joltbnLMvA+uvCAlHLaYC4I0Eu/l
QpzC14C6DAhwbU6Fz/yTag6UIsmHjq88qrgjV+ar89fLUGjTd0J7YKcRuYqfk3bTtSKCP6J+XZ3s
mKQ1gesIqjzr/stsBPJ8jn1KhN190qqnM2g0Ua63alOKwCur9sUWYDtcQxrrrBB7gf6/hDfMAQ5G
pSuBaLdpQ0ikU839Urhkwm5spVNA8rfGUHYNZJn0/5eGT8pIGZ1DOIm0r+1d7v28fr44uBZlLFjo
J6x6AORPbtEzDSkLnaqTJ9ieXH1bQOvt3CN95OkXj9oeKtjPD3iryMl1moPUu/tXrRcPYW2kWCQv
Ayqy5TeeT9fZ/yz2SYXr/icCWFonvA6QxmMCWdaI63WhW+L0km3A/fbZ+c/sUHqL3OGy5r7ePPd4
/fXcn3oDAgLZUmb87x9WOq9MZpXQA67c9AoSNvaV7oEjhsi0yJ+4muRb7CRHLYa9CX6HTEzO/W7o
bkQLgHeLv7yxBjcD0q/xqZJJSl1u1XHqeqSLDqw585AhFlEYiA0Tm+MFbXxd4+rbVyqzeyUguBa6
wZVaw/Ug4L3iDcg4NvKK4fkDzZ5nIOll5m0QLmxbBpAXs0tyhL161ZWrB/EEFzJ+DO1b1PfUV+5a
uf/YGM0TMO5mQvEPrCslMiyQprDhHvKOEQp0Ya65mhiKw2IxbqlojQutkrwhYlsZ4gVluNFmXe/e
ZABdiX2qh3poPLv5Je0YYJJKNvcBZZC5vt0H3n2bJiL2GJa++PfKjHTdpjsJn3QtS9OjW9JsIr8l
MMSJ2vE2VTB1198UssxSuf4TkVZz7Khb974yaEAEwLCV+q+XbhJS9rOKaUEw+plshPTB0V+j/D+O
/b25QghOnE0ZA7nqOOt3r9SaYOi72MwR4sGPXw52am36fOuVUdspBaVhPb5g+RwOJEeS0RJpZXI5
CxcrlcnDWc4sQy61yIFULBrpdK5L53yEiZ2t/7pv+f+m9jpdKNFSiAj/9oLsXiGpQ7rUHKphilFc
t/GYIpJFU3gNugTGV6DgfPWqqI6e0l0jAKQvdnrGjRlMKeORT0mZiF8oAqAEZmxd0QfpAdACmwvu
Rb/0MPy2WQw7l+RiZSrZRwnfWBcWn7Wp+hkg6jsWYKEUCEIkGYm+tio5sZRb1rh09LUVqcJQ/4GB
G5pSCJNnaav0j+5JK0MNdzP9+WoEKnYsyFXD+v2+YWNSKKRzkrGWYXWhMECLtFyi6Ysp0FpmrYGo
VVwQnil1Cj/NXLwy09h33wn8GjW/6ErdqaypRa+SYPBSlqrg7qMAyGOXD+eSDdZYjeQsZPICmoDH
k4tDIMmZQ2xvd6Qsa+PDrWRiQvWu98DDdYhofz+v4rFNjKNj7LQvvOojeCXQ4dGjcvCxbqyunEP9
1ZXrWi0Yr+LiZIIwtOgulmZybnSB5jLFCFJh62tLBTHWUhRtMjRpiQHvRcj6EmsYR5gC4pr4Sxtz
+6gO1Js3ycHuqFzo5lPPINwjjqyyWf3KkocGfT4w+f9vAriEFAPDvL9INVjhVCgTx/J00dDUayEP
z2KHiPnkoICdJZ4nrj2HW24fN/NBE4qhdP7frfX9zlVXxDcFgDEpmoumFL06s0a6gwvewU6Id5Ym
JXAwRLecY71uG0TbJGEV9zzes7dVBGherl/uHV941E8Fp3uHV6Q0RC9n2uPztHoNnzd0P+5XV61w
PCdelkmlC8LdmaTuJ0W7CEuf45kjrwA+BJjt/8+GI0SKKgpczH4f/WEk+tjS4gK5d67E78YS3ha6
r09McPtv/o/M80OoPkZD8lj45S+UYAWiybDXYg/ZwC73rlQI6oYJdC6vhpSWrK4aN8FBCR359bjP
9JwP4l7aBLVzl72JFggVvuSy7AskVvyWADmXmIMyqOzcCQ0jmo3DIK9QpbQM+HEb3Mm+oyNqfQt/
rLPj0N57XrQ3xpjK3dCrBnoKVF9/55i4vkJzslYUTvpE4i1wgQxlx4bSqqZyIqxC0yXxNbMKGvOs
0MNxbBgzlSm9NgQ+I5ephrKxAQSOW4tFx2hHNt7c2ATPITgoXRxTlnRKZzKTGd0kZMMjB2CrfzSm
QBrKudekM97bG/9mnQHPWjaa8PoB5ueBYGQCRAufaq9Fps37I4Ryk6hoWe9fEIl6AJb/BiZGhvof
XtrnC5WgYG3MxDkgfgyBRqtLry0rrkp+jZe6KoCE287P81d/xXe5XBXRExy6DwJfJDN1DpMthkh4
IUZLmKfAYjatmtAovVx9HhR7tC5jylOgT/rUNPYIwF2NODfQUcws03XvORdPNbqwV8XdVdViRsYs
HfelvVxl+tmeeQxg5+SHgy21Kh2CKtXFVymJJxzI4a7xQT5nkavoEJrgEabgbhQig3j1e4gqaH2t
6uanCkmh0QuuEBCeyzUxucw/Reb1h/nOKHr4PCcjioJ7EhaOElTOuqqFSejMS/hZWA6vCZ0hemPA
RJC43Py5Bo7C7NFJ1HSkkj7jPIZOioPdgj1YU9HoJBT11QE1l7/u6HVW8etnpQQodPT/EsNHDBLI
kz6cY9oOqNDy149S2WsaAbPDpCgmJugEimfXxjCPe/uPZ+Do9XgF7jdlwi3zEfkCAyyuc8b/zR97
tbqnEYFc8oByz6BeZOEzQ62BCbC3bFZfTRfUGWbJlY1/mxmdvMndsoTb0wXlGIS3+nRvTkqHNdXB
iMjInIxbttF8zBYlSlRzVjgm7JpGubWLEWHUgyl8tWqfp78qpwf4fjAxBjQxROCf1Esj9tCcFbiI
WnTtY5jWl3Ffig6oZTSj6uyzKRpUeD6PmDXUFh+CsKKK4vK2vwkfkmiJdaH0/cXkP4nNO2m7XBJi
U9Q0cjpQO0Gd6nvohvcviQuFSxujF6yH1xTTzakDBhrkG5Df1mA2PDrIkoMFPaqQoKM5n4st41mS
DPjMEGNd46SiQZEOU1mu86vGOW5x/fQcrYCLKHy6BXSmWNmuZVgFH5AK7/ElUIbjPRaVcJG7Utpv
DLYMGbIaz3tMk2WU1vKNMD5M2gsazhZsBqzLHfYVs7kMAuSv+tl6qXVL9g2FsGkBr41EhGQgX0td
jHoc+wuO9bQFYQFVx9bh5h+Af8fzPDycEpKcwbyP3ySEqBFfCqjNfGG69WKx/Wjy29zPGDDjpEaJ
emWMNlxYWomSq4RrsJnVeWcgeLlg2OSc37rEkztQ/kBNPqh701YXsTwMRYTg/LcrE27UmlyHNKsg
DWnxVP0pB1b0NowkMRh7PokaLYNxEN6OQAogIXGdBJTCRk/nqO5JFQ9K6j1xL56wJsitjt8OOVWm
ufkHMGiBk6LTDghnrGTtww4i5bDRC+soXv+1SnRizmELCkHceZOeY8G3GWImE+u25SJXaOGBYEpo
eWjrF9ch50V+N68vQfiHvADC8CZhlpDG0Gt5hJWO49jX8bCdkBdJiAFKH1s7Ru9Ud1+uTWxhhZEy
9bE+Zp8cl+qS/77YSRgo/ckNzQybGH/98LCxWTGGUqlR+YCPmRcwWpgxZwC56efc2FKVDfz4IigQ
oOww+he41O+7kzwnDEbBT3EyhUHTC058d1DPJKVVX/Gx+FJb4prw4IurQPqIRvOKRsZg3ji0k3xP
dxlefNyasUQVR8EUcgiWuHov+/wSfZmMxzM5O/J1nuDdAXw/kvZ1XT6IBT5C38ZnbzGsbPXirafn
CJTBRK3jIX+dqHiapetsEsOFs/lRgoK0ClwCaWwSp/1gIXyeBz2TJ6BH2iR8zx0bHNeDfrJsdUnY
nWDp5wiQtQnPpfcSC9N3TofWplchjp1Jm0YcTksMFIby0MYNms+rGZ2lPgLpUcmw1A/RpKT3s8i2
2qCrBq+PQDciIrz0T9CLDNHynjp1ilMo3+wsM4mB3terUnwHJIDc+ISX+7doZ8Ki2KCIzChRgViW
hgFFYDtyxaerd2IdkYy2xrkojJPMCYaJAR22fjfBE02Kfm4/vttZBsl9U9eCtQI0x5CKDHI8q1gy
i4T2jPapootNa2oevK4N3BkTWlBG5JLyI44KgKEJdP2ZY1Koyi7GCip7PLEQDSRAgvX5+ftEuO4B
57AxZPr0QL49Jl5a+4EDkWFD3ejFBiUJ6OFJu5BGTq1lgo8jNMRbkUsjuD2xz1yK9f7qFqpvYlue
ELcxogytc1pa5OvrWP3Ur4xq2dk9UXBxtio/vWfqj169zQyasQmTCk0VSNhEz61VOC9EbuM04atB
MK57Z7rag2eul+bCgLW41Vuj5y1BLOjp36xMFgBMr2m1/HUicqk+xprnnJRhqkstzolzajweVeAi
C8DXR+3SH+2hzy75RXgBM/WM0Knhf1ohWysXBN/4/whuzQZI3BXzZr46j64ZGTzmZ9kcs3h4ru2x
xeecB+tJzCz/Qx5HzRkHjI9ENu2Q2NxsJRENMIXCWwYv+CIfAFd52WuCzuOcN55ca5OMieXxSNYX
0rSe5B9OB0+wUWAc8Y5u+ThP5ByoC0ZpY7UJTglBFaLu2lmnhnSRRXrRxkE72T1UCUAzr5CpPGKD
i2o8JP0wLxYQ3aNCxwC6chNa0xTntZuYvfPKRziJi2/D4QoXqiCvi9/SY749e4MVQjHlatBtmBG8
oxxabr8dtxVkFX4uDcSOgSEKWTdybGRpAQyA3QzhJ+GfFi+KYdx8MyEHZa4b9JzDt110LrR6oqIS
yck2rjgYdOoCqZ+Th9V9MPeXMzNZLg81/Y2BZoBbrrbcHwzzS9VJOQ/ec2FIVFFcleJg9mV9QS2I
Fz5z1zvfwdi9pBFeKHBOPcZr33iK0R/nIlaJFsqXVQByIlbUXIA/4vIijgbpNnkacR6RSeLVJj9j
uHc8pWpuSQW0qvLfeWqwOU1Xt9Q8UO0knhN2w5e+pvW2mL2NJ/GigHVVoEE1pnaRCcAr/eq/Mcyu
Lda6d5Bgz8I6mhJ1xcll0H2stpxspAnrcPHKXNJIPA238MOxRjmViuJ7pzvWl2gfZwMA+Ez85wyD
aIXu+QIhPmkLEiimtrOr50L3efauLrpwwcfr1TWwiG4HgLiI8cklOgmn1I9TOP76AFCMAKE9NzXQ
yPqJg2o5S+qn6LodfJ/g1ulww5VL230ffazO4Kh3FZIjfhyPrh2QF5z/GZgpjbGbNUaIBWQorUq1
/9gusClxlHHY6DP9oHqXGbg6XJ59bS5hnfrhmAx4Kv7rR+o6wL7hkZaaHJNd/r7X7cFPPVCqHmCV
v9iYVTSddTp0wufTv9Y4NzWElo+RFAnxgFT/2FXrIBg6lr7a3KDgEHxBOC0Jaqidg1XSDEalzEFD
6tYTwKwS/292uNyYLzwmvuz95X1DLXiAN7un16WZLKR7rnpOG7UinbCqH8y8BLlV18hluieQhWxl
tPd8sLLkfiqqbOsRtruyUVNHWcb1lcpFq1J5awAnN/2oBhJkBMi0sOGGvcHiIZz/jW8EY0xdMvR7
X1ofjwu1KSzAzZ1JDjyu+IAuQZnqRXQZz0aPdFASZ7znyWvHBk8RUvLDyPMvZsquBO/X5rCnMA8t
tbFxnnPJu+P3F29dKy4X6vheSdbV6VPctJwdbT9dba9vUgOmC3q9Hn8m77xleQaTRG3uEWs4VgDE
mjt+Ac5iOIPS9aqJ2GN6OxZOpfSMLzEuvI0FJmEpq1/AEITHft5jxed+MSdkTTSr12/Ic3CKh4kk
EAcf0LMNCufeoUG2anqY7crcvxatYVY28gXrmuZDjyIlq9jXi2+9ACJBzeSzM4QKdQaYl39cVl+s
La5AGDyIORAtwH488wzrfMFPHO708BYmr8hCbPvPzCHdMWcFGYXbeOIXUFIzlDNkXaFvXuAafrYF
yM/clYKoqtZRkja/B8H1Jmboy7oed4+SEp6gz/oowxIraec27fcnu5YKjYLMYH2dJLQZQAIXJG/a
qqsORmiURIK+0EASez7QMGFEJBmtgSSPsoaEVW28RI5faifC0mj5zdojQmpXBSLmOze7lhlulEzw
Hh1J2aLfW19WxfGUgyu6NpZsx0yQMdUNjopiPXX09hLw3P5z3CaIlIRDsddSK41fYn8OdfrCLIdb
ng3cSj/IJd3rufVdaoMIVzQil/hghSUldK010p6plbT1x8YYKO1VocKBlJ3+cYSvyDM9Hl4hINMh
n1leL8jOYEgnkRiq+pq8yPB9zeg3QRh/9FydWOOSEhzZYUbELGubuFUJFprChqQqyrLk+AuzHO58
xHEdlxfcdvMbh5xqN/WQkdnSK/m34q30SH4JuVjf/Ti8l0F0DX0nMjRFknhtmPtLLEWoiVNxKbYV
WVvnkhcoAKrfvq8uhbJWTmlEYmTY62ofFWesCjEwmX3D7Dvu6va8oy+abRWt6d1Ga6cziQNsdVPR
h21N713wm0IxYO22II5yQj9Cz1DuMK3AlH4yIcgfE9hpy4QiAgcRmft9s5jrZvw4jg/siBbHkDUz
U270qWVhg+EPWtvh5BieYCn37VcvUv/RjpuEoLvGC1yoFluwySTjKOxhLTYLAk20SEudhmuoIPDg
DRFnTUwzGi+UJEVLjYX7idgiTcOvCwSVgLy+4VbTXea5oSGulcr1/9VZesvak65sgAZI5QOWpBAJ
rZ+mYXnbKC7d24zADQOu2UgDflqozLOPPZIF6PQvKo1wqSzkVGRwGfNu705JOW3TfMTGbcyKIO43
nvpB+TfGTJkcgDsIa//WoVQc0KfepQZc29KRDgSS4Bpiobf450khOLDuV5CN18GB5SyrNwIKQp8u
fadO74Rct/nxab5g6XTtn502gzciQSPkGyFkt2uot7Hpc0Bh16tbxl/sCwmUUB0FKvUS0sjJKraL
acIZO9TvjeKTBGNCwbj+FxF4/RvZVoMT99639bPPyDBuIHjnP4lSuaTWmFPGKz2C6Q8VroeSCXge
8DpLYGpWL7gudx7OMp06k8F0pmeylqbgdNWwd23H3Z62Aq/XvxHZdhMzR0G7Gp54a9juvUxi2Qfv
pWWIYEs0511cjpRwLwqIXTk8+A6hbmDR1VKWpxbUPatPHFcyWeSKGk7QM3NYXqaxSHg/3irqiUJ3
P6HvpyPZkJHKzRB+ETy2s92kTGEKG47zl55BuihEuqfZvIUGViLyHXEmPtJ2ia8DV9+3krrGbP/H
mOqdxMsmDntnvGX6zE4mcV0nBilF2yEkboEN2t/tZ2xmtS4UDY5CS2WBnvgsaOsnVbpC91VUmhEO
NuFfsEf0tXciTqhqKVdMCrSapzgX0m6EQllayqvdS70/b/nyJ1xVnR/aykNuG/u2z9JRyoZGDkpD
OFzED8ZrXScPwIuKrVC2BkZg2jVUwEMjJi5M0eepib4yaZc1d6NvM38Z/L3EtXJi1oonOVLwuGIS
LodhpkzM0cmT30tLaRtKEQME9ESu7GVVQPcBM28C712dJ6ojKr84uRsDw7xRLtyKKaieTRskjpxW
jQ2rJHxgsH9UlDdwUkRJZcC+rZqqabXsS9yH0Xr2xLbqyFBzrDeEmg6GKN264u5YZodJ3WnpjjJx
FqtaX7XQepE/WCiWpsiXS0QVvCdIYCBnupc9tQM0UTK0ZB3p7lYY1gdBHVr4CSGohL382lW7C0MG
ucmUk2VMmGZVAf1IIyT8jaKNlkCymaNa2ehsyRUZOg3IkEZ1R/k24rhcVg6vtafi0WvbcEq6dkGu
/ndkM4EYk9jN+aLpNoR/xlYLT9BqEXBBcTc9IriA9K0ks/oEOoF73xuCdRlkoqUlwnCUXQ5amd8a
iow0c5CfQJ6mYMthErRcJXMkxGMUr9qI0MzLkHAr0eN0XWxIL7xllBYTehCV+oE4lepPp+6JajcO
a1rzyuxzyONBO4WV2cyQfOwEWPHgTPcUAytYwpSuSP1gVo8CKn1dsSPUECpN80rIGx8AQwUN+OTZ
+49mqtxpfpYFM0MhNxRiCpmuWATY8FOpDNBOM0Evg+7iTfJZQNiTZthTQOZn1dTJuwfw3FcFatq6
S55VxK42uyMRpBmdZjNJuMOPDBZxATLetbZHJpZsaG44u2Sw7B/wkk+dQmCvNpJ4tqyZsZ2SCACo
FwLsg/kskwGCn0rKKmedOVZoZXlMxx6s0MZPmDuNDQIsmeTpPyFu9lJC1ZPmJcOgtDvu+Wengu9l
IyEvngnvNgz4EG+iN8ka9wMwbTluAQvHJza3nuzNwts8J1GlJNxI53WyR7xhlOe2ovPShZ+oJy/h
3WgTpSxkkPbBKjVSZJSovdHosmjo6V3CFMssaUu+WkULDgnj37g2+AZ+bhcdhBFg7PmJpmP0XKVT
K/KU1rMXVXq57VMma4oFjqCrerWAor3dZu+/s836YHaW7Myly3iNjUHzoqQOIFfAUb7zHqGAeUBN
P3G+n6mItSpNJjlsYbnE2gIACrtZgAmcje9IyCu/HciQjLmdGySvClVYEZu6skuPGWd9bjdOyhas
lUV+WUzsPR+Gw4/XpExwoDHuupOJ4LLFbXDstloK0oTY0Po4SVi6Ph79Q4dwbuio5IPSN8O/hfqH
UhZuMvqgI9/SSGj/Fnqy+a6qIwPvd1ZfKoHa+gH1G1DBZZJIX44TnzAsHWD+CctLjHtd1HQ0xplO
8qPFDXn16+Z+1ZVrehXBfBI6+G0Y9pyG3FqrC6rA73uUZy7DI6Ii3kpAyxAbk3L+ERiVTnGeCaoP
gCg4mRoI/SWBH31w9NzmGqEvCkQYyQTRNteM751uoFb1W7jF+li+F6CIAFxXq4te4JXrBc/xvMPc
9ZnYVeNYk/q5EPsU8tlKI37T/YMRAT3CRtLQC5zHmJztdbU5RDxzYa82jA/A8/AUlQTDFT4dEjXz
mFV4EM3P4CJ0oOlalyorq1Ucsl2oq9JgYGxSIE3mWNOFYMRXjtFVT48frX6pwMLEyDNfxufA/9YV
cEpgG/+wqSbZNrbxLJvqB0eXM8p2VfdvbOHc/c+3f7XY8AfPbOteLevAS3WQMVJs8rRWED1oucHJ
fDMSsq2SeOhtE2BUGbMb0LqFLtUDO4kPXBO6ued3nqBWfeNsjJmHAa75H+CcWQGwPtXMqHbYzlRz
0ZrtZfmKrOEIqhJmWejJU7WerxAOY7IUw9MeN5rSLfxQ/5VYjKkemqCgVTeLMHQ3M4j4CFdfreDz
ofRGoytKgF+Y7YlvFjFdFrbcABe6EAptww+DHyjCCYu6xfOZnq7CeU0HWg9RtrRw07D13/DR7QZB
v3Y9mebZkQxWr7qw3kHRey4O6HIUhOurt6UWNZGlOhk1GWeOcEuzZx9HwoxavBgWOv904HX2ZT7Z
tQMRzyHvis78o4j0yQYWbObqG46uFfDHSltN5UMikMb0eY2y6ChG8yAsYkloifEOBpt+TJ9XXmmo
ag52zrgt2+tCAtOVJrFR82X39M99tPrjQ+pitw6dj0sqnB4b7Btxulc87GdNM1KVQbQzJ4p0fbzb
3RQMvHPV4mZBT7Bgo/DPSWBsMIawrOIjffpyqQipV0Mo6VzH4x7PPK5AN7yBEQ0vQzP6dY+7cyBw
pz9qs9FEm36rdqZ4QHQDphtdaWiAUjtWUH7tm2ppbkSgWEfmkKtmaEi6hKx/VYv0TrUWgTHduLZ0
9ZHY+XTqusROcpPxh8NGb8bhNQkUolImhi40f85qwL//55lDLQlmLni4atBRKS0VIw4GQoNRSstl
IVaMwKH5GI8npQUTP4C3a8bTaZ8CM5ObXOdKY8UuAXDCm6UumnFGJ5ZJrdfwCtuFY3igWrocgwAN
EWnhxnXVFc5RmY4GZ1dm9BPUzpda6QWRUsMIKA+/JaH6Og+vIyeUPR9k9ZSJnaIQ45PBA8Bb7hWB
KCF6F/KCv3Zh87i2Y7+Ht8Nl9ANCk+u66I3fVIP+eI9ZxznkmNySMYBrka9Ekd00v2SlEbkwfmwG
KmcvXb5O7O6xrp9KYOkDirOORznT0MyHNhKpJMe6pJpYbIEksdKh5mDQFqUOzFHdTnx3yOdAHBxt
wJ35N7SqxVoLQQybHHRlCpliXxb1xdnvrpKYs6W6pYLlDvwICppYnBM71SfyMpwzJJgYL13WB1Ji
yy/dgWZxa7zgC7t9bg508SzxAgerEGKXGQ0pHR6DdS3WIHC6QbyO52r5D4HC25oEuIZkV2pfIx1A
GDIHIbJYtmSPaZ70DspLZMVtyohfRI+reNe1DlNxtaG0/mJuW2l6NdHnXvQMallGgFd0pbn93Yqb
SmPi5ENb4H3GVd2c1zvcOy/Bz7LQFD/5qT/BgFF/LSKJ4bzyioQMb5VIetqQ4wSJ3DFau37QiRTa
cc7ILJlxFoYMVWABx+i/+UwRVaEElke+thcjSf3QAgvp6hsjh96SBi9XubzG6xFRsovqAIKWecAK
E8W8dzKR9jrhd9lG3+LE4Rj64+MfQPiIMH4hYX4o3CpWiGNXrefryGem+ucKZP30tgGh7KUZI2x1
9coroiCp20ERIPmHv8HDcveSuwvm+NakHdMoboNGr0xKjHexMz29Gv6zpCIHV9pa1XRckIqB1C8c
pR8zykSiTQ+g8mZ9cUrxI37ktOURE591DAhuLGguuLZzL/jvyBqT1Fu7cSQTTzJkXc0xzbtKEwdS
/WXfjiCnjF2kVWnGYBEjiXAtNPOEKxy58Y3Wu5SkJa2yyW/n9oRv4VnC0mIHFagX3CHf3NiqOxRt
+1fpIoWmafqJ4+HV9BF9c2L5x2G0E71KEFwB7NC2zsVTHWD5W6c8oLgKmTDf3YCD7OMOGGLY+ag/
rJeSeMX2l1fobgX2SH7iPhnu4Xt9j50kiGvnz0eVCK7+MhgRMp9sF6ZYEHD8UfIctMpRm9b2xdGu
FRwdupc+6ZQDqtnM2s1qXMYiTtowGVUNpWXo06gFtSO/nPo8BsPDzUqQOrzgjDUd7pBog8dRIPfU
ftJvb5kmmitoAmhCZc62VusCAnoQW2O7uOuv4H1LF1DOSjjPHO61/dTRvHJA5J+rNXssGwmEdU06
3bjUOoKf43DjrTP4uuyt5TfPiaQMli3C07eb2gqJRohaQpMeWrv0hqOhq24VmcrSyzq0n5D0sPJw
dSGsKrfw7TbGMOz34JPZC7RxAdiTQtRtm1kLrG8omBjviCn43uGDT0X7vFfEuxJXoR1srkyfKTsd
yj/3eoxJ5u5FOJMWWcayRaWvmlZM+xaMJNqw7R4Y4dQRSm/QWQXqgMfPh+f6QFtZL0+liEf+pOXI
Q3au1HoCx1KJRQJPHRqRt1LwNGYDqbeA+LmaOxmqxjBlNKzWtyHWNUdWryYQKWyg/VAoOx+oEEcM
elRO2SkkT5n9ssROBxsXEOQaO6dyI/tgvyfrlv7nlxj99IBYhvYOAQxHXQuz0TKO4rANfboujK63
1eTlWgobdBookHeNsK6d/lzZnxikSzD2b829wteEMsjGwiuOr6LOY6S7cMryoON1PjrThCnKpyel
Ycu7WTmvF8IHZu1Qtc/VQKhNa8RRuQeAiNp8qQLYnvPNc9+39ej3KN06deBTwIANSb0siJDJCBJP
sg9krucWinT/QaKlMrngAteplFEic+e1X1gEy7dwXhiXHgIK//nZ6+QONdlVavcowa2valEeO9FK
ZXO1UIs2d5Nk4r+KKbFgdOHG+LqAdoDhNaWm/woYuRFG8Jc6U5/F6390iYqCgHT9b/JEfpDQRZ1u
imZt2JuNVuerg2sqersylZgWdbbIWXJTCCg3RN4M70WGVte9K3x3YNr0s2Aao1WC8OfkRD2hMHPq
alu3Cf6IGuNXZJURbTVGxSo31ncQ8oVNksiCXRJpeYzBu0e20bdgXRL5X7ai5HOaxR8RI2Ov/NYE
8PEoOFfuVAHqtp5X8Q6A8DoAWQcb8NRw8Xoii6OB3G1d2a/9hpcB0ylgZUHjJ+CfeI17xn/UDzFa
HDjAyBVz5m+anq6jvXeTESVRIuUePEoXSrocaNivswxoCzsybML6Cx6FxbayXICt62Vkx9rTaB6P
IFYdrB4d/yiiZzTxNZkqBYus2MXnaK1+NMkiz8xu+wCrUHF5nFQCUGcRgAaSZQYbYxsWbfJe5Bmk
F71ibI8N7JitDsEcpzIg5NYRTSRR9CDLh2hXTZU5b1OXgLNQ3Co3OM9snLwZ9EpB4rX1eJp64Iy1
ipB23RNWWBOzPcreTQES17NU7JMFgJ+a+cAsnY3m+FMbySBuLERMxUPzaaBtUQbdu40/dqE50C0y
t10CQqrnaR6t9OgRhRaUbYa/l6qXGexbciCTcB6NWPV2ZhF2dEdYqaXEcsV1phOT2FAZN8TOY2Xv
EklekkHLrba0t0lJV00t7dpr88U57AvpaXgqf7FE/lvmVjzMihssb5ap3Np0fTUszgoUA8SgSYAt
0sG22uqzLul9Kvv9sbtudqTVSjGYPe6ioEozyTJNihOuLkbTZiwVEJZ/SKxTRN2HfrqlgCS4c4pG
4V/O/DW4YkZFv39wmuBd6Ky7EAmtlClrhtAssABiLaOYd7d4aRPCmiommDE0m7TG+o5Od9wDyoSR
HYqhGtL2nCGptJkaT7/Hid4yWQDoaPFympaAkYEMPOJ2YywDB67CU7suzEE5FAwR9WEfHMuJLHla
qBH1Sa0rhiw//3hCWhWd6Ld12bDL2E+TypxzchPHAt2/c0nlQUzHejZSmEIu/QGQkLPiV/2vV/Bg
mQ6x5OS8IJOsujwQuNmzWcl53hvElkBiN5JSgzaHuD2nYyjLCyjj9qRgBtM4kFKgSEWkIAFR6Drm
0an3pCgyw4C6Z13XLmrM7Y+Ik0Lm3TkfjIuYTymdVK1wC+zJJEZjaYRyU3DqpQZciyOL0ZQgbRVu
F4bLpxqM9uoS5E4vGtMJYrORtYPSxbJ7kfByOtWPZPa9g00AFMxp9RMCVqOeqTY9C4fJiZJr+EiN
E4LXdRQp/zF6YkMhZZbBSMsff+sMKh8WTKnP/oVLt2XD0SEMcXyJwjH6gvYiajMJLYZnUZ1z7JY2
Ind/q718i5pdTTokFpyR2ziVwKebr3k7UjMBTOPx49ihWlvRlUDHm+KZbdmZ6UqR8cFpvyNQs8q1
bdpa0Sn4hTf/wo1Ect40jcM1xJ13gTOJTGIIXTnn2afrX118EmyZRBsADBo76nAZZBuqrT27fHm2
+5URlZowUmPwNtkMUeaFKvAVY1M0BtuQ/rX3z6+k7oHVzi9YBDPx2RyQMIVZ3kzzlHBypJmiqoYO
a4VUFy/y6lXc5ce/04wXWeEO6xhrv9zEzwEm3gP3xGik/xv1E44FSn9imYPJODhg7+lndnPSevqq
Mf2CBfOsg4nlGb7PS/8Hb9J39rnrPeBPUV6YYQ2lr9Jfrdh8CMAxVe2KHTiETTevRFHm18/+PK4k
LuWKCLxD2ncrTQ5rkk0GsHB0aUq+WWWz8Kqoo/6b2MpJB282GrCx0lOOLXv97/nQlTTX959TVR+b
/IiHuvcLe0da+AqmUVYUCLhkosbQhKctKB7nlpNSAjtYWWzNuQurn0CG9N9bAjYmQzI0IMkDJ542
wDCNmdiOWtVhq7nubV5JgTIUuJu8lQt8AJhYdeBPp7r1ghK/CXYHtJizYufsKG3Qy+FSDBeLFlPY
VcuN7Cx0RmpvSgEsAupTHyBzK1AaexreWlyWHHtEa/hfkAGvmTlgpZC/U7+gtQeTAL4uKbqz0byU
3Xj1hDr5EitaFHk20l3m/Q2yzqQJW6rx0OlLUqT+NDXINNNIlW4MiVCYPyw/TVzimDNxnDqb1GaP
KXe3cptibN4n8Ee2JbfLtfu97fg5++9gqYhJX7HGX7FucnwfSK2IRErbtjrkqcWWSJNfv5QyDNas
qNjeCqgk1DRsJd1Dm+PKHzz18lmyXuRMeJiqSq+/YrfxoBv8qL2FdTmjpz6y0GQiCyH7WAOATxWr
+6MB8elHEsuN/o+ZuVMza0Tli9kg6xlQi29ryOyGAB526DsqVj88Q7mxhlyIl07Pb1wJkDnJzMKB
qDilcJ5AWTcNL41rVovWvA3T9hVSnXjD00fmNz/Zo/OAketZGcmkZLN65zpu5wjQqdAiTG2hP6fN
ln/f0uwN7VMnDktOTaM+Mn0bT4fxsYnVD8TCLqRBsXvOrvU/5RG1Q053VLpS04jEhmVx+hdhxebC
T7LRR1WDY3F6u/0vXBXJGqYVtYKY2fPzgO8FU+HuxO1OG+NAYcQ/kIKlrWSvZjWHCWGptDF5P+No
msPsD9xe6ePEP/vQz3E4KG5rzRKg3AjWvbuuXiHQ9nUJxE2W2zT2mmPRL6HT1fNTVZAcQZ/4iFDq
ui5myU20WOLXTLyIwZT1pAxMc3SeU3Y2jOpSCFSt5As/YSEA7AS820sSmxLDoOr6Mssg7ikhpGSW
HJrElbwZXWEStr7EWskiMQ4alFrEGkRnbsCiXwiBEpRSs+2z+wUHCc86ACMTz0YPloIPulSZ7rus
cY9kk+ehzoaOXMgaH7WESbuv/HlRgb4yZ2wsEDkcxsxL7ke13CVpNi6rqYELC70XOmOUYMcV4BWR
XysqZsvtCiDh+3p5iC4o6C0/NyUD0aMO5iQ93kvoNI4HUjHEc8se5R39DWnJ9DHcaMPmsh5PoEJE
iA0J5uQeM8tVAtUpeYj0Sl3plufN5S783SWgid8G7cbnkQ/y/fCcroE9OeFJFYIkidCE/i44WALa
41OzJBWjBDJzwx1s4saAxaOwhcFkl4+6jE4R+xxDJ5+UTeGpSPd2lr4SKqhdSdwdqh0qb3VMjoAF
11czkVQsQevaP41ZlI8HajLV7Qj+5gSAKmH2zWe1YrijSIivrhMWoTSB3nURzJNufg7LMiOqVeNF
TnmsRPrEWmsEFy+GQe5Yr2Y/Xgj358jpdkhvtKY0K6WPvNvGIasP39SDmfwkz6ZRlWX3EshCGDT8
Nd/NM3yBt0e5g63W9P+gvPhU+c4HTHrNQY2qXx/Ypl+edBUDGnj7iAz0ULh6JXEDY0fIu3r50Zkt
S6T/fMrMfbYedtjJpLlrcZYxkzmEeidteUwHAUNkE5tFVn3JNE9T8JSbR/gh2SS4AX4uvYG9hqPJ
z2ic2Obnn74QDoXmjM3LGpTrVUK5d8QJB8cI3zq+SvHVBi3/uGgkkydhxotkB+wyIQLYEUKmKS7Q
qx5zpUBT8W0YsLj3LqmaYnRTo4rgOFZ1RbjfX260pGruj695sfGuPRrBy+/H4NUrrvqs9wuTIOyz
ymhVfnAwgnGsLcE8I71NxM4UZuLyCFRLhZF6/eAFPSI0LOcRQijslBFVMnWhznOjOTebH+z/czf0
ftYvwh4SCvF8g08r0DJOTmH7j+PsY7tbPryEfuFk2bNT0zmmSIaLK0WDV7PfKY3RYFEpXwi/05o+
w/cvETOPio57XgCqTE2wiRVXfCbbqfcSQnMdYFrfRr22WX8asbd+ras+uBH/xGRxJyT1Q6c4qGVB
v0raX6flQzmu9s53Hr+ZskROtzCjtRyfUSchG4r+W5See6B0Mk+4TQZPF3BcsYE6EcTTxPdN0RHH
x/ey98Pb+uhVsMOTT5kD1qwbrkLK5+lh6E5h6o3n8ode+j0iwevzxLD+VffqzKnWVnfI7rvWW6hz
C23JAUquTCoKw2eeejWBuW7ocmF2UjEIr+OPq3UhNcAqqywK9OetOYph0H84UD1JwvR7LyUGalXw
SzE07xdoOYZsijALHyphHIt2t73FNwqdTnaULdDnFoyPb7oShzsxyqyLo7+BGXu9BCOxMqz8q17o
G+A/i7Cgbgb5aF2Ek/JUGHLgk+PIAqXOb2rluDy5HEv/WRKCMncb/flNtJUaGam18I5dN7F1aZwv
wva8LJZhXulGZbppbY4JrNHxPkigNwRawSkoKHYM7IEXsXZfFbNbgUDtKo3U9RthhUEXi4//4aXj
tRKR85LJSxrEjLa54xDgba2NBseuFQMXWi4CUTFFrQFnXRhXajEZW8T9J755xbtIVHpuq3IglE7f
pJpbf4BFjIe1SuSJrQv4uFIxTltknngLn1oDAlzIE252d3+1vcU8Vl1n612sWBIU2vg7DAOu82+w
TWlRYAr6JJ/sYtLtbM+hQ9iLdmqz8JpIdeKguv0WPhxwXHMSz+ijpWKp+1RCXQpizJGVys6cP4aC
UFyFNvfRctCMXBZQExoTOwktP+d/fVllQZBGJQUvLheHGMjP1BzBic0lZE77BNBwNV8EbC2qZ0R0
AkDq1sRy9ClC2WhnMHfVjFPKslOB+lhBMYNfVNtqwO4bohHI2qdcuV4IYZU/FfNB/7XtP1vbT2Fd
mxRmgs+/EQUuQY9WwOI2qmVXVmAfLzxXEwSrSYv3vqO+2PUCn3iDr38/zOWMg96qneEPDjc/oENt
HJLS+tGcD9aGoUEkHvMmE219RqFju4+Ze9O5KTwPEozpgsQ14TlUIqTmDe5nySg5rrdBLqNImA/X
rmJ+KxXHhx0iW1k6eJ8ldTfQ1petuQ7lfwZbQojxJETea9X6c3C/mqQXhmLOcggpf4aYZw2Bjb95
8jTqOuAkWggxyhpayCyBv+fXcHsyfGhCrNnFJx0GbvMsWHFwtFOYFR9B13KwkByXXuczvFkw+K8y
ntsYZzoDaH2HJxUfhcali2r3/GR89+Qm6ELHYvcYER6B0n0N/qu4k+03EOXNgLBm75S2vYDJi2V7
kZaq76sXC+pqvGvdAMTmBk80S9p+dZ/V9wcHIfQtFIxL2fjI4qijM4fBDhZsuBCpmbJdjeKC/HGo
g7+wcVz0CXlOgxoAu8VCojMy422ZZQINJgzH+/tHJFKVe3q8T8I1r6zaznF717ox2JTCUZlLFJcz
BqgEPEtnDOOsEanfD1YCxJii1iPUNNe4hWh1Xl+o8fwvgOq6LzZRjVkj06gGPt22JGjq9QTPc7vd
pCtl/orgIUnUnzvrCZsFIOGEvRtoy3Vs5Eu8M12v1TgGdZK+ZEeaq8ylEfNtwxrTU6wbQqJjEmLp
AUduc4wlQjwCUXl++mMOAoUXQlahBtaqgUeccTrluXPyrvHH51umRscArV/3Bv4BOR9R6tZWowik
g3wnKlBvKURJuiU5BAPMYvgZ9RivZQt8x0ztSKSEyxEU1WDJLXnoDjxPiswHjppCwy6YnSotxvwN
eij9UUL28mv11OjFMJ4ot43DSlfAAORGQt5p6i8x69M5MDuLaMbt9e636quoZnCiqud/UwTW+uh+
6Apvp0tDSdXjtSANvB+9mKDx4Naf3nKqS/5nKlN/ZMpH8swEyGorJ/6qIabbXo+1ZFvuZgUWNE1J
RG7xuZdHvUjkMm2eqBPAomCXGuKlNMzT0zar2BuKZY7h96Kc8dsHJYs34pmbxhAb84Fp7MFhE2AK
dcdyLrhEK6gfPt0BiENfz40yu1xEsB/b5VOSCB1UryC+Gh555bd++SL9MuDhF7N0gaIopyqVgaHX
lMtQlTqtjoUorHOpA+LwC2DMlezgXQoFxxxgJEryyzN3IUA1zVEqLhBGBsavD6DYrU1Ich37UyQR
WX6yUzSaWHUjE2U9fOC1551nMFaW6PKn1NeQAzsX5z0qOViV3YEx7U+1Bkv+bgZz8yjJtipz9SPC
tFszobVdTTHko8lLUGwlMMGlR0NuJVu3GC3xZvR6b8jHCCMnml3FiOZ3eW0qmtZMaCrHwvvL4sB1
9PRDkizSahTnmbEUrCnvEbd1l/b8cgbmlIDalHzsu70wCNDemJjfRcsEWvH/b1F+L8JkxfaOo2vf
brc2b6z0thf3Ovrmuy1ZIU4Cng6moxnUHXnipxfjhjEo4PLHbs8hMwSUGPR0tBW10w6vUoSmJohN
KDUPVOaWGWfr+UEWgIm/j+nc9hVmaYNTOU5+OrBi2imQ4gvg0RGeVaaeKUn6Ble9v6Jl3OEf/S5l
q7jQ3Nz0pBLyCEOPph/fbQcf/Z8zkjsf4MMr3a12oMADojSlIosFljPGcuK9bGJ2G05D68PEXUtS
nHwjMAbgBIZ2BP8OvVVUZJQ87llPTyv29XGxUX3mXAJJOlco7Bqd1/ThE7d5t7ZXWLlcGRmT2LP3
ZWqobLCXOsvYJvZcNE36SL4SUOU+J5gkULl4yF4uYIZ5QXK3MM85MxB1Ntv+23fWX3/DgHHFIWkd
9LF5JWiC0PvATdR5LhTGnQMzqld9fdWWt+C8SI38LqVqoyLxO6ltqRmqFVwLKM9s65I00FOe8/sZ
RYP8sdePewasfFm5H02Xmlj51o+wr1e4siaJ6QVKe2Abt6dvQbpsV/Y/tLMVSX4PdmkSI8K06FG+
KY2lCoUA5I+lp4vZxq+d5RBr5fAv+8yvmlic8M0rZF9jjBwCN2xkcbxBLojpaS5bPwhRVR/d6Cz3
qQ/zVc/8fqftjG7jehEgaldd/MhAOzeEDwRSrFojzniUulZdQRIv8Ydvrqd8uBeJIuKkBPY3ucgE
GhiFA2mMuHekisBbmu+M5WSfbsGqf5axLCX50cQYHCVFrnUsP3b5+z4zBcEnIfCpluNKWiJh446d
UdKpnagRjDH4hOON52xIGw70IIOmCtoXgKsXK/BMoYeazxy8UnwNwJKKPInBhyHqVH2uzfI3sJRE
PeD5YmxFL+EXEyZCGKCPFXAvEqlLB+49GH5KAcWzc/3/8dvDLWdcmPb+G01GUPJoH9xDNQdQjNfR
pieVFYciey/theD/zyZoE3sh2LmEjPlmKoOTnX4FnL90YwvLyBFcV0czQ69zsI50Uj2va59nwM0i
YJfYxrHgjtCo4/6wd8H3Rh9hPZQoUJJRsy7BCski6gPkL+Lh1oowII5wRDtTho92ZLppShzamceM
Dh65SpPCF1p8ywCEVQs7OElkCj4aVB6Z/YX0cki/z9HGIhidZTjeQgpEQYIV6bZLwwsv1uzHMSim
tnOPPfKqC5AnrlGCfhpr6Lw+QcVSejB1p2gdntryj33+1wZMAnxwThbDI054/bYZOj+OhDmyZdyk
xSb7KWlpndRJP4M03Y9lzrXedprTwM0Y27hNuCjp/catiGeMwWz0M0i/puZcmTEaAce1m5cVN6+Z
Sude3qnF3ACfJCGth2OV2hahuym0bEuWv4hn466bCAySKwjzkySSIZP/oFgziU4Vd/8wy35o6YbR
igUXCWT5zoHS8vNGUeZA0auFKZyk0ovmjmhF7ztxJMFZ+0btu+SwjwvBKpg3aFj5d5cnQsPjtkoB
6oyFFH+Nh0C6jRRYYeinoMJVdc0N6/kubDco4VW47x4PqzieUwgUZapXXlqZFEAQijcoNCdAIne2
KmtYp97+zkopE5BLQea45a+cXPTxVFgJFO7iNKxuqLc7aRxhAyO8Ei8tU2GWEA0ZiWci9jIcMp5V
8ldPTlApVhlKgNh6VpewQZe5jKPx5ZK3D/grZ6R8EQ4PRaky/H/1KgFZwo7LRqYN1SHJvvZ/bamD
m6vK2NgvwcXKMK0a6tkxNpD98/liTBhj8Of5rYUHidVnS4tQ6rqvf8z5/Ni8jF37sA+69WNfEAd+
tgaSHlY9+t9/nIhbe6/MYzvhlNEQwhZZAFM35w/INxqbxkAeM2Z/gVPui9vmUtkpzJIMhf2NQjLM
cYkI7scRp1lMmfQjfD4ZKzVU8v8LDlxQd0TUadbaMxLT+BQWf/NBeM9tcCK3RfV1z953y8gj6i5o
cuPsF+zeou+Yh3Qi/y276aBrDoEHsAT54L9n39iM9aWBpbsZqKsNMTwcX5Qqj9KDmZWNqaT4mj0n
wLGvegEzeoyM8S4pjH9jbSwln9DjEmyZCsCazjGyYLPp1Tw1BHBIeT1IHa8c1Ihrq3BwT/j8YFwS
ngBW/JpUp5BpVASLF+Fwxa1DalabX2RMZpbwm+Oc8uVZAsu8kTSzZWbD5fdTsEcOH+tnAdRzZcEQ
csiRSE37Lxm9pAVxCPggR+wt3YKgG+a8/z8+axuqM85TU8eavYM7/cOlwbRRysNBGZrGZnulKuVQ
W90kotlCP8snf9/+ipb7gErKIlnr2Jx4d+gSKk3ulSpwqeUicgBcQqj6XCTAZ8P+zYHKYGEfU2rE
c+3clFfME3D9ZGLiGuTHoS87Ve/hlPfxBUeGKU16UGc6KJw28YO0tiQca4uwrDyXZB+sJgW0AC8A
7HSqPCM99xR5gC/5JyDjBVZFLunn6EC7hX/MCy96E+G07JAbdg0LDNNCuzPS8KTanpFMUl90Am/h
TCVWN6chU9b326VqpJQ5AiOi7pYLbtFFzstHJzLgMtCdgPzo8TDzJppGKygVks4ldtSE3kZESRFt
evLnUwv+W7MA5wHk9niVaTDL4GyJtm8xLoURWbci11qi6oOfeWXEC3Bg+JYqNHPtUNF4kyUNVtI7
pry8/yWQ+qJow0hdWmqP7fPNCe4JSQyDoyVs1dyvQlPpHj0mnpTZ/dJ1j2fL1vRw0NHS1m1+vAX0
QDLXQtFtIwfEjaLKq/u3y6o5MLdwDgyBUBUfKPruaRXdpF56BX2PS6R0xHcs5Q/l5JGxUlD1G5C0
UWb8kHpbgucfkzA/9PZGH5bSt+q2BmWF2UtzZ5nbiX+96u+hYQSFC7LjSj7TqfUqToMpRLdDwfty
QjJHmmeZ0eyMOSnF92fqt2gK1LJkBdH89BfjMw3k9XNHEM+PM7UUdPOobAVnbuuuK33izMZ4j7tr
oJSb5DS648LHgemtayGQLGZC4broxU+R1I+fs5KWh0Dl8y5oT4i/Vi2A17UppzR6YUNHaqk4LkQv
BWMKCdAs1vebZsn35PtQCg/aKmsLRk33FKDOvYz3efB3Mft5+uJQjOh1Pw5A8BZUMSYBOy0E1o9u
TOkh5KfyMVEAc92WJqruskCqe3QfbdPlW/inioR+bts89zPwKaUkxigte6IiYIpY0rblqELX3Mss
xPtiLHBrtnw/eBDkSD83eNiWBHzhLsj1Tky7t61AxFQdDi/MLKveKYiNwSRTSwnDgLqpP68jo21I
yiLfcK6za26q3mbKUdO3ccwwLAWst5oxN1NF2S9C68zDngNnsvhch/at9syj1sgwLlHlAE8MrvOP
tPIvzDsCfUztl/jYhgDTnCd78HP2MxEi7zjhy+yeLYcYTwgpqS6AXvZBiuPQYGCR3X0vJy+QsHb1
iWvR5EX5v7GEK8+A/FAXoZa38Cz+XKyLOZBAFTNSbb/6xGNlhHljQw8JjkMQ07zFdCq33YzS298o
SVClFaWhv877c32EoT2KDPaZ74BjmXi8YMYxrHcn4F8karMw4L6MTCediHiYST5i7WiZr6OhuwGi
uOj5GsZUXvF0CtwjVgIE1WFHiAq+UqrcpMN8lYPgEW1jgV19TZnI9yANRWqBGx7/ik+F+5BGfesT
vKWqDiRVgw26nyyol8NPYmOvPbEnlDZ63Gxvo8ouYcO7d4j54b/2R0kL7grHaFVXddlzbAn3TGtx
D98jL4Tx1Q/+P+DLMfnjcnfWxPcyXzhiz+zZ8+pNrt0cGY4O2t9hn+V4W979gtWsWvZmBrOcWFPh
ciLjqvEkvcivK90tCxGlcQP58ET/jNZYn05ZfniPDk/ndfOYpQyvr6q4yc3+JjUbISk1T7dYcn0d
6gRxnLYv3PF9fQaS7nLyrIPfHMcnmDn8yXB3eSrLdwTJD42fx1hUKGWjz1KVJAuBwL5YdsrG9jRh
U9pF3sLaMdiu9VeXYFz3Z7el/oZ0O78sE53enF9wUUPBtdA4AYxrN2a1ZS2weWcszjyF6TGoQB1B
ToCLUzAVr9RUxHhKcGYsE8kKY//gOjhYtfEukj0W1h36mz1A5VwghoJaZrEEGWLneJ5Xcb7bPHgk
Qn/1RRlzbSHPX6MV1eNl+IFGr8sXfa2V9AE2o7R80hP/TSCDARD/g0qErLSxffoARDRXyzo+1gFU
ZKWP8TL5F2COBnjWaYZm4x+O6wAOcVM0472sKUFrDvXp3MzZKK2X2akEd3RvMJhfS7qghMgvxdVW
cCzq8my38TzohZOYpU0F4uK8PmNUuIisA4reC2DLGZS7HQmAgEGAfLbI0JtbE5gdXC4lCUYkf6L/
Wm1vw6caw+/VRaM4xqn8Fs642L4AnQZ495i+06b8k9npC+VK0XEx/7zAM1SPqR7VWW7CRlpDOYfa
0O42obJizpNmGt0aFEKWj9mz0MBIiObr27n4jUs+GiSrhRaVWfc05vzQLXmE0iVGF1I8G9xV/bY2
QES036CsqrUFRLdAcd5MTKF7ILgfwV3dXJnxfPEI1o/1t09jEKEoC1lOF718r4qogu61VEWOW7c2
Txdto6y2zxyKSIuNdZqhZiHsY1DL9MZIEeAWD0yaD8PxXxMG7U0/uu2QOfStc2YWztYGwch01zFR
vT5xYyKYhST5icX9dLJn0eDniBXpSPabP915aHFv0cmIU5h//ixAPJpbF45E6ZOknC7fZLgBd4Qo
2VJGT4jG51/uYdsuIHtC3qJP/yEg46qhCLy8VjwvqrmzrW/mIwAAirULgCUtJYhFa+loAgPSpJ8D
7eHVaJPNhgj7uBFZFOQ4ofGeLMDa+Qw0fVkJDdUI08Mgr5bS7Vzk7pajdjy4Roq7PaqQa2LrEiMN
KxNHtX5PbJ7XCZi/ie4NgvAKpSmhIQ1n+PC3uPEIbaP2izjIwbTCWbizM6/KWadqT1WqqpQ6OU0H
fstZCPLelTN1qWf1jwV6lUo3oDPCd8pgxQhvagaEqE17tX3vizjs0Uc1PyCQo1vfQogeZ0L1ufF1
isShnH4ZEdck7F4Hhx294N2mJ6fJ4zQqi7Gq/akirx6zHP6zLxP/aRKfcORnzpJLR5xPy6t1Gt5m
ySjZQ7TJGzukXGszO0CXTfR2PTRp9wdv/hD4kcAMN5djnnBWgsjvT3GGyC1aK4BM2z/faWufOFXg
GaoD/9JCTwkB1i7kx0AhABCpfhtvY8YFu9HeMdppGvPSt8bcB5gbeAqXr3qLA/UOxCryAk5L4czc
D9y5MTPuL5rVTR5TLqQdrNw2A1Q6MCNSc+4nmslqjXmkvqG181dzIn0vC//8L/E4dbAXKw1GED6j
eOyyZOeClQ9J+XoSxLBWF0863ED+GB+qux0VOjh+A15gVOTDBBI5Svwfx9YVofvidltlT72St2U1
okv9Rr963iLz8yS0zzQ59tRVThbzrJERWijswT4xhWibCHRAimQfdL5AqL5OJmlFX4cILwr1ibu4
gEKnwnpMWRqBmHP6StFuzdS/FrfNFX3UN2XkSqMwO9MRj431FMqfmbGUzCEsrE2hzbyc0jI7jaa3
gywWX87O5f+bWJ/Cets85foynWZGBzLUDpVD9DA/YMENHBaNt//F9klzHzetqYgAb5YgEnEd76eJ
Mo6aVTF7zVjAaW6f3mbfIBqQkYtyMFdRSJfNjmNnSHB0QUnXx1Hak0JRfvbIVPhCPZ7wYAOzzfx6
bo6j0T4Brcu9blNFNucaN9SfAhGKAiAcjC/Bjex/FfLe+51roka2QMbbIHxpP/eKP2eCXhl6ZPu9
csTPWQV+47E7pz8RlHXNplnlzVHyy3zGM0jR1oj+o38qxLP/5P7w6JHKIt83aMpVcdVVJiJpYq6Y
I/yG/11g1SFQueIv2fDlux70RTYnrVoIjKsVhgvzO5LXD8pULLBS72mQGvIOy8YGrIIRIcLsJvNu
9Qyd8tupqWyhLX7QSTbmBpl1bTlkH2repTQzE034Y8rqb5/rWW4iPpvsdit4V9nw0qzMZOp1etPP
1oCL4YCPmODMVmWqEcwcJMIYqZvYC/uM51OcZypauOoUHT84c12VWSbjnfhWcq6cc2i7FxHPS0DG
K+kI9x1YrUFpatms/sxZk08JC14UNwKL3fcaKwSysbcM5lZ7LD3MAnM4kRRmIkz/IbdqpWMETFkG
GUSRGsnsnlRvU/YCLGrft4Rp321VdqQl5FJnOAyR7AqATRqdA3io+l4T8AcJ3vkEO3vm01twq7+o
zUtOGRJNSp7oleQYTXu2TWPr6lO6u1VJG6LLv1rN3uOqRVUF4KzBhAdwh2je3iDTRLzsBZTIEqXE
NpDfa+ebdnOtqKqSa+4k7zukJgcZvJUYptB1AogTaMzH3MmWMVKndLW57gfDJBXcYvIN7RPTeXUz
2v61laW1BQoYC75Y0/P4G8SZUlenST4hxc7BNsnfzM5em45uxw/bPT6ZzTjr0UYxt47MVxcAC71F
ck/yDZnkW9d3fCI8PqpwvRyk0mYXNfz8irZGH/W7kw4Ra7VzaOYG31koTMgyWb3J20V9qoRa2rsN
Ed80DvdfusE/vMDitkyYU7WmBDAvwzzjx9cxOR4ky6352oxk1TpVHTQYXv0qPQNz3hg/96wXED5a
C7GmCuEu2oWGC+afh5WuucMrFmvaJXRftK3L+ufcSqwR5xvvJQkwD5TRq3ZOjPRPL5WyQV4Nqi9R
d2tFO74M1zTjxG7VjAlx7o3cYPutS+92VmQBE4VJkYTTkez/FoFyyWXFQNLbN47kqQl4Cu+WYAz6
AgTp9IbF/uFVZ/lKuzvdLYK3XuIng6g8QMwN27fjtwgOFDI1Sul6CGGdWjFe+JyDERLpXoeP37Rt
tjNfaAnHXAUhJWViKL6cR4i6WfR3q2R2BT/0ZW++2b4RN9Y4j8Ew11KWT4IROmrxrjNCywu6jU7y
MdMvSlKwIdBUrR3x73zcdUug4JXb7YBV0bJw3HN8dH8hISPIvMlsAwPOdlH0RYVcM5X+UL1AnZa+
2qaKFw9c64uvNUKZuKLo2+CE3mP7FJIIpMnJudyxnzNhkSfXAjdcfvOdUEZbz+Ik0gpYDoazF7ZZ
MRWGqlDzM2EF2euXjL+q8zqn5DLrWMfXbZ49k+QrGDoPgzk3C8Nr9ykEdtesZbKpKomHRPcYzpmH
21QNm1Yeu0zVkZK+a0o/W/Duh/bNk0+it1cfX8gdCRoIWUkD7PSZkM/MgBU/k/3Fi6AgBUa6rpOV
XMFMjDPedr9/VVoUDYie8WEvJo13QKy2/dil91EJpR22nnO+36AfCa4D1GqTUP69pMQhL2vvISCX
a28qlNm0xTQw8+UL8Pvk8y8z7nS3kdf3XwWpKjdU+IQPFGutDjURy6oxEEYyTEjySzylwg74gMnD
MZ4iDgip1NlOAyFjFsLOq/ePeGkKsr+bb/0DhZLeNpLpSTlQxtxdrYbbJtgxCUyUvDSN/1F1iFdy
tq48HqOVEL4ff9JE3LTOrl0NBScKi94SWliiZT9M9i2WM/iCDt+yfGUS2zJQy14fPjPtMKd0k2+n
1Cc0a7guHFo5/rJGKbIRvCTPONuW6kdarw+w3ST30/K0+5J1I1GfZBS9KlDlP674SWuPH4MweH50
eIQNJgWyzdiBGgnA58TzjjeXlSaHa3AaGwQAYNOMlSyqbrTwHCTMAQgsMuBMGtiOf29QLGylJrMa
6TXKiQEEc0Tn8NkG0hP6eqZfREnmAb/KAs1kCmyWACenJ62s5vR9FqP6YsGUp0AGOF1h235mhEv6
bUd5gHZVwZRZscvmYUQDDZcuCSeDt8lk2SI4XyKinzNQsQNRQvLODEYrjbfFjd1i6fglm4ouKeOR
WZ/Un24dHepo4WWQBufwVPtw0HSGPCEbgb5MLsKJORPllvhz20RkGlrlOFFqasjHqctjwF5y0aQQ
30M4aTtDDhFL0XzL8HXZ2LsX03DYOoxmWWadJYOTnO/9CUlhxJVhBjzAIzi6tQxT9W2isoFW1EhE
J5m4ovNSADkNAOcOUY9ONm0YZftPW9NkvYjSMkHblstWL0o/cvz7aSMRUu88BqhjikGjxzLU0RuS
zWINSTSYczr8cMGfEJIoPhRp1Bbwuuxlnf1Xd+gS7G+UD/GfjZc875fJs2NbhjkMRQux1xUTNmGP
hZfcExo3akF/tUD8JWzrj01wZEVW6JoHJCoK8ge0cFFmFZFKKy2gjGVjerSYsqK/vH2rICWDcTFM
TdytQpAufX9FdaYy8bDKbYt/UUl0WsjH+b2j/Sb7e/lPei0sDZdZeV0sHCM0v52KJUV6gBSKgmnN
Wf4e7c0rOgbcXsKTExPcAsYKJc7+84oJ7cMLq7b7NBtWwrn2TKIS+aIeIgQum08BmRf4CZ9tYlAv
O3F+wHZiTk7mC9pXQWNpIS9g09mHnZwSWRtgCHWZZpIxlv/Uco9abMpS69DVcdLHU9bK1n1dlVxp
BwQ+CZtI+ANegWHfIJTiEHisGq4oCO4L1ytmKoPMuV4lfvSYZsQQaUWy2BoactoJbz4DnJ5eonD1
85Yr8xGLeMco1GIEY/uE3gfgrZmMLDOauEHTUE5/ZTlQ/o+bxM8SY/7mo/FyWjjN95iMQXWTW62C
My/G3q3fBTXnT7wEYanVTIHWk6hbx4cCHDBsloSBxxZR0XsWc8r5IJPnOlQJMonxQJBxfhAKvWja
6fTDJuS+ItHe7yU0XK2sLT8qLVjaxV1stbMdQdhH37tyeREPAxD48OWPIgm1OUlxiGBrdcXaHjmK
i1BfM4L60KRHMKZQRDn0N9RlcJwiHRggNUUqdRMQGtVnaSQz2tQm1rMLXvhPA1bNEdcj5kGNoCNI
vrrDXOiJRq1YO1QuM8Xo3XhC/BeLR2j7Wlm1xcOVpPpAVjUo3yMDWDVtHnTrjfgGzjRR+x7QdleR
Dog+Jc50YfZ3ZTug2ne0Rq+pyNhCl6cw8qOgUyHSzQnu9f37WmZC7qzlWI0dtDt526YKq8O17JCA
0DPHgOCEeOcST/Q/se2ph93eDTPBHn5E+KOwuuRREQuRH+38zgFt49zeYqom7PTzQJIKhBhvQCi8
MUKTSoRK0XR1rNAiYkbA5fVgyPw2ora/Z+DkRBZLBSuW5IQMyqbdeXNmZQMTQ/PtaQ9NKz3QGcpf
hGbkw+3RK7a5CkoGP9afuvmMKJwmR+nGdjxRFIaMwZGGv9bgJAJy/pwPhxTmOAKI9F+fywMvXlLp
njaulGh+xoVhHmWFcM6T1N0o7jgFqklc4mjdRjKv9CGSb7DnJWGX0UUe/teEe9u/q6vj4Siwxvej
PVioEFg2AOWCjvrsT2ugBgz/mvOfELNxKgOm7oyhjtcwaIbw7C/uGeb6Rhc5gIKGHUix+ZZuZTxS
7txlVGKYRzAL3+sYmZRGVFNcSi0Lvzx3SlIklc23PxlK5qT/bXIeAjgNcfLY9l4rB8dFP1f1p168
apZKB4m1J5+uXGNrZZR0snZcfnG1AYWkgwZOHz1mAtxU4DCzLowF2sZbPUwLf/LMj/5Z4+t/zFW7
oeRIKAWFPwcycYXIO1Tb7CXknHKFhFwTmhMvwUgBjyHtcs2qUjchrhsPcnkp5hoN3sW1+WZZzaXc
w2CORMKWFZnXp3VvBwtSwvuw7T1G7EcxU/0K5fM7jXOk1egBRMnKhchpUWkxgGHLNOf8cOV9BW4I
MPH8zejGPSv3x8V+GLnAZR9fQ7bSSPl03a21DbsemBAGP2uEI4CJqLDyPGyrRidaUivHZcN8rJlb
otMWR//0E9stBuMCUjwfBo9fCUtFvUT/lPveeV9XnCExr96Q4et+0RqtYD/fES3b/KZ+YC6JJ6mf
KxsAeoaXMWqJ5E7ZJaO6NtgzhhQe396xvthfVrCIyYJcbfGRn3IZ9KMG7WtoyPTFRMAlj+Xl9nzm
Hq6+RC5DtFN+umtdNK1HCV1Kv0NTx9g9j00hbHB9GPuiEXb+PPf8Ittqp1TZaWSp24YiHfKbk5Qv
5Zg8Ts9i7LPc1oGKCOAlWpL/JAQEibIcdA0Aw0A1ab2HTXT0ybnUNBL7cRkWc4G1xtM2WY9/S3He
VXLgY+7RzvAkcW8MA4blU5NtT9EmwdIgf4jy4S5X/TZTqIjhp5HJ81u9ovUEtYpKvQeVQMXzBJVY
wIDcA3pvv+h8XOTZI20ysZtThFcEzrIEKzmFC+UlYX5OFqvjxIY150cWMPTyLJ844pnebhqRLXYs
c2dTKMIo6hUaXC+TEshC21cKJsLKf688kRKDsNJoONnSYYUo4z0KFG3hL9HZtZHJpjZrT8mWL+Tu
5xmy6tX2NJaWhx2BB4Ag/rhR/4P7J/nVO/sytq3HQV8Rl2CcEzjbm5YHMKvELzK9vtm5ipBiE0NZ
6lH+JTutfSEXzGWdCCgTVhcar7D59zyvz8B0MAFt+7yz0kf1+xA/z8gU17xwva+xBhtEmE3YBh/p
ETdHZPSH5iNkkkrOQkSa3/OPltOnsCfW+OXwyp6lzy71kSnvgJfpdMZc4VVNZRnBhBuWaaQEnlK6
bpqgg/QGNW58Wog689TPnYDYdpbB94im/0ZbvjFO20NXHNYhyrorbd0ZG6mUrXwPI6pHIwoVHpsM
iu/fVOWYUycAb1Z3NcoiibyjslHhE8dw6oj94vOXd9/woaCuhUmskCY5O1jiWs+A+Z46ycYODdEC
mkKrCLoTKZaJ/JApW6S7UcqNg7cnzH62TDoogtVnb/K0U0AdHIhnC+zbL/p3s3Yf+kBUuFdWNf4h
z4+oGKoE1Dj802NSXI/3HkrcJNCfsCLUjtE1zTU8NKp0FC7hBUmcZxn38CKuK0hBCxQ3iNuq+Ckg
bYcLGE/3GuFPSGUwjJBX+FScNnLfoyojLStbveOqPnuYpl5msIQek57s2lzlMtLyxXUIdKT6mh6l
54hcksuWU2ieRtmfx0o2ceWCMf53jBHGSBn8fhVzWm1+/CPOxDFiJFYyzgAmmkHiJz9RfgO0FbVG
i/WaYkDNVEv8MIH2xs41qXjfdT09zaMqDXeGTqNHMOYpbppVPARTc4Ft1Furygpb1hM2FnnFrIg5
qQA72lYf8wF/XDXFNSQCtQWaYr0C135808GZLufPVkwPwZ1JeezrEsKBD6J+UaOnhEx57k/rhqza
7PunBK6cP9uWKPDLt0395cjw6vsNhB3TKwb0O/VUtvq7d0NMF0+S/3DjJ/XwMVKKVbwmOaJ/jF2/
jvwFoYHLOxpzUag1BdW4di9Agc9su7N0DZtyMzxl40C8Bx3T8ki89AI7E1grmtNbKMWZS8UbN1AD
BdejSzGNH7qRVg3EJDPUqVY5sk8ysNfjBS07EH0hC1Lzi2S6k1g4QkM+3dEx6dlAfQ2Db1sZtc2P
YvEf+gdzV8ctqY/z4fI1LZbo7xbjqT5OPbo/yumsIAQl3PcaoZjPqvTx87ns9m/PnKhNAp3IBrxR
Nmj6QsYvX3dqKleY7lNB4wOrMrQYRw2riyJmSyjpsuierFVBp49jCpAqIBbOxIfX5kqgDWeMWn7y
2/vUg4GOTXOIRob6EI+ojmkrtLik7cwdJFIe9YBOfmJxdbxuOCPwB5if7b6xPU7ULEargt08Wut6
URfXCIoTWhFasMwpIOyifhjnElNCwW6cVwp1K+lKQVT+dSXpiklTffuRR/TPyQQ/6Dp5OMRPdkvP
Cx3QtA0XL9SNGIdv2GTAFPFZ3jx8wXknHG0NFSMqjLtf7YHyIDJjMZptBgqTduFIoNg0V+Y/aOJE
uAU+UrhaI8f4b7DZhU6Xtd6HfV05MqysQeuSL7l8nhqryLZv/EK8shBXISZ+hWhdKhFZSXvMNdS0
ABgaSONSOAma7qGMP/kZzdLIsOblMBKJUYxqbzizfjPwhI07eTunBWH9jOgWHj9NbDRU0jmow8P1
y84W+xvf/0E1jbDot1onmUVNn5np2mSY5tvYwHoTT5faVTMEQqonU2AHKMp3nYh21bTzZv7e2O8+
UN59s1NmrHf9HnsU+Ye3IvgInR1wtU0DMNVoAbYSKlPGravMtgoPORbCcRaDI+MHV7quLDyGdnY7
6oq+mv0eONKq4zUOn2VlgEqDqzeHltkOOSk6UTT3VMIaRsSNjVQpr4jeeaRaRzk/RNrQyXmqZQXR
2nhG/lBkRN/+UNZ7r1tXCwXO7x3Fbm4jdttbcUuKrpy6nz5+ogKALv1H8IdHJ+jcFkW3K60cZBCb
Fy1aVbxz2D0Lh5/MrMXhNaEDKFCWEgAdzXG64ETIi3b6OAQuS24DFCXb4KgrlntoJIfAYndv8ltK
APAbXBZr+GMNqSHAXWKevcWOw8IKvCxltkTSz+bLT1t/+jNUMlDllnHnmnNYi9KbGIkSsLZXDi8s
NYJzB9hJ1shDuTNhyBRRpc1CsPfZlLuLk6DvLX+ZmgOp9azey2DTt9NIPSxPbq9rqjpv+8l2+wsS
YuSH/0tljd4D7ZjzVdXp45uvxKpoD8+hI9M3zjyvX0twE+dQeTG54UHdzpVB9LNSuvp0ZtkWJJcG
eJqecsLeBAqnw8d28cYnC5wYrFp0koRCUPeVWxXk4TyyxOCOSLKHdnmus5BG4dHeyx1wgIfu8oVc
Ac2jz3vjNF0qNAyrT+QYSPx1K+rUKRUIHBGDte75WpkJTfblOJt7PwPxKDR4CelfknngfceIRLC/
ldWQZWF2fhhK6abO+OEPLtcYfMZcQMli1rlzAhYoyij8hg7X0WJ5FFdaCtiKJswwsejr9wZaUQQQ
mm3qcuazVbjdXBddFFswE/GyzXEsquUDhT4UARpU01d4q+83xhDC+drN+7z2dnlNbUbkoupTiCuN
y/2unUZuw5qur6TB7qZXo/ugBN19XtSvW+k/gWpyAOKG0KuCwfSz5PpEbi2JHZlKIjURsZOk7bqd
Xoz/O2+tN+DvjQiIoFoiF0m4jepE/Z/Wc4L07DNj/DhTORqoKbcxaYw1uuKKcbOEofZFNJF7/H63
0jnuLvxO3Jrnt1VCJw8l5fX2wKigusXOUWkytjgNPwGqFtBr6tB5MqUGojr5zd2yd9QaEv1cXCFH
KGyh7fP28iT2DEXs0v/mVyw/C5nqaaGlkfIRwISiQpgmsFu1LEW/AnhULbIzaxFxamtVVKHUl3cq
7U1EEwidrTh1Athd/se5blWr3Vle754hIqi0gQeLd9gP3Po/LzXPGYibMjLLquJhAGhNzCJUTH6n
4zcOszpE/6TTq1htqfJNudeYrpLZ07ROHUtCtUXeQ6RxmsRHf5XQ0Fh0sgLAfMHPt5rZMS6OjX5g
wCqE5S2RU0D4juhUoW9NpyGovIZ8YZjep47dz6LfFhwEPBn+ECs3J93WzPbJryr4D3w2zOF7/FM8
H1yJfMPJL1KVfnQrpotI6vlLWeuYZ+8/RFnTX4OPG4koQMhvtga8z1l5W4ww3cRm94x98G1GMY7Q
5wzQt9SXoB/GUCXKt2+3Vk9rc4nP+yDKLtVf/WfWZb6bLOMbkDvp9wQl6FiTaORsmFjdlh1GwuNS
3iPbiyRa7G1188YK90cOhHSRS3lLTL9BJ0Fbh1hA6OeGpTudqZ+PPdTOIWw8ky/h220j61/JjHpF
+alFPgokJA7uyNr1kHr7q9GzyiWO71pinZrNmDeA+wX8ZY8YVJxpCUbtcIVOKZFu+jmoBsFGGSjt
pNiZjXtCEAMUiBsuiYvItwkScbbeg/NidedFB+vlKTjzkwj0l0JEyIDcEQTh2sjuHPlAAMPSxsnV
qH+6s2/AuCS7Pi/b6/drB6Nbr//Nlh+tfCd+voaTkslcpXgtktLPCeTw+kTYNAsPgh+5LxDRlOJp
+Ejt1a4B9Gn1+wfDsahez68TQQHryrbHrEW1KByQv8F02NIcOazpVAkZBLJf9uO0d/RFjjtaDV05
XF+Ja6baA5CI9O22M0+3WSmli1sAlMmdbj2puf8qUrQwU2gbBWMt1Y6GVTYWhaOs0JDS33fYEkg6
usFFdJr85t6cxRlwMWPNIrdx1L8EYaFp5DZ3OpeVWfhdydGD8JjWP6k25vRD13K83Ga1MpuLi+Oa
uDo4aK9ERuVTP14snESWQhzkA3v4oyw802/aVXhZpUlwMnvOidsiVlFGR6n1CX5ZEx2mCE+Q2a0Q
ZAH7arfwVE0RzkiFocNmEusak0vxfGmwOMajtDjSTJdFKldtihhT8M1UhyoxBlEVL/1rnXWNpORl
scQV2JbMQ6OezLOEL9OO0L5WWxQmbeYhTY0cAdIrAR9xMKhK43FEba6mrdnLOW7chJ6IE8iQc5S3
by1zqFWYN7St5gcaXWGCKQQJ6Q8JgF8WaEvwOTsUqem7RCOrcBED1iBWCrXaCrP5mM0c6U3LKzPV
j4OqLNcqSgSErfcchPZkusUM+3Myo96S2uVhaPEJnAvPxLl6wVN889subZ8jjU2CUKQ6Tqfx6h/j
c3vuAU+wwS4oKtxpwsmWneuyrE9ta6dBMn9lRDK1uqhCFApDhuqqcPyfqCehwk+/v375ULRiMXgo
FkAqIGNSnhyha4WDoAk4m+RQyV4y+qmwNE/VIe+g9cZbTfmHwVLxEARZz/+Y3+2JTPlNr104ZUOp
nxlC+avPpQbdW8zn5HNphnMMGmU8TlEOZf1tynV3DwljyH0eKBAr9ANmGRyWE229gqbO3fPSIdhw
xmX/RItnQUzke4abzTyCCCpldnjY0IfWs92PN2kqUEieXJEIdLrloH4vDhzjjU2b9hfux5J0JbWr
QEDRF9vDYc6Exzc6KKAd604jkPo2XQaGfhJ2okme2AgLs29GUXR9jBvdW2H4L662vz9O6fhc6su7
kH5RqNMdQ7ZtAObetSvJ87YhqZlR98HJyRJfx3X50Roc9cQvg4cIFE7nHbxe57RU7YX2sWNWN4Rc
KccB9QII7yTqbYDukQ+00jFdntHE4+w1Vu7oL7cZf/AiNtO4xQYCsDudjXSjmdWZ1wpCImKIdv5Y
+IgXnBLFC41s9OEDJHUqzY69Y+2+WzSSI+wRAYM+6KimRPBhBnwTsMdbbioIg5bhPVpdAHKq3auw
UeGBgiZR/CcjsIGkBnOKtmiupzhTTvT/HqIO9EUGWyDGp/mx5/yeSr2JfMYQCxJQnQhGt/N+kPbY
TQTvNBZdDwqtDMv6rDiec7qJj13izeSwA4X31Niqi5XH5p8cO11a1AFaV4oxi3sdgHAiySrQ4uEc
UYiUQVXYTY5QcKSLmWGx/dohXQ+89IKVtVeISofLW5keW05iWFC3i5UGkVLv0GTLHDeRBGH6WyJf
7jU6EkwHxPpWsjZrsFZh8XcIWG27hj/1ZIrLP3J0gfaJeX2jLfvr3eGVBjD09vq5mJBIPitMOpMI
b02sHHJ4KgWcG4Lx/At639wPt63U4S+hZsiAmt9N3ARwBZgaMPHCorEMmf/WSUzPLqAATqS4G0hD
KXQnkwyzJgTJT6xfA4Eq0rw+gMHfGHGg+0tJ2fS+R98nkD3nZ5jFXwvoI9Q6npad4hyNPn8/bh6X
PGQwJM3xiFZUA3YWXRhp4+ySc2mohhjEIYtBs8PwdJ2+qJt203L4WTZXQPz3ZvqJ01HdAkr0TYbc
j2q2CUPbe7we5PGleByQ/C4KeduBUpA0s2ra89MMtkicemsChjMcnvNBdlxXMzHjfLCbjoZLJqXv
S7/62zyrfcyWfje4pvfzuZfz50VmygIMyw0Akbbc70H7/viGj0caYPgnuGpyNp+5uwt9ZWiTK/X0
rA9eIrtQkOoEhGLQaEe+sEq3ORSGUgIv5ttYGG6SXxPfalhhCgkI13L3QE5Uy+8efI7/jlUgDyyq
4eYRMOw7rNMuFcsYkXB6vMYRPXOEHnFVAlR8H+lBzGx01288AVMCxq/XWWGxYUW/ci9dV07UILlW
lBKM9lVTxQju4WbvucWTg0wjq6uMuqkWeaVGzZfpSPKihlZDI4xgB9gqimMbX+D5kBfhlej7yAAM
gXGlPq+6pCQ/JJynp0Clrwhmvx8WGcm7nnQUR/jfte1rZLRM/ULuysx02JpwIZQTjdrNaDhelpVC
xwvIClAJZqt5RIQ9n5xjRfhOdEDdWiHaFeiXM6+Y697yC0HY9xXdoqsVmSLMrSuo6r0lke7cDd3z
HwSrLByMSR/YeylcXr7ovUbG5U2TRCWdauL16kUGF2Ek7OHKmNvhZSnQVAL10+VCWK7PFm3vIvn2
28A9ZyWRxy3jhLmB00RDxXlpAE6Qhofk9lMjoJyibvaj7dvjLNWsUXYIZc+h3QSk2JkGnqbCg5uT
dnfOSmpwhkt+BNCRPfzClG2WOtis9s1nbu2iGdm+IGAKHezuPw4+dZvRnyPkiKvF
`pragma protect end_protected
