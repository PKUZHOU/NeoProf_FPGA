// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
FXN5BFxxg8piAx2nS79mPX8OlPE7ImBFMQgDwr1CD7BJetueY6v2lFRjt3iZD5km
3RTvIlZZxYncfMyVYcplamGs2zXoD/A8xcwIjB6PIL8veT7yaGZVMOq7GqFEvGwE
L4OwX8LCe14TwUGiwoA6Ez5zdNLvfxiGsEewjYLDuwE=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 8496 )
`pragma protect data_block
q3Hmrri5Lgf/n4WqbqFVsyOUuKqP7Nzca1GJ8Sm0AwO83fpOdeyIQ3GKsgusUzS1
/f14l0yzjKB7M37e7ltI0cWnGvz2LYbZ8eG6+ml+IAt9/EIb0y+Fh1fX8ohcBx6i
MxgJtuSap71TIO635zQvp2TgRbhmWJcxF2KahXOssfRgKFhbpXxLA/kSjifT52rf
bR3ehlK2XqsEk6dEIyYUXNpv1F76W5Gw9d3pQeSFhaHVOnKcOsdV2xROpaRt4Tt5
dHnnXN1cvFARccj/upjID99kBAYuWSeEC9em0Dp6NlXSAyf3NS6pzBXo7OS2fg7S
rP8mBvQPipY7W7BhOan2ziQb0fW2PZHv0FR0X5yGpDd5FjFvwc6gVeawxn36u4mI
/cbDZKD2sgLXaPHO/MzH6+Sb/VBRvexYM1T91EXHWFsuf+4fna/vSUtzZD2mwuCc
B5KeA4JlciL1b+h4dGaghGjZ8uBld/E2yH+orHIfiug66+tGHLx5PdYB0fHz/AAW
CSNyxHx6spoFmuKhFYgBo8DYOM0S1s5gCLVbRe658n4nCbP7tE6NBU0BNOld9nHL
AF3/daDj6btoe22/AF/UkuWMrdpMh1Hw7aEd3ZU98ePgRC3LLb1nrQABcf4RB1m9
7Xly2IY4hes4bdnN79Vp24KtDN5Vz+FXwxCDknhwYO1ezEkJNMN59feK3X7Q7tRI
btQzGQKaT2sSFxQDPQGihiVQExI/ZLhPS3vnU71I3tvOrw7nCaTureWYxDXr6qlJ
uJO6YjARQ57ugvEaoqe33xHARykz9UathVR9CHP1J6MydNUgWh0h9CW7UKTjjSbo
35i9/fNtD/DTTCkM2S8b25wlGfqelycoIxQAdew9kdG+/Zo9TBU/kD/65U+gTxvP
b5ZZeG5O4ZE1rVBe9pak81nwu0sMieXyRjksFLUDmv3oELLpzHbDoPMfiOQaa8/V
6DX6JOG54Hg1B60C5yd/XaYVUZjsSzNujXM2YHRthp1nuA2Nnyj0pL4wNKmZaOza
CLZMGxdBPNnGdkDtS0+V+DGjKb62jxWLLdf2FlJj1b/kj3vNOKKXN2MbH/X6CIEa
A2jV0tmZ/EG6ZEHMa7azvFSkdWkRZiHpG3/6IoUhP7iTdJ7ofDXkEUO0f6QTHbWV
5WSv1tNiQLm5dH9fhweJLAGF5S6NPEDPE8laqaKmFeupn+vkjXg5iEdAqQFDNMi4
zGKP/eDcE+gH7SwzBspr34+3owOG98sQwGIVfZFBMvQPIDpR+smLyTkweq1gtlIZ
o2zYcEo7nSOaRwzRg8ZQX4VOR0qu+LwQueqB40mzLqNqxh2LvUCO4u5k1c9v91Rd
4V5E8MplYRESUTgroIcqvD3aM1RYLTgBLkGScoosr+41AAPzPsWt8kbC8guaeW0G
UZmbeCMDhk+QXuLwCL/crjFKQjizvx5fubKd66NjDiIWGcKCGpbZiDUJ5hefMY+3
epKKT9H4pzVq1XZUV8HUjp+zM6a6AyIKyouqc1jdADp8ueqeCMJVuZ82INnOllG9
47qglNiaTU/SsiybiF8ZktJm5/OMN2xcoNAwq3IuWHYz29m38xbVSq+dnqryyL1F
JkrsmMt9DMPiP33N16O13xmmi8lL9stB5lAmHE8N1OZHjMJ9jHIuW8QUWN1Cx+6B
r5PKmXL4MJTte5yCx9qXCciQMN0eA4u6eYcO3hnsDHe/cuB9KmiVIPNNM1YtVj2E
nqX8aNT9CjTAaHOVrvpBtS3jVBl5s9xQRWPWMdaVtIpzkxuJ1GmB5AfljnEYxvHR
Lxq3EkRQXt3S9PAli05xITPhr/4f27+OyqrRKMPo16a8AHQPMx8Iosu02xNy4lPk
dH8jMDenSVrx75Ad03mMcEhqV7kg8XaoitwpYM34Cn0iHzEEjxw8dpSJ3GxqiL1w
77+xV2xB4X5ozYiRX9D8NebxmmwIVeFcAT+somOLJM3sb8qwbMAKOs7Fa2JBZjJw
71lR0zLeMTjL/Fy1haGuk1WWqULJsZ0oNTF01zFm/CKQt4Gvm1ZWjmIflUsJ47rK
ZFYPuyTTxLOboNxNCxjg0P2tSFkwEkKtoCoseg28ckrbPI2tcjVteapulgm3Bt7E
9gt3CIEAZe/m+OGu7pCYg6gp4bocImTV2queDGiiAJUjVu1U6nAQ/PZZ/RvPnooB
rG7ajJpFjnLRUzOPsNWH1uvBO17+fFLIuS0WR1Ct0Q9OkpnHC9CIeh/kcvCnvIFz
8/ykhVWrUSHUyEefpjpkvuAqcBADg5O+6bx9n9q4gDXxcvbIzjcg6ftAM+YElqOI
ypprNxCV9cunqTYsXuTNWzoT/B0ElZREZdcjAAFC6lk3ZoxGEPBW/gjyWt36sTXQ
YEUXsI2xcLKM17ZZa4xCpx+zd0x/cVPR4HtSEB7072seHYymHmsWZkMjXYrxRKLQ
YOY2EOo2TUsbuJcVJQzXSjmJxcYJ3keYudakGkj26mck56zHPTWznZSEE+XeFk7G
4BQa3Y2uJEFPqlQhgBIDtSW1vFPZjFTXe1B9nPvmPn/uxeItUF9hYKHFp6ZTjs0M
hu5Cra/Y8dE2oV+ORHhdMxdFeNY++jbCqpKXu8XnBB96dWna8KzhtRJJQF2Rm+1Q
1cP1HVHbO75IK4W5TOlUrUCwdW3Dsy1/VuEoBzYX2/fC1nlpAABVz8DH8XfxwT2s
7G7QxKpLJWzARQqoRe/tnWh9c4mpEvaTesT3Q+peFIGfMOSBnP1ZxBdWXf60C4+5
KK/vMlq5ik2qtnN0dA0Hc4N4YVj4K7TqgkthmAXKfGU9dnQQPYAo19mDc9ma+ocw
iBHteaxxTd2k55WBUXnu1ETLiH5Av6ewimiBE7keGviSYVFAO5MYhsuIrjny82gA
givdCn3VEFtVcr0DwjO5HpbpIeKH1BCxvIerGuqBAggm+DObcpJLO/xotD540+4U
tpKtyZFuAG6diI26983U/RWyOD+Y7nl30WXJQ4ytNaOI1T3IN8gfqMso2wuTohsO
8VgohB9NhT/Wxsu8GlnOo29b1ggC5L5+DhCthRKfm6EfVfYNouQrnKPurcDggBdI
iZuphCXRuYDeg1+Yrl7MRXRbQX8SDcsptZe6A1RcQsrHwTH9DXMmdpCWKHBdbMcr
ZNSOuAA3xBYFTxdX4HGj3uHTXH0gd2dAqE4tZJFUrcgM0ycDjOf/KUn1EdQBCJNt
Yqz2Xzfrmnc0v7dj+oAnpPnVUCtmFVOgothSI3lrHLierCY5b5PSBwa05UjVS66v
JQ2g0+JNjlJw/MMp10hYr4iKKX2nTR250VHZNJqcevIHk4uOsTKh6uucAFMissd3
A9PDmUC43qlnYe42Hcp0huoPMkEiaRIXxvId3GJlfeXn1bzs0LP1kh4XukeiurHe
OYey3aJXBCh8SSbOKp+cQdtKa5F5lkZ2jkVDV8SVpsGdjKyeFnn7gOakXKtUA+y1
UiWcURJQi0i7p5uPdDpaPJu+U5BGRYlghbq1bCxGk3uy6yNKVwTF3Sj3psDUhd/9
V6LDnQTx5qs6bmTkaB11K3Ze0sVQlAcG7Rw+lw0yekOszhHpZx/zYzcCfl+WI/Ig
GCwKhr997Un5grgn1CQXYDKxC8a9pGfEp3wUIOV5KtZSWpKSNVBRNgvpP/20Djhn
ASGe5RnESBQx63QwPot7glncg5ThPbVI7MVds55ft1EdStl/iZWAE8+ULfpooI8C
vdcIQ+5/REtKo85rmNqDGpO9qYYF2w0SxxFm3oKaIZ2bU4tmCTLxUK3O0w07ixsG
ixFQ0HtaNAb4We0s2+pFbd+T4ZGylngaP/cXDIcoLRmqQOv4L8dkFEW3/aUlRA0G
xNC32q4SZW65vOndTgdvESlJseEqiacEpsoEfoThhn2IESI7E+wpQ5/Uhs7Y1lis
hAKxeCPNGQxEmAow3ug7Mgy96/x0GO8ZE37T9/hp0H4H/NdoDpfj0Co0dDbnLpTN
pOQaI8EZMLxF5fvswxPzfrDwrv0LE8qDa50/eQh55MvyQRnJPBkWUsXlwhK8Ku0G
Bt44Tr870u+teFAhcKVv9Bhxp8CeVkpflJC+8pljS8PpxocSFGt91+OqffXdiJyj
GBhj++IqIegEnAI45EryowbX2o+ZgJGmAGPskPye/eCGSxf/MTRhIbM/KXgilG9J
bQSKXSEhlH7Y48H85ohYUVfLZI9I58KSnpkBELOe4TosAsXTyf50YTZd07yMJHvV
zE2OI+wexjfdNeORc8xh6+97T2Nfl8lhatN8YPTxBHKf3najKOgjW/ya2pvHbq+1
Ud2tn/kQG6Gwu3I8csbYOO5qCQbGBy/oCHooD5OOWoR4uvvbC5+hasFKVtFxytQq
xGpKo4+dsWEfAuvnoI2QH99DTthsECBFIZ6bIRKGvkvFHez8av6g8V+BQf2i4l/Z
Ap8Dp+rx0BhPwJGujQNxkIWIcBGyWEPDK6ANbpz4gQupwL/RJcS+i9Z4Hqx1Qq0U
SAoTClWKziqLTsBZ6Qm6w549jSir/yvxJXHbBfc9hYjWU6QNTYYVOcSaL2WTQaY8
Yr7fmSxFNBL2DBtGnKyGIU6yoRGAkLf7NWytBphlEgsDu4UXF8ZxTrW4A3Yh5AOn
2p7bOKOm09VoiwgIA52WHWXtOB9ANMltOy/5B0evsDeHA7tw2YgBCFQjJ5FpmeWZ
hKyec13x962IxN3AkuWpr3ZhhHlXhpc1CNLLPUWYusQ+ZeV1bqpwBJ5yhp0MndSr
Ndmm1eMqwDOLlEy0OJXZc3pGOCvybpSjcfCDi+8C5D91HsS46bsTDcbeJjeA27Og
eunbxd8Hury8CloWSaAWTsS1SBbAzhpHnY4jiqf5imcX0gFnzPS1whTk7vQYXwMj
BmZ7oPofCPeU6PppAwYdIMH5BGiHVy6iuRqWN+ZznAzna8Zr8gPqJl8PWQ4K270I
oF+iwGTqYKn1os8//1pEHuIPrYXvHAby1Srkf6ieYtTT3sTB0XaMJehte60Y4vQ6
AwRqK6DMzkfeSXgXVGjQEMmKE8E6Up/uEBQCaI/5HrO5HsB+GZW5JXHcbFt3rwEG
ryZBHIrotHVPTbLfDeO7CSIWXEXWc/XDc9LtqDsc88IXlJBPZqG5CPYZ6I490zN3
kqcPNxHBS5oJCCQuTsEIst8XIKLdGc/6hf9WtNhZATq/oJUfRZ7vifNypcdxiqmo
lMfS97yt9+hU8NrUs/c+HV1b+4M7LH+lXyTKWtLJmw0Co1iK0++dgaq7LaO1K1Pr
2m/8bHPpNfpRmy3DMpluz6Eh5d97bEMwY1KO1M/j61MtRIYIpiysIx3hPhEgoGKg
FkqpnRfwTWbmZ01YHey7dBOA/ryVu5J4AOkSBWJsvMxEgSfmDhZ1R/aphnfTDOa6
/NO+DZCn3JEXsY/HXD5fFsdvi74irXfLOGrtPazcNN/G+m0VA1A/Y2OF7soeW22+
BuvSWIcXJspnKdGQuCD9IiMY8hYCESRyFgepdGLaKCXK4Z3L2MkYgt1/r+WyMVUZ
qTFYRgI1EMCbbRCYzwpT9qxk3UTwR1u/J33r8GoS13WOK2s0YUiLqRsyjF92XYGv
IXdJQnNoqC9sjLVy6duu5/VFUt3a0MGPwpPuAuawbUIDWy5SnZsyJ5p6+li3+2rU
0n9mFoOv7yLrQgPL5IgexgN+LVFpKgBAgYYPDaQwoDiTkPvo/hoLgfYJHzC41ciT
mxj/HW9mMtMaPGeRIUGY3/qS4e7ml9cIlM40PGjiGLrOS8zAEhyR+PTieBT8CwcU
PZfhaw3bEHftKmXsiDsLstTm+exLJz0nU3Fke6/DvPp3XfELFTfasrAuYWoaXbau
rQAek5fPd6zOdhbIz+GqIvKPp+afgyXzxjy9XN2pejCQoNBWKItCQelXDA1Alghd
OcDt8yBsHQbqjnEnUafC0wA/PoyAnmrHBMBqy0argfx+bFdc5vVDqU8R+gL9KzHF
DoCkK5Fq53gfDxhzo2OdPeX+gYFyM7KJ87gq2HgEEhagzf6/nEV3Ox7v45M/7TDI
0pW1s7tAoPaZtneKaC5jLgK2f8qnLu0orDN3UyOiGrtJBc0Ifa3vEh9gElU6Us4n
m9lyniUO8kQ9Gn0jHhnHXZwgp+YGSlCwybc75kEn74f6pIM+oq9gtHzWh60DoICt
kA+tKR5NQAuFp+67U5MCZ/HBGwpb5uZ6Hp/aZg78TPGtfTtj1pcSlVWg27sPZS6M
5d5+dsOgYFqZP229kW3/Pzdh7Sb1TP2L5dathtuFPBws0CwgdFgWSyTUbFAFNfOD
VbogEbtrMtfOB72JZXpE1Ze1JEfRy8D6OTdyn47SsmL6atebPoH2qBGPIwRXenyj
tZkDfMGFKUkNuEXq6rWz+QFBpcuVKVeeK98uy/V6n3tccRWZLq7pD5LnEyRlTJ0w
ij0XYv+pmhb133LZydd6EycutkMam15QOxpMBVXkw29S4xt6jWKEqdZDAbz6qTI3
nWtLlHfbg/A5rR52yKfPRNwD9gM3FqKaa0gJpXgr1VjP5tlHPs/A3WSahjUuhF5c
VzA7mqBxj/H5N5UhndyKUgdPC5mfh+ktGlWZE7QmLMWd7uiav1Wls2/O0ilwbVUW
BXfZKUyjUF73UtyfLC4tuSGsA6cJM8QFa5Tx1HkV2p8BGXbdCA47AdbZmnqNAdcF
VkMQkr1n0CWAZHl27E+Ii0d5tciSGdnq9bkf4wXhfzKSJ/pbdR39hJbFsY3lSeaD
e19IkDV1oesJ/fbIKlP7d1FtPqbs8dFb2Lcs2K1sceELtTFucjyJuyVtpBoj45kQ
soentChE8A8vsIMjNyKmkyTVSaMznbZL/nvqFegPMytK0VT/eJK9zj/nKkhUxk0E
a7Cs8D7Vj7gWdY3C3xueEBf3ahVKZAKNTKeKrDLm+KVgISQVg4h4ZU34E9cCxtns
Qxc0NhxG0NXlJ543Po40AnaIIkONNQlUMdGJYIcPYOcjpHbLAU1ltFSoPNDfG9ow
o86DwpClvlSgzJxGxGeIwAEW+zcDeZRH1jJ6a4KQ3ZWr69u4JxxqiNlIorgeTcsg
fQ30DV69wArcVjfNYryJ+cHFO8VrpSCxPEbznYl20A56HXod3YCmZ+AgkUryyQmC
VWRgqqbTNr74wCaI+2nnKNd1mol+IpfMmJzyhuDwcwhVu7BBKmDoIbn1yU7PHS7b
GAI9EC8KklEAcQGeswjn8VDEU1Nbng85h72pK65Sy7fihsmsPxc3ek1/MF7dRgGp
itfa9rbxvWFEQzVOpVuxNhMZJBgLFA+ulSDScGOElYlnrsC7IFfEpeBBqgwoTrWN
tZ0mzV24AxsY3BUwzMzjCxFQU/V2K/z8HMsbedl+2dLi0GriODb2jfvBWFxc+KkZ
wYDZ6mWBaGTqzJlcZNfTvo0WV6yXPy7OBNDwOqHlXguOcyohY/9g0F7mk78+F/fS
Mf8CPhIUl6dhIFdVAkEL0UmgkcqjOWNaF6lsjTmBarwU8SBGFk1axQJPe2yIhQ3U
yYuvxfpwPcBtbdpfJZn9xxcztuv+6IvB024jO8rBHHFtPQxwYf+1hZJrCMepR2Ls
z5Y9q1+Vger/CuERjW0K7o0eNkVvj982azcEL+qxY4fKzuJfH5XWf7X2UGj5xc3+
PsK5sFlj0+GD2D8uJVheVRQaFDpDLycbDeBEdg5qf8svitLdWq0pJRWiwdM8JwFD
xYq7SiNEh+voMXmPQdg+Yl340ytmAWbk4u6dvjdnzBP8gxSoCxAgSx6i0nXDbXy9
tLytQGuhsbCIY2UQGb5uraaIRfmnJKPFElZWfCO3xoit8X0DPaCzmW/028Z9tEi8
9mhZqyryNuG4WFlltj+0pbUTIjwWqf6qk8u1K/57KkBz3MxZIaaX/0iUa15Has+I
rLeQkOn/Ky1OjdZkHHF4beA8L2wG3Foa4c0G69JB7nPBW5V7ZncrTatRw/PMRQi0
m/tYNABAANj0fhjI0xaiMGi/7ZfSSkfiOWc8M0u0zzF7HmAJaCu3m4SHz2bINw7l
c1Ad6LyvlMmlNm24arIG83nkyE8lMmvg5cN2y86PGFfNz6piLFJec9o7bljGh9uz
fUH2LWp7uSO1Ut5kgn+dH4yJEuoeP6ELdWn0IaIYWUvX5s9qAZmiUTDe02PhXxXq
ZUmt8RDxULmh5r6bmYtznu4Qsu9gQBAiODebYPuwmjD2V+zpdjT0ewSMRqPzBnA5
btPAsPN6GiSuo+tGEw5PbX/L7GCFMXIX5GtIFVfMmnBG/tPfcMHSPyvumVQ20dts
4Yk0NqczM2JCrNeQFVBW9FIkzm0KnX5ZowgeFyxU7hJlWx2BT7iM099jFzaGWopz
liEDid8BuDP4xPeAzx74wlXdQUdc5wq4rkujmiFV6uQMOSG0SEOFq7skI/REu/82
JuYxayLKD4sQ3p3VLF8Dt/zG9uhrTk4in1i0Jm8dhMI+mYEhn7+XiB8EDySw3rPQ
otQHLRHA5SpkQ+WVQsJZInT2ocxb6pCUw2guZiV2C0rfoUVAbtxiCcw9TdfxmCKv
c+ZOY3Ct/m7Y+d1lPJJMyBrsPaCwqqifzppUcuzmtMmkBq8uHiBV8435RaMmRaJ5
IZfEQ3a/SnnMmmrvv9HNgAn7U9ogYLCNV77GNBL1P/oqmRK6UG2N9Hjv10Acg+7K
pmJLwkTTkTgXcEvl+pXI+Q303u0YRmnsJ7gnM40hEdHTewRAIYJtZl533FkRBi8F
nE86t4717N/X6GIEagsc9wucTGDWNANm8A8MUj5m6rB0i8fgjOisrtsU1mQI1xtf
if2R1oX/k657oga5WJV18V9lCE9kA1T0JfF9rc9ZKaDBJHZorgcjpEM9bjZ+VkuW
wEKDGwg4ZAxaS/HRe+4lC0l8NgIYTrczohqfv/c5wiY6BXWVXh9EpbJZYVpq0oOh
QEdAkvfTHpbQ7MILSa8asjz97gCrLnFSZZj9xYZ4+42/IbiKRaoAva7V2hdGvy+H
30gffwKs/M4QBciE68NuMWxiEsMMj+bAZCHtopnoHYc+LQ5gTTOkiX0SRF6ZLNrD
lOe1/p83B46X2YGclNaagn8UQ1rR4KqwjL9nS8WtzQ7x1HVkaqqL3n4KLkuXMfeU
XwBfMhmPwPW0BIuhA8xdwbzSM3ibrdey71OLkUwB82Fitl62tB1eiHnW2YhXu4k8
wkIOHCuW+MP6Ayo47Xg876Y8+uu3GG+/aMy2lRVhGbLSeRi1DXamTQgo+aIzvnsJ
KbLewp6ogXN8hmRl0l/oFIyIi+ILrrn/tN4QknVmdtWu9KI54Uk26eU9kOoXQXix
te4Rb1B+eUMEvQuqsjo2lQO77tPD/hNVNua3mytsjXUuPuu26F6sNcRJ4VOVDzx8
tokVlPQnPSDhUfWDPFIzXXg7bwJG/qnTJ1E5idb2TNEJm+WB56iE92vkCQIGZ6oe
uoq0Y3tdqjMxBBJ/yxBEVf3ubje8B9knEIRVoZgwj+IZa37UBo6/pCobFX1EDGmT
MNkcjHAKRmoqmkH/MMqKUXConxuiT6tqBYcdtntu73C/XzHXWsEAKpNHes40lLHE
yx60h42PwvzpfpuJ5rQijSBdmfA3hTWrERENfZ+qkZzlyxlUvOQt95YSV6CWrRxY
y3tcAV2AmvArQwnJWrzg2QnGqg+eg8tUcahNBIRHpVWbk+HeZXPaBb8IFuhbNVK8
8m8PzyE7+FhtNU5boe3f4skrqik7+lbKo4jncy7S69ZmHOJCVjHh3Jxh6QkoJX/+
oeBYjDUyqqxfNlRVSyL0+P8nIyavKyTVu305Iipftd/wVANDvhm3dfAmcgcyRVXS
nb7MK6GnzRrToHs67/RZNT81RPuu3hv81gFnY4PBIKQl8fp0wQh6dfggFW8GFOos
vG3vn5Zzx4ZpSsM4Y/3GUdfOm10V2sRP/4ycT+/xLMMxSDizTLk8Uxrw20EL+9Hj
/JkO2KfbosK6gxK/oNWOhzN/+dca6NBTPLZmqzC2BnYiBT3B2iLuIVENqXgz1e7k
fC6p7YJZicqjLrOS+7GpikssmTRWmIEQfJiuz7W4+cV/CKZh9RjZfqG1g1qR51w3
JhmD36ba9m5qvrVVs3hPXCgNyp4faHdF6YFHxE/gCdo8ew+W3epx6YFpqbj8pm6n
b+symgdbDkm3FJl30eTshXZppF4EZuzj46DGcZa3m4NMF8VJDSBeXgQ+lxNqoBvn
Sqrqisq2PmhiIOZxpr+9VdYGNY/uHPZIVdFuDrpa89yvmjpRRuwjPiuj94Ld8zB3
HE92/7nKolwdQcRGqGyVL524Lq1T12z1HP/6fJEaAoyK/cYHKAhQ852xYtmR65YJ
dslLILfZ0JhmxoI4UEMVDo1sQwaqB2F4jsTmXGBTgZHOcWFKiu3I5hB98L3kf6f1
0oy6RMTjNCRQyHi7d27oOhN7jW02klTg2Q5hKA5N0sRfNFbRmww9KiIlTkHhAJbe
t/s64yKvfSn4Y62HMbVl2J8Pg43xd+l0uoKofcBlizg4aCgCJ/Sy8f8weEKM2GY/
b9esOIi/EgFlvvXjqe/OjmoC66OvgXyy6pjlknA6BEqsdGy5qf/HMUKUayWyP1fV
718u7siy96oEfVEg2DO9IRtXN3cB2CIj+Q/7wzwYYyEhn7FyfMvqKG1Q1uuFrFp0
06H+mv6DJ3qtIEookwAvwD7w9UaTp1ptYuPutGtpmQwhCr1xsVeQyqlMUpWSmvWv
6lRqQxCgIjiaztmVUDD0ngBKoKXnLMdTgx/2iUkhSof0WQggOzVfRxw4owueGCg8
8msvV1mu/nN0oo7KW/OcuKGM4/MuCXedr783M2pcloKx7E9AQ/KFsyWsd3BNhAqN
15R5GJnzB5o5BtEimUbGE7maZlD9VxP8PMuxBFKWLsCDlagxVY34ob12Af4V7iJX
0qhuumkgsc9amGFfw75EnePa6sQNsM9yPdM9QF1mLVf/Kv+T02Jq6s0ZI2L3t+W6
WHE8lCW1H2rcEFuFwoqYcyvPkAQ0vuHeOt0Oh8wHHkO+LQTU3flbSL6n3UsMJozb
M5GAKYIoD6HwnJ14hGbKirbOp1ro1GVJJZu8XO3woGpivPZZ5ImWY8pkJbLYEw2o
ZjzAU6xw2GtmO//m1u0le02omwtusMOrI3wKxXyCKctZCtKnAIKO9A6KdMsW1rZ5
VU3V4zxuYqL5fRzMPMR8l5I+TRC6HgZ4TWxzd3jFi1BC+DEK8kecy8u/vhF+9N69
o77BtRxP0+1T/S5HckZ6K75jXZ4OJAeqs+TrGrC6FeXnGgz/7yWQk9BR8SP1hka8
I5SKALQIe4f0akpmE7e92zKU4POfbrCDXNDpHIsbcCT4gk5+BcWRZ+txrwImO/bQ

`pragma protect end_protected
