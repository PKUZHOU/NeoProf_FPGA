// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
Ci2idbs1b+wo+U/AHl3sB16O61ke+FEQ9ZMOF+TbVFM+/pHpz5Aib5voRfqa4eRI
8hvvYQSf14RF7GwzKpCjEvDFtM9gXPfUJIZOhFbAMImhcxVNI5er0iH4sEF9AWk9
HpTDGYCdvquXVvULKuhbA04vMFACY1smpkDGHtx2Aes=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 8640 )
`pragma protect data_block
WsnG4kZJ3AdQHi70WCER8+Lp7ol+TG1brvxSvRiB/dVxfd1mGv8uCJWtJgTIttbK
fCVL73026kDyuPTJgGE9mK0MWr/ivGFlw7BBs1bC92lPkj/s4XyWXTXk49n+Jvqc
rrMZ++XyzNxJCGNwyHazQ68OS9g9x79lpqVovDhzJHPM2LyMSXIasxg9nwBrZCmw
Z4cYGdvT+Lz2VZOfz3Jxg72Ed9LtlpC4mytSU4utShv7SiM38ZicskWYSIoOv7eZ
Rt1176ZNPToDLZGf49QIltqyytzEzIUKyUbgqtnA9XyVXxxO7qhbP2/9QxRbZbjV
uPof7HNs7MrpmZclltHvUbJO4hRFHGF4B0EldYe9dpD8fgYOb00PT6kJG7GOdS8c
BpHFOTBRfvVIk3MzaKNshTmCL3RfYJM/gUsn9IKOyTdUyaC0bDFanhbwdy9jDNoI
/kXLCiGEDHpKKF+qK/ivhlqO35xo2mYK8hnVVVgIKg/yIn1Ac2AtbtPLI4owNjvq
V7LJbodSsN2dj5qtpZPQqKduFslx9T2l55N6gSu5w/VJe16qilpHi2TSOCboFfLT
XOrn/e6EIryPVftD7N5UZXZIS4BK1o1o/doySTKdPWCpm/bxwQ4Jv5d4mmSUYPhP
/44t/dJ6fMoFL4fplZECX7z2Gs8JbXGbV9bQAdKQdbD5zoNhMZ3HJqKooZHOqB5A
9E0PxTlKpgiGEXOnH1/t9yftfTbr1Pf4r14X7aKBCQZJFhbjn7eU2t2HrZ+Nppqv
K6xyNHecQjksmpoc/jEGnKu5WNccC6+UnWS60csZiRuWXtzuKLEBbBftl44V1dx7
UIBUVERHAOET03yGco39qldQeJC6RKjpin9bUQ4eGrgRIMwzjxdWrYdeYQpJCsjm
YRi1WbfsYcBeY+/vB5ITyQl58P8QLFJpuIFmFv8qt/hqZMUbtJHzANRtQu9K1OU1
kE+fyc0PAa73MHAZtDCMcZy7NgURzaTCBxiYE1W93S2eHdJZbATUu3HBDWpd8IVX
t0keorSmzscHbM1IC0ruWAJq51qQkazgMPKF+WnhHm6E30aqIuG56wxh+vQEAqBr
YqRRqFoit8vy7012qp4ijXDjK3aiHV80SwGMscERKZHm7efQqvO+nJfesBaUh6ND
xIQ5bvm9n2A3ECp4GXm4vbbrKA2qQN6vezpurpZ5X/LT1NKkA9/+rn+MTxB8kLJJ
RtOx2Ff/yUuvbjVloJo+s4uQ9PeaO/ED3Dg+zsoHmck9a+x+MhusAl1HeKgrUI77
K46dW71NpsNZOL/SNa4xwSxEMUYGXU/rARNvlB2YLIVqjwOJdKTFKJX5qn1+gx5W
WZusPGQ2Rc6ExsJ4ZHHrOqBghHQYbDCtFzruG3TiL84LUNGLTeAQK+e52RRR+IxI
V20jXHXgecQrT8WUK8E2DTytgRlVxoffGLSsZXTiZn60vRyIeRBdvOYS96dAE4x8
vyWbjDIYbCLfH+ZJoe7qH2vJGzTlz5UNiPLBORCeFEMQVlWaAKtEmT9VNPTWywGv
aGXG4vkhwv1zxVbtDEcW1TOdS167w2miinYqy6m3UVcS/1hMqhPLlg2TDz02SRiA
QdtMyyyVc/cAtux1/AmfLNSXyG5+VWHkz3OwFbMKb3wQv06dHBcKLV3oGICSkQ4c
UqoiO8XGsXV/qTmKpuGR/wDNEMSm6EsyXeqNdLPHK0yL8svFbg9jl0QTIS4VojHc
u3ua4yKbuAQ+C5qjujMkn7osP3WOrvfWyG+N6YVMOdlobf4xt4CEvnDJbf2j0FFO
DtmEGU36f/QlfY1xJnb/6dgDKDGblVdPzVMH6fGwHrvKZP9GxpTOyZFqSkLajntY
g4a28XhjM0EVTz6KXtOawWfjL4UtpHPy6ASBpvGKeJ5qzmO72kroX6WiMVyXFeoq
ynY8MTaPUJvABfW7abdt5fmsZgWOWyxAyghVGM9yv1OyTvRltu8r3anJk2ndGdsh
hB/I60V4uEG8kO5KKdS4nQr0p8A9CghuZ+Ic4XR1+6u622US6G6GQlQgMwbpLHWb
uJodiwsl8+iT702n8DmA1WkP38vbTV+XrdufzpaZbPVqbO+KXUPpsMREuwH1KoLG
lUA7hDUtn8w0uktjQtaxDMzWyVgMwWYMVUNk6DV17tfkEA9Yfs8GVDq8EOTZzKwr
JckVWJX/qUbjCu0onr3dCTcqQ3G8Dbu66+iARoFLHwTOkyiic6+7VkWKQeD5LaNF
LuDt/8RqPdj/uQL9g4qfWlgR7nYT/M4y30K1ByL+AOxFmvh3riZl4r1aNPq9HPYP
WtssvDlh6DQuljI0L8ux35BPL53Ya2wmdBrJD16SyBBApoyAFlYlQ4Y6C/FIo3Bp
elYp6VUHF0xC5fPxKNCQuFtKjC81tu7P+0Gna6zbSpyHR6gGaEtSOBG8R8hpgTlw
ihBMQjAVQaD8tQxItu6y6Ck651CMDH1aDqWdZPV2d4eIFI1D82ePAnhHXNiwgwDw
rerw5w/K0dO/WKpWR4e5kWuRpbiZKf9sAXsuqTeBIpYl9wMXuAD8dhXf3+7rAySM
ORQDMFRhMxj03tX9huUj4hQ0jRj9+q+iiy67aqZr3y5nriCbx28GWFVlSM9Jcdy7
07osivrzKMGdnnl4bO9AJ7LKXgm878QsgkmSBDCES8n+caUhIcmyNrHM6eamm7cW
kqqG6XpdyH9Qrmy1QgSy6Ra9ohY/OVS1V6dJYUDYArVW7jn5nQgTSWA3/fmTsKpb
XY1Bi1P9Q/66EwjHyhPqln0XVhq70IwHKJwrJKMWnFNSeFON/V7Wcy/skCcCf3XA
vAMONp0eWcs9DnobxPIZxammhT5ugWswIC5KuH241BdLYRE8l3WOeUOC4XEMaQFQ
PiEfjyklhpmyODPZJUOrWSSkQQVU91yGE73Y83pJ0UZLlUZe+pjr8Lgj3LtjbHBp
5ANIwrXFL4IQ66Xgd38e4wslju1GgQYYskMGydTqeaKflUdYpvNm8qWJhkHX2rAS
7RM7TgPrVcn0MwSnP5yhzzasb+QG2y48PgmTbavR4JS4IGvQEP90bUsmHzGHb4AT
31S1JtdBUYAd0px3qjLWUDbXkPuC3PZBjTPp/zkBgRtnpUTeLFZMOuoW06Eb7dIJ
TEvHRgwvrf9FWJksTCDJ9ZHnqdSG8+nbr4zLeWUknoawTNVe6GIm3lcAFDsJDcX/
zSdAXYU1V+sRwaMQ3ZuMk1vowAIOBa1G5O2/r/QvVjRpUHDP+KjDiavt2QdlL/zl
ZFG16Rw32LSqsLg8+zViddtsMhNHtNxerAqWwOFRICoGLQXTs+3kKMyCe3Nlzj/K
5qETDIjXnnEGY1U+JDD4U0hjFo+yLJH0pM3dAxDhLrpMM/Gbr9/ogqSyavIBv29a
tbdE24zhOjA+u9VDURo3zcAuTLiHTRv8wCuKQ+NP2RV9IA7Az+S5qjU0CQGifML4
JKWiI6KXiOdyWOY+y2LPD1GV/QC1G5DMOlet9QDbKX2NsFigQFIa22AtMNWBw4V+
gG7uDKtzZlxhRaoOzJW+DP2Fi+oDqGy/2tUt6o6peZjxdyI2hC+UHIJqJHyZZuzR
TJe3HHGlCLfLcEvrNMLSf1IpTNPZulUwoDKO6U3GVIVhc5AQDcGrlhfQ7LhKg+Po
rQdghTdLzIr2TPYxROh5kMEeNRtBQK5qRCEj8sQzDb8HyFDvy9QEhWYhhd0sCDhz
0rwfJg22NeXN0QlgCFHxRqKBG9LMvmyCdrYsxbuOec96+1HuONyduCrcg2pszdqQ
jhYSOygp+V6bSj6lN/2Z/c2zWM3zEPSfXpNNmYio0AMtuoZFcSkd9S9UARo8wGok
DsMQlLPWR2h++RFgdyI/gIT6M3R5DaKs0b1vcx0vfUYVvXIR6Y8+JQx07uXb3uLB
AC205lfFjMES5ybXM6DFkOUuUMYdLwuZ8U9VGWGy3c2SdTp9UHgZY8Dl6jL8OqIY
pwBiwH/FBeCrQA4K0ZQmKph5oCKgjQ1v3Z0d3fcj/9Y2dbKRcuHnJkyGkyepG6Z3
kpBg5CRApUxPkY9gaKby2mr1TVG6dLSoP0/6StY+5DtfW0fLYnm/7SzOvWunnQB0
at7QLvZZRDjAIUd58WuZowt2Ek4lNcRW+QYDEjD3uak9McHnJSz550F7y8JQD+LS
cd5nuJGRNwjkHXcbn8s6iow5UPihmFhRYzHBZR3Ep/QOi4r7EcjMG9aaFSnclVCi
LDaTeYA5Mq4WsYlgZTkwVfy8+emcnb12Hqd/uJaCZMYLvdKqhEk5KlfJPWng2XH/
hrWHkd5bZUt68bYe+fxMczOeAfxyD6GFN/fvzjqaNMHQmhfkGiw11L3P8nNK74Eq
YPVuj0zH4OjWLPYsTEp3VX0kiPUlhki93YmR02w8J2/HcQMuqfqom9k1DJgH4gUE
dkaeN6gBwQqSlVxggsOlUwJ9H+E8rcNaI2THCSbt6ZabVnNKs3P4IRS1q+mQqNnx
Cf4gBWJeMXFQBdJjzX75rUU/O/swY5VPa1dP/6+pyNEawHnicj5nnSMbVYlLxJjI
Ot9/C9/6UBdX3jk+k2RdDZAcy36KIN66vGGUDq8+2hc5zo1pvPDxMhjFAHDyaaDT
7rxrKfV+OL3ohQtwiKOsyqS2hT3kehLww75f57qY105k3odanocutxcEiQy43MNa
p9YRHGJ5xOL4L602oEfEJdmy7JO4K10qq8YsPQWWdFR3tH58iDDy/Tq5Aj4p33k2
AAZ+UpzOrXjfibPvThoidmTd7RSvA0sHIEkHelFMwtwPBnkdKgjHPR1DqqQQP06j
9mHrFSiKlCr/bylwt3BBgUp7BycdRMdxF7AixlYfFeF5zgZCpvxwyAZA2v/oiSlf
Cv1LOn50S7aZci9UXmUczCnq5JtmZZ6v2VW3FOK+H4WiWr84hcspcCkGGinfEJnJ
U1d2OUj05w4HRg1tYYrwX4ryLlRWVCtKaZ1HL511ZpaMMT7JN8Rz7fBhmxTfXadr
rxBGhYr+AKRpdylMsGybSXUngOWcImJeofhc0FJVkDGGRuDlApI4zWFeRYARLhpA
93qi0hgYt22RdwLj+y1bfrKDclj7u3+IjuSO5H5O0Wx9XwbPd/5JQMy3xAcoRDHT
roWskiHk40w9skgSq3J2uj+UEVwxrrUMowlUYu/E2kBYwKXKYZ9TYJlq+0zKvuNJ
dg6gOTkHcbpk2B83mOXW10uplIWVXm5KBUTbskyS0A0l3OjwAdKSGJIC1tAt4w4x
5w63bdAVszRA4vSbkvPDsd2CoYXjBVdho+DO3niSM8uFzlhMXQNVYPXIsZDA6awN
hOQDqwa+T6W5HgAId4rE1ud/Nc/jSInSKpXr99Q/vFCXbek1jArdAWVI1B3amtWH
VND100fP5ptCgHH610u0oIrJJpAmti/lyUvzEfefYb1syfW/B2f7ONr9g2A4Yxv5
KUzBXKPY9CKXYZTvi0S3GVQUbLA7dW08aYJ5OKUCMbRF3rGWzRYh3l/6bE9Q4QNr
VjNd5I6w4HxvBg4jn4ezfXKARygiwjYABY180fjnkmj1dyDN8ntzoqCDgBxsk62H
AbSEqALdiK9lmpV9qwFC8uEGy4WoiXXyfnvaR6rTQszbiXEWmuFxYqavyQJsKgRV
4oPpiIcCerIhhr1XW4hgCTD5vnN5DqvJ6RhuBjAvC1hpd9IMGFDbKLQxou/fndGO
MMyQawvAcr3OjrMJPCRt1x4+H6701EY97Cfbzs8Q1ENNo1577NabzmrTUt9hwdfD
LNqTgfV6eNyapDRhDR+WvGVYZKoEfUJ+qsak2mFOzVcYNhSkEmUpzvuAIVBxqH3p
q82vd9/fmxE6sII3lOM5TRuCnn3d6L5Ce/CQhlNuTDbPYIG3FHxilGMKsEgzAC58
tmp5ejHysoZyWXyQiOM1bjVdG2hqZ3F0+iToNVU3Ie+Kayrs1Gwp4qXSkLus+Q1s
8YNvm5S4+v2rTbSFHDf5GSFxZZ6qCNSEdGln4ax3ti1QRC2uW+CysAg1iPrECpla
inCqYgKWJBcMX3k+gc0EB81Bflt7NL6nEaMR7l5F6Xn9qi8qPlgHnJDxokRbCjV0
kPUh9xFgctzCZFeUDimdkMXF5qJH7jUQevA7/89pnIxcJdAYxIDcm8tNzxNrVH9i
IiN2wm37R/6SdW8D7ePXZVg6f8/w/A9mv24hDQmb8KZZxwv/L490eVw3wx5fnX7e
i511QmEQb+fgdIVyTKAaJiE3sdPcYeMMNxBQmTnZPgmLOvSkIzf9geAKCoxvA6OQ
3rCnyekEWDgmpO7qAwnOxyzwCyAyVfV08vVmvFuAG+qkyJzcfv+b3jDg0gXFsNTX
Pw7uWYtMVgdWBkDiSCRE+FpkqPGPl8WtMIl/DQlnntB9QxrJ0uBXPV9aBT4pqMvj
ZULhluUmA+/qwd9EJLTJWjsCg+YZx2Gx1Hy2pvxWAH6d2001/q8iUkLepZV6XZce
35vdWohLqqBt44JqHQb2lWtxf0STPX6yPdYPLCbxgmkx1oL62WtvTssd78i1rvBk
lYGfeeKGQKaPjinG6DIwDGbd8rc652HoQwCEX9G1JYFTwVttzsZTlduGm1Efvg+k
fVE4kT9AnLQHHTg1ih18+cUIx2jAorhXHidwo8gr5sPsNHM6T1OkrVzQ0QcjE6zl
wsLIdNbssFVmNSPQaTERQHfOaT5fHET4uILxZWRX3ThHE+g1HpOtG25ttVLNhhBd
cCoFbpikz/Ix/IVPqxsBapzzTXgBeigghUzN++F2k4Z6AH+g+T0Z5thKQJ05MirM
CrsuIxcII1tPbcXI/o8BSKxhpvJRKLwCaK6WKf842G7wZCtmY27U1tTMxqQm2K2f
AFkF/yJ5F7rWe0cp3HyK+1xBLQyXRxJ5tIDUK5k+Az7qHF2V3SJ9cFhTkbnWBoiv
7V68D2HCbl05VSWXN+WOW7zUDMqfgZ5hskVQeyNCsNvigH8t1/ZOjPaa+srzneUx
GFZmGticrZVd++RPxQSXKc0yV3Dar6+FmV1eogjwzQvcQF6zXGB7H8F49T2WJhc6
7sCULTSI53ZnF7VaEsX4Lx/eOBz79fbO+LiUrLtQqc2ivJVrKzxstMZhtTlb9ZRQ
9rKVSFB36hMWHWITYZnQEkQo7kmuBp8G+/U2c9twfqlu6kE3Mk8IRCEG3ZUy/z67
h5ePtCbFy0otNiBa9VJ9LVesGZDtj8nF0YIbwm6zY+sfUtI0VY9VpqEYG+qw4bnS
V1f53hdw46MlHlyerqlsDZpIfT9rhGh0yaoGGjQDI/b1DPN8uLrP/eh/IWaL2lpf
svq4wDyORMEKqSkXPM/eoSFJhNzziffaYnIWFxmhkMS0umIOaVePdQbkKiCHPvrv
H0l8C9NaCZv8PE/+MXVz0ZJ3qecLtNbFk/05pQ+1dxlAUrkRMvzc3BbmViHQ+cRF
D5PiayFpCXp97GVklnhTBgFgmcSC7rrCtm4FEpkoS/oNGRa3GnW6LN+ADSolMmvf
97GBGNS7XHI61PYYZKuAdi6GDBMLJcAVapBU49ObFlR+5Upwl+u+41swJ5MJxKnQ
3zHDH6PIqC5wg8L4ay4DMwsgSMtEtONClzD1Jroyq6WejapIdWZuE5a4Zlx9PHV+
qRe0auE15DJrIZ2nP56qfJT5FtwUHaD8c2oc+cyqG3FD3ss2neoRg3SFgHdW7FFJ
aiRhlevxzNge2vHWANtHwXUEXxoXndtVVpfCFdFnD+HP+uqn/BdvItRpNuPqvmeR
s4l/vTUipRy+InR0LXXurjKBBh85yttLU98as5fmslKdL1CfNMUclaIVA238QmzU
xh/hIxlMXvCL8DtW0AONhx1dbyVe48IVB4sftbHOwKnZQ0X3W8/5y5lVS0OkSLPI
fSSmP/8xFLJE+3KoKS3ggGwPP58b2aWOXP6s2JE11ucOeM5eZb5omSbNFy++IJBW
9M6zD9l6nNXikm3i/oi1vPSECD9vpaR0hgGPhlHgCQhgOTjrLKGoT+n/BJKCTISO
0eJCZPhH5LJkr7zZRercXrDZbIUJWhXojEolKoZfLulYS0DDcOR2THoyTk6a84eh
en04y/yD3MV4YMMY90DGe16c0xBQoF4cZeDZ34k65fT8+aqMRLqDB4s8sqSUwHC5
uEn06OxiEvLFFFaM4JBiD78trVFKm1dNrncbgeqiMfKER/kQqrb7bB+3TkxQJot4
o/FShMK+Cq4i5Hd4JcLKEG/Yw47toau25Rwe6wB5ITGQardPMCJ8Aq37Lsy0AuK6
ezAL9Gp87/CChCnxt4VMGUW4SOl65aVrM4MW1V+fTXAAMYxrw+4Lrcp8HEd2vuaD
6GfLDOWQwsBUv0YNbFy1qfDD9PR1uMHcqNerumgGt1OE+6Qm1Un9Y44yDYql8YPF
2OLEDODUHKBaVqf/NqNmAQO3vPXYCZoRoDTo/AprWswAkvaE7f4QZOfOeaI5wsfq
v2+Ks3iCOxHKxErlHdGvm54+nIP7cA02MwZorv5ssTMQToyftrqJQAqTgDIM3wbm
zy1QOgYi9A1R0fbmaIiLvOLmlhAa2f8LzPWDSNgfX4tDObd25B03qYL6hhRBX0Mk
il4twzYQJPAUE4n/3n5zp4JcM7B6o5oaeqhLyH+x+OmuT5Fm1rfPA1ZVg7GUOxD+
yQw0Vl1xZUZNTW0CuIIX6gUvud8DvDmnKIFnABzO7X7Lw4EqRuzXEAxFGwsLMr1H
Rj9s4wSg1UdJmrPLlZu/vD5OSFIh+dLwTNVucjGPTWOcrvi6RYbBuIV/HZqHtTW4
l1wpsYmyV7PgpTKxR0wHBsKgUWFxGbkomRWDNwKGeS7PIueAJKotmFko53XrWG6C
dVkrcZkCn2+dE7mSqd4uGcrD0chN6fnYHwnrme8COx2/RD0M+CTq+UIlYkEYgEIO
7CNeUsV3bBNs1rQqt1qRksfBPQ6jtEeK4cMJubcxIXaQypgZZDGcxL+AdRx+nwhk
xWsXlDwKveyQwG1f0q69Us5jI/wvhLaWGLw2gLsgGbqZI1S95a1OopD+/XXyafSk
abOkfLwmeIKuZrPIcrCgLdNAtY3A4mc/WdjSnLl1iBhZWI9hAbgx227PRIvXOQdH
C454zPOSyuNENe+wmc1WxUPCCUDBUtO2JLQ7m9Bn17tzDrpxpyUZhRzF9rZfXmFL
43coAj04AtSEmupyHk/W9zmDiyE91QuTixiQlOlZuzzGQMXxcpm9Pbg9xTyE9CEi
qHMIupE3dPxBnVGoqmE2E5c6ghon1tJDdkUWFMPnAa3WCdx7nJUI2wYVJEPjbt7/
W4F2Z4mW96NLK6ye/4Di3EtW9ZFklKQHgqIzuaHtt784vnIFoS0y+Y6OrejalAx4
LmXv9QNSjXtdcOtNFo7lKdI+yfUGY0QWF2LqZ8lJUdDKJGtVE1eKyX//c64ghBnl
O6UxCxaNxqZcuBAgKxkfLHpxVLxo0XTinbCK27VqzwvaqwXP5F3c8GCrkEpasz9u
PNyQpEv/cLiUBvlA4I3tyPilIM8bqd9wAa/TPd+q5oylj+L4mm5vvKAt9qWHQikZ
IVNsSWzItSMJTsIYVlStmP0Vfx7aUo+kBASZoDEvr6u3plMdRhkf4LE89O8B539i
fG+Q4/kJHGU1Xz/UqiViY7PcUGmHx+31FTZlPXNkEoJx++n+P961EinUSLbDUyo4
YlCWrK5H/gGBFASM2wi2pESm0ZnVBh9j0EPcf9i1hRbHJZq+1FKaZoCk4KjiYcf1
t/WI29L+g5J0AsTMgfli+fM4siYHh1mqhNQvAYoxokyvH5hY77PA8c3LRJF1qcqo
sthfySfqsjGJ5XFbeWp8NdculdEvHlulULfQWgYiTRDa6gGohXgCTIsPyLww3ewW
M8WYwNm+wRHSQqQO0Ru2YeXzPrsR8T0tR99pbgm3pxcRzGh/uvyBQ4a2PfciijiI
bcizwZKIFYlFksr8mCdZpXrdhOL8jhGiu5xaz+rhtgLVTrh7qEVaXNKnvFFwd3KM
27Vwi5TpmhyH/eIG8RRnu2iR32LFCwkJ0NgR88QZWXEWUmBuQ4ZiiA0aZ7vSn0WP
Mp011xsxVkDJYl/5qoY8mU2ACu6lP0HqF+K1A+rvZpe8bTLDPv84FCJbwbdgDc8f
qcebl8GTX8f8o2HAim3SJzktn4wk6182eNmfdc07N/maE9HA2C9zkSsVKF3Dg+OV
6gUsuefiPJvcUADdft3iLZ6GWh3f/H2cm9FfY4FihqAzs8GEmpR/YGP2Uihjsu31
zhWCr9JuEPU6QCJeXugjl4EG5L+EPbN8y0htM2xg/a1MeTvyKAsZCtLOVJwekpT4
X1skzw9yP+wFMQe8LygRIWJCDEk0jSmpMQXkFYcx3lIIbRHmqE6JWBNDIj2DA7+G
FSRGktgtp6TBsBaMQcU4sT5dUKgVMRSW2sTE12qQiVACIvJs4VxoBqj7B8Wup6zY
hAOcWYfvBbt/kMY+OPLu/2Qmc6bF9hhUnoN+kusr9avjT/6jvLp8ZT8ytoD4dLQE
JWQP936UOZw30ErPOffLxbEHzMUkQSKjLNfhudY5w0wEuDvmI+n23FlQ9xtL8/Xo
rwALBDN1d1H93lbmhXwbG5Z5XZzGblo+HMzcyfRBrKj2G+oiWFvOg3gTfEzBl6ad
Nd4nTgdzWUeAsgsWaCRtdKXlPhjN8IqkE+CSZDdvZA2yhyLc5xV0I10a5AYeqmKb
c6mZLYwsVDGnPkuCdzYxJ8qJl8kU0qSendwKFAwcAZygCJ+HtOfIIPGZaConEf6p
3g4KttqUpgv2lMsLL9c+i1Uglqj1krgRCZHR7zofv2XigHRUxduTiWl0CHNT7lj2
cpbwre+ttkhihMUUZDe1VtsfyKKpahLQd1MFVqw2Mz9vpQmvo4NJiASQtU3oHmFx
BbU8YspTN3m/1DvEQwmB2gkZt+j4sUi/pA3yyNaI0RdfYCAXcrUzqDdTIANOYEkk
LbFQpF1BjcotL09rtiozDw7xw/xY7GfXaRd0+x6WeR7hJ9E2+BWha5zQulQceQtG
V+8Z/LYqzFaldqDT0BX+xFMLYq/VIPM6pTWcQQ/b278ryh+rOdxWrkOHNeEim9rk
WGfyMHGN1n8RKBCct1P0JJ4oRtJUAtfjFyySez/IoBScLNe1HGhknIsyYUIM0+VX
VZlM/0vvURka/pus61o0jS5sWOA8JyTnSOD0VwzxKfQwfEVKpncxxFY6FzWpbCgm
0Qvv5tvCYGKm8LInSzwaOb4YFaGjRxS+pV7EFuvo/NArb+Vx8mKqcHphSBIKYGD4
TEL+zhsTebghSm7x0jb1Q8biFsalLA+vhtb3IdZHBIlnc4gmZ3Z4ZbohtjhC5BqL
y3ZMeEMXwS9vS/wSnD8ENolmqxu3QvPyfC8htDtZWJSunCUlOUruYkX3gAxeFM9n
WuoQMQoMR+pCHgO/w6z+7QbNRF+YLaNuWg+IjL1FaV6SUe8/Po30/juN+pYCsuNG
W3Qbuz9lx/saSvO5AWhP98qguXV/D1bMiM6W30NVXxQ4p8rDMQBmUp/kNU6VpC6d

`pragma protect end_protected
