// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HuaM2uj5Vdeovl0Tuc3UOGmDT94ZzNQ6GUy/RnLBm+4Vg9ceuEwTG9QTuDUv
dopPJCHq4cKQ3tdeKmM/QGAsfZnSFlHiTZOf9H3DK2TkZl0q223pfhxyoCNf
5abeceoJhOp0YIEcMIkeQfJoRjm+J4jAa6g5aeQ5bcpodZoivhHU5UBGOb+9
D9+tLAXJMQWbVy6w/1mN99KDV27PeUJAibxW7UbU5AYqPxTzgA6veTtuvZIJ
3mYrwZBSXzt3tpbo6T12Nw+cGVwr5jUL1OUvJoJ1NPLvqQ0hAibZxM/5/yt6
ykjqLDi3N51u7qj2wcFTJmpGuvX3QvAHgRMKgdqAAw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Lmak3KcZpvkmKmAf5JwhsRTzignYgyCAARnM3I0R3QyuvgBaxm2fQbRdsk1h
y2BA5dN2zvdRvPdc2oxYkL1sYPMz9KkDlTGZ6AXkv0H9XBRdcTuSS5vh4/gX
keaqrrM/I78aj56yZxgWyVly9gzvsj5ZnBGRhYh0/ParfYhl0VVBsRHmJcyJ
wPcwbRjPurLmRetwdIaKeyBMJHn6kkOYAWtm9gpnHmmzRFZuWtmppWbHoKD1
7RUlhNRygawqp9PX5QIebCFV36WOgpnYkBQTT+DeM8dUqyEawKyT4OTpGnkG
b+RV4sE8r+niG5AmosM4pdHlBh4ItZuYXRmvXYIvbQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
oXPQEX/Rl/K7qFscXlUE3MDGFs5HlnXrkMMnxJtSfkmB/SfpTMfU3mqjS4c8
qETHEI2jE2tU4R9CHadDsLJXVMB85QMqOl8Nct9QnzH+XkdP0xQK/R4+46PM
DrOCa+sObNXCHr4Z6/vEGqAErIKc0y3AoIU9jGpHtp+sF9TjBpI3i/YqDhgz
i0jb8Z1mkBMigVvFTvrRmFz23BwKsmw5APioi93aCf8sz/v1yJrCFWnRLJj2
+i7mAKjwRJRGgSDxs08TVOOf2XTjGKtOq7kDx7pKYqBgxQUGyA9G5f3czcRA
FDoqwjxkLNi3S/wQ2MSXx2XVAOm8joSrrRF+Jz1znw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
QrsERKFwkQferGJKQN6W2TR80rZRmGIPKId73ayXBt1q19Qazkt49kGsOJ/o
DRZH+krjrt2E+bxZ8fgir1bquASyNsrFcTidxPPfA51lE5p3zt2nJj0UijL4
/ncZS2tokaOAXQR5TfVWzPxNJC1PwdIOL9BiEcIfcMkpedDwgkk=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
w1Xkk4VT9gVXKx4PQ30hMNZyDf5yZlnQKjInKsPCfh0SQEi+3A3Lm5RH5ejS
ZJ3PT/5Tkc+yWJowuvUy6P0y4EHW9iriM6rAo1kdhAHwmCQUelCJWwT8gidt
Ybi80xA91iLchVz/EPAjtvauu6+V2YJ7yCyxZfNKaunvWPR+r6VYy8jsGcc2
/y2GX0kEPOq8UFcKBOFck8R2Yzxz4HFshFfK0t/rxXzVEnsEoTaeS8IMhkUs
z2N+g6MNce3IP53Ce30XakGS+DdXZyLbUva2BYDFs/Hvkrhu6nq3Zp+GCDTj
0SxST7nPSA9DgV7xMJ0cDrW43bPYdzWVcECBTIUym3lU+LPJbYEUJ8FLdltD
NmdbzQrJjYmoz6I7VEYAheLO6X2LdBY+in49Z1xe5otR9WTfez/Z0HpBY9kN
NkmrDcA6InEM9gfPuq7aV8V8P0TBms8p7zXwtQhqZjfTAIDrTVh/jQZFprz0
SRv0hBkF1DSRukjvDLs0eD+Q59AcKcH8


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
B5do6ZQfhUVtCG4M/zuEXqVuoL7go3WEyupHcN6/SvdZ/ZZA/MRBcUukFdO5
3OU64GeuVCsoUnWEUzUc5rM9mNBnmNjA9bZWn/WCzN1W5pQN+RA+CYS2gim0
TLNCeEYJT1tbLwBQkES6s86v0iYROPCq9NDwq6+kCTDpVdMdhFQ=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
fM3+va99WN5DpnIhRwebHo5wxJZ7sRsvsIDINR8CVldB5xIUeztMnFO9K0TV
w3WKz0OfDYvg8gQ0N89GbeXXJkfRn/zUn18JHApBV/s5uFmzFrDZVYrT7vn+
aG8ComgHSSza1NUiJbYbxnF3jk2DIHP+oACPaXZWtydXHVesUo4=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 36656)
`pragma protect data_block
HVUo430JFtKrga4XH2AOOOZ7xYKRTJF4dlZ9HctTOEzTLM+jltv3RDSEyiFN
TSRg30QcnKYlyZCrRyKzWbZ8PsngfQBvyJrdDk/NZQg3mKR8BvJWw6ViAewg
rFPjqfE37hrXAfeBSPJ0mj1iZGErXem1NUcjYUneujgVXq+TorEwF7qKnuOa
kzpLjdFK551QtrwvXvkx+kX4L75tEiBFM/LR8uxPf/6ch6GM1GrtxJATukSf
Bg3GPI5aM+RvKBHZStJ4tVYNfsLpzkTZuQJF1HcpPKgIbPpWaiZCPJDKxCUH
xBgz9BQc9Y5TmOHT53OKS2MTkXTf8gq5my5Fn03i64Os20vulbUtwgsEy7n7
i+rfrPCouFlSJVQiQp7j34fudpcSDFyXgpkCoYfIDlyDiCcjOMnEMaggnxIa
T21bd5CnKydaVenMrlY6OkcSOF/K7VU3XJyw2N8KDY3KUwvtn56uPXwTSFcU
yl4sCwdbRhC0BEahOSjPZR8DYrtU5WDzR29a7LhnJePJs80UzezJlx4d06or
AYof4PBUY1g/cDrqBB3HmykiuyhKV4cD6iDPwd01UIlQbgQ4oUtI90ZiyKQD
kF6CYdqgRyN8rsDk6Mkwe4yYXIhdDc5Q9WrTXA4/W8Veb9oHkHNicIq8dShm
9z3CBSzYugouz05TP2sG1b/TUB5JOcvv5mLYd8VQQrkVQjf1F6FiH9pOhYFu
/AXQmriO9vIEs153e1nrXw5d/nqE3wvGg0toNa406hC9LzGxkXj2sYWzk44v
r3K+k9JFyRmuEV0IAVzXvXhMMiBppx1Luf+4MSbHwV+mjn9i3B1/Y2s4kFNO
W9SQqJDsQ/WQJ/ITN4p1/VZpqV/4oc8La9B2mZPzRN6cQMILmKXWTuxCnovk
wOd6G55oeCiKj9B393hO3l5pSJxAOFFdHHLf17IvIX4uST4sa1vRHN0FeATZ
RYptWVTQCx5kZSy6+DD6pKllJt/h/nhxASl0AZBRREHm9ycbQO0fc3ZHG1Pv
tjLIykSxLSXeBn2tC8xP1Je6L88YX9ZOJljIaasMfcD9v82+EdEn8L7IsKM+
RHMWuanEfG5Vd7bl9emVI9jP7utqGKVE7daoQRLaEWuy3DW88JMdosUFStF/
lDan4He2M8rOv/49VZegzfZ6TBJGUZ6f7cv08phxJNnquQ/2mEGgOUfz6a1X
vRqqVjRZP0hYu3x1K/19DtOiToQu6ix8F1JW0YrTZV6kXT0KsIOs65GCpT9p
YRSOp1YtNP7SBAZ+1JlZbsOr4BuE/zpRRQMGW4ghfgeK3IsO0p1PYn9ZZRo+
n1Eb52/lVtrDKpFCRW/Ont6iCYNo/pjIO6MuZkx6/ZdtOoigfCRDM+iurngX
Qv+mrz1G4ynVJXnkZteCZfF7wT3FtoT7LkZWDkQFg/djiXxSB82edGC69dwS
B4hM9Hen2Xn0tcFXz04dCX2JFcmg4RV9OY09en/Qt9ZpkNiPdTHKvaoUzwJ/
v2A3ew3zRCX4/k60VqBDhi3wPJ6w47oCLvDwD7pESZrR4IpxxO7LFCkKkJIt
5JhPeaQhugZgc20FEg5KvaTiH5IzP4ggRuGfgAc5jWL2pzzSlPiJcEJNhft9
i96JZW8clPqpj9tjT7A43VYCFeFouWW2R0dPA4sG/ssFrtsLUAvZyalJLbwK
0WC+z7xZ1kOJ+mdE8fNZsJHH4PrW95HTD+7pAe2gCiS3JUJP8nZKxUli8pq3
Y5u4ZOA8xYAPL6isKiv14RoBDjJmyE50kfPuvLwwSlE0T6Ck2KVPQho1+QLY
8PuIFIzDqB1lvId5E4otrAMaQEL/0aseAwxe1JSdj5owVvTvYLmdHhNyKB+K
b/SQz3yWK7oiTX/s9dOR94O9CAathE8irO8HQQMUnZcyBZNTgTsszhFaX4bU
TuZlnTGQYhGoUGDSdlZ0zd7xF6n2AT2p+eDXItjxp40MWyN+iac4O5Ankflk
DmQF0cu54pIdjpL0IBxKSr8zFsL2XUDQTfuHwCAAE4g18Lb/b6XLU+IDqiYH
jVybdWenj42P2DqOaTgo436puBBrkURthxeTBC5JhuUbmVPR5QQh/ESRFoQb
MgqkBR41jhXAkJjgO0m2G96KtllN2zJZQWCpz1ei2/6qf4NGZCNUUPgQzcWC
ZDZ9ck6XnSoXDOfiwqdf/ZYdzI2Y6eT7C7QP9VeEnOThJBSCBxZosik6Dp2x
0BcBPPJ9oZD7Kw9CCI29QGpcCWueKfTZR3r14Nx/LxPcnl25nZug5ikhpEoI
LfG64LCKF0caFGsy0mcq8Jg1ZlFBOAEr2vwAWSdDCVtrfjAqqa4jLZP8W5YA
ReYlJ9fou+zGt+bDoFdSKs021iq9FVacwXsbJzjT1/PG2hI99jRx1cT2PY97
ruIm7iaCg4lVa1TnqOyfGaKyVgCpEgBviA04/e8WIfcOuJLR08SZf0CYcnxT
9lxFO9KeYaGC4mEKvWKt41YW3kv3pv6TbdDQRpnpY1nisg6Au1A5wh6goMWg
lQ9VymkbWXE4F7x86Y4udOolmcv+UNOgMkmPZypVHpjm40CPkAcE6gzio/7g
YYgVGT9j4X/bEIO9yowKMw2aQUVsvBKuAKP2kzCQ48mCyBbXYa+aT9J7vBbP
l3I0GvRx5lJuG6xd4ZHHIltG3D3YmTv4MHQmWM5MLyJCoXD2zfk60L8RXo2W
h0TCEt5WOMazodV8kYg4y0oCMsBleDASSyTbuVa1RMLdVYCjyClfUimMnUup
Ifj81bh5ZUfkHvFvk4kK+sJB8nTrozz654BoJwzyFnTeGSvbYJJqy0LKEdqD
FvvdceGtd0k3wKunJU+2KxNlOa/nUDUk5BsLl7ZCD/mP7hDZVGJAKb2KPCc1
Md6+whMyk+X5Htg2QYohBFtD0cZxW99NR3/qIfAo/ALUR+KhTZuEZOASyU+8
uhDl+4/lFfTINfA3eLPMzL3ZN9CBpvft17dz2WuVLHsaoqSI65/CeGC+NqnB
JR5W4N5n8sEi3atYO6Y0DJW19TB3zGqyotaxUG5x/6059xDZFypwIInkwHJT
HpsROYz7yAEXCnIQr4TpHVwXV5L4+vkDQzkyoDij/fmvBlhxFqTtLeQkhqTl
x+LlWVTzPbTFaRjVcPu2j8Bp+Se0QDRqJAk3JuOqDPF6e0vGGbrLqXcZmmas
vA9eqRXeuQLth5wY8rLgZmuJDL7qBTdM72JMcW7FQ2TKkH0OxGZ6Ap01iTG9
/BjpCPTSxhGG6T3ukm5zIT9+r7qfcp/wnUEYxUW0aV4YinsRVQOnt/uSi1XX
HJdQWyRmDosbe7AxDhlX7/zt3YSepO7U73Vj8GfO2tzpC+LxhICKkV+t4x4u
APpBy7RYOXpnwX+5ZJ8YrODCcbpFbCx2nQ9an+6t5g8NSsF52pLz5vyaa+1U
7woT7Kdu7WZEbrDNZoDvpx/3tL+EazH14qG+uxEJ+GBynLulA6pcM6S2ZBTg
GVrKe30Nc3csG6AYcJtsovxP0M6mryLMCTTLMtBOtrzUxZlQSOLF5SllXzzY
BW5hADgUltR8KE0vAZ5NHc9AK3bX3rW0m4l4oGP6M9EgnrAVZBgWrmboWXQJ
xSmiFxhEoZtMtmIZGoKE36xjVWk6dwkMyqaLIBg+PMdI6eFhmdW4ylFYHDn9
Vr79isasKx4/G2sPPq6avFtwM2sQU4wOzgOpTnprz8UFkYAEqn452CqdugDd
PxBnSdEteHWv3FFAIzK5sbUxreL9CjcI0qu6hegsZCeKNPT3TY2riVczhGE2
Tl/++7eJxgkW6sG+qbFkB8tUgjWuFWW5mOC1Yp1Ioee8vRvUQve1OVu354MX
IRyZjg+cl0dMhhl3zmlwZrmtKEpBnA5y8ymlyIwhsSyF8zC/w7Pfqz+HwudU
IHVnBC7/LNP7aMnlV6n6jwP5qbchSgQrcDdWjytHlSKAZw32+xLi8bzc6VgJ
ssRpNi4Ti1Kvx8bZNDFAT02F7FDlE4Bia/MY0B7Kghml1R744/NYg23sQqoC
xJ9AHqJIHMs7yNuGS33Aojcymz1OUTBTKFoeaLQ0F+JzS4wiLVgj3t78LK+D
513FzF7m+36d8op3pht/hM97LWTOXuVBpqV9ZLVmzfmqAlv/+qe/OrxcVr4+
/3L4PmTIpHNnnS185J2kILShtnL/TlJVTynXan0Bt+cKFdhlYyFJqCdd2kj4
mapip6FmdAlb2d73VBudMztbsy0G2SRXBejawkBtPnEl6LH+f8MyKkD+5+Z9
Z6T7rpb/e6jZP3IDk+Ef79krYVkxdXZNwQaWFb8CosjNylzNw6phKPLdrK/S
PjqNXLCaLGRat/U8ehxY/nYGq3TNyaj3iKxPPJ1oKz98jAzNyrzv3xyzY4nk
gV/2C12tHLTYXU5HAk5OJR4qjDUsZ1Br+ue4Ytil4O9/uptV+OGr+VKMl6uv
sBQ9OFFhCR+xSCqc4K/MTkoJAHzEbqE+0JIust99o7yc2DpEPxiEKMTvTMd9
fMmkn8vFNnPJMjBNgmvNLvAcD5iFWT7yRzymKYQpszkIH2R9Ov1tfROSWxSX
4p7n6r3FRzG2ELS744XbpEKgbUwGLz3xbxMhvXBihWrZqReIkV0WOBUabthb
X3Y8Q4lkMobdvE+Pl5EorYQ2rti2y5RTbktBQEWb34DvNoO2DGIaxOYtm0IO
urTlW6F3tWuL7PG0yLkNt2vYcOezsGDbHv45/0V/ekWT1Ksncx8n9UYUaNaw
ouvxyQzb5QBe8S6W/NYR7wNvvXloruFX4IBkndkXwDLA7OyRYllvED/imxxQ
Bv6YWZBEVLtjf2ffME4Xos4bYEkzS0N9+JjlYqM4tnG9Hg+GbAp71/obPocn
/thn21VQTtQviQNpasmDwfHZ6WH7oJUQGIwwty0M86VikqoIHtiqkOZymkID
reEoDkSICe1mL2ZvxffISzCwOqC1c208LLn8jNYw3IMW3/cc8j/yazsBA/3c
C+xfJyINvL3KRJr8RTPV9tXBjbUJraFYcPxGj8h6LKeW1ZcZYrxbFNaMzLpr
wvSMXc56KzuTy11rU6pmsL1EF4UNYT+U49sDd+DgDLPEqDWyzSiDPkAxK2+T
42PDgxp2d4ubYoQMN/MZHgeiHOtcFMaGX3GalDB8vIoEx6Dli8tJzgY8PFDi
DHNE209PUaDGiGrvkzqO5hjwDKKvp12vT303336A3d5JY44nIW7edE+PG+X+
u4N6vBDj9gUsDMMHZO2qfXZ2XpV+8cwl3qpO6VPLyk/xlbTyW6UKHOLqLus1
irIrRol468SqHGV3JHPjLYjMsKl+v2a+Hy7jd/+qXmWK8XAiz55al9Jn2B+S
hIpVImdRxN33KFP5jzBbfij+lXLszHSDNZBU6I9rzdul1sgXU+qPb4spks3D
i5x8rpMhbFqB87Cq3RGrxwTsqDywSC3/HNM341tDMO77v0TuB+GjyMLWYUeX
/No0f/Kpr2kE81ELZ5U7JuWhJZleS/qGTWnV1fJP97beuuwXi1Kpsddx7vTM
zfHfP7gOf+8E7mnmZexR2OWPvoB8ZmtDNc/K3fJ1K89tW/LChA2dYW/VCogC
BxwtuRMPP2anP76o4hQMcV0e3kiTJGo+9HcXoN9mcDcjBQOVz+h82TsAD54k
zKs2pM0zYOSeevKqJlTPW8aywSektoOpS9YTz2LIvJzsVXsLzkfJs6xyIX7O
lnymNGYpzZORHEtucwUCaAzUX470liGG68Ariyi90+L9pnSmjvQzRZMLuzSF
wd9hXSCBBI01Vkl4kmLhNyPRJnJV2VMEiJ4AJK6+9iqmPDqvQ+U16F2IhiV9
11MsuNX/PU6fnaqR7TcczfkgrcHO4oEUvU3LacdZF+QfSLfzk/Pfg4TS/ncj
alrATzyYc4PC75btDxwuDee59NE7b3iR6kvQ3Gka6Xc3MMNr+1JBtR45ramU
tAfWMDUhb8aATBGurb2mVeTUAxdHI1yqGLtWVOp8NQKU1hKd+BvJtPUlLosN
4m0oTGE5wLJyreanX2D81kWx5yZeMM9dA7JTYb0MDxp/jsX+UuSOFygQ054X
wnVnenG6UzwS00ZAgDtIyG+C+L+gSymnK6grFyvX8bBQDbL9UJPXPMGZgS/E
BMT5q4UKNFnFOSHttyzXYw1o3jzOafrOQu+AjFtkVbgqX78Ln6RDXF792WFJ
5UrYx1DH2ZqPfOpsYKzLSZp7opsP+M08l1YgRRPhfHa7csXB0w2Oz9eIIddc
vpXoIBaJibteT5zEVQMBdjm44n+Cb2eWdLoXaw7wnaSTs7jKL/Bo0dqWITVK
z8lnwrt69qdj9OttJ9p+GZMNtqbZrGKM9BRRKzzTaLK6Urdf4eFlPjFkD+O5
eSnlbx7lt9yUBslyDy1YZqzgDnTBaZNVU3P2nYOGHvMBP7Th9EjOf1F4/++H
GWbzW5rk6aiDwlIqz8spy2OWyYY84A5ATjhIqVuDAvsEp4aVkkLlW8e6Os21
JtRudeK52Kysv2V0Erio0Ofv65ABo7koIKgdk1+uN8aNY76FyuXwrwHv1DFq
QZrg0he3Rk5I7vzw4n6hI3MF7VYCprDq2Ibs59aZOkjx/e4SypiqYpFT99a8
HS16J54ilmMSvpKFSEo/N1YEPfLm5nkP1bFuTUgoLWYC1tr55UwtQ8cxxXNl
NcYsU9/UvjB4rKG5B+grn/aH77RYKxdUIckoTPbZDS1uNxFRzDgn/nCpBCaQ
AztScr74/sy25X7WRVWB0CCGzsbwTWj4iHLdpee1X9z8aduU09T1YfwZP+in
yD14FYfwWyH52sfiVwH8igi315bUTh/8WNUIXkU4lv55xj0bBETeTF+43Wex
HP1og8t4Z62NwFDeJWty5eQ7/tvwzN22Emu3FEIJQTNGvx+t+apF9JCogyo5
q5D3b4VWwU5hCo8Q2+DF3psZ65bKIaYmnh5uvDCmkYw1pejaBgTt+Mbowjw8
v55eBhbalUY4oBbG48IF61Z8LT3jFJmE1zNBya5hV7Mefb+pd41adLv7JINe
s8Qd55GQftvbHfllK8jOm9a4Pc6XpdSYZZ0Fvqn90QDwHUCKIIKfTubMNfvz
ewEVybEY+T0UuRvFu5RF8KMhynV7WE9KfjnmOIP3Z2sZsVNaJTEA60NBsK27
bVOZC/+TjqnzVA/UqnyK4iwEfg4hT/4MEbOwl4ssfToXsNKa49rCcyC4z12p
HYN/wUTBD0uAKwmtPe7aosB/8ar4i5/K1WoYiB6Wi8u3rOND1BX+nYs7LGpR
d23fPDXSLe4mqsgILuwbETH9p34iV83W6RTjg0yMbbEQxQssrjANNBXADVHj
bdDdj6mdOMI75ml1p2BiniacuoccMsQOmbfIpkqZjAt65v/DGSiEDJQ5bhXO
C/uX0TXW8zJl/CWJ7quQBQ/v4rc0mnosUlCd28JACicQP0+ArF90wsAKczAM
Qc6fFHDCot8ZHaIDNq7baMfYuqgRKYJStIYPdJ6IntZMKi1Hafx401i8pect
HEJou4NJ0pQyEocZGHHMCBfa2ORuI3zXcytZqoYMO0O84kuvm/m3rLFM3LNI
usRIB3FJEEtA4+CcpliXrMUqBglWRxoo07dXcO96IxrWBP3QMA4UD46thpR1
fjjFLQ0avx4A8j/CAux/3nJmvIIJnxd42IfTYD2HXugiALtPh7ZvBF3iEGYr
ij8t2L431dOatCLSY252AJBNCmXGlofttMtXpkoB0D/hqzfGSBltAhT8ocEl
sE/5/byB9uBosc701rBP/bdD3ee0ryZ85f4kQA+t1IRA/PjloPRoPaSGUEf9
GAKWgdPWSA1LY9heQuC1PJLVFoDWSO2WithwwVE3qaJ7Ii0PdmFrazxuKEKc
qv40XZT+YLLOkZWCjgH6qnUQ1JUl8d3UZjKP9EGnT0IPO/q5wpV5VA+Ii5TT
4KZGaMujJ83Nqi7rI43r4PtFMNlH46/L2QS8XnvsNWaTF9FBG36WWqw8Oc5J
Jyu7UKv8Hcm0vQ2dpAyzDktVcfZqZCcK4ZCqdkpBSHR4061foBhzFH3mOW9C
atx63EZzIZEh1bXEqmN0q1tRP38HIJZdIwd0JdzHwknMMhowHpm3lG2RTZti
4QjcNx2u/CqWMcNgq/ATflELCtlfHw0xyiraelNEDwoHmxCKOBgw5twy3soV
1fbIZHXhNip7CGoycNCuijOAHuKY7tVS3buYileuD4cYRiO6hExEJczTh9mj
Idp0yB/OgKIPGucZx1cc8cikFr27Y+ZnSAgjwrrWp7SWhrPldg0mbe3kcaZ4
+2d9IOXf8Q+VQKKU8LUuTMd3vUFmOoWIyMxE9XIVw5evS9u+O5kNqZ+ZFKh2
/MVo6vvFn8fmD/V0AzRcvMnGZ1xWJ4Uuag1kUvnJemQ3cwtVm1W4sMVMICDO
WNWx6HXQs0g/I+cZVcGi7hAFyf+JLdDaPVJhsT/4IMJOpaPPkSMEdnCHOVbV
3nhWHhhNqvRcCvA1fTdCQJWVb9mVmZMwJCk5r4hSHHTG/N6OQTsdjl59BEiA
kQ3TPV6lU9a7phjP1Xa3zhdytDrc1HTZv7VnCN0HhJZkadMrjjeCc25+W+1d
8yebWnE2W05BksGq37JqeSsDs2J0VkoUrwdw+tcTDV10qSaTbp2mkX4R/SOQ
W9EdQ7KhuwBsjIe6HCgm/yf3wpZ1fPNjet/d8oLkxOL3MhV56TFIMkjDSSrZ
1MNOYQW8USUZukvuAoIFUwK6MyICyGFQI9zE8PA8oTHu3DMVg7bUDzWMNBnw
2NWmLJ4BAe78f5agu4pP0aMKzAbqZkqTtgRA+6Nc4h9Oqo3bGY2TVRHjViaf
v6A5GsMZ0VDt6Kcyc1N652TDXicbHcGzITaCCeSCeIB5cJRK5EK5hAjCzlXf
4mPoU9DoMGz8f4smueq+Uchj3WoOV9gSqT0udtMKIFrzkQILrJwnR805TUNo
fRpXg4ZSczqgSE0V3bFeiCkHHIAiW27PVEF2ZTr64uPiBvquxgPzgLoEU7QH
hvgwOJy4dUc5sB427GiSlfqXmKlDHZkPSUUXV4f8JzH4qBwoRLdcePS1mrW/
3YCLQ36xdKcChjCzuIHcRHh0H+TxuyBAnXBOXT2V/0uW9ZrJNv0XctgtWREL
xbfbjYiXy0U4XGR4fdScjUNCgWl1s9BU//N+4T5FUQTX0c+e0GAtZdOYNY7f
l+n/ygK+ahqUSJlyXr3X5WpJBIlpPfJxFvpr1DWssWYYRMMRE66g7HPlEjox
vfkjPERsWRgTn691SL3E+98NT648dZwEy30rUDVRJ4cY91GlB84vvG5qLzZ1
+ErU509ybHjjFjlzGsiIGzN/WS4II8NI4Fl9LOQcsUEsiAip+dzliiTu+F4q
FGejTpXP+uyQyuiF67+3bdfErSKlIxSSGWB0eDoCcTbDIUfvlGU/g7Le6bT8
tYZzNfI1HDGT5Y56yojqJePg2T2ZhWDzgJKrOFYuFWVnZHiY3IGfiXC7RbMU
RcPhwdVq2LXDSBqmb6NrW2s+kuVgHMZ1M5EIKm6v20bgIaOMW+RWONVyhlzn
zdefTPd64tspeY/ugRpOn0E4zua/hP0Jkboyji+lyXJpZuz58C0X0ntt8YXh
LaVTzPdvrR0ttj7nCKzYuSxr5nbs3dCcqNljZ67KJNpwrWv6QygbsZ1sswhc
XiOIZFkH6JSrmQlNwDPs6f93ZfbQJX/SHXZI0kspIQ1z50r5lhXMEaL71rat
SIP98T8dhUbwoJQ/rrmZxZjotJ5D+UbvERLSd/s5mZ8xpIvb8Osmf6ULwMEj
8obBg6V7SUN4Jmhu+v39X+O7tYcsYqZ1wCbzGFeUIW4R5JqZrVeJOC3E7bcx
hooYEuTJ5GBxRubuIRTSFVOjwKOz70YbMz8IcPSqI2LFq5Pd4AC9Hau8x4Z5
cfe0mR/65f/Hp+TIRh70AYb191ixoWckXRN0Gi8elgXfmjUAS6FMPkm5/lg/
RB289+g5FZ+qPUtf3fRpYcvAeHP4/u+OwxIPd6o+wmSrxIjHnaS23ah/efxD
wMAZ8RdDW76lzN5O9B2KZpIL+hlohBgv+oMb4dxQc+WXBxsRUgZoDlejewO7
6J/hjS+WaycPDgmpF/JytenhcCdrham0pQqoS8M6IyFxD++27H/XqcFqoP6n
WzNZqYyFXv7KD4ebBFx/f8j69KbeD66wBqlty7oy4m6Xo5MGwkx8Zs5La57T
o8ElgoVHF+ALGrOkmndZqulHwgfmszsugVgKAqglG01BEjlyW4Qi4Ubjn0KR
qwfE8ACa1e+cWil0iIzimjTqw7vATGuv4Jsr5bt+UF/nUh2hDRq8APgoMrJz
0movvQHPGu/n0bGrChbDTz4TZycirgveio+Y2yHH1e+wBnyFvrF3GgnJzeJM
S7TfsZOty8sC0UJ3COGW+KwJhTlQaZsF2uFpKaQ9THrDTKyMpOQ/ODR5FHgH
xGnErLB2HCe/WSKjwud1rimauz37p79RpTgBdzvZm7n9BcQd1Ghae4et/ToS
QcwSRn/jKz9AASUJ7p9nC9aErsI5ia3ceGUrxCdYCw/mdANqFt33KWO8tu88
4OmfPy0rxZ/638kI6EUouCZmKSHntdoOrCy+udVmlQPDxiOubuK5K1IpGRcd
YfDsXBx3MAigdQ49fINsZe1gRvJ3r3X/AfJ+O4ytrB4B1LUfrKILA1cJdU2V
zk5f0etCVVJMgulf+WwbCrErJRFd0IReq22m9wihlHxwAPiHf7lKDt2DicdE
pR4DwUBFXnRzzAXgwtGubYUTHocaZ5HAO0+8TmvShtVWHFysRkWgLOqIY/yG
m8DoyRrAW5u58DuTBFwR/C2lpwXuoUWyUuRG/hsYc4ooq8YpxP5uKEixQsp0
H95HJHFv5c7sBDfNMkVm/gtGlnQRfxTsanKYz5IFkYc6gpUGGjuilMvXu8Sh
p9ICeBDQJ2f0Kr+nJ4Wpij6JN1/rnD6lEv6ptyHoqEUgM9bgkjf+76bSF3Xp
NA94wx4vu2Wxbk9dwgOklGeLKyqqnOCMQt97pTpxpt0Q+Oms7cwXsW1dqS6C
fcaWxJzhL6hb5OEat9RJMtWdG6vRGSuOVZwRiuGm3kswMnOyCiHuaIJsOgoc
MXCtntqkJwQi3xjK3cR3uvpYmHLOJEW2fLNIimlakwL8RfUcUCFAAnizOrMI
O+0fFNnzQyRzZx1WnNa0BHJXOVFwup+39bbXssa+YLlNsY8/sNm25cKXBj0n
a7+5+MW64k2e3CrF0ej44ceZrIprLlz84IO57ywa5zo1trbWgHTs13u64xrJ
VJtvLXYR4ZHXczdISibc4O5mqXdU9xhKTTuY3RjIk10BNK8d+ydz+2ubhW3h
KYk+K3Pu4Tn1gBw4laZZsrMEBH4ccQvL1SgX2FUkFn8dsnOR0VfIlJZIwmgm
bGbw39xHOSdsMVf8/Ui76NisgGOYZnyRQ+MDhTfgarJRaos1R/9zXjoDLx3+
G+V6aZTSbMs4HMRj56ef5TDfrvVO7aIrdBan5T92iL5XOhx3o2i0sBi9qK9a
rpzpgRBeaHawQZ4BlP5OrDn19JaEZtUUzbzUMBRVKTYKQOpyU3FCD++K0ndQ
6RRq3zb0866lN74LA/Ctk7f4x3rckDmM8Bq5DfN23FKRShqVnU+evWF9xXtU
SNlSt/PwItPk9ga/wrN38DnQ2RDaG9qNI5FSjOyYKoPmBNuMq84LHJ2KV8yo
1m4kAucEpXHd77+jAy7oFmg/+RFHDr01TMmKqFkFbrKQ2TsoTIel5jT9X6aj
oMvOG3EmO0s5tXKB/RyqqUyE4x1Th1QJaGF2vb0IzzLLexho3WQ9Oo5sucFY
+83hq4Uf9jOaMfWTO9Q9QEMuhQ1iZN2TUA68meXwJe8hOItGtFl6df7cHDla
0I8+lZeI1Jz+GVTxgOWgGOAoeOnrRm+F7kZ44WZYQDuXICwNZ7caaR3qmbqY
HtKO79ddF8GJzSDr6uEAbd8GKuX2KWKRRY5NFPR24SNqOJndNntzvE0ufsj/
6UBApZjOL+DGS6sczHE6yUoSjhZvApW/xSPn3iTrnOAbSZCtzDoJFYBAjBNc
dtOm8YqMnJSMUTNNhoN/tSt3uBI9dRPBeUk6mE6Ipc++EduRcrUkPnm+E8hw
oRKTCNhpZ8whazTBc2sbwvul7g9kp3UzqcdyoQJiamNBZM/6AjP2ECIXAgxB
hFHRSYrXnGsTn+zRCKpL25jzbjaWQXHK768FCLJhxkhcQDlTR1ZJ2NCRSc94
nizdufsw70sF74eSF+UskDmO7A2Ta5Bjd+YmXIRA++lQXv8FhWNQccdbns6n
vniyIYHp6yaqsJUH8AP1tr1amA5iFXN9OnxADYJuxhVEcNeqXVKtldn39d/a
TuMkBmbAX3kljVmcd0NomOOoD+H332PZuf/5T/ptnKJOPHMZ1JLh83XgRI6h
21xDSvgNTwef1JolrttR+2Ehr9RTY7OcO4Wag2okAmNuzI0/aIZHTUTdOwYU
B7ArqaRxiG0iZVpYuOHrPRJS87g/mk0fmN66EjAWYLbvrNUzUl1jJ0t8Y/1i
1z2iuNMJR3SCUbhen8lQEwfrGDeM+GMT1OxIU6xKnJD5DGypX7sPPoN9aaxL
rZgaFeSje7RnaejucLP5qDgiqiSENB8mxUjFajQLJ6gZXqjJiZMTvDuyx39g
vNkB4CDr4OKbj7X+tlQYbc3IKb62gsN6ssGLnu8LL1VGr9vhF+u0ey7r+Po7
SoRI1RnlLW34j6qeawj3VmYsEBdH8GgOpvqiRh/SxEt9ZUa+Fd1y6QqEKgZO
99QALfcTFlQj5PiaKo8PbLdSKRZNG2eskuHbulJRxeY4hVE1yAYGXVFKY6z/
FUKaci22/iKdBrhn7ISNitjY7/FmsqZynayzDWBY9zf8KLb/nwIZCB1LmRE0
+wAKFtkzIFUEprDd/F/2tsvEytvVZoipz8oAHsIyO/vLLA0iX9PIwjJngbq1
vt+kQl4Zo6p41ozp4d0gMtBouxqJytEUTCDM4MEWlMXxygtbzf9KwAadOIdc
ry6dCvgbD7v7p9P7lMWYp9XTWsA8qjc1OIAy6fuMg+4jMyB2VoqNCgWrP4cq
VVUfyCSfaEOweXsG4DdVxreEP4HtCnwC/trQ1nyau0Ivf4SfAiTIqr46WrN0
08144T0HzwFNXPOP6WH8o9vtlZ8xfPEGinpcCSR9tIeaV8WgHemsqQhbEv4G
roxpbqyCDW6oIjrqN9smo20PAxOxoo/hcUHHH3mk3ppZncSzlSqa70YZ1Kt4
CB83KDkXuxjY9MX0aQcTRizcWruGNL+Zfvt9F5pbcwz2a8vt4bQ4UW0HKAiE
acgbJtgStLrA7/mv9960G+BMHkxfOyzc0acVkKNeQvTR23bA/6BJGFecAkdz
vzPDJUq62NTI/Fcrvr+eMLQsXX9K8wPbKJaNMIt2FvlsMHNRE9zIqMMWxbK7
EEwKvNc7qirtFby5Atdlp8b5lTz8AnEqNHMoeZa0NDpIgc4ZRc2C6FEsj0hT
W6BvDqBvgJI3GXCKl3SYhsKs3AfeVT34goJVxI/LFcpLDY0u7Ij0KErvjGT3
tEkaB+Rn11BcHLD6oYQtJfCJkRq7HggtZkK8kinG2KtbHgHYDI1DFB6zfCW3
gbPMAkFCeoGJIY8wfN3EMvnY4X/FYacrol6fMJhLrP/+AIesq5mEJ4/YbHoJ
3St1/T7ipI7iF9NQOAV5Ierhbbd59OMCJFFknr687kxwkvp5Ev54ZvaPURFw
7lkYxTXIlSqoc/DI139nZen3yn9L2+BtnlArBR+foqrLIx7QSfILpFviR459
MKplThvhtFvTAHSf3A0HvpPHjkzzlDIFVP3NZKwXAmXVg4OIWfcBKwTkS3Vo
uoSfWt7eP+3Sqq7uCSuf+yyAgoCvywTsAayrWC1mA9a4IovFjsgRVJBGY3rQ
s/IWhejcK7V6dqDaf2z0a5megRLkqOf8vgdeVdPJWORf9MZGxiCRZa17V+f2
laroxyvA1eZbRAcWzlgNikIkfg/TZOOYoBWINCC6bo4ZSPK32W4Ddj04VB1D
3TNz9Iw4vHvFD1FwZJtTc7atJw6/x7iXUqLH/M6kkW/QTAz0/EhuwIrPihXo
cnygSVp3KC8ABaXlcVQt9PmrKrFOkyumPIhT5FjKYPMTlCibYUSksB0HR9L+
ItIVMWcICJJ+TTtx3dj4ApFt1pi2ZmpY/zgFgdUXPdl7Ls7ZNkgDJrsMr2nP
Sc+U7U/oFKf34tn/yHgB2lxABWWAQtwkf0RI5kjih4BodASrCz5dxkjUH5wC
/yWDCatA5olBo8CzGZWh7xtwGGBvkmIxftQUY6NBKHBKgzLtMtN0GGGPcaKQ
RJff0SJG4EZRRb9LM/ugwNVBwFrk+9G1+6dx+aI6+r0ZcOmPsY+q2FPnU5gZ
5GDfymVTrdXCizRiyLrFAlpj6x1ImNw71z9T7mlw0pMCNJEK/HQPifZV9smJ
Z1RvEzkZCw/kwSJ3JS+tPixlpwav1ZviaRxTjPImGufEyQ7curNd1DiPZzdL
KwR3BUsmagIATL5W/fNBxUv5ic9b8eKURwM2WpyrMQr59QgQdHQQ8N3nJgPX
W/0D9BZUJjwfqVBObMXv+HPo/66NiNqbG6Es366Abw+NLMjHVGKUNtIIEG9g
QVQt8PrI00Pt5ewZJswWaWClQxZLuyVKEBdvK3s2vaw3glRoSI01zByloAph
N3K7Lu1QRCzp1Toa1PjLV41ocYE0eU1hw0erd64CbC0McC1ZZUgJT82FfbeB
TfQRKWIOUm5EFXsulsUkBJoTugXAX6EBvY66PJ7oCWSKJxXo9ZHpauwOYiEx
foNYw1Pssp/9NIKERl6ZsJy5mUxEumtpfIPxr3qDeKYyhX3BSkqXp8u/IeKI
Y4lBvPJbCVZkHSPPxlC6VR3CatFEPp8FoCry1o6qxsZvOTM16hX7Xikfqpkc
kDRv3bGAdh9HlXHgVMhoYOOu92ulHem6F+A7sJaDwQNJU8AJFs3lX/wH6N7M
CBR8BNcbxPcWfmTfv9n2JNLDXurErDTf+s7XjXH3jD/KDYlnVGRdPaO29+ql
xQVtaZAmMlnj8BhZdFltO14X1Ua4mxGbwequuSC1/s83UsL2axUS5pM3V0U2
O8LNWfNjCWvtVQKMpZQZ4JkQIzXsSfhWWzboEA1plfJ8KfiI5VOozBayIiI2
KraW/xLn8lCszJyCNhDES6eNGfziTL8x3LQjaHbQ5ZUDjr2HZpDoGQJaBiU1
yWj9WgIZzA2yqppdHGkdP732zfmGDzflt8YlzzD4ymJNCVXVFDhcSfQQ6e5N
0TTpn/LGISi3DdrlpPi1XTY1IPj89jlTueOZiYk9Dg9ww6gfNG/ls+sRZjSJ
KPF6oD2UZKeQy7JHtB4778N/9sN8TzdD8/sZT4aI/Ks+gd1qJ8+pFXhBdMkh
mYjBBzSQ9uhcYTiecAwrLanqdZ5m4eDWFULsTG75992CmxkDLwFg07rzWz1j
tnjskXsb6dxcX9zD6rq4hOdyYBFm5bQyDGCefCIiUUPuEu54ivpzHgpjwOa+
DstKgMOVl9s5B4xkVIH9fhHTh2Mh7ZzpSzXrdQ5I8cTqOL+P1UABKZP/qSNZ
AaJHFUILHecteEe8DJdcw3NH9nW0rEKW5sl1T+mvmF5mPgDugHUUKoe+yDTy
F/xbuFBfET0QS2HEHhOKWEa4vDzWxxy4dLlXKpTVdHQaNItO7sJmObaDAcDI
1oPTurwmX9sKg6adwEvfFv/CfAOgXH6C40nCntEiJW4GU7YN5ynClVTq/eej
aqp5wKccrYe8IQz5CO3uoKUvuE0BuwkFEf+rsCvAnDjn+4VthoCjI138JmPX
wRNbiuDvViqeoeKmh2vgymgL5BiMhHJht5pTvSZGy2y4s7cofJHtaxgcxYYK
Ka+CzYItNQ5TKJvUsGxd0+IUhREl2OvHiDV9OJV7en/gv3tvrOjKCrykRjOE
ciOMaqoohzuzfG873iv5LnE93UbPeh/L6qHUditgc/9/IXmyMCi4SlhLOVU1
MNl6Vy8XkCOyxydRN4PgLi55i8zhd5zOpAPw1bVZW5fXwYgM42tg3x51o7w7
utoVqZ6yS7yW90Yop/wgtNbBDNqxRSnaJmQM8OEDOHOUUxQk/8bK2lqY3I3k
TFdaKiKQeXYt3wGdCg3N3KgVzf0D4ls/wnhRLo/ulz+L/8rw7haDF3Qb7kSB
mkmi/lDsQBh3k0pM6xKLT87c4fhMhmO397bVHtYjtVj5PeqEl1Sw/gZstSR1
S2rFKIVOPm0OrHM+ooYL/Wdisl8MNTzhRj1kG1/UrGsJhasFwngPwjrTxAK1
kfGbOIa38J0dHObTHg0WGVTVhVFODHlEMh1YY6pn9Ml0dPdiB/00xPIm/gAx
hATumA3m+XaLaWwXKiARVKEt0eSFSMz4qnbhtG7hNyz8UzcpaD84zEG+TGwK
/Yvc4cL5u3vVEIAXWnPxL9+X2emc3TQPZqnglfl3vjWQQfXfy4PVdmVolJTF
RBmvCuu9ZxOI23KH4tzyiUL5fVfwxuQ594rou18ge9YVDZgTNjkdXr+PfXIJ
ntJM0OrcxOwlX2hzTPRrdzX320PXsQ3e1y5IY3+H2kC7JA1iU0Bw9OuDD6xS
bcokffHYGGBdKymn+QmJovQ3j/jhIxULkmO4OXeci33uNp01O8JAYx5YyYhB
ssqu14RRCC9G9Z9fV8t629IbBUMwnrPPG/1OxOh64KgcA4T9v/Ft4oob4N3a
St70PCFNqXIdVogaX3nxkPA/kWlHtS2K9hXuQ43s1GBv3DOx3mTnw5EaocJI
FSQyh8aoAqAYAVHtrH0077mPiZNDABHmGaWsgfwOc0oXJVdzHeTmTOar7gFu
sa5yByYeenw5EAhQ2XF5Nm6BaiLvrefuMylLcG0UVhE7/fFA+sTu9ytmF5Fr
yQyLLiHF0Ckp/cjopsOJZZVQHjpG5lfGTwQC54UVPIzBZUAILjFsYQGhIcjN
zdBqVGs3PQl6vPyQrk/mIkrdp7Vyd1+U5AEg+htg+QxolOZeEgzYFzA+vQTm
vBuMEJvmnC5eFnOMgkUAUBgbTOwzN7veEWa0x5Eg6lNWJ3xdOrHePft9Rnvj
eTwQFMwH2AgzR5K7Zb5qc+l7EZKIQE0Cf+xfdRECfcLGnhVux+cyZWeSGLOD
7zxqHSxZXRlVxxCCwCNYJBr74Fs7g2Y46Sgl5O6djdmhRwVIPVO70qQLt27g
n5hEIvx0WnaM4i3lh/2WNRQSMYLemVRwOU+5zBdOWH0wc7tfWjtgcK5LjOYI
6bPTWZLLvPVCVBHvKUjOqx8oO3X+S+gpdgja0B6o0CKigUsDHNJtaMbhbs7u
RlU3JKf4upOR8s6TQrKhcAwgzEGnnc2sKhTvY9EkEwb96iuY0gyGkbohhQ/4
abu+ku2A7KNd/NPwjFbseAyd/QqykdwTBXAiJj9SWCT6eLTrnbK/rLE7zmWy
96+Yr66SzMLshIX1M/gM6Kp56I0epDVmmCh08oCQBgJre7tYAIw3Hz9/z/J5
+zIMtnzmKV4LBJlGL471yjURQNQ0Skti3YAq4omPizfKCDKKb67kV4v2tuD4
XhEoqhNw2WBlCun+1hC1Ff5jvKfPOs24qMzGoh1rRBRxkkPedWvVapM5bux+
jd8rgTDE08bvWRqW2pEQ2Ftc3FPOdQ2k0qfI9+fAppqfKsaEmEwT9okO/z0d
Xip9ibwufH7PF9UDMA4yXqkLK3pJf4DSSqgkr6CFlAxc4WPgs3D2G/aZydxC
jNKjO2uqQ4lhDH5bfQu1q8M/12iBMiI/3soFWtha0emqbX8JBJDTdEMVzkrT
3vxl0d7ABfh+VGVQC+fWQn2NkX5LxK9SKMr1NDucbQ/YE9oEKDUhwab7cYKt
APqbktbbeoBVLlE3dL2VBxEsdKRIsu6oC/OjzAFwO1jBrAHYABLq+yzyuWBJ
sDFQvSUoKie57cKYR5Bw5mD9rE2ZegNXkeYDq1UCeqVze+GsagU/pHmwCEhJ
9xjrplI4qLrSvjGEu49Ti7PdVqIt2FrIuTqfm8LnHGZZ3qzAk4KK4Xl1UiLA
t44y4ecpBbPdEJKMezQ9EYNTfjf/e2kgpetSSHYJUNN5UrPbW3ztr+vrOLLM
VX/C+6sS/s/TRh+qP7u+ZUwNwSez78sQnG9J++pTFxg8oKsDtJiD0l81IUYV
EdbxvJ9SjjaG6363CfrOrANXsYq9qQ7mnVBntPgfR8CjNrEl5fvmbgjKGehI
US4xZkW+hBxDSNl8QuBv9ZbgyDgcDbwkvPZ8oFSQLrkVClK5KP3tJYXTx5Zs
jTYCTz7enq/9nXr+w+Cho4j9mvrPPI1zI88KKc0GEkf19zM/yJyV+zbxgYUc
sw53U991CNJsnJPUOeya8+WkKiy4/IAGdglF3ebovVirRVm4tWHnpJGln5r6
wCqEqaBJMyxRi6t8q5cqSHHACPmXBcRdp4nn1/ZJc7KruTh+ojrjtJFHVN1n
SiicP0eH5YmS0kt2nUwgRAMkuZw6gs/+dc25nXKEXMW4VFaPJbLTAhSkuwQq
MuSa4cHdHyeYtsopEeyBVqLxW9PNGJilvfFIjo/8bwJEBM3WFhUbPn8ODlYO
vBYxzcmNWPc/V56/qdEbfAcnoUiiskxHqqATLm0odPtvecmoRNdBNi1sdI/Q
NKcvoMWOdzhOtRHNvbBrR9bsXSv8DoOM5FD2EfIMIfs9lAg7c11GbHXb32sy
I3ryDJqPcrIaHOXwV7pZ2d1e9iPIEXHUN08UH7wS0vf2D+WoZhmjLQ5Q1xyD
okrHZE5SwsesGl9OW6mmX/RzGGMgPupmpCloTwtBKHMTrdA7gW50eeERHGWP
a869lPz7eTbdhvpMZ8zXDoxW9DJgdMz6bNxYuZQ/qvbiwgDIYKdF3bjB8rHw
y68/5Wsxvm1WiFz15Cbad6Mql7kxh8Vet3D6GyZkDUzEPqGycEBGRdSzTJoE
TjHKIRpTM1gsyovfzdcSZ/UOLebBxYCAqsKWEP275JbDWUy3DcOEg9HLpxkF
fsTWUfyW4zSJR7O//XKhGNwtqiDgAPr01P+lIGW83GXFw5JFMAn+7XSDmGfa
z/FF0m0a/hpwRGr+XxTFbY7U94t8CAX/GXOmplg/wfMe9VHeRsbm17rO5+9w
dy9U1zc3/5ugogGGyVrofpevcJmM5QH47huU38uz8fcz4vuPVZRyvWsaRfPY
4XXuhwauatHfjHxlRQ7Ll28AHHLZEBU5sKaTc8b8xgvE8wIstcWdNdk8OvL4
LYZmb8x5/l4xAlpXPF7BvdjXeFny1T8Weu0RCw5Om9pv6p26lhL+x7v73/tk
k2OcksnXIYv4KsbrQIW+dtRMPrthJu0En2rQDcc4JPAMc+8zL99wgvbCSXpT
cCU5cbJ7dNHVVIf07d2UGCdB/RLHmU1eRARTXkVv0lk++VhXQQho2GAbQumv
48k0K6zY//pejuLkYgp4RBnEi145CN/KE0yA2dqf5COAEhm5n2bei5/puanz
gyXmye7oUwurc32DZnh5Us3FaDjCMAfIKPKVlPuRkBH4kGsSWHMxcPxdUd3Z
HQfP5ciVNMc4tozcp8qDOC45u+UrAY5bNN2LVQSrNd+qDfO+U+9Q06km7kWp
coAcQ4pmXAgWVf43olCzSaIgJLZLe+/mD8YA2OpwMI0DV/2qTIWO+G2ixc52
KNTZnhvj8CYnqy9ACWhxxbqh7doNKnubaaoeA/DtKdIly+VmT/0fa5KceMbv
cdhOtd70UJ1sCJtQlUmGLJfWzCuufpuP5d7k5T5/cWqBR3rSjwx0ntjFIt9v
6vft5yGqW2X/wBUXBbkUVnNCDHyKqOU4Ag6/87Ga/s4B9w+6jBLcL8YkDyk+
FBebpGtLAvQ5lguLidrfRYl+XNcIBcxJMoVqYOFWjIn9XNr/jdIwhioKK6v6
Fw3H2J9kk4DqlE7LCYo5C+Ez42xO0FHNa5M1qgGrFZjYCsWFXtSWq6qwtDYf
qP95Xc0HfAW2LjFNPkDxYqxJ6d4xJj8MsbamOpSXlv/gl7QkqGBuueNIBCO4
o5daoplbdM+WcwHA+7VMCZRIcHUMpfguvNksrpFvPrSeBpWzDUNRGXGgbC9G
g1XsBnhcH6ZEdxz6DLAc4+4EbbY+Veq96GGLIZgtsVnOF3sTAZH3Y0VqMDqO
Oc3QjPxeCYm6r79ZGaVBbK61tNxlCMZDvEzXcvejzyrxwHglBDOWPFZ8unkG
WRKYIJO09DMZkhXIVvxEmEaqV4du/G0Y0APHMs7P+KmghuAR9dzy4HCvHcNN
OXxKGF8E+7nnfUbBsny9VqsrYF7e0QjfvUYJOYdv+Hz0x4n8GDv4wtlkraco
R+SjuqtMM52k8rMdMZAp1ci2rhMClLNhOJ0J4MToM9GkkijNRNQurIw8xftj
y8S49utdakA8g7jcnA4X8t61sH+Gz5bA+wsRYxCJNq73f9nKNvWOFaTOyX03
pXPPhsgOHgcl561K0EKry8RgcWnFejUbSDvIyYN2P8R7PpO48K4/MoaUooZq
U2bizmspjl9bpKRpOBv8P1k0NFItxGB54v0PF8ZmdiWEWSBSzZGEH92Hueow
bPlof5OEGS7GjTM951ZU47s2dPSnM0oyvxCSY1JoI+3Hl/ge9Jk6ZMl8cRuP
/NMsnipPVGYMy1Aex5gWXFM86P9gdj3iCwX/VcbeRMGW3EbVeLKwS04VfWwl
WzvgcC6+Nj5y+9Ef/5FO1F14pJeS7A6AzMl/9vBMkfDefK83Vmd/+kf62OVp
QzAkU/32hGqd+v+b58YvCLHlH3cPn6vCalYvInY1l8wp0paUYdYt6Uk/LKPq
9vh7Smg5WTvgx7/GGV0fcP80XGHne1YqZZBbZCmmVw8amiYhDypwLeR75hca
oPNazI2udl3G1jlBmhVKnvZ3Db74deALEpC4f1CtZbzVxdCtRv/fJBFedloA
D70BNBJ/G3bQJTkaDPwk+IgFhcw9d6Ft+aKdGuRyST7kR83uiFrJ3dHtn1X4
MisXKG61edBmIm7YUZTTNe895PrZFheK96OPQP83R3HgW3aqd6ECsRAHYatY
m8aHJBuLa3YseXuKAXLRJJ2Fa2CQGCAKGgQFgV945AbpUlm2SWWdsdq+khOF
l7RtYuXCJRIayxAdqzfXR1bzhS+iNU5CAqEHlD3sDjlKAJmfGzVLsk8bz4PR
HqVtFJxa2Ev5dAAknupah5JZJ0QFAXMryPwJLbunNTbL5eDp1v9sxVU3yFUu
aZIVQmwsg3+EKxd5Mjqd+s8VAxapIRVxIxkIfEDGwRlNggbpeZRAT4m0rtup
QZPJomd6VUa0C+iBjqen3PswGaUVsGMAlIn9/DWd/S+sgGFnCq1Ij4v0TeNF
rMeyy/UPuk9gjw6CYqNiUG8Shfm8AdPaX4arAfu/lTklSg8EbPk8pbeh2aQe
+0h2c4exNxC+jBCakOidLqnkpGAU+HYFH5/8Bz+h7dAAmuirINDqX0fUyOoN
IsTiNW2j1NRoCRYk4di8cwVJ7+yyxnkhBfqWq38y3T+lw0+RAOSO5XQKlexe
WR6sDfoN7nz0IQ/yenlH/5aIkT1BdOLouXogBfh36OchkgHGIcW8yoHnAmAk
oEddo35wWMpY8Amya77oVNk8XPJgfbLISpprbOgTw3Pgg1yL6z3yWkPvCE5z
ciAUV43I5LTuqeo+FlzRViUa8OzL6t8jBYGeJErUtmvXf7IpH7uxYolAM2R+
MfXiHpxodURWXMY49b72Oi1u3N00DNWx6gBWSDbqeRduxL0rI2NV+N5fqIOE
S83djd3nGglTqy4COzUugJ+41uNSWVMmrtY3cPDp3It+1FM6UDTTh2xpyMO/
vLNzyRO23CQyU9qmS11mGMyjjxEU9wODDzsXkhMlbz7N8i4VJQnTW4ehxqQz
IKyCNFbJoO0fgqmOzej/af6440INnC8kgMU230rbzmViK/glIoIMqFBZiUBT
t+JDjigVO/SiOB5VtNW1LJMoZ3G+LlqfxydUCss+BIVeLyJFL/vmWfIwM87w
yW6XKB4zCSigCESPXQXZBKncXnFtf7a9OEyrW7d0noGNrNeQSNhAn96Sj8qg
XuSpEZ25uxIDZ04JdjHlPwFrfmEC+m6lL37VnIUtv4xbimyAVqQzFbUuzWrg
hWB1zKX+jKNy3uXeAsrRNExORXrmrFZ4/2ZAD6H+fB3vP1/IQiGoJJWHkI+c
aZYH8Zrg2rnlBMvtv5mmotoehx+oYbZGs+F08LIawRyDpA9RBDHu45TFmPPP
O2h7hVbMDNTIIESoKHMHjqtMCQtU/RN7IWVwX0QK1TEo7sVk64y1DrXJ2h9h
jMGg0Ma2nQrzS/35iaLSjn9H2nypBkAU1HsCVJk75FkdIljDhCCKJulVb1SI
RxkvuleqwI5+k/f4CSsRD96g7JLdr0ZYBhXC8+V8tpraSUfA/8j8fPFiF7yu
dBYNN1w7K5gZ9GdHBoUWP+1lJUFpAJ5zpZ6C6kP0SkOFHbASCLgOFbj+WiA4
jeW2TpWrw8vUH+YBY66WQrkdm2dsb/D/XzR+up4Fq4nzEXMmSOuVfeNcCUjY
OG+rvLJohOLeu+G/uB+Hk+QYETsiis4x3ShkdJ+fW5ACE9hbhScuO9i0jBtU
Rs1rzxAAUQqtDxfTGk853TNjP/ost4qcFoy5H262FydMq8i1A11X55MSxo5T
MVr37bia8gcBwDOuYodZ1P5jpbVigg2GwG+CCw4oBADmCpOhSawPxresFqAj
AwKV0vS5IkmiTQoUoMZ52dNYKPvnzBSskzSlLpz6eInbKkY4x/j5owS0sChq
z09H0VAkwmUXYfb7eum/iZ0Qi/XemgRti1scpNBjf+Qiy5iv2Py0R5lSOosp
b8P0FbC3NH08bBiTRkwuZ+oPyKAh8ThYAEKDU1i8nUzxA8WLgvj16poejTU2
dQBLomaw2ciX3/OtqO4qNxaCWTtiOpg0VkPe+OrMCrVbfuH31GhqW6hLjK6j
jVaRq9e4cm1V8Ye+P0NmoAfNRHn7oIEM39w58fWNHbW6zdF7qZWLWJQYqEp+
m29JCmQUvDhHwz58nylT1U6d2LNa8zTYNMMHmEa6j0w9UG4j7wUwWfOBCzv2
Z+OTp+H5sucAnYeYsVqUmvq6pgj9bbCWiAxplWqAnDa4WlpHTxLfUUVtvpZC
vLi+SM5C4tiz/YbyJ4u4S3xOPb8sCdo886LcPIjB5RjPKggjZAh7GjJlKizG
XQmn5Fy/u4ek/+SN730Oa6V0OTwTKJ84eyM0UOVIGwTcXgX2rbQUexROLSIS
lSlQRlhOP6ISa+Ezgs+5GQeqZqzBo0Mu3IRjQ/fQKPR2/JLzF0QSVSgGlvcn
nuwZ+3xqxJ1FCcW+Kn3WBqxhWddCJX5wdMoplFefu2SYl94sPTScXdfwvSoW
Jg0PTEG9Nx2rPwlzL+abhGzBab4hVIEL4aOUifATEb1Wk4TGPlT77WJdLAAi
juyE8+Tk+tS8wvP3F24+nhstaTCMNagH3KlQP5JOjUlz1WiHaz8sFmlgrZ4O
zu3qq4Qh/Cfmfy5cbahn+1K0ltYFcn8hXjd0eC2xyU5o5kbw5RmeqAMyXSh8
1cmUrZl6RaWHAFd2ZSBZhHoLmJ3DBR6MN9v5BhFlYCfjuRD9qz1Oh0t4hkKZ
mzeVESsiBl63Olzg/uRHteJFV23C7wZWyKDcjkcb8sdYHGfmn6FHASbIC0sH
YAUwOBshIJokXaFYxOfU8xGylLNpmoeV07aPLEwiEpsDK1NrqJUMIIZrxb3t
wSP1nFA/53EE5lS9nT/gTQxcXT/PDaHndd1g2dbgsVUTT9RLBjrQLDZtV8ba
786X/JFIqS5CU1YQuBwCtjH+03HJV+lHlTE4ZwROYMDmTM125D2f5eTxtUvS
Y2L7pFc722r6xnxu+ITTY/4h4cTV0b7i/2FNBX+qnG3RuMAmew/20VtgkPts
b1Lpo52k9TpobqPnPiLtdHKLfKXFsXq7sbyb4qQQGKlXODERiElOdVSHbOXr
phNVroSqNM2rDP2IpaFFDTExrOBrzXLVz86c0wnf+vF32hzjwGbTkYqvG96R
tYP6JtppSeAQsIBuOWcPXGtZyExT7o70qxEqfZKtiRdJrAeO2krrWbPntDPO
HCwY9fVdoyIU5QKI4aM6tCVkRJcz3iw4wrhqimR7vCcYD8YeM9b7tkMx87FJ
4m64819GDsvTr/dc7pS5Igg4iA8GAMUzZm3PY3XAsyIQlsiOE3OU2uWDr9Wo
Dsi8k5+84BntMWC3HDcxpvz0U0Xo01F7Kk/aYXXO6iuXjupdUwE1auLGp+Vw
7H0i7ci3b9qojN2SpypAn0z6QpDBq5Xafj61pbROE8OCsGNua4gXncLUpdn4
YNSVwlTIIMBHKz7V1XsxbBOyVWISUYazUnxYftFoevRYG2uxBmqbvQjC1rrO
GKtOSQ8kV6wMbz9uQpj0lz7KEFscWDhC8jpRJrx/jxkXecOlJbJnKLasgPLS
B5wIyOgrrNOYv7jPz+nXMGwHoQSbIzMunbDnCPfkxzxqNMMS7WT40F5rM2QC
HM9YrD5oHC8pTHwCHKxNLFmRfGeT1W1HJmyQijV2yyBlfrWkWpHrjcBrWb0C
DAbVfbe/jQ2vDXaypPj1y5dlfE5n2TRGeaud2tMVjSbCaIjEl0xhuOE+jzyl
ri+LbxfAXNZyEzAaNjIkSslBfrBGstTLb5LmnOxExx66DC81bAKCJnD1IGnP
NIIDuQN4NnTo6gPetFgpbJxu3Pp2gwONGAAcs+R2+PXS5Z5yPROTyZ4FyMVa
jM3hKz6RrHXEcTJZ+ZVnkp8ZtUt9ibp6Z1skbVbaupFaywCs/npZUVyZjIz3
abbm4nnIh8E7ihOzCrq8wvq6gAi6Z7zONtKOjCRYwrgKae5z+txsF/Ya2JXa
us/4HB6NGURKhcJ+6lmt+cifoVCWkO6IlMZrutNd9IwsQZPKLI64hLh2skil
JQWg9OjenE0htfHWQO+3ERwAYrRDQ/sm2yrl2/ZEO8/ODGHUWxQL268w8MRr
+5X52WG5GbDPG+G1Sjf0tsX5Be7ydU8fRKZaFHiaTyz90CtohvnBvkjhouf8
nMgO2vTSYyRExiz70OAvjJUz3Em4KUauB5g49eOz8kCGNcVPFQoYZPXpORNw
4UmoHmCTVj6+hKHo5ps9QMy92DNNDn4ElkKlUUBwEvb6pJpIYqohN2+3b56b
IT72NlmBM/O6y1hT02V6hLi1q/eUoKGQeOjfMbmKDsFFyFyB9khHqC8H335w
i9K9hceDNyDfv3A9U2VI83gC7xcxU7bjLn7qadXWhM5Fu5KgRMJokRbQfpkn
0kknuAEP02PRWpWaNo7okM8aObSVgGJHcnD68+AJ4/FGwdLV4DgxUGCy9Udx
PE1XdDJ+w4H3tXRB9/zcB43gerHD5F5tIa1cQ9QMEdqVVMYeCUCx2AKwhnyn
lugTY+L4S0niG9pBVUdtJ7k9qgXlahKFM4cwaLFIfseAOnKM9NcSIzeODTCy
rZjggUkfG4pB47diTH/WzHya8z9wxjb2MHC8y2KaJjjNCPqRgw0Vx01hzQj5
q2b6yANfx5PxTvNgQkSmHCO+P1UCZSG5xPrBQxUnqP31VQQsBrobcMoOTdWk
7doXQk62mEe86GsB3x8j72QFpiAUaeclM2TzRmPQOTzKj5SRrQUP6gS3E31K
w6ZqJPDGvjEcz66OpXGJ2Y7ZCigu3jJKJGFPHWiZS1LGMKmKx47e6y+H+I23
qpnNLU6EEkO8R5OL5IKTpCnxZr5i4+pN7DZD/mI/jsKtVca0P1SQujP6Wy4L
f9ixHbzaYhqJMqh0791ftEahlabe+mlEAm1QZTol1RjPOdGG+uGBEY/UtvOI
3NfP0pr8M02h2rDo6sOEouYL1P6DV5zlkKcbKEi7cvQvcoNKKC8A3ESjfn1q
uK1OISd8Ju1MM2iNC+vBsdJALxv2yE9zV9nqlSSxLg0pX0Eu1gqENSwjhlu2
X0CHEduIvdgJUIjB00Rqybpl7YYnq/AeRInFmC7d9fs1awX0Me5PIz8fgGaO
9Fhw0U5M8hOHqC8vptyccV9DkT/I/Ss/ZjRs17rkSm2hP1zoRjTPy9EqlFLP
2CSy/eqQnvlL5C0U5O5pAmxbIIKBk2tT5u5ETZqwGezyPPpmiFC6MWyy1HXC
lP1H1xE+2JPPGSQaHXXA/6vpwaVWOFO3yPdD7dRkre9aREnwGDbfw1ZJjUDt
L/+hKUFS8Xytb3ZDA0vV5D5cVIYIVrYxLPr3jttqz0JdgOBQmW58eocqL2a9
A6AXP+P2CVhPMLg+8pYMvilEsUrTs8Imil1j5wSXHaummqB3fkKPE3cKl3AD
8gxDSgFuov/mX5MFybVZoMqUWL+iLIJtGPhrX2nb3aAhW2+LucP6+CTYndX4
ylz9U8RXHbyTPf6jzq4/KSX1JevuNc/i+Q+dyKpq8/7BoxOcdd17s9NeCPmF
dNlltgfmYivq8jXcVQJxGlhNgAMq0VHS3Kj+Uq3CrlcFEdw3Odt7o3y673yO
LT4pjAQlhEqNILY+1ugrf7TDUuUviEiB1oDWU8+HzjVWspvkSdY0hZi5gicl
y+gOsSHsX/lcFc/NnoQ9k3oRhkvOFrxm8ct0GlldMuORRwyCWnsqcUI4G57e
JRA1KmvTcD+cbBaMctutXY/N3sRIenak4tqetVR/f0mdLADqqnuSXsB1gX72
HfhRlX5swsgNUQHPtRevTYUB6vXHmoX0+NKtpG2n61yB7lzgy6rqlC/QbFyU
ciDLhpjh5gPcPH9qKIx6CGM1yHXAe+O0ymdCJvIif4m/1zUOIKgUuXGZdaUd
pmsrfkXeVrT7dkek4Ai23U3KKxez9Vk8wdwIBcHD9555i0YeF36vu5sE0C6S
/dWWJ+Pymnbg6bdoRM5fYcLdaiY5C6BSLmVUZqTVqI8q3seWtpdDrbbpON0q
Cpor2k3yyWgz0o0XqReo69SzI7GyxJcyOiNh1NJ/Uw8nqaEu2jNANfWNP88n
tLtSfPVCLk/SfIDpC2wUO/bhIYRnS3TeCBXOsMOYbib1FHbPHBpvrd9vtisS
aa9kA1EWZcZGM/tFENDvui2nGjRLIO9MrFz73w0GtlrcmJVVLOZjdlx6iDn8
jtrvCoZYQVT391d/Py2S8BCSA6pF/n0+dXPafT45+wcImXFLvqhf2UwQjeWo
09JIj1hUW4ZCiTB1F52TjGNLUJyioOHAug4UPb3NeO+tg4hyUCpXPx6THhwX
jdJcGihany0J6PnktWrQvpHedS4x+JxJXUvUY05sxIKKVO5mYdcQ0Yfd2mKD
sJZIuryf6kv81q7xhjcfLffKGi6EcsRUF5b9BYdlULrMdom5M3R9j/8MNufO
z7VXOO1kWnl/ofPlGBH3e3ER4Afmb8VIANg7i9Y7KzebV/9wplKAYbeu9qnu
Os0scsBp/obw3qFBpbu/SiD6mvCLdcihkXs+tWdxQjjXlBBBdUb/pQQumjnR
gVvY1fTYCXnJKoC4K0kiKK4blseXZ9g0sl0jn9pXWjQYJz/fRZSjF5K1AhLb
wgYtViQsv9wruCe5kMt8vjpmZ5vaiy7k3FQhVs5BZzbkA50Rkbofry3l9lyj
ucpncwo797c0t5xTjOwlsTyR614MYKooRv+yTrOzRQyssAM1iM6TMAfq7elE
Rko08WRFT8ptwhQRyA8/Du+F4SvK/hMuIwV9d6hRDX12M4m/bBD+wsRcnENs
sJh/bgKVeH6NFDcpuvs7jQM9ZRLF/CEVe+CuoKBUoHQzJD+oQOk0SBr8g19+
nusw2TLn7XzFHgkTh4eSQa3WZvSnUlrXnHc/DigP9R5zkCAFdYKuEolSjbcg
oX6EZ0iKbgHwEbSq444ixTfv7+gqRaHq6yDbnAXTgPzDdUljXlQDbb/cJN3T
9djza6Zt/a9YLGBo286fnHKhenxPcXzazttYx/+nJcfXUe5VKFlPJ3qj2xBh
3MxEYymQuNa0t0oKBVhm/jJj8it/PMRWOp/TjBPiniCbVJCu2hJRMuwmaLe8
KCVtDVAmM5wHxQ/homRUBVYaHLiCw+6ZoC9BMMXNeH/RTziawP29WBygx1Iz
xw4tnV3v6dWXoTAIazfHt5jTMhiF9ZvWH33GVwRs2w8q0axSZyV8E9i7Hndz
GJWICh7NDSKxfYk68mBxLEbChr7lou/ea9zGwlvHIDb3GbFCEoE2CYptAfkl
kuYyI6o5MxIBZOSqavue9XPmd/cwoDmbwKJURxUiuW602dwErPlAzXpTsp4W
zdrIhgWQi0rxNwKpOo80Dj0pGtV9e0OOWViQi78jiwufssaiKw4UNjm2XBK8
+noTHh2YtIC/02FUixwHQYh/rW8KjOkPevByUGporLoQfo0PgxLZnaWaPnAF
u/wXSiE9/cr3ujJrAzcPwzvll7QWcVq4wYTne78Dcr6I55uPHHPWSdQQB3+E
brthXJ7xqmEobiXcNpkW+FtnKl1qbqM+MZO0RU9BTWAbul2MLLH9tNnHUBfh
XKShlOxGu+lwdohRHwTmenS+pvEytFyG9beYIuWFjA5QOvgdaNqlxDGxFOFJ
91r7cW8Q6UVZ5JMrCwI/a+EUE/zbKmjGfdww42imkU4toIiqNpHgzUY+kJHF
Yy5JvuTtjRdQYtWYNjmlsN++zmDljPCNKDM3YLuqGGfENyn0qTgJUvAADSKL
l0+o2GxgM0Djq4Lw7R3jdF2JgjQm+GDa13DETpj5hfNbORmmD9xvHMGcqe+d
i2tulYoR8uKdJNoS2syEBh+867Mb01pYgi0oz7D1sWWDAya+a3+hpoB1rS9s
OlLEaRKgHksSHFn2CLQjRhEuvUO3jNbW1+ra8qSZDZDs77nYmczKHlgTE0RE
mhUV8uQfVRvyIHKPcrrHx4W5ED9KaX8GVydKkWHv67R5n0OKqL+JpQfTo/i6
YZLgpRp2lot7Zxv8tuSOhmpkr+QvnVRXqSRQEVN+7l3bQVMPElc0oI67n4N5
HQOCiVtERO2K5O8j7ZpE18Lwu/X6m1agZuTh2cU9JbXSS2aN4yWKpvt/HV+k
3RiCCfLK+BneVmDEPM9pbMcwKDTaFUBl9mfZKnq0QQRrYoAdoWAEgExINJrP
EIY6bd5ff+HkUzxQwilFS6azYWMyxizdQZFsu3zqDDD0VHhOh20MZSHwaHnV
QmDg8sP37WNEahdS0b/4WZQVCo9BZ4bG64xyNWqejYwL9c6bpWXrjcbNNNdX
lzGWIl3Wnemb5OV+1w01z7NSLbcFmD6/puYFU94Uk8KfXtoEQIqD8vUqWxpA
p0H7gT9jzQxIgUmizqefm/bLfpUTD6pTJNHlLJ9xtIDrHcL8gaEwDNhZznmh
f7MxGr3gNRso7pIgtbSl0QYbCNXzATPVytx9e9A0GeF3xw3BUzNW4v+hUdVF
XCElszN1+CJfrj/vexl4GzJ+NeTk/wKGc0b80eP1+mVLD5ih/ydjLRj1QzZM
+iDkgCqJ6LAJDTOY6fGUPSSdDz4RWh+PzAgCCmlGkzotzX3JbE4CqvW9SJJ6
37BaEOKAklRzGocm4KFpIu+Z1BBXvm2FfkwZvmLgWNh77KGJfyx5JXOn6qhZ
3cyMiqVHi4sQnq/e99bLDTekG8myFP2wPYk19WcwAvDCN62V0KXd+1UgTlxy
lAoSCgDzfTQR2kHFSk64dMk//R4LSxW92L8QFgGpumfuZmZCZbgnfbjOL7oQ
Gnx2gjAgnKG47FnHe8YdD6jJwN/0KEN9UPQs7o8/Gs0HvLFq/WYLj4/k2Cte
aXY//VERTM9TCpiwd42Uo2rEcLFwxiO8r8EHnbxSvtTcnhavC1Uy9RfzIMEx
irGYBb/PXw4K3+4OyJvmnz35OozTf8tdK9WAsSUDDHJvRuFU/V4u183ersLv
o3Ms8uAcuGBNmtNtGH9y5KjvGs9isxVnOAbAo8RN5byrgHo0abdan4JoBWo8
EeSr6ddhG3rwqNzjhxoqEoMK4SXkseE38c6Wkh/SQAWq86sm0f1Ve6jjoFYv
Ipc9tXWF9Gq3EYsVEIHkKJsDTq8oL92L3fHsN7TRYyQRr8S3MLhtU2JPXzd2
2h7TCQen4vqdiuh3T8xCz3MJc2vOj1sznmp6xKOyoS4UuxjHqGAcVDYe9KIa
1J6C+BEoEHz043RMO15ZniBxDAmREUQcIRymOKEW2pWPC35by0jLNn90qmlV
gHs21lipwc0cJeHyFFfpwBRcIrH0FMhmy+VJLgUuJFkSbqov3RZ+gnYrVBzC
UbXrwb4KX/sntwIOYYhZaJm374Oe2LbVNoE7ES8PSkCbpaMDJopTnKkEZRD+
tlP09MIivwATsvFaht/2lJhZf3UWxWpvVm6uQfh6aZuonLGctQaN0YWdGJus
Bo8WejyCMf43V+MD7SrJV4ha+Z6Ciokp0wm+/f5CRM0/jlxeph8t6VUXGRzr
3JNjmsjm51E0wFV3lIDf2RH+MPVkdjWm3GC/lBrysOVe0r4qqHijvOGOeNY7
evO+lqmxFE/3RT/JOWJADQiNFdYtdOrTCuvrr6or8ZKdMWs1nC9womvI/RKl
Yl4M8D605ueI1lE/iZr6+RQv0RhS5lQvHJ5Hi++A5EMDI+hbAG1JACeLCoO6
22jM92tkTRcUzp6hM1hf9758h56SEIOi+J0ynfP81ApA+eI09LOaO+X/3QZ3
u/K5i0MLcujOUl9aZPqv0KgtHbwTHGcGDgdOMNdZ06rRDlqyiCSwU9zBf/JI
ZFEufgPoEgsQWGCap7R8tAxSS2JE+eY8s+bCoLYzvvIAZj2MLWu9HxZ948Fr
0jHCUacArJtFH/bLzzv6Vy7LgSGFroHLxPT7sCVfIHqTJYWYoSTtczKEb4cA
OM8QH6esni8tvaltsrzX276TiU0MkJX7lJ80sB8rhiO9ezSEhKJ4RDFcZqD6
fqqy/+lZTTfP1ZwCNoBrLtt7A3Ng8G0SEHoW5HxP3enqAYwTBEERo2gKBJ+M
ZM4o0Ex97509JS40bd3N87JpMNzEJqIECpW9t/Ma0A7ixmv9pmH9/MKF04lx
l1oLphRm5xQ5Ydf8vwfljnCQQE3KUPXdynT/vG6m0zf3WOjMv8VsiBweGUsV
VTTzdjlksDJeNwpSytK/xljhuISnR3atSoVcbmP0IM0KRvAJhcQD5o2OXlkq
JlT5HvrC5akugoDdiRYc1ZG8ysEHK6Jp5R1VuddSa/w62jPw/b/xfuKrcYby
wWoEyEePNjBONCNetwMlxqjtPhFXcPsLc/73tOwRHmav0fQVN7665I7sDGFF
D0Z0f/QfSIKT/+nFduTKw01v2Nkx2v89INNCEoLmIkwL06G3rJxzRfcItMeH
Fv9FZaq7650btKt8Sof6Ui1YK2H+Jbp4XkqwFaAK97ljKOWrqh5Owg2I89/h
HdRwNQPUwwIvb/DtpqAIW9RKLCH+0r/AMR/VmlJo4mIJUPh/EbXM7Qxkg+D/
AGt0SxpBUwZPF994vMVJ/lkUqiSagkaJt9nWjBr7LX53cGU3jSX5foDcduAk
rcDxCctpnblEwqR0ECTNsw82jnfo6rpCda41sP2/OjpUhntGibV5LJY88KdB
J1PE5bD9QVTOG7Y2+eKsIQpFVzTybiqEgCRC7E0aenco5hJeB2L68i1nCPDg
rynB3Rf6zbViNFbCqUzKsYNnuDy3SijDATA9TFW6SCyYWMs3sLioIbDZtYAM
IcCSLvUTy55z61s/MPimwCmU0tjDY4ry8UaPzvV85/el19RHn1WHTvNDEBQ0
PO5ngiPRlZiHwufj9w2JMUvdUaW/sdxxRO+B3ZeMjUDaj1l2pVQe7AC9Lg4T
zM88ScIEAoIV4PAJ+Sat1ZsjOvv2tFo3K3GdRk6EUW2suv7MscHOFGwN3GUU
IVzXZ8Vjp20MjfVGW9ReKTiZbEgGCLY0Zah7YfYcvMhvdan32XuxGVBUhyNa
PcNJgkYygW0FRWVs5/+tjPbY0nV2O6pMCN0smM3n7wALz7kko1hvExa7RQy0
svoIew1xuzFVjjIMBmBY13IzQ15qMpZDm/p+tjXML+TNcOV6SfegZJ6MBgIF
0HT8UWwmnk3+VDMBFHFNG10bwIReFRJrj9r4KoUipo6+QW1Qoe7rRmaCvKjo
Pwk0bHwpqtN4UyMKEM7Wv2dFlCt4vlqBm+7jDj4RACIKmnKElQN6L2w8JL5p
HBb4rApGjCxtKCG/DbBZ63d1yeOXPSI03oMnUN+z+Ia647GP9MVxlJiO3V9N
bWIUG9vatl1DXCczH/9XREcUKbtZc3IuVeFGiZiJbY5QIoVdgSyFEzFJbCd+
PT0RUKqeAYbKjepv7oRoh8nfsmJ7KQldoR0vezos8cYYYdYrJnDBX9rDrTDj
VwtB/T//8xc3VC9vRG6oLa2tMA3j4yvATZA7r9myQb4aE4JsYzopklGdRSRU
7omDqOCuL6v9xMKlSBClMFtjcYMQpI/ZYvtdYhXQO8SGs+PDr9rUwImtnmvD
dOwwbWkN9/toe+59kvpL+mA6ifAp9GUi0w2zmFkW3Uro7bvjI3AGpWZTfqp1
dHzOMezdLxFAUFjkhe2KsNr8nhtfrcLoQzLbDp8Au0fgelnBHrTCIvEQbbNB
28IvDFU4qv/JdRDyyFkQpfkL/k7d2HMiMA8y1LwETr7lWObTI5465mVNgDNk
kN1Y9+ppNJtBdcudIa+NhdRxkYcRGaRofcR1qV01ddSvyPUYFYcJQKcQBkKy
PlfraCxK8SA1cJEN32nKtOX79cYtSQl2w+lrp3X4HffYPz0nzl5cZg1Bqynj
3w+o2S02BLhq1VKvX1F+TveVFppMhx2VfAJrCQ6uqoYmQwQWZnONez1Gt0wn
N5oNpgerKyJtupGXj44GtzGYY7+jU2ZeAaAHx4um1J4mSvcC33P+S+60wL+Y
Q9L25T0nji99CrnXslp1Kx9zfVlRf+NpTqH/uEv2cCPGVpolR8jKL12M/Xo7
BCfmovI4QYZ3Lhe5gVyt6MS8ovORI30SnfXq1VT02D+AxZfWyeE/7pTyvXId
dkDiP80kxG8zTZuIh44ly/rmT/SWZqzLRrs4JUwsrwVcEtr+J6c0JHE6v6xa
l7uONUG5uj3y47Y0CaMQLXZNBYqNd8NfYd24P8cHgM/WyzmKgWeV+ytirmUv
lXmjJxE5Av4vaxT0Ml4zuc0wkrR/WndPKdz8oxawu9Q7iL11MKNRHoBAjiD3
qs12PJbN0l7ev2yFysmPcxZBW0vzeXfYYTKIyfW5srrP1E+Kmv4YvHnny+WB
TBz9djQiZIMAvZPvJsOIB3InC1kpyY30hzELEYoCfkYNhUnEj7URuPdCT6Aj
QNgdrfqboSoEvm6t6t+8DcOCW4Wok79eYo/8H0mvLlLHKRaErzpIZ68RSrPp
v7aWAtjCcGP1UIC6HMKcLnRAemNtPARGBtnuSH00nCqlLtUdSiknwBlrpBV7
pAtdgxSz5+Wwj2yPZJOQ8qQ7AP3VH7wM55ZSoTomrfBM/6Ab5bQ3GAGaQ4BB
bMOFDxhYoUpYLwKa9zS/DIT7VzthyVbkOuX+Wv05KGzlS5OSW98sN88yGf3e
HitdDCB31A6toMCNl0BaW896JKxJoPAwgxaSbbTB1uxIhJMPrVf0IPG+tGxF
8zuDxRMRtwflK9rEjIJP0XlCmyPzcjoGvDmm/hp4m0m9jBlZUPU83BY9nPl3
+vDldnDwlPS1j/jhj2Y4XXCrAze/z31oK4sw9v5dQUCKf5c5+G1/u4i3dzf+
+h62S/9r4dvMlCgali28Gjo2dZm206x5YxeCqKfFR+Szuni2vh1jzBeAtEFj
ahU95szP15O8SpUPeAV7MsthithOaY0Yk4eOcFsAL3Wyb2wboVskJ7co2OyW
qvyvOPQ/XUIjgkCI6T7rWj9DHShcq+Izq5guvq3rQcrMgy/PslVcC2XIJbrr
IM99iJRWRpcna+PPgznWztVaiTuzPZYleEtRvyihV9BjK7m0G1niUPatTMLd
SasgzOAjBJCsn2rNGQNoJ6EACA7Iv6woFZNBGpLGxrNLiN0U4npIeAbIsFaZ
Y+QwfR3uqhkLGyNsOo0l8K4SarHrUreYvEpnm2UJTSTLJlpmgKoMU1fIBP+c
LuFB5nKnOQy6yx1poEF+0G9qogjn+4Z8t26pkO4mk9lgrkNAlAnBt7ZYI+A3
L90IiCLd2G8lgT0oKBHKPHnwl6kAyTCPtyPGoG0c7sUOpgD+SPA8xJv2RQVC
f6ApytIRQQltbLig7nLgNREoO+SJSm4xbK3WPAiRcXyBhWJPNLG83sqRfzbZ
/LzPSyjDZA2GPTBRRemOMmkPVftuTagvPHQZWDChSJgnqrIO2W9DSRdkNJee
2ZjUfL/dcCEQKea1dh2I+FZp4d3PQKRCV2AggCp3Fvj4mEP6k/n4+0Dd+7WX
nATYXDLOpoI7Rk8hVPGHcfHxP4kqvavXH/7u05GQtDnY7Xh6qdCcdLqUuDsb
EJS9ksDG+ylI1KV3vrTbwcijG6Vpyb3URv++e3ncaarn0tO2a0fL1f8APcR/
rDcNg/FAept2Of9Ln9wpemRAFMtfpJUvXhphQIMA47VI1MwIZNAQo/lvIMsG
02V9+IfGcyJkGbDzK7XzFFLVsp0oSB0FJf7vtaaJCO4ho1a4V196s5P1eEVS
Z9P2Cp9XbguUdxWlOjFHYkRO3S9gcUEEv57DvzS5Aq/vEn5zcuQfmlfnbxOR
YABr3dc54iVghrb2HiGSn909aVxYk2+hSWi+VjN++zGUGq9bmg9aFqWRZYS2
kOsTGsizdgd8VynFia2w3IxO9F1mPB903YTOTptlbr2qaUkU3I2E83IL+jNF
NzRTJhALp0L16mTI6jQAIN01cSq4FVDjoTfOhCZPcGLjafNnEFpog/ZBkl5o
eWRhCCK9y03lqlpmZYe4hjCgniwM4RKApHdwEXQb09sL6V5O1fVhhp4KJBIe
sfU1VqZXqNDft8Jw8hkKbU4XwxEMVZCkmVLqYg7hJv9ArKvu9i4ehXGw/miW
CW3ahJOayXv8v3Pmil2lS+rhkz9rLWLeDcwPvQuqqTiPhGbNYAcePHNzF2O5
F0SgVlFTF3t9ULtU2UZpdwod3/foIztVCJOEmm4OWBXiRsbj9DHoddZdlBe0
1GPt/Ydi8pGjqvQSCEb/jDp5oVQcZJZpj749LfbMmuK1n4+LwfIXX41Q+cm4
+epCY6eSvxPHY3cSDB9iVhfUVxVfRm4tDJTflesL5di+aSxps7HTtQV2wsLi
8Zv8LGT9IyOtROcaL+Yqoxk53FqmDcBXH7gWGU118jwxtbkSg4a7URu+oQOR
S/PAWXhAhyREG2TPS+u2X1t/9I5pgwEzLX0a5R7rpo0euZB0sbu1GMRC+4LM
6ZCbfXIELcS+fpNWWhOz06i65dQBREvvUUVUX+JZMprDGWs2rwMJmKsblDpT
V0oFY/bLBK2rsi6Tudxx4HE4qKtVtbYHw1XqZYrc98AgjFpVpy0hzfd4MaEI
7qoXaEPGRRbkCvIZ+Gl+5jAuYGVn3vcxwTQW7Kr95dkEhRW2EMhqxnPsv4Q1
haxYDdltgBSKH29hbZ0XJyBuM61cs5CvDJ/jRlZTb6jnmOee5FTdp6GS5ii2
mJzmpkJlSHM5k24Om0lMth81NG48EzEOgdi8Ju9UROvzpFV6L1DzsaCO5MFw
w1YouOP4a/eUaEM84bogt3Eu80GQYvN00hXG1nmY6jH7W0oje35XQa6L08AE
6yApRxyyDeTKKf89HtgNP4AKlihsCWL2aKqbR0YSMm4LznvEisDCdruNeyc+
edip8A6VO/mBCs9Z2ZKkI9w8w1tvZ1slrhEWvV9v4LKlKxlYo9QBhJEXI5hp
s/YPVySPOPB3NEzQZnk6CpHsn9o4kzzuNdTwQX4G1PkjlM0BeLiNu1cVmnaX
5g2xGtMBqxU4op2xa7pZ/DRRummFroSAv0x6oa7dtUd7Ke0xbQ/uAbsnU4xh
IlxV/Hgs1YCmpAT5FFEbm2oTR/6XkGtcTGZrfj0k3k9qbv8FHFbDbhqE2MVU
nXaTXlszHEjGf46loq778XESS8EreemgrnTn4C5UQWVovEWabVep6v4CH5hF
KOJT2A1qbZdESvsl4XTPPs+XPpXuP9esBPRTdWDq1cN3V0Bde+CTSah5I5HI
e7FOcKND5/Q42KjFZIqqSl8LuAiqbrm47JhYqk831PLOpvtPzZUpqJ9gt7Tw
AiVRB93UHNyq0lE73MbG4LaMfy5ceTnMdlLpznAIkp+3J79mA/kQUYn77hG7
nG9cIERaL86dR6QXszFO3IIb5d4aZQSQnWaJRo4lVg3Lk85YHmiTVsMzp6PC
K9iQn8eKSNHXgfIY+CaFp7ipl0AgpDYx5m3blLHpk0Bfesigl02CkRYEhI3r
iSrney6JEc+nY8Dbucdz2SwTa6iRmySn/mDxPiiulZJwcaGhOX0M6rRzU77p
ZIt8iIzaj/1mc5cUiLu1AhpjE12t0c2YPoI9VTPFs7gT98hw8JGFS2WMKwJT
ZXzK9TOkyrCyN3QR2I/xHrj0BUe4ARS5H3/2iX1Rlz79oo87aFoKLNbOnTef
m8/wRSkQZ6iRNmbf878XjD9ZkNgh1lO2kP/o6QLGpB+PG4POa99SmakLpcRB
JDsKhVKpa4zoX+9WML/zd0yplI8QbfQvUBNBZGRkWxGJn4hTL2RdEC2pjK7G
MoixrV4fr939PL9UVq+e/m1H0WLvEOhptkAYZHTxP+QfXucNvv5vYCqA/+8A
LVgbyxvkNB5UNx9vLIu4V94qq51yq2ZZ7TYnOJ12wgt9uDJSAg1BfeVeSyzf
z5Ke1lLRkLSGMY3piRoyf1zqKAi1z4d7u4dzgEGv8BxmCr1kt23o4K/ak6Op
yOb66QZ+nvlhot3kJsk7eYHYsa1sCDR2hpZ8hAsRIFl9XwkBT/0LH2dw0iCF
V8XqytDGHF6KbOziM6/tquruf+Q874rW1CHZKTzvnvmNzhCi1VFiWw0AmnOD
40C9yu8eKZ/V+4xB5/yx2BtOlpeebiK1cEAILCuwI70EeZmxsNUK+jsZzfJm
QBHkcVC59LykQpxSH9Xi9JzM2k/AZg5ffxqETEqKsR7h1zq8qKM1dFaVk8jI
eKFXCwAy/OuDnLsJXwTGbXXPuX7/Vz/+11IgIlCgbrqP0j7aQXNw+7aBeCEt
a6MARBaeiJ70tuJppJj2p1OCfUtUwB0wgrcoC6QFIg8VKO7agLoDlavOJWz8
erjR92no+rYv+Eg1qTtqsY/yUyuFD6rPnL9/iogr7GPtnWcBZsAxPbIGOnR+
V0hMXfWbeDoAdREOvM0mBbDEzQVQ1dYE5/eicub775Amq7XzQhhtKXb6PeY/
1exNfxB4685FyCnYJPl3AJAe8cBisiHTCXONmaA8pm1KuetDdJVmMI2A4OMM
zOnbv/B5XJ6MKatxzymj1mWPaKIdSzkot5hlBXEKuzPYOEvTrWumt1HiMp6q
DaG6O7E5/XnTVjTkJ3BC2B9a/U2HFEoIdYvwgThjBux75xTYvSaPAb+nYM2X
knyXBJEXQZGOQQbWtEE2dC8ZVPgE7LhUrEk83X+XgJBLlOwaJQm1Wj3i7d5U
IqWHgzOJitRPC53dYCXynCKYjKnzDk/Z19Q+Rfu2wmhNK8YhJwtOOLgOQkpG
DQy3vACFESE6Fh/bJtqxSaDQIJ+193QLNvDY8EEyvVtHuI7mhSYnxiX1gUKB
raHNK2g9pUy+O83vv3vZR1cImKDPpCfg5P0RWI8JdB9y+CacYNeY6BU1/II5
pOmuGvsvJrC1At3MFUYJwC5GLaeDSiu/FSbSktTYYY5faxUjm29HKsnge8HT
g+qaxZdlladaxyoOLkP/FgPb9TyOWN5VGiWp3ikf2HxxNCSf6YzxOnJrA+zO
uoi2FDWL7kiXax4STl7Tv4myAwdJILn07G+BJjFxqnNNzQvZPEQgj1bdKgDF
8cbXqkORK2ubGKiuxOaCHGHGS8BpyzOvKotef7+AVV2mfJtwsZZ0nD9MuLYq
+ShjL6tp3pB7OkkH0TGFUnhAOciBqDXdNWKU+GPDPiI+nt/E6Kq3whK+g+ml
CYMjLqhj3mMyIwAfUubvHXXM+zJwzLw0OEUSCTkS4AbR7B5kytd7sigPcvHv
q7gCFj9XDjzcEACSMv6u7bWR7R28m966HOrISsxSGWkEVXQk3a9tMzE8tvrF
8+8JQ8MYeHEVFNYBnaIj+NoB9Ess2JGv3XSHWNRCb0nUX3H19v/CAGB49Cdi
stYnzXu6cJLZEtSy+0JeIS+TlhPf16F5MfCSMPa0A6EppYEHsPVJ/aMGT1dR
+eQJPZOf82GOo5smLL/FA0nsgGr92N/hU94WbD+DYvfAbx1PuCNEGkYRNxXc
XJOBNuuanwWtG2A4mWeOYSXaevTD1HTRq5dVFUBaiNGSF7K9w2urSjCu1Mmg
6bXzKrEB0ODUT2+n2teqyC7HzRpLXfeJJjIJABdm485EZiKBodS2EuDgn+WZ
diJKuC4vzO0nQttvWENg6gvlcY4uAQOjs9ZTWQIaqXS+gJL8A0xVgUDi3gfb
BRy7c0jpXqW04nz2bvczksq7/OdVIZrgEW5Jnbuo4JI8qIzVKeq0aVtSOZQ4
odAt16bM4BJs9IPEIOAwdaO4tWGTO2r+IUhShPAqSucMDkQNpDuYxtUJpynu
CRZZcwc0mPsRGkcXNyQUu5kVViE8chIdcKcCAJ5EdCmTFnuUwkQWE8CW2Log
GoAedl0Y3PPyqgjH2qUyXoyOGLe1P5LaoY8I874GfH3LD9IzLucTXUfqvVZb
G6lWS8ibW6AV0KccHhibSDA3lb3uTbhjQ9+3M/zITyijTjSZX+WB8COKaTyu
mKQWbnExbuprZdc5DshTdH8X4Fo5+NsrcK3GPIxMb8T5yCzmiDfJN/3OrvJT
mkzjHr/d6UjO6/8S1F9HpWmTTZE5NHVj2WUi/IBzKvlN+gGKxH2EMYlOa+v6
GBHb3MgByCyHrpp7v0CkTI405apGbdNmVPdhgdAZbK5Vk/MLJ4rTc12bi5oX
vsKaEq8SoDSXmBCXQbDl2rSvgdtvIBdjhB4eVXzrmb7UCIEukITw7qndfcLN
cMcCu8itx4X3rttVrNGN7TqwsZZ3pfpBcmkaFOO2ESQwzkxsgDutVScIyMEp
Sgi6aE/Ie5hv3Ewx3cI+wD2rOc0nl7gMKRcA2ySk+j4UIwbaxn8atUIoQGF8
K1iK342uf1on6d6bDYIoK+Io/xMC5BGIGB3SCi/kYozttO4dwjIfvmToWb6/
3lWwRB9IN8CUPLcxNeOMYEm+mLXZ3RsvEbX6nTRjplPzu3DtmTshMmBtfFv8
UatohTfwtZ61yS6riq/FQ+bqGmSj2LdCNUF4oHkfENIiMbwDRIc0Fq3A2I2q
iCIX0j04d7ha2N+DROKhxSh9p3OBhaICll0eQLUYKzAEj8LmluTS5dv9XxCS
hWOfmDkT8ZdzJUPC0R6EfDJYYU2A4O642FH20cOsemI1JJ6D9o+GDilH1zQn
a9nvEF0EuBDILIVx+hC25wK4X0vLivNWW7WDAHBPiUxMlmeZ76ou2MSabTl5
05zFGt7pCX4LZnhXlPlffzmoeVlPKY43hnAkj5Bu6RYi7hic1ZZq1IvpslWV
lqk51/4LQZ07vZTkDXwFSWxtX2BLBY/nrZYEVs9ay+UFJkwl1oycNzslKPYi
Qj/Jvf3l2uELytwqJq9idhDFhYXDkfu5u34Hq+yfLZukkTZwT1kuJ+zs4IGx
ZQunaneWQEXJ91SXRhkSnb9c6xe0dY6x5b/jeNwbQto19KsKxV8sztAsgsKG
0tNw02XWPIMYUuJVP15z9vuPOkX36uOX1i4X/k97hf3HNlFx6kETQkh8NPML
Xkn571o+1tm6foooF8LGLLX8neB4Poy+Dwdj3BbQey73NZXsT4Y5o1TOyWa6
y4K3QIRfGLk6Pgo9GwCiXyaweBsWtgZRg2lZIgkN6UyD8/FIO/PoccgPUgR9
8H2LL+oT9l+ptD/o/kFs52tGPVe1xcO+jeO8qaSk0zBUpMz1A/uptdLcXiCk
g3LQ8B2O5DufmTKP2NXMLutfhlJ5H06kTEmzZVyfWa1wEbHXb9sAIqdQaOpc
EuN52jUpQOu75rhmh16PcVHUQm6pZKVDQTN+ZaJNFamQKAV2G7H6aOYXN6d2
iELzo/lRiMDcHVMHjKsW9AcTRuT3WmXJudeBVuRww2Ku6tL/QwrDdfoMEwm9
/TndprGioXYrzY8qbd0rSxdv0tKXGDR1V+b/FBrD5oEmLFuz7kW8iC1liHSv
9I+szMrET2E58KAX1mBN04DDzAGI/e+O2Zbkw6/xfXuwQl11v+VoONfRKoYs
wJHPI4hh2NhFUHThAr1eMwEgFv7CewNKg7jG0BzmcwOcU4rOq83Kt5zjFV22
lVjFFANELfjCYhuKaL0cS8NBQqErvAM17+bwuQ1vexJF/9gZeU410lw79nhk
QxwMBp9PD51LK1X3ts5RqG1oeHevx6Q9TCJvAPSvoMjzvvznYoKTbnPPBZ0t
DhJRATvGWG0xLxESdvPA1fT1g8YwRY+5Z9jcZSvMJefMcI2/2ElAGhg+TkFt
sMWXuIHD/FxXyq06G5upRW6hEHh5lwoap2K2KTZ3+eZBkxDtGwWfVkzR6plV
IhgEEUc59yLclDGpsDGsRty3dH9aIwQrzq0gsGil0HIU8bFE4/8P5arwtbuW
zKX8PpB7aQrjKZmyjLqjcD6txdGc0lJvKPXJs9JPTXXEpPg35Kn6/lNxd1W7
9yh3uxoGbVkBghyH9utuUOLVLHJf+lR1Ri9j+brgcnvpcVhMKaHbHwWvGSkZ
LqdAe548IWFVM+3LfqOLqGCmgffNE0zC3VldJQLG2ArHBjC1NxpsfKyInqDt
RidfNSrgQEFvJ0w5+SsgQ8xLFbSosWvuQhLq9xau+QQT8rEaAOJminulKwEx
XoLWqhW7oqE3epPVPis+HW+QR+5cxuf8tAhZkkkoy8rgsV00cLsGmtffGkEW
GeuMZNIeSo3e2H0KJ/J7JIM5FxRrywu6pjYkmtqo/RYJXC3WoVxsHK93NDLO
qtrFNyek+jiqn8c8J/j6UIra02rtN5A0YIZKMXX8Z0yodKJmNqHs7wcbo9Lc
7E0MHsXIE8MMSvPtJCk9YTRerep9LRILHRZHf59nZLoAjgjZhS1oR/IGr/ne
lmDH/fa4E/OXKsfKNzv/d7r05/KMGitAgtBau3Hf4fGNSApO4eUjuUNqMgBX
67YSSn2dshkV0cgXorEOUO8W7oYnyUb3IEuhbQse8H6q4lnfLfbmGtTnt6Ic
gFpJQp6itCFl1F4x96bLAk2mxXdJ/jsNQd1oMMVI3ZtH6nfFViUYLG5VcuTb
hpOBsSYtJ3zOCCexl3tGejIChjyWXOvWNqWa214kE5hsGzxa/OXlAld878H5
db0gdzwE1+23jOPqepz97TIxf3lG1d9q6wa1mm/SisXGQpw/OcWB3979WrFo
cjoS+ICTLlEnBmBDALPjfyXOLbi0oLBCTnzFAdVTuaMUQ+Lt3zzsh8OT9S5Y
eASE3xYsXpyBunYDHVxlVjDApEsl/tzDqOYzaD/uqwCZf43m3/srCbqV/1Co
+ZCl8xd7nb4yYt7YvyidrOBUvFOPDjaZZnhhkcLfa1Z1E9MgN45IxW5ZOzR3
K6boPdI8e7FTzb6DCJJ49WVh3oZVd8aGdt4aIKrbRXm6/e2K4/sbCK0HrU09
WEluafNDz3G913Y3F8n8Q4vuuZxf5NAseRMyfEJffIYh7r6ukaBL32+e3YPX
1x49vEKUihYLYu/xasFOHDugzouth35o+9K5B+x08A1Cnpr/iBeJka20sktF
L2xvz270p4+SbNalLafz2OfyC1+p7jejiFuUzu/789qivs9JD8a82lZP5Fry
rHukT2md8tOLiP+6iuHXCD50F5sh8mfoTU11cMEOqNNSoW08awlyARwmuLa7
YeqgA4hwgLWbmnxLJXxsgdjzhAEuMnGNN3UKUHJLJf+aGtDCHkGR2GRgYiPE
0SNeCfl+pTSM3QS4ZTvTVYpU6bdKKoihd+NXeGHGBCi5XyKQiO6AZC8zQSo5
W4fNxTKaEydhUPp2v67UarD5kpXtUDFIGi0m7MYpMJw9u4aR587cKjKWECf2
i9Uf/4P/4gCK+4J/K5MYG1w6KX+bBtPRgcck/NQ6No73oXlxWIhZAs34LVWp
bLZzUO7AoYi19QsOMmmqmKJHDmSl/E9jG6j4Lf/u0b9QfWTBS+Rbz4I1jOud
DFWTdAbs8xcAosfKNJdHdr/Zzvged9uXZbz8WVWHvUysnTD0e4XFRLSaR/lD
MksFOZjcgzouNaZCXZy+t3Kjv8H2bY8iqQPX8BcPQJMmMrya1fKvGMF0U9vt
LBEJZtyDOPAAg8uBhxrjBjAI1wh2LVA/2/SrJtpQunQReTMpIcPAm/4tu7ll
sLyR2dqXK+oKwFHWnPA35Vf/q7/B7B/+VD5l80R4HYmIpXAfiPGK8ztLVS4u
9Xg5wjowjM88LvCLgEuwF+gv5gGi/m49YINuqGRQw6Lp9pkYGLcGspPMzkFP
i8f1xQOeCv5Jnf2ZjI2UwSBFEJ+lHMnNkkh9/rxgy+Aejz4BlNNTcGKQCcF5
OKqRQ4424266Hj8o34B98FaoMjp8RY6FlAyGfzeRttupLwN6RGh+5ZkMO3df
MYcDQrPK1EFg0Fdo8du5CFqylRE+teCTf5QeOhGiqM0Gddfpz8dxRFgcRWgi
MKrbZ2N4jLlhstndtXVVBD18vXaOIUFvEm60BN2otQMfIfNwFovJtpgh7OIU
+VO1nq/JJJlPM+OxA0f6z0fzSYJgcfR36jzLuWRMUGX5VyYdJN+yvL2QeCKF
pdi+Dr/RIf8XcrFmmZi4MR4KfJ3Ib8SBdCffgVUq2S3xMlZ8eEBfLplyjA9I
4vLydr8WNRC8jmKDN7xzqQD5PRVoWVzdNxzU5KYnrABiNo0+f0g6Q/aRPHLh
FUbfc7t6u/FS/6Gf5wy0DHX/k3DyUuL6r7Nbl1uDtqkXeAFYEBh0dPKoY4sO
Mz7S0QaejVmq3vK27t2qgYUd0I90y17WpeSKz4puznd4G52ERHjtufh0G5Ea
t/koYuN7PCPa8x6ZfQ4h3wRJef2jwxekRtKwsskJ4C562t/9h6TZgpUiYWjR
b//g5W+FmTZ32gZaTXGF1VTkwOx4fxjM6s8clr2RemJUaZIct9vwd3Mwzg6N
WrwWRLjOegC1DD2EHyDzAnuBQtKsydkmUIgPL0bD1yXxl1s618YbTBaNXsYl
5qY73JQeZ5mjBwtUcd/J0az5D66c2I8HCbcUZC97jGplQMeJMic3C78jse4o
rg0BL3ItDwUmrtQvkeZX6bTxp9tfD4SyRMtbq9Oy2Id+KjZdGYTCkvZu+59Z
tG4ipS7N/J2VsG28jvmMa/T8gx+G+AlAc/yvutqjqZ7RZ6EKOPsFlR0LeC5l
DvAtWDScF1C5ctAdE2OScXT5Q6zPRShggw6k0XAf9Ezh9SsL8PFc/jJm1MjN
KrEgnlpkv5DxEgpZs1RHRfuoNFCvrUvTPoE+O31yyO6WQkw+NrjQisZLaK37
NxuXwua3hk/vojzaTocI1NH9Gh+mWUmAuLuXnK2edEMDCuTK/400CrA37v4E
yzZwf6LWGc/9nj5Xbl2DsQ/Jfa0oa2o2/JLEiE1pP87OMe2oF+xPKuh4GfqJ
3igpFtDwWTf83dSJJmgCGS7Ps4f4GOhkdRUyEkov+pFpa5DNCtxpQsytWGjq
I1f9YIBB4M37yYxY5KkeUA8kZQtoPoGNyMGBeC4iHKnPhbLjs3uDL+Vqnnyu
GR4um5zoX+6MEjf8cZ7njBRvdexd5Zd+OnkAcp3rm3/ERSs2eUhhazf7LEjw
ULjGVeF4M0T/C/g1LQzJzWk/uNk3NSmErN+BbRqabXxI+0fQSiRHo/O6chaZ
rqnhvXv6HZF2Mq9tex61uQW4HA5ntwMjBjX+ftea3e7cwOUV3GHIMxjvpLnd
UT/0fRlVUfns7+O6C2n/W31CfachCT1y42QAsA4IOAt828fDtWA97aG9+usN
9Gm7rgtIiJ7cnKLmI2nYArxkBIMnupcGtwlBs0rOq2tmQB3cXU4YG4Wuz4TF
3F3RZhxWNo2K1FZH/BDHh36Kya5YIFD8lKmWWcAkvX+wsLbklThx2d9dUxER
gvooXwCY9jnuZfgdEWVksMlxFqg0NthiURTUFkkqZhVYIXBJV3yZn6ziLEzi
1zopBPm2tDav9QZmPWdXy3Hga4qMakcKfsDGiZYDXVujLaa02coWu2OEDhj3
37BYlVplZ6Drww2g3wynnSyWczx53YMT5P1l5yNkKPC7xMNGV/p1onrtGFQT
yHw2Po0iTWDGVSzKyurGhVPTRYIdoshkZTB477Y1slfEC271NTvGPhClX2tx
DM37ge5t0K5/JjBmBCP8K+98PazfmPf9P3Bu61RKvHt/kMM/t6W4jyQNyOvO
RfReDGzm/Mj3KHwYi4SA9ps5sqsWURyUF5s1EKL2VTPiFXhFgrxoABQ7+uEd
WBM3Rksb5lTW18BVc4P2gDxS9gMz4a7U7XGT649mFxPuLmNavYl1F3IqO/qu
xrHWiZ47Y8JVNvU4/xqj41qjIuet7j14wo5wcFb0HKWE9CzHGkxm3f0xcgkx
106rOpuN5WAqAGPVeURqoMzkTcvq1YhNrALtu/cgrBhZMxvhzBVytIndyIOm
0rpEGHfNtJJJxbnha8pdj7Z3Zv/08UAMatoM0Chqa25sqG30Bvm13bUJXMrJ
aKhL1dbVu1v2v4M8ONsqRZo/3WF3gWDsdTGx1OSKRdIoFemFukgmNmKfLqZ5
EQ3ODjzHQRGvM1iAAnrRizxWIj+hkHmBfXrQHY2Nb1R2Ss2ammduZdJhOH6i
Gw1lbvbXfq6xD7YOjmOVYJN4kBgR6CWrINh4Xvv5pdtKSwsz5WbYzV0+4PZl
t2OzMpyy+KNftEqKf+hy4CIVmzVQM9F2cWZYJcdtGWqSZrJUANa84ptGMyT3
YwNBWFT1zplDIERY08iDaBXMTBpCCC3dNgnQjKAVnWk7HzX9fC7OFL27yWGl
89lCp1yf0BZRVI2pwtiBb6CDlRDKY43e72F02aEi0YRKwREfvlbu3cxzHsXc
ZajQN5b2mzCdNFipuSZCDYqgoBRCcN4ZIbE4kxGC07PleJ/4xqolAwzHLBr1
lMalBJZzWBoI+IwrGb9H2d+Fj3qNaBYrkxjt6jD1ESceLnitBKqLecRxQoa6
qDr9ae9KP2hqh/USmbiP1x59cVrjDJL08LmmpdhzUVMv7WCmRyzU/yafoHof
U7bZTZIMtH4wneyWQFoii617V7HrdLGwPxFlr8xfHhGp3E+XIxR6XBUuBb8V
u4fnNdv3T1r+GOlYf4etkboDgcbq68qce2C7amUCqaThaJf3syCDUow5OAbK
PLNF6mT/0ndNw/GceEG2ZNHM0Cmi0eu3ke94qP5INWfGyQ8D1LmCQ7XKZ/FI
pQ58Y3c3EpsI9CYsS5oSnl1B4xdCPNAA5O+VKt4UEOUV0hT0zDiti0Y2c20t
SPrr1+qL7vJt93TSXloGxZ7TGRVrBlstV8Jhi9q5DOpb2yP27IlU3gsITBTO
Li3v39CHvRBgCIAYlquFnS2PagD2QEQqI6+Uad8NBhjreJmyGavAO6MMsATB
UFIysfhU5Yl0cA84VTcJJHD4/Hnqf7h5RC+gFU1MBp4hgbW28920gFNZE/Mt
BGpO29RaQ923Nf6G7ag2b5Z5XIE51p3r6nGahfBMADOtJ32lav4iz4elm9pi
3t2IRmWnUGgf15G0rrSEzwnzwoZDSsN9ltnUjuZIoNlpgnNwColmkYNf/itd
RnB9yqVQMaWEQ8NGX8VbX7n0oCxzKfqXDJ1OPUn1c6aFemNc9zr7jd5H43zy
3g7ePtANJvKNKGYE/y/IKGUNveg3dthwltNaoCncwq4M931xvpOCbhWNJT2/
BmhtAZpAmjM6jqpcGesArM3RQWg/9TF2hq038Dp5G/VAcPD7ivwpKD+Z5Obr
2uKGKAusQBpESIkIqnZXTUalXkWqp0uCndv0mmlWBzWcc1u1KptjHj1zmBKZ
D84SK6OqZxDmjBlnWywRJDyHDi23s2pDTmA50L8Z/yhYh8RmccNndsOIUXVG
cGSY3wXQnN9gwtlvnf52yd7kIIfUF3aCuXr0ZN8n+8Wpv94KTBqh3AFUzcRf
rXMvnSOAt1QL3DNMCypLpVnDkL/GdLveIyaejcSLjiu/+Yn7U/XhkvrKGvID
ZLRkYhCa0yVk1/J1Yyzv8Hhn6N0OVroAC94HZGbwagRApD/ozya90CkokRk6
a3YB7j+Phr8wRBKQAgK5FR+A/vOPVh995m7gUrPa+D7uCJhy1zuV9CFzcM86
K7Boj9St7TxSH7DtB0yJtnPotMjFgGjkkNZUjWoIiVps+ehUW0nGVRHHv1qi
4ZmyjmukkKyt5aUyjla8BFjRaSihKuQpRfeVzlyPt3DSNYXmpXfzTPJPcgo7
yE2faGpsUW1JzNORacACzkzR8pvmOhZ8PaZm215KPzVCKsIxn75rz+qDLHso
b6dbb7S4QF1EtH2TALPpythTnMQNlAAp2Q9Ntb/nV0kJn8dBIxpLzpsYLNC+
untArFdbpI1O2TYri7HgBJnNz8fjFxxqAlUmDaxL8xK+3XewltuOuvMJLuN5
3l951LNarvL7r4HW2o2Tf47FF3IWlvJ+5qgD5267IIm7jtWMRpmuiqpH6x1Z
i8WjnW6pDK8krZvFLF5KfPmji8VjoDnXhMGyiSos3SxZvHIXNDjFnGSvszEu
oRXrSeIq99GjSHwW4v5PEekg8Lv+KXfefRS50Dlrml9ln02V6csdBMpPR0wu
PLjkDwhzzpZHON8V5lMXX7VR2duP8LUC6Y8C8a9j5mllz/bXOjpD7R1OWm60
e7YVNpAR7hLd/MCVMKZonR+uPyslsCI90nj6OO4+rrSsLpDBCh354Aj1Uj3i
TpScGsedclGpy9QVcb8Ve0jsQ60YC6ZrUW+zCSLwp5mMYk6COH6r2pct9Tzm
5ObNxTQw8/TG2RkG1GfeUpktKnIqr5KaeaNsHqh/zDyV6ts3i1P3ks59mK/d
pf87MTcz72VZRGHfgZWUICn2WQI19/VQmUSQSoFwRxUp3p55t9vPBw1kDM6B
eD8hk8SnwnIt7n1PJVJ4zOSR/5HJhTQRkPe/GfbcQeHqjmo9JAHAV9sGJmCn
44RonFBcL/ToZ2WtanEELerYtL5lSCGD3zvfw1QQmDleWxUYCeGz3Og57nEr
JX2CBKfXoXbBuM1f/tFWr/yWlmTqlbAzmM9dHQ/CqbmV85XRXDLszDZBRHF/
pUMA+7cRI75FpWYaqlGxiEqeBiAm/1kA/KNwQ3z6aTOuD7TKMdsSTHQNj3nd
YYRlcvalggCRqzFjqWfchhbbFPrhOOxCznvJ7rDHyibD9o8Ibfx64eigGGc9
5zzIvsFTqfPCtKkAf1DXspxyXGoYOmyUWMIvasmOqQMetpvI6lCoJTk+7/cX
7HKUS+a04b6uSW1VNEwIgZOeyk9zbUTUogBWMAq6pyRTrwR/s5nZkZBSKyx3
wJzZ7pryJRx4e2R97XBqsJ/KkCPpH8jQtP2/gdWm53XcmQ/wFO/7JR9LmJYo
tYC1pYLlOQETuqmhcUwmX5i9zwJAi2Mdn4SuwCSN2Sp/eIa/qZkajWood0Ni
Lj3kgECg163QJFFBVexWgUKWmTKxqbV7TrrnQi2luKk4jyZG3uO0znwzuSZa
OKu1gRapIsy557/iWCxum5UxgGJwQLk/DPVquL1twA6ZAcNdmtuGBMw+kgS5
zB65gSWlFfkQb/85EApsTHzNT9ysq64OLufnsje7XPURWn3H5LtjvGBH0awE
zBZ4hi4ui77qyY3xADnVkH0pnOtp8S46Gp3q160OpcTSzmlPzhsuVrhNdJge
bsaOl9IWdFqSClUPIduth9HzDhyPrbaD0/FedzBWO3utoZ7H3b/pKPxT0R2/
wKNQNcsnxnsgt7sjaVogu597snmVaj9bv4838hoL6htl9FoigSVTrL8IMOb2
4ztrHdjx1QUTLIsz+8G8Qh5eloJJ6EannUD+zEu+yXWUFAFeILOsMQ/vzH22
3jS29D8+lLFZwrortBdM8B6Ipz3njxKmuLL+y6TsT6vke9KsfFKPf/rVciY0
QGxK5WU7Pybe4WjLOxycFQBRHLZCRu+ftdEUqeopgxjfSuacr9mGNs4plhlb
+mZpHDaQmtOeON3TeoA1K71DIwL9Pwq7uz0FjCG3BDoG3TO1Uu7zoxyEEQD4
jg9WMJHMgD1KaLmAbKZGP4XgZgDgMbPlpt76TyJNy5k2n8zoBGqKfhoEl4V6
F519GSiBnwmAfdzz8JXNOM32LqRgQaY8Nl5shKcrqqKOffNuA05HZzEpAfF1
OMaAvsuiiHZOFC2B6qhWp3wXzqhMiR6sRLrw+kXT3GiQXzqEcrpNtMsMenZ5
tKr4tVG04LdqarzTMs5EOEffabxzU5swYpGZobICFZs77pZA5XJ+ZSsGk7KW
oiKVD3+LLYIWs6zPX52gxwHdUg3SUzFRT3sCcL/lnfFD9y12stzcKTOdc24u
LOe/myuGTGRVNRq6PmXWZONMF40j5V7CtpNmzyXQdLPwDPfnf83naPPHguYc
4bqkuID5kmG+I2R8l8wI150Tr6WngPvIK1Jd8pIhOeshHK3+zwnAbr+rRvnc
B4wDHv/CXQm5TGf2Yr0JHeZ2pwg1xO+nju6qoRq7YbP2qViyzJJ1GodKHcRM
/2d+Sn6GhrWXt0dUyfQjOz0BmRKDxZq7uOHeBxV1OfLIVIEaHRU3VxpimrEd
Acanji9Fv/Ty/9kHxUKLufi24H6c2+pyygI=

`pragma protect end_protected
