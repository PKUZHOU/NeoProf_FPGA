// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WJL4n3cxsGna8QZKw7hjg+ls+1B0sbGJq3XFQj3eD9xFv4Avz/wLo4Qm+YpA
m5FFIpPoXRtgSMF/r9XC++CAqvlI3OlsztGpwjnepQS2wt5gjj1aKnMbrEx5
5lKBtQ9ZEaiRfghiKVi2KrUthPwENnWqpdTSb/I2f5Mn3mTSyY8IGSJRYpuY
VzxJV7f3AaAEgTL35YWCUPEfOUfp3HAMNuV++Ir4GoHzEsf2dwxTk9bxCB8T
h9YT9xnk7nsaPOtOy/MftGmy8vECIu4INKG7W633zD82Y1Jt/CcvduD0Kc95
toDoTONFd/Xz5EM42kVIykLFN6Jg32b6cAey536meA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
JQdiAlJqnKQ4SE/seRBIrNZy2xm7UXK/ormObLgcFl2JE/5KttuntBqevj/s
z07hJfwOQvbrdp9mzSEo0hQ5fSsADEOGRhkgA4SD16uInO17zE8uQI08gnxq
3Ew3nZysdYHU+8BSh641X/wtcUMJtL6uMYmz8lkK3sx8BKKvoLk+Ct7wPZOv
HS2eN9Ih2Wbg0zSeX32aziSMmOVAXCC9kiwaQFnWzlxx3O2b2IgvqnRHNoGr
1FxdJp46M3tDXeVEGGyQkBXqTgS6kcTzRA0K3ywdK+m6nwgvuvR9c80umBXt
rpf+poxSWMos1WUJ3Nx9ETYBVWkHNvs0smcWPglvzg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
a7HXWw+52MaAMG00N3GVOpYm4EyHmD1aGwrb4MJz9vT7KDPp7eFRG4uQL3Ri
jcZKZlfeigdmVZkILx/1UDKdwhm02u7corvdKDbQD4PrNTZotUqMwrxUjaxE
Oxc0YyV2mxkYgExJNFfFizA506D9rZBmDCyCSDzy9f+S0CvZAd/KwvBJrjvu
fCHcppRHfuK58YQZo+1Z2zEvEMFYjGT0lS2NGsF7QrxNJI8JokGKEiJ8tPLh
GHVJjy3K8iXrly7F/0s7XSfyVODVJKdNAi7iofEHdaQHXGAN5oRhPZWQ6QXr
7rv3H1G3pFv9xqU318ljgl9v7ScOwiZoiukz3SH0tw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
kW7O0wyFbJgxyScD7jQ/cOF1hmx0mBDXI9x2SxT+0MIFIK5RHKgq9r7Inssj
FM1UovKVLn7ZXKqE1/PBGW86y6/mwgTvn8A1v+xDZEJ3Lzd34Nr5upeDGf1M
YCO9TRYvhxtK04Gd41XuBxXD2JiEpdTGbhc0hAhXb/kcAizWtrc=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
MYCzEJDJlIt8fNg7ocJdJjoZqJ93eawgsYt2MfEssOjlZfzyzqGloxF+cUjy
xHqKg7VrUUOFJwdqwL4fAOXqkBicxaWanuoPl0RO4IrGeWtdl6FfCt/GqVgx
ONKI7k0EqYyiqHCWMbt6JYxOQFftdm+9U3gEtOylrD9XFfzxNMb2Ft7FQcxS
aG4qsuX5B/YLWs1f4UKSr3z+MVgfrgY9PawL6ghnCG7Q2+f+LUt3Fn3/a4LK
M8pjovMa4nnukLAFZ2p5ESkp2rVOEoZAaedACzi8fUqRWq4jGRMi+XmHnsVw
wf/sXCPNMKOrLMZDM1IxtFrkaLYWsn58lhtGaBDgRXlQLDywsvO+dfdeRjrC
6k/OlUWMOvCh7/LOUWCg4dQbyJTJTco+zMtobvaL2ChJDB7X/qhKTRBJTsJl
BsSSV1Aku23HCKiuDUz/Mzs6UX2swyNqpBqN/Il08EICbV+0+De2qhcFBmxt
WezqHFVTAdJaOaVTalmiVzdxW4T2oJXq


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
gLKGdGL+e7rOidsRO9IRPRPnjekK/7HoehmSrSm1T+6zbGEFH4K221eTlvev
Gt0SEDfWbVq1Z8ILnGT5vmvOwoJgRQdi1A6225waM5jfRqUDiQdHGNp52Eho
9/W2pJ2wG3donJnTe1lSSqeIvGr0egXtEyLq6hU9t3ZHsOLbUCE=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
QE3b/kNf9s9jdZFKqEdbXUGH3qS8s4IvCUrFmvdMJgYyIc6dmgWfqNCbd3BO
At97JZjxgPNYsJ74GMZOZXZ4h6Cclf91C0GNHLr62RHZjfaL6CApZrwYi5ek
+Ivi7O/OqahoFPKV9dEt25eQlT8bVMdFAVK9cbRrOFBzN6nxBxA=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 83504)
`pragma protect data_block
ELgJy/aM8RQ7MQNzN++cQLs3cXRJewVDu2d9WWm6MV0Crh+WDwjv99H1ocsl
yqwSr1kCFlGkwyyQn1dTgptTxs5THgADE4BvUt1LHCqup0Sku+Er/prqa/If
qv1qUrpDgP70E8KJvTrVDINVupDlSA/V7bZSQ4mi5AgUXSGufRLjDj3qHHmg
velxOGg91/pKLtFYlJ/WJEVr5wq0E8bXnm7VRbbChfNNGoz9wS2PQAsmxJtU
OMcnFu5i43l4jLVAZl2q94WmRj9IUpbl+wT2yGUQCeIDthm75o/76Z6esn50
A5OQVdlCxH/jgv+9d/qyxo6rWtUFDEGpKZfdkRhErVeTOUbKuUGVzuZKuoJ2
os9Su/5GtUWQplLXc7raRcgm3R6XD9sdwpJIIjkpXIYSFq/+xgd/z+P5O137
IjLYNT61IzBp7Nua0Zsv3PD4o71DVdTPGxpvvwtPraNvhZYwl85zFKpkpzXn
V3TSYi7Wbw1jWx5AMweUiCpekqcoU5zf5uaTGx12QTRu7oZAhZs/C1o+CI9P
8bI/EvO6NuFKzN/aoMUn2UjJxa7ftE9/oivp5mjUpaE7VoAcLRmYj7ViQrrt
KTlh+qlQyv8rMoM0Y9Y/bq25B5Bx8o+E3iupQ3QvBLEUtZnxDfPncRlOXrJk
Ced4ydIJ5I47nvwV50pmAns7hMt9ph0e0K77frc0JpuTyjcC3yLz7a+RyYqN
2TCaz1Ie6+PqEdC6OVnX5hlyJ60wH/5KlnEsAcN08HeGZPacg7ypKpuOVfW7
rMQrCoQVApr/dmPxhmXorCltJWMq/jWuoc66Ygu/jiDjqED9Q1MDSddBRzYv
vkisrR4NLmiE31r+b3Hxq3jVLzEokv747t+eJIKBguyRzF8uadcXL3tNnuHY
+5UpD6e4SslApUsFjz/M1xYbghBb0GL1oFJPrph9uH1cUdItaGf2JkWYziRv
VhW3Z9FCsAkKJM69OAEcdqHWsyuLn6xBI0mYUUPhxZdB3iB8s40SrWp0lxmE
G+UCVyYJdPtKAx866wXUuhmd2S8xf2ulv5kJcAMEjos16R86NfzF2u4Q6Fve
r4Y+UAhHlrh6rPgGEXR7PUTj6Hd0sJFchv02hoQMR2q+nzqgu3JiUK3g9Kb+
HCnlR2Y+UDQK2hJ2fOeQrQeNk6DGTfjZKUqyLBw+0H1o50Jzt3cG/62bZpTg
6DsL3A6lfga6pQzHgXxnGMZVhI/EkkOjdhMtbHiukawnJGhZGv9+GvFBoYOL
j+fOv3BJYdo9a4aXNIz+EzabAA0rDSSUqYEH1vd50jk8/oif12Cqou37ZKOt
fAfYJiYOvpwVWdg2UBT74gajmrbkG0k4pJtBjnld4B/Y6/DkwyVyl62i3N/b
5K30j8+Fb+BwCPMalwIUSr5Y+FIwJB7Fjoolv8iE+Pa+F3XTurkILsSjE5Cm
jD55umo1NI3MMCbYlsT/vwgkq2JgsvZ6+RUB0tl9DrEl5eI6t9Mbbg4Jop+k
W2TJeQh3nquCEf/9QdKMVhdg2fYpNyjdGsBstxXNyS2+ZaEHMdc/awmPjxG2
xHdQD/quBKdBaQC+xlZHQvXHDrWgDFcoAkawEfYszNC2z9t8lRdo44g9Sjdh
N81bmlAi6Irj+dBEmo5AdSeRrwZVg9MqRkqY5u/fX4yCRI21q7J5rzVhJZCg
IS80shhW3Z603vY8sWHS7Fu/LTkzqDbCtLisrH4dfIcEdzZguDhkncT6kUGX
bQYTIK9UJhdU5HO4sX15R8GB/1vHIovK18n32xyurzSVxmyFCWxzWJzn506g
dRVJsUmqyuxs2wIbtmxe5pBwxeuIaSw5mYjPyOij3tdG7bp7HNen7caL1Goy
JKUQo+Ggh6sNCk4vXYAqS+0VX4ToJc17Ty++O2ICiHRrFCSco+V/t49wQhyy
Rsbi7J796B+r5u8pV2vTt+2Ia5N8M+wnzpqkZ6k9rBGbj7dzTP4k9l/Q785H
JgumvZrtqVw1JaxzrXFXAXrDY9M4LDtrC75twhKdF5zkqZ2VWFvTah764mDQ
WYvBwILvER3XaLDhjnD18a8YKDdvka/GvrkmvWjtuL08y2+RsYFgqbj1CSto
nHVewNdpjMVun9H+bTBWy++eAs/MCBTSZsFA4kBbTCDjPA81h6UWaaRJpHxT
fwxEpMHo+MOxpv42Wjetq96Dss05XORdoHUs6wJIMf9xk0B1sE+ewPfA/LUF
VJ0U8ek9BDWjTUGJkRs+Z4U+RRlwVH09qQlwoZxaWanBOme198V6henbYHfm
MRjeihzDbzrusuZp+rFjmLxxw4UcntypzMyyiCGUHxUKpLJNTWY6v/lPt6Jg
NFuV9l3jdxjxowa98HM2Iww4meX+PhZCne2csYoOo6kMGEy2g/YDlnWk5iMf
uz6Fd/KCUaHnE12t2h5XtWMZrrA4DBFiylOtVDtCrP5R7B52W3i4xDRHZK2D
OhOcfi7dSXqrjnGBDaPBE0pwZdroAtxqOUgB4XuJF0FcKmZ30rWw1b32E7rC
TJT75nH93JeDOUBUQTGwvtI6o0w46WQaZvpi74eP+5fYFGmFwIHNltnPMb2A
TNwu4Oh4CEd043pCFzcFE8lFljf7EGQzpbDaRP7p6WO8HxcJWy7Z5BX/mSXj
i7KAa+YGxbzs6JmEu5hTg4y2EOCtaNACiKBlB6CBszga+HICTSs+PoLQTh7u
PbG9VQB/zg20LofdeMLRSA6UCtcCc0f0d2xSKi/jCs5u6caJ+sm90ldOz/Qn
ypGM7fS2nZmQkN9uef+z4eQMaZ6IxampeCDH+Y8PQ15g97ZVxEb7PS7vmaZ0
bd6vYfotO4PEjjlWMhjC22rAKi/Cynuke21QtIAOGekXFnQO1G90FPdy32lB
L+qMHFVDeqGTyhn2C0v21TZhrRTEBnKEVyzwnBnak4+zOxyQcIQV+xZuw1+7
8AI1BwZyeyl1d7qs+6btsjU0KQn9QEqMpJFcYviGPXCqsKvJQkFi93pwK9rl
+AXVCkEW2D7rhGb2dWSr2RfaaPOIjS5+Czlt94DB8yhoxlRtK9BmQ5p+xdh8
EGg9HJCb9ewqptLktzoNQf/XlEjLuuVPjvi5gjATcFgy8FzAWeiBnPy9v4b4
N5f9+1HYnozgFpgqnhxWOPVoeeTXT9lJGEqlt775VqF3HIiUYhLeqlMxaNmL
LcxLvKaNIEZ7w7HRx66Ss9WJnSmrJU3an5xIO8cBj2FqD832bDpijyOYFxK6
rRxS+7cIvpuKZwe+AM+9TxZlekRkdrxoOZAFOpnwJmFM/tSirTS06blEeNq2
WNMJhoNS8OQsAbt0t2WKWjYPuElN3Sk7C8viI240ehEiJ3qAM3eddyAJ24qW
EobZ883g1+tYls5IJAgkvjrZYHED1C9H8DPnfFhx2k/3PDB4J+rG1kun5B8G
4TBTNIGHlu/jjWzzCWYYiqa+qzg0mSKckTK9SKhlZx0wuxW9CIH9vnCJLIcM
T9+eyuMDtycae0sVfSQ7mSP+9k+UQmlf5wgQ8sRUboTA0y2ATJ6K6z33Kq4z
nI1mLqyJkirZJliC2VZIlbKHHixCgRZ2cU5tOhIh60yOgEOk5WYXvvz+pLGO
v3e3zGVYU8dYTGd+iKruwzWtTccCXgV2/A4g765kskshHFSgQT28cRRAXNX7
tcHtHL3N6tKHeCKT/FPJNUT1K3YP66xdi3rBoSJGzCsJXxtEl6tnfRM4xQfI
XMu1y4OZuHDBOdCSMFbFZUHElAVj1Mp8m0jncpmgv3AOjyceuXC7XvDodvgZ
ni1JMpwGYNH2E5GgQySDCR/VhB/Xy4xuEYaLbtu0PicSs5gBnO2mRmuEGAfr
euh79K8PCuEWh2aiW81wpdBf0y4NNxQ3MjcgkeeaW808Hrnb4q9tIgJ3X3QV
PXIa4xUDAQn20/9yQkPpiFKsb9RfnXF/1YnmUxffgwGeuwVQWYcIU3IQwc3o
3nH48I+ZTIj0qq7FNPM1F1ijCl2UablHowW+L3tj+xhAS8/PKRJrH1uIPvdj
EfWklgEXL5Z2hpjvWDKnB1H0qTsLWMiRkmAqEG2pUaZ14wNKeOUTY/KUkGrr
2AvBr3KXAm3BuGdL+W/bgP5FAUcHZxKCa9cwYo5PTH5qbo/VPa36k4vNKbG4
iBWBCD16a2K5Q6AxXp60InfTrSguF2QR35ISc++uLVwonGcGzaAAblhjZPXt
bBtjApAAFxH6GoQS/Yg3+ll7Le2Dl43SKERJ+wueZtGydbi/Z4TZCrCvFQvn
bJdHuNgZ4pvgh0YFOhfo+UwitelDwQWzMwD9m8NY9lVqVeyHCycHex5o2Bkc
BHX0WxqacmNXupK8jhCbcyjEtnGJ+i+jOCk9NbfmMNz8w/umNEQ6s03RGs8c
8TY4oAaz0mug26GznZ4JPRMODOZ69jHbmsKTCArdYyWCEmtRvCSN6GM9i/vN
yNoUOsczV9KhnojU/5X2SMLqSEONmLtKkQ1GpkacKVeK8pWpBZt7OsrWg3//
2cvMeLCKH5G7rUKz3tSv7rVfo7yWJICuKhLLnEv+Xrm0voWPfi3EUoLoD54A
qM6VcL7xoGqAlTdSn6KxDXFfhf8Iuj5ESnd7IfZhUOwuEOy3Spv97ZLF+e4N
8EncogeCSbQ+zmcUlH7mUOid7XSh0TE1NvQS/MPjrkZguBsrR50vxWIxQpuR
mzV5Dn7kqjdaq5G/X98ZPfYjSbL2v7Kc2VpvTES/iO2WTPp6k7Mpm9TBFNWh
88SM0oZ2TCIryullg/rcwRPIPHaDZlfGftqvXmLc/oFdGEl4opbHdA8TAcqZ
VbSdk+KXp92iE3tCLBbOsmkkeS5zuqsQzWqJlOKfev84FZ8DuOyzPX/fXv3m
3evtFxBNVekxEDFxr2RGaxBWfYN07O5qTyxwQY/mCAG7v1TCPE1ASb7tZuLN
27UzsvWeCyVM2LWm4AtDIlSD3KX5o2saSokGaq/yw6DLFaRp0YiYj9WlZExL
ne9p9RMb5Gg7pJTuCtSMOk5Baz2zT3SBOP/13k7kdH1chyVPZ16c5Nnl+otj
UBch6v3Tf9S3QMM+WlK2WD6GkzgYqkBlYUDOq+Z1bOSxo9LgHf0AKCTqzOid
4ITbIjIRe6aci4d+1l0SlbdKvHhnasCa7Qs4nImSQoq6VRZvrl7rthnjlPbB
qt2EsMp9T8YjL1R9Dxm2XYLgskultAjKE469kZhWMw9TPlj6ZFJ4/8QS8wxF
R3yOO6ZrmafKb3KjEci9PC8cHCxB3U81RCtelqlCJg7kK6VzyhFgTFup2+61
ivdOsGFzA72brqEXnvW8qQNKQlkcApDatyf+CKrFcwClME753cgq8JhxiExn
/P7YUrDL8YsCMAi/RVxv6RQjYAX7QylqUq2Y59Z1ARRMIB9XimFbONuM+vdz
a33c2tzEb97EFZ9rEElQ4VaQoWowVO4YIgh34mvPc4RgQ3PBYyqv2KOX8YGT
AxECN3g9UF82LvOjoV9O46+18HsZf28KJPmsSpQVB3028wQMKXZbggFs9y15
fuvwBxoUaQ8KlrbwPYE0eoaP4Ulw1k9wKictli8mYjolQnWgi9Hj/zYVYIL7
zYe9e7a2v1SThn2pYngIhdrs+L7gPKGxawizV+53mqXygTLOh+5SLGsZLUQb
Kw6qD/86zaldbgJ+R42Klizou9Q9vo9cNLxro0kCBcyppnM8uFeu/QgfQFzK
D/J2EmLXT+utaNykyS9Lo1WMIx0zsnNRL5rkpLfOqj0Ft8N3JeV/HQVam4gu
F2CFE5p0c4AMdh3mLurlgCX/azESMsRIxxVxsv2O8QJfLMJI6I/c4FYSIerj
ntO0AXwnfwMOE9ZyhE0kxxheAxIkn9K7qifLr3Yb3Fb9/uvR7xfUrxH8eQR4
hK84lG92BDLKKOu5bQzpaepb3wUM16cGQS0QKxFBXvD0bcaroZYcstjFCCMp
bxBsYxDv1qixQNhz7xgOKq/yn7i2R6V6O/3IOib3otOFER1hCxm0PAYHkmMA
BjFcJ/YiHvJW8q0PRv5eWrNh5Sx8Z4NF8Pj0hBAH26JqoHJ0nf9BxgCRKp3h
vOEaEnOatTXrEsOUn4mIjPHci1nHuDFHjdd7j70JBvDOi8+MkeEuR+Ns0EK/
G211mkD/SRRlX9WS0PcywF+7ydeBJCjNgp6eDJFlcgEwST5B2G3Y/r0FwNVn
4gW8dvGqiNm34Od+LIR5dgMVLB5jz53Jl3gyZHFBfXNTpnxGjtP8fX3snSgW
nTDvLjagbS4MBIM9HQ/gtRQvdLT8sLwU1oAS202Fuz1xQmxknIgVA+9E9fCC
ktKv5u07bZwPFcVT9VXovlrrO5Ec3gz9Atms131h/fexn3iN0085xsacELUN
8ro7E5SI7+vBI3zTOSy2v7ruredvsy3BxqNT2ImAymiYYl7lwRcXxvzPDKo1
pwufnqmfyQ9InAF2TpMf57Q18Jizn/G697gsjUPLh6IEdmLnTpkhcpbzIW2j
ZvV15Fmf/VjBl5on7z5pvcnU2q0jDnHPxcv8XX8CobApXXs40rKyVtvThIXC
MuGe9c839fx6ykdsqrJVFKjucKqtDLH54kt7ox7UyWN2s3kgmM+Mdq1kx9nA
2ogIJCwCinsFJwWZ+ga2Xizlav/DG4QyOajdvzeyXSrv5E3Kfkz3J75eIEu1
EHN0TerPUZRBZP5z7ZuyyqmGj9JUUOIH9grrr29UWxsX/GBGG7RPSE6knjtA
1uAXeeceiuIQJ0SD6G7h6Mxx2s+BjD1frOfa/K/lFxUxOJqA/2mCCz7RnQ1B
DTbVLzP5tKD6w+nUBVednAV5iKZR7ZBPUIFOKxKJL5AVhR2mQm+9G6wh3cAZ
LH1GHrI3Cg14D4c6vccXWz/5ojKMMxfIi6AV9CZ9KAoTPyKVWTy2GhNzyLja
uTq/+b9jGez4dhqUwTbP3gKTNTx47V+3AfJs13HElrE5K4qZ/EXgMjLR3OUP
iPG97ENcMfMo1GfY68vSf4m0P52rzX5hRgBvn3mQ4//q1g+hSvUGokE/eCCB
c5lNyHcXpsRxWisvedW9OD3amb+EOW66Mx9PnMvR/il7I0QU6D6dYvBQ+H0V
o4ZB6RmUzJKOnw9R7/9GTIbSzUq5d+6q2verUQZyKsnrc+YK5otDn6wj85Am
nOS/DrrG+1oSbc6aqozMFFRK4gjOS5wU+Jg3DLZVX+I6qsErWq8uD8Bi/S22
v/LzMl+8x3qyca0xUfJyd6eshFW+Dz+hY00NbKMu6GmYqhmnfDa0zc8YE5jd
H5tQG+/inaHIRfYh/9O8ShxJdgMvOZdxx83OMyUa5bx+9ii8puICdD3GiRIR
A15W4OqyDP3nIcF5gPwyaYAZ6M6CC6PRVx4MdyA9ZB9iZ52XIan01T9FTM4H
A8LvGWKmfCEhNRv6u+KFDx7HCfRNoXvrKBBRY0LwGCwZB+CQO0BXsmpd8Ncj
s14OVxNP0x6dTKUjju7M7mP10wk8vIYscs3WtYjbZum7d/aF9ZKv6+ljYN36
6jrlIpzEAdOb61awu0n+ixBe9e4k1LA1FKuXADBDwDFeZfn74LnO7dTfOEdp
R6f1e001Ps7ExO9a8zDckwlIOUycFLFZPQJ93xbE9WMs77C9BqPKRgtzkDU/
MYAazrpDvhEgneLBkf4egLzgAIYCjAO+428r48SItmdN4IVyeH3rwAP3liAj
SH6Q3tmqGEFFi4TK791ml7MNn1PK5B3d70zIduVwQqTgM2xOGVI0KcPmkEx1
6ykRmYruXj9/1NIvDRXEpAgpq38IP1i4XyLgG4pjom9PhIbO0w51he6e9W21
h91t44p54emyOJ0wUB9yK0Vt6+Hpqc9EI42WNm4LNtSNa22FSV9M+6viYMYb
wJl6XxCf0XIIOR3/tySqJ4y9UkqeyP3nBIuzKIUJyJsW5yEl/k/bueA9Ptj8
m8Tc35MRQBCpR2gDo0u6LzmQ8S0BJUsHlEOWZxM5u3gFvpvkknj5FKfXStG3
GAPSY3fY+DMppmkRHQqEkB8Rkl6LWI7XNMstOKhZNZDV32kZnzZOALy4NxR6
MydbMcdmlQDvRqq0EN2n5fVQv2wx3dieE9vfD2US41/glTpssngdO9EA4Dix
LY17qmLaEuaISoCI5QOrTqY9qyZlOXG1ZJZ7rIoYka7S7ZofAUCf4D7fWuOH
1VdMnnYr78niERTxihq19UH+yvkJrSrUXr3Aj8tz22l3s7RkcXPyMjC86Hp2
E87CHAeAOoQz6nLWoH9C5fWOXwnaKxdBgF3C9i3uxRMXOti6yMrnUvAcUNq8
oV7hCJDUNgFTGI95JfGi7d/I43Tjvrg4046ujNK5vh9L5CUrVJjVDHeop48D
UA8aS+ZGGf9eErZD9IoV0mcvXXIUTGXuFY7mTP1THNOat75/yL44lBJxb/9l
gzMUm/xoB/KzUV+JLtzK5Ey+WbGPRXTgBNQALzIL5YU2ekQNB/cNvfkNAEmO
BBWBVFLPVXAXWwqNlxSSsJzZ2DTaP4/+bl0NJ4pNnBMgLAaQSa4SYxhxDtDV
/PR8uVJlLzT59zCQOUYUCKH7hGcw3/o+Jx50bNzWJYHIs/5NjhBr540QxpwR
9k/NBUt5hvxOb5UYB++CWvYIctoTRiKCJAiVuFiPOkfN4PLs1E/2gRv5yoS3
WGVvaHy1WKuzd56PuxPf8/FSDvYCzRJ2+u3I/0MMWrmY5RjZrfqM2Z09PRNM
EmiUCtcki1ewMoO9T5XevbqvAX3rBT5qRtbYhlImZaiY5Cnl3vmKy3/+yiLH
whbHX5zrodsvjluVMyVP+rHNf/t40lf0qZGzoAJnHgfH1OQTycCcZDQjeTLu
kWc8tlv/dflrkPiEXf5hNDOmnZq9ym0cnP+p03MGXqXhjbtwLosMGwAYK+K0
tAOLgdRv6AQDz3gUoZs9JMVtjRfwFgw3+rRAEsTW0ESgYQS7Dm5fb4Idbws4
hGz3pX/xIyQuevNjz4zZDC+1z75HwS63So1WUbJ7NDycy+MDAjSDaEPG0p4N
VNn8c+94wo3057DiagPVrjFJtPaVCZX9u4IWSsl+2wreno5yMRLpXRp/FXNe
OpS6S13hepOZFaCYfcWSdJJyb0paVO8fUM3idzSAVwwt4wokXiVrThdc6mes
Erakda+ZgnhKVuxXXJpYqFNvrNSMyYl5ggfszLAaGOJCvoZ/DLs24ZB8+jOd
D0qQGAysW5I4Gln0GPQH6h+4mDzdRjZ3X/glVk1ceXRHs3CxT05GdpZHJk8O
HGiJTkFvoLRL+DSWMu90DvG649vVB6CcxyE2ufi2E8t4k/0fsCKj9muW+819
zkDKn/wtLZy5eYZkNsZlKjdNXk4OKegw3W6wD6rOSJL7sHR2Z7TkLfHuK1M6
9KDdGfblbu4aistgGbQ/o5A9uKDjw/Etu4YTE2i8ArC06b9RLhYP6j38oUf5
SFc8xNu//LIiK3CRE4oCDXrUQKbDk2Kgph65VQUgMTYiqv39WC9Xy9TnuMKZ
YL8+91lNS+R3U3oaTQqRPAfRjckUf1fvtODuXVhQaldYXJjhr/q/B96fV3rM
YZaIUl4LBWIW0m/2HMy0xBJ+sVjuqjuD8+s+TEnhRupn7J4pyeRdl9w7k+VS
1Q26wKdx446lSFZfu1f/DpAtaohJ44fysidTCdE5DOhf5+o8nzoHVv6LZubW
IgHyXhWb9H0ZQU090NBbJcYUeMhAIa5cVWwlBdpz67jxledy1hTGvpvdmywO
uzsY89dHHe2dCJgRoyPXIbFerbDA54dNmNkqEaSeukdgzk6YAa55/NhI3Wez
iDGinTal3d2/8QzVq8yjXIRwS2/SlbHAtrGSTsWb1uLZ+bWPmKSyYxJYdBYu
BSvceXAmjNY/CHDmqcitaYsnMmVmD83aTZjwnALDkiCO7m46OFeV0L1oG9Hl
gbGr4jNEzcXoQ1RF+YNeco0v9rrLFMCWJ9cTBEUb/S1G/U0RZ9CfOCDR51Xn
teRlZxm0GTz+Q4ayQqpKOGTyTMNibtaai7E+s1VHmDrEVdgQN7luZAOFuYjz
HQKyCGQF15+k87A/JrWC4clzdhZXw4XqGSxw1YO6M9RP4Q+SB/8sR4kbVDgE
FtNquKCKYDiRyKOtIKDffPESyZS9QH6+38PQMGjLN1PbZPIsK4kngZaFovzg
fhmq9JaztWBpt5vTNE2f5XfDaRxRpVr7PtNMRkn7RcoQE24ThnEK5P34OzFY
G94NoZfIcBlpRRg3eTt6u5PciEqwtkX38l9zg9vwQehXkUcGeXhhoVGJaeS2
n8c2bZawon0l3itGGM0liZ8ekE1jj1WnUWLwhLXVuHLrxa5bt8d4o5MsBivy
2Z3m3DwvKeoxeOHoE92LYyad3IodeWXOA0oMNC8p19twbSceiD/wD3zni04F
VRfW1eyi0MKqiaO7kZRfFWMj0ilbm4ilFmqtZ29rOH8e/MZLXFffU9/nh7Fh
o1kkifRKj/wrIYYWrvQizpMPs2K1ap+B9x7zBTJqvcKH5oOnVLBVqI7R+745
NbCECdY+B1lA5tqg9iJ2AuQO/L1K5xV6obN9qpx6Mm+B0U6QDR34xZsYjHPW
ies12l/150pltO5a4IctZpYOUXbQz0s2MKmGUzBGIUYZKWWcASX+9HgChGJD
zEdfUEAmR5M9+xxoo3r/1Cie8egPQ8Vzybo41WtmV8liNFYk3bMkyxDMXRF2
rqbQaE3MiEX0VcIp0eUS9udHsXLHKaeXEtiVg32eDd00Zyi3EFHUxH5q4I7Y
U7qV6NsiXHfKd9sfoNSf9aDxJ84rfe9eGbg+oOZOvOzEAEtlNzlCGsz/V2es
HIRqZBmSSK+YtjqSa1E/EYL0KDX6imEgZoHYwHWETwAszVFFPzenjatRYbji
2qSLxHfZuB7zNwfbTxPDm+toIpf43xNDUUQZZobg2POLaVAOpijsMyFsYIKz
CLAwBE7qTfjhgf/746jgorrU+ps2rRXr0Ryh7HT9j0bJf9rxmcmPZ8Oe8JJA
bNTnTLLMhQ8S7e7ekwzMgwM/j4ZwPDRnm6UCMgAumXsmzASYYuxCrhiPVNr/
1TtN7KJ15lFe0yaJVleGW9e/0+hRs21lbN+wMae5yEswcnAOse/gEFTE0Qx/
diKdfp2fp9X/82uY/vkhA7qBdcnVsb7pKra+z50TEXMwXVtkcd8JhsUNoA5U
H4khf6I+O+gCNsyt6a/MAY2YmTv4PVvS5ASic+m+ZxPWHa6Zi6oz84iqvh03
0AIs/0GpmDw+YnLOReVczhtX+zgrng9vPnd9263O/B/rUzWS4KhElMUSTiZf
VsAMYvyiro1pex/mVPsWBwhhFPYwozkRhdah39hWGyLTXxs7nsU9C+Bydrii
DCKO6m5BSOBKGWE+GOeH4w/8fqUlNaYcDnJOhX3dbeAdan4i+qXFnfNUQ7h7
UZmtnUEOy5cN98LUaVL67nva4LwOaqfJXy4eOgz3MAEZKRD18Pxh6gWvxPPV
XpvawWuGcuAAvs2ldrSK9FujNhzXpamkNNtau7O/cpH5ICiCBh9mqmBw85qk
z4iW66SuHemNtqNQ9oKzOIhI3+sQpkvHnpfvomfGNqUfFM9/cjh4a1acJ3nS
FardB0GKxPCPmNvWx7vDdIIQKzK0ObtxXlLyAjK4kmCXmT6PYwDxi36N6kOH
2IfHizzimZKAJgPaaYo5Ao8Trt6pM9MhHL5Cx2Iu95EI6Nd+VV7MtxhRRw42
q+1fmCM69N90HrY0uKUlov9kGcxsJPgBljVPcJyKr17rIaZmnugUM9ExvP/h
FTiPaTUOABkiWypLtgOpAjnEfBttY/T8kHybGYFPowD1er04Hew9TBSFMteW
/KhZnDlut68DQjOynNSBG5QzHuekL+ApMRyyQojxos6Qa1PB+MVM02qcDvyz
PAeY5ZuRFVwjFMR2uNayfsk+biEIqsaAsbd84KOifS/t80+WrvSHoeN+/qzD
/18xHsc/m4X5L3SFcnlLLb7qu7uWJGXmcogE27Y761l0qsaI6dm4GMLKr66R
d9cZ273QlkyxlGfAxuuisbeIVB8YTL8Bfd8p/wcrBnAW7oRwr8Khmm/I//+F
Pbo0UnDq7IQ0XuX1sKmJ+etJzz3PnYTNEXl4oQGD1WgElNdwED9KwQ8iZrXs
bFLJaoe7ZkihlWXPMmsf+wtQ3YK6p/hzpzX2Vv1KwUVU2WG7yxLMH1AVI22D
sNw+dsiUSu5zdZSu3svqN8T0yoqIwYASv0h3L5cWnOtcrWHsE3mj/Py3OrHB
7rlJzNLs4Rz67Bi9QTdHpO+vWMIYP11xwr7NdsokghbgVCRTTfRe/4iFZZbQ
BHI+ZpDZIkJvZmMwIdqiu9CQ4EDoRxBQWDWsuGPGZuG9SP+AFBeQ3+n+E4sP
VcLOEJf37qRyuXm+Nn0Uihf8aMT4F352c8qWHtGlmU1lzsA/V825ApT7wr+g
1yraj+SO0OKR6UTOvllsrkyT1bakIOxrOXAx106uDEHKVO7hTn76Wu9CQg4K
QQT06YJzwYgFPF/Qj+juhv0umjgixT814utrIBuNl33nBDh69buAoNAd6d+D
OY5S/dQE8L04cpCdpNyyklHqnRw9TXVaiIidesMfLbf9EYgaAjDYJdgkuq0g
9+2JxEA+QorMUaO7hA7umZvQBwYt4mIaEsm//MtI7Y2mKmQ3LrAXth1X4QZR
4EQm5XGo5RS8aIigpoJVhcN3lE+VADxXt0fPxUXiN14MR2y8P9gSckRv9MeU
XByLqe90QjiCxiLaZe2CCi6jQa3Pbep0ezuJ7fztuc5GNd9r53MnIyEqXg2C
p83BLTwLFe1H+e6kRzaPTJ9ECqotSxErw4zX1G8Z7mbPB2KRWuLAQJ14Xol8
i1QKquLHJlEwFGCfQbWpaI3am43xlfrnB+MqMnuv87GT3XKmPWohhgFsn9nl
UuGJK661phbkFMQYK/nCc7JJ8QCnAlJUg6wpkMX5wtzx9lW7Q6D7gfX3wuSt
QAgrW/PGhAgEIAXr6cYHYSQD2s8dJ97v0axtOdIRG101dVatdtz9IZ6i46f7
XZfHsFx4MEH/LINMB3sBN7Bg6ocOGKX39HEtt+aUtE77xG2Z132v8v9QStk7
pO/K6w0xtuXEtCqX7S5MZAp6EG8mLsGr9PdVNUql3E0lFxgLKy0Ck1PwfvAt
oOXn+7wR7302tcMbeB/wtpbJSEl4ZqVmOgA7jJ+bES8hLx17d/Cwbs7bUDc7
bj9EIK4HTelyXv9EHPgXOZJDqg+CUYoaHL8fH2iARgL1eYdNv3QNb1RCXYXy
/UkA7J5GhXno+tEBKwiWw+cXB7+A/ZYS8plhZcJmxM7eF0lEaOR5BT6bnFNr
z+EvMg15nAWvc3rAHSh9QMUgbrbS5S1JsFxjSBgCgBUIjAwLnkJJ9pVphQEl
Sd3w2fFWpId9WuohQ0hBacPeLEKyje4aqKxZ566M3+Y6T0Xt7iuSq1Pndwix
MPO5qsjgxReN1FqOrUj86f5Haf1Pu8ZvvHkrhl7oiYoYrzBq263Fm3t2vRL+
nNWV8Vw5whpshyr/UM3ZB8uUL1iaI4WpxdJ+1+BYkuw0WbirV9AiaDL0m+ya
yR7wgEMsqZP/rHJQkxlgO01pRyGxvAANRGl+aS76/7L4NomKHXN9c0r9CsqC
7sWuomI6LoTOREjxnPR3kn2ujyVRV6U0t7AQSSMpMo7Ru/yNd5B9EKslNn8i
/QIIPFAok3ku+MnviZMsfc5hyJz3VFTrcUnlsRqEmtMvuB2NeuHBpaC48qGv
k/nbYetY+wiVi0ZuJ1aTUSCBjGSSWlTLfMsexP7pt76I3hW+LoKipnc/wgK3
zteLByQoQlAL+Nr9xI/m0GyYBAx+O5+p+aTm1N9+bOoX7mEHeyEyy+8j0QsI
psZ3fS7emA7U26VSy2svV2E9BhU+RoU+NKLwR1lJ1+rrMHjKAhQaR9eqNi33
u48Wc/W1elaBplyKSAcs4hDfZG9bLS2jgh5UmpiD4E4NIva6T9+lNyIVOCp1
Cki5FRh2AnuO5wHszpF/iW1KxOArRKHXzh8GvfUs9rRGHZ9zMV7SPdwqwwSU
d+VZGvavoG9RurrWSEJPkOHjbqz1tTu5Ax3+BGa/p2W3rb4VFv+ZMK5VV1nx
3DcpIWcRdV5BlKcxFVM+jVW9OlHKIv4TMfKaYZTSo/xLiyTV5+RJCx+UoIjF
CektVOv5LyE+Tf0P+weLPVbGh0GvBIMazkQ97Pf02RtkDLFOgWB/d6D5PIiK
ebGEXFNRGgdrzeQJhCC3NHT2vXm9kLEAEGBQByP8zEWOLcU7xwUxgkSgwM8B
425MfOcPAEsEftzKw+1bLUM9DDF7CnsmaRS3DK2AWVd8nRFfkjK/hHOsdpgA
uNcdPDlq4O/eXS+hnUH7l0oO12aJU2G/e4c2DrRKFKOWj/oX9iwO8k9AxkL0
Lb03du4UJHjsiY8pGtc74Bp1Iwc09Gs05iV+Er0ykP043v40jfdDdwJtRpHb
Ot2Pi6EWf2Y6QPDkl+XAdx7tMYc83ZQW848Rg7W0rxyrdkYkBbKu20eoUrwS
y7fXvOpZ2r+j8ksS9z420l6I8itO7e2moK3wuACsnU+7E323jQFik+n0qTQS
BZtRbmyN7OKWMQMRrOie6fpDID28GVKHmezi/fafnINdGVduUuigltc1dI+G
VTiXldrRQEx3fYkiydVwzKOVHy6G9aZTLVoFwUzy6S4vdXGV5zs4yYIU40kZ
7w4QTvOKIoR3vK/d4Q8HOOjTjN+ttNUoXTlZa+T234SWj4ZUQ5ejc6u9hrh0
mKBT5yrCXA9smzm5muhw7Q9evBdz8sQs21JYoPv5TF8wIbxuI7IMgvxxyw/1
1JwfZIXq12KDhPZBBsRCCFDOq2fGyuLwL3ReNuRj2fdEVpd/cpN0oztLOSt5
UEjXVfWljseSS2euFFVUR4J2Izd9T88w4qxMpNNwNFxsALe8PtKZfnAVugqP
Oxgdwn0k94bvVQ+t/nvUlUoAiKa0QdmakGqTdh4xW/Kkck4m9h71CAYyOox/
jeW2lnEYwFuRl8Mu+wcrkvvbLZ2aABNDUXgLxXLOMBTxMA9JdHwRvtYxo+zr
REL2gRwyIL6EgPuE/oqbAiSyyoIln13kMKw8cAQS6A5RpWBj7pUWiLzn/+aQ
t2/KtxSAoNHCWYPUOb4vaD8tD48xt3UEMwpp3fLPekJja40/cKGEd7cXOTM4
did1IlLNmLbubZOHdigmIlrT59jUsJeze7hEas8nieXcyXj+xI1vxtMC5x6B
WnP1Kaag+SsLclPilA4fInfLMwQOkc9TtQWs+YyziNsLQ9x5LUBwlex9yD4i
XSIoPynxpBKJwAdz7jiPzLKtim8xfTgP1mQM4Ah12oZHcD+LpOKm8N6to7IM
Ga0Kj/z03Sb9hnHfAAlq1zyFCJhzu655EZuzLeh4Pq8ZVz5FIKP0VxVGdf6j
cpbCVQCF+AXWuiDleS69osZYQV5kkfZ3cqhcYXeGLWzrMC8aM7HZmIgV/rzg
qSaPmKd7b8L34KOUAH7sXySROrIdhdsjpJzyDb635+f3bg61BsimdV28V6Ym
CX9qQ8l2/ImfXl/vprNYtc95mxP+Tg9n5vgUIgt7ISfcITqch8pjjJ5Hzci/
CVkqyiiHPTdtechNybsLzV3JyhLVVwK3rO24eqLh/HGG+kEtjbZN47da3OoG
rr23iF7aKgdANNh9RjOBF8jerosPvel6p19MeJc2/3HHu8fIRYhQ6L6bDtKn
3jsjHnWn5PQP81ocWGdQsZetoSSgT9KypIafjrSayxDPD+5UYSmbmu4DLFX/
jDkn+HVz5BexZ0LZhtVkXVXeCyZ/SEfxYJDQ40MfalgwJmWZsEDMHzL+Xo8s
0MgUgZAtc1fK/fVhdAGpleRvlOlqUea+VocFIjwzKEuHRCCeFHkZcveu0oyJ
bWbTDLt0FB93Ttvlue8s93TWTMmrORNxNHj0Mbnr2tKzqlg+EZ+jvet3gslj
mYt5v5BleHSjtSoPujwY8cBM3ZbfvMedq3Do930LGnh0aiKlFRMF+f0yyunY
OrZ0bv3VG27/FL4iWBPLocYLUINmPT7FRNyOlT+pNW/T2jxxDG6Ijq8q8dBu
VP8UXdG2ww4rVhknSqpnwRZQ9Effl0yBMuRmb1YRzKXQSX+6Xmb9AIcKgu7P
WIjJYSl+6y5H52q4AahjcRtUq9VmJQwzsJ0eL3jO466cwwkLi+bSaogvZyVl
Cbq6uRSAZqts9hYSA/ih4u/mYrg0ZmODqkOSM0gXvhsV97j1uaTj1Cgd96ZF
skQ46/q9W3Q/UMM8xhRsp4I9risWZmDm0BbazsgsDeuKxnDN5Ayzcxq1TOoR
HXQDDqdhJahK/Lq58As82z0o7gMz8lIHMPcDI+ZPBNJM3TZNxj/c/SqqeKko
DYaMAeP/vPkU9FhtyHysvUPYsdycnmvX02KzRFFYegQEN2EvjJNAZmmr4nTu
mlC1TzJh6oHC4QekQSL6IjFyzTsj7Gc3AlwpWgC8gdfhLFa/Nqn7dkw8w4hq
cJqmO6kWHeIDoySmpgRCnWuySpXqXvZPVqrBUe9ycJ7tkVzkPRY3xMF3L793
Gv2ltQNC7Oq8sruHniVaPR9gLZTEEOEt3vDsdYwXMyMy/MjGoA56ynPilrdG
WFSbvqrdyI5/KQLzpaOrj7N6eZYyjodIU0itmBBFWSlW3OnRiOBKlk2YZxBM
T8dYKaZemGDVqHJgF2R3xFlxXgy/cMZwfZ7aK3ux5f4IkVsJm4Nv5hr5c9nY
k3DE/HJz9/7aXBKq31wrDMSk5cUAPXimBTOqAhFLhJDZ0Mld2sj4eb28ZjZL
oAUsj/YJYUywvDWV0Ul5TdXRJxN9awYYc8aHV+2P3rZ49YUHwPQ/lHtxeUv4
q8wGoU6bE+jOifMCBm/hMqGNANlZ6WRnN38Y+thrTxlWgyWJg2w/wuWPqPOx
XUwBDDXkEmSIQ9/wMdH0YcB8EVzvL+fQGLnbNF9rZf7UgZWdu3DnKRQ1hvf2
xR9yAmtl75xLA+Jx/EjapU3mdVWbjmDKr3Qqt+L97V/bE8GwEC15KQEx2eE7
MSO+XhjaucGBKVr4JTwuhPHRr9RMHnB2BgCA9flWN/ITKsFBH4l2azqGRvSb
e/HxddgrHu3qPFyDFrze/X6kvgnpuE94x0EoNl6eTe18JDVoTHNdgK/SwLsT
2ciQ5DHB3kj/pCA9bja10LNTqn80/l7B4M5J4zHdAW2NpKmWHlJ6HOaS4sLa
AEtUW94i7ULQ8ddriinc6fgCWf9rhwt1dxjLNoEoN9mFXAqFZrzPzzNDGbmm
Z2A5M/OVQRBmPyo2WuqK9sJJ4uqsYC3BthSpzDswRV1HJfMzr1XUlbycbXsJ
XB8h4U3x98fWuzyFKfUyGbz3laDSUBgzhdAJoB58QMn6U+a6d/hjhqkd3/We
MTWP8c1kmAG5o1VmAkahdtK2vTMWiDBPFw5B61Gr4x+H509QWjm52/5srKr8
1J9OpGFpFw93Z8qUEqIzDbD7lwxpCU4P7NL/Ym1+Qcuv4HrP5KQGOR0yFVUP
9N59FwPfKX5VX0WMySfkdbEALKJSyr+5PL5YFUe+W7qZ51XD4YCxhc6ZVCyg
dRp6pmR3ZYrDBdiUMeEdvYCAkJxwoaMBydE2MxLNOh+gIYSmWokirZ7D34VJ
KqGVzrEShoGWqL1TR0qN9SHPXwg+uVkgX6v0MRQLog8S+mfeSps+CiUoTg2c
hkbyCWQFHOakV8osePtaOEaCZQAJSYl8DM6ycQT0ZOInWdVJxG2cNxbe/Glz
dSISxB6G0NaT+cc2qoKBs/aPpaO2doJagbm8DZo6YggaXi4RLRz5msFropZP
36QaRYfCi0h+iyauVLu8FwFZG3f6Rh3ohtNSsyz4bxV22LtpFzpOCSv78Eat
FkK38cArW+LCEW9QBAdwSHZszBs0FKiEUp5NbydfcreORUTeADt3n7VMZ0Y/
4L9VE6IJ5CH/PwhMCVJwkvnsPBf/avFSrmBphcKlFdczshgsGzEJ+39BIn7W
L8li1welRFGO+ZloQ5EP3gpITEBoaBb3sL7sQxq4ea8jKsnJkZ99LtAqlzMK
zVLA6PbifKlI+IXwE3IdgFFSQ7PRTn/OnwKO8gyYRmAFJVoaeyTq6BLg/9EK
qcANdmTbs4sGXaerH03zcIJHbiLxvLkI+GbZx0KbP+P1Dupm7NYFgLN7TxlO
SAuapXO8dn2mCl6K6U6YFJYdcPZLngJFyCahqMcayvS+NJpsq8dULX2IPNI5
o1RxOTGZ35Mmrw95OqD7f/UKUpdTebu23qkiboRgX/cq749cWvBI2V9eUwWw
vtcbDRU+3skz9zw7DhuEZpBaJd6XEYmaeYNgJvu5hwnBcG6FBf4gKQcyATfL
UwBGgR67rXNcGY5vrlVwOZTHMCqCW4QBicx8qvFQGePlWFGFgx7GTXZYSfx1
775sn/p6WPU3+hAdvWMDYF4LmIF9foHIzGr/xn96xZy2j1b6n7XW9TJ/sWJg
yVEHepJSg9Lf+E0UzOl75vy2thi2z/rJxiY2rxichNPJWFsIAHtEK7WlwIGx
MG3VP7BdOwWqofvDA/udBIeKf4rxA4iQACPqfAXzgnORAMOeO6A4D97bZeUk
rg/CrjAFcVuFVJhx537jWEgH6ezvIdDJOVNIvPhxX+8SgzLyzRTMP6t7jdNI
QyJz6Kmtv8M28MwZWIb5ttxUqtcWU2w73HdR2leTYvt1eJL56qSByyfTuRcn
aeQ4iY17kquXBI8xFDgPU7mwLwBh4K7Dfz0V2n0M3wUsjqEab8ccY/aD4PT/
h7wyvEwP0mxa6VE7Het27pVqSleaBya9EQ9m9l0mwW7xgoeelveG02iTsngU
3eqWRjmv0dBMb6vXz40/k4AYgnQOh6U3jJgJzJrjPEYVSiH9FgegcJJ/Liom
VHOWT3/YCB6v0qTU5JQpr4SMcDEC+1K6viJb31Ob/BtIQsb5X7g3G7w2CHWz
xWJhVF27sux3J17qDOkqC7zZU85zb3H+DDgRvhU6lmU5VriPuRlDMgFUQx/9
b9wgvwDNjIOwmyokwsjV2m5AGf9cMCHTDIs+WXKzQ1gEOxoH4w478tWaqor3
uzJB4NIBkFwJld0n0dHhgDyJIHfofF7OSi4hrOuT0yHcW/QCxKQFuJ/GWGPd
vjTW53FLjv286Fk2DWPe2n9rJ73Qy/8BnZZ7snKTG4B30DZG0NoLOPYPX/wQ
e+2FdRkdDJiTOtcpZrw5Tk+83G/HRauBx59G10qIHF2QCww1Yb/AydYdWhx0
6oCPHFWD4owwxm8X3DqoTwbeOUjq019iDX89VKFMRQIWViJylaYcAlusOXUR
PH9tEwo+Hbx7SntjKcWvjGZSqcozAKoHiWlI5SrQNjDU6ce3q3KJoVrGsc5v
9zh8qryhAWvxpqvckbTaspiaqr9Pet07tT3DuKPDtvsqB/v5QqVgvVJBtZCV
xGbK9Q07oMv/1PGofcOB46kSOsBUhHM63zAJR549HzMB7rjmtR27mK386ZfD
1fQC3eLQbfpmIRTCEVKBNppPlvFiG0jWa1Q8zi/Alk+4yYOLa+xI8Ldy4Nqj
bcF2uAoJKWDepBRtKcO6wMEjmhf6wB3IGIZAdiR/lJ8Ye7butzOBX9NK0env
83f9+CFxD6Ggf2CJZpt+HwkK2OJ75PEhndjUw788jQNwjkmLAWYoiNxUH4A+
Gs6+Y9t6cxTrS6ntdEgdqGZ6HKeW2b4pnYJnynkXLzbd3pm7eBcW8/DwAvD6
M1D7ljbArqr3MrYulQ6uuaBTFUSdBu20Omh8A7mPmh8+nlEUcsbsBWmtjnjE
YP5TZeYvGxjKwylbHpPLqevAdyuagENc0EtEGPkZokrfA2qkCnbgap7DOm/M
KMf1wX9RjR9ZG8bfDFCp1rZr/QOk0H6XJ5CzrX13Ylk96f7HhWmcBsaOFu69
G3e56jr6d9MNqjUO4qgC74d8mxiP0hR7MSaKiDQGPw/hNEVhulP+LvN4r7ND
t9fHkx0vDlROt4UbGVLfkbUCAZ0YhTHX3YgEgH79OkAgp6sn93CfdBjXPmOK
pIUIytqC/2uw8DAO/3BKma3+QeUFLNn4HNrXVJNv1IyQkcmaLpYHN+/iWIkU
JiE1X4rliVOh9Zzys+FMeqzCuRox3zdeFxCAx/xBRCJAqunw++/itY0rTbkK
v/6awgysxXYK3GQB4tdVNWdCLodbBTI4uT2A8y0NhoIKHqITmBfkBuw9qvSB
6A3h8LqfsOvvqYVTzizR5AbemrmEUJpZJm7EWtec4fGrOAV+l/LeS9e2FzF2
hGmgNuQ9RvcH5cERoS3xcb0SzPKGqHgi/p3bqIPLGH1zR/IF6roOIWPNR9lI
ovezv2//GTocXTJnSepzucQ+lJ1CcSiExb+F3DBBidYacQMuoQQBTxh1Y4S0
Iq/YGOjsv3OyEFzP3Jcj37/3h47S/RVSZrVTR1pcUjr9KPsui0w5/8CTOs4u
aOpg1MwTAqxfKxOrJazGEdYBEAwHAKugJvFDSERCMZPy0EyjlMDLzZO3lKNp
s7AKFrEKAQvuO78pj49BOxNJl2U8SWomAdjP2VAYM0ozlp1nBFQFhaAbjImg
/q04ZvcS0RvjtMbZLl3Nq/jGcRTYBXQjCuL9qgVI87+xoCdmdVD7KdGlq3mO
9ZYZ/Fr7DHQLxZp+0P6lskePahWH9HYQGhsrnsYkZiqHyAF8SLxJjBfACw7F
ykvtRHpOXbiFBapiHB5yUNoHN6XFMPmFEX0a9wIgYsPbJVDiOQYc93h0ARP2
plS2JZAAkV/3KdgjkNdKcT9oOPmYe5C5pISawLr0mg+keK1FItZaZBHJKqcm
G4++eJhr3ff9BRXoAsdJSIGwVb9qIa4GczkbQSa4DeQPPGTvi5SW0C6L+9R1
81PfyUKCf202rRGkt05Uble1NnjThuMR7ZiZRcHpOi/oYwY+/Kw08Od+YX6c
zIuTkylFeZvz4nJAW/XduL36JWLRMWR4CRpHr5P/CBztB9WORMTZSmQuMEfp
2PrYTCMh5c8fY6fuNEjCjLS94v3RaibJv1q1EfuTKOOH+yYuyB/+YfMFn1c7
W3FNswXDtrWJ2lobbPuj60zKD3Lmt0Huo9U0EFtSKJxQg7wI/tJ/VQdLorwN
uheC6nN1PoR85r+wbkTRUiEie+jOJmcrL+VqL+Q3kjQ/3LrgleP46yIH4Q4T
MGFA7KE4PI2Vhbb4RRXCsKBvL5dZ2MhhV/PBB6GUu3xswnFuJcD8i1CL39Ar
6eg8eLWFL5nPzCEWAhgliUrcNbvPE6CXq/pgjHCJcxnaLJ9Kn4OsMVNXXokg
Hltr1VNNpRCApRDSNO/BJ7Q9MnWa+1vUw5Ipc8D4BYgUgwEByS+tILF7Wm1B
vqrmKTVB2qAdZhqXCQDc1bfJCW2rKZobVyUIozf1D+iv9alLXtb8yUbrwPDn
0ISB58Fb/8ieh4nEgTeDe4hvGBpHrE+moGFGbhomo2Vo3SaPXuHJAnuLYTIM
d10eLauKzVPychjVsaC9P800jx3rQVSenEdGJx8I/LUWgekUvBFqdsN1inSM
yvoE6WtK2fAyi6YDRySfwHKgAJcfsm3sUpbXVy9pl8bVX8ffvFbBNTTrbI0M
NxJwEURitopwbFY/E68Iy2u9zWABR5DjWjNuBrx3ay1AY9naNn5yHY8lRCS3
htXh1m7MU0TvBRBdhEpG2zxsVic7Fo9yaYSxJsSX1JQWYZDBap8LzC1yvp82
RR/1HN6bt8R3IYjr8eWMQJeGARijzn5gga8j0nWZyQRQl1Gsg3w4iWNjRi7X
BqrnQ2iFRdiYhD0Qv7+AeEDtyHBnzqiAcT61/q195VGqeJAEiEd/zDCQNGaT
0IJUf4QdfWUJfVoLkDCMywJVGDuv7w9ZFNHQ9SeJcnQ4LabEbA86jgYRTbDG
JTz7L/V7ybc+82dBgWgnpc5s34Giy1rI8cHdIrQknzTMYxO/3S4+v+IDrqCX
zY9lP0nV+bSNjaO+LHDk1EORZhqQX+x70YsXSWTUu+iltnrorvCwkuUO74R3
S6wJeajPMB7N58emoEwH1Y57NOncEzCTDK0aVa+iv1aukhysxWttHg3vVEFr
agqX43PQMksvx/GIS3ILcwW7peyw/Egb23tKJ9gXWu12uVuhimWvTT5sAtzn
mn6+EBKLFbDOSaeE+esRBFnDd+kDHKLxWRNHwbUKzrV31J+oFpYDmZe69xXq
t6GZJMmb28TpApLaX5FQNNRsr1HLmseHItxH4SSngoOg+H3qB5bOu+TYlT1t
+GAcF6OVVbCt2sRJe+MDTNd7uFMRlc5zp6v8+SOZB88QnsUxmf5RwQp+WsI3
4EIWULnWE+Ws9yuA3XcPZP1rwLPOHN8LgWbIivQmJhKrUljAqzkJ7NSext+e
klOZZnYkdmNMZNzBxXLbRzPYu6HTl3XdydjQIay1OmwOe6eA6Bs7sVpcUUaz
4s/0ibbmPn1O1MZwyie4U2OzvVNOgm757qIqXP3xGrObuZCd5e6Nl03v4/yJ
zarzycAQloJDEl+KT/mOjhb0deH5JqphIaIY0d/7kBQr8uxZlN1LWT4v1fho
UmRuq9h0txY9zXJ9vGWfkTCQp+YFgysbWTXUa7D527zonHG3ATcaloKaQOjp
RM+MncullxKeTjNTnuRaMVgon0AYzb2FClXYKHJO1TQg/jZTraZewvQLI0vk
K7l9nkGKexJo1jXMOCC2oq7kenecl1cDEqI7kuLZzoecgl62pIKHzvzon5Q2
Xpo/sNmzDZHK0d5msmE7m2021OfLun1H6OehPDemTNeN4ElhfIl1ag5zgfsi
IbPj7fi43+JM2EXjQO2PAhUU+l50mrfb+799/n3FmUkTgds3S+f7XKPyqGCs
b0HLklwwyB+n2gjHwHWq0TMpxlih62tXhGjvFCLPtHlwxrJktVXi/+A0jmq/
6MJ3wmaMmsMzCjNzlI7VsqhMxuXahsKKAk5+YugO9EGaxVIRwRHwI9Wc3T9f
tNkD3svokrWoZOLg1g5hGA4pyRbgcKIeldFCswRk8qI7y7DBzNXFrMfSLEsH
1x8L6QfYubEAZ9Q6ixd/+t92fmtRZvkQIEIIyIQN3CUZBr3sIZc4kyAD5IwW
CLYvKrb1Mqu9iayo/hi7UldIxBg/O8IL+rHGGtk0NKoScA3kJ4RUrTNafzrh
nEegTOO1oPmfGiHzDJSc1v7NhtKVld9DH/zV06PGtHRIr3dj5sEQNkXW5FRo
1PPPq1Lbq8/ehITF2Lu80FJiKGuG1S50ztd6xe1jyGzw3zAiAmgKFqGD5GLa
N6zhWcawQoeLtIWZfr7u5uH8WBTDz7ZUL2U2Mh6gRSpQznfplvxHK2gNnYu+
DFisU1s2PPfjoYtt/RFP8OGopz7ekiYw6IeyZsZKBUYUwPWW3/aTpmv2V90O
Ye0yJ23+4QgSrpV72MVwDbFRTgaypFZBwllRWw3UQykKldRTg0Ar81k5W8mz
+gmEIw5LV623NdGuCovzrXQsK/FkBPrJ15nN3Z9BzOarigQJEbYU99f7ctlA
DIIasRskRT8GODdwI1a6zkqdy9Rr6DffsJmr2nOZ4svrTqkiqht10+IdjvlL
kY+4O5E4cjzfExyn813vbudnIs3HLs/8uQo4xM+6GUWs6hO8ocVSNxCYmdbP
Zg5kbGNNsJz66icsMuuiDvoGxjvqcJFrRqVIKupl/SFMszft78GhPr69AaTM
NohQcUXbDSUr4PRzUBnR+A3WxVu6AixQQkvLNDx3oPFisWlUW/6xTA0blKVC
R6G2oI+D13XGt7BU2RGQodtfrbGMkFz5mV1kkbp4L5Wf5ct8Iyahkh5lU8q/
hEO4rhrzipPPvbJd6B0sPi6LpkuzXIbABlc2qYSe8eaX80luWNOhFYes6ULV
b3fa8PDDtiSCE0Si29FrFg9wu18oIv7s2zhjQlU2eMULRQ1Rz5HzMeFckU4s
ZFzLEcYnVY2cmtPLFSBIhx4c9i2zzPeCo1WFTCTsm2SNMpZMNaRcr66Xe4RE
KazXXzjMoKIGQ/Ku5rNYXuy2SCwemwXSrNs7drz17RF02PRm6jBFwiko/sag
mLUmt1D1Z0XK8j41pIB3U0ohmLuEyzTJGvL766jrS26VTVGoSQpF/fGu0GMH
wv2Dril/eEWm39VzDyzAD9MDHatp2eiA0bjBGInKraQU+D1Yf5qxAAm6Ioej
OkNtCHMFRfp4odo9OuXTYoDf/Dy+iMJBbarF4xDTYjgBcOTcwnTtdMSCPkt3
EjTJLaRtVvLp8Cj61t1r0neYBA538iLG2fYSiGPu7+3EGjQzYJf/QcMBI/4S
pGV2wizw1kcPxugHpZGRejF+osaZmlDtFB8wrJwyEpxbjVK9HsWTJnkR5H5Q
evzsCOxKxcxALzubvA4n6VOE1tkQDiPp2jpsaKn0xBfKX9McGMMWqcrVjOgs
yZ9gwtY2RNIdmq4JpQmGFj+tO38x4HnmGKQusTKLOCmDW7KxbJTCGOFC89ku
lVGXT5xdX7isL//ScuIGNrxRE0u8gN1/6drvkPmbPKbO8vDRCsg9rYOebY20
2l0u+91SkuIX+Ti3MjmbK4RajIgGiT+Id6CkUm3OtbtsB+4OEK+hVaviptRj
KDvo3yZ82K0wwyUFvJeLZ2qjEvNQHbLWnrxf0Xj/Oqhi0axhOYWQqOHjGU93
GkwCxjC1v9IauO8jmwU7JbkZqZ4c3HGoABy44y7I6ExKY2D+0xHRKybhKAEU
PEtuewbErs9Prm3cAPnPLc6iJgikkv7iMt0l1tq9FGC4EzOLyZb+QttO3yRg
eVn0pS0AXzXJlYGtbw2ZGoN6cQSI4DTi8hkQf5RdJhtNOZ0FCB1glyf5SU34
/O5cdHPORtlu/BxTUqTMkS+OEoOxHfkeBGYkX6co/9feWDKlduRblKtLb98S
ToHS/zRNMSbjo19pT+7pNWS00jP+yEsM7TxZDhdTLUS0jDMlhlOaVEeZf3sA
tQwMBcGU5c2a3DQjaJxY8ydCx32Mb2IMvx3+pwLPJLoXjeGx/wrQKdvrAvjo
NsM40nIMhdmhO0Ipj7cfpJ+PS/s03oek5nLwTvYvmxMzkbkGILxjAZoTSYXu
Ce2deHqik/96b9PlVSAVeW9BuCgwXIWo999OMCbp4C8yi+6e9qzDXXcq3ESg
l9rhN5LafPMqGIWjmEJ+5fEcNx0+MNxqb4gYIfp55Q53PJsFsmEfIzNYFvj3
Opzmten4z24XDProkPZw0HexGG5teiJTPhm4kbcl8tRMo35R8R0hCIRd0BLK
E/NrFsWdPqADN+9o38xaaahinMGbMIcnhCwcvMLLCw8yW5fj1QNNEihTe6g1
5rSMy5dYXiCuCfnl7rwlviEQHEdGWBxdSCa0zmQIEKHZ+aNtzz5NddjAE/3B
ZjdibWO5QSh3I8d9M9i40EZ4PZFWSp8nw17lpmZCTt/hZMP5eBV2ANEafrZo
0Lx9zya04Ul/4yclRicEOJ20xtBKoD7Y9b+ZSsjlL8YAWUq5MYZo+BraLnhy
tiMZvmEmgKyww422Cbs6m3eNpiAY7y1SvOajldJc5pdwLNIg60xXn1fjpnq7
BS3YnjJCcrGHDj/L/K6YVkpG9WrvpyaF7A1ABwcURlIwk5ejRtTzx6XYV0Sy
lYPGd5AZafPI5ownk10rlQbKawXUOE528lJTl8zm12OTjzVrjf1uyzT/R3KB
PJ3akjOErch0tXxl5T9e3tQNQwJwYUDtTfRAdyepyAldw9O5sTdd5brlwsnH
VubD28ZNiMyIGGNOg96FYRqy20ATNa7jazv8Wx8ewKC3kxhKglLs5Atjx//B
lK+Y4Y36ViH4SWUfUxakgftI6j2PHMcQTqW0EGyeIoz5+aeL4ZcxoEK1Hm18
9dSgzmcs01DppMnVD7eHeBavnryy2NTPG9XvfMSQ7H2lcukbndG5sOdQlqBL
8VcXepuowTU1c27bCbRcTApZf+fmAEWQ3RcZGKZ1rJ0p1mP+yhx2Ulvbp/b9
zNftppDHdbGxINpSSZtbAeuGD/a86/3ojZIspjQytzkmLEF8ER+AEY7j57LX
vjVIPQkAzAaz4mbkOdaKJLpNzXovz0M8ILGx+F50nxZ8NyZHF7r+7LnaTWsM
k8HSN6c/0z0sdCgKNE07GD/bOAgfStaPTxvORs1esst8kdBCpvHlPLm4xuWT
8FPjCKtlgtDzqwtSl37r++OscIpKqEawe8q6YHUGmuUThVEqU0ExgyPmYsbV
1i8o+eO6mbvHjyib2sHO3H8gTYT/SU4KM20i4uJZ9r84sovvjQ4Ds8lfORyy
UvG1InrgO58BpGjRQlfVvBKMfPyHm2yEjJ1xHPDkNqKSxd7W/mryr7t6QIzL
yXd7dO6adwiqtgxWdI7kDUaVeRRVpYyUFWfYerOI2Bopr9F6FYkdewmsaPIW
Am76mVSJ1FovFoCq6OcfHk/D3p65KDTWzSIa8C1x2YVN9dx1uvAByZv1eC0E
b5cvri6vtPeY54xyWD8QbkLKR91ACJRWr1+X+GkHosIDyyf6W9s8q4ww95nf
Fv/UbXPU9LKDWtNhDxL7wG0wPiGSUyPhZ4+iPHEOxHyMw+RBwN8feCjCClQx
xM88yOfT4YD2xi0vypNnGMY0MaSHZ8kqA07ymC+3ULdC/qbbODVtJwW7NDN3
wWPL+F0VkbALBmQqAslykhDt07vW5f6OYM6fYyCiW2Lpct3hcinT9757M9rv
dkKcVdyMpOM27WPz60p50Dtj5FnjVMIssn7taLNSm3bvCudp2Q9oROUeQ+Uz
Lct28l9oWV0bVhmMIlt1EYMcJRpYgfoc+iv9vHcyyMadWKjBTjokHGP155Df
2XIbtyEoZyqwrvthM8Yoto7LTBJhmr6AJ8PljXB6FzdEjALnkmPd4QDuvdSo
Z7tr09cuAgpC8ZeWC9LmNy3KpN04WWzEgMpPmFuwH3nHR3Ex7xUF/+BB2xup
XYRjTOWAI+62JIK0cTnub3cnM1CfdaLGaq+NwGmA3Ssu0U5aIsQEwGGDTG/q
UK2yHXmEKQgw4zvGxeKxVkRh/p3bGa5Vh1JssiC31m5A47/DtXGiK+bSEkSj
mCAvYMIFFeaCqOyejkZ0v/O8Hvp5euIz2H/Vv/uKvCHaGf5DB7O/aeoWSGgb
B8q+4vaZRSgXXkaUlZsBQYmlorzxRBpNYDQNloTEmzWNd4cqoShlmgh64idF
OfaMTFE14Hb9DhKM+w3+ih0j2aaz6fT4QsIANTOyOWHv91jtFckcx1uSt0GE
GU49lqRYYcMwZEB+eHs9hstGiG0Yzy++Sr6B5yFO8Cv9ziQZ5ruTiRYd1yEl
9zyrAjQQBP3Ob5Klf+cFnHvtG9NJ4thBXhSHyDm389v/+cJ6IkQBRNg08zW2
HAZqOkEcTymnEkO/eXIngK4OXjqYFB0qhQHx4jQsOFeDiZJm+NPZzghQI82g
cVOcF1guT/CKUFSoYQYR9GtFPb959kXokkZC0BnOZ7SYgT7R4XOjoQeYqfbA
Dhs+Urgr3uF4GJEKwXpL+jlaxlzHzyWdi0lehGKzNEd+OyM8FKjQkJVAndG4
MfmdZCHV8z8w25KSOgbSJ76MOaTS951hOPfSd9/ZlkWCurHqYYUs3faqAp3l
25/nucDAr/J9/JcTTgxsQfTS8yyX8SjSWtL3lxf7Ln7sCvbWBDs0OPlyssmE
EyK4U/S0kaHWYzqlwLcNCb8s0Oyr72AKhe5zbLY0YZRKHj8D+NL33D8j+xnZ
kh2FIGaSi26vvHs0V6oZXPgPAiHuAsL7HdUBlqtqApVuOz92YhqjJBB8DjT8
v29T/f+33ACXYpK+wxPtMIRiiq5n93k2IOGzcdzSeo/JL59Wm7lsM9zjRy7a
MgUbm5lp1bxMdJk2TeRcGivwlM1mHYfFzDSu3k8D/qazI4E8SHdmy0im+qyR
lAmS4w1F2MOx7pzmaSdRuV9eBsGh+dGPBJQATeGGlvmpgA0/fRO+it/Q2h9+
yiGdeboFeNc0c1h+FaF8ykZ1T9tqvheyLaCwQH3L3/My9vNAjvvspvcZwOvF
T6LgSfn8oJhwt01x8xYN+NHYqW542X76OOagGTpP+vgV0J2cTaf0fcHO2BfP
xSCZi/Kq8c+Py4eEpiVtCaw3pAmhhfzJ2cSR1zdOSJGbIueKjzAshcfiQqZE
c+PTizfYLMSp9MD6w5orvRzaKwTo42wvYeGvSR4U33b+r1e9OKNzPkuHo8zx
WyXiP3ErxEJQSUD5MIFM1jtZBF40sc4Llf27Pn0o6+MWrTRPQ6KHAushm7Ap
DUw4jMaVP6agrA8ygZUEh0KtMOGNfpCnZpYCGIBanDg2NQkFWoJp2a5P8DQ4
XiiV3ZmbYZ0RoNVq5Rsx8DWW9k3vYI71jhXBoZH53OcfNY2RHWAC/7PO4Wkp
xkJlez4P6w2JEHV31JK0jL6/Ldl0KXTD/qIFT3iLXPPFis4Lr+HrnSSOojcm
3k4tashmEnIIhbHTIJ054OzW7PAaJu+vdbPaT9HZteRp99nz2l8EYSq6ct3T
SU5U+HxumE3yqlTrnUhHcufs+ikizoMyNaBOcZlBsXnA8uH5Uha/bb56s514
XSkfSty+F8ZUiJydeacTc8WdhOQlbhPu0BVHa3ZhiH/+8rhImlZpgMG81YBO
6n9IWMC62nKO7YorLspB2F5paXMWX7RAxtUm5JY57Cth40GoDmWSNy8gXTD2
vHk328LEMnsOxGppA6IGb97gCskBLRas4BUd+Y5H0HAPFVsMrHvLJ+4UqkuT
BeNLsU34YVyr4Y88T9z9V++u959c7HA8Cqt6WQCDABlXBbBX4wbdh4gj1dPu
ZlBLe8p1ObMAkvsjAoOzvulVlQdGyOz0IbNkpdRCAY5yjPLjWp5hnfDjsWWB
II/JhOJ0pixlHwUdI4Bwvhj3BqHcXIpPPs45tY3AlXRf8EixrR+ExPQa+ash
/fP+6N8zxW+mPz3ZnX+fxIsw0A6iNkSbxXy2M4LdnesUx490JF77CzTER0o7
uNHaYxKM/7RCUmnnU/CFr0O4+O6I74T/iqsSG5RDZGdXb61YOvSLkXPK3pxP
/uLD8TUzI4V3ZZOo/Z9lK/xrqCgVNCiO1KYFh1FYsl9FVIyZm8Xnx1JpvrRa
NiK/4shSUh8tajRr/LN7p4VvwEaVw0k7MKSyKYfor6EuJDqfIBjgKM6HKaJp
W1OGSzGh4Zl/1e35CfX6vDlZC/lRTGEoR3wLs40u0uMui59oyv6ActKeB9zR
vuOop+1AWptM81nhrys6IcSxxQVMdX38FqftcIpZ16Jit2AJEBYtZbiMTC3h
xFXY58kPLAMVvIqBQ8zHNHbbBJh87iAkMnjh7BH/3pJ8jiMG+Sf8jZmasS8q
F8omE0aqw8Z1P+7G6o7+CTHcQe5wlocEr84K5JI2Ww/Whuf+2zAG11G2aZtS
1ig+w2GBYQk6KNfBsJMQKOURQR7v8eMtOUOO2Pi7nTyX8x1edovl5MF+cOo+
/ihbgn7L39RojII094ISsgGEW9t6+ZGk/YmpgK/jYam0O0dAYb3LsyxNW9eh
Y0H/+QFKRIkAwTdqmbzzMgJ+F187GPlhZzsQXdX3Ga9AMThdXauVHXq5BCmX
o+/Y3fdai0B5G47SISswDvjpFu1+wGktkvslmJxbg8fR5Q8JWbFrU4qOQDow
ymF2zsG0mavPDKkID4SjSqcfd04DvJRqCVp2U4HG9h2ip3JiJ1SDK0UKM3UP
3F5az1IUKPkvih5BcSyX7O4DjgVRhEVFH7CpZWdpauAJRlykAZ7cEJyhRP7x
Ier8Hw+VLD5x/dLMCf7wZ4wQ5nEG3bBQvXh40TnFJ4Hfe3ABrXqlSbsQ8zTj
238ufqkezAhYz0I62fl2GIBjtELsnLUNtQOicA36oT7hZpZbxLN7F1C5jQAZ
g9fQLCLrlwm337L8MXEzJIPvAAolgSfW96bZuz9jZWwms7/HBPBJ1nX3y2iw
d7zssIRnAwQ481mKkzVla3FEvX22sM4CqY2RdKuEjlSEMmR+ZIdt7DWd31me
7GPUP5fjjHvrQp1i3+ar1Aic7WClmvIIUjJ/yniMDRWQrTPu4z/rzorB/3C9
0Vh7cX040emc2l4EyNULpQD/JHtyeBcbOo4fSkb/8mMquBS8eeHSBFj1J1kv
b4D++vqpN8V+YL60iPGyZ6t2GRJt4nwUbt73sas6LpU+huuQS6WjmIbOwSQW
eGfoSIUA1aMtldqSKOTxDCbzRVt5WZnVEGoxHWUr4eYVSS7GlafhxNZDEmV+
UXZnJkdj2moMCDb/lEQEkYVIZk/YKYYZpFhui59TQoEu7HS5s2kXCipToIO5
efRZDZ6VqS6ETgfFcEQX2dL/OU7G24oZEdMzjEGl454PkfuVvIpNdZ9H6a5A
R6PQgFrwGoKPE4ul8OempLlXAlr1SgoNr1ZAxqlcGDaCkIamMKjJOVKt89NU
/3DxTYd/KrQWyhJN2JPF9e876wGicir3ebRvz5oHrskBn/CJObbXgCS8gNMT
776HyvyNXIoIco5MX45tznsi5AV7r+DJ0Ov70YIcXQ4EB8hOtD5+mVCz6Oyy
uR0QL8TeYoZ6QkAIuyr6QIYGy6CnGr+vdHM0betfim32mKt440uJ826U+1IQ
o1y+M4rvTclj5d9OjUE/43OFQuUs+g/efmPNKXhkRKz21s1OzTAJjq8ITTxW
8pbLZEsRZWCNvQ++KShYewqktrKnM4LVM0MFYR+Trp/stzQ8BjHYtEndlfZi
F/YtuPu8VF/EaFmoS/4/pOViUC7cvLa+kkPIh1TcZDdmWUXGP8PETEAkilUG
kYUvTGoy5fUuL8O0EENyiAKZOGLJVK/BMd+pGPWFbpFjTYjH59wr3abLPNW4
XuLrhAvDYJjyFAI6uyQzAYgzC/ShSUxHAfciw7MuOCB/nIJ/CgZtrv0HAP0m
MTmmLBjmEd9L+rUr9aIojd02vvFL5yWq7dhOor9xhKMAPy7LntCUR1oe/dAt
Cul/O89owBmcogb4fZngEKkj0TX3yUmOd11SQ0RZC3WMZ+its5id8oJFuIdv
1y8WdDLGs30zqiSo8E7ZU4l243hKkTpduJeFp9DtOUDJwBvxU8PXwwZENOuQ
Ja+lcTUrXibD0vtiv+JTkJkEskvCgeNno8fB25cLMpGTY/iAh4yApl2WdNTE
dAW8c8PM5wLGr2RERMm14PeXVhCKuw7vDydMSFUdm1Y5CkdQINNjNo8b9rmt
Lh5SFpAtRCDS9RPKB9mhZeE8okKZE4cUu/Qq73Mw5hRXabZnn3FKJFw3eZJq
YyKH9Shxx9levtB3BW8pgVbGI8bEIE4Xf/4IQzbSgV8Cau5ZuMEGYWLXQKK3
a+WCWxNaPYo/JtAXAwDcrJcm0o9CQC/lofpJJeWanzsUTQm6C+zJ8wm5OBqK
o8wg6rMUfMeizMWxN6kITSJzdlNRaIJh1aboUVJbLCm87Gh6SpP/bZ5MzP3e
cym9/EpgqZfbyMa0VgU4uKDOz1UWDUmJJ9RxEJoPNwny8nmyk1KJqdnOeDdd
RKYcKTwcoui4/nmWH9h9X1JrPgsFUFTAum0gn++pnaFb7/Y79QJdXv7Q2TFB
huegslEIxoIzKVyODkvG6bh9+XVXJn8BRz0q7/fv3tsa6NBqr3ZgD6R9bOrC
Xcj0ispCMh7VFwqVzi2Bv4AgyTVmGC73xDYw6R9D/dMU5aWdyltG2sIbPYIW
MIh8oJ73rqFWcaPiXbZCfZ+2CnJNG409vQlSbpBRmkgyAG7SFV12x/7gRi77
hBOkWTbVlc92qBP1S417pZuhmO5EZBwfJAJaSKfl/uTUXbcYluQbd064+0mh
RVynL+OGkahMVofrwPyqH/4JBgEgTJsoFgB79yifjmi+gInriYDeAT+d7DEg
WnPGa/Q72UphqjERPGXm6OkN4F7X1bRWFRpAnJkflun+BsbJ0VsjuJ8kQcWl
ziGVPB9hzMW6I1v15IuVPR01BZjIe8GaS2++eb8jVV0HPDHb224S7UiXCd/T
ca2iyuF6Q2zBrXWBRUwyep/JyrT9HByR+wZ/LU7u9l8FDZp1GK8tZl3BBaUV
2/5LqVbM3nnC0r1vb6c6JjFWKBOcMROqoK7dsE8asu/Y4u6ezytS4awJDkKL
Vb+/SxILPIrx1IY9Emdzg6bhtWQjWENSuJSnZXzXqGym+hFgUVJmeWqcGUOM
DCubf7U+OtsP5SVVsuEzeJh5Jqlq7Lrd584+r4dQAHlVSLOTOYfCQ3eje0bj
CO8QomqctnfD09NFdHj+zrFZZjhDV5sL7SHg8PpO7G/sOzohXuyx48Tqj1do
Nva6QfUsWsMZBb25fDgQn1vCYM4VHV9shx4KY7EFWS4BTAsrIUBxm3GOgxHP
lOhZXawd65uNR9heOJgmVzwRlwC++L/KcQwzh2YIXaWX+HHp1IvkH4oFCKLR
u50W3HVJrpr3CUVhIZwmjh5YVqslK3Qbzh48wTKobB9r0Clpmzfx4YR++HKL
rSenG62hRneFTK9ZA4SiBE3iJCUEWkrHQJBFxvJjOlibULVYUICx8lKuvF32
xAcsiOAMPWtGi18TZDU1YCez3nkqdfXFPGTFuF/LiZR59efyLMeGkTbOy/Z6
8fuoIMF7FQ8fsUjmYuD5YW6u+nEfyq+maqzPcJy6+LagLYl508CszNteVcnS
qPQz39LeGa+ijDRSM8Ve0NxnHThKR+WsogLscrxpgtq3tob/EvA0VKf+3zCc
qyjnwa9zWM5kod+tWsuwQnL9GNZ2i4oX4f/kW3oil5cuM8/8EI7HnOIeZJ72
/UDD/QV0n6S/vPCw6qTmhc7xzDS0AJYB/NJe543tsIuOpCfUW9NQEibfx3Ke
F0DdylggDsaFBgyg8z6pTwXcsraRse2kiQ2DxDcy6B2KXkkaT0yiIzVGzTBi
aVbD0j8ws1DtTkwjdVxKJxYgvh4wwRbVEMMk53QtHj8HJb86JWGAiw1vt9Zq
v0/gH4Ki3/ZKKOnOAX4xeAxvIFtIDvdFU27ptHAN0o+OBEsJrT1QZZ9SSwPQ
4cbT0NVnBEoxet24tXX2x0aJSZxW7LALl2LpczD29Y3GlPnvIHmplSz1cgKz
mRH5jLK+tRfolpWCKLklHiiEk95q3h3yVhDLKoH+1EmGdEc/2KyF5PmInUjT
z+Ra/pUnYPJa5N4PPVqIPVPVzzzuR6yF0L9tdbCC9ETGu98p8KYpEAPmejNL
dpgo/BnKzmXEGG0NQ4fyU2NkOM/M2iq8PQtzYmbacUAiR0N8HEfiAztGCU9a
B/f0MMl6Uo3s530ILJA3X4IuDgqwSHw83HwkruiA7iVBrjRbzNsDHPL+6+aB
m/bQbt28Y0YThQcZX3h1CED9iaDDfsbE7qeSnJ38YNQFg0K7FnajwUOBK6YC
Me1dAgKn+cBwXZYvzAN5uMlwDfODrk5BlEK1Kb5/9FR4ROkXe4warRVkpHUI
emNs44teNGdq4NSlj/ssqbmtNU3vSpppYXCZN0ZPYn9cVBPsIqvDqdkMeJb7
s01LT1CYx7Ju7pKcBB/AL03td2USU0bA6zUWXQJZ0IWp+hea6ApxG2NN77sX
n9iC4euIawmidSdnfOlNI73LllDW2f9kaunx3JWrcb35yCNwnG0L5lR3eKz8
5FN4yATbGkvcYI7fcNGUVdgKhl1aqJ6TMGyP1ZHt8SbiO+gqEfPE2+zoUIK3
pfJOAbkaQ95RBus0MYg/pDpEuqBVrQ0ILLH8Iy/2b52liLlpsMEGBKH9PR18
UoHmd1wvvdlLFhijh9D5UwYIoODWlI5XDTxCwHgm3t0fC/osaDNYClXRbK2d
RD0c4h+MKqtfHe8XqM0jRSq0IAHoAyRDHMmLSvdNc2rRw04jwJqp8Njya5g/
+eXd9akIfBc3eXViFo7AWnVFeoFLq4SGYLaU00MvKDLx8Ezpdkq1WBCTJRTU
lkvXUVHEwttMaovjze4aAY4vrYYtpmtx/a6d/lqbLqbRknPTbQOuBwZ2BbrM
Oyz3c1AHZ3Bqo9y3lQaDmeFJq2vIbaNacL3DuPJtSNSInJuyrP25y0Ee3ZZU
/PCGME/dvqyLUTOcflhTNKmCYga0cuWDQcFYkd1+5Gpe6R6+rDeSzTFEIzp5
1EiCdbn9jji68OUphoqtwZHbgLQylZtyHr+aeEOCMv4jl2QBsj73w1Rlt1N3
s7l3RCg0aQRrBiRVoJYNxxerFUInWCVhhJl10dN6uLFD4cE0vdMuwOOeu6Mm
R/DXfRqtfn5ZeDwzlUqEPdKSc5cGxz/mhlS+7fTeLXnw02xkVZD0i5QeM1fC
CKzbu42ndu9pkBJSupTf5u5AOuFjvpsShBJNL9MLS9ihfDHTPMOJBwwuAdFB
yxYVqtsAJFO7oNTaUwAG4EUw1IR8D6NgQ5bt/vBMwFP/Cg+1ZSpkm/dwQ6q8
nH2f1ovkUFxMQK6VdkodzsG1eiMkhaK5igi7EUdC0s1BV4LoupXvbLwEKyBt
oMTWZBnUEVu7AXhQZbGVsdrxyokBwEIHgZGofx60t8fSQM5veSFjFppIn6Qv
qyui7IP9KWSFl//k4cXAXRtP07+k4w8ch1bmX31ISgNzh8kU4ZvtaDEaLlK3
AQU4o1nB8g6ijoYStcClPy8GaGJzLO7Me5qWSXpZbPNOE2fUUWijIgCXYIsI
D3v0eR5/yGrcvaSiv+YWV3YmjY85GzZ/luS9JybcTgZRyg264RgxEmr5Nv7T
pasy6okBB2n/SV7DfSUzP94KRCtT/ugQMhbvfnXNoJw+BYjZ5sNhJX8YelMv
NGAuxAIbfrDcM807EDfyzckGmwTdfwzLH0oTGVY+kYCjtoqINinaIDIwfvtO
no4Wo1/GcCGSLtZ4/2LetclAf7HrCTYtnnHKR6uFMeG65orHc/O8iiWtI/dh
iw4PvdotCxn+i/giby5W5GVVewm+5vESg2wwKO5HtSyi1Yym3RaMHbYQjp7o
B36u+PJ3LAg9YYUBeeW0XVv76WvVTHwXbYABDhi0fnOPBAh3+EzSDOyBsxnq
Ew8lL0Pd3indk0l1UxTH67bnGCFiJQ8Uwsqw14vITb5acbJa8KjU+eWtBOOm
HnihFLNFMHzrAjv8B3Sgrsuie5ehXUcSkdjZj0yVTfSgfuCa7cTpNMyWY8iN
2VVFNvVDJCxO2NwnDQrM7lpngAjJxbXdVYoHNIAtQeNvYcAqQdS+mpCkQ2GW
5avZ80o8oIExD8eX11QvsVdG4LngAH3XwLg938mRTB2t+GrlO0seoQYRCA2Q
/i+opDleQBSl43sNjMqkl7rNCAGW/1oyd3x3d2eLI4UQ4y+SWOoPmR5nJI0F
KjnhGYedjsKwGQM98RJ+2qELSIIs6h/EKlnTZXo5HEiRx5/lHrL3HwcKAkQZ
oXA5aZua0G4QLGks4tvx5dEZgeMwMFBOZnbutknVvVx1HCmItZ7iAN9fhuSS
bUE+sLnktgZU509QfSWmqt1t6YsKaZeKmqnDpvwpZQ16VtmxQW+x+ueSYhSB
rZi4F5kuCs6VksYGITWY/Jn1U8CHn4dpcwPn/+9Wu7YFeW/R9K9atLdMvFWd
oAmIcqwPHj+h7yBMM/bW2gzsL+t/B7gGi+XHMyUjF5NOVNdzuX1lk2cUtxq0
p3jULT+NoYvtcfkVNC01US97LBEw8bfR8QbJxtgJdgS/BqXSOA+24XcgzUGM
sF2CQT+UHg61XyA6BUSJp7M/qC2xlqCWiWwXf5fTSc9ODfw7NrXpA5mygWFB
FDLsF0gXQzxQf6RG5ZjlKU/WgOUSH8Y+hvfZEdh0Oi93L4ZNxWaMh6Y/bBQF
mxmvNaFJ7clX4lL+IXlYstq7suKFCwO/KqzTXBZDyP9vEM88VEvuYsrvX64+
Kj1BV3sgCluuK/fMv9QyxE6kxkhd0vJ1QjCW2CEWeHI7+pedDyEHz4sjmm/s
+6yXFm2jyd5XsV+bE/1qTAt221GU38uNHGdxiNQBUM5TxS86P+dH8wwfxvcX
MQn1IwKLsJZUcn3lmGk4+uH+Z0bCPIo0jJ/DtzgGxTBVSGv8aj4YDiZ+HyCq
wOXJIY5vSUwx5tPFzvJG2yivEq7TwqUlwxxlRVg0aQdOgwVlRAFY21jgDaFc
r7NOQPbzCMJs0Gg5BP052aBmN5XKWYnER5hMR3XO2cYDXvzP6jp41ZLULzMC
d3mxs1x5ztsqLAViLdSLwcYZb3jqL34ps0zZI1W8p0De4PfPkaX8OwKB4yss
TjIShOkJX0RwnNG2bKE8fIERGnyR0+/aW36bqEjQhpNcjaFNc5jGhPnagm3P
cuOKK5ISHvEnkaM8Bfm7zecAQdN4/eHRedGGBVc/z3BE5Kx/F6Lch1NORP+V
9upGV4pqaCF89WJCcj7PdIl2Vax92EF44s17unv4WkIimz0JdKNkend46JY1
fjzwMl+Ya59yWSAyfrlu8de8f1V9qUW/zlC/8lH3aEORaldMtsEp09O7IcPd
Ft+j6wXZFjBoCCyVxG0aQhH9986djLGUuJg0cBm8yomPROE/BIG2hFnMOjXy
A5dN8dsepzHzHrJLBakv+TH0zefeDn57pbAmjCyxsHBTegibqhdxiiJs79Dq
QL2uESiTUebw30NrQ3cC1gryM5gdPLwuNq+xfuZ7zohlsSrUApnnDzjF30Rq
jPiecHjuYqcoFnMid7XZl3p7C57PFauedm0e5HvhAXRpYDeBBD65EFHZV6kl
YceWKV94amymc4gzABI11uf51AUAg/tKcjHLza3Mq/qm15EJNLngfiBYpuDr
jyHE/IpEEi0/5SyMQZQL/P1Z5ELB7vBnRp+ZHUklxWZCkpeSKqAR7u7qIpoX
6miAvrEdn9X3y5X2cNMeWnVU+dy9N+4Q0Oqif7QRvPHV7lXGWJfiIuOrQiHK
4UGZebt+ENdmruJ8OWEPnv5LEGPgvZjPTzsQHqiadLKFAawY84PGDkLxey38
F4WOSDbrxMUhnq7dQQzM+0+kuSPXZuDPVmODYIAXENdB9i/zFOhQYXm4F1t4
py9Cgk9iuwCukj9UM+RdK87BIJsPqU0OJWFpLVmkvpN/6M8kaHj4h8c/rbAf
QKlbsOga6M7UkG8CvGQKBs2rmCZeKV2Cj/0T9Sm8PV5ZmkUBk519DjINXvB5
TPcQSxK/ou5FyukceijrAAzkcv9xK1EkNZ6F/K1F3J/jgi/uMsPf9ac9G5Ev
2C7uM2zvLDn3NHLa+DdHep/9I8wn/AiLqhVQFi6AsPhaeUv5VmqviCMphLlP
MHYTgQ8DxlDtIOn1kdG0COUbevw138GrKYZTSRrrVsgvwNVKLJMgdWTAwfhH
HfJy2/PWL9qErVM+AX0QbuXv6Mc5PCamH46I3ku2AIuYRmlf/KzF8j5tyI5T
zG8uSTVz6PyeXTyMk0u65IpkX6rDzmwiQXBkIDu/0qOaN/3FqUOcTUBffUtR
hWTT9SeX+b/R3SW78H71AvQrPaiP+Ejk4rR7iaXfP3yG44wnYwmqF5lgVup3
YHv0yD0FHBR+96kHJyXU0dr/2qr5ZcjjZnzxS3g2FF7RRofg7pAKf/iKW+HB
lYn07HsA1Cz/ThoEXKLuyd0olmJyjuNPcBiS3FRCrhmOyoEqEfWh2R2Ykv74
xRXGJVR5uuLfD6Ohz4oqvGx7hRc7VyI8NPPjCnclitGsK2lMaJ4ZK/bKMkRt
NjArBrwkFU2ZF9GL6V0V+NYmsCSk6rK7dCVS7wGiGit9R/d/xVE+GRWoVRjE
uOkdp0xoV0InpHbu4OxCwSdZ5XarnIx7F5DDNIksYF6peDpe4kc2+EVzPExs
aTPPqGxdRiIncDjSVCE4BCvZe8hs/VPAGJExX3T2Pq2AutJoczNgKCvjzEpL
XiKnHPpqlXdweIJ47t6gVdWmflimpHc2lhwyzPTyWCnKHmnTyHHKnmLf+kBx
a555npnPHpZOo7w0+oJ/h05BojzyTxSqcVggSkFgAqv7l/es6hXTeTt1veWY
fJ7ggBWfWqmP22h61WjHzzASY5TFowjjCNS590EdPzLyzB/20DKdW+D7br/l
xrtZXt1uo33Q71H4v3zzLPYJSZ3EyeMBKfD5EU7I+VeyBHrPwz9yjmgCNvCJ
+A6VUe/qOEV3cdzOhSXaFq0GOqp4pGTDSvDHGtW/KXS5Q/BvBol/urXiZbHz
yRL2424kd6JhGDZAL0LMWxShEpqtfif/qtDaqj6X0XkYocz7u1g+cNi3MKDc
df/T3555A+oRHBkDf9IMLjxAvlX3KDQtoDPtEPuxmHejj3ZR1Q4ih87m8wYe
m9RHIfMl3DHql1vMRNoQzt8ZrPsK8cKg+/oD6SvecHd6ctjjFaZ8JXezo2BR
C3oLSUDrDGcH1faazi/1a4ajebQReOAAZBsaMUZRask6tPfp+thHUERBdifZ
vPuumeKxR5mpnSGgAaBYdB0/SlhONFE87UTmw7R+UWGBStJCT/IIGoWdlKsj
iHpl2CSFPsUhoTjiwBl3nlurAuOXxYm+cDitbf3QBfH6cyxqSHgYosQgv8/s
zLATy7HCMPWvCSZk/gFH4PGrLPCJefjXqeMECxkD56yO6toTpHyBtgFnbXnA
MctxkaNyxlek4+57V+X459pdLnQha2T0o6y+4sflbY4xy4pGWom3clUwxs53
gLmMmvgP208U+Z5s1xcLinSLNEhpFNX+D3Fe/imVntI+GCRJacapIYajd8hQ
p6W5R61uHMca17oyryvIucFmTuak7rsenmVE30//uOLzPLLEaNEuJvfX2m7+
u43HuScMHTz/E0sqB0d2vIkBBhREYMeJwIkDhMJrRx4g8h0OnQNMpYRb2/Pz
x9AedfTjOa/mEqMWpJOoLsGYMAtgPiDKymWQLEY4NMiPRquA5LctQnge8NLV
GWomnGw1FFJseFIwL5EV6Se01wg2Db8HqK9F/UgAor/dyNKc4Ij1BZJ1Ua4d
15ZhYh9LvFnNNpFkSC1RBTsSiQMeC/+yaem1U443bewPr2vD8sB/nEAvegB5
nCuAzwJEINDkxa8Ne2VB1Lnldx/0vSnK/8GV/fGnCIkUAhlRGYMeTi9DYwOk
O/zL1UiWxg9foLfzQIX6HGGee6N+N0rOUedqMjjS3AeTjdq91yyj6JNTOMmc
GapEnks6FB237SULjd0Fd8GhK4w1BmKsTfTd3XigwG+xJws9liLHeiBXskuo
PK2mAhK1YejOB4SRX8EpR5iimF9IljNiuPgRdkuJl+C/9liSFYK4vnn77dHR
qgSRD4EisGhwSI92LmpUGEXRpWVIsucNBziM1om+BlqNdAQ68Y8BUcFMm3Xh
gjuZWTxoU6aX6KwoPpSPCXESdJEKsTasvD8ZcrdwQyKSXHcfOd8L2B6GrElQ
FttitgKsdCnLNB/5CLl7jj9jyfbS0Z6sReiisgYyxTSDqTNK3n6V6u5QrBYM
G0nuYVQwoVKkJUBx6uyo4QpKUEh/YqECkkOKXRezwFea5RZ6VyHZj89WrNbI
/EkPTKN/xUGZbDUjhjOqIx6QHr8bxFw6mZtEYy96K7sHgB1G4HNy1SGdY0iC
SFFa0PW9zQdtB4WdSa8JPJpi3w0NYsdLp6Hcf0G7bC/Fl2tkH9zXlJkNVa5h
mboDmhZywUkLSN/EcXA+WtvFlKlEKOxX8saH322ehdbeFNf6XLlVp4dhhV8R
Tm62eDYraPsT0+R8Fi7iM8CcLkSYX+OddUBshkWGFFsZf90FMxRhzAoVGPJ6
xrRM0MpVEYxSu4aCQAh5eZBNu0rZ9gT6GjedGR7ZDMtEigDonZ5Vip0qj5DS
d8iWO4X8mua9IotFtTLgTWTThR/GBwHdrf2xMA2eilZe1sKhMz9SofTUS0LV
HLKUui0oFFK9nZZcLJNMd1TPhJFPyFLYK2K1gHQxID2VSKS7iaSMMu6wqvtq
PKev08pxQ5LYNWLVgeqUPnUoXIP4JaPMVwp+ulPabMhQqn4L3mVv5CUMW3U3
4xWA/C9VqxEmdDxKdWDC7yPS0J7cJo7KAeTC8N8CMK48mBDRWqti9xxwg+ap
Jh/hP64y/BoJ2hczld3FXSJbbNG9D/2seXdoNO1GzTTPBk96dhbbjwDe7cSb
XGWLTaZfgaDtv96M/sWdUmQaVgBnC32VIWC9FANSRPTO2dvFGvcTtIDLJDma
kMkn94xD14Z4DkLkDYJgH0O9S98D45KsK/UPULhmzko8aZZf9uecU2YqMwVk
fxCXo0MRVkFSOaCHbYrlcM36s/oApZJrZgMK5XU0BaEGAr1nVrAn97F3HC9m
ywsoq0jgx2bbKeq2ePH/9M140PbisxOiNQ0aepKZT1x76V8NHByY0lMrOQXh
T8ECauentUm9VyXJv3Bu3jtYVvNwFxjZABwR/sq3VgZm6QbxrG2XtQE+3YvV
OpeEmEcDTRYVPhXOowy53dIivB8Al2EZBr17gsL9wD9xMqP9GnH6jbjLppSB
55p/mD9QAk4U/CKV1DLW9STeWi20qIbCtbTMEy4sYOaD5zzKgJO5glKfQAD7
e01oj9U7OVcWYZGaEI37coTVeXesZIumB12X1TeUofh+XFzKh89KJBLHA6KP
1d4F3Xcc4DEyDmNMtsU4B0Trl7BcyMwpTeYp4is04ErzXbk7lRhFZy5LMa/a
XgLYVmcoDZzKcfjiz8ifdOJ24p2VjQL09Ba+mAk+i8hPJFipce4LtjDD7Rjd
V50DOCPiEiiABqllLRLbKUCoFaQM8O/RvVgJ5rRavm9aTaZWYTw3cYH4BVFX
pMbkq8AlOLWyvs0Ww5B29Ees7d4gPGDHG/Ytr0xBmmJDr/tlswCi2pdjFiSb
cczgeCxiBoV6F04JZ5abh6r3739VSX0yrjKgdq22FG1yQ6s1zQRixxXpcldu
wlqssXQ5V+d6if25vpsDcA+iH4GUSuMft0y/TLA8sz7zTPUfo3sfF3E8EKZn
c7Tatcfez6BnKYUhQbTAHW1IaWl5LoE8ZuwtXXfK8cFPAfJ8jyDnlnCGgqaW
QomE0nMxxihO/+dFE9akoCiSkXwE4gor9mqdlX1k8aPoQwAm20iPXu0kIWPN
qCz7Xhy1gjWhHkOJ/RSoMjR82pS0tUp3LU9P5xiPJHzttDsT5rHqpRd8H21y
LcNRGq6ZvSCRMPkizQaxdGBBnxPVHfcO2irrhKnesOAzTqvvZkGP0fjDBQxd
m5Q8dmhGFLOOZmEVLdJedw3kbjGxqiC9tHLnRmlPGZdQ208Kymmol6Mt+qos
DzZODEtjRvYEGv1fGA7oMVopRk8mqj8VuI/+CXvXL0RCqDd4aWGO60jvJ+DG
/i/v15zIUO6ApvE8FbVZPujSH0a28PeKRjMnHFoXQa+6I5iUHxGuNyhfzalO
HPcUh4Hvq9Ni6IJJReGkM1fzIfuzbfKaYcLj5W1wBJ/wwwf4mpGxf1n6EI4y
u67D5uUPJUup2oBsz24kDNMmsmvhZ/B7f1MZNsaTfwT+ZLn1ah5b+qLJ6X98
FbjL4XDs7l+REykpobY8Nf5yCAnmVkFSffltVmOliKOXTEvPsx9jLedzEZvG
k4jVoNfqDYcvd/bFXweNZOsE5WqODJNRK6tS7Z715KF2gvr2AF16E5IFBc+e
vYgf1kra62cde6OOZMWGQVkYE/0j7O668PAj8RVl8Q8ae3s3IwKuswfU0L3a
iSiL9ORINwWKqrnt8B5Bjsc5ES/pAdjPn+G299sag4ZRJWkV5jbvKxfNir6C
Tu5QVPxeDhKa0lZZUl98vu9As7ApER3nQm2STFBp3eRkg/mz86a+DoiXmSmD
639w10qZyetfrIERVekcT8PvFjvZbt5EcXee6ONeuujNj/LF4khcOgBkeZqf
8l6WrKALuf8kyJZGljbca/ion2MJYyif15xOXO0hq2IrnlkB70sJBdEl8AqR
JVedGy0/GvUI/EvsaJ10AiJ0Q7rae5K8fdjTfQ925ks8DNcqTXmtDWbpS2gn
EJFQg/vwJgUBx79IgMA6Xx3jLrp1qzpwy+mGiXtAGbplmIu3OwwDhyxfXatk
5Cb16FqhElATjvaEHgg1aNcDLBZwDgnyE0o+41XgadbuOjDDlCdsUoekzeRT
RA0z3x34CGhvbYTR5P3TCOQSZs3S+R5w/CFTQN5aSiqZnKw4IU7/32WJK1dq
rkSv5SmmQjhGtldAm0Ep4bOxIy4+4e9ZP4Tdvrjbpth6e2HwI+t9I/aVZHtF
FhvWqBZ5maSwxgJlMeIrbUYbEQDyiVSrnHfa6DnLNen0xqgDuHY+o7f4dbLv
rYkCvPl6oNbJc+77ZP0yhxoT1rggGXUQOJbTRrS6UhaZPawgnyHGIJtowweA
5dR+HLF1ftRydw8qfcWPOr7qrwxTz5IP/ZeLTK51M8jFBaVSwaKLOk3T8YNV
yXNj5R8ZY7Ng02TOS0OMjqa1G2iBBGJCZTYT8bU1I3bM+BhcDfQmUxBaql5+
oyhot+iNWC/l4nHSBEUX3kDxkWcVELQufVe7TgajvvX87KL49TFfxGV/+Jj7
NXAyhPs18ap8+FURrVXdNxvn7hMC2SfVtAiBOaY8xgXdUwzHdkf+9n/SSOOA
F4rsnlRxvPhcNN/JenMpWSrTUhPUMuWPaimZ3JPwpYo2PoUPC9jzNzbrjFJk
p81201FnP/10r37iUBmcf9goOaLPuz68dMpKs+kEz41iPS+uLacAA83gw5Ki
uUiwA+YU4b4KIeY6LUahNDLYRY3GN/seQo+izrhZ0/UwxnWCfZpP8uv8Qh58
QuhWVuocW2tA1hw/H5/b+l8QASkALnbQbhCVhnxJNHWRTJaOq04i19M9t1UA
A0Ax3dlOG0Ky3adaAuYifYpIWf2gHbHg0Qy48v4XB9Rw/KT0E/1dAmvCxMKG
3eTto7+uBJtdn2Ky3hDjxJm4OwFuUxRmlTziUqzfNk3FsvYgrpLbwZG6xsqw
9VD1eN5YCaoN2YIyw65PQk4+rWDOQDezTXc5Yqi5z0SdBcxejEic1QV6w/Q5
8YbDMwMMOXndmT2C3j4WXF9yN3oGogsMHiPtWCatAB4Z4aAQpACHnGJi0Qyy
00eUCuBJzxJP/3d55/CqZJ2kbiC72pFZChv2Dz6zXQpDg9WR3/4j4/SwvViz
wDHpP3R/YOpRz1OeMZGoBtWt2xW23l325rpWfaatzTFcFBkDRktW26nd9Yck
advrXnBDCn1Ke7a9Od2Bn/2y6nn3oCkPQx3FTHDiCGY+cZBz6LqZaAHEXnIw
MJDB7Ja7rdIKsxYrW1+z8IPu9KxZQ6Sqpu8YdFBMxgTYhLXYzU1sGY8gMtRS
Sb0rwdL9gfxMO2goER4js21uIJFoyGzg20/Cn/OMJq8pFRASdEb0kt8TMJeg
YrTjed9E+gTfwMhmXZIxX+Yqwqt2UqS9yWH0g/6hWu8X2mKhKlLScHlCHG53
UtgxulqvtOMAxZEaBTaBPrXeM9COIB2CBHzssLrzaPOO1JDjNIyWytoLbXwG
Pq/S1Vq0/tRaYg6JlEiyZNBEUykmbrybvzpSZiaTO2FRil3Q1UgBHHK3tCRe
X+7iJ6C5SIiFuyKomz+FnlfNp1vE8oAbpXEg7/WvcdHf8vmNC93S56M3WURN
f2SgOkMPcZQ+EozHbvtUAjR7zD63UBBp7g/RqJyvPqJTnZ/7ji7pRd1vAGJa
PgUVbLvwD51QU42goQFmnAGmO3iIAsUSFZvGuT+vYHZOR8KI1A81Y8rkqQ6n
0DGrGiwxBRDYFw2QAt1RJEYDoqIIM8OuHItlGGRiXx1FazOvztqAUfKIT6yJ
6nOtSx889n6aPD+YyhBtUVGedy/Q+QVJN5irE2euMv5qq9rChKT8rmri/vXO
//z4KkLVl4SUH4/qak+i5/Hr7OKHmZZgqrjisZwfmWipj01HgTkEf+1J5pIR
4+gUVBPbsKJ+0/CuCAgIrZ6ZrhNTDW6Xnxh79Y8I0Hr3a+SfEhBxk61W6qTI
HWIL0Xt2Yd8jBrDZiqLUoJAQG+5/Wk4m7S61/v357QVkoPslpDlV2ySpZEDT
aXzdm0EphDGlCtJZeYumk9ARVl2zsN0f+9VuXHlAP471mVJNMO1MZtnY9fSq
nOrN1xai8AJoOvBlIbplMYCBfIiCAKmYQJM1qDTu5ixM9im4ptz3s7d30lRL
Wuxl6/S9FycmPDK2iHZb0Gf+Fp0WpoVjiFiLSKYrQhDM/PwXWk0Yi6yK25L2
o1DxxSXDMmOuPvxNev2FXa1u1ZnyIKvnkPJsEk+WGjpVFiPRr9QQZa0jPnSX
R2DiDCFT8W0C2r8UB5V9J10LA6j9eMwy7MCRKg7Dw6uCvngvAtF0tdQbCW+o
jbMG1HU44DxTJhpVJxr02IYKNtp/OvAv/a/WwgyFx5xsCrya6mWNcqAwb140
JWqAoN+xxPbHZ0Oclg2IG2X7p7srENlAcl3JSiG2GvHyrGK7EWWTFMhqoJyL
vF6trbTWvPf9UzMGeFmqqPTQoeBcMbTcXLEPBEnm58caOMgcwhQ8WJm55ZFk
T1Uy8uEQFOmIiUHjgDNlWHSIsmBIZ92tHkM02WWgRzOi5/wk9LGAvURBgNEa
AVuuvXhsn3LxKuOl/IyciSvCZ2GzMN+8S93K2DS/ssizQe1pGSiwcelEdXGe
mYBRD9Z4lpTDwBpS7BL/KyqHDahBf9/VO1BxpyhnqOslSu4sj3Ric9DjubhV
DA62SIqbgNSQ7T18Pdy9joyMqhu+o2IWoG8bA5id5XcEgKBTrqg9GUfYbNS6
i5+9Z5cKEsYUyGQCETXDxHbQspmXMewoDMzeIqJebrsP50lDc/zyztIyVRea
KZyBHG1la9hsXpBtIB8uBH+025rBo/i1s6YEQYt+xUebEgQt6daqJTN4gnbh
v4GAc1hIGDGP4KWUNw0puDPp8NIwroU7dl2U828dg2lH0xhGDlAnUEWY/xXJ
g3IqP/KHF+ofuWeESMtcG2xGKt2HC1RGMvImsf/Fp1IxOuPuKXkVayBmO3TX
/hHL3N9vo0uySM2jKktxDHB3yVrWZzLOXeLY1VBzVsTBzpVLPjx9WL93Jggu
ebQBw3Vpmd8xZ0er79Xa+qESSS1P2rUMkU1hNh2v53b+tOiTfh81H2QM+IDX
PSOWB2zyb/eNI2/NHpMIFmoqqMfAsZWRldLgTg2haOn/C6nmKN0evX5YVsfJ
e0A1FXD02+YJh7/V1hoj49Zvxw54NUHLZL9MMpDej6GOzSYNaDvKFGBnmJEh
05MmjVW6h+ZKNbXvGlBkTTvPFN8NiDitwIluAN4An7OVRDp612g2JQoNv3yR
kc7A9Wt1nkzQUkO9ZK8GsqlnxNttGle6AWscom9Qij3UQl1+YQpIz+JUlc6r
bJUUUxusjzoa/RmH1nUWgfh1vpexZ+vOAibvPTVvA0mQtWqY/l2TnqbJifXw
I4RYU/1oWgsah+JUVHDatgGBzZhWYQ0lkZzUVaNZISANxMYR+u4oHQddOAjk
66JxbVpMTHzdUwa8IegQEnWO6S04sZ7di93qR+Tz4d1FBwLV/DJaxeG6FsOB
Nt3O/ulbI/GGs/GHSm6ZLFGOx2/bp3DNRzb52UZuG6xsIhFQhmLg85FbRrcX
NutQteneWkAHlri3vRJZytAASM6uiUv2A5ZSmJq1HktZTSCMRDNPig4lLbB5
wj/mRmHjQzS3vM+u33JgEXbeXh4qV3guCyLpN/rEBn+F9qJyu4brRRLO6sUy
eiq8O7WxQ76S/05kr9+4Z5NWF8OWdqZXam7seYAcVlBXZtsqYsweGHnzQY8V
n9rJuHxvnEUT0Asuix6hxthDiO8BbV5Zpq2YHpULOurWxmLCGQaKWu7gpNXc
cYFTKtJk/DhNSz3G859rGkGu/4pWGwNR4AC0kb2DUyJhKXRpvlau+PK0meeS
Evg7+cg05MC8JGN0F5UgfKeMVyN8mZ2Km0HzTbsHCbtxTM/t/C2aEvrxzCZX
EGBBSjHrIbX966G9vnSTstyEhm2PAE1qWusQCX1KALkEEtJldr8i6d5sKQif
WNofNTfPxS6bm0RoqeRGnKxslsTgR9o+pXid2LIvksIXTs29x5ENWuJlg3Y1
9k4xIBz7rdn8jy+hl7eJY0R6+wAm7HufW+vTRAaLoxkpNeHHNeYYVB6f7CoQ
UTB7fX+E1FDaI8/KnrH2fxoQ81gxC/NrSMiLtN8D3xvYp1W2ynwO65uN4vJ4
l0SOZR1FHWFq49fKO7JI6cKLQbP6F9B/61sjdEG2y3O7BABdQ6QXX+OWO51q
Xc6n10Fg3E7yJI8lTOxVqhGQ4/+TlQEhxtvUDnjlw6mn26T0x61hPNqQv3By
L2mMP4HDEb92sy+yfKqaPwIshgmah8zfSA5CEMav55yNGFzJFoRt7PpE6LAZ
+UIu+sAs4nW3kT6ZrHt7CXzNqzBvS95KoADeXHVInwidqIZisWoK1vLwngNO
/sG3/8nMyQtcEWjCJCSv80d5H6oMFIpzRTXKIQq+N4I3BR5DDqbXOzcePy6s
/nC6ihrYp7c+UEBlM7AkfEvATGA+7GLG+AHnjK/8vJSmmsgyH9xbAsM3OacZ
HZruTmx+3AfX5mbh0qXyJBdLOlh/HeHhNqvMOQzkOX2r3wDRvIqQqw50C4kg
GICVmyP5oSRWkoXexuijXoOBaOLXrXd3TtEnrOrzJ3mmO1v5ulixSFDzWfld
JPXCU3S0E2XPRhzV6JdxD3OaqBlE7XxTrpU0DhxpGRKHzlY3uAoNkqa1n55w
GVc8wCAt8s/5n3EvtWAPVlCCEZHgjehqmIAxVX6/dytlWda7rrQj2wfBeeXt
EJCwIJ1LSVJBQzgu0NrTqZwJc/mCNWvxl5yaEYaiydS063HZoGWfIoFXxV7S
6nsFjfB51p30rDFjK2FpiPNwn8wWkvr2ZZhyyKsy2t/m6E4AVZgziM81wYQM
TtAkOHzA1M1qthX9iiJCqhLsD8Yi5ugkNJkmcl9Kv6vmqt8nm8yWgMJ4a3rV
EXRlUAoa46yzsiiCGRSgEolJT7hHI+ldlskIk50R+kGd7/hGSeIpetfxvEAM
6Uq9qvSQBn/hU1uqW74mUM4twAqOAFwW8miQJlRzLAVsPN7192PAMVt4P6Pv
A3TgPSVcodbtgVs5ZaBeSElyRydCrxYOCqyzwfmpLjj09mXeAnriIDQP4q1z
zjq+0a0OMQhmRyuBfAcL+ryakTlIbdPy1pVQbAX8dR9J62Avw1P7mqGz7K5r
MiXhTbWH2zfg0g4FpWS0o4eaHA/o9Zs0pGHZn4ks3fyPGlZgG5hxxdotO2Sp
L08jNtMULckZI7t8xXLwBrBAInB3GM01sU9ZQwTIgoJ7+HxFYgX+vMEAxz98
jCjR2D7UPXDeQISNTKJaTDm4fiw7NpdpxB2fApoq0Jx7d83zbZxbsTdkJYPE
lFUHLoNWIPX88Lzm56cKBI1TIGFzcY2ZWjlqbWQcT/GZkDedq4YMiz9WHRtX
le/gfbKsJtIW2Ypvifg/iODLzYHuKU+4OmjTuBtOa0HbouWs1FXYLjnFumY/
L2yRIhTP7kyY+kf9KziSzSPKKEQrbBBDAzfKlW0O6sMazMcWzA5JRWLCd83e
vWGsAzfu37pb3R4e83z7ECivu676wjo4DXYzlJTITUke7WxTTo2lO8OOj7Zv
VmnsIHqrAuA/HPnhulK6GoXfWtesOoOjJt90J+b8z6ttVEG3x7CRNnMAqLGw
ASBFZ5c2yqthq2WW+SF8YbkPXFOR1r+KDMR5d2d6lIEFYtJ0yG7E+ZCts+KA
jKo+bfYWevhbYiBNqU4Af1eUDgPczcROh3XRbcQHEuMw4H5XL+NV8PSdrUpj
knArEZk0WD7hMQn6bKA5XDa38YSBsAiySsMQviwdeAvuROdm2DZVQAQvHwdO
ZWkKYEUMEF4MHpL6E2HrLzCoZGeZUujgjta6id1R7b9+YIcjtotiGlWhcFJg
m39sUhHcQir4neeIopOGYQvoWNg7CwGnmpkuWzAif/17Wd2iVpjv9SD5IOfu
CrfzjDtBeM/AjcTRoLobzztEPFB6q2nLJWPvnsJQOrbw3qo+dgxswW5rHAVO
lRYSn5/1QvmjBxqjeqICbjVtvU2OKQkYXAzFHS1k7ptJaxXkXkwJot5+41Dv
32JpTCenu9pLPRizt+VWmyLcgBc86qi/MXK+2Mbh+i5xIS1H1YjxlcPLaixt
9TWYRGCmwlHBcNMMxoukF87a8jVKXSM0TEEToMeSxO9PbCNlZ6Ck7pLFnJgZ
F4GCRNfC99OtrQQtR5Sqogx49eEhKJEecy2BpK9amliY3NXul5oPrrL7RV81
/TYDcTpRoWO8HpDbr1qcPE+IKjIegi1Jv8P898CC83fon3a8HnsdhhBlySxe
vg166/SpFB/IKSlnDLGGvnF9sEg0F8TK9ZhI5b7sccQOiptzBwOTTUgq+o5w
HzD9kP0973zQP0uRp2eq5T14qRDsmoSWm/yFTk9ptC9I3DQ64GTncKQJ7ulV
Wzuwzn2ti2tV5+A1MFDLQzFm3k2kNf7wBmFJNN5T4KD6QFE/K/XZRbSkJhP3
RCIG1Lr4brsp+5qAygnzrdzYs5LD0Tk7HpJGlDalYfERlLZXFznwOpYP1+Rf
+RZYqSc2k2Md0m8kf+7XeC+MXu2KZwMnlDBYEcfgck0Iu9p06T5Hu3A6liYr
9mTldPMMl5O+lSk7nc0CWppyyn6fpVVoHKrPbgNfbanXTEe/RNkk4l73pHqJ
aptf/GKF+DrNJ3KvOoXFLrUgeRg/p5jn7jgiQfGTIFo9TYpi05BiBSXGzb5k
O1fsZckY51JrvqddyymEan0+GKkI4+foDj354o+XJSZa85W8kT2BMucNIYTt
9cnvJSXWzVR/+RBkAGpWJFhRFeRgxeUEoGIK3gsSWx1lhXlB+3z7pfIy/tPD
G8S8BQojqmXpNluZCONtyCVL9GB7ZDX71PHxj0cic1EJGozn/+xZYQM5iMn9
QjuzMvsRElvlttWurTAb0EJKuT89J2Xq9YxUfeMr6XB10PM4G1jIVLy3uRpV
0PAWGDK0xVsMJoZuXV2VPV7v4Uzft1qe194i0Jg0CcARvmVi2Jw5Dh5Xz8Hr
BLfFqquyG2c0hr7p4bQaBh1nrHb5TKTxL+6gvFMUBRPHdxZN7KhPW9/wgf3v
3ftuwNJxMorhHTq09BeGrSDzUdMor2QzfRiMgpdWkO8sgYGyunyP8WCuWgKm
jGiUUYx8tYB2rE+HI4dE+q3Zvt8SiDwBCKo/LoggAHw//L+JKOcy0+Z+T1Rl
z/JsJISorxP8aAecrKrJBhM2GUVmX0tAFg2kPPHYGcc1qWmwSc2R5muJcFk7
7BwA5gYutQ/8/ZTuEQ+Bg0OZIrtS1/O5ehWdSWca2f/HPHg9OxGJAotr2FiT
Mr7d1mW0rv7U8z83qxSoxPoiTbxB5J7T5yZ444FO/gUBl45KVHUBmNICH3WY
RDoclqufL6bzf3tUvUBbhgVzbe4ChuxRj8jE3SOJ8otM55TihS19GxKQB/Q1
GRalFufTB9DUDPhaRzzRrHanWJIDQnM4Rf7EOpWFjjpZdy9pf19v0yzP3rMI
ZiLofVPozh1y3vkMeSydQ7ulC14kRKtBsHx5NcMLZXOGSc2EQLHuezwX4L/l
zmWeUA8vxDGLZd9Eu/fJcOyHrs3MqyUmDFlX6RxPTEh/CkiCQUgOV45IK2g5
Z2jcg/6+rLCCn5Mi4AJohPrM0QgJ7V7LiEkB0WJurt5T2/AX+cAISbpl4aS6
Czp31NPXRHFLJO+vmT+qnMWOKul73xvF/kmlcTkcOyI0q4DpqmQljKT3wqo1
hRof+sX8yN8aF+R9aDTd+6BRn5Xr8XM1jLtgastRPLkOxs9j3dDDeoWLMhS0
jR5a5L//393FwOCrptNsmdw5TBBFPXLTDwXK9EY6JlidKWt2f5b5nUTSgDst
oiNRSorCRAQkD8JKmxDNnv2hjoDOPUzniIjlrgQkRZCrzefTXet7wPiehHlf
XHOOWIHOzEKO3kN38OFKrnCYVeUzXZpohnVJChbB9AJYCAkckjQMSzvL7Dob
Do4AmLo27fQrix2foxi491YgFKjIPUySr9ORuHvllCFyUo/ytDSKGL1G9d88
Ddcucd6KmDlvjVNcZXCAczK32L31PPeqOHBWJ94H7dwu8F/DwsLEKbBaxVYQ
DJd412+iuDHPr9S8nTFDQHC++E4khFPQAaI+Bx44Zcm+KNvD0TRG+XZqKotq
JnfxCjxuaZVO1T8+1Ny1oo6tyuUHmaKC7qnolN9VwKtacly4s9ACVTV2LtFu
ODlbLznrU6utN902ZYMIGhsWXrB9AGjcoN/PCWD2ppv+sdwk87C1UomnYHqY
5mpyvwLVaAeiCZ4Oky0/rkbTEHD42u2/Q0VhtD3Z4kqMBCsV9Uz71GgHMcWj
HU4OfsdTC2PgXcUMLzgriOFk9GW7RpO1vNA+6GI1y0M46tfA5yV+WGwC/pkn
gP71SkFC5SeynH6nCab1XWr7Vf/X5NLVgO/0y3nWlUbpM2V1MPZGchSvutHm
oNPszzemZWbfX6YfGfoGDY6zPmdYZRXhFUlZ/ql0Q0VHgGWWEuoROo3ouTqe
D/BUUMwZ9TFgwCCerfbfTz9ZVmqgmQhHByhlo2c/4wzjKuhVPVWUx+HILnRU
P4p153whPsT3A9pOUKe2T2Nb9ePc1hCynYhc8WsvcYEYu0Dkr8XMw0nqpCdi
gsfbga6M7hTx3/Lhe5sVvkmybWFqdGaR+AykbX8aAJZZaJA1H9n9+Bv8BEGM
ZqgKkwGf+VYZurp4olr18RlSs+28GDG+P3BIzAJATps2VBkthvEtJe3dhOOz
9g3LXQN7XQlsvYl7VPw5jbAJMglLPzj1/7DFR2uW9+U/obPQVfWtKVr9vl/X
HDYinPrbeAPRxAau5siEGygiQCdNYjaoPG6M4VlH3H8jsSDwdUg+eQhFnk65
ziIFBJ350hi5kbdOnEtHbZwXmXdTWG5tCMbcI7Maz5PF1d2XpSRSqZqo+r9l
1wKwV/3bkqJNWjkTeYeXDwROiXgcCcMUfAAOn9tXxH89R5P6CCVwv2udNahr
S6tc4cDuiLdzvI3iEMMIRQxU4UsOFFnJqa0XVyNKYiQEZQBBKbtDbMVQjttS
J8J/S7qQaqFFSLy8+vcV3ddte37MN+HevN/7c3nzftQ67xTLce1Pxgov+PMf
Yl4/7iA4JnUO/HAN/wweqr7NV5NMCq58OT4fsec9a2GqsLNU4uEwFTzRyATZ
pllVeEzG/WkRzFsWDJI3yRoRAgg3+3RVzqdb8MyNFPtaa5gXLz3BxzBld48/
8DGggiZV5y0ttPcwHlrs3kS6TQTFzZvkFsE0xqytR2zOZ+lsEXIKDyBSxmGC
q1zZrM4tCJvidhW/wMt4V1vGNai5EmB4kmCSny0DWDr/aWaawPlrdNN0BnRO
ahMyIXAqswi+YEeTQPCDkE3xkXvHPLvXEiLd29pU7vHpPKJ+X7nrRdsMAezX
wBsQ5qVG7qo7TX71YgIM44zXF2ZYAGyeF8CsxOD/Lyx2vWUIS8fHwCWNBE+u
I5V9e02miTOgaO69SpfGlxGHsfJAgLj3R2RP5KyP3wPxWt2IKQdNZn/vfoUi
UE5N95BpKgCQOveGWDaup9g9O7lNmp9T8B3Tus2h46MoBZ15eXMT1a2KjBAQ
oMMbEp/0K7e93BdgfBW8uouvvEuHd6LYp45PaPDu0YmRFeTO1HULB5oFAwus
9WslKuz2hewxdVAw5IS/lcUDyldMfl45drE2JtFaDNvbO05r4B3TQnVoov4D
o3AVfT/mdDFdZ+j7A4R6IVLU5Axhu9gZ6Xw9fK1gJoBuhJJNGDWHQ0tw7Zt3
759qkSx5C6iYlLrKphKtqVIQu/BZAzBrtu6h1n9jbuNwTz56uMTTVZoSsTl2
bMFtsjQtxnzPjRT4b6VhAzH1y+TIxSpJRYqu90r8ZrWFvzdYzy87ae5IkwlR
NvxEg4wqAmU1tbMgVXEFLLo1wiZGcZNQhmmoq9GM/QLhj+knP0asAIodHBar
9vy60Ikr8scHJE1WIlgkYiY5W5QXg61y2n0OiwkDI/f2t42uP8+dbN6fLkah
3xs9Ft40MW8wTKLoItyiESEbngIkNip7Dm9jGT9EvgQxkwXUSBpND8lGmxTP
6EVhU8rxo1X5JI18l28fHfYReRKUL+6nY4kY00p3Lfza+PxLqV9oS1v7THVV
JabWzaCCP9BmkCFefQKL1HDNxzFyMfg5BNI/dessDYQMY/A5VFgZSi1mBhzA
YFMA7e2iuZb2sneOtprY53OxYygeo5stdPPKl4dw5zvYoPNW/57PPAlTCh/N
S0kDRnxyP+GPqx/Ji06UFW/sjffFJBn0oHGwSBQi/4jSmWyHdTBvqYm54SmM
lLdQSRt01JAo0kkcNuv22aWmdGNNQjicYYUe32zPuXeZa/ZP8ueW34DG7D84
BwxQRMno4LR4FClesTFFtzq/Uv0ygZs6SNJ6YOGk6sl3NMcnlx7MhhkoqTRf
9JHxtAbabiv85cc7KnlPPH58mr9UwjCO40DTZgtCvOs4eFvdAHq7BSDUL3RY
MvH/sqP37V0zqYCi6WAqniiFO37jK31PBvxnRqSUCxCVpuAn68B7nqSfBg+5
DS1qa5dKadr0Qm5LrrDKBxxgUpxI8qNPjgEp1rElQHPhVJci3GsLPEdl4bsG
NbV2oK6l2tqGHXsaX8HWudRPwEj7jembQZKAxdzSCLH7NBlCUUGAJ3sezprn
JvMSgqCseAaitOxXNGx+1vNy2i4SMdi7qisvEH0zRk+vdNwXgcEGF185Qqe9
cvu2ya8zAaXK2sKZjjpIxbVHH3kX2VLjCw8uOmpaGGNX67ZTAWAMD8ObF+s9
2DRAkaSSgvLv3KjBUW7yd0kb5tRj6lRt2oAqVgCveRXOslCnToWVG3f1pTIB
jg14OObnZyCr7nksW/+YsU1X2LgXE06/dM+k6LxWBnVVMhJiPOY0ANnkgwj0
mwkase1oheNb6w6sKoTDITbiXQiuTfd+UxhSs/hyjHIULl4SYb5ZRvqYSRAZ
uGfQXHQvqiuyi/KwbHNfMlGws6Cj55gZmL8RGTcym0TOUoemFR8qJHsp/XUI
Ty2HXR6sBNoN7nDWCWTijgGpCQT/qkxH1cgkD4Ot12KT1Luruu8Ue4ROfX9s
odxQPbfItVtwcekS1Cs2EO/DsTyan7MEf94ryH+DOjZG4ap9Mm5A21HwQpO5
3GQfIbeyk2A1dmSsiAqYGBdad0AWqHD3b2FpZR1eKRu4QvDnWdqhNKQ5tOuB
2RlC/NowCRG7hxTOsM3G5FXJw1NfUizL3gqvf1nBnujHK3KL787z1OboMIZU
MvJ4RlnfeU+YOyjZ7j9tZthI5QXbT9Pu/qvx9EPaHKRnlXSaAotxzjvakTPQ
0l27F6iHzfhPXYZ5h1cYaW9RRE8WhD8hWG5Hzer2V0y1T4f9JaJIBhWyvOvl
MGtbvLLZOqXmQurf/BWct1a/B8T+46JQ0x690xJmiORd6wlrtfMWrcrnPzPq
lUDAEbsVaa/bGukHv5TYZAAR5bJGzrbWzavqFs/SVnZWEXRPVqSlWJZulS81
XUhE0muLa2IE6kxJ02BbAeQ/cC5BfgarkkQkjvONtsuXeV8akhPC6AlvAbkb
DEA/UVdptUlX/XWg9yWbLfFjwgg8cG4BCJZ7uEc8aD+VpRJWcebe4/jkIznz
lDiK5RMb+mOdcYcJR/4LJDNwFPSYLdcY3xx0kb5hxdvvt0/q2/ZTpHhMYp1l
n/gkU/LmnPZqLIiGxdMz+0b5niDzQVVInDyM3QXuYgfQRPINZE1C0uuxdh1s
DcrGovXgOpuQlwDGs6ZaUJAYydIv9jDShiloEBbqqF76NEiqY/KhQLj37CCK
KWkIA8dK70+PLznC/XzkLQps+UBlDYSN17qZvSyavQbbBs9nNIyhRDLXAypH
+dyxtPJHk9lMwSwoh1Rt7L6I4W2DZY7Nzsay7Wy3+zEc07cIjLnz3F9fC6kt
dkB/dAOsooXItEo3tGgMGhhUibEnI1QxRAUJjB3DuGxeacrcDV09ZsHrYTpk
XnxBmWtWd3/zgGfuYW86hJgS3gSAdoEKV+SDaC91ScYH1wjth5e0fofA4DLk
kX0FK5yLkbP8V1wKxFEwMdy+vEsPI42BAHGYaUkrEYpJf8UuaGP6IRpmjTRv
ad1CEiF/4WORyZ6YsaNT+OQ18lKSSem4pMpd0VT+tYX69693wU50qFSzcshg
Oh3tnNxbRE01PJxL5piKs0076G59DGeHylRUFzZJKbDT7ssUuC71ZvGm5QlT
w4jKcRJcT03XNefIuOg9TnIR2cbrYLyobWmIzwp0/koW+b4RgVBRGMF4j4eQ
zahKb2ceS8Mdnp7IQ3KxOlwZ4HhgxcNkKJNWezGH2HRRWkNHwILPv34wnW4C
C7xtFaTVWVzVeQePUlsKB3aVZlltsr+eJ3SssFLkrQjpEL4LuEtzwHwqmYBS
cq3qiEPsmiKi/X0J47bjoXK7b7h866/Bi5DFfr1GMIRgxtacyKAQ7aiyDnem
Y1AmGsGqIsCzlvN9pGsk84i6sPs3jF76W/FBd0lqhMNDqkdWkSU6XNUYFsaG
dGgZjK8nR3mEBPtiTqzePVkX0Hj2nMP9hgPoFJsWiQdBuv+iooCzbEzySDZE
Ne6b+3e/SVvHXKlAX+ofA3OlFcat7+yrCuzXU7HthlfRVdHnZ0ECmmWnRnsx
mtFDyWw979K1aJyh7wyz2Ao66hAAYVtAxg3mYoe20aUcZ1c7tU0I5h/L/Rgz
i1bZ6LD6MzGz86p/R/r5yryOP/vM/Q64O44lmypQh/FGUVN+DqjSxNHL8mua
/sjSistdqgx/GKvb2DxnF4Kz6IGrKpC0pqLaoL1PsB4M/XY6yWtQ/m5du/2l
4N43HNTUO2YpxI/NihpSsM6giDg1sVJbYkgvLezTg7ZXXqQtIbSkHkQbVePJ
p8BwBPfNsmbAsFjW58pziqAPQFTv8GjHEgA351GR6Jo69RYzgqiSngEhCGc8
C9VLxW8535W96jNivXM/iAcVZwUQ1D3u6JQvekjmzjzFqklPk5VNVtIu25XH
xf4acYIhUKphj5w/pB/JFrtROZSEZXgA6PzHdJhvUNOJgGOM67vuFUugrvUb
eFZIc1G8CvbYxbm3W3L+7veC8A7nWmhY3N+JTxMKxkAHJlnhgAZ/7IYPkaBD
ZyxNm+nwc+rokvA8XGOPzL88Z7LbmaAdzkN778DUImscEjdW5s7tY15vNdC7
+2fxXK75ELw4oFyKYbHl/YNwXlXREpYR4NLRRKB9+JGjQRJYEyz0FDuUBXdz
YACBfDuOJGIJrYHqz5lh4XGg2tJjs3LRUD5NZGvtp4TzbB8+V2p94l0vyPwr
lUNmGIWSsdoLCzW6JPYo6dZDSakCFZTNuBO2+EeBotgJgV5FxKFMRm6Fy9E6
AAyYbIh72FlP9Xd/pL8vV6zhJQ2yoevxJQCncA/lQGVLIPNIXyFdsZeEaxBg
Q7rRToQq1lx1p77m5Wh5qibeng5xSoevavHrzvdtlVZIGEYDq0fcJwjgwWlT
5Q4d7gOOUc7ZLhoeEeoaoRPVXm/EBfAZEqO9S1r5kAuiCs6yRrJQ0SvGPBtC
zZbBpmhEeiyhPZBPh1QU5n68gQmnvk34JBhL2i0dUZWG1UulxjTDROyQAfmZ
kiesdeBwxuWHnBELHxcgjVxa+HnTWuicniCuiVh7TfnR2ph4qCNwEAQQRJF4
GeVqkcMdYCOpCt+l5F7g2rZB2aS/EW3GWkdzmg+fUT3BljZlGZ0PPrBXm2Of
ANth3Bl1RxwmVIhv4MC56fdDR0fJpK6u4zVKRL7v+RvaSVbFEXLGAYJPpGh8
bNBN8Nl+qI+2qV+x2J/R08wW1eLTmk7odDcax+zBj3L8YtG87L1bZv+wT3Db
5ZJi7o1yROLrlFdLughVmBwgUQ2bfTJNa6+IW1fhQPegMXA6nysEV118dWeb
VGQdcpsaj0H0bumCI1ISuNZOunevcjCTnR5OrOUCBr7xs/Rk3MUn/4yLp7s0
S1q6yk4cPBY6tLMfihh7gBL56+k9X8s4kGbnMTPNvUFekUVr5VLhLkn8fHqd
1yp4ZSgOF9ZKz98A4sHrekGenjkgVfbu+Bq+2BC8sJRxem0kXSFEGcVlr5/j
8dWVQJxATehT+KN/g/7GS4vb44rXbjsvVl5lhxxP01mzrGt7akV6VO9Osy3b
K8LWJLJ69MoLmSpc4ItkLwZOUbuIKxSvkLDiEr87mOlNnfvf4yio8SdgSIf9
s6fpinHvGJuqJHboj2tkLkj209OgU66xVPrBRpAE/V9FP+M5uwyEPcWtAGyq
Lu2Qp+fBSSUPFLqLlsoDnRlC4h3yQ64KvyparTZG8vjO3WoRmJMYiVjGnm7O
3JUMEcug9Hgv9V8XfBR4ymcP0J0poWrGJwRT07uHo9zxlm8wO/+0aYUK37ju
DoV19+KdOOSIMo8XYCZrE+qeq97y1iNPs4oE7dwPFyqAnL2hol0r0VIGdiQL
GWwn0qlN3aa7dXkCly98qVvnZPiTIHz+bLF58+0bLQgpmK7WQrxF3JExd6h4
1HYU+qGnO2vY2autnZCf2D9GCtdhXtNjNBmKGae3r+jX9Z7l0Ter3a/UCEqk
BM94h4sDNzsu6rgl/KPSqOqDdQ2cyCgNqDT49dli4ifRGcpd6HhmUmNfx1IC
HvKCyGviWSCg6KDJIBTLtxPU9GliU/jZLa3ZHbAMoBRTRp1GXDpWChDbEdNh
cNVMXFRdTqeMu+2ZfTw/45zmUK9g/ZMbrMi+kFkUbrGotbYLJ58DxbbKOMzN
ph9pLO2wEL6ZYEjZOUfUGGzto4Vx/F+xte0VJXJ0DO2rKSR89rDoqHIcEebo
T2TVhEtPMBsUGkpZbH+vI2kMFYgwKRcW8vPdNd5moG/+PzNGTp4QV1fsAuJr
iuehCcJZzotwaUCKEr8F0+icW2bXONgUofygNett9uW4ggfldwPnj2r6x2+n
hITqLp4JeMJRfHWnvEOwi5/gAwr/oXr41SSjWtnqn8e6shTVNTUdYiNC/GLc
MLUAMmvvUz5LrDsBKEMMbhDBkMhMEQSe+AtdPsvZ0/Aq/Eqt4rx8sYqHODLp
AEh3HqYR/F5WOVEHEj0W6HBGV4igo/illc5abo20WhC3H1ZQPM3DGuJQSc/l
DK9fTTWbXsYVYOZy1KVjWasONn++h2Ze3cMbjDz+NoEt6pd3wA0vpS4cQxou
bsGj/2diSpbwmTyHw+alLCzvVYlrkKt7HfplcTztlAn6+hN4MSFWdnDxjgiw
hw5x9fFTD3vL7ToqgwV0hIty7HwTLktjt5vu+Cu27FZu5xhHbcKrcyFBt4Ff
JFgboc6PiFp0l9muFirPP7YxlBL93svXUlIV4E976Dr0nsihvjxr4wRfX9Xx
cLDpUSujMq0vi/+Nqp09LYTASRmU8kCylSMKJwEl1csabV4BBizn3BvxOBjM
D+8bhUBf73pnXXr0LRumgdoJQMrJYnikDchkEim4iXBJiJ0MrJeCfaQfQ+BC
F+cKAzFGydO3x6CUEc1HNaDVQCQU1sDTR6j2px3QPY0cM5rGxsC/114YHUiH
JFrTMCyJlywiMoA4phTN09ykS5Ra/L3U/l0fwFOoTaofPpz6GCObBZba1nLf
i+VUi2qjC7Y/f9g/jZMzQPItsu6AzsvbpcFG8RiV36/BXyMDwiScW6MRCEOi
rbkQcVkkckj47PLFBCw/RvY02ktgHYjZVpKHfwjKdjb3PdQwv6CbDbtk/GUI
TXQviAleyA81lKEF1VFka52KzqQ44VP7R6pOqHTV6eT/LOVuusNz/KXO0sbW
CsGv0EGABhNcHLl0iLmjs4qMP3bLxqOXeqhYIPkRhNzaT0I/i/1h/6bkA8kp
soBGJsMkf6ReQJIb4TpEGqLXrvwFw9eGKhpI7O+gVrB9dnjrl7R9myH0wvLU
5LG5ICCWOpEJQZLITtjMewfLjR68ELFh0Cv6wHRHSsBX17SThdlvE2420Fih
3/ZiNQd/WDQN4X1bd84ZSBiN3SltyJ1N5ppgUtXUk78BnMQIBCtXh6bA1qOG
RkTsD7N3cnTfiSXWP8/87Y4ZegEwgNEgr2UAN5pXSzcJ2s9ZP9e0wP13EYLh
BytfqXnBnKGw813fu+sHv8RPefT5786s8Ce73kNfw3oKGuYrTTnuwgXKh0KB
7kwVcZ51mRpkTu5q0LIWBICZmYOJSRGIgC4W+unr5Dx8TLJc2Wf/LxckO8Z6
ltGvYkLLrkpwRFnPeH3LEQuGlBbi9QdfGClmcvaYSPZPKzPFdTGjbYAMLhcu
TGgZO/eHNvK3729fs8743VBvRPWWXtG97GudSkT1LkUAxOdsm9f6E5+LA7Lz
0SHOBXcZCayslJcVC65SWKxJ0QCvLFZDk0nvJZn6YNV1hvc6JUBlEj8q768n
EzgwDr29cw2yrYV0Ow2dcCUIwOzmMcMlEpvxJMqaFxfKQc2N0UfBbbVTlzgw
KoI+FD3F5MeTL9LG9pXsqQMowBwFG/QxR9fyOEAKW3VEsbu2nMlKLDujD18J
QR3lJBwvOOcFq+HCIOlN8+e+845mi9T9rgyZmwkbiHNzOrNxzlD3l23+Jkzx
/40WoVmAlTYNNguY5uFb8YjUxfAkTjIhS0vhpzHTlKUossWuFwaCiXLS8dXA
VXqaau5Q4TQwm0KJIgR0Ic/s03FGCQcjZPRP0ZhhqATqdPx64uZikXLTTzJg
1Yp/TR/WH8pTHuTFuU5K70MWLfz6j1KjX/By5FhuGwBeTTfifA0DSBUq2KLi
kcM3mKllafTA+rk/7E1QUPNPBPgDaWBOQN/8o/1t2PNI2BLQoqd/fh03SwFu
qrbkvBHDWNcsmpbdoxi8vvD2k6lS/M4JddUtIOYQsVLJo3AxQO+W0n5fwIN6
Sg3rAg5QQ+c1o5A/ig80tjvzZlEFpWgt99i/t34JZNI0jrGsjpy78hBGNrAW
2/aj6tppcxL+QRPFYxLg1raNcoKgz49NhCWewesryx5xqpNWHG1cTJNdTywP
0uFl99i0++Qm4dkW6xiAaEIPXHqwNpWOEG/hA/A/O6/pNyAw9MRBARP/gWeZ
n/pfiggnr+G5geU3xNEIcGT3h8+4JOgewdFXN4v5suaK6tpv05SGOodezcf8
SdUYqIN28UWOiaZ7QmOwTAt2362pz+cIp76UIFPR5paE9DbGiW9uhb3h4B/e
UaP0Jjxrz/zTdtyx1KPUQpC4AiruM1R6JigGZE2qbU7L1JPrqLTy3/kraEa1
CTp0LdSmnveo/hBz3/LPmR1E6BxS5YZbCC574+jWBNr8NnccwtT2ASwaobDX
wNgUtMKUC5KuEAUjlbj1wT9n9699cPDOOf1KQtcDi6gbxmV8OPVv5jQ4O95h
ED/RsPiX3hnEU5bMx8qjQQAaB9OI5bkZPkJ5Cqz12XbW6BlWHgIWVNDz3kkg
Ek0iaakahT+cFWSO8O/PWojjUwcQe+Y39TZKTbrvfnqKrvFOCwyDsbzbg8k/
Kn9e71j4Tz4B/JCtwSX62YaGAo4gh2UY8GLfl9PvRGYqJavnXhKleA1cuIdk
kytKFGCsUuQKVWyArIWubhuPcgBn8/dB+DpKndX71WA5LzPzcBb+3J7ddYN6
P2tgacOtNktf2hLegRDcOOpdv4wz90143iyGGgoiAKT8wDR5eSA8mdR5FZhq
a+LoLndcE6zJL5y+9XP7sp3qBLpVpBGNtMVTLYrUpNS1LXHBNpH3jC7jNZK8
JIcxCvtYlg2cXUf2g7f41qKMW4xBmhaeEvCvpXrefoOvzM/3YCFj5Kq4ys7e
DP6degzuYz5mMUzrhm7/xVXvg5a+KK0JcW9Tk4b8tHIyfyLP4SR3yBr3qTAk
P2lrXlE/5Foi36UmSoebBr8bFxQSJChKEu5yJ7SJyuYbu0gKlokvCJJb98uG
2shcorw7rvX9ZnQ8ufpzM84h85oFGw25njcxMbxhCCzJQaOazBFVnuAlzOQU
MmYDM9yeBOrwG86JHep6FM5H2FkVOQpHyhnLiAsP360HDznvm1ZLvL7/O91Q
56AgjgAFXBzrMA6KENIVDVcko3SvIIHARTGq5kM678MfqoairL977HKpsU/v
udEEakGwRAjdPAN1pglY66fzDqHIckzFsmBYrYJt81ZT4tSoudbVA7eWXXTd
uZZIcwgoG7o2dMfxmdWzcOSfhKjdqy4NRYSTvCB8GBuk8BfCToPF5Y3RWGVk
/UsMFtS189cKuVYvCqg5AIPCHOcMCYwpjtBUIE1OvWFPBqhIXDLNuQdFhPUL
JUyyqPBYmCY0Y69sC9rcvi2w8/g/U+JuSSBpr2GDWm+eUt1K9H9S8FBzo5D7
wFTdDkfFgiQ1uRmqtPx7S0Ox8oYlDoPYo3Z3ej0Bz7+l2HFzYLb532KSyLJx
s5d5nauIuqTfPfp/aeycAGF9iMd9dhaF3y/0Oc61CxVI0up5u1wJCODrAW9t
9+PAA2Lxj7YWq/0qvUSO0MTWf2R62i9R73Fo0Bn45ThQ2/mEC1Qk19jH89z+
f0wSle3BXopurIzD/W1HI0DEsr6HfldkUi1tI+iA6aXZg7/C8Vhf4ohqhqtk
8YkXEAa+GM9A1ip1JPb81D0TbPDLkQlTn8HuvNi3P7Snj0YcDmkX5CmXhXVM
T2eqvvmaB2BopgnLsvRnWhX1IsYlw6MoUID4xiFCMnrX4ogYn3iQ7Aid72O6
453voaT5dj2sGP0h9Cr16klhBSvV3CFDaC75nnXD9l+431RkfvsZJMJi1m26
rEe8o3SqBhWJPaahhqnGC36ziMIvpjA32CHxbkIEewapTn03xV2Pz8inHedZ
I5xYSMMCneKfCAvVxrR/Iu8pMXUgYz8DnY3QqLps8arbcASaN4GVusXDCpG2
/m4Hvg6vqpijVv0A2axiiu6/OHTh3xgrlJN7L9xpw9WlpoYgcj/n4bstqy76
fupJqAUioNVWANuRNzQj45xp4DJalEwV4Tc+lXAzaYRPzwaXQixE50uGz8A6
W9x8ou18gCw58fLysvFLQVtTsZhkUjto5oFwyCwmxrxiCM4JAJwcbpfHIe5D
ZuO2zF8KCtXcrEGd4PBrmA3/HLE9q6lOkjOm4X6fK8qBMeTMrTF8mBR5BEY0
pPbvh1l1OqIlCSxDdsmNaIXBWnWlXNU5+Iu7uV3DnUL8GrZdiq7bD8NInRpL
MIVLp2y2/ZD1JcppT/tTwpn5Gv3RQc4YahGtCAgjrzy7+uLpz7SLEba1BNhY
n2cfHBcLDW99jTNEYybbuBp3lvLfhjx/gQx37n89e0DcKnv1di5knqcdaZtq
OV97+PF+0lPRb6nnwIHcPpQRSC3PT4dBZT1CEhJUamVYrupbf2Jc6GPCGIHg
Xdy8tgBw/KGjmDbTrTOF6UlgzTpw1C4QwwhROPd7j8rD38VCvurS7TV0nXFc
DhEfyM6XucZapcq2lJw9hJvIoZ+U+6uDH9D+TpDi/Y2ubXyE6oVTrEMvugTZ
J2R2b6MYuoOu2yH8DrxLqPblORHBzXObtW0OnEocNCFrYceUeOhhbC8uJXVp
iJQEqDJnULEt6ugAaGq2C84bhkNV3/wCZc+t5uBqFpcWQ1SUvPP8U9LaIRQw
A7vMr+SHylhKOsxRGuqySPwM3X7wht5vjQRGvHAhfIiMmY4VwpGZ0x007uOf
CvtYaO4ALzswBZ58JhchxAeRmUbBllDXaH3I3WFwpe9VcqkIr7QfbncaOMXv
N0Vn4kfmxDeocjO5fjYJmn3WXp7IVq7FlEclfVVaFOIPQogkvm3eAsQX7RGX
5uBdwgAWnRU40TlOSZsNU/bEMXKePLSG6dXd2dFkCtsXw7lJ3m6CdGKpUOOw
Gh3HXvjOyKA84RRgyuGDesnK1SQh9rki1L+PS17IusdVxfLzfWyF9emH6HE4
5NQJAfanX62NclQAWMJMVyLP9s9KkjC9JVOHNf10A5rFW6dmiLp2ROn0j6mT
QkQHAUNU9SWbWYsGAcgsp7TF+6oXhtql5ZegaM+GwQqp/VE599tmZmcHvOXP
p9FHTeBQFDRA1rSu4UeOJyYGlM+q5ryfE9Yn7umPh7XEkQAMrPwJCNzVDJaA
QZlERjNGrid0D+qSNMIH4V9IQiL+GxoQLCxS9hiJ8+Y33pmN7IyEVI2r66i6
tFBzt4xBw5JadqBBgl186slzzAIKg41FAu8HhVk53+rx54VSz9nWroGEI6Th
Jx007HlDhiYliTbgsoO922JaOOwVYK0i+vF4P0SQLD6cFrveVYgoRVZ+tq4z
WIam+t/XgelgayLmu8Ut5sKBx8LijdNhEdus1TzSzizMVJ06KrsHn6OJHGo1
g7dduQRLvDzNCav90Jj4RCv1rVwMsTCnVH1CHImb80C8+mmWamwcobbYY7fo
/+R3gU7dx9SYUY1tFvZl72iy3P0ymHpkC6KjI7ytz5a96nfOtQW31VxvaHAo
Rf+fSvOmn/iHled41Emixtt4Y0HODK66NIRTKAw014Xbz5CoMfDVCI2vNaFK
s7CFa/aQHsFY1Jlf4vF5noqB+OvPuzLwWsU4c1+Zdi6+ybI8jDkV3HfTIK8n
plBgwLimo3MEcJyAywwQo1rEFbda2wJTbdwYHuOMwW5U9HrdHtsjiONmIgeq
kMO+rJ3EkVD0Vum4/3glBLjJJgFfSClluRPjjtZcZWxD4LBDBFCeU0x+MXEd
xHjrzTRE1Adj+xWNzWumBTvP0VmaIdRwRl8gaBSp90VwY4SVJSyugHqi4zrA
F98JxdkQRs+BR3XRFOnppKD6YFraxqTtjl56KzdaeKp3uGPp9URBKAEv4gzC
C7zIRJvcXfN13HfGTDzQDgly4D6JKXGU4AcIO3NB7+AYTtVSp8XzBNBnml4A
QUR0LAdIfu/kYpKtzqQ10kxCvkMI5Vc/AnTDLufUUio8+68/oj+L04v75+Cx
FiDlV3JPWek9F+QBTD/TUqSFSFa1oX4Kru34Z65+w7xed4ffUY+QVWUtvque
6IyeFSSCVFXYcptp55yNU/uL/25mR3MRY1xTBW6JQeAUtIvDJBA6VzC7tJge
8PD2x8HhZ7TfOUL2ErrK7s2EKhy9XIkWmPH23bSN6uaUXhFLZ9UWHKu68Upv
es3Ih3w/Ay6tYCchGbvNY08wlteDFZrTar6w6bvNhrQRpLN/Juu+7RTRryNl
6a6q23A8WJtYAC6qC+RUTBH8dV0DwRMIA1OFDWseZVyVhZxnW+xVl0cZoeOW
J9jBlwIkDQ7X+s1ygtFnebLyN8PvxEh1NjUky/wkMdxmJc5ZPW4m/VlOxiN9
TgSRYzyrh1P+ujFjxa7CEqugV/002Cdmub//mitkP+3XIv6dOCXTVgGOMRvU
cUWBTYyyf+KC653jzXRlIQe2aem63PF986J8IuqRMQNh2nHgBwJQKXMguRyn
Ku3Ehexi4y84F3fGCOCTMHQVfmqipNYbedt2O1YDo2ldXuc1DutepqlDz5KX
yS3ChBbGOped0o5BdyXvAZfUzNSb5ApFIUGoTi7NmD9OAqlFl5Shua1mU1Ev
25vGiXj/EMVfTyIqNVXgIqn4x2fHZmQKmjD65cnfNTgpXkAv++c8cFBzqptf
AmZq0VHNCA6b+Zls9yVgTRkNiFkOUJ+oKMUssBwpDE26JzVogcw4EnS4/ULq
2OuVGW0KUUu2R7veRwHZDZJN0g7bkvCgsMcTvIzmplYCYLqxR2Xcw/K44wnu
ubexW6/AkHI6Jv74XOk2ZYS3ga0reYN6rxHcreZuo0MN5tL+Dfpgieq5yWWS
Wt7Cm1UVI448ZZu5TG0iXJVNN8Aw0X22L+vH0ZPDaDpvb3NygQX/HE2IRRUN
H7bkKtWRQd4FdnNGrV42AhOPt0mBNk27pj5fm8dE5V7499H35rNwZiSwGDb4
oCSoWwXN6nCVAueDcIycCskrFzY6ISdTEEN3EtJrPAKe3lYdsepm92Yo0PsK
sRDNqFODfrYXNyPqeg/VaaldZ9Q/8fKPOgZvU0rhZydM3JvtQTXET2nT3KiO
ZPv8sbjh16T2iRYu0/Ry4tM7vP38q3ywPKBAzNXnqRLKaAgMuNQnKG09JL3f
K6cH+fnSKkBdq5SJxBZaMLqvc3x3GhBH812crq1LWw5rDHrQCQZyVURIutJY
HJjvlmsKS29TlFMlMqOMdtIE4RYq3C6qBic84t9CeMYAJuR8qf717ZNfUwld
LfxFbVbtQhs+w2JW8Q4UlKlwoHZZCijev4zNBbmHCOHbiMojMZEmerX5EgZ1
XAjPfYrfFbrvwij4TEnunl9M9ltieW3kLMgPnwAUnqJw1+4mXB4fu7na6SFT
oJyai3hVswKf2x+4btrJE2SSw+3i8+wznwgaYu2DmHWGfhj4xY/5WU0pdbnI
Af3k2vKA5GTsvg0qSFMQN3jof5A3egcGT67VnE6j2qq/RsIwr4ussij5ZPAc
sQY3OX8w2NNON2Cdd4wDb318Eo80Y0ZtzEI9W20ML6ZRQvyJXZ8MCbK06/og
AVxFT/q+ppQTWMYGuF7jKUTFGMKvngki5EscrG4T4XPZE+05VzQvkuhk9bNZ
GTUr/J16v9HukMfXT58igDHXVb13ZMisz7/e8/Kx5XXnW61D88kI6C1Ts0AH
sIjdPs6CYt6Ac0ucUo1cg4JWewJEXIsHe/cJDbd7PxNwbNAUPinSxM1Jc8tg
5n4HmmykWpcfItBvYrrhl3lHwl37wSRtSrdT76Rw4keY8s6dXyoDMlhNOUbV
SAMQ1cwiAzjiM6QV/3ayUJH8Q0sMKWhZW+tZF9OyDPRIZ9Nu55p8ePCpz97K
aPCjtWhZc9kY8oFyHf6VdcwVOtS8oBL1j2+KyymiJz4VN2ZIyJKlSwfbThO9
5VxhRgrXgDnsYnEcqahpduicAzVA4rHYY2IGxvXTlTjoPKHEOtrzdYaETZLL
gsx363Z2/pKzOtLF5J3+zQ+RwHPNPGBlRxaIVQAGfWD1wtv9G5iS0GtHRws7
B3Bw6AZeWmqkDiM7H0RkhNDFQNpE4VG1tthu/4+fKGkvcYh6A16A1wQ27nDd
tLUng98ZKI7+OcDB3pAJvz+UJ49Fu9wnKiDWP4F3XPPHU9sNX6CCaKJ8rv4J
GTsTOXwlUIB/enpblvLehWInXof2rigH3mqkEafFAR/GMj6GsM/BK91Gdoq/
1M2yue4Dm2lqK1u1GKS0h7qOBPDPFrw9WqDqfLYX6bHqgoatDWJ2/uW+nOja
9c5PbsvstdHmWVEtB6oaDKUNf4SAQcUgdaKXZlefQJcsb3j8nsCwmBuMy/Ja
jQSULwmZiYtxBe8dsJel4mDWY664RNWCCuDHFm/2rsaZaHB83mTMPFAXJ2Am
yqwnvF4Nu9DFR8GJEA9o7dPxLTPxeVWvvr4vt9WXLftLe7K+5YEsoZzJx2jy
PEhdGv6mmKzPczFjVdZ7u+fBhQQAaq0IKLp7WM+NZ4BjitJViBRF7QcxpyHI
TIjI1VeciHOzjw4nVwDe4iFiUx0zdZVHMxEP7s9By4WNMTjQ3fSm6p4fDKHU
Bc6PGFgHtHkHfDrVoOUR7IqRJ3oxwo5OdRrml4mutt0RS0Q/0faYDcTjlqPT
yw6sRsPwKWsy9FCTIjCJXqHlyRgLXbyyQfZcV7OBQhZ3Rx55ZruohKZ6kt8W
i9QNi+aYNZOaCzefJ3m9OTaTHHq1VupJ2bF+xw9NMUy6cFpE9vXvL69TiAIc
cEDLn9Va9acgP9BoODzHh6GtAeVzLAX+HCENDnmSNpvA+6Av8EmyDOfmYdL5
MwscotG+KBoqj+QGsyccOGCAwkt9v9dpomuHMl3x0HzjBGzgxJsI5dlSfFbs
lTdWxCyhnusb1P4bZeiEXnXaZTio6N0invpy2L8IzLiW0GzziJxQQ6b7Gjc7
AqdUZXNZh+H9lVWCMw/DpRNuqGv0Eaymj0Jyz8HsJoxUiak8azn2yNVS1gup
5IJKbHuiLol+158pGAysQiQ2wtMYtRnJSmfuVuVZrOgdJJmkBD0o71utPwYJ
GJs2jDQ1YDJR36pnatbnrKmqykn5o/3MVdxSX1pfqiPYoN/mqdLAdrRGg8ln
+Dlua9ZenXySMMP9AhF6o9aG8IX7UPT0IlHsjO1FeFy09OrX45FfdLf/8g+6
fQ9NyVMy9blA+36t0WUTaWJT2nAjjVGjpuxtNUzVBsoUEKSzG/3UpQ/J9XFY
PigYeRQqcEa6bEHabDHVN6oU/szA3KYWJZ2/NlEGIPzsHFEJlwT8XE89ZBWu
98jZ9aqbtUw1XZAzjfVcwj+qj/S2AmYAAziRPIkovIysF+DYXUCKcHYTG8CP
bLIgeSMogJVoqoR+aWdjwlOie1aCpfvns5sHGl9fEjFKlTm8Bt5BtrJQP/Sh
NGPIMcIjxdEEm4jA3NREtB74NVDqTRRDIMkhLvpaeq9Rb8dmXSKLroQGWW4B
2WmleQjhLYK6VBhjFP0E3jggOGHFlET/53LhsbKa2E8KeKW1H3G5z31iQIC2
sxva2cZZCeZOH9K56RuW6PkdVE8W1P3VucaRhtwPGhO1xGOINDtLxc99oFFQ
4FOVUI/zM5vaWalZSkxLs/XJGKCRJhoqaGOgCNvCKLPI2Wp+hXSnHXVgnWMP
2zoBebS0V7IuJAgLocHUgslGLdQJwpHLeH8FGOPbgL4uKm/QZE7qSGJ5MgyN
gnQvQs/NnaievF2E98s2V+dAR+j1kkBzvBpuFj11pp7O5OUx0d49ga7QKXPG
FfGBr5QUCFuGluy1Bnkd5vZiByWQ+RnWBDy6kQ1TWSWcQCdjIuWg5JNy7gM+
Z7WaxDcrRImYKKVqPSgdACNQl92gazoNfNCVAsxKSDHyqMJkaiBGP7j7pb5B
JsEJdjpKF5yhq71jHSNugQ3VpCW0/QLaVUQ/2JYDXbB1HfVeIAIrz0cLzUhE
3Odte2ne5V018Q4kKISkXePnGlBKgS02sSZ49rGRQ8ZmHlEZrOtraNThDNpZ
00GpKzKOsJgME/SUc2Hc8TEHOT5sRzaSX+zP/f7+Pcj2xxvl4tmuiW/Hh1Sh
ZNQrDdDamkgb76K2sI3JQb2KxgQTIsC9QTA8ZZtClpzLRerk6zOMj0fRAyqz
gEdbTFKKTheQCRIWbtlDdQeww9tJ/ax/zo6I6j5O4Oygq3X3hv2wSBYZoXiy
9xO8DR0tAxE/O+MUaEK1yp5EQ8+OKNBI61YHqpHRdehO3bD4Hhbh36Q1Lrdm
U0I51OFcuyEXMddRnBxkGoKHozLsbot9oARrfZM3j4St/PQNUiOFrNXMBNCK
yAIKJF61yXezzc3KC2yXPjReYQNuPDM723WyNAMQ0q6MjVRm3kFbE836gng/
yJ4HHRHG3puPA7yWTzFuT8KHOucHZ13916+mlfAkY6e/8KHL3fiSMrU/OQuD
M+sdh2lDHp9KjlYZbmMTJrH92n6TmveXvbQqkKNUaYOddUi8yDWl6JltIHb9
05xcbo4DpGqZ5pciuTsyUIVSxWDup46exyB7Zb7leeWWEhYRmGPQ6h1bkpK2
JHWCvsaY7zUY6W7/cdASR+TzOomkjok8JoU4+XxV903+jwxXcJKh7H7sRZoV
YV0runHcir2bEVnf8qVvheEBWtD+9qP8asUGkSQNPR0SEh6BUhQY6mu9X9wy
FGGdgTBwzriB2jBuhEPIeXXYw0UpVfUZksHXmu/eVqb8+nlX7/uFq17dKjP/
F/Che0+ecNIlp+t6+pYnnKkJLlOUL7swU85BGovcqfrEoGFWqpWTCu7Vw+9D
w9RNlNsyg/xEkoT9UgboFq0WwyYaoRxYitYMAvi1yNLM+NHKbSqB5ZvSVbxS
qb9Dgny1Ned6ls4iX5Okhiz35royiz0g+6FKJ8CJaWSKXg1vPYUcO7il0mRv
XqoVuBRLK33HKSdvVCuIywV8tyjFtCTkmyGJXn3hV9RhYWEbsUlCUDtzh3/U
5+0WoWCPuTwqPRJBt3iJkbqMg4oboiKfoXnLmfKrBYY3h25xQPeemfDEFpSx
77ZvS+o972gMnr6Kh0tcb/OYrPu3zdyES4ToCN+nYuJPD2EuxdvO/+kkNJVs
BkXKUTXtMwvlUfuDAAefdEoDBFxktKGzKbzQLUy4uS/6u1JEHQTDcUbrH8fk
LwiHf+2tFA/n2WmSHEgLOiv3m3pEi/2wIA69I3UVGivmqrxKMBSSCxWs79UY
qj0o+iUkB0f6A8J3HgO9hXtMxJlgTs1LNjr/YzPYosAIunrc4PEW+Y6dqES8
5vcGnAqpn0QOR+doCGD2roHXBy8VzHldpNcqIF78AvPa3XKu23BwpUeBo7Vj
rQcRIDGzgv94dORm8oO9FSRP9u9jmIL96uykJpbqE85liWn62YH+YxI8AHD7
/tcgOiQpw94xtGC+jywUj9kKupd17Y49DM0SfMbBI1HotXUXIzAGcVBoeLgR
zEAaFYNi783eUwOiP+2tGug18wJiNGikE36/M4wMpEtwWxiZu+xv6sAamneS
9ClNlfy5SetpEjpiz79XNcWoWAZaPGERHAJA8yJVnXGMuaPh7nPAetRWz6a2
GU4+y/E3Qq3xfpMa6h6PnuyVaqucNoir4dln88zsvACBfFt2Oks6TyknQEcE
ZjXJ4GCVpVF8kaw9O5OBDp7b6RIzPykPoXtI7e5ZXyObmtzdHce5uySWLxTE
McFQD73ZhW+l+VphB5HEERSAkTMbJG5+cDjlomGwrwR61id4d0FMWc+h9uq+
N1AENmX0qb/2OycvacGnxlei8gTOjtLmnpOoBKWLbIRoS9kz0n/L/uEx6Nlx
ZyluRLRSpPXRGFs14DEcK4D1c00xJTZc+r963ZsXzUb2XcNfoUN8RhaIsYPv
DyIxzonK1aetD2R6EZa3qovj0rs1tbnryEMx/kLFY8/nc/VHO46c90H2kaR8
M0Ehb3pestlMMI/jozkzVEbLBmrOkXvebKtXa3Es8nPAiX1esN5cE8kxmGpO
B+ooMcm6AwNfC5vVLoQThOVd8GifCK2B15xsExUieTFoRShwrY5Dwa1I+Do/
RUZjjkknV9C+S5bWik1oi/4qJ628SYyqpQ7z31nNeBGKbaGMIdd6lKFBwIq9
ItmPcwLFa9q7OUdhlJ3idOQzLYf/UfUTKfzw6aEhVMbhPGU+ri6zSPCBZ7Ir
lUczKjLDTbxcbRyvSeQfFhislyUNfeAV0N8fMDk8KlqDWZnfSmL03mVTkyUQ
MJWrlDz60NBwptDU/OvLGEr5RNmtszbivEsoDM07KK1Q0g5CmtGW5Ei+/WAQ
Roywwr7/i1U5tF5tVJV/BuONq3WOYzaY19fLzirddspGMFPSkESKHSZHGUYY
HJJvdUb5IL+rH3CgMP+4E2cAte8h+nqzcaTSlmpbklZ7BUriLBSrPmYaBZvJ
R8r1O8LR666eoCvd2mCphXIEuuHUT0+6gNIDeyAcNK54LUOXB5iw6qkO3sYk
pq8px4aISwuqWMu0VvTLPxsW5LG1oPCLZ2eLxaVPJS1FMZU96LcXuMfKJ8g9
oGgQv3JJ5csmJSgJFJg+MNiU9NIxoWhPQTguMDEikDFqTUTwW8cu2THn05xT
Ks+URWAEkmH7U16k5bn9nkEfgH1u3FP6llUJZmRcBjBcwdyQ7HzWpiQjxmji
ICHrP1QjazVYP9/evx7Y3HgVA0m0B2c2FQ3VVX3osO8W81WOgh1SqW+y+xiM
nAb0qHLTAtPKmefDpw55ZP61quZKGsoDD0ei4YJjYEgY9vXCr6mNoi4vwjq+
j1sBoqDrn3cUWh76sV1d3aYk2Uvlq43bAWPYJGheqbOE3ou1PtfthFSt/+6+
lypHHgOabWH3MY62kQPWpGXIk6cR4v4NHoQLaSi64Bo0us/pl/jGx6tJyuoo
5Y55rEmCFRnuR4u1T45B38oC4k5FiTmiYVDhPfu10FoUqjJp9xFj3vI3m8U8
IHKdzrDRcCoSEsbT6WDSwflgYgErM+QkgMuHA0hjXIAFySHkK4ibw6kLQNFJ
E6nd7rn4bC9BUNXdw2njQLxdaA0N8267WOjwCn78cPpHRRPLn8qgwU7l5z0S
Fen64H4mNSGThi2GGRwzszHrvXUJ+7xv4SZGbZKFfqetlsef7SmEtorg3Vlz
CCSnOXFzZJBJ6q6Zu4+IwtIIhG6b/IpviIbEgcQ9Wt6lMn/kOq/4wkP87Jr7
OK0l9VfUEFHh16sbY7TaT/D5nC3i5eIIZGWgSiviVc6/aG0sin+Jl1Ctl1sQ
y2BuW4YD1qfLO+AfOeRUaTtoqMydTKomSGvPShevpTAGVJZ72mlRBD+toZhz
uQlFtRmh+FXAgkMCoWBPcvxCUpnchTBQN9kZuyQYEybbdKFq9P9nf2dofppG
eEBMcGLI6wbPU0PTJgr7To2Vjc7DokLEwhMwrEKiLMl3B3hAx1E8bHzV/xVd
ZTF2ExAKJbp/6YdPWdjO23e+7ksr8a7BRDlE1x+CPujv9iLRQwCHj2sEoUBB
7gBf6u/9z5g4/MAvSMM2W/NjrDtkADzCT8amhnEVx0TMjVOTll6boI4uSbF9
EXsx800OfvgF5gdh83u9JUtk5sCvMl0zgsOBdPjxG1xWo0OAE9Cg6el3l68c
fbbZjevWJB/xd9TM5dy/Z426LOASalAbhb1KV6Hu6InhtifGIoYLqFT2VHDV
P2ovGfP9Vsirl0Axdv8/Pn/ncip8gPh18IKIKpZDQ3JN6m6tnFf9Hz4AdkQK
QPrdoWoPfQX4vcWU96QrBPIOu5b54zOdSHxRYp+1wKedorbW8vxilWYBg5qE
5cZ3Qpthw8xXw44YZ61YWjmtFmakKaHwBT2bladOCA+qP2qXC1cu8Dfi2hwA
ENUOatWGeJuIgdKQiSC9Y9d4ffAnHQOTdTBLsqjHAkUTi3smxSbnHbtjigjl
mVMmcnaecEKpMHPzsQAdQ1t2O+sqe/h0v7y/qkunhv4Fha7DpGg/W+CDH+qi
f4wU+idAyNN84cuDou/bhWGUATi9S8AH2QnQKl2R7bQurSfH4tkhP0M44FE0
6o+trv0oGFDuJpibQezpUQ2mMnHQFbs5F0Xbul8sLCXR9chh52GfE4o0rTlr
3g6HWAd38n73ND+oyBluVhGBpE5QzR1kk3PgIbZGomcRMiMb5c7+snbKUAdc
lJEzpo+KD/jiCtdlS5V/6aryNV36ZMiLemw5f6k6NzQrJ/OUPATIvd4Vt8yT
dN4otygzcfVNxxOAM3S6tER8vz6nM8NQuxn4uetEfIkM7l1lQTbfCk17SM/H
0oRp67+iLZ4R3nbii+mDmB6gIcy33jbG+ieiIZIe9j5Gt+AVgrwuBL/QgB17
jv0TvLIK91bXm7ksRrNex/mLJSFaPiUHUXjw+LFmuT+ObZ78e3hBnwt6pFWG
y2zH25EGmhMZdMA7VTgZK4blrYgQVtLSJh5z8PO1diH1CCuUsYTmr08agQCa
Yvz0agP/XxjpP65jATWuzjPn5mKUyEaGEjMyz+jvd7YX2EtQAPvtXGg2GCw7
lJigfzu+dCO8ZY1xolebHqKizsttktR62aa0VoOwfUKxbnHeayApSHHSx3AA
o2wa/U+XsJ1SXH5ZPky1eqZ5pj7uL8arSjHPnK+RcGUwFnYRrwTYSMcvXED/
odEQNaqxG70nuVs39p9Wy9agcr0+Wz476gFw2o2WF+CkE2IKqyRd2HRAM88j
G629+gdDpVfvz+HXMTnA6SSdBZrea53jkDUuOiWbpbFoH0u0RmHXqjb3WMc0
aqvlEf5TgyMBKJgozsjAv/iEjcR5YHWs7iF57+yEKguybUyWd9r1XvW0BSQ0
YbvWXmUnONl8+XT19hyYt/1t4wdq+RYa+AI0ZRnT8mjtX/bi2tubfbqZmdpi
JkVOUVPeCSlxwtGsf+/DUVuiOvHq/FyNAsIboR81F36cxhANAidTXRLnmjKx
bxB2sMRgBlYgpMzMv4RW/2y7k9fe67QhGEopxWxyckvAbDW0xzxN/iKsF/tU
tM3qP6QPJ+1wKKXHLSU/nDG/Fl4iHyXJ4CW4gIleCOJAkNJIJEr7gDHZtBM1
NGuPUePjkIRtrzWjjpF4RsBAAbej4kJ2vgQARkp5znt49BiQhYk1k6y4Sm6z
BTlpa3e3YPoFJbiXfjrGA6o1BhyyR7vdqJYHtd6lUl6tjkGAfmQC5PHm2kV4
8FfcICySG3XBH8bpG0lOhzl/0a2lWF7Koe0Vk4iEe9FTSqBxKR0SvOE2Q4AY
tQfX6uyxX5/nRwrI+4oJBKFIl0i3KktP0oNZwCWOC/ktdG/ESU+RxS2zeKcn
TrxJu1J23wUVSKhoVEzRizQO3OGy9+FL0AHe2aOLXw0CQidzXUy7Tbbv0QLO
2vr0c3N4OmGB67uZGdFv+yXTWFILvzTGGRW5nKmKv4++siome5aZRa3PTfEG
dEJmQVkn/BjHxc3K6qnaSxBbWbUpashEbGPijKKda0H+QpnZFPmq0DXi60RU
H7IhZ+VChEkWZH17oZHhBl3sIJ2QKrwpaetPAYfd8NrJal4pv4FDSRvTm0y0
gtXuZW5U1AW0o74G68rw2xWIoIm1iuycD4MU8bgRXjfDkQBONGVBQk8RZVbA
RZtydKba5B/qGdZnKaoozSmk0UapHR9hp5xImTygkIhKg3mFtiAJQNAFIDo3
lH1/I2l7y39N15u4VVxxAjV4h+DOeywiA0qHNGXS7a3kbJcifevdnXlj/JwK
GuqefKrBx7OlaHZSZq3kcPY9sGvFvTZD3XRGuixFfzzx3IPUTHZ+MltNvfsa
o3lOM6XuDY0otrEv8Jwk6LjkZeyRh3PfR+JV/J6gU9mr/1LOtmj8a089L8y6
h1OkfNgXushTHzQQ6r5T02qqYgSOO+8J9ciZ7VAXDG/9eS64neMVCXB8SKrZ
fsn7YGD6ChJLv6JJObYhvUqnXCuNwgxvA3HQCNut1RkgdxmKT3VhNhBSS3wp
6JutOos8uKSpSGOamREZlES5Eho9pBEfN1d3YLFxEzlFvL3LZgLP/lls3Q5/
Unxr7kGmhkV1w3FsLFgV00KX0rZAPYILnsyxSU/GkXwTp5KuutJoW4gP0SGz
qtTMSHUeF3eAPPrkdSh1EeKlpZsbuXVBhNmqh5sefFWJaeI9RZp9hDj85oq8
OdwSzcFx3rJDkS5WwFblo5HU8QTeo+YP7Uo6HjY6+yTvyM9g67aYkJCHu4oI
M2LYX3hm1iaYnLnklCdJLC4H9zRHXW3PtiZ52fcfLzDar5OSjajI/YxNWkEv
yqQN7lkcUSKYJXjVq8joOcbsiZIvX1yOoKWlzCutq9dfBfe+oiP9UywSjAvn
kYcEUiwfCHph574KulvJB/u//LXaaF6mNMmthZNa2+3D4fGFy7w3iv1U1KQ+
ItH+UmnENUdJWNcbHxFM/w+ph7IxVtZlDXcZQRJPjO2B6He6dAwKUbVU30DF
p7QBFjvTZJJ8px4d4wL9CB8Zl2UvNQCgqpwephcfnu6EO0FvbzgnVcz+pzG6
1XNk5o1a1+4ld+Za3/2VbX+xDM27U3CPZz1xXBI19Vp8jruqHpl05CNJReEH
zWt1N3OZLTAWUpL2MomAL0XCZi5RrK5zOJiqUqPh1XFSliIsroOcBDLGKSHO
9WTpPVxXpkzzrNpmn3jX8z2oBxsMlRTyEpONQyRfzwUQNp0x23Vdgqlhsv3X
gcZkLbFlAb/BGwPvMrjwQktLjy9+n3XPKTevIrYYDN7aCLzAKuzoTf1sZFrJ
/Ff3K6jnEFIfI8hDlZvqoEehlybdPtOR2MHUc1MUpx60LFhEtQ96Vj2fyDf7
txVE33FfIx8l5D/VwnBX4Xd72BJtWNCBRiM8NjuH9wNSYsRCDjQjhm+xzyWV
GuEIXekgYBztiFub8yNfwQZg9jN7Xe0f6b9G15N43bFeiXiImdHviEzTs1Su
tZMkwqo+mhG2ha2fFOIvAjrozJXwU+3UNm/HFFy/ex9OyplPbLwC1oWaxAex
jpzmVG/ghWVP7rNdrUl3/3u2Y1J6KkfDxuWQG+WL/agk+wz8vnOByOJJ464o
HwmjkrXwjszX4LatRCy3Pus0Bm0HsysF3kZrSyEAVxb0PE29udBzpKTTvSNr
6P3XWJwaFz/UQXvR50MHJSvsiZvULOaD3UtwIvURixb17okj54gxMYICW+aO
0qiLI0ZUZYb/lyHgHd8dyAB7/Uxlqo7A9Ux6CY+wl48H9o7ZHdFhkqo2wUTO
R9FGi3cazBOiG0/S8XrHnCFd6tWh2pFZFWzI7bDkQ3cTZqRzgcg4gLERoQtw
dm4juewCMcmqu+UZxmU/a7hwp7FUyrEy+Wlz1y5X0DArXZrudycsflHsB41L
3J/483ms2H1fv2CLt4zU/MdNIO/70MAT8IZBUq7J/9ERjCvwfqxq0x2Uz6jf
guSMPz4weQzuHGKuDXVHwgonNsM0M9wRNEFwIa8z/lMIcZ4XtiiRr8EmWfFe
kCBxFZDxtba9trZRixG78EPPjEodjw4OR89a6YnqKjMH+7kClmr9eEuUmeG7
TpZq5CXqecy1tnZotauY/XFzwPHDQw24iO2ja8a5nIahLc2V0KFxdwzgiamy
TvR2X80RV0NXvuaCaavDZqBoJ8L5Jqz3p/0Zg798x0aFIKfEC1kv4xNtkDlr
Na5gNcGZWYhew4TdLNkogmlbRt1qH1g3slB1bP1dZvb8v/Oa/HlpMVGVcZKm
LCoxTg+mcndFXNAtZXoodlN9V76kAyVPxTWS+30b/TIZ8qnkIhUW5/SSL7TZ
DyBRffYgtMsqLOskueiAm0KZc7sJMcAxwTF+nDwNhiXScF/rT7060Xs8xz12
WqZV1Y873+Vh3OmxopNIhJ19wrF+vHOLjsVAjdwocsToFWcLK4yygC1SC/Qn
P1lsi0k85s5qrwTMTRjzmo4PXQ3MIDfrB1q7aMEhyQIOD/8ELRhhhLR4Sy5T
Iur9q5acM5bsJZGi4oQVU5gX7WnsIqavotFyTafaYh/PwI2PdObkxblfuq5Q
j61vgjSzuUsnoMjT41dsef2jWfVnal4rH3Qn8XRMw278grBVTg0rPZx3B9zs
W9iHIX3BhHWDrdCOsePpfRG6j1kJ0jhxCdcj8+S67/jLzURgBzW5p5E8Fs80
IDeRxUj0ocHdWcZBQ6MTLQm88hvgufLdD+2vF8bX8b/L00Ncn19qhSIaMjz5
Og3zcNUjKVHnfZY7BPVR7cxbDtbfYqoAL7CM7c7cZIczX1ee0RdhIzbYtlLr
RMOjn4HswpcArDLhYj4ym6FAuuXzD19T2je2PXX9GEv/6OIJ2a6FbspBPn61
X1Z8axWKaTcNuPPn2boesFX0jgtNXAhJ5pLkVzE21D3jV+dyuzGy7KIUhe8O
xLgyFiCb0JOAg+wr8pIBkA0rC2yn0KDuaFhoH3VPC1INJVMHEkbX548BYVJi
MVMywAFLjVODYqvCeyyLXIVzb4h6minAWo7/ScrtSFAykynmA8VnOgP+DgyX
VHdwk7b42X/MWAxAZpX2i2IUKgHT/Umwauu5C17itHOldAzRtQpo57fpga7p
mC73MaHUyYjNqwG0XBk8iJsGEVFUiIUOonYmCAVAcopOawFAmnR2GY6oyEdH
bXdHJcoueAT+jd+3BUMo7N+LfWUDjgg66bJQ226YXUNKTC6fhvqRDXjFSgx+
cjvC8vePnEXsW0YfxMvC7lQfEFmlEyOHFGesgXgFaEvXyAOOhfTQIkdk2kZ8
aqBndNWQTyzKwc4pdKRNa+DaahEd8HeViysKzmnuOMaPjlchYsdT+gy6UBWd
+mpr1g2zEBIXegTrj765EZ7fu/rH1yN/eb53hQEFlLM+LFeaEQCdpJc5RSdk
H47e0UQQtqcoIYgJJoOdqFbS9UUI3GANDqIixKAai1fq/t2nQIveG9m78nIC
gUqXRtdGUBy1VL8929ZXh7Hvolq+R369RsXdZS/oXHb+rG2UAd6Sfiz35RfF
Yu1vFlbQgl62hE08xRCYfSaRsQ1CNDCME8kOhJEE2DWuUkrI29SZFW32CVVM
WbViRIjBJ0LvTyjVNKpzjcKTB9hY/WmfBhCQ9ru4clpNxZWwycblIkktsXOJ
qUDZ2/p4Wm1BPEQyQgIQnEIEsF0MKqaM+AdmOTno2sOuEGfquVNWxUS5Gl87
vexnxLUIAfR4b6sHtGrg4AU+nTqwIL7OqLxMV6b96JvtTQQ+eTPw8FChpJKE
CGEw3W2QBhKHWOEPUUJzQy8KDTwQOLx7XHy6dzdMl2fYcIf7OTD80tJKihO3
QGEkuOarV5b9VhXw+p41c/C1ZrZJHaHKUFT+mSxt/0axCtcpgKdaftLVppUv
K1B14q3EpB6+8XbCZ3yE1ZxNEblsuqFTnMWirC7i15V600b6WZQ/uRq8wgVq
8r4LmvHqv24BA+f31AySoDhk00JiTVpAOKIyJ51R7GnxBD+EkDjeHqX9LC1/
//bufOeHleYGX8EDj4gWYyFf1Rn/ggVANwmw7aaEAzZd/EP9v8Nh9pBJw8qm
R1SGLzPkSPqUqmDP331Jp5ktJl5GbL0Hl+9vdehW3LCySB4lLIVEvWLIbIcV
WJtpWQRm+Lt+9Tfg3Di4cUfrXrTsdNPwIv+APCCFnev5JXlldbAdns+kMRtF
T6aqq327V8UghnwG/CocAl9msYYR61ob/XG/olyZNjfKyiLxw6ZCoV/Cft8f
DMHNFUiM4XsDDaTGkK7jn6NA6SxZtv112pxp76hbeU8FgaHiQ/R6u7socFWS
Ew9l2KXbGAbNQgoD089Y5rP9baMt4t+bbgEkjHIgvSVL7+rXzG4Fp3PbFh79
b0TsY0ptWQnR3ADcGxffhcC5PZYXBX/6x2+N5Ukt6d8BqeVVODBW1/TmRchK
RQ9DOCAaq27ls9VXgWXs9W17ODMyk7uaI7weC6TZ+0NHdI1ksnnMMBoNDCce
XeoGdbCbotUFbxJX7pbWbdwDJeHk2ksT7dyDWwhZZyvr9iS1IIYvLd+miUtA
jJJ+bh1pFPCelxOroSmkbqyf/1YSZqHQ0BCjpL3VejmXm95W3YzMUL2BbOzf
d4rKJRpTsmFdM6al493JhUZlcjAEq+b2KSPfttjTKDPXPTezLVLmPLD4zDTo
ufXg+GngWh19hrGriLlJJ76IYOu8aYvdui/fL0r3epQje25Xz0FY7kydFj/g
w8hIwAdPkR0oXh3LkWSt+xmSqCs32y8UR90V/Tq5NkkbMAqVnrDRCR+iJHsx
UbL0O2U9084cemkx3tFjA2cEPo8WirXAH0iuPB5jVK/HAi+DoJsp1zFTPIpx
vEgo7z08zrxe3/O/AY93uTjCodauFH2f67gkOEWRVK6BICI2GNyyD9BexFt9
duOLywoHhejHfGrEsl+aaz2xHA8TY6XbdH+J8ToteKTLgjtNNaRL5VYhunUY
9TyBcJdMOGwxcsKXg5qgwbeZIg2UHLhsiyyPTMGRLOzvEL36kawggCeSYKBA
sG+IiQ2OCzy6HLGm8uViWoiKx1PDtNxjMWEAc6Un6nBsRo73j/wvXHaK3aNo
wffP1WEGGJK1YoNk8n3Z2lxmRPjm0OJVZ8k23XJDn3+kMEuPI7yHQ1G1j8HF
9vokpKF79WeJHokV8hkxJnd/r3kkscSBl7qOT/yp9eWDc4zMuPmcw0BKnEj2
RdAmpkDFc40d/1glQfvRJKZ7OgL7kYuU5ipeIuCYEkjPMsbeEWPhgcF1RPG0
ACEisD4dQXCV+pLWCJ5kgvfJY0Vdq0NZ8dx1Kzoa99pEeKTe1OguCilom5wI
S/a7tsRgTM/U6tmj2bX2uMeMRgyHPPB/UVi33HVnrNMDQiL+9Wip5dlNsA6W
rIO3ilLfe5NkHvLu4Y9pksa77Z4YRbtaL55+78g6KZiFuCNxls27WsXC0vMT
Bzpe/INbtq9/yVKfpKEPLIvAd+pREqZn6iRtup426+t2bXuAvI3yP+86R6L8
xMI3NT5elfgrnIR5vpig/iew1QNcmLpGHtiyaIuWX6miLfoXS2+EM754cGi0
TFq//L14ez26Bpo3tYAskUaTna5+t09MLw8RbXZThSQW+0oBRrYS4OjmmKSn
C8hCpTGja//EvLn2vJT44dTqb0Ikbl1oOJ+K5qjffLRU0veVcOlBcI2khaHa
cm/epFri12mplsQwZyHoIKPXODhchb+lVz2g29EPmCojqKvI7qMVS9alIYIX
d171k64EdBUBTtKjRMvmcDRMgqSy6GDzGwmMvLzvGFLdD7CHVQ00kZ8hvrfr
ieAvLn43+0J05h8kNENhzP60lUPEfFrnvTG4yyti25lD8Cik2BozA/f6MvRN
P51rEs7lKuv7Tb667hw5ke3dSD1Ju9ibZVfdzq4Wk2YEgaiJOaEr3lM11VGQ
XAVGwm4Zfk1OnU5JznkEp9GU/neP00X6oNWCbANc41+yvtrKSt/YL/PrATE1
FMrmpEK20H8nkAkr27xAi2D+GEBegHqxkwd457z3e8cvtEL450apAaY+g91E
rfVSle2HnESszjQt2mwNKOVgHQkAxpCG4u/xynrHSRPZyMqFohry5IxZxr1P
uuzPJaRux1rdrkg0eyIOaAshSMDc2TOtu0/EmzBVc6f9arrysH84ILkpC/l1
wTKHVtfNOMHdR4AERh+gc+8/J/pPr47Ht1+c1GluRYjEVEqdmdSkdFdXbcLH
cHb0rgXBgf8TzewrgiXTV+MbVByYjpZNJGgb9GdGFK67ILrLtuqA6ycFx47G
qSJwaXrPbEWNyvsoP/M8YGe7LgCkETMJLPc0HdsdfSg3awsowaWGRvIQIflE
huVKInrqkoQo9ina/hNg5lYynwAYCfw5wuVj5mIIH7jMi7e3loNkWuBSTeRe
1r3e1KBwjhl4mbivR1ObxC+1TqYvfvMjN8WGt0m0HOY3wj1rRy7BLq4N7FZM
TqiKZwMCO4ZSaNsk5USrt0nFVj+p025ufkIQZMOQAXtv2VjkF7C451SeT6wG
+V3bNcGHMLloYL1Fj664ytrm6D8Aa09KuSFpmFlxOJH3rvu0Eu9dBKYcqhXU
rF/MNAFHskQAja47nAEqVhXun+zhDPo9Fs9FFvFFv3tFkD7jnAtJ5YB3stKz
udhYDVduJ1jxoeWDlwieqvv2e/WGQPf4jyhJ2qZbi1bvRWLauIUYJRD8HTnR
tS6u16wYKUl+l/CiGiDaQ7eJpiHZakxdJSs+Cq4kVjrbW+Zuumf9tJ2Gnx81
jneNN7M9cviS7Y8HqJiMI6xaMn/fekqR2Uj1Rb6BxWtapSX/XGYxZbSl5kqZ
rQdJTZ6yQCbllVGiEYvydn6XjVoaJcc0q6fXaMhz4DesAJFuBZU881f8fGR/
chbb25irhV5YxSeqgFooa4QafGNKlE7x8MTo7jYegleUokWTRsYn8f2PYPUc
mcM0ohzxSjNVGoTVMe8p5zHA3lmWik1No0eSPVRghzt71plRt+23YiP5SiZ1
62qEOQW+iyQzFn44b6beIqjnKyzes4cO3ECivcqV8PF8wtA8o4mWSBrlqnwL
hmCLbwNw5jyIJeVRUQCTnn1ctSbT3NfWBKLDuyrADNjvrxVLVnU6Sh3lI95+
VvgQeDoazueR9p/VaqR95fKUKuOa+eKTEp2/D2qQog3nTz0K449wfTP/Atnt
3N2b4MBrpa70MNhmjf93d34y9+0wETuCITIvPdWZ64iGRnSINNF3Tj5Q34PX
0/6xXHRLFrYkLWiA+Got47LmjIZtmTVeAcXijlmzwqz1T8rIYYlXkrhNgAK9
ZSmA2vtG+4AZzqGgvUT3svpNhn+FDSu81UY3KSMk+gzVKfoDbbZZwDewJuN5
ZhIiPDWQEmlxLZJNGpLhHYOkDrCCjM7tq96gHrZe8oY2u/onx7hie0bFJ0d7
FyDGp50rTCDiWj7rlS0YVUd0Y8HAJgC4g1+PEKz22Ban8ZTUdJ67zPmeARa6
g7jFvtj7Ml9oipNcsJIiWHmvuPD2kY2Bpk9ZWVFBU9rDUPYvy12aiycBv0a4
w2pzun5DhrQSHqtSuImKiL9CnD2kOsGhRKI/GN03mnesjeC+uMJNaw2ycvLM
p/0Jp3DQ074tjoyFPgqffRVksUZStgmYL+VoSWySqyhM+XSnyryA68o0PERl
Ezp0QOxuoIOQdapjUXaAOmD9EC2qoXQ9IrmspnKWUfgotO5WhHYiczvOSPeq
IK7qfgJTMqFWNIHr8kEUTJ+aXpIreMs0CSGSnWp8MHq2tTGXZTSF6ry2YspM
eK2l9VZxMSBaoW7Gr2RIUfLOTpt2wQdnW86xqu0u/5eGgrSlGibjAP+K8q9g
wZgQ2m6OzIZQodTY4u+dY+U9FIIZ8xwNPO+CT9OkDOboCVDMWL5afcek0AJY
ciiIQR25QSwep6e5Gwt/0lRKy9LM7ha5ybpKqkDSyO/Oz3cJfweBwUwt3vTD
yuDaPTdZyGNjSUBvFEldddb0YXmu+61iNA8rQKOmj//ZegXZ/0S28zYoBqXh
rXICvaZQsMCvOhKjXgJUFu6fnOYXT5oZmWAsXLLv9xEOSxloO6A7ur+KR9xf
TyLFz52GFUpJis1AUDMJy+1aWY2KGpuM+/djZEMLDPC1am/GftXo/QQdQqCe
30hL+YxV/Hw/Mi9f8mrwToF1sExuf5mNOVnM869GcbTEVI3XfSN/bRmFnr6T
NHc2dTbs//OGkylTrrbAs4b7McEcorW2wJuvN1Trha8G0aIouDnhHYccbEhi
oQFfmBRjOXrtawa792aiNxsxo1hfAEKh7iBsXZJLzuu+J9KCUmkXLz+0ZO/4
RQ6OeAV6Chwt15PN2PMOAWufaOhCY4FU0GxPd1uiW47+/hIOx5+yiN/EBge3
kY5OoT4BedNHyzjCmvsJTW+5Mm1Bbjbrf0qgU7PiQj4PNuVhRY+aYOLRbIuI
C9hw+mU0+5yMQOAO5EVNit+cg/vII6JGxIE9uib78Et/n1lETa4PhG0rUhA/
cKNuz4CLVLJZvL8/cf3NoDrfJ/I5/ZG/fyN8wzYocdKYA0+ql5Rn0cTuqodi
7dsRxkQYWUueCmVf+FyzhWRSkBJKghMyi7JtmeTV7MBad2JlNIk8ad4fWFVS
ho0xMKJbznKGW593+MhPa9IhR0PKoCleIAx4kn6D3wEF8NwlQ9sTqRTNAEJV
3x6M87Of7aUaVCH9zNDSdJOcPBMgqgsZQOZH8kYihACkoayoi1GWMqNWp6Ac
wUkPyDbJ2M2eQILjUSLrbkYkMe9UXoVvJhwiBL35Xz3z7dTckUReJlZbG/fc
8Wtxq6tC9LW57tpIJdMQl2A4mtJ5gnRx1kHnyvGKtyRJl8h2yAniCaocrAxM
1ADt2rgaJkMXuMyEDcIuFZpMCjqKWdbQuknFBAm7krIl8jywMsetDTXyxJjG
D0/Qo2ZCEkJmo7EtFnYqxv0wbeb8LISwhH/XsPmYDowBC3NbwGcWcEUwL2IM
qWNoJOPdDDZQunyGXKPi+vJpHTmiNKAHDdvZGuuj+f5KYzpzhQoyvbzBKl6c
6kSlDVZ6a0+hLYQdCZ+Kgr7bjcXcKymJVv4tH/+t0LJk6XiPD97WUDZB/PrS
56nzcYd9v2xcWSs6iaRG6DKyDQF8aof92cFk9S4c3xDf+AAkTGkCM3XZZuKa
W+D7240u+YBUPTkJvQ/DvC+Krso7iUxlEI3ILXiBZ57lHN3HRy4gAAZHYyPh
VfZ4aj0lztZNpWYXpw0a+1y30L7FeP2BVGtdMqGXtrWpvVu9F5aN3JoVOcZ/
OSDK00V4wlCUuvjJz8/4NPAmrVhhJp+/1wuWouAsFHY+lU7XURrWIk4+saC8
xYHRkWN7IHFtOfCkmG/fqBI8oXn+ZL7+ixpLwbkA6cgPCA3Rt1+ByD8S27bX
UC0IvQ6X93Iuee7ZIekAVBNfp6tXlOkS59O2dCNPxIfFtWeqzElXl76zZipn
eEYnAOhu+yqzwn+RNAzFQ831sr3QX/szmG5hdU1ySgQMFa3k42yv7fQMVemx
MhZqz4FOAx0BIASGhaXBFgWEEnxqZhW44EUr5IcrCPgauprC18fwvQ3ulH1b
PgrIPlmjDOeHOdRuPQ2/lgVyRp0HZPyet68IohA98QGQYudZLYA4APWPzpXI
ITn/sTKFVSZ1Fvxl6V+x06u5I2siXfV19TUj4RLYBWHVCv+MHiN2aJV8X7gR
gBdPL5AAR2hDjbrQ8whal/6exNCMiDRGQ82RFhDQdxJ2HGirYRs/yWNbaQvY
6CVMk8ZqzTHQrmxL4pMaAk0v9exNPcYQ7JStlq1zaZIfEEJoOq8S6ubax70t
fMVrn3tbsNscL8FK4ca81MxwEzVcHCZgo2HL0zj/JeRuioaypNrpVFL3o0EX
HePwb6BGtDcBDtJo+X2nGKi/MHWRHlAfMuYAM5rYh8uaeZ22pgCd+/hzRFMp
ln5Z7CRnP8Q+3dPJdzLjCVOb5zE3h7fK3WVAkqqLUOxzULDtiR6buedMzaJ+
LNsQbwAnyjjLASXWbONXQ80hn5mZalklkUDEdPRfJbtKi3oS0rX4Ynkx+U/w
OnPJTqc6oekhIh051+/BK2ZzSdnJziXigrDSHmdg+GsMRdqw/w1a4c1g63Cm
aNgvOYiP6DXSiuGEBrFzUbG10zSAcMvCHgWth+NOlmvSU88oGNyIxeBTotgH
m2RK9ezuEynR3JUk+FWXPE0kYhhWGOBVU1MfOwXofACKhRdsw7W/XP4UJ3U1
KvtLbzI9PKM0LSL5KP73AXdz/VurqLv2ULbmgnLiYvicTXT8C23jVfcDl4S2
iBvb2FJUQmoFCCTRWJXIrPw/WS9yhMAI+JCKNe76v8445ppgr7HEXp2cK6/q
U/KzSMWeX+gHa1Nk4MTG13Xxp5TK3xSpRNTFH7teL1XU4+IVm8wGqjTlbTWL
KZGULP+RnNuzmoHpqXnbJNU3RIxM0iWOPFMGJYhLoIVxQ1XUBfYAH98/PCa1
iBvmKKDHq6cKlGwBFGwIy0y2nWhiSH+JstuzDY3Xwgg4kEYLk36abo+ev3L/
Ggkhta7yGMcC9nzSfXhjMT/pZnLQG7uwsMtMai67+yhBTQMuxkjrOzcG/GR+
UkYU1O4oLXdgylHG8aT8HZ4oQYKTDmkMMWrweDzG+p4KYjGMdM8s+3SRuQq4
vKeXYHQIV1X4hKM9PRfts54j+Mt20gYDw5iq1FXLZKrlZIkp13rtc+uNmeQj
7PtAQPX5Q3aBur2FizUVw3/X008qZbgcxlYr0doUWjUpHQEd2+Cva8qv1FRr
f36x+NI5vmUQw7XODGH30uszqEdZMEpt6tkJbCirVeFJrsV8yeBQY7iE68F/
QuN37uqro0iU/75W6R1/ls/dBx/qw9eqvNqfi//H4SRDfKjXUc/d6N/OR7md
96/7XlbsLf+lCbv6YIlTZSyyFb58XEGlQpslM4QaaIL+gqIWAD6yiIqjvXbq
Fk2wNPdyRKMRoviuuoHTSg78BC6/mKnjHgd64ki31xZJqGcm9REM5OGyBKm3
i8S6cn+B1qxkkHYTaHm1ocp0smieLVYxIE2njMn0akwq87/zgoclr0mEW2/G
1NjwMHoUOG7aY0QchSK360j2KZRfB09U6ENcwAMOyOO76SF5W+gkXJsnYsGe
5uG0OhbugQCir7Zf9iCEAkYTETEm7fiEZq81Zt0u2sMq7g0NfKIj+BtAyX+8
3RpspYqQ2AmVZyURA/FTB7wnWS3GX2Z2vzIonwNJN18hPRflu5lzGqf1RaW7
Bljr7rOAYts/t88uJ759JmuGxcW971ST1E2XVGJ8xWRXquxuuxGF3nm0NdXS
zw8rbsiu8RJ7gjbiRYA7zon5pQg5K+5nykOrkmg2sr1oksyogRfVA089Obxy
yrhgft2Z6SJmMlM+pxb+XpcmAwyIFFpZC77c4VAZaL8emdXNKXzxHVQqCdql
fUhq8X+qVYYRfQYuOjKXKYjK/XftqISPF/CvpMtQcGqVW2nJqm7SV76kojhu
qbBS1vDN8hxC5tqXgJpWEOopOZKOCVY81uMZhMD6DIA/uhYgAsmaiT5EYUuG
vsG83yjSEuzX214jbcjt7l5jL7a9YJIKGiy6Rk54dEuURA9wOuKIvFphRVgy
pE4Frx2uwk7d8+yzMn/UDEaB857UTvFMB8rqEh+odCxAF7ltErnAzdwrWBFr
gdwhGwEVw+hh6lkQwMgwsMPfAKPsmyX0gkHxMm5o/8ewDwZWIHaISgxUyfEL
Cb3Tk+LjIJyYSeS8qyau8q4vwOKuk/gYK0F5OK61NELM9KEayQf/xlAtCy9H
Q2nCb1XiTz6Ny/XTHNRItFadZC3dXghWzonNcVERLYrWS37GWW2Gtz8g6U9z
SvyE4nfJE0UWn2eUj4RCPMa8yEDA+XMkpCO2ekC6KcIZU00EepxJCZzYsdqv
CFuFG6we7uMqzeHzk9+daIo1i9sOw/zn01dUDQbZWIPf0QUkumdgbEsj+Luc
bvUd6N5rhempKTJBv/MriodIKlcbms43SYcoVUjeQ55ynR7b/hGIc0ALY6/o
BIN1pL5IbyZixoZ2E7x2nwgONHij2/BF8aGh7kb+gkI/kT2ShHd3AbbwpIvZ
82vC9wdNZnEqrvwRYA7tDGxUFa0k/g/30vlcLYw52dSgkoXZJa3frDEvwpaH
75J/QgAy/2sNXHZIHUIUq6dALsqDJWSjd0LHGN41cGZfRtVw6zUSNodjBmE4
CvZJ7vgmEbGv5Fl3Xb12EZ98cpb5bGsnyMFPpsB6qHZ+MDfG/4B3eIaIVE6i
v3BaHGYjZTYX3/Vz00C2Bpwhtodfbi+Yv204BU3SKP0noWUtvAIMkX43eNkD
5ZngvUx39+J5+Bh4qM7ccFT+dOFWVF9O4PmWe/pi1xwc02rszQ2YGOmzuTtk
vz/hcClIAcvm76KJC+ic5W4UO/dJBbRElQFX3vW+/uH10De0WUaCuMN/hDyz
dbws7+B5B3T+4zp24JXWgUspj0NZ+ddCqJsOVlMmsFHBVlGBM6WqvzG2l0Cf
uVkps8oUUGeRH2AEuqv+KqaJSv3sE7mmf4JC5yBXkKMS6TitNMj5MbPdacsO
ysv7rS04i2mGoghzKGtikydPFYcXVnodzootYzWqF79I9E4Flh2dtXNeAV3N
ZRQy7/ajPdjAX5PZ36kyO5ZHCzRNr84Y/+XDLVb4+e8PApyoxyosQbjrhnxL
fZGYu+/269t00Xan9Mjin3nseagJM9Y5YKYktKh4nbpn6EGIWahUVhdEBJgn
ju4sNH62otZ6ym5ZB4OIGlOq2KNUeXBPZ/yHa6HXwWqeVJLvsacf0l8wpqhJ
ikeuHhgb7/IlwnPmZZZLXwOIHJZJ+aj+uvH7C56afygU68Iid1uUJJPts3H1
ugpn2rkFHob84Q7CuI5Xnt5Oh32BQHzCdD15GMJ2Ht8r9sc1gopbNK6XkK9u
8oaFpSC8IXV6k9PMSUHyo68sjS9FWzKiLCo2BfPwUU2va97VzSNrjiYUZLZ2
rSqEH4+5Fcybzdcp3hyp7BquxsOxepnk+LahvwKgCBHo6V5YSoydhV9rIhdR
/IkZ5DM95rxgUlBt8Ux7is1A8h3iEhlV5QV8GpXZdo2bMPxs8eGtHD7LdL58
uH9j2ES4OkQxrkwWnqYHIXSlxr1N3wKd9BAE+Xp5nUM8IUJoj2x9DW/91mBy
vO/2MQyH8NtUgUTPJyWAIVXhFThIHOrWXqJohtDNLFtOXdXy2qZYvtl7/zxL
v11Un+ZI+wwnppXFLkWOC2FeI9+/CFU44AIr11aKznUroGliiYWDBOicNGKe
v4kQALmHjpzfA4PIQJqR2PvSQzrIRWiKad9hifgU5THsxG4CBVymsMx10WWm
vQADPXpPMzkPrt9Dia4Ztg4d1A7SNYh8Q39NhIpjEZAmSjXU82RvKUJK7npY
hkA1jAZ0FS/LCS7rDwvejhr2CvGXWtrf5yW0oEyT/I5hCmPco28HvZYusxpJ
Unai1Z3yrV+oWCEaK+jkrzWZIvLi/kp3O1oG2XzVPlbeBeOG5oeuHedfEi2o
xstokpin2djRV8YE8Nd3Nqx9NkQKhNEiDdU+hibjQi5wGY2lqu9KPpBo1ur1
lxK2yzVfGfaZ0tkNWz1BY9imCaw0HxJ/XxNx3DOpIeScJp7kbx/19ncRgVMn
4rBCSMTAuCICElXDNXLJalCUnIlPe5YoAqm/OaA3+NsP3KHv8T8zmgLXNt5v
keKoL67CnlhXLu7oToXnfCQz0UZmEfo1Rzg98bU9BfWEYncZrQH6zY9JNu9Y
Jfgi20IJinjpTeVxHFP/jQOvsKLuQZECtrol+/vhID8a4KgvS9YnsquMHzB2
SquIC5tIlNV8uoISCGqrsyZWp2HAAHV86Cr+6uodf7Ax8wv/XhY3L07PMMYU
zBcxLKnfmJyigIrIyhh7kMRSSIgB6NGIyzvxWpaEkap7IqII8ZkdNiLUbWP/
TqOOpdknfLwg5eCU77A5gTok1UTqx4nPc9L8KBS0IkIDa92tvEOlDQ9bfHsM
NE+BMQBgm9/n9hNE46eyt7IYTHWI0F+i7J3RPRME0wElLMTqQ/syhkmY67TC
+1uApBNbM4O6oSdBuxSFb+eG2SV/5mSJJoKdbGSAdVpRFk1TigA95UJbyThs
F3wfTdyT2sZEw0Uv7HMnd0sJfefRlpnlybOsP3G9nuiM154sYoaSf1qk4/RK
ugs5KBxa/iy7oe5Vx9/+u7QEuWi7l0ebezKSB8xUei+sH1PWhJrEbVEaMWNx
skTZoIayrOYKkctlf9fV8gq+aLHJ0foQrV/IQy15qBprNuUwQNK5Wq7IVNqp
v2y/URh1lGLqZWOf1vcybYCwxMzKOyN2K8fRB7E75+G9svTtK7mclDankgPS
4FAJ/EPClx/jNFqDD9d91l+Pi/K6adP4A9PMI9Io+h9yys/gUC4qUqN2F59H
ZX9Ezwcr95nT1VUuBHarz2fz1jFUyvFfGB6Pg8CHZ5Q1YiFTCu9Us+FfIGew
SYzHRAbJ6wsJZKcV9tMYoquFUcYRmKW/+G2a54QWqc52d34jmi6eK4IYQYTs
vyXTRyEBhQ3nBDwzXiqqVZal2Ri8+3ihRCdj9TaRI0JQGwvZruJ2zip8DZ9W
qI5TgsmenAUlIFgCbMpP0BMcSTHSSVVAJaX9moywYo821eoGSIsTzsJGqPv6
PVBfn03+SHDYcpwqGOjnrug6gHdoLVW06hzb2oSQovWmxKCx6FUaZaVf1u19
R8JqRt7knWGEh3KLCFz71E8OdhfF8JxEkpk7gt4DcFle9bUpSt8wJ2wm9i7r
aVIjJia8ZMb50J3wVnmWrqH9za0qvTp40G7q6754HobDlQYGPTa93lVXZuJR
XlYQSsMKZi3ceoUz4i9AsCMjZDMTeDwVSpPqy3fEOZaaL8+bE14V7ktTmQn6
rzw3okR9SRqDS8iSjbUAGeCE8o6Q6fxEAQ4t2RruxyDKeUXjC4XwUnzZcYyb
wgscTrr3rF9WVk9oUXzaQ5nedUQOl1G4CiPyL3tBiVempY9jz0eCvnEGHifU
8YVjJocCN2vTRbOyb9LBYBRV1g0moqEKb5qjJYr5SWbfO6mdbVWghoRVq5/e
m9sKPoW55Jzro0TRA/whqT/QgPv+dsUnDIHIZVTSAJX4UcX+d6PeGqFmR1m4
ihaNBthvKo7JJMXoMWvL23fIlB/AEfoF/Hz9s22c2RpUgkPbR/ybZRGWetvd
HTx16/I9WMa3KC+sicO3962nRAfDCBHQxDvwZkdoluAatbYJhkZzAvgsGnYd
RYvxnGRgzMoRg07InSGFTLIl/xRb9JONUh6UnLxpbZeGJE47wp5ElGcLkP+L
/Txp5BXZIFrTrNKYpm0D+H37drp7z3D2/yT5ujvup54peecq/q0vMZAkrKQ3
lBi+hYRri2zP1g2akgOoRwUPmNj9SdaL7rP2qowYML+Rz4bgVxBthwmMYug/
jPWbq/zb8rYLAlm+fEf/GnWNBsGqWW4o5O6KcP6/uPNJLXvUB6S2xREkF+qW
BlWlyN0CyO4KOGgm3Znsf16PEsgiizadNMRLAVFBUqIRlwRen7SFkk0Myc1G
kjrQI/RZISZ66iicQlhxKpmcTuOwYkMuoWqyTInuFgtjSJedvYrnFT53oa+u
yvcMN4bXeDK+PoJU/2k+FztrF+ut9ya8ok/VLISS1rLnKNTNj8M9QfPL24UB
VjO0vOH8wHlwoSGe6G5gsTWuomyGreAzcVj1eaFx5c2zEIIe4n8bvUOeIa96
CM1D7F+6qYoNESQBKwWOg/dR0tXZCf3+rH3TnPFtIAZvEkHg/21c0W8bxq6c
dbAv0EG1TD3UiMatsGUmxQzvv2Z7Zl1ETCQLlgMjpByquWrBrjR/UqcazkvA
t+KtLVzNfbSoSWvfOiPFz7JVROIhBxhoFKe1ALyHfmTg0QsSG3FwBBpFEfPH
bbYEEpTYMegFqLQOe6ih9w1XGl16dGrxcwpAmn7SPsHM+KIu3Rk1z/xev8pI
3FbWEK8VQU/TGvy9z13Yi6rGJ63GZ+yQf0IILlYL545WC1oqlvy6hsr/ykwr
zBR6dCgMyNptScKE6GwtGxpLqTW3GxhIq5uYVWmd1mZFX4KXbZYHiBXMQec+
12OTmOvqZc1vBa50wJgbaTMX06mbEw0Liro00SoZANydhpatdm6G73Gp6Jux
WCBUrMy6jLDmBjNO8oftVvu/qfy9nJxknBDitJzQ04fR1MoVJ3VO+GpJ3b5G
UafAryfvl1n7Pyvb852ypEbW+cjx/pexvQBfSOAxdM9LdT9ex1JPEQjiNucB
DrvgQWW7qKxqyaT9kcKYVAqqvnl6ejo0mZl3whEtsBxsywOIC+qSd2QpSOXy
Fl1zkL7xNzQ2rVzkbxRcdI8TtxZh/yhkA+l3W0oW0tV1z6tRLO3WUWCvr0TY
GkiM2fyFzwk8NsZEZUbr5gkL9Vg4CaypjhCDrDtSGxj1mkhYGMhd6L639NIk
SEO/7Oqb6/zXx6PXf/1r/zS+Xs5gsf2SSoL194eKdXNQxKaVzgBb66z23LnK
GCcsuiksYz420rYcItbAtVpoj0RSUEJyAoWqDVvpU1eUE7bq/JdRII3kExFM
hh2O3WvRm+zNxMl8LPYXF0pCcreoesJNMQxqdO4jXIy3NlcuYoUfIi9NhfFz
CoGtT1sDM5O63k9xjYOV/CLGFLhjjt0mXVlUGvdo0IYCuX9CXl53XC0YH0ng
+x5o/N9YnN0JDBgZNjaGNgfdGFuK6wva54Bm7AOyGT5JaJCl41WrBBzRETZw
ohiL5k9gZPvLCuKBf4tjxC5E0yEr44DUG73JoWFUKsEYBasTVMKE+S6P+01p
QQctV59HLHcftIJncC9h+MGOPfVzGmVX1cd2tC1d3GtoOMSCw1I1s+KDGBc+
jHpzUd9pR0WNuzyU0px5Y+vX5Z8lu7r+f18afqvPSAnn/JlXsN+WG0u0YQhK
LW8QR+0V5uBQ7xxGUi6hlONm5HgO2aRzhMbhVhtwZp1D+CHxK9GgMtCKTkMD
w7khO1w++FohhGT0dtyCEqk0MrsbbwSSsVK8UP+W0b/m+S7MDLfEv0IkJ/Xj
x+BjyZSogi2k/xz0BzKY/QsmzyUPdkX9k3KM7kiOe7t5WPGHroo1UmolxJ0C
9W2lAVRHYNxN9ducTbe0WrOxaQyzSihyHvg3W1IZ1M50QBufWNZN9EvP3X4X
jXIQKSyMePiRby1VjvmNYvk+fNbKZ98upIyThZPHCVtrArl728LtODg7c8mv
HFLtBWY44Js3ZJL9IND2aaZcZ4CQRKgT5stg92tb6ntB51K3Mc1Rbpv3EKsz
tcK1I8annO/uEpoq0bJNyjb/5P/qM15W8oqz9IZ2PFmGduawlCip0kcNGY/3
kZL8uhyWZU+p0heeFn8/T/UggvZhDUKpCYI6KI2S3WTKn/Lb4O6L/3qZs4cE
7i/hamKWZ57JdxS7xfjRIX7h3hSIc68o+zIep+mh3LrPoZAOpajnax+9ac09
8K0jPPuIRQNubih5i0oxLt2VtwyNs/Gt2ONE5nzqxPXQHSX4APx5lJvQAxEe
vZGrPbP7Yxp3muKoY9C/m+oI14ojuBNZ+cuaHlg4KBgaUFguXogkPMJZKFie
nQn4k9yRBGknezYAx81D6rCbh32RHsfhaVmU8G3BHyvGEwNVgEI25I7JuOju
KX52e/9nGQml1wad+0fbY6vCOdDZdlxUQReTKnO16LlwRbcFjM2CNUDnphWy
MA2HyxUm0GZs9DVSr9HdVtCEQjTJdCRPDyBMKU9lJQzdSonKNU1j6ecBGlFB
Y/QzAcEpk94x8XDIw/78/u6n9P//jw81dXFRkDjGgj1c8SZPBKfrtUVx30+W
6Xj4dwhTR95H4JrZ2WiVP53nzQfZnyO05D6kkV8FawhmpxD1ONGupkuu5ObY
Qq1wejP6/CIm96UReyM97t0zbvmZL2jHR/ZkujkzFSf01/zWTMh5FwUzGHiD
w7MoGg01sgEdSRGA8eBAS07N23bq9Rc4DxR9dZQ0s34ZAgkzzXh8t2EUlS1o
zT9HUZhWvCt+jYsd0NIetf7lpGInXztuHQs6bogvmzYyDe+zhhunNYjOieMk
Yhd1Cyg4523zW/Z/s9tpU5Wn7GtMETWnhiwX02XENpS7kHAIWRzwgCwr7fT+
a/jrmmsoRaJDd4MQMNNvxIlkNlCG6xZVeE2eAxFFMCBUjPoNLH/1wDi2lYQW
jlZTPpLa1GRic/R6/inUbVtD/VNQGJfHwuXqlglCYa/QOrZiKG/vl4QuPD3g
rSb4qK8qTSXmTZ42xoXPQ0rHVEzh1tY8jFWb/xUm71m/wCPQoLyy4g3tq/No
M+ocStoTHQdDDWhpSrJbDC4xjZ/p0k4z6vmjvKxg3l1UOZGYB9pfZAEZol8q
yqTJSHpvxpkA3gvc2kfIK7PkFHL19lOzzOnMO6onMUyCMb45vjSrOPigK2ke
RR6AtySc5Q1lvTonRjNdfgwAgvgEnQV9JnYzv7y8ASTb0Z6HYLOccGSyRlXW
GFpfSdLdXTapPabSeSuqZPGOJqx1ExquCVJuxTw2rQykrLr9HDAYRTYWDI/m
LbrKOhHjfjChuVEefXA9nB1loziGNi/S5sw8cyLkSNh4gG0RwqtIjgXB/CFJ
qa4LrEb3TtyxyIp438RRLgfpwWvDjZquvsPiJAZg4LuSDDWwljYtX0KuXIl3
vFV97Pq+K2jN+eBM35xUwgFVPF9HO/7ykv/pSwr6NSMdf3dfGDqKrDIWxpUJ
6Nt17MwQN9SzlahchWRjVawNgmhZ7NBAN1jnHrzj6fBtv4dfJiafo5SNCZJu
561MtEU+GYitienQm/NcK7BukK7hPPXX+iIdxAlnpzWmJ1vawV7XQtILGIQP
Vzyz1Kt8yZ3JYtf/iYPpoOqsjgXv2A8vRHzBgcATDAcbza9KgQuJGfCJnSVK
XQ1iG835BGdgvYy1+psvHK6XNQKzGGoWQqWdqsIA3dbVmLtPonT9CyGEEEmI
kjPPHZOkDTzXEtG92aAEV4aFC4lHfYGdS/1oKAUdXeE275qhentDri/HdgNf
2sKXV9H/AZNsKRrHGeyGYuAWpUZpLIRINQp8zXXSQW3M+qHNapUMfXloKiZj
ea0laKn19X9dCWX2RIjPZsMQcb21g+g2Dcn7JFOhnVvAYCcM430mqwUx+Ggk
dY9agrzaSbBtAGY5MynmG14fQvQcNG49Khve9b2VQYkOEKEU2cA7IfxUWu9o
41tIWexRAWTapIlfskmxGQsiKeIdO+VVsZtEcwS3XBo+GQ7jBCrFkIb2GSTP
PoyGaPyeTOuKDl0qLMGvAOGzeMbXpxDJeRTJicIjIkHHiZnnkuOKYG7qAz8u
dHdSnesZqCxFpzfyJtNCbRHoAyUDbQbg6oLLBqll6OuAUY4R+fIGUlySYyeq
rqzM3dN2fSQ3EapH8wj9hc13gt/Q0InxUp4/mtuhyhcIxAfMXFQX7m6xRZNS
w0n96rGhwGCwppE78VitTYU9tC+xlheZdNNHq6XZTQKBML4BKUUtH/1o9pmH
otsnlyqORIaM6NRrH4XgRA/jush89N58k/F3fduR94boA82CaeLk0hvb5VVD
5UPdZWyf3+KH/9Im/mUif8Zm7Mw7T6kawe07iHdyRjS39gOptSL+Hj/hD8SK
0DUnhKNA2Qj7Rgv5PI4XsjDA10OiaHLVIlsJbTE/pLcso6KCn3ddykMGMHLC
mlCGSUK09E4+kZtNhdp+ZOuIl+PtSpcxuO6QxaAiLcKfovoPDdUX5mKvzXYo
KTOUVzunQZzLA8I8qkor2/YA0bMHLF3cw9yoxarB81IBNkgmce6zOfAZbcx2
XkG5pvorKtCT8UzVO23Ci3ZpQBx5Bg/zLty466RY6yFq0fNO9NbvdKRYS1nB
vzK8CLKx1jtxsGofHNJgYGM8a7DYH5qBrzJJunuFCqYQohLPfdLmF2o2mIul
qyqD09EsGy3D8GmLIOr9SexHnMKZXzbE5mRLb0nu4Vk97lLzT6aP7XCk06Oq
k88X9jCScH79vL9Q9NWWx7y/sDagkXhZC7wmCXjb80HFy4IV6cFYbJGPgPlT
CQRbSGcibsUAe6dao27L+gzzgOcplmBjgxr2BtvHCmT/ldZPURF8vI1sFWLE
840ifBLl1dJ3udktuco0wfHUr0uV6UMYUycFdmWk0iah3i+7mO+E2oCryIZI
DEKDn3a3STbXgeqVDOs9tJSisqajWrkxip4deLZ84Zudq3JtH1+l6R7olbLB
gyBXpFEmsJKrXfD1oUL+noX9ahGNcaWosxpQh43/cPysTxICJB9WGFi9HdrQ
PcCtmJhFbeY3lhgmNOURxgZ0eDHoup7lxwXeFtWAggUOMYmXwPlxmSyUJDtI
h+gU0T/QmWtLyASfg3LVRAtjbnuSJfPRBabBgVqU1ngVBtRzjROJh4XCozb6
kgJkTSacKeiDeiSoIh7siwr74iz4NzkX7yFnVAKc4P2wT2nPEUgfrKkaV0LT
eaqPTWrpSc/j4WjGtgU3ET+lmBJy/Q3YqPuWg9IKrr/hvbF4CufYvkyHHqpj
u79MuBVPQCyduDO30jzgCYTfKpUvzUXcQde+Ri8EhK5seD4RG6mXDPbH9gk8
Nrt4h8apzVndoXuLTyjj1fGnYxHHzJ9r/1rK1vjtBig9eWSK1e1wuIZKzec6
zO13Ly6zY4XnTyBsQ11c+nHnIRAb4zXdwvCFCmkj2ooqTt1Reirvxu0YzZAc
tZ9KiMT9fKgaQAPx/kMDlD/HA9Cv/tl3fEohLT3AgdWdHp+01iFWoNLKhjH9
fd9KqugNcX+ASopMW5JgRhPRoJSzgTs1nBp5YDu0qupTANtzJR2Au/HBnBN/
LS1hShoW9aqHsGYbY04mI4NwCQ1NSYBBW4FvLLbA906wWLB4vkqzvnahG9Jg
a1IJWc7kd/T3YA3jtOA9iOVGccvy5CBDBfjdZsqZJ6I9/ngX8iokW+CwSqtu
abTHzWRcsigTIUlZw1AWAvI6fdIVA3ntxPZHGG+rf9lB5W1MoomEaoPzxyym
O/7XtDz/T1NIoHd+6HFXnDDkg1Z6LqjOH6IG5BwbNYwmZgW96pn5bV9ZyRWS
8aP1LxQmItzD0Umb06RfxpqUTMCv6uo4dNLzF1YRtGsZ4+VeFBf2tNPFjXdl
Egl6BWyaIfAS8CZCZcnu6mgtavp16wNDMR1SUrOt3lHYDEKXdGTRXSc02O0H
m9k4kt1qxXJzOrtZVxKdlmCCx3wwUiSxl7z3+BNEPIFBmUKdi4iBGHihFwMj
6PKjT8fFcLiCXhjqZZujkSTebdJ7YcbPI3cn7H/c6PdC2lPiG1+MP1obKWTx
kFCx6GNOfJILdyL17fdXZcT7KMepDGL+42/j8DPWfloGpTGLugxoZLpKU6/N
vKNiwFRj9IW+hN97FmIIi83Uo3mLUOqgOyBft1grNDjiVAEbnp6Y0wxWtbCv
3ESmKaUGQxS6w/vQ6qCCg025quss0jGHNaeUL1NhPit8+9NtjcGBTLKq0SPs
eFV4SiUexop8qlTzjkDvtGw+/79FPvB9AuUCI7snpidpqR1zUvkT8guQVVJu
wDQa57c7Ix0DY9258uOVrFhcpPpCy3hWeaJlSwcP7+2ovxmsejMfMLQDeLvp
mmLghoHYB3abHjvpqSSFfC8aAYTIiP7RWpzccmouYI83cEPuuwJsbw39MjaU
GTu/x8e3W11u5amu8EKcnfKiZ9WF1US+q1Nae2xEuNWEQW7q7c5y9ALlNC+Z
bpqVTCBJb8a8o4nTDjX7zbrrQ52ZHLjgQAvITCITNHn+2Dfxjjr8US6t3ixa
gTtQiAZympjEFGZ6ei/65FnP5R/f3mGKEsfpWnRL1a8qhzHon9l+VKJUOWv1
JJnCarxtBzkCDWlKxL6SgLLk8CvOmmzaSeNMb2/USiTsbiBJ0Y/v8XPz2T8q
iaNu9c3KDam51PuH6zfuMEbZ2m/xtTufofUdD1StXsr5sd6dDm18XmQ9ii/b
AKVtBBOL5cAV5nxsZgW0XkOKKRdmgQG8Hrr/twNRFlwgWrzW+AiEhjohbFmm
6a1r4Gc3LeowCW7n4UOWpzl51GO5uPPtg9eKAkyUBzAhn8Z3DNnqL8EZmsWw
gcmPTH6KI4SILlPAGM3va9bkGvvgJswT0m1k4wF5eMwGu9KzTx1n3UHiBX8R
IravCtiJYs8nKCKGzPY6aCNdDjugVVo06KWPOn0U5PkRk7VNZHZp+Qou5rpo
kJlPjwkp+TvsXC0uzPcrc4A50kZHnpQ1Y10xY7K8eKH54pRCLc5kSI6Vpa4Q
q3xEfi2CCLDkS+Q3o2u5gF3DKT/cnlHFdqwIABJBg6Ra9pEgEJhwhTEizM7t
211fxR499Yi5cOirSbPi4bhovmmswPWXAu32wGP0UoERqMQcmpt8X4nicXye
wybo+RVtvt/XjF+1QZzwmbMhvcfgCzDAzy6YKAFR3T4rwVKWH8po74ZbG+0B
QpjY/wQp/rtRk0UD/cBlLnCLMQ6+ku3cdVH5tV2cbIl3oGb5dFPCNlBTjb7x
9VIEMsvuS5CUWYn3Zq2Qh78SouyVbIUUV/R0SXX1loSH6Kg+ypvw9/DBJfYz
ZZtgsi+f1MZYUno5TSS1MFTDwMUeyPmFAG2hV8bImnpH9wGMuk7VECZDq/zK
NWEQOyyCZiQZ9ch1g0WgbAboLnWmg2WfcfTGNoD48yQHJ/tnseBIqtPL6iHZ
Ot7tJ0EiI6/e2iP3XbAH/NYFsB15NxcXEtT5BIjrtJIQdJNw3zVBJbWvxF9P
rtuyhgzjymRyCSsK/avvtZ1M99mfV8eyr4NhjupkccewUbXmM8cN8IbbcKHw
UCS+PiahnxDH3STxBj8gqEYLHn9v6hyoXVGC2y22OoKEEFzI44SGdGBSRvvQ
ucVZfx92C0+wD4SH55lq9CnO61rqCEE+xtq8GS4n9zxYgsuuO0RYVzrB3Vd3
hwamm4ruP+aARRXJP5yxlscUetJo3qijyY11lDeZNxsTS2AAF8e0VhWzuWAJ
pVZ5WIvbgFRCJ0+OjWXEn/3FzG3UXd+SUW9aPbkO4ROrbzjujBZ/tOw2SS4L
Iu7/Th/xCp5onFl4F3tTZWMI3pXe3gwbB5bFmOnWOHFmUJDpXE+dipXjpwtw
g83qXInFDhB11N5TnKCsJShjgEJ5wePBg/tGsK8wFNFR6DPo6NwT07Wm4XPe
SmmhLZZKQzOUsa5wP7V2LGfeavnT+/Xr5RqnpYM77MHug2F4IPpLZSOp9imI
vfE4g89SsQETk0Qv3DRnb0xR6CamHiAQkPxEbpYvaCZgysDuwcEhibUX0uRA
N++nqSxtx1eCoFPHiuDL7BhlT36y+hHNTjryI2w4oo+60ZCpeu4y4TFsV5HX
Mc3DQp6cS4oq6aOfgafsEIoeR2baHN4YihR6MB5AVA43yVPENTz9Spay6h6n
GxThwYSDLmTXsQXP2Jfk1SqsPgoOfVWW6wIONUH1FgdoPJsxYkHcXQKRdzPP
u0JQC2+fllwFJ2U40LUYgD6MDWpiQQCZnpnVlnMvTlh5JXghYlip45DUkINP
RTJIbZhQti+/NUI0fVHoDaComsnDCdOcWj/eFBOfxjuGyY/OWG+Z06sTydhU
3uV3t8YRnutbpYsbAdTtBdNX/w44N+XXPxWLbcigM5TFgYUe/1iS066O+bat
dE8bgtMGjBOYrL2FXDGGfapIjf4m4fXNXXX/oO/2el7tZBMkRhpVs3EjJWHw
TdYzFWJWjVgypcmM8fcjdBIBAppGjx+Mc+Jj+c58i8oWXtTyJYlLEDC/agsu
Z1NiKI/VfoG1YP+G5kPCFc5hEiCqcDMCYIQH3ouYx8QvsdjbubTBDbGikvtp
EJrlYTh+9m5HUYz/Wp9ZhRfX0h8ibIZ7grb8mOaKudHdNfo4JpagZrK3BF+X
A7kXALjQJcym2b4axLBxBTCbPR5APlQVN+uGX1JaGWUs/GTlU6qLwCibFszz
8l3e9wJLnnKFDf3TgeGMLxRnCII5BP2TjG9wtIE8fgAnxwZpMVKplErIpjwF
kll7g/r/Qg5+iLuL+9qoNFgQxeFMZcYUQMsWVIZPNUnrEfcxbmg5xGF8s/JL
ue1baVBehDh5dKQEiqBJX1Pg/xOidJOZAvirpJBrYCZ31KdRxGeZQHRdqtsx
Vdks2Efr51WeSHOmDng1C27PFw1TkLk+KtwidOorYoYso4AY+tmv/WZYTVfV
QyAG30GQWk9VCcmX8v8hxYIAc4yWZL9XSu+eMWyh8VPfQE892K3TwshUhFsT
TCJo9fVxTRQrwASO/Tq2+BD51eD/Qcw16aMZo9pYECQuopL9M/Xg8FDvczXM
P+KgyqDyXHq5A5uL258Y98n9qPDskwawFHpU7CMtaOG2YVD1ngbIkiBZtDsI
7nMDdoEs3x5CMJxz3Pz4wy/F6YzerpI+BwHGktLaZwJxxzlQtCOkqXbKW+Kb
H4/lM7Tf6FUO3e1JhX/Nrc0cC7tE39xtodh7RdcUmaPUxRlZ2LSqnsHOYPze
gdLhIyUHBb0SHrQY2wtQR92CvG/zcjLLsoYd+m5KjHufhGXlG/EIDjPfnviK
BCccVULKB9pz8fWut5ojqxLMyG/Dfz+ED+5f6H1WFIz1K5M7B1EGk6VNKdeK
WVT4reaPNfg9bSvMd9TnpMAjlDzjeN2j2sc1SgkgSiEDjb1xNyh5lPuZ6y5Z
Rpf0fzRVl1fSuL/+OVhFkgx/k7pdLsNM2U+q6FhyzrXElntLDhhq4cmkzpO5
Vm4Ovpa05TXW9KdD+xn+g2aX0vknAvbtzBi7jxbi1APYb9HKJCHxhnOBJlRq
VMWArwqHV6IhU5YkXTRfyo2cUBz31n42ryt82y0LmtS9sXHMiE+qWPoLqjqp
E2VGY82oMst/yWcTGpJ+eEkViGSNv9CfS2hxa3x5aQE0kEQsatFacNjPN1wq
K8mbb+v633eXLxTHkWzldpNjZehHF09ih8Sr1cO9hh5vtgIyHgg70+h9PjTn
/YDEbxgl5TwoMNIbYvxAzPlzISY4irtflnN4FwMXlbDigWIMOp9A58C4qOsg
ickzKx/SCGtKoXHsXyz+l7yug4uIjnP75dTPrjE3x7jyoKmyVmj3rePcT4qg
eZk1cRrDL7sx3U95iNKVIC4aP+mgU8KWLjubDY7TFZ55XyX4dEBVSS4fHBaD
Cx7y2BrW1hBMemdHx0ezzoZNsAXIIl3DoMJlpgYVB3HRwmDjF9tQAKMoNmK1
hb2+tvPM5JKKbcN0Qg5m3ED8HxN2jmsX37oFkha0bRA8inQyxugnjlFNrLWB
oAL9Fp0E++R2xJQ6dmnO0fCalql825wLbeESqRQHYuFZbpzVZbAYtXhEiIOf
lq5XuPuGyjp4a1O9ND/Fi3EYWwIW3AiafMEkdlwclXoq0+RnMuUMefWmeFZH
MlhhIbxFeQqMhDZ90hw0j+oul0MTdegtLcJrLWmLl+21iSBKnDaos1jQJ/vO
P22RwECkBFNRuQAz4LjqnZoEUfdi2/WvznUygZ18U5nQSUTavVlFEB9o41e0
jDFjIX/rXPdnQ7pbZ0wRjGp44gtE5nUFW0/HLVeFEwzsDa1qpiJ4S65MkFz2
j+ZozDNIAiMe1d1yg21cAhKm+2Diyc5iMd57/fi2drsLuD0LNxbf9q+bjkNj
cRfxs37It7Y7wwAn2ArpCPp3ymB8ClZisMmV57qoUynQuEYhyKynpkIi0Kus
2ToZy/OkjyKdJonmmTIWBCFgT9KNR+v01A1v2gqgyBFLWPa7AO5GNMbuO4i/
KnWWLtlcc01xOhBg7VtpG8N6d2X9kyUxzZUNkzICXLHD3K5ohdktL/qtkrWw
uinp5ME441EJFpeX91QZQ4Vz6vAJ51e+/0Yu8NWaq3KOmA341Ab/PeP+fAmf
bsmYfOF2H30Bg7lGdLL03Tgo7g0szQ7V0dklvJp5sCAQVCouquWWLGcI729X
MJOSWOqMugsyTZLOa7cKHRBY8d0KnNQPFWHXQfKrhKb8v49E7NzVUo9jigaC
t4+PnCBBmbTGdnYvddV07WpK4A6gnEV057DvMElmBsPEfYXj5Rw1cZReOVUW
dkTQl60PvV/UyFGHszd7qBjFY9+CVXEdx/pVirC37a8SleCAjBG0FHKM9YcR
h26l/p3IQobEEdJptWgrouR+Z6hwPYnNTR2KOfov8hI5iSUxnqJKHM5gTV/v
VPE4/uGvn9hF8RpseFXd7uIQq2U6sEL+csgYTctP2BYpNuo/Lq406P8OT6oP
ljcs8zzurDsbhjQGpUxCxGhZbKPawSio4/44HxVYE79FKKOCcgxpnoCoVPv6
lAP97A7EOe4S5fbCmAdpaqV0SISivkeHPsIYlbNO9zwJmInLu2fqdXfw626/
kt0htfXiRM+MxoA58tVugigdpdO53Yo2sHu8UEUrSKFtO6Q3kNHiIN/5M+EB
zk1lLcvAyoKVak3pRV1rkjNFSUxJOH/Qs65J4n6Uczo7GR686WC+3sR+c9PJ
Z1TFmqvuEWFMO0kCc6QaaGSgSZ/BfGUCzGSpRzymNPpOdEkQ+OJZSBe3i4V6
jCVe3VWY2svKPYdtzUbZbhXtO3KUjbbXXAAQNglUyG4hsF1s1UiLtHKrekYf
VqaPQl4AK6lI+kAGQLbwo5ti1z9omq6XN3ceD05K+QyipfPREeJmQ+Ibk4jG
OzX+kHxhA/9+JgLEO1kKHaXWKita/dsA2mHrYcFf0HWYjTLOB2T8xn5c1mdI
uQaH62yv7dbK4o/bwD13lpZpdXF51cDeAnYnz6uEy10lbsU+MGF1EM6Je6AO
55ZyOet3Qy/WmWh4L9B789H0cH4VtIRH+OnxaKra7MF0Age9oaVSDIDAVwqB
4CE/s+3TApQ4vXXF3qmuAN4sXrMOqNiizKxKEhsHWH7JjxOGlNQfyj/L5zFR
JqSYR/0Uks5RbL6SWgKXTMymWrzxRAUA32vEP4gUtTWkJZrodxsmonI+6px/
/1uHzi88qklsCAW+KE8Ijz9tWyhF6hy743ijIj79eNx05uSwSXFgkZ5TVJsi
HLnGnUJ+FVQY4BvmX9IuMwGA4yAJNXJVIUxZ8g09RQJqn3PHXVgUJrx6BN+0
RYhNQNa/oFMZsS5YxvcPwQOZPCSWRoRS+m4f1385aNa+sgtRr2RoedUhRUsT
ox/iiSOxa1tgUqC/6/aHBfEv6d6zZdBBl3/21qFzTle+zN004HDz+9Dnuxnl
+KuZ4ILUTO/3mYgAE2JpOaECSqEp5xDi8kGpGLpOwRtTfkQHcjMc3XxrD4Mb
nS1zMhL5fNjAlFKtFHqH5otRP3qSLzEQXJjP65jtMhOXv4loJFu8IFa/vzb+
QBtE9rnEOKgqtXrZmHCWMeqUtN/nBJ/z8mq80xRf9yI0ifM8146EPh9AXA0c
8fNKureXXkaAFyW3CLqpjLhAhtopSWFUQkzMokcMxdJG451mX8x3zBwWF89M
oYqcRPbEPgvvetzJEA+qlGI9fB57wN4CR6s5uj3ssxVSLo/NFGLEynft0hcP
+GZSU0vMmXe+XdeOJYnUmu9ZcdLLmlyLO27HwxGTTOhQaLNpp/ZrMlYM5HuK
4256fchSVD/Hm8W5Mp1bKCHSTkz23Ry7+5GgJGjieq9w6sdXY1S5O+TBvLE0
onPw/rWkNrzE7P09VXkBIRaazHUbmsqB8AINzG6/js3cljpfGljtPDyCxSSP
n/gjBCsQ93hZVWc5dqcHRYPWige2NkqnuFZm5iMXjD95GPZ97Rpkl75ONDJd
W5PI4g9Bd1sUNEFsIXyLsUuNb/jOrmzJWTfPOUYLEiaqzZo3U+U8SRuPT/c0
yiaac7N+RGLKtFPs7uZDxyGYiIjIYwWNZpmmZPAYMXnItTPTFQu4BG12D8na
TO5QWGy+R7GgPefN2EXH2D4dn2G3YVa8Uqg8XID7e5woc9W5HX71mT5dvf9n
+hRR/excpcGW01KYqXZTXS1GUHBpsecsTEJ8k4R0MIHt406VOpZWmrxWa8DS
dvxNLhRDeZCIERQoCmIulVzyGV8tSUI5ibDVzQ5Fwr8mbVqZsrfmFEYV4ZWS
W7lzG/VsX6frTVsp6w+ddYxlitx4KltrhlKSU2YBRiHjtrpwnQraHwtfByTY
hWg9e4KdxAEEnbZoSfyV/cyqIbPt5cCAj5F/BVGvRHwESNpRHLjjEPb0zBVF
XpbxulnZEQgtFP2lw/zbfQMA4zLMhd0kJKijqFwrt9cUO7GG40QFdDvmgaXk
K3NvsBJ/21uSZGOVawKC55QOQ6/ZDVh0JpIzc2ImxtbIxdKx++V/a1gl5fXG
POcv0Jcy1OYPbve4N0cXZRMI56WjimCZnbQY3RejoS9etmoA0H8pfVAMXOcz
1iKlh0nsgl0cnlvDgcB5Yfz+NB68EJBR15TcdhJN4k/yHBGHVt9431zcU8g8
KpIxmMbAny8O48+lNpATU2tXBKmcNo92iEn4HNXpo5fi3AAUTcvkHQh259Gh
iVRNaF1Lsh0pvmZ/FDwZIl4Zfyfl03sRXEBYjewBvXJR/mx1iQ7hMCU+EY0D
hUwoNUl3AJDqKimg4M+P0LutXHx5nGV0bTbDJJFiZCV+nQ4N3ce55RIRjRIX
MzD25ScEcQEWGCufQoUeRQ/7W/Ov/P3dzBVVB1mu/UAsaU+Mpx6sEdhr7TVs
SfjeT8gpoXWXGaT767kcv2HGPm1BU/L9DPev6WwXBa90MTJOzubOjIOR96QS
FQu9LBjrMb+NzmVjlfRHmSUPDAH5bu9Mha4n5AJntui1AwIL/TktgO79lMb6
ey8UAgSC5KCT+bxFWACibBNgQea5eKOWU+fkPULVnX7p+8JKHWc9d0ZzwhIA
GG80tLYCXBsfgqw37SJ8roaOv4SxQfF5mFBV5xDx0NnI88kTokhuQCAp5Taw
ZDlvTGxfBBq7fxfmFTA+wPe1XMYa0enrvp3EqNPAVSKkPnU2ktH1wAqrmdb4
dxMkUn1E928FFEMbNqqubow10tvQuW8D5pqLUtrF3ugQf5GQ1P8NNiu1iIBO
umoe1EJIx146MZwezW/DLvTHm9q6TpNbTJBG/InasJ97tos0P3nQooYaTeMl
A2gLxHKJx5UJaWfmIuHw4Yzyuo0dNuolBYZT3tLTIfFKVa4c6j9P5cetSZEy
8++aeNV/HvhoTdhWW6F5xLLHACueWS1evXDfP3EEL0AHTS20jqnWhUBRxgo9
VIugfMCyUQ/tffqBh8BB3eV9XYWE8klBkdy5vhj0T6bSD6H6+26nFVKPx49D
X/7NJiYEP3e9iz0m13+f06QBduAU2XXSzO76iZXLjqdKPZ6ofHKJ4gAnolFF
aGDrXENf15OdACWENsUKPl0pl5kaQ14dsltCjr5IuFXV+XMcK/+NO4JSv4T8
V6By9TxLBqdhbthqUpCRfc1TCXq30lNBwbYgjANdsAOzCZFFNUYk3EgyeRqW
SWqlvBue1dzy+v7sboGpDwj4+6k6YOPSBEi1IoqVSKg5wD0zNVfcT/61GhMb
xnDmCim37tZ181lQvwk/Q1LhsJDnc6C2Crq2giqvobO4x7S2CL6Ib1faXb7J
l9pXhPLDx2rL5g8mtGI47lMeGfHtVMJlSkDuSR+JwO4q+3Lp+LG7qF6yvTQC
cRATIqbUcZtqMm0/KlPTisaKBikkanxzP8qw6l6hKKU5LHKo3WNxbZIS8AEd
pnqT9NZw7zXnjkGN25lCxuJSc/zThLcROUaLLKREHrvtPqSUJ+YAaSJChV3o
iC1ZZRQPl0uuI8UCqZXsDyF+Aoi6bkmQbzrupJOD7nvQEqCZj1+z2tzJhXHx
kNb0LrQssN/TqIe/qbLR7cgNTgTFn3Ef4n6jEscfpztpbO26cTn7jt7XMBgN
MyuzZLd9TTnl/J3ICScZsJ/MiYV6QgbYOXBLEr8Cjx1VeERXCmJuwwbNKMmm
+efDVGEt8CTyyZqus0MkQBj4Qi4nD1u5A/hYZxEAz8dK+/VarSCjHIrvz92b
nCCRXULdrdM+9+oESqThql6/Os8JG7bJKSd9s5lXwYXm65wbfdfN4Pevr8Rg
Nm2pCoZSOSbGo3qxAvxXQRTQPJViHqxmE0Xn2yK3LBRMQ6Bzz18fzlgfObf9
iXMGXdZxkK/g9GNEIlQXAK8D2A7wEaGSShR0oH94anFrKGKpoQN3tyAXagXZ
6OXn7E9z9j+euLIJxnzxSmB5gJ0ikmITngFSOXs90+aBnUoa3tHBh2cj31wk
HLy1U0dsfyO2JcXsEHfhLE2aPYo0A3NEpEaitIigDjFXOteE+Xj2JDLCpol1
U8igmeBGNLTBCjCaRnKCpUFX3oQP5k1sxGS8iN5QysufPZNCwb9BXKDjJzp3
t8XFesoO/R3dKmb7ByLoXZ5Fpc0oOj4sOqASe5kOcxkkYtsLFxAV1JKyxaFv
JRgq+iGKbai/sEyvngwnSASDa14bM41N8TQKr9h+VE9hjK6rSHiHCZzojYmn
Q4egkdulFxbmQ6TycTVeIVn5NX+nj1oBBDcjcTfJ3BWORKniOiiqtU2utyZR
7oOl+tCa2fzz5yrpi1I6+58YD3qfCSrrMHOZf1aJ4F9dTuo+wdymSoxQQ1FS
w9FJDAcI+xKs7X1yWPXGLT3MC7LEfJ3P5q1Px7pTZMIFBF2D5xkMJYE88Cth
ag89mOD/19tdcX9xmNPWQrbipX4kQEhuJT6mCISl4TkJDd9sBNtsw/fYNoaZ
ETonDou4XGrkmZpN8dr+UBV7gdJiQxhRf9+p0khjBGiPznc3VGFIHwv1F1Ee
O4H5mVtP3fm1CTfmOdn/4ZhiEElq07PKemkHjbyuhPUz0ZcQ2r7SButsv9qq
tsQhJsDgZ10GM1ANxUULH+gYLMTLlkH+pR1QEnphDeKbpItthe4AYXJs531h
MMxUMq43BFIVbl1s4uNMugnkQq4m1lWh7hH19udMUAlVvGyFupnLkuZaU2Yf
eM3+tRPxtwOQRml8qUYDjKc4mEIrfoLvIM6GGCkcF3f2ibbibaqUc4/X3RAv
AmN/VNimuUIT9A0hqTgj2oR17ouqSkzVlQ8NW5TGHqZ9fbW1rUY7eZf2LiI3
cHNhV2j9tYkpuw6AbtvOUn/JivscqEHhe9AStIeVNWFSmy04B61mX0ym5j7s
Guj1gFwmWTk6cIkmZtUBbLbSyt/hIZmFEKtytK7HW/Xr2DXG0oFKrCAmSB/C
gFsJ8vJINmeU6OeLQXlVD792JWoBspzSBGJswCyOmwCAkeVD92MvGH0pULQB
lcARg/W0quc5kuQc/J7kAsku5kat0k4zrsDhuwfjODGKCJ+vSNxTM26Qwhoh
UXnMGARaZ1h5pDK1B2hZCN/3BYGm/vsWMhCxiDoAM76OHofLegI5BmwjpH1l
YMxv/zbQcSTajkhq2AsZNalUxugoTNIrjlexegwYxTV9leNKJdj4UOaFpGus
vyFIrfRIi2hQYpEqStmWCFJB4QanYfO93v2gHl7zaEYUWhKtDOtJD8/xY38j
IjBgfqjl2wBCROS7rvTxXundFyFUJ4N3guGt3cz+8atbzsjCt+2T20BDPx1j
FKiCgOwUU3ntMjxoBAGY14Aqlqnc8EYs2SFZGLU7z02S1fkdT277AqM59YTQ
5mXl+A/0BhwIj8GjkNY8mHFp06ZbVazxfZE3rGQCn1LJJmAIHlETXWL+DwUW
9Glx+fHnT1M3mCvLfnIPBDZPRm6KGqqiXGhhBWzAw+cKTJdp1VdIp7tSG8k1
8ltHdVpaclDaVBX76Ie6eNnzKGZZOXe1nfdlSLaJoPk5Vg/TEMtbo1May/Qj
2g9RYeuiF1QE8Jh2fsnc+pcYY9jVWVllfL6TPILYm+Xjc7ZsrWrRe4wvEiWB
3N/TZfgwjKFWlem3kAY88UnIvsdxfTeQpN00jAanFX5pgRIkSffvQEtInsD8
stVn+toH7BK+/93UwmWVijveP5pUFwPaPrbxrCQNuJ1i/BCNrzUTg6v1Reeo
wMmhV5PhnX9FSCBcEHb3LKCpgXpaHFIJ/+BDFUMnIcpgX3n6V7x+WktFd66A
kcX+MBTgN8QV5lvb/Xyt7qTPpNgR3nFGjTX2Zrw3hOafj5ErQ6YNWSIqNtL+
u8Hopf8zzD7JmiTMJJ+a48jrahHIzaxuHYQXII4YGhmwpKqqufkPajLGQR0N
pMOB/tubXq0ixZtKtzVbuh15Ean9kUTfSVxvawZnGdNjBnmURDD2aIg3RalJ
dCT2zVw83GzmHNSJl+mKLF938SpIgN1RT8rWMFtqHtpK1DrPLKEJ3Jg86P8i
WzJJmygm72qQrkC34hfLxz1FQwCGq1DfkkMCTvk1c/dVcheSXhQExG6oO5BZ
FabSKObct4cl9aurnfVeUPhC08dKYGrWAFfLXo+V8ROebphUP78ESx4PyR7m
OVb2EJseDpfb3KjoMg40r4tet2dQQgm+pLR0FpTWOh/eppsTB0PMTNjs8Qlf
KnV4SQuFZix3QNMvtqZFbB+/MKX6U8K3TfEUSrAc/71SLnfTVWqgPCfCM/zc
lf2VcTgv4sSFMAFi7jM+1fZyr4pYNpq+xeIaPjMiqi1EYbmCNTAlGht8TUPb
zLBHgfAqqjPyGLk/bh/tDm3q4jrnm6mtBIrnbMKi8PB3s09gdSEF4SpGydGK
u7EuwV8GlRjT54xrnmE1Q9qGV0EVh+fIF018S+cLUxo9HHQgBdsdBDPKgcR8
kW/kDShv7S3o0vanak6gdX6yhpxACu1LfUr0vMmDrcRTSznUqNgjj50owC6U
JsRvXMSrjB96osji2fMfrD5Vfq/5Llb2e/BSlv0AeHhSu3ADDVrxcdq/fuDp
eJu+WRQTh1AZjdhUEy6aHr+GjfX4BEUisw+YNQoleU2tkQsQA6j3tmpeNMow
+sS4iaoD9B+q6Gk3JkC7t5UNRQooY0zQ+aRtzUi4hgRNnlCZuDKMrF+h2pI6
idjVipdp5gP/EcZ6+W0jEAIbYfzyFjjxM6iZA8zff9goLIfSiyYEQjZXt6SM
UQQgbhsiJDJ7V9wM9C0xGcjzKTwpOf+FkvaaiGBoewz+SqPM9rSlnaKME262
3v5Qdo2aor7HJ08KLO519ahJ9l/nbfiU2wrE5X+nqNpJbddxyqYxvqhxgSR7
tHVGxyW59J5PJFCu3e2jyHLaTMx1UgnW+1dwPr3xkoO0fGwxK27Rlh4qBCZQ
dI0mUm0946l6lnRjlmM0J85y1qLN5j4Dcn+zDI/b+MhfK2tdIIRWC3P5ue2l
2OqFIg0Od1Ix5339cCHHwBeKiFFVaMIBIEpZHlJYvFAbZ6ucALpydG6gI5M6
ioNoQlHWJgHt52v0VHa7f+ROt8Ox6ls467kMxCTZDxyX7zavtn9ybGjf3Io9
j3CleI+xKTPq/b+LvrR+3f/XJoFEFiLU9BfYU7yZQ0DKbN9phIIIMu7YldjB
3H/B9z5BRQPJwJE04OIQFW3LahjRZqcMveSB7OMf0aRG6njlHIRh21yeEMmk
pYbRNxVLXTUq+6gIWFhppnag1MoT+AwSNocpJOrTPliJveCBT+RTsYWZAwlj
r0qU3Pv4Et6Yf7baTowvsXdy7NV5xngvCHObCuZmyTECI/dtTC0/A7m1HsEu
2cuR+YHKeOd0k8dr9NFaJIRxfq0GFpFVtif+TnwNqhfQXYKuXsC0MKCmFYDV
FVF/S5c7pVlkcsy84UGvt6HAQTWQWpOMdq9j++JuD1jfDbI1oN8S5AUqyzoK
N99jDrpYe424e/bRDh9nJcbft8XraYxbpPnhW97O6wcWKyX3ACKbvIpjGlwT
VA3UOTXsSY0xgars+msud/SNbdysweb34dezjUBYtDA2UtxYzHGflKIjYxtd
enfRPMEIwbtUqyrKv1F9NmkW4pzI01v1fZc4dRnwt0Sah9xbjB6c7uIBM5f3
UE+XsSYcWl1p/fGPtFFP0fk/SFBHn70AwFDYpc5Z4qi9uKaFc3YbJzW7r3Qf
fSmr3fOAXrQdY/vaUCRvCEEFKwDQR1sVAdLap8ibvmP1yEsHgHOCKytD+lOu
lKv43tD0SJoD2noGs58VXsA4j2bOixAwixrOOpdIDahltoMZ+UgbSmgXsQie
BuwxJTp6JLxQMJ3o6Wwb1DFq830NqQq9bnRiU6dAesyvYdvC13qTFY/2PZQ0
F/UrA/gWscfFjm40Y98VYslOZfJKfN2T9RgcpodoXR6rVPlPi456FLdnr6r1
j0W0ZosYgfD6H5JTBDYanWAeqUWfc1onqCgurP1rixJ92/vzV02GKaSUJmVb
BmV71dRTz1eCg7aoKlD6KEqshJU8t1SCdm/PZZsgeyxuQIeH/pfmTmrueo1W
LUVnDDHCVAiTdZ5k/CyStxPgNlZZLnoUoo1zffJpo0dr95r6D5I3HtO4Sl5Z
f+KoX0IMnTPMqOiws2Odd7UwRv0k9CDrGplOC0rfh3C9dBGTcml6DVw8xBrh
8wlGVquOwp+dBw/0evUbxy/syLqHPloZYo6Y3wkZAtzaA3KvwQTpeLWs1tp1
4mCtrXJkyvq3rTk21Gp1QQXgZc6RZLe34qMcidDzX71NGJ+0asA4OMx6l0CV
Ylp3Ziv5LNF86Ofkw1zkYBruoZ1NeYlqfBkxqkCVYockTDj9baF7WDqzbXKA
qoC9uN8vjJZPMdcoyafTKlHwJE0fACzhFUcb+d/H6Ifb3vR9ZZf5o7/gpWhz
Bm9EfVM8DQR08IS5IlZP88QcN4Mh+ZPIilkJe79GjJNUWgbX1sBk87tyWPHk
Pd69BHMOzEnn6OrwRc3lEigDPEJPakc60dFPtAHlO3icwIvcISpwGgP1azPV
SkB3BY478ufpEtx+85XT2LMGVcX1B4fLkeJxeSEBnl2kXS1onoRnxDWEMJiC
G2JZAv6AQyo57Ve2em+oBzJAvRiyxnj4RRiPGFlubDar3DQucg0ooIE/yWud
nZvqc3+AppJcT0TTKkMvqrpnvYhgvEGvbNQhFXODWbCmXtiWk5cxdocwtzFY
/nLtPzAJMOLOX7lPeeaU1svolbBMdw8zFwq49kKB/dXVBoxQf+GYNP/osujx
zsH9rgZJnZdPtM+WMtV+fRDdIsJH4rXvPT2Y6xvYhnpisfvZXK67najtOH93
sQmUAxnV1BZ8E/UQ2o0ThbSXqOwVzzaxiszR01ReFUREFVjPd6qghI49Rgp4
fSlAqJnfZ9Si9fNqdtzN4hCuJ+KaFEj9TCal8BPuQhxprZP5KaprANuUrrgV
7xQtGO3i0X7FcZlCjC0LXYRf+Pm3fkx2YUzE1+XJf2yHAAhS8n5t/87QwKJr
s+9gexoPmGAs2YUZ+tAwnFy7UOciRgys8hOLrTVcrJuHTa9N4ZRLOELfZ/nx
qRJzKtdjbtVbX61XaREF+gJUKFumHDpNAV4Ffb6NrQ75BUxJtiPIl8lSVaFt
OB7MO5dfZWFKroN3zxHHCfzOIi2gjjfs/ZsuV+0PU94DeTMN5dsoIVIZKD4s
ySYohvCEIyifWuA8o27W5QGzZRBfS2skC+ZtUqsjBEH00cfNXHMv/9wOkUje
8hW9nRhYOF6LvwhAULuTt75DsuQ8wMPcIFt+uVzsvGEEzyrbAxEu/VBewNzZ
XRLOCRxI8GonugrSnitJw3EU9Vy53KL6HtbYNC6juCdhV13BiO0IopfbOajk
gClqrJQO2uPHO0/HdkNQBavg9q9D9FR6TwXrsP+7ksvKuJ7IZstm7RbM6mnk
0qx4s5Inr/MjF7fR59l2dJHgBJ1oQnpmKg2Yz1AN3ZF6qZubBzKAzOEwyZxc
N/ZKrJYQI0ToAFjbXvDC/Vn3wKNuPRGJ7JcOqT/m/z4EmzQnHFtQkLnwo1F9
m3ZlvQk+0HDOnjlAhssVjuLDCKDJD27wI58X3M3NVilPZFeEA6cHrYR1MwC1
fyd+dvEwolTpYeBqTl+QtoZUhm3oX5DIkc/llYMPwBbnJs2hJseI0ALzA1uV
tlqZQpWDAU8hO4qkosfS+iwz7HdwrikLFqft0fnIoRTnnXcOR7k1HoyC0gVD
MuIffRSIuFuG9psbcWjm7slz32mvwKboY662cegoyKd3Ky5PoMcVgrITWqMK
QGLbJiaIopcfXa02BURDWR6ueZXsUWUga4k8VX0BRcxx8QJt+VVyhg7URMlo
y4rYEKgLhGo5E6AvMekMQPDUwcIOlrU6e8JV5X4nsJC/8vq+zY4MkAI0TcKT
0+KrLiSSwL8MPneFVDlz85kzgHQdrnHeQqWJKWGkZIha+WL+191/bYsOr9I6
O3W+vZRVB625Ohfy7RnOeHV0MnI3KIsy6xORZdG62DeZhsZQFLhDqosY1pPO
sa5SM4J/w1/2BjiyBSgSkdgROdRGZ0W0HPuxXWKbv4rq395eUiZcGuGHvBKT
u9DtcI21TyzhzOVox9n7u8/fjnT4MyNErd5s9ZkzsKpCHBMgkxKA3nKZMi/a
2YVDBOyrON7q3520nYFdSBEUcjndjZgNOqWbN8ttAwSRNaOZpP6Ni+SoNfnH
7V3ezXMoV/N475BLzDgyD9XFsA2oWizLINZ3m1BgJOqFbaOkxdW3pcFW+WeU
CjMOlueiViiVxAlyGGG+0xusHQzJ3RbG6Pf0UBbWt+kujWQACyFisFu32XZi
mMXkfMORyTfATqphfrbUalwcCjGg2kUS/9J8onXrzNhW9BRHlmaxy2ufXBiE
yhizRFya4lWlV55G8KZBN0NhKzc7msqAl02lTzCozje+xBEtOyggyPdwyh6R
XEOfa/xe1hys5InWGFpKrWIpqPnr3SCV5ENs/aujLSdD9OHJk/I4BhHR0KA9
VeaTZzz118RIUuw8Rjj2zQXy2NpYeNhh2/0RRbXQxXr6uyY0TfWVGnype5t6
Pj6a5t/T4aNdDmQ2WTBxhC6hAZ8mQsUBdgqhg2lbGU0qJkotfsMEHhbm0QN8
7ZBVaLRtoAzSo243HKxp6FBytWTjWbZelC+waNAzoWh9RDgweZibGa6EP6WI
U2XlEyz6gJov4tXasmhXn4ssGGA/zAqF2Qt5cR1ZAtOtdxgidCsawvNUCNwJ
24WAEQx6vDi/oce0uPAXhQZX5xrn7UKB/lb78Vti+QFWgTzw5JcdNWZDpp2g
mrgT0V4KemfFFbswKLpyHpsbmyzadXpBAzxlf/rvRNPKRJ0hYE7xqgSctaWv
SHTb0/pK5z6H0F0e0x6tJa37hhqoOPmRfU/UVBomVcqXSmP5bmNZut9omWPQ
hScLtRt/D4ou0kWt6IY9zfzphR9ZE0lA5UQvjGjMlLtUg8VVR9c9EylN4llW
QBBtAxEPTrT1Fk7fkgEoUHmZptaE13AAnwLNnOAVFHtvLKnEGujxUvzp5yAv
D2Khtbzk15arjqEpHbREPuz8Ec6EbiHt4Z/yZabYrNYoTIFQjXiNdCMQUVyr
W9VYxekprPIPj4P2OZqPWD8huqcLuC0nnf2JZXpuv5pLzjUyAzMvtWDUDC6z
NP/9Ft9dSz4L1clYx04nZRXoOmPlQDsgLQbtUtbKQH4LI45RcGSpGL02RNGS
3cA6UT81LsvYyyJguThWEzEuoczgD1iGmbsh7HczzTFqOzIBxnK6w1fVqSgJ
mszm5jfvJ34852D8Ej4rs54bk3cF4oHut8SrVUm7Ka3R+bgA7sNZMPJTRbQZ
lTPdl75tYd5paJCUev+whGxh8Zaf4YZJFPw0jtpf/YgyXo5kz/mMA0rTweZg
Y3bArb6UMA2FeLLMxv+Qo7Cz4kXe0RiHFY6LOdam8TcRnmZxXgV+rZiNDBk/
oaEgEijRR7/VbZZDF1hNnkY82RgStzRpx8PrP/8DmQOTTRF3ErY8/7EVTdra
lo9yav1V0ZMljGGycvJh7UFNxkEX5y1yCwkEoihp5fuxcqq8DD47esq8VBRO
kMe6hY4EWiShXTKYCxLdda8Pkf8LQTL3BAYA/goe/psjCyMQGlIXR3I4MLPe
kDLqxfVNLsC3BOgX3WM0j3+ycRwBOBZUtWS2upEYUBoQu+uWVUXB175B2V7D
hSqps8AdPALaBcvTHLRBmoCh3gx51vyBsr3N15IhXQuVqPMXg7YqnrHKpqYG
sSzDUVl5zwyMeQCX6ILoAxZyxiiiLF3lLr9usLZJJv3RHlQeDUjFFI0Waq/4
+sy26wZpC5lJVQqix2R+nvNxsVHG3qqz8KRNUIHt0QNOWSVol8YXT5CKtNw/
P4okuUkDXm4e12mDYsrRVhW5c3htuOOI2aLxBWSkoCoN0JinxNLy1kJuGVb6
vsFp/CD66HdaXO/qojJd4vbZZ5giZKcSUAgC9nLPEEca/NlsCZWuNGEFfhSq
vuGyTLLtOWCVF+yaN8uVF2ciQMQqmLtHNe1H0yhbc0yzUkZzSXpFkRHIgnrc
mzt56f/nIzhaI4CWjA2t1h1quvXvYjmQrBcrzYZiaN3w3JdV3NaVT9Mjy6nE
iiYa5IKSkE+ABW2uY5MSPgsbbwZYjejMnVqL46PtIeEpGO/3kG4gwnCQz/lh
rQnivzD6AEHfC5gOgTJxRI782ZKqdDqO9cNRl9gZJmp6snXN79atlEQO5lBE
PjRAHVDdN2lvA0lH4bWTtjlPC818GcXhdKb5w2BkNs/3RKniADq1vSc6eNU4
Z7Z5UEW95ihj4HGRNq6KV6rE2SMgO5Rf71wzSCY+rnAWOhnFIfIskLdWxB5s
itJXoQKgAQuNBcwFmJb4c7S2TwdxsbHVqI8gBfJeOUBWzvr/Au2DlcAodB0N
7jy1F/qpkz6z5YTgLDHkLYJ8ghBqWKOPEsW1nOVpgDLaMlIh3IY052OOdOEh
45taM0e7FwruLYaTGIrI+e4pWAglqmN9LA1BPKqfhBeLN19KiYpkqVaQH0Dw
TXtNUCP4Xq1EyUcief8E2dlGkdZA2CKWiMOd9D5cyVsroYHz0tOk5Cd/du9a
AKLmyFByqKVjztF3CIzjcBAhQ3v3HshYCKkiADhXUKJVS0bYC/fZq1A+p7X/
slfA2WDX8fBZ4W+ReWnfkN/ftsDjXIbfhNUtvW4KYbuRFR++7fzY0toe41Y0
hqTgNK7lepwBVhv9NzU3Nq9TDHNUyeBStaOU8kKCZIBvkweDkOQSUctXnSfx
5XTssU1JkN+3J0ZoGf8r58oUH689a7o+XBWq9+s=

`pragma protect end_protected
