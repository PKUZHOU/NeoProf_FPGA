`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
Nj/wUn47GQFrVFo8bsAd3DvMSNYB/TDvpZzLXTx/4ScUjHh2neOwjCK22+kBdogD
oHI8+aCIP8NG2q9VxDxi6AaQvb3/CUNo5MVl6RkeyKfuc9ECavfkcKNVTfd87YJ8
WSmmUIgGztHlII9ewHkgK5HGznJEnDtx/QownlRj8l0=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 20080), data_block
vZQYmJYFJ4YxYTn7+Bk6YZVvbqn4B0UqST3XiescElbL5+ybBpbdUI0TFkUypwgc
8CN40jSmmCIX+9n4wdxs+wbj+4oUsfLU3FkEtOB1shJ5oHWCoKiWkrHjBNBoW1FE
t5TAc/+0t8Henc8nncv4zDej/v9NmJjg6pTJLNWxujKw9wfut8xZySQ4o2gMEnUM
LSYixYkpGjVP8y137jMgLtTaMeq/W+0qlUKG6vPLf0uYii50eWk47asH0k2CLiPo
h6RYLaQgoRZBRB+GQlyRmuddXt3b62eUoxBuUyH9VjWoEfPwV3sEcGMFHgXguJvR
Iii9EmqmkQUSZ9cvwFfnVuwRTz3UooHc90VAsM0FuIf2+lGiozRxBcA4F2zZPT4/
riFTA54DUiOz1XGw291vNAP4JbJacdN1NMSodEhV4sKwjyuHVJ3KK5EiF4SbgK41
kI+ytLn7jxEbQ8ki/JsAOwX1kQ74nYDoQj0+Dul+vB1s22HurKA9zhSO/lwL2Lcm
0IKu893hPPfhR8RYhn6Sx6ueAO5fEjpJvdVlF16y+ifqtrBmt8isUy6IUKSNNd4l
GD8g8fOwixG2MrITwhN9Ym5wgKUci5C8QH7i7iJPjjbhKGfZQClgUlc1BpC7MOG/
uBnldRgkVCqvRZLHUuolSgPAUBPEfk+P5JFnrKAffXdgRzV73kTHY9jUr2d36tOM
WD1/VLKmKWzFtcPKE/zjqCvRKLvQvfRRSvbKkhJJlXbVy0H6/dRGYZK67sWYO41R
8sm4dYl++/ppOkOX/5S6OfDJGjT72ThQJAOBr1+BKS1CW6uDvy1wx0KNpcm5N4Sl
viNCgeE4tiuuzzMc1laCe25iGQmbscT0Xz3GXBlTKLFxUpiRN0MKBKyjKvzre02n
pCnw1whv3jundATKkKT2D4mtMR7YIwXtqhHKwc0ywDvn3JwNEVDqn/kMjJupVgX0
CJY1VW+fCzHDvfK1IRYIkOKhItF0W7XEVq2mkXJSavBcRy7n7P6QPOeG4ZEAT217
Fp03DXZfrJs7svtgUe6ClnhIw8Vww1e8EBtt3P4nmxjjwcShzjjWm329F16lrMU7
KrcthU3wYSg9Fd2Q7i0al6Hu/mZZgf1pqh4EB7rcoKqLt/eP85uSDJFiYXZ+vThz
G+LW4rH47ALkeZDGlMo7gjtGfX8LnsagaoX+wzD71siprkjZFBCZ96TK5JRhRCuX
3xAH+1xBKse4rXgR0t1e2ENlH9GK/yZNAd3rGfKb9Q9LrydmNlBgMqKCQ32YXvWU
SP9k2qMLz4ghFPfYPrmERzq1yTqaR2TV88Zvl627/Bca64gYEWa0EBzJBc/+JDmV
gU9iQDYaKQlcr+Fq2V16dxi4k63iv5D+dfK4VrukR0U1qfe5+HigY0LvEgH6itdM
zEuA+5iMoYwOZsiDa+QF1GL8iN+eYgutU1SdtQxZAaB3JhGDg9B8HjEpwo2P6VZG
7SIVRsR6UQX1ai6lMdvyXeq92YJ+U4IESZJoogorTc4nSmdSF+G11WY0h3gbzDSH
tEsJiCKtsTfgc1MEaXCUuHBzJDGI4IIHXlpUCAE801jLmFtxJW/qgsM9VcFCKwj0
sSsOUYa9M9jgPkkHiPJHv5jUZhpA/5vglKXsD/2domgL7+3KJ3vh7DsNN87DT3Do
eXYiAa6gwsJq1ksbdxlskH0BijrVwo6afgQx+uDBbBInSWT2vtoNK0VeW2US6DZ/
2O6+GZzJuyhKzTMUeDEr9BQSksaFLOwfz90CXl9mmOFrvjOTDMGybhBsH/OPywQe
omQnfrUADQ961vZnv9CMqGCPJgYMNXLZsllapP9XmsCQmR/g/qEmL6akmQQqClcG
h5vqsEkEYll00BXG9sozO/IIYSno5L57mOWNpyqUTPXhFvlbvvDbZV/W3/hj6zVr
iiZTow5Dm00ngX6MOIlGGZd5+hvko4rgGlwHEuAltO9coQYdx47Bku3b/8XNW7z6
sg3mJFnY/DvdHL5VsjY4lbEdIV4EAsu1iAH5sP95NV8372QxpcneXCkUEiYCnwqo
tEjeSB7frJOy0xJ+jY5cUIDltijrZEJBKchEXYHnnNxyQQq4iVbPYMiQEZ/6tTyS
sKYpvP3DQk0aMPuCz24R5O9mItNmoFf3tZaDdqId7lwDQwhwLgqlSfpcbwrvWy+6
c2CZ8y+pV6rW4AYmPn5taVBj0SQjJTqofpohqbwwU1KPCGLlbx4pPUqZdi5q/l18
7EA1r9uMzdYB7aCszAOlEuGzNKjIuwWpfVRR5w8P4qQo2nTbDC5WXD05Olny6Gnn
Gwta10CRPJMAQqasB11rJrWioRSTFhPqbQt9qMaG7qbZuhF0VYK+1sO+Xx4ewh4J
O6n60fwkQO+xeKOM4rxYpxZYVSPsMAQhqNKiwEqCzE2n4AnADA5t2me1QD6YCsd9
A7dnCtsPtzENbiwK42tzkFRkmsaWnYuR3xKX9bmuS/hhKpnyVYJ1octRJHb6HAnO
PBlY4cXZbTgvCRXDWo9KctYmQFB+oAbYVgKanXIA4fsOD5mNkCgCbUV9dULD1h/k
abU5BFkXnjnTSzxGxt06T97J1bFa9C4KHPZptq3vef0lkTeu0HjZg3MIE0Zam6VM
Wv6P7K4jqWmLOBbH8yFe2Pjj5UEdLhJWnWYPjB7UYgs/OwUTXVBGVk2cKf6DwSUM
sL88AneLQ2nMJOlB+6bwbvxl3AlU9qQvYv1RQaZPFlGtoRfYPmS1u5SiDIHndsKM
gdBQ5o40NvVwuFq+qsjhPuAd9qeBzHtpX/xjnN3g8mURejPD1BfVM2fYrENC8f6/
5p/lqlH4x1Vl+U3gWhKr3pbA+GEtTnOAzjTTwUh1zt3tM7ZEm8epJW4AYMeTxvCa
d50tkVMB5Dn8By4hOmQiHhQ8tXlFltbehme3WcOwv8hFNLoVDol0ycrSSAA3ZMwF
ekfpqllBeQSoY7Edsyl5Q4VZo5YynJdEMhx2V4FEiUTPj12GqgSxJMhMVgk05Z30
q3S29xs5IuhKiA+7e8ch+C6E8dc58BuJWIk1KaiQ9pB0ycGmVcOVLmexUlwJtGGo
O1P1YB7EBFZ6u24IzY9r+kc4ZSwbTneSoNRH8iv2eyRMiRu542RHmh4kKs7gHN78
/zs4M6TDZ1HFPPS0yjdoWupEtj5qNE9kE2uLd+6L1s285I0ZZe3wv4Xp3ekS6c/B
OqhLx+b0MDt/LBFGJmNmPx5u8x5fpsBkCLHwvn3E/gs8Mok5mjP7pUZZdUI/HrLi
tCpcwlpbwiFayM0vLL1MNn4jttkYgLeaxTsZIJhIVhEBp1WEwo6PkgfIU6XS0kqF
/SpYmiqpSnMHLCu5VIAUWsuSL2wkvJAKSm8hPKnEnn0F8B/uO+Bz5cRBx3NoL4f6
mDV3jPDnqWZ9EZTDPditE9h+kQ9SP6anKK8p4Bgb5rlw1Cr1fI0YrUgXgQARJgzo
QDka1XqpPsbzAhtAE/tTilB4X7zd1h22QWKBzfju/38SfrmQ2DJ4/dtCGfIhP+b8
+f2kdehoyknmS3cpM1zrQfK9LWetupwRnFs5aAa1jd0UUHo8ek68MhmoQuU94hew
mosSX2d8HOvjVzQn0WQy6LdTNa1sR0zYhqnKOawVJhmZ/1DynOvfKczFhxdJn8vU
XGaa0GOQYuD5rESyIHu0kcJU6CYCAYtVtDoPv3vGacBwjQQWhx4rl3Qks6nfY4iA
CCZEeh7+v19xRDeAZyLuNVxCHvb4fMuOSQw7EvnoYqstAHN5WhFEyoKlCYJ0oI9b
r31jx+UxQf7n8P/l+NMU/MYmhtymMwYjSQpZL4yEEBNqAoyyvWDuhSIVRZErxZ20
DMTJBWkMjmseRe8ZsfP2mBkrQPbOv9XqigUKP9K6GQGPiaqAhLltJ22asaaqXEmH
TOpZ56IXF1kucLfWVGvQkHeCIvEEM0ENluej8jjLqkuSSlPiXbfCk+gRLEOw6m5M
xHg4ojnGJes37bHYPkdjK2xnY8jk/5JPEhVLYZUv8dTKUjogw4j++OAq5S4Wo/l6
8Kv6qqyIyMOo3qcwkjccY3RNBu+MhJ+mB9YbzcwJli2qgJHcuDAwA5pabwRbVc7C
wL08sIqvG5JWIJMViz9fWhZf18jpTDrxc28/OdbRkm4nYM4agFq6VVMKvfN+tvJT
NBRpTUc/7gWYivW0oPYuPlcoOZWyndDm4bBsc+v8HQXFUbD76sgeZIg7vlQqvAz5
WNrwguoPW8JHad4pVnlHUqn+dZr97vdBW+L4YCnwsXNSKwXGmcrGkoFJDyCU98DQ
aeKxTQcjDPjdTBGT62Kw8VSuqPsg0NORCX3jreMrEeD/oKl6TyJuumivzmuZ6T9q
AwLoR+jtuqBCKdVWQp+38nDssBzmy5oN/npU/7xNp2BtNFnI8g6Z0BvnHuIVS8Gf
QjdZzQrDMtLEsccjO34E4g8yY6xNHsSgEqQNSZm7G7MGn9tjbWRwqRBhUivZq/6C
oxBVPqzghlCUbhSOgkUlAIrUsXeZao5JeRK4IZ8Z74XYdwjVnV0SyIATXsrb2h9V
By3dtSDHLxkvLN6vg3mIdVg6pv5QWdeFNetFLIfiP9wxm6hgBDV/wLaXbszAetFw
H6nP7cH4imrrdVxHHydtzAuuGhFAsW2L+MMAoAMmyOLTTJOAp+Cqz1DMUh7gQjEO
akL3DizYnt9/f56ohPqN8U5Bq/mPz+DcMLkRKNgutSBLZ8gHlTytiNkBDE+etm9Y
mwA56oMqfKO4TG2yYeMdw/7IF56x3bzzqpQGpactDxFgV/IaraFLujPy54sephm3
lX6BkmH/9etUBjbbW6hPRyoE9fOcLSNPNIutiYERXmj7eyg+3RgAaWUrU1vM8Dum
G2V9qGNOZNXO10eycBXUAdlKBgHWyqbqCHP9H/Eo08+GGB1y9Hxd4iNSHc1/Lcvb
EHxy3JMHosznuT8jxA94KdIALDRvQW9W+R6TeHQWrMtay3eOhhNKT9hZ2F0pwjoS
yulG6US/Azt52o5o50BZbC2zyR1fP2bmnljGTJc/6emNrsyVJvDEHfw20AMJ6Z0c
mn5BHXRddbry5aN/aCuup8dfrBdegXPwSxs6E8aRNWsNH4SapFBTJ5Yuq3zvaObx
p1WzwTXTwDslBtV3nKGFMgkqEohyFaebiMzOjNPv2zI9q7NNocPYajnYC8lPNVzi
2xmtN8WmUivuDOwDv2IntqGzgHhh+iDXu1PY0TKvN5RFMinQLwClWoWnUg3azxia
LM4NXvS+tfiqTv2E4LSYAhg1UjEgd6tQxf1JPp0baeJyKtkkm3gsaolLF+N3LaBo
2Z4/di4u/IQUNcyHrHKfW/9j+GI0c1CjXMPdq9ZhxjsIZy1kUX8ai3igP0qxGwdP
vRjG276KQqS60eUrgPgaGclY0FNRERogHiPQW5YbeTEGSl6WkgPzBvwVBRVG8ryc
ZtL3+fulFcJF22RQ4QNN8EChEbbQvHlGpvImgCWW3yc8rKpW+01ff1WH1P8o0URI
dVAOZM9Zz6+1du8Odd1iLw6qmf5T4qN5wNC99ZFJt8mNuFGdjN0edKflsIjRSAub
5dXBaAAdGvCU8ahPPHHXcAo4cEcqB0p/uqLt/unN5VOTHYbkLQYlUtFOE54PDGB3
OQzDB/LHRCKmIfDQHTYWYczgtDmEszuaJuQTa/iuvwrvTRWYkp5BynyEGr+j7FSv
ZWT0WJNzGOOJ887PRdZmhYP7JIUdukIj39oyOFjLp2zKOBBtjFo90HuSodVVWXZM
SdOSMwl9E6fRH1D6BeCRCd64r57GIT32RR8Mb4xNqBPexCVkwnssIRqYUrbhWAdJ
XAZk0/uOHk8hHWBuLEqIXtFz/aH8msHatNSnVTBE0UOTWkUxazNTATa70vUr8Uli
P//ps7BE5uppUEip7fHoj3msLofEx6ORaDzkAl99jKHsuDS+EMnxBpSdh3CZn8Wu
nVB8wzO1mzLuz6vEbd9NMcJPyMfRAMxUGpXDNFRSstGhYLeLUNKszcrBhlgB2iPK
DIX9ulJT+Qq8lqYctxga4CnlYAUHLKGrCVPcuakc196g9pziR5FK0VzhG7RAYQIp
I4BGOtzVh/+zGczypVoXBNfO87ziQBDPc+Ry0Ndx+SLWhuesTQnBo5VuW1brZ1Wz
6Fzi4rvGgaJqh2rolvHOL3NZhM13muBkx6hC60Ouzc4wvWQrybIErbW+efjomIxy
cUKWMlIHIiEcbHswWVVl9iifsi9GNO4ZZYW/bBJVOPwrwZ9GQcvSPobCHAksqobE
1Gum7RgPFY4YR35CuZJ2MrMsRo08h2UtP3hS7ZZ30q61sYGDugK53BHa6pxTGvEq
44SoEVOMgSLf57oaSlchR12v69E+w84zmp0L+ZIgTozcAV6B3EnzE/VJWzEi0Szb
WLOXXb+FH6cuMniPpvSOr3T8ZeEoC3B/VK9JartToBKsbctWwGN8wWGIuc65H95+
jfaeWDNw2XF6HXu5COGZ47O6t5/38raggdT4jxmtoqgeLm6ih0hm2dIZ8XH1qlgl
lqXAxjNoda60Z0h1nBg2F6yub72GUG4yErUkJf1fy60EZfKXuCB2Xg+98ty2uaqL
UO1znClfO+bEiVlYcxIyXVluKWvFSTPB7XjmKiCiJRDvOO9xIpej0iH8/oV6Ulp2
Afv2d90rRxKlddjpA4vcV8mRb+/V2Y2uM+tisixr+qoivV6t5rWcRiCFPZSmOKVZ
8AAq6+HF6CUcS5qNSq+f+wYGzoBqoqKi74ewG5PLCuEdARjUsbnv0FfFgbc3sh0B
6W5vKqayg7TzCSCJT3pzG7SOIB+Id5mTN6RXERAg7c5v9Perbbw9dH9DjnC7N7r1
Y7JJ3AGV08OH5wwgoYGKWs4+N1qL6oqUjT3x+DGJ+rgaUxBdgRiN0CD0ov0H0KNM
FU/g0afemmeKJIVnAIqPYHI7oACWsvGcvdC8PmRQ4BheA7ONi2Z7Q7A/cYyr/fVd
QwDet5NLUAO6DGXz2v4xEpi9DeBHJmeBJwbjXaABlKKjvxOH7A9+Hg/eCHWgx8mc
Unz8YPYZW0ZuE6E7Dg5YOfxOTYSvRNGZDqWCjowbHbJ+ctJrbdq1UIutZ4d6IvCJ
F1KKT6CLrVWTFxPscf3oC2UXR+93uvvwd3I9+KBQu1hj1HgrOqjRudn25BXOaGmx
9xhvgl/Bx6Gpr/VPf6JJ7IjlcRcS9dD1UvFFPblGY8DR00RO0ubHsYk8nJ6ef+kh
3hO8vsPmsz8HCUQTHhEpP/hxvpOnA73siCT8jEAQDGdXuaZKpzSMaHeVAwke4tEh
PlC4tQNRYXunmBM+7goxHviwVIacyk5rufGrlQWlQrvBp3NSaRBxhnrh++HL4/hh
NbbZLg8SoVVaDOLPd+a0gWy+y4q7ZZqM+jQRx+FPjM3J6jCUrViN2OABFj84hKOy
ZjniiKocHfqKQhvzU/nb7G8RVSJrSy92QVhw1Rsj+3jfBMiH+Jdutb78/JVyFF5s
J+cvkcpwqlBv5CoWKPvuUReDAkO/iMYlvNguKU+Z0IT1BZ1MIb0p2FHSkTQMsRbf
wcwLFunvvlOzBkiln52tnbpYpAMTb6vBspd2O189gc7bPqxOIWwlzGQOEX8QpF5+
DQ9PF8WgUkFIelbLMnRuXzTPIn87hA0Jhy759+BQL+KnCkTNrXBD6bveCvKJStqq
/tyR5uoNDJ33LnnU02uUl+EnNKKQhXVPi9ACafp2kK4gqh+uB3CXbEsk8m4sdJCF
sVe0DjIgGunc8dDk8RqfzdQPR6Sj1+xagVwKDrxmc483dzeigLQh7+imfNyq4VoQ
LP752CjOxHrcANWvFx8OiJRTapj2td2muYGmSrzlBHHVxktQIG+6tWRGnwgLpwWb
nCILl801w3gROgpUGd5VyC3q6mNweXWJJaYrV+g7WCQnfOAccaVwslQ2YMSau2k4
g7UG9T+JJpw4EGJ9hVw3KVAck9iyEFP/NYaGM6nf2/YC9agabTJ6rgPgsFzA+xmA
dE5t0VNisOyzVLIF6ARyGMpMKYwcOEQ3BRyL4mxThMGj/C28kXcre+2RCcQPME10
E/qq0G4ixWnBE0pAwkPh+GdAQdrzb9hz3ehpw6r4p1E5rZoYV/3tkfK/fQtJ8wxa
p+w3R0oN+3YCXz6i+wcEjPpxJrBZijb9aU/p3ZapqZQK1kt6mVjPXw84HDdqOLKB
Niy0B4VWiJfYjChywrXaloO7xDyxWsNPy2QE7ZwIunrSxLNDeMw59Qp4uIOsEbaZ
5sFucMFlnAeJhrGVIKhiW7zz+6jpv47A7uSihz3CSmVsaoMHMXSDw24NNEi7F9Kl
4by91V2dHg2KeI337PJvUFAgWixYu9LwYlo+9byOML+kKYjJaXzB1OOzDAmG3fsX
8yFUFicOdLpIKVhdZf+VPgxsMXPAA6KFikPFl+CUwkMHmFMFB3hvT/d9Guqa8SP4
54lJou4f59ANtpIhNhAg95nG0KBZ+Y1GTPUtI5DJ3uLmzY0LpuzUoKOkAYhoo4t3
gLv/xOzwQjQ4NEEuYrzOV350d9sY6KbeLUM1YnbYbDq953MjxbDNt039o4I2nbuE
67OOUNiict6qsDiVT+mr4R8fnlFwQpuOQwq/kRzRmFEgGulZddBqEeOGFZfTPrms
LvLBcGU6TKKVtJhq3pb6lYzC4DSXHAuzduCHvZ4vhihTjlBuw68cUX/jVDNcFBD3
IjtGd807NgAFWJGOEg6/2+cFJW0RVSfqP65lMBDS2BxNUQqMITP3ra/O7rxOjB9+
FlyAL+myMIpc8cm7qFQaZvxZw0wJ8F/3fKK09A9xev4UoTTjYhgjgtCB/D4khejo
7PmztJsgwha0XrhGRac8ip22wy5Mz7NjU1r1cdNwZDXW28GhSgJTWeiQZnHcpA6E
i8vBceU2j/I8q6+08c5iN4B4Yg0NFm4UvKJQ1Qt1dCsPrNpunPziE4asgOSpKq03
33fyWD/2J/wtSMR+Trqr//MhZSSpbEtK6gqtz1RnM5BCUH56aFG3/JPcR4DykZa+
hMQ9CjQhUzHuGhLhckAhbYuNjo+mO2eOOzd4wWMHPfP8/EjFTrTx9tD6WRvkPuJs
hkhpoLbwW2x1s89tOZfzdwNAMt/uMuvJdk9Hh2zWG3+9aZQKteGZF+HqRCJlL+I1
y+Z6BH6UvSNfc2dOO3r2b8T7In1yHPFxdYKyu4jwKDD1fc7BNpP8TA0a5j0CO4+C
QdGdFFghwlI8AQe7wmLUjAFRbRBijlxZyf4uqfdl7FhdD2ZTHkeEsSyC1yyYcdV7
kBbSLfsHBwehU3A2ph//bZzqgm/TIAzoYA3zLNmxtSJWWc0MimuQF53PcG1x4XB+
zRRAtWAdmBoi3yuf4Rma/Ck1R9BNtiHxTk2sc8lmPK6O5NRNraOuBY2HOKrWb8cH
Yn/TYIO9AS2RzliOG14IlxzMuvGHmicT7i6x1CmnV3Hs0BNSSxjahzmMe/DxIWfW
P3PVPUzpYeOT0HT1OAZn3IoTLDoOKivW6EzmI904rplNosfXq1VhqQS2lLGKO337
s5Yp1DjxHvr5/KzchJcs3JYGSHtSIionNK4KAuz48OlCZtf1Jt4O6pHoaRj3+DwE
hXX9D6ClSUB66W6NvpudIrQuIYGvcMwD1Fxea3YJX87fl6afIpAwIrXnBAOtDEIh
CzgMOvzvb9hL72JtHPjfe5la5ZUe/Gu1oQ/isYCZD/IOtwqSpzgbfC4Dwyfv4vZz
UDcHW6MhI7/e+8wnifEkoEXPZgR+egQzRqsnxZPrSTvF3klFKPfUfli07a1hqPE0
MvcCSn22Lv4eTSgrUL46BSoWVLE07p175egZMn2akFckoYo8U5Y8dL5VcMUlf3w6
DQQbzDpXQSOh6u3YZbwqy8tr2D0WOgH+n/dDKOZV5wJ+dCBNcG9tFREr+RlnJtNp
IXO4zP8M4qvVOZkF9mJ/SWH3Dc8VQP7i1Rv1mVzUK+TQ+cMbgZpG2w20TP/BX4KF
Y5IsADwqztEYjJPW3dIX0wDnnjd88mbOFj8GuTajVPX3pPneoPoT2uMvAx/XQ79C
tW8O9W/5oA1cADB+KJWh+VPhGteYJ9weZRaA12heLu/bEV/VPx0BaLdoEb1CNLKF
WEdGnL3MLhH53TwQfT0oscVGEO8gY2HCcltPnmYD+XLt1lDwbqI4AGggyQaAIbXa
pH1OB0KSYb82GycdeIR40uZpyFtfvBMnzKrLDtgG60nihEcYhEbRJifNcAIcbmvQ
AV6mWmAJv/lYFOEMbaN/PG9L6xAx/Z0HADFDevg7OEbauaWMIjAyyEbrqh4a9JJR
MtDtCrlVuYcFSbqNRk95I8DjgWtIcBGS58XZooyhqCDbbK0V02wjWzJfH+VQER8r
h4ATimm87HnmR2/fvJmez1Xwyjyzr1/4V4pneApDk6s+OxORSjiH0uSM+NB5oP3p
y8/GGTxE9rBpjOsHKfo7rdaLWwOdxdxUMlTbAMc+clLHz8eNwfQpZKlRzeQSjG5k
CSRYP8AyH7p33EWobLDMAUOQADVycc0civ2X8UrZE/gSr3uPn+ymm3Lfl+2bkyQn
pl2iT2fmG5WfTiqOiEPK+iQJPCHCIqLaohrvOUPELyRHTGlUHQvBY/03tKXL6Eix
DG9ypsynQG29f3A2Jjgxg94MLO6Gk+BrNCCeq9RH4Lw3psw8cnYBC0DhULOJs7CA
vVaivA99m8wluzGSade2s4u+z8t1k1BPEbQOEK2t6pCWd5FR6R6NUSAD3zG22Oio
7weqwlNAlI8gI77r6uNJ6A981mhmrDUv1cXFUkGYLdRolrCnSTxPHcRWaFLJ+IUT
UR0hEY2iZozTAFxoPdU/qChrEw9NWgM/SoSGw83D3nCUY4b6G167WIKBrReoePME
RrYq5sGkXDVQHpgsXLLBri0rnSDWK/beKbpbajRNHBAOojhlXXAVoGnWn2K4dxw3
i4NIc6tBekebz7nxK0NDR30JKP34pN3y1Kuo1b/T57QMS71U1Fmp2qm7inWaeFOK
Nit6me9aG7vn7U7LxvqO586TM9Xp2Ll4QQJCG1+qOHL0+neK79S1/sijg4SIiBK9
Tzievz88YC9uUTVE5zBoungxhkoculLf1ZtMWSGSEcOgkEf7if+5HaDVxbzs/H5A
qn1jbCvdlTdbEYes7jpuXQR5ddQE5mD1G9eurq2UG1bz5VxIj1+GG/TU3buOuhv6
TH89ywXTb6z8t8nPJE+IoOZM4QtllnkoqTO92nOiUgCHMwgG2kfMsxF80o+H8Nac
CaFJyOtzgkxlauYfd0nkX74enAEKC8aRujkYhBRm2CkrmQR3YE0zaGViDkNe2Eow
+xbd0NEMJWr1QB/BNiIPu962fOFopqEVFolhb4eoAbIOKvSY+vKTxB/HSObrJIXQ
tnfc0LLeoMggSKl02HFo1AnfMtweC7nVkQTe7mJ5vf0GoelE7Dc8bdArk3IOw1Ol
zp+XkZGqsEpC66SdxJ2+Qz82eA8ECKiZ8fFzAvAJBD5F/VwEJ57lQafdYvDkUr+h
JGUbnLq4CUv7BXkxE09KdqEpOl8reNtX6Bq9wQDYuTJCNrPrQFRa19+5LKKahB4U
JTnBh6OuWEmzy8AVr/1OVvOnUebeFtrY2RGLRCkOmXlG0ImHvHEHeQ28C5L7Qckc
dhPoA13R4aJW8T5poFh8tUt6vFExUwOlxmoSPh8ylnNt+UZSdKyTUd5Kg76oPb59
3cV5EjCaQP0Jpmzvkeh9onRh6cUXkuogcisJRAUENn1MP8+eCoa0FeaIWcRO1eI8
cBjGezjaWIObChwGVoGdIWQyJ0+dh+wzi2KssdhzADBjyL10gLoOar9yHAVOMVtJ
jSAyKo2eApLw9Ex3bPDHBsfdPZRZEKndT/SmVTP/w9brx31+02Q+HnopLoygh4TI
syChvg9L5yTgHfsGOPRCAwSDhDDjSOE6ayBQoiaELQxrg6cu9IUUOhZ7Fw/xWuuS
tSdrfxWoK57cJnflMy+io7j7oyNWZR6PQX7zvXieaxwHpdKWbx+xTifCq4Lv7uwx
jh9bNSC2UtOG1myGpFIa96DgWsPkOxh2pk4mOlD/1qDm298ZVVasSq3jQnL2bgcg
CU6UuxWigztfpgzvO+WYGdndTfIiS900jvyLhFJydHdpAWz8PbbkN2Uc8TQectVS
KjsKGgcy+Slv83SlE4hlfAkIAs3HPEbUi70zFHbWUUG2S1WJMXHcjgzQL+hNEqzR
q3nF8Fjn+wMOttlRLh4eOkVrdQLh62FibauIw/FHYgVhBXAihzwskysm0lvyvt+c
wJc7UByQXLzX+vmifbvvsIaKZZrtZnkjbqII/KpsPzaPRpGtuHODR6T/RRr/VUG3
qE6SZX6gp7vEFeeAV4P1WElgQApGUP9N1e7y68tcOonhfZy9NsJhdrusRzdM7Dv1
M8fPtHtD9zceVs/vP/BTlYcgddvSJlXNcbKGwPLwGW0YDImknWXkyC5e0oYPjbw+
OqyRJDg1Lb5JpTXk3BZo4h2WL5TtJehTfC7WRRd03N/FfHGRY3pPRBXL8TfYoSFB
rYc3OSH1u00Zj0WXASiI7XUjgHsyWZ+7puTGp4oXQzpDdlTmSCTkikndtnXmIU6a
R2ShIOpH7qKd9H2xvKwqSsvFePI563/Rg1wRcvHb8Ws3Xbz9Ef3vE/hBX4I/9qC/
bMaQdKb0LgbNoW6AcbS6U/bzuFebsDaRBLWXJ/RXi8QQAxxt+3riDbGyQQBPgZ/k
C5WsRvTfg7QktMgVAdXW3dLdqiCyYyMhNkb7Hs7j/rCsoy5kL2QYCUqT1Z9Ed9aS
OGy0B97MhQUld/lNN9ZRrOMGO3dtJP1buK7FIBeztyFGNcvgzTHXV7EI7kBkY9B6
IsloQ57CwCt4yBFqMP+BpSSYqlQLsezv58H5jCmlIGsHqtHW+8eU2eeSIBUfRO2p
4409HAhFEFW9J7E93zHDn4j228YcNyiHdJ/C6+mruj6qnWvye3S1ZQgWIi4LdPQw
fU4FApVxU0w+wBaKcnw0kdKlhrfZ/LWTby3+xAO9JrLkWulBthxH9DAltD9HSPt3
yFeaK9+J0UoTKI0R6JmyaSaeOkIpSLHwf1Q1LvxSXoHjSgt5+/4LFZTTZBrA6CYW
ss8dIJxLgHfILSXYK9Vzzthwp6Nhnaqmw24ABGZplhV/N5y5XzE20Ecdrpvkfqx5
dfDrMe5DcadgCyPedWsr9WURdnf/nT3+Okvlbjsl7GFPzHHjPDuy66p+n299+Tlz
uPKCkOxUwyK1hWa7jM9Fx1AcJYFcgtYqUih4+F5j3OqoG2PJe6NEyABIlozUSuhz
AZTpNGKCqScO/oiLp8iSz5DBJW5C5Mjf+bSFD1qPOIbudIg+L+9udkpjHLA4cD9n
+pOjJBP3jI8e94Ed79ITAC9EHMApn/c9p+hblSQGUgBaKglzbpgOXJtja3xzXoFd
s5M+O0brEhWl5euAHEECgtGO7Q90GcfIfSPp6MJf2rOPZNBRrjmu5Y8qBmSrhkgt
DmvKUM7dL+vYSaQZejtaajDmYZUGq4RLPYwNxmYH4ufzHyWN5Bt39dQgOvrHW3uR
ARIwZhqQZkOaA7psS8XzErRS7umE0kaJ10PjGIZjRc/BKnKcLzn5a/XohE3m+6G5
YvxIAi2fPRKZe1vvquobd8oH9+NB/j5HghiPtlODL7rIy68qlr0yF0LcAJbdDXmI
y8lszm8G3mVGoELjlJvUoteCQ1l0QtgJy/jx/tX4ejbz0TxV0JEcn9/zteD6yv2C
EHcYh3/dTKz2jWlXQel4iXjFe+gfrfL+6KvfhmiBfEg+Ok0tRpQ8KDr5Gmcib6CG
6alahesIrB+aAWls2jW9JMp7GDPBNNbTO1TIBBuZ2ryZeKYCBGWNYN3tZXsxPpNk
31HHMMdaEB3MleYKpv6ugskpLOrU60zJ7PWJSYmgm5Gr2BBgWGCVpQWgPiqTS8QF
714OArnv1DCl3yQO/K+KiVoByNtqLUhRzVz6KkIOcHmxNepIvLMmjhiYeqR42oJU
UDAcWKsB6PMDZgf/adCgOa24ih2U3jYh1ArFWRS7WlHfFnWnF4lSd1/2/CmcWB46
iqEy//MUk+cbgrkT0W3ZYWBZU5SxXClWqBUIi8UZK8cBTfrac1B0+ERTC/kYzG1j
94T7aK0xTf1rK9Y1ObSnVL1I2l2jCHNUFPDQFYQNn22MkTjtrzArnEWdmEEKRh7z
TxXwkWOJYSVLZyPyrIdZ/EFJFB3/tshtidIx94Q9KnogHYnkLQrCtZuheuQ3Q/Hw
D9leCfeqrVkr690DYlX2r3y3TAjPyhySQe+Xgu2WRdsFRnjOTD7sjI0VQCN2A0fd
Ta6hxOnXZBMl0k+m/wAn88jGOLbux8yAQ0LOg+vkTb5+gWYhCtyDyN1appPyUhBx
eY4WEqgFUCKlG83exxvL0fHjJ7GTzMhoaOjN5mC2ecCRmVtfp1hq0uvPimNXoDIh
/PbyxRFdiUBEATSPLjspbkneqKtnnWcIbKLeb1NuxFrgIwlQwPkMiATBfOw0fP3W
Mdqdxo4usrsjT2bphcE5knoQy1aCz4ie7Ivgh26B+Vhwh8pI1cnGrDmdGbyCEzgV
cEJ1OmLOBAh/PKOt1sKmfwOcdZf/79NgYmvijHlJJX4NhAvgpIZlPB0huxj/Vumm
FEtLZVI9+KGhdxmghCR7WRP3NqfSXpw4UovHfRmqo/0r4J81p42uIX59TOt/W2+w
cV2G1rLGI23sftS8LLIxeC+xBkP38C0SpC8UIdWmJVC01MB54kQk7krS6jkdCwBo
y/nGX3BnLf6q/k5+unT7/1NltCu8w4gKuO4unBlM06kWGLp0JDUTzh6NJyDalIH7
ZwUm5iBi9xR/N0CrQVRH6IiGrZppy7fsgerlWrMAL63YEm9Gl5oQvorvqkwzDLiH
aXPSmq+8xzTyAmBxbwotVln+S4dnjx9WgpVmL0LDtX7iqagRFuAElniTWjapdTVY
t8cvONIFY9NpX+ox9dMkCVMNGoeSsydEY8w1Xu62cUWNjuBxD0Lcym57fXOvcLan
YxLvNJFuOKDQ/pXKRDhNoOegrDiyhnsmUnxmDwdTZpVVRJFt2o0HzDaish21cDC6
Aoe6Ic8DEpJiyIiG9k9yijVOtdy1/MQTe3ATlAhjApEtVXMTTA/C3V3SoUoR8mHg
6NLCv+1mvsOQOBRKfUfHzAaaA/zmluNBhUyR9CQBpc+ZWqSj9WSqH4WPUQkdd+KF
tCSWO9Wzt7XmTLxI2nAdAFZ3mL1u3bXEZVRYueD8VIfsQv6mTCQYKaxxtSnZJgjK
L7xC7e+wQynSbIOXVcAgLKktl5dGVJbre4GSIojOcn2fniau1Ro9spTGVFPn7nqY
KylbTv5RlGHJMcv/l557QH9OFN/ASfJPExj1ga+B6yyh4pG3vVsw3sYfQwAUpPoS
5Fo295EVD+aWJqOPHYJOaU9H0MjoNIWLIJwUiHP8MjZQ1Y3mxNwG7qIQzKutM+5K
o0tuyfPQLTQo0A83TSe8cEOe7KoX17lhzcpBQ+VrTCtGBwrCdTv3EGBlLr+Mv6a0
MKkdiIKNMUAFbmbUwZmN4ZxzORsB2c0HPMeqS3TQvA88RWoa0Pig5WNb4p5WGBS5
YqkTlKYTfwsWGCjrLxh9+yjIntZlOKvng3yUU73efkDLTpa1+NiqCQhH7H5MHuc0
PXbEJNoREzw/DdmjCBH5yoBQTxSjyjztPUSfvKS0HnSeLTPhU8CDrdVu117JtEaY
5/Th2LkUq8lsViHFnJJW5n7SgkdjPOgjeoFy+JFbO4W0JFuGpbobPG9fbPeSZc0W
6NGIYcfwOaeENgLpoD/xr7+Lf/yV7folMrmB9mZJzAeiSnFm0wr+yHamtJuktR33
iPjbNaBTaJHP6122iDmMfUxYVGRsSZbvgdVcoYNi90wqHF1T6YDwnwfIPH94++pF
sPX4XHE8Hm2r9Wps8Lp8vK9ozzFyyJXg9UhZvJbZWU17UUQpLGi/FPp9MHK7qf8b
8g0GfLgHJ1iS/mhsYLYtXe/YkyBN7CCxCKFBfwbkexhrrmIt5qr/bFJWNPAUdkYy
hkovoHL+6re5UFrB8sxc6mqQz55Rki04yklKnBaCBik161AHAs/YVjMz3p/jigJk
D2LUJiQwrnPyVHLq0iwlKiAJFNLnxw7q0TH8HAJ4Y0lWfO0tR5pceNbMJOvZUzbI
8RFEBJ4ibwmQQEa5heJlxs6w460eomgbc56LSr2gK22sJsCs8Xt5kjq+gdh17vqi
gAjfriKm9b/HKFB2mZF9ew22q2O8AKXnsqEVv8/0D0c3A9KYVrgPyRsWf6XpDGw5
MmPPP1ydTt0qgk3SYvHaZtuPhRiAToLlyXBA2wR5OWMs/PbcnrYAckmYNa4wx5eh
CcFcWv+p9Xr4hKPpiCZW5ZgpQ8XNX3QOQfNtVP2W/q8zzX1p8DD0b3cCFWR/f1L8
C9yVi0IqGC+pNcIxzubt8yVfhGGh/WejQ4JcafRLWhXb5EomyFDYFPTQwcGXKYv+
O/l3vG6BjU9GCst4gucfslAbiiyeXvp4zVu3tym7J63VfnqH9RkMiAmVz0Y4PzQa
SOe1FUsEFnvOV8caOTkwWYgDi7MyiGfUVdO6SHm86f9um/gCjtVamo+hPzhbzt/X
mCihxn7LonbL4UNWC67ab96uMcgsSsAIbg7AYYA9gkrvfYj0rNFSejBT4o4SLMIc
+r6otNggzfxolGh6YqS0iY7XsWPWDUOga3F3chKoYcvGQmh3ly3cI4t9QHJKHizQ
drCiemFbo3vLOfhqkTw2TFLu+vBSH7nxsn0F9nUYow65KppDpS8Tc1ro1+uuf0wq
B/O7ufrYANfnNCduUlbJzhbxL5+nEGxOc4d7OTmkxeGJD3y34E5Tax+NKNqDS8lD
aWVVlNF5S2KceMge9vgt7DLyRK/osShSKZssu0Q9rPv8IAcSHGnXj3pA8iRV1Iep
Vt4WwuWS87m7W+3DPPXnIjSUyIoH4AeeMikqZcr12wAZh0NqBG68ewSjTyFeErZc
bienbHjCt1PsrXExSOJy+yMRJbB9r0Y6813/8fyczE/I0IQlTegAfWNMVbG3mxFG
Af6cXbOF7KSy21/oL5GxtRiSQEYeCnz9rsoaY7v5Utb5W1UZb9edLC2UrNs57NMp
EPL/0B402AtKKh+PrD90CkgrNzHuWySnH+lfiVz8XpqUZOV2RZDqDQw39ttjUqlz
RYKCAnIeH83nxdeest9AY+pjNP0gGJM29QuOeDRICij3vZQVmWCw/QvqFp5g8J+U
hjRPCxaWZ8SLRgqTX+S4ZrpLHIX3kMDjgx8Ql7KMpfSdMiFh3OsgzaZtC1Nze93q
6/HhJ2Xgsa/gJas0T4xm2cXKlFwVg4D49l9E2tcXmmqR4SChqcNeitXNgo2b7G63
ZhjmN8t5xxeHNv+62n6HZGRW0zYnfR5qLSG8GRiTAo4NmQR1uWCM7OBYTddnZam7
M69cM5oQwzM2QNmnAX0UUbGiNVkxJgREjCOrCHJ54THwSNrskM9UU/WIHohgz6gl
XV8UUZqJAwaZYA/GuWoEd66P3gdMAGd3UBuXcDn2C0qwsdLoUZ/pII8j0WxEGV/D
Moe0sHWtRlyRuPDQXaYzlbz66bDsSm4jkgkBaSt662BoZIMYxhdn0lzpaSq6ta8h
elXwRIJhF/XKBnfhEX6B6auroaRhfwRRSSv8JU+ckuclyAfJBTkhdFld8dyR4QEm
Tkm1fOxuhyG6FUHY7foZO4rYjvNaM/UfEnr786BuHaB8m/65PVffvg67g+goqSHo
z815m7WWdhnbYDqS56VRdiJjAlyLfmpPWpLj5Q/zP5fL0X9Bl+ociHcfay5StcFu
DucJX55B9ANPGxho9Kkt6U2Y+hm4FX8RKkJMfwrvSHPZI3BaAo7XuWktN4IhSXee
d9z64dbake1tEMx02h5xZ3/4jmauiZkAWPN9RXW/XUV677Zlf/WnFUHIL82JE/4P
dbSmLR7N740t1+5q93ibURurUciIrv39oIrc0pmIdAZsDgFlTJluvV7nhn/GhzvA
MryHglrY5AEPwXZdKvr8G7OZRF1Us2wG9vSSBMDeUGuc4M1PWD3ULjeptOwcYJ39
jbUVcdF9XrBlkh0Ax5lmC8R2KymZSl/oOLDCr0ycW9bRecEI2oRcbhdR9bbBwlgx
4ykTJTSGw4QMhO3dZvzOsHCrzBuXZcWr2T6PmbRFJBndefdWre8+OLiy0xFvbENA
yfht8IPdt9ggqEg1dIqzN2TZ5AIP07szs7I6SzAqNRYmjOY2c0B13NoRBmu/3gy5
0wI5HXCxZMpEEmfwE/Dr5UJoT8ezTLy5gjpnphw9t2haIEnYPsFqb6okZQWbkO9a
Mh/YrWlIdDfN6Xu+TBFfy+bEpmbbuhNnLOFKA8Ygw9iUfCWbMVssdnB/nvh7UlO1
zLupA6inO/EulEedxPcC+FeIMqByh4SqgcSOkMJRGgzY32kjBYabPmcsQobTUEKq
hfLYPlE8bYpXNCkHOgO9JgZ5KTBBm+jZoIlBYvHdmRHswwYAVBngEwwE4bSn5RAl
yCub9oYCcPdcxtzW/P92SzUjeenMzY7yqtt7rchY6YWvCSfhumnt/6UJiihz1HwU
wUguIXxdEIMuc/E/toWJfWT0znSpBlwgtdYEIK06vDKMlMgaK8irg8uSqAKp+P5o
U7EODt3/WPHx2oONQuUhdwD9IMzNt/7WgjOikHKA7r2XNW1dFEkGVXmT6GKU7qfR
ymmDTYimv0MQrEBa5YnH/wMMVjL/OFofxfln7OOll4VYYBI4cnlUfCblzDIOAxIg
rY1aLxHXAwnQPklJmAufqi6NTJvdw1SIuZ42xkRiSjTuCY56BVyoUeMk0GxfysOs
tyZfTWgZwQIvfPbBqyAxSDW0WNEHkAnUF487bVY94+yfngH+w+zCXHOp/uTP0W/f
hu2nsx+S//6XOa73weg9X0651L3O6Iwyq75bq0Y4Lferfw5PA7qrhmRF1kHSr/bw
ftJep0riUXuY5MTdJhZ7D5kkRz2Bj8171kZExum48ZUIibrA32NM7BIlksLzFR6Q
pPL+d0/22hJOTpXLE/5+kGB6pKu9TCIQIsnihnckfvrR8rt+iU8TuoHCJ5ohfMJ7
R6e4LBYWmUNFjV6FM3DiyRlPXv8nQihso4tv04i4F9wYv+6SA6oeUMbGN6GAvvqw
CdHQoV9CQfmN6hpevt/I9uG4xPSDvtedq6H/Q9KzAR2vEW9gfdrNqRsPPgbQCUmF
eE/vZZE52SyBbHwOcRubaZKXzndaqUOat/U23KLhatddW47VRtvpFhQb4eiD25bQ
F/Z3ar/LhfZs0mrIXpEwmahZ9uph+M4Xaxib2wHIZTB8IyaKZSKa2uzTOVnbPPlR
agosO1vGIJ/eeCHZTCJfc1kd/ofija4PU1x6gClNL9NHJv4kgxSRGvy1qUSQjd9p
kwswikefIN3O4c9BUh7qVgOQsgICPt5tReWntCDIxmmMINmdGUF5A/18zOUfkUa9
vS+QRQfVV4rEbumZNSBGpBeadPDWe3N8jUUgam2a/nG/kAl52bSLni1ODtAgv8+X
tynli2SBCfaJKhHlvX4312UhuoTo/+xio7PjV1bi+2SZOXs9MtlOD+OOsEUBqlrS
nOyb6IWcjLc2yWa4fOy9DvC9guTOh1//1SIhzWEBkTdP1bILQY3axabkUVlx6PrI
SmQnNI2u4FG5l3F+tqsN2twMeuC3WggtVJ6n6G3gvQVmEq1X7GX2y9UlWquYy5+g
hBDLgKyVGH8bD5iOBl78BNr3M/VKK9EKAO+N/9Hf48KfhZGLDNHuRJFUKJ/DluT/
DYzioslKLuF1kM5Jn9QMKtJMNMbjI+CVwv8OUr7OdxZiLZK7BtrC8dbjLdAJBtpE
tFbABFRXSuK2FaVgRvbDLud+a/Hl8zC0qEfizUFHDQAx/KdIQzv78zb0JpN+LY6C
XhT0YBFUb62t2BttfSyOrb5/NxCbgtgPnIPnErny7rzKo2PUQz7rJ6ocQEJbxfQc
CoSXXyFV4tY/Cz2UVzAhn3f+LYLkb7X+Ih5rOp05NVZnNQ6uR2ZPI4gH/uPHbMmC
voFamJWLG+MGmPkDfLMD0/Fns8UdhqXGWvWdaS60nKzhxE9DyiIVpXpRRDxgFUG3
69bP8Jdaikc2q8xLSHKvYLc1CxGyB8Dh5pdeYl1W2zqUAzrdKG9aPF6xM9sLm9iV
rECZD5LHY5gfmRjZmEdTt3dXn5ge8KvRdUFmhGm2SAxtku9Iv6DAk/FKpHNoNP6h
xMfujvLkppxF7IzhKkaM+9fMLjyDmFy3TGmG6eQhQVH0EQeuN7JXR9lLlzvxc+In
mlYiKAeQ3kfSY0hiAHTveSqlt+vX4s3lWOm3NYvQpkqHUb+pNrPeatT3w6nrqgoz
OWs7Bsw+6L1pEEUCdvmA9KhLgMDlqO39h+os6hPPLH0JcphHIK7rvBLTSY6V85fd
njizFDqXLUfLVFEZRZR6GdTmpGrda8wIOI/xLrpcMtI0FnLXWB8larmHzSRd6C3d
An8Vsw+I0xZQc+65khZpaVMk32oF/uUeoafeY8Wp/6W8jj8/ku2nD8MafFWCuq0o
LIerX3zLcziCBuRrxQosR9L/AixhBi7Cm9PssO1cGLDVFEvIRNT1f52z5yVN7W9O
RrmxmJE4gn2x2tP216OZSXTKwUiaGMqqH5hi6JV9Y0Tj+Q2J6LtbjF4dTJPlM/0W
bFwAH9RfWta1SNL0H/hFwl42ShqQsK06K8b4d7OfxsvRI87284PWX1nyyiYVh3l1
Yx9MtZMaP4qUKG45TnzRb/FZFOwJ7m1lwcAFhKluqNs2ZY3+YZ1fiVZFBEIzx12P
ouQ+l7mb69o2klN3XbhsyaltjQPd0qB/Um/y9h2lPFypgtM4ZJjEY/2P4GoPLWiY
JqmWQq8YcO48GhWlFCV0CCHtMKVmD2k3HkHifxM5QbhXXvbvjyZsycWob36HEoCY
Np+U5sCxStpBPBqfnRRpBsjku+O7OF5G2iAKHcYLliCLW+3Qa51HzuBEB5xxi1Ie
sXfP10B09b3KTziElHMkxoo0iNERPh0Blbuh/JvXkWi4IJcWYvFGQCFItxtES5E0
8VIU7k5yfOM3kalckeaB/+N0zx+/pCuXRJair/29obOTnijMreooB9incYOkjr2o
C1Rvg64xoLn1CuaojtZNaPGW5iAiYkYVp1yJ+MxWbow/g3f60/WBo0mHJam8Kxrx
QwRP/ppXm8uNZmiLpB//gpedjQCPvvJd0p7BgWY1u6ld+bZ3dyzz3xNlG8WjJARO
TDkwu02QN2xNzgnszwBJwLw5gWlWptkJAQ9fxU/fPm8zblZuh6iTgbDEQFh8/vTa
GHNP3RxlKYkYRoxvdzo3OcOci3tuR7ApMcZ5Hr0Og1RjgTsUN2VRHHETiVtDU2fU
Vo7bQPxwLxmMrQ/rDaw1dWiEbKhYd0941MQemrOMEq82uFcuLEdHzVrDnGkLOgW/
btvUg5QgDMkTbU7pixzmCRR2zyOR9R6m421NzwWbfh2C2335A3CvxcZ4UVIetPRS
V95xp5QJ0XhSvPsBbkcRSTHtc6xlvT9ViMgP7tavFehf9NH2HYws+OEmpp0e4Po2
iLox/aeT5B5rHZpJvN4oWkZbFIbGj6YYOv4dAv5RvT5Nl73/IdNqLjGG1Z/hQYAp
RMHx2MhCt9ZAei6FJIfDvCB3ZMl8wB49QOzF8EAn2HVhfaDUuCZD1xWNztIaPMeQ
fb3/RB2SwXqVMFWUiWEb+AbXsyMvoDHQzj+33K3/OQJJMFrLISceZDozhr3wTyCH
/IUHQNLp6c2gcQOuejONweNffG9w4X1qBdNHvs0cwJOH9eS29ZSYWR9HwWvkA0Mq
vzrI7nix1In8LYwopP7nCTOR1vBz+5o+c8kCJN7GIb5YuXVFbpwBv+qla509LzGK
dn5Lfoyv5Q4K++Qm64tjvjI6NlQzKPo6vH9qgDbAPKtwi9O9snmZhfYHuH4o6vVE
Uk9s6C9q5QgTjV6QAp9GvS1jGQs6opVALx5Qrb9Y/gKcvqhwWuuedjVDHG9I7Iou
qmNHHcUWbubSJPG5b91j7zKwSea7klVItmFi9sGSIZX+zHFnGm3KOAzUnRMJEZCf
FgdCpDZXamWDit0vtQtPRDNJwrnwowVjptg24iycpOV8BTRD+l6k0yYW+e4H0vPS
n5avoUuBwoBGqzQueoUbX5MVDmZ9OjAfJCJuT92vjmaUdV59H/pQj7mIQkNknQME
kmEqNCpi8LdGJSRL9AwE1wJY9s7mviQWvirYQCblqij8yKGcxz82MAV89mnWTMTT
Q60bhHXZEdyQffNp2kUXCn5I9s+DGWCkJXC8QOApP1/Rnnr9UdRoF/hKR2/rSSV4
cpqX960Bph2uugcEHycQyPnZvA9hhT5Fy7AOM3LPzGPLk+nQ5BmJIzt/rwU1ykkS
ezlHOxO3sI7mVGlvY6hMjY5gHx2gr93WsLP1NSVozcIf+dRVe6rHJq2BawpNBREw
MEDd7mRwD1ErxnyqCWEnabUhd+isxB1DcQOa01+y2wytrE1+kaVsvmOlcJDdXYrT
mYi60wXz0xow3uyuiN3pgJWe3/Dv3YtdCvArY7HeUI3bag1DTliRzfxTGTfdE8n5
OJwRsRl141dEOe7mvQMYMHj4jVy7DzSY8fPokGo57Mp6KQGK96PVGcRdEvHShkuP
lAIvEQIgtzY93g09YcvA1mGPvecuPDLkzkj/GG67ThItDIgggSpYE7X2dEesQIwP
wbZvR6nJ8j4p6Hf6dPmoP0dlVOSy3RRxF8CvAUiCMOYlarQlDERIgDfnfQRdYwSm
YiXtyEBlwBheWbCoWlRSOYOiZMA3/vtP7CazTAV7fSWuTjGZFSuKzvNKaeoc5wtF
hDdK+ZcEmXdAUlxQyNZEHBsuXsw3VTv5mXKk6RiJQouNkkG+XpkK4YuNhqIp70I0
ZhBEMAqnEfFFxa/DPrUjym+xgxaH/5cgy3sgd276v4/9TGiPHBgF1WvKHI/7glSd
8w34H5Q5ueWstG5PK6um+YpEpJqQSerdIJ3wONSo3VdyHEddcVmZBgzObARmDHCy
ebsrjKBNAWEEy1zSSkjWP3NsFIozl30DqyCS6GXc7fQ8Nwe2zhjgqhCI0ePZLD7+
1JByAFw0lAo9RaZfxHoGw+pFtvY5QZi2qfgW23Thk2br3574mHikda2aLyZX23Wc
gqB6Cy9r6Il9YWKo82tIgU09y5Mb12ww5qg9K57u7RwhEC83m9YqPvlMQAxMmkDO
CckHP1TWMXgoT+gH5qQQZnSge3GWyD9fL2qhnTg381wRT9Gs1ClyOKF7FI/YtdKi
SZEE8GcJYZNIx4NL8zZa/HSur0i02uQg0pxOlqA1aC63qEtzf7rtButwTGc1q58E
+qOnrpmuk4BVN3BXHNdlDGOsjiYKb2VxT7ydjmI3OIHJnmwKcnWuxn+FFlEh3WB5
8jvceYMWuSzD89f/ayGlXO9QC1Cp9+Kz3twGGN9wDnca6jexJfcymataSb5FiPbp
UeGLZObGsdWTjxI4t7k8lwR8EfHVJEU2/NqkJsXB79cHQbGUhW9vNP28/qr2rm33
N1QBPbh5cf9ODiBrHMCo8idfovpMJj0LZzRJmYb+RcbjegLKglTyseCofpO1a6ex
BPhvPEf1lOsJ9z0mMcmTagO0nRMkEAcnWwT0UL5wnlc2ydzEdtzoqFuxD/wfF12H
8Pq1WSFVczMw83l1P5iJ5ZKn0Ngpr71xU0AZ7DE5MFWaalHBE0BmlfiwDNex6Mi9
YyaogO6a9MC31gjKRaTb1tTpSORm2SDOYXApsdOlCbpw62MuUbeRaOK180K+1cdy
X39G5bNBA0yjAss7MjEUp9h3d8l3UOfvtFyYr25nuVBp/p1inB8S+qF3B3INOTEO
rZ/PAkyq3UzW7/27MdQRioyNEaWh8nhA2HxBoU7/UqAIQ3SsMev3rh5E9BODXaR5
NjFv6vt5B+rEsLOyDzY+OmO7be4d27YkfHpIgj+pbCVNqGWuYfxQcdU5KIyXi14t
rk9jhK3OPicH5JRN5AhcgKnz0D3puL/Cy14I4YVH2m5pLz+j3891CEG7DqlmaaMW
zYHLtcBNZa55hh5j9mz11d8+v8D6TOhB2C4AT4GAX9jHJGe74BQgYye1qw10bzDP
dkkgUR7zxpijORaJb2Z81gAMtU3E9bNwW4qSCVx5+eKd01GZL0rj/F2YWejMHhlG
sMd6Xqv0xKr0+0fSGE/m97ZUA/t+Jum22ZH+aB8GRapvPjLRFqIhYYYK5/0zHo9C
ifCCoI6jQBZcGhKG01xFed2eklmYFN5nShidt5l3QJ3Tk1Ldeg49YSRDaEE1tOH5
fq5026ljdrLjpW2jn1N08nSrwOet5BtoOu4I7P7LPcgUIow6TPaBuKeiSUZ1XvN/
zjjHfxCIFmgsCgsbv99M2k/nKGgUG1vkmpInUcxUCUo2+xmo5u6VtFod1lShL0+2
KK1ZpPQrNl4D4+xUFIMHz7rSHGU7b8Lv4bnCBXQCqYvfUmTYjkjLkEfzLtjdNwDQ
Makago+gbAtsFsXHWXhwZDULHxLOG8q3w58tGO9I/ZeZK33RaR4D34GwR+BPMk5n
EtXL6Z9wIepcJcpU2XW0moIfLO07aExMx7ffcrlo4dsrV3ovNHwTaN0CpY1KtFqj
d9C9+dNgumjYIV4kDWZpFGsdoddaLWyyXA2uKL3kIfuqW6Ryy/AedLtZvhg1NVZn
m5rEpBCvrkVRmhb0dhA0WG2ufhrIERzKW+l0RSt+Oiruo9oCpgxSQgLeZCFUrt28
DVeDAwttVabI2SbxogJNZYCU49FeyLZM7zpRgvXy7XJncsZtyG4UGlulfCSl/bMp
M8liEdlPYxNlZDY1uqMstkPHR7JI1VECXtSfjSJ4XTwKFivBkDKbdXpc7snhuMmT
ir00HzL5bJMd9qY8QRZ/nfFLhkW0oU6b81K7RXNlXPGeXXgW1YsHb1vm4Xru9byE
cPBdRJX1MUeyR30T6K4nrshv7PNWOlhw0dZYbj0hYM/HPu2xek1kS3R/mscC2ucR
3xBnITq5fZ/bynRxrvkTTeTvqER+smRxQVey4VPZG19NcZTYG40AOshH3BTuGArU
rruAE+KMmojFadNZ1IfT+t3CQ0G3YQaRUf+cGYpVT3ogh+aUESeQ6MXLo0/5Jkl2
uyTx3WLy++rNGDVU2BZWpC51eB2zt0HcDFdcdszEbCFRzHssUrDo9Gt3L3Mj+YOa
FudZbTC3GmPU6RvCQhwdf7OtJ31Th/FzzGxIT373CgFax0mRFI3DimxHZZFwNYYW
3zz05J2pd5qe2jg8L4IxLLhg/YM72Jpty3CoSC8bs+b0O+BtEplzTbN5TfI5Jbuy
yqWxaqp8r2ZOMLicmP6Jk7mpoYM4vPy28hpw9Hhx1v5vnPzxU9kNP8OvqvvS6Uok
79d9PKpZIstapW7qC1OXQt+iGgPHoAZxolu8lglK6NYNjE8+FAYVlOfHauzTB+eU
1b/NnhEjgTg6ew6gGK1q5eo+s9jiVzp5MYKc4YFH3pJq8tL7T9m31yH+CvKNuTip
8kN4jqy8e8HC8hwxl8gsGRvfZzlbERikw3wK+6wSsi2w8720xNAHIOCQ2SIFgOEO
G5pS8kktzEYTv1Lsj83ho7CiTKbWwwHYWTcM3DY3qPZY146UZ4jyiF7WACIwX92I
+pIYvQqg13poQaGtzwFSOlMNScR4ST98xZXXflUbS0yrvcith449a/auCG5nJ7Gg
PJ42+CfF+GZnraBDfLz55nM5h1gQ3VMaym0jdLW1nKS4RxHZUBcEaI/yPiyurVEj
KiMb/Z+FOCMmgOgcenvb6WeqdNk0pTz9dSmrTkYT9dOpsJ+M1KSLH2hnCHRQ+AhN
B+79SoL1ZdfEC0h8sCQMpOfB0wRYQLuCIDlJ+FbaOmwpO0zdTAAXnUA+oRL29oqV
xP1fPUhLbKq9IDLA6CsehcmeBgyxs5pzUrSQH9v9asY22DiQhhFfAI5PulctAgXq
DVxdowlQIFbKSdoi/42D28YA5og5NcY7R0ojfeLsuzmIC1b5g9/LBHIS8ojTl9uy
TAL7/SwbREK0zdLW9geQe3YchRQhvCiDxZRrwsvOY6YTRdRxRScLysGUwBEv3j4p
KvrEwELRngUAB47FNuqB/AjE7/oCLm7h+vOZ1j9DSGH0N10IY/rRMFgVLNF9FJP/
K1NBxC6KX0X9ZsCoLHVL5VyhV1X2Ge8Zc6gKdxJgvyp5iZkWjeUhw6N9f4Y8LTh5
X6GdF5CzrBapDO80oin3UZnJbTlzc6RV6n9NwyV8w0iCRUCRpXpz6+ngNWWeKQ3G
cO/co5x7IxeMHtTLJkgBWQUrB+54L/XZlG8zhiUU9jOgXwWnfIngDJQk5sPSZLNl
69arcTT8/MGe9DgZud6TCCyCPdt/SRosPW1cqZVJdlVQ9QuWF+hAm/HR45CTkEZP
2gQh7YLHtyCw4tI9H3WA6E8TFV5BmY2uP6fTc8NaPiqTuZVmOCphq48SQkERyKBs
OHMHiAnGzTS1ERF2xOTPT5hA6hngAkJEC/PI/n7txxmYSPnnkjAJtXjsjqDHZler
eLrnViN3uyPPtHVWVquY8xXRuzSsh+CjOKN6B+Qe1HPl/HjfG9pjBsb1PQr/WYxS
R9e9+qMLCg4k3/zVRoSkJ1Tw98+7f/NxwhqoRMgYexHYO8b9LuijCw5O7lg6UU/m
AA1lINEAFu1ZrMSLo1Sveg==
`pragma protect end_protected
