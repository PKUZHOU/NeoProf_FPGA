// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Q6ahNwnHKuMdzIv4fXS3W0Tqe1LjjDgbfoZObOFY+IiwUPfPZCQsZ1RloZc5
czoJ7mDFCZz+yBQhb/TZRaeqL7VUlk3/ij9lfUUeV2gir8p3yJD/j+etDjnH
gUca+Yw1QK7foC7+qbsi7kVHMKUzrNmWjd0iTLBRejKFombHeQTdh9MbKEYB
VvA0pU9ZD0mKE1IXz++lBSOeOOmREEYEr5qNvDDM2GWDAFZjVnKJ/T2Y7BlN
BJqVoMYOiHCqFCcu8ZzoRomeW0z3or/aATdyW3pNqcnX/l3+TkGpSF7e/4O5
a4vgr+LzyZw1zSbvDfLDbxPKR1ImAhlQD55On+JWBQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
AJ0bv9GbsU+9B2ubeE91Pl/x0r3eEuu0YEncgZWKU/L1of4gfzRi3USaxAFo
zVOa4nxtsFn4Ovo84OFAWI6hHwlT2SnuUQqeQ1QXnDkNw366UpF64Zfvloks
W0p6JIHDwruCSMapKev4TDm6U6mV1ZaG6eTuEZLxf4RDYcO0zyOK7NBKvZHN
R9mF+hoDaxgptlchFrn3aerrlLiNl341d4m7Jylj5Usx8c+Wo2gU1+PkEXd3
bPZBADCsh++lDUSIqntjyyx1XQCLDjTznaPcJPwqG9atgnkzhTcwjXwqxFIV
OetFQW4lbI40bkeoDQq0baLECtB6e+bRO6qPVKJRtQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
jS++pdznZZHaEof2tMleaOpDsPiOhgLpJe8BD2XHFlLf7l/5Ay6wH8AwOVEz
pIH2q5gt8FripmqeMdlWlPENCeR97rgvhim+QB24cJn8AlQJY5mt9cXThpSz
XxLw9StlW87I9DErICLbUSud1aCz3wTkZ0NGN/9+tBEPH4oKDrmsXjHNObib
TxRBu57qVFUL/cK3TUWQfJ6TIoPuGIYIJ6HfDWVPUQQLbdDiIfD+hfCcwNMy
D9URRcFka8GQbmaQIcGekkq48cIiGyyPM2Tr+Ky4zbSiyC/3CyxowwHG/33c
46thvwli29lw+Kn6gVtBnE9+288fMIEwWn6dxkwrQA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
PLLdiBbg5/il3L7o2Js5I3YhqDmFYsPOELWlCUb5/mAnTdCMNmbUBaQuZoYy
ch1HAh2tOHPVOonDDKW8m66MCTl3/aDut2nlFTvdrretp6MhLh2Ig8g4vp/2
pZHlFB3BXhWuzmjYX1Rfova5tTzXg1zAcWxuT2dur8S3lPQnehU=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
u1lZ+Xdihy/7hMt3aOwQttVtXg8PTQPqXRO415LirOwOtNjlFF9xbkVRwo+X
LGlJnQBTwKtSy9gAv3bUbd15NHtpkyCegPgQcArKu8qnm768jhTrXjIh1j4w
8ri9Gd6iCWVnxa9Azsp8QNgB2BEtgMFpUTg1MbSqt9RY+bilWw4LGmNfjEfL
nFOb/JvtelqQWyYdjTZXpfh2ix5oh/Wd8v9A5ET2FfDHKRAjxEwTAh2Vav6m
4BYiSER5hkoSE/dDLTp2+2ThrMgZj2TnVjOOSkWB5QNB2OQUCEjwn0pfw9u7
wgTfkSq50imH5a8jxdQl2+yPVhD6YeBkHBFDRiJHvJohWDacW9oGAB3Mwn52
HXckWBYzOqdbk16uy5wWn4lT4a61oBR/GLZPaF+ZkspjtzAW3qhLknlc3ROA
EHtH5r+pODvF+DO8a9fWNmrS3LtT674NS4T2iI+1AMtqy4X+Nii57XZRDjxT
RjjeSmryHSS9EpsXNm2aY796t/QNIMN5


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
pkJ6uVrVZoixWIwnF8M37BHGKL3eYZz3960wW2zD7iEpW83cjlpSUopXkEZ4
h1HLoafIs52b0zS2DrdtNHeyQ3Z4ZhKFqHkaZuslQZHxZmCrZ2VsCK4dQM+D
JhHieOYi6/6vEhBMJQckihHqG9DKgC0kQDUxD+FZFGKXWLICDFI=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
CA5z3h+qsDXmkPCQDzJ/5Eot1MSVaRR0D+1qofh8LVMvKYQqJoOY/GMaBNnB
txv7H5rlAkuNXbby3jgR7sxzd3lyE6BLwvux7ziutq+mOtg1V+rN8PMS86AY
m8IHyubRUIKWqCahtp6CkPcdXHNhAgy0xEnj6EKnpnPe2g70z2A=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 421024)
`pragma protect data_block
tkB8GRyu/gs4SSAojNjp5vHA8lO7nmgDrjWYeiqTC54aT5LUkQlWavUqFFg+
tywKCxdBHP7p1FVbyRB7h2MXgcVw7tj7nZyvISkzc0pk7skXUtMeTWL/PW22
fauOYc8ycpdv2fgtdfgWpQxMrDD9bgl6+ob6EX8CUilbDhNkZ4PUGrhM3Lny
Vu8eMNaxXSF2GtGsemCaoNep7e3Y4s0j5QrSreBm4YI+quwZpBA72uh1a6MV
RP5IwgDguznSmYwppKtjYo1RhP1L3MypufeEFVI6MpqUS9h8l+KkiWuOwhnY
7TEHjoh4cZr/5iSXF0RJoYT6AwvJT74G240EAU45mWBB522PpztoZDiwAoNG
7x6O6erptc2y2rOZ+NozKuK1sqfCDAFxRWhww4xxXQIHumRsUTePF9VKMIzD
QZM+FIrI7iLI7VXZcNcKt+YulKfelIe7Q+8j/HweZcQU2n3/1p3FTGDO+NWW
eiY42V44n1P6lgCdqcj9S0I4+wJpx6Zxw7FmaPdxrf5x+c2LBokNGbaubShO
Esum5sFHdAosINFLCoyfM60KeJmQMROz/BMVw5jnpsifK2fJkXUnco2GkHPm
VxIKlcjqi3JOPp0K125FX56wu3NcrvHYnoe/SQ/9mL4kNh1FR1VdA0kyN0wY
hQzNd1LHiK5zSm0f47JcYo5RQ8NXpQOwg97vy5uIE0ibQLmASVxpO9/Ew/DF
sOU95aWUlsCHjxAyGZOY6/cCnjludrVKk+wpr6jHN/OLGg+YsRWXXQHfXytY
8nD3qZ4MrM4XQ/uSS11ouu0znCeIswjBakgGnxIYqBnI74S41AQIAHkryPsy
tSJLIikq5Ea0n53sfBEjDxIULPadrEIPbIwRiS9BXRgZfEOSV89bzOsrxQd8
avg5oU9zRGwdrImxP/TmGsXaNj601rykQZBkGM1nGB+JASdhXZtMDbYibFCo
LZgXx+tA6ixysAw8fXs5NDbsxkLFntSwODTy5ZkgUWu9ZuR47Us2cI1W7/g+
HUp3wd12+wqjLJBbyorLPmY5HMtne4M10PT8YJgjenf8fzDACxw+cFmRlNaH
NkhLEXakDgFQALTzb2l1oqgnneEgBKRjD3Y7Np0yUAekTSl+/QiHdYfytr6D
cxECRzMsLKt9NbXBRDSdlsO2u6u3NwMtOr0+Nj3PtsCwd29HM/P4gf2MDpTj
4ikg0yEtEez+WvoO+6l5eMYemDgVC9dHCTtrnF9n4BsM0qcDErQddN9LzzgS
ppwgI6bwfHWERFnCSI80LtxxSjpelgWgMPPA5jHnubDqI56DICaBxmrsBoba
1QI81SOsEbzgK4ll7/pmgP5/wcBHlLvWo0BjYn6pyPklHouY3zCiH5SqYC8+
U8dR2EEjo4ACLmV/ux/FsU3yFJObk83Vlis2tJd+sAtsDUz8qJ/uYBX91K7K
8TaMk5fyKW7cA3wcBsAGSGnzYAmNgoUXgA+3XmedDPw6+PnEzuku0AD5Msra
XpHh10KolGTq4oTrqfWFyO0+juziH2PxPWBtK+wjr61wvVp4cYcDe7g3L7P9
nMr37DmpS8HyDr3hd8xNLLS1Nt39ZX+ducd8gM4g7Oa8Xcs3QNF+gKQx9Eqv
nZ/3xNqb92O8jD5DfwFjltamvF1QTLUnTcIYPHxSyzzFYLEncmrIxMJgPeQS
CZj7Zj4FNX2VreYIgWOb5QMyuQ7g24rXXo+UMTjJgQcUYQtAtI1DbaDcmwP7
qLM0XJssq73nc/g3/7LblsGNfWLw0Ld3QF+m/u3PYIwLq/JrI0y5xC+1eRy8
aoJhjiE6WcGUcE10GesSukxwj7WgsWzb8UevylYqyaeRW157B5lzAV/aqLzO
hWq5kigWzFPurD/cjFe6ZQSu7+wtPYtQjUXtRPB7saoiwA5btZIpwt3ezfqH
YheUo2lH3UJrUgqj0QR+S/jdrY2vH4oynaHLVVEFsTiQqQ0UcZW5SMkUNyOS
TmvPrTXps5+ZNZ8uCdXizX6hHPKwlRLDm9MyeWUsQv3R+Rr8/UgWAtjB4pfd
GanGXv0YCFmjXvNwyAssm80lt7A8qB+vYvX4M4CO6fJWUB2GnCO8aoIEfbZG
exwyWCW32PET0XbCU8NHovxix4gsnghRkRQ/nERYsLSFPxPra/H0WewoNcXB
61zL6QztMN08TnmrDq2Z+beh+ZQ3uFzwVs/HtZ2PlacPi8EkvOrEllywbjR8
zkuB93Xi7OUw3npR5Dtwc14ejEwp+mwLK1gZfgahlWoWpR2OX7Ojo1qYn3Ib
th1JcuKscH9IScbz/h88HRGWqiOXQQwg1Vwmmq6QCyGSt6qVV4SDk+RzECmc
hbObPqcmfvPjJ2o6v2UOUztX4kIsqxXnnX6ycG9w3ppjvPQcsvLCceua+OKO
cfmGX4WeSgF1UdhwZkTvZ9cp07GWcYDZBMCNV0NgjAJUOq32jGrDCeNieUZb
z1rxtgb22Wok28ZX8XKSOJB50XKFVoE8n9LSJlRJvUXZiWCrmX9WuykxJSBv
qyOBbDjSU2bvUbwo1fFiC1YguCmbN9xELoUpi6x03tedg6SqlNQr8C6lmPcN
NGkemVYOnEsjZ0vG7YUyHJSf8XhKPMkpcMHdVstG6GBezrXi7HNMiq5p/fbD
R+DWI9ht4xym3m2dCEbDNo5yYGsJWs2md1fLJtzF2g2Q1fca//qJamJ/gEYL
Rj34E4n6j54sTl2HdRAQnpSm1lqq+uFwZLFdjQ3fJnBA2K10poPCcpbNbZSC
nNeTQFO/C98WExIRdVLEgq0DGDBKdPuhmf1O5gog8EzNrMam4ROtRuTUPNdj
K7r+NNe1rSQKEiZi53TLj7TC5ChVjBgLxVtoR/72kZ/QlETuvzhhf1WuzgCC
arXQ9rVvRZ4VbOR0jh6Joo08iGRgM3qoiYp0KEkeu5P+cQK3yJU8wFitD5U+
L8cgJ5NUbTTXiwbC31AdhVxz9x3f3ZJLOf1yy0MkC/2jtd12zgHADLsDrwYw
AjQnRTif9Mtr5Tbh4FSQqXna+EPhFTi0TMEWtYGpw0wtx5RnZupeerRfyTVJ
wdLu1Sia8/3FREmMqEhXE2FflqtUEhj7+tk4Dux1E7zWXGB1+3hb6zqLoE0U
gFZafa1bhdfLhZeVxcPIpLWZR+ARbUhmaWLCPVYEYAXZVlycl+NzBAhIxqDN
kMHQwj/JBYRNFHCR64TzKXNNRDg/aSJ7qBTPIZHRiHYO51a7YJF09QedZXAi
NUw6BBSHl0mHxpnmOB3BEBy4rBrfYMO/qPBgMQ1RNCU5VAOYTUZL4qvTQVPt
aXPvDwOV22VvksNcZVjz6y/lv0bI7msCiVo7olezxdi3uhlze1Du9GGlVyln
XWxiGyMslJvGpejyMM89Z+n8WWStQmnznaLiaHuj9oGO33eBTKVe/Kv3V3Zf
VnTCgDod2YfM6hYuOiUr5dFPZxj4ktB4oyi+7WRhtCxEOSYVr2Zr3qa9Pb2g
+sZNMcYIguVrpp/QFMvTiC56O3tem+ajJJU5rgHpG62gg+IGS6JUeG5sSoTA
0PKt/VmvGVSDy41mwIwa/vwEXlmbu5YcfPoFEsYhTuiE/RooYBe6Ozuom/iA
Ec7C/Zsmm/hluaeNVwNqFkiO3GuZOzklRQWaOupeW31vsEzP9Dn0lbrbH2mS
EJRXGQBCkQYH2/SCzZTfGZazgbm/VEv/pKv+bwBzjMbOtafKzubEdtwAHFWi
+F5n0qzxP9JakcI6OdGhaOM6d+35eHiSl1BUfrHgqpGnMJ6TtkbQe5+1Q1LT
jPjnMhFyd+x/u9xBiNY8SFi0NuI46YM5VMX5MHim42nWqGH1+kY7889QJTxG
kYhDljWP2G1F2IuCAE/hLZ+T5KD1c4pC44ijrq5mCx8Yp/2axhdHxucuo7CY
F7ofh3bnkpmOKQlsf/D+RVpojuVOcLoLYRqLP91QZQrSKyf6ycH+Al9uKIgq
41t3GxC8zlb8BZn6Ie1C2VTUAURYU88mnsYsNGQ0ku/Q4d2AQLVDxElDhP4p
3TCHOq+gD6zUHSbKCpNXnNKz9VpYnDP5HlbDaIqj0SULM15/ME+O8Cg+5A3m
R++JGXpCP/ID8CG5NqzhsTE94X7vsrm6vVLjgjneKCX/tugV9lY7jX5aFB86
KmefI+khyJtCAyyIz/Af2zF/imFfbcCkAEkm+QVrwjX73GG9tYNwn1Q0QP5q
5wTZKswIszLDdSzal4uOVZuW0FIVI7DB5AukVNzVp3fvJWw8oVfDRPPCQ75R
pfWAHd6rMvXtukEs2XRzCqE6vtJmobpFBKtPAPAJD2xS2HWtnJmAVAV9Q+J/
y0Tayh7xZ/+E8Ike+iT7FBqSu4mLUgCD/9mc/BBLwKgRjNQNIbrjsPJ3Hrq3
+Mv0/d6RJEQgDLIxZFlW1AARjGH5E4U8ZgBuJp/U1xdYTV9wSk8LuEqg6wPZ
/hMcekZpdMOTCentwtmE/2QSs3jKDKScs8OmzDkhlAKvzOaxCLjb/b82WctJ
TLgipqFhX9RgMbT7lXVluh/kgL26OKv/I0BMCkeVGzz7NLfx+ioCN01Ma8hQ
LOINGxwCavqy5lrd8eyaimT85gemsiCnG5b8SO93REVGHsrZ5fvjb4qumXY2
uqbl7SPuaNTWDSI3ifJksJxzwYd0O6XpNzSzLXPbD5LWCNZVd02HNzwhBVb5
0HjOl2BSZUC6ZTcaivCeDIGNxBsUFM2hc0Zm5fIby3On1W+X55UhxhGKQlyd
lY/V9MohN4JEX7miV2qjZwF6cpX1dx3ZgfrEkiUpeRCD2KXD7qI1uQLAHlaB
HodbJK5LQlr9994w4rrhznmQ44S7hzw5TrcSIyh/wCXUvHL8lZh63d6Ab8Ij
hOEkAvN/xJV/QX6u29S6vY200q5Mp+YjjZRtTZ+s1aCEFIrQYuXel85BB5hR
lPLHLiy8jJk7vEL83SoLre6YnimtmJmQTWKz+Stj1ewnyfhv1kp9kdPK8sfk
4c/qC+r+leBndGSd73aIBPqTVOdmPCuRO7oOzaA/G3r8NIxZNUTSbQhz5Azg
uAHz7fpWBhfdZrOI4kqMsOsPQarz70q+nXZ9RqmmqfXvBP2as5/5jsomx3EN
7uUmCHk64aEnXm4pmicCAOdySG4abPSYRwZJciRp65uhAnj3nhTRCa8LziXC
ViK+1m24/YnKlZGRXRDn9ys8QeAKxLJA86u4nGYNENyhqi2Wmc1KXGGIsx4u
XqMzl6rlPkof6lPNOj2bIM2AOQxXen4r1j785UimO/OEwk2YZNB1nlYSFIWw
JIp2rSZLo/0D6yf/nrlcGcq9In7HAwe2eb/DTRDEOcYz7li2W9bSLr/4NGSd
K8BntdMYAYvw6tHHMbgjOClWnQahgllMkDdMKRvN0zrVvnizFvMsa3cAlulk
NMyGbfqDBt9WvKN6/ta0MCCCx6dZlrzlRRhZuub1pjpt4RucBbQ4jETL167j
zgsxmeriB9c/wuSdIdAVmgjRj41Lkog8fQeLjbE0pOg3r8S/9bZVTCYd5kxi
/I0sGO6jWscClDCl9a2r04nWfAWG/32zoZOCmDmQVd6Gaz7294WDFmTez3no
5+e7gSjq7hhBkKgRri6oz1td/RxnkSdnrCVbZliiozOlo+h/J8VwwbBP6rvz
6VeNzzlLzSGR5PgC95f4JLNIlcG+zX9WsGasaolnFb1eZTNoLCvUSKisylh3
MVBCv0fw3/BLhxRFLvyW6lMBZmbGxJZwhgQAYyqoA7J2iwx92HIPaqQJQVTr
/vnZ6OfUyhrGyJZt8CrnSbd62s7e7DGnrzIREJNMRIbz2S5gldO4XPFk/x24
Vqz/hQs85dX5sFAZCjSHvRHXKjL//2R6Bk8FNjwsziVfvW9+JDXXqZ8ilyYd
SzX3kAeB642ZD4yuGDhfZ3gtlwb13HjR/Sa7ulK8PaKgZO1BHP/lf6el2WhI
Mp34Ioze2o/ACJr8L7uxcCujy5CYE67E6vRk2jQmwTl4yZKAstJDmevuiCi4
FVUO1YMuPsSo3NwYa7VoiCH5qL543oF6rVOjCj3zhwkJWW+CLGaUiYAXHAPk
ZNtDjGmlwrYQEvaysUoJPNjVl2lmSYuTXbw5ZIKGmiBaVEsuVrOuKnEUeBas
PGEVZa3VcEj4B9B6D6qTzzLth/7oKShaIh5MLvfUGL7PJc7hEpu5C73zoZ8W
8Sm6qDkeTH0HVN91h/zDfWhqjt5AdymfZtvsGs8+AEUOlt9OB3tCjheLpaWk
LO4wXgOdlDpLI5o53J+AYQcRwqKyjYooYpGniAw9XIDuHDCtSBiNpQMw9Ndc
NC716pgsmcnabKg7Iybn1bRUHq6SdwVEj4e7ioqjvpx2/LSmOkIGykps/6qB
7V2wJ7ENeS+pQGaBF/mViM3TYs9BFvTJzEcMfCLACpMiIvmQeeKpSH29ya1R
vQcVZWTw3TTN01MTm+K4jYUPsfqgpa/jmyFXCUfgDplX30I2w44Xis/w7On8
sG8QaiZaSU6gMQ3Zj1liHA+dItsivQb5k69T2sVfXfU5+haLB62VexdS6uM/
g37VTYj7LJ5/sc8tg5WxFXmiCZE5GBAZmykRhqpc0J94n3lSRiX7USavQH7H
jtntr9c6X5O59WSHE+RarcYyHxthFPTJV8vl3l9BG745Y6bgvhFE1WuFDprn
hG7MTjwiVcwlIPTbQOl1+h1UtqVom3mSprLW4DkJOjoaU971p9aKjt9oNmz8
0V64cbX7DBmSK5/e3hBh3Lg3WZ7VmA5J1J3MUp7RZgBCOr7rC5Vi1wd9ia4Z
MxPUtjYD+D7n91sV7Vjwy0QGgxUSEIki++EKecEQcCSKng+Py7dP+e/mTaQC
6otNqumC0zFAI0FyngRtiIRnh1dufXj2SJkx4UVbAW1flLGtVS3CjYB4mm8j
iWud6YnU+4tEr3CFEyoAqNQuoD7ATTRTQVmIje6GY1027IhbILrHfVIikJJt
fxT0QHG8J2xG3XrY1Wk+ZsmZy760Rm8bcb3yP13cO5lqFYr05SifLPVNyKZu
9G4uGt1/sxrKKPbH6qyONmqldNhhPUuPijuzcQdZo6FHIUEk3wsDw5HxA3Vn
QN+8NBi98pX9a8Z+JITDDpG4YwbPXTdPdLmxlCUNLrgZvgUMjTZGNyBMffaa
pjdKnHScHDFc7f4lnk1I6fDEmqxmedllg9panpF7dFCLtsMy2bPhHgJVYA+U
JXyaVR7hmhI1vqlz7IPVQnFjz1d4gLmbfg4z8sJGFvBhsJD8GFXkqamkWXNt
zWSTzMIkqduMXZmeH6/jcdwV4yk0wxk/6ZknOh6nvgxHqC1wXBq6EaZao146
LqwBlHPV77YdNYVWXPZuLx1TU1OOJM5EUyKH0ZqIQ1f6M5gr20kLcRckwbtk
MP3bJvWnnxAs9NDeRvkyXT+kZw5PEdJiMHgQV86IVhZkNrjs8Fuqq5gb9OU+
aWUvrLkAxU2Cxlu1GZggWltZO1VV5XRi82ktkE9ofu/RC66twxQk1yHRJNzf
7t/42NccWL/FafRl5+QiTi3RZyOibUnxYA9q+o4LDBlIhjgGFWbnydihdG1A
w6DbhNhoBwvcqxpucgBuYG0XiXJOhfAEPmxO9kiFQWcv88wK4zPOZfDYtEik
tzgwtzsbkagWpITHPbbYtzSPtCuFclEBv2IKSpGv5Pk3avfH8DlLAWHYCEpX
lqo0YQiK0n+cmrLj509uQT4mVoSnwCtaHf8bDp6q4krqMikG1NLw+pCGYtq9
LD1vFbDI2aLWfG67W2WlXG22AJr14ZGp3vylSdslK2XufaNUPGgMfgpkGAKb
nVQGxGud8RGpi1xzXmJNjMFoG4ODG55dFL3Oe+9ZDSrMsWwcndeM3yE4mLHE
emsuGmcV8WEvNWI3nBfOtVbVdeiSOiYG2irxUJ72CdmghU05WNZGkP+Lbbiv
9WMOEcnK+KJDnu676c1Wzqa1r74GOG2yIv7mt5uFiSEcq1zWQnvBHD/VmTl5
Rz/rzpZwJOLiL+DOEczeSprS+orlciHtEy+0j3cFJuTOWbcOopnSKekgbO3k
0mJa8quHxqstxQL0rngdcWcXJDTAaxwAP/ETnNr2sTyLjwkd8q+BGIqVHvyH
Md6qOsf7SAg9F08NiuWA33EQ8l3G3CxqZ2h0SCcWg2ItCXpyaKYDzuNg7G33
zimXJaAMHQmMEFlKVd2QOBQJhjqPdDUyVa5FCzr3PNcQNyMEnk28XKSNdIns
NbnjFOuYUvmKeOjaVe9oB9nP7io0Jaf+8DAqoHSas38WnBuYSYwNbaIp6t3F
g8GKYO0kgNdy2f+PvkC0WMr55oj9eHTWhEmFRNYV32138bvnawTOTW2mxHIe
Kz47UawtgIAY79TzzupCEFzkxS0j45p8dVw4t4fLECL1KRI8PxPiYRkRJ5iV
II22IXAvMsKOwj6YnS75oRqIYh1Kg0xMjCHaOc5g/4QisCmlQn2lJJc5fUDB
g5kNpTJQM3B8VptKREC6RBMjdAKiCu7+yVYIio71+OfD4DEKLzg7W0GadeIn
Ey35NcuVs4ArtIT+HwR9jZ7djRqf39peVuek6iLEWiS6s4I9jwWnikIzkNOe
4D0W32fhLDaIUj77JgIrXM9HuZUYS9VB7Y52WJntdTQGlwuu2KF2o/l9YaA5
93ic0As8zbv22HAGLUhADVaync7Jk7EFGKftMja3+JVq5QZIRUERSpHJ8Qy4
fRga5bpVPUAB570CYcmzfqb2zEeeIqQTgwllXepD/ENLmMcv/1ama4GhSNbZ
BwL8ULLv77d71xRea4U6XMnHnB+IQGuxj/iTEoJ49J/wfCeY3KHSSLCzS+qc
gD6yYCUOlp9gWEzJD7JUV+4Hhp24yb2pS2jbq7aDS2VrEJmYS/bhTOe6ADwA
SauzJVW3JnU4etWTnqFJAlKiUXe2wpOcS304oxN3xc0lTw3MUHn6x+h9s1c8
xr/xgVt8XX6q041O+OzYmmkRYRJ4H22iCh8DFxw/SIZa6iD6J+qJkcw5sDcG
99Sg5QN4/hoVWlFSKciQAcE5tG3fQGA1kDNsxwU5ZX7ezdmjHsScTFGh9YFp
C6oXMn7b+7d4PAET/OsFSxHEOpIwJc5CsLCrYM+xdtMwZx7IAKocuIwRQjSD
P+sZLiU/eZbSp+hfQ2fP0E2bl3vkP7LolilkZY1RQ6Rfxn1Xv7MN324LXDh+
6Bl0eVoX+Qtie/L+hj3P11LldJWzAH1FFlwoeaqsNCyjEuGGBMVjavNpnnZ1
v/Cto+c3KYkTgTxU9YPIuiys73YOX2t+o98o/fJ0F6O774kTIXGudLtggZep
JtA0tRSEdBa4dycT0hIWPivmrvpZXQNHZCoC3DVzuwGnehw6bHQs6XOBVx9v
YSvAd1ai2VC6RWNsaRaJk720hyqc35A/ls3g83QgyIZApNCybO7ojZCqhFgy
+EoV6h4qsmZn7Gni+HO9+XdhyGvzwoHcy5jwB+pxaMRzywyUjUTxVJ6zXBhT
5SjcIAx0eMzfeDlQpyhCc7SPmUpT6AxLjx4EiYe3UB8T9xe+QLmVUN9uArtp
Egunf2/Rz1neBXBuRPzwY/q8RiGsyUEFuudltx2FnRJQaOo3pFBT0vBAiYBA
5cTzyGw9il5X5mbtnoxYWvsvXgURDnFyuBCHQqLyVnWi6pl0t7bEb00dNcMK
gHUMLgr1HWqeKXcZFrLAAhuMUvx7/0ApCa4tvyLqtT6+o96B5xoQzUV6Tmch
HNbnMkyrBrhkWCKpljGzeathuCloqGH767QI5BSW5x0wiWGm2iY+I5ElJjN0
Hu80wmTS0L9NcUpKi/CC4ewtPTAmwcMz2DpPh3IfK64ZIo5lTb9o0alwvYTD
aETeUQZFLym+pfKuyL4RcN2p5QISTgUVjj/z4gYjNJdBbXTSDiXCVOuBMvO3
iF+nqonxcWxPukWjH4mpMQ7w7hmIdd1A2sBxS4Or5tJREwSng40XgrQ/89aX
5V+7Y1ExTWT2B/6gM0DaL/WdHbuo7UoAq9Rd/nQe8N/mg01f9283I57foA+/
vl7a0cEPypUVTMJfBZZefjBH81mVAdSlXLy/ZpfsV3aNrRfeKCSYwRu8B3KD
BQCPscyxMCupoIaCU9Q3iyAmtPs0Cq5NPOlMfGlUCzO96QvYKDOl1ChU3Qnk
2I4N68upq7bhTfk9LOol4taghlqXTWwlSM7Zz3X1G8anuPgk9FTX3g5xNHJU
Z/k9JzAp8Ne2s0z7wJgMDWJVffQsXr8qz3Q68mosGwKsMMyKnYL8nQkU0+Ya
bMf/rypxZPEhNnm7c1HK1HBJNtjVsXYtsnqn94ysfMxBCf88fIdIYy6p/5ik
E+qKCTwPrRf9MP8+qXe6V2atM0sPRTJJcjGVechk7dEF2Nknq4KqiQ+4cOMi
CUp/lw8mJVuWjOEGFQdFdhQ+rzu3soh9qhpTNfRaTQ0gVutDTxspQ9rJCcho
CyywE6GeLfZjtap9xf3t0hqOSK9KwMgiiViqnKGPK0mrnrfMiW+CO4XXiBg6
h+42sRwEUCQMQ7lf6mNNM2Y5TQcW79pthR5UoA3xAIxdwFBlr1u3W1rD8Uyj
aRXCGitj9jnEIZJpM18o4QnsOg/zQop5bHEYDi9NQ6RFNVD5RnBjAehzUk1F
I9XCfgmGLytAD5t9GYRv2PEeIO+vViIHKVuhnot4FP1GtZfgI/yl8IbwfZrX
A5wSUDcUsb2AkEknexEO5zaUScNh0ZWs4pOCNKDg1QfTmCUAc/CMsSwxAUcK
PdIsE+U1WHuqbtoPEEoIMKifFpo/pBy4U3WuMCZd/VQ7W+8hQqhkJq5wODvP
1+PqudRPUJlHmybn1AuF9lFb2ay8eczhsyrhd2DUDTakTLEYbVLfWqzRIx8i
koRz4GRQ0SdOAHt9QejcQeGDIeXQEFr+xhBvZtwE7NpdqzCanpUCImxks3V6
kKVr+aqVD2IbgnQoajwfXiWuqNSBrFs0qogbLMK9UiqfoZCK7en7YaKyQnwY
q799AxLKfVpBx9U0p0pYUM/9caRKwKR4564uMsJWuPWNzII+dJ7AG2/se0Yx
9uCfWFqkh3GCAFilrQDipDwhwnbY8R/d81AqBNDBPv2WblLEBAX310nnq71/
b98mJD6utI91FdOxrq72V1bHaF74McdzOoGcKIvpaOb57jLNKDg4fzde9zgS
oVLoZYu0op1zmsbG86fkLa+oZa8V4WV7fqNkQhKoPZ/pbji5frxbVkgQvbpE
dcA6je8OGWGlYRAt0SXwsZo9XwqKSHBEY485S/zSl8Tk03tTc3COziDPTi4u
5mG8dDlNXbCaiGmy5YTgIhVqrApnXi6PkjDSLTqSOYkJ1Sb0an147vzSeanf
bIZrs6IDK8ozxpYmXbxmnpRuFWtyauWugQQB7436WiUfRC099LT4kQUZJ/UC
0bxt4TR8VDbwdAdunVDHUyPDaknyjCYS1d/SLuWWzid3a4iyO5xXkrFuZpGV
+Slf4x/yiW92yoqgSG+6znrC77bxrSCeML2KBmSuXn7l/25IMbwvCYULAnNb
jNfJ2tgvFCD5qDzeBcm/qVnmSxJiFDGOPggtx4nCfLNS//SfHIf1qT4pLC3F
PXY3R18yNP1pk33ok5IYce+hUNRFWq51RvFevcasltYLwzbNY0MRwL98j0cH
7s/uvRlhhSfJaCtDlh8tutJ5NvdyAQ69AXFKNChxySeYlPj471io2QQufx/i
9gAhlKr2gGCqW2nPaWhLcY01AhlSaCaQDjggD4DkGboCU9AxYvGYwxuehV1v
1Tg4xKv7UQuzq78YE1ZQr+Vnu/8itMQbWA1voXgVf4QglahQwBGQ3OHdK5Ts
pTLzF8QEiko6B37KXk7fyDYL9X03OKXLdSKaiZ5ehlHaxPmPWwyMGd7yqBqf
S4oXYr+gtXd2r8T9pxSVQIVxFBfKatxLVd/UiOn97iBsCNDe2L2Bv5ipOJn4
TjhaURynstWCGRpk4kqC5pbBiIe1XjhSC2O3XVuCkqETff/cuzVX/AeobCTe
U50+L3uz9dKrbJq5BeVbKXofTaOQJBtqKJrX35DH2SYgcU1/8T46z4eF8q19
wKFiRxiY7z5codv09wWSB20svxty/OZ/2T45CZSNmIubaCgVCH9xvGsZNypU
YiFb0L6fVK4qhVO+DATriwUa+O1wcje2XHM9UsbNbmtOC239dCXHulrqYlbA
H5h/mBegiR4EZR1GvsLN1X1u9r6a9FTQ63tAfMqQFY3NEizDhgGnSF07OXOB
hPMQhza9BLMPiPVG4za6/q1QJS69Sga8hUJYLPRdzxlTZVHTjXhCR98nAYC8
qpIK9nSISC0WZGWu/jOQnNpWtGPuLmWNnCVgyjNYPNnWk9lQ6IvcslXfEpRQ
wU7/eiiSec1FnKjvwggiXo2xqT1DASDxMLB7WpdTh1ieHM4D9uxLNgCXk3a6
6EL6XGiaeES/uDx1ZG/VG4jmnO/q31ld+aS6r2f2WeztZUsJ5pZhQqm9N2kZ
8GLRrMeNnZSNr/rAC6wqB9PTUN2dm7Zg6M3zgrS0ITEBeW6Jq1kLVOOBwzHF
uMpHz9BcdC+yaj2GLQcSOFv06Z7nj27AtkVyRO680HrMc9gorokI5eglEo+e
GL9BH79Wc3s0RrM3TAfOnHCahnlFiwaDi5g/IsKJBQnq+ElfYfeer5MGPKFS
ebCzyJ38cyZ0kQU9OtH9HQuJ5+KBBHJow963Wee1BPyqm67uRGzP0r/cuNwV
n3xCg7tANcHSJZDm994G+tDj7E94n1huZUPykIqi01O5xVnRnDbwT4LMrR5V
v2gC+Y0z19qS8pQ0NEm6BdqjcN/HN2pZ4FARzSGef+Flog3EGZmFlEnYrytr
yHohwDVwJrGnU008spnLHsB/YbU7euDXGI+kno2USYF/e5Jc6Pa6ftIebAOS
3g9uvcxnC8OFk/os1UkL0z7QnHfWG5RNdMaL0hra2EcvTSr35e75gU42B69+
fHgvXjdr0o+NE8x4TrFIYULNhxAopdnPIZ5h+jjq5/Ef8fve6cu4nwRhiVE9
GADwZC/v5qx8mJkx8FfGQwaskcKV6F8kqY+uBct1hQltEdByelrc84AZ74yn
agsrtZRQF3FN4eeMvO/MWprqBKp75o/H9lAEXzxh4HCwhPkcU6Phz8EC9+Pz
eBGxitgdnqgKJRzQIKc6FH1+5A2JTEkGnnAwJMHzX+nR+gIQq/fegdhglrKH
j3g2UeTeVYkeWZ/XmDkQJL1E2OlLIz5EuFSWlpzyDr3oKTWKvaKxysa2fygr
WxjX1t6KFzH5jSI5Fhi0KSgi1qUv+OHw0D4KS4hz+DCuF7JxnT0GhE6apwEg
vhkuA17Jx6WH+sIdVpS/YQ2X+GbH/0lr6uqEiNuIpzWgnO6oT7EB01kmvdPL
DmXJZQHIBnd15qcrz9IIrCMd7E/TnPJYcAasHKTtzP6yd3uW8cEBaSgGYZgZ
qFrAKHATQbGyOOukjttx++TPr2SIUVUoLgJSzR0loUC5tDlfsd9VxdfaIrTf
sK7AwFdCZipU8gvvrfezSdzoMyzXBUMy9RKPiqTl3rVTM6q3nLGZGPlZbyxk
PP4kTbRx4Ll8F40SSD1uCVg/5WyYyhr/0GmkxhZveWwxQZXFgzC5TErJvDUM
/HowdSYgeQwwVjzMRxDsXd7V8oLPYO9CZzvM6gEG0IiJYftA9ykCSR5XYcE3
36kesVe7D7a4JTW2yOIUc5sSOL5Oocz6E7dlazT7YkB44/oOJ3t+4mLExfgB
4B5iv0NVUXbuaDUM52CexCs2IwzHvJCoZmLSoCONMHVN2IoqjXGY8jSzM7ri
8JDEcZcdXbfEM/81eXYnp8QEbatjZ99MDrypA6uJE6xEzzcL+SQzIeh2u+Iv
jRqdUhihF+IsVNG5qJxPVcqxyC/kKxsgRrtk3Ve3tLIOYK8b5deOUS5sxO5c
k5FnpZ396fhBPGDspEJb1vhYgTSGxG43jpZp+kGSgHHA8keuMcoTVmFmtm+E
77YpgQvkRS8bZl6bZXT23wr15RChHAWem1TQjY5IeQB4HkLMOHRXxQPPYAab
cuxK0dNGoAhPdvkWors4tdS7lEr2YADP7x8ip0aRoutcF1/n3uY7D5378iKK
JO31yAKpYgK1Jdg0ncIDiwMv+XcF0JtBMseW6fSnqnqw2N6tt5315Lhfz8ih
ME78n79KxQlBryehj+ExU4iZFVM9Fcn+rwLTv5lWrsIZ6TdyXGIcb168LN/i
6HqPtdDeY9eppN0ujh+H7wtVOAkiTul5hER4Dq6LPwkM8CxItsUCYL9a4ktM
A1IM5SHUXv5wviJaxlUDzTyl18Uk3h+SGZewXOmH6Zgc7DB8Sn6kN4rn5BeB
49CtUSG38hiF7WbbN4mBuB8SQ7L9HO44cbxC00m+HgTgragnqOjtPFfYpuPP
Y+T8b2LkMaYlPskf65oQvR7I4nu1C946N9AmBSOaiKFs9H93XNNKtM/Q4+LD
+P68cpEkSVZv82/HkINz2erTcJUoGVfyhneGh0pnQlH1BO49kAOxm4XYii+m
0deQ+3XTQEAwS8erSJ1/T/tDf4uSGPp32fsQWZmRGgvpRYcO3Oz79LiN/ITF
+D919/HSDZsnb2X3eqmN4Png+0tq9LEFPT75gwHXELmoyGSkJcqSUZ0frsuY
37q4LjcjTeEZqHVRtZHZolLvAlRcay70DxOQIdDZTINZkT8Lf9+5741AqHYT
clnDuM+hvuK7M8TfX6ukRSHEAUvVZ75GouDQjBhLHNgQ4gKa02is7Ont9eRt
zqT1Xiwzqv1MJ0cI07aCBrSS2AkxcfSirOVTdGzuEi5od9NpOjEbeyziqJIx
2ZrwukUfRSnlUjSfqSTSo3RfsO9ehKg1dxFahL8d3dr6rfWAucfEjZjheLIx
HTKgffldBR0AbZrchhqZu03uNM+cslhSgBFMoH2PHusROU0WN8fla27ajfGD
jHooJXO/wA0MsYZPseCzkmV2LxWnKQ/3FExnJS9UG47zq5xiGDksall2rcNh
9mYTzEn43xpqVRlCTsTRROAhrdxfmEF8307/rJ4mTRR6n1Zh0PwaEXSuxYQ0
p0gX3NRIEj8OMC7Xs3X0YDosx9IkNToN1QCKODouuPSr+HVXtDiZ0AEzafQL
UvbkSGCxu0s/mtPsU3eE/ZV1RzOnVSAukP5mN27J20LlOy/QwgNWbtgsvMHm
9q8JGImLlBKuZ7bKp+0LI5GbzGYB/3e7NIC341tcdaQf0GOQWysTAq6RwR1Y
joBttP+w8XLUQM04ELK7L/CpMr7/gAIPudyB5XPNot0WKKL4vaH7f/zw3z2A
2jX7qOmRL5mQFLPA5RdShgfP1Xe4tP5gfFNJfnnl3Az1IFRP0xZd2O+tUSx/
XLbJSBFzuZVQpX/C3nQRvVfwq8aA5a78SAlPWCYAoH7DBLvTYqGp+9xYv/RQ
DbC+lxEzGQldAO5sO2fOET/gHLh8ch00/hFYD1ZutwMnk+CyNgjNLLNKyyOX
rxXeAWmEpbd3Vvs8DBKVvisK2ZZERIxnkpYkAn9nZhJzgCc8EyWcLKVCCU3H
owk+rapeiDsyaxqgOBThSVEGAUVN6lQnzI+cXh6Fb8qaBTxBN5H6RCZAJmXl
cvOayzSp3xsixACWGa9kr5qD9PR9Tt7ymgxwWKXVoITlHZOv04ADWWC3mEQ7
zR9Mdopi20dC568NMmRsPGYm/Qwy1J2575Zo3bUyxXpQsrcmcOI/WEWIz7a9
P6xtgUJ77tyi8WKSRgPOS4Tbvn2wEkngq+7ABwOOVBiBYZPDuLhF1FHuCecJ
gibTZk43yU9olGguJq/o4GizYD/JqG3ZREoPBRsu/D78KMhMr0LZLq0L4j4C
SVh26sTnTPn8auSrY57lQVsUyPNw4MeJfB1SKbFg9dF74iZVSvTdzb/rVt4v
46MlTw5xj1PKqlkfFuxcIGggTbzyGUhO4Shxr72vUiie7QWkHYWk3kyRxIZ7
/Nc3fSjNnH09hzv0lKzQ6tSjGQQnieH1JKYqol4Y4o3g6fbNa65WWpETYxsK
G8wOQ55Sd4y8a5lVxdGWkuo+JE9jb2umBCMSIcbrbtWPaqJitMpyE47lNrpQ
1MwU+4MWYKCRTaKhN+eWbwBWjWZnu2PDxgBZVj6obUqS5SkaB0d58scGuaHy
VTPaSn5duyMsCubvt9xzCdclKpJ/VW9FYRu/4WoXUtpKX8XQJ+ely1FOoj53
W5lhQxRcGHY3sv+o9RGTksjCVlN3eJkpo88CK5u6Z7IiMR/WcOS3+w1QfHVG
LuiavblZlqJrJ81oPpRko895bnhfUtTLXT+4f4H5mMJY6aKZKLLqR4sF6Gid
xmoHBmVPQ+c+fL+cDse7oUwfsWDYkmetHzGc3bU5eoNr9NQw2YbBvA1vEtyB
N0x8quwEtu6gfeqVXivpl3orwIGlxkhZmzPs75oT8woBmiN+SWAdtu3TlD5D
uVEZr9Jr31dLT13omVNtC9U5P4tjpqAcQqzN9wWPFhuCuHSnoWfGAwc1Gw9v
8N3qieN6GTM7POmNi0+7n1mvquDvXtRVk/Tpw+0DhHB00dNDVVUCINJUzz7s
Yp5CUcxEiQlrZMRYgx9OJ5T9CYEriCmVnhIb888/tEbR40GvcKVA/N9xFV+3
52UGNrgq9SfZqi8tytLYxPA8Vx+5FF9r/Zh7NIHijalOirew5e/d2xvO+buG
xAIbQmDGLK34KbkaIqAk4SONgwPEFfF5Fvs1IYQ0zpjbvnDUEpQJDZmQ9mV/
WmpcKf7UzDHzJcC7ly7couVmvDygmtbUuDCwagGxiEc/XgM1UUehME81o5f0
BZmkSe3E42P0fggQEKVCVJ1f+L6eVlyU8ojsGpAq07oZ6rC8XdJC14h2rSmn
2corI6FeuyJEwF4o2n7KD2m/8VTJ4PqdMy0kKg0MYxEAwOFgxuqGWKq++i8M
og6HRUScECPTSg/GccgT6djEwLWGZo7xc/tDW7kPTJehraOBVm+v3x8pg+8Y
3lntWNEghBSp+CGNgts+g+y3ITl9L1HPFFoNqgeJgyewuCdf62H/mfm5iCmt
JwVs3SkKHcIqEb8EJLijWMQNtoNjqhLq0RLdYC6gQE+EGV5cH+TBOpunicNx
hiNvIlMbvEoekDauzRAqHoaaXxCkihZwT3MFe2rvfkGmss9S0/v7iuU6fm1U
8erEXilcSH4azPvQ2TbUaQ8cP2n9uxlTTPSwmTGVALu5MhMtDc3S3jHN6zf+
IaR6JOHZqcswFMMXIid4JivrcSERPelIEy3EVBBIWyf8x16dUywbN7grvFYP
YuDCLG//k6HrLf/sgP68YjOaoPEriYXZ+CoKgLGe+21pRfzv9nDplQdfYsYq
NgvZrevK8SfdNUwgOtmMHojFGgHQyAIaeO1Nm+WlJ3qrfVrGcpoSe/pNu5tX
ez9rzZdCasIXkoP3cJ+2K7OhB8VaezZeaDuMqIEWCaEThyyNlmiiHch8v5/P
QXYms7RhjbUVpV3mKmLAwd7ESoAGjyxT1nbNXfvGMe5RdT71Q9+VQoNK1BdA
4+rE3EMcRgnubPZk+SCM4jJFpXKmj3cJeVpsAGkPU5KnauKvFAfoGnugu+ZG
GSLEry25kDERbKxzbdtFV5lBsBahnMxNXd0xk2KfQKoUT6fqQgrKnfuPLk+i
VPH2a7w/q+7ewRVFm40eEqwsk8GilvSIj4vTSk3GMDHz0VJePKxiIy4u6BWR
7qg5t1yflksgB7AurpAs3HrufYJB8SoL6R6V3uTMk/fUmM1DQFFwxMZaVIMm
G0YLuASnSNYKx+yw7T/3Z5cUotZPHs8BOuz9V1v7Ib0Wm1hp8Abi8vRwmQ4E
yuGM6TTeZwBbpze3wem/i/F8JZa5a4iJDG7NFLEyU4QJgAN9anD8Sf55BW9V
hmHjXz4dDubzHpLO/12W5vMVksq+uc52KLVovYpv20L3HbMhkwYHoqSEuWe6
bEUQwdgs1tQ7WTqL8ehJrQhC4AT538Oqhn8v0+EgyWM5gDssZkZ5t7G/OpWW
CMHxzA9S/qrLUoSUHP5v8xLfhqsGUc/Cjdy+4QwHLdwO0nLuAwHhkJCis1tL
1FNKSoprw1jm3gHfHHnowf48hPJnYgkoV7AaSruOdbk/MLAvNj6Xynkrt7k5
0epM3qpS+45Tw1clg0TwTEopfwN2LO1nqJEdHNkN0JHMbIH4oTG1ktXHVzbv
3o+7LSWYUlXi+yUfjiGeHXgUUBf5iZhyPVrcSc3F9sWWIC93NCL02djNqJHc
RSmSMGh5OmOoeS4sTPQiaRjedBS2RF72KyccZ5xi5P4pknnzjvRGuKFitosW
zSBeGcoHniPA+QWAdtVatJySuiAKsTPsWyn/PF6OvPekCcg7TkD1jqYygviV
x5CWfcoX6uq+syE8ZzLiPg7PrSGbOOp/PbJYr+PWF1rQuLKJtCIPzXQC+2dd
fJ3ydVsWotzHJpmaKS92lDuIrliocCXwvVdIT85nB+6ERd12VdMOe0832xMp
Cpqt29RrLgiOg3005ZqM1kfq5VMOMlaTQdJfWUbVen2WDKoH8/jokjKtKETZ
yQq01/maZY3skhP/FtOcHNFQymkflaCWCGMpddDeuqEEqkhVESWssPAarLQ8
4XsCpEEkC4YlgUyqVqWPnlScG6G6MOlcU3PmJPxe/3uWb2HZt1AC/wgnmx1B
ZxH+GtSshlxuFx2DOH2oAdLLjFNoK5Vs3wFm33thD7dDAGmRkFsCxlXf04pB
/Na7JyjPt8nOKQKxzubM6HjiwMXeYif6qNcKsyx0lVNNI775zKjWRrYN2cph
+41yGw6hurC5Idt1W7z8a5QbTS3UQynnsVGZ9GX1FpLhUK95MPhUZt4rF4C9
Y7SGt+PDaWyDvZ1ujYGLTE7fjGMyDscmYlWTGSeH1ar+3TI6TvjU74tvZ79H
hx/ErNkfgQpFBEwBMCAu9nxHt7HDBDJiHOvCOUyjrg+3Bd7bfXvv0PTe4q80
N8dggIElnT4dOlqQHRGzpik+oOpYXPJ8VIGdruVhK80bYWN53A1N0Zk/PFPh
RYjCeBNUYWkMOD8cjcJJT8JftPle7S/+o4y9nFALjUMgd+oU2JaTBeF89upu
TEbBcvuvBeVhlIgDKugM2DJlK2ZhU6xie/HqWj4TOqqhaSMHIpJeA2o0TN9D
zG/d6k5bY8KOEPrDzhDrcFJET2t0ay8Ho/BNb1Qzz5oBOSBKMuFUK/rToy/Z
l/nLfC+FOKqw4muBXav9vMOBkqlNIEqAkty678s33Z7Hn1AsRtoKISXqQkO0
VnHBBtfdO4XDs7GRnuAzOWiUDyFCWrCNZCu/YCS/+492dceoA8J/j+Xmrilo
ZTdjVT1G00sf4bwOpc/bTmE/Lkd2SKctbZLHKGurLroZQJd0NOTScL15arGz
UfTSltSDckNFfJxwKrFaOujxWcnDIGHDder1pWOHTlRDCwU9l4Ag9w7klhKB
6yHKybnYACjXy9kWuakCCliWpdkredvmPE24Lhv9rbIFewA5sDPD0t3bSvK9
b4I8xDM4cYzjZGUOQZJoyNMBbu6tcU/DnFXXpPUi0TooSTmYy/T+ZhDslMSh
OhZDtZIWzKs+fEq8t0MTc3jbEAEiR3jrEDuLGrk8v6YArKxFujQNmsJ0xg27
ruK0MmEDfePNmIc0D2q73FGFscjFXpNnOaf8ay0RXkYhrhildgFnq7fekP6Y
zOSdPFi/laLmtVfA98yJxW5yOaNJkMAzQU7DFFKvq54y/BpjyoCROq6CXhPR
IlueoKiW3mN+AxyeAltnrJSeQbCzs+Ike4/WpdPtEzB2kTxc6JaMVl06Vx8Q
FqZRbFAH2y2EDTqAlb/fFDGi0AUFfTVb3aqTr0c1NJeR9gDXX0cDw6m3eH6n
yi+ObnYUqT/mzPNc4jaKclTOm/sR2VlPd/UMrFQuYtkdFGvIIOXBJNOtTdXu
fONMS4BdUKeVzI52xrAJ46LH+3xd1gmR33Dv3r9MQWDzIljhpI7A0s6q7vf8
WvzeNi8wnyee8BY+zqEWfsPPrBO/G2I+n7yBFA7hCXK/glNyauf8HrRl56Pb
XVuilvlY2pQUX7e+JHoFWGtU9V35qjemk3ieoQIOTuCk+m20XighoguSlyIQ
Inu16H4YA87OZV7fMX9XQN7v4y2yjLedL7xj+ayLhlTQK+AhDeVa+QjfIYpr
yNvkwJ/MBCS2Z750UH52jS8rhEaWvn7iskh9oIHMZi8EyfDogUjrfuGF8/v1
drN+MxGQEWhK+/VQ7uyB+oI3ANlzLUoqIrIG01FEIUwCL1fouTwyXwrK3qX6
J7rEgs4L2o86ADyCNhlf7F2NgcBUnh1jvN3DvKuZDIG9r/SN0pwbQQNLwiM4
2bOeoO6m9lggJACAiIQlZy0YdK+tWgbzPJ4hwxXOdAw8XJWSej3UcWNSFKEm
fMlPApa3K3hxWPpA4gMcIAbB3meE+cY4SgQt3KoUneJzX2N1WWWFrBP+q/Hz
FJmXCdL0x59KezIT+hmhsVutIQ/FtnfeD3tSUrSs0t51v8KilFxP3/tKQg6Y
hBAheEx5VtMaXD2pk60NjS4eW8zF6rRSrngwwXCY0bPk8q9os2rRDD1yn0uY
/fPI7/jrnsQ2PR0J7lAXc6n/X1PsFILYAO0+kPX9L1qHIeawaXw4hdgQqj7g
4sAYvJuO3UfivbvHFgevB6bZjmkEO8M8vU0waUNO63J38R+QgJddiX4nPeF9
+gcCRV91CWoYg2xRMTFaXkWhlsTeau+ZyWlKt8kvMVAnzuqXGiVJoJuIx3/E
T5SZhNK2b38c/afgRhAOd3Bw8j5JUpWD2ARyMgVjqukLy8XN/GtSXN3TBo4d
E/vOmRev9IiGtOT8SS4aIqKE6ohGk4EoBzcRbZ7uQzfrQ4a+Z3+6ouhQVypa
o/EUaVcCmFlf7xmlBxbqMlFShQLHdCx/FBfDrKUbMhVzbK4H6GhD0ANPou1y
2jPhAe64b4OTfoQjlvugEFD9xMBJXJtwstFE32X7vzkwSMrWi6PfAajKPL0x
/c6mIbC40KgNIvmIoBYW2m5Iaw3dTYPLOOhQ8S2AALPBdIABIP0df1CnL5X6
gmHYkYg4gvoq4F0kYDO4V43U1a2gYswkBLPL5EIdwOUXeazjIkn01dCfwLFs
rK5a0XeUWhfqxzeFpwjzuddSoGp53gbBvVdjWWa6GwVoi6MoVp697RxBa0B+
VeXWLfvpxyAxwwiNdD/V8u0Wjfrh9UUM5CxSkhvlePIxHZxLkASuk9DveP6g
lti2177n80ps+rAuxXoGxaODSsLInEvaO4J31kjo0XcL/jB9XBzOgAk/NEDa
nOaa2ajejJIQX94/edmBJMDqesRV7GfD7xOU422ORz5uPIHCxsHeYfCalcdN
1qkjvWZ5sKXAfuRPCU4iH0dMcjl6d8ubrBMNdpzjmljOv2K+GQGNbvx6+sak
/xQb2J5UAtmCIWRIp5TlNqNkG+lkBT1/AMXggV+srFRPfxLz+ioV2+3L2Ldp
SnCf/3qiUUwCc1qbYrxNO+CKRgsNlOZGZ7UQdMWJx05+6OZBr5RkoCfnMGUY
ffxT3MQKdKo6MrH5Epc8GqotOYd0Tlylcl0kAH+Bjeqk/2lg+RxNNJ/Q42gZ
PlZEUOSTONWr18djJ+BsbPG2WH/bKnvUlG41vea/3L0ksiWlAV/WQmBMzpNY
f7Xa1nUsk4VfbDPF20iJTdkDIsObgmuX7J3hfzGeUCugapuVhZrl4m3s+nFh
lrhnXEMpEllC6IKolLTQJwZuWmX041BfIo/C08TEaOEWsFX3Yc9MSIhhAeU3
Pj6uaeiJMjINoI5khYqHmyt6b/wulFLJGDLnkFa7BfbkgoIvwQSvCVVJvZRo
mCyyI/0sTq+VQosQmr6d3UZrJw18p7457EXaLXFenL0VlIVVq6L2jMDbCM6v
n2HVRifvokDW9XXbw9Z6rzilCTDwpQxZo6L8/iMwutGmdldwT2zcK2UJ7FMz
0BAXM20sxHOz6fk4gL+XzHM9zdB0Gl3ZyD81sMgT/Fs7ZqY/HfG5As5mqcKq
HmzAKwXvi9JiDigqpkOVTwawpavQ5jhBZusxPu7Vq/4omEOC0fTxx/5+/f6T
d1F3r7NFqIjiCp0fkwbSVirUINAZEld4ryBHe9WSHJr6uErF3n9EuFBrOEdA
PbbTUG16Vs63b+TCXOFlgxPWPZ7sHwojm4n4DLbTtGRjE8FtOAgoCkIMTWgx
HY8Iw069JP5EJOGnArSJ6xH0WxpNwjJ/UOTTYejPCsUwA+octB0ASdewKHdt
7CrFhzgE/i4v9RGioafJrngjTnUeAhxBUtw8e4tKDcODsgYMN0xhhc+CY1Am
oQ+Zkpn66gzVeR/47YvtdQaqQKnY8lBaf8q0uytbHavuGBZJfnZLE5C5172U
9A8BZ98FcgGcbaB2HQbvJig/5qCDLGZM35vd91AcGvmrRfHnXlHEa/xpCfY6
4nnHeA2d2oNExI95cE7z9xnMOu6DDjIfTmSVjI1OK6M2hs68WJkt7udz+/OD
hXZqi6b93BLqV80uBpidVeTa+KY/UkyX+V5HjQeVTV0HaHDZgFMMeZiM2s5K
r+qnZzsIILdYiOFuWYmN7Wqu80SPi+Nv20tsmy5MXU7++sXWmb1frTS6p0Z3
bwS2dOVPxfokUtbh8Gw3rTW5elzP3OI0eSaz9hyetF1dPbqOf1kf1bYgbPYX
G2y+TMVm7vjTnHNd8yEAeAS6r/8BTk06SQdwzDivsFFDD1zJmO6RgCa+7OMQ
JkrR4xMQzL9wdE0/tsZAF2Uem0+YLT2sBnBzQCX7kVGbNN4QZ8ynGfljEeBn
mlopAwCJ4F48Hkq2wFCP7XJ/0dE20LkLSnWG526ml4UoSRwXHv8GqGAIarVc
9Tq7KUlPJ9pUgtDWc6cZKs2WL3k1WWQ3FYau++UeoOgA7rif5QsNapaHmBx8
NTZAKlyH08oZkV8IFg+S8Kos3NunFl41cgzdVqYEaA2AtnG1RtUXVb+94WsA
niRiJJGFZNebZJTKEeSQ7fX4cIzJEZ+0U3nslxR+n2NofxfL0tgLsXJ0zj87
RrR98rPT4vN/vDbWmLxhNijHUOzGmI02o0Mq69+20jDVknAxcUrWyfl0e1WK
3hyw7tLoylmbUstBGA+DMNIhBXo6TtVFg2nZaIhsH0LdBsOJQsqKAAXMN4B0
Qo7exKRwWxw9JN1h+BnJCdQaApTAsMqi1KGrghg3B1CFMgcQ9s0KB/peKkF/
fVRiqFuZKg+q5flDBUW6vaelWfXlKkcUCJFryuch1NKvzl/DRYNY+l8eJogq
YuNZfvVwhCdLpD5YTROA++NIqOt/ayBGT0i9wZY3yKt84I6rtvrdtNpET3BZ
MB3uyTNvKo1Kq3fInhwu0lL6sAVDoLkGYXsdeBPNajgS4lD3RI2Rqg7yV6r+
BnnCUHP5dGkMGBs/+4QVFvo9nSm66Jq8WA8mfTZ4jqgF2U9keZ392bfkmPQK
ss98uWi0c1Y/2n3elPxIUTAcCKnhDmvf9oIt4+V+wpkpnj6RTWQ0hxBCaTbD
uAWpvxqZfqO02UZums8TFy8LB4EqPAiKpUBzs5LpFjqTUpIeLDNnj4ZK7KxY
H5o9t2gKC1NSKdHbi9HJFRwHJuuZ2upW/8JqYIjzcnYdzZMiHtf5Y/7DMwHs
huNtW6/lsusfz18NcY9Q2LrRFSjoH9qCp2ysvOQbl+iKjVbiMWg/MFKe+Xfa
o1Q+Xbd5K3PV/ToN7mCTq40RuWNqvzQGHTaqQY9RM3DKDOZE/O6wmGSyApGS
B2bOmUEPtzcAeDIfXvlMpOMQ6tRmobrGRbRZSfxDWgzRQ00LHE88w/Ni34xY
s/8QyDEzZ+I/gtqXdumwv95ja68Qhw+NEifIoi9iFUK1LgSOjCTJCGfJ83yB
kJvhRN1iYFDcSg3TvfB+tJG6dCT/9Wrh2y81Zni+C3GsAFRjSaW3v30Kt9cl
ZBptt7vXfH7o8mrixCAZ2krKJEpj0wUSlk3nZ4Zodt+r27i259CxXYn+2svV
IRZxuVsmeDAY0wzuPPkj1QmeTr4+9vs762CxvqKOsY9+wjbX5Y3GDIsAPLLf
hsN/t3wKtWvZ3zp6bxjCpq9kEpx17Ou+xnEWfmc1BPKhMA6H0MJV3kSFJCgk
bPM4ctnXzTWg5PqdPCHdTU6ZBmWluRW6ZBhEPJjb+319CLMDLEq8FJSfsZJJ
v2pyOb+BcIDtxuErcQeLxNVtEQYwwjmscXKftCYcypXivzyziWfzPyXcG7jI
bdXdYEWUGeQwdSkLWLUnpD2pM4pmj27p6HhRBMQxvlRAJARmqdzLEScRu3fh
bvsBMZTOfs1ZuuQc2dy5Ruw0LyUgRY3Pq+3OIkENQnsy1lLZh9OnS0xgIxm9
7ubC3IGuzBA5mH6gYTgXB4rQZZ09wtqm5OzOsbsr/uw38pV4sCs200IJKP1I
rKbzIicRGV6XvZGOzR8xUOZ6rbjj2Koibu6Rr2kugsbFTRCctTRcKCKv2NUO
osrmu4FqwqdisiDrevAlj1erPG+812Wft5I9bVt8IPkRet6fHv+2Gaj4aljM
6jLQ959MPGCJm1dlzNiibe1sduNlWPkG5AME7hkXitfhF0AxoZIJkTg4j5Dy
RVp6LvQhBEHE2zqpEpfMlybphL2X/HV4tL29hmsPX03dbPvO99++8V+LqyIy
xJ5aj2j8lk9mYLm6uCeKe/sq1bHVk4XG3fUeYck0gJCfr46m6VkKuIEiwHPT
dbxcjXOFSnZvVZLwMnfVnC+KrSbIRf+E1hyCV57IslAndl3DUMsHYVgavgjm
HQGaM4XcPTLMzv1gzFoXbPm2Jz5mhwpwftjOxYGhgUSc/HOXSbkqWzwLqfi4
ns8AjoRUCRbT75lsUM8hkI8nwR0pPVhE8Ems80Xp7LXVyhuWtdyxBuXtG04s
jHGZxLDqL0OiLxnX2IicH+2ljkQVBvX+5arp0fsfuGGLpxpIE8Dn8FVXTfyW
BborrfV6o1T+fZhgiTxmfixVUeWwEUoi/JBfrielNFt3iz9baGlUGdiYFzZf
4RNmjRWpqeHvAU3oFP9DdexCgHGEknBJNg/VqcnCkSU4x+eXmloZYja4U+Kl
bEnbNYkb3K0LifsNC044+lzIjeAl3vTuUZv+ca7s1i+kirXNOi+F3XfanuNi
dXDGtHC0KBE3ZrT4MeaGPnOFUIpMNd7EmzGhkV4uz6lbrOxQ6dvwxlaMAtFy
a5fifCjVurzA1OXZyM1HllSYrmVriKgwGIDDgSkh7JuuDc3eJ9sYqDwQ1+WN
/ic6dnBUmQobY458uvsa6bS7/XgnbbEFxWfEhezLhJoowDKBUSd3w/4NBRvf
BFOJGAkqtgkFH171ZZiSQDrZHHL8+nctgkRJ/FjxwDRTeBr05SCRcqO2ntad
eCBoIW+qv9JMokyZaS1lTEaDKwgGAvFmbFWR2Qw2y8v4wpKE/wIcXVrxkvGP
6hB6Yk2OWb4pRPmHZSxi7Tenz6jlQZpAILinwYlKYbsodb7oJLJ9eNHawtFG
rTBjtXksI4lKBjRJsyhnTL2oNLTgTaiytKhcRVT+4ygMtN1PpM8wqK42MGqa
N1iBPA0/yAf7hu2gjsJg9kgcEg5PBc3cHr7Nl3I/uuJFXxz5xc8UgidocUWI
LqM622UsmvA6laFIYSt31b1Ehg9e2C6saOhplKaNJ5X3/CWQH8pypcvY9/uI
eJDDYgakTQ4pYN3b0pKsaqC+VmKsoE3sMBFjFAse8NWNK75K9gAtULvWW0/q
0XNpoCLgpLj3rrFN2FazpG2ehO0EGIcPX7E/DS8Y2Aqx2rm7guQbwFgYq8/W
45jnDLlWGrfG1S5QgLlrWkYB/sVzg0aM+5SMvM7Ot6F1Fx4U0hVfPODK0FAs
4Gm5E2W7ecPrC/q2yh/+t2b+6KcZQuQPw6UilIs2VfIKbEtKYBuniyZUtl25
RnqxolpN/eJxzPuFfghd65j2TfQo9PMRwJLDeSk/J088xtl3K0GaICrxtY5S
v3Ebo8QsdTjxpA/7/XZrSrVUWehWlFfnuROjv6XTZVcgTUTYipiELP59dn5i
eWb1Egw3LTQpDJTUbZcO5L71/ONOKl3NgDLyFrpaoKTwcMdxPUo2OCONb4V6
kGPsizOdySCS0MuvhQni1z6bxbdc1brMmyud3eN1CQp4KdAI9/hl3zEZtWsS
jg4JHPZv1tauGWlcwf+sqDgaqbIcJi6DG6xn5JjS6LG8mGhfd8OWbYyGYS/Y
O8SQWrNE/qNj4+cS5BzRqCFYz8OZtMD8/YtYhix0j+nNVDh11RnLlu71TuAb
vxPfK20ydt0XU+CsAarC2fJNDF/2B9akfs3MQe9L0Xj9NX1IjqtzTgEZ7j65
0CV43+N8jTqS/923jlPQj50HU1BX7DftRVsmnrJZaB9C00URgixR15LTHjPG
EqsBJKFfj1rCy5RIEwIXWccOE2WfzARPvucQcIDx8j2g5OkCZtT6gvi7x66b
8cUJOKRLOfskMtCGkb8T5EK83424NJFeNr9V+Xa9mAkXzEm00MLpGMYIueYY
57eLOIINlsELng4z6WX+rKCIHCOADLd0KAWjzSfPqWiWNihZYSQGpjyvL8i8
S/zfWjnMQRhThh0Kp4vS9MwnQL0z4rC2RFkI4ZuLfNqXKd6xqarX8fKq88kc
Icq/qVZQUHGzNl3HJBw8R2Y1keEjuTWkJAyZy20rnl5SIpGBExh9UsdHLlWo
zKPtli/I8Ts7PpWZPSUScMD97aXzdTT7rc+o4/e4nX920sYzwdE1wsXjtvPF
qMNJPDCswlLR/xLtf/g9yADpD5FwZI4xPOFEya5NIAq5pXzONEMAY87A4EOM
hkhHceX5ahaSoZRCkOEvYSBNRbXJKcoUxzqC3EZ1bdjYbGng0U5wCy6EmwMP
F2ufFFyflPMLSvB1fE8FH55X8OVzlFR8UN10rPWpKUPJWigqpvaRWEG0Ut6a
vGCT0PwJ1+HWqu1F/j0bsaFJCeugDJ6lxBlp6dbMsrH9NEDrae2ga5kuT04b
6xgCknH6TPnDeNBfgpI9XvSOZAKKTB0fCLJC131S2hQAjUNJcgJVpoJgYDmc
3tkWzzhUNJ1JhLsfsCuhXR0SSn4wHty8UK8Jl8MCv2JaDSc1mqReGmlZicyn
wiG+2aSac1Q95RtH1kwkCfFcgjqQw6OuE6vX5Psv/LUSUhj0/uK6/afiUQXQ
afgWdXuBlI62XvICvJQkLcuaa+KoyvnaQ5cz2FCXtJ5MWFagmwvgbTVMNn99
Pdntecx3n90khBn8FKFsNmm1Bln+HfXEljgX8957kv+X5CctTmoMCe6bfDWo
6fmN6a9f/IgB3RSA7pUikMBARAi4F3Fyow9uDvOWY3H3uE6XmkyYePHkzpSM
TfQJ7b1FK2MSv0wferuGcsVItKk4iMEtlt2ywrZAdVNhMv/jXplB9ug3DsC/
NuM89JUj5W0vc9KUt0UkgZhGchGcbXanmvmFj9UnyWxV4JuD4Aks2yC9jDzx
B6JwwvfeyZ0rdZB5GfZ9AMpAgIVLIrrN10HUVOhfgLFOARXYOvHvQaghxuwW
5Op8C6u32qnERM92mC+xrxTGbrEGTg7LDq+tNslKuxHdR8zzaw4YaYzuAaOZ
LSaCW7wdeI3m3g604iqScNdWsyq9/m2hacjD4b2kTBjOGJqM211YfomLvy0g
X/p9pibHKk2PzyjCcy4VgcHJoC3QFqQmLY0tEouovkywF6k1SedeFRvon+Bp
H/MD0bjWe0azAq+3kAZ5axCpgHwoI2iPaD6wWZT6jpUDkw8h2pdhCHAm6Ixt
ap8o2XrvYm8/oDc8995EKf3kE4C9r2kjd0qjYqh/Zavk0rw5zbOEzivGFoLE
OX5E3vkdXNYujHqV40Fxnj0qqPnwGMYMx+MoWyHbTtvNfCp3SV0sdHGEOG7Q
94aMeZSx4SekwPiaKqHFgiCIw49Rd7hco/em1eHd30dkPYNbN/RQ6LBJ5EgP
f/Vv2BLAf9LeSBt6EtPI94JfOIkP/zHYqkDJkst2dXZtGe8gwbErjUKXaftG
EJ48WE9/SHcgKXlDT/aRDjchzqsD9613UAj8QIP/BOCSuc5n5QGxHP1Jn1KP
PBczimGj64DT7GXnZyDw7Wypscvi4WNZ7iOEpSpm+HgvRKHVQdyijc8f/iOr
MgTXHO2k/7ceCYiLfIFRKRWo10MpR4LtM2W7Uyl8YC3B6ZXQEBgcAODbHABD
vOnalyGh7wnYdiyVuUzEv5TqP2awepyoVCDJHlNornarpIkYvd1T6W7eu2f4
L01/fUQS2+O1Hk1hHOMqWnJIINCVDmEt9ssLn3EIxeb+WUKWVCVXa+0xDVah
QHWd0MzLabPkSlqqsOAdjuc67AT6wbtaz8gdWBS1204nPb1h+MKendtj+SNC
Cl1qJYumZqaBN4YGp+ocuc20DItB+TmR3v9xq9j4RQqolYHzLlScfZQ5RCJJ
NTvbsjzkxYYB5MCqNCrAKQtdtC9MD81Z27K1SVp3mDS/Ybbfggljs+K63C+S
u97hNHyZLmgDdGHr81CjKQseWR+bQ0jvJhK3KNy0d2Vv/7DR2mNieqCQJKYG
HxGf6lMiPc3WV427H2DTVDHEAUB2Ak2Mt9znPTN332eW5qDXWjqRWnGZhvh7
SjzmX14WhZOfBE6T4AuvTz7NqsnNNC+fx9j7l3WVKFOtDU2p3J6mexmbjRJZ
R0WJvp7e2bQHPw7EWR/6Bejbq1Y5vuzc/r2Jc/TSjk/SleZ/9ell/oYlb1aD
bIU/AjZlfpKxAuEB+6u2+fmh8eStogZFER0jwvwmSJ0BcKCCl82S4MTEe2RF
XycBize2fnwc5fbEEaqoUdmPhhAkW3Kc+aG1be02dOP6FrbgsqnekBoV662r
/ajh6H96jEcSFngjNDavRxWnGezkdyuIXQxOE6uuYS9kvmvqBpM0rMHWScEF
BjArNcEFotpxp8eXECO6IkrrxMZOn7epw2zo8TzafRYvs1UExYOoP6nvilwS
jBo3n/o5veOe9W7ODThWiUqNaoxADaqBHCTI8tlCD9n73e1TsdfzP0BhzW5B
7L5ZmtERpCTdjNil3JT6Ewkxc9/y57S+355KgVlKY7uBjmyDGdxDgbjx0dP7
x/q6PQfoGcmI0g2Fp1yTgMBneJNnjzReViu9ZStSqFS6/DKT2w5iAr5Jq8Nd
sOdO53oYp7UlImeuOp/ubA+5DKohRQPTkroe+hNRzJE2iYAQoXFBA8N6qtd5
oiAX3rP83d8Lzf/zkQw0YQUGmn+0VMKN9GD082FcajYD6MUVthkzcuxCLUYZ
EriNXccDBZYbQNm9CHX3kaNb1Ln/y8B56YR2p/LADRfv7gd4lBNXDHFK69Jy
xQQR3KMDz1c86BtSX77FLkEn7yrIUrjroSx+KS82jQPFXXWOE7q58EijGIUH
I5Z3nUP4o8Y0hEUhp+9AKOfKUZiyJDwub/F8/xa95bVBkyH9hw/6QJQnXbDO
a1dID91MSB3LhK6ux5j4U7eoawbvrKjnurk37nw4JSlAFXo2jdDkq0TBAlRB
Swdx7guK6qg5daz/ASCaHLU2p42t7tekm2Zsa4Py4rjpgATgNiDo7KLoC0tK
AQCBzoAvHvVRnqQJCa2dhcJYiSAbj9yzH0qfGHGm7bEHK/PM5ATmW9Y6dj7k
W8qqo6TYtEyN+nz9rF4VvveD2UumvEevRQHF03fuzljr4DCKfGSiUB8t4IpS
wZnOfuFrZNgl6t9ZGB6IeBQ7T0A/JzAlQISrms4PP7ugi2cPkywDt2yGQH4w
ZqZnUXcBVBcbzHnG5ZrjTakqgqUGbRgYd0V9ZNgxqL6CSxhjwjtEbYRYTCcz
eXi1Gg86F87/J/xENSGzfhsD/R+uoJe0K7Za0QLTCctuZuo9W6U0lxRjXoi2
lu13zTwEdGAgUgTQ1aXUNQTNUvJobcjMN3VeSWK9FcdJTG1l3lKllZsCszVY
v7/LQSCUCyTK1PrESJWP8yTMGoEpaDgkUWW8xw8tzJGb2v9eRddhqYgLyacj
beoID7FsDwiua1F8RHVecusKCZB5DEsvuE03UbO3+32r4DRrCEp9etuZLgyJ
xX1gUhMV6ODD08nklp3WnSrUTuQgvgNEZClp6MOhQVAE4F+BmjJO2L9OlrxK
ozZtvo88InjG21gbtJA1E5WGCHRVZSFS+Mf9GerOYJdMnp419dUacsnFddvE
b9I4UDJDX82xllmtmtNzhJEpAwccv3Zh0BNzSY5pJzsZ79zdeKrzh6dP7+17
YLFDt1S+xOdb8tfVuaQ7WuGggc3/pxqgKjNObAJrL3uNfZAjeGZ5idvx/jfG
fLrpzV52Y6wosILi8RaRmD6poyIfyjaA3UbvIrWC8LpxgGlS5am0361tsvQP
o7Sj5/lsoxGz+EIej0w3hdSf4HQCEzBCQkIMnTxWT5rJgS82yeRHyDg86wIR
9Zo6afZy+/qD+Mc81YvfWbAH6IIzrynQNvvHPyOlBmnplJAfvxnFobOi5vr6
glxf0Cv+l0j4LNI8aqnG1H+Fy25+gQahuQeBzlRGB2d3Su2+JFvAYHj1cjUN
q7etXRq6alD0DI8ZtgiH3Ds9GobPQKSWsc2CeBvifyDJbYXyL5c7E9do5pUL
jhM7+d6pxDgfDvZSXSHt7PtT/emXSCfRHnU3odic4gqB2fg0KtSYAAJmaKnq
rVZ3BEHOc7bVIN0lg+2hwQj+sr5YpkMHxgL59snp7f83PdtBPOAjgdKnu/gV
61lDlcjUjpXOKpNMu4Ci/hm6joc2Wv1jYbDTMvDOogU5EnSWi2gY3zEeakvq
AeFvwnVWnOykDb+LDXVJFEJWegfeTjLrCJK5ZGoziHuzhdOtGSjX8hnoeHLH
lF1UrcMdilfsdIxW+ekYjEwJ69GcXimLfOCzuo0mm2wouDyWzE9O1X3C1lB7
eblAnC3JkBLZtNS7+ORqQBTi8hM4MD7XY+5hwJ62QaFeyliT/dzJGOrWgxIB
Yr7HQkewzePVADY5crCzjc+OklaKRyxHNrGIPAiqAyc8JgK8Afp11IL/7ppm
paeOUKRHw61FuOx3YdeDQde9ytX5JxtWoccMdOOvGLsL/DWgXG4brnV2xdwq
+H3Njdrej/6XLxZ/LyQqKIvNg9lIl24iSRKLC79T9UkwSvVUahanRi2zH/LF
9B3sYus+7PszFp4XJMa7elH+XzDA0w1jaYNhoZ9MERAAATqxUiPBaG/DDW9+
p5DtqWVhQmrCA59WBCT1MDZhLP+Ev//uZgDDDkg6UV64RTCaf6Ib6YpZZiaD
0JUUwRlIWaoSdaQMloZfN6LVQlvUJod8OU69radbuPwfjKhr/JYiPXdV1MTH
U7edl6wMnElZPWGtNoIFyD/GA3ZggyFeiwrwVudsWsXKsP+e0WKrK1tUi3ap
/zXMmBEHZWGe1LhE+WceJXnn6TChYPnCjtMtMEe4DRtqdixBZnibpRfSUA8i
/iorym2CUHGBDs1XTgijqoEgYjEDDPAVkbe+1XV6i4ugcJwSZ5sjNVp8R1P9
iyBT9HFoI907xNMXj0BBLgCHL/dT1booj+IZCXpNNeu7TdA4weicFarHeov9
l3O4U28oGeT2JOB0lf0qeJbdCkBqJbBgo1PA5XX3jS+R9DrFDYFXBq/kW9Ah
JF9vwIWSEPvNMOApbrFkC5+mT52paEYF5maZPXgHSvCXNvGxGbQAKazAUGVf
tP/sdQKedO+XWpDFrOuLZxmbMm3Ug7Joo0hMgnodMdOmn4t+ZYdYcovRAjBX
dEOUqNWWnWLuDC7axtRZaIeYLrR2w6A0ihLan0uDp70xJQiIWOA7bIFFupLV
YXnTn9ju8mqTKrHcRfxdXdQUMXMGAimAY1H7DU7US09qPFdSO/jinNcgjpAe
so3dArxSQxdWW+wEUvh6RdG2fpBzSxNGtQq7xSGVNraCRxKVQ9u9Q/F+izjl
+SAQiOU4duab1UxbAzDx/0TaDMxCquzG+atkSKafDLhAJysboJ6BFhqNB05E
wuWxmJAdPDuYZwjNEqi74VEXv4+GSdj2+5iY/ecGqNBXwg4seadimllwXcVx
8+gizo5tcThQ8qClVMshHLTGkxdzPtFdHF6aZxmjK+wbjKqR+cG4KS339RPS
WMDmmft6B3WjTWqjTrCs+mzdALA+WvFGBNkMm757O+wB/b8Dz/7fVe5uibDc
uE8bsC+kC+tEUxBAx+jPG5G7ygPKkC3LGJV2RzsDPmKA9X98NpjwF21rV+i/
IhT+WorTfGzTgvXbuP8cBLWBG+ffxqXlEwFg0MGtzlzYuQysF0xBtEyJQL4e
h/Oq4FNfBqg7B0IRbNSiXT1Zg8jh47LM0TaidVXY92FFL7Qh3Ix9PP2q3ZDq
om01mBxsA/phxU6no1x8dgb2NobbsZ4zfb+VZ7kyNVx95sm3zQ8RnqjBJo+C
MBviUluxstrLHSES3mIWCuMJMWAxYHqB60t3Lh8NBh+OT/bEWxg1ebM7M3DZ
1+TsJQwdeqbZE6F5b7RFNDV+9/Xns1l76YV7tMKphTfytDJWavpIJNDoZI3S
KO44tl2ffLEtg/rib/buWtQG/p3i0F9/JNdQj7GbcdWTZFJTygFf3heO25Nn
msngdWINoW0QYHVZFMkTUJCU0z9RsF1kT4mXrTqi2A+Di0uWy0zB4ug5iXyX
Sdl9gxgSw/v69NoSZWGnfVsS6OyqHhwoEYdvLfWdBC7NJJ3t0I3BqCXHDiyx
gEU096Tjfqc9tzbA/jD24URDoI64d1ojhTZ+Uu9GH5rlX8F7n7qKt+cgWmhe
T+AXWKIbDxGJoq+EwghNdGANFh8afJkmd7MAgj63/Sb0X4XmIWaQ9xzx9UYy
mKWndd5H6K6Tkeq6ORswTA7/8qxOn3ezeh/MMjw3OViBPwxuAPHXicM5/9RK
WkQV1MaJjcB0pzQknV10zVgjUZqdJevf8RyCZi9uDQiNJgN9U9DzuEvUEepl
0R711xz4lVOt8AQFazUmwLJT5Wj0Z/iFuX0TWN5KM2w+x8feQyQutvAky/6M
sAUihUgUzOicgi0pVatzcDSzUbGKqzrvsfdiyCEGTfCTZb+B+tddvAts8xst
ALn61Buu3vY8o3QbJdM7LteqoOYR2HZ2UXzUgN17XEOgzFYwKpsozaKz96FS
x5n71q6DapNq00FQel7CvtGMZ28pn/zA6Jl6btAj8l7QkfSkhw7TxRnZhE1z
RTAmuxL4S3ohPilZtoKhT3G7wYL8udh1k0THVZhg0DaBSoBCIMlcvDC/Ywir
67QwQM6vYp8xKRp5jsx0o1OUgFSZ533QP6r8UmK42FAliLflH5mIX46unRH4
vYutxfGl6AMI23OWLGOJYgKEko4P/eB6XUiNarA8pzhQZjvfg0AHWYfU9r4F
IpTaSFb+IvYMRw9VpHO/aIPdKad4HrVoZFtEzAQwxp2WTOy/T+N+Pp+aF7QD
QtwIK6/d2Bd3TL3M7ajFkAdzpkvVgxVYSf7IwDxf/qcnSudmy+aDwonTQNmX
4Mrn/yOTKe/yWDXNsiZPiVz6DP0T2MuyK8fTvUqQbW+cRSZnHIOPXf4qNyXl
W/C2+PcE9iqUC7FalboEaYPTJBGCaaDUFX2nIoaghVdz5+hFzseu1L/PS1Zt
RnRjb523nQ3IPwopSmCiSDj3gPucF9jdVcIjewWYQag1yQnVhcxheCIVLG0s
tPOIOhk7xTk38wSPssILbif/vxSyn5Yt2K55ycGWfLwEofrTbqTglmovYvdg
tJGXAco105t5e9pURF0k77DUMHwWKiKuYENmBpo2Fddmruzeoc2KtQ8ICwq5
EpCZv98Kzobv4cVp25GNHRJSSw7LODGtyb3QJn4o934TW/LsV98CIPRDyHGr
22UTObnx3ylx9NcEyQo1tOrVKn27TbNMUoYo2K4KrIH4BZfFrtEtGKJWqUBl
ob4DCa/jzYBvo7fE1J2/yaC84rFKFIpcyhohV+vFYIBtSVoSg1OB0Ybf2Qig
zs3LDNZovl5i4rT6sGp4errZV8AeMz1SFLEZ5A4HuVxRbwvlFJbPfVmqPGqz
F5Kj5/WrbCQN9uuHnavF9dJyOijcS6Yhuo+WBrMXQFoh1BSyhV72/zfI6z1G
zEmpHl8xWfk6XyIXjZp05uO52waz8umMuOLoD5I7BfkMtOt14v/nXriHRLD6
rVkBij2Eql9+SE8twP9kvCquI91TBR++nAOU7yczjVtYzogZOwJwl5ipr0dd
1Z7MMcQhzh2uBanfpdgZeDIvSTxy6Acrere7Q1nI27K9SjekQOZpt8hiuOeC
cv6HJ/nHmaZn52WBfOkyxNN6YxcosQjLPQOPlBYkuiYC43tR6wvZcBPYXTmI
CHXXHEL34F3tI/lrBr8p8KeHaEEJCv+vPTofIZq5VK9HtHZiSDdZF5AxcLG7
ycLc6iGohAaQO+P5wzkAc2/ctqK03Cgm1/mZenkjy+oairj4kdTeNEAsYc3p
iCvSPWifExrDXGoAzCfFiH0KZDvNpkI8R96hm17TkZkBClkG9IMtDl0Za6+/
UuLGXO+SdLvsDOuGQ3+iAqWTpc91xe1PHWVhmUdLRviJC3UfnxHlIVqOk6+U
BpibTqkYXHqeaOSaN0yBMWxJynSbneFRChuy60NuN5XCmm/SsgOxavSrissk
DMDak+LV9uGh0pZpbIN8Iv4ZzzeXgQaOE1mjJDDYOmRpWRmU6LSTgqBV+CbN
jkEOyDOMOhjLOEZZi4ENaoOjZYUMEHGh7nSm9DD9UWOrxcPT7djQHVnoqFpd
ADCgb+AcUi49vyQ3orBFZ2yey3LR6XIQILreimwTmnmva4AyPang3njt5aQ4
Lp4kKtaHdjUvvCX2NQ1tPpQyb6aOBN5MqUjNyia5JRvlrwM4NPFJXILq+S3V
1Pbrrj0+vkhwtnxRNl4uyks8upSNtxLbLIMmZNcHnrmgAB4c6sq0YSq3bNOX
tLwEDDalS0bsghvX48AmbTHWiSqcM2Y9p5J7GaAODmI8Ro7UA3gT0Jpehl5g
hOa7HppXEyKGgfC5Fzu9VMkUr8pr5DjswsP+cIdtmc8tMO61/cbsGkSG2ioy
TVP23O7QtVNEDeacghYTEo63mAyvR4BP0LtDfk/9U6sSsrv3Pf7kpxcMPHg5
CiFyFGY0IBLsi4Mc33fzDoHWUOHcBIYj4/TUMiSpN3eey2S0V8MgPLgem9Fc
akmzlnP8Jt9f7lFy3FD5Q8HmTEoQ2Ih/K7CXbwMyI8ecMAYkv8vTqYdMsRAl
ooGnUkvY7RNV8q8/UY/mLpWbYh7MHCcmfaikWj1+LwWhdI1vlCZQ89LXO7BV
Zm0aW3hP0gYzNoBd525RmZrTMyrMEnYi+Yw26W/5eLo4wiqY1NpRN8C6L6pH
WYgv3z1Mne/CTf9dcLC67znaUTiCA7z4OEy6atiKeunWg9cf5L+qspP4dDlc
2gHp/fSoVY10SVCuSdTUi4ArtO/9hMdk5OYz9nozrIOMZ1aaM0mQFb7rNGJv
JPIV89ngHEcEufqfFm60HnR40bUxfIW+meEPY4zpOBsvtX6RFUzulHGfUqUC
uqiZdi3FIq0ltvCDTDH+z9RVHTB29In1xILjpkxY7wjScStHyJvLWS+9eAzY
m+oyWiVAAlO1Fc8AvkiyMi4ipfdAfwFQbTGrk+qZOC+cQxhG25OhYTQf3sns
V1txuA4SyWnDB+s7e9au0aPYMeH+XpxMMY5xffrYSbj4Hzzt7rvBi3jo/xh+
gyW40noX0d8Yf3Pg0Ldiy5j31Gn3xG8P8Q81vzZEj/YOWZ270gFE8/iHrxWE
7OkecR/Xg08oSUyoHtoIilBTTuir+c695B+dosaEg4qshr7CxfVto0xGj1Ox
CzPaX8HeY6oyWkq0efvlZ3Qh/5qORy2UzB9R/Nb0tgWpbNCu9Syu2sThX6Wj
u9zNr3M2xS9Pth2KeVLE1KI3udeh39aq4+w9RIHUWAnZ/FRRb918+aGbFEaJ
jl8pBQMM3mygXbFXNXPUu1VIqAngoR72pmVgnBuujDVSsC6HJzIPD31bJFP8
f8MSw5fMFhfl8uMnvdtvKvm9aGuEWpm8RukGyNAnFiF7c+lofx2QBGLa0QgF
tEEB/ydencVRdrxS+mTtExOCBxbUIF78qptzIKGRNYxzfPESWokxNONtDTcX
MKXnaiVTStz6WaX96upm+TshClHmJrKFFWak4981JBAjYASbqvRrBnrKGLyC
o8I+W807gTU+z0WQya1QNb93FyLNugFY121tMk6DHcvukqumX8de4UkIRhLF
Uc3PJGrVA/oPkNF8niO22r7j68IjC5xvyweTmrpQfyl9lcCW28drD6PJgwId
8z5Uzjw+aR/PADFN3/5bpXwZd5SKA2utEgqwExlHK36gQPojw6G2zw2DpDl1
xHCfvEcSmtF4fHz2lx50HYlQdyL2lPXoppmL6iHyLSeA2zvQpyCSdU0oCAbr
AQMQvSSjx8cu9J2iXVWbGQBsmk1x8+/gEEVfb/xNFqT9hByT6f9Va7ZqjpL5
7xES1fQ1g8WVmzvs3c7kUKnTR0FVxNmHX99VFaye9xLEN/vmr9kihKfRjKv0
VYmxojLoMx2VarNlx/GP4pLIz7b9iHHT0bKTDGk/EH2R3MaOaCe0CSiiXJnY
y/55fsbxOtY35r1yJQ8SMveWOwIdSqu/c17TUeebhPTbWKi/jEbqkBYH8pQz
0aQh0RcxvdV5IgDiexxyRZ53laemcem+5uaRuQqvI/ODytWUHpVCbAKr9lYr
J8ntopST0L0dl4jcI/ZCJZw9o+8kIVE6JEw1fDDQbZYr/b1ME5xAmiQA9udg
D7sqw8wSVWYWDGfauvXt+LR5MBfJRXZRQM0MKXO7Wmkp+qCHSWn6VDT7ELau
FSI+bTbXbkvVbvRq9SO+h7Ma38gYOtWcATcx8m4SmM2eu1ZzoJJTJeEPETzr
fDVqRpiMAsDdPwVw+IyHElgvWh7zGVeoXl7558cpdHIzGYavvIssYOfdBdqe
m4iDis8yVJZYSZvjv0paO2Kmk7wwf5jLsaYDmu8uWKrKOpMQUdEZ4reM5nNY
rf7UAi1A0eJi7/fZl0rRyDMW7NdIiWkAXdMxleA8291aohMslPbm+OkZ3Emp
gZtFQj7TWf2mp9Pv9aS+pIHYMY7o0zu1Mmdw1sgE+DApNHAci/ebGrCpNC5V
FI0AqMBeB7oyCZXrIpF1FXElcoj0u9TqsS/sMA3P/KcGCmJbnfZeViTh2thN
fAPERcKAIh3XwIub0jpo2ye0bKOmI0kcDGbxR5acppcag/iKeZv++U+DmQyb
dA97PYEPHknjF+ltp72an4iRtlJ4mrb7NYG57lK/L1cZO344mGGhT3P3ctZv
cxuHLuG5dbYUv8oXVr/46A9j8m2GnihNqgI+SvwpglYNJIa/2fi7xHKn2+3L
lI4gesdpr7OC2tJX2Vqs1IK+G+oSqMonIvLZmuZA8gltV9fo5MtamahcPPdU
M5yPLBkGu4MgO3AFkLVP12HSKFwzknkC52BBeS6J6rniIuyefQEcnz70qEJe
zgggUP92bDBLiP6NvdNXL8hVFVMAd7MX470PjcdxggB+ir4Yl6mXV2QAEyCS
ZfWKr9ifOvF8GKldyn7tjxBo8K/kyNxZmfPBdsbESDiCtcx0gE1nF4hqEGJX
PsUnd6fza1fvCaN75SVR8dEMSwOUAv8Kv4d1yG9237Lm06QwOTwwXYY23wSx
uYUfzcyC/oH3vZuEdCWLDfqO/jkIlFH5OPxG34WOrQY/r0Iw/UBK/xg48Sk+
657NPhevAToBvvajZcC9OZqPGB+sqSvfNboEh6XcrJiTiS0tgzEf9Ft+TFzA
fiR1XDdGSvOFnBjuInYVhht68mO1vZQuSwuEjvfS2gkZr/V+0TAQfl2Qo2e7
XL+6D9M7VfBlSXWI8R2758kO9FyEjDlGQzqPuYRKhLEZX2sELmASUev0nojd
i7WsubaNf7W2iO5qJIls2tPfyG7/zfZpKEUNNsrwCTtEgPBQyGBx5v/MGFeg
et7wRoYvIZ0aK303OQTXagyNcDXbz2aktHqrJsh3fH7v4a4/ksd6NxJlRPHL
+iSwpjdWXsy1JrtcZoURBc3HTBlRMRIlhoqGw2BYzbAWGK2uT6UXeXFUVAd5
vUOWA3HrFalLMISL4MTDYO5A3rP8ddhc1lZdAjB8Z4FiL2iVoCMsM3Ptxldn
2VMP6WIF39ZZ0wVeCKtuKJoiFYQ0L2mcr/ggmGNF0qkjLARl15P6eykeimKv
a3URjOMst5mE0vlYrq32XaUHaoB0S3AfxRlx115kpEQRhGozRnCg2rK/IElq
L7i3GH8q0/suSuh1W9YxQMiZyYSiwRV8pdYbvIo9q2VIvdURCd3cVNP1aMyc
qDANomR6ClUwUW0mzUS4Nv8VKY1Ny8ZfnI4Xg1LKu9owMfokFV8p6IuVHQly
jGKROaPK9tTmU7K3yNb33O6YVFPBUOLkxDpOM9+5cRgg7Qy7j+nm+Veuz9/4
neLDcuhUnnPIGod5lDbf1+OTPaCF3ngrp3yzxOevUNyqcTqaDJJGbmuLZwf1
+sKBGYbdYPFAyCH7dhmLac9xYsIYGgD9h5kEp05YL7MOvVZH2eMx5tMWh1Sr
gMq5hSdbEu11bgQWRM4PyZ7D0SeuvtPmCDdhNo8aHWGvl2N+baBueKcMnd7f
bkHPVgETxQgbryF64tU0XZ50SG8+MBcpWS906Fta9uPZkibZkb4fGn93ef/P
+nFVbIrQ79x44tBTeI5QVGhQI1Jf6Vlk7gvFIWbMTvRv38GpmEqg8/G4xZ0H
h4gMnh8+vymd5bU3kmAa2khFweUO3neIoj6icJwcy0AenBFMxzdtAjQViCn4
uGGcThzZi6OVxwUzBB+kiNBawDRxFYtyn7lLb+BpZKBwyy7Std93TIys0pII
pTXwBJ3jS5Kz59pCDrykNe2cbV7/iGScrXMNv/CSyj9OfVrR5ZlPuQF1cdPs
lNyrr+r2r9McWRnM3UaBiW2xL+tnhiMGTW4jbeJRjFLDzZ48ObViUAO+ZKRN
rw49DvivKUM8nFlzFfq+jhjNg6p9J9xVDu3tcxPPvyBTGCIDzjt/CtndoAiu
QCX4zcxCAXEr1VmZzJa7Hg0Nf9T+RAkJHBI6sob/5KlvG0/ylyi06wM8MP6k
uIqVaLLq6ouj1tkcJOyMVC2YKVAcuIpyheHMqNZavvCjvR72ZB9Oi9d7Gq/q
d1yqvVZpSgpXABm9TxtH9c+V+M925Q+yT16hFphWiCPJoR55tmUwL2S+arcE
BBagjHy/2dzs+wxHZi1FBb9IIxFsEOj84yObYsrGkqWqOOkC1A03iQviGhQO
EDcqf98LerYA6mj0gBIxF63tu4+S/aw/mk3wchm8/YsjPNYVqTbrzkGuXiYg
A+QQ+7ADxqV9eRoSUqopk08kjNbqLAPNHK4OCae252QXdUwLSGswfmsYeIsS
EDSX495tUSknlxDvGCKaUgmusE+u4g1TQ3pZIAIsW5nCXAQFnhFkfHD9AMOW
egOnpMqwR2BYILHTdpEbeJb/qEEWqi9E9TMMWcLqtwPVCSVgDy92RWP+U+fq
40NOq6EvqbfZfmaF+lJXzWX1Q0m3jBP2K30L/CTCFYO00yUeLH1N0DYiE/Ka
CloRUXBfZkU+qqXCXhwbFSso17JqToXXMR33Qe2EA+nYSFkTLCCckxG11kM8
QzkQq7UlGZ8LggVVsvQDqrAChRhggZB6gGgVRJyf3Igz4M852+6wXWJjYquC
vWABtdpvaSqUbkyATc2WCE6OB/MHcemKsFB/6XFad6qbvJ39r9cM1h8fkYOi
/nUn94/7eo1JkZThGihDGo5XxqOKsfhE/DoQ/pOEk1s0kNRDzpn98Vuia2Gt
WDJYvlrIy6SGnWkHflH+iwCmPh4xhuSCdZWOM9D9D7Bmqf6WqZeGxX3C/a1w
vuGzKK5vHlsQAb1M23WsnUojSotaQ8mxLM7ZkVsjbiRMuLNMcxXTWqmLexG4
Zi3x/oRDWh3A3av1fFmzIlVDBi7L9ZPHHuVbGDOA7TkM+2jqXgF09YkcWjbg
SU9chZ8eonGAcNnVGYz1F1lOU4g3Q0T1VjZuo543i+pEzAMYrgkpfvDpl/fD
utVEBiOnCl6MvNs2w9+cIDwQqxzI89eeqIbL1XogBDCJnFpLkef/QFIM8Iue
cJ98GFuDOr/RPQEVES0Sst1FKKj1Z5Z29PGyLXe9Yc3MJ2ETe5pOnxjFIuh3
znYJr/lCCC7pduwiNWUxnnnO2fmg1qpkGydrVM5EUjbVmC9ThRUaVBy2gwrJ
tsbOD2bKjCg2xNyIXRHgej5kaU6g89jtpi5tSYthTiXtn3wYaio7g+otDbjY
UOZgFRin1OtQKenujnImSkjwwjsoCpea6LUCiECAGNzy2TrD5ZVFzasXWaA+
zT3gLNKGw+VE3HHSnEBlY/7mBJMuxCVWJ/FKZIq8DNrzNJQqSlFLTqQXTS7O
QBNhFW/rEUtFfXuD500Sww/oOTcPAQ+oGBRDlphwi6/8KwVDa3Rj+VssmWsC
MxN3X04LyIzV+1fmXcNIHYURS4l+vKz50BccWGu2PrkYqIRdf6D+5mTUIgJT
tIanjxSNqZzy+GVuK6q9YrLSYYq0rjQBc9KR2uWyJDRzvtbx9Ka3mdGnIbIf
Cnp5prCMU/M1MjUdrRBrG2ZaM9/IXk+Xt3kCtQv1Ektb0OVa3vIdWytjpTfM
PVYTTwylu+YA4kOvxXvq9/MaYulTyM31XmAQZTuUyTJ4McYJZYZ/WZlbUMrx
YjxgkWh/eKn+BYYDppHKflvewiHvbHgZHtpswQh0EkKDBRyVCm7itXP+aj7e
TBO2iRn2ObS2aJxFEd7zO4tF02I7DvrVS3KR4CjYk4Un2UwjsBU+M8qmMSWb
HFww5g2vWQGuJtTifvpE1OiH9U8FXEY5b9EQr4mCH+Pes5grlZKUAZWS0Q6Y
D1XyttlrBY2qLBtUD4O6F+5uzTNc2UelmIXOblyh7St2IwxvhzN+M5BEp2ye
vZQ4GFd9WKcQMYpnXb3yFdcqsfD3f9lFoySP6iOyRLWNqoyvyd2AWbCmmQUJ
L+jZ55+WpUVPv4YTrwtUIEijQJoR9oVLr1d+6YMdkSoi6uxGGMeq5xtIHRHs
NmLoB/QhLMfDKrw1wX3hFElxJf76wxVcJ8SAzTCPk4y7ow4/JI6RaUaEq9PN
aJp4Y659ob02BNk/ztNIiaEIB3ModnaSAceVyngV6ZTWfy6t2gvh9A9OyjGA
qEu6eYK3fA2WT4LnnbMQlBBZwIGZt585QdF9e94j3jzaN+YBag6eeXi3y5Gi
TPUNv0dxpT8M7jvauFYpp3ZlSgKKI13UrQ87ZIqUaVaDmhkw005HFMaJWTvr
oVATS/Pl6IVDWUZsvLAdSunYBncopBOT5gwFJwFRDPa7mwsqcfOBayd8N2CB
W9MllmH410p+zAB2CpNc/hzWhdsXmR54BlILkZ4Emvq8WVxA/OxqgaP/gGeY
tUzxjermA1wX0+5otbgNfXOK9SZ3NTb5Mcb9/jpQKxo4DinRUVagpw6aUxZs
ml/vq2b9TinJc+mgBNMQ8cTcfu6S6sCoQELtWqah9wEBLu1eWWaZS4EWlpgR
MPOMQmMe/2K3VdPGYpdSYxK35DfM+K8JyL6oW2seZjnotEMTW5yjaXp4Phfq
ficF2VECbzOqsKAkieoP6wjyWdIAGx/XH8Vf8uqUy+F1VQztoF0ZvtHiQv2I
9xgPEezKiVkz/lLJTGIm3mGXYO8nQf46xpsj39MEwZ+YRF6BAOloVJEpmTxW
WCsnzRyihZJDpoaoF3Frrwa/IwrHFhU30VJ8hZIIF+d+iwXTo6Hxc4m0HAso
13khYdQWPiJCz7oJOoAQ7pMQQd/Lna65KKs53XVt/M58Efa2p7jEBker5qxj
rgxCoJpJt+bUQ+YkFYy8uTFNW63KOx2Ra+Qjmh7Kzvd5FNDgoOF8WoNI0TtC
lMROCRe7ZaUK9gnUKFtNebdQykNWobNwEIJReIHQnImG+lEPUTuilUAVgbXB
PcTy9/DuSo6DHwpkhGwrRcqaSW3/+lgs2KOWIRTbzXmaFdQFaT0ug2WIAJPO
j60GhYco/Q0ac6vX6npDgvxQE6sFAfYW7hs4O36+Kgn4PzcFKWYXE896GZNT
1MJ1Wl/n++vSwJ9Gbfgigvqh7GiKn0cY8o7TkPvTFuP3GDwbJhyt2RK6o6tB
q9YdcNhQ1Rs6SsCnT6B37shm2MoCz/IwKjRkUAU4Yi7DR5Juc0zNcoGL42bP
hHUcmp/agm0BxBPET6tHVhoWa8Dj5cIPqqk28qGw/qZ98j20WDuAriR8VqvT
sRwf7QYBz0Q+vkuZ+9akdqgipkKt3BCE8e5VQhmOklp1ZW7dXc0h+9KwmOml
ct2crrethgL46yGfUxBIxSgTZr9tHj/9lkaTpCjX7t66fcFi3oZPB3God+0Z
JK0r8xJoj05bg6ik3rbYIygM+EYrhC6F9XzZLXESns0kP5LHgrdXp8yqAUG+
/zzl8p5RC4b0RFrX+9kzbOB1FhTPbziY38FfahC6S0nAwhKwA8fGP+pjZlxL
VjjOBBayACNbXBblMBMXWEehSPDZTdWQ+29nqCQmm6Fx7Ccd7oumx35ELvsQ
7o4m1vTZtWHl0noYM86iar1fmqJEfTZU4unZgeR1pWJ9wyVgFYR/CPxk9vie
ny7T+0sBiibW0InAmgsbjmQLtS3a4+oDqzjOMhg2PBBYo1rpLpoFsnK7XNrP
9G1tBNu8ZQzVmDlRlPNyY4wBDatODyz7FLb67iGpnFhk3U/jx5deO9YFaWl1
xDWArMNLf5YCb5WHXjr973Ze0zm/fskjIvlBdL+RnaIGuGIa9xzclaQnFsC2
jZ9y+hfxs8d7HHVG+9OMOVMn2jZjZmHZcjhsJaMGKVZGgJF7rxCF/T4k2pkq
nHoig5S/QbVKBaP7gAEtKUUNsubjcwhFiWeSll33juYzerIi8p4iD8kcc6dD
HJlbNxV60rB6m1fWDi+ZVdoC+RlZFmmZWEhHAvV15GmYns6yajoeVcDD0P+Q
sMH0ks9gZcJOM5HVsP/ASRemV1PBEEZQmFMnyaiBXz6Fw65dtuWi0aq/0kc1
m361lY6+UGx5h3lhHVui62sJDEnokV23ZMqr+3EjJUe+CmjZ14mwBqR8MBTf
vdkuQXDGdKzEI5cGkmcWHwHPw68KZDH4F/JcYIyjyKKLUB98XPwhnBrYxZ9i
W/lHEtIAGtiqBzyDaUc732BiMXGnHk3Kbt2LpiTQd24FwIpwX5nXGJAz/Ejo
+ju9kUVUnUGcoNntkhkTbHIMUMeOx1bzlDy+jttCbIb+y35Ox6z08ZX607ik
zcmAfdIAmzM0kiVJoFSLK5i8Rrl2DmJqKeUuluaBkQNr6Kbq9+YV11e45mlZ
QoG55aZJvtdCnA8XF/7W2/h6omBTybMiuylxl1wnczDIGRbfctFnhCDFtaGD
Ul5WRks3cDRS+w3SOA1vx8nW0/aYzNWyWEGL6korNJDQrau9KprwkgcC7kca
+D0lcWzMGgpe5Dhoe+gNY2WlE1Jz6EAhtE1KypFiHXwaY2TmNiP/ucE8y0N/
iXlm0ziQqRAXoF6XsWWWWReZjsCLOKCUt6180YP51Sb8gd1HGc5XVnpxxJky
S8C+6WJjz+mQrZEJfGAgn2oZpN8EqbSzjJjdijKzY4shoGUrPK6m2DtWeTEK
LN2s+gw48wN1o/3jm0xp0riFiKgVuCjkQ31bl6qseV0InbVPl8/+0k85LW0J
w+4Td23SWVYgtujH8odp4/D+L6eeEXomnhJrthjcLChTlETx5QuUmmkDEvC9
ifgVuzp1XUoC1QaVqswWlQ/NG+h4S7w0Ca7+qgtcsur5mEtcjMIT0q2XtEHL
CY/kFdk7WNznIrSVpG1J0pBJ6ZOrRXGkvnsjNgUR0+9rpVqz+Nn9bJDS/aa6
mDuub9eb1SjWPb4B53DHVmLWlPQCwR8A9SjiZlmadIaLXVgjcDv5/5lT3qFP
Oam/VMxaR8UgN7J53N2WIR6dHn9vKOgMg8r/G99uIUIVkMUAtZnR02/jAsM7
B0nXzZ1/MFb98cUeJKDyzEKE3hyTo+s9x1f1xqFS9YM1uvMdaKchzPdSIeZ5
YyhLYNIFsHhkdVbLAF8oL+qLSbSBSb4ZWgm3rnU/67UWD5vfYynr/pa9AQVr
oo/fL37ZQnhVhrbyVGPAH/SpTLQ8omWtHgXN3KiVkApxEbSN0YLwFlTQrS/d
1A5cAhi8C5gdzbm/2zqyW+F8FmWg181o8V/YeyZgXjVFUbOeZhYxEGap1LZb
EzsEClcrXqkUReHm2HVgWsiejdy6pE0UMM9Zivhk0nbOmfIuvH3AVJRV2Fxp
1XbAF2WGA7WFAT1O5pgLYx4wk4pm0zVFDMSXVNGqNxCiyDXr0sYcyjYCN5vP
jog3/a18wSvGhpA97eX5VT2eOgReD6G3WiEsKQAzJzn+2WA16b3xdUTjSDSX
xKWC3T369JCTB8c+nBeAy2LLWDFva9kf8+1E9HhzNBb1MFj7/D+P7ip7YDdb
pmJVQMbVK7WHEHHbaT4ydGIbBAkTrzda9qLK6vpVpJkfhHEgcEW4x4/Gtfhh
O1QAi34xpckYOyi1XFVD81CLyx6TI8sCEFw0sDc/i118f8zx7xDfV5tIWcjL
NBqhpfxWmK2+BOxWrPmhOWt/P5ScaqshGjgaMQpGAKp5gvsMRuZBE76luKSZ
iJz12JROx39sB5Ut6KVghyd9rj/ksszhQAQoLdbR4mGUf88ETkDK27hZGVJX
hszR7mj+T+1CNgqDG7kly9JxLFPaLABFloppEYu+5jel81dL9cqMC82Z7al7
dgP5n6I57E53r4YyyKkg/6hxjY9lzwOZTainySpITZrAr79OTcqqzl2/TOHr
epaxBWzGlGxNl8xKicFEXlw0MMm/DucVsTc/pLV62w1G6X45NiP3nhAeCoZZ
WUq+ukdsg1l7jjJ5uVQCQVopx7QumjNZt5gOtBw1a2vAqL480Nn12Do/WC87
47LjlHfaNAjmcLti2DETnTSBnsgmU7JaK7SJI7PN2bNJxsPL7ODoVIJ26iRy
4iMfstQ7WXvxawWm26d0z6onZRm3tfykAbCmw5Z9b1K3hPPXoHp51sf631AF
ij4NkQg5C6+rZsg9eIKXgv6Vfu4c4seG5bM4pHCqItsYvnkDGgwbsiDlvtaq
yrxJ9Yvp4ER38eaf3XxyyY72ki5wzs3j3DSeSz8/tPrMvdZ3N6U2zvk6MgSi
QoELorWQTOpYfcbyTL2fXBgU5NbtMLg4wwig7mm3CXYaQWzAvqyTTSx2o9Rq
jatn1vsrH6v1tQN79uDU6UtzOHYpaAyJJdEThVV894RyUFLLWk3qIlFHQYmj
yVXH6woWOl2sfP+XzaZPzb7a9Pen3MXOv7a6DkjAmAAzJxBuqyZk4O6ni1bF
CV2wD2alYoZL9Hdf9bUFdaUf2doMRSpiIhxJAjYbITm9uiqc09qwqhmdp41M
gaW6cv4xy45kS5BSVH3yghmmcJs/3YjYlInOk/a/UIjSetfktqD7BvL/FEc0
dmgelig77CtTr9CYBZkdYr7IzHKr4ICxPEQtI0QD705+x4Ms8z/SUFm48pvu
PhuofuYvg+7VKzOs8KCsVJAclPEyFE1n9HQzzUHBKzguRyLW09rCLUBhsp92
UxMG/6sG9CQ/gSAuLPJdsRQOeBI7plXbHL2niiFJ8ZXf7yNb1zw+4IU8kSiB
sM9Tn/Le0LonS7CNlVmrTZBuNk7fzNPC68oroOPkIelTBT2U+u997t72txO6
XMCn9wp8ddhB5PACrfyvC8ZOt7dIH4K1DqqNJfSVLEC7mLOmXxmoiY1kRMd7
36KRwd7ENrL0aXSyvJ/eUbCsBL0Z0nQJndoTR+1igtFiWDQNTfy9OLpSuikL
PWk2g7/V8LVd5qiZuYOgXe9CJnfD8Vax4shgR8E7ngR1F6lkrU200NXDHHDN
WkvP+UVbItTbaUxe2xvu4gWoAzW+LNsD9H94admKu7iUsLKq9dxsW3A5f6ET
Y/W5cDk+3gxSt0LvTCd5XArEkvgEort0VjccLvwmTt5gzovMx72Kp97BRsj3
kD0V/8iKPFBLQopow/hdL2TVlJdRpGYHBHijUFyY+Qo45U+4396kFpndWerW
R+vC6ykDWgCd3idtskPB4/DO/ToaX/4JBE3n1hGWhqI1W0Ud+IYCxXJO6QHL
4/NrWeuANMVbx69T2hMgjFyVicjR+ULxv1gzo6lcSdQPrd2TW64JfiAyVujI
B1PcZhDMQyOpcbAQJqM8ga/u0oIZVrTw+WCz/bAHILnJlizUxLWoFV7pNxrq
cgkdnI6PdyL23GInAeh7zADBx0Bjsgyn4QZI498EZjHGgDBNne0XHlgmMzvF
oNdFmELXsjlA4wNHycLCiNAZC/PgiWHl6o5Y2AoPZBhCAYUOpCVn4dqk7Wv2
Y6+2soCOpu9o0hIY/wkAR8hOvlnmeVPESvVh6llNf9mExmD6KysQ0uuZ1mXJ
7td71aCDbm2Zjjn3OfU0KUTz2eVjCfvYQBInrKRi7ZrYx3P4XuxeerIfapl1
ODlHJZ567WQ9rSdnOzYcyhceLGxbJQ1CRx1J03SIUIyMJVOncIFVAguwNKaK
FIpxn2iU3WO9LLYYPyLAedng98k/wIcZe8xYDiHGjSbwCfPnEw575tuXDxvm
uUgVRafVkfAUemdDdviebQ+F8v9RyN/2Q0KyFbzPrGvEKq47X+hzjwJZxmmN
LIgLftYCn5XOhr/1jDWmqhGhVk/y/qVDM5MIwpvQaLz0ncIkJfj355FNAfJM
AuzKikx9aoVrzinIGd7VPVg/AUjbOL0eCjBxdQeT5upHebJEy1HK3BZxa3u1
W//nN+2xYHucbp6DG2yAbfCd1fTt3tsi5T41BtcjQRyLX4M6D2LQ3co6pXPN
+iBi9BcJBvpxwAZZB94MlFLD6oZchEqd2xBbf+CvbXqu2BDZQrq+SA9cp/c5
FfcPHz8iwvBluinx9TS0iCLfyD5hBYwZMtcVWMFBrAaT6w9idvl6TdRKDGPK
DeoZ800j2v9o12j5PlxDaIXOUBgzf7d2Cq1sPxkEkQWNHs+SpzVssicqRR4f
0IheyMp9pDpMMqP4/ILwYUXmHiZWLtBwt9A2jbMgw42tNmkTTh4Gn6aMTlAv
86zgoDFs+R+TnHQsm83TpJpF7F+j0KsXDOvTpnbS07aqUyH4w+hj/dzMaPxh
nmZcz7DekvIii0Mo+z3oSb/XXbUQO3zdoM/gO2keGwWtYu1BLtIQvI3uYiZu
w2WGj3b65j9GDo3xqTgbegJ05upgFNw1MzxI+Y7ISufmcjEQDOYYM4lloiTk
a39k8iuEtBaihI+uU5Jc1m89cFguasbYFgDVm7VZpDHT8ufqIln7xPlj4XHj
cO1Z3KviVpZ5ynZ0Ss1b9T87glPWTBTjoyx4zdWspDbA+cMGriaI5coe5P+e
LWBgaJZHc1GXqhqVUfsg4kMwgsS3M7MUfRYqPx4GcwT0hT7IDHFopKheBRKc
/vTtnxmIffxYUp0k2CUDeIXKmgGdr+mzt0ncC11fLr26Gy8B1x8IN38I1rFh
432QvOomnUgogfEkKjqpy1mDm0iVZ7Y5xmvEY+z9djqShsWexx49RsdCEmuh
ZeG4bwyppJc76UeMWYjGzNAjO6ZwFL4zIUtQeuMiq5kyjnZ7lcFnc3pn6CDE
GBuBz46l8DI98nCM2cWIZzLm3mvGhmvHdhgDUj6RpDQCxZdaKuhHrA7rJ8OH
/UUGJWzRmS6ndo3J9rBrMz1oszxADpzmkKUKvAqZdPg9ks6aOlm1qkNK8zfO
9YfteOEkNWbNGY+1OuJvN8d4Boaj66rnFPQYv87dx8AXBf5Otz6soIIPIz02
NoxNYfyDz1hhB7D4ga2vxkW3htuBiAKBr/O19Ygp9Dcmfij41FiECHP5RCHL
LQtmEKDHUAdWD/QGhhZDaplimpPdO6dutVngfJkyqcHrYSy0DCPxNL7m8Mur
a/5JR62FZPydy8uiyCq5EgaSGvMmlxfLiRkobPqZyVSqij8EEHrkKyqFWkVb
bssCuSOpthvjuE9PI0e7ILu2vsAf/HXclw5nHv59B0g5jzjfb/eoRIdpXWo1
x2VjTXPq8979nUeChexLWNE3VorvJgkMwsE5bwABxt7ZWkpPSDtZAHqKYiD/
XQT8zT8p40phFcGxk/ZQmIqyYp/WXiGOv0i1WEgSP7BmB2t8yzFz76KBkOe7
h+VZiMJRbQbuyFasoHRKgFaTX1/81pU3TZYwR03/K941Qceu2pXDa7iGTGmv
GqCxQ4q54z2n3wD4srY2h5fMmmdxcYcpI9zLJvgaGrDJJT2MBdDp6/SYYQtv
2chezb9UEAXolpFWdqVCSkyYtRE3xr+OF+VWWyntWgaMVns6oMBn+gauhbP2
5bdlz/laZlH2EtfUhSTFKyg/qDrc1DIbcqO471Xn9T4aw2yzo4GAS3UL9iGH
s66fhu2jLJUw4cR5V5922Lk7KkHIxTZhKqg3Ue1+9R16I+LTcO+Ev1wYV+ws
uyyW/Al4xfAtysTKaWvlkcwinik5CkNRl9XkDSZshdwuZtzxrj1jdJeUEen9
NV7LByKEWpc6XAVqeoKEJU9fPVCcS6rAE3F042glOXOf6rvg3vRH/BWDAg3p
vOf0m86wpLjSQJ2ukQZw36TWX0WoehIzOWRsPPKyLWOM9nTbylHHbbCW4Gva
zi9ocDFkSDIvDidWcLznMyP0+ybp2joObr8Wfwb4DEBjymUz+qIdcJ642tM7
2KKD30qVRz+NwCLS3ALAGn1hKsIuTM8a9PPjhC6p0ARdMIyzx7lWrRGSv8uy
xE/kBxuW3dOVEl9DaJCpuKBWgOyhxNjAzXiAkwa4edeJ+u8eH9jof+L5Zq1z
Y85zkOD4AWBA489gMEgeTizVP/SVuboH4njKmTp1YM4+e9alif8SUEIHNW2V
XzqLUsfV+tTdwGgDHKNJBXvfVmetk6Lo6CXS3EckJaEqBrKCa7h3fYocfUmu
Yp4FolXaqTQ8JlomwlI8ibWml1RwiCELC1UySk2T/gIkhG4SzK0/ffuF4qdC
M2mnDu0cCqq9+2idHxZ0XGpUxUXzTpJCNCzlgTVeederqWBBVE4jRPgxm0Qu
GLNgdTbxLmztyxsRld9QP9KzkKGn2uRVdr4zts9OxEcQ3t8HMi2MG0qeC6Vi
NeGc2vBImnOoAUpnTkAHvAPVYr4oHX6ShaHeK4znNLOXcOIdLfsh7zKsRNnd
24tWPOjwHdST5yuLwhe9NKaQdbFGFh2ZqVmVg+m7OSqcVMIo2gAzowBs4jJJ
MkD1xIqG7E2S2fsi/UbSeZydY/xH6A4DMAXNPMY4KJ6tNcV2HgcpfUatjvOL
k9Iq78SGVJTW8LdtU4pkVvhqGBKZptjVV0bn+iODN1MKFFQyOUw1u4kgawS6
FdMj8JHJiJh+orT4E7+z7B+nXVd9OrMHgJQKH97Q3p1DIEac8dJ963IkEVx3
YNum6R25XDwukCBHqy+K0iPR7BtEOV4wvdzWV2nmYIBgmCEOHBXC4rsXvN84
g68ok1FPO2LAPRxADiQogX4nE3Tq2VVpxf4vdPO03B9fc77uF5gf0fP+Stv6
nbmHIj9x+ZR4VRHjuWc0S1kJvmT9aKz4RdCtEarxH3qKRvpW4QEAUijAIIsB
TbGbzUEMaREsRplpuFObzI6D4rw0qYk8MBa3Z2h7bC1j8Kpsq8pJTKa03pV4
mJYBfOyq0X+0HBIcrz6QousZ5rA0KdWFii0upv+0bKLiy69xRnoZ9O/PZPik
ldRFJni1BQAP7LajWEEz1N7rbvMNxO2gASd/ZvzeNWavYLmDHt7CrQQCXs22
MW7mBeYFFwbnNIVMKwGRK7yVzmtciRuoGqpYfB7x+cuJ+d11k4LUP2Wn3wiM
a/73VPGNjQYB4Dh+Yoww+0475hc82k4LeMSOXat0KUwkMR28Jv+rxE1/eI0N
qZP6LarB7G8PM5YmGtQ/xGRss9oAYXEOZx1fYmt4F0dbqFyC29vpPwHTFx/M
u56Jv7Q+zHf1Vu9RL86ai0t3vqbcxedmUHfQr71xDr4XUHkL0YgiUkrTBRsP
f1Vn31xR8SwQSHKGg1+ixyle+R2z+oh18Okj9Mnk5V8s1WgLzUsgbEWfFpi1
8yr0EznY7KP2G6y6Y4xCeuL19vQJKKs3omjwry2HiYY/GYIYkJZ/jWfrKiYc
p8sX9fv/Buh/YmsvBl2MTQApSSQ9C+jKvNTBmRvm0vHNrkI5WSMOfvTuN+H9
H+GJRLvVaGRPkuVktXH55Ri8CGKOJfTnDIgiSksH9zhiSNKu7wqFmf61RA0c
y9btKqaX2lAPycCVKfqL6brXi8lvUJPOF8En9VqsFjyKrQ4BDHRxwOa+DOkX
doeJ4+9NVdGSvEPGXTKvKReyfd/ND5WNdieSm/rmj3Jzpl7s6Xn7ihCPcLuE
H/cZx69TSjGegVPyoC+r3EWxMBCv3VKmbVWA5l8+iEsEdFCXZxSlINOiP+dA
zLgA01yyTBhL9TZAqLsK0D+oUKCk3ZDrfzHosNkzBQS4SwiSlkmhOOiB2wbx
YpxdpwnMyS16NQ3b0NSyHrui3aX8TBQ/X2+Qjcl1cngZuoqcuHs7g8qleVYR
jgD0doi45QHurXIbMRwgzWQMDlaTlI7BGpkLJMKCS7LvmDwCG3Q2KwUtR0Oo
v0A9RHdcIrHGcdybhmvKqHL0txu6dTWi+wdqQZpxoA8gFpd7EsWXnsQyRrzm
VZpsAGLBFtOjFgVERscflHFmiFYqW/JLxN9i3dIHeph9kcleZGveb2T9cyGQ
kuTTrNvjVXTaMiIcWga7aMoNDbe0b1tHiZsm87Dpbqybv/LaRUogGeGhNNgS
iQuuRpZ5SBzCuBcHdJALTwl8iVFd79t9pdgyuqfzeNAA2EovqacAW1n8358X
EnjMYCbCjGmskxqSC3MQYsOGYIi3KAbhDTS8lwhjE7xZcNs1KM9WfaaP0MOP
WqdC8BQUrpI+A90v9cJ+YQbeP+HR6OP3v3xLK6432+xUoNYfQvyP/23q0VvU
yx5Z0DMy7BzpTlhVlHL3VXPsLnv9A2fdXIa1IsRDFbdFqCu+dY1vT/lSYihz
1B8P/qboEZZGyTzDedjp9QWoX7tfv2gW7zTjBYTrdnI5aPSzQv3TfymjzxAC
+3CGiT3u7T3KWYUVZGGXif2WfvDiIiVWGG9rhxcK6roYeDzjmp4Wkgltn+C1
FO2XGb0/9+khdJLoBJqwPImNqfp0ywUYyzieea3iUHu3EFyVqLU7kS/U6jyy
B1ErIdBtKd7W6xHSLWr3Kn6HRrG8ZFE8/PUW3lgkTMlMOolsn4RkZk/s4JYn
6jJfEcY7nwwdABk4dfgKK+8TCJTTTGLIZReJGNePYya+xV+Ut12W0vOKBoaZ
qJjcjvxqYSbssxN3BTJBME6riywINJN3skmQh6UQ8ZPp+vPGPFHIyT9shwv4
LC0ZYvhZH3s5nwEJsFOFN6yfXu7j4Smd7R4E0ZrUQ3T1QBCGc0jpxQ/Xz+OV
YiIyKeU8FrOHGAXo7rieT8qHffvGuJD7fxT6mImS3n68QcDtfKx8oike07M8
7VzUiARK0wPaYSj+6IhHWMett0LRuTjhJ3v0UqrE953biHHyw7gBX8Q/0SB5
20Qu6zIW5k0OxAlyctg3ieS51T3p8U5q6GsWw6FpfgbxTcsBzj/4OVuda9hd
OzkjWsnJyPDkomOF5jt00tIlMOIQsrUsqJm0QpNag6gJcH1gz974jf3fa+Rw
i3KDxTPu8d0DH4nSK3SDh8MrLv84p9Myowr1XcDuOFO6aDrEdP28fth51B85
2YIU88Yt/EonrwLXDRZI56XoyiRjznKpe57CjgQaQwV7fMGnf9f2mDj1vdiV
sslKGxx1KflsnmFVfbEQ99pwSyKv/xyW5KV3hv2CRAk0Ppmj8suJn48JHNbS
jLPpo6TaZcRKbBhoH7NBDh4C9KBTmqv+bQOrRx48EN7VP2yvZQXwtl3nbRHN
5XPF9lZMEBYtkDzdYgLokVufqMeLIdK73uklI7O7aI36sumNahmU4pG1bXxu
pg41f1afeM24iNxwV4jY7iEGvJ6Kg2zCgO4mp7ZxyRok13PYJULc8gyADvB0
2xAJVQ4mJAK1bX2XksHAQ7ZMDF6JguMBzDQzNq4oR3IlmXFjI8YbIS8ff2Na
mYyMNMNYt6hbBAIJq8RaxA3z+lRogM6tpnxkL2gvPvo2SQ3oEIBLRYWegm4m
Q+RNKGgQvgc3XKlromwznXDVAYQFhuavHCtQi6bPIDeu2MVhWAuiI50BXkai
sAxmouJ4b/6AbsocHXZao7iAkRKqTrEHfAFsdhw2oWA4bQh4yNpp64C+xMeE
/93BnlTPki+HXzSO1M7b0G0OIcKzXI90YK3sxwR33S1MdWDHsFW0ncWf0iZX
/q9VTtoK2HrCQiTpTHjGdforcvvuApMBbIezSc4vahMoIV1AexN5SiS0oEob
goh6wtT8vOnL+JwbwxyP/lsLUIYVydt2yDIuj66uwPHi7bgeWK/Lsq3e3czX
p4UwwPEyGob5xwIu7ksGybmIGuzRBO24O1/i6rb9ZIQM/7ErBHVZP6UEiOGE
biaXihsPGb97IkxZjXsUnfinf9ZVYnWZAuG4mmN5rxaj3UBjPKaWYloXz8YL
1OTtJES6/R9Lkc5R7qS2C3JxuXzcXV01+dN0Rk4irvExA+datFv6Rt0Xd52N
SKfPyz8BOiEOpPSrP7+uhepruiyBxK8jEGNIV6ksO4X03sDSRqlANWSNLdGy
ILi8FxRGZR7wdFSMXO8jYL948SFWTlJ2Yi2iDB+bUZHQyIikhdoOdjOMPU+Z
C4KEOAWi+I6wlDsVWOdMHek6HDJ59A9qsQDP98/ydiYbVqSQSkYowjqNNwW3
xWseHcvanJfXErwAebz3oDVY9fEA60jSwmDGUpStJIY8aiZEUcKjcFG34IcI
yGuuxRIxxaCKx0ZsmUQqKDa/nNaoGdYf0v19dJqtlKn72Ceevqi8zAFJihG8
oJy3KavSeSQ+pH9wOIdLpjDbV7tXzA8gkQWgGRyVAJTMsrU+D+ex26yuap0T
viAnWJcn/TE+Ol0FfB+UgZPYYsywNNV5ZuLJqpCdUJI+pspXKyOEzT5iV4L+
BOEEVMjG5x5jPBIID70bf98drx7tCRAPf9E+WHP3dJP78eL8hqz2S8pcQ8b8
VWMGOpJW5jee56W1AxagZrDkOF2idPhQ05pT1R8LtD5lLboccYFVhHrkQYtl
+2DIiAjzKDrGcHOPotDVyrmBA3kn1hDYo1qL2wk0pF+F6PK3x/hX1v72fsXU
ixofMKqC9wsYJXkHzYPHoOiVRPqjexW69Q/VGwystIPV7Rr7/+Wud/GubbHG
HgdbMwTpKEbSPRGPMqBgGtYio1n6hd3YxOqMvUGuTRzXURZu4lLPud4Be5Ox
+WJgMMoP8dwBoLjTzo/jQjNB8vduRibc5X+lPxjEq8yqQhR9Z//3Va3gQx5H
ES7Yg7qsjwnSaiw0ziMwC/v/Cv28EhMAMDAod6+As9Bx775+LJGz6OG3JN0k
awLz6S+AorQ22WHxR/aasNktjxbeRAjBm4391Juvbnhm3PvCGrc3f5I82moJ
7teaWg5r7foRMoaZBDt9/VCeiKLsy1oFh4JknE2Izj0PNbXtKN3TF7XiuIme
Vb37ZF0FvOwXbomYaHqB5kCa3/QbYEgJj5GjmvpUDHQaAhnXvMKEP36iwO2T
cwR107/M5Lpg7AKudohde/+t1UheqD75wvGTnmMEEXU8lhsmtA1F02Ugiy/d
qcK8uusHMo2ynKQZuUXwxTepEJbdlpo74+QXzsgUGv1r1triC/Y/ZnV/qX0b
jhWov7K3E/NnTLpYONzUBg7Pigh2FlLhUWdTBtlLd7sXN2TDlA8ZV3tgIABO
DDhL2JDRE08Nzb3uMTK2lIGvYTxMbjoeD7SwccHxaX2fo7j5fEAD/xLKxrXi
Vm/YXmkNtmc1V6kQ0ETEgxlBygY+x7Ftk+R6tgGko71s65640kCDr0Xo8umi
sQLqiOYQ/XDJWfh6cEH+YGwJp+aF3UxqS3ecx+rkr5FsgRjVgSHYk6iS3Oyi
D1uuzDFmGsuU/LCAaGL08JWlIAvpQXFnxbLG8sYmP0wf8SoXtcqRddlV2dlI
VlwyUc+Y78cVhaS/xt61MGjQZgPVSAdgx1VDg4gHg4dD/9mgFK2V+Fnt8rrk
eIGE7K/hzHQUrCvinN8lq+zkWyA6iq0mmw4okIUYc/He3XP9rzKt+El+axUG
B1j2dsftQW+H+9gr6rwR33XQwtpcKHs3KLpz9/o71NUuJuo6IloIGkg/RSVw
RS32CDJFngZux0c/o1C87gxUPky1npkK75UZlA+ZV0izfL2BRTWPG/SWiVQ/
MkJrB8e0cnoMV5iehz+bRhW5SttlBX5pAvWwA29OXtVMprqcxYgypCtbEAb0
+NHJnwrfcYBVTOTDvJwuxMDqaZxUzNpd0bQRV4sG3Dj6AFiZ5/YAp1dlaDd8
4krBg/vMV4yWw2lfuKPe6e4KMJTrG9/lpeaYGbtDHoxULFemxeghEz1oSYYF
lbZgl1PzyQ+gZgx/JT0ANowKRta/gzyBzd+OaqEz4/mgHHHKq9s5tezvNcvR
zhCwJqZTa6VBJkxV+NJKHGQ/HSbSGBGtmcdjcaqwhPYmQJ4ayfL0Xng6z5dF
KUxR05B1vtdTPCVL3I/aDDVsl/2rnC1L/p26SnDNaOUNhItudlk0jwaT6CWr
kXQqQ3oUAZDUE/wfjoJHEMJX0jKkXYTpbe9/JvP/T/Qh5r7nNzgK/C5M9dtk
M6z4hfBdAtO+IBwV1N56DKxb9rxpVpDQIs/PgK+7V7U0EOrxN3N2Kg+o4l6S
tvJXyV28bUJiYIOWYdfocE2VJk2kFsp9d/xkkmlre2IPTGdeP3lcKep/lRJ9
c6rh1AQanWzfbWye1N5QHjo0VDYDVr6LLNtdtaj96boU8SH7EX34TTLw8Vl+
injt2dlxviJUAwnJ/5k+3VGb/0pIBmsz9S0jAhv/Pg1kvnKodFPdIUKdaDFu
KYKuy5MEB+EXv+cev8khkLLz3ZA9MuH8L62AAW+mHujmJnN3p6KKYXw4lBaF
sPkZgKnyn2kPJ/3wYUEDgmx1wPPn8I169F8dFvtSAGcxdNO8iOyzQO+52ERH
NJOxj+fJP7vY71roIcOjRNUTTHFuStCJ6o4ml2ygfK+KpUkC22ZGM9nrGxjK
SATETSlktfXRijxyH2ga2PiPSOUxuVXBVl/KFnzAqewjoVnwFINkUBlEaPKd
O29/WQ1qv2Zj6j9G5TRO1ptsXqhdaXiPT/Luy0jJkXmDj3qBFXfz7nzGOB7v
ZLQQhk0EoATN0IKlHHKCspibcfvEJ1chdIMchja/J1y1hzxnFCzwhJsdiuVZ
QD/9ZgBCE8fUkiLSIlCzAlbYoyNKKktbj7jRFV7PP3uQibzQBGNSO5ikSxzW
M8CDciUHV1XZ/pSFq0UYFxjpxNQyn+YN56eHxe/8ZYMo8cxfol6oeI1BzUkC
u6eTJWTVInicBbeqV4Uj3FX5anP99rxWqNMbnKtlO4/psckmhr37RGBv1i7j
pswNP5TPDXooSMCplBG2iBpx2II+Zh1kSyTIA9z3hF1JFl42zxyrXRrsIS8n
Ba28xeUjK+Esuc3ATZDtzmvxo9mcPxMAMqEeikagSgf0L4oypmFxwDeD29Rx
q8Eb8i4Y3cdOTuyRiWRZIw/vx3+eN6cj6FJyxYTJs7OWzLGsDoTAji+momHO
mq1FoU39heDgPIhfwgpwT1vddk/+183zYY91NN4oh1rA+3ryuRiFi7FhZStu
q90tO3yZgvHXQ/oiB8A7rX4s0xFNnK2EiZuKseIi3D7IXNnScEo1hZMEqk9+
keWfIPQoBElAQ8Eu/OAlHIWmTIzVEPNKeMM2m7Hd1mE2KjC8Uxx6JHRc+QAY
8p7OnxqZNXMwAY4UjMTRwDe7UbZlST1TSLAwkve1eggIeL/JB4MjUMjhA7XO
yoi+n2agFiQwCO3hWyWzoInCIX4KTodeeq+yx9dkO89nMGx7OMpK1uFYdJhM
U/rULj0TJRCm+6FcRzHvSvD0siITbySCXMSLrSQ+OL/YdbaBsfSp4D6Rr/fu
cRYUtL8lg9FN+XjiNkfWNW71m8f7Z8LIclBOYGYqM6fzJEVr4kodqwFGc2PI
uaK+vGz88TIvVr27WKZN7PoP24ONyg801GvYAWP5W9ns0hzpeuGlNtsq5KWd
RyJcedKC/4Ibe7I+Uxav1YfLsztZQBL4w5lU5aMQcFyiUDmcGPOt4yzjtFzH
WNZ4AgJ85To/OmSv34vBt/NNX8C0xZg/Zv+yvCCXT3wrUnX0KnrDt6Ksy/zS
8t544ujdzKCMTdT9UiToplPvwYUORVSQ44w/78yu5juy2/kZQFuDFjAyEiaG
uQuobQmRDCVjXHxit99eO6y/d0YpF8+MxNG/9sqeOIsPwKolqnkmHCQ5V4qp
dLIc/KR0Or7SLbLltQZcn6vfxMR2xaxdQ8zVOks+vwwFor2sbpwjoHhTzOYH
X0z2CCETWfa2Ook3RQkufned/h5oUR1XwwGvZQ+ZVLsPyOvAY9tLD1GYdewx
swdNO7XI1fdXFUF7EckqiBve7zRxIz1bK4GN9M0QUkLobNsFV7N/FctceZlW
TAqj5OS/fsYXYmL3t4mZRHLdTaST2qH43aZ2iRn/pfzxqciw8iAbW117oPi2
qlIaIGyqxAH3CrK6DsQdawG22zuU9tJPwjogKgQGhaIQf6CLQOqiosYMt0PP
SJ5ZB8xa2Q2cOLNuL9Y7B17ow6cTIV9tL0wnZ+quF23YEroRMDiOqDVUOGsq
6idb6XteDNOxMuk5DVT06QH4HgFKtwkUgctp83mxxx0JvbYbHkPARGT0nIcL
v1heSsBYWJIMRBUijZyAm3Msn7kpjdKH9TQV7Z0yt1kn6/P7IA7oBln7k37M
CoycgKDR3ZhOTsbyYwm8ZRV04qoI3f46TyYa0JuYreWRDGTXU6pqbZY/7HDi
V5kTZz1Gsz8TR0IjuF46JeDZ8ayxbpYTcccpieEvV82mqqGypWBBhdvlJ6iI
zb8j0MI3IXqgtSNq6DJJVAS5SY+5TEX8VmfRbvt9k7QRLcPiX2uPNLDO/aEy
GyW7HdMIVm3yaIUz71hck+JECOh9gf/3ZRNnyPCjQjJ1VnnfsA+RnoNOz/Rn
LvRm+EcnIYziBHEhljq+yWrsKovjXcqfKlMHRQNcbo1nxz/j33P/s1CIZ/L7
ry2SNHBHmUB+FB0Ng/oTrLv6oQfnz7MGGXUYzf9FoVDQqnuf2IHAFl3dgxIn
p78TrBcqGQJeR5TF+/ecXSRFXfmghBfGnsJ2jJNIFsQDsn8DiJsRwQoSTifx
Q+HHyTC8ShnZpMYwgfMLwr1p8yGRvitX/qRTjwhCfV4GJJ6wKpSTKPh3pv58
wJZ+dzYtwqMPnCOCHKNzUKmj2wGQtNRnGRpkv6kTwFEE3U23AXQ+/8nzPlj2
rOHeI6byaLQWII1Cp392uVYJ7IapP/OucTFXHTJ2utLZETkAUiJyp7H6+AN/
b+qRtTj4X8qaf99j/48dVVdGSoG0LpY2+52wQ1WePKBwWvaafCzAurawEfKZ
8rMfLzUamZGwE/TnWpZxR/io84J2SHPqJHx5QjgZBeuxh4YHRaLuunlIDdpy
6Fw2jfQcMOv5C6UbZhLhvJa7YZU2OXnIvBR589S8PDcPba5VllDXCJKrgTMx
OX34/LX3uvxhJ+8f2QUaMRk7SLn0CMw8D/IDm1M1DUOe14nSNtFWwWa4Y5kf
zvMYakeHoNvfSYB8fuJWUSqmtaSVPulY2KTDuBO1WI4Tkzu4qcQLuaRvg/UA
TFdGtRoUimioht4HH+pWYvJKXHmQXlLWMM+pv/mW3PUlf6rLTLbz6wW/nV7X
YutjMbESsPqzIcsReHgFeWwICwH8sd5/aZcFmr3LxsH+75Clc4wyas33sZ/J
4O626a4cxEykK0l9jaRe35hGuRFpuLLNQ1kRufLALmv7PmtrhKcOOjRETnzg
beqpbbBNa47yFayidAM/Sxn/9lZFURm24DvCCo5CooHSZfkss/8er+BEQfwV
bh5A1Qt0G+miKuAaLa9qeSCMiHWb4B4fe2zB8O/3bBGuFZQy1oEx6wTkzn2E
mx0YX6LLzMt+NQbVfrSGd+QgERXi37/r++4d1xjR+emrwfleps+8wRMgMaib
mu4QwCN37hF58+TXyOLMC2aTT7yYz2kCiphy9JGSFOgqlLF4Wx17DlqmpcbH
qNr15ZDPMTrcetUMb0kfmlzt03tZ1a688NEiFQM2zoflKsj0qBkvpdtaqsUf
kmJx1KX+mbiYbHaZxx5d64HDGNfGccLyZq8jONstniQ1eHh/BvEPyr49+rLt
MqkKAxzm47ugMxx8yB+JGZzSxC4u7RkzvwwrXVNEAgVk5tPYqUxVv+Axvszf
c2Ppge/WZxK1FINHDFKktUbB9Jz1CzjJ3S2xONFH62Za2rjy6gZqhIyN/xTk
qE8b0eUBcG+1NrcN7V7U16fqyaXusGgRBnT8svcVja3NSbJ3gacfvK68qJfu
GaUQVQCm9tyZfWRdjhLqyMslUhCfgp4zmJqRfgHe+9RGQG9fC0bo/65vwBng
V+DVIl1R7Le9zSPJIxT9Cemnk7NBvXin/udcVTAkxXgXOb4Ljlfv+vpkPM3T
nxCdMeKOtZm9DY/c7T+euQBrIN83UN0qRDsW19k5m0bj63A9rQIbPIu8Pfi4
ry7w43x2aTvB3z/WtHIYVxXkEci93ZaX8rpdEv63sloH23i9L25qm8TfsolL
+AzSElPuw1Gdyl9gtPyYQgypX0ak+iaZyu5HzDwwWdX5LCXLG8jHRb92OOq3
SCpD3UhIq3STsSS6oJuvpb5xNjnjzPN01WmGl96L4Zy5Z/7Ty4fM43/3+sUO
eqalYizkQh94uWqnAmgsp1LMUdHLI3lruCEKdzj867i5Q5vgDJqSJ+Is3F+d
qsHKCL2kBV4Gkx6aiIltiMnTifMHa8R2KyAjVjvzyDDjA4XpMvmSzm2QWf1o
03sNzrs/JmkaPLyRO+j5rc7iVfnyWhOjFHY2iHrhSGX8MumDvqR0agQltk8k
zJlXAgNq4LhIfKrodeJJJc7StCTISihcxYTPNC0hVBkAxOB98tissy/pkRjz
DkMq4/+UHJdhtIEL8zO1cJPHJGwPvO1mDvzgrwMGXY8mrohB3GL7uInuSwl1
E9PvvxyoudgeFkosM8RaB5gRfi/VegFdlU3muwjy7A98MBhB0sbxD2Eu3Cg6
1GF4H0z+SVdDPSawKnI33D7cCeBmP301xLjn0lA9+sR9bZwPNgBr1lZZRS42
VTX2rcS07UqlP90GIGxV2UddTyghKCwl9/JKqPeWJAsjNCBL4VxAYoBdQghf
BGYSAH0JgHKiBKewm2d5TDTEYM5RAJ7xcpaRFtv51wo2sILal+DGMDXAaJFO
Aoa0n/IUWA8030mZffeZvQTphVdC5BqmxeYfA6OJi8eKkM7e4Dx4V8ifv+Bv
ghxT603EVWHGGPEcL9hwPNc9nIRIsDk2otEKWywVu9oJfza/EYtmfFPVwSKe
ilmP3wIFcAp5xnBg1EUoB9zg/Oa1hPqwNd0lAeLlkeZvzN04FaeO2Zzyhn/z
TiJBXKiDQSmCbfPLqYz/XEYE/3I6vh/GCyiJhENPQMtm5n6Ahet2tXCYvQmr
XB0w0dzlUXN51CBtoFWvb8MCktwNSWwUP+CIDuYkGGPCH2NnVT2c7vQ//C0f
WoVy47evNWK3HRuF7qa/vSB/Bb4FfMoRAiZvdJTH+dV6gbSG7bKOIJB3PDgt
bbjcCsxUMyspDANab+Q/l4SNKPW+aZNQDON3ym6BS2qC3BKJRRQIsDMLPvFe
oz96VL66PnTNL+u53iJfBbEldoBzAMuLgIRjNkKPMO3ZARBsBIuF2gJxl9IO
jTyH50r7R9JlsNAHHimZl5yMkXqx7bYilsdrMzHwBLVeMkhddzNOuPHgDZ++
7g9/k409URtqKgkHK8OGDvVX/NeKFE5fKT7ejNzNQPoxLecLBgDGFf6PUMuS
vOdCkH5JSmtjOQqMbdeHvSnjlDIQ9BDu7gOEa9fX8ToYoxigxYCgIp95Eap1
q5NiY0BOFSZYrHwBUueuk/yLtbqo0CT1M+SOHt3/slVPrBzK/PBCw27OX6L/
4D/qwzXRZQKq1ZTNw2HWUW+rGHbsct9URmd6OQnvsd8qevW0aYrkEjrQ/I6P
GsFZtyaUeI1uZC/BvaLn8JtQNOtpq2aKIT5BJ7z69JEygkDRv3eZ42HDwiHz
sr7mVpfN7XU0XofhQYRLBWFCEqT+3gbIfEstrQpNF8jfFoLSqBxmb18x7llg
c+qy+O7IYQqgC6f3k/sISrRo1V6rnOBNtnCmie9tcuLu5Qx2HoZgQ7dd3uyl
zQIc9lKjYjPpEgvTyAgwdnyTPBD61jps0YkJdipKkQAWoK9MZNm2+oFrYA98
O4y0tIU1AiSFmXrX0URZOL0Vfj7/8jLjHCdjtSnimPZpbipOV6jnJZ7pWrVS
7HaXJUtLWmxoaBOQ64lMI30S4JPedUZUh2D/+WY7U0tlb1dDw7lSHg8o7+LP
Nuyfw47lkgOoWQFx47zbOCwfx/1SsaODtQBld1w1XMetY56TLt5gIkkc8/ZQ
zTqqyPK9arPeb0fWP1zbCN3sBRPcZDEuMRQjPECHtxoylqQudDky4miswcMt
Owv/9glk7HON4LV2JVdjzV6qthwP3cofOwFzmClI20Q/Uea55alrNxvmZQp5
FJpzUcRUnHXOMyROf/2xbvJpJi4cZsvS0/k9DNpxL8gd2N62Hz1oW4wN7kXe
mRcukd20fweh2AoGYKXx/+d3a/+XKat0urHq5Lbn+1Momp3bUZ16jlVQdUO+
bF1Y36FuGFFF9VaVhDon3auEB1CqpX9wyKw+dntcQX4Z0+m+iFipwzAZkzb+
tM0wOzzJhX3dH5cnZXT1uolbnnR2LfKZL7O9CYo2Y8DoJLTTahuqSat0bgvz
LsE1E+X1LfGz5G3AedPLMIbYiSBTuAuGxyCrwME0FaSzyR4NNmCNHbf+LQSk
FPmVuhzShPHXtXb0y6Dts+BuXEf4592bhIDpa45KYa5Y3ePuesqs9atK0KM8
d+4JSRNZctlUttWgsryvtOz/21DAZk+wREA6qi/xv4vy3n/0ihwK7LHinfJN
BeuOf+STgCmr5AY/0bwhI3OJXm48pTS8hqFb8+Ub/QzHfLxDcFtYOgRDohyt
wireQFYV+ZSbR4u4QqvsEDf+FnykATofqPX8zqFco8SLHVpDXhgRfZvdDZeg
zxmQ2BcEwJ4pAFmonYBaiJd/YXQhzbBbnJGvxpteu7ZDVWq902v+KLKpD5JQ
u9t3EtqpBsFphP+SZUHpyxnFpBaNkIO7oq6sHzNxrpCxrobsQg6341nPU3vU
4gruaS+WyXlV/tt+MHwnr1PAtGuuYczVhUer+mmgZi0CrlY4yEhKRdRbUe7s
/egvo5nx1v0W+kcwlYluD9v11OncMUwwhyQvvq4SsXES4XPf3gIg+eb0rJhg
wxng7YCjG1e+ALwTWDHEybFkZr+xGGO5gzNU0NPZMFkt0pbE4W6qkvcY5ed+
+LUGVKkSDUCHxCET5mXoTUBHSg0720ArkoBMzMhpoFnzQftNhUai7T9zO7u5
UE5Rzke6i68RdV5nHiWzlZOCCD1nAJmVoEMH5BBuFmiMIiUgxfO3nhaLnjOH
xrhX/Io12ShPGz39xDVsJ5tV77eqYEdH6Q0MFD41krPsINnKQtx9cxo12oAF
YIEiNTc3Vf4FwNiKdjFrZ3CnH3bQ/bPyKrUy2PgB5HEM4VC+BrbtRfCB7j1X
m9hYde2rVWuI8npqa6BvKn/3xMhQhwNY/GClZa9OIXGNC8a38NXoiFiu4sM9
4bKbsuE53HqhwBCW6+DmkJTVjM+wpQIqN+K8zBDiRfXPbEqSCXJpvD15ALSZ
4boSHpU9tBgFjSOHN/dTiOhDI1+LdFFuby2OIWIfJFWJRUFTyd0nMriC+yUw
hga4i0NU/NzOxBzboyLkh8fj0PVy3yaMcYrpLB3A2og7QBy1AdllpWGwzO8c
eGpRjY3+xVJa1DBJ/u9orA8edMRhHYu1i8U+cvWka57sotToPPGbApOh9TWV
1LyrNM75NhMYcvNlBZFG0QC8knmUp3/BBP99A8vGRgR67jygpKCXc/44CgNp
vZw7dq7pg5l3D9XSD0mPJF3diYQC76/Benp8koSqnRtRUINMwkI0Sacgd0RX
15BOqmshq+OdvucCLOVsbG/WbbG3BT2Ni/vPUHJlWuHs8urniqQdQgeRfs8Q
MAp6TXZmsMbr8k1rc3pW+2ZYthjQoao5GJunZNKU3wmHwtEqpXjh2l1sKBYw
dKxQqwSvReNCZ5OMf+imS01vBuTWESfeZqPW9z6RqEmRrPaGpWwtsZhgC3Y6
NOkRseoZ0ufNnhNvD18Y6dOWbxOpQ2Psgjcpaw9yWPWqS5xpQjA/FOeWrFEJ
Mj0uuyV/MNkVJVwSoo2qG2rP1/IVqGCG+WcEw1y3jmb7ATTRCZSU0QHfPWTY
2poTd8/XS/lZ9M5tFRxDB2q9gEClleqnbdD4TDZEhBFo9jqxKlGv1PSyb/Oc
y70BMRk7QuF7RvqmleY+cpcbI0BDrx/iIPumr7wDrvSVvl7jpEF44SdDAvMZ
vR3CtlzBP2qsHS+QSqWPlhLgKHTgb4RRuG0jtv7/Z0g6yRcy/8WOL5b7luOf
S3aUMVUNc2A5MCSR8QPAL+7PlflldoioFgyyoo0oSF2PwB1VOO4D0bxVly/h
mugdonX08vWnUTjdZUg/ziHzmiT4E4Hf4092Dudw6d9NuA9CtlDvnQO66qBq
emqPqGxPAa29Ro1LMhcZpezN7OJdCU/WWViLtMklT3Ka4CTcAoqQaMBYyYrd
0Xxrp+0xc4YC/rSCDuT7csCmnqFOsPbXMo2ojUHpHeYQGxq79Sog29U3bDAf
gFFltg1c8SB4JTqGq0lsRVGoB9MdxaFh2canCZLOALMj2avaLK9AIcWCJTt2
IyLWbMrS1TWElcznofvXLY6hwN2byJ3BatEJ80CG2/XGlV9TOQioBENL5t2N
yh79F3IfbxueVitVT6fGvJPzEgkB2uEhCBMqg2IcdQgGQMvfdJDzh3r5b+t0
xEbmJ8ajtNFInmY5BtIuR+wrGHko/V5sCGAR/izUZ3uuZ80APO5+cppNT3Iu
uJUytmVAK/6dOVx4fpALCnE73KXwimCOoCWCrRIBV8skMIcTVWvposUp5AJy
GMVspuXbBXcOYXsz6EkvyQph/CmhpbC5HAELl+mJIjeEkDvn7iQHNPGIaa5a
cBnJ0dHFDDNyjqq/ePqjpfkGZgoH6ceBaJETydJgBMfQBcbB0CI4O5SN4Z5C
PiJY60Cwa+ZDcTatHtCCrLL4njtjjdJj+w03fBwDm8+OlAgRWlfuhBdx+Csz
mvrDbk84kBel/x4eGKBGYruNoojCG7fHgGF70qILGzdvh7Zf8RWATD5Haj+C
YK6tS6W9mylZ3aUvBLsJN5IyklgakfQ8DRxN6YWaMGkxp+v2dVJeoTLR772r
b1Y7KclU0eFeBHxXpqXnKgXX9YoDU01ldrKK5rWT51zvdtBqSxkKafAIS2zu
8sQvdfKhnQh0e/sLglcThFvfyJcpjXoxmwbiudhSiSUXbIY02Mgb3bMsr0XZ
6Jl5jdSK6BWEI2xxeP+AED53EoIz0Wt/oon4cYkHKcrzUTHTcMMqAdONCdfo
SYuEwo/BR2Dwil0VaWWBelwdw4isx75tqYTfZs64lHwvmjMfQSIVdV6JRdDl
FFXgA2lCxrTfU7XYZqz+OkCOQvu9wV1Oj5o9UUoVNNaq3TOJFiLExexXSGOH
FalWKHfGQZUr1nMQHqY4cXzWOV+9P21Sdkhe05m28wLigHLBHYzj6Tj8VOv7
pwHBhddYQZNpxNFF+/KsPpX6aqYN/2cSFDE6DAxymq/DNXLjmyK8EqbhP1EP
UzL6ppckmW2UMPgl1xk3wtjN50RCQW7Ns4hDkipvLiv4kGcRH8WwJrbSN7hC
M53Ijl7qn80mPCJkXLvOPj2OIC9XEa0wvfpZGRKiT9CVTHjN+4QXMeiNn6bk
VmPHVcluQxKiK8giE2wgNaWIKfD4L0xO5H7FaEVESd30u/Ivfu5thhPw0DOM
56oxlmauJ0yV03uymzvCzXzWRFBZoy9Z0wIq0zylwwvR7MFxKDMpqwKQ7/Gy
kmCpPiTFdD17mmT7CZUMJ3N98h6Z5TbO0Hy7rG3BNSP3I6NdRmwcHtI8oCpb
Pn/eUhQUT+Ia/C+7MDJyrAbcAoYCyWOeBkRUT75ZwZXBLH9NfEojuMWD/C9i
5iV0rF6c687FtUQPFI5YvS3mZSqNSP8y+mEqPiExCzqZ5jujK0j1UUzin72u
eSlWZqj8wnX+FyO9IqsIY0b8+1TnI+da2TNX0Lw9YAgL8gerHwNf9W2/fnlE
8qAy+TQkYar8MJOyulhbz0WoT/WwVZ/AAl+MD82wNjEFa2WiTtUuE0quutj4
uiuwHArTq31Qn1e4g0ne+qZhzIKyQOlyVGpTeeybb3MJ+DUPsqcnlQnsQI4L
p44d9Rc3xlmhdVvIr7TXwekkJBR6XVlcQ4r3ES1wDoOP0BZIT8NAeyPwHCHy
KzO7GCI7m1qZKCgx+cA4VSLws4w358VFV5cLh6xPg/p7EGrI/HMfjylX8nmN
50Xmh5yzUAPOuX3vN7ChoQLFLFA4O+ilxRg2rN9J4ifyZ9j8vcjStHuSYg7W
DiCJsscwj6fNBbwUImT+DNl5n6GzyVSPUJnffL+SjptnSf8a+Ca/YMNEn254
K0+Rl+c+b2w5movZXDBqFH21nDUop2vEB5xAB7oa8T8EdWZeIAdGfiqXlFZF
iuGmuE/+WhJTJ3dL+GXnx0F4Mb4HZrrYc8j+vyonnCIGmHzYEoOio/R+11bm
YXvpXDlW6DWYm2m2mUsTvBt+xd1h6heKRRq4WEp66FQ4LD1IeaTdHnKprW/7
jQ8lTD14P3knyiVBlQTtsLBeXqqBbvOO7ipP6FlGEPgDjEoi4OgSq5kpj7sV
8q2FZh3ukfv30U1uEOCa8k3lHs67ouyCCCEaTFha1FXP8C4IVU8FPPRUEV4c
xWjfjIvT+XMDppK/GeMGNJ0+rjfnrFVve+hXc/KIcxOK5G7fErkEOjoG3HLh
DcOpCDUyHtpY74l7HCJM3LwutfgyaP74X+yqXncnn6FqlkgjprWJWnEoiGGr
ydAXDYZ3EmXL1NjCSmXNl9dmglv66rtfodOj4PL6wWa3+aYNtsjve+pGZi2t
M+7peDpXMXUUlC3C++3eKb4Cxa5u8AGBWxFESB6OEeTP5B/HKrBnuqVhb/Ym
F/VsAuM49eNbeIEX6ghAm1j0aWTV70q+AXFS7cQ5meuuLpQdVDKpKLhgPm1A
Z2A8oL4UsGPop+fa/B3z4N62XdnROj8f1lpKNnHbjleIzwQg05sY3lfE1M+k
BjaLOu30NZC0R6zIf0sE0xTFWGXEjh80b7wGbLT7HzUvUaQQwAWuFyDKboXh
6SKg2huubvBeo2I3Wn4M9w54VlPbwQQ3mvQvyHm5bwcv0xN1pttVt7Ygv8WF
Dr4fU4hg8Jn35/fTmNiFsI4bowuCckuNCsUL19Bcd76WDuAGQK6sYSpNkn7a
kgqd/QaZRB4YjoefCLykDuMop4+X1bb9A6jzO3QIO91GkNAJwyCopFSeYjln
wn9wZZZXUfLY0kWCyikSYXpwr3QH8Ie2LdPXpntUdsaDYg6Z3rsONxl/PLot
H1zfgZznEevvsGsKUJCVisKqkTsFaDoGRqiMO3Of8Obz+1m2FO8asNJPBAcM
13Hoo8X4mkx7ggiUEyNQMV1fUFWxChH+3Bnde7fVXBq+rGosmR8Cy2mWs4UD
jZNC4hLUTA448GcASPpfjIv1onfc9gjp2eEyufgv3IU27qidBHNmi2cbdqmm
NwM7fLE7te1FliMuOlfoX6cIHDnwwEYAfgncZkYWZ/c8RYKEo8lzPkmtf89w
w7JthqrHwNW2Eid6sdcyZHcbYjdSchLKcp+XnUC8PpFIKGx7Vx8JxLgp8VCM
74MBJNdt9R5/NknS1Y4SapH+rwY5Xvy3Q/SoDrAN0G1mMag6qRxG5Whw2erQ
+eqjowmdd+OW0ohR23H9wYqiKobCJHgcYACuYN4D4FLT6yOkbuNsuNp7FIQb
ouUSuJQ36sSG3wguTx02lVlBt98Kb9/y81RbhLhbMbFY/CO47eDhR6Lotd3R
MWk4oHrkSl5ABE/s83D5kV9h7CJamn4Al2j9khkcapmwYERUq/pYnsdESxGx
ZjL/SPLdgSToVqnIv5iYlE+e7RCac47WDm8C8RLMnVnT5l3oP5e82O+jtuFb
wMh7XYx2nOgXMStxOsAXiJgcyvdAr626FX+r4LXKYWCo+Js060aXR3O9U35B
/uhg6FZ5cRwc9A1lqwpftLR39+lw+Z92j/SZBm4ZdUJLuv3DxeCCigHCjoCK
XOh3P/FJW4wzU5Z6JouljDljDDgCv3jxmtFFPoyzJFDgcVEHN5yKLxICt3IR
rRW9VqS9weap5TwEquxpdMj7yr+I+RaCBoAaXCZDEZfK7xc9p0v5O/CMYvhv
43qkAx09A3Wzyvzb7AIK92X37bq+uHZnYPl0mOLg8sgMBYiTx8HUYogABmwb
FZLlPBreBj1e3fazCY7Ly+Rxd+ZIFAwLdWO9pfXbItkjKxJoGqkHk2bXYDt9
JvC9GB7rii0NWY+oddMbDX5tD1HV8+3JT6tciKhjOG+g+9sV0MY+Rgstq1IU
XCdoQyySWxtW5BuK1BgAe9e0ZKbLJ6Nni1s5Z1+45RLvD/W6G1geBsyoAG9C
3qLvYocrv29fQCUnDJQJ4LOYHD+T31GF8zF0M4NHZfmo4LTpJmkyDL8yYpzI
joBe0yjgq/VbhIIDt4F6nVjyktkOnYMnyjUlhLZs9zVp4t1mw8GJ0aoPA1Kn
gumfbxFVz6zJuhi1Dmc1rVGW0xjeHzyX9NmFZQdXf3KxTfYgT5jH0BxAfkjj
ordRLlrpv5DDXYlhb+TyeKvT7HCWDdrhve90IbeDKBRD18/M7fPJ476DPTlE
BWmj7UmVSXxprlq7JL2uBWBh2JYBDaMIL2C0SxjOpGi6Ol0gJW5hfUlj+ZXL
+owRIlVI5f4QSfLTVTcdhPLmT2nex3t2o3w2d7SKD5cZAjvERp956strIa4U
xs8yemo61V8xfSoyspItmZjVOJEmIxYTGBpK1Qjm9/kmUMxaAzR5hQ81i0NH
qy4hphUmecOftIOZ1nWhMaWtFLPJ2oZQhOoMjHePmzISVHS74vW2tgoMwKqR
ZBHmsLQCyPTEfMU9b+nwF2Q2STY4294s1lnK8zQXFR/jGLRMV0PHrQGc3/JF
wqMYKn1gokM6hfEKmTb3HdQeoBEN0hmlUE1jLjMIDmWadglQmx0MTXMyGK5v
SvIpGh8oMCU1tASqiX+tSphZkyaj1CskGSANMbnwQIipgYep6DduyUNyFd/7
dBQKDIMrcxcdCYXqq6JymgClp9xCK6tFSL9f8AlSL4g5a6iB9LMmNjP+SqQi
VOilkYImoNgH5RapRjgoxEJ7funIeU016pPYph5wjLRbgQBdShjTrmvBomSC
3a3b/Dz+JshnB2Mv5zlDPeKNIHGGh7aEkbbUkH8a9/66f5ep8CHKxJN8neKZ
eHoeiS8fWf8PHqVg5rGhmveZ3QJ0UkdKSR3e3M1HgF1DlGbp/uPUM3+ghwxm
dvGP6eEQS76SQgPrSs+7wpTt3kWKkV+tH4CwvkyKhlBlG7EbNI0inuZBncRW
MtAVp5p34Gw0S5gkwsLk7nzKEDR4Z7ceT/oxAHrriBD0Ja3xJYbY5yP8f13a
VsPc4RhZ9lYU38q6r2evuYzTIsAtOgSVhXX5iSggo+HrTVCe6zKymKbNoC3t
HvNY+8Yclp2g6i976Z5K0rP4nb8fblSQsFnTlHccj4Zf1EBIdEpcGhRZLBht
5+1JFJX04syuJaxHTJq84EaAhzrTFgZVyyD1clen79eDb/wS1ibG3uAZYda5
Ne7yt4UATXlOT8BBjd2zz2pLLs3Uisku1tUlOKOJ32DcQ7dvUEWPFZ4EMEwO
q12LutyeiwADFYjHIddNaBuOjzN7n/v1eW+Nj+V/NuCI5RzppZ93cH0vvQWJ
anD9+yX+gk7szRxfCDxlScD/FJj1J9mKBFmqsFZjGCr0d3iHF52In3x9Duh6
zvoNH9qLmS6efWLzIlotiPcqvoAwuDcPSsl8u/f2LlK5s328FDuKpMuGJUKH
fcX8HkA1GUDvQb7v+YUKtCmIJuYwKEkgl/iZsk6hwBx4hvaVHVBQx+WUpXuj
VKOe7jixw9uwDr8SPBIhK9bhS701woEqGoJ97TeTN7X1lrRoIsGx+nxDMeaF
3Kfl55BAV+UuLRboFw+4AkR2EVpUkygKKb4SbKzIT8zwWR5H7IlfBW1F/weX
QyxkkDdiwTKRtwEz+IlVXe/JySXwrcPGpoLjCgT8k1lwbX2rwDOeQkvqx3ly
9xEpB+gqeuiHPkul55nq3C8+/VbGtUqfDTr6+GNzKvst148SPHFezmBERLEw
yGOrnrYLmHXo61c+pxwwDd91t89xAX0/gETVuOpnp3Jv8hCVyRllnMS4JYoL
CV6axYvJUsSCY2xwCrjjbSXbDpNAUSVaQSph/ppyd9Qhdqnx6BvyHZM/UXk2
XUBlM4C1+s/rBwl5lHCg8+m8YnsIrXKBOaxQrVxppTPyJ3rKmEHE+EW+AG0I
BCqS4Qg/XjlfkHuJ5pAnJrsfIgAGGBIAZdIr47IMvQOswtkYr6c7sicRL1Oc
AXfw4rVPUfRQjyuDnnqVrmqbkeEx/FYTODuqXZj0SpnIg9wXXJc64mse9gOl
GKmeWc3l/vJ46fazqRCgggVGnRSlrR1lSt6NVkKhANsEeZs8jDTE8kb5XczH
Cs50eo59yLfu7yBPhPHXw1wDTWJYXiEgAldVH2j8yTIixVImJPnSY8dBUDEJ
IVIo1oLFrrTo/OJu5rk350mLC2vWwVwDELZ4LRW3LWr4L4g8Molnfz75SYLT
f4ryV9MhxTG/EHaZlqkrLf9JhWLVkqK3XoxItirlYSJj70uMfm85Up4NK4GW
QC/zLd+J7lcUYFMJ4jTJ+6BaBfshe7VcE8i378e/ExxrqU1YQmb9CrvlXpyB
MzPHDlRxb+rAj2IoJBNI7FVaIXWSWBiwbVtdHzqq9OC4nZ4FIEsul+FhvljI
0OdAPDqxzfIS39igsAY3sR5np7w3lNg05Tw+IT5uxauYAXHbmAsgHGAU9ZU3
fyZ6sfQ4wtVZjTfjDwoeXx+HHdOoAw2oW/GaP/cUdpat4Iud2e0j9CaN/e3B
y8DZcLNnwtQ2ctdiqdf9vxEPscxPTxzNzjLeeFE8hldJnwk5jMNZCr54Qckj
DL65zbfBJykil/3G0yqTYQcQN8k4YL4BWz2MujLN0lPoPrpBWkpByfcO/dp4
6Q1zLn9aKKfGuOD4bmpM39+SA7x7mFX6WL0+ylFhgY3Yk0KwXaDji9RVL/jR
VrjKpNpAhQB+IrEETY/MJS83aGcIvWFJn8LS9FaHfo1ayuJDQ/cLtC55kK3V
LpOlzObwNJAOahcrLaEVWL4CmC2HMu9dfQIINgSFOvOIdlTUihVYolgVI0m4
eupLJHDk5U6tgNe4/+Ns+8ZOZ5UslZrSLHxkJO5ySVTTvYfRwvrjoPbXJHht
cm11C8nTJjXjOF/nvZiIERV5HuzUELyxE8ZHGGKEVNdbmR+KNkHZ+g/TqrId
YjcaMj0KR/JBtW1OE/ycdpqblS4aqvhAo70hkmAKfEHd68WbgeLpt/v1kcW2
Y5Te+okjtbF1e5wytEynp1JV2IOQv1lWoc/AfaWd83d7phC3uIKWD8yaxqNv
Btl6jk09KIooU8t4T742U7H3gYpWy9R8poFu+jwwhJaZS7h8caCWBAR4hmB1
kSQKcorNnfQVu8qBeOVJCDyArGzDgaLq40ZJ4vk8A7vmzh07/907fZpW31fB
l5m2eQ4RZBpxDNzn1XCEhY8Bay7+5pMR/z2/izduOoVkGCwVz2/LpnF0AOGj
2StGMm+SZPLfRl+G/Gv8XJjLPoL/UTJHZnIOB3cbGoj8mN2Cf0CehV1w3TRp
T0OH8pd+Da0Z9UWp1F1WWF8+rki80kxEiFn8dslfoMDs7Ac8TrtVXWXrkEO1
Z4aTSzLWN59/QmOVzmiw+dMkspNFmKwXm0EhKwdZ2Y6AhPwPhZ93JH69BqvN
3ikP5iN2Q13A1wocOXo44CYJLMeTjVVokXRYkUtpF+syGPyazltywgWdaarL
00+PEu6EG2m+HdJiAqlNrv0n0cNx2MyCMZd5B2IOWKy0TGI0DpmA88rrlBwH
qAD/ScTGc5/2CkRJ02FJ0w4FP1VgeFXC2QUbKi/g7oU8xAupwYg0G8OSDw5X
3qpRIjMgalwaPklWvcBtcL0PxPfGM6LRrdcIBeVoSEJLyqkLqFxUYT7e5MTb
zuOIGYym+3gZc8QnpHBBDLeBmQQd2hzwBGqJPwK+9aHonWgf5rS16UAuMdIs
TznHYeL2STYYwST/EsihU9Ip26wa+2sMxYpBWesuUSqiwU1LrysX2mr3SDtK
J+7QVQZCehN8x9Bq5pTcOX9wd5Qp19Vb/XLBNv3WthgJI+M+FmwTG4g/O8nF
CpvbaJ/DS6fEuIZYyyJOBD85pkCLTDx4lsdFpzV55inlGo11JNqnGO63FN41
S9RGctUaSLgdsCDbSG+hIz3R90eklI/k1hgLq06hoq4Sq2V4PMbYS57NfV/B
xNgpJ5vhnSf0cqFn74qhp+t4BUBKocUXd7Fr/M4YRyakZ+S8KFryHU7RBO6U
5tq/U1D0t+1h3hrAule84DVU9DxMb17wjoFQ70z8ZszS0dAbYLyEao1LQbmk
MaiVGnthIVFupa8rnWvyzPiGvifuzEnGrVzy/OZhC6habyug/YoWy+gtIN4/
r/mmc4XmA8s3gHfFUv7GtbXytJAdLyZtNxSiziYzdmh82k0HMMbkCWA6I9PC
AHTZw2zkAtAKe84THMWkgYgzFMgF1sjRFw20UYcmrt9OPJhm2AxsrDBFs4TL
wcSKERuihn7AZ42eklVfqR6AFHLQ71nO+RU+9riK7/vXAJ8d+aJLYSQ22zo5
UA5PVbZXfaShahyrRdzGZ45a0AKKzNTVEFp7upBRGDbu/EEc5Nvg75QOrXhE
7fv8gt82v7yDh1GBAm2UUHU7pPRPm8Oa4J/r7FslWOCt1PQ1LTv58AaYeGGQ
LRN51Wd2iPv+GZyW7F3QijkJZXMnMeDcTy0WuZjoRAXVsxmjOzFfHS+8JK4X
B4Gl0TbubHv0nhh8iaDPbRo29C9Ul23HIzEmWGHfKhJSPT/iRUmPh4tl6iE0
dAnPKSD97RP52eXz5ZKRcJf2pCerz0tASkNpE1BQNz2w1pCN1w6BkoMJIKKe
uE5eyehv7eN40iz4zbfP9agp2X2f1nETgQGPAYRLwL7IMFON3G8ZldUUmbWM
E2Eacj9+F20buUPSqpxj9n4JSyqGeM7SWK4ICfzKW/55rXZItRXoQCzTCki8
yaVQFHzi+P8phAuGwBSCD+c1BY/g7NSCNSWF7kT2ptwOJCIJq+9NVMRXOMcY
wWZMEveAI/POx+z2+YJZ6e2LFVZrluq/i5A6WCW+W3G0RCypvIBJj3u4DOHc
vjcUtd6evSo68BJlc7aH9DVrTClwUnWU5p8HE7oYx1afMCkbM31icqsmzPt+
PF2e9z09B1fpgfr4bOuES3jwHmbgqEtlR4XaFm7kNWn2Oo0d+wjrcSsk0Iaa
UgY8Hg0nieVPnAb2nRYp0v4uP4RUPmMJ4/CAqP9byMoqFqBJI8P8HmnMnLiv
hkbvJiXd5V9b+LUJRL5n2ARsGXpxgxpnw3RBreHHadmCERKfaBOZFo1CgPbH
okZK2zQB6gb0j9uEOKERIv+nW6p0bGyVWSfmy6pqtOjsRFVhvqUXjKC6HEBd
JOaETWES/FK3LA2sJUDIWlnSD8YuHpPqBUTwbQ0LZh+NgZ/r/o038a98WXGY
2Naatt49w1YirtN1ABqbHD3H+PBmfe+TDioF0LtA02kXhU32nhZfdr6NU97h
NahDfTcwiroPs0khUV3rtuoOixEhtbvhc9x8q18DUhy6CrvYfNaxJ7k7K04a
Kc2Bi+JF5RXtvNMV7jXWg5vIrU97hxhn6/vYNskN4HyznHdHERw99ZjVdR5e
xIePdi1qAEXUb3ia2od3Lqd3J0sXfdMJER05sP8/xRbBj3K+YQ+iEndxR7cz
b1BFqOIlEW5ANHTRPq8GfMsjwRCP1cdg4EfiTDP159eG/CXHyUKEuHAuC7bH
dhkO8Nxe7AKR0HSGvAZ2bKwSrt6RGKu+lMwKd6Lb3/XyQEa5agYRkPPKs+93
uJKTLwmnrylQlZuW4AlBs8QEljmr/o4hnMei7eXIscnM/q5dQEmPCRbYNRV+
lOvQZy5oo4xPpQ3tDNd7YsLr1nLckiEP5V3T8ykfm3tx1/HDCd97LfjEaDzV
0qsa/8ZnAFPSTLK94B/UGq7Faen1grVMCMkHaOxHfFmR2Ygl0e9DfPEbGzkG
ZuDJL+q3vF96XgrjMwjXR5217ErGL1yMZVe8S37A5KBQpTjmhGXKXD7smshL
/NmrRQT5B8ml9mdwZOZNAJUIJl2WZUTwYjjZvxOIotETE+Ra+g86rT61i1Yx
CRYNOpY4j3t2kophz0hdze0IMFsaJmDwUBKWXmUCYN4mXt9OX2aYWRN9xLid
z4jmNJG1MKcJCw70aeQQcmIj17Iv0bKVBkw1VH7OiQgy2HAaFGL8UDeG7vtB
4VuJfbxvjIfo3b/5xU4uayMI4r586m1qAqMgVaWWRtAyzEicrUSyObvtsaCV
WWNhjnsD0G6U0IEQIRdYnuulUsyhn/6mjbJf9QbvJH8j+9n54dFbsHPmauVT
0t5rMcdwevE/1aaw8u/Eg+k4JmQELZyGC3Nh6ZN/MU1kS8cDj2zCK391rdEG
UY8ocUnbHV7dX/5I4sIdigheudcP2ZATzPqqv6Tn3AY164TrF5RkHVZeIxOx
o+7cZSrIGdaHwJKMgxZW01B6O1+uJrDjR0QC4jVu0/KQI9W/1mEuHaWCJ57S
49ycNyKdTXBzSiz0h8Bx0+hZIe/I1i/EUieXYdJd4jerojZOqbDXgBNdGa2U
HOeEOSkhuQPdJP7J3VTUdP1Gh/Q1MJKEHSZcCorl1YnCPga6kFgiqORSB6cd
nC9leJznW5GZ2LPutOyGSEvYwEL4TihMkFhp7AG7kGq6+UmCS1ivyKi3zMxa
fhd4ouWN8g/2xRuKHFX9PwXdBOYuKmgBJkLMk2u4GeOey3kZPK/sPg39clD4
Xnkc7F9eO6eM6bYa+SbVyXBaBIL0G9t7Ja1bLTbYqmFehOBadJnU+bhSNndq
fyLL7qoovpZXAbCSY8qXRdgSSi3Ou7Z0YvJdV0BH8xxcuOMCD3gA46a4GbsW
roJ/xI1VFUBdaJLPYUWhX6EoCNg5ot4fscQS5dR9wG6FFdRpYH2n3oiSv+Nh
pRvC/bnWkyHqNaaRXrhFngTWbmDyElVXF9T0CqE7/V4LC12JIq3gavVGJwGC
6DzEp3uyfv+JiAzf84vggCt7JMJ9vOkFANTF3VK5gQrC8KIzz3sespuL6W9+
1SQcnItx5IgZX8b9olfYImVoD/6Kx0JURL/esl2xZqSRj05qJKKE73T5i9ER
odlKbW7g9FD1P5SopAKU0nxBQTc3i2x35mbFr///zVHp/5gdznT6hjvO08yV
A2KIecvm4e0wl+xKoHCCM6MSVfpZFVN8sAX+Uu1AqR9riernG4MrnYRjut2C
qsuoWesZ9WSH2i1x8qQM+YLhlJzZCqY63kCeSINKN0/iyXXCxAjtY5GjphQO
buspxsLGHzUuW5XoDKE5bHfeobFQzNj2tq7tLy/UNRXWdXJ1eTOEaGyWfVzI
tAUvm23Bs+q1KZg3wpv6XvYtAHygwtjDc8Xo8dY4ADyirkVnUxsLDStAYs/m
1hVJ4DhPIYlm5/61abpC861FsqHCMLC2Y5qwky5uKOsZ9cbobZGqyqQzXQMn
LRpUhRUzRTaW0J3IfX8i6+ra9E9GES5Fj+PNRMBa7GGYrxVEElGwUVkYOJwJ
s9h5ARck8y1tXrpybSbGfo9efLSiSu0smOmB+09HQBDfU5ybXoNziUZZ2T99
W1dIvT/cDrA5sWeDJj5EasPhFZzfSyKCILQ0kcofE51lWZf2uaO/M1z+7KUx
0DjulOvkQOEVv8DO4836m4xrcccLJ2PzmxHVckimss84ROwHlKw5FI47guZB
hcbeDUmr2q+ko0IhmZx2PZsD5F9Nxdod0hTH8yTG+PodvY2bx/zIxlCFOAwE
S8KH+kGCKQewmBr03uAcSM6TiZuPws3ZdrYds6213qtoXJ+rZm66LjjtcGkl
bwI9fxPuRzQJRhdN4mAN0Gy/VRlD4r+vtgTU4G7AT2CllRK3onMLcBfzYlxV
4h/8obcB0ACg+Me8/Tx5obKnJMxgtQgVk+9axoXuX42kB0P6ccf1DuU705JN
Nz+t7n65to+kU0VF4VpJpKPdS2iP46vy7EWauOiBY28vyO/UpLxJP95LfeB3
5tvPIo4FJzT61Zvq/Vxc9kt8HL9DM++awUctmQ1IXNT/GiyeFUtO9ByUHvYu
egcLcNOImsh6FRdREdDg+V0FMm1WNcSAOyrLUv5Vl2rw1Ez/Z5ZOliXajq/d
CEA4VLe/sQCV9B9ysPLMFmlJLQSWgglLyPBf7xn05pcu9T5WQx6QViNtihJx
HBEXG72UhwpzQ8d5ejAA0a/tNrjxfrsHfgnKohjUNvmJLqE+Fd7QaJ/oy8m3
2MfTSDibId8Eqiq925PiEzx4I7PdlqvYyt/PzoLWhIHfNHUPZbPqWvgaLxgY
bqYk6KEPSInuN2kr3GTltljvvIUqguPP0QTUk88bh0j1R7yb/v2mWcbUtd7s
sjTNPKUl0j4wiHwGvO2disYSEcG7pe/AW3idN6AvZKksyxkXAUZAhZUxtrLp
ZH0z6cF7V9/QIwgzWBJTuzmEGrec4CrgGheNblpkxRBViYEyaDED5BCAj3Po
pwrgEUyN9WDcRkPgKS+ONx22MN9Q6CBsNcHN4Hwx6q7X2g92MsAorluVGuhp
oI/h6xBiQ8dwetd01q5eWFCDxbVCtQDXoLjoqby904ivD5xuE489HmeCqJVP
3gRPw4JYZGVG6OLmcnTHgt9gBus1AVmQLyRh2VV+7f5aQtsUgihcIjOEPF6M
LvWCXcRLlCgQsIa79mJ+LqggE0qnSDYFaFXoEHkmJDjf+rvpPQXsqSHN+eir
MwJZN8p86dVCCiLuLw1kqToLmBC1QJLwuoETrR7r6PZ2YW6OPZueYDTQj7LQ
4mniSv938oGehjA8xZFp6p97/39ySylIjRsAnVzBW40VM9d7yzrQuZcT7qDp
q6tP/XFbgetrl50/uM7er9MtDQj3yhAISZxXhRx3sc3pYCxia8Xzbe0udb8E
DNKHgf7nqN36XU+QpI4y0ZEPziX0Jz1ml/YO2HaBzfgtfZtwktxPHProunFk
2Dyz3Ru0R8DjJz4ZFtKszNg3fhe2upmduwmaCgPwveSVkdZzaH911ZjCcgmI
Ii+xJbwGZllvGWsGn+F+MsK7jdGnsg3gTQMLc06QoR9TjZHWbBie4tYl0ZSB
NF/gnWWr179Kqr4jYpf2kM+4MZPflHUcrFfWBP4erIzGnM88wjVaXm0kbCGL
byl3F5rpImtJWHzwvYs5rs1l+5WxE3V3S8O4HQ5CbqcK7UbIMcfTfO6aAgKy
7qzM7LGNQQxmxmPGNhd+bs+7ez796pxZiAC2uk/M6PmFCm4PkG2BQZKXaIsn
EOYIlOBGglUR/6ghbD788He0U96NABzS7JV73BwyjHfjna/3naz8kE3pQU3h
Jma2sGA8Wu5ly/M80WMcXlVOksP/07cuoEsZVmvMkWmCMSYZbP7v840lnhlr
XPCJY+EtDiZQgQGVKOfWJdRsg6ghhfAehPAeCqNjbGFw0ORDY2Gbe98o4E+r
3iODaLp5wa1sV1KIPiSNiZRnbnbqhzDjxc8LHoNOxNTo9uwNUHwDPk6oj+zC
Wd09x/1qnX5WMbY4DBhx+mKO1szvnWZ7QO+RjcXRVc5GSCJbqHt8oGrZ31m0
+LpRyWu/fZlJyOsJzPZyGkEtg5smOloJrPg7Rj3eMPVYb+kClCAJEhsmOncH
4dodlp3bxkZyeWlVpiDpSzdRrQzbYTgi0JZ4TK+Bkrcj0Mw4Z8lTNbXXWOzQ
NzM4c1yWjAwX6A7czpotvy0aihQKizBCLEgusybpZSfHa4rYMnt960Iba9OF
SKJlQwRy3mqrdpIO52pOoG0LhLH0Sw6qsAWp0foRKgS/DaOmVQoY5Eb8OrBG
kicSYQ7X6LGFVuMRE+NARZxTUdlCeaWX2Pa6zVTR/jvNGJITZ+XUa+Xr32Ha
B/gjs6xqKPha0RggINB6d1x5ksDTQVFVJ1NTZKV88dOXkV5umNKk9+ulofbm
48plwycRM0stgPRcbapQGaebJlEsl0cu+Z2C2IR30Z+uo6pYnSfrbAudqg6G
XZBQQrlJwG+79DNCsosVKs1XkajuIlxNn9sfvXZIGgxMvSyZ1TQ3DrHqtDkF
dCtdP0BLsE5Hm+2ib3GTBIb/TK1huIvPkQ+11v08vm8TrSHPP3t8ZHcZb0ir
mro5ydlB/brPdJrlHFxIUe0M2loXmlkDEtsaTMXhfXnKqySSIFs3Y4MI7xaM
XwP4KCUOOENqXZT5qHNpYwDYDQB+XkYU3yUfadPKwHj13o17FNL53oQAjZ4r
J0z/mzCZaDvDmOnMRWXTACTZaFsm6K4QNOVv9CLK6oWDfXIQH3aZNGSShAXP
7QR4Tt9KKHFxKC74u6SOnZoYvJnOHyPBgn9Y56Gef83qqaI5zVfx+TJXnKVn
ncrYJihRs0Mes93gcLxPswNofhi8jfOR5cjTN1MCd8L/4/b3ui1la/x4eM55
QWx3bULuknH5UxAjhVlwlBbIz/zT/HfZ14G0V0bAGOdomg2et7cHezAoBvZr
PXMZ4MDjGxFCdhjhLv6RWBDw8q625GQ8/kpUimNJd3k06HgIyROn15yVEAtK
fqopUdun8hMqzKaCkSBObQFwomA/RGSKMKwJv4TdEUGBd0XGt/bP5sIBl9Yq
8CnpDvxxOLewp+kOBz+VgnegOaQ6JgUkWV/VN1HwW5d2ZgtRK/7aZ42b7KQM
MbYNOD2JMnWkNhfJVkpNWXeBvvtLGIvtp/LcrHta+McM0UWI8pXL0bY1ftKJ
2g2MBjLVy6a1c/cT4m8CYuZrre519cUrrQeKebZSgw9POlGPPR0EExNffj8e
kvBTF5IRso/7Qw0WKCoruxXjdom4uud7oK4EltiadxRvVR6K/yJPznpo4/XY
3GSQs2I5Yv3xkV6mPihnAfVkuXbwyR5BhPLfAjhxOHHtSX+7iYkChcIP8NBM
/qNUcsOqXMLQUOhdwCtEL2BEsNjHJ6Wzcn+a03Er9AnPzTi3DSL2+vUoCrpt
o6KoU1HWtk9Zh1+X/RzbZ0Zd6/fKBsL3wc4+1L2ih60XTcxvGM3NrxV/ENe0
RJDvtKfX8e+3k5Nzjhe8c+e5aB1ttH4jbIkA3xp38h+6sANvB5J87xcV4Wjp
SSRMddGxn9kmTzW2m/5c576UfC5WDduB/tTaylWN7QbVf+MuKPJWcsiEjKae
B10DcGdrkrErt4xtrmY/BS/5S8SsfHduXiUME3Mrua6JcWdt8A55KhedxqnI
o9PjyeodtHQvvcuEqwjdpUSRfxbyjTcXk3q3FWl/A0SM9EEbjsb+fcI3oAgP
AFhOPREhnM7GrxAj5jAfjRDXeF0M5ajkUTFG13UWI1+NH4mU6fnCpwVXwPmJ
fI77if8qd3iCOq/34QLC+WSe72pUZyM90qJe6QKZVmuXXI3j822vqbW/Jg0I
2vkxBUpGICEUCz1RU2E2JuTUVz5lpVAL0FV9k1mBaS7v1clNYohAaZZRCYSd
M5zxkEPNw7Hr5/7dYPIXlqGY9fw/qEtT4uXRp9nH7Uxk7mzpYVPhs7BgoMPk
w5+LX8ZKmABZ71Dk/bdOfP37o13RRFXFLbKfBWlCrSnoswByGEBTXcJY13bP
JshVT61JEjMWo0Yc4fXo37Ws5ejkO5d6X1MbcYlPplz0Qjbnm372rDbrMk/V
i2aK8JrINP2Y9b1z/dyCbutE+zCUy1E9jx0umc+0d4cnNpTmFgqwAcOn6vRF
Bq2oDtePHB94jzA9iijSk9nFMvmtaIBPIrb5FDxB5VWDjlEq2iJJf8ezwH+H
LPHaUB5oqn+vDZ+yB8PV8TLQlCLJFCpH61Nt0fnEk3a0F5i84seWUErtN2aQ
bhC5l5qH30OIVr5JC4/+N3TkoT+1XAOEqdhYpbM3eANN5pB1/XUI0KOZvpY9
DWcp5vd9Ow0imzAFpA7U+jDbMtC9mtEBfLXOqFWIzpeNpy4P3X2LZOHhaa52
XkhKamiM3ErF2oUMfS1f3ceF+OuwGqiX5f7TwVJnA8FwFenmLE2eU2+x52Ex
a9lcuLa+4Exdpd028yyui3YTrWAaq3oYiKSUDozk6D3O6ql1zrjr0da+G80q
tQ9NxCopG8etyq+RRcHfJXXFaGCKtv2AWo/BjfRzYh523VvIdHm2MokaDCl5
GOcQEpjoTrlLEqP+b2rC8CD/esZxtlgPM4urVuF7b2Wzf4diwttivijl5YJu
Dm+/kVgqOTldIDJ+Ap+0Hdb3qcMxWjoYE0+rGJwhyEZdbCarISQIb8hSs6Ql
taIxfMB8DxTJNXfUwZEq34ceaf4bTSX1nlLMjKpcUH7odm0zzVr8X0OuhlGz
gv8aprGVMG0C76EYrpys135mHO1k/zaNt96nuAcBfDYmdkwJCgP6Q6qG33wA
QHldqRNRI9k4MD1LNbxHYZv+LQkAPUcvidsAF6QxcJBhyp7VaOF3NQE+Tmfg
jXg7KHgz/9Xf/HBWXRzbmD7i8l2tYKsjI9kIARuAqJIdVJIeHiyyjdSqdMgD
0KgcMDbyo+kfadPBijTlPlhkuQC2r0cbV7WXBIJinzr+0X60W7JMhtgaP5hR
8wibsNb5Mx7w/kfGR0eRjwO5RqQwRUqaQz5OqWxEr0EyZiPdbkwH4SWlrNTW
UaVqkAtpJQaYMSgkXelUsymLe9FFoINViXuOACBsFXSepyMEwTX+fs2f38j6
aoCstsugHpCTa1//ujFr2XEUhD4IxkZB5KrEspjaIxfcPmSgMbULnREwAH97
KVOTGG5qzU+jULAAK/gMEeiH4OxnmynaWKaZL1xH304aNrUFGVrkRrSjPV4m
lbzqkLZ16U8DdciTaxyO63fBn3DSTHBqKdeUciv/OCg9a4zX4V7L6IBCb4LS
+gPyDQdR4FI9gHX19GZbAsV+GJT3+i5VG+1JM9FF/rUiyy0UEq6BUgpw8ENS
OiVrJU/GckXg1K2hQQkxcgOMLvRJHBcA5sNHMHL4XJxX4kyhE/YvMHGhTlzN
EKh0Nwqb1gqXx7HM3eKGUyXWVpK/L+cNp6E4pNnC1+l62zpU/1WCXTOENq4U
GPzIpUo3w+Gx+FI83uh9BMjYxQTLdhiGtO1TdCfkHYjsG5RGX1JsGk1KH29t
rprRCxIJ/pwW0CGFici4k6+ITGqJVmo5fQ5JvelvKbznzawW2kYUFDZc7WJt
8mtuB22jdoAO/Er0tHLZ4RgwJPEnifloh0MYYrredY4gRVTGxgO4QYoYDbxI
F2w/hDAeUaSpSGsgaWGVr97e0AxKawNbELcNH664Mdodoc8XLwRjrZgPi0Vk
ZUTNiIkb1X3f6+ai3OlzLKVEww3ln5ugL4z5DkcrEXzFX/1LGR4JpAEqMSCP
ESoOJabxV1quXHmHcmv11aLFKOOh82MsGy0ILcCjTK1VKph/Krzf3m1hvYE+
CY9FyRE2phdMw0j249mxstbUgepBK/4bOS03Z0L1M3ZODh/2yDem2G5pGlag
yo6HZo2ftMEIJQWZJTaPpMd6ZWdSVej55gO9AHsxJSEXtiZYIyAWG9xj8j0Z
4SZ1U/o3JVu9okI5llk5J+eU0th1A+xcN9wavu5k21fKqJM3lkCKYTpE/S7x
yS7Wv2hixFsLCjZPwYVVLAgo1Ty6+IYpmtEuv5QYNpl3f24b8rw01/a92ajt
lIcHE5HxCFhYJ8+Gg4JsqQ88LH19PoKSn6yOLPzQyDahh0XYbMJw3tyRQtlq
Gz6782/zVnA3MB6NHP6CU/pv+z7qIjPld/LO10kW5fygCdxrzAJwOfQ/FB2D
0ZvEE3boevKsJFCpmBPT5DnZmCWdZyOGfgVP/GlzlmaQMTNByz03whqHg3lj
dnrCwV+cbd+oqhr/8WDYjWhu7YWMJnFZydSLq8UF7zZ26Dp0HtZYlmqnyWZN
cLMDgWTnWWaxU1H9IELtdxDkoYmcpo9gMWms3OBHEEv4eVtx9L/18HJVZdaS
peqVPSk9LNbLvB4Bcc1nJ3ybwK1hjcC9LVR7RdvmsmJfGVmIvrVt6qOiLXhX
RKDiazlzMkOGryBXmzRJHNYGicHLSfeGQS7pJOB3W0EblKnr03rkIbZixyk1
n/duP3cLGCubzWXsyNrhGZhvF3WV8U9+Qlxogk77uC8dlRj+SB/xNOfXL8i6
qenlqAzQBZ7rydIAuYQVH8rX+rOuCIFW2jo7f2EDvNzYGSpA1urnALSXFQPA
MAVYhVdCrYHL0JOdm3WbP3HajmRFPxAzeeXLjGq4DkaAP2DM4Gw7FtitNNaw
9WRbRZTItKJtVJcNCym3jCdBYyWyjtI3d5TDAnU/Uk7GG9Gk9rzQoSnb895g
zC2n+IESyLY/r0s4BFE/I8GpdXgunl0trMeiN5tZPecU3TP56YE16ftjxmrx
V7caGB1YHDMqxrqEmg72L4s/7jN/zAOhCFAOhGPxmJhbuy6oqXC3yprzzlrB
vtYQVTfHycH7bBRFcasuRDCeIKRKtBOpPQakkYvKK4CmKPY0NzE702JajRfL
ciRiwOu0KFskzOrJWktddDxEC3XcUTQgSLsBpeXj6/O7pDlbKF2yzk1UOutx
JIY3rWAsHDKCyJYwFP7FyD+1xJ1shIZnmfIiCib/fjILMGd/yl0RX2ieTylp
jA0nx/1zwfkWubxp6kAovHnuPyR49DqzgKEKKHezj7iKc/7ml0cU64pLNfp6
WiG8mfgjs4YvdCnxd158t+s7at3fpCpvdzeqxfYLYXdZAwdbz4ec0HsN9+ZM
2vbbDj7BvXvNrPKhiMn2L/40LzMOuaL9LcMWXncymvdkeovBmhUv1KFdJXTN
8BrGAv1DNIhVmuGlzVaNu5jX428hU/GwG4GZLXLjlNvrgczvP2VckNr9G+jS
UVb0vHnIIxVmmRAJpUKqsfYDN3wl/Tux5Ra8wzsAjSY1IRLhT8sFzbHLPS7O
Apw7pKmerHefEkIF+UPNaPqtIadYHruBjtjoDyWu0Jt8WxfrAa2xQi+vwm/z
jyqw1MH6gbugx9BL9dq46mTak0BYyvjS1wSSFQJA0sYeuTBJOqzaa1DDwDpH
wF8v6jO+vi4aMk0YQbDAI4tTkQ2LSspsaq2ZNGNOeViPiIT6HwMnTWg3093D
0xy8mEU2/ciprLxYndcRelQ58ZFEmO7g82OiFE7xI6OwYiw3TXrKRvo/WTgZ
MI8OVIRqezgpqtyglpFI3Fa+t7INdLl8zB2ulTtZ5QCByK4HfXxF80+9obMO
1Jb6JWLRtEqgiCpV+ppQdZm7/bWdV125ZlX982sY6msO2Ly+PieOYXOj+b3L
JanLcoKTGApB9OPcID25Xb54Lrcy3uBADYiayfp/Ll+ODAmE9KQpGxpGZaKP
Nakb+eUztb1Xm8cfydX2G/6Zh5GcewgkfxVCWVP2enRCdLWSnPbDqptrLBWR
Ps7GuX+FRA1AOEIUPWcnR02vVt2///B6gFLlWstOtmeHeKt8/nZPulxlAXuq
xxFapbdC5nx5gvKHmV1QLE8TdVrzWpAHI7wK3ejbpzKhdPfLnBu15B2h2H1h
7lgOZqW7YDQpVPWVMUmMgF9MXeCQjsy4VXRScvgBZe8b/m8aZIk3gsjr9ooB
dAyhb4dVyxywu0vn7rbG4mU9vp7XHAMSzQEW1a7XWgphhavC/hXhpvF931wC
c9F4Di9ZSnCBJGxpuGqVGifKh8pMYHqgMNR2nLCTeP7iMs+uYuwMqPCbC6Q6
gwptrTNRwv0AWaSB97XHVmW/8fIlKfeQV9nHr47rMC4dY0wmXXyyujDOupJx
DEMGJjhA+0HdinzK5vrviJIiloKFkmHPMYnJVA5HumU+1uloon2KGaWi3441
U02E//oUPwAj50jLheeczgsa1F/NIZCJ8caGJtYZDwtZWNQfVwhWfsey9Lao
4mbo8iWxRGbjR2KH9APvaDYMSZRdT3dBJ9td+QEe6Ws8wrg5G7rxw8OtwGJZ
U0onk7PWRqlLkOPLFJCZVnTw3g5FVwfvuAg6Ih1YSkWxfFvYyWLU92zfp3mE
aOxQYuHuDfI36vLEqtnZgZVhVI92b5yQ2jp4jPX3UUOOTtK6uY5SKjqGPjSx
knIG4k4kLrkEkj3yEbejKlhKyxgyVYKgQgRFJdW4qKAhymfheOM9khIYNo9h
zAfQY2jVaWQMTT2sFCPj/6JE/LXZHU2YHbk2t8xioj/YHmdzsbc2tDmXq1cN
XMc6nU7q+Sg6gRuJSO9vef6NTN4c6yWJcJLxCmw6Zrm6cnPOiAfnQTgBRirW
16a7oZuKlKcpx+VxNKL1U5cAiRRLqzU4XtvgZqFBHzzr7a2v9DqUAnOB+Te9
y2h0HLx75rI8WbaQnWMKOv7ZmVQE+v6R5M3cwdLVHeXXcZkIIEQic0BzvWmT
Zffk328HX5P5OZH5UCsd0pSoxR0FZjUlx5FeFxuQdg+uYqfghwK1TKOQfZ1p
SYbC/tT2igHnghlNIdj0etZF//yQdBz9RNiQ60hRAmshp6kbLjc6i1F6MnVL
m5AWCw2wnvxNtT544iHFvjS7Dw+b46WLfilq0Q8WLuVaT4bg+yvxZuf2smLu
G2KMWUDKN0sQh6+bQSTe3xriawdgyTXdEAFnTgj/qF4jRb64gDLiwov7Z1G1
u0p3rnl3gdyDGSf4PC7KAV6ndEiRxZXzZZI1kLKcyID6FU/WJIF8ByK91bJ5
RTCvGoFwwyy9PkqicF7U1fnd5vYXVLQUQ7DlfOpQb4X1OAK0D7QmJJ82BEjI
kEpAgT8RHFVCLi8pAW2QUOxpfBvnWTBO+r1HV4SaQSJn8S/PdFAPSRhii4P/
yU7eGuDZxyNFqT08Opp/weq1XWtVuicOgGgrp+NUwmjTxDltgqV5DLqSjA6N
0b5tReC/gnApfzVnbtLed7l1juPu5vtpmWbiCxI93rYkYcEscJbP7VEdI8J7
c5DV4qhLb1bAorPjFhSEhFoJxDrt7wErcZmFa6Kjmyha9JIZ295r0ZUC/5Uh
MenrAis8CHk6J8lF/lfHaorazAuhZMXAPlgjJ4+IffrOefdskqCswp4ckKAV
Vreqfxq0vl8KZGUIcKNDIYP4kbSG6c/6txeUbHsYc+0ao1vF4qbekg0wp/+X
4VyBFsF2oD82Tc3NUy/cs7zZcDfYfKrM8CdjRfCjY/8RtAs0jLvK/y8ms4rx
zjXPRtsEJLNvHrqQmwzejWmPAoT9aePg0CyCB4yRKCTiZ+Tz0GsG3+8bCjut
lucdaES4E/kqAXtOloi8f1Q/LwRw7ZJtzCLPCott2jg0j/LoObaIae0zHxSq
gq/W6HUcDCATqFQkdfOIKTJPw1ysexykVNFFT/miIur3TI0BSqoKpFNNQ8tT
D2ZsOE84visRn/iyT3wNCEeP6AU3BWwfZbu1+IL+2xv/6Dyn7PCJyaNRuAz2
OIio6h0RJEPuEgDezDRRIpnbBOjjP7cCpTpgg+uhd10Ie8QLzW8RkHZ0MqOU
C4pR8ePGFq0IjfZqyZ4bVkOkAr7WkQgHSQW7Jrmxs4ifQF2mr/BAhAg6pV0Q
X9KEyUAH9BwqFf7VVV7McK+JDQYOJPv8ujuQj477ZFz1iiSvOs3olqDdDMdv
N08Je8lSYYFqV4KB49NbLbzDo00GbYN8PM3zj93EAKKcajc5f2ZvDp2g+XX/
+/WhKstTZ1HNtzJE4EUvaheXmWj/jSOOUimbfi+zgyxZVQ5jI2Y208jfBjyk
Jiz37aheNd1Bad/kJ7t+g40/ZFPBL8ziHJXTRPGsVLZAI3khSxDbBygI9Vw5
HBKI4Xf48sEASo/tZXgZ5eliWop7pREQ7uxuWe8L57yo5Y3dBxdMPIckKFkY
CTC1Gh41jnzXzSvYVt9z/0eP+2wkLqb7HvaHqmi3gqfIjRNxOjqfIi18pSOA
8tFLzpo4cxlB8jn4JUChEX5YFJfRsKAbrgtVqQpy04+FQbp8zF8N9IQQhSDf
gGooVpF0pRNkFudSn8+HQieeEafNeKEms/vL1AujOErFjUVaPYgbJOrCeXWx
UvFAK72/0WqqQPqXl6X+Gq5CRLFiulF70rqLXJEO2Pvh78SQj5XitcwkcT7+
KIvpiGS1ki+PBXdBeiV5wTA+TN7Zlhby5LGtiSjdFw2aZMFFJHG8exSRUM9h
CCsKURQf1oCYmq4j7i/qydlFvsidvmAbMRDVZC4jeZPsMvMoN0+JJ+H9Uxx1
nqGOzN3OMyr9UHlfaajnmOYmYuGW0B6YrhLhS2KSqoK4cxIU4y3zBbPZDVcb
0S5ydRlquj6R4XpFn3pNPWkonXssPxgDBB74JnLfwTjPckGf7VZbcVvzWhwy
jGylN6CmO+UdgM44xfQhwwKBMbRalTMYYmP0WfdlUwK5LtnoJtb4Ui70Vc5c
QtvVNI24a+bTD1f1pft1rtl35v1BfcTtwCQ5bErWvx8EUr0hy+S/q8ydzg/t
TVNMn+72GWFr01jmTA4PXQ9FmxaBo7aAkYqpJRy5b+DcaiiMxST4nYVMlUeU
nZGy8f2PqaPFhbfjb/Xo3GOQnHXv+Xb0fIfFdyXGwmtrZouDC5K9wYc1OLDm
bBfqA+TQeNjH4iozZkZkupRGwh2Lmp1Kpk2RoxnZXUvGO9cjOhJ+kaWW2fnH
6gv2glDU6lsZLFAxKEm4J3t9O5yA42ILJN9e3YckzOF63goBVlA+Y+3dbskU
TE/x6FHmeYoEmiif4ECaIHeqcVG0/cWgwB0p6DJdFoAE2G+h68xhmiLG78sU
VkUcQWu1xdZOZOS8ZEBdlhjeGzknYLtyliwLrrvTTkkJujgKRhF8pvpq0PQl
aP3Gq+979G2kZ3rCXY5dyRy4NdcPKCJDFu3RV8U2vLyra3LBmLNprCfU5Sk+
IVsqGahDswvB4b0u5ElxkFe0SxIGQ9u4ce9IoDSf/r0eSv476/pskLLo+uvm
+jHMtHpmGubdehC2fHJxB60VYx/m2FVq8Oku0t8Qnh5P7Yg0mCJad2VKqxgU
dSE6wrEOhA8hwFcqpmDMWow+FTxAVNDXGc/gE1RPBpM0gpqZltMgFcKHXn50
HCUtHLpigqX0LVLy9L9lRS+O0znTxJSNH9yBP4tLKLWRupTmB+qYYnO9zsHn
mthlQDTCYbY9fXpQ6W9A7gq799V1dOBEZVL4HUpgXZFVBgWWC3TWmmNSUdEA
9kcPYtsRCYD00ol5bSP+a1v86numFgMLdGjTPLWMjUyCFmvckBdCfaDWyyJi
KkZ/3sdTZrpnrhMbVxEEhOsL/tKA+73BaOs8FSTOvwcP9oBaKKSim6gX/lrV
lO9rVmhvSrXdvvxMJ0SZgtpanPhXiRSq4OqQBxCfpkCctsKZk5sa/4LaB4/g
IfX8uG/E2nDhjFOts807+y+WCRTqqq3e/d2a7tQs6VYEWXUFBChyHL63GuV4
AGddn9qIyv3o14ZejwJaEn9MrRYANnQGdvdgd5AcCqf+anwEWOj45Pi9VfWb
U0YAfX0SjSB+jGLiiCM9XU3Dm1H9v0yr2tahubmRL8Qi9oaO+MOcAZvdzmIS
AOcEegXno0mF7cG/blYg3SZaGoXhbdKS5Kpa7U4YTr4yt954itDitlCfAxrs
qW33rBx2HoEtD1ZIJN96Tw/wxrNPdaCt1QEdRzn8c4KYTY/FYgbkGscvV8iJ
d0mUa6pufXSVVox0FDd1r9U3NvR8Tj5shxagM9WiDCknJBHbWhqldpQxdbOn
g+7voAWCEtt+SOg2/Qo+u0p/cwkWS2t+bzxGyPyuO35NBhRFPPsXJFsgmFeh
VPGKSvm0PjJ+EGbaRCsnunNUpk5q3qj76xInZRqbW+rKYZ8dHC3N3rgidDzC
i/EGCR9DdHoHENTL2GYmnzgV3+ze0WAm8z7GMj42fgmyGS0Wlx2Ki5hRaYqG
HfjwpRjmSAr4yu+lbM/sKKn3SvyDaOWLp2UVQnZeNcDZbljA3QpEVdoY5HsW
8D1ftw8Hw09jA/UA6xm8a3xiHtzMtgF+AUwChSNOXRYKjnBS4k+POtghz7uz
sx2mAmEH0tKCexhUAnmSaXX3/N4WDiSDYD1oapdycONzKEYn36TAgOOgAq9v
jzUeFkCnBYjRrBQGoY8qAu/HjEt1wQx295n2EfXRkrcD88moFP34ywm+leWK
VducaAaiKrKIOCJL5aeTF6PtRPSqvnmt96mJLuSoAnoMtgAvrQZdAbp1P9NX
9zOdnp4DxEMRbTSCN18kL53oGDnndCB9VmE304726NTlN0z9qbhHBQZh74EM
I3RgeEfdbH37pZiKQ6A0d17/beE64CL6/H2+Ix8mJhpRNEZAFIUofpay+3pr
zfXo6wyN8IS99Gq7C0vYSM0nSDYcwDgnf3vNpgJcOLV62Tp5gLFCPRnW37zS
v671GsAs8dvZx12qt70FBl431s5hJKkLKpuWECwBSE4lkiCencA6cwoOH7Va
VBwWc1UEZ4TFGhvYJOfbiRpwg+wDRd5jPF5cZBTDYe8aQz59iNeu3SQW9B/Y
1pfwPNT4kd6LpEgmnt5QSPfjPmfq3btnubZl8dTyPpiFR+7UAOMQaFYGsAvt
y8Ey4EPz5pAOhcQlCE/dKEbkvoWqwd+86gIvTCCV71qO1xEn0UAYh4Y/4jYr
5VRLNN3m8DQozFBfmzTQs0whZsSVJE4msJKyzLyF2FtmBx9FtRencS+G3q11
Qvbx2IQlEYHJeC/pQFwtSCMKvAukp5D5iNuvFFaibRlisy49l2/XQEaH09XF
D/xpfG/kGXVhuHz4G/tw+57kmzx7zTL5VKy4hnaivDN3tXkJbijzICJ6CvBr
HBXXSSfzGLddpBa4tK1ud3om44mCN+YbjDS+NHC5ulAsuexRwWbhiErBIaON
aQQdEZJuD2sdRZIt7ZYD/nm1Z1Q3YP0lxJ40gr+t0Y4v2rqn9jyQesuuqB39
0vzfZ42bwLbhdg2EuHzPlf/kDWnlF5jyk/+S9mMJYoycMqbXoFMtQ5wKbKsg
wrPqSEmhtc2vUyd7XbfT/0z7bKu/TMdWQYcV/ERas3lkHweJD0oglgS7YWFn
NUGFSrl0BYA8RwEgtLM4XjtTLoM8lUA7aT9WbKswG+MtWKyT97IEU0jPq/oc
d9SHqSznyFKOGu/7Omymen9wgB6dmmXzhtIkH+bPbUcv4OKHDkkUrQEChKTS
RI8O/6g9Fs1dpQOOTMe2DV4QnL7c9xu4fOERjTl1R8qWbtMzbbTCR5URV24Q
hASCWH1P7BfeykRug5wlhF/rO9LZ9rVeyyY5AuvL30rMd4K/zfAT2BbQIlAa
wdSpHWhwfzpmjueyHzf7Ekjyjitnw9YCQLKzbET5vq9VDXQc/weVpnOFxsR+
gsQ1I1mkVufbbGwI5IriG8slhYUSjJPrZRzK3J28iVKFmBeCOJEfPwFXak58
GmOEFPTR0q3osolGAJzJU4lQSYuU2Eo4iHY0ZNHcEFIwzMYRc2qMlPcDlb+O
M4dmLlnpuCA7dGsC+AjuUorB/yiDafICMisPBAuru8lPxl04/1aZtsgGXIvK
CuHE4qYUuaY3XaAsUgksFrYNPiTahS38mAIJZalC7b9zLhW83F+cKGCmd6Qo
+tjFwVjJnM6t33jBsgPtx5QUFa2Tn8GZDvigCU+9oi4lplGAIC/5HPHuXupR
jid1a+edndjtN0XrTLO/r6Nvi1+H9ur1djyHGLD2O0o/HqJMI+j3P5CX2Gac
I39lY7fmtVqX3KEjcPk0MYTPs49f76JvgnRQuLhc/dot/17B+GsClIBYeoUn
uDrpXi9hbrLOt0G2V8WtZvvzIL02Pei4MfeeWDHpRoo+fZUfYYby/NcYNYzH
vUROsHvumz2/fRJiV2Sfkoj3jC204R0qfSHAWDbQ4tOOVNf8EZXDLU2Or2li
zLSzOcMyrvVlwoIEDN0L/EK4Hft3rQCLvM6NDIhXQQSivrqzCW3XCB3ZuZxs
mwpDPXwfevJ4CHLK4VIhEinAta4HBwc/RdjFSMPF1ue5GudICz/HTxbcuOv2
WZD0oc4uHzTyrwR83HuB4blytuTd3gFyvyoEtH7RN/br3SkApjFiA4mw8RXQ
Mi/4or5ZMdlw0p65Daj2Y1fM6xVAQrTY9dXBOWlP2qwRQTXF9AeaTZbLLkin
B9eI9klgVTBVOyXILJbY7tm30zPSd6IP57gVJgUjzp1zqjdCmfh0phgjOblR
NG5AM/u0utZNooGNp8dd5UmwaGbnPkx5BtLhd9Jdb36FqgZs+u1CcX9GyGgZ
4GluM52IN1iKah5ux10cmwEo0RrHHsJmUst+dttflSYnRmyThSPhbk8bfiTz
z8DJLWS2QjU16xAfnT7s/Ux3Cptuz8wB9EEYN30JocuG07+VrIDSkvju+RT5
apuXtA/29AOeYCbLi6OCcd821VSWHZ/0GigHDsnYfCnuf9c4/Tx4hOTzyJpI
QNjjCI/LvWSnx8QRuG+3tySaV1QOuNGrS8LMNppQk2rB9ngY6WXcEp/Oe1iZ
ED3xvmUgd9Knes1ntxrtpANaP1sWMyXUAGMOCiOJLOjH7jzx8UCCaTZOLsh7
kabRtqw5YmOkF56l5kyBo4swt4A9mZ4cCintncIvphGP+PE4h0pgubmliPzn
9A1B/BLi/7HyQkiXunQWJoXBQN0UfYTYg0FABHlVn43jI9WUOBnGa4FTEZfb
PubD1YGHvd4mnn406fbAO7RbEFcfEtrr6xbhoSwFR39ljNOnYvB6D3Xu6jyK
loeAtKCzvg7C3IClwwUlyqHg+HPUWz3gUFp7WyyZX9qsaV7dxzfQW/iOgh3n
xyZTGIhVrocKmqV9Dy+fsnWTc63iGK0O7st3/YSu5LxYJRwDUAXL74gJ/97P
7qVH3Da2wSUUyvt2+81elHIFfm8v9RiPFUFzyk9Wpk94Y5+fnkNci8XFtwoR
rPsiivCR4874r5ymojypNuSzOZ3YmnStEjssnb3zJLbPkdhMOVqV6wmKVJWF
vQcQriaOlHEO2CrrAC+Vt+hli1ZPMQ+uMiJe/vAA0bjrDTL1hmxU+ulsl3kP
g84SSWgRd+EZszeYqQXuzRsgHidC8lqd+9Vir2IHJsfi0+PFl3ZweojKndyu
ygNIRVVY5ECvV47qmYhwIoFPQXEMtgPaf+Ld4ntYfZNDGGphRIueL7cj8xxL
fH9dUNgwFkiLxpESgezVMzNWy2iAH9g8iTFWQobn+dVol9Ai8whpB0dATW5Z
ReZB+mtupxL97fpcYDwQoMfoP13n0s2zTnxMPZVFgjN/utC6CHXShY8s/N66
AxEGeki8Zk2kmOelj8QsNx/lRSwbL10/eQqK0TiFpUBNbEsl2TeboJePEDPm
MQGtUS9hsLfOhllVWTP4gI4bs68hG0O6NtJda0LL6khfl2RIq1D9mrNbvZcj
FiPBzlIiIesCaC+jOvFui6tWy59lozvKOPulmqse9bMFHB0/kFtUqvdWVm+k
A3k0qYlzPvyENLJ2877shHI+Gb8bMTZ4a7auAB3z3xe+BUIGCjtbRTpVZ3GT
BjWM/q/IzioXqX1LKAa5l7WBzHu4w2qPzlcvWn3l7C5sVqgx1NMn3JbxxU9x
PY5GK9myr3i1fqqdlFuHkMgnM3UqJMgdoStLL5lGatKEPLODtNW8hlWIIk4M
igAw8iYYsW5p9RI22mboTGZQ1HyR4f+mf+j+2dp+ZHhrz3mY4JG4FGjwk9HI
sD4CH1WqVVZjzGPI0S6SPUYtIQMuIdCpz0NGPzPp3TUniUx4t7E+t5ANa9G/
wHCp37xoAVnmpwF8SeQGu9kABIJEUSpOf6zYuwQtDASo4tY9CjF8C3m4KO5y
qQsp7fGvEuVLwd8uxZ1s4go5eFhHBstsbkZPsk3N/eZ4XxENiY53tHv8AczQ
bzSNXcVDc4jT8hkSWPJ2LYVnF0N+WO1dAUBpYygRSUHV9vtBppb0iWgrTjeS
BY00taMikd+62Nc8lu5Tde0kCLL5kFm4/0T1HLzYBziKuAJYhgWusaUMwMLH
Fm2ALNziLS850N/08HQ5cCst2yL4ju6Nvyi/+2D862Trt/khCrrk+r84nY+p
aHEuOGuIpWbHIlFpxaD8ocB8HoIS15ZTJjryHoszQ1KJnQ/yPvGv7/aTFTAx
PLroW+aVdNBEv1APH/ZHb5PW736Ak0NKvSKjal1cuzbuNp2to3p7lRwbEn6a
A7GvdHls2Bm3zguAX5bLOOdlheEopU3RXDFhdkVIaBRAjfrH8gXl4paVcyvR
emdC/TRapAz5e208EMyNnHrTWp8Kri3oKWY/utx4CXX+EudfsGjh3Ecsmyg1
PbWQWdjb2PTzaPFmI3H6a/P6cNa/L35gP7PfuPB346lEAMqP1MzXb4bR3gzM
9mWN0dSplF6UYt75i/r3ur7oGQIV5q1p70aa7YuJOfMqDWtMgBJTQOVkQo25
kHx+4deMgqv+67r5PvO3J9jQI9U5ZLdQcvrBdBLPDCBSIf4lCGQEyxk+kFk+
AtUWQA/zMej1zvxZhwCzVfXTHzuzV6y6PN9IqTC9w8X8MCa0Sfsmgav85Y8V
drv947uZa0/VWqb7bp3vp5KhlD1ibOYAJw6Cdzfh2FTqQleIm0vieRbRl4rz
HdtO7yfcSEUmvlnH2PYjF0au2XlNbIMRpptoNa4YtfRwVLBBeNXC4Qr5n1Bv
YGPG/Hisjf4mZKetmtqZfXDimQ8aMl6PacwUljn2Oww7dAiqphKJSAlCz+KM
jasnXPWZp7LkAYLRTxQfaDHRWgKaB6i7LjfTZkssYqvXvdhPTt8FJxcof+XZ
eqU2QYxVQarmgraaAJ4G+3L6BgMqdYuC73WfHjRrZF4biXV0uT/3BW8eKA3d
7ls8PGWKQrIslIvPYXg2pkeHdju1NNcr8TdS+XjcK/sNpVbE9eXy5i8QMRky
NuKAe9lB0TzqQKzRQPuZHwKQaXbJxAVM/MzfBRVySbXyg3U5fet0LxTtMYV4
N0OlQZ7+oPk691B0DuxlJkn6H4LAqfoD7fiZng0O3Yk756vdIxkJ6rXWivII
Bu3tj0p1Wp9/6A8MTnPZFW9VaifPUtR9WGGJUuwlP/G2H365a8v2Ds72R1K3
1QcIRo+lRRXbJViLDnn1JHFqrv59GPjb0ZR2N95D/m2Hc/jdF4koQ5kTAjV4
PvgcQxdWnGCAoXzb3HcNOASdUNUqJd0+/6WmyQKmmG3Jq0afC8rOjX77hdgP
8OyVxLRGDWY6WaKaqhEDWjWbk/59eA0wNbffbX4K6HMumbW8YPji4vTEQV54
9WylPrphRADT6eInKnKt13Bq/DLNhZQPWhotKzhwG6h8jC9Cq61bR8dE/BeY
DMlT2prgF2ZmgLocSgzxvgXRvsr5/yymzCgjNyu93vBdCVxTkqs2k7PAVVev
govJpFBLKDwpA+StZLXgtNjlHB9k2ASnqUr7h7btEEn9L6Fzu/3LiLWC4uMK
zKRM+44K06orKZKOg7FQYMrlKNkQj4DvXWx1EwikNaxgS+8Oi/B4UlHsdjYM
fWkHpemF6CCM6Qa8f7FMigx4kvTu4PB94DZh8WO64ZQq9wV+9W7fEi6SG3lU
yuixjoTBB6ZIcs/aEuf20gUcNQKlYT2idhKh+xk0t/9Xba71ZoQYiTC0sYx2
HcipiIteHupIbnV0q8/hqQAOSNxnrnRTuJMabgAdPupCv7xNvoBPi7DnNtki
3oC8v8l+lFojoXnRzImJ4PcE0ikxy1Cv9M8JVqkrTLiUe2AqbUg64dzjADM5
5FEhA+Wbs5+AsgZOV+Ue14OVtVyog8MxGocJDgDrcLOmm7Bt/nRqvvlc1Har
/oafDusHZGIVDLLvKkq+EoMgdE3JA1H2mI3o3EmArrOdvavTQIM37PevMpAn
iZ+fWjpid1/7qPDsCaEsO/73ruf1CNysyu0OukRHx47oOXQ2Nrp6lGwhQiIe
jrrmw60olHUzM7ucZsMhZXyJDd9MshqBJcB2ZK0OqbA4yV54yOdCCFxKBkZ3
3+bYOmuQ61H0Tqf7RX+FSf/McVkSLw88AuqfzCyLVRlcLxcdm+3DEOraIzuB
ghKklWLqzKeXX+TaL1/lagzzs4HQPhaaYB2PBlla8DuR4mYH/F7BymCvO50y
WirOGqd7+owWkh2gNspnq373OlTM2GHVlkRVXHQ3/ZyyjDeLwyUxFF1yUHA+
T2OehvwsPIJFCN0BVIsgNl9L3mI37ZWuJ7MszjigEOj2armY93dWSjPuvhN9
Gxe1ArOEfBccRIXUO229L2qrn+SBHFpBLYtlAs85zYDEG8WfJdhTH4WChz1M
vL05Qcb4KeI/bBEAh1JQ2aSSPGZucLMFJsUo2KN/PWwLr5ftkiVxQ/JgQtDO
MifN/6T9Z7sE6XYolikxbEb6g7MC7JKPrZ+2V+aFKkH9JeIH90PCuoSD7a8N
hkBGDD5CyHmf11TzpiYXUvMLKfNwOBFXKBlP6LgN37rPgzK+CAebxqQHryUa
fKA6rD30BbrGPCAF2hm0LzW3y5F7rWRPA3pK6lcQ2Oa/JfWkc615AsMGFXwb
Z8ViH3bhpkwQkigKIIYoynHsiBl/tLzDgbvoDLxxaVtbtS1L8PP21cQKNWgr
qdViJCf3jRtC2ImBQ5Ctp3ioP2tgcfdN0OFrIxRhoBEwN3rCHc7LLxyIZ/Zz
oUpIHN67V/osWT4tJezqosP4TR/CjI624m/kZr1mvJbJBtFmUPKUMs9wn3+Y
vABSwlgQQzWWp375juy2WF81RpPBWlZYKugc74bdg7blqUQv6H49ntnIeDtt
mGITmf+krW1i/VuJqEulVKBnDy2v3YCaO1xhbNVxf45we6Fm4DwfieLQxxog
oZhCfsJW6GeWwwk7Akye9qnCpuKHI77kfYhocSsrEo0Wt42SpFqa0xiDrmEG
ItBMVSKctOs66JrNoXvqZ+r1D0rawpj+oTvSRi3ck6jCkDHbOUu3oiUP/ql6
NGO7ad5OCShO/UYSzaz6T3W4SJsvBL0dB3qcpWnjPuI+V2bQIK842cssRmAu
4GwNCcoosA7V4nTH5aqf/hEmUezlz6/em6cMpkZBDevJKfeWcTxwwIPeu4HF
Di/sP9OxdKlZDfGVq+TMjDnen3K6Tnx/3QSlsxpvqylQhR+CXhwkPp0BzrdR
Uh1YSD67mCTNE1XZqCYzufk1zoor9zVzM1VSDm/0+AEy+xPOm+1h+R4xf8pF
IvHhGVL4PGeX6Pc0KPAvaudOQMZXukMWnBHWsxFG+wmnTjcjsDfjU76y7qyS
z4ejatf4f01Y3aqJrQhC5r8PhrGcHagqxzYN2u/G5btcQPxBGfJ2lYDdftog
wxBrwF1W3KiEcstP1XnisBjeEhSJ+ySN6PpYBclHO8yeE7nQRVX97p4rKXL/
Jtzrb/wnHnG37eEjMXgYwk1W6YkEcwQm2At4ktBzn1PBqtQGCSQWnf+FYPqK
ZE9DgPnwBioc/e5kORCGZjEH5OWmSWO8tXnXDILqtOsasCMKZAiRe4S0H4+x
wMkyKHaN+tT+SEkqCL5xLGQZ19x+4Vmp39orprAh/g2hnqDarcft0qdjgajG
gzo8LB1RqLCQq5hjCv9vnLBEqeRwENfu0yqvdDDMDYuAcY4aw7cOFPsj/RY2
YZRUjPkiU3PcAtvyIhHfB6uMnseolMu4vMg++i1e0ifQHHEpIdRVepYV+386
nbALIiwhhU0PlL/eRr922frkhYcA+OnW/hg5+El7p5kKjBqQZCfRSwXJBpmn
q6qd5HE/Shd6xmC813xDy5nJWeJ1BF8/h8ffoXv1iczQcU8E9gG5CpdUUzH1
4CbGkEbsi3mQ36+fFwoxItKMPmclHIzz2HC/dm3g1VRBJDEXsMbnPrQUTF/v
GJSzJ1V4ITAA6Ko5P/s6ISYLxtpJb1zCMfZlcg9+hB4UwhOpMSoTdega7QO3
uRvzwcp3+gPtJmCNh53hm9DyGTyvHh7YUcSC1y7wF10I29IkMunx9M+Ut5zt
QX6cNzx1KCVCd000w3FJ+8EzMXU7oOKw0aFu5d969wvMT5QmtY06MdmBpLom
yP8EE1Yr08/R/9jyWewU2Rn7HtJo+JL4JB5S7W40Y0ZzLnMQrsM/HY5naeo7
NVn7udgjYQAFPbzsNruciSme8/eS8+YKS+BYytOhYm1buF7pegLHcf2pb4og
qDnxOjKXOWd86ts6l1MKRzAFuDA4RDWhx0+phYjY3X7HzQfHkBvVw1vGf8R2
sxFPf9KupuPWJPjeYIVE1P046Xd2Wx1We4BgiTFewPGECAKbRjQx5PPgRKJD
pqHSpWbLqczzJnc0WFYgalji2A8LLIizJjOWvXgNtPdCkmOnOanCFsBn9un7
buieS7hdAzVDHFY3giRBg/Ttpt5o88mJ+ficBHbplvQsWMCxIGOUtN0Dzy0b
kRILEXmAMvo5amJhU6JXA8bgIvojWv9ShmFVX78vG0qlS8Lxd35U3PbBRMSk
nWOdDlOcC8P75ztBLoS8PTqPLgGinomiaurqlZ98jEOnfR0ZJZ7a9MAH4yZA
2MdjAO6IGssn6Dql+tvPTSI4YHrk/XQ04p0fiQ0OOLHrYkjD0XP01YataMxs
7JAaX7NEmMzqPmTZUHY9K2iJe4z4vQUfF0qZ42RU/theU2TfKJfHGXuwUq4b
KZLN7aBqHpx1GP0EN82UKTwJBeOnWdd3O/IHZOuItzCYJaEMLpCHWYycGjJH
zUCRlwXRzxBhfO2g5GvQkGPZRQEDG2yjYPS1rYQ80eposH+OgYE1w21Gb5vE
fw79kjA1LOZ4AOrpe/2BTkI5QMUmYkSrBMk/ABjHOFiof8k8PVYYnTp58Zyt
zM2y4138XqgfZKy8/U/DK27nPSsL5kNCpf4tDv4Scs/hiB46yUKQaLpbs6Mu
eEsNNTt7V8Y1NwjGAB5kRq5PSlV9DpFVieSmFX2YQ5GVM6Lfwm/D7ONu2pjz
oDBVWbuRhoO/b5IlYEwT57lbH8RQy1JineTOy/Ko7iQdCapAls5TxdhGJ3uF
ME3M1tG8+oK5753ngkGqJJbc6YKYsaBqIPRAbXfnhPBWKuEVTnAjHP1cTrtR
kN+22ynn9ynwV76TR8mbxDuVHaMsCVqxES5tKV2AzZXPy/zE6p5eHvp2pJ/B
ajyq1WDqd6YdPU2moIe5OnkLlMiFvECAxVNTQu4YlkdI5ptdVdZfQJls96X2
ecrz558YmP+pSeSmzLrwdD0EFHALdYgwDreBHVyQXiRdvFKBeGhv3tEuGDBN
ryVxMzrdgr9hQL5/ldzRPYhCx9gZq/PxmVsi/OhkfFbBDBrtjOrz0FxVACqT
eG2BMYRzcjwssZCMsupRj0wmo/Zcccl+hULgBIfX5X3z+rRun7YJvrw2+ML6
a6dvVTLscffB05srfqJ762iC+BPbtVrXfx0X1h8I37qu6OgCYJEw+G/DTkD2
+PjVHKk2x1ibdA4kItk10cBzk+cjNX1SlwVQdLLbHuopspPfyBAffojbRjSa
2He05+frpxDCp+CsmaEqs9Hg6zT698IqvM+9B55FQeLqIdQ1oy8lHgokFt55
uUVemwgRKuHtTD8yPlEmT352qkxj9vO4wpUr7TBjbMPLMJzuHNI2fPqbwq3g
VHl8nHEuJ+LDiOV6RftUqgZ881/wVhw2PBtdkzTBSb2UiWhcCKndfx6ml/60
IH8PCjVKwxHPnfAqVfgkvYNT7nFFGfuaITHRVULLMVOdv8N4axd/Tzlpa0QK
5Dpcy3IdKS+xkY7KVshKfi1b3AfSBWxvs//oTXxvmR9JhS7YE1AVmZDP/rxb
WdRb+EOwCKu+KPyiJF+AucAc7prLLwTNkTyGatT6yHnOUSzcTjG6z4SSVv54
DNwht/7P375sUUNsHXIeQ3MuhoybePA2CE/UWNacrLfpkh+cm9sAXPR5Uy6O
kkxP5nVFrmmV0xSZ3ns6lxaXVKJhUEfvGCpXmTq91YtIGaZJyMolAaDM7xjJ
1LQcrrOwg+p2UVnwxZf/7PZdEloe8ojzvIPa7cKfCdPJQrJN0TaJYKgUfN0Q
XAC8OXON48TEIKqqQAhCAyqONWW9KolhQnGDJSxpGn0+vYW6+FkRp3+UKkRH
5RYf8cFdtVmWOV3nMiZR7nDH/OXdF3TeZ0QCfHDHSiIJD2YVrWM15O31pgHt
YGOcAMzjvv9tw1OkmURRhi7CD3CqY9rUA5+P3hWvT9TPImkXYw04JgWA5o25
FO7VgXJ/FB21Kd5oSciADVjCnbS3nF4sb9gsx3BIQPh6JdldVBetdke1tQI1
xdpgiyMVX2a29I7qrzsZgw2cNJoq3HKUh4FhmiqmZ8HgKrZbz1IJ5ficnJPf
Cde8Cz83pAfGMf5JssBWU5A0EM8lmLK2pg+NKqbE4Hj6wEBWcF2IdbbDtvPs
nsKeIHO8W4ZNsmEvHmcHdqUwuevzffmYt7QBpWmQsuztSes41w0k9o6Ri1rN
eDpMp8UtS6Dy5sd8GIN0hLWDM7vMaeRhhx5kBcP21iXCSaXwtsKr1i4FOX8o
vQTpc3DUx/1QJlGmrlueey0d0UvbZykM4Wl+p1cmvDSafb74dxRlwROXFXBL
+zJCXWOqwZA6RtEhZwHAZ9eU9NqY+N3xJhkEdTcSQdrn1rcJqAsQcM0HJekN
3fKSk9cRjSQt3zp6W4s6g5gDHpFZvj8DI8tiy0BJ6DZWQ8gsPyul0ysphZdI
P0/ujBt041TcAsYoZqDaBUnmXfB5loxL0IKodFy1n9W0bwZCVwnoxvPP4+Fo
6LYCuQxhMEXtiXTjGaSudNwRCynIEF3M1fxHlPd5LDq+XouyVWPVsI121CdH
SO41tXtOjyNcJt5NcP7BPXCYXXmFWnENyrMGVRQWmakM/m27TB4H9MVjCWNJ
VJJP08cvysUIOKCJed6ea1fpy5riIsnbXgqtmIUhAOvez6rXqrE7+uRjyiHl
wiJ9g1GYFck6aQmGTlmqufoYU4fkmC2F1sg08kekg5ShvndJfaxCNxt9gMg7
zv9z0earrtIKOGDH8uWhzUQpx8Cwzv0PoETtIEsSIUFyV18W25tmSgIS0Bl8
iXmXgMKgF7oCrk7dm3gnWucaeXIwPdWOaxAowBPa8/XsJ9LDEnUyhiKZqI40
UCI+Y98ARFtMrhSB45aggdkxu71rOD+X7qKZrWFWFq9Ujgl97Kg+KSCD7e3M
wO1xv0NFmqNPK7UGnRkE91uAhVGvP2wKYsW0TPiF3ebDVHve+I4xFMKzGnwT
yzYMLLQ0lZMLc6KEVH6E9l+q4kxtNIhxjn28q30nQBgVGwinWq0GgOOSjPTZ
f65KwR5XQApcd1HO507OuvfcQCskrvtUHusFQBtetB1l+iAkuhCJf9Zfoos5
A8Jz4kKrW+He5VAm2tpyohL6xDgqAb7dVDxNwTLL24pkIhWH/aMC97XT6jUx
5O4yrhOeelE5mvnHOODH5XxSBaaCOHBJhQnYfJifh1WPLg0EfMaX+t1fju1b
rzvBRKTIpIcLzb47hXbpxUWUFTJvJKkbHUHwF2vS7iO/NCmq2AWZeQIRQCdf
e3+Tm/gtlaFfgX3rSYj4MI3zwDqqtEyykFP5f9KbnA1dMRLrXEyO8AjzcqwK
WGHoKw4bR7EGmFpmS1wzVbUkAAq7IhsWslzezPASJbLCDn1t5Wacu6FtshB2
nGsOi24S9rNrVdi81JOuXFbF8PJ9VgwRmpo7iWYwqYFtVTuCI/MEPVn+XQgZ
M//O3F54HbWxjBzprh03ZDkRd2rDs1HoVmj2PUa83KselqS81LNKkP7krzyP
ElPQkiQbGbDXKmRegP7fJ2fPNK3lZtoaK85ozLemC6l4oouyprjPxyAupC+M
bRwi6hWDsC56KvuOzyIn8lQaLx7qAwfSM1FzfzI6cHOeRjVinkUW//erXxxg
9yEIRjaMhy1LLKO138Epmw9hffDp/iHaR4J2sh9Sq3w+mdMxFUMLcbFeuru7
8sqsItPFumabD34uVUwS0+DTS4jvIEfwQ3Ub0yDUdeIv9g7+Mmjrp1k3lyzf
AwMZkj66ogpOi8uIAciE9dZkc94zZjRlRvGiJgGJ/AByVeGhdZp78kLIZaUI
WPfAC6pHgcwgLLCn8At++wdlbj12uo+aEorjsW07x+OFJWmTaPA9s0BZ4an7
ABTIo0BW2dswqp+m+06cBtrDmphIRePXZt1cHGnyNJx2CKVKkM1PSNxgrOYx
X/5x4rrTPeLdGBhpufXOCkvEWdU3YB+72sVJwwCDuKzRNgRWgRYbxeKRmuiC
af1sryMVizLfemUPdiYlKjxM4hb+DNYBFna+ix71ct9kPBe537AQRn1OTNcP
zUNQBoPg5K251w0X9fTLRq0ig1hykfC03AovIXe7Od1Toi0q1LYs4ivTYKK8
IYoiGWnWz1N0SshVXcsZD1RiMxB2s9L2087JgDiI5CvQJMV8AmEkAGUjWAP7
S4HikYQQupBcYPTBeR9prSW6gjx97o0dpwBbC4pJAs08hKhpIoU6kM0Fhy4m
gLK/6naFg27U89eQpMvJaiCdOKakqasu4LUTAUE7OOTS+o82LOMDI9oGTr3K
TVHKIAiXhhdxKBbFvvnGV6F/0nH8Vfcoq38XNmb1AM3AaVHZTg0SPMpMObW0
iI6u67oAYax27o4jxewhsdvEiseSg/Z7IJAVaCq3C7fwUhpbnvJc/EdUD/eh
pjeyhJ+86hHi0719DDOpeosdOOXzj3c61xwyJIIUIc7imjkoP8pLh1kLfUFl
kdqqUkvq+8wiGnWXDxEBzD73lxtQofmVkDWUrduiSKAWz03lp30FLl+100Ob
GpuEbYInLWCt82FzVZfjZil5BupwfGhXALnb3KUu+8RHCSQE3cHRcweCpIzM
8X7kUgMvfs/QmILGh21/6YRmSPePjfuNYyUANMDvFgBSZWZBQlH5xfSzHDDf
biWZp4jmUTBwz9OYd/af1lDGztBgjxIB5TT1gn98WFYd+G98SMJ7fv1LEx/U
Lz5G0eU0Ckrzs6FZnou9F1HTQGnJS+J50O6iX9tL9xQkosE2P+dXO8oM9jJi
pdLeOXl8beheaYWuHwSzJ3KNeC5d51AkyBWYfu4RfdwQWoTSupOXGb4smClI
kS22G0+Xn66fNlOoUIlycwaZTqCSmI16vORbtYvP61aIXwwRsZQ26mldGS9P
GyPoYBYJHmKmcdBHyMNYLKYZvoQ9AF9BWWan+YVinJEfqt+Jrt/Q4l2IcvHV
BDLTni/Qddv9vpo01+8pEts3yOXiOn6wn8i6sq9ykXs6hm/WTH0HxDZJtiU8
LKTTitnMcElBzH02f5mdIc9CxAwO/gJlERbj2xfTIlc1HY+JNINH6k6E7y9T
MD7VHSH2I9asn3MAjqmfnffbBgWw36Cs8+cmNXU6ZCgIcI8zdfyCcs1XnJME
KggLq5rOMLKdizGhw5J40fwLNCqkTIU3oSjllVlNo1iHIuowfAgETX7iphiR
53k5giCz2DV+kczc109OpasXKaM+He5sYfZAy8SASop3a50bFG1C4/WFPzJc
du/bq3ef04zqoFskvEYP6TRL4PlJTz8CODdD0YOgGaBvfregdNDGW/NC8IEh
b4JiNGU/c9nvMhxfFlRMpevNl+I/frQD0tzaM4XQfTEy/tCdBd7HuKoWwp6z
ou4wshs/cFgXS4E61siAJlj7VqPW6oRpW/iMaxpFxjTilr7A2fUqiKY3Uc6Z
HyT0+D8dou8faOk5T21RbTMelNRmvlGraIEYhi2OcTL6dk6zl2LMBpfZTuRU
bHSJJFNOOeqpuGEF6W3oMdLFGSPkl6OzZxH9pWU4sfIKlrEa59+x6C+C/zrr
E8dhF3wbpEeftnKC1ayJ/CqTjuMGFNhKJvMSPNmcAFg2Kap0vFleeUpSS8PA
xoGVNd8BQv0ZBfojIGve0l3GmczVgcw4g3ou3v1VTuSF7hc3TRfS2x06tTFD
i+GwoQdyxvHFBeLt7cIvHP13cRDwiCCZ1EJN57A4t+cfm/jxO+HE9zBM47+W
8avCfihHA29fq6LhUcQPugAgcVZt0wpEtXN2gagE7FuHrbNgIhbsWrGINaay
FxD2hqASyFX0/SJY8pNcSnLTBkk3Of6BVSE2rojRLEzP+D0ceOxN26rIN4m5
mTNLb7yjXeeRBWMN4mUe4mBJMEC+NW4zMYWHytnYrH3oSZWXXFKcv1uGm9eX
NcpVqQOROwkypX2+4j+YwMu2pUamRYWslA18wKuWQ8w5dLbQJ6xKAP2qW2C+
EtAQ9KS/DUE66CioP+dKLGRY22QsvCGZuLNf8qq/3R0vthKO60v9ADDeeOSf
RTzX62V7yuAjYFn4LoIJvVFZuz1bKn5YU7EynkYlVDZhAUfnrrAlTnvynUVl
pS7C6JqXtcl4Cf9vkVGMVsrpHVenVhMa8gBtrro4XmPToTV4bKtwAAHf5cuz
EFGVXCqkwrLQavuPfK/7W5R6NuVluhWEFN2sbFvPXOPx+pygF7UvmjD01tmg
JdsaEXGLRgEEdfIc/TfFSNgcPeSa4QvT26XEaxuvvMtnAhRZUz//SWeGX7j2
0uP+Td2GiYOQJvA4ja0PwTQRewDEAJTWQzCxrEPxPRUA9/7kDLt2+OP9U2HP
doi6Db+Mz64lg7rCrUQpQXWm8GVSvXA02AxYZqfCT28Z+dqGvuKi8vvbURtG
AYZvUPoxzMqlG6zhsu/OAn3VBk21DgD0BSSCYSFr6ugkjAOFjYDL/3joDLcn
K5bbqlg+3tk85uO737EcuhG1M9fFlufxwmT/+PiVO6TRP+9mKpI77ysSkt+V
OMSBzgX4DDRbf3y703Aj97zVwrRc5TlLC7+F1LbJ6k3M9s6lLp7rzvQnwyYr
V87tYt30UX1w+Hq+Hao5tnUR+01plb+XgD4Uy89vCC3LsfdJ0aNwyzuOxRK6
904oU2NGqWJ3M8tuksftTMJRYCNlrdyUEhoM8QpTY5MGydFizgAfYGb4aH3M
+SAPRVjxrG5/is+jJHaSi+bDn6uvMZMmzJPbBf1TzCIEHkAbVHiIXV6AfsOc
aIPP4MNcX8imlY1Vwscs7a/IPXz/QnL1HT2t5qX+1qNbu5jxftB7BR2pJ3M1
2k/SU/YzRAKWuvJCKMyLmHWG7P16vglkUeUgtYHWlctkhqof0mWgCETFuFep
rewn7Td/C2s/YFQ4PPlAi54CkedP9eGS0f7mYXMYYJ9Z4hvKKH5C2AKic0T8
/BxdrYx+0iNn3Gbim46+Ovubt0kNCpIe1x7767oKpbBUMfR1OHbIs383y4FC
J0OuL0Xrmdmp7yHE3MT5E1l560d8kW4r+t5GxJTCcHrSQK1rRCez1LEfNSte
MRfBQmoE/trxq4x+3BW6yD7pN2Cjx0CPzgYczcrfSNh9SQigpNUc/GyJ284l
d9zhegdMpFDleYlRKcHpkNB8FjTyBccwDbNP2ExQVTAbvrBdl20deuKGFHJ3
wFzdtldD9ta7i77pqEwvc4Js0CzBfakAfZ5IJ5HE77xNp3Pj0Zr1WZPHmU61
/YzlQUBRwq1HmLJo5qkUiRr8Y4D9AipYJwUprPvddstJVU0zI9frS4e8Xn+7
LerB+b2dT6dqGjExWW463ZM7PERliamK/qszn1YJ7fITVwdUnc5rUGK+YVk3
hjD05j7Z+UI8kgHw7sIhgSZL5PCyt3rW6Jk7yeCF24HPHNVGvdvnYqefqi/z
aneNEVj46Mn7NodoC+7hoMkFx/r+IZOJ+SzsCwCxUxwFLAlHtujdpqNhMIN5
U3rAOaqHWi2s1TAsZd4LN+jQcGt2fAxeC6Ga8pB3Qy7wBX6x/uQD21SpIuwz
QBjptAmaACBqnKR0E6M4CICIQ4Hjy7rufCYmk2bigbAlIMKTxOdtFuec2M0G
vP4JusJvYu8xtypnR8NT2r4k0Sw9MMlvsEj9YxNpLD4ggDZz6yNxkumFKOcL
naRIOpVv9rzTTeqXp1Sz6qh8Kiz8TNxS85hzGlXBVkejIaEYLxbpOYfVHEbr
ev+3FD1PJUJ7hqpcMi5uFeIcC1K/7a/6gRcXBxtm242iFXTP4yhdZf5bbIcD
6TAqvdBvSQBvGKCTYaFH45f5c/VcJ4LL7/G1G8Qom6TJ0k5pPSCwEfETj0xm
7t4yj/m0kPnxXuoqx7XIRkUERoMkyKZcGX5byCreVot/bdjiI+XnW6PJMu1+
axV38a9eNR+tevnHAat7hR4MO0MNdCVCjZT6yi647nrWZ8s2K6O8N2RqTuqw
cM0URSJKGTsHJXYt+FQU3sSa0bUzmnaSDwfkPfaOdvpAlG4vSZ1umIm3c1dS
faZ2KFU+SjkDCNrmPKzalQohk9uaqxF+tlozpWZz3asd43OXeo8geqDhfapp
Dr36HL9ciw5BVVcvYkhgYbnD4ZzLm5QLNoW6iBt2qfm5bVWcMOF/VXhiGA8E
ygQOH+/Z5lU2xhbBAQOYfzZFGZZsBJHfJ5DfidT1OrriG+KL9wAoNCXx4P7J
n4641CXNebJgU5L8XVdpxPIib7vlTsXZhneGAW6hsaVX6XAdLUC0ezc/Z/ry
S8mbWdGlLE8/hEeVU+fSZY79T4WctE+OXfz1tx4/3fqkJQiZ44lMgjUuvrRl
7DFF2Rrpa43QQgrRLCxeF1DidH04T6o622ConfUCGBDhv6ia5JPi4x5mVEGC
33cgHn1Iywjvq24o7oy+fdfKFeXcbLuOV+WiN5t+tgzbkiaa1FOBUK+7sTw5
vh0TGzWPRp2Y8wUWoGetlnwe+ehfBV6Gr57mwqibkN/xi7USH61y6g1J8F9r
34vcSOd2/w5wThpOpBqwkF719q9wuwJTXEV6+aqqaX9syPxeXY2h46sYyMPX
KTOlZrqMVsvLj7UPvrno0Qcy9bg16/xsiMyOxqvDy1wML7vI71pr8eitxLbn
0nd0OFZ9grDOjZ7XrhsWrlejpo5VPBVTBxY83PnzB3aROdKavS7vSXI4G0Lg
DTxwnIDTZ0qqrTPcYwtoPQ2P7e9NXHw1y7IBGxy2KGwzR+jOzedhbGn9nj/P
i94AZh459/bdJjp75aEwNTevL50xYltU5h/WSwAoMUzwYETwwsaLbZtZ7Fcs
rMgKoLJ/Ze52FdnOYee8VQNhk7o+9BPXbJ5+uclXrDkJM1wAIiahBHux3IYB
IviX4GplQ2JrvZx8F6q7H3ToO67TxqGyhNHNKJmUa2pA7po809rII9eb0aeS
skZxhTjQy5uAiU5rQgfmyOoedn4q7tvgjPUUD/UL8bB049zOhaScBGIvpR7g
oSb0BSw8eSBDzkpO1gm+2FvMUdU/inLl86vhXxrWCbRY81Nk1qggQSUwatMi
g8jkj5c/1nt4Lb/AK2hNiT3xs1lgpXMyJFefOJ3ITCcgQ7WMJBVO6YglQY3M
RAllLW2R7qUaEa8Yj5FpUpzteyizsb+8uJ22hQCYAADVjgGsOb0+YIzDRIhV
eG3xB4W53Jq9kUUpQYa6vTnrcveqbdUeHA8kcPi9kI1J9Z1ebADTvOhRlEOe
QRpH1lTKY0yn/B9Xrme8fqXl9wO2Po0pItKQwK6e78InFrzKyDBY+Yxozf46
xeHtRmfzIzjxpBxFSYw+DifAC5GQ7dQHVDiLYwxDY/df7MgCw6CXwz1baV80
g5xUWJiXPnPZg/OLUU2UpwNgmalVgv25Gdu1WxPjrIXB339woulnrmQ7We9R
LoNkrgT6m/iGWp5ib9RwfLnkVYAg+ZR7pS/UMMaAYKXKSZ6VUhKwDLV7rQ47
mrRPzXKn005SEezUJmyXGXdFZP7DMHD6sRXWjFPapu+eM+t+bMsuLradZHhi
loPYPuh6vI+aV0P4KDSwjGZ+NkMttB6TR/2CbUaTyt18Y+4EE3RdzFM87Hvi
RkeOGlFGIc2J69C3id3aLZ2+DxD+KmI7wQqfMcaofryFNpG9rIb43Ky5F/OW
4R+BfFyGSm6oP/cDo/76WVhY3Le2ImH0EtQy0BLQ9nCBxkN3J2wWr1h17P1g
JYqwPPz1kkL9JlS6sGlgDxguhf7FPBOuyJ+wpxa1rm5uKqUxVncs1gduplfl
83GaY2BFyq0YN0ihRkN0CdzjEqSrB6aEdaLhXqrAP6NJ/4OJsclVmJ4Ry5ky
+TUjoJWxcirjKgfHhWc2Z8KhqqsFMxM+TzLwzCCUiTZrqk+KUnV9NwMCEkSx
OmIv5CIeScDEXfJbga3QyfGI9/CLI39XKM4SY0kq53k99uOEy7Q5D2iMOs0S
hNCOGK9/PwdBAg+zEl55SLyt5XfHA9o42e1HQAhHDaX7ig6ubCZ3yA9ICG5c
VqOGciI9dyqyHZ7KA2OnT7tUb1/bKbX4saeZUYEK8TcpW7beXob/1s4j6GCb
rF6mP4Efo8Jztd6ZyZ16F3yv5NtopRsjW+eHCLQ9k6+aTMbUAHkBuUBxckeg
hVnANNSl7Q1gKRwqHuKKGCCKj+62fY4SoT+8A+nRsmUTZjDLlL2S6NTH7xhO
QjjhlFON098f7maD5X7mVZIT0ikSpKpZPYNfH3h3LNORLB+QkYKxiCkfT/+o
Th6FFxZoIsGgNPUcSC6zYdKj0ph4OsqR1aOy7ixuWrH1UqD3DKVFJDfjj51l
/4fynpDGL6zpXXa5Sgwl09pEvRHoqJYPCw0CjrH7EuCvyZ5d1qogmFdRtYUb
ICAK2q1a5LtuqbmrVBlUDR4m2g/xunR6hPAnxunRxFYyTTkkd3K3RmxbLLK7
GxR58kjrk7M7fKed7uBYNdwRwGkq1fA29w7tPgEO7YoUA1s2h7WUxm22W+aW
zi1pg0yGwvCe0O2zxipgpHbgJUxkTh29AaiRlQ5k6ZgPhR1abtIhcamlVvru
Eib/4DJa+ZcMcxKgLyFXPxliRj3cFKWyP6r460fejJjbHwtK2Cq/+ZgRFV1C
NL8VaWqTmKffBOpsQ0oIJbuWobYpFyd8GXZcnxhu4uGES62PKOjd8WT/n/+l
yYkoX409fK3q9Wdtq2Kd1JfcWFD2Cq2TxHQje0zgC7EGjSNXC+5T9iie29LR
CFMv5QTrl7KE5AtZsNlt8nVqAQn4b5u0LVp+yTNz5WmXKOJD0/ep9HiJtYwL
7zr1KAaCCf9B04d4/g6YSvhYNCqHcoVSZIghmOUO5iZ1OQ5jV3FiaScIPtDT
MDlA2baToF8+a4uen3nFn2rTaxREHuoxwxiVXbs0nY43jGAfbkItjHNIRH5X
C7xvqPHID/h/zGFaXq4ltAPXl25fpO/X4LyhhRVLep92mCHTq03TVTzzop8k
dqUBKXK1H2KQEDV4SgryCNvsqqE7YALNFU3LNPZVfv/sPC7xsQ8GF776TaE4
+JoQKl7aO+5KFB2vaABKwWb40zKUg0Csz/DOAFemAuLvNoq8BDy8kq/PsNoT
WRmod60iVVsgcxR5PfQjEVG+M9YX4uf9Dt7QF7UN1qSLXIHuwPPbv4tOWPc1
YIx1LXIWZgubiTP2m6us6z58+S86JDJpVuTLb6AK+EhgkEYmfpuDK3yaZIDv
Mps6Fy2ypdDhNYdsm78wPL77HeMzHDn3eGVbTMGkmfNllKVJ/abEQX4WLLKD
fz+PGakvjp1CsN47KA7VO8jHdF22Bef5mZvMEui8PRKulkR2zXf4O1Op7the
Hu3cOsryJV5mkwlNpwpy9SU7M+inmno7kaR/dItFJt0LvCdiZpvQHZSGzDNc
PGj1GPhlGlfVCdCONrz3htQksIiJiblpTpQemrJPOJ5KBNbbDgdqTGi1hwRU
b+7w0w7DCoeBuSHRNGcO2qtPTf+CyV79q903Y7eU0iHnh/g0VtPpDvZN+y3E
8UfgKRXXJDp1EiBRiW4cJx3WmBploVAX4dhRgG3BzeTv4SvIbMK/rG8Xw591
pdgQCA+vK1Fcp7WuZjyCjcY5nMmQt1ihMBVAnoykUI1edISjjrNFxLyv3Cwz
jAJG2DhE3J0UAn/vd0TcP6PDJXb1rapCO67MPeso7FkCEfS3q2u/vuFyuCkr
bf7PKa//zUtVZ2VQs7jZG4tWAaQPoqjLH2LB4nbawlup37inODJCX6TI+/IB
Iq6x6RoTZ9s+BkrYpyRLznme2XESxhJ7q2RjFTfOBgCT8z5Lw7Nz2rbAJTfE
+PUcLbVGRh5UqeCWROiDih6+qcfTDbwJTziQTupwH5SeRep7eAAPZn93LC90
ZC/YOd6zY+IeNkwRkaLcQ1/0W8/Gfl6PRgngdFPjEo3qCQL4iQfKQ9JVyzcy
KpJDBptjLkmY7gP86FmCk428Fp4jRlwQP2f8eQYyJRb+j61PWa/cqQVZqgJt
9Y11Xm9zhfoKWk7gVf+ESTu4VWIUwEgnBsmUqEIz51tZnnkWhzS/tQJKMzNw
NS1m7NvlHvd4G/8M/65fP9uVFcCdvEYGTueEjJU810bYYum16R2xPaLERvMA
2Dhk7qAL7YTfSTtthj8mVSkviUBJUx95eLe7/aGikzjRR1UAraFTktUCrH0X
GjGQip5oxaKJPh1iaKiLExjopyT3Kzmr7LSvi93K1MqQOIKmLwB8aCs1J+dS
9u8OvVsqCVRAxDqEjy+s4JDvN7yAsHCtCc6Y74z6AM5jWz4LP+Q6VDA3wbtT
WxOqivLbZ2ar/k9N4FU+6Kj3YyMAvh1SsxR//Cx84+ClSsxw0YYbqUI1zsJZ
rHwR5XP7GFKq/otO/L2u5nZKVijf4TpnE/XnmBhGK++dVb5QUGBqLVGNG6xd
20PZLWKoc8yRywykUSEHbsjL6ye8+tcv9ikEtg8rCiFwq9c9ucu6jcmN0T6J
ElJau8awJ6FKX1oEWQc0RDNJPmpkpLo/H6/rqrALKZmEOlU7rYjsuHfBYUF9
+7PnW6Kk99ROtXeFb2ei18SY0AFuUVh+vFpSQyicHSTeu9k+Nt7sVJC1yE3f
irW3khpUi9eEwzQqdKlk0uoFpfy0VWUm4c5tggVFYQL4ljabKtXDH73F78Gw
2Upe9pweRF4zet3dcR0SRHNw6NFPI+mklcmbzBOSyMNq66YF51NTAxjgyLqN
XiUkuLQPLmN2gaoAT7e6aj6w0xnTB7wbMcuECZcc7h5H9DbaVw3D/iPGlNnJ
YoPL9DWCC3nG28ZiKF7Gpir+Su/RdnBh6aRUByqpjpP7WKNStWFvrZdYUe+s
HhJ9aqYMwA6+6sQvz7OSUoyimm8V6sLA3pZlcSTs99+eNsLqsn39kW3Hyefr
ji9w0+aJqkLK7r/R5xEgjpid+G7PyX9uU98v3eX3tFYqbqcjaqzjSNh/iY9S
MSaY7uDpjpY025guLlcosupnQwq9/OpgdeCkxLM0iTcvpYejJdL6o8Sd0kkY
QIelIUpeJ1CaGTgqnFrtSidQTnBKpKrIYhKPKQDWvdBZ9cnehK22A+7h0w/e
uXZrboDrKqyp6cGrDmqIa1KTgl9CiJY0uYOFTFAzr4B+CN1gxKmkSpNKk2GA
YDcUeSzU9qv1hIOzOXKw+AJ0WGNAqP+B7NixTI6gjayx5weUIpni/4ZVOo0T
+YnXgkC8MDk8skggw1ILg12LkA7dlZzMn2IkRZcs/ymqOR9PPuU/Y9N0dvzG
fKuLfHkaGSSiGhiwh8etjDuDqvnrtXwyem5JnjNY1GRy/8ubx+0i8O2fQIuE
JLMXz7rNWaBipRoICQQS8oFZgGjobIPe4PHfjyzrFWcT+KYYaNhGlBL/GgAw
9Zh4Eqj2NCUEYlFEot5vzIM7h4LHk25zkaj9cTkOvxzhSuDq6JwZL+kMTW0l
PfFaYOx7bFZClmdFGglnsi0vhBxeXQb8w7/C/l1XPpS0JOzIpRKfpUs7+4k3
kYpDY6kixB/e3Se6iMFt3cGZIcm1u4uT/PEgKOJlGbDA114vAX9tYy704lhz
Mk5EJ78cKaUItbUgV4MrxRU8gx3FP2BpK2h8E+3P0IUmRhUMCuOyFzzPy+wf
HccD6ksH2BXCPhAKcnCC0p8d2pXoftzFvV5RWpaaphuo16WGI8B3Y4oRFPry
27zcjj2wNwBPT0fOHna6AUvIaTG1Of9/OGWSrWxIyEOk0/d2aRwwCIZBfa2W
/xB4PsUf/OjJ8ti8+bTKWiF3JVTrS8/Dz4Y9BECyJ0JM9Tmq5tDbssuM9xxr
ONwA79HhVXwI0hkNEj5d2NnaIhhNi8pzxDQYJwosKlNcGGo2QDR6T4RF/xQ+
pHTwMS9bAnA6oX+m1bJwvdBcmrPDqcvymRUo/egfkdGPiW/Cq/5U/ERpENTg
qYuWkl7GxXgcvYoEJg4nQR7IkIXdhZuFDMPm0fjBMPjRlm7ABxaS2081kHQg
UDah6tXqY1ki0odRd/uPV5bYFvT78gWoBlniDCGeEyB5e7QItQHA7kt36rnn
thlGyjkPg6WXRNH8RO+EPlbEZOyurV6L+4qSldomUPTAVWT8aGEFqiq9b9Bj
eguMX+jLDZZ77BgnF9Lys6O9jNA/7lA+iIksj2ZHtFTvOESXC0JI/zAkBegp
TSFYMwIPfL8JhntAEVVbqsYe9AIOwSxgkml/rkB08CEbNQqcjWzRc99XaU/m
CRbGQXpHFKg/8rkqvOKYuEZy9+QYTSiiIBWiqIBT0THOquLisAeB4u7Uq7uA
U0Eyo3a6gs9hh3LiZnCOqfzA3Dq0LG7aZZ09kyasMJ7yqG/g/yjMlrDJntob
fHbXQL28Dda6H93UJxpN6bT1a6/oFtzTTr0pS4vRtWjF5y9KaBfKh8q/j050
vBUIAbFtIsPtJ1dosMDkavGXQsTO6w+VqwL6wyQPqzAHaZUyUEqOWTq+VJje
IFr0vZErAqA5ppLrynXBrF/sGDeFlIPXpqusUuQ4PM9qOsg9F2iYSky7iTqW
ntrKUcHXtm57ZVUxrBmFL1FdgZBTzY2BJBgCZf/m7i4Eksi7A444GJGV9G/x
rw5ydo3187rdfpVXTL94AUU8Ye5aRo72wp1M023/dtw62FS4VtI8JbrFOKfs
8gDyoQEQC4KNPsyXyA+3pMWklQI6cWx/7S1OOEjiyfcAP6y0BKhAzydd0zG4
w9GyyiC8rCwM99RSccMveHBuKlGyXu/0iMTqStyEtDpA50M9Ym6AjncTFZk3
puHNmz0K5ZWqL/izBwX4TLd8/33anGGgh9vNZhej6ZI8BAd0i+hhd80kGVuY
DcLJIahg2FQ7yK+Yb2LkP/SYPfJ0MK6bzfeQ4R6lNyFj/h8YJbBuuvlrMQcd
xFK41vMeEmaN5C06sHkxaXUXoLox1UtnzbG9gmRZIm/bjFfbZ7qWFwbi8IqE
Vbc0rCOsUu/9EBb0I79ypMMtl+jM5GivxsdtiinUvobXYxJYllsLsQZPg96M
01WmqExrTYpXGZqN/lGePxG25L+YQu8zRXQJ1KS17fB5paE0gMdWV9Y81YX9
hAhSAty4zrrrvxji6VZhd6D45FtnWHoSnA7vZOIl4PPU9LJbK/YsXJ8Pec3Y
nb+gGqhNKUCr0iePPonhQ8mlC3bjnDHKR1mPeMt1kc+0HZjsx7VZBh6Iikqj
u+xAOaE9qOXIES52ESuRmX387EphXyqz5KjoKye4XHa+NcJ2Ln8HU39cxehN
qbD6ODzh8CwKSAt2iaEGvMFxgekM+0cDK/o3I4EExNkxS06kRau3xdzS6bIF
OOLoMEn/CCVgC+0EM5/uJ+szAAHS6uz9mqn8MDcR0KYW2c3v9W8mUsGzZBZZ
DCodpW5SJirLkJIrKkVkeyWC8+AViUHrwJfITuYbxUeDkWw1SxuqNF60d0fT
pZ96GnPiO14x9meNaZTzBWPP+5hRKqitw8lYCYxL/vavYoEdmxLv+9reC36V
oluNh6mG3Osy+LXtcgD+s7+6jQtOvkGESukKOmKMVMX0IsuxLVKqdqUGw8VX
tXE+SlHv4/F8WslFBA0KWJSJ1INEobxrDw5Dck+XEzgUFzXkucCNpN6fC4pH
0Geym3j1U0iOy4sstQYVdB5kJpy6qT8bjB5WFpj6IqhTQYlwzryFxFHT32qn
R75l/K3pT7e5XTdyyXgwUgJFBy7dtStO3YNXwZySQTlapemeNaXbz5V1ebip
CVEKOEFQ6t4+O6rtiw/CNnwpXi4k6pWl/yOyuLyxDHribOGBp4V1io5p289k
GSkrhA8Fsk1p/hANINi99QJ7FQ6r2aSIhi8N0F6sBgAp7QWakOehN/D7xNup
CfpzPVojoE4xgpOgam9CX8eLRF2qvuArmWGdERVKWiKSAW2aif2YhlYqW8wg
kNQLQxAlqEoQC11aRlXFKkMKvz/9Gc4tpFRedtNG0Pz4uik8OHNSlvsQH68e
hwbedlO99Yj9ju8l/E3AmvUfAVZDf5Q2rsi72XWLm+yfpMN/x1gTVIXIBefo
PZmeNSIlrWVUEKP6B6koypKP+0Omh+w2UJA0dUkuu4kK9+c/SH/p+EJCbRMz
U+sKgfD7+RZTqh/CfVQu5rmgzmz2GY6aoBDrJxsAD322oU0u/dAaJ64ameAe
Xlz2EQh3OEzVi9C9Ijh1/Cn4A1kjOjiFMAm8VPoAddwD14bLbpf10HiJ6are
f79bLUOW1+fmBJMhN308LqoNtDFLUcKK7jaR1WWcBTjX+IzbJmsPU9rKeZc3
xyxmhEqnIDMQ1wyndUS6Fqibt/R9Twn1JKu87uqJccCAWeg3qMEV2gDHftNS
9x4pd6rnyejN/J/Oq2wyoe54adxAuKEfo9q0DAwg48Jjx9PRDPDMivwqzNPt
cDWDcZ3vrPxWVKCa5gux2KSulAwExglz4w6uquIa+yFB1M6EwSKisHZdO9EA
0eojlqF1czQLKfi1FLmG1sDxaCtZ8tyDabnguXST0FMdwOlsvZwgzHh6cny+
aFiNfqr4MzPnK3jNuYs5FBOJ0TeqTN+c2hV80zNX1Cp0fQcc9o3lAT1d0NG4
tzE5GMcVBjd5OVFtum2ZYlY0kH6qn5oFGCCILupKA1MxHiODg3XxRjKPEWU6
ish1twx5rwtT17XotdG4pFaUgLIfDc0C5ZGd0BUBSdUjLBp0JxGcXM35XkmB
NamQRfdAfQaWdWnyD/WXL4ghmQDlL2qPwa9ahtIxCCJFPWvWxu9mW2wlKlaU
RYiPQMV6D6SvzE+nA4WKhtaRfHeS9n4EjDy/rAPEUqkOG4d94pSdFKzJXVip
uFUxjZ0TaQMU6j3t92NHapjE83j3MwUOu2lbfIgdT0wHqZTsJTr+eNjKeVpU
03X3j3A88qFnFch81E/GI7H3FsFix1NW5lmUKaR6h19D/8T/d0+HQISieDI1
eYIYvufEI7OmhFaT7iYiWxuKHC1ZNWDYzZdsg/MxUv5cJlw+7pid6SsLVhtK
m+aopAxvccskQyRamsYbVlz0i5Vj06s2A1LlFGy5X09OoxE5PoKvsQNXU8mO
LJM/NcmubGMqvkNuMKU85iUsiWsjjAWqoglNGHH9BuMzlUAmL+I/83dOJQ23
aCQ3NzcnhbgSM5PfVbfP4KTTmzWeDPJdiUxwwvut8hQ3n/7oAbdrttwpQAKi
dIZReqJ42dBBRZOaSj/ZJxBM8rGlr6NNjWA5bTkRe7+mcGrr8S1IrVsJ87Yj
6QNWq0cteL14e30f0c8ILI0d0TN7JZxRKRqyVsAN+NYyGMPOExUm2OLBiQul
bMVk7VYHJe5zjK3YKCfA9aCbB8zbZIhm+Qno4KSxU6OmdlWpTzV+ohb4zTGq
nDDWgXZYPn66UqCcW6LE3UQ/ScW7AUYpBFEE3tsNcV5niJaeJvyMJldiRApE
aBfb/tt4FU2I6WlkpExM6Mgb2z+iDQ0FhHgwc61vv3pGFfT6u4vjs6A2eOST
My4YkORxawI/1kk6kncandNQ/REgWphN6qKgyFlQo6vvWMwQ3uqP7SEj5APP
iqVLegE3xOIRTOOK7oF7lDFHQXDggvOr6n5wBOOPyqqhQbGkZ32QKBIqApD7
VjxmypDGAXA+7oyYL27TCXrIK85SKFo8o4P++SAoeU6+n8IDLPKEaV1SAQsx
Hu8zGcqhJd1MqxlyczPS9TV8pDyPp+IQKFZW89iGx/EfwQIUU0OI/ZBUQgNY
A5lJq5lk3KygAoHj39nsWe9jFTSui6YzicwBQXd29MzqgQc4crTHeh3nWBl1
TOlI+JwIjq9Lm8+3m2cI1GxZI/MUPgzHy/k8Bm3tBTuLIAl7actKBRRNBcjw
CKN5JqnirDYOvcFeqV4sqmbe1zxWSiSK3b8UrA/ZraSNC0EZCf7l3HqI+Tje
tAQsuShFcLg66/r/ValJO2KuSXeNjkVfxSBqfRcylu+gj/l0nfcglO86ZGQ5
nVwZNFMlFCTTS4UvFweyRwVIJRE/My/aYgHq03VlzylMdipMFrLbfWftN5Im
gIgS0AgVmuK05M8c86HdXL5qlco2I9E2Pv0iP8imNPCm7qVsyqYAOkxhgM1/
Z49mWo1zcXwnojR6lg69N1FKzJThY5H48f/GREPm1imhz2LrW9Jg5DN3dzNL
H1Ci+QqPMeODK36ij2dRveUh5eHd05CCl8Tfz8dEs/wFyWjuLU71bS3MiHi5
gj6OXiooRblLigatri3MNEbCGs/1PQ8oeDoX6DK/jNTqWBPnlJHPFNSHwcoo
5l/1wtcRg+6jIdoMKaNGx3t63t+ywM1ZXHG5FEGyYYIGlbT151N1/ALypim2
rz4oQFVEz1ZWhsJvzyD0QzV+AXyq1NbwU9se7toh6WdsIwed20MUmEN6+Gey
1saNm1Px3s6sWa7izN6HdGD8Oya9PfQ80T/U7ClVgvEOW9ytkLvHmLaNFLqj
GF/eRELSQ4MWrtlwoHdtrxRzOo6il2/OIr+Qlg8ZQETefkAtMbS5lKYxi7rX
HriQMDemLXPgQBp4jghEluDzJiwGwAXAuvPaigfQJXa/AG7S/VnTJjW051nG
0iW1iXvYO/mR/b+Uc8oOAcuEX2awN0AjlBEYLtWoKY4NRUovPA8BXrABqPVw
PIAUVfW6i9Mt4MfYglEBrzN2au2VP9zKQvFmb3+TDEglDbsmQd1hWDeFj4ZN
SFUu6zpykT3CClfiVZgVqPwKgyYVkr5+EHrj7QvlGv77Sn8ElJp8zzdD2SE5
PvEDbH0b8pdXhyFKiI3MTiu6jiwbPQoUaN7dWxzKJsT+A+rPkYH+rQpnp4MN
Jxt0PPe7hwq7nWOfmVc1u0UMCP5gBozSGrLkvCb7TTB+Cys/BTOPeOl8mXY3
/9a1Lp/46qEmxCLuDl+JK0YhWMnGPGFOEQq5DDpHykUvjsM4lQKneqUVUJG/
CGSqB86W9fGLeeqyxjyUC6vn3hiUvjviesNE2WgOFjN+IKEuHxkW/FJKYD5N
GTUB57iqMx00uDa4WdLD8i8fl/m8TE+hYml59ZdeBwH5Q/HmqOAm8EC1/zMN
WKXA/b2G6KgGGw4lVp+QYU1nMB/6qsgRavKtl/jCCSyTET36ORcPmij/91CY
lzVBWh9efY4nnxsLteVdOMioAbytaRdq2t43OAVyvbNFEJC+EvZ3vel62v+Q
N69akQVIRW0liALtF87Hmq9Vd3CPlyXxlCdJ61qq+nyfza6Gu6xUN7HYdoOw
SaN0vMfOEB5L+tApMZ+1vR9vHWNc71k06DNwRcv2Bud4La8rg4xaGmEHuonF
aTPKMFlS4/dKyaZ6GFvyMuVsggXadY/zEhpnemiLLr/qwsiVNDHEdm0vgdfU
IiA4qeklKUAXSm1RhfNjEFLITV0EdyCQb61oyKISTfT19O3m6xjfBUjCXEsi
en/SOnbBtYfh6LQed3xXPPmI9ktM6huBytDXaGFtgFtJyNUOREhl/NTKORQj
qi254AHxWV+43TWvaKkQy4Kjk4TWGBqZsqWQ/k8AiBMWnSpIEi5OJwdZg7Ei
NzADaUszu6E4b4YqyPYUMuobbIXoxKDDMAgbNapA5GlRzSD7as+IDLfnhOOc
S7WJF9UXomhCMMEasBRw1xVtxPoAbkrJwkErrLeJvsWDFivv9d3x0q0oFqID
nbiJjdf1HUrwgHPMNxh4Qd1ouVvsTZGvWN7MfzecYf5Ln/6FWiN0VeAwChBH
ielzELev63U2HRAVX0Er9ifkFngqbiXkGpsp0/Uw+TgDVjLZIe5oH6n4sf8v
buCQeHSRe6FQrlrAj1m6V+hyi78rRksIZXSjyN92Gy4DLbZ83+WIRJCBdLjo
/r8W/jfCDtj9q+w92MB+PRzxODOYtiXPmd44X25yhJmd19zFrAi7PZAYUGoF
iMS34YGwG+fs2QeiNJ6MVHyXwFdKgW78h43sODN9vTL88Sw/mp9YvQp46NHG
t1fdg9I7usjIiZZpeqVNeV+/FflrJ2AB5qtS8b/9nLH9EDNdwZNKiP91FGGM
EOG3FZ8+8uWCvOUy/NpzH2NE7j0jL88d/5Mv1EIzwcEAdEEQJ9dL4bouhypX
JNLYkuTfuUcaRYhOfRMuaixVwjiKObuPxJm6eDXM3nuk0lDIKhzh1JASgxhZ
Lb1ARfPVGA594y8xcBl7MwKOt2wi/1tOPr4dxLtvV02vxQZkw2/OX3LpUUiX
0Q/1CquT0PByAKI80y3IHFwntLupE8JYnIUC5cKNzlbBftrI+WkFf6v+5Map
WDul4T0GWyIw0Flu9z9LWMvyxXNcXFPAukq9FU/re+YFfaJHmsQXBkEwjTo1
yD+uz39QqBNXdPliSf9lJaFC0qKzjNRUcw3zsXuJZvEY1cVccXtvsFi9z5NU
jwdOllthZdxikjs3eC4s4MwYVsSyb5Geiu7J3x67MRYiN7r/w1GtEhAtbH/4
jhjS0gR6gsXOpvGEvOqvMDC8jhSudfA4huerf/BQXScWRdcTGe1zzFhYRhDb
FJovdNDfmYU5/e/24mdBZxX0p0cy/Sc4VzjIj/6BdlUKDoHKO6EJum/tQ8C9
Dg3YZMORlP6j2QXjL8SjjNf+hhpzb11Gu5Ldl4gpN/BFSCj3C/H/GwlgsqfZ
TLbEOqZD4G0dEV83XwVfF8Fh8KT2KSU12JqacZaVjJY5INX2KhN4b6pJlPKD
p+tpXwfBLLrKk/wskqXrbQeZ6VvXwfsOlmqphraKwL0stbo3BsVhAOziH2Xw
YLNUPiqjtAYF+IWDTOWoiyDwcMYyaJ/agvWtyqnlUJkC8fkOmbKmJ8Agl/WI
ljIoGsrnSy+Km0NVV+qiF2t2qSCz77blbkWU3aaCHy74utyGJlm1f7PSxbmZ
LIq8dy+SRtgBo21kgvliUGPfUY0aSTS/txnbvcrTLJlytsU3egfE2hW4K5i5
EIpoGPqH5VHymbKTtzOGOexeXQ1yqNL4rmNIgFzo7ZuhdxQIt/B9GHIFA8/Y
2R99ICaiVeghqy+jdLjfaGKhVmu4xzZwhld1D0nYBoqx9/9qxPoQ/qQvmvq/
oF1+P2oxvVwVb3yyYxxdEJSDDg4GnQcChqurkuLTS5OjnZs3HtfbPhngM6mN
9UuIZj3Ve26LDXWVE62gilMpMGGAmQeiMyYXWuuaE5GBl2HoPc6wUHgdewXt
qfgM4UNjt9GEthB6EMnt/Ktq1QVStO65mx/dVI7UsyOX4DU3X6nmUxQUC+cO
4Bdw1Zmq6+LMLXG+5UlHYYwuFydYbDjYJHw2UfbgGFOtYbUR7PfYSHxOWYD2
BjozjnQY6qJVjQ8c/G4rucC1kx9gJ5qdKUD+8oNl7HpAdkVrrka/zQnHOsOW
Aixsi5P1OS/lXZyBrwRBUIv8H01LJztY+lXzPWgHall+sCrbnzmbaFtjpAV1
TCoKtb+zsdjlDadXBXk68I68id1LlQzNz7qYgvOI868UCVEeYjFTt33yCJOv
kI8/iYg3uVkUhmgwgngNuZDq7HLMJXmcqvbmQSK3kpcTCSYq1pEXmVOjuG7W
wZuTTuTX/SLAw+/ZS62DXlMn5X0UwekaQdVwTz0y8JfLxDRSD6gIGuv2bht4
765vWvgC2hqNiaG7NSfJM5j+ApzSH0Ly4Ki2wfv6cLezmnVOVGpatTypTMxc
xKO9wSor0UmSeThdjN1s/+6J9z7Cf7amSLrbVO/htE1QUYyx0maEF1doaLUE
uryIcF2ga8FBrFV3RvOmS+z2JPUaABhUYDWdw7YSLFjTJtbch929phJTv9Lm
xhFNdfdFeIcJujh1qNKO68CQpcjGvN1fBto7QKAAGQnRdlK3phD24BjkUStF
28o637Pg/rkt93I6c/WOOTfGvTL4Ux7lYxEqycxz9hE+H6gnknG63vDyyo8E
MZo/w+kwG3I/8H3YlLNL5IngKn9RDnVFlfE4v4mCeKTKPVnfZNwsubEowcSJ
oOlAo9VLKeGNA2uoazW5am2yHDqEU9xDViN6Ts88Io/ZZbrAyvuIk/MzYjiI
FISbpR//4d2lGS7iGxy4tGTBnX90Im8OpvaRCrigfphKoSI0xTcQSVp0pDop
PirN0+8Pg93LigJ82hPD/Sa2Gofn2BNAF4PSyuhmPteMie7RVSXBhB8z2dkf
QcDYEESQwfl5C6bHu2xOW5xiqBMMiGGwcgZgSi1Yv/E/FtHJRGOaPFENx0CB
AKviEVUtZUpt3zI7ba3NswC/j7Oatt81zqs6w/5kqJNQD5eo8fwOlHTHmkdS
B/21GxGw+WxsEKF/yRcfNsKcjQjJV2UBBaqjT8fGsm4QJGImTY4Kw1Jx6Rqg
rGeweXs/sOWxCN00WY1uWalDdBZvMEAHnBfw1DVAdJ/2FuFj6rGXI7IAR6HY
iUPAkeYj1ihpTTXbwDYT+shtM5/63Wt/Kpa4N4JIcG4PzRnLN34kIJNGnFYC
LfZUVtnFGDJkavM6+uW7JYcR3bgXDaIhFuMMvqXdY4YeeP1ztO3I0AKTs8sx
SWnLkHqQwQKzmaWp7irBaylCwHozUzTKnZSOUJNvjLCQNFUXR3sJNizIDbzC
6LuksXpIdVGEp/ZkKRdBVid012cZeCIcEuY6GElHGYLMqITmNBz2HyFmJeJy
1XFngXmJJ6M4sB534igxAoIvCNDatEC9vyvWzVlVPxWtNrNV4rs72OQqCdyY
D71GFN6EwsKpImyjuUQ4PUBF5+ajMT6YDRB7kXaTeRonieZxprAKd3kyWakR
zOkP22dVcP8ZfRZvSYjOE5I+Ark6JzMUFYFZFqwrrSHsTVQoamcO22on9e7k
OX1WcvDaCa7/dRBAWc6ZYVoH/CJ+kwQk5ejseEIqogwh/Aj/ZKSUwnumD6RV
2E7Akr0HPIRpa+V1cDjFVt2j2x1uEru3XX0d+SQmr12E2mfTRuNbMqvyizYC
XCiiWsTZbMSm2LRmOvLcaigMsSV40UntG6LGvDWZub512ZqZAm5R6wzv5Iyz
rbNvNSju1TIjqu1+kcx/PS8XvPHTbstNtSoETEu1XpJXaes5fwRon5crF5Ry
kZGJs9iplVGk5KqA8h7blTh6zCnWuPYX5SskTMKZk30v8auCI9me5EeLT9fp
0417svQQg/CL0CkRS3qzarXlxq4YupWvb0b/JqtefOePX54UP+YP2fW0LbsK
Gz7R34bk0Jk8lknPGdlysYoW9pcN4ZcfJVIGuTGSO3wXWzs31wDosHCPtRn1
+OXv//VSGxUDKSiDjiK5ngu/9p6EsStGNDdOdCj6y6We3un2KeGYmmGE5E79
1lYsr/mDBYXl2TFDJXRTdUU3nzrr4QGMti3LlHaxR3+I/Q0bwoDvaFITqMIa
5GN371xc4SSvQvCBPBhBmFk+2QEKbtuhsnGKqciunvgwFdKwrrUrhdjvcHkU
CgPQ3N9aH3APMijD8jsFryax4bKG8HO9oD61avlhUkoPujMtRxtvrM3UxIw/
mWrM4BieBBuzzLd2JoHjQDlMcbKDSs4eZrnoiPGblrNxrl/d3UmaxvKpvvM1
ruahZ6V9Ye6Xtrk6Ii1IenF5IuaTV3iQ+fgZxOLaRr+pCV+Hde4/boMpC38+
Bib0MKz6jkCN7UXnH70c/KJmMCDf0jO1QsQm4jOfzdDnhOQ1M0wBPBvG9Yo6
naGroUrt+OxmQ+Y/Km4ZmlwryBUNR1y0FU6jUM0iDvKM9VcTovE4I7bMVmZK
sdEoHCzik1cBfzTcAx7C1OqSn0f3JAeIUnWb3IXZ6KqTYeq68jNmgiB3Ja72
xSTYDZnXUCN66ZkZ5EDJViZXX7PWgZ4rsp9NGYwE7Hi9pATIICYvmk5m68Os
KNfMuy6sEiaGuttCjqjgk4Fs5isIdmaeDohQx+FgNDQwy0MwMVRdRNKoQB77
locTfWsSi3wke/sUJMIsEayaWxFY6uXd1c4IANFgKcKjbz23Gall2OLPSgPU
Cy043wW5ApgsZMbD84SKawwtEK1I7+vWjeSG/JPR8ZoolgIGijpETQQynR43
Ub4Wyz1S/HLD267VThllvC/SBkdjZ9uRp0HzJ7tY4HwUyPUPU15w94OmKI6W
7UFJLoIEc/P7/bOERfqWBtubXqmYTsrueYLIHHM5YMDXMAKkq1jz7M2l9Fzd
YfzMd3Gr8Bpt2dxLyBTMSlRsvTkzrF2RjXa0Ch6TH2FwfT3tmcOxTtY6RX+5
7TEjSJ4WV2zZbzVEIzV7+uDDtY1d/RfHAnRa3TvIY5YqXOQf2hAImSK+hWeM
Oocf8PBVCgay5tp9rP5mE5YsBqP+ueHwh6IVTtxc13pKXG1bM0HomCYEoY3P
qi6yKMijh6AVLIZjBx6jf3aSx+BHWw/FBRwBnsvE+pvRzh23gVC+IlAHMcFL
dF/pk1eiwqTBn1rtzoflhZSRwprNNS0EedkKD0hG1PM8d1Kgv2wplrnIMTHN
k7+mzrpDYelGNvbQSmiWP9z/N6f2vquiTYb5CVgrxHKZx92UF/hhniL6jRC1
8r5QLRNIIZVnhyZWqehEk/AQEfUKjPWR5tlhSENhMHNuZ4WnwpvDSvUdycVQ
JDGlhQc3gqf/oiORYBQ4SSQjWsHJNkd+8HMVbuEtj5VlPRM2wUP4Topwq9rD
Qs66W87WVk77ZY/2FHtJWv885mIQwVY2BqK//Vq96vFcN8Lc6U+L/feV+1+M
jGHqoOOEg8F5n2zRMB1bpDKpSLO/kUpAnSc7hduio7XmH5/r78YYYmBXDB1e
YeJwWKc36cHCwSPgk6+ZlLbVjYs3vJPQxKbOTa+yc2ZjtNOouaKdPKYakOlF
47mqHg/kcA5uaADEktckGxNoXkmi6evNEM9HZFcCK1aaHVnY0Okb67ZdAnzz
7jZMXY9UPTrQyNIcy+K8uhAmykqNOtLT9ZqkmgteWLqltOeNU/KX0a9aYpx6
GILdVRqQWDSfx3rialxRc+Mpa3RXQVNqz05SyLiP6jQkGWXS2zesCzRWj+xv
0V1IvWSg8ZRZXXBrlso9PL6pAiuC2NQYkJP9Ea3QNnR83BXIijVoCVlsCLSo
xQuuMQtMQzWBY+lyWTNbfltG91gkEYcWnOHN6UJeNNo3/JQIe7l92eZ3hK1W
lmioMSSklWi66RUiRzrLISmhejk3Sz1zraEYLPC5B+Qxp5SXmraFRbACrdVx
WoWWJzYjQACC8I5fyfGi6SjpfnqnB/sm/8wbdzkp5zKXTpCeETJ9a0GZfY3b
AQGbCIELICKvmR4E1r/KBMF1T225YEPBizoCOMPzFEWApnxjPN4BM57rmE3s
JvGf78CyKfAlJ1MtQJmt+oT66VMBpY/1r9kzcq3cTf4qrPFta0VNaxEW8BKj
nXUYXs92Ud3IZ3Eo7zB2XwSsU8N92qEuxxEfd3ZBG2Ew5RHZ2e4k47hHd7En
go66N7ohdwpRYIMgtJSUn7rWwwsRCvVZVogrvq0ZE4FTDLReQSjodLPxJwPU
++OefkNmvfkqpOdWLzVIZxK9WUdYDIkFl4vCQSWgmvRFI929F7mvfS1QMaBv
7i5tXrKBQouQa4H9UFBKTgL5w3DmKbi1aHF0nUk5Bh9Axo8qUJRzlEetH6yP
Fow7pMgUz83ftB/Jjhf/ACoGqEpMfiTKKzmBKGufzaTzhKf7w+oqmlz5g02K
iPUog2obzynoI6Q0OsmhAvNi5BOueZl91L9w7Rgy0pJCOQjywR+6FPv71L4E
IqRpANNNkwQ9c+bJxom7MBytPLgLWF93evMjtrgbV5aVLy5uuJvKRuY6DwcA
P60tXTWg2aRGaqn77G5RAkaiXtZkXfH80MqLZgkeg3yy6P8zKeeQQo9Yqpvo
VNZbn/fmkZ0CCLW6BoKhl3jGehp79vgFnLRaSHv8JnrJDsTdL9/fDgFIT4m6
XzDeF7TsTA5xL9fUD30YfsoVDBlgBCJRhE+K1Hy+eGM1JkXLBmOtl/uAdaND
GtuHuFBgFOAG6Xfig08mGVYsdfNLbsAJAN+PeSkr/od1Lw39Jq8A1iPKk4Rq
xcJNXAXbXyOh5KEwbAIn2t4XHa8/+VhNqyFKfoDfD2QBSYHc8GfrBuE40VQG
/tRXRtftVc7sqfi4DQS+DGESkRjjHGPVXbuPkatCjZj+Xb11OCHc08Zm2oxc
L4eqfmv1kDIz75aZGdx6ZAfcVObo+GhYZInmH/sn6EPjCPbl6CGZwD6lca+P
o6uBSmkxxceio6iPE9ae3uWsfhNsS6nVMM2nul6/11iIAI/TNQMsOwpYyvE3
o20JNuSzyQtRVbr4bX/9CzdCz1piDlwzHLl7Ca4E6Kb3f2w35RelnKmxRiU4
acyW9o7xe1JTJTN1k79rRbffO3fOKI3sHL07GNKFR8QGyWQvGWJsWKD9bXto
xP/hySPc814Bzno6OS8fG9B4XUNlnqcECQKxTltv7pzgQDWyc8zrdZBx6XD5
JvspO5I/YtEsq4DGyHnTm0G/+Kuj36hoy8bFLfoimOLGftrNcMrf/nM8ClGB
BeWnZ7ZYEDNMxFNpVIwUawda1YrSuxzLgK7WSDJIZ1hlJYGmFI0Oz0bXtYir
AmOCWKfjMvvCFvu+Mrcahnjgzo78suejnWDQiRnt6DzFOHssoFL7VXf6VusC
kVvao/myJpBKZifFQWT6xMES4g5ewyfyNoxaPCU1LKkqAP7Vw5YXyGCQhRBJ
l1jSy4A2m/wPAy4X3AVz1j7PjeENIhjS0sRFgb3yMxUa2nUHS3WtgVEuToOR
qHZlY4z+qq7uxskAEDu53QouGoCvUwDFp4mkxuZr9AmfkSNmdVTZ/Qi0i714
YR/LxK/3XjsT2IjmTRRzkV+ci47Lg5NjDemClncXf7AXqWyAQVdnrIzGBUuR
RPDPOn/WlHb/1rjoO+YR5lsL85rxkW0ZinNKEHlFdaMuHGLlo6JVy4VtsDpk
QxlHkvvVrlbGSM71KwsY/D0qV528CxUavFze64pAzYqyU2/yuwvY57lA5TEy
+wq0hrvUBeiucn/FbeGadPHhEDYq1ll2N5H8wVS+Kph3vAVjuEmYRg8fKKyR
xzf1Xp3dp5N/jYHUurwATga1Oek5vIkbzmvsvzXVczF4QH7S47yDO7b2kObg
Ikyj5aTR9+feYGuIXcvrfMROu7ZaoRBqkSe/rcicrKHP1FTW83Vvu9DzAQRW
VdMWzIgQ38Lk/cMqXIQf0rHOC7y1zVt+TZx7baUE9ip1WdRezn9XdnqP2Ccl
xNf7xwbJZwBYXb4L6trhIyr0ZmI5Bqi7TRadh+G1AMGgNxZg8XDgrulS+KXS
76hIEzSqzJ3YVPUq6uTDOab2Zuwhco//miqckg7HvKEkCuJ0ir3PwupNQ/58
8qYkvoVryKwNK0AccydXpx0ivM3HiUSNTUQv2Wk7+cDNeZpDtuW/gi7CeiuI
je1vHvpU46mMig1v8aGT6WnKR+bp2cR0b4z2TCRiH9rSPeGEHkXsPmJun6yV
tsPMmYS+JWBGm64Ch5wd/yFlTawtsbyToD3oPAQiekKfav6fV/taxOIJeUDg
glE6wzoC1yC9Pxu0HU6LwOpAFlg8Ey+Pe8Rj3B+05Prty+UnuU9hwXVsd/9E
cbbqN8QsUy8Dgr+r67EercEjlGzSqfaKZhnvxUGN4Z2cBHfx7QUeyZqypkkM
0SArFzkuRil/9gbFaPkKJVNVN8BwG+xnBdAXin5Ec4WcTQbywk4pNsy6YPT6
q0WhUPN1tTp9JvPyJbvOEVHmQXxGKmmTkP4W4bkUKc2PQZhw4VJK3SXxpuer
dNajQMBRP0k6wyZVx4w+WqYCCF5tog4/AH4aWiemvJ4IWUvA1p6GXg3s0fhY
vX7gXd/pl/+pbQLF43IZSIm2Y5tSd8hSPrR42rqkQdDJEQ8QhAj/k45IO8y8
+Hyx32/3fbBVFAllRL0ngG75IUUYpxQMsFkvH1Wfef/7l2J/jjFEgtXLqcsw
cLHgQK8i/qYrr2mPjMTn8u93M8cyNyLP0dQDLsaWpKHdMsJ3H9j/Clgyfvo5
sDh7w5mDVMoKYJpuiHzNy6Cx5EImDsX5S4e9bjiCYGCdawmFXYccRsLs9BPo
qagLV1615jHUbSEBpdIyeSkEm1k8SeM5k8c144N146QBwI9AaGfjf+Z4STfP
93LC6wEL0nBITSQmOaWx00fjauEfX4sWtO4Q8wZuQHeYfsE+xbL3bP2dg5kl
1kNm/T95FmMr8BKrqBHblmR4wHZZIgl4j7x6zKGTS+EtCTmRvmzO0POUvXzW
ylPj2aKaMnQUrkd7nQQ6MZC4OKxlMl3QUbX3w1a13iSblgbtzfR9uKjg/IVX
VHJMdIBb14nxS6vuiZ5rZq4VK2fNB8IwDpOUcdR1yLRI1R/NOn8pJzzX17ow
TprvjCWT/iEjygtR0yVIGPTx3lxiBmEOGCd1M7hV2OPN0mFjLCSpL/O4VvrC
Us76YmJmB2zofHivvVaSGXXv+yD6KtN6XX06Ip0cazhEekFHpwloBIkWn4Fi
5B50kjL+miXCDaa1H9oTZWPyOI/GpEAr4WluM5pInkau0th54WNDUN/2L9yc
cn3korlm7wnP//9eA2SAFP3ob7EG66Rxyk73cyQAcFVmixtevNM8mEET/O8H
2oZ+tm+WBCfFwZYJhTdcA9q8a2LZ2C+rEgwYPxOD1ghNoMJuDH9Kj4d0mjKk
zs7LSkCYSNOvdHdVJ9LeW6yS66pUtGlhegMFaAM00LbhvpXBcDi99r+n4jD0
g2OS2bo0OLR6acU+cu2Q+9axxS1mBU8+NjwmXNENZ62MRXcHry920bPaEoKi
aql3cymqcaoePF74kRMfqCloSNJOTluYstr8ZAUpJdQgSSK1cbngJr6tqPMp
1i8ItvbPneYeY2k3RnbOHKqJs3Io/rj3cxsO7fZZXMWUSCwU4gdVBjTam55P
qitfHrlvB5YukF95GI9KjMuRr1ZaC4rZSc2xBXIVv+LUOB5mWnFmzWFXOCvX
ggRZe1F1meOCL45ool6bfA3DDT+KLSn5kAWtjEn4N10TaR9kWqAwNfK9QtqA
oENQtxP+L9Nvs+l3La8M8Wdf+dofjRovfB9rKn/hlTkXwMnoMnYX2XkC//2p
5IDxnVeLjes86nwXuiCFaAsdlI6kQdar5Sijf6X8sYmnjg1RjkMhxXmed/rN
N/Kqy8bS/nuVphrKlG/qW6G/9UQVx8rXq6Cho0VRlhuFyARegUHGLRFjo0E5
BcghrT7g3GQVR6jPuWQ6C9HKHJ/+UDL8yHftGPjFW3Fmpx2Kszq4UTqeLiyq
BCHFMP0DsLCMAARNykB2gJyg+SDCm+EKXy4khvfw86TcGIEFPiGyD4MVp/qd
w6Sh+Ttbgc5X6+wrWCveisgvbVTPzI+cRJZi1thr/QtQzdZr+CneZJ/qiz9k
OW3PujjxcHzQr8yGJ1aNDe09kEknXKhYN898AIPSQ5Ftbd/bkssBItZJiN+O
SbII6FTEANm9LIjm7d2vhl/Sy9BVH3TjekEsLZ5W5TKJkwrnnYPzAKhnbn29
jcxx61Bx3m3em1XP95RRIteYCSoLoZBEkS277UGgmO6m+OwO60Z4vIimXJzK
X6ICGzyj2z/0mnzqFRDSLF9Fezlkqh7ELrasQQDBKOENUew/+rHWhUXl8Xnx
REB3QKD3uH8jDMAiTPbfAjh50m33iFALaFfphdY2AXvM7rPw4/uFcHExTGEy
E3vU/P3wMod8WygOOBYZWt9laokdmDlJCde7PifyJdOKkLhKNXavn3M3wgw9
BVx8VCr/fvboe1JCnUHeS3omT+NDItvOM5uqtVAouHSZo8RAoIGG/tZ7m5Af
SsOBQ3sMsxpiLJ8zbxMxx7VFYLz+gmswlwXbtFE565czjECVK4hK5jSZOaMV
wfLBWroHknOH7qKOuFipZb8oarPc+Mamw7QqMQliBsRyjqLuC9V2C37rS29Y
XT5hPn/RIrF3mR9lkY4vwzuCsx2pgOM1eoo3juBO+3+tt+zCHlAMgekhb4pt
IEYr+ISY3aaX9Lt9pEghpYRhu0qpzH4GMYWFThB3kVndoUc2nOGOAwbDfjeC
N/X6iG9cAozCQnD1YRVcEOyskZ4fbvzisSSED9261RFGmZUhBs9tX3LF/jjL
7a3qAdt3WdM3KHZLDv7W6vmmmEQkgDgcgrGWP/nOrMAxKmdq+w2Fj8OuPRnI
EYcg6cbb3Ny7mJLaYDDnOxbjrp6Q+wFkPVSwN+btWhn/kalwtDS8uQEVmcMF
1PJ+8o/jbunI6hTIPh1kwwoCbLGhL5TQ+gvBj8NFEZwfMdwKpL5m+fviDjZP
kXK+lGoo99DeNXd5nhGmjPw922JxJLiI7S+NUEnHkYZjvcbE+pwUEItjkcvj
997V5/WJG5W6GfcjL7DUp35TydLl/BKFNAzOmr91vDOfxl2vLSs4JbLOPg/+
gTwWK4MFCrznb8BFJBnUuTyz5mUO7LB0gYK3CvsSyIWNfBTKoEIJ4t/ETHRW
4obKb12P/JpuQQb2dGKudS1pE0U8EXpAkfxlKogphWNi9Ob5R1m8tPUSDakG
JnQHzeeX0W7hFsH5o86Zg5SDrDHHVgtoD0E5uj2f8TCCuPKM148oLqi/7E3q
GxVT8vh3ni6zXPgkKpqVxZ4/rGGPcUeFYsAk5q8+EHuQJkDQlZfyQxszg9r6
zw6RYKeTp0xlskvO8n15b01c/Uqf96cRA73br3s9bQmdyBzxUZdS0hOY2/rS
1Fui03d3ISe5cXcXgc5YxdhrgkJm5ct9Aa44t9f6SqYf2YwxmE3GmrnobCAF
FoCZJ1WpLNjNA+aLYlYiAs9rqPdnCRCBoaWjoYsNTjtqVelaevQqgIegq1Hs
RFSW8cpxjChBg/vebbT8Ca1wCgTiVUq8qiRgN3MT0LGF2do2RgbkCG9JNHGm
8dVzYfEXAYWl6si2j0qHRnbXqtMHHmaH3TcZ9d2n0K6CIeyZr0hP3PYhSdU7
k9DjX2L0ZLnoPTZo4c6oGa/rnAv9ytLlu66DrFVYZA2E5Nnwq0/rMVC6ENB3
Dk4x76sxo9kDv46O0Sx+vgD9KNmZJiYA+g5qFdlb8/auBrFM5Kb+Lnh0aaMC
wOxpWFGlu7hBTtl+Y4598Toy52pL5ltHOO2zuND75zjsWGDW4i+qGIaBsBuA
i9/MxHZ8MUJKgc5hTVMQErJbY69NhJbjv95crmGLzoq+nCdaaqhRiY3IcpDM
hYT7Z2OPgUbQ/f20DL8v+zS5UYBIQAQHHBVHWFM6jgHLIGP9jG6hBCfSuOfr
RBWP53/JbO4wcxeQVyovl+btfIZG/SHrEo4jsuPWIbLXim7RvyvFP9WH9Y+m
1g2ThaINyTo6jykBUkDG26GZThySo5upFb6xmmgVAXqMTi69RO89HqgBV3EQ
6y8NB65QdzvidNE4Y6IPQiYqplQHZyTwX1HJl2yLuatpTv4PMmsUM6EZfK3l
sBMYadvSCUwdRC89PjNjICovo0f5zltnjuniLlDESxYvGClaCZ2wks762qKM
hii2B6QYutfE7aIfpW5cCtnvSsj2kZWqaIFEW4Tw4EJdFhQ6cHF8oITtGJjc
e8Sxu4zkeSg+WgkwXxg22G0hRpLkelZcXWWebViDW6I6Jde+FAudtrSh9B/E
Vhl3Dy/zMFuOs/6UhBwgX9oqZ2fY/veOIyWjPfzVaW8gchq7j8WfaNNCczWC
Mam+s2sofdMUuklNTSSKB6FWC8srIlw0PotoWCTyam4ri30E3FCimvc6mwOw
ZqS1NmTRCal7FHOU3chSYO+j2qFOEmc4RaHEqg8bQqFlg6n5EDWe/Vcmakj3
5hB0MewkHQ5cAMSbC37CVH6hfRQPk+1ulvBCvSKEZJ5s7W2Cg2NfitB8+ZDE
HUY7RZaokhdM/Ako27s1PsAG7gAPx2lkAKu/MxuGhJrp6um6YHbxt7uA8Js8
+ef2SWHGAeZPYScsNYKxtqNtYpGoq3ND03Z7qRMsCWBjH1XkQM291cCWajGu
4R0+Kj3JmLrSHk1auhs/fCO+wxKLokfKq0v4Q7iOQI4wimLgYj9JeK+VFQN6
noPeRoYYZwKfi8EC/xMPzMJ59WY+EOXhi1evQaHXYLFY3NxLi0vD7RzCCI7s
6p1aQ0wZTZsrW6WAqMxrOdhZffX0aR8y84W2IKjCWR/vU6J8Kc0ugtWrSryz
Gzeg8CRn18p8UIrsKRjxW0GcWNFkzBC7oAL9xvkT5FDgGbEjFa7UTNnhfaIb
TZGSx+Xvt7goZ5+odOystS/DlI4hchYRAzJaK1P5Qn5wDQE8auTQPPZKhDyE
lA497H6iC+VWdL33/KNhRyliTfdvPqsQErp6DQ0hfHHX/mSifxKPhNIbf32S
CWuemgrCD3zLaYASMyjldX7AnGWfiqvTow8gzU/mgVojLMz9IlwsrCzBhNFc
cR+nshZNnpLuG4QSgN7WjgBs+iGmGy5QQj1zQLjD2L0E6nB2ZmNXMXj7CVIp
9shg2ViNs5y6/XpwopuijrII43NKH3pD9+F8RQoA8altzN9Sg5U4Y/4kLdJY
U5HwBHQEL473ChwNKAk6H6nBf9jZ+kmVxrXnXaLc9fJ69C7pif8/1t/r6QUy
cUhxcicITddziQsad9oBbp34g7S3trjtnyJR681md32MWapcczaZ6DuzA5FJ
CsjK0jNg8ZS3jRztnM4K3mQy1DvtkqqSvBATMtZA37wvVMcuh2+hDvJn/AuG
l4X0Kn4QovjAfQbDnvt+6QXsFEWHFSmD5lT6Cttobd3BlmckqiSV1v5bypNS
F32yTmXIpMu0TR8G54l8y3Eug3jyjLD3GLbVGd6piqe9qhBncwf1A5FBAliO
Owr6QQqG1kVeEYTSysKs1HtoupKCElPlczUDrRaOWbA33V2IaNTrrlpmpEP3
Ixb9NA85f4BO58lPXWSZoYFE/WI997dle5D6WAyNFZOEoxuKAVLokdORdIkj
cg6MGLQkLlWi1dX12RrYJHrg2s48iefpsHIsEfGQJnhNssngnuloEHBoZ7x+
aFVnUVz8Zy6wgCB5ByGITxhG8N++GSoGuuTIDdXQoE4lmND8WmdIigq6NFxi
aPPqhckG1J9phQ4jJx/uu6oH2SXT1ghQyIOze1iziHqWU6QD5CI+Devj60/H
WkLq/CkNQWTAF9xnhGK0606DPJlSeQ0CqlhJEy7bJrL+8qoRAYvKAXUYAQ3S
WsX3qwrEHCWaIKVlhldBDf8iUAgUCuZEYBvejdvlzBsJJjeA3RWtdTBrEWdD
tRrREwRFFjQr7gwvyO+PEFTPwFvppq5iis6JA7IqcZ+WnFRGFq/fk8G1jQkd
uqhjH8WGPUxD4Xl0VEx83DjL4S2Kl0UmuqoYtDYN1iBkFt4M6+1PFm/AKGNq
SGtGSIukyKGZGEVMm0rU9gEFFfxy1lcHqZcpY31qrLQEkTnsHkflgHAaueJP
6YNpqg4onUcpJNHqqZTWh1jY/X8YthBqJ7O3MGsChNSKdtDSR+2Uvvd2hcrV
QfAdW82ktaiej97e8cK2yTryi83CCyrIubvGiN+EmRrXjCppILFsyb2DfACE
um1JQt2jFqgpIfIhiFfWGHXTRVH3f/dmvNfxIjmUKRdphfWsdkxs3YY6zd3q
o8QAPPhUCnqReS3iF3i8i/tkBVoEWAg7avSrp4sp2BWKC+u+Vl6DvbH+E2AP
ENdULsZF+P5wbUbkARrFv1sK4NTjRghvbsjE0x2/wOdkg5eTfwPdpEGYU+hQ
UidSEA3cEN02PbgPcAtHw+FI3uOcMI3z9U6AJ7Oy47kYL1sFZ9DCSNnuC54x
HiVlkjp/bMaG8pqW+V4Mf5VJLm3zcbj3Gn62gsj9GFWEN3uIxNX8pzoMVrvq
mbTLPGCtz54dIdJA3+Cpc+OBTesJClyFo4Xv0OB7yuqTLx35cN/6WE3n5CSX
2mFm/vd3990m4CleJPnCg3aY6dki8XIVSJ70ZD/kv82jKgjK093Q2yakCs34
1qav+165ZZqMCssqwAd7KE/A4LQUZa5wLBWGiuni2u3tzPAXNaPXrR/NPlVg
rnLkOnORdFGZfYQV0Hc59zvIdpJv8N7qGgkKxuJPMpBwzjrTguU9Gu7hpekZ
RyYAoSNmrokhC7DHAYP9j76yA/KoHorXlNXE8d/LhJdKvJqHiUwOV2SnHXtQ
ML1a40bOgoStbVZYtxdsPLeP6rQzIY95niBYHwmkCUpmmJPCi1dlqVljOdKI
P5W1C0Go9aqUApjeEG/JmuF2HGEIJXA+gZpL076rblnBru5gwECpccF1t/Mc
p4ZyB/oma7XFKOncCvlHU1byEmCw3AfiONalkHwkHu/lpwUkUqYkMpdBDMyG
jG+WuVK093ehRtfRl2AexJMXTAcz00+Dqd3NxGexD+cNDzw2w76YFGoSIWrx
HzqEHscHV9oHP7vcP/nOrUqihF6rKTcYxZmdeYtoaDoRiiRIN7Nrrar0hrG0
Qe/5jn9S04NjuFcJrZiTqiP4kYDtJOeZsGvugXVbuMi9mvNiyia6tcguoO5x
DR0ENHx1qcvd4fxkS8k6dWVeN6PmIr8eEdN4Z/WVap+WHlegSzjZ9x5uSaxv
Y3WIn7rnP9tsugqpiR/WikWj6F3/DafykRxf/2J3jY7+sSPbjAbklrAUVKCn
KX6UKYbzfSIqSeM46a7xDQWn6Fn3/HqXKpNEuxH/KhwpE3PaL+nazyqgk17R
+60F4MIQA6jumKrt7anY+nprL7trp39UxJ8q53pXOFScRLH+f6xym5ub9CeZ
1aTEmW/LS+G3UyhhlU73A/fl605Lx17jR8LAi5Vtkg5RDp0zQGv5KwIyQDL6
FP+ejc87+ur4vu/cezlyCtFrHjrTfLyskGv1BuWiSE5wOpPjRXm5Rht+A57k
fENo3K9EcPjIz5U3gQoHmdYRi+Sm5tl7JZnKRvYKS8aU6DI2YBRWmaAS6iWm
vc6hUnJEn5mLt5hU6nQnR37MZqoCGvbqSER60QEA2xsVMM86fWzwJq+NY1qH
KQ1ziKGI2dt1zfZOTQnCAaeVSzqmMh7CgEJIDXtKy55uiJ/ndCRBGCTyZ/48
RAQ+2xpFp2RZ0vYKQFUVMBgjaE2YThixP4P5/1N1c4Z1QWYfQCMDOO5Ab4aj
nuY9UeFM7lmVVhZbc1vJ9cKlgV6CWsXOZKuIyxmXd2+si9PPyqI58h8811Sg
p19eKZESvA4pLM8/dOo6TunZlmUmYvsJWfW24DU7JX1lHLAYs94v85Ew3Dcl
+5icw4zjJ5IAy++GS/nln5yk1cRr6eUsbLIoIxLFg4VpzYibL1Q8C7rY3l41
4/AMUSPukW8RTRubGDNyw46Hdeaeqjpn4YP2sc+jdbBuO3/NNOWLAk4g2neV
hzv11XNvnRSfAomQiaCmnvBgKFEaXxGUGTD0ricyd9VemQN60w+iO6/0tiL/
YOQm/diBg02SysTBcAeG5heXBUEJCF1b888X0xuT6kSuyUJsOyoHx788FXAr
F4abGaczgCtOXPT0ptKJJfwzbpNu0HQbGNtRj7a9fskyjWwKxR66we97Mxva
XQPsnm881ktEjBTzUYh4+WyGIybLAZLK0sXurF1TnoPCrxZVxN/6+ZDC19X8
tve2yEiEkTk7+8vYOqV4T6OP3PA4VwUQ+UjTpnJ4Hnzqlmb1gfH36bb/ZIEV
JFRtDm96z9Y6lU5YnsSnDWHMeB47lHyEdd4Cuq9/DKnMN1C22M9DT2+3xTQk
X67YNClRbFEgR0f4x6taSVNijH0anYdKYXdiwPnWE8aHu1/SQd3BiylYNeVF
Si1XtV8TLTZeHJ1fBrKYipApl14GPZMF38IYubpMT8DOP6n/1ECHt9Hpl+4t
cw7rXwk15pK4tCcLURX0d2Aor6I4YTzQDnVwEux0iYagEe2QZ5xRutZsaQfA
vbAYREsUaE+TVrc13kcPHz8FJxd9cJKxnCFblqZETDrKyKMPAJfKPUlNr0Bq
PUr2jVUIxI+MGFQbFM9Io+dXFLiOugge3ppzy9Ffajf1p0H33C1AwsoWySqc
3bPdR2+RzG/EX2s+Z9mwQMQW45Eqan0RtWsdvz4xK8i9OBPz+QIzPC7RTjFj
mFPyxutvx0wtmsxvQz8V5OFF7GLYEKtoXzo0gIlpOJhPj3oEHCNKlABy/rI2
qXwqsUY/6JtRVj4bjZN2oDjn3m/E6UpZ+FFnKG2bUG3QYPUIZvyK7BULVGT+
FekpsNNsYYrksC6sqTiKv07btT8VjFx5gIRI7F7hH43jzVX9BlE7vYg7QPHB
sX7YOD+jm74wIOSpJIE7GXzPmZZ9Ju8qNJYGTHDSyEoH9k/LG1UhaAdpkU9j
SGeIwtWM4iGW80/hZAaAv9domV3NogXk9RQku4W8AuQRFUs7Qoo+qaFSwBhp
+giqH5G/nKfH4ErVgcE8zETNtF14a7NhYSaYM/6Y4XcIuC9ji4YIbCNoXmJN
+na+3yn/9/na/b2yC7y3egi1fj10S6xmJ6bECQhYbHlEhldTXDP+db46N6N3
TMfD5Y5nqjTtwZbgqd+1zarrTq4EceSQDNZWm3Ef6G6hd2t1OWTvFka37cux
3GHXLLQ88kMq8n0xLNOlurZFB5uiF7C4M+7MFjDUS0Y0poDhStHHfR7X5zwd
l1GaJcY5NXcrnKT1mh6Wwggg1RVPQcHTEHq5VU/PCF1kq0k18InCGU7jsbVS
IZD4KoCK9fh4MGlnyNBmN4G/5YNj2U6qioFKTAC8ytJe+4OIGFOKIXNP5f2l
8O58cjCRrzC/wGdBBWizP3ZyDqvaMhVkSywazbYDOu9Gq9zVsO/UlEx/vZDy
sajJTO9D+9KwkV9qQdCg8TkME/0HcZ1Ras48XQVbMxEYTg6zmfyE9P4wMbJg
Ye4anBnvcpH/TQWdtLh5OwxliWwRpqrZQfwuqdUSO6YxvRMtD27t62Iejo++
GeIGHwE+dXc/Yw3t7xHL/XeRDuGL/jBcAgDuebF5AYB+cs87Z6ognXCWuKDG
Ey0iKWMTuTJLpGd+7Sn3hKF1MkT96MwYVZU7Rvyo3tODjoqv/JMmjo2Nazx8
hI9RpEl5ClmHTKWyqxdkQW/QOv18oyz9qOR8e3i0wbco0yJAAMLur64hv8n7
IPO2cjk61b2SMB0ei3EOAVKwcjXNlpKHyfYSo4KGtnk45CnUD4UjMeulnKFJ
z2iCa7lGQYL5dOT8FLswVWLJSJriWcgtNghse7D6hTdNMu4Eue58AX7bQYU3
oSM7b7tzrPwffyAtX6kY+keQROftro0do5weGwjW6hXYRmuUXRRqofzZX7iC
3CMBwbLd6xiwzr3A0+z8WI3LoHd+uZlgHi6+K3RKNfcudOnMqHRQiym9B0zY
nGwYtDeN+bkJWytmq8DHdMQvqVI8fze4EGW+mvFF7YjpbiL3AlGFtx8K+zw9
DAoDofjGdNEX1Jpk/RjxQhvK3CYrlDOFiwkpQVG6xGGHd+tAGHr5tzg9xQq3
yUJ/YVZDbI4/mJGeRZc2nyQMz22eiuJevnzOf7QqnvLoWDmbTl8Mm8YWTAF7
aQDsaNI07nbRQl45R7eV6oGEawEDmA8hIpgEq6TkXXUc6Ss7PV+xmSBSmGo1
lvAY6aLKM/O27X7s5zEhCkxt+61Vlec/qG+8XGGomssQqC+SKu5ZJs2yUJs/
OCddu9hEtKZUKkscojbgIN1Yv3cTIw/Yy+Cz7Y2Y0dAvvtLp1ELj+SDRFlV0
gvnWU2HUslzXyJYN7+FeD/rcOi8WXeKbZo2Z3HMt6FYMYg9fp7ctSmTuCqdZ
KFzQT54diwJ+cZhhQjaweadngtmmulykxC71XTOniPgmkAgQeLApNqXRAUCa
tUreWYDs4ZYYExuroLiQYnZ//r+yYKS/T+s7rn2v/6Xv8E0xF62UpyYpbAFS
/pH6HTyFCnjZ9CiVyjiMxlhgiXARD/REz/jkEQCjjgr5JleSLCve0aXicDxr
+/QGSwTmEP9wa1Vk+HhTFt77FKIloIygGB1ZGrbRo6RIABUVeuguYpcpOvKO
l3M8tvhmB4dmEJ/0w2iuPLNjidjbZEOSkGiVLwdDbZgvVeyuQh6noWvgE/xI
HzmnASzY2t9/j4awlu3dmtsHQ8PHil91qLULop8vyqCvKP0a1VXDmpp+B56u
F8cyKok/RoKQladbixPxg23t60iP3lme/DrG/6Jx6HWWf0c3znztAOxDuKK4
HnJO9+XptCV34HoWatO+U+QOAxNpp0DHHPe5OJ3OncvzwpNMC8MhFeQbb5tb
QOaYa5n8+7yYqzhB1BsCZWDtxTalKLCBZ5ZMnATW4zZw0MxaeYQw0S9MpShB
hv7fSFKUp87yzJq/N7ltNzU/jARRES8HtCkC0ga79x56wBJ1EwhGFxgk6OCB
C/FuXudkOfp8r8whYtHagiEyfquM/Ki6IEVMrlDjaZoB+2hAiivx0aZOiI0B
Fk6Pm53F3q+cZWT5NvngBKvS8Tfvj5vi6tck0DtBKJjeEtwu6MTLuB/Le+AF
/LiPZLibGp9mEKR54iLi6+CQi8API1z6dl9wcugYmBhBQMCBhwF5pXkHLW2T
aZkJi5dMfkPypPQGf1e24qUCoPed9p1WV6dhMRYMHkUjDLVHl2AB2OJ91uPX
AnpjvOFL0Z6J/gf0MYR9mXJ1FoXJ8WYDNHMGy/9zausKiH/rXsJ5ZeG+egYJ
VfuPCFEirBgcHvazDVsovxo0wpbXTcphRPznvC5iJe+FZTglC/iopbBvz7GZ
W8i3cnltCNbL5kYbC5em8lWKH0sEq3+zuNcTcoW7VRe/VH3MwWSSPby8Wtkp
nq9OslWpnYeiTfwBVJCWyJ6VmCNGz+LlwDc8aCfbqpSayMcvlczDn6DzXY9a
GWyFu2xoSGnP5OnKTc8wgc4ILhXCYVbvJCXMF+maIyXHnDYiCyZTuol7tMUG
zZ7adauSxTPmXds2jF66ZGeUzogaSpTO8O4RXTwuShau98zK6jMPlUSpcrPI
JNGzF7uLattpVCRA1iKRUFJCoeEM7EQ4iJppntBHSDxMQ/TLodAVjA0syBKA
RbB78x4Eeb2sb3RchMGQ9MPmrvfwGpR+f/0F5c1xewYLN/L14/JyPgYFoybU
uBFq9/z+SJpZ++d5sdBWOL7cXWCHTvWakuAJ3MfjiJF+/DhahYTqdAuwHLez
9qH88ZAHf+Z3sT0ldq8aW7MxCtlqwOiO48w4JBa0HMWrtVbycebAHiPyAn1f
icVwZ1SaG2lYpa3gZm56BHP4FC/n9Jg04r2qhDLhTAbieJkXGSaV72JrgVOH
n0T2QzVxW2bWBV1GYRJmmzHPAg8mxRBLNbAzfj9OU7/nPjp+yobl0xCUhhSC
7R4sbiNExkLV+e1WXRV199gdZMs49jNAYsPI2jZe6t0/21hmADXoLU9KL45d
xEPyfkeuZsBxYvvMMHuEaO0UCGF7SHLtOiIg+6AAva5rZ9qxD8fPsv+b+k6i
3oHgjj3OBstlG9xxza8dA3nUeNZy4LbB9u9NQMmfHSpjl3rzQuPi9hVxCXwj
aFZX3QmLJZHXz2/1t19PBoy8qGOoNJglv2yV9aRn4Mx0WaD+3fJ/rX/vpBTH
iOyiXIRHWkxMhM+zGpilt7ZzZlRzRcx8Kfe3z+YPUBu/e9eMykhgTHQIVs7m
Fsy+eTkzBal+FbUnFZyFcd1G3LFddTdcTIZCK32N8V7hcgUhfCheqxIe48ao
UC8MlN6W5eavku9PW3UPbMnPufjA3sRnPiTVq7afC/xPlXPv7zMmLCIQasFi
TRRHno7sJosQrLjRqrsyGvvkXi9MdtvkTg9a8AJs57jfbSSfFvc3wWGF8Jy0
HzvOt4Dx2ckqXkVnvUBFHtv0Phh8s8WjH7UgeAXveXVpo80bj7cjHsP6n502
QMo7xWK+c6BtvbUg5t2mxNolhr+XocburzKwzt5YsFrGa9Gv2+Cx0xH7l58Q
4zL0gr82+YHEj6TvUmCIlCa8lcSTZWmrBwh1shV9tPsralxe70IFHqqiJTu6
04mQlySm13qVGnUhvEFfzmvF1iDw/Y+EaWkVkk/4mTeKBHdnvT4b9qfUrXP9
1UoDn+gKA39flAWU5bPr1OpoTQKmPoLd+FbYNvQy7c8FbyyxVIg0zjMNiy2x
F/OBf5fMTue/I4vixLNvOdjTIyTPdbMxvNNaxv7vkcNOIQ8vUDciD7i3cLwr
N9sZrwJilCmNmcdRO2t6TvQn/3oLj478MIkWMrnBmnaPDQBQF7kX6Dbj21iS
GJxmdEj3WR5aj+rjpExpIbL4GF80+lM/nZSTVQtPNGrHm4io9v9NI7w9hy/E
zc+PqRv3cV1dd8+H9J1isAytQvFpWhC6X6gyBHwb24rFEI/SF0klyITJS7B9
rm4xqnRnHD+GyEeE8s9wruEhK8gaBxJpfHTjWXGMN/IUyT0IIyC12jCak73f
AqSbrOMwtNogaEFlzaJX/m7siVN/cn9rvpVcfug3NvGvwYq2Q1Mymev7h9Bn
UXIziCNdeAqdsLvEoR3+U68YyLRAZK/ICvDNr1UPpZ9/kf3ulULLUaizEGjU
Rg4rfSp31ws3NeeY+d5gROIP5kk7jBhs7hgL22vE08quNu/632SDRr6UY5DT
nX4D0IgYWnRVgtZZGMrC5K1MnBox7ta+b7bYo4zfcvSrhaYZWKWwPkGxvojq
4rapIHklm4qVXt5Q7FXWflyZxrNEeXKJFjStHUSAkIqG/3yfT/1DL9+vSYeX
baqJqgzOKCrzRGLkexmE5lMMCZelAk2kyOlv0S9iADxmGERuh0AD2hbbe1Xw
XYJG/a1OL5yt6nBQRmXkn2CH0nO+/XaX1OcWFsfOxJlMO/nLxezE6/csgEPg
c1wP0k5LgeahzniTIRAEFW18Uy4phrT2NQv122uHvO77ezNtwPzQrqznUuOn
jRPJGmCO3k25cJ5aBpZK7XdV9OYvw/IMlkGibjI03FQ40gC+rPFP4sWTT51v
ztk0FoV3XDa9LhEA8WgBpmbD7vYiV94tV7/exF16j/3MD92pBG9OnO+YhOdO
fkwcP7q5z9WmyCKWvnhz7fo9VPI3K51f9CYkHH3pXKRhVzdGnRbJr0zuvftc
xOwPq7N4cGa7iDDHJ3JIba8OvZBalYcLGk1zbNOzvJiM8FmFLs7WYp48xl6/
hkZB7xFRVaNQAWEVfC5I33m5I6vL81geRMw6wdJaton39nAIxGNnam+TqW+g
J2vLS+qTopIklCXlG2IQpcTYIyHxbNG1pjxYm97eqHUR4jcMgdcJpF/8sdHr
rlCQP3FeaBu0vOqaas/pwrY1wZEWBsukiCQHW71URDe1wzPdyJoXAYyyHbBF
GGOnUAILRMv1u+fdn44iaZTQFs1xb3zvDxF4kO6EgfmySlo3L/fC2QDiSJQC
3JD+96ftO89MASSBe6jQdrFaebYySUSPEBlbeEUa/3k8HxUtWGhN3z+v+Ne2
pbTvu6LXpErqjYAYHfjyg/TmrJSTNLCvwxECYSquoqfYjWR874uGYFUh/Neu
7RRd4thWdKd5+Fgi95UGEfrIW8rMVgWkwe3p29GXhCzHS5rMJNEGu9lffYt2
xtJNzlpOfq48y8BEwT5cgxKTu4M5u+FYwLqX75xY6wqa9Nc9l3zFxPjdn4Rc
9kIUfB7SSq7KwNGYaz8IK+jOjrpkfRsjtHHG8SYeX1e6WNAvHTgvwo8zkDVm
m1RbVYWMj8UYONmpiH2ztg5uaP/Geweg1SkZwVeeG5kEyNwWXitbIQEDRYgZ
XiYtAeJaNjw0aASaDfUiTfbbWyKbqxEltEZWcmxu6cj7E4jcFzYK3S8aGN0s
LYjWKdelHMD/YAZr7rE6B79DYZnsXj6Cl0DyF8x6VP56wr9T3bnIbWfe88q9
kVU0FX0tOrxqq2hU3lft3YLrvIBSgYHtxmS1/crH7EfuiutNcSrcJVpXu4uv
jeRtNZle5sBiPnijjpCiWnaLy9bWSPWaDm5EKRLDL7wpheZzhi4QKT+9Cgxq
tw3oBSFl5tTerpMFZRKDiV6g9fOpRf8x4Px/z2xcZObH3ZAiuVW/DP5WxT8+
1Mqteh2MeyLVp+k/40dSUG6bdKC30g6IqMNHJDZiyqEnmLft0wmmkn0R6vk8
OIFLDCcS9kL11xDH8BRP15jPT/BHJiYf5iSuQmL6n0PHkl6IXNC8yX8YSQyk
mdllLVlg4DEpjzXePovmlqB5rYb/u64pkoyxh7uTinQHBcgR4EHctSAxmM7n
zhRUg++D7g+b4SGirG0TNEhkOsCuLVIL6J8eqTMW2pmHrO3b1CcUE1MTXudq
b361JlFUfJZKgYN0SJdq+DbehaSjNT/HH1k//C3rDoK9zgdMjLNxTf3PT3al
WlxHIpoFitKvt6r5ANOUH1k5+YJQHvmGpsbAgf7w8W1ttqd7/iPA49xERbLk
Rj8T8k8Zzsy+aOSk4Mk20NVDW2FW+olm023t8aXs+yl8AnYBbHB7Okx/Feji
NtmRHVP9/WsBnLZrHNVi5V1w/xp1x/csIAF9HtP2QTb9xdwGpciXV7VRBxu8
H0NiuIEswSWmYb/Tl2RgIjJwvhVWe8QuLqWBmpfXErZtmbeLW+UfHeOOHBtz
DWMX/gEuVx3kr+nI9C6L6hnfTVMjoMs2xqhqU01lHgejhPaqI/WEflm4pyGR
6CTwHBcn+bSIx2Z+FX6Xj766x9RS5uvCq8n17C5BiwlRHyJ2ei0uT+SDay9Q
7wsd8B+19uQAEiCFXlSHmOnyc7EmXm4DfAyCYxXWIY9YsxPVsISM4giSXSGo
VuUlWTtA9kDMGRIpSdESl/30bkZdoRPeF4ENm25MEvNVv12vHrJ/DFfv9nSp
UfiUxgFbxyzhjiP+x4QrwTKnxLtovIQtqrETh6SFHi9sJBToFnREggXpxKVC
KcD2ICA6Xik87IuglgmFBG/CGrZ3e/YTFalmk7cbBQ5EZN5kPl8wSB+FHZXk
x2Sk/i4Ive0GYXzWCqy/BZ7EruvC8C8Kc62kOoe2hMkInePGKuTdwREg6wkH
SACT8211BSEmIQwHOKA0iNMWkyeeOVDucn8DOyB9TFjbG6hJMjT+Jj+YHjn+
eDFWeSvo5F4/fVKF8Z3g7R86HSXA1jFBVH8j6Tm4K4i/4hTp9fUNISP4NhMp
K26WKhn3TWHvSJxTrjuLBCeewB3bLe9kvwP3uCqA5TmHLSZAieBreXz/fbK5
PeV9FiYqFBP/7klSuy/CkSKrg+x08u5ZgrwZG9Yob+42rIb5sZvCqPkQQEJW
hzbYt/JJrZhcak/dyF17xDoudU9vNZEtoFCGWdTHzwJvLInZzbed2L68rra5
ReDs4AYCSK61kNOm3H0v8/1thmpPBCDKpA43cHM6onkSH0cPJAlOX+uJEyyA
gROfTm5Am5GturQ3mhFcmrt+wCT3L8TXK5sNSb2em4mNKD8hvFLIuR9L9MZA
sGO83b7X43RIVB70VqUm9X1bJC2INxvogTRIFf1ySZSrGBymodPwIpD5vkre
sDKCuQJNafRoRETrZmt//nV3szMQp8SGDZz/YekssvJnFuyAkOJQsiK21boK
k2279hXRblolUN2iYYL2y1E1ZP4a2GCQnDfIKIupQwpAWleWhdczfgHXyHSK
2ayV1HcI9MewrY+HJE9w+D2Pkz+iHX6TYuLw7sWQXVSP35k9vYPpb+6P1r25
IcCTiYp2ptN3Rg3J7G5u3S1fv1qcY21yVIlyNiaBvm/ZUz/J9DIzN3REvpKg
m+BGhyvEzkM+QPpwuqvvOeYu8CCNu5KZjkFWDhQyUW2fcNzol/0aWN3TPODc
vm5rQ1Eoq3C2UxXXcBMYuFh31444xnzUsAaKCxZwAfhrlzSijAZi+zFHlK/d
pP/vHxq65jzbGAcaYJeQK62MdjeM1wkCDfp79aB0OwgU3+QtjTD1jBXcO4Fi
aB3Dveal2z3XN845hgHUSaGGIpf0rmQz98RktHgOkB5HHYNup3VcwcOCh3aG
YdV7ggBVxoS+QJ94HwzmHidsyQnr6SvXBDYcgb1qWoCymwnYhOHyd6R0HsMh
kv9s92noMylL/rLbjHXxjVbSFUfHlXCbQH1XNtE8gU3nY6nWpG0Su9MtLLRg
DzT85idTIZOjgQuFEwOFE1/T9lClhBIgTtrolkZGGf/Ft5wXuMpJkNRosc5v
IytE6wTFKpzXcSCyYLl6mYr62XQbnjKLbItqwIxNnYO0Rq0NcBsRG9tgS8LB
WbiB/rp7vfql5NvlEdEpOiA9keoxdAyuwFVlVNEEAw57DeMnw/YDvnGYUvvs
aiH2HdqBgpQk/5ZbAogKKCg8VAsZlpSk+gmtrdaMVEnHlCnID9LaVVhTmLkN
jH4QqgCBlETMReEPRxzGCZpXWK48ChK7p97UR6BHi8+rvfYYIbE4c5SOyxhI
0/OYuvLUPh7PSuhjUOUic7Su7/NFh1mRfgE6w0rBDTERcV6BH3lns3CRT/fD
EBGfxQh8A/RegEj70LnXREfkXCVn2EyNrwXYEJ+k7Bt7NIyqjxAYnoSqi2zl
Du75/6Kz/f5BtxEe0XS5h6EbMr3jLcU26+L9ATzBQ9qIBSBAh/fzRl56/NRu
9DxV5hHptVa4muQMK0TQ+80K5abKcKSf00MtNQJ2b5rkSOEx43z4rYFiTpa+
l/uRckO6EbNdZ3m+JOB0rvspmByvdlqUGLoFMJX95E0P5lrVSItok6EtBuc4
jr1MgMwC+RTVmx46lOLXO/6IvGREuBt7a+9LfN4ZGWUVdu+8VILQR4Tp/Ou1
zFX+Z75RCd+SVEY3FEIR8mlCc4jzpE3MQpZiO3cgX9DJh8E/iWf9tFRevDvO
YbJdiQ5kFIKsAGhrmGz7ejYZervj3/FoneLx0x8LTailSjBWdjKEERpIiNzk
mx9ZGvTHZinK7S/Q+dBBmBdLklzGSjHdTaVuEqdM4eO1CU6vCkAk9fY02ucU
kDkBldPf8QiIDdg2ulPfLJc0mJSmKXO7W5h2632Ho6Ml1ERFA+0jS/dEZRLn
jjZ4YZXVz3dla4QfLPN+KDmJBg37PfhR4gf6T7RWpNI6UsEEj5Ba5GiVRTE6
1vhDtP9S2eAtipyoo9vyhbchXXocrZQ1/i5hRUF6W992mu6wqdXMNMdySrKT
Z2eoAK7XmMtJkWgw3/O//dMeqiM1UnYuzfnTBggAuyg802b6gTE+62rpXL5F
8Ra7A8mRTzcBSTPS/fd9+i5x/d8d9KQN4KH4xxEuzhUb6WhqamNzCVAQ23ik
Ph07YMxLvcoemM0IfqtL4GXI8dc2ztUbTKnKY6k7w4jM2LnFd1vb7/iURCl2
RX1L4QbMniJGG1PSy72C5xwUaj5pABbAehxucCADQtLhDN8BgzXbpyCmiZYQ
huzQ6cVdjl0vizeBNYkedzoTgxvoEz8x3/biy4rP0RiXuFBVSPYqbwBZYJ8K
VkOz2sap1yMhYbUtkrlXijukI6Q4nyalhaIdDYkfE0Fdye49gfO1R+uhN9XO
8RoSuc03V3TLAbGGWMvYeXsfKEeNl40yiQukqDCq7QMpk0+eyRYnLFdtPX1F
pCw02q5LF1oQVy2YGIAEQF58Jl/5yNHyXXvE9THK2h4mKPTzJvpQnkEpd8NT
U5/IkjsdmFwcdnDKQ9jlHKGOmuSY0m1EvF6K5TfA9XifM+0YGQnFFBPpz/Rm
xV6UYTmL8yfyXLJXOvySYdmi6PZSh8pjw6bohyF/GjPtBVtjdVgZMBOZ4+Zf
6AV0TFN8uxuaYbSoev7lSglPq06NQTc9rZAgaevTVgBNJjUyfbIwT7MQOOJO
JcoOqgXSi5blRqV/SnaKxnGa25dSqRkTV6hM1OmKFicDAXWdpPAmpwZUZRBR
JJ9Yd/9TidrnXWPCE6tsJf/Lc9XrBMTdK8UqaecwtqmcP3GUMf8HZgVhHKK7
CgyPOXJkT3zg5xvfysBrIJ0OcFC0TyR14aH0bbxPJpMQpHS2UjM0EWCXjRQk
GEE0882Bh1fgHSBbxk8AHnAVX+lBhuUv+Cn2VCIsJbOY5xviZVzOtaRLw8hD
Ej7HhXYb4fBCUJcgJjjo+VUKPkHmpvQuwdJUxARhsN+Ugn6YOzamleYLFotk
mdoiWjfgSTV4GDun89yS+2VBxGPyeBvSdYQm27z3lIVAQ1dFRcVd75B1FrbD
CE9DtJS7mDP5/K0iycWXwx+AYHpmXK34nUnoZPbHyHfXLJP4t0E8JNkVY6sI
0s326iygNXCaHhIOgrASkNMtJEeQGGuI+vtBlpCQ+MqhxVRg3EoPqKB5ZmQR
1pqLNo3s1OZkDFIAfZAWDMuMAstM3yGkN26SYKgXdQkL6PT6eP0ru16CLqn0
zzqEYAD75DUermSJv5dGPKzM/e1Yn0WR8ZwCz4Zq44NfmbPV+hQoRu0LEa/l
/ClhB/RRmmRVg0ZDtgBU+3y7j5vaUUP31hMDL6d89e+jV+Aaudjrdl9qqMiN
rWMVoWLj1XAwGzXERoSAxBPbHAYZ7zLBASMxA5DwjRfv+sjT51tYSZCzog02
RFFsutc54Th8FE+ZSGzn9e3xKwqeUbK6bWK38oc8zrZMl5HjJ7E+LX/SdSsR
4KLC6SuHmW8oW6xJXUcXtESdJ2/5Z71vnKw1O9poReKi/M5ZmwgPt1pN7FvS
VOUML0TPYIo3zT+i5YZ+ro0XWP1/krNCMBlS3wJOeN0hBe34Vrz4/ezyTnux
NVdEymrsdFlmBdySxwde4xqopiQxRzvqy9vmyKvYv1RobHkfVKxoBCqSVYc9
r1eVK/AXdLIdDtctpQNXN0dV93qyil7C4jacHDAyi1BHnHuIZ7OPK+B7Zn/c
fUpVkqCB8MRvNlyj+ivsfTx4yBV+xGaB7TLse5linUxr8Y8TEtEjqMZuHt/m
rgqvoYhWtCZiRLEf7hYpIHVXad2tuT9IuuJtqQqK/WWv1OpMidM8K0dgjj55
Bj8WtnNUM6wfzpr4szTMe2oD8lh+ja2w1Y4EOrP9rR+vBBPgoTn2mw0pvYF0
JHWAT+uGKWeNQm1f9AGGNsh/laQS7aDLrNbPi3TzBmnywZZlYtAhmWMI5pMG
Yo2NJiz5p0oxi6aICJNI1zTL/BhY5eVn9TVc9994rLqGl7trjuoCkAd8nSyr
o4ebL+55DxJf2rMyCVXeByimgnJ487QOVugW1ROP5b2dO8N/QtpAoF0Q0DeJ
cV0gVcIRIJ5dbNWXVj+qXsGpzdFl13suNkf5vOYk4uu/Ry/tub/YvjckuV5O
XfQFhL/wt9aa0jDS3J12F/X7aSe+kBBr4n0YLT+QKlOBj1zvp+9jiMzp6hjT
yDEszRfgSSE5PRO032xXirEQ2QStjrCaFNjwzBVpeff6idXMwZ85+XCpruq7
6kpNMUawTu/JekhqMQ2YhQAWaqMp6QQmPxdZ53W7++Sm+Uzkitd9P5F574NJ
30h2omPzSARQr4NPfsBqW1jqcIUE5DyVpHdvRGiwRbLObcxYUFAZokjWJHFT
BKXBqy4JszHHU9c3h6tx8zZY4F2WlJEQp6V0OxMLM38dJzoCDMviS1bzZuAB
UUAavO3qP6/HX5Bfcvfm4rDKcRZ/GeeH3sJkMZVuODxIMLa1TpaxZmc8Jd7x
2oHtJDZ2+2CPeji5zcpz5Z6i2RZZC0GrcNYx6YyO/nCCUustNKEsyjpPFsDH
DnjCnOH/h3SCc/wIlQDRcucwrMj9432qqu9Ppxnx8P4rOc22gTjNXyU4YVl5
i73NHKbxeDqzmD3jFYQ7tmg6pDGqYCLOE4O78zv8Iog2HjtdUO0JoJ3xm0OR
MC++Nygi7w0LpPDp6+aWiQ2STyHjcQI5lk43VxkON+US1aFm6akpEQWarZps
a+UknwqgmVuukF0URdNiUJ5M2/jL2f73ghdR4WAHUMxnIx7oOTvLsM2CJysb
vSQUnNOlmm52XqydgBH+CB/RVq8W08lX/U+RTT5E9/hbQWfIim5BQSRDD7dp
Kg7vUlOdt7vihNfOUizX2lONXzTHR23H6gqnD8magRlHLihAZsg3om5Gyv+6
uQEoP4IcPk+WEDWwL0LYJxTm7zuHZNt7/g5E56x5IcxYh5VcLdTNMizt1OEZ
guLwEam2YhS9z03QFgdZ0q+8xcVvZ7J3rm+DejVCyAM+ut5LtkximvLMDHCK
OrB2Z9ykEuZ0kQh8Bg1hcNlMJYHpYFTXFWLrvvOTldRFapqW+JAwWh4LAnbM
8jbZBkd9YfjmvvOWQtvUmpssoJsi0zmYTwEJe5Hyvgw9HvU9Heegu4APyYOV
CIXK82YdXfVIa5CSFLzCFtWdWpiJotfG8NY9jULCGO9u0qIkiWNqHohhMWig
2NrRIRZiCakwtEOxDCPBS6x5pOpXFJ40IXUEGR81RcjnVnDTQTt8G/Zhjw8l
Lduyu9LT9YLllZxQBqGdn8DNOj5Cdk7n9o2Ury9J6stjPjT35FjO90zTdxvC
fpO7ZRRR2zxcFpVzlxe0gROW3xCGCehj2cwfhaiEQzUHdjWi1D+g025fPXL3
m41kyT6Bx26w4JKZh7bE6U/JkaZNpmOXzo5LPGJsU7MVigHrFvkjG6Gj0I/Y
yWgy8QlQIlpbfq/t4bwdU73W04ffN7Z1IRgOT3m/XOfZOK+GzJp+/g1xHwWA
/qI9ZDn3Ka3CR2Z4kusO6rgJvKs7Gn3cCwv28Fg0x4xxri4gwIKYHJZpXe3x
Z7cJa/scIQgS3g5wWmXdDgtdWg3t821s1xT7ZzEymob7fDOymzIQ7gXzZU4v
pjK6re4YBW6dBmiSeBIQSQgqGXJBZnVXa+0fS9sA7UmiqmhRi7Ed7F49zogI
xjJWT18szIju1RKvwhUnAThnrE1GIwauQqw4HkEn6lMgmyWTKRH30Gw/QKGt
7MwLUAqWW5d5pBxPHKMWC48a+CppnW2HVC5mGgoV/EmztezEWbGtHw82MaRv
PJwU+XS2SAJG7BIaDXarkV3CArY1uXne894r1QylGW5kOBSlB4CjZS6G+r8t
EbsZAqYOOXhB4HowYVWVjEAJIAdngPZVoCcjQzKWgdXorM5bYHX0wjDVbues
cw95j3J6xnGNIVp+0aED2ECw8vWMgnGI1Obum4lLl3J9Isj/AdMpvutY9pDa
efzhjAn0DwxTvIuN9kFf1/QC/wCeWL0ASrFEyfHe7MGpKelB4v5Z0QK09UAx
CwEglG85LnOb70pk7EouiaOghSgw7cIQIDmAO9AYOYveZrYT8hpyXbCEMLGz
13xkkCJ2iwyDQnNgS8Rh08Xu5JD+yXdJh6L+mwhKT0jaPcrC7qdeAX/nAOKR
p46raNfbbNnlgcC0E/43aFWb6Wv+yXgG5aDGlzNLiQVyqRsQ5YjJtuE2lGlO
Qa/Uz1i6H/CXwjGVAJxl5acXSixCkPH4Q7iHPfKOc1k5UB7Tk0cnVVC0f2up
vZ4v2cX0TkU1DvlrRChpkrqv5WjuzImBbobWo08RZryCUL48Zd6+996BaJav
k1o0J6i3U/Y6RCEXrihrKjmsTXgNu19q/1hTrzCqxbHcKMnJYiI6NCwYz7J9
wUF+krSjbJEOZzqWz3P2My3tL/OfasBhct4kadG59r0SIx9YYsovzu3ODKrh
/KCq4nCdxF2Yv6Bbkm3GLMDkumgPFUMIAEZ3zL0HknbNcd5CRaKs+v6Q2zIV
kK7KFxk8rYP9ibU3GZf//2yMs5WJMPnEQDHVAXpxMS9uHqnZp1txUJrnncsk
RHfrHMhRl/L4qODkZF02lDC8kb3Cux3kzzC/Nh7+M4rKkQC897HZK5bnWBQU
npnZyka0EHCJgOnH67TZwXV015lbtxqAA1JDnrgOoSH649iInTJr1EoMvIVA
dFZO2QixYn2Vd0fcYIJ4YUA9ScHxXOH1xROC0PEHPMGQf5D2PNv7cQTDw+Bv
lMmsoa2au20EEXb+GZHLUo1GFKhDW89GsVq48mmEPRaBSKwhHebeccK04ogU
xkta3cEA0noGNrpbTdCqff480SbX9hl+TIOKJAOjT7pfPdywfnR9c+JCg2nk
1bZZJ8zcAsL0iDKuOrx+lDbnGMcuyfvKMtEqQ3937slbaZWA0bR9P1QrSsJw
KD3y04Nqu1gG31UV5VGv+LPJ7uq2KoO1wzmU+bObumQU/ZrYs41lIRYb8r4C
9V2tBrNXFpeeeIxAnzushbtjdLrO8YezDKltXR+CtlOMUpDUETFfx24WcBZ7
ABHt5oCx2zbCYga3kph9mHpF11yXTmo66seU0BCcfPbcXbgQdXihINDgmvFZ
th0iWj1WPNGNSzpBJ9W+QkX4PiYUUaLqI7InROKv6l4J2ITOG/u/hrHz2mwe
1ZqSAEgunxeFSyKY5HNRKh9Cr79KkO0oeK0bFyK4iuipjeVjWNTDLxmOlADM
ajBKfzQ6Uiouy/ELuDEc3+4FYgLMtDJudmaGXosv/opc1MpGa4+h6rNFLpvQ
5DPAjWQjpZoakBNnJlDCMQnfAhY4NIWhZ0ce6ekyPXmbEaHbLVxKfGq+dGHf
fSymtk6tHUSXvdoOcngnONXfSg8pDo/x9u8PXllu1PzbNdeayvI4lytFLq0D
vMwJSeCrkStwJku6viM3iukjwlt5JvM8DZFDJHLSnOncy96Zl2n6CjZhOcp9
17WHyHTlgkrv3+6z9MEKkHcyMNqmzWGOw4aK9gHqlWv5K6nlpTXHNeM8hXHx
PkOz2rdzjFcj07lRBnycX9oHULsjYGN3e48nvDFuiOjvmu21yOTIL9qPqMLQ
460dejPHsGY2/hog1fChfoJRn88Y+Z59LWp2PVUrOQwt6MNawHJlfh27qLlP
89TulvaNQI421FWDvqci0Zrwxpg00EjS5I60D3sNI74UsobmWEKo+AThjabB
vlyf9Z++agKBJofOe/Tv9rec522aFsxFslhx/xLvUpHGgnRcNcsSOk000Hcd
2D4faEavxD0wpNkeWzAtPbIUlZ4l4en/l5WqTM1WpBzV3wmdWiYtzZwv5hJ+
1B5V1nKqj4n5V8kJoyCEaALxHlmo1L9O+L6wfGcwK3jxOJk/yzV7LGjpxtbr
Ap8HVyzHo2arU6l9PFvbyicQmYq9TkaRZc0Ur3CZ/ciPG5Lv7nNBQReg8UU2
pMpTabKoM/JTtE8pfZHylfBDuOgy2eHVZasgec8TZLWbznVFBoSBaiRcDgrj
YmeJsSuvWSEAoTP5LcNFvO3izwIUGhU2NNbZFFkYTzXMFdIcbWMwPEeWcMP5
pRXbPs/G1V8YHOukX5K6YXihAe6BvmjkyIZYqIhAMRgoYbcxApz0u6yy0Whr
ACDAzq9cJ26yWQU6V/2bc90L0nnXtl/nVSeSGCHapLMoQy/6pe+4UpA3NacY
qeI+Hvl7PK5vQlEiUOCLSUkduNiDDrDNuKW3TEXIEQ/GgdXMjnZc2vH48/Kf
CmeuQF4AnHhox/IbAAPEZBVkyirpsinoZs9AcTptnX+FHYfUk7G9oLITiGgv
90fxI+uqr5K8nMQGycIctGErCb1Lvm4qD4daJZqKtUDrH9Ti+r7nTU0gFMM3
Nus7pfnjaqPuFNOYtAQI/pgSRq3RmAufi0YI6EhAmLlfHE53GFeJkuy7LIiu
jvaFP04IImUz6t0/9HDNfcZjMVTnZEb8JP8EmKaBNEoY3fCjouoKHXjCnmGJ
c9AQ0xg5k8ZEA7dZdToPr0ze1rJdAm6Aez15eqMT4dcZz9lC8B6l/kB5qnv2
bPsI+PfjoorvOy1PpC0BIFaIIKSisGp5HhvTaEGP1VBvDye8eB8px1UpDTSJ
+fiw0s0KGZuNLtE5GauYggwAHOTU7Se1t6BY3/GquQweINXebsg7K2OPSHP2
4zPRArwcD4SpxWN08eRuZd5TSrEDKC60lyUPInxf800ZFO2cHztro28gDK6a
eIvse96sL+WTOBKZDAWZgpnJBiBNo+Y1NBLdyiAfob5UazybIWRCl8tcyNo9
SkZtryoLKwWNp9oacxkj3LFta2S7axBnH/+GaqIrNcj7xeEB9OS+i/FQsQl8
dcLcUGEK1rCysLaNVr4bRp6ptGuLQuOUqH4K6N7Cn4mSEfNXq/TmNHMHHtnT
2XNW21Z2VFkfMdOXEcw8qIyNE3leVGjlU21BG3LwaaKntCv2/K6ae3dMyLZS
qXajF0JktEoVrpBBsHd12CMUVxLIGRRVu/W/xFzlJpD0eI18BxJynC2k5gQZ
iYqugJqyeOPbNFeXgotW2sO03hE6M0nexy3V//wySLXemYOIolZKxKXhcnVY
KCt8S9qkynI5VbBkXGCjX0RlvtE5EVYLlKqQiiSdDd9298NEXuK8waV2VZ8U
l+XP2ZPQBRNVB7O4yZjC8YjuVHoYj7JxsP4O6llmG6g7sSFPCJlO5FlrGXs4
OWzYAjk3SyzYT86azStxHKUwyNHGXJs7IRX+IqmSaJJmYDw7kvhUbZSQ0AEa
aBmlMSWHSk4l/8WANvoeU1pxXl4sM895enu7sku0NsIC/4EtCTEC6yfP7vYy
EMkiERarkZTF9d8WaCnx1ve+0dAyXJnMuwCKDCl9fOzN+8kWsYd02aqB2gBN
zz1CEzRI7KAbEaWoW21NIHpg8w5dO6pT/3sy/OgakjNN0uXEAVDF7VAX6r1o
jWc1aqVd/xoRxqHtmzd8C9wsp/wNnXYZOk7jei4XqdPOYbIZmOQJtVBK4cl+
byDZAyv+Yo/1nKdvOH46n8/sMlgXOy8C8tkqgiy+YbJffCXM13TVryO/XuCw
OdeyM8F3kb4WG8FMMF0usYvwT+fwJIA5uAWLM7eDe3x+KW4gVX9WyGbab3/I
f3yi+OsN/XTj7xe8ojDDOs/+8ctAAvbnHSxPaclC37gvnF3IdtiFXXemHzMd
4DYUzO7d8w+Uwh8iMf/VFJ6HbHL8QeIhz4jrIFf9BOwJkojPcV/tzLgttpl5
vjejeigV8vpFniENa/ToH831BgdqUSeNqN1/uAASNmdxViqbTjVDBFh9+FqW
9M/C7mS3iqDyhVg71diXHfYuRt1Vw0/Dzrq2S2X4j4SaFJprmHDc5nbElIZ3
2FEKN52WSLpq7Gqy9B5B2S55lsIh8Xp8tjDer/fwPJyVv4W+uAdVMlOabgfo
cm8JBwdRGQFoHuYjZnqUVQecX8nMW3s8HJqAhDRpSuVte66fISxJ7UTWiUV4
BZ8JzjrSlnDL68Yt3lM7ylsmTqpBN96+ZfQ5SBIHcWxakRq9DkcKX8E2UDYM
ycGdFRk6zUa0leuaCkp6lyswvbEn5h/RNrHIUwYCvKIlyJKAfJr0+z6e32of
qqVk4/P1EW5m06awWdM3juhyW4bM+9biKgg10bHqzMWG3QMWS87/KyS6smlq
PEZqpYQ2N1P/f4y0CX0wiQFVWeBREjSRMojCnor5o/5hRfejuExA4Gd3L6j4
b4GeRON8HGe+MkmBGjFmruaJxhcE7TqlLlhpckiNw7bPbVjltcI50MDtadR2
VhQ3AtZo+TsrsH3OZGbtU8AQySyxja77WiZbBBg5yA7/vUMtswLoZXW6gv5+
e4W9Z97xQdHw6Yj06r+CTxcbEpNaYlkuMEcL6BhzZoyrZFuRX8OpGPd9eF9o
Eevmqt9jo8SK4EjcKSOy5mZKLmWT8NWR9dtC+Or1+glqLgibbL074yD6Q3BL
Lvy/0RVm6Zne1cH9yTwmz2Iu2DGN+Jrv7DIFQeD+2+p/p38UnW0RomtSj79i
i2+mX8u7OePvWxDcOpNAX/XsVS+MEMW7+8jlI1+jbqSCmXqbhzlg/oeoIpvi
56JI9bfVUhRFzoaDeqT/4OcEM3Vp9Ej3udgpp9JTChWCiNxG/+wapM2r+fnB
S2UNyxb98rpcVqzkZLcHHq3PO++TI4bzdu+IS0oeHrsKng4pbZ1QEgnf6b1d
5LBDhlaWu8ifsuKeIriBctb5AMpJee2X7c6p0Uvu24teAtnkhZRZOIFWxBfw
wddJTzQiwunEarrsQ1JW/hVhO3HWBGmOj27apmg5Joa48KlqDdRUguKv0uwf
9D5EdQpdapJd8RN5Ff0KsnrZkZggoQni0bQySWwSwZptPLHQHP/74n0cYV0q
tWxew33ahBJE0laFvGkwJ+otwnBY2jF07pCKG12LvVZ+qlFLPRUMwP/DaTWX
Jp0GNTfksZUtyobHeehmdQL4wwsMrlP5fI+TGYEoWGC+WWbluElhALv+Bo8o
wnXIUkVHwq6qvvlQap7yRtyT0q/L6ggZn82Gxvb1ZDydY2zT0GgnompgP7V8
fpLtnA7ROnUE7ke8RWtRP3+EotbukEjom4vJAk+i8QIXhNRlq/FTuSJ8984Y
cs8OzFX+nc3rCmkasa2B57sc5EtIuS81fLcHszKPdsnCgUTzUtQaW4AtCzTt
vNYbVdX2EVI2Ie7QKnIpQJ6FVAWzH6wg67BFyisiMPbH98wiqsrxk2zeHnAf
ZxLx6fqguSrRjitLuovhh5AkM88TpODaswqhhJgB+54Se7mn5YHlLFwCQd/+
YBqnWMVt2VNKgvAB4sPHROumlBSbFyO3LVQO+nEgND/2w0KxnV6IgX3MR/8W
hAERmqZzMH0JxChvWSD1q+472KfkkgpI6aF3J3FrbpEK3HogJjCb5tSF/9C3
t4QPaCP4g6mLmP+b4hUmxh8H2H8aM8BOnF3WLjzmhT9qou1IvzehfHYXPJXz
FOQbKoBAuOoiSPupqiJdbdTyvEcyFrcrr16z9wFu4+L96i5c4dinTngVYOCc
a2P3qOJASl0A3kJ3JsSVDv3/pSKk6jBnhRvU8ur7G8+v5IaHcy9ikBmRm+oR
TobCS0XXhkaQWNa+OdV4FqUTvCKN8VQwTtR08X38ytNJjw1KdhVp6OhrlWh+
JRLXEHy5MYZi0TmCG1Fyo55f+fFuBL7VPg0je6CtoGs6MaRu6JW22X/tsgu5
m+q1KEGVPOHxUrC1Lt43b0fHMuwPQMbLxM0ihaTx7ukMdkh4tGhjArGboFB3
dmlirMwO+xwPPHdMv6GMHY/NjVsbIK6I/u0Wu6cbWKia4NSJOJeJqq7nwdYi
OzjetXTZEbLST0Dbkq8j3qox9cKJnEZH8ntKk8E/5e8sU38x1II2PE7jRRzy
Cpi2sI73UED/W5v9h372G04qCueEZ0S/heHpR37cJMzX6yCnXPz/aX6/3zUc
Imkd8+2lVxmv6u/xMdHU1y5mBx/+PfI40iwgODBVChQhb0yDt30jNk5oEPW0
zaSllJ/bJBTUfYDHuglgqmmFxBBmMG8cYPmdaSiCLsIeLS2cMwaqxTNKlzyu
ZeSFUc4JunrXtGk5RVtAYhJZaAiW6bHLCigsIIIGqz8Az2wfyGR+Gje+OOsG
ddIn4Yvu5+D9an708dz8Z24x+O9C0L8LCajB9rB/HgH0ZBVOa1uAHlOHeBVm
jA625ik3F9cD6JGNY+hwS3fdfgNi12HfpRZK4QHM3eFnWl67CUaATdnCPxjm
k3prrOmDYhEm483qcSBfCjaRxfu+rLjkDYZRzbrBvjWvtMqWGGLWqorewYAv
ms+5YbYTW8zCbK3RLnYXL6C8xjsV7qv63w6YIyyery7ASL+L3kprVuUuTlBy
n3jB67oUWkMesZFG+nGCseqDovMRp2Tv6CahNluitTFIyPMk9JZbzTaO4bQy
Z9Lb6UlJakvQ2a0L7iG05NknLmihQamSL+vJgcDixPGUlo/w0P6TknogUOQR
gNknQ6m1MaCMFlqxEN37nE4xa5G9+yRCx3s5eafLL99rR/lwVBVoc7sjAbHP
eI/qsnbRGlUET0lZPA9o9oWOW1PA04X4ALvGzyS0oYdUAvzEd+aj8+54q8GW
7IrIDw7p4UZBedS2fJlOA2ZXt9LHF1evj05chozsqAG4G2D5AcIKEpvZyswb
UDkiCkR4Q21Zgl4HgCT3jME5n7mjXmTAzFb2gWTKd+SeqrZQktkpRslNXwke
Nq6RY+gKAgTKRuDj2D0DdbkGBhBpzwu5bIoR8M9M7igV2+m3MSyVQK92vhaD
9QYYPdjCMQiMlcwgTxtjHDAwQoXTIFJr/8/ZSMynK/HcC0mzYXTLIUSmMAhE
ofayftj6VNfYiuqkdLC7t0dunRDDx4T4dgQNYfvwx2uZM9p6mfwY0R9AQbEg
IL92JaH8wo65ahzP5dQTJrj80CQgnnqQyNPTywvFntjWQFHMZXIEa4Z9bXuf
vZM+fhBPcCOugzrRvCM3xFlYQqaa9OxEH8J+ss2VwGc8cRpntTYUdKdh6chN
Z+BsGln4kFVMi/AoyZpSFCANEM+x54gLzxqW5DUEX/mU75jGWkIM5rF4ZsvH
aXeCxKPT6xl6zow/FGnh/kvaFfuM56NTKepMPCijoDLTj2D5Bq+yVz5yYxZt
g/dbIqG18LX+l8QFKq57x+NpLl1yG2Iu1oFmkwdGzkd5407yqa73gUhnPbHa
ED19Uj+oM5aCJHCgXgAjv4NL3NgFRZTsRVyPDZyLWRoEydNLFSoJu/tkS4+j
7iYXG+VIdK6dqCqnITdEOFaLqKj2ag30AKXpbQQ8SIT9+yHHPinH0Xdz4fw1
+C6P7Uk5QLQPcADCN2BxgKlCuCfOgKADBPK31IX1hGrYIK5k6F8+X/ztr9l6
Etov2OrWFwG673K8rZa+bqQYk+h+AUUPXKzxHYTwa636wxthUG3giwpQXN1a
raKmyeNYZSpqBPJPlILySq7n6x3gwT0yzBGb0gdnTTFvsxmGaVkDv1cZkNBY
HGryl9in+8Ru7ar5qwQxV8B0Korl0i4Mv3+aL0/+EHrAv/pLW7ze3BX18nR1
81/EDSp4SVn2XZ8D8xt+aaCVdJwNV1JVnn7/A7vr0XGa61nx05sMcRDSb2FM
f3ZFLMFKeN6UYyEHy8uBwV1KmmVxtUdClBDCLVZdQgT7SMyU3pYHnng6+Kv5
UJWl+MgOJ5hAYLos2yFKomLOP0CJDaM/UuyuEXRxWYymaVyeDKt9pJD3E60d
44qok37lgMw9P2p+zZwf6mnnP0PfgwaS0D5QLXAMhu/cJ9/XgYF8zpxqnlCT
WCZvmbKhGf7H2cBOiHw9Bej4AtXuSGQtHYQY0iYIhqc/+gkRZCBfR1ud9ofx
uE5JUnRkzPBKjsCRtJXNWlYeARepRoJxz2nJ2BNja42+n4wy1QZRz3CA7Tzq
59iWf7Ym1ks+gBPqg1fCYOeDjzyaOoI8bGvAJTjeCBCT8tnMQbmLsl4iCWsv
zmB15s9dQxXZHd2fRdHEVK/pvgHFRJs4ZE08lmGHdy79QYlk9KUGpAcL6/2C
5KIJK3SFvXFaBif5tY+bmfDJDYM2QsDjRJd/wqHGCSIkMeNomLY+BPExBviq
1A6EnqPY0h/jSaSZXZE9QdXI4VLw0wN79Agf9rST5Fi9jshls38pSBbAXasr
w9ML5WBSQgc9Ine8TYI+CaA5J3Itt9UnZHQdpyo3h9lrHRZVT1RUVhOYJKaM
sLtJSKCqPKk20Hq3bNkJ1oXM0QukmGdf5ktFiLQR9o8x1gi/q3kmjrkXcWq9
wArafUDXBKwrRJiADcaZayYmRZvsTku+w8D58Iax1ymDqzqkDUbt3z+/UfyI
Qo0WZjDR82wJmRf+xNub5olTz7Ucz3+78qJW0nxr/Odn52PXpuN9DsZaU13d
WBDzCATLhmSPPvbQWLyfqWZUV99S19zM94WPqmm3X7pNhgBA/gZySO2p1FEb
e+03nvQQ8wxKH5k4NKGWTzFnNqev82LEEQkO4De5FRf1vt8RJqfcZ0Wo/HDB
ap1n0VkqNU9S9PoTAL8dAZW//k9o7Ws1MKWq1dalKC7sPOAUt7m6Ujd7ZrCY
ctXZmFwKCiryB/CiuIExylVAy0sWAjRZRI+MPc9sSbzhsutbYbPJ+zn5N1yU
Y2+2ZGQKtx7aQX5flFGcfvQZ56EDwFtjPY8ozDHeXe8NjNGGtZ7x/urAlPC7
4AFro+i05VH6H07JvyPfh+LeNN+6+bkOQx4Mwa0CoZP2yi/7MU9a/CpGMV9e
8Wupyczl9DVE06PHFh6GZJq/3WzVNkvsMuelIqEIcKMux5x1QyfD0GpBFF56
XQM4f5aCuTgXytb7m9N/saFjEOOensIRQ0c9pXwxc8SlSXqoQ+u2A8eYybtb
hVmPkY1EiAwQajKIFvS4Oks+m6/48WAWrZL5efL5EtWkuvWnlVjKUSRFcbS5
NBCUgD8kXpHnqvT9PX/UX0LalBFWBUGp3BNTst6lwnmIncf9r1ZbVLNo/gum
ncdDh751QTlHZBFPTPjWT0RtcdOP/Vh1LdRzyKAQhx7e2jYJobk6di1ctpF7
6jNfoR9PtvpANpwSBftXyty0tXSVv9y7z2bRFwCyXTphVXQPYNROUmVDCz56
ioYU3DVnQng2/6TMpsbr3Satl2Z8OIkL7RyXP3/BFPL1B/66IGILU2AB+Cy9
rbZ65ENFYxIVsZDr3luKe6pTDZfjNHrJcpedzICOg+IPCwuyvXfQ4P3H6SdW
WP5dfWo8RL6Pb9GKotgt0kFZgAtf6e9Z+MsOcu6zj6V0KdvVtMBquVrGUf6j
H/bdVl4qlYUMJpWZ+///diaID9Erwv24ZLPAJbJs4jLb/re6MuJ78/ujbYfm
s0Tqrdw6T5ndZ081RMOvyXw3MLjnxnzhUF24xe7J/3kXoHpsi7EXto2o4+CT
2WturIr1h/npdfVd5r+YEYul2GLWexlQFE9c2g9bHMdi20TbeGjqg9KjVBy/
kWMpoBjus33oueuU4Jp1QySKMZYBYO8QcXVu0R/9goncUcwcjf3vqMI7ij+v
jsyJBdYxJrxTy66jTBKHxxdAAjplstJcYZUqKyNOnJWuvf0iXAfQrp1Qiz49
aGh2UmeWVZ/o1QrUR36wDWwhHCurTJB2tn8quXJAzaD3KBNT/POk+/2Muluo
kwb4jXhRKeBP++BAmex6A86HDAG38vG6cY1z2EOcK4fRuQBJFZq6mf+liZNo
4Gb0O423c7B0AeRyiBHA9yl/XBU1TQU2qSvZKU8Nb5aSmuDFm2iy3DXlo6ze
fdGzpWWsxmW0i5i0HTfacFJe8JqdtKNuyfvKxLz1p/1YMediACtV2iB/Af9Y
tE4caRGE/B0G7vysaRERLQJB29nOek50bpAQjKMfY6jKSg7dvFNa9nM+q5dy
26RfuDQZ9JEdT6D6y/twI4vg3XTRclQdOQ3sns23dPRbsA3aS3KTOpUGml4s
1CQQGqjpv2TFkWC2lR5GHrOGpm5zBy1qyyl8ZqYsq7QyWiwGJOA529pXFIGl
kulKFKMv3Osr5ilK/sgBUShJLhaZy+OUzz77SqaXSSq4tOH461yJZRdrdndS
Oi+08/HnhQbsSFkwgLws39QBPTre0dwidka4tctaOA/Vd6kgIYZIUWJQdXB9
9YQD8dtR4kNKMpP3t+i+m9pAdzaYa/0Z6lGjVN88MiS3XMzDZECicSvGqPsO
b6rOBhyMfBHsTdUZByD5uail+32XwjB1v0R4+4WbiDwsns7g64N4swqFe3FL
irIPmI6HqXV5aETs3ioJUSE6kY1EYTUK07ukRu8tTDM7VUjRf5YHPl7ZBHhL
2UaatiBODD+lEoE0d0doomMIAmExodF0Zb2Ulw23WdIIpfRYUMafNs3EBDFX
jYZaNO00b1icyyzs8lHgJiHQ/gtGxyqYpKeU0Jx4RPbwvB9kl7J23OhjvVCQ
iUw1iBfmBlnnuQDs0wxO2dkeXrz6TDlHeEFk7zjudvYE6xotOwjSSXjoXjiX
kHB+Uu2xiCwRnng3O05//cf+DBZMTTVUoY8a0p8jTd5QBmUDgUpsdc/qnvlQ
Bn1UsG3Nt874o6xTOSHdFjatdLZEKZNcipGc3smVCcbl+3Pvgkdmm6nAFdwh
q+WD7+Iy7iQ2MZ8A+ML7G8zRnC0wdylSzavpQu1xyPxYTOPcznN/6ZFCkP8a
lVtVxXRDz6wjrfbLHcIHHqVXfAg0MDj5ssAgeNDmAHGU7ZJY05D5CJqWFYiO
TOB45h1HRELGfduMqve7pmgmOSVg5cnhlIinzuTSP3xnjnBksYOYBWcGkLvb
npLvo7AhPTMXaGNjzlg0CH4z6EsgUVNSO781DiokRNSmkAs23EYNetr77SuK
w1p8AqYYHqZYMAIS88CShHggLT/eHQbkecmWtsMv6tSJfw5RBBATk+qZxGN+
u8xFW7XvH7tjJd24x7UsOuDm9lgE/PWH9ZdJ9CDlyqJm3T/caUJt5f2AK4+N
wG5LaPYhtOKybIVTUsCXs8XfBXlpDQ9j+BPXdgGubVaOwkr6qQnoxxNS57iS
tp4QC0fantcTesbGpUBTHTSbX+aVuqT5qxHScyUq/iVgvergDysusGV6zu6d
elYcirwdygL47m1xWi7JOtwHTxGdp+uNRkzCl++4jaS1IrGISvOC2HNOFp43
A5jk8Ry+RQuc0aCBUSqMyTbvF4ZgxkeEhIfG0fbp9G3PWgKc2nlOsihuOhix
Dhd5hvQgAycdB2+SwGzlsU/fdnsyDOdXgXWIO4bcN4GTpJ40/C45zrN0Ck6v
IKgnb4D8n0b0WLkg4tDyktLwN4BErDJ+A6ToCVh+K4fmMMErwAYjyW443Jr/
lNJ2dZzPYhxngQUmVle7sA7hWESzAhOC48RiltHtUIebDquko/m65encIuBX
pK2LS9gAcpeU0LIGUifLBjDl0fKvqmI/Zu+9sl8v52FKax93XwqXhIWvjf7D
7Le7E7mPs4eQ5hy/TBZWpScrfZ+qS0dneAZ/Zq0VhdNCw3cHIlzde6SnGma6
w3dt3NIEks923L9E+cl1EVPWr4j7aqGdfjrcxDYdH6wrGiw5FlFk8yYCSzjA
KJg/R9Hz6svNXwK8lk0Qp0kgadgbMGlIdGZI015F7VKQLCo3KwO1/QiocoaC
c5zwJXsBNEwi3kKUW1vWrapPs4Hp92itFrk8YsJ9n+J8o67eUUyCOZ7MtQTi
8YUZ/zTLZgKBeBMR0rTUweK43DIE2CaSGGld/f3eS5i1Da3hN47G3lsPM85/
6y2HlFySlquMHqiZ4xJeO7zuAonTq+/OeyLsfwUNq/32YhDDV5MF1cJh/qIy
pKwK7SVL1cJx50qCJdSiDZ6mzrjOwpJGSwoRE17GR+BC6eHEVFTWE2uqMUhO
6QeqfFTVjl1sg6BXwtuEgW1HuCAJ0UtFIhIN5GFpubi/h3KWTN6VF1PCAZXj
0O3mKFiB0s4n+qvMSATC5Ng3VdXFQL5ZpUTLTGGsOwqQFNcIsg0uzRA1At1A
r83jLt0OuE/qqWBmJLUA45Tim5uqjsdo+BJu2wEwaleZABZLwfNzwZP21MDB
tP6Yo72b8qUgmGQErNb7C+pi2UjGRa+YR/QXMVfhNprKN3B/MIIkgddon/HQ
7QM1XemO8eStoOQTDYPIpNm4GiBQ46UUpfSGF/ogtISAXx86XgRMVR1oxt5p
AsFCTLgftlSdE+eBYOLqe6HCRJMsN/RDS/RU22eRswdxKM37L1+dkarAq47X
VywR9XmoB/YEt51HTivcYPilsVqzdKF4vJnfghsaS/srn50XK5/bpHmSDX1b
xoooCNGsCWMf3KPn1R9rQnAycI3mG+MhOZNq9VH5O+SvZ/ARfBhl18UQLFIG
L0lC4xET1/c2Foy/jsiW8KFKDnWLdajl0oJSbC2THudQNzDg+zeY08svJmqQ
1fxZJjhVwtDKJGqnJaL7keBQemtSGDqZTFjqMFULLgcLMHC2UNwo0OLAy13Y
fWcWse/FL743nHMmUMSusU3LMAS7aB7JWsb86d1qqZ17633CN6isvIgOl1WY
J3EhzuhzzqXAA5rnxArvEilHgrvmkwQfqHtGo2g8LUXoG3zoww7XkjqLI3vW
OfisJVSGPClOSQulSMCWgG+V1RSpPS7RjxoH5SZVPImW1DNPEcAc2yJ9BFbb
B0aqptmkraQOeZvydX9t1+axUsj/fzYgTOhY/sQylah78YVKTAy8v4biyt3G
BBIfoHhlWdZjsqFD9cn+WwfMEypXnycEZmuRVvAjZa8ABzR0BXmlUt/AN42t
03V0DJs+PreTuil6xMiepUrmMTkCMiwGh6cp3phC04ssKxPj3s5x7VWTG8Bb
nT31U+B8B++YN4NG4ojkfteNM+O7vMSdrDA2ic32RF7PXzzIOwv9oS1DMqCJ
NrZb4+UC751Hzr1bSXS5d1O87nnu43xhNoS0OtW5m61gxXcejRwme+HsdihP
n2yRcUez60VcET6chlDwNQl3cPfSyzJlOmBqNrt8vl/arRyB894b5mfyeAtB
cd4IMj+ErlfWusSBweFu9e9KKabpvTY85IXyBrwEucqjQNtw1b4PTKuyGH+T
tIAtgpuGvokLOIuOBnV1aIipiMBaZk1n/IehtG/2JB6RKV4Z5VcTQgSV7EXU
cB3hZ6L8g1zCkfYGt9Tt3PUmtq0MxUfqQMwKxUn81+54W7gxPy/37ZKk7czn
23Ouen+ZinpAW+tatJP/VRYvlP4BDcRQqwLLSHkYBlCWwULygBtWK+yF0OYc
6USVqHFfITyBbqJedw79y8mp2hdwDbTagjbPOqrsDww9vvzvvguOczl4z45o
nIXI8D9DRIiEfRMeVZeAYNQufYv1p3xQ7wg1sDSZudJnr3YjlmbSDw6UCHSb
JZyxMmL3XYZWEAmeFLk8CPhHGFSNWClqEp5YEBlogdG0jiXBeyRukx/L3v58
0SO2GMuPmEbHuXsX7WtF4owIQLiPDBQLq6/Utf2HPe4XLm45xk01vuPDXMVk
4nXybMh+txk1gaBBlXhNV3xNZ+XKngoYSDD8VSwVrqoVOq8ZpRvtUMW13kHF
0RHqVDJHdxXLRM131T71MOOboJsSSlGKRzInd3D52XQYpC+xMM7dKGa12/Xx
kJtJ4hrlnhSiGnG8nZYNo5pQ5buecq766olWecj/C41UeU2D1E+V7k5GPYpa
xnWFeWxd4U8Jo/8tK7LoSmnmJh551BWa6nxcg8sJyFK+OrMqVs0HGW9AdMw1
EptasLUPUuhXXudNumDl3JS2JPW9LoMBfs9PeuP/ojnt0wKUnh4EjuVmoxUC
6t9liFZxY1driwWKaAZxvEILpWaNFlXwXEmWGUjc7kP2Obi28hJdpEdatCqs
fkfefbQHrCj3Iw0L5YvXI0KKKvD7GTAvWsgPBJvhERZ6jH5X+xtf/qzX3acX
LqiaCSpGMIIMjnCmH9VcD3ZeFHW5Qtaa5e1CuL7/13dbrEOKerlcnyHZRYk9
VmG/VyNWFfAJVs72Q4Qn7pfurX2+nVXvU+j52HQ9yvZZVev5C0dT2+SzMHi1
3zmLqG9WIxPcVMoK3QJ5N+0XSVufwbtyVzvtuZtmH1ObTEAx7TtNhTuSG11y
eiEbhEJGCzpGfYglsvy5Hg2vlDhLtHneJN8OenYu3MK0OPPA9zMVwljHNzu9
zL97d2gJSkZluYrllPYHJWttnBnh/b1mYtCI7rcxxQC41t2Am9YQH7olruTu
rHAi3BKLMAWfpSalcUpagJOxXDTiUVRhI31ten5h588c3mKVXoCraKYiI6d/
L428xIAJs3nMkM/n0p1vK9zsuOljuWZj1BBZU8Oxj0tx1X1qTuYtkmiL7+O3
K4Ht0FAYGxPcdJSwN3y77QxfJ7YZFiwxd+HkpJcvm5ccO8RaCsPh0PMnXTun
tT24RqDeFeavTLoF0ivz1ZAKtyK0cWYS5mFXT/G5qHXPuyJiz1MTwT7C/qFH
/EKuWGhffOBhnnLYdoyHFGZHzndiyFQLX4UqyymDSQlts/Cz4WaJiI5Qk8X9
EHMtJ93OsJtbccZmfkjqk3ZJDBKU/WLas44FNFdu6LcujGl+WFVdxQ3zP7nQ
Paiqjv413zPFmK0ru+ao+YekLU+oIY1xol+reDsEwFeu9ivdBkA97YZqw6bt
xnWx+jQ0p1SMlEpl1npsti7i2XwLnaUzwVKd6hDfTDFIEM0O+8voYYY4OK3M
7KkH/nzpu+NveIyh/O8bkALDXIVb5TtKILPvCK/iv8kEBXLJjAfsB8EeBqX2
Ib2qEml1l75FfV5as88lzOWBzougvqMs9KgFFU7WUgRQa3KOKJyUBQSG+mcZ
LAdcM/2bzme8twNg/TyUSpkliw36P5EhTn/d9Xp5jIyC7F1+dDwcqYLj2OSO
WOB8vK7FVYfbuL5G5E0Bd83X7KdpoLX+OHBNlCcutCq3B9AhoMHnHkTgF/CR
zH2tDLSkmmege6UmvxWkOXv/KUbE38n4Fhn+VMpylzPsbW8YAS52Vj/9648l
QkG1Ux22M931vFlV2pvFL3MrlB0KFQkvGeH6yTLG3r6a2Zk8wBO+ohOLafU4
NQ+bUj11J5oF4XEaA5RpzBaRnTPqiUn5oEEeJcUoEAtcmSFRdecoblcc9uOP
DHg7bZCmulrHhp1zQ2fJxV8jAI0HFaObEL5yvnym23Ldj9AJE5CCFabRhyPV
J+XjqkNGio+Nx1OjmFvt3wh3iyjteCxhyacNAtVc1RH3e63CTa4GVareueVl
ej1v/u7VPxh2QNR8XeSXP5pYoA4+5tRKIzYBUj1fPJYVSnWNUbSYRMGQoDfn
rIAOypz148Gvq+8Ce05MAMQG8ak0fL3oKKypQnHf57Bq4d8z+hu7aCYQKc2+
9KOySG0i7lfbufEzFMMLmpJGrjjFztl6SEyVn464fTBqeSmoVVTJ6rBjCYBj
uMEron1VIbu6X+/nP7BOGb5jFWFn/e4tsYJ1KgOBtyXniBzj0YleswZtVSna
MuEyTGGq/OD390O0NHQgd9SCBMZgzBw3qXOSSpwAcvaeNiX0bPbsPumE1rVS
2Lccc9CTKMrmn/2woYUMgNvQ/9Kti8r0OVhks5mY7KrikfENhIv/sx0qG18O
q7emXOIaqaSYGz5UbgAiMGm0NEisRoQxmcVjbkQyo3P1GouFFyNm2lrj1Dxm
n8mSf9KhMBXqO70FbJ6eCZHVn8GtSEFHbGinAjRAJCYlMTCqRDi4DxezDpJV
cLzM1BDDbeNicjn5u/fMWLXSc4cowu8amLkojATKtzjzFBwXs3XirZLZsjM1
jtfroH4daVRl6zcW7KP2CVNnudwBEGFZhiehL0MrQ8DbGwEmowMhV6Ftjgls
3QFShLtl3rJR98MokRiYnbjVLDDN5UC6eeKnGkMEA4qs6n4FL2CpTzDXZFlJ
maEGmQfnARNdRzWrfMeHYXHr8BHDDzl9xpqBcS1hQnKn5ufvpGQ2juD5VxlC
VVUnDV16dD+nkjRqyjGHhlKTpvKUFjY2VYX5tUtle4VWdziv+V4tkm92GBdB
WaOu3NVqdcPoDVM500tYtik5nT4CRVJMXPsuP8rvrb8zzgaAuPUargUwTkR3
E9w+LFYEzmXFK7bpVmw/rHCM3UzP4C+GSJWA6XRuqmI61AfTYIqLQe5qfGbe
3K+M7c/1B+vCLORzpxehkcR4GJIesW1hst1QdqhADmrYkFuQVfWNn98+jqVC
rZUJcOwV05Hioa9yuCAQqaSNRhmO/U7N2haTc9tGBaos8bCE++R7w2HCFlBn
T77jZj127E5R0sqyJoGZe8Ih/FTyBdw/DYMQqEOYDNH6+JGnZIsMxV5UatiM
FPaP0ynAc19qlNqTZAVi6G1g9A8Tp89BHXYruW+NMPG0TuIMYhLT1x/SvNkU
CVhQt/G/koHcJGIh+iI207AeVCxdDDkTjaMI7ul0llxFEi0tqlMlbVE0Z9Zn
Ia4esclXjpPPyisU6Geong3a2dv99eRJ1wG7gjZWxF0tywpTDyqiRNyb6+hp
qBAQIw117iJ/n2myMDFU5peKkyjpq0/Yiv/wBrJpv71Uc2lOZzaZa4x5j0zb
psTDb1aArkUcHgL7w70wbDWgLheB5TkQJIxcFLW4yHLa7zNmhikEheqKpuGo
AR3DA8onIkK9f+yaz9pwK6RRRVSKxlGl13OgOlr3gZsfUuQUBmBxi2GjNszg
gYMug+t5juoR7Ue1IbRRtEYpfgqSYrnZISlrnNAnD6u8eiH57OrlJIGzQQy0
VN0prRgZciju5GtAKENgiRcGYn6YJcSHPGm0aeLbUq+TGlhP3n6/xxmPA3DH
awtaR4mUTHBg1hybGR3qcs8LN8LS50zaXYlBAvVhGV5Auj7yG4QiPF9JxWWW
Mb1LC6FnYMuzLGI8XOlTY48KhjS5vcNT7nP7uSKpul6pwUnp5fPggfYdIYSK
y5sdBCfYDzc38PKar6VfBmK3FSGXmFxZI1ePRUPB7hxzSp5Hp1M67UlaxZyV
ZuodZKu2oL+av3qgRYz49171SMzW+a4saOCuSQP6B2hZf+ZorG6wmNNUCacD
bNZgbKOIlqsYM4QSJZAwgMANRcJ8cem+P0ALRGvnwmSPoSvJMhYbbhN5tUCD
tz9ju/fv8TbwNqKroRcvmvejcc0M1BIOYa6bdOLB94VmzFu4WAPzPBGNh0s4
MitoWjXS5mgHoxpQ76dgYzFIabgFFSTIC70+nwMSPVvJ+y81LZrQ6g/aCaxU
JEiGAYDf7McCAEmlu0FLJEp4znGithvKDu5F+qhk1Bgk1i5j5GgJJEJCGZ/1
5GpORbhwBz2keDXZmsxfTrBGZExcAH9hlooRKT7BOetg03Qff2jbmX2gV8Zj
6t1glDXETFwFaDXxDGxloqJBamTjzCYBSfqjtJSgh4Om1MYxytWM3Kt1dbEu
aOg0Cj19NzmpXE8O4YlYjliPVSPfbsN9UGnY3HG1s5/PxmffNvr6xT/4Me1U
qe2E7dfIQs6rhNldmKJ1ucWi8+pRryvLGkgiU8/8Edp37ck+Uafi3Fl3bcGQ
muyhxXOLTyw4dbBCBiZ3nlV0yMGcvSqOfeS59kWZwsWH0Y0hTXyjY49Ldymw
LtfmTAUgUg9L1YyTUVtOF4NQ5JN0AzsOqMB/Oga9XBLL000MuSS+dLAUwBNm
fZLaUXYH3pZEAgZlFmmsmWH+w4Y8fzajFRwBHV3DcAldwl1VcnFImH7HzCUB
aBKl8eslStMLP0hWWcDxI5qkx0OtP+A54oAV3U934jHdloUGsxr+Om3jvCEr
qR+8GAqXX9qiUP4Xo/FDS5mpSUkEPzqfIYaJcbRaVrGy3lfPrhYe7VGjs4kW
6qGP5oGm2+Fe1WAdbqxOQpNLb+/iE6mPuW9hJjhGCArLd9vbr5Tzwf0bmTsp
mFHFrKzcohZWXWLHUxRExmrXCKYQ2VbfkKidZZtS2fti/MEU/WnTZfApv5Es
L5OnyXrlaoVdAE6QdM9GpOE3q6/+RFzwRk9VW7i7m96Zf52wM4TA0HTGvih8
lejkrxd0SBrrpZjrCBdLd+WmQlgbRYAyuD/knAG2CiVhtiw2uJaI9rK+SLPU
iM5h+ioSvtW3uNHEVsOpVqz8e/TYHRK+02/YPuPtc+EEt6UXQPdVgtZnRwef
OjL4QyolG2TlYvmVrzwApDPaf1KUI1Rkk4T4LfStW97hRhUJeBdeGlNw4NbW
Wyz3dct2iZPxLA9BLWtZIxtU1p1BH1UMZG+r/mlKwjjaPPvSotcS4S08SM/w
dqGmtK6sDPrdxAoyPhfgl8dppjM9cP7GovbtqO6z26iIIYYYe392EgfGhkoz
k1yoB6IWaGV8pG/644uM+giR74hvVoOV2sUzEQeZGALUBZ+UWTYkMXOmzNYZ
Jz3A///5IP+BJcYiYx8kEHn9+m4BVJbp7/m95UnELRqvWDBqZJ7/KIbuj686
sm7tiBWkwdx+nMl2aAsLv5NtiGWl3swpFun/BxPDxzKpDdOe1EqQJHyjauDb
r1unI3VOzxjD0X3jIFHLVYITdUvfwg7dWKyp8AMh4sL2VeIKUMnTNx1s7qyd
OSkZQe785ba2N2BdfY5VkMHVshYDc3DWdauhxsbUsEejCIHrB2VJGN8QHJbJ
WYRkTF/QCFhqm+KLvBy4UQp/oZRd3NFMTTtVRhtGzzN7WmshchliTNDfuVpK
dokCr8MsJL/0/gZnhQb2SJ95+RsIEH2JFf9frp7sH+4r79nfYwFB3Zk9b0Dd
/1YjgfEEQwVqTcLS5x1VPU8PRuZSWS1LLc41MIa4/7qRCbdHaeD102Ut6mJh
nnU0DB2dQJSmVUoF6KTXrFqOA7iOIObcnjsL149VLMs7F98JYAzmHWcEg5CZ
M3uYO+aasZLJca3eaJBnNXPotCiwQoSb7l9ZZ/0/KSrjX4/GGDHUgj8QYUkG
5Yas/F41hdWfXa+oo3pl8DymyKxxlTiajCievXVVxfYJ3Wf9aFHx2oGi/QYf
TT4P3X1sAHPNPz/fT/rJBo/ubykUC21IUCHdBeYT1HJ0oZqfrz54/EFLV1wp
Ef8FdWOl2vPIC2QPz1KCqUcDffTs2GPl4GZ47WPosFLrmf0zrO9VcmKqjKz4
LeKDptRbsypKDlqqoNXw/SlDCq2QeP3xhGYV1qEwXGsUk4GtNnRV747eJwAu
JnOsiv7IjwBo0osKQfZ45ExuGMUxYU1FMa5iq8mMfoVax9msULFusPuU034z
kVfv5J+CM5xUtvZfRustqd0RHwMBn46iE4ZNvTeF5Jz7ithwZ/h0CbLiUBmq
kTGbq7AbV0TzHm+j022dvW/P4DpNoLSRE5ScIoyReauU/PRdLj0LIqIBGKAP
5aTWFwEaNpuzaR280TpgVvY2fHMYseYzZbvRhJb+JA+GgH1813KYRtSpPhBK
CCoXEO7vMlU0YdpiMfwgKPEpkBO+uHNHm4plkcyAStfmL0d4eiZYcj5+KZQS
ij/XRzQlceRuj6oEUU29PlFxHXDvLj14bkXim/sMQja3ZTtZKDJqDtF6zG+8
RPgHnMNqp8crPUs6pCPlzMcJElUxI2L7OFa9pxgDvZKUsVDe9tyXYU1bC4yC
jrAe10MZ8CnYIlaUOND85uPm6lpNbIOHouvPyWQp7qm6E7LdzJGZQdMSEVb7
KMmQ13IJ3rS3d7VqKpFHGcMWGn+onCh9Rl781lZZT6smAljd100VcOqJVIAa
hNxOmx8FLV7i8rNt/PhkKsuUdsRJDmxzZ7wSlgwivTpdpIcZImjSCV8j/4xW
XHOH1efYuUYdIWtvrju/O9M0cQ/tRQtZVuhxbEipkQyrING/rbT8BU3tJj4w
GxIoC+mA1Bl4wNo9mdBqcJ9ZDmqU3DJTqQzm6VEwEPfVs+V+PuTkM0mqWbUW
EvJpGjZbSQbKr1EePi0rHsiGhrZgCpqeeZD0ZfTqcHo8/bl3MrPQgGEKJ0df
4mJRHbzsBgC82/rQLLEON/kAn30yuZquv6ocVJRlGs69g2F8wmD5hjnWf8ok
C74jZkHLtvzAdmEoMoX3sZdkbu2ND+oTP7bDaluo4vq6UFUItNkX60r04CL7
DBjhdF0TGr/ekIdA7tEOdqtGMJ03qPsOi1M0+FKKpCdX7mPH9FjdS+T5cSkA
u4W2rsmR4Hh85a1KbDBOfzNbUN/Q+U5lDCc0VEUhRbV6r/obdrqjSNjbhsom
0A9PwaXpoPzt0MsFcpHAeGWoseCCBwV1zN7y1SQggRZXYJaqLO+pR6XarSiO
rTRCvfkpS6710cd21E6enobj+6rXZy69A1Gt9aAIMPQ2LPL8qu0DOIlooiMM
DN98FDYpg2Xhz3FEdzoo0jAx9ed61HnJK4nB4tz8dxONQdCKl5M1gC3b33g/
/WrWFpNeu4hRapVh5vHybVNnb8n6qtHNSUahjhOIlHA79L0QlZlPw2fvM+dN
Cpu+DR+JwK1XyyHGfE3RYZiDVVaUmStpYLITaVGgfBSsQug2IWJhdgBOl6Bc
HAMfKOXjXMhRbNiHkBLO+eadM/R5qlIjAhaB/fbsDTmCou1soXArSN0e5nh2
CG/NHwaWQaNv+rRm8316u9j7BufHmpRgJLhgvGvLnLy47as6GStXh2VHqYWa
j4d1bpxjzMdvQ6Akz6Yb5VL7nt9gSsHTbujAhW7ZZgAMx9oGNWCCT7VUZ9dL
zxU6mt89IDG5on2c+na1UaqtzgWhF+lwvFt19D+A9m2g23SmBudH3WrhvtPF
s229B+0CBHs8rkZAes1cHBFJSucbamxhPj8E8WMOsVO1njl5pV2O5ShIruqr
Qgej1yr7kVZeIrO/EAmzw0AcUiD6xK9741CTpJ1lAFh7EjvcIHpYXKn5Orfa
CJmnYsjDgFar+EJrcwY99xn33CigIgH5A1qy59ISJjKFzQWZZ6IdIsnYYsAv
GHgCGmEpZM9b0z5HWP5NuyF6yG6eXdY9YZH0ChqCF8qY0pMmIXjKJuKa6PAy
tGeUz6njDJCn650161XL8PHKfQLpWeRa53N7ELGaWeN9yEyLnX9voeIRUicn
7XfEenLoFyOKNfyOJERfi/zii2B9iZtvIDlCezj8SpBxIMapx9FbN2pnlcLx
Kur8TEmxRaKdTBL9ewwd4eTdlSTbCfcnSmn8Hh+XH/oizys9MZ4Q8m/iz3Mm
Wd6Oo601xSBLSZRTBVk+CQ7vgItvqXsn2gLkS1/4rvfoSzP7w3JYt+8AXXbM
aIyVqyaueNiLX9/DE2rdfFs68L00XkVH479cItKwCbSrBx95qdgza11Timal
G2hgABezjdwr6OZPp1XtC+EM8yREu2TlSGlc3JK5ytBE28jJB/V0fMkBInN7
GiLv8U4mzwwlCC6G/tnB3wyIAEV1R/xfZ8SgbVF5xAn/f5wNsy65Ptnh0DNl
D/Rxkrg6w59RhYczHgXaehbK7qLAI33/K/UMLKbXdLtwCtILR82VCId2mnU3
/ry4Sjgj11hKylQAusgNZAyPTEV58YxCLa5gEGWmyxQTodvgcFaRGs9e5dXd
3VyxMWjuUQJQQ0M+3YwjJoD40ie6UM7qWsdVdHKjug8tg+1fLlgSzkAZCeWV
MjErw+Xh1DOcg1uyqeD71AfMjb+HJJrEWlFzng5CsRSGi1kW2VAUz+B//Zpk
hFELf3m2xwEiWhisQxTF+oxYk6uWlbWZ1AEb6k/931REMpiNGC87Q95O13+P
4JZSfp5T/fcoFSByuTOfpVa911iZzwG/WAOfCxLMlBDspkqiVrZDhXyYxHyk
Z2M4s9rtUCOVFSNXiNQ5D0MrSNPCVe+f0rTF/EEGLfBmgZNJmvwJzqnFxk1i
Eh0WRdmpbCP9VvNsRIM7rIVtARHqc5ptZ3ava7UkxlRZJJMK7T53mC1RtX9X
1p2HyXLvuzbfadZ+WCBnFSOuyLp6S5NJmcymEPFc1AU+1ngjGhZPoqBabe4W
Goag6heN21msOfJWdmof7yFrfZ6+U2HK3z1MphhCqHYsUxeVGW0DpS+Ifhju
ppVlFKWCAR2hSd+hTh6nvrfMv497bPtDQuIJsYHxS/V/LOFQdo9TXMBAWeNt
DrW169iYHj1AnwHXICBDdHXmPRlglkpY6VBT1zpzAb1NqbAhN55r+yCAnJ4Z
RMI2oLd7oVce4BNGVkdNr7bPXQrIonBaa63WhOReR4ZCBuu7sswZ+53+m3ne
RsclmIY1t9BhIUK2fFborodObbAzbev6R4xbi7HTtoz5R0u+kjUdVmh8eFJW
hO177kOr4/k8Cupi7XMtifIbrWQg1/Kv/jMYn6dYN8XECiosF1MBrzlTf/Ln
owy7wwDLLabT9r9yN0BLLE8zpPZ/5hNuLyarB5BO3mupY9C836tcV9ko41T0
aDBqhESlOzHDpwvvWVv6satp4GwlTzqEniYxDdmwZvSpGGm27b1v37SeRX0N
fdnq87AAlHIz9CUIXmd2ksGyPOlglykzN1mLgPSyuGYworY7Lb9+7zZA0Xoj
nsHXxOXJv0bLRiIAllv/m+hp7dcgSMJ2t2vPO1onli+ESNvxE7DZtHJhcxEp
IWqwc3gKft+Dh3E166CwJSjGD6jGYMH797ujUW9Hk8P+IjracXWoxbvRqMM2
jdRd8c0l2IQI2DQgruscfJey6+pV8/ryeBe6tDgbUFOiAu61v8XlUhEOJPy2
6awsaEbqV+vrKjKAGLv6FQjO2N33nmpGgV7bMysbrdjUbIYc9/VhYn6qPVu5
I8vdM8UnZwtwyIDNUPFQbPkYJTJDFoiHQD60vWz0ulWWjkyYdYFn/0Lt658h
aEnML6CG00AHfOh9tA/Yv3Wa1nPlhgdXO1Suvi5yDBM1htxwe1YFhJBXuwqd
CXA0W47AzqPvZADmTpZi/1XRrczReN4UhAzxecHXZyR8IPXF9RW5i26B/oOQ
ejzKyV82R1qTUA3V1WJWe/L4UkVF5fEgIRE7pA+M63ixVVH3JDlirEZGt8lY
BgQwcR8SCuXvBEwOQOV20kSQtSZPLTHiz2Wsmc1KGqE+3QbduEzUfpibTc1e
k5XP19WRB9ncKrguoZTossikx0kOMK8T/dpBMckLFXDq9YwjyKa7tagdWxHt
JDcgBHLCjw7+zuWaFiOw8yxwH51qTo7WTzsrlsm3rHLJqN1VhidztraJXJTL
wsmVOu5Oi1qOLfyNaDwe29OWFOUXMAkQpIAAGPley1GpyDPMpeotG/L6QTxG
3Fooaoftl4eqEdUL5lejDsKPLo6CiER1sfbV1IrMYqw7IdHQCXfvjMaTCa8V
YrxcefEe+JfFKlLlFp3rqSfFuWnFWRL78PEpRxV1EiAYpl1E9M9TBR2yVrEi
Suzm8b4nrAxmMyJ2c+olyVnOMJqOn4dcyOSE834br3O3m+CmIXTGI4hpyeU4
NiNYUEX9eX2Re33EWyGyE1V4eazXEqj2JdMpPlok47TZFYNvyK4gINSrIZro
tecsjippvpuSKz41ocOT/da4KXTjuD8eHw5RH/ZnBGd9ID2nlOzc9WvQMc/3
+ZsYLMeHSeZuwRNKp6rNvsF2vkhF3sjedzMJgwxQ87s5GUd4owvktvr6XkkK
OSsvmCyXIguzK6Hadb9imuh1w1u1FDW+OhGqOznjjpq0u+bGfLBFoqPp++7J
xxcPlgINvz5jar9/oDCdpbt/JykPKzafpsXAuN7PdShCRbJg0nfPd3HtdlGk
zR3qOkxlmzA1SDLDJXLLiAxlUJijLfH8v5NHMcxjYn+o932ZL0z7ISa7SRrn
gJbAXZMPoxwInM9H/aFzKb1F+7K+b0UXDq2KGUEINAQMlG8XMneb3FyYxr6F
V2RUhojbAOjPkBvrlCHm5uhmk5tumUl/2l0RavA0nDmq9DvzAoX7q4f0BHW6
KOjxzwB76AfS0yn56YNg4HOaC149k5QD0/uZYHYUqOjmJJymFmP1DFjaNa+i
udu119TmZchb6hDL0jY9Bc6uitJf/pNqRYngR1fSFEQ+Plg2kYeNcQt/Xmbn
9KB/ZbWImWP7ADPlRk3jQESDoPJdac4sMogtCzCSR61S+qm9gxg93s6x7k3x
gZ1D/L6wYtWyTKa6l4isDhjfruzt4Qj4XgR2OPtSh8BRWO6XBaeRDYzsNMJS
RPfgD3tzKc9griuoN7AwidW1e852x7e1hZUXca3HEPC4f/8mzXMv4QqyW+Xh
a9e2FOzIHH3vi8e6xFIKGIWlZ8zEjvAAZ+24kCqn3QuzHiv6AuLr7maR9Ngr
jTA057eALNAA54q/W75VVOQph5GPXaob6rbsed8hhE7sw7Kyjt76nrY5MVca
JtFrfU0fwc4593Kk9YMuCK4UsjFFxsakMirjPpmOr0xbTmdS8M9CeEV6UzAE
uzk/63GXrVdw18gdfOWj1N4/Z6T0rcNtt/c35cAkX0/MkQEaNCi6CeZUONZ8
U7GIWNGuR/LdQBNzeVmsmum8uJeWxOh0x9AWYc6j6TZmkJRpg4Rry+zATjLs
Gp7B0QGlaiSwJ7EodhKhba3rGEmqUUZ1YZvJsGwACNDSACz0GCevKRYIQtrv
lgJuZ01JGWHMvOs4WlD4/YvFkSNwIwUju99w+DKrYFuH9feX1Ry6MmyPSBAD
Dg2lybapLrtkMflx5bhXPKBNhhqtmaRSEf4fBz2lHy8gKF2mdbiAC5qI9z2W
s3k1w0GoeViLCpVYQdPxe4D1sDVGvJN4JKjtRI52O/+49Ug4TLcBJHx2p3M/
LwZne6uzaEuz8aOYj0TkHbs1CzvDO2sWBKhZouNCZUUfpVHP7TPlYKnzeat0
/IW/u4YJlBNTCEWNu85gjzlW7uBmhgbJ50bqlgfQryr04CHDnJGKQOhvA53F
5DJ5nAMTkaKPoeOaEjELOl6ejN+3r6cWUHUKtbVsdWpE5jYZAYd6pj/I4fGk
FV8Vi1UHipaH7knuCzvUWkd/WJrpZqzrhsthKAEJqcQpT5B8yhhHC7SDnawT
A/i//Nx5UsSkDytjUKL2nor66R+eZdrbk7qldszw34ZHrKV/8hBjQSYZnvOx
zr2HH+XDXc4EhhfROFW+hgjug3x7fsmLWIEvPf09r0SHOp14SgFAS5jW2ODK
EpFFhX2urGccwoIathjYQT8YUS9TZCDn+G2yQLA0wy+Uw7MwLGpAzT4P+gim
1MmBFVgBSj/o4DRm9mDDS7+ZFzhZYfOhfJsMnRxu4ue2ZP1I2OUZ6FdTyy00
vNo39nBgDRuUP4G3Vg/f9gDePN0X2ODpAJCu0ukfOVRSCHfD6IiUvfeBXx8C
sTtsC8EiGEYozLwU97nqK7B8ANA98QznIZ0ZmWcafCg8Dk50GmVVwSBHf6EH
/jX3TbLsM2Xx+xWVsCBa+AnlZE0YOa51eCjb64RJUyDy/5HNzgzNJDmAc1eW
j99bw8D3x5bjDTqAXbAc80gQyY8P+EQ6MFX3rB5iUfvjZnFnjt5K2hegq0od
Yc/7nJdeLtrkwJ/ay6bOIhvhfy/2gCYQtb0zGYRXaFk6gup/CquBkM4h/5uf
1dZArtBovp4Yp4uqB3b9CQR/keV/GTlC9+Kxe0KOeb5yPrAgj/31muQCA1qw
tSLUbyuOKfYaqp+dYPN+Co2RJtPXkz/pvzAIOL13zoOPZUVxUyCaOHQIYSz9
ra+MAenjLuF2XId6pB7d6sBNOq4JwLDN6yQ545skRoTlYW/ngiTcAjuAxjyq
JQGkEn/jfwWlTZlQMCqC8PDzBR6x64BLz/XvOprckGJ8d+LMlMpra3QwtL57
Z412c1dmqOm2utRHamWEJaN7Ocmrx0OKOukJ+VR1WAOeJewnk3T0C01Phld0
aBnJXZXVxQP3CDihvlEdJsWmkRDAh6XpemR3w34+3iwcN40/MWEP6xeLEe+6
vYCQFlHfGahtFAEgMVMvGoPa2F/bYqVD7hI+yVx3bCA91gcN8w1hzYr236f3
u8dG6aF5qE/Wm4LEyKu+PVAG+MbN5p9Wa4VSw4W1iLIA5GFjlU6MBO7igS88
XhxWybK/T9ssUGb6COLUEc5voz2iVCfD6acMobCnXmg3vGtgzTJOYQp0rc8l
NkVrjIh5esjhMc2y1854anwTgnWDR59NvTK6TQIFcGBAxAYaXIbeOIcWvyqw
r+bJg/vz6JPEPIUq0O4OLKSbgNIxJsf78hhWqXA41FAx+GvzEN5BrpNeKUMp
QmudvHLLoTLQA8Jio93f0wx5ucXM8mPhw31ZPC/lmXNATsiPHAQLAcDFxXnr
p7yY8t+sbJYlbRlFP63Hh/Bmcp6kxzMRnnqinpeUQrfifLiKTkmxMEKoi9mg
+sVlXOXQJQMEHZXEep0mpDCn/LB54jZjFaFI4Yr0yZtZgxRKjhAjryuMjx8C
p+9hI8XZcIHfedrpmU2oVTm1d7L/+M11qux/6Ev9KURufFmUfPlPdo6Kk3HX
F24cy2CdgHyUeEc8l9fHL4aiHdtuqdrHYnNis3554Skw+YFxSqGBH39uM6nk
AqXoCdCOOUhfUFUgq4l2sWOouz3TbIyN89YXqfZDAlH1XaeuylpZq4lUvRVP
4NqlzM0C6UEXq65vRpFuk2D7bwtsEZMWOkm10OzglfB+OxDXjq6KqKc/9Hm5
CdMtv6KiCRPHGyqvfrzS62tM18HUC0Xjby2ulfPMoeZONznjF4kP8MxrDBBK
TRxkXcKS9YPflmNj0ZIlK9Z+SarVOO1i1DFRt1to7w+NoqBW4909txGK38gI
wgeJkJSrqP0e/+75BU7E5mxRatovtUKLQLz/I2z6F2fBJgpHrStMNldrIzxv
rnk/LaxAnq8UBDI2Mr1XdWnJOpfFvBHCW3bxDhBYT0nCjAeitomrEXoWV2l0
yZ8e9e6eT/SvyxnJbr/ulKDmzJH8ccuMj2xlQfV77bUz6P00+CkeViQup3Q5
CghMR+KrAbfSpaA/txkW3Pq92bwSYQyr4lltzj1FpEq6H2xx1w7URZVRCkkY
9wpq4z0GvZP1raBC0YmX7oYfRPtdkylrwNpuPT4qjhkwQcpOy8zfvbpbf3Ph
HqGO6lQYU0eSAxoCmJTYvUX9LjbrkHxkc6LkeRdXG5o/B683cYq0qVG/+CZ3
j9PMAFlQfBln26XUqzWA5uv1T4RaYPAmHhUbIpAKFCftEfNgRSwvNzagOs3e
VkmFZOnX2hc4m/sXdU46CUPZ4v0eheKU7SpNtbv+qK3I6IOvW/grwBh3FUjj
1LxVgdyUpERlsRc3f+WHf0eeyVOmXwTS2k2pCSD/foYxLDa/afFj2Ql8YffZ
L2p++y5oF4RffgHuoKyh+I5SsWpP5lF1QHlTrmvNmSicBcr7XKB1AMs2mGXU
kSuUynBT0bda/9vJvIfBi2wVoP7CjPI4Or/REGTYqmjbe3Vy6u5b6/xHeZji
2YqRKcMaDVIJi0fsq+utJLOwIx0D+nKCX82CYYKhyhhsJGf/eceR88FlHrlY
DA3VCLt0on6Jsod0plvm3pNpE8AmQV/9gXUWbZs9iU5VB98AQ6C0DWB4/k0F
ff/X8RmrVLPrevd4ZKQuy53uKEf93N5lKqKdpUsK4C1+QuvbhcfTQyy/8d2B
b6GkSQ1t2kUON4SXwNNRJTUb/NSXuNgA3FItelf7f1K0+VKzRdQiofnvk40q
idXmXZl6FGzXAMkDDFH0J3WXxiL3gFODnI7wlUVNCDUZOP5MQ+pF0/g2fLkU
cnz8whKYZkxEk4TLkn6I/nzHZzX88wybyGO3+8IlvMvKoeWZKdJ/qAins8Tv
RHWgCGx7mm90rsha8pdt5aTsLaw4/4WQZc50kEPK5FpR3G8x03YK9zANLTJe
V8/iaaVBkAlIBmSga+1iOKlKyoDBBBxc2tGpGHp8loetlgcwUafeuzuIlIyX
rXEsbCwtsBn9sj6sHKUTJ59YBK2B9aq/GBUtUL57pGdam20xXp4Zd6tgnwd/
5O1PykG75TggnOz7AQuxlqb4HmLMqKIIxhhecPR0YYvhYTJ8NN7gd6oSfA4v
8OAjUCF0gXqRjrGygtQFAWu+Y1XuaZdww81BSuMc9DklSx4G/0qP/18R089/
4HIpB+KAPx9HLW/6T3CiKQPiNGB8totptC4Pe+Io6wMX1IXFcxpVo5kAhceY
NKfp6in6rUhbNXEXTmvazKm1UPYwuNDipQpmConVz524MMUnIRj1Lrs0UX6c
apGW4t71tN+n7qC6N5y2evJ7NZzrMP+46BL+yPCR9vodi9py5naVJJ0Y3Con
Lp8sI23S1L5OatH9aGfLME2wXtYhwP5b+w2bOUQIRw5nOF4qZumrg3ftQkWD
DrHueVK4NCDrxCNg8e162IjLxZ2IZt50g+K6J2CK7hE77yGNGJRt0VPyQdoT
oZw/DfOW6VXN5bhnXQ5bvjSNL1lrpTcu36Q3NU84Q4KLzXrEtBbJuKEhmMp6
Sk1LaI8uXtF3P2hqp29x5TGln2mfZ5GDJH/a7MxZKlLb0X3i9SYmAJ7MR9Ko
jKumnvMGUloJbbISn/h/zGS5nMBnuo0Yh4qP4RRjfqLlAd/6Kqv2sFAZtAjD
GqeuOlOVynObC74XLyiHnsy6fN4YYZq89S4nPrdfR7h6OynRusp9kTRnzMwr
+VzKIPnZ6Hsrdxx262AlQ0rkF2HkBYc8lSpHcyo4JfJlN+5WiL4Tw6jGWXpJ
psEQ8SDaVkWi/uN3uPQe9/Yep/+3VdUwLe2whyoJUMU2j8Y7LMbGVhxPlvU9
0ZPTZSU93z5RoW4OnDKtk4GPqK3tf+eJLyByneCRKnwpBEtG1aynvRaXnZRl
vsLzCGsAKJAU5VlAQoaxabDx1+xKfHDECGcDOa5DJ5rFAw439gXXY40e7xfJ
i5hquCUJ7f5F/wmQY2R9DgkvVACRCidJLQeVxU2MIGvNVh3LinNtclpNfYJK
icn9VYuq8xcZQkmq8ePDCXim5NE98hlZtzCRH79nW+dpBNE8RCauOM50dr+H
+hsL2Byt3qC7UfG53jjSmL1gMfS27YncxI/jwDa4WwQcmKoBIYjnI62o2Ocu
AKV6Ke3+HOlbz15ZV/8jY3xebZGQUi3y+pUbwHSOgOx344d7jLrXEDYMIxQT
dosOPuSQds8O7i78f8NRYmr5Nzms93oshsGhlZhlvcx56zuKYxoDEw+MHUKu
ajefxn8C2mJpU2+iAlPsMK4UJwKTweHRbPeQkL1kr/5mKxfGm5rr+eWqC++H
z7imnftYfGjArVi/hbOtedLx8V/Pg9A087ybnWNfh/p4UbqbXHgO0dMo7ioX
rlNgUSc4Ps0ncb3PIBEWBRkuM5/n3jdjEjnVVT+Sce9b0DX9bcofYvOU6Kbq
mniFtEODlj5bgK06g7d4OBtco6HMrchPyinwpN9NRt9kDAuQXL2SNbXSCRMR
or4Slj+Xs5RBxI1QreeMNM3xuEE3neCTXDKai9Hf/nbrBbuGTxs94XIx6yzN
j+pNs1xJMrwSYl0UVSJP5oQlqa1Kg2U9BEmQAgxZn8BapLHgw80nOx7UAtXA
Bf+VgLMjsLQSTugW4pciNvJQzsDHp76ngc38xnB2YjhDsevJFVlijSBTd/p7
iAScr9CkDizHHRoDMzqS1LqxqCHk0rNrRIW9hmXpE45YtMNQZ+eu5Ji6PhIx
aI+xUoqK6e6cJxbteNrOt2wGIyxN0uLntZtxQqeVKYQQtePmrjb88EL5/LF7
A/O/p+8e9iW/N7LTLaxsKRyCxRC60b6DZe6jDTZvK5tJk+gQp1RsiIjeAIOg
HNB8JzBwpLqOHJv6owYlY/nw4FFgP5ILestgBDWvJxG7VOXbMl/xESWTTbYz
/I5mnrvHEBKBDJDyd80wQEUGPbRmjoKI3g9MzFDb4IJ/kaJV8l4LZr3MiTsY
qfyNSrcaItRfA0K29TZjMp2mJN/7+g26rv9qzbjsCFLdDCeiAbkGjot2g0Jf
qrDuzLFzByhJ2S8cMmleYEljM9QYhE32XME/UAzMqSUJu1gQu44gty31t0/T
ztVVO+eZpyQc20A4AglCL6rgyh+MoPDpjJ3W9ebgIWIAJ2QfCIzD73t+1mGg
eYH9T1ZOLdpmEToW9TS9P6BCCIWQLo0LF+5zVrRgmTh9tBSE+bE2uuuvMuzL
eATShrqRThLroVzWlhCOkTxhrIVLCaJ5crW+YPF4EsgA+xepJ62ypkR+ONtF
zAqgs/m4PY5Zo1D/2aROwq6yL51s+GiA8NIphynogXQUbQ0tktovwzaDXIET
rudZcW2/VLktFWkjR4gu7bLEiowxgs/GRYD/KSP8w3ahfLtBk8ZPyZ7I6e7j
EUZK35XELpKON9e4OHWT994I50UOsdpO0jPzkxUPyUBuAlBHU7R+AlhM3XK+
oFaegVHbrhSAlVGJOqZUSxShSd//X+dZ6Us8hSl2+A8ZOaRglO5HNTv8kBdR
hI+G5+Ty9/Z4afgUcsAcEFMid8E7e2td3Gk7srMeGMT9Y+AdxDI3zdcb8m3Q
DQbYbxjpytl+EIX1ijrul7rFjq6bo67/fujdm8C0D5sbnEjiXjcFZdQIj5My
GWhmTwXoa5LjZOs9dZMr22xBZU7PlePbp+L6+4uctTTIZYYJcAENV29urh9W
N1b3EeWQxdBow/M5SNkwlAsXKIPM4cWooX8NxoHkUXcALgz/aZCpfG3bQ3zF
AdXma3l7asFaajGloQjSpvoXXLNwjlX7nBs8Y5cV48mjW/SGCWRjQDMhY2Rk
LJXBaqIe42c2JwkTLUiLbMV6KC8SNFbB2z+zgOemBZkKrtCwdtwdsOt7wQwF
NZlKS3IT0K2UHF3+sxbDwiO4NWZDD+pUnkqWAWBxbjs1sMsGyF0OtFFvunP+
jdvqkgZrAPzCdhkLltYgtiQepODvI9Q+3FBu2JmT7zanyebex7Gmt+vYCEbb
ljsJnhwLt++pb/46OwSIndPaprmVP233gzbAx65IT8aLv4MU1ASoWfSCZn0g
Xzx8qfqcloeU4A0HzsYivE5oSrN+qbsqrk1S3aJNRfSeJnYsEDIEWFqBUwzo
nsUsKt3CzsWyQgOLrkUceRqMdoZtrQhtSMUG7Cc23rJzFYT9r9b4FlwNaGJ1
jxddMILIJ4HCqUMx5NVWD9uQu1VB5FOWnWuRUed9WP2v+Iz+vBGbw5B7jZ8Y
gBB9jwdd7BMPmOL2ow5fV9IcMCrm+BaTOfhCoLyrAixiB/rWbtlfS4ebO1pq
THTSvW0G9GWpiV5PRuedd1EEqwV9fj/KWnE7XLGwhiqdxFvRsfLoIqJNuuv/
S5FZKNSTX/zlUSX2X/wPDmoyTGH8xZhZvGPd2g6ZIO9u3JOWEmTID0syRHys
EEaJfwiPFATsmQtU6KJwJUW3PRXx5ZOu2N4O0cys3S/dePq6JESBgP+l/zBM
WW9viTIsTgVQ17sb4I6QnJBgfveDEuJlu6r8jkNNU2Iku322K21zhGfGTB4i
uKy2LgJc7ZfOOl9PemX7zvnDTQLG/xlnmYiif84uDriVDWiR4HOHTbZt/0FP
1qbs0yTR8czbTnw1nAU9hkQYlRQHCKGgvU/IKYJIVX0Qhn5n4QlNrZmWUsIs
IDaEoHnmftdpudqVFoume9K4WchUysymlmaLUgVDq/Wm4SLMW49IF8IWaqCk
UcuxdT3jTd6sXg4vfGNrlKzfxbtZJ9F8tx7WwlgqdHgdsYLHzl8+2fgM4axS
J6BG59hXU14IBF267HfEOD1Ah7UQqelFh1GJbj/J7VVq0vV+LlW9Gi4v7gQF
V7paJ74tN8urlf9YV4Rhagd084R4hAZohx8WG93fW+MPv8j6WSqx0sM10qfl
lEdXRxYHoE6S5u5BI0AFjIdCUx4GFRcFK/QexD69XZqT179uy92YvhFqa9YM
zSNEKGUV0DJ7vUVkgwDCovz2KZFrMdolywadzR/Ai2oKDy7UZ1fTfCo+M7gX
pJrINdy2xVhwi9PkZJj02pMIY0IUXOvs11EFkltquZKjeHk7bOm1Hq0nvKc9
iwX3jzlX91BcYTTvkXut8wCb6AGk/9SpoYoDPBRcXGJjwnw3eYRI5+pplA1P
Y7lmzX43x71GkdLryDoWAlgGYPPInYQBXto0l0tQMCdUwcxDNF0NbDjeEzcB
DeEIl+LI9C4XK8oFEbqLQMXzuuAAbgWOSUV36GhzPjCzBFIpqeC9Br0akPwP
LoLzU3P+WOAdhXUGrEMEuKFo1v2DigDgT2P0NAc+FTdkSde2tK0dNHiDL/kp
xvHfSFQFnGtN7To/mLvud09TUR48Sntz3ZVnsWVNSHFvNTP2x/jlF3l7xNGn
1g4Dpu2/EIARIsdOaoDwZEzQXF1stbSOhfYO86nUILbgs4DlPr7IzUvw4suE
MuQDi9BmOYpr9QVWt208foFmrIEZR82BJ1HEovOT0yi16eZ2Lr9qAYqJTUxw
qwSUXSPyj+RezBT2Nu5fIqlQRmNEfBAJEi8iIX3kJ2TgvUAMebkUduTBkBPG
X77Y5Nqbc7NzQVsQLwPMzIgwG6fmEG514MW8IvVc/u9cP7g6D5mZpaO/+dXt
7zFY2YTETLqNZOLMW3+6fxTQzW0VKxcBDaCFx5xGnpThNxzKSnWIGSjE4q2W
pFIRF9UfhcgRN+gA1unP4u6pMYQBld+A3KbfReYeKhi6b+kTL4f3efRX7Rku
A6IClWGZc/+hnEuL82ua6dxctw2fyYaO6sE1jVq5dC1lE2VWvNHHbpu+rpf2
TLb6v9P76fEKb9EPNBRRI5EmuKhd2M7POyYLxrn8xD9bIo8I967wYEfKRUBq
Qh3g9P+QrTlYwiPlPQEsD9AmzUOTUUMa+e/egpUFzbiETGv3+Ap6dc6QI1qi
uCNAonLF1dQsq3szRExwP2da/1qH3ass8xnbyu8YJTgGIWJ2owRQGHASbG9e
om0EiO2eRCO9mA8PlaeW8l/50Xdr+Uvub51OmBDuhv+5Cqslmw9XfdynlhCc
YQ2YCB64p0QCNNAfD+BO/WTGbY2x1/ZROIAVObi5xyCgwEkvhRoYXEIY/7hi
w9Ea2pHJIH6ARYzpIzHZoXUPNBlWnwXXazUEr4E3zKkuBGFq7X0RCuBMmVhm
gPH18siuQHCWBV+0amE5cskMe/48ObJCvZCq5KTz7A61X6hunSSXuwWxHvTV
oGFDK+NeeUBhQyPwwtYQz94iP5nqD3AigNsMDRYUzbBWXdVykqx+U+Ux4EXq
6DoCeY4vcu5DmEQP0uLmoUkY65KXEanBLrn1laCEiOmYLz26hpM55mTadBu+
OYsIw1ctnEfYOmu9bTxS2gqYIk8rFbLQjOeMBy3jrDTVW3Zidb1XMA/OgM93
jYQhWVIBUc/XuoJNFWoa1le+eTC4+cMbRYZQ/qgwK9dlmY7YD1ozcAWSEF39
IWMjrMl/wZfT3Uu43dplDBc7mb1PNnoLhBXpArju/uE8wK2WS2Tj93KS/8tc
d0swMXvp8P1mCpizqTjd1PdiJxr1Yyw28LNbx7OoW4TvIDqNni8QcFKmWpFK
Fji5HB4qq8g1zSzYn95aGnP8FIYnnXTuO7Ghxk/0DhKJRgyKTnaQZes6BK3Y
L+vUzXNJl1GVGGCExWMqFjEBRC8yX/yJMEfAWH4y5wI8Nq+eR5tff006KfN/
uKs0lte4fm8tTsEIpWOq356+3Egv4RXmKveEmZACcV7DTOBHzbO008GFiAWy
IEyWpNSODQhplc+hOQRRBideS6Z7BXyAspGBgIuH7srKl5YAQy8zkrElC9US
Fz4Zb/t7DIbs7V1whQKQXpwZGuC9DLw+u8Zn79PusEZOfbd1CWyDuzSOO0l4
XQkbQXXz+sXGpORMmiVWhj7U3qVRqpxCaTu8xAEenvooQNLou6AAl8dB0vtJ
b1w1vMziLGzrVwxl5PqsbvaQxss5EWUXrXP1JGJsXSnJKBXCuRZD4MQr3C30
x3QYAsdXnTbB+ignHEoUg1LMuOQjVTTzZ9xI+SswNBMgZWOKGOc5Bsfr5XK+
jHiLeWGDV8qpF4W/L6P8j0RoyWO8POMxX08s8uOti5rdkRa1V8JDWcSKEO9A
/SurogDvwgLaCe1XrwL4DeXQpbUlbO5+UbaCpIieWU4fmhCKoU5vhLaV7+zm
m7O55sXJc7ihTurSCTjkNUYduqPwA+c81JTdz8gXTjvOOddeNKoe/OSEU3nA
vaAPm3Cs87pSk32MzXDGQn850Cp6EQeyoOtFDr1RjlFR/51IMKqV1JyC1MhS
pyRgusksptn1cxbE3gIf0MtUUwSN17gW7L+9P6UQuE1ueH/vyAopzFsD+rZR
D8EAFsgsQPByjMNfEpai1ZEgXRvPd58bZGr4G+Ay3l0Ai75mQfFaauVuEXHC
mwzB3Ovzjry3Gxvqrzd0Peu4jSyBvEghD+s/njtUfk84egzXaKCiyFbm4fwt
aiOL/zKjlwnbbQ9lYR6e0Ud6Vum0nEtz32zBtSztDwjsUK4+KxCUPgES8K0p
yiFufq57LKGHlaEqiq7n5EBE8Ely0Un/t4u46MvMwRJeYQDp4+32qNumfyy6
Lu4z+PXWl3l38/YTEZnIXZlUNvaV9lmhzerVJar0Dq41e6mek6F/7Fd48J36
4mSVZTHTSC6SVFGSZmHIfLOe/cDCnObiJG2untMLHZU0KTPyBrMtYS0yBhF9
ugjlh7bmkTsuDjVILbducaNL4upJIApl2I2xpwiGsxElIoFRLsnSRo1ujmxn
65nuqhIoqMU72dlRHbWCg4bWz+r0O94r1EI2QEXZKE6VOTJY3V9+DFkBvmLh
E5ca+Mi9mQMbAOuXp7KIhSTM3mZup5hhEmw4Hm/xywEsIkXie1w0ZB1Y9Nka
tzQGoHDu099BMGCBuhj9U4T+D5+mTnOGnHwBAZa3LhAe5SVXqe/6dmfma5Jz
pGfNHLXvUddEFmM/jZ7tSLRYP+OHyhWSf6251kybJ1W7kUk1MuKaQZjCAlrT
2TlVBkl/vE74zo7cyejMMlxAp9evBhMLpTpEsifu8LcN1rQmn0Or9+iCvP9Z
qk8RHfAG/RNLsADVNHesb0TCje6017ed3ci28IGWZ9drnQwQffjoYoAqDVjF
ORjeV2kbzsFre0BrtELmhqLuR+bQfANP+C57XvYHhphtEfHp6ci+PGc/wToK
OzVqB2mCfxEEAKGIByz27sfh0sFNL8hUnuw6Wjiyml4G5MRl++/r6rRAeuY4
ARw5KDjBi7GewIEpmBcnqtY0NAIGh79jkQkIbzI9Cw4mU9E9Nq4Tl5+dsBah
yfaFWHWIOSWAFkKpV+YmIsF0NOnrBB5dSwIUvtvv9Fq6vXredPjzYyXn36kU
ClPYOc4kPUgYgaNOm4QEhbBPBUzJ1TFNKziDEy30Xtbv5y3+EtTJ5isTvCbI
br96KEHeDKrqJYIB92HqRrwYmnHDpReOvXT/Hy6PrOeDgamccNKulS+uQp65
Ix56Agjf8NPmcsjO8eRvzMHxgUk6Q2cwX2CnJWKj+1ZgPcLGest5KuxI6ITP
XVIW7HticegPKvipCrwfWwWQdzsmXpc+mmCzQkfgG8/rWZpjdp0RbW+tluUV
TLFtUupaFPvZbgrJziD6cylVa1dK91u27Tjh9/PDpVg8+j64Yc0PuHMfIUJl
uGcfg6w75Als/Ce0DAZTxwKl5/rYo3Yzu598L5NtWVNEJKrpSoa8dOJf2O1f
TdGpuY1pfNmGNJMy+hITR9UlkNauM1uYVFWUc4srUD5BRfH0xoAQBjnGpujH
iISxnhTllcf5D5yd7zjkr4I+FIBkcyV4rPTVpPGF3ARgdIXqjhP35J6WZolQ
+ErA74FFK7RUdDYTNtXoxkGN80tUmkokTNpIOUlKxf5c+7+6UKptsrcFnqA1
n/UsrkaJFd5HfWJzC2eCETJHwF3iu0RCkGWogSLAsWfq03GOlR7aGkWdaK0a
A0/o3ICTUQmXmma0GxFCTQI//x8IA85DlebeZ1lrxleA5xABW8OMfCHetsq5
dq67wyNyeytlnQUJVEM0Ix2n9QcktV51TWE8VMmp/45lLCYAaZmiYbKk0TEK
Uin/DUD/o/T3YWz7osogl4We2WM3jkUVWtXTMbqQgj59NXli9ZBH1/CgrI8l
FtzAx/VfFQokWObEgON9pHrtBJzPdGF+/uJwss5IUK2eEqzC5PuNw8uhYMF8
bws6wDkx9NGynyPEqH09VxBl+yYk4R+mb3K1BpuXG1cjUL49wJdkSVuvti4q
sbxNQfFBc8bjgAAeTEK6EqWTDsEQPSjPIXUwr0De9YxcCpBN1nxKp4rYNw1R
ucTVKOpYzerRd3MGlmoLFrb3rR1OZoxlM4PxTWYK94Qr8rCVow7hJ4gTdzPp
4DoKVta9h7zGGHkB4B/ZYD4LIPinHGhRxJgKK6RM/nhpwaB1GoEra5pSDWAb
fe1zoyBLDdht5F0BziMXqb6cNi4snQEfMRur7PND/7ORXeerBMYRl8UdxPWC
+JfxVK/zCjHWna9FLvDz1eUGrNJx987/UYacrKhrg1MihzCHHa7LFrJYgVQN
kM8TWBXe8n4VN1MDwwCuMf+nJtalgWx5Q13+BysYJt4AHtuQbJ53stQX+8S4
AfFKP5iufOlRUEt2bNNPh+R7KZ6RfEx/xa1CanqQgSSozVUm+EZs7xrZu4B4
ysZ+DEE4Y0pbORknBiqMMKgOVNuopP+GAe8YulTrfEi/CayL88o1/2+A7vG6
9nX3FbMENsDUcvGjdF96DQ6mdpErctD83Kv0oLdShyf8SZKHFToDYtQ1L16e
MmrgXmEcWVQljSmMrERBjhKb2dcOeZsQZ0xvVNiXAf/x9DI94rGtVYZ8I6aP
vdptGQqNwbuLd3qO80KurIUq8mLcH0TyUOFXu/k82MWgYTrFrV1cUac3EGG1
A7iyuIN0kcKuZ5uJ1XyGFJCKZWeg0WiN+mfuE5Zf542RjzC79HKvsVNdUN0s
deAoi+UENVo7i3IS2IcCZxJNjDI0fcovzW2ONcQOK4NGhGmvQ1G0cna045A7
Y7Q7gBpBZYrsIbc5mMhUfSJnXk+H/XTww0oupljSfL8txD8elGsm8w7CdsTx
XAmKn4ViVmYUMHDd1lKyXipiq4ZFBXu/AYMuZ6aCB+dXJm1lwW0RM+vkgCu+
ExmZyrWwZPop+JMbt4q8uzuoikVVktdaHQMtoZET8M8pFRdzd0F8/lpeEF5J
HXbLKlYZI26umUy4bWKInbwijRauvIccc3uhIrWlQ5q0fep5OVxbUb6A4Xz1
yMEskIazq7zhpAYZASdvKiDMHPJdMySfktgeggWupTHk6r6WFshcvc8dJdow
ZlbXiMX/LfURhJpDZ1HXTnmBENNSQxlk91UuRlx5gwAqtkw3uDXWH17UDhWb
Hbo5DLRmfMTQCkJ6DdZ605DSpcFaXOYmhEpsV5/DxXVFfBu2loM2Vb1dZGdW
KHAXHsL2MFyM/dn7oK88ZqO0L28pdC6mQ5cHgOVDaoRm3MIZLG9O27iuulz9
hmwWp6vYCgYVLnP3Pk4pYlJUuOLZV5+Kp4qvmvCqqU+kjqmKdJg8ybsRU7v6
Lw6e8GiF5LbPHqN92D3HrWYn12+/Drsjsl/FGsEmY0nO7SXnss2GHievpkIh
sHbTC7ccorP1HF4gmFqnuI7GR8qCI5Izq2RegEJTSWwWX+raLwkBtml0yUUs
G6MGo7UtQ17x/fpQ0DzSXM76gWE38dRF5iy7Um4KuJX+hbpGSNEK5txt9ZjY
8gVd7L7E1YeBrDq7rgEQyghncTCM82zOLK/KHg07ttpI2GP+XYIyni9A2J6F
90YhsE/hUHcfgvXOyQm19w/EtQBM6KDpewIVFFTpAuxepPiW5819MbmVN3aE
YkqrIdqzLi6BcxTXmh1OFeQGoOdqP5CM4KItfiT5HYSoMjO45daysnC/XN18
RcuijWJH1OnAQfL3fLPx0qMp3UMsU7aBuVJ4zJPggoIWl4Afi92oHwxd39ws
fnw1pKIdzoJfLAc+srKkL1nghc3bB0sWvOGe8J2CAJ03Y8YHdcatk+PvlEMp
YRj/ITmiMKG+VK3SHqD6277x13TI/ORGe/mq1a5cc370/CoTKgUJzdSLkXZ2
nHuWpIpqbAS0U2L+qxHRtAHjy0QO/gaGduOJPEvxsJbZe13h1ls1Viin5qHM
f3shvD+5AWXAF3sjSd7pFm8DUHnT/Od4SycP0GeeBGWPfX4D4FbULBn8ZHN4
6/+C1KRC7CqC5uz8VhNkRZXHOK2ZDaFM2GuolJBauCITgOZRg7xdkP1dyA2s
Ig2nDrjoP1DWzeQFPyeWy9I7/ly/Uvsf1d5gRzh+yCWnxZHTmI8auxQ47UY5
mGEDqxoqO5neGC8yjvOda+YTkcgHTdzB44lnEg5picF4ncO44reNef/HkyYn
KPVUK0OR/zXlF7DZO7CfHZM09MqZKedvGVNOQSl0qAbOzIO5ePqI9OSw8IG8
BYzrFZ55dtOALHZJTaHiL/bdd3Z0b2Km/oo6Gf4iOMw86Tg5IK3+irb4pVDY
Hg+0NheKgpNNcq+H0ZimqP2h4bD7U8dYHDN7RbINpQxmSy9DzAwpqIDHXhEF
qsHDi5a84kdLi0dXWwlshRPSUTu76ZhUyihh/pEwdnlaO5VGCQRqWUfeEj7D
/UN8DtCP1BWwYIek+Oe2/wUZo2HmKHh/zJmfi9eXYfsToeYI3+cDreb+R0bk
2PhLvZdsR4oHzz9Nq4+X/8hbYKZScRIphIrwUgz44Q0wZsvASlbOiF5Zj6iP
5P0qSUrfP3/+bfEk5qaLhqBXH9yKgfqzmyEKl95ASYbZ65o90v0K/6SBKSX0
l9yhcFo+aPEZfL7lzpERAkl6q1hqyk946fKTzgg2kkQeCImBleVK3Z0jTnGR
zKJRcpy9w+R9ywxTXEBIJZ4jZ3RW63Znyewvi07sJ0WOxGdmNIvcRGfglRdO
Gg7bCzCu5BOsHPSUhW4IRi7ctmKCi8IGvAzQzTL8wn4Hd1qsksAUxWkQyURL
pnEdSMA5ZZXYdIccpYK1w6ndNSIvdrjeLOZ7k7Lx/jhfwhYwbQgswEHjdYjy
44sbwMFeGaenbfBBYoz38zQ2Wke7gm2CwDuX89+pnFLZEuzk3ecXSzMGiz5c
AWeX7pUTZp4JDgvBpaTvA4hDxS1ZZvcw13mBTC4c4AkfmylAuWUulDaTnLuq
dvoS4ffcFKpwtfsUIm/PicLUcEgNJ+ZTuh65ZjiWKE+199iHwvUWJlmRasP2
8jGTJ85+D5UPNSjD0DWIu1SNU3CYJS2wIrFq+CPMTd8qdERWM0QMxc2JrTrd
UCOWDHluY034JKvPYWfxa4JI9AX51vuzH/GKxyw2z0qEwjEvocWApAKsZSiP
yJJcHgjCvZTlYjqnghYF22EF2etZ+HmHLx4AqAGB1eqz/7v34xr7FU1FOhcC
eHqRbVCwJn3ItPoA8hBbKAtipGcYAF1Q71XAkkpNPR/d/sTCUBudCQTOZvF6
8VSR7HLK8SI0HW9v2PpgPHMhYhgIiGuGBXyJ227TgyCSEnQti7fE+HPtIW88
nNNi4zK2VXpRCMMMGKtc5UDBNaRKSwavRU/VnljE7p8SZVXV01bK5BmBponU
SfJCvnsL4Gqdla4NYjEBANWoMKhfAusZLoRbK4EUgMakgzY14g1aoNc3qh0J
CwgJV9PxVsr7NFvF0II7tbQjEfUDKNwgV40tn51mqYbR4/oXkee+zduuj4SF
BrcMVkxKDvMKWwBsYZE/pNa7O7x23pP2i5czCJqC0/RqbhY8dvkWIJ6XE2vN
POc9pNkIyEIkh+HohtghXbPk8gNoPkx+zsyUHZUT14D3Obzv/ytnralVCCRP
VJTEh+Bl96vBEsAoxWCUzqxu0exOSoWqwL0GlV0zypjmK2Gkx6KF6F9ElRRZ
f7h0Jc8HPaUuwkazHcnaAegQHX4bxgWRZlrKy//FQhnEhKSyl54igYdoR1/d
ysQdkvfZaKuW2llN4WSJbaT1FT782U+Q4jplaTDz8GmOXqfhcT4inU0Z+WOH
R3EKsw/0CaDF8ojpDYuS5PI5V0oMuyp/O1f6rLza4GfdAbk8EaJlb5uoqinz
vQ+8FLFqqDCBkNkLk6oNFNTsv4smztZZBgYguMqz+e43+4PjDzerx5z3Bkk4
GlMgKLoMeSkfysDFhU6AWqh2tNSzyQYg1wZAJisXMLWnTfxpFx03seE1GS7g
qJKkvmS6JFvyBBCiC201+VrCzGaKfAixiDay4y3ZVoWaRfwA6QiqSZT4nNw+
IMHd3a2JR36Orlp57gNv9jgBBQxE3hDUhXB8hxF7dWpEf9u97UdGykjI03CB
7FZvih4pKstJq0mjV/Ay+9oFWUEE/nH5SA3DLkMlqCso/sodbEQorRni8uOR
3aMhdz3VwizvazI97zSaMiKj1QvVffXDGLOObZiKEMjzGbL7GpOC/BjhfZTg
rVEzyL5YK6L5rkLXAq6EL3rh/GlS25gVW6bqw2e8yqezRYinIRdepxld8gue
CMSq8++RTLJqmfZ9KWvn3Rjdr/sfGsO59r8K2YwB/I6YMi2oE058zconekNS
QeIUHi54Sa+pT2vCdKsnVHQRzaPE7TKycyJ7eWoOgciebnV1+0j+0LHLYBTQ
HXEWB/qNZBbP5vrIIOde9e0bwG0yvpuFErU+2IduBa0Z2vKCyrqKLIdNdRsc
Utkk/odvyAglcbkMhARU8tMs0O9rFXghShepLxUTMazgFWhMO/HnSRbpOcLo
bdT6fRZk64QY1m3lTymP51pEAwLWF12+GTdnOvaNaniPf0n+NaHRcmWdCCRT
yCCHMaRTwRVAPJooLBb5XnB4PjBmJfO9dz0Xls15vVjS87ltdocV1hHnKsSN
XKb2uly0HJdTIjJ6BK8UtHKquPjAeRETNq78I5fGnMXJ2/Du2pig2FZDOmJh
RrexvwtkNQKzlGJcSRFEVdNsXAQx62/zVJX4vX2UjgTtHPEfo6pXseNOuXcJ
VtUUdJdnXqfm2Q20suKZcBkcuetNxuJd1zIyxanlVvCeFEx/i0hfIfNREZWS
Wt45+cVWQ3RA5Jq1R62VtSbmX7Hz9e1ReCn28BOANmTdOdcJsbyFZxkiLyo/
ypDgF5WjN5fxMRc3DxLJJyaBUkZBJfeEvP6JB086Q2jk2ZkJYDstfZxV2XxB
hH+S8oQFbiAm7vOcsVMkqILA1pqgNPm/Cxstgc6FHAqi4H1A+4JKiGwquZgw
R/r6vRzEpmEn4UxlzFflsjmuqAtdFS7rNjb7M0Gvrg4UCYJOFgRkjtkbHS8A
IqHq5aoxnF6p9llUxbfSnBJ0JQWErkerN7dyuBJhlWqCGjt7cHpx6eZ9XRl7
hi8tlDkf7Bvu23pKcIWAygVAs4IoOPtlntfcBwgUcCKVt5GArMtHG2BIoyQC
EsME5CHjfaI1uDxtMONQCPoQBEWE6/fofFXE2l9zXl3oaF+J3D0DDG0Xrxe6
oswDvdNhWx9uMEDRtWcHNpbEtn89LK4RfJFUV1UI0VouCqCe+Mhn7rh9Tplq
RDmfYHZsVvwI51qc0i1Q+V2LOdtgYqs4iS5ADwmOUfaAy02hSwb6eM6FDKAd
GkYC83blfG8CMJBmq/YmviFW6M55yo7XQChK3QGp74rY4Dr/Yh+vK8h7N45a
ygFDfQsD/sJ+CFgO9vNNuM98eEMtdE6IPj4BhTGIs7py5nsx83a+AWeW196b
anabB3FkE6GiC50BbMuo+FJ8KR/Y58X0JPuBSKQ5dJQVgsmeY8OmSP90u9ar
6K5ukdP7FUPb/yd6UXep4WY0d3eL9yh3B7LTiB2PTOJQblQ+R8IEdRLuAAOt
6WBv2nZtrGrPL92ikzGeoPgLuXqUABY5D3S+QiZg6+LW1Vc8xLpmpBy3UW39
gna+bzWtSkXPJxgxJqLakW9EGBvbfvcVC7L8iatUEXKh+mkUCFSTMcOTRdRA
lE1QlONbbQGL+W4c4z1N0P+rrrZoF+Khr4yTuId84ld8zy7JKZcHFQIiUXL4
un5sA3xpQMHH0sowXhM86hFqvy9MD2PtiVhWJxcv9cnoQi+i9Rzc0pRaRR2Z
fKPzy0nNE/kMq28Wz5OPhK2XoU0yDZuUFjrRvbOPk07hhwDLu8UQtwoCPD4x
dMLJoqUw6QzLnLiYGjXoGHKhnI9BFQCOnYWoZOhGrOofWcD1/JSV6MuVYarp
lE19GHvkXyk/D2Ar6xPiz6w1+KIudihWuyD60YVb/h02C4kX8aCCOen3EG4h
KaXY3oEVGvs7ammPkzk5imP2PUiLFoJQz4Zk0V+qHZzrXfXidMTI2CWgAE5w
xKW8SZGugGqRXpjx7SV1gxWpIp2N5Ld10jaXtAt3D1wW1KoHtzIbS2vm9M4f
I0LXiEbd8LM/IjllnCkjT0lxFOwm9Sr2WRCbnLYSkw8JUBjhmGg9Nf1b0ITv
Zxy3SzcsD91kCwZoaq/w1mrG26N/j9hjT1oWDe+5yIh3DPAYg8PUi2JbUIaf
m3iiHHEANosswlHV8QrOrKIHEU9Txry3dbC5zR9yR31JQf19Kn4JltdjuOGm
IBkPq7Iwpw8QUC2njnJhBjqJC6dmNOdAzIjajPYbV+oI497Qiw3UXPL/oPMs
E5RUVKiFXUZxsawCS9a0sanayXXuLoOJLxRiDutfxIZk5WZoF5NKisddEbsZ
XQVpsymWrUJoi4Slly3OqHL2EzoEu6GAxUb0vNaNbu10MP8aPLc+jwF3E+GS
Y65ritKOEvgIffldWa3+tb20ZUNAkl7SxZgEYbQe+AAWUjewt+pJSxBJL1/o
4vp9LZmncP0xApRIW0LQep5fQ+tGHhALbqsvx3w9z82DvZ5RD5jYJ5+2/5qg
/jqJCD2079P9Xm3XOdAs3CzvyVSAcdtAcONiL6kBzAudO5ht1A98rnPpnSKj
xEXtIGKvl5iEX1kfhYm+g8JzYw4m3o1rmwajf+dRhM44cjrUrMRmn8GEPt/K
28s9QcOQR/1Q4Z5ktsWFGoeNtzS1Un56fEDyxYIlN8MPkZTiXchp3ZjfofUF
plBbAWUXWGFFeuIHAX1mYB4Ca2vY16m6zd1j1tnPyX7MLWabwIr18LLfEWqb
Qznmzy9V7trBJ63cwhAt8W7h0tGlA1bpTotGWCPWlPVbM10VGWcExy/KU0YV
heBSCIi+uFTZzVYjVeq0Hj1+RwlFPkx/3/0JAYSsLdB2M6SGOeV7AKgohjwR
Rj+Hpbi1m7zdS86RxPGtRzICI+HNQeVJuFuyrSHysGLKDuttPTFtwlpBREkG
RQiQSkGszsV11ky39TI2SPXYD4zdSDh+EjHTxCMZkp6oFtDXPj2Op0CHBTnT
wuTDgE2bPxj+E2nwzozhjbZCK3b/kfFr7avd9D0/kMB2i6LWCyjPMmFnG58O
13qSTxN7w6EnexzpbvNl5nS3gs5Z+VLXchUQU9YTXL1YQ4hhwxstvj9Q3V97
X9YrZIUVrenDnV2z9mjiI+xWL/OGjy5jS0XOPsPGsgoCLFcx5jFzfbRtp82+
Be1iTOYGeuPsMHojvQKeUG74a+NkVOj+EkBniG8s6YhTbHpB/GszIHK8VLJO
gJxyXraB/FMR/R9gFRZ6kgRvkDfy/j1LOfcaQAzUMrw9JzKWgmk9Zax04CRc
64EJJCnHNSJmOS1apNRlZEXkoCpRJCkBsW2r83etbN5H+B97sAv/7L3hBql/
ww8j8qsG9nUxnuS4Zs/7NMiGx5YPHdwrFJlP5nsUByJRXeAmf0PgIFIr4ngV
RMktvvXS4ynLyhRgplrjWAhdQRtcCL/uYtXy/2UjHvcX4GODrFpO8+m3e6k4
IX+l/n3DandD2tA0PyR7p4fM/uD9jrhbpkYzcN0UdGAVjJ66mhB6fCwile35
S9UA3JJc7NbtfLiBbiKFseE124SWQPNBuO2dXyALHIrn34aBUi3Mt/3DItZl
6sMoeroAYQA8xRpeqzn46KGFg7jct89b2jSd1foHDfl4opYZogrHuDKQtwMX
Tp8lka0rDJNkqJCNPK86gQQi9lUie3O8yJ2o4TTeoxbwvpImWatuNn++W84C
BOiB059BfDe2APabC2rAjo0Cq47vlNw0Joh4ga3DHYAphKEy5HAu+RmazPnA
0n89P2OMa42QnPg39cLz8qMDVicbRV46PoJ0UdOYGf3DuPp2f918B87gAkVF
0YbPgkHG2fyynf6APbxOXkVHomUerh3HF8lFuU6V9lxnNTc1daVU4xU1zdU/
eP7OwR7S6VHon2xguXRYbIg0/Vu1lSe9xAzqTbiG0w2QRHiu7jR7ryw2GiQl
PF63LsXGhEagLMSoBpsj4DviZguYxmCESLG4ACZ4nAe89RsP5yi8xkfs1nJx
x+I9qC0AZtlTtsy4FNKfFYr+KaAN/uxAC/HTbcdSXeE2RTvGapugx3FcIK8Y
F8xk6NkDAD4A+SMIxp4znKNcZhVXVDSBG9dqHYWWLQVHEmndUDs6dP9mUmLt
8t44MpQ1n67SYQTrwNI1AVVELga1XfpoJ+0qgwlIKaOi5uaqsXDfHiFWCnyg
sgbqznvct+AhJoggbfRJV5Cv2CsqeNH4IPGELXiisNtXnE3/BM87y58hnSAS
pQhqrNqitYxFj+xUs3dzK+ioZY5uDnFZ92oBcfbCH3t9Yplw2vbsMm9/NkSj
TOWB48kbmouZaZ3Wd3eSt19QttOEHZ7EZuajjFkTGeo3/nER755umlKuVIen
M8dgvIFrd2+sW8o8qgnxbPtIc08tjiihwl7/rVBfumVHAPZyG37peiV1zm9L
E3BV8y0e17Kt5+/edchuK31oAXn0bkvAeUPTD6aSzsnpIri2R0rvaGtc8xWl
1HRV2GUV2d7Kd445EO1PkjVSsD9yJAanUaop7re/43FsbzOypZsRBZSOZvqw
ahduE4D3V+86EFPVbPHd9pAIC1qKnbIdVcQlUcxTn8vATF624FbcJD+n6+L0
ScqXTtWs0ak2Eg1VyK39G0afT68QsaVSW8setbeueBagfo6R16VjsrM3RqT5
eJ8VlbNjjaADrd+GIy8WoGQ+gdV4yPmaFp1XG7McnrzcJoR2XmlF10V3yEY+
HtDVGeEMYfnEgVRBjgNV3Zn/v9Y6UrFHABuNnf8hmHVXLrUKsKhpsp9Tg1GL
b7nqokmt6iosnpBHu8UxqfeqWM4dWewbLE0ZeXIyHJqvQblemhP7kN7zliRE
Pjbu6cWWu2IxHWl41fUTYQX2XYW1C1zL9+8d6faacfgkoVmWgZ4ebTr+IVp8
s3lwLLYERewGhyNnSM8NEuOPXAPrQoZF1BSiMh1Zsnav5dvgGem371HzBbp2
IGQiSTYqf3pRDp/FpjPyLptKA+axnrL/FcLFG3EL5xNUJbDes/J3Clsx/NJE
I4wHZLylZiLAzgC3zZaahjww88OMnqDE4MnIm2pEf6iQWgIcPPu6aiFi5qlX
d7wYhy1xLoirZX4BjpemjZGV3lT1RCIp9RgzGEpe+2BpBmnp/JMHV3br7JeG
j7pviSL/qGZGSscqrVHbkKJmFHKj5HYa+JnEgAQnjHV2o+rITrEXX6TO/J1E
phMCmAAC47vkogZ0x5H4mvCQ8O6Z60sGT8Jkml4gC4Uv6bxmJlWazWctCrJb
6k8ZBT5rRodm1InN8gObVDz4GnHPlP3wgf4SWi6rVqdQn964hn0IcWvbmL1p
0JtikWVdnCU6YJ69B1f+EPrvNruhw61/wPokzwZXQ5dxfzTkgpytOrTbr8m4
kcVA9K6+/rE1wVEMAS63WtnuqdeItSCaL1+f3+QUdTtXaNEheWH727NpiIuM
Naq6H8jzDdZqjvPWXKoB8Yr/cxWm9LFvIJzeqMzqToLH7fdfxqzLpdQGN6xY
tVCHhMZsXcxWyJ4LobJR/mFDm5vPIEOEsoOXKGtHUIbxoQ7AmyTlSaD156im
LW9LQRFjYnK+B+3YLsZ0c7nJ6mNWluSrbdhC7Er5vq1MFwb/Y7GdhDOguYVR
DAimou5iAuPZDUHtcNcRMASJaaXgwTLvao8Qcs36xsp0gHUG6nzl00ICy2WQ
xkvyqqoGDKMcdEDLNN2iDazalG7eIcVFCzZYPoBGO1O08Uwb8rjcVLqzHdpN
D3kPnDw47bRoJzqYvURW86KkhSEbKa7ESajKYB4WA/dt2JfmlP/uEM4yQBrN
WZcE0eYtQ/WfqKkzbU115P9dHmeFpH6LKX4RX+TtAbNn0SPClzJUvNNYXB+2
7QAR85eXlhdTCCY4rarPTe0Uf16AD4Q0dbWeZ1XTeh+3JcLiEaxuM9wInLqU
Iln48+ISpIqxWl8M9CilsDNGHrdi+XGr4vxsipyGcn8IdnbHB1hWpjkH67lk
x2qc0KOQ0u6wNGXgANtqohoaWvKdFepGLDswSj1xp1bM+qRaNuavPf0Fzm6H
T01OL0MQ2Aj3QMsuRi4w/mA/FvAzosS2oBXcxZYsVh8Qcyavhqa0D/pEb/5S
vjL7108YGqBX1g4hxZz+toAGUUg8pDTnAp4Y/ItymWT+WiIVw793XEvYa0jd
0mKlPZP+cZoWnBdBI6D6wAEWV9Ltf/T8gBCRJbtJ7aOk2nJ8rBkSLaoNP4W2
xGqfKYBEdkIVSrKuklx9OOx0uSYqO7SdbCXcdTF3oPSr9EVe5w6wW3Gs1rf5
8vPCf+/qsMbytnqHM46MAxgE2PQOJPVbo+YLk0QRmZUM6vZLr1Gfu2XXcAUN
9VhKNDqbChGQpcL9OYCAEYpm4HH7SaLYuLSyezoKlnFS3N+1XKRJnUMbsMNC
Y7aWDR3XjsUTB5LrywX1SlKx6nMIbtilaCN2f1cuKmK/pDAD5v85qybpzV8s
RZDCQHfywrq9jiO+ReUdnUWmuDi/XsAuFCwRM0ZEYOo2HhjGdepvS8nZgfuq
N5cZCJ6ZAOitStwlcqQn+0/Ubc1Ze+8Max6TQGUNFUCFdU2u3PDu2Xpx8NVT
FYC1HRQ1yc5A3dMmwaXPpmI9GRc98dfl8JFRAy/JdjwExqwzwlbVF37Dx4mf
x/Z/Cbf1KBh5WxijBTZgllb+088UM1BuVlsk9pvSBza+tocnP86vJwNbnxWe
JTKW0yL7qrOH3pAFghbdydOvimOHh9UpRIx7e3A9PL0e/6HtJW3j/FKArSek
7RJrELDLbzrenIFJcPxCH6GdMsW8CFzrE9VEAU07c+ly9Q/Eew7lqRrvENNo
gDi9vk9W1VuNJsu0sRB8V/h/bQ953/tjMZZrR1alneCZi7ZdaNC0e8elavoS
IGFxVEbp4TvIqx4GFOPnjg/hHFhbZqvvmrzRCyErglnmibqm3eEyEvhcUl8f
OfSPoolFo5kJNzUf0jCU6gDM/RINRVhnz0rggYRiVDMhKejb9xxeUOa5kScp
kzhKpb/YTlcbLigRNVUidBAoAa4cp+FhozDyjvNFuvIMGEM+UMJFxNY/daTh
68ZM5lRAo7tGdx3u6o49qdap5LWAoZdsSIDJkLYgiow5CUwx+yboJHMiDrVu
o9hcHbiaLyTS+6cy6HGeNWHvOKRday+QylxjM6WBVlct4eRZyNCELLMH32AS
eUJ8+WSPuIHFgFW5zwITeo2/0BRu/YLJRSenlw78nQJun12e90R+lgj5AEK2
ZZSnOdMP+VUnBn2J8R8kHHTphpgUxtUBl3xKOebG+ukhTG/AQTYPNNmvgf32
c2geobrcq97PIf84GFkFLb7Bi5Z6mjQA3xQmKrCJkSxvGe7SuNY0hJwsBM6Y
qr3miYrnf7jii01fUbx8tFMEtcHFD9U8Ld0GOu6f71bbuPJM98MmjrBShIpI
xs/wAHiXS+oJz6AvWr+SFSUwS2yyCQao3suzj5HinsvIjfBv29JkhgPUGdHu
G7Ta3dnhOs+/EHc/65clZCLl3Ehjg+uSrHMLV5byIW8NNnbH9nfR398NRM0O
HG4qyyyu+4NmZJiYDpywI8VpMyXI8vpBWMLNeNkRNfVmM9t3g2glBepXxcHd
WRg5YR8F2wzXYZYEumXK3aA+gH4lBDFIpw7A2Pw3zMhmS+gSjn6uAX86pX4H
vL04VZGsHfJoNhZgtvAWyVr2VvKX5lfSR0Q6M2vicFx39NQkyFFec/TFC5Zv
qhGCe8rLUnUdeaNPNfNnDfe7/pJ2r8Rjsu5tfuXy7Edgzq/vQyfAL+SlchSX
oarasI/AUOiNxJ0fMrFs1BbmN0Mo/MY/sAMh7gtw9UzCXYTD5KokPnq7UhmA
xQODqHMui73NcbbnWke0e68obbaNdL/xpCHYgQtOh7CJvUVK1Ego1FZPdv30
oA+N0WjNfsov3cu5VBiBh1bAhCfhVBSfK3sRxOvXKOZmRVFkeEeBa648RXRq
ebL9eg9I3Zjf2XMTO9w0d526YL6w25ja58iecdQoRT8Ct6z2EbiBrEic+Dhg
OzD8AQvmo4oEgXHqy7NHSsvluR5NXZnsSCpfQ90DJL+FVngBIcPNmnb+yALe
1sU0ySJ77oANjVWum47AP1ieEo1GxyppYsMW7FgmJy9E1/5vDv9XjcFB5fIg
pW/91W6f8wRPppdvQOFnSbT/pScKwMLVe8+bnOBDBh/Fl0ErmgNWw+eC1eS1
nxXRpzyVPKeABCE4Yp6Zn4I34eZ05805c2DMMP6mxtNbGWGZqwIE/wEwfYlN
YXOXiwb2Q5E+Yo98p8LdCAbN3yj+3AWqZWvdjsRnhRvo8ZbC4voGNhVnRXZ9
Q8nZtpysDYxJuqaqX5FznWMpROMpgYXUlptC/5DhrUCSDijCfQEIsZuUmg2c
CBDrkDUyVdjKv0tOiimgUlfMmqN06hgGpssGOrlN4b1ZWe6ycrhlW3lijDhM
ouCavB+JJQWoo9pCmMweF0ZaOm4nWcGe9abprDbp3UB46OoziWSpZr5BXw3E
4HLrLQ+t65Ff4j5Jd2dieGnA7msMRNI2b5BvMx8kHB/SLX/DRomiOo2e2opD
OqEd1r+Z1sfCTmf+DU0Cf/4uWGVhynupxlSOeTZduKVCgVM8/WKI9ZuuL3qx
I71slkeYcVCZQzJp26a8xpCsl9uMSJlnyIFwqX1ED+1lkG2jIKIxbNNL1qrf
/vT7g024it2Ayr4htAJoxu3y+hDK6zKVGxSoyZ5vq67C9IVwL0w/ssEWVk45
YMI3HPJymSGelu+GTZSp8mjMdWgHWdzO+YEEkYbRBtz9NpFcwYv3XAoq1lbT
ckA0a8wn+l/0Ho9MYM5GOY/mQNFUawOBuP2ugqh4XfNIgQQEORNx9v/TpY5W
MC/XXHK3v59mtVXW+igHft9195Vgezq3TT9INmMfXhoWsgXgp/avDiVmWuU5
+fhlXy3pdtzi2b5WUWJjAs68TaO2SQP1tzE+clb+dw4SUKzAYtQZs19maTDu
PGLOtSTbzKl6i0nGdotatdQR7CoxVZw3KYckoaLArSjY2AQleja5hH2sg+a1
nzBIc8WEv57S7fP0tLVMSWgamHS2aqAX8F2u84iW/AiqrFok8E0iIg72RaBt
qzOiFSjklQBaNpVC+PEwudN8f+zRExsaMwYAegpHpDVKDBYyzjLgrbl3oQcd
0tTud+83E8RUNxUFmQLMfbx6tdhGXEzgNFV0Adjp1uJH1f+2FJvrc1OeXnEa
R1oiYkFsb2yJ+PlsqLw+2Oc6oTgI/9Mfzfa9r6FV8XE9d4qVzu5z1eN5IvRj
lJGcPicynBlbnwCE3jJCFhS8j60I0+RsFLyBKN1w1t+FyhvmV1P7MF54rN3a
G1hG5sB0xgVdMOb+fOdmgGI74SDavYQoGuXTODgA4cRh/FG20AzvRWSQyWtH
KwS9THzWl877WdmPjH3ELXFnS1JFpLqKfW8v0J6hZa9DtjB3DJkUEFMiLdGm
bcW8x39nmxBSmfbX3IpgwyApKbrIpSJ7LG4CABqXo+Z5DZU+xBd2B6AV5Yib
yK9Fao40UgM6i3gkRCqP/u3twUVNE++JuIOwhfQrjh4wqEhuM9huazKvG//l
mSURq8eWsdSLMDyV1DH5uRM2hskkU6M/+byAa36Q3+IjGPgCgSkUW+9GWaes
qZJHVoKS8qPChx2fDyy1oisoAw2Q1H3JJSA1FEKvOP+So0WhDzGgGWV74Kig
xUPmhWbJrFaiK7IVH2h2czM1Cj+Q+s+gzFyr+1XKwk54cKgI/HBFn+UmGZGU
S1Bl9xAMsyYpp9h3DM9/PhheQxRSYA6as8IFdCscUfX1ZsxQd/RIy88002R/
A+jWeYa/fcaNLppfh3xUzJYsN6Twk2axztUkos+SAgORtb9RTZDyEm52tBEu
awvJdTiva1irOgN7TpmGFSxkj0Ouw3rGHJgbv2m8CEGMG6iSS6ADlQv6too7
NQovBKW2lpQfwTawdbj8bGRsw126RDrhoj6OATwoeQeorJ4K6ln7Z7ZqMj09
fdwFSnmOF57nuNEVI3H2FmhGW9HpeSkwGMKMP+ss0lN2EADroHqbjwjwRy4N
kKvsC+rNFEJ08SyS9/MbZrLbZ/u4ymXT2f8/QGE4hGeq5hRx6QxYcxjIFeVq
vseWb1swSS2Fu5lQoAYJhU4WxpXt32mtw/FgnG/Tl6aPQaB/vsEMocc/68fS
gms5M3T8BzbBFUXcHL/uyyDNEvPVjcTwDBVvXpTMBoXBJ4pS+lDubT2Vohqb
6H0G6wakfSUiN2MSBLhLWkILk8lQeqGrmxfKDnsSQTezg9n3wfxPkrsfy/oR
KDYj8aqzVYV97099hmnjkPfJsKieYVSCe4J7igxzN7OSibvSzZwFrP4Ndw3M
lZ2P8e7qK5RUGjbqEdYdQ9QgjFG8jMHycII/6VwKTP3EZGUeEjlm+mNLwtaC
+KyWuS4Iq3xIrsLHzjBOJ0+GHQnXYcmSlI0R4oztQ8hnGURiKxExzaYDV1xc
fBorfeP7pmZ/PGI+AJJg6z4Yn0YYQbh7YQll3DhHswfucXX2nHUfsOw62ZiD
zspm3drDbcbOksmzYGP0vyD4NsyDQPrW+bcqPLFdehzs+iRUvU5Osg1M2W/l
UqPqOFiDAOX+wOfBoxukqzUK9cQR53IogQvCT7oA6nFTo34c9inijTirSbMg
L2d6Z477pKa1BM7ANRfS4KMAznUPCA0Alir3LPyfwg6D1is9Ec2YtrsFh6nv
7aopoaeubYG1TaICcJQ488X1HNoCj+6vtt+Kk17i1CVyaHElUKubrm2ifm81
x+SW20V2wYWKsyinoeZLmB2Y3DU0dTMNlxlMOTtJ25r6P0nC9Cq12B1i0BX6
443blL8Zrz22pn33JFjGliKVOWqYGQ5p/Y+NQVrNNR40VgZCIsRtlP+d5au1
nYTslDO4tqEGJiu4jsIIRALpDBQ5/sb6qtCVhBnaSVVGpSi3kn7yyxCMcRd5
wZIlzghJoDwY3/VPq2iWYEL8QPAKTZ+oqafCvOrnCGJ80BcoR3CZyWt8B9O1
nZsTOzHpCraAM3mz3mMVTbdXc8SwomH6vBwzjlIrYzyEYzAfGI4e96nAt6GT
Nscfh0XPNBOyTwTzkJiAEG8uujaXdvDYNc3g0xTEcIyowNG5cJdDC0m+/mtd
6ARc76jD1LwfpfGDBvJ8w7E5EtqGCtRI/qGJNA59vxqPO1nS/I0aPh889hcz
o6wfvQCygVH6nOUmdG3WpzCk0+n6i6vZ8D+c22u0s5gtf7MZBajXb+eyPOQR
xZ4Sv9riEXwAPpH+kKY/+uJVouRRk3m1FGmCU8vz8laNkOHkcpVvLAYU9YLY
4hsO+9tu/f0t9gvYBSbpxU+PNT4eUf8whBf1tfCOvzSxh3jrh79dqOYgxofb
S2Dv+DJc7i7XFTIM7npLc7ECeUFOxymAaTtSe0wyNkyK9bSa8zIohK3DqWI+
1Fl096y3p3JroLyM1AmEoSa5VRfMZuiGDKCYHC6GaFLP7D/0sIH81SrmkBZ/
INrrqTFiwPPQkg4mWXj4AVda+rmQDhKp9o9VSKANMizsTSAsVpd/xQbVsuKK
nSyKIlP1ZccoUttmvApj+tv4j36f9rVamMfHeKozF+AJ+u19gc/IJT/aUyaN
nhwlggRkSJ2tDozX7Cn0tkFYXgwIHNApgAOrmWiHHLIX9O33UNhCL/QcQRLB
RkkuwCVkCWszRx5N3pQ032g2UhJXBvL2bUg6fOnNprka8j2SxoGe9YfLQ0/C
YH6/ym7enlemqH2oPVjLl5ACcCsg2mGAvemm/ZTbXbJUsFpEy1JGZPjk03Pb
dHrUzK690whyXbgoSXnUOajThXoFUgWTmatkJtkrZ2Yg9dCQm/Uyrz5F81a/
ITRVsEaVTn+53BjRD6out4JZyaV/YpnsomB1SUs5rOrXrmSnsgC0z73ZRZr2
UmqL/mc3FQt9XKf99+UyPxRf5gOhzHqv453O1/ebBEoff2EZSJ+6yNAVXrF6
skxmEgSkPdTOMYXMH68YPJmvGsryj9d+y03349aK6xf4Vs8tHXAeyY6eCM20
N6AHj9c/RQtk+t203r9yN8etO749gzKscZABuPm5wKjHrToAPP/XeoxPSVDK
MFJmxmZIIoBxe0mC+nzhLK1FgvzLY3d5ypDZpHCRO8ovBPu4Wp8vFjtk8lG8
kpekaErJBK1Wp+Js4JrsCHR/0D4TvdcTPIpneKVRPG/RLggJz6xp3zyrYHL4
lr947XnYRNpsOmfA/Gkt73N9SDDf0CDyr+v0UC9Dz1QDslRCjlUKCoaY1oV2
XzMoJWpXNJF7hkkZFw9EVopw+by7SZLSIdURPyyd7Ou6lnJTGZFJYHjAy/UU
mnUAgoeP5PxZ1lsy0wyGEusGNVJuWiCVn6V/Y4bq6r9kQ8qtWd0Kj0dF/Z0g
S7q9wH3OViPHtb8gqsjY0HNwis0Jw4nAer3TcF5Mofgi4z9cM6te1Tv8+nHw
nIiX/P1vIFCWBFncJ0s/xOI0SC2MMdOwzGFAYUCJVJDKd1LuwLJ2MPf/mpAv
z88JNy9cuRUu65xLf+ikFfHPx1ss/F9/wZ4Y4zW46+6mjaKLJnBUC590Mihf
j5uD9a3GskDS5PlKaK55G5QwXakPuiHubXkE4K31swG5kPfrYjW78eHOUgIU
zbPubI+nldVUuTsU4eHfYrOXdqH4cw7ezgGkfjywRxoakAJyFOzZqTi9yLjK
2AFc57folg2xHF/TESYw8CvGyLrOQd1soSfu+F6dpnTcLlQtkPCrMNIzMIWF
vWFSM3QcGeBILNf7rEyPb1/V4o8R5Rz2KlLlSKo0ux2Rw6/GJkOS0wjRGQeS
Hinwv+IMQsZBoDXQHP/b2a9Y62XcXrkWdPYAHhABsE/ggfAmVr1Clc3qVaBs
il2mFv4p5gaTvwfKcwzUyTGtLI21eHBSQJdqGWgom87XbC2mxDQST8A7oPLE
LedI23keYRIlCnYD5ETLpRx8o9H4867eFcLdGLUus4Z4nBWihEsH+At5vrcD
RsY23E/YfpsvR4XAuFBsRqihJN+MQFtk0xEwmdmAKgl1WuD3n+jM2SAFaLg5
iiR2afTryfz0GYovex3082A1C+Dk+DaZj+iXhHOn2T2pwhVGtiAuDh0nu4PQ
Gc2Wkcb2XMqdsgMvgUMeLLnN+yRY3IAwuZNtgDMEXCWROxk/CksXCTQJiMmd
a04h3je/z8lY74jsjgdIWQa+Xe47ODo2JNld/weH3G2GmL0Iy+S2ndwL1hFH
2PHClghGlN6Opj/9zh97eWEzb2vj3h37zQh26mL+lRgI1u4RSbjUDOs25+mU
cQuIkAp4dWSRa93R9jQTmS+sCOQrGYBhdIH4Yk/z0TrOm3+Q3N4iCidFMwvm
VHDViqetqtEqXb/26TFADfQfbVXw6nRQ6XH6IxejGuxjai/Sejmiym5CrU6Z
oznUlRoe+gPq9WKaylbVQudsU2sGjDx6jrLbTx1DpyJjl4XGquLCHwfJm3MB
zsk9HPOknZxDXgE+GiDAn8x8uQxYDjraryn7B6jHTLP5SIUHU36cRjlHGj3Y
K5ottcx1w+ZIi2DSSbm4XEEUkkhNnDKPBLuig2dnr0ULeTCytoKOuv0JRCZ8
djrBWgcVEKYZuiHnzMeZuGlGJQXIPsBscqQrlXJrG8IujRK2dNMWLEcj1DZP
KJP76NBE+XfYklBrhD3cmypgX+YRgu/UEm8rlqM1glehbxDcrt2aJ2UUsD+J
K6Tk4z0ZTJiZ/Lvxumzz06/ALx8giyPP+YiI79pI9orPmB44dYDe9Z3UWSgt
2KUqAbo7QTftRDY/pb6N/A25U47SVGHOzK9L+9+FUaE9An3HAL6jfxerejh5
iFWdxoKB8IFDDNRSrkKBJiAyAN+yP5ktcRnVjh4hMvP9Hsa4Pnw8wwOMSplJ
tjFKAc4fqdbB0bnhxFNAIo7fXUBSW27yXOyQYhUbdYmR54viVenPwsxW71/w
VnjfdeNsJiQCK4dLvLCi0wydJwcdkOlgH6M/WnYMuLzqiUm3wqIqcs2MgpRD
iZXpgFrZOwUfVIn1jBDT1m6RSUuS6djVGvXzbydrk1XCA1lLv+zODnOR1KtC
zEfkAl6R6HUHC0LioOJIahwdT0bp2r5SovLgMgrxv5BHWm5hH7bmqJ0zIuGw
Or4nWGH9PumxlVEzrPBLJXGhMS5aQm41EulOLzWpumXdgI2bJEnDfXjgvbkn
pUe2gMF0e0PD5YO+eY3mLPacsEeMeBIPX3twYAtYg4OwUrW1akwZUNSjji1G
+HWzwPW3MkYbKMCBk41h85Y9z+RgpFSS33nOI0dDbL/ICf2+vkcIL3nlekye
oN5c7+w9XWtsHgIgzNopjL+R5NgDbMsAHvBnrwyqh163DUmOZ8zZVsm0xVju
VveeFR/aH88tkcj9PZjiiLt47oiQ+hzEdBpzzJdnGocrXk/48Vu0P8Y2YMsh
Q+1Kcmx1vUG+DE0BFCsVSja5w6OYZHUaW7BcdUE0Ojq4pKULpa24K175VE7P
MndmagIOcRqDPStkzRdllO26J9OHW6/IK5q7mAzUIUtpSMSgB+OYVqdxTNXZ
iFLFD/+hQ2N+xzj3V6ly0MA6QDnzXSSmWvOhKruoZumXTLHzP8W4j01Jk1sh
9l+PN0Jh8HVLnkpL0M3dQUrcwlQw388JlsiGVBlbWI87CFRUEoh6JiwXmQMT
WJZCePFSddPYrEsCREDLoX3NZvLJ0+n7dlK6+A3RhfktvWScA5GG7s9WKFUB
20dj2F4gUh1ddrm/M7HMTdvPOQHrQoS6cJ0hGnzijp/nClBfu1uucL1wLgu+
CwypjVaWT3gIvyoWCrcsiDhk+kPnfMGpMeWNwNjGmwhRmdPMHtxZ/IyYBcj+
/PC5E+svYRrhwF2K8jMIrT0ffjf6ijbzVWb/nqfuacqb7HZj/JFe6GaDkAY9
U1o8bXJqFWu+Q9tCiG9La0yRY0EUrDQ+jkLM3jqj8IQa8IS5HsXxazcaE28+
KslSfY+rclj5xawFDwn//jkXPLk58X7Sd0RShQ5795ZphgKVnklWBdlBox7I
ZkvFhDxAyrcSlJa9R3XdgFYp9k7nsnWLPpenU7uhliQXC9aqVs/rO7fAWYJj
nAjfk9bTyFHdtDxM2KtZpBX7b8yvRSmQX9ZLSn+AjBPugwfR+98JImom6q/G
9wrezDDl3V8IuPt/py3uCjarIBj4kNpJjs47uO6TL0fHSqfceWGzkNF6EfoR
XFCBHT2nLlH2ALgPR4DG8JAXWE5bBCaZGDAm3KeroUR1te0SAmXh/7sFH95D
dVIWMQ+gzx7p6PQnOgGuXFY316J1s7Ol4tDlQLfzF0noHKCg8UG5i8CdAeGQ
TZcz1WUN88vaKQIrIhnUByGFLNGcXO9DMyC2G/fasXo4K4qX/skUUhVb9o1t
ma+IROML8vxceC31ZLt8/bbWMahYm+dUMIONeLHAL1IcHYcm8KB88OIVQQKn
JlSrhkGCZye2QbPK3ovfOKf9JMr734WhfaR9B1XgaoZ+dr9Yz0YejtCq4G+0
i+fMPyTrYetaTleBEgiIRXU8fhLsN0dsWDfKQrQ4Kcj/qTjRCRCJabB2yHFZ
sgryR2GcZXG/QHbR6oJzFVuyJxJTmRpbguRSomV0wTvYML/rJpgn+oNODbNt
aehGhiPuG0XnNgAfXWPQ+nLEfw54Iq84ievpZ1vvpv3Cw+Sq2/g2bnPcMlsl
vMFrECrNnwhsHDLhjVAMBANCqMjfJwv67V3F8YyiaC7w4koOf16avqr4Uqr3
2MLLTQ8s1Z6Gn0KhKFDD8qpvk87j6a1QUOwt78TdY4U6/Vr5m9BL2/WsgdTt
rUFOSO9Nt1ASJYACWuU0XVD+mEta4WYsgkPQHQUqOWCL/E7s6WIBemzoymaF
ucB8ZsFDFzLNlNIj45x9Y9L/kCVYFQimgfOZNqlMhz7ok5kriZAP0ZIrwJPM
WRnBr0nuai/g1veTFhPMw5MbuXeOwnhhwBU1y8GNGdj2p8RkCVMVbdqW35Jr
jJLlYuVKWqCTKWCkc4W75QDWCyAvHpjaLcbxVoAXg7mDJMrTOHkzASr8NV2a
XufYuzSNGqK1t1blQH/raHMZ4ElBSui5D+ugQUo/8dY8GVnc8nPgdXtba8uh
eZMP9p1u3hI4mOGm6qY104/h3S8Br2AxlWm9AEIiYRsMj1mk6P7tMM0uxvuF
mf7DqyMokDk5lLtIgY5mnGyflL/A9fXI3oRyeh5bESLKgkc9RS1r2JbV8UiM
Ep72PKu1cSCixLFAt+k15qfy5fkzr3kltnHg0roda2fkQvsjJXH+iz6Ua2nL
DB5Hvnvhvq7sqog/wYF2/25Vi7h7ZMxvS/kJ7/VGkxWYAybtArRGpsXo8Z33
NmnCJvQ8M2jryHT7jAmFta6Eb9FnI/+b3dGKgvxVxU1JpW0vOOMuNdbMFWY2
lkwNExBm8FOzsEXltZM9XG8krpo9p0r87hajC0U4noJrFLIGKnljOwaNbbIy
sKMzBqvkKiAGfMaI/33VUy2hwwNCjsnQBGmiq/cTNzP7UI029krEhz9XgTrm
mCONwEaATWPPkDKj7TbX+LsqbY6PQEWv+ss8AIRL60K+/fBMj1LD5/BrL3Wv
v/4kMWUhHITEis16q0jRt2JE3syBHuoyqin8urDpt3XVEeIB5wpPU8bQnaRl
Y+sKfDP5XkPLMQWuWlnxm9lB77c9/+aU+jh7PifRlnNHZRoUY8hFontjfqsZ
eCaLRnioKKWkUbB4hia0st287kMsPIlGkqvZij+tnpPMoNH6Yzb6N7MGRxLo
Vfokfh1UODfxfxJPMdba1hGcqmbYdWqiTjhyIYT/8R+tPhEeCrZfIZue3TGU
tJq7YdLD95dfqimTnl5cXOeDkSZdvM6ptU8ZsZNkbk3lEIUzEUwBKbxBNH8W
tQCj2jLI9Hgrd4K5yASohtnsuDCvM/dM9Dwh5Roupadi2tYb0IFnzgUSbSNO
U0h9Qvl2fYRUQ0779eg1zwuBzCUwAz7baB8r2b5Yr6CD00nrd6TXfegfDUS4
/X+nEHgt4dIaSPXYPaMor6YwwUOe0fSmxLElQYVKNf4Z1TFlwr316rs8427t
eLWoldKEiysIBfVgQ+laaKNPymxuVhbMqsMmfayx+ff+Jg+ui0uzODlgrQYi
UsUvXvauFYzkmvT/ZcJ6BYF4k1FIIohmsn63z45zloWTJYexqOPqwWV5pbSx
7EFnupWeePuIwT0pFI/eFOP9VnMm+tqY8fIR0Fqjp3sXhLRp+lH/gCWtvjtN
UVzUG2n4tSIpNZzThbUbCR2tJnNYAahdiEz07OJBKs33GlF0IZrPNP3rNtIp
gkk0BdmsefifXxwxiTf+oa5dNwRqvSA+yiGx7KKKn0ihCxoB5ipP4I0VxkWH
Q3EUJ81Wxu4cRMn66gNJhFmHL1CVSgg/jzTYr2uhT8IlnM4ewx2S1xjcclJG
aYb+7hO+v050OVgEXUnj4/W9DA20XwmiObSCidnNxNNXLnUQB6DvJsWUly2j
Q8ZJvlCngQNki/N4/dYrMRpkX1KI6fbQYFdX6su4lCnUl1FuoBvAQLhqaONy
FZqaI0Z298D9RqpeU6YY3x1of8tOY1q+XE0cjv96SWLklnReZomYkPQMirg2
5ZEP2rOJOBDOAl/HwldLNWLLGhC74jsijY7+hNy+0HsapIrm7dYX0yDHUGG4
lEvihjw0y+PoETvwF16OCAbQqGBR6Lfld6jeipwdRALXyEgZj1i5uPpt0187
zqnra0fnz6EbsFsVcdfLhNBGowORkCk/u2YKL9tXCCYhfP+Inpv7KYev2LYt
Aa/uoOlG74pWAYkuvhsOvysUJnA5ZWt+0/A0aEh/23vZBKT5Kphy51iK8JC2
nruqAsiq2h71+qhqGK//hyQ7zroX2F0DVTUo7zZ9xDpRvCY1TCrUu2q5Vod8
GsWwtUBC2g3K0y1F5zD6+4iCAtZNVGSq0Sg1xQP8jRecynLCM+oi4zOlLTIq
wznpT12JO/ojklftUFo68bzbeo05bET2jdde30hDdXO11VVZutSRPsRon60O
M7pUDfHJbogRnI1UC+FSfwRAuefd4qb+CwD9xo53mlq/Xvh9tkWLznCI15Ui
5IaQqc/uiRtDsYiow7msyxjRPVJXvAhckfYrvO4pHvMk284I3Vi0ZIQnLe8s
LB5CvPp00cv46RbksCGS4tlDQ/05CQQFUzLQ9jA0Mh0JXNReR65hZJzoeaN9
YMr3gz4hXT4Eqh1jk2sy6VP8xvMwKwRBQGbQEAUUdAAde9bdVBl96CIPH//C
Aav8LPzzE4CT8YfholoISKFkaGnO4nRqGKpRnIkYiECUD7ynapwjeIPyEe37
16k4SKRFO555+vgAadpco1Q6wqYRxmYgGxXn+cHMYT1jESCAMwE5rQ1F0gF2
2Jma8aTTuvH9hKlZ1EBK1qPfdIh/FIZOtS4PQfNyM1OszpGiGUMMDu6IcQk8
rn92NA3FKp4QFoWENFC50N8SKZxE4EexcsECwG2jAxKqz+sN3iWXBWFl6gdh
6BDrUZWZunZarkEuddbM59Ce2NaXSi+A7vK+DFcyk4JsPz/JNGD2XtCgPx5T
voc53BpgHehgepgHeceuAdUOHocmlSvJiPeru4iJ/cNFb5Tud+d40MTQLCcm
uDL+XLkXNIIBT+KIVDnUcl2Y04qcty74EFMmcSF1sXiCSTZ5FD9CYSL8oxb2
Ttko0Uzq9sXBrgszoqwZHSIPS9wsFPn8Ki76zV+yv4RJhmXmnHQ4Cag5oqwM
IAQm9ebKEGiugVFds0+CkbLkSM7UqOPc2s4fugKZPUN8HBz0poGBXjVjUs92
6tCTzbAHf5wQzZndBI8WRrcx3KIStbtubY4ZWxgqPHwdHNrdIgD69IVObYQo
LCFwiYV2wJeTfCiigesgRISMiQF0aMB6avv/pSgs9D0CIubqSKsIDmpznty3
05iEZz0PIBsS1vF7xox/VjjPA1zqyd/GCl0YToTBqYtREOsMiRcpW8qTEg8k
pcJbzqdW36tzOGQCSoudE9QybSMSiPRfOQWb8WybH1RWvK6BOwuPQpsJzkzo
gaY30mh6trxYNK+v7VuXgSVRvJ3tSHKao2zjS+JfMH66aehQ3lfhDG/O7ne8
EWzTXQ7Tks2CpCETdO3IWKN6yy2vwTtFRXYGb1StbgKAPpOLYKp1KI7ajol2
k6KTInAIbG9gfdiMn+031gVrB5FU6PNJvrxig/ZyVVHT8MWjMsubIxB+ypKl
62alO9vThXqVWlToh5sRsFj/oHQj6K09gsmDSypTVvqMHBqYy7jiwGYP3q3d
Im36r7uNPrsN9CAVreC9Moq5zNvfv2lmYIW1x+ledna65RLHj/3mEYmBve3s
xc7DksY8KTht4d+5PTnlDU+IZYAhvAxMlI0dzpvTmF7JUGlvH315JOB21W6r
c/DpDtLiP0HlwCWSXX9NGZQRBoIzsk6moGgpod1bL8MKzs5w+2LkTKOgc49L
4rsxaFOF8ckztpSJum2W9x1ruptEfXtns4rCBxZCodV9nxhICDEaITULjEzB
1TgAQYEKGki1CE/nFd0acAQtZa3T1I913dWfXhHIz9O7G8wHQs0T2jjE5hJT
nrhmpZ/nR/Kkiq++svtXsfyTeSNA7eOCoxQLJSFzkWdm6225MJvvxJhGpA5y
f2SwL7TNPDx2AuuihvCKZQFxEIR7JUNQ1MMlD70wAxNXUAfEbZtnyjsnpSnp
1ISA0c+wYDCDPkSfYP3W/dqKtJ2fHoZxFx0VjiyNT7m+oO1psM2U6j+y1hRA
9Zg9mQ2c/hIxsa28d1nnA66S7KzFzowfx9raMDB+ry56/Tt+/1kiCe8dUj3K
SbFPppPvZtXVsHwuMm7asWNhycui8wSCkjf4dw1RWP1q6Jh1sXIiHYpVNmFl
iL3EYtBESxlzy9TNsa3+HojES6JpUskEncvzeGX2mY5yCPMz2OjIZp9xLT5b
jQ7v0XFKSqmi0sljCxRw+yfKUtT4CZzbimwXt5If0R2VXoT3O7ZRHLRmViWB
uIRpBeziM4QSU7StN2g2zWmJ2JX18qZi1QYoObPPWUwVNvDhVUz3ofd0hXqF
ngdjQwXvLvgppMI91xhi+29gw+cXV/RCsqs+z+oHw6/mHlQ+ElPKX8+UCigz
YTXyz/Uf+YwfRtqt5uvx2VqeiaX+xhK/nAcZ6bE4VgK+5HPn4sJ2zzM67QfA
1WAP0yV302Nf3CvkypliS+TpJgtL5ZLrJmZZvao0a/MDVJENIRfcEVMG1gtZ
QxGmjIYd/S0cdtH63kz06bBTDcNxipopf93pu/uz4KRWfOzpZsH4hnH1xUbt
dYEIUnaUw2OxBkl6GpGCBebFDaWzSIFlURzEmI6N8Su8HABaipDy+cw5lgIQ
re5MHOkSRkXNZPS/AVBqF/7v/nS12tF46dUSix//vEU0dH6UcZmgObuK78Zf
s4NYXTeKYvvaC2LCa1gpnd5DUxu+CSUOoZC3+SU7Nb69/vdmOFJ8bjHelS1y
HOv0Kh/Xz+Nc+SaCajMQow3Y4dZGmhv6rCHr4cAEHiLgRHRCpA2cKG+ud6JR
kRoI+DrwP35SOxb0yjmID8woX+HujP1at8DVKP9qbbzm4u1to2QtY0+G5gQ7
yEnF8PemiTTf+z07tw9VqsF+ltB1EZmzs/QTRxUbwQ/Fc0Dpjwg+2XCmkUy9
TRKj8Ca6c/214pR2HreVi0Lf9LytOL27vNUL0jR/vuRTu9NEQy+x/KaWprUH
yAewqMZLZXE33NXykWO5pfMdkvYgy0oqAoUnSO3hRYWoC63JvH1gOy/A4h2t
TqdGp/uKi/UTlGJOvs0Qlq+CkBn5iFPWG5NnzyAL1uIqZUhVcM0I4zKZiAlr
ikGp908U/itf/BA1Sf9abmeAk6pd29vF2Lf9kM9+tgBktTOICd4DF0uFLx+X
o2CfNLu7ECGWSfuIFEIC1MqUSkrG8nTujWpETj9X46+53PgNKHCxL9t0N6l0
GUaNNgjBpOFU8eAg9EKb0WlYuzqng2CqPNhH/6ntSar+my/G47oXhaqYRNEs
Ccx09isUHnZrQ9H+vyd4czTpojjPfTvSsXGtFe5xT6hXXurZw2Jl8e//yHx5
gLGIi9R9D+GnH5FF13A+asJtcJXU3gVQfTrrcrhxX02l95NZ8iPE701JOC4S
X28hfweUZUVtiyiC9HxPNksxIyTaI3Bqh92zEgW0YXL/WwRJJiRonQeL8rIT
/ZRuETe/xIbMf7INrbYCErL6Piy9MQVyk0II3vCYDwdM+vcS5t0yQt/NjOee
doNRN9nclzkrSExVg+0Qffdy/U6qrE0/4UnbTxdH6BwAyeEv5+CPPG9j3xMh
l4qBVCHtR3Q++OcEhS1gTbYC8ZLik2SflA19tOqIbW0dTJaSW0Tn2WcmF7PO
CAUGE44glO2fP4FPJLAGgky/Ev/d276NelVDazasEURM6iGYvCF1W0oAm4iC
nwOtwb0jSK+Zm7TW8Mo7PQXhuA/NPKqHkn/WUxZE6oC7DxtMRqYXFKKWgkli
tBLqZGll4NezALjUHJIiCTVe0OKVya7jRbWAhxTZT/veA1+i4AEfd86ku3H7
McOvjVSciRWissUzBEvvWPqNl0BNR3p17x++YQY82eibuZ7xz+vsd4vAQXSR
BAA6d3gHtRPKeDMLg1D7xcDH9kb3CV2utvHk0q+/gyV6fvPdYEpNeIZug1Sh
ppQtjhJsu0rccqWgd1u8/zvp9+gkRs24/WeYmLJD6WiUrkMcgh+Gf0RLgGU5
XIlgnhycdkYIxfgYILd8Or1yOOL+MftjGxsH034mcLTgtgY4upikXVRQk13c
YkryiU9MgLZZhuADq8WbdxUNSuY5+W7NcFarFVvzRCnpdJExDymBiEFrlcup
B35C5dtlb182wmuBMP7dAjLNQiD5wEQuIH1y4gv0cRiorRRbuIgU1df7vPeq
FFwUllLXQedeaNFG6F8aN0aDWH24B6Snu3di4fQ9vBgBKtPhSO1EAt5760Ps
xoM8FriqiMIdICBjbMSeyZUr+shlmvOW89QSplYqK12tI2NWWBWb2pvQRXbH
A2P5RKz9ZLdiDp+nn5/pFuszJD95LQKqIFuH1jvAOwD5nPAoFkITKBMxEosO
i86MO5DoH5nduSIIfxI8DiinpWl5HHb27u3OYAyfdSHCY3lROVSxX6M8mG6L
TbMsKQqrxlakL7LLT595Mt54yqJukCVxV5wHMzKyjExYERZ5bMOzguSW9jlf
62WvsDQskP2Mh1TiRcAsKP+qtQJFT2uGkOaShTLwLt5cGG9h056QlVD7x5Jz
d/vFYx6u7HrHvKguXyPzuvtrt7VXea+2nzQijmqvgGJlEsNV/gz2I3/e+9fZ
ADYBJj3YFYmaOWUVmptyf+o80rauunnzKbIZOsFsFvGpyCWji+W6KJlIA5lW
0vcE1AMfiwwUiTlCYVHK4HhPXms9KPqC2EeEfs2ZMD3FPfxBPzFc9DwJksun
YQiMqaNASJAPcO5lbk5kI6fpn+w8Ke8NjDqDshu8/PCwRARYh51doiwdeku2
zmVtKhb+zPvMv/Tg7+fG0jXabTMfEHIiwlcmv42cP2GPaq/mgUOZ3GqdYVH5
ADb5FMSIo9F1Yg5bmkUx5hrorK0Ybqdx3oNBam1mgxmVYIyN23Z+npVLIPfM
cfNm0rwDywm4Eb+MmD0uD8bDQFU95RdixNrUkfF+Alo4uIZ1AYmpAscPYXbx
hxNm3nq8Zq05LNvF43HV5SKRGVKdpAVYdUYRmc2GY6LZZ9thgTUjQLHxCumz
Kf6BOXMVBeFEivNLpELpTDkyvfxksi+3Q4msrXsFyZJytNK4SAoGwnvNcHhj
ZxCW3tfXh5HxktB7qqpJiTbWeggokFv2k7FJuU76yHD63vAN/SX4SnIhS4Qx
OjxpVKsrIQc2UN1HzhhJDVRpu84MkxSREtmZmNQ5UlVMQWcKK6xhFjjsFuPW
5eMUIZOASUpBZ4vJY9eqMnR+XiVpXxDCnLDmRkVJwp3RptVcX/CP2IfPUd70
HI3bgXmhzSdFZ/0GHEQYNkhFx9NKU9019ZEQBJUGPW9267Se55fNxV8krXRg
L3CLkIKVPDdFJkOOXCgSgyOwDaUTyDQdSH/dbBZNF14g69MIihdAFxh3VjAL
EDDWHruL8ogKcOajckbZySJQDWKf1ViRJq+ikh2MWUrzZJ9AlEUIg6Wvp+id
DYagyLQkNJkKtp9IVnXUX7RasoqqBN0LKQ2WpsKSiqm53ynj58Xdhb7ptwhs
UEHfCRaInwnAE8u+/An78j218XkjwvvPiztNtjNUix6yTpy8QW2CXRkZ9QWC
20OU2aCqX+Gk1MopFwpfxc7Ccu7iudJDEjXZ715EHMuxKg0YiyjDbEIaC0Ut
L0KJVUBCQ05kei7GeJgo2Z3MyLjydluyj2rR8cxWU7r8Ga5IPQvP4wQ/XU3C
EpVhNEPSlvKNDt8GUw5mD96rptStV6GcCxsBjqAHyQ2qEN9XOCnzM0G+eHE/
OysPZtX6DEEzwSoVa3a/j9/n8cuvtPF0KECyiS6s4z2aBdOP0BGbk5kLzn22
WZmaTj0Irz8DVDxed1tS0rQPcj9l8+KFLBMyxx8k5ZBtzTiApfGqGPHebQ5C
7+3VzU7w1SFdy7wWpUBbkFb9qoE9nnmHxwnCX5AEKalXP5f/hot3YPv/2kHL
oueujB0YNppdH44I8OU4S5u0FUjh8vZW5NpmfbJSOLPiMHTBC714UOvgOmFP
hOSTbweJC5FvMAmCLp33r4ZnYm+Me+XXnXC5ozEBfaLlg5u9u8FtDI8L1P63
NOgtIM24Aeim8D7ZYTNasSea1vVSb9yRB+6r9M+ogKD3UiWDTr8Rx3Wn0pZb
DQT1u9cx+CxfQFgGwuROkN+xD3f5UTzkm74B7FpjZdUQpjKCrH03ez/rpA3f
4lvXn/wHMtoPutlTo+85lmb6Jwx2fAmgspFaRjeGw+XTokI/GBU85WLQqnbJ
0iMNklOW6/q3ZqEb/OpAByW74IK9U80JrySuNrt3rXRTlHD/DlxduVu1kjBf
XlwukibH5CUfLV/K57SPRQwWFdkdlr4xWbo3mujuVY6wnWR8Fmzjl52llrz8
vmmynLu4Ee2rWdd+PNJlwjXrRx6iJ1HtQboXrmKdh4vuhuNGI4dKSI2YndLy
uo5wq6fsZDK1F23wzJk6DVv4qddvcdZjq/4taG7gRYmka9fCBjwZfNULH7p8
LbWBkzJjNHs6qFGV15LdZzmrOCEvQ1pgtVEHRuTo8k1vozeIlYIoLcjbq1h4
Rw0MnC2qmfL8N1g69JmABUdi0F0ONe1W4NLQ/895cz1qjK1SmLmdjUuYEy6r
9gyJJTeXRCnIGO8xDG0rSjomoAUJCRiJAjEF2T4sDC6qA6cBP73pM3Re+eQb
kDumJLTbapecghz6/l6WsFGKkAkDSFkYSXyxQi0AEFkkh4BK/SSNRw9/oM7D
9mYekyeFj3HizwJzJsTfxNh+7suhSX0qQHCTcjKWnqP0vFSHOf/t6m2wyl7p
PpW8Mm4o4Gu0Bm+6yzVazed2JOVjYWn1ECxqlaX5u7pFewmFtT+BcPKXZNUX
yEt6y/N1KGI3u0Tmq+KhLVt7E26F5AUdhkraU7jVSQxzIaIglVYfmnT8gnKj
RZG0PWCd9Gwu8s3Vz3FFU1DmotjLRmQuSbRNqYUSXMmd0dL6pOTckPpV0a3w
obKOnx7Z3pwuvON/ZwgtQbC1SCMpS65g73rSscBilmHF4ZbVYksaQLZSPXpu
ucAJsvYoyIxGWG54EXYamXcHNfk/LHg0EE6h3s3MeU9zZ/q+lTn7/1HdJuRJ
Hwm3AWtMoHrbPURroyIPb94NZaphAaJH6p7rR6JJaWBW076Zla/aANXo88Zx
EJFRZbNhH/0MS1kqC8eaZcgyR9IuRFLvGqbwBNhiCQo4RRGnfI3HqLYh/Ckr
HH7AxQ41txkKqkS6ACdhdudYQyYMOxIa8ReK9ivp9dwGy75IyGho2pSoF5C/
Xob2BuUpGn6DeQiyzSFSMCOthlT9cwKVCaExEy7M01EpUtapLxkDFxjIgPd5
G272OQ4fhXFoHCMiM7Q/PM2XKwmnvpdeYLZHTPE7ws8NqRtQ0eeo+eZbu2ge
M6mhNFluG/T/50TkqJP0i28VOPcoCQFxztmzDufwdE82uZZ7HaOmz7tm3fzW
fFNrn8IPHYS52eeTJRKT7Q4jQYKvNwnS1IS4+UHDWp32QoEepEUENzfN6VAg
lH9S/X/iKD7ygh2uPDa952wdqxjJlTKr+ayh46tN0ntBQCy6NLnoyvjG0ONr
zcQVu3umCWrXuoUhQuzwCzUd2uS2EtVCuHZVY814MM/kf/HGSUsn14IxokGm
SnjoeW8I0jbFDNCqYIpaGgJXFbCBwzr1oy+1+fa7TAEnFAsvSPgdXL2W2m8J
BWCaawEawadg4lEC/LLJV3C0Kz3JSRowsjh9kcg7ur7EoPxvfbrIoxCDsi2I
nPO+E4BvGnQCics0VwCPNZvuTtOScteJUtP3JK0zysH4OLhcxs+TMQif0BUx
koMSQZPRq+SSVZavbfquIkhMo2ThmpCOyrYYVKw7gucw+pAZhXEiNqpNU9Sr
/Q5DPbw+vVRxf38MT8Jv7t+100FIlTHI/CtH3z+YCeYF6Z+xi107hqQG7x1b
GeH11GqfCQyY8eFGjkscjVENrczrV5Z98E2ePn/9JVZ4uqQE/fWnVTjNk3K5
Mnlt0JwhBw+LxMNBroYrJpcQPwK6I68mAxH1CjZXF2bt17aJ5AUEAC9FnIFI
ZOa2wuI3Ixs5PFQcrZHMvMDqmzrdrOiGjEwi/tBD9JEi4Uv+Ph9/8UdBpTL6
dRECWkHY+1RChB91mVHiIWgtqquu9MpIRdCPqJArE7xXf4kNaY0HfgSMzXPD
m2PAYg+yrOaoXyr1hMZRdiUSZlno9oH9ZBUCwmMFcY2SnuS2jSk0IQGDpzLK
nBE8YnZwoI43CrD656/MerHtJ0YzUhQC6EpdXu1Sq0L1zmcPMhGM26fWrucV
ihFw7y/JYWMJvwIw3FLKHbGb3g91h6Br5+CfvaWblh5fxf/8zo9rZIHUzskl
77MJ07Q3Ty9SoFxCIa9Rt2PPsiPxgTq21GG37FZMUZoPeFqY0J1gZmFt91Wk
JH8CpuGTJltMGp+tJ8b8fA95hje6/EMFvNQa5QptJdxZmu9D73nZvSfRWgwy
1ObKJA2Hk3Ztrolj8gn6bQbF5smpC3WpuBnI63Oc+dEZRTdCg7S9UfmUPB7f
Fk5jFQET8OTuNcxIcMn/nHZ4/PCxjBrYSBYfzFS/B0lB76qgFruetGTQ7DLH
62eyu5cvQabsf6ZDNXHhsM3buAzci4UQGnhlQFzvJhsCeLngokiqLv5DYPGD
i1xG+BgIgoPGhfpq/BAT21RvKGtmcSE4AgW9RVLp1OBxXRhLB7urFs8F7C/7
PnkjvO6X2FW+Y0Ch+XHbetEVLylg8aN7doUseFQS7PnVkTLLL1jHvgdSzr6A
xLbYs1eG3zmHpdOE7wSdfw2oYfPHYQkjqEJcD8bLFdPIJ314YTSb7b2898mh
dJfBkMI7ePe0q4SgIGai91ElBO1MBEwwEh+KgKolZY1EBzLCsxzxlzIoAdRU
6zadeJduRrMZN3WMD+AcisKGtCyeET9g9o7dIqAObaGP1tCtRxAG+MrKLBoG
ts3DIaQvbjpe/HoOt7q2JDLHjXaqOiUSl5B18T5dTc2WDFOyvrBlUtFO4Cxw
E5rONFRwRpXrC3xSnUPBeKwoMLfPzrV/MdIroLHQKeHanr3wDKVzfKrrNS07
OUoCVBuwAgZtR81bn/+dwWFhX+7ZdG5d5VaIwr2Rdwbf67PyShd56PZ5bYFM
XNiZKi21Me2JcQZ5qCX6HGQc/tGRxO+mVlQM/zb2s+nSVhQ/i9Zv9OR6L29y
tPtvuCmH0wAFhBdHQ+BWoxYp9UtscVcTACscbm4TLFe8R3jqYjyx3CCPQwK2
MeBe0J3JwjbVYAbFKTH8nGZxNd3ygbnfRSKT0BOGw3iXXajDaB4Sid9/yVVH
U4mWZeC2BYl6HZvEmYTDSe5zwG/yvP9YKJrnBf+L/zWHtjnRObpEkPbVsVBx
md/HiJaO2pdRkVWc28jT7OcjvJ38tU26Wp5cJZ1bZgU7Jpdg7l1ggqIPtq1y
113+BKcF0aB70aVNgbhBL5bNS2yAE+4B5Y7xytdnSSzqt6ZfsMOy3YfR32IV
SnNC9MY1D8oHOekwzvh/4xJV73Xm2e4fnqnIxtCCfsbDXsdJ6WJC2fNXEmuz
OolO2bXR/vSPvmsM4Sg4lQu9n55h48Yb4r/Rn+RNdOoc1nSfApPho478eSm+
/mjXhwjWdfNUGxRcxiXV85s//vLnZqjSS+l2Gau1ZWAZOgcY8/lB9izqpaQ0
VouBz3ez1IBOuq+rMD8AfhOV2WWqinbSa2aODbIeGL2mzj2yM6fJtx6Ord0E
JU7p2cuz/BVXdc3iPb+jpbH0yaHIkXoNjrilBy5rfAfxYKiPF1DFgVHMlwi+
pLu6dGdPEqiysYohHSiZT5TJYaO0sA0jR0AH5FrG0nvYXhNP14cCC4ryIjYU
708rR8ckRa7BKJcuYgzyWQTkjTq6zA0OojI7NflHxXL/JZhxRdot93imz3WW
EBV/hYmJQnB+jFdZdTTfugtQFFMu+EdhMRC65WIqvl1IFHAg/rLDHi8E6nso
1q79yIwGOiRHpJhvvj4DJi+BpAfoDn6joWpCunDKo0o8oZFpR6kAimTtHzIK
lzCFclXaxtL+m/f3WIL0l1TUn308cmWtmXG2IzbR4UK3EHsef2umVqe5fFcn
7qbNcd8BRioXlqpL77tHrQ1mgah0pjh1aoVrtZxaxa5iEp0umHKUQ+U0byqP
JWfE8t3U+3vgUY2T+E91t0iHuLSKqVnWPDtDXfLvHguUR2KNqDVB2G2BEyF7
6Y7yXj8F7hlUlO5HJEK1zk40WQarXiYMGi5nZtSd9hklDhaOBQgYhLxWr+j2
lXRRg83iCBnESR6mdEeCACfyMaKPEOCEYWa/ZFKxcrYBCWJ14R0p9LXISqu1
X9wCD4g+PQZMGC6DYIUVrHdccEueM3m0awVBBFFCR0YUY9FiFYmLJjQLkQf9
WK5KuuArxEwQ5Td2krEKRBn76Hg9GQ0l3HAUd0OsTxSZ3kgWnczU3kdsgS4W
DMDK0R0rGhTPahIc8QOLSqgQbbnSUbrPAkPvlR2nnNQQ6Ubu76Wx4qbHwNi4
Ur7oJigDulypa+cNuOVKly/YtDvCXQKJC0+4a/unw7pxmR+WuGeBgLCojs6Z
EEmOLeJ/MzYCBC8gSYiF0d0dAZsxsGlALWqpSq7NIF4FW+Xt60LRa2sUtd7t
9UbAEYQv65eINn2xPVvMkslTp80O0OVvJh1d/ZCapDJcthwe8QFM3Ft/wWyi
VyI1o9D/E8R1r8xHVytPBRetGbOFYcRpPVm9fQ4koq1kBEg6OmNW1s1pyS+h
MJYww0gfBAVEzFzjLh2CknNs2IasVSesBsXXfyXi2ZalyzMMAfU++2UX+r6A
daBtJCclQ6kPidiGujZ9YNvTvmERXZiUwqEOMzWEt633e6O+Jk3I5nT9eroF
5jhIHdgNkWtfZzqzXvO62tfkupFt0SVm1djrt3GvJtUOFPjqnfu8RvEuZ6Wg
gk/EdMPnhbk019FZMNduPxU3JwUxeyYc+9fePC5aYXtHc3+FXS0xCwotdj9C
amQ1z/iC/0V8Wmw4BkucZgnTq4GLhBcIAGBm/LJYYkT5qScq108OMwJKw7fL
ZWGvtxC4wXxt9QOyvsv8MmGQIBxPxcVcooH+jK1+ZVVMIFxQ4YA+K7pbNLQf
ScBtuHrtApkfPkkiW1Ks8gR51Q1TUPTPnizil+b/ahFIH9+RdgTtQjUmhRsM
XOkqTfRU0VJFk0qVBPXcXE9NImHIWJVmvsTzXX4lHAQ+wd9aFV9i6n88ppd6
CMidiS9DO6fZXsMW9l61NINxiyl8se4PYsBvTXeCHhBxg6AgqMuUIvcJR7Hm
plMy3D2nBpR6FdtJjO3yVq87o7h8kp5Tdg5p7jT32vmtDDdSoMt5hd2iCZQu
HO5sflM9C26hz0a6sjcTIV/Tnzr0sNF7exp9RN07+56RdxyTfBsgy5U0uwyv
RCPvNGQAcUaBT8XEJZKvNi+BtkmcTOY6wlcohkNrEovXQp7aEOiNTvrSRjNi
SYYTcImgf+kcCrYEfBnEwdd8ns+C7Oq09uUraX3qlwLog1TI+4A5FBhn6YCN
qkwB1xUD+C/ym2TLzEpzB88FL2HkWXmsWcMX7PTStJ/nQyTFAPKzHW2ZJZBd
LXZeTWJMUOSPKpsxyVMUMx3uP14l0ePem/7onBiHQxwG8wJ2ZNqscx882tTU
5UeIdqBilkKL1Afisc/GDvygPlraXS9MystqOWpurKsP63Vk6fw11fZRHE3o
P1iuoR4fKj50zDOd2c8UVIpvEea2xVtmv4aPcLTYiubEqRz5dZ6Ku8UCqEcX
oyKavai3GDolZ0ZHYfuW3zpvbii/a/THhG50rqpHFSKgvvDtOz3w9HHzKKH6
s4vkjBhK3fj92r0DYfrhKEqgAJbs9Pn+ou24Y3bRUoUE7PkhKmrqrQAR3Ppl
E0OAq94eouGrsJ3ITj3e+YxmMmUkhR2WWi+HUiAzPceX9g1abz5+sXEuXnoZ
D/zp3a3jOMtteyx4zrS79453biANMu40sDmMnkCf4AxWvujnnbFJ5L1OS9gU
VCLUNIBNmuIwK32TOtbi4XBAxZGXq7zf4frZyQru90JWuG9EoUnN2/U7ejf4
xmcNPaSopZH7TkUbQeJQqyBYoteSE8g7SrDuK2SaiW4lBU8nzFI0d92WRzZF
4nN1B/Wt7IrhFP/ObZRsE+rNNViBwDcpKauV7AhWkgyT9Wvut6mQcbdDH+7M
CseEgdG9sxgaxClHqeqKd6LCvz3y3arF5a1xFhQ4VAxK2ZTWQ0GoTNTi9A/C
qRYEmp4g5ozy3m9H3+rqhpXbi2vW40vhP4ggZPPmv1T1DSqyfxQgxqCOrLMx
XkmEXjwYpTAPS/SoahU6raN5aHbdNf2uAN229cXJEXoZVlsqkq6zirqqeI/e
WeoJG37Llqn6Y/70g+EalVgQblZC6dWl39W4HHHCHGbUF+jwEtHMJOk1NC3T
Rx2JsC6BFhfh38SeZNhxD3zsjbJa8bFlelzdJSjuGyL1z1bWwnDseH+7UJ9d
aXnhoDMUVJK+d5mPa8Mx+S1cdH7pLIa0PvppwBOksvS6kj1+Saek88UjBsCC
BTkFUsaUtORn7HEBUZchVViA17p5U/o2G8jt10sVNY0dqv1ZM8VumefchRTi
6LQXM/m2j7wT3zSDcyzA3uFha04y0u03NO2AQ5AfdeKByfoLOKJbAB7AlsXs
4LEEraUxrjLpBz84cSCC73anVGLD1tnliWXACnFfOMd4jPZTDGBgtMuwo955
upBM+9Ld8QAh8yN9Ei0U+P6h659ILSk8QL0H7PqfLVz+0tGqOlMtq/bJicAo
P7yXawmyUimXkEcHsq5bfdxagOvSidrcSjMPhEju8vsm9R+PFlOmEfKnUz1j
KT2qlwvykjrnr9oeESDPi1QbJrK7JNBTAgmNOqoTAOcIZ3Ecf9prdLSsZOGf
Te5JRn8ECg+BQJu2i7uWolfWnNL/YETUXdrBzD4aE+I+IrMqowH0GrULZWeM
4RG6NYKdetcQOh0lNoQH2AA8dlDaBeigmcCJyfMmJKpNHEQeHywttPNmGkyC
klaI9KPpnrE7Yq0AwCD6q1w5/INXthBFW3iiLsbFkKfMuyUQIzSKSDsGtmCM
ODe0WlGl3xbTBdVFezPbbiaYMB8CYyli0rZFtqgHhN+PBr3DP9u3QGy12peW
/XKhjLu6VdtWkrMO89BZysMAoreZxwbNgdwKMdKZfyk2IA0kO5rI1PjonOlA
2blRo7H9mIkR40wVbIOLRq4Qs+EzQV+IteRS80njSr28Acwe7mWNpViy/a9T
YfFKYSZV7LGy6k2HKmY67+QKhexpewocQDR5OaDvhsRso5rCIlDszEatdJyh
FiRfci1L0hgUQ1tS8dOzSs7yZcZWUSCAW7DbR2DPtaup7wgiwY2Y4hw7FiBO
jNpqMufb28aeQG3hylx8zM0u6hrbzhot/T0g1epshx75mx8kg/OwWyhJ0unz
DrSayoDJJfmPcGsp/1CtNjWDQQVpdfPG5oWkP+WCJqI6XXDnIxBbZA20RU93
niV+IJjZPc+VBDDk4UWIEvlUiCaVaZdNvZm//DDKNe/KbzAuOmED7zLkebsv
hLTUZLVypZQEmD9XO7N1mLJLe1WpEruYf6fAPwyzS1d+VZE4mDqIr2zl60b8
NAKokSk+lEMkyp0Anklidr12ryoyziegsiw2oZvz5jp50emcVjIZtYFJXexO
6K2PoRkYpA53x6BfMu4q/M47FQldWavy03gptRgJLYLOH1GjlZ5bbCnHKk8o
LQSn8F5oJ4cSMOmNQQ6ou0P7+2Y0vZ29FQFygxOx09ebkJnXCus++3NMAWBI
/b9HT7YeD9rIxpPyIUD4m5uKwYwemhmSGzG41Khe+Rtelxb3hGZ3VYMFt5R3
+rL5YvAW+/ytVUdyLluSwtc59gFE8/S8kVVnY5YHcCI0x42oMq7DtTuQNw6j
kAw/QOy0x43hQVYNiED26WrnJ4QtrEKFvEGvRTUlL/TQ3A7llqTq3xKZ/v6q
5ORTwBWV8ivPZg2Y5K73PwP9PO0Dkzr8Y1MBnn6/ogsFaGuaxVC/tORfMg96
dqwSKcUv7URPkbVNviISvbhUUUUp7eXcgNcPFBPYnOJqukPbiroQrFGojkBT
e1wNWe/7CbFkLlqTF7uTFYNBsrEtPZjMW20Zi62MJeGglGxvv7UpqxrErb3n
PP156VswD6OXEiuHxoAc8IWypwG5gOQdOAbkeoDCW+I5e14tBawNxyNfzwWL
F63gZBWuMsGRunCljgfiqCG4lwVM3fDw5WNVxIkVDe8awJuoiX64zWINmai5
u/6n98la93SkQ8A/C27ns9KicfEOoMxThjmnaBQfiPubDp3jE+8p0O5svbxL
WsbIw2xKOlaAmpAPxn4lozOzfXYH0FejkYdQkoz70vcQMmxWo6E9O3keuKyB
FsTyTs5ZpYjLwe21tQl9MOhOUGpzrgICGsVgUcbSFOG0wnNb/X2I7Ng65Zgk
lxAv+W2DXUX3vHOWNzy0T4k7zmaBGC8t6KFffw8G3Z+jnzFkFQJLTvoeQ8dl
YT1cYWvKt7+AiVY5L0hw+0qV6mtxXqf4V6k/pAhS7QgN4IQkVgS5pzTx2fVp
Uz2R8wFK99QNmYfVx+ALZtKYjYA9iOVOrCyUL7NJnyJb33ytw7nl/2lJVst1
eS0W0nzxZyFcfqge+q1gfdPNhdbywyMWsNvxkx4TbbXMz3ZOiMEotGy/yQlJ
9sjSumwgzmhdoR37kDOqtH1EqD3LY+RVBEUB0xuaUKbaCD3gyS7AY3q/rWD5
QWC86T38IodgD4NPM6c0Q7VDT0+/H17ieyHTySY7bK+ic9iuFPlkRw/OTkcX
IowuqchX4Wg7Cyo/eEBPmm5Cz1YY2qTFxZRkNez0rlnfJs2m2Hvwg95EFsg0
aPwhEtly/ksPK9pkQJsO1NF7VTXNhvk5U9R9oXJjxtma6umYoWO81I4C5hBS
XOeDLatqbycz9RSRLMRy9KBA5yVLZtKiR+R3sESjlubRwLpEK8mf55i/81qO
bfHCUEB5AGZmwo+ZSfR2cDsUY2N60wiLvTMmNgWD+yeITD58KvAptZmgo1av
zWHm/mjj6+65yxUz98IMO/z8tEcKm+mnZ9VLV+H3o23kFJwXW1G+bqXwDKkT
/qbQoC7C1LI94bAAnqhQwpAWBwSA2jBiapG4wicBAfEisKv1/bKrWCsERV4Y
wTA8d1BXKF+DjQVs5ur+fzQyTPD9iIYIzStlpDVVkyqoX0Z2ilv776g0URqc
BMKEPqK8m3dAaJ+uGJA/H9kMS1sRtOULWbfiWInJG5YGROQg0SciPIZecZyM
UdDaziGDOPge5OinqxnwE75z0P6O3jKOzhkOENzBypEYm7bIV24vJg0vxZ+N
NTm2wXMb5wrbKhUVi37Fk0a3hRPEk+1RlWKCkfDTTjBZCjhiyQhBAX2DOk4p
K5JuLABwc3Aj2sOX1j6Q0g6F73avlKWcOHIlllK+SkIwU0kvZ9Ix6iqPsmXL
a8S1OhP5zF4dyYLBUOnYQfMBx6sKZpJvBZv+ChNZnR+6dxWLa4uaLswZqqu6
l8ffT0YbNRG6lJTVNKYEVGqX8KksYtS9mrkoZgobdaCKTqEvQwG7XxSaopSD
0gfwKLuaPDsopn+LZKKDKiEAa7FDM7WWb5rumQs0cVAf4nSgHKtc5FgnKkLU
huOFCOf4uh45oFKNbTgRWYVLM1AyvxzgPZEp5cD+22ctTCpQSYE1I3oCQRnc
rZr0wkuR/8H4YO1ki+51u+3Kj6fyvEEh/Nm5uitcrxz7rwjjormsuFox6XBw
jB2ZOtf27Pz4Rio+wYkeWWiObIZQjjaQWECnG/nese1zHq//tVfK3PoWnnAP
Lh2HC4/sMLv0TQhjnnZ6CKJT4ZnJNkh2WNvna7OpzRnjaGLBkYtpiukfFp7Q
4cuqamCyUIqyh7ktPHJBJqZVLDPjBNcwcICOCvmOXuLYxYkAraJpvk8oMC72
ltW3zbM45NQqAvACmwZVJLWq8lMe3QSODxPiXQJD09hlTJ6pHOfBddtnKPTs
kyEf+6DUhGGrSMwf53BbudloOEYQiyY9GO8qZGnK1CXsGIUqAWqQopBGMdct
zRWJj0+gfzhA6IVunfwwUGGetlTDE4ZZwbHGqIfBYfPnHYfY5d4Up+2lMafS
oM2KirMfGNtauA1SiVxxVHiOVqWqRDTsJ2H94afNYcO0QOYEp3Ntng0JtyWD
QC9OjoAynwmoXUuoCFX++Fvemh6npn7DfvL63r5/Hp3tCHFhVqASVaJfMtfa
dr/gFZI89pstdaJ2ciNrn9S/Dxj6s2LiOa0SHvvQw3V+TPU8kA26v2TYqEiJ
5JbcK5JmhB3NcwTOi8+6vM6blmveTK2ZrDX6sPozOUM1iXXCSf/0ovGGTiIX
gsdqulM8RXNXkt3N9zB+jAtOuSGxrIl2EhCm+p+H5BdIwqaa9y0+zcwPKNm+
25luWnX4Kqvvh9m1Q+zkRUAjEktPZBvwE3VGUtelboK215c9iBi2uFuJP/D7
NLtom4fyT/yQOLJLvjU1ykSZDivPRdu17tMBL6y3NU7uoLqdxlZuIl8iGgji
GmS6RRC7q1+feLBcvMkrxjWQilQ4ee0sCxo5PJY+ZHOpC1tQKj57uG+N30sR
kXBJiEbFC8R79niramxs4OkFfIKQPw6pZClaJ77IAiP/lP6PeYYXX5eBvtGW
wtpe0/1UAtekkVIxwpWFyqN9XLYQ4Cq5wVB3r0YlYlUsWNdk0oNEV02ReBf0
UftUGffXXpNmn6eNlwe22gTzdIwfXGdAA2d+Jnbo4Xyq5h9t0MXCe1nkoini
832uYV/Ho8afXUPvCfJe5pXjAelT5oywJir1F0nbvjIFiluLIIMJn1Qe+TqA
+ZdtBIkZIhHRCDnjBVna+4vwwXXdjqiJoHrh1Hfraqx20Hb2kErkTnsTPVk3
w/E3cah/rIEhAHqyW2sLMGOGJuMzcvahXhqslv4Ezro5o52Wy93fXXiBQJSg
1UEIGBQy1Ag4QI2oKji4kYfixehA2ifzxGw4Es+cUG6KuK1hVK83oN51xmt8
C0lZGgafuJSXbL5/tWmPHl1lamAf2D+VWGP7us74ZQYphFIyqgo5fxP4iXnF
8cnkmgallGBXwDj7EOs184YjXpeEQB6NRq/Kv7Y7z6o1P/lrl78UZGymjN50
RDjvDO7rNfMgrUmsmB/zchepFV8X5R+1NJso5i5EZcSoR0Q/8l+IkxTWmZ4h
Rnnr04viyXVsfsucl7cl291ItVfaZEVeEz59SRaabQp8BM3CztoS7FbuCIFm
Vzr7oQQhne0U3sLi1A7uYhOwkhuazgyw4ba7CN+WnZEuwA9Z+R7wVyjVCm5z
fH2Ne7f9wR47uF2D2giuFzHa7VYLyoDYJttnaPbeWn/M6MSEiyvkQdrdXMpe
wrdpbiHuY1U1wL0ROJUCYdb+jsb57cdel53z42mPVK2Cus6Yh3JasrWW0F/t
X4B7TlpP+0vre08RxwfAI20X846NW9AxHdW1KcCDenf6IRmd7x3nWxBQfoRL
uaPz2AcxcedNyHi/Rg95j0SNaatWJwU4NXTpQfTjMpn+hXE4mw9bSc//RDVM
LPlp4IsvO7Dzr6+w46f1zoG7t3Lkc9fyh4NiiErbNdzQeokM+DlsA7MA/Qi1
etNoX9enUFwF4+s3qRNzulHWxtK/Hea/LzcJqymIU+sLD0LaC1gkuwo4G3H1
7Ap1OD1zqarncMx0/GMXhsAZXkS0kzyF5yzXWuuFSDvfTFwT0AK6pnaYus3A
mMxOWe2bp35C0daPbaoJxrYy9mOFS6kXduK1VoG0wQaX1JlTEwulRfRtKrXI
e1AhLVfvX8+n23cgs2k2vj0LGV+zhM7JfGeXTqgPGNJeaCyTEZBO8aljw+fb
AfbuNoGPmH6XLAhXy5+IfisL8omOVMXoP+hnSbv3FnfqZLK2/CzQwm1AKvjL
oSu9qK/3+bEvkIn/hrmK7ROool3Xnh1eY9OX12jZZ8MNLNqf8xqN1U+/hy0F
azkrHnWjYED7nWrI58eTR9DHH9KqBX4lBGEnLGFY0B3zEi10jqQNqkquLhCY
Vlj1MrM59Li6Nf3h6bmlO6c4PUAwraNxp0/KYc6eUtFCuRhb6d8/Bpcr4ACc
SN1o51X17CQ23qEWlTpO9/Mmj+4wnvNDvxxUPs93VSt/kII+/0XkqKoO6izB
oPn1N9hfBLnnPlevb4VrInNx7zCymOIfpifYFQOnHEwrUagVcGLUI3or2C1M
b5knRi0tAL1ycrsRHE25VA9YXigpdmAJvs6q0SBK8juSB0BsSuKwT/c0eniz
RvqefwFTXjFNIwpv4ll0pNI+C6o7Bs+64QSMKT+NW7iJ1X4iWmNap5UtLBT/
vwSnt30bkJHAeIFyBQg66BUrn/2GC4MZouYggOB/YqjSlMvXoWZDTqw6wUWg
u84IXjH0UlDFPVpn+jtr9UY8KxKs2SVznTrYSo11zqIWHx67ruIahHa07KE9
T4CDN/6dfzoQj2Dci6gQQho7Ky1KtokJ5QXcsydzF9Z4qJd95Hdyv/4nWQZM
cJTI+aDC2gouabdXxBTzk1yI2hOQfXhVZDekm9SMv7VKUkplbmwwhvtql+6h
FPar0jGOZNEEjG6TxJGC715utM0x1Alj223hE/vb2noGwqvAzQffawtVWQZq
WGfR1IPaL6ECqqJQuVtZpiM9vlpNMxfvvTymd0RqyBnwSjwyC/n4lFaBF2gx
8/aAMmCvYv9TNRoeCu/sZnyiV3gNL79cWmrARlaXCb9R2fOH/92mr2brK2RX
X6SOdYK71sJ6s9z5AO+IhVWcU3u/p3Dw+eN4EhEjZCHj+o88uvjoq7fkSch3
Wv5gxFY30eu7fYtNn8jGhHTbO9peUrMq0PCiAIKGM0HFe42m9aUVqUOk1HBK
AxAwjTYIlN3ZqZOczh3lqUsGe3rH8R7s1KEL5JbQ57cqt/NDgTLFbX0WL3oH
RkCooj3LufcciCXb/wzVKcvWztd3aYfti6IUflnggQdYRUh/TG7+vM5rKFw7
gCqXVfa2xSNt8vbmiubKTZhqJoF1Ce/SZqfCMeCQy9HB6gslxnU0hf4VUX2z
TvFs0akcyF+eWEN+KoxunZCYEC1kuxN0rbnWxc+WpboNwtGC5Pz2lLOWZvAH
MQDeSzX4o5lD+gOHJ9PTPA0t5yrWlwbsGMoyb/rrkbMmjXY9w4B5u+ZDIFUF
oiegx9RNtA7zzHIqxT1EAceKjd/+6RVl1ueAzt03jqknTSUh+RTSdA4U2zwj
T9UhCi2hydoebyHefBS7UZQZx63s2wiJS4aaf1SCsyR0t5j6DkiQoJPbH8UD
ZrQ+B34VEsvYOWrWFf9EEz1vrGkz1fhlhV78dHt1+SQW/z4igQXao+9RF+Bc
/ziL7D8ZRl/+tJr2j5anHFgXFLwHRbctvg7rFCGoFrTycXiWpevcyxNF3V6G
uSh5WHaceZ3N1uhChGT7ysiUi9tWOz83iosEwpaONmSBe0g+m8emRl1T5pg1
biRVaaH9t2DXjfJ5laKByC9gQx3nT37eKqO+Vb8lELxdrZ4lKAcQWGXDkF0b
yIqJeRwZyjcY4ejEwdxjWTXgRqiUBw5juLxL6NpPblGNhX7/urhtplU3wJXU
Vu9njZ+RQ1vFiSXQqZ6dtjnfCFdWoPqaPM77uzYj620PQKxc2hzM9v77QVUu
n1YUIoRLTeJ5kXoLixObb04ocp8nOl/f8aEzSgNtD75Yyf7v7CUCZ7d482Re
ON1dERoi3wdzZRamMiCskckElwcN9OvHOIl55kTYqPTgStr0QYUk153ExNPZ
qO4hUEUWKcE+KxJItSrFgGRYAUjnx3pgmG8meM+W8cIz9R2TIcui4zJ8nEcs
wxUEqWsUbcFtLs8Hpo4OpOXgFc36l5qhhAu56XNaunNSWlkbwBXEiIjSQ0pK
4IQ56+B4HOeOnf1fY/ZLAXTgNFE1UyFs3xE3EdXeDzUtRv/K7X6dNdxqL5lX
CAC8WiGjZ45IkhtytUFgsyUNmOs1uckHv4jLzw7xvA8IcWQbtB6PKptuI6o0
5omdvqi/xiWUBZMqjxtLrd5tSndRBKKk87upuSLE7bAHOnNV7XBw7O7uQQEe
AN198o7tsr+1FydZJU9DPiwrtjjflzTV9zJVbburjU1JrMYPGiZBYRx13dMg
9rVmfTPsdVAqwz3R7QUtZiISEra3UEVwFCwEYYerHOzZCHJTNEU/mISUOuxo
Hg1J2nkxdWiqW3aqK03VPTB8L20QtL1yKClzMgl1I5Eb+FtvQ/2g9o7dMqqx
vTBicT1Y7XSfmfku3x6qD5A9A8G6Kv+kZFNkj/kIjeheNPiTCYT3kiEFOTTH
l9tu2jzR5my19kXwnwieWdXNWdO/Vi+h6B4HF3uAdrmBqP+rX+NX4RoXFZab
RNWzCEs0HQFBL9X/dKPOWXzB3NVyAuathbGWqK8FMANcPAIMfsdL0Pzx2Gmw
yDwM3so1PCBrjGJnKHPfwRM6guOaRYv74CYgmOqDOuwMjtxn7rctl+5Z/VT7
hegVdcPA+XGoYIp29JkSNZvY9lbcoa+0fXA5Xw120stlDEtjHJrfh8zL1tGZ
+otXP18y/icSd6rRUJbnBAO9kMwniuhwhbAwr6C1TctllpCvrEc84b1Zqhi7
RqCswwnZP4qA7/f+pUoOGYzTnIrAbxxbhbaEgvr7PuuOa7dR0Mi5gAK1uGjf
a8ITBve8bAm42F0slDz2ZJ3F/ICJ1N780pwPQIAVdcefJzEam0kwnyeaCZxX
YCcGUKFb8B7GBQ0lklwq1ha+9/Px5r4r+GWvf3pJnE8F/NSQou965lKEUMKG
MCoPmPPgYObZPb1FIWfb7aPH3wTsiV4ytU4I/lGguDhD+lA4wj3zwsrxvFdW
feHcVUkqQIVJqy8dP8JzCmDF7m+t1Gj5S1J/+BB+rdSVDHdf1ySj4HexW9lL
peIdqOU7XtRUNm9Osv+/Y/CllhrvYPoxvftDQg9IX7qV4sYdDqE0KE6P6cHe
N6D7jQSUsERT44Yh0Ng5GqAUpWqCu3Wjvpz5zQexx8xLYgunLEL7FfkTU6VG
waWGNAnXAAAU5JByV1nYFqqTCaEab/ZdR1MXFr4Jd27+wOFQsHzU3y8GAtUA
SRwlOwJIIuFr4og8ccjE/DV5dkV7g7cYt2jrlofURZDU7TjZkQiTNnEVfOex
OnBOqefxmyWYPD+CaFmmRHuBtWGTlfK5JY0r/BhoZA2/kMjzB6jmT5mSa8/q
Ru7F/SnuTmWkZlKq0+BTF29OJrIHFs+VM/Jf4voAwOvLMQl1WKxUJxd8W4q+
5BhkEkZ/g8ojaSTdC7dUr+NZpSaSpP5cEvPch48RQlorUJu4+IFuhI7zu6h7
LMlAFwbjVhAcGH4mtTXHFeb3EJRBLpCkA0E0TpovjZcC8HifPbUKnYj+S6dQ
K5JCZgV6aFvkOgn0x3TDXRNmgA6liMOmSXjnFXFQBYtJr0AOVWjNJ9XQkZEB
Nv9hWwPjeuVxaQTuEgwk3QkR010+xtBwFbVStsUIfgLKWScnO0F61YAor+Qi
Opd+SGWM9AZ2o78VLy6T0MRsMDB3sh7eVoH4JWSZCUkBhuf1QE9KeavX5hGi
HhZrT4GKROMmrou+H3uBgn0tI0fXXlqboBAK56ry+zzsW1RDJbC4AkjoRovH
AQf6ehHmB3PKtkkktBbuneuKDwta/YqLUgg0SwUEfFiJbixMuU+PzY8x/cr1
lmEkDcl5R1tjkPld3bZKG0ZOiWG283BW3mVOw3MrsIULLHVoEo26MOnxKYbR
s1m6MQikzDYWaf+Rs4M58S2DUU2yZ5pDdShJaBqs7Ej3L5ck5VEBPUAHNBXr
bI3iJFb/bO6KGgN2V0LBITXKs0KZSAc9hyx+4WcanFLzF6ND22CB42rbEee1
VN6m0GZFSLJC+Y9WxfO3ysCo1nrhWjLAK7xhelJFYvSsbcRTeOwf9mrUYMcx
0mpWz6AC//1e8qzHqwzRoALS2rr1ZDewjyZ9hhqQXGCjO6mNmQXT2fYnlBQT
vSY1CvsDrxLv7npQzwDTrMJASraT9PcYT6Sb7pZDxEHJ0QD3H81TRkrSDkyi
3zfgmKevWd/peKkEB4FqEdtq1wfwarHAqwinZXnfTpvcNGJuC2nnQiQNnN3Z
S/lg3Of6pU5D6tYdTHXzslyl6VTepjpJfBQv7qhILNajbh9CGanwUwC/UyG+
YhNRDmaqoTKpGANOgmM7XrO2sGXEO87H1ZUEWNqvo+JViKZWEUTgtAlCqGsc
Lbifn5N3zOUQSWUg0gKXmeZqw6XrhwMs25IRRJCo2Y00DYwlhyTlMZtU/39d
10ONf8NgH6SDoaPWUQmcW2Z15gIhvl3aSeOs6SnRUTb9oeSTEjytnN0VnXL2
v4GBEE76MhQjirCMiAWBw+is71DBJSMlep0I0eA7HGg9nTdivWwemK6DAwdB
ucJ8G/P1uVIqIyLuVehLjEtjDEGxVJlA8GyOKX67NM4joEMCmSoIx5lRkUxy
ZnAorNx1FrCnMyTQa+K4XLUFPiz0+Md9EPZfgi0yt/Nu2ldwQ2bkVx1+MpHD
xAxGJWsTmcQG+VmX8ir+SV1p+RCtp4tUSmpNWT7bWVGksuitp6mxe5SLzTd5
JQDl6d2Go+xHyDLGNIlQ3saRycLEoKSuySUxShQWzBjAspkeQKIVQuQrh5A/
RdanMKi6p94QUq+idaNXPqLzVHHSjVrqMjMDUbFvL8BhT2f1mZ2z6pW8ArkG
rhbWxvsmRH+IkYXZXTjo8xASCt3qAB1Uv7RJShHo9P9O0NB0FE9sry4SDhML
UWZt/bVmYyRDAcvHNFoRMORPJ5b2QzjqsDOjLLCPB4JlWAHOtHEVheraeF1u
FL3i3DOgdZlXrQ9jzH4rXbKLjLttyg5l1X2Dbuc2Du/0jwQ4NE1J4T/fl5GN
etqFjPtVTc10PyTdVQkyfNM8VIgvV0+rRXP5AziS89JD8H/69kJVscJMsHvX
sM3MnUFbOTZRxK/mGkgPa491EVo+TSygH/HVDTcxtEZMeEix48EsLCtrGDKX
6e3Maa3QbJa3Bao2e8VwENeDE1szdUfMowmaFoWSNUOIU6JjjwHj9TDcJrIg
MypDRYEuja27pt5HeX92aROqsahlih7UOZyPBjdTH2+UXwNfmtkqaFyYc3g0
dzZInvHpfsE6z2I95PP5UdnRXJHNHxA+mclB2CR97PRD6Gn8t3VJktIvPqyC
ywSvvXd+JMG84InxNBCpD35lCH3ThKvQRJfbsQVxaNtIHvQl2g1KIOh2qvRi
D76PCUU28yT86XUgr+osfErg8B4XUdesQ4DQrDfCQzLHWHCYJs+1lLqG2LJb
6CvLoGD4UYfgmbeH18dOb9fon8UBRcW8O99HYjDyC/6JWPwFxkCMa6MC5Dca
rBSOtHHIjKJaKXplzef+C+CGF1bAZn375C844fLTQ4OMm+yESq+RS/TEo6zs
owYsqslQimtVW5QVR0SQ5Tnt9LQznTkODbJiYKXtauKRfKhL39er1zz9vh8+
ew/vA4uE3m4FgvrFYUtSb5J5J+CheBXD+JAN6XPqJJKQP/15uH2lsMsJ3plU
UIuZBTNk+vVmZlwsnr0HLPWpiIJsWNAHJkUxucUaUNPsELuqkvr9TJIhicUd
3QZ3TAgaCrwX6/ppwbzWGks/mwVNxRvCOJFNsHV2gnUGsIDHZX2YcXIIsw5a
gngv3DDDgaf9Yx42F7l26oA3FqsBFFXkED1mNsp/KH61XUKznQUjgkkkrSoc
wO5kjONlqXiCYDtYjmrIn4BHQjs+6QjSNWJ+HHNZvi9bA9SzWOmogn82dADp
vWL7KCG2Xin5ZMjaNX+3c1eOS507Lp52MA/PiMV1pY+p5dLCFdmaJsZ/qrOQ
WiKJZHRQwPYtJ9Ij4VxSDgQ361b/vGaHEvv5oJR4wqwiFag/aCfrSw8xX9v3
7bDfkIQIqBMPWe4FYfVT2M4UVvE0yCNyQvk66SYeZCjxpYo/tmzN+yDJAXrL
M+6HfK8YJpEtHRwi/KW3JX/82n+kx/GP744c4WrfSsa9dHq4RhZTAZ2oyh1P
tqejFAG/6TXBgSLAAHv+BZJNc8ZMr5LgJ8BcHAnXFWCVm837XgHs3brud1vP
uzS8lci1tvoxxR8eRBW1hWO/dRT1zsa2Ladiybmz0oNYW+6ajTHyOQrdXpmU
y3M187eiQMES9vMqC3ibVYvQuoPsI26swAAYMI6zPp2VJi9j+tEDH5Enb+/p
d8ski4LbGSG9+uKbTqhoi9a7ET98+7TINd580DUXnLWR0QN5vRy7p3sc0JWC
gUcXXlD0pXGaTV1NPyBUsayuJVjE40We88+gz2ShJJ6H99+JmXOg4VAIr8jE
/c9kkCN/UnGkgHxMts0NDtnyfxfM6abULWpqxqP6GhBNKwWEXIrds4mosTlS
Q3jjqot0zrBXznkmX26njd2s8PhNjAA9roy6lhbem3+Q8BcgiKWSsZ5ichy2
T9t7MJQsoD0r0Bd3Q3oJGQZF/fpCxIGfe7SnXREzZQJYrE5UozoTokQI95yN
KBeL7F4c7YDLFLpHVOQDuVCaDFTaS6KPxledOcd8K9OzyswWE/0/CXr9QoZh
4gJsCqH9JaQ+cb9VwwHZdRP8pPd7k8bvJYDB4cpoXTYHwndSAgb7V6yU/son
XUduYfeA+hQT5FL5rP+Hvtyn0ydngidph5rd4kKYuemSfB9kZAu4xm1BaUIf
8r5ts5ort26b2VFoo1zFxsF1e3Ct0kfe3S7zeiZLTm7Q11ihTELxE1FlAoMw
hE7R9UlSJ4/4yf+Snk+TEXDNVma7FQCFVJj0YVz+64L0ejpEhpi4TFLOy6LY
/4b23x3tdS5dYLsZNehY8jp35YUh4XHiUkG9VIcbo6TwyzTvO9Sp3a57aqKq
h9CI+7CC5inGQE2FrfsQYevR+T4P6HS6gXidpOVTUSYf0QVb/rypb/zuqYW2
qf54kMFNnA/ILxY1rpuwyBnNSocrPRVxlAy6sW2VW3uz3zim0xnl/TQn64OR
5USl8i4Oe76XQcHHqfZKVwSokfyw+Mfzu34CsIcjdg4ikgHd/6WMWoIqLYXm
vNpk+Jihqpz8FbZsgTN6mFXPhzv/Qh2emmBpY6cufe7qMbq34h+edjmPxnwo
bu3okDQ56aAixSpP0uvPMb21+a5fev6bZXEa+/mSrZjQR1e+dfowmGNUIR9D
2TydRohoTvnzx0v4ZrP7RLZjQRk8UeXj7OfKvR0RZQjfy3ZbE73XR1vu66fq
8gBgJoZkXHVg8dqbd9cXBAau9ewMonIUv8jwVo3Nsz5E/1cCrOSHM9ozep9y
81e6cgHmnV369LJJnyUjlZHy7P5zG2sc+goQvKTHwlFcCSJwJdwC+g4jHafk
laXEL5ti0zuVCEpOyUQebJyBRjxcmDW4Uy5gDMDHcvUjPa2khT1I7x9hAd4M
CQ8KweTosqioBZKFA5sdB0ixW15GTKBRVM6xgBONBh51pzP6vz/vuW7rAsUn
LFR8mT7g1GmvRumj0xiyljGLq5+AVOqTNnNNVIWoqNjTi+UpWWXkPkRuyDtf
j14Ngd4/YUxHKeBTfQcK+4k+bvz3CSwduT0TjcsDBP2wdWM+JeCa613eh6Xh
Qd1iC275WkGCjw+pKQZbg+gk8NZc+x+Xuwh+yakxv8q1cdOaTPhlPKrFZxvo
szoJ+yZqHgBKYFR27XAvp9e4FeiRHebanpZlm7EuxVzFCr6piuPDTfTyKbwI
YLJIWp95PLv2knOzFCGanQfykUc8OGBg5BozymOJ32aEY7MVPa5eQpqPCpWT
5oyAL6HrBFPkOu5ya32LZYR9YC8+i/Q6vCabwS4tZ4nwNaUvZUSQOQl/LsIf
RRCuXbWOzdtsIp1M4UeTRRRAKABerdpzA3hry/fhoVkmpqyqQ4cST4mLDI6Q
BuzAxYa3lXhq084/zfZx3lHz7mt6X6FR1HIWs7xb3vMmdTLOMgjqSgFwELEd
VdUxOeGkM5O9u8AuGEGPRP73D3ySxcsrmxzozop1SyK0gJqWgdEhOC7coJFC
It0ERxqgw4MR6t0X3n0kNDuPPoI02h7VVnkuWG/xBxDqT3CH8OpwN580rwX6
IJ8WDatBlP9oyUJ1c0gw8HFkARjdI5z0seSzTvzMbeyfnsFsJApKGgyARQ0V
ShDNXeQaaKzQpbiwJuposCmlnKWWBCNQ/1BXblrWQfDUsOeXDodqfi4xdyoA
ifLo5ygNYJHWzBn8dF2T1ooY4+m7lYLWLkTG6nkqVoilzWJTu5JXzuBIQdpm
TAqvvvdpPxnykWyCtQViUVpHOAWTgJgSodnU8sxTNF8o5K2Ly+zxYd2rL71H
yhwxtHsl5JwmRi4TiV4UVcOsM4PYxlclW3lgXAn7O6/QqWP35/Lk/KpLg6fh
SLhNXz+H3TL/EzAOVH+8s7q4PrMLc6vR3ZNUO7Xc33hbmp1Z2RUcmX/Y8B3t
wWURfQ0xk12UHBgdZ6FgtXpvI1GkDqzd4/RaqkPwVJxBkgB2wA4lEdHwQ4vX
jRdTaM+UrOy1c89YJ/zyh8CtGMz+0vq3Xff7rLJaRUqOBX32HT9T/jnNkjXV
LbEBDoICD6HrUoGegPjZJ34xyyLaUULAKWyGwmHegfiHz5yDMKevvVOByoOK
Vk7NzEprcuhhekwd8SoQ0DKb/pAemspgMFDE34udBJ45/3MEJ4TZGGymNUcC
dyMgykEFPc2UQ9mpghzHjv5Mdy/Q8XpcH8JLyW/s1R+lC+CUSWuvTqOGoIH3
bY4LiWkOMWypfMR044RLWknRYSaiANobDNdwhZFPLYUN4r1jCXXSzUTYP8Fu
0dOlJPvWmIo/m747/e34eGpXjp+0QqCxSKuM/roYwZAKa7eQZd4epHvvFjBk
xSqwo3nJcp0G4nXSLmzAeNcrvPWTv7o/sZBctTkvPLdMNBHyakTAsY5DEHGv
/3oHul0w4LdU2RdglBBMqwU/vuYbu3zwAcRQ4sZBZhujwA62Cep/MgorDvRI
5BYYwm+tPant/Wd8MpvF8sEHEKTDuwfezfso2zM92TB4A2e1dy6SLmlO1E/F
D9RJSssIGROQjiqG6nJwLeHL+mUO5IETbjOJpBTjT3j1uqsThkuvJNFX3n2e
8hbvWyLYSADU2BMZZ1XbhgcN/z/YyexkbyOYN68MGBBkgUkir44EhowPzK3G
EjllWMFzpNoBuMRKtgPfx3rHtpnLnbcZcQ9BBrlA5cTTsy4MaHjKIGe7TqE/
Nm3GQXXonI6rZrmnLX6VVl/bGjZfG/h5yYJxrvHcPNKjdVRDU5PdbDS92EAd
mBZVmXbI6/7AYTKWshpS0+1P3adevZWSGiPWjtK6jrpYutSd9Wykb1vEEkAT
0Hnpx99m89x2/jFSRLqX2IdXnbbMcC2Zq/LL4wCypeIcryn/3Cz8uyXE/U/G
mqURLJQsoIeSZ4LHDWPISb2PsQMEs1u8gD1YKXzUV6y3SSeVcBheaoWRbNiW
Zn6vbCv9Q67gZy4ecvh+OAr76nZe9jgrinYTS5JjJ2bIQd4h1rqQ1ojfwxYY
a3KcGtPUBZKYHBHprlZ5y44BhgJr9oOUY2yISlJt6D+ikRXsZXHnbHxzAPf2
JGtgfnnDeI+qc5oZxAdGbit8S+Az7HwaWUadTs2hwYE6F+vpPA1vwZvZt01H
Up6QNZJDC36F7j84u5OEs1xdIW6o4mzw9ScLHmAo3UhxX4Ax9RX1djDN6TMj
iavuE1+F9nyZurJBklJ2tAEqgzpJIAo2wpLQxu0+XxwZoTDG+aSs6GNsMTbo
+ilbQhrswzaYOB50JivZQP7v4+6PK82XQJtDuPe8HwpEYExY03K9zx07M8WF
vjeyJyjKJBz5a8D71GpzmrAX8gly+bFF5KyhLBpAXwYYy6etNZZokMVyrdiE
PD2qAU8wCWkqFoI1nLFGMPgTWPwGcZ5v28qTVg6kdrNATX4w7mVkHTOsoIO7
G7PzPuCx/uviYlirPaR1e9eTRtPqXOAcqJVwjDgHlyHlyV39V+kIeT2yBjS1
ux/cNq7hHUUWeU4daFqx8uflS2D0DNg/NVXBGCwiGNHhbjCMu1VJMEysjvpj
X1GgZ3gYBnRQu3Fy8y6LkBMzB0AnyOu2FPfadtsi3ywqrP0b7U2kG20Dq4Zx
2+2zAtjCDt9N4V06VfkWPUcpGTvybZKYXi6Hp2R+s2BpZ0wu70N1JE1iEgwe
jp2iqrVJgcuMxpe7CZi1PDqizo4qllcuFY6FWQ222bmQsEzdBJQIGrY4tqXv
JHWcuw/LIPp1VYj5ZG3MBed9ptevjE7VHceMrsrg0UVdUubO0wC3oi6/CSuR
nUSMUda1B4vUkS2lDi2YXqLxqsFEXvzXEj5oubcBzr9vb1vHsXassaTHVE8B
4Z3y+6xMa+E05BVU5m0kNzRG0SL6jSbDUZCdWodSE86oQMmcZeO3nbjkEXut
X3QkEQnKuTdrlPs7ICi/BKUfueA68a395mlbOtvkI+Qn1yiQ6gfbBcem+HBF
n7CQMmHHN/jQM91bJMjYv5X989qZjG5IfJ36bHGWbsxNIL0bWAjIrUYklxML
ef9JoERmCS0oD3BLZg3C4MmJ4oJd4mFczZcKGcgeaw8Y215lNZqhb05WEOzM
slRPj3nLwUOiKd7a5gMV+kamovLhNVtWXCv5PdhiXxqr/rPiX2dVCHCvuzEd
PFtmND3jYE7PLF+cLwYKAIVeghBwFxPXqWV9hIUXxWClt8Sf0xq3yGKlLQ/K
5OSE+IGt90B2PBQzf+TBUd42TkRIuh6UazxoEEOi0eSZWu+XPP1vQiuNX6cM
v0Z+6bpf6hJN4OYb8DvGdCN7GDQ170CQltQMZktEhHt2E6hOoyTo2e1kBc9J
573zdn7b45FpyNK95ajS6qLDL/Fzi4DgLsz0WEDtvqz4yarnI8gS3dR5VSs7
E8dlCeYG7nVmaI7b4LR0sF/BdR2sTVmdCDx2VFubG2Sc8fo8wypf1N0FBKnC
Mae36zSg9s0FdgbXLxs1lOCczmNLwpy3z30AoCYSmz46QehdKcYU1Xh6Vf/L
unHXVyyN06nm40ZEkhI+KjmlxphTCa9y+o0R/UEyE1MqNHMbWKbM1NmMYvvh
IlMbs8F4fuscqKfFIjoa0/87WXNFHSfNYQeoXlKBYDySyVfjW8zbk9bf+POi
fJ6E6q+XHgOj3QU3fzpnNAFCUgX3g7IfUWJkyBdOY59SqcHRdnE2qvlWn2pg
yVTj5lnAmFUtgxp4lQZ7YV/Je7V2ES2UsjjFhCpnSNUABC4JPgML7FsI83xG
9kbHg5gY4cUgWUBBI3saTUudQAipscBHf0ocYeIV9WICSJwi3TnOod+CxDBv
oal4mxlc7MPZeqRacBSsnsCGAOZjfvmak0QQDtffb8A0ytt0vKfHDv2cPzFV
SON+E1Kh+IZL20+uuvG0uCT95mYibonPgUBHklbVX72M8x8JFv5mizwjUh5a
0Pp5UyZqx5OzFLDvKWc3zPD14hb85udSsAUMrohlhkmQlI69mELObJ/El84k
7sWwsBPXYbrb5FvM1X3hQj4xKEDeelZ5XxjKorvqbIyWi4ihBrG7iFkBn2tT
/Vn8KOkNFXsWbMpsgt9h66jS7uL9ocMJm5GPgfLTBoCKsqS3/F2N2EspxfTw
x+pFh4S7EUW8zWBgeexdHXgbr6FrO7nxa/+bk8SHpUjGNnFxGvMPAm3X2ldK
i635RyLG5WnkR0s4I1lejPl1RVvoGxxjCyxWaXGQn2OcEI+Op46Ot6o1Cbis
O/E2tHzK6daYdIOzC2FkW5RYeYrtvKYkkTB33TtxDKfrZXYKXiNbn1fc2N+P
sZCCKTUesunIRTxdUCaLgjMKaH519pAcI9FMACOvIPpr79qWVAaLxi5k8PLl
cNwc7AE0qXww7UZTnhtEymVK3QVtC0m/YI1KhxUyRUag1FlHgsJVp7EalHsT
lkb3koHqaXulaRWmMNvfnrYgUByp9ZslzkU2HAvUdgUvC8ea9xvfzkpCzDCV
N2AKfUwE0gO8wev498/eRmtnF70kFFmpeVfJH6vxO31t+NTxICRPthDz6EMX
pYpb9ZcjrPFdKxCz796CveOhraJFtwdZXYptoCiyiP8UikPCaGPSS3riwdhp
+fw1aTGaFgLb24kI9I4L/z9gDR8jv+uQyZQERU89xc5yMTzc2jRp8sHA1Asi
IcYTsThSqUHZ1PZxDeOsqzk/6kIn5nNQi0qQ+afFCmUU+loDGYtMsk2+V4rU
YaFIcXusCZHahovB5AqtVvLGKoPl2idwffhOo+UmsXieb4ZHesZHhMPedY2x
48l+c6eeiUU9oP4XdTeqT59SyoR7ak+MSTWLhN9I7nc8RN3sUfovH4Hx4XgM
XgEqkAffXTg1HVSC96GvPz4QDzYPcPiFTdHkFXZXfbPgg1D+2pWLknnRAVgl
EThRqAmy/4ucA5BKA/oxncuN96T/S4YIwlzU6aX+HrCI049yd8e/grMq1CCH
EZQZeO/nbKLcAxtnlmpzgA5c5TspYS2Cfoy+NPHQPWtQURGYLrwkPD9KgNiQ
+TXC9qnXtaakt9UUThmKEmK0g/0bkvQRKZMyPZR0W350XyQLOoRKyDXK7PSv
2jCnZ5aAJObfvoIF90R0qUVqHDy2A/3GFlCwJpuK0viozVoQkItuYEKXUlKS
pz8oOsTkAVT/iEiGl3XnCOTEFLhabWWF1H4bgRbaGmEDwqQFsbBH4mABsh/B
R5/rkjlQrR5cD/9Jy99iM7dPTwWOsQ5UudfYW70cTk1Is4jFUsQlsoHFOpia
743hdbFARbB0ydgcbifeafqda5ZweD+XhgN65iVKsng4ZKFYCiqAub/9rwgh
eDlCnaiOetlfPYnC6TdZDGUPtTWCEqeOPJr50w0E4BJxvfTmt+QpKsCZ3pib
/u/z794GkesxxsaUBLyHtU5Q9rmDfCsf9V2sWlTRKGY4vy1AcONeOQ4rWKJc
fXRg09/JmEmK7JEuGlxrmXcT3L07JMuF1FrbnB5KcvbKP3SZTjsTo3rwvxPI
o6ah3513gxg7l25/6PtBO905Rrfl3nQFfs+3pdi76Jvjl8TuFseBT5VO04Vs
ICzuTURD4Trc3QjFrjdEJbOS0PNkZUBz/8wdep2J6ncHq5InzFDXIUSK4R4n
z3JuadVaIM4Q0NIXL47XxsbNJMQhJfVlznT/5UJykwd2KElbcf7G+2OCQqEs
Z9sehXNm4dacPOhAuf0BWhvZP02yscTn9lwu26CaHxFCO1aaemUF3UpkjynF
7Eh4/LYjdsE28n9Yl6erdcX9W9+orknFIm0lR4sROzMi5KG6XXzRpSVHFDfj
mmNIizaFLfNvUHlvKD54q3cuZzRzQWtrH1ZBNgzwPL4FnY7L8+4tLVwjaFf1
hSS331xwsR1UxUFqOj+wiDU7smrhKJHWJKScU1XMRD0Wuzoe7AC3DQlZfbPk
xh0yOogvi8cTmmeAgyBy15azMPN66d4dzN7dL12dZz1l0VO6tM6kXnoNWDyj
hC5uTa25eNuPHp33L787ecM7+t3cThSlfxJH91sj/DoNlQE43FgO+yrpr0pH
bo66rbRW8AfMZvoQ9aszVaITWV9O9q8l91XSWb7zoq92OiVPtTJWhe1gj1SD
ZtFhCkCcffuoQC9NNWUkMN6vpDOX/QDUAfOC6hfAonpGGd3woOMX+GkgVg0y
DN51rSU+RX5cL93Vy+mlD7nUYh17kI9OmefMYDAYkLGxdAYiGzSEe27qzamW
XTFefMT+lTtQXeH/Wv6/6NMOADXtoxabmH8eE9SyMaYWM8ElmaMUIPvb2fa4
XnoEC16Jl9bxR51+vGMlHADFxYQRwoK6ekk59sEcZR53FXZSo/Jmf9rgfrgl
K/vQnPkrg3ZZfjVFI+ppnRG1kbRQH2tNFA33rGgC4pfgE1vw7Y+nZFq66E/9
2Jmmq5Mq4nga8Ly1303lWiOqBV/wiqCKw9p5AfZmuqZLq6DzXgPHOx5zh0LK
U3n+sUC/hbuv+kmfgpLY7hlgynMpnMysEjhVjktEgH0zFsqqpRl9KfnWE37x
mVLiW6HkGRni1kE5b2ymf4QE9//crgSS6q700OnKgjIUy8w6jZ486r8fYo0M
Gmo6YxJ9ljapmkpYzA8myHcrX6U5CNrPeqAXUw4I5vHKIRsvBSTXWXiNSusF
hUvgnRTe3zA6YyXlBhgM8KUuVcndqOkkK5PrAEs82Zmvkqm2MG2FBi7IT0+W
SVhJVdV/qtrWFDsT8OCI30Gxv8yX8gvyyHC05m5I5NEmL6EnLF2rqyauLRXn
Aj48P2AC7zNtoxw/XIhQyJTp4mUsctsRqI/8FZ/8QtbVnz5jy7NZrAsSjFHD
V+i8C0JFOG/CY301rib80PQ/zr8mR9Sv+GtKOFoqZb/Mf7RM8RaEYMxHki5F
O5ueO2ibpbrUDmnDDExnQ6Np7Rd66OGZYq1c6DgkihYVCfFUbkL0FoCgVNe2
VLXxfPPCEl3l+XLT4bMlydAVtBzniYT5Z5k19Ke4/XsOE+HgtOG4zWavqeUA
NyKtEGgOiydvtwWv7RnDHSRmo/Xqfr7VU7ZuxR86cyTdQDn1zQEhpLb2frK3
u4bbM1mlsG2pgpi06F4fOW2ZH98TVQPKIK6auhHGsGzTCSysPXFqVzu0FZMa
oSx8nDYRDn03Gp6synVluL3c3we7DTXtZ4HAL6DHEGetWdtzb3w9Qm0aMZn3
Y9lWWYeEWfTr8Bo0cw4qMXWeGGiEqaXu08Vggx8F7HYK73UzHOljHXRY4TSK
1XEMo5nFSPsfubSH2UrEhJ6jN6p/SzamT5YHjULzuVdTwkgnxrziHYdthfui
7PD5bcbQ0yMH3Aj1NY3IDqF4AlMr30deCbbhPBseHKGxYAZjzonJMMEILCN4
DJ1v0VcGdrJwIbhUxOmOFkWyTs0dgt+z6oTICVYJESeVom7/kVXPf57kLlWl
3+R+9BuId+yt8FpUNrVT+oTBs9O3puJW1dBg2Gkb9qvxOfUTAd6x2KjTnbBi
lvF1rsstIAGvEnxUx9uuuT63Cvap2miOez+T1DsPCOumlwN4f7ivrGJZh4jW
qk4M7CGiq7sgrN0ZYXV6CMPoGeZYS6/KKmpbRWDYqEP1mW0UUkI5D6E5jEjJ
02yEcfHHjfRKgVdFDFt2wep0Z3vBj5bk8Cn4Hu2Ug8+4iOIuTwCvgTpSMcPM
O9Rwz5SF5HMz38QV+JENBaWcDdiKiGn7fBd87b+dbc/kaqY98dMRNUpg39l/
Hd48BcFyGoAiSWFZnWdQMGaAMOE5cP0RCSgX8yqPiFNMDDB66YkmI/i6VYgC
WK0Sw992K3VVA0UNxXX6eb/8Gk2HKm9RDIf2HURQNX/VmYVymtiG5mqSYn4X
/wB1vFtVp/ru/StVRrBeylbwYnq58MEAMtotpL1TImmp735aMYVJ+jo73qGl
YZl7CsI/htL5Qq3KcK22lQU1O8ax3kJG2QUlpVpSxdab8RhAbIVf7GEYfU8T
iP/OvbyjNkrbK5p3QCnoQ491P4ckth+x6VbjvhSxpeUgbAw47RXwXGMTYNWC
3vKSRowEBrspNTDG/YVM2kEnqeqduGHO26Bvol5jIrPhRkk64SytTwuYVHZ9
nTEix0rNABxI3IN7Rhru7cudg6Ylswu79PAki4SJx0iXXkts2/T5ViZwOTsW
6uXsng2BoqXUa1nNTJ604XmqbV07zzN41RYvB8ZCT+8qWRliLRAxL2S7n0UZ
UxzuIyOsukenWjYnaG+akBfVfcJwuF0ak6HZJ6QhfNYU4b+VBc0HmuHDjEJi
trXa9j0nlrT6E35eJQA7lyQpIeKa1nWSMXqfIy36hB+qxSxn3vnWG6OJHh43
oKaUZRZnnAGyHjdNMXKlaYTsLhjkPU5FY+oHcoHyUY2G7eGB6pJ+r3N0gSs1
sg1Bd/z/7fDO25/NYgfyKeizxGPZh85ArsQ3jWGC/cEXuoO8Xb816h1x6gTO
IGAFID3nwVEptexkGwOH/g5G4riEAFdDbrxiZYflVBLD34ZElJudugL0vllE
ACDJUkX/rcp4kHiCIH1m3Ic+8v6IGMOAthkF8qYPVXQ+Dfp4xJ6XNaBdqgbx
aKhlBuysx+dTwIzlnVbPgjUvF11LeISxCqMX1MESJmx6nbnkpfxbGe79u45L
YM6NNjPyI7D6qtaUxLlc0XrwR1NqxSBVsoynHNybFaxGlyuk2+bdCDjxfcZE
j4h9j+NfzyEEaHSz1zrFW6z5Au3MEmWj/xq0zUdR2xIbUDYDzGNvSWSNzcqz
rdQkGJfSKewn7DiBe88sVjh8pHB4UInLSWxX9NOflgwGF208ssp3KNVJk04j
cQeHfSFs6+tYhaQVMtPaBVDhOvtndZW8IgrgvZ4zvLwOUF4NhgnWihNPwQ7i
ToCOFMBbnVPwW3INZUO1jRkPgIsuQ1ZrzpoyK+RBtdj+C+2MXQ4zc8LZ+qRk
TtKruFf5++0fX6gB1rH5cBJwmMPBRaD4txuQPOLd82fgg3wbi0Qk/rgbbBPI
QeyE2A9rsUW++wXmjVdubnwrQxVAhCMwRTMu/23cWgA1LElqKHQ23j9RPWSw
JjJKY2Ah++2GjAp36XSpXUdXL4QHswRMZ5FurmRbKN81T/jzfOgGJk23gePd
4o8NW1J1a16Zt1RYfDcRcB1JcG1AptXrFbVbNAVk1fUegdZpd3ITN4JRhjEx
vbx4gVeaN0YPrI4NJDFSZCZbcEXoI1jYtQ8ebkGqLaBkBPofIVYVwbapWGJj
p5NGA/6NqfklnAQEy4S+AzcUkeMI9NdQJbRu0ssU5TvZSmoG1CZTVDE+uYUI
0IcYQ/SzB5+F9UgKsbZJ1bAy0P0B8vodbZuQyN2jwYUQ2z5pUSzF2sfM7vMP
pBQUywGahYUtmiiwvGZQbo01qVbzfmPjMFbC7Bkh6wBpNs4ZyVZW9SOy+Xr+
JvqGEJ/8tWzHEfvYlGfXELOCgh4l4PQpLE4mZpjogLjNPqpyqWXBiF06F7E3
mXz+PDWtxtHnN3FbCv6QIr/vI5CFEe2kMYibCgitEHG6cSMQa0Uc3tT5nEKw
H4Buo8sKwuu3fWmxabOu2+OnsvsBraVu3F5cVY55qYjX+I1xhgGeden5Ye3A
4GMysmeqbEXy7Z4Rbob3DX6IyaVQXslGuLoCC59E4ncXhr+B4nA/GYocc4at
73VR/QNjIVb3hyIlnECwEDzt5v1uzdZfCkTGW57lKzfEdiQCmoF8knblK8V7
1eun0nhmhBJe6x3Rvn0Lrm00fnx58rfbfIY9IwMmbOpTZXWsPbtMdKQpcn+S
p43qDz1992ZLakSAi0T6opywe23TWyaQzZqryWqcfGtyUkcfbd4twDa/c2Nq
1iiOhgKwoM3KOqDDkznlfYUx7YKJUVkyxqRa29l0M6H02EU6U0BCveQA9xHE
9AybLQIGwCeZ+G6E2e9WBXCWQMfJo/fmFtK5iVsb3F+ag4Dp8fGL0Wuf0cc2
r0UGsMLsqkCXck1I9WmMcM08qRrW8FgAfZ/ae8I4jZePjNBAdXyPuVVf/9vh
ZP8tDUsDniVvv/D++p5GE/50+xUk1ErxLloy2bThQcIWRr3XB9DrxGMRlig3
79LSWYSmGqbb5GBxUfsGKRwmS6vhWvh4yg3gh4HzmyJ+j5fO1eG3XVtzwCY7
tsraOjyEWuqqpstu+ke1nR9EJvQMAhdeHCGgGYgFRqQWeXR5/GdvLB1897/k
S8nFIcGXkNsob09o+uqwIg2JWvuSkwsiHX8w3nY51sDZqTGQRu89gz5dqgNw
2RKLqgvcjNSkiAN2E/XDMcg0ZAuYImCrXu6EibgiXmBKZDGZMadZe6EFuimu
5dRGpsuB3/MNKre0qqC+rIpGNiEGYKdEfAq8zPaQ4K9vDGMRiHX+z6GZpAJP
BWAqJOSyvuxUHPjx2I9ZCmfR/UuOP4C0MTJGLumjgRiOq19sAr+oOjOB5qHX
di4UYWQajVZCP0u1jCggvT6+c5/sbfbv4L0qkvrCgyAGtCReklvP665gidl5
M40vjlLMkm20H2EK4Tr9XT3c1iphKpC2OAxmOa6BNeV/tgFcpNLtPI1OMU9C
Z1moOjWno0eD2NLgZE/JRljks4dyLzMiTtQB8qBTA+0uaMhrxbiLQ3cVBpCn
Cdsvl6GVHBkOhtWLCvzsbLlgUpkFIFMeFmx5sEHYVoGuRA88Sxks32JVyGu2
6i52V7mzZpQghZ9yxbRxr90L3kz+h9qQpsMDv2kjWT6VHMPbWcYsbTpdAkzB
Da2pW5hC5ltaOmATN8Ii67SOmPi2gXdYgZHjZM3sqfeFlIbMPzsfFkDjBi3u
T4rRJCr/MF1wEeLMYulGTX8Cp9s7xJq3QmKoss8WeDLmspW/HXZc4/mXwZPK
0mX25lBg11G76+V7/adRuD0bufgCd3ez+hNQA+pXzX8dS4HQMYxTU84BNHae
eSydrOcXesTmOwhl/mwlYgUT4XCv2g57hD3gm6nMVZG2FCYoqa7klRp7GFtx
mGSwfGlXO0FmtJv1RwKPIlIIoCkNUsk5pGeNQ7M8rtNWIOcxnEclFmVKoj1/
vlcQow45gZfm2SZRK91zJzXPcG5sn9J334ydT52RjvmKQJHSpjR/ZY2TfMzc
jS74Kvur+65bpKWXY8fGXK09TsZV60DZ9klylI10Yq7jysxggRecyhjA/N8V
s6donuvmwDYV9In8NRcAd4eQqE9DPrGiyYzwGyb4OLVg03j5PnSz+aWGAA1+
FnWGBcmfTbLeM2hQGCEIPGl0UhTNaj6IY0jMqz3EBa4cLPjXY0rhumZ9V0Vf
P67oNZrBWk8UPSHQz993BOGxXtIv8bT2E/rTPouNt99uBBFgHLdXYhaPI3nQ
zft8uVvoCL6xTec14aAH7lNo4g+qUA8oOrfQhaPaRR7NjJdJJMjDtfufzriF
FTpGtIqUw/TuOPl8rhcl0jicLYXNf4n0LNrz1r4vcLQx4Mcf7MDVIYLR/RnV
tJWRr1xJEhjCc6VnLg/Vq5mGx6XvrzTkqfrY2C5nMtF2n/brlA/UGFhzX04p
3Ft3lM8g28O7Pyzug40k9Y3cFAO0CCGoLH0wbsZeNP11sfecB8YJ4jLzrbFN
1c/G+yLXwpDKncddmWqR4lAA/CYQNc1ns9dafv082c0SMQZuP/nnIw6bP1gG
O0/4wlfcDCP1ZBZoia82UNEhM02idjWCX+Mu+RjhHneeN+tHuvWUdvuL0LA/
xA+mYoYWiswuvvfYl42tJYOtULSwEP4jYNfAFbC/PDEvBvkMqADzVJRf9fip
HQwQ8QETclrWaqG9QJUHL6fcidgkdXPvmNLrcAollBJh74OhBT6rzaIFfOl5
/Eg5vSmfFALwZhHHtY4KSaOqLWX6+DgmAq+CmNkuQsfYYYSqpdwPq2N+BjhS
LNa96ZBUYbxJe36ROHGlk/ubTBPGBZ9YM7jafyqO68PZ2PJs9V2yQ9HBN9Gm
6u0MkKwzT0gZL7Y7UlubP8gWG/mXRR09DlKJ2Z5YvYqKv89IlHZ+wplvEHK0
qNzW0PQS7iIucZGILBGUs7qgrPc+r+s1mMksiTborOkL/5hkqedv9545pls/
LHFEYtfXzGcNoIJ/GnvB8HY0BYKEevQfG6s/Yx41j4pUbofZq/kGBHzr2t1R
Oc7LFejGy3D77CMfhnwDyz3v9gjogI2x6lLLLJQjKP+LukXFbUMm0ER+7XbH
uq0JTUxUNoFBHJ+NOOn2MAMqnONmO/yr9Luqtw9bwJCL48+ncBTGnwjAL2/B
kNZcdLQ80JupdigYYTR/VqVd/fNRbaO/Eo8nqYcOTXULaLstsjfS27h/d/1R
Xr4NYWznvrUq1dtbd5FweBY4f/GZ9v14rHl279EhEP5kSknDU10qB/mSyxeK
rEwI300tx+W+6HIYLaQmHQCXeyvj4NS28c7YTHxEio6MTiwzjffI2syw73Db
mlRwJNla6nucnMOqgo5pfNXq+IR4cmyZ4pudIsibjjBIWdPw6NPD7oL3w299
mQwVVItjdjL5YNxYhTeYMkExi0vxxCc7rXt3je3AI461gBRlAha62zd1oLI+
UGASBu6JMJeYmwREnEa2MPKnmelviu9xK4ImAaJ7gcP9l+ZY5ScN4oWJ8iTt
vzFyaOmMwdcfnP0cOQhHKnglU6R+3/+eVIkXgSH5hbLoYsB41W/YHP1bDdbz
PpMEawpfQWPEMF6dkBh4agWLsjrB7fgO4NgYSIC6p/VQlZhUfHLBiA0zYuzA
xtOT9zDW2oxCXrqMDSZOjaBpFNTD4jW6YjhyS2STBPF417pxWIHygJ3aIiRc
Q+PVMBAoo8lzAs5yda+bnLSDiLNWwuel6wBgQmhsS3amntkgUn0EudsdKcN0
4bBi3UBpeD0VL46DbbmKPvodRaDEaQ1My7zHOSi/t0V0wXsP6qjAKziW5odV
vDv49mJNdwly//MhHfGXqxLCqhsL+X4fSKF3qfkBcd1YD0Ocxd5o3hZJ18dD
zHm049Nm7KymYtvBXJBPfRPRwWqatFA2cR8w4DBBSl61QZOvnuyPlGMjBNB6
yqweFmt4b7MstYlnrb5ArWs5m78DjPY+biyXnGRnwz91CJXKIv4UHyKF856v
k0Io3lzgsqKb3hS9XshHbssWxJ5fvDKfQnKe6CGiFNqSLaRCAEzr1dkh1rUA
pKBkGr1tb3d94PkWNlOllzddY3xmz6JIjAfTwZGsrW3nrt60SBDGbfgz4yzD
116K0q4+nglkJe+Pp5Scu3WI+uXsub7P+R/0KhBVuJ1TAhk3bkMHJKLwD9N9
RTh2RQJR12XW215qBfyyf+5fxpDHCIOidnDh0Is1p7PFOTI0LwPGik/3cWjA
vSrOQke6Rzql4uuSjCBkBmVan8zeOM1Yi2KuIk+QU6831bgeLwtNrKQeKbSz
Q7EW+7gD3FJ7yWEb+Fee0t6AL8g/NMGemAaODjqZ+SuPp4OZzSQqA1q6rG30
+XPivCioLHS2eKqujInsMgXfyWlApjpd71bQ6aVCT6xPvgZLGUuPJ1tmQ5En
nxvP43kflVU/sLu0yZcLXN02kVGDeJ/0uIjZrerHyZSNnb6LfroFtzDDHlqC
mpMzJj7rRTYN9hjdYFDbLmRuz22eewZPf0Gy5OuxivP8xesiSo0Warkx4mcr
iQNmWYHa02J2XXxLg1Zc5GipZW0ly5ya2ugb0MiaYh27DgrHn0afFzMKnIH9
COMBAK4fy2mo2pbizeR3SXIY+8ZzmJBJKHZ9DER18EP/dQT+b6pE10gbA2/N
LAg8YNYBOmuczLgnUflUko/3grnVnC2QVNb9uM6vQfVcNi/r9Oj8ZwjEW9VO
lOD2yDBB5lD0pFC4u5zGyN2tYkkSoI0EfoB0B8nFWxfmstfSucp5t5SYgbPr
SCyPoMqnyInpmGv1fsKNP9CmU2rgE/jedSp5Ik5cfDLEsjMeBcC4179C431i
OGCMms0hYcb/dqUxTPihAoLGjPCHcJ25xtNd9qRULuQ7ekgQeCIqcIe5Mgt6
oq5vNoG33K60qT7FPVkDfADwUA1CVKfHfYKNl3IgVuOo1x2WcB06oIzVnQw8
Tp+VjYx2d0k4FF7dr3LsF7gIrpbw4PVNl/AexfPWfhBe9nge7R44enRpKe/M
DgH6R1KVQUjmRCdwce7idavR0+/l+3KfBDSuVlN7hxEp4eNjN00cToFJ/XlN
yQZUjvrSBjsPQjI64/BZuiPYClE6e3cyqZO1VvkQKLGqMCaGmjT+hhBaZQym
59mZqhAiepfg+zrbn76U8v14j1SjcVivsA6LXISC75k0hm2Hi3/cNXDrBLgb
3FqAdhdTwM93XJotV2u3291RC2QEOgQ5QA7Q6T5Z4BaT1jgVnenfeOmbyyHL
MGmJYDZpc+COop4v1+TbGoG8Us/AmhCz1M0G1ZzXClLgwy3Q5xMSOUcQtqPq
YslYzL58zzpdcW3Xkoxl86vN12wVL4zg88BU4LeiRDyhG1Y3+Y4aifpnvUjh
VkSMnRmftAfUzr/LKTHxDy9Ng5tGtSUGqymJXSWMO7kJ3GhLDAV3o5hNe3kr
2upGeujNsqQjLPwvt2NlHaCV+Y93OcOnlY0XiS7iuMytqpKogrOx5PQN/N9H
gVHRHeImOgH2rKJPBmOH4N3YHmkbQ1kMwqXl2lqu757e9ud1M97q7nQlnHOD
ib5N59xUWh7pCqyc3k3oTvPaZsHD9bdIm42f3QkywZNqDA6s0M1zwj1wjgic
od5+SGTBt5ZA355VObGMn7FdOdY0cJjxyoiTpv/vitwFgDpoycQLjMwHHBBq
Ql//mCQGO+P1JEBoi97nZFg+eo3DDAoc8lWeTBO1XynnHSNDL1fjEHTlP68D
dxgw9e+RftXX6V4Rf15B/neZkzAnwWTfzrHLqd6eppSyOwos9Tn9KW9sfNmS
2xmFPGOfKPGg6COloa1vUbMDhM5wYum5y1toP+q7AMBNApB8yo/0JgnYjJYo
4094J7b2LBUgjViIlvsLceZFYWi2P5qs+kjQ0P+GasFsSpFY57L9GWARSUUg
NHje/fgCVy3uc9DCSc2zvtAq/t3bNQzSQKOiMuy+do9YIQOXMDTkIfhHEXz4
rNzkbYSxN9WnMu9Zf1DnLNuqNGDXVXZyOIpXmoWSZLDfXwewgJg8LTLRsnys
8jJtZc4JH+FbeORHw07HuhwLyCuDaVp/Z108ZmlpMPu2kBQMVAeOw6fGsmjl
zWjHFf+AysUbOiTUI0KnOzv5qIkijFDGoqapfQfixvtkrcfNJ5BbBy8L1O35
Lkr5dZn/+nZrVCrv7Nr6GX4ufbKJlNWKSeW6zbrx+eCzPbC9P9eaV+l3X7SQ
XSatl3RHvZvpDziylNGjBYcuBbHZ+6qoxAhlopgXlrhZiVGzVIQVQRSMW85V
b0W0i/mMZGtSKbbBz3eZkfAjamLOFNHwOz7OBlyh5rOFBWknT5BQfmYqGAHY
Tr+mznd99ONwZYLzVkDVABjuEDMmUs7dGvvwCJWbt4u+cdX7DiJ1JSIuLGD5
xUlD+gXluoMbQpRDcIhkPrMIVjX/t7RMK5U89SM3CQvQDAusSyIQL3pyrlGe
TWZepcqQsv9th+a5n/mV0NvJjhQGQyxmtnrwNEbpslwZa6iwB+pndqSDmDPO
3rXzyFpvRY82jzygP93L1J5o1jsQHRCfqHcVjFxCaUMEKs6BGyKEuZWA98kX
PNyibXoJAxGyLSAv9htDy1foTEWedmH+bG7ZQ8F3sNC3PzKEpgMNgvNWuHWG
/IlZe/ZGScsc7oCHKjsJ5kM0FG5ceyUvxMWunlLab4sPmXGp2vxknz4l+Kss
7YeFp4yTMBpk7Y82VLGqiAYcN3ViDH/0LN1p+Oza+pXxx6Hvmn9ozP5no8zz
BqGB9YieysQf47GHwLyjaS0SEamRdXufD3WPFIXccQF510J72P4qTw+epYyK
iOc9O5Fe3glWxTZK9QbqBHTGzglhhBqkqdoR4mwpc5yIhRuB6Dj+KDnjJYob
LP0zZL256CT67nxiLZp35CYSPCrHth7rZ1QL0o5Q/8BKV2ZC52yovXhUW58u
E/mRDq6bKKEUcyr6rbOYUFFTWXDK3480EglG7Qb72v8mRcB1VX5xpb6JjBWs
wtF0dJz55MIwEueMjV5MJJzlIn17kG48FdrgagdTuWymoCHUEI2U+A7ji9fW
9Wm542D2qNNYJBBwhyo07oq17rCVaERTkldH8/iEdUPsTmJ4fyRELVtmeKvm
BxyQwVRSFObbaLHMFEdm606fEf9iVrau6E8cWo8bxxW+wXF8VcKbd/thixdv
iRSut/X9kS98y3wm5Y0yeY9n/tXU1WjT9/Xv9sWPfkrWTiwn+Zr2PQzkjHuh
+JY+lS1DxzkaQNq5P8JqU0zsjrrG06vG6QcLmsBGWXZbvoCf+JERjxov3BYi
20BXEJQhdNO3EmNhX9RGgIu4X9qdrMMKIJh7CX/ttuPi/nHikPL8RCBvB6iL
Xcfz2j0PBQRaKz7Hw+FB9Pi10IeIBXun4p6bw+qTisD2rdoOQolPm++j4cG6
HQija9pk0jFcDG8L0tWYvOH+9aJN2+AOeLDnxtnLAU29KB+mJLJ57aAt2lbc
FLemmXAfyQVG+C2qtUg+LtSSTVmmB3UO+dUBx+tS776wAJ0qHHXwAoH8gudU
cCaUHL77u3Ro+PPFHnVMQMyOz89hR0O3T6uRRMw9cX1WqllKYMAeAjB/x+3r
VeOMX3vaXZ741kOKCJ4Ueo8ufk2PG+2Uu/M/9b/0930rs/tRY1GAhZfPLDnW
ejCNTaGI+sy4Zu6ZKAc+3TGPpaQ+ZTF7U21hAPr69PpzVvfMxmbQ3GvF9D4Q
1cpPsngWblT2fNQhAEIQvavX/XbqI+410ymfKlV3eNF7LYoPhTk7sGOTe0yE
th0Z+3rCSMR5YIMbg5g+vT6wkL2+PLtzOn7wuBJ91EbK7IER6zaXHnnd67IF
Cnbm9BHXpbIv9UPDZtD02XmgACilNfTHPMiX98MMeey4Bkd7A60xhdWtt2o+
0cP/DkuwMhH/myKxWFZhm2yaipRKnLwWJtkYRaZzq44BNlmbKst0Gk0xE82N
KO48yDYs2p70fLDg2tpWiP1Fovh6lrSv/X4voxiZRl8rAXXhULhuQjnyEbfO
/Y5B0M6cAoJ2mnXlZdNuJYvIOo7WLpK5bRZSUAvPl3652ySN1Jqizk/gK4WC
t1kbW9lANwTDpW9dLxc6Wd+bG3hLYK0Xjw+IF1YoHFtBaQAmdOWALzDeXDEH
+scptfctHbMtcVNron4nQMp9S2WO+2xAIcUnWZfwIWH6vgLBYhtElTYE/Vas
QRIXLlthYcBewAQs9lULqi8IUIx5Y9KBVgDMgrgq2XVG/sRAc/m0f5+jdU3R
JvTb2tCHSVFe+5jbAZP+Si2HzpsXtk1MjfLfNXh+RsPTw0nR82Mk++QbmIHR
bUa6MH2MthIzO1BM2QHZwQsqGxsmpsmvU0I8TpuJdpfaKy73z7Anfw1SNCju
nKMF/aeHd0BVfq7eLh7dhGbdk2UPkWf1tckunePanx5QqEvFrrHCd0e0qEDP
SsWkZQDZQBmmA8IGVrbNj28SXcWRseib3XHEUeA5LWUb/SG/mCx5Q9WZNvV4
f6VNOXT9M3DZ+Rfu7CW9i00L8AkfV8vNcotozrGO4Y7O+yRxQTU4Ev3MLBha
IBhlS1MQ+r2I+QIFiX1V6Oq3ojLuFMosXTZc9q8d3G6n5RgcrQkNbNgmLtTK
HPC8BvfR5JAUG4Nm1OX6p7SLgksFsxtBZrG+3VEecO/+VtzGZgs+ZfZY4WP3
WWhjQruHbM3fLnvmEEiaMXqmg/RLFkNwY9mg323opXf6D37JWFCPo79B/YwH
uErRWVNWP4ES2DFduD0tMdQysYPv3IiP57cdz1o+ejTmWSaMwdoRmChUzTCR
qd85uonxYYjs+qVM21H7e38wqYJwHYfEKsW5VrfM8Jg/rBzJZLzoiEkPVB91
iw2s6Ofmfa9QOd0cQWluZCW/bV9Jla+/ZIbN6NuD4g3CFXrJzFCzdrFuuLak
vPLQX/JVsXAqo5zaPw2LbafgEM4/1uND/JGMQ1vTEI5hoJpxa9Dr5DF4pUyi
u8WO6eSnQoA5klQhSHrqDLoLX4SA3LRXPCrEOI6V55S/YQIqdfUVsjzqr2uL
aQvR/oVgtfiOJsr4UB+KwJANJPT3RWOrt6FotSfTxEsSmlMVpg7SXeQ4dL1C
dZCvnuu6w2cVGMETlhOtsMAOcRNya1pnQpHxglof8izBcpFFfKpz7a/z/BpL
FWNBM/BZ6sxUaaVOMzgwZzYMI/eA5ryHd2o6+8SQbTi1PKdeuvV0/0OqUWrl
C3c482arewj7llC8bbDPZdzAr13iZBarpFTQMRGY6ZEj1MP7IOVFGVIRCny8
sADc4ErjLWSMhFY+HmI0THIobl8222K8AWPjAq7OTVV9jdxHLnUFiMYvAzqx
PDYTm4OAXlupm40I03G8fqEnEH9SP5L8vqj4y5xpNfaDeECuy3N4mIqH0ZMu
eN5uZqeaoyMrS8iqnNRFyJQ2XHmaijAzFvNAx5CvI9CX8sSj5I6WsURPS+iB
DJp6IJlpYf40QQ+bT+t6rYNgUGmmrgGJvuwKfW1JFeSIz/+vMVjCbn9GM1Fp
Cf6V1Xgjpuk5/awR9K3H4j2cevXuPC/TK8hJdeAtGTD6/Lpt7K36P8huksBP
E1IvaHzqXTU81wBSmhwS0ey7vXJKedOvluHNEoMmxu4Ol8B/DmVe++4iP7ov
6LqfmZ32rIMa4YnEaCIqz1nhgUtR2qJasEJYpQoXFb+URc8vScomZsY7or0C
1VFEx3rl55FzHxA8maCraAcV9xKsRQcjHtDN1wJgGhFmITLuPtf/gseViaYZ
KINLC+U3enWiRsB8oUryPk+gM/+kjPuTi7orB7hJkuABJFIbbbfrUCu5qMlr
cXcl6xtFw1/gV0QlwAo8wBzFhG/lNva76LqPidVXqMgjEhyp9DOlFuLUt5NI
Pe7D/I4FCIYW6ruSXTudrp1PY5QwNeLDMXVvmvKbRef6ozpgRa3r1hl8egPL
ywf+BcamdxjzdSlUhw1V4gDovBnpv2D+50EdmiuMCDzcvg51G966gx/YrWN0
OlJFW6EA86Gyab0J/5yMBVaz++e+K7BOEMIVk57hFfU1d4BRYPrFaD8w53kj
QNYLZUvpCmNpTK837Lh3XWwlNSa40T1vUW/1XjJeRoL0tKKlfnVzd9MQ5qYe
Ncp42U2wT980JvKU/IeY3aOpTbutExKoN0cju/HixVtQK50fFHfiEthjKkRF
lohnT7ayNSjFKc/oGb9KyUP1RKgOp6wQ8sOc3wRQ2jDjOpjWpsQRyv2iNZQT
l3HV12oP07Ly37TE9xlMbCGcqA5lJWPcQyfqFUUAeLDoPdvjO8kW9vQZgCgP
eSRzHdJWnnHZ81iaBGKM/UNbJ8C/5MVMUni4fWzpXvwdWkoGthPagpVVxymf
bwK1A7fKAhYJBC4Lap480sCf3al1NwVmnEbbdq5aQRXRlHoL/NsDHAAwxvSe
CZB5NIrcUZELA38FxoIHSz6sVMrJjoxnGzj5VFvOHUN7hjApvJos5Px/c3RO
UYEzal3LATiFhqySWSqtXkZsGs+9vz2x+0aV3PxnXtZtFgLeRYwePQkJN5ET
kXs/KB0O4dY9ugwG6DX4bFsQqORzozAFHBL0OeLJQqhviN5D+eWeeA1LIGg9
N5vC3gE8LbvzZ1c3P7KtcyD6dmduVR3HVH+MGcDkgYdu5apdaem1dni5Gdf4
kcoQvvtPH/Zkd1Y+yFuYX2dt5t7RaIC72eVJ1QGZpc6yK6MYomKwHuAwFCjF
WnnU4dFNoBwoKaJxO+jVScwTzxGoIYfeEUiiRmHHqQplqGim47hTVs+Aubf/
5gt8/fSy8lKJo13jxHjswYre8yltQPyXlSKw9o7KrR4ELQicyHUHW0OOirqc
hkLJ10PyUG4KuNgaFXf+TVDmoBSJPbqKuz/vVr3Hagjq5J7vSaTaHDvGip3J
O5HKjKbzqL2DN/MVS2a1Va/1W+zfwQcl6ovGGUWREGXri6d21O3b5UpPuUP5
AsEE9PGU57bEewG0DpfF78ogUopJZfRcRFhp09G+khZwesf3qtDkhCNm9aKG
rY8HiPQLMQQB65gfGGb1EZu+7MeNG0ws9YdFW3uE16DiMTtR+T1aztQ3xeX8
sVplMMfDYjZb69Q+6URvtbWegKL74Yk70+lUdO5YATbZKoBtmS1cJm7pTsME
bOL+jHEyTdDF7XphLJsYn9HY+XWSKMtSdsorKMDTb6VnsG0d8r33P4/NVplE
bQo5ur21CEZamFj5OSAqGmFJJf+2ox5dFxgx3uMziZ4lFrrlDc7S2XNzUTYD
3i4gCf4GccfoMdEIFuPStiC4zyFJsk1fzwu4YqP7SGJ9WjbnDPB5vrygtzWc
G6copOvn0VfyxJ6pbYnfmGIqYqc4jeao/0bTY0KUxGifFPRiub2bEidAfpSS
B6HeOheK3ITQ8C985fBEyBaCMcMuxi+LZi6mpIZImzT3xvDHBRBIgjqrzkol
L+ngZiymTijiwiwzvYnqK9NZSyqAAlgy8IHjHTW0CxjuAtF15QVoMFpH3O67
bWRlJI5zbbOeJkwQN9tRoTWbigA1JE5IcKQWyNpnQNZI2CL9V47XDyG41WEp
cOkNPUIg2H8B03ePr7x0j13A2ibx6onl+1cicLJNu1XGVsITC+S/QnDF7CqI
7CnJNiYMgZLjD0oc+EkXmKG4LsdZnD+TkWNfy6dYApU5nUU7k1efSvmdoZ+E
2JnUMpKZDDuewWBAciCgnF9L4dTpCot7KwoUUVj1l/pl11Nb9iNk0Wp5s0Xn
xosUltbyK1a2giohrFyyF2CfdryHVH2J64Jp25aDLwitcBAU/gM6LTZj+ajq
vWTcX2G0sS/YQkTihj5IBsqF4AigZ3m0xByBfvjzEtNgCXryAGBdefQbVrdi
1iCBTSzYZz86s52xqycZTneK4OE0Ed6RH9regFQlnJBuMxa6sUoYttnSu7zt
CwiqTh+2/v0U5wz74J830bY9ykNmHRr7Cl+Z1FCi7vqKSi+nceXe56fBOuer
9Y/kSheVao4bedeLActtxKInr08i9XK2MVVbmccxYmbd5AVWIGI1+FgdB2h8
bxFzvkmZe2gWd6njsjNPnG11gTJkN/Um0OKxLQVF9RmFtzS2xPKPIBnJWN23
CMlfOwbpdHoCEktNQ83ZeEIWqIHYFBBRnrJEG2S1WhpCcBbh1qS5W8bp3yFg
wlRcgIpdb5MbldPWNH/J5FZyAUDf47N6822V5VD8h8rKRPIVVh6MnlI8DL8Q
bNmHb0nW4RHD59sMJiSI59CNrPF2+8PsXuHq719MpCbHDHUfvO9eIYrxml0s
1UJdxTK94BFs8Y0p+CZdVnAmvV86EttLiFnth2bQ2BfZolFWZVEf9DTk7RBA
Oa3/Cy49+/CmaroXmU/hh7nwvZ/0fRLeVvrmuPb3TGNDmX1PDCCAF+CCtx8k
fiROsNdtoX+MD+0L/RTXDPf9irSjfP8PAr/uy4jkGAZ1U6tpme/rQYTMfMt7
zJRbWiDTyIhYqafCNb6rq4C2zGtUUi5NatSG6j5ahVvnWZ4fY0AiIKCiCmSd
X50+/bw0ja5j2m1RFFb1lb6QZjSQPVAuBxKRvUex1QFD7MSEYaZY1q9BAfQk
gfhS99ApsKdjvq8K3/4oxT9QalRD7Eu3oq3XiQ5Dp/AVC+GfnbwfVNQ1UStz
K1aeqq40Evl+7tOO72OCCmiSvedHdkZTsLZ8DLs8z7QkjKK1JpNq6Obou5fl
98DrlrLGbNL3SSPKOclW8QxleUplPr8z6cIR4znYQ88EO9Ftc+CTQR7GAXxg
GQjTfJFLG/+ZD2QrFUNNkWwdzFmC1z4yzfaqtAQabppweSEw7II4SC30F/90
XbR1MoxK70CuSriSoBT4L5+xwrDlwzyihBTQ3ngAQeLt2H1AYj54jawLWlVL
r+X/oE278kyptmiFBYQ0Fx+oUGdmHlnbAYGQo0PqZG9V0v6f8YVWPPwemiGP
fx4eL3RVC1ZEjMUqWNWOK7Rkz/gTZSuyo5x7vKQPjsCp5AtL/N8AMIzxWlun
5u5NbmIFJqGLcE7+kT1PuvSLrcfJ74AQQcSmBQD0t0/CzJmh5Dnbxxjon0DV
ZqPgwqlZR27B2EYy1/xrymdb8YtUbhxWIXd6AZGebUR2ZEdea8EACLA4Tqok
m9XMrtXIS+RfstihmSNSLrjrfBGdKzzyEicIu45+M6h00Rp2LfqsoGwhDsek
rrH9K5QwanXoM+WHxUmVktevn+EqMI9r9Hmp/1enQ+ao4hxiXwNGiDu4SaSK
lffsfQmTH6qHDRCXbuS/D0myJWGr7rmen+BvcO4OKCUvZH0VWhery9EXj93D
hyr4+Gsh5vjKeNpa4JR7x5K5iqHHhH2V8CJimc9q6HrtBDDVqkS1in82aNZV
kAehcKE/BZRnPijEvC7CDq+zEb+miTRHdL7dz4OOSI7jTN9fpLago2X49FcO
1gUecXQ7fILpMvSwIYcKOW4TISoxDIudbCJF8NM3iwXR+wgXcUyyiMT9beTS
Q0uhURVUHMo9w9LcARDy6TZZYEsTgJuOx3oipE35mZj+nQeNTuicxq7ZWHl4
AkRVCu5RybFsU8tL5Ts2Hq/EWM6Kp64Q2Bha+nLqfn2x5EGyCHK8R6Cvyx2N
GIygegOZOg+8fkl0D4R6c+75RKubLNx0hlY/wdwoZTS0YiM++sGv65jh2Pa4
NZB23MIXXEQNZIe3xH/L9Xthdh38Z3bxiTOAv2SlFcS4+tFSjLgx0SiRKj18
/dymDj8UwgSM24kbcZjxrb0hq+5YJXPPHggHJqa6qJ8+/egvbhTXxjbVMoyE
EJlN86N1hH1tveNh+ORCTyVQ45GPAbpaLv1y7utFPOsqR2l0uSLB+yl2kuz/
kof8DcYAiy4UERrJqvyrHJmgIShcq+yaH+/nl7MRg7yNOSU8weVrq5J7MTAL
pDtdTZX4+janVPbeA8JALg7NJw7IbbdYQf75Fl6+hMgxJkdbwZjz89lgUPOL
DU0gVqZ969CxkCUv2/HlP9NKgAxYJReD52ykfFSyp1j2cXyBJCk0zONkVSFw
gl8c+Ydx9AkhB/Ilqy1HB4kE2Eb3+0vCNn6mP8TdZn3LCDRN9rGdSmxmRgPn
vEXCxWA8KCyOiWkcurazvqodw5VzR7Hk/ZwWu0X1HQ10M/JMZHZyQSTIv0Af
tgXBYskYAYdzycFDcUGkO7F4kd8L7/1Nd1zkp2liBOU+R/H/alrayqHwBmhk
XrTFTowWxH4kGLTI0Ojr0HH1ENr9bbFYWUjS5PIAQl6AZQ+6zWbltoDOdsyh
AsYRm/ZkV3kYleVUhV7qr0lopkGhIFmg9Y1+mCfqP03asz4IffBFPnhgiqoc
Ue0SPFf/6/dqCWaTSGyH99oGPLFwXMyINbHRBtoV4FUD5fd7ant0WtrhwQwX
Yh964kuNj55XBHibiPwxIndfPPdhcLfE53YyA7uuwLLO/3rb54gyo8juLJCV
5XiylsAu2fFbt+u5wPTmNhTnW66jyMtbsaMzcVMuQEhxt/qsb98v8Arq8sPN
jjSB8nyujDJkx6puNt53fW9rUizq/mSuYSLt1GbNMnsoEAskpKKmtL123YHx
QwUmT3ckWm1nl9sNFdgEN36ec4lPMTa2pMXkLw0A8nHF6JIpK6poVIhfiiEu
n5COgatmCl+9b8AF1QXz+XRIgd25mF+j3XucRTsqhRoyotKyy+etK9g/bPg9
I4mGJ2UgBip/BEY5VZ0bAFqGbizFu/x8Nmbki6FpKswAsC1p46zHDlcAbgU3
807GNj6Bu24sOv3936IJ6g3TF6h0CWRgvMzRIPS24CE2FKazbZememVh+iTQ
L3R42ESMfstQ//LwKcRXIlQDvCwbW9KVzLTvQCxb8G+Jvec6JEoEsL2SiYsv
q9pvdbBjL2AFBtSB//pTTw68D/rBVI5brLxOAHViIHIGYlkv9RC33n0Oz91b
xB3s8kHcGAkVKGbYAIYvzI8bX2zlmWmdzcEqsgEP4w/M2sAPlSTv1ffX/J4U
kdOnYf2U+PqOV7SeRmI2KQhpIt1UyBLvheBF/QRmegfovCWbbF+SX1iXHBz5
/GxpqVsY1Hu3nC3dDbmCnHevag5JUWKaKTrMbOjHkWFMPtOMB5xFLKDoK5I8
VPsiF7dvylextOC5ZyM3uQDH8POFLCyOmjwgUGcfzQIJF+GVmlgyd3/ubhuJ
mSJo5V0NxWxJg3x/wWQNP2wE65Z9MCydxgpwUDddzj7G1sYL7nN+xSRQFY1m
I6YnHOq3/GmY8813BNxt/5W0Zw0/0DlUrdEEkKMDJsP23k5DoSb2CJncPf29
STsDAuldwagauPP9BQUO6vRDp6XH3nkJVzu7p54QkhLobuCZ8HpiU1uLfE4H
EFwMdIh60ytt8B4ZRA8KRQiygA0X8+pJ4NE4TXgFwQ2uK0XLp7FlK2DHRLsC
A5pPvH6gmmTeQVJBQ4dt2BGkTF+oDJqTiXVQlp8WcmhHeTghY7XxoqqzbAbw
5DTLBHHZwHvRKEClyqHyc8kVffhKaD1gf+E6ATet60ZlFjfriiqD0dELf95r
rGI8azGZnndyG52R46AulKfYUZSciwDrlItrfPSBBNyW75pWI3p7sj0sE8nt
Z5VwRPR8Th+6WuaFV0sw8/zPj4lcA6XpM83IvdHjdaRoJnjAP/jXUJ0kGyE6
bC9A1u7yse2DGOE2kg5lLsLobZq+HQ66s9T+ySIwzahGQTx3EuTe7zt0fwMf
8a9GLkHG3goIw4W+CR4vku6OSzgmVtcYQ98gd7CJ62tpUnq/6ZiHtz2GrFLN
p2oxWA7U6B6JvxoKRTIx7NqEug8GlYNWwvn/YTDgF9yROAz4/0x0GnQKNCZ+
OetqFM7tAiw+p8pTUplTkPbVUWkMKZcMlOWuLEL+fhtfxFP2jT9+N5UlxFhx
lutWpGmctve1MbgqfJBZbN0E9jzcbsrFkNYoMUNKqlHcZp7Mx5cC3QDXy0sP
BRFODtFa/oOsQL3egS4lJmV3fef3Gj8U2fbIYr6dmg/Y46H0yDpGld+33R/e
LeYNU3VdoEJEdLxlFoIkU6gkwWhPXGNwvnXNE3wlDJNeRgGsJrxlD+YIDwc3
OeJQLKmlwf4xFvjq8QPWhA1zLXB2i7rZPgBNluKU4WQl/JPJUETjkMZHAP9s
OnhZfugAOihht5hnBYaglM49q7R6s4TaRumOHiDm0ipAY+SkjYOJY7S64FCx
DvUgB7Q0V2RC6UnAtlI8qEv9+sCHiaKeqgwt+sYSrcPYtsUEHCv6UVVZX+nO
kcDvyWQJGzOaZaYFUelgikmMDYpDWiOZqlmFDo7OT5GEdzkAmtmTlFil+gyx
HWw9K4vP29dPFBDXs0DNQR9o+qmm5CqE6mGTOCNYkE9ZM/1Mle/JQqahhvFl
U66VwosUyhyd9imxyKwPpngbwNkix0YuNj6Zx3DN/pecJnbrqff9aHYYQ7aO
WTZOiYYDLE2+lZD86bPCf94s5X6hv1CuxUSfVpLpjd0Kbu3BdYHJKzy/K8Bf
8Fme5uscaOO7lxukrppPzb7ixIsHNniCsE4ARio8Jb9WqFbGQDX0kfoPTm/b
vc3I/DsNiVvArzAyl6ajcc1+J0I/aGXaua+rarMf6umHebwxTBPzDp5poeAH
cJDTpQPTQqS3kSuiLrk3g45G8QOtJ3wwP06S1lkqagozLVwkbXi/amc7xr2m
mgc50gvlgzQbcCnTvnGCc9n6TEp0iZ/2ISNDYAqYTmOrn30JeMNY8y43diXU
YDTiepr60F20k3XNKSVLMwW4jMdMS2guX7b9d9hpxUWFMm9Ho6AXX7Iu4p+g
lTEc8WMtrfyldFm3U45kZO98s0YPHyyj51C89apjKaZSVso86+LDjCxn7kU6
+JhmH3joK7e/77Lt0wmuVqdTGtOnjDQgwxQveInfE8dEjTBDyRdY54P8jcgJ
lHOEhYckoMEMlLJTPy3MD3LTf8OKzNVbFYgD/bAUChcRqf8QOPnwvkJMDN5U
IxfCA8zxaegDAOXsDlQP5bRtMBcMhLAyEmZ1jhCEU7Hl1uB8HYEm/lLlyKgO
hHfRDpNMsjzYoW/M3C/S08fWWOIJl7elg2HgT8hy9w9f8J4S4pjgDmbuZ/ob
7keq/JmbWFJVRBnO5POtHu+cKUc8dFZGQEjtkx99c6C8HyJcUvuu3kTWzbn6
CfgnxK5ngNeY9Y79zmtrHkd+4WsXp2uwiA7LzDyanhqIwt51Neg5dzziO/ky
FYHhj4xnRRCLaKykzmSvgT1N1hu7Wztq544KHaIBZs5+RjPO0LhUxANy4UCy
JGeDcIutncn3vuDjKcwkCqD6tVfZttGAzyqN/66WasvoxVaPBJ9N4qzuKNNV
mowiV5wibFOdja4Gp/9lGW9dptuC78g9uamMskm2zSTwNe2KmniNRxACAWi4
1C/84v59S4jLQGOqSBl12NIcPohP1XPQouSjtMfTBeZyoW7+LELFx8a+3o2C
8oDgmUswGT9bHYsGqYk2rfGm9RemA5mZ3/0DXInKoGv4jwYlbJ8WEhvvHmeu
N5yrDOmOamAyWQoqBno0MxDAMfg7RYMLeBvhvLSkg4+DGK03K7cSNqr/GarV
vSyStG1gMtnnq1gwXirLEmg6tD3BxEfdEdZAClAXx4J3Ul87v10Fx4KWeR4X
Jm156NprGW8fyHLE0T6DSQOZzQZuWF2KF7aHMq1aUnvFs+vpRCH9yfsh5Kad
KwN3cvKbtFq6j4uhdLx7c9U7rC7Sz3CCeE7+GxbwKNZrCrr6hR5Z20HI2s++
uypnxozlgIMlqrVI69BbBj7ZGz0oE1Vg0tyHTwfWCdmByB8h8EldBkPbNhcq
vfZUMY1eVHRI8xEsFs/YOSSNa7BXpTML+ifjbjxe9v+x7PnnXT4xgTvB3ds+
RU7a2XepPHeaOMzf4gzOS/nAMOciyjgaZPny3Kz82yyAMLSCZPcp/sC/joaA
7+R7nMdekFiCV/QxtfuiUl0oxqPeiW5FhvfUc5nARU8BXEdXxCW+19M0oAc6
5e+g9ZfYY3UU44KxBmjXtis8ImiL9JbJqwq+wSjiqBGqqdBep3PRCGNHBTFm
jN/eHpdokmvoSMDDneeo7RMp3u0gE9wUOnECTOw3UI9AyEhAX7Ugxfpewe6o
PlCMzBr0Tsua4tyZNhFEs951Dgt+PEceG73UrrivmUtY0nhpo9+3QK7yunno
D7XWk0X6aedDK/f32DySiF8fJfv2Bg2Ne+larZ/AavvJNhkWTNeNPTtMyMrT
G/76p2Fqf2PXt/wypQFunArTEn4OeUNDzbAlogos3/Lx/7+G1I7AdewTb0am
9+H2Lvkpm0bajda13w/pJtmP5zRansn8eU7fsivqSMU7pb/d9Nt/qZ3md9Y0
t99R2mnKIYTbmQHjgW0GpGY+qeU44UEi5VEy3gYoT4/HoANBRTPPOK9UpyCM
Fe4Vlapx48HXRuOuFq/kZN8vno+QyKK3z2Cniso3rR0OLAG6Ey6VYkCaHJvI
PbDc33s0S72hWS3Dntn0so/5W3cZpPMF52cg74Z4M3bzMdLhQVbrOOmbw0nM
jCnz7on0go1h5qi7PyNIv+JYNHIYoO0qCJkQI2S9h30sTT/XO3nWumvV7lHg
1Cai80TqgVyaNE4y/9lIOHJcvLMGLsm9N1G0U/CmzjFFgLQtfnxaC/Rn8WKv
GBuGr9BA8mxNdOOhtBZuqBUO16NKdJgWiyVUcjDgE14mH7JzwoeIRzTqJ2fY
qPBB7M2Q5BcVGGyr09MZLnA6s5zd0QTpZAeciIgSBzpRgxujj1/3ZlBShhOn
PKbgxf68zzxkLd5690fI8uJ6rcTp4R80+R1Fi91XlrTvfPFbTLQJfygQ2q6E
TSQOHItD89z5L+zTtj+GpkIcVvh6+VSSig30BVSRNCaF6SQ0iNNDZZf1Nc0D
DEoeH0Dtw4LG/Hw4ac9m9ez5nOvFHNky4ReBjY726pBFKrHvznWLr5yHqrcb
30Z5USQk5nk2sCLl7kfgYNkhocmYN05Tpgu3Ov04Ouc/eebmuBiOwiuoEgGK
4zvpihK4JYL2lLGlUwcV5m+Gxh3ouTvXaIpCtIKZZcBKY4/Uu82aWOZgnr7v
5SGc4/sM9RZEAcMfxiGvFtjzXT3llEFdOj0xLyfnUfJ9zB6wNysJu9Cv+tgv
1n7y3h0uMh9LI5E38iR5UClfE64GIqzJoOVr5vtjxES1fnFhHPuLGf/sdISr
WrfC2Rg66FLyGC3DYpDPXyjrOvB5NtBVDo+zOBGrSM4owb6W1cZa3XuLXLbP
n/J9WBNm/K0EPtui0KDJ+RBF5hLto64/TP9JDLdGE05nf13PuEuoXglZBbL1
682vGcuU9yP7auo4LAwJMR9/LqeC2flNmoWute2XI0cGbjOQ9Rybcli17XKo
+mB5Zh4q7QsMcfnrbij/8GO/duorMZaF6D5OjwzxxvDhgTFn9eMPYu8WKQ4j
rPiN6cESx7xEv0HsQIt1Hz4HwaupoxK5RLM9G5HezGN9M9cHRywpLBoewMsW
FSsOiCQUYaF8PT8/TBPA+PEd7LYt3HaUWQO21G2KcvcqamnPZ5Dnp2ZKaoKs
0RFNIfNdoPkEBy80x4Ek0j/wRZtZDp+/A25BQ8oaojn+YqbDqpo9XZOm3e/c
f4NPV8sypW7d5FoLpaz7XA8dm5ZaXFXQNvAX38zRiqKahpxlurCjpOnjaEgc
chuL62Tc8elq3iJaFC+tAqOzzVh1eSAs05aVgV87G6ATeK6UEnzj53ysls3V
8x36MygBLFhLzKuhXTEcizW8OZCVrEx978vWFaSzRgWQ+kXtK1QDnqFaElJc
QyCdP1ENC6L5VVZKmgDVLdbq6VTJE26NEMRGiCCwV3/bpPjkntA7jMuGB3p1
g2D0VkqC3dkD2W+2mXyQau1THT+YN/hhRqG90NuQBw9WXPf/DBznHehfgqpq
OYKPxXZUZIEqGPwPTYrw1aOsg4GWS7UsZbbKUzWGP/NCqnLifNN1+on0wNQ9
A5ok8rMDeAbN1KGfP+tUGDhbNoQhj10IwrP8kcQqPW4//J8IBkqhA/jmIN7Z
ctgoM7zepSoCouEw2P0oLPV6nTfOAcdY2EB8A3cnZ88z/plyQ7355LBpPW4C
QNpOELbjEIwA2Zp57x4r+EAM+gjpTthJOwazkNIwHHMcCI/omzgxxx2RTDQg
XMV6wXMAVTqSBElXXROZGMEhqVaNJ1WogjJ9G1gxFXT2OLZnZEK/LARJmWQ3
oT3WpbPZCWueq9hpnufEzfpPST+o4ps9FD+iXh3oAl3Sk8POtwT6iHjubQ0U
mmLlnMifn7gCdSfmVaU2U6eV3t9hQoNqf+I5c/VZ4ebxomp/c8mfwIKY/DmK
Tz7Ok+lOKpOLrXOieZCAMhoem84/i4EWM0uyqTvZclyzeVIng1J+TEuvoAdu
RjBc7wKF4zFBwl6Pw/zGpoMpqPg4jOTtwXTjXWeNhzaWuSFurzaUzSeq4vjg
jtzo4VjY9+UhqfnR43HcPGDTRZxwZx4nA8Hu8+++ZWoPegl2BzFfNpuRjkCz
WSRNBuf565rF2NL2sVyLBHvCFCR+siDzLPStZTG6EBCDo32/ePh32vDctkne
OhuvM3pXgRyTaSJMoWEKCyjXRAJo5zgwgqrlli1WquWHEitj3GJIUvLo9yFk
3dJFeam5Zeutvi6Fi/1KuOpl9Ev1Neuyn/jYt79sUchNLkxvamFZhdfFr6Ps
XD7JsdJ9DLbXLv2biItT1YkRJx2GLQ6XjZn6rRxbnz5CDRLYzTnj9dk6d0Lu
daA2s6TSBxo4COYGcGfuJuc+LIEFEO4/ZaVaqXtfpZOxBI+IE5yzgkE/dChp
AJer9i9q+Y/UtFQ1kuLC7EI/D5e/vMmSP8B33HLOsKBWmbhp5D9pnt4DY9jC
/v8T7dxSk7RV758S7u4G2zf6QIi3HIn6KbKhpmRsjzQ0y0VAAuj6+WzFeS0R
YN0/thuxcnx57EUcl4ooRCUbmF7Ow+SxLXnMtkOzUMrlzlbyBTGWFakYHAVY
tyiSeWai7NFwNmv5ActJpvtsX7OdmMwfmABU2YtTf0d3n+86UEVteaWssh9i
XM9w+7m8CEu2yoI7YHVE+02zbyOTtyBfPJxSD/uRjA6rx0EdeIO3ZOpeoKS0
dxppT3jxsq1wHM/FyXbma2Gl+4UCbYUXiZP/3ntloixWCaptFIztNrs8dlBy
pJTQyOiLhcDGbvrlCWH8AMrgnysWSTVKg2RZHSNm3o8qVfIiqwzsdAvBpfkI
h81WSXE8dEoOZ1FzPmVpnyWLYKvIKyfFOSJrl6L1J20raYLUOTGdqZFQe3HJ
heYQ9tTSRIkyHq88f1O4q1BqE2gu7MP6Bkde6+1qUiMHKL2razyB3Pr/2DCP
qsU8UxiTKpJcITQisZGuugHHH39b2bFYV2cRh6j0pv7UiQekDohzL++UAyem
7AvMFORzI0z0G/GQwcjdRzlpjOiPYw3wiCD+U7f5wSS8rr2DfRbHvl4Cqv5y
Z1/H/czbvHeX8P5T6p+73cdutj5iQHM3/jtZE5hTDumZtf0+HYJkwvq1qlPZ
5v5pK2X9C/vd5gr/C7REjE5yqHO4cwxa7B3DCJpS8XL9U4LRc30a6kT8GtiA
Lc1RDNh3PX41bH2sGm/QkwqZzBdgcdb6F0Rs90jxtxPXMWGT4Y9giPBMpZ7M
VA/zBiCRIf0HZlnHqYtYvE2uZFQ7EEUPJ50D1RLNbYvkz9ftIPxvBcaIaq+3
O9r1TCU2sXik48hnlue6L6T43oYiuTGNyyZ1ewzCgFJxlgpaJvOT6LuL/C1J
sWoUUNnxAqTNMB1LseXaAfdRr4itVp4nxhf+XC6qfVSd1hoYRqjF930/AR7R
f1T9zMTixUpPvQJE8pPqKgFwsKMHdXB4a4qkCdeWXhOxAweUGgfsVXlybRjY
waZhqyRoHI+BjS5yRvmkL2rfWU6Ftb+SxZey2StoFbMEI+yb04JqK84rmLX4
45ZtwLAnfJtaUMYyMLJiLk4RdCTsB1M1/ElSOUobaSHgLK1uhQl4igHB+8z8
67WKQEgrBXzRE9MGlKQophwV8pGHHpYzWpmka1mH0cDGyxcHDO6aOMqOZClR
O606ShlqgDsqNoeRFGI+aTHeCipbC7KBJ2P+IQHiU68ewsuEn5LylPVD9A2H
cZFXyOiMUJZl9vlyCIXlCMGOGpA7Uqwtx2gGvPexE/AnoleZfi4EyAimatsN
yAK2K57lQCjmyP6HCq58sEoc3/CyiHjpCwAS7avrTWnJ4aDdgmO0x+vXVX3b
rC5iqOC0hwdXDE/JHJ+2wV9gApKPy4Il8dOyDJLYKNW0pRy1rDTpRHrAtDJj
BiSi3X5wRMtgNhFMjbBOjkErk4JE1KWhbFgb/9HXphReC9nmX3BZLxu7hheP
7sry+TX/DWrzKQttecvMfxYquE+IZosh0o8LdZO9cZUz55ZEUx9MJdPrtYT1
P41SAoz8dEJZqPGDEd0//xSOtdLO1JGt4shkdNdodsQhDggJ3mpdVBg4khsf
p9g/1T/OdusrZCrSn+sHBg09nJwb+ttkSL49s36WgMLw2f12EBEQ4xTLK/NI
+VzMACEXralXhGthJJqDInC19LzLCiKwdxKg595gpYx9yIyFtN9ZfQvtu2JQ
TaVYSud+RX3yEpvQJT5czcjh6NGC+uzvsJhodU1B01cp/9XZpfiZAoF9zjtD
w4t7bfNaZhYLaDi49u9HCwg1jXSDtIQ6aqvh3dOM1iVjeDzM3qSiXl9Pj1DO
z6LKeiKUFfsifTXD+P/4I0GR7B83M9wygefQZ/fliqTYT7BkbxXtemnl6wzv
/lHvyEaIoZQD2D3asZZK7+93dDEUb0MraPWZJvZ+/XkXhYYcP1vF3Kd4jB1L
WDdw3xcOijxZcUQVON12p6XxRzMJh6l0rlS1/vevsx2MTUn5hvAnZBzTbSdJ
ueK+h4p08qORVYpa3mcDqNQjcYkaPz2zOP64VTOD+JPbxogwv+3Z1nTa4Zyu
bS64DtB0SU9EcV0dx5FdOAfxOck3VaiEYl7qtyqgo7qOnyumXKkhboSJclKX
re6aroZ34P2AbBS7R/RkKVFOHWkuj+c6fU76SR+RMzvgTfUG8koYqhWXeyjB
AfeW1FarKXuEruXq4TWYFP6BGXlaymySQDFr7zzGzXxWkyn5X0E3mTtbZnfp
n8X9qARja0D1fDoP0pfSmWkgOWx0L1SRJCG57RIV/3u/qeAqnt7H6+GY2wn1
YbTXSrPjnJlfZKhqb4hmfbisVS7ESh3VSVVew2an74EMPN1rkzNVbyCtgSZV
i+qE8ZUTWIFO9x8yGRNjclqwkwU6o/LxQxCQtjaxdgZMN+9HHPmORUoa1EjJ
dz7QQdP8Rjpk4hf4O1G3qFmcxiC2IZCT0GamNxi8wZ02w7ORCAZfXEXIumzD
15896ZyQZLsi9X9hMlEuoeWWomcT/UT1QhCyRgpoVEOcRKLHHjcGdZqN2QM1
Sl9L7g8m/4q3WTVxMy2h5lAFJxZhUawYC8OUpraxuIORL3x88P0P9IKYFfSZ
NkZ2rNGP9aPzqq5uXniUZ6628RRSb5PGJKIoXPuq4WqwtNHpQtLp3Qz//rW4
AyBT4jwbpCZaSddfxo/GbpWK7dvv4Mj9oq0jGwRd3arBpm9BepVVy4e3OzaC
ZDyztqQvh+eSdASz5/szNt+KW4N8DvIbD0ria+Ac8ZhQa4cmtTqugvUgF3EI
by6rX4fGrZebYJSC+hU7C4HFKyiFqtMTc5L2C9VAkudGscEvBWRqrmTv4MlK
yRu1WnwUnZEJmRxU+Q8TtPm9aDVkryi7Ylwii+RS6HiCiK8BQrAFoWuRlF4z
neGHJ+GAb0N3EzCI6CKCTPTlF16GUGOPXw0yrRr/A5O6g9XUJbazhofyyABo
QeKwkHTCDqoduPf7/EYsyjaGVVnYiX2LiE1L8hHgIs/Pf2qe+jqTN4bSOMRs
Mx3ED8GbSG8wSFUHKEpOuGTwi96iKtoHfD42kjnnQKVe74tHSVktWV40Npn4
xD2dknQa+WuQjLhmllcGErjPMeRNSRcdGELTR7a1OPK/Zh5rtmZXo8d/pPcv
P0tiwi2Fs8+Zni+yC6JXrhKI4bRj0Plm8kFI3P4uraSgXrrp4sEqAmKXp+tT
9mFbzVHXbLxRkvVgY4bm8I1w8zBSY8gVheZxmT4LeDaBfQy1HOpuMvEG7hS1
iguokS5G6AuaPCPZBDmlKarj35e2I6g54sFMRXfGA0pD4Ijdd4hwMwUpFXCZ
UX0SZ7HvBYT6TPS9rJICgtN6IZRNGLrZpr5GALEpUtJvwMICtao1Ktf6JN4d
pgBQIYjRxq0QrNOHhn5PwMWD/z39wvO4S2sZF9HDK/d97oRn/JpjLmJRIAbH
Ot4m+VUVnhtoVSjYfv/uaRvutjYPNlFckvYXyqI+NKeFSs80VC2L/foCenLj
zUPvv4n1zCX232jICo//o3A29cXbUpStMR+EkfE4DBhzJTvZKcOKsXlsSOVn
7hzCwRRDIpcEMffkR5Mz28QWB0BNFmrfBP0fsMoXiYB6XXAz/jRbcaRb81BD
JKvybGIXOEzj1+bZ9NTvSS6JzULj9354/chj+YaWRz+pUHFK75k3SSIuZYVK
+MaRKvc8lzABRSGuX4rZwHSNHzltGXJ7PskuGA61swfnrJXQSaKa77S+PYED
JfUQ9XD05woHtGgjgtzJX6efNiP2JsB5KIV+2wqWE035Mu7dqczFSyZPTbXh
Xq7x4M0QXVMHao9nn+hN0VahF9MXViobUAhcA3a2FeyYGY3U9vzTQ5pOy272
xbrVBu0AAY10dJKI5drMaAmRwLK2eii4s4lUuwAgyww9rJ1/mZeRW12Uc1EM
t/QTZycPVLPCIWwWH7gaNS9rmeNudAtMjZpiaK9Ug5J4+W1UITJg3EgiW6T4
o9KJakdrmyRKtyVXA0nicZTg3X+f54SJHlO4wiYSko7GFx1F8hR6Y+z/O+cs
Jk1ebwLHZkCUCse6yh57jtUxK44B2Oj7y/GZtA25X8O2FVjvHqGQlaH2y4KZ
DollIwU9r5txs+EpWnTFweDwmdVOgyB3YuhfLE6e3IoGGx56SCL4x+goNNB1
iR1+wEMrhj9VnZioY1PWwGWIMi/vy7fGANVosxD1Z/fhK8oYuYF0WvayYfBU
XMoTb24i5X3sK6VXog/Ejh5OtF8D3jtP+dAi9SO7M8a6WXJwpjkZ9L4hUhOz
WkgGFbYWashB0wWbbO9hd584suCeSWQuI4hGgqrWzhMqfKcovKx0mH9rcBYp
M0otCrOZX9HrID29d5mCyb8EmcRJ0BRD5u+LDXJN7et2q0Nk5i9ENvRZmBjQ
aNJerASyCsNDEGHWV8VzCgqDn7KsQNRcj4D4Xppzwdmdvis0LxYU3SXyZnhu
kRYGzNxQxGvxEXGoKRkIxQy8fM8X6ptmP+5YEGS6vwAZBtIcgP78WAjEZnlX
brwdboIWtqW8OZNRub108Nyqofvh+BZSDp1ql7m0wC8/HC8eksP8/RrwhELB
hPWpnr2zJxStZ2W9crlf0ncBlvCoTV+hh90+82oWeEXbI74cltfPnP+M0jSi
eklI0IXTggU2Ceie+CPm9vBbGriHS1u8F0UeL6uyxIoti7YSvXDCsP6xP86M
lqB7jvirY0kiYymnP6FNZoYnn4JyHqJWrvkYuDhbdmEtUoIz+wuk1Rgm/xCO
3ibVDBV3oA9+SR/ZZ+X6iB4Mxk8pjiEYxmWsFbAwJwtlt6+OWPsr38BLSZV/
0jcgI62c4GNcGQYJA4D6MkHL+T4h6zt7zlnMavPF89AlZIeBmOm6/Y6ICSwr
3jnUfXPKj216h7an0Be26JzQwbcqeKDBNFbnPEP0fIBqw4QoH+1uobXLCktR
woTMX3r86ZC+OOFkn4KB4WDMKYcxclJhCHlGD8coPXP033jLSCBq7am8p2gJ
lYw2eTj/1Oi4dA3ryl9q4Kbt9qjcxKoQCBRMTC5wasQy+v2/tGKDgddlpQMD
3tP2G80yoH0N2oWyQ7VfBcyr8bo8MD7ZwSkrDlCd7RfghNjVurxxCOIEdeRo
F8VAEYJM8ksPqv+OgLumgvncB/qk2oRe+3KvbiJp6aqzf7oAlf1lA1hHS467
o9Nk9egCisECAtymMuBsRPFxrZLRvMRnWHLdlMFEQyOeSnzodKNtKPcqykKv
sEKXJkzGiVw8Ytk06F39xYo0xNlTXMAn7kBmw3ycsj5tZ34yGpMFeCM851ux
4cdOLSV9nVtJfi4pAuXGkbyRgGJtz+mbZ61aCn97hICAQ2IKe4SIVOhO9zyg
pPYuK9bXdDE1RgMDxo7MhRA34s7btWw5uAs2ZPkFMGZnidKXyudZd4MvEvfo
iWVI1YSXJFXVhzJ8UlAsbPTeJUDdf2F/9DuX9gsaFIlQMW3lEROq2V3N85Yv
kH5AZRhOHyY9BqIRo9Nn66i/jwEWh0ulDaDSlo/ZT4lDBXwrLuB5jt1stBh8
YPjDFdZPaPcMATy2foK+h9OR0SNoUq/rHC9S5DSghPMA+xeX2IudmVUxPLVn
ljclglS8KC1GQ9jz/aXWoY8us1NDk2Tth5JQ9h02o+p5ASMrX3ePUUJSZcX6
eU0SfXvcpSBQ0/ahK1nZKRdKmV9UHU2/iLfL4Z6JreMmGUaQn1i9T4rsVJ3N
kupdEBwPF6mM4cqQca45K8pn355etrPAh94p3li32fUfamWGMnsxPe8Xfydf
Xtz7TbrrTOMbCWnl489G3Jt/JVxb2TKl9LPy7G30xuxfup22Kgz0PDifCLr/
zHXyRzsvknL8ECNZfYFcl1O2/3dg5vgx0MUV0TZiShSiw27xxoA5pds24W37
IkoLTsxByGRX4iAL0BxzWT8APNh9kNIv7WwiYgGYrxgZbiZGiK2aRwrKGKXO
oSbPT7tRGXbf82Qse9A1LRTsIySHftF0moBKWPnlqwneud+fqi0zxSnY9zU+
vNJh/XwDWYjJ8y5yYwq4N1rlkWWk8bTpLV6PDeqgUdPdIssvLW7qOSwCMvHq
pf3Ptp/oyqd0cdlV76wOi1l/brfllxA6NJwyl7eOLflXeZrBO8QmTn3YqHiU
GRE+JxtYipU4Wh6DOEDvdWISukEfPkUie7vfsqXR53JIof+oHKPQqXfeqgAV
gBwkLY3X14abLxGE1Qmr8afgxmEZjITnqgobUPsYxWS5MpLAxGVS/5lSiHUK
1qWtaRWmWRAkmYUDBI3Dp8vNLJb/to8gjPaibgdVvNzW23ePAAtJweWoU0dy
3Xv/aI8sLuz7e1nztrinvEKJCCQIt63BOZUbKcyHPC4F9PCayaFT6UXkBn3q
QOPYi84Z2ACVYP3ar0qJDY4J14hiXuRFkBEV/Y5cKioFyzMZMofn9cWVyob7
XEZzoV698CE+0vdlfPHFehpedPq/yKe8lPk3LsQZb4zlRsh3EFCoDnWu5ZkE
aUmeJ4ip45I1g9HAaBazoQKYEfy4UWcvh9gmkEhwE9t/GynSmryENL0qkzVO
Vu/0aSXbFmY3KA9XzRZWJ+dng0ic1M5NyGSBFVEEXcNUP5Zq1L33UkvbLbOk
pwpZl0FivpytMVLAGCBjMlKkeZ/6gv53VQxb4VwMbjOU5NpONxG38dCJyLfc
ygYYs+PN+XYyPpuauOwl/CGhudiVNbf9qce4euh+EL811lqV1fMbVeQoqgUu
0D5qi62erZ6BXZ/UFfTBnOO6J5HnAJgZeRUM84TwbtEjq0O+94Utz/loyYsI
VGKmdko6+VhT96jUTogHr1PuBYAAyRMXJx3OVqT8r/eGzXeYjyA/V6aVU3nE
ZjkVhtvhH5wFuleBnkh/gZZnURToc4t/E+XSOfOCO94ToOZUgv0cQh/ni5g7
Ic0ZtTIpTTfSKLA8d7GsNlx1CTpC9JVyp/xtrDXNNIHaahdg7MyOMnymIEhL
0ydby3ifX0uinZb8iLEHVNTOzYsZecDGQCwHmLNsJG3bsp0EcNeXY3kDWAgb
tIkBRw/TutDtRvshUGcl+KUybKMXBBC9dQmo1cRrc8lKSMbLVE/LlAwwWyFr
oo0UBDJksYrM7AxRfkH/+UmjYKwAePfoP+v2uhvwNdNybMpbS7kpxZ9RfwBa
6Ew/lpyG3BFovpT/2VXzlPvCXC+fwUTRBoKVdoE8CvHpBFPK4mgWw9xPCjsM
5JeHUxGXnzKLANvxmw9VRXSODCshZ0UUGNUh0tlAtR/TNy9IY16S+311SQS0
9Ewskij9fQXYju9uQqI2bStA7CbDXHzVI9ub8BextJ5C60uelv1L1L4Xv5o7
6YU5JxGFbihsxlm3pDxYaDAJY5FK3JkDSX1TU1FhHMTtfJFQVSebQIAHcx1C
zWgqehm6YVFe/rBzhmzX49QzfjeiA7LZHgFbUZag45uvHraI1X23Y/xJgAxa
sizqHF/8IAut+NErtoAJ23mw3f7/8M40XZ0W0RXT5LNkDmhspafxp4d5l/fa
pMxzNi0c+mz61iqHEcdI5Kds9gXJ2ri5vN7CMOQVOgUCzqyZaaVfsCI8CeV5
eqM5v7Bc0KIut5gAqtXgL2bOUNkue0v3qdS2s7W2CxIOKHF1rFplqZnGDWiY
a6RmAe1AWGBHjtEw8o3u8efVGUnw1gX5BKb5mCBSl2MSAcZ+/B1+nGZ6tH8j
ZoH8U8hHoj4ZJ6lS2nD0CvIUrDW69IZ7ZmBpevNUCDt8eE5NyrcMgI0JCU+L
DzE0SeGqg9NPE5XkY1ix1cniKjdi1SlxVnHW+5r73hRxx1YfA8p+K5iINZ6k
kkC9FvdTV8cecQb1G6PGg3tcGo4xQlYBRap7yCvvo/PTm4VWjsB4Vod0Aotw
ymdkKq2fdDBsiByEULZjcE+jv2KbpC4toLoEM2gId0BASp9WwA+d+bR5hSgJ
728UXPSbMwxH0DLcDQdpTIMmcNnu+UUcrvS1Ofk29kfZcHyqEDct9v33Gnd7
OImOlSPX9Kb88EXrqAdSA7Yuu04GKoCKyUlDz9QVwdaQC78MTFLu6GAuVtUJ
ixpZLwgWgmvAcwG7eY+NU3apC7RPpfUHLx8NHVzX3Hq1xo256D4rUBTQYTOo
utze3DmB+AGwUzrfAWf/UNZPlXLB5gIJVB4vWzWgI2Q6jbseO2jOuXnci3+Z
6xr0maH1KgHTaPPIcvFzGQvuly848tO3ycycuy6dC1uQo7kv2l/bHRpGvFGR
4bwWA1GdlsZs01EGJSxyQINFDCEf71nN0dxaVBNl4S5FvFSz+f0S2s2oumNt
QA9NJxRWUmHr1gYbiX9yUN/F+4RTZ5vCcG+uYP0XdsRUt1U5oIWAMMJ229jh
8feruqa2iXxCeWet+L85mpTjwlEumVdKyShrkZJmT4BOUxtnRmZ9irntosEm
/pOd+TRNB9wRwTm56nzp28e6WuXjRsXm/5TuhtUl0lHbR8jK5NOkLAslAv5y
jjKaR5S4JPGoa//xvAROgqd95O2Gynuy31+GG6sK7G9G3qAudbsPw7I0mmA3
cAXmRZ6FE7YUGMhD3Dhquh8nhML4oJvEHWqs8dAeuNcu9fv2RTPrQlOJ+ZGA
A0r1ajjWp9zvALjeR6Hii0MSDuTKLFUjQxubIjd1cik9+KvoQ6ZWDf9F6gVw
YL8lFZyX/QVRiLyceCs3v8Top4ePWLhX0zinkTpj+y0lLGFADIOkkjNCzr26
jxZbruv46P7fIIj7EKVUXzFc9nLYWyK4A32rnGWszEzW9ykquyEq1zh+dDiO
cF0Oi2tkUNXozc7FvFuQKoBQ0eXfum27WMVMOpgARklMRTQ3IhkvQbiROZJ0
aJ/n35GVQYr7C72C1TwgC68NkHND7QX+xaV45DxCk+zLiQy2GRQmPMCDtzZL
fG1WKtRY0xuY343MHHO3Gg80gFr4OlAMtGtdDSWr+fTZWzP8Uenwd02zU/y8
8Bfdb9TzPI3JJfZNnrpCc2bwPoqBDi136Pxmq0iunxALkDoA2AnNOukyLEpC
GnrIFnFm6fjbD/pD+Y9ztRsSsUPxnFr4Il3GI01HP1mtH1j/X8XFXGm+opqt
uTPNTV0jEuN/JrpoWOZ5wJM+J4pqbSGf6EQMAbcmN3YAiwB9mvs2hAVmCAjN
DoyWmrbcq39fcpNPmy6YNBKe9PZnsD3C0Y6cFINcBaszkXiCA/pyPRLjtv9E
uuf0ptnUI1zeW1DAfW/SQR6myaXA69bpOuPm10wgRKOcQ6HmEalplxF8WA0Z
1f+v5kj0LahVM/xzzCh6XnAuHghi7p5qs5S1jxEWrT4YTPLmdWwU1qODv9vm
JEpr/YT0ozj+RBcdjsl9ywgS6vknhhxqT6/zikCSX1d0PrPK9rPRDfpWUJXY
vhOMGhdNLaG1dEIgQvd4K289wVUinhvDkfCrJqietbHpqEt5S7D8CtRhWuLI
pmqULipK7EVwiQ1smtbAAFxjuKZ+nDr/uuMNZbb+96YeuT40e3Gwi5VT41iA
bS2/ioDHI9KsP4l4FKmHsiOKluC0FrRAclrI3jMkJsIA7OCoOrbccECIz9oS
dI2XSg+E9brxIncc+CnUSxFB3SU9NlXaiCwXRPrqm1b1ijekR3Cq08ydxTW8
kUMIFhNZp5/oeJZdh+qedlTz6tW08YnbhOYL5Vz/mjlKzeX1GSYXBvQ/WWuy
+FE0N/HMnWKCk0gYElMA+yabweqmOhYEpvTMPY1LhvMnotn6a2xVUAZH9RxE
+EiuaAx0z7Pj652QvxG5WVLR56IhvY7ztdMRgfRwCNmP+U5azLzdbGJqF4IK
hd06rOzHyohO3PKJ+ThyT/Ou8zlX2eKpqvyqxL572hnXw4ke70m2MGo8PxOr
1RDldh33jNKJEe+hGyPCGUEoDJruX2pymqen+ittZllJ69Q53ep96gJ5gh7E
4jkrlGqArKTPcY7jzmMNuTFfjOgbqNX9u9fQkA4pJHH5PgpeRo2WHwAPYK+X
43DyezrNyWIvd//naBePsAKRq6WMQLJQM47nWirbHoevDz0wULl28zqtKBxL
DOUIr6KyZEpRfxT+IhfgOrJ9Rv6yPErksHLPvjoWyEQ2cHFhJBmZzWCke2Vb
Xybgav85XZODHIBvAlWhv0QckQz2ntJStBsvw+U/Ff7xGJKu/d7p3YWg9X/g
2Q1Omxr3rzI9jjU+MnLXm4FBo1kUJPKDTTYN8LCqVj9G/M+GripHCDz6lR7k
UEGenF7xhFlJMDcPYji+G16sy6EXhkRCarKc3dYbCuL2cla9P5SOYI820d+P
TsYdVdYrOstGRSP/1ln2nEyNe8MpHEa8tt7WRQb4GaSsS2C6CizRJ1oEXxX3
90sfTm07vJdBmT2nZ+5Op06paf82QvF3NQbw0e8QQSQT7/SHDuO0a0+sDZHw
xbFP6SyqujmBIuagn2XGCU2tj9AvlbNiEKtHlWhYZ350HDQBeqwbV8Ph0J+D
Mlf3C91WhkMdsI9eZuHyQk2YQABjQOX1EI4uHPu+7AB1XsyaSQzCXnEslGFV
qkBiEAMAVnJ6sgnJBqI0B+B6qL92GcRGmEa9OpIuDJQAeloaPstGo5rMA39z
EH77ANpHldzNdurqKyiDdkf+n1iqhPSCn0r2tYOFHTTA0vwaA6uEfnbLysiV
y3xjxnqLw3DDm2wzqthKog81dQkg8A8QqhNi1knTvfTNX9n7UfPl8immC+vk
SfODwmJb8jaMX3sHlVpJyvwrpuCU8WG6oyWxLhDJy8U2ZF6drh5Kyuw0ipFf
mxapWeW0czqdgjj17Gj+bVEUCN5ZvVEjKKwFtSpqsOPslDNRFdtqkUfeTDF9
J4CYliCqFyLo0AGYnUtjDa9ZjoMfP1oPnaTT/uBKP16n04/iUmNUUXrjFBFm
wyE7hMRBJHFF7l6V0QfaAVBh7mN1WsWCcA0MHuEsS/yHgSaRSz1Z3UET2oT0
aro+ydJ8dyXlOnlkpQQju+VJN0n+KQFIcAHrFdIjiR4SJ9dxnq6lLTkSFOpo
EPzsRNp3YyOudsR7JMRKKNrCLFP4Y566pR+nP++eIu6a80VGnlSe/JXnrn9E
AW5szwjMKlLMT2pO9KeSfqYNa+5PJnnxFlKlhUcDMwbNhWNUL5KXnbptZREz
AzFL4I8ZDj2l44VIHC8NeDdww5R0oYy+eHAu/8EbO0COL7//Yk6h9Obiqt8h
30FIcTxdDIxCkmoyjhmRFBwfHjpMg0gKYGQZLpVN3DELcEfP0u9Af3DZT53j
D57RaciYYLJbtkGBnxq93E803fxt1B+seNJtLjYY3PqI/w7i/6nnbl6aZt+4
JJXU6NoWWDLzMuzPkwYZXlM4Vs0ePSqEMiSWNoMIbTilRt3k5yofvtDES8/3
39Ld39xGzju7ilFLbA5bsEx3bpsR29xVbAhQf+8cZegJQiv/HkOZ2hoQyg3R
l451tPMNqHE6loQgF57fb75h80zYbggd4RFlTJePDeMcDffZH6LvJtVNL1JR
eVpI8Gkj+A7Pv5VdnB6h49KcpSIkPGn5R5V0e786gwi2Grt/opFI7SMnh6M2
jRr2bJoC7CKtN3Wnl3Tlw9apTzvM0Br8batk7PuFULCy+NiiV35OgrtrtSV7
uCkWgFkyuDhVbs5zxZajV0oZoFeMYNPgH2Qyq1SpM8ivXcaAaFRC9QKotP6Y
dMTcHql7fdBI0drKGimI9pHkxQzNwY+B3BAH/CB8BSFGUJpHT5qO56jcDjy6
jOc2qEJ38eaINZBS/SeWxwlNZbz0ukAANPIt/SxFl/x1APieNpCTTsOXjXew
pXnVfbfhEJZdBiI7J6Ig48lr6Xh4zf0+yEurMjDc/9l4pxR1ZUSCoXQAgxJF
8dTbEUDk3S6DjFHzNHIJ4fzKnEtX4HrOV2voS8g14ygGjUMJ7MZ87tCJwvB7
E6YAACMXT/+T9DKMwWoMPKomG+8pZZOmMPxcRYamAv93DWaN6LzTA5maCYUT
aRIWwdtyJpZeRJkiY6BLyKo6w2XABLWVFTM+I2++mR41io7eKV6o4zE4m4HC
cTmsSojRQJP14QGx9p9iGnC+0oisqo5yPJi1/ROazMDIqBT/CflCDdvhpSWw
htnhbCvwHPy3OmAydkWyyt5vU5NM9Qktyga5pmpcyAXOlJAQUNNFO5D22qLC
+vENCJKuxh5ILx0Q4cFWTxdJ43wFPW9d7LIeZ7Oxqx/pE0eUT58HQY4scIC7
mzVl0/b7aEGlvffhdJ1hp56XRlgHbYf7tZcltBdIQwalFgsY5ttpRZcM6Bcz
spuuZ6O53Dq+h9S8ULEvGCRT8fbWZWmUNf/4YzZT+8n0sc01RnFHG4YGikr1
9anHEu6hNRKr+QY6g9d0pxbAxOTTeThgyv+EEFd819SX7ERpgRgIR2fMLRjS
MywCac8b++wTAWu9N3lg1BVAPsSiEQt5IxHBDYiqbTg55t56ltDadxTrOlit
BQeMdxjmshVJGoqPOnFp20vloH0LAizLCSYoQEf/9EXGdrSW+Jpa5KKajwGT
vADhxTyTY9W4rox//riBBNyMg+b87x2EX34/5zDNga4pV4wqT2bHvVgy7C0K
ZeqHFK0guVAhk55L9fmWH+nZv7QAh5xYCllTYj0Goc1Nnr+ty9bVOq1J5q94
sW9MQDc440dwUskRC0F42KgsL0pcAOwqkQOpgZ/GaoJzQuoztdr0yFfSHNKc
hD1tg4HaMYbuJZWAGx+uQXBzR/HBhtgNN63YNSDQCLYSJiMigdLFx8tim5Zi
57igk10a68BwOTkr4BtBPuDCdF+vXDfPEUOT/+5oIlJ17ALMo8cg0QKs4AIB
kV54SyXUCCRiLvt58XlUuEAKrBuzC1po+tHX5UXpUfGvMJSJ+R/8yMLm2LEB
LJTxv5aLyvuL9Z9cWzVO9SGrkdU42R2g4+ExxuXqKx8p3WpEiONIC2T/2kL2
mr769/rdPFC+MPElRvr+lptfa/YKbXcHrYHJvpvGnrff4B5frLE6iOvXuM8a
ukAzE9m1yAW98RA4X+V+GWpEEIby4s5agDzUJbH1KIqU7f2IX79JhcRw7H8s
YmQ2DRGpPwJD+AvTgaZJPB6IvAmwbirX1ZcLNj/lx9eeZVvq6MPtfrBPodZg
fv4a9y529Ns8B+qfcx2edLpScEzRK70AqsW66Hhsrx5DBCfDlNN5dHu/L03I
S4SgKi36FaAjjGvS2V0pcny24pMaO7avKSXGhoValDKeNgY1nymds4F9+wXX
S6lXRZTglPzHLE9u4vhIQJtO9BEEs4E74aW8ThPW+d4EC4QZC/GseKhr7F/C
zzTUhfgPwMEApSZiGk+jQ3Ap1+tFvfzo0Hh9yLIktFCAEhDnxJwPv1UgveUf
x9ethxiD71mY/kmP7MqUH3+SkaAsqHcoSip/HE4UX/OhtCSgkRWFQmCBDYCJ
baNUWie1zmLXTtzOotiXjfMmR9YyDPinn/ZZHUlF6O2Q0wVNEXTU8Q28wmc8
bDVH1ZbU68X/sOgfs2KPK/IXsoDftYgpn69lCzeFhhF+UgaB7sXojTlX8KFr
2NqJ+18kI2wJKvoWQ1HJb2N2wd48hiqkn6x3v64EHmyNF0CfAvExhn/Sen1I
OCT/9AFPPoZ7R00xhB/Z1V+ZSM63D8l+sQCKcAZWWwLju94gDTmI+44uG+ES
270gZjFGba/zSKlfF0I01aQazzQGSKPH+DWcSUd9aubi4himLAv1dsz/eMls
DgK9Bz2S4v1RKBB+GHWPKAkyb9s6JTziwNix0dxizdcMw59oJz5+xIOHPZsH
B1DvoSBwKKyq+p1e+rP4i7diwCpN8SnEX3dOYG1Irne0/HqjNPPpQajZn9Fn
yDrSbvKeKkPzFTZeOzL8sb9ATZDtFqb/iss8WGvsCOOhnm10XS7kxl4y9Kxw
mcV5arDg+gW3UtoSghbixlN7r6KBe/G3Lc+O/6PEb/tXuuEGBk2FRs5b/kV9
IN5/Isy8M39yP73H1DhLMVJVjm4wtp/pwxL/YpBoMgsKZeLoz/3Jf3DT3gHs
xi/gEVu85dr8WuOHuEqvzBKT59cJe2VbC/qd4UulKoxJhrGHGxkfUaK4KZF7
LboZgX5MWGaOAoAN9varlF8TVfno6SRpqSvd3gejCw5gNt8Xo4jlp7jwGpf8
RpMBFDfOO3ocPhZle7hamev4YkQjtZzeL69xa0xMEpRau0HSeDRDBoMRyzMH
ha2FDv9uhv0s9oFHLbZr4hDnjATgFcO6OFDrqWKofpyuGjmYM5rSv6fV7qfl
ls7VJfKTAlFnru2ySZZp+CJ7B+VAu5e9872s8bbnrK0Zpjmtz+dpqjGXFjQc
IeCRaSt4rBdAA5doLzO+RrsJBa80YvLxgLiudIA0xUqyYE1UHY5nmqkBoCLt
x1XyTrqVRXhT9dZ/p8b6dL307P+4uZE0IfB9QAq0/Kg3zALn7gUU5CiBFNxK
WZdwNCUmAwB6qg9iwKzWkO6s2tbP93VqbyL7hViRSbjMxMKy+qHYiSHohcwJ
jRVt8hJl7X6J4b19LIAxK/iiniyrFHxoKOIHDJvSx1BkqOtvVQdjkJFiiALm
QiElPFALdzH+PNqSieddyzCXsc6j/1InI2Ho8fJI36KT2GlNYsWecjd1Fbk9
RRaRosoAo4szR362jBLZRC9ZO2tlO99YwTVLWlVqyP6CGF38llFuNftrP1cx
7wbaH5R+UNhY7tKq0taDm6U/OJhS0IMrC+MVPHEuEbSOMSYpnOJ5vukKp3u5
dR/kes5iLghMgn/ENC6IRw6Tv9iFISGLwPCkXkfnyrUY6+3ACH6A4Csg7w8+
2aMQGJnasK0YeoNbiRV1EknkioRI7D6YefhxarAR5GBwDAnnd6OEjwHw3KOK
DUAP3RhJ/ABjle4rOrHqGuYIYnxcFljAC+IhVbFear2oFJyhQQC9QZ73TJtC
zwUPnkJc3PUk0PiAQVjlpcb32KGy7occxHuR5mcEMS/Xukei+zpEWsmUKlVY
2SKjiWVZ/TVbHb7G6pNiS4nQTjjpKeulZ8S5eTfcBRez76A4XSqJXVRa1OOa
nLbtyu5/71iMJesGtuYr36CYYu+AEl1kIE/oKPbxWRIFDQBT5UMzHLsz/ya2
3pgAmuiPwTpF72YvprkqFYv3JL4PdJ/FpyDrnfTeC6QnPYOswtIGs/OdNyRT
+w9kU8JgQVPFiEJUjuI64moWIJOQWJrb+OwugKoyVTpmrrGrYyRTYgStLCwx
vtmcpFvJ+BnUl4P/dG8NkG4Rsr3I2eKpqRmZDQN95G3XQz+uvYB/eXS/53s1
IiBKK52281avcw+lcQridXpCLNvCgEuqfuikUk7cugq6ytAovWTyYrnwQ2aG
Rr2HQlDgLupF9JUVGQKsbWJoHVm2jPo5hgdDNCiBMTNjaN1LcFwhWf8L7LXn
KOVJf5UUVbTGfF7A3KKGNfznO5u20+M9kl84Wlt3tL/Ffwx6qO/1NYNcnZJW
1AHsc3XyFeoJ3yJIRU4RriGdAojCaBuzpukoJMT2HH5Hn1VTk0SW3Ifs+iwM
b8whJXJPG3gbyljXZMGKOL71y8Qs0x8ayuJvdHeBhB3cuXJTKaqKFAe7fFna
7N5EYAKjDwB98ksYdJmHytyEnGRcWKOjrLo4w3LnLH2lVl6g33SPIlC4daQM
A8mluxwwvYrdbGi8OnDK6ZyauE1M+PpVVTn+9FNzigeBImEp2MX6lmTACMlD
5VM+K6CRu7GI7LP9iwQzyc5N25jv9SmCyN+icWYlbMddMzj8Lcg21yQaJXlO
KeXNlFQ5iRTBt/ghr2kJuTI3bOEpY42smZRphcUJtFnRdvWAE3QLAKMNOhHT
dW+sCk5VzniqBI2akocXb4BaBzKQeKBy6BMjNXxThFkN3wSXFn4E4+PsbcQN
uDyUeZ0Q+huEc/MNyu19SQuBoq+ndhebvaN+YPiMFXna+/suh4hJ6J83lWso
akXwAaMYbixBEoxjQgCXsXzYmSTrJEaHBbiQw6LOGAM82rjyZETEQMeyqV45
O/FVRA6zTLvntSPv3ydx20qXiOXf0mlxlpUIzLw1GciLV1+8U0lvSY3DM9Iu
b/EMMnigh1MNCgeVEd5FPx0SEnHBMA9vcKuFn8NODThr6Lntp+eAsfP/tHAx
KVp9mlc+F74Y0tXC9/pbWk2e+Rmc6DSl8rikLjsDspwLiS1sCdYBCMMmWoxS
9lXYbqy0Hg+lMy6GfodVm8cJIGmUvsCUxWT6rE3uUgURB4BcIfbEivuMpo9I
Nu+6YPWzfHubWYxUci4otMTXXeCleJgF+eKF/Tb8e+duzoEAqzElO0rCFasc
QkjUPZbG68K0f7NX4L1BRaYhKYquAPXYNR+KSvRfHP8eHKW/N8KKkoBWCPCo
ZsbsrFq4yseMcUDwwOTiWSawVQJbVrG2hA92/cbTMXTZ3Ajv0TqChVCKrMfC
KtyEQgDTwsy1NHavlgZc3/Bd4PQK+noiWfBmXp1KYWlMMEyR5sPmfNVHaaxt
BsCn2M9HxQoTOMXvEVY8ZvarlAeeC1pYWs0qMxA8T+gs6KLJK/QIbGBd+99i
0KNXSBKScXJ6BVpcvskZOJ+/C5sJYFdIZ8NuABzm6My9vqWPLmc3H6QZvkGH
ba5S5Q7gvSdMLn5fxcFlh+GMeekA8dv0RZGfaOU03If2k1FvN441CC/8zEWJ
4KZ9mQ1LI8Un0YmN15Wi6KUBhqg7s3i8EgjTuzH/jLKURA0i/2s31d/AoHyy
QVroWumjh7Ds89suG+zdzSfBnv1CCyIL+DXITBhnTJHlfS/bJfNYrtdLs8fA
GWDEeLXHhpPFcqU+pyRyKD3rmVI5Qvrc9nQuEH3nm1k0UavFU+aIHuPlWCah
Q2S7yJEKHSXbTbKRJdK75cADsDQpm0rNGbzYCp1Ygd/acXsvIXHY/oU0KUyC
MKysu96jhZng1KnT7U3o8W9QH34pjxYE7/RpMgwLj9iXNqNSoKBR2xJe+8HL
xLibEGjhs8/H92GEHdsTZxXPKvtcqsJZhpeax59fKOv3DLovZe1j1A3oFrug
Ve0cbnjh8JJhuJev6VQ9N4d+Q+CBl9pXyp91fS/KysQObqBc941g/S/THhzk
KNDsRKm6tjB0n9k5mWsSo4kxnSKn6Impi6xAg78He+zaSYyz6H53ONkgNPpm
cT6XIwYXzF9aMLW7tVarjCesoPrBZU4ja2mCda5uYH5+NCBrC+5JddG0T7H5
O6aK0Pe/Jf/CHxwq36hjNGU0neLCxulBq5idG7+zxcz9VNOzV4EUGv1wUuB3
tlgC6Q5fTcghnDiBTtx9M6kVGQFbEVRr9fTXozlxoTgvQsszMHu8jHAuIjdc
BTQ4z1FlAa1Ekv9PlfDUj6MXSh+wP2gAYFBfiBFo90EZyo32dMx0X4grHzQI
CTRrIC3GGBhUemU6A9qjjw9LjsfaSYYelvP6mk5KS9479s0jNvlHugCIeA5W
ajsYe2qUpes5U5A2kthYxVfkghnILljIBtp40UcWpF0O0xW5Tz+D3hMWD9ys
hkyoqQ6wRX0mfYhTaoBSvrbhormSB3xytBjvosnehJC3sZW1ebav7mRPl9UU
FZpWj4Zw5SFSDcuKAdHS0rOR8Brev1wjsQdrGYWkKmZcKcAFP75gUFErGyt0
BWrmOSm4BIOmRlTHHtYKy7c/uMjIIyceyz8WDW761n90Fzuj4v2TRvacBzf8
0PKh6f0RZYuqrj01FCHAaAcEJs/UC480yHuFcSIEU30xqfj/Ji26Y4CG7do3
g47I76waGKg0sXlaiYFmDNwY+Ra3y7upZMCgUpT1pvTu6OVFnD5d5f+Jc9kn
9TjY5k6+FuFQZPV9rSHODJmlT2dJIqwXBTFsE5xHsu2sQf/+o1KkKVkDFF+c
ayXGIjND8vMEJrKVk1F7XjGDVCzhESpedqErtYybPyHkBBiH/3UUQl31ysZH
mVOlLYO5mcQDh+a1ORriaebbydtT9w4mPDR2WpCYe7OF0FGVpyrBAO4tke7p
X6BwYXKUELlRXXfALk07CvUB7Csq165W7b22WToIQIi66dqo5vxV1oEW/BSh
Vx41hiTwQJATVkNhPtJUCyuPCYxybGFXnzgzRoVFpZxyck9/3kSMxXH+9kVR
BuZgdfNLRqpAaNHStjgRbrNH7I5Jd/aCyFyvSyj1OzkSHBk45DCe4urbevXX
tdhrdZ4Dfe2kZ4uA2BE7oOel0A36rcmJFsf5YOyV84CbXbru03hh1lz0p0Em
cBan2CvOFxa9Cr0G/iUiXrWVpFjc0dTJU2XOlRaPRuabwroNz7J8ymGHNmnI
5dbRDqnSaKnOmnAZERmZbw+og9p1wdWGYFx8mY7NqAM1tc6wmHI34p3LpMJL
tQLJksNA/u4kA6BfmS8v8O5SkVVp2ToN1moIRdTdaDvUjnWmjlg9aytZFpJl
HmELRWGw6LhId8DlG0sXKCckDTgLkLhpRIx7I1QVrYpnU0DUvsGdpxM6ctwP
BIH1pSDvfyZ8foIdCZGCGm9dd0gknBaI1aG6jNScqq0vnHKLg8RpQjhDcIZC
U94/IqZHsW1vKVXowYbWF5Dn7id1B3DeMCEwzkr2iZ6YkSFCVvQzfMNOrJ6c
pSylSnp25U8iCCwwKC9uw9OfGWB1AjQVn4kO4QlDaOzCGkH70hkLmaUxu6GY
64jiKAyxEiauRBpVJJ0VhROtnNalfcSbKwcK96+drxsyvegJfEc0IhppKGb0
+vJ6oV+rkylY9lUoDxGr58p+zXbgKds3C5YfB9SKw181FLvKJDGPLILW6BIF
SqdB2++rrC/WnMAq+jT966HvRyUH3XWLfMGhP0ftzkdLLge9pGLZaplsfe8J
GVczRbQx+uYqVVvJoAkhHyLlGGSiyRJjWpQb3+SGCjzPjAPJeL7kufNU/CWv
i9UyGHfFu/WeTz6NzQ9UlUH9eEUECMBktIe2DexUKcTMMDk+6n3v++5XNJg8
fI/lhR8lmjhbXHfFCduWMr12zdTBuzsWo2I2OZuTe02F0yg3DJ0vVkoc6sCz
ixijBjTIFBWESgbnU2tXfpmbhEd8576myTlAxJ5ppldwvdiRN7QKX6PWLman
Ud26UDKPkb0Pu2YqMGc9lCZzyNZy6/k3HYJ4A239fSVde986mm09lN6g+jQ0
4g4xJCQ6XiRgylwAZ+KsRbry2CpTtSWNtBXrJHAl5q9SwWWKUHIVdd57BIYr
VMAlcmgqxMOz2zlPBNgW9X+L/eamRxYyJP46iTebkr1QTyYsI6CF9aaFinqc
HfKsbB3q49Nws5y9bcWosgplrdYE60ytlCVWLLA2REB2SrW5RGcmu56ZqGAV
Lm5DH98xk7r+RSTV6xrfOKjyx0LcyKFLh6pKuTWnn6z0SjJQdMkQGAkTFzJY
sgL8YEElluihQLwpT18l9EbFnjWl5CQWUMYyrLnnno+4p3GrrcAgKGO6A2Gf
rq9zl4qGZOUVq6S9zBR+u5iHUDpQsLQm21oXJzn5nG+Xlohcnzdw1B06zUqg
XKefSpvJ/47WRWfNpDRE3SHGwGxnikMGvDuuLnC0rbBjXLowKCkHow4do0Xp
6I+kGwYORrKQM/aCFHwQHo/q+DoaY3mAqVbNjgQTm1+rqSA5ZIk1E363D6su
ZNxaeFBJlYz7QorgPATAWp7w1gqYJ2cjmMTH/OgGH6XHshMmPI93xNNcvBsh
4tYnTXVrnIeAZ5Rd8QbCQru9y3JtLDeym97V/OJKMJ5MdrY36Y6eJHTOpfaN
VdRoIz+IdZy1ui1O1QP4pCc87cplaGGKfCLBwTTBRN8+wOVEY3FHAVwCIqsD
xXwOotBndi7Ekvfik2/50pg6QsORobe9gQ9e5BhYlNzoUV8qxcUUGwi3q6Pw
8+rGX62p92nlbnGMtpgPOrfKbRtdJvhLbUYKba4nvXGPzL+9RUeVCOosOX+b
C7q6wXaWGgwdiGwibGQddmT1L1ihGJQfWGF6hbfr1CE1KVczUBKj0mt5rheK
s+pV1DS4pVacaiJUrDDfAf3vK0dBgS/aIbnh/roP/0vyigX9YXbZaQNe/8ev
8s7HrwrCnOKqx2QxiV7BEMGMDZLvk0WUp0V1wsjowVjZRG27b78dgYbSYift
clmK9nIZ/jAtffV3zRh0ae+PFJfTQpRm8xopsHm/v4jGZq2lp5BzAe+0nh/c
duh+U2NAbiwx+ripH5my4bV+bJqtwXui0Tl+rjqiw66tqXdcxxWEnZuM1ayz
IN/rpxbOkYn0Hh176UN7YAvjKTXWzbcz5gL+TrwPleWgimf9J8cMcTENGVAt
T1IBHte7JRC56jjV2JnXUMZZtgm0E+r8R3waYOV2nDOr+vgyaCZ1/XppJRWR
tflzdPpEYQHdHgAQxTg/SMIbzf4pu2cGmaflXTVJJ0dgXA6zvAW9uOcxP/gV
9pU9TKApUOATNQHtBmHjMguknaz9OnGqHBxXx1tjMF8SQ8xNfOETxx4gcoNC
nLDv37y0jDAvr0VCN814C3fNqAB/BFBnb5DDbBakPNNWSJ+tNayh9/+i5K/P
Aar2y+a9QOuNuyMYTq7jA92CRL9WfgvxpyBKIC/C2A5lA5ShcSAnyBpmvsxX
4EDXjjGtC7A5jl23z2IApizllylMic37bcqR/vFB5Id3WAAFAnTuL70t3URa
/AnJqCNcyrukHpUPX0HIV5oeFU+H+H9ChobR6TYuOggqQM6F1o9K7OfN06xR
l0DHDOpYR5QQ9B2JnaEUHWgCOdGiDU13nlbydDGVtepSeqphiZukqZoLSXih
ygUjy17w95m7rpOfQN9mlTcVEzIyZ0H+oNER8HNDKwYDNTxbtMDCSJ4rZsyf
RWNvmwc0QjTcJF8BGB4j7tcCkX3Efe4zRHmKYFd57OFaLcrpqDio2UF632uw
pum+QDQ7TewqVtq1y0v8vzkVjpa7lhtxKwUfkIaO/UCb4scWx4wIAGDks0sv
JjxAA/Yxwe9hcv5rAhlHelou5VKYjOdehu7bYRz7UBBWCBuN/U5EMxABXgNE
1g1m/q2RhPMZ84sBmHdtXSExFsmZmrYsSQLLoCnQn91t9cG8fU8iieWsIPs/
nIgUDi2DEfKfP/tkTDU6sccLcpCvCHQPSL647bbTh8oV0tnhqGknqtdsJNPP
RQ22mPWfkvzqMkeA8toEzEgL+ctEBps7SHkNZFHbaTol5Vdm9ieAdSSgyIfw
H+c3ZVvdLAaLBorSYVDFcUJuKg/m7YW16MGoSeJrK+TJgFvzoxQSsd3TXZTl
v4iF1X4s/voMZxZyevdw+dN/lWzsTM3l2I6LKLHoiyolnk9u4Po0OzIhp0Av
JVARCFgIz1ucpYCRpJNgzss80D7AyJaBJFnBr0n9zxqNLQVZoYgqZ4fHE4t8
JaM7JR5gbSCHwe4mv5Gz0wwIZeEU2VYSasA5zKgcgQIMV/EMl7fx7IIWaxHS
eyIqsZO/D5GzYOERZzQCjO6DfHPYF3zqiPxr4+xt0ZebOmg89zFha5znuuYk
RT4MCZKIfrVToLQyEqLdJscDhES2yCBBUwJAsU5ki6YYEh4ejhVAe+wfCSut
OE5jWfgD+Ry2YsHspooMrs5XWRfmypCWpk8OzKLbTlX210JMWB92sKmS9wbO
bK9QPUtPVkmYUOOFdS6trGprg6S3CYq+3eLy3gfRbnh/9HlbGI4njuslk7YF
QbV39ZjzJTG8cVl8b3fnaJdUTcHNdJm6DYN/qJ32luYvru5v37fTYGcIoqvB
yIWYnMb8tpyCUUh3WRfsTOK6zGgn/RrDUv5H2/Ai9AbHT1XMa/Tmx6xmbYZW
X/VUUfeGDqq2idd2NGd7UKOJXBdKUoOsbxp9ApMpDfzJb71uYFrF0YS2ysgU
zfPE3WAZ+imKxodmWPHRUMPJT3yGE7f/DD9b9QOPqs+69JyZsTda0ep7loV3
Ij8VwuIhsmK0RJAKY2nK3wfLSudm4aB5zv0tURUUrPXQWGEsqb9B/tZ0n3IV
Xsw9LBEudETNjYkE8w7+xSaRPEhBuXeSC1j8meh3iVShhRNg5gCCk6R0NXDv
DdoGrOaEHQBLe3cMUX2uAc665QCD8RtJC1OsdIRS82pVewkZR9hzK8OSTUyv
sBVYmuD+AIHsFfgDP1rmhEa3TkKviDPccRWqcZxuDWEf74XXuuOsSoEjMrlB
4ZdXfhLxj4RKoU5CFPSyMkrQ6WHgapLh0iIR8VhMQe9E/IzVOGEaSnp6Itvp
VHy61z/EZ7KPiPMOPfYESt8K0CPi1jva6E0qbEErF/XVBLS+MNY40Jkht9D5
k7lpCLlbfBgh06H0UugilMJ825hxxiAMrt8EjMZqtUgLTWQjb1PG1UX7QYUB
Q3Iuvh5PwbaQr0G9ta1wPzQU7nFt5UWJYFHLdbVsfPKK3zPqyNV14j5bzyyl
0UkiWC/r0CFEIy0WdP/PEpVKuqxcVxIa9aL16r1L7/paiYoSEI0rf5C8ciuS
t9Pu33UbDYNvXgldUVbmO/66KC7UVZGYBAzCV9O5JGA48SZIxwqaD5PSeR2L
JNYFjsgp0lTZrohoEfMO2XWefZiT9mBYjWefTYoGHVg8VG4/p9PdZfnKNb9+
KZ7TcMH8AkjweTtmIk5/RoEWxjLapEw6JPEYvcLMBphWSGrjeRNyzdSnoDuN
phjpKfNcpzfDWTFMYXzo+m/6MyCafJeg2kDSbFUu7kmfzlcchN1+TMsuC/xm
HhJmDsnwfzdz796FPBXBBjczSHvZnwm6gUrtswbxyZY8HiLpDdEhOkkfGxE8
ChLH/x2efwI3ZYfLfo4xdkNudNyicZuGk5FqXWG5o13vK8pYj73tjl1ay+2a
ylSoodIyTBlR4xGF5YStvxBsZ8ihvk+N4c5lXK7CBESd2IPLp7C1lQnF8tHV
MxLnvNj3JIaVoO+vW6KK6rUv5r9G00RJqsx9LPi8UKkNJE9Fq3yQYG1y2wZt
pW4CcnF007xDVXgcjqLpyRpcHDP/c4nBNiFEIDB/OqRYZXq4wOwlvhp7vGP9
v1vlFS92UZBjE34g6r9E2CZh9xybRniFsGlWJjgsMcsiw6u3RM81j6qM2ipD
wUvnV2Wjd0+9yrxQfK/T6+ekZlf5XiH2LEn9SmsNQt4Oulao1PRpqoOtZXNo
kxznaIlMAnJ6bl19spC+FgS5zsooozxh5AhcVvbz65BWSx4QZLXrvKmgff5Q
8j3UjkkRKTSKsGA+AZC/mZ6MfuFrXpmt4k56ZVEFCiGSxzZ3PoHu27Ha1/BA
oe1bayGWM1Qk4cFG3TdwbavUrpp2LeQPkZ5Hzi6vOXdITEXi9Aw7/Q2T6wV9
8GoPbj4OX8VH2m+F8TGGg/W5RnOQQ/+PBiWg/BbqsC14qZVAxJ6QYDCGYIMu
ODvIQ8X6NP9a0821C1cXpdR8lD1MOBtk/cjPJfnQNNimcGRx75ABwdU3cC7c
qQAj6JK+9gyICMRXwsAH1cVLhKYl0EAtpnXd6RQyiu73beeIz9qimgsWA3fd
o/fU9ktk8fygaX6wUW7SAZMrPvbfsauXS2Loeh11RQqWpwbEWWGnYNgI5FIt
G8VpUyyV+2YfOzF6IsFzXvFyVbJJFWn/zrNd1Ak+o6MOFEqAyMP1zEUH71fo
bp0IXOHS5Qkpp6u1ASjJRsOPVN1bsHgICgndLkhAZoiWA4LKrGYXYZQ8F8xS
7MGM33dVtxqUnGiQKbqtdNCPr1sikkh0ZMzbBu491dO7b6qky4+RfaFpnABt
+cxBx3axntdcRu/QHTqZtKjBveSVurwoKMrKMVSDIYBD226Jl57qGYFNFF2M
x+IzyHMPTvWFkdoIcobKJZL0IxPABGikB372Z3ZgllmvcYISfdrXrSOptH0A
QOUauglOCaJNt7ECOvnZPlFiJWs+yIxxjN/cgYqc/XZUkTtNkTrpgZ3s57XT
Ejrw3mFiaUbplMRYvjET0K8JBmmTX2fieDE0/NT8KmfqvmA/B5QsrrNEVKfA
Vhgep9uWcjQ9PU2sezz75eznN2cXpa7mijqPv+woWI2aFrKl+YoppU3BpxXf
S8hRoB8MyT1IlQYG/QevY4KTwMCcBrA6B0PyXbY8GinKlIIXCDrtDM+KGFXV
VOqLC4Mw9a20gtDcXqKnYO4RI+Q934AlVt2r/7hrGj1Oy8VMTfPclX6bdYQj
zaA8Xu71xf3/W+IspOutiVJwN6v30hzhPzBMikIGngPpcx+S/8y9bkenIkbk
WFhxl4WSNvNoxx9uI1bf4QmRRYBZPpCdcPjb9UxElFj18IX/0KirXE4tT155
cDFMc+01XV8p3u1k/e5TZwR9TnL9AXEI2WyKWWSwMRZIA4E0UBkchXk+h1bI
b9PrRUMznSsm3vQw1x3XpxQQ7CaNmsFy/PPUoqihapN0XUgybyIjkrRb651t
G0FJgAOQ+ogS4u8uApOt3H/3jFk7BP+wsHoFuBUzshKd1xaowKeltoNVSWCx
awq4BUOujTRXsJEAJpH3IhIDclwxbTiAYlIKfkDSlJReHw7GBByMSC234qvu
IbojRqJAt9ZgbJVtwIEd+ffqwYvrwPRF0mZKsdn0Ulxoy0PIV+WVBThimq52
Qt71dyhFNOUmkZiIbpEsntQsl/eAtDtDR9PrXOLP4GsQ05BXw3T5qDRMXFDU
xc4iMUAOrPDKes1E1KR7HYNaPZm6mFAeT27LRM6ysXpGhohwIPRq73B4T5XG
l512zjjT2+WH80xS29IyX4QY5Y6/CNscAVDRzQDpbcYrASL8sruUd4fkIJFW
E5/64eMBslVAYkQInDOFFf/8jiWSwNBn2KR4M4ZfJEmxVD7FlAmR2ootPdpJ
9KESSfx4ChEAYTKxhzY0Mm6TR7mV9s3CjxXeGcSS1D8fTVWkog790K474xR4
s8eahgD/GwjlWlGQBVj4kPGYZ8e322PjWE5CBCyN8vNPf8G0v/d5wlIOSbr8
Bk295RMdXxYzxACZwb9BhYvnVDAY8rSpOgEThGIImEP0eyv5gHxvHnqj6dgT
fp9wprTb8EXq33Tzu4pwsX3/8+6foEkmKu+G11g5asJt0Rv5TPAeVCzpdrAH
OaQPEluK8TroowoeqhfdbUsUkRfI64gqZgUNWV8Y3JCL1wKiYNu+pYOQWxGf
lOJz0yOV0HEUveXM4TlPreKdlzBFF/qzG1Yi/VN6VUm9q8m2Q4+0sC2jCtFK
M4iNFXc4KUxt/HP54ljYsXFpsFnQpT/8+zgyi27dcD/y9VCdWlccfcQ+0oRK
aIvGZ8OWpfAgoXE/jv8S4OoLTQP9WOAi8jgNKIZiNN9oVTj0CW50/h2MoByq
kady1lw38I4mXNFQv15cGceGj556RkrTo9TKdKleeu+Kr6h4mfnuMzTP/PNn
4N5XEIQBKVOgKxXrP363hdFYq37RPl7Zq3fTGrQCzZakfBD/q/nwEpbYsX6x
WKNKyIGNcdGR9GmghCzbEFGXbHTifXTHQPcUWwdxWwipKfvMspExHZeFGzux
ngtvOydHfGTXnkI2ZcoKSbyMyuadT0juoKgnfLTJSEwQHLrprfuthHcC2+g0
IhOhHoy6YwfICCXPVCld3MzJ4CB9yU4kg+MrbJ2yIKvaY4+1mw1Y/VdDR9Kd
CJFgFYmjjQZy5Zl6VKJToL2q5tWDyFoeuvhiXwVRkf5LS8jcxUlrwSZrazzt
gN/opOIbNRzBJCVNyNeMCkI3LGmSOh/98wr3tKjC3UGNZV2vl8ffEQjfbGC6
sPLQsCT4/N7CeXbWoHU7HAWTC9etb/+h9KNMc04abfXH9EZV7DL9QOhZ9mYE
Kk4aPFNwphRPb0IVQ5fRQKX1ylzZU8FQTYeuwNvytZcFzggl5ODir0mPaK6a
JPcCbKEC++0n1vjWrG5FEPwEJ2T+BXdjvV0L+1+R+OiyB7Bm6t7RWYh3d8lp
T7IAPF5D2RAo07hoDK7gATt9qDkmy0TcmR7KNWydZ3uRRoXEjy1Wj0yDkjoj
ajsYhXNgHTvsc3Z6MZfh4J3MKmcX71MhR/XviMgKWr+IH3x1rsPuafg5nEFk
pdZMSQagVTgt8FZz++vJD/6RWKxXOjpnBkh+XCLBx8u0PTDwvypBCzT/uY1v
8PSSuLE0kNmFivNehXOAeHKZLUEVO9h8WI8xMT864IZopZycwsIdtHCeL08s
ztNzWQGBOS69ZYOTf4Y0pJuDsY9MrG3D6J0WYtXAGWVTR8AcKE89FMrBOQaz
zYQ3B6AMKT5+ZWa1LM27gaeOpTZ9gLT2Qzeh//d+brD9sfwDES1zBZq/ATTI
EjC4YzY9ISSeHOZQK6atWNv7XSiT7u2Wxn5loDMMMTkg2KOdUEHIGhJfpmBK
FTL/YXMTxrwNMDzMcwtu7eT/phxz4wchVMYVCKgIdwqh19lVNj4J+FhBDdn0
n2MHqOSdqZpwt/RdVdzQaUjka1SRg/HbG2HgeLAO72V0BsPiQGmqeCGjvm1E
U+GzVq999NBuzdRJuJYlx6Ncotv6XfiUB0VIg2E9ygJOGow8F/ZzbPPy0HnW
oKkkb+CZpqmawTdnYPGwH5aY9+dVkQ8fzhF6zwS8z70nVf4SJVoQtfn3olJj
C2Y6QD8mFavwVXcvGcMszGKsO+WMG5D6dmpfonOtu6KQjdFV3tFqKsG9kJSu
Y+56g5eXqtkblZekWeFn0f1R3uvDd4cRiInYF+hRipjtFyRLD2a0bzFpZjxU
DZmP6FyejdKKC6wk1cTQlcRO+M1UfpXlUL7K7GENRCcklja40QRf6mBF0e40
FH9hC8gGlbeOCrcUsAZt6KdVd7iAKyCRKGIxmms/YfZyQqax/4J8tRWKPiCN
t0RLyqx9/GnIjjMGdQ0t7ZGMo5GkzoL73zDSVLv/NEG+YF+ia0Z4u6bFf24u
lFpUGCGS9ibfAntCi4ktWWw0/wT+L2etbeMXtoXEyQit4Jmeo3XD5SN9gk7+
sn3f9MuouEdiUMiAIYeDYHkLXNAYVF6Sb/3RnsSZkOiYlY3vLcSwnszRJmp2
ZIHQrD1rw8fByKU4cLHvBn/TrDGVkrw4WdNnPvF08URytqb22CQwS43nLiBe
x07wSfU6v5rpmmNyjs7SN4/14OwOPR8VOhirpjDpkT5rmRJzL6NBnX4bCBgX
OC43sLuOqafI84DikKbUb/N9dA90XBM+dzbku6/0KC7jYxXsEacTZa3qtyrA
zs3z66oBk3VRD3ESxyJetsYyi2X206pzuiLDLolEowmi+ohoxrjW0xvx2ieS
tBJXxmBKJpqMsQOZGN8/d1ENmdT7FRcZpwlVR68I1c5naB8QqoyZVGaqNiSV
To23xEQxCYXv+TgR1CQtAy6VjwWAUzkaFLj9CZFGtMWZWQ8+LLiM/NuiwnTr
iQsOcAcHVn9OMqOox06SRpA/k1GTYNSVoYKuj8LPDyI6c70+QhXXKPX9QkQT
uqdpp4kFKiEj7b4xkP/H7MuWEIzJGsAUZy8ceiJxNWVEXjv855K/69Dl+6OF
bN6RIaXSKE1AaHsi8OwhOBf+6HyC+tOnvjYmbkp+jZ+YYA0bVq2p5erFMynv
xmeYBxevl7wpwehaLB6FVZoesapPdSJV6tkoAgULD85QjX5ctn/YrxJsjLfe
LppZAOg9A61LXXdclNeGz42fzW4W4MCngFbjJcY04JBSd78HluNYOZl4HPkB
T2oksVqhrkr1W41JN2PLpWr0fhZTJZzrW9nju5ReoBWK3QPa2Mdw7gwXNE2C
r4S+2L6vfhrnvjQLHoePO+QnPfZpxguIl9/Eq1/81tO4l81DUxyt6LzZPlVU
8FlofIp1wYRxuqYEEmSnv44Yb02LO1HvPJvFht9BthwHQE2FqRzkRurbX724
fKPZ/usEsr90M8v9A4H+Wl7TzR+Xju3RhOhYrb9XWTQrQdUTHcjJmJLcvPxg
5bEIscxCIj9LKDCeTMRNp0/Ig7/SVGuAlWmhk5DeUNDNUBgHL+zH8sxmyATz
7/el4YuC3TXGVdWcfFcmFQli9r2QmZtV/mT0kgIk5rQ2wbrgigSjMsx9+ObI
/MT8ev6capSchrMVd/bvr/Wu29vrNpmkJdV6AtPFkgnrkJPKTG646ffCc9QU
7w6H2n6oMnWfuqXBl9YKo3ubc8ggfJt3hhtp0BcX9eTyZjJlfjtrlS1fg6/2
7qDLtpzm7U6+PubxLJt5GZMz9Zvhkh2DCFGcyOsT4VfJdVUvMGMX/U7ChBcp
347s6xEBmGlTxk2ebRlpGaHgEoMZlsh5whrf0gt25p3dSuodjuUO4+ETJRf6
8X2aQLA58NONWS7OhJbgo1zZttdwj+dFdqTGG8wjmFpFL6YeLic684IgdpPy
MWyZ79pJNzeYQyVYvOF0RSqxl7CVqWpWKV9y8TfXsPuXqUlrMCkCtnQmYhMG
TtBxV23aax163iMAj53ZhV0ZWAUpWYVcm9tQrMJz9ZcFupk/4Oe0QdeW8jIJ
YxWgn4iSHWHDYvmLxmwGi+D96JPm5fuQ2/01/wM6DKajV95Zw1SMoYu9HxvM
r422dQnRHv3VSwVzwuPYTTkVD31FyZ2xA6YVo+YYQxlrI+a4e5gXJZGwXHva
6qKHJTX98KogdZ8BjZf/wNA3mCVd1lOgvSXR4tZn1Nw83cFAuafsavfjZXJZ
WyoBRIrc5C918Xrhqef6QWGeFPn6d8xh7LHLGL+KLp/zNLaljJA0gOPehzAJ
FUfWdsGDqTwv+am8drEB3XFfQlMYDaZjMp92rJiQjGO+rmeOBtNwLFJnGanY
kR1HmDL9/mQPDO3uGWI8OWC+cMt9sOvLhsYwf/OIf4kKj/pfaEw6YIiA+eSU
SuaUjuRVYFutjZ6BtE/22l2NtG/TFop6Mwh109cxS973YKPNcFGj6Wal2xeT
SdO9jKZPKsd9Uf0TeddReitJWUDVk67GknmjEBusWrGeuZ0faRFdPKhgUGyP
4e5mblvjcgcdoIN8tpfXVK9L2yDpxeZF4ypF6Id2C028RYilVhNJLWWnV6eO
PkxMy8SxH32c2s6hdLpz0YSUo50FMRTJyNjqsYkcSuqGx3mIqX2rdcxmj+hO
SreWXKnXs6+X5E/9OnnuRaaVXgbg6gqrp3w6NbnNM8Gp1tm4oaaywBFs9/P7
OzLW4mrrH89goY+o/1A1WiIdoMbO5rgcJjWctPOmgdBtt0hQpQFXAIymeIvf
Yz7S5AlNeYaPbob5rjSWE2e/oGewRw6IpDt5cX/8WqRfKZwyp5l7Tsl8W/xd
dE04u8netq+aybuv9Z86OcvFa/8WnIqZ7quU58+q2CVUZX0oH8peFbys/lEu
09NM9xEsrQm7X8DZtLJpqpxGbiBNPsROk2ECmey8g85wpxQirxzD8d/kHCy5
XxM5trPepZS2issqKMtdcKYn/Ezet4eDiU+yfwNDiVyW8Y0A5SeZuHU4Eadv
kpYFFVPsTiRYPon2ScxY1rcQcv48/DED4325KvVLq87X+cGz6bc9ve7fnwJ3
61MBrm+sOzg4+gBLh3Hq+IX1koPKu5KiUCwU1CGBwXZR7eIYl2tXjZfxZBXJ
VGd9bJi1tGZCg15SpSqQIOoHLNLBWSefA1DZPhjS22b6+CwIe+iuOU2O/D/X
cRz16fPlavK6Bkzr/TRJI3KUc/ru3+nx+TXYCclDR8aiOkrQ8fHvGoZJt84w
GwpdM0Z3dNhqeDI6bvhWDVsSAhkyIFHvbzOLenMEW75zOKTB/7KdIAtRvi7G
AKiPTwsjKcb5KbFlsqM6YJpcdq8+rEqbFsMHYpRSrxq6u3n/+mAjl7LJ0Fnh
BJIKmnbmOGWmWhczEadI0vP/+JbD4wT6PyhA04zJhqkWj61LyyGJK10a38WV
KyFsQHMd+SCTCJijBZfEG34xobP4LnAX8nsPvLx2hGTzWTvXNShI9ZLu8A11
HcJQxb3u8hOylaj2PjtCvE7V4qkDoWdQWFs68CeE+QJxHh7xnuwER5aeGAB3
NfL8tKIO+h8dTA7Huv1olZrBd5wVkOd4wpFkiJ+yqvYT0qHmd8HqiY7LwMAe
VYKDrtDmDpgheeUnk2oIENuTk6XEXbzJXFJfKOwAnfLAIKiHS9md+rkc0H6l
Ey6WlYrtioz5RgtHlD+Hmph8Ful3sA446Mfu3tBlehuBqD6WyENGZpQEea8l
d2NqJte+r8sbqNu7JdyjDGHRKjG0ZrhO7CJTms+cA0iwfQTNobFjApxN2Ac0
LOODs4jVe0noZXmUWDCn/CQm6dCaRV5p0sydKxb0yhZ6jHS2MgyLRy+nppdF
3NaBdNc0m2DemHu3+wwlNzui8mr/2bsVte73Jm6MjE3zIfWl1V13UN8QQaPj
tLcGVZkXHwxWMyTMvqVzI8AeeGpPDsypj3Ukdax2g8vv6QojZ1udg37Ntds1
eoMwG1soie6rFvvKySj3jcBse7CCc1h/0aorJ46kMfnSa9OKcQ9K+11K3LCv
x3nupvrMtCfNtdA8/jcnO/R0+tVEawuDY3qL7FJSz8Lkh1eOZJSpan1o4tZp
0KTk7uWte/giZhBDptkfbRCdNXq3xV5LcY3KEJs7DvIqTzb5k2hVbPtCSOB3
RIK59TsRJILEY3U22MQb05jGlmYH4VVeQ6ixSTqC455IJYEBI2IfK8q+A6bm
fWH6jsYlfC+Kh2wpA4nLuyhGyYNSkbjQUKR5DDTyzdQxP1d6kpHC2tNNXVGO
M0zT+3Neclr3mLkwVD+tHkP2fv1iCJikdhyxwiEve9FFHK/5OWyMg5I+8Mcw
kCJS/YLecrkQadmZe/M0A9i+4OdJP+jeu9Pz8BNrWawW3hHI27QNDXldJCDe
WzQbRf351B329XfzCUrt2N1ZX9tNvxhtWHDqvoxlfidUEC/SL/SsR2jM5Wpx
3FSaCpzFqTB/7Ohk6x82z5Uia+01urXhFecWXMhGSPI/dXStMb+0xruTP2D7
58EGHjdlk73+jmkmaKSCS+Tf0Pg2Gtem/ipiYmAVRL8WeYY1DzscBvFxMAYU
88PUePmGGDty5Opx0KOcXIIQKsl8059ZYY0OmzZ5+Okew0P2DnOvY8DopbkH
ym+o3qxYZkRFlSCLgrIKIzK+DrYGCMgJFxvwXAFl5XdQvSCCQxiIwKo8K2xJ
IsEqBrkANTZi9Un0A30XukwWSwd19tju8ojobXqiVBqmkhaylWj+/R0Kcbyh
n18ocULEidcNPeyDHbRl5cZ7/j+BmkS5XVoDOjM/XNbmnZA9DajJhY2DRh6I
BQwRozQwpiEile6PIQdIjgmZTJo4dt1lO1uZLuMAHSmThKozvZe7GKm74kOM
/6GYKp37ZEDMHrRZtapXuvEGtCOsnEBF1neCCWHc0YXkapVDuU1sJ98Z0JHx
0j0Zo1AyCVdDw3mUWK8v71C3RNrAk+NQ94MqWb6dmFCfPXhXZ6HbUf7uwh9l
XJoBxId7aD0ooVWErYzHGua3TG6SkWYWKCFxO0YUuE1KEjBwgzJhA1GP1PXd
2NwzHcgtVlsmYoEKd+QLH5lyIbVbHM/yEQ+JHY3eOP9ktCA9NFRJWv1NeSPg
d3Rqq8toQ+UVS9FRb9zFrgctmpI28JZSg3Ex4wznPph1uScEs4fK5wvSwrEC
e3ZhbrsFU8AmnaIU1x1/KCn0PTDZ6HCj1AAcy4NXTVVXFe5XxJiEp82hWuOz
XZl28L0Uc/8uHDmaTEvzMyHSgosWV5lDbPZW5YTWc2K5GqzUUsy1VHiYQcXS
rFL0eDEl1KIaLdyQzt8393chG8XQCCXKqhP+1fnpedeK4lOC1CkSfIklk/mD
Rw39cM+wc2831Q80ICX5hldmYDCfKQvsfWMIWUW8x5/MyVv9Y/TyeB4jb4xY
7+mUmXk+rirvi5ea1RxBNwldWcqXARi69YHMpV2bChIwwPLOVrm25cmUu4yh
MXAul/Ar3Cow86vj4lkxnWWZXFGnLoDhFhIGl/NgKcpUiWZLhitWpw0DAh6E
/Giq3SnB+Ju0RhhOJOHqKilNZ9ouyoI3zvVd0sdJEPZLWcI8mMJ62QPRXdD/
KJJakuWR7ta/zdKxkai3aCUGq1btH3a2gJ45P5YicyQm8k1GzmZ/vO7vbI5/
NvHzKNvHZ3az3Azp7bkbx9YBS45JNXA5slFaW680hBMDfeGXuSebDFlMgox9
D4CBjkOF6Tyi0d7gS52x+og+CM3UhhPSJIAGO6gDyIl0b4XGlszXXh/X8prz
AGeZuD5qxuMX+9Tuw+xycQ3xiqKcxmGeZf9IMS4+83qwlJ6jk5R1N19XNcSc
7mBB/60JrpMpWeqxbEV4qzF+FqGzd7bJBW0qO6TD90oifKkOPftVidF6r0pw
jtZyAjWIhC1GotveWkohm3BDlIvd8KDkuL4Sly+A2Fs3zadzlEo2E9euTppE
CeuakyUi9Ayjlt36049yJoueVcBQFEo7zUyB8l6m1SlSBSYo7LwfPSDDhS6H
2FnzmBBW9VPfFU04Ni0bReEs7BYbc9WPaAHvbtTIgiryvYVbnRCAwuOplxWH
kiatcNzu3lA+bOMh6MI+JuIXX+ORPlF6n2zwLOAlXgkIS52dUd058KERU91S
YCQm7LP9gEkjbbpTbXceXOKtb6bIOE3RXO+z4YuJOKBaL04TwhZirlvr3HVJ
0Q94Z2aXWifJeo1fesX2BCCi8abe6iSNayEHdZhR9kfMch36EbM3gnHKCAgL
3ccYy+1yl/zNMbKq5+5DkvwrpgKEnFgWMp7P3MZ3wAeCfdT7xGR7HnQxVTWQ
r19hf25hHOQZTZzjSUj2DqlafZTG68pckf6OzYnj+OD89fzNlD8eTa3r5/Xh
0cSoUapMDrJkHdkdqzA3O7EbGmm97EmPNh9DzoxtC/wl7Q7Xur/Lq/jRqWjR
+H3bPaBTBEiJPU0bC68uucKH5DDqou9ah0VTX7eVqbfBZF++tvPzolGciKU9
vECD0O415MuH7k5V2nYz8uOfViyx8lJ1r5bi0kaU2RGy5Rt9YVtgtRNciS5r
5ZaZzSHjIp1vpCCq3BAYsvgL85SNBkfhrq+gCndm5U2Hxeuznw2J4crxiqZi
TZf/3L21c0l3/u0hic2Diuq/ktdHktfoPLZBqbTceduqKbTlsnUEO3/vVGLg
wwAZ007ZA4LYUqx125CxsQgKx+9fZXcoN1Icw7EtYtcd9Us2jPupUVL20Rvd
vW47PkE4yUW9WGHSUymKBpPI3grAPNkMpNDh5fYEAaR8VyVHTu0Ze8kuhdhT
0NeIhUF15B97iue74ghSys5a1aBYLfVwwIwi6i46/7sjfNccnQvcK3yeLo+I
OWu9mY1VwK0t/pYIUu7rgj0bRj5mJazq+6QC3/LBReFUqFu5G0ANHsr2K/p8
TlwE/MFSK8BGl0+f+cvZwBV1u5MSBQeaNh+/rbtORKode0R0xWBGviwh0ZUD
hwOTUeM9Vb7pC6rhgRujZ/aR0v/yD6f3hZMOr+aB4+1mCrgasky+E65Jv8o5
CR/Tqj25Ugawh3MZmPC7RisHqNVbHrDvqMmrzvASQVofITgtn4UDdX67GUGx
BrY0wgM3arNqBofLEBqeRJwy/yY+dPro2393xIdQCMHLLZU+QDeNNlDIkHAP
MDuvhkXG4an9Vmo1JBMIIU6qF6SsdcSMYMpYGN1yqBEklO8HQZtTE2m19rHZ
y8Tt3AfMfZqErKpRSmps0LkXsxviakKAjc7cqNxYS9AjRI71fLdd9G50he4q
aZC2KLSuuBKIVsTmF//AmyCZz93P+/IxJDp3BzbgqWNYpaw7feNzJgJKtTvl
XczAhiRJWbE+1as0pGJ4ym+Ma/poEkINRgXEWMxDhGHoM7kprsYNu5jQM3b4
PDOL9OVv4bKi7jeybz1nNcEZpBP1WzIF/njfgvDIvKO9n87YePJCSQ1nH+At
wKkbHTeux+R36LFjJ8d5cXLW235oVXJDIxe8dfYRVq48LEyEsqOYAu2mMWmV
PwuK3UnC5SY871pMsbo8uh53TNNu8jiqGBxYBza+rJB/+pSRcyO/mF7of/o4
/PBWU0HDSFGHrMrAmijkIAm2ajvJsj3vMCkrjI/SvYIE8juT97P2+D9Auz9p
XrQTSvpE0gHy7zx/bwWIvDg3AkZtg38W79Znfuhks9sYNMsQBRdzgsjd5L3h
4gn6l8hdSSQ+z2Dsz35lm08tuLVymlJcx8ayW3G/dzRaF+gfJ1DcIHFZTuqz
zjnBL8vHAlv2g1J/bFd5c9XNmiYWA3ut7awrKvQp+eDLLAXVqSXpToYZMRn8
sXreBbbQeRrjSJIcvLaFOX/Sgw9wDOlrhcAIwoFf00+rCsIf/MM5sv6/HLnn
bbbgHziZj0j65J8ilm4o9YngUkz69Fy84scFf0hfWsZGrMQfSRrJaZ6XV4R/
482VDDzXRWEMehpWMYUuT6s34CQ0gz7iv5k5DskBfKJ66VJBXNop4mpJahOh
rPLkW1iRQWjkxUb9cjekeLorALrJCvlFGz5AGZY6UJmTs0dgfVHwXfMOGfTH
kj4RIYGOFWVsE4Z23yBGeTh40J95JmMbJbjCBMTwpcwrvYT8z2avZ+KsIsPS
0tpbwymkQkqxPvxBLrh86B1YPXgN8KR0EWGREDjl6Pr0d2l/oPM1omufkjE8
HBRhDIS3F1rAXPUFdZX5vTWhi9yswWtmNSfYA4zziKICiR9o6Ly4pTu9UuvL
3oeVXPzAPzxoXhpb5IyyZ/MjpWews2qxHUIpGLKUpACb3vJl2rrFPxzXUgvs
otVWGyUDS8GhZA1J6eo34Pwe6wkSh2CfPwIBaU211zXMncLURtzqMlpec7C+
fTQe23W/CxVtcXMePEZbrmJSa7CKK4cH5TiqPcPsa6GcIfKzWaovrM/YIZW4
+tOYpB7aLI0kZurrXnEtxWkUxrKy3oukcxjOgHGByf1V9kpwZYg7GGJZKeWk
i4tlUhRr0Tmz0kOluElQp8kgXTyKOHmQeYkw3FpNL2OAnPpEX+lqTXRZSkmm
XfadH43x8uTfyonoEj99KrEmWkbY+iOQ7rk5k8JpC2X5yR+fSUQvcAdMp8OK
dXb5hy/Kr4TutduceAfwJxi6dmF+Ozi2cFqUb9255epYq1vOE2SArYlwRlH/
dtYgLYi79xXmugWDF7T/ngf170EZ5y9UCN5sc7be+ILLP3CoF262xr3K4eni
szDOpdB0aolR5MVJxY7j+I/wX2Bdxpim+f67KoCjxZLfZd1l1TI69ne9acca
ce0tuAqdfLJTnjpcdp1FuktakCCG+UCnb9/Pigef/LOgBkC7+9R/QimwuA0i
DKGck/yvkoXqzyPooEGMXPozg10nTE+M1UGLrn66NYGWYmpFA25Lz6iM2+Wr
mZkfpGjDh9w+PBGodGHW8tyVFt7MSNm3P29RBZDY3iL7rTMshxPI6Qx5grdA
ohK0UHFPH/1f5/3ahY2LDtkQaywSVapsBzYgygeEQiVgfC3XSVmUub9jSaD8
41l4fF4kpMNAp0fS+9yIzRDJOthLzjbeBGj7fyRtmS3YKtUXj+FB3CPECxa+
SGrFp2thGuLKosCOCOxGbr9k93HoMyQps7rODWyXVBkH4+seI07ZZYUIh8Ru
xj+mj1HUlqyBw6yBRHXhfs6tKp4aOjc4OCahiReyYTBT6QkJ9Sow1mIcKVsL
nSK5yyIS/e8Pn6+1xBHj40/UUsuI2wMbbF6DfWFzX9GG80YHfAGsNKdDyPWE
x+bP/hCrGfcRBv8W79SxexMq+ZffJEDzDFXo5REVvQzFcYs0BUFJX7nOtnIQ
P6YwAuTa7tsKqNzwZD/26NubRHl6P2ZNRIFRfqsLTqgZW6ZxnpSaLzwe3hR3
xH4NVwTejsD7dlzczffp2/PJmgxd3X3fB8/I+Qgf9Ow9ZgHLXZ80dwhiGBnf
lRAKqzo+950gHVmyvvacqJS/wFUths+P/Au27G3w90vt2k+/yZcWICIgXIiq
YpAht4Ti1kNBH56yniFe+CQOxaf7mihYCQJ7tfEC1x/yY6r6bmwpW/KHln1z
l+Td7UMdDSG/v9dX/RmlqtAY/+QJNsaN/x5OjeUpZlyFWJ8CMKsDuKW1IwPS
Sug0P+ROK/Gu84F1YOFsjJG+ExstvQlaeesFfutcssQPKIAW5IYs40+ipjjH
4Qpz5pbgAYyxFdoXKNx2Ny2BtVHBoCMJu/v9F/UQIr27TJa4GWmqCUUuyMGP
eNoXYl3zqAUxzl3LDg23hj1DKcbsTCihgppY8uw9stOSFiZfCtKIon5kmWIk
Wgq05SIkDowkIrWzTcfK7MELHNM3r5DT8s5zYEt6tsWrdXVxi7qwmDDpHPWY
pxfo/39eiqpyyyOGiPF9Lc78wNsdpn9cXuoxGrhvlQgfbe+SoUpGIdrM4rOR
1/kTPGrDSZPNqZBCHc9bFFYFam0BaoywbG07WE1nmNkqXsx1PYoxEHKEgDoG
aSrA1FdkiVFUXE+LJMphYVGy4QvFxSKxQ25wBPg2DI3ul31pzGYtBU6nuTvK
N0WYYqtUaHi/2e2iLd890T6Ju5bJQnGSdG3KFJbeayDTCVDShLz/9ueybqbN
zfklBrjM4dPHmDMEIQ8HQLlfoqnkLLXuWsbdmxKXzo+gDGF16TP/8pN0XH78
4ZH2CVYKtrXrzH4p4HK9Z2MKyJkfENd+vSVIeEA2KEUBxJwejbz3b/aXUAoe
7w24KMNGUduC/lEu4b2q8JjlDug8BRKd3Di5rmThu5kc1E0WREEE1/pV1NNm
z1FWJ/cpNOdpuF4mIB3dfrrCiP1BgIZfHztFm+x+YAeYOwBV53luwDJlhUiz
Gy8FIEC7Eoek/kGdePoIAzQ3BGpGCO7TRBnYno1syMtxaQq6W1c/3nsd7BBA
KuZpEJsDV85EI9ydRUntJVc60iqT70SMKH0T+IQnIvXFUDQ9fOl0K5fl9g2o
nYSYwM6gzjnobx9OsmGPLePnEAKf2LfDKoIDFPSzMHC8jKaEZU5YinY6T5Wk
rKBYvPKLIU3vKBjVO2VutyHIT4NqSolZ2zrqk0OuVnoemdI04YWpq+64T5g5
1EtNqpW4I8bC+vRfYro4Rk4adzvZyLhC6EQpZWnGCC4mW31VhC/D2EipoAKo
PySWeKAw2+MbPb5mkbCGeKlze65uXLVzU37nsqOch7Kmz1rKKBf+68EdQIIx
chzO8DnXze79fJpva6XSRRcdhMrOl1yRQaSAvCYhrVXyKf+eweDT+3wZYr7d
AdAZ/JXlHcJoNqwRAISBAHxSd5forhIdDyeCZwlNO95ZsY4QF+0idant6iib
gRYS34OIdxQDFM/espTFDZsp+xws/ovUUcGwUr1XSf4VbmIEqyH0TLn/hUTL
tV32C58fj8zJM8uUqJOlTZlty05zrjLO2mgekPKa7XUyuEZH9Q9XoHbe8/RC
vLI06UsjHVhpywJVhR3WXI5Q6wS2zQOqsD1kz/MRW7leQXKrUE9iujqpfG3s
N1rzW9jOtmWLvIofvRf9T/+AMyoSkoFAJruODOXOCXNeMRBIZMM6HNQ1FSF1
ceDqyKyK2WBXlz1DEq7WIG3D9boFbhs99MH1nSWfbXfnnD2ZM1Kjy4lOCEOw
wMqm09i52eWxH7270To1TrJZQDAliP/HywGLJrW6TL7nbZVL/CMtUWV1wrTL
xJsj+v/Iul6S1QCVXXLsQhFdrXJmCy4cQFo9TwvTPOP4VoiZj6xDSeXSeU99
h4om/XFMjnMkiLF+23kkoBYk6+eXuQfM1pZjusZBPYzNPCkHB1hakPFCudJk
QDI0yBhSi5r7DB8iIgaHQCXLz9oxOubVYvkhgzYnEGHkdX7w3rln/SPNUJ1R
YSpIMLxw/LM9NkwyMCJWnSyBzgQqnDqFDhEFNUy0ZUbiJuv5shmw4sz5FccA
/hifSVoS5/xe72cOLdG2PCCdKC/Q14J5u+alJ1PqxSJ2pCClP+KBYJ5qDSVL
Xla9if613eb4iDMhxsKKknN+fIe2GxN8M998Ph0dz80CTTKn2zc09Z9y9fvl
6mgPD/ihFlMqX8cXrc+NBU/464OQeY1ZwrwUudwB/3KR1Q9vp9BkavQ7DHN+
DhTXY6rKmyVy8CSZeTPGNn1Co7a32pCu6hNEl9ak5jGpC6fBeJiS/aNjuem/
bd24eiUyraQDJjAJxkekzFUSiCn8cpPLXgjbnUsB5ujfDHW0qCBozo0FqhTq
yPj3eeqVs5+9Vq5J7D9X2PmTB4U2O293xvXlkCAtnmVW/Sd9NcHR0cqYIjeV
7RMnNfWM24QBXB4FhZC6wAm95iVhfiVxc1zPLnq04/X8K6Zz2EEdOHI7I2we
Ev+otCROLlIDNkA3CifJNvSgCi8h48nzJ8C4Oq0zUeIEXjqcfxDoXCPAhuzd
gxKHioJx0bw3uDrWBRcbynrO651uRCw+RrG6SokPssS1LF0jvefPtyn3kRwM
yvV3Sq0F0muT9iZB5rzIzbe02ZdPmyTfBLcOXRKPPJFd9+Lx55kSGVjRjfBA
Gc59GU52h7fg1yUOrzJ1fUcEbjzmsLpGBD1moZFZiUJ3c7VbEP1e+2f+mzWy
4XjPL1zmt/xH1duYprWxsoY2Pwrzxwcr36HqeaFQQrt+XP3KxxvTaj0zJXmz
1h7Kyhlkj+4/wuGS5bObO2fzR4OqlKUd9jO9XMaK/gHMlgnZqAIhb2CxJbET
c3UZebXRmj7KyNQzTWQ7KrbFX5u2S+VwO18NPLzZ0/fxJ4ZwONFJ+3B6qGqp
HygbLFrAENkBIXEbc54cJbJET2gkUN6PSrwAhvNh8rg+YAcG2/seCdmKAZex
x7ZXxvKe2pSIXvmnQ6zH9/wrZkRet38RJ5dzrJ3Ku+FtHXLO/IbMSvRwQqC9
roS7dbp5yM1r5uB1OTM9M1wvFkweeaw0NWPYDHXBKUwGr3qWSGDut1qRSh4E
JJMf+DgRkgacdrXRDZItvLlMED4+Kw9v83LpYt1G8CGiIVjSQoTGrmpSeglQ
dik/DaheITkX4UFzFWkOhxBnuPY+E+zybiK/gML00mUvaOdRsZHPiK1lDYxC
3EtnQ0l1/Bcp/okB2hxysu5rKqIYcYL2ypWf2VlqMmS5n2lUEDzi7hYuGfBy
jHozdPmr7M/s80NPGUTQ05oJVAQOhNj0YCIUdOJzjx0/FZMem9owomXV3ERK
vvrHTjpfeRMEqtLu1LfP2xVMbtaX0pku6739AHSgI1Z1atOkZEUNZTtv/g9h
NvEyThC4pOTTs4UePjEl1qqmo58vrcRkKvGaRejhExFPAtNlza0p4qUj09wK
ZJMVM9gCaZZve1eT8Lvfmd3SQqmZuLO+ztPoDjmQ7nRFlUY8Po4JPf7pKpyX
8Vv2WI40ljRt4Jl/VERw5i0AX3dPhkABuyvsTWr12kDcHjrflGteiCM2DC9Q
y7Tz1IeWvRHGujpO5h6AoGPmUTIJXBiczkHczWZz3ISTAkiLxGjJElzJY+44
nswmn+8ChXxs1nrxDFmXl2rfJE3Spfzr5BLf8e1iS+XB7Bo+00nxGxamg+vr
iTBb5IDHJ4Cz3NW5rDp+8H0W4YI7eyv6kB3LQJVwcFw1lyctUC1JRv0ykYhh
yGXukzTMLhw/jVE15H8qNBqu9taWfKearY8NyX/3e7r2vWXDcGdZ8W/4smQD
IXKG8BcBUyA1lH3F6oWiuNFU3fWHDemWgCmvdmw75H2ZQTea8JzW96jp9eUP
T6xNE4abb7Q4IrY2jaCtGfNkbCMMiEH4+PNVVHu8yoyn4ebUBG3rVlr9IGr7
pIvMListoEa/4W0v69lKjpztUoKfvwtjHktTqbrhIVkD2COVAEwlVHrKvUGZ
fg2JFgW7ddbj+FeBWR9tn+UsqonfvH+c1SClCTgCKHKo8UuD1NdxQGkv1lM4
Ew9Onoil76QScIDtlZ/V3WbnInlO6xeTaEgQgEA3hKh3WT1wrA6RBBu3h2Zc
Z8QZqUUZOCz3aNgYnRiURLAZjGXI+Z7lDRqfFoKsEpjrfaA+cflE6/kSLEaG
ykerGLQ6J76jRx3aPFSzXiI3MoAdaEfJFfx7FMEmkgHE31eK3KDvwaaYSsb2
EUwxqUdxuVmlXCi/UO+Kh97lenedI1+mNLvvNlTpcK3EF3yuRFbtrOBN47Zy
hmaR/60zLNOpDW3AePbi5Btdouv1VVmXZSWdNhXSlC5inI9h3XxUAgZTX8n5
A6Y1bEpHHSYB7hkZUOUsd31WWIRBSGunDUcZyLFj31xQTUR6/8egE+OqQ+1v
auTCHtqSHGRI6OMNsAg8UeibbVACxgJ2NIxLeNAkYW926aBQOUAFlfpGGqiG
ee2mu/DvO0rVpwoxjaRMAnjutVLOkyGa/K9sqTtX4G70tvFn6bZZTOs8O/bH
DcxSqdjTDBwxH9HaTscOgOioeigEBgfyxr3m/nbrkYuSyy2/4IaXJkIkpE1c
Q4tfYruCHRlpaSs+MtDpK7GehZNjPEHj9xAPoIAyTIQReewJTk8elPOvTA5n
jhYLdKe7EO8FId2MQvZ3vWo2NRvKsTJq2GqtljZFRSpiPqSuQ4cBSRfYC/iJ
Wf+6yXYD1WWtMvXL1thKXZ7hNkPZUYUCWMSgcG+IEPbm4/u9L+6ofFaElZer
K5Hge1Ch07Mf/bpAJ+R1F/yFfwNwVRvRV4OkmxUoqWzBe5gaQ1ZEgEHGUUVV
qEiSQdaZsL+1b70F+6znak1wIPD9WDspTGgorWUOLv7kyQGqGhCkzvQBsS8z
Ez+Bbll4DZcm3Ed+gQBTkC9+QNDjVZSxj6RPHBfWPUjH49DE6Z2YJhRtnL04
dLyW+7gktQdZgYldV7QB3E+IWOncYUDjWo3xEr58Ax+4HnLinXwpasW/boXo
zv+zMfXyHS/dPWpLpNW5cKyKMkhfMil74+EvRORVjBwWNUPzjwn1y2YETDFc
MDitHAgPU4G7dbVC539PThvwR1E5Jr0/DchAIC1WqnGBE35ZMODDH0HYdKR7
/gNov9nK58DTzJCB1m+PEgDlL7CO0zJU4F9j0KpG8nv5xz4tdcO+TDUwA1tW
aiyCIjss0M+0cTu1EeGakVtwzNR1s8W6XC2Y2/TJTfcyUARWLSf/cSTN5YV4
nPjT2lyR5XpZwSdsooiaE4eyVxuET6+rZ3EnP/pe9WE+xiHkVrQSY3JSwjdS
SyNa18xna6jCwgtXJnUXWiRYedcB5YxiwjSmKeLUKzvg0+hdEBgOJM1YAsRe
SIBqCgUSKGri263yRr5uT9A85mTqT4+AIF3S11nn/Rjpc9uUMCiy7/nItJTU
c3wVbgy5ktJZd293hKjFdQUNQAMMUrKb/jIhee6wL81ae6P34RKVBoJhrdI6
fgFNCAxmWnEINj08Dz7VqvULLfKI1wHxoZJOYMU/pHZK5kOrX5uA0xashqNI
cn2kM5nNZkRs9K7NUzue/RQAofulqPZQ5I4pOi390tNH7ce7mnn+2r8JwGVh
hCzggF0/YSPPmhAv3PW0qh+pw0Csmuz7WrVQtPk3u84u1VpPQr0HRXePbM0/
3/u3ybrUPmLoQofCYxNTGI+2AtxK/o8fI3MYArJGWK+2WlPf5yYXHI1FPGRD
BK3qWZPd9col2uarRqEz2IwY1UIwt9PmuFDlsVZxkYd+E3fHPpUkCRYvG0SR
65jzt9hNpvRjME3890EV8pC0IcqMSMxQFfHrQ16uXvS09tJhqBj6b+NNJBtO
9kk/WTTJKVCUaWp6Rfbl9ZvjLEnLOqok3Bg4ROzYjoT91JtkbM/6y+McUY8W
MvggXw1l9fUXYV9O16JsIf5NzCVlI3lTq+HFQMYN/MRx0H8BU+JA8POq3Pwp
5Ke8hme3Dz1e67kaZPjfi4qEuKw1n/9l/6ADaUNJZd5TKamyKSZCvAepmKLd
EbE2Kd2qUPYhZ7nLzhyRnXC7fw73uk1PpRAka2tP3RQkXTEfSmAxL/BV2ntL
ksBUuQQnfBZpusEQVWe7l8rYpCCv+kfiPcS846zFqwY/yK16ifNOZAuJ1bAj
g9YIeFn1XTj6QjL5WbfyPZ6n/jhk7qEE87juBEBn1nvc8tTCyAd3x4eDjc84
5hQwustIZhlHdQ6uawx10dm+y1AvojrXkxF3V2YpgiZ2PT+TS3Qq8ZGhPRjA
L/xKqG5GK7yy19lcXtV7JZ/mpHCssFRyKWa42bOhO7ENyyzkyh2nQhlHznWW
bU5hDzKXWEglg3yvch+Z89/Wzx3zi2G4VVqjCj1bBxzAvBCYpr92j7lpGLZd
ZPcb18d6d6MjpklHERhpK19auESDr9JMHfGAiSitqWzwALeF8DZ0Ouiw4jj4
Th6xM4a6p6x1osI4EOtVsTrK5KUBrAjW1mA1FwiCeOm6wC8a6TzRY5dhnbZk
YLzwxie7xDYtjnQ3b8PgckXOLBwpbd3m2wvg+9+AT0U1nGXXPdGpZ5ThKo9g
EfKP21vMKYviwWUW+L9votNLZriHWAaZCNGjIB8bwBVVGjlLDqSLBqMjqRt5
mnT+EyaQtWilnCdhvsGj/VxQzfGE/3KYIXLtnlwqTotFShWx/3/JdJFdzoXV
3G0gBNt3AQsq9X9sIqHu67UXrXoK5VpenUPFdI7yCd8rpqHdunYnzubywAdM
csThclSjcg02CYhVpuQNVZOQfVDSwUScORPmurqD2omfmhTDR2qPjTFaINew
JhSycduAs/3+B+2bRagBkr6m8xD9DCNJo5POdgOq+bQNhG1jcsxjPjL/1dZg
Ld/bQ8lLxqyNLoZ4dJEMcrFXqR/ukJnghze85q9kZwwdyG9wJDJYaUvlmG2N
ylIGXeLsJgkwiqr9dKb4lN1Gt9VTtmem1f8UNuhQ3LURgX8O/S1pLOD6fnJ4
jnXaJjZP8TWQxSExQo2u9m2sv0nt80d2o49GkIyFeRBdK1gYmQu0rPkbMjyl
8yRGicLZg2Iw/QPnvysIv+YsVEfx+Bupud2OuhY2X/L4vPKIxS3emQI57vh3
AuKqUIpcgmrOxjQmR4isV7N+RwO+u36z+ZJuXx+ck17oHTD4hLJ2FzsRX7zV
t4gLGaTiz4wKLn2pzm27mvqO4MVpM5ORWeSWgJUEC4IerZtoSzNTaOOFRZLK
+ct336SP9f9is4bXrJbkPtRSx0USD93/aghf4MmGslo101M3tXu8Bvx5lnwb
3R2oz2Mh3t7k5dK3T9lJnviCu/Q/OXDijqShq5Ae75sG+CcFvgqTpqo2hYqm
/LV6wA+4vxwpdF1tGSwJ6cZeNahMXdvZcLq26uJdmID1ZQRTZZvgBtdWXcb0
wmOOJlzzR3Y9Dd08CJxQNyyT//fCsHspTGdmj5T0vxdWtRft6aF6DRyTGaff
sEPFfJVmyQoc1pqQLTwr+uFCD+yOo3F6+AxYbFnUOu+qAsosB+NssVTtT/Gb
LawsyWZHtuS+I+5FdVm68p5AgYjEthAQ+RP6kR/2tnfmWb28jElg2MhQw8Gb
TJqx9BJMxIXXp+nFZrZtNMqkT+yH5yf82A/iAALXVApGbc6iyCdNq6ac+9Uv
Uc0rgQNI49OFH/CV6OOxDVHnr0W01vYO3HqOHmqBXoYAcudKEfecQMSvhVdV
/bNgvfONlwuamNgL/Kspi03xV26/lZghqcZGXYQ0bAxatXlTvSR91wLg7RNR
qeA4+GbnF20VoXBokHBbnzTzJtBku8qW8to30Z/r3UnvKzwJ+xYsuHtT8zSh
wRE2nTmBLGuxxEHtQ86RbKWy/mc1XrVYKlGXXZSMi4A9+TXxjUumlEA2xfAd
8LGZxqhUxP8azgqmz7/AfHjDo8dDMRvcfsG4q+JByJ66CgRA+5vCnRGlszMW
HKz/9rZXI2WYp41rWxOtCB2P/d3jElorXwVFA1PddWzz6qwddVR1xbGJts5G
1//TpOGUx2t+IHIGexLUiAnkToltFGRVJgmdegtB1gNQtIJ4j5mw0I7YMNRn
yEwQCwINhvIppappjPOkc5k7KiVYtO/Mj+Kfq0Q8FPzjAMNnCXdrp+1zK0Mj
81HXDPhneU1Pjei1UeDZYsneBCMBuJiNhZGfvPhKX6H5IV0V9qdmbvCf6XL3
faJKIhhwPKR+ZXGwEoyzop2BQxhs4EQ5vblBYphHfoyihuBirGBs3gjAF6CZ
ughKqW5iA57qEAFNTj5/nfgK7rZ58p7BZZ081N5mjxtQAQvQ5L74gMRnOXiq
WsBwTdTQT50kOT3+b2yGAfoOZkttWmhTh6cu1qHN/2ZHJWRUG29mT7rFKiy2
Lq0YbTi9hP4YlHbBhmhM/GPXuXjGVl9r+bjQ9q0HukxCRScpC1xUqSIqcEEO
02r+NYfnu24LGwwS6v3xgOI3MTkQ2/s5+pgYE9sKOxwlKwBn7XOcI/zl0p+X
gh3sfIK1t62bawJcm3MkTNaNlotofJZIwnp2vlzRdxGL0DEoDJStqi53uCv+
GszWmykOiXXwe6x2AQnW/LryVO8qI5OKNh94HLXg0IdB/UJfhWj/402CejJb
SPoqpU4U6aqPqQIUlPHftcu7VMxnU+fshUT8Lx9DfQZoNDovk5d5Zdca0vBM
0RXBiQPMaDCmwHkFwsqB3K5riZKebS35e5MRdTcs4GYv3GnpPpnqrSiPRNlv
Jz3Vl0e2roYIpKLNJeVp1nW4d5PJubqR7IuTPGFliE17pDfIp5n1Bufti11M
r6G+S1LC+ijGeUDugqOY9IHjzRSGMrgXTFHWCFKlvaV4AchJ8z72bjDWxtO9
ueB36CGUz93kKCqlzm4pcqMEzNYKOU6Lm/XRXG4Tyu1Tcs7XRedENT19J25I
WULGi1UYWM+tL0dHfuWXQXZSkPsq9lIb0JwA6Cnc2tUd/hUVlGOLL5svw0Wh
6SGdeAO1BjlTlI3ctVYXokebPb9xzzwwCIUK76n7BBPwv6xEi7n6HxunjS6X
1TF0ZLmkCGvZLq6cC2fPS0LN/dj/MN8BVl4YArX1B8HDW3eASYw8PaIgRuke
ZYaj4Gp8c8mmVqwE/VparALf+8NhEwLvC2C301Wj84Cevcf/uIv3vuTE+5Vl
+FEyo9xx49Fxdth/CQBL1GJyX/dTvXW3eeggH/jdT7LlZAihJ+MlsAv7h4aI
9JlbA1b/Xj8uOikkjrZIfhp+qnWQwrJru1QsOeJ4EQKdcKIbOB7AXLdo03DQ
s4lR7QryrGr2Y1p9CaPHcC/HSvhpnshoQIFAnNSQ0VB26mDxH/GjDY6dIf87
PfF1FY7XJ7BTv6Kwm6Icn6akibTjAUfNhNdtHFABcNdzm0rPfQ5mfdhzI7Sw
fjpMvvnZcoHeFpGj+2xPHGSSxviXgxhCyTRc3kNv5LKD22YiuqLFNp04A8ap
vTNr1ivRH+DdtdOzHQvvmD9il95nTF++Mv7mOIMLnKSul245p44Nmu4K7vJD
h4j4hkzym54dlFroD/z3TAyvaL/UepLQvQzDUQuUz8DjK5NQtwCujBqi87q2
JMldXKQEf8hOPUgeMVrnfqgjVNrCgSz1Oqy+wYoWceksdD+KUA6QdtDmm6S+
bMN9aVZ8T00ogl3SQSY1ZtYyMPzRhWzQs8yQbyQ8RlbI4r6p3OLnO1LrD9sv
fyXBd6vhC+YRlEMxCMDvBj/2erz+H2pFr+m4LRMw3s6bELXNHzFl6gfNjdAa
PDKB7B55R7leZREt2POJ2sfVeuyyivImJJwrUzW3JKFcBl7tDDGkSnOdpA1I
9z+LluEBeTjmbknPnUpAW4r+saJ1CgEE7LNYacL/67X9bHgL6Nlju7C3yEQc
kWmsoMVDjR77e2MUTNrvOI5rLk8SbUC+9l/HHkrgmeNQi5t1j/TzIwmATKH1
NcyKyRiMvuJ90dILXCtdlwOpcyZRG/79vYzVBfQTBqv5U7vp2UQYJtWgYJTR
ozzJnz+pJLmwlrLlHaAaK9OD6jCdWyJpEsKsiHtckJVIMKehQ+6vh0SGyN+1
SwOAn3VXflUaGEXf9Ciz9Wr+lqk4ULAMAXYbBDh+Q97Pf7li2McbEprkHnAo
6YVXAeAexYTHIqtnFMgbks/DtbxBnsf047vPg9kXGMNmPN5Q+5+zjXodSBLC
psWISiqc8j13a28SjjTW9xqvXWHyI4/FkA4jssarRx46XjfENiDZ87aeUBWC
Hywn10mg3Fs2G1lItJEVwxprfQazQLs89jvRVglWNVxIznb0P4Yjxkx690en
pSi+a6uAThtH0OC+gpypxJf6TGmHPlVrSE0q4PzwqCN7E4cQMu5Q+erR8ENL
xk2o3MV+JQy4YN1YXnXJQPSLUNt9ZQSplSo4DQaObUrT2hWxPa2lpc0ZTimm
ypTVjqUmdjxjdrpBEkQVq3FPZir5zdFpUrOjIaxLPq4b4SfEHpIYqstpPCrj
o+zTKlYag3mjC2YzOBlDSZkTammeqKMkb0vkAho8RIFpo6khK+OOpuSa93nB
7RjpFAOzdvfI4XnOUh8cGypEWLh9zLaQ8cwb9D0ICyRRfU2/mYdAsKt2B2Ww
KzWMd2rUr6cY7G55ZEBOKd+AwJMTand9+vGjXxNpgyPMPiDn+iPjIhXAG0cA
V9Z05KKg5m4QLSu3JXxrP0ce2bccNOLU9w7YS0/sOaHev9y51mdsQyGjGY4e
kV/2unYH74JK3zXXkxpgViGw3fa0je5fnJ9L87jOwprvwFrsSVOGSput0VZl
4hjjIbHhCc4MxRpsShfne9rE5gFXOOOyDrPwsjIiFZDN88kuMHnw2CJpbqZE
x5AFQk8Gp9Q/UqHK374euLhubesbLzBijD+nnaXXcra9xB4WQ1lZMrLEQe7u
7HjBz2qJn7OeTVHnWuzLi0pGr6NbXS+Xj24+DDamo9Ae38iEXarhcXdNTpyp
2evAPaUQz24wGm93amUIpriFutB0s1JL5EmuaItNt4X+JN49Lgd3y8TCF17q
MGLsZDTZ1h9iRG/MtKjTcSMj/Qg1MrloXlxe/XQtD+jxUoybuxVcxvUU8q+7
YIHsO5tO608G38socD1F6NiT6rpvImUoQ6O+/FFY0gAqDwUDABirEVTbU9zc
YPllPAgxujh2lGwxLzMAdxa1c6svdu8sQeqApGSzi4t/+FbZH5k57Uifjoaq
yqatzQDQzyv0gXcLETr5g687GjVj/5T9HTfwEms2OwT37Qbs2TL6GHz5+l0w
GiaLDNA3du9VN59Xd/aTX77pq2SHe9D9UHqP4x4R4PavU2PmJFcdKi0ssIIv
UmwEOooWQQv7O6BQrUFFq583jT78WpIkVr6gXnNOPh7J2ChspyrPVxtsA+Fa
47Ye14IIJBQzw8DKpGPz/jLXCNHMIaeiQ2Ci2OyZzWuK2/usmpWVM2GsaNnG
58GXCqaIxZFcD8SkSf5qeszXS5d+WiqBBjwdyd4DyfnKER77HqvkjDg164On
68kTH2h7Dwj9OBaZhnhV/XTlNI2aG5ykSjnZhCo0Vgs3ZayzeNGZdmqtGGV4
/VWvLRaLtPLfR7ZW4m4nL4z0nXWcvtTmQ5nF7i/sn+hFbdeizmG50vvMWUar
LFwKol6jg2pjDU5qLCFm4Pis6gTfkj+6W4kpQtWcGEBIviW//wYepKTPI0nR
TpuHm/RbzdlhcJ0ClE3xmVjNoXr9FcxrYJtTpd7+MQHyVftC5K1hjYiDzALR
jKgDfr4Rey2zefW6z8mx2SHgxXKORCkYj/pisX0S+nprd0WRYbGk7XRp20pH
30MIB7oNohLcHlDhZM8LvbP29dU23hdOP5CvsqsGdhxkR1D56Ib0BNvobhU3
Pvj/2wBzKs3m1eUd+YLwgkFb74swayqokKOUKP8nh7FBarykOriYveFrWlHA
PjH7Jt+UFjErKvb/54ajHAL/jEOzT+6o3GBRR+azbRlPCOPbwe4pESeRW7RB
P0eUVB9MSPET/dDC98RCda5LyATokDDvOjgsxXXKT3QC/NjcadANqTihIbTs
VUywr+XdvFbfFMsNLTSL/QuB5Yxh2Q4BmxkKS+Agyjv/QcYhzJzctGP6DX1h
sLPw8grmj/Ped6moZp2k0K3+T8eCU0KFOe/koW+wxvrE334Y3qwc2v2TUACQ
a/T9mOx5WJVZFNDsm3jU6NJzd4DJY4NHGQ6NKhbvDWeICKEtSya8w6lag+G5
HdALbPhq/NnLewoko7g28cLE/1pd8CFIDCFNSrUqgS0rn6FdYtJ3y1sshLpR
EV7S4SCB+5/8hHN62y2pj+Lwn86pwp8GJtCSbhxXwx7PaO1hdM5jSWGsPRXn
6D3CatPA4/zVEuX13PNdRZSxzxHYA8L8XmJ9XQlWVOIfVFoX/ZsbLaTSlGCE
dNRRvLJiQzjYygo99kHdHEEIc+a9Kb2P2jHOsM7YKMBM2pnklj7fuLoJjmk9
b0YkHInvNifYte2XEhjyOdtzpVaHJvCh9P88wq/yUfj2wT/X374GZ4VtlYYt
N3mKUUoVxTMvninfle0MPwVYry05EMBwW6T+6QLQ4/N9xrSMYWYZ7OHvus2h
pDoD2p2EtKE3Mp5Q2TA2Xmfgz1I7xLlvm+r2wz2fES9s9OaNV2DHBQCy83zv
B+vXvwLFoGcpbdf78uPc/B+nn5gnBC3+PvCT5cofpsi62pnDobKgsMxgzBQq
cLRMws7xlXcuMnjXvAd3yn60MwWVUrZaxTmtJ0JqCheAAJ2Bt5V3fNBCl4K9
bpM8JMIZ3nbr5YRIaXfp47XzSM4OfTEqTQCm+4TA97euIwi4fyjhkgLTOxs0
dixkRD8KMM3Juu3momfUEORLszZBzfIWuvHc8GzpYIREiCwDwtA0jqOhf2uA
ceSJcA0cCJApcUr8x8TqphUx54lFbq1W2AzLR87ml2cXf1CLF9cExtBiSYih
oRQGtKeMn6LtJN1zw4nmpHiQDInS6mjIqO5FrpVyP+2GMFGIvlgCnGs+IX6E
BHG2MTFNSG4xaAXE/4p6ZSlQiqHJy7ffA6njng6vcNnDbMyo7/WLO6GBzuHN
Kcv1pPkpSsW8X38E0vhYljWGfeJogqCo+S45b8BSCibXwWrme7ltiN9SQcx5
NvDKDDXwdiJa5dHRPzBaU1oXR29geiB+vc0ZJfqiab6GZHKlAlCKmO2cIHNZ
HJ3AbkjKwTnyrugU+l1Mf+MVxeJksRVAzRmyi/jXmkHL38pScgJYb/o61weM
4yxT6S+ie6JCY1JuCcWVzOfeveLaWhA8opnbiePlHdfPDmjGDAmlzHqt269O
2jz6LCiIaZ7aycmMTBcniVlSElBDQUHSRMYLJKd6w8ss9Onepy3VBx1lFAeP
GpEDCzhzBkX4qMNozRwIUJ6oMGcf3qm0CelmTBRRWgW3l4ipdSkhaw7LS1uF
YMvVVUyNXms0EQ44NrNfxTbGpCZCrwPLCHhMjS5IiEYEV3DZDDJ/7BkVRLoL
2Pp9yQsNbEc2kDmC5g4TFXrTqdUusjeUFT2+hn+OBq38ad4FvAiMU9cXRSrm
I6Cqd6EWSh1l+L1WfF2rriA0Xa6vU7WdD1Ztl28dI2c3xyMMG80oq2hZ3Ut6
6Y4EAI4YLbrhKB7hfciLG1KQYyUKD6f2+rYdIodAC3hSkRiLKKxdGQ4EYbUu
keejOsqypQtNgNT1dXUaoM6C5m0WK1jRZF41qhUP3hX8R+K1D3RN7DbUNQx3
dyXpZbzTdwy++b/46difa9QtBMHCjnSVPugjrzior5JFfZGXiuSb44Nm76lC
iRBj8m0HYIPYRiDGZWvdF/2lkEijIVFJs1ga77Zq9GHlAuCvtLfqc6HlRIft
Fh3jxvIabM+++xA7LJR47vZNcFPb2H9cXbK3S5u8gRQP6MTL+xh+Ui2qHA//
Jqk50g/707YS7KiRBSmsB/Robfyjx+OF1NCddzNjtFOCw6DpXTB1h+8R5FVW
8x3N1no81rpczjE4IKMkzZAElIvhDh9zYY9jEHLq8mixyrzj66vpf1k5Bz5O
2a5HwW6+xKWH9p2qhWBFoLBi7pntvyFZg1JBqosdtfu/tJmCQ7akKy+Iqhkz
JhpWaSsAF6KJIPcOpbWwzAUnwrJQAFaOrs8KJ+52yNdJBwCbhowcFbMemXm2
kzkoBvWpjlP+RFL3fSgoZ0SeebN/1ckf968QL/z2OFOHtDGHwjplSqBvtQve
INYpuAOE2leT45de8jFE255q3u4ivB5RzZEZc7X+vr+j75DUM80td/2TRga0
CF+CKlRCCOgjRokoYiTdXep2I0ouEy5TYNwg5dNXMb1MNPklqGofKXO9jhRi
r7HbFeSYGjKVprLZ9bd+yY9jPBzxN0rpJVCYIe1NacR6b2dYMukg+Ixyd4Fr
MiSmJg5PuI8M+/RI23HtNo0zn/O2DTQAUfRaGAHXTogzlyoX+1Z2/mVbKtDD
9TAFgEj6uhdyui/U/5W38kGNEPh34YtCvERN2IAAoN66y4oCFIMjd1mmskEz
G9Qbry9K0JtNux2elVBs6YbMcp5jPeIj/gnv4ANdOIsNpZRzUgsm2O3eOW5y
5E3oFSnJrr4zhsBBodhe7Pt8fpqquW7TXtOkYh6b5WEiTjvSTKbAaE/OwvwO
Qhzt4ELrGVteRCRtlCur/TqgzeNQwCwzKbH5x+rgm47SqPnMW2eOUt81Y6Ll
d+uSMUgZrWWgGwqIA+9S340bj6oti6rmiY8Pylv8L1Vj8QHZyM3r6S9EYheF
Aju1TXOGHJI3V9uS4QfRAAakjSRsGFNZY8586iHk7XD3LVksaOraor8v0q5B
pQvZnF36hxGS/Ii/cWxm+d97Yt+Ckq/7fQv5hrN6JM4uKeLA+SDSKpYQMD1r
UtgDupwJ+IvFlwAMlA0jaMVep+4XXd1CKZ8qY8DSmqSLXXokU64oAf9Sqf+2
mi/1uWjyH3ZJFiZpQFYK7mM/tM58sB9vycey7GCVOY42VhCSQVnARVDy7foy
CwdowxeSKBclgt4/StYa8TReS1U4IuegyOUmjO4F7o6vWDGyL2AQeVq+hAEN
ZJpW0sO0t8/JdREAz/hNvHXtQ+CwG4mQIGiJ8MvT5QqqrztOhp2inF2tk+w9
/j533yQ/gG0NHp9ji6dzS93b08uMVNqQthIjn4EFW1GmZJ0Uw28DRLnRRprW
LLb3mzSP23UpVuZ6uuTUjb1vTVSNjW48fTL68tBMwIE8pEsmSwDQwOz0kAb4
iUN/T5gNox5GCnIg4dlucno6kcXmWwNyDQitLqvv+Q5LnZfekmUoB+GeJC2H
rttssKn25VTdBny9Vv5iGeTvabcG0rMPrUHfLInfCMEaZ5o6LbYk3ovUiYBd
R0GnpCBtCejc5i7IbE2Ne9T9+P5a2lsMhuKMQ4XbL3QP6QP0DckD0ptHtl7j
2G2FiVQPeVM+Wu3NKd7oDl7aSb1HwwICEy9L0BYXp2kLOBRmWtj9LQJQMWuR
DBJu8Nol00Br1qwaqqXyqfLs2nPJjA3tfvqMXoXFx6zaXGmTAKh5GlMJzIAq
dOFnNzNsj5sUzr/Bvmse0DOVZU9UmxWeK0km8u6GrICTY8r1uN1O4Ez2SPED
k/io4nj20475MxYjf+Cg1mMVksUihDJv+pdRS4LCgSjw2g32QQeKcRP5HsDT
Jg7wm2kHgHxafxt6T50wko/mBS7lZCaohU7T/Z9OgbC5AsCTWB8EsLdETgVG
yk8e7x/ZymQ76acue9hhExeJGVDShAX2IK1wB+VRiODfgGmDHL9U3JlPIajc
hwaKrIV0Eke0Pca7ieEP8Z9Kdxd0O3zU+tzJ+ELzrxz0zg56x1V/QaqJTsZA
c4zk9GxCEPdvwCvjlXLFUCQLaCtfu2uM9a3q41V1Abytr5epkOUqZ3mPggQq
7xickNOKnnxWpnZNDFGsXl0aGJu6nqPAzh7X3qc3UqXBikWUTmaNPXOs004G
8Xydiha719ZhkijvD5HkERO4GQXYZK5S+ju5X2KWpTvXFbRuQhr4VSlcN6VX
/Kg+/VLF1h/Xucf2nl78GDQh98C7N1UEAoUYbrQWkr7cVdEHzXk0nbkWJP/h
LBRRMz8mjjGw3g8Dl13nfpIsOGivMfANuAw6m/ycrtMZrBCmqpi3PYZuvlHA
15hPu+K2/HBPWz5jwijwumRRRUhJPK67ILw9z5yR80f5wi0PxNbX2D1cPg5s
5KQ5zhfZgKu1A/vQ5i+VjKJKAsyF2hTMIcbUJ7Ws97UkXYcihJKMBoBNmJFW
1yaHBJmqBAUCCMxFg5XmtWIL2OJK4+bvUGa4s0Jm+XowzeZ5IzR4HBxd3Kxj
bpll9aLReR1VdQ5h/upFFSKIvKfcUkJP13pQ0VNHPY/dt8kI+0uyoBKzhkvs
3Fqp9OLb8rXQPDGAn2/3g6L7fOQETC6xw2yYKZawG30BQpFgQq4IQUx7BybE
7va83xKfEVKK0qlCf+z0WlVM0B0TMmcph033XZkCS6f0mLB120ZnJ40bVPAZ
5neVq4K/38FXWqiezSMa8Zp619ZxZCfmzrS71DojNme5Jy55XyIwYXslbsdT
MTL6YjIP5s3CTrxCmb0jML/hhbLQ1/yLcbwWvQxBfqYJuuUTnIeI8OOwN6Pr
OWxqAi4yypxgEbusQgSoWAVAMLjlE5rZtlofX21pgWQCZ37OMgExu5a/QCLu
gpOjx+fpwuV8LmS6Y1Og7eK0ZuMmhsv28wtI0MAD1urq/1lSuYcXeXTinZC9
Leu+rsbSpJT9p8QgEkmRRDZUgxJ1QfM0uHvTQ+600vDMgHBX39jkBoMBXca3
TVKlI7UgC8cG/977AaDzobRFPRJKoOFQXkeaHM9UROIz9es7C+kyXb3vOhUy
X/RsAxBhJgQHGJzwlrGW4tu9Unnv0cmc+cA7tNYotcb5IkrVrzCeY8t0q0qV
UIrjD3nyYz4l32LKsHsQr9bRtqXbn2XVPYZ+WHazgsYVBF/k67aIMdxlUS/H
mbpPKzuMZxRHk8pL/5m3X7SNzAn4ql38njPZmjQLpiGqiQC2q4Ch6c0btjig
1wUeDpcL0fdQdy6M2V32R5LdjSeUMtvaUp/mKkn/LW9U6xtTGnQyaeEFvbkt
Amvm35Mx+Qz1/n1fK5vRIux+NoSBCriyRkfl4yyPJtuIouMT101dim0SblUh
oEJ2LcX4wz/MQw7G86Zs7APC9z5Z+AW0gWXcQr5qy5i+2c5hagmZvcMEtGpB
9Md5jaxgEs9qY5h0YN6eH7rGNJ8fs3omTpg+ECKSO437t6NS7i9W+7b0H0No
NelPyM3HBZKSzVJg1Ff2pXAwZpEUedRZzPeHhwey96nxXS7zlMK/WtVnNxJF
OVfenTQ0LGRiFE2T7HxN+BQIgFwatR1myDVBBfLuuvCWwNUi2Z81OM2dbabe
wYLcsqPrRujSbeCzYe+KwLiJWF3CFBLevmLwhxRFx0LRCVsppYwxQe0gOmqc
6bvp8qAF8G3SptQP/04a1oNev0DamNF6QTAKq1ZCksHg3wpnanIgSmhYRRJX
MvSLCOdoEVq2Qj86iKZhrOqZd3iognv7dFo0Exmh1KxzBIn1yKeA25fSYl4v
GNK0whPVHTUnpthfzLPp4fM/tgx66AQ+Jv8gXUveWEKrNnVbuZeAK1oKHnpi
NV0Z9awvXg50qoU0s/b+vnmL8d2eqnKIG7m6fA0SNyp87PdfDWt//gRvesXQ
SXn3Y4iDebKnE4P1HE6ghYdYghbBCF01D+BFJIZ+EHSBrrCtaE4oCdOa66N8
BLbQaVA4yHoy4cSo2QtkL4xNqfcONxpepdAjBbanJZQbdJCEylFrOCTckIww
sKf9RYlEIGs/vimH5FASLdvfwsPykW6h0h/vbzDLhE/4nswT9qeAtj+IL/TH
9jlNRzLY9PzLnKLwPfpqKqw0F2XHvsUIzJPP/Z7X6djCwcUxtSGiz6piA3Bf
HMveCoqv0WThMtp0DZwLYX3YQdBXS+FGPRQXls+RcglFaIqk4z61K8998n4f
MiJiJx7xBMw6QvxzwG3iDuQK3gnhLwv+LqRyZpw0HgtBQo5NZQ6/TC1fjYO0
AflWE9iMwrepaB8I/VD4UHYPHiPvF6buofCjmLSK/rFlMni63N1lWc9W6dIv
QqCKUp19cdnK5wgvVpph7jHECHOYLZz3B9zkEQbmsQWltNHf1TP+J4Jzrklr
J9ZsNCPPlfYoCONw7lCiHH/TDvN9nizC47B6/W5hv5k3P0Bu8w36ghWl1qFC
kVmU5Xs+xy03zDPt/za10q6lUFGAdR9M/D399klbYQTcYX9HqDqzRa6HgjFF
P1im2mYvJvlSErA7vOQQq4ex73H++yxR6/JGh7fE0Q9pqA+WsA81ilLoA1Xh
jNz1nvKG6Y2pPAKjBTqgNulG8g4U4B0t8PWjgGqK9+ZRsStlBj9hcEZZ7C8T
y5Jp4dW9CK/uz/LIjwiEfn7/zikUH9Yny51ku09YaHlEQAZQhJ9X+cKKzLJu
Ytlh959OEWS+nMpJdXfIHxFUVbCyatDorsZ/lEG/euBkXDDS84MEheq4K5MJ
GPALyRScE/+/SaYSZpeCDyuVKq2pLtjCKhNpgj2AMxvuEV6OOLIzDvY8NQxb
qQU/HmXKh3lV1AtE1XYxMwK+T0xmD9c2VXgwcypHdftXnSt8FTx+k3UP6yEF
Kc4g8jnYi9KxgS+q8hXlQs6Kvp1o7ATMNopTqPj+KU6Wh1h75Jg+ARRthtbe
qRzGWSJ8iaLhsV8LP4e5MAQ/7loW0KnlChNeETd6JMoWWd7BD/OlFJnDlPD8
pSSTOtzYjJi+qhD/RJA5YA9WS8hLdoQgTkyxgm7pqUAUEDjmopgKqFrEfbMo
n06gRnvoBU/tk50++35NU/Q0p8kyhhlK9IABDeHjO5TfDDRpjwaG+2HBxMhb
XoLFySaA296JpCIKTWO1l0VJFnPOp5qP8Rz3P3P4j3k8wi/UQsUov3kNFSbs
ymiaMPjuvxjqQkk+DwWxcGvUqctJaH/BZYxGtbTJ5sOqow17gzgwnSyDriTv
gPQij7DUMsxyNwiQoK3dAsjFwHqWMecbneMN9jicwgy4EF4B/vZ21Y48sw7J
vfQgI7gxdzdTlHKOShDXplL1Fcc9+tylqz03pXXVI5zmmX1+PVukx+nv16i0
Uk/XQANUlAnyrGMfAK4HkoI0ZxNR9c/J3NiNoMvz+tRIvxw1iR+dVe6MijGS
HSBDHSvXan8HgYC9dxkP50UUihZiEi4w8N0PV9jrJTlNaz4hOhUOR+lbJTM/
u26zaP8yOG3WA/OjoeaSd64pBHixG+Ut0vwrn81ZSieuz2juT2eGsLQBddZO
/P29qkadFeYdMqXqIITHhNNU6EMfpBjVMQtR4WQBdfenxRrXYbIfA55YIvMY
vxw5wINeMXb+0XTg4pxM0PnKS5Q6B3iKwLJ+vXLqr/vmVN3KazSyKzgRu83W
mI8GWwDe3wkU1unJZ1nJEVeIkpwCOvXbAi+S4YFtkyY+or8ZfxdEcl5LW20f
EKHJuNamEoB70CPC7t3bfyINxFSCOEXpPP/f3ae223tA1gJBdhT/0aPcdrFQ
lKh4A+gZiHbsDQ3cD3UO2ZDw7vpJPysuvLCa1wPtdfA0PUnCUe71ucoTibiv
0IyPoCz07mcNdObSFz8MbFB4EHwPBWJu98x9mjVQaRgocrH3z9ldj4+7VDbK
tKVkug/kY7EqBKkVk+WjOos756Dgzl6pXqr2TjcHDSC8nC/dH+aV6bkfOUne
37uf2AnD5SFTkYIYiccbvNmz1+3Du1HxelQUBDhiL6ksnPZcijtzMiX8IqE9
WS8/SpGo2m0koXx0+UdBKVYqbJsIZAOnfOML40JvNyO2WkzTHtPqVjbS3osH
FPAJjXqB0u1bUihgLVD2b6fqDrX2iceXWvP8HAtQvBlP9fD8tG+yuLWRpxoj
QImXmpSTIIQCRNJ38vJwM75FeG45r9CwuYgEves5V9XQK3dQIyg3GdSYRftB
Qk9nTEwDThXixFHr7ILfRFrNy+88lA1K/Dh92AlfZtb4wTsN4kBQraQlkECz
t1lJTzP4MWmoHIzLxClXLwQbC0a/cZa4kQg35+d0qxUjvtTTYM+OweHudVxV
6E6dRKzOmVOzHn00yVKzoVqRJT9ckLJa/OEYmAbkgdAckcWrYH2NL4AsvWfC
Snq5D6gDETa5IHBeK98vwRRlMg/FqyI5pkjKhAHonvXEmEcwHDxjjio2peXv
F8KFgsZqspoDrF4qKECHCQ4A5egMqcFbH9nbC9iI6nWH9obDAdqX8HTXuNjc
NyIfQWiXRyP/h1o9PSbkeeurkxa28Seg3DI5n549ldgW2sUfuNyCINJl6LQs
qtWzhw2iEXK+puVoyZROwj/FddEjH3lujBkz0tZkX6laQmSugFj0lGOb9IDq
f4llOuorcaNO1hFBQO2CJfd6Csq62D5qpCMAobH9qJ8BvMyneLclWeLqDTyP
Z9+rOljPTYhFjTaYnGgxVt6yN/USYpy6vkoaseCPrKSype+4EHmQmrGuOUqW
NVInX5MAeGLLtuhE8wJnJ85oFp7LyvALDLcUiy7ND6nxpitlvfezePkSjaSa
ze8ocqEyz1PjJaYEPuq39K8qBgDBtEISsxh1sATGhjTLZZY/xxYU6f2eNG6A
rctwK1Wo8Kk4VktTQTsMjyP5kuwc+SnlIO7+juBDfp0ITEh5YfuQkuf3pgU0
ynZXbnqWe4ya/nPG52Ze1isCxLJM8RKIOGjM+678oC9HjQBoEd53MpquMX1x
QtnL51XNYhLy1U4MouVmHxx/ndcdB5k3gcxIlmQLOEGJ3VlszcNxU1hewWdt
lxUXTypTqycdA0+RzAzZbDgqR8bzUGIpokrmBGTh9WSDIdt6OL+bvvBmFkrG
GymkeTEAVM+zUkhh+zhvHTDhAjXz1AZid2OKd5kLQr32wm/V8savA/2af4nD
shjK7OcY1x7Eq/QtUmJHRZ8R9rpHS5COF3eim3ha5k+dlGyiQz2luEdgMQll
6S0PNA7fEgamImAHA+2uC0SKUrbEj8SAx02MtXYIToRkHu0P6xzfE1RL83P+
WHtDPgjMLB8kQoE5gIC7G3IiKr8fhE6vhZCf9E7v8jhkAGIxTAm9+ECoyRGz
2YOlXbzNUIxyLCwSdnL+7pQFtshSs5QaAU5Y/sK/c0ryPCE5+rmsnMIkhN5L
ifXdn+y23bMOE9K4YmGkhUhYOwlteYZvXCkCVjC9AV7gdnjTXaIzHAt+RCrG
zEtLU9jRsKowPIeTitP9XqLmPhz3A0O3IPjZ/ppV89x3PmgOjnwdx/7GI5oS
0K+EKAP0LWkrAvj2ctdd3bkev4oOhcxpoWKlyivz1rTVHA1Y/Tbf/qBysMdU
V4Oa7IdFnjjxaeGGNHFqRtez+6kIO7Yyme3FaEN9ii/1Q/ec7O5H6g2uvztG
N5mlGkenOPMhaQr317ONgYiD+7yOwGs3hs2bZOKC0iZS6vA84MM9lx9i1+xN
yGZWzIFAEiZrBz+chpypLFfOgqbqZ3nU7YHclWszrJc6bZLIm/ncPav0SvUx
gyJoK0bbObtkAQ2rvEobQRX2m2slR+6+sHTSffk3mza/R873Wx6sfz8mFVf7
Seme4j/rtXBsBBV/0n/kv9Rdf4CiVYM4OpMGu+8FTh3sGCV0vM5CuXCBKcrm
4QbSIaAqb1exNbXHRoSix8qFpMd0j4J0uWbtLmHkPq33DqUiDzzXWFHBOrfA
Mun76Mne8cv3fUShgXbPD147fCcEb17p5/pebKpAhtZ3aBGUZn3nhx12n1Nj
rjLMlcshD7zzFPKquc3N7h7N5FcEA+iyWaQ1ajGZHmg7hyF2bwNdmvlXugcw
BTy8sxswhMZFpyq2ZHEEe8La45Q9lq7OYMFNCbH5pJ2brFShIMeo4zOQeKpD
PUtP7LAo/DZsiJlc5kxjIMHRtJ8DEa+H/VDYa3gABpJqWsoPYfIf+wvqkhhl
0iOhp2W61GRsCH4uV+KJN07375DaBA6K6dAdVSZWrVY7bazB9uFnmkSmuftu
EWWosgQREvVzysfQAoV/uW2Urn+C1CpWPRaSGTBFZ+/5S825q0GBQx93zmWJ
Ee8RR+olH+TTvaWRyWzle3H/zTX4p5B3mxwglMnYok6qU9QbUckCjcuU/Zgj
uq4jD5BzFvKV4uI5fAfJY04z/Bg7QoCSqsVS/SKep+/NaiN+0buzeySZf+hv
MvxruyzEqpiS3Z4n1NfSeskU/vT0FcEhPJknTrHtI3vgCl31KxRElDGHGTOy
Yu+lL9N9cijpht9Rk7THwzGsQWvAiF9ADUi8HBNs1pJ3fU/4peeZ80krxc12
DMVWDChR6ipctiVHwV8YCssNnWazEJLq2IdERATugz3hD39DMrNqa1G8TJYv
NN90gzzt4XBT5TdhzPwiwkO1oDepP8xR/b3FzWjxQ+/Oo9yMc8E9CDoXf6Bp
pdgfJtdela/KVnon52vm8myM3c+luQr7SQNlycGSIYmgV+9BngA7+uij1C2d
vYnn7hoR6WrfwZe117Fl8GVarbcphuZu8NLAIvqRcUU11IGMmsYD9+PabjSL
0Xvzhu4C/ZH/yPdoemnNet8y7oip1gC86cx12MsNrDYmQXa87mragpb/gcvu
gyneWW78NdAW6tMVVmOtkkHXLB0fu/P39Juxh7fDXBt5tuSIikZ3+SRIo6YD
7O11RyHn/wALi6t3yPajvVwiITn4czbQO5mvCX/ly5FB1pq3TKDbdqiibQy4
r9US6Zsq+frCjmVnski4gtSFJhZke6P4Vb63aoDABPfhjFAwQtHcY/ZGrxdk
U0mZvkYmpZbfqhWQmXDd5c2Ww6Vh/o6cyH7WQw1YU7XaRiLMEFzP5QUTSomT
sm1j5jB7ifald18f1kmHAP8KY9ExtsoOgEnvmLVM++M/PKfkhz2aA9oZp9a0
5HuPWfT1GkvoxWX+gdBQjpye+mU+dTFEgxOdLV34ydi5XQzrd0LIUtYCWtQx
juf5Wd5hZaoFDV2M+1T7bnosniJAWVZwJ5fmZitHEsst9kqMD+jQFnM26R6G
oxFOTdtOk4DFXwCkXcmvgPppOT1G7Onrq5cv37YvqrZcFJEktggBYXDQf6Wp
N5y7w0biL7eeOYexqipD9HkVPGgNzTbjuoFjFTb/T0xavpMd8AQaHVXD0Y0s
WcIeCrmvOwHiiejpEOkidK58yZ2g7caxpPD7GPZ8p0Sbw6CyQWkDG/UHiTdu
0YPJUmtkN67kWJPFbMB7YwFOY+jXj00RDzllNCe4luiigAtRqJMMd94oYL+z
BQCvuNqZsiFISvJXU6/Ua/HvTRgKBVFgHPDwfKZuockdlsqwdXxTeollfWWQ
y9ojOUeUsMau5hrDAJNfXhmxCT8zBsoGYI0DxOzXKynZWqWQBUfkUYEcXJ9f
YXKBaHDJX7kIfqboj4mXO5oNCSZXOij3ZYbf3BXAdEqnUqkOv0wubyZKM7Yc
FkZ9Zx0K0wfwrhb9moyWjZeU9JlDV8+5aYRX3t+j+dgcnFF2rCdxP4cBFbsd
WIJs1ZbcHmP60Zt7dZS10d7nrtg28A9iBrRzj9OUL4x7YvgHU8gsbxwwg01J
jCLBncsngqHOmRSD6W5zWgonGC7KpO3qvP1UYL8QB9g0YbZqS8VI5+EBYCO0
s6JWZJK4f1xlU4rdTns/yHed6y1a+vF/WE4y1tfuobC58CUINYFoz/VAoB/E
EHTjD6Uj6bCW9eSajQp6RJM2hFSw5yP3kb6EsaGeNRON/heStEtW7AfvyN0N
zkz/dEUnnIM8DqSDvqH8icKp3bDbCZu4uKDdxUIA9+WF/Lk9bqQu6wJKZrDn
hzoyPzuYutAMrdBk49VWI5Kg53pCYOC66XoGjtHu435R9uBWM2DJHO+edn1M
mvG5/9gFVKwk7sHwN/SKD+wvtcwerPYzdruI+P8rl2jWJarEz3JuI9wd3iDY
P3ZukiLKolGHOzkyPQDwQJm2cPl/M+/Xgihe5916Tf9rk9ziQ2yHsdZPjNjt
Uw4/d1qihspH62zyvZJRhXXhSmvbPIaSHv+dy+6rPq2mFOCSV8wgWw+qHItn
7EJTZ6Y7v7NEaaQl/JvnpJXQJX6HIp47TVhT2JNUzNVxNqIIIrUGRD9/kiNA
f5dFyZ59fugOGb7cBp6Lt2WMbqya1GqT4uq5l0yzlwIpLF9CTP6zKFQYPUw6
OUC7Apu34/31OlreqXu4esbNyYyxaHzC1sXAQI7JRPmZ2zVouf/o0SMW8dRy
gjUFxvM2zGZwqe4gi6Wb2WFi6VQrIZWhtb8dvPRDSEUyEVQgwvGF66rI48Il
XegX0khLFsjmuIKqG760f4oCVtnxjujzBtQLrcLdzVqV4GJHcXexM6fUeYHg
J2mSgdf0REjbvs75TX73/8P9kv4dmC07CgqyswNUPiGFMVAKiL42xVvQJ5Rs
5GILPgWiHN9CCxHCCtlKSCZgWVlpzWA7EBByv2oUtlgreSAzLVdg1hXPfL+t
MrPqmfijbWo1RFeXPgnuyUWtIAnEh8pBpF6mOFe4MtLaGZj93DrY28Ysv0Ly
FTSECG9wIYxjHoeKCDmkSlX2VqIn351TQJhv5JB9IjmxFE77rGGnOynV5kA9
Aw4CEYzU00meag9m5SN1CFIreSPVRamkAFTDqXLckS9V5PS1aHjc91vGfp3x
Dwhexu2y+lZkVFEuhkhN67BtBqpaUsXzleX5Fcstte0A4jOxJCOdxlF68gjq
E+a77vG4tc+t429kvqhQedRguqZk9spHJh5DOgoY6/9kOzmL/V5JqT7CclSz
FQXhcsleS7MyzkHT+TprhyhJTRCX4BW/SHfuTGs1e2z56MfGr+Y/awNLKwC8
pTmgbARakfLCJqWYc1YJazyQXw0AV39vATYRBtZQ/0JfHAEnn6hgyuQYeYBa
m4nUvrhLwMN7Qh5nwtj+5L0GeQ3H3Et39Fghxj/Fw/HWEAYrQazb70SiTKFz
9SbsPtx+P8BmBqNL2fhXVPcKbdiMplIcBtq2P4fwsPyvZXlnLGPkqFL7oY81
fpFD6IdYo3hhEtILqymK3PLHVW+iU93Yf5EcCWD/2L3eYyirkhfrBRTnptp0
em1/4rDmTVqKPr50EANLBLRoAmjZoVH3dzlPRZlDXuw6hmvh0dqscjiycJoq
bxXiWDjwPebHOtFGR+mXjlkvKGDa81WGcy122+fTW1lTErMCm/ENYYlLrTAe
3AOcoBlS06DeDDOT8lJiou+cSd3ylgTlYLSYXoMxvPHrweJi1aW55aAGymis
AehpjJr2dcKnGaNxnXei1l/j3lpp+gHg5lDlsqjbxTZVz9lW15CQFzO5NiFh
R3rxQacgJrTWPE+UdrNCdiUgXuE6CLsOH9k0QHoT+cJa5W1jNa+jrPlmVsGN
UnZaoiHEYhnvwFm0rjVFbvgW6bSKXA1g9XyqGQ93ENSEqjBOYtP/RUcXtfDi
HOlmiTTfzL6cWKxr9is0+keLa/MJMaL5dODt+D2MXZ2dOgyLt5ZjXiBDUerw
dEG4WbI8kIA5tZzCq5zMifZ/VFr9mDi/ESkavUGXJud0M3qUHvrCXGoPhv3Q
RGwnOJj/epQ8YF/MXq/z1UQOvRbFBnyfabOqBkM/pJLlTYvMQ5D34iGbh+PL
yTfS4LmphJQFkYxjWm521Xud61Ra7JwO3f362Vfz5afFB0gOwo/OJGb2V0d6
IqCmPIE8g9SMr1icw3XxOSDsO2TK4LBgytuS2amOO8sfc2vgSUFQQtFEzcRb
kCCI6bGRo9XM7iR5D8eWBQJPiMp9h3ghwaJMuenbSR4pkFcl8fJQ1CjnyjVQ
pGo1YbxjYDfenJ8zLTeDD0LGeUfdeDBvhVCLX3SV78VO7V0sW4ZsFgo4qnXz
K1g5dh8AM+ZouVPml3u2ym5O8rFHxTt4nYDPpZ8Y3RGHN7UXl9yP6pEOxyne
6ktAgNpsxQzdypCeP0akqAN8Pyz2fZ/UjWuq+ENA0sYxZHnmlshPiexGA1cd
j+fisGb66BA2wZcqQTnjwM38fnBM0Yzd7VE/3WzLT2P3usVViD1OiZOmxfkB
Uyi3z4RwsfZkkYowmLMc0WosxM1+E8izJ+DjbCUeoZj5fmW6OZq4D6IXpz/G
Z7WVkZYwn2OxP/abTzXrNisSaV1M5ufQnRQKr61QqEL3ObzwlfwqAg8Xj33k
UaExZvd2kmuAT6GAY5Xou8iRMu9bzodQr55ntura0v6riwy7EwQsKtf7rjQ6
rxBo7iNuWqUJpdb/Te/DR2YYyU2ZGzlyzcdPWXNH1w8CCxa40Bl0t9F5yvwe
9u0OB3mh/egHQ/1Ve0//EzG2IOsC+RtUCRS2j6PQcXovp0tj4BilfNRriGS2
KDefMa133GzJo1uJVWodB2pm3dySK2T6SGOva1AEPXESV5nAx7n2qOoJ/cAm
dT2GcPNNbqnwJP1TEwVtS9993QNkEY6yMNcJXQqwzj/rdS+6/QXvy3mgYysd
uXxN0eiO/Pcs5C3AYIG6AN0c1bY5dH9Wo3h9d9eHwD9gOtrDxfH9e8hD0bQn
86a50tNAe1c0gfKgdceyVFze8NvvWryj1tVtuq/7GAD0PpF9uXHj6Ph+EEep
RK5EghQlGcrPrhI+U1tNwtWrpSu5yc1lquDtd1mA0uo6ZZcnJBsjSn+DlHWE
fHQw+XN1e0ZmkpyK2lE1OpGvgfvwoEVucJdFcD/nukWurM0eYc5dbAU1ibt+
gMMDLbm6xHDfk1mWyX/49kHSenJRudsImGjKUuPvPJJTeosbSaWGJ9LquIhy
1Ua31fnsZsJaT5ztyJiC97EVLvdjdoDP+vJYWAH/mZmWyD2z+0LY1lD+Le9o
vm+kZ4NbYivgjNxrg+F0vfEcLQ3qI9Jmq8EA/btBJ845Ctna/JrBEBFyoVis
6U6yV54/3JRDe/RmxfuUbkFct4v+dT3ibEpsdhDHcMBAWq2NFu9y8E2MyyXr
vh+mr6NsM8ntCPflz/XHzC5/m7Vhvj97a8RiszB3ro71vpLTa3Y4deyB3EI7
U5+xi2Y5lZW3eZ7GjQLmWZ8SjU0NEx86cgk3ll1FqGiLGHEwBZ6hktcN/Shx
e5IsYhKGKGwxuX9h/MUV/RNMnB724LhtAztbtiGDL2TZTG6Un/hjckhPA59h
gEl5Z7I2EsOSR8tl6DOPG52RFnxJ9wDBsQa9f4KKkU8kgvl2oUUSR8gewLSz
h6QHM5yTYuS3EKVOgKLIDuFLPjVk1os1hsf31FtRuHTBRIxCNRjXB8GgI2F+
E8/2wMhkPrRmwyoveXzSJdg+K3Sa/4T5flGLzwePXE6VKIzAW/PQKLqoVZNL
/pHVkeD8OfZdqIkMEWh/MX+uuskt/8oA/Sg6quk6cEShPWgDNVev8PrkdOx8
KhExGD3+A5C6grZlWa58e6A5jUobJcYTjadRJaqncmKnNgGBjIm0a817FOao
kz/ZGbx6UDE6+GGahJ4SPJieZMA9irSS1YPK0af7b5skDWMMgdN0+vI5jRws
ALslMtuBI66TACsPCVvniKeL4pCof3xShJem9arm6iZV+jBMnafTJsNIVpNu
amHFYM4lVFB+JvyX5wwBzLa9NnZE7R7BKKhq2VHfb5m/8/fE+ir7mHFEKI/c
HgXo5JYAzvskqeLMbaBqj0ZNQm54Rx+/6GFZJxAwy5ObVzKs+MP9V544fbko
wX3e6rCrhdkHna7syingrsH+x/C/d1ovCkIdFfJv035I7aoP0WrG7XhYGn3w
K4WRghnsuNYwiKw9jHaJmCM1cCub3FeedLTuWXHmGCfE/ZCOOo2MbFo78lNd
2NbCTMxYQqqFkyp3U+aEiFnRRE9evsObwaYabvMPXVLW6OO2ubn2Ln4am1GV
jDHl5pXCpRCa+xhqppv5sPwtb4VUTYPYHX679IQCRN+6fn/agz+qjPt67k7i
6wP6DIQ8bEzA6j5RuipxhJj1EFepniKF3B7W3tpidfIpDDso6HwZuQ+lbZn7
kz3gnXk3h7AyMVlG9O6W238sWkEeFy34Bamm1uc7Rzq1lLrRT6riby7+AoNu
MuHn2CDUiGKcHLrJqYCatuwgt4XWpZN+941Q3WDkSL2zpFtLbOZ31gNEjai0
/pyNWwv1L4cJcitXk0XSYEvWom96FBERa/E0vVBUXIG4XOSAQE95z6MgGISu
ahNEg8VvRVRtm9d/6yxStzobwpmmaqHRQ6g2kXkKiSnpDh92Hvg6x4ve2yNu
IzGad0+N8h1QBejLumHl5TopKgEcZerdeVxzmeadgKOlNfwVIgbmzLMc+Cqe
1v6DUcbg8qQKlvrx7gC9SCw4Zpvl2O/YFvgo7fxNI2foltc4gy37udIBa8XG
66WAn/1yragvgJqw0jN+aRlF/3wi4MSpTpcCQygpSne0ZhENXVlpWHLj8k3m
RKO278SVRnlnRjt0WL2eNXZI0LSRDeKrcod9qoWcHWO8if+/iVHdyXnQ8C7G
OARlxRjC3Sw4l1OT6kkKq8LaNMHJZBDcxEFDNaupQXTKBdbwUbJiZEF39JIS
SRtiCaN65w/GRNWKrP5hhqALNnPF+OT+IASUo/dCfeBGbEVzQtEfX7lP8DYo
caD73IOCsUBXLk+hAhEcSBpFQEhgHf/X30zu8xJfMCfDssX3KRAnKSbrQEv0
ZysOKLYxv9aFCFVyyuuSqapfzt5HdiDugx9fXrtWW3HWrbCGpGY8TypnphGu
YihOOSUhnyG8fo+3BtbYGxGs2/1uddWTroiDhRGsc9qBLh7PoL7en0S7Pd2/
+pg3LTMklda9EqWIo2joCGbV7QtP3CjKsgbY8lzOeZaW+CVTp7/pw3RqeM7k
KexKrJH4lfrK+V2QkO0q3p/H34XHNWT+h3iZasgZaZEyiCy9WWd6RHUqYn5k
Ls24N4PrFfntDjd9a27NzMkziVk0CfUqwNkLBGX+FDMkvG/caZXO/JK+nv9O
1fpEqsJpgWhRn4/Jx7xd62GKWGEA8tLMJxKQar7Tpe1zWMydiaVzDVYn/O/U
taxVJlim+74mL1Vr3WXFE9m0ppp0FuKeH98ZkFzKVE7OsfKsJwX8ykklODBq
ZShXNjuB72jctLosfLLZ8+KZC55xlh2vD6oUq4dWcK+ZGKcWk0y4Kdh1Pald
4/GN9HsAczx86T53gZojHmOKhPawVUW84/wIgbDLE8RoGuc64KJPOHysDSWw
Fy1bfiPuh+TNyl7j8dXjNYri0voz4vXXxpYCYIQyPXrwRnCJyrxCy9ywcSpk
Tzx5bl68oS2SyDD1pdhVGoIaRQWRiPhFKIDh41ogLFT7p2PWjrYB/gA1iU9x
tDWbQ451pWqlhrVAhUv0rH2lkcCki94AO7p6hK+L2Xgzt0bmV0fH2tW6Srzx
HAtk1Le7H71t9h4APqVCsWMsAo+p4F5ct5q0wJ1sPxzyzD8Maz/3E2NmEqlD
tYYhJ2JP1cMY7CgjHnagM3gZcSdq3sTCirhSK/4Iv0KNWEfI8UpRtyNPXtfb
l1hBPoUw7+TPsFg1pyAjV8sOf0rOcj0MnOyUP3q8vhbAhYZwGaj9TLEHqVJA
ENxUMe/woijFN0QIPnp7zkpzt35P6+RlN2m0ieqszfAqL8sILevUM9W+pENe
TZdwhXuL7CImNf9J+he1EQnWj+tIZ4yFf5MQKv7kA9YDhiB8hWYwx4amapEN
7G6pE8QrAzi4otL5J6qe+4vDpM4bKESog1zQO7PCukpGxMV2O7IwXszFanxE
39Ez9FBGeg7YCtWmGvOGSsXsTbKapgSGHcKlJ/1dxSb/o5R70uF5qRcgWAUp
/aMQs3p84WEgdMVeDbPfF39+zl7MUJEusZ3AcYTueQQO+1lD9p+zpna/8I9o
P5DDO47Az6C8h+N3xTY7I/qXo4iGlMwdrt18XZNX+S03LvrZFjzQUVnP8BK+
z3bh+G9R4LCuZa15X1cM/8KFH/z7ewjyBaznuGMz02Uu+Kl3uVCtc1m+V9p3
ZaEK1jXu/MbEJzEykp7uNGY5rXAoaC2yS20UnMMkQhhbVXfgLYdGoFd9/R71
YCsRZsR9w/bJOPy8nnspUTMYGwCa2UW4yQirWlhfSaVdtG1n2Muh7J7GMZ+n
yxQtLgeTmq8QE+3UhviSKhtFocFq/nqqfed4H3Q6KZWVjSbxqxfbpvhSY1p5
Z6uEibNXbCSxICWi7qWMltM/CbFb0qVVjK7j+sLhbQk74IjgN1AwLhqYkk0K
1xkFPAiHx5u3OCXMieuENHuNrhAXZXi1MdnNDXWIt8JABoqlgW8T/Ja7PBq6
4lUVXBKoFunOAnYKVOJ3CrAHHXvIqMhDqtM7iwjgPrXQBll5ehsffj04eYXk
Ku4THPu389RViaqd3ZOqKjU1koJEia0+WAExBUfXpCLT0C/2TER2eLs/yVtv
7d2yR1Lht+BR086FsdGi9WjdvaKKi8zDNtCZ2NrbZMFMTgnuMT63DWGNO7AD
LIpdJ0pMFSwJtUQqZ5orj7sJ7zo1tV/BSv6et52FPeo0z98N+80KwpzV8x/E
2vjWy9q6M35fq4BKeaYj5EZK1t0hcmeAK13hrpACHb15w2lSRU4ZQrNVzVPH
bHY3fHQFXUM5tU9mOe+nbxYHAo2uanzm4asVWvW1+JF6op/47muvfKyQlmo0
JHFm84jaU1VGQnpR7eUO9JTidZCTmkbd+9UIQUimbGq6/C0oa3NZbynnav8Y
pugD3p0y0xabIhkBJ75Zlqi2AcAirImrauQiO8PoctvdD9p6xsKtKZpBpvhk
HX6usO6+inUzR7/H3LZG6vPLxB+8x9npYa3ZyjB2pY/glbxOfqDBrtHXzdFq
EmDffnHf2dIKTK+7uHTpgAuCYLA/k+zx5XA1qoM6/LcCWubiVXQ+xQiPNYM8
7PtHqVvHL9Q/BV7vq38aHZ6i/lQbolsncpQnffguvPDjoo1N1AWiuYaMxshI
GnCrdhfQNruvBs/ZON4NaWKIhhX8IBgkrmRd7g0DpZ4Qn+Nic2w7S7XFv80A
iROo07xhOAG0GVUQduaRIhAbqiCXuMy+qSbQQ+X4Ae3CowMcoxIbCKZl4JZ5
d+jrGgBVVuy2Nc5avs5xioQ7fBVSWjukdY2xr8zW/2vZpGd/lWBQVRs5V01i
IgtfSjHzwChdwMh3HEXHm5d2l4N8A9E4uBTqqamr04OHkUORNGU9SxrrjoFj
f7fh9Gp19vRqRlNmJenUUYNeqkSMxsY12OL1JtsXmQA8XoMRMIOwmRPETc2G
Kb6m5oRAj4Rj1Jf2ml3RvYa/d5OclhH4qwmnGrg0mZmXkV9MH0O3KseQw3m7
W0IAm/GJN7JF4CDSj0MJtrOplhEOqIvUHyc4t0q5tyo28PIwrHk8mX3ar0/8
yzrYWivs4o4VgKBQQSgHbBXdWqYp7Y4taJ9uEkpvB/Ex2CytddoCFG+OZG1u
u0mH7s2Ym4gSW7ocV4fzEsSbMrwDRNTqHQRKA/8uWXiGx2W8OqLC2W+s17BG
WhUxWeVB89nnEy8Zdbh2Dua58e2h6eqKIuN/fZtGuIgiSeIZezIwI52/amwb
l2tUEbXciYWYvqGcaty7VCwe/GDmRk0onw7PDbhAh7TLhYk4tAvsBwu/+PFi
p50viWkMPKF4F6oY6nBQ3s4wM+FpNGWomCLndkOTJE7dp6lqilWK3VEbZ0HM
1CFkg9VvOa1uTQIndLQdel1O3py9EMvlYn9/ix0oT3jxWuAIdF04cU7OhgFY
SkOBOtzLzKD6AX3ZG/kucqmbzgcmQNBCwQUVCPaWHuStflFABsZo4ufBCfko
MSnGpISN+vcucsQoTFi5pdqmycNvPb+8gffXJy1LEVgUKYQp6fElqjo4RrcS
GTdr4A2w98eDtIOgAa1Hp1oot/MnKHDSwyKpT3WsVgb5y8sStLSCWFvhJivj
Yz9TxYzxVbIBXMoRxD2tBqe/jO/etNSyYOiN//EPcljWom9aJwXB2MUKmzfP
qjxeJk8OfgW8GX30Pmsxk2bPFHbxeSR9LzbjS9rOY1zpdVakI1pBTCUbbzKu
IjUrfkKViqRowNJ58G7u9KqEa+XZLnFCCBD6dp+JWO54JfajtiyLXX5L9nt2
VGU8+A8he4sfM46NoXKrqHlqQZq4zgEkaBG7/j0KdxQ8sB4OjFwf+VuC5R/o
8XB8Yfa+TGZ/eV6vlOZSDK72axMgT2VP2WbEVt3PjqOKeDl+dbwqW6P0SMXO
QHdau5egp6wCoqNxxE1ZKGb++AueKf/eb6BIfzUC7hVVxjhEAP72fromjE/Y
91lG7A8Z1jQ+lrhgUUNe5AiVcuLOfm7y3uzzxMTSd2h5xenfSmx9Gh0/eKrP
oZ4mFjpHhcM5/SKGsUTCN0s1iEm/VnI+dUQUtf2bmHzj35SAlKStqn/cCljX
ji0j24LHmSotytRDCuE7Yi1jCU+otAe27Qt8n/JBX7Yi8TjGpYoqKk5nFELg
BeG2RQhseboIbYVX4VNxzuaeXCCYpLFnw+OSw5izsdhEWo0/2OAP8QMqEqIc
qe35MEcaQgZy9vuQrGV8wEs1/A/lBwSSUWHQvsuiAm3jwqvNkwoL3kfQF8sw
dT4wlfyJU3lhTdCh35h53zyo6K+TUtj4hvtNdUPT4d9Vdb5ld72ouD549FzO
BnDyyqOq+ei5M5gdVeXg5B1x4T2wizRSfkZwdzDUW5H8cAqn6XNBCMh4ZiTs
eNWD2OoVLbVZQN6cENNVuNSh1PquBgFwmCRCygz5w+HhqNmBvnzZZEQpPOex
fje/j5Vx3VP393w0KEXnzoq5+CUsKWO/f+lIEcHEkMvFzqn82+iCAjYbZX7+
kmaMtkfPCPKrGMU/12yYi/GyqLIG89thYe6NurNwmmF8tQhul3JuaVSxd3R3
xeOFhF5rcOw4Q6DFDeNsocpB+3TzIm3ejEQ0gpYvxi4e6RGP4VaFnIKzqUCw
Iatf+zSghuLiSgdGh9RewvkJRYfEZ4kKctz9fuRikl+ibIafYTtJRDOyryFq
i/VnTeCNa2GTNysedwElP0/AUl3MwaMh41MmuWnBfaxfi9gw1HIqas4H+hZR
as5mV7LBcjH1Kf3UL4Ins4CSgUzqJ0RjWRmIsFEV3qjV0nH53Hjk5xhwfdgp
jUxi1ZRsYRBMW92NPQhHZGL5wrpn4VQI/Myj7mt4N+hihhqGgJaZ6XEiC5V6
3IvWu8GayQKqNeH3nra2po0Dh9itulqDTONY41pRsperimqbyCJcHjZSV+Qh
oWxQIFk4GgG2Tx9ro2PPynCQcGLvClUuIv71M2jOUTdB8I7tQH1IejLXUF05
wB5mJSp5kLtsqyhU/Bf4V6Ie2Z/BIHbUMWTrv8z8pymSWmnN655i4Kwgv6IC
m2C4u8aioLhpoQSVJGjiTbrm6sRP1NTHU7k3h1CSMrNjYwIpFJPSiCQcbtJb
uiWIe1PrUv5xIatk+Ky0Thu0j6uiTBrztCJBhgWW2VULnVnW+dapgrK49qgL
oomXMKjXS985d8uZVfzEzZTPIowFrq2Ms82hVeLdX/d7YJXdgLdZne84pgXt
ooW23FV73XSJ+T3Oy0EZl9CuUZzRMmRB8V3k/31OHybXVdgQvQTwo/eSBUqc
JXTcwk5ruc+EYVNhiG/SNhQ/iExpsAZ5VCplBgC/hYRGixS4sOXE1xe5BUGo
rArJHAUEzozy2tKrNuuRDAlZkf2ftE4cYut0l+SvGrFW2HwG2XgIIzobyjaq
CsxxtEO81Fl9BCMpIusfEpqJRbH5fX1geEr20fEqtTBWxfuTWyc/McL83FiA
KO6GlubB7p50Fw891coWXBk1BsQiG6bz1a3sGWKwqN4K9gHAqibD0/AwJn/s
afRIVOZJDljy3MvAATOXOKYRcXWhpOVcPsz9Ba12UQonHdI+CmKljelaxRcB
lWNMi+QY64QUJzfT+x39u51M2SXFw7vBCTcWyej9Y3I9WEXO0Dug5p6jdrNO
74G/4ryMbOlExqIXaCePS8XUZozQ4a+l0kfNIKFSnpDvsH+cNvQpEwI5Uq1w
JIlE0apVk/KMbU77bd3VpmD15Oyj6LVR2iT5BGcLhTU+SOeCalfvmvWZahfU
AWEiHWmQKFuJDTAoOpIeuMSOUuUkmmLYCG+SAzVSGygDvvWIKojR2b+vmni9
TuIu4KG1zwZK5MbBsMER8m93QVwU7ODJ6aUK2JNDo7rq5tGPw2P1nYgMVS0K
+5qvHB9MHSXkoZXMq0sZL0N7RTUzUU5WX0oQKHgQNvaoFiT1k8oQPbw0UGhZ
MCSRWEMwP/Tm+lAAP5g+iCZF9TKZWtEnKMQvQvn1VpjfgcTx4IzR8vbrEFoA
waPWCBAVqbnsUijM94zNDLjHcfzEChiI6yn+Hz/pba0tQj03NmVgq4kVCQx+
KMe/OhYKNhe0EeZRzaCut3qjxO6DJS+hxeUC6hI1ofmLI0HVdazlTev219zF
GzEwP6U+m6R7Vi8K87QdMJOqpc/zFazx7kIRiuLxidRdgPv/yzkqg1lxwn/q
KtCCsUl9sas3qHAjv5Cltc1Krw7wKFWrWBYGKJhpYC76nYbqI1WmpGYINdXZ
2Nqtd+CDoaIp7o6m03t9N3wDEnWgAZfCgQYkWEvJ3sWcClHiIW+k3o5FElJE
KZ1E4W5KDReMXyRR4FecQQKd9u2GdgpzXXOijWJGIEKlLKPrM9nwXlg3vZqj
dKkOm1SqIdE9HU4IXczGBw/AiEXnPMcglRWpjUcVZIGSVvpoTEzegdUqGTWh
o6bvR/0VEVsUZ9lAPKi56Q8kcizKgj0C7yQfiL2j2k3dPIpQPPFFvT8Plfe5
nC8atCscJc1nwoaxbhwgQQp/DwxXIemv9UGHlZxRgvv6G4TufkMFrBNu4lp+
iEZ3F5V8Iaaug9rI0I++/+CQ9+O8QnZz+dHP9O+EDuK6Bxgu1HntFOPgadaT
C9Khfy2OvNC+GJ8W3qgbgAodAfHIeokkyNmEZyeiN0urqlrXc1FomYqSOgVJ
WXbMbfQ3ZYKwhtz43+viD0TNRNyIQkrg3A3M7WjESDqVoI46ITuz7fqjrorL
QPI40+lwYwWaiwQLckJO5SynhUcGfW/NqmYx1yVRVqn2KDIqFKARHRq/wIu7
xrXpeB91Roz3isf/EI+AmtDK67oM2PBXRe9x+wgFVgl2D+PZHOdBNZOIZBWP
vh+b5yvTMY6AMxIo2YEkGYj8oFQtnVojUGiRcTt+RJBl8lDOqHDRUbSCvr8f
AzNkg+ng9651HVq6itslLzEewAxJxiGtVRnFlHRPmmAW6Q3/Iogb0+pKArue
SkjMywGbzSgfANSNxJlxnQ1dnk1c/sN0FtGie07g8fS9hRD8/8h0qUyfC9Nq
Uyyn7/KMD3nf3r1RH80fq2Acswy9PpI7TeDbIEMo8C/F7jc0o+WHId+4Jf8f
NZSt5/bWvh4sKv9tURaRJecC+sDwRlSocx28Q4AHTno4uefl97R8IgvrRIi2
dDq96FZgqp/8OhffU+PRYvm5MnYYD6CFekJSG2eYrWSwWnFjyQ8O6Emw6761
my8BoJOG1SvyNQWHYqLjRrW6giW1wwEoNJxcRZdwhthSokYFZIKHxWQIdEHG
4baCjxarIOQLumySAm2PbEjr2eNcQQQyI+sPA5ZlpeykK4GBWHYj1sDExuQK
EU7FonebLgmOM60HJHtkjGPEJrvHYhInE76Fgeeq3x0a5VGVuWYBFMkFhTWZ
kvRxIRpAwNNoPMzJc8KqGhq9KVPINgEuPy/1j4rOg/G2RPKw9hCEYnkvCsOC
Q2vt+g35q2vt9ClTun1BrgTWwRwMZ6vwKKS+X51nu+7XVCQ6c8q+h1CgNaDX
iRcxaYBH0EvsJEm81CihQ7A3p0mOEZ2vsTArmedzXKae50YeTGMnhnIg321k
QZYToN1VNksYt5t5TpNik6cKzzWkdEMcKK/EEybGtIWEGzwY9PKvU5tzHv1A
BLyI6pmJgXq3P4v7qg/CMMAUpKeFK9YtTb866v1uVrjq6VZuCU04fpWEyGGs
4HbDeBc4+YFVo0+isrU9cb+G0WGxrGvM4X51oeFeeiuiTRetf3s8fm95QMz2
PsnU1hrptIIWZomG00vjey9kFBG/TnN9Asr0laxGKVhJDGb3ilK1IdykVqhC
D0RVPjJmOE5q8jWSygeExl2xpbN6sDyKgoqFBkdyg1cYvO7kXUxd2vXFWoEU
pWC4EMwi4fR54VM7MSqtTh4rgLkBkwWPdvO7UCFGCnpnJrSrnt3WCf9HZaCi
0nYl1Ir4DPKGaZ2Sw5bl0VSap14gylAqodiyIchmBseTKwy1Q25Oo2dfRQKQ
F0a5xdtU76UInvEwN/eGNaLRQLDFwVUu0BO6aycm/CvSDILAFgpBiat7xS5q
UNGCG1/cwjK2R8iRgqWJp5aFzoP5rW3Yw7QCoVeR7rcFz6btf3m6q64LE1Yt
p/3Z3k9Ad64atZ0CGUjAyVauAgtJf5RzimaWl2ivLi4jP98ffHlFlRWJ40mj
XQraiegbxtb+o4STBAGWhWccycqSe8mDJiPdiOb6hzUjcYbYqHCMbb++K1Q0
FsrRD+QeX72Clbe4OU3jojjFWcAgRoXFfsnm1D6rBByHZmo4nCIpi6q6SRjy
TbJMH+yD3SHuCP5mdV5qflPweWQGdD+JuDpUzHqrV66jB+2M4KAizCmV0sXg
c6n+s/+Q8xGpxv5PAJTGyWQca8lyAGdXZLDLSEFjpMzqKieWkAR7MYbkVY0p
gVd6Pi6dQ9/zCsR0RXc9Ei9SZoR2aIhpMnAsqVTT60LCk85vuSuNcSaArENv
uDjkTqbeKf1QeKXfL9oDUlmH4N5xkXVIcCvvDH51PsfJoOTQJU3vpj7NU57N
eewbFfrFlZNjDYp1GwsHwWeLjfJR7SxJ2NANWNbJarq9hn95MDEAfyVHnOIW
lfxaB3vz+NwEyQo+bNKp6QIgWXIgrUaSSOPLoHGhBuMhcGxQB34eHlVq1pMU
xZ992bUuM2O0lrBud7POpnGxR0315AuRm8W+W+YtzpxAIjYiJ7NAHDjs7OAM
RDGMdfD/VHGRPbjKQZ0SuCer1AcpA2bgjsE0EmGCh07HsP96f8o8fjhhqWHF
WiWzK5KlZgGlLOD37tBW7B/n4lx+FM/ZBX78CJkPVg02LKnWp9ymwl8ppdmQ
LiJTudD5R3ZmucH4ASVLl79lsbTfH4NKcouaj64QHF/fog4HSg7yerOhgqUK
Ro0XLW5dZ65psdJgfxnB3M4wLZiliWYu6E6GIO8+ofed6wJ9DP77lC0VE8/I
J1OaKbTAIeH9k82FyiBFPTaZIC3R11bbKFlrGRldH48cYXtS7VpDB783s1hy
vfkesQvEqA91/pnRuhspQoLejNafhwMqJXMg5C9OvKckH9gGItUQWE5ymWx6
IUwiA8ATNiY9Wxjl759g9TrKURW3ke3lamCvFhQUL1nnU6si+SmLJGiYxA0j
L9dwy+EaNdeF8l+yXhO+nQx7sbY6S8vYqt8agKOjVgijHTSnzGEmKtNiPvgq
NBthnvw204y8CXHhGPRiDLlLv596zHWZlTseCRCLCKd8a3g1hFdGI2TDzaV3
0fPTR3lcVvBC9jd6KfioST2aPvas/AbwM26Fd/K8JyfE4Xy/RWJv+hsL6VGd
4ylviZVukdPIUmpZKM7XZNwfMPsPNcQtRrgR78acWRGudGaOwO809Gyv76kZ
0jpfn+cHkxzvZLC6TS8Ut+ze+suwI3JjYZQSNCfKD0DBRhPpIrKmetroIW9i
ETIUq5hTs4S8nLSpz6sKinWncJmM4tsR4u56EnCp+/nalKQlEn0CheqgwkTv
O491dB62XMzE/U1Esotb6JC5tmISrH4diJVxeLIPL4DEP/dQRy1E3yQXpB+C
KbEUHn8ISwEiWFddWhxRKjtQ17qrkZXCSpzievis3EHQfr7A8Ai1RT0ikQGK
s32HCEWvTu1dSxFHqcqLuiX4ywwV6yX9fxOSKttJweZkDnBsLmZMNYR89v1r
xECjUq1lkkFlZBRRj0RUKqtqWBhLDzAV9aooAA9W5jHnnwbnIM/G5EZP67Xn
imjYKi2XAQW6rBt+xbh1AT2cKZlmmJC+8Ka27fMqhNVcXBb/SaCqSAVjH/zK
zlUOm5Ufw3P+SBg7MousrFCPKpl4wYTDCLkOhFK1llxp2u/SQ2EfB3XDb7wN
yxmBJ2fdKTKiuekdOcWQxkzHlnHUEjklVRRALndzY4/t0nkqvtth1iF/NlkN
UAhPRpNN213QcfH5URbUdoGDSoAutzMdez6zkly9G4XOXvtu0yBfdZTWG5QH
NFBygQYJl07HFWbwnEjpdqnay8iK75vBWUXLNGtWF6gWQAi6g953fcUtsEsm
mVk/pwJCWCbp4d4nXJ7yRmAMqwZ78MSDXUSwt6uP3zMljg4+pD5ba83nuJhx
RS3jemV2AiSv6qONM45nSoae/8F6EX0PEDP1Sdpdd3xLzKN//nJQ7SfmgYXk
5jlJSCOM5sYa+aUYGP/Pqh+th9n7upKUvOkELdoA+DCmcKDCKOdkcnezgjCE
NV7CepMzX8UwqMAIM6w1pa7RAD2bcX2ktqryfuY/pkAbvydZtKO5F28zwMkV
SBINmeSSDMShgYFfnwa92jjvV1qvbJvVSl6u1pPVmbpaIN1pH7nbIQWMJwj9
LChVxQRLrsnYAnbBy642idaJKp/mk98gN53Xq9sDO0iXq7uVHzKXF1iaqBzx
/f7O2MlpOFEydbAfcXxHvsrSVv8onGcHKUfE7WpLu4sQXhrkHZFjgJRIMwO3
XCwD45QiAShTLKRAqZa9wOMDNG8vfJ/KTi/qcLX6Z8hV7E8tfP2a291C8+oW
m4zf4Qaogu2DQHj5f7LwvOBBzL3yb6ntCSu25USzKy51o9xRzrQLuZx3GZRV
f8DBvwz6bTtLiQ2spzSHBQXWzW3xeW6L3KYhTafiDnbm2HdpAWx5mdtK1yJJ
itOGV80qYjLXLqiIsNwKp8NyNCpypOcCDYT9XTS+jFbzedr5CufWbsAIjOUT
F//c2lJbL+DydVSB/lg2XoeoC9+9EaGzEpJh+OYg9kmJEr/14M+CJZjKRedK
4vyqdL+cAWnwyri1uN7Ifenreqypd5iUh75OM+ZzWLY1x3tbGGQalARElizX
AYbrz7hFuYt453Ij/vYsNy3PzoSypKFiTt64NF2RBAlR3r2PXfv8koOixGvQ
DvmafYNtcH12gYbLeV9s4STqTsAa4ukmWyPWhyYEjQCHhq64E+CthH5KeiM/
TwxuJNU/K3EW5/mNfYGtxRnbkMYz1zK3VwWxYqwYx4nuBI+mB8kHVPOEjNXA
fSLCzqSrm24vOvCkkcoyBpCxOY7yuVxpdVweA0VYyit4QRm47OP4S8ObLom/
R/qKGG6++uNWL4/5c1zrihqpbwxk89DPsLR8yaFzrwdcccIc2XrGyUEAox/2
RYJLk8Cq/8j8pD9+1Fimtmd7LYwClLVB+xkkRC/dMtEoV8+bbUmAb/TuT2ij
yOcvAI6fHBikETHX/ISQHQopMSxkAX23cW38OtcRgV26JkNUI0hmDalc0NxI
ATxkui3dOwKC3l+9e9u9sQjKdef5NAL2eUTUre5E8l1/tpBEPGjKPBNtb0+n
iluY0S5b92dDAtNJ/8klBh5H8CY2Y7YEJOdCbX/2OLWU3+np2kde67qS0lEL
dTIrrW9sIRFUjywSZb54oi+XjaBM3yOQnMBX/eXTT0UQudyPTFSffJ1EwHbN
RcWx1aVk+30NU9IiFeIPLsymYyaxA8AH5cFuZvbtDM+B6JsjOSc7wPh6+z6h
ok4xJn0PQ0N/aOYM29E2is5RIFbrSQaaRS/ObOz/h7QCnQVFumTh4yA1x317
I/sMaILodNNKg9Dz0eLpHymUG1ne8rwvPQTV9DIz1fB6ai3NcYMNHBLEI4tD
TugvSfpDZCbQs1pv0bh5nLiV6SPlLkqfxeEEeqXtulwTEVhHnJUEuj9ScKIP
ykWnYGJopCszfoIrafGtJ6RQl3mfiYasjK2uzTWJdOspdASKAaKmvt0BUaUb
O4ywq7WhHb2t8xkjnKn2r5IB+qQbpEP9CE520gh3a9aLV4sZL/L2C01Wa5K1
0UPyD7pR6NTr+9Qs/pr9N6LFMl6M72JiSKQDHxAeEVf0XN1tww95GdF4Yj2r
09FERvIJnRsWOrA9LogbjnYwHCnJNMqpt2WYhpkFCWpvATnOJLE6kWoLDBu3
F/VWtVY7u00eMLckloxWnH5D2LEp2j5dWZYEmm7XZr2pSXpdt09UaK8d+4WH
3pGhKMCh4UplqVfgTgwofWovqhkOaYE17zcOKytEJbhGqbtNv0zJa/dEoYu4
mXxhGV0UURjSRutVncr9c27VdL4c9cBpTMJY6bxBiJLMPpZ7J4st3W/sVJgm
X8NtpX4slebvBxKFfrrElce946goksTFz+Y8diQx8kPbO3qYXkQZCr6qbL9a
Sv2m1o6WFFEhC+HywxaC4BkNe4fH/Vemk1G0TFlec3xilxX8GqSBIxe9fk3r
nBs4SOwdRz5yoi7W0BNcBaCIsbKLpgBdwYjuI3IghWO3M3k4NyjzSH634Xj7
1Y7QMdSeZsiY5zqcX4FLn4JP2yUuB+s7yMv/0EsTBpwhe3i/RRfg1fiu4fH8
/4m/3jEsd2r3f31APXIJS/zehWoFUgWUerrfrpYaq0bQ+oow4jQRxlAJwrp1
SBj2DhtQkvQ9MXxEcIT45qMamRmQKh+pc57dP0zyGdbelyVoxhuBr5eIyhcm
QtJ0F2O76Nkhgd1ROCEDkUwNaLeU5lpL4PamGVbQRb0Fp3z40QupezDjS7Y3
tcdOa7STHnV5Id7tf/hI4rEsEZnN5iv4+PKYIFz0dHYuQt5Z2z03v3xoGgCz
MJmMOwmKt0qq/m/ZrHEc24o3lM/7vFAOjVW7tGGg8fe+ihSiVlchxPnovYSO
/nchTgND+2JWKGuEEWFAauxDWoEtG8P0SETqpREj8/+hSHwnstIniClvykLD
/hSLpdRiV1icSYYnHq95EuPDJaJ3y3PXCeoUHanOElk6pLlxqQNq78aXquku
gK8ZG3e9AZpmZrcCnTbKXG+ego4fuFLUUPPLFGqG8fRBcPM9PPvW+aTgIHU2
h3l4gH47zeEPcvRV1dG4495R07Wo9XwhtoRL8xVQ9XbMVeU7MY3xsIYPwPrA
1K4eiljtjx+4ntvhkgi015zvmBoprYjGvcmti6a1I2hsusk8aZ3hqsyL2BnJ
6ff9OcfLlWa2PvK6Gq/CsWCcjJ6k9pD7Q3GFZwolXh2U8Yxu7eU4g0vQIeUO
K4ak/bn8+gdEaI7Pn8EkcHtj/iPYbjRIi4ZhDauqOGcPCsSi0gYdgs34UaH/
/r7k54LTmeMj2OeEu+m+uQFQ0qjjUPicU1uIW/F+E7l23PVBPciQ23e/BzVi
xOSHjB44meKwR1uyQPEezUCTLk/OfMhA9zr5CXu3jNj1QSbb4rv0TNp4E9Ox
dShRO+HqVBzWAVN6hJsjIB1HricURZevWrGeiD9FVe5rA8cq6WnwLFfMgWeJ
wCbG5BvsJuCWhhPQo6QCynFu2PPPDAUal+IZ2fkJJAS9n1n1LijjZW2CZJ4C
NAH80WP41E/PceDuhHfzz5Jgb4jr8FdHiCg64aFk8ibl5X6J9cgfw+XLH5jt
RZ2Vc2Ulnvw7AmGR0agO/YEBFcNJRqSLcsmr3p4AiUfpRD0Nb91yYWFv2WVb
hLWvZx/Gyva08pH7W0iJ71E1IrDF5p76UCxxQOSAi3TNkttrk1EJHK7LpDbU
g4jhnY9DQeC3aLUbRk4oIeBU9W4kr+0OemvUwsLJnqPKrr3RVKRxp4gyp6ru
XG52u+cW6ttGrrCmLoMPReg7iLoTROwQPSsNf3UGey6iorJ37TNVpLaZ3iRQ
pzXcOe/fpkIthzOOwaFtner4TdD0DPETkDyMxdqtFHhZMNruIGKfiV0Byy6b
FhrVRVBHKrrc5Osnx/3A7B6oE0MLjo3zADvJCPkuSZAgeR0fhLNDvZeVCynT
v9GYZsQVRy8SvLjbDiPhYSdBFrgzzFPKk2HIbatpdhAikMEKQRN33ZET+8Iw
HXyr1471ckq3QivbqbocHO1af2L/2kqeAHppWe2kb7NTzEhjub1DBzY5NHlV
nfxhBYGXnt9ON7t999+4bAW+xxSFEbdIvYXjpI+ZzW7q4pUdk/iHiDG2S2T1
xzWTrRf0oYXrK9qgsayjgDmL1jcb2TQ4FtbOzFhRE0pjUoO7mSgVnfZKT+k+
9JS8I9GxMyrnP6KyopBA8MvPkYJtX2+XqqwkWM1xUdTJ8ZFiykqM6pdZ417G
07lVWugxrhqHGJp/R6XERIEOTFeqwX5HNrmIhPM53B7k3/JymJqWzMFIyx+v
0s2Rc9tq4b9CcMZpbDZGwp3X++Xc/cJKqjxPnOAXcfqv0RLYVWNXh7HngDY/
GKcOmRy4/kOQ4FpeAF1cXBVUbNtOlk71yspylGD6Qp8X4BHTy58UOLxqxke2
tRHZTKgUtj0KjS3YulMu2mXGrR0Q2nfe+ifEJyXkYYYPYRYLm2Ar6SvYpn5e
ki603gpv9rTAYwF991n9t4Ssf8XNqgMydS5plQi30DAXZqfqT5wLyLmZm7Ok
d+V7CdBYgEFQERGCXqLRBmjHIhlwHwrVF6hyyDH2YDE/9TYzY8znT5yJxX8A
AGMoQENrmPIENJvUICvrPCQstI1r4y11Nr7U0tAWRwvaVbMafefaHrudEeFe
3etZdHT9Ep3uL75d5DSm0wZsZEOac04Jiavfhf2eZPkaNzCqZJZVEVWw/fao
jWwEPg/wm5/T5WOQo6VDPar+PCwnqh5a0Q+NmaYkYtbpbJ8KhgtAZZE8WXqP
v9KB29PSINrac+dnU7V/LvpMPyFm5iiXYFhkz4dNc8uczNcWEjkFURINiojO
kiN5outNzxHkkAjFiJAR0QgUHmcvMJlkhTEofYWTBJXYOPhQIECR47DO5rl7
gRN4ftqPB5e0RapcasFH+sN1+a96R+IkylSS0AtPct4t/37RCMGsWv69rscy
fukH2krXpYzpW325hDXAK1DCnW/RH+TKgtzSs01O2vMwddzQD5tPsBd5A+lf
vjdLq20OXWPvemcZHSOLqBs1lejNhKaL9ccGaqIseiOjPU11AkdPLPWz0gbU
T5nqHqyRWQ/FTodMf+dLWkn95FoEVQnknbprc4GoYKMQQf+vJZ2DJIlOa8Zd
+E5dRdYTrvA0XVqwBN4XaLGaB9mSFUjKueB/MVyFNn+L2/BfCv3FythlvjmZ
z3J5O2aBRSiFSCrsAZeZr1PBTQuxQsufQRcqVu9ZaAwViSGLIoJfJs+6mFAH
R9wMt3S43673+uWZ0FzIvCss/RPz9LWzR9eFouWg3OVqJCJvFbcYS/NvhKeU
RU1anqdnbNrfT9jlwPU5ZcurTMjzmnv1hf9UcA28IwKTxCv5kJlc6bQQf8Fg
0fM0yfFdCPrXG4Tsp5fmHBhQsZFIOWibJz5BdfcfmqWSmam5qDOJuXn2SsIu
vgaq1zteElNgWQTLCvH+2zQBh/mD8AyF9hUZXYCkD5wGF69dsia+z3/I7AeN
gufQIMkJgPqLHaKYGLlJhs2K2bmE/lf4z4OX360vM5tJpJpGwqX1c2ilegBX
FMmirp83Om5X9SMjLE/KlQeZKdIJnBk6tEEmHIPt79A+/b50okws24eP9Jhf
Q2d1GJpsJZRvfWjSYn5rL8DucSdV+OwCthG+CLkmnBD2EeRyqFZ1O1HfDNgF
BLuXJHgCL28pfSXfCMS8lFBvOicWhJMHq2xVRitJTPWTCxJDAlwa1MD8KIYm
gJZumBUs9rWgXSNy+xINpJI1UwVQkikJ3c0dCNdGlU4GAf8rp/dYDFrmRJ/N
zVgSljANweKYKT8orBYpyr4NHSqum7dR56yXGjBRAmkxD+GFi+f4hKR/Fu0t
eIfqBgXQBiS8g58FiNgf2TeR0MUJwjiLWF/yl9Vxh3Mz6ypTA5QWjPSLWFad
PbFfoYN3RJI6wvtLk+Z3MY03hPN41N+MSgM9FU8C01q99ta2R4yU64558wGW
P49p1ftzwVf2vFDF/yaviMHzM5ztFI73j+WPpi5ozFHZryXOeiqGSPg3aQ5N
WNk3+DYWM3h0RVetnTG8pO7ZCl2HDGZsC/T/swaqMkAetQKyac2iOVBrbRv7
Lq5ZjXsuY507AzMhdwVr/md4T2ee5OVaZ+wwJJMeCLf2fCBOuCRm1M1Ypx4H
8++vYh85OR4/yaVvFcw4YvddWssoUAkgWCEqtSDmYJnyacWrQGlrjFzemHu3
cR2U0t7ca+EzR2RodPMyAgMpL0uWYm7HWrjnbmiekW5qzaNfcLXCzQUKuBg5
DSvGuR/VH9BfTVRSGq9G+6kJlg/9iF9NJiT38ZOHJ9yJDUhUdfsFVLQ3Vf+E
dt2q2Uwg5v1Ii0Spfp75iWt4EbrgXM4W8Cm2u2ogl/lA2e5+czs+FnoLDzNq
MuXPEKnq3Tt0FJVN8tfLITPpyLuFR27wHEkd3CGgfkaH5ev6le07nuJS3jcG
myrhIAi+bzdnHmtOpOlbWc+m3vjsRT98+t1NDwL8kIX+xCntALr8wVqaXUns
LrwDoUowxypfwJhFBTO0vgrnClJymyC3trL5uFWNLunKLMoHA91c40I9lMpM
Zad/cqSdHr6tUdIIsXCbGoxVMhw/kzL/BmBrCRgcs09RJy9umQ4h93iPBwzj
rp3/ZsOAybLIVaUbPSvh0a8Ltz8h09F4c6mOOnDWBK5qn3qT2kre+5c5MkT8
8r3WLWmNvdx/NoxKvS4PJAA1IeG7tRVPZOGGq+2gElENC3VCh5ftttqWcOUf
MAY46mLC+jsk9nyVxgLTwu0bMy6vSy6E2tejYHRGLdXu/QiMxtMdDOOnn/Cn
lo/6I6NCDB68h6aajYrb+Kaxc+kXfft8fGTubdkZAGW7daM4+ILslnI1PQJM
U0W0B4WULf0U9wqVaFpfGGfTIFaZScJEvTFH0RIBw0t5Km+Wavr/fXo7lL7k
0P0+ZhtI35Q0Zvx8RBeFb30qipqP/r98gO4YQEzmOvbBYVBE5pbK6h4t8OFc
lVnHIRRANSZ2Altx3zp9supooCCxNJtmZB01lpEyO0Bv89C95x5xtvd6SwrM
+aIKUVZnT2aYmA4FvREpPZUUE3GhWQxQvSBtzCK5MKxke/x5bIRfbYXj8XPi
GKXnt+v+1ZsWcwD98htnum2oS4Crt53snPR0ooiZ+pYpKN2h6dEMGiaeiVI/
H4Nj1q/Euh+l/TNEkE++TYCOagN7H9Kgf46R8CQ9Wdp3uvUW89YyQpIEle9h
4Lqtc8kOIuW6usm1Tk5F++yDDYaKVgIYs6+ZVmqjbomL9AmLaMAS2Hrmt0CC
2z+cwSLMffNBeCQ6H+hZhntWvJZLWLVRkZcZcviK1RttfAuGuNfy+TIiBEDR
vrYAgRptRiQNEw400W/lSV9WVrGr3666q5xtOtP70y2R2xs7A3B1WBKnqWLN
KED6hPpgn/nXQp+QVXgt3p9UWsBsysReBPdJ38dPOlfzG9XEZPz6miJU7eP7
+TG74Vc43YYUYF+010enJ6VqvX7OVzg5aoRGJWeaRE5Oso1Do4JULeJImZkZ
as1yxr8L00Pwr1Y+3xxxO/GsJDdeQgdPEPvcmIZMzMqjyC+T0Kszk/lQmq9/
HH4u9ez445bEUSNwRllT+OXLBKPP2vC2G+xlHJeyLOJxkkj+uO5Wjm/qN4rI
jVbAkoEhZT/bs4+5QMtFcARRepZgy8baBBYEhwPrT58w4hlA133KYZpJ0Skp
t3hvQ0DdIh+HaNhZA8K1krVWMjDanJGwizYqp6bGJLr5GbKnOyA9RiCFuCzd
Aq6B/x6L6/jJ3soQu62O+J0LiArG5GVe+SsE2Tai4j+/jGVG990iUm4A7EHO
dYEQVon/pALlg1Fc8Rn7aFoSX4gZ7EsdL5eqEu05JeGg5wexrKNYxn4qbZcr
D3Ktv3rDpOG1X/0ZAWNpNV86tfDbEYX4drpNpZ4ZPN75zuNIeJ1SvY8PRQS/
cZHyGWl2D1i0xuvvawK2a1RfXFNWjpb+VPEQ6GvgRiO0dbmFDE1DXlmre4zP
OkQIJYLY3zg1Bo1nzGKKn+pdu7yHBY9uaKyxHxIoRMaM4KPAYE8XkvEeETCT
Loi0LtVm+DIvlgCt0RbLMR1qmh4v7rxo85rlkRrWVd6omYPHkF4USzWgm9Mu
WHzQS4J7NORR6FNtmLpe1Q38vU56BBU2U43Lckv6zkkknsOD8SBrbVfiDowp
bfPfJxoTaM26aWULTLAFlC4EWlVNF0UwzR7UudFtQ7g//PYyuwI16jeGivh1
AUzzaaMs4zMQGRt79LwhtDw26KpXuKtmR9ujN/3cwpjDd7S8BcNQjp2Ao7QB
zzjrOQnBCbTov7p0H84yMve3uT7v1haJaNNJXwSs8QorkL+IDIwxK8C0Br+g
/815FkqCYPeb/Ot+JZzbNAPe8e1a8q0UJgoy8P/3Mo6zMyswOWrRs/VnHA9C
QfmlMrQQQuEPXWj4JrgEGXeNVEO7YpmB3YTewtBSfiPKso5k2bTijmkghNTh
kODUhw1hPzdcEvR35hmT1f3y2h9xBP0MzwCX/BMGjVtJf/HWJH+ZgKfQ6x+O
6UbB1Pny1b24gvBmD9c5hQcwkkQY9PjEfwYztp8JIRithqz22gbF6ixZKy9K
sCBmhYGNbUpP/X+O8Pz0zC4Zfm4Tw8Az81UHCCDMEMbeZt+A/VUmySDFsHhA
aEycF4uMxGmsg2UXfTB4dYFfWneOvRrQG4lMdvb9+s07YUVotYpexco9yFAD
sXA0ZLr6+4n+h4SkgD8FVphJ4tTyT5v3FMcsws2rwqyfGKuoJiuRUl9edLBc
5ndmNh2jM3Bu8Fi9OHIWzZ0zcjAckBfvuPlDD8Czpf2918UX4qKyHowpkREh
d/TwScQtSPoJHg6dEU+ifH0NH7V5dGn3RMnDhYgTcOnSPwOVqwXAqk+92CKO
Z9DnTTrM7iMnhQnVbIOwq6is2810sDQTMoJI7ysOjOuF3n+V3TZUUtdVUX6r
AHyyxTlBQUZZUvHxemWTEFp47b6wIES2Se+/1YNLXuzlPgpWqvwa1rLijWZm
xKR306A3nvskiHQAQmHSxKrmm1MOyktJiABaBwHE19QA/aTVwZQSjFXsA8Vh
pALA+QgtcQXX4z0lOWvGJhyyTbm6bbadjGd8niGZAXDYLeg5iAHmFhEUROh8
uHcQQ+fXb7XGlAXAkP+SGdC3+uFKycXUZPQ78ctZhrAADkGj+oB+2fgDdfoR
j/XYAgS5Io8B/ET+GiW5B9mnKQIO+jZ4p6sDZBBxaAST6lwqNTsVhU5K6pKN
A0PZgsbIb8hl3e250uCtFWkHdgE3suDyEK4wAk+iDaj7BsfVq6Kkx/LqCV96
xQFjVyMog5GIejqC3IgVDDfNEoAN335uVOUHyPL+AYb8RYTEs3bosgGtMN4R
XEfhy3eeTJxk6ocmLaOsVNGp8xfQY2dH23SF4P0Gx9meRFQZLPHcG3e9n1el
Ots3gF7sQFu08anoAyhFctp0j7HKZQ8/+mv18mzQmWgnxYNmMwxdD/7cegUM
a6UE2Tby76nuhVdiCeLvIkzX8zrMKaSZV3j4griCgJOfd76QDqE39UDtkESx
wKa6AgfOviXXBLWurl6ViFOB0snU6gDXqcuUHyVqCTTIT3WmmTrOl+Vp75FK
fdnVkjs1Ks9EHjol5EnEFkjKwT1f1DgtqfYxBLuF11HfVWGrsNwFsm7h/vi4
j7a8JOdt0hOAU84RsMCPoq74OYWMWTM5U0nniazUixuU30WLwPkL1mxy6nm3
G9Ico3z1rceEgns7Pztfg61hMxASV18qu5Ar+DKEVzBZBYkPjckCCJKUmvBL
sjKN0fkvWeX8fpFBdATDWtWpDOeHQd97jybrMjsJFDGtK61Poyh4w5kMgvd+
yZodFIlPJon6kpBHuBkOVy2xejcjkvXVHS3zd/mkYYZ2O5fH2PzMBtC3bwe6
dzNrwqw+WyTblJtpbvS/vm1vlCjCssPE25fF0UlWxEMlISkYtPnTp0JzmYXw
I1RLcUijcHu35QDZ0bkOKO5xaFjlgyKLKjzB9+Y2ujUb4vBx+BO8wmDy9q2a
Uvpx94+hJASJKUS+//VTuuj8xQPhHOiZYv8IJkInJD+c/xgzA6oB/ZOmBzIF
+v2jYpjuVAZ4bOwRVLvy4icvfRcJtw12jt1R9b6Daw27gDsSfOf6T/c5mkSu
iiVenLAHmBDVUcNEchKc9xryD6npRvi9AUyuf/dUnoOgoOCWMnpS4XfaTlIc
FiDWf1bIreeuuKWTIHQOY7Qv+tlixWt+cSloeuYLVbgWA1AT8eZsFw62aXuF
dKpUK2PH0kwAXeC2btcfAs4iI1vT0TEHA2QPg/MSKR/A9ocnrqw4xeyoztCi
2yMSVARKfzKy9U+2efSWPdyvRVh3BzjqviEI8GeZHPuzBSq3KAFiYbcUyrml
IOfSOaQFAEVBLiDSp2es5THB4lBjYXYjVPhC8BM/zs7iGOmKAaet+0845yWC
1TwbPRWpwImYq/DCHH4uLjmTVxG8BqQtxrBstcIMYfZ/L761xMpiXF+iiQ+X
CWBLB1oXr7f5DbV+qpT7fC/siuPMiggAga3GpzcdsQjH56RX3A5iqmBmH39s
d/tupO0OpsntWgnmIckZvNRuu8FSrIfV1uWC1qQWoopLy8+qsdba7wGX3YMC
FP6r9U65R1/H15cm889/sWy0cpjYmUVQSElC2KppvqkMKovaCWjjHRw5uJV3
0zUDM/Ut+UJBi9WIh8aTFlwmGoVXmyUEUN2yoAuIh1AGwgtYLDHGsCddz4g2
dgGN9IgnSvCGwcWAk0HUbcFShpy39Ym6KIdJHA44hhpqEGqKLf0YPr4Dx+ah
7Z6g7ms8K8/5OlD3RMuduRbT8UF2NPxRXvGyt4yIBI9AiHXpxfBPALDf8IE7
+wPbfi+IkFK9awkBxy9RUqOGpqDjaig8Se6GwmiwSmOVEEzt5SOHhgnpM+fg
l2qPMyPEeNBT9X5LdirWtQpN9BYdocHkjoP0W1b6hdz4Y2BxsSWEfinggeBy
v2ZXyvxGjEw8vrO8qTCAAFFj/+KR3WKSVJskDkn8ddvevHEU0W1g74uVliTq
FwjMDUUIlGGf0S3ml1t6LPMyHq/1ZPMdIEChVl2mPNNnd93QZIAYqyOXxsFW
ZXBzc1O23bx3TM/FiV4MMINLQBT4vfguXYHW3uQtBQshCBSE27S5W3TiqXdb
g/3xAsPpvspqd9n63ZgH21QyDH7zZIFcGl8mdMRsV5Cfas+rPIRBtD/ZszKe
y+FaJx3RI7NrEyUfctVbdHsmEebAZC8FChVswK6JEc53QqU2srWqWHunWPZa
g1ozgmuXYGY7HFryDj10FLFD9I716cqFH626M5jZk83Dvlsf7z4KXnOAlL/O
yCYNA264s7wWugMzE4hp+hf/fQ8f6M4P+QK6WtSU1kQr0PaIl/SbYjohEsXE
Re1wmjEgWtO/A2pXIkenmKhcgpM/K+3HDVyQ6z0nLzlKTfzV6Ur2iu/Xesp6
lCwXgSroQ+RiVz67MtmMW8cKt44QqFaertPnZKT8TTq+3FBDKEy0x/fnD2wi
B1g77Yg1U6h8dlMBGPEP0VxxiZbNd5aTM/T/ScPvPV33RHKeDb1Erv1QIg+X
NBGEWeQnWFcKC9T8p/d+eqF5fjh2vmwA1z746N2nHaEE4mrdqmSnZzuzGRbm
C6aYbDnaJXeL1MvQ5PTbDDc5wB16sWOCTKPz1SIeDHqoeHwtjCO0FZgW530s
mW/zdHm8K2HXT0FQQWVBLPT9G4wbl4YUT3XJYtZmRT+OEDMzkFTCsFBIMwm9
N+w56dnUPnODJlnplQJ41RewpAgLu60lnO+CvJZrGN0j0NkgZDfqege5Y1xF
eptBbZhV6Jxd6QdFt0jjJz5M5N3hq5uo9z6y3B7NttBo3mTgeZCeikjcKWFd
cIHLS7VQDZtODJOg5YGzOyiziw2+Z5TDDqTY9WHH1QS2kqAgPZdscLo45MK5
rlHxtQfOr3LwmoulnaM5e3U2PNHfKwImNSjl6S4IwzZJNqZNUUtPiDS/pCMe
huxRx0NWyc3Q7T/o/zKgRPXCOjGRbG9PzvpB1u0T7QOdVLFvM4X5viqootTg
83Wf4N2wVLqfEPM3oDXbkI/oF1hDI/ohhJkVBsjjtYbmqlzIA50WePWUAz0E
OBacS7Gn+Dk8nmGrk2DeXRpShsh98f7xeMHnRF4zbXg6/S567p8VQxFNYF4w
+ZVEgTk1odgrmTGfqeuJY8rYX/JdR5n0wJVqMQVnrMlOtH+iYYEOnrx7L1/n
/wO4Q3fxuBIaeBrnzXKCPsDo7JeKSE2od9JG71TboHmYuZKjva3ROC2ww5sh
jWexw79agKG/uoyMiUXoV/VRCMHHP4wWNq5vJ7S6IVx4IeA0ikZYZ+hweymx
sj8H+rqo7GNlwz03iZgrB8IjN8CjSp5pZ3yHH2hquM+xtIxKb0dqJXJvl9NG
Nfpr636iEefa/glRmWgo7JooLDWorOhJh9xAJOrIw6eOb0S93Q8fWW0FlUFp
86NvsM0ZgOnRj6wv87FKQw52+bftUP1/hkMh6HHRSd1UW93GSdWa9DeSOED2
Ix5VI67vHr5oA7yL5p6Xpu1vVNjdiTNsY0lxOQDwkU5ah8TUrQFp1j/bJjqt
NkpEy73IACzwooo9yvBl5eHxIArryRPkHKJU0Nzxe6d/o+9nAn4WNoAFenGx
+0G7KVu/C7rQxDgOTXHGUbRNLnmohFY99k4xW/6TnUiZQg4NGNQOqCMfqwnH
fooxws24R8rz2dC1RvY30RypPID3nFeW9xANZcEsMP9xtlGrjIFyYAvZf5iI
JMn2rLLWj3PYhrzAjBY5FhzAOhmfecCzlXa69yb7u233CtgATJeOndqzMDd6
6tfYmSkOhMOlnh5o4q8KHVxn7zk5SEXYKRxV/NIm+ZNUPRQ3gw0Hwzav7NOE
QUfVShbcyUZclaH8ZtPJdJwupFXB5KdpvgfTfQYY5P5EG+8EFTUUzbNJPwix
mRgjn2wa5Vx0yTXJK1eLA6bPoldTmAMCEZoNSitOy6gx9V+FSX0X4uOuhm4L
Prb2rceU2/Djg8as1qcp4o9scojUxF4p/dUZv+Dfm4Or3pedJklYce8dgnB7
dJKKaNlxZcsBGS+H3Kd2r5RgFsxIZq1Hg78/r8V7Mz8wFsfmFjv2mL+aaz8B
rxHZ27MbzAzyL7NfpSBZbrwxhmypTETdS6A150t3LXMpOHnc0sLFjE/yoT9+
6/Rgvw7rJPrEJtOLXr1RGC05SWKH344bAjPMT57ANP2jqYlfRpVctyguW5b7
ZQkaO22HhxD3evaoOBUVGqVZPxs5BaSQUqu7LSSsW/4iZTXlIosC9ieEmUmc
Hv/N4K0qH6y1zuoag5yuOCwcgcbciIW1l7Q+MaKWHfH1PfCFnJGKtxppBzAx
uxpFAzG3vSau+BqUVZGq4FEbbzPsvsWIFsi17c/T167ZhVOm0pUN6lOKO3dH
75zR05hLNeBAmej3oGTmYDCiO/D13eFm/mkDCe4dUAUoFzXrsE9TwaGbRpdi
tFgS7MSzkQ9uUWxq7NZdvKXRaLKIcge5T4oakFGfr/61QFJ46N31czgLpSo+
2cbIOYZiLsYTbVdKD2RG/TsrOfPxVve406lHHUpmJVG1zX9creTJvDM/xsH5
U41fb1uf4mI7NlomGML+3N6K9ivVe4IUtlPu74jrdVG7FZVdrsHz+lFVGHd3
F5YCwF/ZRpvobNq3rxVIKpZ+EdS5NEUQHSKQ5LOoxCGyn5t2QcubG7bv8hZx
g/k/u+TciJ2OrDa5yO5tPIcEIcfQ6jkMyVXcK72gbGp6lap+1LZsr0RmIQM7
mvCV4ikHCb9PPIEYS7u5KqmaYOKw/mA1mzLbzsEmbIZkPRjn7L/LFgJrm3rU
yFSqHqVLuBwKxkh8TpXqNvGI0+O6uIY13MpoLtt9y2ozsfEcK3K7MSiPCjZ3
rWUR1Qq01HypUeVUOrA4H07CantiSMq1SMOV8HRyIdZoFURwuvYgz0IYSryG
TeUNcCyj6C2xDWqhDxMtvvqFV2ZgG7V1byx5y3RnolgutSWbKU8tpA0fO10F
u5Xa31Jjb3R5YXdEoBvnF/G65VsKaVIZPOSNUIB9d3WAuKyVe2IhptQrCMQt
yI6Og9G8Bz4UEttTloyDyMC9NCZBSr2eKUbVr17Tw2uwy0pkJVFZizmMGDtU
oRdjDU/FdObkutYy6EhfiivQxC251jYZ2kd1uacOEg2AGSD8kwOc3l7428QL
zMvx7GeLc61hP8+uHEt2Sjgfo8cQRqXYAVvjTPtjZiK+aNKomcWAmv4wBgNt
89QuW8+E9NFWoAI3fbFCWAj08O80J/2vpveecxmBCxRGnmsUqwieNyqJntPf
573oA4cRX4bfek3j2vAeZCmW0yqtdGktt1gfsVwOxkPr21Moh+MRZIRn192E
2Dh2FnJXRZk+28P0O8QKc6u4Wk+VEKbij2jVlkBGgtom8dBvt/OSWKNV/qHR
a6mNZaF6NMyYKCp/667i085cBeHsC7Y6Ww7qK15lqSqS5ad1MvgH4eJWFFAV
u1jbd3w9cz9v2C+sKm3g0bC+BFMQHoZiRfG3TEW7Cf4yw/mrkgCRGTQnEcs1
QCcDIE9r8DQDV8yqpvpu9hj5SgvF5JSe3tD1wea4ok0979Wifea2LmFyj6Bv
TR50AfVC44o99IRIyBvMn/Rvc4tK1ESRR1S/LNaymmpk4PMT73hox8faHnX5
uwS+n1fPHuR0rXXXBAs9QHlTVJWQHJOejW+sIyY3kwuIo5unJYqSI5C2HIXh
1fuyuYO3a/11yfgBhAkoquCct997WZ6EjT/LHy6+JUkQMu6brktU6kCnu75E
kNWAn1yfDV3OToiWGALnuvehGc12W6ZTjn/cg9zBXLY9pM3aFmfwZSCd5VdB
vpLls6Bt/JUOhyp48qYsRyg2GiQLwS7JhQJsuyibHPD0WQbmu5V88jQJukdF
OOB9cCMWsvgXc5Dq0mgLs7A9zNYBcrAF/IDyaFHi/94NbdpJzY60BXKwamyF
E6JYazeB7ePDmmcCbkBcBpv8jcFuQAqwrygcujZvM/jqUsRPC4bkTGydB4PS
JivM5xlCFAThQn5NnrmLrWGV8RVqMziWVaZTkohzxSkhpINC1skPiuPryhR+
U6y7Z07oyUyDPwuO3K8FDDZeb7dStVw+W7e+O5xrmdTs0USqrpcy86vyccNH
Ztc40CsGR3++Ft3b0L1EQmEd8Z9PuscVm3d2sEr3I3DKxuvhjBEgVg1oyUI9
lktQQ5L3wlmj4nvKxqQIUJZ9KOg83x7LO6bfDQqk+cYZxKcdTEXoz3+6bYNt
p+s0L/Jnf7y2+NJc8QTGn9hobPcy43c6OsTbnDiI4cH2Rw3s5IG/Y4p/D2S+
Rqc9K/ndBd1W2jDW26k2h7tcDVyHPAnotuCsHd3BhOD16ux/wGKCyF+L8pLd
yzS/pnO+La4po52tvD1Zcs0yTE6s6gIFf6sAkpSb2xCN82MndoitSlg4UyPu
/wBGex17bCTM00KTGhR33YnNomMw0LeCXTYj12KR1CxTxwqKa8Et7tp26oWh
jG5EGLj1pUwOTLiugoyDDSDPw+CACgeuDAb10C2iOfXvQyfmZXPU3VhaYyea
EHS+hGkIKsfQy1F8XLcazZfo7tEDs9qmR+Hx+1UZGnRzhfyZJetHf8p/3voX
QxWISjaLMWXKpQs+751xMZ8M3QXeHqH+WuFzIsiBMSCNorUOW303+8dI2nVN
s2fr9oK3nTmouBfnRkwxCMAcEGP9bSIeE0NUtTSu3ch6UFT79ckMGMXvnRRz
YtDuUsQo2i9GxPAU6msvw1poUdJIudfjMkfzOAw0UDbvu2T0QwG3rIfs59wg
hYmP5ycPzhbiDfwRl8NZXO6uhzXvfCj+G5vSO61HpwxGlgj2qRfzqIYC4fRL
KIW5rnKMBcC0CletuEm9sayR6aiXqHUNgLc4DnJ9zH3oACJ1OfWnMnbdTuUD
iw+75007idIaL8vV4wHb26VE92cp1cB6/PDFE+QBh28ADZ9VXo6PnKTiN6tG
cBiiQZZqIg4WIvCfp1vQr7T0hz1NErqHtT0Nu2RnlSTCapZO/jEjuQOCMAU6
YoCc2cR+NFAzBfOJo+ZPtW/fjzvn9h3Sbt6j0opc0wPMAq3xoFfTrdaHJbRu
YO3bRwkUVJ5P4CgU0rveM5FXqBpOj28gsXka5k7PU4MSKmU3XXNj3IkWDqyD
cRw9Nn1TWVjaDSqlLWMx6mEwNnuojF3ghMAQ2RUpD1G5LCXkVVbEtGMPe7+x
pZGEPZfqn4bxtlYbbJ2Gri0I83RDZPtW3mnNjr9Xs6GyBxn0GnmqqGunJt7M
Sk/5WiA2btvYiIlC/WdjI/EVeVmwMtKiok4Z9mMqIYtKliPmNWmT75HwcWFd
vd3C6DKAq243fndBLi9UL8ed/huFa8k9xTwBWQMo1lt7xT5gwgfj3Dlx/kJ6
NyqFgozuglLqJyKl0+t9D6QSA9mmR2AKHIvjyOkLXsmWaz3vB4Mm9mA1wAH6
bwskIlZCQOXPnpMjF8W/dOZmVfdZnGmLKjK0BlovVA6/4VItV8WXQ4328dwu
rhVLBT3I7BQzxzDGNOy+EbjbFu9IRkoKb/LhIS0nEE1nU/1gYYlTuQYWhiI4
9uRjKFTuDnJd8ZIBztNIScshantCuAOWG7bQxCJ8w9a/uQ2EUofulZ86Zzeg
RRlc5+jO46knbR14/6Lp/pyJWfXOPV6t9BtxhfFU6oykEmTITBoOOQchhdQv
J6qtX8SzO2vZojpL3wtHSJI0Lnx+4TqpFEK5ZRk82sWJAZCvyXScE4kDCKeL
4RgWYru4F4F/vAG6Ko19dHJdNjZN36dglV4zXak2B09J4f/zrmfHtCHsZDy0
XkFGNjHQwrxjOwcsRSQOP/Wd/dJp4TgWIn/knda6/6+jsQln4mQrvy+TFvY6
Y7UVlvELlt3ClZsq6/OCiHrkJSLxme9kRdYxFkB2I6Kl8Jrk8RGXkLqVEn1x
AoApI30A8mvQC2NV09Q0IWJ3mx+i1p7Zekb+cTGLMyrq6fWNg0fn/889SAwZ
yt0jNUt2u+93SGS2eZ56B0LpOnWoORcWiyIRgb6dx7+0ARK+1ESrjd4ZQwZM
xWJsYY8OsONQZqlJr2TTYi/GujuOhvSqQc7lTSs6/0M8HpevbCYIbAvVGdBg
EHFV9MugCHYu9TOzTB19ccAKHXozYl7LV+0RCr5Ynt/fztfSsrLhdGyJespk
C99aMW8r/wFcpOri2ooes12lKXPbf4z4MyIvvsmyL04ZbtvC8cVw7jMz5CXl
8wUI+0is2cinZ59JbQyM+yL52nepCL+iUq8Jsb2AmKMwnsMCGBuXPlQxRgxz
MMWIpgfOgm+Q/9/m1qEb3ve7d1tSo1Z0B4olhMrDToc5JR6KkHgbKsokhIn+
w2Ybhj7twlA34PP2xcJSIlMQ4c7zszvxzIihpr6of2lzR7dI1vg7wUrJzytl
ZlCOixR9iSFXCiiAM58Tj/zQceXR728AWEzCAnFRkg0U93oh8oJQdJFHIrI5
eSKmWtf86aiBCu70PjhTO+dp47GuLTLPLvXkcKrzt+p0dBnqtLqIG2CI4tLf
XaqmIWo6PnTqFTXMWa72PFs2vqm37CAb8/7FU/kbB01+p1BBgrYskxdI4ZOP
0dBDPoP1k/HwsyqrqH8DO4eZeT/BXQMowRmeNZMKuP9gjEUGIU9tyD4Ynez7
8R5yOMyAaSUbYl36viiAJmPC/tzL5Wck90r0yZdfMwtU13Yia0hIK+LSPzcv
DMS7Qkz+dV9DukELBK4Acqydwg1QVeHjRY3U4LFKF/Vb43OzJXjJtxun1Dmx
fNRjA/FLQMsJHQWTslxdns1+8aqn3DOOhUsFY+GgO7Fjxcf0xIKcgrCUwc/k
gKJOhxlHGOwjMHPKK7i4DDV/n7qcnA33Cnph3+5JWSJQpJW1BlFBzu6R8c4F
de0bsuVXbh0s/gyPVogqXnpgM6PDe6rs5QpPb5JbGvG87/7fegKMg2HsSxrP
g4vCivcGuX8HLn74UAoGBDcoPfNnjeXMz+AHOzJdC9/msYZfaKPAmlE8/cSv
An90NEkqi4ht6vf3FCFg8mXCQKlC39DtyoUru3K0MO0g/EQAM0rtlje432eM
Vqxb5uRedlC3X7AfZbUzTqBjFEB4PiS9Kf6lw3GTUK330NvI8SCplzp/icwa
Bj8g9wzg45Qj85Q3GUMbVK3dkDtOvWr+hiJxyEXcmDxI4gjFTOCPs2uhX3Bc
mGLx5l40+LIlVhEy4CGGtA1bPAp4GY7GPu83lwLocmzS9fOrSpEdcNeMLod1
vvW8lioR7hS/wh8BBDTcUN7nIstz/I2owngCOt4EYxv6mYFI9StnaL+oBYQF
In420GbuV4/Ol6ixnJ5A+ChKnUi+BHZ68V5LjS7afJBBiR3sDcsMPcXZvK9w
3GCpRxgXYmBF7keRJN8yuKXWG9+X85/p8g9geC2EsT64VwvNRzY0EQsfX501
EMWdrZsKHZOBARpZHb5UAUHplrlqgwazjZgldF+d0MGjluE0teA8fkZI2lWe
NERfHH1GiCIr0HOSqZ3nD5KHLHy2Nuf1TN76ZsvbvetICROMcZmfNn+cTtBX
vJhp10hStSV8L4MQO3kO8AzYUHJjzykeW4ZmzCz3/AhgwW7SG7IxpofpxdLk
31A5Ct8sa8TVg1WC4lHcjw/q8i8MQBimX2WRX8QGA6F5ljV2htUYUx0OrYcS
+Dhm+hxOKRoIXxNRWXMzQjMCF1L4x9KQWMS1hb5dP3Zz3IH0vgmoZMtDjtMC
RjRGDSXZhIQOnj9038yKxnE3dMTi12BStzJpZgwHAjNXW2UKIxqQdkdqkdo3
rp6hcMkA52g0p7AmqtpEE99+LN9t/s5Aoee6erblbuvzdw8s38OtsF5YYWjl
KMy/fMhnFIr5o0cbvk1XVdE1wKUE4Ad48IYkXYqObW5h97i/pvGB/qS7N7WC
ir4Z9BnJBloe8we3+4L+w5n/Sog8eHuNesDg/uDRHJuytQ8NRRG1pAq+2Lgf
zzDT9VeZ3gshB1TVqzxxubLtUpKs/oN4YgpfDa8TCLIL6zgwPsvvdy4rYDok
GZo2cG/SAI4YD4CLISptAbX4HCMsZ8X1BuJW19cjXqtgD0RL9R6d9P7sY+4R
GLDDazaEUChi6svxMUawnkN4YTv7RwSshv9Y4GzrCXsqkAnSUm365bUgdT2O
w9ZspQXhyacpHhf3gOCaAZFS5U5o6Cyqlg+gbslKK6SOumhozjOktHohX1SN
X8XSjqXAR1xmI6sMXzkSXRepN8krQnVmG04MfIO+Rp4UomIVSg1SuxdOT/Pa
o0fdc+RVYR5YQIeKdQLhVdVRExUFeTEOB0F+ZOTvGbLoDQ61alN3Da0B0zUI
/vX9wZh8vtF29GNZ1vPMbckBx4Odp3cSTSDroGbo2GtG9A9DT6DNMHZ/jdaH
qBFaLsiN7w6mEiU4bokkHkvLlGIefokEoGDwRyKcBB3nZ4oUaPIp1ywZRC9F
pzNZXnHLo+sY0TFTOFe37/RTmjKvKZYWLUf0raaWNhdnqaWzwGuMmpk+dIuf
k1wEb5WBKQy0lVpmykaT134VeLqqtKFVj5E5mwizUNRgvhpn4bx85iVSZDqq
iTkehmtU+Y3HUW6ZbYP73aFmsKIKDOBVLN9+43Eo9reAspmaoj57ism+ByPd
XLNbi8DZ1D0X+fKJx0aEVkykfj2P4UuBOVmrdP8en48lVv8UCPk4zTiVgJVE
ef+0MHwCv63Jnd8EqypuPiPh1G6Eb9AAU3f3VMsgmACT65gXTInewPxQ86ro
VsBz4g3VxxxocWS92zx7MZp5kcr8mR1I2FJIwPHHHpO10HYbF7zHHEhmYkTE
4Xn/CMJuf1TcQ+zLbKTTkvgQ3BvcN22Zc4xKNwyvD0+ayJbpD0rHGnfVlUaR
HbC6wS4grij8JeJABPghcEXiyfq1yLm+mv/tkSJODiUfOMJSPRgACCfl7lKg
hGPHhyoA1USyiLKZ3i/ay5j8oWUVOOjol7+wJ5fh87A82M4CqycAml8Tpk3a
0hafSrpYXx+r2b8BHd39ogKduLsoTCb9aaWh4IsVuSPxuhX1k9KGXbmDISjX
qdC9evxgZVIzuVzJvpDQhLlffuPEd/BDnvabPbmIt6c04b0zRPNkeUsoQZBA
RGB7Eiz8BDl5JLPdtsecoYjuJd5wlnWcxcUsEVJMcKbFlFRaaPqG5cXHH3DI
4SQUdZlnxq/e5mDnUOixLKmhzIB9AR7Kmu1Jp1xVTMLiNUNepvnUr5nhzaRM
n/K+aG3laOdrgI2U1tvDq2VqftISwVKeGXa3KRYEMCe9/jz6DksgkciOpdIL
jccG5dOdNdV+Aw0z4qqiLd5jVZNAjL6//GzBoUC8IailvWwLGY2wkhq95g8t
IhfQnYkaMZ/ETVd1E+T9wo5Rlo3b8Yr7jCYjLYvJykDxEX113vZMoz4Uwt0U
6Wz0zaEndx9tif8fHhOVf/JyS3fNWf8eOdewM0EnCyuqkSlyJQLW+4LOUUn6
pmwvRW+Vy3HS3Z7cS7NAxAWttOgYpKxhosNLKG4oAeN9SWfk+NwpsyVX5X3L
YWm4nrKO7SXUts4hPV4u19mbQfAuy7of2MoH28DOXvR6AqisDelgzN8gTyJb
XA9eJGvpc0W8pfZlpezEmBgWlw8bw7+6tIAMXwyon6V+O2Q5PBeXAasG1643
eP+4+l2kHHulZOP8towr+Du8RnARybQEYICsQmQq7sAr8M3hMyL+ejX6ttYh
QM/YtERhi8d/5JmUYe/VfL/z3MTAMxvvx+DV12cD0K9gGnxCrWx1zaQh7pcB
rjhN3PT2rgt+7rwxTCoKnE728qknFgmjZRYy3ms0FNRC5e7lndBe1rFY9qEv
ZVsmHoXlE+5fSOShM87U3RP4tsGxozCUYdN3k0XiZ+A2G3zsvq9/puGFJdS9
H3P4w/DFEXfBc+YhO72Eh/qPz1OX97ObY9Bfe72S4CHBLkLCfIDMfx0B1bFR
KiJYS9CwWDzh0yWRa6FyPYmv7C0gwiTHzM5GIBGZwlLA5MLNZSHnnZqCMV5A
INmvVa1y8bzb7HdHPbxktPXxaSULYk+Um7eVx+AtblszbrZE5KEi9At7cuW4
N2ttlSG3r8PbtK8Hcg+k+2bNTuNefCwm8L2/sP7D4IAaIbEKrK+39tmDxeyI
BNwON3pHIjFn29zd6H/oyHdk7Lv8tgnYaoRXvoRwH3qCpc79zXfqXDUyhiAO
y9r83XppKlf2UE0WI86m7YufwO5qi6SnIcersWXeyb2Xnd2h5EarXOCgJidI
umGsBtfiAs99gjyKy/FxlG/iSHKzGnlJryq47/U/I+dXRdWbpYOvJ4E8imxL
vYYE9bTfxqIA2eJmTfCpw9p40kREGSDP4omOeC3EaHe++NxOHNXv4tu123hS
mqfTPk7dmYYzyTMJgjxHJBKz8CCn62HXKfcrkhnN/iQBxVJRoUuiSwroMZ6g
qfOrk1lKxsSaGOnW7ymBXTFsMxfK+o9OanSg2Q1gRRjG+0HwujRA7pbAdiDv
pNJhZBfG0cslOh79iInHHzAT45EHSWBErh+aa2fuqD+UYyxW9QrSCoNRw9qS
m5AFFQ14mc/zmXm2/nMjJ5V007+nv8j1rpSq2poU1nS3UZf1a0DGO4TV/mwu
uekext3At9OF/fphQgpWTa43z8sc+TveaRPir9ink09570sGRi/Uo39qzLuS
mXw6XP8JC5PymGTMztJ0FdKCGUnsa92OUyW2wi+ECDNffjg09+C+sE4vPVxH
rA48/yUtAnud3M/Vy2cpXGUxbYYlyx417js18qQ2jIKPASRm4ETfamfdDWvL
MI6bgIbzrB2e78lHVRqqhLEeQuPgxF1OInXsdlGQeHvBUm9qnINp9q7SmpM+
6XUbZJfB3eK/T5xcdEQYnNzaMA+HV7Kok4xSXBBBKTO1oikBmdCFZYuAYNzH
WwCm+DrG8AhXa2JLR82drV5k++s3mp0YNdiuw2gdo0KOgNjucMR1Ll8d+ojp
BeCBsVIHu4+x8YCaBeoDDMjMTNacLXKMpA9xiHDDugm/eeiOYXRKGcC/cXE9
yNjoBBb3B+DcU4cDZGYQEaLCAxYzVzubRKnTsS+iep9VkM6J8nFXBbBWSOLH
xN6c1UlpoWkO8Um8jTuR7bGWsNwH2lmntz/H7/c3UkHwmjQmq2U6Pinx59hf
persDEcGHzBN9Jw69BqHBzh158pkSB3HQZrg6Q+G0vcCVigwtpJfpsAwwxTo
nDaaBa4b6vvlclV1GAih80Om53fyhhEOSOzgBiW0wH1PhVCorAucBbIsj8bB
J/HJDm3D0iVTzPSF0gQ5YWwol/dkwz0ovzR8fHJXnm9t7fbHqMr/IwIyBCGy
fRIrS7FSDd6RX5DZLRFM/cet3yt29uP4TG3ebb1wBdWNUsHRJ17ArjIgaXau
8UkpNMvVwm2gkIbIJgUO/6VJkXzRfeGWn7fopQ1NKMtFAOqWfjdkYh/fEDUd
wRShiIhuNS/NLVsc00cXJMR3/EWd/QMsCfoIx9vAx3ae3OxVcJb7cIqR/eF4
rmbon9cL91OV1ALbFW5Fa2WuSOzX4dtonIGO3w/pbzbf4h266L32nIxtTycM
8HFkYkPzlnWNfbAlzTPlyDn42+7ptY4kDDTBNQKfnc32t5iekz43g4uQcqwP
/AQbrYsusMmYWzG3U3BrOLzDop1YyuT/C4qizjIQyIzcNaQDl6TCylfvBX0V
jCY8V/pytTrFIGoI3HDcWxNY78sdNlafH+LMOUdZVB2r2ZBhDiORWZcegENy
dNFV3tkr5UdBaVqRmNgsjPjez//h47dMDtuMfjAoHpPDOsMJVTdydY/bM85C
IiswkaRA8d86krmiKXYuaEzaqg3jirlxQ7fVARJflw+NCZEDmh2Hep34Ea8v
C+0tzLU/wwWzdgg0VRzr7Pht8tzmrv7kiK6pi9Kqo/TAJ44RAP8c1+TpLIat
oYLEwFTBZA0NZv2aQy4lgOBzDk2+YGyTtqlCwNHhgbXKUKSrhT1ODYXjvp2U
kp6Ns+VMHvIQ2fWhAQA6ZKJOJ10e0VPAdJy2Hg3bSvOvFoROEiQf3Xvo0H+n
br1JAcHQrKuPGcD3hZDL+R1O0sBrB2MrRtLOA4IPUt6gCusqdI9LBM18JJVj
cw88XJdvxBFGr3S7zt/MQv0JyAvGM4f+CYhCJG3kbEBfAXUTcPsj8yFr1qBt
/lYVfV0KnoWdVj7fKKzKapjGoHVlpreEhQdeWURuYbe8RSOD7Au8K0B/IFUL
1Yb4nMZixupvfI/5znFN10dxeThcNdlDGNjT9o2OhkkK+gm7xmB/Am9pUnTX
WBSV6bTgTzfezrVELRBMXtTmvHQCh17DAuKjjbI/dfgBuGn9/LWQb3lkJR0p
eGut2Qx3/+eqChB9XatVD9iPWpmOHrduQ6X9OCn5G2M1xXQ988sjTJ8hQB/S
5l3qnoR05fkTfYHNwP8nfIlARatJPrQT5G88WG1zMr7njxPQTswfwH5sbrxJ
na9NMZxxEOy8dlUV5o66nnrPkrHXZILuk0hKOHcD9itqRzNJ6QHxwzegQmdh
lXb6x97QC2sXEuxwwqMyYLwzcl5qzJfZrjDDjXeJyKwOkT4IMgHZL9ntlHGT
tAKrYkxJ3UWHyP1FBCYYC7dLiIlbfUQEuK31VSkuMxgCkrBhKB17Dgg42RnR
R6RHjpuEgiJOCk/S1zi+7S3uFe6XpQEr5W5sZUq2FGPfk6xzAoTTfmW/IgsR
yAaABLA0pw86TKPuy1ynfC3HH5WCNzEAu+EgrZm1wSBgRTEHcpf8E+YxQYEF
OeEpIuQP4ZmqOlm9X2xu/rBEWo4RHhiY9285HoWq2/39cl3pTJWgYiVh2efK
KQYRVEjDqPcIQ2h2nmaJ9E86hv2YrhQTEG6IZWlWvKMYwMs6ycbDTy4qgjB/
6Qui30q1373N2bU9w+AhJ/kss/eU0kVYSx+/QcZP8k5jzzOKJrYbDEY3aJ/W
Qzyg0kQD4YGq+qJE/sTkz6DT1fYCx8t9S8g5KS5fsKaOphr14Y9i25oHk5kE
0foUkZ+uebngc3kxFPc3/Bwjs3kQNaXEE4m9dXRBijn4vjqme4ZHPO+2y0Uk
ymsgpAcJ/moHKH5q5bgy/cvBxwEFpVNiRFs5CvCihf4Iru93xj8Aj7R8xtsH
jYxiAzzSmbcmuoxLVsO0Tgx79RGKlgIM1RKa7Fxns012nOeeK04ypszMhYzo
/6grx99SscjF67mU+sARbrXNKYoy5P7Ml5gG3lmy0X3tyVml4OpEm91YIf45
foxFTWvgJUPPVj2Nz9gcsTIMgpeI+Ux1eHljY7FxNHiaB1cUWN4tOLspogoH
dh9kXAokB3ruvq7o5yTUtuFvRreqg4BsfcyEqbX/07BOODjAJORVdnZKS9Fc
dbzqbGTf8OkU65rW4faCqILMRfUpHqmcvJkWOlDYTJ4863x0JEm1KEhrPLQK
OOWPXWa2YkgKkpmMuAxoKYZU0mkjUN5PeQAge98KQzZNh+c0b0AFQw1xIxHi
iy7KvluFcAqxfgtI14yrSjkTLDe8w3mmOyybnH/jlA5KZDq/zhSDDfuW/6aX
Aworv9No5rfNaEDrmr5ipao+IwOlp9wLkzoHhrnVbN10Uk5WIS0q40JSAxah
B9tdWqDMgX0BG26kIIDceozd0ral4M7y6fJbksWISx3nHMUVVGltKajGJ/mD
Dc9whHGWolvecO/v+9cn2p62rW7T4/3Jw/0Vv/qUWfh93l/mFkB/4YNs/kQ1
iWqJFJllNWZhTk+BEHmpVfaNacieT8XAPTGqm5AhK3mp+ZHqQtsRrVYSbhmF
G39N6Fks2cCbgvzsCT+OEZay4KuA1xahdF2BcSw2wBAYLYq4RIvZUIxpNmuG
1j2xZoQrpoyaZRt4UsklBaA/yTer3DyX1bSuY4EJMUZ+upKrn9oEtxpsfuda
VjnVraIqUeJs8DqSGAJX2CQdiUB35vI37hae0vSiwLbixbJPu5gh8tuI0U3O
Vcin5wHw+savx7+b/R5aUsrh9oZIQ1dtKOU+bFQia4R702O93pW6jKM17PhL
kam54LmMg8S9UcEzhEbB25BJTU4mTLqbZjZuh2+Ya+Ii/hoCj5AyssG5W8n3
ql+daDS+4XuaQE3K2KrnT3/Oeqmj+zLKBDIE2DW/q2FK5U4J+Y7kRcz+rjPI
aRinDdLF14075/rM1xzD8NPiQuaukcqLjUoi7feIWExF4MU1le2+muxfhQSk
uIMaNTUQSpE3YG/R7ZRrazrse4GIYZMBGzu0WYSwk7Qj9jyx31LkUH/ifQ73
MIhy5sIH5u4s66gc6ZaaYNyzSLZqTqysIYvaFOTd9IN243isUMATHgt6D60L
hFL1D614xzrKJ/3xOyVDa7MuDX5HPd/W9T74oUJ64KUoyeldLd0/FRRNq0GB
VxJM2EYeBWLFNg0qXDG0ccau7ogo9Co8jI2NiR/GXlECL7+OdhdllYQdZEBx
NwlYY05Gb17PxFvnda3eDDodvsvegYu/jb7AuHmrOmYWIWOCP9/zVLpZX3tr
yx2q7QwRWjCHnhr5PE9FNsPWAdFTmIP8PjPFCreunAF6GqhN5DBhTl1cuZqL
yANwfksEHM2gP0FJYZLffV4eb9GouIum+HVhiGq4DVk4ExjGTHHGcNV1MUQF
QxOrkwdW62AsRkiCOzB2ShlFExEfBzARSwqu/QMZ5VVsc8M0BDdbclksviY1
xmibDFL2TzKG1kXy/CrCiJ4VDNC+EgJHv6PaOvMmYn1jHA7dcvPDzBZHLXMB
KbaVHEy3hhQ9u7h3yzmkHzOHymCSHRHNwHMZiKdUvoY22sukcgMvJTUxehmM
Hu/qfK5UldzXGR0x7+JFyThpnBtQWBj5qXBQKDWofk4E59NbijGv21pu4wv2
KH0UKMmS+81zBxlZcClNBxrxYo4kJSxO88Je3O7pYpsooDt4xdv49ELMRq3F
utbd6N9Fq951mJjsbJhq/78i8162NziTKEP42U5ChcRj/nCm2h/CQRos4bg9
Swg7mLwZbtbmFMmm0YkDXin+ZKmmPsyRL3bMACFLu+dfLk52Q/c55vRoAoXO
SRi/T1Gs7xLVohf5ErpK1fW9khkimgucSZ3bow/pqprDLFQQU8nESGOT5u+m
vgDNHTQ5N76L3qHZaw5+NSBxvPFWaPCFJ6dKwcCF65+H814/sQYvhdO/CO8J
UWlkfZh4ucpjVSmV1lXbmsY9bAtlOElNukspmIau+QMOKMfyMlz7u+QBftcP
Pq5m0bSnZG7SHrEIZLSACDHD73Y4e9z4Ohhm2E2Vb/Rj8xZFl1gd3bl4zd6r
S+cB4FFyOFpZmVwxsRx6rM7wgRhIgOpsbZFyI0wR9QUkkk091unsw0/RYAjG
gznwcq8Xpx9XLbJUJvE72JHGo1QHr9twXbkX7PIy4DdZ84Hz9eI+JZBUW3lM
bB8wIDLGbRFcsniZ4BeTwQTKn1MfqQZNYRarK+ReGW1eK/gYKU9UlMv9jB13
lLJhESHOXQenw0KYXR4s3La/jjYrm1i8UYmiGbbY621mzTxqV7yB3En1scMJ
gIfNUfB4T6j0jg7Iplj+OIqXup9WklRIsEISmFEdzPIPDPTVwkMiL4DF/3dk
RTqa/cWanoGL8rB3E1yOfZr7nQW1mq5XiWTORJTgq/cu9U9ZJkmFQIFd9WIq
0FgZHgIi63Zrd0WiD5tQWf+vOnyO8dtwG4MdRBg14UyFk3K3yeayrWdomnls
xAeC1No209csaNuM4ZsTy5b/1QnxqQutRnSnGAqTIYynqsU4r0BLlUintyaS
lNJkuXfTqj8Ly6oKbYhjwoHovmb6Tvxob7AUHUj7w1iBXDGX0CDCcbRN2wEO
cGj5TVK8aolwK2xCdeKJxZ/WSC/884elQ2dVsyDtxGdblGu2MEo+saVEEmGf
gOZwlvQv/MC5HHzpsRfbIYjuUTBdUo65FhUfLt8N0ZqW632zQZHAR9KINXC7
e6kWyJhIJbVe7Ee7Bk0GCJwYyESh5gXapTU0fQDDv2TCdQqlAodwrrljj7LG
xSsricZ4qTt15r/p//MpZMA93gRlwCrjTVjeTskmsE315kBY+iSYW+0NfE+S
1Kyyut7O2NVsmwVmVBTzQjlKT4Da/HIIIiHf+6sGKG+XZXAWeosg6i2KXmXO
J9/+khhNKJcog9eXjyUfmC1oebYVL/iOShQEZTsNH/b8AzAp/Yddaj4G1wwg
f9KOMFMFJiWfRvD1B0TGNlIQqQmxxfNhYYRrlwk2aE0NXkMbEJXexiLS5baG
faGSLsMTz4vRZc0fnlCg5UZAL+vTYW+GiEoOFzk2uuoQpaA8Lq7rymAYJYC6
nGurpPXn1nENhMhowILMu4dl5RkqPP8fRobEnyPIg9jdrF2CRcrYoqMUc01b
xF9t0gnW8pl9dTRGU6Cc2b2jU6uOOr83GIKhvd3K72xQq6qDFCI3pzRn+j1l
EE4DFgB25Ku3/EFmlyf50qtvyyY1o2LuuePU2KJmAVMpGOEmW5EXXZ80T4Y0
SSbfc8gLmCYypFTaQd0W7C3bb1HkRk8X7CVGF0prpw69ulWQ9gKUoPEdPs5h
kXF/CF7KGZzGukfSsjzuhkjItQjYTUgizhG8wDMnHRxAacIfyAynvEt9Jqdd
ZqqTzb6z9MG9VWUYSpckxe93YoSWHZcqHMBvDkw6dJN4pwnFlx/T95y3wKAX
pk/zVkljy+fHwYOpl9dx04xTeQN+ChzoEqAbiIUrNMyu81azS/7+EfFTDczT
q8KkaysxLBeS+Iqcvcq7XrtmGk2AOL5rXosjhsnPvrmOw7ZbJm79igD03XlP
MKgsbXDn0hXMTHBm/j/txCEypMxgldzW0Z+CRtCo3kMc7y5UjReIzpApT2Su
Edr3tImnv5T1Mx2dHLoIaCGk4mJGwWIykk/tXMZ0ffV+TOG/txP92x6kaycq
dpLcf5hS+xtifJmFx5lf/EOcx5BrEewK7G23FwAtIW3LO22nqtvPD2KLBDPC
WjW728istxzzh75fqF65fqvZgEeOtsBp6j+PaXxT7GyVPoCC1n6QsN6z1Gsa
3Wz8/oCqMw7zGo/MvhkwzVPIiqUh0iGTzOQfBg9B8XTa7hZnKzXF6i5G9+Ic
t52wPojwo6O1ljf9m0kRvvmz2I2KSr1iI7VR9vbcvPx2+B/ywsf/wtoinwCH
na3Ggdo7DirMSCEPFRjh/n5W27tdwFbyaTPQSj98dIwGvf638z56t/QAVQOn
gjJR3PvYkVxfTXj6dEa/Xa/EcxHvXc8AACmGpjklFQt7qDD+jB/AqJ3Di3eR
cDtFQQwASE/63L+QEzVjxA6Mfd6at/KZeN0bpRPLHQN0CVOP6+6exdYAZt16
4y3nC0JT/54syiW5vMq6/JL3c178bi3Ge1Xmv8Smaxz4zODw1MqIdwJ86OfZ
NdYeU14yTnbvoJpYq4kMFh9EusbgCNMPLxLkdjfkpTG4ZhHao6MTovcyS2uy
6q//dL3REPcNqTsZea8tk33qbBYukjJAlRACm2EzhBHahQ2dPYPCvbHKSyEj
3WXL4cUthgKYBINrH13eNHCXtEzv8CqQUTFkYDTKr+lIImNoUqPy6iDFoKdH
WxmhVCOLwzpiEMtiErJXI4dVNLukGZKE/eLMYPxfzHQAtiMNJ9R4v4LH3SZl
c+cHVRNJLTkVpVvKzhHwfnM4H8CzUZyUSs1E6G5fBeDT7cDSSUMARseOpRzw
7YArnHEvigNUHdmrCA979xpZz/A6XmO9oSHXmG8EF99+KKwWSsB2zAyRpX7y
A0Nq72vJujJ1fXUzyrfIwOrE8+zRvlf3yzHjNMbo8RS0SLYujpm9I4hQx9Pk
UDqtwcNfOd2sWlaS9VKKDxsZ79ZUu6fJmu7ypQ291Y//BQ3RSyTl0h/QAbwX
6jc5WdPcXB52n+XiwCT/6eBezjHcHf1xl4a1vuLTpxnXTuCIMmzKoDrfG/JJ
nN5MHdaFGFj/gsCAo9unTlabu2CNSra4FcJB0t2rBq6o4ijQPTIv/YyoRN+E
j9lYzkv8bB+N3f5DdygqzIdt9813TVgNrL49aF0gLAH0teG/TSZPIwNQd9+A
nVKnAUlpfw02RGnJMlXAutuTPyWPqXxoqN8PI9OwFeVRRIz5LNF3MLkI3Anl
ia91c4z7n8+7XFxPdb+jacsmJUH/b7qX1NFHHmBBz36d1dRqHKGY6JXykK9n
bZLyZHptxgZmISWzaC1nYIqmJ2I7r7BGVO6DYnkXff8iV8m67RHiZOCveTbV
Wx9zSwoS4uIvRTCuNGJfC3AEklFonueLJEWbER6pcHUIiaFtXrT4bPclfrmL
7Aoh6fqnhRgJ2JJxFz6oKUk6V0O8i3yOKCsYGZiMzxfxvDTp6W9HRxTT52be
s645NDM43c02UylLh/aKkiKkxf0BoSLMqaPaaH5xlKJY0ZJAANjgbwDKczXA
OOBr2n5lZl6sMPlQbfbIlSqjY8zSTWD7+eng2ZgOAmxSSEJeMQnmIpB6KdiE
vTdujVMRM5M4HenW/OQiaBXekThj0rsc5CvHD6QclbZDxq0QebHI+M+uYydJ
KPLCVDQ/Ylk9MPeu1ko5p5EKD8eUfKchU3e6a6VgzDX5lANAHDkLZgiBut0D
DQOF1lkzpcdVq54C7e0N+VY8B4ges/D4XPrvRVKIMt+UNpCmSJSziA64PPdq
btg73n6e6urpwjp9pmqumYhw2/ZITWmIK0VabO2BaGotlDu/VlaAZNXHKtih
LU8CFxQK/L8YJwVST5q6kLtSL6dJKv/ChxWCHtWPRIhtyjhsjG9TDAbebta7
uEozkzaX/UYpHaAuWa/FdxgiWuYCC4Dsj5PT/M+HtjRhHVvOePQPkgcSygm2
LcQQSn+cO1MmbgX7idQMOUXFzB2xxd6Jt13YOA6Tf2bL0qiHRvBvHsL4zEiV
GRC48/IhD2noslj5rQx/NAZVGzr/3dcuaQ1Cv8DYM+KnaHOk+g6wWP0iYFfW
k2+oZb4GAKcNn7kD/qV2XfY04336mSlSn+tubeS+LRcw5hPOrcs6VMgwEB2T
Yyc7j01RhAxpGSXvretUL1/vWuBAA5eoauaRGoMkfD/Wm3XP9pVR/NHp/dRD
AByNR3gbWEeC0ylhDhxiFv/Pa/n0MabjCNZZZCInLrKD4l9lFkj4EVk5l9fW
5bCoVz6I3Fgc0l2QFYv16M1uPDI0x+1c+n0v/5zUzsL7DbAeucwbxIUIWav2
WaOJQK774MWYW2E2TMx78Am+WQLdbxfTjiUpus0SDvvZN6V3SI2aBvyXkM4O
GMpegNtURsqdd+n5FqdtnKzQaPR+4JU0Ka6UbxWUTXhwG0CaG7qga3R58jCQ
UiD1gKwnntn9EKReosckOuQqbLAsE5uwR91zh7hkbbafzBLN+XQLX7B6t6yA
GZ3hCDBLwuEBqQqKxSXCSD3v+oQHs2Wfl5VaSamdfh9X3PUB+vl38obqZjj6
GY3ubEq8bxoug52H2T9j4ODREVokQH5cszH732W1IvhhA+OWrLvWFdr40Y6j
TIZc17lPtQcB0o2Ss+V5R2L/jbEo6yMRdhqPvYdWBSjqYcMBzGPpgbV3Su9v
NlH04YwjK4pBDKUhdX7OXBfyMVOuBMl+ZiMiW0LSll3mm1kKy4g+8RwESq/D
nQMUUI47cuhMCZ48akte8FBMcW81VZzHdaNDUH66F+RL5OE8u51yXHyUO2y2
OnEmkJxztIBNCydkVewkqrc5/6nDk9wrbZurUdep3/gKhOSUmQMlnjPpE8Vd
s8Odkkj6htxdCJGAy2/dkOB7YPwJS7aoBx3up78VSLX5RMuBCN6lxWq8+5fg
akUDjauRwQSm3w9QQhvAqvYKRa3DHCrPin+hheN8+hy7tr+uh9LVKguwF8Al
kDvZk6oQyGLk2aVG7BZBpfFO6Xyok/vCN0yx9g7zX4+DFaKOYE/FgrsOHU6b
YcZFl9UYl3prkA2HF7aaQqqXOuiF1ZQ6rZPxmby+ypl97r0Wj5os8Mgqvu3u
3MgDvqR4P6fHKwKxcqF3fKxTOGUTjslMXV7TxqHG/IH5UmeBr0dzvv1K37NX
k7u0TnCjfWD1z/EZmVrIvCvbaejPgGUE865p+bwUNeeDQXQvdgz91ZAUKz3y
4yyItM2SvFP8FBOD46Ou5UueGU2OlMvXVAzU/v1tQopOalCf85qhtCS4DsXu
qoJ3RDzwYLYEf+72v/exgd8iSJ4bo8aNahzh5MQfq3VXE5N3ZcahIvFNe7df
KXdVIO9uLGm8dIOe3dgxuhJbji1W4i7XzBlWfcZO9sc+K7AzZkyBUGkpj5nj
q62xsq+ZkVcoVlNLNGix8n+SMGuiF+gsbYJJ6EChvTT/qDpIg0z9Gin6Glo5
OPVWfFs8JI5Bz2aroZXOHlHvDBC6hxB+QhU5PJ2ZHZOdRyt5RkaIrM+ct+Tl
G425TW3YLFcxZZU0qr78IB+E9d+GEugfrYTFnEtlsStoKIDi/GD/1QegmSSv
QqyZMs9M/ndsCJ6L7PpBy7X6zpUsVvGeRpYNhJk/TygjLtjsAkRft5JJ5b4N
RvFvzaeP6ApScJMfU6r5j6+mlzZAesSxcrUOKor2BdMpwdAEWsAxOJvizDjR
Y8N8FIpnJmcVtEtzkdaBDlOvX5k6Ry5DCOvINQsP7pPJ4R27ai14GXZE/qVk
oivmYyYb7RpjviL1oBCWUnPNfJ4/zy1MdizWweYxzSDf08hzk4w7Js/oL8W1
CXj1zefxS2c7ouZcu/CDzaQgyATtK7PdEqKkiWbscs56V6KzuwVxxxGiY+1U
4nnXukqBPu1/fPQGEUtR9yWquLrhiDs2s7edRpP675rSjczKVMc9WHEHusDM
dL1mB57+hWTg+dhxEWE7sevdGrg/4Pnl1mCzyqluWR6DxkKrDYUXAxqm0xAk
nYPmzmKGC39dsB8qgiLzKl9J87J/OUa39lnh04Dl5PHAgKrTdKE/ZZyr3D97
xtj0YPUcxtYr2pkBCvoV7mazN38pTrEO7WN9eU6zPXCwX4b7g2TVzpHHtt1Q
PCF34oOPbB91e5ZabRsRVXxviez6I+pGhg6FX8H3O83lclTSN26dfzyebb5P
iRyoT8b7VV4mjpWv4Hj4Vnrx/GbJWnq3DFXNS8VhwvpetXLaYpW7gIsKBlyc
O4MNq+kQ1oxL6s6L5W1QLtucPVFqmjrdh3507Wp7XRgZFkZ9nuAiXylk/ZiI
P4T0qPnB+KW30MXaVYZXUT3w5Eq8XwRK7Fa/cxux6BLgMzqTHhEb/SPUF/rk
7ReDTUQ5aZjSBqdmyvlKgxIleyq0pgTk50wSpt7d4k1+8dyluP+B1nP5Qcya
aHKpIjO614I/bJAya3z7fSAgwezrLuRIdv+AR68Dw4JyIP5FREy7d3rMaRgJ
60RCgZdCbG7tF8Vx2QQiNysQZleWMTKSNujiDWb668USUeXK50Wj4i7Lx+go
xEzTO2kHaciE0+mr1l+I10VZ/yRI2R7jdpFsSkWBb5SWdbeZuJCOUzqgHNii
9Xw1Va/bpqnMAarLC8ikL/bbk0Ue9lvnF8TRKVT6RkPvqlhwndOpUQ5M254a
NaR9bcCRvXkQ8BjnfUFKZ5fsGf2XM3iQk5RHF7aD1921XnuglR8FpHq0MgFL
5RxZ1mWDb/w/jRX+VvXQV3h9hCKwtc5CoJqyiDwVymNnELNM8SXJ4vXtTwga
1LcYABiMlKoCQyCreTe6xRN/X6Hd5QI15c2eNHuUSA01Ft8CCmrFd/+q+NX7
mc+y7PatXouxNAOmkaNj96cwUQjUiVfxmuIrGzXqZ2riV4AJcAWT1lvvVtyb
TgzIcbVA0QLMGi1wLs04Ly6oijvraZ/W5+vnpwBKG9NYNQyyHWgt/HLbKgSV
5VUNiEUM/U+ulg0jiHyQV1gL+UC9qKCNITIlxbx0rL4K7Xt67nYUcEOR/a93
7OR23Bu9OE+MsfOH3Y97iRPwtNtD1UV0hzole7PX4aZCwVzPnBSYGJUxdmXx
pp2qKiENn+9T1hQHJimRjaZmtL2aNT3Q2Bz8oOAo9kwz79DHs2PyLHGE9qj9
5lLva48XNomJQmmA34nawGpgypa7+JABuDF8O9FPI2bldtASHTEMaD49IAKK
97Ex5iLqULcV09Dn61j2zJzTmnu1/aOKbGlB/ZquBQhwEpriwqQAJ2CCuwB/
mXOuMxi8TygKJwfbxckwsFNFMWr8e67qoEtN41H69mcEs6AZOuRsW19Pim0j
LIHsl3BAjOlRoBs+IMkt2/AyU4M1iV2xw7YDuXippbM/68OhTC6DyuAkq1//
R8RjRKROKV9Bb1l0ntx4EjSj9VczEgJd9uqyKE9YQKFHmD2Vk+uV3k2hyPIA
ku//NEKiglXx6UbpArj5UO7VkmXrypwccAm9RZKK4fpoAsQdcFdUY7CVk+hf
wIU/zDIOgW1BlRT4P8k9HEflqt3JfxeZ1bJFWboEkbw9HRLUMIktXMQ64SX8
ji/esXm3duOeTKWs1W3TX3PqJcbY1bmweI0mHhfxssDMV6YKmLbOJFvlh37n
N0bk2o4cy6frHLIiEbVKmE0zhr6X/PM5c4cK27Jg6Mz0N+A7Pvil2aVT72uK
ghsHEaTenUr7hl+ErKZp2X4YI0lRg2NqJVjJCU/CoimXVFPAnrr7XWRes8O5
Nn8S2GQ86LRCWmjzNUdI6OycGOoEx1lYearMflf14q6o+Dm1HjIUTiB5Upq8
jv0C6HDnjmp6GqaJP+qInVWJXjfXEfjPLZqOnEzXWOdXI4qtgYnkacS8RRDA
smNy7xn+J3q3kiCbeNtg4T2uF1A14kdPAEzEpjohkLbiSwMGpVTd+IvptEdL
g0fjfzYvCQ2LV2qn9O5iOviUznYESbtiQt3GNUUs9K2t6AMmbTvlRMns33iq
U2HR/pbiKjm7mhQvLEvohb5ncW/6+R3vkHVOcMQtVf2NuadmZPM6/DMpRpaP
qBrEz/nBGTxlL2x6Af1vzm9fS5Usl7z/06pKoTdM+KoO7bj7zPX7/7HsngFk
+DckwEJv9WI+aZj07z4B205r9skgOilKIF5Tw/C79hW+yblMvqbPaznIXD3N
Ldsio4vAIbLFOxPMvSRgYOKvD3iCWT9NJLbeJJlpEOvgLHiHLEdKIXv5qDBG
rIaBGolwuI+JKIi9ZBHropmvioDxgh1J6ndoJc/nIi3OKHJ14qEOJmmadBv3
2OWCou59R5JPDNLi9L3o3dMxzJ5bIdUjjm1X80tdioxvdNCf2MLNqaoQ7cnf
tskL4K3yUk2Bf0zj7qP3Zk5o3lXR+dY+cylTEt9PzGvpJzMuYNOG4he4aM6F
YDgSLHgtSwpgzP1wMPTycukxN9XnZv9/22DKxgJyT0WL5XTDVPh/7P6PnZVe
wkNEdDZ/UjVkgn4Ypm9z5j2gDW+R0rJ4Kn2jmrfKj1aOueoQkC8YGIe25e86
KBA2PUlpD/hzDKsKg+mdWzqssId2+XK/sKyeSHQtvhoP1zQ33jwLRmd1O1uX
QA/FIUkhcD9/FWoWG6obKuvGqVkEoksC1iMIdLTQMmC0/Qryr+ubP7ZvsFZ+
gyQS5dcvvKofojO+fn3tp6XSGRR948EK0k5E4IlyYwkSnhFOzQsl3m0wwpvU
Ww4rSoy3tgvmqDgQtdnQOIlxLMhI4WWPvLVe6Gf1hJJfvQNgNaxdyZ6bX7kS
nlgHAI9LdL6ud6Ts0pC+ZWl1Wo9+MlYOHUKy3kwowxPS0QuCKdubjI5ivs8U
+Lr2hzPa2OA+4PL8bgjGqYqk4wxxA5ClsE8440OrrLBNYfasPxEt3mZfLWhc
uYwHFLEAAApgC6OnwqKZVd08GKG+RrKcSn2rZyjkQCctDuyCqTOVLKwdcj/h
D/x2hmEoGJtxTvtdSGQ254mr6/24Sd9Qm80weYYJyzXn+zyOLQfz8bjKgnvd
ULIwijzAF1kihpJjeTB6fvwlP1D/rJyGBzs0F3sSF+OauzHf5wOgcp0ov2es
LbhP+4e4oBRqj7djKMXcOYbFVPfkkRtUkKrhr2LP5X0UZDXiOiq5dvcUK/b3
5L5cMV8kYGaHJd4AFiFMVEY+p+qB/1wKV5wZCQP5YF2E9bkl5mp3cybYNkts
eE4aEFkb6fWlKzVIFMzQKLl9qtQIhqzIV724BG5X0//oGzMABU8dD0nWEjRS
A31ESt9HuwTZ4roJXigodcuha/HqD5Q3BOF900TfZdQ7YH24Cm38Tes9Y4Et
DNbXKP6M2MYN/ZAH4X4q0c7SO1MmKppgua8I9xDdgLYjyM/tAMBTh2v5XE/z
8IYgbIDoCITaOx9/BpfqmAE1SS3e1ObH0jTAMQxiwR/lwfLF0lIsHg6bZGAK
iQ7EqbSo9NUE1o9KkKmDMYg1DQEVgOKYIM2d/fXZczgdM/XCQW6I2noCg1eG
Dvw/v3MaDu3eXb6crS7FOI+u2/kronOr3B3Zn99HEB9P7qYr02rvQPwfyTGF
yG+GJ1rvJ4/DLfvGRSWWeT68v6n7hQRfR0vviJPXKif0pazYU3qezMPeODhg
sE0F86vSBVyCVJXwkSnJM2eAOXo/sXTbfTwKLdwBEtpA+VbXkNhMFtG6QuRD
T00Uw07GzkEnG25ubstxoySYl6Jku5CQv4MlSDckiMmJxh96kwDMvWmddQ5T
l18PpdbG/oIcbE6jcj6yHgCuvoN9srLmRwQfBTicn/HmAssAYOuPDW9q1IHG
tLIzCtZP7P9jneR15hD0OkUCEhl3D144iVJ7/2gW1wY9g8MkfsUAwIWgIXFc
dlcpOAJcbyoAejkAlzFmqlt4Oe0ELT69cilaZObu4IcnMpVrtm+ruAsYE0ea
5gZH1Hi9j1YQTGKqeNRlaW+tqtFdQbsyr+Ax3CotamVkN2Tl94AhTd/1HQhg
0Sw4yndcOervIpvz4+rYXUhNds3IF6bykGyZZaOS/EHvypKgCkjhYuyTnHos
ePJZ3vMfL2BrRbwuvA28gQ8c8olv/e7fyQa9ho8hQauQG74dRM8Ff606X6yH
pHASO9B37TREAQo2DTEmKTEd2LA5bFgou2UAMZoY6yXTbSwyoirUsnqANbNV
yO7kOyT3jKexDiFODQWu/47e2N7DKDiAwhKcjDL9Qgq4+JQKWsP3vHCAGl2v
BhrnZwOx7QDA7N29cjco5JjNoI19c+YyjXypUqxXNljpgeHyrxQJv0G9nCJL
lhVDYeGxOKSFFUvVLtpb0L8jphoO8k0wc03o9vmjpo+6RpDHzw3hOEcyqXqX
cihAwJa1Bp3LRxDvnNeS15tFOd5Ftlp/gpaWSOTdoIXr9b5FKBHTE8mEE1dv
hKqoyawoufk5Qo0/mMN1TkruNMl7m1uk1xQLHxsxDrqoxp02EUgam7qDG3Zc
nn43wHhCT5w0Bc+G0+BRHL8gU7HKPRi772pUYdY62tMQK9/F6YMdRYjwdta6
uPRygqtzz2g7FbZNOqs5LZZMSzF4W/8qDYaK98UAD4m8MjiAxiI5izPQYKcb
E4S5t13bWljL4/dtpVIb+wC/iFrA7Jp9fnc7ZgW71RzmhrpPbM625jFTvKtP
2vBkO4CoWqlpVJxA4t+P1JfxiP5lQm6K9iR4ewRm9qTEZbsK9BIxg10cNpUc
JRSZttiEiKrfsyaCVcX+K44CrxBrzXJz/CHlEyGh4tnoMWOGqrRo6Lb+NXp1
T41ezyTuudz/VeRJxcquXR/WQ8bQP0xEh/w1t8cPg1nGT4/UOE+X0jM5mGFr
4o/XtSWnyoRRR7j6EhSprvqy1ym+3n5LJDuP3mCgdnSDcnDvEPb9wvFkbx2A
q2EOr9IW1FVK2nxuhfYyvipnbUYBagMP1K08xNAifCyXLO2wA7QEL62d+wP3
Ew/vVrNKy2U50MyLFrVfUVnZ9pBxqfErXV3S6dh3IRfTPc+s5evM1hwd1y8T
3ifzbvT8t4uPbrSLCqNkJMvZxF3NI68AzkpAH0+OZcCRYxPQTthmaUrmfAiL
t5j0Q8KZeOliMmoMpCl2HIWUsQwRbV4Zr8QxC5+vtAb9GHBjB0LoYRcRen6w
Tzz2iboA3VPWcVkGZh3PdzawJVWJdZtXtMI6V16eGRFZQePT2IdeCmkVW3nD
LO5WvyWIZ50EkH36XW9IlsmfVbiktJAuQv5GFEzZnTJmBGqgtgQS96Y0s3kk
qDdbu5qnZYNi+Hkw/uuqL3a4A1IkQiqCX1rEg4R6SXFZ5a+tpE9cfyfy8D/Z
+XtDHtroyZJMlKrEW0GJ1GmW3XfTFj03zLxX6uloc5ixanmA9+D7Ua+/4c4I
Zmnjl+vcj++RR3wC0wZcP8CPM/WCXXz79tSnjZskMymJLi2NXXkH5PraePOE
FJHiL0lqBo5930Q8xF5dM0wJCXN5+PCgUzolk8pnW8R2fg843kQZwNZ/N0tY
BP+ZyoA1Du0/wvVcxNTxAeisOd1Ob+uWi+i/aZQicXZ3GXvBWrL59zHd6Qm1
tXkrQqEBd9fNExkx2tnDxhWnwUH3X3aMer1KfsLnUsyag3DUe3L5xD+FKhYS
M0t/WHaN7vyy4DR14cOstS0tDTxqW8VTfHp+2j4UD+XThjf4AyZSexX9VNCC
Pd0ldG2J+WUA1W0zkpvNl8XE52kCrrGXaiylqXawL14tOi2eT+ytqELwrA/d
Xt1NfWjUURiYkPLGaPKXlXGr9m9dGf4HWg4BYZ5O+wbISw3TFcnzvNqoyDii
6FYQGHIkDDMFigcSO9q0Crb5lcVeVDGPHWCf5iAqoxIFbj/hKCqHO1y/jrQu
hK391BCzysQvXo/pfwThhZTnNkwmh3bBXuGKwL6UV4T5LNzwa8h1UKyaSFC/
l6luxZaBLoigc1SIz9k85lWGKibCAdtAAidffD8dPkJyASmv2yfmJa3IukuL
Yg1Vp+8nuOGaKxLc17yXWgOLZqX/vWFfcMOmWcCCCDrmre2BWPx4dcgablAD
KGksmGt6he0Icmm7cLeggBWY6ofC/gT/CPq0DB6JlYoSuaYmdWdFrpT1wHzs
Lia19a2JAd5Pi5b2aLgCuD71gmdTwQ8NO4LGpP+1FpakHCJKUS/knQk3ts+X
J025KAohfjhPQLP780v7/nh17i3K2mSblRmGewzEecITPBWXrvFCQ85hzk5Q
SuYseEyDafBn9zyF1Ij+lHfwU2/4TecuOwn6ssEl4bBWmYfyDJyqUwyPARJN
eZhFjboH943F20uiVpEqp8NHUQbxAwhe/dq6/1xoFVPvNi+sR33JpmV9Bmsq
Vsu2KVesAHJgyJ1I+Rm6k1xF4+Ezvgll25iXlPxHCQ7NQHIqhRmryHiObAQ0
2+8DGnyVJ5a3ZEPkzRBbF9LgAIoYAFsn+WbuCVV+rGn8bNGnjXCR3M1hu3MS
L3WddIbHHzWlNR5IrgcaZgOvLgIKCm/wgjDPbGisOR5QodEA4YWYrt1kNWz3
EI0VL0PTWDMkorsOmG3rarSPg+Se7w4DCyrg1YqGjS7txZrrvvFqdSuxYbXk
HiDYzH86h2gDpHCytoFLtV0KxbzAxBRtSPLde5uSUuF6V5/m/9n2EWLmjduq
IVslL/AoykU9yG/WO0O7eW1fIkVvzQ/JXnbeEY+iPlaNzBuIWZzBgbbv2NSe
oBS1zptUiXCvgJqX1d+L0f9ifkBmq5zkK7hgX6gXe7lp/aU2xLqVpUYIFpC3
JEbQDSN/I1Kc118kP5MV+VhKKPU6ASQLWpCO/bRvR47DCk4JIwn8Cik+HzkE
4aNPWM5o7IRkkiAlnjOHK2p9p3d/RhUyhCUytW8Eti57oqEWn2/OgsqTWDh6
6B4nOuyYJOEODABJl6sa24L1Ig2/tuhAzk7yPwkQ3foGfC2Y0xjv0+o4O3lR
QD52zgiN+/YqT5iuwoTRf3O8NSO9MMq1TDvDTxAAe4GtsT1LMERbdG4rbXse
2Xftv+uediY/N/HFKYJ9A7XWOdtobZlBJd77gSNdsDxQk3z8mxMJjkXCZE+m
uSl2GNPFfh8YX/pATkXiY0uTpzqQMY2NTY0/BvbxpHtiSn/+j+yRI+frLbzR
ZHlfuXFhmqbW7Xv8GeAWiDqncoPcV9oOoqoIR93eqmrIzr3N54o351T5FD34
b1Y6elkUW3SY5odx87sDzfkSMh16zD4H5+fkBTxSIYVNU3falcO8B471l64F
3N4T94t/TsVH/1ZukJxSR/cjgxwlJdNUZujsBFjbxhJ396pE7Dl1VIK7SYUC
4/C39hPdDhTTfK3GL5c+whiCl1cEADaOKSnYlLCPgplFCMOhUfE7e9t+GB6d
Tjbql/b/09X8avTtt7U04GxJCVm7v0AqXOZNKvwMXgIWiBBlhppUZ0uDSdwS
CGK1/wfW0IjzfIbNea8/UWTC+tAlEnnCc5VwxkCoORP6RDrTRY+dx/PdUWuw
LOffKLXV56zP3RVN7e3d4c+djk6f5P5d8PTKrfFLNwEeNEtfj6kfet3ZwkPr
rtyaw84czyw+/YczedF5v+PVRSqtpExprp3JkDr6NOkWrgLPM3OecCK/pPcD
vuoccrjn9hPG3RUZTWhZQVYmR17TF+raGSiDWyK4v2+NRSBi2SH+I3MtPszZ
tshSnnWytzG5/XIXA2XkMH2Tawvul7rAV5Wzd7o97yeGHuNCfv2Su5qJYcY7
/rVWtKIDWfXXIKr9EADjZrDHgXrc92g9OGqiEHB0+x1ngiqlGB1EM7ZrWHLd
bWJwh0ahNSf4BsKt1hHxfnXftXPEgaHimjyOCLKtQpPLd2Fd2EaUvs++7IcW
Ovxicz4xYMzfWgQJewI3NrZQfn15eSgZqSSet4BFmxOg0TQn+hV64uhpZ5eW
wHwbi+GJpPZgQltPeTmodeSW1AKszTxVz9lQHE1KLpV3egIqltq1KLMDDyDf
TFe5JwHbLpqDkTJe9q8vizjI4d3n+4oslFIUjZUqhqC48lJpOv48lkbaxrQZ
kBjGqyR3tjjYW5LMymCGumOlGrQ8zjtkZjdoFlwvV+fjeyU/ZRUpqZqn2Zt3
pjTzi5gvg1WOsefhLovZaPq/BGKLTO9zDeB+Lbed6FJN3f2Uc3sKMGlpwJRk
HHOMPYVcusYBuDHvQaovxfADSCz//dR7MGYKE2gUfZiKEfworh/QBvurR+st
aoc8rJUSYSN7AsiTfQ8o7vIXLdaglDGMxoXS2ktJqGGhbFjm5Q9wsXECTDBh
D9F4WyPkBThfYnWJwfwQUhUy66pBMqYmg8J72pN0AdTwF6zHzCjVvsPA5Uqk
7ZQU3uzENfqBVQnZh1zskKFHI/oieUudFR4tk3oOtz2uKwPdsztx6sE3kHu6
L+hYiLplrE0wHmouWfHzPUhw2nfGOxOglcxw051E3+HYqIYxfdaDTim17hn7
+b4sCTyX1+O0WHaJ0tKuVc5pxjcf+x4ky5m//6coS1ZGNHrT8P6dgJGZCbyt
0UsjmxWuMD2GgQkCx0Vpm4c89euKqOcAdMNE8OprLhsKTCEOObzuPQg6TXBA
LSyEfBsMLUlBvK0HX87AEMddYBHx/WOPc1iDnPvOwmpu3eR0DbSX0ztB1gzI
kfx/5gUBxdZ8rAZ1jfr2xF3/74iicqGZkXdNG+Z4qO8+KBc+culwIzsH8U2j
UQWpiUL+VGLY8pfNpThbJRvaQkHPD6nHhb3y1tU6Yr6JFIauhxooGYhnmo76
rmzaMRj2jfAtG2oXrgJCgGb+bmcLpBRaJrdEKgOs/gsJhDt+attdLmIWf1Wi
9noUKHqLo0h1J/YQ/kT+/1ah4QEUmxUkWEeOITx8WbuHiFbGMmzAs0APt0oA
Zm8LTTvhpUtN2g1U9x+wZXtOhut6y2Ux+yIXd/JB3lNwk1perGqGvwstc5W0
uPcakULZSgHIhRbX3KC/S2Z1HliXjh9MrXYP/leJbFR0nmcAMhT8/VmuUk49
C7WXEb8jbUpI9leQJj75HA9uKemo1ZIZYmR2owSxyGVSqx2bywDyA4sCAwEC
/RrRAvgNgqr/pDD9HQxAu2hmV/RzUC2xhl5vJ3yBDZnemuHbjydWUOl5zjc8
5b4+907gfuMyEaYdZ6MTgtAMlMKbvIxZSvf9+yPTahD6DRDrfCX9kcx/wEI3
oLIXjB0SJGVzGyQUp2x2BTDEfo87LI1H7BRKveF7H7ayFZ3RsrCMk+YkRfkv
8mL3hUOvGeNCqyQMPFe6fop1fGtdhaV8eczeU/wb7RHTIQqjp67j86SwkqPW
MIpN8E+iYE1XgVbUFgqjHfKn4LrKU7MFzVB/EyHIb/eQw+/MAPXjNMtHBYGl
uzZAySd9CXhVBcO6yLTBbsd7saDLSB/JvLgwPBog1dKG8XvT3fZDvmFZY8Sn
0Yg31VlvPZCUjotpIZ7rxVetRJsXq5AZGBWmxLyZCzAMV8j7sZitUQW0/bN4
3/+BNj/iV7cZQC+jdg8gXTdpGEdVQHDzdO6cA7VEJ35uemYuiU9i0jMMcUtB
9sDJE8/KkHckRxIzgw7YOmUTKvu62BtzaMXJeZYwhmJEXfbVgLw0w5iIEZ5p
97Vkg1XlVR/9+7S0nIg5+sjdml2Dr/4VnoWxY3G64Q6w7xWBxNCLt0f1YND1
0CeCX/g6vUJeoTHcOkdG6IBlI+6ew00GEZBqOUe7MDaK45V7gTX0RrkKL0Ie
qmnhQou84KfNc/KmjAikDHmo7ezw+qZOWlIX1jZ3zBHP2WaUr9BAXBMzJp6f
jks4C0uneJsmOMEfMf25AR1t1gNfHCxmQEr84VZgHykvxuoeAuDoueV6jmHS
Aoc67cfOd+xHsNEJlBXq0RYD0P3bJY6A984t0YWenVSTKJWu8iT25SR5+Vvu
4PV8PMbDvFONVcFX5PR0gU+u1fiep4Joj8Q0q/vgmam2/4fCq0G3LzGG/6RX
xvjczE1ZHj4VSnpFXuGZgolERasl4GFAC9yxgfBuOmH5sV8Ct2u8o0U2uvJM
Hsld0wNVA3KKDSbAlLnoFXjO4DDIXDx6qxESxoNFBBNrM7IACkHNe5pFhlek
6V1l9eRKeu6IHmsOlqnEaiPZTM0A2c23VkqGddlhwfGmk0tReaX+J/1FWxtF
feVu2CQa0tLoL38RobUl75cH7mtF2c6MsqPWoRbWKwOAGgluIBTr0Lx9mURI
DGCdIweTeNLISv+ur9xG5/WT0DiB8rxSoGpkw6OBxW5etL5bOu27Tzi+dBqP
ZsEzjmW0icGIQ5zjSGvgTTP+q/Lofc+lEeLjUeEs251YlrVw+Xr7r9pjXLJ8
KAhl1HxughCZxhU2GeZP6igNbjBhEFlCq6SN3sadU111Q+Z32uuV95gq5vG9
5Za3H8OuiAUrrXrBtxGVMxY1/DCB3YryXIXSLEvfcL4Jz9cVelQqdjO8ivMj
CsxQoUU4FItJ9j7v8SfOfMfpeiFExXKO7+X1SdsOqPG7+vLFucwNCmeqOG72
7vsLJed2Z+i5+q41yyRKcRcDBkL+8akLy6dOe6oajBpDyEVe2ymoqAioE1aO
s9cOKQKlOSIBRUvl8LaBFIVnP/TEmqAWw3pC2cOhXSUmhDFJ8p0psuIORaaG
KKmfLj0X6emLd4xVr9u8iJwGp2tffGSn56RAR9t7Qs36cmIZoTCER9p8lg4f
YXwn2DK94V9bAD/NhA+tMlfAKN4GU5diXvm1AgO+LKPSD06yu4pRXglEQ9Mh
scBWdBXiF7GQs99W32XKKcsAK2whSyJlo47N05msBikNXigDlWN42yJKAcNr
CwHrL6qYOOI0M3ePN3i1edgiFJ2f9z97oYWM1zlEIru7mlmuHWitOHT+f9Nj
x7v/rIGY89Kry7GRPTc/48XnCHmREB3z1mNcICYbfPyEUzaJcx/O8JWVTVHy
T5mI39jdh/B9eD0EEmB8lgrEFm66DZqfsXi36KNtjtU7M7s6RaBc1uTQX3Qj
DrQNJ4s9kpAFfEMUi7/dFAZQgUfxhWzu9QPWQCPp8NCOBtSe9H4SyE0uzea6
TkQSblB411eI1pRxgWlRixSckLnfbSy3cPcSWT96T2psD5awuspmdGs95idA
yh3ylaEAtR/HmSEe0W+wvV0dg0op2EPwS9ivqQDQ7yKeVuOHfzpJz/Nzkpqt
OcM1SnCJB9YcTc/WhgZRIjtqRsmdGYoEsTn1CH6WhRyXYQKrd2mSFb01KfVY
PqNhdBdrta5e8WFiFyYZeiASntl1pra3OJNCmP70uLEbURKGLBedV1/IfX7T
n9WYQ7nfifyzhqGEmrmcuIoGoQwISJVTUsVyjtDt3OlYoPWRwBfmMcOl/Uun
V9cRFUsu/3SaP1UQYe3nIpurznQPKXQRUxMAMPhr0kLEXbiGMHmttSgWuPop
UXDHS6kEfj3A5scGm0ajO0Zi1uS4dBf6iMV3tgq2JrMZoi1bOnWYOj421b7W
4SYAf4QueOZHv9+Kf4h1etEGtiOW8gC5LBNvoQRWbpjYstzBKYxEqZ8n3hCg
GE+/wyoWyrhhOoulcTl/SM+Smmddp/YSdjl4DBIceIGQgmmokBSQB2ft587U
TrjH3p4LxCen8sZIeMlh5a2TOl1ta8FZ7kBL2vkGVpE1Qp05Dd26X0VTRXI1
whWgPQqvdjWd/BRieqsVfEhjGWYu5o3PBT145CO4ZApdDkQl5btRUbVghNLJ
XhQVZnzQA8xtFUTqYEQcfAmK22M7DAl00qyLEOQgiw8nyD0y5uqYnfVq9xxP
2e3svKoXGLxL8lSGPtVtuL6btsDCGDwC1MMttAZg5LtokKcb6g9c6wf5V3Ve
2vmy2mKqxQI4YU8idUhiQoao/BEGi6iD4bO1XrkB/k8aQCHzB+BvLeeL+SHk
dxZCkl89Q3GcAkZq/DlxNVCIQIXIg7Bk0EmaItPe1kQcnTFsHYSlXm/ZrOZt
1BzAP4PGbD6bOu3gN2WJPZro0xr/vgzYbXxdfHQy13y1mNgCOH1lb9lgVyHn
wLi+gVmDU920eBBUr2IQ3xwLjh7/VXitctfuTfTfgcfYhk/Sud9YOAb0cgt8
Ak4W6gLHk8AqYYrB2x72aU1uZJWspryboXx2/vdmRWzzB6Ujtx20yni0h4ql
0k+jQSZUroBivBMwLV4vl+TbvkpSXrTohqZq4U6JSZCLQ/FTiA/OR+EcAZ5n
Kj3Khzxa/x6zCkdjW+gOCyr6DFm1OhF/lcfv1/GyyKnieMCpx1h6NPFZzmIO
w3gg8TPfOomQcmX3Y6H2hPM+0aE5I2Qx8l+oogEqTFCw1mLxRkAXYhLwK6rV
xfr8MuvRQhrI3LwJrudJ4HGjvKfBFWE7QidPLJoyVjbtEKufgRnYCt8QoNd2
aKOFGxXfxRXKdnLpv8ggEaFRoWTVcT713g1Pbw6z9khekE+XubhBALpK4i1+
mvxsyg7xFGuqs9XagcN+yr9/+c0D/512d73qSels6OpXB1ehQOehkuh4606K
h+ri3MtvWPxrt0xCmy9yTSEaTBt9TSV/utu0kq/gRX88LOD0iygAbT58Oicx
HoEGL+jS/siTfWxAnbqg0iG3Rnpq+rhREp6SwkVlTaBXyP1MfYAQqAWenPnX
sBv3AibXkKewvrymmoKeSs++q/gdyKHftV/mk/fStVGnYaqSVqhXzucqW/aW
MfipOIuB1WMeFdWSNQg+YvUpvDHIzGQ0OeZBQPPV4+9ZuPhAGf5O1DUt/Fr8
urifRNVYBmsHSjusmxk4uyWw2apJUrZym6CHT4PLbTDDk5oCDS1/KPYDqoU9
ysPlUXKSFnbiRcBcCe49ysMLixokM1f9Dd1Oph/QInL6BsO7uCGr+kj/faNI
X/8kcuFCPL6zGY4qA6WcUurRI0EGUHOdYPPr76htC0jw1BKmWodi1/571Lwm
03fnSyekeiV/FcohwkU0MkD+Vb9k9wNxXHmARnoEJvLKir4lPe5p4Bdym67/
da8VKtxIas+Srup8vNXyZYrMAUV2chXXCCuHWy5JXL9CFGnSZLsI5Xge5FFe
2QAWYG+WVS0nV8ysoCSAm2uFKxsmNRlb0scaaA29zMjUHHqLW79nubpE/hcQ
Own90I7Tyx7AHFsxHHtbZMqkBB3er1FbpeMoN5lQiyjAuFbPw+/WcDltGw7e
suZ/3EWNQpFMbYTtTG3lrPMwctF/GrMKarFIyJT6X+C4LB2go2OC3tGz45L3
y7M4lJ3OpKygWUHwM7mG3F0MMX/O+Ghrxn/4iMB2ujYtJFY677pB88cng9iK
Rt9Ho2f32JaX51tHVh0veJGCqO2Tp7ii1dm2atgua3gsyjUl6A/A/gDm5dSW
XxdILgyKRm3WDml2+QyJ9cerUVIgu2JAlymfxQEXsBdm1SaENe5hLiNg3sb1
ngVDW2D0lZS+jsC1+il/H/nuh6UJdJ5u8zg18v8A/2SG4Bz18kzEvlTenfL5
Hb8Dyw3/1LpI7MhNOK7eEbj+Pl2z5fIs0v+VUvchrI+atpbicghjwnqzlz59
4MMsBziC5hlmiXaBbr3MEnDYdmb6AsasBEpcQBae8nKKmDMQAwi54ci3EzT4
ZXqhNlHx+esKnjAomI9ImXwN/rvjxzyDXrczezxco5Tz3sEuO6/lPE88BSQV
S9V9Sev75U8L+TIndVBOeqUe5Q3Plc4G8/4VBbt+hdoyGHLQZTpfYzfAdtUu
uqAP4gvbRf92J4uZGwdfC9d7xivblNEi/A2W2/BFPSUwSdKFzpSmytkQfoqC
ulF1o4hLFVniSyAimH3BlKBALB2gac0Li4YEUzjS4MalBnwZ40njQUZohuJB
Q2/AmHkXmvEVdqZaRF5YXMHciPh1K5RVD7vosemxT4Vr/qB3jT8u5hNMqrNK
OwhEYQLCuP/1/N60DAcrN7NaGK4v6T5Pk92oPlG2DZ55WFSw6MBmjTol7Dhn
vN+/URPJN83LT4izAO1EZ5FApMCsjRk8Wti+MRbyp7mD92TX6U+2SoIGNF1f
xVqAD15LFfswRoi1E9W9bey+NGZSsUHUIzugoN8/m4aCIeJJg1OZb8tNEYw5
IpY8P7pBWh4uHKKc78FyvDvVBBNGxpQu+90Qhpe85tjrIpcyvbuQ7EDLi24K
PTSFQt96EuPLOSa3cztVIOhgMsiK60sc6k/CzfW4qQuyU2Ix2NeDXAVM7fFR
A6pfLkwdvfEantXyl1YkOXtnY574Uqu0nv/e5yFinwSJTsrde7LQFvWVmGcZ
U1qxfqjDUBQhYs9qIHCWNHjgxNIjL7Ml5imhs8H0Tln0tFn5JVIenxJtM/A8
u2aH2K3mLqhOX2IY4wDzb01AJkOfzeoqAemTK8vMqONPFdwKuD0LYPKiOVCb
Uq2SpEsltyycAFl3Y8dxAeCb8qHgpYzOgk4nW7vMY7AYHC21f+wNlNiWcpBv
H6buGk50DKtWtJxxUqAC3vgZDMuDlzR8Dow8RUBHQnFyKh/kICYHDwW6ao+A
4agb7Ojt1AHAVRiktkMip2ATmNh+J22hn0sPq3dcERU6P5zNQwSN0Fag6o/F
uIXNtywl4B8WTeL5Io84EEur7AWcNWnZtCg//kI3tMJYhBsnZTBXx8mvcJfe
6U5IOJLwJ+D92aoijOkbmmRDrtuPND4w8mFK8jQGlmw48mkVwf55OrzbTFC3
HGtFTZN6BYtHAL0cwCXNf+wzdO/aGIs0Uw3EHV5EVYlVoqk+2NUp5iugrXDv
6ESp1eT9pR/3XZOT4tWUoc8kKLQFtdnWAjirgbDPowzWJlK+CFZLiHxo/63j
T79a6wgb2TOBUpdcJRvHv6Nq3yz8Yg5BO6k+/Riq3c73kX1PFJkW4wsciRZT
0i2IJlfwdaJn3tGOYQLOkNKYvIQXnlXMUkqfUmIyyZt3rVKGyLUfpiWD13zZ
3bCpZ94fdFYhUWp6dTEW+vTEywlq/8zUiimTgXw34KdcmtTgw9trVC8upwCZ
st2opfuCZ51FCAaVqHJY8rzzq7XnHIIEZ9Ck5soNYSIJwCtg87bFhQf0L1/l
+PjEHd5SFduwu9vRDVfKswWinWSh4Cnq2jEPyf2sQ23SFsrj6WdwARHuvC0E
kVCOxDCuIHVtQsdk2qJ+o5WL0u7effZNiCThHk94sMK928ZE6NV4T6ErgUSU
M5TmJdTtUCFOlzpviOkQiOiGbgpUA5hHzPHpvk2wRRJaopABJQtUKf5wgAA3
x+krQbl1ylz6C1mi7n2nQaDt6voUJvYXirTzxEaxOEYws5U64dCROdjn8QOR
yKSSrATVZ55aQXwArdeSz4gHNdKTX23Xvqr0prYGxP0MMVUqId9f99I0p3JD
YrA55IkWLucqJttiKDy8hdcXbwz+TolX6KtSxTjuyueaBP6mX7UeDp9kLldw
IKTqCLrVO4O2UYsLQG+kKKQmL7Eg4OW0DJ4Z0A4SksYoruf+L2W0jXIpfPjB
bkOBui5HPadFx1jEqSZxGPRB9sAmTx/8sctrigJnnFI6G3aqdcbtlPhEVs2i
KDftUlB/JgvxtNC15VEcM8NbDefQW9lrMWd0PButTzs4r/h5K79kuFp59ESs
Rgy7TrPWauuBphmw7jurmxEkQBYG/v3zS3UrSDO2n6bi2nj7e6SgxdhVBeOY
uTjrT1r/m78M1PsEwNWDTemuxO4c7EhuQ6SyZn+rT8C6IK4NlxhXm389Sj9g
GwDjXT8tCZV9V4ItntFPUpcDttESLu86jJ8NiDmyepK1nQFCM3b7j6p9nL6C
u0paY0osThYw6LVgiPEMBTeoe63gvoCxxPGPtR216eUpmrPEPrVNcqLz2V/W
QBFUN2urJ1uhWdnB43DjvYqL70/mr++AdcLh9gTfltidmD4M89QYCNtJDskA
87PKvm0UAfbCFQgIyoS4yo4vLNJUFF9V7uH9DML92USZagGM/Z6ZYkUKs5V8
5oPXEOFSR1hry5VoNAgF3AoFnqO91tG6G95Iit7R+02eIZZ2x8HJS7YDDswb
F28iMUOSCMDA2JXz37v5yPFE9icyjMSQQMFRlazearJYP82Ei18SigjzcW63
zDbFZ6df7VgZuR3SF5tC8Mr8djfS8DWxQ9kMU/2OWZkp22dkn5vRbqaPBFEn
HEmsINPEPsDBIyKRwCCybqw0KNQaAQBAZB/JYAmmDuVa1qTXJ1CuyLtmMnJv
bkrZCkFwXOB5gPfLaM4RjMWTNhZoUKT75ISSKYf0GPZ5Z1MOnhxDz/KZFCDH
0510YpZ4sPfcaXSqWGH81QjwkfnwLaK8gKaaY/Gl50DAo3FJgwSfRMkpJ5PG
al9XlAI3IME2XdM1ZznnHJHWve8Iq9SbqZdF2IK/wo0M2P1j+RbxCeEqBFAY
OwAVC9l3MV+CSLp5KZS3zMZ97Hsm6zHVaI9JlkUxdOEEk3SZhVX2Jz+DU5vA
foZbicK8VS0H2y/yzDkGDwoDGUSWim9iO8tzi4poTlZ8I5ImBCu6pu1Z4YS5
uICJXDEX0zuZ6drnVVfiNSfcnRLyXyLs2jUY1+6jV3HvGt0K4zWx4VGGo708
jY9SCnfRVgGgceE91olvX/vK7PFuayIvUt8jL97/1rSpcC/MDNpae4QLkCMD
nEX59eLbWPoOrQ9HCouz45o9MptTbxTe6UOKgWG+cttjP6RdS2aOumEy1CLb
ZfBuyIfqaNh2iidU1hpaUKwE/iXlhyeRx7xS424/sXhwGs/o3MpHN4VeBmCq
0j0SAF55MFKPfwLCqs2UxsFmHRgorBNopOTzzqv7rvilQhjMfoN2dK2bZiVv
pamV8qkuwyWMn8LzsRWnlh6ss4qB/jFUmEiAiVvQGVwcdip7c2fJq1nHAEY8
fqAyl5LZ5Mi9DtHvr+tKBVg6VPjND8xm6/mRsPS6wQFygUYHALaBTt9jspyz
6DrZkS3VAZM4SPq+hhHoyJi2NofpEG3GwKnBaVh+4GmigBXabXF6IdyoNrjd
SyYR65z0/OyDsx31fRFvfK7sJ6FWcxv9gfLsQlvuhSawCZzNiHli+SxLKiJ+
tVWDKiLzn+TM6tYTcXy0OKVu27wloEDIEGXxouc6La5/z32dSn0tLhxO0Se+
pYZpuCM6knUP3vQ8cz2Zm7FlD/Z2u689viL5VrG5IJM1pwrvJazNH3fMR7Ha
yJJ1WvPJ4U0rWXX7Lq10iddGY354ES1Pjob3TgHIdagVGTsfUGeIO5rePV8g
h1ha3Wkpavd+YSGjrCgmKraEtDiuKsqH78L+8yBk/54Lwh2krRl6sPDazfG7
uUAlMkU3fDMpAtPOAlqm8YQBBWNcOWNZI703HK2R1io6856HHg7WTb2UloYG
o0+/pGZZuiUeaZEDi7P2gukn2eDGa9TUBJCun+u7dkPkXligAr2FH3wDWKKc
0JhmoKWtwMziubdfE1MyS/96ImPfKaYaKl/35h6kBtuLWf/vZuK4mLv2xkzz
9tD9+qK+TIqVMkuOYquPFNEfEz72tj0J/WtxdRIt5nOnIPkoSpojhmmGP6zg
tvXfg+OR0eauefc1sL8qar18PCLDUIqwrE1CiG9w0dK5OmUXNs0MRgbbP1zd
AcizF3wlp4ls9glXn6gzqOiu1rTagKttJu2RVuScXz8Mzxhmpp68vXnM+YcS
T8tLH2/91ucuvfqZY8/f8o82x1nrndZEOyJoSV5DPiv2+KNd8QKASB4qEZa1
AdN8tctsd1iNRgw8soaQQFht77fssQ7PPTUPAyp50dRkZUjEeiyhRahFU+/C
HC1i7nl+8Fyx5GiiSDmv93FDiOiR/9ZfLhVIkayuzoM3h//RanahRu4P5oYm
tA4I//MDbxBYoWVBdfXS1ZUVwYxMi9fZ8udCltn4HioIibPfxpBbk5B/u12+
FQ8k7cj0W6SVpNbUVCulIOUOo6ABLtsrO6hzexHFBUs4FeOkEpagMyP4e9Aw
bOeykPwXLi4Ku6xjmeFjQEDrWPPaRQ1JeNSNuxQpF3wp4F8WVPCHbNam8FJ7
jYP0np+r2OEjieXSwkMERfa8jCcQJ9mKjO7yqN94k3dWtPJtMlbhzczciLFg
0jnpN6/Xxvk1lO5Ovyw+gvgyndPU9r9c4QMAThMwXjZmxmE1jf7/4FCKirpx
jQQMMU+KTcNjsxPahRnxEhTJmFKymStfuKw3Xrw99Dfw/MC5/SOF2r612cqb
DHVLI21F45xJKszJRMnlIXWBIWtEO7aaXvQ9VD7bbv06FQ1Yb+r+hGDDfLz8
zoh8i74XBoKk6xfQl2TUp7HMG3QxbFgw2HPsSSq89Pyild7Kvjr3sXaPxL+M
5HJ0XpD1IiRIqFz7crvqrh57x9QmzVNjRBozMG0LORQxK1zE1apdoDYPaTf9
FswcwVilFpydAwznDf4CVIpwNVs321rF9WbjlJbWCD4/w1cEnNNSgJoThTFK
qgQKedIdxd5NsnMKA0wiWDy7X44cb49Mbyjr98ndnSTMfEj6IdZDaJ9DibQA
YC8kn7F6+XdOxlnW1aR5Uy8uge9z0IjQ5gNiGwnCXAtqvYOdgINktQ7774Jg
qYrSiNp8Alm33E8OpcU1gjijHUy3cgzd4fDrCVCFOkv+7FG2G71StepAQC+n
VJxfhO2sT64u5T08r3jWIMV9zGaVWlIOJdbErcM0KcnwVAj6UPaFWhqZ/sBt
XmdwPpVHZubBAt37nyVt/BbTX9BgF8sr/5avAJzQLsbDKnjypcQmmhkhWXMx
byrvJf8uQo2jppcW9D6kjtu8DdaK8c5Gxwd1X/S2D+RNTs5W397qPzzJqr9G
n5KgnNcarglRa5zv622blaM4Io5Gn9hhp2m92pMRZCOODyiHu1QtOCqi8Q/Y
XyqhIS4dvLA93AzkeKXncHTuVKiW7AZfzU7LyMc/MusG47BAPpr0J7YxCa0K
tslqpGyBcOZJJcUkkdUDWLepw07CbvgWWpLc/is1mogggI4arG5cm2uB0c5k
nAkGCh1bEp7xguyRyhEMtYu5NHgyrQNqs8Kz+0/bV2fWjSTlpMjAD7uG1cs6
1syjngrEImMtfxVxPRGRNWHiwDDEJW0vyQOmbdxnaqmpBMT33Fx8IKY5RsV4
PCMK0bj7rvqt0MckywFuiYy5u5rMkTGDWM2UtUb9hD3Se7V8HF/oRDg2Ce2s
s5NdnRxa7dY/gc1Rhd/Ss7vKUmtZNOfELLDWTj6ojbv8Ll5zjQnCclXIO3jB
pmJDike18cRQS9imLvZSDZgzINJ2d1uGLig9Dn6QxnWN1fpTC7n2s166eIsJ
xwnHi1P2GxJ1EjGZyPnikDW4ksZrIlJbt1vdf1uMjQxphkdJp/fOYn3VN3hR
7GbWgggWAqwGe8coe1wqsX0XGOfHLTw0Jv9xmcYY7XkpuuTu89s1WAgaMI/J
3F+zTZ4tNUR2XFZiL6riX1huDNpaQXMgdgwHHUca/T4yoHtmZJSDymR2j0r7
RiBMe+bLDap5LXNVZXM3h36WGnIzNON8Xo8taVYo5KnIMRsmV2DKPKB+kemr
dbZxUocOfTmaLmMkXkyOylf0Yt87B4bMnPlPWfZgbPq+tDz81xT92alSqG4O
IZpiWQFO7UvpWvkw5+y3jKZLzCt2Znhn3iRe58jjGtN0EliYVoB04tAybJ97
cWQ7TiTnsXQqGIJNKOHpSR9wrtJr/BNXR1XRvsuiD9XFOo9zHPCaym3MX370
UjXwmdjkPlYOBUgIDYq8SZhrK1qjXKdTuZ+MNeXKPNeabCjRA1ICKuTPRAY4
8vXmAieaQ0GDaF5YFRrAn8yYlgyLOvpfDT4NeEf9RtDzN556DDG1Clo38dFb
UhcOwIoU4au4bKUcOySjqNmy3t+QHAFUaySabwAmtugn9r0hrW9ocopVHGwv
4DO/SmoUPoOsI0B6k3ghH48lkSlPtDFcIDTMsPaToSOxbZR0jqf2IfvtF69f
VMsobceGGlNOS7vk0e9gF4e+Ef5WlzSrykRM6/3a/Nrd/r7Jk4ZTBYXF/oVK
s5g6f6EpKy5ylXd+kWtl5sSFcPj/jWVFMu48H9qZqRKCJkARUvXI01wDwJjq
qJcdrr+E8TDpvn0Bw/jX12SfL5E1xdxDPU3LXcnjvPWLaxTMJXT4Cct3CUnN
O4S6/GYJgpCFlrJDpaCVVUFamywd4wlZgXmNGQ+5QNkh4bQrNoCX3SFF4gCl
I6lDInXIdoKWXOzAom4I912/HvBMPBoSsCac0rCG60KfOSHmAIRcIlfqpGRa
G9ckNAky5YvPa28ecNJfHZsr/enQA0qIN8Iqbf85+6waiWLrVPBx35R/qwL0
0odSYbHOYAug9ZczCvmpxCJZJqrVK+SX9OQMEdsG8+teYKtXzZ9xyevWNWf4
A6h+lSdx6LOmzrleWu4Tr0vFdn6wTKiJXCzBtGU8XhnIoT1FfUxd1mCQp8tm
wjSK0uZGPW0cxBzD0ub9DnqV8LFHe0bVrBWEEnBsFlnBAUeQr6GCuOVcC4Cp
vFckjqFylH81/L/A4ljmfyVrC/4xt+06VdhV0yfDG9PF/0Ub0kJnXHr419WB
NCbvWNlwDDqynUd2nKhqWNJ1S95Gyf/xVajt4na6+Ep5MonkH0jkDNj2nnNt
7FTB+8Clex0Is6W2fMKEoqXETC9lk3tuDVq5BUZPej4HPKJdvdYd+vHKiBwU
yvC3GDQ5kCZPKoqGoAbD06MPZEdk84BeeIs6IVyncQsmD0dJoMvc8QkoKuWS
Cp97zNm3CttkujzZX5HOOAeD8yonuOKtBCx5FC2FA+YzmwteiHXt9HChsFix
NbhoIWfD7ufkXd6Kpr2nHzDsVfTx5VYvbuGlAsyuWTzoAzV8AfsfMneK1Fw7
BRjCYfeCfB2qaGLRjBoImMW6vNK2jv1E5zvwlA254gdOyEA2Lp4VwfUJIkH4
hnlmCulY1m1XQEugC72Z80bc/xLlhEN/9RdCHGni/ME6rd5/FPmj8vPxdLse
4Lz5lRTyFToUbcjlRRejaOoF+sX4mWR0vCTcstv3jqRwmRgrA8mD+V6BjxLJ
20ADynjFwbBHl2igyK0xSbj+T3yjO9WEmqwPi9S0naghRN/tr3lIdN9eqFzB
8l+/RVjW+u5E5RwwmG0xeUbVFH+6GoHxvxg3DxHvY/NnM3V9IAADDxtCSdHj
aE1lH3bY2pF/8OxOQtZg8fteJahVe/paZzbNdfMO3lv+s4aLTG/2aYBLaoBi
MVaZJSLIsfJgf+53KAtxHSxzmxoRJTL5Hmo6RIyLHDP479U3IWTfvQ9lyoaF
yIJIx88j5bl375gmQTcu/LgLOJByoar55a4rOvjdKakn6ZcftHSz8DkZIT2P
Tp8k6Yw+kjqtnNtoYsonlesdvrX3e3E+YC2WgRx50y6U/J9jDBb9Ksect0qD
WxnTnv5Wb1G3fYIA10MKe4ZXIMo6AkpgQmqAfQzs+Xjg3crSB2td3A59Ax6h
Pb7kZfVxTHZxKggEUt36J/wiC69ai30ihXzPUAdeGYsINY57EA32DF3EByiS
yI7LZsN3eOo1MRp4My1j9YRsbulI/C79cRn1xHXwa6oCqZZfyCul34tgwfHh
9mu1PPdgbFsRzeAHgMNwE2EbQiROpfCrpmB8meuk3c7xnKBK2kSbALIMw1Qq
dMaVM4yUnhxwlbzFG7pqS6Hq+Y4eusQWTQrzI65BF3PMgA/EavQS8dnFjXdm
AUfuT3oD3hxsyo2kIq7Amh8AwY3Ut5hJzwiye/N4ElPMkOHlyRDkiIgCb64w
CxonVsArKDfagcB0K9Ut+LWA+TfGnc4SkmZN6ECLFsxO1s4NImkhgYcBoQ4W
+wIZswv5kHI+pm5yOF8vSEH4nPfiQ7ES3oqZ5SqRfcBiH2E/UvbDj/4WoIJv
HIHB2P3efYcOAyQLkHU4T3sf4S+Fb3alY7SPeKm6HjlkU1gY+ji9l1Posf5C
C6L5D7NvH7Vcpkw28typUM91f6FbHVDmWItxSGGD3eJ8qqG2gWQeOURtLMuW
9Y5G9U8KvZhWtWzpc29Q9BPB4Ko3eY2StSJ4xPpVjitu91EY3Z4IFqJpqM3C
z1yDjOlpNhZT27CFe9fRITQuExn8hcRGqCGsT02vkayyhmlQSpf3d2cgPyY7
55KFbjabX98mVy5Xs/Zok9/hx+e4HJNBRw/2lSLCLNimbADl30+LSpn1L0Eb
HTlaoHTj+tZy27ouRFf9BWDEnC8VinIh/jLrQ9zgwPjKDCsiFeQPotlZg+14
JoI8kYzxV8+kag8MDwb9n8Rn/4C1Llx1EORxNzGJcw7rOnNBNeN8fExo0Upm
g7ra2JNZTrSEeNjCHUjpUP9z0H+4AGdhbKzGhSeH2j/8N92xXtkdd/wVIacb
hIfsT2B2fDeaHM0vV5xv4ke/zsHJhfDZCBLZw0p2F6xmfBlD8ses0UsHauby
5jrTiILI8QmB5wGh1p83R2Ev1TcMwnOtdrfmC9i48PJOQKDaI+yc9ayioOkh
iy0CNDdi5scFKrjnNfZ32lUzraPX/Py6+WTheoikjercI0FOePWOpVGY9e+H
nEwj6ymXeVBTPO4nNtui6LOhiam9DKTH+pllEucUMyeO3ri9p/x9ij2/sBKo
EBdfifjpVigIxFVu2tINDYP+5LXkVHzplvxmnHZ1B703bJsO6ZUeyMdqwr2D
5pBhtwsRU3y2El+CTxf5IUK9c/jKgpQJCHbr+EgVafMrzd8ZEPNSybZFtf2d
+aiycExvqK2I6Vkg815pYmyXLpgsNUt098v03lN6/b09rIlFKTwySxigHY1A
d/gZ0OSs4+kzFSy96eX3nygaOOUJzggxEbT1vnRK3r1j/NbcchtQk0hNt9PD
wuOL1Q6im1+r23Zy0Dckc6sTXubPmuxwNDoDsFH+TWpYE075jGANV0k3LiQY
soDaenkBaQ0r4x8oelrhQLRSjtVQuakoPL7PBqY6ONTlBsVYIgArUlFGqwSn
N2AthNEJTVudoPysuzTXPfz4CNKmUbEmRtt5VZK2A/aPlt6PtWNQV0QLY1EN
pWs+uleLDu/obxlIBfFQcyPz6EfGrpbMcqT1EYNAVzoHbs71VqfwlHe3tQzZ
joYhukYkcyKaQQZslpCJqC188QZ87RM4iChs00CWiBJYQOu2Qm5Wd7/Ci1U8
nlXiwNzTUO6VpYumS7Qk9rpsD7NOwEpcWmL+d1s9St3+18stpBiIhvIaq27t
OEku3RnRJdBbtzotbnS82dSJ7mA2xzVcJhmB7iJMWfKIAZUx9zN29yL2+m7t
0eO8+8h7LUsVdF7cxDzYwzc12a9B5BJV24tUjO+XCgeGJBqTHXvIT4ubtja1
DCk4lY14D0juxmEoJC3wXfqNjXNtENm2nhWdl1JZQ/hHvwvyeSjPz52GTg/t
txn+5m9O6m5n4iK4B3207toypb+9T3QMWdBWX/HrSEzIgmD0m+7rNei/uSw6
T6z1ogEqBSk01AqQ9AtWvO2MW7mEmWoeKTCDFGcwtHakqOV3xPk8pFNdVp0T
huWlkSbCk7FcAWZGaqEvVGGf/4BEwIcJtlne+zdD6HnYo36WYtP/b95zLvh+
VELLvQMOzvoqUZZQb6kToc63NXW1sAAK/yW0yynDZqW2pwOUscBBfdP++e+F
YtitNyaBGpNMtMHKCdyvOikcpgtLjwxdSeTvtrkwHCNgomsTbFloVacdK3N0
nKCiVPEMVleSqQyt4jnufGm6rrEGf62DLU1gwdssjXGqSv33+1Cc8RpSCACS
Poo44BSn8eP4IxgpYkLM44tsOF3QZ5n9OLWarQTOsOdpGUjadS1C+HVfjX5Z
z53o6sdj3rBdTTHhdz87KWN93INSAQA2FgDDa+ugRD3ii6ethbaFP8zKJ/6F
uBNjAUx8qxzD9cbtl2ZAcJmOIzeu4dbU+TCqd6YTL0GraLABbX+dXDVUO/de
jME+oFVXEwgNK+LW3dfxEEZW2YAlW+RWOHfGD+I+tu54LXJXDrshcGNlmrXG
tOLgjel7f6IJ8OcJdo9F8/X/iccrGbNzZ74o6b9gYQYIvQ7V0TB7DSwAeOqN
49JPLyO6JyUM7ktSnZiJJ8m0pecqLgv57n7SvzZmaaEVLSzdpFPnSkcbL7yD
BygLr7miUmRh6/pVqUzns9lrW7+lzL/nbmh3vuyjktRwDD3j5LxBItcoB2dI
x5ivcB/OWTizDM18O52ddXTZP7J4/49oUOTJJ8x0tHfeQhszjI2EZi1lEX9p
SsQNlbWZcpS6/QlUyh/Yhcar5MAusvs40Xj0bM4I5m99fygFFJg5XRk1g67F
YTUUG6PsCpNnyRPm0bC1lTuQ+EF3xmiJPlnylWip+HR+7LzIzHxAuBvLYemT
UQevP0GAxKmTSx28JV/gUpgFCi/gm5J8Xl7oFX2HU1K7VBIN89JVZzQ4/UcI
diJ04nRjcsv15XM6+dJw5IoYbx2HvfuTA6SisZFrZiGQs8geCj8Zw04ahdVq
nCcsMaUQE3yfjhBVx/63Z/zTSViKDLn4MHQHXa/3GNir7NCOi4RXIIZ6+EcM
8VVweFUepz/aYLPgxyfKxigrITzMhfOZBrR0cfT63cLKw3r2rN4QmpqcMQnH
251XAksWkFXF766za2KNxAXlboXMXQBlFyrekbqJY1VkYNTp69MqLCsXfyvP
hb9pq7b5D64PBexzb+plpu7KyZelqKX+TjubSu90eA/LuGTdwI1PQ4dSi0R9
EwjEmtixlqOZLvnnIcQUxAftz6eZNHIMFDfhkrHLr5+yaZR5V1I4UxOfs5l6
QiibBAJ1PCdAykkG5qN3SXHoQqybl/sJLJ3D2JlA20ANRxYL7h15SD57yKj6
18HLWAT9XuBOsBNzDdcTPp5mw2lC9upNsqvoHf9y0zn2vldrpDqnRc5ZTdcz
U2HTlNFBI+VuTdWEt0SB3kHYCdp/gZh9GeVg3F2h1wh0vYl246W526BLmoOP
WmnhXgCQicpmu/kPF3/RmGFatBgglF4v8e/666CQ1nCYzz3FL17g2MpdwgWe
6TWUtT/cqTjNCX8PsCfhefqIaeGFERSTnDa3YQ3yfxrzaJHKxGK0c+6VKLzk
uQJWvBkQPECeI4DPShiL6+OWh+UW9P3ciw89MdhxPBzsI+mO0KaktIW9JG0r
ifkUQVGttPrAoVYhI7EGjpLqN93N5+Q7RVUz05DRExdXvLxWjo2zPgGksH7l
4wG7d4ZIaFzVJNpbEGVSr4BsTWeD8T42SM5xq6v4bIDaoxZ7gh8TugZZt/Y0
fcuB8AXDbejTXz0sZf2mwVFpqQman7Hp3vJ2nQGfgTfPaOMzbZsWNJBoRYle
NCwAlD5BB7M4qsb9JLKMRPG+4b4v2XlYbDuTPpOPSP1rZoINPduuCP53/8C9
P70TFiqJo4rMfZP4zb6EFN2zWsaWHZDSFxPI5O8+9gf72UfDWKQ4Zvx/dVew
aEU3sDrGYQ3lKZbUKNDIdXxvs7nCCbMiOvbbzkkPWA2CDbtTxTQVCtYlvD8b
Dz+crLORB91uJo47FhQWkfOFbWf6aSA/1lCzwdf2yQO8p9aJkEfzlBjVKKw9
HdXLfQAh/5AINN6Ei9PJehwNxLQPjVTSsnP/8tCNeBHbdxcNVrKiyR5E0mQB
lNRefOy76Ub+f4NB32fg05jjug5ymIxZBM/3UE7ZR07QDX5jUUTYKPctwllp
+g9XyXr89nRsetrGXLLHDp07bwNTnZDAMDhgYqePaHjY0xp2yHa8bLb7V/lK
fgmieh0pk5Xl0ZExTTd87qn/1ptZ/8y+CHPlYXT9by+uz6RzmIGM3dEHW1Rm
vBz1gWciuAPokYZA5E/uYNIiUmN/KGGRBpHdH6dxmlAmptYx8s+owo8nGIyp
18qzzhc/SjFaZ7HESv9G9iAdUWdRW1a5fCgNXZiNJ31nom5VBBTgHzS/kzU5
D8JPEhCYIjFSsZjO4LrfF2ewZlaON7/ZDbJVM3/yoc7j/72Ob1wuSllBDrQp
3TF0F4b0T1KSNBdKpfJXCMqtSHgOxNSh0vEtFi8TpZtak+QFP+lTai2fD2rL
Wn6x/WarWXbEsfzVyzdlDm0keIewkPWj+n/4oYJcwQXm1af8skv09jYLeXEC
ley1OmbFKwGu7ltoJSRCTxqJ5+mtXuCSCQspP61+utPhk+SOaD5+q5Xz/2Av
e9sri5vr5re5XeApI2Klm2Uh8flotDrrOr/btuffWUYVmun263sosimFKAl4
5LftRL9bIj0m6HHi2xuHwZ6BWWxcU3Z07a+aTogQhcE22CyikgcZBdT6re4X
4hV6q5u0WN5qO0Caw5zr7/lvEYJMQ+8n9aMQqpxdgZKxTfXmWGkVXqz1JCjb
WBkAiZOf80xCn1nmnVvlBWBqQJpgokk5A/ydveyiG5UA8hZlwSpgpgpa2taB
gzoGlzVUj8Knw4J1On1mgiDdzrP4LtjKpgxzDPuGOpYJ1nnDMb0QfskRxi5J
0WlF1vK5fytrEWw6mVCVmV+qpPwgqjxfPxZ5KMxwm3hfED9oe8E1loJCHmK2
Nh6VExp8xfppbk1YpOWuhgw5BaiNOwyCMzKFSeH4am6NKCAycP6U9QpAbkSx
ltErpznd1UqHYkTxV4wdC7IXeR0TIOCt5zENystL8JH1nA53F2fDLd0V6akJ
rI6+aW1GY/XsXVggEAPOIBUCfh80a7Qb7kTac4vdxDXbeNXk/RhfsVsStXxq
wDzJGlQ/kdckaP+DplPJ03CvM1PLoI2xn219DopIX2LEt/k6uVCORoZNO7uY
/kWQv8UNosR26chE33ESE6B6R0qTtOFbq32APdh5zL4jhpnqcQQP0HFIu4IY
FVTaqixn/nzH3w1TrwSOFnJHaakRX9G00CNskuBwtQmsyYG2vOcdP4eQWQmM
P2jzav2fHaLE9QKHQWnqbBG+kLk+6rlAxfdBfuuL13QMZEyCNT13xYI0cdxs
yQCpZqEWLY0M4BRAdhP1c0y253zPwawsOxbIRIsw82NOZ7fIUS+YGngPqp3A
m5IHe/RAvUwPUOwirYd8o2kWKHk3bgGjUcKAkGohuWPtzqeM+oyP9qqZ7K6B
P2GeTbWcNSWxswG1ka4Dk5fI7DouKbBNWDkZmV9Vpxi+/Kpvp1/wtiE/xfES
VZ/f/dgNj1hbBZFxtsLtvG+YhXep6Fy11iWbWiujPOFsCR7hPvRjRwNLkKxa
3/qK8WXL75dZUHlzCrAD72D0So0kZPDJZSpqKx1iOvRwz4sBXoBNbbg46Qrh
M6RqYFAQvuNktGJNpLxzrw7M+xM1sQFFRD893Bw5U0eEf31wefGvpESX2b9G
lh3SB1whgR6iip5iutQ+yo07wQ5KObWuPsJQFEvDeK9hz2M5NJVyj4U6btPX
LlJb8CrZDgtzaaZVrgRemSROfrPiSqvWqa7qqdJI4oG6/3EI29pEV2VxuGQX
75ucmxptCdrQl/SawmssTajmw7FZ8tjEIhBX9q1Em8RzpEU+yzZGHO8kfwUd
YjvfRC98WLg1eDW1BgKcJiQOgJNVDAEYSx74irout7Z5KIfEWcFMRLsKPZN2
3txBNpByOx9AhtEKff17aOVgMvdjUWqDSl42O4d5DWXnN2RFILCktytUnEof
BToZp77F2FvrilkhR/OvyE1PCLhRTDrXLFLdYJYJ4FfxRG9tP+U4XKpwoJRW
Ulbe872ACShImEnDa4HNVFFbWaAYRtnP1uxuT4HJ0jEbwS2mPE/qxX4zak2R
9GFX30mJW0VObPRarTjpdMfi0Tp9zBAUDnC5FBplcdQOM5zT0/zjpbvgLpDk
DXnA7/ALDSffU6I26Q0Y6rFB3Pn8QXlCafRc/W7LJ4G4lF33osmMB5V+LLeX
1s20C3X5AdqkpdQzO9hwMUs9Bc8t9ovw7uqzBYBZNW5hNRK7JiJ4NucLLHKT
bi1cA6th1E9wvTbUotJrvo4Ov5bqfWTQByRzXFYdDxD6tHJNWV+JAHdjRx5R
QEi5kDRRCgkPIKu//sXiqVs+46g1cHnt+nsLSKl8COLxjcpoPg3SaN2QWQFg
jqdNyPDGWmPhLrPI2dTTrCVM/NdwwLD4SPyzRGn9L1FNvlCg/kGpBm5LySKO
Lv1fcNQeFqdGE136KUYXdEhRz2ZT1IRLw2hBuTYHOQ+NlbF3UClgw6g1+6z2
oMaaPbhw1ThNFs7tpxaPA+7mgB0tGazvnjkdN2++YAPWp/XFci7bOE43OaK2
dC6Vb0F60kUIo4uY1Qf4iZ5Sw/nTKE7W7cmU/6BPSpevP2VWBIXuAMXGNKGj
UzMHZh8Jpe57A4RC3WGX1n/NLTaJzFJCopabARHvlxang6f+4XYCRWDtOj2k
DXwEUanIMfkJ39fb2xaGSj6WREBFeeUVeO0UDXYQseyROwoZnZ5jvhDyDNLZ
E4INXoO2MVku4p6i/EW1UOg5KOaZz1lsOmLDFq5clpH2oXBLuYZYUiBE/8pL
RT3WWLjgDUHEx146Xb0WmGdmtK8WIkW9SpPvF5LebrMO6lrrna+zBof6YSp3
2fA3WVNS7iUdVoqkLBLwvWSUbFFcSAv2j3x+8fPr7eOsROD3UQ46up1KdWr3
LFo/cv/3paf9yPHqW8GFEPuBEsmHyjEKyPU+GxP7WP3cqX1iIO5cYl6S6O57
9tlbM4+WGWzLE4uPhP4/OvsUh8Fu2iJOynj9eWPPtkXI6Isy0Y2Q4XscS6Tu
zeet8+1t+1sB39IcNGjcR91xSbNZEfTWzShrd9kmWd692mgJskcsTfsrficg
nCVfXQ8pTZCvRLCs8cGWH0IuWJgtv/6BW/o1Thi0qQvuqWMP1QBcK7SilNSq
D68rX3o1WhFljOM6yZJgDfARf+cBUqs3on9zFBMfU9mpgCH+yMDpKnoMdKHU
Iee7YCzoRnlFKP6vkOmYwLZwxS0Trtq0IODhx8Z2wFjOmGf5d700FQhxveSx
pkskOgq+dpSA1VOE3Av5Xk3IXp/+3UM939QvBGUrjwYI7w0gg4etpQmfPZpA
pU2gKSQUDmXKovv6U5faWRw5tch1+A3tir8FkUmHFqz4zhlqOnzKNTtKAbUZ
ySYvgI0InWVcgzZcakS1dRYdjJF/xJ/LHMnczFs1nChr7jzAudjYGun/jN7X
B5WeMa9Z+kdjqAo0YHMbaVvyRuSQLDNYEPQ5IAQI8x4IEh/Z10JvHh33iAiS
RVHTLaCtS4oNPGCvQTL71xEPcNk5grltks4rLWoTaOXsRxPH7cqmtjbEnZ0P
jgFy5+sZ3JDSfGeNvWzP1pzxNMBDn7B3UoLp6Fdqays5vAJuEw6e8JN2C9qO
3/+7dNJB6e0UxfnEWOROKBLq1WffqHrAZq9cm6YjoYDKfoweeRDyd8PW2S9i
R2nf1l2xQ8ENU2itWJWMV67dzwQZqu9A7vk/Z93/VFIdXsuvcWSsGJjw8BmL
Le2/DoLr295J17Hs96xPo0ft7ieeijhpXECFgoYZJl59Z1XGMFVMsz3GWzXU
rH2rzLueNsmCpE5e92/zMmFJtvgxbHxurYvv2KCjSMfL04gKzGPowBm1K6n1
6w14EOIGrRCkEq42ZcG7u6gRD7V4aPgjKyzOLbBOEO7F4wlP7cZzd3kDwrV9
30aP0NLY7F0H5TufhGzgbLTwNi3G6ACth0F45yOpVxExw3jIga4JbZH+045j
FTZIZOcJ1N5V4JQ7wz60E2EnFpPPbl7GmWwk8w59tHSjTfpvMX00HHoSTvXZ
7aH6Hqhqyq8CVXxqB4ylBogcDTfgWlLjlcXROwCMLNEI+URiPVQFZ18KS7wM
783jU6Abwf0dPYUk5AvfpZMelb9inrDSma4s2uj/JnOsMIV8i685tt7YqvQZ
pXioke1z9AWuFM66E4SwvhkrgM3XBuULZri+F6HeLEUFnkQJfEVWBO1IKh4Y
TvQVM2PF1ttJ44sdtTPuQJU0PP923Mw/3lux3Mjt2Uw80wyTWXewS4SnCUlf
Tj19E+PYF4O47GxJMdYxdnDvYBPf00F46ztIJg4BTC/EKyAQEQIeNHWawJh9
IwyQCfTx6XhwjPK+bXr6wDRHFDfu96B23KuCRGFCzOaUylwyGiQ2VN6SKOkk
MhOZOH2V3szdfWfZj3zTiMWbuYt2GR53iVhYcfRQrvFXhVR/+iRnvuUoFBOt
nlZnucAL2d9DT4YEwJbfwk+BALiAD3jnwrrIlyKeLPuL4SGUcvK5zfy5eYUp
jSMvDykkNfnePITedyhENP6C0EWThDlSYv5Zt24HPirh1mtG/H/Luvckf33C
qPHDGWEhZTjYK6Erp1tZruy//w/qZTfLwfukE0rf36JSk5LdGfKWeqDHtNV/
2sZ4mdnyEcc1NHyk2YvOkrHtndN4WGO0CvCHoyg8rZ3kr0PNZCQPqgbX49j3
jBPDsBv0QwELx6AF2MnrRZygFGsNUb6EgdtN8ZKSwKlxWtcM4B/Qu2uB61CI
k4yKKCSV4cKRZ2OLE20hz4FnYgCDiAZ6Vp4oTbFwzoqMo9IkvgZBvAIHn/vR
pAe5Z+GQYsEHWkw8rb/nRZ5fn2U17dB9XIAiS1Hu77eciRLUFxF+M9SdXGnS
KPsl7snjG2EqEMHMGbE+snPxDfyjmelaDRPG5cLwrXg0Pv63llQTGsK0Ay7v
I5OWYhuuG4hXt+33pzVj6pqiH7AevsD4sPm/MuraE+1DJnQtWwxNSwX+DYQo
yInWBH9VgoJCzkAXHnTqwMCenRq4uBe0RlQU10o+llJni9lT6VU0Q9cui8GE
sWDn8q1d5sQ/IRHmIRC9PEBwjAwc8hsaxL3d08Z8eFRQcg8BvZEGOUXFUfWC
ERlRwtdht1w/1xP4yjQPxcim71uvaP8JwwcELvA8LDgew8MlBhyJfKkZjRzj
IKP1SiN9JtlPnpjhbJ/egDzwQ/q0Hr1cGlYG6f6T06eOexAJCs6vS8ehVSjo
BrT+rXFBq6xbBZM90FNc2TIgroR3bA36JdzFUupYOGtWUzoyT5vqpUJG6WN6
VGNGaWPkA7P7sDJzWu9JJ8lqnSyvBQFMvA+W3hX0xsalSYesZO+X85MQ5tg0
6IOau6O392u45Aqh7Zs6MT5SUGvlliMulfnyU1obvu/YYtxxQdPvk69cJwQP
W249O6eZSCraIQeyXO14xvEzD9MwE2IzD8z6D09MZk2buPjKKBpC1qAK+lPK
FNG5Dm0mQ4MowNpQu8tmQePeLrwhfug4MPZwbxoSR+tXNwiAFJlF3id9JjCk
9dxrHWV68kbu9iM/s0KeiWi88RqkrHGehR4lRzqvHzPScyhLkDiFcvT9my5b
k2sqLm7wbqbPOUUf9R3/igljupai73H1eWYIhRmtbJqa2GX/o3YnniLaXdef
yBs91K9y5Ftiv5HvdLcsFq9m3SHrpPQldu4BSmk0vZ4bGWG3KlRSYskxzYND
vquJOdaaq8m//J5Vhyy0idaPZHKuIhrVmZBhqabIA/UeAW+7BVvsC5I7Dnwv
iPUTAfWDbJO8sKRQprG0Cw8/rFdeUQ65i4/89SrpylhMZ4zUrDBekoycFAzj
1iePmVWriIw3zZ7QWyLENHI6Y87TyKYKHAKmYKyn5JqDBdCVRFLo6I4wUNeV
GyQ6e60sQKUlbXaCnwgCGF7EFdtlqm+CYHesl2NWSu43AM6q0M63XO9cbKTL
9mj054l+fbA8y2A6/h/VEbbMrXByi84v/lrIvip0s2tXFFoLdFcg9/9Sb0+L
773WxRT8d+XrnVsEwX5tl6dBreAJaK4hwNbIa16+WQQ1Vs6Mi181+VKRp3Vr
CINX0tBSoxBxPh3i81yADgWecHRawjzBl/TLWKjUg9VsiE8Yp5LBZLXDruXh
aXA+idb2IEBDs4ligTOC4E/jx8NcBG7CTp8fy2BUzP5tV85JGIEcGNlczX7F
43z5bl/irqBK0DHfHndxSQAr/1eQXA15H0U1U76pzujxRg5SRolj/ZZSX9PV
1idfQxbBU+ep4dpLt5dYgyQWjTV9b/6XzYH3X+rhlu0FuPwzXEDGUMKoG1TY
lpjWm6yS/KaZ8C9Mt+/FrlOA2AXtOjpl9z3YxoNa4X18sqxQmzkL67ipXssh
MnmCHOx73WtMBRqF+iqldvTuvMywYgNiXqomwgy1IXKMcGVQEY2oMz+n7gFC
qdDztBJQk/mSTtSs5R9zlvaU+6ErD6jFf3ywWedoVTEYkqpE919jQSFEH75m
+LrdhDhl64+YLPZnv4R1s/Ia6epYs+J+6izcjJo8yTDCfGsrunPMIaXUigMA
JQAMgDdakJsOiq63GlaBVfxaPx2eLxbylT9SYzu9y+TSk3S5Qd/KKkWxHvV6
kUg0SCVKk5dKtU2QVecs54eedG0t/ASP2Orekj1mi+iuTEKq1zizCJPsz9Ph
hW9c13iTTg/x633fkldr23NORG5rcMKJgApYUOsKTq3SoANDn9+pHxgl00RA
3+4EtCfZz/5+KkYFssnk5IKQR7wD0j2Io5yZb34DIkkytdQhFjQu17Exz3R/
IWZaAcR/d8I8BLMFZrFItfA6AsA10/ivnIj+NlW3a1bWtBr93YMeA87a4W08
WAEl83+qPs3XwXLyKVDuaHqhb/oj6ZKtjcAY4hz7LMLZIJV8pq9b0xUKxGJM
U/gHhhxAWFnWGQpx9REyfeVo69LQYWS3pX/5mN1DCIaZtcBprTP7+sAUuczu
QITmGWvmdbvmYPuFNC+niZlxmm3Pd1DiRZSHuRukIyhUD8+rt/+8qqbg4dLA
8XMvLPENKKWNhQtaF5bd4YlYUCxRc2j0wRlTNO719Ik8xViXQ9XSEem507gq
if31yikkSkFcqJTmJi91cb6ORffQ+o0kH3DGa3hiKqCgqehbJ+nuMIOJw3V9
ofGij3KjU4bs9MCptrRWh17TDrctTxAQbri2t6mkO8gbj3Cf+0JY3clv/3HE
xGka9MgIqtnSIRiIWQi74vauwZkQpuYWkuKJ+0qGwP6GTDDO5qjKAcOMhu7a
jBhK/17GLI3a4A5c8qbyCasZOO8DOoTX48YfoFsE+B436favACzQhTGumNkc
HgXEB5sv0EbB6fC7gyMtp8mdHg6aOptCkEV2JJdTteH5lR2UMneqVW3Zm0+M
5tVFjG5QK/hByrhrIPjFwpmG3vXhFvFbSJsMy+Oq/q2fsUmPekMILTo1T2/2
38awrQgkGjDZq3s3pJMBLXl+938+RWvVmnGbDh3lmiUKO0XcocGOuEvoEJUR
U9C9446M+CdWGT2qGgjVV8bmKHimsw89uu8tFSEN9z0U3FAw+Oppopbgzmcv
LtvzGXiRk9fTKLhnGXMmFK8J/JKJZZLkOE+ZAT7bwsE4N9BniBZEhlur5GR9
hA0FbCEaifAUov1YJPObmTvUislC3/qpSmn01KGPdezygajcpLbFtfJfHBHW
cdxkyx0mBeZSAjhwm37pLdQLTkom0t/B/+ZOKoMUO2IEgygZGoK+NIz7A1Md
M/AGfr3hZOLIwxd2aNmRcnzhmcnPIkRIaIFxxoK/F6jIgaGFeEPyvmkxaxIv
i9c/iyXcEnyZRJ4WQDWsA8ZtbTNS++pneMbcyvIR1LE9XUS7R3oCgJ7pNsYO
rcYYMRax982mawFVZLSFXk9slBdkI9qWneFX2cUkqnusETTAVbpO2VYKSaZ/
el1pBoirQc/2gjbB1wrphI9p6inDQzB9DEcBXbBN1qWuob2qiUyZQ+GKGUPk
SHryZGx7wjjUf2sG+A9LSM7EIe5G88St6SYVoRmjonqruTEMutwFRei/Tx+U
SOwGKH4U9Cdx5ZgUkxVCjNTano7J+tF0ttj8RzN1okr9zXQOGvLh9zwc8rp9
zaKtNpEVxknKrjgOL6aTNr2uF5dIcDUiM+kInQ71UETtVk6LdBCjElZix1Jj
DPWm0L3iv6ejZWZi7///fkQiunCounY3Kr6uTy9u8u2Akz7SUbMYbK2NRDZI
HK7pgJFNTY00rGaU4TSIAxtWeSyJMRZBzjaGN+lqvdcplq5TT3Ul+VWozXyl
DKIu8aPt7chCkiPeFdxjOp1Z48kjzxeFDvx71olyyeaRSPWkzSpC7eNbMffl
LPAhCLDNMTFItpH7SHmjM3sO4orzcFP5/z+savA9lQOgL8W81mqNm5BWQWfj
TeSWjuP4SQjN0/MX5zPyMOgFGZyxLqQtT4g6h6VGa2QsaEVgPQrhhg2qzby5
FkJsad+gTnism0Rx+rKhXSRysl0Z1BcOlSiKvZTenW449jagjOVT4tDkBN+6
88H03+9r8yI0zxvQOJ/ASspB30GNQ2TChbXKZ9OP1ReP+q6K9hivUV+JvGba
xAFS2syp0IMOP1ibPXijZYvilnp22j6pVX25rj67Bo7cE6rxNDT2PMe1eXUG
iST8ejR2SBb0wsJLLXcobqPTvl+KI564MsMFaxHeP702jOex99wX/mvoxzTX
5oWs4QXkhCEvx+5MvyQFYirMz38n8L55FKgbIvoWsyupNsrzocOkYD1J1yDP
TccvT5HHA6ZAr0FDYQH2tQmzw8zeWjMEUkTdY7GzzTIMDj3uHcx2669Q0I0Q
RvwvrALJt3FU+ZcwO0GhkKcQDpAmFOpikr/l3VQHtKAMwkjSuil75M49ygk0
sZIgBhUZ2HvHCoT8vhr49hjOFhcid1zvIgiMlJIDTTmcLvp8FBQVIM2cWKw1
WiQPi/pAvuAj79YGW2BZhemE6oRLv4dteOkn/vx+Fm+wzK3hZmqHGIocF6W1
L5tZsuvwyludx+0TbS/L5V+7JFC3RbnfLcvFHwH9jsnhE+a3EZfLcHvxlOoY
f26iFOOXe62EJuM6KJbSnJxOHLhVbgygct2m7e/kc3S2yareL/ZWObnw8hQ5
dw76WEXqWs20VYCMrkVNTFeOpwsF0TIwFLYWjmBqEE7656PTKlqol8CPMuj4
utUu+duBROrEMYrowNE8mnsMtDnDtni+7m8cAZ2NTXzTgEK5f+xnNf9MFSzt
1Y2NI/BB0ze5HLnccZXncwcIodxJJQ0NxltMGwm037YzW16PRkYV0FiNkXci
CuxyD4g/z49q/e76Hfacvb1AfEnc0dRE5q5rkFkEwaXXrT9iotnMUhPrLIdO
rbTFnMhV9fDczXgHPoR9rT8h9NlT2pQCJ9I5KTslV2gaE6UMe35gENKfMAth
W5m2W1cisetzjZaThQAWc1UF5L3K9jnrsAk6QBtUvHql9sHN7+7KhKmjxESU
wV8omVKXDhQCyNMIQnVgzd4oOyD9MsvRqNJwIEwpYC5J+Vjpo4HIDks+BisF
qmMg/AoXm5tZZw9wolPX7ZNZFA0lrT3ox21MpddeAHQ9MkOpU0eAG/zFQF5M
RJVl6yXQYh8bAz9cCJhRYAL5U97Wk5yNlkiTBXfbW2ryqFfo7qO9AQ9C5P1D
s64rc05QfoQDNenvHj4wkZS+Fiwz6ws95smzhxM9nQ2uYYwS/ZlWryuBlSpb
ViWwMXWDcweBAoAJhEKkLSJcO994LpDBtikcWuTXtLSNFGolfRxjt0c69iyD
F45MRbiV2Ot8t+Ny4cTeuSRBNErAmKTEafT27+Jb1vMIXn60RGPyd4lWGc/x
RkA2O6f8iHFDeVNznFJU6T8a++6ps8U/1VGi9kqdki+BVl3e+RYWYT/ee91n
39wcTpIF0pI+0zLx+kA9NhSB7bXl3PgLpADn1ABUzxgsK2Ajvff0aZvDDhkr
xTpgiAWj6y7K/gSgYizqu2kgzqU1N/UdeQeyFIkHPB6ZUZ9MLVNzPKmfNXt1
mlGrrKuSunJ+ND8sa/XmOb+sVAP5yC1ixcXuvBNea9tisQC/sYiZW2lKQm3x
5M1Utc30h8OqpTieCuK2qYi4P0v/Leyck/ah8iwLXTjRZj1FF+dIS57s7dOx
BC6QjNL/uBajHQKgaG8JfzRqdCdZsYF2xdTrCh0dzwyce8jjXqmvqE4hNJYY
wFX5Z9JEaDq97QRhnSYsiNxxY15Nj3vHK7TdxfuSRH9Uhtqz//L7MLdfRAuU
t27sVSAXA+UljQH1pk7esltQ+6B7yMO/a4m8Khuekk7m7V5vJj5inQQUNn1i
yQBBtKLavVz2wyEfHLbwi2SwARO2iV3B3F3K+VgMC5LX9OkspMOkwS9HSyLI
mdSEjMWwFBFkJHxZZtwbLZ+Go5ZKqJheQqxEq5Z46/IXggqYkn0yG4UvJ1zo
khe5hTCfnhToicpzRnTwW5G7hdA1dqq7DV8ZH8OYaJ2OL3Uwp6cDhdMHeHsJ
NggvofKlAGVx1BRe9Na47AuD3GwZtYfAY6XR8pqK7LadA/94w5CW8MwyiWYO
nludYmjobEhuy+yHnBPy+7jP9FgMBGhbxcB3CsNrGqBXgbo6VKoqWcGj32RD
5PwolhPQK5nWdTbS/GQ8/xz0Ql7pnUBl3ruMxut+5FzWZVDqDIxIN3gGjgfb
qPA92N5NG4wwPf1fijgUuPtNYbfdvmBgoJdfo5dHauoPbCN35Z6QxCiyveTr
96I30xofHLWxU2ZEdr5sE1xKIP9ZaI5Oypl3O/SgwaqKNJpxgPc3jSb3v3IX
HawdiyulAtX7OL1uOxnYTXOs1W7Nd2402KkQN7olEBybXip04p9Sk7yl5tC3
qsGyQew+nQCQABmXvvFNcY12bTD4+JcqeCxLoUnTVb2VmB0J3P5cSHQfxSot
+fHP8VqkFRKsolehSFBSkhlm1OPjVa7K9E2zhgQhFdR5wyR38csmo8XLhud7
AhcMjCuzLHcqZ2lCDo7v81nMBiWhIkAzeZVn2clPXdUJWJNTulewttjmv9nh
CbOw2O3EnSJMSF8mi7lNuMPjfUn/UVOGg3L+fXn+IE0A22UYQYn1ZarndUQz
va+I7W9HIbGU54S1PSn0l1JeSKMpptgK8D0Vo8I6gvKE1sMD4BUzVeUdsUi2
xLtocBEuJl96TNgr6cOp72yHRFqfdjwl5+VhCTOmvMigVS3RM+PuECyZ6mVd
T8EHtbAjkMu+Pr8V2flkMajIfYlhyA821PlrbevszepoVV3inGLJEr2HZRb5
gcbCVlFwkVjX7Q5xEhNkJHSEq7XQVK8To0I3JPeIwa/Bowhc8g6b15vZZN9h
PYnp7dRw/1Ce89UHVdh1+yr+YmUbIGp+vAbEdVprSkUt1LU634jjcFl2cSeS
lk+MKLkWJ1AK4t0ukjKGZF8jPdFHXXuG8GRUs+nAtkUXBc9UKP8h3pE9gxLU
43EkBZc7siOhILqM/jOV9dBh06w/bnneXYCzKGKBPy+BBlChzAv/pAgfLop9
wQF09wFfj6A5LVzvbx8PdkHwEVsqeKFSuJ6aavrAb2abcTDUQi5xPC1eOnl8
Zc5o71PBh8XgNPrvMj4V+ptvPSUxHkYFGNBpvidMx4QkQBAf6rG6BHKxVQAG
wLzIwHMh3oxemYP6K9MXrMTXcPcx95WBR3fHxZvqYUt+MPcwmBIPNwJ8zNcj
ZBcEpFWoBJ8dLDiFtDaf1Vj7fYGZSs/U25L7oVbbepHaniHxOWgV+sWUNo+Z
ADgBS89KyDY8Hr60kca1sYzIfpoBxTbjCPGphaz+iE2RoNObV7ZmyfnLEVoy
MLMOqw/khtb7dEAXyVe8HkS5wiyod5sqFMnoGS7FOgKqkt4fbWgbJoa9dg5h
Btquw7xo2irWPk/dppyDYJB4EoYGidcVWkJZxYZyf/eD+6z3yWLS6F8g7S/E
Rx4MDHex324nzT/cwu91w2aUIgIMK3lzTh1wpCVfB9Ii+ghA1OOc5ZfhSIzH
WkCyVhEOI1GbAYq2yNgXHiFZVljfPPaQTK43n/TW28ZrKo3iom3QjyLKsBRx
OBdyj1uyiwUcQg6NpvSeF8/+LmSXT82KommwMxOVUfogV0t6H+6I1CnbHWny
inUJrhvDn19XwhWZPi8CMowhGbMjPZY2sv9G2TBkdF6xbtkev9N66O5dfuZy
xK/hr7IM3Zh95kEgqSaywN5bWPNiK28c0zWNwSvZcJfJqdIhc0SZ5s8v0BzD
cHrvDuduxI+OUvFDdfgYXUdk8OJEto5iCq4G8TWZ5oX9MJghUQFVKKKDVd47
6myYAOBKgF7Ory3+G02jBULrZu3Ulz6hzIm16938Pg8I6V1YsoPlSj9bDpYC
UwcRBL5xYKpHh3mnvpuZzexY4EwFVD2dS7dMsfaqw+XVEuvyPSRZupPMbXUc
WngwM6ogVeaqnJK2lNkoJeqqfLqsa1SL/8i86/sq4oDeTIuktVhiMwyUKnkM
EuEsdNdq9x+8tvqr9Gpfr/nAB4dU1Op/zTIn0GT52U4jIh/kSCrgosC5tcxU
0XxVDURfVha+fJOd3FYk9QqwO+3fsFtuITUaorQ/zh1NjjLIMXem4d4M0Qlq
cB6tjFYhz2Avix9Wzx5mrqrx+n8gueBH7wq7uQzNn6Nhu+ZNsJdNYy766+bi
uaW71tI4jnmxbrCRxz6O76il4HgyBFYGFFzjT81kh/z7TMPnD8H4SBctaJkO
+hLKbGlU/5a6PbszUa/MjMXu1fScCSI49Za2trbRyLTRszE9BTMEdcI/m5+k
oYs+bg5iMIbsu1AmBzUmScpvTPySVP3G1NXVKSdm8s1cYRTJwmsLq7d9nWBi
dtQKqaEx1zyseKCvp5OxFzhtIFw/cgBap9ryyZu3yAgzn5mbtd8OLWPt1Ach
xaALxv1E0LmP/O1UQqwfE+7uwn/eKYALqc6sQFnjEbiwN6x+qEh4A/iWZO0R
pWQjtCpljPQTkIbr9HNhXBcIJgfOtStC4I2la/0kO8Zm8gIH3GmSpl/XK9la
fG76U7noKJ9VCAYwwcjCnBzDdpqjvwJb0H9nbuFPCKOPVhxyJp5DkRFEl5CQ
rXEjgIcgsfC/LRpIU+6Rjx47u83vnx0MDu/hVjvHviNyrWFBbRzCC+lwncxX
Ma/7JbiixZ5djD/EkGzewHdmrb6VxsHvNA39EYc1CKU/qK0cgqMvLweWRtHi
kPJ7ua3UmF1aU0Yfp2YCIhXqQb+lUuMO9qt2ILpEZVV8pSOgQcfoLql45ZTb
AUSA3ZJSbh9hZZh/lW7CJehVZv6mlGdh9dIus22SdSVvsoLir5ddrZ4Yj2N2
rbmD9EN6C1YljsRqB9JxLOq7BroJkd5x1nQkyV3F7Vdu/PQ2M+6tPaRVxESf
ObSCmBrmdp8lBLTYHm8CGKU+Bz+r6aXipbWMcMoO1C4GgDNpczCwrryD85kB
Ci8jqw41vOlVMY6pA4W3JvJh7zLRH729M141g1IixSahVV43Ksv/QnJoCCES
M96M7vmqnobsM4kh+4t6WWrSlzBL4ds7ZVHW0c0CzBYH4M3MQznQ8FQD1OZ8
vHE97HbQgIRDxlJyvsHbo80yV9bYrzSL3rib9wTOSVdFORK4TW+EcwnpXUVd
7pD0jxPfJjl3EsMXa01UNyf49yc413+1lDtnJ4LbmHtXJbsvlD6nZBHxjjzu
36431nzLQhMJpEVwEJldDN2dk5OTn+qpfQC7Sbl+hRInJYVV8LYWvm0qqDUf
MYQS2KRxODbxQRWg5Gz+hUvNjSEHIju+E13gfz4908bW+8CdX2IGK5TvXjnp
7ntZla4A1Q+abMLDyDYSqpAhxciebpwIh8K/dgBngjyKS1BYNjSezWH/RAkl
FeBA2WDpb+iH9R6Dy7ew29ALnuzaL2Wg75I8KJcSvFtsMtaCmR0l2f6je6As
iOTIBpMNJZwDCZneFIZSobxfsmg1vG8QAZlw+CO4MbpRDx24FSZErwMEoZ1G
1cQvfj8egoGWtwFEh04EG2rZxA/dBUGbnmhHMUzOeRf2ze18iLIwptA8NhOf
JmEpzA/N7duqw6GpEe0kAnYYJ85ehHUl1QVS5SpP/FY9CSZiviplmAyqEwbF
ukffvXm+xzAjN9GaO0GtvskPG8F8mYvmrdpPzYVxzCapunXdnNiz4JKtJ8X9
1qkJgnSDQ1Xc+kWqsvfXk+yEvCgUx9UxBgLvHhOk/fyWWDUcKmJ0tBiTcph9
/ng13YnfHj+qpxfE0tNM/X+typv709XGjaMMMfjI15Xsxl1f0QFRXAByUGMx
TOAZ0dvUHYz8rwc+EInvAbECZQiusWcExoPP3rnEPdpqCB1jtKFhIXosUQdy
5CPywOeBUIgk9i239GEpC5YnHRiYB97oa4QCAtbiOJi+CpDfWdvfu03a8vfS
rrJItu1vhMW0kcS61IIXAIJjD58osfVEeEw51dN+NQwo/hHeOPIqzeJY6Ffr
Y+r+kKTJ+88YtLYZjLs9h6T3drQBe3GxF6BuRx/iDuJq6x5fY8sOQKr6Y7eO
PGJGqGcgTmNBiNiy/H/OFX3UOqQ9i1Iu32liIDVEo0IwOBuHGcnYcSPdPX7m
8u03FVqwqK5Xpgaw3nIy3Icu2mfCz9dfI/YLXDs5Q+dq80VmX+qP0tlW59Kd
bEr4p/KOHs2o1axPVmJM4cnZ0dqDwp2HoJ75p+Kg5EsknwZP+kScvlqwN+gJ
l/R5twwMIhxew7vtHIFOrMXpmXgz3cg4Buw7KXq8bQ4nalJZHvVo0Yc4uhYL
OPXIYP2HfpA91yy+ZmomNIrkRR/F3ugTx+QW/1lQ/GyUQaxpJdmx0dS2RF4f
9kY75Y/IpePLjEKojKOSoTsiqKwMPOzn0w94yXpQEFrKj/tHIkKIRq/0qr5w
rHvyhXqckUI6U9EybmOK1XeGqPNgup0ZhMQkwGza5ZWLTZnYLBLgMII79Ibj
ePZYEAZCBMhnsyOyDDybs7YpzS84eNa19cQU2N6w0wKB8pZ7MIWFA43w2MfP
Q2HCrICGtRcT8wYEGHY5Gz4qe8BCUu2pJOjmufTD+ZgDpZFiH8AtfF+nXbss
UBWk5LyntLwa+ecRwf8baLmOvC0ujyQHo/9mPntvZQWS2XspBd3cxDWB+v6Y
6GtyFf4gTUAmR4HNNq4fcwGWFHv5MhGhuHK26pgs1WqP3KvgHL+feHSam7vn
PcEExGigrz9fW9C+neOJ901Z+a4xZkVfSADebFQzTIH196pppVK78qqviV6N
5gzDARru6ITUYMvNpB+xgKbFk9RESbszF4Q8jZSXbvnjjZIjUVYs2bI/fDqD
ItBs7WA9kjNf9q7uSOTOyzwt2t5Xhs15xX8IW6CtGdw1oyReYfhcx9iee8Ji
WKVn7V9JYZNNQR4qmlCW+pVh64DCNYDko/Tv8uYqLNXSX9szqcQ+oF4hpQs3
5Va7E+Tl+mnCnOh0X6Bsx+adkjgP4oY4jbs+j4qbIJ3Z+DnoLmfl4EUcO0nv
J5lNRMsgd3XmeDJ3dN5vOpbT+Ob8pr8KKRjhGxOTXFxGcKPPiOPSGL2QRBAV
SdJsZLpOZwXfgRYjdahyd6SfuP/N02zN07A70l3IVpcSHk5ec1kof5r8yXWt
vB1/i8kbbk/twmOrnNdO2fRcxIPxq68tu0Rrs99opmAQlLJkd8Oc+6qFHjev
IzFjPizfWOSv6e8ZmSe9KSqa8AsUxDqLGR21a5EZf0C+rjCTRrenOajP6aai
tCiWtyZ7v6H2pWr0ApEWtF0z/Muj/oSVqNmPDL6V8kpN+AwBv1A6BJhrPVa5
V7tu9WhBpg/u4DwQvKTVhhcen2B7kFtjw14LtAJiQ0Zydk/9pNgLjhnZbx1o
/ab4JOZRyqz8xppFplYTcuU3a5Fvf3b9r7M2atNOjyUjAKuE0g5PCEyxS8Wv
uDOe5FTcmYxD0NDbHhcUXERQtv+4pOoFdIUBtRBjeVKq2mKEaEFV+Z+ZkxjV
ZGvz9N/OjmO2KUCSDFWgdLTTbOLXXd4/qs1E9/FcfYJE0pF/CnoevNCAVQt4
WgjLIIB6FaZPMt3JRmTGpt2Ry2bJzYa52XNaqFq+0f2/uYamO+sTr/ZdIiDy
/sU8VIbW5ZLB/XQhg8hKXYw6EfmLsFR2KXq7PxeVHj4ZVgCkCE6Q/CdCb/L3
N9+SRzf0hOFNQgWsCJWDd3trBYoq0Lq3N4vO65aOh2lnsW0f5f2btFSm6HNW
b2OqbKczL1EQ9F75IMFur3gzu6czNuMwAgQGaado7fODyCZw0OSq3KZHPFpu
EkF326WCrg3joY/KxoNf/gKktb10SmvreG/ZWcUv6rihhxJumjWk1s9P3vtb
lx9lYewJHQ6T0pmrTp5GpRkcUarnWLxijSeO4oyTVljzZ3lv7pm7sYBw1wkJ
LhfSHGv76JMOTqv9BC1OvrdutpPfAOE4/EeW2dR1wss5boRzD49751HdF/GN
K48/iNHVp/AM4TKqFvqRqXTNtgytYAoxQjYLYimheExAUQCO1tgXWbkXPiMU
ZCvPbDgWSnoI9zMbXRMZHgXdXWT2YD/o28wEwRvRIFjMpKnzn8eNCxrRNVTa
hbJ2WMsx9wMaPQHt8Rtk2P/wLYScZ85Rg8f8uduT41qne/qyOaJp5aLId4qG
LrEfvKz45ZVrtSaCYQ75Q+P7Op/+rRZT41bEx1G/new7Z0LRsV0k9GUJQ5Qk
O3gOYaOCEIHiYDzzdXoaQ7lzP90+57BYJGaqJ4JjObRSdjDoenjmpwNLtcyC
JDUaoaJSZhZXVbfjZ30+2H+utGxRu+I/AhqkbWrGDBuyL8UMgwLeUV21XPsL
2MbdqMcgFmKO7UFSepFsZWiij9p4vlzBS/0i3dJ0csy+jIB+OuXsln/lwWbq
VsUHD4fo6FprqcqlEaWp0YaWbXkwWaVV7JvBqHKlhk1vHw+2esL4iL/N8lYJ
dPo7zZXPHfA0bF60X9VkhCRIXWOGggOh0Z43nGvwvf4PmG2CYqI22vsA/5WZ
YRZhGocc0wpABp2AP3i3yjTLFcpgf0tStGMkAha+pf5z5jzLlJ1ArjBMYm7m
1dGCovwM9ArawcR3i7K54gJdfslApJb1NNloe7rWBM7qKIOEvn2vqDPaAjV2
YDYe1T+L4d3QF6neoXYG1ncp1uoFKQBBm3SKjTd24XA6Su3f7RUWuNyPFGSt
haddArdPd9M8B/q+6SfEd8YeOludtq20EiyFF2harR5jbeshbm0lUYYmNXHd
q+xvGwLwQBt1UdHVfzOVc8eg8LXAUXmoGFmYGLJuk3NxG9o4qDI7UD1IsBZr
+Zw+IbOeRXwAs+8vpZcNLP6yD8VrsC9lYdwuthJJVOMNMcgukm4CjSTALM4B
wOaNadhMPXMACLmbSaqcphcGV3cKXtCdvCIFv8udnowSmarOg/a6tPhqDL1B
aF+nPgxlSypbt0fsjy+C11z2pjgvu/zPtKK8np9APbfNpBGUWhWBmbk2oALM
WnOqmiJSki5tzFdv1y0P+On8q5oe1yS77WlInIH6BbsOTkZb6gkOwnRiRvKn
ZP5WkeOuBWxbfYv8hs9QLd3desp0Q0hibskDl2Xjvti474ESV9GLRdB4jre2
d8vzT1eF/5qEh55Pnr4JZAxKusg0PftGrmrJolyrPA6wWUtCmXgVDCNVRZ1k
T5+NTvT/YCSA2VY9w5dQinV5288BN7x3O3rozVPDUTSTS0H/Sh9uxxv1CpnO
uCcGM3hIQhaGUAitkd+uoEevRwfOZGrFt6MLdMT94tIAwZoeOO4LkTy7iIhY
sp6MKE7Dlnsgm22qNT4H0Cui521p3KAnwjz13Ph6IGLaA5hASzULRBN7M0sa
+j0ZG7NQMJevXtmzHjILaeBs68rXJie6ME4b9kpS2QxkLNht/e0wxuRlBH1Q
euu7/KLAGyDj2vYAq4MdQSuK38vRGfy+R+cT1g9BIpBEB6okDiW5h5y5BQNB
ACK/0KzpT906WKEuqE9MdPEVXZSlbEvtyIDhFgfTTP64+DkiO6mrQI5DHPF7
lf4cM9yWwVi/R/EAmLCu6TT7PIbeBpMgXrwPikBfzaieuPKu4PHEgtDwlDi2
pGtIop5WqdcAu11ORt+Oxk9Q0/p5OtFHlUKulPndW3HZ6JzSE3XmjwH43+dZ
noferQYOluwKU4Y4sWY6BSvAX6rmZctJ1CIccgUJKeU2WYXslEOBaGHimr0R
vldEfYUitKK3nliCYXpFSiQvo0Ch2ch7kKbsrc0bS7yLIHanYlC3DCj5oa8X
qX6M3GESznPZjqiHE/RGdy9LLQYCHa3t54kHyX9vjROBO8zZeNyuL4xrPTYs
IAajuv2M3gnsXKrvpGNDOICSKaJZNHL5h4g4XWYVtyGW6/516pk1+XLmoSc4
Gdsj1u2lA3PzmEbu+GnsFyScXt3FEi/bsTc9WsfRQuC1kIux1mWrX9upHWc5
7jrQ+FR7VT5oFw8gEtN1k4LcuFH/Q1rSnB/yAT2fTISix1htfqHKFxQHVCEn
xjFvm3GO/OmmKNiIIwInKB4CF+yoNHztubKHIPL0xqLYzzTJZweMAR/XEiro
b1sVQyOL5X+6jjJX2NFcL9w0DS8EXSP8H2dUavQ9aQSj2/STxqHj+bI3NmcJ
PPxH9tzDUE7ng7keLso205/P31o5mROQkLE2fqNd8hm3MG1OQTxwgFH/S/oa
j34TlspkjYtpV3USa4fToPkrEv5tWsSdVGJyXZDLJy7aGQitqj20CMIqNH4A
+HRxM8vMddXnaS82SZ+7uIRqPZdO22sEm/12SkrHy5bN8QOtSs98Wd5IgcMh
3PBp+ZqJOkCBGrfqiaiyGbx2jARqqZmRdCVLpnKVdBHjzsMPR16ej3e3wxxh
FfJr9CSS1ewjr2dYLK/nvHHKpD+z3fCtvPUZqpNNV36sTVeEmwoNrSPm9QLd
ca1bpWqcNWs8jd+dNjHBKcodfkvy0Dxh2yX+uvuyihEhF/lvYIWbd73l9S1Z
qbvxqa0yinhP7JYo+PIRBt3LEfagjIDVoZlRXBf2TxD84+X11WO8yDN8dqx4
cEPwpp0TNRY5ID8vkRz0E0zxZxRFqxani7USr5Lg0MhUHFrNBW2OxaGlUSq9
yoneIFNqN3ltJmUqEJtXLxqmDi6Y07CWI/Ql1hoDkigVvOtHrT4R4ZxPD37a
YSesZ2PseoIr5ccrY0uGS6PokMVIh9ASeiTBi/I3iA4zPyEDOI4lT+/91ICG
AeeyCFlQIKiMAtBcHErnx1Fj8gf81F+lIAmVMDjoYNkmgAcSUPcI75V8lsBL
RUvQ06NDDfxMfmylQFJYMHTdofGK9w6SC/rRi8c1gIlQv4wX/rjxMqwKmEqF
b9b51fitCu+IdsZskrzy3yeoAojMNpV8Sw4kqJYzmG8hWFr2Fu5lFfHtNVAP
W0NlPMetbGJDR+CKEdDeEYs1NYUXXDDFCzEzOVPb/M0HszTTlK2TttaJrG7P
btYrhKOOtsAwIsmz2XkU2TI7wucyCkJmqOfN3JdGlGstdBzM7Rq0FKwDc7Ts
4IFs2+OZxux5mos4mTKUKPkrngo/3N2EQX1r8+fIazm1NJ4tyCMP1BKI9e4A
9HZLTNuer5ykg8GnaxgpUO1OIjs0gnxr3Pb0KLX1QKQoux1c6fV+3/+7LF5v
RyutGiIacZBL5Jw/VZt8aiLDfMsP10f2SX0AKPgs5OhrRy8kcuQRNjnGb069
hk4KIBXbli51ye0Xki64mhuD4gasMhU/59y/Kz/CaJ8xGpeEQgaJL+iPtK61
e3YFLLp1TPa8XJdfgTT/IuF3V7Cn6wCY1dXispNVunFmsp7lnYFtc8ieM4nV
vG+hbmwoHD4zc2wMM/AC7iHl2wonFyLPYr09TFblXAZuOiVVHGtnc0mGx+0b
KMGibNBp/1M6Ntl+WHti8gpeIpG3PE4njx5JlUWvNhkrMvTI59su++S+feAW
MRXJ9ABFez/ZsHCNkbDm4dMkwwQy4A61DluiN6iu9H2CgqAnQ/nSgGcMbgsZ
s3Rjrf5mTtL9FfO2xsTqzalV4Yj+2w33Xml880Bzme7HHynH34mhg5EOkxIy
xY+YGjVK2wjDC8dQwdpoMHp2rJlnsXiQbny1EqCVixgxhvvGPJi39OdqubjN
kY7IjrtWFHSRfPBJ3BSfFR37oSFOfVpgNOo5axiHpCFlGi9l+nM0E3hqPDpg
a9Zbh63KzBvtZ+R1AFBih9WK9GY9Dc97ESliZZqFnIk0rLtWB4WhsPz5gN9z
lF+DG8/E+4Cmw0nRuNUu9d4jT+v8NVO4BtS6r7i735zGiCYTwZRHVxqtRaOb
TyP28OM/W2vv+kTIZT7/BNqeOTjK3wOX/qDVhIOJ8c9st5MC3jsw4IvW5J5t
plCBpusEURbRtCQM3vQCHZzUV0hMGhj/LJXtEtufi1Re8FgET6hUc/bbFrjN
+nIftgMbNRdD7iPpz6XzbTQwh+8/9ZRY9dqo5aFtVJHYgLKIhT3qgvn1NLNZ
iLs8I8NZ4Im8dphbLRhVbdZ4YGUQWxA6ludBve7uANhZreU0YucrHIKeibsE
ZO4pBC/6Tjys7G9Hz+lsHo2EYEKPOHzK/UMo/rLi9NnoXabS4spnIdm2laWk
tVwuIMV6ZQbDbtblbQbK71/c8gIioI/g0TeHmIGnUsVG+4XK8jnTtoQ4ykxZ
qxCENYAVdF868MrWKsW0o5NwlFAZKxuh8emdc4sACLI1/notxeBK2Vb/vILQ
FPLob2/OmsHJH/Aqp27QWQoObE6FD8XxSSzC0IFyHRfd5mYebKCCz5qmkUgm
kc7xqsosIEzab/1H+cpeYsHJQ7a+7bH8ox9dpS7rVyXi7QitaAqjksxEcbUX
RFpYWHeJ/Vc/5CAYivNcyp6rnEuZPC2bvOvU5d9t/+o9b3d50e1gFSbVX/Qg
YW1Sh3inww2WhpeMMOZI+M476+Og3kmegj6dnm12YOt7eO0c+eUhgAtUTpwF
kQGYHsJZiBpMJXyN4lij1u047yhdEFOeTD+bIiBM4Q4LQmI7aSQ1UETDSfz5
3kNtOM103lLFW9k2R8FCEYQGV59MiXgZK6AKgX17LUtyIONhWihK+DB+xlzw
XGUyuijalSfXFPwyEPnlaikxJ5YmCeHdb+gurTN6+N8PX41HyB61T8mMvLgW
A8AdJFkUn2qYpmL0plw7pk8PoeikYQx8vk6ZeqtAlx4AK0gqfxFrC+ECdCo8
Vyz1BLFxlblS42o/t9E/KmX1NXEKE5Yeva9ziltdlzshzpC9QGFmayYQ8Vxf
3UckIAhJ/wwyreVFbb1+ad7+t7O2qbogIhN/5UFjp/sxprdvkpzXNjUscAlH
ZFQWwREQXPc//Wm8fV9SPEg05RUF6mSjmNHkM4OQzPq9O4J2AEF9byp4NLtW
Cxmtlbi+MYr6lR3S9jx3ZS6JUZqESSVNMWOpMrQopOJ3RmxvKSAG9LnGk6HP
0EjN33UwDKqOfCsgDcrBLif1jZVimyNyX+mMryigpdkV2aiwHl9jwRC6TQkv
YR8+xiTKUoJpVgkr/O5ywRatQafEEI+aSllTQNW+T21coAfSV8ovK6geymhb
AzZLGkczI2t3he73sBBSZvCRnYigd7P5qg9UPh+WtvzS759aCntZ1dsDD5RC
FSbmdW+TeJckc+lAwSrvZXnBAdhz55x0XPMWTPkEll9zdyKoFcxXJEUaZV+Y
7HTMUubTofDnLORUhI5VhNQKrnyXlsXujfHVlKb/o5vtEFtoAHWJSxJykbSR
UAT2BTH1B+1iwLAJ+ZC4+AcN7Os9sQvWjZi5jMkt3cBc6Cb3J2kPTTIGaCwu
YuNHHv10TavNdIyj4qjlhpWpVvT3Ed6GUJIJlvLiG7sldohMfJ0yLvxRcbp7
I1qoqnPSVfxAm7afWCHwCEUEWdbh9+Eg3k6R7qK1Ea6V+0bZDZkD86esbzXr
Yk4svCN8RxdG7HSnrJjj8lt2Hh94a5wcYfy39hXzeuGWmui35YnwXWz7hTXE
dTX+xZPCZxCaXrf2+pJ5UChaGApNuLO54kJIQ+F/niaSZJN+oPafS+U96h0K
5oybeZPD9jOCIDFsLhmj/zm/zsMZhIaSQxZCHWOxLT5ZikKDXkepEsJ4sKXX
jhi6XdEMRcDG3/zYCX9AG2PbxnkqtTHCPU8vEUvLo37d/vEnABkH1qbGQ91Z
EsVgPujdQU8Sv58DgAjKdPV4FGdKpuasu5ljYrFOLnq3x5cMs+GOTsIHE1qA
DMGNyjf49TSGscpIhZGMl8aPR9WwLbs31bRJMk/ivDJiRx9bVbxBcljlm1Ni
hwUppE7kkbOu+Epik+L2Lvv9LdE7//FBw2oMUZgq0u3xoYBEMMR4vKPgk9PR
a0e/CTc5NWAf3hYljkrDwiwQ9vgEenDTUtyus8qdya2IqCPe90BvX+ap+phj
+UMqsJFMjpqFKUM2No8aDmfzuE/AkiVz8V4LWKMDod2MTjMpaddD+Xncii4w
H42K4yy2Ejx+8OcUiKYyq7uK9bwK3UB+JEq4Ao7AddP4td/DP4wvI4avfa5W
YiW/YSqZXCN5RoausiNOiMs5pb30FXHqcR+vMdpR+S7rUoFTd2q0SWTdBjrD
7AUkhE9ND8WdMqlRYmYbmH62tREKrG7ZijOFdDdqJtgndWj2sfK/uWdL4NMQ
qSiTQEur8ShRAwpDaPZ6xPmhPuNlWg6V62VHpLb7d2L0s7VPh5IXv3TtDt6y
/ed0K3S3Xmn0QzsFh77qhtx10kpv/dSct4T6FmoPNYRtajRlKMq5iUeLf0fY
EizxOUzt5Xz/l15t5WsFqV1GfSI9HlqGg+SYp1jBeFWAgSKYgTA2OwMuGdut
MR04HjG6yHrqojWYgVH6gnj+6py9DpohBdq3LDRhfPKwLdnvNvsZC1vp1qZN
kJMh/mAKQwswpSeFNWL71WemmEyvAVGcyxX7j27ouSobNCjYT+KZk1hmi2rp
ViNbp2a2wsj8voAf6dt4KK5ES1ioSBtZ2CXbnO7FzvvMvS9z6HkFQ56Iop3m
Cjfs1A16EqOWLfE5huvqngXjMSuSByIS54lCWaTIk/1KvNLVDBH08E+xmrYw
d1ubCmXxmdzfYjypIiefAs/fKAiWa5ausuQm2/4NviCs6L3F0a8vjCmZFuOq
D70VptG8Tk5D25YkK1Rirme1i0YDtHJjjplHlWH3GVaNKkz67kd3kdCHLNOx
oR8GxfhB2ep8hcknIfWcayszj0Niw5+jxmc5WKQpUjurcIHcmdneHjwTxO6K
Az+fJf1p00am8gnYOAt9DNJb3W4PxrGkhhbypOJX6Qi9q53Ruouz0mo9sxTo
ezTtKsfGNo3lVX/u0m2pL3lOnU+HO96GOMEb5RFvRVtPnAK0+80f+dmsReGH
ApSww3baCh5iY/PvhlQ3/GbxNudHEFYP0P8TL2hc1cHQK25nKheauqBLJh5d
L3gaXb0sXjO2QP9mz650KFSji2VnnauOAB+q6J22CyCV6zhdTWEm00xhTBCO
k0lFUyj0EEA2kgZxW7gJAXgI7MCxmOqRnsWCzRyoerB6g1Wc87IZgyTVR6+v
k38Rfo8PCADQE/Yv23MztF03q9H1/ZhWhPIQYbFZeJSWymcc6rPggH7YQC6t
MgTINwf7G2BUeV+8w1A6dhjk+Vxr4e+ZYsmVwVJTbp6yWskPOGfXJgm8w8Ds
WlNjEVssL31jcPcOocJZdNMZxTXWP94A40L3F3ZPZpWzQK1XROEPvL1wZIvh
hFVSH8frmb+90+kkMY9ZmsYTeSbnCembUkRKKeUdNoxjiw1Oz84qEFBwpUZY
dUhIleF9IlMbavebKptm3qaa1J/JHL+oU0t4DWOAl0DlCGZ7ZfF3js8ySFRG
YQybDFayw0Ao5Xv0LS7MepQG6aTA+QU3zBIUyrpQ+k3cNS3D0a+LyMWqdcFZ
J5zC/gonmKvzX1TBj02uIdg9+jwEyeoeSkz5NdsI2UtYyw5ROMVy9PyUkRod
MUtPUorCSSecK+WBVZhgg+SxXlWnARQm46cssmxzS7TJ5qmIBKizeRlu81h/
vQaBqaLhkd8QMbocUXu90ZB0e6q9JPLs+ndc7D0w8rh4KQbWSnD5I6azcuz4
7sQVkH97iqW0u6vWCwQEQYVl8eD+04fqOddl4NxcTprIrMM14+YPCjc1PJCC
+jU3635iDW3G6fpDVkBurY1sdVbOVySSHJMsiq0O83KaLuq2MyqDs22rc9Sq
oWRK3ji0nUybAlcL16Ah60rkjjxFsFpQC8nvHoxvfthYDu6TxypH1fZtGwiF
rHVNaAaegL1mOl9+644X4HdiiD1cqnZ3Z0NulMLtU+Eeo2c7p3zuksjDhtzI
/JIzt5x3cBXlTzHPTX99Easoxu/uBD45dizefLpzO4YqoOTRf9yLDsra32Mx
NckTLI8taMH7eVp2BjPfoHuchcXeMuulPrMDwOu4tz6etlre8+bOe1Tcd20a
ZZN+h5r/y4yVQxTpIJ+Pl9L8QS5elzvny/UpiDbq9fS6UPRT++bSrJMTAyNU
s5E6SjQxKOLGZnbeF8ts+9vF5Vgsb45gCCIDS5/t5i9fep40NGtpTL7r7zFY
ds1KFtqwrjOOyhB5dQUysrFIDcy882mfDwYy2cdsM2TivBPLL0DMCjVtw3qF
yM92NAHSmAZ+iQvg3DvCkZgmkqK3Vjo4TKB1XS0P69kh6FBjQZi522gUJnGA
Hz0dVob/ju87XFi07a5uiV8wEV0Uxrd6QufZMqjxKhhM2I9H6vc4bFApNXx9
viDEF4WSFmrQZnjT9Rb3Df6wBu6c6yzMQcioEVW9uRy2a3unhh51LH3rhUvi
zMfHUprLs9GSP2dYRDhBdpr893TTz2ETCVJPJn224QDDYp93ueZrOMHz8Zz8
R/mAbEQDGhb4iiUL1xklJBZiz8qkMuV+qkduLtgg6Ot4yyxEWNm/Lgne132z
D/iJ7D3Fk7IVBgKxA2/KOOIVQxGEezZuK4aNdlhet61RZ+R0vYo6hnszU46J
G3+xIgHpz4x7ysfqdG4Mhh5HcVkzM1Eg6ZYzOQgS/LFd7sDG+Kg0bFCp322I
dHa/YedlY+RNxb6TsBvlvd5Z1D6EzW/G3lPMUTkeBffCJI6Alb9B62U4JAlN
JvALiAIbm2MmiZoXUCb0qDGTUwenML/C8XEYrFwW9mdXdpdSX23gCvy9mPR1
pNcAbHJHcrlHr0rO6navUiLeqPRS8oBwqZEIBY9tqC/YJrdx7kt4S5vZEidN
ErWW7oc/nB6PTONCZAPd99vgpf+ft9oEtAYhCLWHFEC3Dqdk8EX+Sq6KbO3E
ffuZNkYF9LMHXoRYfMQnYkuY3ehguPj8s4nF5BAMtuY33kieWUVhm37dLvbG
ZJDPxFW+RR+fh9QuEb9Aa8efSaPorsYbi//Bo9j4cdCS3ZbciIS5rznVQgSK
FivqixO2aSgib8bkafF4FKCbyDi5KCx6cViPjTGERXI81kU37qq7T7veIAeB
NuUtRaO8um480xjM0rzZ61e5xKs3N2oRwhAci71M2nkhldIyNLRhFmJqo92U
5kpXsLYuSAh4M/e5WdxNztjx30Sd5k7EvAmz79E84yf6ZQS/skb7MaRJCout
UkhU/xCxZP/fYvX/qWgQdLCGmzhMiqqRR8CPmPTKyZdaCyrY3BTX3k0U140/
dmOq/H8YwZPx9dxNPxJ3dwGD7bMRBhQ2a50pCpwfL/My1fHa89llDNwVmUom
idoEF51xRefBU1CA7DzZOK50tfPkdcGxelvBzeggpNzF2ABmFqBeQ31edpzL
TZLF7LE6A8Y9Xo1Odz+ZDbbf17ryKxKpZ55RVRozcAqlLNoJFqh2MYgWPZTd
PAaGOKgZPMak6b9wsRyKxJuQ+6UKa9vPlG6H+MdnAsRmzhy+4jSlEFoaYl9c
0hPMYpjyknQNkxXMd4xes2FOqrYwAWFAtbrw1+Uap9Ororuyi+0OPmHQ17li
laBoj2cNsoOlukHlDKEweEvDT3C/faQ8PTPDckwmXHoD2vZwlPgd+spuiKzj
G14i3M84F9NhY6/MFh+ydB+I4t4HH5rYtDFEPvdpli4Gmx9TO7y7uR1fs74W
rCm2LH7hzwhCl8bUVlXRZzOhsFi0BPqXEn7rezP39EyEWELPcFSoXP1mSLEU
xMY6CtxHX2Vciq8NLdZMvCynV0fEPl+Jlxzc81xD3n8FypL77c9BKdhz40T1
40s2/dZf3mkA1OVGMVzLoRb6t9J+bAKfi91YFXa2LlJeE2WAg1L0/UofDST8
l+OGJqwmG5J4bfGoTrOA+uBipRtIR+UEalJTaKbaxN4qNXOqzWIg5OS4bH5M
l8z1ihHFR0le3bBDf6vLBqdrZqiR3uMeubQADGIiQg1wTWZWJi8eDpXMP7Qb
cRd2C2ue6fsbgISnxcDqLhSMDgc76imyWg9Trti3CJleA4cDfdemwjIVCXAc
rmttMynYW8CEhO7uj5H3zSBRQwtbSZvxvtmyfCODi0LpT3ik+d5QBafR+cgE
SJEjNLJhtGfH39L5dPBYPEjR+CpZ/auh1k+vUIz/Xr1CC6LpwuQ3w8MN5+f6
aq4NGJYM6HVsg9PdVEfPibLWH8/gv7BxVh5Xu9Ljyv7JWWtdn3oE4uAXYykI
ENJhXlSf4nijKgAaEPcLw3fDMqffleNJ4tqgMygZvRATuDSL1BIgwN7qzlMK
7b3vpD72QNfkhWD4dt9YFcnQaFf8dzjwugiJD9zLGDY60DZEHRhj5LynDMQM
Dpuj/0YjmshjDIXSRrp2NiiL2h3/7YakJbaGh18893SM/B8CWQyzBXKHVOTy
uf/lQHJZAs1osYe6zP3Q4Cxm6EmmCYsEhncDVgrcsx7RIW7zUtJcZPGQf8pn
EgexzFpLlkhkrlv5K2u1heIJxbhJAaapagNwJev5J8W9/H9h/0goQhC8Oaqg
MrGA9LuTrTLhPUPMfRELiIth9BGMO8Ldk1wCyOiCtCZS+RCN2795DNzePYdZ
o12NrR2Tf8ua9T+fO6CJ8Xfo0WlAHAtwZUgpiKIM8UeY6jwipwADSODJKXWV
oWBLTOCiasxRwS1mbf52NVmCtjqWB6275S+z2LzkBiPxSLhRPKHF8hKUUL0q
DQY0KagcMlxKjfdugreTAWVb6LS0YNPtOipm8JirL3+gPSJu+eLbA6YgscQt
+KwX1IfTXt6YwidKAIOnALB+KQSoyah6tkEhudfbCGyqtXPaIvd4CBrtj97F
Hp3sn0ZxhpaIQ5fbTI2kequ2pM8W4Jk61hgw4c0PIVz3gngAotHiIbhROylr
SGAs+aynQcG8B4ZMVDs1YaNtmVlSkv0P9b6DfysiAJxGybAhPmzhQmDy+Qdz
lAuEatj9qSJBYY7hUFHlSY3TIqkFuX4tvqbi9z0fHNK5eg42hkmdPKBPeciH
o6b8rKtto0zV0hHgtP41Ammr2l/vUDmcgGfhpUvI8oRlIi0oj+SgH/ViV7Gf
yQNN0MWU24/BXOzjYYpwiBrH6Q+WKiJK+VhQyQRAZc6Mw75UUJ+rma+QJdLD
0pUhAv8fsq5b2cdiHHmxRW9czkv8eultxhum2CMV/cfrHmXw6oYJh+OzuV+k
oLI7QS8l+7Mby1g/S1X74qTkzN4C3qyY856YRBpMr4ooIMlRkSwkqZn/2mme
oxt6fzY/sW71d/fp5+yI7M60ykhifOe3ti7xmdq4kSKAoPiUikTOlrTOvsQL
SEDdX9GlxDeRk7CXPnnETBqWeEgbQHX7OwrpV0oNVuA+XvvXbVoRgs5/A7mj
R44Jzx3kcuwcOGMoAgc4OBx4Aeqhc/l0+DIQscgjJHfOU43nSEZ6Y+/63pK6
l8S8hVsv3zEcMI4xpIyvI2jHXMEA6xpbH0bN7YS/6/FgSIqnnN8ErgOGYXGv
kOGnmVnpWjzKWWa4YEoiNNiNjUvxKMvZ4/3SMaUFDFZkxDODf7BhXEAqvkPb
+tHLZtAn/I70kgZDU2T0ZgEaJ1UAkoApk+vjZ9cBMgROhb0IlmAcogdRM9JQ
onDCjIlpqKsYxyYdz7qcbRiZ+2W22vDkwdQifSgoo1dMjekKilyl2VmVHVH2
qXvDI7iQTfQs4SLT/wAuv13epJbJ3R70ds8yNCZcHj2hggAkOWge2vhVKX1Q
eVVj97KrExNJJiHTPa02jUieOomzLT4m5a76ZPmgMmmksKDjY9rC/Gt+Y6uU
PAqIxxqTwQHnpbiHeiiXMljpSXcKCL5uLJBoIfMmbRmtNXyE5S2h/P9BrZCM
k3h4DDfOccy9y+ozr7Rq1Y7lKS5o76rnZCsXUPUMI3Ti1VXv5XbfWri4nlA5
u4v4222EbOqI4lajfZMLBfPeADDQXfj6TzKkpChyy9btaum3fAWg6qEfEPVH
TyeHJHFz2Daz1a8j+v3QVXFCmG/JNdbv1WoXzRzwZIC/EuXBb/6FPwF3S7Rc
ZlZDsFVcZVIZY1QDWSG8GZCZhE/35lpyJPtml6u8Rx25zvK1fPagZACDFy/n
gAqM/8yL9pYnVcOSEWNQ5LaMgvcYLa24PIFy42Vb3dIOwFA3lra/lIeamL58
h/H/MCh/BsTCpQH/Z9z8MZQau1XnzL7BJDC+etRvj4si0ALps8hief6Q+kJU
tCtrmJo1VeTQTr2eYSGWnSDsAAE+FdVauL9rzDrHTb9YQ2/qr64AYBWXCXAN
ErbtpMfR4sU7oZW/HG5C5T7UJ8Vs6j6i/TZihUKnNC2CQpQQ28DfpXMSypAU
/Vc2jCVx0x/P06QVxYY4h6Pyet0AYrRd9pnm6jdBLOlZ7ONfEj3NLVK1WYFh
eT9cE5cZDLZThFFkXACHxzqYPnezYo3oTvH+ZljRILNbtSSLlt+ro0JUQoxJ
eQNdwc387FZsuMjbGVsskTb9u+0nLIjiEsFQH2iPsQlEzorZzqHTkia8B74T
1VZVegedwDcr4JjbGaYVkJX+jCznMAizXY0yPW1nO8zEZIBmiCq0ShfTHm4u
zU9XMRV+PWN6KnhKcx/DfpSlIAOJiQchC1qul7Il0w0CbpWxpclDZCcLlyKC
9vXlBMriAZsyx6dI/r1cfmMOyirVEdA6CWESetOFcu7wdtIXs/F1Tlk1t70S
//oMH7YjEl/aCnEOtoUH36Wl/xe8hrgaQVnZNYHIKo5xAMeF91Jr/BVC/Yfp
fT63+41dO381TrBWu8+yr8mB1n7B3VCvgXcxB8yS1dRqCDjdZWS+tdnQFSiO
rK0Be6S/22pJ/wlGqxBQTfa6qoJw682p3NV2fSb6Il0j1q/QAv4YabbsIW+g
foQ2xqwG0M2KBITXDyL/JhW+E0sLKO67/uLh8BrAp43M6biQHsDK3bFsXBA1
rkeHRWOctWo/9p3Y/4GO4GQpDiC0Rwuc0asUCsMpLWJokBuv7w2b+7zQGsMN
E5F4Qh+rO5GO5Y3PXCdqSo17V1xAO2KwyOzh9UsDkp3E0AyptENNbZXno6vF
YkRMvOKbS30nXYpq4fVGPt6g/vbKiENk0ZnM/ASAZh7kdD69jrnCCplgGAxp
Jcr26JEatEk0IkakKNuBUoMCT8By7VjupeBmQFoqBIJ82ImHJynYn4X4bt2R
lOVEbgNf4TlkR9gnd/M7pozdYXVlruMSTAaeuErJwctKrCflI0dglsPStI2j
QT3HFlKMgM1yRJ9aIWm0zSCH/dpoHP5jHgxCHZXoSd+di6GsLm6xM84+vJh8
cu6g0kTFoPB5Po/vM/3E1ilmiLpJXddMgS5sLRiFC1PZPOF0f6y7MQ3OCZ49
mqv7esPD7h6mlcyaVzjXY4rTDWhMttyQcoZjhSdUUdAlNIF1O69ebRRbB51y
sO1hC9Zib6zz+MLxgqOLqKg2Zputs19a5qvRjeLOqZU73qsKOOU8fCAhggYD
6rB3DTkUHUvB5TrmZ3x6txPMrCj6gylZNZpqrxoHuVFg9szI11flbYrSbCaM
uZFuP7PDOOa9JFQX2kxiji/ssFjsFJUSWfYQwapMIN2OL1R4yvSruJdAovwR
JtKn5br1TWult3Lu4JwQ/Hr870USnxLcabi2MsEqexgNq5As0454WT8SFNLZ
VpkVT0uF3ph5G8ecUa6gaWGM9bF/Fp6tdivawtMNA+iWh7wJD0QKcncZYa9S
Q+QTRVxakliK0rF4myDsMLX6j4aDijcfZrM4TQip1jDJPF75MtYqN1SSZFjM
Ardch+eFuy+JQ3e8K6XCFP8xyHhrqIFLT04myolCDdnc1zpWd6Z9nTqkTChC
sGuGTo73aJ4CYrL3aO6kL9btvMgNKHleRsFlUiN5P17TC4jiU7tYs9mR2vIe
oFvPNSsWQgLu7pzF/FlQsxI69nJX4ZdmZPjn0PrKqWESJnLT/ojkALJh4q7y
cMAnc4U6BHtITo7q/S37JbIc8U2xEjZSnyWdIlOS7RfLMp1lXh36aVbisxdE
P0DGouVbo6av0hGHxpj5KUq0RUMuf6EnEQZ6OVmNvamPX/Fv98ViA5eyiG3l
Fk7SkwDFuLaMDc3xzJl4UZGCd424CgTB7WSWGvnxRSveIJvBDfm9iItveZ9m
BIs1rlOrfhfuKNueJPVNkff3OdmtiJqexirXv+q1s2w8zGT8oBVpJ5m0/0rw
ASxKR+TF6LuK0rutgmgv7iuKmwlBtswaCqu5LtZ9WM6SPk3DTKJz4ejIwIhZ
eOXOCznoqzcx1J/sqMgcxT7dioDbJV8Uzabd3kmqvHQ+sZ5YS//7+k46zS65
uwIrWxsQiG3d31WLM9i+S/g8Lk4OXV/+UFtNtfOSzb+B+70uJMG33yroQtQ4
H0/zcSLrDJwwBrBJ3yyT2rq24eWXZDD6SQkzLn3sAiYrSF7p8XoWXroWhX/x
1zZU43Ma2RUvbJ8ykKRPbzfZtPdnkaSfVIquStgo++eTzWrUoXyboHa5LbR2
Jwcl3e1QFgxdk9zldf56A4vCnJNyDsn1Akd2WutdlCwizunMGgys/+34303I
ua18EvFX/lRpepVizSU2Ul17yX5tUaAzFIimMvnhVuf7zHjAXFr8qnw/kzOs
LNMVnmhqPgucApXhXdnB/58EF5dXFcvCfDXR4+RnafQiGcMOq/B1XY+YT0kj
EmdcuQ/vUBjjSgsbhaRuCAFn6VHwGxbloejZS0+eBPanwvH35AZoh2Lvbdhj
1+qDNL+dXLWnnzx8CTDyecTS2tK/KYbQQJNORB6qp8JavEIRN7/8sdKathg8
0C1v6wdqj8tUtIeil/uru7vVWMjz2Bvd8RvkJfWnY2zsyxu0K22jEdWTo6z/
sy+4aCbB3SHgZcgSHIzcAwxcr8niTceCpvpxr/RbCo21D3+ZcTkIBYutBtjv
m0Vvwz1pJaYh/6IQNIhSw5FL2r2XBKwp2XlMIeC/TR2UBenoQ5IEeMLbQQfv
6CczwrgxnrmpLwoTIB5WVnvdIEWR96YCxGNB92TGiiFXamW+R6H3AbJe9+IM
8iExOXFybVkMo/xTkv2Tj7nEnagLAO26Tn1EERZcVne28+aiuG2yacoxB2tg
793RjL7PM3as3S94J75WTEKXEC1OzN96jQNiXxirHCLEcOy2j6OrbioyBhpJ
XhtSlpRTPcy8/fqzFMxRbACiDVaiTJnPWRJgq2/uGOzpayVP7nqRh4f+icVg
hdXWMiqFvk5X9zP+geqgZZ9vAKW0lqH3wHJVaGd5MxHPYR1utXU0AHZPk2J7
UDcEHOb9FmC2mokzfn/tFxtkn8z6SjW5ZICQGgCknvXQkC5uiEN9Gurlzokv
3OqrlllUPu+wZ0tJl9Fm6S/vc8aNTIQPh3ZGZvoBH4hkt5HFc5CqAyA0dczo
5qlAIfJj3rOtYymYkZ26/luTXdr6yGW4TfgS+4U2H5rXR/fXN61c9lvaKTWV
/GeKWoWjki2nhiJJym6P+ph6YC8mfNUJpdP86KCKrpp4SKA9Z7j5LYE6QLce
2Y8OBPO13nw5tC0xK8yhkLIBkrWx3lTvidBrnZ/vXO6KrOMjHgTkcJq12+5e
xHw/JqFYUkS8KwMhLsIyVjUwv8JveImoSrZxIRN9fnYtvyn3H2aOKhLlXIn6
lj7QJzbRtPThEFPr4g/NpJpZCCpeWarOw5qaDzlHsT8cQT7SjhGI6inpWv6H
blbXbrCc0BNsT28qitdK8Z5c+MX7T9gOE5lQKvWCysCeXN1VFw72nHouS6xP
1Y0AcPvTT0eUqIbIUewHVwOzqekW7xyxOPoAgpV15fhV1QetHCcNWNJARIgq
M4qloQm/bDQpbyL7XlCFMejRjM9U5sUGWab9nNuLz7+mFpGYrNtmdHs/LWAX
A6bxIj4X5/Fd39FiwsiCFX5MwqBxi/itcRC8Sc2/InAo4Dn/WiaRP0hgmwKF
PSqGzWP8XVbm3sKfbyGZnsqLFUDw7sSBNqT5SwrnZtTn0+/oI7p3GdT8C/2s
y2YETLp9TgFmoDTy4ik0MlaeZJuQUfHwgI+DMP3gLSvNnhGiXz3Hju40NAOG
57TgTvpUqkgiRZFkwgSMqjScMZrnhl5S2dbHv5VGYyy7jBBXcCIuflbKhsAV
akKJ1AhfOugRNV69nhzLauDoMxdn91lxFSY1MsH1ZU5ghZwSjfglUW/Jg/XR
HLZmvwfnmKWPKGf4gM9ypX60kzNrGpUVa2/sN1RXe9B/sL3YV4Prt2EnHp6G
VjtzYbS1Sa2PIf3WlX0pDmJ6rEZDNfGVv/dY0AR/sGIEZszZG06DhAhIf2Sb
dJSS7QvWfCJ6OCP+u4jSIpYrL9ARcnNmfCzWzDbs8MSTsJR1Pea+Ny+DozEY
b4SnVXucO/aUNEHg4+FWDwoLmw11GOB2fvvhvV0uRtGoZ7wXUsq5EDPLnvIb
1PE/mu1bgxl8epC8uowTyJu1Sn6V8nsuskgPRl0Gd3Y5KSjnnbDtrSMAZxxG
boklKyaJPEkWT1FxJ/YqkpDHt+7i54sRLXYjnT2VDb7WuRiZFZogF4tbPQi0
eJ4YoPArQmd8zxC+aR3GpgC0LkRit9QdeCiET7W38mG4ZdE+pIoeXqNd5lx3
cZ41ICuGhFoe7lWnQYz/NnR3sIXyEQUKrcUY7HwLHDtMwTgJWtzdSXZz8Gtc
LQbCyxeWWUf0ety8DAvUGoQJCmABXK4fUvlfcMme9j7ErzhL5S6lrbR7vNU7
4YTKECQbjWm7gCH63ormsJtLMsplt3EsXa64P5y057RHIswyQrCNMHmkGTOi
3r+RXwVzXauwMzZQzEMiOJi1pNPKBomnWe1py6bBA6AA0FtCeGI2Ph8RsFhA
+iO5Pf0xCGGqgAfAt02Wq8TBkJd6T17hxdtB/1w77d+kAV65Wp9DccoAq6YQ
+pS6xA5KKG1tX0q4Ws5WWauTLUNDEzrk2rhI6R9tvPZw6WWrV0p3uWAJ1BOT
YhFwEb+JH4jbUCRqAwUUk8H6R3wgKgLRo4MDS7tmi9hUNSqMBDZo5hqv+gll
oq4zJolUcSRQvh+Evlathk8rgu6cZ+LnP343/NHxA84CQI5oC4Spy2Ou7vG4
f0QtfBK4HmF8GGTrtfxehsBRyj4Wo6e13dEpNE4v/iVYHI8eGvJGS+uLHBCR
o+KUam6vPaCBu3/p70ae3ORcbrEiz5MGkMRy4w75FG1GsMl1X8YyQUJYJL5i
vo91Idgq2O5pkpDPdfEadlnwsL6qZCha0i6pdI4f54lQllrKL3JIKYgEhMQO
7Uyr1UF4th13NF4xOHNI40oIn+8VN84MPYooEkl833Htbu3v+gIHJqS7V8VY
5pGIKXl8ViK3YEDZSYOMqcwyFKNDUnA9Ir1jnPMSPzZZom2wH+Ib/VwgtOoo
ktxfsNf/8HFW/NS+4ed2fy+OoPYUGzC5xsa8AFLeOSTL1qllygYlilQQ2Uwf
kVde2V8Tpbl0IoAx4YjcFV13KdwdsXOzBjMlMP7heJoocvMuAHciEpZVoTw3
RBgghaBN9nOHlSGSy6T6IDn8+xZM5XjcJa1x2LetHkShWkq+kb+fEn4VxiCx
O9JNUke+4t0y6xamX0iqZnpCC6l8oUNXfynNt/HCc1Kcz4HctL/TZzqnjFtQ
8D3yVdnreTAEruzU9bZDbD7Snv8I/10TuykF/+Y4JtVIhcN5wBrzdJ4MeKLK
l1VfnfOAittct8WtmolK6eMkw8TsKtP3M8d/BZUrE5SXdkM8b3k9gOji8MEf
Gz/6ot/D6FhrVjmiMznf9HRagyS9BmpdqhQXane+4Gq3MSymshVrNYYG43Ky
INGU05xndehAHE9okd3cY7J9Pdea4oKK+XHjoEckwiJ5vhuUbxN4xY5gsy2h
IUVJgjihAXn5fczs3GyckXqdAnNrlovWmuSQn/ZJEht01SRQ/+26DUraBCBv
u9/dLs1Bik3HUSNuJjOlzbwYUpJT27IxE47wiKzAcqWMez66ilGFXGXEFf/H
kNE5yzlaIgLriOWMj5k/bKaSQT/OBTX8nfAsuAqS4equBFh9J/G5794EJFBD
Kp5Ljs92WXgmyyDQOlrFjh93Vyq5eJnXS/9ec+6SRKimrHEhsKT3vdIDL5oe
4xFO0XlzsUb8jDCrPZR9WCJAzu591MLbDdElVGuwEUoPisv3Dd0lgHVee+wT
mwaDZAFF5FbI/qbSlzeGyZZy4YZ1UNTMzALYWEQSwraKxJBBn7oRPm33qhRq
K7/sndvo52uDQ4K9658fl4Whd14Y07iUU0xsHAOwcCS0zoAU1JXzLsJ6743T
mgZodTcerpUgfOR6xPodf0biDsKLoSsjY2+xyKu3/nXiVyEmegM45iMsIlP6
4pyFwWpjoR4jdEdJ5nRLC6w8iL0CCtRE8gk4Rr1RGHwCEk98pbdtVajXAYtl
y5aUYvy+W7fpFUS4w3sDVLCGStcvT+bCNc97u4WgtKhBMLLMspRD2hVqqYZB
FvXwJ78Xl975uplE2hKKpBkCnmThZ9+8BWcKnenpxBtKJbz1bslr+UrfTy7A
uibJ7xGwPIaecbTHdHvA+KK9+BJJOfv/LT/fUfkngY6e22BHzDob87p/dz3w
Qou8STTvP29vWnKeJSYO1slosi/eMuo1vN51brw/EbiooHMAMUpZ4yVCzyJW
LpdP6oWhP2idPXYAH2kfm5UdwfyiW32RjthCFNl6VhvdKzyNKD/X7m8Bywir
NFSIO59tbTyhOvSA6ZUE2R0hIgfHEl2oVlTXc/oJ9+MlwZGl/vWNtkKmD1Tx
fZFQDJYFwuPy+wyUTyG5nZG9KdRFmiwqtuHPEnfN+UZ589cZZ1KN5nEZpODm
E7PrPnY9BbAGPkTFw3Y7rXcfZRyembt///DnlZqjofOlfKr1rjkV2/4LJInM
K8qjGXrYgir+eHYeJo9PDDrxsh3RQos01EyWg95BHAwK66J/lTn0ZUGf0gtA
Xo31ypGFjCtyNxQFrv0RrQGVd4bJqzgYSljuPVAIbzlsedQdg7Czl2YBY/MH
6B5ce1ozgQJ4yaqaEQHpWAOu/jiQxBZe0XmuXPIiRUMbptc0e53ZXhw5UK3+
Xsa31+WDk3Y7W9qDbd4ypdfSwfvXerQBlUyiXmWmbCDKKK0W5gJ4IdF4Dxek
JL118lckihx2u4yq0jZRci1KfqV+qQ2LYZjw99W90XMNaCAaQk2AKZIM/JDe
xH6wPhvtd+Kpo/0Il5R8MbOX+m/PBblxKCPlSNv672zIH3OyWP8HtODAbT6F
tRvGbc35BJ65yk6Sp8oaFR6/sv8Lp5aFPh/ZX5S+nukj4Vv3faTpbWZTVqji
jmdSuPIzkfnWqWDcpijwWUMohhp4f6c8aqe9AJSDDd27EElPLlcqT3T5esn7
ImvUzR8q+A1On4Hk5DKy1yM9m8qDmyTBSjVV75pNKR+5F8uXYwMZG92lcJS4
7qnq4kRfXpE9JrCXMV8lwtKjLd0tFj22NZmXskDIOj49uScIWsMxZPsTfsRp
omhz2afHWEMzJjqY/yo1EaBS2VcHd2dJsj/7qZHM2CR1QEJbshpy7d6Q3hcW
LEII4cIm4R3etc6kAah+fM1SBMAFBRkzTVnk/NWzr8dam++3WZdQgKUAYHAL
1KC233p/HMYv8WHfWdsdSBzxJP1mN4Dyimy0TQmmEAMkDaK0lOJcU9LxIsys
9vEHvfJN5l+lhnXsgSItg024pm813VHQgpsz/iXXdr3Dhb2URe3i5JpZMY21
HsacJiWKQFxPONsdkFcRjn5m2CFphpdwg6qNxlsanpPxhJHe09wfsEkE/JPk
dswl6g7FliucdJ9uzGyaCTj16FsoF2AOo/xaOmyl+pJrEcwdjwjv3Ox8qLa3
HY+an0TAfVX3anJD5P48k8GG+zvqzS3rIrHTueYqaZ2cT+cFFkDLnSaUwFAb
qJEPAxVwXwS0iWugxBmh1GwW0V+OZfx68fEsqY4VhQbL7ck9sD0pu6W99bHV
29kgd0mTFojmQVp1Y5xqvYIXoL+gVeqWRsxlKDfb5+MB3jgBGWTYb8fAD+5c
ofXCCLJ4P2Uje8IvI0/CwNxrtroM9q8ow/g+NVf5GR198KAVPZ0Ng8GTpTM3
mcqtKEohYCqyXV2wDob/YYAsjUkIbicobF6FDWBNxArghIelWXtsq69snh9O
gtoZzvXyUeartDTNUghsvmqzwidtPX7AqfhaUMFt28MgLeuZZ3fvB2+k8jjR
rMh3TYIPMThR2bpci98+xwr4QCjRpeEwSeb8S4dI4SjilFwINIjYoPefNirH
+qwK8s7X651XoDafaA9cpC80r1WM7spKCYYNZ9GUg6B/T+foy2s5CK/Nsquj
uofiojIHp+W3Pv4FMvuwKLRlXsZxy8nKN+e+nsGs/SC/RWvERW74/i8eZ+D1
Hj27uxid5j8aGwmDr7L1jXAWxqNqSs7pozQLtz+q5UTxTlKmZsVE+luP/DPM
033OYpimscM4ynNmeR+qjWaeAaNTvIY8VPuP2Q/LpemMU/HjWeMUsVI9ggGv
s/Ih1zmHv0q9ISiqBS9nBPgoKH40mO80rwqhqY/ACUit9RiuOfJEZrnoU8J6
aMMX3eYFuIETAFOrkHg+QcS0ntP5ViLfm9f3LJpwl1FKbvB8xJXEvYXpJgZ1
3aLpReiEMNjMJO//7dLy9RBA2uFs6bgRzGSA+a2nDZD+J9+eWmOLNvO95L01
uk920rAi+iMcfN9efvmJMRuwDFaCAL8zaSa3gQG9A9WUHGw8SamL1nOCGKGA
C3Em3kEqWFPPiaHdNdmIHjWP6f5Ot7olCHvTP6TvmxopSUM8NIivSl5Z+o/t
OOwiU+FrN+086ymCXiNJLIFRLhMAqOVimSsVXlWMR9p7g8pYh+3oXn9wdpwP
NrxbK4AcKy4SYjfbwnpAlvOT6+jtiM1dUb2kKZkzCwYdE6H/W9XkLDTfSvpO
LGz5HbLb+P/+R87LP+6oD5j2Pzrrq1bZMLRt+wCy/RokRwaH6xzpEIMGkEZ0
2SstOrjg3k9FA786F6h43gwh8quBikSSzoMucCrrr8mIQaJ7xFnkXYd/Vzqw
IWxrPe3QS2w4HMD/YAjYp1R6Wip6pClz/JWzadMZlIUhX9uMRsRg72eS2QCJ
EJDmkAlEO0/KXaYYlvA0UNPTChQJxWIQNl6+X2e2QYQp1uJdRujQpoCj/aXP
TvP00Ur6XcEYFcKzGI4MVPGCqpRqr+ejcnhe2L2qy/lfQgBt6BF5UvaiOF9a
bLEQYaJykVtEdNLf6obU+OK1D1wRFdsI6GZKY7vMfEVejiiWGg3Mp9WcwWEW
m+czLgdVclEkGKE3j8J+ukdE1BoizJiTW/1bSSTsr9UbCG5jK6hY4YxVXnqz
rAQsYjM4vzNiCwOILDXg5NP2LeMFbUk5fbNudTXmet0yxJmBTs8fLoWQ99AM
AVbdeSTGaqk2we49t0kKSgbUnwNc2kztVL+EWT3YsMJyOzjSkBBlv9lE8io/
TWOSY8/rui+t6rEclLrA+MjIuJCBakMiWy+MIdbrNA3y3WUSZM/9ref8+qUK
L3SJzkSOlpiYBipmWrg2XifCWmFBvDjbBHHY5mOzxT4jj2Ho0whApGujQyNm
8HFr5oucgPEFpItX8811Pkd7KAuIK61OJUQiFf1oXnBcukvTnD+CEyaN/Wb+
ncMnX2HUZibf0otZ/IbcsKdpLQ41tcgaeYZB2HIDP6QiOSC7JZKsjOnHCGaO
MYB9eX6qiPanqF33pEFkvSlvTAfbdibhPCET+nU9n5Jp9It5wGTyERHByCpD
H+SVVeMPiFfJfjk6sdMk7LV6+WSCFO/uAE4tHGhnxmQ+sDto7loVwTd3DYYp
ZB0/oqTbRbEpbY3ArA+c85a4sq0rlGFMFgVemdkOBGd8XftkC/IyWeGNh73o
9iS8deZ6IxBPw0ey2nx85CX6LSuea9DrJfnMXV4KCy1G+Bfso9zYc57Wg6Zx
fAo92gvPjzWRuAafS0zSpsy9a4K0i9PEkJ1Vm6XW7oL7atNVyrRXLyq14TJW
0d0i/i1eMnvd7n375i5BKQSqqgtorjGOVqRISUiZeFrO1Psj3/52fNT+3xWV
kO7kQL2RrT2wjV+wiE03E3fnmhy4OzLPXfO0SDN0NUuD00gE5pn5JwZU2D73
CXtkMIMrR9R4jbuG4F1FwK0phYv6fxzQCdoTP/b695HzhUnVJfvvzu0JTKDX
e3DmdUDOzKZqBJzGqsViV4AHnuH0wPZrQrCsV3rgNU5eJQS3yg3jbJPnXrtG
xKdp5c4OGga18zXC6Sj+KnSCd7BMR1dKxKUrC6O5EqMZaSK5AfAwJEU1bIkW
LsSsmvwtZc2RhluCPZNnmcnMlY4/CoTOdyWgtJWoDXcawXhqw77rodFZUfBP
it903zbRdQ6ziXlp5Ga40Rc5FL81URu0xwhPM16HtlP2kUgIQjhsdLXMoxil
g45rb6QuardGETtxkwxLC2YPFpQSC/YcoL7NvnklETelfE2UzL8m9TWUuCQ6
6lRpsdGffjZf7U0u88liLu3ziOfMyQelbKPZMy7QAAK/mCEQcE7Omm2ykfnj
OB2o87ASsMqaX6TCW6NEXYGU2s2OJqFPL+NEVzKFC43bzUdPGH6gFcZKlgnS
08sutL02owfNdBniqPyDn/TcR9JBCQtPCtRRCLe6uyeiy1CNqe9xocctjwUp
cGnPrGfXn7epOXtV8BM+5zmKpMy/2g56BZwt96lmdKpo3Vf2Gl5kVfIWFH5M
3DgsnRAiEAYtHTOESupIHmeJWjvp23SmgFB1UqA2TGW8cHviYfx+Au17ybMP
ITIys0Ele8f7b08NJM+4DW+0GIjCyu/ACGt1ij41WPDfE9iR4+rc0lyH/WOp
WJaiLNETXDuMgG2xnaTWH54rYeBxjeJaO+G7lUS94aO8pqs+ilPLjId4JDOw
jbfCus8F8jmEuFaLGTlnebis5z0zPUOI9N52UIe93qxGNmy7gfYwESUhcYzN
k8prbdOF1w2gpVfGd02hHk9pajoQr53C85AjZvN56EcIeeUS8+THeFI9neJW
wV6HojfnFfA7ch9L59H1vxLbksYs1PVSIwZd3VR6Hz03f9YtecUUmKhRTuV8
oixL4iHQ/8yWFQoeJoQmpzBV1TV/ukGb6KTwUyjdyWPOD6OfpTywSJ236icy
xUtWF+ZKlFqftrsSWOxkomk2/teOM6hfMQTELjJoDLhfm8CDVxbzQpjPRwVg
D3nxfinF/94S+Iwt7C/PJQLy1XkEOKsLslu06gMJIkGrAHi/Lshah8m+jOq2
A+JtN7id/7uM1PJXVmCH/7/Uy8lXI6TK1Hw7WNgARpixKGD2137t9M4vjVim
rjvko5fzr+q87mbgTs2+ICuVyohbMelWUj36byXw2mM1bx7fFfXbIighIvM8
5DrxmsMgGRMzCRRTzXWWurCqdVn1d9+EAO4Sa1prM1HbYKx1vEmiNmXa7wZg
fHn9qezRia3HWBk3MILVuvBVEwGwwEBWcqE+I+0Xovgrll4vf6EJqZFI/3N2
WwbzHD23uj3XnP41RauliCAxc1Tns8AaJXZzRP7HZRYVN++9KIYNYTPtt5xN
FcvEgxiXjrT6q0TBIL5OALTCbYTfvCc9LqeSBKOt1sDLejz4KhWCwjbJ+aAP
LyxAPQSu1AmnlVX0j0XBSSaC2m7Ij77zSDT3qw6W3Mb/E0nnMz8O1mHW3tpF
+D1ncxgVNhgJVgKW26l9WDR/tTjBotetvPIWE0aEhMFr9Hh2msqMg6Ye/JOg
snuUMa5IuGSAke4nYIBkfbqSnqYm0sdPTZnS4G59OCqcUZ86NAqbDRLhPc6c
5JSwB/opy5IswQ67niOGpqIjr2ZhFIeSZiNpi2/Uz9Nq9g0jOZvGocR0hnlm
xq+twXDylpXqxBKfesfKmsTqyIMd9GSpHgIbuFFlC1eKVoZDKQiIyQOCMoRM
ImrQ9XIxvDW4HYI7A9lAFQZ4s3uWc0a8bhkeznWK0NfTWh9e0YWKFunlvFwL
HVpZRa/ZPP8HWRu2oufAH1bwCcKILirdKS7U3Y+ljtzNjvx4YXzpN8nul1aJ
5+mLJQLkgALTKXMjFQY38RrNWljrVojr8+DGtYQKGJc8jWgNcv5WzM0iyNu9
PP9Rc/Oh9Tf9BxBBBypRJCLex0Qvr/5/p/x3bZnsEEeBfId6lqjlmtuF951y
cJ18zMB6n0dy0pVqWlyvBzIMWqM+zjUqh98nHMCIaZtNPVNq19tZFEdAwnMZ
m86uEtLiRTdnqIouDes8X+MD4nM/EjlDLOsv0dJWrkpuAinZa3ZeIMLmUUfo
hy2iHTL46k8nxxwFDTg7ljhQOxtdxmnU1Q6nmT5fEDq4dolClR8zQcnJzzkl
mklB2Y3i/3PLcXfeOE6+hx8TiOsa86+4n5nQNSHXfoRdfQzW6bD2jG4fEt6M
oclmXuC5w90Wx/6JG1xtm4zlzDuLM3FdD2xZOQua/ravFWrjEoRNW4xXUXF3
j5B6CnEa2mKtQQ8Bdf//OwyYH2ACtJEPvzRb1axX3Wj3DrfHCnSMdqPUNTLl
n5mzC7N7jRWCKGKmHo5m4n9iGnqRfvYAP3ZnK7mX/JZDsuUa5Doy5psJg/Sl
tpdtcXXTmk1oAnEGNCSlsOe6Y4+5SV3U57YGYUFhAsGr3kCIEIrvL4HMvd8X
bIvFezImkuYngJBlF9gwOCXaRasgJo3HsaYte183xwjCrGKbE02Ggcrii9sZ
j+WrBl/N0mMemYOQYpDdxb2UujFNI8RbJ/wSAA0YgCAmImB1L6CV76RIrFht
q17faoSkqT0sN2gvGsC1yKCgUpfmZ03s2WJ6BsFc16VY4+bOVvOsGj2NPE4r
MZGXPqzpSm1BkwM2EDT6o/lAIgA9AgI8zkr5qxWvktzdIaYsEQ0LfVAlI5j+
RN2Bo8eSOWoB+3ubm/BUccUZQv6+Z7INoyyNJq/G9aq+LZAZWZH6tkQdGb+5
cjRaLas9Wjk06IAft/bP1EPgBUWpXvtEMdCbMiiY9NE7tCEi0LkCAWsALPCb
FGUsLwrT3Zbna1x5wdzZ+mEg6U1/tWKMTKa7HRy6fuihqPppVXfTScMoJ1t2
vYi4sYUk7gnO0m6zQCkGpE+dWLqaAVMciAep4jx0xMXR72fhAQRsdKc56RHz
q4XYndcasOlzBoHBKsfcJA1n5wXhoPfcKeU7/W++QNR+o0SV7CL2JdWQUiR2
gGjOCdSAtGqZW0Kkw//DYreOxX1Uukc5QK0FQXP+G/686mKcaNWEL0Lg6qwc
Exr6j50nmgmHvuaOyOVCpvV5tbA3a6btrGsEBI2rQiq4GII+I29e3ABFjdIG
iaVJYG802YOnVdYb8dk5Es7oz7vOvD79D549Al+2Zf+ibN2NG4uE8Jir2IyN
LzzTGwJ3BqGeq44dee5zKgkI6BJl+b9FB1wvbpuXEYni3XftmCmN2r/Khmi4
HE2BazE3BJV8mFnSJ5H/Bhqx8dl3+ox2AssQFqPG5eTqz/xjiAjU+pzTsnky
pZ8bOoliPuMLMfz6vIAhdJ9ykxj0j6TqKi2Gx+ql6hySGGmllCDMLz6ju8xp
Pment2tFfc4xMCEdIYrWiAn77D89FdvBpgsnl5KI1ocTNekl+ayTQLCCcIdn
vC0GfR0ao8T1omnCeAYYbeWBB9JaPFaQh1QddtOYlxHjXAWAHD0FhEf1cRhW
vU3P8t3jon3GFCKhvW9HtBGkopcN/7cGZdJcGYlLZWWFSGzvKMMrrJxreLCx
ECJE7iF8n0ngV4cFGAFplkd+lwBGZxRdH5xp+V4O5NWgPip+BrS46P3aXZYe
toPxpWBcFt2//el/M1If9j5PwawLV3QhzOcMJxXAnoOGtHZlH7Gsl0WGcEOW
H6MJvZuNdlUobYRH9HSu6RyhagyoyNILKqyNeQWGYfD4xZwgf17NK66QXQ52
Us8xWVOmkctM8Klrie58uk9piEXFpGYYCLKLfYQeN2ZE8RDSdIyVbNPNehO0
XdQJiInBF4HxIUfubiNx8vIZ2v5ATN3PTfDpDyq8OUXpkIaETC8jfwxH6c9N
UkFtNrZ4z31/qUM3XZFdTLcdpowvhdxjjP0S0jSQieVVpDbI1kufui6nK7Sg
PhPKfzLmSL/27vjZssGZHu4Tjp+hwwyk4/5iNkwkCKOwzSR+1L2PnQAjmC19
uWpoeGNlpGhXQgtv2a0aE6eU98p/ZObzKeAT4bQijAKrtULdb+pohDRbrv/k
+UqEpe8NZHXepGT02hTFexbsSFflUomSLHbNbUuh3GjeFkcVdW9Pji1UIhul
gk+j+1JgUUD8LvIJGT7g6zG2+NXYSlRVfcvVNrEFQuekvzJiPQkV5qIClX+W
6gwA9jHuH5JyPOUHQz9SbtmxyfAgS2XTEv+WDxf/Q2ypV0KJh3naJA1mJ5ZE
rRelmND1aI/H1VpPezJbD/UpnTuJnsL1Q0HyJBcYxJp15CYrboPgRnO+t0ZU
3fO1GBYyx3/W9B59fAeK8ZG07a/+9nxbBamA3fm4hLp77m0Bkn09vh1CvKqr
iTD+OH0Vq/Dbcx4Bx3hqyz8TAdWzmpiLcgCYT35ybxCrYKfQHP3ldec1GY1V
/UqO0Keei1Jgae0CceR9LmM2bVWYyPUvB0OaTxP/K4vzc6o0ccp+XeNVaQb4
lRdGo1KZ52ZrKiQIRK3vUrUc2JY2KIqN1eXpD3yRys+xEzSqLGtY+q8BxLWf
3mNl2I+hikskFEjeH3do3tu6ObOzniEZ28Ta8ZgXIyCaWCuKubZjLgMf/F6P
4Al0DZe7yC6sar/JYkBaxW/AZtca3akHBPVNkOwTgZjCvWI5ithaMOh9hTqI
CyRE6oqzJwYepXm9pL28DOqpI3x8+pVPAkDoo1C7XLQG1gaFu8DTgQDXQlnn
4VDXXnf23Nmc2LvU830BZT4LfT2hruxI2fMykimXFGwT7QP31ZJnwWzQXrhb
AoUlDy4nX8RZPU22jr5U+QFjEerMgdP3IiZvrgHOdP+blOOIPGeATRmpv6Eo
gyrjTLYoL0pCwWrLZGohW/as1t/P389sQ+njZOaIVeCjrVFulOtt0IcxsIFs
Cy8IuvxTc6om1eh8wSJtKkZm9CE6w7pv1r39W+xdEmusA4LZNa1mLLhbKCTN
RZ2ex3Ifi8AhrB/X6VXSKs4pEOXnglNl5nY90vI1sk0e1dKKOn+jHh7HIv3E
IDRolpaETH7DYJq7TEg/ySAifvRsCIM1iJ+Du3e2bUZwEgxYXOW3wIj0iZqQ
lBewsL5s8wQtR8Jkz+A5UOOd4s6cSqS+FRZUHcB9+9ksri05n6xXM1Z7D1XU
lCOmiqZ18xG1d8ehBmsshkoVrMuxmUlpD8nYDpyw1cULAMAypQDyVIF/MQJ4
krnC3R9jienlxIquKNEnT47xjm8rXqnNze5dBxkfSFeJK9PBf3StPQtvceIz
7QBDi8zo3CZvx4V2028fahkhDGx5Sw9RhrkyWVngeW0yCCsafWCTen7wNx4S
mdBP+v4MzSAGCdpm7Tu/meRtvfAQyK/cirSGD1/t/rK8o3dzgSaRHicYkw9+
GdMi/36zgDtecWLmJR3tN4mrjEK6KWOK4OuHl3qEmS3ARCjuhng4yNC81wtD
OIWnoL8jzvJKrE2ED6MnUfMqN3bvwGn6OUeNNtPnGjVUN7HIQIFgu/SKmpAv
PkanCCHm6PNSHwvmW/QE9V5vQvYYWFegAvbJCg7WdV3aVnsoWjgkJ29QYCFa
mUQ5Edj7SWYqwUNC4cjd0b6tVXnOWMxCQjfIFv7rEvuc75R5Hmy8Tp4YtwCK
O3EoIL4fSLM3+rN/wHk8TkgzgHWvMk+omL2QyjFj/NcKTXgenH2l6FoBpm9E
e+5tRZixfiF/KWqS3SxAzyHWD3jNHRH60INY2F1I2L8yguwgmlsdftUxeGeM
SPZ0NfpYR/4rhMvallMg7FHvMcljm9NYtU5U8gTlABgYnG3XwE9Y17jEZrRA
BCGDfoFrAH01cN/smQDdQ4KVTu+2qVDrw5OKbIVA53j2bVJUjkt3jEK69C6E
0SNt85i8kOG4OXqa5ewrVsaq8fId2UEfMc3D5yw7FI/eV7oLlGtVWCfSWdI9
e2Fk9cj9l2xZ43wEtOazZ6NPvfgA6T8k8eaTKYGK+QDM3upPhWLQQ6Fkh7vh
gBSQ7tGQsMWBBRCdc+gfMQsiQEouKVeg2SkJx1po9N7Tz2dU8C0IPvPZcAQA
4m2nPa2XpxFcbYu4lR3ovOOqYuR3GDjtwPB5lE2V9IFAVtjtSv6/SmSCyETj
gqdg/yY8ZwCg4nYP46c9mtVGoUyoLXYE6IdsnhmvnUd+NlOQ/3YWf+l1KH0c
p9jHKDlWEI6DJNgK/XP29p35h+rp11fEnAXKegsvtJTlb2J7YOzUa0iclsAB
wfhVJNRf1HwUFB7IbnffGs/90WPlpkfX/RtuPUHQN8kq1n088lL6cpRw7mQ9
GMBmhaZLkw302UkNC2Otkb2P4Tisbb1tow66V6mFK4hOKmP/ywWn6r/7lAUU
Ue94Kdt2OKbhp1wbJYIkBIM4JTvXTRrhBgBJDpZv/cMxdtSc3KpiO43LymK7
tT8Y9TYixNvsT8ZbsT3O0RVGjtAZIWzm+8TXmCt0FnZP7+5swX+xBTnf3t/6
4xNgxFLEDpdoroFz1ws67ckAT7jHB/Iq576myNHouVFRe9zhnihm7TiRDJdl
8nr87Bd5B1zmwOCqXD20KNOJZtj2YlML63RLKpZ+pcPm0owWIEovAzpYdO1L
/x+LvfYQE5LBJBys9a9t4sbHMHt1jWtLDaJZhOkf4xBE7koIk+Kz68JYflV+
S/FuMjzV6ATG/P2dbmG0NskDiBMrQlaT8j/VzwBbZW6dhbuDjIbt3ciXiuS2
V0jbVD3AYH/5yKl1JRFykugs4VA9Gsienhicmeh1ZmraVUp3JNAFhP8w92FI
mHAJ5GGDFaztIHG5oEBxLMk7gOF3hoWFqxA5ivEUqDqNBEbE+4i/CfEs5Z4E
83GidM9vzGmGAy8QDEUflWaQke3N/UGpk879FFQn4Gc6JZdmsN8VUYCC7Wnl
zOb1yRx6CsgWZwm2aRF+kco1IsAKwNrgL3pL9VjBd6RcUYDdhzVK6BncxrDA
Rig/Yc+byAHpVf0TJ+G+wtlN4tBxR5tn8VcHyCkWLfj9fLwrFox50uBAxQl6
qU6U/xd4ND/qobWU16iHHCoYGkAtFwOsj5++GgIRr6oMAwEHlDygmM4YEc7K
Dh571gCwZu7K0evfkc5aeq+rwUPtZ4HO9E2ZVGpA/m3yBLnqCm2qHS9b2620
uxXEWcuvaIDzmum0XQS9jpkeXKuQkcVymV1HlZlPdmIevQlseMKXcl62T0VM
DHvQBK2EreCgOThywLlnKB2iFIONvcZqbKq+MKyq6TPrDnORrUN3qv6RwW2q
UAq5/BvG2W/j6weFws2ZV3UmrIHzT2uHT3zDYhn9rjU9gs6OD+okqaN4iIlu
5GcU2SAYlzc3FvjgxDSQz2WIiDNzNPyYZTUwnDr6nY+eNRGaagSp7IZ8IQPZ
S8x32EeEoGVhkPVHKj7JkPttQRZsjVwkIR4bwLItL8Z4z1hZMPMEbWV/gvXU
kzYi6x3ECktwTCmUWtkwAob+uSlcM3Lv/N0nGxbM2bBoa9rurKn+iw4AtVwu
/UUpoO6ui7fKglmSZAx82eDWSvkMWgLAHGY6pcMxqsBnC3/22MztfVl2q1rC
YqFag1X4oEXcktJNClUpdurmc8MLFMjloU1YDUOsLLSaQQTH0fZsYSID4GTU
15ggpV7yNB4AfceAkrFaoCQ/U5NtHczwtLxfTTiX37Uze5YLMJf5+zs24Zgc
yEGgG0EbuZP5HTrfe8eNyDIB62d87jCRrc154Fkwjoh1as49d6UeY9bVgEpe
sISf4aiKyyEvXPjvrI/83yPUlbx+WQ04Fn5637NBY7EW1YTmbCO8vuGp66cY
RK5msV9iUPcT78KsDkTzzoBiG/nam/hbMFn+im20zamSrQnsQGeASThlNnLw
84Tuaz0KS+L1Ol5m1Oxu5o0B71cS0PFeuCcuMv5IH0CKxAr/Aht6+Z3a44mC
4A0EnF2EmThvlF9D+ObEdUvPBl/WdGdJ8O1OAFHDO0bdwbzcwcY/zpQb3xHT
lTZ0MjhJg/6a8ua9Vp0F/ltGfG3edi4XojPCgpc857jrAyIVRqCV2nB42ar1
rBpddVc89mI3iqFTVQFzCvfEDR5AVSB+J8npnojWBF1W5xjx8suz17YEI6ct
x7ptlZGhfCvCnwAhxlny4O9sqHndHt27oTcJQUAZWDcS6GE0NRZO3CMTVjCC
AK/beIoe/anOVzfoNpU6/NkDgGS6P09I0DHjoekHWBQ8mu+lMUFE1/vGViP+
sacjJQzXRSJriE82yFxL/1kpJEKt96aXRZbaJJsOP4MxvbUhoeCpK2sH+xkJ
Kwsp9oN2aIuGyyRt9o3bJXYOBYLHKMxuPxf3In64RQHUnscgfKmHJiaezuX8
MDdI4HxI4Q3kLwL6HCiWMxEqtO9d3CoQ72F5ZRpwyAb4EOhRB5cEhP2pHQ5o
GFduqaDyj56nFAvVQwdmgZrV3t9X3dERurWDiwNMH62T7JftySS3/AbmJoBa
9X1KUveMRpw7QKePsAmnTEb4WQM+nZ6kSsHkjfSdHzEX7aMsTxTkyPsjgT0M
PaiTQ9fwloXHeRXCm90Cpg/tPK34+6WGEpMTBjTqDzHY8VEuMHQcV2Z226cS
Urg4zgc3TAGPfe1DTxgsXGmc1UdD8PItwbsHbtD5oMeAQMUHHbl+fLRJGRjd
4dF5k93PClL1X7Arv85vokF+P8ZRcEUUXFDSGCZbKI0LJhJBrTV/A//74jFd
hAgHS/dJHa0xAH5hCgUi1uvzr8aOjx5Dggei0W+D4ar1GguruP8mKYukCasV
h1JnEjLcvOhaPOewtqfL851gYXsDbMcep/d52P+C8BSFtnQ4+yhLS+Dlc88y
RGPIXaVgg6HQB0PX8jjFivbtDcDve7vMByIHaDg2JLGPBAmTnlkbpqsaEXC/
uF+AnkeDQUUh69q4oJrysJ9rpFmSNkmj5cqB0xtRcaDVNKOkD6wq/gX2FSC1
vpA47A/90Xk6MvwIDiQDjTbs9coP43R3o0f1nQjsIaiIvQRhK+cZu/L6+/Xv
6+v+nOuSdJQ0NV9y+doOUka5F1BTHiKqVjh1uLMoEdsfdbFKUr6GKHRbiVEU
izaxB345mUi7d0VCuTJ6BjTEWD+piHI20UZIu4M1ct9KlD45fCTVQkjo0GL0
axpnsGiyyrjQA6DCiK4hsHGlNBwZX+liuAdjkQckztlQf6APytuu2yAHvzs7
9bQnK//a6kvARh+E8g+CUahJi6jywWI0Ddw1lwpURdT1WGzFomVI6IKuMzNR
iCLCvwUrf1aCIEJUmBI0RGtK3xBpNTJ5M/MHhDEAANtUY8dCLrmLUNiBvUWj
PBLJBI+Re51AuBCWQaHS91YlTnANJ3Sqz+iahif1wfV93vtdDPrv3BgMfMRO
M2lMRIbsuDkqJpBbQ3qOCsmYyQvqkhQ3M8E00Ia8IVkZ7hN/cDtdes8hJrxN
BqCIv5jCiNjyidecOMuzdCj4rEZRVmWCBb4SZPHCV/1rN7YfihBsvtOnSAzA
hjLdIrJmFtruY4QOVAzvDsfsNEhUxlgivfUBtv0mVA4ktGEzQeBzyda4U0Z2
JaIQunJ6JYIHN3oKbYhuJ3H72Y/zIdnvcFv+tgQDD3ISc18V5272dhPpcouu
kR/tqmzD77OTnVVGq1sc1/zM3mRnVbgvrHm4EqU5JR5meCTT8TANeIwXeQY/
uSas+wunDFwZXPRWck+zX29XB5PW1kaT382FAWAC9VaTQCA6dJCi6Ltm1ZG9
VDpOjEx0/kP95e7vYavqoa6Xa8V7UmvVbk4QwP/laVU4+BbohEZARdDDE7hc
6Vf9iy4dNO7mC1d1/wufLEbLcIfKrqMLcz+ZQPONCAOCaPg/GHJ9ge8Iti+B
Ow0finKZNp0yXGtgr2IBYTQnCSxwR2TDjz2DNiZDa9DWyVkBfrqa3SyOooAM
ezIY/RDov6GXWaLSEqx0EVSlGvzn9Qx0cWSfIo06IP/qsi/QiRnZNlym0b4q
dAJQcietXWEEgecSnojFz2wLNscOFSGsksQGanO7plfbAuxf4TUl0MPcEOsm
Iwk1uaLO6/htc3uwsJXtzsWRCb68g/NKRj4J/AuutdbNVnGy6Vqki78KRNAZ
YabhnGgDcqxiH36BuG3DUP5mg3+ujfuliNnN4sJi8tIh/1rjYqAR7ERWV4U+
GHG1bYziSO7Dhf1NU6w5mn+1T762YgTmpscGJULaoaFopgLoNnfcrqwL2vIl
6t013bHw4sdELPsMOkFn+Audlq/2Wp/21M9PxryeyhDT6fhgNE0V4OrtskGC
ANE7AL2QztxPwqRjLfxRrcjGXxav1sUmYvQuGgyS9HRqAsa3s6115sg3B3yS
+ne6fp/yo+pvRZ+OBZD/Qkv9MuzlgF3cyrbUAb9I/UN0bDul5Xrx05aIlY8u
MT72sxeO50Uha/Hw/k6/3Yth6ngCCzI1nklQchrbI+0NRd733XIbPMBfVM7c
bwSTIHwb7YZArbFNXS6md+55Rg4hqxgVAA1NzYuFxjwcZiztruLGdvXppoRP
dqBqf3n5NxXPi0Mi6gvF4R2w5JmAWQ1V+Jm0Rftjl+f/Elq2XtOkuOT3FEdp
EGOqyX7masnkT0+lOPlP5LkZEMSvJB26XuezyCvz4Q78fWw5TsHfqQ7paOd3
d28/w/fAt5zi9MCtarKYEr7weqUR+rF09BgpmsgYF5DjTMVUkvkbhOTWTM4C
01rT0Gk47Y70HVGu+bE+brocvfu3+ijPQ9eRrUD+qYFMlVhblDtzqAbYAxMn
PX/61zbs9MWSFx4cXSoKoXbi8kmUZQS/iAYAm2E2LOLO9bDVx3S9ld1bW11h
QJr8TxFdjmPhYQVD6Fqc1uqVyMnjRGeLfzKyAi8nIir7mrvhMwhAo4nnZhWz
45SbyYf2d5GldsxdUr1bCixo4jLqhoTMvI+xQpuafgioRBqICSBaQQa3T+YN
hkd3LiR20kKgMoo5EcDFxPGIUeUCQo68Z0SdSZ3x4vNRpYSbaqv1Fw7b5/Fo
uqXBMyPv+sRzUMhy1iSx2h9H6oVcZYIo8AaZzRRFm/jnO889+LBj6ZFIsGxY
mtTtOpKWYCgUDlzTrTMn/PNFk7puw3VG7sh5NDIH34ys7gZ8ZzX58nl5XjQS
Smxw0TpRfbfWQSzdaXy/yJaz2aQhF8jZZ7yX8/8a+Z4m7FYPUNaRPPcgz6pi
TJMLGuZ8Wk1ti+AQLJvHuTocIp3WoLqxbUIECxsS/JaVlgeNS5sR0aPaEKU3
PUYdOi9NB3FbmdJtCdCdcACuCVLE98Y9y+20fnskTKbr9tSp3GPogWZG6th/
PwSBmXjdJ4vEXzzDe4GPRKb5wHmwNBSv5XjLGIwPfxoKVpss5QNQxiu7wqDw
rDIITykIwUNddyq/2ZsjNm3SNRwGvQyTbPOKijQkwZ9RP/UUFHCtP2XhKNOP
9O84HU7juVoZ7A54u8hN/tNK8D/WFShCS+p9gRPXnKNFcHGXH7eTVvE3x4ks
xRxORpgxYxpj5faxxoa0nznwVSBMCfse0v8VwtHTRb4DGTLRHLu8UAH9XS3y
GzLEHbzmWq2ZontKjv7274svr4z0nWhOmAhxsybyDC5BviW3Iv8aEGRGFfgH
aS7/Fo/drlB3FmTQQztM7WUwERlzXjMLkW5XeZDDzYWKHCTWFWTw733ZHWDl
quzh5PXy95ctAoruuobL2ef9qwknxU7EmOA3VxmaLhg2UxKdNd5jrtHZoQWN
j1wJz84/kZ0Wl/DwJS6gAXl2oZDkmFLg+1erns5IhEO9CKRWRYAmNXBueo9Y
nV5YNc09Dc6h+nyypFeGTYjjqItqmR5m0BeO98s9DZu5W574e3KQH6qLVSAu
bihTRC3pWF9MAllGujMPPM6DRehd4VEZRfKy7jcC0dCnMXt30WWNEE0U16le
sKkOM28j1ToSqY+VXgaM3pLMrOuajTrO3Rw/CRh6qzkmPQ/F8kcMHfujOE5V
mY/XK2GyLVQI1Deojx9RQf+tpLlMrd+JxnF4Y5u0oqJoJ0sTjoPmLpLbNEoe
mkf021thjvU6b/N2N7aoC92Ci8llc6jf9TGkBaFezZ9HgKwIU9GswT0t8JB5
SeyTDNx5zgN5bhAzWCi6/xNKC/PQ/9UzvvXSWFjExHZCn3qFx9M3qalTznZu
Lvzm7aaort1Mg1n7SJiT0bEZrv9x3DcsJbl0V7HtoOkbapFr5IQ5zYAsnKAR
T5UdBmnCrPvUEiGbwAgBWO/mdWwgx83Tmmt+1sig3tA8MbZaIcPwlahvE545
am43awpLraQahWKadLtFGWx2E2bHIzZygPSvqcmC5qIp/uZzcyaBNburLVxT
yUKepiSlSkBfn9gTAYexfXJCvGl44rggUhYI2Fr3OLJ3IlC66kRvoYIkMVxL
qmIieWfcGNEZ9N7wNiJHnHd7bLSOfpKX5H6wasOglTiW4Q9Jn7B15kah/YVX
ha8DkVQlJ3V3OxEiJ14o8rXNDPV0f9l7c0DiWZvPhObmXICM+vTOp6YfDzn0
xmT+tYwQhzWLcAD8Kwu39+7psYFTkdmWYOywJMjyi3VVNE33c3ZJ79/CCmJd
BuFnnK4vaSJb2lnvknxHt07RQBJqcnAK5XpSLn+mJzCfS4eJ14UEXjzCouUO
uMc0DRqOTAFuUa6uzjhbXw7+1L/B9koMmO+tTLNUxIX1Pjkbtz+PKjtS8buI
zLPvDozI3VsyOkeV1IviePwmdoOKNcCGdu8FSGte9s9fkixnwcykfOKeCLBD
wzXSJ2qiohr699oJKVjJbFmyU7Z2wfDB6i4a1H8cxCHmW/DALZzXwWbDpvH/
7ooVats4KoBz1aRXv3TN4tB1yQ7kmKArUPq0qddDGEh/iSdUC1m4ZWiVWaJR
T5ypAda6MziaVKHtWrcdhv5+DVarUSNrjk0Ws0nAc7idGn0QAJHc54u5xb5U
1O292poC3XbwugNgXvOEsFI1vf3/1PJ37dHSU+NabAJ6yeZCTvfNqph2C0OI
SwK956uiPEvcHFx0ffNHAx+NQDs/zBykf4PVrdsATLjvoeexQKIyjaoUcqAb
Dg5oADcs+H9weVDCWXken6KltdoSsEr2+KxNCSwWiF55R0OAFSXU2besV1Fw
8wIsAPEpy3zoQMEy4/dUs68qST0I/utWHQZ/jxq//aejXRthJIdx49FBz7iL
Z2b6zkwzKoj/rUWeBjde20FK7Th8nB0ixDYO8JdAMbEKiSrfcpDXur4WyMB+
LvI0E1v0vocdsAnX+5ATUnGqF7tyR48lmJeHbg6Tr4CvLl2Wtjjvq8I/zxTK
cO9KREtREWN6Ce3CsrcCiEYlHu5n8eYCweusY/OmrHBzMmiexyZ+nRaqoz1t
cmC4FIqzeAJmthcC9PeBVS6x7A7uBOyQqxsLsymPayqCH+GpeBvGz9QZjwyu
VBujtP+SuUwgJvGxUFMvsQRmlUyjM9f7R0zdlNWeFXT6aD5B7FV7RUGoX/wU
AU6a1HbTlFprDk45Vu7ywgIHg7PH44bC3hAmw99lpEGkGac+hfXpZxds0CnE
rFZCYu35+7A1EW0rjtM/m9LESbxhI3QRnYkB1znujQOQSXzTYg55DLKmadqx
jE2IcMb2YJW1h97diZGdwyeV6H3+TJfQiB602jG1e51GYCQAvNmVBz4aY07X
vAzVp4GlznN++A5F93WfnQyp4rZ6p72aJzLqQd0XAVkEQfl5gfBo/uPvf9NC
LqtFjTQIqAKfRykKacf9T+rwJ5ZAPrphovqCOsAkeaS+CFnX4Z3lGjiqWIkq
+iwrxLEBzYBQo+wVPTDCpgfeBa4CXbb8R7JyDy702vVrEG4qVVTxnnkgY4Kh
vKSTVLAdpChINqCuDP0AomTWHDFgQiM2T5/kLnxqGx8Oo0mc8DfBza5R8Epp
UDDkCQ9TUtOp9BOZgdl05Q95O6bsmP+4i4+4TE7NXjOnNe6F3mfMQJZ7RQjm
/XTGbCHzOP01zNddRJF4mAwXpqzUlpu/dZS8jYhWdqHODj05I/IPXJplLbFI
mai/9kA2oucZY6mrc7tfsiXNQ/1i/ejbIVFV5UQrbuiFh2pk/eIhOxOMpiMG
DdjqXmHLgZKyRej6qYEIi/kMEmajx/SA1AqUbQYBUI6EIHS5/XO50I8NkisT
s/a13/Yfa8YDgai8grvcnXxmwKIPzxWY7wCwSstPCCNLVPC4DyorZuybjNLs
3XjrJKj0WESDpps9BKUB1u+9iP/p8UuwFFW4pzy/gdHPbCxQLlvfrHJPbNbA
MXY0Za0zBcE4fLahH9UHgnWMNzSXY6jAu1JNsd/+2gKRk50EEd19WyTOAzYf
4DaXzgc9htFxwQ57EJO5eZwPnv2HWsn1ydHWJZY9mVSRihn9KZfeCi2DHkzl
+TwRw/rRESBbjBLdblhjTrbsxlLEcxK7bQy0Gaxq8iZt4I/a0lG7vKTSPgJH
4ENUInjKRXdyCaGPLcpyIEV70fiz3CVC5Ijl+gZNll2wDl7iI0ojypduOUQq
52Wlg4GV/uHBksweTGLdxb0IYxzqzylSg8u3LbVIpOMQ9JmgPEzAmHWA6+49
dJddIb7npPsJI9JPg/w34mCTCAfb9gsF+njJJBLpJv8VxrO5nTaeaR/cH3Ty
khh4P0Sj+N5EpE1F2v+vVothTmsRM0CZ8+a/MM38ZZj6qGuggtUMA41OgA2o
e66MitHe5DDJ8B/Jl3ddSBx0xgkwrBem2yDQpQG/0TXTf1BCk9TaElUMUE6y
xj0NslKXw2e4wvjwBTraJNr8AFaIau2FW6KEYszqm8T9EjQDI5wZ0R6p46Zk
EJ04/4eIaT8ub3zEXTO2WCNSq7Garrr+Dv+RpkAxfsBjnWGOWYnnk5zb+R8D
VEjw9qYLUuBRcQ8uq7muxSWTtCKPQ9sLcSm9jQgjv2r+iR1cnel2hpog2n5o
nbcrK5pWXe5qLfUEQdD7vIebZy5vjbWPlvueQXVefbGeyhff9Ynm8FNal3ei
yNrYMvsp5K/lAH9eRGF1DPAKhHu4yhgk2PYFuNvqAmVzxWrB8D4zDc/CsN64
eD6MxtZw3fvaRwk186HB81hpOVq6gNeyzEd+rCdM/lkBxgtxFJmWP/QRcACz
RopuqUl9Ofpdop9xaCPIkBUMY2ITM1OPU3ohZMf4SwXKptrzdOsCemjoiyF/
vW+BOs2KzIgdGJrqyYkLykkxdwoltZD54NtVZqN5O0HDeKGJs1KVGHbGldUe
SwIcgbWu63qr81blnnTh1gdIF54JF8gBJMjWUuIiha+5qScsuENB+wmvzkJx
NCaMoha0g+0nTb2sYLi9simYbbqlG1+GG+PncDFX8210V6vtoe+5TW8LYemg
AnL09sT+Gxp2zjSwax8owMY1OkLf2xH96sLPylGi8zlWNKqSIg1ezoSJaiy2
7IzWqzW20UxWzmXdrj2hFuZOECf5l5+oI0EcfSOjJJuK2oEsbgbM4JJu4RBI
Q0Ar7wVSulsZZhDO8kJykXTu0k4ixUabNGA8Ofk2TkDVSAXGDZUKP7HQLEBk
HbU97GS0xDySQO3OaycIQjbn35+GMa95d7lwC6+69DHK2ZLt7CL9NCudDmsb
yedSHX/NgTtIhMCCSVgmTIMYOB+gUaUESGROd9Vcpw0y5ZKEI5LkC2P9+58F
jv6mNk79AxmeuEIYHb9y6/RXvX4ci+M3iFD/eVBKUNHJTtI3M3VZtDcEYbsI
38BXygzXoRg67Cy3Gpppkp+PTWT2+IPEzlfpZwoQhFydA7fRv3ufGKCoMxFH
17+b38vHqVrMmhjnnsByaGu+U3WpUHE4/yt4bTcnCGH7Y1NjIhsf3ArP0pSu
y6tnx2z8NFArSL0MeL/gsHtMmACzWfX0jFxjH08MHVCTsUvZ8TSnter1oHO1
W/n3HJY+NZ+4qUibmXzDL9wLZKd2wPQlyUfT/BRhITOlb+oZRMjBtocEwtB6
+waxwGSsA7PilVM0kZSiclLc2QY+UtSNann/iGNHT6JVdS8ERK8SftbFnSMu
vrIV7282bsSvPUWCHIVfc+VHma7/pQyvmoc7yo4/t+Re2b09zpw3dfe8b33K
N/nR8CDFRDGRkKnbfJ0SUftXvikASLievWww69Twdm2M+HgIaIIbTXc6AKa2
ANc4qqcNKlV2NyhqosKjqwpS2GB9D7UbMGlQH7Yp+8RcIIbrZDbxFm1lyavB
ZZvYwaQRK140ByTMaEGjwQlusK2f+Dh6Q0upy661yvhbvjDVe79ZesEHZ56m
X8SisnlnVXJnx6ieHaqCsnZqBPzr7C6XdjkvY3RRsrux10PkHooASmx1ZfPN
6vr9QHRLrDukzdNGy7GygvDs7QNyZbdBrx5bfEqXLjedl8jruSUu/dfwocQ4
gEawtWMu0Xzmt6p4xtp/obR7RFE9987xgrF5OFHKFuBmdcT5PLV9j9GOEhPA
gmBZxs0WSC+m27TRBIGdzwWATZ5c1V2kSOC8DU2Iv7CEQG0tIcr89LbNOgQz
eOqJkm824m65XVHNeL9TQW4P5MlNn8vXSfuulU8fzyi3ZNBySIjHEv2U5mq7
lhMkY55szw9ruKlyBc4+XT7zybC0SRF6zipAG76OtFwUCqD/ll8et0g8bcjt
ASPcI493pHPtaOr98RGqj1sHZoCGrh/RQ8m3fR5nMxAmJNII60ZoTXsPpljY
calfQXQ+9w7wZP6/kqrgS6eBVT9c0npUElcHz46NER7nJnakY1tcY91l3jxl
KyiceiMMrzz6t3+ziPA+o0lHZf/bXPti+9jY2wxZSxf7Qq40k+6dqS1MLxv3
ZLOypGBJ13nA/4/OxvdaOw/cFa4CMt6DV5D3DOztTM1FMCCNheXViWDfc8cf
wJ5pMECv9QbCWuSl8ha0b/EPN2HiU717qlcviFhSl0O1KTvlIuQMjrBveHmf
kFcda2kWKo2JGlhOhnlh84f8KA29QR38apmsINf91TUQeutuESbaCn7CVlT/
W3NFZk3X02D45vj/FOmZALvaQZkxo8xu22Z5wrdcgP7HE3uGIc1m2dnCImNs
P4GLMzdq25NTT9G4VliRLeviBJYA7a0ck5of1H2ZZik92IwuGnltaPRBb/Gj
d3XovNJkeN8IJYhNWL/TzBMeDA/jNMPtsaYtbb1rwjuMQv7ode8Xp33OS6cq
UNxiuBfIeu5HJj8slWv8eVE3NqzYUxB6+NTfjO8K1CqkFe7fkgyj47pQdQf2
PJV2+w93qq2gbk5ApBya43yqFBFzylXxqhKDc3w7giV19t36S/yXUA3uPHEQ
D/C6iwnzzjiy46PFoP+mubB9rhMt60OvRJWTQenflbb8d0Jb3P35/89crqsj
2vXEvd4q5zRKGmByBcLjpk3FQlxmMcImx7E+pkOHY825CU2ud/XTy2VoAqbY
QismvIqf05zJ5Lt8zMJc94u1f7QwR2mm9eiDxyfVjAoOZ5aG9wRF/AQWw02L
wfndUrTH0KBzUYwBkylIKgd7/AanCFRkOpG8ZP4OgNfRTxz2OIdfrtegwcJS
KCWE/GkHzjbK6fJAwgoEVCv3QSqCl4gox2KFouFrok4npMF27MPRUGGeqGFb
lJ4dTCPnOX1cTvYWQjFkHLTUbh9raZ01TTVN+h8WmV7tN2xYaK6LLaQJRoaN
3E8FE0m4pobBpSkppexim1+uSxOxC+5Yghy/ZLSzbhwxMV3pHehKrS0mio8L
elAZt/ApVUMa/DRjhBMcRTJYNIexZh8Aw/fkN3XTYF0D3SoV4zO9jcsoxgxY
J/oknTSqHrirUq/t+E5jO6EFaOrO77HNcjkRRKDrXk8so+0BkW/kRnQFi7wv
O6h/J9iZD+CyMunekqMPQLIr0HAMTUSAqvSvuaI1U88uEf2fQD7wVD87xZ/7
g6YilQPqA5DajSsUru/OlX9V9JP9FPwmc4aBW1aG3ik5vISxm8eNFey9LUdp
7pOyNPr2IAPtN8f1g4xqdqeVBtDgt7Gf1f8C65uaw9EuJX5Jjkhl2/Qgd/HP
gd/eDjy8j1Jsp5uz4wro26U732/lJErdF+ihGNjYnUazk2yWTnb3eAWY3auk
uUnwdJbdf38J604g1Kpp3XjkwOlqugCV+LtSZKvnwSRDE4F2DxAzpttJu3i3
RqHNcBZZtgF95f/UqLHAvKcP/Xvv6j9eWwgfPD0lFdIOw8sbTGLdvFImT0t/
EEaL8yJMbEDuhHi/HuI3k7ZVDKfF1nUyBJblNrBO0sDju9WfkbGy17quFZGe
AkTXVgKXitj+QGIWNu3bni+2qjXw9lQGLMgwCiWLEdjTrl18kr3NKbBBwSmz
BeIHGUxS8vuoutTLwUwAn3nzBuP8vV6acAr8lvWp7jrgJwbAVfQdBZ3Ad+oI
zxF7dqZWQZVYezGR8Ywt4vdVQmRPWmLDRT3kipE8tfoDIM11TsG2rBHie5OG
W62pGm3VbBQZctfK4JV5X2IV3g+ZMAUNrlo7zpk+HbRB8PzC51/IT8rehyK/
WEZIwXtj3wc7f2Ngjaaxttnhc/KT+WSwPZd7pW7kokt5d8IHZo5bt3GfPijg
xAKGk9+R95ybgsl3xU9pjN/Log2W0H+Sv6N24OHuk1sOqAcb3w0Fp5aQ3pS1
cmCLmsp50fcSPzb8hRsW7vxCOx9L5edghZcLH9rxQeKUrNjmJ18CfjbHEVmZ
8QZQeIf2XaZZuOpl62pnH+0IxTVfiMwUffWTrhFuokakv7h6dQ/fo1DTERY0
MvVkaR6CdMBTz6bkkIfUqA6ZDG1lKeiwjrm4IfBHCh8vtLTijqs72rIaUM9D
za6zo4ic3eSjIZix1T9DF+/QGhfeDE8iGQtq9JXH+VKx2B7On+hSD1PAIThu
YjUeUdOL3iJ6Ccn9dhbcRF2Gx+nvZIsxy58M8N/7YRQCTfSL+MFJ3cXGjP97
4sGup66V+VJlvcHEHzDZQ7aR18D5HTywUYP5pjX2h00FrKmUKinEa9rIYaYm
Qxi1Wxk8nvQFR3YPtLeo9jF+gvqFxMNVHiq+iK6BUQZmWUPj2Li8BChL9jHo
lvmQRscdlp9Ngxnx/iLtkmTqvssVZ+MSZKVAaqM6hooeAnjKjz+B1xLek8ye
nHOaHj1n1YBsW/72Np61NL8GHZd52gJEUIImsUKMz1TAbsUvkHGNhCyiaHyT
umiO7FOEQyqqpU5/EoCNW/o0u0A+9IbaMUJ+H/f+Jz0Fp1mURrHLnH7fq4YR
nwH0SbKYUOoc3rtx5ZBG3nHsSeRRe4/JBPdIpVusdspWGdwVH1jV5X9Al218
+2TLBQcG3Jv4ZKr93OTGEGqI3Lp02TOaMApDsDAgkbIbyxFCJBvExjkFwGUv
yFtBBW+dMzGnUM6DXKm6K3I8r30rjF1bYog0KyKgLtiSQ7KlPdV4/G12rhui
ycp8OiBeIvFG5asc9hreAKNuZ3JmyMr8ck7nHOl4Vw6sK6GXIc5BCmEX3YzY
WCTojfodsNuL7fgo5sfgAP3t/oEecI/i29zFZKzHWuIdZGSossNBTD7N4LZ/
YYx6pbtM77c5L8EGXiTLgeBXTmJYLtqNrh5mAvEUQIrd8yjd2Ef1bHk7NYO1
1K0w2yRsb7pLnYTNs+FFsZ3tcXD69HkBpwicM8ryMTFRFN3R17+Z5S3pvGqG
aiII2rtgr3r319VyVNmrrMrpG8qFkLZaXDhvSspDU3cosuJA5/bmhJCGHx5H
vl1YcVdFEF7n6DSTWRXizfRKerzafNytquEp2YqNbuYGza8jlzpxvUus2uGx
qNj2Sqz5PzFcz62Ovc3G8TNZnbCT8si+oC5dk/G1i0T8Z9hLLu78B0/FGCXJ
pffBQQyzgnIbzsQAnWuZBoH4/P1P0eYExcq+hhWSKADliKH0o8rLd9qglbkv
cC0x6WPkRL+vdBSsB0XOER5ux4XED9HQeRGAc4zIn7A6Z0GXELpfzllKiXx1
pC5Cn+QJHkkbVSExB3qpbrJtRipL/87cxOyOUSs8KsmPwPHfKnRNn4bH6MgH
6tXkrSv/2UMnbVdUwtcRRRdL/6d/8hrn5MMkwSTrLSuabC858cwozpd1+VVp
EaaOKzsiK4Erbg9ZMvwY2cSQFIsfZW0Q1BYF7MNX9O+u71v+vbj5cmD4Bd9V
fwjQhRAv1iy7jYFDZo6HJmCuSr5yyXMxPIAN88duy2Q5j8oSZHeghegKKSit
N8IRhDji3jZlkJU3Ox4ZB7Z72t8ZkWGYj2JxvqsacFyWe4U2DaMKnG5WHP1t
1qFWy8kMGSAifyCipdRwqhlZCF69hx+R0onxyNyBDE4TVwmalWDxUekQrgus
ItwoboylxF7LFI/LjK2OJ56eIOO/ww25tU5YaCOgmEdsGwIpAghCXv7qt5nu
Lf0phAOhWYm9WqNZxKcw9wn0AE1iiyksxNt17IuR9APBIYa4z1RRJPQc/y8t
HMsMWRKV/75S0RUPFVp0kxVdB8jDt+rq8f57Xg7tLKkDOXzXFByJz8shtT5G
iRM51UcgrdbYXyzS4UvEDGKjz87/pfnyzyN6hAtQnonEzkRhaXaELu8Y3/aq
2QVzfNJt2fmlP2/Rft4puxkt0Y/qF29fqOe3CVVT66crZj/VfIPRDuutOSQW
7FgtlB5LU8oKM/fAPlDuU5FzKad0EcjLCphq5RG88C928eKkSGxkIt+TdIRX
+TDU8utOXtGSJUyd0ustQdy2TJt9WyEAdOKMyauPDHjb2e63Sn52WX/2AS/V
U2KnwSWJxby/BRomT2ic35dav/oWb3m0f88slKQ5+9UGUf4y0aaVC3W+CPO4
kRQNmCQk/MSE00SFRfeYKtI07z9KRSyc+xk07PWUTy9ARu+fqCjgbLG6aK5z
Rf6mDOsM3q3a525/WxOP30lXjmFPh35eXpRnH8Dim/P+ID0kjNuYvp/AtY1a
t839NjZsKm2mrpuP6TilzjZhWZtKgzYNNg7JvwrMHh24GLQtQXMqKt7kQNTM
38/jHxRlBG4qpJ8H6hBNQCvBk1oOeoqPB0scI5EMg/KF3B/a1QSKOXOH0agc
emeVQwL0hVqIY0MLk/vwj4p4kOojk6uRQEdziQNDnQRWaPu83C0mAZtk2p88
wNuaFz6khJYP/d5IucEkpmq4I7t38NYVwqQnMR7UUBukwMBRqzXXjjruUIVT
aydSODTYIBizIBWCwcCZGpJ76qfVYjx9xze51DlvoIvcNe4cFd2FKUHl33TK
D5Ts4rKwTO+2ogAj8UYZ+PxeSFS7+A7OEN+Dk9tulFXYSBE86L9lJnXgC40m
dtun1WcPKxFkWvrDcl71iKEMYWsGHdhmoWJRjCuOyzKjDOxwONH86c8G2JtG
TIWMqGfZTQ4SZ0zuLrlFym0UHqvpXT26VYwrKqMoC+KIzcM9fL/l/KtkfCbw
tRfgVH1kvwVE9dKQWyz3LpRCKNcvi30SOKLVGqBa0cxDRGfAODhUy+Q7jepB
2o1d9eKHpVDjw+u0mmfORoxU1mYnXabI/9mcTwi8mB2Z823uhwR2aPakVj4e
smJDlsmRBGdNEYxI8bM3HrHbMXsUcgCDsMZCQnMXrlv5qjwmra34pE6cx9BM
mrVhDq3aeXg5iFbNmIL3fD3uLYRoysWDWb8+Jy5u6GyUDx50rOP2DT5ze+kT
LEwYEd20AmVYdraIbE2rYoUKxSaIC+b3r7iYPJNOcgLpi10PL6X7aaDYmtFw
wt58yH27hRQgRT2MBYHTEDUlzpA7uGja62YWJTWSn60BMpMBeq59lWFljj4P
1C51GmxPSu0nu0ADAjv1jaoRT91TJqeshyUXp0RdorAexfoPJBlG4HsoSLNN
4OR5aCUmw7ijlHL8eAcTIi153W6TOqLx5VychA4uq7ZP5A2Liu9gnE7PjfWq
ingbuTyTHEjHuG2vezOBgYoJtZSL5TykVREFguIk4//1xSyvxUwBFgN50+x2
pXtrQRjqT7b3sexfFCI0Oda0KeG6P0OgfPOG54LQ8cUuPh9Kf+OHajCOmGL0
aLyXlL6gVoFG6acTC76J6uzVl31mXHa5APAfegcZDZacmAxaxYNFRhjjQ+or
Ce+igG7UFSHUKJ0dDfeBxyLFDp2H+2fo9IOa6eSsX2SQkTNL8ANnVkw+qALB
g4QfQgl1jn7CnEZw6NdcD3QSBct8jjbXsffdEQcI+zXSumddb9xiQsLKXSku
820WmK0Z2ck0JY4rMXjgG2UtyF0YNVtI5SgjofvC+eHEHKNZuLPk0o3tPMWA
zx0u3HY6kw4kVsmNmBHkXrl/JLVamQB115dPWjGXrlv29D+oySHUK29yCu9g
JHAykHesYZ6E1kavFE7FK+yKNA+TsltoK7O6L8uTHpqyak5OkiDqZ0bU469z
F09YTXcv6mSyyuSGShYw/7PiuuMVmjijVm+vA7sf+WiF3AfsgZw9XaTEYAB2
ZiDphNIqZWEWNPG+heGVEj5OkyRdTbogTlZnYjMlN2AXrNykvuLOc+8gAHJl
xJvtKm03VO2D7Jkc2pkKw6yqusq5nmaW1tV7EksrawOXozLy2qr5y780aaI5
IYkVsl8znUTx4h/zpP6oBwd4q3D1lhnJm0i+VIGP3x+toS1Qn4EuhnyAXgDX
dm5yu2qEiqO7V214bgUwdPa1dk/Y64fFP0Xw1k3db7vXVoHgohiLyUNtQ2DL
7mLezORVAnvgYhzQZ//8NIowFoB2D+QFstZ9+8n0Ce6ktybc/Iq6jOwHmppo
XD5tVjIF+7LrWn4Vy3iWFV+0WzgNR9Jz3opG0SAy8wAQRWIFjDwsF4AU/uGU
snzH3BJmmXxNHrAusjclYbeFqASfaWUOm0mUvn/kHQhc4lokd3HhZMDbSumu
apDuC1nlaPPqCoPz12KboB7PGZhBORy8rIASXF0EkcDLqsQeUeZ4ChlXuPLJ
SaHqwZ5sQsUBTydDucx8d9qHBhRtpjt9nYoFGCGMDp5u+Pv0J9/s2Q1kP/99
b+NZCSdt6YZR4bKTd3/3Exww2Co2GJT5+UrhUxDnC1PYY3qNkXwd7yBM0ue8
I6mGVxCtlZYra8uKpggcw5WxnD6F1mlTYJSr9YHpuskHwnegOTUo8TNDkZW6
QD8FE/lgOdOOFvA2go6YWZxNwtd+U0oJ3yztjM/WGGKc0HWviV7BAV+6Lz/0
JSI0m2+7iKX42U0TeY2YZMDRI2Tq/p8h4E5uwdIgC4u+V6Xti8703tzBjAmL
WDIZ7JuQ5sayKMigG9RByO16hqGdkCZAU0Fudvb2YPhak0DZd++7re1Ok8bQ
yl41TkDM8zdSEaEOPGQf+t47GhpRXz3uzR+kx5s6SPpEII5RlZ4DQM72UnpJ
5I5uY+OiPJcrhg6Hh8/6l2MBjdp9ch4aEaVjMNAHDJ5VYOSTzpgKz8nmeBV5
m+npSL7ZNVDf0x6SFjGti9bxuVaLblT/AdRnF6iY3Lu4whFQ0TaYCSbZDhyC
ipLHFfetPCKesZpBHI+8y1BsyRXew4zYEujXYx2kft2DscI+a2lLiEN2o6Pw
yqTGF5rXChhkMAyGBeN8pyqqEX4vcmhoxh1oqqryGtAxvhZ3bVG85LdJo6Ec
RQVWqZ696lpuLtc86FJ0ZpvJQuT1sv3Fbv/rGnqdjyKbVYSHY73/yY6CtYfE
LCq/ua7kPe5KgV+mba4f1BePYR6LxekaV4S7a48S+ZMDSfQu6x+LSLtUuGvS
2+98F7K0zza70//C0lmEL6spI28Mi0NVBoadUnM8WoQTq3AqusBW8ELaQafl
bru+P7SIeh6ibZor3FqL5vTDJ+15ZHZNpvC8qdhM3XufeJSk6hsWhCx6qSdt
bhswJqkQ/ZRhrVdXEMl7zMIBddKQA3pqU2hdyCLBysrxdFOZzh6BFO08g5et
8/R6Xr3Y1WqPwOrTcnBAiuhJozXDxl2hTz0UdP0/IvMi5wGXeWf7uKHoCnf8
eHhcdNStFx0de46Jfw7SlkLY1w8TDh8WwrzEzKW9QRtJPVXZ7BTfxe8TBgHN
0rHwuGLadEB9mhocxyT2MdWTm9KAP4WAV570loqumpBAFWPeeln1L4rnKwAZ
B2j8AKgRncgNonVNvrJSCX7y7zSDVWsneGKtegcCEQ8+fkIZIejx9LTL9Onr
Sx1xUZL7jB0PtvjRuMWLwrScfUN4esJrVnEuanK2+R/PB6ameSV8QgnRuM82
md7RALlf0brxUN8ajY6E+pnbnWZm1qva1IuEZ9Jysm8I/pG4E4Bw12lTqkwC
CpMsAJG8aSjcVasAwc/MMwRdl4FEimssY+iUDearE2xMYoOVH335Wb7L1Cir
7Uy4F6/cOWVbm4i2ZPDu13nk1QSRIkB6nRCMoq7WUElr8lehuMnOxKJJM1k7
WBMzedtKun+hAvegg/8EgRSks8Gnoj2Q1EDGfsro9zJVvPME72A5VIW3hRcl
UGs/Pp1+KGMYSzANv4kAVN2jnGJxdNIPUxXeeKQIx+Hym6PWgiCLbYoaDjNv
K2YJq5bI/oCINm7zUINIUx7yV7qcIT6fZfZbVCHGnZNMzVUcHfH1PwHlP+YK
UKXRMnAR3RHgfZcrJm3d/krDl43eU61DcI3BclXDbmDSUl51M3D6Ke9j5rJT
wjR34toU7O/TJFbKPo5TxZ7LbEDhbRPNiOcDw/wJemmbQD10rU1zD1QppiI0
9f3wsTKcaI0jdrLTczgN6oBqZvftcAmjPaEEQmG/CL7qyBpTMW6w7sEkUzRE
gmbayaSMtq+F94HC8ZEABVhDCBG0zd4sm5bVXurBDNxCnarT/SDJE29Ol7at
pSy3S9DWnIE8orG/IyHp6WD7M0q1sI1DbDfI7GU1mKba6vSw7t40mn7CEba1
NcnJfgNWrcyO3Iy0COHj95nPUKNSBRHPvjrnjWWLjnw//PBkOFYb7XMFBjKV
2IpjAeu5QA9xCaChrvX+726brI3/PtTxVO+TZW2emY71Isj5ApriBycq9XU1
C6hOr9AqLps+ljCxfGnk5r89YZseC04TF3apg9W7Ai9drn98t64vaPHEPASd
KtqRv5c2Cav4ztHFP2omD5xDLSRz7pHirf0WYri2N+Xxu97qmx2k4VP9Bjba
v41Y8HvHxDVHXCS+7lJk/FLaMVCb0LWtDffLD9LpP3G4budDMNhK7Kv4LLoT
obaOJ5oEZqpKZzOxiXFW30VtZ2ednrhrwAHFmkVwexSU5Ej/cQ8DcViIE+O6
xTE2WJF4kwe+/QPuU2xf1iT6TratlRrk5JRgydFrInBbWB4RuVxFyIUVMM6d
v+AFDnrQWzfz9V5UqBvthfnO0TbUDGx8DMg8mnluFC9z7d4hdzCSmJiuIhVG
py8RiTycrEvjZgxRTWGiDRyqSChbgjP4PIob/a+jiI36Sew27YDvag252YNN
mbES0doNwt7ruhzeYGevCwYV0n2CmMyd7heibPgO4hw9czKe+ew14VNIMyd0
6zk9A68eARbsHmrrPH1h+8ucCHnAtINyaHLdoqJcBbwr08ZOUoyiY8Ieu70q
Wea/hHjhydHoQaaQOmLjFYGQLtpJlNmeI8A+dSk5jrM+7DvaiGpsT4x0zEs2
g0wo6yfLxEsyr7MLcnNOYrmrpVXGThvWuZvjAfhU3jAHcsypGqaLhEycS3L5
A1kJDwbc05W5JXNfRsypFz6XeM9VTQ1QwNf9doyiiXaQX/PNp6e03UjWRlNd
G+TqsKwLam08io88A4d8v/9UVK3i/bqlYdCWRvtJDyUlweY5uu5zbVa5ENgl
IDqfm6fBl+339qH4iEQU64pPpiP8Re9RfCBYgvr+88Q5kMY0NCigtwkVrz49
vhcWBFwsgf5nATI6kQbHOi2lyq+AU5IiJAEjHPzWuWuGehga9xYExAP5JoFn
lSSe092PJQIhkwF4xBincBdfioL+tNiNU34dg81p1EF0jUlHw+wxxO4OnGB7
WNBwZcHfo7Q7s47d2xlWoIn0qDh5Bf4S9zUYqRb4yl559pdUdNa8ozxV3nnn
0pP3ch4LzW8VJgtpDme/LDl3UlKqHmc0Kpoh1r/HFcZuOzqZuk1yZMgLYs7/
TgYOpNYMsh+hKVmQdrzmcXt8+d61qXWad1F0wsB+j0MOlZATRofiJxDDWhCz
cOvCu0JVmOvFOKsThHARYbI9UKBiN6cunlCw98IqsuLNHSpoQhctTw10A89k
g1BaCDr2s4M0SwN0sy14Wf1IM0PcAeeYDpCKVX4CRww5PDZ6SqfpDFijhphT
hG0iTtyrQ3OK4eFMO1drKOWm4F6WfHse6Uw1629YX3Qxt2NNIwAsEpZnfh0v
ZxKRnEhe6jNqXvoaeI68kpOKhjmTKtuFpfmvlsmjW2vbFfqrp+sxOLTsaqkg
ZtxEH4OIK9zT5DMhDIZ56p7vq9YUDzcGPUUM/FCfCLzgypJ0w5rSH4YtGLxS
1TPq7G+hCPUpJLO+Iz1gVbfShRaIpRM9WyPPwV/rk8MHhDLgM8EAiRNuhX7p
qckWto2TVKY/NNka+Vpz2hQd76Hyl29NcS7YC/95fgR70qrei0xEY5Ury2zY
k5lmoYZmwBPCiXq03ue/S/uwkxGaLyQBGwBFjZ5wJO4Msd9xcP2xrN6vA2zu
BAUgxXy6nTnZ9NHk59TZN7mPDS/uWbw1kRn/z4cwcLzDyoGpL23Ar7i/UDGw
KXqp4ptKAZud4YmgkdoFT2Ga/bS3hHEOI1mh5Ce5d3XyuBZPVVM5Ez1Hogsd
yzQmFNWmSg+rA4QEdS/JuLJGa+WGzgLcpM8twbZDvFwoKhsRrxz7qPeSY16d
TEaNLmtH1KYYQtW5IiCHdKdohtwoPVGOY9F1oWgIVOoD9Wn9RPeuZw2+u2Ls
xIk5BAbbS7/CBEc9e0Kqrv/bx0bqW/+J26S8mmMy/uWtGHKtnWkXx1uby8gM
bIx4i5RBAvopUW5dHXHB8cPT4VJLZJagyRNzWR9CJPaIZbnEne7eLgEvGa6r
Y7OgKrDD6exPEsqIf3bO74Gvohk90N0SiOs1bILB2JKU6ztJYfJ4SY1yzehv
WlPx7cfGN0XKasOy1PcgwaOY2HIPKN/Xd415B9UehgTzNhHjItaKoMnKBxeg
whj1lQke0GlRuUSLJhFq92TLYfmp68PbDLblMfWs21XtcYP9HTKleW8hwL5D
3cZ5O0Du9VURygJnuAIuwBsL+dl2nsSj+jZlzGvYA0NG3ywkfpTsxoXLDndO
8AEXOT04ZzvyZaAJ85v3SupDX3UDzC5gPnCjZinBQ5Cw1LaDnru0WK5RjRa4
Ivp9kfBtrCYw4I2JMnTa+n0z0Fnkx2tpF3wRuEorpO4HGyNNkWH9c7qCR420
mISHSukZUwhDmsq1TaAAKc9FWpemnGr9tD5DT1+rxM8TEPgXAEbaF5J9tMls
WAydvZzJvtGU4rj2zS5hMygBS+P0zw+DDbMBfkPDaR36S2DIxMx0zfKdT5ex
8tCiPoJ2PWzfB6jtwmfLkxsnQnxAc1Lem2djQiccpLezTQpFrv96/E93B5ln
qRVDxT+Ry93OnwkywtvaYfYdUGy67cLfdVPzmkAvmO4R25u8BVHntSW6ta4G
4LsOGVZzBQH1s9RlbnjkOL+XPRVKGghHL8tPGY9b/883kWZfJMAaJJ9OozHD
CyhvjrraRxuiwo+TUEcRCcWlZpcfiYaBAUdlmPFbh5ah/sXDMXv0ostryViw
R4LeI+qptTa5oVWn4xY8yC9Yjbk+gV5hRfkgLU7VXvbsiQSVaP7Ei9iTCCFp
7d9T0dLifRFEb78Nirp56js8/UqTFD8G5eZtABrh22rG1hTpi6oh8aF3ZZ5H
FXu7Wn8MjIalAb4WtqJYtPVVymQ4po1P2DhYT+xCLMaCgd5m8Z4d27SkzU/8
YMTDODmj8jMPzR468eTxt9yvWgfA71Z2gDX93sLr7zY+pPWp6RQcNqn8bP6R
WFeTuUzg3efj9fejJIT3gAWbTOOfKqnelFUijn1nbOhm7LYhlz+/x8EmGHXB
BaOlxVHEGF9d7m8I5Cff4NPdV6+eSnIPurY7jIR1cRyieslgduK9LOP2C10u
NALWPFtRaR03uujlBMxRuzWyLm1sH4den6ePwaRzwS6VcSz1FDEoZKM993ii
1jUxKJvQSuRtLBB+PCigZUCCJN2Wpb5O9p0QtmHfo0uOU9yKIaA5IQA0PWH9
vQVg8eZco20WhbWGFYDx1raFAVq5WJ71FnxHFQS4NZBQVYM4Z0MFNMtc8Gv6
xQNvAQ3U+Fjy7FUXMZCpImI2uv+jiCMn2t5aSVpKlANP8Oiw7gPy/lLyJ0Ew
826wIyES5zWvO7aL73EKaDLu+asYVZxQzi/JPt2mznUgs0OrTODH7FAQPB09
7ZmpiW5UXajZx85XAmdj7tSlZz+xhz1q3v2+Ax0XCPegI3jb/2rYw1nmqzd/
yh7D9L38AueVd4+qkeGZ9HsVLKs0E5V+9FU2KuMYEhNcZktke1pED8c8LS0K
wPrUl3+NsU6B43i5SYRGh3bDDD+eXv68gcAlStGK0TOl2HPpl1btX6V2iNKX
YrNwR6sQhDFcrDGVEvX8WOEQe3D/8ehz0WpXA6yAV+Hz08zPWIxy09ssjMqz
ozaZZFTg0zgiyFukdUYO4tUjJaohpQbnCUuodrEXu4n2bzErfnQPHs5bYm7D
bnuc5y1w5otxX4imzVyO4jMbn5S4DH5+icwltKiD5DtO1Jji+Y+XaX4iyWts
3nIHJ51MwXXg3KXqRWZUA2P5JsEO4W4Fp/gU3dRvyxZqE6yScjvswAUzWr+1
yMV7G16kB/LSV2J+bIofJPOOG9g0lHDcaExMo2c1J3+92SRmmWuy+YDGPxuN
nYG1Sq8QfwsXjcQnoJA8Q43Lnkk5vfdFSlgFapma7nfLhUYOox8Bdno0YBPT
babq3cQBv0+ARR67bvgiTGWSZozzkoD7Ob7Up6CBJIGrjFIYOqRpBprOnf5W
iZzx/FJvbD93V5vptMpWC1m7DWrfInggEXDE6CtuyuqDdcP6MXPot9AQQyhP
LwuE5OAh74O7g4GTFzHQz+INylta0vv04XdPPUF3KUtEF1+M2YihAYCl6yzw
31JOpH7KhrjeDfcIPIOSsIf1FUehb35B6CE/o7ocwbrdKPs0GpUQjVGgAJ2D
HpZ4EW36JhTvJLkVjZjlPV4iDKJMs4qZqlU9a5+4Z4s61oct6sUNPFZjJ1Sk
AJXzdLJ191W64+2W49dfjVbmPZZVC86pUMmbhA6erZsRDAK14ojxrYNNqwTs
Gr9My4TSRioqJX1BB0CWdHGJnQ5rOsYN+Xut178G7c3cuYdUngsiLxK8cQj7
ZyMnNB7RY49kQLQjDO6QMhe38zhm5itQ9gBV/q/p5Sjcp47CkLdD+BCty1rI
8N9pkp2CFGHYVxVtC8WbAiWVJXf5MObcXCzXYLIYRIYVZ+yOjR0PptGEsPGL
csSqW1qKpB7ub0Ym8nXgAcjx0Ah/yLOhf8YTVnOJp3RiBUNPCr/ge2aJ31tD
4+ISnk6GfDmq5GY+P17j2dZOtHGxT3tG9+SbRhh5DUjG4jwl1CyVACuM+NKW
o1FvjVAD712321aQrE1J77fLDfDjPDtxUZPL8khIJNO5FUbTHVzbsWeHvX1n
pSQAAXNMlnpeQtqk6TkWDY9POUrm0AHZyMZWEspohiVU/2jrBir9w/9BRK5z
N5jZmBbNZD33DmHK6wNO1mPi1fu/vWEXua76u1mWIARfvibYpiQBWzkbD2IX
Q3IfizoQ2+5YQ0Sx0s6839NoOcWPPqquxAaBCAJwJ2lKFbI/rF8Wno/fjrFs
kWqhOjmuPCLPJfdwOFSq9Iv9OpR9YgxaCfTZm1LHn/m7hgQFwA7U2jQ9CCMQ
ADWRRwOHr3AgN15vzDZmR9LcxCC4T5VWWtfLQsfd+CWUBt2/lTqHhLeE5BWo
E3rrzuNACZliOz5qFkv+SmqAhTEPSKrYQagFpJhIpFLhuj0guofsWIwrgA6P
BIh1HZ37tY18jndTeJjhabxR2Xjoz7AETd3WkOyUAYTVaHPyPYSavi4za00/
xc+BEe5izcf8Ps0/o1kjJGsoaxSoBMVIiwm5T2+UyguEOaiAkALfBT+3EXMv
f4BTL55BZrm7DQv0/j+budnwzbnVSfknuy1rB9L4OyE9fk7E88VX8uFCWlaL
X0k75QUOVUt4KGGCKe+x9r+UbnAgEH3diQyJreDUtLJNMs5luger2zEatUfN
+CkCK0Ni4szJs/bQNnAIarm/xo93bHLJ/FwCWiutRVko5ir/Yk8k2W0Kdk/Q
BDJvFNZ60QOYw9taVfHcrleb7DxVB2PmR9Y39vACMRjlII7bq3lZbHTRgwdb
VVfwV9pp54M159g38j+zVrwpxGDbIEaQOYYzQQZZpgjYE15jZ/owqaKcHYlI
dBQZQ5p7CSTxhaQ11AZuv5fyt+8eBxJfZNIeCIQmL7vb2dmVGU6INViaxF1Z
oxGhp2KH71kwJhk4CyX3Oigvv0rtIf9iIPOdznWJ8c+k/VDukLFptlr7y5fn
BSQTw9+6wxuIV8+W9PM/ZcrZWFPX/ROXr3Sv7nQv987UoChOKFs6N+j4bdK2
D7Oet6flhd6zNC+2v6UU2QBjNSpQpv1+xEyOJDussOpg3+MM6oU81q0Jnshd
OZmgEG8qOr6QjYDlz26YgDzfvi0tgflx7HQBGvLufgi4hMSPgqGHi7eta7MI
eefl2jQItYhQM3mA/6L9cCb3dz9j4+3vlHlTrVnpaQHL3pG9cTz+Z6D6DVKL
w0mnmUe1ltoORQ8VuAlfWqBTTwIy5PoNKoBrZHTCWwR7RrQqKdBbu46cx6GT
KA3ZThDK1NyWrydtzqX1p9d6tOhp8rOjk6zspBxMS6jxLJCDKAKuv+zH8FEx
7UF/IAthVYzaShxy6Ps8BQP2Wt4mrGD9vbuoijHqEx6crIl2xAJLQq3rW8y/
SAkXKnEEc/fv/5/fzIGLyoJfnJKP56kZLVp30qbAdsHNlQgHlYZ9MtDBF7m+
tokGu+fVHRhmVvHgrp+fLJZDnnvZIhXkI6680fuqHwCdsYTNm9KLS0vbzWFw
6XYd/e3l13vIsjcIVUT0B4McVswVXl0H0jeN9FEtlRLTiGKXRPIdWLpCX7Qn
ah6dBFQAtDaQNaWHElgES5h7jOXffr5W6AsRQIInFdPF3xqtQZbXZWo5CVZJ
7HAQnMPV5dJf6kImx088DssujnknSBu7BtZk5r6ak8HmECQT+L6dnaEpALRl
PXlZpdt4AzoisFkA5nO+hNlaQJuWvlflG3F2zIqt2CiObKvwFeW2Ygk+OBWt
9FNzuw3jkfS5JVaOUHuQO34l5T9jG+0NDdr0hmXtk5dKcJV77uTXaJ1rFv1l
hOegznj72Uha98+mFataGFucEUXjJ378EhiO5JXGNbldDrXflKTEG3fhBvHQ
wKmjPs8OJAgKB9c6SkiuJm0AF5AQmVKiZ+8Z64wPkBLXi64Ui+WtTZ/AYTNl
cj4toNGqBqMRNkkAY0Q3wW23jMfJ6LqhqmfriB9oYnBk+lOnwMXrhHwVQJ5U
wB4THy0Avz+xDe2PINqE/DTKu5yubrOKTR3yN983z9AOOQOExtTOP8yLeQpC
0SJFoq7XzViE01xW2hswE7o4l2v1qGBLas3L2Hgbdj2/ayOlM9BqC3Xjtz83
vFrEJM5OMKCrfcnyS0+8J6w4m03dtgUc8z10Ea9+U2s/QZRixJzfcTdDailE
/4QTgeJPinBDrgoFwE8KNBv4GQgzAXc2TF7w4avhHKfU1H8yXPmrvB0bYEPc
yHYpq00+H8T08vwMzTbD7CuYLu2MRL6gWKCdP3RynrO3P0JOlG/wG5dLYSl1
7A21O86C4+7PT7MqOz4yODwofwyLnkUPnuIWZ3sZVCAgAo6qStJ7B8Qxfg82
a6KoOUMarXrlDcf/EjtX45lDmB7HsP3Xypy7skL3pCW4tBBW8dJzR1Kki9RI
CAEmsHkiIOq5nLCcvSqWLCSvc76unAGvrIzifLhXTuR2N6cCpEIbTRW2NfM6
AQDXHbznteq+fiZvF09MrjapTarPSd1ADPempcVT0Owp/9NmA1tAsoUkaI1f
gP/FwZgG3m0ov9PYHmQ8/ljsCOQWZjnUXa0Sdw7SRI26hwaKY9uAAGDN6eKx
DHFUHqRC2TUE52XZt2QXs8PfEULxXfLNR/OF2ssm6EHuahSnPRKdQw7FUKva
GdHAUxzm9/0qkdQ2ZYzY/GFEpKZ2dyJ1ZXTfCrfbT0NLmM5wzheUI4DcC8IM
uYfarXabLTSM1eFpm9VzWydRBmF+OcSBC21SG58zG34MzAcKibCb7uvzbpNi
HAMImx8RNDjVUjT/Rx6f4ZIABFWHQo2oJ00r4azutEUrWePg2y81FtECgDRL
PntV7cURhwz/RDzUR5a/ll9H031rTrYEAzIgRhfYD/pjE6ykN2P3QDHtaYms
44hNWNTPnBCtBi7lXQbredNJy36rVdJnBX/UbMBo9C7cN8fYeny03AnQ9zQa
s/7j4DmLKKKR0AUElatAV9a4lmPgo3e8cjGnvzRSIXEdK9FrOrgQOT96AhQD
bhuwDkhNoxN7mKy/6PGDwSA02psoq7Z2oPsmM1sjnvMh5/SAG5ic5YXKC9jS
tYfIuTfPXscXf3ybcz7spvXJLbvRx3r1hoSfX/mZSw6cHPZbQycm8b5dvC+q
k//ZpTDuD42hJaA7qdibD0r5+cvN12Qk9xpqqC1S8sGlDmjRJzoBf8mKdp3Y
cNel6ubTa3782L9eX9cZ4/gR72X3PLHiT94iHJTxxzFnlO9tFLMxStdPQfAD
+A0uNCvdC/aKsa8HT/ZscqNSSO3Nj9WBHJPAHpgt6WRcNiK4V0adgXgUZ7iH
+IlH67o/NA9kCN/j17NPE4fvB97/YjcZ9KZOfCAeoNeII+JIXSXoLmWqId06
OppXhqtXia7N2rvjlhxqGrRefUw9MzkCAuZugIiYEmOnEQ0X4rhY9QlJAAyd
cPNa0+d4s8ZaAanXhOAoHQEd+9eGuL3e97Hvjr9IuKF/beMp9/G3X+DC+XwB
sTDu5fQo0diBl8n2BVZcF2KGHWExKGDw0p+yZygS0EfwI6BOlQCvNKfEK5rE
eYh3DZhQrxURmiJKocrMspF/IT6OYzrIzzijTyLElew8B9VZ4P66PX/59ioW
F+bg8UUR89ekByHj3jvHkQMHvp+t0Nuq1Ce4XEJpNVmmiEZ0uOEU65TZsqYr
BWPTmPQhquR/HAYSv+4QzmmMJzWSwlPUAPlNmNcZ5pUxMtqdbzcF577zKFb/
9Ii1bE7C8fxU4U3ev+p3gg88/qdky6417inEXz/4ZOSKMfaZW4HhTcOM3qsU
JfwTAvNbqa4u4pVfKM51JpQ3OLOVlAC7N2BfFjYb3iR6bMshZouUtwHIzn0h
DkgYo0KqcWtc711i/JCHM1qlIT0yOkJ/XnREmc7XLzx/hCwWYtDPeQWemrNU
jZ/J7g+NTlu6nXpDFJazBfNKfU1Jn6zI7/u8NO7gbxNpwotJUH2oAK7iUWmL
1kRaXDbkYpsqAGbzP7Ygh5bIRPpORq88DRIFy1L8tPjHRaZQ+MmBxOg4h31g
hIIkrDXE2VtoMnpLAWdk5WW2DyzR2E0aqDB91X7snOwYpbWFfBIgGYxqzVT6
qRNtVcTiBbAXE6I62EV+Vs8mCepWSmMCxwoNgms3fzhAZrTyUwv1C9Glq/xn
TsaoWtrGAd0hybAnALEho28iFaLYP5fYCNKR6PF0J+HbR5tHpAMY5BVCSlkS
botmbcShnwqSp9AcnfAlh1CoXR0THcePF0WLXj96w2iaWtd0hB8SJeHZ63Ds
siye8CT3zJNLUZwJ6/4dG4D2JiSjsIPbuIZfyBSTtbDQfQU9HUDGE4XN/cOM
MfzEZJAf4BK5AyLcNb+dFE13VFD11UAICo2KJYB96oOHfoEwQpmgev7WEDeL
lJ0poM6wtbI86dxZ3p1FobcKeehyLPGnbbBpQcz4n2tzA4yBo5v0liD/v+sj
OkxmgaFHCUPUHz84WCaTu9Ds6t44pYAfadF1GcivvmNOsdbTiMcvnzYdT3th
Na0G/zZHBmikXtUGpeMoTkVlsSgs3XyHwFOjOsYrMsvBTIfIn9kW0cZQt0Gi
NfIfJJ7a4C4GP/ByxSSVjs8EqFsjbqB7HzLAHWvOLlduAYibfX1V06LIJzAT
MLy2Kfbvdh9yuAvZOKjJmkvHMwRFoNFV1kh3x1gccKHOSnXj30Ud3fpscgae
KR8RKTXTt/Geupd8O+3eRkkaFsT4FxfTbU3JPL+ffjLcWE5hHfd2R34VwnFX
nnmrVpXV4G1hmGpzC4ibq3SlVrJcT+eIEK9GOKeU7lPo5xO6hSSfWFCVKrzj
eYfIVI44uqr++W2P/Aa8uqk4W2jPdtxb45yc+/Vp7uOKkyn922idqR972Vtm
XAapdtfdDREUwws+7qsjfJEj88IGvE8Gk0jk6uwE+Kg4PqKtPoAm88X2KO4W
wdGr21iQL95ncPBiz/abwdZg8xnPfkKhvvB8ZQ3jc9UvU0UlTedr96SDUbXS
2W9TABinOEtjPupnWuh1T6akZXlqk3T1tg65i4l01B357Nt14L4oCS926rPb
wjd3MwYUbg/QmfHyaU53Wt2H/IEz7Y8WLJCkd2Va6tmuiInbNGjvQbywmzuf
euIqAEVzOeSseKb+fTHAuNBdKa/jo+XPUWMteVTsqvuHNvGNHhpdfrgshSpy
9xSR2Pj+Utn2LWrwqMCPyiS3+JxbcSoUgRYfNnKuxK/sCEujtU5byJbqzCus
CTs5QH00Kwhkl9/x65iucu4eccqGgM2TXaSx5QUj01TirEtt8EAEFWtnDoqX
lst6KTy5OLpmDIW+q+0S8BEQpNLU8wGA5lt/+aA6kScsiyLvUn/3mtAnvt7/
xM0jgeBeVIhkFTmoGZgI/4N2lZUXlxM9Q7st1DggL9uaw3KxzkkGNTQ5Y6SY
w0wtkrK/95Cy/iDpvu1CSOafRkx1yZBPjRQuZ5CIhVp4tL3AOOW4Vv9A0oRT
mZxiBNF4tPt6vzgJIMmP2WL6xAHpPTj0g6kaqaUjQ4Q8n23sZBcINEh8DHta
pTPc7frN1/39s+WBEUY5MhbmYNQJEwh0mxH3an1DH7aTjIssEx9JdyoNecu0
aDQdUKr9V6nND5uV6jfr0HF+2vHQ3zfRWFE5jSuua8xithnuFGLqfRYuG2H3
z/P9+Xnvdg844fz9sRC/gsGcojOrKqHensvB24Nd3+Hk1+TNNcMyS2wSceE7
Iz5j82t3VpN+4YpEnUhCKbebku/XDsv+ogsjF6AisReWcvNxGfEkeCyR193q
fTM7nBuUzRbdmsCoMC2HNbr9+0blD/r8wByA0OXNfo+JKOn7JpCYA3gxWkhb
iumUMgWz0/tRd4GNLOF64eeZyFckmO53gDFaJFYSXwaF+eoXRTvnD5Q0pu4Y
tDOXIZ80ipQdQyu6/8kBmvreH1L8J1d3yjUq8w2uODZcvSgpCtBHk2a0KCyO
vpKfUkY2qlnHWDqo+GtEIJIjE3p0/oR3lc0v3Ng69dD7/zXFRMNRmdWS2QxX
niWTSqyrr26qzrtGX5gdVehJbWFZOQFTfW4AgmJ4d5yoXO8ueK0nSY0pmE6a
l9hdklI/HGnigGBqy6DHpaBYevoeknr66ly+3Wbg2kVkvUDN1VRe53Mv/hXz
IMt6JydRkP/kZarcWR3lmK6tQrE1i7cvkzb1X3inA04eFB55DYeUxYMIEytc
Cw6CTwKPGSGIakCh1rx1XRPBRxkDAdMgum7V7qmNkbUCzqOsgQu9ps8Y0S0d
FnlMbjGcWcnfEGn5JceG3cdH98UDvITY6uaGgsxeQOoshBdAecYR95WRn/i/
dS9Iz9lzSIEkyZ0Ey4akn92nPFsCMXRYBOc4092DuXfkXNh+UDz8BbddTiov
gEecMq2luEFgk6dicLAuvSUyRIQA6ICa6ddAQq5yjM99ru1Uyweeu6Iz5fM3
x3jfCLMdXoeVtwc6tW2ngj3SSFN4SS+wOAek0eT9ZWu2YfA0fWqPhwu+4Cnq
BJKpsAB7Yeh0VLrcfYJEQVUjhiUwlyy8HfYK6JS16p/v+yW9kMvwNpZ4RcQC
dcr2s1tAd70cBD+KAFU45sndRb5wlHt2gc23xI9AG/8ZGXmxJClCIl/lxPqK
edDVVwo/YojlqlggKGrdS2a1yEB0bYROEJg9EWM0yHhkkfCSP9n1dsNdB7sU
1W4S/t7zv1eaNAJKBvIQwsKHH2Bv7A0hnJfbbJSl35m3oKATgQFvV5/TtglL
yHanWt0LjLX3wE5I8LmxP3s7qI5mmuvRsORokUtxh7viflZLjhiwZ1qd0yEf
oy6VG2ZDCYKb4TtNVePICTe7i854TmrvyRz9D2jVK+0CrvQiN7sSJjfRRnJt
d07jRY1FHWC5feGMUPgl77oV7H5bad6r+PR1a8nTgudf0UnrRuOZBmRNWONw
SXtrmliIdGuMtGbISJqBW+GSbsdbK+gw97Cid/VYexWwDO1LsEAFtaveqF0S
iRbj0+RkbrDf5Nx0h5SEOdPTHV/W5cb6oYIszcPHMMW2k3Xc4LBMleXkGAIS
y671xW/v/wFhVjGt5dbu5l5XHBgttqSazOzjcO9ukxljoI8hYJ+PIFJdYcZN
WIev4sNnECdVYYRx/QeNdQ/eLN1tldQuspHWPlLTQ8LOISHwZf9maCXokLS5
ijxNMNNO2bxIRk9zdFLN25UzqMuSUtzB9DjLqGCOFqHMtqC1/30CtMFhXxvb
gUk3wueQrutaKKN75w681F7BKUoQr6m8ncVQtYCE+ERJpOhiMTzjFVS5f6Ve
sO/ynb/8rEjX5CpLJ4C7ortr43E0uad16JQmnbGPyPHy6CYKPzoy/Llq6oO2
41RZgRjaBnfuz3lyg/PvxI1E+htsef6hKGvv4ViCCqIWAT+gYTpRgxHkO4eP
tm3wEwKFQOVUrp32e2eMmLGkEXjTK5ZId1N7J1lLLS2cLn9/nmHavbEJj6Ds
gYegXrisnnA3T87NrFqRp2XpoiuM05ovL1YVCV177zuG2f4AzdJX2oZR/6lh
1YOD6pOMkr9tUjamDuzuulWj11gdLa+ulODggb3RGqLiGqg6djfYr7HQjOZi
C2LvjJLk63mbtB7Abc4s7YYBZMLKjYTrWIYIk9lcknbLY2B5sPaWqlF0OVV5
VF6NzLdg9SLRon3q1jpmoZURopECI94hnCPS0l2a+tGb+Zt3JfzqO76eOfYl
bWpkKNvjfSau9mxuGKH/l2c1nBfOKg6ry4Rbm+VcDQb8Be4qHxfDZ0FFxmLV
MTrsXIUTn7Md+I97ckjXS31g2ynU3vBth2njc5e8pUbe9qM0VViwE+BN1GZw
R/9nqvFLBt1E6vqWSsMRhsQUiFWRvhJw4plOKKEDWktNmnVMa4+07wdpNdVZ
bjQ3n/c+FzcCKd37wyxFlCxHxMDETGbjNk4VDtVAyYZSKeZ4Nt5CEXUy9PAs
kwTXcNt2dUcJK65dDpM6rp7OOu5rkFEzXm44C01FXTx2HXUp6cCIp1CDEkGA
nIK3wjt0zezsYeckMJsH0GtIrJhPtG1RzAufHDzqL1p2y4LnElb4XzkvgrVY
Iodts4J4vMQylSVcKt+RzlvmG2x3YVecVjOI/3CIs1uh60QVkwqLMJT4PsjN
sGmn15JOGlyquz/0LPbfsSMhJaxJu2m14H2CRniZjK6hJ8nz+pDyV3TkcPgM
RjX+mqXpSqZfIdhuuLwZWI0NW0/F45i+XlYXZJ3u/KKdgBfn88U25RnuDc4r
d7tAGvnjJidMAUYFTXepGzADkgKnhkom4I4tChgWUh1eUV68ZQn+vyh1t/5L
uVGtMXj5+JTNqCJfLObWPUNmT6dJGwoQ+UkwB5oKdP56I5H+JmDTQcqhb06x
sJxzx3rEBs/j6mzk9Hyr2mb42SP4JLH0pnzbOyLkGyMaOYxb4TKJMUrfsXmc
kS9u2mqe+d1pL5jP44+3AMoFdkELuFbHgxDfeJHxoEmoHmhTKALWk6HJSySC
mHG9RwJyavjoKHvBNsEIrMZaeaZTDMqJSomakvoKDd/a1Wne2CMtJJxW7uDj
SEXtzYM6kKMM5xDi2D+663KrT0LXiL2zFoS/Xrjt4vNEKj7Gg3DIJG/jV/Jm
tZtTBuBEwvBtzmBbdEWeOut3sw8MC1IjSta/NQAa4Bc4ZrKUK3YwDaaAt/RM
+OQMTYx7+wVNHKn3Xt1P0/HW+LZdkp19FeN5oGRsZ8TLHB4yaThVsV8HxFhp
yH+Sf4cl48Z1xksOZ+XsooEPPKuar02llVe4y10BbeSSMG8uNtSwBmASnEHK
7svdsDfeZ6Exa1liWwVeNVK6wZ1kuXKGNmc9WHIeqywPTqaHChzqZ8hJh8xU
zvxy8r3+CVe2bqqJPT4zpp7bJySJiqk6KpVTn4yf80Bm7povxQuVgVeGyTD+
Ti/P67ukuo2zRtKsLuhS8AmtKD0NuSTSuvEnkA9pYpvWK0lCxpbzukZG8aLm
EPGAhbQhnSDZYfrR6SpCgKG0ucIV5t9IU033O4VEI0xpUBw7VGRZRoMD+Gql
GFPYVCfnt4w2rWzs3Uj3QyWcyoE3mrSlRvDN4R7bm+rL7SExfgw3Nu1P+Z91
xBz9KAhOnZsv9SxF9ove/PGmVReTUib7p7yi6tl5jwIfE76Vu80wNc5U6OPT
nDfM3POCBOgGZGy+g7GD68fxiBMGIn+Y/0rnHnKFMSZtyM1f5aY8/ZqPQlMO
ilC8FqONNp0mgAdqPrgAq46CVO+ov/iyEBCLZKQ9IgGn3FMHUhxKBa2ZhdRG
gCOyPpcgdtogAjCOh1DIZqaUCIqiT5V4Ms7HgqZknQ5NyYNckIqjVgJUsnFW
S6HvVRMTWuhVO2jpen5L8gtlF0bMm9ZohLTTDm/tRdXknOpgfWk4F1bF5KCw
E8RvADDS63ZuyGKmIdoy8yedxn0gLBTLoYoy2vxqp+AqV7ACLhBrsxYsW0qT
pjDWG++5TpoA67poURQQXkLzAycnkG86h8iwiFXVNyFc+ms2kYkFFzFQNWXf
y1TTMUdpWAbEHPiL1e/qDFfJLZtctEInUU7cO0uGNhaP7eDJ7A9wzfApcU0h
wl5FOf/wU783TaOUzpiitrP4zjlAwqVyZpE19bSxYpVA6+SGEQRakot+wIQs
lkt4wM1lCcTDL8HsyXg9nzZnOy5oWvIoeugOgnAEPgZ3AX1M+UmwK905cVCj
dMWYqfdR5K/OpZB0/oE7eAQy4FvJSJ0rSyxI+4NI8q1YV2bxTADmj17uk1ws
Wo76tfHa9WUghC0PhPkHyNJyN41uzRP/4RHLqkmzFUNA6U31sK02fe7BOtpU
Ceb0Aq90JF3hPDh5F8+KG6M7RkS5HpTdyxugHWsgxt8wwXy1hQ88/EMTGnpR
tIVNn3qzjTaJZyVT3Tzy6XuFcX+kIDU+ru8Ixf9NsDxOzwPVFliOCuvO5bl9
wYbKXzsWMwL9oBkMRvmD+ISALWkNDSts/wewqClixMH6TIeAqfagavDLnoWo
q4P1Fdteb1tfaUEn3nvXEEbgJTL50Ky984Km9NSUma3CWsrgn4BcKCecRGuV
BvtCtLngZHUFMwiQ06qXGtl0nR8DsxdTcHLjoVaRePG7nRT5Hq+382bjnba+
U+0qNz9NUxlsarHzXyQ0IKm/DApbH3k7AqfRg2uveA7QyWVdEzxlFaS9vN2o
eTXY5IYQZoLdNSkqsYfYGFI3V3GPn81w1XMmiVLXpUb3GUgdycBbsF2D2ylD
PioYefRt6kyPbDp7yqw6/95OFrgwj6/AhzNmT6PZITLTxMUTpJidNg0kAGZ6
GS5O4IoM+wK8MQBf01kP6WEvY1vlWvvKdQnXzAcUOfBGz1qJ+OtZVScLUKqR
Voh587V8bmk0jnlR0LaJreyorR5p3tmJQ/r139+JFPROHn63cyv2MxPbUpY3
TlC+R8Hdl9mxAACxZT0mE5bcf5URop8qqqzqzqNQetN/IWJa7audpIvcz6Bd
kqrRfUUTARnLdav9KJMZZIGZsHeCV7ZtW18enYvzcaROUYRg79+9g8kxtfkz
B1xXo8rVWlxjDnPY46EB5NAdE6/iDop6+nQW+KOtZcRzu67Dy+eEHdVXar/Y
HdSoEZ8iXNFN/vpdyvKPPSyRFUJoZXqmRzgRZpvCs5jE7YdqJs9mrTB9pjGE
KWuLgIbVPmSB7Xa9IjhCz1in6Oz44Q1uelS2Qv8hWqym7kRnU9xutHIIXL3z
4S0FOT8tExtFMa2pjlWXptHjIZhGgC0uv3zVhwkwv4bCZhtZ4pHMRiyCrztf
8Mog4z0jSRRChdP1QCI53BKZEtsGaQpcNvQa4JaCzdOeaksKwIZl2EYCjfRW
4vVjg/aD9LlyB/famlO02hjMWkj1EFa9X7iIRUWZGf3VlTSu2SSMxZoS6eGn
e3opnCRxJtGZIx02RtCrHkhQR9XebYHSXMOBBKj7XzNfvSx2bb6UZANXMd8b
Qw+HZ4MVe1ykxVDD8dooFtiwqBGYkBn2pDECUoweQjGx31JgQIlJknSTYBES
4+id+P0AyOEiNL2FkBIPQqrcyI+2gWYHQeN/49JhUMR14LrFlppl2liWUNSd
oMvsxRXctVmRUzDToVrovCFu2oGD/s2m/ghPON6G+CY/n/HBEaGw1sqXwTeE
gIfJuqWNvbP3phUgRzYs1XmuS2sMoQxC6mjgGLzzH4hGoPmJHevsR80UlPBG
UoSnLvkg+CFF6Ogldro558OGYQqgmoDvzoHqN1NCxmGdWj61OtrWBktVfysy
M/hxT26NKHEScV9Y8TfFR5yGkjJUzeGpN7P0Fq0czRbyGu2l825bIK0vZIH6
3sd5Xuee3aotamv5Tumd3XWoZ7pJn7HHsUWu43YaG0p70rj0rNPwnlHqSUAi
3S/iLSTh+Gr5ra8ll7sS7WfWH6BzNa64udGlF8NG9Ox3XRuFRG7nlQPtNbme
D2jDJ0swa3s2kOfAKQHibebidCwJh2VdYxfWQCf0x5oEdDlkX1jT/rCpjtKa
l1ZzTksmkPPnQ3XNJWDbMZkUVDYUMWtYWuXiU/QBwoR+dP4UtY3upKgXS0kM
R3sp8+rRbqKft3O01MZHfCab7pCIHYikTU7atJkci1tWpkMjSAIF+hLUxv9T
bG+hcg4Iq2rSc+PJUzI3VoAGfMGFBthPUwORV6L6BfuDApqmILcJhEPwlXM1
dxrNih54pRiJ4cfqRgpbRfC5c4KQLEHyCYyge5mofWhbGZaWpMHQ5j1zU63P
yM1e6iIk5qcQYwMmWrQ8u+jpuBt+BI/aki6qU77PVswyh7zOZ9hN6y5z7cCT
q2y9OP8xW4Mekp+KVGqT/3mi7rpFSbQVSeJCy7w+PiXAG7nqHHW4QqIGZJTu
VR4shKRLu1kBy1CKq4e5ZAsnzEmnomdRjHmrNYaD4VKF1MRG3vjuQl8JIWI/
j+CY7InXxE8ZEApLZbcMYNCCBoy3774kpMtSOxffiZZFJDFoZiW0yI+tjB9Z
7Oo8HoV9TwfhHiwIlO9yBrh7htyuyABxU2KwSerznJk3bbl86AjVEY9dxJL1
Jle78pfUcxcetahnyzY3+w8iBrZh7Q5w7bhnX7PCPS4PkTKuKxrv3VgLF4Tj
9LohSPeD+aYJwLTaLyMRpqmm65vaN+uSnK7sf1xmDiOVITO7FpvOoyeJg04J
T6zJgYwr7XWhT37b8qkT46ohnO/EhoUXk1KrJ15jSmJWWuVDYgnj4Q3+oKQt
WtMj8K1KFuSrzc5yDFJwjageqVc9XadB3uZDSUdh8CF/hLBZqnJgbS+Bbri6
ymnpzNNLKsvqNcrcAqhH4Y8+GCexTq2RqPsBl2y5tTGEunXhGuQKQlw6+oQj
UWKTVEdJnMgT9p5sSTiWljtAPXPqaNQcdd5vbvKvdRq4/HYtRaWZffN6aF7q
6ketfBVUiUHXYGsNtICPlKwmLlGC8SQ05eVw19Yqtbb8cFSKHV4Oq4tGApoP
5O1CcJbTnxWdSxmob//+2zWkkFM9YVIdTtAzH/P1MjJYQLqjYnUmWi0uiKw1
UlpJPAYCFOSGhx2GaQ11jhO3TVbIZFgdGMeMgLQqiWg3b66nkbnFz9Ls+iuv
Dmf++dbGKng/+LObrn8q7QxSkA9GDwcMaGUESGpGgnXo7SK7R9RWSLt5eIEI
mKUBFCZFPYvH4aH/OFPgjNeBv4Juzjrli6B7uBrQY0ZWEAN2bCbPQY1Oee99
gCFGrPXG/YjhLZzkDrsL7bUAhVQhaEyydygi3LUzC/rqENHEblciwOVVZvqE
dw2WrtHe9TM1gl3wi7jjzdCzuqIM7OVCW7oY8v3i8YfHcgjejGafcfu+A9MK
tuqkt5aYqCTx2cqCI/MS7z49xv4fqfjtoAiU+NlyBDWX4V/LfLWyo/Q+DMp7
0gr9tx0O1m4Bw2jRGhKueV+Pu5VM/OnpmjfVtsvQiGqMXN73TT2Ie+7vI4+n
fXgHuBKklq0dHnbXSG9Dy5USVTBJ0k+lLr8IgCjsjFH/sk0KGAbC1IIYi9VJ
YBCqWvlE292ItNrNHU2XycnRUmEMwHZPrPiY9jW7S3Pi4PI8SGy5VVcBSlPg
hNZ8xZMwxut8Gpx/bA/jx4nYdWvRrK11fyHcWYei88EgVl3C6Cn5KAR7eVCa
JqW8O9fCsQOqhZZPF5Slji+2Lbu84oPUTSKEgzO+iIDCvhVwsUYWumtXwhqA
T0lL//q7aEHk6XiKWL3EagVvoJv7KzitrPnjf30X8P9KlFct0HTjvo0NTtG8
si5xIsEmiCxDYJxlkfUH9XtJTZJse1GXVmZb/r44FxW+bh8ku9CQVt7jZ3Kc
YuWTM+tjx9DAiS7haKKySdhL0ue2FdCw8nMxvWZut4kDo8dk+UYFLDST7cim
Cow98CALfxd6s3/osxU2UEHiix+hzXDnouSMkIcgvzjgss5/ddI2dH+tlXhH
+LrhX5GbjHNpgpgSvIGgxalc7IJ1gcLpXUosatVUwMnlC4G4Oz2otjWZAkb2
lO83FJ5FDh/hgnaajLWQ7EkmpCIkH5nrxhnguYq0lyUzyCp+w7rccd8fddBA
W1gnbtyHr//gs/x29totQmj8JMprqmTDFzt1onEkfbWLPZgnRKYog6z5XQz7
FzEwKfrs3ZTRwc4AXwn18IXrJKq2ad6Of8oNWUMUROpDW7ZJNUFr/17X7Cja
pvLK+YzD0x8F+c+h8PP5hty239CbwxN7n9Y9r3OotEhpvDdYXHY88Uf6xFeG
OhbbeprwuT0l8i5y57QuWclp0cwqMZbkrRoyxglmHLTn2R6MCuOGcH9GiYPr
ZAr3stLcASMkqE3Y4HybV6rhu5apI35AXGQQq4HsaCduUDPAbEFF6Mmb9UlY
ccucDJ5y8g23PEvQ3mSwJU93x2ezZ3C81DvXr/RRMMv2uT8EhaQul7GVRnbF
lurrUpIO9h1cRoGB/Yzvmf9c+z5gdJ5xpTjVY/clkQmR+P1X3qF+kveE7sXF
vGBfGGpl2e7OM4o4S+9w6uIJArisjs1XAbmnBc6s7Ob/a9WFn9rboxzFCHK2
WREoatTaYlmts9MbMxDewYeBuc9L99PnUIdZFxkNZX+7ZAEds/7zL6ZIRVvi
r3T2DAjVFJBcB0PHG5SBRuqBLRspYasJx+fFJhCfu8N9p1/Z5vnXLK1hU2zz
Vwkjj2lCjFF1Ofsg4qqib/rZG1WEs+yHdMO6y+osSNULch12K1O91iJ0mrVq
AUO9NW1bQteE/P0JbYCMTHPQtA5fWx++4PP/9/GY5yV6kOjWDXEp1NsGDe3r
mAtjgMDhWaCYpvwnnBfNPD8xUESBAnGnmGpCRfQ1M6tm0n0WaHk+84ljlX8S
lMAv0eb9b5CvlRWQwku3QeCtvMq6pHR2djBVtkgjqFXYSSM5/eu2dOL8AuhA
mm9XZc39YPp+0bsuveO3fZPggol+qOARC80g6erJ/Y8I0ELxXwChReSsnIdd
AbfD6iYZEr8R4UTKmXN7pzEdJzKG4ACXx1fqGWTRGYGAM7PfelRSu+T8BycW
IwEXjLLTQTq5Q/7fhGYAoTg2CrtlCpbiMEwbrhWBsgEo0YgjmmrRqFo/UdVP
cb7qCOCeiHFFcRDUIeVoRmIWkOgrm4lN51v8UbSybO6P1Uf/E3GHd/c/D5qD
1OoBs/yQEMek6dTY5sG/4zclEpre8rwNT/8ueSD2ZXh9nB3SvcpaWZbxuuPE
DD3nJZx3j7iYItB8o0V1bHyHe36SqE4wa5U62/3AtePi2DwUD1bjQvL8HAWk
j6K/IfFKrpUv4gyxdErDt9rtxfQDPJkDI2VIAzfbNn6jFFKry2gL4Mcs7YPZ
ibyC9whPOjnETlR3TQr42C+iTHeQcwWrQMQiN7ymDnYKHVq4Qh95SRLIA+hU
/aiMgJRBnPfq5ExbenJhwSEed32M7kUm72tAUDZCTz/EsIaEMsh7xBqpcovZ
WH88cDyCqP+9Fk+BZPkOyw9nqJdU8Vcq70cn3UgbDcWSt5RDlpSY6xD2a21Y
CJIlk0MlBeITyaJOyJMosR+CzkrJ+bhelU8rKhyUMukkWTvQOSrAh7XVcILu
NN37Y1o3H19AgbI/nnTBscjARK2FWb7trdT/8xBiu97Z0gjR9AP5hYwqHwfT
i3ZwhUXkj3NcMsMnJ7LlkohHXVR89HfOydkELoBGiKeE2cJ6WmnF8+AzBvYv
2VECPZp8b5WpzosWcVQP3fx2LYW58K/lu1OcZnqmyu4wfaqXWQKXSVph7RpL
LnMO69jLz93w3EVuQQavAGZ1PCbcXVxb2aN24hPPTEvZs/Y5e118LSw4veTI
rFzhVEAQ2D9wwVZZpqABG+PoNHCxGex/GMx1Uxe/JnCV4XMqapS9iGvcyItU
KIqADQdZaYfGRYrPT9q0bCgfMfCZqkTNAsGPsrY35UjykT3cA/jJ8Suv0a5i
5v4Uw4DECPuYhpIOJi/jjiDBJRxIjgGHddRIxOaqQajqfn3pEZE+Z/Q5cMn6
384zvNWWifHTmYKTMbAIdL3EhrBgVMcszp07SEcWvypaZBtx+o0X4P3J5VHc
h9eDmZB7GiUCPJta5jS9UOucTyJsDpJgBMF4o012JexafQDarivvl+1Xl2Fd
mQstYkS1mOoU7QfeQHVaQBD6De/ZLi3Uy0OuHUXKYhLJu3nNF/UjAI4q3L9n
osCwCcjvqSHo6SQlf8J3s8J7abBMYpGgXbAwskeBveg4kvQIbLalbo7hbksX
NqdkY5uvmtFlzcoGnMgba0CN5hwibGQR6KXN+3OIrsWxhrsHELXMoUVOWMVm
J3hCRzYjyhUCNUsPgASzpFn/Ttg+Pk2GsS4fBYqrjd3iyB48odNIFdzylZbq
T2je7tRvkY5qdTqyJiaiaGslFBdL8+QYe+ac+s1iV98UCvyzSwG/gciEe0tT
9BjJ91SS54pRvkBd2lZ6SOjVeMufNMlZqMcHHur9hTO0iHCXnpYLyOkh7EWV
XkaGEr9JqV8rlMC+N4LQEjBqCAnVyP4Y7615pjWP6lIrxC8Pt6LlgLAQISiJ
R5GRiGuJGRvo3EKvDs8DmjT0xNlFuFSGLeuU/BQ/jHx+D0E6fsVYxt4xh6FY
zPVDOu+3uaiXx3F12evozA1poJ1uYB7czyCKokldnfYQOheU2BLM6T0+wRzn
0HrSkTJU9XuREplrrpM0q0Rb8ZT4iO5XaMUnA57fzFHnsHZSJDCMQeZa6N0W
itPgaJfXuO+SI+odUhtpdkIB1zMvED5ZA3Tw8CGOIRGzbceQDyh1ie0z3DUb
jUKEueKzD/glNE5MugpQ4dtyFGi0QpMU9xXDHOMPN0chrFulyOczieX2mi63
5qaQpAbvm1QcpvXIReqoXFpICCrsobLFs6A+i6+i1rQ4QrFuodxYeHgBqzNF
D+Ij404Rn9haD09judiJp3/yLp0Op8LDHBu0fm7U2v0shKLyE8QyZjDHpUxF
3w1pFOjCL7EBh4D4gbXzXu5hx5KU0teutCTPrEvoPSTx8qcOSCBMOKvw5HYW
cquZXO/IV34cyEJNRHBvqdiTU00SvrHGKo2Aik710anD91BzIiYjX+p3oKB5
s4xebX8g1OynYB3aklEdi+9jgwmuTAU89RRtFqJ5y9VMoisYJc1IlklsFcrt
zyNKnWnMbsEc8LHZxCPIPoQd8kJBQV999qJXd6geHBAcXwxRPATnoKcEQkLR
uuQ4iqAqR2WaiDgFbt1RwEuwJbq8J1Z7xPPTEfgg6NWG6SxxAQJhJrkdwfF+
ksFKd38/TDqFj/7cmJyqM7VmZZTzEYvDCTgzA7GAmcrsWhoFt8ykRyoX1PU9
DK1F0/y6TUFXTaOhlQgRCzKqJ59rh6X5BPTBE8YyePbKu5N+5gJnscSndhBP
MEE1TQjk+59fV3YnMrkiW/OgiR3VAK8nS6w3r9nuwoNGUrGUL0DT/u3umeQb
XHS4Q/E/wVbbURxCZL8xMXxTRE7fRW6P4/GH+/xM9flqwnY1vrc6kES+WCHg
mwX+34U/swFBxvybVY1+Aqe6HNLQoARRUdUHZL73uDtTuKOMoIN4a94UXhAk
XChzEbetBbrwKrT/Y2+DA3cPzFDeFlaJuDcp1y+BQA40khZ7TjUjQdmauq4S
sERS22X01n2vIjkH8tVV9Q5M4CGh0wykfx116WWfyBlTj7eh1kdjr+yxYY6W
AAV9sfs9ma7NBM3RRTiQy4kwd5PxF9ot6ziobz2nXx/dOsin6LHMxq0WdcY8
9I9NV87yle1h/TNAIv0ShU6yvAkMOK2KAccx432oCtSzNNYewPsJSeWBr0Dd
jzcJP0ZBukVL1Xo/RwmEMLmtGWRjxtYXDgbj7Gi5705ToIP0HyxPdoPnbS9z
hj/+sRWOVzu5gRAYbM/GXHJbueZ/iU5razXnp5bsqtuGc1EURcC/EM3sT2zJ
XVKFXb2ggGZtYASrl8noGEI2HROp7shY3aB434xu+IFn6deBJGTR2o/jDKRF
N7GP0Bx6M7S+PkYi90Vr+h0Rja1EogfPE6XeVwBgF5czHfVVZv3C6iIKLLe6
yO3ua8bqGJvAkpMDtWKNJmOMLbdkuXMNFSAyY+ALE5WJrzAOC18SZHOtqbYx
dEN6YzBbxR3i+dtgxhXITEKhOdqaJwi5+N6Dpf6tLzZo9M6/ERVWTrIWmAo1
FFYIkJrbFKZkzf5y7XoFL3p30WcIhV6ndfU4uQn8tE5mk6vjsCA27TcTEoJ1
cHB+MiMUgLeAFeMTPm34lz8WxvRI27HwA0K1uFeuhFpX57wV87UOpIEj9JqC
BOGEipIfhvaNq9hFLAs1CDK/DQIHJUyRVh6ghpe0xrsDxnQzq6rGE2FG8G/Z
25LL7KnqzEKsdrB0qrzeubnPtnyQ27VuCOoraLLWHOOwzLAIS31JOQNI+xdU
Z+AAVoD1jkBfPrO+graFHa+tm0MgMoVlp9Yov4KNzj/li290uCdcBHmKd2TE
mc/dTl+1pz3CeU1HW2j1lo2bDkpeICFlaG5/MFQoFqHmkced6UaKFn4X9LvS
sC/BYkyYUjXX9UGaxu6gfj2FddgfDbyNOzQI0dkmueJRhV26VllryWTfY4HJ
83EgCzXfj9m4nRbymlBKh0UwePfR08TYcLjUAMwMtZNPnKoNgokz7s5Y3qNt
jBVW5Xjl5qHBVFa2Vv8tVydWKCNxVOUozUi2jtT6mVUwiys4VwUqr3YHzkeo
7bbU2/hebz8MNh6ZnSLx03UtUQ5gJqf2BjZrL/2zQThyWPnHk6DOEvgUTZi0
3Zg2p2CsteSQWgT6UT0joJeaHhs/EGKNeDxhZnbsmiwDOF6M6/EMv1oCNenH
5DO54DufwBcAZmUs/zXh7L7nPargINYU+IBImJxOawbzM/Cdryno0bbEVJtK
mZsRnksiGNs5W1N9Y/6pzP+/I6mCzmkm6Wd7zcMiFvgHSQjo/PSiffDK1MRl
Y9lVMSWeLxDMX9UlZuYfDKuNtEy+ij8o3qrNIqLyWiVYhB8XkGTcOg7LN+gC
b48t8Gfrqv+izuzq0QbDrk/nVk39Wxqehznl/027QOuo/DEYTdK1gKwwZR4J
SPcBkrz4miPmVnBYsDOoxgG7Yf7pyLcmCvvV/UhnkSffI8JJm5tpPxUAkynn
mIUv47sZsWTDySBcpe54NoT2WJf+fa4lRvVLIj1aVG1ngg/RnLl+c1MibUtj
j81ksJwB0uO16EIBNqMIHnzhliCmP4cfNCiBmEVg4CuwUsnGEM/UR+BfQFFk
zfvgGbAK6cjnhTjaI08KHV5hbWlQh11Mw6JMkUjxOtogCV+Kz2rIlUCubYn6
ozBYY2E+9P4ZP7ynyN67+4zoLnG8U+whg71l/jm1YQF3CsPQGdXLkV2sXBKa
IxDUsQZJzXr6r1ku28Awz1owYB0oBD4iZfT+Sj7QMBSAPe7g6JawnrqKy5N2
bb6oMBnEYrEWWZPDqa4qxogavoIQPGz56as+XJnCwKAZla8bA6ZYQ+/wb1N1
3UBXv8M86o1//zhNEOCuEWP0oqylrxwkwKp7q9Bslhtn4EqFGj5F4NFB2wcY
+iuxzOL+AC6PEOaOLOSuRd/la2wpxA8LSD+Yb91aC5esLuuD6OZRo6cWAA5M
ZYQT3/2YCdtq6voNNy+t7g6HAPosKPDGn/ovovNyQ/nUFNr2DYQ6SF60AMFE
G3IZzAYBy8oHAe497Zs//tmn2++CBKwmJg7eTJ1kFKkZpviggfa1+Y77RNFy
e/c93LrKk2si1Ui4kNHEpPpCvauzZdIpm9rXfQQ4C9Bt4NeaZ37Ht8uhdojh
ccXvqPtw7Dur8AI6NfCye1AXFPMaHbXCgubxWW9SD3sqrNGSXLO0AbmY5+y0
JuuAf77qTAM39PEp7c9WIS/AQFjCwnnExEJi2zjp6VxRrrHLi8vx0g4OaZrU
0AKc41J6686tU7G/FQZSoNWc7RhL7ldDftvmB4suKsjYI6BWuBBk0334rpFh
lGAGwYvVj/z/6lvYyhcCx2F/HSq4cYXyYUmgJ0PYZbpvJNcdHpvwSJtA+cJo
LnQnBEBtCpaYRp+FQFcENi3zaakUpryFGZnnSbq6GxsdhfX01Yl3mSoq2MKL
6U72Vg5L0ihVkdHP22SA+L64PLUh72X6onIp7665MgFEfEsLB0lKUgY1nETx
Cyrtbsc3KeoGd4KsXjoCURXqzUnHXswGt0Ge3UaPQSuuTJAwIgOxyhPgMAgP
b9aPFH9WCwuOzwayNklwT9sRlA8cJco/VOrfpbPah3lAvGFx4Guv64+K/kLH
UJ3fObHwb39G/ulMtYrQpVsRPPpOY9pmTOk2vMm/FQCy7L514uBboEs4x5CX
Y+267Jr2uLg2b4V7f1loWlwLWtg9T2sgSvflbDeSjmQFo3v+h8uIykdx0s1y
AZBxIzT+qGMsLP3JLtHEva4e1MsRQ58GkJc2UcAV7zYVz0aBPc6xFn4c/ykG
YVOQp8RmUGKbmz6LhgeBduLPcX2gfaxRHFB0VmS8LiDa9thH4+qce1pv9ehZ
ERUwNRbXxoy5EbKlKigunU4E0huAuiBByOV913X/HXyjP6yIepfTt3YBnu6o
9rAqR/MuDcbZp22q/0NpqCwEdruVzQnhV8pumN+5rAEEFbu7U6aHuM5vAd8R
iaDM+96YMAwekVjnHnKNuegfixwP5N9DKqw063efBDXpDN3n/YEYuzxFli2v
mTeOo+V54WoWE5OuInm6t/ZWP8wanQRrjMlQxk/C8uMl/miBfz/W+fQN2EWk
JK5XGUFFZCf4jIhcweo72uAH8OGjsZ/nHhvjoiGvn/ZURes3ijBKfQ1I3eyt
NobrM6y+OOnFJ1gNUJYG6/8sr1I8KBNg11I3gEF5zhRt/Or9uz90z2qZSLTT
VT4okAKE9tyqNymfHSrcg0JzZm1oPW8sSZaTo7zk39lu8xYINymrvDk6rt0c
Q9Jg4QjXyF/g1tk1UkAjwOisd/bER2eKN48p1EtRSTsHW7I3zJJFHvew6UtU
i2vzc/nHfQoAFYH4bpE7ispxs3Vipc5/cOXGlaYfZWMjHm9x6IjBfTrP5qDN
4+0oxAGVrsuIVRrXIx+DnTEEDrHkD7krVxIyYSnYM0p5JXgriig3jI+SPJjX
TE7ku/DC2wycH72Ey4JcQTAsu28CE7vkMDebyFYgRia+1OJl6GMO6xJoMpdH
eZ0+juhsQdyFR+mMGXh7LYle0iPRmtXJ5H2c81ny01SG9JrUHj5TY5R3jZ2m
Pnlc47vzI4ZUVarASg/YUsfKelKvKm2LdHJbnfBBye+C22/8Nkmbn8Fg+YXO
I8F8VSgjNXJLEN/f0H8Yw/ITNOrDQNoPxZZx7NhJG8B5jKq6PwGr9mY3wT7D
J0MS1gmHMOsYUpVjon47IrKTBEVFowHpZWVqIsj0BBV5BeBZaJl/dYaENJZU
D7pcEwixeuImchMIqq7WNE9Htyw4aDMjEmjAXaeFCbLPGfOfQ8CFg+2k1Xb/
o3gqzNSc9R/8emzXF5EVijbFsuoZciSt4thUAWGy15PEVo/KPyn3cl74GKmS
BsHo0S6ucDcfIRzniVDBhfSYkX/KYIKkqXjZCJUjqFA8Pu6j9UKFxEK03CYL
5IPYESi2WrQCY8OlCzAXn56vzEdNzRqgOCv93hrXDIogGpj/8bsYeC3AS4S/
M8xtUnmEFQHXZy7SqLXTOxs3JdlrBkd1xBiZTjQtvCwizPLAdxh8eJ3XndrO
aAUjLuoNKmMOacyiFmeU8/LppqJYIWdrVoMtT3NyzAVwHTh6sZF7tls3YJFK
L5kxAr/92EZB6J85mNaAjixqgLqVYsmuQ7sIFpW4bRihfivg2fSyM3oEeJCv
v6qj/fkfRZ1hdSdeQdfgbrWFnXB1Ur+S92KK7GsSrIo+GH3HFc4LWdd4IHsn
MnVTgst5mR/9kQ6eIa1SFWSQl2dRvrzhGHWZZKsG5gY4TFN7Mrp2JrbeeGNK
XFLcUtwUY3PHwRSc8a8v71EMMbPDuRPqMQriBzsmSu2IrE/1CWP72PZ+Z8dd
+v6/sYGJ7ll+qIir82reP/PPHorLXCmDsL1Boc8Qw9JA66vHHJRL/SQfpu/5
dAgooZs9ZV4Jxa6bkGt1SKnFwodtAmFSNwC7iibH55ahIA3Y6Kk1n0ZLFGGx
/fMEOKkbMkUnpS/Go4QxmLSSAHdtnczimYbAivSIPo1y/vf+xd/v7GwxmFoq
EMCfJw5z0db0WTTDbURHt21vMiYrfNB/aJ0+si7VF7vZL4f658gVU619z+At
mbOHU/LF/ZZWeZGrnXvG9tRk1kBmaKTQ19hkGRdVxxcyUsx/wUO0AxZXoVzi
eqYd4t2qcPcjVk7HzCZDL3PABo1x9BDqMZOqkegULg+f8FnQsBXVNJQZ54ko
VDIeKLc3THLXRe8dGKboJgJAjoiv4Q97KQJsYsG/zPCkMWTN4oxuiOuQZq6A
oGG2qJHJp821Y8hIa0reqm0PV6e+5Ty4MRQnOEo/PjQvF1GOmG6pHJlDDNJ1
75lQgEsSsMm8RH/n+zaXejtrPXYF+HTqwvOzbkzY5+Vvg1Y38w/jS+Q1N9xL
CjfU1cL/+kPNLxJ5fWCNDTYh5r1CbEB+TzURR1JhpkpB8XNKfNF4u/78cDe3
fxgNOMnzv9ncdSw67camoM+qazy3Dxa6m0WNzHHbpRUr3CwK7jmr54+jWGL3
JJoVR0Dznxs9CZUXw1h3QWk+mNBAORW3dbnP5vwdi0kEkFKZyQWvei4FX1RY
Fnw3QNkPk6PQwCGltE/mK1k35uX8UF7WbczpYgGGxmTu9WWtsgF+nNPihXYK
0WnXNdN+99J7eAkGdqr9W5svxcfwFDbRK8nolOUiirigsiLDohIvnGZzttra
tfarO9ETMBVzzNGka3/wBDPVVT0b0cJoQ7soe08TMFnbdfRVgoGyAopIeo+M
2Wvr3GTpJrXEWNe9Hjyg0SOJM/qcKL8KyuKMBFAD3MiZWS9EDRT0LSL0fn+G
yjx+z6c6bNXlPDBhnGFHkug0ncZTakWakQ/GTYK4cE0dCeNixLa5OaiqLPSl
g10wXoY0sXWRO9qc/QsdH8i/WrTsbJYToZxqgSSUG2Yk5bEtj+IKKts6+ojL
Qm4QU9LKuI+PxsnJhuXTXxR1iYDQB4ehpV+kyOHPW4GcazooSm9MFUrGt9MV
Q3IWr6mw1Ld0SdoEwGXQclsU71+YK/6JSR9H1xheerdxRRZLC7DGwOTIZwPr
MiY7HPCCnj02PkZQ23mj+NL0q+h7aoZbzVWmuV+heLU6nUbKMspWpW4IdR61
lPNJiPPfsgEldWTJcmzCcCcC4TlLt5lwguguIGOWgK7z57xOZ97jO3g/CANR
pnA2y4uVR2c1ltmm0edlDgqp3XsYWGqvfFPBSi51ZosnFSITFascCSVmYNdU
VhPjuX5k8EQjJ0wMSkno/AAykSmImJ4c6ldlEbHKCELc/QSmTUi13K4F1eIz
uNQvvO0QB3w8neYiPGXuhJN3XyXJVL3XfOYF/5N6jW6rR68/U4ro0/1q9L/i
/st5VCUAS6WwZDn5lC9Y1wRimeFkj6Oobt/59FRMwkRoKTuXLcRhFho/3dAc
uAI8pZb3NcmagYebPBtXTrmNtFvSpO/uMI2/56t6E1bWBDRXHWvzTCa/4A8w
eoml2nqEKQssjhQyjorqqIC2PtdATG0wyfQVO6fTxgj75Up4hgdupYijoaKh
FpDDQ7G+iAJ/GlLkxZTAmGfky2sFwk3+IsaC1TVTfRtUHbII6EDCWjkjs66E
V7cm7x31Prwu/zn4366C5TAQTtN8PS5nmxORSFW622cHiNVNbJZnw65iSkkJ
+Z15G0idSw0mJa20JWHgYKQqbKpo2BRpMy0d0QAoyEHfGRndY6pPhqFodprG
Qs2FYh4cAwg0D42QCFSZLO3w6mq5Fyni9AeGRfvJ4Fx731cnfFv3/1J4OYbP
aBfCxPd9BfUqWZr0cgk4biHS5yZ3w2OFb1Seyaq9Jnd5GnAa2yBlcmYQxZYG
eMNQjoYGQN0NQd07Xu7Fg1zrEGFgualloK9s58FRbzTqpF+5LQvDBRsaXVAX
MbSkpl6Ek+vSlyGscPco70zVWCeGoPVscpBmSDpJ0wSsQi20L1UR98/gu6mW
7HZ/3k+x8P92i0j6VrkKJ7rsWLuLPMVf/0EQOPqZgNpohPvcB2SdmxcCoJ8u
ExDWCgKo+3nMJWlOhx4vYF4NVbN7OPmez9QmaME2WQppJMBNncjjJZ/QJ0AI
RDp2rGtM8ZP1AoBomdZqt5ZEBBm+ZI5yGa1fYKct5L0sTWpTSQpqy644cj8n
Q9Ru6TOLWIDSpUklONOox/lzlu2DpuqfCapMdtzuuU9P5R1XHG/SAdlMAMgK
FB4ZLVAwigQ0WsP85t2y4lzDb1XwTjdqzfaggeVnTvXNncLhLY1UxpHNoT62
242g7NkaFGgRvPA4I1K1AsIC5jnoN1SXTUvoP4Fo/lzgvDx8nmBzu44uOMrn
U32Eb9YDIj2QV4CzpUyBTAw8g0Jlv/sufX3hPaeu6G/L3v77/8aLi8bzQu7T
SRMahZ94ld2rLK1vnh6ak4f2pyDPcbHl8mIwNN40KMhAzo3KsUA5P1giznFP
yQaMkg8g/q6XKHWsnNLGZyeFbya29d4RdjYjivCAdQCpOBDU/g415XTFAWLU
mHMq7ddT6/WOMA4Q2PWCHzn3CSuwzTz9gamqExkZVG6E2rf2QWzzCUrqh7ox
PikE4wey4HIduzyfag4xoW+YMTUu33tLdC36zJMXOK7meHrcexGTkc00O22H
8crma20bx/8zl+w0Yu2W1TrTaZyczHjlVZEGo/VlZV1YrD3aacryJ1pzxzT8
u/mPX4me02thfNEn2PCJujGXOMTP9MHnZnUnQiSqMkAOQNun0QV0fvEb0Mrd
tm3EjuovYPloMuuVl8F7453wPZ6Zyc24s3uzVpj5T3er2IlxJE7YhD5NkRTW
SpKsFXi8T5UGnFHrRWrYq30yjDEmprVBZuAODPsyl12P1QgZtwKq7PCPyQft
k+IQgazN5weSsGFt1cAR+KN/FEjX0xrGJpx1ntP/jKWvXFOVuu/A1JB2z2B8
gMW2oNBCUcoxnSGWIbYZXoTMk6d3gTHJF60/LjPs7o2l/JoQZ65bhDScS2VV
CSZsTw1YslOvJVRf4B9rw1Osc0IgD1r69fGZfRCjA/JB4Imk41SYlYzsMkXk
ifTmNDp7tDSn3xaYRgTx7lw99iOyUat7YN9p1NxhP9PayyHitQKbk0E+NCzk
EO8f1poSS/aKRgYrfNWdi6TlSXz3xTXsV8Lnqw9/ZOGkck7Jw1HJsgKcVWAD
xjzBDcKV/RbNRDy7bajRgzwRbci0qyq6S3CU+KwRtY3AmEBiZU76drkD5MCB
3uIhss6HLL4Qz/DhybheIgiNSqLLzI5OlzYjaIIXusKb7uvcTTzK5ddF4YBB
Vv65qgw9KH4wmPQArTJXF30/zTZu5AF5leki2t+TOKN31A3FfaAArecS1YIh
yFQQpF+6Pu61vAtzqOfPDhxNYioRtbJfVZUpBgnkg/xVLsuvd6xkreWKTEWn
YBfoH3wjJ6PBtOo5WAI4d8LyIrpPwYTjQiXKy7ED4cCK14xd7LrmXBfBY/8y
RjYz1K3nfMiKfVNzU2zQ3jlKBkQCtibe9Vq90KFsTyAXq+BfI0BE4P3fUk16
RZ5w1L0ie0YYkNz1cG4SlTuQbeX/UPHa037FD5cKFsqLQTyvfz4bJIBeQpsd
e56HGmUnT8JSDGb4KidWUXEbcCsG3bAFu27k6cRrJSqP5prlHl7E8POP1YaU
Q2A6rXBbhOtFKelruUWZOE2j0Dz1xHpPsegK0pGaap3ffHrKLeB3XZ3pM5Lc
lGqc35VHFIHYBl5/yS3vEe5bRIRvDEHfZT69lLtvZj7tnM6expgwLVny4eT8
CKj1qwcjj+YA/i6Co3erwp/8pxplhPJ9coBdMtIs2Tdc3yZhJhXx7z87ozO7
AcNFDnucmsX2RZVxECOoJIAw0Si9vfcj5napDGcigW0MWWPuNN2dEkreFLZt
ry4GzuKaBXIwIh6J61iyepf1e80jj7yH1JN34cCY9biBPTeAY6/okDZPF0J8
9AgxX5t3zmvZNqEvBHmprxnYE+0bCSrHLPpeh//utvr2u+8BVXwNOVw3rZvH
bBLvjV0g45iReSiw22heS+P8jMxOOnNlSpiUTNN6VujWPRACDtufhcrE5OuN
4k/xZtlA6xEdxYkjXfEqR74vEZlamdcE9VvgRXCv5X/LRsIoXida/zMfJUWO
8gnOHelZ8iIOHTugicHMOtmML6ysmc1HOsGywQbacOPNCg0OxeT+82Syp08W
BaRrsX/wj6xjNiAluvOU1ZhzZ3MOiUQ1n3W2cE+3K0DvBEJtejOgeZdH3X6l
5q7DVP13Qp9Ml/cY9FTJ+B8HN3INcXPT5nv1npN1cpQzBehEkOZdy1Yp6tNk
NHDx0wNEaOmkGFXU6YNtDvDrhKQRXet+TN93KPVWgiUXWxH4317V2q588lgV
RdrZLwDX3jEbEsvMItFSSvMyTr18604zOAmAxA2mSk37EstxNUsEwok2XV0I
WQUBTBxbX02ZFmgeh/FZE7PSw30OjyV3OhIolkI5D6m9x2GPYAg64T1VpuMr
0zqj5shcxoKFn4t4/UF+ps1RuWv0Xyj50aFRa3Uu/GM55byM/8pZ6jYpDuNe
QMDeZ58gqUTKW1BsRZ9qoSgtU0Yr+iIMfV974xLlmViYKcTw3fYua2dZC6/R
K9Ppnge3Cnz4S/Gc0elObXMa5HHSJ8y6id9FmfVwb57ll+UWRBuKJOjwVRGL
Ky8TaYHx3Or5pmUObgPEa4b9Av3s2oHd+o9LwNuPh95ca3PDXTy5K65fE8tN
3bLEMyHdyEi/lcO6Hiyo+OPjjNBlTYQhBFwSF1HRdnwt5OhxYGabaCave9Nu
ScxzeX8W/rd2rH+Mab4D3fNMsVe0Jr2UBUAyNgJyfnMITewKLIMhmXzDKEPK
DTIeLuTsYTUCYEmk+THbkVjTnQNzl2deJFIsHgCG7faw46IpIcgdgfflFfCf
qObeku2zTreEuL+ILN1CI8upjbf1Uk0Eev1R0UHxa1gL25vo45BJsh+jCzMB
383ymM4xm2i3FMXxq47DdEhxgflfySFiulTJNOshoYW+xFoZyB3LzM+rRlAm
E2N+r3yt0B2f3ARqmFXizZ+zRQ1DrCIOujfxGqCeN1ZrIY+O/q5L5V4K6Q0j
YbnrGShCKqHyd3el5xsto5ResuOnUYOK3YYIHlaWCbr+nwtL5zejNl2Bx5Ju
kBp4JYBH5xdb3Ji6aUFrJKiNqp84Xg2NSTclZh5tklUE2KvPIfrwMytHvgR1
sLi3A9n3mJgbfWi+rR44JvUqzmYHEJCxvvpVq4eBUBVHdAUfpduHZkvOM5EZ
O+4+5jCMVf9jK8CVatm7uyQuq9dvMjSoh6lP9+gDH0NAqKlwBY7or8B74pee
RNErsdMMIsKHPWbZH/7k31gTAHSFV4W/Ow1GNvOR7rKPODiMo1Ujy8KkLVjR
GTk/uoWXstO0gyesyArRuOHQa2eK+l78rUxpKN0n7nMK6/+u09D+OjJDz/PQ
iH0PwpAuuGKZ4mu0pYqbf3h5p7aRVid95duNyYiQev9FizP+pJy2DAXCBpca
DEfhDkFOilAmUQb7dn0KsDJajwhFWnydvGZJ3K8SRns/Gllv661qD99jehIa
+lYGHAxujbtZf3xtiSkkzkKOcALcPWiHzXiUw2qjJZBm+bCN7PdxwYFCzgBi
P5zi+LwCCOmYIwhH+VU8Oe/8NloVRvV+A7grMtargzL4VFXQL1VXT/KMfPCj
fLJSGZePIAM/IGpMxrg5hmw3e5Ya/7u57EJ/kTx3Amyd78PHyDMkUGRU8Y+e
CDdQToxxsxxfyvrlWTP1o2zLtga4W7vfM/6RzEmwKFSTNiNEI0g53di5PFi5
/vS2oi5Id1twBxmKDXhTcb9fFD36c8deKScFL6uwf2P5dcu6JDNZ3dYZBOiU
Yx8/qWXoy0swHKem+Wx1EDjFlZmLYD2d/3kbTGKfMU8dcy8VdZ98Yel93e8X
/M5HAOammQPNsjaD+38sUVE1Mzjg0PSDKik42JAlcgISceSTj83rMcWzp4gs
qF02w+RTPwrb5Nl6/pA1JpYBll7v6DCqleFto+DEy3OTiUOAM6vgUPfSwIoc
0u03kY2/t+4cXeY7SBVrE8RIZ67EncSWstQNvCYysuuUkG1TTCamffbLajWf
Bx//czOPPDKah9jfTgRUIuu4s9aHWg6rCFv4176I//nlav9zWZuH+phaieqa
4ZOeqt5gM2P5mUpERPMyyLJJEg8pBL0A0Pgz3YcS0onL2NTHDDwU6boV+nRz
2g6pJuZoJEbXrKukkzHzFqebYcBLPA4TkmBn68eL7Loa6n6uVtaopkVmXHRH
ja0BlQKgXCBUkA6vgPf91GjpKLiahq9mJdKkrt4BEtuMO7rTPYM5T8rrkIsd
P+i5EYqAlJSySEgJV4IZxfhIT6bhTWhNTLDH29CeI4SwP6H/cYc5UbhMzKT4
Xwi7wB+mNalYRcXyPco0o8Nk4cBZqbBKgcmH6khHL0TwOKJCmIjrHzH+CWDp
PtbkRfzCf+IU97tPwL7QKmmrbUxDSNTYGl8rTv2F07fHQxz8NC2rwLNRefgy
EjzAO/P54uJvJX+xgbxjxnVVWINFUZQGD7r1rmb1T787ia/ed8t8wrcU+O9E
XwUsuo0K4FslqCje4Itcjc/KBr+jlRCtKR/MTdRMVrkqkJVgLCBxwqzIapBB
LN+A/z/dgxx1jC+7wRzaCGDJxJB1PPpJOYZiw00EJhcCH/97TiCjWM3B5evi
ef3Q0hxDOH81usHsSrUdo2CJ/47m7lDkS4t106AWxduTlOAsDAmQHhySHSaL
7VwEKD2DDpxCpBB4Fyl+nQ+TjOOfmq+EXoozT9FmsIaDoFDlyYFfyHwnGT86
3S/db09F1KKXKBYA3X/ln0suKDonxbSNjjbphccs2RDld8LucQHcmakaQPYr
/WdWL74H8WUBfL4690JaDNscg4dgwTkzPHNHRdyZFbUluZSBEeE7xBVukai+
0gHHhyssFha0kATTroM/3nn5XWYdw6xO5s8dlQgWCpZHNEu3rFfLuCiaMgIB
H3OlC0IDZHzaJZVgbQBes4Ti7dfBY4+wJBlzF8SVMiaeBWvYuMbHNMqXkx11
W44XyjtBIOuUIH//uLM4E3E2iW7L4kXxs0csbQBUeonokllmz2kK509weLiU
aLnD/Bch+W1d9VfbwtFYyHXhC8lb68NzenTCrszFAldNfLD3tt2NWttHpw3W
81u8h5Jsg+WkIOG+V7qBfn7R8yasdwvWf+CznSgzTIc94cTsrbMjQ6VGwpPM
lMSIGXCNGyRuDQnD9Nc7AlG5xYHQivhW9z9wB/XwrzUrO26Xc+fJFtP3KtIu
WOX4zP1UP121HeZl12zfGNmF8ZxAzh7IWMxeRES0WBuaCcIOR/bBvGn8nKW6
5pIeigKery5rQkzxNnmHowDVrBh1cbjb0fwNJLlKpueJkE6wZVwjab3H7G+G
Mq4pqcNWSwvdzrdLk3nObwez3uzFm8jiYLq4wQTYp0epC9IYSznueK09XAUv
R88kZqKXsXyqHswoqKuAw7maHbfTxum1qxCvJr3LvQioEsYD1RYpIO5zTrwm
wZ7nhyw9FThXf0O1ohZzWKebRHbsvmwzupHl5jOmLXJCHOCHmjNNhoRQjVqe
PrWVJpXh8gwWeoI7ds4yUiem/BeGaQ/qTdrVcLKIpI3BV19bMHO0k4rnXKxU
W9mkDhf6qQJEI9ePpLTg1f2hfzimpdcv7KOtAA08JL7aoKqt2Wyrf55z9sEn
2vtNKzQ6h4GALiwNEiE0zPd5jHCdw0g2+JAA+yfVO0BVvGTnezAvWThnEDtW
naLpDlMm9pWScmR44byHgrJzOqHolBmBWrbHoaj5d0CwH4GnhNZis+G5oMRo
YkBx8icYRbLz6ceqG8XNn0pP2++KgK6dJOXhf638Su68P/FAdwLVnPnvgEUN
7tLB8GN27oAHm0bwswdzmwQZxWF/5nEQI8j9Q9WlLQYpegg+WGhrFGdEirtR
yPSddy4VPtLUcoFbVhBTM07+i1+tsjPbHNqiZ9URWblWtNmevAVT1EwwjsEU
uQk592yBxdF6HknpyZXygsGsEWcs6j9sPMboFDunKZxF10qZ07Edwso/M5Qr
FH216Gyf2QZU4aRf3ln+5fDA0Bm9Qzbjm9rq6t0EaIQWDgeVOq/yBWKEvS9H
p2Q8Br/Fq+8q5k7cYXx4no4cx8bjvcOe2A7xWdHeGizhdtzOWiROVzTzD2V5
6LexDLdmAyP0KiV9U4hQU+Jz9ua1ByM/cKRO+Tms3wxo4ZqU+EgtSF2iyTkm
mK7JSYtunvgf9HwiKgiWPzHNZNpb4i+OFKEO1MdH23Lhg2d9nLVcBmUq+NuC
9LtQbD5I2oEtRw5wV088BiABmu3fjtj8rD6YTVZkWfwdqtpEv5jkqQ/RjYqX
u1yaOnm7/AVKKd4bG7dxnkApyUrJz3neD/jpH+Ia8QgxzyOdmzNEa/Yy5yXg
8GhrbJyMchwK1t3J7GtT0myZZ/mPQFQ1waF8t1HLNG1MtX5u8GFje92REpjL
E/EcFaib+Ygyu1u55Y2oo/L8nQP1Fs1pAdwgJmRp3okCvJQFNPlRC83acZeP
rHvGxjDPt8a3MThNC0BtuEvJoeGy4a1wjzYhN5bFM04rFzkdwTuoI/32385W
BWNCctI7EQZwAIs9xS+3QHS9Crcg8LjI2lOs9+Sb7IF7B+MuJe9LRdu2R9rN
RwQzkUQr23g+ZXfvheBN6bpLSBGgNbHj1OkXsR6/pVuvhsx+ZBVK83Po18TB
Euj57yJzKlTHmA7VEdKCtyHeay36ZsjiUgW0EClV6aVszicivf59IR7GerrZ
GfMSXmv49H9eoeb8QdQ3RzATFwBAjdjFErh79rVlWNvz73HA5jpC7h7dopFh
nkCC2Ju/nLSiNEmWAdB2WvKUKnt6bxntItr3cy4BTKpfTuBbJv6IF/z4VfHT
9uE9qaHpSMfcC65wGRCjqZf7yvONGUYE9rzmUJ+7LkU8qYWy95W+VUYdaqpP
+ZtwISe3HLZiL0UHuXSDkrX7RkSXmT60DzsgoxeCFMs+OH+CNIhkRCCVTYst
P+LGW14K1GH1w6XLRjANaIZhzByq3i7HByDyJYL4+V5OBiZB1F/Xq3LpRwKD
FRCGpvQquxAJ/vO3oySQycpwGxJyrcrKdz7PYUPF7JzEHiLm4WS95is/RNHJ
wbSOorEMFt7E/CV2SbLpiOP1l0wNmDzhawBI/sodHdOIZtQY4b0W97Z+71m/
jQ6AAsVdY5+81fqGZibhowe2naDL4l+cQ6gcBkRgnpM9aN9Fbj6alFz9gulU
XwxjL7GI50Lbv+X1ldbkN1V4DUfc/Mkwj0G/MhTFCSlSLJhM2mpdxRMu9mNi
cWQCax9o56S8Yz6b1RsJ+8RPRwAW07lk9r/TQlPNafJwsp6k2j7+HlXdh7rX
u05Yd4pKi401IizMhLQCD1PyLGipXnPZVtI4S+YJg13jv+6y41NJwxcF7Grn
T98LPe9a5gA3h8C5a3raqgk4hTqggQQO0eRMABbctncSLIMHAVuBsIdPnlJE
NY53qDtTUkwSrPQh1dU70sTPoJrZIRKf1pMI6sYbHY/ICSEsc8v9U4vE7pkv
8lA1s1xtAad1iKKDCdzcUFjkz8I9RHimD8RWbUi6R+4QphVeu3OQDqFG3/Q2
Adh+GMVnpo5eS8e4BrpY4c/98pmfnYtfzDwr1pc1WUT1b4cNkpnx1aDNyPPY
8Gck5Bxo3zpsHsKPoHwJwiTKN7stLpB8Ex7nMFHcroQMoIYbWYr+KBeL1pIU
YDawWcCDGSDjnwlIFewN5qRxsx+U2rhuj1RDbZoCaRik8S0246MxtNNmxMoC
cVQdjXkqdZ9xQH3P6ogJW1p4y9fFUsPxU5BhfRymqhE84dPqaYid+Dxc6jxW
eI3eynKJgqdOZFOEQPSmHPP7f7Rtwwq3g74afrV+q2ueKgTveEYYixN6u4c8
DI0jF6cpsWBTNXys6sebQbkaifFj3S4rBhNlA4o3AzvfANc1A2YPi/rwKm4d
I4bc6UQdlcq2XEU316UJ5yPxz7p+K4s9gciDl36t2Nup41O5JYjcpmhZMBGK
edb0JmePYGv45VgAbONE7HCMK2H6IQESSiAAfPXkRsgtQZ+2koOtgmrgcYsX
4ddHpTk3pCwxJt0rqWeB9yPynU9TR7Ep7SXDt2Jt4poAB/N/Mq3PgB4TpGzR
L5hY5AvG3+OckAXe8/fzm/5hTeOa1/XltVblF4uBPFVMTzbyf10FUO7O2uKX
RBqY5yt/NP9yzs0d/0UEWaxvZwR6kjsMNSPAjNAam4wNdfHAoPpnB4J4PRL/
zpTEvFsHvWl990Q63xxmrFfjCl2Q/ThEO4dLz0ilVUiD1PHT3q8Urw7NFVsP
3yqh3mR0aZlppy/SM6s7mU1iFFICWx4T27DE2MVV0b4FDbsdTgLVeZrQ7EB4
RfuKPuQRSDu1I32KqVq4QjrOeiEQsppqloDCFWitdX6ZnPwz+V5O0+XSwe6R
iEQp4CzUCjmrgiBj4x1SmzEGejQYJgaRHmNxpuvAkmQmUL7O0Fcc1bm9pV7L
GT6pYIlAlFls45TGaSQt37SWU14bF37viv0mArUdQifb/6pHpKF3+KpBgWC7
k3LXM0y+kn80jx/cNAlqgcYuVkvxKVS0J/R+UT9D4FoZif8/yQkYJxbJGNAD
bc45ZLHsS5pfXCs0kqeBhdh3eMwfWHAPHH7eZEBTAI0euhATwWZ70X8SnR+X
8Txj164z6/1T17aG9gOQilFIsRMydbf5m0mfU1VUCVZl4CujF+Lrfytzn4EY
2upkCGGmW/s1aUOKZbiGh55JJ+AORRop3O766r/tBEdbgH8eGWfsZUM8DGyb
+mrqXx9XNvoON6mYhBUdwMQQoGzn8U2KOBzWzI+MkW2g2goI+lLEADP/mCnR
Q0Py3qfnUPgGphXDUuPYQ9WDJo2d4oOzI7EF6t6cqc6HZ/XlaRjf+7vNXy8N
D3Qz1XbvbgX+uU4uSvti49vGO7lhtQScr5XJUZIanpN+BT3NKLjWd32nJ3Cr
/AlSrGdKrxNabtJJSiq64Pvx61APjN22NI2wrtqbtTIbGdVvmwN3KurPWXzU
KAXHbIcE+CUF+q90W+iKuNNKrF5nu5bTOeY2waVvxToAL4ckTQNR+PXLvQoU
UTxpwuqEl+sfza1pG1m8R1LiOOD8ByivoIETUJTm9US7L3BjMYOzzjSh29N1
RapAgNDkrI878HlXf5/Bs+xjbckDKy1tUMsX7XoFDWV8jq8lNenmDluoCQhU
XgJILYMcVe/P5C0r5o50NjsaWOFDy6D1CFtI8zfUD2z4kpluL0kCvcX3++c3
I430USVD3rfsSg35FHtA2rmnBbTBkallj2NdPbjWp0K1Dz6J7acBntEu94eh
DoyPpATfWMLq4AX1MEMkQ4nKOsUU1++0SxGzrQn3W5T1aVeD4WviN7PKHaTY
8Klj8/iYQBQ8OrJyBMBDNWVs8xhv8rCE0wHuhapsxwGp02DqbkiSKmd/1DN3
pVVUVWgW9yKdgRpIiQdacJeZ5nTR1aWfLydBCanvwVtOF+yyvbmaD4XjSM9A
SCAphj8wl/pXqxtUgphymax4MICPU0dTMRW0sxTen5eA0EIcqHTM41+fHpCq
IEigx+ok8ekjJXGLNQnI9lAw/IcGDJHBdmGWcsHh52nm8RJs3Q0zxj/KIdJ1
7bulhM3Oh6YHf9zyS+lmeeJD0StUUM2Xi3z83y6ylpbdjarcI98ieFPKtx8S
YfikKZBm8uk82M61WlccptvNNZy3jQQGrJvXzboy+UZQXaCo2A82iwXxT0mc
xdAVnCrvjhz7Rxyt6IZ8rlVIBrMiuxPTYoF6v9kfQ3B9iVF2+bp7IFcJ533l
H4M7Qz1vLh8YHmgOvhvuEeWKHFA169L2jurNSUbBDdcAXx8jHoNtgDB/vSV2
qmv2cFc5V1D8nhO2GJK9Bzre0cAFjbzfDwCBFSLgYkCEw9a+jPWWM0jjd09T
eoJflW3STZj/k/+SKSZp7hftDbvpJ8L16IsHtonKCpjLyZm8mFWpC/laFeTo
UH47Kxms0xLWPld34DPS+GWwlJS6AvOspm7IKMlzHvb2+ZLD3JAmAH4LfrFR
Rz6/RudmKDGgJxx7nSs9foC1dB3OW2X5C5kBLdNreRM4IcToURdQ67lhb/4T
RmvnNoswxYlyGcjllVafMaGPPSD57PjVutw2m6daJdWMTFuKAARpc7Q5v2pC
hRThuOuf+hbwsXU0EaUAflmVAdPXxPu0ZQU0wzO8scG4cFHeqkjCIKpxmvkd
VIaaa3WwlaUO27yGqefakgtHpVeOhaubIADcuyNijW5+kisRA3vgDHRWaQT8
LIdVBmItIJdadm26qj9JVnVVwtScwveWACeEWXJPMxztwEthP5LTh4IPdpWG
uYZ82ldXyiEuMpvaa3f/OnIlbmMIrofcwwZyv9p+DvJqnkwk1XWCUleBc9N7
vVDGKHaVbnf6xgr9PGOGAXEtSBBjfz7mFxmZsriZW6EUTwplFZZxtfjQh2Aa
6nXEst4T4/RXpapw0u+RfxfS3sj9CcsvWxg8bCBkCNEDNO79LwxYdLap8Cj6
b+u8Qomu5yVZvXiR3f2RBvA+pE3EwBSafZv7EJZmE2k3Sf7kYUDMXZKn7wfp
tsNUoxE1C8UHNjPcLfLfHTFlBfE/HMwBGPKSaJesow8wi8eGAmiIigaKf7j5
M08S+DbRcErhNpuUISHJXhj9apk7OmWHiZchEm+PGRsE8UXGHt/xs53taoKr
LK4p+FCaHqQ9JnvMQbfsxwGMEEKJqF2Wuz03RVPX+kySXYrx1SDsWlroZiW2
c/tsTCxJ0p+8j6W7frI1aa8dDC6mhGECoMGr1HMOVHrf01mpJOqjy5VSvO8p
HOUaJyd3DxB8zIqhupMR4pP+XP0gRypgd3I0ZIZ/9X1IlPQbQAki6JsEb8lg
J587CucaXSr/C1gkSi24oepv6y7uRi5NkO8jMm3pQFyP/AYYBLmu/U3yjwh0
HJhj66f47HNnyewNowZ6W1HlrInCBrc3eH1yPt8wjNP3ZMvaDZ8qcDGAmcHI
WeuDr1dnRqFYcUjh9S+9FBg0rhpSKZ9MiQmCKtBUujp62K1YDf7RuUIJzBYG
I+YUIVXaiaAdFPn2gsxAEtmQeQ5w6fh5gXUsWbtJb+n/0X+w9MixhRkNEOeR
PmVsrY6h1wUpWKDIGnFHzk/VEz7quIhtyrWj4PPOsc2aQwPX7YSailLK0HMz
W1BOKpWwE9SE4xxzHUKe5gsFpS1/VApfHjhFnGWJJ7uvFKg0yfCTpqVZo5sF
eGDpuu1Agl1pWQxRyZXjunvtGkwYto2VYxKK/mhjuyJp3cwF9HhmKtXnhIyC
yleurRJ4s24HwP/V2mwJwkpnPBFwAIJ6i0dH58eTf/gTq+HWeK8RZLv/PpUB
OfprQ7H+xmPgRPg+XNZFYUL/qGJZXWpsfZxZt/E8Geo/weq19umx1CmtfQtQ
t/BOMfM/a5BHr4dcWRztGMJYn5gi1g5WjKdKXhGPctPOB5Rp9tfMdmy3/ZdL
aSikp0/lPp5xFyMze3NR8MqXAEO1dM0kEaamJcKuTv9RouMChyA4n0kJN0gK
U81fFIJgVeP6tutIqCHlplt8XXNPTgGkNGe043fdxgIZJorABwUn59YqRuem
2sVpCAj36yEQQcD1LUpemlOkRGxUomajgfmNj+wZ+qzCIKAmiYAbjhueS9Ft
2VZKPruv/+QAquJrL1E8sQDSuqcdyz+cE1sw7h6vqMHDdQW2BEQBEPmGoskp
Y7mDV5d7qwYc5qUT/Pz+BweTVLHYq1UXp4oCkIzBsFuL/Ill/MkVQzoxmvl1
YjewOBN4yjFN0K3xEIuFYcZDGkNsC22G+4QSDGSkAEhpKEnOwz/bQ1X96VIr
PV0GQnrKY7Z/LN8jJP7zg5REjwENYW5ds4pGb1A6O6/aYztlmnhgR2b1kCwH
qi+5CNFagYy9DgOmFROjPN0TpqaIOAWjZMUwZyuIvomfk+0deukas7TB05Km
ZctieSDOwG9iYMOyzeKm3jmVjQKIm8+uaE6Qyx4z3Y4GqXrpJv0h38OjdCMi
c8o+u5fkvw7JhDVYrr177M/eHGXz570ZQyylJjjGZnqBqrat4wmP/2qm9P+K
oHKnsR+qwAbP/NDjYd05HHp0V8vBMeNjMBNB1L/bPveK2+0ZIVyM2na0ZluF
6EXU8twmuuhNNlwyva/WKD4Gm4g19FnIjLj1v1EL2X6ImafxcT4yZUyaiQxV
EIdnF7nuuc4C4itBdYOqGXUuZgp7uMMxFkWfY0tNs5JXjQYVtMwj34oOdYUm
7RvTV9ZojTp8BKq3H3xg0HyOQBa7osqhtmWNgaxmCNfu7INEvodkImDICwK+
LGO+uuhR1IBjyAjGcMzeonFdt6ZziKTBGEL0yNPL9wzD8QqzE2HzsK2/1Nzn
kCD70I64t5WUnivtCj3c7yXByQ9DSZjXceVsRs7y7CAIN52q930Tcjhu1m1Q
BHmzMYp0qGsvdcYJiQ+/NFy6VtHU4m/h3vjkvNzuk4wvTNb1L/jX+oyV3Fn6
QHVMMP60xqDivijQlUvI9hdaWxVSLKSUu3wRqQ9kbi389Hgr3c03ASGpbXUt
H00CcoKBUPpMQQPgEnv5wFiJodOBI1pWmCungKrW8C6ckLR+f4BmFn3kRH3y
hpvqpySmcTVivk9ceR96Y07vPdHx+CWQmQsLncsXSVGC4XXVswOhh1FTX8oU
d/iTwlT/9162VYQRtGlluh7SPwKFFwX7MtFGMYV9e4tysUD0/4+a9Hnr17E/
VAUiP+lh4rXiBkYwAX1Pz7DI6GSqpRZIKpY52T+CfjY8Vwihz2TSFn/PuzKA
RzkuU0wR0BzkvWCgoUTUCca5qOEDfL5HLbVCs0mi3t1TmhOrOEsVTofD/0kQ
xad8TvoOq7V4ddiV0JJn1Hm4rV04jvSypMjNzpu/kqqB1736WcxirHC0FrVG
lBEzFuKYuZlSRAnsomDWdBQaSQ/tamRWZRzw7Y+JBey/BRY66skRO1WN1r/r
0H0p5LxheUVgba/ZL2z9eG8oK32lOs/3OKkEdq+KLTomvsr+lbBc2Uj7Fv5V
kLm00KmxroPZBWgzWB+EqDQaTaHoWBuzizScQAtPu0PjYQ7pa4D52fzEDtms
Z25aSd3J1Gy0B+JiObSDA/4WWj9TqeGO+wasE1dMcTCutzUgzht5J6pwwzBo
ktP7nSJb49yXaPyssJyLU0lyhmHCXvvE6E3ETAMS2wgK7y6n5w7SturGx6pp
KKtBEbOGp3OWYuCCh+zhk0jCQf9uxmJ5ZJAdVjKrQKbYevOiVES9WK4Zf8rI
McMxRur/n1f53E9ggDpeWkSl9oKavivExOHR23yRuLOEiBs3t5VPSw6XDqPa
bKZ8wVeg/FbBzOHm+YEpzuAl5Su8lTq7Uohz2zywxX3aIgCX1mz6RTM2w4Qj
QrcaqhcNWPSzA0MnGgQbpyLKcjxl9/HlDuPhAFlPn7WpezeEe0kkUPfq3AwW
iTUFRdan+RRniIVzoshQieM9pBnhyPUQHZ9sZCObLYkH7yA3buwvmqBiNhuy
rGgPWLUyuC4QuFuCCBkbhxFz4YZBnV5f3nx/Kvw5GpI89Y+RtJoAoZlVlFLb
LbpW7/is6nelSEYvj0LaZiuEIRZI4tZ4WX3OK8GGoxlEy9uNqWWj087O7Oui
zXIaeGp4T20JYtlgc2LemLBPLAnfRJfE5+J/RdErRQSjlT69GGNIdhWFLHB0
17u6j5GvxmXM3eE3BRcYsZhRDHWc0tUIFoawIJvz/dQzCnv/oABZu4RETKkD
fwWTBuCcQCAaoAiO2gVE3SUakBaSqLkxp7/0yWisic7P9d/mroCevAxFI+Vc
Gq+GE0cqaCrNmUgIXtekzqimUqfptsfUeHKtYvuvTkBRHLSvpIwLVpsrI9Ra
W+vaEG3OgIeiH/G6RrEk//LUCZeO9WewBthYzZwvpGCHfJBROkOoYWQ9aRre
672doH6OSJ2HzG7zD+eN2cVOLsAhBaU3kyN2rt6Zi5Z5MLtwAUduiy6LK1oI
HmsBL9paT3KebExzBwW0Ho0OZ1tnbuXKvdw6a4Ee7G/vx5Y67n0VTzYdUvL7
UgYZwyR0tyN8vVLuHB5MYS3DQL1OAeWOwKhNXQijlkxBSLqbSTpWRIrcuzr/
fp8/yarQKv3X2Z8cRPRMWSjWGrIrp3WZRnS1kT37SLw6oxrqzwHYHDr9dSwq
SidvEfBockcMRoC3zQdtmbFM11UfDhpY726pnGI9hqmVdYueNtWEdjKqAEk1
ZBzVXj9SIdKNUklW0387vOByTsOUpMaFK/cLGtshy6k69+uKP7tyuvmrAKmQ
HPiFy4iJxYVmcKqf+fqR3NGOVZPybgaWzBGpZVzs72c1vKqWf4ECs5huf5Vp
Q2kt1CBBMeOxhrP9vyQHMcYlVUUvq2EKCbM75XBPozWjPV9sN4KwVBEJXjLm
q98/uxXBH5gnTbysxWHeaW0HOPFuTeF2/5sQlOhLDW7kti5caWZv1ybu+FtR
FBTVcVNb5IB62fJXvN7kOdNSFwu9K+aeaj1nkhvRabreinWNJQBDeYBlxEY+
S5TOEgXNojz7fLm5VH2Es06RKWhdH/41GFS360qnjSGmpFO+AuReHa/qNOdT
P0L0X2/CQsxTKVBTrwwxrPCvkVViTgVTpmADYrW0c8vEFka6Q+rPUsJp2aLM
7IO3hRDJwD0lowPhUkppJ0Mfcm5Zam1/LXRis4uBVKV0/W5wvJe3LU5lc+jl
lw5K/ryjq+DRBJfTIUGAE04Wm7sANHINuJzlDKROxwhSfsL+lzD+0JDnSBY6
dC4QxRpsq+bwt85RNo9O+pzUepA6CcKNnhHETg7vPvbIq6OndQRMw82caEaI
ZInIx0wejCb4H2lEFBG5SIk7qZo56LvVHPP03cqSHoW364HwiQhJzWnAge93
EdNkioeWN015VprVAWaO0xEs1pgx+3+Mm+3oCB9Mh59XLP98fEgic7Yv81EU
QUZsMg7r30BfZYbkurirDiangFfOwClXGXQEV2qnplggCT88rZpqJ2AX/X1W
GQwexnEcaqe62y7q4sqW2QOYHkLsKwUMpiTV5l67f2trOqsBNQsI/U4xTbT7
MIJTVwAZl53Ffa7MomQhWPloeNeNjknHPVhk24QrUzrMl0CPx0My+mggr8qX
F07ZVs5FGD3wn2JHZfJSpSH50kCqmNLyN4gE7l/kUXqkunBtjrC8AR5dzS83
x/SPcJWZ7OgtsH2jbQdm9oXk/qpqRcQFYEGOmJxuU5ZJvP68bSQu4CAFk/uB
//R705l90Whrtb/wYy/EzI1NRDPNOc7utB+gtP+IfYtzyW1xGkJDh1eO2rFn
cmY/+QQq89m06p+kIWKJdZiQWa27M5CzbMIUx1lE9DbfDxgmdgKm1SngNico
awz8/fKStMGq7tOyjF0OR+2rKy79urlkFRt0eFLiAj6Muzr8brXiX+0CBuhc
QCg3Y24sAOIYdWzzx8i8Gy7vX+iswSqumribsT0Vi82vaag3a79n0zvI208c
r/75YF+SJL15NH76+ijGkMskkRiwS/4+++0bo/KFs8AtQ3fLqgX1/iiVpM0+
lwdhyZBAaSXuBJbwq5BqY4oGNKgmsDq6v68E+LQ6Wm+Pm1WYh9i3r2AMxMtm
w7f95mlbAuBX3IlnTM+nmMLNXdpptffzXNN4Ijn/OGaadANU38YIX72WKw/e
BTzKI8YKEfYKN/LSPRlbULurE463EWPPzree+XwYpuPQgItwb+ainEEXJ01E
Pz/P0JrftpwAc7V60IKZzmguGusct9qnn5lRrZMZy7PdlGjW0zXB3kFFv619
AN+a6pkGXGcln520LR2oWO7wn3qtW1xhY39xdV0Y5CT0vAYtXTictZbiI/nB
o+LA4GrmjSmAWOvns3LGrjdaya4B/OISd1BO9QM35iHy++yCtmqVB5t1VHMR
z1YCBMNPqXZJS2WoVAeQ7V948/CGGb7Qqg0/1mmQE/uBaneAY1ONpeMFdOFr
E/hA3MkfQ+Su0b/rZOs2ygo1Ouu8V45WvPP9WAQI9YfyTZPhXea5K7eVtRSG
L6dziQahZS0szVENoHqFZZ0vLnN01BTv0SHRfzYxDcctyMD6k6oz1uc9Eg8d
nbe++kOx8zdFtmI60nZBJfLFcchJ67xXyF8kRMQTOl+XX7vaNmamOwIW+Q8t
Fx0N8ao6Nh0zho+oErTUzCQ2I84j+ZDpJMiDiWaMNVMlPPUhx0wWeJs63zVL
9GPjXRXClT0RZvZxLUr4YBADroLUsqvPAY78x1/9AnsUrRrhC1QVm1iznAlK
oqpjwQreO6SQLNpcU8KB3AA9Afs61TXQceoACaT0PmIe6jXm4HNXi99gqK46
Jl2NO/1z1AFyMoAPBfoRMJWzGWmjmAlbCAKIcWI5P1K6bvMu1pI0EHaTVUcs
CbdYRjwBA1SVr0LaUs9a9I58G5Y1hD0UPSGLaowAeJ8m0xnrlyDKAaoxNzhT
ikxJzhrl9OduhG9PrBKS0jD6iQmfPxpNfjXepLlYllklJq4cAgTtUCrkSSvD
wwjK+cqmlPNTWntsi/yXBQ7uPaAbxlyp71Ac6RcIeYsyRJQ42VJr9dra3q3C
+d3bJmcAleBi6Cxh5bXTsgLTVGY7Cmoh9olSaaaYh0ZSxBzx+fYKrMxLXbBe
qWoPK5ldCn0r8Rc1crB8iY6igHl+ozQFTmwdBblga5QVeqhfAKHJwG2cB7AL
85l5vzA82GMO5TlKODCPRrxP5tPfML8+xKSg+dFCaej2gq3VyOLrV2YYp7ed
fCHZl5mWsBNkoOsw/6YKK2230ejCzzG1TrC79mtt1GB8IGGOWtD/9JNvaSK6
OG4I/E7B8+obleRdENboz/PFIIQrQFFYwyi7HT2rPSGbWsL7ckZSQab7VrI6
f/HdgYaDUQAH1QWXZq2OayUBwT/FvopjhR+JG/4umlGjb8/aXTaQs2DkxZIX
+NNmIM4+tunP3Jpokz+JLjdUEYf42BJYpG+YN27kJD45/PcEYAr/KgfJ28Go
UMGo8djLwQUWPaa2Ul/SULyDDxLb1txa4c7myPVUrdDAKWekR+KjWNrYfuzB
A03M4/FnZVRT5YlEdn/LE6wBJfB8cVQY9Ol5uuFCosA37w5Mheq0zoiYXk4P
8GEYuX197mt3Quj2DHSKi7PftqrF4b4UffcTMZwNgESeKBl/JSy91J0ohvAn
0rrOpXveDSSl4S/zFT8cX5h1cVrOqdfwIKZyQ44z+78O2DHJ+M0hUxgZI6y3
fHrnSU8IWmzrl3yR+lG/wPwBX6kXAfg0sUlmj96bNu9WIC/4vVQ+v4x2iWMt
WkcPfoa0RCYxAsuaPSjOZd5zAE8wtASL1gKpm2rA5yBrecc6iYCC1vmEKsr2
+fxkk5MC3aMhpqZGUhjE/bJ0RQBIG7PNgFLbymCpDD0v3WUL0I+cF7AxvTmk
V5qMWT3QJI/FNgfaTLbqBhHqkpAxaz6E1qiA3loHmZ9JC4V+l57g+tlAkVRd
S9SqQgk2YMrZsg+uvUp6EM1JIVX+hIw/M7sAP8QuoheQ6UNJTuyEdW0MBodV
qvhxFA36XWo1X2lu7IWsmPBXrI+xBjdM8o2r6cRQGi6cQ6Q6Fvjk4DBeY5K0
zjcR4bPimC55auiFgFsG9BYLIY5PL/cSt6zhrV2VIyZJxPHQX+XQ9uxqS/Ay
JGF5kI94o0r1J2nj1qs8xJhsnjwiFBnqaKd4Cs/AMvkbmZYXX4QzataQFCjW
y0m2jS2wjqbtxdv3VeDXAHfGuX6aBR2xwH+pWRwOsAxZU5X6srSyTu/Ocaa3
W2ClT5Bxxx/EJMT+XwrzzjbxbGFJJlaFpzkEQ70RseFaGw3oa++H5OtefKe+
mDoyyOrpHHQxqHPQjt6vO0vfYwj9Y5yWtYPjrpJYkXpC08rAlcz5RIEHrFPQ
7xJpukTnVzCB6qYMEBVAWbM6rSqH7SdCk6Ew60EFnfjJg8rfsx8boQbKkUnQ
FPofkAT3uAtsVTgwYL71YEjMMeMmDfI49SLY96dK2F6jTuEq/cUi0c7HhmCn
f6r5YFVnEOWiXhsill2iwQVVvUJll8DZBAF3T3Mzqiot4vsh8SngHtHchM0V
t/5Z7mcgDzZn3pEELCjhcFgOkqaIOrhyXhDor+1c9XxuCndPNpWigfkA+6+P
bUWCgJ5EgJWseeZqk4dnC2cs3BYJ0HTskafG83uzAm0M6xWNHUVQs8Wd3cSg
dsGl86d8qFjSRSQfkXLdOpanlPjTe/MP6f+IxdZi2PeQYHeRBvuHbdPbFIZf
6v6dYnCqx9LGqrGlR3GzJb5yZUbMvsCKu/mzGSCfljLBYjyI3LLLDbQ9vlj9
gR2gPrOfRfaTZ1WPZN+Qs5sRNqP2b6iZpI+T2J4zxOHNGJ9by9tfq9ighp4s
8JhG3rarwJHCO/f0aTM8P0tfZNp+0pzco3e77teViomkq9xBg2t3szGfrMHe
U/qFv4FWYcfjP7jbfFcDU2MqJrDj7l+Woa44Pp5r+/qi2rh5Db71Y1IzKRU2
6cP9nKJ/omILf47bDiO8jrfXrRsQuNOv6Qh1tFfhpBB8BndNpvLBjicWCn5N
EetSd/5e/CW0Xz1jgAMyjxEPTDYlBlzVeb4KhE+YfAlHLQh4DdvEbHlD/Avz
+clAHdgLX3we5VMKmLDtCsajGz6mCYFGgTlXkGT0dSKWKi0NrbYK5FF8gQsy
XRJChEx5YoABm1H8l6NuK+Ljma8m3E7wNu0xIFhsULib6zOfRDlkoFmTEJrE
Tew38TQoHNX6VKmMO0WmvKUMKTsLhscZzFhxm207I2/ATJHL/OPoTrnLTALu
jCYf5RmaHDXtvYcTKMqGXbzQXRvp7j3MvIJCKPR/JeJE508lbEAWvd2oRulJ
NpdI/OyiWb//PqiudI9l6IPeXFUOY8yAKbvtIuCp5lbeZ5rfr7f8sEnT3NKQ
27C870+m04jW5JAFl75IR+jJF9fiEKijmHqU4ACiCLRsHhmN/6PFpbA4vKuU
QDMvMhCGSowYBxNqpBjRSp8yFuEQ1jGuFIV53YWJcq67tjVIDYNZm3AH4f1l
P09eLwEmlv8xheag/DFULroWre3broYAc5GadH8fvLmCXXnJqMpVy4DGflZs
gkM9jAdR/6jSLnfEGLq3ndyAq94igHy3PTP3oGzsTOuDM/vx4530wHS22Jxm
QkK0wnCCTpvp3r6Epb2fHyC3zJm6A3g8WwVNOcEMiNMcr7iWvzbjMewXL5T2
IogRkzNr6tnrjRiPnjge10ZeN9paW562oV5agObccjQyzAjb1OzX7Dp6IgmW
Tu0rJToV2tbGXQMGpmseZcH2igKP/85qyoL6uhPo2aa9/fWdFSpPvyQv6H0A
hs8ax3g6ErTNtNrUlTwbc73tNEdGW9cOQwC5D6MT3UIx3QHc4KS+KGo32xDX
OhNYUHVZYD587KxluoSc1ZIex81LTYGifJYW1dCV+53PVsVa8LUijkLrI973
XY8PEydKGwMvvOhaqF6hXq6oIDXk2qN06FCqHH35JNfhfagVRIEBiqXeOFxn
mZWAR2caOEI54qppi+1B/IcMU/MNoRqYtiOewW2M/GAn3iqOiHd6nUCwm/2b
/Ynj+ZhWKjWrd0axtKByy8lQjLs+84J9/W+id80ZWMCkL5u6cQtsLQuxfDoQ
HCbpZypYlRuiXUY8gzJgTMSFOcGv4ytC0v1kosi5WkruQkiW0SR9r5VsFfxI
u++s+piN/3icYjfNElEq299pjfIRg8VXQJPJaSjjbisLr8PRrGo8cUP2naZl
pf8Jnnd2lOgddLN7wq4RsvBxFZxaGhpW1SQ1bchf2s97VXQw6zf/kKFCf2vC
SeuN5nA5inEgo2dMMrVIfu0DbXyxsCNEJRgBXse5194DP90ZfEVX9Andfj0J
B876YR2Pu7ZOolnBanNukzidNNYGSIMKNdajPxtSVMCWq67IitkFe0D66uXj
14gIVTj1oWc8v4cKoK8T71sjghDNGLEkJmusctwK/nRD4y/zcC5GXUSgjcs0
ywkMTT7SEgt/LTpxGgXeNhgtQ9YKBo6ox3yA9rVQl0kphOhrj9mCCcpkwSoi
Fw3j5OFqVYjWkSc1PJzuH5WIUOVZxg2L12bC0v73e9/iXPLlXKoRVUnHGI35
CE3b55fnpyW1NPreZ+9IzBYC312mYuzD38F8B6rEQJ/tufHUz2bxVcw1JLXC
sHrcZGve1p0hpB9OOJ7YS3qzAaTeWy4txvda/+yzNNYgzQDI1rZ7fbVWSGXM
JqZo3VzrZYyS2ZS2xR1D60K/SQkk8spSGT0BW+MC/8TmqFFtT4zb//Ixjmzw
YCcBHfjt8Qk8UNOH5hx1/l7s10fy0PpdHMsHPNpfm/l8RiIn3WNp+jA2rBgh
FI7K6cUW5s8Rm9rcW2S9LOkqqaG9sOwIeLS/P8qUxHt1kES0+hgjv2o+PPmu
I1bLMlCPMqoAoVM1YMPGWHwGtIjyPG//dDxHe/VEf/gJDd5oqG68FjsO9ZsL
Psw/moVRiF5WRxJN3ok+/Ecl0zPu/EG3z4XArdaGfd+YT7I6RMAIwSyo3Mn2
3EHVkPdfJdUaUIIZOIrVSP9Kg8FBNacDCBAdWzlLNGWEv6rQ7aLfvC3dYv55
yv5gsrOGS3rgTfoYP9sJKnvrhWMn0x76cGM+RkJzMeVBZUBYqeVXl76l+wCf
TteHb8hwhY92JDhesRsSMA6imwHDzt1oMTnUAZwjrzdFXvn//221GLUOXgEG
vS4TRjkZGtbl/gb6JbDgS/r+hPqzhkShY9ML52mRGvnIzABb2rnZmuvd4FJ0
rUX9ZyOVB4iWGFBaErfjpVBaLqFbqSZCriSYdNq4iNWz/KTbMTQ6oQbuOICo
EoCjUaxXkBiFuJBte/6H9R3QacRoD5ykBmtrBegeOJPgnN2BhS73l5uby4FD
oYIRHVSmHHbelEWGd/wW12k2eRaTnkaiijOt5irqRGEbJveAYe8o8W9kGGO6
CjpH4tMtjkzHJ/dNO00G6M5/XVUXO7nTawBTXGewGP7gIHAXXhaFiXjs4i0S
ELVfCKAIYrnHI6QVJR1qcVw+kzZLZ0fv/qRq2JJm/Hoxcia+pSEYSDD53saf
j4tvxAvEMCpOZxq7sgjBYnCRcKeEAjbuqaMoI3yjWm60cr/ljMgA4lzqK7mm
A9+ej1ae3/rE08p+Tf/Q8R1N7MwYGOIxuj0q0s4P9aE9cBbzjS7kl/pI70FQ
y94C39uWGgtbYShFy1ii3NQW8Tq0WrAwhaSDLCJL9mgxdqyztWrQvWkwM62l
7yAD+SjyrXXwJs7i5+uxyuHdl8iaWpM1dsW/dFBFSiIJOxxVrFW2wvFWJ82J
egLa7HGzKwTD1hyR3ZVWCr58HlLIEyVfM+rlzQHsUsMw8/+IrKV6msswGwC7
cqwuA0AtjOtjEmMjWaDuTfqToTmLy5YYr2/OiCQBBLdstlMoqVC3f9Lxmyv9
/2cidgKsCIbvRE0c5U5IlhCn6KDuU8HBuXNNet9dHICwlCJOh7ADPbc8bsBE
CL8wSxFwbTt0jK7jIi5asQKj00+5m+Sp/RNKFPN3LNUBJMzyP+pfn+pF/SET
mQpVT6yNReGTGxfHyMAa96V6SbaAeiAuDTVpXBED638d7Fv0b2WSuvtqqMux
E8ye65LGxFNLrKaxvcBi7/uE5PIKRahMNtNSwgJwWmdE2PB61qZN72qz3YoQ
fpkSR30N+ul0WXZFikhrXQ5e67p0nTOdIrkCgakNP+Cr6lupMgcEoHOkvP/T
uDLajCXE0oo8YqPq5IuTCK2fPZzTCnm6fQFN6FiuJtFQSnLCffcPopEFWMmj
M+n0Lchnv6ndMqY89Y1MzKFvrxJCbx97RljFACTXbabl3gYDJAIURx5WuztP
EhqFKax6WbAum6xTzZYNXns9fYPNFWgV1I9VJYOBab+WAmyOcoF5F7/GTDT+
OFaUjRtvNsklTJG5s+C8BV/2NlJk4u2pMf7mIpWkdzs4mCU4PyeCv5OBcqJu
LaKDz0nsydm28sjjhj32ypBy2xJYEvKqIfyh2IBf4JByAjTnjHIaLGGXU1f+
oYnNO16s12XE+HRz3hbLuC+Js7ayzmzgDrxs1dJqoqyUl2xDb7QG+9qhelNC
DrIRrJkPMOLDuZXeBPonbgh/WzQCTvF7NwIT5MqcEZZLWmwf8x0unGW8LHAN
XH7M+vMU1rR0JzFMFtYe/PSA712m/6T/gnU/i6hWM4D/6KBaQPba9zkYHXZw
mqi9mEc5Uao4YNMjduZItEnvxDi9+1McjcxU6osJGINjNpiOFIpvjgOSMMK6
rQue0PUzgm9rGuHPzQotNBGHlRjy/yvVWxccZMigb8FU599lkXst17Da/HGj
bbA5xw7WECX9pcuERmVHlzWzalbfGaDoffVnGybHg7/9uk9b6FbTL+OxlEij
tHoYakCHbwdW06wQSAUpy+oCwbx2czyG8c6WlfvcaAXbP3y8NNe4TC5EKpXp
yVZyhaME1VVbGuIayE97iy/Rnq/yEK+r8PBoK9HHlqftpbca6f8psakD/qzG
F3Ztzi+YoYFZjqHFskAlzVWmjvVrDdZxsKlflDJiTBBZLMjPu9Blhm8f+pEQ
QDg/KtL514bAPOmncEY+l2nUFXSSBTqa63TIGxYUkNxc0TxjMtgHA7BaaaSf
1gnxW2XHai57HVpIIHh8cysxRbuIbbIyYn1TiXkah5cEU+/6SMOM+gLmYa5y
mbsfnqdWOK+q2XSkiYZYKuDN6TGxhSVoKOPm6SBqDL+NXGXRRn4WVtFfzaI0
M+nEabeSBks3Td5DjnwS1jP/UALOunRNlIpYOWgRz94I//lf277aUbNKXyor
/ulC5iFG5XQf8rwg7aobHjizAAWjc0uyDtb8rvhl2087oZsEzufWwznUM22r
zPXYJWEf6N5YEgeJIliPu4c2o2RVy3B6rSiF7axXUU/Ual4C/ZwNiGzbmGNj
QWZxpt+zu91hCchKvfCkftOWgr31F/KXM9ymj4MyUjxC5ePi8RJEmKvVRed3
rqyP9J0axR73vEXxOo9KQ43F1bQlg628DeRIOAHGrUUpswK8Diio06gi6y+q
2CmWMVZJvxDZ3CRCC6tQjR1Wasvyj0zcossI5Ubx3Y2vg5YYKlp7w7WgTMIR
2v8cnzcIwk3I6ZJzXJvEfRIc4qzH1wDFvnyerHaUKA6zDQGmqGfNaOEiwC5K
RoL8F4dc7lQxjZVbALRqcuHGvOKQzD9PlL9sz4XQRWBLNA0A5CeAV8Asv0zZ
86SWUu6pdR7AbIbCmbsxLZEfMB8mAudEclrcGHcyiBTRWKIRjETDY3J0GZ9s
75MbFE8LbJzLFtgqRU+Vuy8EciDT+GInINwvZB1heAOIuPlyft7nMyW2cXgf
PR8PwKA4q0OxN9FNpxVySsRsucyPIiqy78I4WlTYDkx6YOgxNnF80dgQSSJi
i+2dJ6loOccUUzqwzEtUkhVoV2KySRQZnNt+OFzZ+3T6JlTD9r9Z5w4Auuom
mjYBlYJ5OkfUA7PQcmqPh7WrkYNsXXlFhKyHxoJk1q32ZcLC/y4sLrIAhsz8
ErbrY/yyahCgOJzlmuGHaiRFR99J/yLX9/dltPHxJyumsdp87U67fFGnUYjQ
t7NEomdmEupwujdy9/qvPRCXorpPAhVEn0uZyG4D2XQaDVYC2H/TFHQ5jBMi
BjGuTj+ClxU73p27se5jfDmNrkv1gZVqInWhEHTnKPZR4o9NyMzir3I3HhRA
yIYKXVDcy0wB2TLRJJftxj62RVWtyXLWtU8MTNPfjLVEtc0T1CCSxDnc8PpS
dDZBVzAsWyJUXFj/KMV0PfXfVE1V9PiwDKYar1Fb4D3nuu4+VV0yCGKFojDH
JBNxpmCGW9aIjYf7P6ulHv+gFoAsu4GWX0s8FYVyqUz0TBcGdOJFrW/MH915
QOTrlt/MwBob6U7/LY64+hxKe0IcDAjfj9iUB8y/VqJ9gBOCbLCPOmK/X+YO
74GBjY/onvPQesBvtp73KjTBA2C6W7KbHKqnhnaDUcpcOxjC+Avn8XM9u31k
ZMYjDevCHfvaDEkrhIZgo77ixyrPPy1oyIXXMf43AgwDEBsSInvllwnkd7ui
/hkoQXdqpOsfYQ4lnBFvzWFD9ownZ2nJkcP9vDG1ywLT6ayQubPBTDFKMrDI
E7w8+Aip7ftdkZPDervkwCWs9cM+BtcgQ8JVSebjFYpLMDEmtDjPJYQsylly
PxehzPLGahXM0evY8C4UBdbnoTDQYa+vpMil+WRG8grDZRu9qXOREk8mv/qR
XBa06Co8vdRkfpCvMBObvp8Mrrhifx2YU2lphFIMw20EhAMcUKDBWA5TuuM0
SfldygXZkMvBG/mGq0ZV9mSDUHl6/O+IuIH+y3sUc5YrrGIaRpgkjr4G9Ujd
oARJCdGj4CfWkDlhuvMTJ8VVYuUuuGKC2O4IiFiGt/khvBoDbnX97s/R1WvM
t2R2D8A4+7QSsLHMhzM7F05Zl9OwGE2DEi3N16jl3gUdZuML1nm+HtVc9AsW
Ntjt5EEn5nN72Li4eB5LDU5uAafX2eCW6Y34F0TsXWQiR+HKLqFkGtCkn//v
CrhM4/Zot8t6sM9hZLain2OFKX36UY37xxEhSmvCz7kH9QqnX7+oWBOfvqsX
SVgbw4VbUBYz9ZV9SPuFkIs+c3A9pyyIAMNYObJTCiZ5ZrUknKUynXlRLtZ1
OkqkYhKLCG5xDRcMWy9jlmNA6s1utgXqf4js7L/g4aa0I9Ovp2L+59YNz1zz
j6ne1ta7YXQnf1r/a6cOJhOdqEEtbqlDH9h4+A5bjOlvA73NovZBycrlbUQz
3bKWQSXcDwxgJbWjo+sJQEdKcTuYJ3uA89N0x0SszV3lMAyUS43zWTKKTJ1S
FN0eZvo+fzMC5beGPJxKKIYgdw/FFuYAqBWsCsjPpIX7r7DjEb4Mu9M3qjFP
9dKVnVSM+1No130+rBQLfBM6Qo9Gab1XdWOtyS+HQJqYjsU21fCPDekoTRhr
nRDkKyPFYSkeUTAS7a//O0/ScK8UfADog0Ij2KcRZa1TCbTSwgYUW4lWxoQC
vBro2W0ey9FtVyizlPlVvmF+X42w+xB1Kb15e4nsisjBlh66f9vQM4RYet+Y
MAhcstFwAcu3fSY58H2U/L+S/VhA85q1h5Yk9BahPKC6cx5b4Kz2nIAOHKfx
vfdqAuafUjqKRqrkEaAjZZAIzIE3MD8ov5FG/YSPMVJWHxxMrdwPbykdKaeT
6bHm3WHsxheFcPd231NOqhOM2P0VnOpFANKaH85HnbsY0ob2YVJryxKerkRG
b8oPdggMLKh45KkXrifKPYbCN8wjWrbm2GUU+D7YY8jBBN29rWrzUb/z5LCl
LyCmqhvOA6eHkHbXLHh7NT0HdSvQrO8Gf8gysYxOojwX7kvVYX3tdmnxmbOD
xUWNWdZmafrx+aNQuun9/FrtsvJJSW3OKkoluu6YOTC3APOkxyJhwsSmPEWU
kenWlZU+OJWmZEZbL7qjH4HX1227S+PjpjcZdbI/dynCLPMGsVxP47yTTFCI
gcxfqaYzwkhws0fmmhR8SIi8AkYt1DxGCYtknFQZUqQadjgbgfb/RmOMoDKy
2+G4fonZ3333lt+vtKRHzzKwiNX4XfU3E4jBl76xbOcqANGT3aiqWQqBQdn3
LP5w/R2PnSGob8rDLhFbzY9SFqu92vl1Wp1ApDA6WRbdREuNVGriQzWlqifJ
iX7/Bq0e9yW7j0eB0J1S+FGsqvyuBlQolcdKT1sCqL87UWef83P1Xl0Oz06q
jRgB95mAecvZ5w6y721X5kx5gZDWGxalpY2AX8GStEyiJcAKqKI6uecRN3C/
luX7vNTfeTVR0i7agozeF6aMOTBSPnPgUiuzKQGVb3s2QJfRsi+w409EHb6Q
Po3RYR3I0r1WJP3MvQ6XXrXwTdkxg9L43jT+HtbKaadF9sjNCco4JxntOV5F
t+oPSTJOxv2DibHcM+gxlRksxyUCjzAYeDU/zH3q1MgOv9xGNoMSAFfDwkfK
biYOM4avJC6C9+i4E0OLUnIYIgwqzGxdVOBu+1pRgeFYiSLbL36l+4gYQ3Sc
W878CDqMcPv2ECBOWHB7JlugAsLLM13qHWO1H5tfrteVQh7n6mLMqHfa7fA7
KkAgP1zLfPlJS0/6Fw5VFdVH8YoYlKOW3+ENPXz0tHPnIilSSYPGHQE2jKi5
m+Tq66adQN6t3jd+38MUBircE8WUPXz/8Y8t5a0+Uiusj+elLgi/s/KLM9tI
/Z6s84/KdF7tdTRK2xKJ2npiwUF/AcyNJ0s5vRQrnMxeg8sBo92zPviU8Jk6
zt5+5s7CcqAEzvDCI4vT/5UEjvdIigxs2/YScUFxZq7gynviZI4PX34vKszQ
6sJIJYUbi4F/rtZuXxaK9gBgVb1tqr4cOnozwqMRaNF0qeQBfIlbm4jrZpld
YbbbzK2YGT+MavoAJoRvCMFmSICuUJFOWlgoX2O3N+/rVNsQs+zXOihpV1m2
JIXtao/NKLoIGxmDd5EL6EEbobB+nctQI6p4OXkt7bDZKtuZ61H/n1CV1aIO
sXm5IGvl4ZshBHaM7q6TmKSJUwWYmxgu1+3tnbWk/NBx2pwwmLWf8siCkX8P
cXaPAUtzN9dy0xoSME76DurZLmqWv7qynjI4e5bbTkluP5rsMSCO2ZwRd2BP
aEfSiyf+ICajZ/GRWLx5T57gOppuIUMNemb9xyDhM74VcJJWFDByx7icJgr2
hXDvQXnGJmK2CVHA7WiLEwNiXK9GntOsoWshNAhAB4wafk7a4IhdxAuJjz7m
ZYTDnsOJ1ND7Wm0sF7ZZkBmEFIb9cw4tGbf5OUuuajOAUQdr3wiUE8nJ5kpW
nQwU6wZUf2nwWDKwTfQhUc6ImmYkVqSo3B5lIqtnXDhKBg91rhvAkWDlooyZ
PQQSdiVgiF1cnlTWjxIq4wqXl04sAqzW2BVUI2F5RkiYXUGNjQ/bR58Et31Y
q90PiLqiAcd8Xa90Ks76muBTJPrWGNqhNoEIkzLlm0U1sW4WfPq9nzSUMdn6
e/Xj2Iy9yzvyQdmNGi3EXdqLXeb/eJdoWOorRJc7wfB5Atgpkn09BcyjYx+5
Ep7Url/+03uEUesxX1/+NjmG8M3vAeJKWLWm0PjNsGCM5JSisnSv8kcAh6Xg
21RU4rfoUWXWGtNuoK3yBWU7Kj8Unp5skSviKLnWDdG3V+SPRHbUe1HG50iC
CMXWH61mBeYV0UyP0K/7VVXdID19JIwx/8SLWvxpnmJc5r8zSehvprqTDg/C
BcMRHlnaHAip9o4F/JCRwExv4syEXoTkQS3hKIxDYPj+H7vJh3dQF8FSIh9N
Q6zkyA4iDh1RW5pk0KIPWmdwKaA+/v89Jj/ywDcQJR1Ck199TqJKO0Y8c26B
2DPjuGr4C3bycR9dGu/ghCdVTpyuNbTJrTt312uPheOshMcTm8rryLASlW1q
we9CAw+ELKCprzkcS6mjRL7NGVKCLTIXHLT1/musQdQrcEFOezHQqCpyKgfS
uyWEmTfGoDj+MGuEt9fCKpnemo+CESOvXq249zh8cefBi0H9pdDaanju1rGl
ZzUtX44ZvZtQpu7R13aSlBFYOK0u7/wzHeHIJktuVouaWcroEaOMCbb1dQ6n
pRBsJYTFfwHhRoeZV8Jz+MHVi73I4D7CXAbDW24GqHwC4I/QoASOt4Fqs9wI
LWAmM7rOKWL57/pi23OVR/fqBEcCoY8quHwJCjFObTTAcCc6lCRkGhModEbb
EDiOz9NcP2+GRJWzlkxFF5tgZqHhnrYrtkdJW47WfZuSo8gcfsLXhvIHlhD/
5opVupbh8PqrV4jBcDDoPKOJt+ykYlLTGlCroFkbY/aZRkpJVlIzH+Ocjbpc
Lx5k0bWgKcJUjy2uo7JQj+QdDHJOzGDPcrjQaF+BTq7+BA5lg6TJ4MFL8a1M
cV2fo1Llk04jUz+La65H/4peuDDZmp679uxP2VjTkAp8d0+tEquDa/EcCxPi
ZxroLwdzX7CVucb01da3cITRQKj2DZSPeVsvB0J+v4i/4I0e+QJKdwK+SZP7
4WM7j6+/gLCBqo7g/vsW2q4icQ6w6+aCZ+NiYFpJqDObrCcg0Gu33ZtZhiTK
VT4CivKrWyP9ABNPGRnHTZmVN6sx5ga3Y+fTLb6wb8AzYTwOw1OG6TyEF7uo
cextDeLYnmpaHbyDPnGw8Y1j1VUfpd1NZOAb0yvB0uiVzzwNrfaPTdMtgPOi
kJsUZzMgsnBz3prBhfp6nMM0/NsohnQ+yVFL6TtkkS4st1ZWSaKG9gSKnpjm
BIiodg+TlZaVIdLGZyvSKUYmItFOqxCY6dEYMnyZs9FjaxzsiztdQxI3Hayz
crXuHA7tm8W1UlX/JmTC5Y4nlxODSLVb5jFD6ysgM6+5po/pxSd59nvwjEFf
x2ZGSCSVHHD3RA1jzvzdSv1Vc0lztpI49qoiVw0g2Q/XCQnoWNkl252AzGmI
h0sjShybrSKOTqfw73ydArCKE6M8O4yhRRmPHsDXB128Daj75I3CWUD+I0F+
9m0+IUwtee0D2uP2FiormWIV0VG6TG3MMh27ZOtXP62Bb+FYsLTx+dc01Er/
sNsDneOtP4ECbs9x/3klWkJkJsXWG6klw3E1wBv6skzxKJf17BKKP/VR5cNB
PDnHK4BH15LScxed4/5fbwOKy2HsediqHfQJZUDltjhnlH5SZlvc8C5P3/JY
tGPcBvULztyw3atAmh6crST+Y23LBhKLdEY6lGmrXohD+yrRUTa5nlOxRf3N
QfCqLzzXys38rlJ/hfg0tOOgHrb9li+YsKnTsrxZkShGqocVOkMaw9Af02YP
1cFctI/OgFC5CpuD+xzmxNDID3aZGMA4reaRAY6w5r+rLVE0Vsgis93oZPLG
r9nTsve1Q79a21wheVh+prU6wsyn3Ji1pShysom9KWvB6fOWerNOIARqvGrG
t9i7ND42EEMWuGMc4uYQDnR55lIyKcBC7p71+rFL87+Y0Hy/7732KqHTB0YY
aSedUiIpq8RnuECmV06Cnoc7HtbG8/q9HfbamzjDzDbKvgQMGtUot/K11Pd8
eZahme1w4icFLbb7HYcFNtsoGfplEcJ2GxmXtMt1MXs6ENq+3MDRa++WjdgS
DcRnQvTKs2sey5fkmBfYlpUit/Ehmv1m+ZctUYPOCWQLhSeGAItHKV+L3BFU
qFB5K+RzcXavGimhIoUIT+0LrqKN+Y0R/8vneJyhj5rgh7zsu8yBW6Fbn8yn
cvh+TC0PHm+uMvSqkdJZK5cSitIfrfMp2y9SU4qJN3DlahdzryXbrwbxQ5OG
PF/Hqbn0VVWiKeNPm+sJMAyALuuIEbsAIBat1eqF5HJP7dW0wH9C+un9LoAO
Qqq4F5AJDUD55VySXrYDLF8PsgXha77d+MrQ4/jsOj8nem/WwDDI1uDX6hob
05uNd+WAYQNu/YCPKvmDeoUd0CJ6iOxYtPT/Za0dxBL1O4/LGrS0lCAyDYlU
gSryrucWYfMldb1QNLj5BJ0NbhdeB2FBpBrjndGDX1GTW4MWtUpscQQWVouy
XPqqkj4l+fGxleUYgUpplBU7C1AUx10tBLpvi/OPHJhiQUXbfaAixFKWvH9y
ar+VGZ06ALoHdt4zFB0JPt2PA2fqjiHu1x9nkuGWlkL5xWeQyoapt30yRTrj
vFbJxlpYXThOwlFC4h1KV3ASvB87MUHbDXcR/8mojW0REBrF9HYd4gQ6ycQ+
thMrX+L/b3gXUdKlhFtPYhJv9YHVniOq6KQMzqsqen3Ppj12jh0luDApXK/G
+lyH+GeL0EBfN3svWGKDjki090RD3u9Px6h1cqMJvwz8YeANdyAe0fJRFgUJ
rQKz7liWLOC3uO7Ty7Ue5szHigNA2fHOADaY2ob+UVjIikyO/7gWrAlvevp0
K7wwo38iD+6A6YBKAaKuYUzwtUDn47J0qwaswVeZlWgFRVNdXUESjq1itw17
Is11mhKGP7CBXeYRM+eTZu5UyFU2h1Iu4LqSzgLgPAAg1UypuhbDFHxR/95i
/NU6PY6jrj+rOWxyrpRbIDbWHt6IME6GphtTVPhiF6X/xGbpk/juhOhj2CkM
RuWhQfB1zgYJ/kUpPxKfbqi2TGYlGvwjQPGc0AkyeznNfBA98+eSu63VAInn
e6r9yEMbrIGwosCVx4RALjv30+6SGftcCyPa3voy0Db34lYTqg+kKn7uEvXQ
ngCdfnKjk/FENKwWKu1fJAUEO8EW5PeYHZfpZKZmMPx2zG2F38QII8X7ZY6v
9AEU/s6xoaP6RFJ5QUTrTUEMGDiKQJIIcBO+pUZ8tUQyD2rXyh+XqzTL5ag1
z31NyZ7FkZkINezzq/jWqlNSdmU+jxVl602ishMjQqAei0mov945cTjL6dJ2
EYij0EGFd3Zs3aA2a7o6PK34muSNXPlyxyxOVtEVGCJypnXj+WBM9sLDGfav
veVaF9EJPiduye5hLWQXYA2NZhItM2PQh6NOSaPx0pqxr+xdFj6OAX8uv6wv
N2NLevZqlaFYUIfhgauScrzqh44CAztaR4Cg9ydLxyGgvn/l4KtC/VBrwkve
aIspdi72moJ7HenTXAIHg8ksNFF5aEUKxaPt7PpdVVdlEcFkv/ox5fXjSwIL
lZFAIQTLj7YYgQ68VA9TNksBKzeAQ6piHf5J6pMz9l+jNtRzOvWlf8HHkerX
oApZ7p4CvVzyb91BXAaHhNH/uorwCKO3oHNPN4vw+JWbl1e7Jeqls3vPXAzq
kGgDbNV4TnaF63NK02ydx/1rKm+/Q3DuvsWYVmPmTpwvr7WCkamVq2RBggRu
R5eA87z/z/VzOaZVvX32zpM8L6Z5gB/tHU0Y/UXGWCQCGHgQY6bA7X2k4on3
dp1n5VqI0MCWp9fo8ijGHSnJKqUcwqkBMZ7Gg/e/oV4kD7YaKVZr7529V4gE
9FbJ+yoNRkUmmLrIgMWa3woa0oOmLs3NlD77Qw4mxwoBsfZSZIdHD9e7OW5l
nhH/p+j7oAedNqAbn4Wc/QmwqnLN/rB9osBnj+4HY54jv3CCfq7EK0rRqOvs
hjN04nX+fv0AkJ5Z9ecsth2SeunOnHuFJnFjU6C5oiKxLFFxdEW4BOl2Nx0k
4uCwlPp22IDDgXTeBkMVYF/lkOZtTcWtdCGqsT1qOkdldYzLkW675WTuLAwI
iV+GVP+pt0IObAUIH6jAs/m647MgjmnbYHSdT7HSE5O0VIobhc4PdiiMCGlE
NbdGn7zhYkU7W3WlSDG9OW+zbZfogolgRLxZlXnE1WnN5APJY/Grl2weEAat
ClmMOy6N/ZutsoLCLKvxmcfjaFuff9MWPuE4EWb0mS+W4IeVesh5fQuzKp6W
BUmFYxknkYC/zcH1ztnlS/I3tP2sOgKiSI36OiNAZhS2ZnUJpl58qcdxk+m8
/TEXZYf8vs6S4KGY58TEV3e9YolxcbsgUqOPADdpeXeqXJ6GHWMHgH9KghZa
Jw08Q3/MXrgV2YOag0HAKg/P/qWh0gu4stAPg+0v6HrK2m82Hnncf48Y+Pxn
FWMlgOpYJyOXIVoahdio2oMpW2CT6sAdYHq0aRdLZgNuXr9XhKKtcZHxDDnW
amkdRnyJvnuQwxy3seof5HCbP6WswSMXrDaF9Abonw1032YY4U3dO2nPaHvC
f/d8yZJkOmwPeFr5UR2fkbDPSeqP3kgQiSL1cjF+sGWXdfxIf8l9S9D4FVJH
lrOHT33haxPozhJ0yGaSkIe2paiTroXa0txATf/z6SBNpkK9p3KT/RES4TJ0
Da11KnknztZMZqscmZwrT9DtLwnpd1RDzs4V37Mgssd7bFl7KD3NasuO9+QV
5JWAkGbicO2AJmqSy1nhAcqoxN587vyqjp80eAx2vXpv5kRNhUkBf/qNB+/O
fnTl4sYo618Nqj5NRRKvLvPZpldO2cmGc2d9TNv5dJj782e6oaXSou9PLjrE
ZJ5O2kzY70LBlFPjLO5M7FGecaH8xdmRuDrposJuw7JTf8emm0LUa1gHLf+a
dDW8pfUc44RXdKsoIWgTGHrH5B/0ISJJpiwJv1oNhqHjDHqxd4Izq1+f89Z0
dSAkzlT80I5ULhriPCcVqUEr+wbixf+ilVRiWOY0JTcKnSgi/d3zKLlZxG0+
4uuhdXZ5PaPPMElIjo4mZmlHyB4vIu5lkiW9uTnjD6CyYjqHu5LAt/0sN/NU
hwkw0lo0/mT1gJNQAqWQoRtYTRP8fx1h3wrut/HNpuvn+49jWL1uoj5TldAF
//IXIUS8SV9AeQ+uxhy08dq4OZe1BaULg7afLLI17gXicc43Sre0t/EMjcjE
TRdDSj4nkF6JKI4JMiip2vUMoZ2IFGV5EYY7SpH33EdeTeVtmRb/dU9DbBtJ
OYV7OrtKQqfEt1ZxIhcZMLYe/c7D1P5E6H96We6w4tiS//2Xvb/PJ6lnauCl
SI5NcriXMlYFhF8Mzk39gLoT9M0gBgsqCUuAbjXU2VdJAuJgs7ILAZtJfdhM
YyKQhJpx5ev+lCCjuW/kVbfXqjZxNUaxhEHOPVuzkdEOuOZekVz8e391fcDq
77Hu4IPJLlo8KGM2QN+tCfs/O5+KCVz//aFUdVnxfJ9A5kWYA2UU3JzEMWjh
5LvKs/Gtg7jjoBT1w/KefptcLiesZeQtHHalnswgf6AhAqZDo6Op3ucmVrVt
TJcuyJ3dDXC6A+IJ444XFqPn66IXq1Kc4yzXjZmxo0jahAUB+oLvp4bMfgYl
DDvs43g0h1AHxIPERdHBzxwzuLIlxNzYod/pJ0biqsJUkerh3piQxONMl400
+q8PY0qh/zsB86dUoliXzebf7bm9ouSnRcUqu1Cb+gOdVsJbyug9Qk/wb/PW
hf8eSnuW5RJBRUq/VkDTcoVm0o9towI7g11V+8FOdydEScN4OXuQQfU/tRQi
7cBckGwP//03qruz+f8rsNzmCY+9KSuJZJk0iM03SxwaUpSn1OhPkbD8op3L
Md9Ku2DvqwN6qwwkhedNpsa8tBCHiOhsAjtnhef8IClIE55fmIR1Q4dLMm+B
jsynhI6Aav9VqdiQ1IfwMl0lNaGJyYigl8WatzQkr5b+jttViKgaiD7jxaDP
CPwF9+iHJQLVxcgxy3SBEDn8RrqfVvB+ME9kq8yMoPTtYCMRRhJbo84rMLmy
wuDekWtQiBL2L7ODcNh/6JEuKuqxLOCocM0eeg2OawqaCsnmaTul/xBJ4CJR
W0X433dnUmBYTsbZPUPTrv5fJRk6NuKbTX7NprToLVGDCE2lHnKSI4G/LvwD
jSkrSjCiS6L2jsAmzdLyZ0fTRLZY9XJbPv17UJUbIuELeYyqfD8bJ2pRyMSN
IcCQFGaR1o6yFGM/8ZITO4nO58VwQbLjuAZ3Q5vwu78hLf/GPzt3Nva95mP6
pGzPQeS6tJDPU0qlu0dUTkbvO39sJtDpLfjlGus2rDlsTadM+JYsl+JOC/S5
sXL5CR0NAKNASiqE8LJXHymnJ+7aS+LTAQVfhFlLDA9p2zL2wsWD8GtWQFmD
cE+w817xryhyU7LjttPOLX3WxOoYyiu6hS2LNo5wbcP+LGZVcsa7qER1Rq6X
8rUWfQlZiSyPhZEUIruNvfTFY+XSLp+DSwBujosRpaSWFWlEgBBepuBKrbhM
cGWMlCKop8IswFn21mf4Bqa2jpmKY15qiksKEk08Dbwo8jO50ZrXkL38S5ql
jiklcnbMcUXr1cwIfOItvS1VmNqmfhvYcNEhw9u7QY1/Q/5keSaDOOXihj2j
cXZDqM7qGjlCptB3koZ5OvphxnSzHvp8xIM2hrT2fZgQUzz1pYeskzmLMaDo
NQBM778FYu5RiLACDYMkhigwZAkEadYI+zEiEFFihBVhNeM2NBQOAROCpnDN
NITkKeFF+x8dDsW+BDmMysBi3wGWGZKO8MYXvGXa51gaqEywIFUxnP7/elB1
4zhH+O+RiJneP+EXvH+ItiwfxFGYKbO9I2odHTq5RkVgT+XPNEv/3TqDiUNh
HhY6RvVEV1t3jYB7EQA+iyJgUm2QdxTu409ua7fJ0tblnhThYzyJGkx4Fxgf
4d8QsfI3kTNkDWT7jaCH1QZeXanEtOuzomAnTt2mSZChELugM5oCmyWLOdsK
kZv3i6nWiKslR6kxU4VNyOmziN8O+5QMrcFnqYjdvN54ZWc0rHSbAUg3SyOb
pEdAl+0pCh5ZMUF+9s5C4HQF/SPEwVjar/6+ISCyoW63NsNFtdp9XcPj6Mtr
rmjKBIfu2Aho4U3ofDea7lN20oMbo4AnnK0Udz223fLT6AjXt4RS6TLzyfft
uBIUYGaRgOmSwfe1uUrg8/GUtIjdTpHDrKDtrTsEkCl8M4V+3kpS+/hfzRSf
9qKuwXKi3zODtDG69s3lZru+J695m60aLiHXuAVAAk29vOXcqEvXPA5+Oi4X
ZpjxkCO2eGYXY2DzoJJCPwRRRB2UbWvWkgFHlCUDYpdnYkZhZvsv4S6ENDqX
uoNEPR4QmlNDknDVuuAFp0eJFCrdj4Ic3CFzSd7+2F3niIjXEnuFdMpsBSkM
KkcX34AhcJeGWq376rY5YVOoYU3PwqEDsrHLuiANjHdIlNuSVYCr4g8VUsbJ
uVqqO3uhItMy8uC5zdtohv8tDBljwYPxnWHcIASk2aj9QgKQc0RjMkOUr8T+
1STkNBCwJeBmysgyip8zbaaev7l7feF2SC2gux6Wv7McIIG0oI7XIHEHn18m
UesSXSE4q8S4D2ovYq/Y6VaVKiHWTYHGAgupGSG2lM0H6uw4ZnEerJ3lTfxH
4RSvbKADH5CtcXRZuW+heehP2Pogp+b2ea4f+m1ofPSetuIYLqhylBze1xxy
M83iyhfJeMTgCH+lJRvgoSDUEpwWuWB69hr9MnAYD410u6Yl0r8SrL6fYkdL
Ua2/7g7e8K50IDHdB5yBbpuT+NUwtdr1QjvWSaDPEVY/vtQzBOW2TOfgOPS5
PtV/dst9D/uw5qCKhROZaxMZrXzbMlMSRWz1ELulxec+PjVNwJ0V06wngSKf
KkI1YJEK9PrO09EbOrfJUZHwVPgZiSxav0K1vT4PsaUsZnoFbldDenCm0gYH
FLXDa5D7GFhoBGAGefL/7Ddid2kNuDyl9vwKks8+9U1XVCZuqgyiWRlSbepf
72Wg9lz3k2Vu1UhXCOhp93YE9DE0+ojAWV0//PlgPRJ+8sMcR9BNG61v2+hD
HHqrpF+PsGGLqOyNiFvQuO/xU0VhpBNzN8TX3bnoERQxVLGZnCMjhIIDWoGu
iWOZLTnX2onlUJnL97PH/BxydZ7cbHWHy4aYUXmvfUeCljXFXJbhXNTthHnK
3JyRoTLzsETg7rDEqmJOF+dx7HaSN4EvBX3aKZZzvjsdLXSVy/WRBwg0YStQ
vY1dt6TTxmP/iBpkDfUaUjC8erNzAJFNN6yPMdzYv2i+3f0FyLB7aQGg4tnQ
Qluv81I3VJ0G4imN1gqam5u8e7jYQ8vMIppS+4ci6NN+IhZhsiLIbLtuXPfT
7k1y5BdpNZusKEJMwIrKSDwe5id8Tx3hgPvKohAerXoOHMpPc7FtVb0ubcGH
M620UjitkkW3p2ucV1bx0JgOKo/i/k3Qmu9ECvJGxV9YjJN6UOOXANK4sgn5
oh1ED8RvuSq0IGS6qKj2wYB4765yCNr+1Zu4zqzlSL4tP52jPNm88IshhwG+
GsK+wkDQ7wMp3NaQclGNlKZ7zPVwGuswJNR1vgMBTuTohKjnFeQ30S+XkdEY
ddpfrFmaK+1vvypEP2CO/1C98Bp6gZ2iszTiPTaFk0N5FQ8otaSGoe4HfUp+
Ab3WHVQXY+XJGdLwLfwSu65OBy3/lXZR+0BSa2KDJNfXkdAZp+kojCLfGq/C
EKSpe51Awe64SZXUm37WRJFaEfmpxhZEn/eeQOtlpE7+a+MWsRzULGjUQX8X
8p+llm6Qm15F4gxwAbzOZdoILA6t8zBLWX4Vazsu3UyOvSTANfwaZQ0ZyUcM
uXJhIBhiyNjtefw4Q5fv2f2XQD7bwBPZIBnkgGPRRoxaFPZPiRg9Ypic5zOJ
7nmCXiGizTwrNNMYkjO1ZV2OrLRD3eByStKuNEifterqhnd9iDpnxojJs4On
VUA+cnBQuQrgbIsCcoGLCgvETF6WJf5Kt3vn0yNz8xRFHFCPb4AggBQdLCPJ
SxW1BwL79bUW5JGXATDO5oZ0BilsTvaZxFzQNc6+RAjXO3xfeP6NgeKLe74X
BoF5vPVeW4lofXPJMu7HbjaMquzhPIFMZOk7hF17Ecl2wqvs9rKF2KHM43S3
duhfyeqXGG8rIgv+S7tfTjtkSYJTr+JiQ/cMLthOFkclqlRxxHITV6lhrOPS
MJAz+XGFfpavi1ToGO++mJdPHQpOvlV6mtgyFpQmKULcRGFApFmKAN2QGnfQ
cleT73G/c6anZhJbY6qED4DSVRLaxrsHXQTLCANtRUfD/PMyLqJaMyChc+P9
MRkWQ+MsaJPtg4+qhRFjs9EK0QzOEDUVVc23aED9FtVAcrg/GrONKgNIjJxR
7MQNiezHPsOTm67YnXIkjZC1XAQIOGjU4Wt9eC+Zj/j14041TfTPEaL69z54
ZbcaM4e4FMM6d/d87NwTGcLMIJh+PgmCkJrL6DuaVYSsy69VHmxfYjA7lHPX
1kU6hFcjpGlCqwBWg6/jjPCmMSkC9/n8QBVdpM0a/s4E/8ugkJrZRC8CzmK0
bCvuY+fFa5fVqbAcXfL+Z+jOhO+xIWNhdIuiVUsBZD/55nLCRJVmUAtATHCP
x/57Bqiqj+Tn8SjYQdmL70K7fQY4618tbSQ8o7JBE/gDUO+VZLrXcwp6YACG
PZl4i7jZNVKvhzeZTMNiIrP8I00cGcrzzp5ZBdN5RjMYGvg7vX7w4aLjyVGU
KR+UsfAIpmBs3YhmEYZKIxqJLzLn4ubGw7OZyPdet763MkAmxZTlCK4Pzi5L
3svyDan1Ipq6zIo3hIrFL9Sm2yf51RGUjFnCNgGu5BE5QEkGMyh6cE4VyQ9s
+cFUbSi9K05LkoA08LLkF0Jyog7lWXopBkXYptfKgfMz+Pw77wAyZGyqdE28
TejhtsnHQb6IxrrvVMPG5iqjC7pzKch9i7YE8hkmXITUywUOyL3l81x36zpj
WWz0xpQNjH8P+E6Yxh4jFkJHY8zgltCR3IXTo51qHES1Nm7WSqPVMvTa2WbD
RpymcY7CxpijvZnnFDwLkFGc/5J+kezPwBh1phs20sSRf0+gXD39Hhxckfwu
uXaS2a9xXwqlEqd+DKIWu6lrcdVuy3pl62CN3kLhInTfO8kX3X5JQ8zXneKX
uYDiuLmXEuVsSe83VJWLoveU1/ImpOvhS1WEH2kO3/f6x6A9kQxA4CxRZaBy
fbvYmN/Sid7zkZLamymdK2hOId72gURtyLbuhQqNRfQzSXhpngpX/jvZ0wlo
vnl6bUHcE5Fuoat+kDKbQBGRtMVMS8bGnOt3whn85cm8CQsYdY3BEKrp8YOQ
C5J5VlNm6cnmpNAOcPd1Y8jRPIC69S3A/FzvH8XDpIJoCsRgCe5uBW2wqgQs
5Yb36OvuINVox8gQbWkGozVx//SGAJ1hWo3zoecdkLU8bj8ms3HXFBhfVrx8
1lkEnyjKchwGWeFOw9Q42R59g9VZurKx4Ipo8cwzEBALhBfBN3Mpulef9Tmi
5lhceHPNzAKBxGSgANnj1ZfZQc4iBHv2opy5W8DZF5AJrDF6+LABXqVjX8vY
oiMyq6E0ZBpMKVmAPPEL1NlA0KgvGO2WfVWgcRemG/HImAIpfKf/95xptvMC
JBKLD1pYUi+efXOOU1jtBSfer5xskWSm/mRuMkfPj4VlQRAorZhiB3Dd8eUQ
xuLetbj4Asmn2RnxJpAeEJfPlyNIix4w4et9RqRRCwaT2oR3BiTelLOKm2b/
FW1QhVliXne0AzYaiXx+WuzeEDwYeod83z/YsiJ5N1U8U79zXen0fuTOoSVf
S9735Mz1Wb6atkmAWgvfpUtqkCWOVI6OxmqmUCupW0lYObesu1m+1vynFiFX
iV0vtrNDOPyqzbmO9EeOOxYXNg0UnpcP5vsRysVKI9rwUB7uFFzb7wpC7PH6
E8g/YYPvlnQEup8WG8g0kZlA84gphxM5rpBQlysMt+T0ydVqDFyVXNSeHoiK
Wpd8L3X3HHGxvagP/QnDSeTqalFJxki3u54FdQkAp/P72ySKfIzYzAfsxOX4
VhKK1AUQuogXddiqeyKKDn+k9vvVXw8u+bEyDV69+qoNn6rm/bpwfBO5NJmJ
/M0qXqqRLe9ln1EM98VGOzMLXn443hk6GZBx4gWivblWWd0y4I6WETB8WIcr
MfuvAiTehTtBx3l5lz7v6Gge+SuIYpp5c+12diyY6R5l3YNm9MxljXMvWjfo
mo0uf+aWBpLIdDbwwd0rE7uIMFciPnBD3fYfc4V1GOmfpRfNv/NqUQTZlwbH
tAzWjI8Z2lvnLWxcvSRn3SSsrkmOYVyfIuvm3y5c46WgxqXcM14+wEslK0Rl
nPI+q65Pd94I0fSe4EcGULWw3V0TKw0NnKtqE9K/VhBVzqTSkVDp1mrpoNVk
48fAu2+nYoGg39r+eolns/uBq+JJ2nwjHio1tFMxA5zyQTsmsB+gXNCPqp0U
ZXNECf9B6CfYK5uX/Ksh/DoDiizaP9p+48y6rBKQQI/40ZNma3Pw1HLCw/ts
AaxcymUZZyLgJHePdj9BimqNmpwZJKyA4Dn7Itf/I+AjqN18gmxxrzBcakZZ
oFfW+sm5GgCLToz/vrEocGHJtnKH5xpjHmyAq5NDJsAq7uAA3ySiAHLGir8K
GZElie8ZTzq+vFn+n9OUQoXINnVfSP+tM9jy8fZfuVCt9JzhlCn1WvdK/Nwi
p6Stkn/EJFVm9///XYQqqAhhwviNDCOFK5B/6pXnn1s1moAGB7NBeMIc8+bp
dho03yznY8Df2yx1HvTql3sFTh4C5DOi9hZtPHuZEOqxHs6r2mEKVXwAwoYY
B7Soz7npJN3qV9nWiMMIt10wkLX2HF76ZAAoxYn8XebV4GD+yCA7ZbVh4UYk
LJLNoXw5C/NOS6yduDsltF4ImCj7v4XJh05bNB+yhp9R9VrjkNqIhVaQpGeE
WMXmEb5ItpV5f9oED1F3O5uwlzN9SnswOPhMoEMKb1jt4nqSYiUXHV5rAUAg
p7YjgO7QMvzhCcmY1lDngcAmAsjs4RRz2/oElsVLXcVP5gWGXRAotpZDBzp6
4ncFb2i/6AooboGaJJ9+C1g/xHp6/iM+v79rR+W0BXHkQauFBm0iVXEOog2I
CbLTfZ9eYgcqxAD5JK8m0yWPYZ4szmNQ4izSLK0f+AVdv7kCODgIP7QzAd//
3/d875N59OpGt0xToddHIwrmAnOU9AhpRFB2kohR4vkfDED7jepGXa5Mgt04
z/mY/7NiD9ejdFLusj5rVA5g2743KinnEnsm6MgVb28/WaXfZ7JflY2o9dfw
vFbGiRub5TZkYrZW3JB7ocil9EMnVcA8t0cAl+bleO9pvUB6aehBY+pkzjHC
CArsH0+ngK7Pjd0unZfOcB97g6+KD5ufgczZpAP3gnFgIHZfUXMQbgVFULTL
/PtZCAaXFido6TU1rvfflhxplfvmxdUUuVXkwyobNWQuKICaqnYGWLOs7CYs
x0BDtkKBr8p6LoDcbfzYVwkZ52X5gDb8SzIwXjMdbNdazuv72OMPRLsnDBin
A8nszubHAvUBS5waaj+YxciXXHNoLkYBzxFTRCPGqVss7CPiAhuYqus0h/Uh
92ci5ed3bDBzpUb4jialuvi5Pbw82KcWKqwrdpYoL45UQ39ULiKgqeSOnLfU
tzELRiCZjWrb45n7VtkKTf9VvlX1vPfgSz8C+iK1afWUKMBB1roiH/Erq8Sz
LYKLbw/Ns2rEQ93Q0+5DZRBMbQfR6V5o9vHC87G9c4un4IW3XEq/BrBVp8kQ
JK0SNt8ftTK0JieIa0jHuHuwbcT2xeigPBU9aP3gF1jv/TINEuV4zMMIr36n
j5JL7IIYARLfpSDqFXEhTTCN1mRjjP7ie0WOHUCCuefnqquedqphJXB9+9A7
uq7jD9HP+keYK8wVRER81W1MZmblEoBhg2q7ZEJUPQlAX6XhAITPJ5UL4xrt
lnvGl5L/OCAzHkqfKWc0ksO8SoLKLovoV6b0xybsY4+gCRECAtxYaVuY+dTX
uiITWzqMtzOiD9/VZBFnLzBW15drBs8GUpflttJeaVMz7pI8eDCkbifuqaQb
sSAxlcOZfF7kaZ4eah2C4TfeT5+CArdzXnUDk84KcAc0I8PHXr8+6WIyLOoS
stzBYBxNwr75qcLsGdGRlkjEFu5s8eyCKGZxUy+5dPGYvYlwVu+zWfl8Ikb6
QSJv4iKl35+n1d8gU6WMIHhBqQyPm8fMge10CK9kKH7d5zdDgBwTb3+5RbKz
AY7EBR6WCVDFoxJNaoEpeTRJY+R+6Qx7Q7R1N9A4+HePdMdW97KcEHQLBHdd
NLT+4WEeRWEEjFGs0ezwaBYs/hS6MvUE1ZZvuKmnFLYVRDn8NSBwlgKTwZuT
gykss6KPT7j49vsjLJtNwwDbFx+oUH3/deLaI/1DMsrjw2jxQEwAQrvt3saX
tdl5AO8MkiBsyx8hL3rKMMY0H8MqUIFbR4DpmXjyI7WoiDpNAuPzOILX9w38
u1VOwVMUjPZHKIvTXg8sXKKBU3Y6FXgS2rDit6E+7h8qujw9pGm8czWBeI3d
iJeFUkbebOGP8EnePqU9kk0GjTlT7lKet77wMhg1yih8TyUbbxqQy33HPCdI
Fx34Nfjb6I4Xu8z/BAPqrnAJHKc3H1N8dFTwYgf1RXRoMLJV7sH2pPCN+Brl
qNa3bKuuJvxDGOc6KyvXXONn2jadLENBeM8ipHAZNC+b+mpgRwPN6EryTw/1
7Bpi50TkD4+ALGW/3OEczz6MFbDWUVfFUWg5RCifa5nBJ/0xAPBDLvRIOMUg
6iRXQsDa/DJNME05mpac8KhDPmACIFy0ogYkovHZuGYuWWZFtzoUckCx6xVC
/PpIRh4IdNihb/nbQeRf2xf0Fq7PADj3nHmbsRnGs4xpR4KrVONrhQbKq7lp
qyc363PBhjZVoxvy6b5gFDRx+aBdPuN13CizhZCx+VNVn0qjWLrd1dgbzS1R
/Bip3oKq3CWXKBNZ0eVhH5v5em2XizsFR2kmCcT+KY0m5obj+/8/9LdXcowM
tMir1DcCEEVXDfEKzsrYMwfysaGbkyVzyBaFh+wNCKPEkFSwYTidKoyt94So
2UMtv6Qm/WQ7kkpqUwOXrnhxBm0/E08o/W0fq6ULYcumWMVROe+AH2dZgddQ
GJnn3OdKlRhEzhTXScRC4hPWy6TVKTWuRnfJPHpnTXSvcyQ4wTT1u2L+m8W7
DAh60XEohz37/+YaKVm3JNDp5l0zWn0/tLyY5oSy3Jf8QegfpoP2bwt3Zkoa
bRzzEWCkcEs4l3XsYZhgjdspvgaoT+7CaaLyD7vWiWXo5fSrWX0rVppRsAOG
AjZYXKona14g/0t5dCbx8f59U8NiS+XOhehXjDecLBj1gef/QXirJgdomRTI
5EgYii9b6sImjK5SPzml/9jRWxOQqkxXf9rrYo+5I2ozgmbNkXoHSD7E8Dcu
y1WZiZZqHkP3hu0OBDbnU05eOfG0w8wd6Cv9HaXiHgfA0YaVY8Pso/TWBEe6
C6itMUR0jdvpSjpRlxA7OthGZi2CtJOkLKxtu1PLtPHPFUToi6kCw6oj16pr
tASmSxG71+e9On9gBN0gsaDVBA1LCfQv+VCz7NLSslg4CgTKTb4PfCEHR6fK
mO5TY+9kZxjT2j7mDA8x0kwfQ9I75i/8YjZYk6Voa1Uglfei9zrtNLXV7EtR
doJgNQ07BwNNzXPOK46AQIIYE1HoILOr3XjuLGUAYyAzUtszj/vAFihZDuGD
4IkfK/flNoM+CVEfCtmaH9YDIS1ZAiGbUPunVpuit/l2lPGUJQotXLWOvgDh
Uz+BmnIe3M1OqfQroBZuHBqZFpwbS/Ez06bA/eUYLY42CNKLmyBW5JJ8Ms2D
2wAWSKCD54GdV7HPARsWI0dyLi3qTqWUaaQtd+LT9JuU1EIBNn6sCkM1ea+G
LuuMkVAhhR642zF90Vk/f8JDqoL7m8gA02t9Huik5kBal7MqH22nJZUFmJDE
6nxGmM6MvipbzfTYvH5LzhkAi4KzdfPhXvAWBo/uw1dyrNBdv6/6RWbQzdJt
7Da/Zm4i6XIq5wKrEN6xbYz+THDlPfklnPluoKUfAYYi4IqVE/pQX8E/oKkb
SX65QFh/kYk6lBBVN2Poe2M9U2rhbn1/tEpHAggHPJYtDytX6N5qMAn2L5fK
TjZlDCF3u+KCg8gPEAMpICWD8emZ9/1H8NNDcyTIx2KlYQoVwQcv3HMtoeuJ
IEo/ziMUtXlpfiggNM9hy/Q6tQikvPR8UxcRQy+tpBrS7K7lHVAqnSt1cUCR
LOH0UXGhwzBeNQLUzdghYzHy19PSEhEx6GEVfVCD3qUvfkVjNaTpVjycMNdq
5vH/FSe9tA19jIlgHPXOgflpMj3JrqNe3m5dHUDP8QBh/hx2TUace4mLHFch
Hmbypf2I1O4gL4fauCuLXRI5bZxMYrcItMNRLw9MLQD5DVu/IvTb2KneSk7n
npvSw4gbrvX7Pl/S45/pm7oGmY+nsK13UV2DYdMeD9t7nsOLwEqwjn8GAAIr
ljQ8qqjXFjOefx1xRRzY86yN3Di6Q5bqIdacb2ETUn79nEd+cwWK4jVVqQ/H
KZoMpgBeHfOCBNAwJGiscpMUE+2v3tAG7XcAzAGAo+7+whyO0oswwN1Bmlfn
sLbsblqUX5vbJ0SKVnL+Ndn8ialKj1dKlJM9KTASskrmR/rtIGKm12p1OmMY
o3yJ/vy3NVu6zrneAXQb2L1Tn1o5EcjO36pgniVEEzUmkEtiaMehBMdHbmPM
QUu0N5LY/bKucI7R/IhXtP5a/Sv70RNp7LeYCpCAZmUQxyDj4fPg+1GtVqqv
+pu0RZ2N5RHkF2XAdBIE1qQWeWH2cdOyVGkygEXpXED5FIfSMn7U/H3XHR1R
ckiswjk/YUdlB/yo0JDt/IrA8Mg/ZejpXPutY2b6jDjLOTSUG3eVs7bUYSPy
QGnk+TG1m3Z/t5+cKgJrfvuyUiW/4W6YxEJmbURUPhlkKWoHKbFzCeufYGVq
x0DQtQuMb7ZA/aoAvaDbVBVuudwPvpq00dRcy+9hvJvJpV/a8PaU9HmsOJM1
1UnZfdx2uAtnzilfD9eF4Sg2yB3xbKNKj0MngyjWP22uJVy5TWWgB0E7JMfY
XyFRmGk6AAelSTsEHAMLKC2byzki6PWwdXgLUmRcHkSE0nuAzRRacPhv1Rzg
bdi+mROlMi12ojEXhUOIK2QyeNjszeXVj8vmqQHlsJY0c98QHH7qThnLyIfS
JSLsPgGoYkOU+X3czAWSEDod6ttJB7ocghXubh/EDMhgUNVBxRemvAH8H7W6
/lSpjfNLXt//UnAnfrag3qVIGvrBkiOR6pNpgJurKRzl4ZysE+b/cElAAi3F
oeuz9H4EcHNoy4oX0fg8UNEo4TeJL+Nfvrs6H1toflQkBrn4XGs0P1TrW/mm
Aeb7FoEe4pSVc2wblNUJFyfmaE2fxVDJIsVMNBBfo79XhdqUGKDFldy2k3pw
eSpjd9jDH011+V5u5jJvROUflWLrhCXBzv/PPL/ku4cY7mKOtQM58V5KYI8l
lk9ObII2o35yEEurQreRxCZkLFYKx9W7oWcMynNLdO966yCeNk6LNWGyuLhT
FFpe0gygWGlBe1kyqaMga/hypJhPNqG02Y+1lbeX60t0udq2C7cxOct92i9E
aqCZ6WRTIW2g8rHK7/Qf9aoxLsUbKgQ37lgSXvWfhFfN2ppp/us9Im6yZbtd
t67gzeC1IVWeIojJ0UsviFfb5qw/5VO7KVFzWi1HiASnwwZywU1YdnhEP6Oc
4y5RNPwKaM2ORbD5tipaXqGrgmi34CH3G4DwD3WBlL+2rAvn9zuKeBuBohcz
ubVj6ep/zRIlgNVZnNga7xfY4cF5zFT1EDlujPxGFrR5E8fNkcbBUsrpe5Ke
bdKDjLtdUtuCYm1P2P7t+Zqr+Kj8F6HIj4jD1CCUD0dYXDAsepGXHRzH7Tm3
fEc1UggRk7EpN7ndMDOg4oI7oIrsQAeM/qbAwtLqRdwkFGcw5Vobev3klbUj
X6XfAR+pbi4Tu5G4Yv2FtV+3B5QyLEfCVTYHxLH0DOb1TA3kvK8UOkLmJr/2
XccDmVPhhmWR6tWMW2X/y1inmEyt3eodF7sQZI+K1rG+voRmkBWbd6pToU/g
osLYDHLG23kRjFLPazkN+529yWcq5vfLiIufXa4SCCMiIuLFN6LWauf5iyEk
RmTyqg5wsZJn2S3FRdaC7ElFqHDDhsecYdcUCAu3pJu4M+9I5qT/pqW6ZVgZ
GQ9wgKhJA5mdDJhrsjme76FmZ2esCrJBUY2Je+vig7Cvhlgc1IOhuGJ4daJ/
8NBAKd/fOMDP7mawtIjiUmfTMKSB9qzCDMAjXJMWnDJAUrepTH3C9lFN6dBB
xEn9VIYfj4R2/CkwAy5YWVFVEQVcNOWMHvUTNs5RkBGync5G0Bk5BU1XBdV9
K814GOHVgWQNtwRtUQ/CgmTy26cC+xsOP81k4qc12x/6MU5VuzylmnmcNMAz
raK1FHnydwAhbXJZXimih1s7TAu9AZulU4ZQFA/0tlzCJwG9Gg11o4XpNVKm
YqbTv512DUIFdSp7of4oLSYseiZOiKPtyIQu5LqMpnEqYE8QpP6V1C2CZWbl
iH6gvgmZPcJinKjkd2H7HIi+xvon+zG2G3zEmcc4cy3tca3q5TGyzth1S5SP
czo3bjoXXrb806fIslv4svIYnerYJMujzYhSHdfHGC57Q0pLb7JuvS+ZHcqq
X7AKrDMyi8HR6v03U3Fv2xMx2D115zVDa13uqHZfu5Eq1pYHbvXFgh2Y4U4T
jyejBrAMcDI/BmKi3IXg2kLmrwDqIXyHEIQnZIJaxEufs/VnZm1W3/UwvFQl
OPkZ2YqDnUiSBtV/E7nn+Y/XW7CuoT8aQ9Z7FiXydl57Yie9vZkN8WqdLl8J
7AYAb6QLsnES8/n5F9CVWApwUh3trxkZXOjvbKIx5GgJIA465eEF25r15t/K
TLTsg9D6iI4Sn6KSyY0ChHnBUeqCzMTgWrnOCcOo5lRd+DsOqg41GmRgnd9b
QibX/hYdYpH4HH2dkQFjxmjHeA1ZVCG55Wlmzr0mfDdBYNKsgswePFDyxT4k
2ybB2qKAbbiDxSfDM+LFlo2iirE8KgdhKEcILkYtm5k28GyrMroO41BVMJBh
ZwrrpWZJR6RBoHcCzUEZoOTWcQGWzfly9Fr/HUof+1fjDY+5Q6wQoekPPY2b
XOSOnoCVxrEq8Vh/Rd6i5d3igPoYy1yPpuPm4FsWQMkuCMmoE0YdnokSjwd0
bWLXZDftgegf2HBX2hYSrzZMQoIcR1zFw5fTfMh1unWZpFCPji+fu6HLa0dN
S5SsW+OjhKS5mfqYBwFjrGI5OccobKmJ8nltVL7MC3gnA0RljeICcTrrFQHD
0tFv1ka/I/UhKLtnVftyIfMXDwo0YLiNUzBO69lNZ33KSUdAJOkTLvl8lZgX
sXYSOFCLBjtJ8ZLZ8RRk77FUERXLWcqat+uaIslVJW3Otv/PPdevxML5HsPG
zbhG38mX+IQIR+z4FzSa6RmZOMUplWWi9nmYw54uzF/xipQbSKSNnlkDu1gp
TfK6F9DyV8hQMt6KeaVO4XHIwg7nPhxIcJKYqApTl3+XFTMBsArXHgdJLQFH
n5G6AqS92oYvBqaTLv2qRO4QFSeXxAMlhWaUshHTW/Lyp4j4RSfUI3Rgks/S
uHm7ndVWKcpt/UoO5DixPlOtHnFet6wK8Dcj5uPJbU9/zh+UXtaV2vyEpooV
zlDwNF3CGEQdFv7QPkyLCB9dC9o8avLyZ2OaM3QPUCiCDhqxqkKRZYgqgWZ3
gujdubMiK2OxtjrYvNmdwOcYplemOJTKvRq9ofQ3v9nLO6+6faqdHyjqsZri
v2ygW/VcEejNpUia9V01c7guluVxiEXJ6jWUCI7oRyxZNMHkPO7cN0Rc7kxd
E9DobpQDFO+PQvdQv98yRVvFh0w97J8GrY1d4Wl+6Gz6H1+Lli6ZSRliDMIA
uyjXO/6McxQyCkQFpFg0k7m2A1l4RmqJpXwXPb85BVQhpzP15vw+2UFNPHBy
tI5RgCNDnkJNtniM3d6iJPzTeml9OMopLw+aPGw6+D6l7OqJt5BuZoUHQTdY
Mf/NHbfBU/z4E88MXrFrEIvqbNtckgegp9Qv0jbydrY1Fx3HvJhWevzo8sAW
4KxTthI4N0agmPa/iYjahngROuy4rpXtyB5b0SPClGzyWJbnFUeMlV1+1LW5
EvLlkVMdP03BgGDcrdvPBnPpXsL1T/CMA9YewnSKH9D5keLO67//hD2GHSY9
OyxC/PBLgb+O89AX8NAcc5wnL9MJ7Ro6Y4qz95/IHI5c+FT+wBix2wEi2hrx
XVQ7u38uG9hnaW9u00VW1EpNpz8vfa/99lgLkwFz4h7OYM4FeXGV0l1znpb0
YAOd0p7WOWzROECMJLTdjGBghM37k5oDvEWqFTlJzWXQwKb4m49uVkD1b9gO
VYay5zLc244v8TAe1Ea8Oo4D3j2KyUbX/QM0C1XYAitwNWIg5fUZWrFl6yNK
YYxLFghjcSSTXj2Qd3kSMQR3Qz41eZAdpyjj9Zmf42tE0fWO3uR9q0/R8RtX
tKtj/vTp8TT2XeoXitZpgjp8gvOA6f9clu4YghTbR4YcAlEj3i5UGMKPMUmk
GEWs9rQ4EFHIMUHEwki/hEQoDVMtP5K+yaujv2hGLy+694V9euT90p9HWoG2
rR8+NuvzTy9RWRHnNqRen/CxrbPnsa7dnIdYCtoad7qBl4Zy+Jf+mFM81k/P
q5ivUXuunSNqXUz/XJJ+KeTjOA33p9b7IgP2z9vjzJ9NdZlNRvc6TU1hcAva
Q8oN7MHS+yinzRJzoNR4mA9bHqB1W8RJXPdPu4OUXn/2ag6u4/h+vR4pbIhK
hR4AmyZTX58exvSEwoEXHvWe4K5hgKYBdg0UjP47boo5o9gCqVp5AwPwXA+q
ATpvsKR/h/3dDetcyHnaSxZ2Qsuhp+s7PsjbawHcgJYFdLXq7p00k13gzE+P
1u/xqa+SbRtz9f8HHWe7qArgm2KQgkD2wvfSBUzklVurcGvEhGqbXPya0EzB
Lsi3eW1E70KMTlKuPlunTaxg0zwLSieifIfMwWbc5ulLogsJKha+q3dbr6zB
SthZ3JqB9DY3mAtunw8hED2eUSDa0MSsHppE0S4aq2wuBUvLTa0YIfXNEg2f
K+75BVAJdGM/sFATGVGTyb7yt5HY9Q14QOwqqEAOVw0ROqttUfcZHj8QQruv
6YdwpGmNLvJsnUdz+3gM2h5cX6Gu6tlaJb/NfXwO1QjEffsP+rMXrg0rHXEk
Wx3cQ5Ey8lNn9nc7sD7ltVLjvyn2lbOZfZTGZKyqvLdzpEpomu7cOiDx7gdB
ZLHEoU1vaydDujVWLEs6n0a2PK1M8CeJbwDnHND5WTPBNZK/LjSU9E06+95D
Hympt8WgDT9Z5BA397q9xsIAzplQAN1yv3BwmmRqs0RGDEipf1UXGdtRj1ud
AWHUUC0fTDRFvEFM9TFr1nDhFLsoCgfEMXSbZ4R41DznFfbDCbAZUJb6JU1g
8hpjZdZ3Ee9eoMjgcEFzKhyg97dp1G+65QFPLIhMiW1gxavdsbyWkW7FwhP1
6wPq6k3tb40uiM/dcd3b77hTF3VFykLfwvbr8W2v8B68EeMFpDYOGmg6y1/f
mRnJWyLGHEn2LXt5BL/ihmrutT+AQK5yZIhAN69RoAFk3Zs4WP1G0rc3M6ph
8YVLszcHvKI5CztWViDlOZww5zFIeSy8KaqbVvXo4nhqByGsfR38DWYmqsrd
RMFb5+oX8TSsFpeuVPQl6sgc6ynX/+hP1SitQZ7o2glsq7Rcm/FUBBmnCLtN
WToC10HJFiywu8vMoCQGmpYl5OQuOek6WjD1/cVZ+iKUBZwT3vGvdwaBRhre
lHWKL4CPKSsbufCJsuVLuWwUvLL+jjNE1NrsSMc/k7BszPWUKjhJEhaLsOTt
PzoCOIJ+w1IFJMiFVgZyX39UeHYwJutf+UEgAa/gMOY/uxMwvlql/F1BARAu
jYVGA4MpKSKo7bWPHlGHHbS6/mpDFw6gF313p144pFHtm/K/BDEZrxi0VzNN
MNUDZxPaGrYdm6BLLEFb6QATLGNiNMkc5HqZx6yo2IbnrGTF1T2xjRYU5pQ0
fzmiTnkgOuGFiDODOX+8HQNZCu+K1rv3Vl13u7MQQAoCdrn/j4Y8mS7siZCk
dTNI9CxZY9qasBI8pBppvtBU576ep05cmEojbaBkK25RIOYwK2SHjQHT8/RB
pNqRukoHpGKAHaOMNk16hWtMVc4KO9yh+FDJnZSH7j6QI9l62NqtmWQZQLDY
C3jmOs2ag5LzNMsHgEoyk5YUJzZF9hr46JOnXbvtLfnHK3icMkreT1sEMNt+
qb+3UQ2vBQKyh4eyW8ByYLB1dEmvmBo0egcs+kG/xyoqfcNTcpx6rfSV9Kef
UB4IizUqrLM0eAAuBLSkcRXidFsQ1wgBBH3gYljC6CHaVAE/WxW+ug7AaYVq
ge1kPXXK4Hq+47Kl1CKGRKht424S9XLgJUDGUXiChCXFujaq3d4EajhG61P9
gANzMTcp09a0b7riDz3OAVlrjvgpeaU9sjg+5HolXMEBooPWbOHkDP0IjBMD
VlMY9gMQZ7I2dnQKLYaqEey71LVex/AIEW6K7PjYkHbTgZIRF+qZn7aPqzyN
ofIW8Hgu9Wip+aJfN0+RzRTRVC2OiVoIL9hhvsDUHqdopR5gtgcHqSwnfNn7
UwmIu6B9jeYhhix/0RHH0gAhAfo0P3ed+VLMcV59/NuCSE7WQZCuK/iBRmec
uWADQN7TeAgwLUJH4d7UuLvK4AhwKVQcyzV+rKaSJVzV2cJSYm2gbH0YYLjA
1ITOsOGkU2+JsLnTOceRw3t+UPcHfjsryqe4q3KttRg+yByV67McOuhWSwvS
MklCFHFKVRhREsgaZ300dOLoOKoTKdR/A5ScPE2yj++8fO7RPgmgF+DDd0rx
fdlYeztRNX4uLL28MsWs1QCviMwOF0L2+YYSFMPxRr6HLZ6AySDndXphbU9U
N8Pe3JD7Qat3cFdGIjye3CddTTjCGbJZbnJ9O5H8FO+V8ZbtY08dh+gpijLU
BhgZITfrpYo/Gx41sMtK7nNxY5vjqyHllw8awoSTSq6Dp0g/lkwvu6elwIAL
8kFf/aHx4KKVBPsZFzRkjx5fXlBYPnO4inDxnz4YfsYyhj79LCgPli/Cerpr
QOlLzuujuZCAzWO6UDAgDUOhH9x5h7p2g9i0foCgU2uh1RV8bxjIAUQF7Rm0
tXkXOjIMfB9pWOb2d4Wv216E8kpuE98SVl52idwLO4R75Pju89vsjnRfTS+2
UPxl31b4H+22CZqqhRWfQ5Os5TnyvzgLfymoEZz1FvgWn+xUQ6q64wf8pSev
6oHwNRglkkviLC78rOibGQBusoHGgREragd5ZXsALsdvhuGKPqIRdEFK08Yo
yevfLZhz4i72SYXrWP/UCMid0VDXhDX/GYvLjvJhSYQM8n6btmJaJNz5U+Zs
yNmRElISbzYA0xet+FUKQXleMEY0WrA+YaCj2HTHAq4PrkHXrcnmr0O7mBKN
TC71tlyG9VPw6JzPbWkPy6LEPdAR+OLo7hGz5aFRVIaPRPoxnswHx7NMpCNj
e7QPEgP3HOehL6mJQKoSIYo5koCk285dTDy94fu4oYCY4BlUYR1/qe1pmlKA
Z8dy3b1Rtovg7oDRcV51xUoJ/NgQq6Z5IsWbJt9bP+9rMg4vvxJirhUCL4DP
bsqTMZR3Tb443EUW7c0NWX3UOCHYI3vyOXux3YimR/eKGo+PM9OmtZhWnaY5
pyjLkUXpiNr/FSoXgdTwnH8K04LLqELFfQkWAsww9ffA95T+Sl9Du8UbHVzN
qciFEFJv9rDZtUaQcbMamxOyzjS2Ex6LmhlURRT4nOguI0g3jQry+0Cfdnf6
3Y19BuHpyWpPFSJ4J0hR9Ch8ecyDFKYFAVX3LcBBCFSUzopJE5gKjZCkif98
WIev9vbT1JAZ0ZfzuBpN0qYz9WwbvslZw4dtTlhgRE9oDDyBNVnj3Sb6aVvz
HADIsXKfXqtPak4RlyknZki55LpQF1RKCfBI25hAUw4OPI6YbVDbH565hApT
0auXZweuJlFfguOTfnjE8Mr/Pn8vBpym+uM3s9GTPs8lsG47xukAxldTXdsO
v9xbdA8Enwru6e9XFzd1IK4jb3xVwHJmr10oJZ9YTXb467oQGle8vOcVAe/4
hLyEZh9zNdLFP3tmoiF3Xr9ZAw3nPGY+gXWMFaIa26SAZMHRJn9za1A9cSaG
8qrrfRC8KrBFl30iK7hCL2BSr4naehCz+4+G2plLMkk3XA1V141twlgoo0zu
R4AvWwRmS9B/8Vehh4mLs2EMtOsHkJ0uP7mnCS7stPoJsa+Y6eGN1VCa8SSv
GHWzlK46MSGEi8JjZIrCt2PDpXpyhAVwiUKnd9sZfRzvQz8xmLYmUs+w6Y72
vJY+RAdMuJmXjkrEt4r45Kftb3TGpgusPPUnsc+FI4Qqqe4+iGg7hJjiVDD8
6yZ4cvsfLEsl7WofN8Kk06HWPpRwNR01YwAbuhyy0b4WseiE5BeB7/MN5yDz
wemAMjc3j36i8p3PHhcJ3fCE2uq4hc2vGuUg1DU27UO7qaAdh/ZfASU3njno
NVOFIxUXjrNWioSLfG5HWZW1bOqEI0yetuQfxNU9Rj992UnGeV94SkVdRM7F
pspQ83K4YPNsldojy6p69RUeCPrpEHIlHVTRvUNhjd8J2ns4SzMwTmpqwQ/p
Fyo42ia37BOcf8bDIPbb51YbA8RPlQYhzxe1urx7dmcMj0goTI8Y1+hY4XCm
5JS/0NfxGRlJ211ToW9cVGzc2ndNfATqCvl/TOWQfHM9p1eWXyncJUwVdbGP
aFIyGr2NN5CbdroE+ZeQE2uyS/d7tcmqAzCZc1ya9/lN030rkww7PfeAFuz9
2GSbRMf0tcQrc0sAhGWYdQxuE1WwoDRATSryoiibLvtNVIk2xUTkkPh1nS/d
D3LmuSymkne3126Qcc1Knq4QCm7c6Rb4+h8YwP9EVcZ7NZhGbqUfMAOMVXre
fn6irL+8OfqO4DBh16W1o4MMqJG4lwF1dT7ExOOV55CigsAUwbVqzPhBHfus
rbgv7sjUwqnFXpEdcJ1I528u2w8qwpxWA4o17orizMQc78prIfkwZdZKsdYr
iN/c+OvvM8A+TwzCKvBcyYXKpoM+hpQpMySl1/k1v5IsaAtRVMLhsnONbnGr
aVGkGa1dl2Me08NeVSZLDs5WF4NU7PsOe+Ufb1TZyE016OqednjBFBvPbSLo
IndSWVCo4DiVhZchatbv3z+GAjnieuKVoyyPc8Dt0hyRgmpsoGHJ5derpa3P
E+sSxakSA2BPcC3z77S5qeYboQoLQolctWJu6ODV6HTvJORS5LfSwdBoD1aa
A+oP5UIgp8jP4LHsWhtSlIsgSHRWKIuIyhSGAMHh9Obf6Ytc1KjuhXXP1+vC
mZXvkuvDLKyTaRQNAnwh5r7Z18UXs6nEMFf12kXz/0LeZcNTYF8pRMs4QCdW
Rzw2OyHyTfvrBFiDuHELIEa0Ft3Vo882Rf4821a9UUGDlmRILeVflJH7MVs4
/j3WOMgm0KsjOZ0k4bYuxtU/HacR+KzQ0y2ykb4GAP43iu4GSe+9516pe3Go
dyRDeLVwf41n7NhufEqbxYdJTSJnNUzmpKFAo1jDtLj8a17P3oBrtsIj3J3H
ww7JTZR9iw60Xf3iFVyo2PV9pwEsHDdPjwOqYbRCXHsD449Pv1mZCZ2B/wZu
/GnXNJqjBFtGREQ7iVxdG7b+xEc0LMu2XuhFxtDq1A1+3/8ZVqhFOMjUfkZi
IXlqf2MTc0kjaL1gNf06hhXz5jopEyWKZ9wMx84mpuFs/PaCNO/RajB6Upm5
hFoWBefBlyLxLDVWfvvS2gbh8v56HPSqWg/toSpyK+owNEjYhTiOyfo6NPCd
gjRWbgP2ZLXsF0qB7GQ+NMJP4j08cjvxtXG7Mbvwy+ACmodGVi/rucrd03Tk
iLHJtvuKXzfwpkKKmY3wJzYIGfB3LeGZCb2/UH6CgXaB4CsPUnEfonByqPGc
ij0fY8cam5Uyy9v1vncobQYnQGvYGNXuGyHfHJapO+lvo6QXyUz0F6LzmZBT
dH98RPj9gnQH/hsL/rCPXwk7/q6Vaf8cIU509SvsjQLRyhNto8OYs5X2s7bD
d3PcZZiNJkkt2qODWtOVm+PdJdaHOLvPltaj4g8rryeRDGX6pl4rXgFoPBVF
7eRKrjNKzPJpkOsRIyYH2S+iOTkgY00Kkn6uAq9xN+Fpj20vaPlV/GfwPwQV
GvR0gfaQTaL8wMuExuCUTPZiKDaknYofBEFJ35bYGFCfAL6q9FCbV0Eb3pa9
oboKzF17N+lO34jmbH9QQgeec+cGSw1Sgr2iEYDPhsSm1NXaaNsJgCRjsOAJ
K79F/2VVIqIIRliJU7yUAU/1VcrQFneVedjUWoyBVBtBmBq7FvpgodDYrPF/
jSmdmI6Kx8r2lDsj+0RFT/3CZV6KrCWHqSsLvIvLAWLc/jfpDawQOjO/8tHN
JbUjqfyh2gtK3/zXcNVkQgRsbKApHrBjs8IdWYXQj5PSpufZwE8FCc/xEyts
6BKReRHf585vlJASPouEKWbvpwWQB5WjLMqga+qwb7h2dvLF3o86URmEXJc+
Mp4z/59Aty8l95G9gv8J+AxuzBASOOERp6RTH1tkzMubFv6FC/Go9J2sJq8q
dKoBT/DrwbbMEKuFcbWcstJv8oC/zyO4bt400nUzdMd9f5a5UEFPAsyJRYFl
kD3+lsdJhqiCKB7QTeFbsFi8TkW951c6oh8O0v0QQGvSnyEN2XKVHJ+8wlzx
olpLGRh7vkTqN7OciK5Y8rSe1gay3rdFP6hW3RQnkGEMqJWkt7CaeggVxGZj
l6SJmpv7jfF4sL/mf0ERK0HJTSfonh384FvIg2YsIEg9gtt8szugjR6L3HGJ
4VWVbNhDRgMOshqO00+sq36mpm2ulaxCBcZUmURHtiHUojBT744SuUdi/YAs
8cxlsGuVaj0GOcnmzRNf8U8VNIhvzBHo5cdRdOv+3RuCsQofyQ5EAKVD8Xe2
5xEpvpiQ0YiRC41k+8cST/0u6LS46BaXlJxnIN45l5wBx8LNrV2M8uIqmEd9
ki3hN9i/xjoMyKGSsxGDWGjU3fUYWoQWjLNviKCDyJg5Q7tnE+cfKz1g+BeY
Z7awUTC8GPJ9Hnm9Dn9rw5gBGZ087gVc46y4GsXThV2QX1Wf5PluEpmMqXrW
D3r/RzMJiSouIDp4giVnUC1FdH51OoJ9EkS9xIcfiSrN2flYeV/82gYXGIB0
aFM1oNdOMlr8Qmi4UkvzNKhsrCwkRWOCcY51PL3AZ98KRkUWJ4EL/IUUtv+3
5gok/Pg+129btaHw6oq9CsXSLQzvVaIrNMbcJ4AfELjadLCh6lVgoB+qd6sd
O5AcGcX5VZXMijV1QRBCzfGNVDtItUQ15pnoZoR4Q1fiVc3cOo5wHj5QMWxn
hNoBXx6RBtE7/xKrgzwgc9WtuYdKjovS1CbaI0USooZWrDjWbBwt17wQSdgr
Ds7BDWeAndpai+g27GK+YFGSDwWe61px9WoYlofWbYohKbFu4vQaBryyiegn
5u/1jRm1fm7lQxXkLDZXK1Oms4IH6hR8TkipwOh58OCyGSnA2lODd9DjsSat
TZIjAE3Z+7BxNGSE+272RFCVRd7v79jA9Gu7uGkzpCSYVRsxOFpZfB0KVOCB
pU5a1Vc0xHTJCJncXV4YcFkV7YGqnz5+Un8xaneiyS7acrInemVv3oiOcKG4
HenBxxRegu0yjVvskclU/vAtsLfAM4adOp4dVpX9/C8U8TCxh90A3oGiXrVu
POwwRpEy0YS6bm0zwCIzgUpPQjg7Q53+vS5G++y8Hp74lODOBIn4ttl1EyyM
hecv9DRMVf2bnDNDgx7WMYP4TT106eIngIyuRKovpFDo7MULciwyl7kXUyC0
tzjbqCHfuDN3sTfGvt1+9e//6Pe1DJJIcOf5BeIAdNIaA61aG2nEmi7xVmS8
xN1kmaXiGpf5RW2VOGy8uoQs5znMje7SgcsrXBmAIcFPJBnPFrcCVm4s9GjU
ejLIs+hK6et2Ge6+28wTcIfyZFofh3umdOdFuo+X6ZZ2Bl/gDz2ACwMrfr6l
9RW2AzeCGH7k/2r7QLw/Y/ap4CwHrK4z+ijGQlYMAuL4Vxbntg+YcqKylNp1
nm5DQQAh66RGeVo9KHO8b5GmlH8eI8MNjTNpPg+KXfp7XFbE+G490IsHoG+g
g3wsAFu9dTDRqHHKYi6yYj7J3asVR49WdY5yboHzzl3WZWcuD4DWJDBb1P0x
z0JH1EJKQUuD2s0ft938CKAMJXULYwCRd06Q8NtfKLk17U9Tu2xEGiczla5y
fsb69NgVQgEylQrtaU+GXJ4fYB7RejUPFVzVoo3ZHiOJ1khjxy8WxNNQdez4
Ove0+rMmz09oY4WdJZHX0Sdx6Sp4YjSzpsI5bqLAdN4H6Ti9W4097A/DcQ9I
gqfrEu0f+b4VsZiZ4qSSai49V0aDCouwYFZRugSABEz4poIclqDxHZqtwa8d
C6KNLIwqnijMzfIY5WLPfB/4eabJJGicElrJa8UbS5ty/ZZI4U2UI/Mi0S/Q
cS9EO/dlBMRceerkgqiTKDa4PsywlhtJmtCPBL9ZP+limctdTZ9oumgwRsa2
aEJzPhLYUnfJeiqCMnlKjI1lYOBpAPP3D7aWFx0siDVH6dJr+U1SIX4/9FIt
nDMa2/BMbN6S8KR/jU+cX+yQio6wECBXEfwUkil0XI3nEHYdKrpKzIcKXPuR
GMgnSSoCHyUSSqOeJ6SEnO4SjZXFNDZKO9Qja7Q6nPB49FSV8Mo7mANZKIGH
noh4jwqXrMmu5AL3hL47e84tMYDlA7UV4XmGp833/5Lmy11Bdfg4YFAjRgLs
3MzwYwg1DMXWtzW2DfjsMLDC5N+BIi/Vzj/D4LJByziK7FEnJGLrzIqfFijA
UgYOcAEC+4BB5QOrmk2H1WzQksLALVqvvBS7damtK97un2T+xUkhsUlH7L8U
LdrLtXRLuoYKCNgYAjXqldVCETRpLMpuEKTx/Hc+DZgIvWUJXJ5JPhC0rLM9
pPzskjoBYuPXWHAPA2cd0oGGL9SWYDXQ0zg3rn+95oIPhLrlZxCcpXNEepye
ubyerBSsa+7hdB8aow5Q2EQDXhGyoEjb0w/XBJDlVpDdZWW2uAX2B+DfEK63
IJgwahMFDFVs0EgJ1cMwMU0yPdL53EbaEqtfR5CCCgleX/DYTLL0BiH1+brJ
/03nBUmewbVwTZPxoBOy4sOzGodrokAZA4d5pmJSipGq++8Nz3fK7QcKdSDs
H5/3seBeS/Gi7ixBuetpCWI+U4PVG7iF1er92fSJw8fpf+avd2FryUHqUMVn
w+pjgsGiWmk+rspfRtZDYo6hFA/l0T+M0ymUtLWkrEuISf5sUHkZntMJI2d9
NtcoWfokHdRZOU7bXMaTXIyoG3Ha1eYg+k47RTQpEYhU83tU8Xf9y2HlXMXv
io6JTDnFFRt0J5tPPQ4PjGwL6uklhIlNpqysrflFOhs5DG5cPsAxayxKWE7P
JV6Qwf0JacH1BhGJEqKWNfNu5VehwIhAY9CfMjsq7abfHp3WwfuTU9Qw8zP6
zwSITSJqVbyeocZ6vorT4kHgadki8yzhsq2Fu0ry+YAh1y3D0GoSs4NI8dSe
ePVNo9LdWOraoMtuLMsc54BqXeeDIjHRoO2r/Be5qCd2CF23I82DP7BcuuFF
89PgimIrlNsYc4vZlDtuu7ZJwdbqgC3zZR7swUVDI28szuQhuRTTezL68EPF
qAMaphJPTl7DnaYDD0ohGCt09HZzCy4oJGPDR050FGESJu6i5cUW44gcic9R
beFVJlwMPLe6IpMoXK5QKIOFM7aLbpXGmN/DzZKCf8l7hIat8zW4qTwrxGK2
MN+GCCLGvcujuhszYnI9+Gas+nSrRTh4AuzeUCAmAl9beizbiN0VtxXabEfc
rSvzkfVEzV1B2zZMuSHoRFi82FlJWIGRf2Kk45RU+GX0Vo54ws6FDN+lRbh8
o0/TsedrIKLjOAJZ1ahzsR+vlNC8la92/JaVMCzHwdxbpRrU+OSe9simWBDf
kdm5MyhqYUC0/5F0lZPcU/45wdsQRi4PVwTYezyWvCLdMIrVSGdzhHXx6Nky
i8xSJuT5k5HH/HZ5fsC+Ft9z6uipRbC1jtdil2KMybbN6fHNLn99LVjSo/dM
Q9kioFB4hCPn0JFJGi4rJ4nNufjMiHCkqH8kq/PK3YvjZb+7ge+F1l5t3f0G
N1n7XwIw7G6vb25d2vZmqjkdN7GtsZeddtju/UsFVNnLVzp+0qAE76rzaSn3
M68pK5VAi1QgdEyAoHs1c4yzW8zMoWdqTJzS0Yb0d2ieWzFj8igayj1VPlgf
y2U3fx7j/rUGM2EvXkkkLQ242kzBPRgRSMYJY+L8maZYHJhzW5HUx0lWUtQM
siwTNGMQ+HPbPJbwf/URfv9srW08vh0YPmgkguvxHvufZ14fZK82BopC6ih/
3HvjwmHidlUQTgEpYatOxoeIv9Vs7BPYzjJkYLVwJVtqO/NY/cNbsbtX9i3C
YCwW27f+N9nIVNnDAe0NkVQTrwcO6xJdMLVFeKXG1bxd3ql4CTasBju5M9IB
nR6DllDrhR2q63gRfM0L0ldQWUMGsmFaUOhwYTh7maKU7lOc6dutX8sYi+pg
NJ5ih/mOLJ92h0O+n5y8lYPorvMYx16vToXBVRMT6CzSu4aeoAur+t++Gl4p
mn4p3S7QH7wiLwX2FVdLgvtM6/N9z0hWskpkrSs+qIl6OlAsUHF+nYeGpfBU
Cnp0Lw92YGNQRp7P63tAqDh16NA69eKQ+LLKXvSrZ1/9hsOVq+z72QTCAY1f
UJYxAeTYl1osprWaHIJxYmzlNZfOtiQ+lbjUaLYCMh8Zlsm/Wblyg69Lo5QN
x+W95TNn9DWWkukAMVF70Sqx28khSsB+SXRX027xE3C3SCCgEXY+MRlinxAQ
nDZARliD8FqE5S/h+wYuJOkKhqhaJb8SXm2TvI2bD142uZOCjXh9JCnXe9ny
PHnS5/RwYeJQpGGF9GfC+sd1PzhYn4fKnbjk6zHq/nQD1tE47fkxtYYv4lDY
ZypYFWSk0NhipBxKOgLIl8ZZuiFgVnX78WkAUMBMwK7tdr3IaLPJTmOCLrdf
qZTEcQOz/tlULDCXCPqAYRiehVYUR14d+coHaO4RNouWkBJHmeCDRz7OYJVM
YsjZg8oxxjfQ/bJUwj/XZ4Nor74rKwNBBhjFY6QV51bavcQ/S4kh7eInee89
X/kx4lThGqMs0oQsNU6kFmr+1yi/vATsH+DEgDZZwYBTTEDpGk4k0ZWGtUzX
kK0nWsem84HjFhjA1GRlYD8Vj59XsakPQ5/A4quMcQuuTfsCYdHQyQEh1sZA
uKPyx96qlbcks++y512daicG+jURN1qi6q/Ci6zDPCTyLsgMEC/cMP6JxZPB
YWKG/u32iEGVa1r7VjP3bLta0lQbIpbA2NMTSTGAW2f5trEuCPZsjkTATHUj
YNJoOLesHxcWg28OquGHF2hXXrcZzhi4VC0gbIWjSZNXJwUgkbDOP8gGXjGt
Bntx2hxBYNU1e4uexegzWiNjvWol5Q8O32Yqi8LCf8WMn6t1/MpBhH2pWY5l
fdf/AzdzKoAeresZO8OBtu3vpvgFHSgt7M4jlR0egNl2jhfydXnLafeaPbUP
WzmxdPt5V6D1Te71HTq6n4Fl9DvfcYkVPWyFvh7Ndyj3XBM5G42iwWk83ypt
Q9r2d71TB598kb10DBHUUMOLwxmxSuUzMBkGnWBV6OdIR8HowxrPy6EZItFo
qw7RnKLGXow7myMtjCx/KJnm6iYpTthTx3miQrbakAUT1OYKraoB4CPGqOkD
oGv2YbqmWFvju9DhjQ6BRktIwJZiu07Wl0FDRfX78k4p21fQFpvqf+WGutsL
e0NzdvodcAF1G+ShmCTG8wm7mr+3LgmPHSx/RJCjd7//m0vjyzL+ndlayTNI
Fe649R/o8djbSniTf3jBEo85jdTvlFkoimiPyX7m1qjOaTmdVXl0Bz+woBkE
2uuioDpPOIzDELw1u2Yeqp/z1+JOLux1r7ulg72qsXXHU5PbzcAXVftDRS/2
8jn8Gp/dZhwZ/6qec2kuD9fWzEFyy7LAHyPOPNNvw28fndC8fO9N6NeCGeUQ
8gMsdZh4Qh1Yo44XLdgb8CvqDExeFnmR9FJKtUFcJSZrNefr/2sRGvWYIP1d
wEXyBgtx1hNfoUuS72SPypaRvooekRn3dhxPmJUndSQvxQVJSgqwt+l1Fce0
pIL4X35gMqk2R9/wRcsaUWWANXOfdMZMKnGJ0TizRSo822HW8VVPbeSe6ELp
3w4FEebD2+2z1oeIiaxFnINr7IZ0W68dHCy+d9d8EUeGTgxvYqhEMEQRQSqT
xDWbLJrS011cqzTVAcStUmTjmvs1MK8au8/nqMp6bir/gCqkqQPZHuqeCDsu
dDPCjaKFaK+XSRP617gPRjdZRbR7wUb0srQl19sdXlfHgKEIBb1rz2A4+6lv
nWFA+k5MsvLM2Sl0iwZjmF0Nxsgpk3kdCJWE025lVs5FCk/30tvPmU63USme
slbp0wfQmlYgSC+u9Yz5UwIWNrTLryo0U6LzettlrG3kvoTDOXhDWiYUVS4L
/X8RVgZciVJ+E06OrfjPAhCb+D4U+yKubjuNfmqV4Ki41N/JjTXFZybD84XE
2Fa1JMM6zxzvBFVfOhHawJAFpQw0YC5zbtExzB8XwwWNL2+RwTImLLfybNcc
yMkkBaqmomi1156wrNoCVnpEnZraDEQEI0pn52+9Smo6jMZYJHQiyB2fXBr0
6KTpAOZtrsPVuM78H12ZNNImRNjRdv96fFxCzPcV6h+jhJidsFcqKymOps/H
DC4VCdCg3+woR5/rq8awCfa13wILNfJ8Lwnxud/kQZMiAy759tfVH/Fjnfnz
xFytFCRI+gzq3oj5utJCyjyxPod/BfSvflUZrNzMLsPhmUmR5tadyHRF80iU
l6dTooXehjMPIv9lttdOJjnHeWiPCP7hleo28MlxGU1JSTzTPKIvQsIV4qAv
+WRuBi43gJSXDDUq8ta9vi8bjOHZWrL3Ny5yXXykdxTzNkQGnCMQpAVeT073
Nj/cNxX7AVzrC6vpbW+06XxboL/U8R4NxlwwTcpg/02ZyfpSdT3y6RevYmhd
3i5HLICWlSnapEdC5Q47UrqSh7lFEQU8e87ig60efi8G5PRxEaIobb3Pl8if
O4PQzwaVo3R1v5X6UTpCr2drIrDDCOes7V2gXA6WlwuH+i7hymBjFK0wYSBI
XW/wGqfKZrS6WwwQbUvH9xtOkgxdl85dIGeagh5Mseeoj8NOBjx+znkeflyh
rdKltsIuvUoyEjcjFAtUu4URoaxg77dOZtNVqet5OPmLsNjrs+zJWOvofv8J
Ldzj6vPbDxmySm6+K+J5EdQ5Kt3ZphO+jiCOfpGGIlic6H944m/1764lLhck
LB8YC59wddhL3b0XbqtRyjZKSJ+E8F+bfF7aYzr5ss85wQ8QhOSSbb7aKXDK
RGdYpfyOD5S5IId94IIrbwQxPZ9/uMPj86SCcrrDG0bGedcjyvFqOHfP5Tz4
sZOR/qaWl5i+5XLJx4HwQEj7U3zPJbbQVJJIiH2NkVuEBG5ouD+x59LZ/zKq
0WqGhWLIJYg4CquLAWdmbCeNXEcI4/R6ck3OBotgznvZOj+MxO27l2tvZ2H5
rIuxUyHd9yT9Q9e5wpv4X6dnlLH01dT3BElPNqR++IwkgcCsbab8Xocc6H63
/n1M9Iu4F/sBPQoNL8hhfIZrK7TSQf/x8XUVrbfMiWQ4RP1W9nBKZyu197Hg
TZtf1p2FCiz9NTEaftzumwygBnzZtAvjBw9kHPeqKsZrjVVV3zJEwBWbCi6R
4Y+4mY+6nN9l18z1m4U3rAHxTXzsXI5pMPSco3AFhOKUWbQOC93semdkBtyl
2ef2PhT12J8NFhnojxUvv7cDd+LIF3Du7Q23zR+MqnJm18/LVQMW5zk+e3Dl
bDabIRfM4GS6OJ01/JCfLBq6H+Kk0RbCzU0l+WJoKIM8FW5FX+YDMmgCWugf
NZmgFMzzUIkkvWkgZaHhqBqF6ZS+XcNnvOINDNuMSgX4cONOisXiEqb+ETs2
aE4yFbN7bJUkx9AyyG4hiR7RpTEoRaZCO5jiADoZMwY8m1oGDstH3ESihCHt
djjLSt5drgMpedhAW8UdXKXti//haXijIsZHKR+YEaIa59py7nTE3owoIw0W
RwZ/vu2TB8Jc+NAdiUyB18QYwarDPKe6s4IGN0xPO2xFqUOXLHlmvL9ykuQt
8HZfLD/W1mzvBKNvwCi4kRSOEvyLG8yt7A7OVLpaJEgY1/p1P1DR6i4TQpvW
wbARL+6Nzb34rCGO0NkHCTSDMbkO8WGoRQYsAzLglk4mGE5Nv7A9WF7HgXKR
x0eeErFb3wo1rWiiKAnbw8o/OeoXPttJHiPuhieW8yoE97YVyfOfFeaQ+sNn
KGxtU7l4hHWBfCDUKUAVOLbqwcbsTdC3cdawy152YHPvVBucjv+y31C1y1wE
r1zRRI2KBbBFsv+5kRIfAN2jztWOYVQXvm1ax46FXrpJ6PGyovlBIacU1U5j
hgZrRqfrgopZSy+O8G0DWxJYqb6pJ9B5vQ2MmCQTWg6Tnjo64LmnO/st7Lbh
D7cQXkdLhLfJaUopClGuevRYYv5Cw/dXDr7J/uMn5jmQGk/MTl6B1WFzBxVC
ZwckXEy+0gCWPY4JlJIgY0nqH2hYkETcnCVMBZMV/4RPmluaxiFZrdm4fY9Q
FPYDLq0/CsbriMs9gst1y4V7oXTXs3tzu1//QuK3q4auSfvUUZG89BUzHR5y
H45ReHyHpViZ3PD6vTlL82r4XV8brP00Axp7dKUExHR3GgZ9qKv8IdbQKZg4
hYES7eR7/+dTN/bH1PUlC7C+iqRUHjFE8K8JfpSekeAbHgSQpLw3cgg5cAqF
R3wZL7iGJwEHPOao9/afcfZcf7Ll81Uzgdns4lV4WtwVAZtXc4viNT6PcKXD
TMTrzNXagKrML79qA0q3X2x4AI7PGMQxXaoLZxIJbH81xks1tydU9quy5zxf
DiGYKSxfLgZuXhCp2icivmmLvTHzaWahocErj9gfybdU8ehZjFlbSlog8klD
fXFIEs6s8+5iUpvIIWf1FcOAiXB2/XKEyiwDzNNzsSo60svHTxkRKzlUrXYb
I8d3UuwSjM4VknHEQnJ/YNHE15KtnFphOZJY90hLetwNr2uOPrqx+BuLCNjf
dEwmKDiNR1MaEYOBHa5Yy30QcE6KkAF4lnJwrKqIvzw2+l93NwTz6TIe+ZDa
pFlk7J8zBotFNZKlln7IU83rgy/pttuEs/Zqe3noCy4Hn5IBOMv+q7JIAuMR
hSlc96tRGbq8iZJCJFCmJKoOS4X5jachZtT+x3vJLmNrpgahrch/FrVqUMUQ
5jjx6TBsQqUT5VNOkkTozXz3p9MF4vqhOcrXs5+APlTIahJF+kD0h27qawtj
fcjVrga1MxCvbCm+CXub9Nw7+vAqZpcYSaS2OP7WiH02mCK0N6XMhqi2ZKm+
Q2MZlLKxI+iw62+r1rxeiz7hKbsjx2BDI0GU9Kg8xfRASUfhHHYqs5fbNWGJ
KzYyboh+dyGNmf1pYk8KBWWkEbYR4VRr2szyLjv7sC8wvNT7xpkUD7B95KGN
Oh7kJn607vWHdUvqXhR+oE5jI+CL01da2zXmSUGUFMXoPVTnjkPz7SETpLZo
ilzBjmhUMPaDjAjSL1DmB/QaKkCgwbrXn3zMSEClGNeuk8tcuJla+Tigf89d
la03sBOAojlHJvxP41UVXFntmQ7xx0eovvWwvfIMQsYuWZvKJBMmbPB26fBZ
0KpOwgEjlnEWYhv+kkrPIgpNYLZ19DBo7Dy1hsG5KUtozQ807cw//iPisbpG
zWXH2VSlILlQVAvqUWh4LO7QRvr7UtNXX/MGGJpcBlpZNhSfH+SrgSopDb3q
VJyBVQ6X+QYS3jZdKAFbl6U3CQCA/Tlwjke60qVF+0CF2+/e4vtpAZ16Lh9Z
nJicseFwhxBZpA1ufmuYEzVHTMTBboqeXYlmHTnUJrnlo3BgABnvFa1NQ5FO
Rz/FlDk1nJBjzq3cOJEcsOZm9ilD8sCKHz5jpMWhMRPXGIZbU0fkKbzx5vjp
0Y5Bf9BafKp82ShPdp9M/kCVdygjA4O+U3M/6Ci8umhRvXaz+g1xYfLT7cXo
78xms+g7hzLilvSWUtCkpxdJjW2Gx5T3c4KRCwobJuc3UjiM6jQh7ed0paIp
EcFzGnNYHff6jtwDBKsxh89q4sA1xX711eRMb/eohxDq55vUE+uFh2OddjzN
HoTEN8klaVxxhSLSJMlH4Oa5e7A2jUlPi//HbArBUHVhaXuTDKHJ/x0vkcnt
DHOtLVZcKq8R5QX75RHpCQOVIw5PH+AoGhcjgztQ/riwKpTorfO9sb31S8Vl
+LyZvHwZyXzzlbOa3P2xbh80WuXkVpPQUqpAOdOYtJL8rVsrTjsxBgQbS1Iy
AMMuDL+UZqEmMrKbSqHajC4acMI639DPatU4jiFV0ajYnP4jjqVWoibJQByo
qZF4OZWTManSZ60Hz2H3MpNOTE0YnrUs+tlUOblyfovQQU0gBXrkZWkLpvRz
PHirpubuHWaJgXeSF091x8P4HTI+drsr4IqUEhRyKwFEHBRznG2xuzIs6gWE
jrZr5Jrd2zIQTyjLgz25G8IuRepiOirDdhak5/O7Axkmmk/W+CW7ejDiOmQ9
b5o8qNgcuG83DGvU6nSulQkKAO+Fns5HcN6iyZyDWU3VX/XGbp/gEI/wPDHq
fDOD7DZes2+64pwSsfbB9sKOfSDakV2XzQH88GAj9scqaDZDZxvlLOhELoIN
2HmzdJgPI5QC3wheWTyoK3l7vNHMZ9eJZ4i2LEWmAvoLOetUdzNmGptLxCBQ
aHAKhDyj6DkIN2Q2rG+lE+zb2/xkUtuqUgDP5mHtcNpptgP7A0XQBbCotnT5
4VMFcynvzAJ7WXolkUkr9UBBkFSxtVyZEVGlml8oR3iAec862hR4fRneI/Fo
wtLEKxpk8/nuZrM9DJll33uZEvPk/QcBaUUexEgXLwjixcwYjW4d+bbVtXcX
Y2abPHiy7WitlwuSnEism3lNpesyni/sY90OYphkU7FxwXwjuVNCjrziHRgw
+sh0gtU0KRCUztsCr4gdJ+exY71/Hn5CUBc9ZaTU1ZizXyqfGvhskCw6pZLZ
qD+R6XRbrqeo505ohoFZ5zJMSRSu8law1AgN3hO9nWRXEM91sTVKrReFlgxj
OTHalrUwfYLP2TkX0SCOvrApyvjToVlbobD1WOov14b2ajBBz3SCYDQV74+R
zzHl+tbhRJQ8oGt40LMpln67n6QDmMbb3rT+pVswJ7qEbwaMuftvcuEmVLev
GOcrIZ1yaDOxMh12GI4Ix8oP20gdhnv9xobH8kHQ0+HzvdA/V/Wk7BLR7ajj
H1wK0Mt+mXKhGY+wXDmig850Oq+KNIX/fIfi2q6t9NFe8AnJ30253S1poup+
s47I4wrw2Nc2MdAptVjbH3x4tikl7uQHSpA5JXuX16bo9lWvAlUvq9waS6rh
kqqyV2z4gzRzAPTGuVbXSbDpX5NLGArw2wYuceaklNwVR5dzN0XkFck81vxS
FtdgAValvv9KSq+4C2R5zgXEC7pTZKg0MReiCbeI1+ljKbjklFq8qsD5oW9P
Gd6Ms2Nn5K6WFHVw0hWrFkj88gpcZuHRVSX9BjRO7UEHDqrBCR6syHcb3Tt6
A1/SXJet8uRoqdTzHQQa+TKGwPldYvvt4JqVyJmFrtasOPEi9JFbBtErwBO5
kj8Ks9rMF9OY9WAWSD1MULAppOh3b4HQSYcBxu6L8dk+pYKJ0kUGe8+BeWs3
x7HbcKNb1pB/Ip1idxftam7o1EMqPmhYNs9E8LgpWPlbt2LOk6j/8X3MbVhD
4/Kf8+EfqX3N8Xt7w6czBEdLTIIgHIB9pfOan5Vb5PzvTzS25WgPhF2c3TTd
rHhJASKy/FbT2Io9mw+4x7E7YoNc1A855/RMlRrM2M2vKQe6n1sedNjN7zy6
SUap2k8abvRyeUAhY5K1jR0vgrjTSkm46+xtbI5FaD+3MzYXfPSifkdukIU3
O7lRLbuLKkx6SZNupz2CVXWnP5U+S0cJSJ0OTLwJr8mIKtsyaxKNGCeAGPjh
9FxGB6VawR1iyn7Qj9IVjDgKdbustTbwIUo7T/udGcmeGTCmt+SE9Udkr+qI
MmckASbiG2AhUtqsJIQi1hFLZKr37TyEweM08qFS0Hjg8JrabxXalUwslvap
jq14bH/T3fqDzy7caZzPnCifnhZZBoBm97fDJlnx2LfEHmieryFcVy0kBT7m
UiH6H3ua49tMIKirK31idkSsz7dEyqDZ1pSZ1iqmp85YGia4v3pRE0r+FfAR
suxK7JwJb43wFhuHjR8PkORh8MsR6Fcfq9XEzSslOkYcL3FVLYno43G32lz6
wTm00kZQZL496p4/TArVO+UVbI6Lnm8TXlJOJgU79a6Uiho6T2JLLW+1hQnk
PZFgZsP93T9dTHu0SpxYZv6+HpPlaAFLpxkQm8nmovNGp53NrCPu+OGBjTmn
1hVIUNR0iQ5nEUMkdoHp9YLlMlIkPj7fFNY07yf2/JdWlhL0Un6hvniQk//L
nqfov4/JElUhNUu/aYO2CBtNrf1szfs+IsPw0/MCpVRoHSkj2ypf4qwyjMJh
OJDChD/6u8/TJQJjezXY74oHqr2AfqhKGqa/FUcWfeCSwmAHEkiQGsgbwTqW
kvqUVok/8oHJt8LC+HQNnMKlFQ/KFaVYqjvdNP8uX3WrAxck8rCba/hfmpDG
hA/cx9vuGjW4Bm0KgO1j8Gwq1+3MzoOH09gwcnPGxd0vj50dF0nsHAVC59jB
0Cy79XKbaz8iUaAU2oc5/trxJPfiepENSHkbftxTTAba1S2DpZYCO3HnsHN2
KoQIoLA8GPrb3H9g55kEJv/Z+BA3n+dZuHAefvwlkb3znPRVz4FDtZgtzpPI
4MEoH4jNHbUQiBGXvEvnwhnymhiVZmGUADL6HPqTCfhXXE8oTOFSfE8DTg9T
OKYv4hmfl4fFFWgn6Su5DlB8vtWid+38Gxh+R2+E36vLdizhhr6phtXlc9oS
wDnElWakuoodU98KrDF7fTLcfoK6gx4/XdmUE5qLC+g8ptKTQouipcx04J1b
l3sgyrISxeXhWDWeXaPn3++n7fYryWyv4VjAZjm4abzZBJw70rJqHzQ735a4
SRHA80ES92JdHoP6peX5/LYoVhwLZdx5TSTVY1u8F1YL0QlWzCh/3+9Jxlm6
6QHokoDFUn/pS7M0HWRKS9Vo9/O+KYs2NnB5mGywt/JpmAKbJDHgYlodHWPW
mxUxUMwphQAwKnPNVu6Uig9lzm97x7FRki0YKSXJitWpPp8Y6O6F+9DmvL3s
/WA7fGxP0UrIj9eGJmAPU/SyvCVlX5dS5Hwm0qAdP564loRXxGNz/lQXrRcM
eQdQZaySZaID98TwypH5m3U3ott2wlsGxpS4H+IfgySZHsbTfc79VTvNfeEw
gdXFtwoGKyRFTi3wic/hgYFvFpDZgmTcYSuoxUASkk+KeL7xR5H00oqnkomJ
oMARill3+8foZ24LRegVwnhw2eOSE9siMrG8EFBec2xFfP3MQyAV/sK/DQlf
IUzQRRNU01O8/RQyE6ZjZCf8ePYTDRb6jD97l8i7qLKmbISardqYg15hgq0m
xeTra+EQofHEKWgr9g+Ez85MA0WgG95iuu7qWv+Skj9BNYAymfIbQx9xUw4P
G5BfcgUnDPWwfIBfa5bO1f9Bo/fexqTYFJrgV/JNQ9cGpoK/02ssa7bKYma8
fkvF/LnHiInWhRGw7x/mk6IDJLw3urQXlBAvenfng9oLHOpVJqtfH7WegVm+
H4bPybNSK3lR2O22LCfr5xxG6uwyo6cGbzECMQtGHesae2YQVaLOeSB570DL
hbuBaZ9gx0v4VbAP9peIoGY9nu3NncmHSbOF10w7dD1XccbbIyzD+ztewqCz
Wah3Hl5evBRu5bGfPcxqgBuzIC5Iif0M0O2rHhLWhjq4jutD++0tDEWQqMYf
LPj8bU2iXuOTXwJXjhE6UskCRfsXxoWXN4fJlPdWSUZmLTxse3mgsK+N59+2
jAOxU4VnQQTy9nMh+0h3jJ5Vz8mWRHME6rCWLPYQpaxXQ+ug5uU+U0ppAno1
eZobPjjxXfJybjgT7hJGn+SAvwAXBT0tjldOXYGwSfhIPbHqgzK5KQ5f7LPC
I7vQuVxx4Ke9aWvsfexkKrswlGyyzVea3pA/Ry9/PsJSthXffCFYykxDKt9f
yqcnhIYfTuiUWpIpZtgKomzlzbtufG76mAEosE6pHwlwKVCfDDReth3C3bBt
03PCUA/+kT/Ywq6kF+u399oMFI2OD0qLTkUgdhL7H19YqB1wRixVAfi1gLbE
u81lMEYm0Jj35D7dihQhd2uoVrRPsHeutgiNYEJv3lTtinyZ2DHykM1SNmO0
QPGHFWGSTmJUpvsTXmLeYXuIs5EBvBBnUjjmQTWlCvdajjK33EDgd8M54/kb
T19S5RlnK5z/1+JEM27pej490Ud2o+5KvvWTqiRAF48YJOkpdUCHN8PmQByg
y9YHr6erLprmctEIdrEyE3f9/oisGThdKlyRL44caQxL361eh0O1Nwm43zIy
PFzhpFaov0Yd25ivAWbjmYtqZWe3BVmQltS0axS/hPaq9ndEBaPSqnK5froP
TEv0sCnb7aFgvkw482Xt8QYltydsx/6BYUn8V6j0COaP6rTHC17o5Cle+71P
A2bby7yI5NabjN7GNjgiY9k7t1gm2kZfMmz62u+jI3x12rEneqiHBWManFd7
KmwslFH3gdEgmsVUHkAKeLoZkFgwXLYpBHiEz+Q/AnCe1jV6eL9AbzuMLo7I
bJr1THB+F4gykmnuszy7HHJ/kGaeCX4B6vYRlOO+lrvJVHy4/TykFBLlMiJy
sZSg80Z0JXsk68ypzraBG2NMkHrEU/CySR/EeFmpHMSklMdbMMwJZWDobOC2
DBhrJhWqqjeKesfS7ibN0vJRUXeBjvQ1DF4vKjDBFVVqDso7Hw2NWX2X8x7h
cb/StTUrndaGja2ixRqWUu3nRkxaqOf8IAlSzzsNgzH03h+pUvBrfvOJ3m6q
aBKrSdZM/saeGUq4Z6ky9Xnyd6xmdJSR4I5/+5CqRVjsIZfCTV/0q/2wYSvU
PpJcccCaVrqVC3HjZVMBeRIxAC6Z6qTrL5NrlwwcE3H3fFNq8oSj4RH/Ov7V
BABFckTCkFVODgfN+kdZQx96taxJq86yf2TlJKv8+jWG7qcsHg2Pm9bL7A+b
IdzJtLQo83QUXYBX5eHU0xfhVSBPB0pxmtCr47vajVr41/dGa7kW7z2SCYyz
2stsiEaiETPNIK7mYmBZ06EwvASUfGImF6Zp6dU2rHPv4aaaCFTxsuXr/bfw
PBAqKTrm9W/uJlZsoEIKmv7dgk/tvf6ZJXfjtA4jz/y4baMIX+KUJ9CRsI6F
mVcMJEG+nTUySh733yi2G3m3Wg6Av5axu8ntl97v9CNSgOnMYSsz+U1yW3UF
WJuV2g4ilqdgH2vsHQVH2BQBvMgjbRYLF4AnT9bKa1HSHFipmiS/forSAY0Y
zH0FXZR/ZuDt/qR8lUKTUzhPo62Xxg8DApy+aX/sO2PG0tIKCqqGKjnvl47e
tLCANeYS+NDQsPolL5EYiqO99UNLb/BX9GkSqFDW9LN0RIVotm5pQI37wCPM
OrY5doPK7kq1AwvYim7gRhBjtSx2CvMwPhSctpS5cdNmxfFv3DFZlbcJM/Be
a9gvwBe9Tuv475YJkAGkvwhLbG8S9MB3/cisgT0wcq5VPkJVWPnyts8gDSFi
Y4G5k9u4wn3d6pbN2qbyLd54JOz87BwRQnG7xYoKSlX/IUl8rhnMjxrP4SW+
wdZ4LSTnNpvd3fDiy0+IhNKmHQzBDPUS7d7Tz+7hMHMy0qUZe6QV8jKMCk5O
QjxJK6pDmLbJE5deijaZqMo1yrM+w6L0JP0helKjG6XmcNCKmbMd9D0e+fLA
RO2BhRDbBCDRyYJbXGWIEGK6bK3gOwKYMbriVt3e7EOieUfzr6gBz498WZ0u
Zg6zp5YU98SFgVwDAxVUIsRTLu5Qpyt2O37c/7lyfkriPBdINnczNMwsoXKV
L4NPf8b7HRDD2zWF94NvOocqYDkxZW3o+T1gtV2FsEZtUUvvo8YHpFe5sdHt
VSwhXZTwiF3zVAXpBhpypztDmT50QxM9lOfjBY0GtSup6TdrBe8Pmsfwr512
N8uQemKqQXznKmPAs/ZitAO8B8vDYoOjVRblXTV6Fv7Gb+haxdVHncCI7GAS
o+HFF5XRAJt0LRNEcSGosCd6ZtzQp5NK7/JL+WMCh8mAqUxtHiDW3TjFMem/
h9Mv7AVhRPyJ/lMs5j5Rg7GeNQQZpi2mrNVWlgBp48KXZDpAoSQ8Be9rgDYw
SUWRGKLvy4jNi5tRH7ofTUcky3wjShE18wPKlii0z3wjae6HAUm9yzPfiZrx
Tqvq5tYilAX3O5KW6L0NyrY3oVLvY4QxWgMLufP+guJaEew0xCTF5TvQfD7C
tb6NZunC188YW7EEecvCWgOdNKfNgYvgwbDqReESSkqZO83Y+pifkBKMM/8u
tpBVbqvnC1ZkJfRXs1AsQuDIQzbwJtuXJ7FY1Zla2pWv45wOYjs7RzAG4Sfn
Cv9Cd5mj/wi8jtHsfBZJCPgaCCYeiqUJIMN10RzFEKKa12HXWCoYqNmIaWiR
0TID7kBsixSaIbVoYXabjLu1YKUiywO4tB5S9D24C0tftfEEFPJPPkBqzn6w
R5L2AHD1RDGNqI22e/s9dE3FNo/G+MZcLeop9+M9GZ9by8sggppzBPxTQoNR
czZm5EzH2EpYTc2BGdSkOAZcUErLMRpmmG3BCuuXCi7m9YGgx38njd+XdDhv
4E33zc1SmvqsjO96lGE6FRHzhr45SUT1FWuCBoq5nH/cWVjhNMNYQY8r+oCb
7NRwin0Kibr1dpJaKYUgnhxgFjXGVRkgPj9cHY6UNUQhCfibOOzcI4WwoS3V
KaHbEYpJ4jlprw7Qxm6PwtE0iyyMeKlPOTqpXEbF4Q7mIqGjeW24D0refn9w
ipgrusFRDleoGde0gYtHJcxZVEoR3Fl2oS787TYqGD4hidsxwtRGOyt3VIo1
t8/jMne6nvJn/Row4dTL6EU/k6pIS311/bXPXATMe0xToAksY9Dwd2XloxSw
BBYAJMUeewc5H3aP7Lugyc+CRAfS17GzpAyL+wuj9MrbEJkWN1gpUq/vRvFO
Ne1BFIHqb857pK5vin2F3OEuta9kO4a/490DgHkjXg17+hXnjJMOPcNV8HrK
dOQtwtM12KYVMGwSXRTeR22kXi1wg6DBgnS6QbZxAP+E7hN1P/eIc39uMgpM
Hi9Ji1LykqC5BhozK4CHvOQAxVjxPDFXxCWWntGBJUwnEyT0wx2oxnbCVFAp
8zZED2LDwzdixCVzj8DuKqGZVcaaY4cKI5hvXSQhea19WgiPPJK9+EDxKxpy
go0K9kVSSvy2SZb0J1kuLMACnvw5pv41ncVsVJ6Eh9CGjMofxG37emGZenPO
9BfJURNMdljHMOfZpResbIj/0pvyeodBDHoY1qfWKMT+Xaevj8DlKDga76rU
qd60FzWWQsbK6OK1ScNlcaP+5KOA6w0JMxWUu4GKEZrqIcjC2tYcZyaGoKiz
wdVsYv3ZcZuBb4+Ix1tjhmCKfI5D7/3DNpJN6KHrT4maOtUcAMyped2aOGGp
1aUA5H/+EvZv7GJ24h68slcTLqsrJL4Ecah/1Gk40nucvJjkJKorGpojzoDx
AJU+G9UI5f+Ugc79qXTjP9+WqtpixHx6ZVuuPaIYyCnTxvMhfr4O26ACf5i0
XGa1ywfaSEDMFQ4o2BWsEZFsCW+nLAloN47sV/SPpQZXAFHIUcVNsMyXR1XP
RgwPfZRaJ5aCG99flcNuqI3MsRKVXz5dPjMIYXoOZsKsXfkGBMkHsnB+Af7u
ixSTK120fF3sACA3Hlua+3XXyajEpwcpGzlq6vzjQXprTApcLvUaIiO9k3no
CGkj67qQZZN2T8aLirANbOuKph8Cwr6A0t9huQkURL1Wyx0Ws2PfEYL2roHw
KvD1R/UFcmr0vTI4J+whlFSrOKzP500QO0eUyV1KXLcozYMFzbEPtZS34oY1
ryVLDURmCcmWzYtj62Sb0VZ7NGn0oR9zTPpAZyltReSXoe8I8/qWijzFeCda
2jBIEs6fXjsJG/sJ591JKEH3oIWVr0iqmxZDK/oyk5G2iX0nemONipxeyt56
1ycLHEvD9ImsDhomN9aj6SihLC6uJzXITmSfA/fEEPF7WQu/gWtixPic/3Wa
q2pnKAZyMKi/BykFn0DqLpCWRH/X9jbj3JTY+lKOl2eiTzisXE+k3LZrN3Tm
plRTdOkZyYGQmGy1wQl28O4dm+1t0SPt+6W3dAlmLiIZySfPIJus78uCXhE0
houi+4RHEt3U9Y9JHymQKyY9T7rfqiKjLJvPkGagREc6YjtL6TufaanvgUQh
/L4WCGTF21RwgFtpmFuXWF/hZNxKBgiAb3qCyrX4gYYxoNfIJudscqz9a26o
tTHb/JfHUJyTzhtFuWnbmTK3ovHRZSlRMFtqwglMyu7Q6AC2v4fOyQt6H5n5
uF/IL9A/8N33EtybA2OPr2cqHtHQNQZaWyxwXhP1anImZxOi81j2CNtM7xW7
J/hK9ylFZxaO/W4Cg8FKkX8ivXW58KeZbx1SVeifBxeoMe/yXFkpFT9u/4NJ
oYqkc0uO84506L3wCtXkN68zEB1rtJBBbs8bNaJ3NSXF0O4ju9moDJPqnouD
XxqKJO6kY53TrMx86yTYIDuqM9p508MiTO/+U4XKdzKlVeyplRx4QXXkdwzJ
lU98TSvcOrgQ5Yv3unXTJOwTH1MTURGXOqmkEXbOqU5EDrjfPK2+wo6jj8SH
YFK0+X2o8il7cs85mT1U0D4g9TiAmsaxJYBYstV33il0DWPYmpyZfNq5lkBT
m2GBGdSM8x2efSwCAXd9lmhdTOUBdfQu1F7sD0vLrdbJlSGulAR7jE8kMxcJ
gPUcS6yJvYhvJ6bTgtBNKunRtsMDMrtSXohhbaXoK3LhxzT36w930MTNHyKa
9UVhF9G0RZnF3uLf2fKtLxJFdiWPQawLNMdkOXGRauWPmJKPQv99GoucSH5V
XE3S/bhryMHNlB4aawQN4DY2S1FO8nd94NhXQtif8D+E6KuiSATPtRDv053F
bZTz9WEaohgpt8q41TbcShJETiJZdswlqgbPstFReOvF4xr7JKl4xXN8at1q
S5ShGudTfRFk3WDfNVi12D2CXLsmYRGMs2l4t1F80b5L6/J6b3/8LhGBAThm
UToNA+b7JO78UPrn1JcDdt7Llq2aW1kn3VFWGk8Uu2ec3qz1r3RtttQLK768
z+KzBHbDCYAsffcQSKZbXJDTQ5W/1zVP2mtrXklff1+cvyuvezjLbPInhbuc
5lJrsBjR7J9XOYFQEPY+P/FWyXmerwQtUC9G2iyqViIyhZQw0h3qen8lhPcw
nnamshQVwwzo86nYJabQtrj2g3tEYlamqApxlikFpnyXBm9fXUTHNcE/Ev7i
dsvjmgou1Ae/KHUg5zqBNxbpydepUlcWmKZU6Rqv7OmsOg31utGrtEJo4N9V
eowMRr/6wXQiyijNVA1GnQHNGMg3EcVpHowvarIKuKk6cCUn5SnSKLNwTBIL
J5yuYU+bmvJ7QBmsNCKyyq1JD4LQe+tMpK3PDJ/I5dcP3hQP2PRtyHGGcgMN
Dd2RWdg1ilZ0ly7j8ZWKzrXgHN5JnyzUN3J3QnkedUm9QAGtbvQr9SGi5Aiu
+40nkkrUeTjprYDIigM2ci/ylVUXxivKvNtW0EyeY+JimM0Scqn0NSya4Q/U
AkI4adGKdMkSfz0ylgU2omxA3dJ2EnqugNSOPmhWO64Vf26Ei4O30arSmWnK
zquY1Zw5GnD14MVaFrhkdgI78kjJxguHXxvfsrvVc5RHqENQ7E4UaV0tYE95
I8paUvLNvC4UFEVkQugscE/z10RBly5uaTwR483yLWOq8cAAMAWJn3Wx/Pjx
mZ24t1lHn+yOlRPmp/UcVpZ1ZuDHUd+sQKAiYb2qYIj3+0AIEeY6NSilQTwR
fU6g9a5hZQPlZlfIvjDYh8C4487sRiw22dxy7egRkIWyPiqvFcAsZZ2tdNkq
Aw3FtnbVTOHTwKKnyU7QhJhesoV/VMZzodutzfJdTNTg1Pd1bzAfCwYYg0lq
aqy/e9h2OKXg3O9B4IbkH9PipJz2Rtb1gUURZtdYbuN1qthgHWbOvZUdLe4n
tarO2Cyd2Igigrg/Xg+3+FMA+k+coMihNEXi5hye+CakdbKCIPkzjo7CfsUq
pX4adYchqpaVPCEOszB3wta5HgUGVgbJeSW7DdxQgBhn+0GIo93brp9C1Qo4
qnhrR+EluuN6hzJBKuGnzvaDrb8NcNR9xq0LFQt8Ff+k9R48CD0T1c4E92hc
vLFMcBXTUj6nQdntxvdasPaHlssrSCIquiTYzbk+Bp4cAek61MxbbA2ktECQ
XlK11Qf/9C8pU3Iik6FZHGVkNX964oRCDhWXgRSPV6PE8ftiwpatzjuzHtAA
co+ma9V9wlG24Z5zv9VUzkolm2JRoXgSPUxRROLpZFs6SFOs4kyDQFuhKOdb
FbVnOdehdWqxC0F3PBDsc7rqn5OK8GuTdN32GuIB0HC4ZSSO6To/VjJK2K6x
2vTFotSytKxHdx8FOlBo3Ny1s/lLw+6YZgmQDMtdg9wcMSbrjjQ+AOfjlYvI
x9KtnE5GR6krorjWizS80Q4EwJDTbGcbxMv1x1IksA8UlW0IdPshoUBGZe6k
UHY9yiodm5XUPvUaOcrxoaLTK6lRYIHlrri6KvuEae5z/f2ZMzhyyjV6RvNy
AZ5fpSi3YMltx8fseYZ74bf2ZYkDbVmSyayJEWYtrIRG0l83RjmGn3CwtXNX
QI6usGXwu3ZReLv6341nJ0ovVlH8nSiabC8jVEZ/wIbdDcSceEWcftj2VBTw
SLQm/Uygk+ZihJbXRF8N53pMIZQXo8l0AB4IBgYPMUHOuwjuYZ4uYhvhBXX3
E/xmxqtJKcBBMNX0kMHsARPGW/eZraYvavjHsxxTGhLUTWTtUYbz57KiVjYV
G42nXTymM1wW2Ee0fILcnNUuTy5IpM03e7XfzxZGlTfTbPaVrVtBO8MgJWLU
dlNY1RqnkV9JRVI/iqbddh/kwvAGaKY8DFmKlFKRCY9GPgTZAAg8sdyDI9+Z
W0EKje2jXhPVSd6XJZaEFlvWlm+cqZelWIZJj5HKTvGaSmSYj7Tum0Zo40QH
y3FoLcCIsQf+KnLyre2Ours4/EJHdU9khC0kWpBud3KMwlJpb8BW2+r6hiry
d0q7fybRboYKpGLgbgm0GfPEwWnaA/mey03iYb5wFwKqXtucERjtw1dcCbxm
cpZ9agoBnnfkgphNGAjPBqCgnr+3poQnINO8fwQR7OCnEzHm4iHGvXszwNLb
PnVF+cMPeEOnT9pe70k8zUi6I14SO0YCRsgTwqwpO6QWnQFn9FNCqaCh5F30
Jf/JFkQf4x3BPqlc5I8UezYd6Wo16fHSbGG9Gs9cmzTIbLLaHkU81DRb0gKN
bFxxQLJ9x4Ee5//61iy32B9oQMzsieSC+QDcy0MCLDb0g3+Tu+B7OgGh7gwk
o408km4J5cs15uqRBDkHSPvTusD2ctWyrMFciMsRIDhltSgRJaAF+MK+3a69
jWUaXNEW6xbRDj2m/m59kXt6mTiLQD4hSuPbqMFbzJexY6v3b1IrKrUPiM1+
dW9FX9jKu2d1vBfOhIoxUH17CS+HUff2fnD808n9h3PfZj3QZz3dJRU2FMxy
Dp0k1W1oXi5Ujrhb6bhDhx/530Z1lKOOv4e9zc6PcvYsVjr0QkdRJVIMAAZg
Lrnf1u7hXfd7FGU1pv/9IltufbeKqeH+F9Z0SWK4sS59PzzqgpsgKPbiAjDi
R9dRoPeZq8ddNiW4wKdsBm9DNAom077tkApVwlNQB0LxeumIQKem1YUyg5NZ
t4QuJ7QWjFn4o854ahNhnaMz8vLMEi1btPwgUvIWpphw4M1XhgtUib1COQol
7Fd7YwnmDCyG/Jk7XxtCiY8pfsMoVqleQjxXzmVXsNpf97frKRrWnAqKUTR0
i6NMRYMKMcyQHESdDKhYCAsCuebGP3ewuiBH97etab7zf9hlOvg3F7tm+1IA
khMWO37AH6Y9+KqWlWFUOmPW4Yv3TflxFV2eqt+oj41eIF2J9AIazr//1n8H
IrFRrLD2F7eXhQINq5wSQq8+gBH1YarnUj0psKDpyaObR346sdxIjy1jxABw
p71bTTru68FvoMBQwMqswjBCcoUbOJYJ0FGwZC8rkCH8V5sdcENXhQsX0Sf0
WHbnI3VV/T5vmW+8HJ6ZkA4pYMOUecqXTXDHQl8XGvJMxl9b00R7wCfVp28m
c/MtahmNfg9T+DCAUu4fI/Tkx/HTI8dH4aMKbK/8XOgjLKhz/9kyebZ7RnvP
ylcvbh2JLAFgLLBhetSGkQgxMjSciFlUBFQrwkCegsI/M4vHONX2WPdnyRCC
G0xU2kaH6TtaBe80Bq/5A6yMTPdFGkgWT9XYiY/CVJFx41+w/99GaKmQTBHr
tUWPH0OiDwk/mbPgDQUA/qmcgTTbQhfmI0xD+F8ib+jb6Q86j5vyDvBCKQ1f
YDLsclN3XIGGUq2OFd4tU+m45arAX5odOrjE60ggny4QaIO6YxdpuMivx4FD
SbgZV48b4GBFtah0srdmEeo71RjMKmv4bpyhxJ5vgHx3a4BNPOTQGBghDJpB
ldg0MMe3LGe3vvoTdG2GvJoLAwL9EBWev7tYWaV66kTSZ3hqcJvqZtaSQerx
NfyzJZQqvOTN9/DN5o7PKScW6BQEN7ZmMkUsfNVShS7U2A22vEBB91ICHzai
rtHdoldVP20lZITeDMMIJUESiNZKdF3h7mKiqP0FgXaj5rN/lp0DqBTSjWlN
kCYNQ6BK/lpTopnKLzLiRO0FJWB31aQxmPduWrfWFLTl3vOWFxKPuLRLIdJD
wwGKKnNYitYPx6iSzHue9V4OIom0mb2thye9ynyXi7cqcz8kSM8/hJbS3vgy
pvhWNd3HgLjrxoNbMbQDZCQufrkelsNnuu9LukqZDOhKBlS6bsrJiaFBUXm0
oVA11I3bfR/J+dfz2fiZVsolM1DF0n/zeCYGcC9MRU7OBSaNzqJyYnDShb/h
eASbHo4piAku29dGKlApw3CwCOtBe3Jn5ZpL+kvdB8mD67XG2Kn1s2h+ESz+
dPB6q+5YaEErD/k90T82oYfnQnbtLxVvTrEmLuqVCUqSv3u3z/rt7ePpuk/4
LAtF8ObK1sDC4DiN/AqMu4C6aW6Cv3Ub7jkTmVuUhipKxOEN3MTtyaEY2cQc
jOIb6dzGlCW8+4DuVedE+5XEvDjB4YKXoPm9FyqBmc9iuN/HrcvtJ/975EtL
/7AyJytA/AdSw4ESDrvWYN8aLbhExmrWI/TJ+InOUuHB2Y9IvW0iYGawvRE/
qFThk7D2yV0SQiMe3kGxy9L36X5T3F62cQIRxFzyJfIRhZFlmiX16emEFC6q
xSYyUMD3CNlenu+6+zPT/ddtdu4kibrrZNdKJkKnQ1JPQaiT5QMQW9iOhnZ+
QmffTjFo5494iy+dI4RwnHrTAuScyme2gGapWS1WqDY9FyS5njawfODt8XuD
D/MCbVSFNGVx13DFQiZOJdb+ggyFVfxF4bY2jHaZbEfSTMXGU2Kztg+LgGyS
vaLKZ7Wr6d+PypBPmlC7DjZLF7Mlqg6XTB1xLcal0uLrDEYqt+HJ4cerNOzi
pxqAKKI8aUngHCcZxfUE17ASZ9hOs0seU2+6bobWQWFTv/8zObTYUpJsQ/P/
MBRRgS2R/m9tYy3k748xbca7l/lnCVnSIpLYCXmLLjvQ/eKVzekSP7SzNlYk
YhBe6iKguk2eENHw1HNXOSmhta17sgP9I2nFFWbSQHfUTK9dj25Aea5XAKgV
zyfn79+reiCGLVj4rEMT3g4a+nGwZpcmuPx0bblhQAKGJHBTl0bxHAT7Zpqk
Gjz+/8MCQASig2u2Hni2Q9VknI2iCLZTTQfLLcIi6s8bRAqE6rzdqdwWpdnh
wC7ZdbwPPDZAVQWRCXJC921KOrahosqc59XyF8l86quICvOmJpEqrjADZN8a
FaGafW7dtR8llkBgtM4RJNKOSWVPm7CiVdvdwrWxN6t/Nqlp8mFt9kLQbWAu
ivXmyY0wn9c+Pz3Jpmj6lfZGEOjyaLIZd4Wy/g5AUI8S5wZpXqqPSpYpXVFN
2WQp5kfu/Z+06ko2wQovxOTx8SjwAtOg4GJ84pbYp2d71fGi1ealY1V/KZL2
4Qun/i6XvHf1b+F54EfJ6aWdK155FDChI8v5Yr8cyK8Otfij5OYWyTtJXCKj
2CyaIZrOQQs6ug5JGf0XtOMNt2lGHXBGhoY/SApLpjV+ESxXNuw/HWDrnnEV
DyaJypb5q4jTFfyQA6VenBMoppj+jPun415W7eWY4wMgJ2aSTsPaK9dBLVgx
t/kXJPxLiaTEmIBjw5jcUodSNc/0nZt5bKL/KFiyCZ+8cSFHW6VksTtsyogt
GmFefGoFQ9ULLDRPnWMscVLzfvV2T9BTVLTM4oRhwz8aBr274KzsM3QPi6KV
zAmjG9GV0i4lldAQDQNb3b3CYu3wquYB+AKZWWSMFzXF2ank2RsSgtNyvDHG
vF/wEq2nlTuEPFn7iCYzeeHYPwgzxN+QUhbPkIzNLH2TF3R8c2RVX6JQxwkj
fxUMVUZP9E8JkH3j4NDD2LY7v8YkUdgjN4VadXoH6nbTWd/0VQKdh4XCA2zk
paFpQlpTu0HqrsEjCg5ct32oTf4kRiy2RbYcafirSrvvj1CpB3A1svyucBcL
mCvQFqofCMpqKD7S9WZPvm1wnOpg1OQLyecrceOB80VI2yt19gh45PU2zzW6
HO6KEb4FesZIB8mUYhgNWk3MiAJgo7Npif0ddvJb3zLHAUJYguEJDIvkwudr
d9ObPM1iAGbvoe7gswn93DIKvrYATuxLEVwx6Qg/l8RUdlFF5Tqm9BXFfcnv
iPsiScc1nP/1kwRNqKQhCgFAqAGTyka1os6MIiTlqkANjH5EazPFk1n90iKW
bBKOaxDT9fDK85jthPcG2SQ60C1qStvby1wyRWHSKBnrc9epvnX9rgiAYETD
MQMuM2WXGvrm5pYUXX+3Y1vr1xRfQgl8b5PEa7JJfFsk+LLylB5DmsrM4kKm
+0i6ino9tgMzRnK77TJ7SWMurDGobQph5M5q9mYug7dUS4FLyVAiK668WLj3
YRdl9H7P6+LT1bqeCBnXPvT+TUXjODRQ5XP2Tkeog6Ckqn+hT/oa0rgWeJE+
aSVfmb/DfW19u6O0JacPhMDMhbbfKujgSKGtQPOBpBXgRtZvboOLZvt3NnTr
LDJVLkMcz6K+tr3Th2/YMMgwFi6g33wNYIdYw7MdgbxK/5aloXOje/jjZYtd
96HHY70+zbEiz4ndhiykR+X+//pR3iJQahxljFmjcmWoWNreA8Hgfwss57fO
OBpkRpI5n7qG4f4yGgFFquXWDSME0lDZfPY5IJUVyDNqLFa+8kuqq8qdImis
IttRVK1TaQKk7zQOfUuWoEFD5lV4n/6Uaa9xTu6ubkcFpdxq1rkL2MUMiQ7q
ElD/5ZbhSPMgfPrqLYJrTYpzisF8bovAs2tFic1S2V+qtu9je6jNGOf2uACy
sHfS+FOnORCuA0lCi+lAhUCStGm8iywpeoSeCOzwIm7QY6ZgJUGwKyylO77D
rwRMr2R9/Ix0R10lHqLIY52GPNcXpyOotjAjqfeG3iD+ChbBXT17SJn0w+n8
MPp6f2yTFQwiQHBCiph+AdiCfWlcLj0CGvQeytaWdEkO6cnlIHcSMLa+HzPZ
Xvx62IyWgLMP3MZ3SggxgjGW0Zuu2cy57ryIwNdw6Rt+xEdYDpoG+hfxofE5
w+5vToeB/KbEeOor08WekDt+MLm8lU7sk6KfPR+wVwdaoRtVMwKwMeKa1vmr
7Jq1aobFtGDrM4AzFhVOjIvNAxgfIsZb0GGZjoIOkeKwyMMw15V+RQLQn5/V
KoCC2NZhH6iqWpXFDlpAFX3MtvrUXpDeD8jh+LZgbpXlsjBV2TP3iVCQDY2o
cQXKbR9h2NxTX/4x1vzdMZe6aorPOFoaEpsyit9Js9+lirAZbkUVbCilVhTj
LzgJPoYOg2EtGN1A67t1A+GQTWscBAIdlLMIn92WRAcgvSk3r9NM1K+8aV+7
xBgRHR/Udq6ni9RJLggi6dh6/qurhHT3BxcmHMPWRcipHsNJuofWeg2zw353
9hR8qOfmrJtMBZJG6l81zky3U3DNSbzTUHghlglXryRhE28QNpeOC4WxnqjZ
nAzirSnpYdy3B6pK0KEd5+h7GddjhRmTOYt9nU10GgqpFRT1yEnw6dWktqy5
XM++UZSqYeG1KTsuPhIq5FjMJtxHR0aeww7BwBiDNnwHNupC5hcktMiHClzn
sh6uSykzVSxHuo9vcTLy3+IV+g5/ABdEWWuELWZtgAeoY+g/bIKaZjJlyibL
LVisCRN9lKtHTePAM3BUkWMHqddaNh5nt+DsqHwTX635NAZxB7IGMqmNDpmc
A3F7b2mTHy+YX82VMXT3He6GDVjK1Qtja1Vipv7oZraxMv3R4zsET/pPyZWz
HCv8XC6ApFRTrO+CXVnWKyEzJwj41NpkscIAgnzZnGhmeSdZRzKxxMiimxAJ
gO/psWOGSsyn3z8P3Zbrwu8y0gfV74SkTpJoHT5Td9nAfH9D+n2B0tkiink4
ndNHJT+SYt9RixQaFVuCPVkUEka2dQ2Q+UgW0W0Amp9k/GdTk5aoYwqj4SoB
Q9M+966mJk49gXIWjWQfWjRiwAdQeEPq++w1Wp8g1OMsjJ8OFhR3EmQeq2Dl
aGu3KSLJgOJHC90VrwZyXmnMAegi6MizEPWJqy4CwHvfb4/o9vnY3Q+tB//f
juP8Icg41DLs9yiq4Afv5DLJVVqSNOitRb/df/kef4oGBB+TyBvLPdaYN80C
u/Rd/yqKUGSMXBJipOe6hY9gyB9/Yf8kZpUfMSDy93enB/8Q65x9ey1BVyMH
w4XhyQ8dJbwOvxNsnlLxAbSNwRIDmRDdbko/FVwoBTn7/RRzZmX/n8NNwN8j
ZQ+ScRhECY8vTu2FybwEFyKgHILgTjtJPgANFwoR4251vaGLugEaPn50Ty2S
jdPlcJwfSqiUcl1LwYh1zHLFkYAJvJHyqaWvfzvze6OmJqwa82yI2JZnlTum
P+QqTwzjtIjMsYFftf4Wnle3jdaEGpbBRV+G9rD1Zr06zM+ToHA+CYMP+f13
teB5JhcXTi/iR17Z1YYsIBUHjIGOYe35L8Z8BaHA1RClnnanjwUUFoUCxIQW
KjEFOBn0hrZHTa6S6pHTn/DCQiJdnk4s9pWJkiUnO3HI7E8Lc6O2UF/8kjLm
Sws4+Pb5xwnTuE1ZU0IvFU/PNJHv1hn8qqpwZF7yCJav1eTOXNMZNBUV7B8o
ho0o29xGMY67sN9LikiUN1Asy/ZOjWjF9f6+E4j2SGcvEQRxX09yOT0Vy0pr
EEQ1h3il970BNRaMwvggTXyesNsauxC1T0Nh2xM88V/HIUSA744LnZz+vs5O
rnDpr71okj2aS4/xOGE2yidkbfK2RY+vTu0TJeGYG7UfnX7c4WHZb9bsWmUH
5FHBIigqJs6ZmA9up5WY9UK0OPmONgMrulEv1+t/acT/otpiorS8qhJa92Pn
6OthwF4Zc7ZgDXmKuiyb2mpSYXvzMh+Kc57/w0w9PLPNRpjxNhfXFBV/mtAU
yVtMmyG29dczFdNbec98gtM6NYbUNTn8GJL0/G+y8vA4uleqKxM8fRWf9GA5
V6qvOqv88lqPDVuwBgew7RpqrT1oWA8tSPHeiaqgprX2zU03fHbZKb7bT4JF
nkJU+ORX4a3T6sQGIWlR5HFnXMc8dqwt83LJVAu9iuB9rYct0DYP1/qomTwO
V+6aG8cqcK4nzwVsxFeAap9OCSc2WLJbyqAz73ceG7IWDfd5tY+BxZhLM8Gg
lpeoBP7whIcsEOyz47IFGHeunapYmD9hoTTFan7Pv1odWmuG7PqqFYEg593c
2aIiqAcgvTDG0vSN33+QRpRHMD8YiALLM/uAXNFNDbjMoPh/5Z/O7kYDnU4L
KPGFKsieuYdlyfmx37vpPVyRNLoGIOnyU8VKcEVbOI1zSQROLhdL9VvdlGFf
ytSS+YJw4ohQxwxr7l9zymZ0xq2bGvnYK8bVLrcAbERFic7jaQzZhWKcZzTi
7jOk05yY5e6DyJtxg78vh4IDVTv0QAJLoufpu7uXHWKwpXb9BXcQMT/8oNe0
VjkUJZPudUBjnZSjILfmqqJQGr+UywYKpx0yl9oXpPX25mNpgvfx+HUakfVk
OAE8RAVtRAZvH1jVY0289pZQ5L6fnsuiSXVwKisLoMxyeTHKqXIt8kMR3uNn
KevAuLINwULpjeopShQoWxn5c8NMX1/ApvYsMHv5Td4DoU/C9E3S/FYYwcVR
oxgi8hlA4eoKG5J0rU74YxilEd3a1dwcNUFedZR5pQAFRNjIr0VSW42ik12k
HZ4a7t7Rjp+Gxg+7wzg7KJqqwqrXTW1SNtmDbNg2KQj2urmCIsKupeOBFRkX
JEyDUi4DbFpRuVlSp5mZKLPmT+icXR6CTFrY4PR/2KViTPfNF1H3LK1pXQHK
hkI4fef89oToGYwnSSN3ndWlhUSUg3xO/q68j5Fc0oZEiTKeHmbZ35UZW/UI
FIF7kEdv6c4s3co9VsfqpjbTiCcBc1i9TcBr83YTcCFKcGB+l+l1oDmvLto4
BbcywRXUxxFYgbSR6QZLFcUb9cXSaxzyQtFXKlsYpvvfJCLBDq/nuLqhnYHe
zRt3rDyT9/afefOHAtOlEi/8AMZvj2mG3hYKfIgdkY17jyWX61l3UxmayvAF
AuVnnc8KuPpTpeIkqzmIU2if5QP/hv90wv+rnLWUhkQiMe15Qi4ilQaK9MR2
Zvy1P2a47buqz45QGpGg5UEh6Lj/U0W7PHNjdWLozn9/hSeA/b8oBHLOWbz0
0dJTAVUxmpwKHsG1xISMnjdzf465sileLIbr2tkRL2LY8v+zREN77sNUhvgx
6Us3GX2Y0OjJ2Of16KFtndDADGRRza5moBW0iMr8bGdjXQG+SpsWVBJfMle4
l3J3IQ==

`pragma protect end_protected
