// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pKxXnROdQOaAUu6QZ/FQwHTDrfj4dh0MQv1GARLbWgwEl1erRZHF1hY5lcIY
euKzizpuLF7nh1Z2K0ZNisAjT0eFSMoj9a6YZVtRlYWOpgOFo/ILk9jKyPMm
5YMd5uIUrG+iO7NUmDdOOj/BvOfUtIbO2WtLLscOIKK/ygl/IbCiS8ogurNQ
0GxYKRw72xhMeOP1khHV5Qrj3VtHNaA9ge5lAreCtnP7xnJGa1ApEmEgCa4D
MEglM39YTCKMM58HWJOEVE+kd5a8DucjTX86xNEV7vkAqMTNMwUQIZGdtOnf
WrXzeo5gPfuub6UlNElsx+pCW6kGhRP+mcDFW7o5qA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Q1zSTk1rQAlJjV1xYMN/k8pRsCevpFQSxUglMVZBooGyEX5asKX2i/sArsFa
KJ9e0Wuzg1oOznpuOrF5wCMvyYVGCV7hXWVKa/14y00VBQpf8QWhaiqxVMqD
AMQOO12Pc7viLu0A/k9VUsAmxkqniBvfUfvXeFlz8loXKVmrGSwmjuwVwQ3M
6FwmQLlqvjNZHGtCQolrC8xed/VquAmts6SiDyBSvm7CF8XP7K8A9ZOziYeC
p3OSertKX8UQ5HumraIWIcjwvEbyJL0WhxWvloLozluBmUta7C00+vzDs9D8
g4hnMEYYwhLxDJy3BI+TJ0bN6rDwig7RJE2ijYla7Q==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
rjxl1QHDYWkRF1PvQHuFkYu7F25UT3E5gWxADGVGvl7NLmH1m/gOya3mbIN+
IXcRGH04aGjQFs/fZoRSFFfI2WKyjIsUr6S8IsgISo+65MWz8mJ26xfTUJGC
o7mEoluyJZMiKpY3eM/Cga5F64evfrx0OSBtpSBDHgpNknePuh1n6VVD8dFs
xiCO0Rf4ulfI2IslbHteRHyHXj7OI41D75dTx31fhCpRZ1axCAs+lVZO2kwq
AuDxlGFgwvCVA9sYazHURaIZzIkbkIB8leWeM5hxg6RPTkZVnYbI/YjNAr0L
vDK/JzfaUHmApdjtofu/ntA7Y5f0+JpQ0fz+i6EuXA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
VHXc7nCE/GwaxR10G1YfngkiuZpmJF9hNlWI+Nk+NbKR5BE3mn1MOsjeZgyN
GNaXBOeetPFZSmEk2E/mBnznvFiTKUzDicjyaSmrWZDANi7oEYFMBXOmDqU4
NzhJHtFHpJ0NdFKjfZRPk+L+CBLcjDH4hbVs9K0kQDbFHCYmLsA=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
luiS3w6puMPMvrJ4eOvOi6jt7p/BAplZ1WLc4CDqOj+BHy1Tsa3tWGf5AhHC
5mPgWTuQvpPJohgG95Nge7ZBpCfGEtWNCyvSK5R2meZZhx0Cm+sfP6GDwU0n
EPLa8/77lJmEeMuZlHQtSDYPmDvyKaVPLagOTVieIximbswIlmCtO5Id8aDw
9cIkHSbQ6V6HQNw8z1KqBnRKMA8rZfI881V5rcU2toVxRSeZO1nMNlPD64K2
z1bXUjeXZZeWQxCAMJbRq1EHVK7eSmHixNwZwczazV1uFxt6jxigU9eOb/To
H6NiKtUGJx6+JiNd3r43OFruL5GIlPkbDdB2aGzwuD/odrqevtHW0P2rYNbo
fkHoyMv/rQz3EjZ6vp80OEzSy1SoUe39aOPVZgDITPhoESPVmutS8IEKSA09
QwSdUPa9Jzs2uwfTZpU+5kidID1dIsGtzkjLVrVk5Ry+7c4ekfy9QsCQm1EW
S15aw9bwwTB5zTHJVqqN3lSVySDK3fgR


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
OjnYSjOg2KdffaxtUrMuX1IWRPiUjMVONJKjhIwvbNhXVzG+tLEzErkBSDX+
QQsdscc+LeQoJnTf8BRSzwgEL0dqPPBYD2dHfmEOv1J/dLBb8Xwfk2mdeubR
j09xF56tULaRt+t6pRh1AI8bfqb60GdAwPC3FI4j2Hmyks7jlsE=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Wj/F0tmAO64TCnmrzLyHvg48+3w6LCw3fq8yHksa0iqPdxDfDZkfzU3coZae
l7apSwBOoDhVICk2q39z7Lsdm8IYWtr8kWPv+fvB3nBeHSeFt4IiPIJ2loQf
Y/hANdnk2oMsIM85X2rSbULMWY9GS/W4ifus4htHU9HFXE9t7Jo=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 2784)
`pragma protect data_block
IbmJ1C92oIWWd3/qp+97J6Y4J6HK024D4/27Q5UKZMdgxnVoqUkbXxVCkbIP
k5seaW8LJbNDHQ0Ghs2pq56anLHtAV1rptq+GnO9j4RvRXZif9xaY3vOnSnf
Thczy34v6OhmoxR4BN+BM9ea3DOY9C0hKgDPoqbyjqAUUa1Zzb+rjmIqaC9Z
j2Qnh/4N9L0SGXYTtjEUn6kkPsqHzJ/GUhsQKAxSaXYVtTJgnrlBc8KaoBic
9zo+gXNuta1IP+g9M8Uy1bL82OHDOs4NCOPV/KO4n61cFzsfLN19kw0MSpHl
3//wGO47MTUyZZwz7NVBJpJhGQsc4xzx+4htzDVQvvHXqFKsI/FJly1mIPOm
1rSK9x3gl0kmoZvz8YT+GW0P+WXh3lOYCFQpvP/DHiFFiSo+aZALfwzxEg1U
gCTMYG6/EuzPUZTNUIWJtQwSCoG3UORRtqxuKP+RKDozUevjUE5xDjDdjbyK
uj1n4MIY5lAycrYVaIzZHbJd/kURr+2FdczoS3fKb7I3z/Iw00UUQDOuLdLy
kLEvvxT4P/XVwlNg//vuhdxE1nnQYItWOpF5MlBHaxrLu2OKDdmG9dBDdwHt
lHaN4kn9H3Xw78FSBFm3t522J6Fy+/a5V0mNAiqmKlvaXGro8aCYuJhHS5UI
iFsxKIp6ie2Wv6h6goltGGzcOugWsf93Jby2Pt5c75M4mqPFeAJXy9kvHVmk
q9t07nLwJ3dSyeMA444inGVaM0HtmzV5h1iTnyxVU3yb+Sci+IFXaGCRsGnP
mKVPGNJYUSTQTO9N+ULicKR43Fo43Ataj63nUUOVY7m/rql/LSjbm2MaatuO
T4AcTH55s5BFbpdGOSqCUvWCz0gyGR8kONTuWA8wZ2EMSgq4+maamGByPICO
z0jvg9xzYcF7+2kKYz/zKLL8XZZutOvcMIO/A0PAAJAbSbGKjzh1UG+kK2ja
l4QsJeEEa2kQGOK17icMv3YB3MwDT7a7HGXXhR93nzsV6HajmnCgkl21oXi5
AK+V3HdZLDkZ4v/WlP0sSDhB9JyxXk1BKfDlR6drShwN//1ydUkjPIz4kvVW
OXVen76XcNZxSEtdLKlwKMeJek8TQETAPeOSDj71WfWQGHgcgkYsTRR9NyXR
0lLQgfYXqbyWuUAQ5sb37+cBVfwqtEMLeBt+hStfDsOVmIvF5Gd5r6epwguL
CTHrpKXLtb4jujVefazfUsgMOOz6az/HVy+H+oc3pxqi0Ov7xstHnsFb8q9g
nALt3ygx/JwmgOFObiOITp5TqkK/ssVY7fRbwraLhTaH6XAybHoAUGtS2FFU
CRQ5ayepWih1CVZbEdmhGVtsVQTg+Q8zWWGqdXYBKzaZ0E4pGL20lTopQgPQ
ym2NZC6I/eLeUypSROu8+yiC0jJ+rcBYcaXaHfh7iTWcSOBEEGJSS3G8OyEA
0ZIKLaARAH7+JVlVp0A7dLD9QbTT/y12JVk+DEmF+mJMcRyhF0Pyl1RrPSGi
wWNw5SYi4bcwBt8E0zLVTemhgQ/fTEdrISqrs0LPAz5qI5fJVdDdFOuKQMru
PgMEMqYOFsz9+uMpFPkFcO9ed8v3vGL/1FuEaXwj4daJUxuvBFo3FVu+isV1
fSuTU8/6wHmb+CRfo8mI7Ze2tOn+nfsF2TLQbzoAGAq9/12K0wKyXt5J3aq/
XSPaRvGh++i1ytoY+G3PdWuf8lhNS+z/SqqAAgbHmJTJsj1ElAU8TOquEjUy
g6cGI0sLZSizDNRVKVs/bkaI0x1uqO5BQUv7V/SFII/T1ZQ7FgF95zVnCR5L
v/1k/sbtoR16KPsb3NeoH91eM1DMNtaA5Fcm2P9b2lrLilpWcsxejRU/SErp
KB1oP6oCfrG4E8oYxUdmwKtx1HJPyi/Kh0BvR4xwGYSLXCgJKaK6npsAXB59
mQfaRCKBtiJAnzlWIzR8JsKsyCuf9XMUN4/y0tqlYWFhWSQw9bb8TO9NjBKU
a3nLsdboebvTB4B7sOwHkpLK9ZEAhuXscjH4eM2dJ5UVhH9UVEEYcqnLDa86
rBkkZjWBx+WiNMBBDwNrnfTPeV0k9nsdgDKAhXiWhWgqjkql7AD4BAxLA5Lq
ADVfS7KmNWk2p+7T9x+fPdEosVzitZnZe5SKpQ89Q93tmYQMxv8B1iY9PqAq
QvcOCYsr2Pwgdmgn2Tkl070wDW84wa2iw+td3AIXcEQWaKhvMUx7v4Ey4Vfm
vdu62rmqfNZTBheUjumTKZIY1Hj+mRCEk1R39deSCGa+iiV9/NS7vuT4U1K/
xH3+FJDYHcyxrNqA7o47dwWKO1dpyZ3OXpI0PdLvTJXrS7PLgJdLVz7noUS9
PhiJFqQrufVbzleIF0wZ178j3A0p6qiJyHKfQpT/etuvL+a4QZVc6zHeesh4
1nHTP7/DVLrpFegV6GJp/PzQOGE2JtH4b0ANhSTqqiKh5sJYRIee35szJXZf
nwhyUT8Iog+JRpd7ZUvfQm8CF15BjZSDZkIGZp8SWYtvlIAXyqTKlJqyUuF1
ENUJwsSeu9tX0Rm63wz9k/nH4LX1s5yL6X/PRqviwe6SWEeU7glR/oPhFvWs
7PXf2zDb8HS1TE0dKKRRVvUB9uRvIw/39FB8oD8eckBC1GXu+dt5Ye30TyT+
xgSPueO04Ps9pp3YPyHf9h/CxhcNGDCrPn/z8jvT14hKmpB42/xib2AHRTMQ
jtH7/U+ApuDSFR4sfezkrm/xnm+jsXdQk1Csd376TLOrKaOJvquFakJuIwXL
Xu1nD4lx5o1BSXR60KH1Etsyevf4PBh+ox8CMdG2yOQQOKVjo2oEbwqaO6PN
ORtMteosEfJ3e0vaydRpppB/79BKbP09rjTyPGG6JI5FTNzZsDpNtwx+nJu0
FxN1Q/3MqGEje5E20mJNPC6VYGpI201GVzYz3Bq1bJ4DForW1N/NAvWU05GK
TlZL8fNtgtCdF8WnsXlAjCt5a91XBBxYMmX2u+F6PVQQ1N7k48Fcj4nWX378
z15qCRN+0a0PKGyZe0i8+FyC29vZ3RDMXXzIRxHIok/5kQpeoWC+thD4suZF
axPgUIl/CqcxJnM97QyUbcjo0KZc8gYs8M3MN3EUOrKSzl+SVY/QF+HCVomr
SY+ZNnORjJhNflSWyGIH5lFaqDLHDui7aztO1ni2ka7iisW/UEYcH1UdukD+
/ot+IYtlcivEVqsndukqgCNAm+3fIfqMjo4vSLJTvPQjgD4YBcQp7k5dkPI5
/vIOKvXZqiasw3zOssXdwp+BVgX4oO1ZgALBJnlo1CYi3eubxi3VDZIVfC89
T8b63Bvwk42NPSfYnODvnyAbKLkVR0M9B/rgoCVJ/++FzMxXKhZTxjT29Ua5
VG8rYjsolFDS92IeZNxZiE9XWIYjjy9meOI4Wj3bh1G0hXuJnN3aJIbvf6CX
u8vQ02/e2FyiszLGLSep/jmkZZ6sNBY6Vp0cE2ugDKZszFI/MtqDHAWJuRWq
KCPyI3mg5VOzwnOpKX29EJ9XiyGEUO/YIjn+myxzSh1icAeukmVfw7Pft3IJ
quFc+amNDogy7Y78nkZVHyrxvlL3XMpGUpkoqVkZbj2ORq29tcIIapPfq8kN
wECOTaxbWArOWNv2osBKF2161B0i6VM4rG9Htqja+0VT0LDb3a3cCRz2t4Io
e9ffK2jwiyaRfp6gCyPSpIwfiMRPYY8nTp8D6muETlQ8y6DwbD1D

`pragma protect end_protected
