// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
vEXonWzNm3ugkF632H0gRvWtw4w6xLMAGZJAmBfXDtNWskGBqQJYdBXXrP8ANzSf
dnPsjVZKn8Mqds0n0UFfjYfK6jV4wteBg9LoJEikqUSDD7dkhz5G/s4GVvzspGqq
ii3KlyER4AEECbng2mjohBSrP/vZkjgKwu05YuCI+co=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 38896 )
`pragma protect data_block
sQWtyCa8AViGz2DrRapk0TSTXqybYofdYrBjqIiFrl4b+TfH0inOt8BSeHP4iO8z
YHcAA6zY0aJa26iVDmfhNEIUr2wm0+Gf6A5UKiDbp00vKPhXhgl6KJVhO/WsxOmZ
8szfcMHhpS6fUZ8RluLWgJPEkH1d2WNPMyuA+kvwMbSeZlh8yr9/UC9I7Q3eKXk6
ooBtTxlN78bq3UQcUZPUwz3rcwgQ+5BdiFTx2A42bxptuwyxPbsKbvfs5SjqCSSO
CU5APzkx9ARKZgNff6vjDXgQU1THhEKYRLsoM8C1/UJJMOsya4JusSM47aJW3CCl
hlZ+tQ2IXuWiEN0m4O24IR2VlHhdRDr41qwz4JV+GW8EtV+c0jEPX/vyDHhHlfaG
OCkGw7w9IT1TReub/a/9YYFX3eGX8xuKfv1/cVU1x1f4X4BuVn/NKgngUiMMIo/8
unA7z2JKugNhBcVYxHaWnVYQUCG+Dkxf3XpWLd443Q8Y+0p5gESFgAwwJggrt254
VtRVQk+q/fJ4Dbs2ydVFpzGvsvJnCufJEQCnzTEbpNUIJuJWOCCL9e6TtOlScf12
Cgf5DfzZTS/abC8aDfbRGsESBsb9Kd84pFvAAEYw5FNWRs9Dp3ZKTbeJb+3pv/ER
ojR5cFBZlIJH3m9Gq/jxB3KTpnW9SB7rzZFsOIqnPWO1sZDIUocxXeCKRtWOQAiD
1U/2IbBf8brJQ03oQDYw3FVSOa4/yA7SzPRoEHstUQ3g8jJP5dCajDKXYuLv2QeH
+AiXC+eAhlKCoCeoSw5aotu5uc9O8u/BK1NG0taMiFBMElR8i7Qf0qjCqloQxzlI
QbAolql03kOj+LDD72mwP8N2h0aIaimn4YRJbstMkPnZ2RAJlsnzfsTgAfkrHfQB
O0kIKNK3lrAQVQV4o8R98WuO0N00leV8BtK6ijsMeUaoQfDeregp4+Gf6rdpQKuI
2u/YKW3zXEbUXSKiCBoYLP/N9f+H+U3EBXdZqC01JvMn0vIFKyyB3Zi72BSLylzv
5xxB857W6I0vtvhCfmV67JdQXGbPga+dttkcxjQHl/mkSsrP6PukwpBKbHnIhih7
spWzSOswG2wKQpZ/kJnQBxFWc6I4P+KlK9lQmueGPEHk6CD5lFeK7VwmydX4Erw3
gzLJOdNYiWsBcz6MDyY1ZuDkz09b7MCo48tBHHXPNOUi06UTTXlsfs8zYoYSN6AO
f/1xXwUv7GwzfmEt5AfnmEwEoxd8OaVLwP681q8EOJol2s0fmU01tkCUQ/C2wW4K
7FC+Sr7WwXLNuDpNCl88O7tOo6Us33QTMebbNyjyxkTp/7KRRaAjf8LBAX6+ltZ0
fh7z8pPFlRG6cONcHk9Ph83uwviRFoyNdDhkfTmCoFkqEG5ceY5xl9W+UdJ9kOiM
MpheedVHHCWe0Tfa6TYZJRTq98Uva8CcJLL3dhdWSNJ5LKtoKwPtF7QCzJVz19WJ
Afx/HNb/XZg7D36R820VNDPW080/QoFbAHGxcz9+KH5X50MqSgQempUNl094uEWy
sQ1Iaod34qyrDvN/IU8v9PJLx8HUhfW+7kRD4LTu4uXq62x/V4cmMoyd3dWROVXz
g1jyeqnO54qdGnHPsxjRj+TvUpYnJOyeUvtN/5mkAE8YQ1IkqCEVaHuL1BA41YF/
/8OL8bcWsGSvTrhyD7Rg82MKoFq6bTbuc+UxhrlRL53X9wXAZQhWneHtHE7y0ktd
RsQ6gdTF/NCa+CucfnVKLpx8cTlqShvX4VdaDLA0P9+ZBLA1w6EdafZSVAmixXes
8uhTU1qfC57mEvYdoucuGB/pb0JqQAZK0SmDL78jzJVdkAbTTanhvjMCGIJUR1jR
IdqXRSSVeokvAsPCLn7V8fBXY2zh5HH13XMhp2wJ7rWWWY6EFBjIOI7ZqvtMUdfm
Wk4hSYBmv5WjeCOOXyYemPP+iflcllkSTa3j8OSj/Z8lr8OJeCROkCCMGpBZWXj+
XAJ/PV6aQM311yLHrk4SL5+87dCfqdvWGCMeWU0BjlZsyo7ACt56LMcEbSMD0L7u
CeCce2muYZ/gd5p6Em/Md8xSgAlkMJQfB61XbslAFFu17JS3JvMk0t769qsA3gkU
ZpBykhv77/5j8hnHk9oeE+38bgVLya2F1flf63pDHIO5nREWmvaXIHD/gMjgYjSP
hRGvwG9SSDK3CLsB7qE8ZiK3YxA2k4Y7g+1R1z5DulM90mWxTZHs7OnKBE7TeeMp
zRMeLa50v6uuE14u3W7+uZVzYZEboexChmW4MdTVjCY+koC76Q+TpmWlKCxNOlkh
djp5MlfoyZxMwpN4LWSRm3G9AtR5b7lR6OwlPOgaK/kLIonMXe5ZYQBLrpFBDh6w
UX2asszUyLz8sgd9rbSdR+wFjqbRFc0RYvjuuhYBr8J4ZE+kDm+ZK2qo8/0J/uN7
N2Qj5e0pcY6ANcBQvennyg5kCx9tlUH/hjupsdy6J2ev25yTaWlaPRNlMiWgdu+F
D8iTpC5wXn3sbGBy8fjIGxuO0oU8kBgQPlbkCfWUgYIMJ6n+79qJTm0bD64gRtQ5
qJFSG6qY8oWn89jDr/Lo7LUiYkQ8PGj8Mjme9gNx7h9iRdMT2VZP8oSj1vJ8B4XC
FYO8Rj2WDZG58gTfCwPY1+IfBj2BghjSUSalEd3AY8H+4PbxR+vvvpeAh7uz3b+3
n2fd27OALMKZhBnU/WDHEAbwQDS2kL8f/FOYsw7O6eGrzUI7Xza4CLPTn4AhsYFV
aeVOj4O/RaHpySe2Uh9ACLOGvFeCn0vTH4svpjYg0oR+kFA4Mw4pudJ9QKNR7eKp
GNw9iwIqddkmZg+bdy0Nwi9xweIv7aRWyPjg4CukQgjpPGwPXmF0dqgkVqxwVx7l
O8+/ZYatyV2BPr3R6Q/LDOb3phOVTfZbr3/SLvZqdF1ADTaJqSQS1lFPAMKYEc0E
QV684YttF0QECGRBVcoQMXEpIRyarRF+D8u1z+aedj37hB1HsmxOxgkBt+19cfrm
IlzijNchCTJ80+IXGsqd4vjkhc9dRz2nGnDy+gIl0dUajGZZBn1B6+LRPbtENP+s
CqQ7whjkvrFgEn3P03+k4iHfrk4h1oQTxNd1WtFLqlsae48QI4XVqm9pDE51X6QJ
MIQLWH3uYMwI1DLgCOB4NIW0zHOWo5GAjiqRFkc9d/uZGqnJnqVL/ZYxWlTsdbuK
DS5qRkDz47/7MEeTZ73enx0iVaz2AG0qETy8Ewi1DPMWxqAK2upQHgTiN8LG69Kr
7hZvLlfRJ7mvliYdxHFALUIGoAAjNJuYr/BXPw8k2kWnP0YLAWH9D16q1Srkv0aG
G7ptgtZ7z1lADt4rPbJHQFGdQ2t1CAaWrKxL3MUPo3brwk8txSIbE6nmr6J4oBSB
12KkDaeXNgRLBD4rAOueU7dLFhoUVI5b4zGj2m/HqZMRwUPSbzQuTmolmvgWZCKv
deioJ0wU3jD0F57AKrMK08nJIHgVrCBN+lbwBxTqV18s1KD0pna7sZjrcN6KQang
rp4BFVIq3VIy/lrUQTRP+BxGpLiJIGQYFceHGIfTWWyzZW58V15yr8EMA5L2GAEx
eTYbqz2zB14YViqWLra8F2S6dwS2rcBmokqDhAok79dm1LSCQ+I8YCL4bl+Ddmaz
uaiZ9kKIkvLyTM0i+t8HRvrWj6sjTh/kBIKCkFfxYBPz3Rswc1vXT4XmSjts8qhl
y+aLbOL5cMaP/tO5j3/5ciQZDk87Lge76v5uger7kIjaiZF15UWRkfYuF4GoMJ9k
BOOBs2D1pRZRj7I3VjofNZzPN27XvWUWZzr9fVhsGVo0k1RHNxnE4rvhhaneuHGW
yF0+hLRhZcFslp+LYWZGST6J9Mahqpk36YzVnU+DszXIqH/tU/Qtfv5IjvDaCYm5
GhEY+kefx5UMljz39S/13eeAzEEyJy+K/9pnHtVUAXWvuuu+Bzv5muiJx9tMrN5j
8DRUIjMeH5mDlelWCZm56mj/5/ur7q/HIbJ/5q+brrDidr10ouga8H1Ys1gJW1Qb
vAuyRz4FDov6EuwsFQpHP8ux2+lgXi7OkN0HNK9Z+5VjRIWDojhG3e1ASojoy6iN
on5QyLG7V4b01j7JHrFRCPmg3FKWj7Af8Q4r3ilU5ZYObl6AVTLhNEXYm2tolYqJ
HWsrG8QGYgCud/ZBQkQ2H2LwQtWdxFWVM3m/0hu0/MJ7iCg9T/IljXHQGfu844i/
/UKmXJkQ9ihtabJwnxshoylFf10dka9Cbbk+xXey3yeoxSj+fsVdU3uwqy6Vkn75
kFiu9sy8DSRHo5dv29VTnMZMq9oHgH36WAygSOagKZQ7i8XCvmduA4j647CBj4S3
K4EMv7VAs4sz7QIbUQROatfwsgErfNvvKyDQ0TIOx0a8XV3F7NpPOE5p8zCfaj5y
CvYt/UPeF3YXT16oVpvOzuvnyuKLXxuam4a9ZIy0Ll7BVbW4/Ntw0GQ2JSrH00cg
WhD9y4lfR5s0MLqhtN2IIcq+VuFD57JRxP7Escsm5mHkQyQFKUtCihMXiRpgLcFD
STurX+c0+Uz7Sk2TyUzqzKAzC/zlsZUFYAkOC1D+EZ6n3s0mmqxCafRl8r3rMtAO
uCMqei/WmKyYd14yHzfOM8xwSa5D0pZ4OSqg9WFvDd2koctlWe0NcV6vn5xJFdh3
9ol4oiGAixAbO4+A5+NVTpli2MbAkqpAq/LGFot06oAg8SuHJ8nvBbrgPE1iRyW5
xfMhOBvf65D+rDs+Ie+2E/o926UDtsPvC+2wDKSfHRdh9ndTvonMBSgLGtQncxF1
poqvcf/qG0TJk4LzfScRLc/ll28Gc0afCysH+PD9KDKyuMF8OZHxjq81gZ35sVNZ
+16zYqB65AU7wGq2HaSdF0SCGaTu+sAhoBTco4BZzbN8KLNdBDOViT6hB0qEKo4w
vVSFx7fd9PqkOC+NivZb3J+GdqnMqcxfl65xPHD9ThgMtYGKLFKwpXeOlyPny9V6
sGmuyUwu6iGYOs15yT4vw2OAvH8NGvq1iYF+9aUw1z26Jle/jfag5Xyt0nMVDdxp
9BVSdzKnScGb8Mn4hRrmnmATXMmBkNkwvg9gDFk3AuC/Mz76iZANlqgJ0kCc6zf4
oUF3e2o1ovWyi3pXpn6dzhk8DwaP2B0KzHU9CnvgEqhViwxEqqUPRAsrMpot8SzS
/hoi0/NRbOT+obEu1aP2Z6gTmW06LCKjV5XdbFZmPNJM60ERZTDTxfvVDP618910
+lDt9iTIoXINR3RB32yA1OjKaENOlRg5RbutGDCZquyBOT3yo+zEk+PQ8HnLAWN5
1a93lEcpi/kd4Nu6mZDjFq2wy455PNsstKLVzlcPaErz2AxnGuamDuBq8YJGVyGn
DXxpsS7cacObQnCy2Y0XiPZMe6uaIpgJMsCLDy4C7oeIMPXZX0axF4v/5YdDZy7h
KEXsHdxRcWQulaUHz+WewSqnBCFIV5iHFxZHCOE/SgH615uLoWrlDUXFsKbYnqgP
vrYnLcx6R52jz7jeA8XOWn4Ls3UrtbLavnBVLwvowOGqd4X05MzRStYUFDo4Qdpt
yIfLKsuBJLOfrbS863ok65YPe7v/LKysWNsApvQbx7EYwWUrpDocFVyUCsSo28ja
2jBREXX11kaE54e/nM+Q5ZymdaARMk6MZcas/R4Hr4ZZ8yKcl1t/KrBgdKyz5u15
n0GOvKky9DPheQetvH4nSWWw+hkuXErC0rjvu9+0wxS7cgrrhi++6Qbqp8y+6t49
v5HodPVBtyNB7dEIAxNxaP/Oim/wO6+wxAEj1yh17tevFO/7Mf2WuausJw1YSZ/I
HEnTfor/1nSjzlKDQUrzvBAzr+hTuOR+BN6nUp8/wMG/Ee8+7NZHZhqk3ZDE+w3Z
0Snqhfoo49SEtNeDlVr4I9gIp8DrvomBSIoe9cTykMsWlGrqJfljxtAJZqUvDnCH
j1Mbhu1Qdtx9IQjQh+sNmYhbvSKFsSxKs6Hzfw52OD1ryCmWPLOLnlEjqntBvlMD
3e3kctTXFjSmeabn8jPcmhRHrAAIF9GJuXQfH8pvTPzNVUwAA/t/1S63wf7+bOGe
Crp2iZuakIgsXv13aV/3qdBLsJXZ22GhsqRt1M6qLgHxTOw3oZ4EZCO+mPdbB0rw
++B7StgjJISG8qvD+8VZFADeoRqAq4HUY6tpysPY3T9i3nd4oONhw9OeJWO54b8C
VbpCNWUU3K0d95OK7dIxqvltYbnfxCr0bwxcXE9+N8VgjS+IeFbQ9QS3qcSlU6EI
269ik43nU+bERRAYy+ntfcrlS3OK/pJ0EHsgIVc51mK0evX0Jpc7ZEFM/LUjgrB9
6Jjg2sGpA48vGfiMW6jkZJTxvc3DQu6Hxrk5pSRcMuSp3ZIrna3nigu18YGsSzPr
e1oi1XxMdqs+fHIo3uEHpqzkIDuPklMl6bs/lv1hsOr80ptsiUKtmkLUP+rdS4iP
FefJ4ufjC9yZINd8WEhIuNXnFMuZkU9ofZfodWnrEaNdqYk66j3/1Kx2Dla8FInd
6pRveSnVxsSkP46WktOJA+54xLULCB11l0N1HxRKre9HzcEG4Ae2MwFiINMH5CPZ
KsjFFkFGF22+nhO8k38medG7LeJ2vtg4YuDb+lLmxPqksFJ1pWeVcZlFHE5GGngl
gFak+9I38wj4iuBKlwLp3hca0L3Nkx2r5WGpwUjmc81jW1//BkiLfBgQnUsFsIUi
F6dOWf2+P70EAWa9icOwKGvm/N+MQuiHNwJq1+k4KHikYSptGehAIp7ICoaF4BTG
26mmuPn/M7M+1+W6KZLmIasnXe/2pjUlWaQO+KX4iR90FkH2RabuzYoD0z+H6Al9
/UJWiG2IFhk8USee6jm3EmU7JuE5GgYJkG6dQTtCXvzLwznegrm3OCk6H+/oVmSe
uD1BhPIMWsZEk+F/MDWVZdvCICmTGzyzyTzOya7qkdKml8y1wOAbT9yyAcrDGLNv
dgazZl9oeSSOuQ2rLihbI56SBUOQ0oPFZy/dFVGNYcrX5VyeKjMk3cUrRbWxE6Em
xJD9SLyuZcY6zvzyIVhhAykIJwV4lSwMf3gBdINhMnSUkRcVQEDpiVwSnl2Ot1GV
z7EhgvPg0yrc1Z+aQSCTanbhIf5wTd9yx8yDy0SMNAW9Q/PtavxtFiTNw3Yc2xZ1
WsgyMew51a+ZwvZhXqcCOyoFOgOh05jn3QKxnjeTKmBZrPILge9P3+xUIL/C+nkJ
uTHYrcJXq+x/G6/W7EJaVKJxTS3YozMz1As8irx8ducT7WhCRw6bzliIxWDU2IA4
0A+xiKn6sPxLig+TV9lVgCxCnGvOZy21x6jAq4Cs8ynu34clAqOq2XdP3d61i/JC
gi5c9SRpi5d4HBJ+K9JO4P3ycV+kXlMvDs9ZQibfyAZ/B5x0+U24UVopudx8sFfA
Hky+AAww+n7mOlbQYnwVu8+/1xxFdUDvhHcgLTGA4PxYdmaoS4ql8kx2ov3k/fzT
i4tL8mE+oRb3I7pOW3m6zv+AbKj7owNmpLatwKZzjHyfn7FRd9nyj4H50Fw1QbZp
mjdokAhqi8N1E36C5wFhaVsmChX/fn8Rla8yBBY5SpKUWB65C0cOPpv6DCJnKECM
q4KHg9GmbPbuPIohYgBFbrBrsYkYu4ddTZkmDaAAFNLii1LXAIXyUMKOaMp2QxL9
6Sb/iALVbLTmdft3V4B9UujUGV17wmI3+B2gzPEq8ccTTrSJwGDh0QO/Xcd5Cpof
NJOk5yqQVjbW5+nGGQMFqGWsfsWr/cr00UXvXAtfGgJREN2eDtqBNXojCzePIW7s
dOxFfxrc9e2/3sqtjTzZk5VIJSj34G6CpvEFIJ4wkVWePcG5y5IbsuFpzEBU0n5X
mWhK+p0FjX6dF8tZD/kBk2g67ihwrw/lNazfBNKqyaPUpg/hbfLeRQK6T5d+iETq
R6JLogUOUvzAElsHgB0Nn0KKEM6hb0dMFyhfCVDMuzUpnXWsulyeP7SrLoFzBoHK
Seh6NOrt2kC5uEiEXwaguqdpR6KFZchQWcaBgEVfB28zmk5dvIM9se/MWQJWcTOc
Gwj4Qoi7q+z506ou0UncTciDAfeX2u1urbWre0b7et04pDA/N+rM1vqh46FQgBU5
35iS7+kPx8iGTfWHn0YX/QkGXur1vaxxnSo5naiqCgwH2tKmGJI5dLNE+zCwmeW5
iBp9aETcx1hZkqu1ukDUL6JqOPyBm8AKhNru91Y46zC4nxK4g+DDLpTzdZ9NQNfV
wjuVvskIOX5O7aws9FFKxmEagqK8xonSg059PX5xj2uD7CejdW6ImujNCrO6Ml2h
v9KOJrMpcSshUVdPtNbLllcDfWGFWEjaV8K+02nByKEZQdLtwKxMp9z640dWevoS
ybqRBjgxdoLgXPVuzQBqT4BkG3Ka0Nq1PEUuJyBR0IZ5hBEW1tyfUNZDeVyf7J0+
4dOYWap5WgYf/MsZDW7xWZ1Mr7ms1jVy73lwlnPSfSUmWSsbVxSpNWmGA0aU8yLt
LW7mJ+Dg3U4Y6rTjmuCPS61C6+i3/YOlxlwZC6rPPF8FVzXAunbhsh06ggllPqRz
6J8F4PabIKCMpMVjIjawDZlhXtD/89nhhp76RvI8iWzeqcPljVZ+Sso1Ozm1FKfk
CfD/3E4zrhl1nbX4Djgi8ONrGMW4AHy2zQSw5wK3YZvWAXccvMse9QDcpCPQ3egc
ZM45KPbv9Sif5zUSMEMwehVPDXSojQ/Q4jsyE9PiJSbJabQzV1A8FqPlzfp5tANm
7fiRNBxopZxIh1rFc2DqC1JELNAOtxa4RqptA7Pj8FQhtv6mLTaOej5o55PHfDbA
CgRlz29DUUWUpJnegx7RIyXtp1HYeYaT1KfSxYNcepCTLvhhQZNm/aXfycghE54k
84dddoozLxYZ+KgQigQeMTaqCOP6cX0C16gl4AUg+OxEcuCxlorrzYtiZJq5cGTT
88mYIRfrPTZzMkA8bOYaAfHck2LI1vRDWct6fiIEWXvlimI3azEMHkbc82X5Q8RK
dSEzc0E5Xj33zgE0ezmMb1h6XAK6UXdavucyD/JtK0gyoJ2nSbRaOayQCFmRR/oq
vcJKNj4KSkJf0yqzAOEdUTgnawCqhqhB3LjSquJR7qDluK0LI6Pv7gIGPJPWZyGs
DrXrEMxtVULBDd6LEIH9yfBwTe0tbb4doqrUzInezbpHnsbbjZQg4YnrJZrOgh0t
e64fyUoij1o5v1k4wq4XTn+Cfl6uqnCs1gOF25T7BWH8AB0aYj9oPjDyEhC92F/1
qt10VEtgW1warVbB1TON141HXNSpdz0gJ/gPYxg+O8TncO4SR4oCOCXGhxJEaKAl
ZZUA3FjraH6ZEiJjxK7VDia6DhP1gGGUV0seBvn8PXGkOcxUuZIXjO5AGAIb5IKF
a6rLKVaVtVh3gAlp4rwcPckxt3nnuMu/i6r5U45QSCFSb7DAaStiwCtcKk9oLDZr
8R/u6Te007/zEag+u7OqrptRTa7VeSjLB+qLKa+Hn4/0RlpTmktQ1FKPPPsbM6zX
7ip5V+4lzPiEIlTQ2OuhXSifXyucn7WgfIBzfyQ0lQMfovInOdugdQ1bFHqYqLOL
+Acy2zoIBHPqfSNcd99UC5+9bUmpgdqy6RXqECCh7lW6IIUiy14F0ChMhcsCjV2y
/Xfygydu30ixJ4AhlwZ61l/1O+VKU9O+CXbgqMzlEAhSnGMl7qhmpMKsN4qj3t+R
7Zp+z18I9E/SFKFqibubM3RohfUxmr9qIpMDD1UdCyfKmVfVxggdBwgpSUoKsQCm
AEuhBj5V8Rgdwk4WB8OgY9/633olphpI5S9QPu2UJRZ3VemX2hOHX3ArbuuMkius
HCImpH6Rn2SKbZJEQn3CbaASpwUnfuG1XtWdPB1Yr5vO5K3iYvIgYmkfv6CjQaWM
AwiowpqW/vqV40MiawI+g8tCy4oWXIdV89RNWmrnC6EejIok76bIl4NdbHJW2iK5
P1REye/DITg0v+5tMm3jEauD4zLkXoIVjpEGmaSJqGpyUc/xqqbrPJQEA7Rwq32X
6YUiLG3WvWvcFlHqaKFwUQw81P2zS/XbNNDt2B3/wAJ5yYJOpdNBGwg9wJkY7M63
u0wRQ+l02ZNT7JeujgEKGM7xGobyZQX9/mxpqrrejkVbjumnRHnEwCJ79JHFazm8
Z3flBSaAXl9xYF0oxdfg4FOJnXJTeNmbYSrRFqR4LMBFWwOF2IjjWi01slaKgtQZ
v8f0V0Ehb6B/zbfwbdwzCvqmn1y3pwtoFVhzI5H9zln5s3NHHThgOD1rinLY+4qi
iqHZazXOyv0jqzOazeJbyTnNFwCqkI1uoE9DX8K9PN6ThaKgT71kGJeazwwTcGSe
OtUCYzjRc/3EVj26ijfFlkZZVmlDlCpVeeljDoUTAt/yYKSImek6bwEmNC74s135
75HBy9YJKbBzT7Xd07MGTsnPgpKchQoorMdHwgH1YJm8ENOer8lQ+aNkYT6BoOAM
BCulKA63K85JOdSPGccg2EPRfIaJwkX6o2/ZAkJlMA6hrZ1LcTznEpzwAEgVJLwC
Zevxudt5HIbTJzUr6zTQiVLJGT0+4DVpXSc7oUTNr4cgiATioNTEHCxwWp8HeYft
H9WsDod8mjXCHDoHusU0OL3d/H+MkJB8eh1EaihYSBldlaQLDEG07+AN5rXcrCMk
+KKukIEbKNklDSEimRgKZ1Weld095KbWoBqVEFWM5VaEmMDtbFU152Ka/LesTE3u
jnMPk0Tbm1OHvWjX1HDroCM6I2+vvYSssOCyaroaoZzDHUU8TDnpAhLC6XuGqJmG
jzGk+fkDSBAOXrP3PME4fqN7YjYuneixVgFni3oW88uhzUqINNEU3JFX+K9R9eC2
bhOLhDpn+iFFGikt8hKQX7LD6QgvS6c17ihFshIrDvjOhLGeFHu01IW5z9UvBheV
GWBZaFQCCOveIhNU72fdXHPw5rjMo7uXVeY7vKkFQn/crySP6Zq2Uo/YJoJNL1lc
Ag5L2lRalJptz3y9bJgapqQPGMtMZ5CfpHI5NNyp09GJnao4HEvKOB1rCCy+nWeB
GeMvCdHZ8HPYLbNutDCLMBM4n+Q4crYVwm/Ld67kcCH30XXkzTGUN9PfhstOXwQJ
RxNGUtBs2JQwUwh81FAvhpDaBK7cOW5rlAj79uw01aBSyuwg1zVo1e5PnSQqXCIF
laMGDGrTYdy0foNNKi6tgKGtgdxY3z7fUmABR5TsttXzQrSeOtqKr4GdEfCHqNyl
hxrV62GV4cGmoPXjevmoCbDeVV0aFKWQ8TAuCFKmYGNqUsy7o0V2XQ14Pn7cnKTP
mR5Dc3amAK1LrL3h1PbAe/rDsY/k+I11zD+XGb3TuY0HOfsVGPnlRuw1n9V2b3ry
B6wgWe03YhWtuBXNvCEdLXsBzEMcHLsZXGTBDWOAGd7acatoQx0FQVwKbw37cxeI
ix9oQlzfCcH+H0zatcBEdrqRe4/gSwmcXw/C06K4JlOQAXW9+RBWO4RwowL/edkX
yZ/YfLP0W0rJN6EpHRqhLmybJDNfMGq9hXpiPOBLf8IyZXT2iSVLFbBXHamduezb
KJFLUf50GBpOG+XyEvHhNtkZGe6MqdyzJc0/XJYc+yZx+Tg7X07bZimN3iyRgve1
a46eQX2dVArzZScPWfS1fYjLhrzIN6OsFmYiQvIFj6QpaEyGY1VrHkjMuXsknDm/
/pR39RHJS3ugZS0IDpjRR3zzAyT3FXNduj0Jk8QRRNx1l23gm1JHOXHjsLOmkglk
EDhWAv+7LXRuHP5j5MKJ3rj+UFbGNoi0vlgXqokX2PEOSuF96iu+idHPpCRWCY6y
LL6s/s5z3CXW9NUyTNUnp1lFgkiyZ5f0TJ0Q9rDghWn7pZdAbTAWg6bDoA0bIlN/
j8Ue1asMPE8XtyE6p4jlptkAFmTJ4J2QtQv4ensXp2EY500IkCwQWUc/GWMGTu/b
B74FX7Ocfatty4pRFe8BLis3f6t8rRAuXPHlM+Sd0g4Xh5HusiZ83iFU5RvFokkY
SO28BwI1J492240z0Ft9gAf+5ThtliYu3dopeLVSBa3VQHdxSDX+ZFoUS8+4WZXk
NuIyH/FMxcyPoXIpDSiU0c2Dq2b5OguDKKTRPeZcHnXh/npLa1Cldsxl+5JMj+QT
8pK5bDS+lEel5PmqvJgXTx3X8gBiXB51VFjEOb2W0aeKNiqE3MAR87/xxuFytPKf
FV/uJbVm9OiltHDsWxbjaIwMQv+tLi2yqKbA62+b2kaSeMquLUVdO0JgIfM2/cmK
O7dqMOiNj22aDTJPG6w7HXTkuXDRuztsEyTxdJ8aHhuCzZXsBn8C7I2z+ptm9MqK
CISTEvAV5yJhGv1XyecwuqnoXVMag6be6IgEyuP9HAnagbeA91AOaIQItL3oSCq+
/d7i9sngrurF/mp+T6+tIj9PvYMOOvIe7rzgxQ7P084GeNYzrbohbmJsZ69TzGdj
Ngrq7Cyos/T30bshqpRB1BorGW8aLunfKugfHnrioEBgO7vQAPTab2g/XA9SPX4W
eiR89l4gGD3lBxH2kD74aIWSqeE6QRYLp9kO7AYesbVj7dVt2ieQXZZAAeCcpB2q
1J23ytuSK6+qxnJJLQUb28HK/k30q8IDsY+8c4ek2jgrIGMw/JSV6KlSS4wMbvuT
6aE3PIHY9WouMBarVF5EIdEFKDijyMTIlDP745yxXKKwzkmWq0oW1X4f8SLjoi1R
/U30s6R40xmpcfQth9FUzrk440+S+WsLP5qO6CZbVzcg1Jy4TW10uiqOvYWjmk2e
mnYinRe9GWuCeAC8ApCrc4rNV2yfjjnVJXXYjaaT7O/gKKcC4DoD5s1ZXuV307Bn
W+ke/KGV1yOE16WPZLvRdEMFgxkKQNK0LMVu8bdvkiwfHeP6EzBLfMYiVdx9kdl3
CxnSXPQ7xxiD4sKyC00LgFgGTntkkjAmGJ5bKIv+rff3WuHm8PpExXIyniAaSSZS
QitHd/zz4Hoqr0hzt5O3F3RN+llXTiHIErlEfSmI7dFgqeEdQ1kWuP7uiw6MT/Zh
qIsgkSyI1jFbJro3A3GKIzOoCS9zKf1q+PoaWtftvcNygBxEP5TyAB8Wplg1O0gn
k3M/lfag0GGcrWPgZpObbHZdS5KFUgQaUs8rybyIMZiqJWE2fBNs8/TdAizHSBNE
AcvHWXqH9ow2nhr9Rb4WxUcFAYd0SOTCyR9528kGRDAnL23JL73SDSwwQ7FvYqC6
fgbUUTSUb2wdFnK1W7gussy378LlIpq8KUa9cAAhvROmhxuLuBK1rv9GpsRdDTYI
UM9Er+a8/PMQvqcO1zchMYBLIGf4xLW/TM1NfkHu5xso4oTe7zOMyIbJ3bxLTOjG
eadvZWRUDaSoTLD94gAe8d2CgbKbiI5Oizm1Y73UbJXHN3Wf1IvEH+OBZ2OllpST
gidZcrvythvxi608dwCAUjfVB+ryU2MixTmUFXiiaqscPLgaIE0HU8XuTHhl11zR
U3yTeirzAVKwdFkU0/CAli6Tx/t7m8oMCvgwFZxwidZHMOy+Egz/jQ/iF5Gp61wT
gtTIMzkZbsvlTmU6xz7QIBRu2w8eBcpmMkavZHf0qkWRUFc0vd4mAs+09WIMar5U
j5COYnRVKWU8KsSRtPEFUDhsf6NosyPg5WhB5+gktryL0v3L1Z0S9N378dsq3Fvt
YyvV3ouqbYRTdtfTDakOmnECpbYuqcjbpSU6DN5sIKLLWboMR9hy6p1DP6d6U/hN
XuGuBOBdt19Z0a9forJ87ZbTW1ufHN7k9FY8EHyyXiwdUAEzA5GZ/WzqJc/FXtPy
Fuc2111soTDW/QSctBI9Trlv+fjRkaJv/7+5tkabEaSYuekh1do/FCfgyZc03Tn0
s5wlFH1jDtV/BLUVwso8k51iKdyRGfb8uPwtBlbtOHQTquoQIhSZZPv6+uDhIVqZ
9eC2BzWMdX1+WcQ+q5S2Q5OL/y5RlreQdBmS/RoU7NedY3FOgQ9eAL4jsegR6L7A
d3u8l0CDRrz2TWEmdyfMRGupyhpd2Y66CIw/nh3hr5hc92mRltxNCZp7WJs9nwH8
I70l+OI4ppyCqsQeisK7vFeBlW2ZsU+JgoZ0c2JHSL1RK81yN3yKI5okShyCF4PU
6HrU1Yu5m4bmiBjjcGC+3Ci+TW5qAVEVpEVgxH4npaL6p7Dzecx90xn5qZ8W3+X1
thMPK/5nblSBfXvHyYrtT9+yTrYxOxD5R3pdx+oOCCOfjVqQinHGQnt6V2LghpVs
cdthmAgsUB62kT2AfqKTbP/uV4U7UJ8uxFvyWq2XFWDSrca20uwQOmuKfq9ySrio
lpwvOf2jTQlJswxfyvobSlWxMJbgVaof//rLGxirYBepvoW8JILyRnlAjdb3NtxR
fl3pRdzSW1OO4XBsTTsty1ZpE4Sf55mPYnfUUAGZvjgIb0UueK1FNgRGqU0ssl0l
NE3Zl+Ylz0x1kTkhkLes60MiuPNmju7/NUlC/GFf9RHjC4VXAyzQp1zkD2wA1PU+
6LYu62nfWRsa69ZiFUBTf590oAmKl+w3qQtl6VRGj/33izZpkM7/thSLHbekPY5c
p+3kfmGbTZm/aNewYAgX5bB6geRO4TBdHEFnMw9j3RBQFT9UugKp9LhsFVUMg1dR
YoL32cxPoR6/+AD3r8lQLSkTYBboHhfFwcrETku8BSgMEnyy7Lcxc1L/fi45dW2/
wZlAprFLADAGhtqIgc75rcefQdJsGmL2sp5oAF+LnJ4cALZHsZm3czMjxGd5QqWd
4N5KMesms8tCjCpo2PMgLC9/X0SOS+MzNgjfKg7E75DDyRFzSjyzKvJVSL2PXBmh
uBQKUBIOUkJZaOxXisqFpe6E5olIStpdX4mg1yWhbiU1nse04FNMV0Erx1uWIi3U
yahtT4nmHUGLpcxPwjByxq0JylfY3cVXIGwlehB2y0aY8ZnnEJSR//xQVs0vIqos
IatUOGSnrz+w2Yq5ts6Yc5gZUH2WjITJI92EO41lhWbrgLIxVpVD3ClDfkVSJW5k
Xhb60HdxGcs+AwX1izHZ3wTCgPzvXWxqvTx+JeXTZLCqP7tE2f+RYHVqQ2yMkG8Z
NzvAI2pBgucv9B7lxHrdo3IDYsP4hR0vPB35aG8Mq+pi2LVpUXpRWd9c1yDNtfYe
k3ltbLmgq8xpCcKStfVdBO+3AVfEdyqnCPF715NQrvJWa4GuMc/NnXMhXABVZWo8
ZGRuroH58HOKv3boBhOKpt00nPibHlk4XW3I9X1u0p32JIw8sQ0hDW6PmRe1Hdne
bSH4WWjCOSrW/dbN7OYxK2futrJ7vIseoBHrgMCgiZiP264mSfeTSOJw/Vf9wyX+
g2hoJc2sW+ukWUpwheUpcgO3YZCT3yKJ4PxhZauviswN3OnxzyFNvA+8awC8AfjM
mF5Vgf0RV21S/mOJOyuFVeZZcM+hfXV5fJmoyXuIuumVcsdPgmSb+Uf4pG6qmrs6
9RXozqfMLD7zcx/DU1dR917Ioy4VQXpdTnNxgo0Y3NfKV6qS6Jvg31CiMF+5wfdb
I9Pz78fU61WTZpzY8NapPGM5mhxQ4UY9izXF6NHprs2nIQtmYNrPtF0ws5vcfhON
P+u2lbEPWIZSJlHS9CZt/HGSUmY7bvTFYMmbZUP4TNg7WncQd7gdkVt+mmUjGFsc
SXhN7xtk0E+JkiU8iD3rG6a8xiaX31PgQwPp9EdF3Y5kaETC9YPQfLzZiKcuoXT2
6wDdIt/tmFj4t6B7my2WxwT+i6St5JW1aBwCa6bL2QBkudzm4hSRYs5BdbUtoRaG
A44k+gH+SeN4Ow0hA3xc08uuNFK/70iJpuKC3ZXyunh4kDmz5+tYKPO1JaSfM/W0
HI8nlxKSuA0JvbCxIEQPlYtUwk3GPbj4+V/WksDMYDEMgcvRJ8MhtOT/6tap+ZIV
CeFrlgpxcPRbXFMXYcVX/ePESAnjNTzDOT/fB+ZRq2cY9JqQ7ZmLT4pwUepaorer
cORo24wUqx9zjutK3CDPVvP9GnOoMGnDd9xygkwcNltr7BH1AaQrvBs84cX9RUeJ
Ffd0th/WSUITUaHW6YiVEb/PwJXdWzAoncGLpZXCg2lFfRQpA1Dju45E7aQIwriV
taH1NeuZdHUnWPTe7nxAex258zxy+1AHOkjXgLV+RLvI4o94N3Leg5be2Bp/g0w0
Nre5nCZVWkOO8VI4hAw5uAg/mj1y2gKW2s02jz5Q8U1+HEaOUxI2g8B5J8lLjQve
ZUq7SK91M2jbMW5n3HqO2hLhBZdOnOfgA4WbZ8GH49u5I3CFg7jNEHJw4EwUciHe
pqlQiqnPg9DQhLqNMoxe2mcXYg9tVi17r43NcoKAMpppKQZMrTaxyLM0AYaquR4Y
XrXCT5RjMKGT3i31xMAl75C1XSlVvCnITcaqmy1JDcQAjADWwCTp7hwFffi/DaOe
NunLJCorM1IOgOCHP69kYESYisvy2s5tI+bkyz+Yl4zh3oLwClfqPnf6e8arg2Z0
gg/TGW/QPOQPguU1zn6U6hKHgG3tEozlW+qVX9xQ9Mn059y0rOZKiQLoDjuvcGJa
6n1ALCRY97wG9WV4E4mzRbvpKA8qHxRh4d9A0vKiMYXN4q2pSNxGOhp8H1FiNMj1
FjctLTMTZ1ELCSSdzF1NeSdvq6L7cVacoBiBpVfd7Wn+oyAyxMKAgj8lwJpt42q3
BQsowJsPDMpuXYCx5SiPZemOvAOBKwBAQfx0pXMsnKO1xRJWjMKOHZ43Q0kPhTGd
0AXdocBzrHw7HBW022BXhINzpICheZrIwlLAWtruX+57PhQxwqNfK274NLsuskgM
epQ6WsEGcFw4VAIopy8bZ2S7sTCu4IssNMd8RRG+EIZ4inHZ9nv3EOlbY/8kA0sM
aIzEQoQTDbCy54k+LdRrM35g/SvdQ6WFX1NPgk2/XDsO/eaHoY6pb6DcUecV4Sd7
Tj4fAn8kI2xUR/lGEGO0MeaQdsbeZP7uWR9p1NSSGEP6mt32oD1mfMlQX+WUTzm8
h5ob/BBFULI11hh2h+dyTAQ+8KLulA3/tZnEH6QOgGO92HL4bFKYDYcO62lJuCs9
awwHYgn+WLN2k48mRKeZkzL7/Mustw4To4GbojXWpLwIXP5uO3wJb1Fwx3P+jCJd
WjznFkPycs7YXl7KXwSW4J0au/+vFfPqxdfUV9/dhVcHNa0KZrtJ0ZUSglNzOadc
LDU5exz9n/u3ndT/pwryQaOsxJuP0CIuHIYDbeqLFoKo3xeRRatWFyVb3BAobrXY
nHK0BCskOTrWR5cjnSLScaLu6aeL8npMHPQVxVSY0+k+cQLAiEKKYSBfrM/+yFDc
kTrVI48+TE7L/aWwLZGIx5tgH6+WPMepbckNZzCAw4PxlV+zXyufx9UXYI0NuWWv
8HshMRIztVHuQh5rg+HnYk/qPoz+OqLY129RgNvQ8G+XLtSfea1L/qRY3GdHghoH
hSrmChEoF3FwdqOhOOoPdUfo1McPBsXNqxCeKnsPS2M7HSuD25F7W0+Gkxu4PkYt
aF8jvDUdQGR+h6YOUvtKCZQbHJtuUdCAfQb9OWHNrlRrKGt7xiayIYq0SCu5KJaE
1S5cExQq9V8483BOVWA6FStsnQAxDLMmE3ErmK8BrcExUDTkZfcXfThzAJWQOmsm
jyF17iM/uU3T/0nnxDiwRNyYwS2YfoAiSoFoSDLyeQFIUD9QapFMCXfRg48VAoxJ
FL9VlDpVFtf6rCOFArnA9iICgC8CyIaKwtrCT5QzWJUJ+Kz1jtSr1EIkAahNszU3
Tt4icOD2avfAa2OdY9KChixxuUQdWGsctwdtHraC/FW42HzYpiN/+CejGpQBQtIC
RiWqJsMrwCZnVQj7cJf4IcF+zUq8BKplDW6nfWk9nFeM0sYuv3UBgiS+SMJVXzbk
3E0SbBt2HTNKbA9caQlhCLsLXdcs4UMc0JNnCGzSx4tEqclFjmibBbsEbMKyNvg7
spsOlPwXA6nl50k7U6mGUSszNpiyTMlwA5zRq8mPI1NZx/OpOgxO4GV8r3MORObO
shbctbe7qoDZ6WAPG+RBNhfyRcQxUi9AMKp8xAUY82j841S/eDgYYYEPiTOzmdpw
It3QtkbE6bupjUZmB1AnIfFPATtnRSlZxAtoHhR01acAIwSucj9PHv+m2G5/Fz3J
rBub9C5Dw0gMU0VRh5Ykb/QbG5ng6k/S0AuX5VnDBAqftt6P8E8jqJpAbMEA+lVo
mOECWs9P93JxOoBCPxgxRemZcGGsvBKzfl71JnyRksvAmQ/IUZb+kdMZK2NRI01a
wdm2i+jB9tQSKOMefihciqFwCyH9mgvXSRhVPaPaN7IrEz0iPu45ylSIdZWzfRBq
M4Ca7f3SxLdX8m4vMMBDiZfa8iHRlGXL5IFUcHRSq4jiS62RVDsWaiOrJxp8T1O+
AyraZzx61o3XEK5kGNAHJa4GkKIdwAIQuF30TLn8EnSZcJZFCZdOgMNKO8x0x0dB
2K7YyNdQ2FDVpYNiQIQqUGApaIxsp7xXk3mRCgBkS7dmq6wmArhgFJFgDek0AkZ8
WTVQ4y7opi/WJDFVcoEDMhUelFiUW/0JAI40V7kAvaZsFDPb+CzsyGpcqMqvcczl
TlGQwkvmC++4JvWXWaEb8R6ursEDoP/4vbnbhOXdaiAS/v/ThzGwCTyYwcNi3fnt
r0fpKuDrXFnKCkKzkI9Jz4NorZ5nUKk7Fsz6qxC9f3/AZf6cpQ/8KPO2eTf4d7Ba
kpqTuwunooEVItbJbSSVc4UBM3DfKLzULVbzpvklolgj84pYRvAtjR/phm8mDFEx
JYRzgRd0jRwgLjlt8d6waPdl0mq4SO6MdcnPTu4TNpqDt9NTJ9l6Mo70G280nMm2
dBdQP/k6X4p0FynGsq9cImUR4ysJBoZhep5qWFBcZ4PeiU9cQCu5Du2dOIP33XR6
KBuRrq7qoEUMGt1LET/ltmM/Kx3ath5hdBWD8tl1RSoEdFeHagAJHf0sYF9yHOvJ
OLkRyx5cK7EQ1Vr7ykbYgtsgKtY6UST4uXVFUnc+36j5pPPj4+3teAfT/bqJhW7c
NmR3h8Ny8p/SKgmzBBwNIw5I4xBm0gmteLU1zCJVugk7bZYRO95PpixhD0EGh0D1
9mo5dpndiAG85r2HTZT3cp7s9Us7kUOLgNDPMVOIug/wA9SAGPheGxpfrSOYmQa2
5XyOU4YbRK7xmWJh7yB4bHK/Luii3+a7LCor+nJY3e1eVjAOAOtFLz24/IOY3W3J
TWloFMciWQadfanq0OkLq7E1vku7JGdEqRcR1mltTICkRPu9kDWyzg+PAMu1maQU
mg4H0XiGUmsuhr6Yfk5tkSudWI1z5+k0abzQDQHJwIaUu8ur8mZlC5iQW4sUeoAA
5FEOtYzrhgdlhrXOdc2xslpFEdUuT2GADg6pvyDuGmir7l9BlOqCdI6g1sMb/3h1
qNokzkzndZGvK5vgUjdM9b7o2FPz5SVAZBT15j4hQ2w/JwNp5oU9Lyw9GKl2dlbv
PdIOiehx7v2zEPTxZHdFnKv87dYUE7AuvIagVkT886dZPxo93EgXWN0bM2EuXDT4
CaKkBD5bfo+P0KXU+fZA1+S+llBUI4ku4038ckmtaeoRlRJP18aqaoA3c7Rw1tSI
67NaE722jJsL7JEQ8mvKHLTGzZeLITi1x9LrbFY7pN3bdoB9NfaUBcRpKfHFAWqn
jCd0KTaGbC8PN2PZ0toWWz9xbtWiZRyDIQ8PzRTN4IjbKjGE8TFtwyNAobCDhRzs
2r9Ywt1wzN+5ExF0cV3alCc53BCMg3ebxNyh9eXV8ocvzBRGiVk9FsCqT2M0IWcn
9kts0UKo6S0V+TiWHN4gUU7bDlYZR7dHbdnBcIjqjquc+IAs2Y2EIsUkOJQwnoIR
gRU5jX4jchR6STEFZ697kRe0QyTbvJ2qjNMVu3tOWTgk+ozWoZxxOX9mVzfY68OB
EMioIkJTy+PCQ2lr76V/Q0/sE10UwPDhcV9M1fHz1Z071hO8wtLB/9EckNPMUvyY
szUjnQVYy1O0LluGmTVl27Iv+ubHFV6KP5iqWapUM3AyVEaMZBHKi4UOlUV2Ozcv
qL4sNZ7FJEFg3AQSk9yjy/WetciaCv8sS7FX+X/QjWAVNDOxTwuVSuoaaKvyyYuv
btAm0rIfSVkGuRj6yJ5wcaqwtCFSpGUcn8CoYZS95PcGryglCDN+rXhbnzBvn+Kb
aFBynzqz1sHS7gvwyZ/QtMQnWhnpFOtua8VC1SQYm8pgUDYHKzGp/uJfT2Pv4miZ
JkpK7o+6iki/p3l4kZJGw8TPPlg7gwtic+CI6GWKHUeFDi/bv/j55KnfZW9TndHX
ewk0nsRZCpyT2OAyaZBP5/lnABbZkjUm2i8dWWXtL4O0qEsx/DO5ACP4nL0tB1yq
6ZpsOUe/8/iH9q5nX8OjBa6Aa6lR4rlwr1NmvKjd1px/hDbuYJgM7es4kkrQ/u0f
P7YoNV114xjSUwXMh/m9pKI7TUKrudNsLmLL19+wNLlUg+3vgN2nAunEjGtnr844
VtzvS86aC6HrK9gHNaiUOCiNFp1GC2Ga6Ob6Fthw0NaJ1bhxQkPcVMtEXQ0HjD7V
BKa2BVhs3Hu5n+OeqdL0nUVt8rGPdSW8XbwSOLI22o+foesabNF3yHWDEj2kc0XZ
qpWBZ70WasWj/76OGmVNjBxyLcfS6J73V/yvo6eJSj11B9fjiwYk9oSplLIjyF8p
0W3vBfdWmJEZEqQkRGfVa4Us5OxCuAF1Ow7Ns49xa0D9TKHfgOe90y9a2+IsuBOy
uLruqwVsuyGhRPiO/TKjML3alCFC1HB7KU8L/I/mq4TwKX+x88YCCTWRZi0MT694
n8Bag9d0jI6PDisFTjO1sk/WBuCGSZNwBE0P3bADYriC4XChn9x+A6V1S6EZQIiV
1xEWzHbsmICZ1piAtxSHl2bgOO+lyvmRKul+eA7KgQgsX5oKR06rYyEbgsahhuzd
ar3fVRHRZLkv6b0nCJjVig9cIBakrdF6AfYI0uQd+dVZ/wkRmffQzIjQ/0uyI4Hw
t6oqJ1+8Bf9D9bwigOPkWh0xM53QRorVSvoAaSPG16A6rVpKmeJfwHRxP4t4aS4K
EcbIVd5cTngrtDjtwyCqQTjXhLryx13qC6gzJWIxTIHC4L9xOPw9xCVKFzEcTmfu
bny/MMSyIreBdB7OhcLTZGJQUOihfH7hCgavJYUqV3PnG+9KsyHmi9RglraVIXuA
U1n5EkW02a1JMWVfhVRB28Py1AQTULGhoulH8eN6vKcmjoX7+lAbNwbXrPI7NJr9
i9twOtLvYRN4mkJuL7xU9gpdhhVb+1WqtqSmGg+pOEsRey5TjAsd48rvP8bBe/yA
FTC17FwXXi8bmtYK26IP0HPCR6fZja57EKt/6QrZM0VAN8/5R2xON9WYa6y0sWML
FR7JwSwEvbK6Z83NlMIE/TjwHxLwjemftuAGdTaWD9yqTpsJEvW+qpz4f0mjgcgH
LPm44mfrGMj1QdfwpmjPD7elVbOZrtbSySiGcEt4mam1ebXf5b2643KbhCGxFReD
pHlvr09n+S+zwKceT+LOHF1OiTmiVgZA/g8c5zypM18UxY1hvLzixe4+ETwLHu2W
0zjN8DA0Np4t8HZ9CmXVXGevsQ6VDIe8hvI64cLCsWbIUSXfz5kob1sKZlcKPUMO
Pxb5DK++SzcAgqP+evgdw7Qg91T6/Z8T5SyZ15KlvplcBq5WHXkfaP2zGNcsaEGm
vFAw3nC4/DOvgO5vA3dOZSfj2BVpLG5QeR2IVm26INht/wzlf/5rSYhG7jBR4M5U
ieeRt17qpB2fidYh2PCx+PYlaeEyZvDQyFXOpcdhluhC6uK+wMQmVwqYtePTgWL0
vi1SyKWgotTPr9EGjJ5Ejo1RdJWiDM8e5PYe09I4HpdPmIQ8Dr52yX5JolnRbDpR
lJ7CT1JkZ9BDU97wfi1xqdLRNbml+E4//GE213fe88+iKTy6QzEjEhzafQGzodVW
3DjbeXOTd8Tw0cW9sOZ55dp6PkjkvC/JgLT2d1BrpYd0pGKy57WdyugGHn9Ysh9y
x4PMzbuFmbafwVRXHORcMALy0KgIC8Q4zPTPA+XFxV0DVCoA4/1OID5AJaOUsGXO
3+1P5KN+ToIgnzKiDhIjfRjykkhoV6QoLscE9iVQ+0xzLzbWTuDlvhZgcpbh7B6u
Ut34GC7sVip4f74qDypvReGC/VyS8WZdF7ypoJhYp8ol0n0T5gpeAwMr7MA2jSWK
kELFerRddBgmF4wFh0tUfQvyAG6ZOxmHwH/wwo4J+jMZ+haTU0F+sZTv/KKLleRg
/iDxo81Y+FdBB6CV2gRZTwzF7fSQT3Ae3Z3BWgJQlm6sXpZ1GOWRzXuEUy0h40hU
fT6dB/bFdW1JA6dzRPBov+fT7SkrcRpzxLUX7fEXlAZPWJXP7Df5YQF1LUicKjWT
7BqGoJwbq74d5xhaTAl/xB964NU/o0/KGMCK2NneyHROXKtPVsa0bz+ZDnYfGk/m
mojRidwTulpsE88XQlSG2wnkSC+RpvhJlQELKuhM1G2WApUzfdhrxH91p7A3SgC/
2vSKAzENgtUyzkqDZKzFfmZxv6zjh32ILJVUMgVS9Cgz4fM/IQm/SIFdSgvZlKsh
M95i0hQavW1yOijdUiiJwsKMMNgkZWVHIvKmLnKM4ycNjkAlAoJRXcJcx2QjqrfT
2MqXNzp2sGsGxy1tgPvweTMiu/NG1q0BPAXzrw+pT+fxGkers8Il1dKYdCI72hOJ
GqhlpHDl6Z56E6YQvsTxwkIeexyEOvNDhDroDCs+hfJRdv3g06KAaOY3VKqJ9KZK
hFN4EiC9BVev9juq48DWJceYVCrGc3AtxQ5rM/l/NyeNhy0QBcWbQGSd8TlFNXJ5
bZ/dQvzw4Xj3+cwVp22tP5aHgzpke5gQaLKQP/QNz1tMGuykJKOtLsvuc1Hn9bNx
e5sGlGMAkFrfp4bA1LZ1V+0XFgSutYtS4QPeIhePHzSMbX2DVz3zdXz2QAkxB5Jo
/0SXOeuSZFUXB4hYhs2D2rmrLBG/67p2uUKAsqS8j7L46F7171yO9rIywUv2EMic
WPXDDy0pc6GxJsRNnJy5CpLV06IFzM7NdKJjzKSuoyk2Y0kDDfgK6fHBdhIcZQCk
D1gJTqaMYy21Z9vQSmb7My+dtkPNkCWXDfWEgWjwUrrG5XdHXz6UYdhlg3oQsqJI
m7/ABP265/J9XKYlz3ISn10ric1MD+3TbF/N6Eu4X5jVLLG3bMtdGNZHBJkCxR/8
YAyUbj1kY+s/l5R08GEyxo6/ixYgJpP0D4RXFUmwNuuoDBGVdzvMNjP4yfeTVfr/
tNWhi3W5UqBFS3C84BAwp1VkoJF13WEYkndWTrYF+Tun7LG3W7yAIdTHITsjYxht
qh2Fbnj0Pq3HyC2kqAmf3BsaFO7umBeQTLqL//RgXHwiwe0cD6VxkK3ildHnda0M
2OzysDuzSZx8/g9xSLOqYusqFkLTNTBUYuNcLtObepDaoOx+taQ+z38fCtRO0/IS
v8oJUlaEfMp5oTQgFiZ/sIBPaZud5TUjLSxz12e1TEt8Gpz+fZai63T/SDPHKv6f
sqUx0RGq6p/36mS18jqxwetSf453e3dGasS6ZmZk4PhQG0/begcXP5oBmh+iUikx
P+HeLtcsUgsp4siwArlVpRH9My2MyqoMNZtUZuV9xsEj+tkJudBvnRqrBhKb6k6b
eJt+cXyGE77BBaoeUT5UMPZ3ZFM1jfKqT7s3QagAyWv4ZBDdTEtTZCXsRBhAYeEV
jKPEwZZn+2Ky4+VX81E5U8GDwjhSHWyDvqFSJq55dKjUqn9DjTVPZZQ/GMSgxU8h
E6EQ4n73KEPnIdoKw5vw7QDz70CJjgtu3K3tXyyNbxNgUARjtOmUoHn5ckdh7kL2
dDJiZHFzQ7l1i5YrfcUep0ch3WwOpcrf2tKjrn/XX+02i2+YVBB1Ydu9EMAs6+DX
N19U82rHNM1OirzMsA3LEdhjRcF43MTH2kje+/MQO4+HoRz7cwtg0vi3jrsAJXzL
UmHhYGe4SMcXWam/qCKldYSVo9vXiLnfWNIQ1/Q1vX5zeWlyoQwMsa99h8CgqWph
zbBZAc0Bph1ZUQ7A1e9RLBgZ0YD8n+nwXwQHwLyH/tldwHFtiUjZbDOQotcoUEUw
BUvTxvwjXSBbMgD5/KonapZRrUgYahFdKghohqbXGoOfSXSEQv2tmeGRU6qmWIr8
EvjgJnISpYHgIum7OfRxFFjfh+dN7ju1rxVnRiql8MFD3whcJ38kWfmllPj7m8lY
4LejQuhgQ28pDNXeOH/O29Y6hyAoPGHCDUg3iE4bh06ZflY5bhpnnkutCeTMOOg0
qQdCxpbJ4DTg2LCZVLRrSWTpUKfAf6VwBnYIzzKy40GwB3Pz4RkyTK4D4Y0ySTfd
kTKxcaFLavgzdqcKtXti1VsWH1s11asoGhn/jqZ9gQWw35ZkyyDdCU/ZJNgsOMvo
IveX16owiCFPi3MCw/USsSM0V6NRpuJ4FMXrcU56OS9eoThZsCTD4LiC5x9xOQse
8w/ZWiq3HeV78tyZQVBbmYj8J5msf1hv++UHKALZAswyUmF2aEubcqNlPl/5bg3+
+PeylH20avyjKy3ur7VhM2SB52ddBm1+Pz5f+2rbdnhILhc9WrLEQFfzbqs+xfuT
uDp/OGwUrfOlTnwoFjNbAKVwolS37GRJh0bqinrfAiFC6/LIxVBuQMzdz5joV+M4
NMJJsPSGD3V16DYiNCVjgqWkCSVdnnWEWP491qe2XrfkTCystIYA/tcAQla2HREx
Utb0zEGEwoN/3od/z7MvcmYOhyqEyfob4WZfjpcV8hrqPrBW4WJguAaW/STpoXjJ
40SwMj9T6A+SXk618+zqdad/ioJfosEjlvvg/6xOHUsJrqXBgDSeDiIHSNvRT8t0
rjjIFOCjiIBl3ENoGhUz4P+4Z2lj2zQ8CmGOpjWesIhp6BohujtmUj2U/hUxxi4s
s/spWJAeOSvolSlzlgKwTxTeEFBzOQE3p/bczKQyJGMVGKHlQWhmx1AFxd3fZGYE
fJNRqCxYl3KviPc9iOK22Md740D/kSbXObyT1hay8w8jTIka87mpVp1RCYaDQkRr
Tea8BLqKTE+wy5gI8hRfiLhUanO5BMgJP+opfdYGMa7wa61RkN4jq+83cTFC//sp
AmuZxLDnfDAjyeGL3T3zef9rEdI5o76vV9T2wELrCVQzuhyZpB5xgg6eqt7UcK/Y
5ebXVCxOw1+Lua73N1uUxRhHGV+vNAZ8vqxa1j6KfVzmuWH1y0jgOSBXRL5O8PLe
kPfTt/juVgVO70bay60VvtqYiru1U+M/wIp66DCivJ0GehnuGFerM7w00LVk+b/G
4CVOquea6bz416asY68h0/zf2GQy67sbNr7Rdg9/koh522pRJo0YCBBzd+qG9r0i
HFr9dqDaySjhD3z6dZMEJvUvY607NH0eBFD1o3OuUWI+97HAiDcEVVZzJIxxdZ+/
g2jdlCw5G7X/SMb+mZYTva01jXcBQuWdgY5/gFH5YcQSVDrCouGa4jv5ZfCnKotV
uzvCdBSB0qAppLOr2kT//aL3zGmdT8pryB6G9pgYKUqYmC2k4ByAde8VFlTOIP0P
PYzmCs7Ip26+FIIYDnG2ItHnLz2v2d4MqKCm1pqVv+KDaQdxqF8Cvk+ElzvjkXPC
XS8t7dwGikyAKDQ7ZPWSUZ5pTNHg+Ifjz6yposdXk/BnKZkl5T5JxZh7gkgQO7z4
pNWQnFLJ/2Hr//FVpsJ2hz/cW/XOeGtwLCIAFotFNMIwLTzU+Dbi71Q99KUbgLgd
ju2PBXstAU/8yzgNyoclpF7fqtwjry6fRbyjoRjHHdfXYMgltoNT5IUFfZfYC2wf
tdTP1kfAFTT7C+MUOT0ABjV6mxPzG3RqbxquP9iiobHEO5ioqREHcldeXdQCqNsF
6y8Mhi/rElqPnELZ8IxzpzZeCtjdr1CFdHDq3Cq0/+7QAmnSy7xf4+ZmTAahUfYy
gJOIjvsAuuLQAH55YLlXrZhOARHFMX99YVuosExLA9smFcnokRAD7Thh2TnrFr0x
kpHAohw65qespTe3XAexGhH+zRq84vyqJLpioTWIbtmyjkVA5AHvnKJom8xHhVws
DYv65zt6FTYZ7c9Rttmcvz6+iIfWZzVwGfJ6bK0Z4ErgM/Yc9/FKm2x/ErVQTF3P
6BvqmHAIqgewL0kcnP4l8Yuga7fB8lTd6VJsJf4ktewAh1oi/28foHrpDA9/Fg8b
oP9LPpIwvvL9/FfTcPz0H1qHJZXo1yOA3N62Vm7JQF6wiMbH+KEyKojxmvkXsEH+
4cRifnOZWNXM3ibUuyVKNSXBCo1G2gIdCpkJRzJC6sVPabj0x5ylacuBc1l4Jjty
xIrkyKSifctD/dErLYy19ISoSE0hs6ygrsgrVvtUMgZPqWZQ8rNcabGqjL2KkKtB
W+FeugxqPR0rT2No8QYIOV9xcb/LD4PX0oXEaYQoY9ceiozbPen986fWZsrlm3sl
lfxMcqwlFC8luSUGiRSehigPvxWNqZmBWlUBxdXnKw62RLCdGzwSH5D2jJfxGS+k
TS5MbMeEUlnuiAmzwuhpRhRSNJ/vHe+PBxn70Fwz4Td7biL+sAWqm14WtKiI0Zyw
qj9ZyWLy+2hhYiDMzFHWi+2Y1z8ASxeyDhSv+TOHNuJVLNGyiWx2IU7CQDaSgDtH
Tm7G2JNqo7T3iNygrkRE24F07Tt6tRZeswCZoF6ieAFZtiZ7kdsDdPiAPnYvoZ0H
oa4t9i4KJSvRsaVTP3PUKf1C9cQ3h7OilL2fUy/5eI4saUuLaIYH0CPKMMBXiQvQ
O+YSolLp+ixMnIu3usFHPiRkzegQgpDWtHx1dBXSg6FtJgVApKiMB9AsPC9B9nZQ
yAxqdxeMKCd8iduPt9KILFfwkuO1NPL8N88lfFEqcbNPbe2IT3+XZg44RLBIvMzd
oVExc00nHkrh04SzTQQUnBeZucOF0fmNSo9AGqo71MYPb1GA2qsZlw1nMTvVJT9L
wT3U0365Zo6DMjC/s6E0MdXzP2AZXMiMmrW0C19Zl1gt6cBbUle0FvSsBfzWSCOF
mDYF7rhu8Ltdwf18ZTW9rhxIOvgL1RssMD0Umm8k+WIOSNNg6q+nSgVwLp0gsujU
l8UlaZqGTCBWq4vCHzJy2A9qMcIfoTnWAshEZ6ek+pmR5THfXYb3EkxgmoB6FMlM
sCY1/SD14UGdS2oIod3doxseuSg3u7D+hIoeYRG4Qcx8lRUXfgs5jTGMQ83WJQSs
5M0mJk3Gk1Jeu63zPOyKfHZ4SGRHL0tRx+/uz+5mbTPolgBv2eN76bDZrbdu51OE
QLjs8rwHcCvi5dm+VTuRa8tb9YLJQ2uKYri1GWlgM9zzT8TWODQ3GHTMb6nL2hj/
z623YzaESwrcSf7skmP+o+B7pBekYhj0bqPmEk7AHKeIcoaXjtxAFiaIcbmBLi+J
0VfHCQskZVS6cJNj8+Y1XDcLnv8za2TdDB/XFjjIn+Sx2WrG/lGWbKaC2GsWnlvM
ityyCj2aVve75W53bTkHhXNqnGRc5fMPXGuRz+FpVGzl8rG34Q09qDraYMqoidRW
UXE29NRFEg405yI3FF4wxvEs5sUYJDj9hf0y3pSqtC7yfuiHTxgHjmzp4ud0n+go
vXigC9LbL7a6ysyWYZ4xKR7CV0w+r0GG05Q2SIkCS3WY1K5VxB1bHevNMVl/0zs4
YmTXOSrLkPV4HKJlkbqbrQjJxBpEJ03mDimmVVKe+czI/JXweizVaQudZZ6ZFCr0
VE9XygOfcZqhc2dqU2084ga8R3Gi//2BYDRDIOcA8VVKHwX6eMPULz2fVKTI27UJ
SSrTWnJ6hrq3pc1VoKPtJjQwP8upE+c9Gy1VjJIf5mQLHT/QJDDdE2rgryocx5K7
nlIuXB18RUigNxDXKU8EC51WqJ7jMQcOhcLPGkRwP+NYuybFQ5wswTCxQYDWLpbj
I2SOel1+Ljfg/7yZrhVREtck5j+MW2pu5Y7WJPQZCKeZyUOGMlXZj3SbO+uDIdCQ
yRxt6v6P9uEWIPnOoYL5vnkbkntDqloUCnMGsuxF9hMy5gQNFNeU2N+Sn0ncrd2j
NWB9zHyi4NvdpMZYlt+7KYIOSrPjptxHNIwwHIRM9u12W8lGe5G8rZzvEai3EH8y
T5rkBDp11cH/AHZZc5psX9XEHiHoD6YWY4WN098IXsu2sWriynjY01NjWwO2sALX
4mEuXtCmzajiBddtsSKxSF3LQFNPim9kt/xrOaQL5VaK2Hw1+xmN1S2dw9RRZLns
NePALMo8EKS3iI1JLeY/IEp1chmIIWfnUYZMsNp4lsjIq428bA98yYihT/02eGdh
jOgah7Ab+L46WTLcvtTk3rW0xMrcsrKkXZ+yqfJRQ/NCS9zbCT4a3qN8lESten/M
IiPQmqmoG6whmA+UK9Nw303RDwIEtkwk14rwixoGqfyhMh92zKvShkzUkzIslr9U
b6Vhmx5hYU7ofzhvveOvahqhJaV77eN8AwcXzs7Sxx8ztUxbBnpFPYH6IA/lvG/2
iZtIkx4sHbP0ohfXHz9UHC4xsOSCGLNtEWmLXV3+rIMTzDjZlxs5bm9C2A0MbC1c
VGwyH/L71oQqEVqCMRATRBouGg3/kcjnnOhtbiadcnt4qA9yeMljsGUBTSYKJZCv
z+HN5ktiQVzQuYDoNVpe5nkJN8zw+RROxtsEdyVfkngVgM3jZjULKzx9popqpPkf
rp2G1Y81LYyOcX5D9g62wLDxwhfbj32wNhIeb6Tv+TWmMXp4ZHjXx6F6tMTTXvzi
l0NDAv6zqVyIf98hqM2jWK97equ2jnG9UozImo9q5bNnp3p+azeRr6PchE/j0ehT
4K+xqc2GWJP2w/c+2T2xlrMeowkW99mXzg/Q54wtuKZUv/Ez3XoPifCEFHzQXW3n
MXVR6FKUH8PpiCYLL5oJ2EXHYo5rBiQGSbWC5Hrb6Mij9TcmM0311tgCpiJ2QaDs
4eBVK3pb8+vt5RWZVRN7ikJhNFYEedM22WQoo2lo4oR0+aiquQRtn5/uRFm1D0Tg
ggAXSSgJ10laJhRff5j2wtTb4JI24xahu6uEV0I+znmpoIh9/LHTvNPe6ME9qDlY
Dr+ly2Bq7P5sK0lUUfsQxlYJQjR5zqYxfssa2e6NXNosnVGE8kZHGgf53KJBJos9
XbMKAZHTHS3xnaZlEqCZ1DS7uTaU9cZLWGe9SBh+heCmrCmcuBUF31wVrrAl09d8
8MHPftSfLgGMw8hQu50HVfBPEqAA5qkcVpl+QxUiGYfoW7OTxEe6bHdWut+dtkuJ
cL6TIdnVZxHtp6zl9Z2LifD4jh2tpsjPaVNjXLdoXpbYY8jyJrkaTseRVHSHHO5A
lpCeYdz9sGNBEM2t1uPc3eA9lCsPLs0Ia5oRFGZoRUyAaydE9tWbjrU97gaBgKbU
96va9kRvojLZh55UI6T8rm8QjAt7JX3GyptFVQf0KhZelwzjugr9x2qpfztMVla2
FfvxJbd0qHu2yd9G6o0Fy1vaH9JgQJoS1CbuaTuxCTLx3z8zR+0PoxYkASuD5ALm
cRscG3/QP2YmiwH4FPFGHYeGhD0bG7bnCwAkYfoaoDsGT9SDwxIIB6Jb1mkqh0nM
MNxubXSRMoBSnJbOisjaht467yi+0f0M9kkD1zp2BhFgJB/ltXbM0C5YjgNtMLya
rhDvgJJoF7ajkJj59sNSNrvtKJcxCjeXd6akd2afetACEG1Y2kuzRRwCI0PId6mm
UbBWr9J8Ndd2mzg8q+RxN8Pe5EAnTASaelfjqPGDVB23JTi49fRQnFE2j83GyK1a
2kgyXGcfU5du0nX1UqYH5uiTY5ELJWNh/edXgcsvUzLD0GcRXUK+UptpBv2G/Sml
tqoC5fJavSHgCO5q3kQWJ4CQpy/rNc1R9VB9EG5vI+B/PNTLH8mxv1VAOCqpn2Ta
WNMWqjoF1IJZxq8gVfkK194jkaFhTCtcLlz8jllx6uhpxfzcz11msQX4iSxs891I
WMLJVZrjhDFzcupVHFk+h/h05gMR/QuBKa4HNZQdP9TyfjmvS0Tv0Vlae3DLONRi
D+93gXAyy3DNDlvuuWlAeDlSuQTzBCe2TPIqYnAO8rSbXQ7Db5EOeiYvw+vc3VLT
x+p012rPqKTWBh6PpWvr6K/0LS1pt/Vf7wx97KylS168Dlo+4mHa2tMVGg553qpS
zHlsP5hbUwA/NVLXDfspttCwlaujgaOdmzaqhxL09u3F9iqHTuz45yOzmXwGQ7PI
GJ6qlnpDPHO2z6oxtLt1WxHovcFWFtMTBPJM3PR4vPbN0fC0W9CvWS7HaGHxrlBB
UO4aGypk7F2Nol+k7JSX25KS733t28shpcFG6IlNnMvblbtcDq/zbdv05Z3iDKqK
xQkZg617HMCelB3Uy6pcR9m3ilpXmyR5OyBvvuNOU3qaznbTwcTmdd3SbhyQ/K/i
GPAM+7apBNbTWsdPO0KfpZu2PEaJkn6iXhsq1jaOETR6VGzoM23p/aOM3ilR5chI
/PB4X4UIorm/0ZnnyWKigUb0Jn2W3kcf32cmpQvu9vIACsIvF4SNLS5AjJYhFsvY
r430RJTr2e8CJjcccIQN9ClzwVJcgGiq99/7oiJ+Lp9rGq3qfRFTLKQfqZLoqCRQ
WIRAdK3y5N296pyOHlcQjrar5GLtFKhCplgKBiKsSWe9jEiWQ0tS116+jXeOtRJQ
apalYM+Rko2O7iMlgfXVkUiYMCZjodOtBj3jPf5dTWoUXbl1iCoJxBznALGF9ja9
q3QZeBLfFDXz7he0E5QEOKZ2XN9/Zabxx5Z8Vz2s2vONpJoHHj9p1OvKMpX7H7Lo
V86K1sf7RP/YrR4kTm9OXU5Qyt3rkXT+8PSrT622U9zm/xsEhD3V1qFyT4JwtCw3
5WMpUNHGPC/n43ZrSDtynqVzGZFDde3ql+xtXg7uYFQE8NXzbuu1m4WVWsWAtGVY
w17CX4o5MPcYEI5nyo2EoSj4c0FjI0Nm5egxFY2oZgODjnM8C7tpK3lu9Iv4HW1l
gZ/FVpk3cOa5fg6/uGbtAwOD67aqIb/RdF/CPTIdsxh4u9I+uBXOYPtOyxouxRXn
lkcFYfx6Z18+IIalchskhChZVv7bi5X1sHygO9APB9F4p155YW7LRcGy0wxn5OeT
cLYGxFXwYSC+nJirydAJjc0o3N9ZmCk0fopP3sRfmtV3dLFPh/iLX7/U5ZJt+zMY
2bkBP44ivG5DS3RGdhTysCBC9bguaitbLl/yCm2DM+tWdMM87IUla7TuYfRjgg2J
p8W3DgFuIsHHc0h9llhHMMvpB9wYmSb9e0h0L5Ay4ZDA80uIXnbooAXbnXHqfB1F
MNEcfiHdq9Bf6dUNMDXbLfcnbY4sI+S2q15ERVqvJB10EzMkNsD42lKuJoEwPCzt
1KCbDSXshW+VdB40J20uVCEiyaZKN24UfniVFFtfEldbypTkz5cUG3l4cFjNuWFK
yEQ72Q+6EV0+cvx0yDV+NFkfzpkZDNOC7MgbLTAm1qQ91YqNDYdfz5ggGWbcNKzS
Gm08/UKsWx6KIhJ1HG4EWAPbeP/cJPQuGZaj25kwUPLFDgYae9JBcDjckN6j2W6D
NHr9pCeXQvaZYHNw7zZfMz4sAsyLq76NZTOtf1ICvUAnzil6aJjMBaXBNYQjxyB8
e+wc/UPVB/goge/OHXSWXZDLVKtrCZwclbl9ZpuHF6MOP612CzY5T/vTqalFZWFX
1jIF1iqp4mNCsThV64OKrPn48l4Z5wIEdbAPSiCqxFVNGixGOr/7FDZxUEWqtEUn
d/IwhjeGbTpZ60OldjMakGmMM7wS1j2oaDOgiP88wxPJ3QpQgfcRtchc9zyHS4l5
bdNmU0XHENaYWC1UGQUs6QMouc1AqPT9+ZNAoeWB4H0u1xr54EyUiWMVrisOgpyM
Cjda2Sru4QitiZAll9Bllhj0cWA0qDexJs6m+oJkfshgWnElrqpc3IollT6QF4wy
MlNsD1/ykMR3Gy9rp5TTTBWJvi/1nvme9Eda0m4IMd9wEIHyqJktvfREVlzHIiGx
MPdBClp4dCCa7MwsNB9vLznovdaZok8helS2aAmZMx+EfIVp8fVnstbUdnx/WstQ
ic34UZ8pFRiAhkz0OdXA2H+xNi1nMsIzcODocLLrCDK5DSPYiDWnaW9wdBjhVDqn
CZyxqdAwctoHPgS/K60JcGO7PUs+27JycQlPLs/B+cOEbOuW911RqOEkaKsJ3gSF
rsF7ZxClHkLOlL1xS66zZtAIKpExCCa9KWwkKW/wg2hV2MpxK2g/Wi4IFLgAn+fD
CiaAbdxep8VaHxP0lngkPYoyDQ0QrzJ56o+N5Tg/kor3MiH6zX2vMV1SR2u5+RPN
QtR3Vl7NbPluzWj23cGjjJFyefPkzs4YrE0SwTtvNmZK1MGy6X2mkk5HPoJ2vRnY
sgRBLxYHM0UXILqtUYdgq3t/SkLRkvRPIxIvkbtZ92lDK266pz5Aalz/c9Ot04Re
z11YXVAylftrY0pBt7u75eNfjPbTudxCXbn2v6uYVUgxOOSYCea30t+Ma4dbJYxj
/Ky7x5BLfrhnA71hB4O9HqVg6D04UWdfyNxwCuJiI4H4ujqX7oMX5Uu+2mFSGFFo
V+4o/SNuND/2mj0TJQhJhIoidybsiZh1SEy7jLMMm/m2LCmH2BLFntA9MqBQrQt0
E+P7g4n2rh4qZ9U1BmyrUyVtRGauJ/dGf8Jlxe063qvykqarbFRUJkufxYDGnE/T
PW0nFGxP+Js/1++C5jmSOIQuDwpLylX2MleMF5Iy/6BRRS3iMtEFFVg/9fOH0w1t
Hv5To3mA5vg6tgh19W9MUbGl9ySNqycG7dE3uB+7bzNAsC39bTSu9pl1P8YfcE4t
QE/2zKH2xzz3clMDc0qJTRLhFbp3YPxyghUUcktv+Ok2PJZo1BZAXwz3vklHWI36
4BW8JxHgfppr9HLvGByueGw1KjlKJxY+8iNH9pTER8E/Ka+I3EVw72rM8QGbXgcW
SXNfsQdpQ4OkxVQvtP4i/W9Kek9X/ltlNtItVzRHk1mAq2coIvzQgsz8UV6FkDe9
B7MLFxt0PCEo0WyIOu3BmwiMwtCpwxw3Fkm4hebJuIKYrCmivWVKyoBrFZNK26+/
lW/LmoQuDcHOxdw5AtHP7iey/Db0jqZH9Pa5IFxeB3jaxvESaMuHiqwFn/1bdnby
OQRP7Oo0b55Mq4drAByJh1xyGahiklzwuYua2embo1O/haHdR/k2Sk0Kz22mxEw1
Mziy9ceLKpa6Dk+vU0jT9TNovQtC9wlaLaKbTrKTbceE2lL2m2/8+5u7N0F9JsDD
+Wj+bR0Bpthyqb437p/I8Z8UQ+C7NTBliheH3A7ylgp4u03nD97qxwJ8udrEOX8U
MrFQTxesu1xzAAv6k8EbUl2jj+LmBwYrBBnZsi1hWnqL0PlE0RwAkq0LGbXvTcMS
mZEi0ZDQgRoA90fO8EzlflibDcpgkU6FRzeQiI9vgP0UQbOxhKEIK0PGzgwMZ0yL
51NiNQ/WPaKCka1kFYSV0HJb+cKGt1glbuI5tuH3Z+WbdzDFBB7FiKfQins+6yGP
Hcfeun9pWb3EPWg7ycHZWDWoIXyLiyzvoWk2uiCapeakbqGPV8aUPXHUIWhEvA6G
47zEtP8OW0AdGwY+DWE31hD+alPAy27f2xk6tu6725wAYFH8pnlc4CHIeIsCSLAa
FoNUxQmK0xu/9MrBZsr/WxKcQR/YHPhUGUgDHHnOOq+HxqZ+TmQ5ga8NetcyqK5i
GSMXwNGWVrPoshIQ4+sRFXwXjUvCxDDmGKMrbpsdy34ct5Tgd3f7dOwx22ZhBx/n
5ZgRsxe633YrG3oF7tG6qoAh4Ar3DS0xj+IHc7N+61Mnc6DER6Z1QcE+/2RLvOJS
kBMmji+5Har/0O+4MAh3RE0UZ6bMqCMpUUjnCnpz7/HX5FXzY8J4vhuuiuwjJV+A
ezuWTBdzfWw7myXDbdkbDYNPEc7ZABr9LQTKVkLvqm1lt7C879V0LWUBgwH0JVnd
xPKAkA00++dBCWqnRR96UqmQ3DgF9Paq9u35RzmZ8gCZu1sxffXAUpYwK8N23gMC
C41CUbYh4hMDB4ncZPEHOnubbOyhU9KcOyFrv62zhTfjcwp+Phx0NhB9kyUrNS4Y
jr9XN6RpjdYyorbX3FYzSwAeHiNyHDQhh0IGWoau6wS7QLokXHloHiusVNok4C2H
9usfUCtK4UUnpTgDOClfM+w9oR7ATorfnRzLD0Jo1LNGaYAtix6Tvp33VcbSK3VL
+tGOJXAeGfAui9CLoS/A7dKVqp9n5VhfcfgNQBmfg3mVEd2JMG8Fqdxi6iX/atbv
j0ONLwrNypvBLAB2hDAEkI8zuTMZL8tL65bZn7vd5itvq/k1xHLm/21fdn31d8Ow
hCX4fPwLH0mcD2kBfvrldB9uaajkOgGHGX20Q6NaBFEV8BGn0k5hR+rxnXTuAM86
E0kpouSS4/UNlUIAcDniT8/t8aMmLNwdJIWHzpZrWRJSoKNRW6ZdZby2rmIMf9TP
DOM4VKRZur0s/r3JgtQVQmqcUsfIWtqhw490W0PcT7SkAK3C7AoP7IdvDQhmK0Lu
cm2/WQrzPGXtXo4Mo4m8IiA1OROBssMI26GqGiZlYgmiT3EegMn1dYCvDvlTgYSR
WVTM2sYBm9DGB6ZR7kZGYS4UHmCCGYc4FPA5/ap47iH52gj8y3QE+9YSFl45yN4t
hl/d790hZ08yIzC6wNeCKsAcMxvajoa7dzxNrsjdLSXe8B+4qovBQuY5JOHogA0b
gQH5BjEZ/QYP6vBPlS6r+LNxKGjo3JYv3FzjnIJePjzWQF85qwVFgkxEjm5+9GkL
+zvjSGZBRY0tJUKDh1ZWJRD1EgREkR3v/j9wOD7mnEW2XnvOHoW4y2tnWmmjVA1M
3M8WKHB1NHGluENNFs59ROWVLXcMZa5joCWrAcXyf1FdZH8t8ghKCbDReHz+wzgd
4JTE2B2v3UfFkqyiUoWhhNP4evvsj49COWEdPIE1vJRFzSLva1COLQqiYOI/OQbv
btLobHiZ/ZIILH28WkM0/xYA27lAHvJAe4Hl07ySuvlUM8s++GtlSzsYjGudtlA1
lWT/VUuoeczy8TMgi7d1DMdkJCV4Y0GosJjiB0AcT4tCH2DdWxnIff1WXPrgh6iu
jfKwZgr7TGomUQMVZ5jIwcbDMU/cuf3wdx4oQisez8yP5CSg2VwfE/kwrtVY7M7r
i9u6RL7r7UL6SsnfEqq1ugVeu8g28Hza+avUbKNDfSRUr/ZjyurXAFxufbTNToxm
XaTJ1P8WwPhC0Oloj9n1WlTrEiJmF8JcV774Kr0J7BWtVYK6Ao1KrBsYZs3M4GCK
VUV2EXxvJnAU9oX72TDvWzp87WePXLtdGTdWlniFw2S+i3AfdUzEHsQ4wuo2o8bw
pf6m/Yxz8WU0yBiH3raqdbiPsZLsLw066lAffKDOBN6R+9b0Whw8+btB9dGIDQ6F
8TqA+QxqQfBUMkD/o8BoIenGTRMqUaKCBLogBja1uQV0plctclEO44QJxR+9z76A
Ls2pO5JSGgCSiMP3SXc62bXhwsEMkO18tLXtIvcrN45NzY6mrMvmDtwLC9LlHJMm
ZEXbi7Wf493EDSxja1XzivqzqvrT614W0L8d3CB/FG6HkYb5zQ2ZtbTY7DVhr4ip
ipTAt9DIW+wME7g5O7sB00VGN8PtVcnhqBL14i/cgPkNZpJgYO0TsuhXRK7SE7dm
MAh1sdY7n4LJKjKG1m6zFHqG/u5F6NFjAKDb7IxiesN/n2eKBf1gt96vkJJUt4Pg
5RsYTGURPuBFKPk0zDYJNiKohETLW4e5Xv8PsfqeTl1634c7FoYHouE5+X6RikG2
rZ6hlXZIKRtMsNqx8PpjCNsnfZ7i3V2HqDZp1rCFnMkZZLFtmoXLwRfpgEDccdWu
x+jlK0YCxs8tL2LTlZjpmmMxqDNEe3tuMF06KSKoRFuXlHow89ADtqnCzxz18lXy
q+1WSQQxrMICCW4imLI57N1NLS3XUgrkaruie23FJKwj6na3Ya9uw/Y+W0UHe7cc
oZkTXrYGnl1fDIiEkByM9H/B5OU3JLZWjsYbfJdSYaYNlNY14QB8CJY+uWGC4s/Q
jYirIMyZsmAfB2uJrjVr3TdbeFiyvWBpyp4fx3v7c3V6akIfSolmadgxnR+MN6zh
IgG8lFbHVBqGV2HeJlNNpQWodiT8m9fLe1g4ZQn5KqFb9MKrVlQGD+V93Sxexk5y
LI/efEVLiXOVoLB9eIu9cyvoYRZQO6SYOLC3ZhdKJv1ZbDOdzi9/LNW9zZDEVwfS
GcNFl/B83iYOow9BGKBN4lWJv9zxmVpcMwaN0GF+I0zdYJkSvFBj5Zsswy8HW5Ou
aKMJN3NjipxYrPRyahlLh/E7JTq2WflZO+tj1aAXPqAbk71zQdImDy1iP2jxEGh8
xIbZsf3apnlM46xmLGUgaYJ+/gxj9UGAwjXDNwEd1QHrWnxuRFTIkHOeEtvIMgcz
0SI+Fn6wOczttuajMes4dZnz5l9iDcXSjIKFNNKmIXymXbHRv3hrNMUM3djSSf3F
6ObaumPjfgMX1f6yiTm7ejlHzz6IKMdA0O9PkD0lTBwHy3qNUd72rFO4DDNj37jh
j8S0/umYWd6xwFJi4DJTZMxRPAFcl1+wryimFoVs+gNYQnWA+KS1jK46zJXbdrv5
xCoivLhx3DQJQ0YyWVyGTfIGseo3zpAliPlG7G6JKKLVawKeloraQWyQR1DGdPyU
0oaIza8MScyHmKRYwk6HJALzx77mNSYZKDbst39SPcykwrTnBNjIuZ3flIrT7Tm2
q/1XtPELtxAvpxHmr2WxMvxDU9n8g9tgzef2+b77fh5kPefQhxqDevOq9zzOZxas
Qwg+fwGC+6VEIU0ukiAB7lVZ6438WmGHRaNz18cEnuDkVKzPRcwoHAWpgWg2oTeu
2VNs3+oLTJIap1LaNk1PLm6hSKeDXyUODm4lRzw4Y86x7Dk8l5JOfXlC7vxnWEVK
nPxNqGRi1G/38ZJimp5o9nXIVVX4kLy+IddTeV8EcOI253GxvJlQ99cQXDFPbmi4
0nr4A2UGrUcNNGkArtgJIPGH4V9YSH6HYQiybz1QlJysYqTp1YvytB5RlkkOg7tF
K7UgaosVDVE4FVbQTDaFabGaMNv6v/iF73t22jy+qL9BS8tqEBbiQlP7RG3eUnAh
7enKG/0mRbfOkpoc4+RFWAafeCMqibyZ7QqI7cRKNEO12yAABocjh7CedEgUIUvB
tLQ4ekYt93uBaUbom20TA/RZeWGRRp2SRSj6h/5zkuzy5OwTLIj2Hxba4PQFvBzM
laHDbkNX0Dqv5gNcAlkcdVI/BKldr78F20PP+AujZwsQZFeAJ3IrbqgJZDwEggip
3jSmjEN2qEnj+Xbux3VOh0+xcsHF8yDSLCqMJ032ujjiUegcufX+SQ1x2zqSKjTp
ZOz2VTmufJgp6VfxKkVDn/PR95nrhtXqWAds7YWuB0GTwpocpKQ2svHF/rMo2QFj
PWH7/84n2bX6vQyB0yNtAzJswadn+gpDJWOFccRzOZ0efp6U1GHD6tUPEDlydLHl
BM2fUtcN+m5Hw08gYUN9HFg9MapltUe5qk6fPIQMsZVEAEnnAX7wU7l0zCgKQmCe
AhO4B0MUE1paUuNfYiihaTfdqJ5mUgKMGI+Kt0xD97WdmFnOFei7gOmTKs5KNrIw
bDqwjb2DlhQK9Gq1HJFAv+03znqsORXkqn6K0hHLBHxQiYwQtsomP0Tn2LOf2ryJ
OggDQ3YwcJEwdi+bj1UuCihXwDXZ5BwsHltwXp46cntuwIZo0NEWtyBuQfPUEDNn
bGtwN4CHbAohc/oH9GeO79txZINJ6spXjZ6QtuZjgtPRqyH6OpY398vDlB2CS0XD
JdnDPplwia9LIWkk1OUaPoyUdunF+JY40oga+hvber+L8JZFo7rySQJUK7tF9Dvs
mI9wWAJGt7BMz36hf/9JhgQ9lTOn1LofFUf5T3v4mOP7oRWncNrjU2fOCnbMTPL5
dnZi4EUeF7x1sOcfrptvO9YcfHanoLAlDaSVEYRuuKxaqFJTWHGMDLDn4ee+BrhZ
BCHyGq6TG/2Ci5qbhDN6eZZRzcUxdgWpEt4YwbDtwY0p7LBQ/AAm7MpRYY5ioWpT
/Htze4X+vLJdKlBZrGXFeDhV8VKFVf3B0pEmEuAo0AXNgB5reWaNgOROEEGuWEOd
zJEkBJ/9vyu8Rl0ITPz7cUM4sSEkryGfiu9SOoLq5PXRBVxFEeMsTWmYxZEwndzd
ufLqslOF0o8byPIsujhefWljP0pqPOrm5a+hfeCVzO5OSYiDUZVHnwWnI6H7nHH3
zDuBnabo0luhf8p5mc65VZSuoRspihfeTt+hDfo7Es6B9EHNJCQT+dTjEX+gdqc+
jw3vyHEIR7cv/hHXxS7azyncCPTXRx/k9RrziGC5vERN8VBaYsjAXDscvQs5QvZB
/ncGWZdZDYlkhNgqcUaKowO4FjICHmpoI3qnYE/1K6/C0g/5rd4BepkhhvWNg0q1
2/H83O43/CgBsQj3a7xJ+euNnOGVm96dpyb48zfvBfOtVKmahLTiOzXQyBAAwabf
IMA102klBQI6UhHK+32kp+x7xe+1HAt1yT5xppRBwOQs3vpEB001b9g7QLNoB6kt
8Fm4iEaH5PLE90waMOsIaTSdefJVIbB4+6UH1+eeA99yYJ3kIQHTbqfT+nu8xu3M
VmKanA1cR7kHU7u9kmPYzmQpVBsk3+78PuvqwdiW37FwcIO5ThMCG2mki2HI2hdU
IszWXth/i5Pfdos0sjFzJtHDijFyJF65XrqY7t817dUYakT67quJjVdAq7Avj6C+
5CzF7Okcq58ggXGfAqzrtWxUzho4b0NL/w4Q22ufIh2qRGIpGNIOjDxOLjYHNmHE
+kmctIKuBBzjSvi/8dED2+1MRA7lZQ2uRG7lfy8IVvBwXRqWabjye1wM6s7S/jq7
74oZdfHqFQQkPMLU8YSpicFYouxE8lRZan/CAmAJrsx3wOlkqliE2Ck/Q8I/fWKs
2/gccWujGAPDY5CAaCwgIyGMU33tsmDHP8OYwdZqiUepQY1nVXSBNesyLhtmGbA+
pZu0RyBnRD74XDvihKzeoDdVWY8Np34NdCBbW21pvrKo7A3UfJlhQOHZASoWqpve
p7S5ZeSmxq7p+ZLiQVpcdLR0L16NK2or5rjH6Z5v9LsuJ0FxFYgDLVoqfvyCp6cY
+vTPVbtq+Ixi8Oa0hg7CqCYxhRlYbzHeoGEFCWRsrkaKCSwTvCfcWnGFSwyCZ3pV
3xpfMuNIRPZj1mUJvY6sphjsCLe12vLIb+exwkibuBFhAh6YFUf5HNju9QNLMMbn
rxXIV1zzZ/wqlLWmXz3qdZdwdLbYQ8c/7TDHxOMMpCk6wDsoexH+G3lAQnOnQJzb
EjBK7c1TdQ+fQ8IHDBJwVrxRM3yJKQvjjm/zuzwORs2O6hs91nzQNM66tx4ZiXSu
zGTVrar+jlzD1yoKrVlpdFgcRgPsA9vGev5vXheGyJRlpWnSlBP7lfA3bO6laZRQ
beuzFIpenfVclKa2eyGOEqKSNcnnzT7A7MtDz2h9pIpaYMozL48WOt2pwk1oxlwM
09HRJA66B+B2YlVZZAjnjSxhzoOR/mF/5nKRSNvVhmZq/YQxr+Ii1ecgsnZ/U4hB
T/8XIKCT8S1pjBUBO/8oxXRJm6NQYwkUgE+D4DHJwCcBOZiUNq4wz7AZTwsae9Dh
gFkyIH/kyZaa3EoaDkvEqvrHJiH1RU31oTxhiZduwCTZU3ekQS5GjbqldFt5Xald
E2V8YymiwCqlV2B0dvftW2JBtowgezCMPa9PP92yuTnzHcmEtlOgj2ASM7e5/fBo
DH3+hMcbSX9omlnE47bJiBMVCCB7+pP2u/BX1Lr2MaISpRPe3CTnLFlgp272ysP6
nlyt2Rux9v0AcgKzmRp06b1EmgXmj+U+Rb5SSOyl3sZi8m1EziCOsgAcQXbtHebL
2+EBjx+lBEHpe8ONTIRK823BEmt3MddVzTz2vEVkwgUy1zQEBuGuwmM83Ej4967s
HSqouC+hi1ADx+TGLOMhPFpnz1lNmJgbyLW33PVMaEOhjfF5UbMHnDqHPeBut+5N
qoN9GYQFNLdtldP/ADIPQtcbdwcd36pauONpQq4P1LcXg/HCqq31/AAPWQrR37gH
DqhVpUZVCq8sQ+14MNw4l/6zjT9/XW2dhzvI6N/OYhLGHxs3Q/SjhDlt6wIu5B51
PyhLDoWQdnotXHyfO1iWjCPTIAOF4ViZGG0JCVwA3dyXSOouIoM5VFpeNkB+aJMQ
3xdiRLTEMTlYZuHQYgQr7PrEXNWZr6RynNv3VEcSpp5IYngfhel9pCXFOgE+me9d
7O1Dbxu1a7X8KJaFq89En170p5aqRmsUzqvAsKlKmAgF/tLdFvEPnzw1IhEMpM89
OZ+/bzqZxARz6Wf3X4o9OPdMDSAX1fenrmKMSOxeLcPMvynqbncA4r0+JIzMFaxq
wP21UkDyg/JgXJrhZCztrYU1fXr0DRzZJSXWYbYBM5Ip9ij5n/6mQ2/YC31X8fBw
Ljsc4Y3odGzTocDqw0XSwF8dxOdGW7waGo2DYRuGa6VJTy5UhtWfDmQROmoJkgdb
9j02ebWUyxB4qNwXqTdjldPZtB0ydG+HXWUmelmBw9bYJsa2xZUVEcY+gEyg0hKN
hOXwNLkEdQoIhPaXKDPf1CqzMADKNTh2ENUtQgHBcQexAgdGnLhHaTOvT8dTerZi
MlyRj7PohRwpZ1W8TIBU532qP7Y1N+lR5z8FiudaZc8oDiU3DHwDUL2653HqOiX0
FBdDHVuVlhdHcErVZPe77ki2cXGnCh7LY4F+HnHCu6Oo/o3+X9/BdWdqotk5kFo6
8f7GPK3LsDByla00bDl4kGisXriMbMTOsgW5NGESlPSgkaT8OYp4Lu0nHD0gzSOG
97Yf8uQfl+I52t5520OlNfL8wUbEAb0sOspDnTHYrSPRnXaYWUq8jZ6xQxLgwmXv
AxQy3DeXL1u7+SG+PU2QgkcsCa2MJq0pExey0vyEhtWQ7COwWWXlJQcVnp3X3xZt
NjfvAP7jw/McqGzEh//HpHPvr94rcokOFB++BMcyYbm4PcoSu2Ovz27aZrre9tLb
ComLyTZYMGvv0c6Ps7/N6V3H+HRFgMAl027FKEQA+UNlGAbBxhEhLT41iZqonof1
MdKWoHBOEDhEEYp9A8zBW7Drk8XNG+CrLtqeiCJ/iWF8F7q8zutadK4KIfEu1bkv
nEFNFdihigZpLYZNZXSW1fOysh8KhD4mITWFpcPLNiIzJljzj8YtI9yrAaXEXOl/
2P3vZE1YWUEWbiXr0FyXdDD5QoVga7ec8gQ/LKkbu3D2vWr/Cd2pw73IfWcBdvEt
7Zv38kQbKCcnNSIt6HLW9FafaJi3x4vtYO4ZvN/xxqn4nH+f8ZGKGQUtdvFucceC
M3/YNejlRusr5ksr10RVSCRfiJuwbMQyHPYLuoMZG+cTQLsAElQeB9vFJzcHHqNP
GS+5LSM7Uo7AnuKjd3dOZRYqgmkNZOnFHF2cntQZHgFnJbh7XLXqtIR2a82AsEuV
gT75uDQEt3Gs30L/8C1mgmGaUbN65uN6HypNawFlzSY5N/5KEjIOwYXAwREP0nbO
6J7yJmIYUeRNO4VdJ/MmSF9yG5yQfFg4plNXRwJTwcLAPYwYqdkc1c3rGuJil1xh
qh0m/jHWu/3G/9zyz3yUPgbrdWryVS2nDc3A1Oe0t/0vdP34plRpfaPMmyj0eGIB
TdFy4cczoZbtxJTlg9AlcaCrr8/1XdeQszyhk7EW5G6f39/I4M1/joMllICcH6v+
ORJT7j4ZC/fZAchq0JONHl+Fka7KyBqh4KRjeCYO8VMHRQ9Zvrs6X4hhYa7bMBzQ
QW/83nRP5GoqF+6bGKoozlw7Wh9byWZfXMGksZCbcKQShZEzLurQJptgmTgy1Qvw
F4TSDpHOgaOa/1A8pIl7UuTi3Bkg2KmREVJgy69Dn6fteiCTIeqm/cZyiOJCOx7s
GSjnl5GQWnFtOLcucNz/KrffL6tOmQpvkRswKSQanuMdwIV2lCd+2eLvIIgG/GVD
Hy1/C1xwR641iF+k2wLqqiSBu/lnx1GgeAqOsl+/pXmz3uarGXQADYvtfbQHoh8E
coOQDT9MEBvrJrtVdZHX+EEt6V5yA7zLuvXt5CliiIlmMarQk6668T22iqt0gD74
8O4VYVXHBTiJ2gogvWkLgnXlJXfrJ8In4NJcUrx+Ol/pAwXMv2agLHZCgJ8QTwdl
ENWKB9Kz3MCD4Sth1nPUMP1WmLe62TWVV8CU4t/ZqmpWBrwzqmfsvujrFKv+kaaZ
lyDlDr9J0E8G3bpYdlfhzub92BXwANIRJ2KYouea0CABX73FNLk9eYCiUpNHfUke
6Wso433pE5xxkeMw/uOA9saPCziJA3BIYl0eDmIlA48tHCuMrEnTIP/n30qq45k3
/0gznuGDWhgh/XmeOoXuMqGr/Q6ohqKH7HMPlfW4vpFQVIkLf9A4Y3Xa8AM1odHE
QVAh5TwNKAz5tG4H+mtHXpvVbFUpL3Fx9+ZpedYuJQK2XDHa5FpiOtFbqV/B2QBV
FCCYMVvBdMGC9iTN4EpFgw99HeFYJhdbwx+qYf1r0sVD4GKmIT+S19awIYJ4c5XH
Uy6kqICQ09tD6B2hqN1t9CY8fhzdYnh/Q7ZJrHJQSyl9+OZydqY7n1E9OPLK4YMo
k7vQus7gm2DWgOFVgyCCAlzy/Qix7Wj7qSkerUzbesKUR39dK/wl8ny/7m+h6EsO
8hSB+4iTOVhEDKaDHNkTCPRS5f1ESzr8qEdAZ7z3VDyG0ng2zEh0w5q8g5k6O94n
K9KrwmNPI/1yg369LsKDgr/nPLLg+uuVeVMlj0Dh2M0DdPLAfBZHK2+BFEpgTO20
hOPQkkToxixZ+fUPzNmzFo2Ix4eoM0ke1FDHX19LBfIvRH0Pdz5QHVgYXlFpZbCq
xCjG2Z4hB+BhzNuaIyayC0X+NasQBFtevbf/Wa5+wqbrChzOoQBS0IG/3PKhq/0i
7uo1sXv789kzd1iz4vK1XZLKx/jz6joz4+W6OJdjtoMjYHUwl4jOpCa223toX2X1
a/h/x+MeSOTme63COZXdmFpvmqYyd9CpLl9AH1pqiZRYHw/tCrb4OjJLHr2aghTf
tv/cVF9QSZ9Clvd3B5Mqy6Zas/7QWZC9KmnKbu8j8oN5qISGK2BbMB8P99+mAYDY
iceVbYo7K0w2NMGqCpl410R7mEYe3jszhoAKfXnNtWnPM3aHvMyYbIO9ZCGcFu/N
MgGTLP9i6bUlw7Ln/9iveVZtvDEC7skYUAhUwCdGsz22A5V7JOTdKUmPDq3R3oLj
5/zGZh3xJATAiZfHJ/nwe0I5CFEuIEYqtjNSUEJac4HvRJID+I7EjdurdPHCRzZI
h9Au9/DQEPsmALs2zOLwWiszukWcqdiFcP0zIOKtXA3wpPmP6aOssIN5RTknAZLF
yc/fehFdA+CDVyJodT7jIsLDDJr+Qdf+CYTr3X+tvo6Ffchv6JzAY89jo/PhdMlc
ykOMWYLhcxz02A2iFQ+jM/8zBrZP0CYLEymoOiojoqKmtIpeawMqH6CD9OwoDBIR
DEt7ciIiPX6CeOqQf5gFFXmKW1bk8BMH3w5GK+2j+Lc2nn11rb2Cpza/J6WL7XkO
Y8vBlfAkXh7UkXwQru1n8yWc4m9J1ASZ7Vo30XeSYFsvzAXJYVshXK+LaIz0ku6i
pfmkLSKYI6NBjgMFZuWDfn66w/F+0emv3qv0ui2Wsjej+lkhGOGXUxZQTk7ObCdv
Poxg9EhGjlcm0RiB45Oz6fkty19f2v3R0y+esEPnVBVgPwmToQUWMwgeJVK2dQb8
QWlJdEOpWkXw/b+FdUNc8P10i/Vg1fHid6I0CcMIlux39RM6jPt6ZE9JCMHzDNBC
Kyl6kWVGLlS/TR+o6KkAYvGe0Ft4AKyH2gDkDuvxnY76NbcMwPRc2P3Fn72hqH/N
hhRPLkn76nQjSU+fvoM3MsvSgYgoVc77/+ncvvNGKj63MmebRIx7yCIcXuWhSeBN
Mxuup2umM7jf6NZ2Fkp+oE35ZGqMT1K41C0P08PGRatL6e5wXm5c6k1Y7DujKdBQ
YBb51vIIj7yOBKjsfPyrOxu/XCN2HcrnSMxHzxpL2hj0hlUtTOzO1OrcbORWarjZ
y54IS81yky8AxwBlCXzEvnCIZFLklXhmxWRkAknVThUkJ/OitSMyo1WTtWalzyqb
1KxX+JYwQkpQON9yMCnWd6xtvllUUWuTD0E97mx/RAme7lg/qMIefrXOkoPTJWRD
XKVbm3uBwoImAys7S3J2So4iXwPZjmAAXmlI+oVekOFwomfkOMFYsVm51aCUT/eO
P8bde/fJoRqMIHG+Srb4nwmDahyuZn8hD4KSdLvmUk4+udwN8sJF1IZ8ejXtJlIi
XdFzuNpDyf7HVIE1wWtj6aqpMRzgCFZKlb0Mn+6D3DDShKAGGS83mNyHsQzBKivp
7+YFwr1D1VflkJRyEGCznizcy5at8SyqpPKJFSqBk3lyovDBX5kJmdvbG7ZxBbQJ
n3tPW1qO4m0aufJLb3icuyOOmvF3bTXMCbhA14epCH6e2szRKvQe6GiOpZRdcGXu
napOTFA5+2q5cx+cexFc8GQ9U+NT+sdg0Tpcx9rlw0oYnlsulVjKcu9PrkadSQth
+DNCK/rXpkvFWg6hE+/Hw4MKqrgEvEMjXyIBpHbStdg/b/pi18toM3wt/GUoZd6g
LKYP9YYBm+8r9TXkgLczlNTZeUWKlz7MIfq9k9jav5l2QJ9SXyNCRp9YVCcSL/mj
L0nN1o8T4Ku6d2ANTk1hS8nj5hOMf7x6UkrGZ2NecKHL4LSHtbjPSxPrcpBePArS
wyp4zd/7jBbneL/qp66HWRtZVTK/OhLi9KGVccJ4JzXNmNlC69om4EpMaM3xIDSG
pae+Z4I350cSNpy4MfhkDAr1BMwAEv4TDXrBIpXYsfnXN9Qg4Tvp9pndvKL2IjdO
hy4UgRKDCwFXjvmUKbD/SPt6t8HWuXA/xHk9bJhJ8Pac0TqkVWrA/jaXNUU/0kq5
dMfbcm8JJIbPgeX4aNwxQKs2oVQgkwTL31WDHd+SAj3GsCIUwMmTMmk92bDnibXa
ikOkay/1vJFaEjzPWMaO0zrTREPatgcjjJCBg+4v0YKBqrfEDFgBgmbPJiBVui/Q
fHI1fBoBdolRrOzUrTt6sSRpqxhJD2VS8sF0umjaYQxkXjHbgCO+2NN1I5KvPjO/
mGjRBY6ZuFoCvOi5V2dhGi8L/VxL/sIy28mc9L2Tov1aQegFR8Nv/n/skbmWPMRL
ziZ2cExighWWcRz1jLRv2A6T4AxbteNezhtUAzIFIpVeUztdWjwNkaLfvYUx68wu
T8s8lS8SNs38jCHYtbOxFTwjnBShpBxdw9gfAP2TrLDJiqf/QEBq+FFQGCQqo3od
oRSGE2QSq2pVqjMz7G5qI3rOUnVd25cdqCk2m0CexG3ervOOB5pxyaqtXkl9iZC/
jyOohR0I2SO9c9M69mEhRiM9Ud371kTMYLTsO9aW0ok5Ybup85X+fPSLH0tXG4oC
i4SJgKvyebSSYr5VO0cSXdraOUoA8sMJe8IacDI3C8LvMYWXvxEhWZFQ7KFAd893
PwROmWG+38fdaGkPVbcNxxSSCi/M9eANhlQzrvxDrL16wwvkIPLy1tuvNQd+g6GW
O/DEJT2F6YiNfve9iGmPOWClSGvnxza+XQwKn9BvbiLzT8TFNChzzSSCnkh3tKTV
bu6X+r9IFq8NHXFU7AZk3gDz+sUDudnI798e3QQ9CHNqiu2bLFc18pDKfSCbE8BB
AASJiNsS07FKmCtIto+OwB9zMGX1CJwEZ1bA8wWkrKGcYmgUwiQ4txbB/qJq1GB6
enNFYQDEFMxlstP2LPwMDPEtXozvXpe1tPhPDcQzZuYNH6I32cC+WWdWRRu8oA76
HgYW2sfFrckCwCHunjNuikaj44E2GNiRcynqyvcxQ17LyKg6Aenxi+e5VdswtpkM
mSFuWLOrVAFlsDzhUwC7OTfe6Lfcy7PwknzXhfbhvWiYElqCrk1jWRWfeE4Gd7Cb
v61sI4e5qAM300+ZkVOLfXDAkXVabV/Rym4AkseI7GGYeFL5/TKmRudqBFcL1IxI
2xPQfDO609cKQR6RdcpIAlY/lccWze/e3q8ejUkID35pWICUed89U6qX621Xop8r
TI2b05fq4+lvOC69DunGGvV9LbMkK+1bnE6Awm2BqoIiCOnimPvu/8LXGh8IDcPe
5kKclnRtMaHMuJiO1XzWJkvN1rZcLzdwRHn9mXICAG2gs++N9oGgGE0IA+76TySa
Z1BsLzZUTBNtMYHYfybmrIIAjVFmqyyJaX9Mp4fTHPKCByh9tVuhJ+inWWwjjeyC
R/5tvItXybC9hNoJjUiJKr1vzlp2YckWwCfO9zMKelPu917IjKl5zzwsVoa+oFnB
anXmkOO9rq9iWWl2HzYht4q65li9OJNr0gF5gsbA3TY2qKU8jAaXZzvFj73d35P/
BXUcQu37tRPyv2ZzQhz/YhnjzZImgP5Q/79Xep2I0GbK5z4EcIWL+Py72OJPVm72
z25HGBFsVWdoSvfjOWQKZ0/cN+ctpmctgs8pm5jsgDNcuYfA/D31YIs+wS02zuFV
jojlfyt6xD2fTcMzFezZ+uCdqCCvk9AuBwOeFcNiBPAm7LoGV293OFXH946wZ9r8
Gnii/afRKZNwTCEQP3qLWC6IkAoJIj7AqcU0PB8LGVLf95dK84gZHJAN8OAtMX++
ziYTFVijmlI+OKcz2IsXfEEtitYmTnxRFWjalX3DOfwQo42/g7fnExNr3DyW5/bs
K/FI7/Ut682fZvqA+04wl8X163423F47TRldEzyqitGbggZb5pSlbOt/4SMmBdy8
gwJL87vgLdqDg5HFJ0VNo/j8dETRqjU+u+pxC9X6J9/mHsnLI6nKuGKCku+clHWu
bmdYvydDxyA6qw2mp/NMu59mnzxRZKtDr+03eYy+sop6p7dHrDcYJEnDBr+xBOat
892CBuEt2xEFrHinh8KczJZcRZ++qvugvoomEA7yxre+ngRNDbsx+F+POl+VrQ0b
DDwB7xje4wVOnbEu48UsN1e1tXORonj4h1zXpjnEmFVK0XKaQBdRYZ7UCYqwggnV
YqldNrFrB4mSNG7hH0rSNwQExofNLRJOumuvA890d0zdYVk9Ze5cxd79MQpmYsER
MEmFcUu8lB6OpFJIWHbSAC+L/f7F2rjXOIoKNp0fanH5eS3uh7KVyMoDwwfKoWC3
Ri3axdgBQZEWsK5YHcWcqwe1Rr60LCXQ+4PDPczMAND8YnJ1q0LNx6iOWW/ljsMB
tkIHGkcdtn8jKa8A0Gx5hXUfflVSPf1YLCfBKjPCiS6ZJv6aiuYGXbp5N9Kq3Ymm
YVkyo5M5ph/86P/hW4/g4rnshB75E4b4H408d6jtuAFVGD2nnyfzkcLJ1BzaXHH5
mDZIY8u68wsXzqPupgFWhA7ZGPhQLV+gRucDi2fObN0B7NL++281ctmS16koQVfE
cvR7eZLPRnnfWMlKaTve2iBYfJaKbTDWUovNhcI9Vsv7d8essMpit0MdgkJspJ1J
dnU4qShUtqdmaikYpB3Aa8WH5XWHhFWWmuDi5mCb6N5Bq53/EhTrbDszvTwxS2kC
XhU09f7DO28kxwmcWEr72on6tS39RhIT4y0//n+DVVNAZIv7Q5/huMpxMxZEaFhU
/4PSMeg4dmAuVy/c+pc41apBsoz8r5aISBmFDETTgNoUbX1oSPSqpszJLXnFLSvS
xfhgV+WnogLPKEkfJYxW3hgRy3D2cn4gvTxkAE5Hx8GvHtp2CQrXJ9Z4pPIUUNJZ
XJGkjGyyiDopC6uXf8NRxenxDNBX5Yj5TnXSdcMACDVqIxC4bQtqXz+8NiDBBH5D
Rk+SmBLppshgc1MMzOpVBOf5HO68TKE1b0iHwEL75/Q+SRt7AP4+DPEoVa6ClC9Q
IzarhZ4C5AmySbi2VZ3yxI2QC+ZeJ20K23Wszr8zmTVnP83jogdljB70Nl5LOnfV
smCbE+wheQpZOiK2/9aD8bKRVPnz2BecRAT+qwX7hmEpKyeheRrSNfh8BfFJKfRP
QBLw14a+k/DUIOhTugyZukCrURy2BL2ku/nnYyThdKG4MHMAVMRwuM9R1lkGzAcz
MRmt//Y1LKNa1LITnek6Kz4jFzwz/ig1Xjg8mUOd3QFp5UvNgJmJzp7FGDTmH9YA
MUfmZEQYSNVYBsBZEkAVjsdBBaYuRqcx6h5rYThUQuUoYxBKaCjGlWWGaBCG97a2
CXerDZ7TWBRLqvdSZbjk6kfMvT/v9pU7Iq35t7Zxrsdy8RwVsTgphiyxIZSZ0UuK
bcquz53gFzPqFfYqEif3LiNzn/5FvQwP+4lyYIXm6Ob/IVKJTZHoMerDAFDLAyMf
zMj0eYYPaCMldsUWEtCFT0YgYb2QBQKDGw8cs1g/2phvvCtS2vvCRlD7zxE3p/K/
gaNeV/UNRoYjHrTqXkLq6ODIFClseYd0oombihAqV+wJIJIhWiFxHpZY5Tj62dAK
0vk4nbo+h1F6+0935uykUGd+D6UNsthL3/Edd4jFgx+neSoDWWhRT4guibZT45sE
hBm6o8VrdhirPaO2y0sEM5q770WSxrpCOLD1IFnHnEKiubiWvMlwzPSB4G7cWPyj
IUsjS1uvX47731TX4sFEkARdWq1pdi1YVB0Ni1jDKn9Zm6QccmZAxZZIWSYdPYx5
DHOfHTCGu13gAhfn3kwBt12Og2714qANGyNEmIDjWc6oOEWxev10x8EM7TbJ5O9y
q5ZFSPDOYwrNzfQ4qrYk+CiCJMl/8RTtBlwT+uK8tiPn7p4KmtLIcBOTcUjRRcJI
cxEn6IQCcYTHcAb+DgZdWCEFRx4Xix7RUPz25Codwl3GbqraZHwzTylVDTh4J8Fz
yb2Pg1+WaoJkP3P+cRKK6brKgbhHlJaM3J1GX3mlsiV/Hs9bBNxQh2yh2Y19MRWb
IBXWshY1u5gnrlt/yY/oCzXCLA45gXG9vIxpbnK4C1mueradjiuJmDM9mHxG3xxz
/DhQotd3XO0YY1uhQnEfGGu4KN69BaVkcd+430G++XDJLn/gMHDOG3ufhrMaGGVd
ggKeV3dHZhcwu90lWWls8MCBJKQiRLbugiQ+42xAjKdBBlYGSRysVmQgVsK/aR8e
Q3OCtXLVbFKeqBsg8SFk3bWyKi08mbWXBWBRkAH3GADvTYEE0ksuXo4bWQ9pvX/A
x4uDbYrUNxt5la4cb7hLvu8uR8tmSkI6hXGuuEQROeYoNxCCByw/PU9fieRf3m0k
+tcv5jzKBRrW5FdRRWe9UuMkQNf9m9kNMVZd9b+M9v8TXv6MG7yrylUjbOr0I250
UglzAHG8+6snmLL1yAm3qkJtw4i8xRb9SjSz8Lxrp9YMSqh0G4hHI45fZdkXA3Jv
4Glxc2CoUMnj+0jWDsCJ0N77JB0N4/KiAj/cvx4XZBj4wtzP0W6UREe50tufIvzb
38OO/UxWjNAfyGn/CIxlEvf8kK9E06/vh6U3IzYs739dtxi8rE/p0EAs84WHq6cF
1dZDPNP2ICPoGNJroPNWb1oCY5HexiLA/+daw+xvXgFIzKojZySVnyrxs9pWWY5L
1q9asopRm77m93DbSR2/L/Q/gsgpTWaujXzb0rxwYydFe48C3gD0SBBovXJEmAco
Q4nfQVYNw0gwlk62gIPlnIAsuU44oAej5QguuJHM/eZNKFw0G0EALl8hCGfdlY6j
OWL65LDMWugI3gx/+TtbHJJDNsA7taMrnpXY1uon9uYjGWSyhmw44guz3EYB6mgO
K8ZlKjJHy11kto7pzbf1RFbNNc1ewLmbQbK8PzcF8CwNptM6m/FXPR1D0nzu5Mo+
ZvVHBeykq1VYK/7A5fuRkukMzDaifmT4EQ8H80PEu+y44wy9O0Do4Fojuj2ZRWVV
ktVRGXy/URwxSdi31IKi0nA/Ay/Vgx4rEMyCGTDGN4D3yVDc+WPqOdQgz0WBpFx5
FWfRO04KGInCqzZKdfGX4PtEn9Rcyj4KWrZ0TNJXd374WX4iIbPz+Bx+2aNQzJYg
mlAoA9poxuGwNbJamp7dASelN+mYHmn11Rk8cLLEcez93/u8hdwCXYotBlloyGat
D3pUo9qprxJyEzgIsEHYD1mEF1Mxf/P4zVQvfa0UKN2oyJCdNrZM01ZSmQ2hkAep
LtwsnleCFhyVA6BZzeW2osv39Cq+xxi+pvhSga66n22X29Kxsro6Zrl3+BiaUoOL
5FlsGS1skj4gQQeFOVHvfnhw76tX2iAX/SrWWnlOAndgPGWBBjDxEL6TDmEcLV4E
mAWzt6QZlGM4/ZwwkCbIHgoA5DDpYYw/yBl29jqzvzOEpogRv0y50uvRxM4PBI4u
jc1w5JLjfOSQUomVo6EZryXwn0jA5fEY+6JVAdtW7cNym3Mf2IWmW+mOjQ7LHnaQ
YM+Sa/RmVlEuh0uBPUI6Ry1yLGpOvZMHDGSSNS4/ozZerZVKrQB6RCsVjRulJM4y
qySBN6F3B4AZ6h4NQnlB2A54la9PbSPLZGDSG7ZGcR9LqAIVUY6sEtThtnGB9/EN
jqDRDWUBZ2+o9lCDcStS5B8l9CekYGaC9FZtMamUsymdZrCzPWBSXiZr+WULBYwz
UWClJ7q3uNLBuKi5RbU+LZR6y2eZ2ik/Q24ghteBuM8RzJUfzICB4z5pGCG9z+J3
3asbToa6kkjKssFdeQ4+wkAx2eDpEEts+Oa32CpzcQRbKuWfPctK+4IUFvmkahxe
TUsXCqxfHIZ3klB9nHSTN40uJ0LtxDtewzdDR0mQU5xG1qJ01LmzrOr2xJ9Iisdh
xURW42D94h5M0h0wH9Sq7IhvtX0Q8eNrFcJ/UCQUqzk92sVvDHNN1s6PeJPO8KQK
0RgH1ExWq77//sb2lUZh831MJrC3T3OsrwDN0xqdd+uoVHaQVmhOrsBxnYchW9I2
j+GzCA8h0eiSQygjCD7simWBvrZADur73DngQ2h6GApAbgC5l4P8C9XTV6ROpH3U
Q+aFWBqLHjLvRuWqxpkkd+wsb6xBdFwspzWDueZvtvvUx5a6S4ichTPmR0i5DJZ+
HIjb6noMTdxL2nKl5ZqDcxHukUaDKAnVS6i+f5o+aFZtvphbodzww9nxXo3BzaKG
EidjNFsSziodT8SvuWmNKTMJCP7+A0ad5+ZSV5+ApPpdk0vDdsMaAY4ItGdZg1WH
lHrWuh/pY/ScZqEw5/jZjjmNd4+OtYSfFcUmy+hWpoWBfGKa2jD9S1PGilUxgv5K
SDfYjAaRwZX+a7v1XSZc5UdnAWBiLyxHgDMzD/AfJlCNfo+vvrq2DpI+0Tu59+Zo
6CmeotIwKT6V1lV+lFO4nwb46qRrg/ha5M4fWfCd57RagG+2KMi5wWAVd3HI7xjw
Vz1Kr37WPhrUjTzOU3l2XLpb9VNeaCaBhn7CsJtx0yLdmXhwtogKWy8YMTjjIB+X
uUs0k561hf0M8CqwSzH8ea6trme1Iih6p19nwpFV9c3mKBKMTH8mKQcshoigUcfB
X0RPyx2HXXjYaaO4CZ5/yLPlPV+w7EoldOOzaQAdr0GjiR3aHJ2o0PWTn5BEj88J
mq/9RvZ/2oZaXkVcn5ScuQ==

`pragma protect end_protected
