// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
faWRAA5dCFQ+AWYhieNmu962FtiFK0z4CM3lGWRphqGjdgf6cUCwV9wK4RCy6yP6
2uDXLajyEfUk5ud7wX1x3oHjyfSMOAMaw3MGTF2kDnoZ24V+tMarVWzI8keT+vwL
PVfdD6t3jsOLn3rH9IbU54gU0YEHP/SjIYDkgZo9Yqs=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 10656 )
`pragma protect data_block
nBm0rnSimwdfg/Bx5NNB6yMaV3UYcp/yAjxMPO8dLBQBe6XMGQEu2TwWS7hybu5b
w0WNLlD1upO5SA4ZDkVlAHY9YjKX5fdq2lBFtRgdw9Jg85EP63MLao/2QfcDoXlP
e3AX3u/m6ZVSY2HRRXXxfNQ+/BZ8YFI/4SlJnIBQnjlsKFHIIAUMih6Q/zxuTHV9
mAshxyhgzkkf1b4bQJV2FtS25BI/CdXUjYdtcb6qIwN4/pPF3PSQI6zXRgFUZd9/
05LNVRg/PyHcLsfGjjGAIihTzfqVd4vBE2bX9D7TrDf33QyN0YehD9IPN4zgFwIP
ADFJN2J/30zS9SaRytv3d3c2ORIWXi3MKYsc++n0AMX4AGyjG5BcO3l6QeX4hhs0
S2vSiYlulZfMbh6NhCMPOCgK2q7slGa6pxI7Ll5LS/EG3YhhAqT8sw7WramUmWgG
VvxQkcCgMWOkIA5dBiph5qQYxTKElCg8aHH9KMJsF5RaDpNQasKqT8krnq9Z6jQS
3Zr67hJyIeNZ5mVe9sYspDBvt+XU5QKXe72aLE7pgoPa5QTGl91Zq1Y46EF6Df5n
kevhQEe/a2d1OgbRNIQy0QY/EHukR1SpZfdL+ez2b3icIXio1Sf+3kWuwcWTgd4Q
laTmdX9DTsWnaqsvWl+nejTHLlX2WQIEiU641b9CSrIDT7qN+u/uLK4WGY4+5sR7
eYFiKmFznrIRu9X1vfPN3UBTC8z+cgD/jWXbUnL6r91B/msjlrdzEWdmjasfI+FA
dOkdyTkSbtpREsRNjy9thzlE2TO6w3LC1o4vot9G8ql4KkqwsagDeo4wCTlpCwQb
6W4a0lrju/W/fUwVDgDFQXdYWoSfIMOekK5Q+59fJvgDGRalNbCdd5KphJEsv3kq
W6R7WwQ4D5q8FOnYHUMQTsRyVia2D87JSROkCBe+UMSRjVlQqWn9SWDI6USp18OQ
laezIVbETB1EJjmMrqy/faWEUKb+kllCpaA2MLLk6ncj5Sq2hyaow6BO3I/Q78mA
dijwoRQl+f0gNY9aAxkC520UMUct/XnlIrPe755HnKnKk1sYiSWNZRfmTsqoTifq
hUjQf7xpk9gHbvq/V0nPzWzaKZ/x0EFlgqItHNLi2QMoTzhFZp9Aum7I3LI4+p4g
oPG849ysWQrHlQynSjrgxxOqvVyGzTFk41By8Px+fFO0ZurwDi4uuvoVxQRK3wBV
rnvxPUGpfvDkEMFcqSd6PHJlpVesH+B0j0wLYOknx3rN+9deU0iJ8evzxQ7Bwp1y
l+iGvXtRU/npEjrksl4bDDAGWn0Z2Ny+Usv2g0gwlu6qOqT0jfP3NMgt2xk26VOd
mE7oZQJPC92SE4jMqexlvmryaCTS397cb2ulGjCQ38iPFIBWxmflv2bpyvEvvyhn
wHnxC/m8X118BSCa1aSikUTAQxE3cTa/sSzXbmG9sn8NdOxuKznTf7IDqTvyKWbR
s22RmV6QHhwPhWczPtukM/cKLOqHr6zXmGI6hPg+mYsDwRErET5eaUXVLj3op6/6
7Aqv/mHmeFnVHA0eHWDG8x+mhrChKf2IIL7GjXZS1mPXellQOP+9v/HA2m3DgWCg
yRtjQaQu78iVYbca2rlOVaJIC6OcAfRK+EG4YMKvP3mfQ6+mKWGBN2vQuDMq5eze
9nFtTCIjHYPWD0bYnxLsU/eXDi60v87Fdnndc5mg6Aa4xToEEjYoOyETlK8goKwF
DWlD8DQNQeE3EjoaJ2xEyWI7DcfRsbxMZqzeryFOk8u9o0lyZm2asIgcyBNmhtAs
rQffWW/uBZCjeWVveSM7FutmBUlwUddsMCB/OciI7fwlx6XVtjGkm6hZoA9m+Bsr
5TxfKFvs+iqpr/MmJHBOky4ku4M6sZVDdN6kbpEHF1QxDdV52i20/4tjX2xcDc5R
U2VjlJAaQpM3ZpTVTW+xaS5KMn6hxjvAWrnrxfaizgEm1t4oB8fDnSTaCuGAEMcb
HcJJhLjeLAapkX2gt/hkZ+Cd/bHLu8AC3hGnYZL42n19o+8jp6NPUfK8s3SYcc+E
btJm/sX+LUFC09ZvJavp8wP3pwGBybDh6jpF3BEh6A+7lsIBmSelJ7nV/sUKVJZH
R9S3zU73N4F1czQXC/qkzBr1lfHoUT7VbasUydBR/jRYeMfKa52Zs4WfR/stvwss
VQFKuQAe3PUkrXYw3v7KPtATgsVnwbwdoJcunWl2LN3+V5+V08Sr1Iy5ma3aDIIF
ARg6QwMtfLDSPQ0e28HQBjaLKKXels0DSjcEVhzYOQPtgzty8I/yFQEfiXBk4wIA
bsWfIaUDYrBJW9Z/ZyB5wrzXJsJWw8QXKhXE8eFlOvJjC8/mXpx2Lw+6NIR1dr1t
pMaaoRMTgvjJHNV6MQwIdkY33Mxp9nmcJ45fyQ/fPoerCbkZWoqg5QtN4DKwBdXh
wPqXY30rkpGqYwpKvqTZLWdAzmvWPeVsEF9SXh41KJdqJbkjzK4Fs6CV14/BJJ+6
rbJ8aLD4s+MfFbLep8fU8oR3PX0LUcaPyCJS/swsAZReXzYXEDWOTjj79VoiJTa0
uBY3p4dKFOkwtCJc1zvGiaiA1i1PD9HAnRKaViTysTvBekcQFB2cikG1yVEjivVy
Ic57q9X5r6bRZidM8l/riAyx45yaLJuCFP6s6cfTF7fjTzcyMyRjekgt8AUqqtmi
ytf+ZjON/ezA0YGCJ7nuqh0hYz1hgGjwnDMyaY613khdjE2qesqrGDZ6s1wEdzOw
Ojmd7odSEENAoNAAx7EeiO2J8VTV8WuFDanV6dbZs/qBdpZinl82kgZaSYrAlWP6
SrQh6jqto/B/n0DK2GHDMRib2P4F4Cmv+R6qsiUcXx7yN4PHIE3eW+EFWWfDu9FK
cb/k4DDUe4GjlXtjXcolGQXT81HMGHZBmo4C9/sSXSUpzcDVWg/LTfP9HJ/5mZXp
cDTUh6sFhq7kT7d28cTaexiCyXYVcdmgovjUHuesHoI5OYjtLySjip8zNp14jKdq
qwldyQ11KVTdn6Cxt2rZQJkkaRbkEggHkc22F4JK4amQ+bw9RCIg22eURbmMEqgO
EhJ/SD0ITfxYi8ZMZUpb9q41z3j47hzgrTMJiTRkgl4mXKO9MEGXekD+MusFIDbq
nwihWEW0FNwd6GeLvAPnzpGTps7t1P7D5YSHClbBQ2E8f6MqQ/seSx6I6ylU2c7U
wsKEzrZL7vLaWqyvSSWWqogn40y+Z2d4saXuNt4uNCaIg3uoMpi/MkE+SbcfutF5
r3V/tNLzQ+pchZIkDcOuaTHiNypjD+OWNtMKhxgWQbT+f1RVyyD5DrW13t1fjckm
zr+0Nq2thzAdyFPIHTy8cJqyAa1N3FXPO2/yaBsDP0zeChBVajJz8MACjMY2knxT
i+d9f799+qh0df5EFbH2kEpVh/4tDiT0zoNOpo9m6jnnya9rENaJylAPWjATKTrY
5y73xaDjCYXaNrI3HyrCoZgYU7VOLN9uX6QF2YMUxvf+G30nzQn5GYiEwujHJDvz
JzMvmMlBfgy26kSM90S5FHT6nOVFS9tnFUYFyDdL9yMgDStNSJjkGygwG2xiy+4r
cIE9YqMMpM1VpFAHd304MnLEsknu0J9lagB7tEQ4RtO7LIYlskNUQG80I7iKck/U
GPP1DXkN3gZ/n31pjrEnIboi7lsImpGSBaq1sO2OwrgvT9fl60/n+HwlvdW8hb+8
RngiTBDOCyt+v08PpUSNylY4Nb3uFqQELlSuRf/qd8ILZNKgFwq+vIJJrM+2MaMf
4OYwjtmNdXXzoJ7GC0L1pK9eWv1kq9AwczNCskLi9JcDDQv0/yAw0zICiESuDqL0
tC8MEP8laTfi6LXqm9U1NO+Bu/StJ6KpQRSkGFU2NEw5DnLcr4e3qGsANrVcIFu8
zzYs2DHpxngtMW8QGKaPU68MKpsKROrrNJCHwfftw2++FYy1QHsX3SqyDW9KcdgG
ZsZbFKkT24UolPzc7fTKp/SrM000vvUiCZ/IYlnjJeYe8EhsN5DHGLAMujc7OfSE
s0dgvvYBXTXLJXw0rwNErzJQPds1YxvCygjC5wJTYTR2ONNL9LhjJyMV3ud6Q1ND
vJQGYrxmnkS457YeEf9bJPCOpC0ZXunhCT1izi2R79giLOkeW7gByAPmhdkSBxKe
WsASsDWgyCjkR9dJ56MZMp/VsBBuS6QklpPYGWe0qxJI1hV1nE2JaQ8BuFRHVPFo
wS3BCKwh9jbXb+/vro/1nmg9AigaNKAHfoThIPY/MlmS3h1pmxv1WHIWP+R0ra9V
OtG7tZfr0WrYCPQ9CxZ4K9U6FTpg5xnGZVXNXBOa0KSir8MQ4BYR70H8+8M8S8Fj
s813SmlwrnpolivcSUltL7XcvACZGwRXfC7oWmfTwYnbO9lfx2N3czV7r8kDJv0F
MIDM95WmPdVi2tNE2ueDzjkbmocN1X/qzmqMb1ONFCKUI7jh3CrLjRPIwdwNmNVu
e26mZs8PIPuHBTUsS3HBixo9oNlfQqqW2wOHa1n3BW9gselzPMHbDXGgHZi6DF8A
aE7qKKu6D+5NXRtS9BGiobvABi6ewPwMNuPblJeBN/7Vozw6n/N6Qeh5EGr00SjF
Elh43aI1rPg0NgAevnuInr6EvaVdsQ1GGk29hrcCEVTaXz0uW7T0c023uQfHsJu5
qDcp9B6TOfLzKkv2Mj9FlwMGCCl0W15+Ueap9/tX4NQN1SIZDJoiAIhm87cqMYqK
EnhJ5TggIttBjHFOMfYEUofViog39FCsBvonUQNwQda+CC2Z7w70IdS7twboCdtT
Y4PGFlNTN0bGfOwOgobs8A8aHRJnlPUh6Pv5uUVr2G2NDznEwnzqD/REXJU4vh9e
H/12vLmCN9EV+ikJ4YvJTJ69U2uV6tPTv1G1rQxCtNsX9X1OxCLhP3FUpx/kmP0y
0zxAPpcYwRKTmbZmWdZyc9VTDRukmLxv9zZQ0NZ7rpLALM1Dr6C0dgqMRoejJVCd
TzCNjLh60F/+uy8oSx5Hu39GS7ImkB6dAKxJAUGvPlNBgdgtOkKlevC2HVUuUiGE
Qh/0z3JqSmwECcsV9Wi/taDnNeUvTebr5jpdEUkGk4jgyTu6UtWBH+rxDR17KWYD
b66EKaFWvxsuw4gJ8ORNIxBKP9WRZO3eM6XOfvWmM51BOMaOarDy1o2MXw7BuHoA
daWZhCuR8tn6I5DsN5oGekE8ORqAOKfKQdNdvAeI5vq4W660sCGZnQZx60nKBvzC
GsXQe74NmhVldNMPP82asfRPF4b3hpLWZ3mnxf33sHiKzqjg60pkOCxPp0UpufEr
VPhO+GO7qxOr/1Isyzd9ASSBdeJ8OKBbPOXL5UkY6rmnUNIiHHmwwUNFB61fiXG8
ZLckOma+M+AZiswz6LObJT0uxVNzpzJ9hlvx8vlq5GCcr3xhikg+Dmwf6RR4XHFW
ULkzxV2R1m3Jyt57x4ixrBS3URTjMOvTRicrIdbpqpIxtzp++GuoW+RELQbu4r8b
BNzyRARLbrwhrfHwUr0ea5pzIWLC8hnlmKz78rDieZJqShuHI5PA5h/Sa5MGhaCd
UyqnR6AHtx4++nzq2exPtRSkHfJhky59vMDT7DsiHlXK4anH7fd77FGSzZ7bjVaD
eVFaQyDEmqIgfKUjpT9WYkLCPorOaHB/jnrnb0J0qMm0EISuL0cIQItnxDLERx6Z
+rGlWFfQ2Mk2icaGL5Fj2EelvuqfhbvssW5rIlZqMwgAjwM1c0iLKOehotP2+55e
3L1cm2tNXp1khQkdqodGysFXzXk1yGTS8ZHNhaNGFphxRTXOh29DAIeVWo2ngAQ/
6ynOYFZPq4hwmwY+0gC/eMQ4dCuxBYXpeBOksy+RAkc3jLDiX5cYqMWyRHcr1Ov9
ozPhoS2mhqQAK5rRB+2DIzmqgncSNkEXGbd3aGlJaWOYKCNhufCVKOvSHHmPMHZT
uI/G9gE715UPdgKoQvwCHOVzdYsFOlUFaNli4GgviHsVbc5sUIKJKvlBMHYJlsym
OCyKMPuP2QHQjqEsIHRlzTsMyqFmhI1x7DaumUF56zIPreVWvKH6eK0vlPeC9OZ3
v5WlDDgcoitzoGvstEO5CNBY5jdOi+bN/D2aVhiE1qrVoxvLpYG8qy62t8v08teS
qDWVP9CwnPXWYL38AAgLhuvD7IKdfLLKhMl2qcUeSuEGTUsQY89P62u6KaoquR/I
Z6syHWmlS9X4drWVWaP2jkHAW2a2B8UscasCwXUR3SBw4SLH+3Lwgb/gUa9X9ASG
7zv4r35dYk4CNFGSuXx+HJA7m1xaKA3X6YIdsLxNfd+8Gsq6h4iBcVh+Bn70+y/a
WUCSSaAMUdmg5rZAXvY/hpfMZGo5JrVtMxNVHOSsqe3wMX+vEEQD8ia+a20CyiAS
KiLu1yd9j7vtRpsSZh0x00OgfdlLqzFph7NZAGpeyluurlWI9uwMfmgY8eP8iS0G
u4DKqelaiAHRqhgmH1RfNKPm8hZC9qMFZgACF5oawF+ukaiEHfz5AZu1rGx53gMz
L0CUt8EYX2TK/EezgYToYdjqjTmDBlgwlmvelyui6UtFhPd11XwFkzEC+sBwpSWN
TXT3jgH8fOtsb5o7kSByfmMtQCUa+UxjeFcKPrtEtaDSuOUdxqeddWy3BqKHSZkM
LeVL0by1sbYw2sfJLzxwTURpCTKw1NKVarMTQapHXqrN0ep4H0+SHZERpf5XdgQ+
oU3fN9H+pbi0+f2RM/D+fo2gUkvg2lBHjL8tyBhCRU8riSvp1lqWEczU3NFbWOsk
WrdzWclYI+VejT8qXbwL/6dM4ZEE4gbZkOByvIu0rEttR37yQQu3IWChAfsLmMLt
dihTga2NYIBfBJyReFMifVKGUQiQPab7NVEmbPDzKG57AATgvR2+jWFNmSpc8ug5
iX/lScCSh2xfa3alixY3PlK+Lvw3ccL/SyIvhEAp8vhRXUcDOMmO0qHOOSnvirG3
js7W1CjhJlCGqm5rh8DVxHPDKGUHAFhCTCrDF5Iu5KPtImoMSU73Qn9C1fo7Dfta
K7yvw3B1UqJGA8ZRm/0iP02QCFEA2vFQfbkrbVkfhI/Zi6d60UEnzVHhZeOvZGBU
5MrHoDQulvFG+w+3KtmxJqkPUQDVEBDxcDm7EIsE0zcVW6wI7l/C1JIdpnxVd8BW
PTlOWxFHx1TbVBDiQAAn5YMzlWRFFnPcMnNsPCAs3AJVpBeWyS4WcoLeVt3CA2YS
XzaTHn32jwBPVJe/ZoEwngrUKp+xiiW1M01LQ3Yv6cgFT4K7OCQPjA+Ik0K4EUVv
K3R6gBzgOLKXFCAsCFmKQ4jgcF3cILDo4pLbIrl4atbNXVTeQWbNqjAlG58slCwm
VZRrvONtlTPLLbPezGNDGlV4PiYosZjHAHAq5apNXyZ7SSAahauvymBa7AQjOsu+
kGi8sO07bBAHt5LDdF8/S7O91wRF94AjYAac3qiUx4d2xBaWYINOIfoX0YujO/iU
Q9TsiCu9XGS26L0qjmsrq67gJQD1ZM9KBm13wkJ0VEvCGxcFNme8Rf8XMuKdkpA5
yj3i5AS29Bm2LfEFzi4ZRs3pdxJuwu8JOQ+4VZ1tLKE/vz7yab3j8oXgEOZfN5gE
kn6xmnQC1PefaUll40VaLL/muUA0f9VIyZXUObAWYIwt7O5UciqMCDIIQ+4aEExn
FX07yU7wRnEk9seOo5U9VCkwYMSRDEQ44OBPFL4GkarWFv6weD9kEEJXbRdDux2L
h+BGz3/1uNV+1PkeqyTfd42y0UTFGPoPpxELuDrarnrkXjAq8wQw0hMUYGJv7Png
KFpPBQiisX2VKiiY3BW0KCJzRbu99RmtweuKLHLNMXm2yEntHj7UL79ru1ecvEah
kHO7DvmiCCFWajldu3IvtLOjZEQpRERv7T2HcWm2nrghl/FmN/xatSK9pGEwfQDT
u1ubHimYSPCvEI39SXjwUPZB5iMgCXidztQO12qVDgpr6MyBb1mLW9AIEBU2gjmj
gDAfr5Sy9fHhCZsYRch9hUVqzxZOo8TTgELDTWOjy2z3MBIlkV05JQ1q3l6PQFqe
QVlKeei9ZefaTCQ3twd8ELDHmVagH+uRArOLn19lHwxz9So9A2F7BoqhcBc+X+IA
CTQdq21cVXbF7NvxES3jupLbk/GEaZC5o4GcxVi0xyh50frNH1EF9JoDG2Vi+21V
ur8rv7PGj/HlkkheB92iMfm6/ZtUpzXOElQnqej0+LBsd1+X13N3eWNecQc050ns
YNb+bbiHJu0DC/A6ZhSbDUIBypXqCr3Bg/RfxCM8v2e4lpvG5kNR2wc6w0NiV1ed
ygpfhj8YwVI/oFYaD+uTTZjSpT6L6lIbItv8AulbU+YmlhnLSjiStpGh+1uRfTz3
xIL6wMLcYU2iDiXPu1nSWrPIWlyF0O75qNgX6bmqzTOMlZ578p4MCyEnQRRuWqD/
GewEyefN/3+bGjnq1Q3PMw/9h+Pz3xN94f7iocDrYW5qvW+OI1hAjM5R09koEYgg
+FrlB/IazruwLJ8yw28GHdSftv4VqaK7w337C3xQz89CInlUgWbWJyxff7Vshf/V
fZ58bhD/tPtYzQ2BU74bVC/8jHZnTZ5Gpv5wtRKhnLI8hptIsHkFjG+gbeAU8lVt
eKW2z4DdE36M/vH4gDVAOS9TA0gxyzfYnLzv3u3YhMDbdq/HvCEYc447bhylcbrk
vxLeeNwVcmSXodzZIFB3C0phQzbQtfNgwiHT1TBV5X19sAy8FkbMZFmvvkO/nXit
BGuDvB+MtkCNOhH3yiLSrGsbAgnLtu1iEnb5jXDMSv9s0Hqdjx8H9sQ+fXEP+JmY
CmA/AHcFIuvHjQ+pryFj41oFqFjLIf68sL1zgkW+OXkgC5bnxDE06cdDGXJbME/d
YQ/2iebJFzJAVqpRB7sk2s/iPHBh3QQTQd7tZnvfIFZWC5PTldvLvKqfICBwYmuu
xviDNdZz0+IZs/fPn3F581UQwqd6k1I2yvzkHbRjinI/JIAH5XfaxOViWOQswxfd
uX54EPQsSdcJAicsleYD8/AdkLs6imRuGqZYpHadfa8NfWKOaMuA5F1PeHZLBlAb
zDDge1TsO1fTwpNP17387NHNXhAZsedbtvNvabd4s/0iAABIpTf0kKlQALDqHe7Z
Kiy0aiSuezmvBubeKyaqNW+wWbElL2wMNP4XG1QiNfsVDJHA2cHYHbnLwvhYHEDm
vy5JyFjmEGz9sbP8y8G+vI7rseAx2LI4orJdfreDWAMy90aVUCWt3t9jdzsA34Ly
nWM6CzE1YING6gZlDjoEodiLks1KYgBZyE6xeFCU7KSiU5dSGie5TlBhDinK+snp
Qfqij1mtkB3GiBGoA3YUtuUzZPHjZFdtBxPnNJMsvr0zWiV4CUmYqtSxTW4eNQGh
oeP8hR9bIgw/K3Lj0zk6LxL69eTWhT5HHO5QulFyEBjEfICtUnJWjNsRXrcfZOlS
cyNWiAXu99zxrXJ8PRnMeOiqU1TIPWvTMcXYaBePSpSH5luQVCy4YM8Ef7pyIjxl
AvGJk47GB67C1+1ZzHP5Z5Dn6IuW7fuAkxFHJ8h0pajKC2s+e+4J7QbB7jufczf7
ULGszhuQ1cZ/xGN5LuWjvi8AlhAwMUvr0BlTefhAMuchGru8srr0i2vu0HHRoYTF
sC2L0++Pni5jUzkurKkzNdCw3TKucU+MS2Xl/RAtvVRn4bE9YKvGf2Wgfi0+nkD/
OWKH+vMevbQnjbqlxICTJllJsKnwnJ5OGHuhn5R9bmtPadDbefGKO5GnfFCgXG0f
ghKAAQNSm3qO0bhc9pzQ82d40auRJvXR+XtvaSizcF6X8mIUFPTnlDwN6DBPu4+o
9w2UoKeRX6gT+OUIDAQUBFPmRpwwHvyfz8l5Rxlzl5nY/CDEZ9Dvi1HIK7xzwTqA
g4A1UgzNacENu8zc+/0N25wm8zkLRTh8I2INURudXrBqojULo/CRyGAkC1BAKfpo
Pl0GqMT7cGE/nWvYd1DZiBZO95YgYt5zTK4i8mhzSAePVaZbj6zQDcqRnjzuRyfq
1K6YBLqN4qYCJB4RaE9i7AsuN+Ruk9IdoyEA36oHPId1DixdI9sThJxE34xG/lWH
4HfWdRvOub1QBjbi9nAvoOLQqZqrnKuDmmT4SATbRdcfU4Bk3Y3EpXnDWOTKmxAf
H62qV6wmRlSHuDLGTERrtY3VMQkccMiHp7QQdLcfFN7P/rHTNsX4w6Qnb1zVAVY9
MF41g/RkriwrM8vIL/XJJZu43CtGo03lKri3QSaUC3JDtUEDvkxMz4ylb04fuqaF
YN5DJyH/KxKyacdC2u3IAnOHATPyh8m+5fcZxRlJ9TAPi7baFKKlZPnWQiqzYI9B
crY4tJ5bYXj81tENNs3HDvfSakKaCJ2jNxa69PFykBh0PsmHgDmFT7+aOmpp/aFy
m6LDqqYQn32EKz5dAtMQ4zkBJZuAlvrXz10UT32wDCumvVgzBdkGMpc1ulPhWV7H
hgRlKTMYGeAFhC0ZonQdoqc1vcifj4Rztn0UFkNcJ5IveNXzxXXetslaWONOwuDI
7KjF00yeib2hjzWFtUSxtd+BY9cZSnRC/eJHwrLt3W8FyK4+ScyVslZGMhwMvFpU
6smR5La8seBQRV5dE9kAjUBmTjsvlqAvcnymUXlxRhKfazZ+ampNi6FSd/KAtvS+
o2tk4grN5KlR834mECGZtieLwlmYFCC1abgVvp9S5EoNRd0mS66wJBKt3IIi99Ug
C8WCZzqe8NFaFqKxpr3KxPMP2KyzE+zy/Wrlph310uZ+CqFlZgMf5zbQy2BuXHHf
tGJGcd1BKW4fCRmBocSbbzxPM40mY+mon254U8A1TcrP//HphrqIyLWmySiHa6cW
lXlT+hKoavnTekPTmP8VJSd078IjW1dgItSfUXQfqIAstTFjmKTYI/zfM0g9nZy4
F9RRurbd/iq5Pma2z8g/fDXMNbpaty048+BqkLf7tzog2m0YzorrTzLqVMHl/dnc
aF0UKVB3HKWOhBgQS/8qJwQiwiNTPuL5Z2za3zzTJcBjQ8x+HwR391naoaSMscLN
e+OeBBCxIAOXDnv0/wQpRetUzAJ3jN2EocYa38oogUBBYzej93LAeeSynUYx4n/K
SNEGPi6XVz8VE6VqRkuWUVZWzwUQVAhAaSONhmeQjLQXOxSBIqgrl1OHtFoIolfI
fHEsUYRiHtfVDiXzp4Z+9CfQAR50tErty2CSfnyzGpRAR2Mi7Mb94cQEV18nDdmc
cagbLwFk3BKhkKXZP/GXd7OQK1ekMP6liE7lJnU+OK1YX3qUE9aTMEMd+j31jZF7
arMQU91foDaTpje/1Ynqf6T8pG1cw6ZRBhlhmtC3V4SCPMozRtjToJEaqFUs3X2L
gHRvXavEZ1t7zqvxsLZD1N9BhmLXM29oqI9rB8i7yi7Jolt0HNM7V/Z7JtwvlNR4
7KBuz0gx1z1CPnVA56pkCgD/0rUa0oAWkQjqf5J7DBpxJ0MUDASnjAhhWi6KNpPE
4Y5uidyngdC88065REoMKdCUpBqWtjyOWiQK2rIoMttHy83lIWXa0Av9ZcnR96rd
3YjaiYOZTeEurm6Yg2mmnuyTl73KF6JG/rXLxS84XBMIXzmzJs1EgM98m6kimj3Q
0PcmBSBGnhvHifAkPLFxlFxG1CwfZSv2fpUoQXhWZMM0ccO3VUCgHeVxREDa24Zc
p7xoPS6yhxUdqS/+0navX14j+jqrx7DXVjAfL7cn2UFL6JorCPLVOP6uU0FhmHXJ
pyKE8cOR0AOB4Obe2g1st0XyAzeqdvPTZHRN1DPVXalsa5QzRibns6D0yU8EwKoZ
kENYp7toOkR7rSu7uJqj2WH3XRqfu4gTIiZ4HkiZILP+3BvJISGJ5YYwD1Dr+L1J
Lg2B9cYKMWD8Pl+Lyt4axPJpDQF3fAb8OwSZALhDw9dlO7Zug6gPGHM8K4d9x0SV
8WC9vmN/yfTsHfBmeLmqZOB2+jS99RK0jRrTGTTFsR7+i2Y53e65wGd8DXmKtNEx
Id8i2iod8vz9xWNLTo8XeseW8ri7hnk8OnViCEj9jVoNcusn3Q9X4mq5zq/OOovR
dw/gvyODFCHd16+VoRkigVMIwVNC5GWBF4e9z62WoGLPT6vFMQM74ewOxXKzulT6
I0buA9xnigeHhOr+/NSOy9zZ/f4woOn96/U1EWoPNNOmUeTOTb6l2dWS5cLmLQ4B
2yICx/iDsjMj08O3F/SrnfJmFNIM5GVApl6b5vX1eNod6yHiLReuFo98OOeXw5cI
b9LouocZJxIUqDsXMMICSLH2q5IllndN2FKaa63jufzd9HHrX6xe6psuM02pqSgQ
BgP09tUPsYwsDT2YKtJjwLEiPPFSZwptmZSzPFbBoFUIfHuVkWEOLWbnX/FurytI
ru6NRBtIVOPzIRIiGaG+m/E9SUSAaz3tV47KwiOuq5dfJSZPq9FJWRcQgTbfbEBq
PsdMGgRAFYQ6b0oSExIDqnGCtfnH0mgvav3NvmxmeAptET1VE4BH0+fALhvE3LZG
5T2vfAj6bRlGYbT5P+ol4ZIn2t8oOWWZxsGnOYEYoz7wdJqdud2fckaiVuvxtVKn
T2WvmaZpLn1ADU9QRfhFxPlWcNzywQKkvKiJKXjThRAVzuamgQcFeySskl6Fc25t
T6uMBMWbpKm3ccoKR/TRVB6AS3J7qNosvDd3hdeiOQbfOQBSTGVBzpGUxU5HEM8I
mm8IdsKCf3xYF4pgxh3nlPG6VU4W6ij4IH/lrIX71Mdyv8/adG4qYed8Ik1IlOJY
Ai/laoEDTHqPaGG93KbCawp0VrwTfXdU/+kMhPs5X/TlG+yQtiweZHjqLd71DErK
tYuTMpO7ehsWgWTEdfpbnysczCh9jukOsVkr3SDkJcIJdiQchj4xA9gMI6DX97uC
B99Cv4Z9Ki9KkZ2OqaGeLUo1oorTe9yB7J/D+la8ghu5bxNK7eb2RuIse9iAe8Zg
ATB2i4uGRE5dfqxeiyo+fKh/82rzAyF7Bfqsbab3mMymSXH9GYpJsb+JE414I0cF
VN9KKHUvYA2tCHeIiKz3K733dDm6MNohGxiSx3m/5M/N86XK3QdSsPSRS/45/d3b
XeJ/AeAkJNPWD/qqdeMcqanGDfDTaLp1QSu3BWQ6+ONc2lqvq6AkvrMiEWzU7S8Z
XEx4FDTGuqlc3nZFCt47in2v25//HiKY8RgFjrR9hPLsVFmjTWjm5BWZbIhHkwAx
rmfP8nXoxzqD9/ByBeErhc7iLTiafWiD0dkfJfVZ2mC5Ck1ArXqjDFV1DWeINOhJ
S6kZSK4a4ItCo79VKRxyCSNzaegmvNN0G2zawqY/VBOIKMJ7qd9SPPIMIfgEv3mx
xRQirU+ujdl8IWGDiKDGRtcRmqIKWe/R3l//1S0DY/+42/ICeZVY1+CIErgKh3ao
tM9t5RDc4Hzi2RGt3U7H3eZwiiS+dNJaVGWB0fngeev6NjCjFySiwuWTNc+qkR5H
WkeYgngtGtu9oM7tRchlNln0FKoF3zloJDefH10gyWPMYyVUbRcxp6DwJFAsQPaG
QpFTd9DZOQdnO+CsBXvTQDSZYbi/IyBWdPB1Jqr8g1RsYOQCDaeVlXuVfTNn+gBi
mToyv2hnpe23tg0cqb3lb0FKJvExUcSdT/V2hA6fW9JrsIwMq9ly8OGPuHnWGe2y
WwvxFI+m7eCMc6i1CSzdsHFlM9Roar8lUbTTrDbK608Mg4MPOS5/NswM1MrIhH51
jqvMyt0cgPTZFykh6Fy4mG2CLXR3JMHekMaj25K9A8cDDoWgixzjf/oB8VtCnDCx
pRLohyA0kaTtqd+7FIilBsuQ4LavJxcqUU5V8Msr70hSBcEKOsI8Zsfgncg2GCpT
0Y63PzbGOlvhbAcVR1PoKsJlYM8SoOpaz5yQ5Oz3mUoeO1AdG8QZsFMEyx6Cbdyy
QwwBTCLVNQV7fY94oqkht5D4mpV+2W5R0BepHOPqPsTFOOE0jeUr7YO+7k1htjvT
3uTo7y1YNo1RsC2ZPQaXtzFFW03A8RiwUnS4SoIAajeQjrR0EUUTC2+JXch8voWr
4Y8/l70S2XnNRwC9WTsh2WofVePeuLV6Wri/xGTnpnoxux36k3kFn2eEdZS1heeN
oZlaB/WaxgmXu11ukqEbs2JM0Oj+COHAMslem/CyOebWSf4AVDv9iqvq5fq8nUYT

`pragma protect end_protected
