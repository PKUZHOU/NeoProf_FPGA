// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
kLnr/gx+hO+Xw7U5fJI57wTc4Nhj86hmj382jrRKFU4qiDjERZWI57g4cbGNTNM7
b1w736O9rGljYGN9yE2qjhB6nTLABbe2PZbEhyFWlycYSR9BEnaNmSU+itWKmxVN
DBxn96HjfqueCD3zckMQ/iF8njWhRF51QPXDGY7pYpY=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 71936 )
`pragma protect data_block
TbprvfH2IJV1dyRn4ppwauX9wSTLxaFo0NKdnLOZFsk8hDxpD8ldsGW45WY8sX41
MB2irf8NPNUSpK1UO28DzTqN1UTlLFSLwVj4smXWOktJZ5sCcjbGxRPOWM1BEHYX
3Dhx+151XNHVDUAct7deR3bXBIxBsWdh9oMVPHThcT0ERlttrt+yU/e+FnuXJAFm
Cz2x0UBCtl1xrbsAF1v9Wfr+qmUaqtc16Fw7um8W0T+1XgmKAq0/vGkY4skq/ULo
/apful4YZMTbZH1QzmxynaWDc57CWgHHft1Zuo9HYGE/40QCTEu1fu4iAyGDYsFK
3k7nD/1UpeB8j4/JgXbmQkzpMMkxyVeJzJzVkGIzUUtTUTpe73MI+e/s5y+DGZKN
Pbi59qcQGR/SEL8eOhxIX6db7cY+7Uuk8nee3+zuDXtQYdzBAzAXftJ0nAAtq0cd
bZWId4uqN9gcy3mQXWXsnRgFZtQQjelMImxbspDnBh9i8UpHL+Ld7bvar6iC6NJg
Gooi8s01iTt0pPUMN0/ZJghz0p6VA0czamU51me8fSZWA93+072ba3YBd/eqI9ir
mrgCRFcaoN3lYErZglH+4n9x7yA1xvAVdH5rzxOjlXFIJee7s8GKZQiF0dWpj+c3
x38QNaE3SNLHyvgDeHZiHuEjIFuuxJB9T0MAqmyVmBLPFGurli75bw8LQdhTIdvP
aIGpsAqPdiMoeA4fxpDipmP+CsJeYBXEeYEI2Nw4AZfJUVDTVcPPK+DyQVUX8p0Y
EQ5U8foW5COHStfKnZ5rc6B/2XkGqkF9P8QOyCqymvCigH86Es2DrnYbp/gFsEP6
sfyKW4mnIUtA4yT/96ywJAp0kSS9plsLg/FeNZzX+7ge31MjgHrga4Vg8yuZWXhP
fRvqdLzhtiIcvBS51YPRjciaGOJh76nx8iC75+Ki2dcghU70cMBCs7yZ6ikP3Gdu
s34kpS7a0C5u4p3HIbceKyCJB8TkwZjBLKFpAFb2mtwE26Z186j4o6ICsyogsMHd
x0/ydB4SA4dqA/VAdHZMFH+35X4eb1OvYoHjdN4jjJe4oo4YaB/eyjLplkG9kOBg
YbuCAaMklXH1baxDH1eTgIqsGohzw6kcguApbHgHvjIrB2ntqllxhh8gV5AJZOkv
u91JoFn6QxgjoLXVB1b27Ht4HgpY6DQYTRDskId25zmoTkRdoIQ97JANHO3O2KqJ
AliugWTh+jQR3xzQYB67CW8hcgOuARi+knkMdnl1Euv3ceWgDJLI5twNblMLv8tg
xFH3TmEllXB+6OQ+9e/OHFbAthtZzGvqzEqT8sRmgwptqjcyIkC1KFXwACOCAv0l
CsG3Sw7OEnkOvt1nFQmR0vZpzl+X2Q4XBic+HV05IYpJOn3rkZnillD3+9O5pcfQ
LljcWEMP1vYRq7CgWPdo726oRSNhuqcnuPQ68LIKfZzO7OmFJYXZ+2/W4cgSSUku
yAzIjrX5ALdj52cV+nrnmk9vVZl8DEdnB8ILoqeZfJwZpkHXo6cM47e007MLoZVK
wpk33UKuE5q7L4nW2zlNbLn62DrfX+b3EY1x4b8sf/cfP/+/Vmz1ZLjBUvly/20Y
NDE+4G3fPKK2DuJyEF6qD7/lSrVEkGT2qIv+4UEPHrKy5zb9o8O2XbpGgRuiSPtB
E8/vlozrifq1ztTcjggCDrXGwQO7xGsDb26g7suL+Fo/Sd3N8v66EFeF2DGypOXF
J6SMPMvf3Wv5MOrVi2JDOOaBMhevmg5WjfqOibWPvf8Me8cNP+/KPyf5N34RCOnD
5M/u6IJOsCwe6uZKLSU+TYRshRRdkLjhAPlCQkZe0mU/2a5g1hzRVP0gHWzsrIFa
qNHKDIdt5QTggwvmjrhrJE4s3kdS+TmWGdO8eAYPXiUlprQRxatyVwz7vePLv1MA
o4X/SN8kOBWSYfbOan8OYLyY1YBIsInJWSYw2Nt2mNcRUZOMafOEupPrNxM0C0jW
mBmaA8JhOvV64pYHeZhYihEs9veSr65fIXm2FcL2dZHSnUrQ5MGRRaF/f0PyeIYD
6C5vO5++ThUaDLxYuHRdlC6SBkaySDcBZ2ZbHZxi099kqCENqq0dYaC70ZspTzQD
OE/X+DaJuG09pepg7LGbpdMPH/WHpbPH8QPAeEEiUxuGxVLkFga95jRMqc3GbYPW
lab0kKCQ5pECyesVcc0dKq70F4+5uTvdI2wsWm9IDeYRD+uL9BWxtQvWzOQXcHAb
Pf/7MRGi0sJuAxp6KtwP2JBUU0blKNJ6qitB/9cAgfWai8OLrhAOmgh6iKJq7ORn
D5RO09I6xbAzHV0DezVwmZ87wNs72yt4o+INh+CfuaSe3x2/O6zH6H5uvszJQSI5
syoFdexlVCxjH2ykQg/QRy8BxA1b1VIeztWFRFJIVZXVG/oA0yMXYBlus7fdF0ph
HDLdGk79HCblqdqiiAzHTZ26MInzQYotJOYUsvPAQYVPZpxT5L+G50+UBnTnHRU3
AZmbjwjdVhCg6xJ7iMCizX2su+wOS0Nb2ccVrYuK/s0KOKWAO5OLOldXp81IAkwV
7G/T1oE/stVUyQ9Uyy3iLiBHMW+aHJE87/DjvDiQvI/9ZzAWAb9k+ZzGbXoej1xx
tjNbpZqzHVbH8A5peBnp7ccDlYTBFK+S5LkxUIdiOyNnh7k32xDsf4S3/YH0fZ9q
wYp6mJKl/JxzP5OCK58RzkS4HUBsTNxjBWNk6Ve3uzQbI8Cw4iveLv0L1LfKCZ6y
XR16IFgwSf2qluYlriFUHgOwx5HaJBL26e81bFX4NfdsWbSttWxwk3YRhMwibvSD
CbOoqy6EHoqll+Wvntkvrly9s00uABxVbSfp3m8e2136VZQXiN0B2f5i2SzTYIwu
xeQMKTt1IMqtutTRDqgyD4Quod/VoK4vOI+lCFZ4Wj9OWKYoSv/ZVAT4GMMCVHyz
H3QBiGHIb+geud7oU7YISYE0Ci0XGfRrc7Oz8QX8PiEWcS2hvYVAnkEEqUt6vqSy
gvgn7N9kxHCakpsakTDxG86tqxD/fWW2wu4K0WcWndbZyKaEJ3eIJN5uZRqZutaQ
WYlzWMPabYr9s0iydd/t/GA7t6ArlmQAwVQAn3O83H0+gZcr3eFx4dU0aqYNAhn4
PdjlmzLOejzIMCrdQ0pVSJOisLRa1O2dsW06DuQ+QEgSMLGRqgdOP4zGsGppEB03
QH7Kkbzp4DelpqCt+LIDHpVw/nMguNjs7OkGZ1Jk7Oy5/5HzsyrGuDdFQt7+inqm
oX3aVY6x9vnAJgR6SW2GyusEffyYtzLEZAPTPcU5N+k9NA5YdMPg18351Jc0FaVZ
A9+ljHBwJfCDHUc8NUUQSgZ6D1mkYz27MGvxKIE2MvxhsGLduQZiylIRTMMCb5jP
C9ko0HB/ttZG1LoGgaZw7iy1SOBOIH07NgN4eXp6U4SVwh0WGbvjJFb7b8zhnX6N
n51rLsXRrQ1Wyt/R0qYSMuTZRTWiX8hR4lwkv0FqTh1+uIBLRpipK+rBT3ulJSQb
eaMrm6I7mniWocE14ZC6gQSIeqOradFDB+ofjr1QiT2ggQxb4bd3qJSqAdIovEeQ
8r4NrgME9o2D+BpiKwnadS9JuLJAQmzYQS6HwpxUlWqhK6vuYdRY/0ZTOF/wZCLl
KKy5nZ9GNPn6LHn40uk2F2hNgGtTknOAIDCnP5CuP57ICA3CP0FPf5wxByj2KoQE
kAh4unjm2cna1zxzxpY6YnCFO42/8xXrS+AtAW7F+gGMmK5Sjc++qzspHj094iGG
vu+16ds/bPz/hAWrlBqq99mBz9p4VoxjyqrF7hDgjDcYrG3nM1tsGkvo3JcGwvSV
QOidZQvfAte9TE18itbLpx+Wuf0hu4ZAs0uggzx2Bk8oTwygamf0+TN6VJwLCita
zv1UYRsuS0lydEL8/phbvux+JCfLfXztlTFcUtdS1nAVPFZUZwa5QYUiCBJuelN6
uysEl3cssftRa+1YDczo6Q3shib4cyAY/kNrVyZ8fuWr40zpYAHpL/rwsTzRNHGY
SZpK/vgJuendcjKoFsuPiUv0aq86fvjwQSKcfqq7q2PzaMzbLWz4WBwCk3Y8Apmg
p17SrcP9srqUgKQ2nT3ion8M573yMxtaKLGmligQWS+d26dLXTKgpZsz/VA1HaWm
tK3BMPs1QdAp0H1qmTw/PUT1G2esP9XAEMLV/eWLvoFMV/ZIIBwFM+4CDLqSbMOh
RfYtp6w7WtMPgqXec9deD1mL3TaT9iUSmdD7xgGgOHVuIlF1HgqJVI/bYdZAgB3n
e0yKSxFHAzadiL2haQ58UrJcl9ztj66DZGZHJFbBUVLAQij29eZ5BhfhVBp08dsM
3DToXm5acFMCAQt//4nVrddtbBIyJeXzoTrEsXg8t/BF/zReQaX41QRIruNAFysO
ooVU9M2BZZfbwbzPH97NHMC0cji9yo1aPR8rAtHUgGlLrCleHuUnUwRLSQxxUYxy
KSANWQxky0+fCwhtXohGV5OYDU4k2s1637WvtA0dPMshrWWDd9D08qDw3SbHHuYp
3x8f4M/1o1qDcJ3coNVKKNpKPhsEhIC2VQeKVeXkvnxwm+iNGWg1uQ3UaGVv75xR
sygzi+92fFTt51AIi40G2Nd3r0oKb93jHBk5XVGSlY1+JBAsRaSJ1cGoed8KAz1K
aroK3vJD7hJkji5mPBm9XKwt489HslAlTcl6rIrMqtTzpgDl95Bb5oWf0BlqzG+C
hZYzagO1hUO3chfSqSzy+WZuX/B34tv9uemTy9V4b0UOZAtz6QHYQAO2CCmmGM9/
g4KH72GqLFSD2aI3iVO8oixv5AkZFqx8hDexjAanW13sOxsf0C+wlGqwAw5OLdE1
PsX7gr/7UHdj+6zDnOqxTPg8vN2CJQR2EKJIKphQ07zeuNsCj8tOKzW0yu2GntsH
QOevR71hkGu4MFtcGPbBKuY4ZEOc01/D8djoS81nFH5heEQfUERpQCseNTnvL13n
lpz1rO2+O2KldXZKlQXHnhIZNT7W/ODQoRUMNyy1sbGD9kOK4XyUWOtvmnKlpyJC
3RMET6o3X4KaNF9O7OKV1bC5H3/DPflH4yicFtFbisl4laPUmhlHm92EOgAGbd6U
i3tGShn/r8qUjNNeVWsthxMClDdw6EnbC8e7QJi1bJb9WDbjmv72oL9QBAvf93Ou
2JzYi/oYDViQKILW95PspLPdnyRlh70E8xiNPnI9naCaQPfzl5wo9expA8bZIN0x
iM5V7ugCxprOY9N6zA9AKnoSDxvbRRh2kHir6m54wswILO2Y5CHOa9PWi0QsDvvo
7h+cvvsSRwB7yaYFscS76/ug98bVeQH/KtVBMn9wNnZdQy89MXxmP1hG3Z+rrKKV
rJlyhgwkaV9dUAazNL50IP+sLSb4UWsDIBDnei+uc76Xdtvq0OKDTUfrpbkcBlkg
CX+qH+1fwZ/c286MJ2l4TIIxDNsejw0fi/YIjS4RBmFP3X6lzOouQJhVI6g0SnO+
kPrtaOUXQNT2RqXkQ6gx8sYnpI/uevLJ8ZT+fKEJQBY45c4Nze5Nf0fo9P08FmhW
P5kyDz2717MgQ29+Mobe7Hh26qhpzvLLucLzLDWaI3qpTMRPS5yjvbYdxASzxmed
LO4fBw7hDea2kSZvioBZpRzjO8y5vRgU7+ZnzNGxpxQmA8uBihMv8LLQyzsbvkZH
2quBV72i9aWq68UIlo/g9rEIU/Bejnk6O9ej0Uo9RjdN1ghL5TdviLAL69dKGuA3
fGWm4mfua7/98kuJOj7vnP33K2Wbh1E1EXc/d64IZ+mXtXQorz8wRdV6hYxbFm+o
Pzp2pOSEUjyNj0rYHIogiLiVgfIY5KdVBx6DaqkI5yCrScsl7nhbZ8t/aoe1Sao9
YpjmBVf1RflalsOCA0aUoBlE+aKVTTjSKB2Dts0+I36R8G7D4GuNgMefSKsJQOQk
iSe9CW0/a1ZHO8pt98dWYKOUmeHBoqqljCfdjeSGzj2YrPtyoAi+ZsLT/bk8Vwxz
GNZHsjMoCQJU70CoDRVvpFZm5/LStPuaJmayuTTuN1JDuHUiHcD3yV+0ph4p13bX
0JWgiKu0gyFnAyzCnwTFeVAUXzIGLUFu5RHr+Mv2aUResl0wkxrdfYAns8Q8UPmv
QtwNeSPwoNU1+8EIB767dQARcqE20zY+het9Gc9u6GAp6fxnzsK4UnzyzvcTgD2I
fCuv+8PVKhB3yI5n9yPe2cZfRzaxC2RI6DpONHpgRIhj/Jaa4jqkqYWWAaB1HFrU
aXx3n1CKOILbO1OJFxCNc9zI33G8Oy5Udi1bMBq3Pi4VF/ru9GI7+BWuHoKCmvB4
WZrgx1BwJJY3plTKE9/d/nCduVPNqlOzT0XqswQ3QZ7lVRKxoDYO5Zq3XNiYG4WG
Cri9ceR0vWspCPlksc81oWLKnGSbFk2bHIjNdC5apeMI0P3zQxCe4YWyVnL0xCht
TvnLtWaSLgDyeZvi3r5JNLz1/RTGIlmt1LgjXogN6tn2zzzAAuE6ddCqf69QEwke
Qk5o6q9HUrue3C/AJOa7K/+UBPfFoHJoVsPNthVlNMIIXMG7pjpbmcSM+wfzdEQl
Fuqdao21XyLZpjMfH1dXYZJISv37m47708DwMN9qEGQzog45iLRdZaAq0ABSMD0n
d062+J8EpKAun359t4T9plxN8q3wHEh0h+yy7f3hiC/Xwoj5id9edv184zJ0dgQB
BB6CtZVI0H/nnMS7X6QupQULgEc7M4iyLyOcJu4oRqXIVKLL72VOh6MvQ25uJZAQ
pqzF2/tQmVIL21cz2vLUcGv4x9B0mHC31FNESWIUmcw+z8Bmth7f3uPhIsMC1HoL
5fwTFQeuY1thuvZjn5Uj4hjhsRKfv5FgPXFLPDkZpnY67nlCjI+quQOFdH4sKPR5
OjBfLo5uw95qtXQA+zTbvu20kAGg1GXxzTe8Wj/YfZ5qRz6OiGUNr+dvZxqfN9Oc
gYq+ILJfjqK6O5fdOg7rwU00IP2KfMKXKdrzn+f2FMIGJENkp7ok4cUwnIWknjOL
vPpE1W1MqdsgS2Zxexhb2MJQcfqWMX5kV+2dyOw5Epn0/NlLjBea1/Y+6rg7/XUk
nHDroNPpXtOwwwhGsEn9jdEzbjKrR4AtQoh8PCWQKLJAUwx3zldua1iL7MO0Snz8
38/gWD06JSfz0NW01Mbz1sIK/MzSM8ihIYBphRq+K9zDuOwfJG/spv2SMKsdZvX6
EpQnHS3EJp8Zqj83ihwwa2Ia2HZC2MH0qXHjy3g7RC2UzQvjNxjHtEymcqsPEers
kTFvb8nkUNFF4nqP1STaTzYPIP5HrggrjFDu4TTbNTlGKXDt5F08fc2wWs+Tc70p
YUtfT/tt260S2QSycrB6aERHrIzE+j5ORTgQXc26c743U4XfKvTwQSVYrmnpbviK
TJkpJgtLG0JuxMQj/yVq0offX6UYC2ilCHJ2V36KBxaKlEEP+nipe7OOr//hgIG0
w6gNYcFrlxp7pt4iR4eJjFyiW5pTfjvMS9thqIZ5CkUrxsMqEvSvwtrjh077x2gf
WZSgBbXWA5lTIyr2BcD/vpHgQXEvlOHl904GSLyRPQC9zPHPFNQejb9Jk8BYDAMP
FAhPFzctIXnIcUCiQ5S8AkdB5NeZxd0xu6U5SKiIuuBHjCI9pL7J8wP0kuaBvr9w
+qxUIkPd/7j+w3ic+y3Yo1c8ZQszXpQg0ItFvsX3T33rK3YP8X7M9zNLAAx07aSs
ZBfkFCnRtj1t1sDjKzAJjBN6mf3aK9Y69/8deu19N5YoKevAvtDtaQHbCQkq5dQy
t3UaXalBMacYNPCA1ArUZC7+Gx4TUcxlALVYWCARvRV6bUPMVpFWBWBzSDM+BzKE
H9kiNk6yANVweqA/WB+3dUKZmoMss9MH4QixjYkn9YdHQHTpeArr1893aXs8c7IX
LaC8uac7Px9XDOvBWUT0KmG5muy9TPhZq7MN9xYT4d7B4klB3AQpCD4C8Q5TiAXh
6aVxJaXAzuvYycwTN8gM1qAV03X2lO9987aQLdp8q16olcTf+m6mqcMjOuRACo9/
hZ0PvqDYiqk38KJAjEmFOQhUck1tdqUu8PRyV8lvlpaEKZBkSztYyVSgPtBbyXRm
MxG/KsUzb50GlYbC5xy3SpthzWgYWnmNk/5O5nd+wl+Y+izKQgsyMjBL6s9z8D6L
0bkaIJaGYkgp2s/ruLBIpR2XTs3yBesy3U6uSWxMO7nZCHCBPg6nArukxtxoh7uV
JmegurU/KKUBFR9RiKi1pU4Wtbso1uPwHfatxLHhXG84QIEUMklXsKdUGgCgduvb
9QLbLmbxIhkqD5qR0YC7R+u191aMN/9cXAzTMXW1nNHhqTfiHP5a6DZBkqQUKydG
vmZK6VokC0d79j3psCud48QkjHxszfkus/BXMZEtceXJecwFCKISJq59hSQsxJ13
NTbPUajzDPQYVt1ZovELEvCAzieZInpfgKmW8w+rokCctthXI2EB+Q/Bzx4z/Nql
m2Dfl27+qSMYPe52wBic2jTbori4CJKZRgNaArjPMFSdLEnkWgd3SK7Z4kHue1GL
XBdOOaKULiLegJf4gNXuTNM+gjtbm3VnZKQmcTTESLPEvQv1kezWvucRLJ2f0jCf
FUknyTgRkf/G0XPvPIvGsRFAU6h4l/ELpaIdf4bHvT8uSzTqjmlyrfU3qM0zSGxk
ibIttiIcMhsBv9jZUzyRNcv7ilEUpKbOJ810tlo7J7oucdog/41fIP2Y7PIUTg80
d6uwSj5nYbjvQeLjsX2ZJWS8g7g43/GFdYld7ErwoKIH9/Jb68bfkafJZorJSMwI
i5XGlc8flE+X4NRlZfmifgxNlwzMFLI50FdZ2jr1lZocEmHsQAh82id1h/mllzbA
kSoRajKgnbYFXBjLYIH/kD7W1+3E1nrGQEwkIvIO3CJwmvA1kevyq1mJXV8lk6p5
49Jr/g4Gxo7tZOevjYk6rcPFxxqu8V+UMYWO44VZ7RTgRiYIJOYURXsOKAn1jEs3
E3yIY3vLWv3ufPOYqzjLWMiXtox1PEGqyA1X0RqoRbqmZUZbj+Ay1tF77w1dZxOM
M3XP/qlzG4YQ5W2g1on5tp4VbYZDtHhpx5suldOp+1B1dh/ifXRkmto6Z8roxYLM
g11jvfKtxwprcPuEz2ooUnjRDw/qSAA1SD5Y2M/1uC9co5Op2X9Ch8Re2LSwvdVy
8Y9YbHMs6eFI5ZcP7/oZwhb4LqrW1QA9fTfgkK/Bgnac0cOQHrypbXWa1mSqeeUi
T8zEEI+4abPnt5etbyT7g7BSQH6yKoqHRVUOqw4M3Im5gS2jnQsjvHR18j2iTvK9
jUQ5VLKmh+kM7iTgp/qQmhBPuObqIcuJEUgjlbVCh7BmJO3uyAmKtZiq5y2vCdNf
LiJU2r+jwOeNfos5rxNtNG+egoUlNxm4zJIxw5yqTXSHrZdJN7ssy30JlLeoGINT
lRUi+iCQHihRM3JTmXYobSp5xcWK8C5VTXxvNHlO15YuFdV1mMss/tfEJMbovZsy
nKiJp/eVLaeSbfCdBTtPDMesPjmNHEl8/6Ft+4UCOpHMVutOPpJ1Y5/UmTSHc+LS
374Wb0IZup1MWkvZ0WLaI6NJ5XevncD3c8lek+BAzNQviHYheLqCVUOmFqcD6R2I
KQOKFwp17KwhXnkpdrYqp6xDB6fbWDnVh7CDqJUYif27wsSZ2eh3U86ARkBHFkTs
6pgeby4y9RyXRRFLGL3UCCND4Sf4m2AJAndCa//ru5dGkGSsfiACvI6G45VEdqwq
iraW/6RQw+epjBmTwUOkQwsDU9XUQ1yDEcqbZram4YMAzCsvcnneQK6zeAWN91iw
3HnXHUx64e9/3YT0ejKjrRMW07F5Wd8yOVmNhyq6wUrpnPlPUhrNoMhjWidDuGIz
p4oYBn0NZ8iosh0a0UiHlJ8r5ny/tBf2+Eehm+8RBGXVr02UDoi1uf2sW++b/EF7
X2+aoG/CJLNiR3mx6hXbckeH05YAC7uAyndXApLaW8iARvemCRNsdQhJzXj6BrRI
hhulS4vfsp+Nf/KxPvw8NrO1YGoRWASoH26QUbzc477fAvr8lrPLuiGVbFKLQnU+
yZ0Uv+q4nKryr1fkz2wYlyuZhiJdI/igtNtVXwpApEFvY7BBX6bg6kh5VX4FM7Cn
qWQxz8Nb2H+sSZ5NCye8NLvnsQObqMzgcl9d8H48Yq6ATt5VZoiHE+UL0FlDlJoE
00oCnSVz7XR8/8bib8s8O+ht6jp8xao5kJa8sbKpKiYgkYWDbE9fB9Q/bRNCHDYY
qbNbUCDPnSzKnR+wZeYoxa42N3YDMlc8ukn0RZR6Wac3cK5yAbT+rz8nsY/MKH4K
tTVZyDfKo3h+7VCf6jOUuHojFAiDk7FApaIHdIviCCDHDwiobs5qGENmXxK+x+aU
lQfhmJQ8q7798y2O69SxbCTanFfONwAovcX8/m1TBcLg62jBjDC9LQ3qVBT/gXYV
/2XD78NXxvPRbF2KofLnL/6kC4QSJDEUFuPo+MMlvnHxFIl81YrbohZTeXAVJ0oc
PDKSC329c9wvlalidMmcaxW0Ds8Cd0opIRucCjo9oBQgZJ2F6gqZ5pri1ZN8fwjD
8oMT8XZFnFB6xfjeKVdNAaHyqVzZcGB3VZLO9WvpmR4Vixkgve4R2HUdO672sf0+
FoZuOROEQ7ODMvzA19LvlsIwk4vfE/4KXB7j8EGivkOjg0PR0RLccF5AQfAv1isD
LvGys1bXq90HXcC0U92X5x8Eb7t9+NFzjvk++KjbrNGsK6IfM9ZUSZB/INdMY7RZ
TRRumw4nsCHSqdByEjVZBaumJ13ZYoeNsXS7Du3BlXWXfoLOGP7zKSWkv+F8VKKR
z8d4GQEjaivmHRsRmeVR7FbrRR8adajhL2OpWuzNf0RcbJCLVPeMKyojtpGeFGOT
QB3dUfnD549QUIgE88UEoDSb26OAQ5fdbvPJwRKEgiTMqiAbfNsbPVed/t1tJmh/
w/NCam6ApOnaRajCSICym7Rg+qGx6UGol8npyqq2p9CwO4wsN52wwyxaH0/VXfOM
93W3RTyd3DpXqJ7q20mB/LqhYuNDioHWsgZQk28OR/fPU7Xfoxbf4UgtNDIGmIwy
MyQuogNl1RPUYcU/EGk7Qj7aAQMA8pGtAu5PXF4EQ39MXKfMQ9oUNpHr8mX7Vlj4
OFAA6XDwACDrTRwHTUAFhyRrRcJlQaqdP620GT1nsHeAv7ePZTpADpVfPxFVmMrZ
3cn+ufnQAbQKJjjS9BpL4lvZQdtHipJgtFGGx4ACbxPIjEEyfvJmLwKjLf2VHCW5
t9SeXQzju5Ldy9ZXLk95DQIJrUscsqJXMv9VndT2uUNCeNVpxFXZdfbCVZqw+mil
vSQWTSgeM8JW3WB9WTDt0HWnhaVBTKL3x3s16uQS9wuxwewCOLDQeontqMKJn31H
+sepK7osZuLLKzymtIGsb1I83t2Dwx5gMh3oF7Kkhwnf4UK6rCE3mmkgZTDDQINZ
yBJzIhn8v29bFgLVbWtROuWWyb3azljWugD0MjFtuom1LeopnNx6cq5A8+W1yL2X
zDZVjT2rnOwkcW+e/pDP3AAc2UOByxi6gSynwbNJQ/ydKc4MQWtF0RIfZ1TypXxy
Dytawt2zm0O00t5nqQNmRMu3uYljFBUBaH3hULOfYinktbY2htLX1N2PiVvnXR1h
XVFbxnWvwBlE8mdJ9wSEX8turmzcQGV+YbXSuUEH1Ob8wCPzgM5XgMXR1wSppGPA
yO+5CoojLnzb1fC30MNOIPGoLSjkfb3/0c2nDzYV8OCJiu0tJv9kGEUoa9rhaBYO
SHy8GlNvGnpRgQACrg6hZZM7eFGc0HN0ls1kTvg6RGauNZ+3Je/MJ9cUMr0UVoGi
uURSn2kZVZIA3TqXsOo5Phiu2b4X1DaNnn9gPn8KTve6FpPykaH5SdDluft1yI33
2L1Y96PYl24cZ8tZZBFho1yY+bz/6FgVlKBevstiWyW3pvGUgsFpi10lLBPIaZlZ
+PyxHuJidbQg22Wzhi3JQmT4cBWvKipAZ5G5cuda36k8m3gKvy3cTYBLzhnMxpvr
eFONi7X9X3x32CPPEN3B3H7ZCSSqSsns1o4QWL1n1LtuZwr2k75TpAuzKnK/tsE7
c24f8JbCrPyqcxWaEipjzwviN3Hvel5Fre/TzQAA+/6u73mDXNH1B+eSA15UmeB6
XlH1kNY0/3kbw/uGDlL+LGagT25xstCnnahN+FjFj9uJ72wdmW70XIGhd1Ng2jDp
tn8nFdEd4WC5JAlWmQcWCUMyGTuBouyTTiYLcHKnKaoDn5q7xDv/xNcSVjCQsn/u
VPIweORLZ45knN9i0tuv/LL/0QiL7NMpqL+s2gzDoGRJodoQQkPGyeqstzI1qPuj
YDiGTcCi1QBxqE1qT/t+5K/WuCqaYv9NG+66WR9EX7tKa99xko21hV9oAssOJSkI
5DaIha7LvmgrkpmvNLSPqENB0EaqrjDmpoKinqQ7r7UEC7x2SzpqR27yj3LOdPIE
QzhNRocx/3WZa9d9SHZFABTqYPR7CdVBG2KaxLmI15msvu6F7Bxk1sT6De1IynEM
wpii8rmOFFd0ukEqPb3Jrhhfzh0++ZW33+s8nfRQmDg2QvQS5aonyJeoi83+8FJt
Uk++I1PVoTyJPo9R/ayakz19wyCnFozSjoQ/qxKRPMjiYRoFgbPBiSOZdoXcx8ln
3NayO6V8xrt+wh2nY3Yjge1Yl/hqgNbyhFh3+oXc+H3bb+WPPqa17AIigQFXpv6w
oxKt7Ji7pOmys/7o4NDjRlq9JjnallxrevW/rQoxiDo76FxSW8Biwrqpi22Wd9JQ
jnZtJsdGOt/hgHXdykmg7/B1HraTMVubbECLzxV1L1PBozSnlVv3Zio0MG5p6JGk
mneDomjUyxBgzVhWN4BQeoYPlPRmY+g+c0OwJ0x+U08ZsCwi4AM2bmz8quA2hu2K
z6HcLgTlK5IpkfB0y01V08zvGTi0QSadRmXKfhCOFrV5x/UTtzUEv3b7lKyUPmNc
CDHA5twMjDEGo02Ur2XweLWOJv9rbZiD4JOuQ9WYpyXkeH+NyK1ifrbR77qARFL4
tMg+JC7GJcnP6qOXtGmIywrpNQIis+Zc8bPLtv6FlJsirevrUMnqQnsuJzPdo/fW
BUB8sGvZ05BfKOPzWpvXqDdIg+K38kF2px27HiwgW+d9Nww30Wdsi8nKqLeTDvmU
4oKVzO6vld06IegpMLvzKrjVVmD/64ITZm7ahwmFDNGDCPAJgdDeQg9w3Bnm4Ffc
ZQnbqASoxdeo2KEEISYXci5Obad68s8uhoX/WgHPZIMdyqoMQyMvwLdSQ2N9RZlU
9hC6eAz3aOiQfGi286eLCUwZFTBSLVYYYMbCUqdlG4oPE5ZxXxXvae3HCbNqWHN5
IxT03C+up+zgKstwCYrTkPsD/30wmrn6sAphkfPhbq5XV6H2azKK9FR9W5JbX0zI
kotR6U/+xT0BQAaYCIt5BiRUONZ9zWAQowQxQtdNv3CDZNUPeska2CNJFH+Gok8B
VDDbZv88SWY8FB2NkPMv/PYVbpdD1RxG9kvs2TOOOaYFe3CvBlFrjTxAPKqhHGhc
8MzMsvycZAd8iBpW7uDaqwZzsBdMzfg0eLeOSEOW4A+9alzss7nYCRMMNPITwKDH
ili0382Kw6ZdUi3lMVi1Bs2lK5W6LVMHOhPnKP0hV8xDJ1H40VRQqHAcUxWg46Kd
u+IV4/P2XC+gABqatE2UMuOiWZNlm1o+CkKbzMk/C8yJqJt/r8Q1GoveVsA9JoDM
nKwaWurX92G+iqywe/i1m7x9b0XBbrodFBQWzrro61pTdctRYD+2QxIhVy8ybaka
ZRzU4TCo3zuE7zvVpQqPjZoCQsKdZhgClaqAAR9L1L83H9TCWCsljCqo9SIzFvWm
edaydpCOrRw48dLtLy1d3h/Y+ApZdPpEvFIestG1obwwfFbSyc5vr1a+XsV8YoBZ
HA/WQvzb3GMq6NK2BiN7lhakNHCbqcJFFFPIaqXt/eE2OwEXchKmNbZ6qcMwIT72
Pi0UXLfUnjq8mMCj6eFRDozOCJ1Bdk6jQCzXWrXAuFluLD+U3mUJWuVv8MRX4Zps
m4HasDmZhYBfoMA/cY+TwQAGk5W1luND/l+v/32ksoFPvOBTt5nHRrmM6rlRkv9w
reLnEzlUsbEy9yu7Duu2bx5NsaOgfbbkT4pYxwd3zKZJk6Xzk7MOckMKB/hwsZJS
C/xOAoV87QMgRg/OO+se7oCwURmA+Hxk9C8Gsbi6o5XB9Fpb0tFc0+dlyrnxQ5CO
xa13j0B8fNwZ6YDm7YXbSERaXQyVGefoMM0/4ZhNExIzVjMms3ZutddIRSHd2GY5
yFwPOb4EYD4D/Wac0FiIwScyoIsNzAVSaaAU8ept/OlIBurFZ1bqmZ9cqWWBBNEI
mDqsU+enIotzWgDDy9etjx6oMoSa0TW+SDbJY2jahggjamUJRnvbiYHcxy7ZVAWN
oaDEkCkvYFfpbQEx6VxXVAbxHAnbOqWuydva/JB2HLcsPiE6EqLQa3IDXcBPs4Ee
qmepsftDTXYZpjl/5z2+hBtCoCTXSy/ycBtbnCtKDX+ikvDMonF+HGJmO5TRkbDb
cAL6F5FlxE7QK/nY0AcQWZmAYcfykF7Pu/Ubm/4wuGiRn5HO5ItkYeXklvlkNJP2
itwMaWP4bXc9TuRULPqu1ka3QabecjL7rEFrdQt8EkQIhqbplaRT1ZZX5W6Qm3aF
odT75rJOgy+PPSvNxPq2ir6DfxvbF3Rsbw7Fzl3Jgvi/fEwwZz7lZEF31BeVvIHc
Ae5vfj5HR9/EdlsQfhii6cNa92IuvoBoLEaXFeGW3HkcBkDSA+O0+gT6OnErCxF7
3b8VFxn245Opx2F7rEMUQQycZKmkncTfSHXlb32OFUvbOQ9wWK0vYvs7iOhAtUQ+
M6bmXMv8dkPe0tTPRYbX15swXUKqzTM+Cc8FdY8DLUvgbEGRE79XG672qa68EsIB
mwooJw6/M8yW5LrIEdxQ0gr2ioOhe1WVj5DGacfWUoWSnclpTdqz+tD8/IuN9SEm
+ERubXzqoRpIBHEts2sjwxfxsSyt2Ek2yK8cJeunas0LWPi2jN9BzNoAKHr6cMIS
BvOKpKuT9lVqGYTqZJILXJ4k0jpfuy8KyNdnJAF0PET5svSLGcjeA1cEr6AXDJGS
ABKox6DwmABsZich+Z3i/avj/wMhM9z74bEp1QuTDfXfe2/66zkXIBkYS7BKF+XH
9g+WanjZx7g+TPCKDTfAIWA5Yexd2Jh5EazR3QnrZ1SiNe4rEsPGUqXtIr6klL/g
yZ24Kiio9DrcyurdACxrhlq769F7yX9VUtgwjHo11fdxU19Rtr8M7LjhGq8lgY+N
20voPnBuuCdXGCcu3sXNmILr72nKubihFNgXPWWrEs9Qs8gJtaYzE8ru76Admyr/
cv8WEDnD6W6YMSOMN2lje7tSsALHSJ+xSBX4y7FLWNqqGBJamvk1rBCR+RW++kS5
KPawt8epyZGLa7XqLH6tCidQZB8YYUgEzx1RDDVGygaGf4XoRMkBa5fzXVGIKnHg
WSgjWhJCHj0uOue/qEAj5bcdQfuuSjuaTrap6nPMJwS02p9NLRC+J6X2R4oXPcs3
71NbbZ9Mtn+D0YadShUFneyLuzsDqwheqvSIbSDC3bvga5bgCdElc29fsk1PVzML
bIANYdLna9aP+ih2hPtDAIZmEcPDy+pwJlz5omSk8Q9C9+iCAbT1KPue3ePhheCA
GKvUd1ygoXkznJgdCg2+ktLLJTgMod79FVBKz40Bicgr82qNxgzvBjhY8gLVpnpg
slVBV0fgoEI8PMOK32TfWziQmPVx7nv63c34925WTN1qA9OuECcpc8xGJmWW0Y9W
YJ54EkZ1dcoqKq3iUOyM7ZoV3+0twFEvu1xNARnCu8sly5SGTLPgnVxtiqAcyQ+g
Bt6l6JQ9HjOCnDLUw/Qhd12PxMEAgqgBP8VljDi91qb0Q/F0BY5Wtm3ol0rjF3uT
672JrJEfvuMPm+Hso5wevcBKjpoEADyyW/3KpTFy+G+GZ3X0WLr9uetkt+ZEhno1
bDXehhJTqV3isp3vdrMTn8ksAXl+hQis84s9QJKucNW/SqumRyLJ7AnkfD2QUm6m
xaI008oQ16L/0Y6GsHrSvsl9DXcWq4cAxKG0Ck2H3dh2Mg5a8OBLxu8ROOGrGVML
H3u6HA+I/7qkD31E1gLXTr4ZxVhT6hPQAyIHIJF/rlPfCFeHO/+0rNAjldCqZnRK
UBNMsyiDkKZzGMEeyrP2KfkA6UqI8wSc47JI+yr/XdBIy19lBqG+/wFK8CEdz6yE
2WhECLze1RUDY6SuMY2HFLUZnOvXaSdTzOlyhjS5wGv+kOMwuZenoxvvnuZLUUog
Ao0HWdPhRQBku4tQ0R5CmAbdDNRUK+/ntS4ghMMmdTv6HPEP0a5ZiPuWiUpmtNjd
MyaPV71aLOMOBZAj7avUXvZuGOR4ozo3fe30H32Kp8Usu0WIiNayN84NmUK5lH3+
A7D0Q+XnFPipacDcN2l0klmTYfMejPjHZwvL7VsBVO+DlEDFhB6iHy4seY92r/QN
83suqgj/PVlH+dJHBxWe1R57bk0ofR7g5pdzSSsYQx4HegzF8g73euxGr+Zo7mSI
bupnMFdINx5pwTZpf8wXiwPsuYU59Cw8P+gqCoAiWW2UKO08KomEhr8JExsQkCxF
urWdRpdVqjoigWWWy5ODmh3b/4rNlKuG+uHswk0DTALLntFhUwM3+M3ry2Z88ZTP
0ESWeulUwIDmPmQ+cg3MHXhSm6cbIJ5bQVjGBMAJK4tRyeqwJVp9BJf8oEqkpJeN
jPyAVPSk2Jj+OjN8j7WxagtUDTtJhCDMtWDKRPkQ+TK2M919T9hPg9f71Q/+LHGv
LOH56XMfEXMp05/eaczcQgZz8MS+EP2WQJNqYyhPesny2KDf1Wue33gxf77gLdPG
s9XmrneM63sK+7sSU5ywQR2Yq7sh1AtJHt6K5YpocAkuotMOF2k2qhABeoc1eUcx
JoeSrp8XtDdqULP8bjg5Z74tYUKOTZ61wWyVR0iJth4UMP4J0LmgMNATl+V4yaZc
O/CGpIP6mDiv8NURZ0UN/F9sR0cvIeqtfT1kw3PXehqYVvuwoV/wyUwa7VjXuN8d
Eq79oyH2CWKbSTUwUyet7NVc0fhaGj+cE8yVeVuzXAP2+coocPii4h/9H75xpKYk
6HOr9mMJr8a4vtlx5NZVil3uNE7hIzXjAUxL9MDiy/z0rcF0TYu6X4vDdRtmG2NG
8tTQoT9QVG/koxJsIqv0oyKUqyR+1OzV0PoG/wV/b5NccyHT4lMeLWGDkJlHByYc
2/1kFn7tsHES5QlLeqoYSSWURtma2jS8nJAjlRBXUAumDq+YWnkEXXVYeZQtu0yM
dFnVZ4vJ1iCd+AOpfao4tqyXqhFuv6dKoYmRFsymsST7+/EfSznO0xzOXsLNiuVl
H4L/iDoTyFYfdcfQKbSB+DWHeA5OE3MCsJr2C0xylz3wDE9cJDnL8BI1+u2athbM
0ajOkAnMaxJJhaHH00At5btDHCL0Y9R28fINa6GnE+NTdt4m6yGdG1SU4yeVv7XV
06AXikytuCusEj7I/MmoqlQ5xdHrv/Udqw9MfT9USnMdVwDGi0LLOhQ79NYgTyfz
nd0yemyp4XBiQfUl2pMokfnchy/XLsElV6w4nd9AvgagwP1dHep7euX2p4vudFxM
ZAuZzvN+0V7cCOMgG7QLxGPPuyNIJtwrEhuiaausUf83nldr7LPO9E/F4d/sxaFD
rK6bP6ZiBb2L3pN5PYdA8+bYqr2kkikXopxJgmHxG8TjXU2/JzU9LZpYXwls7HSd
nbbOybgah5/HffsBZcaibSSYd+OcwThgE6xY3e27MUTWb1rEK5LPLrT3yjkI3TtV
WFIJK/sSsxQxtWta8GbY3GTJ/bEvqgIs/d2cIgMWB1xL6RbQ0Mh3imPWfyy1Ivcm
3TNYxt+Vk/vc4LDtBOJeCTjlOlO19zBJsnORR0IelUETuNPkGc96YpJWT6hJNTJ9
cW7+4zhMK4TRblQmemUxzptfXtlQYCtsIB0HQ3mqrkXPYLbW/FPX0FHpMTHFYoo+
otmyxClKCpabXkdMyIscnmrTv9e/lts0Cbgz/a6iFIYHlBXyQtidpOLq8hiEO77G
x6xkqS9wU0qjp7koGfxTXaDW4PoQkzb7rvAL0pJ/LuW2cm9MoQ4niqFaKHd3tVJP
1Y8BUtblwxJBKuBSMAvm6I79jpOYN3AfgRD/zyDXz7uDfaaa2JDIH7L12jKn3fnU
BMw89JcmrjTXBWANIdSF2UYlcnrjleb8g1+/Mo8e3y4VM4Ky6l4ZqSpaiC4mYxMG
cvFrD/lJFzN0Iy1wWexvqqSP/03c4v72UiOjXsqiTn+NpBsI7ap40c9hligZvL/M
2ii1jZEqT/LVaIM+BFYNTowDJ/oJGrz+wIZAWIKH+9mqUc4lfQQaJoFHc6cCsj5R
H/Y5Tihb05CH8XWqe96+zg0eZ6gMKKc763+N7OmGglT/n7ogJIbfmCGyqX/AyWTE
CllZRfYyKQXswxgb9YOF6kzIV2lyupWZ1IGBF7Rev/aPtmSOLqrkB6mYiuKeVskD
7SQZzc7FtelDeeJC1Q2wiMlgY4kaTUzatSPLuF5beISqGLJLrUahYrb+CD9FxAL/
r/ftN+5OEcMCJxc+onz5a08Q46dlwGf7O5b3/hHyY1rZV0u+uTAJR68ENXEWZL5k
lp+CKtQVeaO4LIYe7Cm0iOwdg2xgmeM5sfM52iInk7UBSQ2hNUiwTBe+7ZErKXME
JFd7beqT0VQ2NPHbWSuFUXJGVN2uZ9FMW1EPWMrdPhPJRnLFAunYnWko7TM9KT9z
RqMt2XRxlKS2Pl6DAW0yzwAUkv94Sv8/4zgFaJLKokQI++TKJDYBQtBKKvkqp5XC
BylMiV8bVdbHM704zH1bZzctXuE6km2ysH8jinqi3zF+pUrWPvZMdgDXUZVxHr6v
feMdbq+XpUz+3C0YQmN+mLg4XKww+KLM6akkOlHgONz4xiafYMONAwFGvZTBeOmH
tZOm9THnNGFL13K4RhlRBLpi/3UoywcoOtepaZihEE7HG7F0jFyhqDbM2iONGDJz
MWeSHgbtJII8ZgSw4PFrjwU3b05MFL/EkZ6m5Os6F++qI9RgpCoPK1WS4Z6QBQ4F
OHm2QHSQ9+53enPKwgpTljLaga2WRFyjKlAqarBftKWqrqzbEDRjiu1eNp/eQU+3
8wce7Ru0J3Lvs7UOnrJV4WctBpePFH/E5sAYrQnfGiUFWg4Z7EgnGGdOkzs93vku
9W0NNDYz047FYu6sZiO7zyOeHMt6H0aowPiIOrn1sXnzfyBKMWhrK0bdoQjVXZhX
Q/hIhpOu+3pVUC0j6IvVSZn6jQ49DUsWt56qmusxSRPESewgrTfxGT/yMIna/kSz
J3nUdEMB8qJ6hpVjaJtvgq7ZGbk1cr3Drjl259/azCJ8JiNb6+TTDNVw4poN9z4R
zZ/WX378vXWBCBV1gTis3RLaCP49Vko2ufrEiqRMxSFNrT/1A1QiDEqZfDKMjEPW
2Q4ktDUj1X9Zw1N0V2nZusyH8NxEMgekLOXZVVf3iNFxktMil9gBzphlIFd7XxCF
YYsRDcKldc+OiLvqcUAFKzk84RImz7tRLwzVtRXv5bDnavM42okyAku+7JtTHm5T
yh101b8Oj3XGbp0Fvyq6SAAoRyY5kObj6FhGQUKPHUlH0Oj6JddA7/GLoE8hswO1
mkHH+o9rDpjIm7G0yEMYmUi3veYS1E/Oygy8S4mPnA/f5rbSmc1+vQy5tiMYAZM8
oKOKZrY4dIHL1nW6OD07KvvaLksZEglWd69qirO8henzXxFkTyZLGFnGcF7FP+yL
Y76uK1i3ZRVuQHseaq+LsWDcevfpWX12XpkHLtY6vcto7RR1yb/dCyAB+xjZVq4K
K60AjB1RzzpkpsdANS3Dd5B0ppBMNLAbr02MQdSF5GKDieYUELGhCgfE+b11KQVX
Rfgdc78Ng2mzhSRWf/1ptjx1yhuq9Psxb4XV7vaIMF8puh0+rWcL1yVYGUP/MWom
e/nd6VuxYQldQgA8fTgOdNvySUY124kjsNVt5NSWSWhG8utivKCV2bQiOIH1SXSR
PmMLRePM9xXl27bps2S4SiuikiU7ggF7jzX7XNqzxYdSF2QfNYloLsFsaxpbFdl7
64/KhFJ9X1vpjW/5lFPBCy2rkRaJmamPvwopUJnZH15AFfDvFQxtwOZyYzVOuuDm
LsaS40pzLHs8imtgjt3DV+h9poXV6py9ZorV/s4keMcRV4QPmnmH6kQ4AbhnWScH
MVwBNwBwYYyGvag1jqn+UQYxI8QbKRxdvO1TWjYPGkTWP382HaSWmRLBLVZAbckF
7TgMkZ72ACNTx4DSohtlAyYPnnTc3Tfm/qVCxMddQ74V/zLZJINxJD+qmmpdh+fk
/cQlK7XP6NH21mY8IPCypLP7iU2TygNCCIYi/otTzzdwE1pnJVk3blMXTKzTlDdN
Ct1WkfDr7R5qDCTSL1StXaP7512PhdvBSq6YOB0O0u59w7BC76S+2ttQODDoz9Zo
WsSBgsqzJKz3Es4qGW2UNvoz5W7/KbcFIZdytJDaPD715D3PSvRQ9YebC8gTLKU1
iKyAoWSAuRn5aOW/n9/GSXJvgjUptzBLFxzc6SAFvf9w+C34aQT5sxE0wZKDpmqu
lNh37d6P63dAyI29Jh7pMJmXMNKCB06FXIze+pF79vrzudjKG/LR/R4sXal8szv8
pPuAfqT/DNvJ06QhEjR1msKJ99OIZ75Phr41Eqk28oqVVaxB2fHXcHf5+EdgHXCV
kRfCuquv3A2irgDrBGj9g42GYua34LlR7ZSAPuIjYCBfjt/Pj4eJdpMi6VGOR+d0
CWil0xg+/DUGMekefPc3v9tOE+nrzTMKdWFFAv7PKT42ZBjW3Lm2VROAOerdHrma
bEVL7571q7zrsF8Go0Ebyqhq8It0MUj3E2V3thro1ejQBEN9Gh7zx2lFGimmvpS5
rwm0QoLQQH6evo0NrPWodKfWRqdq80NR5JZ0AxxQSnSc5TkE88TlKIlxTLT6CFai
3zWN+o9dFmwbE7EHAzfnbo/2W8yqFD8BQ3Fl+ZQe6zgALKljLL15rkaeSGZXVC7y
Yn9hmaUNtIQTgI1apG6zxiSRWhknzP8ZLW4m0qu6cgW8RKfZJF6y/q6STgmPKDep
vnvhpRgbuitpBygkDC1gylKkYKuTVUbajadOgBwk0BSZB0F7eHjnl80UcZJf9Em2
yxHPcjg1Jl+uIDD+i/4bnYW3g8u5YpK0fNBamMhfLiTQKQNe/6YDN8wmNQh5rNND
67p3ZNuPt3ealUkTDmSs1SnustnTT2uT+1Qhk7MUBGYbKJDnYPy7n+mH2eXVYF5m
pvAULOu5DmXSdusp23JJ29q59izTl0IaSBAyFk07W66SqHna8AbrzwFlOaaFprW0
BIB3Zs2l6ZaBnnfYnDxX1J0JaTuinbWOTFFWahp6+Lu+yvst+WLEgwjQTYHdUcEo
U8zPpHZUaSQRFytSz9EwNklIDBkhPXrSQ/WiH1StVaju9YdGQByBU2g6m61DRX6N
R04dD6NfIwhWDYjGipLP/XaFwTSHB5jhfZGxPWhi9bOuLsRClcX3bXi/HdfDzQ+u
mOnR9lEY4I8KprZyst+YLRR1vm+K9s7+A4xwfxXEP1je2X2oPGGXZOjPnlMF89UI
oFgHsgHalT5QMosuVVVcWoXZAERlDXCa1DU7O2AqQOMF2TmMr5xUJEnOVymdKORF
/JsYxWVNQT31lomxFYQbrKayHcz+Wop3cKKoFkiRIKk9MORU/C6ROGBPU6BV1URB
+3yzZH4INnRpF05nwAd2HSLgqg8iP9/cFzQbUUV3xNF9IuMc0huIQ1fdAgL0BnHK
CTFxhMopYY7jp56UN3Q/ElnalYNJJyLfXkDtsTTPNLpqCDk31zEu13ScpKbTu0p3
N9ocLT8maNA8Mj20+Yo0Zda/YLcJMGaU5HY+sBMlVUgnPbSJOMdwoKt9utSv1pJV
Bg+s+N0AUAvRLMXaUAmvksXbFxN3y0oPw9CTup/aqUqCiqw9h7ThHGCYKKtuEeSp
PWtqeaa8dwzorfSjcARFhH6bRFPqmozag4gaLatNtn67Fi1TqLnRQQ/4u5cs2CQi
HRay4rijQBrPRG6JR7IPw6eXiSie8oCNS53ULLkfppruHMtsnyr2trtO0mtU86SI
SByDzycA3FJ7ADsILc/2t2IldaG6MV3KHea3CxjxMGxR0GdUk58AEzgi7ZguxuNI
YpUc/ZhdlAbePLkqB41Nr93FSFeR96092uXDUoPYk5t5wIQMeNPKXn1JXSWJafuM
k6F3b2ifDoFzvEeQ6RY5BZnsNJKTJNbFQ6RPob64TnJMmZv+Q2eMXY3/kuYROop6
KKORKRzzVVjUg3naQScZF3NYDVjYZxoW3slnbLN0TaKLan+BvTN5wVdmEdI85Onp
mTxbvTHWTGAhY40t57xQ3gnpsn8SZGhkCdPaPu21BDul56e2YVt8/Jk9PAPPKGrV
iSr6DF3Y04dqjF5VSRvjx90+XYMZn4FAxsaMVx7JH/c3mvPoz3xRScTNO1INjXyo
fcfR/AMJ9IaphyzvIdJKcEi/p8WmrrvMi6xGYLUdjyx+UH6OLlt3OnE1v5zDOlL0
37Y1/vbFWAniEzU8SUEKQ0cRqtHOhECIUiz3LgluOUiEQ1t/DOFT5z7JwFmsaQ3Z
CofbWNk5I+ptIqpF/3t+YZfVXMauexck7g1APTWnH6UvEAyMoH4nNtAi65W+tA7q
Ob8QRkaEVxDbXLKcj5VjRSVhLAHMuoVOBAtu8qwzD+nN7CcroifrwjKkCyRIx4//
tS8KbE3opAYgsYkfQ3e8wKY1pjL8aRmDkzNNGhaQ+kt1PUTXlA+y2fEBpCgtJUtp
1pikRKX72ZbOBl3pntmmeQWyrcn14JN0k8weWcZIh7tJ33IZmWsFU0ZNZ55zaotp
uFsF+R3AJF2eSkuB1pY/Q1RCpnTWgzvyunahJYzh7gyMqEPN3zwRGQF2CSvE3EG4
NoL0kYTt4HOuwx+WbjSNDZaTE680/mzbyMcKwOw1wY78zqrFz/28ZQ1FMvzGinSs
AiKwH2/YrBGmqAufnckGWzwpKzd5ca3j7TI/KMp0CSlrd2IJrXQNSwsdcrKlVGjI
6IS476dg+UeA66x2dQRpAmKfgmLFGJOj7e9I/d/WdYs/gQ041dIlw+z03l3cWIIt
1yniXj/41luyRNF9WJjbMT9GXM8KZp0fZNoMy/3+5GeOPFd5NJQktlTKWgCJ/XlK
HNR9yGscwXarIWhSTkjL4MpeNxMM0zsaKcRGCKRAcDIxwvsi3y++VmcQCUi5VjfD
denbHRbQMWtBWFFX9uJp5lgeuMp4JbjQIjU7p21O3nitFZIAp9KQc9+TjWPG0XG+
fwTOgbtwyXcy5ONQrG1HhwotncJ5QnQbHKX7TmzDaqDQjHBvXSBT/A+vhQSllz4e
lR1DnuxW/aFTY3DeHEPtVlyJz2pRT9tOXmhsOSWykJHY16Ys9pOk8v7VnL9PLaij
ssjjmiH59rBwVG/z2E3g3TM5Tzdnw0LNcBzVsD2oZODgUw2MAabaD5QDUkPhZGBU
n/zeDPIgMyMS8ZNK3wCcmGc9uIScTzejZIyecGuuxULwcldelSy77pyMF0REpSja
E7JNLr0PfHdqUSPHCNiJFrFGDF3pIDuYnlYXDLFPjw2wSqc98O+u2yOdr3RinyPx
fSrOFri0luu6i38tVB1qm8ftF0pcxcWO+vUYSn1ZzwFRLMH8Gc2bCiMeSdWUkVUm
1DEmb+88rFQdnN+Gv+N3KE9tnfHOOgMbwdHsGt6D4nsREhc6l9RQiaf6aukpWkMy
IeoM1xS5J0LIAxVyaZIvshXGdHOZB6y2lKPHbKtpBcczi9XIe6TTVtmR0auPl5C2
UqRsm9cgLflZVq8qlBNpC5Pr9hfYxVXcVTikrCwACMN5PUrFLkbkjPk4ikMmk9bd
0reIGj9X2Avsatt9Ahm2o0ifyexCqM1NpH7NJehOQdwVIbYfTAMZ3MCwdAvILtLk
GZuYFMSHh13YpPbip68t2S0dLjDGKcvbAcHu7QpPUcWah2Svdn1NhrT3vhPETB+E
ulTSxL3bYTK+rXAHCQfOk+kmVdgye7YsQ9r/VH8qkX6l3iBm1VOWrXg+SQU3olov
5fqEdi5IIda/kXXYmTwX5iTowHeJ4ooUXevg0ExmKpptNDFTheS6dsHYHPhQwPqv
lXo96BXPJz5NRbGCxb3/08b9fEQwUAsy8lFF0HnPUanlicB4D5ZkLCI2ES7f19gW
jTvxd97aTJv3b3U4vUaIE6pKN32x3WUlMPl9V/ioZUJpXtLmIHaLLw3ihoc4sE+m
2of60C8/SfIkgyGYmRrI0NOnHoSP3VHu9BkPWzHIKgZyVTGqbE5GCrxbfor0Vhtm
JZNtHLriouYqse99jEMp6A05rBJtTujEmsmyXF7aNIcQq2HJMgkFBQSZogRVilwI
c3pddemns0D4jVd7ZrkXyqA7Hg3DzQug2hMgdYL8+pmOBWAlFcrph/hu2AZhA7wT
EyMtQWRhxz5U9dMrtWFNLcdqTTU7GGrCMX20QEnNRH3f/ggsYzeX+rDbbhqCLikY
sAfXZnqXq97a8M7TwWb6YYlR0QTMWx+hVWpm4pwZ1b28GLlpkjljluNs6tm9O8CK
alFgaUldXiIfqU+9BT546UFjtU1rxfcXUGPCU2u/bDwfr0duSHSY1X6Z58uMDKrh
3wqKvkuEUNvkTiQhTwkzlOiHWBGyGc44ydmwJsisF9MPTsO0BuBRHagMnB8XoWvI
EYNmSyy1jHhGpvPbVL999COP3yhevZFjaO7v3XdVrbfkTDd1yVNTf7vDC61KvzHx
X381UqHsV+Q59GNnxTc+S+pZ8fN3Cw667KXf8Oflx2f4XRPz2g6wgtIflpDki3JB
qgmMOwmjJfv2r1TaYH2FoVyDlJYmX6MqLDYX12efCU7sO5SgK7Qb8/sZ4Ejk2dDA
ypdAruaDUBT4eB4HkmwZq0UHIe03wkT0LMVbU3LubrYf7wlVOJrnFw7Zq8fN7Ech
kdBaIZqJ2pB+aW4IVdVbxpQZnGKZSKkVudebMzxJ/kg45Bkm77mu+ht+dd5LOsAN
SdLuKK4Pue6zAePCNgqJbD9CskkpmNa/ruk0ciBifKOAptcdYTqyblVS4xp1m3f3
Z2Q1D1ssjk3q5ibd4nCu/eAVG47SC+9/ZcuAxOKYlQFkcUUSytgU9Fyk8qs36e/4
IM+shFFvH72JcPrrmqbc1A5bUY+Y+seWm6NcKT8wlgU6dSRcSLgp9SJleDxfrHze
avDm4IgeJ3SwDz/rXOW+UScDi2GdHnuTVyBQKeUtLgWELhL/hy+B60v6eFStLETa
kQvjKUvlcviD0JRjQhWk/TQSLecc3e9H30tn+XR6Z4AYrM8XXLuWxwROFhLYgA7i
+0nGleKmMLgk6fF5Q84z81TxjMoBVYj04OFbtYaNA0hQNTHb7WZ/G1R1jjfkMBld
IpnC8woQZg5+Kbmli+IuTvESfakYRsQv/f0N6m+yWnXhleHtzg4WA7bShnRyl+z+
7CDaneZhgeXPjaHbBe/LN30XHjIh4J52jzfZ3veFki2ABZk6u38schU2/W5krmjj
yVoRL0Ig6JpOoft8Shp/6uqlcpZTOC5Q4fTW1V2OXoQKvAWtTTe7Hgp21+vwaNlx
QCCcK5mY7xBh7CpzdQOeCgft4Zgglk1tLlhYFGS4FgS2ZDKXnsIzQbpzsgHLdG61
1Q4yfyh1tzMa51V5cSS7NoqmdPMv5fiGmRCQa+RGCZSVfvLSMNUPddsprY1aMbLh
p3xsQJBqURZHzhoYo1mzowgiTNVRwpcezyzjM74xMYfeVlsVJGr0obvddDbixkZJ
7UspvjIzgr3KVp+ma5Ys33IQRiAA3L0gGTPbzQTWoAkahw0ipttK2hlC9HQ6jJef
3hdLx5LDNsMCeEFjUZKZytMC1P5UtdE6FyXVd1dcOLImPHP06Hb60z7RzIKYa+9J
DVTHKBIQ1kuUdlabQBpa9M+r4cR2dv0Dw8rnS44jHmcX/wTWEncvF+PEVImam4/U
NmCaw3wAjzmJ0BvqYRhgoh8iBmFuzY3LRdiUpNsx1slhrnH9DxQjgEvY5Cbz93E3
/QHKs7b2h9t/qRfllJmzBn9xl7d8yNKGPUWx8kpszJNHQJSk23nkQ2nK/pUdc/RS
/3g9rDAOl5eJbWLCH/mfiSX99EoWuM44x8LzOc4606r4Zb9nGPkiky/8qP22FCkN
13bKzJMpVnt4i7JHLGfk9kiKoHA+9VlBBa1vpvkEqTO1Kc/48qL6Cy96XrfOKqgP
ZNubCB4OBszx1KYr4n9+dfLAkPaD6iqGuLbhMtxnRkGp4UAfRdXs7vjCp88m/SfF
M4lnd5j1o8mBOGASf1awM06PIXyYCbXpf11k7A+mO1t0LgG0SQ+qWYRatmBaJ/RP
ZzCbnpF1AyhjdqB4a6clOUhgm2cqZCHYoNK25Xl1ploHxvo2F8h5CRuBhpHl/Mh7
LbgDUred6wFci2UBVLsbP0hBQgQiU7SL3eig3DAGkyWeBl9+4S6yEbTOPYNR74qA
5e3EEdeMhWnLkMJutAu+LVygZSbrx4lANDddSej8/qpykf2+wL3Lf8X5p7R7HyVO
vlMamtZ04XJK/aoQTXSo6F/c7ThrgLBIdRh5T3r6m5en0TSUi4GlifzlG6oTDpVc
Z+oHopvJN953E4hlljO28KMdf5+HCMb0ITqWO3CZ31GIKnzoE8js8vjYnSDZWbQn
vZhflxBCoXTm7gEVx8kGkaHPtZQUX47xLqNbXbU/7eiQYerGOUKDqLge7+pCXGap
cpM9pow3U4no/kOGatlhrOx9TrLDYZDoYEuM+3Kr//No3BSmlSkjmyLeIEfJnCYV
61j37GGHJ5nBrV9vVbp6yBaRWIwiD836nvOJq1WCn8sZCuL6zcn5g6tPgtuidbRp
pc4D1rs8T8OXhs2rN5+ezIyjssilM591XYKRENfiRax0Ugl1bEVD/iNksO3TXtYY
PjxJ9bUhrF7bWW4N4O15B4odR1/58tr+UFAoUfoXIlJTn2k9lVOPgrZYaMzw2Mmj
b9YjIHIAQhLnmx/UlQ/mXz2BWLZFVTastBkoRN6T7bXiCsVqSzQyIL9lPeK50h8B
kVZ66+3tih3HIowLQLwHopxbJUes/iOTzf9j09wwSHPigx9JTW6pCDLLehVItWKV
UJJynSgpYpWcTli62jNhhGIdfMOjBI9jUSrQTPefxxRvmh3Q4/4dO+SwTTJcNQwz
JOEycXUZsjhJJ+xIYrH4ffqH40ndB82TfnhRaCLTfSUsc5v7Or09qQXh6/WdfQHH
F9cxLGXBRqHhJNPlKvIXnUokeTn11w0fRjTxoYAaO9FoiIOsHDuDxtprY5RpCO4w
vazyTWc8W971p9HwDhIhiyq1oEqPy95fSgDUgCN/yArRmMn7CVVHLY4dqdRfpLYG
CAe9BnRt8kfTZtVXYkWSgJA65txORBrLaqG0mn7EJ3H8AHI3AIHOEsjrIRLNHBwh
yMddKuWbayIMcxBkL4H3gN31SZGi2Ndt4T8fOpdXe1KOAvp4ksLfpJUZ4aiyJsuT
taZM3i3SApcCrHZv2xALiu6yzcRdbDfOXVD2kaAODbj4cSMYWQ/IJJy48no+j8Vi
DJkTRqX2uZuuP9ihC93mK2jd0GwzeC8P5E4w7evS9UHeql+JL3bYRaFdkkIF1EZR
uc5UMcOp0GLFSkxD8tf4rVYZcEahJOS3R5BnZ5M0NLx60P1cSfasibh5BCtRoQOd
/PbRDKAQpE6MBUhjvjpp00afObsqJZhFnv9gKh/0ty3PHSwV3qXWcxVzs5ZbT3tO
ZhfDCsUVjvvEwm0r2PK5yqNMm+XVokLOUaPphn90CNoMsm3+Znlg+5oOvXhMYtLu
DIkz6As0/4y19GEZ4TRnmFe3l6flsC4s1bmGrRn2WDBMm08RbrP1uiCQYw8sw0au
CnFwtvyFOW0mXwhUcSvM7YcLmHV43TI+YaJTdOZIEoQ9hh5Y4Q9fjslYz6ibqnkp
4hwlsWayUHPGpRK+5r5EIOc1HHjaBRsm1vTZCPeiWfi7SFdM2GyGZu3nLDfkGqfD
bSbb6geVaRFQA3zL65VT6GLQZr2JuItf0vRBhMvDvT0yb8ZNoPEgoO9cFm9tRLbz
VHb1P2r4Ea2wgOxIAIvv2MFQ53Ccmm3DX+qeLTydgto8ZrRnuxtUPTWhjCsDQue1
zXTGjJYnC1+giLOhID2Nml+zP6//3wESP0jrJ0yD5257TErs4Dh7P0o0mZ/HclMe
4v6tkeH/BMiKd4dsbGyUputktrBNaqD3ZYSjc52MbCrXoytEcb6avOSp+vxJwdCn
dYcOuRC8EXrvHbDGTRTpNaeM4y7K0epaRiPUZylTgq1KZdl04omWzzJYBgiLQw8Y
2YQL/SqqKKPR+tEPwl0tA+/FN5jOPM2ZrZ1efO2zg/4Tkekc2O/FpXIBW4TPHa8Q
u0Bc1v53rNMOGrY04TqHRPuI/qCVFDE4cvsLSzOFnKzlcuxe02WvexRGQOpu3w/p
ytWhnL544vtojun7nPGbpKgmAuEoU4A88J7bkzvFM4amOsmQtABL7h+heP2+E08P
P/QtulyUc1yBb7vgalPfgJkbjqljkya3ppXkeyqxx49jk5zR2C1eaHa0njlqRcz5
qgfmACjlUoLBIRA1MKZrXkRAANj0I/0zCHHMmzZUi2uCWW4gFAGUFoHkIK1pbswd
iwNXqKpJWJxJsy3cY31P3WGG1MPgY/dQdPl8tnJy0Q16RTHUIsW9EApC0KyysNOe
B+OOrR7YobtRuTn0QGrGwZB+NqmNn1SIvvM9sdGrA6qH5YVes86oQYNjSmPeTKwY
NpjX5svMSHtUqj9jE+49IBo13SbItZjT8BkuoxeH7wIOnlCYRffYYCXRBK7wOeRS
6kZhR8uCtThxFFrSi+t6wbPhbSxFg57HAo4DZWiuglUqpbyiqA2j5r2+tdFoP9ws
u9RZEhEm9HORjdWutAeireX0UAcxuQ5+9rdKlMpb713A5vAsbfj8IPujEipBWh+K
71E7rIO4fBcJl0r4/9ClJu26E9moCSumdpjMWW2ZYSMQT2v8ZTXFP05uJC6ccVso
dVhSrL7sVuxNPwaNTcuHg9vo4oa+xCu1mjQRrIhj+m6cLErNOGQsmIxbCoA2on0R
HjMAX2Pz/oMhoioqYIqAu4f4jdUk+cYdDeThKXREd80T1rYF/wY4i9kGig+hcj+w
+xI7AjgiH5bkQuSMz2b/tE/Ee+6WjUW9LzpuG423XKYIl3G3hWSokyLi1puXLGAs
pT3uaNmhn7sRPJaQJe9qTJgolA4lmsP8buJEi2lHk6N1qfTz/yUhPlFToHese1nn
JqbYU0CE2TtG+ChqkwqApxN8vb/PDylBiahs3lisLIXCq8JKNcd7XkyenHVtkKo1
UmBcEi+ZwqA7SLt8wC21SYiuZ3bPXm5h3pWMmTDWnQJuwAYzkIaSiuQEjo9XOehd
206sZ8kWX4MgvJ8wJF/Ge2RnSgW3l6aqiCWg+Jvgcp50vvRwadgzW8NXps2wdkKV
dnrtmjCwyBM//7q00Oa46dwSUJqeLw1GA5KgxaPN52RnkWGEY6YG1Fd6cZRJzf+l
KcS1MtZeZfyEImMkm3lGPuLfUq7wSo90ca2aiILjnr9g5zIEuHmW47R8MRqjezWb
EjTtmclJxO5qnbhuFJ9AJ7Q3uJu7xhzoQ7ZC1RbaKMRs7oigw5/nNHUgxh5hD1Mj
ZE0t1EAGFguBSc/44QuHOeKagSoqRijENm6xGXTwTm5Q2mYd1J6e5myNf/9p2jSi
Z3TE2O6s3uAda9tFyDuxn4YKWoP5Y5du0H/O66H2WUaSe19fWNNeGT1ruNdVVYqw
cY1A0t/8OClZrEkahRONlyvDOVx1tBUEy7VesZ4kyuMq4jmNnK9teFCLZ+RGY56v
wRKCn/5j2BWHIeRDXIc17+RmcOuCWbaJLN/WrzI87dNYE/+dt39mrBjhYBaeCXj4
HqVBT6+caweel/0XNG/fWhYy/RGwcCfdbFG7tJjZxE2EfIjOOWqWc/jgdpeQC/8j
3MmlklRpPyGQmZ7GqH+eIT2wRYQFdelOmWneaxR0hmHzCpET2OjjHzYR5ApxCKfK
XIUsYgi15FYGSGW15OCqFYTiiMEXHh8XrmVsThyTt6Ua6KmcThzoHNqU7kPlC+cn
WpPHYLHHveMHftFvCgH1UThm+Oxehi+w1P8dCZ1dkiWf0OIwoRFCLjGiam5fqA4X
k4Z1DdAWy6wRODYR2b5/ctf29YjNWp6CuIbmjfsWxW0jMdrbFf1aL2ovi+ReNYzO
r34xjskQH+4tGYXq0G5kgf3pHZiWDe+IVEzEdl4nrnPiPuayKLXYgHI2FkVVytPH
IgIn1iKTOzoR/+aTFy58BNdx5Syug/vsppS6ghwr/DrYqjjQi2kcOQBKrF+I9LYO
KlmezAAU6RD2/NlxJpi7JHUIZUHx1E7TWY0Y0HYyejSxPZmNRTgFuQtOcrghEFUs
26vl2+r5ThUysTR0/bheUYfvI+I+ojfO3XpEctR3fI/SWWbI04AXb8MCMANf1FUd
qxuSmvaRkqUHh5jWyZZz9e4h+70x156x4KOjYlAGVQnbuIlXKtjSw+IDtzMXZAYF
qe0HNGKsz/HqMgXL4QlC79+02hPOXZwrYU5Q4IRjpHytXIfP3pE+2CVc3/br8BlX
KHKW6h2Ta1Zb6BZ2J5gfRl+tOpSs4TGM2axdCmhDO8T1swZX00R7BNGnwWGpNSxS
Vvu72achBy838C1WPcZ9cMVoWPA+otjqdGeTZ0wrM5Y0au7kFJidiuWjMHUsZLR1
myxrzsCu2adnAVn5ELacfoIGck+OwRcJXMhoslQ1U06Vc9MvJqA++Pf+0ss/+TI8
mWQtMBn+2wVauT/KpIXtftJbaURTuNpjAX3PXA6na2qyMdJQCLb5J+Xgn/MZFZqD
Mw63I0/Xp9TGTPW21KHCcD03FF0yIU5Eewa3T/zLLIxGvlve8S0kUqcFx8//EKjb
cT9BmoyxSoCBcGDW3miF2OuddOE+I5cjME6YxLsge4YSQ0b9ivqsHLxKfuFzGwnO
4noYW+jm4W7FPl3A9ljMiiVmZlrcB5zs2kTxP2bWB6SkDd5gJM7AX3eJp6Eis+nA
OhU5v4SH8UttHCnJ7zT1nwKWwLc0zJdJgm/+IVolc4MvSXapgi68/sOGzjhb+tCq
xUAiV4qylrLz8POjIzfU/aDiP84p/8KCAE3UpHcPEmxeNNNySb6rwgXDYAe9Iu9r
5feJ4T3jVn2SRCnSfvak4pMBruwp5SVrrl0eKQiL4Wn82XXClkz5wDyt+7GuUNJg
k5KqqnWBpG1zg/pfock5MrI1TWDn4X77Bc3x7kvF8HPoQR1LMvzFVFtE7kOKSB/r
nfo3XPiAEW8q53Gd8feTuJJXQw5XAzdhLEV7Ourhh98MeXqqIxWdJnvWg5Xu6qtl
CSeIDJ4lKx768z0y7QNj2Vd10T99XRSR9rICQSPpOlg7iqrdiSARxhtD0OJrT6k4
CrE/11Kky1XaX/d1riNjzuBhgaxLLbcKrLePxXUbGizKfQHNv3FyjTqdkYeeS8IL
z5rseFJUANB7SMsSzuYiz1YpRjhdlSt/2QaE5EdqwFQDBljb2TFGXFFF3lsRkOno
P2VRbPLF3x6ULWzXFd42blPw85LH5eS7LE8zsCxD4qlS55Z0Rv5XenIda+TNZYJa
biTrAdjrRKR3VLJi1KL1Pr5Bj9fUCf1+Q6Mqc8ArSIop7jwjNZR34o0EkI5aasOB
Fc8UhNvgwjh3Lf8DRkIzzgYd7pRIzlK/Aw52XWkt1FIS4agWwVEJhTaXH2PWk7Ai
LGnCBybAvZd2Sp+p2MZvbaOVZFbfl5iwis1mx9T2kqjQHb+ZNsoptedTs3r4BMvN
L9zhkI0SVhVwq+qSXmxDu/IGJpR0covxNS83UQZZkCfPDrSZlf1TcDN+AONwOoGp
yTcYz40Dc80xCyz7fLXJwTquo4lZseaABmdmuPldw2FTK5DMhh5NLreM+lzbTzxr
Ns7Buk72DuJx7+t/MUv0LNYSuomJPikuVhUEWDKlX2YbB9PFk2GQCHHGZDKjBdcn
DzdZamZeAUDcmQ+tKGRp5C8Mb/olzAckHe99pTMLoRXPyPaN+NrAwVJ1PK60q41T
bj/hSG4nOXuABwhTwP2oMpWRnBbVybOHVgpI8HVFGwARTP/ndhLZbiO/FQgQVOIP
7W8Y4Q7ivbBJIt8VMyRwEddIcsuaOpIk1F29uD2gJNV/YttYzWfd0CIhIi2SyIfV
pvubtSKRMEN/x636JkDtP/h9obeC81+TkKchVp1c9TH2/YE9mYNMtaOg9RekES7/
aDQjoPlZdvIZgpMqnnb2jUyV8J80IrflpGBbe7e2pXpSo08XQVMvbfTKH8swhKhw
7mxczdzG+o7Bi3c5OBi9ze0yI8Rh8beoPyaLzvM7va619JrlTzdZ3J8kFgDRB8/+
jhlBJ/IMhLqrlxJqzuvxyskDM9UfOkEqFBANSWZL/EdQxh0C4C2lUZb0zSNfV8z4
WKHDzKqmtD4BZFIbOZssyawP2aGh5i7SKr6cdek1Wzpb4CtXrynQUQ/s61UYIR4a
nBycZJ9b5ky5fZ8FAGuOhjOYHxqE3raGzjbCrz+rMigJ1S1+dCbxX4VXltTu8GLC
qxobkwZM91nTkvhs85C4yX7bn2jBaI0qmF8LLVatOGP0zKOlSqAp+VDSYz2/S7py
sQQbibdQvRIzRaAanKdCL6obPdKlrXGdAaSWKJKv2O6ATeEwXyill/rPEoNxG58P
MCNEnN4kpqDFiKQs6261oe83JtBua5wOVwyFKIn1cPnp3HS+glKb28d0kQJ7hOnD
zrEQHDGViZZr4ZQ22lttZjfahQ45a1TmqQelhCYM8f0xB5alOfWGvJrlpbvmw4Se
A0cxIqsk4NAvTCPxo93PNMOzCk5AriRPkV0cUMwe914JPcEkUNLfg+YKxN5xozju
77H4O00Q7E4dgFPMmDCzlYgm9gYtYz2y3sx6G9xlHArp24+5NGS24hwoAjjuVnKF
3IZFCYhPfuZ8njH0qtS9sV65vOg+DRTKZXfmy9LDX6Az1i8AIEIJ55sZaXb1BcIZ
/iJ8uAr/YuFnOuex6lMcIWTsTMzELbGXqdehFHdpt1lyLGwxZzlwVT5K1l0vE0Kz
yY1LbmzpSrS/tReMRyYW7+asUUg9fGsD7xD0U+6A1p5U/IVky2yY2W6Ya378DjA+
AHpBFPILb5+qUDbd0lOnwZpI4gc4IearNes3G2pCx7c8+It1vYfq8yGTcuUEVcJ9
9yPB1z/eXjLtjJfHYEseUMKBhLpgbuDLdRXKPHZCJ+I0hoDzM3FKzSMtDzgiz0Rz
D92tSutvdPjX6/DmwUKBp00nTGLxYaDUnr9WKTOYSZlsR/t/JqLjbKEFaWH7cY/q
3Daq0Opk5S7z9cjMuvmv14b4EyVgk8/XHy2HF+CIr06BQaNBcGtK1C6w/ULCgCWS
AEo4Q2qrhTuiYNAqAJEgvu1/AyJftDlwptuIBK+Gn1lE1nUKzbA5FXljquR6lpoh
QmJS/1fTTIAolyPyX8YGdT54GNZ9Z/LhmNbGHQ4gLaCcKGt2dliftr9Mh3DNxBie
7LHzUmQEKv47BC1vY5TT7eqLVkZ/XAbeoirp/bYaH0/e9b0++Xv9IyA5c7nimaim
4NWZaFR3Z+0TqlT7IBMHZgthGpiRwRFNm9RHKQb76ywQWBjDfx2OYzvjdTFHD30Q
5X241NLoGx62byfjks+GtWpofn3Oom/8TWw5Xzok8XdvE1JeE+k8uDwdgZN+VN9O
049Gm4iXM04x3gX8gkKtjIjxOWT/Vw0MeqDC0/0UXhkpT8TXoDWqC0pZuvl7L5Js
yPPxK5sq0DEFyU+GjP6vk1d6v5B1LG/pE/z3Xqd1iNsuoyNknUgRb0DiIGuY+SFF
9z170Ko55F+CMqsJWG48AoGZKssGu72rNfyCoZMl49VQmyBzkblaEo22fkPhRwoO
ojq6a2DUNIscrLFGcMoRleolmUycaWYnz7hYvpfI8AzdhCh7kB4GdQNr8XLM84wS
z+4VeMkTj3TQCr2W4BNFg6RZVWk1iQXSTyg1lomcPA82lI7XovbrUMLARRAWMdrr
wfVbQ4ttRzIaAvPy6iG1ZZg71o1wvwzDdjRkCWcQUjkyhkrXc0W+eFvotnLQlYkU
pm9bLyPvzn8qmFuGsiAdAnNfQBb+jtrjhc7cLHpiQmu/WEAnH1MW3RJhtwDLozx6
zoDV88i+WancB5ufxErtROFA8n8RkUilKk9diTxWEX8ZT/Fua9pRlHzToVtI4OX0
bcgfTW2TG5gAu0zGeCiPvNUG+Rl9o7T6JKEdXksCtca6SyqelzM2sHMY4IKSKHGd
PyUTBTScBLDpTTWJMLMC3k+hOaWZtufetZbF3QUIgyFfOm9C3ZkmRolJ4q7fV5rC
qzVgqSQbT7/pN27afzCFbbmCASLjXSnJXW+NUxlljiCZnawDULFrmJDiHabfqNvt
H7zCTvNnXO38UkKjPhXK8KmQkXW3j3pufj5uEWG+ctdM79S32xRdq0mNtFD8bitu
ZrkOkE43PjX7sfW7lW5O+E6Grvqizjc+nWDzmJp2ZR9IZhBhkx0Z+LVZ1g784il2
++GI2D+YlshLqAQXCCZjo1ZORA9L1+Gtuy2KSHA+2kMs46Gqjpzdw54n4GxGbsKr
3YvPHvvNwQUKGWHmd4OMAE5aDfFHr63wL1fEveKRfNHEcozDjBeceslUO8SWQCS4
SfVy4ZKoZplWfnHBAydf9hF5sfNehZsobr/qovAVVUXFmJb3UB+USiBzz3ItOkCw
qsRLqicFdBaXhtBcqFBfLupiZuq2U6gN+ilLIBJ5b0Hoovm6nkDsxvDtof96EDCg
N5OFxbp+n5QCVrQ1EmdFb6EffMbQzNS05dLWXbPdQ6AIoux9NS7bKJZV0Yx4+TfE
Q31FsWyp/j/aNNLsjw6p5PvGD00RWRtqTAqXT/L3Fv3IWhLC2fKMET+WpdsC1C96
tnJd+aWk43dzIv4gfdukXA9KkFnpc8Il9zaZWtyAHwep9xXj99/8z+fH4NUvJ84Y
Ab4slJa14cMDXJCfYp5FVfMxtCJ6Jj/y6RQ+OiL0x9FJtgt/2Xgh/JcLwv1C40Pb
zH7VlNWsFNOrW06U7LCDvK0JOb9T0/v8ULqxLfmn6szj2XO6SaUdwMZmclrvGkEc
JQGk1l9vqMoY4gwYETYtCJaRaNYz8uOfjl81E77tr7QJ4SLxoFHXsDHFnkySE39i
igaBqamzrX4cwymaSbhuJ2glaBFU9PZFQgW29R+C0oFr7azYEN3YLN65rkwJX4Be
Cskjb3t5eyE/OfLoNDmrwEv+naoJhASMSDsz2a6X7HhjLqO//ZPrwjh7RJiieP+4
VxzDQs3Iy5zmSvj3vdZBI0gyNElijpKj+jjKFEXI/jJGIMmDe4bO5RoV3t4TC4Ei
h0Or8b0+qn/ggabzQ87G7Ihy59AZwPwFzBcAQoM3NNzKaBF2ZP4nbeGsgr6yutlx
Ry59XPFWnrAXDKkzsm2p8i04I9v9HFNTeC6LufWs4rOV6z7k4KWcwMtZkdXFQkLk
e6KMM6m8ZpQmm4NnFxNpwM003PBXEjbMl2q/vSK1A7SHkKLvIS71OrkLUaKD1VII
ug0feVV5kx6NzOukRXfRxw/lkqclg/FfbD8OIQ4pj8Gv9XRZDOlNEVLe9Zod4IuI
CHm5YNFKFO5bkqxqcQYyuB/IG5ISBHg77LRwwyVsxi5zHBaqI7jD/UEVAEJewFcW
8WhioyT7B/bsskqjKG8F7FLEpZ+mf/HAN54l7l/EfDUL1pldH142EEGuJk19qftc
qMhRmVRXcmgF55uYhtSiC60DKdV69mAmb6uM78fAhoCYePcr32PMvxik4Pk9OE5x
Vto5HWophUfXvXCycwQJ51vX3N2AIdEpvueAig9mUHc1gq53vmE4bR0Ex0Jb8qmH
uTJ0wiCb4Cpr7ROyMRrSxjI7mylNLD+hVovVP+PQWI/73zjlW68EY4GTFNOvymw2
YBSsWCGxhLktllLcvgQfy50Jm1cZywVIItrNXpEym8gKRq1zdlu9lqzVuII7fnZs
Ujjy6WPcb18Pxh2dcMp8+Jpo99WRThPsxsLafVzlszQjg4Fxv23jxFKkjngnippk
OOEm7WUFAVWGwJvgiKz4Zql3wjpo/NO7+0S+Ui5mZeCXc23aPdikWEH59zZXbzki
oi/J2IvwvYbQbw7fDVMoDWMP9MhbNWfHj+x/bV8OLlfmdCJwJPNjtvghZHHBx/z1
vZD4UwXykzuzMx97o6idg9KcD47t4Eu2Sz8BLAzZRIqE6qwSDwRCim+BcIV9MZvq
f+Ju+uR759WoESuW5VLTFyxupces9Ii9sVaZcMpnT8QarVDyj5NwGMs502MTvEFg
lJBhOR9ZuzcTusXaGYth9Zj0rV7EDxUGLDONUFAxD4iRbHebR2etDGLsscQxTodB
iV2BBEqN+k+sNnN+gZR6JxwLei4lV8AaVw3iMCjJOGWMn8G9xIhPJsbP7acqTqau
a9VnplhXofunZ1W5yuCvSmB07SPWVPQIr9zUdoVXlf0PNx7Rt1aITogAK6wA0lwp
7Fx+k2sEAZK+AIAnerraY5Rc/Y/MvHQJr3H+FlGXYuKHNAtC2i1ATCu8O72JFUsP
BmUXFcoWAD0pKL9C7t1jV41/vauUMxmJ6Mc+D4tTwAHpoXkBUCrtMPY3NUUMKmDg
o5O/SNfvbpC/9I6S7mENYNmS80h6rLA+U+V9JZQCBLbTfvb1uPZWxWgOG6coR8s4
vjYevmEvfKdi8fxSOikWaV+Wj7RalSrKusvKdAZ53onNb1hT/ZEViQK2tyvp9Mmj
yzC1J15ZLa2cRhXYctUia7R3Ixkn6ediYwlFK4h/Oac3qBufgDiiUs2MtSqfmX/F
nYBmoQpuzxH5QwseVuFu7r8cMYoUHcc86XUrupXaFKOsAVbJbOJq/FUEp4Tp85IG
gHWzmnFlV6YnqO9FqdEkVabkjk/KFaA/1Og7P5Xs2+Ymc4XjgAJaX9pZMc1BusQ7
BxowR2iV33a3QHnDI2GEEDQ2cNHjeuweJf3Invh4IdgZerDLRBghADF0fcmmGhaO
9LcfiR6E3RdQZIszvThtvgqfm51chK+PSKnQlaB38jGMSwFmCYJyZnrw9goskHd8
WfjX0tGcT/f0wp3q2bbFBDHdMYH03GaWv8Vqoxu+KYyJ3E7ynhI65hu0G4/o4Hw9
7km+5dOvzLYdAkM/f/Ph2VlWvih9qLNe7bvRIat6j1hYhzlMrGP7CFNX5pwlze5z
uCp+2fDyY0aSasD+aGD+GW6aheiA/cqDAmC4goZrAG0jCQpZSuQrnqMG3MoXTRe0
JcdYwwap0pHVR5ecsd0OAQJOqjOB55AgLVJdAUxGiK4MCV0RqZLufLFOAh2zjJW7
10dP95NGIS9GY8p3GxiaBXDJihLXMZxhjCIMC5/y68ovA69XE0aCVatlwkqPBJHo
ppo1ULRj1FIuPoWVoxrxmeh/S55YRjFAuGZboL+Fmjj8KQ6okuGPRMc2vBz+fW6Z
QjCCw6AtzrnzeZRRYuH4lotJFY1zo2WZbs7NiAVo7y3ybVNr10Ebzg7PVrineza0
eJgZpUUSH/R6oQjFEl3n3JZg4Z+JOvd7GoSB/rAtKM8Z4Djosev9m54+UqbeqEGO
fOe2n5/I5oOGh7QJFegsPtPy5ueLzYAB4y1PzSsyfnsJK1gEbcpI7kA6kPwnrmW1
KxLBt+GGLY+aPRiIFLcD5KzPWkXoOGYZdW0ve/JMjIUfISRJ3pzfUJTnG/LcO8DT
jb0BZViWEBGBKMTc0nrmiooCMh6ERyBFIrkElcliQJ2IOq0dlhUUJAbD4z4hpSSq
CRYGISrL0fdCx25I/ehV8NSn+ZqoTINZRESTYEFTUzQkCx+jPbWKmeSbbjwqfpeL
QOVSBI0SM1GW2mQR02edZQZGEXThw5XDEcnZvyOyBQEf9465N8CSWPrwkriBQ4eZ
Svxv50owqDB+HEvA1pms9JR+Ra10k9YZoIN3wPQg/I3j7QYZM4nap7EmzTrSKsj9
qftU6ZQO8vQwS+c3TwpUKIMuxSOk3r2DptyEyg14dyZhCiTwUMuxvxQWaguiGUjr
2HsSeceP8+EyypsOt8lUYvf0FTqyVMTPAkUmf3/uMsEAzuTSG5r4vksnetiUF9ri
UEefm30fWP41DKK2rSaUfKHyPGJKku800L5NL3LgFizwHEqhWZ2WKM1r7M9IJegI
pUVCTyjr7oQ7cweb1kdSmmkU5QD3/YaW7rbN4y5/rh3KX3KizGqMyWMY0Z6QyG4D
ag2wJoF3NVyg46NCYI2wZdZ2daLX38GuF3aQLh8cT1sJkHmmv/fJLq3LpIYVDEI3
qfMMI7Lh5pOa7IMNQ8mxiKThJduzpOOCOJlZMxEr17CRAEsAkGeP/P1jNktP+NTI
sNxxgs1AF1MRsJocKfaz44v4JAr3P/iobOY+CjgMbgKuhbgVuUiqhYxbIHbc8jPr
Uw7hf4G0Ye6tlzzweGraNJuT1kzARqZ6UQYzC2QVH/j7cGDGYR6puAue+9zSK/ve
pv9xU5klGG/zvukt/7ErWpzBBeHCMHlCN1hC+JKcwEh/8CgGvWCPUnCmWTHRdnjq
fPKXxyKekVvxF/s8Y9f40aGba5usj/Sg2+ZSNWHwRtBERI44+zBi1iwijpvOkaBS
OW6cvZf+0Si5JKEoZ7HuWzXrXRkCJXKIlCnyesynq0CEdbl87BdcrWn+6CcQItlQ
7tH+APrUyLKvJae5NHrMw16vRNHAhK9n8pr0kal8E+gl0ObYEUwP8bHPeL6sZ7Wm
9zMzsCDnvpqAh2HqVufp/xHOQdd2adWmc66J7ShYRLY3THHnrElQhbITH0fPcTkg
rq9k+Fml/EuTr9UDlwYiJKOUc4NhudDRTpnw/k+4VB6pcXT8oa4iNMBDCwTozIYM
XC7/SykNlsuQ7NeVLwtFQr3k6mmNHHWqcc5wZtosHhIAV2lpJOigsit/EKtsEDAm
uB/9CyFEmDH0ZGTO8ShCDG8PU3Uizjl8fbvjC+L/Ru3hqGTQ0JGZ9nGAhrfFPGHW
s+MsQgmatwVHaYp71MKpghrjyCwayiyIgZGdu+3BsDvtyGa0KyO7T99ZfAsgzsYw
lgpOheSt29yFvjWOSJWxjoZsYL+EhtR1nMwP3beg6w+mYYUBkVpDhFTVceHwvzsc
MXbwyLvP0ONC3nh1CJz8cQYfT6u+9o/SF3MRh1SkKBBbr+yyYFVvs9GoFy7AT9M2
Ea3/aX3i+xwQf7acuY/fsx+F1aNA+8lbmjRTZpKvogfZ3FK3+Fkaf9Ti1LXfWoKN
ZmFXFdiJ+Z+IcI/G4TZNjea6gK8drqQ/C4UnaW8lFNTtu8qfiwUoPmFnUqa38Nl5
Kc9n2eymR09PToQsHlnecITAb/lHQponshQ0aq4VX41lDOASszYwudIVsw2hvN8s
5EMKM9sDRsAVbnr58//ux/mhR29pYqwtQJSBLVGu9TIJEanStkT/p92/yK+RJsUX
mU2NeiM54LqNhiUV9IirjcXgnjHTQQQgKitdza5C7yDbXgCPAyNn8+5OrX43Qrff
RYSc6byjs5bmvoBo6E0YjaEo3Djr/Z9byYl76NUmDHqTOOt/hRKZHgr9JBol4GNl
zILtui6wG+74xr7DsigRcA7GFdup6tW+GLBhEEnePtOC5egIsQh6pmtCiJhC6JrY
OKIZemO+9Cy1zzLKlFXJYqYbvROnLmuTn9YO17v+5wihJvy5u8Sa5uWrdChXiwo3
DqQBV1ZtP1sNDXGDsJYsJuDj73qf5Tc0u39i8dJl3cGR6USDHX3mmtwBe5fm+ELe
hHMc/lSH782x14DqCjQU3jd+U0U9NLvWD26x9pPgFhBSBRXGEyjyiDQQGsZEhOMw
WAURCFeD80qrdLB1i9oo4KUeMwUJX++1m+bjwoQgDYJIfBPE+nlNHGm9EOvCgEE8
/x5/f4conr9yDg7f6nYJg6Obf85Qt5mBMSzuVmTdlh10bxu2Oxhr7VRilG5zYO12
/gHYLR/m0T2SlmwP1DRJpObk5MXcg8xMUoGrI3W3RgxmDJDPJyFMriJT85QgS5RU
boFThfu8oH6ynN2vaU5RWT7dx+EiW37iMEXC6shrR9pV3TZUaxS0pqmQEDICSH7A
FuGGfKOn1zLAcpCI5zF1qxYjOC48KOmV/vhaBNvhu0MuFUQnIvOVRy89I14kJrG5
3qT9wIRkcECXz26WFu5iaGgsR1YsZ0OO/9k6y7EUiZgjlZDzTTYCKeb+trkyH9qw
ge8bHE/vThnlC1SKpJv81SSUvYjlV5yiyYhMeOkf4zMWuIvDoFZQCzWDRiVgn7e7
DeErf0puYoYeEQfI6g/GLn4oAqn51OlsvVI+fidYi7DoUWvJKGWcG08RSycfplog
bDv2PC7XFWZymBeVQ2gAkKLvOnYt3JpbgWpFVUoMss+7kLVAWhwBjIgw86Nbeapc
+Q4PJV02XI6PFsvf8VaT4uSFmqm4p5PGDv+cuKR8fa7djhEOTTM9B1ElnoGKTq+E
ISJ6qqWPJ9pCH0MUbwNHa4s5BmrVdniUS86abrJMGPoh41jJck/g/EA/Sszl1Rtb
wNgOa3nANMCNdKZx2pwTyGkCHf7AmKbEwDyEUgve4dGgXSsx0t0hQceAzeZaz5YO
nJNYfuiJDx8g4ICC9/5JQ8OYajyfsxnSIiusw7fVWFHDSa7Nc4c29QMeWWfW70dh
oThsbNe5+MrYurqsxyLuw6LD/SLJkSuVCLg86m+Cn3r7SAgNsk+VDD7MANZf4GJk
amRFbNF/kt/8xy9O58FokUYkSBB9ybuSsXATgoiva161NxwnUPjdxMtmxTBKuS+1
X5UCqIoXpR/i/u0BagARNenkbQbN5SepgIODt7bLHwAFdpd647G1MgIBlc486+L6
M/Kr7vEJAi7kvfainIE+AHAS06Vh4EFB1cvMLcct6/bh0QJMFITAtJn+bw3gulrP
fWc3d3sWDV9FnjgaAeKBZcUQKfLf+d59Sym0Yu6cOZbOYInz/bQPAdT6dgTqLKlE
uLC+PG7Fa+fxMiTnNG2oZBl05y0CZJ1s3yvKz6EKDoPHHRf0sGAsczsPG4qtCO1E
ZNHmts9UZkT2VatnUzi6sD7FI1YZeIHD1OgZIu268Shaq4MyVon1t84PBh9SAdXd
01YGk0Isi+OZ/NJf+45bJqCkr4pA+ARfOlOnUBUGsZ8Rpjf5oi5+f5l4zJdAR3X/
W8mZANcBMCeTxcH1x2lmReNxcg2ZsEjVhEiaWIthjrwiC1bDoeUOmA/87Q48iYpc
W0JDS3jlJclpUw50Ks5IVa/jM3v3Cg/dQDMfcJfEzhDnvQO4DmBwp74zq601e8Fa
+Z1n5yuLj9vmKW+OFnGyF2fIlA5CSLgVwW85+oBwjUPxt1Gegi7Kvg+siDbowFCW
8uLhxFGVTp94juVIkWXTtpNTqh1g509WDyTvcMJ/PL7fHGrch1t2yXaKoGsLuMEG
yuZ4ECvG4MEn3dnfKXghFoVoFTN+9yRaURbKyu7QQjkK3aaTIlY1YnOUrQJaYdVR
7+2miq7aNFWG830kPVTKnQGrsDQnkHkQX84G26X4IrdNTWvKV9j73OfZLDJy1Xk7
yMgnALC6muJaR07mJkpABYb8imzSkAjuO3+qfSztkw+DrnrYp8fHvXH5VVUWCQM+
rlRDrnzlxOHfHcRo+pXA3hoTBpdhNfY8Srz+pzWmrlMWEKy+R2rt3iEQETTiz6sL
pV5ZLHR1iqXrYGkGny87aOl96Dbd054x6RzM9037BDFP+N6nsY1xHZ1vRBuokSh1
2WrGCGbSrI0huq/E6zr+zt8q/6oOq7onpEcuzWtSq3HNJ7OF3AcLpOuwN8jZBwFp
BHZqLFBqwzGHvwSVh3hr0SgJaTE/l5Y3vXeceYgZtpUKNM3qGZWQMlCWypsW1cF0
szfrtYkyb1oHEsHXafGU0QsTqhFY1Uuhny5t5XZ5LVucSJZVBdFT9RcOXD/IE4RF
XqSUMA1y4khSyEHIt0Ch5IDO3xt2jnskeJQi1sgyhxz+JQIdad9gU8pOo+6eXcMn
aKPbF+hxi3v+r84+VIKsZ17T2NkDAKc1ZWv6mekKibbM2mctSWeTy4Y9DiygLtVb
/kUQ9rQMlfJP3k2MkaPPb7zvscQMb6PJkXmApEmQBWyOcCrYn6XaVKNnz+qE5VDZ
yTZDTapZqEqqANWOu6a+uvh4XnZA0SVH2BXkJ+YR59vdYeymvP75iKV91lIF2QwA
RJFXnK6TBqllFni12HOz0lv3kEv1Hn49E3HJbOb3lr87McpdlSB/hbh10bM92G4F
4L4NcKgvBHLnIpkMkJp2GFD1IK6vuGxdWpsHv7tTqQNfgUM1XIy3tomyC0H13JBk
qvofo4yWDkjCTuQgsWjZNRya3RXWrB2/Dis3tJRq31FqpsV8NQb0QsZJw75S5SqY
crqXu+LdDXHKZd5qQp/2ISYz859JOoQlnjl7artJDt+1JJU9NnOYB1NIbgL9CGjR
Z8G0KfxOabDSurhiveErGIlS7Okn3KuVcqZbS9E23KmdIKIdK4bISLkz9NQybr3Z
E+eXAz1tVvghgUqccK6tQV0q9LNvu/rMhGS6d8JzCBui3+N19axOJKKCaj+Rzco8
ZKneKfqtl+ZNYXUqCc6HbEQEhz1oM9S9ZNg6WKhZnWoQFiR8O6h2OH971n0CuaAL
ab0RiFkq+4N+varNufUOQ+4jyEf/AEhMVEJ9cUEXQFW/SJ+uLmh+15d3L4x7/8AB
cyFUwbF+1qyqts59VNFasocJvZt0bXXCoxKd1GIpS+o99d09NaOH7b0JmOCU8v1t
ms8/pi53XqGEQKx6GyXL8zSuMYDzBKJSQ4RczIo/OmmHdrSJNjU5rBXnPGuIYEAW
mxqTZdg0QYlwKtCqubMHeuKxJ5eg2azr75FACwr3AdlCEf8ej25BTuO5RuP57ZKw
CgbK10tkFSwxetM2toEqffG9njXPTje8qhfq/cRHcC+CsRVkeCE9U/DYjqURZ//R
iOoYg2Fo6W6G4adsMbEoqWxqfMvn7Zr/TQrZBrc4/xBi4PPgxO+SioYXaLY8dKmI
ZChH7XOkz2u7zxdfnX0Ac+apX++cqNMjkSVfKZP0vIInnfi6E7lEMJ1dBHCBZ8GZ
T8+CrMRURuHlwgQPcGKNpU8lC/LQK9UXaU8ykWMtwPv+s5355V0wTAUgoyaq/Bhu
faNb0jW/8QybHgOdw6kZzpslXwE+4agLT1yaPrRKigJ2jx1KksQ3p6OTJZVd721e
4vDoLhG3hnurTe/H6iZgSTHKOvQ8WcHfzHBwi1HQdcAJLHbvX8u75XS8ECpGkyUu
482YNetPUCMuSlqI7uFfSY9ZfCasKO9ROrduTmnOFYQCLulXPFZq62LrrhnObjXx
IDDzLt46JZ+pdWjcmJoBmwAV48fhnjwErkJqr8E4pulkku1sNmA5/M+RTyxEbiuX
4qWpA+WQ5sV323DVYnKlHJPNpP3RhZ7QZq4jV/SN+TrTPNkEwZX+kwhfvmEflW14
f4e+e5saHxunpKOK6+6PHcjHVAB/dpTlh9+QJ1bZvvCMF6cWQ/HqXc971TVbWbj7
i21pUvqn/JSqWRPVAWnyuBmfcflgv3m9FloRpBizvci965rU+QEcPkvzqCCHtDSy
x55oCMkD4IEbWgHaLhLAPQESp2ZsHYZEQuGCPJGfPodSpcn0AMKho3fPseRrSOc6
bE/QHVwfSzqjsY5eGWPHtKTy1mUrxKTivQs+g0ZyDZgw1/Y8ZT3So5YqNNCHaV3l
MaxFTIbmEfusQ25pZlqF93/gF2u/Fs3ES9tkWj3E8JtL343E4SmznJeinKD5xQQU
dIiPWZvSUbSWdwW5O0nyXccZTXZO1aGSPzMCeLhJvhEUF0seW2EQryKhdhY9u2eI
vaGtFdOFOMNciYzSv1C+avD/LVmsJ6NbbyqVVAVn0pun7QW3pXa4PIk65ixLDqDJ
y1NW3pvXjaHeKE3Kyc1VuRPTeP9DZ01Vfn3xsHjQ2lj1/T7SAJBfjRjVI/Sxnzs/
BddFqGLlHePSLstHKXRx9nQ2o3RMEewniJ7N3lDaobRV9Ha5NiPV35xc4JocErUf
GRv/HZEzNU4tIEoeVh89q7BJhKGPMx52UyjXABnoEgc6sMNCCTxmKNNd9UPzHens
HehaAd4gpr9VTTmMv0mtf0+ASU0izK5AUHTuHnyq1PPu55ahrliRzbrmDTwaHu1A
dKWbsGbceW/PpZUMpULECdr8WTxauoPtHjyBz+5fbCgpGLszqqtZApIUHJvkM2yV
AYW+oMnji5vl6K04aDZ4nzrfj8g+KwZCxHLRIrnSBtvtOlLlnItm+zqgf67v1DTv
lE4bCvVQri+tQjCJzB3m4X+/xCllaRzJEFddbv+f7wapTpWghhUJwuOYBR1xpKqR
gGaumjosdlz2heQWKD4cYUhOgGYmbbcKcFiuUjy1+yJwuYWEEPvt7JvaCkXHV2G9
/neKLGo3jI7pz2zrsIivXuCciJRklfvgvp771EQdIOwIaK+uJ27vwx2/QCtNJBk9
7xqHwwSirHuz5kiZjosW3mOr/MWBP7mJVC2anTAiLto8KPLoWfoiZazbY3yKbusU
MLnsp45BTTj2QFrpGppJ2ClBvWDNf75i9pauleaWfcReNMLhFqfEBvvCsl9yqLM6
hlhz490EAN2ofBQr1rlpAcG0cmJAyzSIfPvRja3iVJ3r4lsoHR/iY2dKJPypNpvF
1jvKALUeuvOGupkuvzncMoJiv/xpKN4luYjt925Ygqb1/eOPTHX12ni9dwvMCwI6
zKj5j88T3yIPdp9XsMnqBCAurgn5uOrJTAQCGsx6Hj0l+93eDrQU74gDGRqsDFfw
eG4LYGRmnlwJ0+GDWCdfj4+cwJ78ws3SFMRt+RP7/NtTkHYwntrt05HowOCQHjya
xtW+u98Jn7rrSgPwSOZlTVoZE/llNCzB95za0SG1+zAwbUJKWVgOEwy4762z0yKi
GQMXrXmbYkcbFozytR2XjNjGWaFmXpsD18slr3KA7Q+RL3k5c2xw80efQj0gYtwi
Lg/njEFJjArK4QDwW39OBbMhTx1+nGN1CYk97J0vX4BgXjGmW22RyHCxxHjSwkda
F2y++p/tIq6mSArUzEPHUust5NJiY0EWiH4cUlk3YPABuKnYr4sS+5vnG2GtjuOM
2lxvrapp7JpfKiVVYJB9VKOTZa+S4IJi5aKhQ/6ht/4V4ymiUnAnFvaWrGmTiqyH
VEg8q5cQ2jX7agjXrwVFfiKzMo5m8Errp93Ob9iD3Vjm04NYyHA0qLjjTRI8M9u6
16W/E0OjUvFxbed4WIHtq4iVC7mlfQY6YhoKR5PIsgYf1A0jylIR4keK3eYaOcc0
8s/fcNFBsHdwYfOaMEJttK3H2lD7reqqWfewhxOF3+pOsdN+45dRzaPy8hWcF01+
g2nLZ09Pp1zq5fospOHyoVjSrJjl7UYFfqpf+nS3JuVxqqsAh2G+pLPRbPq01xar
DU6z2yQ9Kzt2LfXHStwyUpN6Q6DNXY0SweQUmSuv8geLtr8ARHuOFMAz2PKePtvw
mu5VRgUd5Q37vGEdjkCVO8fmN32eI/qOFa20gXpmSICvkQ3py3RMfkAEvOH1Kqkr
Cfv9H5+y36Xq8dhFQ4OAldy7/3mswhT8SHNgYILLLiZ+DQ4WT9+nuBE+bjqWeLeI
YL6BrTvpQvFAe1aHzTpP9xl1CAMi0Y1JQ1EMLiG54ewvZoS8BGYvvjd3a6+W79v5
nVQ1B1tTtMjZtmhVjpBErZ3uU8qL7I5eCdAdDmrdDl9yp+ClhSBvV71hb8qf3pL3
2CN8STUrmo4kKsrLH37Yura2t68NqAjB5DhMxPu2l8E/fzfxz57sL993NFLv3S+I
D38QMPGix8g0sFm6a97ttc3dBRUF1ha0HZMaK+bhGogdEymAikr5FLiG495puLRr
dCE2Qc/Vvc94dLpNe1k3EbxixQMpifJZR8nUa6BGmuBBZyMv7pyHbVrXIQKusKip
stPhOTAidOfoB4GKK4uW58hdLaDFrb0BSaRAWzMOI7KHCZt+iMtWloU35pzGzGPF
Dh1IQWpcIBd6vWBWBDgKcrp5DFs6lRzrQt3XIpxyC3U6CQyRSmy69kH7OD15zsOK
eA7Jp25zUKPBj4zTEEJSsYM2T8vgulQiW6rofO6l83fEvnaFIRlDhffbk+bbx8JX
vOpyNBoFfGf5jIRcYsUIhcaVl1iYq/VLWMHOHidQfLitrhGJwgS/MPDGdGGLZdCG
JeldryBBWre5Z1toPoDuentdNrmeDGqt24TF287mzgGbE7GI37ngxn9SyKUVLbTe
AtfXw3MnDRhzEzYPnJrhmulCwmTCLqtiG1qdeHCS3l1nDG1cRY93KhyW3z109ikh
NEvFCELGrPrJsznuvp6jGzKHyyQ9zJigy92A/KJTnhIgl01eFbuYiYaMZHzNgr/B
SYKnOBsiJAeIfyZeg2yGPZCxkpOIB0sTxlEXvLRsFOO8O6jmGXK3y6dOp1CDn8Aj
zsUPFt9HPhL5AeLboG16fhIhyGHOBiW9HwQT1tmP/3g+jYy3Q3td2zDRXj+yAdJA
xbhxrRlEowmmwGdlGSKTaAFLllIJIp06Ml8tvJttAXKu6b0OvSHJr2Ae8VUq64Tj
YsXvK8ubfYpEsifW+ym1Y9t885GdiiGJi0GYutf3+IDbBn/cHIaMX5vDaUAX1F9r
UTn7eFsqiubJAJT2bg7f2TEEBALhFs1FBbDEggzlhUCqeDB/et/qtqzRqF8mWiHz
dFFm+I+ozD9ysmWKARI68CVnswSg4YHKsH/CPYt8KTM2jS3Q8m0slcdRou6eJFuT
WizVGcIKv3bC1ZZEYUJyQFMazEvVvXZcAvVFHTlemg7BOY1+XP6r9qVrB3kKnWoU
y5nah1BQ2oPxxEbBSQUdZcbHV1rUNuf6Zz4wmIDu+/FZTqcEWirQBFH7J4mlXFWH
Wiqj6ec7s8NSxmv5BTgDlkzl46JKU+pyAYVyZgbZ+onniDbJB0UQlvm68T+TX3vj
WG9shQ/xnj/c+5tLDtxDv5f2tsNnV7JLSC7ubPFYIEZRh+jdo1rMgKnL4z5mbZeW
U7/fbZlm7JJAzMj3VBYl/FOuryH7ry9SOKURfz3QgXvlb5dTlVHswFx0UpVybJ7h
0sJ5yHv+1PAt8L4DHqf93QDy49Ov/s+gEbN7Zjy/T2z8tk0JzGIa1A66VnBsGx2X
XBhkKw3nyqANwD6i0xj8i5bzNdbv1RmZdi8g1tbKXqw+bt+3ecK/+XxFPFGkP2O/
dyGlJzfOdzRqERRiOLDxh54y2CTNSSHhSebNJ8mbCKaajYSXfTt/kxII4ADmihl8
8Vv7omfrkKRZH4UHlcBtf8bUMFsiDTM4K85nsSLfxpkm8YSNRpjnQnbUJezG/0ow
PMEfIXobWcSBHYFymJ9H8gC3khSIVZrspEcPP8wpdJfQmIvZ8XaVQolBIuOPEEii
2LcFby2XEBzoPvLAlbO/KXlNrcHvP2k5Fk0VoM7jOnaLW97zWCxiVtGMgk9Ebm/w
K4+761mSUXYjpWkGbd2MbE7tpvPZjTDB3JARlpCyIKIfM9PQvkrYJM9iYrJL9SFV
/ugHWt9APXxiPw4U4bGkppmeQqAwCIrBmQKOyY/jp+xrkqewJeIxCzaiiEVvGBZ5
GOBj8oNH9PJ0CECzsEu2Cx8tFLMTx8ODNrOlbhC3v4Ya9WInGY4Pk8tFcsieSQKE
6AzvxWY+xY5hbmUpwFK4S07UhRJ+velfuj4O1k2j9VntQ8KIMMsUvxcUfHMcuSjI
Vz+vc+UsSfbilM04456h+Z9fiWvafp/qR8rqTSaDqz1STpHwv5KlFlBlGIw4oOWR
GK5Kwur/XPvdNIoyqpetF3qvg6+VJHKBML1LqEVqSiIEn2hy/VB9KHlJv4L+1ds9
jiPWEAD4rvxDJ4WNbqYb+4OV3dyim+tYjhTHTOMfQI+qbpb/Kx4k0mnYHPV20vEd
VDLmp3I1eApq/g90m7dHt5ZhY9EhToV2LzcI6P0KN93aI3zXMne5hSgahYf+LH2+
h9BPPL+0iMoNPrhjrieQUiDl5SmmWCCqoRxcUoZOO0O3+w9+DjJb+zXxYLTz3Eat
s2BLzFFahj/o4t746JZyEhXCgukxxm1YrWr773x+3CQ+F0sxnwM9By0gh5rOT3SJ
QFCwo/aiuFdoLIy2wdZ/Doq1xeEv1smrSu7GpMhvkLbtG2AR0oTmcm186wwbzT1J
LhNv51YHDh2EPSr2VEZOyT7pG9p5KJ7+L+rawxwMMElSndA9Go7CS7FpFrDu4WGi
8LA3saj344lnX+pmz7MA58DquGHic0Sumb8ODCti1hi7bmFOSYYfpGkS7stzAeEu
1wzJsZWT0sxhlX6lwAguFaWlu8Cq2wvjFYH4gB3sTCD08zbHptY1YOyVKK3dvdM9
/uEYVBBdXgZ1aJWpy7ZhvkstGXtA9TpcRnk0NafuiL64AIBdDLz0/haxgibnOG/U
0e8RDj6XZzFw+KHQOCFXCFNUmmfrKNB50rhvYQq8DKFgdLb5QsfX+MpzqX1JUztW
Xt8zrYiQiNeuC0VTjlCvDFY2moczs4yLjOfR0qi3sqDZ9J/PR6vHsdo6UG6EAOyJ
SSIwIgj2V89ZqUB5NR8/Ar4fdGJHMWLggnVxad7h5RTEaPmnl58z9tdZSX4pvo1z
rMwou7MUtiYuGFWniVTcFY6Fe9AJtNBRemGdvsfPW/amBMt2BoqDn/jFa/PnqHat
1XI9cb3djfvmDEqRx9oML5xxxkHy0elbIdwxROLfHUZ+D7DjoVqhuB4zkdRBrNzU
j4gnb3f0xexZ6SHTKAsx9ILzOWmIqXtsVWBOmepHLerlugaBfLt+P+6OAnh+f85C
/2B727zIuGChS656TnUyxWIFA+BUy76fx0XlTrnZ14irjFdZwrIx306hrxtur5R8
dMEgP7MRwmroTIYh9BK881VZ6BA0FF2Q66v/mBLNw3ZpTgjiinAALu1Dm1rPAnDa
o0kzWraBXD5P4nP9F6hzKWiARcH7nPeUxk1rs5+xS2aPDROfuiMgvgfaGQnBKWsz
uArnFxsJUYemqzzfJG5iNbS8jiPuE0FFfI8sUJn/hcKrxHhRhQvpzJCZHsrmMaRy
k/6BFapU44g4+/14lSDSP+sTLrj803C7WxdrVAeMC8bIe42XxnI4UeL21HiduNIy
WK6WJdVqkIx1K23pU2VtHQ5+hghDiSG60rNzpeGSiBkJuyRkz6rc6UmyPnKoaDik
Og6U2uwHpLcWBYJPxzc2dxMmEJVY6bzbGIYsN9o/bTEtc39NIzXs/m0zmdNOLU6K
YKXCS3PJ7fkGHWHffeWiHpiEc24zdPnMBAPIR1tuRJKIpeeDd1x16lN3ZwIygh1U
AD2j84k3hEDnzQUv+6I8Vn3TusTugxVpv9hiQk9MzpFCTBwjklBs+8CNPi7mnhVe
u+SpvVOF+Lre+ePo2fCbMF3mllxnLgDvR9AXv9O50M/iJTASAHvTeKe2nIjcLALr
qf4Gpg9KUiGMpDAN78sapAEbS990xkSc036gvYBe1emsMMvPs5FvbmgCB5fdDUdJ
tom1WgpDCEGxSAFCVyGTKm4wMBb3EYb/YLJ9LO+lvK7AmGvPDTx8LjBH5m1ClXTY
NDe0u7z3HhnQztys5lfDK8X8LpeV5QINNuodYQAQwhAUbGkBYWg3e7+nmGdp4R8Q
1I4huOaEHrUpekz5ebb00zcxWHUycjH9LISqnb2io1uIe/issZiWDidVWrCCSRPX
j6Cr2XJxi3yPFyv1aOcXGeHtt0jbQXE7QvyyfPTwyrn9+vL9wwTgg8kSQKiOlPI5
3GVJueuJTl07G/TJoXpenD2pnXH162DQqSes0YrTD/xqDQCfdbYfNws1secA8/TF
83U28cQw6h39CNjRF/2Jwqbx1wrWPn85knnkKruqvthzWAn0wsGADEQHKvSMcFuM
BI+OXY9xDo6d1E3jbxell74B44gkcw8dTYLy315BqvQNR6EmZIhmQ5FNQJuZQsMl
kZWVvA6El3MSxAOnoHSEP6xb+yEVzv90TcNbsASx1DvvmLC8T9OMp/C2nKmjjeDy
0Q/AbP58R5TaXr3CRiHdwuzh/xPxH6JJZsbeR3TXQ2fSwuooIc+ElJfUo2Pa5+9B
awq66bgtNOgG4aup+1Gs7yE51mkd+nWeYshAP+9sg7KWniTmHlAmCwzrRTT2PEpO
mrDX+q8NkcCKrgBCWbf6AB0AzQ9CCaS60z4XJlAr1+updeAA9wBnwzGx+1KIHVc2
9fqaq1vauW4KRgiF8aHyez6REDO1D6Ur8ExW9ByUeFGOhoUsgvKTBTYMvP9PyVRd
k5ocAVZrCvhcHK1lFOR2Y76gk4XCOfKAieWfNKTuVKmXrQvknf/XAzoT18Ip7nMi
EC1S8sWWP88vwse+PB5+0KASWlMOdRoL9ajtLdjmfp+dkyClmz7IzoFM2lLNvg0S
4JOyArVfw53s+/9A3fPDWc8tBenxX5axE9gJH8e2fmEKTBl2XaXyvLAIeKWXFdlG
DuPAxpbmQMJ4AwSAY2ze6WoNRt/y3zO/Vd5DSnnHES5B5NMnXcG4ucM3ogFngxXK
ZmOcu6XqMg0x0ASR+E7CEWb7m8b4k4/POSTwyjyuYBAOtJZt+y2/K0XMIawhb0f3
75AVUqem+nHLCwC9XmK1L00et1Ia5js0xMUSxdhOx5xzESEAdsiuYQq7RKyocGor
GSyOWDiKaQBZQEQPPt+rL0sUMim67wC2G+CyV4aaNWwoE71jUiEh+5jcpMyZdkkd
EFjV73IdJOpUkdCA0pKgUnJawQ/FvNk5bRIlMoErWy1OtI2hv4NdVJ+fxg0o2BOO
JTkylBTSjZH4k+rPS3KDfwe/RCPEgznyPIjoIr5IvGWCdDSxDVYlu8U/8HLI5h4Q
z3mQZbAHHdVNnqRCvi4HagF9r9G0sLYpXG8GVBkHPSSFQrW40UR8GDbOtG4QljGj
9YFSP0y8QRm04iGXoDf3TpRGNR+Z1zbGXSXMVkSb7n2NlwXJm5sleeT2W1Ne61VD
cJ7SKbe96TwxseHEPJil8oShqWnN2++9o+34SoagtYtDSLkGnLc3Fv/WUwHmFzcQ
S0fAbqHUIc3OnoaHCTxfL/GnwB/Si9+OW7/f4NP+vLmnPI0+4aPNrZh3k8FgkA12
HuirgWwW7pj4sfYMIo2FfMKvZqUTq0WAeNyFI44aBKu4Rp4c4RphLiJVqDOp3IbK
abVBq9JvwPIPSSw58DoPMGEABYIfQX9N050t+fDW44WOtUW97klXTjcStO0Nl4Mg
7xklrpNMuhIM6tpgstA3WFiOaRJIuSRTxHC3FtsSnLz9Zz0/4RCBuEFmvYjjgEO5
F6XtVO842DL/0D82daEHHDhlBk4va14+v9MbCT0nSBbuzwlzJRWTEBIDGE8QCIoB
r5p99OFzTjaXRfQa6ojCuH75HewHx0ukbb6p8/5rwuHipydyCNTt7y4fHqmrmuKV
+XD93RFA8lgw4mL1tAI6XKpu0fDOVYdAGtYbXR+9n4TuP1xkVm5/QSNBQ/O8KWLp
VfAoe8farSy8tq71PBbpGCNSt2oJwavvxJzU0lRUtgMLnhrdjCGP3Lnc15leP1B0
XrGh2+V9HB/LeMHq5sS0kP/Z5d4cCUxdlmRmZghXHqYl2qfZHXvOHZiOa8gup9p7
dQyolk4nN6yDEti+j1duvdgFdrqgr7m/zbCCjLo7KxFxKJfWBmWBqcMluJFjHQcX
lTHgZPXaibWrdm+luUsB40n37+9GmO6biMR2B+jCfMu8ZsmXAF6ki0prwvmvzVlt
hVN6IfEQmHDqOsrFz2LENmeKsic2Vh2fAsVI+9UjrCqQU+1t2pUB6GdZ0Me3deoU
4fOaS5WHS6tFgkmNSTBnNFk7eG1ikxRU5JEgfOucz0WNfAx0T73nBufE5VR9rYh/
fiZbJDfytTv8MOekv0WLnEcRnvVohboLApTSFUk5DqFKm/fdZ7D8O5+cIiQGcYKU
RZs29Jfhk7IR2KS9HaJyg85WvD6u0CPX99WpoIMf1FemBlf8LgM1W/n1UozbQT7M
RrfvUatUoB0KPoTmRoB9OiYE+RlWcOLlYNRv+0DHQcLMeASdTzqoitVIJueXpoxa
5wCcxv8/2yym7CcY9gAaSA2/WhH/ATCGjdtxKJOh3q9eIu8rCL/u3g9XD9Ux/3RH
A8qBFjCE+wId79xaqrFf8iEVUhfHusWod8kRUPrdAjfxHEQpKP3U0+mMCOCzk0rK
SqYVJBZV2ZanRX4HQZXGzyVllEsZWvRufMB2htS6Vy1y7yp4zatOnzqHLRqPxTQG
WfyaQmHDOeR0JDut/yW7/GFg9o+6Mj0P4qygJoOqXvEW7SXT7wyyJSOqFL7sScP2
ufAwm69RI0gRU96wqoXuZwMqIhVQZ+XRQ7SXh58nqt06XZOHhRphmARngVc0cOkI
aXF2f9UjFwg44NbgrD5/a4P6B6HVLLBBMSrUObcNO7ZIRKooOK+6HgG9oKHNt+Qf
+eidiBPRDVWjGCLP4GLt3TxGtefnCNhu7nB8HpKQXipsf+FpHP9DPOTSjgEDT30u
eUkXS6NcKXA6GblPwJ4zcpApBT/1Vi5HEbNcATe2hSxfHoHEo8cGGgZDz3SY7Y4d
3kwv9hAWcnl73oD7/kuMA4O9XPIRpEUJcjaMrPrw3aOpxukh++EfTo2xpg/sktYC
FcExniR2Q4lwFgbNc72USHy0QCuWDCQruVUXs2fBOe/J3CmH5wXiShZ+nPjYjTS1
hnmwkvGcadz6RzcogakqLbkTpLFuc+A3x+HGJn+OgNYnUvaqa+f5qK2m0V747wZw
8lAoSAQoNuMKJ2KwVIxxsmOao/JvNOQ8Vy4O9A5QgZcYv7cI8ZAUO8lRJ4xfuxvF
akS2Ps3G63rxCVmya5esUccHIdf5mXhfAYi7NNrL3Qp3lITxlILbA40zg/1u09yb
RolHe90m7LtFf+eApXuHcxUKGC0p0nOPDca7WC4UYxTeL1MaN/Oayhwxluj591FT
9SS+eAKTj0i0W4d6IfvDL3FzdG5n0JL6qt61vsdcUqUv1v8i38vGLOeNo+moYGgI
+Th/kHTjCLys52oQFwNlq8vYnZcTUhILvnsM77nk2DRNBx2+8iL8F8qMm4PVPD3b
SJ6z4XQn+xV+sJKITW7IWOSIGu3eOu/L3PfZwTW8gBs9Z7o1grq44OpJH0RxGPyY
mtOGGwtHFQNy53G3bUjMIG1PShVi8jucPVr2lenPsbhVMuw3bDeWbSpifMlmELud
0iZDdh/ZN+82N8+tsw9kClkODbTgu6N3sR3VAfiOaPDDm7bSCCpqlmD/HgpP1tHx
sH7ZSp4el+6PaED+ZQiyn82/VcYDPlFvT0IvnqvC4MQ4Oe62zKofraCNk/C27FES
c2IjuibGFF8K8/QSaPkJ2m0DVV00Ijpfu4RNOte9X/UFvbNp6JxK9dFUBBLdNios
r+hznnDCmhNhDMLbzsagUT4TyzZ+BLUk1VBQ3Q5Sff9piwA7FHV8Ar95rsAP60hi
YLTzFRcA/qPtsAqBHIxDsns+bePubqrzP7E3Zxkodxy5+TwVqnMWjkasFE2VMRWB
kYWrnIrU4IxrMcXsftNqfDH8CRbSpEBVaDEfKBa4UoScbMw4wsfefPHlECEBmKIT
hrd2xsXmDfQBBUAGmvLZ9ojDtQBXqWcej6cVK+w0xq9PoXL+Nfif9l+kk6gncB+X
1IWrS9AdE59Cm1B3gpkmvsXmNlM1rGQejQ1t8jh/mqs9emO3zoE4dxDG6IrWbuqv
TsCAd+IWTRm2YCv6mYZg+oUJ1uU4MUWc/bo4MP+HLJBTHFfPGnijwmYwAV1Fj5M8
F1L3Fnc4Y445zWz4DAREkVf07PaEnsxMHn//LVUnMHR7H/jFGjaBDeVISa81YWj4
m+OZl8ZsbXiQQY+zuCFfPYeOthCgRyQ7Hde4g5WxiBHSmBQwB7e0C4EwPrPj4Q3b
ZMlF+aGx54mVu8suY6bS6qYbxFIV1WkgHUEO2bBwC3N4HuZTDlhNfngKnNpiylE7
MMt1x+Dh4/PaEALew5ORFq3DG9w1tNNylzc1Pj7H999ui0l2a4GfKvqawG3Ugd3S
APYM+ujQ6zwwMbY+0XClmuCbIsXOyMZ0r6q759Muh+hHGwxL+nwp4015+4tX2wJx
nhobJ+7hXjSLs30G6Z0TY5+BpXRxsQSAyoBCB9EwUmMBGX8MprUCElktJ12KI+/U
zUTLQk003jJqv0IKEHEv3XYdI8eZm0V8p4DLOOYZVKQ9fga/Ytyrno5XlFVAn1Yw
azHzO8YIfpSWXotKc4z0pBUuMjRazvX5RWtCBLeI3lX/vNf8wIqesn6OIscQlLF6
PnG6HICFFvv03s3gST3qUMDwJ+8X1XJ+MLjspkWmHYzZDhqhGmc9YptnFicVHPLQ
EVPKMUgUXVEwX/H931hx1TLQCiOBq9AoiCNHNSHXdiwa90yVc6hL03k9ErigjHrr
SWulVjWZDeToPCne3cxKrdj9CZmdo+H3WMrOsESGUUVOhWRu/PdKblfHTfIfsv3e
gmfYzqrxFCIX45YaA5MMiAywEU5drgAirEOuraSOETOagIna8X3eWcvxLi5X+9rg
MGs/PwbgVHqOUnECa+gbyP1cEPSbcY+Xw0YgjwDGyiQ0ycTaslpSqqsniyU7FaIm
kpA/gMVFq+gXlzVBXBAV7ClS+6ssCkVgw2YnlVK7vvtCcHT+aqZ51IctvtSk/JT0
8/DyP7lhI3eGmptheOi8b+iC+ZAkIMakSq65qNoCE7hXwthA7WHbnpIXstmCfmUS
ngFyDFtFMH+0r9y9m7RUbz9s5eV2/4We9gU2GlIQlw51RbRjXqnp947xKGh9cW9l
yKNjZABApl0wnDIVFaZc0i+HrsgYrLBHkOeFYlsHF3ZOjaHfW9XYfAaC6JsLkCQ1
aYKNIu9sETSieTurNZFr+slmhZzOVTLTpglLKhoGF8ZjnTR/urjkebMcysoibpoI
Ias9koEfHgK+7O6ftCh5DMlj+zpy45oQRPsrmeZu2ujZ3cLv9x2o+kCIF7+Pf88w
o/oPtistkmv+iL4iOXalU3hlWv9+XzENsJJsDcnXzlXOrciTZ4Z9Q/klqlKtTPIw
Cb0x6DvQv2TTRrw+L/tKVyGJ8rnKSYBqy9AVyZyPBO5cKdTVGdwAj16lf6/dl7vA
LA3ucxqa64Ag9VyNQxcd2RLQVyPNS8Lt350bOrDU3FvejS6yBuEeAEU/0k7osW9D
8YMqro6BWVIaErcnEedi6bSfwXUrZ5WzHf8xQLIZoXbAL9tCiMCHgD0T1Gp7HmP3
/IzvqXosH5GZE6VOOVw2vJvvP3CqEaDjaouHyUNndkgkoJSv/rXwHwAGKBUoM+hS
8cRHBfPQuAwPMRhIfe29zoPz2UgTvFdDEwLjdq9hCud4UOyy5DpdsEY3Lx/rVq0F
5mV3BTW5cQYXCECY6qdPspLdWXnUU3VOjg71dV+UZqXtBC9LOAM1I+qiLrs3cjkJ
jHxhNH6kycfwL3PbPDDl19RBlgYZmT0Ha0NSWSBjak/CVEQOyog8xoBg9TL89bNn
tlpJn13HZb9Lofa/v+bRFr53n6TIflf17XEbjuqoMDqN8J0NkoxjNa38HS1ZACjt
mGnmeGIbdWfepX0OlDUCbJKgLb8oCKozGAkYLs3eL/5GDUn4pwMe5comJjW0yfSO
+qqPagsukKyzCWPSpKJ2pBRzIcxdbEDdxXUnXrM7lm2NXO0bburIK/A5KFPbZNlD
88MjAAqdEDCRbMJKJMQV/cLu0Lyk16S343gjCvqfJz+EvJ6LJo6DPw7vXkugh77d
GdF1OTmGWvkZY7PHqEL85dqcmGE/5gXGBYikGGIgxlcId3dHIEnFBNqOpU85MKqt
B0bSWBFloIlcEGmsDjcFGPtlIed76h/IWTWDWUHLEapG1lMtTKfJQmjDgMXn4Frm
s6quRRsvadsJ6Ok175s7+tlMITgh7/vhwjisK33pBTe0OfWE7ZPHHR+Ic4lbBDUY
GqwOk5jg3ONU7yQqr6NUW0aCS2Oyz6g1iQlqZyAHX5nvPzO64Z7UHq7MQbvULLMi
yX+BVkq/dh4sfy6nUBhRs5rV3tnjkvxZ/yxwDrMj3WxfODMvTqW08gn19sHp7RJj
Ua71/39a0MjkzWcGBwRXfMJlwoPiRHxy0+WCrK6j88EdD1JQvtipeW2NKoT4kzrM
guuFdMrUSKQFHwmBOgxg1aUuBynPM8/odpYC9PooNAaah+9uFP2MPpr+AymgXxmO
KPqFkUvG2XpnDIVTLa9oa+0ol2yQk8QR57gKzMamwzeNohUEiNJkjw8uMLmQCBg2
9/cn4kCHpZ85MrEaVUt9z3OESsXR+4xnU6AScMH4O9IM07FmazLYbMojP8Ki3LEk
Yl59bej1lUwdyajV8ujVdHZHFSPFUrjYIHl1fGMLiru93yJaZlrMm2xRamN629Cp
4TCyvFHTp5RDuT5B4SysNfXRZK+Sc+FMk1NtObRiZetXtzUKTQOExqQxB3uoCQ1/
zOX6oN1+gRy19XrBzRQK/nfs4XLNsnKfdO5KtkcD7ddvbIYPwwXb5mnUElmKOKEm
Q9njIc8I2IfVIXViplX4HVXEtsvaOk+2XheD0g8L683PmX9q9JXzw0ha7MlqcbhI
alI49kkbiLS92zF6Tn1PHSMJpg3dssKwBW2lOfwmjqf5NvC0czhbzLdIc0N+OY+Q
jl8XUUILO1a7vBn5L2FYaUHIdq5cEm9sryvVSgPrIe/WdbEwxFnpv+MSNdnVTHpX
UfPneiLt6c8RYVbzbJ8Q+y3p4rJfRyzAWJL47VeQB0rRPMOPkeQoi+XgP3AtcW+B
B+OVJJwld8ZdWXy2Tevm5Mp8dJgcv4tjUAT6qD+w5dBozlGN8CA3QhoUucK87ycq
N/mHNBk41jd45s5/Uy37r8bmpCfeLTwk8J07C6iUyyWKNaqIUrE1/QeFjKmA+3Gk
14r1+HZTBrUUWbqlVaPIr93GoJjJM3agkFhopLI9hnph1etIkgAm2kajPwwRA6qD
c9QZBFFi/IfVyENyZWS8Z7LN5zpKagBde5Si4dZCTcd40/423xHKTOon+37FsRiM
iGPpKCrx97BNB0rrKS0jiAluvCovX8eOSkdwbdwkDJhxnxlTy6pqHg/gPE5tPsw+
B1E51KTX+dFJxIRrxlO/EIrieOkjeo8WhZzZqhi1Z1WkqDbea/8b4mmT0VDyjcjj
j5Wg5ZCp1G/rLWy9WMe4xOGDgXnK7Ff/KMywu2lp7MT7wTm+OUR++0BFNAfgeE7h
4rjJLxAXKhhRau5Fw77s9Uq6TMLB5W7Q8eYnAjXh79SBUFM3iUyoZMo56MwOiQe/
BM/aSYkcP5sAffIjPdHaBy6L55TH8/5E3KnXRLs48c/Gm5Khu5GtDAcSjOWD5EXo
j23R4dWEQ+q+wNsYlSn9krlbjuy0OBcKx/5hDatsPkwZ3q3/Mms5s5sq/q2hifcg
314cnS2CeMBaBY+mYGPWE4q3pYfTJ+Z/Q3PjKUMILkrguUNS23CAzPKa4djdeT2N
LB/jvIAH0tlO7Ap4HnRv1uvqLd03p78RTfnGcKTcpIrXHZigQHXJ2G8iidfEbXqP
LqfQTYQBAcJC0QjN611Pbqk4pdAuCra/j2YJX0RxR3UCq5lbNkeD52aXEogmLLb3
o3tf3q2MU0JmdiWEIMaQNlRmUDEB39PT0FLTO+l5i+7kmRggdpGQGHHcGn0XEW0U
kWnLtQjDnVv1RCQd0cHI7DCGpXeuYNcxq/pBf+5MTWbNkYBW99zYOSNuUu0Y17rE
3d9I9dTAYX5izKP4XEESPnbWqfcGuo4xxS83wnhTzKskBFrcaEILWxvTA626fsB/
aFLkHO/OwoPv6cgRCJQnUI7ekMmtXcDl4CJT5QQNfK3oUrXOW+EePncLchbzWbkW
Oipej19KMHp3xwA/b3g6Rwlto9bdtdCszof6cMXbLbn5pnHLc+EhSmL5vqaRKcZF
H1RLIUWyw24tcC+fgd2QfqBJMhSLIfQMBSLBAutm3Wrkp+9hoxzYFzRa5H3HJV6C
2EEN6Wna/wBVMVghV8Cu80OONQDY75+Gz4yJKj+P96J9oqm9Q4QjQdIdd/jy/5rN
bUaAXwP/0XMnQWeKvnXo61brmCHxYwyi7kDE1As1V+8SpbKWa7ksITSvk9MqFlFi
n/iAztGW9ScERrtxlys3ziejlkU5I8BxuEj5iBgPCCelYadnSgm2N74zAby3qCE+
6BbuFiJ3uwNXUZzLq0eh5C3LKy9p4NxqUCbpC8G3pWq/rubinwdj1R/c3UJOlcXD
lBEQhUgbchjmhEMY3kJiA/KWjA+Bxb1Hk813fvtLgS9+asoRsFmRH6vF77pdYQ14
ARTWq2wodzkwvBuDopVetOARBKhTE45JcoMxOYwoxENtKU4gycl732YS+3/+oKUQ
1xdyZiTTsFFMD92iKAZnvVVgX2JjUo3auQkHKm/w9BMn/uYSt2K24oWBVlaq1qR6
ndWd3Uu12qVkTkY1e3TqidlbMg0VtfC4QQgPP+PtWIiCuyP3wWQMM2WpYz2j4qiW
wrt8AhTDQsYXX+KEgQu++CzkW9n1o/GgpAm0rd80QZCkmf4ZeBblWJ3yBXFqqbNT
Zaf37u8GgM3QqDQQb9wInZgj9OtIpINWDy5R4M3q8ve1Ow4jkcU1XVPIiaeH90Qi
0yGV+qHdoaGLS9AoSoeu1h75J+B7Rc1SaCn2opaFddZYLNZMBixwRfqYwQ5mE/9m
HNxi2n7wdIvrfLZJ8k9REPYaYlWoSd8JvDXIXjJVUYKwzZ+4+ZPZvuXzWGci6qN4
gHUNUo5MJj4zyWnJGQF8A8SmvHHjSdbNfn+Ud4TeEvvouC4LN9CjcG+AkUFyrlu9
1q7uRP2+75rDDe9Ym8hoc2AmpGV4pP/z8XoCSOnanjiBr2hQnrst2EdLXBAatDIR
/E0pG0eF+B6njeZFCCCtFoe/bV4UG/N04IgL6MCsm+9uVEwco7M/Kka7LsEVoznG
/NBeHGRc2dzIahlQ6kRTIKODmbtVcCnf1gN2pNWRkTCuSSuESFo7gq1JfIkRCW+8
EE2NpwestsYJbSQmox6lDmAgwgHUb/EfE2Pc4WkIWUktSpCX2ZHlCs25RdI3glu1
OXdK0TEqWHYDv6sYjGODmavVRk0+HZY9vEhSRNz/xxKW1MXvSNhO1slgXG908Ko+
F9p8F6wNYfhesychZFXREAYNEnXOx23BafoJCKZ6VsQGlNBhL/OUWAN+yETRp+w9
+NLQywtYiNQZb09rokcUD02ZHqfqOJRnIoMjKM1fyTrcYqB25L9MAUtI/3n2KxGT
kOBirmgpGVJCmPt7OZlrQZNR9NJBmhs7RjG6pcxVxJle8M0sxw3dGN3BPIXJbad0
lV/9h/IFiSuFFKKWeIj4dOWfoLYdNcPpo82yT6SrIlLeTQZdqkVXoASjqpLKsKJE
3xlFcAPPE3V77+P4eoLknaWlamCcDA9UghMFPCg8P2NKxTPXjLgP0JWRlXcH2Jds
Se/Mxfhw35K9ISibLXryF0gxnXapGpvW1e/Lad1w5oFFgORcEHMsCBPVNTUbWJ5/
2XJxQEeHOeaURKZwwfja8kyEVuEO7iz4ScCrmyhfAf4MH6iwK5xa3sbAfXmmZkSL
YrDugKW0vd3XZpeA2+WB7La4lj1HJD7g8somDNF3VygwOSYMlzGTjaMhv2mQNkBm
QxTt9ovlnwM6T35YWZMtVHQ/Rs4cx4CNXmWaanrZkaUR1p+A5JqLhF6q1Xobj+46
DGzSdaiNV3/yJARa5ES5kaQmQQKrxZjWzoaNbhNYIRRJHXIHyqDeK83AHno5JNR4
nIMPAvmw/YZ60z8hKl4jdc9FJQUQ3KCjX1WoVDPCP4SlIFxteFpmn/CrP+lxe34V
Fduryu7HFsyxWZTVHQkQ9LSNidKIGxwtNc0S5r9nytvTbauZVhcvy+EAwE/2Rziw
kwUq4x/CSnh2MjMvpeYHX2r68IDwvJUx0z2WzbmfD9xRVnUY5kuTAbFSYe7s8FF0
qy2UM4WFn5lrjAeV9lUKjSCB+TjQ0ShE5P99dP1U353prZ+//UC6QXwcquOEc0Pq
gxwfPtbemFf8Zp/CTc9apbeqKKVCocTHtcNHyAvGeJiosiXN6nU7kQrz5WsY6Gs9
yFczaln5ykav9FvvjmXlcRAsh/rQ9fwXGhN9igpZ0SQ2oHL8ylKeZAriqi/00Dr6
6BgjzOU2EgQZA/LDSR0p4HUSthSEvSk0IXP6zVRdfMdqhncGj3dbRoUaywpw9nXM
bgXGtNBus/n9MmbuO3RLf0ncdNuMii8WY0zS/EaZWWY6YbyXRlJs8HapCDWoqlJ5
Fghy1oqSIxuNiTF/MS3BQ+3tDB4T7F1ZrXGQf3gK4SpbALGmTG+aIxPk+yNh63cT
x23/utrv8lfGBdve+FUcAkC1AS0VfSf9HH7Y6wnCdYMVmTIq4d59uMd587m8oWdH
ma3s76/jj7PMFBEu3lGlipJVmDawDKV+GjfUYN9YYKkkM+nL1VzRjUs8HEaE8Usk
eExtAA7xnt1IFL3n4kLq1ddOmbrS8dX3Hopw/LjFdZSRl6mTlmgo2MyzXcq55Jk9
/Pp9k3raaiaIVkcvFkWin76+n7Y2XmHtsPJ1uO3zpLBI0BHNmndnlMJaD3UKcU56
60oqvlHuJV7xRHrxYnLuaUBM2jofwcBwEtBCoJpFcWMII0U0V+wh4XpdVXvDl0Q7
oR82iHFKUA5RLl1pfqa5JgOBaVabrciplXIeOxDHTHnx4GmC52h4BlPpEcjNjuVP
3GIBp7Xm0Rg19E5qgzGnP3Bl9Sm+mrZaOqbStx+RIixIwtgTqRXS8u+64clpod9g
xEjsnjn2bHA3ZnZTsZFy9zWe/lR2+ZbslgIyRB1xWfpzRf0qSdDbz0iexNH5fEfn
YloOSTXCce5p4ewFBz78YobG5LsEwyaU983VhRauhFUyASbxybyhVVw3nABjPvYK
/EQS9XCvNZNDQ/leLKFdpWdNZzrRhsHWHACXUuR2q91u41OmnDnSf628C6EA2Ep2
AiyTXsEaAig7JMDtbKBN1tzi2zkioyWmZPOdJ+jx9wwoXm/BIe/T8ACpxyhAuVIt
p7yLB1GNIeMIYt/rXleY6yalhFDshpf35pYbNSFxujj1GD1mRrXIpm5P9+Qcux6T
6Y2pIjqOn52ABRXCjC3K0Cim2wwlJG/u3aoFNfot7kdYeZZZSUrjuQuMClWFrrCu
PvzY71K/LKu/h4k+Iaxr8n3h15Sxg6R5Jf73nyGvntTf8Pg+DesIHLolBQSi+PrE
8iaauFPtXxQKVo/lWaYiDy6GhLwOjjO8OfAkefy4B5kgTosHnye6NQECFTFnLgjI
cXEBeyL+J1tsa20kV4Keo73ol9cLP0gU04UOy5YvmiJqdRz2n14UOHyTxr885shF
EUyG0r774mt9u2KhBML1Q7O+TAdCjffMLQ5W70JOvNZXTP8/I9dVFXuq2dYyr1UT
IQm20TWqIAm8clTCh+j8xQvdVTcdyIflvInAWnb8D/k3xp0hYgi2rNjw1bjLncR3
amcJesK1sKPiOKyawzC/X8+fEufg1XJVAcucSiEF5kTJkL0awia5OqVUJkPQuvTM
peXJITBKrmukJRaBrlksZ5wdo0I3XeYkIr3rCaGawBRBE39XSduSZDP5dOG+wcqe
MofvZzjeeLSszvTkHC99lIIpA5kewbbUn/BMNtwShv7oGxGmAfsJ8iT7wT2MHWhl
TsKETSiXpryy3g7N8wwNKA7bNs54fMpIz4MYrIMTaLisLMRbPQ3WwSco6ndppNsy
XFEYUVMvm4BP0AjkamFOuNhMOi561foDmvJ7AXMuuEQSNS2JNhRlj2PyFul8J9zc
fQm7ozAF4L0KPRXkN2YoQAR3Jy8GbNSMLh6KgTbjspBB0idsNBJ6YTlDxkQOOb4o
yBegrcG9+zDWuIJv5OwX6rRoF8ttVRrEuF8IE7XM98gvHvs5M75SojJURukjU4sr
YKNZU50cDXEhOj6p7nY4PTElBQVpjB0ucptZfO3HVSw1N7KoQCe9MATsshNIEEiK
t0ajGkYbXjuhqrMYZGUzYQo/75Agvl3VfuZIOY3gGTyI5qJyi0BM7wWRj+9Y2TFa
4oVyO6P+Sxg1J3DtviS+CAC6pAH055WWe2agNk1Aui0bk9qlPWzx/7j20qX9Axqm
k3X69GfC0rEbvD1iLUDdN2FR4G9mmw7x/Pt51cfznW1dTdmN+puPxVO+mQZLwF9r
+xwS6vfP+9m+1irnX0oop2FTHpRsqiqkyi0UQS8cqkZ9HFfm1/Hx4iB3gvLbEYGe
eJHAhIqVnGGDnC5nik7VpgT+cCbmCPVP9Cc+15/EOOEcU6scER6l9xDVe3G6MGo9
1Mj/EI5XaMjQvEs0GH6vTVy3++LJ6zvMBAkPZOh6WS1yQ1AjBsMoIE9CbEp5UUwU
zSZbgaHR8pKMzhhBsqqjk4exjJQyI0Wxyezl26qmk3+eV6bFcCW0qrLBZVFgOBTK
CA4dFAT74HkqdRLqdFy+vxTU5QlQYnI4uFPBtKwAqqM98WaXTaL+jjwkjgtk7qya
QNSQRGvLOgmOrwTbAOJXe5MSKVa8ozMMlVvT1pF5oTJW/i0n00cTMFLkU49pEQiP
815AG+mWJadET8ZuOt4505WxBRTxhel13ywjUir3qW/afTIZn1bt1ZHxrCWor5aW
z665U6yzkBeemc77ep1qWeLwwFmpOdiGF+c9mpxgQMM8Q7XTNDmfAvqvBv6nDama
YMShdTNvrppp3sejqg+5cb4n4nNiwtZCGtSRFmMCBgOAHavTp0xOtXx7ysf2iwPy
sfvpyIJK67UW2I75YPSG5wVEmRj+9Clc5J0HiNHSDjiS5FAsNLk+t+hSxHDIDYLG
x08eVldL4d4onn+Om4VzeawTlT0xS8EK0rprIm8bVOavJEIzVqQtB86huNECwupg
X9rwP92z66xKAjG/++sg495CnMW0pkeYBVDwC1eJBMANVWfIKlwzwCy3u7r+JBNI
MAGBpdnhi/ovo4dcrOnNfhPA5aB7sKjq0nXUtI//+lZPARChQz8IsEH3Bmb5oFgj
P9pzVRq2CdHBN6lAsxO0717sY6uZ0lOLop0yFewQPEh5dlrPdt650ONSO8yXDkrs
Rb02eCxkPkqF/M4VqI76uhGMzeGzTNU51212thXm9NR1xJbD3bhcMEg6+dkP3/6J
rFpbBJcOlLUOERCxmmcZzNIiNO9kdBr3B7Htsh40+aMKG6iEPvfnFBoMUkQmrjer
XVyrV8na0++cEOiobRL9pLx5yQ5kvG0lXTr1Av9yvXIMTjKFgx+BIZzAw6wvHBA3
0EA30ORPPa1vWqYNelWklhgP+ZTymtwpG6UE4mllx+z0pvpWzkv9U3IWdceSADCX
3V+x0k5gRSbowOEVdPckIMhTxe8aptLzW0ogMJQJdoMyeY5CW7ktGLmxBZpBzVhr
PofBwLNxrvXufB6y06THaVOAGWYfxSIBdpApMr02iQdZR9Je0KzMuX3OASw0dnF+
RpZnr1Gt+Iv+S2c8Zu9B9SONQz7SpOW/JCejvYeX4kcNmDkpwePU6z8S7UMWC+ef
g8wn4ZHQXk0ycPVQRnZl/jhhakeReBYkLmngWogNjSo6Tgk0rkI03OGl6TiE2plx
j0uiG8IBq6AFr/BwDGzzVeEo/KdN2oa85g362M2MvpxXJGLbF2rVQMYgHhuL6Ogb
3G5WIqh36awjxwJfamXi9E5c3+By/2GohPZka9mVwbzzeWrknmmW57vOCxJFRerb
bW3FAAwf821XbcRCrcD9wmcuqGEz1lT9GE4f4LH+DzJIKriM0j/ZXUED+G9f05pm
igQOTbdBCAM2SgojWmYMMwq+kPBbYdeBTIYaJCtGAlnG5I2O7Egk8owNtryXzgU1
/iXYdQw/9b0gsxehQSHgr5WVV30zsjClO3jcR+IYf5lJPOW3SyDxziXUXkuAagtK
4CPoD6j7VT+69eswVzGsRTYHM9yRStg78AkIiYjdeOPT/IY/cBuQVJIo/RednBzM
RuktqiQUImhh88tg886VJsqP1ytEZbSgE5RbAUYeQGn3p3wjdCmQzyEUoauiYahq
aIXdRtEI48WSKmwrk1HcTbw2CCxsbL2mO1UWfQ5wrwT2MaDBDcSIE8YWOcv8+aRg
bYKdjfk9Ra8eyW6m5Jq572p3bzjev9OVIPnW1KuMRNBa0i1S5dN2iLG5CAt2QvVn
f0XgLK3S6RHXMmtLQTutE7krV1ojveByToT7m3uFxGOlETBcElghlNKSdhZitFJ1
FsAX8u6xU5SOsZKtoo4XM9b/ggT6Rz0Wg40bTz/+CMIPVOmvGpGR3IXK1c5Q6uXE
qOWycagnmNwv7gb1H0ACQPSltnqJ5C/6FTlPIWua13SU+IRsjyEnCWJs0PzfqG0u
qcMUmZzLsLcOGTPuDv8jPHQvUHYO6WYFhZq4TJy4OTkpah0TFi3pyddXcg0X+KUB
qJlFb9/u27kEv0Oft1zPPdZm20v1z/bRLnn3odvCXTtj8ILORe4RvavD501nljE8
dwEHPXCLk/LMrUJZkDI5Fl5fGloXpEKinUwMd++O6qXqDaOZYMnElvs+o7mRfsUc
O5vtSNnL9vngmcIRONzNG3XkYYWaYe0iabOG0tcjrMO3InSihtRwAmCytcGIJPiD
Z90y4FjyGwBGMEu1xPhoj9FHeX5Py5BDEUYUazLNUcGLzXIMhttMsfZZKzEQUdQN
8fb8Nnh3ME1UAXL6O02zeY3FzgCTkESKJiAmjC+i7p79c355E9NeTvSWgWVcyhse
HWD+SxCmVRpTLZbwUjCDtI2iv46fOU9BQD0RBnx9RwVO+sFkh6rw7QvMIrcTj8MM
No7WZc/pN509tkHRxWnRZ0ciRYWpYc38U8XeOQo6qes54LV3/p/vJweCMbaNUN6f
GSs03Z3LihM+aOv5wrBKzpE2z1mmBn2BCsVPUcn/00gD2SUzBbzP3blujAf9uhPT
htn0nAjvmK3szOTVscEqpib7XgTp2H9pON51mfM8a8uZxUJKj/SZoS2cAeIXhyf+
gahbQ9z8QeppXE1UNhdSQ7maI8ePcaJ4MRaqlQ4AWwvIz3EpV6RBH/CJat5UPcm/
bAdA00yM4zPbAManljLWN7+Epu0nzrRCZdDu4ov30InqFIUH1OxHVHoq7nOjsv2a
P0eVP426II7lL4qM5uW6MAn3dZCSwhB07OSc9TXFDAbKIlwVdT80hNVuJgqd878K
9yfpTDe/DycOL1D9Jyjb9IQxENRr+V2HwA0vBc3weEW1R5gJgyFokBY9GWr5SlN1
Rz0m+6NrXD/YLTobFFtvmOnFo00+LNOBMYUB7P6y6Lm2FLexwhW509beD1JBmqc5
E8sLX95TDyQfBw7mygYABKfqKg11iTwX5vFO6OriK3eyOvu9J9qklh+od1qChQXn
xjsLuiXpFWSrIkUlhq3TDAiutcjXyecGTBrqKw8zWRYqgsykb0jFd9YBmMzeSS3u
BXj1+LqAsD4EonuGZoC+F/CR1ra7Z8yyv2rBQz0Q3bVN9gl7DDQI5CWaE0+VDx3Z
DcIidjLzH38v6BgGPLtU65JIdOwHCEBmsJ7pS9bWfZ4ekW3IbVUg5VlbFqepmXO2
TW+Tb1P0D1zjm2NK/PRpoGmJ2MvaDaGTtOiJk/nIpyoXc/KQj1xzXf86YG65HeyN
e0GV3uit9E5UnJMP2X06tJI9bRjpgoJsl0uKzmWEBpKljFoq3N8Ht7v3xobbwVef
/ZyQrulAC6SIUkyuZ/ZpXAX16UZ/javV14LytQRydiLFHUU1pJJXRqaIJFCsVpas
sM2oPYru73wdkuCblSyL96GMpolSCjmtsFwx43TTqk5Hj0VBFsZXum/EzKO1ePFB
j3cGiXF+/7WTGqpWhml9CTdq1kOIh0v52X5Z1GoYqmCJ5smgEuN1bLlWtlqcRl9k
2sF4tlHAjQC3K/Zl5BdQU2JEKB5aQgm5qvOvuud6fAZjDRSTv541ledsQAFMo6uJ
mCc/1PnhbgMAXIeEPQqMe7eqiSc2gvPY+aSmf1Ut0GKXXm9thHWLWYHgJgrl4vQn
pYukzqWzW4MWAXmI3fXvL3CrOzc1TAtIJVNjWmNl2iDj/KW9M88QkZnCW4aJa4mW
ql2riWHO5fgiG6qN1wavIXIjr1k/vyzDwGj04HLv7067t3zNhNtk5EV9YDFjItSo
4rRImG99WvJPSMFFXD0fIPdDa1YgZM2d496M39YiWn4FFqHaQZJJfAIIV3jQjguT
c2Zj2iDj9ml7yhk7nqi1VNaWTK5Hqk81GpeLzCMaEe3u60ZjY64k4L50IgP1S5j1
JQfTBDd4PxF+ShTDxeTJvsRzyMm8UMkyt+7a3hUBZjSBBc3ny4cJvc0gz2Yxc07a
tU208FCT8tdiJzXGNt1+v5pEqZzZzqbrL+N9NlGCyQ5ACMVaa+/rSz0lB3hCcRth
O2vD/MEuFSGzbYk86cEvw4wjKQWi/G2RLC7bxQtUI8XpOcBZW5khXDiwShwfLLbQ
D2PhEULCTVMBXVJPIlIxNHjrY4w4g+ANgodM1Pw46MZhgt8g5n0v/xIlwAAkDxAC
3U6dQMx/eReTkOIdnbpISIvs6yqLrvQc9fKKqFQCz+I0A4jEeMXzJtr6nWK3wntN
lkTv1TGAZvzkKgV7ZK5mqHDAzKJcakBum3IVMB/rkOV30gkeiNWbcKErl9fYAnY1
q6qygyY4phEyxZ7Z1T/mCtH1XrGHJFHeGdlAIJmpfs5wUnDEzHOcxXjTvXiSSBSa
ZWgf5Un9Yo4ux3tQ9H7Sqc6lEJlBRl8wVUuZSe2j7+arr6bCyfsdCdXWVpzBM7KY
739jm7F7c+t6YuJoSzGOf3oBntO2HHctvAfCCgvK+bQMdfciITzVt8pfejMH+CYR
VgCX2tqNGcfBqJDRs6OklIG0YTYEKXl6mDJRPa2pGvNp3A/UWNgwcZM9q1OAW5ot
1nG6Fj/JlT+YnF7d30V86RvkXyZsHTP04AQc+tUJlslh9yP1oll0AA91+a+zDQO/
JGVZBOj1EUH1mADpJVdmdPp/sWgX4Bni5yHANTCSiKEkFObWg3MnCLsSj7LTben0
7ozOpqnjH6/H/ZdJxyzqtpHOGBefS5+E0zOp1/2LyUqvKiqIA86QAXrGJcJGyDB7
4lXcwByi+5lGU7vc52N8FDBVW3dUmZTtclheNLFPZAz9/RkVlWYqriYDIj5lL0kQ
3QN0SAypZldMDYKexqoB/5Yrz44Nucg7lS3C3MoQtnTjTKDoP3hULfgcdOOx6HC2
qiA3wCo2pRdwF0PQ8Y8co8yA8z4Yi/JF2X7SgPQ5QEGGS8pqtVAtWqrYCSsAIT2Y
6N2grIpOvc7Y7ozRJsPnd1UBz2jpNlLzAkZGE+oWRk7pi+yAMjHCLGPufu1RefFJ
XN36DCej+jaxVxcwJUMq7hZb4dYVhQYmRzDNECoM2JijQDSm6VygAur8Bamt7jKD
16tKLLZVABac0lAtwEHhpKlF3Fh4dUc1dckdT0pb+0m798puZJTENHxSaf++3hzz
/a37rGh2St+W2kO/oMXEJWgoizVSv1qJdbyCM8O22kDnp52GsKu7NZtcegNa66w1
YcWwEDmkgiZtw8ZkLI7lceuXHgyCzFrtNnA9H+QatwSBIcgSSwlHTtFFrDj3xeMq
ARx1KX9PRDveRDSu7/95bw6IKV/splmE32D2QWpzFOdZJGngdELNQIUprQJda0Ol
b5YdhnSKCB99cmiPhstqP6HYYgvjzacbuq6jgn7/XxUMw/c9le3aaQfCRd1ANGvI
ZnMwZjZ1VMFngm7apLtt7zyA6O+6ReNCpT+BuwR8074yZ3zwc1O4nKNu/u69jC+h
TAHhJyuNh1CEwy5eewCdGvdFOmeD207aqictqzNB4FXZipO5cyV5U+7tPDwelRjb
t+cUH7zm2nYPEPACMtyGTv3g8DRK1PZwYHDN8EyUTs/7VPRga8wRgOrFTPRH6ogf
CAeRe2AjryJnTq2E25p6F2n2Vqld6dApHr7eE+6EY4cw2yhyukqq3jU8WiCVzsCl
y6BMkql4IqnHR5TP3wZx0Btm4+Czjs8L5KKrKH/4E2XPw8K23tzAwy18q66ACcPY
FzMfxEE9PFSCETtH3Xvpla+tnHuMauk/eSB2Z7/XwxmjSVYiPDBb+3uN0Ys6CQQv
jYlFzUkzC7uH9EhXGK/Im6u98Cgm5ZLQEixMZ0bN7XZO2CLHMHqHR7xQcJJuZTGf
pEg/I7rdq+vxU1m3bFA02yBKROrUl8R8q8czv8Tt7BvsHfx3yZ4To+Dg89Jen7YC
86zywxP8zOiYvPwh2AXSnO1yZPtic9HyvSsLtb9NdliM9M687nQY6MxZLZcGVEV8
xP6xBgcXZUNDrgTpUYRKKB8cjhOzO8BOXqyG6vdPlr0YZs8VeKc7FUGxLyX5iQrR
3zBodU4ZxJLjgi3hYJhkMLoc7BKhfx5VC2u94iFnxhBEHt65UqatjFd2fGBzPE8x
aatkp75h4EnRQ6zLKQmCFlL85SBSP8hHL2mHMS+UHqPhJg0tGp0I8g12VaD/52rS
zC1RJTjxHx0WKeZb9Cn6DpB08q/Mj+0sCZT1Xz+ZpBKeoubi93+gxjj5C+ZOIIYH
RQ7SXSFt9WmNGDQrdp5LwCYgLDg2xIeBIOgqfKL5XfrBMspf0kFjUKi93POYqBlG
isgJBcDnMmRikC+65dygUj3uusNeZJfPqRysgSU/QfwfYh0LHNkUYugTGXfInd4Y
x9GF1u2Cq0QQu3syCD/TBZzkmHHaaM68evuRcVh7hFVbzdl6jmGjTUx6cgKcpEA+
Jk5A/Mcv5bZeh1AzOpZmA/PIr5v0d8SQacd2ADi2JJprjlzgyuIxl7e0lJO3p4aL
O2W2yBJ2EBauyjalgtGAdEG8ggtHDFz9bhpyJeN/ngP0J+YJTIbHL0NOcLzMyGlc
PinMkNtA6Tj2+o8TwtN53Lf7m2C0mEED1zpuAycBkUXCvEiMj9xLGOtSPb+lb3iZ
TfH+tDy9okah8k2PhzSkGicQc/7i0C2QaSrSwuzvJDhCgcotcULrKqr31nA8kKQc
jMDlGHm4Kh4hVxAXEPsNzmtscW2CL1GpmHyCkcWk47ii/o9Zs9WDWuQgMp91QByQ
j7j7SMvS2pOtIA55+jY5GnjQ0LJiiF7zlY6lCbnxamV/SRf9XzFhuRwz1m38agSX
HVxhPjSn/8LzV/FOURLqswLybPHAcIGpi/5dkkzLFBdQvtrVqCCt9eGdEWAVknvf
0HIvf3bPpDtUuDT4gogeoNWi5ev5thkElewFtSMqtIGTJWAEztxNYJ8t15kQWe3i
9NHu3F2HV8lHav4V7uUbBhuQX1sbDaeF5R5/m5e8yOXEPTX+pwAUQ2IfUEgybQar
nWNUxGOcU/AOHb9/f1Fj1o9wY4aTiT1xvYJVRAXm1ZUy0h0EUjw5eq2UfWnznd2A
Hq6mNKSceDfU92CQCmkEQp8jiKNj+742aK+/Eh20wcFtAuRjr+IYGlmH/PsZDrUR
lSxov1mTddrOiF/WlnFEXPEFrq6yPFy2VegPxMbZHL3oBc6RjOQzhtTQh5ZCHcw3
exBx6I3zwVvHf+J0fBHOSg7/0cwr7F8+Jza+cUkNsUemd5OnvI9UxFTFzA6IXA9J
dmBNqsvGM0iAO7tZgxveLOVZ2ugm1k/zVAXyDVPQCa0Bb0+a2trz9RYkMqKHMqJn
qI+lafcXa9+xObImGcX5Ddi4edB822rC4FAZf/ygTVH/50S3VrkK/6kGg9KQosJ5
RmR6W5xTPTLoXlIBTTiGjmdWfxqV8MLW/9wQA12KWAABwbYHtLiuHLpciyez/zXD
67Z3lW6bCESj3lVWwsT5ZuYKRWczOv0Ci2ZVeTW/hREejHZcTxbIybiN4WFdf2FH
eXndb/D/RACKAMzCcDPnVLubmj6k10NSaHkMMQsD5KXWp+7h0o/HPRMHb948xvXr
O8jKdim7ZU9YU+817/BrSh7mHtcaMFZ42ZtJw38pF7Ka9RJ0CfSRAsyL9itbWpwx
A84VI/GPNqQYa1qVhYhN+i8m1mbEywMES3hOhJwNXQQ5Hl8YNHEwYfAYG3IMd+qw
nhM5E1zXfEgw0NCbxbmWxU7FBTGTNETiwH4l8aOvYesIcth1eP4ahpAJK7MOz/4t
3sTqf1uxbHSf690GODLHvGsEadR/6LbOleyQWybIkfko3icqi/SDDhNigurE9QR8
FHeT9i8eq/c4ptg6t3tBc2sD1WHTK97GTijrTjZv4wHXlseDSs7etWDN4eXyRELD
Y8HNYU5zwvFizjnJyYRuFTTMqu8nKsIXeLqahrySZ1uB/iDJvtdTuq0luOwIeWnO
j2wvxmPmKZK3UCHH6axYOcJEUR5DNrWvl6PFMh07UcH/mBFsbKe9tKwiEliX8cMS
mILMO+OOltcK28NNCkMboDB9bEbY5sjT4Issdw3bsvumpRCvvLxvDKKZ6PErAUcg
4imlmYVFiy/zOn+DQ3szi1TY4MY0k/tmCh55W+tfacJb7bWx2DbPBB01MRW8g4eR
S3tjkLzF/5iJt+BqH7ZtlFpsTdv6NKZtP2N1l2WIiznt2DKb9UI2PguYJRMuIQfN
NSpvXG/EEQ/KtfcevjRLePQU71INW/P2uG1xGwV8uZ1ZssNCydW9Q2Uyht1RLWBA
YD15f79Nd16vPlVYLwxQvXN7O6Iir+cl4vgZmHP73sJfQRod32Q2tGwFBfbA40Pu
GLqfgQFu8FA3SBHyVEygeHfFpAvZUpjKIPObr9XUeMpde1p2niHc4MBcz0PYdgfY
WhXxY4I/FgLQzYH5JGCaTyTpfazo99jAnIQx/xxg2CxMsAnkDE/ipCPn3rjocxc9
SATty9nK4ZF23XUc+LiGjeRIYKXxJ0l/Q+JhAWIpBzj4yGuo1KZ/yG5atrYpHAIL
gQ5OlHJcIPhs2MLRvP+ICW8UM4v2ij2gokdnzFXSwwCR6cdonj4g+9cK9PHMYnvS
wFoXheEJ63r+VatgmvouWdFB+j36kH+nIW4W0zgrJZdY5r/QqMLnosj6nK+i81/S
RcDQ/EvEuLM7pvjslp1UgUFLjdFjsjxC3d3m8LGHM7Vi7S9GXGj4ykFxsKJPYu9X
BxX4gKZRE9gaK+3A3V/C0p+lMSMnCASs6uxb6m0LdO/1YiqIbuWlzBL8A5AP9sku
n9lls01YEWby68r/ftoQZ2eG1pBTbBSsfeim1sLlmQnNj8KaN4KHCM7NdZxMDXgE
/oC/+wuTC5a+U7dzLrZV6pILpy49KBeOQS4Y+Muab+tOwlHIXDy+pT9W828GCAL5
10C7lLpseRn3Gme1ZIQvgMJl6nQ8Qp092sR9cAI0rcOaxkR0rfT1kBA4FJOSRCet
DoUhDFrQKkWPKV0znXvtIGgwFj+DPhrQJ+XX7kU7Lv1G0Qv1NCxGzDxRJaB7LmrH
HOG0ltgqFchdhvRu4P29YUK2SR9kpVdZWcsYBx66r3WtNoD2avS8Cu7dI54Duku5
f/HVn45CzAebLZKb63M64z3FZI9UAfzajdQvlh8BUQ/tY28FtDJRbXdsWrOkyDDd
OOA1wR+gsrS9jNt/x/fYQtm3IYroPLohMxzNXM3ETUccw7/cCQx1KizCkkO+qvkB
uduXS6qUHUXMzvBAS0S6otOwlf/ZEy4T1urTYQlOLKlBTwkSvQnWzpPdj81aRL0L
SEpGQ86PwHQbbnN/AX5SODbUAZWNo3DO68u4y3aud5B7mnWl7Z6cqIEyGQt1TNrR
wpzZNzpQJx+rDabWrRkdlBEXHLvjGjd/D9x374QmDYUSY7ixQboTc6SHoDDYk9Md
8AtBIk1rKsFOpXhC04Z0vnCPnw9PcOtVGXWX2XL0siOrze6hJM/fE5TE2dieVP6C
tHf4ZRA5bJd79LNinV9ZzJZI4wJKJR3Fz1c/YFlqhSlJ+H1rjJ+4VE8rTO6x94d1
/u+uBrw8rDJP+wcYpKujx0IXMH/PrkTyVgN82bBoMvrQgw0WqtqDbZcXq+QKv6ri
vGaZup8wONNpEuRc4gV7Y5S5BqvqRSrXouQZDszump9/A562C8+4jJH9kkKxYeXx
jvkL6EKGelJipWDQb50YzPHPkRFZT0VkUFwcD0XuRsEhfz6ihl48KeZrrAH/ZQqu
1JokNmU8pYQJSsKMhyNLPVvygfR3g/8ZP5W39Ul+2zGeiA46aL0JB3vcAhXhxEdr
Wo/NMspEkJOwy6UFe5AxcoZ/SvsKMft9GrhnO+41ugqfFK0zsgS3Cz7viSZIQ8y5
Txnrtt5tpAa6QAE3z9oqqocNxSQHJBb7PXLxHfErKRFqr0aiY2KToibSPiZIb9XS
d/ikj8kkYI04TRSiVfvlvlqIsev0aZe3twGBBnINgD1+owsLlnKU6ts5qK05v9Ap
yyLPvJvl5vu7qIF3EkmChKdJYBDAE1ZRFSdc8vNaETHIAXOgGnb3Tmsg1lO55XXF
tNOdbR53DDokKx1DrShe97S7Hrc5nv8DoPs0MXWWMdWSHp+zWr0SSkn2uU26rcoB
j37MYOiT+YFnwm9lun2wYMLjos+g6GSC4hSV0gZtizy/6mwgCT9HyStoajkYJXQh
HkVC1wVTRJQX3xieogJaFdmkkypOMUDNJ5HPpYd4EBgFqYRIbYouDUWmrp87k1wH
JMnvbdT/RVMOBb5QV5CpLM3Mxtjngh21OwWKmcaWSpfTk2dd9wTeZc4KwqMlSTMC
XJQSHhGGJP02NS/EFVhoJJ8/o19cItOq5/nDecWsoT9d5hyrRekE6sNPcMXnz1a0
2DKW5qiqzHo+6ZG9+BQH4STz3imRqhzNbqPQBFxUazHog2qVXnQiItwx+GsgjSNg
j5HfjFhfto0VyKRLx1hw0BdPXzLwfOLv2Jf/rm50dkW18SzHym2qI/phU0a8rRt7
ZdOuLrhsW/u9P2oOhOT4ps2TcsLlXlw1awvtU4p5w1FCSxuarRgdeYNNo/y5zwRk
FRdjMEjP9czGWeP2FlIUUJZIUu5xmSJG/cwSbKGOKlejWLRfPioL/c2pcOxUDz/H
irXQdbu6ATNQeJU57JMllaGC/cSaG4eE/WNnSrIdlIn0kOZ09kstry1hsecaALHN
CDpfyp8RlS81bEjG6nI9da9VJlwqyLGnuWURN2Uc5cf5i1cBdY4NO5ZW+TN/UitA
WCLPCQRoh2Z5W9AapbdsuYh2bz+fr1hmAXEJImH9zQow3wF6087/r1ayQnhUMSqg
wM0u5PXYpp2cQuUWFK1nMjCQqrfUTU+yXr+yfFbzo4BuBSv7RX45fcpE7foLVOyJ
H+Sr+wTw10vl/XP34WtE5mz+6/YqyJDxM9A/XLMgs9gCTrJXCi2VDBJcInIwUaua
9jWObhPeQp56O9O4lspLvdY2RIGhIj9rtQuMBf6JM2bp2n6mJNjKghbpP6NAScfS
wTFvfVPyDc03fgXUBXDbhbEZIKmh3wRcw1l1/wumxlLRCU2aD3o10GUtsUbqjOMJ
MlcIQX5WW0WFgffrGP0AJPwXTkBcv0ouwnQGl/zfzTJAqy96jUCObbkxzUqWmN1p
9Bi60zlBGm0iJ/6N7uG1BKuyqAbpsMgMnZQ5/aRNpQsG3xMnGe3lVMVHK2JZs3Ih
/JkNCPud2oYE5P+ZuiCFFngbcVR8jz4ANL1xif24+zBlSw99GgZR7/yaUUheFfIo
9Eybc/kpZcvoSjfu82Zmf1l3a5z2Jui7wQT3l5uRlyiudy6LceXn2sRK80/Zf6dT
Okh/uKkKZTuU68zFHOuzcRpl8aQ/y5HUk2aStO1nS/aW0vJJ0W9wOehawHUyvIll
+Jg7UIfRkiAPKl+ELw9gETmDqlSELWFEkqC51H8+RxWjUxr7YOxyUbTh4tN+VGHo
csTT1wbfVPilaTu5GM35NdKgqAol85TXWgwF+Bz+bQOXX6iWax3YvZ6V7DulOUHY
E12afOA0LpvBp4Pogf4HSTnGwAeoHg4VPLIFJd0ejXztfaKlDyxDm6apuYfRXHRR
OlNn9RMaPVJkC+LITnyCr7jXg2iVs4xxfznvbWzL2isr24xfUsxUt2SIURrTWDAv
7Q97uCWk0VMGP+EM6BzYLbbz1bxvAjW192OyfFr50s4HCf1PD4hHgaHJg1+qH3LO
QFaEy763RxWbZJ0ulV1UCHaKtG05qapol9oU3u+RSlXxRiwBfxesgFK7P76m4kZh
IolPl2ujQe2Y24wmOQhWuzqoA58URj8zIdqvGFtVFmh7wPp/Ihh2kb94hOElzrxt
MmcuIj5NdoPYYSmTdh9+yzijcmc/vtpA0GmsrvP72zvyO5JLkKPkHRmIbXLlDPg/
o5/c1DvDh80VyWcVd2OEAL394ZebGQCymc4dGzIh/VxjSLpnET+dRVZA72k4P4Uj
QPYnC9JYNCaxsKrpNHYCzAaiyuLBxLcBusGxennlI7zcqy+iZDCT4WtBgSCt5daL
1ntLIIqI9mr3wB+GMuMD3deJyZE0jYG1CyGEEy7PpXXTLI6VqwApC0SwEtU4e3Yg
aCwpJHjwla9a0cr8QjvjaIAT9AQis6yIYaRftlt0/uNjV2wRa1MpX8DEyYWiXZTn
+WFNeiAJf+Io350NWeM+WS1TjOrszgrNL2pEEsvnSY/cDTaBGTHr911wziCvfiol
/Hg7/iR7zNQLkHKZDulf4Jgp3NoncwDycDEaeH01V/3dPjsaUL9tBaRWWsvn6QGa
WDcSMM6jANfIzvENDP9QtK5/khb4dS5SZesLwXPzPUQjm8t9gn5dKNmyqLLJ+WT7
64HsrhXnNcYDpMJl/qGI0NLf9rsuFnmsjwa2pGbm154tqNO7ddStqYhZDs6VgYgr
ynQ+osr5p9USpjs9/ZtRlMrDA3JuLP4DPZyU/yecJdVIqKpq0XeLOmCFnXF5800S
CMS04C0RFYlcH9SwYYdFAYRO+F961lJS11lQm3k5Nev5ChIPke0S2rfKCAFIS3K+
kqEZ6vr9pxNUZO/1FVhS5aL0fcsVCjjNhPUYkmNV3qPlI0+9elqQy1pOGAGdCfrV
BBIw40zmW87om2m9Q3FhJTs/GQR5obGDXmkTHoGX1c1TKQSaliXDvGBMzv268OGa
TjZ+UB/nrJ7/jta0lBRnDaMy8B4aMtdisy8NlsjiBIq7sD8GJu2ZJoUYJPx1m6EI
GXClwPXjxnk4N1ILQ680FnGVLnFnQQ5MBjiRrTl6PdTlUSCflmByM+WgDyBVjl0f
n08ZjWLIqKN2g0eJVxJSxC5DmlemcDUahN6C6hJ6kGGbMDW+Bq4CNLmQaBOT5iAM
1ckWOnqvNVkoUwvgYe+rwqXqRzNex4QZWjAgm3eP0aUa0QJqmyhVOwB4igkWBZ9p
/T1hUsD5klF+WOZAZd0n05nhPbc0m/Yve3okY0baCfmMg3YuxTBWOmDIQQCJOwQZ
qqReN9OiPt9P+DubhTIh7Hg/+L7JaMaeiM4E7V8H30FJ+PSVXqzJfZmHW6M3PHTJ
sQzsR/CBujwefO8agLunqQkGFQfzqEndWFoN/sPuwUi9mAH/4TKh5Adl7VA1IuG8
XRL6juDSK0t3WmlkyOqcUOFQ9EFr+uX3lCk36JPi7DKKhf5kGCb7c5pqYWdrmEBl
Uv2lAGd+oOdtXtajtLTTqbWfZXGtomlNa5dEjs6CePhViQ0+gFGUqmlTTwDzDnWS
ps9C9ueSC3NRWOOfwQLveO/AsaGSb85xt6dfodnngdXuSu3rWPMYwioOW+056z9u
0AIlQDq82wVu2EnbT3qowwWNp3NITNqZXdv2OGLzXEJRo2dF97OUWnuT2/tvGdmV
eeOb5LGQexnLuP7KYAtC8un9T4KczkWpb3FTQjGLWgQEHMlE+PTM1dq5TBghPQgY
TuPCensC0lpHQwALOTSf6Y0LKubdX40Y58cjOWGLwYV5jSFjTcF/8mj2NJvJwPRZ
4dEVC6gFRMpbPgsANG3vuVKCKWXJ7Un/VttBtJ7UoHXNKBIwNZgHuBIee4kNkxr+
F3mFeFwTigo0bD9xaNmSaJDJ+dXYncn9ZDb9BK/7JWoEMZe3PTAEy1f9bk/kiQ9M
wVD1J0hTqF0dCgs3xjlmJ1nmKP5f9ZiFsw+ZhKvmct8u2q1uotaRVSqJEmQXVWUN
G7L0rA1fLW0XMeyktLECMeU1Tio2RX5EGUigTzpIFYjls1+APaO3KQ65ds/oO6rb
0J2zz8fuS1s06AQdbgyugc1YmNy2L0BeHjW7OrDx4ixWn3AIaOfOIVOwGtwLm7+x
O6YmKncwaifR2N8tLvTu83pKwPsjgcLaeKYiR+2gSbk7I/ese8qMXZG0I8BVC4AH
ZwRb8Hf3h+HVZejK6xrhyApd9palR9yHxjgsMtQ/WkI9shMlRVxi6k2Ct6jW6jvr
OWE0l26a22BGxH3xzelF19uggjuUszWyKt/M3IyLXuM0Xa3lpHFTwuyoqHXnEDYa
QaOv3rEcsTMsuZNXzmg1ACXpWxRRB/G7f4zTBQ+Yq2l1fn2vjYtVN6c68lAcLe9Y
1xJlRZgD9Ebdhc16s0EpMw1SIJzvt/RGlzP0/0VrXJUoiaCuKWzC9LxfLeqlD7aX
QLgbFD8R/cHlSp6auah1hdTYFZqvhUqQTUW643JOvnnbYO9Mk0FyBZHebGeFnLqr
Zx9Vt8V5ym5LRzTihm3Nttc2z/jcZnBKmRuIzfKflpqfHEfsdcdI90hy1Zp03Q+s
4TQSp8gl9WX2YFmmDSq747nDlBQuQZMmJeMrtiGp0OnjnSJ1Qij2v98gYhWq3SFM
GBgTMUeqAyvhLF+kux4L6KV7eh1hwPRAYg6bkdXGd3rqLS6y4hLN1LF7h7HmHkWs
ckTDmrb+HCLXrWpBtyX+WQqqfgkFdg6ZUWrKPIRVb4qgyBPQ+1k65iRlV4Bldwvz
T7r6yIb31K8GR8xQBjoElJa7oQf9FtpRpSzvfh4CPJrTq363sUhh3dH88qzZSEFj
/a5UrbZ837/BbFHn8SrGpkPcudqrudpZu3yw4P/Etmq0lMG432RkQO4QdWkDBe+t
Akx+HUBIFGvcMZkazxVnh1bAEjtQjLwj7H9dTOMKEJSmNapo7P/IC9fLYPyF6RUu
MiM2FN8hSkByeu4FLs4SIUh/MxQo0v72mTSeIRnB5ljXM8i+kGLw7qKUNsIio2ha
z/TuyTdh7wdSS/G7Ug8UVWjHG55aKffDGjpX9dOgltWncIzU5tLlQ32a1rFrhEGW
4LP3gqXIRjMw82uJyHTrSxbcpSuHK3f8AmCcBaBWMn8QSr0fTmkZGySfW2V7qvbq
GSZE+4YPREXRDLb8waVWNDhheCTUV0BdDIRYxzgmYa2NHP5pWpOkFoZ0h66FMKJI
Q9oJqxXK57VTHuBqIK5ExP2iUYy1PWWpdvJmFmSmrVkF+LhDyAeevBv+JtceR2o6
6WMPfckEPEHVIMbnyaT4C9D+D00Kpr0UN/DmvZTCIAabyM2mHI1Pja3rfF16qCau
6xL7D+PDZsuReTLv1nbUf4SBUsG3wgPKylu/btlS/XEqaifRZgRwTbi5vpyICOFH
Mmw7/zohyrLMx1+N3gQ+L0RNHdL7lnIqNPAqC5XMwvtV7Dp2qT2L+HyVydoEjny9
omI8qdOkvB5deWtbhT14Fhb8AcL58WO0llwqpU5r8lZ7BijRKh0CKUa6l3BRaML6
4whhbCQA6JAOHkiTF9y+LkiCZUlH6I9RfOr3Os5OSdYHJSvPaEbPhKH6tu9F+Lhv
lyBKB+Kj+cijSmUiWt2Ahjoj9wAfpqlODxcsTEhoG0v9rgZfQ4pNP8IL/4yZhSRb
lUTIZNfU/BcFicg/XH/+QYVjdVYAj9Ph9peyGFBPCZ0O1tDYbw5wTtfbx8+iB7bu
wFZC9+FIL6RbwecwxMfQZi6YDDnz7PxRFAy49Lkhg/5ARDXqGD+0PfMQlNl/jNes
ONXCEF9anFUEsRgHryoQM15DUe4O1zbaJviXxQnF8wiN3FSQegDRSb3Gb3TvjDSa
KJzfsphPLR48SoUZxsaOzTBjOSY5f58nxJOITDB+14DP1jHi6ekF8OAt2JvhyBTl
eAubKOvURcNL4JBhwNeoyKypg1A03Ik8rUIm04YAg/iUGXEIqI8JRzk5x4xWvYdk
f/CM/EW4GHYnob/IF8qLdZVhgbf564z85gldTuVKyAexGeLqaqO1rl1d6QxKjQHd
oc3LuXVPzOzl5ni7rJvARv2CBU5VrbnTGnORITOM6m76L4Lu+ekbLiK/6eW0Yd5k
7U04qtJdCmp+lJJXTCFVBhfaaEXB2chldHPrOAzvfUSjbeThqWgWDbEuwr31qHSn
DYewTVNTrIHIW0L0VVbXAajFzpGJIfFvnHrvdqSs+gbRFiCRGPnLgKjr8J1p4Fd8
V//nILIiTnyMGQdw8WeZMMDsBMQEScY04KaECqhB6S7Kp+t9bkzzEDc1A3tDMGAt
mvRa1eA0xoZ09v+AguSuKZ3Pws9vqdMSuRAOYiqk1jpibeZEYAzn2MYGzP0Pdw59
+W5bxmJjXPXi4buVMfk7PklP8ldABvcxC4z1ilBGTZ3V0yFKI1Lch8GLJsQu/Slv
6K3EWnRelOuKPMFtrlQLbEiNBBqVGt0F0Ks8aD6rJz74RAM29bjlyQWlQ79Uz9dU
yl0/74I69O7YOy8xAtbKNPUmrnJSAXlgGFHDUkwbS9Kk6uCv/34RUJuTBE14w1S9
Tt4O6rRxoB8jOqSwTp1tGm87qw8NpES8gbk74e30S5FDdg1/sdp2Y5a4yUu9Y2cM
U99oW56J1HX+KtSxzouzbiS2gpD+guDfUdqpbwFZEfekz1ydesQnLcjLHOmMcjRn
8Urb+ekeTQORCJltJm4bLRp2wkg4HOljJuXiBr7RuZ+nmqsYnIEKevW04YV9PwrW
Aoar47HRSiiNT80dzDCxHC8kMPpDAg/81CnBW93qnOVNp6pw33XUjrmIV6CV7GKQ
JAvWNZ2z+W0O2MmEG8MbsXLDG03Lx+EbVMtiLQO9DMd/sySJW9eJk0y7H+z+MlrU
HLnAZauoVyLIN68ubpFWELmbhyHLF5/nRhGTvl/LBDqg2y/YntL1SllHmjOGDUYc
jgLhy8IFamS6EhMBaOp3AwFlwerrBoEmbjkMcAVR7zjVmn/XDSfBBsBItvHTR2kT
lY6LDIWBa/aiojPANw4ucEA0jscHn9NvCguWKrS07l8Vey0lXn3eUUZ0EO3Ltqp5
BKGxn55qetnZEsL2WakraEYwyL/zG+7btNj5g1oSfcExN/8Xnr8txMps0AMYoMZZ
8Zb9cugiTO25Acor5g5Q3CUTVYiqCZiQfY+8l8XeFTf5hTS4Er4IKUCW82UXWuYt
3MQB8i3CuPAhB4exiZI+iiico3Qk6aEtqS/6DHq9kAdYQ1qj6RdGtG4nFIOUC80y
mLt1B5BHaIPtWJcmtVH9Dsd50xeFug3BkGTV1ktXueq/i5/FNpKa+yB/LD3lfkJB
dGi1uy90lpprahwZRkkfv5kxJvK9BZk8QnI4piEM15Zu63D9D25+VILwU2oXckt1
bXPcUbK7oyTcqx05Qk4jFvfaBNriaPTAJFmfWBBXIC5JkcnAq4/Bgw5bQJDk28ld
u9xBU+2nJP7bcipjV8athQ0vy2YJAiJy4rUBi1YgIxMy0XREGyW5RbG/dBMsbHHh
+/af+1yo/jdiOI/XuXD5nwgnvzCL5nItOJIEGEe4CEXBsSWK1IHP6qJezUSnZVl7
nHNQoyY/vcvtMDQj5Rr7OmNaLQA8CnCajuNaquPGx2eXOSYRu/fI5lQE/cdXPmFe
grsx0wMEW+5lDmnFsS8qb+fvz91HiY/RcNJn6EeKvZq6vrELlCDrqeOcZrEPfT8J
7luhv0tljFxRsq3scnXUjcUqjT1zvnkgM14uSz1LnwtrI+5Yq6a5rOD9616KZSWG
EwRptFQeGr3g6sJTRl2jydk4klQc+iTzRR7OewvWK8zdkDMu0/i0b5iXZjFYCKrw
EHyja2AwpuT/n9gTRZDq5jQzLjReVlsTpfPudYHWd0TfOxxO4aijrnXw1b7zlpn6
aHbjNVctbB6ku1kBcsc0Wm2UNJLioPhAiguPw4vILOjupxoLnPuPN1fYAlB6lMK2
Po96VQAf5elMZ0mhvbULyPM7Au4yyDAmzmOic1GONA7sEP6mYbXJ1Jat4KFw1FRV
/+sxQ9F+u78N4cTB2Ua5kAWK/gDlEN9gtf1rMdBefXmIQAkKKpKowporIVaTsAC/
AnerjE6cCHC7J1fc6Lwu35/dHE8CGbKHU9wwpFacaNugjFcSlkaSdkc/PSBBjvA8
LA7EmoZ9KfT2RM3jbbOCfyDCrjytwSL53UWA3leUGmxueWkwtpmY7Dh2Qxt+eX67
aBQH8ENn/Es6aYVnNennwBWXxH8/owxjJapmHewUCsMfcLwB0sFzv3q6G17RGK07
69wlhCcrSZ8B4PsKmahaPyQtDhIyLdldXw8HIBMFoHzVImNSFXOhQsI59ccHJc6d
1VEU8BBvUW/TjHvUmIf8xKHfi5RR0yj5Rs5p82vZ+htgVx1Mjt+hb6M5E7cSzl08
c9SFI+AatpB3kcq+zRfcSpT3nmysrhnaGfpGI52V6XYDTT3f75QtU71LpKJxEAoP
G3/Skrz4RODgTh4CtxcNSlC6JjE1SfpvTK5jA+wI1SZUSG3IFCSd3yEx/oI/bhtv
Z4Cgy72XAEyJf08fOH/khjd4AvOPZI1d6DWaLDZ2vTNiZzS9BWJuyjerPHvBhOnK
xQR3tzQWqlQjIncqqYAoXXkEb4NGqT9EDobOjj0jEWEfnx8bugdq5Nd3fN2bEIn0
nRlrIhpaQu9j9TkUJmq+isrAQwHrvgiSdvdlJCfkZ7D1wJRZtHeUXyEg7+0rZNkF
QPPRvnCf0B+Z5Qv4Q1VMgwafTic1R/DKEBe4KjmnNAmAXa5x/GSE3AUXppDamXrK
YKZKpxnmtxpkGLr7/2T4vxreAmwTCdIEKgpIGJBMijfQzs8vK/bsV59P5sBHv44h
JMmVJwh0PHOb6D1kv0i5CihTxYBSqhVsYCXh4uogjU2OeOignfB8CaBIA7OQJVcG
MI+b+tdAVcmGxBfuoYtFy7l3Idec8quTkypeoTGH5AUpxI0YKimfdZ+cYK5DmNrk
fYai6wPv5fhOXyk12cERcxMKVkkcYsSL88yc6QTrbIQQAZzxWmPU8Hnpw8K94Kh2
yPli+a6DFBHwYvnj2pJMvwfkKuWWRD+xNuFO5jrM8JS89RgpVaqgBfEILbmRxQoA
eQWvm+EthyioibV6ArR1nAqE4yLrTBcCceTV3NdJ/YNkVTh1WK/dDHFOGAqtccGW
A/AG5Sc8EH6r5lP6cryPq8nXo9oKvP9uWmEsnYlbE0Gi52aFtuEHDs4i20NQr9L4
+3Gmd/MzENwyBGyFxOZ0RTky1ykuZN7jmkjBfRa/AzpETdvFtaJO3wit8WLKqtfZ
vyvqlOyyyItfd9rV5+W/pUqsgxvCnNTMYDjlP/SLPrl/JzYyOkORQEccKw0Qe7tQ
f5Yo8d7jdnWr+YB+yxyA0YwcGw7GEXUFJ4hakB9P9VPO6aHj+3LTsM9qzwa9MZYc
i22hKPnVrynuH+Ez7ky4angnFGhHV2DlykZjBew8ALqFqGp9/1i/qO+cU8Rc61W7
1s33Ebu5QOqJFkNeCUaLRhQk4xI4Nhscw/neLuVYzWp9VnFySaz1v6LlEs86OhDX
esl+caNRdXCXu6WrV7wb3rvetN0wVnqAisecnm0RcbJvEFXjq9/6uL4PvN93aWQY
jtMfyW+52OzVm4DaYo+k+sM4ZXfhpNP7B7SN2sYm2Gtd/ZWFGSmSNmf2X4HWorXd
g9C4TXvWmNLsh5CtB3SNopbYiZfxC9Bt8fmTbAC/l8VewCM53SMJIbfTsYd6fWYP
shWXZEhPI1woyKSeIdxQc65zW5QhLvqQdWTRAbk8U8Z6NE0L0Sw6hXuiIs91cxCQ
2gi4fH5Uq3YiKshrPWL+KhTYkEKN9ReQqHMQYalfA5T2JwQz4dFzhprZc33qBAPQ
hIUyuIxjfEPIBdkfiV5dFRn7cXTFgET2EZgJRZAvR5rHrWIpHl/LQVdJmku830Ry
/esM+nhyaXpE5w/BiReo43HfDqjJKFxlZO2TPYI9CVRLss0HiIttuGnCCJwC+swJ
3j+Q9dMlz3tAjUIH1LTmT+xbVYHNkicwtPcERRFpL/W6PR9nT45BKogb1PKU6hCr
MHKhNgKP1J9XdfTjaqyXLKqgcZznPVXFVUH+uq4RBbup0xQmOjBT9eLz3KWPAb7q
swwbAXr+k9FeRFi2ctKkJX3ictO7Y8g4zPN6pZCv3CfFfrQe6wpLFgkAInRefsE4
6EtfJouSEYCbVkO5vc4avc8hkI/UHpbqtj8ku2HNciOHHjGxi9lWzYU3k9yzf1JG
usS+6gzL9tWZUIDYAvOn4lkbbOGTsFJEav0WEmBWOpVLh5nIgDY3Qs2j2Y9ABixg
Ckk3vH33GbJrfy/mEjP0PgUmGBgEMr7fTM1B2PotLBB8Brfx6u1n5uRyB21Pa8bd
vMDesvdK06pKh2Z2nc45/DMve5Z2F3JfRjV/AqO522oY8ifZrJJ0WN0Ef0c/T4EN
71oVV1yXjmrt1cV/T1hX69lTmuU2P58hdM2l0CnK4EYkLz49uTg0t8HSXuAHu47m
jQ09zGhvQduhjk7YnFQOnH9jIgm3r772hrvV34MTl3kbVdWED9LhrEXYk4JNVsE9
CrQkE05jVLT4edIXqU7xwilhlNdyCjT+YqcvWgO+UjbNbKxYxrNtMjDEXHMswPTr
ZzW8RvA+PEXUokyY6ONLxuWcYhmLRuMfS9ghKPemZhsOG+CZZV29TgolGs1yCdii
jBIfqlK0sfUBdNAh6/LnkheEnTNeDjWvyN7knMTsBHgpvRfQFALca1RpWbmTAgjP
Si0cqojhuZsp2+wi8r1HFezx5zLvSiDJMSqST9eLXY8qoo4+H+6HEJLS1bKN/dQm
6CfyduswVMgHqrp/Z5pwvW+mKoJ8wY5k2lJSLYXxLMReQa3S95NhOFQPaInJsFDT
ZqgeS/aQKe9fonxKSLo6VzTNq8/U9kelJe6aa3VriPpt4kRJAvL9EGtN0x/pD+8+
W1bB0jsRqWB7B+bFZuIbQrMaV6RbbX4dDbel9DyY4U2IdlwcjsI16aUAEJTT/Eo0
IBilhy5TRtmJXmd+sTyAOBmLy01R6xy1RaT5S0PVrPeEucx1kFWIE0UKi6I5dRvC
F6GSejZU0D6E4wCvYy08kMNl4juH/1bRCsG77B6JG29wTwnga46HrcEb2v5C0l/P
YRuQtGbR2Y6St1r68vLDGvnNlDwnyK0QzYXIveiji2AfWzQO/w2LxA/T1PAFV8PS
XcmmWlJi3i1IXA3kdXRzR2E82Sm9UxfzHC9rdB+GOoYaYGnGB5DWwVjr7xhI4d5I
p5jtfeZdfbMxfZDSNIEsEonLMXxi61hAtPJyka/XnClc4xLkJLj8RhfqzsYCF2by
amVWRMLTMPhHzDVQ6u5ZS2Nkr/Nv2e2n03GGTHW36YU+A06FVxxaoJfaeia/H8JO
KUT9Lh1wMhyB2IP5+BMZ/5m2uJAYgQ0D3wzKS/YXUPWn5Hhazc65YvtO0mq6C9+H
/fIwnDIoWoFCYvonb3rhrcrOQTVi1KkSiIjLbqiFZv5mYirhexNIpZNfrR0A25Xq
mRimWW177LHsbf/lnxpPmzjKH2LxxBbXdogC5WQUaLve3ddZYNFkc8+mkr1qxlKo
BFkg7vLqK4A/7J4cCm9lsBvotYJZW2ceD34nPFcAZ43+VipiCxZtZhS6gQek6n+H
/ZAnxiR0OLqX/Tl2hhHIY/LZq4jOMTScbldxJN5ZJnDDGrYk9qmUukCvTqvqdAmS
Mdo45b+ixdQREpVzyLawRJVSPLFMQrQnjNRsn1vVoLXdRXwbzBvvAGsx4wMg41Bb
RSk3Hhd/E/pQaJvcrrIAUbv6W2gYHInRNH77yoCTOsSAEhLaAXGfZcrHaJf9usOW
FvG81FE88Cqwhq9eNYcxasPnIEs6zgNLc+8Ii8/URo9tRQJiFws9mZ+mGzb3MdnS
5WpmGY9FE6RSgbV12oxJT7SrIde7vXX+47XKTyqHX8t8T+8nMW0qK5vRpgdHzoKk
0znphBXkorGBtYskH4FI6yHYXJg681VkIRvNURuYjvTuW1zE2yLbaSkJuOKoBTdj
j9uub7huqvgHvLv2vbCEAA0tlHp/A/rhRgdXYolzWNU2wo3+1g8yiFbYuCjHaJKu
Sz1OnyOwMZ17WLJJgrEgo2eOHuPTytUbwHd+dKwCyhdTWYihbwwuG7G2qGemhCHP
Zjl5V/2XxLLrJb3kGWN9R6m5cFqtJ/trinmjfH4fe1UT62MUpZLHTtV1nPBKiiYf
W/g933U0Cusf9Z1wN1Vmjxqi++AZcAyLsULUpDiUW3RLCedy0k341zQveyRCKO/d
OrEEnmBwtdaW9PFHRgS93YQJ8RpBWY7eTtHqMbRSHPozhci+0gPzm2zLwB+KtQYY
ac1e3Vb3sod57qxNQPXW/Ks903TmRP10FBT3SGx3m4h7km/FqRj0IhYLUDiQzReq
2G5Wry90OhTr+x0nXLpg7V6uTSIUR+bwbcIw7MnUFnf/bdct4PGbSufuUs1J/QUM
gYirqXGpLv5xvic7zVp8FfxdpeW7o2yF2G7rtZ9kSE59Sh711RqbeAR4gmVjvmIR
Gm8xeVZ8qqQPGvdf5KT2TrWXXU3HTHMsmw6mFX1GYotFjwhUX2NvhcHpbbFVz+j5
5qEyHIP1NQCgTEr3ceQ+FPbEJ0K3FZgoaNKFZBr5ItfTlXT/hrdJRuV2nyOWFi+u
rlCWSJx6f0eNpmHItzHrDZq+4Q3WdBbSkuHp7xU/sWrQ4tIScpgZpiIdGgCvL9UB
l6IEDUHYLcOKB6yeTqlM4t8iRpHRy/VlUxZomfTdlmq8BZdZ2hho2atBlvi85zib
iX8Z32EbKIYgeQ71PQA8l+1BRzAh7jMLE+jlpCBkVO8zs6t6VlB0Wd8j07gRFw/i
P2nM1DGd7t1sVj8M0GDLIu+3taiGVzq9AlKL0IuPdxKJQFqnrVqUrKq3055LHPDG
WwXpcwCgP9WvDmaxWQXjLeKtJChEY7lQgMRemQu/YvWkUTWaBsOu3QDykmOH03uN
65pta6tuWxrNDkk20dYHzmDHiRpE9WF/PuGBoVhwzPtnUQLFT9Y47DYnW86MVO0O
6RvBoVabwsusLUgWpp8gQKMfy4Az+784LbiKh0KFFXp9SP2EUPURdNykiD/K/Hn3
nBFJyv8nIi+vqZouuHMJDmlLT0F4isQShors5yVYZ+g81Tkq84fHHDoKJqOvH9vr
CKCC+R7RzTriLY5mvSNYItTgyoWzOdaogpRgU6uK7nHBAkdkQj0w+nbF/5u5YgMM
MyLmyBwzQkPOuN2lx2MjLM1efx7TNeoF+BLREBFqmLi3bGi2dkxAApSOvVgdIbER
mqpQUaRpufBJc+d9tRG0a3O6eoP0M0eR9OQWekHQAj4s6EmL8ohmH35UO21bZVrb
vZ3j6LzvLe5/fKIBT9aJoKGIymqNEfZkNnRfws2sSAEvWPI/26lvhFZ4WZgzuhnO
aVnkyDs9penZRorObYiCJibbu0pvEzHfoFuFsCUfv4JSND0WmvsvzmVbFFu2XyTj
pPg4uEhLtFhbwQKyFywL/8aUvP4k7ziGdzUlVwQk2CeOCgPPJvJUXDaq6M3UCGJT
3aLyKvaQfh7BdNCCwmHN0FWLEfTI4/DgZkgVFSQqLaIWjqRG9C6pj3J6PyPjRLdS
dr9swEFj7KnSWJMP83WUH2RG9qz/MSbeQejYC3dKwxMFUOg74Us/Uq7frwEVQoS2
usZE6UY7ug++T/oOFuO+Tqhp6izeBBT6WEObBIAcr8zsNanAayLiNuTCKYSGy2mg
dgacraN/qoORQyartUHYL6pCoDg14nIPMU2uwYb2dCmqKq/XnWylHhoOnntsscJP
fK4iEIm/fNQ1mWgjAX6I7QreSW8dDDHcWcQ9jEtw9xeXSOsL0Z1/Osg80n48V/BR
9lDneRTJjk+Imgt/4ycll1s9kus+gVUoWVZD54j1kNFjM1TpKExLXxkafVxYg8uT
IiPp4/Y9Pp5z5BQMqd/YDA7uzJhPIpixrEwKj+8gA8DERiLQ4h4jufGxslk3VlqP
bn0pqqVNLDGj7DF8oQkcPgOabZnw/q8ORJeb4omq7naUAVvQfzM1O7KbRBkBn0l+
riyA0tNLplJkPKQx7MqakDvmnQnbCiQZfi2UhVQc5OJTRshfp4zy3U+XTOj1FtTm
uRnsQpHBJg3uZ2WRb8GSqDKi4EfQXWqWYIcNSe1ZyKD5Koc8dW76oTVmpXTjxsEJ
hKQLl34KhDe0CxZhfU9j+HnKtlEWG9OOnP3OwewU69Dcn3vOGAjldnxARBkqpgDU
Qk+fQqQp0itCrmXpuEjig4/RjfqsSG2XRPkxZeaQsMvDNwzalY0nuPJIMhbHBaqf
iA4WJw+HjyCtwVp5dMp9Hj02m5n21tL7G1LZaTTuEkjfsdCBCm5VyK/rdFwtWgfG
xhvrRb+bonPn+wp6i5NrRM45EazfLxxLEiQk3fIkD55Ej6R3orDwRvGWBtwHpa8a
gteEuIeXpId+vDrcOdOxGpXabJIyvLtL3y3HRqSue8Ed/+RaNShHao1Ajy3t2G4X
GHhve5ctUhTtwGu6wbHDeuXU7DGVIxY92Uz1PEo2cs1E5BQLkwWYwgDjmv0sy6vK
2LQxbzbqcDhimqOolVaTbVTf4Y8oHa+8b5hU586WPE8K/fIfSktvqyS6sDJ0Suti
txLIEfGBrQIaQv5Cp59blif2H5UK++wd0pBqnyNNDdScRjmZU1HYI3CG/66bQAZb
PkDDZQcuiFqnBjnoEXIJ9Aj3L3yd/yX4iQYwd1jNyS85KT0ySlwrKc0/vmBldyiX
0R5tBOwFdvyZedOUtgAuZlbN4viNgCupzU/nh+8Hvgq3vhbB4Ii2OOnts2LUGHRF
aGVr4vdDnVwaApHYMf0v+GBU3170Eby9Gc0+Af1bIJooZa8xxJNaeo2fhB9rkGot
L9h5JrJN3eFk3/UHQxE9A+J2ioN6vhLfpyNt+j2TvtKhwHKtJmxvL84HwKuoke7I
WVMJRolEpXIO5Ug5eJ7ieLKtxMFEOH+jqUqkCx2Kq/F6gHJ56ARYGiya6SpxrxB6
/e772/NSRZNvgnJWVBoPieBgJdKIGgUf3BmkafAnmVTiP8rw8AEgWIGCgIDr+trT
kNUHPw9Qi1gdi/hGIg/JTUfkbCSOd2Hpm8MArJA82FVGkPTV1zp/E2UFv3ZrWY+/
vmE6sR/TXS9NKMLBwB7E+z7RABGhm6g+l+6bSBBpAUcUVbiACzxk43pqeC+hPpK/
F2D1KmXsm+mccz+stjn5M0chE7Hoj0xNeHgBfoaoe3aGK8vDgwByGS7wKJdzA/sA
MI59Lco948MPxyLcRBRmJHdGmcyi+pcCN40ttnhvyFquZVkplQI0qxJy8XFg5DEr
p95cGPWleJ/2/4Y5o0Mus6n0PvQ2bTNfCltGYYlYb10bMnxBoOU7dAEj/OjCbXw8
dmS+P7HhEg1SnanvnPWqeB2FLCoT1EJK/gCOg7viz5bb5IuYcUClXn9+llJp0sse
b7j3r2awMPE8LbMgkkUYHjVJC89VxldAyBEdo0dOCwNToQOq40t0R61kLQnSkDpZ
Gf6E6tayQwWxgCKToY1Dbb0cPGicu/FGXWtPJ4nog1AydIflwm2cfH2GUZ/5WzX9
UKLsyMvhJrm9r2OOiR7yCUh9ovbY9yT91x8Y5GIISAjTJPGqVxt7i+97YWvXgZog
xx+HAGLCaSi8e2hMh+tr4mdCoBNxrbf5pWBQ7wTrP6LEOPuslOu5j2RJ6A8B5Zkk
zTmUyvhTOSNC57AIxD9gSpyclexm3hTUNlfzbZ4XiA8FwewQt1CWgDEB+tQVGuqv
5eeRfb1ccqXkbJzvUYFdX14LnUmgzRmMoahucG7UVoeTDgu6Wd1QAH70en13CDXm
1dm8AjfdNumHu0Fu5d/jYZ9hfD67TVzm2AWaQyE71IqOskuZ3JX+MyEY9mKHqZeb
5FDDQQ/cYysYV8EZoBmaYLPM/pW90OOxFkE7qvm3MFIE5rsOvTWPDq3SO3sAOjiu
8Mq5YYdp5tq3+gcK1ay81FZo6LzhtDQiWUgBuhYf7AHIy7sj+56syZvo02glX2HG
1yQ68QbVjlK5rRowyB0Yb3Bc/q8/Rl6oNWBREKTHD4XTWavUKM4Ryu65BFJqVLYx
YNhC7ApyIE0Q5lrhwZJrq/S4ao2G3ySI0/9039FdcJRIcFJlwe/vk5WggYxRi/cW
Aqt4iEBQtAB5yFh3qESJIXiUM5MHUQf86U+pMgfa8lfQ/OlVKBCuP23MUEMMfgL4
km80yE5YurRfu25aQkMM5Ffgw3aTJ8ZHv+9WSDAES2l8YJe82QyXvJSTMLpOKnll
tQBXwmCUza98Ye8SsOe/2Yj/5+SeLlSP9cU5In+I7i2ahlqrZMdb0gjRbyespt4r
T9HAxZfvaQa9kMOuI6Zcb33Zq1uTtup58IRehTIGH/jgv2EkbQLmn8tRGqaE2L1c
kgpfZqY/Cj5RMujUbFY4q0TLCD2DRbR68xsaIttytdgUpPBtLkBPXeMoG+H6RB9c
POW8QmQePCa61DgNVwLmzndvHu3Au3O4rf7cClHRuAPeqsfDlA/iylFYNuS6TqaN
ufLQziOCtjnB29YzI+9Gi1M3TlSXkiyLpLjjeai026Y3nOU/++uhCrN4Fvl0c42a
DCAQW8VRwsMR5z/lNZYNNAi6m9fWnHFhaY6mJrBi6M/Z3JX3+McLwlqTs99V9VhF
IHKMyHlBwbb6l8rVWN3iszEqTaY6MInR1JG9e6J1r6fDIh+RbpgepXAh8v4s2bIf
PTA0inlt3b50VmG/yQuUkQz6Rs6gFCqGPJDnSWAP1iWaUmbM3YbkxCtNlE0zEsXA
BPIFp7acyYu8z+ZyW+6Bqeo4RT33qAu1toHOplOr0TLBfknpNtrNsMdGn6hSGi75
f3Mcerr/761E8jt3jShwlZDmxmG2xyJiGed6zq8KZbpnEYKFZh7DsP9vtZYLXN+3
RNI5Y9gockHzdcJGA4hGzDykC9nmY4RLV8VFfm3qYcvWD4nrQaQ5tqzSFVdKndgH
HKCmY6K1x9OJ7+jNuM07FizDRR17UhcMGnMlHBhWeiEk5k71CxvKVOMNt1yYhr9P
gmAhKro6trxJpv714jSPu5I7b3smFFxWNvxFGxtO+OuERUY9xzuNHSayjT9lSBtV
r1Gisu2D1vZaMbJ/lit5uGyrcWrq9EtbzL7mgoi4okejZTgYLWhwSfDDE6xklLza
99PprcTP/2X/B8gdD4CxioIiuqt9GfGIXZNuwS7rJ/BkqvQOiW848Q6ndk90vD0p
+B6JbTO/yWg5X3+CFp/oVkvdL+OX8AXJ/hJx7pDWXGPnKwPtJvciQdC+wN2uHG9s
ZiRY8oreIgs4PwOOF/K9qHx/mKrldGk2oHZDacC7sQbNVD1KpoIHZCQrP49BX3Um
32HGeq9MGHPRSKQsSrWVuwzAk4ZARDNRRNO+DQftp5n7Pxe/U8WFSDWYLbbE0i0i
hnL4MM09I8LYrzdzo0NQAevYiX2gBk81qEOQ9u1zEowWFfuRXgz1uotwwQj3uU7y
TRdZ3eMTOpPWdtTYADgW+eEotQfaFW0zwrt6ChjoJ078kUK86OqJr2IE4ZXk5aRV
7+fpeBogWYNljTSkj/LsWNV3MfphO8GKxIVpmKZInmzWEZlnkeGZUVQ9oCuX2nBo
muOKuKVuXuBRBb2UDA47V2R8dIS5UAyxT3mNQfNvc7HrYfqkrDKKpidGGclYRMRG
HO/VVLq6M1W07uJOeGEWT4OnT63CuOfo+ueeqGCVkKpZYOv8fyrcRqL2ZTH3kfDN
pKfYF7ut+qKXdx61uEU9ilL1XvTdrShmr4JH1zZ3HqSzjvGzz8ZrCN2WTkKiXK6o
VjfIk4bgeEIf4BrjX7kIH2q/E5FY4nQOQrRr9OePmW8zi0HcZvHQBoK9e6OINZ4r
778pYAzUPaBUhm0OGW7kf5dpkYPgrQOzhqhW/Mrz/++45DzvxSs1u//24nT80WLj
io2BAh0cd9Ar5JhKvSuR9j0EqrKf7g5oEYShTzUhKfU7W2eNLedctD+/z7/Loa0t
JNFmWgN5bivY8gRp5X+95K/pPZ3Lz0Ti11YdMAcBMO7Sve+au5w4FBd5wSvExd3g
ZEHkl1x7hVMh0ZjE/Jnliau1sXqL+YIHl7ivpAz2BcXDxPPnHHmuhG1twPxptI3W
DMw3DT3JmTcuXZ5qgF1HwRXu60mN/otn8NgpfcAbr8TAsxG9okUZXszH8B9X6Hir
/RYqUdzVB2dF+dqkD4jDoAKAePWYryCBNs/ffnor7Kio93NgSVjAiTaIyPX7kWC9
hvVAWp1rCuYBIGuM6SHIZq1gUkfpaiwVEkGuaBIY+yXIv5oYD3gFtU+e397GIvoh
lllPX/9fnywXA6UYnJUyG+hyfJVECJUaXDlC85JtTGYC7erp8alnqAi+3w5XtMwX
4OqvwB3Xjajzrb8d28B6+6+TI6qOQG2t6uyTCYxqbYd5Ci66wH28yj/P5+owMt2Z
9tRkLsr3dYW7DqFNwwjTUvo5dmSDE/pPwpNCU/ELxmHXC2F8t1sfJKItZjjfkXmb
4zl3EVZKvx9mmT2UFnms11EgbQwrBC3IRzGWbT0NXAetrTv4N0iP96ywZf4W1yyF
V5eM+sw6VA26Wr648c5l/Uxag8fQQTtwNnge+7gQk751ZigSTYi7C5O4TZ3lwa6N
0gb7SNOscgbMJmLZwBJ7DX1zOQrcmh+OL2p+ze/b/3pWbY2Ala3FP5+YuKVrzm0n
FGFj1yeMbIda3GXVetfGxSaDEKkaDw6bgjGFVz61YTxiw6y0HTQESsHHnBQl2f2q
mf2rrTq29CjaU8OaKubVKYiNbaFWwKcYy0pU8FYxC+hn9xRk73jnC4s4OJMqFgvC
hrHedk4biBm8CBl3vXqjteVdWP0HSTuoDKoYcmNzSGSBsfsl2IXu3TON1ZZmrF1K
4y3TelyPTHQ0HlCKeIh25+bZoujoPsSV2rc5BnpJR5ISyy6F9QzjYb3xEMMGALnx
mSIpflaN6F30Gar1o2rRBmVTzxHHlq2pMLsKC6jCoW7/pYh/7qXA1NYy8Mq2UijB
I7ulXcw9xq8eC7rh3pdj19Z9VqX+DDhjhm+1+DcHteuN1mWDrOg+5Wk74+jN7YWW
zHPFw86da+URrfVMMVrIy7KrweIMvVP61PvK+GcUxuSUiC3EhGFioJKg/E0B5Pnw
FpfvUNkwEYU7MIDbLw3OBlvF6JK6rRwImnGWIBsA1QAp4R9ZpHisaEK/g0VRLiDk
z9OJmDc6Rt38UbOjQl5d6PXS4rfxquhyVKB5OBBOLGJdNRry4lQiGyr/lIzHovFu
MoDdebMeMlvWoIf27GhaEh8xkky/sVB09kbg8RR67rd/aGza4/lS5+w56blPg3mV
b61yD4rRA0y+JADNf2k/Qv1dxAkz0lDFsPRh1GfuPXQpJJpXP/RYw+WgiEpdS6dE
6ug8eB2/QIwUDZIEstKGW4VhdeWeW42wrULgcz73UMn23Rp3Lyy7UDRGPTMarE1U
CUisVJ95BoJ1JR4Sd0vBIPyVPPuQKi70dYj3poAq0EaSfS4t606fbmotnCAYM4Az
hd9fOuLVhLGNv4lDY9yAMlPo/ZPL1ntuRJp1nqPDCp1z312PmCdziKAFODdYZaO9
jQcxS8qyzroXi3ItF9t7xWUG2ZVMUHoInCdHZekBc6MaWbc1gj4VIFEzBg5vuy+s
2OcSLPeSmCJtTNzhFlNpm1Vdjm6E5D20fBS49TEfVQZnyMrNpdUFo+7VzMdhPj0+
uh1ArdL6UqUw21f/axOF9dQIFcvQmLakxhyXjZt8iaAPf+A2xh3l8FAPuH4GSzGn
1HkqcP7/KHhOyjNZwPS04RcgvQTKi0y55tANi9OtF2WAlPw36MRMHaRRC9O7GJJq
xnl9W9k8lMq7GvKxv28/CPJ3+nP9STJLeaKgBf0Jgai2IhFwm9RxayiR1dFVP03D
wNegXfGJj3QrEhSkwvPLozSBU5erkEtjFjN1cEeQabj4RdofxsbWHSN/jaXxgD9E
J7BEPGTyKUyDQw5gebq6QjljDavDNO1XSuu7pSLo9dRCM1h56E21O+avCUhCoydx
WkiUy6/kExpKHfHvlh3tpYbT0+eikBIf3mZWTSbYbtp5mWfgO3mi7TWeao1I4Fyo
Afr6uIAvuonq/kLYi3LG9tXvw/joEtrv7aV72yZx3o8ED9IyyI2fjXAwANauXNkQ
iXXMIiIp2UiuGebix4vNEvWd5lQfyDNTLfSBIdtDo6d11iZeTMOa8NGwu8qw5zYv
/qzsxyBTPxWVRD2ymTMcLQxZ2kJwCnHe98BlCefVHbhYeBrF4OfOY5GXFa+M6TLK
uzEp7Gj7IWIwUa/c6rCET3Aw9C36DPRtFkkjoSMxAX/0szr0s9bghNRjmj79ab5J
Z5xJkqOPbsi4XlSNLROa0GIqZGdYtO5HBsMY6/Okk88XGEGeAIjTbydjD4FMYh5V
mnUcrBHigvqtLkwmJdeldwvRZjZlmTtd2qHWCIM0nrX6RZDws8Y07CQMq403zLuQ
aC3jHe1jnPP3IVHXsWih4EWIYWiCFVqVBDQtF9Wo34ecQcJG7/EJJLHRYjelJHqF
rckeDdvKsMhA+cb7RjqRrzr2++iVzSDqPZMvc993kZg5n5aq5tnQ68sDoSxYOyG6
dYI0+Xv8+Bvos2RYD+x495fMuN4YqVIGBL7IpXbQebBnmCbOzlWiyictXCp+qbLN
0nOroVZGZgV1rlNki43rpaf6xf+suXwi/0iANGAXVRdV4SGtnoQL21uQcw3p8TNX
8EJXloG8f98SUULeNUBScFzWe7OEGntbOP+oqFORDuBofTCuaA7ywqdnvvg3bj3Y
tzzUFRI5JCc3j59d48uBoOKbbRqXnIRSwr3YLGvLUn0L/L7tXECIuzTFQXbPPLvV
MsosvOpm2nUpgC3VogH2kVSnsLzSPtdE+Nq6wKgVzeCtrRuL1Z5vAuBO1k1/2Jt8
rqRgjGfXlz6C1yqU05jpCdW16zhUukDx8QsKwi3tvtWn5QtdEb/nvMY2tsNC0KY3
zkzzydVaN1scB+BHrr5epKQdFXTZMpPvYqsRLbR81rebONoJfGezDaBwUsN1PTg4
ZEGD3YmdGrQsB3O/DSm9X4TzaGOWoRHQ2Ybo5d9WAS0rw+wFoyXW1305Ln20CpS+
8W4r4sR2ektJz76MaLP01o4UJXa90h8sEft4PmZGnXcxWpXWAkFun6pvufZZMqLH
MjMTDH4isxGj8wgkg5x1I2oyJMo056nKToje+/l+ZNwlr3qLkjh/+p99xy7MTiP8
EQPtCvdohCx4A0Ahg7n9VPe+rH+8sIy5ZXd4AbDo8WQzW26qkRwE+kH7uE6eDkEp
Uw4de9jgcwGN8V2TRhn5gj3rOcg9r6Jg/gnDYv3I3TxREEeidf3aZRezAV+nGr5/
FiyR6xAS0VcLIjNkCHH/D5Egl/qX9k7KvXCNRWnxO2DzH0+a9ME2HkF5tJ/IF9YJ
QcFiLZW5cum16zcBwNGaXIdEBZroVzmXhENh+NI7ZjIGX1FpoSGVU3e+yw/VQAyl
98OhT8R4OPbFa7OGbXBWU0tRdQu4z0IIcYEq/Vf0E4BLJPkegf4NSxdbU7XkBbSK
F3bialB5IceAUc9a7hx4OLx503430yXTD+VlVVT2yTO/Tqf0/S5ntCnG6phbrReU
hWr6ya6fiXOVcYLzfcG+SmmLlcL2LJJzO4llXc1+QHR4RK7AlUkb4hhdscDKJC+G
KzeXteWaHLMzvNSelRACg9ZnWv7Dp2nGj56yR68OvZxaS5e6l69MY0QiNIfdqEUR
UnplHQRiy/azU+rLAAA/yNAJX098ebcP9WZqUngy4USS26fQWUtaa7q9X/ugZogN
N3qEGAUxiNgO+wfI5obw0MkXyIG4oM7nXbDkLXWpM2NJA6hP16lx3mIoMMbPxWUr
l4fULqdB0Zdd5Zq+bnT+RDdCyJO9dxOBqdbxf7KDsat9IQP1UTHOsDlBRkrvuFCE
p8IOJ4QKTFFLlTq1sMdv1IcWUQBN7YpWCVpw+1twKqITY27CpQGFSmLobo5zrAPc
WHvJ6TmZSY6BmHn93cLEjNt0zgAE5VtPpFFUEg2TDttdh0k8bCwYeG6L7SyunYnJ
a9eOnuBkBJF6N7fziNx2Sx4nK0j3U8cIriPt26T0wNA43h2WYYWi6JuF7pD6Z3hu
mD0kTHlbUVL4pJmLZCpFqxcFUlFBjNHuEu+Tc36buEO66WwNq5CygJXlRotoxks/
haM9iCOjLZVkPwY/vkk2DY+BsgfV4B2ThjvAxLUb/pCkqii8DZNY0eY1uBX+V9ki
S6L+XAnjEcnGZ9ZjBHuPSFv94IMKVvf5+eJDsCp7bFyegnciOADRL3zK6ht9jELB
BJ0ArCO0ajF3nXni+SsacYyxcCS8qKttaLgEGlYkiyN07q6o8Xhmt9j4W50z2owp
D7kOZebRPT6u2afTc6pkQ1vA0wAybZG0g5549H0Ses6IyRlJqPMFx/orVYYoPyZo
UJvwVGSDkj/d2vc/4+udGueYT0eH+QUBJRazBzLJHMrMaOx5UMoqRLX9A8EJ4bSx
1Db3O5aWxod1AnW6jtzViulb6JFHn/akzFM2wkm3uksclPmk+DH3u/YVrMfuHlN5
DrBmHaLrBI+ZKWS1BjqCOKcA5yNuq/coF8/djZvM5TvJXtjoN8Mqtj9pM+diLnfO
XyoNTc/BfqJjxQ7C5PI/29wjN9a8MDlFQc2Ee4Dc8CbYEi1CI4K/OeP/67UCGDii
W73zGgSY/MJBzYqUAuYV9GKsSgU4yLyVsZFjEEnwo/esaBlk7iIwtYR0INvO7dSg
EnK5dmADlAvbRJd0bMsb8pyX7t5nM7z16y4dAV5bP9R7CTDI5Nfrlt9NN+UhypP0
97vmKqpjedz/DJj9HfX0HoshHp+G+WOVMPPDAQso1vs6oU3+N1u8aVwvHHf47Vwe
aqBiu3ULpTqCQFZrW/GtM0/Qgj/sSzbdiab0UGRDhzcQqbZYXiThN8oWt+p4jRhP
X144oXaWb4YEpEHzPYWNX2Bg1sXnt8yAYN4W2Srv1pHUHzbMBc3BqKL/AS2A0mw5
vXYqOS5fLpwCVr6ZKoR/EjYsbOb1ddSf7ZV/4eLtTf7AIk1QWdT+1Iy9d4HTTfIZ
x8h04vX/K1ZZS1s6/QAnkNEqM2BqgLtGB9b7WgjFZfTq1ZS4btm3NbiidsiR2Xfw
hWiqBxDjhVVamz8Lh/VE+tRXudHAcDjep88ZyQ1r4uMFH11p8Kb0OxPsMetCjw3S
LPtSVY8rjhg+8nBajBzsnLFIErtGSLXyW0T6x2ry00E=

`pragma protect end_protected
