// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
BnHFFgDbRfUcKKHhQW2GFDHsUH+jjcrLIgpqmNpxba3w0mHVGC615PAL+xNn+0L+
M/uxl6YGT4TagEJ9YpBHmFkQpchn9lcweoip0Rr76nclkiOu+meMIQAQKZgcP+Ac
UMU1+YtoaiptN9Ss/YX2VT/tM/iwBcOdBS3OsQ/ZiG8R96lveechvQ==
//pragma protect end_key_block
//pragma protect digest_block
8ynDzWMnKrmm+xcM3cnPUXycO1c=
//pragma protect end_digest_block
//pragma protect data_block
bObSxbziGkJmzTxyjCrHARl0R1zl2gpgBng+hOj/ge26Zx+Z/QWIpd2u+fxDjziP
T1Nu9qzddW6VsnfJ+NQgio6Fvpe0CyzSCkTWzZvrrIj0ehIBkHzfbOC45Be1afS9
B6A+md0SbZBSz6C8pB1/ER+nXliA1qeyvKLENZsOa1vm8EcQmH33ZUxs7hUjrX0E
/XeIXfcdWek5hBF403777bnJW+gEaTdnQlwLYavcbdaSlGLNp7Tfypb7OjtOZ9OJ
dK1Vf1eIm5NHOtLm1bf1kDVGBPdz9B7nhRYRy8otMRQhUTGDAjQiP7tG84IDEtE6
Uxvxje2RrLTQuK3wKJjInuDVxdWwU05Ph+dh334s9eY9Wix9BzxzlGr1qfbjD9rl
2CXCEp1hoQgJuueJXTalZbMSX3KqKy6bTD44nFYFpF/3G4B24PDodHKVQ/Nl33cc
VMEW1g4O5vcw5gpWlAC55S5QNPhhrmgarGvtqSqu79prpqnw2m9jgc+u3j34GqSJ
RN5hgWvD0RxXqr3c3DSs6hwPuWgRtu5L0U2ZybVTHoPZ7Qyv/MCOMuPdP0g5XW/9
oFYRt5n0KtXbSkQUf3UibulGQQ1q5Hhuop9/x/2r/DVmhpiGeLq2Jz5HBd+fX/rn
CtCkFHSyNdxSPsqRk0LVcH4YIevv55U3cCbbqhtLlaNi3xvsZJrYTwmH2F7f7Ugu
GEHsVa8ECW0tlVm56D2vh7Q3zNIPXS/AJ66whvr1uP41pDuQ3H7AgHKgnPgRtlti
45o451RsLhGz969XN8xeaOWuOLOJOH5CnnWeHCbrpQdQoVjpcE/YmJhsXJVRyHc+
K4QKatHc0DPaia2gvyQ7KDtR8VVzTkAor2vv/JESSMLGxrcUjS3QnQf8K6sm4mum
sEELpZP8s0WBd4smTdJbSdqtmMs1rDdDbDHbouDXyEx2pkviYoeBnYmgsar9zL+W
9ZfhGJHDYdEepEymv29NF/L9M+U7CwfnH5bcLxU4uo+Z0ZMsafmiQlgAwyThFNyM
+sG76riXBEE4r6TI2j7DEKXTTBOdC36qOC8Oydn4ehfAKw3cR+70XVpBqDnHxmWv
Pq4F1fwf5lVssCYUbmUyQK4hCYR7g5S5BGyF9K6ac8TJpQFtbjcf1XlMJzBDYIHs
FgG5fUklmoj7TeOTAxQE4yLuXSimMNSEDxcefjgbqLY1l32SGqpv0sxfga+0lmW0
akfJhBur8TmzbbOomT8f7ndWfBhock3os/+D/ikuzPCYjYW91WRc3aAz9J5WbUsb
nC1CtAKQukAS1EKpQjKldmgHb1WpJEVdfm9eCFUaEdJqAZ/by1JbUWQWK2amnnRY
MF/x2Hx83N5mfZMHwEFAzie9KCzByKmBgej60rcmz67isqDysWT0qT2UJbW2Qd9y
yJY/qVJFQnFSX4HkSCvU+pInrtoROeoF+l84Fl1dLS25tTaMEfGiQxzpYt/rWRwi
FXw2CNMAlmNj40qkRCV2NjDASF89z5zLGjLNW1kIuDmjVv1vVzquZLQprBebA1uB
CNl96I+A3jhXQQDkAuHrHulDhUMk6Gdt117OaQfn8Tfl1u6t3Nj/GC/XES3EQtor
iFcLFBXWaVv6HPl3XoXpU+FM/Mu/IL7/sju2kZ0ZApV25laIl2N/KF7mWCWbOk+l
rInWhZzOei1YCCHdVhd00PLJx8ahFu0EsH/DLKrtNJpnb5njdZ559VaN+N3qAv7C
sSgmX9/DpmBrJSIgmQ6sMXyMA/HWSFgDLMkCO53GMjlIR4QIQTrpELE5q7M071Qv
UaFLLDncG0OVW0r4dXL7J6Aoii+Ki9NF1fpL1I9zy7KyHX0Na1gQMuiIxAPFQolg
71qgXBMAi67Ps0LxlFbnmV79D0IYECZLLsM4zVoHFJN0Ofu7A8zYpr/tHNF8tsEe
JieKfWHNpQa8tbCa5sBGhVj1yjFR9loOaev4JPvXMBWF21ptNv+HhPnu9K1jfOB+
e8MnNaa6KTImX5Xtf6ZfJPlMS/cKrhwXjl1uqERZjlokV9hvxHXwUYpbB9fy8JI9
qI2PzXHAlBCD0RTbwFSeS+g4zvxCXgO6JwDEA8L+aNZQwjRq6IbCoubAQjG3atQD
ER/GyH59TLDJJTwyWkwQsWTI98M5kxp4K22u811g4oDUURnGPNJ3DvQ3SM0CB4MD
OjZ4JFMA6stTPPNF6ds7e4Mu3xZ7j8cHKFxD2K/RtKaSOX1ERNrrkfmPzZUPNbSP
plwQpG1OxBTs4gNLI/YJG2MV5wkOuR0fcYH8FgCrcxPyYMrP7ULbvcjq6KBXhCVU
KFhcBrH5Cmu9KHlSITBXnVtjRqFMYhrz7sVzkCxsqrVREK7OzUzE8fG1fpq+B86r
deaXG0marEpL3b3GywCJgesKUlbW4xDKSX5YZmbxzWuZINGFaql/hp89dWApkwwU
nYA6sDK1yypE3j+Aval/82BkTBEdaCqNzCi4nMZ6JGIQMroV2e7J6Lo87qQVIZGe
JrgkoHLqwTdIkp1kJhOtZrgITm7yVFhSzbj1GIWLlmVloUclBfaZs8rACLtHhq0k
PQ3QsNPlkjWUiIWmZQZ/qxG/IUi5lKCnC1IQI49srCXM0Qy+DVp5XAlpvWRITQJX
BNT0DGAGcbon/6TC1yLBxCYXA8vAEEN14vdsig2uEmAeB6+0/8zeAuA+R56D0C11
BWgfstnsRjhrHG+IBVwZJGxYsN92pFjCwUfXgx7ZBA9Q66wI6z9HsNOWWgZ8kH7n
Ug1pP+8HlOeOtC0Idgea52iZSa8urNOD743ngcYwPe5vyFWSoR6cZJJfpZwyMJBN
o8ms5bCBmfyvi8y0D8hDA/SJ70UKb+hSYuCR1Xc7QZuCqCWj+tMt83ngQ4Mja09S
KTmvoxSG3R+ayGLRp6NWjCZlN/IvMPJ7IJ4p4rL6XICPc76NShvBXsZGlt4d92ye
A81QnKmGpgZQoqnwj5LLCw4pg30zlSzCTYV/l42Rf6Q7i8UVT87L8y5Pee1lItfG
2/6sxqiYjVlGZpfo75HQC7xKhy4ZKtQK0ZgWAtaHeMJIrg7ThcipCttEuRkrsPdP
DGDvoF17BA72dWqKuqmNvXbiawkWiRWhgphutkPMlxLoVTNXA4n/fjBdI0cU4G0V
hAOVDnVuIYBuaozCEisCfuW9VuAHR0MRNmecpnClPoFRIdrKOaDvoAWNv1w5hwiG
xOVJi+fJ3ihK0ij0fWU3NxPiEG3loIZ/yn4Eij5uNQifmoPlU9U+/7LKwRO0Do7W
idpVindTme4ce58gyrnf8lkO4bMO9gdecaDVTNxSgVcxWAMB/Prlow+PNmwnhBtk
51oNC/bl+RWySGYyRawnZRqppN4AAvxbhcGPL5cDUBN82yIDtSYChsMazFLSwkTh
E8Ibw05AKfKkSbYbtzqykOHWLLPFWlpAOzDek18bhuWZUKkL5muepOhj/aMkhazB
tWaXtbfpErGo9GsiTuhZ9ru7B7dJYikK/0Bi14DZefjFSoxPUVmi/+u7Zl6/SLew
1bEokyE7MOJbpX+Gah01UCPzvJCIeo6pKFHuk4fKVg2+itDrv01MODMFvIpd7gD8
FafgsRNxqAyBcX2DV22GGxiPAH6ZjAXocu1UseviO4nZFOTlY/szzl8Sq3glcu1z
RiL/1OjWdiX+tsGdKc2j/VrxL4hzI1VKA4/iFf1mJih+QNKiFkYa1jteAwbdAAVQ
AA1FPVFi8TZCer72DlQ0675k4XiO2nzbz3cximu/ompySk3XzBysOPoqUbXCyPV+
0y4HFUqLVDt0Wlih4b3LdjQFACWdke+tOgmc5KG/0liymuLGMAveufcj7yOXmVxi
YCMojMWk1xOZr7Ei5Ogwd9vEjciK3EQWnylWaYSnegMboUdiejIHjC02HYSQ4Zei
cwpzst/3jvhCd7nXO8anTHj6ARRcaDavwu1nXtWPmLbCgXWGLvMCwAMyP5CDFoZ0
1Zn3W7PcPO7zW4Xp9NLGF+eWZbMoB47sOzzHkUzcu5iKPlVPFBQesRcNwDx4Z3GU
zG+922siPEUlY0V7QmIVcekcH1IhU/GTz9SK1S4xgASJZ69aofqs0W12R5fxzD2t
74VX+F6JCoFQksKzrrpqd5qNVuFUAfJlOdJDeJTYtER3S4NrO8wneIr3FwTCgW7k
J/tNRefp3RKZN1R+p8bmm62mb19CQ+gRO/IDKiwyS5hgX0NuT/XreXwV4qjteKyX
UzX/sYEYL/r52hTV7fU6id9/0q2WgGzDLGRr9pghipNFKl0miZabDqaW+9mnb6fS
OZobM4Y3ASWV6Uyo/OzCaJ6/zDIL1ueWO0WZiqG+h8nzg7++6uOL8UTyEkm/8AFx
86yk1g7BCewyPnv5JHIWItb2ikTiZ0zpEhK7fvJ3pdBG+zjov/k5tHpVLG59fdFn
NZbXT9L2FHPRC/JF97EJ1pjS+/G39xEYwETM7YVD45csD/uXYR5nTTyJmBVr7NTo
k5Gdldicl9eK2fWhemiBJPY2Tji8TRBeMHBMGkcFI43LEa/PBpNns7Aly55Ao6uJ
tbmxIOwBZatqAVYCE97mD/H7va1nHAHwQBo9MrodMMDAfp3+C0DQ1y60R1xd28e4
4K8PxbF1MrQDYygo7rozpwJzXRKRWEfq2/y9xsWccYwABN8BKJPihF+hNq8JupZ2
TrPRJjInXP5F5DA3wJzmHLG8iN49UD1gSwOuoSa2sUDU58p/zEhtK1XNfh7anOCe
LCJbAY5gbc3q+NSQVkFVT9vEXkldBMwnTPW513DayFLMWUmK50LRHImY7eZQvuNs
n/b34aJEU+CGvYsvvUHL8GZ+vQufGP3R+U3ob1YqjDLbzElwKZWwvStbKPRJSB2T
I+k1bhwhx4uXuZN7OXRuvOpOjHI+yjFqEC5GJp8XZqXjzX23Pfyhs/838UK8vhMP
syQsTDji8rGn5G278vulZUaqTtLBmxpXu8PdIJcG3l0Uovka0IAtGb/lkY1Suc2M
sYHv2TvpPL8rp9yDqc1TjKBqGyKjvr+/rDRYITTNDsWsOYKOfrZ63J5CDYv0uEhG
/W5h5miAwG98A/XEKS9GVTrIBN/EUpFAgEvfdLkI9zL1Ect+q7hkAmGf/w+q4pba
8DVMhYwGUsrZ9IZ5L/yoWoo0xoHq/iSe946ALksi//Lua6Nx5JP7xaDj1TYvKl7A
lMK+qbLKGkFjhwMqYDas0aQfCMBd4oS8G3rkSiTk6wcCJqKvAuuvHyLzjMSEUvqx
bIneP8HyO8HzcG7Jcf8kDMoEsRFw1glIJCb6MNewEC13jkNx7d22ZnbO3HLUJ7Wk
OoOhUuCZWN9qGgj4/tVtXJ/bL1vaw3Di4/vKZxik4GWRpLJdWXtC6G+mAzrN9igq
BqI/PO8Vhaw8c30ANFUOBFW/x6uNUV57rW3TZc7jBZRXz1B9s98C9K/xsxnwnJ/W
aO8/wSwT5wlD79c8QyO+wi2h6bdk6L9blbiTho0J99uohM+xUUI875dcKrtoyBI4
sNB+7Q3W4DCPvNq121DSZHSHaPm/NkmPzGYeAl+Mu0RoNr1X9+pM3m9DakMe2iwR
g0g7cRDNcABcQXwvo7uT/b3cVPYatgLD7LhyCc1kZgNH+R3BcNiuRoPn3ebrDjuP
hrYkgKmYDhTwYyphnjSIxz8CL7UL9FF2ZPYMfPvriWtzw7K4byVi9dPpBLhSTHMI
auHo4HR/HR9TCcN8m3VNA0c9ltfPLEiXXtZaXMi02kK/ieBECqVHpIWRiBdY0nKu
UjPw2bsrZul32DZsbnq26tnKcD6aRgZXdv/CIU/BFsTrf+o7AOf0MX5p9uue0dAW
UVSfjvXSwY25/wO2/32eni4N6HQOTb9UsNAR3UV3iTjRWbMi7oODHF4RdJt2Fa1g
d2Fl3Rz77u/CSqCKmbIdYw4w0kROHbgrRQ3JObeVxsssUeqKy3KzoPsWJoPaxTP5
3RSwQmmqp+D0B3xBMdIzDFgGHSyx2WjU5PJPYFsLKLnAkV32BNi45HwQB8EAwzep
pDYzUCm7V3XUmq9Elk7Y06MMCINOtipk+o1/XnpfEguhpWyUWY4ujt+UzJkxNi6s
lqtQzrlcvvZqZJs6N3o3u18xjzMN19ua28R9CBP3BUD5Vf8ctVTiwHyvqpEEigTx
T07rtt+jaVmtZjkvBA55sI5kkjDqdnkEEPY9hVR/CVvXRGPDg+MXQZOtNGW4PCpp
SCbd9RLDZz5NhdqLBIwzLvJ246BmAJm2CebE62AyExX3K6ioQJ6SPxajvwGQ+AQK
WAnofDSvUO1FIzdQZA1vSj0Pm/KJ6jkQagtVWTBTtjOV4T8zfpW3dk9p8k8KZkR2
Ve2N+AZ8RA4KsvO2xVrOpXfyUoTynzEZA3VVl9Mz99E6Ywc4O4j8s4Z1cwDaXcfk
uwPdaGM50pnyVI6sTiytRVGJIPhS+A+aJYRvMda0IqoO1iIcGpu8m+g/6K/2MiIr
9CnUdqIaZNExpnDbDC5xrmL1NUvKGceyb7hU2/ZjKl2LFVd9XqRYCHglQUqTmeR2
NvZdD/7hG53gpuj6+NnqAIbc17k7aeOv4+E3YAr/tUsIWo8CiNR361nkSN/K/qZI
Dq4TQoiIk95E4op+ktb5ebcApuukGlS/bIaVXibMIGmWr6CuSpcuGd5sjCvJL9Ti
XLuxXXBnvx28Ht5uvRY6MEo2rX+8NdLf7nfgUv0W4RndGX1vs4xrAU3Cr9KfaAUt
eyaUBvZ+XbeanVhAuCZpphj1ss88MP+j7irXkctjQj5h8YmH+8xueZTyLukfxK9G
s7akvez1r5eAquDLPJlkz2nzF3ggZRASOccH1NjGZY8BQPh4WPJ9DwHsjLxRR8Ap
mvkFcrkA+fKgi3U3vjLaIFUN7171+WrXe8JGFNCqivUHJkTFRf82azKRmVu5q0fD
NqNPIq4MMMZl42dJRIaA4XqpfJVq85HpggrvIWcUOOR4WxEHcpT1bQuHUtdDZqxX
cBdRX7AbljaoD1UzVPVm3Wjo5+46qrQuZ9P7VtoIq3cI6y9B/j2zRi1yNX/fjy4t
MCQbipamDuDFm4dN0Nc1opND5vbKnwonrZT3k4oEApPRS+JNVQ9yR5/lPTJbm1fq
7sZV3FwEPsPCDfvPYqVRIcz7vHLpMbuPpBzSe8D7AmQwFCGdPERHPb3IsYk8nhKO
h3FGD2g/JHAInub0n4APa4uek2l6FlSJhjvL3RDjkxrhz6XPGaUEWktzJ8SP106u
oaq48vCOIgPCvi9HrBnc2YGJqvziHsJ+sWB/i3/PF7CbPt1CxFPK95BQwy/XQH+T
pyIMcy6RWC5pnFzTqA6dCbd7gW7vWtuLvRuyhT8e/kSOGILKS8oju3vXObEk4Zsy
QAM67Kt5Zbb6VHKIk4OhNZzLXAQ3ddTsVqAUMyGRlFQKR2ELSSxTOMOO0uwKbYc8
+ni2gtE3xyikC7JmMIrQcDTXnm9Lsv5epKTGzeF5wIex4A3c/Bp2k9WF+eZu62eg
+QSjvXxAPYLVYBZiDuAvGHSFrvN/DiT3wgKbbcAgCUSNfeTHLa+Phal/nT7v44Yx
RIsOlZRlVpop6is+cMLolKlP9oU4KxcqplLKXYCOT8qX6iUpE8fgtZosbOqo/+pj
PvRDZJEIwHDYqbjcSlrijGEsP/FSzgmqlOYmv37CLqJ0JA9wWyadj61mLatBwBM8
rilWj6oGEkMBcDk8wXxEOlnMyRRliL9tv6+GMLCJiYAuvD2GgDmEhqHUjWJF6wPJ
LoV0nGS4tc+h/m2pvLvaIXKnfAiGngIwS68KDdAWztT+Y8Agl7yt+MtnMgDIG6uc
uUOGHh5pyA17bAi4KUhJJMqftDVGqZwyTD6w9WZXLvPNAVsd7i+uv/lo3LKjJwMo
B8y7H8KNDzUvffs6H+D1Cu1KYSVjNo5/FF/ZXju/Iz45S/ODbxY2j1zo+W6iU2ZC
r53w58tTeyS5YPBCI52bAbtIltUkiVPt3BxJd2zLULWk6HxR3yYgRZijw7nR0akw
bCm6yek9qFaVlGwinqI7WrNdyD5cPNTH35Iq9RikvGlT2jfpjrhsfb80esgDV/Um
Ptm01yggTLt7/VEFk4sf9E6JztwrjUQV7ZfYef1eICH/krOxgaQsyY07WsmqJBUN
WhQq5M5EwaLome5gKWY450cp9DyQ0urIcsoTmytIy7KslJ113du0ERq3HkJaAe/I
CcK+dHev8SeWdTlMgaku+mflSnl3R7DxJGcHBh8iUz3Ex8yiuIeImCUpoxk+ACyM
Wi/w+gCkc7qrVPWY5hSM4fcBNyVChKnsCdO4TPJNVoh0AtWDBOfnpz5poHrspeUL
l0JI5+HzVSeg7Qp+MvMd0KBmXBKBacD5xtgdrqzS9QlSVexvebgWKkugcGs1sd/w
vvLBTVFgL/bWK7XmbyFx5Vt/SvXugTG81hS+fm4b2asir1EhqCgr0xEKvSieQzgE
OCuc5mcKreax7uyZJAK2Syq8i1Fp4EFAhRVl4MYlCa2EgeG8fpyxBIXv8Em/z1+s
qKqpOL3Odfq7CIZTGbGzROMV+5ahwBA0foIwkbZcdMPSLqO6fM56mQOyVfgLQ/dq
L82KMssogvbCxvG/ehbRRQiaknaQ0/F7M8IaLpIxkdEG27qG9Gp0BoDSQX8/uNA9
PUHQN5MLqx1FldgSN4s6+tWp+3Civa9RGf4KE4hFpV9W5kou0L9UsFEeY5bxJYiq
X5eNSkqQbPDAftpB73meWZtGx0eMepYGdpcGxnbVjEIe+dsThbrCNi30UJJjGrQH
l/CFTpJ+o8AJLWOMqZnFafMePnSt2o8Gq5F3IZ61vLyR0Tmb0b3MqEJCWH2HLVAa
L1ijmHAgvkx/zq1vlcrVgunBnXlarxmeozf9Ru03mgABM/LMLWZc6FtBQYYxTQdP
yLHeGcrCaSTgU7e5SUkcJsxIVvj9hVHsOZ92Kpj04oJR5UWNmOj2PE0ouuSuPOXC
AGKeKxSbDwvGUxo2Hx6TC3Shxq5JMJXrUiGdq5OAeIPhe/P63/CxTDx515O2+vQm
KpTLdHb+Exuxso+D88DZYwQRFzsNbBz7FL7f8hANFNiKSPPCuy3js1vmx680+Cw6
XIvjCDjq2tkYRTF8ZNCq42h761+lKBewgNNzeEMlZCRxTgWDCQMJprwMrwdWALJZ
+3oJRIW7JrE//iGgm27hu9HNXlDc1u5UhKPDKdMHr7vQrEyKmbwdg3HGXnHu86u0
nEUUPnsOjKleRY7r3ptS4Y9l4FbdRVVJkceZbbI2Uz+WKLw8QQtIceJyoUIyXPiG
mleo3zaaukbcG6slW/NToQFF5YxhUE1lgIB9FKYYlsdMASoG27LlqfS9jDnoLiah
8XJybbzfHVXugqi9GqHe+lyVbAsTjY2siqnVtk+6PDNLrE/hIlR9wWNReCkwUUqX
by5Zu+pSFwSlBNn5zCr57uwMLkhRZ+iJHLgqoovCB64b0Ct3f4XIE3Oba2SfvzBi
1p/8Diy+ZEPzyQU9/D62LWUOEHr93aJbY+84/Sdku2uscw9K4fzzz2yfc+SJnwE5
hgaxhgv1JDko9XV1I2m2aXBVUdnkeLgtDX5d/ECp2KVseVpzMbIkOmpvYUIUAdza
a24xDh7mT/Ds9K0G5D049WGanf7q08ExiHA3OiJAesRJNxqfwSAfrUA/N8UciAgr
frkA5OnWq/voPOWe5Ov/zaTYRcrJCdQCNIy6kC5cDGuVjbOGOFcbeC25FH0SwnIB
jsmp7BbEKcVfrHKU+HkKBhqD8+ruLktKwl2cXkIXkNmKCeLE1jVuQavmTZ93NZhI
5Eqcoz+2h/xTCNiGEWcLJAZ8CrfV1Mn8TKe//2FtqORarqlMb7gG8Z1gp9krMbX9
/6LPfeQAZbgKi9OcWGfj98bFUPDXhwqmkT7L0NNm7lwuDhD6pmKVHeoESRv3HCrU
JodFs5cnIF3x3zdtRLOOIq0KFuBt3TkDLh6yJ5SSlxbkyL8AS57a8J8mwXP5ltcN
4++nJem6YFbRwSkPu4FIKLkGo+UaTfC87JSic4rk+/zsMc480QOCPk+Afz0/Ibkh
fPrIlDiBSimMZgrxcSid/6oTXVfQQCHsI8NaPhhfyuRVuN84DoefTi14KevqpxK7
NvV5hRzSAznPHEECqKxdXMUP/QRx77BfDDM80W01xjr4f7kcsRsgPozR4C0mYE90
QT6cHqsUSNo2fBMkbCfSHup3/QzfpE3XM7HmSn5kaPf+SNpjfrRy3SFPFWfrm3oF
P0ySS8UzJ67xCA0JI6dTECMU9lNy1qcFd3XK+lxQJGj1NR06ipjFscOe/SQg0a+1
1y3B7QgoPTfJw+wihZVIEc7EgMtmy6KjkRoz6c5I6lMz17QZNng4m9Pvx2iowYKf
oUHKJO0o9RCfzOPqV+kY524sEXkfnAjn5gt43edWiPj2ADBQMsoQBehKNza9b0Et
mSouI0r7aT/uaisK4neo9p4YzUEPz/8AybDz7uP9YhzpJ+7wXS28p8wprGw6Jk9b
hGcIYoG+2fVj4WRB43OU9V5XcMQ416JeVai7i9nz7bCCQZzU8IHCvEVxGR89FRWa
/o7J1kfbxA355njoBHrvg2JQB/fs+BdQ2PDXTQQaOBjol2y8mgFjyMkjfL/7705Y
SgjqU1QwEk1i3HD9mqCSD40KN7LG8f32IDK+T/0FUhdHgs9YKpX6WmU/kIKKKmHj
eHXws45igU7siW4lin6zl0UFTcVboMdBXs+6qhFx+aGYGGxfNAsIHqksDOOVATWx
0M+ZW94DTXbug7OUgkfqxaXyXlELLfOWCSAjhqKceBvxUfxdCpZEdsk/WvfnNv2u
Q+PBguTcefovxOVCyrdQWfFXSNcbtrBqTvZ4yDelBfUktyWYtu/xjdBLvME/vbby
tgUrQ9sBK0MpBCtdxvgvAS9ZWgSM6JrNHhwPHr6/SExR+QprVHUsVwJkXBw4qH8E
pz/vVv6iWRa8eo39/ta4jfRLdmmX+JlM268y4Z0HNObWqo9Gib46RaqoMvoPUKEp
Su9vPHJh7/p6MZxJUl2vBVAPG+5xmDGzAsErVNP2jACf6t0iswbmIPVLS2loQMhj
mjVAK3OgsXTnJlY+pGeZjO8b3/fxVW9AqJZUdIUdfTr4Ki4KZdxzSyqa/W04lMtV
6a8gRw2LBTvq604T5P19cw4vNJSEI8q+iJedzOjJ+g7Zj7q0H00a/4TkVSzMrwxr
nXRUeh2lRoJpSQax32tRgwWk7UC6cxkKWHk6aTDtGIrLAgoXzKxXieVoSZkrZ8MZ
I2Qn3cHJqaXt5HfbyJhqZVjiSsVfK7I0/XK89b2MsvsDTNiPWr4CE73+7RlOv8Ca
snWX6dL1NVpP8/aIlQcGeHRvjr8ajta2Qz2TIpfV4/1uJ/7p1QrkYVWFkp5sRaFG
26o/AT6s1icljavfo0vFthxinVwgwrljVJUDA7wb9hFzrnjEl0slAHp390btsgBu
zHmeFR+rC9+rSee/G7ybXgfr+YoRZXc+mRJMEbUkJSneIu9vUhMGmC6J/Y1H4lXU
Ov9dE+XLmx5Wecw6Xt1hIbIIgjWVoZN1AZXNcGFp9vLWl/aTfpo7X/CKIJwRHTGq
IHwRY8V4h8IxaiAPh6xSHVbf+gvC40iZEBzZolX2zMIcaE6C8O3fRaRhW1VeVnfD

//pragma protect end_data_block
//pragma protect digest_block
XlYiTD5q33yIx5DwsrAHBteZ2ug=
//pragma protect end_digest_block
//pragma protect end_protected
