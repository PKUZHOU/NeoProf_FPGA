`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
LZq3xZdCz+GzhMJPHVk0cl4izobGipIXMW5LQa28RWwAr4AUoh/+YEL4W7fGNzww
m3P+73KVRiWqrFwXoy4mHLxH6GpPJ4H+KhKuiMBRZTFF4KuSZSLdt1S0AGa6v6I4
wAHbd9sVSGD+XMb/XgM+fJxs6fEVpUmc/TvM9yZAToM=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 4128), data_block
j1WaAQ3UWozYmrURANccF3KKQwea9iOeHrW2XN6CQXbvrf1q48sJRVyWMQ8PyahT
whCi1W+5zrpiPnRjZkEu7TQK09iTexO2pqTcabOne4REBl7w3+6yKAeWZSLpwgNv
C/i7KG5BaC72Ufb31KeBIDX9QeeJ7cCj1ADhKONYudhzuPyXf1hrBAaJ5jrP/FPY
SY2u5kUEYV/2JBS81iirRfY6IJ8aMzi5plsDvwmXe5gYRFicsGCRP70jNpLKysnM
/WqSVdsk7UGlHDvXBrHasDgjpjPkKxRWvxB6gW02136fYMbOrzliWx6lMPLkKcot
wQkuB98V4FlAX20FJ6iFMYOT7VUuXVjmHZp19RN3cAwvcjS0krklmwvQnI7gR3wl
0trFTSJDOnP9ORiIfOc3jo9kijRX6o8hG6jZqBDO2eYYKn9wj+yG27Xnyc1xqDnQ
ijfFX5aEuO1gX5aQC3FwQZHfZka/Ieyfb9pGRNnBM+vz18m9K2h/0elqShL+Jei2
9Qwcu1Y3Z33KLlb9FNMi8Plt42G6XM16De5g01aVGGzV63hTIXWWJBbcjVKQF3OZ
Go6WE9tUlA4UpAYiWqQC5kror1rBDHDKK0N9xKVX8wZ7P23kzhNWucK8VjXKd8q/
hITR5J9/Z1ZoBOLZQh+D2MRzqs0B5U1SyXEDOjNpw3jQrb1osJ4tYAOW5RJFtFQS
y2WmWcXZvlPPdLOUquuMSGwdtWOyKDr7kbKckX/rhm+UnKTquAbpZ/mMO8w5yXsH
saCRioKjezL8/wVL2U1u31pxcfd953razdsXJbf7ehN7Isd2SD5HaexDq/syYA+x
g2YW5Rl1d7EiGA95+WSdiMEOJ1ubE541Ol8xErBYrI5KP/bvrHaSLOishYLt9rkb
8uAFpGbuuCbKaFIzi+a6NbR5wNSMVE9f7OcE8AoPBv6M2Jkb6MuQ3DzvO4tLd1ze
bNo51EMa/nNh2XSY1Pcff9YzOV+YJeoXy3rwN8qv0YUwm0oYWZfG/740/LX8v/fu
pv4Dz2Bpgm3bC78RRYAD3r8Mx9bp//09PvDbTLKh5OAgu8oyqjvAPVZKjmGLA0BA
UGjmOfN7OKLtyOGZ9P8TbzENe2gm9v4i2egadlSBU4KZTOZdjJupK1QpI/cy1u+b
LfNhF+mt6fmqw9MJ8y65mKTGr1lwIFHTqHNUWEzlt2jxKs7J5tPqqDTifxpBcAq4
PXZpjtcPxF9kD40MJMcvnjyhSah+2gE4uCIsEU94SB2hoxm+CeF+VSQ9TTHBQga8
adBq8MvB4QQYn6rQDPxG4KJW/2doK8clCoO20bGUaBoAqAcxJn0//Y5evsItxQP2
VstVdP7tBY5m372TdNGMsL9U+WVG0dRVyLMorcqAswaGwKEv8ban/b2aRH5Ic3xk
PvuE1V/jyDhBtgtsRWEstB71el3q7goG3jjg0QIRM/TzxmotAAMxRWEi5BD3OS+Y
xcobqOGa0OiKKTieaeP+12Q6K5aCvQtvx5hdY8IgWSnbo0zjCqIsMAU5it+3nsN1
ytO8GLjw2+iwXfAXfNDn4tfNp2CI5dSo6zHT39sWDNpGDxGwh2EXa+6aVprcTZwz
oW8IYkEmDoVc+8ttQYB7IglmF4cU/6DjPbkBBkkksbluVKPTryf1aY22jR2PeQsV
5ckTth5WrW1FIIY+cYsXNthqjwe3OqdI9aAS+1mCNZB5jMSiW1HSofUYJCtybEms
uDzeUZWaDoy6Ch+MQgHTgTaRlecgPdV0SMww+YF6lQ2w6v2TlSLFlAmF3uRFknuY
75rsAw6CA6orCGV6R3tgzBGikFuT8r3FMjweXZ7g4A3GdlklJTjEtE4x8R8pSipK
/pKgtPGMFLc5Hg570Mzkvh4eYUry0oIPxsT/IntgnVDbn3q+uI84TdDAJtct/Cg0
ML2yzVTGrcNNBWUZyR8kJth1JI/2cEIpgWdhVsVJdHiBp6ZlLi2SjgrXBGpBx3Wn
YKn4ZK97EcAL1zxOtAjXDOZA1zs3MOc583CbwUviZzjlTw72xylGO9iWhSVYIz+d
/Fpx5IDKF2b64PRqkCmG4fXjkkIM7WAmGZe6akq+cbSqGRUexOUjRJ6OH/8QyLO4
raO517McKTuq9Cw6/3W1dH4TC8LmKixPB9eu9x7tQol/iQAberAUQyuhN0uTSO9/
et615NsqXwCBkT6RBVg1z1nKp0R0sebljFueqAGoeYlX3Clk6FuGTJ2oif8BSpYC
C97utPtltknoVL9Q5878Z/QgR5/8iScl14TKcSvc2oCpw+1wxL1vXgSkSLrSMtaf
yc52LRYKKtQKMegjOO5xhccIjuXw+cbrd30QmixLNdBOMKJC30GpSevXG+uoJqAo
PweNKSdid2jBN47iRPa4zgBuMFDRAiuMU7phH/VMSU6hqGC6SA+uu+e5BrofPCTo
M2kcJndSW9EoOkeQKQInozwODNu7+06E3NeFyV5IuiCJdPGXXRBjPu077PSRjnVV
LQtN01z4d97heoxOQvwp9DzR3cRt/5kJlJ+a1oswO1N6YMrl7/8n15Y0Cs8pCbZk
1T1vXKS2aVh6l2LdxiLVkaCImSuHavfINXoLqEOtfrgef8BykfQIrHDLiWUNzWvQ
z76GqNhwepl3LLlgNgMw8mE3W/dNgcqMObl2TqcF713fM204qHtNf8NZ9ZB4Ti+E
tfg8lvx4D30N+Kk+Fe1YCaYR5GORgYycWoHuSRtgKv/ifjMtxh4grm9O0NuWYbLW
kDVbJvCP0iLjnlWk3D5gePfY2BqsgzJg92acSgoKyvPQal9tD1dfDomR/fqEr/Ca
A3HaVjyTI759mEbmHAC0JtWRIRZ8Ehe5IX3pDjax+WBGQy/pK9F7FsRp9EcMD6wN
Vj0ym/bR8S59gNi6Gke81RzfNCE/GzYWehDw9yUFBYhmX2OR+YyQcUy3v2090wE6
HEq6Bd+0VJeFwI/nxB8+abj5g/5NxknMN1AdDKZwpL257Alodq8yAJmxbC5fWM2X
Xt3Xx0M+Uz6/yUDLIKV0EFkaAr6dba/tNGd717KHPW6VrNgMNAPO8Gqt/QqiSAcI
iO63C44e70Af6J8dy54P6kmmJE6tElgWqubHGy+kRI6LuKtdvhw4DIsb9L7SdWHo
rV0jkkTFFev/rn3WTDpSunNRAElYAL5Ur4z6tKKbnlmFZKMxAEMp+3ZJZDyaALCb
3dIlEMcWP3WF4Ol0loNPC5wf/er8OhFZa4TVu3ABcR/nFWW8ImsSGURjJrauf1jg
M1X56W3Gb/v6KDMOJi40wNtX7aepiVOVA+unV0E0RS8/qyYll/v47ywVNVjtgiWq
ryt1jOkxJ0bZlIg4Ak/t5AJDYmBEiyQGb8sa+n7LAWkkdesTAXiL1Vd9LAIDBhCn
7L8L/gxC8bJI/LnqAe2KK2mDa9X/47AQ4o98z1cUsDGT/5dlh/GEjtnlQ73n+uLG
KFtu1YhcDoOkSWolB4kzOD+zdDv/wz/Aee1hVzJ9flI71Ih5Q1xpWRz18yEbtEMs
S2tmiW2ZUxo0rDF0SWFoP4W5FCKjzK1otIa99MpN8VCLyPgaTo9Wlib9LzQrZtDj
vA85GAlNk1yQWsq4rZ9fXfYatIPNSQfVyHIJxJA9Q/5dE2pydeBZ01XApmX8mN9i
AezX4qTn+y52UIQtq5D+CYMVw94UZ7laaxLxhiggouMzsXusZ8CgsXinYFdnzWsU
pqEwJHs7bjL4/Az228aJ8elvcPDJnwofv8OUsnve8L15rMLUynbjn6L1dgGq0P18
JZEi5uYZ6/BSX31B8aY0J+7xz+qmPEN8s+S/1yCyiJScGe3UPkD8ImVYjjlcdOpK
1T+YZlITJ93ZWuYBH0E/M/pDcxTVhxkWkcNEBB/WWQBOXsXVtQxq0hU09AWO7qyk
6GVRh3ZWUYDJQRrMS4IOBFNM3Kj09zj0nAn8rhrUg0q+VI3DV1Gt6aCWaSnoX0k3
5R70rlpWpryzhQRb0j/sUh2GfObtlEeF57aHdWYv39f+0UMvXifMuqBMhBqUOuQ1
fDVeYKGQLvmanrQSU5CGHYhkpcW7bID6Hbg+LmQ7VpsIDhlP4FEFUDmAyM3LMPFP
DOWXd/FebH6LWrFz+GDv+X5JpXbhytYqXhGOPZF2ZXmLjuXWuhXYebcsFUKm6hTF
lM7Dyv+vybS8y33qSn4VYnuawKlvDikB0ilPt/aE/9QbWa98Dpmw19+ks0Ae+QD6
iAw5ixVUfvm3Ir3HJe5pHszCGsWw3T8jH6GKkLYOGqebkvj6rmm6Ga9R2IVpHsBF
lz+qijyxJ/72X0tNm9sGIt14lfSBZI7N0D3ZhuXMMJl34mZmSGw4aQrYZV7h8WpK
bqj49MFKQyxhFUAWD12cx5WlMTYmWjQa+ZTb8ZVx4dROe17AZoW6M7YKIM1AIgdZ
EBtNxjzqZtJopzjwrbnEo7N7hwXIfk5gajQq9tsHkghAfg1vOiTvaj+Nujk4U9px
BIdZ61EA0hFJniCeouJdwTP6gAU8hLdLI2t/oN5vnCl0LpT0DE1jE8oRi5qZpM7h
xl8/TB7yFGCSY9y5yX+p5ICYADOneEMwEf4qQVkACCHsFkUsFsxcGKEgYOIoFmsW
Vyfe+kYUpZwWVvFp/VoPO5d7kS9KnmVrHCLOTou1N6MBck8BRBgeRhKuPmgbHCPj
Y4UyAeYJPZEL+IrzPgAKn0m/tNufVGy7de2YRQZDmOuXUr1JPE5K4YB11WD2ogrd
GCG9PziWfodSes8MuSREuHIUAN7tXabajitz0/WBzzUT2KEo1FpDtMbpnQPAAk68
BlNdt7actlEO+6W5vSwwS6ROPyyufatruA2x/+V7nW5HqrQBJN50gdARoI4lVcc2
fSf9bABrxO3m06F6fwTw8GPyohEp1YEwSG3+ma2AktIu+sBNU9tfRLHyU//x/qPz
L8EYyAc7NRyzstGltRWP+n+yHrmJt4LTWWuity5a9s7AH+Bjoj1hmZWm9RuMbuXx
LO9HslrQ60DFCA330kiEmoihysPla5hxoG6rBdAGt1f1dfsQdGXNJpaRtLMzLQ6c
4iHFM6RdlwW6pGAhW0ndFN3Mz+yLzNkY6lnBjCIHz2tQISNM1Zkc8bciZtRuycfa
Rh3omanJUFM+d5j/1b/TdnhJcCxsjEQeBlEVXpOBXS2bxGIHuNbDMF/LeHuR9SlP
agC0WGlkG9BZksQxPg80Y5tHbpRxWXRRUD2lzm9ZgQMhXKsxd9eAoIdy2fYUqNLJ
+B9kJXKcwJd9Ilv1/rYoQ9jFLc1BJJhNNkLkEo61V4i/4hUiTul4gGLuEbo9ECSq
Kl8pDAvbOQnL3lp5QSQMhLbDTbXK1qruFwivpv+NZFQ8zx/V9yNJd7f9U9nKUiwO
l+XEUF4d73F+SB7Xre/6CulyDgfuRiyHUWp5cM8G+K2Lg0WZpHJREgYnfQz1EGPZ
YRWH7A0OgSEK7nTYRorWoXRECVWUQ4QVqSkBvd4pE6k55xoTVHELYHJU5djRTPBC
`pragma protect end_protected
