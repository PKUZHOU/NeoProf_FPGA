// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
/wgLzZLc+06hSdtecRqkTpgKB1XFDDvNG+CP+CeaiADbWmlzTLBl26pC6MCzivUc
kt5FhC/3w4XMCcBMOxpdNznNF4tP/VYhq8g3JFFtweBbjfTZQNbWMo7TvnVzUmjv
RrQpCGWgOIiqwEhZzvH9iL9mflVU+i8Hdoyg1caHsTcN6bQwUjHAmw==
//pragma protect end_key_block
//pragma protect digest_block
SanphUyQ9PQmFj0l3HVJjetlcuU=
//pragma protect end_digest_block
//pragma protect data_block
zNk9ICZLHETbY5RA2ciu3QPJ4CORWHj99ubMMW4c2DgGeCa5kKP0RgVXlmLX2fBR
pFUrvdHzr2L062HDKHphkmvQGkpx+MdUI4Uf8qh8SGU9wDD1Pa4IATM3PW+CyEIQ
mFWE0Ns6nr4yn8Avj3bgqMQPhOOu7vHDv43LQAQVHSq6N2O2nkmjctYDEbk5tkht
KvYfkiPIR473nd0YiKql+NG4GEFrvIkwdDP2dMPvS4bEYyFaVt/2kupNiVqkLPKQ
+LUZLBlL3+osNIiSMGi7t9XSFaAd7jkYXtPc9exl/Ba5ZZQHx1soyCx4qPao4/BI
gEjalh5OExL/mQi/MK4Bl8Oukx0f4kvINEted2xzcGIqF7Xm34ppZT7gMYITxAic
ejO44fCQghxH/49iZbgDAj65W61LfZ2tkCdRSLgW/9EIfjcXRzGU9NOlwvbkYh0H
9PUz+wq6C74ApLBh3U56uLRNv4nNyYFTOED6adgfUhEmVQJkAwJ7Okxgh9PuRe/e
vFkRkxe1SKq9UJWHopErhb5hWx0v6BqUg5XictM0mjPofafVGyxrENBckZa9NFxq
CQvnhyFyqIQGKJJnNIU9pPWYelC5uDiz1sDTcalg33oQCCT8VbHO002TT+4wWKfr
H9S71YKt8CqYxyfqeM1gcg4e4KsWiGILl4Xv3a/B9gkk2FP7exDloBySmNePNuaQ
qAS+r4dg2ve+CitbJXBvDbieqPMiU7ORVyEfVhL2jvhioILCQ8EIW+9Qufk/tjp3
cCyaz1M0qlFMCeSXzg4h8bdBznTtvnhfbLXbtDM6i1ITkEJ7wOxNc6rrRYOt2fwn
/KBB9fePRwXP7umaCF6/xl5a/wUpsov5QuzixOamPk0TJ1JJDl6HqU8oucEdD8Gi
2se9OFG9LXupVTYJkb4deV06ZUNtp4HT3w4p2+W8jLNfjjRYiox3Sg3qRcnZZ8HH
Q9c4Yc75ttzOgljpTTq4bT9tkV/FyHJOlKWLbFsxlxhSojOQhPejR21r/n3Jifty
4td9TEH6Sh+0Kxqp2Cjs1MdAVRTGm3IS+cMEvgtSQ8GUenUj6GhFTIJpWBy4O6dB
4I6bzGFtH+fnjqqz8/4WsDnAjuZV6H5zBruB9PjcVv5rVmZ1aIqOn70HoHd/56h1
JZeHzdqBCLg+yw8aMKB4cWvkU5AezgVnXQImv5qNHOdmnxR4L1hZXa459nJ9FVF3
8oQw6i1CB1iNeY6zyg+aj5eD9AwcMVI7///qHcIhd+2jq1pOMmLtb0l7MjIYzEvR
W1l3NPAdihE9mMmodGkv7VIpbc83CB8AyZAIfuoBM0M5lRcKVs57BOQn9MWqZuVk
48BlsS/IzF37cYYQdwiYHIunLYXOMxnYBrBJGA3R6sUANsfKIHfYd70npjV7mSwD
LoMBH9f/tpj1gB6kkPd8MN09gIlrPNPQpSMInSm0yuT7mej55yM/R4hJJWZfeQ/e
PHdugyPtXjpOdZs49iaABMKx78BnH9hI8KTCAVQCNG+tmNe0jWsl8+vH6L6OrevX
EkPK4zaJuGpaCMhiXK5GG5+uYP5cBm5VvvJK2vB54tdpD0e8JDP2jM2knt3rPiXq
V3j/wqdnozEpLyX3eXHk8DDe5vc0oxferm0q5aiBMRvIWNk/4H8Y0BKSY8uwlvic
rrV660egrF4aXt81GZG84dfFahbE2VygqGQqFcVa3G+XXtI0WCHTf09lu2kx1LBI
ktaepaOKrevtpNywwx7kW7bXJXiqO+rYbyvcfrawTDa83pFYlmLl1d15SCyN5Ql7
QtbOFGGZYxiKUKEqVXXFKTE6o/unOlfsvA5lAnrD1wwmiAO9VSWQAURV8jXW/9MD
lnXNAMVqjif96/rEbNtjDSp2P/0RoJMBmuLTmIhDGUWRdmsQjVz7MrlOvchAle0z
vlHmnXAmESpyBrva/cEo4t9mAGmeeaXy1mRglX16I7wtzAAuVDQeNgb2a1UV6QFF
Vy35TQqK3/0r36BaDiZMfkC6IjEpaC9bB5BXhC0XqQrFxAqIwIUtKoqXKbr8yE4b
NPgBKeSiRlgPoJ6gGzNFnBzsMirY8Xn/sfF56J1YkGWPX1Cy4yQq0ajFkisM/Mv9
fr2Zk2sKdEftDDnlcn5v2n3C0TChnACxVNtvVUY8kip7mPIsn1mvmqTX2w9wgXUx
5W/Cw3kFwmSTwNPds6CWnJsm7giiiT2uvDTw1FRESxlV4p5O8aHyK5kvg2/7jgqF
qfUvQKzbRRDKPU0YYEkCcr58bjKIJUXjxVCEHrRRb280p3KpwD5vBNEqUSGRMxd7
9E+gL3D3hZPWmEJBt/+KjTz8dgJ0zGeG/6/13+anYe7Pp30exa6CYSQskEDb7VJn
st5rIHxR/v1s6PE4mMZZO6wAFeUMYtXmPGI2XVHRE/T1GbBdmMzKsIQrsCV13XT7
IpZoLj38tiqwoLxcDiz7VvQwetrdfaUPl5ANj4qdXIp/a7Ewz9NQj9muXeHD9r2d
bJ2lN337vKOQgaTUIPy7mOiDfZlIaD9CeB1HYsKo2/N2qV7YJV+bO7FOfqpaxhc8
azV0uhz0JxJAVq7gpDOqWN7XCiiNeZByIS3BpyMnCnKd4fouPtjVQjMgX31RcFUb
6j8X5Sd+v3HZ/VITg6RvUkX7p8kazgkRGA3VXrAHm47e0EiL+TlD+4wWTHGcZb4p
9UgsCpAGF807ncEiXXdwJ7/Ogdiv29QKjoMSduKusykgcUcuUQh6ECYIe7m5FSgA
+KANPfd3vUlbcqYNDLQQQTudK9T7sC9CGMu/niX2RyMHUqGuJsz7qfIB1bnODm9h
Gtk7Cuo7153766mh/FmfL0K5q49bcLZD6qvLVVemO8eK+BLkS1KpJwXLJUDJh9MS
LHwj2FdEohOQfk+DDD1KeNcFJHJO7TuYNp1NzdxgmI9zDwaHoO89uWpKYWKzmb24
mMaLh4vXJs18F0+/uWigk8YX435xNoTH/Xjp+qU/KT5p7FB9EvBVM7g1p4mS6sMT
yUef+nFqEjFxZs4lgsDkdDD7sXw6Z7nqBUN1QmC71c5205FzTX554Ut+ClYlORRj
I2lbM2o6KX4mu8Ez+kD1CFpXb1NSHTkDTVehQKfJqi0oNoL07XZZ3drsk3ywlZI+
qoo74mwbAKrXy8VyThGFf2IKprQqIefRqoSYtKa+qpFMgE/E2tj7DUyv22SDHNIQ
VdsGaYVJImP8Lb+IE8Vptv898l/NqHkcyQ6qNUNWFsRG5LCuj3+8/po+kjNHMK4C
3zivm49NTEi5PlsdfeyL0o+CgkVIobepMZYS5VLZXOY+JhLD4WixuxsvYXiTeN/8
TNT5FQmu35CnK85mvnXS0+QM0lu2U0jdv+aIPl4n8Vw6mrkYNvW7Q9a4tChh5+N7
9GqPPdUIQ9DkgMMnZ2OObSDZHU4rtxz9jH31nmGGCd9zdu7kFWUQkbgAHg2QajSk
lLzFJV4omjWw2nbCz/tmHoDVDJcSr0F30VI7+eb1N+zMIwLFRulTMkZmNWnWBgOZ
5JJ52qInP1kLNEkpo870ky3jm803jG6rL4vIenJH1p6nBMLVYytywUIJzWh75RPW
wpnN4g0OT8HfpmLbbHq+FE1R59EZvS7IA5mZrm/oHe001ozBcRrItDd9+fvoEYc8
sH/rR6aKPJkMQ4mmwKWhNybMbq9pp70EEwD5WPu/pq+snFg1lEwbKo9xNnMok3WL
D8XEavsYiX+cc1jWs//YkF4z4nOqqEE8QQzIvwZSu9LZIdVsxfbD5qBAWmfo3T32
reS9T1LUQvQ8P4Nn0OQM40KJ5z/UcozmzIFiNRaQg6rS8+u6mFKL2dc6CBnFtXmj
XX21qr2Vh/CEKLefMx4HjXA8qYwInVA//5y/9d9qGyLR/aoyyzBLEeUbF5yW3UEk
aax/TXBiYu4dI4a7gOCctnejGuhFreKre3aG4s/x+9npvClr8dGBBlA9n3YCBztL
D2AR/knR9Pz+XB0+5jJwVQOot4+Ov+jJ5B3WHt8KIMDGmxY6Ofw7YMIXtJxDAscJ
0IlCCmASIwyCe+94qWqEe7PuwrurjSWXESsKBA7FUl/Fp/z5w7y2OVFdFhAnOYvZ
ujo61RxQpHfBEXDQX8Xo7XOxiDTOEmpaCJF7p91x956HE5zCHIwY+JGEQUYnIko6
yfBKEZQ5FFtJTwRF0Kc1Q3o3zvSm8slSpt5YGi3F4cyIeCvPC5vovhVIx6lgcUBc
V9/FMKVFDcOZ79gxVPk9Qo5bFc9ZyOTKRwQu3kUSvajvvpXGUxxBar0R9edCEYp5
hSvWn1yw7tKsw00JxcPPleQbw/98156U2dP8vobuywlE4/o2N4IsJqiD7slD26k+
glq3SiSgWka6wY98IS6kmXZn3rTC/Ula8nlyGuy5/4j3JhiWrpFDqpMDpxKkMOA6
T118x9G/knPam7zML/dUsmOyyY7vl1q8TYWqvSLnJJTqn14XgzcUy/UTjsd1Y0kh
qcq8ajkD2MP8X0Dkxma326gk7l+9hqCMPN6REsolZw+Pj4vMxx15FRKu8w+uHLnx
C5d24w7+lf8e63wdOhm6La+rkqbkptWK/GB58x4jAibdDE+BL4+7M0K9dvDtsHLi
wnqTK7g1dgXCXWubBrzTiGZAA6VxtoLEV9C8eNO4or7n338vp9NWfeFMTr9hJTyb
8stabA+o+aANlLFKbEbzkE0z6zFRAkIzkiAjJh5otPX4lJ7DYTUaatn8dA9wVLRE
2U62Ho4ticbmLOpJl5XVVysexcKAiprjhbsrZONTJmolOzpxRKnhSdZjjfO5RnLF
tzosFeGpIQM3yXAWbMp7Jy4srPBWwViwcxdXxou299bO9PeWnCTSP7LHPiFOjHLR
xn5s8YqpJQynRqTHcBzimyT+jEFy7UbJcwJ/GDdhExOkpJ1OpfAuZCOkYZ2I6URJ
/WtR1TtfcKEQ9LwycPExU/tGm0Ko/YpqXaJkoP/VRtxOfaEezvEogIDq4CmIMc8x
dABKtoyr4A6QPHs6Bfvkwi7GMQImwmlwcvIwEXkcgIYwWP9jft6JpFL5ltB2+pk9
SFu1vxlio+nPEkQ8FUtwET3MSiknUpAtsJvc2sS+IoG5map83Ozzxf33ACXWfpNb
Gtd7hl3QHsB56GLktv9CqdlpRV7kV5tgfdEIDpQIjW7A6h9K1P5/pfxfAlrh8i7I
P0YXTI1UKjsk/SWzlygZ11seMkL+aLV3SDiFRTHcF7aDV/2lmSXDfkLX7zGXXPzl
oMbkMQ1yBg4r7JnDNcew7gd4A2oaFzuUj+rvGhL0Yx7Nr3errOP5wK5tbgFkf3er
P2+dXa0Qmgbgt/ifq6F//GobuA2WRsdoNszIzeU3/MrrPkcHejDsE7/Jql1NiN9+
q+U9jeQT3HfiPUbemFDrf6jYS4pJquRiK1l6MCo8ihu8RoBk73zv0TG6n9Bw66sP
HNrgftPUQNLEoL1s4FeCpLqOREL0hsE99Xg1Sb6kN6k6cyLJhN/2JuYGOmvt3doP
SnL9M2rldHqtkEZUOa8gHgCbIdCa26Zi6TSsIQrjPaoMddhhNwH7jYHJ16yhm+rQ
0AAMfDPS9QI1ZFZuZaUci1a4e+4ybtCQbMJP0yPcG0m3ZkUZXh5RCZgTYKAypLxu
0LmkbmBmW6erWis1p7arLDlZd7kpVSF41Q/MLbRxLIFiVgcTtvB1WmJJb4S4Q472
5UUo6eHQeca27OJYaVMCkA==
//pragma protect end_data_block
//pragma protect digest_block
STY3H8UslupYo7TM8iStEFD8ImA=
//pragma protect end_digest_block
//pragma protect end_protected
