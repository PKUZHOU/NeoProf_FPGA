// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ByYcGh9MnWzqjTrBvnCTh8Szpa+RnBcln1iAPIIowAWprtKMNKobGryzYi+w
zvih0YGdvw5rkyHuqA0HP0NEGSOuIXJU+uPx0i6qxp3Xm7Rxgyp/erPo/aF3
8F917HAqTc1yAD3LCKQHmV54O0SWxHDqSiwg+vsthnZeOuHcTxjwOC/by0ve
pHJ+qJPEIm1B+CzX8yJbX6Y0Km9pu9myBHzXNZ986filoxfzgRaDTo4EIl80
VutTTknryZ9N2av1yMtCBmtI/X6Ubx1fLO1HNYXiu0LgyIM3Egnnmp2GB9Xi
CDXJC/BtJFwMd16l7KKPjCaM3yD7Da+JnZMNJhyYAA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
NGxr/B/E3tR5aAV8oim7kHwaIK9357DG0gwyWpQ/ARK0KZdeGum1kPVncji9
jgqT9YXkIAjbY4U1MLINUS+NClk/5f2iAtcsI7hCgOX1gl5gnntexVkhufxx
a8wbF/fl8ZbIR/aLAubGigIFamwUqEaBUe/dx6wXBMfmktN189r9E9ngWJid
IH4ZC4HT00aCP7y/FYKEZ4hmfu6u8AcUCMpwVQSNqH3ZBQ/oaar9Z/phAuei
SEZDhBIp7+n1CtdcauRjW2pJBa+FpyuurLn6ZbEQnLxxYqd9XQ1WZmTe06KM
4hg3BSeAB56CZAi39QWO/8Huv2XHTzzYm8nkBH7eQw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
S3sXR2fNR0gLjjhSo4YxeNuZ7Lknao82fpdhxg4QvAVhsd+08G4Z7hOiouqo
XpbBkqvxbBiaGAN3X8es3by1ntOH01Qjx0gUVJSQ6s8H+j1NnOqJPBwroz7O
mhwrglog9y0GRA4OLylww3/H+0wVCSYLZ5jJ6d0XSRg8J5eFQPzemIrFge6l
RarilhB+9wSepiB5cgB7ip7Vg15By94T5tZD6UV6srIPbI/nWvPah0IHMOqX
Cwc9wxX5paqAx2Ri8e1Mu3sYMTZ1hgZcTqISEscwrDK7/avSaxMEBgB+bI97
ZlsH4X02cFEZUuxKxhpm8ZDxIhXc83USBj0OkOXR2A==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
VhqlIEQZ1ps1i+Uw/rT+Etj5IZP1uyfQgij4+yHMznUbC0CpVhbhOqC81cIO
YRPXQjxbZFAO60b0FyrcdBoVEmUU8ulVStfhZOJx2GMunOm8Jn2dn7caebEC
alY3r2vlqLA0483hezhXsz1PQDN9m4sGGoSMG/u0iG/UIaVdRHg=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
c3DqJz1A8JB/UPEw3XG7LCbHAVc9W1eoi/OCNd4Brr6lwSH6J7x3OwjInrG5
/RL1e2dJLRI8eUvbAZXXM00vY8JOe2SoXjNr0eO2ppOzQwDAyK1HAbIM/qy4
YGiR8EuLVWAXNIemQzYojOlJAEMIcX8ad48r8e/RqD5iogAjmlv1g4TePdoP
zEIueaPk5EBWjjOvajf1ejeFGxrJqaYKRAmlhNsQ/eB711sROnwJNDRvImKz
cNtom+Uq1ePYkYtLgO3RKKQ2Wr6kTGFFmA4J9JcHV98rR4438+aYZr5LCn28
/nATXxt0a9AuvO4Ki6IKdJeRmPCFuT/oJz7AurFwbRwfgwx07yYW4Hj+4/bv
06R1FTolyEhKqndIBMc1DtzuRwWTmDckLsjIppFLXhyQp8R+uNkGoUNX6Rm8
t2pP/r8FOsEn0T/8LdjNpQCGIUhID7PFOGijzvjQitxchjx1rGeQxiQT0r7Q
km5ggmv+VG+G+Q/ZI2/vMA2IQLVBkmse


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
W7qUNUdLoQlx/Jx6j6QuDQiWeO1VLtHI9gg6laFg7Jc5hDE5yv5yXjeiB3Zh
WHG1JFl5kMVRdKE/hJIwXOKn3V1pzQWw2DZl3omkK+TD7wm9MTpFI49V50m+
qWEO48ueUagCG8GSI3X1Qp1yIhmaXlo//wqH6JvzSMdn1C+Zhc0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
kKz+7yh2OeH9w+842jwOqA/4IB3Q1gMxg1ZhK9Wn6NeEQP8mvr7VNZm+7kUM
CRz/BpTRqEpbspJoD75ZDF58f2xK5lfNTTiz0B8p5VrFvJ/l8ewWN2DursHP
jyKYfRpNithK2C3N4cqNqtvNLae4f2Eqp6y6MN5QKzpypc9+NWw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 6768)
`pragma protect data_block
WQIgfTsCmyng2bF98nKH1ojaBkJ1Ky9oK726kyMQ3DwS3rYFI0dvKAYLKsB3
RwCr0ez90WyBRMRo4Ay0QYrRAW2vD3vkr4zgnC8uFdDeUIQ+4vgWi+NRxmSh
ZrzM+ngrEmOHcCEFGSxAkcFiDODLARAcXiyV6wMq9wkT3lCpYuaiFioGWXf/
pCuu2jHAqdHDD4RE5+zo2frNjVnbzkxOtgYwcMI6lFGg2FTIMZb8tq2KnIle
8sZ8m7gXhOyALA0GdWkPjdMO1vcW7B9B5cmUUPS2OVUiKG0uexHRzUcVoObn
MRA4rSrEHeemr71j/BuFLEGZ1evw8XJ7HfQlEChd+1kZSO0dl6ALAjzBDifh
b9WJuZGQcDnFp6WDYuKemOe2bxtO9ZeGo10CHbF+tK9/PbUqnrm1G9Wk0doH
iWwzJstCkPMytHiImKXPBzFGyiWsVB1c4DOyhR3WwZJ0br7aZbPxzAdh4Q1u
RaJvPgWd6MSS6VBLnkT0SI77kUkWmYgZ408+GmJ+31Pe+Ri6Dw/7fUgb4Nix
47KO4jQf8FLyZ8+cM/3CoOmtNgd+PTIvjjWYaAQgOrl+oHp6934XUDQHzKwz
JQqzW2q829pa7tZ7qFGXjRRPCQuBPQkim/RkNzTApDQiznovdAxTCWS23t/5
tZyfDQrGgkM/+y25wHGDFxdjyai4ayudT+pJW5+QGN65tmx6c1VeKHb5ORTi
dfsxdRcnck0X8JCAiptyljzlk1oOrgOkURXaikEYY8boC+ndI6SqssbbjZsN
mB8IUVjxlD4jhwZd3gF+s+EmVNyG5hPpvxqPs1I4zCmVF9jN7ByY7wn/mLXX
LwG08N0zDwqwZdHaBQUiCJAk6c40WKuIK/wcS4sbm0rKWK9EzGgvadJ5LFMQ
gtvesDFJbRJnqpszUReCzmr7XBZ/Nz+cF/YiMedfnBCNErZNKnTIOcVLqmfQ
sF50muOrZow1MNNe5zF6Jn10J+R3kHvjJOsQ0qx/WhwU+xapuEa11T80yrO5
B9uGHLcCWSfDxRm0hmxo1jJDotzbpDhTdQRwzsWa5zdy9Lw6yt8morfNXNoP
ZRSBu/wtnuqcd5Z1YotFPrbzagCWlQP0Emu+oE/5Gz59MKH59fRJm0YsJpR9
hA8vmR6g5hdlYujfBPtSOvCoakRWbQykbcykOC2ffK/mWDH7et4ZkasU/IWF
b2YUpblOnIbkGrb90NR8jyR0HogaVaoPuEALVAigLcSnqdobVbD38SRDEam3
9P8I/na2JLT0I9LLto/rHgg5vNVeBFrAk4imNAiVPfclIK9zabT3iH5oNu5F
+V0/RAamIFv+LO+XbfUkHPJRrjna3YxKENjsT91m4gjWfYjcjIh9m6zuHHBy
6Q614VNYdSiE9/2BJFaipfH3NiWhXCv7EMIbBf8PQ3QyjiI39F75O2DZoWIE
9Xk6svG3MVQlUm+21PmaCc1jBAE5OJJuqJC6Ma9Jgsr6ra+cQJOxb6FufnEM
SswXrMXq3jq0r7FDYeQT8G4lP0p26B0I8iSRdw4LxncI22NPdybqYi+zFYo+
s7FpCQLVBAnjtZDo6HALWnGIClfoylSGXhbCLbD83AM/qvrqa8QlDupU1GvQ
a6jq1JI6/6o0hnYa2Jq2r8EQ8dwYpFfx3fMGLj1o0iEFI4a5OW1iwX52GusA
PAtKy0nHxtX+Fbm/vV3QG/uouzKRt1t2a2KSFYXl77k80mhIbZUn1I9J4R+u
mSlvEzU+Qm/bfrivTNGJ0ExbAQouhOUGo25dRhX7XUMxBb3HOpduZ+J2CsKh
xbGDyDQWbNHovZPSRw4JSBVFcOmI/ZSnWsIcVE1wRiegUnwUKQSe9nPgYZhg
Qh+NQvvPJzrcAtyIgXZyZePojLHjat+4wLy2wL1qv51Ezoctp5L4ojXZr+d8
AatWvkovBZZd0CFx8gf174AgDEzqavoS6NC/a73ULtNWXcujGnyIzMHG/OLt
PzeI0MR0RiRPOgLbPyY5bwZQWD44NlWPJ5Ig+hHXlaBSOIRPyQkB3rreKH3G
5syZ0Qi3PqxXcwXyamWJKukNfd4TsAFosTBtRe2VKwQQZekr2ldQH0rjZyZW
Sruh1ffAFFh9MxAA4LR3kKbWRCVQwOjoW4I4s7rRIaOugOdZxFEo2Me/J+d8
OsUKxdS54iZXoPwGRyWv/ussB4jHITb6YlbYGnsr7qI9dIVUC7LVkPy9nYTl
byPk0R0Lvx0+n6jkbASJZjd+Y9j6krnrssKirh9PefQkLWGo063UBJtlTRbW
tH/MMQXTT9vy0mkh/aaefg9bsEpMgn4emu2o4FT41E+F2sEppbXfBjPs/qHy
wXeyk+zg48LkrrJRXRb5Vvhqa4ggceN4LFGM/Ft/SxOLClXD93WOC72ryZGP
vB6Dzd4Qlpbirzt+lv68JoOhAMkCLYXOiUXy334pQgU1ircKuXf8AyIIINoe
tDtIHeeiOukqQcAlb8NZs6fKxEe+M2f/7C+F9YgiFADd6nHvcNWo3Gou1Ut8
KdlZTO/jdcJSotWQf+mqycy6SdD4/Dl5A/cPzvVWu/2IyubrvPfURoeVakHa
2/av4UGlJhJgj9bZusMI+/pczt4SMFBZCfCh3jVoRpdpUqQ7hisou8KHd2/M
ZxIPD4rfAYGkt6qnwKvxwrRnElrkeMT709VVWXXRMQd8LPLo5Jf9Fwmtsyex
IWrPVcHHVSV5R33APS9wP4N/GcbbXozR60HlxnQSdrJVnxBt3Uo/TaJQx/g/
R3TwAME/2rfejBjMXFPls910tHLwNQnwvgDVAMcULkffIgTvGYA/5exfwjmC
roG2v3jyzPPxBFRlBbEfVTZASO02Wox4BEvln+jr9JHadgZ9n/iuT0Ln1cEf
PCOpa11jwo5xz+YZOsd+l5yOcoLnv8TYN5aB1iqMUFdct+hRrqbISggroIqb
heDRqnDYQf6/PNNNrj1+ivFm583uSh7zacd0efz+N/vmt5XzA3RCT3SHtXNO
PeOouammdP7M0UgMhE8QEmQDo8svYZc7CJKymookOK9VJu9mVu1Mpd0GanLH
tg609jkTsvgBUAcbK1UjyMihjLGm9eAII5iDGAaM/jkJKca9a+HjyLQgHh0V
T/GkvUksMP+l963G/LWdabUNPCMATVclL59hCWJFiKeuU2Ewc6rwVWthjj5n
6ex3dNoskq+73kJCbykMmEpH95Qk54sRH8mFL0qfKwIzeRjhd499p/WKz7Nw
vdiqMqRayJ3dXV5XJHQzIJYzfKohFudTXxeJe5Fhn0lS+TI63Q8TL/FttXUh
02vSPbHUGL5tzW8GHyEi658mXppSV0HUVLvXTLmY3xaLL5xTi9UX9OJJBE/a
AP8YWHKYm7riEleHmAF5won7l9hCyjyictqFb95k1zng+Yc0sOqtF1m7b3Lp
bD0tt+Sr3iiE2vQ9v6T5YcfWhcNKxA/dNOzra5W5pEJy2mFvNaYWtMYFg8jS
yRNIYKkq1yuJcrMCL+i5vDljAKvUdu5xsUOZIHqjkRZxtxObArT3NFsTWniv
Uo/ZQU+qGFfC0KxRPhO93au6FEkmeMqA/sGMoKyCzUam1X5L0jgP1s+0cFIw
1dGLEpZ9kOW7JmAWWflFQTF5qsWAdb3Lb/+py8oS/Crrf2zankNo16cFsS0B
9AS2EU3orZbjeJWPm95KHtb9AkTMHK8HX2EI2dk9jUIyTwLfl58/3Yay6lCD
E4JV5hKMCdCqcU8HKO0JZoHD27Uh/1ixxPTTA+mrXnDpK9qgkWDjk9UJ3aG/
W/KTJIwai9YJBFfyQPrERemC4pJmVM6RbZlIoJd6xOhN4ImdepgOBBMplfAv
oi5MrsFO4x0bCvQ8Rm+HLh/EUMTRfXOMfBho/rjw9tjLv5iUCMVYFk5KNfER
PRcxy17+wjwxxVaUpWBXx68xNrCMJsJWvSQrSFQXzn2qFispRGNSiUbCLu1U
J2SQMDhmNQX1aMXpikAyp5EahsGfaFQRc3HSfbHEWsQ5agBFfZLINdNlpSif
0YFe3YtkFUIrHuFhiQ+aShQWSaIxCgd9E5IJ2tJBALy3vgdP36sBMeQtno5r
El6SCzv8EXwJqQZsuqSFEg7q0hGchn4U3tb4qOkPRVVgTs8giPUj/IXvwB/K
8ieXybha+DxT2KzO/w0ifdTrzFPs6kCZ+SZfDXUSXMpmlBULfbZ7zjDAJEsP
z0bfB+QS5futv+Bu+OTFUo8SFYkxOlNBHeOIkE9ad2u+/7kMSHMAgEmq0Snd
RsWx4h75QUPpepFuCDG4fA00idnsm/VKwjm6zSLkObBRGUydXYskyu4mc6hk
4bnTfRee//KxsWoqRvMNmkOcHJFiRBfh1/E5jlwn5GfmqKj+sMeFhyCVyYaO
pF5y7trV0P2VsF7rmc2a+McUwt8gT/y7KEYLCy1VbdSZugVsw1xillxkzY6r
+KeolQoG0J49GCGtT+ynj8FzYWibg4UjUAWnvgSTdaqLEqPPiKSBupZHNKAb
xkPAH5gxxhNQ2u1RzvrnAsAU6AJYnCjpVMYFliRkhHrIX/IKlZmb90AG8uVe
PBaqOChECXKVOf9uRLsX5P7juzqIIwmpaYXrWfY+nCy+6pttN5W5zsVNA8AN
lbBw8cTJPbFbMIYlop+F/Qk/zq6GO8IaFlEiAXwESXBM7Z9yE+kZrsj+mh2G
A93dwIi4q4HBWE8ec7G5P5UPbsWFLixuy7PFv/JEA1NH2ky70ttf3nfyoJ5V
MFgK88qZEOh5yaA+WoRoYK1ga0M5FeYyXzjCGvH8Bng7KN3vNeO4XWxVYbQr
LZoHaarELy1UST9kdt34FGyR8VBVh8spR82p1jZHSdI9AjbR0valw1CWcFT+
7HdFaikiSV1Zw1frr+WVTBkZlwvHbmxl9Gd/CxR1FXEyxVwg1AVJfBgKdd/J
L4wq71g69auBNZCB8fSwzBaSlJCxGYcUbLy84OYad60BBvvsQHkXyLjFE4ob
m4ZS/SFB1/3IGI+oF0y4wnE7cWUlTaU9I+AbNbSjvXLVjFHe4DbDi01wJD+u
+RzUtevBUBtJIfh0NL4itKortjMoGBU7gUqEnxJSP01wwXuHSmIEL2tsbiSP
zZ+YTZYCyZbCNl4IjXdmbGxMtnKlFw0+2F53xe7Waa2o9rJGOfG1pNxZZJkq
gOhzOesFcwtKi0Fyrf806HrQOHrooirn+tk0EKwoNXSZtvrPKF22sk0fIGcp
6yulv/fCk7e9tyL2q6k42dRbbXOGA2BatuF/T5vxp3PHWiiXVsJs0PA9UF1S
cEPpKlY+ZlDNV89YhjS36JMYMLWfuAnP9HFopLADO3yc9s9KUqZfEaW7AgVV
kXgD7W2mWWeorbVBm4NYiuruLv1KDoYuj/l3+vwk5FFLepjZtW38nIYZDEvF
MKbI3pm0B669NxS2e1jwAV2h8PV3erFjn5aW3kdlpmt4CWP3+x2KU+s+zHFj
4RZcE5/SD4fTM+c/1gUXtWhmWlJlKEfm+am7CSxgBm3VTZ3M5hEBIa1XI1U8
MasM/7jD4WfpXCXvGrnNHxTeAL/KiVf6VOwOZgKx1Dy6CFYjQW1n/lj8U9U8
/l8oyn0j1fiEKLznSbcnRAni/km+mP7qDyFilNWDhCi9DXCgqS1MaOJvVwZQ
0d9AIuDkHZJCT1voG1QA/N8RWFtsydPQNr9l8ZwVLy4RWfg6nafgK77TcJsn
pt0DEF27S6FLZcC9xTgltVF84HYkF2WeyC0ehsHmORfN2NarYmGevmpHlPwq
wUdqgvTC3l8eSca/g/sc+KYlngTGxwEVDg2A2us8jzKFWA7WJIiQlxV1ParO
6e19/3yEDCzRf9pGju51LhX1FfL65dtkfXZBLIHbdEf0iBzzn4YT+lwmV80v
yluTbbl+bnTdiFD/ssSIkp8NjqZdO5Mwh4mwRfB8PqO/sVQJcFg3QkkcGmh0
OQYbONIieIkqSKNHI5zvwV95Csx6l14tw6RqSt9WQkMzMdhZ/7iCk31ddyV9
iZxlzysChYeX5kxtBjGj9kJyPKnfIsGHBuezTU8dca8eNNy1mTVRNvqRgCls
imw4Bn1UYFqegbgxmpM21W1K8uZUoiYgLVokTbqr6koanjwVQdWzp6A0s6l8
ePZWBXpZ5ZTSFYN2IR4rMpNFmBj/c4P99Dt7p4WmVlb35TPVVx/9gnCmhA6a
h1ULgp1CcydYZitnXJWHzMO4FeObqXihorjdH7/utPsMOpVxb6AxWDFMIGcY
WaFz0gpunJ8bgt719YGAXEjV9LjjCF9LOOwCQspFbX1488l1MuEhfe1hpuAm
RHbh6FvpOMo39dRW08bRDGQhSsmheVmgTZJWU6JQ5er9Ch1e2x8swjfwi8c3
vGyGfKWS99Zvv4T4GZHafA1CpC2Q37Uyp7c8n9ko9P14PmXcDJW8cQZQSi24
iFVf45rDubzwgCYcr02owj07ikQC8JsDLpjZ3w8K0Qw004pX66p5KCS+TCYx
nYiA16do9jxmJvAOXEkwDb3SNmzitCUvwYhvZ/qne473AAf9eYwbBGu2zIn1
LaTdSQv5r/mOABs/0CcV88bEclTsIFbkLKAnwkmGl2VsgB73X68FXOjSf+St
6WC2VuKmTZJ8gWQTgkExFCvDSR/S1CkdrSbzJ4Jqe3zcGHNrRd6OhdZ3w81P
YqYnEJseNrLf1QqfnHw9HG0tFPJYzn2i1UJG1+ox5pjPEMt+dACpjO1c5g4O
EqHPNlhqOo5VCVjwIkLlcR6lY6mz3gajJr5g7GUC0rTViVjw8IyXoGr7s2G6
blRx3XWdLQTcgmtqowCBGGyc3vMYFHmBVzScSfoDvp2A8dSndMtU5yOKxRWD
TklPc91kUZssc1ejKflKxrG2CZHvWZi9+iSfVieYbpzRUxgSxDX5CEto1q5+
kLriQhN4C2tINy2U6VpdEXKZFJ02zpzesaJDfVePq63cztjqSb0ujI579hy3
3fBNYk8gWzk4o/0gcryNmedcYEf/14QozCjCIuNXwSknlsk64jW3prcD079G
srZs9YyjltfwSnCukk0chxrEg8omMgXUfk24TZLaotHZTBvuXFUWaVIv6gGJ
OW0QTeKYNpVihcHzs5dFTF9GxPTBDIsZD++Dd/j0deNI71uPl4wIrbGcTCQF
6yeV9qR8gJFE+cb7DFN+vQfLtGVNYN5fWmlUS25KYhcICcD4L4sPXM9RMtnj
HSUJhX/jj6LFLjW3fzZs49NDFUM6O96d/6EOeQxEV2GSR/evqZ7KJ0yrYvY5
KmDLj+/7oZMiwTozPsyXiqUPvBgDLGcMD9JLDE+Xg/pY7YUfIQpv+oZw0GVH
Wq4fI+mu5f7HXX6jALMz3p13HKe5epDNNTnsi/wRlDEtLl/u4s8pL1ZNdeOq
B2ZAqlLF+zynF8hWYg1KEO8tTCrsnSOiTO+M1600puOO+Ng1YyU9HCp182oE
clrQQj0kpBW/bus3K7aZ6u5rsglm/lOPjS3olLlwie+XYQC/MogxpZkJrDbY
vPCM8070mFjyhRy2fzjVJlAw86hiWc14ED9FlcI0F0ngqvo7gXtuwWvgS0WU
3GuSMovqdP81Gmo/GdQhSEeM7GAuWeWLbMf7KxhVGBApe1cMY6MeYjyL+6K+
WXSpIMTi2odXoOCFbGhz9iq478YLzISFRCYYOozfyiQ59Gj90R2wtLqm1D0C
Rj36NxoY/hHZy/20ZDoBGpnwZGkiDcbrTcsuWmXLrO6kAy9I0UIPHfU4ZX/k
wsUcHE5/FWnWgL6qkQR1jjXkHsP7ISZPlvc2gjAersFt26pWn7T3w24BEJEb
LR5jgXRZeJtYwj6CTYxZQBbmj6OIy6BIHZoA5Kb9HDVABjUrgiyYRhjuKbEr
Zlygz2M8ex4CNtcY7zGmXydCYvF7EGTPEl8STK4W0eLGz7u36RS4QQE8QZrc
WkSBuTz46m9DHKxFVInpz/7xNCnq7Zix2QcAY5VBHc0cCaA+wqa+fdfmgPmU
gBYgW4pD5FkqfoZpWyDg32932pqBLWSqkq3xTf3XBnlmaUVYx5GwHScpQEue
jnfbZ/z2PQKjEWmVjPnMJ7/HvaUy89KJZABvLZ0+cMtAqX0fbqwiiI7sk15G
s1CxAY2OVpgnhYhDI5lS5n9DXBFxyOINaRoWvpsFvsUH8J7UQq3/cyV9vx2j
GoH3iBrxNVtfCAJQ+/VcefdQU9C1D6r6z/Q9yE2QVdBrJ2jbecuArFg0FcSQ
9C9yjZfRuX0JJlp61hiZeFK9Fm++9GECGkhcafOCMNvaizCjr5dJw9mgYxh5
6U0jPYmKe5lPiEEwbF9YgkWQkw6duv+ABULIOtbg6piVV4dBu03pZuxk6SXZ
qVTqFXVNf1yy0Zgxt+vvFBB6vohT3/o2cmtYHOsykQgdtXRplDTyedBfyoKE
HkV2FIh37KJ7jVuSfOPHBqIJqkCMWmKEFLLviUTBsjcNBsyGhfyMXA9FBcAA
R3/OL+NvgiFrBMFz1VG96Jl2VHxP8fhjuzHVSkFnLTSZGETC4yL9Sh/okV8E
nmtEsw3kp1IAb3QiIM+FapLjCMcnolKzn5Gkf8B4xXZJ5ZJQUmHx0uo5T9O8
S8nsBktJPsl+mH4Ifq5XVRoaLnSm+pIzYZzAZ5EU7vJ9bOtz516gIWYpKbz+
J/q4HLU5D5mPRbs5l4BDukieQd1TdH6iH/uQwfXXCLl6J7oujJCuEPwNAqQ4
JU4toH7ijMtf0U77mEqbRDGYTbUWQuQVaGsepnsFRJm1P/v0X8BljTmdAp9N
p1KKj/NSJXERcrnCKrJzgdn+0uniEFmeI/YR8tPJcgpuxG/g7PCGEL4onZgV
+lAkUu/JEaaHRr2D5+8H16cxE7o1QFgzx3JZNFo8uSDzXVjFyPjHbriFnXQy
HpR5c5ywycWEzzvdShjgIPd9NefWT9PA5K73z8h+77IR9t0DM1mQKHAsiYNm
DVZ240udBXN1mzFMIG4LQfqX9xcoNqoLjUy58Qjoh9CMgn1Y9xCa9a9BMFJX
KDFbCjXeU+fb5d0EZMHGNgpw

`pragma protect end_protected
